--  Module : ldpc_encoder_pkg.vhd
--
--  Description :
--    This package defines constants and types used by the low-density parity
--  check (LDPC) encoder.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ldpc_encoder_pkg_1k_23 is

  -- constants
  constant C_ASM_LENGTH : natural := 64;     -- attached sync marker length
  constant C_LC_k       : natural := 1024;    -- k = information block size
  constant C_UC_K       : natural := 4;       -- rate = K/(K+2)

                                              -- n = code block size
  constant C_LC_n       : natural := (C_LC_k * (C_UC_K + 2)) / C_UC_K;
                                              -- M = submatrix size
  constant C_UC_M       : natural := C_LC_k / C_UC_K;
                                              -- m = circulant size
  constant C_LC_m       : natural := C_UC_M / 4;

  constant C_SHIFT_REGS : natural := 2 * C_UC_M / C_LC_m;
  constant C_CIRC_ROWS  : natural := C_LC_k / C_LC_m;

  --subtype asm_t is std_logic_vector(0 to C_ASM_LENGTH - 1);

  -- hard-coded attached sync marker for length = 256
  --constant C_ASM : asm_t :=
  --(
  --  x"FCB88938D8D76A4F_FCB88938D8D76A4F_034776C7272895B0_FCB88938D8D76A4F"
  --);

  subtype circulant_row_t is std_logic_vector(0 to C_SHIFT_REGS * C_LC_m - 1);
  type circulant_matrix_t is array (0 to C_CIRC_ROWS - 1) of circulant_row_t;

  -- hard-coded generator matrix for (n, k) = (1536, 1024) code
  constant C_G : circulant_matrix_t :=
  (
    "01010001001000110110011110000001011110000001110101000001011010101011000011001000010000011001111110100010000101010101100110101000010111110001010011100001111001001101100010000111001001101111000101110110001011110110111011010110110011110011001011110000011011011000101010111111110110010111000111100001011110100000101111101001101001011101000101000111011101000001101101101001100011010001010000101010010110001010101100110000111000101011110000110010110100111001111100100101000111111011110001011101101110001100011101101000",
    "11010111001111000010000001011011101111101011001000110001110010111100101010110101111011111111010110110010110001110110110001110001111110100111000011111010110101001000100000101000001101010101111101101000110001100001001110001111101001010101001001001010011000011011101100100000000000110001110101111010101010001111111001101001010000110010101011011110010001000110111101001001110011100010011101011110010111011011100111001100110011101011110100010011001001101110100001111000001010110001101100000001111100101010101110100010",
    "01000111010010001110100101010001001110110100000100010100011110100001011110110001111110111011011110001011010011111001000101001100001010000001111101010110100000001011101001010110110111100101000001110100101100001111101100001000000101111110001100111110001010111101110100010110011011001111101101110111010010110101100101011001101011000111111111011100111010100100111111101100101101011011111011101101011101000111110010000001101101010100000011010110011010101011001010100110101000100000001110011010100001111001011001111111",
    "01000111100000001101110010110010110111000101110010111111101011100101010110111100100011111111100001001110110010001001010001000000111001011101010000010001001000100011111100001001100101111001111111011101110111101001110110010100000010100001010110101000000000010001100101000000011001000110001110011101001001010100100101101001000110111110001100101101110111001000001010011011000000000011001000010011001001100101000101011010001000101110111010001000101000100000111011000110011001001101110100101101011100000001100010010001",
    "01101001011101001000110111111110011000110111001011110010111011110001010111110011101100001101010000000000101011001101011010001010110011110100000101000100110011100001111111100010010110000001110001111001101100011010010101011011101001011001111001010100101011100110010110100010101101000111111011101011101010110000110011110011001001001101110110000111010101110010110010110000111101110001110111110010010010101011111100010101010110010000111101001101101001101001110000111011101011100101000110010110100111000110010100000010",
    "11010011101001110001010010110110000010110010001001111000100110110011110111110101010100000100110110000000111101010100110001011010100111010111010111001111000101000110010100000011000100100001000100001001100000110100101000001100100111110110010110011100100110011011100100100100000110111101111101110110111010110011011110001000011011111001001001110010010100011100100001101101111011001111000100111001000010111110100111110101101110111011100100111101000001011100011011110100001101011011111110100001111111111001011010110110",
    "00100010001001000110000110110110010110001101110000111110100100011011000000011101111100101010001011101010110100101101101010100110010101010111001011101110011000100111100011110110111101100011101000010111101101100011110010110010111111011010001110111001011111111011001000110011101110110010010110011111001111011000001111110111111101100100011101100000110001110111010010011000100100111000010001000110111101010111111000000011111101010101101100011100000010110101101011001000101001101100111010100000010101000110011011000001",
    "10101110100010000010010101010010000111111000010111001010001100010011011110111110111011010111010010110101001100000011010000000111011101010001111111001001101000010101111111001110111001001000011010010011111100001111011010011011110100000100111001110010101001001100000011101011111110100011111101001001110111110100110110111011000000111110010100101101100000010101110111001001100110100001110110011000111111101000101111110000000110111011001011001101011011010000000010011100010100101001000011011000000110100001100011110110",
    "01001111111110111010110110001000010101000101110010101010100101010000110001110100011001011001111110100100100000101000110010100011011000001100111001010110111000110010110110100010100010110010111000101001100111010100101111111000001011111110010101001011100000010101000100000100011110111110001110110011101011100100111101001011111100111010110010010101011110001011100101000111011110100100110000110111001100001111100000011111100100100111011001111110000100010000010011101000010011101100001110100011101011010001111100011001",
    "00101101000011100000110010101011100011101101110100100001100001011100111011111011111010001111001011110101001110000101001000101010100100101101101011101101110000100010110001000100000110001001001110111100101110011001100100010101011110110011010101100001100111010000011010011001010100011011111110111001000010100000100011100001010101001100011111100010011100001100101110100001011001010110111001111111101110111011100000000110101101101010000001101111101100110111001000100100100101000011101100011100001110100101011100100011",
    "00011011101010100001010001110101001011101111110011101011110000001100111111110000100010010100100101110101010101010111011000100011111110101001010110010000100011011100001111110011010011010100100011111110110010100110010100001001100110011010001001101110100100010010010001010100001100111110101110111110100111001101101000010011010101110111000111101010111111111001101100000010110110001111110010111100111010111100101001010111001111010011011101110101110010000001111001000110111100101011100101010001110100001110101010101011",
    "00110010100101000010111101111111010001110100001111011101111101001000111110100010111101100000101011010110001000001001010111101111100000001110010010100111001101101011010111100001101000111010001100000001000110010000011000101000011100101101101011101101111101001110011110000000000001101001010110001100110110011001111110010101110100100000011000100101000001010111110010011001110001111010001110110101011010010111001101101101111000100001011001110110000100000000111000011100011000011000001110101101111100001001111111010000",
    "11100101110001001001001011011011101101001000101100110001100110101110001011011000001110101101111011111110101110111101111011111110101010101001010001001110111010100101001111000111011111011011001100001111101010101000010111011001110000010011101100011111011100111000101011001110110101010111111100111011111001001110100000000111001100111100101101110010011000100111011000100100111101000010011010100000110001101110011001101001101101011100011101001001100000001010101110111010111011111110101000101101001110110110100110101010",
    "11111000001101100110110111011010111001010110101001101101110111001111110111101101010101011000001011110100111010100110010100100101010011001001011000101000001001111000111011010001011100000011011001101110011100010001101101101101001000001010011001111001011001100011101100101000101111011111000000000100110000100001101110010011000110111100001101111011011100110000111111111100000101111000011001011101001000001100100000011101001101000101111111100100101110010001110100010100101001010110011000111101001101101001101010010011",
    "01011110101111010100101111010011100110110010001000010111110100000101011010000011001110111110000111001101110110111010011010111100101100101000100000010110100110110100111000111011101101110010011011000010111011010010100011111011111111000011100101011101000111110000001101011011001100001100011010001111100110100110101101101111010100111001100000110110101001101110010101101010011110110001011011001110101100010101001001011100011010101101101101100101101001010101111101110001011101010100101010100100010110001011000100011010",
    "00001101101110011101000110000000101100100001110000001011000100110100000101111101100001101100010110011101111100110011111001001001000110000011101010001111011011000100010011011010111110100010010001001110001000100100110000011000000011000001111100001011010001011100100100111100110110011100101000100011011001011000010101010101011111011101111011000101111010010100010100011010110101010001100110110001001000101100011100101010011000010111011111101110100110010001001010010000101101001100011010110000000001111101100101110011"
	);
  
  -- functions


end ldpc_encoder_pkg_1k_23;
