`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nFeCAmfGYh679FNL8x3jS3knawN5tfsSDW4InIdQZKBRzN4kSVkztq12/tMe1NyjxAi0cMi1p1mf
v6YsF7gSNg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nLvd2l9aDcTJcRr7PlbIbTAdTlqSll7rKgX3KRhTm6DJ6LKnYLgujWQn6ykfJMZcvIdD2hQjETEl
AVztkXcemle01ooF9vTwBqEgni3MUKzB3M3gislQcAk8dn7agiNAvn9Q2m3tmAUg8FcsXPvBO5o7
zc2EBMZovl2F7DKN8fs=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TJiYU63EGsOQzcVki8Bdr9VkW2GiYuYjy8cb5Z9/XG8LgsGJYrBmLZ2ERU0Z/ii01CLvlE1YydJn
WIDOCgh/1WFJYRL1ZWB7ohWbB1ugPLKV6HJgXOpuDQoJ0rQ304b5xBjSiLH4X+LZbHURDJ7ORm80
EFq7SNptkst73RTgLss=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fx0xQjMTeVb9mxjL6AhaMVwdj/PIeQwJN/xbL+GV7FQZ9+GRX6zMNlSaQ+s5iG23Lve6Wlz7+6jy
3JExpduc7cT4EK8HgvvuFvM9tBzkfzyXFid4kRz1yyfZ+22KyEzv5nC+jGKhBwdyJNTpZI3nBpBT
YlCbwT/wPFwnbooZqUjpksnu+YIODAUJzuu65eAi1fVwQVd7gEjv5v5TvZJi7pKcrK1ZXEadock4
fqehxkNd6+EzbUcfbXjgplHoevtQDecguFi8/Mwa08S4rFQCHEYRwF7ppgui6vwEZdLOlV0xwkTM
mTnDaR5c9k2cM6UiOolTWhwgxnMhk6bv6k1PfQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jXzUp6BpOygpeAJ8nt5CMi66bQLf3O4FAxzNCP69YWp2qZTZKkN9Js5pUdYjEyq6+T+hvf3Mcsm9
nhmM2NHgCvzt/Ua2sR3CfeS4HmlbUdnhyhBp2sta4UIVATLo0zBFA+I1GVZxCk7QB57WoTaOsVUC
PbPyAXclgp1VhJru0gjc2pDQa/fpVpchYRrm3ofLqy9j0xrV+SWGpQ58OpjhYkUlrc4CJ2UwT9eh
cr7rW4qg5+3IG/og/qjJWObQPgMuXYPtUSSA+xTtAWAvYzTRkirupyuJTtHfrZQ+vLfxPyqmXXUh
EMr2dTZM8Ufm4fJtapsCekBOiCy/LFW6zWUUaQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ir+GtoRS/s2W9kPfZ7WHJXdlfnyH2nh/Z5PLPgYkiPBMa1f/xwfEqMlF9oi3mKWj5qvsTMIuL8Fw
4jIMwjxDs0vpjprQ/Cs2x505GOF/dlCpTBARO1ObdA3UH4Pe0q2oJZLBBHdCJVxqytG08aSsgO44
9F30J+4EcZeFmiSfP3YyD72W1NtIqzXS3jeP/H8Cjr2wzBxNn7Srksj6LVHHFLlJI9kYqqU/I7e8
3Qnb91E0H13AsPi1J+d1p9CxhEzKdeCMq7m4kioswmioKsqbAao6cQdaKKbjyPutVjpZmS0Z50Go
B7ERgW2xb6/18GYTGqr5Mt+lpbXxYZT2Y9k/aw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175296)
`protect data_block
2+Vba9gwH83zJiZjFJBuA5HaFMhTYXjUmexUeoMDTNZmk4GVmlWUo6zhRads9CWlSjWUP3gu3AkE
RXYysiglNrL/DAgsBb1E2iO/Z3cD6XeCJwY1Y7TukYBusgepIdPPp5xmh4Q8qie49ARISCffcgUL
LNefYruiIoF/d/hZ2PrtYdWvoipEO67xEQdSXdoYUsEUBgz4ucPMfknHwBZdqk5HGrynlLoFyf8F
C7z3EsH86ICtgwVov1vDrvNZavfVJSEU677b1x0x5DZB6+YCLFEYbe6jA5OYFOyamF4I0sFfeKyU
taJota3yf9/aKZNYyQBr+6rx7XaKRu07oey/NesVgaYnCqGt9SsUx86I9rKnZfMCp3PK2urC6s32
z70+otB+xVTP60rK/vw5asOivnhs6vZhLJqqiPKQlNXuz1EVd2IiMFDRpEkZTRq42BhKD+boSMQe
76hkLltlp0D/q5JVfBTjvtY8zKigFG4bBR4tp8wjNGJPp91tyUcusvi3tVuDhP9cXHKFaRUnn3c5
JWLcm7doD/bee5A4fJTrZuzUAMkWE0WgqpXRQd9PGmbF+4MvbqQSncdIvUmYJxVAdhPvxgqJWF2x
wJEq9lEds7D87ijDmubO/CfHNc4pfVxfHNg/1MPNaVDBDf8S8Kmc6FF4FeySPi/0KTFYE9PR+wF0
kbKiZYNYst2+AaSQ/qiw1Q3cwPaCQC1a761l1H2/xoRMhKL7HKeXjFkDYfhJcxYwt8derlQqgYts
+T95I5KYXCLHZnEqBz+o3AsgLrOkHoUw6EaO8qaPsR+6n1C3y4kDQM1PyovjnVZjrN5WqagmxAPz
7Oh35fqN5ny8Tvh9YgGXt/Rzu09fGH5RdbAB6q5LPb2aW3WAtK+uUEq8fYrewfTKbT+JC8OZzPTY
SihrVORi++aXXSvqNfpYehftQxSgJweRjtM8xWgN0jhlber9vfVsF2/srXVIhPFZJM0kAqrZuVC6
gOAOX7Hyu+BZevOMTKf23R6Y0WQzOuVnz7mlXO/TK3vy4S+qcjDxm3ExD5uH1P5E9gx1CfSTKhQx
HprHOM4/pPNob6uJ+JOjbo+YKEqeK5X+m96wrMZicxZT69wH+78Qi+CFYiamnOXbLJFLLfZb0B/o
5I1iLVlo+pAjc0I4wGHDIgrPKx2DSoaUqC5058zrlqbrLdg/5jbus5cgBnpCEIuyy2BlvxUa9w0C
CzF99Oa4DK2dBFzqF09liCXO41XAwlakutzA1chtBaygNFbqgU4OeKABJkNDe3tpxL2fj+Gmg/v8
a7ixjAmxvgPVQfDihf9pFGu/TsIWGcZ0imS38ho3XbpsYPKWWMt/4PzxUEBgJXWHPSUyKPIgQGTa
o2qI3XfNxzxGz3r+48agN6BTyfojsArwnm+o3DwMLqramuNQR6T+SCdRwaepvvyKFimdF54a/ypL
bJqeIZbZ6tX81G0HZgKfBFWTZaTsXzqOU6nKW1EC6u7USmh8uUL8c79QEZEmysKRqcbqR6+WomSC
gTgxvm9ee5UymKB6X/IH0JARzkFc+Qa4qictNm9C+P4ZZ3NccKG9nFGxEgG0G7t9bMzE9MLfTlIT
kJZ4SMO8ZQw8RgBJ/Sct7+xIqaZVRc7jnS0ln/KNqLGjerTSovfcBcDlTyHqXADSsyXTvI/NA3M9
Uc2XA7LtiNixk4tH1yscq/bxnX0xN4e0JQP8QdNtlGpVwSeUb9MYwwllb6SHQQYcQPboSr7B7ubb
OOQ1RRmOzWjL3hDl9XSexuWtngs3DrYelfaLqZRS1tPOghEZuRQKNpMtLBFLrKHBCO33zOaQ9Lru
mHwsTW8xhnVq2Zp33DNy53gI9tJf0/bQuHyiVfrQ2IbJ+hl2Is6QGjmeboclb7ccDKLEejnb0FKz
DkVhNuS5VhatxkFf6WLv2PoiyNn6Xd+bvXZuMTe2pzdsW994cU25i7/wk5oa/Kf8/YlPPjPHMy+5
3qHhytI+/Vhz6R5+FYjwUDCYE3Jemz/pBd8UYEmYjQ0MqLTOFI9pFp99ytPWX/HBE7bpGm8BZ+mi
6noGwYMAVXyhOQz+dY7Bb5JsoxltRc5IZaU4PuOVhfZk+KC80BXWWWOPO3lqkw7fAU1zEwhSFsE9
q/6fGqNansw0fKA6pHFXrlTnVMIlKn74NEaEusE4uifAqA6PS6tvWBKWp+yQuhhmFN2qkwHN6BUw
zbsKU7SWJA8H2z4QzX1u5BeHYbsc4mGJTn2k6XDn9gw4I9Adzp5CW6fHWvgOWTCHCIFIPQ90xUEG
XfDKCOtcls3OdBjfDkAjieFvXyNqJsPcOT3AzhSEgTF0dnprpmpUcoS6v3My5DZXs1fk4T5xuBOs
GDZH0vPJMg6iQMF9cJxoR5LH6z8TUfiM1H5SkUWDTiOki3fRpOvRkrjS+7ebdzEwf67gtAG+D3T9
/uG8lQuaenIEiu6+rOg5VPeKti/KODDtBlogGnwKYgMU24pOmTZI8ZHFei05ORxvp8tz+x7b0H5E
jqM9kjGnxBCbe+7reTIxoYodecxJ9A1XyFQjJwyoEGqL3xljNIxYo85xepZc/QEucwtTOcNqbJ9B
jtanAvHuUfkNnr8lY4/ZEV/T3p16zqWA3mqgpXsKPAXnS4eP85ePbsC//s1KYkwQT1JHnXxekAU7
8jLK8+0Rg2IPBJ7Tt4ZxqUcfShr+0F5lOp3kz3PqSo3iVIl7q5fNgT1zAB3YnDcmIHl0hUcAY6F2
pC8SHjNGr++YpKSOZlA2GBQjEZbcGz/cLeKHeYBBMbzwZy+HV2c03abVIH6v7znQkKycYxupzwSs
PFovfvebtjYb3HWBIKwOHpG47BRq6JGQu6rw42DsloWl94zL34Dl+UA84UmUnRRXw5eY4eLJmtre
eAOkwzfaKZ8mYoRU+RtgngW/Mtsyu/qR/1+b/7ywvjfCsYumnZ1iVPLK2EAwqGG6AMjC2dAZJ2nd
H9XUxR3M8BcpcuatfuTTpcX+hvKRRIldjJOdXE3Imp9BuJjvhgAknU0ix2EwXFVLJuM1Kbp/Lc1q
v7soneWlwishfZoKoHd52oYkXd8G4P9KMttSnInOZeXKxn1/wd+xZl3hhYJR5Uu5/smqfBg0ONb9
mviU/puCnZutNTm5bFxAP76r4Cg0tIEZC0bqe/K7+KJzvQDldso17axpBUb361q+2H0Yb6tY/zqn
uixi7Mvj75Y77r39ODsFF8s9jqflGahLJAP98ZoYukOEknUoTKutHJ2TnBa45BrCao6Avf6cgXkW
c/r5ZZTJNcX5NK3S0ZaRtEu8dq5JPhfji1jhUsnhy51WirIuhIps2N3mIMT1XlzfC2qR0JMeJC/x
92j8GmC+/i9dxzPm3G5rRAvkUWvCyb1yKk5XUrrEQquPz9slQVWkiBQlp4oKpkrHOZbmOkYbSBdB
wD8iYVEFmogCAck08LKz6bDfgx5Dk6co83dcZ4jJ/m4cEec99uhyCo+eCem9E3x7Jsv/Iptt20A1
yaZtOzQR84Cptxvnwey0DF0TrG2B7ZyJQRAgtDQSI/xoWKGh9t2r0KJ9MqpCebGiIH+VpkF3SG8B
VJJ6S7fDDnpX/w2M4PVpa78xp9TOEGJMhZz7aON50DzczVEanEj5Y15Mrnzu3HAbQ0WPHB8a5zJs
fWWg+BDhVzAo0OlSrbSE9rcULmGRzB4xX3F9ntaN4tORSX2RVlmx7a+S3XRhYq0gzVQtoPK3xU58
NfVuhyfefI2rVEArKbK/bF0IgvUhBnwXVw9tcuT3qi2tkXfhMaKPlNBTckM7/P+Mfk5aC8MYsj/P
aQe4jOLYcDFA0EeE6TITXRb+uN9mfVO0COWuVdaUB5mg+4bAkNrR0fQ/sCrE1lzlelwzuhth582U
MKVL1zQcM7Jimvf8FlgKPQpZdoBIvCBTgZRUbqskINbA4a6SP6OgmhIl4dgSyaUU/jmaXIN0XXYo
kXjBHWESsT/BI9uq4wf55pdyrPm/uYYbA7qXqaIQujAzfJknv2N0fzGrJj3LrZxvmAIJQtz+uLbu
cjPTZp2P2vWJmcvUrp88CVk7qukr2np3ryMv4REBuJuM2IjGNc5S9VBMvoYturMKhyGyWV6qign8
mdHEaRftxJpHnY/AfRgYRcIpt/3Zo394C6mr2EThZOVMSFDDh0ykuLfTuz5c9PZ79O/f3W7BPE/3
+qbhpQztepWdJBQA0piArDq3a0h91G6aulXO3Cpc7pNzPmGxG88jnTpNZVt3PRIJTHUojMY3GKcR
QWQOdw4hhkrbXyEqXZiltrTFo1qLD+v4XJ1dlYgkheU3r1OP1nAJ9LaFXWUSbz0NH4BmB+2AvIUp
ukitv0609QiYj+X0DKAHNqvqtIkdsQk8LLN+arB7yOOXFtL9I1wjCLstTvw+kHlVq1sx84Q3uZMo
EZsK498bTPn60Pa5AUCgN/nUqjeFlM/2YL2N4/WY10piE3fE9DUeqpqfqq1jqmM0ni4hno9I5Xor
1RKFnePDUimwEey6huKA9jC+eAipsDOdRirpWpRLP6NndKrYHxVrKFCd/bgbPo8UBxa79dWqdFee
8PBKqKLVpNqDxH+nW9mAu9+ofX1ZWz8wrymc0hdJGbk5HlP3GbZWuUDwhem0y8vj0Cs0kYjpITOs
nx4Yw1eYCcSBsHTCgRjznxqMi/vhpAPz/M8/DOy9kkXVTjm0OMeWzWePc7WrK8Is50MhwHNVoQRT
qnmH4jEDS00xV7RmhHVzzxDyFluIG+9/J3vvctyi50a89Rld3xsciukekxBsAQYhpGVCo1PtNLcB
itaaw3KjHZ1k4jkHsgG4enJH664VnUeJ2apiUGVs1bZpXwJtZ+uvqn939vSvrNU1KXeyL5NNRyyT
Mm2+NzS4l/MvJR0gZKqVg3RfdSVzHAXl+P73ckSFQuDt1T8ijvBZABHWM0LuizzWjYD4Uie2tgel
D4vvpePLfWI9/mh8DBREaqltI3lZotee+/kllUeImErSMzS4P/ntdG0M6JvFC7VrTN/apoxw6FfY
SYA0dYaPVGhOyIuqTcoC16v0BFYWTQ6LknW36hzNJGUy1pJ9semx/114ufD5ukfujZqFiZSWC1qF
fP8Bk6oX/EOTz0Ck2LZN8786snkDoRRLLNbfVkI9TWgXyYbOARcgJSVVUDbuOO9NvO7xk+AilgGb
g89lhO84caBdO+1H7jF5OsYcJBE2oxQ9jj1vokjIhH5uDxQwYH+UzJenPjuVa4suED76wKyKizyY
fSgnNDDP2klConyratRLI0b9R8DZy31extE1gzuu05IqMYwPf3i4MoWe3Iw2+xdhOP+vJMTEcI2P
XmoMyuZRlWPPTV/5pCy0DgiYVEkMZr0u/mLMZCbuKsLOsbgW6yZVHnGWr8kr1PJwTpvvxj/CKDVj
ttS0tSvHVX6WxfQt5/hvwrhL0wUN02rRZfHRlBnAD7f00YpBngjP+Ua7MqtIlZuorulU0picXb6F
NQNrMogYb8b/HA0TaxfWst3kjSGYPXUA/qbo8BfzEroQk05ExMWLMcMTUkrilDZFP6KMVEqxb90z
K3452bQpozmFPYVbSy74N3FBNDqviYNjca/kg376IQnS7L6etd/fud/MP9L7QJN034hjrcEJ5Aun
RePkqXm2xgQM+k4CnphsiQFgOGtzidPYRBaHD+aNSfenJsOinBPdX/C7H7v7UCb5DRnWDR1TZQfI
DnRk6m+a9VSsr+khpBlU9DlWgRldo+zHBPRxevqq261ojsIQW1Suwe/WMUbbTVJKB1NPZcldS0sx
ydqMqasRDlBr+JkqGQq7ZnaT88oCYQ5fBwhHtGb+KMvch5RdW6LzRJdd2LqhWPkXHkNkt7S5C5Xy
TnpBLFaS1lg/YKD1ThvTJqWt/tHPUhYEVh8uRHKBtqll/yvHIqDyiq5Vs+gMKoV05WBJAMzZ8vx7
UAxAt0T0Dd9TrC22mPTMebx/qha9tsepcC1RqHdmeDatnWNiyIVboDlrYKZc6Ln5RdJh0idKa93T
5eZ2l5BqkmRhO8iMaO5kDripiko/Y710y/KRBHtk+ZOHUMb1a03f5wOyJVp0+26rTJGv+pv0/DzA
uoSc90r+lRu+wx2rGrUG9SGLksBrYtRZJ9c+cSF2bd0rc0EkzxENXI8D0OswiAm7Pcs6SVCyxGpP
/0nBlAafvjal/yqaDry4ClJtLha+0vA8iQlqZ6KdTaFgYnUT1NR9wTZSslAyTZV/IByRM2hVd+rj
dhTlN3cmeCwrblplSN4mDHKjGuGexKBSef+aBwpHlE4vPH3zYMX2SDcsLrD4doI8wepUlWoYct4L
owW1kTey+lQI1Pe6MzvbeZ788fSzYArk6hgcfYUFsNYZ0YrjMTsa3V9yLXfiuYqRfV97cip3Anfh
8A8J019r1Bsppp9FJ77+ClcDWDJBLuBX24fZvYStDrBZMIqpkxm1QxzvtLwJCsB6VO70oDpz6OnK
4QEP53cP6eLVuJdD2Lt/OUablZu7D+m9gvrGIb/7CSqK1L690aBaHlI/X9q0V7GuUWN5t+wMIH6j
jK3Rmx/JqlmOANeU5rDNI2k7yuAXrsCYsVU3caYH/1Hlav3fRJEEi0F5Wp+bRRvNZ6fP4tCYCYiv
1VY6xNphP3Qfu6v48HDCCqaOxi1UXCT0hxdsZyMo6i4c+ELny6vI8Dujr54BuqfXMWWFHxJc4wuN
aHUnWUG2WMOmBimQlMkduLxYh08r19+FbuVXDq8HAvj7oPFlcb/IMSsfq+MOydCaXpL6PnVyNd5U
iBvTOxguyWtBiAHnNnllIqGd9tep4tjV9yRSKFAjUiWGCROFr7O6YSEd3BLHymBhuuswJx/Y0dfJ
y5anVn1z3iF6f3VhrX1hEOCiSfczxOqJoNS53XMfd0ql9ymmpRCxaQmfk7KlVSRKqREukV+Ak1Up
XPi0eXwG/xzm/yZCxTN5e9hHcTgNAp0Jt9xtPhRxNeT2Imi1L/oyIN9C+fxOW6M9uiRnc8Gd7cn6
N6a91lZo49DLHGY4S7claHvV91LUxa5weyqpGZG+I3OAwxKQ41Rnvr1WqqSor5ARqCRgvgldp3yX
sHJopMPeag0i1qgpa7ifOjNAUs2L6QCVoj7W+bko2F2MxSHZiWUy6wo7bLmMd/FIhw1NooKOJ27I
1YKcPCf1N1wTqOoH1lGGGzNjpMDE5DVuUGT2OxLtuXT6V5GD17s8C9vy3FERAEi2m535kz3rmNay
8bolFjDy634kjdiGttMilsF7zMpQouWXV4ZLjgEVm7nsMTcDcHNmwraoIEVJMXAyvmOnPBW2dCmI
yYzVqfWctkZ4j1d2YsHKQ30w/M+AWxZsKvmiB3wQlPwXyQiJWv3PzyIgz0svNXCS0avUEuE4r2MM
7xKqEtLZ+VoxQmdYeZvpIoqN/6qDHNdopms5WYUnlhdTb3haqRpe+2VTao33IVZlLPipvySHD9JH
Hf1QnGiT/N/1UM3EPfvtGKHnA7OMo87IJ2RcMWok9ESwqPFtaGgYcXR90OvtMXiTxcK2QxvXvOTU
u5GyDH0wKpA0KGSnpJ5Ll2yTiNIY7W7vQNijmip9M2eqxw7Rl+RcgoQFpEOItbs3yeK2UREgFED4
iq05hNAecPNrQR21/U1sOepz0xDq5MNtjb8YkIGSw4fvsRhsiwJ4nuozDh9KyyKYCBMRc436Jc+u
iZha8HW7GdcNcqxV/scJ04zifCGUs1vj5JUnxRWfjeWfGwYxIyc/Gph+w8Fx/na6Qs8D+oxfADa4
TPlKCY338Vd5Me87ZoysK53iZ1mKuNxtemET1D7cXwLAoaoati6engZE/qHo1oUm8q1eBc2NTEmv
XuL46OG6eSEMZmECPgrmYMP6pZzVbWejUDh95Na7rUhJULVCihwLfIl5EWMMciwYK0XG8VO5zH0/
oRc/UQyDtAyFGT3F3vUXMShT+JgxEfTwrAABjVxrhMmRD4ZqHt3x+d4baNzCABdgUk4ReRGc3t4v
Zn3t1tE5fXTJv3E154Lzg60y/rCo9XokhJ3NxzuadEOCEZXZXetkX0g5SB0ku77DjtwKAWp+oq0c
QrBUCk4gy8qCRqGIpvvxSgmDgGVxA0kiqppoXLJcFT+FHWN2ZtT+1Yf4+g1eh6vQwC0XTkmK6GPi
veFBqgfHvFcIY/znshTzul+bo6k5R+p4pFKHjiFPtLN3k5QoJikC4p6a1MMjxglqNtGf5KyXw9xg
q6No1mKmTCrQo8Eti4hdOgQ/N4I5SMrGxE8JSQjWz2SobFiHJTUQSibL9mV1kEH/fBPXn5aXWhN9
VP8VklsvO10wEuqxSnB4mRJ/0MDlMVosJltkYKN3EmkuTkCcevWgrYE+h8R5vNOIayQX0gINAIpv
JnhCpkUyzcrV2udUjQYVyPDuRdi+qlFSrah4mLkFl9vfNIKIVYrbLi0AM0/Ob5VjBOIcy7hpX1Fg
yrYeL1YWt+Xz4z837N3/jdi7zgQYngSVgQilZVMKvXQe2V3wJ/LERgDTrw2GUPAdRUQW3t9FZBrM
i9rfXqb/1MeT5buF84uhB+9YslD/Tna5g4AxroR7+9qoGd8t85IDMeYyyOQLDkOB76MTt/TC/ml+
etwufrre1zfsj7SI77ZrGreJ6GPUavlkVhjI+qsT5x5Fq+wvdT7Jw3hHgiZd6k6x7CflGDjKTXdf
noM5jOPsEJMVY4o3GXVlXAN6sxlkpaWa6hw3W2iPTPz41QKqiPXfZ3JlS3nQEIpALKJu9UnuC/Hd
pCZTGaMswMYM3NV9EikSzqZcdnZw9emStS5bvhQ/x/pPrEmUDXN4TC5wCN/oTSFHv+RYMXfF+bY1
fUMb4twushqRIL0avw7VozoISJaLBu6XhLWb6LUvCIkdUxKBnRrqMJFckXU5nE66qTsSIdF7uPbB
7RvvmpoKn0q79bk7xa4pWMkKGhDJOejpyS2UOcwotXfaXBUWMWusMdeZ2/R8s8qJbJAkxwFstj5t
qTICgRtBkb9LOSXJFB1f0M/DZyJk7pWVxhIWLyuOiUxHjpt0dLxmGL1zq/hZ/gv4xNnSu+ls8p69
1jS8TdckJDemaA5MpYd1ADM8I/VgPQ2sUby7W3vhGg6QbRYW4euV/owbJrNYoLEL/ZScQZHEiA98
i5s0jWb35UDvvTzo8mvDadakSizJVmvEfR+uN347ogXsdbYlcQHhYwxijz0ul03UIGevyE55SZ7V
Wb7zWKn3fAWQcxncWuZKvENhMZBdJJ2WVW6x9vYZ5/atZV+8XpCsGHZGTLNtNgvmW6a1lvsxMjea
5YqLcBiTcSkJCn7aoKnfw+syfisbHUNZ0sYRYsKrTShrt5BqAHeUV6QRfOvmzdpemI8LUpmY7WaW
fHYz5AEBk2VH4iOD2HEmmcR4IcnrwPYWZbzWB28UegGG5Zi43nFM0Xjgy4lo+B11HSSvqJgsUrtk
96/qhWFvWpml0T2ab1sXhe70BLUwKEjximGn3Kqq9b/mC1hZJJG4P6oQVjSjNb8l3DcI9tsitW2g
9sjq4wWY1TkkajuQ2pge2GnYjy0OBc+X6nxkQpSLyiZTdQxSkcfXgI6tJTKlBNAutJhW5MgaJaWp
uTNXHrwORrGKGe2qDMRR2uo16O2bzcTsx2ZEDbXEMU9QcAK0BSEfGNZZXaFTaLRjSYCeQ541AQTt
t5CV7VaguJ3FyrHxinHEZvHY6UjtVikK8VcUMN6v6CX46mHR8v7MwME81Ij8dyf2AGrKop7hnPxP
NmKqCuMcgk0sQf67KlgU131uu4LOk7FVXnkuJ/+Y7MDl8P3E9Mol6j8etQ9izu0FgQhI37JKyDon
u1NY5zzGybeCLf8mB5y9lyE2vrk4SLer8JUll0UJn1HK5MjINnays7C7t2MLOdb3fhyIENZFBJhq
KdF4yi82Ujwc9u6dRqhmktZmBTykrr+T2EiXK1DA8stB+NLV4Clqa1PcByGikuMaeMLtLUnA1+5/
05sdZ5k9OsbuFhFN6TipkYiMGO3wTqFi/5a4GGHKEoPuF4GRUkOf16xFMT34tFibwra4Pdc/HhI4
x82Q7hLxe8Fjc9ENFrACF3wz4bV8qgFPvb3veUE+fHT4JpdDVm/aoC0w3ltYX9p4QvpkR2A0BMzP
k8stY0q1vK4bNTTxW3uhEe12Fy3sv8Mwg69fynoO0WHmTt/ZxUhmoIRnfYJFdGYaLDf3D8vvfKjx
A7G1LgY4Z2ICbS+wjO4k4RYRtHMucRkOvqbTUw/FU7EB4HkzqGk4liy99QNqhtU+T08EuAvMT9AI
Fv+9xcHTh71jREGDAWOAqoX5Cxk1QUME3JDo0lcvmw543KKxM8nRTU9w/f4CBHbDqr9is5yIb0fx
NBSBI46fqjiepjqSPOwrO2t8QyV3MlMviPwoDVnTcJBG+yERQRHIawRfHh+bjQhFEhDizHDg57g/
kyIB4F8rDvvw2sSMCn1FzTD/JymtOEkBP6+YR9YsgEHHyJVU6XZdUAdmMZ9Du4zJ6Zt1tz0rAR9W
cUMSgLucUOmBt9ldUdUhi9VN0IXZSb0I7uG7kSztxaQ75RGb47KlvzXLCKyR5z3LB+PgUNAVngef
MpwYHnS/AllafJXU0WLjPDiGiWaMT8mj5sijmeBXAsGL6lBuQzk6YNxSr39CzCnBHD132HF+qkt7
Cv0dDhzqpgC4umA+yyZPKR/azpyF6pQtLyVgobo5TGS0nKOt22ATjJ8a6vUt24U2UjiepINS3VSo
Ruh26D2XRPmDGnQq2VX8DRqtfQqaZbjfmQU0hUr8mpt2ZS7B6x0tUT4bUWIJ166XCLZGx/rnYpam
TOFmy9L6XAXAcIJaY9Nn304M823/MudqwmM3Un52Wp7Z60Sbpu8M8EasRZk8FL4JRasxI6izK6ux
wpPjkvStekAOC3vDvfhS5dLm0eRH8FeK3Raf3JQ1jkA5p+SGSv/Rwd4twd6EW+w6Elh00Nm7Y7Dp
CFunxkBLQCkqxshFI9bWY8e1ipaimM+p9tV0JFJGnDGLDLsmV/VaCluPCcWjQ9h50w5qY2mnyX7x
2IvZg6kU3MxzEU1LC7p+lx3ps3hM6gZuZfTz7J82Ym7+pR98CZs0cpn9oaDrK/MbdzDoaLcsVMmu
LWc5LUCgs8d2HotK2cRN26SG9IvGUzJ43kIp4Q5KORYmBoeaQfjMGLpNRE2cysSW2AEMTGhE65uV
s28An8JeUtinjQh6oJyqbYYGXijrBufNTtGbWr8Za5ceh5Us1rvsdgKS81LMmIxw0hpvJAZENDD1
fd/bJILFDM5Kjxdn7qjKTHQRazoKwvDa3+6Ii5ZrbdDjToa5azlTXPSLFq3PGd/KL2QGlIuE5en7
yfT2yoYdd2f1SMS8VkeiZh4c3v0Lcld/Bztwqi8WGvHw2rEzs+KZOVeqc/vNk0VR3Ovs2XX9NCiA
IFgFDoHtIgQ9GScmicWzxq5D+OzZpiV6O0XPi16G9OCsmrlUtXiIcikUN5QnzwM79+V8dlhyT1/M
Ypu+Pf2v/RD9fZepU410k/zOtVG5VYWgTpa5fyukki+JXRBcYVN6YRM+xdd8bD1hhDvVNMlLAyCi
LdNzIhO1oerFLARJ+lw9pKNNZWrnszryLHNammKEqW11Ze1kVgichRO37bp0T6186VtHnU1HyWd9
MhLmcVrRCcEmnz2AyKFgPDR4AZViM/9UU9vpqPRaIG5fwICvFohs9SxxArbJasmYm4LzIJ2x6lF5
wDEfs/fI8EetVxBVK6Hlzff80jztwJjz/Ps3jICaHOk84eeP/JVdAwqq/dufEXQrA9D0bee3t3zh
hSJglnKq2+CddS153zZDmokFuBqpSfMjusdkNPdJtfu3yay+MCUbaqQgvcqgaf6LYC9TuKrtHF3D
vnL/90yowyETGqrWolFQ33ykQL92K1oX8GOGb/sT8ovtWinrB3Sda3SYxqjCg7gjajIViGLgXP3I
D5FaVqcX1q2dav9/gHqD686G7/oIc5ThSE9N68aw4cAeOQXp1rswh3oAu7/Q+p33ixa1zRSpYUx1
1AJcC2X2aiTR77Fm3wfegb2cF37AZLTMVIwJjsm4aWdgePpHBlXiNcODf6t/Dri1blf4/EhtJQA0
WnjXR8nf0XNVnXwsv1L0L6y4AFyw8OCtJ3ZI6H/ULZ02x8KPR2Genu3BTGUcegtrH27/UhTZBVZL
5pRNIaXCQ6Qya0Orb5uBmUH7BZONguO/wUHxbmOSFUETkouCYugGXXDkdUU5vEdgrPipScCYBPgy
FcnzCweY02gmcQD9hyAaElZKYioGPDsVH1xJMEfxMnQtIx0YlScc0WekffY3zoX5MSNk4hnzCfo6
oi2ufCqbtrcTsepq4tx7+/3aU3JGjUbOWUtQobnyeVsKirRQCzUxBfrpeqQMf7hBz3J8DE+vnVRJ
BunehmwR9mMEi5/W/vZCzjUtW6BRBka5EyYBjIqgM3UY3g14qJ1kSkpa9UxTIN6UW4hBZPJRCl6S
R5bHrRjaJAkFfIzqeLW+zlSb0Zma5TYyKbYQ7aEWLJ354JSff7wziJmYt+JsSw9hn4+xsREZR+ib
pRP8dbpQDpAFTTx/p4nhfbas1LH79KL0OKU/a/hjgD76pVHvls0Uo3gaV0JYPPZBmea2mlNxYB3v
aPPgB7EEb2Y8745+kNsjB3Fo0gZ5wKuxa3g8hxWLk8EnPEpymNlvzMRiSDx/UmUhPrUcbz905uNw
s1B9EIygIdpW5ithYNwmm74PNWZ0eOYlMUYu3DkPU/rLMJfWhA75mpV9Zb6m/KZVq3LwtRNRUSJs
2ATyRzxs5fsNLmGWbUY+04jpuexmAI8q98vcr4BDbQkFz8qmuZnZSCBll7Sks93H6CMG0x3ZmuwU
MHMn8100g3j9S6rNOIFLxuYRSy5J13YfqKPmiB4qfQrI91CPTYW7N/nEmv+43gl5ReQVr5GFRUEv
5BVPOC9RG7zs9dm867RjBiAWRAB8cIJ+zjZTea93VD5UkV/YtBKwTQPtRG5VW3gUn5OmhunY7031
nrgqNqAed629AmDt8V68pFUnd5tD6uGJwa2Sd/LVzYYExptSPZRYaiTkn42y59zg6VZxQr8mHhgR
k2Pm+n75n4XbolDLmpy1UoIqRiU0TFbqUqtklgvUm914IP57PFfYc07NWmajSN3IQg+eKmDZ/AGo
qZxMvor8yp8gyGs08KlqQUfJjbSD+S903mKGr01fmlHK4xh2QiR9lq01EhsqRuZznP5F7Gy5XPIc
eDQBfYZOY4kXzYNi3RQQllfMSYc8r6UsIT4NbEKZauz4ouZbUoaw+BACVbjp8RIeno6ay0Zs1c+q
EqpMbxhaAoMRUCWRw0jvXp9IIETvqteogtgquuELWNUF5vQRHriVnZxSWtT5OT+Ec7ZVEzgrjfsD
jU+1x8P8NFhHSvnX46LIIDAPQTt2jEqB24x+KvLspOt4CVMLoVcFZ3NcGfoK+3JekOPM9Ufp33Vc
Tp3j5pn/kJbeaR+YNbCK+YL1ksd+vLOAXZLJffN0clYEDk1nrsbeSh/9TwUifj6FZxDPKc3clWZZ
HYKlDLYCTCgsjOIxjKBAcveKKohg0gnQact6zCRdmXcfV0tcA0E3HP3/RO+PE9andq1MuXfflh54
M3knsxxI2GGCbKg8WQ7C/qEI1BLAF3c/C7/4+LZQXZBXMsgfOIqnVPsTSpQinKyZ9S7p2P8TajH5
cjOneiqLeX3aG2IYmQyQ0GsSEwYXXL+68CV12HHPz0LB6dgvaDGsEf7my6raRSsNnF7fg63N1ctJ
WyAurl3l1jHfauFR2EFQnpcagvj1gW9liZBD7EzR48Fj0+GJ+9loNPspET7U2ZxxvAQU6c6NGoto
8cEx3kAWwMlhKYBXj3nEm4ZX8w9/YDN7f/w+k7Kzp/l9oSPV0W8GEf63pYvY0YxxcRKfTiKn0JQn
US3Kq4Nmec/WaCgf7f1NF1RqElr99CTTI+TLdf8dPXL0bZIRU1mFXMMbmVlI9+fmlV9X8CRqLON2
gkwFRXgL7Os1yKAajiN9q3mn2Xm3IMZjIs0bD3ZG2Ol/2f6bTsc+eMXEjAC35tmIiH/+WscmvsVS
N5XfsVdTtubOLK9h9cI62PzmSWj1qzhv95MQ6ElXvJsP0EyKWUHMD0UQBCss/eIvfRpMGj2sMYJf
5DCtGTjTQkwYbd1jFgiJYP5SnTCE041w90lpTG2DysMMSq98evkpHx8GS+JgmxRO0daN3kffHMu0
BbWww73ttlqxnbv8GDJuQAgpxS9GC0+f65yT+FwIuBqxgmNOeb0Ikemyrj0K4NIoSuo4hFUoOWSl
Y3rCdn8VMlfHd95nS5rShz6IHnYGotwcupTF6TUmit/hpISaLfx+LYTfBMH4dMh4aEZz0XF3fEzV
E1SQRkftx7KNTsQGApyKuYUlZoO95EXF4kbycx93AAh+guTMFjIpZvMZHA7YGHLJEveB9ze2T6NA
nvk3VcfDcFtCVy1NL6Yt+SFhMUimCYCLa5ihOqYNCNcH3Wl6AWPj8TIbXPL4JDORESVqgw+8VayU
pmNoqsSPJYAKWOQhs1LrMsRe6pHbNVkSxPbOfZY5QuQh34gZUwMMWQei9zuTMtyy5Q9MrzjdXCql
oRcwmuwfyIhtW5Ngzm3/G6h2o/pjI4/Ovk/Ew00GXb95pg5nMb3831pgwrAK4AP7BgxlkjwO2U7+
dasXWxmszoSZQYqn2UzSX803yvynXdDT5mG0xo2hwnB2YFPB4Pc0RerLGgdYO89Br+VSdxLdLUIQ
Zkp31IStLLhhRjX1oomtDi/8CFq+pody+Tvg1nSlCqXJDudIp+3Ba4cDEWdoX2uEtzHcPixxqQ9E
V2qYUPI4i3n+IT6gaSMMwepxkdUTwW7XG23Dc0az6BdT6ubkqZ6C9xKWb6FEuMnGeRtN1opgWTtB
HoSCbAtsB1W3kYbNKtA7aUPcGwonbIz/7em2FurAx/KqVwyovGGUVKDZHyJP+Jn6he+s+lHFF3XS
38pZ2x2limyL05cEwOsswv0VH11bM5XSIQbcZ1zoKatx1NdhmSvDP9gML2TIGvW7vw3sK+TvsSd9
zOI1OiMHAQQ9TRxgRx1+5xZ20A/18RkGPLUdlrGtn2F2hDGCqTPTSsknShK9oPgHZRfxs9802Zjs
zDN3vEdXpMmisRci+3JC1fvzF+TIro1f5OmgC9+dyqsiCnN/DXFqGWSs6U1P0B0By8DYjuwFyqw6
wKNIE2Gb/4qXnurbtp6iK3BxPEALrAvj9nC85L3OanEWAyYUJPZ2mdaa06kWIJAvZH0v7PDTw38t
OdAzhfRguRa4jENcUpJ06qYsG1aFzQyoo5NBN62uGiZI54eLLP3i4RbL949t6/LQ0u69dbc+WKpq
V/X0+QNQgOMh8wR8lqqH+lsuTg2AWNNEDUAR1TVRcyRMuQuXEkMScyM2PFauscHVB2kKZZ5O8DSP
QgvR64QUWhtYS/F94XbOvtxXXv2WOACtidBn5aunBFlY7gh9d4XYhOF+jL5vN3u/WaQhiFp2bjQ6
34ve8Mo+G9S6k1u9y7s/wGy/MDzRmIU/qXeJrPfQZN7M/+2bRbLwkTyLy5wP9Ey9TogyiUodCrdT
inkS8vns4Cc6DjMxh7EGG+WHtL9dbiaLC5B9Imx0vFR/7CaJilbvnyHTqcQR+UTncYPigD6loGTh
CwtE5ycycZpPVxrtkwUjM2k1lJe9EivU3KJqauPmwWz26CLGf/6xku2TaCbLBX2tBTvNMbEUjj5X
vI/KuP5ERzv/XrIo6leRLY9KNXJfStmcn2eY5omPJzz0FUkcPguIQvmOCTU/kuEvRPjKzNR6k+gi
WnXSTTeD2nxd/Fm6YReZwlJiNAiEITBqH+9WG1Bgl0JhvYdo1ayVKbRaMYVcwbm+E2B7+/pJbrk+
I99axrzs1ZOvlOWpfHXdz7PoROSd9b1Hj9Rm/TB+GBuSOmFwSh8pKjrsPNJix7yXkDyN3D9aP/Tp
i6OuC3o6ReoosD5OQuAEB0hoYYVEm1a4czDXkm4YBud2hDy3cJXo6Z7fwrWsYQgaI8/V4T0ZzNUZ
y0Xq1bJoniS9MmtmA13ejdV5fgEM4BCWGyVwE6Hc5HD7VQm5sPGTbKg+PBgVTPzSW+NUT5nmbcMd
9vX7Qd8sBxIANNIk0gt7tQjit8JOYz8i9XL31YWndMyLRGYQIP3G/EMH1PGgjF1bqy9jceypL9WU
3lUQ3tbEHsUbEqCXUgPr6mYLysXrSzcvTvLgGvqcEFSOLV9J3VIbu+nydfR4s0RZFAb5yrGhB0C6
C7nyMGX49bRm95WFdpMdH7A5lVZiL6yvLx3gqTXAVdbO4sp3FL1wpwXXDfUXuWMauryGYw4o00W0
jd+hcUxneav98+xuFBYAFw6V0liaYSrAinTRB1ISwN4To5tyldFWPzjYuvyHie/YDRMbiveTwncD
wcKnXva4uqAqVCBfCRS4h3CgzrBe6nuIXZraDtVyIEOvlkR5XrqbZpgU0lwpFU0ySEV6BH5a+XXm
nmz5g1JXLJbxWt866Mjv5AXvrl8oqWLCScV3+ennJm1hRnfvY1hAsq5CbjKBJ83UEhPzl6pOehKM
cl5mWXVB86NiU6un/A1r3dwxz3RuztGJzgQNSxMgei+v5ryTxr0Jqz56wXYqGj+jz4aJspf0rcHF
BoijgStrqhkimTW1Aa+8oqMLRXfQ2kkSrON/tH96r13pakhALe+Hv/kkWdejXPabohdPNWxJJbi8
OT47Ww813K7fNY+opvbYSE+LVW8YEof+09NMpAWhqU8FU90xN3OqulqJzWWYYaI25VwduXKvB6nW
GXoEs1+ADVZE6dFUxWZr8I9YfbmKdNf7hKlCtKsA7FlqGyPJ3+zYrng3EBHidK1xMSawq1yltTqo
nR+BXPQuAjQZ5S3xr/ySXiI86xjbD81vlb5DAszS51mMNzvdht0X7lLdohAhn4QrQfuvgovHZvg6
cqNkAFlGvxsd4oYHtvNDYScM7TxFDUAkriOvetmoaw1awkrOCr559MWhoimJ+2CjkT6gMNXtZ7kO
l+ytoLzUbbIQtZxJQFFJ1mhZJg4yi8pCw536Ag5yiFcV+dJiv9sNzMs5x5jK4kB7d/+WZ8dN0/Gs
+QtC+uy3qtMesFYj63G62T+vXmPfDW1RlX9EDZpkyPbluqG4FA6QCx3MHRy8q4aDVm0XNSnqbFhD
xHupKq5QfF5dHdg2vacwBCgZ20YzOTSKdXVwuHGsMEu8Jao/EAgYwVNeNBwcSFn2ggYI/QWLCDEF
obrBjXpPdLd+5H98SU04kUoFp6VloNfLVFicOa7b/ldgX/tSDEBRXSei9UVdOv7GYFN+rna28UT1
iXK7pjvw3+3DC/RC2trss+jhnKji0a7aBjRSUfL+gi0M70OREMj6SPuMXYo9GnR1aDx+m2J6Q/ze
PO40LUTBuMXeZg1CYqeiEscSn0DNCThrRhbjSqFx72cn3ETH1bEI0pcBQMYYjkwEyRMAaJiRyE/i
mf7fD0FgIpeKaHIM2noDbywwocctL8kKYb//DMqKlCPSVw+nsm7LsQ2iiFmAO5N2fxypzPXY/kmc
ODjk7lzxiD124Nn7+JZ/VVc6VDovmRNdTT7Le+gEqGSf7FZEh9hNLzA4rwu08658aoiNrh/VjMxj
NhhwAPl5+Mj0f7R//9y38vfwFcuSICwx+zeCUWfDU/o4SevfIwGyyFKXFV7PXyYKVHe5Zy9m3LLj
YRAb7L5SUsURtOSRbcvakMgFJhr+6vtsLXSN7RKfAAb7qx0BCoWzBlN/uNjTUcwbqYu4u9eAWgS/
9uT1iBXb4v7efsAXAmrggazWhkdFkEx7EjvkqiVT3VUZuqitRZTW1CZXzkJ1n7WoPf1TzpOpk/CA
IYrE2MLqWBR0DDyi/D9iXnnrYMYuye3njQx11NhmtqjFR0DROsVoQT7DR/OUoLQnAuhJgR8l71aL
8DvOSWliu7b+ZIQGk3vEC9B6mz7CU0N9b0m4sNtu5GV5dHSG+cu5fOgsAh1WzUvuNBnTg3fOjgei
LSfXxcXqZyupuW3yE/D4zH1loHLlQCcstMwspNQiE82IecKq9yZgtEl4Jzqi0bDuNLONH4dGlsWI
xrpNDAZdkb0YNJesYzhOu4tF7zeCY9g21+KkMLlVjYPaFOHxCSbNKT/0MwfYRNsRwGQCZDU2WcDF
zY1c0ZCE/O+CvLuhYcmWnXJ31DPpWFCoREMLMF/eGGyMJYtKgj9Fz5r5tBA9e+kINyURKXNfUwJT
6htvUwLE7cKJR08cfYJ0YCEMYLeCCE9FO9PyLu3uoYRcwRY4j/Mmue5WqcH57sJQ9EXAdtB4Jbtz
cHZnSijYp4KinzE8HMt87QgyTduGOwjCWOFYuEvXZVWr5OQhx8rfqSHfvoBK6idmAtHrMdguDUjU
arBtIZcS6yb/mepEvoaufu1019yMIa787FLKgqSCJ14ajkp5mDkCrqEWaVdBWz10nHm2J9KziQtB
yFnH7EHo95QJv3FaDrJC4xGxiwGJSERZgAI2x71mWx60NKQlYran/A69/zGXqTAohEZYEkHloEJ8
CSteS1IMSzRjW5lA9Utr43ELUWWJQ9Gby9yzVDHOqW1VXms0AgjiM/84Nd5z/mfrolDCTlV8Ke1f
IkhxypiIPeqLspAaGwQoJkMlQHimhHaMNhB8ndwYYbKdwPqDtNo0poAa8q3Y93a4nLdTUwUX6Ail
wGcnj1wI36zSg/9jtbyfgcCq2HHgeg5LgZW7AMj+jH//IMyg2Ebae+a6Dgx8uufu0I5Ctkb9e1CK
D/lH9xyy7Y6wFUEvfIeiyzl6dyJEarKt/7/Hy3roM1jGjTWrcMKqZ9C4NyTdJKAGWDW2cSIV3B7r
+b5NLqt91A81MAzPgdoBFzYdz6m6T0kvZRaBL+VIVp7NaKZy4Yiz7uPpAHhiOZ+/5YtOGcWiVNw8
W74kQHfzqocn9KkJq2v6kDWDBI/9LQbsD51X6fsOv9L64S5Vng61GPJmtmbg5E9WAASgiVdBNG27
4s6XDB8jgSFbETuOMpSuLb3JM4iTM2eaDskGz22IiXNJZIY6dmQRCwMP3sJm1pgulaPQCOt16loH
hUyrlfKl2RSS6Vxmfei3to26xnSfXHzv+AD3H6iDIJciv/9jmFW99vSogySlsExZIPnuxn9GVDXI
1PPvwCRgo2rkQqKhI5uU2aSpP8dgNDpHBixG55MbKuICRQgd66k9Y5KYX7WrTe8d3wqdy6zkcQaK
7tW9DVWQOMMmmdUWcHALaVlOwTXsHJAZxNUcOifwF0oONBns1DoRgFL6/HtvefbgBhyaKC3pPl9M
huRqX5yL1rdvJH6NFQrypIHSUM2/ZphdzgLZY2yPmv/7M0xmnMhJ01RkWSU/tP3iDVBhA4tY9PpH
24BFyGtabFrSqqnlpB9sfjny2K3h3UDib14H4AmZehuOZxJiv5JXYuWrO7aFbttoeBKtW2By1EYp
CO6YUOhEABfIdT88NpXNcU8tn5EdCAKaQc0mBn7bGnZTtzJe5fEoLyrDpnuAA66orm6NvNoWt43w
rutcPovzQmtq4x1xH6yIjv/t3XtHGMfMs46G4F8Dk3etBocfQe787ZHjdh6KQCVFH/LEjCn4VzCV
5cpeVyEtkPVaOqKyfjYjQr1PtkzeqTNJkzMXUBkSxJy+PfF3BYASm8norfuFJlzHhiAxFtmjFfHX
2ot7oHf1eVF8ekQ3eMyPfKVlcAXan3u23akGHu7XXDlzrcItpyXNSMt7+IndjIpM0zzyv0FKA3kn
2T2Yhj0H8lzkJdBoTv6FbdT4P7Q3ezMG6vyFElPofDb3RwjQjv4izkGITck8Xeq0rxaTBDYaEIjV
wz2SwQYhcsuptOnA762aJlScXb/G1p7jgOy9m5B4kjfE7kffY3Q6vA26pUx5CeikbNlyqcfs0vdN
9X15FH6Tg0PqXoZVrdVb9N+iY3stDzYg557nrINLARogI1A8xKJlt7lNANwpBzUG5JIMzpLAo65D
fjdk1nc5C1bND4+744pJV/0jvgFciWvLyeqTLoT1XSSaqvyERTVZ8twxyFwgr89AVuclkBv0joYY
knXUHjZR3aITHOZcD/PY4saBhMcEm+eC8IBHgm/9PpcNBFyqjuRAxqWn6b+qNW1HDZpml9A+OMlr
OQqweO9O9cbZRu2AmDN9aSzV3flFL5ERVyiry8ocBJPgKD8HiwC/7sVLMf8TIZfvoyusri6sPLpM
3ZD05KM3vqmQJQF6MVFyKc1FNm4r61CNr4VEUmnq1eb0dk3NqAeHXRRBv/UzbbQxEZGsg3MBtw9d
AUGeb/aQYHt+xi+sRK04zLkg7rS5YLeDr5Fb6+wtXZ9C37LIEkTijmar+QJ06WI1q7NHX0JOfuVh
oZpJvTTRnTvzToInGvE2p38uGhYGjqirr1jij/q0V30poA35+pZtjkyBJddzK2mA8N6NwPKnUGHa
juDg0asu3GX4XIHM/jqCmKYh2Abpdgveqq95F+2VMpwNspgc5YEFVzNo/yaO9+kWMNHwyx5+kiUO
5597I4mo2oE8Vq59Ekv4CGOTn65PKKgAVVEvx6BAZQmfJDT9tMN3uPiSafHbqvqykNfCW5N1qTyC
o3GVi1OnRXpaoszt7x2R4ZQCkfekwp3z74vyYYhgJNKbJf35X2QUM1eSRUQHxY696zgnSb/O79Af
kWeOGkaNL2mnoqQozWUGW7FC37y7uEfBIPh2NsISMOPrWkEi7YDF/i9fH6sDOfbOXFWnSUK6A1g9
0/oFxr9LqceF1QGq6GVKjbl7woAhGtUuxR9fAQvZwJpfGuuWDXREGwIhs7hDHjZm6FykiFtvYGMw
Atb7IjnlKNQ0fcU304WisT2MQ2HFLCiXqTgkgTKjmKx40QpL8XAFub4nBy84Q1NstkBEFQ003gQF
RGJCWllPeGTr5JwGA8MiujlxcVeoL6J9APsRpd9mxHaNNvlK9H/4X+qkcvcYXVrWPXcJSdJNRFya
uTeTYRfGr/2cCaqESDcZMhbiavKlhN+JVWclsUZy/db/zVvUhB2ETdPPLrMn6ODITqm1XMbP92bG
tSKFhB1g+p+ghfH03rUXGS689qz3SvQB/zKX30mKk32AsvCiie2+Ez4e7PTnpXRV3HJc8rpPj8GG
UbRuEwG0QEg5uaXiU0Dhe7jHf7w2lLaQl+bYFos9Ftat2gKAyPrWepbRlafodeiA1VufHf7A/WYu
Xz5Vcbslo1h0A40t5bi1yAIAXD5guuixzSdS2MWzto37Pw97MEIGjctEneau1/VXSGsGw7oETuIy
Hjs6V/tKTI5Ja1SQxS4sAJNz7Uxj8j2IkehWs7eQgzrk/xCS+gDylZ6omCvYmauWiTTrkUhRvi7Y
dDOVNKjbKByvOqYW7i9b3keh43c5HwRf0lSRiTYP+6QCQGhfpp6we9wk/iwBTIX4iLm7MBJUmW2e
Qo8+hzMOaYAbGXFqLy7WbMb57vSUfvWDxM+t0gXe6p+gUHzSHRj3ekGtyHlbcMQKmoUCjk2dlCPl
9b0aDmxR5SWwRy0oVAWM6F4Wb9iqu+gTgjfYqSfgARVXhiJdVqzG/RepcP3Pss+RPYYyYLHqZvPi
G93+YIvjTM1uB58BiA6G4HYqrC3u8KAZ6PtwCeYRLPdv3t0ZXR5LwtBKw5aJ/yM7CUbkPWRp6xCX
wPAX5YnzSK9qJ9AgS2VEZQHeGQd0Nw3k5lEuyRIoL8yUkFGG5OZlsSAOcBdcv0ZCtVDBEWUPJvj+
MXJpc3JSObKIgBi2cLrmRktlc2kX+fT6hPm21hyOf4BioQaV1ChKiBdJmxZD6qqcwh9XEaZ3dByH
dljtmspdujd4EXJwr5s+tR5oiiiG7mMDIbn72Aau4o9cRh0jaNrkHVW0Zf18HJIK6qGQsPzpWpVh
EYJGzzOp1B4dsfKy7SI9vZ+QUTkIdgUz+gMH8J6kiG+MZodkZk+WRc8JJDj5qU/tAa6yx1VbIK+n
QksKyJak0+AZHQ4qYMCJBkXdeOio0Hvb8kuPTkX9f9Y1zbz8Fe/9BCJWwmdowLUsK24dq9sZYJx9
YPvssh0nHK+y+0Fb1B2Ft0oVe3LZCQLr0gxdoLksslCqAfsFTTqGIEVes60kHFMxruRr32ccYfQa
akQex2PpxTbR+jWV2JNhBmna2owLenpJn2P6mEem332zus1Pv+n/FAqC6D1omepZQXS4c/7ny+2i
x/O5QbnqGpr5oi3d/Q9+vZjY/DFBhsX/G+5QwvSjVgTmDetGSPN89uXj8KB31DT92Yb1qqEZpm2w
Pf+nuNS1HRIMIkcOpv86IXOdOJcicBcgUk1SefwURancIbD2rQvYGAUHS90jpj6fESIrPK+iW/Sj
xxr0KHUm6IFKZidS9drwKGUaR7QviymtQjfD24kmpLHVheS4bsOx341/xzktLrE6GFr6Yb2AcTTM
Alcta6sqaYLxPckrR/zOIpD8pzQAgoLjv5WezWgVNJWJZoZozJoPRaUaWlXPsbeNbe/Rfq/Rt7qi
+8dMFi9p7FkCrb6Osg80fs+0CzH3eSIcPFrnHQBQ3jMnubOKT49IR1hiX50w1Rh0ht1emF33H0T3
fEQAjbIXulZA1K91ztnd6byU6pY/JPNzCGssCfbnugCmX/IGaQmlr9BXfLa1Jq3dRc8aKbSfxzNO
02HX3glo0zfFn+Ft3DVOdHNvIXKuu/06G0o6SyFPxpyYHCdX0a/v02bUHSyl8yvLHGt+CEWef6CQ
csGJuYCHiVtSSTSlRE2qBnLFOECtCKS8sKr1weZ5f3KsP3Vk/zbwuocwudp85QZgf/DDOObkKcqg
tCrOWSBzness9MWk4Xe/Bgr9SH/PJ3jKq31Pka0f/JQoPHJtCSns7mfYaEjAHCwwocWMEz0iQDHQ
cN94PJ9AU5u4Uxa1XGrOQrFgkE1ginsH+kCA2BehjuJqb0roa+pKoSbDASY7aZlQYOiMdiUEhwz7
a4mRb929NmAz509FqIPF3rK7iMCjqHDhli+ir5a54jnS9T/4KD7QJufmyaidOwLb8Mv1eyzmrI/i
nEXYrO/Lupk0D0JrFKVKxLxY8TXyK+P+YkGZVxRYIWxaHxmf1kYap5SsHKMNq3BlTGdspdACZiqv
xzLq4fMPXsUq0cDgutQ9DxRGLy0qE1xIyNmcgXVJyn1MgKI0bTG6Q9G+fAD55RRIdsZAddmhZscb
5yx5wXaMzp3whyUtNJAFfYIiyyjga+sDLtw9uFdvjkoewsMMijosF+W9wHfAog365B1H5uYme6f2
UXc7dXdDGl/1K4H0sT07OXwCNPnGeAqb89HGrd0k2JXroeeZiBRh5UCdEh0wv766YE5s3WRuLrG1
dFzKIisEvtQB0OCfzHhgzwgVgVyL4TUyBRt1lN0QTU+0eiH3OcyL01KER+JCeJXH2nQe86BKgRm/
RizUzmZwqmCF59UoidO/h05iTy6lHqhZEnuG9pDE9ruWVdZnjY8kVDwtJQRVbUtR8eNNTxWeDkOB
5DJLaue5SefjLwc0KYuHXUOQQWNFgJW3+UiIA5i7HLP5qWjvzb+BdFQ9FfrItbZXRQnqjJyb1U7s
VaOuuR+bf5wu4OQ9srIG4pGL/F9g8sibc1l5wG/2rfw36LMW+gOj1W9neIkZsC9bZg63cpyP7cdY
RJZYtSMNczv+Kmv2x4DQgYmwInvhH12H9CqNR2FGijb8qcSN3ywBGdKPND/yymaXGQbifmTeCpzf
PE5vcFWV1KGyqXhYhTF9hJtHqkr/zXBkQSPQ/PvTXHAFus5sJLUY0rQfQbyGs7fJ2HF9v33imcvT
jeQs2hHq0lVIP2x4ZeKNlDO226F86ykMUCOBx0EPzevBHc9UoZGfpLmySAB29buSxiN7kbaFJnit
nu5DndcDYxuQS960DUT3ao+DF01XqgSYBXxf0RlHScK3qSIs30lBdUNTqJ0cOc92rBhdb3Fgol4H
FOQnFkWvuugGX5bF/C3eCO4q08ajcV97abi50x+IS3j+TqJeLmZltqfwz3mC3Trd6N1Uvdl75tTR
+neOYnwfyCwSjdxgVRfLXOLPgYssuZNl3Xpoqhjmpqg0vFoXk1E7HipjLpt+gl1G8UhVSVVtQ117
97uJ0s2kO3CiNPHSowWY2Au7X+nsC+FShW4SPFjj14UUEjxrhR72oNi5lf0mqlB8nh/GiidRQ2Xs
ZBkUKDj1+7of2NUtMFsNw8c56xTFA0sykYdhixALDvpccIEsotARiqpq3T7yAwXq/5CIs339yBDH
L+82kTmIlriFyWHJ/hdiO0TiYP5msFPwXUaNfT6sIVRjdLDoVA+6xQBcie72joewfLq+IMsddmMA
DSCU528qTuawVtiAorLGVkrGH2cYVwMNTTby6/nbom+mMlR1wjTqIJtHWlLAUff8Cvp6WZubMLKL
2SLeywur52jyFREtg4oFjhzLKrrHEMfgb7J+1tUyJ4ZgJ/3jShAopwT7Lgj9w26fXrIOKQaur4Dn
GvzTXMC+wM9rYPe3eDYEcYVDDoiFa/kNHB/XjqoAwjWv8AfvS4BxLAznbGtefHHHWrv9DXfwr36f
487djqiK59G2dC1Vs/Mrwecq2JOCWXB6xc0+1fdN0/T30oGz3FQdNMn4g8VZd6nJByXU1sBmFL0b
47TPHTf9wY+VuTH24PuKAzB1DUTkZbwAJ3el5riuiFzyhghgjalWkGdEFSNRvgXhPqza0oSn3QHq
VhJhMvs9sXQ/bev1EHqxO+nWU6f2e+6dH8j0aNCxI/3ztgdJNzlzKQZHswuKf3LfLF2MajAVA6wq
0smLd65eY7Nuea16lmo+XZ3Go5q29XCBniQTj61cgzDQ2li3xKEFAxY9F+LlnOgwim1CtitRbpij
BEjfipG1NC8Kwle20mSm7QztollpNYTi3F+9RhJH+rOzB2RTR2LZXr9m1gK3w5kymy0Z9lhwyCV+
n8F7/qoksqM+Dhu3oK1O1TzoZduuVvFbTmaEDPfDinkVilwfzKadEoz6PvnAKwpzu5OlgvB672sM
8Xox/M/hBkJ08FGBsoZCHDcuUgD7Zy+YsIUIvoSnxAzjCvbC5AhhVt7Ly/yDiQJycSDvkPIQVXsa
tQJJMPOfau8K2YeQ/PBlLxBA2g5mXrMUVKrq+wYKL0zh28Da7HXm3xpip13g2wEY9fzDjUsRnVB3
QEvOyCarCUUxmIeXY9nYpusZ/9pTyMcCrxnWOaQRhFc4Kkl6M71IACPYV0988qMrypCOpXzfpAER
xYQ2LFOplHkPgxm7QC5dqeMQIhuztBSg9Mrv4plWzoowFGVBuRqdmrTakZ4kdRy9PnMcF4yvT9Fu
OC5qJQP0nPONByMbLZRAHVqH6lEJbfcmK8nXxlJBS51k9EcxsLbgH7hytq+8boL6CnKw9/CYZGw6
GsigpSdeedEO077korTAq7mpSUP3Sk4XvemNSIimHFGdgS/G7WLDo1vubqU/Q2cfHxYk/pcVPJBG
F7EnQA6/3SCFO/WRGivCT9TwcOjl2aKSYRvPgCrLrE1V+IzLW+E3JC6v3QbonILWuxNzbsdTJWBH
ZHWI97qHbljBKnhrxQBLPt9rG25xGkI1WmnLIIQd67blqqCYL8FMPZhUfTPUhQs6ouBk6Fg4pcxm
qw6kX/IIQaGy1vsjQUQZzTTzjHGrNdnydEc2qhGGGsV68Y5qGN7Es+3DTzmPXHyHdlpsGIXylx12
rMsWhyyrH18TNL9ZNXsK1i7NW8/HbdYwoEQre/RAoyuC85z/Q3NXYKgldfmvleTogzji1aaUovlP
H0MEOtpCQ0zx2BEvg7GfXoY0Mj5bP2LnCuFUhrRKuIDmoRoIBu3TC4Ck6kfMpynxq+jGLzrgZzXh
mBlyJNwW7wMLDtMYyNnnsi3o3npre++rSshxEUxo/M5Mdbyrd7v/4J2JmPuYVu3G5Jfw+GvBcqrP
BNZN9RrB5jLEBWUQVhxlaCRlVEtBX9xhqag/G+o1J3qVToVcZiOU0mAmw70MPcCJKttfKpURVZnx
b/8U7e5m3I+QZmtv5DWl4iIg8CfoAnnh/QargAI4ftbtr0Wmytg96dAjtN7QECH3QeP8ofN2dBmf
Q4/3MyblXZsx78Sd5eqYR3SDcx3KkqMjhn40lCHcyTC+mkea8HURQKEzwY1BkV1vcYG30uZFpgUx
SZ6bopFz1wZ/jo6X7nHGVpV9pzaYz2vI6/5krxK29qaptHdObGcRn4wGWI8/5+j17M/qhTulk2Ot
PdhCxBWX4B3IRwbNCAL82rh0yGjYV4vfE4yd2TMQVp/w47OljQcZE5r9E40RA19AkEe3HJl1JU/L
G8IkKTiVhg3cEH45mG/DTHtw1HonhM4WM0GWEMKbmlVMFP3fQK5gFQfb/6RMpuCIG29dDfkqx8Yc
+jCW70h3ewQLJn2po2BzZITCDhM5VSTCRV9MWDKO9sa6o4ZSpKf9uptLSakR03Of5eCnbmhv1lw0
SS1LWZ7Si06kHfutf/5yLyWKiqFuqTnUEuNlyhjw3nbTAsUK6VBlkigNk+95SarIWerUB6m5X5/G
C4dg+pOu7NGShXKnV8oJnPNPS3Un30IpQiDBr4XmCkzPAh/gSwTFa5BkKeRDrLyARdKFUEgcFkEV
u4yERs6hpiFcwQwPKwNepvYS2u278qqKhK7DStaeEgyD9Jg6ek/upUqj3a+7CaP/wXevmsRRQk2K
Lmi/eDIBAdu7K7J4sPeD6Z75Xh7L8ZP9PubrSSo85RbBOJPstBX59Si8wOBCvxTOmql8JWU1E2CC
CeZSjze/0wvnhZT1Zs61bYBbEnAdamZ2DdWfc75uOz0VsvK8q6eUIJsqeSSflUOPUMaXsvV6nGTV
jH0s5qjWiAZ5EIogEHKmWVbh0VEmcS0jHfMB8/FifTsB44rG1zAaVmtR3d1jn8UVAP3P7ncsmX7p
uA0GAr4ZlrewrmB5XRurDgVgLvV3gfg9EEr69FEvu3HaQTTrzafBKvBfJu1xl2B4dxkGOj0hUjbq
aw9GAYAzh0qT39aZ5u885KGHGYOkiA5FZpIZJnt8Mpb98CkUBLp7PAgD0aWxL4DcB+hoGZ5vHgBI
b7HaWYEUnUoaoMIAUkIY1duYIGwHkKF+YEeqU/4DuY6SUnqWS5vSSeVXm5MjbDmZ43ZC+qwCd3jq
SdS6PVGCPi5jgnSnuZDDO9QA4c8dnZdxiexoiRKLyh2D0q+ckqW+wS0wYZ5CobnOi1GEgtXcsB4T
BUjDd2NDhvqskN6nu5zY8bkYDDNWE8z8YKXsDhIiSwh+5gC9Hs7ntuRim0nwiNqey0tJoERt94QJ
ohFGUasvPYH2aBzW/oebhM3ffx8lgUUFGS5P8GdvjyQQtRpG0K/uxCwbb0aThHT6ypysRIZ62Bzp
30uNIH7GDjMydRpldCzlkzmZkyokvlzRAHDI4BeJZicRA/thLsMURZYr4GpsNAxmX6ty3AI6HNkO
0SdwHh4JY4ItorZ3r1gNP0YkXAbidJoCsY5Yd8++BqKi/jQgqlOsehzPFvSygC4Qq02Ccm1KVINy
WFmIpa0IeeLkzeLuYcxAVxp3YWQ6B4Qywp3RYc7Y7PnuteubWtpgyEhR7vWc5aM07dpR5zBY3dYm
6wPm1tdCE6gzrl1gu+NSkxE6dYnimCkY2aTlNHx/+K3DB2InzoCBoWJYSDuyuULAi13nDAWOl8SZ
g1+7tSgQabOJDyq1nnGkSiJZRf+JMdHGbd5EdPWVcM1h+4h3JCHEy17EqRnIpvCfxdj9af4PD6Eb
vpxQSeHu+NRrpKfhBOaBOL3TSfx8yYcTaUey3mO8KiYB5HdVfFUvcYWcKdOsf72qKLvuLbthbIeV
8yvokGGNVhzZRhBZfprOEWkjY5vB9Yn+HCmvQI/Tb0WdNNHAm/2xI+re1DrgR6rlIQsy+/4o1Ibm
mpBWWUx8WBXSyYbAm7moT8CwgfGOFLZQAqWxgUXmkR2ovXeWbF+oFv6zPaZwyIVpJP8S98LArXqz
p30Y0gPwEfWovE3hTjATckkvJUjiiElrxv0ZIu4SXl/Ezak0nCwIhbN3V/MsKsKmmTWxgMGjVyzw
anpy0O0CqqiNJGRFFOH1TXLtUK+2ogXbIPayFvY43jqHbEoQ0GUNIqh0ULJe5CkQI2qQCpOtxpJN
KO+VZCN9pvSwZRPEbzee5Fqj1UUo2UGFkxFFZSBUESDlHZadIzSgI/WBG2amkh8Fo5ODu4WYSoHx
E8bwM7urVo9kVW5ODJc8ProniWk3LXOAjQENmeAmmTXnegemfplIDbJFMV/nmcm46bgGNTf8e720
brBdACJ/88KeqdKu0cdRHlpZYqHLS+fjYurRoWRJ5zBWBsJlyMf421ElCluUvKDc3/17W8kpGBKV
WQ9BUv/zncDNO6nyzVPCGn7t/tz4X4fY/xkNVXki9JpkO9yO9mJcDd0fQvGDBVtON70AEgT6oPpM
b66mDAZPCAS+YzpC6t3Ii17WEst1zgd15CSazLkwzUTJxKaMuNtiMLNeS1QhKZF+1kyC2KtDJFig
27oUbL6NSvrWyCGY76HEbM51zmT0IbJypcyOr/UDsw/YCmLO6rIUFZEdqlz1UJjgBaiJBgBXd0fe
H7q4ahJcSUgek5ebLZvVZb9Ucq85tvtNFcwZcjzfuLGTKeQignVoejRGxALRqqhAfXF+QlTjTX1O
X+kvsZGM4OeM3wTE73rMNigE8/80yqfiDb3RSXfogjZnnDyoMTQgjRA0YXBGWwZORRxuUy9aQVkN
WcuSp9aVXoW9avXEqEznIk8R3fqD+7EN+XBoRcl3C22oVKZeDu4VCHJQHh98lVilUJ3Wv0cuKAuM
PgPFGBQzlnTCbD/GQxEJwG6zoOoU27dx1yV6wCIOJ/l2rue2V8a50ys2nKxhlmAyOodjsZ0bzYz7
zT/Vd+hnBDTPGMQfKaK5SgjiKgQDZwkYU7ejhbpwo7CCG8RMhfRGvcwL1GtpMnMxTj9eAAnmH5Hn
HSIFBFBB7BhAY4PhBQxhzhqrv7/Hkr3EJMfiBr4m9Ty1hMZ4kHZu2LCb+YKbju7H3PJmaC94J3zm
/3Gw94VdRT+pLbMjyNvdHjTwoe1CgRd5Ry5Yo0edhckxFE/mivDhzWvxe+JXK/8QLyKcac/kuqd4
nUHZjGxS2Vqi7zs7IGM0Zch+pYwktlGaRh3vleSSteebWYZobW+26hxJjOeP7BxsIcuipr4UZ6bT
dyiuv5TKEKAKU91hW1cWEivecak82BfbhgWXFbZ016RNb+2s/Mp6zirYsiuC9raCGRKBEVVCBdTa
1ErfnwRkaRcJChZ6cSIuF2+ynurYq4ngFQIM1cQ9SeQ4TNkCVxAL4CF/7wB8g0Ar+RNrQ/+Frc2C
Mg0eHY9c102ilZSvlUbF6+c/Rz9SpBRlQN/dzgEwfeaMVPYDQxFD5hTiNRYFrHXnbuB6o8bFmGnz
YdnWUKYfSx7BeMykhaDvcwoL2I5Dw0ZWy4BuNF3Z9YveVvF1cjh4yBiHDUut0gMc25qOsQLZZDUh
SWIyNjhdxfC+sS2XQg6GbfBE27dinFgMUE2eGzFjM7HAoHo6SVV9/5gJgr4jWBv0iyN4yKrhany0
rybJgnInWSC4JlQf0sf1pzpX3hJBvxn3buOzVi6NTasmHI5rCCJSquE/SLpLOd6q/Rnw/hikQt52
ftzxJ/XZigxc5krVk3GFJjrFX66eJGk4PZIgnHIwkYyX2BipKxaqjllgmzvHJlAZtA95MGxFVaeJ
MUWK0ZumQj7XGgPuN+C2bBZNQMR9ea0FTI3AO3QhxYNUWSNh+YGK+ArSojwr969hztqYLZR3BLIy
L6GXwY3MZ9C8AXRd0gRPn+4AklHNYtyeKkPSC/2okH2OWRtpd5QsoJFkX0Xgii21D0GzezfYgRxG
qn3S9mQODHseYbAWt4hhZgrOV57AwVhh3DcK+efupAutlJpqcWBjiuYbux2HgR1Nradx+C6dQMXN
64PbqnwjH5+lQjUnjU1IjlT9wJ5fGIaGd6wijAL0dULfHoyg/09DWlNKaVX/tLXxKbwMDBw0LCpe
7MMn6d3DhnH/PnB3iYPS6MOLvXenYLVeZmoWXum8fgA9dJAAtxHjXSYuGwsNn2vYQW4pUeCcwopp
Qt7HJBhxZpXcefXptbh2PwWcQFVhcQQ7n0g8EfihHsZF0NfvVbXSAv90eHBRFge18KhwSSO52PpT
fEtrZeVl+cEddgTE7Ks1EHrGVWcGoKFWTtD77d85IQ9Bd8DrWMw9BW/LFC/M3ifBeicHOCKysb1T
smKIkMSAgBqv51I2WIW6jDKrB4omjOGi7uXibCUTFF9BhXI0rDc14gxO8XhC1IkK8JVmhPfY1Leg
2/tPy573EA/sK3GdVrGgJuzIoGT9EY2RGk8bb9ld75nYWywoMci7N1s0GmVc7oZFZGOqDqTX0CPt
ZbTTVQJ0RGWPpDWL5qZVV41Rhk3haBcaqMySF4GLYWi0PLNXrq9ATCsoTbXw3+E/y+agwMCkmBO4
LQsORJD4HjgPRgfMb9s2QIQgqvIj9wLEsmpzvC3jV4Bgi+YdfAopaxNuiOPR86JiXOXT9CCiexEE
nJXVn57u3r/EsomDrTxZ7GursZxRs0xA12TQNYFIkmEBDLHAOMpiWJ9Xxc9Frx4xe4Lee8q5lSxg
Wq+bV9Sco4t+BoFQpeh+3P78GomLbXgEFgj9vgTknutGwTAkWqYM2Ex4GtAgvpE5V2YtfH3er5z/
l/SH2e4xE+ckJ6Dt23d5oU0t6sNwSrEQsaNLMYxvB6eKBsO5virWUIXuQieZDoh+0qirhVHAUUeN
XvtaldUTkYZFX730OHPUBlyMRilRZjDcO2h3Ce6yUkg5HsCaPXX68UELczSg8+GaUKRllU+gnBC6
oSBuWECCoyLC3Glz2RnhfPtb9fFCV+LGmNdM07Z1E1Rj1+Ss7gZfYPeDSXn5ZYHqKRcBsOoyNc/i
exLxScqwPo5NBZOOLtTVZ+fi2eXSULAng/xGSaiXz5pqclEuXOB76y5DZgcEBPuVq7ggzxmrRdgN
jCybO5g1P8HQrMxGKxGZBu3m/KTBuT8rlPXneNMGjB7A0wh8yroQlcl3kyM4f0bkIBrcEuDAIJmG
USYhjbv0IQ8CSbLbAaZCDtBpfkQLlJ5J8AtuEi3fP7XDwWwRL6CWjgKEWwXXrUE96q9Gxi0LL2VA
10m5MbJ7V8X6fTSYlX3K4DCDo+FYO6EcTvZICfWdOc7KO7V+9TbKxdi1Ged1JdGm6RLqgfq/ZQ9b
bgEFrCdSnWUHflbWWf8M0EocF4dvnOZPCesQzwxT+7vIugv2NOcmnQLLrxo0my3NLVu2rpqoxmsc
3uiQpWX7ErfKGNRdgGdjaZrHUgTlwTVHlfxipJQyFzh4imYod/+RO2tyHbApp/1J+ZBY1RWDm6QH
M7n9igLPjsFJI0sadrlUPkqXkuDMp9LmBhmG7Xf16X0JMvePejjmxJEiTZXCPFSxithakPRiyrVG
8nsuOldBa0YYoXMgJA9CQLDcDzI4JFH5PQyaJ6vhgwmzF2v3QjyaKh4MRikmB6XSpKo/AtYiqbyz
JipZXJqd0alD5GcAQPPBXHT55kZgTs82RUm+YhotDLn4Z/I1X0HJALbWE6gjbzpbNe8J/fbHLPTK
yqoHKYsaadRVgV5+w1uU1VjK4/LPHS5QKNqU0+JV058AZJHw6DSsC6g+HWTH33xlmgxYUuN6qNuj
/QNmmXaqOzjyyAVzNDZlTTWlXySifIGZFa5c4M4ltn6ZS7KmveC2P8NZhwxoiMJ4nmHqiQSIrSmI
G+atSxXj+Rh0j8tydUuoTUiGelPah8cGbFqxcLR3CWS4AIHb8798sZRGlmKGtgQ82lP4pEl2PyQu
hfhQMKdN6q6OtrkfwhtYBrW/FQchSniaav6Ndxl1bLxCRYw+Op6UxeVmL4IFqrC1Xhsc2B5A/s1C
LjO+MX2WvEmwcIxyCIpMym1TKLYs9XLjEAOpUlCPRrQo9oMYFJVl0mXGiM0A+/a0UwFMf4nvmhJ3
3X4JZB0f5nehveZUbse0YU8/9f+avGdjauuCG1X6OoRWSkFc6Ns59lzjCEX3ELPcSQXbogMKvfXq
QIBxLWcGKroaoJILl5vXGVRTupWyXNq2Z5fcXSGJ9boE3NOGntX3kY1Gbh0OOP1rmc5fjjeSe9PE
BOWlB2HI4Ve7cbrdH0pkOSoesD1BLd72/NU0rG52RNiVqYX9t9SvBeBrSV61cROREOhazyk6Eg4y
z+8ckiip/4Lf6UEKevpVWINzVC96QM+PwI3HVPDwMCaMjBsZqttRI+EFQrZ4lrk3Wun6yD/ebn9M
tNHYGr0tBiToI7hrGZ0LTJglO3FzaVdvFdAFyyUDm/pdMKFdmdtGhhexoJhFPTlA0wa71qjXgNWh
0NpIIGNNi4QO6e5zWnkQxKqZFl/xjYXfdmE9/uO/gyTHaJRVCv7X3Z8QKovPuRQFPCVsuQDoT+Pi
90uKXa92O2tR9ZndQqAKsbhiyn8tgzDc45ofFQlBxtrVaIkwf0TANf7o27NaxMhUpHY34t+eFADI
vDlDk8kaJWz1Yv7BV5hJTg59PLRWP+P//u0NGEXaiDNkpnKFjh3LyZBVUpEPOZ9TLzvU4q0icR3A
FBhEfiTmtBNI8b7S/Ibgda542FnvALl95vuy0RlKmzKfLSUXLOBhSxsjDn0TSMgl/ZIMO/rSHeRs
czA/Wx7sgsV6bTcmwa103oLv9MmphFTrIOPDcq91vvkgkCeEOG0nLc+Dz/gzxOl+bFC0sM8Sl1s1
lYGX6mcObkfYb+XEqc949Gt624Q1dqSS10zOwM1V1nzlC2GE1x4kenuaAOgZYYcJrTB8gvjyNZ/e
0cFYn4jrbGVVhBhi4LObnNlh5JpoTX3oUTl4I/HM3cSz+OCbpfwzGzitzDBRm8/TOQGecQVw3y7v
d/sU8Qm/mIPmHAIIAEwL9PmfGr3jRL2flfB2P5o48+WF8oqos9J2TB5BCBhsChRpdhWzxgLmMrr2
vsW5/skls3VrYjQtp5v+MSa5HQGuVcACLTZ7vna++jHtiZ7jx4Rp0h+SW00PZzD7EEKgvZoxa18F
HF6hjRTWe/531wGg4kzwXh0sEgIDREK2ZzF/qmokmkZWq/hh02F5Tj5bp3U4xTzyL/e1/zrbUVmL
HrI0sZUET2HKQlXtuXkjboz9LpQjz1dN3mx0ktIljSg3FqRbgo+cgqEIRefEU6d4LjV/XzCSWgbM
MO9gXF2dLSDTAIwBdtPPDkvAhGHd6ndjJzhlDgzhUpMnSNjxo8F3AwMJDaWAiyDxwDN0J98CzbZI
ZnEfIpOWoev8b4Se7Aj6+fD82e2Yei0gYczw4g69MeV2X0Jx//RT4/VghN3S6XwqWBuHnG/BYPUg
y6+PQMdZlzddwfOYHlFa7zj+tHfPr9AHgMZ2V+6ANHygrsWtyQ8MkChaYmcP1LqyTa+A93i8rRbK
Acz3QZtSX0k108rp6HNc5RLiI8s0TAcARVFut5lFENG9SUv+L3ONsO/bg57/q1d/nJLhSiY1InKr
F3RqM8iUc1dFt3gGbbsrMhkPFP9Dill10XOYlFYx17oT0txW8z1XfZSL1dIH4kSUCb8v9bcT3UG8
kvlMrPyNeGFqkSHhm9f0Fct4hoRtqioYButFXUgiGJakYbPZz8VQzX81UWAxyTMLelAEer5CndiU
KQ450YSBOg5ts7ZWUjRbyScUn+lVumW1rkVdHBJf6l5TX+/FAkZb8DxiBWnnYW8KnOjA2Uc+5P8P
YZt5vfxiHj6kmYF+mFFiVf/19dwIghdNgPHYtru6r9v/1Zvjxn7sj7prb0R0FfXesvxVhP0khblK
jzYqeZxhq5E1ut2p8GKNRsWqmR2ob1OgjACDDeoxE/NnKUx33lgxt/kAGISCSnSI+zTcrsRFzjMK
MkfbXvLMFYSwSy/dEsDMHzPZm06JfwymFLeIKBbJGVqVf4mjM9wApA6DfFdPJUqyYDZxGnEVs8od
i+VZWLX6tD3x/U0hYoaCfiakawwMXX0ERdihXYXIFwB5Q/FYZc9ZQ0HIbnxfeUktQJujep58bgSw
vO8z+x2cDI9P86OEreQZMhFDAPE9rGy3nU/+gcQrwrKFctezN9ByntOPlS8JoXaqmN5BR5nDPxqE
4mZwCihY8qVW2KfK+xBlAgY5zj1BSeipYCSIghObzk4EmhFVLdCTm+oBlZJK5nf6srgkGxpQwrFK
0SgcVrbKr2hFx45ulzgHIR0KDWG7IU9RUJ8a+Ecb0Bzm6Yc4bxtbQXB2YhEAkALXsvmuBNaSG3jW
pWU2SAjr55NqI+Ki0XMplDiokc3knyjiGgl2jffveeGd5lRZ3CBvRUbw7XC9DuxcXpxGuNxY+MWp
eXanyir+GxZkJ6k6ODaRC+KjDt1aLUn99IuoMsiDp3ia+w+pmduvZtL9PjUR26gGBXfRVA2gMLtu
gvWgLpu50sjbvncBrWU88GJ8rVi9S4yVO5nd0QdL28xKCujIsMvPAsu54kL6+3qGB5WdISS9nQTP
8GQ33HQijbQRK8XfhEVw8nUYE8VXnCW8l7Ha7aYef6ph+0DiuSYDj6lQhaOdifBfGR4ynp7fKCXA
D/7mlvbVgOErf97Mj8Ue6O21jNoYjev9WqWX177MgqvmiT0KMf2uLZICsjKSa12Twqppan/KIKfR
EMxfx10UpdaS6H0sfnRoIItg7YjSVVzALfPokIUkCzns98I1AWrsFuaP7LEWJWMJ2EW6x2MDmYPz
6DPIY7N/OqbWY3iSTv4HEM00W1QZZazXrRsxrxS3aSDYSl6pVIz4urhiW+K0Vj99YK7VwETyN70z
ypNlUmzIrbQwRy7DJOzFveLzP5HLPWcCR81N0MRwAkD008lcGLuvoV8Jvl6b+uJoylCTVq6ivIIF
Y7a2GMi6n1H1ukJORRCJi8TykOJ9cDVTB9U27OI29gn7oFAo6tbWZRotT0Fo4bDIFiW40dOg287k
5Sy+1xCMX+sAEqb8Vr5vKtpbryE9mFcQ4DBKmPp2OkJugXwkiR7Byku1MJSaixfczcSLqHJ2s3bS
+L8GTK/T1HsiqSAW2TXCstfXbEo+IGM4ceXgDn/Bcb05SUwhatJd2DDzCCu7nbCpnSwaT373Rbv5
0porPkBr9+QgJoVhEFMEmk46OMWwuQj1CeqFOfpqRVBWXJMTwFsb1fD06D2wwu/apSoSITzgdHkA
xNsr9nKad3eZB9hyH9kNJJssbyhOZYVQNcZmo3crdh9SiofMJF7+KczvTZZA5UMltxETI/7RM8Yw
jtEwpjCR1Bn3sZ+F5kNCXuoUQP9DxfVZ1sDdThskIFL0aAUvvxqmi5PobIhYmVG2C8wmAO5+axsU
VMJhJmzhfYNKKT9Pviz4zxIQ9xGc2mIY6AbJb9OqkL/KbYvW/VtPer0pqborof/zCFjSL0tVN9qN
98Y8esepoG4TUlzKYme4UDVCPUH4o6ezFV6y6OJCbX6/c7Ep/be0YCpr+0VRAC5QR6DGaYGx1Nk0
duPShc3M9Y1QxZE4bBnjy2xyaGaKHk80JY30cjlLdtl60O1kstyyFugjNJLFpZF0fAm4Is7yxA1J
oRY3sZ7uZNtOVqS3sV2oM2jvYoymJLqobjxTmAtQ5W34cnTpnxqQD2O23Y/MDLgDbQqNy3WHR7uY
DoKeeefFT0uuRJ0jQnL3dyrPek12S6bAPNU1TdKwY2UEcWtmvRm8Z7w+bLFMbeNnOwdeDZ8FOoMJ
SA7RSziUuAr0lDAPlHXfTSrhokXm1w+inMwGRYn1At/YqqSc5OR/qiVL05M4XBvZ9kHsILP/P5oe
fN5R4x9VVwJ7Dbp47YORrhCccpurhRb3DMQ6/88gUJiyJMXGGihDtbJE3th/IFYvER4CpQuK73cE
/xHCVjBVIT7+G7baXWXi0K7F0ifg4FNe13zGMzv3pGuVMOZO33j/LBkx3gI/nIy1QP9oGH+CMBUP
KNrPzdqf+3T5uBOTeIIUSB6lNIANUmMUkAXoP4bubVwqtO1TIle1p6/dmBj24jTw4asqPuVhoHTX
15jOjSVixxc6lALOB1lgLSxu1sm9Pbt+Zn0RZR16SW8BSeGOS+38CZEXOg1GsYMAqpi0otkJwLmp
6c81IMMsv3RQ9uA9BpeHGP5p3I7ClXZovwCwau5rl4BvbXM+pp7Kz30N/Rzd/UQ+MUtmP+MT/efx
Z+vGQDiWGWW76+Cr/DTG+9Q0mLc6ISk3wKXkGn5utxwBlSEuGSyfzgIzEopkyf5iY9Np6vQrVx9s
/1zHJCbCtFqoLAsGLJXblxiTJ+fzCC/1XZQq1hqUUY6gRMYxQQXbUuJS2+9Vm0lWssF8p19566xT
VdP48XsU9qQQMNy5jpJ4lR1bSk69nx+njJD922B7Kmm8DrXnSGvCpeYiUdudGXQs88aGDT5na62c
gB4E2qjud4+tq6fncAEquMubudtm/FlmJyUGEXtS7/nQ7h4wBfMk70XUDE7bMLilZcAlO2reUIGq
1zqmlv3NOmEwLMDWo+4g9vjtSYljHK6yNZvtKeWnMYeyDuFZqm8+WLBh4ZIdfa64sN65uCSIfmVO
6R6HzK2daOwHtQcdv/qqMbGwIyiUF3vwBVqE7v5lcPI92NNJuvyJYxqfZl2BJIvx35Npq7fvjbMU
OaHL3B5Et8IKk3fz0G1xC23eFe29l/qqKsl0GrpJ45xWVGTVgU7OkJ01EsBCRYj/SeC2VxooeiCt
Y048cI7ukIDIYsWFhz9W3o/L0o8Xhf9vT4toF/xmjrjdFqBIsoddH19J82Xmxpr3890VK5XYzOVj
7rHohd8svq2DHjAe/THcDfCZlAr3UteqSRY2FoiuEahsAxNGzefS5dA9KnyA2zKAKHw6Ua00TnRz
/EdOFxJXRvkA6v+sghV5Hc80sygrYc1QRywnV2mVuCrtTE2TcmV3MlnYFGs+ZDpEaVTvjubDvqjJ
WbIuUhUj4BGIx2wgZcmKcfXAIO0zQSOx0Ov2tpItUOhSLv/uo0so3Jj2l7qKPNBFfvuWP7PrhTXY
1RPjQzseNtFzyjCTAg7cin4ASh+QB2HqTdvXDdugAIN+bNm8RPZbXeQDoVir9AaU1/9PrqBGg7fl
Lr6GARkyg/JI/k9NrT6pfOafr+I1Z/qLuYWqktaMy/eTWM5K/cwqKgJL2+lr6iWRsYdkXyDbGNR3
SK12muJtXa5JejWmHDxr5Wk2kgHPzQQHjYUeQDVtnRjAii06lhXv6f8U5wjLOia0E6djDLtRwbb1
ePcAakhUFNFI8Ti9wLj/xt6le8CnZrIBl2IoQ3qm+x0JZOiQ1mjzVXawwJsC7GgqdjYPyOfJeeqi
jp0ky6VN+cKtCOy7Y7cqTE6ivPxM3Id9yFxZljHamX8jRh8T37VJB5vfNOulwkhAgryzoIQndvU3
x5HMxVKL599hl3Re1jnkecqCcYpeMyjizc5rNZcLGiTvI0RpXH3S+G+cOPCQ5i38A4MaQrEj4fvn
uSNETBCfHNoHoNIvaeQHECNuTRyfwBSGegKvfPC1H59cvMFl5VyaAWm6RPIcYTdDHs0rsr3G9DDV
No2NhHxjITRCGK6/LgZC40HEgXXkXy5FA5XxrF5X/DfBH9jaoyyUrU0O8rSMnF08tSFoPdmNWQGW
fOT2QiEk2CeMcqwpIsixZv+AivP+OEe5SKfsr2pWQYTwy+XcxQi6YXr95ecdIvd1m3vo2XOpHz3m
o4IFmneconN7qzxT2pgOMoXs51EsbD3cWHZKpedleNhG2pE5j2lmE8TY/2MKUSNFO5a8G3Z3OLwZ
W+Gk+2WSyHiPr7+WDGEHO5FKYlcBLh2WC9wWo+kD0Ajud9rhRarojwAweAH2mIFArI7Z3m1DDmj0
eiKxAmQ1ku4UHni9lNOfSqzaS9ia0QDoaBe6W3+xOgiD6s4npArCg9WM7yGf8yV/r8Be2vSTq+fQ
Og5EZswry9/AyG0cR+kFW0vuFXz0hzASUc5xSJnWGA87sKjH1ATZ+6zyGT21FUvj2dzGcf2U5pRc
m2fByoepcDFS9osJYkPkTTWOOV4riX+CVcahepddJfTucaaNkQmQU0KusifNGI+Fu6PzCVaPF1I2
cuOVOMv2KocpvpwuM6RzuOJr65vdQUz1TUyC+XdbE+b8BZvJwC6ZSWpftwfo9b6LV+ojqskvXHYg
fCPy/NVTUS+fjRQG22kzs1wFmwi8YksjwZDTuQRcleux1k/z/vKYTfVLTrXszRbaxKzJQxk6hikH
2nd/7bTkQkEmB4k4kny5vNJ2qvbKrhpq8/Y0gr7+K2S7wQrPzCGpN9kENI1qBJgZYFb8de3/Wjys
FThi+TIpP7Lum4UNSjJ3YYAecOaG/C+kw+qsmad8QGBgkAbWX1KgsNu2dvfgoJ55sGi+DSrTIunS
kZBwtEWQYq+P4mxgS6AX3sZRPyaQrxJ2clHwyvvKVKv+/EcvjrFraut3kO2HESW4XTlWRsJtQQb0
AGmJ1NwmK8tABgQls3TlBPEcfnCHgPS6QI0I0w/nCGWNlSB2KFJs5Ci5HgMDhqv7vlCI3LgYl6GM
AfDP0FsgFfyBb2LrJh5kR7+T1SdBZEj/S2cTYjn86ZSflV8ivZ8vvXKgs2b4LNoEaDW88LQsZg/K
vbzex9KjgwjNgJRDU9kooEXEwYMidp6uZkirqVGCytTNZSyUUg3t1b6uoDv7bxCGy+70l/cGYMgR
/hc63KgWzb88VbK4XcKPRvsPvv1wrbxkz3JlC0ReEpYxJHSF1lua1EjFw568XX5Ai1mY+/b7361S
uo3jR1SJe5K/0tcGr9vzPA4SDxTa8U8feSYP6YQKW1wQ9GKHmsvR+6QNUjuoD42BEiwebPnBSoSK
Nbe+5Y0ZoBRM07jz+k5r2qxhzCpJeDXCr0hhpfSTdcqsK1NiuAORNLNxjX1wiEXf0HyqDKYK031Z
embI/pR1HEwb6lK0fEFjMLrxWsgNd8BmaxtziFeDPjitr8YArZNCGsJjvqLobxX83N0M4lYjjv8E
owX2XB8XG7crSRYrHa8UnKoO2Y1ip33wCqG9Xqlwd+AzGfmV/M1uwVvnhJ4ueunTCyy62yvtjLVz
w3gqYYBHNO3FOM8XCb0SyxKA9+Fs6tWkyVrzH6DF5onls2T3glwntkmIVAh3dHWYxGTib9Ppo285
uON7WYxRn3vbSe4lj7UgB+Omv3jaghMpgNdYTY3cN1SRm0AqF+X9cTM/Rp+D0JrjAAq23xqNnhTY
nERGAiZc8yBfGfJ0Qwi49piQP2+sd1V4qBzT/OZ46jnhL8nHDEs9XGNwxjwhwX6/4XZrD5XU+n5y
OTV6Xng5iJVUmOg0vn96h9E11GYlqUiJOS/pcPxiqS+ceNwFr68tIxihub6KPZ+x+43LzSd4V3+R
p1kBRLJsLOKaWArObMEJOSe7eC2GnGMMcT0pO7XhGvzf/tPFGsdPbLFWVZWgbLGHbPsiY4KvVDld
nixBPNpgSHdR1mz9zBuFM2p2sAnQ2UtWspUqHJX9hYW3hDVUbsUmlOMMXyluiYASvYPdKjsA9WwQ
hFx/Reis9/7oI6ZR3dfWDdOsyvs6fwzfo+ScEVfGQOSCEc6TtUapKcFWZmjVk5xYmD7SFrjk7H7q
k+feGlGCyMbfOv5W5tYFF8DORw5WilPt9nMOWlmiiVaNDrHzPfS/JspAZ/xci40qFw1J4U1gfbgn
zE/VBssIDNp0gP98UTgyQ5myU6tr4vWtOK83CNtO4dDq9xQU4xszWnVSSBhFxV0vTAWt5fpxZfum
yrq89kJ0lch7U5NvG709KEtZsm0VDeY26O+5b7oL89qcd0TJjzasdnAhoh3g1pkjYTG3CZOzOMzQ
nvK4ODsMSFNwGvFc0zZsShGy4QDkrhV9ZkDCuTzWCoRFbWEjgkgB9g1rzwHdhAoy2dVPqmG6A6v2
AuPp6Sf7r9QfR943xIkMIucrhqx0wbAl5U7/8GjwvrZG57H8o8uVoI4sy5xij7QxbKPwT+GWacmU
3ZqbLUtHA5L1IP/OXbnbBOmqMfjSQAF4Sh4tX220ICYc7LlQ0tGUOHcbG1Y3CxrFtGpskQI/bH98
a5BEpG7odK+O/XZv+whK1IdE7ZdZ6lPRr3VeMSXcUes/NJub9CS9YNZILTRcdSfGmNRlQ0FJrach
+Q8nqrBk2UA/4SATg49CvFQoU1DxXyC6BighIyCeQMiS10rPTeBQtN15R6XhrCIw/UV2pA/f1NFV
GbrQgF23oNwD+TBZoZc+jZvAVViwjJn24QU3Kj0WykuWuMWXIw2W6fqZmlQ1gbczJeCZvU6R14sR
BWxgTm+v6MKGjJINN0QmzQmiz2+rJHPVALOsCU3Dk7PPgeLbpaxBW/UMYkL7U7HETRWJjVCQbbzf
Wp+/xuyObcFq9N5vWyASYxe9Sk5OwY8SP9n/UE5OLCmE5z6phuUw5Fv9H3P/BZnPl18bEC6WWAXC
YSRbQihvHsXXeL9TpjhdRspiqKukWUCyntcEuH2pcB+jXKx91rN7nuJPr2M8Tafo6gseEyaTox/w
TDEWAmpUuuYRO+SJI6KJ+40orfxhaoJcugi9+BA+Xxspzyv4/4pQQlSikxtDzsgRGiq1kNaEkHZi
WtEjP/wMywhJYCakEXSjegiazA3BYkarf/0r0Te40XfD6+jNgvyqPC4tpA5T8ha3989GrVjqxHWy
VYhbSIQfRxRcPRysRjKx6AG8P96BxEug0n6V933rv+UdXKpWd9kQgrtrPfam3trle3Zt5ZqGOSuY
nIBwLMTNsDymDOd6buf7Ok+uKzsnXsMqfxD4MYmvtWRnNCiNFr3+YlNpRIttDgPH9CP46MZoNZEZ
zCgQx01LTDEX4FW2HurUf0BBbk3W676wLwZKy9gU01TgPPHpCLSSJdIjiV/M1vRxHNUXdGRU3Ni+
gN1nH/TSnOaf4NvULKHKC9jOcTAsTDRQgnQP6d6coryfbM6Rhq0OgnI+APMyCxoEXVmZHl5J9KaJ
BeYyhbntapdaeMMG29LIdvtC3PmxJ1YgwBiAhPaz7fRI9+95bycP+Log9tFL/DjOTuMdc1mfv48g
u1HBoD1D4furT/U5b/gEjaPBgD40PV/Jv/scJegZVfD/KV4UkZgqeO2vae3oir/Mn1xIeGIvUnt8
KfcllEtnxhZvyMfHtMSkY0VKhudGOUmK3mcHHA+zEte654vXZLdVpoLINj9yB0wbsvG5bG1tYsvC
hdLFh7Dl65JMl4g8uafkeFauMGmDFnvFcuiYKgHmsUIylBlageGXFqdSwm6GfvQFZmcqaiPDp8tf
B+/xhdl+yDnIGPBsc5oupeN2EbUOIfsT/cylQkDOkwi81eD7d4EGeOyc1f8m36sljrm7BBRLX09A
zzmbMLzVgtfRTMwWlbB3S7fVeOyh1k760VB/KXY9K83cvCUeNPL72gkPonwhTaLTpms9+ptWQyr9
5Lp+le4JbybSdIyoIbbGUV0+ylF9QOE7rEx++Ok1hS0bXmGgmIKPoAK2NH2uXamgmdFtwa6aZTtw
VEZKylaTXgUiNEympY/BYQrle/2C2mxDbZnD1bikhC13rfvWjoq/GE1gk5++U69eUSQ5VeEdZZBp
71bQpHzkiaqEnDqNwlAE3bxwH1yw+aHU7t/p4i5VVDIe87HYJ6E4KC/HmizaswYPi7IZd0olgnV8
PoHkMl8q49WJ1UTOGpbNaeMCbPXwk9PUB091nT0fb6Tgo/bcNfaoCFj2GMc033b0uiT6ogkML9+R
sn/s2Sp89CYx2Sbs8rSKRiicO8+NNZXyTYJTFLU9BW4URNn6ZdND1xygzNQWYzoxW6Uh3/Ei1CO1
zaxB4bj+fMO1P6fMe6pce11pgeO+xCD6v9fSGAsbmxWgGFmgCm8WiQ88RLxlHYx4Z19tWKPR/Rp7
j+r4flAcMk6hVNUzXydKnFCBiQe/AvweDJmcfmLaPu4EBZjV3To7s3L0HCvDQMUajatadxeshueC
QjtS4YQNO7IQuG7TjBBrPn4l8vQI3AhFFIpcttMdxkwBwA7TEMTLAhu5U4azdOjprJ41VlmS43Ru
SP9gGuTz/CPwZYQeOGwryitN8sQF2jHGfWgB3Wqkw3EefPlwCUy25QIK/6SrqWzi0PCEProATfIy
cApxFJPC51CTIZE/1oSYq/0D7z5rfUcf4tVwiL0kKLdhleQUWkayMQBFaoV7IlB6OJ4oI8YWzrWs
wfXK2LwaAQjFOFnJ7Ril2air/lvwthHwxF47KzJGm4xJLL8dMN9e60dH6aUUmtHteWtlRYAc8DKH
TVdYuLOVLARnQlBSAkbjvuHq9bdfpc/33tgz7qCE8U96QLs5eIB8mYyYK19gZ/R1N92RJ1Scsmyc
Otnk6Zdk0fHrh/HWUTAF4pORdwA33hneOeJH5NtNzqz1d18/hirsCD4mE2SmSKi1HAJlU7iwIUo5
ayFwPlPhQLamJBP6tv6OVFIhN2h7iIaRTAGi/HXU4VI6dJ/HgFATggG0hO7f1WI/i8pZhEbP9LiS
DaUmaKkxM43373Acj3iN8zdKWVgpYQUDqOfZAeR0G+Zlfl2hY2kNQGR6T+YTE8zszApPpmIqQL0o
D/+dUzPRlXk9F0mZCXL3DfEftHgKriUj2ckaeHG5CfTgPjMVnneGGH1TDHetbbuxEwazECC497xy
uCML45SYyoh0aILSJdFWtiKGq6IcPKK++G75OF4e8QF8Z3SYsuHWiwu04/Gzqk2im5LPN0SdSVQY
MdIY56Uyo/AN0NVSMwE3e2YiOJeHHWAVIHKWmLhZ3Tv9msRhhLVG56iXm2ivoiGHMj58PQTmRi5h
hhuzveGZbLkdWG0VZPdXrfdKH4yvktQkzjISLw0H7xlQih7nzRW65/tUMINrkIT92bFL0DfG4ZW4
2SgAYMefgQv1tJtZYvLScZM8kTaVjyUVH/M9NiJsFewfdLg9bESy2N1KqRbzWnd/yleIxEL11lu6
yX3Z/tr1GVRypzTeU06dw8BDX3ay/eQLczdIyEiYs9kxaQn704DwqX0NOYXhWb//B+6sU46H2lMp
aNOGfxdcLgRxVDLhj0QAen/rEFOKTHuwGNhViml3XyWZBYbog0QEFMtoin6bu6kWogLZllVgD9f7
GcwGdWi0SRWFfWfKgKvDwJ2+ZkBz94ukW3VkRAaEKH7Lmr7a52JGUgCkwLHA2qMlmMOvVJIDe3Y5
LbDqdqJp/v+tZmFSHHPWBpvIBpZJSs/X8hU20RxCi79P3vv69abgPeVT2AovlDjnWiGmYBEKOulh
K6MXMLiV9RnXFOaW1EkzoKAt763oVqRdwkYZgdWwv4zeHqW5WOMmGoHMuHY6pcms89RqtJX9Gtuh
8iR1x3zWYagmxAgT1blYHkPabd5qjVtAUjF+88T53A9gvy4VDyMu2rPEe8ya75cJOwJBUpMz9CrO
4LrZn/g6/jUhX7AAyd6JrlErfIB0sMu5Hrnd9fyhXc/rNRFqRfDkMUw/tDwZKpW57pJWPP00nc8Y
VLqFLmBPbl/ZAewJ7sOmMLKBEK6IYM3KqfG/r677Qy8sKO5FZCFXniDRC7tmR4BWVHzjoHEcCFbp
79tYgE3v7qKiZ42/+Ql10g/Rnzqq74TOsOc97ii8Bouq5YMDOB6e6bt8UVvm++dqMOEe/wrT7U6j
mWnc3neBN6QZySlHh79jKLKjFNnj2NPE13vpe6+skIjsdXWuhGjpxzDec1rg3DlckiZHP1Mjl0fS
iqp5tJ30uNEDNirJhnNnpAh63L/bx4EKdLJdmfnqYMN/KqG6gq6Pahin3VE1Y9JuL2FU9fq3OpeQ
D81s5dUzwKyax5LCDmgjAIeL2Os9Dc3A1SMku/50X7lK5v5pH2dW/Xzw5Jf7dvR9SggcHLxAMaH9
I6UiP9OF1U6h6DwaU2riWwFxCmCBsCIbn1epJgverNUc1th3flEwdOEYr7ok4GY0lvQMo2RVJusP
XDwkOiFkdMLGD1vwM5f54EPKFJP8rLXkDP+W7iaN7MvOX3V6bjCLOwhNUKbDfjtjnwTs/L9UzaH9
gSu/+vQSZIi5MThojMme37QbgWPEmI7WTojPn2GjRY8ufFTgoRBEtDJs0dMBt4b6NMPMZZ2ywdk7
xtRpJjpABHvOoYJ/M0DlioDkSwO1NYnt2EB5h7FhqmTbFoUb+8gPaingw/4o9GoKv62fA9ODGbnF
iXLTPggSlAFiBapoQQp1s2E9TpaUNYXTPN8gA6AQmHIZwY5niJrfk5YdSa+YlcF+Tz8PyZzCLZWd
uVJ4t0odjndTevxAVy7/3VsBwm5D4yFcvyDWBvtKjHDWjBvk9YvIBobw/GEq1E/PE+fS2wotPW+F
NFRmHq8umdEoVHFj0JO6qRUqBgDVvWyGtFQEUeK21JUpOpEM6cvZye2931mbSbpD04fWPznGguGw
1n0MfHHjkKR033n26N2UeFcXT4EKhKhrqJIf7X+SAHXe4EBndxdu5fl25L05lhZOSWpUuTqjXz4r
JalWnuZjc3gAbXsHrigd9s/4FtoOUDMqUt2Q+pjNmh/9n8dmJzO7z9/wOlLG8+q63iHuBg3RggAq
INch1Vaj0jtbzMnZ/M9AtZq+1kpEoCLER/j1cUVZPE6VhTi5ixNYY9dErBwhKF6NwCyBnhywRj/d
CdqpeSrTvMfmqTySEWv4SvSgE2vX/Mycvn20brjUqS43ITDGvjDNPNkU4Sydle4iyueQD+QIWlUg
w3xgi4+myrfq1DWmA5zU655mALRpjVq/23/VLoe/tmAdcoV8Xp/8cXJf2lhjxjK2C2OBbzenaD6a
CNm99JihZtgPHXv3FY/AZYueiE4/6v+hiE4kqkvi+BXWp0tnpcfL2aqVD0jh4HF4UpVy1N2uSPr3
ilILiHE04oQI4lXlklHfDS0gCyj3vr6rrYhrQ4/VIx2/aqGedn9eWF/F+0bZ9ymyCEOJsLFxEhl0
/l/SF3MQw4CKCejYFivKzi82iPmGyvPvLiJZv1F37WS0lo24Cv5rSAkS8y4rBukDHXglhvDA2vte
zXyFPOl5pzsA2k+6DblIYIL5Az9T7mo8oeCqNJiZQOfpwGnB+2RTCjl0T79s3iEZXUeBwfR8Taqp
38w4FFfNy69zM1EDPFsA3EsfW9fJPAUSrtoR3xNpudbnB6kNxB4VJz0VVLiNMxAncQSTZe4Z3MmP
N/uQauW6vFjg5GnC0RZUJ/T4BClNoiXNBNYvko+jkoKC9lInq8Bzwu3oGdySsJBQ1PTCMJywpqfy
8Tda9NLb6wh3PikWFeiJNHuOJ2RRMHXa5uWjlASt7y7hxGymiGah/KP3M6hl863+gS8Bz38Sn60u
P9APSfOv0EeMIc1dLv010rztPv/qjr//VJWA8CSJ7eKMx+/gpfCfpiAQ/Nv5CcVDXMiGhZN0qbzw
S0R3OumxK/LKcg6AeY6NJtbWl5oC+U6rgIh2rlSETRdMb9vswWe0Atlhm58swvQFAmtfL8wj4gXp
q3C9w4/ujauRVmK7FnM2Y44Gtel6spD+tyINgogd2HOm4iIjEM5pPAEYnwnII1wYvRM+9kIvXH8c
YaAv4iD7Q+XMfbpFU3Ms9gYvFNVd7Habem+PP4ndbA+sn16cJ0UBrnKjJWQzT1dlkQgXQVU/sDiq
0PsmzM+QRQc4u5W0vyd2UEbyTqB9JuKtMePNTYKV4bDvohL4kekeLulpog9TfUu+5HacGNAv4UL7
xd+/jfg10uutLhCJxSH0OKtb+EnX6n5XtiKkSXdbHp7R5R0o/JjHM/kVURUtFPPCT/22KTD7h9iO
95RagCEdGqaSJo/I+OvNxyutB7WrKJ5hR7aJ/lFoVD42UaL+1YPVrypqkdYdr5405OjVu5c5v78c
HsLb4buoqJ4tjpaBG5o+JjbdmJygLSQu3m3N2SlwCe6hZAWs+3crJWJqz+9Jrt57hQg6edQ4kjTu
S4n0diJyPN1J1AnodsxwBCMK/k4BbCCxqoS0+LmuSKL1aXnzwJuhHm/DpPkqrOT4tCm3/9ozFT66
j6zQdANvNs/hTxjULU1EGSLC+xz05R71VXRl9RsXljQYD0msvyRhhDi6ejLpj/3M4QLnEnkZW2s6
QVr95u/nMaSQiqWFl/iSvSFofT6RVmoBgwYEJTV2GSv8k2M3/vF9kHecwmuw8BynBJ5IvlTctKsf
mFP+0QcBEDgweLXaXowpeA4Fo1iBDONjGuAeww3VOrP+870HxD+EErx6hb/WNxulvgeQrkWDlMBa
iePxOiBNhOkCZDz/K+GYMQbNenxzUjwYdQgKeIS6nc9rz0cZtlsvmjrcjYV8R+Vv+wnF4TFy8yG3
Yuha3OGbTEP3jd5fCNdzd59bDpl5IlrUynJu2U+C73BsN0AWGijyOIeaHu92ZwkZJdRtswfW33WV
FfPxQyZ+hGpmrbUSZiDLuVQP6MuwC11BaBwpoh75Nm4w3FDesjNmF/VzeEnd9sY7Bxt3Q/euU8Ox
cgzrggfMhFXd6VnhI9QuuTxvFtSNbfEnIzWQprEPqO9q1rqhR6JVXGFn2++iV/pMKDem4CjxsE4p
YLBgRrGoUX12OJf8Q1HNF8ddI/giqSn1jvWAUCH4n+Y2RlbIAMNtDm0OjHBa454Ee2bmIk4If5f9
vYtkBY4yblxUp1kL19Sy5IW+zDCchlgF+oKD+uV7nIwY6CNFIiOy5bLrHpU549a+CSlES/agflMF
aeOeKsENxU9Wn6sXXwaro/w+ND0AOsWRdt5UItEi1wpfQDt74PgD7fTKyK+vlbsWzzKA2V4qabWm
eW6h9OJWJ+AWWqPZQBdu3FOb5/dJIPI99nEOlgmVkvBD5tIrxA+11Gg/rwWVcwq0IM11+G8w5bR0
WjTMz9t9YPbRps4xE5NnzUPA49zYo/LCqDInFtYItHOXh9uf7bc7a5W4Zhh0I853EoT1jbEoKVnp
nRsIWsDLo0tUeYsPtRZNTJbUBr8M6pVEYugyIymLITQPxwSTFzvaNm7Le8KuK+H5syt1uuyTbTHk
n+ScRDESI+2ftFLD0JeBUvg8JYTJPFDy1JACSmEync0J35bT0trLAhUKGSaWjKhYm2SPBUryM/uw
uw43MUQ8IxkXPO8mOBVqyzOD/MU1WYAUDj2P4HenSHfnXZLtGXdRzbYPQSBV8WFQ0CogRoVGW58w
/2OTQvdVdEduKIlR5IPjbA4aqz+10xlRlMGbTiJVwAqBAXQnzxWLUATusawaj5w2NYv9krnsLxYv
rft9xEc+71+rzIxKYgCu5l8ikZitAjiTtM9WZkVshEkZRnKnOwzL+iSd4+abX4go7IE4xJpedarj
CYok9qmBh1ioTseF8pqaEjGRZWy4tbSrRqfX9/qj4TJIVjgCK4bz3ZWFOPdgt3o9uHHxFxthCVTq
iXSzFxwdBmwlEe9Gc7/ogxUvwa7u4YkM6J3kvKJOJs+Lw3KNve3jcp169h4xe2o8N0RQuXGom6bK
nA7FFHw9OEBsRY9hKMMfXMA8pYaqqdmVkYqqViUgM6iK3YbF6IDYSMhz3bXrMeE47hmVrwxWVCAA
S4u4l3XPa9+ybfs9bZiiT3xxHpy38oMzYp9rrOrswaA63DSlwVidn0c6YV7gOnHxVrS3Z4GCtVR9
/arZ427HkJIFW6jfdjHPMQ4eKn3ufm2RCExK1c5Oa68PWqJ7a2bSsmaZHchwz8BxqIGtcoQHxkSK
tXTvWmUFR58LOk457cCKJJHMn+1D/4Q2PgtqabeOGvoE9uuw1biHi0TLZLDwmHdeiMlKzpfCKYaR
77nCODAC65v8jbNCj6W3DMBmC+YbsYGiS4Jp7EjOhRN5OHY8rScyK7Oyu8v8sdDP+poxK+1M2f2w
ggd5EXaHsM+AXbkfppC9eeOE30Hc2eZomnQrAMm/1xjye8MImzdH+ttnGFi462yx2wwjgYLyZAIE
OmkluF9KBMuPg3QO+RSYbc7nDxOFISUXV1kdFXlIZsrTQe2LsdbmHjkjjuL/AdCz+9rvcAAhzV97
zsns6wPUdMRIIj2HxfyTMqnkBwu4/PjgJeEXvXOSSKPgA8iK0ZwR2Pfeq4O7enYxwjycPAwRQ4oC
bRyxzQ7W/Sq31Y2EXCePWomUNdm1KpLnoAlJ91Dsgb7/C6QI/Bhs6FWZTVoI5EoA2I4FIDv7k35B
h0Vb7l5VUy979Vq80HOwkMoIXd+V41GsecAw+3BKP8PvtmQzhquTIO0RAHfdfUW8m9JUdv3EFUlo
KOXhhhGgU9jl3RgUbksEJA7wTvm9UlAIOCLbAdAroSDhYJ5BDFK/gMzITbiYK441ELqLU58Ka2C9
f4jyNRCe7sGkS6wKJgzxkg+xPY2/esL7Tq3NuhWsnc9Q18Hct40QiGE7kuxrLaBi7atnJsxRVjkc
dN8I+iFUnvGB88di3Rrz0laOnc70Oq5YHC7PLt75/mWgo+12U4nHknqjck4cVe7a4odPcn+FUOVn
rGP9Fr6qbi/Jeswbjo0yTXDDnh1keItbeGF0RGkN+yZt32gr5yxFnS8ONqM9eXCNJs3uLA31UhUX
y9JIVOI7N8tsP4GaDB59S19TZmZlzHXUmCqS81qsyzbQhQmSJPfsX9qgSGaDqvQ27BAbk8/V3k5W
4tWbuwCo5lOMt4XLJfIBpUvzKA1vVMj/7kAVMMFDca5XLCm7VfFOZvpqD2Td6HvlCFReEklzCTzt
RZdftlFwGMyketVpWcLgP6tVqS54jgKM04Y/HId8MQqH6T3qIAcrVLUGnGSVmymgF32u6HHGr69P
T06G1YqOudBm0AvfEAF1VZj69d+nMO1jIcj3vPm4i2LYcUr2T2C4yZR+JcwjG+MgcIKPxv0l5Bk0
/jZiTfKPW1aaOVh+0oFdJOj/8FOa9smFmZPcuFQx3RWOtuHpIBJpEPPIunJ+/775iGSM1l9qi3FI
KW54WP1zj2okqazvV5usDTT47hxqHpV3OY3yRLVBanyeI7sIBmD3/8NmTobuu6HGfx35U2Su1Xqk
vZcOlKr9qZT6pcLpmdm0I+adb7UXCSafFD1shFzrGnzbT5p+39+hJ4T3kn00zzkNlfGgh+8KZcWE
sZinuRAcrMH5q5wzY6aTD+TgMfb0j1bDRK2hQCSDk/lUZls4LnHefQQBjWD/BZVcvK/5k331MVbh
PBgQ5syQpKqfzluQcdjHDl7vRp7Y+vVyFI2zlNKyHvKM+1Prd6Zf3nSxo+HyWhZ0UCcVo6JdKZrG
8I301kISwsi6Fk0BxrbRU/HUIccWDtd0TufNt61z7N1s4SuosWKokBXgVfpQ60TAQuaB89PELNjd
V45afXttp2agc0zSczu9p6AGKSdC//iGhjrakXXZwjdudprTPRS4H8RInEbdG+kGMv3DwsG3kgSV
ojwJDRov8dggc9b8EqhxBmoQaFYpiHPB4cAb8yLBmW5o7vdD3lDryrkLUu9ZodbkaIPq58FMahAl
tIdYHuy8644UHvRMIc9oyE6LQIe1p6gHxM42z+Mjw/p2FyFD16zXVwdDYlhI1t8yF+CWogOREEr3
6M/pdJpQnDxxXZb/IST2yXmHMwnY+lcy+IkjT4o10qgScTN/Ew9wb0qDdBtp2YiKVixqxQp8xXCR
jyY3IlrHyZ+MwB9vOsDUt3rX2ZfqB7zqbIiKLQ02DjIrjf7554BEjnLdpCBahZpbSOi0a+WXmk1i
1++W8PfVQAwsLgiBfhUvHughUWcRXq6wVuFyLA2GeVj4OFp+jtiNgk3Tu/c+5O2dWV3VFrIc+YBt
vKsVtTMCHQ3hhGYDNNaF2abY37FKF9PLXV1NEPDkIk5W/WAkdOJKBcb7bHg0dc/YrGSkl9UUug3D
E3Ez80dR59QwXYUNHTqmNcNMxn5CADFx+6kXRwur4PKYQwlOKWFKMioL/OIrsdf5XQ99i5oRcRPi
nLFxLEhsEDl4pDP66cCoM/+aubtbtBht9Cj7ciy84P9WX7SrJ6n61SEZxZvy/ZUgRcoosXgsWLB/
cxROueGa3E5eKmYPUUeE6x8TyWfMgk4PCX8vJOe7CZRp2xMKhjHy1ua3VKH8KBxJm9Zl7DS975Vn
oWO1lyKUFukf9WuaVP3FNntFLMV8GPk19kYGchU+tmhLdDS9e+6zqVTav1ljsrduER+TIVAauVxo
vfwQSZ9w3RO0w55JxHs5kvYF3xQGYfiiY5n8TilloGVgkAv4ax1N919QGZNuZJ9lYb1Jh+0zwU0M
U7v2Cu7c2LYtthW7YTEEYk2FY/RzAEK4TM87wHQcbiW/N1Dh5tDojOD4w3+y9jj2xIHx2XSOagHL
WN0J/O3txA2NNwN/TmGTxEIC/kN1sNvAPimTzS3CHM/km3NFQ69pBiZ5X5bEu/L+e9OYHfFN3vO8
xugYujCqwqYqft4j0+sHTk6VCMmh7FyO9Zppniplof2UnHNU6tfdK8T9uUOjexq70lGyv/a0IK5A
cwPExuEKlR5q5KjLvgxXEm6/S70ky2/E+UmMtvEgzjY7u3oQM3DTwe5BglnScv+iUoVnh5fByxr1
57A6YFurEQ7NVNxdRuWJE6Lm4uFwSv2K/QShdS2krf+0Bo2Ksbo0bRFqiKl5mlmUFuXl/Rwv2ybM
6K+SXL7aOLXS8tFgTgk9NvOxg/LTVfX4qRjzEVmtVu9BgLCqC11tEzQsvc0N8hcwINyb4qa7Mr6z
ucWN+4fOykg8gfQ3Az2QkMHTRy9+xEBKwIkBFwXiXAOM34N+/ZuFFVNdYpPxjWjApLr7mPOHV+Bg
xbGXca0X83TXVGW2Q3UbnUeftl2K5c0t7oM/dnZlyIaU5YMpBrJ+pRrIbuC/aCoWIk7Z8UedEpp0
XPStFBnMLWdOFUHH7xbkPbcW2IzRlEw9LRf8md2LFbXJISb/yAAzqd3fg+0s509ZyM0XUsIEvPAW
aJcRbNsgP+5uOfilFRY4YvheSjOC37qG9O5C73/Q93awaXnnOChwZZ8TbffpNq3pQozCa6r2ehpn
FCpLozWhkdL+7CI9YjhmOqgh6mWZGDdMC1pO7A/5T9uWN57Bk5lE+cA+V7nh9o/uTSaXoeJROxRz
msR32zly2u9gd1Et0lEO+BmKgPSm8zsSQ2m0eswOCKo1BK/YIvguFs7yV0jRObVPHoudrlkMZouX
KjW1wwySMRTuOF1oWtPWKW6TlxD7UePbjy58QxfwMgcAaz6TEI1akQj4IGoSl/jU12O84QRvce6H
NbYYxhQxkaDmhuGmyOnZBEOXks5/4U4B7qx4SxUA31f2T6k7856E1hnG0aRqDBA7C72g7GOoJj2B
4Fi6asS3bbswj6UgZQYM2Im0r5wKwdfdivUBsRdrvdMveXedDZlxay++oIFb7sN6+b9zC5M1ekfu
5INzOov7/OlFqP7qb+qk5aQDkCkuYJnlIBNcxyw0/9UmUaUFfg1jF9xmCRUELLiugI28idHiAYXQ
Pg/5TpUqxFrLSPcMYWQfn+VSpG5F+s5I7yXUjo6VDByUe0rZjyUy0z8H5qOM+dVVpyRSLwgYI873
7B9jwEU4Ucmq8TQFQQ6ZxK0V67z+HA9V+EiDD5Y0JqlWkVIkh6GbXVGjDSeVBaeaxIFittA68PiZ
MPUwBLuUCDgSz/X9ychApmFTu2RWVSfB957GpGZG8aLROVCLEzJL+V/48QJM0DuEgeUHJLRx8Pwm
C2SzV1dP7HclVnn6ptQRY2K/Na1TueD7nT2lmnvu43gam0FiReW4dQg3zJ8rWTl9mrga7NR49QR5
I+dJGCrF3VglndbeMZ2jrgldsiJiSg8cEpNm280VCJu/UfzMV/kCXS/eUGFzPBVYZyihhfV7BQ4K
upg5BM5MapgeggnNT9I9awPUi8SgdvVcPdDnwO16rJZ/BcEejH2I166gQaMpqL0lNApyX/tVkFGC
EBJwunjBLyiacmkFNEzfjWFpTnftRcW2zn1dBuyOvwcfoj2l2uJtm3TER1BAg9SPeRid809oPy02
za8T49fJpbKdZxV0WJgFd5tnrxfgYGplLX3DKLyJctBPDlk0xwo0dlz5zUqHER3col9wNiOp72lD
pkwu5Gk/AGX7vTUWC0xOGtl206t/NJT2+y937uBxK+HHtgY357k4/PX1eQPCQxxDL8OtcCVpuZuG
2rpt7M0sciGSLqKYlgNzTGfTuMV3e9i8ZQhb3oM8KaUSdWA+2JnJJc8jMov3yCkBTYaoX5X8guR3
skY7q4i4EGyloBADAu5Gk9du192LCORMlUn+ZYmFf8p1K4A4MCAnX6OgUspxjDrH3IdUoIrpc6IR
3edkcJ+TJXD660IpLRGZsyMX5MvgGdgO5V8W/8fVRTeDLxH+YzDXzAzci0HdQCKerdnvZC8OA4mJ
yHXBIHhHMa8FZQpCN10Xl4cqeq1In7mo02nYMUm+fThk3wU/5bl//2UHpZTB9983xZDaR7t6LvUV
3jcnPcc62flBhDk+MJC17FDHiMbc1JsmzoQ6h2z1Oe2+EoUzwAWMFDfYwuHtI06wPn/5Yv24655K
51tLfyjXo1FhhjztrSORIC9M7chonOTXv98hG0c+pxSqPFASEGnqXlzdHp1DUXT8ZPFJCNiu6RR4
+j1HqlYWsqSzq1StziHFI6+T5vGoR5TwW1rtPgEHBE3VnkKRLVi1Ug/mrE0vbJ5OnKxu+dIgCsii
KczoXD53JHDy0IwvVSSokOOuUc4wU3/nWzI7SxhiSlavhWQEmnGx8WD5ZE271JwcsKs4dRlmJ1U2
w72wAeXBMVAmvo01mzTWciXPC4A4BxYIbiQEbv9LU+CnSNia55LkN3LQMKiI5wn7+c9IQWOLSHKc
IAHzjm18mB6CyW6fvyaxvcKE2Nx8zmzKbuj2BlIdkUL1wM92GLvTy9+MSPjJmw8sMuk/IUUI98Dl
0cTYcTemiwHiI0U63fpZBkqjcm/OuiEcgFWiPa3HpNQWQx9yOcKS2byYqjeEbiA9WdyZifXJikcO
yIRfzAEwG8QiGtzs1YJPBihCoKdhBE1474am16FVdJ5sb93DSCOpqoDhrEPudwUjyH9sFri9kzL8
PxsAHJYrQA4JcXSz+3yukCAAw9EJkFutf7LJHpx3faE3PATE3qQ/sjwL+WCcXon2ulahezdODdE5
EVMx3/njCKlLCwq/FQ/mkqvsPvBPkjcTpwpl6t+ssFdhCi1G1QHDPAnETIZfxIPW55JGCoVW1bdc
DpAPY1n6VPQe85k/aMZWWbOisFGmA6wFoDBZhubCSb5IIkEku+TqaHukTWsWv8fKYkA/3Akv3uT0
fswkVhyvDKT/ndDRhWc/NoA58ErXHG//TeHRRjuBHIW0iwympLMCEMgyONyx1VxvMy7guGOjQ0qx
GHUMrE6Np0aeRn3CXEkVr+KTaxAqAe4WKJYCEHpt4WNiWy8SUvWiK1ZX8s9inAsVdsJ62VJufKkj
KYRFqDpfpEKDHGWLx061NVzfoGliYluaHLpkwaOBpU5dVAceDZN8Na2ziORN10/BPCnU6Gu3ajNG
pbKfPqb/KrSTzmDEl7+RMITHOQO17SgKDE85gunqd6UnFUruHbbC6AzixVwSkKwi1v4SLbQ1dGRA
ENfBkzVGpOxchhJfEBFgIOuzgPrrr4eDjawll8h94Rn9NHoCUpTDLErQ4UndNfsW4s2u/Z/0tfpd
45NiOhODNtY2H3e7m7z/Rq7x2LYzmSulBVbG1Yy4s969LdUVfSWKkgg7MwYgz+j8MTENmU51VGFk
ryVQU4XOaZt7oV2VrQuUsXdFamJDRYJITqouRASW/x2Vi9XNVQFxL46KFscNhb11jkzOshV0B0QR
pVkqfyXLlUZp+Xhr+A7AcYcjSouSiXqbNqZyh5zM/FIjeH17g9CT2tiisibEuXXKCpoKiEqeRVE0
EOHv1QXQD2KDkOXcEc53Gdi8PK5XTuBP6a0n4v5A4kspkXsCUOkLzU6UMZJfR9bg7Jh9T2a/e1NJ
8ebMppKj44526yDA5JC7Ayie4xOXTpKTlniom4ha4xsoABoX1YCSQlt8eRzRb6c0KS+a8uRTxKd0
Q+3GbVibmdR0cBRll39mcH2C4MTJKdmjQeT8Q+rPJmXHaxqZNzUoFHr8n0uGK39X+FmFBTvn2+5n
0tMkWtFEYcZgzERrjDAltML38ryTjk5XMLlXDpTNbxJ0BFNfgV4+/0j7XBara22r2EqlTda9l+L2
Z7IWWbuYP4Yx13MpvO4+0G2hYYKFB3aLpx4PcjRA35QlcVXUIzebkg3rXrDfKDp9pVxCRWa1ifT6
bhVDBkMETYiiVFibeNl6XdJbn+w30ndnS+ubJIlsF1iXxqQebtK0JzFf5ysNnt2ZYlgT4dYo8dBY
2zmTC5GN6FHpchZ3Grx0YZcNhU+bnCbmOvb2nbutYXyQOwHggIct8C+6XA9EXJtI1uL31A43yfc4
BjLki6FP34U7iwFDytyPkGfyYc2qtikw4x+y2RJbBIkrb+tIX1Wv++3ITmkritbgUr1IFaJp6cmy
Rdirv2h2rR9JsY1YxbT0or+3UH+edx4LjIJ3rog8QNDeYypJW5JgvUWjE2/0U6GlwafnZZll/rzq
VtiOYjFuTCYqNNQHaTUBG/yv2w/NFN3j4yB4CNHa+sQBnhqzRwOLFi9yLKMLMjlkJemqTmXh22sm
eqZDyWctaZ3l3f7ZJgGcfhR/2rTnmtlsoqSIaZWNPjhosCr2b/tKzVBLlj8TzIhjjpQCkZVwk99P
OZlyazy0je9h/lgAokVQ5UWzmMOotvMrhtiMdUg7t+AkK6ZpnpG2VnBY5NXrvXvbIUHrIyoCXihZ
h+65HHdjESbzJnZ1SMtps1MglO9sI6cnhiGgX/fhE7Twwb9vgV/HROhOvYuZgCWsk9LzQqwLresb
wsiRTOE/wv7FHWLqCgyxJIxGsNQqOYYgMsDcbjIihi2Q9btLiB0qiEkxiPatgSTET3aLJ0V+/DQ5
n5ceBK1g8aCUfgCLalvaEIx0XOiZppxsWZteDxmp2x44hRywRFhI8hhnJK1QQ1Tz1F2R9aF8cO6J
HJDIM67Ysu2bsA0KzzcwVtuz7bKMWvSUyCcaa3ZwDgAQw34XV7WWp4rBfpv4wPUw0nfk0Up5kVj4
pTgsgZBsSxYZLO/66BZEuQvzt9PjUFoB5/CIeJoIADdfj35ji1wexjEAKALTub4cHH045E+tn7Mz
SPUTYK0EXSLJ0rhKTrMEY89gy5Y4OOgyvmyuQMeVBVWoS8YuaHgVK3f4H0P2TDsn2UVfX3j1XyKL
KI8RQMKkvwHGrkhHdR2+Hye225SXsyjcef+6/rdkry8xOVDTmarvVySa7AgxyFYkUqLyVdu4xW/u
MwRtd68vPLggEFB3GeSrYl5MkISn+epiRLHWF0+fXtWl7O6QPKFR5071tyYgU82uGvxKzhY1xlmf
7a24emP/8lGhmL+b/m64DaEYymuB4gSyN4OYNa8yR1IilhlIShK5pDrwuPLenaDtcznr/yFpn7xJ
U5lDHHvd1qlHJ7j5iBp/iw1zozBLD/Csauyir3bMy2aLDW+D+rxAkuGvi2/xs5BKta8x8jca3qYK
ENPZetBcYbQ5YzVFjbqIMZxmzJ+W5LnQyYE4lxX5cEnfsS/hBIoRu623fu+1Fz+RaXcamclGu2P+
t4sHfkcUbIGMhehpmRq2bWuzlxGpR8qLZgdwyDFS6C9d1OwuVm9V9bCa4NI+WrzeaElRiNcSTs64
KZFLjulWiDvCA+4azCz3oLiIpbc2SgF9YHaCmF3xBEJKxIauFZwGIk+6S6Ym1j659pcQ6vEa/9vs
tAGSMDpCIdPM86iAfUPRQSP0Fod6o6A7MRXB+fP+8Xg1AEz50yc56p5/aRbaSxLzUubHlEFY645F
TfPqn92LFHPCut76vLLZfdteLPRk1LTfhaqKggta4+EPfhDH1PXAHUQe+lDQau1uvtQhVEkVR3tx
OnVCHCZt8XZrXxexnA2mfucqn+VZccAJspUe9VszzGzuSNGeYXZhjKXtJqr1pGXw+zntupkU7HkH
fX33y0P0yVdCKfwpbr3OZceAPh3m66uO8oWD9g6v9agvhdBh3J0OWXSQrlsO9ItmSgoIf7VLiEv7
CPWMr+VdLUjVQlJEa6URPp1Hyvx9AUKeTrpHWA75WhjoHkQmapL4Rn/FJFaiOAt6qTdJcHoRFzX4
IvtTneqNx77HyOotB7twZdMl/UrPYM9ovOvEUBw1As24vwjAQAFsgs4PfRWRxhqORwNgRonXLMhu
7g3O3YX0Qp0dGM2xRlCyBZJMoo+FGCgdXOzSYN5JtiLBCIx5BMFw/ZR3cNshbHHOc+H/MyJjiL9O
DUa+PgvDatQunCPRT95ia/6pnB/LZbTTaXFeKnYY29JNOgYX8szNewoDH9ThJGEZtijigz1jcTmi
vRwjeyvIS82/CJDCM+edpStC4aBblfBwV1/uy6m/Io6a5T6VKG2AnthKpxyfx9+nG9yr7Jdjnlvy
47qX0I8f0QSi+6ZvQK3K/DPWvHNtHn2DPkyUQ7+QbP2vEH8CtQ/TvUf392LqLkrbo9NrYuOcQfEC
+n7PDLkJ2o8aTtjwYgD3KhSzn6WtQN3mrh47qRXXYi3EEo6zB7RuQVGrzMyR7+Wy8sdAqxLjnDNR
elJc0h5pwnspVB8iQEYBnQQq7BjaK6g15d6xrW63sha60M1AiwQZ6+5e5D27RzAY8rWswyMp+fyX
R+/GzQuv8n26kUtXYeHjfr+etPg2tqOy980fBuFHlBtYkgw5iejYXUlYKk7fIbRFVVcWvRVegVnQ
BahBddI+BnGBHDBD+Bl/8ZpoxGR1kfytlAs9fv4W01/qBlukWrLCiRRZtCMYJFnWZe/UoMQAOq+l
5J39lQsxGNrZqouqQR/cDhoFRDJ6uPixxqcC17lGq8y3hHW/HGMvRDdRm3VPGcM23W82DJL0nD+c
nqpT/Ehw/j0trosCcR5mR6D3QqumkauicW0nfQdi9v6444OD68khcRfa+Wg7qThsfkWZFJvyISDl
7b/IIoZyHZOIRYtD0JIJ64n2tjK+Few+4d/T8IsUzETr7MtoQu2AoRmn8+3Y58eBScQDlOV0bgvC
mO8la+7OK2NRuntN0SQBrAHKQK9JTFi45mR9PuSQ7BgcjEqdZ688Ekxbk3rJsLq7b6SQ7BDvYoO5
TGL2jMFEy5IinJRJP/sz8aEcZ4vWheue4RigFuPdmlEpONdbR6V0fodqD4BFaD0CWAjdwvlCG/VH
iQgrnTyQA2yV9lHtnG36poqZG/3bD0WDJ4BiWLVz03Z9SYJvKe2tBwBfDKD8FhgHGGORtLrmLo+S
NwTBh8LBV9TEX24lbe4Jq8gHBXjM/boJeSLjSGJ4O874sPeqidscVJThbIbMFkcWmb/Moj/X9JMB
RApMPu75NifSN6UNh0Bv1K+o1UkMob6aj18l/tTxDlYqniwJPyZCXGl9w8+2zF8m1SreoOX+q91n
loipMuDc/c6QtG5f9XylyI8GwLN6eP9Bl2mawvHp0WKrePrzers4DstbEfZP2wdeq19uQkPRz5hH
w4hTfLZnRt+pyA5mS7CgvXjOKxrQJing1myCsUfrH1dKpIS/n36xQ08lhIOYFIef08KHvEMjGxcV
Rkwr0LCRHKx42tAvPq0/umZzTp9U81G98wED0M9VkCjW5xNbD7aoJm5ceobItyUXFBwpb8ahXU9N
NlwgevGrRCp7zDMTJyP/4s9f6+EOEyZ5XpvqDqyEQ8nkTUm5rzhXwZI1/ZX8UOFzTCHJW76k+4Pw
o/j7SWvXmZI7Jv6XLyG7Ej/Um2ia7jeo0HuiuE3vl5LHFuMBoBXgfjncguW2Qk8UBMXA1+6Tn2S1
AtU/JupnrAGdfBVelnPuktcJyuDhp9IEfgJ4Q4EIbxDZYeLDBBxH2KeUmWjJcN30TbnQp6Dkm3Mh
yGqdmoAhYP/qs0MTDqBu2id5Lb8r6BpT4LOlg6w/FAer4wOFc52kGxVaX0SUuvIvRd4IzjjAIwLe
9vbyebTJ5sRYCw8+wpbcdXg2qB/vybwMdMsiEYuAnTq5HvYM+7QGB1GvogC0Bfc3cNjQIlz0ubE7
jDg2ox4I5byv7c1Bfgw9B8mSj0PaPoxVcUlkKIQvpTrwzBigPhtvCbCLaXFl9wkEzHzY45KuFSH4
GXAaT5LgcrUMzVP2t8qOn3sAv3tE5VeuhCFGDP+o0Hv4Oe8u8U21UljR7QvQDhB055RoFBnJV7cf
6tQMvKt2mI4D05BkldvqwYWCkCd4ebwuc+2oAvK87koGbhL3Bb1SfZOv653rsaz2cvi0pmCmqxIn
N9ojA7Gl4V6u3Hle3WqdP69NxFAEJMo+lm723kxrU8fPo6s7UIcAnVXn5M0q9UI90f+y94aASSuR
u5K4xdyZk7ebUz9kTf5Klx8SV5pnUKMnbvrAMtDl6daHuEeHRN3fy+D7ho/o1qLuCdU3jzrF3vVc
Z2Sm5ASohSxF5R2teke5nplBCrN/DucTXjtaQfWMshZaYmLlTkUCkJefF8aUfyF/16T0aYvgMtmG
oLa03jTa25GZhcf5t4J8rW/8BeD8duS7BW79vN23rPpc3yVp8ZKnbriXnCv58XX/dRALAfIUP/oR
xkzwsxGQgdaSrMLeWzKfFbzAZNdtSIVssfsRYYFh4Z22shFj9yPPMgsSA172bR9HuHLLb1kizwWs
XCDlKggwrXL02GMVyveBFsMCpULlfjqGMOHS+b5ISe1NqR+0OuH/RdcQmypAu+NVyuYWKETRIymX
8LuyoBwV9/rJZnyw9kzn2IuHOV4cQRP3qsZJ3ca8FDchOoKfCvjHzCrsBX79NJhDHa6gLGxN0WLb
HQ6GxzrsZcLUBW3xcIUVWGksIfEzo5jGfpx7msIwMIfvRTcXSZQCZvj9mGywj61c2HcKu8s9n063
zU9uHFYQKNvQMGJy4Gp0Uzrj7EW5zPfdCjiLju301avVNgQrRgbrSgeospSqXBjw6Y9oZD3Cr3EB
iq6ihrqzBKkx2cMmUcoQm0APEGXwu1Leo5hYu24PFFrDzhm6NBEamlZ8TMHgKHupuyD6EniMRI8w
LBh8DVR4kaCGYqTlE6M2QWyv3/OvxbbDn1rBU0w0nM19vnok3FS+lEXCnfk6mRaiVLJxJmBCS0TB
gwJxKwDudXvic3pCCZjugMA8wPD91nXNcNz9LYZ2mPJMTIY/N/CF1MKOcfVqcmApywjG7qhMcNqf
Hb420ECybb7EozdIky/BHPH+ZGMo20gfr9s+0/id/sffvaFsS5S+af/++d0OXCu7flSrN7mwQsOe
TgO3KQn6xnOLn/bBMx7XRFcsdTa3lqswWbmipU3YexFVErvK2xw14BoN+AMmDKA10i8rdeh5bgwF
RGbHirLaun4fDR3vyfEfPW69nAzBPYq5+NdTr6potj6ivXJfTFXmevwuxA3RG+Oi+21jl6YQOcIE
JNP3F583o7uMHxvH/l3TnyMgPKPxoC9aJ9mtSNAr61451cwYlMgD2MR4GYk219uEQ9sDOtbaB3am
5zeIC4IsfF86bTZucYoSMz/Q14w4UhW6pMwZSzUjHUM9pp47oo84Irn1ClvjBzOLAPwBaTUuyzCi
rghoKcgp3sCoQdOrEpmEErJe0EsBY8sTCBDsMhKoihD7HwOwALqkWuSJ/cGiLdMqtxjrNgCuPPx6
ubrZ8kszcgm5IioY6WiDX9nUwCpjO979mbhKefKKKU79xbu2hKlf5Y/mhqUffDDsJSt+JfPQVRAx
pJqZy6Ebl0G734wRx+fr9NThUcxnCD9SuWSARA1tUc5Suifk/mfuFDIHZ1HjZqAN7O3YKWC+aXiU
bOzcKplQpIaXTbgGILoeO4zPyTjeKXLZnbqLGEyyJ/Ck6dRBAZ00+IgKofibR333HjaWvV4Nzycj
2GNjPq2iqF5Lr1aVrh4iMHmUaJh0gE2bGY74F7Qt17e+gitw/xufjldeeUkK+gRaBdZI1moqVbwZ
SaSrg5bxKeda5r0bqdZ2JrOY98KMIlwP4zRxXEBTVaHQu46GdgkgviUDMkYrDikK/PCdJa+6yYsa
O1ecVguo7W86AB8aKhx2aEsn+q6PopE9ZaV7T/LqiSrk49TE9PkiP9HoLtzuSfWUGi4zSC8zkfZA
x4pRLRCWDvefI+O7ZByKQsqxlNmLg2JlbcWolJ5qNkDFVUw9g+x+7ZGe9CljeLO42QmxboyHNDLc
lXFPlQ7/QiOKuwHsZy/j/nNdYHO3LX540OCyTANR7Xg6LuFCtP4iCPcEm3CoxI27opZ7oYewXZfc
aYKD2o2+7ZQS+wB6oDJvIEJuPd1uHKel5W33cdcGPwPraJZLxRI6i40wkrBpcxidD+Pv9+X9ygxj
5HZvq5mIC2QURF3fYXH99waxqUY1PscutaiJvbgPwnksyotbj/oJYnHa6xI8h4kt/kVQvmMmsGz7
2BkR/mm4Ussxefdu2+eDQsBVv6sTEaFozn7zeKzugP/iB+drMg0tYhM2Yp2orR0vXe6Ldil2pNth
gEL2wxBDPtMLt/cjodRcPyXz7+oLoCDcCeels1WtBHiEAxtv5oYics5zYH81SALiUSFWEhJySkrE
FDUeOYfppv4zmmr03cBCBZDc2eSM0n8WNoUG4dbCNeeFplkAYQlAmmwmuTv7655UJ/zOB2fbeZtf
KN5MKkYm8qn8cYhEbO3eLs48y1RmapHReGJlPQ3iGJr22299jWkUBgN2oF13nvOOf7KCGZYM8cEh
n2t6jqJoSZ0QPCi9HgHnsFV/4xMKUVwELVSH0U/vKsYo3CJH60pwlfDbE8CRQveALeLhb20wDmRC
BoGUGedbVHSW52rECkUw6X8vXBwFfqGjEF568Eayj6pVYfZnVOwA3W2NVUSYxh0/KWqWvWAz30DV
WDKqRfyfwTcXba7SV58n2/Zv5eHVMlkAgcgSNCZok4D9xJYgOO921v3TcHEYXVY3W0T/LRd0Wvp+
DTK7s+oA9Sprhds/OvG2/rvVm5aL+wX2f4T3dKFwcZR5N29s1HUPcMFV+18Ausjqr3LnF30FoZWb
VRe1l4LrZsTvCISwsloQtnJ1tHn6wu6DIzw4Dr9ILynj0sHNt5Gx9FexfXUCe9kLVoD6IBxyCFxL
fHIGsbPdxxMPOl8NdKni+xoTFKYnMYGm83TjQTz82oSK6yJvNmeIGQvm23Uqn6Xdk6QPDbAfTBZP
9yel7iF/7hzof3rFxgkZ20JjsOj/9w3SNRx3V30XckDp862Dh/o4rRZ1W24V1TkuRqMs166gfYCM
u9MojYQyiRIZsqVll3ZMtdZF+FUW0blkJd++aZMP3uxK+69BLQeNHkk5rLeEmQ0nE394LWTF37dN
8FihkV8LZdVxQGCDoIzEvJ5hx0I8UhStQacTQUX59dgUVVirabQgt7vem3a5GYNqcSR1eOtr6NFv
t2rFy09nXKNDIGic3LEtSJZ/7lYlWLIqHmwkI09vTejp9glp0vnlh4Eaxv9fo/M9wZ7/gwVE9JS9
tGu55Src7a69fsHhgOzJcF73k9jYAlLjj65YjLRCMle1mH+CbuhSTXDkCSdIvhCfu1QtUuphBbjW
ByNpfrJj6via3+E24kkBxxi+71QuMAgsAZl/qMd8Abja2t23tOC8LGZSqZFPVHJfYoFijJEdzzdC
O3OWPBJWo0kOfGFWwkSVBm1l3SeNgBlOBxAZq+SxJSbR0gkDzxWSGFDK5uq0gQZtyePc947RoYbO
X7F8lvlyyC31T98C/ybLSfTgc6sp6ybOhpZIdGDeXa+q7XTUMTjO6Xjw861ZM4stenkIREUZ6Wur
RtL9/jPswROO1nmi6oSJfuJq5EBf6t2HiBUDoysSs5DeUZy7orWR4wHiner/lNLedoypoJvGs7UF
q3VJY9pPSIoYENgru5ycPdvIGRH9EvybZN12zG2zMH0jGxn/ph/gr2PDxmJNcBVkwG/GVXjY17Dz
p/+7Y7TT3w/ogSlLQqNRcTd6FgxqPWQy8LpIxn9dWNP4wkV2sZkr7br0SzfEX253BbH6G07OLI5P
TJ/8uPpASZFaTVDwQhA1UhcVk2N9nQGuw0dPSguwsIxFajJTTN9+Z2KaNr5b8QWPUM493bUNzvkl
cyWJ1V0Eoxsgd3QdX3l1mhBMR/v7TkUW7fegp7gUpb+T3SjxGM+O/5qVQA9Jv80DAnI5CzBO7crz
3WHzSjKqrNtwR1hQZETcOihus85jPk7cey3AWkGA0QG3vq0A85oelp50WHoOUe1Jy4or8GuzU7vc
VH1/ALaAfHHVVyviVLuV8ja7AxTYCqo+wUF/DAiiY0nOV1j1CvjoUzeGL6JD6kaH2L4LPXRQEpua
puZM5iVfJ6p8RX9+xL0sZpnJ/0hOugH+fzKYgN7PGMYWRVSRBXOKsFdzaJ0jEAfS973ycyzQSsSK
yZMq4jlT60hyPfKmeCyd2si1pXwqXyv2VcAEjn5CUB3PBfWBQefOYLu5/mlzRuQqH+yG5ju6KAEd
QInjMSmEQNM5UMPihRXkIKR9F1P3kgWIJ1CS32qDfrcvIZane0tZS73Y0whySHLdCQS6/vZA8I81
IjNlQkYi+21xnIogZebdMRWMZhGe/pK+T0FjYCm74wluyAxLenIWGlCeJNn0walPm+YHE8paatLc
VdgrDeVmv5BVarar2bo+kgXqZZbH6VEosmFIxaalRJVIujEU3feu2F1mEvfHwEeXBCf6tbfNOPtC
xU5nOZN9Zo1G4cIk4YCR7qSxmQxuPjWJnLu63F3Pnxqn0gIakbHwmF6AoiqUMW1LSO0kwic16Y3G
wJxbEZwmqbnSZUeArlbGeU64ioJ48ndcL4O48reaurQpyD57qj2g7P11qIfTP5ZH0uIU58Ff4Jcq
HqZABG7tu7NymUC8nrhhPvHKkYjf9NPzQW29BAkD3ItkTLlqYbYZejZm1/s5gr7z/Tc/YEQhore5
wbUjky+/Ula5YMUf50vWJba0pBhqHrin8Qinrdtp3iJLj7zTpjvGsvM+MOsRzULpbYyH3Xh87uty
oqZba0Cm0baIsOvcObGBpThFzqUJ8y7Bw6uoPy5HcpcQTz7YP4KiCx0WJMG8iyVahfQ9CsHUcU47
ihoCzoGD3/1vuzU+H6rItlVgxTXqRlE0PBa0XukbEwu2oV2sbQG/BROVScRCZ1ZeAUR9OFw2+TE7
svwnWpCuttwBCcvCcGQCiXZv7VJgLqgL5+TwO3DgMQ8MfpRDmpMdwnTbzWOgA2aVggZl0ssDWZpC
der+/UZj7HsuWlRUqw0vBY+C6/tIK2zQ1O0rKJmjtN89Ts7Mx1GNzI4H1UxjxOpG/meA4mJSs9uT
q2QRSuOpBAf2QaD+OcX7uhBt2zDGaEWr6ug1DByAzR/09YOXjnmHh61Et31lfJZje6mxqCau+Qoq
XR4g00kV454owZ2nMQz8ZI1Ri8bf9Wwy+Yg28I7AZWrvwDpFzdKlgGvxrSKvvoK2c4Tcj3diwPZb
8+ViAJHcPsLnDhNFzLpO1T9g4vsWfu84DRL0/yYD7SsIn2zjkMtPk//jMt31I8ghcXXerzUUP2mO
ypA1qWScqZ4LZuv71rc2rCj3S+rRKw8OdawDtoMdf+MjgeWtMDAwGOkaZfJIHq9FDqpJXLcwgHlX
y+JnN3fqns1Btrazz5785dL52qj/QqR+mOi0KeUFQgX77nLKMq4Xe+CGCUZWFI6nAz+wmWDQ2ZXI
pxlRWgeKE0ycnEpwGft3yeUUEbaAcRqTLqAqcimPmzg6x0gg80vIPJbVzJsPb4YLBhOdLs51qeAP
+Xp/srjIQiYUittjfe9OQtvQ+ybnaATf2MdikJpN6Jo/pwWM0AC1SZ//2jKpAT8OxpprXo3T9GmZ
+FgF5Sk4KsjL/QHZyhkj2bjqidegLJLdf8do5GeHljytVlsXEyDDvMHolFpcGNKSsWw5BWttNo5o
liY0O1rj4SIv84xWJb2lQ5oXo2VDiLxtH9GN1qSDLL1ycBwLn24NDXP9w0GtAABunNWIsBVQRL5y
UCd7p2T9la48XfJ3lIk9qlZ1FMbh3fAU+p3tE5vnZEOF1OoXUj4yTInUjpYbBw9iFjaS08HkyTJg
ZAiIX5Fkuzv2SkquOm19iVQWf3zEgnE+Ugx2oOqg0ccy+yB1QB/XqLEgjdFmFxAkklfWxiuU3gab
5rDceDPJDgIPyVy9Je+v8Oub7cxR/DZXtEjbF5Wnvdb/8QinK7QZ/1z0iB+gtAgbbGKPncPwISGs
PubYentx/h8sAjx4zlguSjDX2FOpqpA2DHH++3KdLGWO3eQzi9ZtmEbUZY6iC9IV+MZSqtJsihS6
7XLqxA/vE4hQgUGav1twcstsexQRWUaVx9U9oaYF+E56V67Fs7nxYg82oGQpGrCSeF1VM6qMjzxB
CtOkki3fhMMPUQS5r7/R1CTSsLGcaV6KKCj8yCRRlsP09QIAn8uSm7BEBQTwsH63YH4Xl32Aj4TX
Wlv4aL+rs68yIJXmiCnUkf1FxndvAsW1NmF28csqqfNj+WABjjv75x8wyPvHcPV3ke803ciyOATL
0i8nfeF66PY6GHRGPdAU1SmtVFLLnJ8+cDlUk0PS7qpKWK9i039Tz54y4lH51JuSbyAPGNRCgNkQ
ewBJDTklnhvlz6fiKHCYxKXbBSUnFZiYyldehoP0/AXchs0ZyZOhuDSHNoctdLiT4WU292CNUuD2
vEufwvTx0ZWgQ2BMmUPT7pN66lUpJ07gksWlhnlky7eJhaOn9R4A28AOLHqN2mgiOiW4q6HroYuH
eBIK63nBccD1mZX/y8unFD6pc4u8XKqFRuF2KzeshDKbH3YvsJ+onRNHYhVrMi5uPCox1zXWGJMu
E74Jb18Fkc33/V0kTyzZlD0GsC0OrXnV5U4G7P+PHHuXni1TxMmj7sm5qEX6P/vrqz29rJmHHIpy
tKVXFIKHialWqyPOTiBoGkj4/Q9MNt3IBxhZZ+0h4RKTO9kl8eQpUn196bGCMx4DuQ9MMXoE4t8N
0mMZUKg/mc9ft5+MuqZexA1ZbUVTyxSk2Bs+WSTlymJl9dUSkQ/1W4NfBmIVky9SOFe/+aBoRYpL
v3ZUEgmmO/Uq6AK+c9aYndXxWT5Gzr0z5GisUdaTxUJgv1J9uIyKBE2JMCKsPEAZZhgRexZ1G6/V
DMUAOs1/gLADwUzYkyHQReXAQ+Dc8ouRIBvbG3J5wszcBEo+wQpUSqoJ6p+Ffu/efYKEFsYuEVHD
i2bgRF0PYLZMiYQy4dlelv+fJMtKrffkx12+mLUZx5ysFM/VbnhcYMIS9noO64NxEpY1JNg7I6as
2e4TavYZcAg5kloVAz3qqZpjEDTJbF1sOM0cCYN7O3sxtHxhGhYACbj0uY9du90k34xV0mZrRgij
PHlinxrv0KRfGmpqUfy9fSl9shBf6bJWK9isPrLpN8OCxsaloxDGx92hWQ8CEXQUUD9L8nH95gpg
LpW8Utc8DwQvb25U0RnaCnNNFtvuDxVkl3/CdVtgOK0pRfGJP4EAxNOBVhTEHLDn+hPuBx0dxGEA
CMTFTFwcYIa6O2uh5Yt42hwJ5RYz0EpUsqEmpo9QECX8TrinazhDMk0huNxD+xuvxR0NzriehBie
0DtYFfrsYXA6elgL3uNL6x4jekOACD8mvRtCaC+iKR2ABMigHUKWehknnkemI/e/Fs14ITjpr/Oa
wvG+/TBnLsSBI7IdHjU7CMzocAsA1gIOUhn0GKxPDijoMcQxaBL6g+y/0UnQheJViSK/gkJ7LcdI
yP52Vll16Tc/9YHQH1O3ASkGCIEYdeaCxEayJr0gWSG2wRSXH24cKFXEWyl80cmdJyXIO8hh0aPI
dzNm3IwdMPkAapizCO9uDJmpdvAVxP/8A7HgGOBgyB7NHnE77UcchQkSuJnSnlOnB0MTA+K8rATA
RPb35Asugar/1Ck0rPlEBaJHz70QN38MgP6oBseIIoiPCUue5pm3em4HtDDduLv+DoGHZGZCuO5P
0wdB3FA+g0JNO9mDJz64JQM/LKNJGCpvnPeb+lLVURDnWXQpXsGW2xLu4hOVZzq1oLUpQB+0l0Gt
FTrUrNVUoTgsAcc551ZUYIJXTrKwpSz2nS33XqebPP3Aoxz357akgDQSk5qqG7unHbHLhV4/0ir2
tpEttiAD1bbaCaK8Hx/xpb4mZw+Qd2UkAUZzExBC283EWXl4NprEziLPcO/NERreg97hClPWa07j
oQFTi77rpYdpC8UhisawVs2WaIM40mdt6FNTT0mSQu9vJZ6C0UoDMO0O0E2QNvnKyAglPxUylZrs
OrwuycxjwAA7E9brZXyscsiy/18oHxwRaB9kvgtfdJQJOs7A2QJxXaYZ5r/LCWf9xupWoOB0HSdj
0LZ9TvHAUDV/ffUrD9JTe9YGr1pAEf2f/JOggb7mkVwmHIscyxh0jhVCitQH8mA2m1/9bi/DQbR8
ubcX00hkD6ydXkQKdNezJrcMiMHaKQ3vtcpNOWSxN7ekErPcrgtqJU8OMengG9waOk5f5nV/VTVC
w0EWnLG/BR+I6i1ExmDL9uXYca7BvEXB/oTJwkYUZFdDcz0nDU8rSW/r/lIxe+FXSWLNRdk4q3NO
bdD5aQn4nZtrqI3XvLY/jLNQf4Nt/vxceYHvvDogG0tAv1oMqy4jkHJznb0loab1MpITaES8U5V4
5Sypp5PtqP6EUi9x1mkHRQyAWCkYez3InNGhwcL/3nGDGM0m77ZJM6yZrQL3JQGXtJNkE2fRFvul
b1YLAwH3azodQ2eSXFudlwVsUjF5YFo5aHJdiDKwecCwP1m55knPsmo46QzYp6lNjeHmzElKFlhP
l0jaqxLzO+no2y+saa76SXNFHSPo0vd3/bg9wBFQEdXG+Y6ZMYJdWU/t2YdKXqtmFJuigfjxB/Ds
KoCWUUGSpZjDwtJNmezBDVOiIcTsDCAlvugdQbpp+rXpkUUO++jEavVcNaErZ5A7hBU5nIqXPw/7
2t2HJMETYjzAhgTogf7NS5lrYbq+TfqRQrIGBLvYMktk0f6u4yGUmXl0mQRkypxQ+1WSEvZNYYDk
gqYn6UU1AUp64UB9zfylx1kanqENi9zEiO9CCxakDp1Sq2YMRBvFZTHjnvMKsmyLkx/x34Jy3UMv
9CXQueXBazRs7xQBmN3D+g0Td78QHd+p/IFWuRrK8w8WgfM8MHzOb8anTgyBfQ2OpQ9pPeSuPYwm
lxSikeni6Oac7spgq3vWa06Atf3mZRU5Gbay3rULE+GWL7GfN6Dd4z31g3kQcJuZNKAJjtN39pQa
0I/KkgQf9dkPpsiyt45IXimeN9Us5nczStsRDBHYe1L5EGJDbDHrQ6eSWuef6GIHQkA0XLZIz3NK
PBtWg/mJTJvEHqa2MHFoWz6XP+wYCNs7LeJE0Cf6Sjt1MNDPlDLKWOV9k3OVeq+8wWQCYpZBFi58
IbB35FECTW6BJj/tyyftc31LSdxboCb3K1GxyjvtL2Yc0S6PMM4iPfGneQNmfsn/p3qxy05F7qxL
Eih/SNkZrwYMKqPTZWVR+3rlDqfqSUGK06nJ4ttsTRF7ceVkJ81NOlFLFccdilJhqyIW9UYRvDIn
0S/0AeZUwxELIJ+iW1N1mtrgpXzoCVWpUQA0DWcVbTPY20Kvds6tkbwbdJ3wA4nQrmQVDd1Y407/
ctmB+95TpyVNbI4yqqMdPu/IjrFAvoHNhTRch3WiIrdd7dJRuLEs4AD+rh0qnKiNQSIZyVgVSN/X
kSJj7XrqnWHmhbRnHczOn9ZBc7YtQYI6WXkaJO+E2e4X/VvZe284ZpXyERjIC3t2AmEN17Xte2TE
lbJQ4sCiRYYK0XFV4rRDn1ExIZ6tzzhBbrULVI6jkd84qgCBijTqSkDJPm3Y3ZANuR15iVOPkOX2
0fznHtNQQGIjKjr1C9taeytpOn2TYJxfrwlBPVlXGBIVOA+EN7jHSHlQPVHIMLJsWrR0q/vasSz3
J+zUaAWdnM9reb0wPRWud1jPmAJ4tUTHgHU4s4+mUf5BhopjtsaNIIIU30sFT1X/gg6Xa4o2WYD8
qzRIe1hCkYqT4+sLYQcA5XbKgk8pPvEL9lJlcDJE1v4jmd3ixOfUuIczUNoN+aVT547L3ey4Xfmd
WrnfqL1wGJKE+Iar3YHQIVzIfLL/sJY8WlkoW2w7OSeupC2SjfUedVPIu3JE5GUvZWs7sp/ecJGi
eQFHs274J8mMgPgGAwW+M23elL4QiYjsAHGoJvCTi+dqVfBGLapzylGscf+8ZEXYBktrO9ga4JVq
a+1NUd8TssGj7uNhi13FRhlgtQYO5oGQ+K85o/7anFYzRlGcUNWKhrpBLjpapduob2LxlOhyQr1r
o42klZvzk5DueOhPiV2wsqyEus2vXVIKTLJImfHrYFKajKq9sClKZzfcn374MycGVXO5sf2FYJzz
gj8yL3HsQUdGItpMM7U7JRiLXG3OpCZtwItfXQv48QBZXztfQB42xKSCWyigrMAE+L6X2R2sO4cp
ivATZN6Kczr25xY7g6BF1jWxqGvWUhJz5o/sDzjIYdmq3QknhsBFeaHLp7Bv2TY4T2gX/Qxr9Abt
niClyaR9hOv+S8uKLwyF6LxiCnWov0N/+JNrpmvR/SR8QJAMExpTfOLirFoTpz3v13iqcYUCASYP
4mMiofAysC044JZdn5CZumaMQkB8lHwb5wEYd/rg/SFVHmJR8k6FnhO6haTK3i1M4IfpcuhJCZh0
zax777sjw6UjxSehitAB3ttyUstQvJWj6riqUMU8Fcwnodiqdf270bBRSQTQWV+goaEsoT+INxiY
q2FyMppqsqAbh6TMP4UJCsue5GAAAiojOoaGAwn9fAWctipcJQqaZ91oE6LCiMGP01xTFot3UcnX
WfQZR4Aj+gWKXHSAUpq5LX7COJGSekHaQHPNYb9QRrqJ/+OKNC9vd6QnGmgjt8SszUYoRBXAd5Uq
y6egxsebRn7uD/SnoihXEU1rjIpmFT+EzV5OWeRySyqnTEkM0Afz4bxcz1LwWwLxTFDxb9+0AJWN
N3iuU7gymmZaclB1BR/zb/xTBywsqiZxtMbSa/9Npg1EmKXPOo8E9B7bcL199zviyLxkSPgbdv1J
cW4p/D8FoFoiLWlpMf5wuNpbe38OW5XIiObz0GldFS9g78Z+QVMYRFHhprD+earwoGAskFeyTCmW
7+qgZvpeeanYtFAQGaYCBMnGdvenY4Fi/sPbvvLP51NAYc/YdH6E8Escl+JxPPxaGzDZoQwjHKdZ
WF32AQT4UWFe621px7SPkUlAo5CzsHCbEOaS1uSzSIoSszG6CwsxuShcvO0SPg/FuPXnV6O6Lr1m
lIqc/Po3Rxr5mOy1qJbn523cAHoNKbSuacMUousN7DZa2TUrh0v+KHvGpwtydEB5Tc3C2/FXyRiQ
X7cBr1H6UunibbZk4s4kPzrOc1KJmzaO6EmOUzrHP3Pm7mEh5tjUYHs1jsUd+DqQaj+NunWrT6Yt
ALh5vrDogZGT8eILI8iNgr+wparCC4Z6jm6m/RWeVo2UM9zQc6vSGEWJb6i49v0ptZE6YoIWzTzW
n+2/LTMBH6CpiYdroyZUrj1uUfsMkW7PUbFU82m6N3njadF+Kp7FQ5Kq/xXnsHdE1csQslqCJ8F9
aMPqjjk72x8S1OLWKFnwSNmU018PjmPh9xA+O1/854WWexjbuqQPzkpVQ6dxKt4nbyxdUfYo/E5y
moAgPgWsvU91VyPKjVdB6ufTDyTYLT5yzzy3SvHm2frnj4uO5Gs5rR3wQlNW1DUBsdezZhDY0eAR
whvkdfVlQU8ZmxyVSSlP65yMNvaDUPY1OmG51aOjlANBY11jevsahkZWEpBQQyoitXMYic2gpsDZ
pwsUIEV38jUdyCujOyox6SL4VjPnsshuXUqtAQEAS16PBqzbkunzuy/BFzIMuKTl9+gzsAW9RSIY
P3jtJ1UjRsQ1Xf/WXfoauAqrDfDw4hqJAZ3bX1GPMiwoEfnCb41IyKHMWy/HPZsLy05YbslnCWOi
t0sMk+CUWZWN5bPcbLRhzQM8jow5Xnqk629LZESGvI1Vzv6+Gz6kN+DoSWQAXHSfXffMMHmHOO+6
bXqZ/PBx4X8uS0p0ujUPqMuew1Cwn63KwC7/xjRbDiyU4vZvKt7rGhrGHaJ7XbbVoiUZVuMJabuC
puoEJg1Oy+Mm4r9KeDFjbqAuPDf0PKjf3y1HjRotgVjBtDJGngHbUNiSQHFrQNWi4surr0QXaa8V
Vu5lCaBHSf0j6GXmVbmcHE3KOCQgCfa2R/uOm+//POEfcUm0rHNYLyVPn8zJclHXg13i3OSOWgvw
o1XI6Z8RdbFPcIqSmAGjVlYwh+gV29EP89wLSIi/GYiSTzrNbXeTJEKbk/J9sXOjbaYTSBxCGkzB
fHFGycujuxFD/UrUcw2LsLKvEKYV/It6lClMs7zMYwWcaXZXvw+G3ITuyizYHfEd5mw+JyRcJ4IX
xI9oN93NbxAuqOYw+p0GYxy4nuSo1lTW3YuvxTApbQF5EgWKO0pdGUpTfsSJ5eJML9jZXi/TfHbZ
NpFSFH48Gv3a6DVIfvcRdAtEJLsMys4lJ6WfyM0QsxR6xORGg/UlHpFRrA503WUYJMBlV7aNQLmv
cH0e3Ws1AmuNNp/J7PffYJ5EDAmCWCOQD6NQrg3yWoA1YmLKW6FkDmbgks8/Es/O73DYRdnpgLvc
0O6+5DRALLbMfgt4jFygnuvHYkr0uT9mdSbvWFqoGL+Q9HJ40uJbh0cOGTMpVy9Muik38BHKv0kJ
Oph2PyaOrFg9MY1M6RJBrV6Yc84gXDuufsp7SIX2PQ8tgvnNsokaxQpTjC7cAX9ZcFMf/iuecj/2
TqUiJuCECMNU8q3sKYCZcgZFOrLV/Uop1rctJEWfq4pJvY7i3yvzUemxWEF09PkvuVVlXE9wfLne
IgcLLt4SVJpjZq70vN29w7Xx6ghhEO60/1NlZzHASEN4EStXCHmEuzSLZl3GiIYmNywQ50KYAgE+
5toGzzPFhtb0cO7WMWDvP3V2hK2nkLUNANszCHdMQtwUeiVdfMseKhZwBwsInGTih7PKy7YBZVg5
vpaHi2bKzbppZF2TdC2rl6jus3XkKjBOXOpvkDVupWVjHQ/VbHDspF/FX0kdkd/NNKTl32iNV6eD
aVpKavHZhf2gvP3xkuT9khl+GHGGSTpbV2WNo1JgCLkRKiVvM4kgCGMdHVmBPkPyjWIVSj7h4IUa
4WlZwm8qkPbP2v7pnO14S3S2G4NQnTzZXSzcKEbz4glIXfKgN5Y+nYUhFqXtCdJQRApX3PQLQYMo
BHNys8VaJeTgJFz1ot1M0uLHXrEUwjjDsAuzG51svJwTJwqyZ/0aGl1X3HMpfTxyxytRnvF5TiLH
aMYt4G7kHywU7bYdowxEGrB3bOrmn/f6ERAuBUsddzS31uSrEt4OZ61vnW87BsFp07HK+1Fr9mOF
It9mzqiJACekA592V8sL/i+JUMpQCrOv1cuHGsS/QJzgyd4mI+b8KpGBUTvjiQvCKvULxg1R9lTw
HeFauEN60vMd+gEMPnJ7JQW1+fe2ySSmrvMIzLW+M6CUe/7B9uHE5lQkQEtTtceibAv4EIyy1hT2
rDI36w3MbUepEE5Qixsd8PPxFOfKhXUDE6T12HnoW+IErhjcI4FoZ7JbE6dauy8alFF4czd4ZAJB
l3W8OdgOfWDRF8/qNFhN0u9Qb8x8xYbqi1PsCzu32Mvzofkazu8BnHDPyVVoLXRfwl2A32zpHzUV
pqruiaf4osPNN79iPaW40kufc382cnqnK46tlb4GsB/Mrd5s8iK34+JYDS1thh/yCtp76t4bNJx1
1w8BxGAGv4iOsHPohdl9zBryK4SJJMQyuNpcz+jcQY2dBLIrJowHg3u5+Fjqt93YyEMBMnaNLndj
VhqinXK9twJQhn4gcKTUY/FfzV0gMiXiUU+bbAITCzybNyE1pIUpiA1nzwO4t+CcO93i9ocXWco+
eG681n4L6bevVabyJYkPbwykafijq0GmbUjmi9e9xnT5omxPOx6ZjOQydobTcTd42yXzbNMNrUdR
oRsEm/fFCCqAZ22sJPkJW1sJBJI4jfcEJx6g6Iz8KbbWTE2zKvo6edyK8G0t9xZwiEApcHKF7mkQ
/WH0H89FkkBLuYg/cbiiKnAGc4aI+cynnObmwRvuPe0MnzajrW6tfi9Uu3CBsRqB9B0W6GPDGnNF
cjxYBKdYK3gxIM2TuIQ0I5S4hWFwWX4Yrti8OBtWen1QUG8rK+nobCRq3MlVl0hLti+LnckaTlLP
I/4lZ8VoL/fquu9oPRFCoz5/GkxYJ6T3t6vnRcTMUdcZpYQk3gqVmpXWnXmJnIH/qSXqMTn03wCM
Yfxfwxo2YS35i/GPIeKLb9FIdnZDjbQKxu6HeDoKznBH+16s0e16DKxax8NLCyT3FjsVcPNUMhqu
jy2P2KcqaHD7C/taI6zfTJ4fDqOdwieme1aCBujP8CYx8WoqZ+HmdwP724I4GicW3GWBRK5jERyp
GIBx27de3IHhjqDSu1c1JZJBKIau9ktuZlhjcCBsk6z0OMtcGiLlt6eaZCx7b7oCh/ikYxRg5rE0
zlX1SPGw9xmhUO85gCHWzrUfJNPrAbQHxA6Q0g8XmLOaVhuQWWYLQZNQ73m/VQX9EJicfJwXAU5k
MFDTqdGlEpr0tttKpi48zKMPtFmvAVL0Azw8ekUMbWOH5mCfvP5TitzGi0ar81SBXGB2PpcA6z8g
FIQ9CxsimKnTjDGujj+OvSNq7qelMiH2rfqL6OYEN5R/cXIPSLYqgueQYeC2eBFAF33YEulXop8O
YawsAaK95wkND7LacsBF6QHHqSYVljku0u4wrCHHu4yDMMB3aSKBI2HZPOTlOug8vYydrKanWcx8
yKL4KPZimL2vvCsYNEpocoqD34wKrL8RoKHE42JFFtR/TbKbz1PONPiqkhZXbiaWCTBHa9i7zoHY
xtSW6rJu+cr5nmFDxt/pjLdKo56LKbF1hxsA0TW4BX90Jgk2rsvCVKIFjwXRj7kKsYz575p7to35
nbsGCnQumUVW3Me6K0kYokkvUV2OJyxhqCajkWqzrwvwUSQA9pybPe9iq9OxRfqSqa35OKfTMCEx
nazfbatg2siUFh0UVPL7m/8OOgKN3w6FGQ08BhYAizJ0La9VXyxSndK3ETxUgY2Wvg5I/7TmHh7Y
dFxmsZuKZtPasjNbY32OYTQuyJjMWG5CrOyglsSLg/z6R3CP0FkksAdeDAxbMEnnQ7lZl8Hv1Kow
dLeU2/86Fz1xA86jsXVOgn6ZaM3HwdAmCx4a3J3lzuamgL0GGVjQlMDCROq8QOYBifBd0/Cb/uyH
SUsvVg7cQrWKzt5Cv6qw1MArZCNvxkks9gXrNdyjD/mCuBCLzSbi8pO9otTKHBLqvhfFrs3A3LLk
rxXD3SFmKX3ZudfdJmckStHfILI613DjUThu2ikxkf0vHrVzzCDfQ7yAFm0ak9EgXGgpM3/YYnpk
XSJeMnVmZ2IjQrdYV/cc110/fh2spVcTCrkwJJ78N0y91ESgPI5s1W6Ry9QXeZeU7QLHimznmEHv
2HEpvZdEzrAOa5BM/7YTKUciO3dr6XiyWQoHNonFH3a8O9YaDItSBKVqBJOp4MI7DcgNxyIl4zvR
173LXvxfxM/CNWMUlWkZVDTj3JQgofs/I+njF+K34hW9le+lpzKXj76cbSW/RByXbcaXwwroCDhM
YQE4/aY04gaodOw9Mnau6qVJfR+4Xdqdzw6WnI7JNFhiqYo/AHUH1ftAlBQPB9P9/+okLHbRg5AH
vjtoDTlYqFAkeAt4+eieRl60k1hRWmR3Ku2bi7lYsNDL5Pa7qLJq8VCp2fH3evlKp6CvoDjjTEbT
Pmc8mjww2eB0dOPJBTUfIRDtJuCs7N2gGwqGlekX8eX7fvpLjqz3oQAU/LdT9lY64CoVy/WKFz0s
bvwD4zdtwgUqmjp9RfYnDT2EjxjxsyLfToy+AaLWaN3K6ocMZuKE60NrkcPepME1SQwHTl3dNgZG
BedzQfEThbEKOtwvSkGrwd7EG62M+wQwhqPRjX+GhEhCWCPRiovR7NJ5b1U7UAXl8WUj5goGSsat
LHchKvE4xQwzGygYISZVtKrSd9zLyNo+sr2PZMFa7EHmhGsCmY47XUZxVqY4v4Vpq4REZnZzVyje
ZO3PyOBGHP5SCFMBA8ZWoWBHKX2M6ZWL5eYXhuD6hdOhWYIcSF6/cHXTablyhf6QEaHT052oYGS3
nqgGQ5nE335nTVGQKme2l132KVqPdW35E4JuMBGFPlJDn2UMS2LrpbfNW20LIdSygm+d2U2DfCNg
DazoEuNoFGxSJW6B9XJHh+zDK2TKK/sMDssG8ePqsnevAbgI7CKuL0tHiUCqOW2MKm6+FFtNPP50
nW7VG1CAG6heiIh6LSs/Z+aMnhl455549Ao/PdN9UE095dfVNk12xlP4rnGuWitlrQrQ1oXW5+nc
7+Tw6OpActEmMKU5fMD1ihNx6mq4UwSa+3rEsiA2CH/J+SO7EW9cubaOzQhlksNHGhmlkCMXiihB
+5cFmkEZ5BPn/63/PCJAkNXauO6fSf8z76/Pv2mm2qtea5EgXvS59Cl6UMl1fvFb6mQfFi6D6xeY
bNvSZqJjSujEGHiAEj/aNP4Ssg7lv3ywDqdKgv4IE9GboGtGqThVItYscofLvEEYSvHNGwW96/CE
108wj6QUkDKHl5/R1J98jDpoDLZCNOxg//t7isMqbbA3eTfCKHc/dSDvNbLGpt6LW37Hq4arORy6
/CsijSA39p5+PfZ8rUu5cnKdVapU0nhDqLhzIo7cCBYpk7/LWCs8ngwLK5BJpaSZD0G5hmBTJuGo
RLgGgPjA4Rn9S6PQknuCx4kwlU5UCTO27aGWHu1mI6RGcR1DmQdgknXPmif1MpgWRtvgtHYzysEp
tSa2e4QmBjRzCI/+0tJ/G5SOxY10y3oTeBFoQCcuf55h7Bsw7whTJkpdvlxFNP63mqgIjuXAdM1a
9PwUtfDvNnR2ZR4wlADgJ/ZsiASdQ7OJ58MNcKnQlIw4qZn8o34ZUu1RCUhIWj0TYvhCpLtHCsNx
G6B+s7kA4tGOM++4CObrpYuXrb+uq2+apndRptJGiDlJJSw9vkmZh1ZZSu7Dj3kMmr9aIJU4l5X7
D7E5wBWO86gtQbDpsOqNmRad0B+CC8XA70KO7oE/XNmCxbFJ/nlIKOvpi+ewH2QB9NnSeK8Bz2BP
yPl0yBmEYdeyHECh0pESYlW5GrKEvG59DZOu2bbKVBUUUGbujHvO206vOcXqk/ajS/3ZFGT38JP/
ztwegHHKKCzUY0lJyj/GjC4Z/y6C8+ed5VohtOYSNF9epPqhba99rj/ubvWx5zHJs/tfcHSCbTAe
+YeXIxkxXLcptGCWItqhetl97l7qtwzxLIT2sR9yAkWMfah7vTYZUQ/EdrPHRNdU2721nPKsC2ji
Vg2xMCRjcBTuLMi6VskP+xGmPDDOZTNXL/dX1N33DEFQ3bwmI1QpZmewTO/spmI0IhLYnzyLsNN/
bi9Zlhpe6dc15UZ0ld6jiFFIZX3qeNFVpsxnsHMBAhZY3YusAM/OjHECCM0ndJmHLirEUc5KvF1z
wYYUFwoc4gptBCFVfaDMdWDz1WSYmY9dWNcs7Uisjao2yo4ltsNemT3iOnXlLHeEwbX+BdtXNM45
eFxgKAdJid+MqXogpBvklGMysJNs9EISgz2Lml867C0nVqZVvWl00kZwuThty9abljLPNBsiClAY
9cQrSZ0w+JAr4aFOdKWjU+TwFQ57CD791Eee6bzNEutww6dgKhLHNQmHpP3KDEBi3ecf4rZP1yn2
q8EFNcMReXkMm2UVA4323s8v1vFXn6iTGOQ0D1bkpsgM4cgXwZeHoZgG1LF1gCiO+UXWgwb8Yc+O
PbrrrdhVUp+UocC1sSsOE9mXMAIlBMWKbwf5oTTsIO/kjKYotobZKhFlDdZhwCFl/w1oVo4jzCki
zDIlxxegtICGgZ1cpPRc7Gv6df4qUYgmtZro1Pld7PuHuuBX5N9rV2GdYE3CfplV5YcgdbcLZNeH
lZVysSTfc5J/vRCtwtJ0lMmd4H32DWNk+ioTGbvTYFxeQMRAK5oCrRxZgTXPnqWTcWSgQhcP+UZ6
AmYOuZawQ7VUi/Nzt/H2LzBvQdcIJNyR88/gTuff6jLK6vUvSW6Klt1oCDBJkg7i20J+yUuUjzPa
jCHdbxusORzX5hFUBsEFpK/II8OJ+XIfhgvDCzhmAeXYyT6G1P+9DEZMKtAosQUToiubzuNmMOYr
tCStbySgou/BC/giro0L0Lz+lYaXyl21zjYtx9/SI4O3YQTl0gnmK0QekylqSMnne7yic1s8HOJa
dK8aanpO7v0piIdwQY6uANiwwdnmKPfJIt+oKFts2tJX4meAD/7aD9ed/ax9c69roCMMCbZoT259
VRXSQkoNWfvJqJFhryrLJAOblnRv+6q7E22o5miVBhaB8Bb0MNmIV2QiED2zJQGcLPWBdWQ8Hkus
T2/MH5udDje3d08qAA3d6THLex9zXp7v9LkC0mF4xRUzowrxajoim8AGel3AZLkaVfwJZr4Yi2Cr
+xT4FXNh44e+3xQi2Nx6XWuNq0tohsInBzkE2FGfGxSML+nyVwdIuJXwVThycIfvnUTLgOX/ro2m
it+bVtc8aIE6bhNhmE/PO8I1TrhMaGKqlsQH5/p7w/IE1wqMjw4n3i7c+hO9/VXfKc4VxrY1sQEy
1UX8MzZ7sK/2zD1x6eqA9Cosn+vEljjT9kqDuCD2c8HzovSqHOYTXRquD2ddMDf0Fsds3z5EkllL
0hbbfFST7gl0oWz/9MfFD0/yJRxFQqBS9Ub6kQ74d35Nk11t9hNbZkHSL9ag4rVTf8t+aZGx3W6Q
4J/GZN/Zkz1rd7CdC40wDy1IfHK2d0Qi5F5cxtvEtHHVrCZoOoLEnZPeMVYxvX5wdXJnjUzm6p9Z
gtbNwli5vkSf0cCKkn5RdHDAe5vgc71m1UZdWXslF3VnO+SsdJ8SsN70yd2CfURpSvlLs26n24kH
2+9RRwX76Opoc7Zd80Zm8zI9hO/TH7K4UYCkn51LWH6jdA6WgVT6D6CIAqZzbQn8sMk6Lt0sA+hV
cgsiFsTYmY4ilCYxlSUpGRyk11oAE3uSbaL5iLxK4GSUT9gJYLV80qkQNO0ZTL8vJny45oiuldtg
EjdCXJB1y+9bDF4K11tlM7j90wad7a2yLHqQzr1TjEcFII/VaibC0obF6OMUkMOnqpFgnn2XF30V
8oEcGnzKOGFx9qtvEn2VH8pKXxLwmrA+/rh9Zw9dPZAhri2LIoiL3FtFRIy9vCunZvy7klNUIvc2
0DwoiheTQLe8acIDWv1gMhDzT36u0xosQdvvrU45gM/pKd+Jq9p6+AoAWrsrCW4txg6tRXLd9YA9
S1tDagU9ccUG/X7ZfnXsJs5a0YAgUVFHPgWFkxqwRJghhNieCSCPm3yLhToJRCh8ZRszVRqUzqES
UcgfPNBSbL30UPBoIusexcfNzhduPoMzJrRsA0EU187j4rErZ2hb1crhW00xv31MYMMBaPZZgNnI
z/T1/knAsaJYAqDF0adYRpNIslJXhA6iKPidXYeNl3IG1NfsX6kwpLLnOT9sOtPLDSNg0ADZYU+o
QlrxNEq1rv7zY9Lmwz+dO2Ql3qN/XySpqNmdsYEx3jmygY0yUDeqA0ay7E/Ta+IQH2h7IXzYkQc+
E5nIhfRZg9e4FmkoBgBy7UYgcqm55MHksp/JGnas55TP7l1lZA+JUdcPbRnVvM4UyfJB+DsfHXm9
cHc3YMEO1YeOR7d3ygadX2Gd4wncKQ0NbehYs06oUaHIQiwnnxtfACPgUy/mH6A+UkEfK/uljb/C
4VesIiuqy9eHscgb6TQ7C1D8K3j/XVsrDYKMOzxS4O5ztwipWn4YtVcNq2EnhKLx+cFAVTLx7aLd
i5xzhJyc5wAQODFvth5qNSo4rDHp7wXrNS3/fNPKdkh3W2cr7hcvzJalZQcorFw2KwM0D6MA1jyN
SiCxGrcoKCYmpAjzA6v13duq71yDkBLZGHRhbJ87r1XVyyX9BgNtJGROrXBUQxXJ3MixXl0o9+DH
xeQsMqA4nskmmWrV2y9i7LuGZzThEsuzELoIxfn8cBGyGiqWEFdxVNTKDhVl2R+i0q7aqnnmqpPe
ixCvyjPKVtpDg8uxCU0dskEygD9pyPtbBwJu3blhtBP4zHJFbHtNmlkGyyy4LHYjOt11mDBJVLGf
6v7e/VPqvBfXjQddXOXw091SDJc5IHfXjfpHkHDatYvjxgptNDEh+c9pF/sbAnVUhaEifQJATtk+
qVArE39cLSA3ZSU0WEgZjgsAoy9mPjq99S+CKdZETIBHki9pEDsRujROgiF2zHo3DqqRq3HQNiRv
fGT0ydsSP4jcAC7wOW0Z78Y5sRPYrzPH9tynG7qwye5JOBQ/vE+r52XnezO5ZoVn1GRgYzcbMfX6
D21ORdjZ/PYoSQ1gXHUYsVTDFR7zbY0UgtbWQx1XTnqmUcUHawDAqnuc4DcT03fAnh5cijxKI1DP
y/OL2QpY9HKvpR8aGJ0hXoz29s34LTk/ykd6E2fJEY7Pysg9Q9D1QD8M4ROSAZE/BVQWlYrGYD2t
2wplc43tYIJKa/lLitVwITLCtX/48lTPSMojSX9Q2vneJKJ5uEjsULj5vXf/c3EHnvYRLRBfcAq8
a/LAMG7qeoUTZ+oWKc3OCWJMuzuBjvNMeFHi5mVXAXKdYEIkVLcuoOZlfIzTnXPzozgHcvlkFy/h
y6Ij9BVBulCQbI0uMn3dRZanwsjOTWYMDKWyM3fMbfm8DI+MPEGXavrUWfskQLrwh2JIZlZ637Lt
pL/csYBn3kuQ9pamssShtzIzBw7My/QxbXpyjZW0Fe1R8ObaukY4GomEhsUxQJf5+HpYefhpJpd3
mGEG/k1LfppVUXRO4MRFb1k+YxPcJxXFhEj0vrJnjy/cD7dtBSxNPM3mtK1G19QzEdZtziEdR26u
l2+U71pAmu6oecYCYArOMbdIck8b5qcXDE+No/+KzB48wqQ9njfNVPexOIG3AuyTfMTbHV4o1iFT
u7VLT4y0d9giXC+YEEmQmYYNfVBJvoLMRVluyF8S6uwluWA3otKf1x2uR3ktOUS6H5dRBBD0kXPT
6sluH4HqY1PTNrfskKZ0aLec/VE7M+is5DvP5eYBJD4UN+BfLMAa3aufrNcRnZFj/TR92yMSBLNl
JqaRuxw9PGEDEaerPI2hesGVEhi3lujcI0ayN+bjN9Zz0vWZqzjOVttphWQUZgRjVFi6zmHwfl66
faKQ2lSPunelejxYWpX3QtFqcp3TwLGZlEomrUTVa4drSc5NLhku5CMVo8/Yx+mjfZpCG4orYK6T
kRONoY24mFjENvEbvJV+6qOxo8OnWFSPB0RVFoH+4ELc4QEjeTYF81TyPwK2n3ZNuwgUWJ1ZHb/d
a5muFXzzXEZ+Ib1P/w7WSIKQUPJGM5pNX6fhh+0gjcYL/ILcFJm2pt3bFpLfvS+rSDpU0WZojBc7
JMOCvRbSmIu5mDHFpl9kAB+RSXXXIwQaSajjRSTB3ef2y272WK6On49LkU2qu8oOvrdxIBm4PBcE
AEUerqawrX4gdwtUKu0LuMXRtDJfkm/zMsjCMfu/0CXa4bx4HQmhgaBD2g1NgtuJVgNVJgew0Lhu
XAbxJKokwHukxa5m8q7zXO4jHqYpMjkIqnow1Bx7wrN4M+IoyA6G0t4mX5PeXy2NV6FG5MfSFOgg
f+HItpeQ43ffgePmXF6JUGlnTgBPo8GwxVT6cD6Z6Bm3gQkTz9l7b4+MdFlvUxn01Nnpqb6QQJ6g
njWQlPkFqoAZ3OyeLhVHHOK7U6+05jdSNvidTGOI9b3T4g/D/6VRnKBjC9bn2MFT9Zpqb+KlMUFg
8JfqdxWIippYZsYHkw7V5JgE4xqSDR0FNiiBb94j8uGdOKT3kGQ3jkyes5yAL4vchEXIoJwHQGJP
vPcef9Abs8tP7DRySMIo8ZmyhqLLfg9+B6O2RM2lKBW5s7vfJERl3OU4Iw0Ca19hA2Fg/y/zK4mz
4tVwNt4mZsan9GWifg3h5mdDqcVOgZDb3GioE3D0UIN8o1cSbsTUobg238sD5U0sAwHYm5xqhBvR
kd9JnhVvS3FJnJSkFolZCiZLxdivhAtrsfjKQSERmYzrwnfhR+7/28tkZsPy+xjij7H2jEioH08w
7P/KP0vW2N0cnumz4BxCg4sLm6BlL0XcnU9Eba6BhJSTXCF83c8iNSQdJHe/XhWQCOcN9eK8gat8
VbD3sulK7wdaRAZrQfIjum9LxjKP80NADGhqjcUCS86rgQHjW0xQVtkqwUJJ+DQGXJc6FQlVlqjk
Yvi5nm4BDxNwxKwhZyKHle4u1NFHatn7XdkuPbe/H+5lJwSRDA0cQYzhcYkOsLuHva8fazpAzDRX
QYz5dvx941cCW4a4ZsUnA0tFztBsd7vf6sY+KifrpvsIYEGKiLDwyF+YK6JFlS5zY95YSpXofIok
cYiT9frcvURvccy9KzgJxBHHwqGhcOTbHNawwXXWNQxdGXsTdSk0kd9XNKhwr7Em94TESjATbJar
9TVxhei3fe4DIBvWDWNsO+lmDiC0XSOdW710HkEjv+oGtrsKBsLJcMSumiQ+u5FBxkzbFCLdyfY2
oR3h6T6n/nageBiLZexRmjLCO+4WsTWstn3t+oRs9PakXQoGjtz6hGQjZKdEQHO34NDSP5Kbz9Tg
rTewIH2G9/Svg2Dx7uXQuQnQ9Es442CNupbegyQLBNiIejguGINN1PIQAUHSOZKeQsQw93UQETDx
UtBJOWVm8A4xJh+7QPsQakALVRDTpz0HNuGa2CWx09HJ2uzKMFrzCuWm5vmzp82PaFfIhBbfoiN2
6W5qbgNxfWNoGE/XL8mjKbV8K4SHFyGdBHrUDmZjT4w8fL2C/AzQhM9aZlsnYcRgQY+IoKW1L/Xo
k2Wuq/2LJPwgneTsX9/b7zQTspuKQM8uGZ+pqcb3Ig31sS/hFSFlfGXRXoGojJTLvWX1Gw1VGUYK
pYNlkv2fN8V1pWYAn98be5AafzFwbXBPxx3M3p8Upp4gE+ktoR7rMXS3yj7iMUUHjFZy0ZAvzKSW
wZjogqMP63kZZK6dotUblqrB80gIlR82VcfCwC08EBWB8+4xDvhgqZZJm5Vl4qQQaC34Kzm84/8M
RCEEYubp7GcTZV2i151jX1VOxvWtjU0W3jGJRmLs32if1FRHCApCDVF9s/R5crA3JoR2jw0Pwx9c
GC6Iw1+nYTW4YDb/jwJqTuHvGINpPm+aP80bsz/owSOH0xur7oZNQths/US9xxJ58TmYohGQ0p8d
xASLoRC0bpRiYEYLB8CYxkmDvUrjdZBL27O+692AR6VXaAtP8bMjdq90s9JzanwyE1RT2jGVY6y9
uCplzrPMr4stvxZaosEgbwJnoirqsOSsW2X/q3qc2JP2bMZoHgsMze7SM8lBbMAr8mOZBxGvM3eG
UAqqrNKvxqd97gc3D+R2mOIFZK4pJhW74u+teVe2rL3zzelU8j80EJh6/g3Ad44p3ehEQqbrPEVk
TcNUbEec276Z6PYlf7OEmDXTlGsbAx3YxWHLtJy/Qgo9KpfNtWbAv7MWNvjA1HZksf5gl1VJp05L
uxjohCAWmA2G+zNz3kMBOdMU18rG6L+FKHL8oZzreynjbyg4xwUOq20OcBHrD3qc+eQiqLo68Upw
LSRMbOvpHdLCM3l7OKY/OTFk+aGOZJSQB8vy2TxAjW4QKl0kvcYG3RGmTSVoivN1IZG9cJBuQitv
cTeyn8GEf40pe9d5UVc8b4/Ix2ZbW/HR7vONMz4AU4Oxuuc38JABY4+uVZ1XFv7eELc2aY0sASbA
Msp7qzjKxaFFN75N6DwMWhiiCvS+grbSG/D55oLgPKKW5k/VbqPE66Ymk9+g5RBoBxQ0O13+ZMM5
WAihvMMkYNT7WbIpa6/7Gy73m7/jFCacFJyOlFzlVjjRTM8YgaxRWyv/A6RrQKOvxyHxpRHdryNw
rpciLF2H/TkFgWLD0jcBdrutcBmCvl66fGXkqoaIezHPAE17S/tNkttRQJ0eF1hfXMoU/wVr1qrC
HjkQb4soH4DIYH+LoZl+0Z35c1DYaZgxb/D/BrnIK6aEj7bwz5kwqBqSi0Un6izukDsoYoQimJ0f
EmMPDkKah8aIiCfQs5dmS7E4vyPLBAcryl0J7ghrNbD/dwvKiGBV2NVTFYEMD5mxbm64+Tk4wFHP
VUWVvi+T1Vwb9GSi1CiSRovAgy0exPLemFTAt+BGe0Ar0MKhd7f0tupgRdr68dxijraXY7zpTayt
hhn8jJb6+VyiToQDFrE0uOfPlzFG7l/RddiXR9+ZlS+4iLQhr3OawJKzWEQlsnNLGPjyNH9E81wO
d6xmfUFHGjbLLeZcjAkaOxbkvkbAQU4jhwLYoDWbIBcsUG8LubhJ2+N2EcSwZtgqVLB0kQSqhJhZ
wKRx/gkSXzUf10xGGpjqrr/PFqBSxy+ON8k60fYA7mMy+TbKxrTbqs1xteTeqDB4BMok5xcJZgvl
anDqUJHPA6gKYsdBQGgyIqgcD7HsxmqfQDV/IogPSkPFBtW9korJ6CHmmf1O3Y5KGJgKvkrIUFZ4
GcgtxsqUNLQlAuMyUAYmwMzA47pKJrw+mqBfUBcv/iOgC9sj2AjOoA+ymul1r89sK1YEt9HGbG26
OXJBpB2yzYwMoZ5rGFWAyRLF9AZ/c50gRuxlPrzCVHpR3DbDIRSPs83j4OtstPkvQ8ROvVw9ivaI
tXf/26kmzSLJga/kAj38VukthAA19tFwTGpZWZA0JdJdXR/+co032jLXI+RhMszKGoCNd+TfNg3c
y8BZUZqOdJkONf4wXk7yA9FhqjVNlf+ybOnFjqPYCbZxmtqokf+UGwShCnVLcALo/Y+mc6QcDUbg
VGgp9sjZpoWpjmEMUbu7KFXv6bku88u0vGqsuBN3Ya59iG6JMcOEhhza43KbUU3C2z3y59Cf7ipo
Xx+gfcxl6aOF9OqMHYpxOklnr1kIiDlVxEY4m0IvJW8KAveynjDBTfrWludGi0aotb4jV7E438fC
yGNR0Uo6eE8YWv2eknnChdMI3FelpVIXcQayGt1w3JTzmHqo8a4RWzVURr+2xaprG+ioqbm8DBLU
xr9OZRt4OZyHW2HNCKe6KTt4gaV59nnu0+MhejvMUtn3wm9UsGe9bBzfaE+Mn24QnBjvW9dFghhn
VpiwmecdXiFBCQo3Ut3n9JsyRbJsSEYVl1BPAj8xCnpweiagQQLq6WYzVxdD19IPVyQJ0qPKG5Ng
Z6TQ2v7nJRiQ0ppAV0oP56VlyIgnBftTirB/YjfLM6kOKh2cduQ7u77xZO5OuZje1V8tAkvzWYxe
rl27RW5HU012THZ2qLCxXLwEJvq4c7n01xzWdN/0Mso/VwA+0QYPz/uietqBE8LDcPopD//pX+Xm
wZwpW2YdXS6Ufmsqcf2nJu4Ch2JC0zqPMBVBJmZiqTgo67e0QF2rn0ptYtRSyVtcE61JjYG0fK9n
4l48cU8DEuAqGpfxZTI3jbzw8oeIjsTRbpK4f6DoZFbF7dnWKj6XrsiSczv36G45ayYVbNozLRQJ
ycnCy0mUyEw+97kTIVFGlpKh64esjp1yKaMFTYsKNZww5BkWR20MUPfN3j2FTOyTVc6KUyZCzfZ4
i1LwTVgvBugZdsRqqbofRASeS5q5A5X/qlXcYAcS/gaAe35T+G4t4Aj74sn1ITvHwBa8maDeZnEW
5TVA2T7lnChcYAssJldg8x/+UQnZm7Lmi+tlQ+yzAxjjO9Rt34uVOVd+Md7kYMqsCMLHGhcTmVrA
UESRT9KM8qyhLxA4MmO8lCWzjajVsDBUlgtDrvH4qGs3Rrho27zaQqSF6KcTbQQzm9HgJ9yTacGJ
7XLN8+T/SEim16uFLvM6Qh0cFakQ7Kw7WtupG4NWXmUb4G1WFX8CgL/yBVRBzBPFVJWAMpnEMWiV
FFo5PRGWH2VueTWsXaWjHcVrl9Qvp0IkR6GMvUX9ADuZiOfb0dMh5rF3p51xdY3rSbzZgwgijGax
w41W78BmTGb4JvOCJ+f4udV5+1XMxjKGdL7+M7wW/mOVp82/efwmK3DKAS6U8Fs3VlEzrxFLTle7
pEKTI/WRf/UoKqN1Z7EcYkt7pNe6l6RtLZ0PdIeOFxJNbfPaMhQCF06EpCAd8sXvwRgaX+Eq2RWX
Zrzk494XLoouk+SddEpEUbBTPIUtgBsuIYjPWc5iJfZH9BqcggDyadtnAAONBBlb48DlKPBzp5Wi
+AGiVU28V10zZUjJQ4UTsWLCV6sMG6MrivydUqNjISZwXokroN/Wj0LA6fbMgnmqwFBh9pJTd9qi
7Iw2eUd6OIjMvLApOtVYK/3TxlLO3Z4E5BYK6/uVlH8waxXSdJFlmcVGoDjkCK6PWo1oGZVzr32p
JxbScJaOUNMTgG4Bw2Nn+DlcBn+rJ7kLknPr2BnQVLlJ9nCOBRMngc5f38GuyDWVEZvlbAso6SX3
u/5ekJo69P5iELJrxmjpVBjsARVi6EpAUwD8nTvjeJ0K97ByDcM8dRSszzP88FJmazQKSCtjA+kT
+vOhzP1hjU/uv9dnn2apDNltRfVj0pnz/Ei/7IJWpoKJd40QuGLIbnCP1N/9AoN3KsRTPlrC8nwI
v0CjKEeIWC0uP2V5E71vDzvKn2tJO+IPdzE93T7nTVF5BLxJIIutWnUXyzg7e3TUdwvhheTUwdlR
xzFyvlF3lDosekAopc6WfSvagjfdNA9atkMBcdF+tdsMb5k7X4Pv4OXlv8X6i1etmacyitdi76e2
ekQyuVlviKGKReR1phpVozZiukgpW4HX7x1OCwOCSOBdHVgBTfz5sVsEbrpDh/7kjsoGvSj38oCK
Yzmo8r9JOgBkR7LIQhaN6Jds1F0BQqCbqoYylgFg912tUNBm6F5V9AkNQXV5ypq4IsXmrPiA0zpE
xIYKyuIPbYjznQmA8DE50r6uABZxziRNHciQCavcNW1rizia2OnJnhzVYDGFDC+V+cxFcOLwOq9L
hSo9YhF17AJXBsYIBNXdiVwYjNf4o0aza/aT5zGgVXeshmYUL4HBPGDDnCB+WVgZkbykPkphSxeP
L6XD9S22+H4iEOX3I1YPxRFmBA1WMTfhu6/uipIBAyhghH/dq1VKPMeHmfAA3PDLWJppOiFY5dJd
+pcCL7T1GGkrlmbjVrFU3RkNG6huvD+M1cV/PVPDJ5xzAgnshZ0NcaPqhRDV5oNcciiHC+Y9vsd2
uGyCKTLd/Q8r0exoDQ6tqXg3W8PqOgVSjVUO7PDmBddCycIvn/I0hi2h46kT3mP8YZNj/zhjVyWP
EGc8S3pHAMi+DqGXb96Hm8JKnmudjulV40ao6kKuCV0HZ2+0RpD+HcrAn6YYLbQ2NL8ARJbUBfJW
5Fo/UvLLBHkxklpqEfy0R5lLGEa5WoQ/0w4HVMrG/b8w/x7ErBEAlxPRjT4EjdMPVRmH2ScQ8U87
3mIg6h6v9RgBt1oMMo5F2tdSsnxQY4DtlZiuQ+TkaMeAM3DU+aH43SX6ZleC5nuAAVe1iNP4BC5c
i+MlBstm8ga1QdcJGN83SUG1PpKuybHzBX0LQmIYgZXMbj0zdBCfuJrqrLrK4/0aZml/913TMjWp
OZZaLQCUOySIMb0j13BFEr8YS2XewZi5PXZchWBqctMAL7LRkRoJ9DHfCsD7WrcG3IrKpvZju0LG
2mxLIJUQ+dHYVX8sG7sRxt2wdfcjwLnMh/w9kcEPpi67Bht4XSmXjnNI2es3XuwXGIHt7OXzrYp9
zcdeLw0iZPkrSBjL6CLxHAQUkNypblLR9O/YIpUd/LKh3MOdJLmURHuAqxdg0+nefPqw21DpWLZR
RRHo4aqc/Ys18pdUCTm3FbuYXebtsgVlZ834RGl/5MMrnoIXuRf+BwFLxQ/Gxqz2BQp+soGcOuF6
Z3s54OGoFwUbxrbmqnU2C4naWCVb7XDi+AaXXhkPXeEaemjfrcpDAeFkY9VzwHfwxpHROg+QxacU
39j2/FwntrBH3qiDNOaSSsVkM1YOUbwLCAlGRpDFcCBGpB6UWmht52dwqMe/Q2ZaU/B5u14pxx5f
9gbx5eD1Co5F+239ZiS5L252CaMLvC4mG790aGY3Ic3VJS4ksyGAfnhiB8xP/nFa2z5oDQ5MHlDa
503Y5As47kHUH04LP0iP4IDImVk4XRUBuXaJ35V2Fr+zw6h287cCawWkvvLyDWRVdFCyTrxOk1G2
7j93PjujP6pCvz9xJh8V6VkFxprjlVKp/Z/Ld7F/CoeRBFPfUf92By4No0uO3dyBMnM4Chj6q6ZL
H9a5cGGCDjC9sRMePFvJyIGaSeKJynjZcZoAPHINmodAsJqKyZaRZucfIC2Qupb1RDI7DkLU31ZY
bYjHV/SgIwJJrDOrSuBRFZBBpjvu4mRefjT8aGAp7Fmqbd9bfY6kbxjRs/COMcrbgQyINnEbOxJ1
WkBGWN8dpfAQZklqVgbGRMKL/Ya8etr+SRZHPvz4ilH1lXW7II9gvex0xuzSPted8+N5mvjPJKiZ
x7QjAxwb2cQYW9YjMdKmft3/z2l0xyS4xYRK2MWCrIzqO7KCjlH3Sql0hvvhbohgcgeMNzZbvej1
HMnDow1mgW/wr6WUkdmwX/a+zUiQFP9VW6dLPxt/g6hifCb53CExOq4Ovh6ah0GaYBF0GeZsDXh4
/uRjZr7462kVDVZJpRlMMStk2spCKLxHAhVKvin8ySlvpdAoIqn83jEs/+nVr6EoSdvyeo9P3WaX
LRyV9BUwxLAFlWfkmWwgs9ITsobEe0gFCHdGpvkgrveFYgkAXqbONAdk9NlVLw1dcItqWS0++Ksu
0EqtgcSaBIaI1+YB9WfeDtaMC3FJFkIvaGM0zbDPnAkMxyOjf6Xbuurs8ecdwl/LBgJko2ndHFF+
be701OuvNqxQ8hC93QGPdGD8wo0/A7HsrwFvOehCxm4OkvuxHHkoSfayaD5/qA1pX8uXXMMXrq4T
N74+Tuk6/Fdc6Qq0dM5Jp3Qa8Ae/syBU0fNH9LGNrGTDZZOBPqoMDXpaEZYw+UGFd8N3JDRjdNkF
SpjQh945XQQEfKo4e4PH0/MkgYMURny06riD6IKcgeKqGfGnWHoUopdfsVSbWkPtgHXKxxzMn5Lq
aDckBvIbEem0v0hS0wwXcgzQEax3e4SihZiH1SemVDr+Oo5UqRmkJJeYayL0Co9Y+F+1dWWD9/dh
YLLSd1VSqZJATCmun3WjO8MY9LOnICHOiP7ZSVilevvgg07Bf/Czg3B4B0QQYExS42QIyg4InngB
eXc8k4o9+ZMVomARKFuVcOHsFu+whevoxTRhb8PnW34lOAix0889u3/W0pUHyFPHIfzhimLh0tSc
ijMPiKRJs9HViuEaAJUvKxn0Vrm2dtDVFp9YScB1vkheP57NShLzzJp2lno3nQd3Qvj6IAQTQbTP
9t9GuoDuOL8oSZwv+UPxgt2Itsc3zcY9SnOLLNZC97nvwh0K5u0LihbN1bQzZa6bhHpFzjGwwOi+
WHaD9BRzMhWjEzUB+TIvcdlhdiEWJ31twqdJ9KeMjg5hRUfBzOgfkxpsuC4/z8JvhCvZEqm8agbU
p603wMahuz+h6DsI3w1dDJOqPO50GVmTo6ftMNcX3ROC26ztoElDeJjF1MzYD22EK72jgPM0GFft
OfGu2Gf8LB8ICGF00Yb9bH14FcDBq25ppFd016zJMBXV81K1TDL+YcomprTx0tHHxuY4qXbb1xtV
F5ANJzevEHzC3Dqy8kQV5+4BS4HkPNBSPUWbGfvXVhPY801aznqmunb12fQYfFaxW7p8akiNNMZs
sGTOzJ+y8w4WG90I2H4yul4TCnM+4DeZyAYu1OLiIyfZbXbr/6E0XKOIngqjpmTTeS52lO8/mLc+
taWs3UKyB5x9WiARYpa+FeyH7T0mpt+89BzjQ7khXcI3ddzcb+mbRki3Dd2U1YXpB2gZdS4IeEu3
cyiWDvOKlMESN19HShnlwYiGjKl19ltrnLB9fouwzVjERKjWc0tpaf4Mg6WcaFweEpoYPO3k9olf
ILnJXwRDMTFFmVYUTytrAIsFibmpHeQZLxMQ05i8tCEKGsaMdCxblcRC8a5SpW7pdTD0AE376Xgw
EXHrUEK57OFzZLFQV5kYyHHr+x3ESxyL/RWbY0HrP/hKVW53JDiPSgo47mZB0asT0rPDApckaAQD
IBLDYIXo3xbFLBG/sezyw1Wy5W5FsYVGtXjKvGQdPdom5QqLtt/yggyJoSElDViiWUhaHiCsIGy+
5iSZboZq2wpvHXERvpiJCQmJ8NHFwOGSYINc8SDQ7+KDdJ8YZvG2FqCkfL+S36QIa7DqJSAjfOct
5cuyke5SaHmGJuOAjqzIW3MQkGquykflN4wJHi4myjzIC8T1+mmHdNi+8VDrEyrbOL0Z0DKduV23
EdEQdwgHar7qff9knU1re1bouaIG07DFusnE3KDEAqDy9Oqy8xsb1xeqq0wrAxY9rXK5dWa1OqjO
QvBT+zn3GWzzdM/bULhZm6iCDUhnQrELSHaHVOiIlDhTcIN2GYaz/SxRIkPnp+F428doy0dai43O
PDj0L+wepsBVFJKHFDWUy2shfSp6KpnSdPwf5WDjn+Gp+Hy3FLodQqr4fUk/GUkGB/t48C+BpGb2
2fd08GxN4G5vs8pIOw5fdUbFY850+tHkcI7k4nC3NjDO5KXVvQs1S39xrEkhQM48HBoscMt7PJ86
YPNP+Mao5gN8E8gbp2aQTxRd/hkPXeppMSG69bNddYm5HJ6AIpOvzUD8/p/09KMK1xL8iOZHqObQ
CxAuZrb0ZJD0rEerJhjOTVnpXLZqE51Ob1DJXiw+6Kz4jFW4OvR8138NUEFQRRdk90OWSenGcOL1
BNwjQEh98o6m70JKroX8CWUBhQ+Xn/YZW8F4nWMBIVNXUQugJmtLVBz5XujAbmKnfOXr8JrgeAcd
Usr8tdgTYJSnwG9rxP+40bEnxpIBxoT6+I8TGFBirZSzFp7A9q+ZVuGvKpotRZpYoucRFEZAdkTu
3woxTDyVqr8dVMWqiudwUbDF0YUPte1lphXghyolJfSfqIHQ32A6sNqFViC/cWK2cwJ/PeR4zTEF
+ibrqiRlWs3TQzVsv/s3k7TRNUrLorrGN3sksnD+6fnmLx+UGKmnhqZtxqrSABixCLWZLQdgsxcp
YEgbiDu77+XmdrsI0/jbQCSsu6O0YkTchaHZLWo7l0lepixs6SRfMOuJAhhdRoJJ8lwajNTbiGuq
3cpVFX+ZY6McDNKFQCJo3dCMBGMrgdtlIRC9Y//aWJK89ILgG3Vht/y0MBD+scFSZB6EihZnZZ5k
eXSKsCgEDCxPyLl88NfE8bw4K5dWzW49PPlQnEEp2kUhjXQk9F052wo5HqDinzvDsY+M8RYsUix4
GIX+WVZ0+5UW9gFbfShPJjp8At7ccv4A8fFhb9XKqup9pesMP0O12r9xc+Fiasb25Exj0AXg1Ri2
kpZaKwb+NWPkVRMN/7uPpEAWPfKj5sxxZ1ErHHxuiuyqaPDFO0xg2hODzvsiJS+K151xyk7gtKmD
W38qbr1GKea/4B/y/xhc2He9blYhALQtN72B4LoDbOOCqEDC3eRC2g27CyzbblM3uy5MXuq5v8UH
zUL9OaL2tAVWf2vMrLPNEWNEH7vyrW+NiEmAewBIgDBExbFpTUWnqNDh5Ba8eEzUxA7HG6QrfLZT
G4vvHJr3n+vj+aYuovbvT9MPjD/8D0KEMuQsu0ZlirOALmYl2mahhc/GT1tz22qCqfm5GX8TF+OB
LXYS8kkr8zk+LTQXZ5eLpInZpb9rnUfj3JNu4fzw83dF8HKD0w8wSygtSzyq/KyuuXiqqaKqS11L
5c2XRv6GljApz1fAvs5fVOqCoHEjMmu4prkrs7PxaaC7EKed2vQZHk5pWz0eWhpw68r8uYfCroa6
enecTjRXVIZntDzFajzIV4kJDbcOm3bNcqIU2rhuEqpOcuiN74uWYy+D0vmIS3ugElFQVOEcwjHb
AJQzOrmwGBLHp7kF/WJJ8TxMNbjcZ1jeVBoGovfAyaD7SdIpeYykZQnfb6Sb35UeHl6hdgNVrLEf
ovPkVQIAjd0aghp845isnFRVwQ1B2p2uhPa2R6gJyWhV3r+VZG3NE/BeV8xoSYyZ89QD/kGMP/Tx
X3oA7FqyOgYKQoAKi+ZnaRZiqDJrhla/U1yGiRcrNfxleXZDN3LsCspZjYzNPAgJ4GMudTG6O6MN
5jOFhHKlokrL/C+hp+8oRO+tBt7FKtnZKuHczbkXyaSeeUsJj7biMi2MsG8PAViHj5AYR4h436c3
mJesrAzw+qU4WO96emVCXC+rRxNF1sTMUKZu/k6AQP4qcpRd4WFeD2ba4Q8FHGJkEVULdK4m/QWl
GUczYrmEVmWUc71FZvYuhoxX4te26yk2t/nyBF19LL0BFeGeafqXWyAcpBXW8xo2aEpeM8gJu2sv
PXKAZNP405WeeSrSQUCge/PWlyiCtZhSBbN4jec1uccJ8n9ANHXqIzc5+NAxVKpa4l8dc5La56N0
gslD3CGWdgsKRFyjhXY/jOypIzv2Wd/Bc3VKxOkXU5CYlUdZI9b6G58512g+B4Ihu4Ub6qv/YAyB
oK9RI6FUBUc1whRUja3JE5+CymIepqUho1kniMEDCpsoWZVZEe1MJqqcaDnRrOv7QoAPOpxJYf4M
wXFjn1/nfeofux+wSKE6XZPSNvVHTCPlMmD1YAhoI+VwppEwbwGoUa9NOy7q42LZSYv1yo+Pf/0n
LZcDBsr4NmhL8fHaf598DAXYAu3u2vdu+Qhm+7Qw936jKMPh/0cN1jSI66iA4l+0UejcVA2ObYSX
b1GnbVfyTd+6y7MUMcPHFLaOL+NUa/G944ejON52/50zeWysYdglOvnVtJt2APq8LCGmNTAYncch
BFQP9HOdxFOIiOIyaMQlWCZiXJceiA3rjnM/5C5ame3cyawZk/c98XzDSXXHhplrHkozu2V7QEB9
9TroX4fxuBI6EG6yXhU+uZ74FLbnDfGhQQudwWaMV57WYBZLtPJEr7VYePY6tToVTdT5fpLl2Sfs
edv5cIseH3CwyTq0RbxW4mkDtDTxNsDK1e4QCy4Ip+9TqUvrmk5aNmpJnUs3VONaHrQInlPMwOBJ
YdO1sdXoA77aCrK25Yc6PWhYr7R+Lawpnc3ww3kfGpCZ0TTm7E6qRJQ+pVEAdD4permzl5tdtF6d
TmxMEvnlcr8/v7liUckNzZ05aCC255p12YtTF/cmnSPgWJWIlrsqEAaXUhvM4chic5PxflWibrye
ypj5cmFnfz73JS3ATkOnRJn2lybCpitNCfDv2CxJyefvQ+JOSD6ojwLyRXwHrl40PTX9g/6saAIl
bs/8Id+f5AmLy1xQOBtNDLfS6kSKjB6XGvNB7rYO5Td2dLyiwY6SvTYydxnQ4qdKmZ14e4tEFys7
QoQcAJ1jJFfA4w8S8zx2hrxMA7S9vcDPAqLrajtR7Z3QhKNGQ4tUaR4P6PfSOVCR1nFMXzt6xEJp
YWatXHbMrO9hed3kMz70SWBZwFt9VKZKw9c5gpW92SRXUQlqF/y5b684dQTOS+x7ARxX2hZRPdgk
dFQMob3U/tpzBHhSAM91lSPpX2d+emTqZSru6Vu78DXerLEvOAX1lob8wAQPG32qmoCp/l/TZ+QJ
J4E93o1t1M5ZNxm1k8aZhA5AKZA7Ha426ev0DPQmJfERnr6s+li7avqEkjCN16mi0VNb0h2KYJzq
uspwixl3vunfUp1qRXwjgXonxHdhPgan/opKijx8Tz2iLXhhnxrBuVXYzzrHaByZTquVuY7C9xWu
nHc37jNWYkha4OaeCvt9Sze3HWF7eKKz3ziOFK/4qlJR3cGUytlxOySRFwWbHhv7yG1eRmj5z0ut
KSGsIc4D3epZ6ivr+e9PC+7v7qtXDEjI1SKtrZS/6NLXaAQOmatDLDHCwaJhu4DuCLGWEW4YxepY
sfkKgZBeBdfWOGtXPMVpfAFfLb/Ne/lbtKN/tItPhkz8r0nXvbRdLINBlj1H0Oah+RnQxSh70Ktl
+p7sZay/DN8c8UUGWd9Czw2Bao0bcfW/jvNcH9F7uiJB1GcBqQArETXycsXH99EpthVvwEsfwzAd
Kihg8PTWOlJV/bdgjggu6hK8PMkDMbe0xPORHJNLL+/dfNSCSQpAWBAY4k7hxWdmaUCH1LxAstK0
nrNiKqYiFebuKtTwM7SXkjhEykAe9MLgmkdl1Dj1E/6h+52mjqoOHFGKVv/CecvNhR62MdvvVoL+
8DS9LCS3Owwe6E1VQtP0vXBGIMWwmBjNYddQ4l9q1ffWRFS7KcHCSNZxfWGHnTUZv0EVggHQ6aS2
KyG3hQ9O3Kv7+QqrXoSY45tnN2n2d0y+jWxt9CnoYwtdPq8YSB7B1tQy7YiES7NRQoRaUUzDfsc6
3jC1WBLL51GJjyR4K5Nl8igxxIxbZ6PES7lfDqqNYZQVFrzqtBQ9/4ebTlsSgXCN8rmCZfansWzv
uUZoxsv2EOJDqgFK1DFkCUlifwK9mbGRIks65d4xWNbrbJC+ATc4F7drMqagozF2e3v+/ePe5Hyb
SbOu9goMhOLGehOwSTjXrfRB+2co2nbd6hcNPcW+LbNW4EDS3Mg0BtIMwBzcEndMdkz3WnEFA6Ig
Esz0k0HSlerwlnfogVHXK6hybCRGKPMpXCfSm43q0PL5x8TPkIhTgl6Fk3LWABFxU4dMWY/LI1CE
KX/htbyh2V46fzDYMkUblpJ6assTxdLPBPI7ZylQxxBOJK1UT7Jwcm4zH0UWTyRFvk9pw2Zx7Mg2
bw06l1AT4rz6M3uwYTrzJUcQx56ipBhiJhYz+W3T0G/vug+sBif6Rhyby3dR/t4v1NqYVKUSum2F
WDVbJ9UwossEXg8zQm1oHhTnldH4PPLJTo+Fm2F37/RBUpykIZU6UL8hD1rnqmNRKGAnRYav4wG1
bk6No4gJQ6dZceV/RtGOijQ/IHSnuxOLCoRK/NjQX6bKKAiY7aKBxy8wmrLOdvzEl2URoKmGXG0+
t5vHyKBrsT8CZVNi/hPU2s5voSuwsNOdVZKnH7JGrB1bT2tyrqlboB0dksFnZncftjdNrzJ9ro40
wiLjsNUiOJTrwFPoWlD74Nv1fbz0SAcdFMAIj/9sYuoH88USTztW7fDMWusFNsVGm+OWhRv2811U
V/hWGYhQ7cKNL4IIJnCaaO4K8nYhhRWkcNCTq5GAwbl3gJHyLIvefV6x9lTtoZEfIVwiqelkswqV
ADlJIv3Xig4JteF7uQ6554l2ParLMrrc3GZHylQ1bx06rugpNfLCT9d8/hrxWW6w3EwyCs1Z/U3D
EcieSigIuutzGvmg5q7pws/A+Jxc3HW9XsipFfj50fuqj8gdlIFq/+bmJUXyOPGe275kygg6uzWa
Dl9aGuUXPhZmMOSPZ95/Fa5bkvBgKfu/IjBHk9+Ry+Q7xJkFwMUlj+vrlgGK6lbytXFMpREvyVNC
B6NGsrfQDAFS2x2vLeSMf8fviWNUFVafnaWEfMa5eAMiWJKNGiBz+PlTCEjUz7SxFQuT+TirseYc
aSy62ydtst5diktC4oez4kXKTqb/PstYI+YI0ohyse9aLTH9JyC/cs7ydzY4MmQYteyeNwPAQIYG
2eCqcywagZ34JoGsDK5uUbEG/nb2Kl6cml9m3TYANS06hAzMaNSy7BCnmLjgG9jRnM/VQMmrSJAV
qRp82r5gG2rT6J89iXbkp9+gBOY8h6/g5P+Mchb2LoehmMB/5iAi0Hk9/5pMl0iRqYz5IfNKgoWe
m/KdWfoNqFHJK3MS3m79JQk47QLhegyoHRDdadtAO66d8+785lu10/Lj4/Jzwe+xGl5FsEjGE+nZ
TbZL9BBYLhFmRFdYMAiBJWyNPV8SHX5/kheZg5ihPYG6EnB3sglAzlp/ia73CsM1dPLTY8Q5AcCg
ir6z/u+yw7vqgIQhrVFQz47s4Zqy7VKQbL593jWNmYuw1CxbxvmULNf7H2c1xenaewlLadn8v1nx
CvRZC6HI4tfAKLvd7cdjDcDa6hW+WcxOHHh9Icfe4ARl6kE4sFUyGkzn/bSdx+CZ7PAohMLvqu/O
J0u/jjmtCd2Hh1YnDcyHA0VOyZtpoWvEdxE6xhEkcPoBmxlZNzeiWoiMxYDGTRjZj5D3rMdWPjWq
zlJ64zzms1laDh/GdYHoNIXazDXIRN1uHq6snGAuKa8uKh6aTnzFJeyEDcOk1+IMHNBRn352U2Jp
AH2SEf2OOAfI1KRiDwb14mkKLCgR3oOWLMgbKz9V2rC/Oo10f00IYAKrwIsMAzR7jD34x/2GPf81
VtRoR93fD7SCW3P5bG2M9nm+2Fl44DOmAlgrW6Q/mMxv3sAUQB+pjtjBn55vtqR1CDdpdFxsvBvb
S4kWJG1dXo/X2ZN0IYpfN6OOC/E5vqoV87uheQfLmvcUuqTmI/u9mTSR7h8CfVLkPFVukZ4JlbHy
W/PKAYbpHaKBd8asTfPGPAhH1olMkMoMfaMz9EGqIi+fTmxpftGgeiDNqmQiAHxONomuE6GrU+9C
MwcezVnv0SJob3dX4rvAv+bWCvIHhiKbuACmiIFYc4wYBFE1nDzmtg9SLYAKXsafWXsa7RGHCC4g
rnHXbSrtVvOC/6PfTZMQ5rbbkgYKNsjtAIhoSFGZD5ftC1pZ3Y8Vhphkl2KQ2jposX/N7idvSHir
GHKQWljI/uU+41htREWcDYUSTHl3otraoPrN7iSzFO7fF1Hpr4zZcQqAAJE14hR4qYPVXiCXVrgA
TGRdb59u9PHacjYwSgKlgApdoSNEx8h2QRugQyKllz8gTNoYGMJTJgUEpiv5uDTpr4EPP7qEt+8G
iTqVJLfOUU92ru1tXgPT5sNYg/5O3Jvcl+i+EHahsyGFZdrgUiDbFnebUn7viPhU+Um0ZOZ6kJge
Xsi46pv3Rdu2Xcnggwgk66V5UiWd340yqx3NkWZOpRV0B+IPJaxfsq9Xsd81XjA0ARjtotI1jB/g
rgDAioLiTD2LhIIueZqwCIC+tBMalK6lDFlNNhKDoSIHH1Gh4VED/aZCw1THOsrtfe7xrIv9L/fB
kMzI5WqQYSTg4cLtFC4iQtzjUVDAnFDQ74GLf0daEwbRlfKj7jDC6jTdH0R6RqEbqLAHAQNOFmyw
xDDkDjloDTg9oqNLu81k+23yv4BcdGc278CAdY8Urf5I2rR/dufHUjEu71bJeqdNilWHogGvqeJm
qoaz/hhDCMF5RcEidWWKqgfVjFej9ofMu/IcR/zeqy8PYNShxMyZimiN/SxzQKt6xBPaKYMWfyi5
q8m1Yr/MeJP+7bqyf2cMA90ea2rMg1jUvlXSE9T8mqyEmqc4ul/D/m/S1mPr5qmHJrGYG3DsUhU3
Wtnok2rZOdawfC7QoZLpPNeWFxLvLnTLSm79ySpZdSzhYa8BmslIOVt4OYVNfCs4W9otdHAxzam8
9ElabNbJph34li+BlEcVZarfiwl614T59t2LRufzNCfR8ixOlft1La6d+eKXkBnU0LpH8HLSvHVp
Lf1X8ESFhGeczz9uKLCYiRKD/EK1zgN01NXSb9kDhUL4q3foACE4JhOf+b5Dy3wuDnuT+Jk4PngY
uyjNOaK8pgo2P/WE0bWxiV9jQL5fDSguOoiXtcMDDHHYkpmgRF+RMcvRo22eLN9GjNzLOGv9rKla
LgNLSPXSKluyjKdj0nKSwLvF9jaJPua55U4QLtDXCt8Gu081aS7l/NSPl+BAmG3fnb7xJp+kHlES
R34x2FsKrCD0QjUtJfUXolJ9Q1HIhaNlP0ZtN+hKFEGjHzdo9sPnwDc3SWArVZvrWIhcPT6QbTeU
AzpKGrJ8UrSElOEQYHOSrKhrGB+v2k7KWXHpavJOGlO3ZazgagIJnNW4iJIAUbgp3/QJ/N2KVSj/
9iXwVMrHNwJnH28YE7WsLe8kZwGW7vwFxWcthYJ2Epzfqx6wmD9LJZ9H/AGg4UhasvsPE2ufFlHb
75qpcO2OuC9JQpLKHLgoSmH7k1fLWfgAlfVQMxa3UclF2UKTL/BED+7FjHYe/uhDu9OdRYn//KcD
SYM21n2zhsXSTftHOrccJgXVDsj0J+MLZ0Djop8HK0WEXQlDYRVz7AyhmeF7Haz/S3/9pKxCzBQH
deoPSX8s+5kQ5pIUVGyr5JV7jvG6VObryZNAYW2318+xGk9jK43cJigd7tkQK/YAp7phrIlu3BfO
I+3soXebZiLG0gRyX2ta5qasKOsmssQ62k1E8rRaOfk3eU/xR1LZx55zkKsxJak0sZ9YjR91hN+D
mVjOJcptQl0skGwlhWxNAoN1DA9JFWt2KWtiDpu6Y5wkUq9JfQktYaCOLInkmnl+ntku3j7IAmFi
F8ctEUWYu5WSwqrJ5eezh8h+cINnkfVnLF3j7gpa4gcm4FL2i3zCcMitm+QaInEcVdCLix7T3tGl
Tp2OyNecKS/COXBiYr+OzcopOsm9fl63Bhv8dQqPog3ARjXhxnijOLmuvF/cufLpDaiFcSrJzASv
asVHp9X01k2P6WmPynUET4f7p2qEUIBA6g6uwovKCtgLlvhwnMEdM7UmJXOulsaMG4yq3rWxvcFj
aoa8qtl/0sHTov1+vKICYj1TaI9Yb8f8VECOqDWkwWlyMl8iWffwlzlDRdg6wENOPjNbLD9gQo6Y
36d9NpF4qhydEIS+sjuroIoCBkWLqWGXIYRRLilkvlFTruwgqwNMnCIsaulnMh8aM5KBoHBJ05Wh
DmsUBjSqQeXmw1+1LoJFXHL89v7F8FW9HdigFqZetGD1zrmQml89zWq9oPE0soqL1UicUPiT1fFa
FMz/NaW8RjjVuoXXd6m9xfapST0JRxIvIJK97KpdJtdaLxfZgQU+EFesGcRFi30QvwabRV5TcQQT
Iie7DvGyXYRqM4E6KwHTchEKgNQW86e07ulnIoRLjQBdxp6QF3eYxxdv50Y3T3TPK3PmGDjgK7pM
gJEDwoLKVlVL05fv5PtGZlP6m8Im+uGbbnEZ/wYgeaD35iL2UvP5R37TBczFAGDku6zmXshuUFGO
uBbTj+s6grA3atdQsID+eVdzp9IfSwdk9xQUyk/Y7PlzRj6PPhjjD3a3TqeGxeJSQAsTGRfnnnPM
FRqMsxs0vAI/3koddPmkw8D03j863YTjrj3wYeCgVaOormJjZhQ0pFP05IhW7+GtsVNJRu0DV/oA
v0pMH5EcQigDthPRzHbwqd5lYSKJo4nJJxfNYt6BmJmiKfrZCCyGr589VXI91aSyBqYOHFOLdhmb
UomVXfxX0Mp/rq0B7niDpH423pOY8GbZpk5f4R96WLX0pQNSG+42Ss2/XXrFT75jRbZPljXT5M80
EuP5AQNfeepc7FeJj4yL+lNROXM5rpLJadjEHPvNeZCZkVsnjzo0UDOQGhKp4bH/r+eywNNxSVB0
hcCuBhW6N7pzRkoywgDKyS0qX+SnbVOvBu8UOMSul+QJ62V4Pr6Iwj5otdmBDjttJC4DWuYoPd9r
JiDNE5MiUrXx0kwjTcxeTZNd3FTWe58rAbTWqF5FplirBgLYhhFxIL5hKSQmOViYSZ7E85OGexhy
DS2TTSTXcBWTpVCQL1ggauxjf0sVcNBWQTdbrMI/ES4XffRduL+GDRCl8xJdJmvMwPCBSUuEnpfc
ox7zMnrP4vIzLsHrZ1JPawBHpGsWDupJGUPzHhnIEs446uhN+sw5UkCAEU0JfsNate0ClD063Et2
jZQvVLZCEYvOSHRpzps0mP11nfhb8M1MCzDRFRwL+LCrlUP1oSJX+qCgJksws2yFL2W5ovdQkadw
VOGtwiEn4SDXYTno0ihb2Z2EigdxP4G+PQRlbDb8l9TeC6snEleQkOcFRtFgibKTwXevUAhF0mck
Mn/0iwSpdzfPAKy/wcTBUJKx3HnOUjMK7rho+QxcYIlQrF3u8EUo/EtMbZwGqpj2qV3qd583ppNh
vzbmhECiSXfd6rzTIZlYHUxxuhdKfRmwzv7MVGOX/FL6qCVIuYLidd9XIF2/QwtMeZhkKwQdfQAY
cknZ/58/x27qp5GTYqcFPC2ykzbU3zADwFhWZUP2bUQVq/lVlJWu/rkzQ1mLL8QKOIiIqkp6RANa
CM8P8CKkWtFwU1zLOo8zrnHfWLYYKnvlHGIruEg3CWdYL5mUQwnsQckfitTlEPwBjoI1BqkuccEc
v2ssEAhwk29IWwM3jPx76ngKAlKMfk6jE3U+t6joz95F7YXOqWVm0JWqabqzu21MIOt3dZnlUlN+
/oMQnmM99073sg36yf27RKlPjU+WdUotBqcd/a0SV+dPMPqFNFycNdV+fGhKndPo2gnVm7TLNrs4
qXOKT2TtKZC5a5PhbbJUTpmW2azdgvqYeMBss5cnG3Zbpy22903hbN0nL2BENBuY0QVyC3IGz8Tv
eE3rWnd6q/aZwRyzS7P3UFrf3iltIbnnU4sVU0aw9ha/W0dAX+5MhZBdbnGDUFXTlIdLK4wLcjCb
A5/GEeyTOZz6MJMHlKEjIRzng4z+zkHRImiI1O0mViyuhOXqFkn56wrl9oP6yKmNvPdImMuyFg0Y
tjwX80hIBzR94qlOTiC3HaUvlLpvsSEFy0KaZ3SMwBUw1utsD9QCRUAOlz7Ae4pDcZ9r4ikNLiDS
QN09dhckSaaeI0CLHaN67iTmnRwHak6IL++MjKd/Avqa8l+Jgbs563vpdM1aDCvMRwSyNjBnC6Cx
OxTwudZdaQ0Dyyge6G1NZXM1afF4uPdzSWugy8lJNCfYjM3ua9o+VWGjcEwaiqqv74nV23D666l9
0XCOY02MFNlZWiTEPONfTAVeiVbQawyId+TMwlIBTsVTiB2lQHyskeQD+RtsFfwGS6AjxCVjmi2X
1qgviiwtf1k1GUu4h4x5jYGHYJygYk4RhPhorBMQA4SVlJniPauixkmrm48W2qpo5yduo3ycdSd0
Ji6kjDstpcfZX/pSAVbQGf20hk91zQhOjoiVaFe0ByPiCk0QYxTLjbrQrjO/X95Y9a1LV0oEECmr
r5i4+sQnQQ54mct0CZ6tyj8ryc3d+0AEFf/WLB3kSwOMEGN9qM9p2DQfJ2j2izqo4LSyJrV/GhAq
CraKawIb6/XPWV4GVtZ9vpLVGIGq+L/Au9F2ylu83KkTgnhkRfxF8b6igYwiV2WFO7QWwAQx/KKi
Soaf9rbP1q8tzHE0RieMmSnKEo53pzPj9AN700JMdISiuw/wCixj0Mo3cXNcaigUHHogahIcxYkD
//vgbyx3vk9kGRBqz4qvA8Ik+R6oIxN7U/W2ZBR4GRLQ1/waiheB6PXBTV8QtNaO/IQPeyowfCbb
nplkY3kc3/DPCj9mtQhGydDyxpcdu0U/eK/e3fiy5MSU4vTXlgJyVT2D8fKHDY3SlzDDkLGCGh9M
3EwU9AWGj8BkX5CjfSNF/CUYl4fXjwaluYXPPBZ2qGedQgHABpIGEoQeFC2HBTFiRyBmw4/ZmkE1
Ia59uoubFvoamxZas/ZHQMwW8egU101aGixEEAaPdV4Al+tXfaxuEJIyS3bpV4vPsqhRC7a5iaXw
BWgrRXn+JScNc7aC5S126Wjhki/Sj8syO2ZCcqQfmXCyI5Yi7JkvV7uPEK+iwzcEDCNR5JVal66z
IRh4GhAgoo/t3D0WwwTpZLMmFn7xEx2S/qaQB7cO3kDzN+V/gKAvON0tNbOKdJiwxbbD7rk9T1mi
BtaUzHmdTsvpoAviuz856gn8EhunR9+Ssb5AwiYN5PA4PYM3OhJ3Vw5U6TLwK/JTZ2NWwQg/qKmv
5chYcxFsLRggC2qbaxK5RyHvowojzglqE3OwBQJOF5Sn6qdHMM02Fm0iz1quv1Qh9gWz3j+ZyG+9
6gfeoUiZ3fQo8TV4VYEvehmCdxsPDp2baE3b3IYScmSAqodrcWo2A4sIWZq2fuMVx7M0vmuazEJw
zbjTLVto6YYqd6qXFw8nRpADL8UamuszXzAa2EklnZapQmlfBvzfpDMcJwH2W5ZNpw9LSPzZjSPT
uxFdEYN4iOVEZckDEpvfhu+YzKJobCdSOhSBiLMjTeSy89zD87L+tQR4ejTQcCvMu+mXyXqsh5e3
WQknHL4lVmHFlTFdDa98tq2fo/1rShJV4H58B03xai0VTVdQADqXmAkmc3OECSGxOLGPrCJjUAsM
p+8x6pJ4oR78VelMkc5oxAnL3BzV5TBIdpJ1EHKaxufcJ1iIRY456mkxhn/9e+XodMNuPKcDVqU9
kCjIzBliWNdKAhCGLvX4UlhFE5un6H+rp6o2/K4uq1mV0dnkQIWyUOKDrf9CapN28vvkmbMlXlI1
NFLiYdYM6BRfpOkypkEGneM4gCZpZ51r7Sy/XGuNiQ4+rGirEge+s3dWbqWwPA7h2gi1rAv9sNGB
3z7w3dyCTtDeWcBwYn1tLq6FyZm/HO0+2BF+GQOy5MTwFCUi5lmD7FAFjkDr7qYEL6pi807bHuKb
ueExKlLP6udBqmWKctE2BC2gpEneLSiR3Qxy8NVBbiIqTxe3j7+GK3RAJ2oNnYdsn/2V6fMaW/6S
VBgGFyte/b9KRaYAMtCSY+rHT+iTOQEKikYJLYmaMo/4/ax8JDAjQFYRCfBhhwS99sgVkbZXzIvT
h5Xu7Qmi2Y3PuOBLO6tJ8rfUsXyc75xTrtmq+npL1jnPAE/GD1JFpaeMlfhj817SUiJB19s5sYjT
EmJs/pM541IuPzxax4VEIKfNBGkVT9P1MZijdPUtpErNFBPgm12GeuhlMVSB/+lUbNndsrXt1xpJ
j79UixLhOQcUngEx6y1Bt2b8S9tXttI0f8aaDjJq2bBpRsYFQFbZupx7Nl7p1xZTjXKDlr0jjVco
TXronvGv6UknW02JgB94RtEO6Lo4lAPACI3yq/Y03a+b44enSA9O6dFqDFCKjae4Th6414hKQ7Y7
GchwRr/cWaDJr85HfRXdY90NONSD5TkJLTNwWRSgunxk3IcCkOa0wcSFuKZf+v3EdOIVYKU6Yefx
uPQLMFAs58B/y0kLIr4r82LtXXo+Ec6rT5W0tLMHkhrHY1yhVWCGFDR9FhGr7VOFotSkzbu+FtW6
KIdoa8ogM6C79vQs4PRdc8F9khynS2Mh7uxxm0+Y56OHPhPKZDe6nzPJA3JqXMW2QRr5mj9QNobL
DrrhlnOcmiADitnJ+c+3KgLwg4CAcVDlGTvsT5ilbwRDt8TsIjMHsqjneinMiMEjEk9qwjFkk2Hv
wquZtv+fpfXxo6kqMUjeFrbGkWG/a+3tzPDBqBgM6s4hj7X90usXkC+07w+0oHUAmHM0O7oe/L2i
z1dY7UXhRl5O9kCqiNilEdGo7B+gplEHJpH6si3mQslsyjV+uTWR/yMsc+iVw9C3mTlY+Tlq0msI
WO0MxI5H4lYAzhIMDvNNRdEVIoLicwxdoGmnOdd+ZI062hcGA0p7dKLVjkPwQoEHPwMEWtIeDUYU
QgLPVSn54EO+SqAeuj9lHH3cMPQwyAdzlye5ku3a3WCxfMGWRW86KicOLobbOuxA3eYi2lpxwJrx
0m1sJJCebgOgJMyTgH6xcaIaQkarTRTMWNx0lguzXY43yOAAq9LsLEHDGlhjmHTyFRdnHgv4yUxz
x7Li5jJYli+yiHVucK7xnwXQF7ekRF4z5001ASambeM92URzh0VRvpTapeoemwAQCfyhbWeWKWEl
x1qwawiC+s733WOZgoZ12rhpUCj+UMpj+jqksHayzx9/GclTLtCv054/zBdZHOqxTWM+g9lDwnbT
ASlILsqvGAfhl0r4M0psAr7axelpSeE6dZ3fVHYSSmC1DLUE553cyz6qC/DPH3EV6eA32hdSbqUb
/YVwmHbA8+XJH1bw0RQNa3EsyjKLD43+26DvGgMf485sEvM1kNPXZFXRKq2wB2rTNKSOo7YiL4gK
5GTnl4QwkGUgFUAraqHEm8Xy2AW2S+WlDZsZxWvUdhSvDMkqBeS+/OrMiLcPlzsDjH7XCWmE2/aV
nJYB1mc4ed8EGPRbek4x+z6oXZExYceFrfevOKrO4p5/xaMyZcwEDQZGXOECln5a6RL7qBqxEGes
FkrBczX8P09ZLioCXoEEm35lH62UVhr2RnThUCNV1pxQ7yIAANugjBRk/FiT2FHyitKKifwRr8rq
DwtBjQbKvXSN4yRBSASvwvEGPlPwGC7fHmZ0UTBGDc1YI3qkmW3PA3dQhJwAJAEi/BaUlhhdl+44
m/xAemktcca5eEPbCcTUCC+9WDgk9xv5YNzuVFmZ+EL9S0Y07JOo+fe1J3xiqA3aBu1f5gQbTaR2
S6rUp+gp3w8ijXQxV8Kq0INlPilzDdIGoZsr10CFRW77uoigFlDeu9FneqOA8ZsxvBQ6YMvzn1qh
s8vE03wOfcO7+faapHaXn2c0wMbaSPhpgjJY9ybR9xJybxcbIEWmBkGYN8XOhNd0xqW7aRbj3bGS
k/ZmGVDNQaMfBV576eyloGEU2liv+iCnYoYM87EgW/Glh6llmISmauachrUFIrMB5GHOiMpf2qpY
KkyEYFnWAVSdMoH3QAzMpelNG0X2d4zVt3rGW4AOvN3DfiKCHNImDV0WOUppd0ePyqkfkgFGO6Xw
WbJiQZRRv6DYQL4FwcVcIFyUPM1XTlSPI7B2KwB1/wN24LDOmjEIlDHO+s2r/hfeF0fmwlh09sgZ
9CZj2rNpNVPjteTj+xDDFbnYjq/NHQO7Gd4xuzqUT6H77YRBLEfln6EpGizQp5iKf9+nlkWhEApL
8puzyjtjqgi7++flsvusYFR2pVlJNhIiklPY+DbDiMAglI9BOP35QmjRAJaYWWrnWBNIihWWvKJs
G90WmTS1dysymVAfkf5hViiAGAQIYpMyyHs7dbxSbfl3RhqnaZpDiORyGSl8pPgfYaJsZ1s8AOon
u4nD+GhOh1ImTDXcAJhLTRuHQAtgGbGPKdrjAO4ZX/WwS1Cve5ised09YoEwx1fkr8vbWLh6hoWd
L57fydlCZpBc3yBNMnk7DrhehH1iQ6WLOyba88ppQPSN2VDy4uNFl91OUgdGOFCtSsjCZzuHxB8M
2+LKTybCdsVFkF9ejvkIUFG1RHM0YkiqzJnu8Qd6o1KrR99/Lb7YJm3NRsSZMD0/JwF+O4iUgl1b
9Y/HBI2fFgAi5vyAZHBbgTi4oxTgCdaY+zztYd2Sm8D+waKlo4VepCBWEuRna9R4lYBPh8SKjfpq
8fQvTNSQoFWQ7AwwNTLotbgP6moq2eGL2iI+qGyV2COyapmw7hfjlyYjQJ0P2GWYYCDhk4d+lySp
VQqz0birNsXguUs2GpsscyniKHqGimSmAKr71w/ZPxdz4FS3ay+pU8HNZ1bCE6YBgRs9B+mhb86l
7bJ7gCEoGvbY1xbALKqowwRNgOu7LpFXOXojd33EfIZw0tToUZm/BO3Xa5sbdLxTdboA7RP3gxaZ
vSlGB0JmMKJ50yO6QzTittcOB60GEgVUL2TumNHOf3rAiVDtV7RbyOvVxIiRqiUoxoiVeSxlMJWQ
TvqYUtxsmQdRmP/2gqocuf1xDZzMINJY6dppkqH18QODtqGROboc6IaVAeR2PxXC/N8p1TgZ8lJW
vehe8agrQjheiYpmv106sNELhy1szjcHkmj+Nr4exAsPcHd9QT4Anx3dKMUK0C1YmJsLLr4/ZSSK
PlwxvUllXUVQeEVzuz9d7DdwVrontrGvLZw0XB6bso1HmllO2yRGsQ0NOvwwq85ayFbkCQHM8Sjz
VYAAL5tbrTqvw8LOyYAA8HxbwvUigqsiJN+XF2QN2bjxk5JL8lE3N3KSJjwpBreid8+dnCaoCxB5
ELK4ZCFtjzPZcssm3wp/PkWnHIXiPsqzAcm+ryR5sdRRerN3HMVBGVNwETOw6MnRZ0I1vZo7Bf87
CeV+QisWsLyePiywT8YlRtRIjD0hDtVAZuYbi2ughxMoGTVHzGtAMC10wyGgg/4GlxjH3kAYlpl3
v5oWXuZ50Glam8eK4l5bPnPLT1KzuJLysDxY5Qw44P14fu9d3FaBvAB7ZB+PMTz1SWFHFAEHoRiS
brLWLXmqrkvPb58xmOfeJ52wzGUmCdejtN8sooCrJfU74ZKWdguFU2jLX8tDhH1bmqydAiwq/7YS
MLXyJQUyw7N8lbr5Qb/gV/XVoN2EX4XepKLdC+MphHpD0n2Iuf6ExtAK6Kh49l9GgQfFpsmg/bkF
yAvUYVpejTzpFG0C7ci4/r67jMpXqtMjOB2Bs7l5UOgrw+H2t513abKx6zz2NC942nLX+wShBpsv
UpHL8EaPaXai32HCbutE/h3ylnj2gk8GBtdC7v1GGgY1ffw2H4mTl8LHU6GK/xXpNCyTnEkTaSKk
tAwmiK350ZQMG/+3saNpVjKgeWv3YhV9iHk4SdXwXj9urwZ3DgqknHqGcpCKRGB3o8Pgo+IMLm01
aCoRavnfLoaEi++MeiiRWqwTKiAla/q4YU258BFrsset9wwgma9x2JU7kXb9sQQkmF5pFGGKF+ys
ByR9NpeDDftbQXhKFtbKtCu1f9fy7PZwt6GEZcSgLWXk3YP/8BGDU6sDpolzX2SDlYrxyN9tBXeJ
hM2w/X/HbGNbxPCShF721M4ItHIyVu/I6864gn+cVQyQ3eOhm+KmQgHFwSZVHJcJUFEgB/BCZBch
N1dfISo3f61viLj4QVIHgvHuIhGkr2z1ltAHpB5OWWXmiaFSdWXygl/Ko6evVEh4MhszCJHTj3xn
EAwg0m7ADkoMj3u9qVjfV5e90H+oj2ekYI0kQEOqLNSkxFG2skb7wna/LISIbaxadblSXTdhar9R
VU4VQfT9JJJOxDYGgqmcMpf8bekIKP1dxaE/JW6aE5m9OPFvNlrKQCojqzxn7gEts7Y6Hx+OLf4e
KMKxGgYKg4Ph2r20HAOBIb1xFxiJwgY6382DlIzOrGC+C5zAs4cxIPfxr5x59x77RxXN9Xe8OhUp
PR7tl8HYFkaBtR//36151RXqXiSLf37Tgu1gRm4olBNKSK4IAVJuLyxlZSNBVl51H+Iv4tjn09Yp
UTJvHyHGjpr2Yb/vKcd4EfZ98O6/WMdZ52Ddyrs3NHtRIaux5WL2aoHyTb1mjAoiLkOup/3BBseQ
TwtwC9KfdiveiFkTmG82vQUlCvV282PySucFS8PfHGMfmiZg8rdXZYrsgYZMUHLjC+BGMCCDThRH
1AOJuk5sbmuxg93kmhkN2YYwdrMQQ0TQAkstzKoQYt4Vt92r3VL1uvU2Qsmg6sIePxts44AqK0nm
Mi8OfDrWDUpGaXhqBzvyKYGNs0CyW/1X98DkuOFEVN7Wrp/nZpxI22Yzztz+VTWKOAu42P7SRNRA
4GS26walEQn1gaQZ7V+MCqMKLQvEA6h84D2a5qxyvXRSajSMsOwNB+dOx5ZzpVYeIab5772EqUPJ
gAOMVsaP2ISv+57B19m+jpT8w8W405eC5iz8F8fGSz5PIYDlsgt6rLbNCsOGklmmL2JbjI5kSYD/
c8ZkYtOSY3Phx0e3TF6TTX56KHdLTSTEpL4Xxj96OUQvjgXHooyD/uobunN3FAa7tM2tWOStlNsZ
YCTcgNOdl38nrHuWJ2cNVZgG2ZJf7pPUNs4c3JrKqCT2wSGL+4Vb0kqfW/tD1r94i4rcMF3+RY3U
QoUDrI/ian2bLN2OWEIWVPCZkWnQEHkoAiydgXuI95XHkOC4xqWAWU5sZLC4nZuHhm3cnUWI45wF
4wE7kEv8OELUAuB4gjx84C/9PTsyIyzN9uGcem6aKOZgJ0bNcdBop7iQTZhFAc7FDtb8Kaprrqxx
XgUeinBtJfjbU0+dTAN9UuGX2hUp1r8x7ACcHA8688unAjK5X31OMDBlVlTUT7pOxy5n+Qd1Zcir
LGpv2Ys38D2t+Qyq3k14l7WSVPanG9GGBYMbCDM0R26LivVuDB/aLePQuhQ47WesYGWzukLCgz6d
UE84GCjXApCRVt38/U4/xtHjfaCfNqyFnEqHfxGYmCdkrsDxNa6U90Cvgx9J35GnNOD/u1Rme6DW
I9yzCdEE1csg5RsaNf1ShdXgwz32jxQoKB5ro5VzWLFjLB708EA70qNJr0qwFIjYVs2jTwwrNnkL
22jCl8xI9/66iMs/728qrfJRjNyY6kO2Yhyhu27xlJXN7S20d5Iy3MJXaAEnrX/zS1OcobqkYJvN
6ZzAS54YmFRpCJ5m65xnjSEMj/azCmmH7vR14pdEL3ZOpYpvIbOKde2g9g4Jk6RiLWnobAkzQygJ
N+nGZutd2zMKjHiHSCI576/T1nd6RMYvLmKiD9832WviHWs5D2hEmPmneV3c9Eq0qrfNUF+4CGkF
3KzMlqJuY01bxOvpv2Og8vkjdqymRFj9PTMBXi/7poA+yVHZCy9XQhuyxWK6gAC+qMKcR3zkxnK4
w46oMSkL701bgP2V43Cxv86DoBXNsYDQt/oDLWoYOXcC+oGRyRz46Ex8V2KrdLIRmdGflqX3jMfl
LUobI1Sfl+QkdZ/4vDSt5Acda86huwQEUpRZe3wzTGwLkVGsrCjbhPd+3eFpZmkkhz1eSxTiXF5h
VMcZMwdLDUFXyyoeqim1oRgoJqBiIdWcx1fIPyjj+kUTLYneTz8zgZE879e1M48BMGDGrV+AIIHz
BlvFy+YDLMK0JHmlHeqJ4NqSzFpucxoWo4jr3XbpoiRte6xPm43oUl1QcjG1Y+7TC9G5+vGBMzvv
Bvoys0j6SFMAJtjpsF9xzAKk0yK+TXGBTssx4/Hh+2KVaFaarQDZtwxc9HRU6ZQmCbKhP1aT3Mf6
1GSVRnvr98V8X9UGcBhw45dE7KA/K0TQGvU4Y49R8l70P7sf8UPgDhyxdnYEX0WgvXYXmJVcN6s3
W/uw4JYqh++pzPWLbAdm9sZjD2MZxZ7HB/U8g2bg746BuaujPEnfZK0+X+byqal1buU2yS/QQqBf
JOXhJYPVImi8wlLWqGlSE7QOM6bafsxg0QYfi6oDDvLmLXVjuybzUu3z9x1zTyy3ESnwQw9PNxzA
c1Ii6R9s9n/g42WOi7iKHfOXWDkaqrvWC9Fsg6/rh9UQ3J6J9sWDHUFzYXVorR1ztRjNV374cnWM
+3/SxZEUQx0yVGp35VkvYVQY+4auoPfaYn3CHgcbm0UBiXIiLIwdQ73ZRI36UNPpJBDdwU1Md3uR
qXIZK22NyzgoOBb+MMJLsSOxJldBKl8YbM8IcjvSiY3tA4Cppcdy6AL+YEdL/K/Ip+JunHQoTW31
qvvDWnl820lPfVnBORGJiVNdkH0vM/Nw6Q+/I55i1NRrSr8BGwLf+7xUGO6lmhuLFC2U1DfwIin9
pqtipkyG7dBJWq4xE1X/4jbglCFhi7KyfxY+YGnECvhzMr+iWEnaqJ2UtXJGP4YdXPROUF4zDdhh
DobmEGVK78FY/ELz5h/yWP0t0pIX+0s04xSqabvscZVgH9mIWLCI0va7sgpClDGrnwLOTvjt8z6v
5rA5u6ZlpYtcTvP/kOucqhaTzQ3c1q5D1Y9r3/MW3F3fMPYMaPD0ABDZrDFStp2zrd7zMFn3y1/Q
/dBtCZQkVYJFWXRMIFRG2UcTlmi7AcoDckoEzvoJ3a0sG8q6s88Ok4RtOvBQG3V3XcQkDg92WkjP
2sqBCwc4UoTf/KpmbKVQ1xeyTFfRZ7Mm1FhuUBaTjgO+C5kcV9Ld2zm1i02Iy0SQgXApbaRmgmfY
zCGrugxVQzrGLjhnlbuexCDnTjBHDZM3aDHER/1pvjRnnq6AMefvZ87mA8VSHqG9BjmF2y46+l43
kIKmJzzCM5bOtZlXbFU1ZOcjlog7ArB36d9dEhp5Qip65YDJ7gbJuLiAEkSvlqo62tnS3IcEo6pC
YRMeeuZTyyhuDl+qx1/uQ+3PaK1tZ7ahiz+UHk+u9XfCJf5t03FSU/9hp1ZvchwTouwSWwfcA2gi
7UTvUVwkug+ARd3tUS7r9yAZfB8FOVYEsHHnFwJnDAgptRv/4UJhF1rfg4MDw0Di02sLftNFa2DL
i3NJ7ev7vZntD5hL9B0Bj5ASCi9RJChX7O40126GkkyJgarh7NsGyooEbl/bSGde0XQwGaZ10hVa
ar82fVd9ONwVXDDv53IDT0xQHchJCfQoHJ6NzUAaDSZhvUoBgTi7aIfSwSI1PcRmqataq8CGrLRr
kTs+9LMze+AA0DBNe2hhZJ0+czwzZonNwWugab4c8/fHCkQ3dKo/FpVsgb+dwRuScAKmwjsbtfZT
Y0h+0bBrUuQoQTveFcb7yshzg4nqqj/q/WVQqn2p4cbPaTe5rozDQB8stoNZWga8mRNbeT+LJ+lQ
9QvKNsIkh/iF57azR2bHbU2XbNLqNPOXszvXx+gMWigS+OIky5wsXRuk4G+SYkpQFOmCoRJZzHr1
J6eapkUi+5vubOnKFbvihE2d484rBKvLzdeFMnpcfwMP8T8tRRmYXUIGAQ1TIDgc0Jo9A7ay8Rjz
DGDxhzzwH055pQyAGinj/osfniNSfWgpFhIreBf+lHSOm95NQ00f9ot7qFBz/PmwAmIIgs0AU5Kb
k8CvYg2yUn8c0muLXBN4H4Qyy2EQaHinOFKP9vGcl85wkb5xl2lIDO5yBobCDY5qPqAgzHbI7T/T
FaqwXktcqJOnS7orHr7PlPrYl7lmUKhfXE2QKQnBdYgQbpCve06Cg7p2mFAr4L4MClySYRdKIgM6
So05ulGN1pUNNQwNvjjAmZGY2K4cGxyQ+IfrERO3XZvorSeL+8uEFSoB5TJHtgpRfBItvE+tQN/Q
bLJNKFKLXP30FRbZWJjesk1HUFC9SPtEIsKrEJml5JlsH3doXOsSel9Z0j4fx5xCeZ0yic6v8X9w
53zVgcx4ebnk81LVFA/w/BYozTlSlMmBKhj0896GXAWVMBbz5JDSP+lofBItgAFJrg5xSTk+KOtN
RAvtcUBMfXMUjiFR+EPMHYKQiDV39/2fZQHbGLP+XXSDij++ljbgQipyG/gOlAYvjsaTV7EjTXiO
JgcjYrb+mMa0oAvxxeBNyZouNPU7AP/+J9LLevKHHziExrwNx6pfZaswcz9iMjVWRyh7iNbNSRS8
T71gJAQooR/ywjtYZiE8ja9vFhLFvg5+uyhwiu7/2pxLEaRSf3o+mpbX1PTMVYHud2ZDCGsr6bi+
EVlMFTxIaaxWv1Icro6OQXhhgSLtfXGZBYnN1/wti4iv+xVGKme36Jbu7WzdUVFDzV4dH0evcHdb
1pXbnJFfTCL2GkZBFMA5h93+09CpiwjKimxh85unyjH2YiO2zFRrT2g7TOvr1zLnH55hjfttEt3R
KsB9CZp0UCLGwwlkAamG4+gIWKi4ZY6SrMlhLrrp1vi8svrPbXZEwx2SFV/h50moVHTJPKiImB/8
2SXRBM3EDAjTWyAtrQJRJdczTNEmQyqd5UZy+arKzuslVcYHL1f7DDcfFAJYzkSaHB/jndAT1hHC
bxJ6wRLlwQGzpSdTwijSHZSvgEbE0AvmAAgvQUS/o2QFBdNl5W9K+WgLB0Y25fRmAmBSbGbUIHFK
avvEus0YACEZuLD4zE3Z7agj7O9xl15XqkXMBLoeA/yFgeiXJ4XKoA08A8i2e2oyvHMP/qpHRSdF
mO6Ly5fQTLopysOQcEVD6bmCgPeoXR08EbIregazy9dUixXEV4tKXxi34k0wxfAFVxZUW0BgKC/d
FEJ4aQUegVSEirCSVw1KSq9cITj0mpwxSYrhaTfgQ0+lHB2WuBZOPZrQXijIQYuChQKa6ov32put
mSBKkLEGJqEISZe5+52mID4R5SZSGx7vShSF9FAQYngHri7+YaussV6Ksa6LamzuMRl2UwrFaQnp
EpOyAXgRriWXdbVM+UgqD/QHy8MGflJ9NHp3pFv++VcXoi2qviDb3vv2kbtHXzwmaHVPI8zkG+t8
LMJIPgeSJp7PaeSkVUg3kSIO/VeJwheCHg/gNQ6cCJ1TdDzpTHKa1myMkXtsDdvqE9I8leJalcWN
OnkJVPcvzNoGqhUgIj8ZEBNx1+izhgDX2F/g5Y3q0eIn15+0ets/AsfaxT6IXaB3vIXec4DHcNwR
5akXlG4UB+u9kDn5Ip5kUrLEEvDrRnT+D6sa2ZeIV8FgMVv0J7TZphnEu96Lw2n7iEx1CryoS2F7
sLqAgsh5kLp5a5eOZV1QddNCMEXeTj/lCBQPiSVU2EWDpkvmJRIGSDQKJEN8AFlRhdQR8f+/TR7h
GAkl8+bTIbCDdPSNgwyc6FXTFE4KtQP0zYYezVKJmhDbXKXudOjNtkg0oCjLIt3ExdL+/ri/wjr0
RSeG9v3ajZPQMifUQZcU+vbvtKEH2CLyllueMTs22j30KS7UlNhHBV8b/XD7FTnhjK8t6AHNY/Tu
O5JpPzT7HjhTRPtGtzFf1Ob8Aepme3r6ScxDHgBRfVaxtEubs+d8l70akAMJcp+5FyUKfjdpVImg
xIaauO8qeHI1QFktcMNFJgbKaT2dzGFmjwju9HMq/yQ2f1zxxVKCEFo75xFu5Xz9FlK/v5v+/f34
vn/3IxU3SPcknVmxV8p0Sm7QvvHektyW/vb0eUvWy23hQ6KnHpb9VqZw4BmE0PluntGZ+kGdgxVK
IUHKStulionhM2TEiKZ7/Ei262HID4MSRhowb3Ggn56yoZR/WzkgFY5v5pq6b5MEC8XCHx3agZcZ
6mo8xcK2WYsgU4X/4JT4NsLYfcg8BpCO8UmkgXL++pOvgB4n8FWO2rY3fjjjHMZx0J5epzxoFtK6
AuTNv2UyGIoRAJvyS+TcX5LqTSlrzD9o35ungWhQaIvBu25DgjZUk77iA6aiIFvUzlSAK+KqPsfg
3xnb7ewoCUWj4MFMPKyveAcDOJyXDpY/upHIYbcz30/QYHHeX3ycAvACIBAthyrwiLvcVY2lpyzX
mvToYNNnpL7X1u+cOj5DfTBVWHlmeU1F/uEE4uSYUKEQQ0lrzNA+7IH5Y85AkcM2AbRrB8Jzlect
Pj891zShz9IGATcXgJgjrykvnVIgwCVrgOayXf56fvcwYWgNLrsERtyB2EMBOSUuKA+b8G8X7Ln2
H5A+16rh64mZSBe7ds5PjgmcYHi+ROjF3TmpuAT+IRSLQWgdewub2PjhgZbwv15We3EEkV6nhFkn
UPAvRgJYyQK/Y545XIhZAaMeAJAdSpBlZ1ofuc1mcZXBcQiU8MxCsvm/VpSpC6bW7N1Rwo31ZjDH
Xs1izVGGj0kZ7ZczWqop0Sq4t5XAIxaiyxCrdVIvA1TcaM+CEFxfkgIeO9pemxtHafx01xRq+4zV
2qM4WkGTEBD3HyqERCABwa17Ou1pm9cWMhvIBD3dk+RHqyNsSrvlZ8hDOCaMDb4lLJjE7Gmq6phh
0UTR86ZiwX7DDTtCuYui1OHP+lXB20IZNmnNyB3dlcrJotplSaPZpDP2Uj/pC4+IyXXUpltYF4ki
h3QXVl1Xvuf14weFdaSWTem5GgNnTKbql4aiDT/0BvYszxBoUazcpX7GGfATiUw7yS7WReXllH4d
qZ6W1FlW86ph2G47kcl7pdB2Sw3TbrCGE9H1Sd2F90sL1+dXn3DeVdFifiPjeDT3u+anT94kh5Om
k4Ei7BqhSunEMysPJvD6Uvhg4kWb1ehmkcUXjS1R15lC3Hhwx8NnjdVob5dDjBzZohsKOUgBHKsK
EJPjZ+E5SSqvnuuEK+D5fGvm0Hxnts6x396R+ZI7JNly+AacBx7IKdEK6lWovU+9aYGFFfSE+1lR
JF8O/fN+gK/9GxRU1c8eBFaH3oo+TdIiSN9xjw2UDBwTqvNpyJv1/6FbP3wWgtDw/N6jw7e94WUY
sy6lVj76SZ/UK1c+iVQ2wqPf/XsbufR6seRhCMCIv3tuZbAiPhBmAe2Lm0DsHCR6WzTTAAwPcNNd
vtidFRpbGOJeHMGuMNnHW3wjHMblFJgBt+wGnVOIx4rqFvNLQ2T3PGiMsuhMuli11mcRGIWR+tpM
q7k4hCEAAc/ljc7kKsguLsWWKTEBeWdWDiyR8tuV5RPiH7azK66YtNGtPHDChOaPm3g3fi9GP6ih
y6d3hFzMWqJ1yqOwEimPGOLEOP/o/CXnzPcb3jpkzM0CEzcL/SpnB4axp4Lg3ZVpdck8auNrkqSv
cbpIxASmvfd4zzToQmruEBaBKwue8eJRf/rE3PxGomY2BAq81s7PoBMQCX5hQC5RuThPfScKGHua
tM4FMOgaWiFIDCvRCdKFACewoDDKMkzx8hzIPUHGH/7WCEAovvKTzmeb5ai6XikEvTaHtCo6x5P1
/p6c2iRWybBT2OMAebs56cy72hMtMSOgh92MLp05720d6/9r2BkxSbBwlSFbRfN9eTqXFLUL5Wyn
bnyiLvogiZxtGrZVYJTz+mdxQFKwbAe0+zagtSdPynXo4P9kGENn8ZYX/YvFaePIP7VzXSMzKChA
8OgwH25dqMcgMMzZvuJoCNNyuhPYhDWLjNjtjo28KumYIkfq4r/27NpMSwqBCEIfWIzO0ixlC6sk
UN1q0dd3Hv06NN66qz1+XV9SSbyGFlK/t6WY7NSNmHJR34WY9Rk4UwgZXB/OSMAa7Due7go2siYy
tDk0Q1iq9nJXj0tVsMlTgo5ramCnSF3dfivY+lg2mKEefY1QvwWKa+oKVH4h0AIx2KohU40Drk/8
Fo3cJ86l/+PUTXyf0SobMUyN6zwM5//BrVHRZ1RgtJqLquiLCVyfmcmTB/aEbob6qGrlalMrkSFl
hY28FEFeoestoD/HQ4uGRJD0SnVseH+V74JnWSkuKjPiLOw4YTFkIkTuRDcNbTbg5kOOl62PHsfU
S8tBJAQ2191ln1jElPwEDKTAJvbpeSJi/iueZx6xTnPvf47Zzso50jnjsoX2czdOZuvDDA+Vto2O
GgorSq0kGXhKNNgE9rnbYFQciouIfu6VxGdJ67KY4eSJZ8jRkEmZDekBTo3oBLL33Fb8zYwsbAKb
B0pNFdSrVq7UaiQRUhhowfVRLmM3FX7cUPNeZ8CHQaj3DZ78Zgt8x4qtPYqMN8PY4yWi2MZIQHYa
in6aLKGGe8agedeRqr7JAv/OC/h1YM+nqaYwy9cW28FhuwuUlf2wDT/VAMjQFGJKplsy07Feev7B
qcwGp2c4srsoHDJI8ryc5yxOAhmxRrjkF3Ui2F1WVyD/fmukK7tmj0yJ7uUo3aC/CTl51iJFMrII
Svg+E8IGncJPZPkHTx8flUBQCVrG4jI20CfP8O+oJ/hsQqetCfs2IVjBXmdMxPHidAHFbTrXFfaV
/Vjo3TUsQl0Ye4mxtvThISzpJhEMlE5OadPVsOh5LYtj2+vG3Ca0CCZ8Rs+nWuJercB2rRyprACP
E8e60QbSZkBO2atvmmLJ3PjjWHxs+gpXj7qT8A7VBdDnrQ2PfUpbYR24Be3b7bHhGGp7VMUfbRY+
jOQbvoa8e4QqMe3PL+oVlklYlIGxrCyY8JVXP6jYymi2SsVEAgNmlai6cMbsa3dEB9ZOfnhiqhNf
rKiuXwGufERjLG3xJV/SH6JGxn+pxPsBa7agnnqpY6DLlP2SNAABwngNAjT4SjOMJKPfj7Tkd2c5
oxcNMqvFzoD8LnWuc/EBSI6DYzVFdZkU+FQVr5x0o4dR/QzSbN/9yaS48Nw9HIdYDOCvOTSgDPyn
2DivO7xtQ0BXMG5jEVpmhEDP1sPuNGavZQRfJPz+Grbyz9QZuCMa7pzrjYucFcr476cfaMHLw4tR
tXs5HDwt8pDxtZ/vKb5/8xX5L/YgcBb/lyAUxaeOQdsz0U1/7y86dYvwv/jkPrYIROfTzbzSvC5E
eEnhudXvsI6PsNb54kX/dJ8ccYUKrlOfmNZ9e7Xc4EbjVLJlKpgKioBcJE9gIK6P79LYcoRt0Ckz
oTN3YAuaLHaKfF2OLAsE/khfv5DSk4UnTe0XCjjTC3SrWf5gvdAUoxq4igFUao/xw0p2AhPIM84X
q6wiBDzPYEvVvgFhC0a/LF0VNSmr4Vfh4hBFX94f8N8ne/Wxn82RUFJJjw5pWRS5KhNlvbUSkkGm
oh7CeRLWQSmbJ7X8LVI7iWfmCbssLVPqkF1kDJR69e5tzXNQzAakPwOhQ5X+X+WoW+icHluAXdcO
dSqzreDpUsnBm7h1vzZ2EXCdU7bkFLQcbk5AM2thgPVK0uWf0hjvhaRvXWLhYfs142Z99bhukShN
ki6Ll5VIt9AGh6If5Fk/nKGJLpbB8EAb4LfelwVFaMw0fJmFkrJb6MOkHvPc/6lj1RBHqv0MFQ2W
Co8awLAIMGe1exqot/EH/yZH+/fZthkxIFtxQ+7hW43JHNGftCFcrbN9dRZJOTjsM+h4C9RF34VY
axU/DrYgG8uBgr3OVrWGins75IZvwzIioYpJAFQhIQciCWgQOgZjnFvxSo1pjJUsyANyhtyVrIDG
+lvD1en/JAVWuA8zEqjyvdxYknw/ADvljcOSf/WuBHC5DYwHEf60dyaE2V1S76RQJPx5AbnTw9CY
7riLsOhsmgFEEx/YSim4FBAldMAQkerwPlhe60Jk75SVbA+t36Kg7f00jhccMn4SLisrxrMNPtV7
EIbE9Z6FjGyIOK62iDexwgxmR9XNMwAK7gMloHjEd/YNPhf6tAhFdZoEMNb4TFbt8GUrxmnII6ue
ooYjiP1ifpNKB1IzJDzATVD7xEs73mr/pddn3Q0n5NK/nSYROHdSeuV/5RZdZhafWs2rfS8YfOdk
d5+4h862lFmLWNbaD6dDZb5UM1skg+yep96T9Yght50h0Xh+5yVNOI3OPC0AILe4d8e8BSlToSP9
LZ1DN7hJpACf4eVoSFolZ/H0PRjq6WOi4ul5vq30gQ/pKl3317awMZ6rr7Rw5N3qPxhrMpqCzbAY
W8rzrK8YXhxlcsBFuIVjD8WfY6uJx2s54kueEcyZo9xHnjD9Y3mfb5qtSqQIPE870wrjehV2Wgsw
82fJkOQ4SnVf8MX0l6CWMTGWxHTm5tU+qJImz52RMMp6r94KKRGfT/uvv/yUZL9K5YQqfGXIYBMU
44mGFs3SUu1sZ4ORquNqS9i/ReEDlZPkLHaFaELhuHLAlges0NoKvWIiTmlitV79FJG/W0iKzO4L
6J+sEpgg5kot5c4g+yfl96CkPs/t4QWO52iVFu54Ia3RAepq8kYFSJL3gtUoZFeNGs1/N6UGXOL0
RN+clK5igcZ300IxuNmVc9BtsdHcOmrylk/MimBfWK45Y9Xyu1Az8s+l1YXSjVcP0mty6vGqn5mj
RTyTyy3HeG4rk5AJ5YWhbn3OxgP4Dw5hEhz20XkbMk+gd9b4lQvTYo5pL6TpTFCQkvljiKE9b3zL
v4R9xAU/tPtgN0IWrVzvwi50OKXD7pejlpP3RquHeHtvNlgRedX+PUYRoQOGTD6oTXChGTtRhGr4
hhAYdQ59e1+YYrBuI11mWjALHxhOMCHmK883UGcMZBDKWUaSlmd40OcnBOdZyWhRXU2vK2KY9qVC
OtaIuKKzDhNPHZhbWSYvkdjpnTx8EgA1GJiAyNlqQx8N8KAyMOB3nrWZ3jdXYUDy/3iAvFGhQNEs
pxNubxCEBiZIlJSRUOCryl1cD5ssAmEA6Q8C3HAO8VqJGW1QlVLGeqBlEzExXO7F91BH2sMjwo0W
t5Z75935//uQG0MG3CqLgtsRvq12CAeI1GuqdKmRkUpFwXIDUzO37eBSThob9cu4CgoJE4qCIChs
m7xAGYh474GUJ2ezZH/fFJz7xUBos+AZZWHjPDJO8B9kiTdLcYbtRRylRX5rUxtlwohswDUeUyIj
GBQrxaRFUYVoaeCk67noyU+wnh26p84R/QrlmL19Iiri6RmcEjToz9NruZZrbadqYhsVvvQczuxX
hOsKOCghl5pcXZg+JvScA1ekxci5hvx9WXLWwN2z8NdBdRJWnjQrQ5JvK6Ke/ftdpjfxI929z5iv
jG+EOl5DDHHBJeB/W0SNqlKUd6l71i6VK0YVhJ9UvYRW2AUy7kHiuhq/EcRy/jxX16qfVJAXC0Fx
ldPODS15UpThqeM6nxiSmMa8wqkkIR7Rca4gRrM6mVimWlHBeh+wRzPqDGR/HHqEdWffcyrOtEVC
9IecIRN9PaJ7/x4MGApi1PQldHmBYWyLi9On4GU6y4N3UtN9kYjH7kuv574BcGOY+JjmqnYbmF8R
m5Ja4fgYiCC6RYxd/sqZrD+glm/BQeytqWf4I1STKFeTRvWEfiI37GsfZcxrmlvt81gyx2r5nWX6
cI6+9qObnRedI1yHCAsECaLm7jh1E1iqmL+NukukBUpRvqmOpeCjMwfbvFVRvavFl0lJnd2HUGBe
/Rz21l0biR1SFPVLxP0YWqKB4ZRQGZ4Iq/2ggkvi0lBXVR/3soHRjWS4Pw0iGD9ekPLKEvJFdHb8
XkLvd/1aciPRk36mfQsVaOGqmO35LUq6xW7o0126ZdngHyodyrmhUYWaGQA3tDnSouQHDIsRKf1e
uKSz4tXGu7XWLT2p7/ww3H8Ep9Z4WNReEN+Po/nMQpgLbe2MhDyXeSzOI2VKiMdOV3cnqoRf6dZ/
j/4pcat/J1URoNADhkm5lS8umiWzEscU1o0HT1b4rfEkyLfoDB9+tUJv6zwhmnMGqUifRomIo7IJ
sle7MHUwiglr0TiGNqZOvDyipGB/I4+/fsGresFiTXd5q8k9UNdkmP2e4qhbCiqYyAHsv2W9DE0p
y9oQEXG116Wp7qchGNIcESRxJHFl0Fvx3pBYX5ZLn6GpbwW9PHgqHSQz7apC0B/8qMvt2Y3Bf5wn
iPJuyh73NtHPaFw22JHMjVeT3Qo26It5P1JBcGS8//eIiPH5thtRQXEtfTP/7j5mEXId+cMJc2ER
CeRGb5Ci3v5I5caBtpcFD3tfb583mSOxLzQEpx+NBvt6xeOmCr2C5I41mHM2j/SjU/C+Phnn5SEm
HG7sfqSx61v8I9kNZai5NsA0lcBzmpS904DbVLSsYjxiI2abbkKYNd96FudbTKzzOB5Jf0I3IfJO
hHRs6gq83G85Tyv7qBkNPUqheQ9242I9A0eHxHf4LsCVtfLU4XJWKVxppJrSgWl1I8Vm2z/ybZzt
u2/xxwvhf/R187UdaWJdooGCQV7TcNKlnoRsw0FEi4vAoGFF6Mt1tK8M1oMZW/bjafuWhtw7UBSI
+A8U8hYUM3XKck92wh0lKbM0LrA6qWVhAz0bDzvwuMLSagEV+idlGSwdllW89a7ifr3jQgUEaoX1
zKywwO4M3Ug74quAo9BImP0D/2C00u8KdyYvyUIfIBPqDlc+GxI1LypO/eOPIjrAGjjluVAdS4GB
OJUnh9Efm+0AlxICoZZai3VDDHAtLZv+s6+CFm9cvkkIMdQ60GPq96GS7D0YOqpD/t0dpTGJuOY4
KkkNjXXs3HivULsudBNxEHr3Q75ir0fpht/i36XbJSXw4qM9o86ZQAHtFCWe34gM1xUP2Q7pKKRQ
RGQ7OWa68aHzFwxtweOIf3Yx2zTk/QelnicaeSF3aH7+Z5CA9FuXZdydKp/KKX0DT6i4r46NawZi
/iGUXRFHQ9sBLQ5A20qME/p2GwdajzC1TT64NQKIxuEUNTk706Qk08urbziiy9vapoheU+Oivn7O
yCDKTFQQZW2MAoCj7ONH278W6XYhbHcLhCN4bCQAP1emnHaaNKY/Nj7mRI+F7pmGW5lmj5fIUbfh
HcsaF1wv0GzfgKfQqfzscZiU6MVL1kmAXer+sn+uzqztXDradoB8qgDk+jeHMPnVL/WD/p2SNvoD
mcvIhKs0Dnr5I6p5gHtaXtWuacjZoV/mPOCz2rVsWn26T5PjDqbdFHhdkU7V4oaLUgujQ84+7Q+v
iPrlk2vyzfLIEj1G6fmz68tyvHi9VA8VQeHuO1OJjzqJMCuXIyiTJ03cVRpSpbMKSrsqxJ1DAM+P
jUPbNjlhbAYqJGdFTGKRjylpUcMsizsq15Fjztx++QqTGMXcOdpvowdDgVu9eRk4ujtqFob8yjzd
UfedvGhTlfOhIJG0eZGoCkNQI9gdKZyzOhLy0Scx5ZObTLMTqSmh1Q3i/4lrSVrtQ1FIT03DobPT
L3oVZXkw3M5llP12gucfnbtYNA2VqAS3FzpSc51mrYQG8OLteJnOP9Cg/l/R/1TLHBXEojrfaQ9B
7xucRKvrti5tnEAOjaXZ5KxHuvFJtdwYUIcnSL2mtbzdhKl2BQA2/zuYvSAt1IaCcq7S5B6slT+z
/KAFIjPitWAHSozxP3Fa2QIwY7rdv97MNDI7Dv9KtSbwVgEfTG3VkDfGo2sSaSa93zjR1oZatpiA
czzz62bD13nkYrtcCfwAsuotAvwri7X4tpyrrSKoWJD64ajREmKXvX3LrqDOSTMHGWAnaaVv0H/r
+OXU0C2q+Gw2NCX0Zl5O9eAhQnJcezav2XBe6X7A85vfX9pr8xyGn7n29UBx81J6fTS67Dys3AUL
BM/im5JBzrQQVuZLsExn7NV0RzgVKqUnCVpmjm4spUKSDxOIk0LY7a5ElGFa2h1VmLb4KzPakjQv
+aXJ9cJ6wxXsFdnhGz50INxy5UrcuiUCbtxE7+cg4/cav3lQj9a0+FZZsSBbdZvJ2xdk2VqHNt0V
Q3BWOzkOAST7XNyY1yvNNQ7vDu84DR+MAQTU9aYnbsYHgXaCh39TDihZOy5eDeVRh42l+Mr+gam+
vF0dU11WpHzHsLVL/aTFZDe8ifSOaxVV56m7U1jcsWVTPKxfLQu2yi7rIGly5Mjm8uDDwVHGLFyG
5HApPiuRvkvlC/r9nQaMxkNk17amY+Paab6DjNsidxW8Rz3t5CRfzG/EOVgM6iVN9UEDysnRaMJc
Xgb773MinHns87JmVcyH70AJH6jo12ZvAMANCa3t65n0VSjMHPqZtkMuG229VQAypWawbmygHWI/
aPTB1W1qvvhxKf351DqQuTURynS/4Qwv87+6/DasJYKdlhoh9RPktPTSQlgrRlVGrpLXMJ50BUVA
9gqzSKPPvHtaD8vik4DptDlbxwACqx8sk3siyfnnB9tJNvQz3psKPgL5bFbRQStxIsFutoaMD3Bj
N8JvHh5Dz/nIW0VrfI/A25j+hPkGY3Amd/WdPFaLOm63CWxN46iqQeh7mndF+RrBZA4SuKEAMPFs
l7MpcbkspyIuYA71jqP6rNZenkKakQ2GIHHE1X5rQxvwtIc2X5YtzcCJVf/CEyY7/h3AJBO0JUun
0uKwnBQ1WeEXrOTCxKKNkZj2hWwFuF/Jv/WBYoOllmJbEaRNG5Tofrd0OjlmI+kLPAHtOUpA1oyc
bS5Lxjepq3fvLv/1zMm2lSWFthelX8HgUzhdSIXdA3FULsJ8exWnCqow9uamXi03hjg5tZxyPx/Y
np25oZLIzCJeoWzo8cHkZIwFBqtE0H00DCNw8bXf/dTM+h7ZusexgGEVhU+0at+AoXn/bH60b6hI
qRZI9PSEfym9CrpY93k1Ab7Z53d1IQFwDOVtWv6n8prNVMqawBFIpmi9kZczq+PcmRkdGv/3TNBF
XVlybV0trZtTJ40zZVo54vFx8+1MyscNg1Ul7TZcfNp7VXE5QqrlbwQpQwRzyZlFBuHEYRKAxbCU
6szT9uuuqJw19mUzFgyyWkj6wEQqvW5A7RrINFaizbUGhMq7QJYx9n8m1NM4RBA5CRcM4ev5vp/4
A1bFNfEyppvaA2Tn7vT645S386KVGixtGdI5fh+FoQDBGqoaPcy9jIhB46WUe9TSf0C8EKexwl6C
f2ETzmAvHS2Ed5+Yj1BDG/UEUKR3XufN80IBd6g9hb7S+yjtTNvSQzh4A9epa3UR7sT7Dm2+S6Gc
Wxb05vHwvKgRorn225KrgwhbJBFLq1CyEdzzRxv5/6VeT5VPGKvLSq3Evl/QCscj4g/20tUdlIjw
98K4RUl+UoXzd64hv8DqepNNYQueab6mu15UYzEFNbSJKDS6+b8+XsSjIhX2pEBvrHpO4wSOSsa/
aFHO+2Gq6T73/3xDGPM0p5X58RO/fPGnvL51Ie88vnSTCjrZJ0R9wGT2xh+ybcix57YmWF42xz8i
hYjtBGFW7/KRdGxd5EQezUi7Uwd8VvpRYlqKSBfHebMwQGZlZyaptt1lBn976QtPYqgwEy/JboQs
rzuz017CvB3WVbpCSZTUa+LdZ2HKp1WGimzQb/RZ73tTf2Lb65UuSJpVDdmAqmxkUdtTus5okm/p
aYzpjZbV0gsffdFnOwiNin/Xg3cKOUgvcHP7KyXlw2GuXYt6M8Cv75ngeiP07zzqMPAcLBFIb3iE
EDWg6MbI2297upI/pELEKMYlQpMtmXCEsEFvgReIbwHZ8noxbW761dqptYDgzKtol0ISL6AgH6zq
s2fDKHBxh0ZEMypNndFjiTuruW1OhSb/MfgryP8fQikH+hQi/sK0adppiPyhJmlRzQQQNwz0ddOR
WyaaxQ5zw62y9RtZdBv7vQNjIaS/Sm1Z0k4oJdVyYBJldO5Y9jYPOW3vYBQ7YzOHKM+16RDc/uCn
BTdaXfF6cp//MbsZpjDOm2Cz1jB9IJGHod4tbE/srIfRUZrtVrBKo3NCkOUabTOVQG8dkPOo5RrR
yP+XEH7EuYDuXYgD207biiEHQznhpSJKGGMkdOZ2m/CideDdvs/TKVh7jSFXv+nVDpwJOwX4oitF
aSOuKeQUgmiXi7txM+h4LcT9R8uHfMvVOQwY0wKaCq6oyzZ5ZKknpq7PEhsO6OXsRQmX0EmkvheZ
8/frI+DgUD09a8CklhwQxqh2C87UeQxlpIkd7h6kQFDk8jGaasYHMgwG0bVp87586zCBhXJi3Ql8
qC3MIGjvU80pCg4N0usmyP1DZlBtHZGrzU5POddEDoKECHdzuebglYWBbC5WTkCPBk64sZtrwTkb
RCfkY4kgWXYv2WvDAIRzIZxLs9eD3X4dMwRsBhj1qlS5vwhx8OcMIDSFZZWNEQ7rLJ8Qt3sOuts8
l62oiwSUlqKB2MxNmS11/nDWbcU6jMD2jJzNTVO5lORrfaqyqtLBk1Rv0Z1S3BFvUP4sVNCv1t5X
0EB7zAmcpN3X1EX4ryjy7VonuaYcrDt5W6F5e+Ch5HTIbyIaEqLaeiauLP2p7295OEmccmKeQhYY
pBclEsZmJDrKzr7A06SRPR5CN7U3alqV7EQPBbkIukGpD43qvgHXelX9QZGGFLts7HDAWmM++RrX
LfO6WUJS9XRZh9MBxQKyD1gtrDU2gkKTfxkwL0NJFi4Acwyck8nnNeHZz7Y4kX3W/Ia5sr4y7N0q
kIyaU+t1ohS8BaROuqeRu0wPmiTEH8ZlSobUyAYyYYNFs4wZJMVTJNMJDtz7O7WVtFf2I5ylP08N
FtZ/272OGkcZ/c9SXG8Gi+433h2dLOFmV6nsx0GG3vGJPFeKWYU61nDXzG2I11siglAMZ5ZJ3Ou4
V3WUR5Nnp6lSN+SVWOz3QHZzijhQreR2XXzxGFMZrcl2/QHyZsEmS7PNqEfQxx/XIrRI1sMx7vyX
5Aox6UWeBEJaPGcH3HO90pxBZPwlKtvrBtCznpOJuUhIptqqMw99tsqjD/xoffmE1AYTjZ1+VT1c
jJQfujtQcD7mN3yX+tVM7YDMUmsfXLM07kR4mSjp+ugL0CUdJM/CVc+E9+yeSB+9gHxwpbSxedIL
eX/nL/Ly9f3nE13tvQgprOtnELG0drftOCvbZLJWZ4rmr0sL/ArjcyqlZD37KZ4bdurQxQgREHs3
ESUqpDR398209hGDTJ6Zk45/FUNB9PhFD8Ks4ZjIeokYWC94BBNhtgn9Yk5NXHEFtZqruYD6/uXD
7pMTLOlhsZY1mIX8qgin3rGpA46a+s6cOLZuUwY7DKXb17PYkm/+JtMyRPk0NkM2l9fZHovCexbA
NeMvlNZj/J4IOUIfSPRf9Hr4V9Wwxf8P4c9+P4c8sI7dl3+rITWRTSti2Zav1cSxeFFcU/d5P/EK
Qgk+8s4ob3gA3IqaU4gvmWgWpobsrMx7wpn5W+u982oQUwVoz1/G1BhWa7P0XiQmPmw/JYaQ0DUd
Dj3J9f0Tk696SILNFL0pv4eMfXexxF7zNYWSeYNxF2jK3bE8cho8U7awaaH0ChnVvtr5MOz01o7a
wVSiFj9wa2s7c9ltWniTHXP6q0zF0K2HQYPt/tDTQNV94uQwdCItHvbqq9RElytrmmw1GgGYlOfA
jYgwfxHqnrx6idEHxn8ecbgsjPDnxXuMF0CVqpdCvDNUCbFpATaVNVFBBCDh6cwF1MSW7G3WGH+l
BbbltBsWjsCPrSbu+4bwBWEX9/5hZ4ct7stI8KEG5HxAjcTnpe0NOsgiXby5OT8m7Y/UInzDDOLt
U5zGP0KRqYIePmn8RqIbEwmQVbLT1M86NmNZBn2pSz6uYo8+Go2bK+TbgTMvMqMO1uVS/rHrQ86W
J+UDYgGfH1AA14A2bkj3C+qNxpFfxtA0enBKjeKMQfcudDAiFjq5F7ZLtCFPIdnGefXXM6rp8jer
kC9eYwzQRXL2VkhLATpq9n5sqljFBi9GLz8CmfSdTtsUNtVa43RVfjB0hnTvwQe1Sy1iN2/51hM9
cRO911iK1+uk1W2UvK47kPe4RrRWt6yMsX5JGWJ0XBwpmKPyW/cTxABZHFQ2ktX2qzogc+MKpJwL
PTOWq9n0GRf7xBPwXA5lVxpFQibYau1gQHJL6Kb1kx4E78eXEMW1VJTCwTFRX+kuqc0z0mXU7QZq
JRgXxAsH9o2umltgW3YVIILAR2Opgglkn2RzxgJeFKLMoPDczWslq7KapeFDRkCi8zzX6uBjvuOh
hfALXS5unUrwsTSS5qrjjqzhrDQ3byFU9kVIUQ0ldOnOU3jA2gla71skSsHaIl28Hv6zp7BjkhAd
8pXOc5VP8UaMFyXWoIHc6iCgxW5cwemSt/ggi5XXXSpCjKSvI2Kbs+56/ZUBp75hVSKwKPYKL6Fo
1z/6yYWCFeHXZacl99NDo4GxBTp2OfjgBIIm/gJ4IZtMaYjN8QtlH9i3Ydy4pEp4Vbcl+l7/YXG6
s3pNjvwtlOIi9vRoxavbJygyzPNArcycuKPk5QK9yNhfdyBlmd+Qf5wBiizzDfrjBRT+of89WulJ
GLRyV1EoFM4MnK/UlP81m5vpxyZ9sG/oLb0ByeQ5yhF82JZcHcdm8dU1vf51apYeiK2SoT4pxDuQ
61wJW262YWwEutGUY0KhOwoxMUAW9gx2qVuSX4j4VM7AKMNbXDLa8SPLRcJ7GEbDrXocfG5JVqlu
4CRw36W1SucA5Fzxk1EfotqX3ycamUbmiwvp+xhWTId6erRMEeW+KEeWqXAc4LZ7aflET0jZCVPQ
+r9d4gQh/DX8IdCluq4dTAWjn61rEPGcVfTh6yz91WWAL9NcwdAnmZfOFmnGcIFOkg2qGiSoraGX
g2MkTHIm5WPMFxzQPyttucYgngSyJRVK9Qags6bZfInhAD36v6RRDsTHDWLp1uHmh/LyrOBd3CGw
9oClm85oj1tuXT54murd30aHQB0zOMyIOhfJVqaSClW8vOi+jauEgO/N81MaK3G8zbdq4RunW5nl
ruws/OjERHlsRiYOXGItspwDPzork6juAhPiEbe3BAQh9RO3QV8gzKNy1Yg3c+Jbtzcl9mYvAppa
orU+NfC5klAGvuo1ogePzf0McNZT/ZH8nntIxIehRdZHmiRckqTXdNyt4jp3dkXH0Msgop26P4aw
cuLk7ONaYacvsI9EzBfkTWg4H83QyaOVgRo9YJFy5cPZk3GTMYDG2msuKhHn7//e/v0fhO93mACC
lI8/TcNieq8+KT7fhPpnYvgpDNlvxGQeVV7UTc6gIVX3gB0AhRXHWrJCrNU/ebSayOM3Y4XMgJEB
rp2kfz6DYFR2nYOTGWzE1uVh1hT79/MHoUy0mBwnDQh9nEK8g1XHZbqihm2PQ4Rf1FWEFFxbaSOc
RAZeGZRIvCOa1lHOGTGUw3tZqtHkHSIxYHqoas/0/gCyLpRqsm2/PU/105Vci+QXPBou4T83KTli
SrAcIhpgCLJlRqoJlvyZ89cBwHSScZUujxkcP46l466WwLF33N7gAACqPFTvZW91ECW/MlSKQGxw
O2kFQtiUWKkq+ioxf15b9unSUY2S0qviqeFLnrHhEZLt2nqG3miSLZROPZPHG/rJXXnFam1Ow+ir
iXt85YVemPFOy8rj40jmrEhUMop14/5W1NPAf+OHf7PI/Z9iKJFWA7OkQ+vFSktAPPS1t8y4hLcf
ze0WVN7QAxY3QCa62YD6Qpjw7PPOUQp3bQO5TnitEgy9MBGH+2bkAOH3Gbq421FcB28vrX9Nvb/r
NyH14gh3xNnipPOzyOsbvv/lzala7IevhYYkFdz6p4QQ7px5GJTvlaI36QQZzv33F2MLIpSPAyyT
G0YQ6zx/xqLMU2OqJP3z5DSGy+06xCH/cO6zIZc+jkmMvHk8M7D9OZCNCkUa71q9KAOqI/twkqyv
f6IbnAPpkemsUOKy3vDBTPk9cy6Q9BDmMAaDVIJiL61Rtks+sFkqUVG+0sHdL7TXmqqvGJ6wd9bF
cTp+QEPFH1nrJUag1oc7UDTZUikz/vaOq+g44G04KSccTtqrD6DyV/etXsid4SOELI9c+5HO9Ldl
jW0dgKR+iDP482cG7DWnNxTiPJVToBheJ/xMJ0L5VIadPQRAd00LTTo664AM1aR0779jAbrPgjOV
vmfBaVSdNGcArnB3wiNN/wS02lopmGOy57uCwYTB/pGhFlVl0t0VLlEqf7z9dHYjFpUZWu09qeH0
GLzegaMn1FRDIJ8Hxnz/3cLM5MrLGeieiKXhZOR09WPZbj4XV6Y32rnbdwEmCLRf68goz9/+6n3s
9EqiqhcctS1vPL5cIM0R6lqmTbK2+pQdoPVFUC287o9/0k5hSWH4FR87wqxmpYpimkItft6esve7
NPa07UWgPY6vonsR5gqrBd2058pLIHYy6VVh1aU8DVlIWMuW4VUChs1aA1DuLJ+g8l9ErrzMMwt3
1JORrSggmD9iyzfzi5SGK09LXAPJX5aaO3ib9qP/6173dwDIiNUl+NSsUIqbOjU6GW+ncMera4NE
qKQpuvx4NwhCOBNJIHUCzlEhLjRdBtFpJvP0jCjwjLuyHNMQiuJHo0OMY5zGwuciGjkYePNa9W8m
j5Cd2VF8/n51raaoVqQ4jMqym4i/V0mjtaS4t5D352zkThfJCzmfFbeL5U7UJ/8xNEqo3l2c40nG
uJ3R3wbFEffwOoOSjTrtzYJJuPCi/YDv8mQ/JydCwvIVpOY+7dPGPQszZYHwsTJgfKPH/YD3dZGP
E7PbFB5VoR+e7M0zSUVMihCCjyjY4gHxZCH7eJVkla3iMtCHtU0fEmPBIINhjygJTIgyxsMos8am
699FwDw3foHEB3ufnQOMRDdCpme8/Wt41S3mXjxJSg4ayiteBd78oitVNj67guwHlzzjjlFvvbVD
iNIiu8Kv6WTsN4A/6mnLEyFlWAQb8b8dEd958IDUR5bN47iirteEHf9f9oH0UdSxDMFLz1LrxyNb
VyFZY2XZc4bHxVCWBHNXnuK15d+AS4zQGMVneQrPblyiXJcvufev+t04FfJe2+ZKJJ20nhNvk7lX
2OQgASNz9YLRV2TGmvN+0HP2rRYnCaaQH7QoFWdomj3sFR2gP/5jeASZEoFapww3/nnhFZ/INzDv
5vl/YCl7c4fDAi6nIoHCT/CkN/oZoYIFKsQ/tdvDLb8IKWBpqRgOo2ID2TCTd4apNuu7FEqYaqTi
ywKd+ZJ5EhQb0j2dfoJ3wiI+MRaNDuzX6wswTbLztnGeg5EWIEmqrva8+iYYKM4X01kxNZvOHKr9
27id7nn1X5xS1gX/mCXlS/R1gGdAXbPMkBC5WfLcFRhbAP483gtTjrEHJpChDSTELLdi7/TJJi2T
XKIJDboYw8KhqwOTpri7s98kPcEsJrC8YHBCVVlHoLJiIYEceOZl6WOWha9eQqM12v6BwSfpHGdY
MzwNTlnN7BFBvYBp5cenChRDqBi9i9wwjECajhATvROpC/gyzFx4q1MsIs+N6rQftVKRe6x+Kycp
I2WtKF5+VHtLOrRZrIbNmcmY+REYQAPbCmt2t9GSgzXPErVa8vZhHN1daKkwgt+yy9CLmSK0RQRj
4tfRg5Rg0Pa3IUNU/MAl/X8igUuEnNJhaQf0EBsQ9jCQ7hpBHEHeV5OvIoWxXYsqym86P9iuSREe
Bvnxms2KPRqcUSH+wewE2u0vb9GaUVmBlVg3qqo2p0DY0x9jgAG+JFG0VIXdQha+s0pPv5mIMlNl
U9N4JZElnbByi0s63y2SGUU6HSMpU1aV9CcieNc1GVkYLKnZfXtBT1r8fxUz7b7v2A0iK4VCf2Ol
/e7jLl3gdcETbMJfW4yN4EJv6qv5GfpmsGsiNj//7G+Vf1KlYDdRa8EQ3tZHbuvIdauNuenin4z0
z7IbORryI9MxBef1Ho2Ztgdw5MykdPy/+uL9AbXd7bFfc7IznCNLTvBvVKdYN5Wnh1AtW8G+uRE8
bHG60O/oNy2glLo2LxYVAbt245Na2K/bJ2Kx8yMJDCFuafnRrtcH8sshMVa8/4wDmJUo7Uwc0B6C
sgD5Kix9/VJz5pGzTnenV5Qybkj/qqDqclLrV8kQ8BZfvEudHpwlKjGQQyx6TQzE6SLGiNMsEtSo
/LydJsaqvWrNNTulenz6BT8GYt2yy1qR9zZAuV2wSN69Xcb8O7ovlN5NNGSJl+XDoXMiwaybbwU7
dcXYnhi7TKXpVdPTsNZu/lYkT1WWdxC8eXZzsAyr5hRgBTxJVKtg4CrfB2Eb68+ls/q9Gm29hM8h
70Vi8WlwhzjC+4LR5WzrZIyHP7I7Xeu1GN789Kk8bOCEOMvXrDw8kvnG0hwoh3Z0xKDeHwiFb/Ik
lMuxH6FTYkSaJv33Kl/nPZ8KQtEG0o9it9GDq2U6WyyyJDAD0EEgVoWKZwlWn2O05A1k01/C8Oz0
x3BFaS/8XuceGNutTmO19EKMubiZJwjZLJtyfUrLg+fHh5rq4wU1D+QbkVzT8sjgwSH2I6ezts4j
kVPUlxJmUHCfnagzPq6eETbShv7rDP2BI7x6V0VD4FTNXbjmat4d4vAbm3NFUKQ1dpgLjNyJYbI2
knUpP32xxHpa9DLRDilMvapLRgNv/DWKkRTEU1usgg/CQTRZyjSBK3x1PHL6gGFKQlHfzxC3zdGL
f95PPJGwQITUVH5JaR8gtVZT8NL6XjZnRU9CTxwpqclBlfhx+Jaj++mXFZjTv4YGtriLPOmTk84o
w9qi+5TMTfW2TldCIZTjknqD/taHyg5BWyhR5Te4NczsA4IqzH/c2pt8lSFfpX+8OXw1YEHGEP8/
ucH4mdgPnz4u0+k1jd5ZeTuxo5FKLaGfkaOgrQ9urfYXcKgfBS/iG7cNugAofHCzj8ThFDkGhsWI
vzzRAepZnljp6wh43Rc61G15sRHwKHlmxPh/Ho4BSUWdL01sG7qWjwbrZghq3fHfyUgVcZkAZlpk
iG/y8eRXvloipYUGRaDE86SPk5doExg8SNvYf8qGftPRaLgKi7swtvyyZYrZrUIPWsW7l7RDIIg7
zJeikQ8dGjErgsWf2ARKfX4SXr6+VOocf9Kt4IUSGx6uMO1yqmSvDC+a+Ff0AcZOhYHC3Qu+Fe1C
jraiNr4sVaPr16ltL5jdNogeqaE9pGT16gtkl2ERsd4o0GmOzWzdr4BfndIiQe5tQCEa4GQJG1t/
iTBtnfWVi3bzz1fhWRESHVXC0H9uvwUCruTg1RDtRyAkKvZ8rsZmdJLxr8iIJIewWNwtk5K3VIm1
9lsPKTnD8axmw+5YJriTXdPWNx6TG+xYoQTvXjCdI84i/RAABviUYThSeyGx3S0XP0sctoFzHdj4
viplMzcEUmdGl39132BBt/PW4ebpp8axs8NnY5XP3G5atG/ZFwr5cNl4rjuVj4ZtXeEx3wwuHFIe
n8Jbo+XoEy4useyJlWJSJwbkDD8eGspU7mXrC4QEojyhO38mTvU3gT5vR+CFOT4kZHkh1EwgcvQ5
UoD8JRNHAB63KY1TzAIBuUtYC104imilbvSUBmXdFF4SuXmB1eia/SjKWcLT+YLGgrNQOMhk6deP
zsROqSgb8z5BPl6bddqOtSxWjB7ANLOnamTRjkW8Ui4yyYuzxJ30O+FozJY1oo8OZM23PWQehEiw
L1VsrjakiqHv+gBL5AYt12Xs1RSyOInbCTG1mYDKtpG/nl0pZ1Nz9LP27IPytnuQeAsy1V2uvbnU
NzyE+fVbOLIjGLEk6L/Jq7YyfFubFk9XqtiSlvB6FKQPrmdus5kI4fDVqPHXh0KyLFvULE3qnkCj
Ed1613PA6kQpRX88lITGWjEZk9ud6w8t2eiH6oTg9KRqW5DXC9r2MuA5V8nqVZjV5LBT+JSSJ+wu
fyretsTWZyAeNui+7LbdGCAn9zLM5mS96WfCSnfOEbK5abbezUiVqGQM2UBi7nTg4IjnXh5H4Aah
pPNnHA4dgQgLQ3rUVqdIfG4VeDfIz79y4AQsFxS7gVPSrw7yIuiQMDmEFfW8eA6sYbBbezA0/iX6
9k4FkKR9CG3GppRtsy+9eqG7MCd2M588ccYhMcZDDLLaBjrFXdies5Tp6F/Rdhe7DTy6Dfr9DxsS
UN9HjuZb7+Krl8XnLSnMQxiCbaVF9nx2ShkKauOMNj24M6/EH2Ky1Y84vpKou2uh9kuD3xgmEelZ
VpLUSs0vulUtZdOkbsFF8cBavrocp6xKmPnXrDurlH+Bgvk/AIt05FWhzoW5nkFyX2ypCOGZcQJp
TaAWf3COZtxBQ6CGQAG6VxTpIljohOLHG+j4dxmN5C7fEgJmirzGal4vaXTsFlD7LQDPoqs2xSJT
UmJSc7gH/O02CIpE5y71NfYMmzMZ7O92agCKeHSbdvAH2yjEfgSB7E6wFxXVXBBiioj7q24i58+B
+9HRkGnGofazZN3q8ewleXKQ6TT1smDlHCuIf7HwHneZdxmUFeDdIPe8iqABewQePNpaX9l3hGyN
xwVfCZcEsOyCLkOLK7uWx0OVY3/FOabItxpOUlp1sKjl1WrDDBKMMImliNkXugGNm5/eaCegPGrV
TDm8gSzFyOnVqrqwjtPuEWdM1KsEAEmumQemDn5Ajrij/33fDE48dPCpqliMdfuXWNTuWvFlQEKz
f18+fssgSIP+rFcf7mUOn9RqtkwAAHyhNJCN4pzh732nHj2MCBjLicmnGQeEtnuSNpiLc/jqFZEB
XbizNPaAUWmDpZsTZNcmOWlH/nWr862w8qYJ3jDFmlgMaovRF1CMOte4L3PnJwh2eMnjI0QVl7Ev
u6Q3lXRSdYOYwAEytqfP+H7D02jg/0PhxqkWwl9wUqbBFvGnjpdZcoA/ynLnJ4aouSlO/Wy0yWoL
ektMIFJhKcnk0F1HtewdwZ9pifaHMrURKtVdzQovmBfu58FIyFd5WuxknXUjpaXArcIgj7zxOPz8
6b1qemyEqW5Iw5ZC62DjcneaLJ60aZLnv5NJ2aG89I0TPD3+CdtUC8GZ2wbtIzAAMWmS0UWEeSls
1dQJ/8oepKNOhUZpRiUDAWdgv+5P8Iz7IpIT+TsmEn1f3iSLnQMnF2RyHJkwgXBofPLWufZYVV2r
6rhHy8qBEv7BUvWbioqhLLqEu1wox31vXf7FBXDt7cfZqdUsr+1xE4aTzDG+4WkXs1XzybR3jeXT
uZFq3t3/ZDwF1bYilRq44qjVZZnOi71E+R37nU/VHxF9LydNIVpMdxOTnYvW4VSoWTMkbWQdT9cI
C3x1reLXG/Cy1CzvYOpbARpZuzjoVTBSNuCJD6a+GP06ZCtJfhZpo+WGLhz4IlXCRU9RleYk7VW3
2Cj4mcrYjAeNcVAx2UHeULbCey8yoeX8cOzYZ9PtlUrqhDka+UtQguH5r3oZ2tPwl/RNdyH5dsxA
uce7i4wrDyBsWN5KmOQCzRU0bHn4N1FSmUuY354WGAP3AlR9MAhYjTFhG46Ii0SYgxk7GFO8Friv
fzXv0A1YKuMRa++IIjzscv7La9j2mZBrt6LsFfMGKScBwdDcecZns9iY8OIGche/NyD6wUwJGii2
APG689gFWO+DDz8/gfbegDExY8NfXxR7E7rSJrBIjbuNzU2Q9N9vXeh8N9q6UAaNZNZWgqBaXtCE
2HEhsy0D7wGpQYmh3ec3ZRSTD40k5JTwDJiENX5cJGuqTICjzSogigJ8SUyLQ4WrCvg6ygNY8V05
TZ0CT3aKb1xeGUC2QzLmWHW/ZV8XsXB2Qc1Y+HuZOJc8Q5yEHa4y6Pv40yC6cRfmiQqnX6kRe7fv
c7UFDqlA++ilNyFpsyMt49MIUsrkVxWuBmoVVSPOouGVVxZpb5zUx8aLKVcZZyXZRKZn9ThFJI3F
VSuO+vBdYuVcsKlhkQakPDoKwK0VJZwjorqZ1hMJe+xNou8+6VnuZ5GGrpX05OH6B3Thl6EhC1gV
027dw1n1T6T+uSE0kZmerbG+HtyWXU5dVXYoa2YuCbEE5/xs8AxuvB3h6S/UsNC4ICHgXC4yi+U3
LJRhew6BrOd1B8AEdnoYrtTjSf2D6RRrnZjXGMDPh2c1gI8n/Bgyc1X8IwMoa0dCtEI/bNUecyUO
gtT0YsFF2yLVKietarCxK+QX4h+bMBPV3PdZRx2w/4lT4HmM6PwarMEPdZZkQSty7aHYVuMQBc9X
rJDIu1e+JZ3TwHHi8W5YxNhF1lEDbAID5ybSK8/bq9x+Go7Y1fpngvtM23BXKYlqVTz3H6N2wbtm
qLJ2L2tjg72i2vvN7viL+HqXlGBa/xWzkp+NR5ivALccUCsJbFP24iI0aZJvD5t+xJbEzmbo7ChV
BNrEhecpMZ4sJdfEB2NXy2UwzI0ii6Sh/R7hza5fb3Xvd5XiisgAnq3bSi1a8Bu6fbO3/MDfvvNn
QwmAxcmQ+zZ1Xnwwgah6ag0PeUXlDinynnnAVVqmkGlJ54nExZ093O8oH423VqeMRmPg+3xQkg+W
WXJyS0diXVXitpEFF5e0dYQD6AVvwNtLogFoUrembJLPvogiv3KDJyjkK5/ZRmHGCHNrJSrYSNaM
wcqh3wAjXEdB1b38867zN6zkvvgZorTJ/sKYJqCtELu+8d2hC5CzkpVqzUhoiLuz6o/cwPV95LQx
78l4BOShUzZFRB3MMmfy795LMPZ1sP4skwpavzcgWEHHGFjnxAkwirlQMHAGoVw/JNcXPGi/oy5B
XHf/o9HxFuLw12b8Bc/UW0Jj38VpKsYnHG3lAuZxW+NZqajDT5Jc/7P1drXAoRGV/4GxUysItRhN
9bzowTpoqVDtkPqsncxN2bQdQNUsmhdATlUMwBvEWm9XMrcv8h7GdhtUHnxJ1PEhHhY8X+HLHOHh
wAuyiHA0ky3Qc6tzqL97WuzeFMAZo+rJCP2zxiM8EiFfm9M1WNOwzqdZVgJdS2VJGopcDVue/J/G
HJ/5YXW+eb03+ngo+rg2/d3TuRsbUWQJ0IMOyerwOUMSFlTnAUKM18KJdsApfHWIkLkvjSLhZbA4
cBEMRWKBeI1EdOflvYCJCvPdy6o+Jtjiyl2YDGU0kis1dm5l/lq8olJO3QlV1r39GfkIV3PKkF5/
Ovt46ObIqiALoqF8DT2Rg+KdBPAtuAfcOgaXURe7JUURr26IvuDlZXKLXLx9qIw6JQGxpQ6h/gwv
u2wNDi/blOgQ/U0PnX2qJ8glAfD4N9DOWXMo2xUjBFPWpqJuKKaXVRxPzcBwM5s57PIrq6+/2E8D
8DOfMiB+7qd17CscM8z79+ZYbzmpaLJhG5+98hfbhqwIJE5wW2X4B7vwsp2bQ3oQOW5DLQYhFGBh
zo2X/Q2gzu4dd9EtZDvyCBfVXiKdTBZA8BZi7/Y1HGTES3ubDIjRCFAhf3FzQGX3RZp7IFxMPtyp
XGdOJbv8FQa1wROLXwFcmAs3fGT3Ust8sKoPreFt0jrJmgBoJjETxynDG/A/3P+cXnD7ODcK+SFF
hhiImxsWFciptFPetIiV8l3p/6D+tlcWq+J3T1NHWUfyY4Fv33WbuohfbeWffR+82Rcf5Vro9oSS
+LsavFutVcRJS6H62nvgtQIo7zrqLKTKdf4GMkHZzA8AqALe8jZnbI9Gp3UsRi6KgInfa5ryxNib
Uw2Xox2a1PscPAXrD4sbsomJiAB9gsUnRxhOBFqYECluC23+WCeZj9t5xAywUzeGBDWNmc3aTe9M
1SqZmzKOeJZqgFRVjUmMChCBkHNkhVyNi6jJkIE30Tk8nF73AuYLplmfj3hv8doGhH8BtqOciEKW
fOqgNHZz3lNvVuavt6G7nVdBsEc66MyHVacs0HXdMvr1f3NRkuh+KMenK4iC2LGxwD5X1cWo5vlf
C/KLqszt4L+91NsjB+rs8Me0nLN9/Gy6vUTVULnh+YWHD2mVdKbwLo4NGs9XDGwOqat8Bgj2bsep
e6NuicManYO8yesv9X9DuzbG5/x0dyGGnd6byvH2hfM1ZODfyWZrVQgA+esem8iQqGAqNMk6Hm/4
WeSSHbdP8K6mtOLbmBu9i1Rv8sGlRx+TrU3grz+c9S8ZBBXFtlZdXznbx0i0zMfs1daNoQFavp5a
oDcG2fQunr6+5MqcVPIalDjJl00WH63aXxuhaNxu0mMRcmwlV2l1BEEuXcB+70jZHd1YhUxnZ5fY
lS9cAw9+SLDX/jF6r2xK5/RMWxmldapQShrC5ctGiWfrDIAz8a6dn3xBZHhX/IYLSDh9fWa8HabR
aRbDWcw7WPGVsRY9+lzs+6cPjC1RCRMc0tp7/+tExR2Od+KaCfd24OICV55iqhsUIj36d5O+8ICA
JfW0Y8sstPo1DzX3Q8zuCaPG7HyhVm05Blk/epwgveLciSYyDFNuDaEycIjy5/OHI5pFYn1jzZrE
N1FFeFos0M7e5CZQXQcfYIV6X4Rw+CzPrUGLJquSGSnflqGIFsBRrRVbrwTw9GSGVyFwHrpSZF/d
I0+FlQPqWGFPXvZUaDs21UAF1Lt7TQOuglBHolevb5PsN04Q7rZdRFLIVZt8JPQs4lS2ueV+cSby
y8fcvtaU1QDaWKroZzhddqRx4m1dTGslodz90ezxomIuRhhCcJANPuv9pTgM30T6z+z8pnZ7XyuQ
Ci6oB7r0S2PHGt8jw+K/RNdICzMGTJIHsgSV/OwqD2cXQKjPVQqZ/cXzzlJjEIUbaOD9USDpT93P
uOLzkZxIqhczWx7rMO53Cg1iYUxslbdI5H5q/zL+OWpqcSTtQThswI0ZyQrRSuKeVAN8NPxqHofa
XU2u9hXUziFvUiVtwuOmDLhxv5lo0rWO92n7Lw+gzufCMjOe4CoDvRepDuQu1/kB1TTvhFdj9eX0
aDkq/STNdxWTwerHd9Iy6312npaaCFg4z61wrqD8byRu47t6NooWQUoTToB6zq7yBcM9fpzGNQsR
wq441q1oihZ25k4UfHGp8WpTUC6E7whpcWTmYG3SeEDkeLyKPTvY7J4r+PFrNBefjRUUmyv4CbPy
t0NKbU27ey+NLGrmYuf6pR3mUlLuYUTvaXMCO010l2m2L3E6KwiP2k0SFuG4Zi9PMBr9jzhdFKbO
vJY4JaqmUFntTcmblFGmST0LJslDQ8AwEGyy+tKGFO0zjIGFBHfAKh25WmyOhnjFXCUF39l3mf/J
1Mq/nmA5hRXYZhh5eXlYKB1vs37mgfF5MS+3T4qu1LfKz1VutBlcvyDKxtUrhMMhbBVODJhO25dP
Uyf3v9SA6fcqX8RwVtgyyjETAaqY6g/BQzO4UBX+NRCIkJvEyZWOh6zDzf1deHkjXwGpj0bfgqHu
kjeD2f7450zgSeSbMTSS2bgGOvjqAB2ES1Hat0H9/FflbWrvv0c6mDJZ5XtzQi/pEwfkjvxLOS/J
YLFxxzv3S7CKFBtPZuUy1E7p02hcnjiGcLKR1cJlxtfu0bANzQUeZ8mUo7Iod74VGy64Vj+mWVyZ
Y6TmuY1qDVen0/6n95ONx1mp7LYSXKNJBi19hBKwTZJI50f+sjNHExl1iDv/F2CKqp8ReeDTjYnA
2nljXX2uDNXgPNoh0+h/8E67RYAciLMXi1R7HC5ci0JvB3swrPJiHKsKwdGEB8vsxq0eupLxCGk/
sTEkvxoy+oah9Gn1/FS3g8SVqHZq7ksavWLBnFUH28f7Dlz1cUTXcf2X0ioS3uEVkMDBOdEyV/gw
TLymYt6SePd60WlzfHomIaDJGHqVRpWWw4RhAuBI1+mcHmXJiRy64I9eNHFN2TSzQgPTgy8dTeEy
00H1AtgvwKXWLu+ERwH/4ioU2UiOCIXk6K4OKvi0lSlGl4/nm4DgBTBdhBf1RQCklzYil3T1/bZA
Uv3pae8hIVibvilEU4zekzK3e6MeNgfKzVUemvVO10xqTxEpE5Q+np3PsaD706bDyTjYC5Q2OinU
gyIccNbR1LzqM/4vGm+8YLvgVkx9b85Sjyynbz5Jv6Doi5xuyU9892b4wnY4wY1Xu/zqtcZLZAXz
aw5JCzSkP5GH/jLG7AYaBntVhhXQbnu5P7t+Dw+GWwTxrnR7S5cQkWth1NxX6T1bWOsNcVvLuzPz
zRG36pI76h7CLg9sYay8sYEMqVvw8G8dFqAp4CERPbIcxiniEFjuMRdtrTqT4gUxfD7hqXriOacm
9OaA83e9qhIBl1o02879Pe+SrVCNHmavLLP+HqTEMSGhoNXfGFm1YzlgnTHZ1JzSm2H6Oty6CV88
uVE/1AbECspFtbQzMW3qGTPOHaEzcyn5qxhtSI12k4GIM1NPE8mNN2lG7qM9/lZQipFiPuYsc94p
NuLJscmoIm/2w6bbc0msWDpGlA4IDWHOQNe3+uDuUFXGJL3DUz64QNyXOmCvWY8NB6/Sazp/PwL3
HA9udqDBBcGSBmqEEi44waDxPLNEkQUMwBkjWQoeumn1t4qSp2afFQdSRdWuWJwu+qMwJNmBCEyc
dFg0xKM0srbcNfpp155iUhz+8XAJOeb9tMZkdKQHi5P/IJAkyZ+WFJUbiG9m2pIf4/IEQkZ/U7tx
tyfCcnYYQ59YExr4IO3lpT2XNa2wBv358DYrUrTU6rqCzAz4LeqBbuN0H+ll5DoS9qiTJeXiwcrn
ZnM7Vsi+KJsl4Teq/YvOcrF4ihiVPnM7SOlX48EUC9Qj6HqAjmDl4LdGNSvGpFe2aNL57bccLlpx
f8E6w3wlrQkIdCdoGgoxPKJXGkAjbxgqUzUD3WIIerv/bigf9eylm8Gt57aKxpAvBsX71mHPIEJ7
KyoAQE9qOLPQwlD06l+9s8qT2Po1ajTL90VfW4+dKiHzg6/5oP5xHhMfrzjcdyyDlTZIbT5bS2Rh
OJLvgbPhWBJCukBOst0lbcELueTMB8YlnITuc4UfrDf/f7mtd9mkclrwPpcp5SJbpdHNBBuFRhDn
fPNtveo4AYWI/8NLi0IOjSfXGjh2ZgwJ2U2G/7NKxrUpmS8gDus40qBlNUITo7+/61ayhY2z3COG
ULw0Vha3XT29Cy9d0OlHwb2833LH0PBFKglRC8VQjt26fyHGKHUm0cGRGQFCKEON2fCKGWFH1dRc
RIMKOsPjAeutj/qq9pQ699fpthrKru04tmCBiHm+UQ1hZq1akeea2QB6XWEOCaY59RGLDEOl4UWh
uiUToHaMOX7ths82i6jRDEsBxtfLOtxUX+VKCQleYYB9DQd/yl2m+fb7bqLy0TO11aKSPwvRygjE
XZ91+IUA8EThFH3rQ0BaJ0EMqu+Xk9cy87zpilSrb3/vXNOXkeFck4KzrTGRv96SM7lRMiL2M8Z9
zWSUwEqj51ScJNeyg0hIqZ5xOz5EQLIua+0tVSGTlhJIkYlmzCQ9x1UbpWcy0zVcgVVIl/eird4u
yEGdWzTm7gYQIhB4ygkFKd3Ya0TNrMLwNkB3gzCIKXEMutxzBMy7mwk4u/ePPpyVvOjVik4HsNp/
mDaDQwoWCJQfwSUeBPLv1HKFJOcaMQAfT2rkleVhU8MA7eHPMYOEbiraG+8n0URXqUv3VfCCN8Rj
MrnENl4xv8kk+1HkgAI4MxJkJek+ufeBfAZa5OZQfN0eu8Ovn1krin6nPacNc1fezXfOwFDACNJ/
7XOqdrg+572CDVyP3OUz8sHgS5n+pe13JDg+i7HFkeEbxliChtMWbLZXiJ6nyUadfRcfmGQDg2v2
vHlYUOJBnSbUqSLA1Ve2eO9SLh+TBhNEiljSQt4Y0htMkI0O1Tnpazv8uUrabrvrH5YmJC26SO/u
3ZCOKwP3+QUYvjVS1j5rFFWejqPCeCWh9ouG5ZowVwxxD0IfF/qHtJeWR1a618pKKs1onIyeQmjj
Vk0cTjK4SlcP8D+W5gdINSXNTAr6GDXIYy99d+y0oK5R+0lhWrVypOSu1Hz/Tee5jOg7QHQB1w5h
YqFcbIyw1LLZAMftemX1RTMDKydZqLRmcDKWErXS0mZ95lMYUJUkiCzB5dJinmbcKV2X1uF1iHoB
pC3hiAUBOP9GkPbf7REmxDEp8eFIH2pzPVP47njgU/GsPzKmP+nXuHD7awPsMfEoZ816tv/AvUrx
eMbc88Zs/ySkMjX5QPh9cVJxGyE7TygkE5LisAYUiKrdY4xn5NcrC69U7I/JstdTh8z7GvVnT1AI
E27tc6WcmR1Umk/ZkzCcJKm3JqSn+hjeevRUGXnzQLCt5aKDEzzmR3zBATdoegC5dcxeX7df8uey
igcqRdT/5GBDyA+t6Uk3h4JlFbUYsRZYKZrT9EfL7P6qWtmyjX+46BW4C2RpPJo1hWF8Ctf+bNUn
Cu9ffGsOyuS/g/zJGpI3OMsgg4sNQ66zLKnjGDcqfgIe2RbcDR1lSUSp8Ff2+L5F43hyBsi6z4n3
RcyX+HEDQVTp9D4hPJO1xObflwl1NChcGXVjhqvJLpfMZoARmjaYdbfNlPDw/v5s4tj4YPvWix8M
+v9N1tEwABrA+jujBYym5H87KG4VVI/DrJ2mIB4/UyKuDv1rX5MKGmi4lo+t15jqkexfjtkDyX59
IsxpB+X3SFVT1SOdC2SEr7f7//7V79WAk/6f8jT06uFNgFFHu2rdWOaLdoS5tUfgamaWcGmYwsjQ
my0xJrCoHshRj4UxaQG52jvkM0+yUbaaMrvYsDsn+PSiQuHNlK/RbVKjNMrCAUyzZzPWBnku563y
/PpNF4IfnO4YVBNUebeTCbXYu28zntt9QzzsEtUFDXYmi/++PfKA1D7Kv0z7YzzhDUHD/romxv2A
xlfjdbv6i95yA33IhzWXVpbCENYFSW+wAUP/BxiEU2zm0LqMDT6xrc6cT2whHX/nXow36Y3J0Fza
MN/rITrCXt0ab0l40op7Ylq/K7cvLiwgA8FhsyUM3X/aOwKf0hNcvRPWH3hD/LCN+1L2CPqsCx9a
/0glrKyKdsSuYR89OFY/EisnwpfIHHdQRLqU9XhgR5e2mv5TIbrJJro9Hn3jIpaVe4J2SLbCdo0T
zbd7KVtazB2eiZACNM2ps8xrXXwsgcrGvvJ4GwbBSXbLtumaD22nk1f3XpNFPEX965HSZePWlucB
Adgb3BtXXLgu4xci+ZfKagacCm3pY8q3cKSw/GwvPhib+w7Re5m0oFSv1b1yaYxMKg0eaBX3GGu7
9Fgqg+dmmU8DVhuzNTH5nfhyQ/2+iEpb54ZXq4TwSH3hj65ghrdZI36vfcJHumAjD8giUC3FXF0J
y7TCYsCEWLKn1abgRECa42IJUC5jEn09VttPKBcm9DnrS2BeCbDol+P2iaNAlW9wjyR/BJrj0VG0
RRY9mcXeHkEC/mReodWYAyUY1RBhxelKvP9nAoP4sPdwVrWaULh4cvGqPnxiFkcB4CUJlZuuBe+A
BiVL9x/+pgnTNibf+CHZ0XQ6ipvvdMrpUGZjXO2WMtV24CTlU76OzqNSNK1xWkyand/CzhycuxNL
LWbcujdafL0lyp5rbTxsOQDlY2GkLGcmhDi/4vtbhX8Q0EqjpD3wI0mc36t1WBRUe/74/tiiiZhE
cksaYuQlAzPVnK4HKRFCPZiUsjD3R7A9XYoGLdEL/xPP/lGurFJe91H2zh3RZaKfCJMkl3U1JR6n
bO0/4rU3h7mF04vUCN/bY+IJ0KGqJnIVSj5QmUw5VyDHGUcnPia19t7so+xI0UbaIi4eTUtSrAuJ
qzZQY3uw4cnILQ5a5o0q3Jtg7zOXuUcrmcABcR3txLu77o8ENVcJSNcbFbpQnKJcSNUIvfsAoEg4
llcFmnotKECFRFAU99QUhQ4WZoZED9jPFlfghTqdGQpZUG7c0JBd48u4R56rS9oninGBxyOJSwAy
qE+7NiDvS9zFvZLGUel1Wfu4Xw4D2GJuy5P882si4sh2NbqN/W2TpYM06rSwvzPadmU1l7G+crQl
qm4QfK2PN/Nq3uyZEE/oNfGIjgFP2HqvwKVnKFPmJT2nsvN66QFBnqTFoLgL/zsEqqke1hyfVYGw
fl05cKJPG846qj/Gig57MCYIOG2e6eF672uPNpAZJv+BsEkyHiWeWQ+gba37DHhrd3/WW9fN0C3T
sITFq83hTtd+xec5X7H4HMnWq5bgiqIVZtKFuHeFbi7yuuecoThwTij+cUyZMaizJGvb9wWQowDp
rb97i5YZyBZr5e0ZT0FiEnwtaa4YMTV0pJDO9BEgwyG2xn21j/UGfhjwEyqjC/lMZBHHOaL8kNYH
sjK/WtJQXf6BJBfHbqRryuj+rozawfuCjQKBajT3PxNXckmXCvmXbK2SNfzeTHr9C7U/ooTHyEvQ
zL+iVWHsNJwlQmLvijMiU5HMD09WqqLOL6H/DwcDy+5OkJ5NbQZJOkAkpB+vJKg4hU3zQs1Y8cgr
HDLicAj/f5bm/BCeDhWzLNEk7RCh2BXlbPbhBsLdP/CDEYj96iepjy6upiPpjsJf/eGibfNBHT2s
tDit4SWXZ/Hx7PTvqxNgCLlarMzA0lMnHAk38DmWJycUppHyNFXrWyT2AH3EDAEuV1GSTBphFCY4
NZBit1bnPukUjhU7gI0b7NmKiJeS1ejr6H8S0aBwOUvfP2yqZDV+O1sCBjurt3ICbpQXf6quIgTV
80h2NpSEG3PfOUEsDJxcRyqjtwoHlYVer3xIF6hO6v66So0sHPAq4gWG6TbQkDa7OUz+33eg4S2f
/GGhVZKmDnZPt/48V4eysrS85DVukfP8My8/quRMH8QrS7Dc+px9C/mG1fwRoHd7jzVkpUm9pspg
46SBhqw5X2KSFHtIQPmB4hXgsJA+mkfrA7m3E5whJYBfje0owKGVYRCyR3V1ADClNL3B76klFCev
o2VeKqYQdF5zONL2+cx4UeqJveK6cDrWCYnyWklCUre0Vd+D6E5x1nDYomkR2tuxrEZYsJbCD2T9
0ceo3AmQeQO4ktdVNbbqk3MGr2tZhjNMjE0CS6PJsDXlGqVGcucCIJ1NeEvzd24YLdOOiTauBnsv
u1BB1+Yq8tsGYwGBFUDAuNukdr2gIU7RhZuWvjKoZ7Rhb938YUT2PGfRkmFBUOXYl3UdLCn1wbh6
+/K+tgXZj6GdYbmdjGUrtfgN+kqxckRKa69f9v78fGrSBgHnRxgz/FmNjzrTerCfjAaR3oB0Ie1Z
ph5Y0EJu+xkNMxkJloDYPBqGCLWnLazdjyXWrYtj2FqwBofAlq960ZJ0gWk9mRbgrNOmK0OXjCqR
nkLS0ki78K0t+FHo+WZvZZYzr3+HC0e3gyMJLpK8qy8yMVZNEZdUeucPyUfN8qBxySMcHAAiMBWt
IxbEXggdEA7PMJKAxim2eWEp4WcRDDHT2isKKW7EJ0AsOB9YqP8pIipiqa6u8RWBTTsrvEVcnEha
58sFS7iQ9o2/P/O4RTYb0dCfBxHBYGajzPWVj9GivUkDeAgzk5xYNLKvJtDtE7kch52h54EQBrzH
FoOYq8HGf3AQzscNnfvGVjfjV5Zbtyh8t0nM5WTnmhhnlesrLGFxbzCXeqZomD9KD8yvnSc4PkmR
HHdw0HVRNf7zH1f/HRJhEquUOaybQ5gyZ38sIALVE6+qgNFHwiQk7BP3nk+rn0gkIelQzVMj0TZi
vscCrlty7RGk84uZGAb4GpEquDXwCNhxtKV0dAoo9y/kbJgF7HKZdFfIcOsxF/RwGg5i9+0Rsl1u
J8b6fjhiI4YHPVnoU84I1ArmezBF07ZlFTMTWkIo5t+JnVmrK+l1JL/2auH1HB8GQ6EkqtO2A4dJ
fQ6U0mQrFq2v4UEUiOt9b2hRHRzvtNxHslg7Y9FiZgLGPS+URG947bGZ2SoPsP6mRGpBcbGyN60m
ja5xcGztoW8y8Lajvw8fVfOTmUcZ+a05sE+eBBTseuhfuZQFKMg4ewrW2HqFacoQNskSHAPxHp7S
xCXetlknf4V9SGaWumCu2xX1GWcHmke+yyQQ3WWdkiP8GPbyDoz5BXSSHlgT7eiWYR8m/cq0GdOd
5t15P+cDMkFLvHZMSc5V9fvUM0cPRb6FDRJj2IWQD7KmPeIQRI0k87tfBhWtVGsHNQqffvl8xDgZ
pwn6YSNZIhgXCVV93LoG9NPfOSVepq5tMeoNgUHOU8RHyHpjLL3gz/U2/jNWXXAxuKIyAU1yLaso
HOnIYZBhB3dKiSP6DB+sAMhSgDT9Yn5RUsaPmDj3/xsPWHlbWR72zDJnZMDrGW26WRyFaTim4+O7
PnzlWA+zDEbQ6uKmHPhFY8zY7odYEiR/tdvKON2+SJz2WzBP6gPv77aY5CDKaQH5aoH3EMfRQ+QW
sWUj2+jmigVhY0fhtKKvcWAzcOdt2bqWJ2mX2dgcN9rrzFhgNyT5YrGgfWtdsU2oBFnOOGebQyW+
i3cA0W1wqP1maP56Ons8NOo3mNh8xu8HqNkBJ6/3ef+aMuyB9B7DYL+eFdXpgp6HZ7p732l/tPfL
e6H4f20ZhWxowrdgKgVNg4qwNNvKREZNA26PtYFx8Yfx5RXbaLkytVeaEr2N+UlGSdshMSlhwT1s
9iSeJFDG7O4+G526rWV1SsTrV3uWc/C7e40TyJqXyxO5LzqnH/O5rjaAjjyUwTZmBUek3ckg622r
a43sNrY40c9pY0V6youVGDWZNkPKMSi8oPZ18e+PRaMZZZSpSaJBK2ouGrxyXqU4Wr/MJXnv+s94
YlyzaIrE8exNPf6G5uPRb5OwUF/5Ct9QKlZ0v5xrcBGnSChPrlseZsshcbY+9myIolLUDkPB2BmO
nkbQeXbMY1eN3uHL0q9vtsV+IyaYAsofgS1EuV5CcmuGmwDkrqB6ysY84jSCEK/Xqn20AgTrxd7b
Egs/9W94VAVvgwOZV0j9JwVRro4qJ09YcYmWM1dBrrc+5H2B1h/UwZunR7bwuasCAHPUvwFMXG6M
gbH/lBF+v+/W2ZsXK3BCDK99SJALhFLaD3nYwVdvaNZzuJfjECWq9Qxe+bml/0G3DijLrl14HsJV
AG0fT6p2uuDP8ODESccM26KWIBIlsz2SDPeH80cjdUetU+cfIkYw0fkk9eq7Y3AJLY6Opkym6GCn
Xoxf+eLzAxNJGGRx+9eonyOdTuudfmVQi1SHGva6AlAmOa3gMyvQSw6hql32YvxZTZm9u5c8buRa
FnDZDE1FZGc4owiFuKf+Xcf91DOqg9s5Ga4jrYaPjodjLLHJfpnoWgQ5prO/FnndLjt3cyJcc8GW
TSKXLShdQa0UC+EFd6EI46dqnV0GQpdJD2dukj1Mucr8gmFJV/lGwGLkHN73i14oqqOIo69GMi3d
hrsFPC1ynggHw0KKUwP9UVfPQ5u2+zCbTpiAp4EOSg241+NqfiaNPbj/8dsQwGCekTI1LhWG492c
DCQbzkWL9tSgJixgibVvOWM1r/cG6pGxel1NC61p2GP2ILRnU9kX3EX89kND0Juc+P28g0Gbkais
NYaQoTBRC/XMV446k9QWlkzY/emlXK1KjSlb9ZncMeGvG392et3l/tY9fNestK1hAmR71wOf99tf
/wF6g+CtNiSXnvzgbFhLzRXWbzNJdyPDF0v2SJL/AN0zZ6ehwfSKQgEgGwhSDJhaS78yjLXCGmVs
KYmx6YxjaujfQsLZ039TVTORGCMroqcykNL3vvlsBQSgZO3j78SZkHf2Yb46HdGfUFkXbt5I7Cpc
bfMnRTy8wFjJ19/kh8V0x7175aih6NdAk1UVP+DsPiLQO7oikJdiR3mUkGV1MC2qCjQ4fV30HQ02
a3txunqLa7ENiiDRieaTi7yuJ7D+skafuycB4lqy7MG6rmgN/Zr/4AHWkCAVYLTLiW5TJE7LU1xZ
15GZeoYPqL1z5RiT5bsSS9OeUmclf5FHqRE+rpG28q/CD1Jv/VHgfAZqEMz98DKt3Ia2vtAsmmNi
uHYs8tbEivA0EycG1NWr8FvMymOe81g1nBt/ae98d9S+M6tm08weQgJPYqURthnsW37ILXJCipgp
byVrftYp4S8lkhnHpUTs1XK0+6IueTrvDK96yZguokhxIZgfM2/YOdXgUJg/UaGacIZhGw4AXMqS
x1FVjP8f1RuzTyrsO6tT7FwLUHiTSDnpi9S53IYpKES0lIDYC78shW/DO6W++Bk85BzZc1DLq7X4
ca8YwiP53ugI8+Lo+55jBccV2EHA52RTffJPml5le9LfqVph+1OLxCGuFkKFBda5f/BYX0EGmhHX
OrqyvQ/2o2Rp0FwhY7d5g3W+3D8cZ5DLj2Jjc6pAf0o4w8+vI/00xk/pLNme5623TbnDFoYn8L8R
eEXwf1lfZCWBSuDxe+A4F4BKUexdUWMqtrtKpQ7QnqbgR9RK2o5VE7GskbcCqqOUIDz+mJBnKjpv
NNu+efYuo6Gmm8IRFWr2tM7xfOKhhptCwzjN24Qfq0HhMn4TcZc/VouNUg6JkcaqM5vuix+A9rYn
1sZ/7lyCRHlhqqXca2fOHaOLddoGY+j6C95ubgOkv61uaJm1fYF0rmAz9406dVJvHeevYRXWrfOM
f/arTlxOCaOtsmbiboLBSsmadyA3Xa1DoSGmWIls3hoRVda8N36Q8kWKO1F11uUV0ycI3jdpfeqY
5+/wn+LBludOppbFcPhbWzBgTc/ZBsNan319M4w8qtUTVb/7l+HCGr5BcuAVU2v2yZvTdZmOdMZt
POVE5eDg8ar9oDWeZAowGe3bqFq08kPHr49UGnsqZ24B8EA6fnpWaW3aCyJmz3VbXOxo11oBUL6k
dHAGpqoqlob4qfbP7LIp1AbeEJweDFnPRvtyyD795hoxJ0W26AnIw8pvgyE09fmNH8VBz3iEiFOe
JVw0R6QyPc9fusY/eJWo76ZbsbubI4aC25qpZQvzg4xj+tHRxS3OAe4kMWowmqvw2z8rjoxgehJG
7ZxrAGcm7d9KDn0mx4FzSLO5UZlqYoRdKn4Ni/2qnIrPB640sRfxFOc2VjpYKMO15jWT7BpE/onb
QGEV05F1g/wVTo/DtcRAFD+YUN7hQpuvjLs/84DDlhv6LvhZMgfBpUGBWicJh5fOPA23PIgvk3es
nqKJ2QNF/chTVgauxDGdJv1a9ck5WsTwLMvN7Ax427Ofb4WW5ytEMdAu+4RE3GVrPxD621p+SZco
lKL58kpsmMO7IUHGVTiF02sRot6CCPbOKkGUMADS2ZC5jluIHUxA09cptPORHSg3eeDL8J9G8lhS
UTtd4/870SloTfHkofcQG1EYDJxVlWOF4njA7U7x6itcpRJYVcIDyoXDMjYOX24qUgp58w42AiWH
mqHfNR3f7fL7LQtmd2o5lXwEIAYnSTffbuY5ES4PB3RzhtoI6tz6HoR8DPcS1zAkjeSCS9mYOO11
dXFkbDlXiKDIOAuA7n0mb4cd0yizUp+tp4ietpzxfblQ6udAUt3jh7TgdfChe6L/2+rCHL1wugIK
LOfUjZ9MYVYgEkCkeLZ3nPrGnXqIpZkOdeviAqy3h2T7lLTVDG4BpHCyWMdrDzhJt/ACYIDDZkCm
E9jXA+M0c63uUrGEPphrNN3rSBiXgtJYQ5JerV3//AOaAq0cDFDSiSCVMfiiDcpbTVFD6JJt+/qm
Ng/nyqmAT70r1wXD2ObYHWJLtP9YNFkL0dFX4ytwy9fVqgKRnQtI1nEuLpU2wdV8Mgw7m6eQ6Mhk
6gDFWSk7iOsQ1EWvaRLD/j9bcOYq0LrHZHjUpsNvGSZFp8XnacCi/mzvywqOHIBg262XeG545lk+
X0qwHuAe4j5ARa5+FpeJDOt/tSdZfI1WkLgHLWWJp9htxMZsvHLqzSEvIDk+0ZxLBfIt25lO3k8N
iVoJZ4UteR45BA/iVhuMcn4s8kORqdgUB8ge90FnvoILqjcq1pJ1fyPFHvBGPfHPRi/0DfhY7f8R
r7tiTSJO3foYadFJ2PNBN6+9zdAhF24B1dlZiDyou76bTexNR6O7udBptEeGZS5jTuJmqDsSrixw
yYfEl5PcXf89WKpXkZxTZv2kk4ggA6fkKfuh/9P5KcK0eSVj6wCVD88yT0IADS23XbRnWhHaG192
bl/siFbH6NJruBXhT01uCpll8JvAwN+NvrWc7T4hQFSUivNMURfi7O0039mQV1BzGB6Hp8hwVqh9
R1lsD/IOfFD6LUioWgfftDthMiJLMJe3mRm6d6lOZZv4OJ1g6owpwKq0e2ADbdwHTkyXb7ZSXYrN
30YBM/RPj9m1v27aU6mIAr4X2WwOr36FKXl4F5ECcMxLpIjnLNwrM6gayOyvVcxeDOcPqRVkeZxE
klpYrtlp9uNRyPSsYvZDOCCYX0tplWDqjDcmspZLI2KLCX5aii7AQx3FT6pOWiRSHpgO5sGAqfI5
KgcN4IPDS9V2BsGDjwiOgcy/3Kb1at/sF9QTFF+HCA+cwKxSUj/vIOH0GLB98LAAJFNjMDB/oz6a
7uZLAYLO7TE1rMjxIaiYx1b8VhS6UpZKQHIf9RUQdv+usf2rGScnp3QxJqPcfJz6HhfZ5zc88HI6
cj+Mw9GcxAhi65JGT3JPCdF8bkkFj4+xgjB4lt6+xtZ4xoJIftcsUBCA9Lvt+SDA/z7Grjk8OfXd
Kqp2n5vngpeAwJ7wpOjuxSdEoPUdRkDwBtqnlNi8eBYDIWZo66sQ5GOFNnrRHv/pEEnYDqUedES5
TS2K+rX3CeZr3nGD0HsHNWgx14q18//zKnsh87LdRvSH2CSNjixETBGNHR/jERsMNxK01/RIGZm7
TRV3v00FBpcnIRgUgcz9z63Sgp5r1icTqa3giF4deEJrIqbicxHKoA3CXZfIGVLfPedUcyQ2x3WG
SPSoedRmNMr80CL614puAB5yJWoDzg40WesefQSDKIUmFVcUoHNp2NB9vRf6LOa4dx6GuODh6JQK
9G5yG5VqOXY/ygogLZSNOzpeKEuFEYaFdWonukIzz9xmk7T0TpypzNMpwIji9Udh3NYtCACCHCL/
kxBsPLJRaNuQ8beBGITFCf4YnQjlsmRMdeuZUVtU02L20ASoYkwYzYG0BE3pC1c+p31ING80ksHl
cf3oF3PUXvdw4JWDrrLSrcDizgIGNaVzxSTyMMQvm2BIAdOLZxI5/h9FWFMKqzSsb8J68HDaBROo
vRpNzh6VyeXVdNCJFAMU8ZDy8ZAfud45HjpjguPUN50EoAclD+s1Sh93v0x5dDiXgBJqPOXhNQHN
vJqmF4Gqrd6FMRI8JereR62ZAo9PN+dGoAOQNYwwQV9cTKhiuZmrXUD8RJbBwOoVR0fayYTOM8+G
CaXyl2uwtRZhMJ6P/uitRMIjJkp1Db2W3I/RSn3IHpeY5EtgXmWeVILn5C47rEiYlmMYvXga6kUB
4K8S9yTHx10qcdrvvDFUu7eSbYP/4QykqgXdCD4rOkgafHKXQJ57tQD5wWiYxZyQomxP33duZnRB
MI6NoWL/H9NjPEAKhbTwqwMU7Gy++PaWW3z331t38j1eSlc06DS11k7b3YaOUv01BVKQxNC9VNpe
C4P97y5brvMQWrlDqEUuyeUZpcDgaEZP7z3RnJU2sTimukr2kexT2l4V7crcWH4rb6eEFh8U8KKz
M4VfirHKCjb6xdfBOtB8Og6jljVye6mrsRd1REbmOFVYge9qD3SwyVT6N3AJkZTXTa4b95qmUqnU
CEBh1oz95Yc93wxp/hGB97F8rY9W5bo5CSu76q22C3MxIFPNy/pqVWJ3WVfm/LvZRtRqe9rtubTx
vZZnQhzu4LNtqTb2PDwFNoupgmAsRDhzFNNR42bIaKkCPIYJ+GCeOPCN0PhAnoDINvQWkPntVdxp
2AzvQithX/7KhT140iLK2LpfFqsupEjjklxpqwqUveZGeUnxuUl3/QAwf8QBHM7zS6Qxtqhu21Cd
QwZ78uUyuu99xBgQUkG48v/Bjnmw/QPXJp9f+qtjjFIvixcX3nR6FpKF7buisy6DJd0E67qSUtMd
OA1ZICWlq7tgFAQ4Ni4mDdEBRomAUiVkxu7+lN0pMkZIDq5tXDHPZRvXGOe5fPyHQ6v8pzZMqnRN
gIZmFfr+miEEcAcsHt4hjAhf49d7pdU1vEOQL8JoQ/Q20Yms73nf/tiW/+MjzWCb2Q50Gu+2J7dE
zw7hoC1s6RURGKLT9r74CBXPxRi0syfv8UmVhWohgzq7LN+wfLmB/1eFYuUcSvq26YKi98dYMaMp
ouWDfYzRnvqixfGHTD2NizaI6dF6LfoDysrPhzb4ikjVhs2YbzKA63cuq26MvErHBrIUMNaKZY9H
hSWJ6m9JmVekBCAwY0/1DOZprRp2hL8BK82I3gFgTzKXsfyQXlHjvB04UgJBemacuAGwK4yzCkdj
srV7FudvfG/DfnK2oB39SaTcaYyi0BEACSD5XAGGUccuHHg9waD2CMmeWZvUq/yaUOlYDJ/DNOxp
eRl0mjmFDwBNQTfEMJJM2Pud4e+dFckE54exjV1ulMgT17moM5yZcJf7uKeHuiOMHtCsCGZQZyUy
OIWSss5I+ioOiKBUAXCVEWIKLGp1BB8I3cLq0icz0Y4CkU4NdGlv/lLMY2+/EzVvIVCO7goO5SvC
TV+YXuMh0o0HchCbsm+uVIi0PwauvCK5/m43SS4YaTEmb6mprh61TuCxNT28jEggb4ckIIapYwEG
doOaPOEjl+qsoxV2ioRqSLneTKagOkwpsMeq+lb12E2kLXOs9DArEbqSzDm9wUk35lKAB2Ht+cSZ
MzxBpllfm8023kW4+ClTKNeYMFo41k9pKbA8bTS5YGWozGv5l8HeVDsc55NIl96x5+LukPuTzPlB
2eVNjpgScFQDRJspNYg+jh9z5JY+oGjv9XMU+wYsxX1tycNWfs5oabjBmIzngRyfExxgstOl/7kP
SzZeLV/YlfjBVK0XWuaUwerMFRmjizfMTy3wuJdynYtXIDNiogK12bVXj4+luK2r9YpG/pk12ZUv
tseh2NcrKAQGSqlbKSwCv5MNVgZqcgDTqA/FtRmqVGnaaXNTGeu9w7qq394/ZtzrFwNOm81HwfW+
bJZhfDuLpPydYaIvSsh7v0xiaq78fetRZjy8DtS43pJO+iUfUATVbTgnaazc+gagZL7z1NKUPDEK
sGDuj1g3H3LKEAwOKqdtDv9Yc+GAG/KLwPavbV5lgJiFi1ZuThoHZm1WgjzfSqwVWJ4sbzH67n8G
3SUEmqmLdBaE1TDckQIvlsSm8DucrvJs1iLr1OfuQUjtQWjNSJ7DB+LUqKEG5ksXwg99j7qq8VRy
MoHsbMRo4tzr+FeWf2wj/GD8ZoKyj5SLbDnxgZ1kKtTuljgWNrRo6jxQ8Vz6dlJtSShuywZk42uf
C7uboG7XXFoyYONIvFZZvaJ4v3p8dZWacbS1G/R3aMkjdtnUr/PXzNQp0+/W1JJOC7T67RJ0uEzZ
uPR5qF+n2OjHLDra7JS3KyrZPEdYuDZcizyvyn2zw08fgh4gHFOMZ+bBUPsNBbX1UPfF7EnH2wqC
Ucb55R0EzZ5KnQezVgFfR006VkUXvtOh9UfyFRnOcfCHsd9jW+epr0+7tYnXH0ZoDtIuWAQUzG5c
/qW9u1GL2aVvGEj8Tomjc5hH1tHduGQE4xMR1LPlyzI9vD29y+AdG4N5bkuZg21uBzSF5UctHssx
1h7rpcie0T12o6lyT3lnHL4dwY/VEtqj/nqHCuB0uXuVaVAQqn847FSJykDmtM2S68nJqph1RnNW
TzaRUv6e23e9CXv0awikoPtDzJvleC4EpqgSiqBWLfrnIjxBVt0yT7/1Z3me85Y5b2+aOaC3Ecmf
pI7e1jkffGoHDo9fqI5qp1BUyow8wY2EBq8Q3MwtM3GaySHvRtcNDiAOGiw4Jq4bx0Wgt13OtHeB
VYS7y6EG4CAQ1bF5OAEY5EVKUTSWRgQ6A/pFHBZQkqspIv9270sBiC2jkJ2ACFNZns8T2KNfhcz8
GPPAjSU/RMTLaB90SdSiEiAOtB4wciHG+BJi21bIf2V/B4V276LeiJshvG0nffOOKaz3NylmJhKO
Q2ZtnCEfN+AxbQxLy1SDGWGpUBam1rqQ77l8Lwax52QFy3dpxMqcq1eWt/Poct3FsFHAsgA+1Cpk
cOTQmiu0rO7UJPPucqYVYKUC4SxOTN+7A+qruKn3bItzYmRs9/me562In45Wd7H0YShVPMklNpjQ
rnAYLrEqjxMK3NoZirBFmbiun6w6AxESMGBkMD+r9R188Kc1eDDaXtQsouPTequ6L357BUi5H4wc
rV3lP4XgIwzaCl4nykXKDyIHmtZdwmzuyDLhwSOI1pO1I3JoOce4VwlywxM42jERaroaYXXpLVfP
KBdKydY3e0WtlfITOHR0njH1/Hjpwo3zmLNNH277L+zimwuyj1tQtpMJDWmKFSubh3jELZM1w0tv
K82ZgSFG/HRYx6MOjKpDDobC1+xWRtZ/+kO+nuviZ3xJ59TEnhnx9YKxizbNrfl+ZVIqFYAQ9umP
kPYYtPxecccmueyHuRke+7E0hmXAUxmvM/C7gIcXa6nLLrK8JBHiZ+oFNqlCXWSQfinYnReq07B1
HgpjQaPGXg7Gi99kRZ8F4XHxWjZDu4r1Beot0C1Di08hHIakzKrDuBlrDPz6zrBg5ccR+05S7994
gCFYQMXy+Nb9LBam3fyHH/5D3aX8cPAqViShw5n1Juy9NT4dPZOCFVuM0gsEhR/FlY/8V/woS4pj
RATEsUIHYABaZ7TMGUToiUW4hHY5mFTyJx4q2bSTOuCfvZ0bdj6Z/bDHI9lCamwznGHp19AMkDDk
UO2hF1mCFesE+F1qHCSznow0t8US2QnHKXkvDqq459c61hn2qfDqhI1lw9rU+cQAyK9QBipkYWca
SDdIVhFyBTYrMfk7zEstAaPdkxqHfiLS1mRRYJPuKQmqoSWlvOLfVAAwusPI/W99d9rXddUUH6b8
4lR8gqDdXBANll/RnVZsBZpT0tGhQHyM2WAJ/QFoSzTGu5iP6W4h8qSIbXvfAwwoU3PPDpbUdX18
kaIRvmFGNLcHvR/iAwX6yiW/aaMBVqO9Gcw3bz8xqchSz5PtmFTgdlUhKikOkVOuKS+NU6jY/4HL
Zf1YyXlxGmSoeID4faKZmeyNby1yX08q2HDO0J9jyAtcDr8gBiLc39Wvnvj9oBzu4EhqxPY5Q9wd
OIExK0CIJN+2jbeBY89R8LwxdqsZEQ04ib610ypmClbIrJYUm1pIk659ivg79Gc+hCcr4HJt65hs
vFrANmXo89JZp7IG8svcfVniYeUwnDMpQ+bhYvh36oqmCoqn7QRJIsUb+bBY4+MAK8Krdxay8dHl
62PxKwqG9WNigv4Dvdb/z9wzofSgsw/dhIt2IgdkWQki6eK1589vaxhOeXHGlJI3Ue8Je2k7rlcz
Gr3A3N+N1XHIoAGDu1KILoeuetX0liyx7Tmzvigce9ZVR82wpkBftzZXCEiLgMu7gFz3y/mM52Nc
NOKEabfnBfPZkip5lOc0pvhd3HjOIDqHIWmCs4UBRUfDoFhm4PvkdR/cIkEB6Y81toPWhT94Rku8
VD5w3GB9QZ0K2XX9iOhFvwBZK/xT1MM3g8z9k30gw2d90zO9+ohA90ZDLQbVz/HL8ipq0r2MOcwm
rnt6IZLlL35FpPqUxsZuUFfzDJ5svDq7Igca4M9mM31ibSWBRG0JBnRXOdXjUG6k4KHKjWGiNFHJ
jI/ubmq0YVW2pdymopLafdsJEZMO3ZJ4RKFbK0sG4p9Js4+MNgp/5R46PK6KjNleZBL/zWZLRg8I
AIhswICG6UAplCnIcyYG1MPVulo//iokS9Q078GG9HvnnSVB00PcwD93RZE4jMs+rbHJfY2Z0qwN
D1W7a5rFgYwcleIjqVS6zqL2ErlxV09cjWZR6daH9QnsgkfnQceVrm8PCh3Fo9qV9Y+u2dHr/MVx
s/I4JI40XBRbP/WsRLrlgvFh9S3awOQL2IKehGfhJDj0eBxCMDC0EDq/r1G7DXzmQJKUrgJjyq3G
2BJaemkc80Jn33vRgOT6nCcyFDmZVgeSogWpYbOVRbcw/HmVWGXByEWCPyJxKjLY2cODiU/57LKD
mvW/xdsj1ds0PvCW6JiOxS4cNq/3kZzhv8gR4AS8sUudRYmilO5LiBHAhRp0hT529imrEiEaqaAo
/1ZW9/UqtiUzTQvQiZLvUYzK41mI9ffbczN/XS1p+ayLO9ip72oRYwSuSV6eCLzhyXjsD9YwgLbD
Lmk53nRLSEYbxQSEgz33HXAPhXEbXst5akFUK1DIca7FcB1VYMqTwEVlLivtdoYHLUpzYqMf1dGu
6PLK7AwBgUJ5GpOh1rTTWWKz8j3a4YafkR8vClRVUIEcM0EfLybRUzVBlwYdf8Foi4ZZ5/GbId6M
SCSyNNM1lnuddJweyKcbAbfXMsAwWySYcq0CT9A0TO3eg4EZ6a5tl9KNAWk2gz3RgY7V1LfbkpZz
8SUA1ozmykDNEjeFMryN+l8+mP7Acir8gZ+wSq6UYtN665Lms6nHLQKcRARRVDxbDG2bO/44VuLl
IiOQ++Bywi1LBl8CQNmRYXcf7DPxd17Xa52xHY5Pcanzhh/KWXEGzlq/CWtWr+HfDHmvs2TeS4Yx
eNvwWtAEQ1JPV+Ta8RVtY7t3tv6HOTLtQeQsLwzfVG0nVayRPZnWEePjF8xnzy7/PL6aLQvKNg7J
A+ljOq2Ak/3PQ5REpd+WlcIpW+uLfKa4741NgykpwdXU8VVyZ1aXZowOl6f4G0p7FtZPJXXvLuik
NyawihqCGVCq4tTPgvEagzAOeqfMYbSnnG95ietQFSCIASFpZ418xhhualp9i/4mDxVJ4BxKjC2E
+DjntafhOMy4lsAJ/NMiSEa0BEK0MQH2mw3V/jQaQkLxSpQzAHcCnnBgHRav7WSaC3/zIIIGlM4O
Bzuw/OJJHcu+c3b4hfaDjtgzy6iDsXwNls2IJ+fE2xWOUKCqc9es0zTOWKFW2r56DcHq5JIArpY3
YisY4xhjlpfK2lR8U191ykySHmrmXJua1A1AiMg7dt78Ncsk1Y6XfOR9glfAgEiEsaqrcXZhGkjN
XAV8+pJH5ItBKIPcctm9fsq++J39NtLhJBex/lM8sH/NSRz1fuwsmWg9/29nwjtqt9tREWBQGi47
6N4CAivb+rsewI45scFbfOf6DYzjNvDR45/JKWG7wcGI1JbSyw+TTIrYSOvu76bCkI6GlfvQL+nm
2CaM3G1BgKMZd0emRk9KdYjXYv6Gqh/LtyTc2MdcMAM1LDCQAXibgUbBqVNgcWca8rH30L0919iL
8ExnqCxZsTpJD1bIULgnoe3QV6qck4Q76OQwv/KCip92b5xTdYG3dKtYFIGF+HDRXyY3qmoO0a21
MjWnnZ8vM17Uvyu5rZQxbyt9xWWeQq9Z3EBJBTbUG1nCjLwWMuKb+YhivSuZHSEOWZHOlZXWsCMr
/NVc/FMzrlYM6TEwCk/krdYEh5XwM6ld2bSXUIR07fnXivsP2y3aEdSTJWOnLNFukE0fs1wBYss+
28q9RDOSh/l4+R0pthcwxjXvbt+seD6H6l/s+8S+nzrntYVOIFrqywkxrMmee4MzqclER9STrvRw
rjgyyLUNxVTbO7WP8jynTKM81/vlzZkJIDExGf6QRn9B/ZOkv9RI6ngXirV0PHOzdjNc+19hLSOV
fYI3TDdzUShxXaRIlTNRCoxzcWTdWkivoy3XyuGGtjRbSIBfxIhJlW+rVmSguIFxTnraX8wrvA5l
Jd9HdHE2FSM56rvZmwyzOTFEgBu8ozOOegxCkXX5Gbej0In+S4/U9rrfhwRQH0QRnTt/oZ0vbT3+
Jf7Bx+rpSjfOiozAqimQTM7hsN4LAcDKDSc9IfcLyWwhPjB3UsZJIyBTIPHnZKLQ23T9cIJUPnWY
RZm8Gmnwf35FOIitS20jAl9tDkqgbyi9hl/rLfSA8mMpHSqdjgT8bkiEgZjo1lBx3blBGPypLZj1
UZEkB7/I34bLgCb6RjEhoIqQH4e4ZDOiQRrwErOPuMSow7SreDA4+VFp6IGaUdtRo1fg7wgvRmSF
1jdWragJl2oREkGvck0G8lkgVKDfx238g+dDIllqLWh8A5UFh7erD3Y5KCw6v3b+elExxHsZH30a
1es5IHeVPVSUdxJlhrStg1kd2w1djFEKbHNKQNIS0mFA+4K5hTyosRshRHWDeB0KyUyE9VDRiApz
lGTrvximXXvWGP0LZD65DrXhI3X8rhIIAdwy9EHxl+50bAUgoAT5YYTYjbH+bgP4GlZ7g2Py2NgR
kZqNf7kSmwYzwJBcsTwTO8pxc5BzoGRXRvxX1dENYD8zyYHZe3S8BlbQAnhVHwICpM5Fc3Ggx+0R
keHI12an3HEPXIQp0bwZC53uRaV2PYPZLBN2AscNS4ODAlcZlt3mZEo2nnorRhiEkmjhau6SqO3O
MFvj23EaELCrlXSxJEXgFp2jC4+K89EHfadxbUyIQvAhTOe8i9A3guCRb/wOflaycbz7JGbXcffc
PxXb2dLug6HCfS6iZ9hXwiVyTKRXfD+j+TH8C2leKh5i4P0aNP0Wk4MiBLFjFSE2Zxb8Tq6FjmJ7
HXG6qVV9UnJwVdNOpve/0BN6CQ641mMADU/+r94Q6t9pTA4fzXcyLNkKsMAxBvU59o7KvTGotH27
xAPkDCFtLl73CUGUtQpfqljbbQiusUBqYE0I6gMaiTyRdmI2lcQSl40qYOM0yf2VzqzRP8YDvdQD
Uhbkp9shPaYhCCHRs02g2ChhEYbokeksy9t6lzTamhidKwjmTNDVprZzdr2Gn0T+uIMIkQ4Su+uM
j/lg6/Y6t/rfUXNEUc5skaTvs3hJOD+Zj9JCYJynSjm112S0ckbC+OyYpnzsHXjAn2hPpM3mjZcc
SszSO9viFUkHYRV9bTnpRtvCvUSjPFxTu/rc7aLnfbLk7dB8e6sXfNjDjmVoRwlBR4QGOJq6nUX1
7mNo0+0kg8qByenTq4YGqpH2bZIvx1XPt38sG2pLUIPPuFvhHv37mVA9JP9w8OKQkKup+dtjkeeV
Gw0g5hU8AaaGkgse/cIxGn3cmPUwBgTnmuCuPJ/56OMCoytkzuKKgZgpMG3yhv+AbKvB7Xka5wEK
Df5wKT9OJ+AYidB8gqb7dWS/2cbye/0h3IuxUcgmC7ugByqIDI+NzaiqBbGBvFw5iYPVd/JdZqh6
xUHqZYKZL/Y/QSAbZ2q5SZJPJ4tZcTVK6F7HFad/2a2ZopNVdlFy6SkFeDmM7hGPUL2dwD8DL/Vy
i5eEVE2t9NZeiv80ijR/O59BHUKbwRLiItkq6Tgi5qkd/d9ymEx/Njjz8gn7qVVtRDW0X6+q8N8z
RwCPHbOQRusldUzy84zkhYo+Q6YSRsf157fxh3HzWZqVxitxbGfjjfCd/hAv+EkuMfCdmy1N/Dbs
NBX6rLAx0IOwgRVFF0H51r77FAkncpzPNcyaYYrZjzQfz4KD+ElGLO083nOb+U2j3EHwU1CPRgeF
csgqyXnVWVYjWdzc7CVuVwT7UpD803zmKVPgVBGbIRy2sDnE46NniuzQ5FAjVmPHcsxUtfPz4KmB
AF4j6PENEFLZLsNheEa25ooIM04iNWIG4EolL7FOf0J/sVgulQz3lhT4AcVEi0lOapf88XbS4Agl
d0TF7WGwRuHpBrMmnX5Rsz+ZUhYi/xjA36o4zzcpRW2d5jPS05APQKnf/w8DSQ2Hq6hoKxT3uQiA
ViVPwyTekfeS3J7Wa7OP/ll6g6gPhgzfwxO2lS9i2rWHf+ciLuXXM/sMIKiz7A9tolQqcQwFfT7V
8BHH2AIwemVcqDIsGIZekAwjmjDK/cZ4DYsZMftZni/SnBNBTMO04s75DaCrCBTtfaYKtn7UELSB
YcWaG3CMEr+JzW+fBURXQIp4eV3RLQJN527adTEpn3dzvpBMmv3gkU0vvpP6vlOGI2tDb5VyIfQb
RUwespsFWQTed3xyQ5CXBBtxtCJjy+Cjij1s7hsI9JWpGp2NeNubnB3It0XWRLbVNhamHUrJLFVk
cFxDmfX2hNlFHQM8gI+lW7bIx1cQe7/NEvvuul/pnbTviFuWkWdNxR8SQlxQH5NVBQQqYgRvoADM
g6vB4iQ58PKW7oWLMC1YYjvBYSA6vOqMvn92xNI1mvUY78jAwuF41QCjNzc/i4lY3NgfzGo1ecRN
k6wVn9CfR3JEDsPGE+idtykSqTIEORnKX52EMvecBum2P1ou+jr9R2dMFbGAd+Pno2beJ730tWez
qoeObdOVjz5ADMPVXJmihyPnTRw8zO/uO4bdCmvpehYcKo2e4ssu/67KceFw+Cd4oeifJ2RvdGAL
5YZi8pT3kG7mbR50IK0OE9AY+FuEG2WVx2zLiVcRSlYWN1f9t25oitnbuiv3Brc6JQETq1iV+oSN
vAF6916zT7ikCoO9N6IA3qRYEXGt13uagcs/3r5wJ4xL+GW2G7/RzCE7KsVme6tHDGdg/a8jTvbj
ED6yv7QdxKc1ODOL1/7zdvgFKMefCYMIwKtBurHZ783dGS/V0VOaja+iXIOUIL5vUsFoV4153sxC
x8dPiN0fbxIn0h+C3NG0MHNNcEaGSP0ep3rhFxtPHksDfQ4AyV0yTOfOxegCwx2/XVEHdBjyGUpb
ztQssYQcxQ522dSjyhZfSw5XNXQBOXcqwPrO//pSV/PXPWcnicufATuQ1I7ynZZAHjdGn5Dyu0W4
jOPzdYf18WzUepIIKTL/KAyJIuupCDMMtgcLkNy6KHRx+iMw6IkHA4YWaGv1hBIKesrzEfuhRD2R
kMOnN0YC1GiQXy1iRwFfnuy5RGxLQ+APNymd0eEUaCEHXL5Bt9nu9jc92J1RID4WVP8c2KMc12Vw
5GoZMzAflpGe6i2q+RIXbeBZ8o1QPp9xgx98YXa+tzlC1nO872HC5Twd3rGreJW5RNCzH7/TMA7I
azb9tN6jToNp++gKjO0OjMjv3WYSizq1X70n+4ledPdvNnLpThnhzoBiYUVr6pzpmkD4LTsJIJe6
Gf6ZVliNkgmBVopznNaoajKEl8b1JzJCcu3qdS6ot3FkrW8NmjFbsKuDJVZcCQg+WJVAKJMUZfjJ
ZL0pTA0nVddZhk22r9HzGl2yOY4S8O6zryh7HRj02B+eJXNrb2gAeCiPZS2kXxkegeYC+tkCK7yD
NZHbaKWZZWB0J4yyohxuhsPXMoQtdUF+UKlX5eUFO6sqxG4Y4bFUGzyvKoYDtoQsbADv/pTuBxbn
f4meS4WHYJvTW6CgkMbIXik6TX2ykY+um/6zCdr8dxuX+9r4ndObvMCLoPn/o2CxSYp9qqcsQqgE
0jO+oAPAd6ZCIwN9EfJgPVs+yQkA/xL5iuaGFKS48+V3NCo+tKmQ2qbEewbpTKdCJrucrLp5kxA6
Te4bb4ytsdMDl//ND5xg4IFa/4WqbL2w1yj50CDv3ca8fplfP/NoxWWCmsWnB0yGYM1bfvm+MD2e
D+JYHViKpShGa/lI43VyfSSDiLId4arWXNE5CdNajorQ2bhNujVGVBt6nAkqwesiDFoLcO0aaO/2
NIVUa2xlHQps0AI8KcZqo2FLPfGHhoXvTpaN/pbR7DrD+Vuh9/tVPE9CN9kGvz3bi642CNlWbPRR
tIxBVbi/Zn7yd3EPD6MKKtbUmEUsXyqaavaNGYb5ZiMrAJT6W6+FTzmjxpZ/R4RMCUy1Xh6ePzDl
exuS2QSRCzTiuiNDSRqIWQBrtnow8bzUHMJv+KbmQNr2vMjo6gI1z9nMNP+XU0rJkR6p8tVfKBFG
g/gGUMW8xI9+xyA6zhbIMh7zAQJGjnbEFGfHzmxr9DFOjvvRzpjqEu9Y8zrbXLrkSeZkwPxXwFJ8
/U0WRRv+EuQUp9sfAssot0RV067Op+hdS2wM481iMRWvqHgBg8YTHZ67Fdg3JWiTi97raY1OsxqG
DLtZI4ErpelpRqtLhHQ/4emUZVTPsRUj4aaQpr3l5BtcP9LfudomoCJx95C5nBwOgOewxndqDTBM
c0w1s3R30jfXqoZmWWsvwfq2m4KmdlxmL9Cx2TetqA/A674yXMHf6Fet7f0L1KRZRzcyu+iydfrL
B/n1mIFyMq6X7qRa8pQpBgUDfQnu3+EjWpbkIRrBlkkk/7gW7wLVitV5niQNCYXSF49NjAPryCwg
2bsSfiO05gaAEOowgy6d7eCEDfwtgSjLtj13JECSSEA77Rgl7n8t4eSiCQl768pwwjYIdDGVlEIo
nT9oHydPyC087IwP065oHb/wr17ea+yEezBUS8qJbjtmayW16ecdXJ5R2R+yaHz7aS6SN44pJ7vn
QD9KFJlANnwtc6XElSfsc4J9EX40XK0TnTZlZj+jdm4issb+1PNOpyC0yI+XSisa8dt+SNHOe2EB
e2Xt5NSs+u9pdY/gIh1UJwPJhq13s6gsegZLCc4F3bpBmnCdPjhiKpbetGs505Eczo7T/JEx/Gwj
Lve7FxK0OGtpRPr+YwmOlgA3NsKSS0JjkaJDzlMDe/zjNkkwUsW83IbA5pF4QeSD0al4k33hkrU2
qdjvOXmcDC2CpNtO8l/tagJzSQLeCEAXb59vIBZF9b3cSXhH4o3NVaWevL1+IxVDecvlL8CRmIj8
W76yHnqkiilsoih8Wx/IPcx55DaMtcpZooakKmd1zK3O9kLXtCUwiUJI4i7SqgutosVkYOvw9ydq
gH5PAmM2Og92JNbCHoJW6omVP5iP+AyhtpBaz11XpwfbdG2oNwRVutgW9ao7tnYzDr5/GnBXsvXp
eo+GKx6btUmoHaqbNnZjkpZjAKDZA28ONTU/oQfDvj84faLxdf55TU6/gOlWN7uo6/NEkLvq7Lij
EZA00ShVHHvPqeo383XCxs3Zp9RUEm3DKVLAbsWJBHAFMfH9R/osp8Kg8EF5Dc2UuGn6bqYDaLsD
A2aODb56gWv5+XC2kywOlSyJ3MI/N8GTJUQUowAHVOnBorcGMDd6MoMnmwFAqdgjLJ3JpvJRijw2
q5rwSr9DrE6tE8i4XtlSIdvxjjztmZXMxcYLBGj5WPKioUUVrkWsX+H4OpiCM13jVaL8hp4tn2xq
N18pELmmrEPW5dFZfiymnjqEh2ATXCUXsTq206DGoIz0gmLsr/9gCLaTLgcXijqH7zxkRwOuZhPz
DbrfDxwrQdLNXSUgW73wtFZHoEt2oAD7Jg7bA2O6xF4vwgDA9BH/CpHJLKXBM3FT/KDHDsBgCMQK
JWHjEamBE2nE08+SrhMsEISxSsYmOIfjW3caJP0dH0lGXbVlrn2vYx1k4ADeapWH7G0ZKt/W3zzW
+ihZxIesAi/XlmZjMhDVwXkWvHZhUy8lRze8oucvT4yrsR0lmU5bwOFq3oRlO0T0/Fxw1OlX1uah
CqKQDeW7OBVGCMWeLDrZV9PvUtztKlZ3/nu3KJYdIjFcsXBjXmjy+C47ShWaZPOh2FLapIybECQe
+6sB/rvZlJCYqPY/5CbzYN90Fp8RKgMfx85A7Bi7AuFFU5SgmQrwrUyR0DZGIbrGnTtu0di9v5ri
sxJul0siQobCg6oSjuOvJ1N2gyZqKJ9SdMTYY3Xz1sGsTZWx2HU/HS2lSRrVFhofF8iqAuAs6KUc
96maWPNd8XxRtdGG26JekOPbIHc+preJY0SGT8oJU/87Bdo9l8SzfJGgPR40dLsIFbHuuCaS2gZA
7ELCAYYS5VmXX7Dr78eWrFliI0aDvf5VuawGFCNW62+xkj9O1kVOP34RiegCaIeLgoytY87dVssW
I1oxLp2NhmZWV2gRxHKYvTPkXpXAtmj6IVhseHiGKmfxVi7F1IhuqgD2wzWIcsq8YH4m1dVvuJLA
LbdxnctR9vfG5EKZsWUpCdNvG+F6yzty4CJpsc5ElCGWDVBAXbmvjVmLTC2TM51Fcb5MNTF89LT0
HApGIEFcmYx7U8KZGKGQk0Jqdu5sj3nq9KatLuDF4bv8/mzu1L95HfeDya9opQR8HO632exdU7d8
MUmnVEb/SpLMdhcH9eoN/Yg4Tm/KgHxGdkt96Z40FEjJp8lmYZsOVmh7eLWN0a5/OICyVk3uywXc
mU2nBwOQS5W9WZBJFFF7xL5AnUow/ECshSrVUAZXflsTTrS94QJzsR6buWZvM0nuEuC2Cr8i+wpi
/gN1uIbe5gB4jkEMuzGAtnUqmtrZ2IpAipED6g9xCdsUXW7TcSLFMNqJDc6sTkaFWJBabnFNsNPP
alKpEs4ilIiNYyiBnas/KzageCCBb438+b3+AtXFg+6Xyb2epYVuHare+FiqnHdNYKl55wWdl+Ag
6Oy1jiwyCGUpemMhFY0bP+8wqY1PVErCyiHRURnczQByqkN53zUFdX7u2vukJ6jJFUvB81jEQZrR
NFUiG9DgMKUmR8P4gt9hlzRqEK7vh/fJDo2FyZw0HUS0y/ZoSC5imsqWiET7Ixi8hdornLqITvJG
KfPY8Tj+r5TdJa7pvApp6PME/Map6aUAOzh5SgczDxF7vAnnPus4JJLWpyfhQTrEMSsjTRkPcd9i
mrhQxywrGwHqKg9fhFzEuCKcr+LD6LAkE6x5OKnEAi9pPhkQ0jWLcAJGyfcuDKiZru2OK/9wX4M4
dgDhFMM3Srv9oiR09N0XF8GmoQlyLkPeKirVLYOZ/V9P+sfozLpAahHS78wopuTedwFHrfKbJxkf
1V25AlYa3jhLU62dbaBya0WhHC8C6b9lF/sweX1QgbktyRSqqQiQbw56jZBzxRgSa84ysnc7X/V7
7/xSa9ZPZ2V03ewdBYh8Tuj+gBreQE6D3ROanaajhVDadG5oBLnkL86NLyuGTLVB8uxRg1oTONRc
Eg0QPngYtMrAEe007aLTucvBCu9M08R2+ZRXiu85x5lzqPLJ44DORviRRj0uNoGSJMFc2kIenEIE
tIo8GAqJWx2bVwp9Q7d3mzJ1Wb21umumFl3SukD/U4eBTv9/tMt8cR8wIrmd9Udn9NApAFOl7JXz
yL3trq6gerMprriz3UWJ74yE8JLf/r7IFCwJvVIzBTY+ZnQneTDDTFj5HwHX2sSQvBhMFynBiAx0
vYfIhFaAMvFuJ+3imh9ILltKyD43ETQ/rVJijKsmX4J6PlXAiwRs7Wyb892DjKz/t1GxEc1BEXsC
bae9gJRx+jX+CldouzR26Xt6BSmrSikdyk1CEuWhl9Ny7ufr/qUthXf53uP8FZK3RS1DugXBCAJG
pbjUwFygoIKt3Jnr7lvwiOhWUE9NDlbmlDpmp4XkQruselXc93BXMerLZwORFSmwR0MUsc428z+j
84JPD5RgYbFFmr+499EJDkXPL0vLL3B0FSZOgXynZbiorv+rGEPUiAwJGx1Gd4VJPyplJZeavZwP
/XKbXnYyXGorX3rCksIecP3Wwny+hKuO9BptJZovAcI2g/CAcsEAvkxbxd6RVKehl27UWHqxT6vi
XFsut+dFPoZ6ME+bntUBoDFoFWML7IEUUsqwq46UR/zQT4Sffw8gRQ2UrtX5Yd9ZUfHufm+bwvax
OlPuLkG5V4ksg7Sx7n3emzslwlN8kfYah+dcxTq+z5NwiMcwm8vkpI+UyPLwhgUyiXU8gHMkmmft
DxzBjxP7JXqHeoVUkooG4PMnofIKBC0IM229BVEkhfZkRBrg11/wkz7FquCe9w2optZHgnTQyVPV
y0tV41T/vODzOPPDAARHZ5nLuCjJ6OsVyN/Cq2IxiiCUAJDANGVfsMjMFAKgkyJWKUQ0MMuRVPmo
RmOXtYOT88BP/Kn6bhr/CUTDgB1kgex1pjXGJzT+UWI2OYkMrKUVHNhWophVNc3WQf+coZuZOLn7
KOF6DbHhYnW8R7bCBUPdMWDhQWRTYHa7tgs1mPI1FyEG/bEqeJ9HG6uN055kdkLdLH9gZ6bvL3Wz
P8KsCgU6yzOiHF4a3qQg7e2LTQcade5j2YL1mSBiTnaQMfN7vpapsnKx0pJsQCxhbWY8DweUGctp
2S8Onw4Uyz1wihSQMUMdM+kzI0p/mUrMdlX0lULfcLLHE14DOQoIZXKB2NSGMM4gCTKOE1idtFLr
HhTpTb57BOYqyJ1Ul8u8Tz47c2NTjvMmhd89ffY1d66ZYQ2DoI7BC3ayiU8vRbj9oxZ9vgZTCrXb
iNlm2u92/K2EzFRn9UH45L2PW4muNwKrpVoA5B2LNgeS90zgXoJ6Xz7E7pqGUVoiLgDpndm4+/5v
mpce3ZZKRlA9ZbykZau3Uw86HtTNnIJWdz5mFa2r49gLuFzvyBbDnuZPouAhNy/lzOaW3nACE4DD
bPEgZ/oO8IcCmYNJsarmzG6Aj/tUI6bn0/3vxWbxjXZmxLnz6P54p9Vbehhbmzdva5C1sJICc0jL
UNQNXdIAHVYte4I/gu/cDAYVX4Hgu0sp82bpXpWEI62Jo7l6riYKic7dQzKuwncEgoSAPKdGkzjx
qeREb+oq1+nG24Bwkeq0h3R+NAQjrTEf09ZgoeAfxl5qYBa6ZgipeCr0+EVZ3e75rmL2wl7kyb/1
yxk4d7CPrdldqNPwrB+xYtRm7roNUZ0sNwjxSLwl3d9OqTsGy9rQoPxWEUEsP33vC2aZgU4JXQwQ
PgSXnvqhB3s8mZUaRJkv6P0OSLHBRBRu6a4MvqGvPYE0B2aKVGOyqUyejvdRotrvyUlzwLCxkY+I
bLLG0ZsvE+EkxgHBRENmqJwTYxu+7fqPUQzmkDt2yoSP/OPT5YceXCZv12Jv3oCQXnFs2gFtW+Jt
aWUjzy4qX5nlxsu8jEipxOdpwMzogiTSdynUViu9lFPNaTUkcAb9ajfz2no6UfTZCuq9hcpyd5yE
2TBPw7mCAHr5Mu+xfeVUZJQvCbPbq8jofp35Z4CSEsSMJKE2LBnjwlMGVe0JTBC5egXoEu/3OUmH
uiuKOEmTLcbxXzk1SNFY1UkECbmeoNkhEaNtgAU5Tl5i7dB23C4xitmtNohYaHEN++s1moUjOSwO
9g+T1dRre6xq3Ic0GhB9ZmbpG/yXMM7fIxab+K0yzYmEUfIIKtCHvF1OwieUuwJTOGlZHQgsL21Z
z8BVgtov2Cbfa+J4GKxNwQH1Iz6x0EGZGeWJHYqQVNMs7GGQxjdTdNM3UnT/A+HRi1YMqbt7H/sm
/etjsYTk3FCqjC/ygwU5Wrkv6scqMU6FlI+BeQHLvuwWbKkyZJcfF6D2WW/IdLRd3c9LGqj219se
V7aH2p5RFcDdAtgVcELx9cUtgc38FEO+X6MMgK5KohxQ2wYt7aXHS/debU0IQUgftLRisf4mAWS+
qyzUb81MkuEmc+vH+IldqDEq8MtDUNBaoreNV/YOz0gHwmQwACqECglCaVzcVlBDivMNPRfZeDH5
GHrH4c4LUsWuZ63Tkzjb0qRpKsIO3ndpNllCyt9fdXwIW5MIGjyGiIws+Nm8g5jvMu1cbmK55hXr
e253JfLgDvStznVPT9oXLykB9pXIliUMiO5UBCzDhOZJmJvEzG0dGpa5te8Xg+icKgrQR5hM7K/k
/3P9sq+Rmj8wgxPBWSH5lj30R0V/hHQj85dqSET4b2DAwDnrAntIl2hgkj5l3OfkOndOXjk1vTF1
4Sd5ovtprY4KX9hCWhpklhiQLRqzz6Lu4DKqaceFL35tHsGZC8RfkwlI6xtQCUTng6DMkqSa8pNP
LZqRQ1KAwyj2vsX58XLo6j53rcnzZGKNBGZ3odM1NMCkZycVzdPhu9WdQb2B5PB7kxD+M6/XfphK
YyGy/PYug2ZNOVH6m9sUQsNhBvpoAws0dOpWH+4M9qOs3fFoYHXpml12BCRt2AKdkPmQ91KcmBi4
SHBQIpkm9tBn94mNg45LfRqh8ojOjxVUz0ZBF41NWgU+jD/QtOtxsMrPB87HMtRFQ3dSsEk+jUUB
xNnIBQogex/RsEuQ1SCObVCjR92pnS9LwIpVz+VqrJ/P39cwJNtJWXzb3DDr33q/gBFYfncWoSog
EBc+QoAJtv8H+1LoGD1QJYdiqOffQ9bgYAhPRX2F0575MmzdLcnenF3+pUgfTP/DCTD5KeYCbK7J
kHCuKatp403zMXCYKi802IyGQqGF5zztvvQxBg1KC5NPv4hZWkzS00M8qDsHrvbsNn5Z7YbSZ4b5
UTHBJqO887cs3W6hEkx4N3B5kNifvyh8I4IvnteQQnoeIArD9ohLE7GydkEg/cakZT9MKAC+/OQw
mEwyP2IBCyuf4v3yH8Rb1PaiqM+rwShrzEAsyLJn5HBKHn1Z+7hbLbR8Na26UAo3vfv2IBgAcJHf
s9Bjno/xu5vU6QAh4v/g6IEwMYjealwJdsM8ybDZ88/rclXh+EdYfPoKlVK7RZOgGzjjtMe7vpUO
cos9bMDbKtX0SrbW3FPCh3qX6gMbLoLKie2ml6f7GcLkqMsKwx5C+DZmD51SXOHYGZLtwdZ2IHJY
EMxFpH5t1kLkJlyodYKUUq7QoukwHgd3wAMZcuEPujtgP5vrbj6xXbL6qz5DhUJ4qJZPohGwdAA1
fzpV/TR4TwCDuf7Vs+l3BWyhnDaqTko68dLze0bGk+LTDBIL9uXxbj11sz1AmTq3+Oto1IGWvcwy
SPvtF6L6TQeEr6yK66WTTzL9nthFh6/TqOGmuYcFXVQE299lxChGxXjQjM1Kkb7nyUu4WfL4sI/N
MdxzX98biOQpOc5TW2enZv76IUEBiSc7zsjDV+6IdD6Sr/HL7G/2TAwqd6jcKKUm/x6BUarMspja
TpLH2k2R4bmEWu+yufXQHI9oVhfjnB+KnCEKM50npmQMvfty4p77o0Qg3D2m86qMRZJJl5TuhFkD
NdUUv2tT0tlVIJmdtuAPqgWmrFqUNXXTlnnRPzv5ADeIIjSpFCiwMoSUE8EJMVJZndP+XD1QMMRh
b2r/u86k4HPY7241dnYJKJI9uEUfAWSMp5k8GMhODERUgPDTruaYBd2GgMtHfg4KoNfOZK3HNuyb
/TvnTWDKnxSUHHqVanDpQZrk6d52EkMuTN0WwDQrv0i12MLES8JI5jP21zlXovwyAjhEW+eTssZZ
sr500ZCbvE4fYpkCuoL1jHyVI6pjNZz8iB1H++qHsW2bRU/zrGLs46cVs/UE/Rgenc4+LHSXFOKA
H+TmzQ5+ftkvwEubtIzLgwwrkLnaAEFgKz//Ao+SANxDsbmEjbuOSrQQOFBvv6JWWp24J1uZ46KA
4PJJXKdAxbFNPkxQ0D17kKrUUhJgGJvRKh2FmPlSBFCLL0N9+TyJSh+kf+o5KwHdxOpEHoW9Cz0W
eMH2W2lFypBq1mZVVD5SryL2YsIuY7pfIk9PfE3pQU8KTC+wf+Kc+1ivi/UsJEzSLIatk+oxkKjz
GrvYQxA0aGatWHcwsbwNV/f69HVgzgHdq9qLuIKbvynURWUCFbeHxXKEDy6DF1wBQ8Kc3oZ3D/Je
YjKkWPLSWBgfDdz9BFIjpoXwdKmjjjgXtLo9MEZIXOPWTr49dpQyIufKBTA/BRGvSNtswi+1nGON
CouEd26kvtiCBmisyEHUzhfqOFEvMPmbn167BW1IjDNiHNbUOzBauuP3T1waBqcCsRqEMaaLRM9f
SAtKooE6ymAqEi5yML6U9t5unGcYJa0TwLADQjWZOrmeG0+H8bO0yIKGTLIYgH1Cy9BFVdiy9VdC
E+8ik0kdIMx1TnwOTgr2idQsCiSvp10RsoWVwUv3Nz2ugeWo7sK8Hzi9bES+i6apw/4JXiQeNilR
X12Ne0AXalxb1NooYiYCn3q8XD21lL+5HcqdTeFVkWFdxBf651JDZ4XIDRUr+2vo9+pTjHbQvscE
GsS1yRvbnUIcGd5tGNF2F00br5SlYm2aHmr76HyV8H1h0Zjy0GfMmZdSYBsI+BwBuhLFuJLJVwVR
TI9nntwqridHa+Isq6BZsIfJjWoHcGMe/ygtG3I0P8vqoNmxgDcRdF2nfEph+txcwPYmjDXQT6Ly
xzc3Jn8bhSwg8fPCN/fwxSwYVCWtFKNA/60ITRRdLjTNyMz8rvY3A0/MFhUVn+yIqJjsPkRvrx/w
I2xEBKqBnLLsPrcR1Jw8KKr1W33iyVWHDjPXX6a5okoMjIV4Voa/58qumpBnVYbOv9GV1KxWpK6H
lmZHdtMio2wKwVwH2ofo4vaZt32MCgYnLkZQKvKCkWwzmZEWBNEXpJTfMdup/XPpn58P31OubHEn
7sKy09N/yos1haMx6DKSTYpbOYe819uT8neyxQQWr7Bds80iJY5HTBfwFFpokjO4sLTpiZOK9oG8
F9xQXxwow0sS0pdct2yXjhv+cO+ajwEkgIFefyFl8rNiKrRAC7WSJqvgZWPj5twxxWqJeu73d/sb
W9f2tkaT5gMeIwfvsambazTbfDOdHoDINfiPkO8PVTBD7ys1YL0VegYuA2XU25dPrccyrzDeekmL
/ilBz353FNZEmGCgYKg0zIoUzZTkRIiDY0LnCj3Mym7uP7NXB/I1rIwB9eE9OstoP9zMFBelLWVr
P3BO+zqualDO7aLpU5VztLmrsgnXlqcDL6vBFvfTC0ge0UencZl8x/o5OYLd1N8j9ig05FvNvsnq
Or9dU/zu4aGNcS835FOY8yB+TqBR/fNFSXf+J2SLKe7EwAZHBYsG0Hwn0KvtKnuj+e2R0kwBLEDJ
cRo6QDyYlL/TjMySNB9NCWRvS8GqfMZGICw1vcqh6f4HX63KwNzv3Csoizw5GmCAO/s+VI5lwtkV
Y/L3+zLGZteObKmYokaL2ZGKqceKGMAKrVeAifNwKuey5/gAM18uIaSNdlWZY5pj+xGdxHMqgsrF
uKZPhpq9HQFlMmVUW6HtmLfQct3iEIKIx2zESKVeEhWNUA63jo7Y4wCtAIZKBN5qJu50ZNiNPBSA
I3PHRJcq7OxGbDnmLmSvGnaAtNeQy0M/97KKhue8W4/rZwWmtG5rZAXYyXchvBvHkrONyZgXYwMM
lQaQCfnWkaG+PTahN60844wg2zZcnJ2FeVdfOj6gj+FAQVcdxHHXclG7BO3CSw8V9A/VbC8vO5fo
qKf/LStYwoZwU6yjCkw2aQHb5ZUBrn2UtyZnHDiBZqTw7S3b3+AxopGtuqsjnAkdbymjEUde22Fa
G7pGHjEF7SOOv80SnnPmcYY3ojj/0lQrV/KFYkGthvPCJBkXT1OMJOAXETAAtc6G5Dvg9xzDFbVD
QOcgnvNSxcfTESMDC0gGPIkYFndgnwtRtgqdM2RASuXBAV5467Pe6KhJu56e9XkR7jjq3+5QtarC
Xmgo2rCVIhyjMFARxsp7yc/GtbM9qxHQ5nF45oj30soBUv+NGQiYDRCo/AuvMDhY+LzTGhhAJydr
5WNz8DI/I9jzGP9AeuWWTWKn9slQ5wvkSyTknNyMwBBP7O3p78NaRDJ/W02LGvHYnaHfGwCa1OXE
JW1TUYJvUIFFLqm/JIIZrRTQGLzld6tnbRI3ZaDPxyFsHXKwIJndK/mzF0uLetj0ufDE5WoM3AjL
QBR5smMlu/f/0yPiOMJcRkfAx9upp/3c3wQl1iIr/s+wI33E/Nbnul4d7GQxkEC1QQb9bQOhSMGv
PWJlcE5TUwIoEmC/OrtjoYiAzqLvzfvWdMKY9WT5WW6/Q6CgWIox/7WcMbY7iIqslN8VmHDOYuOc
jgQsELh4FWwvd2OikZ6m0aYM29xZb0ZYxSy82vQI6o/s5bXxrhJeYZwIblioeOxiYFi67ykwDJdU
wFUlbp9x8wBsLdLb9vyDUlyA8LbHRyIqMnKAlOR8DFUK6oRp+tjJl7LW0/1IdYP8tSV1op0n425I
fQsI3AATLzuEXRW0O2TZrwZ7FcvW1bH3lsL0NxfFigymJC5CEpuTTxUFWKS6n/bR1w/g0nUdC4ji
R4USuZEJ/EyZSRDQ6XJZEaJrhZvy7/CckIJjD6qIvXdCZdN/ekqgiDrTL7q/NfV91u9wYZmMCqWU
zSLHG9dTMgVa/aXh7/J9pbl+3q0/HVbGFYk6aq0entMgnT+adrBGmzzPxLmITZsD5zJD+0E1npB0
IuuIp28rxWDpkcmMKTFkLpfO4Xr33UDH3GD61wU0LXf5rcnCFpLuQWkg5yyTfUnMJTDUVMLVThFt
WVNVRf9LuFpTC8onebNQ3PX/+zml4++u4Wel7pA1JZNC4qsd8HipEvDBXbs3h17cqfyI8GpPurb+
vOiFK/0LlYAxSJ/IWrZx4M+OCT742HIaT6T8mxRjlCTmckPisATa/44jbdLbvGoMs7Lj3rzEU0TX
9CNv2iUCSTDzcjsYS0h4PpWiMeUat2rHz2F+OT0I47ixS6yDUwJXU7Uk2puQWPOwpfXUM6EBnpXY
tI8NcvvHReIqBwGK/HYPpft2AB8pe5Kzk0Ul4kBALX1hO9UOG/QuOibqYxessfNh4e+T2fDwRkWo
J8CsA9colNB0lsyOUfkyZTBdwjkJ1ta3mn61oeiTWhYgvNOu46XTSWEQwafr04IeB3iOQkNWYSaG
ZPlvAd6+CtJU+Kl8gMtKUTlfVwjiOevOck5MQkxEhIbMfQj0/WI8tFb1Gv8KLikvDJg+26EglFDp
ACsflJ8ib/qpgORBjY3bjWC69x7YDqs718MVpouLyNweaWPkb+dRlJd5ididmRW9C6VOkSWBC8GP
WgAK+OOcFg1HAloCgI+rtLwgP9Jfjug3clT/JLJJ2zQz39DAC2b3y+eH56RswQCv94Rh90zPqP5n
0kueTJyzf3Br2GknuohRsrzwR0kCChg+DN6Idy/i4TUVl36d1wZemi2hn9QARcjYSzy8hNpYjfP8
DSZD/UernUY3o2tsmRse1nK6nYrUe4due5Bd7b68ezAhfzhELxmCAn3zH/c7FZoeZha7LOYXB0T5
T1lPQsxn5XzI51BRzcRQCfsRnpkJXeKK83n6j9QGbx+Szd9SZY5v26AmYj9bOnJk90B0gfPaP5z0
mf1ckjDzsJquR2jgvQB4bzz22Rl4IRVtVVug2+7upq9cFQ0/9cqD0mRGmxGTlvjoA7S0EtUOQZ6J
Wo8ZAZP/ECYGne4YmGQ8x2xRFI0u7v0V3Yc9L2TduzceNNQqUDdKrycqe/jBRcGCR5a58ykiJVaX
g20+oRqZWTwI41whCaMlqz0gnqiiTNvazDufUQZddK7VRZhLWw8zGXHT/PMuON54gijdqRJyGTwe
KkkGeGzWoMxoAy0rAu5zqGVmIGhLy/bEgjp/MpssoI9MX9goXNobAxy7JZDygsji8QSAbZpROaHN
+Y1mQkv2xC6fhhe2CYMrvx2lF/+M1bqgEGGZPSFqDMZdrFyQHX4ULHUd/ITGAwdoeadLqoKnGUOL
mBAsMYFKNxcQ4DFUrF8m/byJm7o7l5cBnXg0e1Cz4vmsfW4xHp8YieBy+oHDGCB9qBsydSAXL7ob
IggQaOR7fmSxSEaYyFX0/6JbVCezbK1Df3j0An6n57mv/MW9f4iUg1x+C4itm2CY5c5k+dyqlTMA
HDSqXdONRAYbHzbyxpD1bLOo3sLjJXpXhtXc0E/QSL3UiwkuB10FXFN4opY8x6Fhb16JMHvnUHL2
0fAnbNtruRFoemjVBTTPUEvx6LmLzgZjDiecVsC7s/wVk4ssP9wDDIdwBJjeo2i9Ry+qw0YWwMGf
FoYzQLI4+KNlv3boE0agS+vy5Ul6fYKXQztHbKTTHV3H4rH6/XdprBolQo0sJDrjBDpk4/3YTS+M
QcA+mnK2c2pGOu+4TE7zSBOcpRPS73fBJSBsHtDwV6A8WAEshfgxdeKZn1pR4HniALjci+Bt0lht
16d4Hr8dw1ys7ACIe3JWbLZXVtisn2+6vjYjyyT9J8nC5a+UkSmQ2ehqu81W2On6pjNFjUudw1eX
P1LkE2e6Mo11ckTjRR/pK8hcCQQgtU0LHWJb0ANzIcrchH5JhQ601av0IgiqOFglVqT6p/gDYFRX
3S+0I76OgpN+QJ3HQvWS9LzF90c1yrb0sieEkNfTMu5faWzoZ9w+Os1emyg4UP+aIEmcJcvbhkI+
zqIGOc3T0Ac69Q6gcPCmgCsmS7Mv4MnALKyw6xNZxeIcChff0buK/Rdus9q+c6rl5Ng4YRiMmYt0
Z0nTi6W6MBsaZJc6UDHGbmtx8nSLydVSm7bm8FNHIs++VJUxCrZHdsBlP1PqZ2IRE8e9DSmKZZ1O
ltLiljXaA3Q+vhprAQs2Ksui0gTiXLs4wBecEzE5YbsYXowu7/AJQkN8MKpcDLScZs9PEpk9dpz7
7agywHsFCWChphSavfhl1r6K4c6OY0KaF8JcG5NlFpx+bJaziIlhxknZNEbfkbMPxTJuoVYyCmRQ
PIj5ihmn3anVq8d+lfNoEvGCNuqcVZM77e4QhZmXjEEW25IBqTkCarDhQurXSAR1wJ8GNhBmO+5s
xrWgdQ5Pj2b4T+xlbLpFcRXSwHjwhjvTt1C8YSumJgaoW3/xJK3J50kkXwDywP3PKajaKHFl6QUf
vZgktdWZPZss1SSA73f7McgEFxDs34h7T9hUA35rb4eDJClLYBmeavZCMe6iwMipkYO7S42JQEsx
HdCjNuYh/q9WlaYodtqdpRfH+lt7cjBIhQ0iqVslp6wx9+hHswAINp7Aq4R+KcH6LL3IXZWTZZTZ
LPlfytdo9UZpmkvBVzarTPXSKDbwrrrryVRSZiUWA/RfxvWvG2mJpg00+9Y/8FoMcUknJi6t8rXB
mxubTjPCScwQHu+4gea9CstQlDz7Op1ZXQeTYzWDDKhV8brtVA81NORebE4aWqM9toFArF5racG3
JjXtCEtp9fTVj1A9t9dMo+64rYUVSAMLbIiZDzUWkLLOeMzjyUUdfk1PBPwEVP/8PqX3SG+Jf9B1
4bI4iEps8i3RxqvtZiswFJQ/Sl0Lo7ntS4sIC1gsdyACKIdEbODGdn64Tqia5fnYMRJL48iwMID3
TkgBjpLhLZVMOiF89p4RSZma40wNoDDsT6LgLJ13ps9n4K2quobZ0tbwHw+3z5pAeS832s21MBhJ
9kp1MQfhL1wRfuXE37XfAEO9G8F4kAGzVvbu2Xw+rsQX05mXyE7LYcZyp14FsZzx/BslQoVoGR0C
mR648b3VGsN5iX4OK/+B94meOXuYEkmZIr3/DK2Uytrd9OsLpRechiqN4mNNAGsrKZ2UNL4YEUY4
XaYQX10SoQHRIlOq/ydmurX9PdB2O/p6gXUHhfd+K9GI7mPHZvkaysZiO47LzxSq3bsX/xV1yTHs
ONUxC9yRUaBM66oDPSG2eerTGZC5ojalnEGjd3f2lpjbWb4WvyoZrNHmNuP0zWBgssZcvcC1c89J
mW7xDGqP2eclrwlBbu37uJ1y3+HxhQPDXGeIIy0f/BzvlFjnKQduRM5PsS87Mye1NIO3raZEe3SY
v3GRaib0LkiIkTBiWuaUifLzFdS6RdiAbBsmJmlOW3xGUiYrBZarpFhCuJgxfY8gQfB/DNhb4Ewj
cAGh279/h/6dyZ69Luml0rUrgLNLr5rnHQkU+xlwsdb2THD78v8V6Q2PX3xyGh3XBKaqYlwCT9JR
QBAMwnoI6ivIc8Neb3/U5DNztSayOCHwuv9v+Yg3zSkbei3Smj8Q0QjDJN0QdO0UgGrfcGKwnGD8
LeNz2BkI4XQkfDQ/i/1GcY5fysycxEV7AJnXikXCR5nUOGaqcImn5A+zhzp5SFzLdrGvOubDEGe3
I9uwyPIo+DJruYoDz03O4lO+OQ/Cv+A1wTXohd9QOvAuuwsDdeA8o9F9/eiZ9XINXC5+8ADCD6vn
W7iMU4XKSiRmP2R9pC2fiJLvEGDdCEYn+QWZ9n0WojyDowqDLawR5jXEKf8bGkGWG9XEmatqv1eq
H3TEDYEQyRJxYpKDfzKhZGy1qzEAHDfC30CyAXizuunrOVaDdZnfACn5s6VmeNQvqfNk2Q5mY7GB
3Nz6I1BfvuiceR590i/4yaOqN4VUD5Eyrcxr77iTlSnwoa50IvPVUhxgZynAX0aPeQLt9fzv7NDB
gDeMgau9vGWmnMo+VTFrByxI03piEDxgTKOgG3lhY+e3I+ccKmmykthMLoZfeUTQE3GC6lDAepF5
dnP7IUKUo/OJ9KyL3m3rMNFqRtmmpA5B5pBczaZvjha2o5eb/rRzXL+i59yjDg18K9wimhq8VB7q
hZzotoojo3kIy+DsrqjwRVBrlmkJkaQmq6T4QC7hN2Pa+/WqBk4Poxysxq/XFlKJcX6AJEBJH8yx
cUwBdtjTihNuAk7i/kG5BdidEhgo2tstvrUtcufd+Dvt1ctfk6OC1bHqsa6NPRdbkd6WNfvdU5sn
Kpoor/L7VXSXHDFbmulyCSGEAB1JD01gJFgbF0TvulSdQNwH0h75IYNkrXN8LV00QRjgLMeR5UFQ
FMwHa2eupNsvpcHdx83vpvuq/aJSksw28DaalNM1LaE4RvGN4FuwyN2XjF7sZzBfJnimoETmHfA/
+vGGcZ1rijQtO1Q4tVdxWyLqjyJYJTsF9cT3dc/8EYww01cYs658mwJrZKIEVVxHemL1XP/fWy/r
HYx2V6qgvHeWGvKG+C4nvYGovbb7fUaGQCLV/6XrfdLyK3/UF8TX0U1W3r/dtOPDV1uDo9rSa4Iw
JZLxf/ZNLlb/fJTSy8IUGSKp6h+rqt1aEBse4tCGsuOX3uNkZdax66rdCLSLbDqq9/Trcd0xZY8r
gkMzyFh08G6eVKCZX1Eok+oyUiv3H9qiXHrdyC5wytS0V/Re2AmrDaYCd0M1BbcrcOtEqcI4byXZ
SydAxAKETHdZ929UrG4UWSP0j63+eZm3syVA0jzMQYzbjtozcIfxwGs1xER9NGuEhxoDm3tMGecU
61RsZostkpVRQhHExbwYy1324QWFSAy4qyEBBvn1PVtryUKpWwgSOSauKqLocSDP50Nx6Y61EwCt
eP2X9ChzhbcCx94v2pVFcL66LfyyOoViRzvqOcIRDTD5Wz7h5Y5bXPlDnEVU3cGKiMCBau5zj1dm
V22uCWlMPdknfUA6yyrmhBa+j2iANeJ+isxgz5FZUVMeG5rHSa1umN3fS91mTo4/iyq/SdG8+uSx
PSUAciKtj2V8FM20zmaZmFdD4/GSnd8mokD0VR0AS8uwwyUSmqivfsHvHnw7+b6Ax88Ub8PxaJ6j
q7DWGAy/lYVLC+7+CWAM5m6dV3AIzsC8Zy4j7NgxxYwp/uuTNq2RPnbQau1AiTQI+GC8srF7FcXY
eiJpw/koHThkY9FVMGoTy3ozh7a1MrsGsgSmAO8ycdaSMMgKlTreEz1E/M5jwcXPfXnmTq78yNX6
yAqkc+b2QPB/No/PWG0akCBIHtArzBsb9v0AWnK0/i2fGM5+dBcHM7OLjmcQ73rc3iK1u63FIymT
aXV6R0OmIIGAM5G8Ektc0dSZVYEhJd84id0Ws6dhe2KplUCIaC+kyLgBdohWwozJMWyLTkM/K33M
qLHlEat3cJ438FD0m3fA3yq8tYuDOZNhTU9HoScVIQDig/UjBWXX0hhX1t1pOV2ui6wSYQIsi8nx
kIdjG3gdw9Y5XdDBqnOb2iOlikEuIXBmUXfVJt9oiOa6CcoDy0qhT5Jwt49pCH99n2oW8ew5pULi
iSYRkh+j5MYuRwtbXICKPyEYt9vLavKKKobOuO6of1b9351ycnfl3UDYCngsPBr75DKHBkLm3Fsq
H9UIbhqk5BG4ktcCKqyMsusnDflDOYhqKSokkhOb/8vyZ6bMSr1wiOwaL0j4V+I7G9RDg56f0uux
738dEBmQG5fOB1xi7Mdt1EEa0xohnifEZR0V0MPI4T0AhpirCdR1fa+Kzk1iachLRIJK+dLAXScY
PENxo2DJY33TzpRXpJpVXapftr7e4lsSuW7hWrjdJWAXPqqPufyXiCmZ/QrBb2Syy9oi9pv+ez0c
6a1ThNWfHsicAMLzwFgq7HXRhe2tyYxs3TJMJvQnUsqRYt75Eav/Kk/9Kx6rz+YKgTKJ4VkuEVQV
J14FjcauiHDf+98JXhd+3K9uJJZyNrhz2ZIP/j5pDfDZyyJmqb4BRi1XNwTx39cDDOZ3SqGMntHm
dMqcBPpXUxSymzA4gyfkOm7QxuAnaf99lZBo+yCA7m86zHHpXUiCUBHvx6yfLiKGQEl+Pak+Zjh5
inrP8kXBSGWy430z4id0WcsAT2iqCuAX0aIEWWSnc/49TKSHtMX/91f3nK2Oy0Znb4e8W7DcaDG4
5h7SpF398DnJdtrfbK8Ig2Afu1L6nZZBOeWkI9a7WiPP79aFpW+zCqPDvgV36WuM3R+RoxwCuY8u
UHAH0Np7IBoAimeDSe6MBZ0uzDq8dp3jHEV8wg9NxL9bZYpBsk7Me9Dzz6AtcJN2Rd7Hc5dqrxFy
uQmYKY5JSuGFp0cwj940QZLwCyBea3O6jT/C7MBgXR/Hnd079EofJ1NQOQuxxi0v0KogcHGXBtqL
yNF6EvKJ5bWGB9S7ZthJwMYYqRyGbCUxwjq2IOvH6TD8nZwwdyM5g+JIJGR+hh072jfk53VZw+LZ
jt7FC7QnKDH/LxYJYsOiK5io+bsvdk+SRQPG4NtAf3odJc46FUQs1/femCpnjZOd/XJfRX/NAoWg
tXp5jcQifkARwPIMNqGKu6GhLFZteyj081xqeyn89B9fwo5GhYJf5Cp/IQJKzS3WEzcbY0I/koU5
T2P0sg2RfG9rrLLmTBzcAUIWBVFJESiKi8m23EKflvEt3fmOOj70Yoirg8sVpq5JHjEVOWaT3+Mp
eVu6RE6eD0jtzIThNNqmZOsK+HxRrG6s7dnY1M+6OirQ5s2Y4yxZ1YiocM2RnmzpZTboSoiKH+Z7
QzGpRODnFVUUjPhAXBNMmEuu+d5cUJKlUfgD/ZQkEP2gUQxt3zkLzLUCUnII+Rx3Y5OfRyPjVcyU
vCqIrI3DyKcPwTP0OvWi87Q+KdmLqjAHsxhBUTBfqbxNJ2QJAs6/AINILEC/8s5AJXeDDwcT53O0
Wsg8h6wEVZ8x16tGi8vjrXwYhmp0/7xOqe6bUEtHQDW0Myrad/iddSeBWk1TJiu1xflWikgiEC+o
KnLn+Ojlu4RRr+8AEeOwXSRC3xTQocmldfoK2OX5J9DgEeapRcysEvXPey0Gxuld0G8iCsWezBMZ
aEkflR6qHIf2aAL/9/UJS7DtJFfW2A/i4zXGQ9xt7lH4ixvljwC6sV01Y1P2QkqGVx1UXdg9qJMH
aD2AMrqXOuuFtHVTRLK8RZ5pq2E1P0PQje21yu+YnQTsGDNQg2uygBLkAc91ID3AFuXGyT1brT2C
kJ74j+WW+CejCXzWQ8JeeVltSVfapygx1/KF/n0nDSoJV3odVuvlr8uIt3l8BvLK+O/eFCGQvclk
7b/BNOGpVg55ih0OdQxdstehZ/4YXGEmj1YospuhvX8egLasm4Fhjg59zw+F+9+mdwvvJOn5+5Da
u4Voe7rgjg94BLpdi62cpJx3EnsEAbpgpB1OcSpkAXFfCNfgYxQwBw20qM4Qee6yQzR+uhMjp2ce
kFaaJwakPSkf7oBu3QkYQx3HA1I54IXHWJzNlWjYKibaZaVVLCMDjT6dTxeg1qSTETYLN1aBq7Pk
8S1/WSADKmmywsLHzIYqSMFYgHsOjONcNBpaWomp0UwsQRjjKwG8eyGUnA0NwCx0NNLq8ArgOZI0
YqCli/IbLKqny2jRt5Ph4NnyQ2TeFlX0A2kk7Q+qKeoSQW90WEV5fZKvsDKaGgR4l/wtCjY7rwo2
9QVIZ19Y6cq1i1ZW4KQLhHOs6/4QhZueDZMpWfqAc/PAFQJx0SLHdtk4OpyoFcoN80vl96dM8NYS
jQiXrgDYudN0AMwjSHDPuR8KBt4qm2fil+26WntQjjfvFzcXIVDXlaMoUdoChjp2ew8x48zPFaTY
4VmOhRsCZuYuqKN7FUUYxrWutH2WHjabQtsg1R9atM+5S5UTwTKuOe+SJ6WSqOcSVv5FJwpLeoXd
D4CjCHNc4sVH+e+eF3G3SS3E/Q5Mq2Cc3yWK9KWEIbMbOwwFUXB6i761tEkvJuD2dNVHt9R29paK
TulRtEMWdiaiTQ5txIn5E/qfIP7T3mwhITkMbydY/Nu+8K4f7w+66yz6JNWuqc0wyiDhlE4iPiZG
yGB4/DOAndRD3HVxH9T8XL0NN54sJ/jyrAYoenf79j06XdeE0OqHYCmrS9zVd4naLHbk9SfE3qNJ
Dv0nYLSqTAHC2oY7u6LIoGlyFO1V6HTeL4gvtTzB4HNbhX/uzJaj8lTci5SZPlB7uxKB59Kn1qce
pFoCRQLRUGzZB5Bj62tZPlGjs3bYTpoReYYOAt+/1BgAzirw8tI+iU91XRTA0v4p2r4lSzStrj1p
plcPbiMB7f8sUyYsDkMVjBctjgC9UTD5jI2DhPNtPnTRVaecFgJ5puiHraCm3DYdVCaFaXPV5Bt9
lYbTgZ4RFOLUGVXhJm6ow99VSy9Ln5Km54ss2PNOhDofNk3I5nTqmoaaMVjb8hUYLtu/HW9hYWqA
3563dwnh7Y3XMzrgxzSJvB3fo1v50BaM8rPpER9SmoGBejK01C/S+wXzOzQwhgERAfNMpzDRnL1A
rtoeZIYTltWtNEP1DWOx2zxKru2aGKK7f/hPe0tAIFgYzGth/QruAGyGFhLIdkg+gGWnDa6RIXJX
hxlAALMZ8l4Im3ZaEatO8xEmrexAvcW342SiyKiL9LrRiXHy0j5jUqwRr4zVPwo/A7WuMLLDN7M1
/Vsjz+NY5pkDnMYJfzOnihmB6MF+kFsIEHFwoUgACPsnroNSTIfatl4LobVhPeF3p58Tu+W/A9Zr
YDvZDpHKtCQSbsrnRiVhI/tmUnrC9ld0mTWqjM7a4WMsGl2+dMVdTMvoa8O68MV3bLOzqZ40J7Tx
vcoEIvxh9wUeJo7ePR9iwMHGkBm1kmzShT+pxymlUsBotHH8hBgwjYaF7vesUTG91axmQz2Y2YX/
0pF7ycarT70q6iqbnWpTj7nyl8TKcaOgGx2C0Hvlza//k7KBjsDe887NVW9g1Z8ht7iyWmFI5xBW
GYWvb/tMWdQ9atC8nl/RKu+6olmAoigehqTlxM3PQxSDo8Crbw3VrpTKm7ODckH8XgFVKBWjEll/
+R7ILJ6Pk7ZjZoUrET1mYkS+EOlHCePIiI95dFfoixprfAHrIj8MgTtvgj2sCKwLi5AflN4S5OPb
VEqWUtdcY3fKuNWwh1qsj7GHnlC+jshLCuHw/PWAMls83FYl8jrheOsk63e1t9QsAx2lgBa7PW7j
AEFo0K3kkiIXH6zzmmC/bXEbGWrkxgoCtoayuxp2E31CcencZ8kPgNc8aO8MdHYy2iOuGJ2uiSbd
5RHjex5WmrJAJ2lNf32zS1iylkZWkmkJ8JPmoETvIu3cPxb3knhZb8xfmkdyeySmaRikxYJ81d2U
8dSl4jx5k/pBh/6FiEMMzNI6chUZ8RVeUsIBDVvl5vBQRr3n9A7pLFJFB8pdp/KZeUtqOkh/MwAb
SmKpY/4/biSIEgHoR/RnA/ddRlKJVyFZtWSW+sCI2WHOOUHBd+2LKXl6Hzl1JX7C19rYMj4mXdjn
nuGgvG1nO7e81EtRLe525KLD11W4fVOn80N4XFvCpjRoBzTUEGYwJ70swdFSU2nR83nakyBSPZHo
cs8Qki0N4YPGRK/6M4/QQwJxAzAYw7+2EjipsOhmKB395FhzhnHMoo5jJkfAxkawdfOjJaxjKIJN
k/cJ98AR2LpDe7fo3soxwqO1uTK0C2rsr4SDXOxJ1DkkEwAagjnlk0G8lAdsdfpCl00ZQ3nRFJeC
sjIEEv5B7NJR7abOgygigwfaZ34cYAxQMpbv5reM0ydk3EXEPaaHDWyqys3DmN7UOQGMBV9F8WHU
xp2EKHeuFkIjkJReCYacJlB8hFRaLnbke8I+oKJVy2FB/7snmlbjfg3LC5u/HFEDjYkPiu/lbysx
dIiESVrKscOU0lvTdgfJ8qq1Aow9wcY/PkP8zN9qyoo6fLD7y2NLVTcsiRo0Ol0CVqWBH0FuagSW
/HUfm8p42CIGqoK7+1iaSxG9FWIaHt7G6Wa8MJxY/5aqGDDDBK5YIcJM99201ozKmNsnJkWvuUc7
opCFMXSDL6OOFuq/PtrPvc4H2TG9EW98yTgEnoapaL1244BsACsQ6ofdo9Woobxv/clkR+i2cV9K
Lomo77XC0DMgkgn3w8mmqKC7ZKJm1c2m1SKIez/3b0X8xEIQdi1JPuUDT1JhxW5nPBdLX3Z4tfx/
Q2I+a6okm6ytnWFvKpTZYTfsPRgTR0bNXKLDR1UcXvmc/da1nCQ/mRAaay9Evs/MPfBoIz5ZVZx4
qGuXwmyrCbCTTdsoGpmMd7hIc2fGb39souakwEAb9fljzuUU5ExDHLc2nF1nTlUVSQdHqos+Tk03
tVF/5i7nzsUI7IhfFh6FYgS4gcO6JA/bvRJebdpi56RVCiVPmEinxD2OXpqzpWv2TPCDdXkjS9L1
VTItmHYv2k25bQ1Yp8E+yr4LSoqkPY2abdC/y4yaAc5Jt9HDf5BYwdN93YB0bxVZ5HQS3SP49/xA
iOKTbcvad6EZB5Rt1ZsBdLmgEfexE5NxJ6OaIXZ/Acw8wwHoGQEqKoisQaD2Oe4uh/MiB0QFQO2M
slHw6ddqnu5gHmHEZNmUE4ySCQu2udrjuvSiwj3b63IAazpBu+LJ74LuSkKznRJ99ZgKy8tq9jPb
vaR3R1BCi5V2Byl0DG2vP5RfIOuXwweu/c+Jy9KnivjAyvcr+XMVVpTvUPjGVN7gEW92bK1knoR9
ebHKwZMdgWe8qxnM0crjCDgDAyz6trqFTECfIt3WbKieMl3KTB7MCKHp98wBMeSOvtzJ6mZ42AS4
XfsUvbbprpkDxMa/Z9Vf0bU8JK5t7ftm8a5zmR6bvFaqgG9c1oRQbecdzNuzrdD4LYJ3znMn2RhS
rOKJhvTLMWIqKvWiU3qJ2BSHW1WuaM/jB6CvZW84s5kENmCFR6ZuBAcwnZdh0gcL8hz0a3MH65Gl
SFydOzD1K+69FWDnTBLvPiJQ4M5n7ZR7A2++Q/jAT98jtXNM8aUif47AEOnF2Drl+bBX8CehuztF
cAM7+2n7Jkc4o0L58e5VkP5ejssd4iEQorme7sG3TrLILXz8+Eh6pwWA+UD6Cu2lJiz1SBvcfrdb
oMMWAaT/3dtFCyOrGAChKTH5oZzuHuVpRsEQ86PkskIenL/UNmWBO58p2O32DEOMk+3KmgFq/3zY
vx77JbPiHQsHRV/15ZznmA5QVXVdRtxf8z7S8idCIf+y9OVzpR+xLsr3/Dsk4qEeilShmk9MZjNo
ppdGZlxmB7UIj+qumSSZDiYpG2VUeUH/HNiyHUN1afTcXMOWMgPTppbh74MkB3j2aJuTGD849dVg
SIGT9JFlDVu2XdSFyvFT92hzRK09w1YA3ZtH9SbPKz/+9W9DSebtWlx1iM3ald3uIh88syJRWMvh
sT0m1sxmAGeCzU4a32IWZxfAFFw7pVqxmCBLWlPYzUN7FBFTOVyqHC4mza9sd15iCchccmw6vTwU
a2gDp5o5ewKV53eKJWINqQms3ic78inRJu5mjQi4evoSf1kCNTAG6UncpaYasAoBNwXGZSddXQ5o
3/PGAU19rQP1DChKW5wQcrzdtxo0lIkRHgk1HfXivr4c47q4JVmwI2t+cEh7olHLY2ukmmWTnJ7d
vY0gFes8tsDmYYyeqEYzSr49dGM12lnx9pAiDVlz9IH5CMRODvotat/w5Dj/rXIQXno4uOAn7tZE
v/xwqMyIGkfhWYww+KksYzhOMNqthbck8WpRn/xATBdI0uSjM+A92wM571VnDkxy9KMB+Bswir8P
lUZ0lsZaxoLK8zasUCPvEMdv628ggaRwE2VKlnixLwbkWxGp7QbiA3KjRIFME3aFRBkzwe8JlTMh
XlbG0/LwkI7EPFcOoc9EQXQ3+Ps1TqtyAoxPZfWeMuAEaJJRSx4YvUewGOtj0WmyY/xl6+JqlXmp
kDbhrRDMgTwjuvfNVOkrV6AsE1fu3khk8FoZxDc6J3CHBhVmGqq98N8XrUnQ3vJRYrew7lWkMfG+
u/j8Rh7/npASJZXPTGT9DZPjxiuRHbrYLAZddyngBTUi8DHftWIlIuF9lmwsTiUmWjfkzjrzZU/z
BkPZ/yFgFC/AwkJCRDZtdxQXap+Y433tLYmiZDzjNJfVqxpwUzDCk48L3xqO3D7loYdCvZKgip4X
Rpk4b8Rsnd6ly77JUtr9L0r6W9oAQDcNYGucmL9DKckLF3PI9+XH4kF+JlVXMqT+6lDnbak4xRKD
kAb4aMhhjmB5PnFZBIob+sIApWCH36xtqn1oW1RJW/FH85fTOBCpPxp5dqw27IkYGRokrPR+HOxR
mlOPh5m/lsfDap6ZpK65DuLxGwyN27grpAw2TySNNEw48KcwxVd9EaX7y2trYe9OdfBvDGU8gIFB
4DvONYzo88b2XqTF+prGkHLDp78iId3wjPELYjy42fNs4PNkuV2BDsZA0li5kNEsmOuh9fiuH2KO
xbyP2kxpRsQpveKhUyHm5kI3fyDhaClgXAW+r6H+EV77nF7FC8TAUOHgxUEV6cPt+EgYMTcuvUst
zb1yz75pIUrmMNaOCHywrOFQowRecNf6mCqKkDkN9LxoL4uER6lOTA0IJMkw9O7xkQ6EUPFPNnvy
MDhk97G/t6KXdYLKUBbo4dL0jy8c9+rlTgbcli4BV8Ejp+Wcpa/KlBODHVyNn3QzHAoELsyVUzQq
L8dDApZZVScwbq/4pPB8+s5q6XMiQT3UraCHRWIw3LwhowOpCT6VoQxIVwDh3MahY3qt/AXoGCf4
NiO/GHCDPW5cuuM9eUscVsuojwK5BHqE4jWTMlAg0Drz8xvBO+q3TtOCTiAr1ie1474qgOo1mkm8
t8Y+D/5dCWYU8V5ILjZNpIa7AR8bEFHp6SKtneN/ZsUIS66E+S9xz1u64o6kUKV1tcOHFIzm479T
jeZu0WXzzOdBh8OoTG4k2HBvWF9n2l7D/ksRcvjDuYsIgVfgQJMnc97TrhuoJm8ht48nDzc1kxwn
pLfXJqJLWoDRM0L8WLc7Z+VwM1XQ28tbU+TZB1LOq0wIqrEAnEoO7vEDwtbNM7xLGLWJ6D+wXMno
tF6MsbAycdLZiDLXfXylbGxTPRDRF8wcbXy133URTRBqf6OcTDuEBzW5pVc3KNb/+pbNAgC3rSHE
zdHPy1YN2WAQlcCM2Mc8I6WDdR+ZDk42jD/ZGzv35Rax+o97Kp4eJ1hbh06Lo5lk02CrAEI+aopw
1Ex05OLHpaldXqOh43xo0qGDauP3XFcqB5ZMQzTXjk4uCCr7WwDKfKaMqI2uwaNdByp7xPbY4K19
tGSsM7rvNnHeObVpJ8dlHehD5fhdtfbCdOfnnUIgq6IQ/DkDQDT9Iw5RFrcgLtZh0luIWMq0d3CK
eZ9IrOg16SnEojMvlilZxxtId0619KbzRDC23shj/f2gAIqwIpQm8m3nGORg30AGBGjpKvQUM/FH
nb6BVLnuK9DVpHXzVE7MTX5wrwEEO3VAMoYK1H0iMg0sUDY2IUcfeA9gpxq0tyL0LXaUda49kYrC
AVUEdMIAsZtxoZp9XRY9uU79OIxYCl63VwvYOOygMd6VlvtA3CExHu4mM35mffGIPHzimiF50ibi
IpqfJihaD31oO6F/CX3gBLrfItNhERbQsLIDmuNy5gcWWgPa0f/yZrQiTjfFiPPSLqvPpWRH1K3Z
BUf+gJ+9Zi4WZ89H76xFBaZ3M2rhwkvzBGw/J57O9urNMMg3vp5fcFjVObqbUglc6FJ3/19Vp9Ui
FDlhLIvYsg6UP4KCWBwCkcOdy8HUclRqkc1jaeAu4Gi177/V8391uR8te5qB/GsM+4TAeTCwl68t
Fm+1NAnddkrs5Wicj+tTIhs4JAg6Ry6HxL/aPEnJ5lI9RfuyZosdeZN8beTKZbvMCRUTwfwK4PxA
68nPqTs1YWqK+3YPl+2GEmcro9cZG/SRychac/z1M0hbMFLqy3bmediE5HJjdHLnoBLvL1Go44lb
Uqv40zmuxP817TGoUy9ISai3jehvDdqKPVPQelHKEnlfKlERQXOQjJqEFYvIuyZPMGOHfxjlHLxn
xP3e4M9RSHaIMKYBwqEg8dQsNoBk7nhBuGrppNUBmAF7WWhsE8gMz4X7Sqs0bq92IqoaVVhWtzle
WdjbL/+Sl3rNymb+tmsg5qaQLE7do2loGNYL+cdWnDJz159yYn9Adnf1ls6qG1O/MERz45AxtIkD
A0fALORcTV089CCh0LQJAchAvq6OvCp0K6VUr5E/180ROulYbInRgcGmfCXB7VezdZ45J6PKXF9L
T9izjtsBL+mHgVScJQmIl8m3bruf/Ev8Ggn8Ht8crDe/jeb0v2KU9F7UHyMCzO2zElBluX2S0l4g
dIxhWTp+SboxCfF9U35VWCWIsOiIWRfLY3hCYlcZFjhmhXupffK7qT0fJo5kCILzCvD24C3KJ2Tp
w/bU9EV7X1z4cE0RNKGe2AVtvUXwMuSxJIaSKgBNQNgGOg5XF/49hRVKR4lc+QSkjXAdlvyWjSvx
lnndIET/TIuuvnqMDErjGrAfcSjRQROnHABZLyymGEmXYzslH3tlc5JGbBEfHgRSyxLdoVU70i4t
4xeseM7Xaz/NElLsTtW5lThG0XyUp5D5pXwUOurGbVey8VpA1azHe8bW5g2ewpiYrQVAnyg4NnkX
HM1MlclErng0Wy6RpkfMZPdRUPEtUUSXPlEIXp8AjoEji4N5eBqFmc1cLlWEymyt9DnT4tdHAMz9
Sr1hFBhRtTVyBJikrjrIojfip0XJEUE5Kz53Uen2vKMSzrjXd+SXx3TY6Vsgj2VecnvD1PW8PfkC
e22j4DR/A2xNFH+1qlAaH2hTF2LH9b9i3RCaoMlXcSThgyJXKJht0P7H3Kt+4XHpfvXWrMo4En1h
begRZPDzx7NodTKEHK0OuAyOlD4uguvZL8w6xHgcLer29tzEReEN3YKP1IuskpggNH9kqLcstJSR
u+va2HAAkUbYrevdSlie5/E/Sp/+mcjgu0g/Iv2PK3szF0FVUYs/SuG1QgyiyClIoo/FIQ8uKX1T
p+ZrwiVaioFQy1490ZLV5tZyy5NCyrOP/Nh/CbCNckMznkZNQSxjnqYDypyqRnsEm5NTpAd+Er86
qW+hfGJuYIUWlZQlO7gVSK5TmKMZhNofcPWVjCjjrqTZg6E/QnqbMUsub2spKD3EGICtPwsLh0q2
9EX7g/Mt6pItLLhd8Ocm2sETS7mwtjSV9NgQrBRZ2eRjypEl4KP5MJjs/sfsFMHR3HFnswlt3BqX
NCoGlZq7T4w3hnQaZVr6WeXm8SoySl8VWzUK/LblqACONO8rXSfpM4FYsogNFFUm5x8Qo7s8dBcp
KN968c3dvGhumOtLDcTs4uLLx41XiKKGAq7Oxi7H2hwfg4qsSfKCYr1UqTMYfc0AFSF9VOOppBzC
yKXTqhrORx/FGYvcEcB/llaujJ3k/Iyad4o2ibTpX/ukr1QLoPE/u47qCypLT73CmCNzed5alBLv
oGFCmOXQIZaZREc0xD94Q3QiAEWg8RSnoSJFXTwTHFAj/cqX2LJta+Yn1GQKGQNMs18lHg5MDTsM
ZwcTGR52zkUhhLWdJ6VsJplxg+M6Af+pvXJ8ipbbssh9PYrFE+g538IOR+p9VznIOYzoHJJmj/z5
hpEYe6sCSZKzYGZRhUsDLxbo6PdXTVSypM9xrB8Z/Xv0FpfV6WVgskMQYIcGdUfkB5hErEBic2Gy
9n4FuOVWeRnzasyDGbDrcM5SREkqhniCwOM8jH2cx6pWoJ3B95QiPSS2gCFLUDwh0yeEhGWvuhzm
tEz/T0VysnRd63lKIHfc5AcwnmNXONw5/WPRcVAlgA35sdlQbYzVJCcG7+R8JFdnEzgH7JbwiB06
4GMdY4IM65NhFo8XSNzXRgeYpJmbok/0xrRLHUFRxbVSCNXht7h7enyrvzk++ps9hcauVOZOjsSk
dgLvBdGuHls1NMfz1XKyTrWnEdgeQi6sdTNWSgKwcQF2wpX729Z/nw89oR5cLk5mTQ6Y3DqRatnB
r+YUeIJAnyJN0JvQoGF/sIWplXZt+CJxp2vGWJuoGkK8OKVw4nIwnhj5vh1gP0NAJrDZ0ZVfxTX9
cZe+0euwIpmeM+muewBLGAvR5GLvjL6vcGtqRW5ppP/z3kh2r9DybDqOQ/vxQpdzOrWCisnhIBIb
yUj91uliE274q0QKApndhcWp6/0bn4JhRXs9O/UD0uTQ0Uz53d7kPEsbfD4wGKGZiLlpeVlql6Qc
5sFY4VFxEmT+cKfU49tr8wV6VASPl8IB0MKaonxR+vSkR9bTzaGO/mYw9RxzWiYq92dhaZs9PZm/
GgbhXZgFIkgVpbKgvtAJpesnRU9LahxnS6tRc+sWGoeukCVQNYJJYsRXBf9F3vPAL6uqlxVaptAN
0gvYEmO154Fnl6F0p+lwhzduZ7iFK4FgqYoKlGmTFX0+2of24ZJ15a2NmULMfccDvldiSOMQsMDo
fIFVGaQtvj2M2A+PCKBOI0N6PM4FbpVcWVE9/01dJwaDwFOdd92OQ/M+s8UXeBc87w/nZ2VZqfRm
ZckHf9C3r4LinyIMjWei9CwXshK7tHq02JUSBpNUELdx18Qmj5nLT5cPjPma+2cXVFlS2dXheAVX
0NUfVj54IVY+UL/QM1G8iXD//Err59BnKzxRrQUOZuMm7w4RJKKLOrxSkhPoii8OyhrMFSAt0Asy
Tyc+h0QXgcrSP509UFerd1MaKliYXpHlG3e3ikJL7C0FJlJqB8lStMObJz8MJ7HMV/wpQOe+xHS8
HDcda516AL7OcOo9mT8uX4BMxEQF+AY3ABy5F3+pMP48gg+sgRJzzK0VQQJ14XjWRjLjGu7rGn71
2i8AvzeozAoEDFhgT+ezET9oFlUZn++4NLwdPGjMkzw009MLI4PwLgyalGzK438bmfducpEFfF3v
srVfIG79bHQGphYIi7EJZ9YkIa4VerGv4L7FGOXl1MumWPcJZPtOhlei9qZUFZ04LCxaLqGTCJ1B
qjpNIOBM0fKKUM7xrD+8XAc9vmzKE3XYKHt+8aBsYuXc2DEi60sTbDueQKqEhoAKf1Z3G6Hks3+l
eJnfGS+Q0pBCZeaQyaUvIcjJDMrsYY/Qm0rF1cYN5b57s/M1Hu79/oxNdj++szbiBchHQo11k4cO
uYD8cxJA7i1OAbU7iraXVGUnKCW7BDLjsqEBMM3bQ/xagiftGxiX57qptKX6rAOSwReeM/IVMdRA
b+w7Y+1/+ez3344bYzP0phcCEZoEdYd4E6d2LtlU+9QODk5zimqI8KmPf981CVW9kS451v4Do6yI
9Tf8kjd93SUS4QFjvZvoI3I76K9rNYSzCAS+s0HD+o4YhiOiAz2XfYdt81VkJvfzJR8flSOcDMqS
qswCbGmW9hT1hsktXAh1YOSk88XXHZhpDmJOFZi0FnX1Kcebp3d2ft0ILWvslQDfLlcg26RdMVvK
U4vzUWIlTdKHvCwsMJcMor7Vde8cBflRiil2CMsyM/ZOB7CcxXVmsxCd19Fv9qELkt0Z8IdAUyN9
dZzg8l7w+4i8LsqGLkXzuGM6g4MP/pWYxtfZ92PJeeTFZdOFXNyI/s9jxGUOEzfp4vLpFMeikUL2
0UTwqC+iWD8cUR1XzRJSEPM8W6TC81CXIA81GqObLdvGXDIaqu0FLixC4OVHyFZT2ITIhC+vkoZy
T38eXQqGrfkclgT4e071MbN68Pod6vcbeMVRDhDOMO+/v/3qVpA9U2BbcWdvc1jlJNZ1i5RcKevZ
OnMfjXowyPmTafJB2Xdlf/H8qR0NHi5NYHmR+3e1ff7KDgpx8Fmns+UbpPPsm07g7qItriKIT447
K8v1pKYHNM2vnrkBtsi9LHQziRtnEpFPEoiOgJimQJaydQYoo1zTmpVl3tnwqry9gGIUdCaB5e7L
NK//BoVl8Sg7XhOsHAx6iprFctYmMa18hqWaLh9jFsI2Hfxsq4tBpn+MSseMKtLynVg5NY7lRkpg
LCOg814ZFTrfXyUKys91AqyzAKXAYri12r1F86p30YEE0ECVkY2FxgWaL4aWg4kcXkSB/L9bBz+1
PxWMj1+2imlJaOr2wNHBmfbjluDLD708dA8BwRCZ4Ztql9oiqs76gFW1cMrGsEccO4S9S4CNizRJ
NXOUyrluGdO0H8w+ork8W4HLODqHnPXhlK0blaJv6EH1EJuX9Tu4dtKRDMcrjqgGNZTdA4EZhcTz
qHs0fk0j6mmT+8vb5cPEZiG4phjzn0zEUMgHt8mkyfUXygGd8lNvs6BBIIMWjd7+MMyH9y3sf5u2
mdpfwpheVrsfh5UG5Wmuntv6VGLjAHJcZs+p6uvCNa983xU1xpT2RRQMWRXuyYYfTvrhgGVUmxb3
FWgn18uG6I82iQD3OkSMl++CctggR/PCrlrJjCJPzASrsRpSZYC+l4E8iZd0MWW/ymMw+4BCK3NF
qoHgZgmu8jMHjHoE80yhv1LgGtbkO651RgZLtsxtnKPND4QYbEhbrW0laL2+7y05rhqfo0AqVhHG
WHIcFveS38my1FrwJF4vNXTFXDI69DBlkrgiGWDUtRahCCL/woeMvOTX7iMNXPxV/6ni3EEywo2k
BpEt00bJzf1cztkVA3yGaetpGliArTLZ+RFJ+kgYPj0Ll9Vcqt4kdkG+jFYARlIICeyF8pA9zglo
VoRtxtxvLScHtetDNg/5u/YmOIHOj1Xdyab6TqZTSUOJw8N0d/vagQVIhSg7WyvzPvAXEMhmtNyO
nuKyZZJoYomMk5ZuxXx+pHeBfrVVW6oEZ9c1lZZYRwHn6N7DU18YEwUENX7tYIvrijsqRov89Lzy
dIKbjXDIKYY1jqWj9y1R7NaTZM88DV4urppYs2vNUS05HsIHrvc+85M9MEVeQk4oyxR92OElaFgJ
CAAnZIibxQR1Nk7qNPZE+NeTFoUAyfseeyoEAM/hWyKW+Xn4B+/cj8g41iy3b6I72AyPhBbc64Ek
vaD5FVhTamMC8yUZlJxoDIVXdjy8pw7Ncq4sAFseUdt73ABMpRBMVntPE1eRzu4tFT9ZvmqK8rvO
pWOjqVHumlIPKykhrPT/OikJ8lrfEtRjHhTZA73NvVMf1wvMkTo8Gfu/j7rkVfyreUEZx46oaHJl
agKEGssaBsR1YkbUjqte21z0FLrJiS3XVjkH4J6bKTkzooEgMEqgD48Hv9wZlNa7/w401tvgIJqq
as+Ydq6Iri3re/ZM1gXiqKjUuEtyirJwfq4P7cKDWYXm4usDeomF84ptIYlBG2k/JRTK/bow2GXi
1rQgIvv5+twtsZBjsAhOz7afVaKcVaQP6rufF1mgKmVh850O+hzGtbMP0UzDfLoZLLiIg3b+S21u
GiFP/xIuz49CCLeOwKhh526H9o3HsoHI/41JemEesLnsEBOpn8HRJu99NW1rn1/roalzjKvvzwz0
UXV7hK/OHqRpGoqU/QWQ3MrYUgOYkxurC4F/a+Z5e8lBM+rUUV8NxOB4H9JsMZ1pzyPXJzCwFhck
zD2gk8cmTAY4a+zbJb2DYeUW3XDEwM5eG6buEuJ0na6W5ctG/UjM5zH/8/iFkVs4nWNHyBCWglUS
+PE+eR0oWcdUEcmZcQnlvPVleBn7C/kmmbPZp3nJxB6f5zHYFCQbCwnQaBeBGrn1wVUKoQ73A/L+
9NGs/hKiSOSQL9v5s9H+lnY6ekv3gH4ycwPfN+iQ1mXvDlMbMqaM6nN1XVGDcCHfAz/NON23Andp
aOjFyWKjaVB/mpy+cPRpTYDrvPm0nCRjjab2+fwUuvaAXp1pI+4o1f7AmZQLno26DtdIEYZvM0bS
Xq36aR7mcQDM/mh24joen6Pld4m2ckN+9S1o+7zKVubx91yeACd68cCx0nhvnheCEvY+l8PeJoBc
/SYsoPay2eFKbAjqGN4LDHV5X1InCwv5jtll2hJ3vzZkjzdwRf2KCPs1gdrJ70Z5iNxnlMKDdGzO
Kv4zwZFJ+XAoBXpcrbQO6OLN53miX0vDEsZh6tvek7TRPEWRSOaomeKhmapBipuSKLOuDnl8WT6y
piGVLgmNk9Qd5iDBxvMfx2ifoGuqfns262Gdzy+vJK5LJtqZk87nJPd/CYusnRHBD6+zoq8DC14p
O0BmYu5g1txuis34thA617ZGJ03GUjkFmouYnCvFiLF210XxNDMfxHIcp5aPdg0ZMsd030fxlAxK
YNtQEnKh6hPlk6xYAOlwoq09+IycpsNYCE6rW+S4zzPEE68h0ehBcl7FHq3Uqke6oesaIVsdg1u8
U9MTZeY1xxnJVX6e0y8nuPoz7QrjLtEnvcT67g8p7ZIP+xCH5gzzzC2XXTjd69ydrjvn0jxDa23v
wx2w12ufoGeg53pV7v647UAxq9LyAaaTqR0gM+pHTnP1oNpncmiQUuKkk559puDHEgRfKqn/Bcyr
ZL3A2a2DChD0zYn6NaRFJKJv1LaVpo6rdSkI5oiu0+0ea5ouSx26fzWgHm/N7rnzxYzwa8bRC6G4
vcF/D+p5Ml4TBZtAUpC4YgEWXAn3hmdvAWiqJKFIAzK2SX5mO7Mdw8IvDf6PvQgvoZ6ilxEEI51U
V2o8w1Xmi20XggjsZzA8hBQfbHZk8DrT6oTBXdPwgwo3MhsKkfZoC+a1a7xRBoQvzMhu4D7G77aa
H4Yy1/IBm1IgtN/8CV8+3gw/isLSgNMjefg95h4GgKLWxnymeKLkUWgzgr4QdfIBdMQN6pS54xZX
+Ylbj+k80mS9zS5GrZbS2NiEf1WVBJRMYZXwUF//sLat2mP1zwWtjKXRdtx4hAZKUW5g93CpsNFr
pz39tGez3mA0IgPYd7e5qzbK5l1sP4hyPk6e4noJCZO+LikZCTmY8NlpdkTFKYFJnR/v6PJx2NG1
VSMnWSD93lS1XW/1qoJ+PEMe0fnIWv08oRxbV6Y1er6/0J02t/PDXjx0uiiXV5bqPkofyY7BJRkE
lYbhyliHFEmdERa+Tco1igMwQ7He46KVke4qP676WV9UIALnFWvJSwoVsQzQ7w7FCnMVxzK7wIr1
jorQn/e2q/SMQXZb6+ruJxBadXRT+PfQwzRG78hwoFtpBZKOTgclAzjARu0efVC9Vsw06m89u9pa
DEgCosxGZV3c5HzL7xtOIZZ42mv28PXgBSy1WTfj9ZuXWTVms2ryLcGQilBv5KvV3qUT/xPVxIps
QAhTyT4jz8jD3LgNe/0QBgetoJtomm4l9o3KSLpdjNdG+dQ4q6UvUwfSBUte1hW6NE1GmKFziRp/
wJo7T8Cmavfpq1t6RYNejDrduVpss4nHlQMFIdqExrA78YxcJgtt/CSz/ZV6trjdbi1Etipe/8Bt
trS81IW5vmXDqQU6ddgpevLqEBg6LxW8LnmQclixU3gBmXnCUdnNmk/BiSFn32XXlm4H2dfy4bDb
r4PUaRBpD6PgFF4sA7wfMLRtpBVBpwXdzUwavixnyS1/JSMTbVY3WZvM2Mc8oMQlVBnsrFRBCKQf
78KBPO5mw6W21HikfxjGx+dQfajNHsoL5C6xXvVsHuIzt5zJMCRKy2HX/dUoPFz1L1gJ7x3eViWx
RG+lCEPkxOHInQe/JPFjwoIXVEnK+nx+HAWhuVUiEP12LNh7ium3i6rGZxZ+OnysYjtf7AK572k0
B7Q1HxQUg+NfeMu4e/52lP+41I48Wa3q+cIFUPph3wcWhcCiArxShv8cbSVrke/AHbX6finPNyD7
L/XUn0+Bj+wEU8Em1kjcnAh17SNPI0lfOVH0aZIdKVqdfb81Wls4MFPJq9mWhdyYAqcF+c/42RYI
HHpwSAVLGMwn27gLMdQJJTJDpB+pMlGQ2s8IFc/ZD78bIyZvhOFSSJ6Sn6h/ogQ1Pgi8KG2+w1mg
K4lSZ6SoUj4DutgWe7epL41rNCKb9EPlUky7Mw7P8JksulC7jr82hws2novqzYfUKDaDPQRmk6MY
BS1sHNEsZQJKOK0Rg/aTONK9IF0hLEnOP+Ypf5mKnEIIKpB3PE3w+XIeLRc3YuXaaVFNa1nx5nLq
pWYEutkc0ZxSfDRpHraYEZWu5yqlMHxVY/OyXg/xRHr+JRz4NdugmJp1yFDxHUVbttOQI3WDCs9N
B4xy5RCEev9un8+RNVezjuhlvH6J2DIuz/ZpuFSqtjU/sokZ+lSg4RwX44kNCyNHrC6/2BV/UjM3
dHd/2+fKn8nKMUOQY4nwfOMTZeAuLEavmhyOQY5gXFeQKbdJ2r0FjmXQA2SVYF+jKbeyLaK4RBo2
MpIdjxp18ru2U9NsHe/JjUEVAZP4S0kZ6EKIEDO3AbdU8eT3AYsi/cz/LnWxBalzSJmNC4hNBRyc
HRhzGiIVx3RHn4v8a1id4aihawMg67Wiw+d6Ex+pR8Hr2Jv7IprXGsLMLwfKVBG3B99Kj583L6+3
0NJPAOAUZxpH4vIfC0YOhiUj0JfxieGJcgoOQdsG6Tj8mnexCcuO5Nd0AkorpqPFySAMDybHe7Cg
1BW5ScjxX1pBwuMplzlNm7RS8THUKbwvn928xtWqvdOZkzD5SNrajzmQLESx0apAEpOw1/zqTQvG
lob2rbq7osuxdy/sZuJE3P8Pmdpaw7PzPt6PgNVBoYgNwoGDgaSRIo7gZEB1tAHwRmTsHYWFsneU
LHIsp5d/nfJSsw9TaP8Mj1jsXr3yrWLSA83ooV64nxpiYJdeAWWOhi2Qf/6pLpa/Geo+SMe/Am8D
iOCg7g838a8FwM2hQPo0UhTA3EvyO3i8L0y1RaKkUPkolLCpj21y3yh42h3lsf5119IEKtughEY5
U9JXbCQPlmiMN+v6FrH4WukYD6awQ/sXxCsMetxWooKfM8TsXtFHZ1ReOxvFqerBdN/zStKjCi8z
oFkoNInri0M5O12izUR1ho7RibXnWr314o13symkJ1hzJlE1phhDhXa0Wrwsc3sfiQo5LfihTj/2
NRHeWycC7eCNTL7mlfGHTxFyKGy2mbndidkXTNWxuY53yLvC2yqCBTZqLFHUD3ecvB2SqUYTxk+T
3y8UdJs1eSCXLs2uxOsULwDtei6yDEoKuB7NvXnKpczCh712S3FnuVUVDLgPuQsrVvX+A8nePuLz
1JrWIwDyJ1tqX1iKo6NKYvc/uuyU72sWMQUg8bdo4oj/BDVrdATzOdiCpOwAFjXlBZ+f6KBgiDgA
/0WjVBlFtjUaq5ebg7t7sU8kgNHhj+wnty6qLCknF9aafFEwOkZPqICQMEZKchIFTrWqBB+Mjfwn
LWQOoj9juRhSIWf/tqADr1JLRLYQvyBESzeTiusVePn5FTpJ32Sda3P0zUmKNEdmEHMxTniRRU3w
k8JAWnhlvZEzfQTF6wqF7ytnVSTKl4VGwKwdB4FZtBmwGd0Yu3jry7NnDk7Ok3b6BZsNalooXp5f
W4cGB09Iclt8I0pIVxEaAvPHjmax/fuw/+kAwiSRgc97BLOC9euY8zU4IJAbUEnr0vD4Oe8hxoEZ
6OlHeGbPuun0mrGcb0yzlDglwGsu7f6Zq3LO2KBBmJqFUSXjPdhOnfPLiq/TwyMq77JUGPRJQljF
FMnNzlRNVRNMvDuxrt7AYdw70qzJiBVXbAQzNwgOUEzi8pIOQwK4yHPT71+p+ENe8KyBnLNVBlIF
LqF0q5W0WwaKc65NWgidenF+CZvwwfQYZqj8Y16EvhWtpz8pVzl57KcQNafk9jzqLDcNHPIr6fk1
YcA43a4xRE0g0BLSMCfE7Jnt+sWxlUcjhQvdSeuCMv11Y11djD8Vn6VTp5btf6lv/AEyzjXg0Mxj
XADPs6Ptw43D96VYdVpF02DjkwBO2OJk5aSUbEcNWttvtQp9EJ/9xXqPPy01nDM0i/hFp7Z19ZIe
FQPOUjGLdJG5yX4vkUWRXdFWkjuli8rvdRLCDez5CdsZQG4vYV+ZO8sZzVlSKoJ+vlCIhynUXjRT
KxNMs05cEDoof5jDpYlyzCZr1ZxSoiGPQx6HAm73ZbqO/vGHX9aikb9SuOMATlCTMLYQG4z5aVAL
/ntNl5tPCLjcJu8Vy0KoQOnZ6Jp3fpv7kl2FfYZkg/VMHl7DEGJs//pUAYiUOJZTGuE6BfQ47yuc
7TJ0llcKNICGxsWNObR2yhD7i0X3vBnJknoaN4dV5x9rKVaT00LL3s4erIqQdg9sSv1hF0Z6u5zE
jqaS5WLhrZs+EWhMVLmj3l3cqAWOWexWBfRJCGU3ColSSP3VcoHF6IVi4NCLcvBZ3RHfSzVDtRGR
yxiHPbzNoGKxmbCpCnbXpURbV4xAJi5lP58U/ojlwGlCK5HKwj5V9f2cPd0/xOeMInhyDwW7Qhj+
rrUmYgo0Ovz5uB7BTWFjrT9kuQBJPvt8D61KBFIuNVM9+InUEbfCtgvgX5fX2RN5bElJagkPuMtW
afI/cE1f3PyiZE4e+W8oYi043Hx/Mj93xM74tKHS55CgDPCEPoKons2J70TSo4dL+94rmL5ZzJ7x
QvsFJt9CKxLA9WrDQZJaFN5p/CHxC7NeMvfLzhSjfziV6sgfaBgOhWRlDObEk8eASVvV8BW3pAWT
QVeoALwlJ6Lj1XszF4fbF+QQpi+N97xzCSgdIIRL9QPk/bSvTvQwdjMTkmKEQhZAb/Ewj/eXIQau
vzZ/Mowdd2ZezX2vtIE897w58/mupBp7de9sl+zZ3BmzP/tj2IW62ouEM7Tyzg/Kc7ghNSy9t9BM
VALt0L3j4YoIpZLlKDMu2i+sAx6ORW1PLQVW5bTr/81gSCo9Lmho2MOIgmgK5hFvCbt380LNQ3oc
JHXIGdhzjkXWdiws1DkG70tluixO+DCjbbB4EQ3/Gpr9Lc7d/nmuFRFYlnLaCcfY2h4GL3lUxFEt
KwWRoTnAi0MivG0+39+X6zdEOkmQFZ+Ii+WdldKNlS80rMMgOSq58eaahqoc+wdt00EIvQomgGGn
p2qIl8HjdnwYueAqmoIm61eYrJsUmkX7bPqXy14ewaOgiY8Dv4ePBHP0Pyqqqq/RxUwmBvW73zwm
yfdtQ4Z4VKJYhq2alZry+KnSwdAtaX44oF+86lBuwo9KepA1AmYmRFod0BkPzeaBo9MR129Aj0iX
V7tAGMxbw211kmmkVmmUBX5VTd33e8QYes/ntaIyiJaOWlo/6Ng2T85pehszpc9alVLdNiS6COSo
3a29Ix4mDIa/c6PrpIvoF7055LiWsTAdCzWYoiSimqHR177BrNMZf3lBozYwhqyHgTHOAK8PiGZ8
hh/vY6mVcQlHkfuHbq6oyaLqz2YPIJHftJK9enArEqnRktr+CfvK0Ofjxa+obMcGzJQRlTnpgb/y
+h+rtgLlxn8lYJeXEdoSLSzju77U/sr0YnwvXhUCqok7mQZQXxmK7fQK1/ujXWZhiSGfP9ymqRR7
3m5tzlTxg65l6kAqj9dw5kN7aEXSE3skivf8MsB84G1Qbed5qt+3PtNfkPyuY0NBSiOpe7P/notx
CUVhBE5MnQePeBrU2lk8eSgYf251+FEkHwC6pIPzPZgamR6GIDXXEW53oiwAKWQkC8BtkYa2cmiW
/59uHH21q27RYqKbqizAeYURDBMPCi47kcdYhUjRmcDWS6v9pnYPayiKOaW+nF4ofsmsuEnVwXdm
f/SdERwTWG5HvPU+1ppR+vFLHE3X0uh2OUFK2YTn1/MM+B5FinkGMDx6MH3zy7PVwaHwBghzpaQm
nTiv0D/cgK6ThDuSvbWKkhq76ZM9IdZ4Tjqms5byHxcv3GtE5oSxja74LdTmnIfRLuohO9hcETsV
hgKlUYC4y/2dMibyV9CaV4wFvZrd8V2SBPPzz1/1/+9+up+yeR6zBMq9WHs6P7r/4IqGRSeatvJF
wGPwUlgPOihMm5LS1gQtRMSS3nOnd4g2yJL3/jAsr5fnOEmQAiZZgKrvwnFyOSlTXHx82FE565ZU
eqH+vp+qTqVCMwq5S+CYOnIzObFTjmJ40M/Lz04Y2b0SPSzOeDFy+uaxrnQOOpgOFUuMOwUEoYkW
lmMEMxf/meesm+f6ky9XEFqm151IsoqSXkLXvQRXoCGS8fjrDxhlMcYmas7G7mxpEC5YFmTmBqf9
6Nj0d1+X+sfY8N3KdrJwIdl8aDAHw5qwDRNrJzJnvsfGg4CM5AiGqpzKVjcnN1Bv7m7BPfZPKwfs
ZjhnmuiaCvBxnPrG0+dui1LPQlaz3URnx+9YqQ/AhruPm3+pmyuqGVujPyB49qqWHFlJSIHBDB5n
Xi6RY3NhYax2HE4Spa1LM89kTcpC9iu0wFk/Z6xqQ9GX0FVbgFcV1D19w3sr/i5kWEsEclABMli2
S2p/8qXRTBjKx4FKUZMnxDFM0+Rldl51lScRGWduFS9OT6mGvxtFOluSbR1sIg2iG0XfB54Nvf1E
n1mYNX4fMx+5Dtq1iQwAGkoluhr2/yPLPY7pAqx2JbyxenmVOyb8gJLMrrXgTUyjFtrA/ilq3id0
XEdEVtvkJyI8oeJn+XvqjHFc63MlYx8xM4YyLOIX43hEifGrRxTLu2nKogVmFTPYEQVIBRW273+V
2D95ALcSl8QNaKZcX0i4xnLT8UFt3UOsJ21F9rwL1ZlhZ2gxxUWUzMugidUCCiCDMo11RtCs2e3E
eoTuuyMc16m6IGJSAcVhZ7hYiW9Yw3BwMBM0fkqRDZK6RlV8UM4qG2OwAZAlXSUsxmD/1dGGTVbg
YA6aDVvsx3pRX13+6zPG5lNTIljqvouAHcjx4WnklqtShzx2Na1sxPVHoIjJ7rJQ74MqWVfP0Ls/
J9dihQlcnetqkdViLS7mPyMOngbeDhPxEnGg6/uUejauGbn4U/gQfdxgTjoysIK67ORrbbA3QLHo
wMrUwBqIINbiwagT4wW3Wy8iZdiHKdNm8G2mJk4KAbdQoeoxjnHDmZuzdEN7WSstJMOihTWLvnA2
tsyO3srHVJtveJDne0VFH8ck70uYusPsZR3NJ2Ee3tx3tCSn57B5u9kp9f1sllqNlj2EiEBX23Op
CTAvy0/u6A4f391/2JL9xWt4jwRCCPgPF3AyX7HHEAEdq7Zs/7tubvF/zmbCmZUlstK2lGXbOESO
6RxmJSyWhZuxeL4mj9GIY2l+BHkdp2wLQhQ5FNPFsWCyw0jScpdVjfD3vRkuyUy5qBEPlQo6DKIf
Fw8fiEt/SVuA/24t2NehoCNko98Q4PUGoeWGJTVY4qRp1nlMGu7vJV0YUkUiieDE60HLEdm9USO7
WsXPIM6q1s7b1ipWPilB5HpXyOvShu7FS2sQYUOpq+1W2IbaURhxIIl/797T/lLivjRBqOoFJbz7
iLlVDoPikHVlFvHKXnp+mmplbBof7I7m8D3crGQm2Wzp0SsMCvnJda7bJYifHiKcaO0dbUROBi4Y
rWxSHHA0ymcFkx3cqF6NBPnvQUsXULYmgzWex8n5vmNt3xFSWZ2mYhAn0ZDWS15gvgs6Brje6iiH
ll90PEMyJMxkEy1HFs1nCFBWgFOoKwFwK1Y0ZshA8AlMtPnEPTGxpOahjUaiZCbasLl1Z4jWfbDY
tS7jZe/tlh1VYR2jPcbfMemwTuYYX0P9104Zv+O82BH7jn2H97/9iGgO0WAGnJ119761a/yv1k62
kHdD2ZSzc8W8B8B9VKGNCN78K7u+zu+p35oMxIRQMq5RqxKwFHcrauXuZJgwyQs679auCByphpWl
Tvbt0trKb7C3SSXZd4r6Cp+7GZyALYNfT1crhHXs4P5qW66Pj18b5UV66ckcnjNB7noeEfqWO5J3
NjE1hLL/IYNQJZxRoVpx+NPl/rd2faExhaPKtiHF/l3sx39zJDt+VG5dG4Ni/U18dBxPXAhQgLDP
GP3bFjnly2sv/BrNbfziQ2lam2Q17QrevBoUQPUsN9TymAxkGO1MuFH5yp/fFhYgvjec63NSNpX8
nlde/P0tI6FGBWaB5mvMUKMYH8bs7IvUtYzB5NJvMZCmHau15eRgjlpP/rGzAgWKWPBHAGl8wt1S
kzjYazReGwcWb4iTKwPTT3xOS6mjp9j9IyVKfK/mfm3Hso9H4AMnZ7CznS0uFJfCIMFGIEhIw2AN
J4p6Iq2WdKCA07AfhfBQuTXmlQpxUR3QQLWf/mIRAwZtHrDYFEIy/hjTdFtIHK2IUJfSMV2hjb3q
W9IrBbmdAp9N5RWY7NfIGnOv3UkFooUaz4a7iR9JfNTBmqsePcucpyj43KKFjRoTOk1KD4OOmPqs
QYfMMElo6ywgVS9hqETNl0aSzn6Z50sKP32TOBvL9Eqk1xVXuIKRFe6exPTI8Jbosk+1/xrs+yC0
Aue3mmvqicY15ZXlNVB0biW0qgI5zGMbvgD0SEhhmf3fRSn1oyDHFNXdrJcK4Vp9idVOnBpXHiuA
/3KFJfuKI97HuSRdPnizn3fwDrXgiRVFzXG5RiZZNkyC1FiVDiLHrNugtagzn+X918vPIPaIF72L
BHWGLN68n1TXeHoM8IG7x5zoPEVPbMAlEKJYj+gOEfRuRG8T7b0maxBPuRAvu6EcdGmLGDv8GA7o
j/6QVW2B5z9abLxWsVhS9VbB5PmvyCs6dInNOvyrjpbZDnO9NKn34W7P/AFqS1ZXG9pfgfIDcICt
2qm0EG0QnWq8+6IRylU96uw2So1z6PGCxnHDwowyotw3Dj71SGU4Sy7QgfLEKlmRASAUzObgzPMI
XUM7wx4ZUu6cuI9oFaGYFjokbNH4bOywzm0IiqdEFZQdRCU+tJvafEvyUFMA5VI16YFTa87qUiGb
//z+ANOA4TQ+Ude0DL1Z4tVPHO0QdJ2mlb8TfZueukQyQfHdok+0vMxF4M0H1zYTlXYoMRH9kJxq
S5Os9Eb0xR4L7BDIX1ehiRevkxHLayxaxhLOHnw8ea/AYJ2UvA8RrMcsPvZRfMrOMynVic+R/jXe
ySRZ4NDL8fHHLlhn87kzpfEtwC/2IiDvnw0rOQbsvcpIfOVV6Mrpsk1yMDCuEa6g3aZW51yJUl0z
aqJdIDGfQZCnGGNrGKAtEE+QecqiMa+NTUfkYeIBZQXZpahDDv+VZWAnJWCyeIhC5DRfm1UMtgu7
l+y8BgqsZ467HChDEstWZIdBTCKhz0RT3T9e4j1rR90skpiXcY2R0f6ANCdlTiBSKNNWXeJj2Qlj
ECYBLoLKVzkmsp1ES3FtQ9t4PCtiz9bw0ncPDkD6WjkgYj0lHVIOwaIVka7ekp494CheQWEhbUgh
cn4pnLtkaa+9LhQiE6UG7cpKyUrEgzXXJlax9G34vqLcCOKWVaMSFSLphwIqT1hvjjZ1rPZD/A9o
oqXYO0sokYmekZSc4a4TYW7W2BsDVmkzdc9YlWG2BSKgxZtxoAdGkDNiqKlpjYCtOXL7Y371IUcL
/Ss0piXKmzLZFs6Tj5GXez8m+3Ytil7r8Ic5mBB7iPd5m7cY90G82/EGUKa+gZnEOqeC8b7r1Cjl
kWQID6D07dpgVeuznOZ8E1WPUh79m9pihi6ceKhSqiLgE2AK/w+/hjdAzUDKAQRjJQLToR1GX9sC
tgOBT4lFLOGOOBYSlV336iqqLQmtm4xst9GN7U0TPUyC+/jOH/R7J6+kkY1vbjlKxbNrKMFNByRn
/wanZMf5lfhnsPQIoQ8gwXysbs9s/kwgl8Wm+Llg8Tjm6i+l4PaUUNG3FWe9dewZ+E2z+AaUFsMk
xZo0tG5qOt+MtBQC/EQkQ+GeE+bLBfzxN8dqQhBebhICw7U+Bviw5uNaxvB5RkSQYNAI6stByVI7
Bj0Ok5xRMq1veCvAYB+RVZBbCpeSu/aOrRf6Zy+miT1Mq9jBZVib2zyYUezbppqu1oxMrpafC5iX
z32jpMOEf4rNMAaMZmFwFtr0zu5GWjgJHciSpdqtm9Lx2E86V2TLBWd87jz2GFCV0zJaML4yj21a
eQvwGLPboTen5lqnpHbV3GdaGLIJaGlftzPC9PLDlSlnrE6djlYQ2/0Nzs3MNIFXnfFlcL5AXBVK
jb+EpKzaT4P81ZehZzDGLeYul9NwqBNwOzxdcUOQytbicx5gxdfcAObSFVqNoDSIJM9tq3W9XCiI
x60NRZ8k31rjUV5kNJ0WIzgxL7hJbyMxuaeoqM1iZ/iV5AaZrFJ6VurKzfIYEOMGL+iQZdOVYVCA
fGa8IDQJC3J9RhRCtwS+E2lhXUSXOvfpzbVno2BQF6B83/K1TtmJ9XpH6uBN2To4V37ZnSKl6eLr
dXyPbJeX+aciU/j/6NiGWCC63uRUg4ol8zzJeuNJnFOkqO3PKntIAvzq16x0aC00int8HSYNConf
a4OEroJMKk0gw86sCxNfRnklFICXPlQ/gaHzfdT5085JW9/O5x+gshWC/x5JKmvb0Yw5pwBpyq0c
2HpsLA5XhJhGkWM0PVkI4u+y7aAlEirO0je6B4R8rKofY8xkCdHZxhgc6Q/squLaLfhWLNjT2WbC
KAsoBk1Mub3H4CCf3t0kiXaOMY9gpTQK/hn8hLab7pJzcJplGM0rlQry3pxISnDis5ylB1PBcQaF
A1P+/1H2brwBtfcCwsd9j0+44QfvCzQwGnmJh+m885PaWUjxadev20Xqr1usUztHc1Z6tLvwCAfe
lJs611x5vPLMpih0WQ38NktuvoOT5vVsJFFjqe4UlNNzS0kCdY/K+/CoVGlaxMwAegvYo/oleZVo
7jxfu2Vw2Wi3Zyb7ZJWwFz7TTyswZJguE4rPAQbgj/OmB1kQhcj8AdeAeiuAGvliKOiERugzxIJ6
amC9v1cveLB+BCeoFNNZSLnmZuNmMcAAYsZ8sgBwbNX4RHvo5WfDpARDRLqZMdLDxqOt9U9dMjel
JTikrRuSBB4SyzY9vhHaR35oBPSor4rNV/zd0AHEH5w2ODJrft7RQ40uqlKbnkQ0uQ7F6wjtHd4m
F1rXIT5QVxBlTH71N3+kv0JxGPdYHj6cRek99aDG7KWl1zLW8NrR8CJhds2aV44FC/tNsdHVA1Z1
ORO3/+v2b4DjMTrrOJj2915sInnjbEdNkTB6KZygH2A7QDpMDRSwRHxrNemdraml1zOG0g2oNR7S
EwXcUj0fsvsUxFYLsArxE1uaYruphbvfRJXwRTXQpKz+GcxD2VsGY3xOk/z04fZcA9/VDmyBIEbl
SIwY7hesPrujHm4M0K/R/xZ4XIrC0/8cpPzI0bZvfms7HjxdTDujocnZ2hNKZO4jbo0FbX5kSyZ8
Lg5pdBH4LqgiXA16SuvgGy8Dnd+aY34x1tiViR7BUCj6aQ7v7ExzGyJgS56YyBhrhiFvo3ZH0ZDj
gYHwsALtrrz7T6NB5MingdjVmHCFySv6FgawV99yqdz5WQu4qudXC465s8mV0kFylqLbn08rWj8F
B4g2fjNr3nx6ysdQrN/1i6EARccsXV1okZmpE6SQeheO387QJCVwoXqk9n+7tDzcKL+SJQ2xt7zn
0/sAxHHDhiXGEykUpMvhoLL0QdWrqkxfUcu7M1PU0OrVr0oBrENu4g5Kc2SBiNHFgug74v8l2Jtq
DS3VeEw256ro8VZ/2vdI14A9twYZZP9saGunaFtVhW3Hqr18ekK+xZzPHHaWSuZCxhswA8cMhkeZ
pPshFYXWyN6+HKU3kOwBM7ogqcVD+ZyPflaLOqxka2ZKMbQPdZakHMb8fKQkdvdkKFLsc+S5Jtxk
eaqZOefBR3vNAkWwPRFuaMGiM2AT9/+xBbGIdrp6H2dJxPdGCG9umcgUD/Z7HwJ8t6qckUi59Wx8
BQAFeFmhhr2gbDJOkhHaEtGdF04QJgsNSTJBxA3dLAM0sehTzUys3xJ8OzJIfzAdvbbvIGg22Uej
SM2S0qnaoXu9pDp/+u2L+fbFyDTeBtC2AhkB1bSXJW2nh7DSESXvyyJIcczzx9PCoNRD/aWlPBRd
c3Tt1IsCwKykOsATBLj8SvL4fM737WhpwbDLl1dfXbgYuXPnO7yCG/6Vy4yjJUEgw2deJ2FpTQBZ
XTmj8bJ5ify5LNGyY6aDUBFrcz+1Tfno0rrWFoA66JJ2ohrmNeKhwta+VSf6XkKS/F+o5wFprcZz
G4yhGrErxIIt/PR2+cukUjQSRzxxRSs2VwvfeXP0QjYW4Te8dyuzZM0b99rBYXqq2ck5orRH9321
k4auMgBb/b9MgRj5ZJGxmexy//zy/Rsvom18SGUbu47S6ex9HjHXyPfCBuak6YY1VUo+tFv0RNgc
wTBrF+GZClwRFxtd6v8Jqr9JFDgE/8VsIskn9NlkAl1xfB8ruGX98fKk4A9rzgFqjQirbagILZ/T
QHmzUHQXY6UJ0tDrM5HenoAe+D9bHdJXghZ0e5EcRzxNkgk6EYqNmu4sb8RuO6CXF/BSVgRnE5SH
XFF9X4ilypzqRTVz7nGWbbs/nGGjvfotylJDqC0NZvW94ky0HCyxxYACcT4M3TzTAYVwxUp4aVmm
0vEd7HH3dCK+Xu62nuChGCC1oWg+DJ2t6eZgvv5hQEb9oikSpjQxIYkNv6PwejhKiR8CGJlsDKU1
16X3HQyNGjCJ2fwrFT2t26TCAr7EsBPV1gM5q0Dy8yOJ/fw576yRPRF6+3w2pMK3Ha/lOJ1x5rCh
3T/Ak9voBnl0qgyTz76S+CfhY/3BiiMdUa6RW4AJaCznZjnvbT7vOrndoi1XKGN40NI6eD+id6iT
9DKMZ5LIru9OR4yVkstTMD22AXZDhVXPGiTInf1pwVrUiKsf1fRm03IW91DBUZYqsmJLeaP3GFHc
ro57LdySgHY8jdgkMtqVo15pYgiLxiHbwOXWfgnkswQiHYpGzMxzd8NtHutEZvSYZI1EI3puM4xf
dPe+m5eWjD0/g87fhfzajzyzh5VzCK/kcsswyzpzuoyHt5I0EQieVl8GQGsnRyRqGlwnPAl9R2vt
WHR0moifFdXXeGPRLq1hxCzbpwZQkffaY50Clb0rhvefgZgNDC7yj3LyYqyi1ZCzsFy057UJhN1a
EL+hafgKj4uelOQGMk4LmAFT4MDSZ4e7IqYnptEzxE7gYOIh/5ZhZsCHI+uQv78+yE1NAsqgKi+Q
cuN4OB+w5z8C1WgZBgkO+H0juPn8llhM9SoZ3OwwPfH0jSfTk35uE8pHc/JYaz+b/qoGZjHXEdgT
dieg9qe1hpkAE1AfXwNtUcgFiHD0fXvcoxfJ0AxYUZbmFM9xwRjVJJlsv2ijhJ3eG2NP6uZAxRFN
+FbFQFM47naJLC60CDS3w5X5+6AcHVVWZ8ZmEBn0rfYf/DwPkr4QXzgvq9kwY39u0vqaVPlwGH3Z
NwQ4raRuaPk8prsfqyo9/ntaTsrJBaMsYXwVzNKrKiWMQB+9uh8I3PcVP7lPpAFAHoHh7IPmwtOZ
WWrRCZVZ2dkZ8QKey5OMmBfKst46YIMmAdaAjxStn21lUwYnaZDgI4AduY+MrIdKZ9+P0MYpkpLC
HlRqwKmG+8uRJ4bwlxNVFLh9OWKH18jqfI6JpwWZPTQBKNDOrV5R1rJQKiihQCjN24U2D78hh+zp
yOMWaPRYfNg8+kyjJbhme1asoSDjzdg2iSRSieaSjYdFcEQA2klq++u/BgcmtXH6JLzpg17WV4Sg
Bz6JkNaiC/Rr7R5+D+2HwwUjwl4XFmRFnyxkBD7Mud5xGRaTykyWVs035dJ0KYBtmgMQet//e5XF
U5geG8JdoZqCsOLtdHr+ZkbJOWP3Cl6EvkjdQrELe1n6rSProX8Rd28eIsV+leDj3tI7WJyII+54
cBlgeLzTlLSYtLz47/LDiUm16ActMrnYQaNMgcdkGEOyG2Kf6C3t3feO/aVLCl9ghVB+AfmbmCnD
LVMIZjjEWePcTBdrU/lpst9FGz7C6J/whaeGtP/EHLg6XzoEQcFF/9UBSp44K/vsCHFAl8HpV+td
BWrTwbaTuL0p44XMu7aRNTCwsoZL6ly96xtB11eywEz0jCMOjPQdLmvO4/aWOxVR7TW96BG8zwQR
sVON7q1LhyMRJSxn1Vat/vn0jPBPXSjQ4B2dr6mqPVvPMUxl3OiXh75f/JhN6AMiRBA1tCIhqvN+
v0ZYR0FATjV1Rt48Rt7PkPA2fDq+RTdPnN0wj9FnfnRcK+WATXHsnVBPqSD1hGnlGOOILtmRHVFe
K/FohwphhwIHz0uXxk9dScUQNQYJ+D6c+/Do6JvpjWivD+zM/61fL1sj+19+bmAGNY7NbULiQZQT
BYbP1hORbkj0JuRI04f7mAEnM8G5qgt0ET6ItKFYpQdTdKrbTg0mOp58hBGeEzU+Oa+jioIil8C0
TJafDaW+nhsPvUN4FscAGYoxQfLZmVTKA7T9cMQLeM+Nwsg/KqV7VpvIDbuqR83EF+MePmnwe4Uw
H39UDoUSiiNzFNhyzZWDWOC7EptNif3hnF+9bXJHCZH5AwFg0k/mq3KpvngGhIBg53+8RU57D8S5
J5QB1YVZlLkacFrm7IjlWYJ7ZXfTXGzZ2TzN87Ql+OcxLCBbeu2vYPE0U03VoFEzVRf/YVfRsc/M
+mNBztWpHanHPAPPeK5ll2QerHA3O4MfvSt3/hqCJE0lYwMjqtqqRvyJPdVdxwMNwH9ZSLkMydGN
aCMQJ+BRvZCCZ0vRIQENfYn0D0lMwlUon7wxIe/i8qRywKk771n7BKVp+5cftANtMQPBWDvQ4ant
7TZS0WwIHWZ8u1XBAAxl/xkaTXzezSL7q5p3NroI91IxD4tVRuwp5RPBiblo0N8S5wHPOWdFloVJ
V5qxu87B+JGGPcno/dcJbcBqX0Sk1IO97oiwIp9sfgAGah4cbUuczsSQnVkhIDa1x5T79F5bEg+1
XhvPJUABUhWN62fQBjKdhzowzUV0hPE7ymuu9o0/ifRoGKt/+3wqGtnsl42kYUAH35Njjcex7qXx
dxf3BNiwnJhLnHqAV/t8welDAABfTsDRTq+bL/TGgaoQCAjJMBpFA0z4Sd0Qd0RY9/fXDZ8qMvoq
2bfH7EA1o3f1lqvcbdss5gyCrubX6L/hLI14H18FtC7Zx85Vxl/wLg6aQbRADTnEooxfEDMEWz6D
TqTWzCFNuPliZT40Djo4184BVS69jjquRJNqzKSQxECI5hAgaIe95GSYXxIQoR8cmOfTILj2NwFR
6D9UxqSxtJazGXxkZGO7QBLXhnyfPEXf1eFdLOr7nt519eFIclChe7ZNVi8553fOVIn5KPgloH5l
/ioR6+L7QXHJuYY8395WmagnapQobr3Lvp8Fg+m7rphIh3k/ikjUo/tYo8Z6jI0Dl3Lhr9WoJJjT
Iz4XLPQRBXc8QQU4Qe5tqz8qwj6o5dhWzp/XiO6VSV+gKIjVc8bnLZQrmiIP0lCzgXo7Z9w4sG85
9auLekEaCsQ6CPnXMYr6iQEzhdbZfrDe4LQecawjBWo5fwbZkKxekday3Y3qSJcVt8vJOG+qVi9I
eKDxwZO/nmp6VWCAxKPd2+2KffP9SbBk+tgtFbgWfc6jLQMdPFlp+W0o/yg/YeyOX5hLxGWh/Bah
4yW31x1rgbBZcgV+fPdKHpJ0QSx0Hm3K9tdlRy37FBDLjPxIWhapvbFc7XqXgDF00TvkHfAUpDk0
SmfOZpMcsxrW2rnNURRSXjqWU814BdyCiVTpxKMkm8j6PYVAc4AKJqSvhgqvl7EX16Cd8plsB50o
0zea1ryfaca6VXWOZMC4yREE57q7RuYVlJYfOZyk1J6uA61Vm7szOmvlEfVGqtYz9wpkoQ+IlEXm
A/BlLBZA0OYh0K1RejpFj+L2xTHjOAIqNM91VVPXoBwwxR4poAGQRe/DEcnI6vayA/gQ7vZ2Vd+b
AZXNNSWJjCDD4gSf70ibj+OFCHsWTmWi1qSjFYfIaEX2GLfrBQCrUVW3XvapKSZk+uDLBpnRdG36
Ruasm5T5tNd/3KKqqt4HoR5O4FBnUF7NOqVIHwO2htwe5eEWmSBdB4A5zO69husbQs6Aa00FOroK
vers6gZKMWd5ErB7MH2qj9j9uXpa+57XFmiFV/Shs4SID7cvxNzLzID1XqdVJ7t3coiGbS7mNiuc
jfYB+7PHgRZnhsUyPbRZb/yI2065RoNpDcWwmHIFaMpsVuxHxxXeeKH0ohBI33MYlPPhrUIo/vJA
6s0htNe0eHmz4zF76MxA3UCAOBiUGw+WW8ccFvzF/wGWgNxUGaM3dIss2FeNlBGqIcr6hPEpfxEy
LrfZGPBKheJL74TLZVyWegXOnNEZI3ExZJkpWTn63b0Kspymoq/mJcCrVVrT68M7+TcF5VibpFdC
vmRc3c9fS0kkztxkXCkE3xaImpBpww5SjELYaJDwX7mkp06+B1o+CT2XLFeskdBNlnmXlLEvv8Yy
XaT5Ktk74WT0wz5Ko1FXRivXsgztRH4rOqZwMQmLn3GwWfjG3K9Ih0kB82kC1alUX6QLg/aOxIAL
OwC9Pl4wCN7Sc8+ekcA+S4hRe/s5xOitTyZ1onnf6XMEtYWj2Vol2W7gk3qC4dGEFRFG4NggDfmU
x37JcAmsPV/ZZHhlTxoJfAw63pUG6RYYRXpBuPHQEDYURvPgH0u2wzK/BPFTz9rdsp0hfV45g34k
x3KngfeErE3qhFIUvOyIWWpazlmnUTP2t1Smyfr/bynNPM9v8AjBVu2hXgmk8le6+Q9vFDQ8E8mf
E7d5nnMWfrGGer+TD6TH1+Lb6j/X7HSRwxwt7rU61tszbVc/pc0P6PwhvPpqUnnJLEZ2gBN8PqBH
lEhHpQ48LLVcOFd0epttYw/LmDcFgKpB2AfsICednhOClowSHjiYpumlKzQxYQ4kQEsMhCxz4Aow
57XfdTHfOXes2owZ37Lqgj5F5oP1Uld5Cus5HeHIqYRMd5178ipdpt9jv8CFCyXxXNxA+pcC3YKA
ycCAyHAB/bAUmbyQHAnSHhxzljkuMugWsN8OUIso9/Vlb6rfIyJpcLt34FNVI98xU2c9fQNaRfJk
2/eOksY+veWC8XxNiV9rACP5XNOMjfzSh9IL5ztza5EJ4C47CcT+oOCO47u99S8pCY+VNqOStg7m
Tr3Wpnmqe3PbOtq+km80gQ6xDBjL3a0pSlh5AfZsBD8VWV+tEzUsnkXR3rF4JS4yXh1e90RrBzM4
5tRdvJpHRfuX3+bu9T7Ij9+RMegtusdk63CsJbJBUssR0qfS71V+7Mca+LciaWFMB3Kjh8lIbNs4
pemTznuxf036/RSbMweYW94gTwisRnGcer76ewimmvVv1fmzmeshsQfgk3ytsandDXcYwJ0PicH9
I50TMHnZ/qLrVGrM6JLyK3F1IUCvpF0KxEPGmtbUCYQdrqKwfbmjTbmwLXliiaWKoXg6yjph8Et/
3ztOq6wPhbsoh7OqiEcVQJDbZ07IOqv4eyhkOdy4tAeAG5oMp9Na1O4x2kZd9u8aoVg4Z9fuj79B
Nnq9esYb47hdlRLz02pEVw0TiK6QFl+uTucnKg9PC/vExHLYePGw4Q67JPn351bxcMBOKvYN3bMF
EKuR5o/Q+dlSy32IyzpvKRX/DiMkKVD1pVzTRQy1OO195HDbHrVkRSTlHdoW2xfCi0a2w/cm7vid
9TzSvHhxXfgDSiBZgreLdGNmIYbBNsgdYNeJyrku0h3excgRlqcStZ5mNBaS7o3oe/0xkv6gsWlm
Xfwbavms4k1msUD15eTsCgBh694+fyAKSva5sCpG7JfhVwOkmk1Q5xH293AHwMENK7r5zGp1rqJy
X5fm3Ew1cLTFdVJqJGMKNXEZrX7h8eGnnqZQxnaRu+7akUuYWiaywoIIitafGpUQwOIdjvwxmk7c
wTZliHPI5Ybh1hBL63zsBPuGi6F87d3pFstYy5FyrhzdVBCxl0EcQMAr46HqzcnxqrWb/3fM1lxT
hvNaOJ07mjd8FzlE+zFy//TV5GSPIdI5RfhkO4uncTLg7IYfLYLja0w5/k3V9tcrHXjANB6mMkFJ
MBEC8tBMf9wecUotTJzSHN/kfzzQ/THHsTsbutd6LjEO8DQIG1dOFlViHRqwVdsY7JzPadGWeBDb
irl+8V4onxIcYt6Sbdqrjb3L8bHl4E0b/3MReDwd/co9P2ruyg1pj7hoCbTOeJThrfxvr5sOVFEO
Ysvy7/UZEHFBnLavnI5326r+jRTJ3rUb6YV3/lZt018UVZ4yCt1D9K+L4JqwX0K9L+nRszYjbNel
31YgkQJrlccVtq+0p3gByB2OyQ5cT1gIHRL/3f0evvYblBWNYfis3DUTnd+N4NoyIZDRRMK22kzT
6TMxYdBFJCtdeRxAoLLLyWMNX/kchBrRFDmvdDUQSMIZ7OXW9toA83OQSr3N6OiQyRZk555b81iM
VGvRMDIejcU+4ICD3OT8D+ynMRPvXqZI7Lirg51ci9QnTaRjIIo0EaJrx8oYh8K2m2i4GuxZM2nP
15CrQGUq6Izjx8S43XkFO4PUCW3nIa60WS8EKSwIcY84uP5lzNJBG8vK+yto6LY33oIuKiOMk83s
RdUa5BQ9gtcJ9vKF0KV018g5KTqY8pQvacd7yimv8ZdlezYKCAZPD9uyrp2uQ5HHldjrfXhn10lV
R0CTkZAqKSKzylHDrhtv5x7RHTV4BzI5MurdpE/aL52dt3Hzovb1ElvHlpUrA2Uc/LcvpVeXL8Pj
TJGBQXcS4aYKdOrI+HZbQ4ig8a2g29L5SQKFGrFjDzVhJuqI/a1xVekPc520RTzmNPRKWOjTx1r1
BOqhCMR6ta8aStiC1fNuK+m55Nd/Px/IYHo9DWfkT1hHWLZMbaVZ+RarvwMzoQqk9hQ36ACSkvJg
eM4kiRD+2xTLqhjaD8ADCl2hzV5zhY3f44HpjjRBN5kMkbPxD1Zr7T/dnuwg6Qtt3WydZs+2ccsF
TjUTWDbxy+YfO/mkM79RUuRv7tTGfMN5WTeOjxLRyxOHRmYpE5Z7HYkTcsOtsU7NOp7HngtMIZk8
fRV0DfLfHSWpKTa8cSoNCbXGBPgBgZ+ODiYJGBZ4UnPT/CjhscW4I/NEljwvqgKuS06nIkIi9D4J
lmlsJ0Bb5+lQdrECMnYZzYxEpt3oArcdc2pEOK3J2Zqs3bfo7liSoOt+jCnnUKKxzUdoE/+1G0a5
QYzUigVkMrgW64aoS9wBuq0YYimEKXYWCwYOPU89XQXViNkwyxR7jwm1WkaONas2xINreeVnz3qU
zfnoaXfDt7PvzPQ2+IfVX01OenaeZZotCqRQxqH0NHnrZa+6lYJGOSPKIOrV7lKYjgbrQ8BbcpDx
6wVIyMFIAKgnfZNjEH8PQhMKLX5DlFBcO2q5NxofQOb2ocBgq0I2kMoogX2VVgYvWUdXuS3oPP82
LjeT6uuhBiZvZUgSgiYkfeGIOs0H8ZNfYIQPQG6teo8edRZmlN8rJ+gVztXjbrPW8+V93Qp8S5MI
a/MR6R4Dy8p7RC7+ffEyDx/8c387yzDjAfpEAZNDKnsI1covRYZGEXdSG6iVewF1717V0Tgf+9RI
x0ZoI1l4hB9I9X7u/RRSjpGE8/Nnlqkl3zq8x7fYuoOknGwF2qH0HMOAMMi3l2j2q055ti5goZrG
NKmV1n4zQZLK+vQ4VJuNxKS18ZERD90y+pd3VPyR29VV2bYS0I+nGixS/30Upudrql8Bh5AIoecw
r1DZKBnPbVsEUlJKRnfcCJ8wWoC7D1LEzHHDIdQncSrM8cnhdIVMXIjLsO3teeWue8VNeC+3GFky
CPpxYsj5VAbXgy11f4ssgnslzwSDU8NPyH6DMm96lVAjL7UzQ/dqE3Rmcf48Mow3KT28SscFH2ns
RRXE0h9pR3ElEt+BDHo7P43vaswgnXyLY8hnmfjDgGjNs3dwYB5EzroYJHQz4L1g2DC00yZasWUQ
7PyM4I5SyvyB6AvfN5ggPcE0cTMK1cXZua9SJLdsuKoXTAUYN+L54P1iKLxzDuCdWX/QLIi8RE5D
F8VgKTvUeAiAOT4lp6E/Lajc21bpwJsUbfX4LV6fETTgf9JnEtaTEWWKEQak5ctF96Gm10GAnriU
8lleykkqVmBpXFqC5QMZ9ptyhIC4f4JDkpPA1CldgSEAoDqDado0AW8Ckcj7RWB4mQdsbiODK8UJ
qR9PveD/XQ0RRdV8x4xaC0F4g1XJt399zmO2Hg3R7YamoA/l4l98zfWPs3wFj95icnJVUCGqH5J/
Yqo4v7VDzYvPowauFmJLDd881at5nlxE9wCKEQCr9qyoUT132MZ4/Yt5Z6Ys066+3/xMhuHP0+u4
Ltw8ag3KaVWKobRS5TBuE4F18F3qoY0IWBIuWr3/zh/5C19LWoBgCO4Jx2ExGANhqOyHZZWifBPC
YBtkhI4A8HI/r382od1AO5mDCrWtm2toyLcn2joKLlKfhNEtO1/iA43DcHYLiqHOvKRmtBfrKi6o
nERx8L42t2s/dnOZmt8pGG1qqVVr/USiMMNSxWURvtiHG1ZCnXcyBpFweeF+SgAX2h3pXFT48x4N
Do2CmGTAldVcHO4Hg6wwiuYh5u24+qfejvkrxROkykFnMj5ZhSkzzNXhrFPHbteXDOTqjTDlQvjy
+kC1A/zfnxLddaBYuJ7TMhRf+zRaMB4AG5XxGV1WV7gEmW4JuLS6/ehIallsqUlBfokVVknV87mq
HFn4Qg7E248XsLGLuBTwkZ2/WrnPavIOgHNaA+5dy8Ak6LKaMvNbyE6rIN4Xzgf3L4J7fVqJwNf4
PxyOitsaGrbi5MSswiNHXpKcC0jMtCvl0MmGLe+Lfm2LD6EkC3jJ7Gz4nBIN2LMuhRae4JyWi2Lm
jfQ27WWj8/NwO12+tEA4xhJp8FL0gEwFZ87qKA+6wCuE6Ze73hCdfaDyXHBiBbYdIoHTmsatKBGl
SO/H3BNELUo4Aq5Q1R2rBnw4ulOlEGo6oWXEo96DQ92ShXP3YIjFr3aU4aJNwhU/xXBNOaSlnOSm
X0kmInhr1tc8m2LwhNaNQqp0imTG1rKqScOGVewSWFy4ouL90SRNSnhFBbpqP5Cv1nK+EDGid3Q/
uvIo3ksecKdh2oByDAuDaH1nzUczmIc0rw8T5nYx8dJsurx8qbD2M6uzUs7F2n28hp4RhCxKdAcU
YguAQDOCAY61eGN+A5e2xtE4G8WBR4VcckZlFVlP0f1LS3X9W+DStlq0e156dF2QGfFHx2aEfKgs
KmmKL4c6ctCot7GAzBSBDlqnFBoYBzuMYH/XYLk60z8b7uX46NBb4Awk7d9zfuMyCZD9Y4ULsach
YzvFQ+Hkumx8izWCi8X1HKrKFYpYfRqG6pVQFD4kU1w+iG0Y8g+DqO1RLpRlHwLjhNv4Wf2+0baF
tSfmTT0oWz7rkXDP+BY5VqNYCfWZBBTM/sHvO4vxBAhdVTkg7sDE3bZD0tRM6NKpv3dvppv0fAPm
dxdy+OuFrpJjGn1zG8FR42EbevR+Cn4DgBSkzuEWMppliossqxwenTOhXpM6OL2ZdVz419BPyHsw
Vnm/ST6oMGzF7Cm8ehL47huV2xyK1FundvmVg4i12CIX/qrxPZXoompHJxhmBEPW1Q0VX03/H0Y3
qE+L33vHD6vbj41IOA/UVyKWG8Uo16K2Se1ZbxnzKZsqgLHiz24FxUO+EEkoz57xvWUonIhhcIlL
3z/D6083rEvo6xD8m+DjBxN40DdLFs8zxi4MdXL9BIg7+qGYSxetGSTlu9O/o1JQ0ZbaFNtQciu1
1zHAEzU9rvAOb94g0jp2r6GCfvFbemrp1EdhalUZ3vfP/Nf84FvTnAu9sQ2DFJZ89/XIaukOJsPO
5/hIoOnLPQeZ03SJ2TF8u7zGg1es813X4hEa/eCS0esWIHdCPZ7QVHZvR235NpyD12stt2Kp1gBZ
IxZCImBUj62E6Vzj1EUUG/8MIr0P6gWr2OOZoqKyuuFWrtZO+EAnxdWAbqZpMiNU1mvSsFzBmjVh
1RXsBkTHb8AGmIgNVJSXsFp70Pif+OuH0NcenBC/lzdacjEwvfeSrykXu/HMLk5B0oGvoHE2pYGb
RkxDT4eXi7PT+UR8H+BHLKJYlgoNzw9g/DcAFQMn+xOBs+ttdRleqfwXb8/nPVsSJ8MmU2itXnO0
PYgBYLRkojYt8FWso+JCylZGM/cd+abt5Td/Ozey4/05Ytsks+hWWjaf8H7rZwPlqjJjm95371Hl
05xeg5d4pN0EDkrMKDNQ7wvZxd2rQqicHcoLbSB9x4QSFv8roMvuUDeZFS/tME2cFVr/xma9pfBn
ca6Mo+OwnJmGf2MIXhvbNxWlfF6+8mo+EjKLWyldbcZ2331ypcXFKk/3ZtR3F9Mz0KsSjkwEBvdQ
93C7cOAl7P3SYcY1mReH0XJz6vduZaVq5DDhT2/v9zz8Pknla2V+VlMv6xmCv86228QFUC07087z
TwgLTjvUFBBS/6dHstuiA/DCFlpp/5XaFa26OFOi+slW6Uhv4nGooZnexaC4/Y6vU1t8z1rz4nss
/Q06IA+Y9OTcmbatRnwm0x29O3yz62SsNuxtfHOB4yLHkdNL1v68I6tJwN8zRCwG9iTPzrGaD5Co
tqbhBppqZMq6mxvX1rgjAH3w5CYZlwKCexRg/RO5ptT709dvRjMd6Vk3tJAdc82aWcrPswalWRlQ
SSWzNCcFln2jxlyCckThkgj0HHezwbdVeG9iyUUlTgiqZ6k3u/c3oCeapbgiAT/XsBMP4cJjSBiu
/BwEg2CRYjYZeqtlJZaMUNfCU7enZA0gOhSHG3fy/tdyuqTilkehpw5UNj8ecNU7CTxqUiDArDOL
VRAc95bt6sF78Xt/l+mkN/RrfRj5Jkalj4Bpu9eWBTa5UASkfRtEf7okug/6PV7b4qzy/RosAKgy
m3qhwrIIcFsxW6peY2aCZj2XPJ7C3XZrjVkxyQQSCpzja5eUF4D58s6dyBE302x28paEdIao6dNi
EeLPd0Mu1UDjoLINg9NhKcZ6ZYu4IGSftmFQoHe1YD+8UzO+S9L+C0wblNB9lf75qx/H6Wkh1pu9
WA+3gEkkkmXaeb7vnSumV9oUjZ2d3VLatoBVoXcxU+N/wP47N2/oXYC4NWwQyV0VFxjaycIQi8qj
Nj/5ukruBJMc8AP+hgZIBM7O1SlDVKktfgYPu/+BG6ZdLH0Xisgz+eTjt7DHHlLtrqEI8mg4AjU2
LhduJCsIG1KMZXXxMFMtPBy0XzvQSYp87QpVQXB9Zrw6zVDOML4bpYXFZnOQf82g1shXMUdT5Htj
KU6RJICFXxOYmRGqdTD00+HXwwSaKEgt7vDWhabeE37J097rwUUiGIS6eDdx+dHQLipkWQDN2JmP
tVmP2ozN10j0XmxGidYRfNHlXSIYcCTweXYytLTBDEA5ISv5a4xN/fOuejnEzT8CbAyICkHBMNRE
jF/PcHU5RcC70/I7GGBHBKIZm1VXAQnRT1ff4Tp4b8HLqNEfvpgrPq9VkvLEptVAkDQT1Ar3jZIw
/SLEV0stvcr7VaogZOAJzPla/rXMV14UP1kemo0Lh4eJgq1kFKGBO0x1wQgA0QvxX/gfdCaV5B8j
jrE0zzRrtpt6qRLpGTXssfMCdj4G9gRZR/z44JGIioQcAw4rq8vmvwUecpaSKzmnCJfg5c4i60L2
d4Y4EPCzuL3fqTetnKoZRvQ3TCFE0rklYtcxfaXSFYtXpRky5UNRiR/Ox2xb70E8c0kTNaBD4PV4
53/IJCjmD3xJJ3PbWe1vz6aJPcjnS6RJooekKsc7wv0RanrpEkoLlb+BouU8TWURo2F3T6ajccQz
OeC3PJKRvIJ2QBGSKn6/46Nkv4sm8q2azLTCh3WSnUROBJFd60RQ1AHAIi8G/uaZ2QL8u27bTX1i
6tx7NlNJhMdQeVX6LUkIwsrSvzWJY8Gv/4tGIGlIa6pb/qUiDTflOb7I09LTmFRVh2oE+Vgj+Lv2
jdlXRSdB51uOLp0vm1gwm5Blewh7M07Qoyey7HM/bKj7jaRuVMaxX20t06+ZRok+yuOXhlUWTzy5
NWycXTGlISDUjzO9L8ak8xnEaLbyPM1ObpFkQqcubxAZ4ccUAF62/58rHpJbXr33mYQsIJzDchhl
SrG/7pNonG6WxNM0Gi62VULp0qJ0He0hot6OFMirO6zd5eC0KkVSGmUm+tieEZuXY90RaezD6s06
gNomFXMMnbkdPxToKwoL6i93LNr8mWYUwWAOeFTHzvZyOaCbXgWBcSpy0s0H4tBJkQvTxtYfMy85
geYRMHyAgt4Hp/K0jvxi6M7yVlvLgJcuyjNKSmgmZAFQg5dq8+CIyIySDyopNudZKairRUQt3wbB
1ImBSTw0hsRmCl7AWYujWAyuuKTWml5lW//VfwcyxjRXziMnxdSgqMmFaQkREXDLhw4Ib2J5Ave1
dHQUXXgIE3tKJSo0Z8GP5GxcIF9q+DRpx+4tpx8uFYRuDJ13ygukojeezhp+A8zGq7aRGcbh2zJx
gocX/4w1+996YqFjQDZrm9apipMwInbo6iKfm3x7e/+5I8qkd10Ap3cBcvFQ+xDThnsApvMSvGxF
y1vrJDYlx1D3Abe6rXOG42UAgvpVd38G6H7IWurmIu1VFmac6rq5Q98B4pOHoWPfWVab05/wJO3d
dypGSjM/QuZHd9fCCaPTW2C7JXVBUjK5DCVRwbFihT9qB1AJU40jmlfD9HJ6inrCxROSRC2v9zPl
UEQGAwVx+CBHHC6XOk7jDCNk0FdD0+6qNBfo0ywE8ouqE1ByMvcQcQRNJ+RV/+sx+d0I7NDnD2Tt
ieANdY9fawwFzOiIjKCRNmUxHXr5j3VhLCSLTt5osgSx/SDknNSh7i1b7itgHuEPxwxJY0MaUOLW
/tvt1FrGqJYmqUXpcAh++7LNDDnGwdnu95gxxY6QkxEDRg1+BZF5xY10ShbMH6RQeQdGpyOquouQ
fjgvwzhDm0h884CHnZsUARZVZx2LDYgWYp3zaPXYv9D3Hw/n3tZMqJHI73InHBC2o6jsMgWVs0ev
VwXSIsE7UNVrUF5dllRndub/sRLen5AcpA1RIifka2YgYK6LOg8eQg4VRCPk/RrdbxEhmVAX5s/o
aBmRvfd5VXPc/P0ZZc3m/7nKgc+NL1DnUqfzZg3QYHpzvTd4jP6YCvq8OcUjewgjLZnKo30iTNss
59UKGvVs9HPk6XzkJ5LoDT8/abEGYSQ3oXlg9PlUrwpvz9+OvM6hfGJXrXtDwB5Mz9vYXCv7ptSs
62ztviiio6OptChB/yA/Wpg9NSq84sHapALciJ8KJXOgLax+Cse3YaTAcvD35JQqQPtNCyq9POuG
HjA7QYU8FDzA8qxBFc4lbxwzQwQTgs5eLrGoXBmS/GFofFlFe2jOcjKjMn13y8XUNRtT5dExogF7
cgxHQkxJH8KuE6j++/SPBBTOV3Yom3U4l6482OKYYPZTl23lV/N8d5xsM+x+Jtm9YiExFuWqsJJr
DxI3H7phWf8JYE1D4c1DJypA6Cpv+soGrY5t7tIpFDUZ71r2sOTjTwjZ9JCl1/QaZ0SREhrfpHSe
6G2FsJ5WT3FZkNcu3pwwb4Xo71Kkhs7zkhCQG79YxatgCptIr+Fth1+PWfQFHxLHwlXq83sntgtt
1nSylb0MiG3PWSDibE2UkXw5LN8w31CY+NnWqbejkL8bOKTc6tzh8gFEJxa5nDTcf2+Jo+v3662Z
RbZLIsmVnHyatsfMQDawgHHI04MLvehFjQrEEUv35dcoEjBwZNk+B1IqaQM27o4jdC/icnvdesYg
lkaCe7N4xT0nWMgVXoSVGyWmNpfQ9ChGw1JyoMfhMfuFkCc6udSn42Lbsf1e8eVqorDhxKufmPv6
lOjr0s+igie0S1fSV5NFqfOHO1nGmUE4SPmpvidsxsyGs3x/bfE7SXNlhuVPkuIKLSjAzyh5ZnCW
PHx2RwL7zgZJpHuW4zxGakdC5t91ruawix7W2EiyXyrjK4AXTdRCBkUR9cPy1Xb+oU56symLGkEB
39g7MlIu9i674x7RI6e6OkMS/HxiQZhjfxLO43f6c+3l0jTci0yW6Z5aQTn6aRf3zXCb/lkgLy99
R0dpjKYvXC9s/604myNlCYbuWuhY6N4kMU1Nm80E4Kno6KlDf1x1UOPO7omP7e26sfSwJK89CQMz
zDO57arnPgtKkYDuQVcUxMyMnE8mz/8YRB3penSqW2Z1FA5/0Ihzbv30eWgoDMEBQASX4d9ks09/
PQG5otjsmN13AHit+DndzNQ73tvmFYqVOD6EzPpvZL1Ifrz28j+VhT80uCU6bVGoiV8csiWHCDQX
wTN0S+tCSzj5L+lQUm+f6nuZ1n436QF6AK8gTJXXADI75ghh1lTzrGUeexuPDC2lJSb0o4U3rt8L
SYLoC0ODXpjxcov7jJyWhI63Q4P5QEtOxaTjLOKzo7cWapUWAgLu3417WP1jb4a6zakPBzD4XaO8
tHG6sSa+46NWGJJ75vj5IO97pvHTz177aP6IAqtlQrm4fTwpiYCs8v6LdCNqjDVDXwHT+2YJZiy5
E1MBHmAJWGyVBAJtyKNlrNUAhWKKeEqqdcl85HnpdLxq4mWVmE1Ss7a6+mBqnVEitqtQUHxDp7DV
DcEP35ruoWjUzKhRZUoBVkhV0fd7mHKpqVEH7akQZ296tXPm+gr469QKIxXEmnxBxSE0TugPc4ov
DhIkTmPXnvxSXBjwVBxgSsGOzDWuec67ynXnx97d7EQyiBGSDrTRNAQNEp1Df1Utnm4yMIOr7ZWY
RRyrWrlfo7FI+ZuZeW2NUkcGqHmX6me4vFg39+zRqH7V1vr0EjONypu2dD4fHMQOgQwWo+Acw18/
6pqHWfOFn87dTt+f+KhZHI7zqWpjb3IqSSWJuJsES8rc5B4biRIQx3CYbYVA+KQvo7xkwxvSez4k
oKbCzqSkJaINZNGiKCa/q0AlnxJj2yu/fQNseFDUc3qY6aKfsGM9QA4rwQoDTTtsULExC0OcuNlo
sSsLdLyAEaKM3xJydefdhmpzCg0lduLbaWKb0JIBks766NKSPrFWdPS30vfsABntofZpmQgsgtlf
isXE1imrLI5I1b3rsN/U2PNLRecRntHPQ6NTSj4qfXrKwKO+yztqwmN3YNnKX1hDV3r6axJrogPb
TB7O4QGnYgeWyP8v8tHYuUONHnK7/T22OW1Sf7Ms5W/h0Hwc6TvfZzaC6B/8McqnkkGalR+BgPiG
xSfaQEkygVl33bJhFe4IPijhslUF6DabzOkXbUsveZZClycF9UmXfj8f1gLzZuZ9D+ir+XwxHkI6
46NgUMwlCh8Mv3Gedci0E2e51E3F04Ejdjv6mVxQQnvI9pxOWmX69XZrJT0IKuySWc+7UHAa1zT2
XXxSLl2BHmReK5gwNRhpmAjNEzzE62r43GNNFRXRScr+ip4AJfdwkRjCbP8rlrK75NTTXM81XK+f
1OMUydKq1pYwobVAJT5qegRPT6fklvmqdjWRb169Dt+zLYYfqrycIM63cpzaDjPVZ5ynmtTyG6vF
VLcgQ3PFSxIoPqDTmM6iJ+sOf9OI2j3Xb8niwVo74fJhUUrtOm3vZqnO6qQuLWRB5OgpWAQu0sXz
BEw3jNjIiiICHCwJeG3no+7loOFoXwuIjz/WXyq/NCECkna95UefpylBcfxvkrAXAgw01jQIQL9t
vxtBodsA6AG7Xssq4gmabZtS7GotgjAx1OENSIpDukqkTwP8mf+/YmSgxwCM+a6HucG5vohEewT0
txyfDDX051LfBWQboZjL55Clniu7GUZNT7zT63eRqsTYijNfi/JLEq2VBjFsSagGcXBa9vTE/IPn
p+ys0/0WDSvZrXOv2zVTEy6RFPMi06zs21iou+eBaf1QXkp4YXBooUVJkcb0TgUUZPWUWYEFN+Xz
bIAqxT3waehjrip5PB/mef9P3eBNAEn2Kk8bpVNC9EfUS2GKJcBrETQsjqZsKaNWPfMqqzgeyO7R
1Wfush9ITincTwbdgBq1D6pbMKlfkjLMpoWHULRj/UDug2ZFSf1JPQd7lyhVxS4Xtg+R80bcVZoa
hpUni75gpXUGp7WIQjGAKGpatLofdpUMo6KXTUFpgOW6pB2xNyByu3EgJ/Ma0DeOEtrfH9HecU5b
d9Q3NZ+VDAvV4Fz4s1f08jIAD+dbaFQC8373MmwILHoB8DR+2fL0kC79evbIwgy3K0/uSkGzO8f1
Lsh8FNcKvvQ8OytQ8H7Qf0Om3d3CBpm/Pusmq0sahffCkernYru931HIOF0UC4fJj0t7QGIGhC+9
wuJfK6i9/X3LWIRaW+xdWEdThjFkDOtR6Hdd4q89Rolaz7EE/MuozsVs76qjZL6dHih91cEya9Il
1s23BQjd4dJEVdRiAFfs9LdZZVfeVvsPXEi7mv4Qkor6Z37dyXA2znV+tHgdDcaJ5WIvxW28/uMe
V7a2138NSet8vUJtie6bdALbgE+AlMdAD3akoJ54vQjEPUFunlOCKcuBDYttg5cG46rE3IHufzWq
dg9AypkxM6IaWe1wBY+NTg3FIu054OI3ExEHMu3W9OtiQYvFTd3wp0xqMfPkc38zsXh+s3Rs8fD1
3unjX8zPEEXVpV8zxOyQhfB8Weo7fS5yRpqZP/SdaGhDM2GqQ5b7R+aZyHL2W+xMQx1PlALG2SFc
KhWZzFmehmE2sQFWvbaNTxEzW3x8Lr5bJ3O0MOVHvMwcizTQX92BeUW/tft8Pmm0kNW8s+G+N1PI
kLU4UmQ9NphXn3+K4eF7xi7t/FnRHjDFWspv20wHrOtwJHgLc/NUfPIfzBzzAFtSoYCHcAIyiMSc
sfUQ1yH/Hv2J4R3zzNuENyZEfOUM8PpSrANaGZ7DyJ8/HVHMKMju2FAcUoh5mJjoWARvjO2IsJIb
8tSp/G16hQMQKWo72ZRcVk/gbKJhoPyUbK6BT7FTdZUCLHRWQE0EWgMVyVTlbF7uzYtjOu4V+Zd3
710xYLUkoRK/vTjad3OsSLgQKxoWUbvL4NsCRNDLeGdcD20LW4iI1nB1a9S6v9POuH5gef58mC/8
0ud4KRDLptxh9ulfN0FKhlh96YyUYdiPTMtxCNDdBvl+F10jtJUV4rUtfpGoCClNRdu5ozb9/K8L
w+dFp+vW00YhyyJ5YpVlFPsyXhH5SNgVWAUXrSusVIFZTM1yNBa+0+EQ6qY7fgFUiQoMwlfggE/H
aLB/0jB270B2RAQgzkTB2FL7xnNfrZh58VgPdlSXZZJ9skNElBzGhCQ1SgzEtTKBXGu3SopSM+kH
420fOYNN9LeoCVa4a06bY+yGcz4CAJC9ToaSr80ok52uOKb2VbrG0W2a8e3i3OOyOBqqG7l2DBeC
Z0eCN9v/LTyFyxkYgqGEf4H/AQVtcJ8DtXsq9HuCvaBjX+j/UptgCOUSfLkPGyxM7VD6HogUJgrL
8r1gKEWwFHWZeRTCz9pjGOl2TOIg4nr6MJ8Ypsgc24gLbassgEFkTXpBIrRm0m2/Ll5qbOx0AD8s
jkUZiQ2j24nG/FQdpmRujcFgaDdMIboTS7h8JiZDWpfgU91imJqTrtkVFc2pM0etbrbGVvdq+G+v
q4DYW0d/9aO7+z7qFReQ3xH8dBWyDd5fdJqQx5BFk+qMXB3aGjt2kU2xSd1xH1G9TTuSPoQk0Dfa
54uo5gBxp20NlxeSVmzx5mDdfMedAnugGDEwejGa30WXHergWdCPXL4LsO0ipct5202fLU1E/3/j
3GXdSEUuQIYIAmB0l1sgPvXgJlH+9BxsGX0iHbl+gyF9f2jBM6KQFFntUwIsLerzj1g9bQLDhW1x
gTFNwM7arZZO+vvViynzY7+p5lgfpC5SkFNZWqRXGuz2rP2ub1USv77vX6uhzMvzJGA874B5jeu5
kIqo/fZaHpxMrvUvAO30enUevFlcbzUnJFxi8n4LbtKIAiwMILUO9DObPBOPW53/UxhwzUbBEL5S
x1rS5yh+/oopH5dSz02ReWbxqz+y0v145D1Nian2z5/EmkKO210GkR/UZCsY1CXVpnluYFSpujIh
z4ABigTAz8nuU5a5qT3V1PjzBtBHXwOMdTJghQ7L1LJOPnVCK+zsUnKsPKX4knml+gksnmp7ypWZ
kEtTFs6OV3VcZ8MFGGjl9CLynRvFTw0RHN41vY7JT0x2mFmiHnq/Ox8c1S7yv6srl6RgAQF3TUlP
rOY3AWeg+e7o/zksolK5auNstIw0diFlOyLtlefDtlis2yx9u8VE64p7RsHocxtyMjwsjtcE9zEV
562dhHr4yb/bpQUeiOq8sHSpM93l1WWsxZMIeEgZcV79aAYt4yv26P5TyOPklSnADuhueynGzTYZ
MR4B5dqasZJQRO5YLJ9THG0va5j+K1OSX58p6qctQ2I8qfxYnY/JZprAFrQ+y0psukJIHPr+rerX
vMyBM6lKdjzAcqO8v+aKeVoXjbbOMlwnETjQ2/CL/dqL2B8avhrG80v/55tHfaktEDymWe1ERNTO
gvTVwJmBs3tsQ3s5puuR1UWAU8VBg3CdekWpoNOhw9ROFe97Mvq6wZLUltPDTpkCIkhsc/lhOAwF
r7YZJumAUqTJlAr9hvSMkewHEM6a869J/Xg211drsO6oJxf40fhBnrOhpxZTPHWVEb8OAz6HlSGb
LAy0jvkkbdt+KC4NEE1RVuAd5eylzO2Xs8bMsxCUNH2XYAQl4qcN9orew4GhaffFunhxG+Ef7FM8
X1peTFTH2yDwmulYCSoLy+Jh96/Y7/xJ1VJv4OaWB112Q/a7mnEBwrW9nCZKzh51TnWUKzZBP1tj
rVnEelN+hUmwd3OiFEO0L9xaWflgPBS2KHg6nOhSrILKMUFqH8YIfAZsxTeA4rRGL0Jvrqr9llKd
pgxcp/hf6BZS3yFs8MIwyiAhldKHeaeApejSgskBe6jLRIRlRmxE4Ul1AirE7J6BHP2mK8E4PQ2h
z7rm+QEpkPY+dS5B7jTJcltpxdgBoxY0n9nSFm7OZHOErxxx8zgXKx24y9I32q4EY85pp9Spp6vF
Gxj3zt5tRqyUGdN7GNvDt6UMD3XTc37oTu7dGYnsvNf3j0locpkYC36HMkNle5vddZ/3YddsxUmN
qTFSt2VoVyF9YvuWXZ+ieGOQnCf7lx5fAY+tpB9oHer02QqV+9mVi8wP0Ok6AiLyF859FGKlaR7e
PR8bDZ2rRKkLrsuyZK+80zfiOJLExWfZaPRXHM7x1Cyeg1djkMrBgVOOVPIg8mAyL5X4/FLn2K8A
HqTpGBuBh2aZFvaafyErEQjwwK5fZxvu0PvvQ+d+PSK/rwGRDBWn6JRk1Ls1EC95ZdwlsRYUCN3U
zUoUw0GiJfG6vqN1wM0xaKgtM7i6SwBfyCbyXKdB0vFJbP5hKP8WU1GdqwbEdY1axLN/7DmnGfj3
wZP78q2iercz0abrle9oA24AG5Rah7RNAU341skxTbBBuPdQPs0tjrtVJg66PAg2lKLqAyp8McL7
DuLU0Qs//yi3GbwBKqhA/QLcs0XqCamJ5ymCc83EWkeoVMEGxmSTKGNbWD9DDG5JJSZUHlG+D4fV
VturlnkNLTZNaG6Bf0gXbaEdCsmeSO1IsieNTRvkBT0zxxfe4xg5zxFy9MMpR+NWOkvWvTy3c4Tq
XS7A1PKLJInVoSYk+7AUy5qlGtl6qqe23wkxLIJTZ/dNgmZ2HXbhi93Kl/LNWZDkkK7gv/vrdFJB
9bwvh7yZSD4ynBkqMK8pwYQEb1t9PYV5jjc5vU2QHLd/OpIIDAwHvertzJceA3hsHDDDibYmasYL
iK1GTpJTxngA3vyDKZsr9tJkfGs8Zex9UG9Lejh0/YbGiMeUIjJXAgOXe76AsBJAvjOj89Pa9ULX
YXnNzafhQ9jkoeTIQ63+VXTm9ruwVkPdzx6EvccG+UYAL0wp39uYtpbK0Dvmqi6Zw6MQ6Zuf2d7D
Gv5LGlhaFCWBIJ7QU3Y2F9zp8vLj4uq2P9ZEWCAyARs9YiuoRX5RP38ZvDB7Fxw6eOdDbovcntON
lgyOeNevCQVK6nb2fPsC9qiMA8wTWSOq0JCA/uwgyohqrTRu6bH9JRV3gSQ0ERMVwJNOAMg+adEM
hPXBMtLzycKi9Rv0ZP36cQYfGLEK7DiP20Ym2UoDrONoU9YiLD0l3RLWfZsfwq1wF56N2LrV9OMh
SipJOLrh8yrsI6aXrXKvdtHzNZwErGLzzUZ4VquQv5YQ1O95JQdus7F9o2SA80nOukpPiwLFeL9j
4lkrdld3+1sb3KUqVBQ8t0BV4BaJfwxRW+9CnbAvFdrY5Lr9yQioR03JGcbks0TCJqokgR7Ji2R8
FQzvgf/s58CnkAIG7XYgUVNyeQrAF2NOyqiQYzvXcShsdEcrtMO4joQjfKWVLexYd0jTI+62meMD
9n3fhyBMinWjOnVC6Mx2SIhLlOSblm18Ip+ub3dSrz5OuXG+PE2fr1DxvgPpu4UvjHmJTFLlkFZh
ROVAO3oWqiFJ/VCFPxWvrhLcywUfhmt//ou36/coiVnp6vnQ6CUYaT6CDNcAOP2Y7tiIfFH9GtOO
ebMrvKRQ9SBcTfdr7YAR7UcAFRdkC7X87GLKVXTuHBF44S6J8IFr/0TxhRuktfP8dnC2rDEZ15iH
P7cjN1un8ky3LDCKg4zaoLuK8FXcWgZkuHJBbH7kICKkNsxPpjk7/ZfDNAFcNjl92WX3H+ATINoX
GCk1AARfYf15mA6/BGEQC/23acAjs8D2LG/1AxWlQRgJLqe8b+dCt9qQiFG0P3Z2HLCez9PmoIeo
WSzUGvIFfie4sspVxUy5jA7mZML3NvhImWWknyaa53jDtyWFmLynO98c50VWmqcq3+mijDgX382m
claZkxIjq3LWOPl94U6nCkcB+an6fcjXj/Rir0Akx/HmHs7mxyjWj7qAd5A9y7KS6EtF1iKSAUXY
KAsQw85qh7UWJ58i86plJf6UOQv5cU5ubHH9dSdYODVtea9b3Y9fD60fIbRIvCe4Wdyz1BiIiEsE
DpJ292KeARWSXPCv77uDZB3FlZTjNZeETbbizcuV8WE23Bw3wVqAAICCm0MkeiRHafnLWUP6CTS9
dgPvcMXgJtB5s/3VGw9tGmGgZ9nL3U1ah8cmTS89mWx25MxmNti7elJyyG1pihpwnXV4XrxzCSS2
2LeiEfxK8wG1xq99ao5yT2VVAFiGz7+ce1hV9oj1H/lQ2csbF+aNIarFJjI3+nJsXmap9BZ4rYBg
bmS670yUvrHuGCfGJmxOuwbdKASqj9R0NM1nYNq+yRxqMpDf5hnM8RJLB6At6iBxNo11NlNyOzsg
WjsNnEsPLbh8NBk+2UxCuQ9y1boZ+wpcJDJCymve+BQ/n1Ws3vDPqIs19lwDNllCQVGJqwxU8nv1
bqQ/GOM++9y0wTYAVqyKPYkwG3gLQKUUzVQSH7Xxh//Fe6MwKEDE6zt39XZoDBSMb16aPZeOd8OH
pgdsdIspRyEa6VhHxPvuGpmseIR7VKBHQy4WFIGNFi6xVgdOSDC/akekzVASZXQe9tXfkgaW+PcY
7ecyQSgULggT2WTZlxFPpjjCh/WXqxDI7Pacqg3e5AIZ1ECvOkwwi59OvOdgQNpMS1ft61zSG8ZS
LkjrO+7VO/1CVxeYgxKuja8FfHYNf5gMIVjj06LBgKI0DCNvjEc3enlmTKUtBbXqmf5RG0HcoYzm
AOA0Z/DdjEnwsxA8D7tMzYyToAoQlQl4A55x1rXN99gDgt412DotK8m1iulCl/EXjqw8lDEtrYYA
741SUyC2HQnLoeOifH08tX3+ioLGVA6SWKG1A6uoGOlxiXnFNU0Y1fnB1+hNPQQ5Zh5K/X5VXZE6
WIfXkId3vpAVPfGKjRblIUcJzT1TQAhw9eOWsffBlfvUSwFNX4qaGgG9cVxnaA4H+6TY99BibFx2
yjH65eMITDHWVt/O66PVMl9ab+W43dCYikMSRWODXOAZoJxpiWC1NPjy2gis9nsS8lAVamhcsMkM
SxCpfcqIF2mzMWg9XWVH97w9Tfgicrs+d49yQnKYvusJCmJNnlRnMyc2R9tlpiD12TVcxaBjVTTp
2ZSVbPz0NDg3QaCnI+r2ZJE08FXKex6qaST43wp+ncf3CQz+utMom3X15lQ21+4GfVh1VcD1IxPF
0HT1/3VaLUTOJPS+M/50sXboDrBFJGbw+0+8StczDRpFyItKB+w3s9dZir66WeU4I6/jhbTVtJuk
dQ5EJ0qoyoqVWCeo2+2uiCwHwu/2fCNkQqaJsMtgsaxsjWB1h0/8gHziHQETRcxL5jp1NP//QETG
pzhZpNEngzOThsjcYr38vTml9jh0dxw81kC7VzGiifNMoQlfvIxFepGDFU9OrNxsoYDlPZefOwPt
UJFmnO8vdDgHCIIwwnSexsTPkKr52XI+ebn1y5XDsK7P4f/A8BFoJiz8qHSUU90BrjAFuWHTJPKF
vh22ZHtWbfllOBbfjOkkWbO8qt/D/61Sy9pIJDcok08hGnGaowzrHObGARCgFFNLIFbvrz9Ux7x5
7DeR84CP6sBMGlhORmvsQezA5RSjjbYUuqlTtW86qk1zJQZbxTHGG1nhqFdrn31Q6v5ACAlJaV22
znZTk39pqU9KUiRM0aUxeYD7/JkPZO9nFUV0DlbGImpkIFo1dLiH9wlqG99V07AROIV2nHzoTdpD
29/Ijy5KASPPkhmoG/H8hHJyzzicgRk4DIUlo0g7bx9opXyIUiT0VscRIbZxZpidVWez7BBrZkq7
5yCiApa+pYUhCMVLMQwwLLfRKFFBhe/3I13UyL2+UU0vE41ymb7i2KINmJaYuze3rOAdATPalHRC
oYLgO46/P2DWTr+kC7vXrCAFM5zUskH1Lcfkoj57705pLJCmeexVMUFOPIrbp4d7psaXZbPE5RvO
HPK0tqlGeBoQU0HofYWY8YlqmyivzJuw+hP85FnpZnGLadyxvwmJe1khw2r6C8LY3zPgRj7UzwhH
PoloFjE1T+geQ7Iuj/MxM6I+cufD4m2ltOnd3M06stLIlubYph1Bs6IQITBCm31CVPrPTcSNn0I/
eAMt6JnWGal0PgPw0cB5ApM6N7YgfxhkG8Rr4O6f7Ex8uouD5mZdlegC2d+AUipKM7gcq5o5t6Wv
I6X9REJyIgueRNrvlraW0PDFX//S/2m5i2tb/AxQ4n+UIrvE9N5hghEgSd08sPlRnoRFaaQHMCgp
XTiVq3TNicDq9PCnk0MZxfVM0oSH+T/wnufxaAQTgqFC8dE8evwn0QntgMRrxPecUpxAc63WrdNM
hI/PdBGxrKiFWt/s5f6ic8c9KSRHGUjnRkC5RuhdxG61cG44C7r8n6mpJkmf+2GcTpcZ4R4/Zf6F
4XeePdlsdspC8CAVUacGIQjFAd4FvYO6osSFE7ey2eHO1KZw/kqpd9Z/UksszeQoReuo9vqm3SmI
qw94EyH3Homi5BjvfAdLXGNP5QtkM1TAF02zPF2ix4gE94NBX1njzwmL1rsNfzKia2DnIEDHOlaA
Nsoc/e2RYUv1r2Vr5JS5cOBL1WvsjeeJP+y7OerZSYnTUj0SoG1m0QLKFZWm1vrMz9x4WxMfLlgi
ld0GMbhlbW+WQgmd9KD7lHC9jXggP+pXlA5fRYZPMU8uWxCxmFYzgPMy8cPMhsr07Dw+NuUO21Pq
atgU3aTS9Y6giYHIye0jQ5JOQ6k/UC6hVaHhSevhDMSdIo7VcsRlL5n8Shce704pXZfwP3OFKaPH
zmGBofnKTAcGszFez1iKy5MMJOvziRmAkfMczVi6k7C24NEaJYjxyoli2cqHy5QrgNebhEmi6/j7
o0Gn66hS2zvhvRE36htOFBWZDPpsvq0k331mRxdwCRIN9U4WJG36LoF7m6bzV4QZbvij0qVmpAQF
Dp2xtvIlMdfb1P6ASo9rbkWKrxh/rylj/goyGDyvYWiYAboQniJL3XWlluJafReilpJtUgbO6Vwa
O8Ea3Ulstfv7tYASfT8SG7SCJvtAFyijNXB7qCEiSHt4NP4degwStnOMU6IZzUbAruF/g92QeOAB
MrwxwrBtgXo+1DhNXeYOGZKEVeqY2qbPohntaCcxz6rmfCWWt114c0niyEavUBZfbOb4vN7jdtE2
xdsrzIlvPBqtapP/2KuXXt7QX+ihYRKk/a8pBFvXgh3LMikDD4BQpVO6COeb0VAk2wAxLi1iz8y/
aSwN5l8urwEClMZeDMioRZjVHAdBq4qaedxcGi1xkhSgi8iwlE01p3LRaZ+EGHp7qCGgU4mKWmrm
qC3o7QTO2+mRpeh0Vn+KwtgKWGwf4NWXTzw4DKK2GJlS4nKIZq0qEFE1o9y7RpMXsDrRdGnR3/XZ
1wyCSFd9ZvOgkqMVRtZQubWaXdaYdNn2Cb35reAi8lnr9AeWKYGTBChwOP+zofZCvukaN8gUAq5G
09pedIclmeP8kbB24V6+ZJcbxv0/aqWlnZIICVCW8IHt35ynjzujTEPdVE93Q6APKkZmagrl7JqS
PAt2gABNG4HlBZmoBAz9jR2kfmzahQXX9UM1PrQeRilPHSFGW9QqqnUSQXPEpeWzXQcPc9oNxQ/S
IY9rh85cm1ZXBgvYWJVO6mAdPtMzxYJUmVC8gF7IWTKxMVN4fD9OprpzOxDTvGiT9HhPdbTW9/T3
XQWL5j/2lazn9fNgDC8Ed6TkVxePj/eK7Cp7LAocXpNQpU0j98f5QJ1EDu9UnNpe1tV8Y28FRA+Y
gBe028mWsn7epsmOLFlfEYS5kKQ3UQA7r4LKlarW+A4dtvBtEmwfiPp89miGr0mUFjWo7nr8Fztq
aS250CF8/KX3rc+8K99dNDR+5Y4ZaljuV6Sinz7casHbzln4vxy5+ou3cbGMt6MOsd3fi3/Q2S5b
96qanG5czIEvl8W+jYGhDSfIManMjnXsYrdlVqF3n+zLlYrCn4w8W6LgfLXEceQwxwyHG2ISHnAL
2N8WD9cp5JCKlgMZn10r9lJfwdZbzbZct2+V+2XS1VhvWbeblaDHq41SXZvE8skU0e8U7V0icRAT
5yWXpdkxR+MFLv4EvRqR1jQvdIydl9f7rkPcRLpUgChkbRA+x5bf44ptkoXWamQipT7juw0kE/oi
TCNXtP+4mNB2l9BBghkHzMxQpw8R6xWBk4MVY0dwRi9r50aoGl/UxlY5SPYuQtHA52BWGScC4AUA
46odwXCDQZjZycZlirBNjAMeYcmGI15iV0wD7Bx7FeQ6x3Esm+KZuI9F+LYsQZuiCqeWdwL5+HdG
Aob09OsOl3dIJseBPg6Z1+qqYAjysG9VulFiHlIJvnNqR4Ue6bp0y/n+GObCscya6kAowRoMGBSp
9azh/UPU85tliCUDcrkZBZEmLKpyw1ScboeIDoBanrJ3fXLRb0omzexxCBv2OeOIcw9yRDJT3FFb
TzAAEknVtSfTSKEEiFPuHxkEUVODLKVv+aSiWQ26nyRMTmHdr81ByYmiqVVVn11o8nHA3TDotya9
eKoFlW/spBa57zfJmWSiukUh+HtA0JY1BtnPhb51wRnAW6i4udXQTBHOsAy3wRYksbkIKhBTyg8X
0kJcyJpYmOIGr+V2dcJSdwW5BNqkdxG0zkchqAtCAbkJXnqNK5Zq07v+njmgaGGd8dGb4wc9Pw7E
+W5VR9966BBwn3Ur6x+BSda5ODCZWg7QWp9wsRSbVv7+5m2fWMhJOFvT24MYDRKWipOO9CCnmZwn
NHL5Q0UE0Vh4G7oIxbUVB8In+PcBMSaIBR/FsiHR8609ARYDDGOy7NYrtrOJYIGKpCcyXbBn+95f
XP9Z9VrwAG2Ptu2c0UGuLStx55hPiPxNxQOkKs/mi/Th9zC3MWdCAwBLT1jZtf2WvAGVZi9B+ws+
BmR9Y7B4H0uhBKGn0jWQkg+iF73iWS/xZBmqMCnaPDu9ndi7H7kfZI1QcIoSTSN92ZVHnc8NTxyy
OpFrpdfYPfy3yxXqZXFfC5OGW7DUJwZe0NUBZ5DcsB3X6ikPAKUgIDfv/kECzlz1fFZ9O20F4plJ
FkZmTxVW0AnnJXBngAooK2JRE4dXpkrSzLMo0N+hQHrIe8aUO+ybJ88jwhT+uGyOZon+oc9l2L7S
Pn9dqfbw+81rhhkS5WeutcekfiPY45DD/DWOSJ61OQitqT1cXp0eoWcow9AH/+rSx1j7U7zo3/qH
QFlfqVwqwcEhvOblM748QVoadR5veTV/ItLPN+3dWUG5av643hgkC7m0qjM5fd74lVet8cLgBH59
IhI1G4zyMY/1t/chrS8NQObj8rawEVd3QvKODGpMKNUnI6TXCsdzgIh69/g2KMrW3k3jlrbU0qSL
8yTGye1iTcANwHqI5cJvwtdBSZsN1ychSDjgpNZjD0l/+ABKupV4GP6m4tLMDI4GuVQaby+F1DAn
WozToiVM4MwHepzuKICyKc2eezlAqoNeKk0w35BBh1Z8+eki1vC0oEqYvWhCBpBasrky8mEfgOoP
x08UGCAFN6SrRvL5XEhf6DTBut7mONFPaWIq6yG7b9tyzh+Z0QQ+GZwXRCASHt75b3P6coOH8/bL
9bGp/TfWQDfTz7afCRKDqOD3kmhbEF2YeujpE5Rk4eiHnQpqpC3de6WTjGb7XJ4w/5dRuqu350sQ
xrOS1DUnGD+F6otxr+O6TzGdYcLjOOKs4qZ9crGFpEk3Z6y2iP6A+QaneBZYsVAHURXKofzzVw0B
XtC4yjNvM/d2MQOBd3izB8SO6y8FxTRreA14Uhgv2135/rkm6lqWZLKrGdQt3zzsW+Pv9+ytwZ2z
gJEArXQLylUcmpDQp04lR6J+b7m9QPbCHohhRmfZK0tbkSts95OowhY7viAyIoZBMeoAlkiZhbuY
aiHy7vpZC5gNCQf5Rztg8R25HXJQF1gd2Yfkuffv4knxedXsuoRztQvCQ9pBKVyOjW+0KpQ5mv7b
hZ4QOoabB654QLDyrwuvQTt3rutGBxGpD0T6nthhdXd5kIESPBV6weXMisD3TPfYAjhlilYyYDac
NGNpEmBO3c8ljPd8gPnS+/SYjo+neJK0h9kn56z6DUab0gqXJNMZdcU/ZYCj6VQNcGs4z4zey0T+
TeCmZLaMGchaVRmGIgRO7nPm5C1D6M5xhwT2LEgCMdMC546DgLc02db0erGqK19zsRFPQOTuA3Y7
4uvAxv8TRcUumF9yvtX1DBYXDcst0C2NzAmBxAGQJrGdxkA+KfsdVjpKxEqahuvNT4/pHdsPm9jN
PwXcYqd+TzHIv1diKLBAybFQGN5ixmUoG/ef6SIc5gPYXBwH99WdO3y551rnj4NJUdtlldZCGS9E
WLwB69svymePIyuvTrCb3obMZl8E+ynfBpID70qzkjD3/iHp7mmkbuWU3uzsZOV9AWYVSw1GGyUg
hX8PEJCAQVT7B2FHAUQ5bvfFD8ZHtMmxnZEn1sHcoypVUyd1ZyyHWRQ/sW7+Xd5oM2vvd1Qm8g5m
78uroSy2jjjnHEvCVD47aFHN7GO+gpNYr2CTMiKNE3KkZYCfilVAMnr3kjlbbszXiehXlD6oR5fo
0qUGbyiOpE17a8lepYUUVIuJqR0NbEKpOt9Nm1BVE5W+dnyYmz50bgoHVw1IvFd6vOlkdq+y0TF7
6qotzHbsIfT52ECSZDIW2onHJoeaMUna3PmEu2HhvDraSCWzLbRUWWhS/WKrEUgtfKUPYIrRojvH
ju7kavM73nSKhmvgOmAuINdP/L40uD13n1sUsUyQePccK7Bu0VBzYlCbzAMriEa95EgTD1nsh/az
Lw8fZkh04KCmND0zEiU3oENzmGSHVDtT6iNRczD5OtPrQgpKfK7nbGqBNWZEp9UHREM7B23JiWTe
SD3q5hjV1Rw55YrxvEqCaa2tEwh8QEb+skeARTCy701YCfaDK7PyHNAuzVE2PgKZeRMTi5ZDZQZF
uf1gb9GUajbz+t0AwCx/6upJ18GCvqei95ioHGU4rgCyEuLreIX/WzHUqPzJUtBzvc42mtu23lKl
j13Dj1FUx2x3QhLIjlQotzYH2hX6h60V+Jz5NIJiNFDlaMmxMG4+3msFqewjPjVAThbrHmusy2UY
fMk/m84FCNXb49MTjxM5YxWQ/MktwfYqrOhyJMYjyqe5Q58NVLIQBKwjlvWdXrb3t/HUSn5eBJIr
5uqCfPcayWdFx+zudlCAgDRcoHdUuIyIvuFX34Equ5IslSEjNXckIPHCKUdk6+reUXEkw6Pyz2DV
xDYKApm9OKw2Jp7mzKYOxucEd3whf7S8IiKlLh23/hSpYIzzJAOUd4TQGcprDc6NrRK0SuyRIq4J
fpurt6glHyrjF4WzTFQoDtrS8AjOaH0R3iFYspeYBNrsddGr34vFC57egJ8LjJ4nkWKZY86MgdiH
ks6qNT5UixHBH9CV/CQ80HXemsULFtLVgv0RgrOnwQRKhzGy7lm6cUKF8c6sD/VDlu8RvYGbcW0q
uqFkRkAZGN4SPHP+MFSluuoyrnoZCq2FWOOxWqzz1EKUg6ut/sMeJiKbfuiBgXFAg+WbVNY+hbVR
ZZ+yTJs5RA/Pq330YrANP5Z3c4Du4f4fCTRLMqVIz8xxkC9laPWQyLa5/pOkpvsKakpdiz0dKE0b
/j0pMq9yZPpHmGhy/NVn5xLJzt9nrejirHEOe1wityAKJB3Q9i96HxbBeRyANFtqUsbsYP6yDtbH
2sawVTUerBOFjr7rs60CYRUmhn3Qe/ccGEuGiHtWydV0VQlSSWEu6esjXzDs8Yd8tQpWmsJoNhdL
v4BElQ8mgIjX0dUCLS16OI7RzTYA+NpQllaHH8dp+I/yALqlYeEk7MfzEdxCYTaTsxDy41CNYzSw
ai1pJ7SSBPOD7DsHxgMQb5Fy7iGHP2cn29FhD5+Pq4vkILiqRu3STwsJYfuhI4WZLNy59gzKePZc
o1xRvCyP+2WIykmSAMvHFYZJi4XsM9+gch1bRMGAiFJtOdjlTPI/J+lQcCJ16oiokNVlyUHqUp5I
dNNwYYfJJT0nzaZ9UhBxi4PRzRsoEgRJOmY7ReaQPY5l1QE1ssnCi4+6RvmdMJCimauiDipqhoZt
CNBVBfFypBLzor3XuxeU6aq1SnhJgjTb+ruYRt6uAo265w1bs8H7SVmkcopgtqL4ig+Yh3Nc1Yl4
KQri6T7wxI+sSOGrT6sX4eh3enGU3IXeTzha8p2/hpNxxljKtC9EBriAtLMpv9A2R3aZ2x13a21L
uZG4r5ourn7osNK9eN57wanYOqISS6eO1gd4QOOErhT1rxwASkG1Uo2CyGjx20Qx0oNFd7B1RQfG
ohtvK1NKJ5mCgCG5X1SFDuzLTLofgezEcjFcuTxhClrEW7ETkuhJ0uuV3+fhZOllrp/lJTmki27P
fONRbxQcfV7+69PN0rQFfAb9UogIgG4dZlrUZtfAvqvEFTHKxo8K1b7+FFbJZXuhoM/HAJdH3z3R
nmucrZjOnGWBk4gl9QXaUP4it+gzsy8Rq7+mCOQwendG2jCjZcXYmGw/NB0/HYBcJSzQs0BLDNlA
gUoQejyCf9vqamzkdED6awEFDx4WXcqDpR2E28bO5LFqnjG3wuvU4muRBOQq6dD/CnwmxgIuNC2D
kwSlYFYmYKb9nfDLA3fX/xtDx9JXjD82wlVzg7/4WABW9JFiKFEc8OHhmM9a1hr+JKGmXSwyw6lN
fKI+Tg9Z4KmrAbNIPKIOyGZxDrcPUAoY7v9v6vff06JyD5hWSdtwPr7XHC9rfw5BO2wOrimhyh1X
0k4dQnFx/Ymi3i5KIFQpkAcaOFx8U+/eCkxRrPZL6qo2Qa+KdTSuAedYXr7NXVtB2RhZIX3hmQof
dlnjS8jWaj5gNMsawSrXkPDIi8VMvO+VGLyl5/GVBwV8jNELQfL2mG7HNBCsSMOws6xq1ogIeeVq
XhFzZXmuZizi2LAn5aKP62jq+cKLpWTMedFbOrlo3VdhMmqfPq1oJGlN3sRvSs0dFXgMrSIq88PH
hQPdxqoImY1gEuBEPtv1UIwGYH/wZbAJrdxJLwGsazsdX10NIhWVNCRssoe8dfzFPgQzj7be1opG
OBb9EcbI36ho6hQhlG/kh2FFv6Su72DxfDdqRDZaAbAYJpApL/Ri5fmQ+MdQBdj/JBQJdIUzuK1l
G/9TcRrle3C6xfFpTs8P49ibwEwOS9tSK4bv8p2yOcByLg6U3pP8oRXxp6xcm4iEe93tcW6fILDN
8944L4Lk55F8GzazjjPQOav91eaUDkWJEfQsq5iHcpf3fhd898JgSLOuGMVwi7SUrKATULLmyLlc
6MckPpCOccGrdizam8T+L3umSSxQGH5D9rJeFhZYxWZTxU4kfBDaU4LCTD1Nn57MGsu2KzCIRy/D
N8QKHbGPt368+2wNu9JOmoWeb9+vgIkW6byNp4q6ko/bWQ3dbXmUZELBg+jV7UwgNggkfDOpwPo7
BoZA6OATZo9s68McYwKTGGmyGIbrGFEjs1fPOYEdzL5Y7M0JA3pp/EJ+Z3RK6d7pU6Lhoa8w4jis
KIye3Zs86V6WkkVNa2iRDc5AdI/BH8mBPxHA/GrzzNOKDCMVikKiP1bxnY1j9J8529B2FtHrbUeI
gL6K+8UMHmhRHBfZ0n4ZuUfE1jw3jrWeUSytBBHrf5PiJDgNN0Kh1dsCJOKnfJYb71nu9lXtkhvq
QshfZ6CuK0yYMqh3g+/rl+I63+ajdzrbmHJk3Nf9iOP+PCwme9l/zV/DCsD+D2nxnbmPo5/pK698
X+H5lCV1eb/oYWzNQh0gZryKFGzicn9nhuVP9h0U/lo6481vf9GGis/c1KOfs57e15laGAIZ402X
0b5FKwxY92jgjxN/jPsUXOdiG8jCvWZvPwfT0vOip+2oAwbaSYge2atfO1ym0WzHGg12Fch6XCaM
FwN9K2ZvybreKYas1FPwm2lkW1VXtfsh23+LB+mNvhh/uG3Z0jbzpc3wsw72GAFNJFgVZ8hQVevW
h9npNtrB19R3ET2JBuN/UkV4X2v6BCYDOfwVk7orKea/VVJvAbkqWeVacz6Pq920F4TRVrxYhzgh
xJKcZA/d9yzMzskNLssYBfRTpT17d+Y0LH9CGeEYJFiKaAsx1tMKEGnE5qBHX40gsvSpSKJHoVb6
Y+tSA+SitA9b9ZQan178VVPVi0Bgq0B8SHoOYl/6D0Iro6FKps1klRCyzW6SbSNlIwuVj0II30mF
LlzRH2Rd6PD7qCUHR4Ma/EmG+w3zyWyyYrWVwLw74esDinVLN7+dbMF4xXw7BlB2IFNZvvADJDV1
LNpmQcET3Y80YkriAPZDPJo7BEMPRgIvnUyl0gCBuUnR4RURlkUbw8dzqLWnFId2E6hY7BtJ0OQY
5yBbPcTS5bXFHU22u1yafS3KqXBGY9pXMeA/nigg4nMrvPt1aQ7oc0d8BZIdC0L4gh4s0+mSD81d
aBaBxsNGEneoyswwkVcyORQ7ZhW+8gp9+a9loOqLKU2VowKXqhTlwptu3HFLEVmodjYUodnDjou2
ZTOLvQSZPFJSsdWK1HX18Jy5uRCriQTN69ZIrVXPc7CfZ2AmScZX1eJPVnT/mpWVJcGV1AEDpr2N
pMmVjTzTbza0Xqidfc5cWPzTTw3uCx54V7VvNZu/rpJcnrrd+t3sXKP2pJoDlg7H9Ep54vKUgOF1
705sfCZdJe1O4kX3QdIvOalC1kYEDX1d8ITRjlgKhHFpOJp77Srel5I9h+wHGH/wy/Evc2fp1o11
iCbme03+jwQnkXRVj+FF4QlKMW9rTLUHfCE/SqulxZikjO4ATLw12rVkutEd+pLMcAqjzmhz7F9q
Ggj0SGXOEG+fJ8J5yJe0gGrh31brnGIs5KDev64UcL3kXa3uYeEVP4RamXqsmG1J+lrXmHqmAbtq
eqNaYhH7AdyTc754DKGvQYY687k0qw8rrwuPh4nHTEtBt+XO/K57/owT/oJHDmPUcRb9ujgFWXqK
ZCuIGC08vUMmE4JxmqnTINZzE504AEyD2hUQYiBX/UPpPsa885SJxFMVwC1Zx+MPd92/igJEVivc
5X8P8pI999OFZgelTPPbsLxDdvdm52WYz+rNb/EKPFGHrYfIbg040bcfbArMZHw72ItnTLzEdi2l
lx2FxqfWx5anKM9yE65BcVEu2U6lTV2oacK8+LNcrUHbrtl+kFsfHC7YxrWRfQJmMzGEBTaKEMfJ
xu3BOJqtwgmp7s/j0MsCpv19AklWJJadROcmLmxMMQI8XcPLcqx7jTqd5FW7Rldwvu8CX/3qie0A
hpb7JbJp44dgHzsYx7ulhNlOJ3dCEuQkMocZv8TO0jvSjjMBNq/lvHzSZ+7Apjk/XNKbT97WnuyQ
7nAzaL2gMtLuV834uaBKos4pnCQFc1+ZncujmZju+99mqGwKBWRBrwJl5oiLxsm+w01/OtTLqael
QminErCvNamI2cqtwstpA6Xx+4bGbho3JismJzTiEe4q6xtWQgfBc9mdHD+lvZ/mN9qwRogLcFYc
JwzcuTBBD8XY/l4RXVh1SXKLmXQueweMPdxCC+74mY7Gs0RY2NpRS6s6G3oJ6pX69vHTAQcwbx+w
2OSVmpmom/n3jZvJrf8KlO8j/lvXwj/9LwRtFUAJpiUbs82E9UdCyqE7RGqxoqCuQgLRY130b9q+
084SceaZYtAvEeZJnUkRcp4b/S+51SezPmrrAb4E7SFcIqADpk2F4DuK3Y7byu/Xv4Us0rZ6iHIR
+dCwkIbGXTbopAOh3c3KSwULnuhEBZyD9DFH7OoZOZVHbZYD81i24OgsjApX5fQXp0YZrXiqfZT9
WM1AheKWtjGKLEXJGaGttDOqW0/4EvaeI9zb9pzAhyD7vyNdghWG2oyCA8ij8Mu9EwHvADfXOJWU
TueGDULX55t9XyNZcQJHjXThT8b6xIaClhdcL6bUl2LfPUzcVqepMhJ1AnKxcICzytJ6tTUPhICV
a8LJMVV0q0+hKHVnr9a/R+7LCDBcrsNvWMhoIbWiskBI+K+CnUWGHpLMRFiLLNyj8mBOt1RN23sH
Sfi3IS+4uviMpcgVM2H+2dKVMxzyH63M64UOUCYV5kfQf/QYz06JLWfnmij50S/Sc5Dasumygb+x
Fpij8dpPXIAGh8GDphvfZLD2hNwfqmguvXf5WNaS+ls5+xe8Vi7yy9OFHe5khheP9ZtBW4U862QA
84n8FNuc6OgpRehzyotpt94TWSgxEiIJVlpmxukQCBwb7h9S/6lKhH8LQmnWKykoVp1rhE3r+Oqc
IXaVw7V38wjIaWAMk/cbLmMB8c1UPFdAafGZs04hEpcOhSQtikqDGWwVlSZmL9dvu00LCgoZD+Wi
evv+9wBgoVc8LKxhOaUFod1jFRZO6eU7gku7K7va6m3lL3YcsoNwQ/THo3kwDBmL09QWShePtx+/
7XV50PZ0Fs44/i2X6CYDM803VJ3X/aWbvzovb3E57xjjkdY8xJZS877Yg9DoOQDeA9zxVsV5XVx/
17lWQMDGfI9oPLSCpOWO7BvqJJ8ZXYR0R4kK4fwFdF3F2RYziVyN8AttabQRJKCUYfNlasDy3nkL
y3WaPouAq3vw3OxNmeucOF18eVQ5lD4cVTuPCyH7/qLsz7FasO3S+FnZEX+OT9u7PLcCCmVrVTQt
4saE0hWjD4JOGd+lWjQ6iQvx5AN+AmKkU0HSARJQWWEgEYi5PsIM63qwJVMkDqP9TgBT/XEg4nOt
R14otsij/wDE5o1rtg2P4a3D3c4MNVxSz8P0vpun/2EGZfN5v4TEXNQw3tSHoZ8UKM8x/9ugR9/v
oLIq1RG6jYtx3VcJgwSY4+sUtFjgwS57j8WHpH3r9BxVLdhzJcd7KNKG6tCvCraPla+fLKQdrPWL
Y8u/i6d7XPANHO2vcyhCzlNFLdbKRej1qY6xMi1EqTznOtcgQ5/0SQoPv0wk3eu4Uk6PQBvMCbB/
U+oFYTn+s9EJ3jOblHUmtZ+UrlB3XgPAU+IIpB8rZVGFVClXGqXMYRYxGx+Wfh3xpSO9H1FWuYDo
PIC4xw1/6M27FYPGhZNU8NBoua9Hte7VQ6byDsO3wm9MpV/d6xWWbJp9e7cS9Jhhs92ZU0glxinD
Aeo9yUD1kmCxrJdSV7wSqqjNMqZTsJea35RyrFON0wcU4HYVJBwfEON4oEv2FRy2o/tMDoX4Y5uT
JjIiu0RAWkf9LwUnGJWgIgeTt8F+txyOb5Kz16t9jlsb43OPz7cvJRidHNdTdeRg1FT38+UJI0op
zrU/JqCD6Rwuo3AQeSN9JkN88r8vngkY3YSxd6DreupofZWgYjCJj3liGx66oeVuTBB5UWGcDC4r
GW7Lodgm3F+vTAvpIGAxIFlAhbxFj47wcHmV85jU/2rQZS5eWTFDGrc1buBk6YgTNpu0DLtBP/qB
gmGXy1w7SKmlki2TU2XMgePAgZ+F9lJq3+ZYcEg3tzNL7sJUWQRcP6i2O9F/6460C/x8lI64hYof
qlo2cWnmC4ekqDG87qbcqJMEu2m7wUZJ1a3oDraluyEVXyTZtl815imVuK7NAxD0cd3Y/ONNHqDJ
by1BSJRjMtkI7YGllK+3N2CgvFJtDS2q3gTWdfqWpbWvl5meZ1TYNrc0u7dol8h/m8QLIvj9G9dp
OQZy/nGAG3jy6j8PlsG2/UwhN/Fz7axsjmAkfCEaoGne1TqJnRqxrbpjXU16Hum8rznXrIxf4GaU
Nk8Zz401ZXfhGgENcYIK0aVT5Np+IbE9PCL8+A+9KYNtS6qKU653wxjwLAQPpsT1gWZ7dMYqserh
pJNfJvp4SD8pnMpbishraLSUt+uG5R9STKmX40a8nRoqYbeSb/NP3up5LnyvYGWXNX1NDJUKsZbU
G8fBcYEK2brDhn2GFttPsZXMe9PMw8MFiL8o09Mqf0gcihmXwc8HTFZ3TwglqurCjpDijvfGVDVO
U/ubfMG5wPcmBblzl5835dmW5vuYYn99L9xcbeI2VHzziBcC1htPSbo9TuG+SwSQG3JEoMi3qvnO
al2dAMRKgFGKlj7j0leSNI4ehdw22xJyyO/LEuliR8RJPHHShQNbvJPxwGrDCloOF5jBN0gtinpY
Z9DCTcqhJd0qIRrWnXJAPmER46UZEJRRKJ8lLb0+FUIUH67eS8tZltXgdqzWnOEpKFnpVjKfPntJ
0Of/FTl9riiq4F8AvNe9paluumr97D+E/rtnnRg7dMjHv8e77THB2VfbKQsgw09qH7Cihfm4+O5b
mpbs151yfOPk/bhButvS3S38rjH+W8D7ke52z2Nk2+Pg7040FSyhARzVp57S7cX8XLGlaWvxuQwk
3Gwfz2h1zH5gZPssgpICBeoS1p4tCvXzpi/Z+MaSUYcPW88dV5cyGuI+p+Ydv/72IGpzfhBq9/FP
gZTcy741fLN1RQAsFKl9lWL8u0Oq6AAD3frt43ZLnY9ZOUo2C0uQTz5gV3rxVxPVqyKSYl970XLM
By/vK7cRMxR0vS/wajRR1SB5vu4rx/lUprqKTauHisGDk45s9X3pkwcbAInoBvw5ZXW8/vY7A1NB
d5GbrNnsDjQIih8Om4D33qhiB5hi
`protect end_protected
