

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NBEaMs3qf2vRCt9CFTGP57HVPZ3VcVCIDCMjXDvQFwX/EmPbB88zO7+RCFEibKSnL6iB1S9uRUV8
6fkjPweJ8A==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kTW8HzSs+TK59Udtx2nT0jkDmTeoDqv9kR7OeIAboT8M9FgxuRhFueLgbroU3svS1TD46xwgjO67
gjud5nWulR/xxnqkG5XjPbXC9RS0FxG90EL87XW+/vq+VOMmh5Qm7Th6oA6IfcClHONPSSuNz5ez
EjyfMffr2SJtq38ZakE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
uQ9YYSMvQJDTKZv52gFvzo+bXLpj8FsCE7/Zl15EjVcMpzrwh1dR+fDhWdLXHoFmtEPYtHUdVU2T
7cG9Jz0GHq3MfhRFJ93/MRu06Y/L76cEgKJ+Ojvibjq8RbviK3gxA6ijnZ7LW1voPiUFPWK/QERz
U+lI9GDjYIRepWe4IkU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JfyN7w4w1mYxh/nQyD+Jk1BAD1YQkJDkWsj37Gnhut+k++yBH/pu3yzGsEfzw627nLpYj44BqrBl
AXv3ce5dfl/J/yqcmKdItSJAPip11eXnFDR0vPHZ6z2Vd8rPI5l39rENGQLuU+QWlNoSMPH1f92X
wYGKLJ8gPjFgwPmosASaiG5JMxsqwQuXH6ONZRK8zp1tQEFGv9ZfVyVMfekvuQJ8+z7Sra6BQjOr
i5MJ+cwyqOwv+rkZl2msvfENIl54Xxowc0q+cAKlVH/SyPntvhalXdVNHvBEu9dRAk4dPnqjlrTe
B5Aq5+m96pfONqv8kPqwgyfUNG6EkktCVigYUg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iQHmyIgxxlgJ32N2NAuClrJcxSP/FFuyNYxcCJHEZrwYdlX6KwZ8sUoJ/UxAPPzxyyiUvuVsE+Gp
a042I5zfBo1vSmsLsShW7r49tWICzld4PXwCm3rW7hkPwcGa9dId7xg1yl3ub0srhvb8pcBhli/a
1bxfVh5blwx3Vx32jWOm6fMWKpKBQawvb+RsmX+hMCsw4IE2lRuSwS00FsoMxkR95wvcviObCgQa
KrN3ili2Xr8IpDiZW5yiP6R8npYI8La2+z2kQh0jFrAT0W0SawlE3rB/GCkxZ8KLST3/CNLW5p3T
6VSbCP/kVOJ3Lqc6V3f5OJBrZ2qJAosHKzjUdg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QZOleoOE/U3kW4+Rb9J1mBPE3ap7T5ZkRXRYHDEf14UtoZXkuILnTdXG2hYCNYR0tM7b6Scfnyvm
MG/YovfRxOqawHhIk+BJ6+QyIsS9lgOdsOzSAweY9l81dyrkTgZ4UG+xzydnWVLvZKrH+Vr7jln9
VWgNHmtYuaDMCgXx2CaYRfdyX4g0isygcG2ujr1iyneSg0TREZSvjMUpzK3Od6BONp9hBynnLakX
Kc/AtT8V986EKKGglNTGNS77Xp2/p6u0MPUpWnPJnPYBAbn4TzFgl8puOZyHgHXMivYWvHJJ1uY8
cME7QLv+iwnVVV9BLtmO/rSOhsc6uN/Mkc5RvA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
Mgj2IR0XQTJSgHArGNkLEjNn8EXS7uICFdHsetKvxnSFnSEVroFMs2OIjw05IZH2aZf3/9GvY5Di
G0TW2CVpv+FxEWUoW1xXcst9zjG7l8dxwgO81swtaRqEfnvi4cAMrPqzjO1I+VyNw/0eUOrkpX5u
UvE/XXUoBCCL2/hEZsYpnZKv3SEQcXjFr/+UeEykySYMP7iyohHk/L4Z83PP0QG5vjbaQceTo2Gb
edbIPh78K42/I/ke8lnryRzJGpG8S/w6Lkmgnjxo7P8LqE4v28zqxXIAd2wBCBbJIJZRoYE3Sok6
O+DUSx87nTFU4lb59kBxbBHy5jLR0tUr7wbPw785YvbqImMne10FKDgWzDzA/cT0af9gqlrHdrCh
fmauuCS7qwmqW39DB9hPIyMCnt1JnmAQeYB/Seh0bVl6SbPRHDjAkwqu+k1ai3UiwsbZXZDtlm2/
9+pHSvd4aCzepPMlbeziknKZUQUSqHTN4gOeu+aOAbDi1kvDWJtTFx7TuKDJ8UOQq0yX2UiWsOcM
E51g6YbzJ4Ulr1JVwHHAA8pSqv5vLupSAjdPE/fud3ELy/pQ3A8MIN/ZqdNkgZeBI7op915q0kI3
IrkDAWPeSliE90frpyjf6Tqa7xRZ43jWxF83fZB2/ELrjXAHlF2J5Xvj9Pr0Vtz89ucTWiHkYnio
Ib9JK6oRbRK4Avr0tzS+mCXExMjDd6K+OGZ0IHTzRL8m/l8zOhp6aHA+xPthXbPYnAAYVith972U
dn5EJqZRoc4+sSMjkMh/5dkE3PUByuWWDZWfqy7Zz8uJ2GAw87KwjB1foCsH0NzEgpId5/kTd6uH
PBDmHK3Httw23hDddCdQCez/H+XTsGjoGX7KkoCHkDcAgNDzwSdsp9aJSx04ip164BSg0fM96YPX
Yx7Z3NxQ0eeCzpknhPTgICL2QsKgWOAKqZGZMFCXEJsOw0NzfnJHZCWuKvpMF12njcxgdk9KwiZB
MZoRMDrLLVGQ4SC/X1+PinqQyEDK5hjP9gLvje7JYvXTbPh/RsQzYDI3D8JEJhGeS9BHxSOknPRe
OUD9NwTjyrFTf6QF18jTaNn1LiKWIYtcqpLxqdCo0RjOypMZpgu15vgieqtSqe+BUf5uo6LFrYaC
npzKWcqAzC15plbGCpa37V1YNxOfeNh9Els1/wbrABIUPp8nkKNFWBIaviJYrdwqm03YJ/YymKDj
h2w56sdWAAWxKaSIEei2WL86RR05rFupYQlBjGh6PnFqllvg4VK9fURZMrsI89aZgPdY18n0WqWo
qkcR1/U1NsR4piP0MZOasZHdj70827c3Mgtd2nZ288WVj8G/OUTJarWcPXec2eyA2sh7R3kB3vyJ
xRsPyWfrzt+OGOZUcbpe8369SBe6qSIQ/aAQuqMpxgS2rT6n4lvMEBvHYDfl9j5aIMjJTPeQoblu
z/vxsUvO3CSjM4EspS+LQykmkum31npbw/0Iglc5pV8bpAFS4zpTglFnu8x2eGvbsRzOua9G8XvR
uyJzwussuIChKhi9Aa20FcexaaTYdIbjyfsX1ZuWfsLRbldR6AD6cIp2zeOGTGkuzlRtXWjvaqFY
lo7TX+h+0Jjf0nt5Eip+PhPft0qcjQqwTuGwcLu/yMLDyR2RIK9Ij82tTmWh7I7zzw0h/yBJrTxz
QhxillZBZkUJY3CqAUBZQseONFvmAFrtuSIgEhOSIZRLH1NOlVPWBJZUw99QgguvWIRkivfFFeqq
Lr3uRyDxVltXvvnF69+ndmqAo2+ne1GDG5tl8x8EF09tMp79fsHPVx/dEHcevdiiFI4ywMOix9mn
cu+bRc5a3SkDt3xrtFyVXoqowxHGlzFgzprnXdA81zV/Z5F7ew0F3z/sYRFlxwQ7cwnISY9qXqLi
vy+q02nQ3jnrC1eXE9tDTVyXQW2teiJNdPzKzK9NMIJIdOmqHupojDz1fU2AeLAzUoQFZfqCBklb
ex70k9PmofcyIOrrY7YoMmXAYnre67y4Pg9LqDgGy6p0FOixGpOD8jn07VhZqkFqCCiMiGGjjguP
D+U+ATFrmyszR8czyNftOcfaklHiuvbMOQqQY4wtV8luFdx3lURn+BDMWDazfJ+nzhg8t/SdUEiM
x1zD6538XxWWpmf49cVet5LbhAUjDakYQOiWdcYaJuP31JGUB7L0T1Q72esOMqeTZdn1kS/3r9Xo
Fs+kEkpAGsogSvWrEbRGXmY4rJbf6iSSpjEkMWgZ405jbiApuL0ObLNAcOpTudKWL3lmfW1uNHdx
7gs5hScqq72+MH8EzCYBu6ihw0f8kOy5R+xkIa1NsgnxfIyhs8dQlXaL88l9RtmDPXJjfgQ8lqmD
80EmO4Qoxy8sht9Di71pEpzw+44oR+Svlo4Uc6YSXrzsjQ/2tGjCD6fjFPb6lERoDU/PAi1DzTXR
j330VbzlJ9Aen8x3QTmrdNUQECISZ8RaoA3TOlHNohxyApXNvMOCkGNKsUP95TGKlUd5o988hsVq
AxzCT2QR8TBE0n8cqO7M68iT1O6waCliyyTqPF7VEY2LYaARZKz6pZD41Hv5VUBOTDHeDlrfauKA
xLUyGIC0/ad3gYv0IdaRFOg2fsIB8lKSUbWM1WTbTa05eoiIfpctojg4H9b8l5HLrhO5Aybw3ErO
g5Erttt8Mj/uvZNKh/CrXjj2lL99yJ4W6p458STRXiwnK2jVXMsHWgbO95PalvMggIvK7LHiMqh0
qqBJmedIqTlVuywYL/Ds7BMIT7rmzuD9+DblNcu6XOWKRqryRJCFh/mU3lR4jmRWf4mYsfDZhV7Q
NwXyhGwCmkjfwfjz64W3XtymftTUpY48P76f42E5hTbfHm/tFAIDc2MBCXMXOpzxQGXuqcJDqMcX
/uOBrP8JnGKDZ6B1syNeQz4sVM7VVhtvAdywTiqHrPnWRHG1/HcdGcrjKzhQAfISryVueb2/T27D
HokFd3J8q+Ft9yhxwerIcGxTtNcGcz55oO/C9aGhBfDmmNOn+5VGSD0BYtaQjeYNTwSsjCHWis1s
jRm9z1uJKdY3gEh6bLvDDDFmnd15Z7XK+L4XwHZejBxObIATcnE1ANva/Os3HxdwQzXxTHXRdou3
4HWx8uItbSuJClYwCVKOG8PI6ONB3UxmmwKvd7d7Uw+gmWQEDKbeqLX6pmh7Nt+V1lcCF7nDpGYU
pTHSV0EEjxSZW3WT1nvw6KbuEFp/41dL78TuAeuk5ddCqgJVFqNBFhKvcRsmXipoN9fNm8e6YNKt
pGbXvQin2+1eh5R/j0vv4cAkpFh6vSJYQTcFPz82JmjTo45d38qg4jIeGRteF2kwuJzDhsKkKjd3
Y+/trkgC2SaLcZvX0qfeogzYShAipRZeNQn5oHgeqZGOAyx8C12sWsK8o8VBN/XrJeL86+pkdvXR
EQjpl0oLPhF8gV5sZUo4ToYY3f2odL1Us1ynrmYUbS96ua+PxR+LQJ9X/aLI1s8IefDhM1lmgTb8
AdsqadedsLSbQYj3ZALaWSFKW4pifakmgSPqOc2ifgKEaR969tJxdN1TwELsiko04FeztPNzz3np
UrJ48yFtKAeOC9sDVtyirvBpuVGDDb+yYONRoTX0AYD4x+NULMTo8WFBbgQ8YVruX2BNqxKPlgg4
PU08WubzZA/T36f9WA4e05OZc4/Oh8CVrWp7FlSSAZyyjHcu00mfEtcz6T5mF2VNxJA5HtrBGmCY
7EQZpQouOiBf9qErtrmlsnLsnCub/q4aenIH9pPTiQAc7Kj3uxkjwSJb9SS5ckGOHcn+aqC9B7eH
RGp92XWTIYqMdQ+lVveByuB6zgr1n8jjXhxSDebFgjJgeeaqLD6m3OiBMd0dN9uIMD34H2icnZnZ
W+o7qakPttRymb+YGj6Gu4sQ3PLxrB2GOtZt8I/PpFhkF+CA9tqdfGlVSkAr51g9MpvXuR4XbAgO
gjyU6DMP1B3N1dtEVXJazdKfEaEKS++zD2LB3rFbraKExshdQB4Auvcd59/Tm3LL9fMGiJNGIwgt
SOTAPhFxCZUUKUcnY/5dfGqf/jGcZZXSjrGmyRj9vW4BEGH4zuQm5R7vJ8uEkBKLzs6ZDSafxdr8
iTuiJUAotJbAvC5ZrKfsu7DVUtk7Zg8v8fGZkHVs9EQRe3PEW77rfIHeEIz55I9aD7MVzQfWdSJ2
vyktKgDhGt7KskkhyiZ8JFX25N8y2dTLuC+kToAsdXfi9wkFv23Ha32Fj2iHljJfkE/LV+iCLLfi
vZf1cC0n8btICJgjYqWLZDKaQMhVPeSo8wQ9XHNZAx7nKDiRCMhW/siZNUvnkxUc+THqebmGgNci
OYhAP7HnTQoxM6mDMffElgAHTbz36QADwVHVHRcYFRd+OILPyNkLN8HtjK+RxXNes7QP2/oBxxPV
fzaUOVL3X9YQohsMapNEMvEfoqIveK9vMX/J82P4KfR1fJM1ljNpfFNi46gxsJBrJa317riMC7Fc
d2XvXpV0r7wcZoZdikarfW6fqQW3HQAZaSA0AlFQtrLzt8Y6RkzNaDy3U+deRwARITb3rd6/2MZ1
Xn3WS3IcysNxR2fyPDKiaU92oMgSHcdTuOG9fL26Ge0UZG7/MTnSs1SJvvg4QOm494Ld1NvbuIVl
FnxhOiGpt4BuU35LAsi5GAZffgzFbDyYzxQn1EHpsOZYedtaXrEPi68ZZWU7MwoyDZ+/8S/SoOxU
rdiLTK8d4gZpkfBU3bKDRusrhLP4u34U+rU+iKFTfymYYiNYYxJwaduntfWG2F6fMisYfHqWhn4a
k1IFcqiFmpaJvYWn+q/ATq6/Gu2IzIaqvKsRHh1NlSsQ9CX4ITs3v9fK9XYEizb0S/UfWF2A/5jE
JdXJHb2QfJ4HvZqGjztFuf6rBUShsmEs9HAyiHfMTnW3o9iVMYMNovN9CXzWdPJuZeBo1WGMawuL
9u6qAicnQlmG2q5Tjs+gIpyTiIeH0xLo2ZCFfTrCANe5JRWd8V7AssY8yRGjX4pF/82n/8RDFg6a
vvxQ0OUowwIk5MPXMqxJ08R+Qt4S9EQ8qTLkcrSzSaqnNJNQbLi9mdSf3Yh1j2rgbnto63hhAwpp
UwBGcZ+ub1NdagIxbbE/rkLX7PLm1gzVW07481sjzuxvw1NcycmTDMBDZtsHO7sl/htsd9wg0hR/
Gtz+btIrE0J8y5s0axLRz5iSaKH8Dg47jfqnObcdrmr3Rdja/1PGs5YcyhckrVsEtDYHdLngWHJ/
QLKtf0vzW7mQRyvtCFZ8K1+CHCSHJA2YngmdNBP+YKbFEktMcVNIjllAvgIABqbXqg6G2tGKB/0t
zfOq6QxD2+C0LA7oTPGCMQKap2HaBpISpYfFK/GJvkurD5tV0Xpd6NzPdlFuNSdDjsyTKt/9vuaa
G3OctYBsKHvudr0IWKFFRfeZiU7xNRKtaL6Zp6o7PwVNAzSo2cyYU7fEUMhWHcBIJKLbWrXPwlXk
JOROtpQFmvegwhGuy9Pp6dF9NVUBt4HpyzUr6j/9gamW1Fwg7IXTjCsGqufRGjSBvm6XIzflPldT
K1xZ33LQBTg5781cZxTl8sYwJL+UrZFjlzrT2eHSn97vNSWXepcVkSagqmE1J1+kd0vhSwbC46Tj
0GW9yefxMsKAYDt9uLUO9sZ6kRKpTNUEkrni1BLsXKbSKNXJe9GokZVvqDt1fSmM22pO6gqiBoq1
QckfDNT7nMLNaHTG/CthPTZwFJFcKl2K9ZBTTDOflo9XFu6hXrY0b69jaMwxCkIfAwWFl13KSdth
9xnsXCyx+qCo0V893cz7heOTHckbKN4tQeJ1fbY4/WUHvZ6cs3XZDImAmb9KAjhBB2Sf0YHAFTHF
m6D1OztmtBz/ZlVCHEGrNF04PYhZ//M4/ht0mB+FYbV427/tRD97iGJ38wazqxrH5h3l69jiQlx1
DSz9AIlYoZBFnAiVKzFlBoD+GTRY0r+bSRntgeUU2ctTjRmJXLvXfm/g+Foevcs/Gy56CsFCFrDh
8xSM/jzmiKfWT8I/bnpZEDF/4FJOCiAsQRovQc4fvuI0WZtA5KGTrnLpIfvnDwYR65RDYErqFkZ7
DcvI6gSDu7HLWVAwt5I7owlsWEquM+i+9Cgw3/EEmroxZSl+UNwR7+d6HE2xHevMDjDDeOX/45T7
M1LfpfTmlf/FQX47spdrDeafdzYKXxqS5nUt0sFOzVfPOjR1wBK91skNwzmI59vA2jjQFMJy+gAt
Rk5mZfgFOzawmDndNaH/yAW5dwZihyV5Ql76qRhLdgkp/Fc+FMSZXpm6gc/mzFlXt+623VI1bAdw
EEekR+pmmMON7KDQ7LdcNV9nJprDQU4yN9fwzicrOdjIWepDgSypat5aWfCsT+HjSaYjC+Vo07H8
oxqlIUtJLiIzidmxUcbH0RMnTgOCx9GSLkN2ctXDnEDEkzd+VUCL7aIX9DyREzg8XejfpHs1WkGO
tuijvlJqZzrHi1KyLzsU1UTkCP8aKOBk4anl85N+6H6zy6NRfbIho8GXZU9JKHpmLkCrhHDmx0ay
WQMwhR94SPRVBgh2q70BlIQTA+289cTuIbvIQEQ0VL0C8t1vTQ1nMLouCnost1UuPu3MSICiy99e
2FV2kSws5wjOw2y4ByV7bu1f/MpcXaMCyFaxJT9QpfQATIf8RBXbJCDXny5w6I9qzMfFKhbSLS8B
qfQZ0LbgzSEE5Vvj+fo8y92sNs+qEmjf1A7q/pMlY1ogvDe2hDBw4LRPOeV2qBdSQ+zAjEYbdYT0
prlNv7N8KjMQxKJOw8tQfQu3nzOzYnj4SOjPbdrbxMGznqJJ+Qn4WARRcUVsQv2bgR1DGPppVOq5
ExglLvMTOAHZuzLufenADphtO4TWDIUpQ2fQXRcLbAwdTO6kuHBudcVlwnYck9UrF1SnnoGF1Bb9
B/ljDgIyvGoxxxlfuAgCvxAY4cRxsBBF9XW09ai2l0DO7G8/kozUvMz1VVhRhkuyjfZMpR55qYOP
rsNTplwr+V70EdWoLWel9XoJAng4QwcJ0UF3mAnk6batbh3Ss/+Ma1edcdWzJ+0UuqjuxhMGRwrj
ZvXVFLT72dU2UAzzbsKYK+UCVC9Z8zCP/fqv3DkwHBQgBH8K6bP+qYMEUzq2MDAOoJAb3Wqj0d8X
gCDfv6oEWTA2nfzs/hJPm7buMKuaWR+ltE7Im4FqXBwgT+b1DNWO9y6M3AFAeuW4ACPdz4jfWd7H
s9UxG7WtQYi+6GQWNtMD3X+sM2W6n8kxOIgoWQB4x6nZxHo7Ix8aSmBmT5E5uoF5u4RauPND5r1K
zEE5+zDA8nuCNluLtosPpwrf406EM3ceryFrkpzXQeGn2Otfh5bN//ltg6UZrrj+cmBrgAHusrgk
AWTt1yduZpydloDE18teanahKq6WbagkeGHbmEUWMX6hpUjoUB2AE3WwFL0qoVVh0PoNn0OHi4v6
Pjpg3LYoyUoiFnvOV6aepZ4YptmbaiR/I6gpGTSeFHnRkdGO42BWlb+anOILmQjtBZl3Xk80t8f0
J14SU/Y5B33G6gETO8kRTAya4+5xqRHiDlNUpnSfZln5UcZNk07LRbeGor7PgVLV7wr+Vvb7ouxa
q5svndGXbXiooF6ROjRfXzcWciV2CIHmEZl2pk8K8ra661ihgnzcq6xyWnPMsj8R+u11xWkQbNMt
DVy1pW+AIXoobB5R2qLkIJSiFAYFHMpIQFoEpWXkphzJrDHW0JzK8U3TneHigJdP+9xbETd0HPH+
TR4imp5EQdAipUwSfHtDY+EZp61XHAAnjaY5nIWIKm4mJb+aZrL6XIa5riUI3ZVa2Hr6xezBjHd8
e17bbls9xzjVT+Slv9g2pZ+VYkrIO4dabW68PEXLdGBjwzIE5U1MslnZpsUQg7HRXctSUX1JKpvH
lP3b7dGShyDH4fygJcTV9IFQYdYA2v1y6qrkYmJXZ7wWAzKNKEr90+RkNeID4/DTGqb7DyiCW3E3
PZKqaQ3/tRtDG74WbPCIsg0qliA326HdG7j9yXyr/Sl7ng8/JaU1wG2QfXlkuVvuBOZ1ooCwytTY
Jnha1z7MkD31ZPx6i9J2nBi9tj6V5wSVoZYBqNlRY+XID6LfLnfN6jj+5WO1PZ/ULW4ePnoNcHJO
kua6SHnBl2FdzroEhOes1vy3nOuTzPdUsDAx/feZ66025+DoURhYPF6SyEwi4RVF+fRynSLZLABe
E9xQ7cRy8efcSE5etq6RirHbE91TNTMzyE05WMAFuZiRNtsdTO8EWxu5rUvYs5WTWWny7ZOGvrk3
/Dy+nm2E7mRajEFiFSMo7wGi3l1CN2OIkQp/YzTwOuz3S/8R75GMl4OAeDUggCZo/DnQQMcQYy1g
b/xR6P+YT280HtvnGEXT1+J+8Q3kCRiF1J+XUAo3jNg7Z59w0nLOsQfpG/KSEYyA4FpxzPI1tEk4
yPdJkUO8PWImXR95KNBf0fJTblSTzgg+y4kVROUTX9WHcfoXe4g1XYSSNoBiug90g3YlOkXVQjKb
FMKbHMS+tB2aaKJVmWjU1pZy4KAWdorDpHILMiwTEf4bHBMTS9yKZ+HP8a2JsSoEpK0KDL1Qmamj
/l3hgDw6HZYX17kXi76cYrZAsvNDEL1RaqMx+GDgYAj78OiereRD0X+YVbNSTRGdx56JyHpqd0Nh
oVBfal8hw4W5alBwdKxeX4QSI0ABTgqMflmwbX7m/x87TsdnTxuLLbjTcQi2k1Nd00wQMy9+yp0Y
CKCiBP49i/EYo4hvbsiIeDw+i40yd2kLvYy7dGUde2g4T4TY2QJYKQBwt1G2EDYH5WUjhojmnsJX
d39/AzUmaFiXYcyMT0eDmacYl/hirDY7N1tZpXFKN5mfymGrpPVu5V2LkK9kftn9MYjOkv79M0kw
oRChoiiSMgeXtBfvWuqHCXyreSITYNrDw9q9DdPnZv6G8Z71Mw2DoUtZwcGFxrFZI8LkMAtBmnlg
2HiuorgJCoPQBPnvFdeFAWKsx15qfyyckkaoiFrDerjRcclsqHpjYdRAEo8X0L6zcP7ekmZMvi6E
UGx0Gxf0oC1ySD52VUUQ5qC9cGsUw2PxHWSQSB3yVP5AEAWq4QIG/aifXmrzCSwad2T/tACgTQQh
zqFdDFvxje6Cu3dT5M56PDWtGkHA1S/MigUqS0/euGHz2x1peoFi29J/hxVvhsoHO12jNe18drNb
Y0pogiqn+AHJ8sUEafkJYWzsH4SMWQHnhiSpiB/muHmIgJZ23U5VkRHwbgXbLHPPan6O3ODhqttQ
k/+kNfhe04PhFJy+bU/jcerssstcOIlAMEv9CZ2CQrtwqbp2mhdbrQqF0ab1E6KqZGoiMoy19nh2
iCyD9/nRi+SKVDDl4A5uk4zdJ54JnQAujFr761JRnEEW7gpAWBof/nMqU1fK/NE/G7a9ZBF2Dco4
pK6Stt2vvRREoxtZOIvzljnHPtFhJgpsuvRfeINMtlfzLnRTpH8Kr7QqyKihHUgKgplqR1OSLFRC
vLC41HCuQxxxlnoHrStGUiWaelYDeI05jhb8q9p71z+jQGYyfw7W4F6SL+s6hpX3VH0IP7N5YC/t
8jOXPnVTuOctZ6WRBuaKNon3IcqhjApbzJrsqFA26jNbNVDGItK9hUFLJX4K1jXHnnEcO2zB4Odm
SsKgKfO5flpjQaEAG4hSpBIB8UnA5KbQO+F8e6RT6DUwC1feXtUa/YWDDlQgke7EfIMCMinX4Q4j
PbkwDWfON0CsD3TUdRcZG+UT2H0WZvymXrOEk1Kp2JRrHL95Uu+iPiqUzahfwO/9oEnDXcGgydUt
KKlc+IyaXqurRe+rbhb3Meo5zvmIZH/Sc3069kPQksvybjBqDT1q8tmvM2Ls1JZPVXNJVfA0UUNC
5FEB365KABpIVjxPw925FabWTSN8oeU2KlbxaIOOx53tf9Q09b5fX99z2naMGyVxxgP39lQlopnV
RUA9B1wtCls1cThkkpPk4LGbOd6SjtKuWvBJIdEqXA9wKnvalvZ/MdVNWBxQNMhm5kPx+Hgu1CJN
Mr7cLxe10cpVZQ4mhxeTF1FPaMMOuNuFOP7x6Rujppo5bgU1D29DmcUipUVtTLTmZN52/wBemoCc
0vnzfBU2+DYZDF7zE+pbErR5ec6V3qUycgy+jfwb2qvgurFQLQQezjDS5dAG5TPdqEAZI73fGFTY
L5bMNjzBqIZTVp+Xp0FjyRYGe28y40D+ZrjxV9Q19T6JEMTrh8xyUkN1kHF0rGCh3GUvpUbkGJEj
3nr9QKP44nNIYxKfWyTSqcPyb6QEGf9qtqRYPywIxQibtE0/8eLPQ2EAP2HZKe8ldJyTrmM+JoBO
Yb+jDSCXkhGFg745Y73N+L1bOFv1N+VZm/yfelIJGXdQM4qdX0KtN5qtBGBCbMrbNKdkRYH/3UAD
dJn0Cj4Bm3DTiqA36ZsmzHNoQtvKboeGFEyRDt+NAEss2zNFP0NZu0Y3ZjsrVxMt0m6KnaRtKGbg
5WkKQ7BON2pYC5YkAd5s2Jss/0H+sZTZ04+Dh9Y/1kZbeu4rgphTxko9UQcI1RCQHVfXctB3jU1K
B6asM8cQPzDguIZuPLrspVvDpA6nkQMRniH23TItIDUWN6w68MYz1EuylW/FtG02s/FX8JSvXbCb
1CgppXGUVUqW3sNDHcm9ie0mG8G8ehBHqXrs0Q+Jzhqpa/ItPn6TSCBtAGWwT3WEdITle5kC03Qw
nRGPBr4izJs5V4eGn1W/NEw0lIS3rf5zWdANiMeNj7Zm3ILfQHhVgyfBQ47DoCdTM3KJ+8eAMgPj
5zYNrLWq7Q3RIyLzYLKl+R0euZMh/vetzUvqULlM+kuVxoUsCtaxunJf84R2iwRKoiuDcRITgeb/
bTuTF6ia8VMoEZ8Tiars/2lFG2hFEs32cAmRdIc8g8JKro53TJ0TZz5nlqquvNonsviXcyYIM2Qk
f/BRJ5Ishb08EsFKUYTxYt8LrR8SvhFdpbJCcZaUBcJMMNvZIh36bh+oEg1NZB7cy5Hj94yaaITw
cuzG7q7g0Pio/ycxD5SxEFDMnlPa6nYvYMPmUjEu3bbL1iecZby0tQtIAcNYf3nLrNJzcmtlsmX7
tAe1hBK2Fw4qCBaPk03+jCtBlXQugi5WTKUluWZCHumlkmvLqyhD35IxZLJa6x3qbtkWrygHnL5n
7uYBVs61dez+/eFee8Uh5lCvQ4FgZ72xSHlED0JV3/SUPHIlsOkJTOys9oGr1wD7Ypmsgk5zwCIy
YvRHv8N9x+5qNu3HAOU6DMPg37cgaD/Wtr/QJaUrTIZ2aTD0Tf+WG/PcnTYBEHIC9wmBJsNCc9il
wJgptvglgwnjuIDI7wIvZuNmULStnjkmVgJ+X6GPj/piRuxzSBFE8xtQDKyVY4mP7yJQbPnDuSMm
7TvE8qfbIVDZq9Qoye/nQdd1rSCAuz1TcwFz0ktMbXpDDiMMkHoN2kulD8++krQdEgM/V4kTCrkl
U4mTX2/vZE/W7GI/z3Yg1C4U5SyR8xGP4vHYUlp18p1kWe7NFKJed8I1LvitJjEy6kDHdQtHBfQg
WM6E6NEKgn2gQ1Sd4TOWq89CpZNPRbxY6Im7xPUTtIMlWF++IOdGsRoW4rcjR/PiaFnaF3ZON65o
NK39xBfHkJfXD/Bn/LDV02mcEXMHn04m7EjhEStuV2Klbzb8wvsE2vJ60EJQ5OT/eJ92dNKegO10
dans69trqtE7uyAiipzFP8JD2FCmJpcWIqvkAWZEweHjYyqByPiM41CJ9JS3QLgqN4IYIfrUHYyD
/IA6IeGcCnYV9enDAyh8vi2/GrwEsPXhcOuICdsLWzzjZ12N0IayftFDH3nMwQavslCmucAC3oDL
292Q/hi+FTr7hffSnGVYJQq5O/9X2pcPKgNReCHlEL88kYoQ22qCvfq4MSElYGsY6WzxBxOQFACz
PLlHajyVyzuJzygB61DYlRWBMDV/NnNT4SbLuqz7sJBnKvQk/doqZK5VY0o8U1nsvPeP4GhvoGii
OjQGHa1AGZuQ46hf0Rpv0aPUHGvsjGjHzmmTyZaY8K+2e3+v06FtYht/9G8q6KKPzIKMZqIzBJaQ
SBZimFKH4bCHyF3mlDobY2f2IwTeTNM9R10cciRYZ0x94Q27+6b4bLf/WQgv0t57SroESHAGCsNl
v6HoAbjuoJNnbak0ZPeu5/zYWCXng9MCF8UuAptIgs885aULgQ9Sy3azF7TkLXvlFkXOFd04JcRA
dj4HiXRnq3hHCMsV9bwjUkwwXna7LGppkPG92czcH27d+rPI0LHOzCz02nYDXa0m2/N+Fykw8nCQ
eRO5W1AgIyF+pJvCLKBEK7BLMfDi3I5TBLkWpKu9OZk9IYwh2Bc1GSCWCOOWNkEH++88YV7HW590
o0Lzt+N67NeMEkejguf9DeBgPz+c+WiXmeg/zxXY6HaW5EjJtaAazX5XM6w7gYa5s9s26D+v4ncv
3n3XveipwEkWygbUjkfugQ4mv4l0RnX/VXUevfCrOFtqISci6ikMWK+FVX1Ej8Ui54WOy8osTLER
ysM/0gEa783vcBLvpd8cyNOqA/UfZ8CBszHONdt441wj3DGJ//c8iDje4znNfKpa348R+fva2iab
FCNtGRwfB9LBHDWAJNl9jor0pQGNBPhOrK/ghAgpyyRpZxRjEW9esHkO7WgBBKejqEeQT1F6wAr7
epcaPGMac/f+0gMwHG+FTHl30Dc5VJ9vOoD33IFFgxZpQ8fjMR3Vy+txSO5T/mvdU7Z7yiyxyPrW
sYgDhdBJMKQOZerTMm1sVXHz6GS22n45sd/DWUnBK7Zp7D+4e+7hziGhyaLklw+DzGG7+qY6WT4l
erzGqm/SHJYzirfkgKPpiW9LikSQ9LJCNBhsGBzvdrwi5pqm1ph17xPd+CM5VvIaejTS/rw3TSrp
OcrA8PO7Hv0t913dByAfDLf6VnUS1O42U48ke/JHNFd2mHkpxA7ZIFNAAW/YMw6fshegLzAnydiL
ixqVffeJmo7Xy0KAdpZ3YYrw4cDHbEWD6clwzxkAZ8voBb8sbysIk9gv1Ki6unQbqrjG21Po7lDi
SvYmibVpHPFAKMBpXNdvKikWHBOnQuymUWZeZ8XXh9xiA6KsKg54V+xDmS+bWprv4Odm1UEuW1au
QsmnqcyYZgZvR6DoLJbK/ryozoxRcSBFO3yVCADJx3QefYyXz/bLZ38zmqrKrkKBp+KJLNx3S1v5
wKHnlPDXug/oTbs+ODo9b93JI5CcG0ZPpYszjSoK+hkPMkHyOJfewmF3OsJN+7V/Akz6INqCmPMy
H9zBCFKS7RfwMSo4v+j/fvB349IrseTfGs55saDWK7PSAQnUvXU6toq9W8dkvpzCbzlFswlTVs4N
f5+RWE+tc7b1KPRisg9xtpSYrP91I3TogNF+Jm66Gszhhy1kfm7kuSZ5NYErjFl/16wB3c63DaEC
Y6hqHy7jygbNHgoGKsge6bsj6Bo8nVylVMquWDcmWozbJaTVUKXqbGJ27iO6dyeJ8RuoS+r6ACHf
eWHwZKltOjkx7g+hx/TUjSKEc8WGbH/Hd8kqiygWipMTUMQvl5kce+a+7Zpy5AFkUezrlurgC40F
pOhic3uzcDJKIJYByDEFRSRKfEK7znrTxwpmkUX8nKpZvuysE2VZ8PBgc2KWixOgP3Pr0xfTYSb+
S1s2Mp9aC22DhPWhmb/eaAkP1OH16eMr54ecyKduhK9AxAH+lAhWASJTYS3IpBA6gouNHNzu07KH
+1WJRAsTMr+N8lBKkCwcg0jvKm83rv+e3eFtYUn3mKPbIGdpjT0XVuAn/h9DrqKos4qWBAu+4ZB0
BSpAlKrRW0ms4WHCOexaybvxWou1kZlV30z/CZ6f5CFHSyk0RdGsyivHPrWeOSZbgoAnUpGTibyt
W0fRk8lz9lS968K8kJNgbVUjFEqMDZtJG3/8CtNpljdXbmfCuGwVi1iuJ9ijnqQiFc/OBJ9W/M+l
PWD6o5OuNfP9ewyuikdg9rG0L3tVOlk8D2VKGDIrtQc4i3bqCSZZqpLFtE73k6KaB+kcb7zDkw0R
5GQOaC3uq5k2rTKLiGgnfEHmUzZfpp4fsjUOT+a7skPnbCs9b5U650GKrWdDnV0jzZ24p4JCEMm7
6QFpvhF4NGG23yoa0j9NPK+MckPaSHK0FENU/xHy5o0mXe8kCXYh0uSBR2G09BN0QT3DMTge2kWV
sgGhYHZYlimFWy8iUWWHWn2mi3H5Hgqmegt9A9Z+eecJu+Tv4dKTN82F6Kj/mj9wPSaR5isseAB7
5KHzCgNVwvyLUiwUW1qr4hK12yFGXY5gl3Uyvk8Rjcv89jGGgTsr/KkPsoH39HLwAV6YlrRAQgs4
uWZtinXk2JYUjxpYH1ptx+Z4BY6mxKpj+h6Ca1cJXesBBJQ2Y5IZvSDwk9Cd9nv1qxxMzE+lopfv
PnjmFfIorTwzJV/JflZfP+QVCTmhHStq4rdrZwZSyHhnUF0CC5ywYbPIWOXsQB9FTS8x2KiAq5UW
+At6c/ksUGoUyeBtyoLrPzUVKJw8lAbIr0YSixpaQWGmU/ugsVwMpa0J0IcxkB7+aUN0FKSLMJd8
WeXAkb1/dRA4ZMup6JPRBG4KqXKhgmfvOjoDET9um3tjxY9+kbdRGZdaiWf/WoMqRM61SoCmLO+k
E1CXyMyZ7Jx315A8L3oa752YRHXmg4WhlNSL+WrgkGn1h6n7O1+FZ6/CUbLFGq5lg7zJmkHptP8l
AYkwYTkGjujsnXYhJSAJl09JprWVB5w0IVx8PL0unWKZYI5SXda0aQrpsLPiJ/R3o+1PhZfHVs6C
mshxtnnH3q2agYLljBtJuMosIz3wGZ95WQSjnqbHSIlr+bdXUFQytPZTW6DNrvG+XdPJ+pnHucAT
dSHlWyevYP/2Dggz8VB7A5n57V2qdnF0fL4HGFcFpyKpzbmBP2Hc5SnKYUWEQlegC6zlJSmtONsl
6MtP7GWy8FUubVWM79GellnMf4006s5yKxeUO/AUF9GtlkPXWPvduSRHOHP2sQ/JrRSEXQlHwr89
+S9RDzbRUs+e+yeTCRaDn7CP7/d3anZxjpzjNoNnviO2Zq46slrjwDStFGSndOHeg0EPVOutfJq7
asMUzDAi0sZL5rcEsi9gywbpCF6kVO7wWMtf03FUXf6JIyxywEc0gyj3a/JwnInO2oGJbOtFIK5F
G9a4HXw7oMJ7d3xIb+7AkR2OY97tFxt+G/zG4RjwmvsWD/Y8JmcUMKGbjaA8uquj0IBzRH23TVVI
zGWLp8oLXJqqQabmqlarjQ3YyATIdNmWQ7K1Rt5SLZ9OMDGY5F9KBXN8YTJzmvM8K9uS84uhU580
nr6FhK0pzfKnyTA7xvT3Rv/5vGEIk0HYYP1BnXvEBRhieOXQNa0n3PhYT9e/t0l8dCNoTuX1x/pJ
plp8nZZkMn2YVNCccsRsmbF1VY/ZeNBuiR926vEem4MxHjJwOnwTgr7XcooRmTX1gEOlm5HUfJ+4
gBiQIyvkuiOKQ42GK0cmcdRoXEAQXJnNnpJ7x68oMpHp+82avWEgKninY6BTHeVzUkSTkTOPEwN7
kkVj346DMrVf4FfrAYB/aChAtUhxO17OfFe1Lk7qMD2A3h6JI0UvejedLEpZVgMT0E2xJNT5J/90
QL2ucOA2TlPYln1M3kiTpv8UiHWxpMaBCzpQY9fuxp/sUSySj5/3wdKDl63HIo/Ytm6TNAEeUesN
WQJRdT5Xz2F4t/3C1dr/hU+cqdh9dI7mdMq4EyAdLTNUEkVYWzjBWA/U/xb69PbafXxmQrPUSkKQ
gRIBvqM9Zkwi7LnPcSeHMlAoiBn5i1S+1I4wrrnVCgS0vBPfLiADKjEEvCWxYCxnrciWi/J5cEzV
HAvBfMzqKwru8w2XrBbStpsyINCuOoJloVrYv8R3DpDvcnNkMCxPLLEMDOazMHCisKV4lom1G389
FlUHpm04nTvCALKnSa78a9zK6KmASWPAPl4XCirND+dWw5m3/YzT9v/btLKlwVaVR8Z4VK1JQPan
uj4785XO3EdARr8GviedYC8AW+mWnhVbzOpwFyB2+XG3rAQvI11kIL0KVtnZEK4abn8LnWp2yGV3
3LvsrgYKm0qzrij3nl9TeUZNvmZGa50IOG50Q+He/OOxJuJoejcHUR78LDK0K/Z4lREUon1tX43T
NN9D7WNwy+RdNzJBHMluEyGEst0ok+AFv7cDL78kM3PiNTQkp3UBg38Y7gXIKfO+yxOsbqkMKnSM
ACZB5qurv1U55LJ4uhNmSxPA900q21yjtZOG/Lfc+pMO2/jWHlhydZTsXTchYHrZMtXc4ioWdYNR
x+K+WDKn+euDlpsvq44DNwVx5d1TRjg3pvL7FJXAR23KIcyrtuN1CM3PjL2X/U7w3G6IyholNWaX
Xtyay1a0/MwGPOImvtfKaGtZ/gPfZyEpyHGQPPXlI/hEksG1qW5rxZL99BpsU5zBAyq8l3JAcP6Z
VN42BFlNOfWec7HJCegzmW2IWBhWcuv7Di91nkANVa2TuVhmOLxWKWnriQNCTAbc0hOq9+s+aK7U
i8a0Vfjt05dhj/I/THkTieki2+lSN3ZEmeXtO+RX12yLMkzRPb9KQ0gAS9L117OUnoO5J9H1dMyn
UwlIDiFQetoyXhaiO7uhxqzNYcEwpEoakwkZ+EOAtDyQPAYBTt/oKvQ8DSPIvoFn0L9/MNSOlnHC
2Rmxo+sxzq8XsCLDrQP7s6WRv9hYL3Ed1CrYNKKyLWueWUHcaaYx42lC7vNzBeU/NwXKZ3xM5qPw
J8SlRQNjbqAFet9bxqGx0fH77+J4fxk75rWcwkvW9rf474JCvk2s5okV8elQV87p08/ZhKkmGgPo
AGnMa6gd/RhNNke5eeQaW06mIB8NtVsQXJU5W31ZMmCz8YPLvea2Y9QT+XgDRkOl85x588IKqOKP
Yip65lly6evTqxvgqccXSLSl08d0IspPljZrvHCm+y17u8nlVkQLtCyi+BdoIfEmDbYi/tWMkB6r
GY11EakiW9eZDDgN68jA9D0A6JY/vAp2HYPF/CVvaEH0FfSVTn37DNiH1nI6B53dMHzt+8uXB0lQ
VYFHieEf/ciKOifZozmj3SWjK18cY9sTcfEtbg7t+WB8EDsYgERfdubKJwQkQ0LcO0Nsu5CX3POH
Fgq9MrfwmAY2zl741WimqLa0ocKglIvisKCqtwSoi07F6hpocqf7CdPbtxmosyzj6uZHldytJnvG
E0JvG1zjdZFeleWwh24gfsNQr8ISQVRc9U+cd+PdoU4P8c8AqchTL512SwTy4yQkyiIOB1+lYV3L
TdR/g1WoOjg38D5XqeomjtOf6WSGuL6gnSOgBO3jJ5fThkcXDui3d5H9aqIZOHILCnTdnpCwY4wO
WTpTYIWLMHFJQyNLqGJxUsUw1dHK5OSXIJM99YfvR8uMnCtE189ESvNQlX8qsXGaNUnH5Ncci/y1
vHKlC/H6A6of/A1xVvKnYObSQUUuwQNj/izyyBk5r3IbMe5WPfsH2BwpgoHqmACwzCiNBFFr+qbH
GV+qW00riWXgXVE8WcskQw+/JXDEirRkF6Ow7KlmJTPTSY39LqKHzulwt0OGsofdH5v9TrbsNp9T
9P1r51bH3xl4ZItLrc50GmfUuUXwofZ7nBJwbJ9hfG55sGzpDhHEqmNkWOVPjWid4lSidgdmGFeg
gDrs9TRz5SjDmNh6PKwJBXZrutB4+5t0Z/9pzeBBr1t5HU8ej82DAtLWWeMRFrZLct9meWfCq3Nd
PtSIBjaQnDJTD/kbPZ7tMD4Cl8IrubXbvSJ70PzGerPgtZQcJvNYzf82pYjqOMKikarClb5yvuzY
BC1aepsSUyJwRCch9mN+8bmiUG8l44/7tiQ5CwTvSROpiqIa51qfXCNAkjevFlPv/rJpCufJtViK
FaTW6cLt2llFaGGKjg2sPS+qzcoKZzxqpdNM2xZiAA4VdbqHkH+jI/td9LosG0KRZuywksI3kSJj
qJFW9R2YRxFUXirIaCsbNICG6iEIMeE8XFy3PQfYZHM2Djaz2gf8VNxcrokKmoN3XhaVHZv9mQO1
BWdVqnEdXiqGnl4vVaT8ye0Q7N6vMJZxy2fe8wrV22QuER4QWNzFGUQ+sX+NH84yVvn2YsG4pi4h
UdnS4EK/CvRJYjimvQ/Xh/zQqrQnKRD6IfjF+wDh9Iy22eBp6psd3s8ijbQ5O9LTPsMwoNKX5siU
8Zhs2YivCAVuMEi1ZJX5cRXHalfQNJWCKamyRYsvGYuuF8LmiSkVps16Ia3AuGaAwqKBhJCYAGq6
QQnsEBa6cGb9roXvD9PZrAXeKx4aBA0yyicl9SQOTR3AJ36B0NUDr++egXTs/0bkqP/yQIcpDRSw
WIbZR6IishohdZyK56ZcRou5dY7DcyOu7/Ih6l14zVAVVQpXi/3EZNO7wOx61v4E4P6TulZgYv3b
oO15suMM+j1vYjz397A0MkBiS4mCLxaMq5XlnoVQLOHIBcMC1o7csr3PW9ObzhFT5RxHMP1Cmpiq
h0gYsrrv+j5wMmKJi24Zq60xXR1neTUgdwXH7DNj5X6to6FslbeUWmD09QSqVVzcRw8Md/jcw7P6
BytV0agoMRqTWHqu2wSeW/ws9h7+prUieShMDxKdIrwqKEAT7maXhH6wXEk85c8kiIpsLDiLVOy2
Wm1miKqYAOOTYbCeQKeken4OGTf8aFgZ0zYbEZryQ6ZedE5vJCnnx8aFk9i/p80brh/5/Iqp87il
3hHSUvdiwob0M4m9IWj4wpn2W5SiwpuBUwVd50dwzDaXJ8cKm8LyAsHvlB9jzBdW2rCiyY8Z5Mrr
EmFLRLw7hmpeiSFIIrIpmweT/AiiIy/5tInSK8PKkRYafIWzCi9d9Nnqd9QHKc2pvd3Ayca8OFnN
rdiZoQXJx+uiYjzA1ggPKF5W9MPsu7lYvqqMjkZaUGBNaj59KM2cCghFLeXOuUrda8QDBfYGSJcS
yQQIUlRJ4STAOwNBSoWYFnNleu2AkN6hgqNFAklU1IbN9DrODUv1cNMJk21R3c5NiAivyPBXP1bi
QSw5HzU9Y5O8A5EoGsX8dNWmxdb+udA4V1T35XPz5I5zWg+VzWpEV0nmV7Qzws0yM/dgSpwBJIxb
tr1VZZ/FgJXr1o7KSfuVis6kOCM2u88buDh1efawhNAMyYQP3frm9eeQsdsdGJqR8yqU7oELmGdL
zWPByKDvo8BZOt0x+hWoA6RIiGwKMRtIR3YEQEv0lv45uux30+P9NK9QrkNI2ydZ1ls5PHdRQaL/
oPcxACccMFOfEEzM6RmIe9Y/6YOANxgwL+J8OWBzfdmU0TqvZofcQVSsQFuz9DmoOIHcPud53MrY
2NRD3Wifd8AwszJEPCxG9PYpBZfWsNN7vK6XSZj6sSvBX9h20hr6tKPDykRkfg/s1LPYCpc3sZ+w
TPuM+SeYvgIYoDxig+s2d49HCZNTno+8EWWEtceK1qGBfOGraIAeqZBnN9Y4mt72L/5E2FL68lnf
r5UZYHrbNQq5fIbfHZWWWY0YZnMwAKe0J8gIOIbr3Eu4KCt2CyCxx7gY9ByDBTZjvKn+2yuZrLHe
R8ZJhOMl2W0Hg3MvlMrV4QMjwuu6zSm34tCRftDgJHBFUswHEXffSv+IfQgK9wptN8Pb893W+KLO
JkzwaGOZUEECScEf5pmrP51ArT9gMS7zqehibnfuHVd1m3W2MgrDBS+WbDIT4nxREOARxYPXAHDX
4xJZGBitTmd/Xw4eU+9TpscgUq2Lyr0YMMInzsTQy8/UTr21rX8/2dKP7XXa48DPofIG2tBv2BQF
LaW9pF3Qck1Sz+bASmXx42X8BeZDayM9L0TTY0LZV2zo+l3mIPWrYXuIR3x+bkh0PCtRQBbVaWsH
saN1Rd995DXZAtfWNudR8UlHvR3PCGv4cbJXyhtrQLLizRz6DJjIFOouEcN4CIHijncqBZgsbB1A
0UXp86XCqut1PBB7XvN19UwaORCk6/q9okIIrGGdvb1/Ge9BRZ2hqH/xCz3g+ajo2epNcw2xG2Ts
AOfPUFm3Hi9IoPtzAK4mk3/vm3sK52ps5ifni4gDLMlmiNYlfecBOCyvaGqra9RIAlh/CR3IATP2
BszX1HJ6UN5aniEyLobjX20EOBdOGbMm08SPkGK0IulSxsuYTnrUkqy/+TqBRLfBJXFHGsWgNOJc
vSSj+i/LtzfoUyk+Hov0z1VoM0rigLTciCmplIHbZt8hVYdkPfDD4YAC+fKk+GMEP9OmVwUR2nZk
x3nRDx7NOTfKKPR4oQZ5f6mU9UfJbJJ6fnwFAPeHp7aM4HFvWiIrG0b/nsE6C3tGMP3/Vz4H3V5i
17DlvWyixn/uKCOAJdCOfEnc50ped/8bO/JuaYWIiAJW/QmFPcygU3Ma1Tm1E+DV84+BffyF46Rw
+Aq8oYDkNqZRG9ORsMFM9EP2LWPBTPmUmGzq2nHtxxxmRBUUmlP3ijvJ8sr0T5ZtRy7I0lI0X73z
ZGfavsZUfmC42dFw6Zahe/v51HFYl/bKp9ZBAIVIXrXSglhaTIPzRvdvbMciap2ZXdfx9wRZfNTO
WIB6VbEMRMNDXfXTh5pSZgae8uhldKKp6R7AnhrEcFalQy5vmeYOQaHrM5idBWNNhvsuNDS9TFdk
kalW7GAB8sPpONgBudtVgdFW6dOBEow0KRAwBj0RJ9JT1jVMgeMPKat0+zCV+irCbQJydtL5V3JL
9IiP+KWbskmVtlRDFOfJioFCg3g8E2Eyb6Qip+ISjEyztKSMeZMG1m5fPxjOpmpq/AIXOqqhEUJ0
CD7nSXXI78rTZzz+F82PZt7PIyg4g163bAqlm5tfmfco0UAzkYweKnsqhuf5P8/pYgPQfY7QQLkY
b+5deV8P2SwAMAzrFrN/biNp0s0lSwH++WTXaTz3BxBloJubrT252ZLGoTqApqI8vv3Iozqv+/uD
dnSXxVBDQadEBXl0/xjfNBz4O8Fao92PCDDwlL/DT4sht9x2gm2wM3dwHAP6Rnez92tAxzx+toph
msAYVu2VkoIstfj7y2HOfxrSi3F0+LCY3MQbDn3pT740DchdQVXfPyIsBKGFP4tSdyqsUftM4MfZ
PM698iD9LaeBej3dzPoRKN0sFgZDdfjYoYjxjK0VCMW9jP1UTErciGBQsAC+r5xJx76pRDhsOpk+
X9rdXDqSUZRehsQEkrUo+SLp3AKzY99MK3nqB1C0AS+ijo96FDupIR/9kk+mdAqdt1rKmzh4+fzJ
mOARI2F5So9jbcXOEIMg+/A1gNVpNJxq15lGRebAgy7ZR6Oo5jGzCLIFrkDg93I+5TtHZKxuFvL0
R5v/lyeAg3aZTSBhtrjFvhPipQCN6aDx99XmXx8gD8T3SMmra3kBXpKk7x1BLKujlFikie06+a82
+Qp9+536x/pH2qDp9tTJWgY8nXUF+9/+uhoJypcdA+sqqyb0NyVkcB9I72lsQPnQc+ilVBJwo81c
xdOhhNUOWULQHhO6TmfmMEAKo7pHalU/bHoveQBm1jVVV8YuLZsQDpBI8NB2NgXYgrmxwwW2XzeC
+9Qtw8usDKeTwPR6EkG9vn2cvbuyVz7zfiW3vESoNLDySk7KLsEzQGbZNtG61kINTGxb99F2Rodo
G3fjjN446NK4XhLW4tlF/RuE8NismE+VHtZX99Ud9pryehkyyrqnCJrquFpRENNfSja4rw5tly3U
v5kE+CLFbN3x7JTdlPbJv6kkPxKKaSXuUO3fYQnq0O0XF3EB/0A/qsJhig8GLHPAEPQT8oDdDATz
j/MeV8SiQhBeSfoyBENgSsUCpXWjfI3h4fwI7jV9xcA2xmD7kGlT1W9AwluY0Aeg1AxQQePe9axu
Db5dvPBf9C/yoEuzs/CX5Kd+a6ZN8SZOE3yDd71fj8KlRsywYh5vPhaX7diJNQYieh/OOCCnj0gb
pjtATHRhKfa6uuK9BXLNpB+F+F6ZbNoodquqJJVIQD1pdy3wZN1dYeGM2wLR9uOReaZQMAwKnGX5
rvOVrqUfFboDNokEiVjcp9Ny8eGIlruiggtO3lwSA38xLcQbKo8Th17ZJXPh030P8rPJ9rvf7xtO
0/B1f0kXp/WlyGpkyx3Fpix6yMAMFGejWObPYVc1hVgOzVynJscmHzbmYJOFbnQplsqFFxoYacpi
M3xWZDOrvzDqvnHPLNKC0zVHgtT0MgkllyXkt+B0cdbQl6DgcBqkD/ruNqqGF8+gkTw+3RNUPOBk
yIb5jVa/7+ziZ7n/i17cJKqABUGBGxErbHFSj/gJ6QnW+o4owUdt0V6mTjApvKophV+hm/7xNGLq
kruMLrtpxGbjhert4vzXnbz0kShDPwrY1guXLMC5GJ1rnZr0VEibRCW52BLLxr/Z9yo/mXY71ho6
Xhpan6whWOp8R/bStIw3psTM9c2zDIg/bSxIcQSiBq8NRG7hmaOcZApzoueakjiup0qSylZY87uV
PKhUaUdtRoN/EdJER1KQiLPygVzN7waD/cVxPi7/gKgzM96wcVTCqo1o7CGmll4AlY/eIgnx4e9E
6EzRcynuPdIfaOK2++weNfr2zM936j1R/0+0hJygnez3B0BLTpaYTgfMlajvYGBoo5xRea6grKpm
yokZTwsiJyateWCMRnrTY7JyMRiXrmUZ/hq9kKD6TlhKTatyqTWeMBCPYCiC3egDrqr2UYwIrysl
cxEa2wQHw5zOjIgRHcNSM8HBkdBaoj/cUMgvkZHSztF7bQYmRDq9glBg5rUZrUkUIW4gKxPNDe3Q
ZzTPItMqB0kDw/BQVVnNJAcKLlrF/3Vh/Nb0SCiUkWVVb3xdT+TzyTvdcQqMVQWHZj4O0mfDEjWt
t8P6p0+luo/g0s0ELk6UPYYIsuAlX5MvFzuj6q8zzFFgaIZMKHmivcHONxcb/sN78Msuutf1BM6K
1WIfbKQRU8f2WO8LjCTOF6BsDxeUDWbHXTLclR37U77HU5Nwa89t+VtsaaF1Xoa8+iwHtk9WtoqZ
Hh8ZwOhbtK4ISl76mLCuJSp/SezIzcLLi7B1WE+T61vanrSONDOgSBmK7ujjgpM3qo0RZpe184Ik
0YXb1LYcyAGTMLKGCMfuhN8g0b/EQOSAnr6NjA/Q/kCGvLTGBk+MGIWX/3P71BKOSiTTi8sZdgQ3
2t3ePXtpijeQ1Dw6eo9zdW7nCebH8voIDtXqjyyl9H3/pbMnXkPR17RSqcCtMjJnNb2JEaTpbYvW
nKE/yJ+ToFQ7y1gOILkCyHKdC9BHICWkkNPejaUYkHXQouH+pnNo5HoechoReW9tN0qyquLTFeUK
fIc/juPnSXyYWceSnz9q7n2+zL30qmoFquuutQnSOAfAaynfyLmCW9lOOvw+/cGzqligRKEHFF2t
GOGbkAm7tBHBPbrSw1/cRuIHyNptQ3ZQ+7VNDhn/gZBlvDZ6/xXCSpYaQUX5qBYCO5RIGm6fhViv
c1VfiWipJc8e8VcvIgMWNBdJYxVQF/+TnQi7/voRgx+8nZ1j9hD/D33zfE02hyyTi0f8XfS5mCrO
xxlgQTxNpiRIysercvNtpePaiZknbtalwSeXP60mxcu4eeg+6yIztEXophA5UVjEJGiRG6YZbklm
T5CpZooQ8wKajoXOVUa7XfvX3EgC8bFN5Pey3GdRCx2RQvrIdGn57zXoDbYhbYMucPiSMmxDcv2p
Ib6LVDE1gWcfjOmmoJxg62eIBvE+0lYXP0vTvhUgKkzaRxDQ7HXV5pWkxD9PkGj6C8m5CHX38oi8
cP8jOSJOUIRwFeE/fpW+IMYnhE0O8KU9TRG2CsdcIS0tWQvTawtby3MHG0n4IyPy61gEazb+36QU
KdBcVNexwpmJWJBLCHO9UBHfU7T2KzQAMdiVrILeIFV6C7Vkrnb8OQPSkK9QyuIkFl+Mepxg2htf
nLrH7PtD2hfpHdTtoat6rYp+H0sfENz7Vnqlb18YBwL7T+4XwuMVnlGLBpW6OWlqh9PkoPjslRB2
mGF44ex/Y7UoSj1GiQnmsoGJsg58Q0Rz4qHJoXua1EQm7zloiOb+0/HlQixb25ZETrnKqOWc5fZb
dMQ++JLr1jUG4qGEiKdep+g5CubBxhnK4xgUT4XypbZjJEAuFnAzud4tfyfWPexCxbzF9HGMX8xF
me9CwoB9Yb/1RBPb85jlLLiv8ZLLuQ5lWTnbdSTMjR1etjDaNlBfDknwzRA2oUZ3R0qhTWldw+4P
Kb9lENG9rdbFDCmQhQGMgCpYL1BQZL9EJLh5apadUs96yxWwwaySC1+T6b1mFzdbvuH6+5FDFNzT
enfvFEWcBVW3GX7KKQ0chbel0D1cixEaFdCayLYgsKVDMg8vhP97cd8E0hKCmuXCtOlxt76gJPfJ
JPU45iAUyPCjyrlQoElefK76Z/vgMhwOTc6TjC1CxG1iZUuqk+NpDTCOQmZ3x7kZnhAX7x+eVwiD
Bsmwgt5E5EBVD0RicgMZbw0fC1Jep1oYNfwscIC0PzLyqaczzzcG3stnJs7NR1XJelmVtbQQxH6N
PA6RpOTmQYt0PlygVzRNzVZ88QSWSnFJ+7E4jXO66iUpBy6hE+2uIUeyD2Qjh0ag+V36B8B6f+E/
ImzZ6zcBg4CkYx1yO7xQndhh57yF13cAmQZ1K4Ma/lVuAjHmpicYqS4DExXEV+JDRp36+haxmHUr
lo4sBH5vBq9U6HXciyomeLMla78pfFLYCt+EzEs+BLJS363gKTOjBHVsu6ePP8Fa1VgH6HcZF9kc
mXg+ZYSNRssLZalTuwgj3IdTA3BdN8tJ1g7zKfZbVcJOUex6EoYxNJO6HdmJJgptHutjpPZ8cPRf
naV8nd45nlpU9MikQIYv9alexRFh3UQhjNvSkV73bfCm/TZDSvaYC8oYDB6tYzsNbdg5EOWMZVH9
9HNDnugA0FYpu4Xlga+T6HGyUNw3lZgneyoNV/iWr8UNmOIgxhWkzczSfTzb9MEE77U9ya3qZJV6
edUeZj5oLntryGnWNyfp8LBFcIrdDbDXW696kDPH6EfWQL5Hd1erYg+xck2Cjf3kqffGCp9ksW59
q7YAFclcntQqzpNfgwugFS0Nddok53VuwYTZhqSB61iJh/PTLB5A7Z1S0HMskaTTVPvZGkxaJiS2
ZDKRXCByc0jhOnpOBSvkO1B2tfbXatR3wxhKr4pI4UTiP7tuoHGrlFIrBd84K8INnNN9oOPdV3aq
Ykgq3Ac6fr5Yda7UxBrvqsG6cQLAaCdakgnp7NAXOK4pkcHicoSsfKpJq9MDweFszNzWjwWdcNx/
KR1MU4AScEGebh3CBMDdS0yZjaY5RUj4w9kx4Of+FfP2rULA6ivJOwqsd9Y0JpI02YFVmr4GPeTZ
32j2tiFbF2puQAYJ1bH1RbfNMHcjKIkltCSKcwayTi0UOJwHm2Kxk0FBPoYdzuVD4Zwkq7GH/cwF
XyUpYc+Os7I7D56WuQb3FkOnH0xTIddxCTx0qtSDnvoJVLmHjgDME3TdSrVXRKv+sFIMUUw/SenM
iXogx9Vs2qOVTXYdVnY89TaM0btpGhFnrKS9f7UsNf1GREFWbDWt3bNOzBjH5k4ALN93t5OYnQLb
MmH4CLRMaIKQFQx63rJ4XC708lKga42DkxWC3qLr6jtQW2t3AElquuFrRunl7+eRCVrEiFdhCY5x
zIpEkMMCPGZInTcpWjzv4w/fM1FNbKJSMWi2lw9JFmdbHe++uTSF7OzOYTtVA33J3aSPK/vDAJ5T
4E/THWWnRmO9HwaNu/43ku6hADfaa1+NtGc5mLMGBH8b6gTRgriZ0DVwbqk1cm5zTxz9QEZzZI2G
t//qXkwxcw5kyGrMqjgyG9tfMnlKzQi90X5d3NkNKoW510fr0/WdboirERZeIHvkYXCiS8uLapO7
v5u19VAEjZnh6D+UeKoideemVDl9iWW/NgmXRYrCyE803XsXGBaB5ADrXdq7rpu0IHAOtmBn0Wc0
oXYwE6j6BbPDAkgRFh0Pm32z2ZbNz8mmAKT5cwTcT+mhE5rPvMhgcdfT198ur//iyCuA8xgbFXDd
l6MqLX8JR9i/41FqvwWr3Uafcr1yXC3YsZp8mty/yUA7eWdYqF1V9fYXluGSHleBTQy8MgOWtBCs
v6GHF7ii2KkYK4L5c1ozOVAU6CRF9iThVT0V6nRIU62ApE1X6e2Rw0jbOup/5wNP8NxU6R+g3khb
mmbbdAzfp8Nqk78x+564i+9EjlkMVENejq6qT5As0j75Qoob2q3pI5Inv9xhnPDe190V0XLQJ1Vs
1zMYOBJB02OR4AD5Yk/JSckI0ZuYVxfQ5xGR4MIHaG5m1BlJFoJ720yLEP0WYYvfOt9Qxz4N437W
yXjtUHaMaNMWT/5lDIVBCjjQ57+ma7LuH4heONXkW/AZRgXzEL7eZr9+QLkIeO92JjeQKNMx8QOw
EN2XQ8p8SfH2xknMWLt+6QIXEzYYw6x2qTvZ8bUbwPWeLa9LZ5hzZWYTGgJKLTdH31lZi1wIKs8k
cMw2GWqavKMRUPMnmcL4cs0r+qrvtX+un2wwPNIZbTfTdbkctvesxeYiTlDAISuGjcLyJVY/akRk
7yoZVMu3PCDC4jNZY8BsxcV6wPY6ItSY0xeK1SpsRzOexqUpzDmz5WsCxCLMQN70yGY16HRscTg0
ruXhw39DHlXe+vXkMpOeBQQJJr6JGl9y/IpVg5EmOKEzU2Enez68DLexQkRmuXidOMXTEltbXc/F
YWYn/NGtV3VsjjjscXiFXiJNql9KtMVlPWmdm+EFTYtMJabxIY6bHqtKqxhwx+bah4c5GT2PIvWy
jbhm5k3fnQ==
`protect end_protected

