-- Generated from Simulink block Brik1/PilotDetect/correlator_fifo
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_correlator_fifo is
  port (
    real_in : in std_logic_vector( 18-1 downto 0 );
    imag_in : in std_logic_vector( 18-1 downto 0 );
    valid_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    real_out : out std_logic_vector( 18-1 downto 0 );
    imag_out : out std_logic_vector( 18-1 downto 0 );
    start_correlator : out std_logic_vector( 1-1 downto 0 );
    valid_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_correlator_fifo;
architecture structural of pilotdetect_correlator_fifo is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 9-1 downto 0 );
  signal new_correlator_ctrl_start_correlator_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal new_correlator_ctrl_count_rst_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 9-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal fifo_imag_percent_full_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_imag_dout_net : std_logic_vector( 18-1 downto 0 );
  signal fifo_imag_empty_net : std_logic;
  signal fifo_imag_full_net : std_logic;
  signal new_correlator_ctrl_write_zeros_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_real_full_net : std_logic;
  signal fifo_real_percent_full_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_real_empty_net : std_logic;
  signal new_correlator_ctrl_pop_net : std_logic_vector( 1-1 downto 0 );
  signal fifo_real_dout_net : std_logic_vector( 18-1 downto 0 );
begin
  real_out <= mux_y_net;
  imag_out <= mux2_y_net;
  start_correlator <= delay0_q_net;
  valid_out <= delay1_q_net;
  delay0_q_net_x0 <= real_in;
  mux1_y_net <= imag_in;
  delay1_q_net_x0 <= valid_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant_x0 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => new_correlator_ctrl_count_rst_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay0 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => new_correlator_ctrl_start_correlator_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => new_correlator_ctrl_pop_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  fifo_imag : entity xil_defaultlib.pilotdetect_xlfifogen_u
  generic map (
    core_name0 => "pilotdetect_fifo_generator_v13_1_i0",
    data_count_width => 9,
    data_width => 18,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '1',
    din => mux1_y_net,
    we => delay1_q_net_x0(0),
    re => new_correlator_ctrl_pop_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo_imag_dout_net,
    empty => fifo_imag_empty_net,
    percent_full => fifo_imag_percent_full_net,
    full => fifo_imag_full_net
  );
  fifo_real : entity xil_defaultlib.pilotdetect_xlfifogen_u
  generic map (
    core_name0 => "pilotdetect_fifo_generator_v13_1_i0",
    data_count_width => 9,
    data_width => 18,
    extra_registers => 1,
    has_ae => 0,
    has_af => 0,
    has_rst => false,
    percent_full_width => 1
  )
  port map (
    en => '1',
    rst => '1',
    din => delay0_q_net_x0,
    we => delay1_q_net_x0(0),
    re => new_correlator_ctrl_pop_net(0),
    clk => clk_net,
    ce => ce_net,
    we_ce => ce_net,
    re_ce => ce_net,
    dout => fifo_real_dout_net,
    empty => fifo_real_empty_net,
    percent_full => fifo_real_percent_full_net,
    full => fifo_real_full_net
  );
  mux : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => new_correlator_ctrl_write_zeros_net,
    d0 => fifo_real_dout_net,
    d1 => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => new_correlator_ctrl_write_zeros_net,
    d0 => fifo_imag_dout_net,
    d1 => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux2_y_net
  );
  relational : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant1_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  new_correlator_ctrl : entity xil_defaultlib.sysgen_mcode_block_fcf00fc5a8
  port map (
    clr => '0',
    fifo_full(0) => fifo_real_full_net,
    cnt_eq_512 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    pop => new_correlator_ctrl_pop_net,
    start_correlator => new_correlator_ctrl_start_correlator_net,
    count_rst => new_correlator_ctrl_count_rst_net,
    write_zeros => new_correlator_ctrl_write_zeros_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/complex_mult
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult;
architecture structural of pilotdetect_complex_mult is
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay4_q_net_x0 <= b_r;
  delay5_q_net_x0 <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/complex_mult2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult2 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult2;
architecture structural of pilotdetect_complex_mult2 is
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay22_q_net <= b_r;
  delay23_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/complex_mult3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult3 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult3;
architecture structural of pilotdetect_complex_mult3 is
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay19_q_net <= b_r;
  delay21_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/complex_mult4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult4 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult4;
architecture structural of pilotdetect_complex_mult4 is
  signal delay18_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay29_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay18_q_net <= b_r;
  delay29_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay18_q_net,
    b => delay29_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay18_q_net,
    b => delay29_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_complex_delay6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay6 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay6;
architecture structural of pilotdetect_large_complex_delay6 is
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal clk_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i0",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i1",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_complex_delay7
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay7 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay7;
architecture structural of pilotdetect_large_complex_delay7 is
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 8-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 8,
    c_address_width_b => 8,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i1",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i2",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_complex_delay8
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay8 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay8;
architecture structural of pilotdetect_large_complex_delay8 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 7-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 7-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i2",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_complex_delay9
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay9 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay9;
architecture structural of pilotdetect_large_complex_delay9 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 6-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 6-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 6,
    c_address_width_b => 6,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i3",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i7",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_tfactor_rom1/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x0 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 10-1 downto 0 )
  );
end pilotdetect_address_generator_x0;
architecture structural of pilotdetect_address_generator_x0 is
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 10-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 10-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 10-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant_op_net : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 10-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 10,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 10,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 11,
    core_name0 => "pilotdetect_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 11,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 10
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b834ce322d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_65e9092d81
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_f84e73127e
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_377354b5ea
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mux : entity xil_defaultlib.sysgen_mux_81939abd89
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 9,
    x_width => 10,
    y_width => 10
  )
  port map (
    x => counter_op_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_tfactor_rom1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_tfactor_rom1 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_tfactor_rom1;
architecture structural of pilotdetect_large_tfactor_rom1 is
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 9-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 10-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x0
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_222d6d85fc
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 10
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i4",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_tfactor_rom2/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x1 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 8-1 downto 0 )
  );
end pilotdetect_address_generator_x1;
architecture structural of pilotdetect_address_generator_x1 is
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 8-1 downto 0 );
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 8-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 8-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 6-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant_op_net : std_logic_vector( 8-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 8,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 8,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 9,
    core_name0 => "pilotdetect_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 9,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 8
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_2b7c6b2428
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_a8c933a1a7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_b4de442209
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_78f34e96e5
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mux : entity xil_defaultlib.sysgen_mux_4b3c2484ae
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => counter_op_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/large_tfactor_rom2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_tfactor_rom2 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_tfactor_rom2;
architecture structural of pilotdetect_large_tfactor_rom2 is
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 8-1 downto 0 );
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal slice_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 8-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 7-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x1
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_2e499fd69d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i5",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2I2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2i2 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2i2;
architecture structural of pilotdetect_nbr_bf2i2 is
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal shift4_op_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  shift1_op_net <= x_r;
  shift4_op_net <= x_i;
  delay0_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => shift1_op_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => shift1_op_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => shift4_op_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => shift4_op_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay0_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => shift1_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => shift4_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 513,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 9,
    new_msb => 9,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2I3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2i3 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2i3;
architecture structural of pilotdetect_nbr_bf2i3 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net_x0;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 129,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 7,
    new_msb => 7,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2I4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2i4 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2i4;
architecture structural of pilotdetect_nbr_bf2i4 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay25_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay26_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay26_q_net <= delta_x_r;
  delay25_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay24_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay26_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay26_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay25_q_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay25_q_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay26_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay25_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 33,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 5,
    new_msb => 5,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2I5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2i5 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2i5;
architecture structural of pilotdetect_nbr_bf2i5 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay2_q_net <= delta_x_r;
  delay1_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay28_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net_x0
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 9,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net_x0,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net_x0,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 3,
    new_msb => 3,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2I6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2i6 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2i6;
architecture structural of pilotdetect_nbr_bf2i6 is
  signal delay30_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay8_q_net <= delta_x_r;
  delay9_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay30_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay30_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay9_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay30_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 1,
    new_msb => 1,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2II2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2ii2 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2ii2;
architecture structural of pilotdetect_nbr_bf2ii2 is
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift7_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift6_op_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net_x0;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  shift6_op_net <= x_r;
  shift7_op_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 258,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift6_op_net,
    d1 => shift7_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift7_op_net,
    d1 => shift6_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 8,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 9,
    new_msb => 9,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2II3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2ii3 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2ii3;
architecture structural of pilotdetect_nbr_bf2ii3 is
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift10_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift11_op_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net_x0;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  shift10_op_net <= x_r;
  shift11_op_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 66,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift10_op_net,
    d1 => shift11_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift11_op_net,
    d1 => shift10_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 6,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 7,
    new_msb => 7,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2II4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2ii4 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2ii4;
architecture structural of pilotdetect_nbr_bf2ii4 is
  signal delay27_q_net : std_logic_vector( 18-1 downto 0 );
  signal shift15_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay20_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal shift14_op_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net_x0;
  delay20_q_net <= delta_x_r;
  delay27_q_net <= delta_x_i;
  shift14_op_net <= x_r;
  shift15_op_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay20_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay20_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay27_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay27_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay20_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay27_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 18,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift14_op_net,
    d1 => shift15_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift15_op_net,
    d1 => shift14_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 4,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 5,
    new_msb => 5,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2II5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2ii5 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2ii5;
architecture structural of pilotdetect_nbr_bf2ii5 is
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift18_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal shift19_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net_x0;
  delay3_q_net <= delta_x_r;
  delay7_q_net <= delta_x_i;
  shift18_op_net <= x_r;
  shift19_op_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net_x0
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 6,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net_x0
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net_x0,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net_x0,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift18_op_net,
    d1 => shift19_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift19_op_net,
    d1 => shift18_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 2,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 3,
    new_msb => 3,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/nbr_BF2II6
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_nbr_bf2ii6 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_nbr_bf2ii6;
architecture structural of pilotdetect_nbr_bf2ii6 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift5_op_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay10_q_net <= delta_x_r;
  delay11_q_net <= delta_x_i;
  shift_op_net <= x_r;
  shift5_op_net <= x_i;
  delay12_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay12_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay10_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift_op_net,
    d1 => shift5_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift5_op_net,
    d1 => shift_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 1,
    new_msb => 1,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/small_tfactor_rom/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x2 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 6-1 downto 0 )
  );
end pilotdetect_address_generator_x2;
architecture structural of pilotdetect_address_generator_x2 is
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 6-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 6-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 6-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 6-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 6-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 6-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 6,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 6,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 7,
    core_name0 => "pilotdetect_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 7,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 6
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_392cf7ce5c
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_4adcefda0f
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_a152b8b4ce
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7d4cdb5bbb
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bba3bd89f4
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 10,
    y_width => 6
  )
  port map (
    x => counter_op_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/small_tfactor_rom
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_small_tfactor_rom is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_small_tfactor_rom;
architecture structural of pilotdetect_small_tfactor_rom is
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 6-1 downto 0 );
  signal slice_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal delay_q_net : std_logic_vector( 6-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 5-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x2
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_c024ed0ea3
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 6
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram_dist
  generic map (
    addr_width => 5,
    c_address_width => 5,
    c_width => 18,
    core_name0 => "pilotdetect_dist_mem_gen_v8_0_i0",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/small_tfactor_rom1/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x3 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 4-1 downto 0 )
  );
end pilotdetect_address_generator_x3;
architecture structural of pilotdetect_address_generator_x3 is
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant_op_net : std_logic_vector( 4-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 4-1 downto 0 );
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 4-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 4-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 2-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 4-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 4,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 4,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 5,
    core_name0 => "pilotdetect_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 5,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 4
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_6a9e537061
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_55eaac7d5b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bb4a1d2355
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 10,
    y_width => 4
  )
  port map (
    x => counter_op_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024/small_tfactor_rom1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_small_tfactor_rom1 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_small_tfactor_rom1;
architecture structural of pilotdetect_small_tfactor_rom1 is
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 4-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 3-1 downto 0 );
  signal ce_net : std_logic;
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 4-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x3
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_1672b64d97
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 4
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram_dist
  generic map (
    addr_width => 3,
    c_address_width => 4,
    c_width => 18,
    core_name0 => "pilotdetect_dist_mem_gen_v8_0_i1",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_1024
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_fft_1024 is
  port (
    x_r_x0 : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i_x0 : out std_logic_vector( 18-1 downto 0 );
    done : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_fft_1024;
architecture structural of pilotdetect_fft_1024 is
  signal mux1_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay29_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x9 : std_logic_vector( 1-1 downto 0 );
  signal shift4_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x13 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal delay26_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal delay25_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret3_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay20_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal shift11_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal shift10_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal shift7_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal shift15_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal shift18_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal shift5_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal shift6_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift14_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay30_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay27_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal shift19_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift17_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift13_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift12_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift20_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift16_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift8_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift9_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift21_op_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= mux_y_net_x2;
  x_i_x0 <= mux1_y_net_x1;
  done <= delay6_q_net_x0;
  mux_y_net <= x_r_x0;
  mux2_y_net <= x_i;
  delay0_q_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  complex_mult : entity xil_defaultlib.pilotdetect_complex_mult
  port map (
    a_r => mux_y_net_x13,
    a_i => mux1_y_net_x12,
    b_r => delay4_q_net_x3,
    b_i => delay5_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2
  );
  complex_mult2 : entity xil_defaultlib.pilotdetect_complex_mult2
  port map (
    a_r => mux_y_net_x12,
    a_i => mux1_y_net_x11,
    b_r => delay22_q_net,
    b_i => delay23_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1
  );
  complex_mult3 : entity xil_defaultlib.pilotdetect_complex_mult3
  port map (
    a_r => mux_y_net_x1,
    a_i => mux1_y_net_x0,
    b_r => delay19_q_net,
    b_i => delay21_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0
  );
  complex_mult4 : entity xil_defaultlib.pilotdetect_complex_mult4
  port map (
    a_r => mux_y_net_x0,
    a_i => mux1_y_net,
    b_r => delay18_q_net,
    b_i => delay29_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net,
    x_i => delay5_q_net
  );
  large_complex_delay6 : entity xil_defaultlib.pilotdetect_large_complex_delay6
  port map (
    in_r => mux3_y_net_x8,
    in_i => mux2_y_net_x9,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net,
    out_i => reinterpret3_output_port_net_x2
  );
  large_complex_delay7 : entity xil_defaultlib.pilotdetect_large_complex_delay7
  port map (
    in_r => mux3_y_net_x3,
    in_i => mux2_y_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x2,
    out_i => reinterpret3_output_port_net_x1
  );
  large_complex_delay8 : entity xil_defaultlib.pilotdetect_large_complex_delay8
  port map (
    in_r => mux3_y_net_x7,
    in_i => mux2_y_net_x8,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x1,
    out_i => reinterpret3_output_port_net_x0
  );
  large_complex_delay9 : entity xil_defaultlib.pilotdetect_large_complex_delay9
  port map (
    in_r => mux3_y_net_x2,
    in_i => mux2_y_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x0,
    out_i => reinterpret3_output_port_net
  );
  large_tfactor_rom1 : entity xil_defaultlib.pilotdetect_large_tfactor_rom1
  port map (
    in1 => delay6_q_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x13,
    w_i => mux1_y_net_x12
  );
  large_tfactor_rom2 : entity xil_defaultlib.pilotdetect_large_tfactor_rom2
  port map (
    in1 => delay6_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x12,
    w_i => mux1_y_net_x11
  );
  nbr_bf2i2 : entity xil_defaultlib.pilotdetect_nbr_bf2i2
  port map (
    delta_x_r => reinterpret3_output_port_net_x2,
    delta_x_i => reinterpret2_output_port_net,
    x_r => shift1_op_net,
    x_i => shift4_op_net,
    start_in => delay0_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x9,
    delta_y_i => mux3_y_net_x8,
    y_r => mux_y_net_x11,
    y_i => mux1_y_net_x10,
    start_out => delay6_q_net_x9
  );
  nbr_bf2i3 : entity xil_defaultlib.pilotdetect_nbr_bf2i3
  port map (
    delta_x_r => reinterpret3_output_port_net_x0,
    delta_x_i => reinterpret2_output_port_net_x1,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2,
    start_in => delay6_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x8,
    delta_y_i => mux3_y_net_x7,
    y_r => mux_y_net_x10,
    y_i => mux1_y_net_x9,
    start_out => delay6_q_net_x8
  );
  nbr_bf2i4 : entity xil_defaultlib.pilotdetect_nbr_bf2i4
  port map (
    delta_x_r => delay26_q_net,
    delta_x_i => delay25_q_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1,
    start_in => delay24_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x7,
    delta_y_i => mux3_y_net_x6,
    y_r => mux_y_net_x9,
    y_i => mux1_y_net_x8,
    start_out => delay6_q_net_x7
  );
  nbr_bf2i5 : entity xil_defaultlib.pilotdetect_nbr_bf2i5
  port map (
    delta_x_r => delay2_q_net,
    delta_x_i => delay1_q_net,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0,
    start_in => delay28_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x6,
    delta_y_i => mux3_y_net_x5,
    y_r => mux_y_net_x8,
    y_i => mux1_y_net_x7,
    start_out => delay6_q_net_x6
  );
  nbr_bf2i6 : entity xil_defaultlib.pilotdetect_nbr_bf2i6
  port map (
    delta_x_r => delay8_q_net,
    delta_x_i => delay9_q_net,
    x_r => delay4_q_net,
    x_i => delay5_q_net,
    start_in => delay30_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x5,
    delta_y_i => mux3_y_net_x4,
    y_r => mux_y_net_x7,
    y_i => mux1_y_net_x6,
    start_out => delay6_q_net_x5
  );
  nbr_bf2ii2 : entity xil_defaultlib.pilotdetect_nbr_bf2ii2
  port map (
    delta_x_r => reinterpret3_output_port_net_x1,
    delta_x_i => reinterpret2_output_port_net_x2,
    x_r => shift6_op_net,
    x_i => shift7_op_net,
    start_in => delay6_q_net_x9,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x4,
    delta_y_i => mux3_y_net_x3,
    y_r => mux_y_net_x6,
    y_i => mux1_y_net_x5,
    start_out => delay6_q_net_x4
  );
  nbr_bf2ii3 : entity xil_defaultlib.pilotdetect_nbr_bf2ii3
  port map (
    delta_x_r => reinterpret3_output_port_net,
    delta_x_i => reinterpret2_output_port_net_x0,
    x_r => shift10_op_net,
    x_i => shift11_op_net,
    start_in => delay6_q_net_x8,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x3,
    delta_y_i => mux3_y_net_x2,
    y_r => mux_y_net_x5,
    y_i => mux1_y_net_x4,
    start_out => delay6_q_net_x3
  );
  nbr_bf2ii4 : entity xil_defaultlib.pilotdetect_nbr_bf2ii4
  port map (
    delta_x_r => delay20_q_net,
    delta_x_i => delay27_q_net,
    x_r => shift14_op_net,
    x_i => shift15_op_net,
    start_in => delay6_q_net_x7,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x2,
    delta_y_i => mux3_y_net,
    y_r => mux_y_net_x4,
    y_i => mux1_y_net_x3,
    start_out => delay6_q_net_x2
  );
  nbr_bf2ii5 : entity xil_defaultlib.pilotdetect_nbr_bf2ii5
  port map (
    delta_x_r => delay3_q_net,
    delta_x_i => delay7_q_net,
    x_r => shift18_op_net,
    x_i => shift19_op_net,
    start_in => delay6_q_net_x6,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x1,
    delta_y_i => mux3_y_net_x1,
    y_r => mux_y_net_x3,
    y_i => mux1_y_net_x2,
    start_out => delay6_q_net_x1
  );
  nbr_bf2ii6 : entity xil_defaultlib.pilotdetect_nbr_bf2ii6
  port map (
    delta_x_r => delay10_q_net,
    delta_x_i => delay11_q_net,
    x_r => shift_op_net,
    x_i => shift5_op_net,
    start_in => delay12_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x0,
    delta_y_i => mux3_y_net_x0,
    y_r => mux_y_net_x2,
    y_i => mux1_y_net_x1,
    start_out => delay6_q_net_x0
  );
  small_tfactor_rom : entity xil_defaultlib.pilotdetect_small_tfactor_rom
  port map (
    in1 => delay6_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x1,
    w_i => mux1_y_net_x0
  );
  small_tfactor_rom1 : entity xil_defaultlib.pilotdetect_small_tfactor_rom1
  port map (
    in1 => delay6_q_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x0,
    w_i => mux1_y_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux2_y_net_x0,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux3_y_net_x0,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay12_q_net
  );
  delay18 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift20_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay18_q_net
  );
  delay19 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift16_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay19_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay20 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay20_q_net
  );
  delay21 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift17_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay21_q_net
  );
  delay22 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift12_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay22_q_net
  );
  delay23 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift13_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay23_q_net
  );
  delay24 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay24_q_net
  );
  delay25 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    q => delay25_q_net
  );
  delay26 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay26_q_net
  );
  delay27 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay27_q_net
  );
  delay28 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay28_q_net
  );
  delay29 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift21_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay29_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay30 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay30_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift8_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x3
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => shift9_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x3
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  shift : entity xil_defaultlib.sysgen_shift_c51054fc18
  port map (
    clr => '0',
    ip => mux_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    op => shift_op_net
  );
  shift1 : entity xil_defaultlib.sysgen_shift_c0cd8b3c82
  port map (
    clr => '0',
    ip => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    op => shift1_op_net
  );
  shift10 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x10,
    clk => clk_net,
    ce => ce_net,
    op => shift10_op_net
  );
  shift11 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x9,
    clk => clk_net,
    ce => ce_net,
    op => shift11_op_net
  );
  shift12 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    op => shift12_op_net
  );
  shift13 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    op => shift13_op_net
  );
  shift14 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x9,
    clk => clk_net,
    ce => ce_net,
    op => shift14_op_net
  );
  shift15 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    op => shift15_op_net
  );
  shift16 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    op => shift16_op_net
  );
  shift17 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    op => shift17_op_net
  );
  shift18 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    op => shift18_op_net
  );
  shift19 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    op => shift19_op_net
  );
  shift20 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    op => shift20_op_net
  );
  shift21 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    op => shift21_op_net
  );
  shift4 : entity xil_defaultlib.sysgen_shift_c0cd8b3c82
  port map (
    clr => '0',
    ip => mux2_y_net,
    clk => clk_net,
    ce => ce_net,
    op => shift4_op_net
  );
  shift5 : entity xil_defaultlib.sysgen_shift_c51054fc18
  port map (
    clr => '0',
    ip => mux1_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    op => shift5_op_net
  );
  shift6 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x11,
    clk => clk_net,
    ce => ce_net,
    op => shift6_op_net
  );
  shift7 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x10,
    clk => clk_net,
    ce => ce_net,
    op => shift7_op_net
  );
  shift8 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux_y_net_x6,
    clk => clk_net,
    ce => ce_net,
    op => shift8_op_net
  );
  shift9 : entity xil_defaultlib.sysgen_shift_dc7d2f1ef0
  port map (
    clr => '0',
    ip => mux1_y_net_x5,
    clk => clk_net,
    ce => ce_net,
    op => shift9_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/FFT_buf_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_fft_buf_control is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    write : out std_logic_vector( 1-1 downto 0 );
    write_addr : out std_logic_vector( 10-1 downto 0 )
  );
end pilotdetect_fft_buf_control;
architecture structural of pilotdetect_fft_buf_control is
  signal write_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal addr_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 10-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
begin
  write <= write_reg_q_net;
  write_addr <= addr_op_net;
  delay6_q_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant_x0 : entity xil_defaultlib.sysgen_constant_1993043fd7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  expression : entity xil_defaultlib.sysgen_expr_ecdb93f3d8
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    addr_eq_1023 => relational_op_net,
    start => delay6_q_net,
    wait_x0 => wait_reg_q_net,
    write => write_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_d590143351
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    addr_eq_1023 => relational_op_net,
    start => delay6_q_net,
    wait_x0 => wait_reg_q_net,
    write => write_reg_q_net,
    dout => expression1_dout_net
  );
  relational : entity xil_defaultlib.sysgen_relational_a77d10299f
  port map (
    clr => '0',
    a => addr_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
  write_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => write_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2I
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i;
architecture structural of pilotdetect_bf2i is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay17_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay1_q_net_x0 <= delta_x_r;
  delay_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net_x0 <= x_i;
  delay17_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net_x0,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net_x0,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay1_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 2,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2I1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i1;
architecture structural of pilotdetect_bf2i1 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay8_q_net <= delta_x_r;
  delay7_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net_x0 <= x_i;
  delay6_q_net_x0 <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 17,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 4,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2I2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i2 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i2;
architecture structural of pilotdetect_bf2i2 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay12_q_net <= delta_x_r;
  delay11_q_net <= delta_x_i;
  delay5_q_net_x0 <= x_r;
  delay4_q_net_x0 <= x_i;
  delay2_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay12_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay12_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net_x0,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2I3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i3 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i3;
architecture structural of pilotdetect_bf2i3 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay24_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 65,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 6,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2I4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i4 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i4;
architecture structural of pilotdetect_bf2i4 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay28_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 257,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 8,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2II
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii;
architecture structural of pilotdetect_bf2ii is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay3_q_net_x0 <= delta_x_r;
  delay2_q_net_x0 <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net_x0,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net_x0,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net_x0,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net_x0,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay3_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay2_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 10,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 3,
    new_msb => 3,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 2,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2II1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii1;
architecture structural of pilotdetect_bf2ii1 is
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay10_q_net <= delta_x_r;
  delay9_q_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay10_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay9_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 34,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 5,
    new_msb => 5,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 4,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2II2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii2 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii2;
architecture structural of pilotdetect_bf2ii2 is
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay14_q_net <= delta_x_r;
  delay13_q_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay14_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay14_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay13_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay13_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 1,
    new_msb => 1,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2II3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii3 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii3;
architecture structural of pilotdetect_bf2ii3 is
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 130,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 7,
    new_msb => 7,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 6,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/BF2II4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii4 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_bf2ii4;
architecture structural of pilotdetect_bf2ii4 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  shift_op_net <= x_r;
  shift1_op_net <= x_i;
  delay18_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay18_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift_op_net,
    d1 => shift1_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift1_op_net,
    d1 => shift_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 9,
    new_msb => 9,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 8,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/complex_mult
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult_x0 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult_x0;
architecture structural of pilotdetect_complex_mult_x0 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay4_q_net_x0 <= b_r;
  delay5_q_net_x0 <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/complex_mult1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult1_x0 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult1_x0;
architecture structural of pilotdetect_complex_mult1_x0 is
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay16_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay15_q_net <= b_r;
  delay16_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay15_q_net,
    b => delay16_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay15_q_net,
    b => delay16_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/complex_mult2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult2_x1 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult2_x1;
architecture structural of pilotdetect_complex_mult2_x1 is
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay22_q_net <= b_r;
  delay23_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/complex_mult3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult3_x1 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult3_x1;
architecture structural of pilotdetect_complex_mult3_x1 is
  signal clk_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay19_q_net <= b_r;
  delay21_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_complex_delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay;
architecture structural of pilotdetect_large_complex_delay is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 9-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i0",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i1",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_complex_delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay1 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay1;
architecture structural of pilotdetect_large_complex_delay1 is
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 8-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 8,
    c_address_width_b => 8,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i1",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i2",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_complex_delay4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay4 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay4;
architecture structural of pilotdetect_large_complex_delay4 is
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal ce_net : std_logic;
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 7-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 7-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i2",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_complex_delay5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay5 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay5;
architecture structural of pilotdetect_large_complex_delay5 is
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 6-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 6-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 6,
    c_address_width_b => 6,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i3",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i7",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_inv_tfactor_rom/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x4 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 10-1 downto 0 )
  );
end pilotdetect_address_generator_x4;
architecture structural of pilotdetect_address_generator_x4 is
  signal addsub_s_net : std_logic_vector( 10-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 10-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 10-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 10-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 8-1 downto 0 );
  signal clk_net : std_logic;
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 10-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 10,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 10,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 11,
    core_name0 => "pilotdetect_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 11,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 10
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b834ce322d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_65e9092d81
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_f84e73127e
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_377354b5ea
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_81939abd89
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 9,
    x_width => 10,
    y_width => 10
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_inv_tfactor_rom
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom;
architecture structural of pilotdetect_large_inv_tfactor_rom is
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 10-1 downto 0 );
  signal clk_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal slice_y_net : std_logic_vector( 8-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay_q_net : std_logic_vector( 10-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x4
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_222d6d85fc
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 10
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i4",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_inv_tfactor_rom1/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x5 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 8-1 downto 0 )
  );
end pilotdetect_address_generator_x5;
architecture structural of pilotdetect_address_generator_x5 is
  signal mux_y_net : std_logic_vector( 8-1 downto 0 );
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 8-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 6-1 downto 0 );
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 8-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant_op_net : std_logic_vector( 8-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 8,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 8,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 9,
    core_name0 => "pilotdetect_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 9,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 8
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_2b7c6b2428
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_a8c933a1a7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_b4de442209
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_78f34e96e5
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_4b3c2484ae
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_inv_tfactor_rom1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom1 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom1;
architecture structural of pilotdetect_large_inv_tfactor_rom1 is
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice_y_net : std_logic_vector( 6-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 8-1 downto 0 );
  signal delay_q_net : std_logic_vector( 8-1 downto 0 );
  signal clk_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 7-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x5
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_2e499fd69d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i5",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_inv_tfactor_rom2/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x6 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 6-1 downto 0 )
  );
end pilotdetect_address_generator_x6;
architecture structural of pilotdetect_address_generator_x6 is
  signal clk_net : std_logic;
  signal addsub_s_net : std_logic_vector( 6-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 6-1 downto 0 );
  signal mux_y_net : std_logic_vector( 6-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal constant_op_net : std_logic_vector( 6-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 6-1 downto 0 );
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 6-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 6,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 6,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 7,
    core_name0 => "pilotdetect_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 7,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 6
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_392cf7ce5c
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_4adcefda0f
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_a152b8b4ce
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7d4cdb5bbb
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bba3bd89f4
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 10,
    y_width => 6
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/large_inv_tfactor_rom2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom2 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom2;
architecture structural of pilotdetect_large_inv_tfactor_rom2 is
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 6-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 6-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 5-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 4-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x6
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_c024ed0ea3
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 6
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 5,
    c_address_width_b => 5,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i6",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/small_inv_tfactor_rom4/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x7 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 4-1 downto 0 )
  );
end pilotdetect_address_generator_x7;
architecture structural of pilotdetect_address_generator_x7 is
  signal mux_y_net : std_logic_vector( 4-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 4-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 4-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 4-1 downto 0 );
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 2-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant_op_net : std_logic_vector( 4-1 downto 0 );
  signal ce_net : std_logic;
  signal concat1_y_net : std_logic_vector( 4-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 4-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 4,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 4,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 5,
    core_name0 => "pilotdetect_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 5,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 4
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_6a9e537061
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_55eaac7d5b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bb4a1d2355
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 10,
    y_width => 4
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1/small_inv_tfactor_rom4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_small_inv_tfactor_rom4 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_small_inv_tfactor_rom4;
architecture structural of pilotdetect_small_inv_tfactor_rom4 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 4-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 3-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 4-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x7
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_1672b64d97
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 4
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram_dist
  generic map (
    addr_width => 3,
    c_address_width => 4,
    c_width => 18,
    core_name0 => "pilotdetect_dist_mem_gen_v8_0_i1",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_ifft_1024_ver_1 is
  port (
    x_r_x0 : in std_logic_vector( 18-1 downto 0 );
    x_i_x0 : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_ifft_1024_ver_1;
architecture structural of pilotdetect_ifft_1024_ver_1 is
  signal mux1_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay17_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux1_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x9 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x1 : std_logic_vector( 1-1 downto 0 );
begin
  x_r <= mux1_y_net;
  x_i <= mux_y_net;
  delay4_q_net <= x_r_x0;
  delay5_q_net <= x_i_x0;
  delay2_q_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  bf2i : entity xil_defaultlib.pilotdetect_bf2i
  port map (
    delta_x_r => delay1_q_net,
    delta_x_i => delay_q_net,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2,
    start_in => delay17_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x8,
    delta_y_i => mux3_y_net_x8,
    y_r => mux_y_net_x7,
    y_i => mux1_y_net_x8,
    start_out => delay6_q_net_x8
  );
  bf2i1 : entity xil_defaultlib.pilotdetect_bf2i1
  port map (
    delta_x_r => delay8_q_net,
    delta_x_i => delay7_q_net,
    x_r => delay4_q_net_x3,
    x_i => delay5_q_net_x3,
    start_in => delay6_q_net_x9,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x7,
    delta_y_i => mux3_y_net_x7,
    y_r => mux_y_net_x6,
    y_i => mux1_y_net_x7,
    start_out => delay6_q_net_x7
  );
  bf2i2 : entity xil_defaultlib.pilotdetect_bf2i2
  port map (
    delta_x_r => delay12_q_net,
    delta_x_i => delay11_q_net,
    x_r => delay5_q_net,
    x_i => delay4_q_net,
    start_in => delay2_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x6,
    delta_y_i => mux3_y_net_x6,
    y_r => mux_y_net_x5,
    y_i => mux1_y_net_x6,
    start_out => delay6_q_net_x6
  );
  bf2i3 : entity xil_defaultlib.pilotdetect_bf2i3
  port map (
    delta_x_r => reinterpret3_output_port_net,
    delta_x_i => reinterpret2_output_port_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1,
    start_in => delay24_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x5,
    delta_y_i => mux3_y_net_x5,
    y_r => mux_y_net_x4,
    y_i => mux1_y_net_x5,
    start_out => delay6_q_net_x5
  );
  bf2i4 : entity xil_defaultlib.pilotdetect_bf2i4
  port map (
    delta_x_r => reinterpret3_output_port_net_x1,
    delta_x_i => reinterpret2_output_port_net_x1,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0,
    start_in => delay28_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x4,
    delta_y_i => mux3_y_net_x4,
    y_r => mux_y_net_x3,
    y_i => mux1_y_net_x4,
    start_out => delay6_q_net_x4
  );
  bf2ii : entity xil_defaultlib.pilotdetect_bf2ii
  port map (
    delta_x_r => delay3_q_net,
    delta_x_i => delay2_q_net_x0,
    x_r => mux_y_net_x7,
    x_i => mux1_y_net_x8,
    start_in => delay6_q_net_x8,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x3,
    delta_y_i => mux3_y_net_x3,
    y_r => mux_y_net_x2,
    y_i => mux1_y_net_x3,
    start_out => delay6_q_net_x3
  );
  bf2ii1 : entity xil_defaultlib.pilotdetect_bf2ii1
  port map (
    delta_x_r => delay10_q_net,
    delta_x_i => delay9_q_net,
    x_r => mux_y_net_x6,
    x_i => mux1_y_net_x7,
    start_in => delay6_q_net_x7,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x2,
    delta_y_i => mux3_y_net_x2,
    y_r => mux_y_net_x12,
    y_i => mux1_y_net_x2,
    start_out => delay6_q_net_x2
  );
  bf2ii2 : entity xil_defaultlib.pilotdetect_bf2ii2
  port map (
    delta_x_r => delay14_q_net,
    delta_x_i => delay13_q_net,
    x_r => mux_y_net_x5,
    x_i => mux1_y_net_x6,
    start_in => delay6_q_net_x6,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x1,
    delta_y_i => mux3_y_net_x1,
    y_r => mux_y_net_x1,
    y_i => mux1_y_net_x1,
    start_out => delay6_q_net_x1
  );
  bf2ii3 : entity xil_defaultlib.pilotdetect_bf2ii3
  port map (
    delta_x_r => reinterpret3_output_port_net_x0,
    delta_x_i => reinterpret2_output_port_net_x0,
    x_r => mux_y_net_x4,
    x_i => mux1_y_net_x5,
    start_in => delay6_q_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x0,
    delta_y_i => mux3_y_net_x0,
    y_r => mux_y_net_x0,
    y_i => mux1_y_net_x0,
    start_out => delay6_q_net_x0
  );
  bf2ii4 : entity xil_defaultlib.pilotdetect_bf2ii4
  port map (
    delta_x_r => reinterpret3_output_port_net_x2,
    delta_x_i => reinterpret2_output_port_net_x2,
    x_r => shift_op_net,
    x_i => shift1_op_net,
    start_in => delay18_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net,
    delta_y_i => mux3_y_net,
    y_r => mux_y_net,
    y_i => mux1_y_net
  );
  complex_mult : entity xil_defaultlib.pilotdetect_complex_mult_x0
  port map (
    a_r => mux_y_net_x10,
    a_i => mux1_y_net_x11,
    b_r => delay4_q_net_x4,
    b_i => delay5_q_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x3,
    x_i => delay5_q_net_x3
  );
  complex_mult1 : entity xil_defaultlib.pilotdetect_complex_mult1_x0
  port map (
    a_r => mux_y_net_x11,
    a_i => mux1_y_net_x12,
    b_r => delay15_q_net,
    b_i => delay16_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2
  );
  complex_mult2 : entity xil_defaultlib.pilotdetect_complex_mult2_x1
  port map (
    a_r => mux_y_net_x9,
    a_i => mux1_y_net_x10,
    b_r => delay22_q_net,
    b_i => delay23_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1
  );
  complex_mult3 : entity xil_defaultlib.pilotdetect_complex_mult3_x1
  port map (
    a_r => mux_y_net_x8,
    a_i => mux1_y_net_x9,
    b_r => delay19_q_net,
    b_i => delay21_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0
  );
  large_complex_delay : entity xil_defaultlib.pilotdetect_large_complex_delay
  port map (
    in_r => mux3_y_net,
    in_i => mux2_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x2,
    out_i => reinterpret3_output_port_net_x2
  );
  large_complex_delay1 : entity xil_defaultlib.pilotdetect_large_complex_delay1
  port map (
    in_r => mux3_y_net_x4,
    in_i => mux2_y_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x1,
    out_i => reinterpret3_output_port_net_x1
  );
  large_complex_delay4 : entity xil_defaultlib.pilotdetect_large_complex_delay4
  port map (
    in_r => mux3_y_net_x0,
    in_i => mux2_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x0,
    out_i => reinterpret3_output_port_net_x0
  );
  large_complex_delay5 : entity xil_defaultlib.pilotdetect_large_complex_delay5
  port map (
    in_r => mux3_y_net_x5,
    in_i => mux2_y_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net,
    out_i => reinterpret3_output_port_net
  );
  large_inv_tfactor_rom : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom
  port map (
    in1 => delay6_q_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x11,
    w_i => mux1_y_net_x12
  );
  large_inv_tfactor_rom1 : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom1
  port map (
    in1 => delay6_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x10,
    w_i => mux1_y_net_x11
  );
  large_inv_tfactor_rom2 : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom2
  port map (
    in1 => delay6_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x9,
    w_i => mux1_y_net_x10
  );
  small_inv_tfactor_rom4 : entity xil_defaultlib.pilotdetect_small_inv_tfactor_rom4
  port map (
    in1 => delay6_q_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x8,
    w_i => mux1_y_net_x9
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux3_y_net_x6,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux2_y_net_x6,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
  delay16 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  delay17 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay17_q_net
  );
  delay18 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay18_q_net
  );
  delay19 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay19_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay21 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay21_q_net
  );
  delay22 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x12,
    clk => clk_net,
    ce => ce_net,
    q => delay22_q_net
  );
  delay23 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay23_q_net
  );
  delay24 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay24_q_net
  );
  delay28 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay28_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x4
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x4
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x9
  );
  delay7 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  shift : entity xil_defaultlib.sysgen_shift_5fce716372
  port map (
    clr => '0',
    ip => mux_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    op => shift_op_net
  );
  shift1 : entity xil_defaultlib.sysgen_shift_5fce716372
  port map (
    clr => '0',
    ip => mux1_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    op => shift1_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2I
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i_x0;
architecture structural of pilotdetect_bf2i_x0 is
  signal delay17_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay1_q_net_x0 <= delta_x_r;
  delay_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net_x0 <= x_i;
  delay17_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net_x0,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net_x0,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay1_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 2,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2I1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i1_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i1_x0;
architecture structural of pilotdetect_bf2i1_x0 is
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay8_q_net <= delta_x_r;
  delay7_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net_x0 <= x_i;
  delay6_q_net_x0 <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 17,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 4,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2I2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i2_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i2_x0;
architecture structural of pilotdetect_bf2i2_x0 is
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay12_q_net <= delta_x_r;
  delay11_q_net <= delta_x_i;
  delay5_q_net_x0 <= x_r;
  delay4_q_net_x0 <= x_i;
  delay2_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay12_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay12_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net_x0,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2I3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i3_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i3_x0;
architecture structural of pilotdetect_bf2i3_x0 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay24_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 65,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 6,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2I4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i4_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i4_x0;
architecture structural of pilotdetect_bf2i4_x0 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay28_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 257,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 8,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2II
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii_x0;
architecture structural of pilotdetect_bf2ii_x0 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay3_q_net_x0 <= delta_x_r;
  delay2_q_net_x0 <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net_x0,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net_x0,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net_x0,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net_x0,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay3_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay2_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 10,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 3,
    new_msb => 3,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 2,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2II1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii1_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii1_x0;
architecture structural of pilotdetect_bf2ii1_x0 is
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay10_q_net <= delta_x_r;
  delay9_q_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay10_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay9_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 34,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 5,
    new_msb => 5,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 4,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2II2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii2_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii2_x0;
architecture structural of pilotdetect_bf2ii2_x0 is
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay13_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay14_q_net <= delta_x_r;
  delay13_q_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay14_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay14_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay13_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay13_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 1,
    new_msb => 1,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2II3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii3_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii3_x0;
architecture structural of pilotdetect_bf2ii3_x0 is
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 130,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 7,
    new_msb => 7,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 6,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/BF2II4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii4_x0 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii4_x0;
architecture structural of pilotdetect_bf2ii4_x0 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  shift_op_net <= x_r;
  shift1_op_net <= x_i;
  delay18_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay18_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 514,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay18_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift_op_net,
    d1 => shift1_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift1_op_net,
    d1 => shift_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 9,
    new_msb => 9,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 8,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/complex_mult
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult_x1 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult_x1;
architecture structural of pilotdetect_complex_mult_x1 is
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay4_q_net_x0 <= b_r;
  delay5_q_net_x0 <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/complex_mult1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult1_x1 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult1_x1;
architecture structural of pilotdetect_complex_mult1_x1 is
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay15_q_net <= b_r;
  delay16_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay15_q_net,
    b => delay16_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay15_q_net,
    b => delay16_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/complex_mult2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult2_x2 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult2_x2;
architecture structural of pilotdetect_complex_mult2_x2 is
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay22_q_net <= b_r;
  delay23_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/complex_mult3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult3_x2 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult3_x2;
architecture structural of pilotdetect_complex_mult3_x2 is
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay19_q_net <= b_r;
  delay21_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_complex_delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay_x0 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay_x0;
architecture structural of pilotdetect_large_complex_delay_x0 is
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal ce_net : std_logic;
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 9-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 9-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i0",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i1",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_complex_delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay1_x0 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay1_x0;
architecture structural of pilotdetect_large_complex_delay1_x0 is
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 8-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 8,
    c_address_width_b => 8,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i1",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i2",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_complex_delay4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay4_x0 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay4_x0;
architecture structural of pilotdetect_large_complex_delay4_x0 is
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 7-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 7-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i2",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_complex_delay5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay5_x0 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay5_x0;
architecture structural of pilotdetect_large_complex_delay5_x0 is
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 6-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 6-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 6,
    c_address_width_b => 6,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i3",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i7",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_inv_tfactor_rom/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x8 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 10-1 downto 0 )
  );
end pilotdetect_address_generator_x8;
architecture structural of pilotdetect_address_generator_x8 is
  signal mux_y_net : std_logic_vector( 10-1 downto 0 );
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 10-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 10-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant_op_net : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 10-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 10,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 10,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 11,
    core_name0 => "pilotdetect_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 11,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 10
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b834ce322d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_65e9092d81
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_f84e73127e
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_377354b5ea
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_81939abd89
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 9,
    x_width => 10,
    y_width => 10
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_inv_tfactor_rom
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom_x0 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom_x0;
architecture structural of pilotdetect_large_inv_tfactor_rom_x0 is
  signal mux_y_net_x0 : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 8-1 downto 0 );
  signal clk_net : std_logic;
  signal concat1_y_net : std_logic_vector( 9-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 10-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x8
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_222d6d85fc
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 10
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i4",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_inv_tfactor_rom1/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x9 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 8-1 downto 0 )
  );
end pilotdetect_address_generator_x9;
architecture structural of pilotdetect_address_generator_x9 is
  signal ce_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 8-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 8-1 downto 0 );
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 8-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 8-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant_op_net : std_logic_vector( 8-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 8-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 8,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 8,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 9,
    core_name0 => "pilotdetect_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 9,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 8
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_2b7c6b2428
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_a8c933a1a7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_b4de442209
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_78f34e96e5
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_4b3c2484ae
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_inv_tfactor_rom1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom1_x0 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom1_x0;
architecture structural of pilotdetect_large_inv_tfactor_rom1_x0 is
  signal clk_net : std_logic;
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 6-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 8-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 7-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal delay_q_net : std_logic_vector( 8-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x9
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_2e499fd69d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i5",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_inv_tfactor_rom2/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x10 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 6-1 downto 0 )
  );
end pilotdetect_address_generator_x10;
architecture structural of pilotdetect_address_generator_x10 is
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 6-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal clk_net : std_logic;
  signal concat3_y_net : std_logic_vector( 6-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 6-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 4-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 6-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant_op_net : std_logic_vector( 6-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 6,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 6,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 7,
    core_name0 => "pilotdetect_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 7,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 6
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_392cf7ce5c
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_4adcefda0f
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_a152b8b4ce
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7d4cdb5bbb
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bba3bd89f4
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 10,
    y_width => 6
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/large_inv_tfactor_rom2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom2_x0 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom2_x0;
architecture structural of pilotdetect_large_inv_tfactor_rom2_x0 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 6-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 4-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 5-1 downto 0 );
  signal delay_q_net : std_logic_vector( 6-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x10
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_c024ed0ea3
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 6
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 5,
    c_address_width_b => 5,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i6",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/small_inv_tfactor_rom4/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x11 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 4-1 downto 0 )
  );
end pilotdetect_address_generator_x11;
architecture structural of pilotdetect_address_generator_x11 is
  signal mux_y_net : std_logic_vector( 4-1 downto 0 );
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 4-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 4-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 2-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant_op_net : std_logic_vector( 4-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 4-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 4,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 4,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 5,
    core_name0 => "pilotdetect_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 5,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 4
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_6a9e537061
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_55eaac7d5b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bb4a1d2355
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 10,
    y_width => 4
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2/small_inv_tfactor_rom4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_small_inv_tfactor_rom4_x0 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_small_inv_tfactor_rom4_x0;
architecture structural of pilotdetect_small_inv_tfactor_rom4_x0 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal concat1_y_net : std_logic_vector( 3-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay_q_net : std_logic_vector( 4-1 downto 0 );
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 4-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x11
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_1672b64d97
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 4
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram_dist
  generic map (
    addr_width => 3,
    c_address_width => 4,
    c_width => 18,
    core_name0 => "pilotdetect_dist_mem_gen_v8_0_i1",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_ifft_1024_ver_2 is
  port (
    x_r_x0 : in std_logic_vector( 18-1 downto 0 );
    x_i_x0 : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 );
    done : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_ifft_1024_ver_2;
architecture structural of pilotdetect_ifft_1024_ver_2 is
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal mux3_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay17_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x9 : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x12 : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= mux1_y_net;
  x_i <= mux_y_net;
  done <= delay6_q_net;
  delay4_q_net <= x_r_x0;
  delay5_q_net <= x_i_x0;
  delay2_q_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  bf2i : entity xil_defaultlib.pilotdetect_bf2i_x0
  port map (
    delta_x_r => delay1_q_net,
    delta_x_i => delay_q_net,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2,
    start_in => delay17_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x8,
    delta_y_i => mux3_y_net_x8,
    y_r => mux_y_net_x7,
    y_i => mux1_y_net_x8,
    start_out => delay6_q_net_x8
  );
  bf2i1 : entity xil_defaultlib.pilotdetect_bf2i1_x0
  port map (
    delta_x_r => delay8_q_net,
    delta_x_i => delay7_q_net,
    x_r => delay4_q_net_x3,
    x_i => delay5_q_net_x3,
    start_in => delay6_q_net_x9,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x7,
    delta_y_i => mux3_y_net_x7,
    y_r => mux_y_net_x6,
    y_i => mux1_y_net_x7,
    start_out => delay6_q_net_x7
  );
  bf2i2 : entity xil_defaultlib.pilotdetect_bf2i2_x0
  port map (
    delta_x_r => delay12_q_net,
    delta_x_i => delay11_q_net,
    x_r => delay5_q_net,
    x_i => delay4_q_net,
    start_in => delay2_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x6,
    delta_y_i => mux3_y_net_x6,
    y_r => mux_y_net_x5,
    y_i => mux1_y_net_x6,
    start_out => delay6_q_net_x6
  );
  bf2i3 : entity xil_defaultlib.pilotdetect_bf2i3_x0
  port map (
    delta_x_r => reinterpret3_output_port_net,
    delta_x_i => reinterpret2_output_port_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1,
    start_in => delay24_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x5,
    delta_y_i => mux3_y_net_x5,
    y_r => mux_y_net_x4,
    y_i => mux1_y_net_x5,
    start_out => delay6_q_net_x5
  );
  bf2i4 : entity xil_defaultlib.pilotdetect_bf2i4_x0
  port map (
    delta_x_r => reinterpret3_output_port_net_x1,
    delta_x_i => reinterpret2_output_port_net_x1,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0,
    start_in => delay28_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x4,
    delta_y_i => mux3_y_net_x4,
    y_r => mux_y_net_x3,
    y_i => mux1_y_net_x4,
    start_out => delay6_q_net_x4
  );
  bf2ii : entity xil_defaultlib.pilotdetect_bf2ii_x0
  port map (
    delta_x_r => delay3_q_net,
    delta_x_i => delay2_q_net_x0,
    x_r => mux_y_net_x7,
    x_i => mux1_y_net_x8,
    start_in => delay6_q_net_x8,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x3,
    delta_y_i => mux3_y_net_x3,
    y_r => mux_y_net_x2,
    y_i => mux1_y_net_x3,
    start_out => delay6_q_net_x3
  );
  bf2ii1 : entity xil_defaultlib.pilotdetect_bf2ii1_x0
  port map (
    delta_x_r => delay10_q_net,
    delta_x_i => delay9_q_net,
    x_r => mux_y_net_x6,
    x_i => mux1_y_net_x7,
    start_in => delay6_q_net_x7,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x2,
    delta_y_i => mux3_y_net_x2,
    y_r => mux_y_net_x12,
    y_i => mux1_y_net_x2,
    start_out => delay6_q_net_x2
  );
  bf2ii2 : entity xil_defaultlib.pilotdetect_bf2ii2_x0
  port map (
    delta_x_r => delay14_q_net,
    delta_x_i => delay13_q_net,
    x_r => mux_y_net_x5,
    x_i => mux1_y_net_x6,
    start_in => delay6_q_net_x6,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x1,
    delta_y_i => mux3_y_net_x1,
    y_r => mux_y_net_x1,
    y_i => mux1_y_net_x1,
    start_out => delay6_q_net_x1
  );
  bf2ii3 : entity xil_defaultlib.pilotdetect_bf2ii3_x0
  port map (
    delta_x_r => reinterpret3_output_port_net_x0,
    delta_x_i => reinterpret2_output_port_net_x0,
    x_r => mux_y_net_x4,
    x_i => mux1_y_net_x5,
    start_in => delay6_q_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x0,
    delta_y_i => mux3_y_net_x0,
    y_r => mux_y_net_x0,
    y_i => mux1_y_net_x0,
    start_out => delay6_q_net_x0
  );
  bf2ii4 : entity xil_defaultlib.pilotdetect_bf2ii4_x0
  port map (
    delta_x_r => reinterpret3_output_port_net_x2,
    delta_x_i => reinterpret2_output_port_net_x2,
    x_r => shift_op_net,
    x_i => shift1_op_net,
    start_in => delay18_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net,
    delta_y_i => mux3_y_net,
    y_r => mux_y_net,
    y_i => mux1_y_net,
    start_out => delay6_q_net
  );
  complex_mult : entity xil_defaultlib.pilotdetect_complex_mult_x1
  port map (
    a_r => mux_y_net_x10,
    a_i => mux1_y_net_x11,
    b_r => delay4_q_net_x4,
    b_i => delay5_q_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x3,
    x_i => delay5_q_net_x3
  );
  complex_mult1 : entity xil_defaultlib.pilotdetect_complex_mult1_x1
  port map (
    a_r => mux_y_net_x11,
    a_i => mux1_y_net_x12,
    b_r => delay15_q_net,
    b_i => delay16_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2
  );
  complex_mult2 : entity xil_defaultlib.pilotdetect_complex_mult2_x2
  port map (
    a_r => mux_y_net_x9,
    a_i => mux1_y_net_x10,
    b_r => delay22_q_net,
    b_i => delay23_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1
  );
  complex_mult3 : entity xil_defaultlib.pilotdetect_complex_mult3_x2
  port map (
    a_r => mux_y_net_x8,
    a_i => mux1_y_net_x9,
    b_r => delay19_q_net,
    b_i => delay21_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0
  );
  large_complex_delay : entity xil_defaultlib.pilotdetect_large_complex_delay_x0
  port map (
    in_r => mux3_y_net,
    in_i => mux2_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x2,
    out_i => reinterpret3_output_port_net_x2
  );
  large_complex_delay1 : entity xil_defaultlib.pilotdetect_large_complex_delay1_x0
  port map (
    in_r => mux3_y_net_x4,
    in_i => mux2_y_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x1,
    out_i => reinterpret3_output_port_net_x1
  );
  large_complex_delay4 : entity xil_defaultlib.pilotdetect_large_complex_delay4_x0
  port map (
    in_r => mux3_y_net_x0,
    in_i => mux2_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x0,
    out_i => reinterpret3_output_port_net_x0
  );
  large_complex_delay5 : entity xil_defaultlib.pilotdetect_large_complex_delay5_x0
  port map (
    in_r => mux3_y_net_x5,
    in_i => mux2_y_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net,
    out_i => reinterpret3_output_port_net
  );
  large_inv_tfactor_rom : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom_x0
  port map (
    in1 => delay6_q_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x11,
    w_i => mux1_y_net_x12
  );
  large_inv_tfactor_rom1 : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom1_x0
  port map (
    in1 => delay6_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x10,
    w_i => mux1_y_net_x11
  );
  large_inv_tfactor_rom2 : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom2_x0
  port map (
    in1 => delay6_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x9,
    w_i => mux1_y_net_x10
  );
  small_inv_tfactor_rom4 : entity xil_defaultlib.pilotdetect_small_inv_tfactor_rom4_x0
  port map (
    in1 => delay6_q_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x8,
    w_i => mux1_y_net_x9
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux3_y_net_x6,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux2_y_net_x6,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
  delay16 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  delay17 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay17_q_net
  );
  delay18 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay18_q_net
  );
  delay19 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay19_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay21 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay21_q_net
  );
  delay22 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x12,
    clk => clk_net,
    ce => ce_net,
    q => delay22_q_net
  );
  delay23 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay23_q_net
  );
  delay24 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay24_q_net
  );
  delay28 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay28_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x4
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x4
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x9
  );
  delay7 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  shift : entity xil_defaultlib.sysgen_shift_5fce716372
  port map (
    clr => '0',
    ip => mux_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    op => shift_op_net
  );
  shift1 : entity xil_defaultlib.sysgen_shift_5fce716372
  port map (
    clr => '0',
    ip => mux1_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    op => shift1_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2I
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i_x1;
architecture structural of pilotdetect_bf2i_x1 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay17_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay1_q_net_x0 <= delta_x_r;
  delay_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net_x0 <= x_i;
  delay17_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net_x0,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net_x0,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay1_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay17_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 2,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2I1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i1_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i1_x1;
architecture structural of pilotdetect_bf2i1_x1 is
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay8_q_net <= delta_x_r;
  delay7_q_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net_x0 <= x_i;
  delay6_q_net_x0 <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay8_q_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay7_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay8_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay7_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 17,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 4,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2I2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i2_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i2_x1;
architecture structural of pilotdetect_bf2i2_x1 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal clk_net : std_logic;
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  delay12_q_net <= delta_x_r;
  delay11_q_net <= delta_x_i;
  delay5_q_net_x0 <= x_r;
  delay4_q_net_x0 <= x_i;
  delay2_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay12_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay12_q_net,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay11_q_net,
    b => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay12_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay11_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay2_q_net_x0,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net,
    d0 => delay4_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2I3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i3_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i3_x1;
architecture structural of pilotdetect_bf2i3_x1 is
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay24_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 65,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay24_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 6,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2I4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2i4_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2i4_x1;
architecture structural of pilotdetect_bf2i4_x1 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  start_out <= delay6_q_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  delay4_q_net <= x_r;
  delay5_q_net <= x_i;
  delay28_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay5_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x0
  );
  delay5 : entity xil_defaultlib.sysgen_delay_3791cc6a11
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x0
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 257,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay28_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay1_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay2_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay3_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay5_q_net_x0,
    d0 => delay4_q_net_x0,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 8,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2II
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii_x1;
architecture structural of pilotdetect_bf2ii_x1 is
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay3_q_net_x0 <= delta_x_r;
  delay2_q_net_x0 <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net_x0,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net_x0,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net_x0,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay2_q_net_x0,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay3_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay2_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 10,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 3,
    new_msb => 3,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 2,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2II1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii1_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii1_x1;
architecture structural of pilotdetect_bf2ii1_x1 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay10_q_net <= delta_x_r;
  delay9_q_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay10_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay9_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay10_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay9_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 34,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 5,
    new_msb => 5,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 4,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2II2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii2_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii2_x1;
architecture structural of pilotdetect_bf2ii2_x1 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  delay14_q_net <= delta_x_r;
  delay13_q_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay14_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay14_q_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay13_q_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay13_q_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay14_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay13_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 1,
    new_msb => 1,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 0,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2II3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii3_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 );
    start_out : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_bf2ii3_x1;
architecture structural of pilotdetect_bf2ii3_x1 is
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net_x0;
  y_i <= mux1_y_net_x0;
  start_out <= delay6_q_net_x0;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  mux_y_net <= x_r;
  mux1_y_net <= x_i;
  delay6_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 130,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x0
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net_x0
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux_y_net,
    d1 => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => mux1_y_net,
    d1 => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 7,
    new_msb => 7,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 6,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/BF2II4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_bf2ii4_x1 is
  port (
    delta_x_r : in std_logic_vector( 18-1 downto 0 );
    delta_x_i : in std_logic_vector( 18-1 downto 0 );
    x_r : in std_logic_vector( 18-1 downto 0 );
    x_i : in std_logic_vector( 18-1 downto 0 );
    start_in : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    delta_y_r : out std_logic_vector( 18-1 downto 0 );
    delta_y_i : out std_logic_vector( 18-1 downto 0 );
    y_r : out std_logic_vector( 18-1 downto 0 );
    y_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_bf2ii4_x1;
architecture structural of pilotdetect_bf2ii4_x1 is
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
begin
  delta_y_r <= mux2_y_net;
  delta_y_i <= mux3_y_net;
  y_r <= mux_y_net;
  y_i <= mux1_y_net;
  reinterpret3_output_port_net <= delta_x_r;
  reinterpret2_output_port_net <= delta_x_i;
  shift_op_net <= x_r;
  shift1_op_net <= x_i;
  delay18_q_net <= start_in;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret3_output_port_net,
    b => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsubmode
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i4",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    mode_arith => xlUnsigned,
    mode_bin_pt => 0,
    mode_width => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => reinterpret2_output_port_net,
    b => mux5_y_net,
    mode => delay4_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay18_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay7 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  expression : entity xil_defaultlib.sysgen_expr_1fcd00473b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_8a1084dbe1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => slice_y_net,
    b => slice1_y_net,
    dout => expression1_dout_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay3_q_net,
    d1 => addsub_s_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay5_q_net,
    d1 => addsub4_s_net,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay7_q_net,
    d1 => addsub1_s_net,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => delay8_q_net,
    d1 => addsub2_s_net,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift_op_net,
    d1 => shift1_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => expression_dout_net,
    d0 => shift1_op_net,
    d1 => shift_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux5_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 9,
    new_msb => 9,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 8,
    x_width => 10,
    y_width => 1
  )
  port map (
    x => counter_op_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/complex_mult
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult_x2 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult_x2;
architecture structural of pilotdetect_complex_mult_x2 is
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay4_q_net_x0 <= b_r;
  delay5_q_net_x0 <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay4_q_net_x0,
    b => delay5_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay4_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/complex_mult1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult1_x2 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult1_x2;
architecture structural of pilotdetect_complex_mult1_x2 is
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay15_q_net <= b_r;
  delay16_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay15_q_net,
    b => delay16_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay15_q_net,
    b => delay16_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay15_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/complex_mult2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult2_x3 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult2_x3;
architecture structural of pilotdetect_complex_mult2_x3 is
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay22_q_net <= b_r;
  delay23_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay22_q_net,
    b => delay23_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay22_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/complex_mult3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult3_x3 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult3_x3;
architecture structural of pilotdetect_complex_mult3_x3 is
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay19_q_net <= b_r;
  delay21_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay19_q_net,
    b => delay21_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay19_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_complex_delay
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay_x1 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay_x1;
architecture structural of pilotdetect_large_complex_delay_x1 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 9-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i0",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i1",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_complex_delay1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay1_x1 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay1_x1;
architecture structural of pilotdetect_large_complex_delay1_x1 is
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal ce_net : std_logic;
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 8-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 8-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 8,
    c_address_width_b => 8,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i1",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i2",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i3",
    op_arith => xlUnsigned,
    op_width => 8
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_complex_delay4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay4_x1 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay4_x1;
architecture structural of pilotdetect_large_complex_delay4_x1 is
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 7-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 7-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i2",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i4",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i5",
    op_arith => xlUnsigned,
    op_width => 7
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_complex_delay5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_complex_delay5_x1 is
  port (
    in_r : in std_logic_vector( 18-1 downto 0 );
    in_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out_r : out std_logic_vector( 18-1 downto 0 );
    out_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_complex_delay5_x1;
architecture structural of pilotdetect_large_complex_delay5_x1 is
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal constant_op_net : std_logic_vector( 36-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 36-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 36-1 downto 0 );
  signal output_addr_op_net : std_logic_vector( 6-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal output_addr1_op_net : std_logic_vector( 6-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
begin
  out_r <= reinterpret2_output_port_net;
  out_i <= reinterpret3_output_port_net;
  mux3_y_net <= in_r;
  mux2_y_net <= in_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7dc385d728
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => slice1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 6,
    c_address_width_b => 6,
    c_width_a => 36,
    c_width_b => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i3",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => output_addr1_op_net,
    dina => concat_y_net,
    wea => constant2_op_net,
    addrb => output_addr_op_net,
    dinb => constant_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  output_addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i6",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr_op_net
  );
  output_addr1 : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i7",
    op_arith => xlUnsigned,
    op_width => 6
  )
  port map (
    en => "1",
    rst => "0",
    clr => '0',
    clk => clk_net,
    ce => ce_net,
    op => output_addr1_op_net
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux3_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux2_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay_q_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => delay1_q_net,
    output_port => reinterpret3_output_port_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => dual_port_ram_doutb_net,
    y => slice1_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_inv_tfactor_rom/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x12 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 10-1 downto 0 )
  );
end pilotdetect_address_generator_x12;
architecture structural of pilotdetect_address_generator_x12 is
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 10-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub_s_net : std_logic_vector( 10-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 10-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 10-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 8-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 10-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 10-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant_op_net : std_logic_vector( 10-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 10,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 10,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 11,
    core_name0 => "pilotdetect_c_addsub_v12_0_i2",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 11,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 10
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b834ce322d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_65e9092d81
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_f84e73127e
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_377354b5ea
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_81939abd89
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 9,
    x_width => 10,
    y_width => 10
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_inv_tfactor_rom
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom_x1 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom_x1;
architecture structural of pilotdetect_large_inv_tfactor_rom_x1 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 10-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 9-1 downto 0 );
  signal slice_y_net : std_logic_vector( 8-1 downto 0 );
  signal delay_q_net : std_logic_vector( 10-1 downto 0 );
  signal concat_y_net : std_logic_vector( 9-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x12
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_222d6d85fc
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_57ee5c1d4b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 10
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 9,
    c_address_width_b => 9,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i4",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 8,
    new_msb => 9,
    x_width => 10,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_inv_tfactor_rom1/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x13 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 8-1 downto 0 )
  );
end pilotdetect_address_generator_x13;
architecture structural of pilotdetect_address_generator_x13 is
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal clk_net : std_logic;
  signal concat3_y_net : std_logic_vector( 8-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 8-1 downto 0 );
  signal mux_y_net : std_logic_vector( 8-1 downto 0 );
  signal constant_op_net : std_logic_vector( 8-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 6-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 8-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 8-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 8,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 8,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 9,
    core_name0 => "pilotdetect_c_addsub_v12_0_i3",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 9,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 8
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_2b7c6b2428
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_a8c933a1a7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_b4de442209
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_78f34e96e5
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_4b3c2484ae
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 7,
    x_width => 10,
    y_width => 8
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_inv_tfactor_rom1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom1_x1 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom1_x1;
architecture structural of pilotdetect_large_inv_tfactor_rom1_x1 is
  signal delay_q_net : std_logic_vector( 8-1 downto 0 );
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 7-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 7-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 8-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 6-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x13
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_2e499fd69d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_3e7267ab01
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 8
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 7,
    c_address_width_b => 7,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i5",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 8,
    y_width => 6
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 6,
    new_msb => 7,
    x_width => 8,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_inv_tfactor_rom2/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator_x14 is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 6-1 downto 0 )
  );
end pilotdetect_address_generator_x14;
architecture structural of pilotdetect_address_generator_x14 is
  signal clk_net : std_logic;
  signal mux_y_net : std_logic_vector( 6-1 downto 0 );
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 6-1 downto 0 );
  signal concat2_y_net : std_logic_vector( 6-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 6-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant_op_net : std_logic_vector( 6-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 6-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 6,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 6,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 7,
    core_name0 => "pilotdetect_c_addsub_v12_0_i5",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 7,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 6
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_392cf7ce5c
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_4adcefda0f
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_a152b8b4ce
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_7d4cdb5bbb
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bba3bd89f4
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 5,
    x_width => 10,
    y_width => 6
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/large_inv_tfactor_rom2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_large_inv_tfactor_rom2_x1 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_large_inv_tfactor_rom2_x1;
architecture structural of pilotdetect_large_inv_tfactor_rom2_x1 is
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal ce_net : std_logic;
  signal concat_y_net : std_logic_vector( 5-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 5-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 6-1 downto 0 );
  signal slice_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal delay_q_net : std_logic_vector( 6-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator_x14
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_c024ed0ea3
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_b172047307
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 6
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 5,
    c_address_width_b => 5,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i6",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    dinb => constant2_op_net,
    web => constant1_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 6,
    y_width => 4
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 4,
    new_msb => 5,
    x_width => 6,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/small_inv_tfactor_rom4/address_generator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_address_generator is
  port (
    in1 : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    out1 : out std_logic_vector( 4-1 downto 0 )
  );
end pilotdetect_address_generator;
architecture structural of pilotdetect_address_generator is
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal mux_y_net : std_logic_vector( 4-1 downto 0 );
  signal clk_net : std_logic;
  signal concat2_y_net : std_logic_vector( 4-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 2-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 4-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat1_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant_op_net : std_logic_vector( 4-1 downto 0 );
  signal ce_net : std_logic;
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal concat3_y_net : std_logic_vector( 4-1 downto 0 );
  signal constant4_op_net : std_logic_vector( 2-1 downto 0 );
  signal constant3_op_net : std_logic_vector( 2-1 downto 0 );
  signal slice2_y_net : std_logic_vector( 4-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
begin
  out1 <= mux_y_net;
  counter_op_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlUnsigned,
    a_bin_pt => 0,
    a_width => 4,
    b_arith => xlUnsigned,
    b_bin_pt => 0,
    b_width => 4,
    c_has_c_out => 0,
    c_latency => 0,
    c_output_width => 5,
    core_name0 => "pilotdetect_c_addsub_v12_0_i6",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 5,
    latency => 0,
    overflow => 3,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 0,
    s_width => 4
  )
  port map (
    clr => '0',
    en => "1",
    a => concat3_y_net,
    b => concat2_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice1_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_6a9e537061
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => concat_y_net,
    in1 => constant2_op_net,
    y => concat1_y_net
  );
  concat2 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant3_op_net,
    in1 => slice1_y_net,
    y => concat2_y_net
  );
  concat3 : entity xil_defaultlib.sysgen_concat_059a3b2d1a
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => slice1_y_net,
    in1 => constant4_op_net,
    y => concat3_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_55eaac7d5b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  constant3 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant3_op_net
  );
  constant4 : entity xil_defaultlib.sysgen_constant_b2984b3948
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant4_op_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => counter_op_net,
    a_br => mcode_a_br_net
  );
  mux : entity xil_defaultlib.sysgen_mux_bb4a1d2355
  port map (
    clr => '0',
    sel => slice_y_net,
    d0 => constant_op_net,
    d1 => concat1_y_net,
    d2 => concat2_y_net,
    d3 => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => slice2_y_net,
    y => slice1_y_net
  );
  slice2 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 3,
    x_width => 10,
    y_width => 4
  )
  port map (
    x => mcode_a_br_net,
    y => slice2_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3/small_inv_tfactor_rom4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_small_inv_tfactor_rom4_x1 is
  port (
    in1 : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    w_r : out std_logic_vector( 18-1 downto 0 );
    w_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_small_inv_tfactor_rom4_x1;
architecture structural of pilotdetect_small_inv_tfactor_rom4_x1 is
  signal counter_op_net : std_logic_vector( 10-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 4-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal concat_y_net : std_logic_vector( 3-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 2-1 downto 0 );
  signal ce_net : std_logic;
  signal concat1_y_net : std_logic_vector( 3-1 downto 0 );
  signal constant2_op_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_douta_net : std_logic_vector( 18-1 downto 0 );
  signal a_y_net : std_logic_vector( 2-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal dual_port_ram_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 4-1 downto 0 );
  signal negate1_op_net : std_logic_vector( 18-1 downto 0 );
begin
  w_r <= mux_y_net;
  w_i <= mux1_y_net;
  delay6_q_net <= in1;
  clk_net <= clk_1;
  ce_net <= ce_1;
  address_generator : entity xil_defaultlib.pilotdetect_address_generator
  port map (
    in1 => counter_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out1 => mux_y_net_x0
  );
  concat : entity xil_defaultlib.sysgen_concat_1672b64d97
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant1_op_net,
    in1 => slice_y_net,
    y => concat_y_net
  );
  concat1 : entity xil_defaultlib.sysgen_concat_83b84ba15d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => constant_op_net,
    in1 => slice_y_net,
    y => concat1_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_ba5259fe63
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  constant2 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant2_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay6_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 4
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  dual_port_ram : entity xil_defaultlib.pilotdetect_xldpram_dist
  generic map (
    addr_width => 3,
    c_address_width => 4,
    c_width => 18,
    core_name0 => "pilotdetect_dist_mem_gen_v8_0_i1",
    latency => 2
  )
  port map (
    ena => "1",
    enb => "1",
    addra => concat_y_net,
    dina => constant2_op_net,
    wea => constant1_op_net,
    addrb => concat1_y_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => dual_port_ram_douta_net,
    doutb => dual_port_ram_doutb_net
  );
  mux : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_douta_net,
    d1 => dual_port_ram_doutb_net,
    d2 => negate1_op_net,
    d3 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_2039aba8d7
  port map (
    clr => '0',
    sel => a_y_net,
    d0 => dual_port_ram_doutb_net,
    d1 => negate1_op_net,
    d2 => negate_op_net,
    d3 => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_doutb_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
  negate1 : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => dual_port_ram_douta_net,
    clk => clk_net,
    ce => ce_net,
    op => negate1_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 1,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => mux_y_net_x0,
    y => slice_y_net
  );
  a : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 2,
    new_msb => 3,
    x_width => 4,
    y_width => 2
  )
  port map (
    x => delay_q_net,
    y => a_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_1024_ver_3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_ifft_1024_ver_3 is
  port (
    x_r_x0 : in std_logic_vector( 18-1 downto 0 );
    x_i_x0 : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_ifft_1024_ver_3;
architecture structural of pilotdetect_ifft_1024_ver_3 is
  signal mux_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x9 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay15_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay21_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay18_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay28_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay14_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal shift_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal shift1_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay22_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay23_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay19_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay13_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay16_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x10 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal mux3_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x12 : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux1_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal delay11_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay12_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x8 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x6 : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x8 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x7 : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x6 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal delay7_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay17_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay24_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux2_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x5 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net_x7 : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net_x9 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x6 : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= mux1_y_net;
  x_i <= mux_y_net;
  delay4_q_net <= x_r_x0;
  delay5_q_net <= x_i_x0;
  delay2_q_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  bf2i : entity xil_defaultlib.pilotdetect_bf2i_x1
  port map (
    delta_x_r => delay1_q_net,
    delta_x_i => delay_q_net,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2,
    start_in => delay17_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x8,
    delta_y_i => mux3_y_net_x8,
    y_r => mux_y_net_x7,
    y_i => mux1_y_net_x8,
    start_out => delay6_q_net_x8
  );
  bf2i1 : entity xil_defaultlib.pilotdetect_bf2i1_x1
  port map (
    delta_x_r => delay8_q_net,
    delta_x_i => delay7_q_net,
    x_r => delay4_q_net_x3,
    x_i => delay5_q_net_x3,
    start_in => delay6_q_net_x9,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x7,
    delta_y_i => mux3_y_net_x7,
    y_r => mux_y_net_x6,
    y_i => mux1_y_net_x7,
    start_out => delay6_q_net_x7
  );
  bf2i2 : entity xil_defaultlib.pilotdetect_bf2i2_x1
  port map (
    delta_x_r => delay12_q_net,
    delta_x_i => delay11_q_net,
    x_r => delay5_q_net,
    x_i => delay4_q_net,
    start_in => delay2_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x6,
    delta_y_i => mux3_y_net_x6,
    y_r => mux_y_net_x5,
    y_i => mux1_y_net_x6,
    start_out => delay6_q_net_x6
  );
  bf2i3 : entity xil_defaultlib.pilotdetect_bf2i3_x1
  port map (
    delta_x_r => reinterpret3_output_port_net,
    delta_x_i => reinterpret2_output_port_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1,
    start_in => delay24_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x5,
    delta_y_i => mux3_y_net_x5,
    y_r => mux_y_net_x4,
    y_i => mux1_y_net_x5,
    start_out => delay6_q_net_x5
  );
  bf2i4 : entity xil_defaultlib.pilotdetect_bf2i4_x1
  port map (
    delta_x_r => reinterpret3_output_port_net_x1,
    delta_x_i => reinterpret2_output_port_net_x1,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0,
    start_in => delay28_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x4,
    delta_y_i => mux3_y_net_x4,
    y_r => mux_y_net_x3,
    y_i => mux1_y_net_x4,
    start_out => delay6_q_net_x4
  );
  bf2ii : entity xil_defaultlib.pilotdetect_bf2ii_x1
  port map (
    delta_x_r => delay3_q_net,
    delta_x_i => delay2_q_net_x0,
    x_r => mux_y_net_x7,
    x_i => mux1_y_net_x8,
    start_in => delay6_q_net_x8,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x3,
    delta_y_i => mux3_y_net_x3,
    y_r => mux_y_net_x2,
    y_i => mux1_y_net_x3,
    start_out => delay6_q_net_x3
  );
  bf2ii1 : entity xil_defaultlib.pilotdetect_bf2ii1_x1
  port map (
    delta_x_r => delay10_q_net,
    delta_x_i => delay9_q_net,
    x_r => mux_y_net_x6,
    x_i => mux1_y_net_x7,
    start_in => delay6_q_net_x7,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x2,
    delta_y_i => mux3_y_net_x2,
    y_r => mux_y_net_x12,
    y_i => mux1_y_net_x2,
    start_out => delay6_q_net_x2
  );
  bf2ii2 : entity xil_defaultlib.pilotdetect_bf2ii2_x1
  port map (
    delta_x_r => delay14_q_net,
    delta_x_i => delay13_q_net,
    x_r => mux_y_net_x5,
    x_i => mux1_y_net_x6,
    start_in => delay6_q_net_x6,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x1,
    delta_y_i => mux3_y_net_x1,
    y_r => mux_y_net_x1,
    y_i => mux1_y_net_x1,
    start_out => delay6_q_net_x1
  );
  bf2ii3 : entity xil_defaultlib.pilotdetect_bf2ii3_x1
  port map (
    delta_x_r => reinterpret3_output_port_net_x0,
    delta_x_i => reinterpret2_output_port_net_x0,
    x_r => mux_y_net_x4,
    x_i => mux1_y_net_x5,
    start_in => delay6_q_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net_x0,
    delta_y_i => mux3_y_net_x0,
    y_r => mux_y_net_x0,
    y_i => mux1_y_net_x0,
    start_out => delay6_q_net_x0
  );
  bf2ii4 : entity xil_defaultlib.pilotdetect_bf2ii4_x1
  port map (
    delta_x_r => reinterpret3_output_port_net_x2,
    delta_x_i => reinterpret2_output_port_net_x2,
    x_r => shift_op_net,
    x_i => shift1_op_net,
    start_in => delay18_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    delta_y_r => mux2_y_net,
    delta_y_i => mux3_y_net,
    y_r => mux_y_net,
    y_i => mux1_y_net
  );
  complex_mult : entity xil_defaultlib.pilotdetect_complex_mult_x2
  port map (
    a_r => mux_y_net_x10,
    a_i => mux1_y_net_x11,
    b_r => delay4_q_net_x4,
    b_i => delay5_q_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x3,
    x_i => delay5_q_net_x3
  );
  complex_mult1 : entity xil_defaultlib.pilotdetect_complex_mult1_x2
  port map (
    a_r => mux_y_net_x11,
    a_i => mux1_y_net_x12,
    b_r => delay15_q_net,
    b_i => delay16_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x2,
    x_i => delay5_q_net_x2
  );
  complex_mult2 : entity xil_defaultlib.pilotdetect_complex_mult2_x3
  port map (
    a_r => mux_y_net_x9,
    a_i => mux1_y_net_x10,
    b_r => delay22_q_net,
    b_i => delay23_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1
  );
  complex_mult3 : entity xil_defaultlib.pilotdetect_complex_mult3_x3
  port map (
    a_r => mux_y_net_x8,
    a_i => mux1_y_net_x9,
    b_r => delay19_q_net,
    b_i => delay21_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0
  );
  large_complex_delay : entity xil_defaultlib.pilotdetect_large_complex_delay_x1
  port map (
    in_r => mux3_y_net,
    in_i => mux2_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x2,
    out_i => reinterpret3_output_port_net_x2
  );
  large_complex_delay1 : entity xil_defaultlib.pilotdetect_large_complex_delay1_x1
  port map (
    in_r => mux3_y_net_x4,
    in_i => mux2_y_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x1,
    out_i => reinterpret3_output_port_net_x1
  );
  large_complex_delay4 : entity xil_defaultlib.pilotdetect_large_complex_delay4_x1
  port map (
    in_r => mux3_y_net_x0,
    in_i => mux2_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net_x0,
    out_i => reinterpret3_output_port_net_x0
  );
  large_complex_delay5 : entity xil_defaultlib.pilotdetect_large_complex_delay5_x1
  port map (
    in_r => mux3_y_net_x5,
    in_i => mux2_y_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    out_r => reinterpret2_output_port_net,
    out_i => reinterpret3_output_port_net
  );
  large_inv_tfactor_rom : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom_x1
  port map (
    in1 => delay6_q_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x11,
    w_i => mux1_y_net_x12
  );
  large_inv_tfactor_rom1 : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom1_x1
  port map (
    in1 => delay6_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x10,
    w_i => mux1_y_net_x11
  );
  large_inv_tfactor_rom2 : entity xil_defaultlib.pilotdetect_large_inv_tfactor_rom2_x1
  port map (
    in1 => delay6_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x9,
    w_i => mux1_y_net_x10
  );
  small_inv_tfactor_rom4 : entity xil_defaultlib.pilotdetect_small_inv_tfactor_rom4_x1
  port map (
    in1 => delay6_q_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    w_r => mux_y_net_x8,
    w_i => mux1_y_net_x9
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x8,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay10 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay11 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux3_y_net_x6,
    q => delay11_q_net
  );
  delay12 : entity xil_defaultlib.sysgen_delay_2eaa039003
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d => mux2_y_net_x6,
    q => delay12_q_net
  );
  delay13 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay13_q_net
  );
  delay14 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay14_q_net
  );
  delay15 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay15_q_net
  );
  delay16 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay16_q_net
  );
  delay17 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay17_q_net
  );
  delay18 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x4,
    clk => clk_net,
    ce => ce_net,
    q => delay18_q_net
  );
  delay19 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay19_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net_x0
  );
  delay21 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay21_q_net
  );
  delay22 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x12,
    clk => clk_net,
    ce => ce_net,
    q => delay22_q_net
  );
  delay23 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay23_q_net
  );
  delay24 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay24_q_net
  );
  delay28 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay28_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 7,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net_x4
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 4,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net_x4
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 11,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net_x9
  );
  delay7 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay7_q_net
  );
  delay8 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 15,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux2_y_net_x7,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 31,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux3_y_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  shift : entity xil_defaultlib.sysgen_shift_5fce716372
  port map (
    clr => '0',
    ip => mux_y_net_x3,
    clk => clk_net,
    ce => ce_net,
    op => shift_op_net
  );
  shift1 : entity xil_defaultlib.sysgen_shift_5fce716372
  port map (
    clr => '0',
    ip => mux1_y_net_x4,
    clk => clk_net,
    ce => ce_net,
    op => shift1_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/IFFT_input_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_ifft_input_control is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    read_addr : out std_logic_vector( 10-1 downto 0 );
    read_addr_reversed : out std_logic_vector( 10-1 downto 0 );
    h_sel : out std_logic_vector( 1-1 downto 0 );
    ifft_start : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_ifft_input_control;
architecture structural of pilotdetect_ifft_input_control is
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal start_ifft_1_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal constant_op_net : std_logic_vector( 10-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal finish_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addr_op_net : std_logic_vector( 10-1 downto 0 );
  signal read_1_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal expression3_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression2_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression4_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression5_dout_net : std_logic_vector( 1-1 downto 0 );
  signal read_0_reg_q_net : std_logic_vector( 1-1 downto 0 );
begin
  read_addr <= addr_op_net;
  read_addr_reversed <= mcode_a_br_net;
  h_sel <= logical1_y_net;
  ifft_start <= expression1_dout_net;
  delay_q_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant_x0 : entity xil_defaultlib.sysgen_constant_734763fe12
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  expression : entity xil_defaultlib.sysgen_expr_c9661e2436
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    finish => finish_reg_q_net,
    start => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_ba1420c02b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    finish => finish_reg_q_net,
    start => delay_q_net,
    start_ifft_1 => start_ifft_1_reg_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression1_dout_net
  );
  expression2 : entity xil_defaultlib.sysgen_expr_a42a5f85e1
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    finish => finish_reg_q_net,
    r_addr_eq_1022 => relational_op_net,
    read_0 => read_0_reg_q_net,
    start => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression2_dout_net
  );
  expression3 : entity xil_defaultlib.sysgen_expr_b4b1b8224d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    r_addr_eq_1022 => relational_op_net,
    read_0 => read_0_reg_q_net,
    dout => expression3_dout_net
  );
  expression4 : entity xil_defaultlib.sysgen_expr_34a27e207b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    r_addr_eq_1022 => relational_op_net,
    read_1 => read_1_reg_q_net,
    start_ifft_1 => start_ifft_1_reg_q_net,
    dout => expression4_dout_net
  );
  expression5 : entity xil_defaultlib.sysgen_expr_a0374b5183
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    r_addr_eq_1022 => relational_op_net,
    read_1 => read_1_reg_q_net,
    dout => expression5_dout_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_5ceae8d63b
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d0 => read_1_reg_q_net,
    d1 => finish_reg_q_net,
    y => logical1_y_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_7a50437cc6
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => addr_op_net,
    a_br => mcode_a_br_net
  );
  relational : entity xil_defaultlib.sysgen_relational_a77d10299f
  port map (
    clr => '0',
    a => addr_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i8",
    op_arith => xlUnsigned,
    op_width => 10
  )
  port map (
    en => "1",
    clr => '0',
    rst => delay_q_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  finish_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression5_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => finish_reg_q_net
  );
  read_0_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression2_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => read_0_reg_q_net
  );
  read_1_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression4_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => read_1_reg_q_net
  );
  start_ifft_1_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression3_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => start_ifft_1_reg_q_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/OnA_input_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_ona_input_control is
  port (
    s : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    r0 : out std_logic_vector( 1-1 downto 0 );
    r1 : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_ona_input_control;
architecture structural of pilotdetect_ona_input_control is
  signal delay6_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal r1_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal r0_reg_q_net : std_logic_vector( 1-1 downto 0 );
begin
  r0 <= logical_y_net;
  r1 <= logical1_y_net;
  delay6_q_net <= s;
  clk_net <= clk_1;
  ce_net <= ce_1;
  expression : entity xil_defaultlib.sysgen_expr_745d7733b5
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    r0 => r0_reg_q_net,
    r1 => r1_reg_q_net,
    s => delay6_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_c938aa3d94
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    r0 => r0_reg_q_net,
    r1 => r1_reg_q_net,
    s => delay6_q_net,
    dout => expression1_dout_net
  );
  logical : entity xil_defaultlib.sysgen_logical_b6ae4784bd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d0 => r0_reg_q_net,
    d1 => delay6_q_net,
    y => logical_y_net
  );
  logical1 : entity xil_defaultlib.sysgen_logical_b6ae4784bd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    d0 => r1_reg_q_net,
    d1 => delay6_q_net,
    y => logical1_y_net
  );
  r0_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => r0_reg_q_net
  );
  r1_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => r1_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add/section_adder
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_section_adder is
  port (
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output_r : out std_logic_vector( 18-1 downto 0 );
    output_i : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_section_adder;
architecture structural of pilotdetect_section_adder is
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_buf_we_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal mcode_rst_addr_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_output_valid_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal buf_r_data_out_net : std_logic_vector( 36-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
begin
  output_r <= mux_y_net_x0;
  output_i <= mux1_y_net_x0;
  output_valid <= delay2_q_net;
  mux1_y_net <= input_r;
  mux_y_net <= input_i;
  logical_y_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => mcode_output_valid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_66bf1a97d1
  port map (
    clr => '0',
    start => logical_y_net,
    addr_eq_511 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    buf_we => mcode_buf_we_net,
    output_valid => mcode_output_valid_net,
    rst_addr => mcode_rst_addr_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub1_s_net,
    y => mux1_y_net_x0
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux1_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret3_output_port_net
  );
  relational : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => constant_op_net,
    b => addr_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice1_y_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => mcode_rst_addr_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  buf_r : entity xil_defaultlib.pilotdetect_xlspram
  generic map (
    c_address_width => 9,
    c_width => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i7",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_op_net,
    data_in => concat_y_net,
    we => mcode_buf_we_net,
    clk => clk_net,
    ce => ce_net,
    data_out => buf_r_data_out_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_overlap_and_add is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_overlap_and_add;
architecture structural of pilotdetect_overlap_and_add is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
begin
  output <= addsub_s_net;
  output_valid <= delay_q_net;
  logical_y_net <= start;
  mux1_y_net_x0 <= input_r;
  mux_y_net_x0 <= input_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  section_adder : entity xil_defaultlib.pilotdetect_section_adder
  port map (
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    start => logical_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output_r => mux_y_net,
    output_i => mux1_y_net,
    output_valid => delay2_q_net
  );
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 17,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 17,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 2,
    overflow => 2,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 17,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux_y_net,
    b => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux1_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add1/section_adder
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_section_adder_x0 is
  port (
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output_r : out std_logic_vector( 18-1 downto 0 );
    output_i : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_section_adder_x0;
architecture structural of pilotdetect_section_adder_x0 is
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_buf_we_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal mcode_output_valid_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_rst_addr_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal buf_r_data_out_net : std_logic_vector( 36-1 downto 0 );
begin
  output_r <= mux_y_net_x0;
  output_i <= mux1_y_net_x0;
  output_valid <= delay2_q_net;
  mux1_y_net <= input_r;
  mux_y_net <= input_i;
  logical1_y_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => mcode_output_valid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_66bf1a97d1
  port map (
    clr => '0',
    start => logical1_y_net,
    addr_eq_511 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    buf_we => mcode_buf_we_net,
    output_valid => mcode_output_valid_net,
    rst_addr => mcode_rst_addr_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub1_s_net,
    y => mux1_y_net_x0
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux1_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret3_output_port_net
  );
  relational : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => constant_op_net,
    b => addr_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice1_y_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => mcode_rst_addr_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  buf_r : entity xil_defaultlib.pilotdetect_xlspram
  generic map (
    c_address_width => 9,
    c_width => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i7",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_op_net,
    data_in => concat_y_net,
    we => mcode_buf_we_net,
    clk => clk_net,
    ce => ce_net,
    data_out => buf_r_data_out_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_overlap_and_add1 is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_overlap_and_add1;
architecture structural of pilotdetect_overlap_and_add1 is
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
begin
  output <= addsub_s_net;
  output_valid <= delay_q_net;
  logical1_y_net <= start;
  mux1_y_net_x0 <= input_r;
  mux_y_net_x0 <= input_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  section_adder : entity xil_defaultlib.pilotdetect_section_adder_x0
  port map (
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    start => logical1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output_r => mux_y_net,
    output_i => mux1_y_net,
    output_valid => delay2_q_net
  );
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 17,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 17,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 2,
    overflow => 2,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 17,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux_y_net,
    b => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux1_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add2/section_adder
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_section_adder_x1 is
  port (
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output_r : out std_logic_vector( 18-1 downto 0 );
    output_i : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_section_adder_x1;
architecture structural of pilotdetect_section_adder_x1 is
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_output_valid_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_rst_addr_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal buf_r_data_out_net : std_logic_vector( 36-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal mcode_buf_we_net : std_logic_vector( 1-1 downto 0 );
begin
  output_r <= mux_y_net_x0;
  output_i <= mux1_y_net_x0;
  output_valid <= delay2_q_net;
  mux1_y_net <= input_r;
  mux_y_net <= input_i;
  logical_y_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => mcode_output_valid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_66bf1a97d1
  port map (
    clr => '0',
    start => logical_y_net,
    addr_eq_511 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    buf_we => mcode_buf_we_net,
    output_valid => mcode_output_valid_net,
    rst_addr => mcode_rst_addr_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub1_s_net,
    y => mux1_y_net_x0
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux1_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret3_output_port_net
  );
  relational : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => constant_op_net,
    b => addr_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice1_y_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => mcode_rst_addr_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  buf_r : entity xil_defaultlib.pilotdetect_xlspram
  generic map (
    c_address_width => 9,
    c_width => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i7",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_op_net,
    data_in => concat_y_net,
    we => mcode_buf_we_net,
    clk => clk_net,
    ce => ce_net,
    data_out => buf_r_data_out_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_overlap_and_add2 is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_overlap_and_add2;
architecture structural of pilotdetect_overlap_and_add2 is
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
begin
  output <= addsub_s_net;
  output_valid <= delay_q_net;
  logical_y_net <= start;
  mux1_y_net_x0 <= input_r;
  mux_y_net_x0 <= input_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  section_adder : entity xil_defaultlib.pilotdetect_section_adder_x1
  port map (
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    start => logical_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output_r => mux_y_net,
    output_i => mux1_y_net,
    output_valid => delay2_q_net
  );
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 17,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 17,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 2,
    overflow => 2,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 17,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 3,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux_y_net,
    b => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux1_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add3/section_adder
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_section_adder_x2 is
  port (
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output_r : out std_logic_vector( 18-1 downto 0 );
    output_i : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_section_adder_x2;
architecture structural of pilotdetect_section_adder_x2 is
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal buf_r_data_out_net : std_logic_vector( 36-1 downto 0 );
  signal mcode_rst_addr_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_buf_we_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal mcode_output_valid_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
begin
  output_r <= mux_y_net_x0;
  output_i <= mux1_y_net_x0;
  output_valid <= delay2_q_net;
  mux1_y_net <= input_r;
  mux_y_net <= input_i;
  logical1_y_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => mcode_output_valid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_66bf1a97d1
  port map (
    clr => '0',
    start => logical1_y_net,
    addr_eq_511 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    buf_we => mcode_buf_we_net,
    output_valid => mcode_output_valid_net,
    rst_addr => mcode_rst_addr_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub1_s_net,
    y => mux1_y_net_x0
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux1_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret3_output_port_net
  );
  relational : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => constant_op_net,
    b => addr_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice1_y_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => mcode_rst_addr_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  buf_r : entity xil_defaultlib.pilotdetect_xlspram
  generic map (
    c_address_width => 9,
    c_width => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i7",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_op_net,
    data_in => concat_y_net,
    we => mcode_buf_we_net,
    clk => clk_net,
    ce => ce_net,
    data_out => buf_r_data_out_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_overlap_and_add3 is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_overlap_and_add3;
architecture structural of pilotdetect_overlap_and_add3 is
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
begin
  output <= addsub_s_net;
  output_valid <= delay_q_net;
  logical1_y_net <= start;
  mux1_y_net_x0 <= input_r;
  mux_y_net_x0 <= input_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  section_adder : entity xil_defaultlib.pilotdetect_section_adder_x2
  port map (
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    start => logical1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output_r => mux_y_net,
    output_i => mux1_y_net,
    output_valid => delay2_q_net
  );
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 17,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 17,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 2,
    overflow => 2,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 17,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux_y_net,
    b => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux1_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add4/section_adder
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_section_adder_x3 is
  port (
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output_r : out std_logic_vector( 18-1 downto 0 );
    output_i : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_section_adder_x3;
architecture structural of pilotdetect_section_adder_x3 is
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_rst_addr_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_output_valid_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_buf_we_net : std_logic_vector( 1-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal buf_r_data_out_net : std_logic_vector( 36-1 downto 0 );
begin
  output_r <= mux_y_net_x0;
  output_i <= mux1_y_net_x0;
  output_valid <= delay2_q_net;
  mux1_y_net <= input_r;
  mux_y_net <= input_i;
  logical_y_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => mcode_output_valid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_66bf1a97d1
  port map (
    clr => '0',
    start => logical_y_net,
    addr_eq_511 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    buf_we => mcode_buf_we_net,
    output_valid => mcode_output_valid_net,
    rst_addr => mcode_rst_addr_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub1_s_net,
    y => mux1_y_net_x0
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux1_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret3_output_port_net
  );
  relational : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => constant_op_net,
    b => addr_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice1_y_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => mcode_rst_addr_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  buf_r : entity xil_defaultlib.pilotdetect_xlspram
  generic map (
    c_address_width => 9,
    c_width => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i7",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_op_net,
    data_in => concat_y_net,
    we => mcode_buf_we_net,
    clk => clk_net,
    ce => ce_net,
    data_out => buf_r_data_out_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_overlap_and_add4 is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_overlap_and_add4;
architecture structural of pilotdetect_overlap_and_add4 is
  signal clk_net : std_logic;
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
begin
  output <= addsub_s_net;
  output_valid <= delay_q_net;
  logical_y_net <= start;
  mux1_y_net_x0 <= input_r;
  mux_y_net_x0 <= input_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  section_adder : entity xil_defaultlib.pilotdetect_section_adder_x3
  port map (
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    start => logical_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output_r => mux_y_net,
    output_i => mux1_y_net,
    output_valid => delay2_q_net
  );
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 17,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 17,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 2,
    overflow => 2,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 17,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux_y_net,
    b => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux1_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add5/section_adder
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_section_adder_x4 is
  port (
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    start : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output_r : out std_logic_vector( 18-1 downto 0 );
    output_i : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_section_adder_x4;
architecture structural of pilotdetect_section_adder_x4 is
  signal reinterpret1_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret3_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal reinterpret2_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal concat_y_net : std_logic_vector( 36-1 downto 0 );
  signal reinterpret_output_port_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_rst_addr_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_buf_we_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_output_valid_net : std_logic_vector( 1-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 18-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal slice1_y_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net : std_logic_vector( 9-1 downto 0 );
  signal slice_y_net : std_logic_vector( 18-1 downto 0 );
  signal buf_r_data_out_net : std_logic_vector( 36-1 downto 0 );
begin
  output_r <= mux_y_net_x0;
  output_i <= mux1_y_net_x0;
  output_valid <= delay2_q_net;
  mux1_y_net <= input_r;
  mux_y_net <= input_i;
  logical1_y_net <= start;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay_q_net,
    b => reinterpret2_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 1,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay1_q_net,
    b => reinterpret3_output_port_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  concat : entity xil_defaultlib.sysgen_concat_df52b3f9f9
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    in0 => reinterpret_output_port_net,
    in1 => reinterpret1_output_port_net,
    y => concat_y_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => mcode_output_valid_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_66bf1a97d1
  port map (
    clr => '0',
    start => logical1_y_net,
    addr_eq_511 => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    buf_we => mcode_buf_we_net,
    output_valid => mcode_output_valid_net,
    rst_addr => mcode_rst_addr_net
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub_s_net,
    y => mux_y_net_x0
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay2_q_net,
    d0 => constant1_op_net,
    d1 => addsub1_s_net,
    y => mux1_y_net_x0
  );
  reinterpret : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux1_y_net,
    output_port => reinterpret_output_port_net
  );
  reinterpret1 : entity xil_defaultlib.sysgen_reinterpret_70f34f62d7
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => mux_y_net,
    output_port => reinterpret1_output_port_net
  );
  reinterpret2 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice_y_net,
    output_port => reinterpret2_output_port_net
  );
  reinterpret3 : entity xil_defaultlib.sysgen_reinterpret_17fd93603d
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    input_port => slice1_y_net,
    output_port => reinterpret3_output_port_net
  );
  relational : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => constant_op_net,
    b => addr_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
  slice : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 18,
    new_msb => 35,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice_y_net
  );
  slice1 : entity xil_defaultlib.pilotdetect_xlslice
  generic map (
    new_lsb => 0,
    new_msb => 17,
    x_width => 36,
    y_width => 18
  )
  port map (
    x => buf_r_data_out_net,
    y => slice1_y_net
  );
  addr : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => mcode_rst_addr_net,
    clk => clk_net,
    ce => ce_net,
    op => addr_op_net
  );
  buf_r : entity xil_defaultlib.pilotdetect_xlspram
  generic map (
    c_address_width => 9,
    c_width => 36,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i7",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => addr_op_net,
    data_in => concat_y_net,
    we => mcode_buf_we_net,
    clk => clk_net,
    ce => ce_net,
    data_out => buf_r_data_out_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Overlap_and_add5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_overlap_and_add5 is
  port (
    start : in std_logic_vector( 1-1 downto 0 );
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_overlap_and_add5;
architecture structural of pilotdetect_overlap_and_add5 is
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
begin
  output <= addsub_s_net;
  output_valid <= delay_q_net;
  logical1_y_net <= start;
  mux1_y_net_x0 <= input_r;
  mux_y_net_x0 <= input_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  section_adder : entity xil_defaultlib.pilotdetect_section_adder_x4
  port map (
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    start => logical1_y_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output_r => mux_y_net,
    output_i => mux1_y_net,
    output_valid => delay2_q_net
  );
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 17,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 17,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 1,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 2,
    overflow => 2,
    quantization => 1,
    s_arith => xlUnsigned,
    s_bin_pt => 17,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 5,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux_y_net,
    b => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i1",
    extra_registers => 1,
    multsign => 2,
    overflow => 2,
    p_arith => xlSigned,
    p_bin_pt => 17,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => mux1_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Template_center
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_template_center is
  port (
    addr : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    h0_r : out std_logic_vector( 18-1 downto 0 );
    h0_i : out std_logic_vector( 18-1 downto 0 );
    h1_r : out std_logic_vector( 18-1 downto 0 );
    h1_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_template_center;
architecture structural of pilotdetect_template_center is
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal p1_i1_data_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal p0_r1_data_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal p0_i1_data_net : std_logic_vector( 18-1 downto 0 );
  signal p1_r1_data_net : std_logic_vector( 18-1 downto 0 );
begin
  h0_r <= delay3_q_net;
  h0_i <= delay8_q_net;
  h1_r <= delay9_q_net;
  h1_i <= delay10_q_net;
  mcode_a_br_net <= addr;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay10 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p1_i1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p0_r1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p0_i1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p1_r1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  p0_i1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i8",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p0_i1_data_net
  );
  p0_r1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i9",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p0_r1_data_net
  );
  p1_i1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i10",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p1_i1_data_net
  );
  p1_r1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i11",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p1_r1_data_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Template_neg
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_template_neg is
  port (
    addr : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    h0_r : out std_logic_vector( 18-1 downto 0 );
    h0_i : out std_logic_vector( 18-1 downto 0 );
    h1_r : out std_logic_vector( 18-1 downto 0 );
    h1_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_template_neg;
architecture structural of pilotdetect_template_neg is
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal p1_r1_data_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal p0_i1_data_net : std_logic_vector( 18-1 downto 0 );
  signal p0_r1_data_net : std_logic_vector( 18-1 downto 0 );
  signal p1_i1_data_net : std_logic_vector( 18-1 downto 0 );
begin
  h0_r <= delay3_q_net;
  h0_i <= delay8_q_net;
  h1_r <= delay9_q_net;
  h1_i <= delay10_q_net;
  mcode_a_br_net <= addr;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay10 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p1_i1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p0_r1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p0_i1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p1_r1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  p0_i1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i12",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p0_i1_data_net
  );
  p0_r1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i13",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p0_r1_data_net
  );
  p1_i1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i14",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p1_i1_data_net
  );
  p1_r1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i15",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p1_r1_data_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/Template_pos
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_template_pos is
  port (
    addr : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    h0_r : out std_logic_vector( 18-1 downto 0 );
    h0_i : out std_logic_vector( 18-1 downto 0 );
    h1_r : out std_logic_vector( 18-1 downto 0 );
    h1_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_template_pos;
architecture structural of pilotdetect_template_pos is
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal p0_i1_data_net : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal p1_i1_data_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal p0_r1_data_net : std_logic_vector( 18-1 downto 0 );
  signal p1_r1_data_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
begin
  h0_r <= delay3_q_net;
  h0_i <= delay8_q_net;
  h1_r <= delay9_q_net;
  h1_i <= delay10_q_net;
  mcode_a_br_net <= addr;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay10 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p1_i1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay10_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p0_r1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay8 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p0_i1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay8_q_net
  );
  delay9 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => p1_r1_data_net,
    clk => clk_net,
    ce => ce_net,
    q => delay9_q_net
  );
  p0_i1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i16",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p0_i1_data_net
  );
  p0_r1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i17",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p0_r1_data_net
  );
  p1_i1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i18",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p1_i1_data_net
  );
  p1_r1 : entity xil_defaultlib.pilotdetect_xlsprom
  generic map (
    c_address_width => 10,
    c_width => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i19",
    latency => 1
  )
  port map (
    en => "1",
    rst => "0",
    addr => mcode_a_br_net,
    clk => clk_net,
    ce => ce_net,
    data => p1_r1_data_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/complex_mult1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult1 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult1;
architecture structural of pilotdetect_complex_mult1 is
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux2_y_net <= a_r;
  mux3_y_net <= a_i;
  delay3_q_net <= b_r;
  delay1_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux2_y_net,
    b => mux3_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux2_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux3_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net_x0
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net_x0,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/complex_mult2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult2_x0 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult2_x0;
architecture structural of pilotdetect_complex_mult2_x0 is
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux4_y_net <= a_r;
  mux5_y_net <= a_i;
  delay3_q_net <= b_r;
  delay1_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux4_y_net,
    b => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux4_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux5_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net_x0
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net_x0,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/complex_mult3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_complex_mult3_x0 is
  port (
    a_r : in std_logic_vector( 18-1 downto 0 );
    a_i : in std_logic_vector( 18-1 downto 0 );
    b_r : in std_logic_vector( 18-1 downto 0 );
    b_i : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    x_r : out std_logic_vector( 18-1 downto 0 );
    x_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_complex_mult3_x0;
architecture structural of pilotdetect_complex_mult3_x0 is
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult2_p_net : std_logic_vector( 18-1 downto 0 );
  signal mult1_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub3_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub1_s_net : std_logic_vector( 18-1 downto 0 );
  signal addsub2_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal addsub4_s_net : std_logic_vector( 18-1 downto 0 );
  signal mult_p_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
begin
  x_r <= delay4_q_net;
  x_i <= delay5_q_net;
  mux_y_net <= a_r;
  mux1_y_net <= a_i;
  delay3_q_net <= b_r;
  delay1_q_net <= b_i;
  clk_net <= clk_1;
  ce_net <= ce_1;
  addsub : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mux_y_net,
    b => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub_s_net
  );
  addsub1 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i0",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub1_s_net
  );
  addsub2 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => delay3_q_net,
    b => delay1_q_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub2_s_net
  );
  addsub3 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult1_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub3_s_net
  );
  addsub4 : entity xil_defaultlib.pilotdetect_xladdsub
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_has_c_out => 0,
    c_latency => 1,
    c_output_width => 19,
    core_name0 => "pilotdetect_c_addsub_v12_0_i1",
    extra_registers => 0,
    full_s_arith => 2,
    full_s_width => 19,
    latency => 1,
    overflow => 3,
    quantization => 1,
    s_arith => xlSigned,
    s_bin_pt => 16,
    s_width => 18
  )
  port map (
    clr => '0',
    en => "1",
    a => mult2_p_net,
    b => mult_p_net,
    clk => clk_net,
    ce => ce_net,
    s => addsub4_s_net
  );
  delay : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mux1_y_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net_x0
  );
  delay2 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay4 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub3_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => addsub4_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  mult : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay_q_net,
    b => addsub2_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult_p_net
  );
  mult1 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => delay1_q_net_x0,
    b => addsub1_s_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult1_p_net
  );
  mult2 : entity xil_defaultlib.pilotdetect_xlmult
  generic map (
    a_arith => xlSigned,
    a_bin_pt => 16,
    a_width => 18,
    b_arith => xlSigned,
    b_bin_pt => 16,
    b_width => 18,
    c_a_type => 0,
    c_a_width => 18,
    c_b_type => 0,
    c_b_width => 18,
    c_baat => 18,
    c_output_width => 36,
    c_type => 0,
    core_name0 => "pilotdetect_mult_gen_v12_0_i0",
    extra_registers => 0,
    multsign => 2,
    overflow => 3,
    p_arith => xlSigned,
    p_bin_pt => 16,
    p_width => 18,
    quantization => 1
  )
  port map (
    clr => '0',
    core_clr => '1',
    en => "1",
    rst => "0",
    a => addsub_s_net,
    b => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    core_clk => clk_net,
    core_ce => ce_net,
    p => mult2_p_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/fft_buf
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_fft_buf is
  port (
    input_r : in std_logic_vector( 18-1 downto 0 );
    input_i : in std_logic_vector( 18-1 downto 0 );
    w_addr : in std_logic_vector( 10-1 downto 0 );
    we : in std_logic_vector( 1-1 downto 0 );
    r_addr : in std_logic_vector( 10-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    output_r : out std_logic_vector( 18-1 downto 0 );
    output_i : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_fft_buf;
architecture structural of pilotdetect_fft_buf is
  signal ram_i_douta_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal addr_op_net : std_logic_vector( 10-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant1_op_net : std_logic_vector( 18-1 downto 0 );
  signal ram_r_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net_x0 : std_logic_vector( 10-1 downto 0 );
  signal ram_i_doutb_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal write_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal ram_r_douta_net : std_logic_vector( 18-1 downto 0 );
begin
  output_r <= delay3_q_net;
  output_i <= delay1_q_net;
  mux_y_net <= input_r;
  mux1_y_net <= input_i;
  addr_op_net_x0 <= w_addr;
  write_reg_q_net <= we;
  addr_op_net <= r_addr;
  clk_net <= clk_1;
  ce_net <= ce_1;
  constant_x0 : entity xil_defaultlib.sysgen_constant_f456e3a573
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  constant1 : entity xil_defaultlib.sysgen_constant_e3fda8f884
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant1_op_net
  );
  delay1 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => ram_i_doutb_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => ram_r_doutb_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  ram_i : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 10,
    c_address_width_b => 10,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i20",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => addr_op_net_x0,
    dina => mux1_y_net,
    wea => write_reg_q_net,
    addrb => addr_op_net,
    dinb => constant1_op_net,
    web => constant_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => ram_i_douta_net,
    doutb => ram_i_doutb_net
  );
  ram_r : entity xil_defaultlib.pilotdetect_xldpram
  generic map (
    c_address_width_a => 10,
    c_address_width_b => 10,
    c_width_a => 18,
    c_width_b => 18,
    core_name0 => "pilotdetect_blk_mem_gen_v8_3_i20",
    latency => 1
  )
  port map (
    ena => "1",
    enb => "1",
    rsta => "0",
    rstb => "0",
    addra => addr_op_net_x0,
    dina => mux_y_net,
    wea => write_reg_q_net,
    addrb => addr_op_net,
    dinb => constant1_op_net,
    web => constant_op_net,
    a_clk => clk_net,
    a_ce => ce_net,
    b_clk => clk_net,
    b_ce => ce_net,
    douta => ram_r_douta_net,
    doutb => ram_r_doutb_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max/store_max_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_store_max_control is
  port (
    cnt_eq_511 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    cnt_rst : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_store_max_control;
architecture structural of pilotdetect_store_max_control is
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal compare_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
begin
  cnt_rst <= wait_reg_q_net;
  relational2_op_net <= cnt_eq_511;
  delay_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  expression : entity xil_defaultlib.sysgen_expr_fb2a2194e2
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_18ba54a1e8
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression1_dout_net
  );
  compare_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => compare_reg_q_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_find_and_store_max is
  port (
    r0 : in std_logic_vector( 18-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_find_and_store_max;
architecture structural of pilotdetect_find_and_store_max is
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal max_ind_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal max_val_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
begin
  max_ind <= max_ind_reg_0_q_net;
  max_val <= max_val_reg_0_q_net;
  addsub_s_net <= r0;
  delay_q_net <= input_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  store_max_control : entity xil_defaultlib.pilotdetect_store_max_control
  port map (
    cnt_eq_511 => relational2_op_net,
    valid => delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    cnt_rst => wait_reg_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => wait_reg_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => relational2_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  relational : entity xil_defaultlib.sysgen_relational_cb632989dd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => delay2_q_net,
    b => max_val_0_q_net,
    op => relational_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  max_ind_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    d => counter_op_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_0_q_net
  );
  max_ind_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    rst => "0",
    d => max_ind_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_reg_0_q_net
  );
  max_val_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    d => delay2_q_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_0_q_net
  );
  max_val_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    rst => "0",
    d => max_val_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_reg_0_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max1/store_max_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_store_max_control_x0 is
  port (
    cnt_eq_511 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    cnt_rst : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_store_max_control_x0;
architecture structural of pilotdetect_store_max_control_x0 is
  signal clk_net : std_logic;
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal compare_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
begin
  cnt_rst <= wait_reg_q_net;
  relational2_op_net <= cnt_eq_511;
  delay_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  expression : entity xil_defaultlib.sysgen_expr_fb2a2194e2
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_18ba54a1e8
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression1_dout_net
  );
  compare_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => compare_reg_q_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_find_and_store_max1 is
  port (
    r0 : in std_logic_vector( 18-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_find_and_store_max1;
architecture structural of pilotdetect_find_and_store_max1 is
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal max_ind_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal max_val_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  max_ind <= max_ind_reg_0_q_net;
  max_val <= max_val_reg_0_q_net;
  addsub_s_net <= r0;
  delay_q_net <= input_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  store_max_control : entity xil_defaultlib.pilotdetect_store_max_control_x0
  port map (
    cnt_eq_511 => relational2_op_net,
    valid => delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    cnt_rst => wait_reg_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => wait_reg_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => relational2_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  relational : entity xil_defaultlib.sysgen_relational_cb632989dd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => delay2_q_net,
    b => max_val_0_q_net,
    op => relational_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  max_ind_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    d => counter_op_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_0_q_net
  );
  max_ind_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    rst => "0",
    d => max_ind_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_reg_0_q_net
  );
  max_val_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    d => delay2_q_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_0_q_net
  );
  max_val_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    rst => "0",
    d => max_val_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_reg_0_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max2/store_max_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_store_max_control_x1 is
  port (
    cnt_eq_511 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    cnt_rst : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_store_max_control_x1;
architecture structural of pilotdetect_store_max_control_x1 is
  signal ce_net : std_logic;
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal compare_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
begin
  cnt_rst <= wait_reg_q_net;
  relational2_op_net <= cnt_eq_511;
  delay_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  expression : entity xil_defaultlib.sysgen_expr_fb2a2194e2
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_18ba54a1e8
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression1_dout_net
  );
  compare_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => compare_reg_q_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_find_and_store_max2 is
  port (
    r0 : in std_logic_vector( 18-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_find_and_store_max2;
architecture structural of pilotdetect_find_and_store_max2 is
  signal clk_net : std_logic;
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal max_val_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal counter_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal max_ind_0_q_net : std_logic_vector( 9-1 downto 0 );
begin
  max_ind <= max_ind_reg_0_q_net;
  max_val <= max_val_reg_0_q_net;
  addsub_s_net <= r0;
  delay_q_net <= input_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  store_max_control : entity xil_defaultlib.pilotdetect_store_max_control_x1
  port map (
    cnt_eq_511 => relational2_op_net,
    valid => delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    cnt_rst => wait_reg_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => wait_reg_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => relational2_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  relational : entity xil_defaultlib.sysgen_relational_cb632989dd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => delay2_q_net,
    b => max_val_0_q_net,
    op => relational_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  max_ind_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    d => counter_op_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_0_q_net
  );
  max_ind_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    rst => "0",
    d => max_ind_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_reg_0_q_net
  );
  max_val_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    d => delay2_q_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_0_q_net
  );
  max_val_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    rst => "0",
    d => max_val_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_reg_0_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max3/store_max_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_store_max_control_x2 is
  port (
    cnt_eq_511 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    cnt_rst : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_store_max_control_x2;
architecture structural of pilotdetect_store_max_control_x2 is
  signal clk_net : std_logic;
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal compare_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
begin
  cnt_rst <= wait_reg_q_net;
  relational2_op_net <= cnt_eq_511;
  delay_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  expression : entity xil_defaultlib.sysgen_expr_fb2a2194e2
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_18ba54a1e8
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression1_dout_net
  );
  compare_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => compare_reg_q_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_find_and_store_max3 is
  port (
    r0 : in std_logic_vector( 18-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_find_and_store_max3;
architecture structural of pilotdetect_find_and_store_max3 is
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal max_val_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal max_ind_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal counter_op_net : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
begin
  max_ind <= max_ind_reg_0_q_net;
  max_val <= max_val_reg_0_q_net;
  addsub_s_net <= r0;
  delay_q_net <= input_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  store_max_control : entity xil_defaultlib.pilotdetect_store_max_control_x2
  port map (
    cnt_eq_511 => relational2_op_net,
    valid => delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    cnt_rst => wait_reg_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => wait_reg_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => relational2_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  relational : entity xil_defaultlib.sysgen_relational_cb632989dd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => delay2_q_net,
    b => max_val_0_q_net,
    op => relational_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  max_ind_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    d => counter_op_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_0_q_net
  );
  max_ind_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    rst => "0",
    d => max_ind_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_reg_0_q_net
  );
  max_val_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    d => delay2_q_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_0_q_net
  );
  max_val_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    rst => "0",
    d => max_val_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_reg_0_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max4/store_max_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_store_max_control_x3 is
  port (
    cnt_eq_511 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    cnt_rst : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_store_max_control_x3;
architecture structural of pilotdetect_store_max_control_x3 is
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal compare_reg_q_net : std_logic_vector( 1-1 downto 0 );
begin
  cnt_rst <= wait_reg_q_net;
  relational2_op_net <= cnt_eq_511;
  delay_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  expression : entity xil_defaultlib.sysgen_expr_fb2a2194e2
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_18ba54a1e8
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression1_dout_net
  );
  compare_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => compare_reg_q_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_find_and_store_max4 is
  port (
    r0 : in std_logic_vector( 18-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_find_and_store_max4;
architecture structural of pilotdetect_find_and_store_max4 is
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal counter_op_net : std_logic_vector( 9-1 downto 0 );
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal clk_net : std_logic;
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal max_val_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal max_ind_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  max_ind <= max_ind_reg_0_q_net;
  max_val <= max_val_reg_0_q_net;
  addsub_s_net <= r0;
  delay_q_net <= input_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  store_max_control : entity xil_defaultlib.pilotdetect_store_max_control_x3
  port map (
    cnt_eq_511 => relational2_op_net,
    valid => delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    cnt_rst => wait_reg_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => wait_reg_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => relational2_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  relational : entity xil_defaultlib.sysgen_relational_cb632989dd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => delay2_q_net,
    b => max_val_0_q_net,
    op => relational_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  max_ind_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    d => counter_op_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_0_q_net
  );
  max_ind_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    rst => "0",
    d => max_ind_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_reg_0_q_net
  );
  max_val_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    d => delay2_q_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_0_q_net
  );
  max_val_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    rst => "0",
    d => max_val_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_reg_0_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max5/store_max_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_store_max_control_x4 is
  port (
    cnt_eq_511 : in std_logic_vector( 1-1 downto 0 );
    valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    cnt_rst : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_store_max_control_x4;
architecture structural of pilotdetect_store_max_control_x4 is
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal compare_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal expression_dout_net : std_logic_vector( 1-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
begin
  cnt_rst <= wait_reg_q_net;
  relational2_op_net <= cnt_eq_511;
  delay_q_net <= valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  expression : entity xil_defaultlib.sysgen_expr_fb2a2194e2
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression_dout_net
  );
  expression1 : entity xil_defaultlib.sysgen_expr_18ba54a1e8
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    cnt_eq_511 => relational2_op_net,
    compare => compare_reg_q_net,
    valid => delay_q_net,
    wait_x0 => wait_reg_q_net,
    dout => expression1_dout_net
  );
  compare_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"0"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => compare_reg_q_net
  );
  wait_reg : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 1,
    init_value => b"1"
  )
  port map (
    en => "1",
    rst => "0",
    d => expression_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => wait_reg_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/find_and_store_max5
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_find_and_store_max5 is
  port (
    r0 : in std_logic_vector( 18-1 downto 0 );
    input_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 );
    output_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_find_and_store_max5;
architecture structural of pilotdetect_find_and_store_max5 is
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal ce_net : std_logic;
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal wait_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal counter_op_net : std_logic_vector( 9-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal constant_op_net : std_logic_vector( 9-1 downto 0 );
  signal relational2_op_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal max_val_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal max_ind_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
begin
  max_ind <= max_ind_reg_0_q_net;
  max_val <= max_val_reg_0_q_net;
  output_valid <= delay1_q_net;
  addsub_s_net <= r0;
  delay_q_net <= input_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  store_max_control : entity xil_defaultlib.pilotdetect_store_max_control_x4
  port map (
    cnt_eq_511 => relational2_op_net,
    valid => delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    cnt_rst => wait_reg_q_net
  );
  constant_x0 : entity xil_defaultlib.sysgen_constant_0e16603724
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    op => constant_op_net
  );
  counter : entity xil_defaultlib.pilotdetect_xlcounter_free
  generic map (
    core_name0 => "pilotdetect_c_counter_binary_v12_0_i0",
    op_arith => xlUnsigned,
    op_width => 9
  )
  port map (
    en => "1",
    clr => '0',
    rst => wait_reg_q_net,
    clk => clk_net,
    ce => ce_net,
    op => counter_op_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => addsub_s_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => relational2_op_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  relational : entity xil_defaultlib.sysgen_relational_cb632989dd
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => delay2_q_net,
    b => max_val_0_q_net,
    op => relational_op_net
  );
  relational2 : entity xil_defaultlib.sysgen_relational_1b89fab8d7
  port map (
    clr => '0',
    a => counter_op_net,
    b => constant_op_net,
    clk => clk_net,
    ce => ce_net,
    op => relational2_op_net
  );
  max_ind_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    d => counter_op_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_0_q_net
  );
  max_ind_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 9,
    init_value => b"000000000"
  )
  port map (
    rst => "0",
    d => max_ind_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_ind_reg_0_q_net
  );
  max_val_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    d => delay2_q_net,
    rst => wait_reg_q_net,
    en => relational_op_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_0_q_net
  );
  max_val_reg_0 : entity xil_defaultlib.pilotdetect_xlregister
  generic map (
    d_width => 18,
    init_value => b"000000000000000000"
  )
  port map (
    rst => "0",
    d => max_val_0_q_net,
    en => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => max_val_reg_0_q_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/pass_max
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_pass_max is
  port (
    max_ind_a : in std_logic_vector( 9-1 downto 0 );
    max_val_a : in std_logic_vector( 18-1 downto 0 );
    max_ind_b : in std_logic_vector( 9-1 downto 0 );
    max_val_b : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_pass_max;
architecture structural of pilotdetect_pass_max is
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal max_val_reg_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal clk_net : std_logic;
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
begin
  max_ind <= mux7_y_net;
  max_val <= mux6_y_net;
  max_ind_reg_0_q_net <= max_ind_a;
  max_val_reg_0_q_net_x0 <= max_val_a;
  max_ind_reg_0_q_net_x0 <= max_ind_b;
  max_val_reg_0_q_net <= max_val_b;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => max_val_reg_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => max_val_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => max_ind_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => max_ind_reg_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay3_q_net,
    d1 => delay4_q_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_92b6e25f44
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay5_q_net,
    d1 => delay6_q_net,
    y => mux7_y_net
  );
  relational : entity xil_defaultlib.sysgen_relational_45adaa63b5
  port map (
    clr => '0',
    a => max_val_reg_0_q_net_x0,
    b => max_val_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/pass_max1
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_pass_max1 is
  port (
    max_ind_a : in std_logic_vector( 9-1 downto 0 );
    max_val_a : in std_logic_vector( 18-1 downto 0 );
    max_ind_b : in std_logic_vector( 9-1 downto 0 );
    max_val_b : in std_logic_vector( 18-1 downto 0 );
    in_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 );
    out_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_pass_max1;
architecture structural of pilotdetect_pass_max1 is
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal max_val_reg_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal ce_net : std_logic;
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
begin
  max_ind <= mux7_y_net;
  max_val <= mux6_y_net;
  out_valid <= delay1_q_net;
  max_ind_reg_0_q_net <= max_ind_a;
  max_val_reg_0_q_net_x0 <= max_val_a;
  max_ind_reg_0_q_net_x0 <= max_ind_b;
  max_val_reg_0_q_net <= max_val_b;
  delay1_q_net_x0 <= in_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay1_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => max_val_reg_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => max_val_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => max_ind_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => max_ind_reg_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay3_q_net,
    d1 => delay4_q_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_92b6e25f44
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay5_q_net,
    d1 => delay6_q_net,
    y => mux7_y_net
  );
  relational : entity xil_defaultlib.sysgen_relational_45adaa63b5
  port map (
    clr => '0',
    a => max_val_reg_0_q_net_x0,
    b => max_val_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/pass_max2
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_pass_max2 is
  port (
    max_ind_a : in std_logic_vector( 9-1 downto 0 );
    max_val_a : in std_logic_vector( 18-1 downto 0 );
    max_ind_b : in std_logic_vector( 9-1 downto 0 );
    max_val_b : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_pass_max2;
architecture structural of pilotdetect_pass_max2 is
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal max_ind_reg_0_q_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal clk_net : std_logic;
  signal max_val_reg_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
begin
  max_ind <= mux7_y_net;
  max_val <= mux6_y_net;
  max_ind_reg_0_q_net <= max_ind_a;
  max_val_reg_0_q_net_x0 <= max_val_a;
  max_ind_reg_0_q_net_x0 <= max_ind_b;
  max_val_reg_0_q_net <= max_val_b;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => max_val_reg_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => max_val_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => max_ind_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => max_ind_reg_0_q_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay3_q_net,
    d1 => delay4_q_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_92b6e25f44
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay5_q_net,
    d1 => delay6_q_net,
    y => mux7_y_net
  );
  relational : entity xil_defaultlib.sysgen_relational_45adaa63b5
  port map (
    clr => '0',
    a => max_val_reg_0_q_net_x0,
    b => max_val_reg_0_q_net,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/pass_max3
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_pass_max3 is
  port (
    max_ind_a : in std_logic_vector( 9-1 downto 0 );
    max_val_a : in std_logic_vector( 18-1 downto 0 );
    max_ind_b : in std_logic_vector( 9-1 downto 0 );
    max_val_b : in std_logic_vector( 18-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_pass_max3;
architecture structural of pilotdetect_pass_max3 is
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal mux7_y_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal mux7_y_net_x1 : std_logic_vector( 9-1 downto 0 );
  signal ce_net : std_logic;
  signal mux6_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal mux6_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
begin
  max_ind <= mux7_y_net;
  max_val <= mux6_y_net;
  mux7_y_net_x1 <= max_ind_a;
  mux6_y_net_x0 <= max_val_a;
  mux7_y_net_x0 <= max_ind_b;
  mux6_y_net_x1 <= max_val_b;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux6_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux6_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => mux7_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => mux7_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay3_q_net,
    d1 => delay4_q_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_92b6e25f44
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay5_q_net,
    d1 => delay6_q_net,
    y => mux7_y_net
  );
  relational : entity xil_defaultlib.sysgen_relational_45adaa63b5
  port map (
    clr => '0',
    a => mux6_y_net_x0,
    b => mux6_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator/pass_max4
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_pass_max4 is
  port (
    max_ind_a : in std_logic_vector( 9-1 downto 0 );
    max_val_a : in std_logic_vector( 18-1 downto 0 );
    max_ind_b : in std_logic_vector( 9-1 downto 0 );
    max_val_b : in std_logic_vector( 18-1 downto 0 );
    in_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 );
    out_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_pass_max4;
architecture structural of pilotdetect_pass_max4 is
  signal delay5_q_net : std_logic_vector( 9-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal mux7_y_net_x1 : std_logic_vector( 9-1 downto 0 );
  signal delay6_q_net : std_logic_vector( 9-1 downto 0 );
  signal ce_net : std_logic;
  signal clk_net : std_logic;
  signal mux6_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux6_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux7_y_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 1-1 downto 0 );
  signal relational_op_net : std_logic_vector( 1-1 downto 0 );
begin
  max_ind <= mux7_y_net;
  max_val <= mux6_y_net;
  out_valid <= delay1_q_net;
  mux7_y_net_x0 <= max_ind_a;
  mux6_y_net_x0 <= max_val_a;
  mux7_y_net_x1 <= max_ind_b;
  mux6_y_net_x1 <= max_val_b;
  delay3_q_net <= in_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay3_q_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux6_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net_x0
  );
  delay4 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => mux6_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay4_q_net
  );
  delay5 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => mux7_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay5_q_net
  );
  delay6 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    en => '1',
    rst => '1',
    d => mux7_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    q => delay6_q_net
  );
  mux6 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay3_q_net_x0,
    d1 => delay4_q_net,
    y => mux6_y_net
  );
  mux7 : entity xil_defaultlib.sysgen_mux_92b6e25f44
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => relational_op_net,
    d0 => delay5_q_net,
    d1 => delay6_q_net,
    y => mux7_y_net
  );
  relational : entity xil_defaultlib.sysgen_relational_45adaa63b5
  port map (
    clr => '0',
    a => mux6_y_net_x0,
    b => mux6_y_net_x1,
    clk => clk_net,
    ce => ce_net,
    op => relational_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/multi_band_correlator
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_multi_band_correlator is
  port (
    in_real : in std_logic_vector( 18-1 downto 0 );
    in_imag : in std_logic_vector( 18-1 downto 0 );
    start_input : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    max_ind : out std_logic_vector( 9-1 downto 0 );
    max_val : out std_logic_vector( 18-1 downto 0 );
    out_valid : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_multi_band_correlator;
architecture structural of pilotdetect_multi_band_correlator is
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal clk_net : std_logic;
  signal delay2_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay6_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay5_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net_x0 : std_logic_vector( 10-1 downto 0 );
  signal mux1_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux1_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay4_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal addr_op_net : std_logic_vector( 10-1 downto 0 );
  signal mcode_a_br_net : std_logic_vector( 10-1 downto 0 );
  signal logical1_y_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay4_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay5_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal write_reg_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal expression1_dout_net : std_logic_vector( 1-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal logical1_y_net : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net_x4 : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal mux6_y_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal delay9_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux4_y_net : std_logic_vector( 18-1 downto 0 );
  signal max_val_reg_0_q_net_x4 : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net_x2 : std_logic_vector( 9-1 downto 0 );
  signal max_val_reg_0_q_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal max_val_reg_0_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal mux5_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal delay8_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net : std_logic_vector( 9-1 downto 0 );
  signal mux7_y_net_x3 : std_logic_vector( 9-1 downto 0 );
  signal mux7_y_net_x2 : std_logic_vector( 9-1 downto 0 );
  signal mux6_y_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal max_val_reg_0_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x3 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal addsub_s_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal mux7_y_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal delay9_q_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net_x1 : std_logic_vector( 9-1 downto 0 );
  signal max_ind_reg_0_q_net_x4 : std_logic_vector( 9-1 downto 0 );
  signal addsub_s_net_x1 : std_logic_vector( 18-1 downto 0 );
  signal addsub_s_net : std_logic_vector( 18-1 downto 0 );
  signal max_val_reg_0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux3_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net_x3 : std_logic_vector( 18-1 downto 0 );
  signal max_val_reg_0_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x5 : std_logic_vector( 1-1 downto 0 );
  signal max_ind_reg_0_q_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal mux7_y_net_x1 : std_logic_vector( 9-1 downto 0 );
  signal delay9_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal delay10_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x11 : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay8_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay3_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal mux6_y_net_x2 : std_logic_vector( 18-1 downto 0 );
  signal max_ind_reg_0_q_net_x3 : std_logic_vector( 9-1 downto 0 );
  signal delay_q_net : std_logic_vector( 1-1 downto 0 );
  signal mux6_y_net_x1 : std_logic_vector( 18-1 downto 0 );
begin
  max_ind <= mux7_y_net;
  max_val <= mux6_y_net;
  out_valid <= delay1_q_net_x1;
  mux_y_net_x4 <= in_real;
  mux2_y_net_x0 <= in_imag;
  delay0_q_net <= start_input;
  clk_net <= clk_1;
  ce_net <= ce_1;
  fft_1024 : entity xil_defaultlib.pilotdetect_fft_1024
  port map (
    x_r_x0 => mux_y_net_x4,
    x_i => mux2_y_net_x0,
    start => delay0_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => mux_y_net_x3,
    x_i_x0 => mux1_y_net_x3,
    done => delay6_q_net_x2
  );
  fft_buf_control : entity xil_defaultlib.pilotdetect_fft_buf_control
  port map (
    start => delay6_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    write => write_reg_q_net,
    write_addr => addr_op_net_x0
  );
  ifft_1024_ver_1 : entity xil_defaultlib.pilotdetect_ifft_1024_ver_1
  port map (
    x_r_x0 => delay4_q_net,
    x_i_x0 => delay5_q_net,
    start => delay2_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => mux1_y_net_x2,
    x_i => mux_y_net_x2
  );
  ifft_1024_ver_2 : entity xil_defaultlib.pilotdetect_ifft_1024_ver_2
  port map (
    x_r_x0 => delay4_q_net_x0,
    x_i_x0 => delay5_q_net_x0,
    start => delay2_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => mux1_y_net_x1,
    x_i => mux_y_net_x1,
    done => delay6_q_net_x0
  );
  ifft_1024_ver_3 : entity xil_defaultlib.pilotdetect_ifft_1024_ver_3
  port map (
    x_r_x0 => delay4_q_net_x1,
    x_i_x0 => delay5_q_net_x1,
    start => delay2_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => mux1_y_net_x0,
    x_i => mux_y_net_x0
  );
  ifft_input_control : entity xil_defaultlib.pilotdetect_ifft_input_control
  port map (
    start => delay_q_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    read_addr => addr_op_net,
    read_addr_reversed => mcode_a_br_net,
    h_sel => logical1_y_net_x0,
    ifft_start => expression1_dout_net
  );
  ona_input_control : entity xil_defaultlib.pilotdetect_ona_input_control
  port map (
    s => delay6_q_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    r0 => logical_y_net,
    r1 => logical1_y_net
  );
  overlap_and_add : entity xil_defaultlib.pilotdetect_overlap_and_add
  port map (
    start => logical_y_net,
    input_r => mux1_y_net_x1,
    input_i => mux_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => addsub_s_net_x4,
    output_valid => delay_q_net_x4
  );
  overlap_and_add1 : entity xil_defaultlib.pilotdetect_overlap_and_add1
  port map (
    start => logical1_y_net,
    input_r => mux1_y_net_x1,
    input_i => mux_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => addsub_s_net_x3,
    output_valid => delay_q_net_x3
  );
  overlap_and_add2 : entity xil_defaultlib.pilotdetect_overlap_and_add2
  port map (
    start => logical_y_net,
    input_r => mux1_y_net_x2,
    input_i => mux_y_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => addsub_s_net_x2,
    output_valid => delay_q_net_x2
  );
  overlap_and_add3 : entity xil_defaultlib.pilotdetect_overlap_and_add3
  port map (
    start => logical1_y_net,
    input_r => mux1_y_net_x2,
    input_i => mux_y_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => addsub_s_net_x1,
    output_valid => delay_q_net_x1
  );
  overlap_and_add4 : entity xil_defaultlib.pilotdetect_overlap_and_add4
  port map (
    start => logical_y_net,
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => addsub_s_net_x0,
    output_valid => delay_q_net_x0
  );
  overlap_and_add5 : entity xil_defaultlib.pilotdetect_overlap_and_add5
  port map (
    start => logical1_y_net,
    input_r => mux1_y_net_x0,
    input_i => mux_y_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output => addsub_s_net,
    output_valid => delay_q_net
  );
  template_center : entity xil_defaultlib.pilotdetect_template_center
  port map (
    addr => mcode_a_br_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    h0_r => delay3_q_net_x1,
    h0_i => delay8_q_net_x1,
    h1_r => delay9_q_net_x1,
    h1_i => delay10_q_net_x1
  );
  template_neg : entity xil_defaultlib.pilotdetect_template_neg
  port map (
    addr => mcode_a_br_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    h0_r => delay3_q_net_x0,
    h0_i => delay8_q_net_x0,
    h1_r => delay9_q_net_x0,
    h1_i => delay10_q_net_x0
  );
  template_pos : entity xil_defaultlib.pilotdetect_template_pos
  port map (
    addr => mcode_a_br_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    h0_r => delay3_q_net,
    h0_i => delay8_q_net,
    h1_r => delay9_q_net,
    h1_i => delay10_q_net
  );
  complex_mult1 : entity xil_defaultlib.pilotdetect_complex_mult1
  port map (
    a_r => mux2_y_net,
    a_i => mux3_y_net,
    b_r => delay3_q_net_x3,
    b_i => delay1_q_net_x11,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net,
    x_i => delay5_q_net
  );
  complex_mult2 : entity xil_defaultlib.pilotdetect_complex_mult2_x0
  port map (
    a_r => mux4_y_net,
    a_i => mux5_y_net,
    b_r => delay3_q_net_x3,
    b_i => delay1_q_net_x11,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x1,
    x_i => delay5_q_net_x1
  );
  complex_mult3 : entity xil_defaultlib.pilotdetect_complex_mult3_x0
  port map (
    a_r => mux_y_net,
    a_i => mux1_y_net,
    b_r => delay3_q_net_x3,
    b_i => delay1_q_net_x11,
    clk_1 => clk_net,
    ce_1 => ce_net,
    x_r => delay4_q_net_x0,
    x_i => delay5_q_net_x0
  );
  fft_buf : entity xil_defaultlib.pilotdetect_fft_buf
  port map (
    input_r => mux_y_net_x3,
    input_i => mux1_y_net_x3,
    w_addr => addr_op_net_x0,
    we => write_reg_q_net,
    r_addr => addr_op_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    output_r => delay3_q_net_x3,
    output_i => delay1_q_net_x11
  );
  find_and_store_max : entity xil_defaultlib.pilotdetect_find_and_store_max
  port map (
    r0 => addsub_s_net_x4,
    input_valid => delay_q_net_x4,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => max_ind_reg_0_q_net_x4,
    max_val => max_val_reg_0_q_net_x4
  );
  find_and_store_max1 : entity xil_defaultlib.pilotdetect_find_and_store_max1
  port map (
    r0 => addsub_s_net_x3,
    input_valid => delay_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => max_ind_reg_0_q_net_x3,
    max_val => max_val_reg_0_q_net_x3
  );
  find_and_store_max2 : entity xil_defaultlib.pilotdetect_find_and_store_max2
  port map (
    r0 => addsub_s_net_x2,
    input_valid => delay_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => max_ind_reg_0_q_net_x2,
    max_val => max_val_reg_0_q_net_x2
  );
  find_and_store_max3 : entity xil_defaultlib.pilotdetect_find_and_store_max3
  port map (
    r0 => addsub_s_net_x1,
    input_valid => delay_q_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => max_ind_reg_0_q_net_x1,
    max_val => max_val_reg_0_q_net_x1
  );
  find_and_store_max4 : entity xil_defaultlib.pilotdetect_find_and_store_max4
  port map (
    r0 => addsub_s_net_x0,
    input_valid => delay_q_net_x0,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => max_ind_reg_0_q_net_x0,
    max_val => max_val_reg_0_q_net_x0
  );
  find_and_store_max5 : entity xil_defaultlib.pilotdetect_find_and_store_max5
  port map (
    r0 => addsub_s_net,
    input_valid => delay_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => max_ind_reg_0_q_net,
    max_val => max_val_reg_0_q_net,
    output_valid => delay1_q_net_x5
  );
  pass_max : entity xil_defaultlib.pilotdetect_pass_max
  port map (
    max_ind_a => max_ind_reg_0_q_net_x4,
    max_val_a => max_val_reg_0_q_net_x4,
    max_ind_b => max_ind_reg_0_q_net_x3,
    max_val_b => max_val_reg_0_q_net_x3,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => mux7_y_net_x3,
    max_val => mux6_y_net_x3
  );
  pass_max1 : entity xil_defaultlib.pilotdetect_pass_max1
  port map (
    max_ind_a => max_ind_reg_0_q_net_x0,
    max_val_a => max_val_reg_0_q_net_x0,
    max_ind_b => max_ind_reg_0_q_net,
    max_val_b => max_val_reg_0_q_net,
    in_valid => delay1_q_net_x5,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => mux7_y_net_x2,
    max_val => mux6_y_net_x2,
    out_valid => delay1_q_net_x3
  );
  pass_max2 : entity xil_defaultlib.pilotdetect_pass_max2
  port map (
    max_ind_a => max_ind_reg_0_q_net_x2,
    max_val_a => max_val_reg_0_q_net_x2,
    max_ind_b => max_ind_reg_0_q_net_x1,
    max_val_b => max_val_reg_0_q_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => mux7_y_net_x1,
    max_val => mux6_y_net_x1
  );
  pass_max3 : entity xil_defaultlib.pilotdetect_pass_max3
  port map (
    max_ind_a => mux7_y_net_x3,
    max_val_a => mux6_y_net_x3,
    max_ind_b => mux7_y_net_x1,
    max_val_b => mux6_y_net_x1,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => mux7_y_net_x0,
    max_val => mux6_y_net_x0
  );
  pass_max4 : entity xil_defaultlib.pilotdetect_pass_max4
  port map (
    max_ind_a => mux7_y_net_x0,
    max_val_a => mux6_y_net_x0,
    max_ind_b => mux7_y_net_x2,
    max_val_b => mux6_y_net_x2,
    in_valid => delay3_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => mux7_y_net,
    max_val => mux6_y_net,
    out_valid => delay1_q_net_x1
  );
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay6_q_net_x2,
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net_x5
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 2,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => logical1_y_net_x0,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net_x0
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 9,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => expression1_dout_net,
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => delay1_q_net_x3,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net_x2
  );
  mux : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay1_q_net_x0,
    d0 => delay3_q_net_x0,
    d1 => delay9_q_net_x0,
    y => mux_y_net
  );
  mux1 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay1_q_net_x0,
    d0 => delay8_q_net_x0,
    d1 => delay10_q_net_x0,
    y => mux1_y_net
  );
  mux2 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay1_q_net_x0,
    d0 => delay3_q_net_x1,
    d1 => delay9_q_net_x1,
    y => mux2_y_net
  );
  mux3 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay1_q_net_x0,
    d0 => delay8_q_net_x1,
    d1 => delay10_q_net_x1,
    y => mux3_y_net
  );
  mux4 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay1_q_net_x0,
    d0 => delay3_q_net,
    d1 => delay9_q_net,
    y => mux4_y_net
  );
  mux5 : entity xil_defaultlib.sysgen_mux_6d354cfe17
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    sel => delay1_q_net_x0,
    d0 => delay8_q_net,
    d1 => delay10_q_net,
    y => mux5_y_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect/pd_control
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_pd_control is
  port (
    max_index : in std_logic_vector( 9-1 downto 0 );
    max_value : in std_logic_vector( 18-1 downto 0 );
    pilot_valid : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    pilot_index : out std_logic_vector( 9-1 downto 0 );
    pilot_found : out std_logic_vector( 1-1 downto 0 );
    pilot_mag : out std_logic_vector( 18-1 downto 0 );
    pilot_pulse : out std_logic_vector( 1-1 downto 0 );
    threshold : out std_logic_vector( 18-1 downto 0 )
  );
end pilotdetect_pd_control;
architecture structural of pilotdetect_pd_control is
  signal delay1_q_net_x0 : std_logic_vector( 1-1 downto 0 );
  signal clk_net : std_logic;
  signal ce_net : std_logic;
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay2_q_net : std_logic_vector( 18-1 downto 0 );
  signal relational1_op_net : std_logic_vector( 1-1 downto 0 );
  signal mcode_threshold_net : std_logic_vector( 18-1 downto 0 );
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 9-1 downto 0 );
  signal mcode_pilotfound_net : std_logic_vector( 1-1 downto 0 );
begin
  pilot_index <= delay1_q_net;
  pilot_found <= mcode_pilotfound_net;
  pilot_mag <= delay_q_net;
  pilot_pulse <= logical_y_net;
  threshold <= delay3_q_net;
  mux7_y_net <= max_index;
  mux6_y_net <= max_value;
  delay1_q_net_x0 <= pilot_valid;
  clk_net <= clk_1;
  ce_net <= ce_1;
  delay : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    rst => '1',
    d => mux6_y_net,
    en => delay1_q_net_x0(0),
    clk => clk_net,
    ce => ce_net,
    q => delay_q_net
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 9
  )
  port map (
    rst => '1',
    d => mux7_y_net,
    en => delay1_q_net_x0(0),
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net
  );
  delay2 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 26,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    rst => '1',
    d => delay_q_net,
    en => delay1_q_net_x0(0),
    clk => clk_net,
    ce => ce_net,
    q => delay2_q_net
  );
  delay3 : entity xil_defaultlib.sysgen_delay_8b3a0008e3
  port map (
    clr => '0',
    d => mcode_threshold_net,
    clk => clk_net,
    ce => ce_net,
    q => delay3_q_net
  );
  logical : entity xil_defaultlib.sysgen_logical_f0792c23bd
  port map (
    clr => '0',
    d0 => relational1_op_net,
    d1 => delay1_q_net_x0,
    d2 => mcode_pilotfound_net,
    clk => clk_net,
    ce => ce_net,
    y => logical_y_net
  );
  mcode : entity xil_defaultlib.sysgen_mcode_block_9f7c19dc49
  port map (
    clr => '0',
    maxvalid_i => relational1_op_net,
    valid_i => delay1_q_net_x0,
    pilotmag => delay_q_net,
    delaymag => delay2_q_net,
    clk => clk_net,
    ce => ce_net,
    pilotfound => mcode_pilotfound_net,
    threshold => mcode_threshold_net
  );
  relational1 : entity xil_defaultlib.sysgen_relational_924fff1a23
  port map (
    clk => '0',
    ce => '0',
    clr => '0',
    a => mux6_y_net,
    b => delay3_q_net,
    op => relational1_op_net
  );
end structural;
-- Generated from Simulink block Brik1/PilotDetect_struct
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_struct is
  port (
    imagdata : in std_logic_vector( 18-1 downto 0 );
    realdata : in std_logic_vector( 18-1 downto 0 );
    validpilot : in std_logic_vector( 1-1 downto 0 );
    conj_imag : in std_logic_vector( 1-1 downto 0 );
    clk_1 : in std_logic;
    ce_1 : in std_logic;
    imagpilotout : out std_logic_vector( 18-1 downto 0 );
    realpilotout : out std_logic_vector( 18-1 downto 0 );
    threshold : out std_logic_vector( 18-1 downto 0 );
    validpilotout : out std_logic_vector( 1-1 downto 0 );
    pilot_found : out std_logic_vector( 1-1 downto 0 );
    pilot_indexes : out std_logic_vector( 9-1 downto 0 );
    pilot_mag : out std_logic_vector( 18-1 downto 0 );
    pilot_pulse : out std_logic_vector( 1-1 downto 0 )
  );
end pilotdetect_struct;
architecture structural of pilotdetect_struct is
  signal imagdata_net : std_logic_vector( 18-1 downto 0 );
  signal mcode_pilotfound_net : std_logic_vector( 1-1 downto 0 );
  signal realdata_net : std_logic_vector( 18-1 downto 0 );
  signal delay0_q_net_x0 : std_logic_vector( 18-1 downto 0 );
  signal clk_net : std_logic;
  signal logical_y_net : std_logic_vector( 1-1 downto 0 );
  signal delay1_q_net_x0 : std_logic_vector( 9-1 downto 0 );
  signal mux1_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x2 : std_logic_vector( 1-1 downto 0 );
  signal delay3_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux2_y_net : std_logic_vector( 18-1 downto 0 );
  signal mux7_y_net : std_logic_vector( 9-1 downto 0 );
  signal delay1_q_net : std_logic_vector( 1-1 downto 0 );
  signal delay_q_net : std_logic_vector( 18-1 downto 0 );
  signal mux6_y_net : std_logic_vector( 18-1 downto 0 );
  signal delay1_q_net_x1 : std_logic_vector( 1-1 downto 0 );
  signal conj_imag_net : std_logic_vector( 1-1 downto 0 );
  signal delay0_q_net : std_logic_vector( 1-1 downto 0 );
  signal negate_op_net : std_logic_vector( 18-1 downto 0 );
  signal mux_y_net : std_logic_vector( 18-1 downto 0 );
  signal ce_net : std_logic;
  signal validpilot_net : std_logic_vector( 1-1 downto 0 );
begin
  imagdata_net <= imagdata;
  imagpilotout <= mux2_y_net;
  realdata_net <= realdata;
  realpilotout <= mux_y_net;
  threshold <= delay3_q_net;
  validpilot_net <= validpilot;
  validpilotout <= delay1_q_net_x1;
  conj_imag_net <= conj_imag;
  pilot_found <= mcode_pilotfound_net;
  pilot_indexes <= delay1_q_net_x0;
  pilot_mag <= delay_q_net;
  pilot_pulse <= logical_y_net;
  clk_net <= clk_1;
  ce_net <= ce_1;
  correlator_fifo : entity xil_defaultlib.pilotdetect_correlator_fifo
  port map (
    real_in => delay0_q_net_x0,
    imag_in => mux1_y_net,
    valid_in => delay1_q_net_x2,
    clk_1 => clk_net,
    ce_1 => ce_net,
    real_out => mux_y_net,
    imag_out => mux2_y_net,
    start_correlator => delay0_q_net,
    valid_out => delay1_q_net_x1
  );
  multi_band_correlator : entity xil_defaultlib.pilotdetect_multi_band_correlator
  port map (
    in_real => mux_y_net,
    in_imag => mux2_y_net,
    start_input => delay0_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    max_ind => mux7_y_net,
    max_val => mux6_y_net,
    out_valid => delay1_q_net
  );
  pd_control : entity xil_defaultlib.pilotdetect_pd_control
  port map (
    max_index => mux7_y_net,
    max_value => mux6_y_net,
    pilot_valid => delay1_q_net,
    clk_1 => clk_net,
    ce_1 => ce_net,
    pilot_index => delay1_q_net_x0,
    pilot_found => mcode_pilotfound_net,
    pilot_mag => delay_q_net,
    pilot_pulse => logical_y_net,
    threshold => delay3_q_net
  );
  delay0 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 18
  )
  port map (
    en => '1',
    rst => '1',
    d => realdata_net,
    clk => clk_net,
    ce => ce_net,
    q => delay0_q_net_x0
  );
  delay1 : entity xil_defaultlib.pilotdetect_xldelay
  generic map (
    latency => 1,
    reg_retiming => 0,
    reset => 0,
    width => 1
  )
  port map (
    en => '1',
    rst => '1',
    d => validpilot_net,
    clk => clk_net,
    ce => ce_net,
    q => delay1_q_net_x2
  );
  mux1 : entity xil_defaultlib.sysgen_mux_148444ce42
  port map (
    clr => '0',
    sel => conj_imag_net,
    d0 => imagdata_net,
    d1 => negate_op_net,
    clk => clk_net,
    ce => ce_net,
    y => mux1_y_net
  );
  negate : entity xil_defaultlib.sysgen_negate_333ced04b8
  port map (
    clr => '0',
    ip => imagdata_net,
    clk => clk_net,
    ce => ce_net,
    op => negate_op_net
  );
end structural;
-- Generated from Simulink block
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect_default_clock_driver is
  port (
    brik1_sysclk : in std_logic;
    brik1_sysce : in std_logic;
    brik1_sysclr : in std_logic;
    brik1_clk1 : out std_logic;
    brik1_ce1 : out std_logic
  );
end pilotdetect_default_clock_driver;
architecture structural of pilotdetect_default_clock_driver is
begin
  clockdriver : entity xil_defaultlib.xlclockdriver
  generic map (
    period => 1,
    log_2_period => 1
  )
  port map (
    sysclk => brik1_sysclk,
    sysce => brik1_sysce,
    sysclr => brik1_sysclr,
    clk => brik1_clk1,
    ce => brik1_ce1
  );
end structural;
-- Generated from Simulink block
library IEEE;
use IEEE.std_logic_1164.all;
library xil_defaultlib;
use xil_defaultlib.conv_pkg.all;
entity pilotdetect is
  port (
    imagdata : in std_logic_vector( 18-1 downto 0 );
    realdata : in std_logic_vector( 18-1 downto 0 );
    validpilot : in std_logic;
    conj_imag : in std_logic;
    clk : in std_logic;
    imagpilotout : out std_logic_vector( 18-1 downto 0 );
    realpilotout : out std_logic_vector( 18-1 downto 0 );
    threshold : out std_logic_vector( 18-1 downto 0 );
    validpilotout : out std_logic;
    pilot_found : out std_logic;
    pilot_indexes : out std_logic_vector( 9-1 downto 0 );
    pilot_mag : out std_logic_vector( 18-1 downto 0 );
    pilot_pulse : out std_logic
  );
end pilotdetect;
architecture structural of pilotdetect is
  attribute core_generation_info : string;
  attribute core_generation_info of structural : architecture is "pilotdetect,sysgen_core_2016_2,{,compilation=IP Catalog,block_icon_display=Default,family=kintexu,part=xcku040,speed=-2-e,package=ffva1156,synthesis_language=vhdl,hdl_library=xil_defaultlib,synthesis_strategy=Vivado Synthesis Defaults,implementation_strategy=Vivado Implementation Defaults,testbench=0,interface_doc=0,ce_clr=0,clock_period=5.35716,system_simulink_period=1,waveform_viewer=0,axilite_interface=0,ip_catalog_plugin=0,hwcosim_burst_mode=0,simulation_time=1.1272e+006,addsub=289,concat=118,constant=200,counter=103,delay=616,dpram=34,expr=62,fifo=2,logical=4,mcode=21,mult=69,mux=279,negate=33,register=45,reinterpret=88,relational=27,shift=26,slice=184,spram=6,sprom=12,}";
  signal clk_1_net : std_logic;
  signal ce_1_net : std_logic;
begin
  pilotdetect_default_clock_driver : entity xil_defaultlib.pilotdetect_default_clock_driver
  port map (
    brik1_sysclk => clk,
    brik1_sysce => '1',
    brik1_sysclr => '0',
    brik1_clk1 => clk_1_net,
    brik1_ce1 => ce_1_net
  );
  pilotdetect_struct : entity xil_defaultlib.pilotdetect_struct
  port map (
    imagdata => imagdata,
    realdata => realdata,
    validpilot(0) => validpilot,
    conj_imag(0) => conj_imag,
    clk_1 => clk_1_net,
    ce_1 => ce_1_net,
    imagpilotout => imagpilotout,
    realpilotout => realpilotout,
    threshold => threshold,
    validpilotout(0) => validpilotout,
    pilot_found(0) => pilot_found,
    pilot_indexes => pilot_indexes,
    pilot_mag => pilot_mag,
    pilot_pulse(0) => pilot_pulse
  );
end structural;
