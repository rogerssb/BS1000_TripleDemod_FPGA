--  Module : ldpc_encoder_pkg.vhd
--
--  Description :
--    This package defines constants and types used by the low-density parity
--  check (LDPC) encoder.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ldpc_encoder_pkg_4k_23 is

  -- constants
  constant C_ASM_LENGTH : natural := 256;     -- attached sync marker length
  constant C_LC_k       : natural := 4096;    -- k = information block size
  constant C_UC_K       : natural := 4;       -- rate = K/(K+2)

                                              -- n = code block size
  constant C_LC_n       : natural := (C_LC_k * (C_UC_K + 2)) / C_UC_K;
                                              -- M = submatrix size
  constant C_UC_M       : natural := C_LC_k / C_UC_K;
                                              -- m = circulant size
  constant C_LC_m       : natural := C_UC_M / 4;

  constant C_SHIFT_REGS : natural := 2 * C_UC_M / C_LC_m;
  constant C_CIRC_ROWS  : natural := C_LC_k / C_LC_m;

  --subtype asm_t is std_logic_vector(0 to C_ASM_LENGTH - 1);

  -- hard-coded attached sync marker for length = 256
  --constant C_ASM : asm_t :=
  --(
  --  x"FCB88938D8D76A4F_FCB88938D8D76A4F_034776C7272895B0_FCB88938D8D76A4F"
  --);

  subtype circulant_row_t is std_logic_vector(0 to C_SHIFT_REGS * C_LC_m - 1);
  type circulant_matrix_t is array (0 to C_CIRC_ROWS - 1) of circulant_row_t;

  -- hard-coded generator matrix for (n, k) = (6144, 4096) code
  constant C_G : circulant_matrix_t :=
  (
    "10000000100100100100111101100100100011000000000101001111001011000111001110001000100111001000101110000111110100000100100100011111101010011111101000000110000011010010100100000010110101111010110011001000101101100111100111001111011000011110111010110101110110010110101110111001111010010000111101011100000101010111101010100001101111110000001111101111011101010110001001000101110110010001011110010000011000111111001011001101100110011001111011110001111001111111011110010010010110110011111110110111101011000111101100101101011011001101001110010101000101101011001000000001111101001001000111100010101111011100101001001110001101000101010000101011010110101111001101110000001110110011110010001110111001110101001111111011111010011001100011101000011100110010001111110000101100100010100011010001111101010101000110110010110101111110011110000010001011110010000000011110001001000000011001100101100001001101011000111100101010100000000011101000110110111001000010011110101101000001110001000001010101111110101110100000111101011100011101101010010100001111011111000101011100110001011101000110110001101101101011000010011000001010001101000101000110001001000000001001110000001011001000110011011100101111000111101001111000001100010110100000011110011101000000001011000010010001010110001110000101100100101100100010001100111101010111111000101000100110100000000100000111001010101101100110001100010111100010011000110011010000000000100100111000110001000001101110111011010101110000100001011100011011001111110110001001110110101110001110101001011001101010101001100000011110000000000001000010111111111100111111010100101010010010011110110110011010011011111010011111110001010100011111110011000111001010110010101011110011101111011001001100100000011001010000010000111111011101000100011110110100110100001111110001001010001010111001001110111111100011010011010001011110011011010010101100000000000010001101000110110011011000111011111111100010100101101011010101011010111100111000111000111110000101101110110001011000010101101010000100100010111001001001001100011100101100111111001001000010010010110001",
    "10100000100110011011011101110110110001100100001011111111000111011000010010110000110110110111100101110000100110001110000101111110011101011111111010011011101101011100111101111111101010000111001110010111000100011010100010010110011000001101101011110010010011010011110010101000110111100101010100000000111101101000110110110100010010011011111111110111010000100101000110110010010011100100011010010001111010101111001110000110110010000001000000010100110010010001101011000111000000000010100110001110000010010101111100001011000100101100111011101000101101011111011010111001001111000001000110101101011000101000110010110110110010111000000111110111011010111110000010010101110000101100100110010100101010001011110111011011010011100010110001001000110010010100001010110100110101001000000100011111011111100001100100011011001100001110100011111111110101101101010010100111111010011011111011111000000110111011101100001010111001100110000010001111011001000111101100011010111011011001110011001010011111111110110001010100100110001100000000111111000011110001000100110010111010000001011010111101111110100000110000110100010100001100001110011001001110010001000111100001000011101011000100001001011111001101011110100001111100110010110001010100110010001011000000001001011001010100111001010110101100100101101000101101010111111101010110001110111010101110110101000110000011001110111111000001100011100010111110111010110100101001010101000100011001111110001100100001000110001111000000011101000001010100010101101101111010100010100100100110101000011110011101100001110111110111011001001100011011000111101111110011101000100010010001011100000110110100011000110000011101110101110111000101100111101010011101001010000101001110101111001101100010110101110101110010111000110100001110111100011011110111111111101010010001010010111100101100110000101100000010011100111010000000001010110011010111101011111101000110110100011111001100000110100110010101011111011111000111010001010100100011011101111111010001011010110111110110000101001100110000001111010111011010101110001111110011110011100101001100110011010000",
    "11111110111110111010100011001110000101101001111111010011011101110101101100100010100000001110111100111011110110000111000011111101110111110111110010111001010111110010100101000011110100001110111010101000010001010010100111111111000011010001101100011100000110010000110010100101110110110000011010101000011101010100000111001000000110111110111110010001001111010101000101000101111100100000111011111010110110000110000111110110011100111011001100100000001010001011010001110001001100110111011111000000010101101100111010010111110010100011111100100001001100110110010111101110001110000000111101111110100100000100011001101001010001011011110111101001111101000100000010000111110010001100011100111010011111001100010111111001110111100111000110110111011010000011110100000001100011011000011010100110110011011111110110001101100000010001011101110100100010100100101101000001110000111111010110100110011001110110010101001001010101110001000111101101110000000010111110010101100000011111001111100111110000101110000011111101100100000000010010110000001110110111011111010000111011110101110111100010101011001010110010100010101001000011011100011010010110110001000100011011100001110111110100001110110111011111100000111100001100110100000110100101101010100101000100100110000111111010010010110101101000001101011111101010011111000101011000110101000100101010011010110111001110110011101101000011111110001101000111010001000100111101011101010001110101101011001011001010101110111100001101010000111111110000111110001100001010010011011000011101110011100101111010111000011111001000111111110110110111111010010111000110011100101100001001010001011110010011000100110111000110101100101101100100011000101010010110010110110101000001010000011001110011010100111100001111100001001110111111111001100011011100101110111110011000010000101011100000001111100000010111111111100001000000111110110011001000001101110101011100001111111011010011111110010010100101100001011000010100010000100100010100101001010001011000011011001010101101001111000011111001111111110100000010001101011000010100000101000110010000111100001111",
    "01011011011011010101001101001110110111100001001100000110100010100010010001011001110010110000011100000000011100010010000110110000111100000111101100001000101110000010001001110000010001111100000110100110001010011101110010100101101001001110001100001101001010000101110100000000111001110010111001011011011010101101010101111010100111110000111110011110000001100000100001110000001010111101111010001011110110111111101000110111000111000000011011011001011010111111111000001110011000000011011101110101101010000111010111001011011010010010111010110111110110100111011010111101000011010100101011111110100100101111110010110101101101010001100001001011101010100011111011101110001101111001000000000001010001001100101000000011101101111010001000101110101011011110001011110000011000011111111110110011110011011110001001000110010010101111000100100001001010010111100110101001100100111000000000110100000010010111010010101001111110000101010001111000111001011010001011101000101110010000011111100111010011101110111110100100110010110111011000100101111001010100000110101111011100110110111000001010101000010100000101101110101001100111011011100100001111001111010111011111111100110111001011001111111111000011000011010110110000001010010110001010001100110011001001101000000100110110101000110000001000000000001100111111111101010000000100010001001110000010111111101011101001011001010011000010010101011000100101101010101101011001110000000110011000111000010000000110100101010110111100011001101101100111111110000000101000111010011100100111011000000110000011010100111001111111011011011100101101110101001010000111101111101001101000100110001000001010000111110101100101000101011100001011001001101001000010010111101001010001101000110010010101001000101110101010011011011101100110110100001010011011100010101010111110011001001011001000110000000110001000010000101000110110101101100011110111101001110001110011001000110011100111011100000110101111101010010100110010101011010001110101010101110100101001101101000111000100110100001100000101111111000101001000101110001010110100010010100000010110101101000111",
    "11100010010011010111110000010111101111001100010001100010100101111110110111000100000110101010100110110101110010011101100100110110100010011000010000110000001001111100011010100111100001000100100111111000110100010101000111100001111101000010101111101001100011110100010101000100101111011001111001101001011101011101110111010100101111001001101100111110111110101101010100001010111111000101100000101100101011100010011010010110011101111011000100110000111111101101001011000011100111010101111010111101111011100101011010111000011010100001001110111011010100111100000000111011000011001000101001001110000011010001011010010111001100100010101000011010001100000101010100000101010000100010100110100110100110110110110011001011011111100001111110110000101110001000010110111001000011001101001010111110010111000110011010110010010100101110010111000101000111010111110110011110100111100010010110010010001001010110011011000001100011110000001000110100111100101010001100110000000001000001101011101100011010100100111100100111001010011010001010100011000010110001111000000100101001100101110011110000101110100000010111000110001010110001010111111110111110011001011001111110110011011001011101011110110001000011110000000011010111011110010011101110011001000010001000100011011111110101011010000011010010101100011101000110010011111101000011000001101011111000101001100001111101010110011010000110001100100110111110010011111011110110001111100010110000010001010011010101010101110010011010100101111101110100101111111101100110011010111001110111000100111101111100101101111001101100111110101001110011000100101101010000100110010101101001101000001011000110111101101111000100101100100000001001001010011111111100100000100011000111001000000000011111010110101000100101001111111101001101101101111000110110001111101000111010111111001010110110000101001001010111110110111101011001110110100100110011100100101110100100110101101101010011010011011100011010001001001000010011110001011011101111101000110011110011010011010011110111000110111000000101110000001011110000111010011001110000000011000110110000100010011101",
    "11100001011010100111101101110101101010111000001110000010010100101101000110000100000011101111001010010011010110101010000111001100101001011100100001000111000011111001100000100000001010111010101110101001001111101110101011001110010000111110111001010110111000011011001011010111011001111111001101011011000011110011010011111100111010000101010110110101001110110110101110001101101110001101110100001000101111001111010001110110100001001110100100000100111110100100011110010110010111010111001000010000011110001001011111010001001111010011100001000000001110100000110100100110100101101010011101100111011001111001110001101111100111001100001101110101001101111010100100111010000100100101110011100111000001000001111011000100111100111001101011010111010001010010010110010111111011010001001110100000110011001101100001000001101101111100101010010011110110110110111101110000001110011011100100101001101010000010000011110101010110101001010110101010001101111000011011001001011011100000010000110100110110100100011010100000100001000110010100111011000110100000100010101001000001111000001100011010001001111000100100101101000011011101010110110110110010011111110010110101001000101001110000001100000000110110011000110111100101001010010011101001010011100011111110110010001011100100000001101000111011010000111011101000010100111011110010111101000101011010101010001101111011000011010001010001110011101111010100110101010000011011000001000000010101101110010011011100101000000011100100111000001101101110100110110110110111111100111110011011000000011110100100000001110110010011001110111101000101100000000101100110001100000111101101110000101111100101011000011000110001101110000010110100101011011110101110100100011011110110010111000110100100001000000011010100110000111111101010101101111100011010101000100010100100010001110000101100011010010100001011111011000101010111010100000111010001100101010110101011110100011110111111110101011110000100110010111110011111111010000010110001000100001001100000011100100010100000101111011111000000011100011001010000000110001001110000101101110010011111110001110100",
    "10110100000000110101011000110000000100011101110111100001011011111001001001100011000011001111001100010010101100111111011111110100100101011110011101001011001110110101100000101101111110111001010000000001111101010000100110100011010110111101001001010010100011001010100000010110000000001111011001000011011111111011110100000000111111001111000011100100101011010100000111011110001101011001100001000011010011101110001110010000001111001101000110100001011111001111011000011000111010001110001010100100011111101011110001001100101000011101011110000001011010101110001100111011101001000110111000111010100111010101101100111100101111011010110011111001001111010101001110001000000000101110110100001111110011001110111111110001100100111101101110011101011010110111100111000111111001010000100001010100101101000010110111011111101010100111110111101001101101010010100110011111010011000001101101011101101000000101010010000111010101100010110100100000001101001001001010000010111101110000011000011110001100010101100111100100111010101011000010011101000000111110000101011101010001011111001011010001011010010100111111110011111111110001101010100001111111000001111001011000111000111111101111010110100001110101101101110001101110011000001010101101010101111010110010010110110011010011101101111011111010001010110011000110100100001100101011011101101011010100000100110111010011100100101111001010001010011010101010110010001011001010110101100001100110001001000101011000110001000111010011100000011100100101101101001100010011000101010001000010110101101010000100101101100101001101100000101000001001110111010100101100111001001001110010111001110000111000010110101101001101011100000100101001000100010000100110001001001011101111100001011010011110100110110000000100001110111101100011100011101110100100101011000011110101010001010001101111101101111000011100000000001001111001010010101100010000000010000010110111110100100010100111101010111001110000111000000001111001110010111100010111011100101011000011011010010000000001101010111110001011000010110101001000011111101111011000000111001001001101110010000011",
    "01000001001110100000111101011000100101110100110001110110101010110100110000010111101010110010010011110011011111001011000100000101010111111100000110000010011110100001110111011011000001000101011011001100101010100111111110010100011101111100101001100100111111001001000001001110000111011001001100111000110100000111100101011100011010000100010011110111100111101101100010110010011010101001110100110000011011110110011010010111010111001110011100000100101010010010010111100111001011101100100101010101000010010001100010001011001010110101111011000011001000010010101011011111001101011001010101001111000111001101101010011100101101101100110011000010100011100100001000101111001000111010111110000001011001011001111101101110010010101111110111010000001111101111101110001010110101110011000010000100110100011100110010100011101101010000001101101111000000110001111011101101111000001111000100010010000111100110111101100010110100100011001011011111101101110100101000000101100000101110101100110011000000111101000111101001100010000001000010100110110010010010001000011111000011101111110010100010110010000001001001011001101101010111111110001110011010010100001111010000110011010011011000001000100010100110010011011010011111111110001011100110111001111110000011110110001111101010111110000111001110111000101001111001010101111110100110110011100100100100010111000110000101110011000010001000101100000010010011110011010011101101011110110110010011111000011110000100010000010011111111111001010111100100011101100100011101001111111011001101101011100111101111010110001011100101101010000000011110101000000001111000001100101111011010101100100000111011110001111100101001111111011101010100101110111100011111011110011100101100110011001000010101000010010100000110100011110101000011101101010100100100000110010110010000110101011000011000001100100001101110011100111101010100110000000101010111111011000000011011010000000111010000001010000011010100011010011000010101010010100100101010111010001010000011000101100001110101011010111101110100111100011011011010101111100010011010000101010100011111110101011111",
    "11011101100011001110011001100000101101110100000000111101110010000110011100101110101001100010000011100110010100110000000110110000100001100101101000100011111111100101011010001100000101110011011001101001111011100001110101111111011110100001101111010111010010000011110011001111101011001000010010101011000110001000110110010000011011010111000001010010010111010000100100101100001111100010101101000110110001100110011101011100000111001111010010110011000010101011001101000110000000100010111001000011110110100010000010111000101000000001110111000001000101011001011001010010111010100010011000001011010000010001100101110001101100001110001111010000001110010011110000011110011101011010101100001110101001000110001011100001110100000111110100001000010001111110111110101001110011111011101001000001010100111110011010110100111101000110100001111101010000110100010000010100101110101010001000000000111110100011100011001110010001101011001010001101001110110100000001010101110001100011001110101010110100001110110100101111101011001101011010110100000101010101001000110100111110100111101101110010111101000111100010100001100100111110110000010100011010011000110001100001000111110011110010110111000010111111011100101100000101011110000011011100111010011100110000000100100010100101001001101010110000011111010001101010100101101001110000010000100000100000001110010000110111111000110110010000101011010000000100111000001000000010101000110010000110000010001110011000101101110000010000000101010100100000010100111000110100001000110000011111011110011001111110111100000001110101010101010011110110000011000001001010100010110101001000010011111111111000100011011101000101100010000010110001101001010001001001011010111100011100110010011010000001111111100101011100011000011100010111000110110001100010010111110110010011111111110011011011111001101110110100011110000001101110110010010101100111111111001100100011111111010011111010001010111100110101010100111101100100001011110101010010100111010110100110011011000010001011100001110011111100010110010011110101100110110001110011010101001000101010110000001111",
    "10100101110010001010000000101000010010010101000010011101111011001110110011111010110111010100110010001001110000000011101001111000111000010101011001001010010101001000110110001001110111101100110110010000110111011011110010101100011110010110010011101001111100000101010001011011001000000111100001110111101110111010111110110101110111101101011010101110101011010011100101100111110010100111001000100111001011100001001010001100100101111011000001101000011010001111110100111011101110000101100110010110011001000000010000110010001010011001010111101101010010011011010100100101110101000111110011101000011010001110111111010110111111011011101100001011101101101001011101011101110010000010110010000101100000001101000000001010101111001011100111111111110001101111010100110010101000001100101110011111000010110001111011000011101111000001011011000010111001111100100101001111010100010100100111010000001101100111011110101101000000111001010001010010000110000000101100100100110110100100001101001111010110111011101010100000101111001110111001100100111011011001000100000000000010011100111001101100000100010001011110001111010110111100011110010100011101010100111010111010011100100000000000111110100110100101001111001101101010011000100010110011001111001110001011010000101000001001011001011101101010101100101000100011101111111000101001111010111001010011001100001111010010000001001110101110011111111000111001001111001001010110011001101110101010110011111100000011010100011011110100110100101010111011111110101000100001110100110110001000110101011111110001001110100100111000010101000101101000001100001000001111011111011111110100111001001010000111001010101011110111001011000110011110010011110110111100001001011100000100010000100110011010111001111010100110111100001011001100011000101001010000000100011101000011100101000111100111001101011110111001011000111101011111110001000100101011101000010110010101011001001011011001001111001111010001011100111100010110001111101011101001001110001010111110111001001101001100101110111001011100100100010111110111101100011010000111011101110101001100010101011001",
    "11000111110111110001111010000010000110110010010010011011111000110101111001101100101010111000010000101111001111011111110011010000000101000001111001000010100000010100000111000010100010111101110011110101010010110000100110000101001100101001111101101110001010101101100011000000100000110000011101010010001100101011110111101010110111101010011110010111101101101100100111100001010101100000011010100111001010111000101101001000010100000010101100011100000001000100101110101000100110101000110110111100010101001110101101101110011100011000111011110110011011100111001001101110101001110010111001100011000110111001101100100010111000011001001111110000000100101111001111111011001011010001000100100100011010001011000011011011100010011111000011000011110010001010000101000011111010011011000101111101011010111110100011101010011010100101001000101010000100001111010001101110110001011010010101101110001111110101011100100101100001101000100001000101010001110101001101101010111111111010110100001100100000101010010000101101100010001010101010100110010010110000101101110100000011100001011111101110111100010000101010000000000011011110000110010001011011000010100100011100000101010011010110000100010100010001010000110001001111101001000010001101001100010011101101011000000000011000111010110111011111011110110101100001100110100101111101110100001010010111001100010011000010001110111110101011011010001101000101110010010111011000111110010101000000010010001101001111100100000011010110000110100101000001010110100110001000100110001000001001010111010111011110101001011000010011101010011011110111001011110000100110101010111101111001000110011100101011111001011111000100110000111000010000100010011011111010001011111101011100101000001110110100111111110011011001111100101000101101110101110011000000011111101001100000100010101010100010111011110110101011000111001101011101011001100010000111001000011011001110101000100000001111101001111000011111110010011001001100100000011111101101110000010110010000111001011011000111110010001111111100100010011111111001001010010111100110100011000100111001000101001101",
    "10001110000111010100111000110000100011000000001111110110011011010111001111010111011010100111000101011111100001011001101111101101101111001000110101110000100111010100101111101111110000010101010110001101011101001011010010011000011000001010100100001010101110101011011001111100011101010000010000011011111110110011101001100001101110111011101101110011110111100010101100111101011110111011010111001011001001010100111100010000001001010111010010010101111000110001100001011100011100011100001101010101100111011001110011010000101011001011011110100001011000111110101100011110000010001000011000100100111110010100011010010000100110110010100110110010110001110011011100111100010111001111010011110110101100011111001110100111010111011100010010011011000101010111010010110011101010101011100000110010011111000101010100010100001011001110001111010001001110000010111010101001000101111010011111000110011100110000111000000001101110100110101110100100001101110110011111010101001111101000010011111111101101111101011000011101011011101010110100100100101011011100111110101010110000100110000000100100101000011101011001000010110001111001010101000000000010111000011001000110010100110011101001000011010110100100111111101000100110010111000001001111101011111010111000101011111101000101001010111101100110101111000010010011010100110111010110010101001110001011010111110100101010000110000101001111000110101011010010000100000011001111110000011110111111011000110010101111110010110000011001111100100110010001111111011111001001100101100010101011101000100011111110001011000010111001001101101011001110100011010111001101111011001101001001101100010110001011100111110001001100011000101011110100011011110001001101110110011101110101100011111100000011110111010010110111110111010000010100001010100110110001101000011100011111111001100010111001001100000100101101001100001000001101000001000000111100111010100011000111010001100100010100111110110011100001000011000000101000011111010011110111010010111101110110110001101010001111110011111110000111011110001011000001100100010100100010100101111010001000111100011100",
    "10101001100010110100110111100110100011011101101100100100001101001000100100111011111011111000111100101100111110001101101101011000010011001110111010001111000011100011100111010011000011001101010011001000011100000001011111100111111011100110100010000110111110000010001100000010010011101000001111110111011101111101011111011111000011010111111001000110101010001011010111111001101100010011001100011101000010111100001011110111100110111111010101010101100111000011001001000001110101011011110111000111111001111010011001100101100111100001110111010101000000110111001111000001011011001100100101111010010111100011100100001001001000011011010001110001111011110101101100111001011100110001110011001100001011001011110111010000100010000111011000001000000001101000000011111001110110010111010010011101111100100010111011100011101010110111010110001111100001011111110101001001000000000001001011111100111111110010000010110011001100101001101001010110010010001101001001011000010110010000001101101100000001011000011011000110010111110100011000100011011011001011000000001001101110100010011001010000101010111010111111000100010101100101001111010110000111010010101111111010001001010101110111100111011001111101000010110010010110101100011101110011011011101000111001010010000000001101001000011110111000111110001010001111111111011001011011110110001111010000101000100010110011010101011101001110110101100001100010011001111011001101111010110100101111101011001100110011111110011001010010101100011101111001000111111111100010011110110001100000000010111000010101111101010011011101110111000010011101110011110001111101110011100011011001110000100111110111000000011000000011001111111110101110001000101010110101000100101001001010001000000010000100010010001001001111100011101100111110110011001101101010010101001010011010000001101000011111010110010101110000000000110001000001100111000111100010100111100110101101101001001001010101100010111011111011011110000100111011001110010001001011101011110100010111000001111001110101101111011000010011011110011111000001110001101001000100000000111110001011100100111010",
    "11011010101100001100011111000110010111110000110100001001011000110101000110111111100010100000111011101001110011101111010111110111011101010110101010011010010001111011010011101110100000000100001000001101111011111010000101101011000011100111010011001111000110000000111110101011100001101110011101100010010110010101001001100001100001010010111000111000111110011101011110010111110101001111011110010110110110100001100000010110100110101111101011001001100111101000001000110101110101001101110101101100001010111011100010000111000101011101000011110110010111101001101011011011001011000110011110101000100001111110010111011000111011110100111000010000100000001010110010010110100011110100110000001101011001110011110010100111101001110100011101011001101001111111000110110100111000111000001100011011010101100100000111001110010111111010110111100000000001011110101110010100011110111110010111100010000011100111110111011010111101100011011100100110010101011000001001011011001101010001011011110010111011000101101100110110110101101000011110001001010111110010110000001011101100110101111000111100001111101101101000110010110000011001101111111111011011110011101000100011100101111010100011100010010111000110010001100000010110010011010110011101100100001010000100110111001011111100101011101110001001010000101001000011100010101010101110111111000101100010110001000100100110011111001011111110110011111010001001111111100011010111010110000010111110110110000001111011100010001101000001001111010010100110000100000000101000111101001011111000101010001000101000101110010111101000000011011001110000100110110000101010000000100011100101000011101111000110001011110011110000011000011001011000101000001111010111000110010000010011000010111111111100001101011101001011101110111000010111101011111111111111111000011001011111001001010011000110111011000000101011101101001110000101001110010011111101101001111110101001111101111110011010011101110111000000011000011011100001011110010011100111011111010000101111100010000000010011000001100001111010010100101000001101101110001010110000101001100101010000100101101111",
    "01110111010100110110100110110101100110101010100101000000110110101001011010110100011101000010100111000011001110010101001101101011010100011110110011000101100111000110000010111010110101110110001011111010001001110101101001101010100011111001000010001000010110101001001000101010100001001010111000101011000001101011010000000000001111000000101001111011111000100010111110110010000100010011011001010011011101101100001111111011111111000000001111101011000011011110101000100110010011110110011101101001101101010111111011100010111001010001100011101101001111011101100001010101001111011100100010000001010111100101011111110010001111011010110111000001101000111110100110010000001100001010101000000010101000110101001010010110000001001110111001001011110101100110110101110111000011111000111010001010101100111100100101000000011101111111100001010111011100100110010001111000100101111010011101101100111111100100111011000101011011111100101010100111101000101000100101101000000001100101110011000111001110111101110110001000101011011010010011010110000011001001010000110000111100000101110011111110111110001010110010111011101001110011000000111000010001100011101010011010110100111011110111100101101110100100111010010100111111011010100000011100011011000101000110101011001111000110100100100000000110010000011011100001001001100001001111101111110011110010001101010110011100000011100000111110110110000110010111000110000101100001110010001010100010010101100011011100000010010010100010011110101000000011011001011000001101110110001001110111101111100110111001001110011000101010101000111100100100001011001001110011101110011000011100001010000001101001111111100000111101010001011001001010101010001111100000110111101110011001000001011110111011100111110100111010111010110111100101001011101000101111010011001010101001001111000111101011000000010000000111000010100101110011101111010011011111010101011001001011011111010010000100100100001110100010000001101011110110001010011110110100001101010100001010001011101010001101110100111101101101110000010001010101010000011011110011001110000000000000111101011111",
    "11001110101010001001001100000101100100010100101111101011000110111110100001001011010110011010010010100001100011001100000110101110101101011100110010010110001100100110101011011100011010011111001110110100100101010111000110011000110001100000101110110110111001111101101100111000110001000010111000101001010001111110111111000011100111010010101110111111101000000111110000011000110000110010000010100010001011000111101110011100011011001011111110110111001011100110100100001001101111011100000100110001101100101110000101011110101010111110110010100110100111011101000100111001010101010101010011001000010100101110110101111110111001101000000101111010011000010101001010110011100110110100001011110110110101111101010101101011011110000001110100011000000000111011100000110000011111000111100100111000011011111111110000010110101101111001111000110000100100100101010111100111110101011001001100111000011100001101000100010110110111100011100000101000110001101000001101001000010010010011110110001110001010001000110010001010001111111011111101110100000111110000100100110110001001010010110100110010110011011110110001001001101011001111111010010001111100101011101010001000010100000100010011100000101010011010110111111110101001010010011011110101001101100100000111111001011110111000011001100110100011000101100101110010111110011101100001010110000010101001011110101111101001000010100000101101101111001100010000100101000010110111010110101000011100010010011101100100001101001111111110101000000010010101100111110000010011010011010000000000110110000001100100110111011000010111110101111001100111000011111011011111001111110001001101000101100100001000101100110000011011011000001101110010101001110100000011101001011001110000011101110110000111111100110010101001101110000110000101000000001000010011010010101110100101001000100000111000011111111111001011011010100001101111111000101011101010100111111001100111010111011111110111101101010001010100100110011010111100011011010000001010111000101001001010110001110111100110101101111010011111010100011110011001110000111011100010000001011101110111000001001101"
  );
  
  -- functions


end ldpc_encoder_pkg_4k_23;
