

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ETvULKUfBYvpKJdYQkTkWlSnvEbePNGdQh7djE8T3h9Ss/WywoAfFVd5fBOhigCD+SiqthiSN3yx
eCWNFTRHTQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
iF0ra2wFoGarVDLaQIrIocIa4wBHPu5oKv21QKN1lZAhxy3NTUfaMnpCbqz9ojy4NzTFwhfrG6U8
oec0gR2G23/FnNqpmkms70IKG2ER70/sOpPABM3ju72YxbyjULt8OUXa2F1qybvUD+2thXH+u3AY
w/3Lp0WSRNN20zDOcjs=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
GynVkEHoyvKwR3nDmMyDxiqfUdn81oMrs6TH7gd8ZgoHjyLQc+hvIryt+s3c9BKmBNxStsWZLqZZ
z/OJwlYNz8jk7BzRRNLZWRHVUxbZmkTAlMrSypXXx1DjiYucMxmi9/uUw/NZ8Awf1Us1XblZbFyH
Au1f+BvzegUa7bV5KCo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
R/oYKs95fKNWDaMZ82CVdXM+2zHjd+/lISntUYmqbYMlgMmX9Bsnf6OoC4zUKoAGL9JgGzjhA1UF
f/+95GFJXgLwfGZ+5l7kEcZtmKWCDcL7WRMxkZqdPfYqafnamtEIP2KM6H9Z9pxz1sF0T3JHWgmf
wpuwSCqSZmV5IjkedEj5cKljmKGshs68ty9K7u4tsDTqAZ1Ep7tBeAW1PliEagd7+YQpZcVT+XYp
eYiv2dROnsPi58c1GJS89Hm7tEy9RwzhG+bj97casYHJAG8V3OXsO/+VhiT8rD2cZpVzZQYh/l/1
BTwnm7xt5q9jS8mC1/yWy1GvkH+Mo1gY3aOzcA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Kkz/REdmaH8/zbTviF33/TO1VhDO2iv0g1fAvgx6nk6gz4daDZ3a7yC8ejlHmZ8R9Koi9FZCdT3M
Aye8agyZGFk0ApD/vskf/BVf+UnPRG2l2oe5DlWJICQWSR4IjrwWf+WGuXKnapljP0ulXC9yEs4U
0B1QeBMig9AP5DxR8NweLdtA89Sm+r9cat7NInE6w93lwOCDB7W4eFBvTvyagMd1nrjqwFEDUdF3
iR6BGwOPEv6tOtZOYLiuJj/GcnBbn8AWszDfzLL4y9mZ7mhF9BdIjgHOsN1BtwnzQhGkYVl2WbZA
xmlHVMdSIV/V9Ks12hz2oRhXjmossadlG8WRjg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
xK/yf5SFYOOh/C8PaaLVxyHQCCSdSwq3WuaqnUmrR1FLdcEhiA5BePl5ISQvgSIX2I4lg8LF7PtZ
JcEfKbd/Dd4k3IjgHX3JnDuyfw3SX9oYm84eKzvAq6ad4XAIilNCe4JXXT04fW6J9XVSWhtPSGnA
U0zGDOIbM+zOlwegT37fP0KWCyVHcERbN9O4jpIjSB2+DoDkZIgTrzW5om20eo/4z/+XKXLuIlqz
Cg/tfDjUWxBBPopw+PVmNkhb1AtWA6I+eeYlXpUW8Ro2wjg8Di9AqdG5YhRj6dSa9Yc9ajmCsGXN
vVM0Pn5iSd5uHmPQgl2rSiSAu42tJIVbgzwZ1g==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 121856)
`protect data_block
g7ish1JsnpyflaLPGK1fCG7Tg+VrlkZgFk1IuNURlvfZUBDJmpOX6+JJXEjsRKirSEIShehAGcKw
aKIiEmzOD98F2ovcdI6wxiIsPtwLuIDag4C8a+/mbd1xRC31XY8NKXxENmPvgwn0/QUI2CNdPFiX
e20S0HomAlKCrfDc1Rr8ZO8ygvj159YtnhdLlM9/IfphrAGe3v+7ErRjHl05GBtLOIQF1u+JnSTp
xgC/CAQrGF9q6jlg5DGpayRMSZ3LZyDcci41zoXlDmRpnaVs6M7lB4J3gCgup7iiqI40AnEGwgAP
pLMJXc4gBOcgR49BcSng2tgkm9cz2fQ+dgcf01oPWvH06WzZIT/+zZ7Ho0xWBjDrUWWDPOeh4rgy
RLRTXyUlzblnLwUfZWw14KyXbA56xTrMhlQamnoLTVsaTMq7qmRJon5W5xPdVBCED1h8FuVETj6F
SMn+aWFF4KBNUdkYl/lnc8u19gRMNWHIiR0fxgmwwjuh5aSflseP6WXrdHJ/u15AmrNeul+gZHUB
vFEHUz3ybF22RFBznVUNM5XTDMbVWBNxwnXQbPX5f9NfQlMC8B92zASqpZq3ufG0I6eeQ3vj9SB7
kCi8CeQw5tHOGjU2KDE6D1fon0OBAejO5e5p/XK0UXeSsEM7W2tJa+OZR1jo+vkshTw7m3u1qD/j
5SVrgc12K3Kt5bh39zfYW+crf9oHftSzE66lMUnXDf40/OlyCnZ1PhcZ0o2g/+kZ4dZZeOuFbWhk
evTA+iLyMmQAXHKVEklTYegSrmj4biU+d45jD8U0wcU7F5hE4m0rkhYfOQq+ZTn3ZoNtmdYsyxMi
Uoid8b9kU0x8LqcyXs2sX2fG8rQhihT/CJUGaxIdClBM6UQKwTA2ERsAZMNynf+BbKFEhou/Zqg0
JnCelLCpKXhxYfmR9kqZFRXxCi1Znqxcf7mQP/Qlc3T7zd5ZRMbstcgy1hNsROj4MJM5/8cMSwF7
m27XUjIJ7d3A0gAFVDKXUYZ52AxNjYxtXvFe78jTWCsi3EvaIIRb/X4v6epeLnbrtV9ImqubnFJe
TrIq9Fo1HA/5006OUb7tGlZcgFzF04xhx9vKm7FR3juX8ohpE3oovRrRK6DxeDe8Ot4E35cj8T24
rxvPTcweE6tG9OmAm1XXIHtxq5FRPSSlXZ5w/jyR+9qn9pzd061pfWC5kNzIKo9ly4939PQeluvM
tPXYQB6qzocba63vyvKD4xLZgc7FvhUyAFZNi5EMi5rUina4QgkSc/Rzw9ReVrYKyXcS2Hfkx/CL
QcXUTI6EmrwVREr7RJhj6n3ZSVFECvt7QBzhOAech3NbEDPfiJpb5NNJWXHNxm/+XpKgLsQlGh9t
lGsC9Sv0Em8BsXFt6G9d3MMLBAe3V9ch59WZW5PeAWGzw/upSloMS8qK9ZElFvrlF3CPOGEav5ee
nFoCeg5bTr5Q9bhvqYlI2kJDLIUd2XXavaPCuiLSQstqcfoyRGC4rogEaomfzHa4gayxFtYDqvGX
fFhLjSzlu+VhZI3a5/Ol+dXwSsJVEl9/0sBSxJiOwj9/g5K/ta/3pR9fnFT0gdHQOcMtRjNFMsJ8
slIT66gRj//3ePzO5yyqAjHDtj47FZZnlILFNTLa6vgXKjiebMeCjZt7udIJmiVwuZk6uqP30wzQ
4SSxYc7n/VlbPFsSqeANGVq1m/6cDHQdj3+oGbeOYRpxx0dxc+1dK7otbiR3f/xN7JOSL8mEF92t
o93Mj6mGEqWiUiaxtrxLt0khPPrg4z1H1EYoJgjFiHUx+hPRLRIDf/EFJhQR1spC4V+Mj+9GaFFm
f71l/mPi3g3m0x6QJ36pW2jd6nXHEsq3pwtJ/K9cGdqGylq54ZjcxBj5VPes7KW23cQ90xHsCr91
4Bb+WzpKlXsp/B+s99RT3yepOR8y6i/1/SyPVj/rFfsZVg5KAMuwchflg3S8xaWKLdqQMjqPhJGt
h4dgmira4SRPkwgM1C8VI5nBzmNbqqXFeUFSC8vuxWEubOZzpjE8KViPlHPahOv4qkfqCc1B4jYl
r8WTChoxY+xVuqgkXH77SHNys9Fb0AcUsfab5P6bhvdX7Z3sLOUnLPY/UQIebKkKH9KL75nlzDkq
Y7NQ28waam9tnKwpBTYEUX5LNZnrloHQVib0WprCWRBaOtjUTvo0n/pqdBLHdlpfgHJj3qRnzfqH
v6Cnj87Grt2VnAi41XODvR7MSgUVTHKhVfKbv52wX02B+QE+DnJm4eO65QctCoQJC+T1wUCGQZbC
tOsN4V93lzRfkwIPDM2vSMQ71Rcf18hABbUeZlEeAVP6rWFqGEZlCJc+rPmMn4bDqJ3cdW9UW9M7
7vcFKyNPFLLjbsT+xsejSth480u6IVnEFitf+UJl96Cypeul/icVSkwLMcP0ynn70YbM4XhV5oh7
teK9dswsqA0GabjhfbYPW23OvKDJW6su08rCs8yGMauUiRB8AV4dmZ+ly2OLSz0o2u5yYOBHCP34
gxTVT3nUDjFtyAuyIfkjIGi0+cU7BVoKBIQGaW0oA6NEJ/G6QDFpglHVkNLIan6BBwiIVWcvuEcs
Gok8oPc9COrCTdeDkprgajzi3qo4P0+5mcfbmx3L3ax/9+kk1FFvj2xhSEmWoZA4fnmMVQiTyndk
x7XusCMN8Q90S+zBMJNXrsG1in0GajVdU1jRlYhlNp8iNprvzohLUJySAHzW0IUYDvVAAJTMk4wx
69Y3CKRreUzf3sDm0mEEyVK8wMtRlgvHzXSA3JXCcelU19NHm1tBVsfQPajkLkhF+cZ9hTBJqixT
90j3VsLAq5yQaM7sriGAs3ShM1IfVMwnlejDN7S3Py7ArorGOCG9ZlouwC7RDpNPw5eHvd6ntGiM
sKzrO0Q964bXcSZ4tw0suGvDaB/ij84CRKy7l6VxZnacWvluutR+ZjbfusUUVcaY18BXLd3Im96g
iOImNHj742M893Rmyh8kyU2gcqw9/63OMn4eCExNS/AXnCoTScjosHR82lwtF3bwsfUTEi7NkcSW
w/j6tT5IbN2Yhw/TWw0Yb8lELkJ5kgMMxQsIe+V7DqB4PiRE0i9IFcngq2g7k4cLRbzW52Cxyful
5z+4xaOi3Yjvgbyse0bjlazE1YbTDI9aDJQj5WlTW4TJnAgLLmDzKTA/n2GQ1vUowxLlms2OCQU3
D6+ku7rHzLJgvRjhcm5YexbMXnBzZQCJMH9UoyHDHTWQgpRixETsOZhqEUqkJW067ymybPQLUbtv
vzf6d7ampPvsjme/j8DgjBQqOUHrEg+9InYWUkqlDOEMBlZQlhXQd6+FNko/bkvlbOBHRmQaKawm
UnbDMHCLb5UefPGNsIYOqHYvxrUgw5nmnnUS7KjvcFPxnS3bkO7fK8h3VDw6CMb7WnJPoCHtiP8Y
3Wxzmp7gBORUUONQUrV+RB70aaXYvyFDTAPkTh+Zbw18bYgg6PcFSBUrpFsQ+cAurQ02cha3ldZU
PYtpxXQgst79aEBt5nKqpw7DEpldPHciKNGB4qBYT6LkfLJvuSNIb7iXuv54xDSvEO2ZLaox6nyW
+haF13PbkbAx0jXt7GHEWhO1Es/Y46rYoqrqTtTWeNSdbzrwXemwWvDPXfFGrcYNxmJFzKR6YRtl
lPt7+FuwKZAjgDv8KicxUonAvqaoQ/DhiI4KITmTRZh8uilG5mq5ITwfFtVYlEidgO1tqpHZ2o+8
69YXHRSfTXnqH3iptqhUPtCr+XlJJJRXeEKoTl3Cc/i+s79m1be+onSmk34Uy5qnxu+cruZ3GN3U
1yK/bb8jCp2+2FE7nDB/v6IeMh20LEvM+/6pOWL7wlkDkPRZX7AuVpIGNrJA3gm2/Dk/Ppw4HpIC
XPUe6RqSmYsia86cE6Y44Ej707V3vtXQVWIdrgT0Ep8YuXT3Nsz8DNxdYVkzFQXUmgqgReP0FMqT
7LgxbB1gbxL8KSe5H2a7WQ6FnMyv3qygR8xQ1i4/kYtnsy5LAGgdq3bJMbLVAP6/8iluK6ZywMb0
C9tFnRYioc7eKlj9QOEmwyO9rNXgqVlJKJ60FbQNumeTqsPW9GydM0QrpGZmOkeO525mTANJrx5x
CH2DJtw5f0cLONcsIqeGwuGEQSYawjkQNHAKLrDZPlZzKrAmX0F23cB5r5sj7Y+RxexX0MhWilpF
Bx0jfua/dEp937FC5nXCs/HCP78HrwCCCu2aPpLZTDyw56T629zBisVYlIQ9jrHJ4UQPwCkYSSLF
MyaUCFWKTYjPcVeH4C9ruTUbnRLAEED8LxxTDKTWKYovu30tQ+jqu/1vq2C9u69WY9RJlk5e3LPA
CQxjQp8FQdSoXTug4ShYf5FNtBxaoEyeL+1iDHoPpY+G61zJ3EIyunwkT5XCYIoDb3F9+49TY4km
X0aH2xiSuAWgPSTGNQhbO0cqdl94/HriQri1TGAcI8MxYglvineOmZeccbtOXqxJEhlbDPnGKUHg
0M39HIgnSZHGedFHL30n4Agk3onOsJ2UbBVlyzeDHK0Dxd9uoB/s4v2x21QUeslOPTzH6KcG2Js/
eqqqeJs8COS5TJD8mGutEAuerhMwjWsi+mCOEXoTOfYu/1Rtd3ZAK9LuI9NSe73zhOiqeUJJwS8D
Jsgo8z1u1HzfaWy7vimJ72dM27xg0rylrX+//OTcGgOSDi3pt4S8xzCObB4PKgkvEqvzLrSqc4Nj
7bbvEFSy8dJFyc0+3oQwNpjSPe+YKaShrxIh+F8wIueZJt8RJyYlKTFXZ2TYuHG0D+4LCDar7xdq
lYam56L7ImWzv28b4oCBNtHgpo0Td/oOXisTJ/sissoXZBJzvjZrjg6UzFcdOBM5jEyLmqa2iH/y
CwvLMA7UvFzmJgPSjnM3zteYrC/8zzajjXcgntjELaOTWBS7VJgkRCkCvKcHWfh6z1ZhghCZXUqR
Y3WwYZ7y/xRQfMaQLeTOfOXVI385d24UVzGEfnMhqCG6/cJkf39uWCpIjxoAI3YvAGr7XGErHdO9
8kpqZbcltNCtZ93hczVU+E2BUHhpSKhgtY7E3DcdmImMSH/N6cYEkeQmADNRvkEZqpxRPfTW6Vdl
vBG85+OFYt5sUf2w6RyGoBBAA9ndhC/AUfVaOPM4ZJnbgFNtkhp+laVpEM9veRs6PWqDO+Bms5t8
LApwvZE1w//pQ31pQbJKhfjS3o+tMDlL9ZgWzQB2dnSX7ezBQn127wK0n8kSzwIUhhnfctQzfSQS
V0BvSyusJdR/nxMEneN3YPAbwSCHuAL+3Br+UNscLDOrQkrCXp8+1wMiopHNFHt9pnCsgQAYTPuA
vMZChqrIfbusTs780RlI+WVPtQa4LEasQT3JUoGoh5/IizHmw0Zl/Xtp0KBuanncMBy6MY389mF5
vGTBDRv3qiFZPJSTcH1Yyhy4J6wjWAWfdgiLY9LifH2TwXnmgwgb0OwmmEHkEl/bUqqIw+K+WS+d
PrLiC6Pk1PXIQnaBRHrsE4hqY/TqIJliCsuCAM6jy33I3ven+4UNJhCL+hrqAMMSTBMs2faoe8uj
HERUlNFKquIWs3Z8Dx31yOBqsNSaIG5ealzQdpVqPAhiUV62FMja7orniHJ81vigf5cdb0LKyMcS
cYDwEyyzZDn3ogHyJOFCLsgGYl0O+XBWY454VbIDue/s40516hXjrlOGU8OZC2r2oFTpTw9QfTFR
6OlfNSik6ZNRae3r+LXXypzsezihvQFL18gFWmFLS/PosckQ6w6fCaVEH5l/25aN3N6aaST4u7YK
RRkbGyot0BtCYDybtuPx+IS4x3574arEbCiu0Xj3xMeLB8K9aCvN8hPocSPgOWtRE9Jm1BcqPBW5
gncx0YetDuKsqPjaT7Md4/ywS+tYNyFg0kL+VsPQWNlVB9afIaTqnP0eB8sEvcbKDgH0gBATxjka
3aLA+q1wgMVBFlW6DqFyAm86Gmlcxcf+7Zku1gaC57fHjzZGEKo1kHgddZf7xNx+SMcZuQX7bHMX
niJzGBHU3hiCupjdD4ob0KL/B8IB3pUpsexnThsoBMZlhst3mQW4b7Cruu03o1yo64m0ngJzVbG3
Mfr9bf3G/qJxYYl/eZMhSZqlbgwIFXjMxAoFnisBU3b0hHdJ8yj4uNfNJAM+y38Qm8l3XjQo7lCO
iNjR1plSpAbeylmO/ToOUXNZeGgn8iWG3iNYtbrk56cNRCFthrpSdRCI9iru9/K62ujXFWNcdey3
o0/J+YtR+6kBwqp/UJzMu+oScYXZog+Rp57Yc96IO50vsucGipaT+9g79oxDqVwUn67WajEUetjp
4S1ZYPFAJlBOxwDZQq/sL/KY6Au6mPdrNt4KCV0Gh52Py2pGaHkXq+j47EUugEhdnaRi8ALf6vW7
Yho59r2AXl0afMvJdpyQfAmWL/u+I/qCimSNgCg76BuFWFt0fcPljhwfa7XeloZSgp9GA66bLIh+
FuBapaieAW6ieToNOnGX2rwLQ+YHxY5CueTNheYJWGXbjpQUgwJuRQSnPNwUU3/cIi+sjk0ZKQpE
1VlPyvscHcKUWFREwzWdmf61C9/h0Yd3hptL/Q1SjCuUjGUYkJpK0zP51CtjyJE48wymLhds1D5V
thwaYW/eDol1ibzrMUzbQTPI2n+HLNuApJMRJmtMITMPYCgU+en6XfsRYq835/DvPPohafqZAV/g
wsPUG/ndkYoloRIrx/2NbFnAArcE7FTyiH1KvmtV0bF7qQlZwsgrLxCpHXzhI824o2wiay2YqNTS
nKUp0u0df92Otcd7SmtKPLfvwUgt/PdJ6Ich5lPJj3dGmBLM5fZ0ZW8CzKnP+z1DJ22ciY4AWVG4
bk+b+KxvPivQFeKpEkhLUotK2KmaC3J+gXSpRjXO+e3T70w7kFZGKFaNf+INGpXF0tAOB3yAIczy
08/Hzpcn9vCJMQJR+NyqwushmMvcCbNjdTJr42OEDLTH346oTwhKWu77R5ggBbgJl6SACtXAD2lX
PhqtXbPrGdX3x9GlTdh2dwW/lsZr1PJ+8+2aIVO3opAmElmV+Or71HHevMXnwzWN74vQpI46WWr3
W4rGcS+4W4EERxS9s2L/0leVf2L3iIgC1JfqdAIG6tc80JSTlHmjgAErS0WryJf6FWQr95HyW99t
rlFTrfkX3swTIQ0AGRcmiV9rZHKEG1EHCawjLZWdGhol9cuP7ryYGX0o4qIRvFHjgiwFI7m/mYIl
UYrWPwaPqQg7ScapVGYD42xKr85JMqSRnL4f378J/pNiR3Bxd14NCJ15+FOEKd0/ZCLHvPO5XpIh
OTFTi4lKExosIm5b6AJcCqPQksWuCs4q5ASKGYZLzNEjhbYf96rHcX0N4iVN2c1C3himNfnT08c7
rpU+tcGr4iXuimvFKzeIXFwS8TL/knSrQkc2wmSzmMpGt3wE9ggQLcHuR789dS2Je7IEdz1jEW2q
yNvcwFc48Vc5icnevVVIvQTlK8+MLrqGcEgzxbokl4I7/TTURXvFisLjWuBs0jh1ZsbgYepNlqp7
ZIGjDNXbsT86IGRgzLyJc7mR8Un+WtuNOKaX32LF51/REOenI/3oNKtJPwBc1vABx+9dZEUfHE4W
y003vN85Y+/+SLDtqmxVWM8hByFB1kw3an8Mff5O4FzDiFyD1wPYUsKT6zFcnMSEEz9HJQ1qMJOt
9eqRlLs0TUn8fBgvjr0VpUNiy5WpuSjcO4rIUq+FWZqRCIJb0GOgXfliLNVdN8C4wd6LEDvh05b3
i1hBAWT8fr5dptySkhF8b+qwNslNCNR+15LkxaCBJLdNgvKgY8K1QAT1ObtSKS5G1BZFFCaMQ0ph
dKdGgawgF3PBDR1hgYtjJmI323nYd5qoO78cjv4yIpa0ysOV63/+H7uUTM48n5FEGsfX1MjTX7Oj
dkd04URmzVOjsIeyaBkFTa1nzA1yBU/APQKwtuPchiybyfrHbfYPLH/47IRoytk80gVXM7LTO88X
PqhAU0+nAeK6EEmdLgezliS+kO1pW9b8tyhZO6VW94Xf5YTu2Chdj2QKTznFFyVU+XRDOdms9y0h
7bofXL64p46DLFtKcqarYAe3EtAkkoMTd21DLdAx9ooJd05Y7mTrxMLYzAI0lhATWWmgFl2xehpo
6WDYV2tVX2JSkY7xCD2MTG4Ffmfzc1bVk9CHjWU1T+7GIuL9I9s9Nz9zj3XDDwf1yLiS3dxsLBFt
wG3vyFfBC6yaJcucrEXRWnvfJDmneKzg8MtI+iV4epfRn36oGNYntLxazN15JmGxHTmPAa5AchlH
SjNH8CzPh8lOItZlrcxt/adYSYkNQABIAKdy13uSkWwZN+L53R2873rgLDlMxUs8OdU5EiABXcrM
hjxEtt5EeaCcnj3XSaQ+7Rzx9p3stzerJeZGqKZ8ZNTrKIvoAEnuSaLpWrmYR5mHyoKA1cE4qNxX
WgFfl6kjvQCilj9m3mUXRyttxBJogBk/2drmNhf9jFViri19jL47qMQBbJehnO4SixhS8Cqi2vAC
/Ykkj1q8hGlMNLQjSXeNbATSAAjO+2IPKRuzdNUccj8G7iVIehRbEbpTNePxSXgOH7AwxEyOYAEL
V6no5S1hw3JKTSVNxUwSYhFwvfbrqpCISJ6SgVXDcj0415uaF7o0V0wyu1bGuCk7EALCRyftyJfO
msI4UGoqTeo2kJBeV5OKziQpZ/UV52cYpAnsjAQbr+zRAA9Ejyhovf3wsayqGDuQR1GHwwL6j0TH
jR4NeJUFMiyqAa+sew24fqTkjy0lci/w6UThAc4UsACwVcX9c73qo7jRTVQJ7DbRue4Rf+84SA1q
pxlGV/ykazMGxuvYTliA2xlVPgvBe0cTSGthaXGRuWIVgm5Opid1RBTQxc5fICWyYTTdZytvn9a0
347qnOjYT9nQ+/KfYrMswRcWKATAI0M7IYXTHhzFUUkPvQ82Q+irTG1bcGxMErCCu+EgJezLfLTI
cqS/WwHlVqqMBjpkWr4nZg2YeQZhG/r3gBImdHx9WHmZ0Yah7o3CRTh0uT+0KFKTj9Ay7DeYGpto
wVFpcgf8+pIlYzxFQ3/e+JJQGZIE5akqNevMbHJX/skyJaS/kmB/jz80b0Va40j1EgiXhlpgJkjY
2lj5D5toiXcLXY4HaYELo+S2hUt2BZT4yRXjg9k8NLXy4D9Dx9QX8A0HpEpYiTwPOHr51A26K8z/
vpmKypZgGBuIdqyzBHbTGyJ3Al5gAfgWXqid8AawHDMLXhy8IPac4lx4V+F0hlbM6Itcc1XManU4
4I2NgAyRAEJdsznVt6aT/et++hcsdPfc83/+OlWKTwohoySDTK23amvl0nM4merprSrb0EoAFlP+
OtHZQ6DJC2haAMUYnqTNyw5h+34hMl6Oql2VD/YUzxX2jw9abpmmk6V5gEOClDF8LlTSQwCsU6cv
Z2eFuZBG6x30vZEIGo5vl+hJBJryuuv9mJBA2QL5ZoyPy0WCCPIKHH40LvahBHnPotghlWMCL7ra
+lK9rxKOZ3OTER9EtSvljaehGaqNXaBhmoxgyFRHDC/LhbgG1b1y0lYFvtYntBfnn0nnr7JGc6UN
faLyQVkMKUzX0EtcysSuCG0EofJopRqZLYgrkytmEUfKWqaaxxd/ezXnXdJUBiZpbFd5TnNdkEsn
nrPLy46q5JYVj4BoJoNNseJElAIln1cKsD/p1UfaYw/aNrD2yFa3Waq4sJybFxS5xryQgPS5V8dT
w4HEozV0bSwr0TvEAV46Ytd0KbsBBSffYgrrsu0BatBAkwKiVUZeeyJtWYj6PRbn/tV32loBzr5D
Wvd9C3j6hngUhvFzsaA2lPhCba0Qz8jgFcMBJvozCrJCfV5eu+jkFQfdHuFK3gM8Osf/KQcBuR+n
uvUH7NtoqAtE6YGjlAHmoTRFE+OLkE8Rz/unSFAou3QCMDOHDnuBbklQG4dgSsRqewGc5MP5OBoh
jZPgu2iBTALxr6y7DS3BhbLUBcq+P5u4hSY/4ihOtnlylCLEfY+YhXFcsfegUEqmG1L/u4nhvx+N
UVMQuh8BnqZjJulEF1WBR9nhRvQkbMYXpyT16HSruAOZNgMq4d06nUK6bWSSynwpJnMX6o41BtX3
xwAitsvTjXw8Eynfv4YzGpq5QrhQ3ckjgBJHrMD9zIJXH0DPxkrz5LtBXtusvgg4w0KQIGblOeN6
3lkCVKQ/+z3XJysYS2QhamDCNMe28cUPWg8yAPCDuKOuPRGQhYhGQEkWnHH9hUapcWEUAKWb2HyT
x7N+eU61k+UcQ8D8Om64YxEk6sT5dGH46EAVgSsSrrDNP4tNvaCnrlom3mCTed9D0dKTqHf4aAGq
0VsvnNw8qS/Je5tmSs9xGw7OfDbm0ZAN6myOvhNHlmiTKNMmkrpZcJWmMHhZ2kk5d+z1PJsSCXEM
IO0gzIeHlmGxhtBLlZMFijQRYDOHZf8/fwZ5TAyi0tT+qQlwr0La5GB77JwT2+WN0g20TYPVIKSs
UG9t6Q4jaGZCHodvLd4Do6+1vUATJ82y6uk0Dz/d/f+hPmpCMnQJ3B8+u6M57nRdLoCsPDVjhGeY
w/hzS6w1XzuokOYZPdj+Xhye2g2UgzvVOhR6Xmw8yWN5pGmWo3eG7L0ZdouLUnlWCcXVbkl1BVk0
j5hYgTIDPMzwQWmDcuGMGlvf8EZS21KT6OhXZKyrgni1oyTI3t9IuV8FIMN0vyu/BLNY9gQ4SPYK
XI6iVdYrvm5uGA/fvVngpPzmoUjiIw+IiaJ3ry7/P9pAfNY84NBCJf2fB2MMgpWqUBAp90r3XzJX
Hj3q7mwfEIB7z6gX3IdmFFhVDe6DCZb0EVsuYJiIFLq5JvD1vp4vBkllyaTZ+dyb4oCHQ2MbZBKr
oUAVniYotitLDboxIqQTanUnUC1HXH3qO121+4r3CfKa1Qc3OGqZ8GQj1pvkSv57J6+Mmz4IOM4v
yXvwriAWe0s6X3baUu4CvnUv8Kwg179zwPR/eQ6tgunN3g6TWesOa6d937ijvo672jNPF1eaaLsX
REj9tf/HDj1bV4XoXA2Bf5diOBhDnpQq8A5k0YlzSOtU4P+Vjn4bHUntsXs2IZeKC4Pp3516AWnz
/6peSqrcCJ/fscmTtsSt7TYBxZnCvCNeOmC8EUUGYA8BihoTgEAgA2IM6tr8mOZWFMRY14k+JSmi
/mAlWIs0+JAfrZPGJatGAsDDI/pRlpRKvsbkutMh2XLpWG47VXpOOE06hkxLhWngREZUzONWKzH8
qauP+Y7Sghz3Zn0qAZCQQZt3pNVzLAmwdbiSRGnunEbYdVvoFH4gkCcadeRsfoIT2hc8Dch+L08W
4UO3182JGnZiai0xfXgL+lFI3oQTR9NmcFzshVp9+FeBPGunK7BywmNL9UbW2w8l0qlbDzJDbDEP
ukOyX4x0M/H8MCoAdS7qoeI35lKuLm1TjfU5cQojeKF6taK2PMFkSPaYuVU8Zztb3I6UiOlKP1H5
JwHlRS2vssOToqjyLUoWHxFtiTfWz2b/YCy4YvWuIymB9NPoDC8iB0NDG6+h4jun1W/yIoNyYOOj
2/85wVb9o+ILwVpJSkyeZVEmYKMTmeoZ8HlHo717fRxs/SKVaaZ/rOe68BjXsY57zVTXstmxOsj+
Q3sBgfxvgQpmg/p5qiSUYGABD51CBegpMC9m9NtI0QYF18NMCzmo20Fk9UKQrBNjMEPQb7MloDxc
h13pstay9JFY1zOWoqL+LmovlgPh9ZHzSADOTrP7L8+EWI3SFPK7kPwjKsJbxENo4JERnqQtZ8z8
Xb5J8arNiAYqLazLyQYFki2c7ya59/9KR6STZUUMoQyjU/tFlYS75DBEfZ1MfOy9RHNWPuycFmmA
I2lEiANmX01wkyON/Z86SENOpdYLdEQDNBWN6+0Y5otVRNXOQwASkdUd0cegB1PEBun6Y0NHIIik
bUeOOoD7pBHSapzIFy/paFmUqixRaFIJBqcotJ+OcCllvVGb8+ea9n7BpJyFY3U1JSUGg0V1Jlh5
lY0ED6PhxRHbrtSenw7JlM51tuy+J72TUhn3N9WhULZUvVv9P5w9m/Rpd9W4RgwJd06kXJfujE/l
RvAqCpy8tjUN5UUQM++JjxYf+HWnx1r9bcfFR1FaZbLpTp2RtixEPQzuMe/XRsrsx2+TW578FXDa
CF0fvG9FMDyBcYjO6kyZwIx4wK1CAiHWNeSlp5uv6uHr37s2hWom3HnG1qjG9vyVJX2LmbVZmZF2
OA51KJl7oBy0yiyNw6YVx2t42M/up10TwIIguOfRBo+nrhDCbRNkMBGcpywDCFkekKXGWCQdclqi
gFlXYE8Pm8BaAZOlUg/lvQ6B0eZlmmAYCMCfCu6g1mpvn51psvEa4Z0as/0IwJNAO0O43HIDsznI
e1/7AeShrX+cHolxIrUJUY3B5Z6MGaAadmoJdMf18ja3IkBkK8Tq/63FLe6/N0F8DNVvRhjXI2wl
ymlciRbZJzH8FPVUDW+OBxz60YGo61lyWUYb2ONbu9z4q2GcJYNxekL+Hb+wCcw1dIsCPrbJsNRB
MEVjKyay5em5hWVLmtJ52kBvyPk9WT8Qmg+MMfeVSULAK04wg1qPJCBEWv3jNJoiJb/3oQoQjk6R
rP9jpPGY05Xj/vW1lY5LWHC11dPZbR/xAvLflfPdqeW6xdPicvesNOvc0UkXMq9ZTjAXL2Xuqp6V
7JPcAr46DmwgATux2/P2o6N7fxG7Ta0P/Peqc4Wg7CF9bgVPfnpROGpCiOPgb/VkZ9RuhMivUlVV
0iEv67PEnb7hY0p06Yj0qGe6rgi2Vy2z5zufSA1+81vT6x1Qt9/MxAsUy32N97HSAY11EynGE1OD
t7EbCOhWkTfbruzY+gDpNXW062hq8232l2wHlPlhN1JXEJI9DErzejFNrk7OLFkqQHs75+kEgXvn
OT+rSC9o1Ll1JvVirzPOmjTozKGHWBr13oSzSpw5CpdE0HU3hqI8GVeR3Pdnkzqzf6Wgg/u43za8
Whw0XBRF0yRKLeC37xvewq0UFZ/QM6uAKTLODn6GBtC+p3PcxGeW44KUUAowzAKT31pgmgeghi/F
JXwkBg+BGAL4gFc9Wf9DpUU6Bqobxkz7JJ7Ga8i6na6aO8593CERfDAXDcsWrfLJMLBGWJf3XwpG
dkMAdoy2n+qhA0I9viR8hU+vfro81ICfmj44f9x2o4S3j1ljnHZvlEMEh2iYKukdlCQEE1od+QIz
o+RvUhT1TsySiZLJlLHsMJGFqeMCqp8KfnR7IQUnoqpC7Ui5PxDD8SJVwq5aSxWy7PDUkWJqB31X
k3TM1k/PUuioYHzQjgcyXR4JMvJxmkkeuxXs2FRMFd45sUw1MVr4kKEEjxt0D9ZE+VqJCd1CnxyI
q199mqgVMcNTZsRw/M7nZzWL2NqW8hskMV+neoqFYFhaIy02XajshDBVWnXf16JJPtOayhuFmTPz
Rx4yMXbx42c+iphUmnHfy5R9yz/8pQC4qVDI5vUAL0xdH5grPLHvqwXz9s0vsyYY0R/eNOaXWj/d
8VN1XknBvYE+UV50J2mJbkLAtVEBximaEZzI8tL3/oaCq6eGItWgnwfqZg4gsPlpuIuE4wMUVsXu
ZJiXJlyGMnM3/iIcR3PXbfEEDjWeZuOQ6tx5aqYle4ImMGiDjpLCRy0YcNyBF7mLG4iGKxXrxl6S
CADc7+KdUXuM5n48yrsf3LJLVvFexgMZAY/1KRz6FA8hVviLLffRVozIQqyVitoGaXt0tNruipwa
QGH1b5rOmB+ZlNv7lWJ5pR9YVeiULlokf3l+5w2rWYjEASl5SFdmwj3sC48ihhsmocPswi1TF3q8
tBmY0DhYe27bj6AbAXCZYrhYP50rp9suPFzD109AQ1R7us4j76FceliaGUSE16H/MD+ysCXMl6WD
Hz1M+A8BP2r/Yt9zJ5BT5sq/oAfNWJkUPnkF8bqXN9Id/h38qrR8VN8QKvExxpKthgdv9r9IgSCi
glwWR3O3luEJMGqadC1dG8+kPYDQJLuFUvOhVCUpR5lolkRIOqSi4KXKdKNtlIAL5ojQRLKyySal
ozSC/bPzp7Z1nz00NzMEEQI9lOFh+48briN1xOtKeeL7JwneJN7wFqZSQr8VUpKRAUI1y2b5HFXW
ytFEVhYfVcqBD8JaY2bKaw7IpEUigCtPsj74ixQEzF7L1u9uiF99NgdEGjlXOQamZeaMhX/xSSkE
orf/0MKZmoDMkj45qdXajR3zsF1B9eX1/hk2iE2DlDJ7R5b+N7980eeQ9q1TqJtxgDxMx1oG0XzN
HxoCvjus16Ktv4A0N5yjfSCVHmzgG6bVNbjZqFN0xNDUA6uG1xIdjqyrQ0AuH88da6qOsUBe3DLK
2HFM23fa6HZVi1GpkgNEVWJJZ5xsqQrvGqVkJu2PAtkYG4WntTXeMO7rz8WWvc3bfPgYeLT/6VoM
eDN+UqTEYE9Baq+Js/5h0A4m1DK5zNIjXoxnmFvPzHS81k+k//pVLHcPXr4WS2NZzNgPPGakLqnZ
7Hs4K/eqpZ5wZUD0q1b9yTgTob1IX3qyS4/9CdGysiCVfMKUZ2P5GnNa2vB15Aq9veMW1rLh60Mo
x+oTlcYbAo0fjxWf8sZJ9MqRtGGozCeLypV8avdJoTRdwTaGhd6Ts+RbBou+eEWFk1omo17XvGe9
DoHX/WDFujK2XZ+2lMMwbk3BYNzZpU0QJMQi/ulC1ws2pdPwoRASMhNg8FTjrJenCulfYdLcmcBw
M4W48Wuk5kFTPLtULdgxEfWEAbmLJzJmz8h/EuCVt4T3+5oO7MctMmSGvRCNaSupNR6Cg8b50Yuj
LSXxsN2v6cIsLsHHllnvXmpqHafzBQ/kva8dXFQlSN/L4Rwf6dRRrzHlbvKOOPxM9HU9OvqR+Ike
ziQYiNwmJyYpAQBt8+5dSYOncQw1UEVobzStb5o8WibOiKXX93Rqx/XhlWdq1sY0Yw2+yDCCRmP6
nX+YiRRnlKKJNyrLP3etCtCkY2ZdKnTP8W13jTE5STeD5SOtw6LsGHlLZ8NFJB1oZVugnGadWHzR
z84K6+uX5Ns97LX22AGrMAlcaSiJqQUyxrIbyot6vr7vD2+OahXojlgDpOh2rFtAVWXuZL5WLIbS
7DHSmiNsNPpdM5OXweaiCnrEMmF3IrmYsNAzmfxcJvSZGDR6HX4/QthU84qR6mwiwW2adoGFr6G5
otRGIoOjjPkPp13BPYRIul6LORu9i4oMmbpbG7BxY2waUSuPT2m4i7S7e4POOR1OI7Kg5doC/8Ik
XJfrCa0nSlleS5fQRwS3+cpe3w+bIWOK+97Wvzn8YMvcGo5aTMhqPXlhl2efZZ9QqG6ra3s8c994
pI5GTYpPBjMAh+KLmtVP9aRFSBdB+SGidp8hqmSKKUj3NxDktwROi/+T2QQuchOkE2YCN72JcpSI
UvlEGGm4wCzQW/v3x4vC8UMOgK0pkNHZDT4xYl8ULT0qeYYBlcCkSf4mM3pRVTZ6AgpZPvKJN2RX
8MY4AkRHjiDOI51TcLtxYxg2a9zNUH0YXAT/BHqpQFrEFAF2s6IzvvRs/ORlYOYb4wBj9ybKKZXj
aTji5xPF/dIPHKhT8m1i8wtam9R74vfH95t3jbI6wzGFucptTaiWp0gSuPb4COiwiYVtG74dZf/Z
FfwuYEuaXszzWtcIj9KRwvQWn82SLKyw9co/vwzYwWohtrkIu7E05JMIfRSRvq1c7KMihbtef7yM
zLqW/JowDn3E9qEA+Y8Tb/v/suVmNWyikqSuNFU684NMK8dY4sfWcN+65lV0h4wGSn2U6C9qQClg
lCxaXkHoSfx+C1Q2coDamBiiWHJ/7n3QBrGIfRTQqPR3DcnkG1PQ8lHx9vX4ZKga83xCYBdiUkin
qvqYRlZS+YYEBfITonfb3lhXhd7sKnXLLzELAxabX9OnloZXkrAd6x2jai0sL+NA+OnVUMVFop9g
BM8eR4cj1wxnYqMFk2u9QiMAwBx+IcfdJ6M9CSAba+6YjDPR5y9O6Cl80k5yOzcRE1W3POhyI4lC
0s2eGQmzGpEy1Crgcqq6wJs2CQIiQp/D/mBFpSXb5y5Ddj7pas/NHaFS/v2iLn4vscPFTAC/KKyI
INe002r3pCiKoWrAPI5lw7+IMLZZjbwqSBpuFORrEm5vxqvcEmdoy9y/F7HycOMhbySwmVYoi00H
orRzr9FYEc2zqvvJXFB7k1Bd9CNt8K9F6BqECMSdkn1LNOZf04DpTy7EiMKlOZZkB2BLEuftUymB
PkgW92X9rRbE1bRcxmKa+6iDdGnMxEmHdPmE6NvfK5XCsd/+FHnL+OLNsBSFkcgxQFh0ox+zTDeh
TXCOn8Yck8mw+ISx+1i1WGAd4yzFeYdh7RqDubqkXFg2hiznWg1AA3CwmY9yIzmSnaRXkElURwkc
cKnQHL1taHa5Sft2FLnNqGBZUIVWa4Yb6AJEnI1tVzCjo/pET+YxIguEzh/rV2X1rJKqwFa9ZI/N
zWPKrJPFcE1nVo/Qgs4GhCHBWQ53+EERi9xxJgDomfcSG1ue77u6c9un3D/m5jBfLAbxF1vfafDP
fzmM+a/cuXupuROLqEUOeckFs6nnUOonP3wYbt+vg6BukykYEVSFA6WhPM3vbQbmNmEcLgQeJg15
dMAZEAFyBGs+0r683erJP9xWr/yD9mVOBOg9ui9wo/JRpKTbYJH8ndV8JrX8HhZe3BBeqsE9u2CV
m62kFAKyZI3N1VcqqdqSCTTqsRyvqbV2ggLTKjo9Oasfy9wbNeD3Q4/Z9vAmGgjdy2eeQEvfnpOi
2svgiyFOOX+47YyIBLorOKDIcmoqOFkn4JOSszGd3rEtn2H3IB5l4Ebqaw/YLRtRsVnsJCZZI50A
neEt3jBIRqFvevA6ojnTesxRsLzcNmlZMjPvZfJMJfUxsqW/dc5+TTMVje1T5fLEssdVWBqmrUx+
/YPf7tMOZ2vQxHSFN3FIGAknmOL8ntU5i0QyUgWhVPelV0c/svPrIvYv54Yn1v/wNbxS6aBrtLPh
QKrEjL+ddNumvd6PAE32q7dJtKnaj+DKlVxJLfV48VI21wo/VsZuwySaWXeJOLHL8tRVsdBeiC2r
BRLoU/wCIi4JzbORFN8NcRbwE9lUOnoOV+bPBTXIYN3sWvcPnoiVuSjgxpGm5ynB8aae82d8fQbw
WLRkLmAfuO7HBmr+ehLinE8zD2ymP2XuBpHK8QZtHdfdUeI9M4SZD+3/EAhRtnvpXOKj1FQt+50/
st4sB84cWZ8JdG84y/llybl0319l2xenLlyFQcq+8gVQlSjy8YH4gQkvW19JD+mxYuksKpfOIgo9
zwScrH1wyvCAhpMkIEz6UN98w3k4BxtBYJQalgNs7Yr5gfDsiVb8/wmsD16MBksGRkSRSBRBFqos
dXGKl5V2azXvzpt68TD6eyhJTcMBZY5w6PMeLAk2ZkbyzE55BhnkEm0DecyJdo6mgGAZ13vJci1a
glwuEM3+RBRnKqLX06/8KA2NXV0WF7R+9oUQQ+NgZKHz5eDmDSYaAMxDFRn+YCwc6/nDm3wM59LX
x3qRkDEgZQNLjvSI3rqSMQgCsMDW9xFnrTn+5HYu1zZLFzZU5Pxxd21R1hHBhbpPIfyEzbD1rlgK
ZWISgE+9VTIliWAhweujp0Us7I8NAinl/oRql6rA2qNKCg9JgkM4wWlZMrsq6kwyCZ28VkWRsz4n
HORT6j1f9h0pHxMRTlc6tRwO8IQlXWlI3IBkcLahEIAdNteTwfXrv7xkpkbhbnb/McZFFC14Guyu
K8J1P1JJdxPdWvI1q1ehH+epiYnqdjmyeaMVThLuVOWfo8rW1GhqadXKGPbbc0xEjYjxxSbgEUle
SfH0N8sc9XB7AsS5TdoioTSU/uqyLo8W6m0WTNxN8xHbgSeSbVravk5b9fHrqGVJpsfXhS1CEgo5
BxxEZzHVxiEFpcDg31Z+8oGlZ/evyOSJVC4xNlIT4jTKRrZgm2vqII0wN1gvmah2NzfQ8Sou1WWP
gRuKtrtJck0AaTuwfU30Jq0hJg9DXlW6s9+UIClaDbxPWFWJxfnDE4dyvkSxb42iRoAjPAASmXYh
4SZgujJy5yeo4V3PW4mqhz8wJwjGWElHldH3MjNkdFD/95rAxqzC/armUE5e0/70HeC56365XY8N
FE9EBue88NGyVkMjU7rMDjNNnMsE3+tn5Q/J1d1TTrakZ4eEyG0R5Vp8AGgvzaUinLn2bHWWGv48
jLTIGEqHmebfdYtEFdJz8mVJ8TiqMzA4lCIO6XU/YLF3eQaS4c5EybiqJS4hX+qCVjVkVG5DkrXp
qk0xMpd2AlUB64hhksFVlGdCxq4uP3j3srOMpTUKcWjJLA1j9mmHAuDJe/qiBhhq+tHJ5+EfL9ho
5DhE6ulnjTpJfOCIN6k6TSIVTpSpjWgSvP8VwwEQl+4MYSGiP5i1LylwuH/pcCxNXNzl5pKb1I46
B4bnPOmcD9dC0j/trOg4suVCyh1tiOcOuiyjfW0mBcrb5zpt0ecH6wekvSLpMZrdgh/xXk6cSdHX
4p57Ikdg4iju5THDS2/j+8MQdLW5xGPNjE4K6KBmY67FZm9BARrIkddowBqik6SbbSAWWVqSquaK
VPDb8uzIW44fKKWssUefzJAJTnmm+hh5BkpOebBphLpXW8tYvmTO706hzOvi2Ou0yH7HrT4JgwU6
4BQAqr3xQaPl75LLdhD2IzUVB8REK4xPO+3afx2rTpJgDsk7vIKaQpuEPsPsmRenm6oqtzH/K4LX
aQrMS8v1IkNM2Hfwr46RchhwJ8eK+WYzwreFP9ylj7KVhTmYA9N1z+PKDptjEkcznA+HJP1zIGOT
SLaGrXDG++BJCdj8G2R5mPHYJmSLGOP9P4/yuxgpP7+tKf31JzYJMUHMBLu3Jgf0IqsoFVxFAQVx
kaask5cyuY1VilMNRtvUEt4JGJkWbwFvGfcKwMiFze1kRC4sLJhBfl0tH22WGroVn5LErB7LpK+C
qeo97SVgwBBwRqqDuIWH44sVq0UXAc8sbjm+iwRhlZJf0HdeVUqddZVqmEUi6YTbCG6ot1LXKe8q
3F82GAVTu7lTDF1bL/sjS+ITaAJoN5X0ck2Ia2KRiNynXvYupBJsUlQ2/rUrO21ynCUrRAs2abgf
M2jrnh9ZMRPM5bz7kAK5Ae6BDQedby23XVbzIHByNhSAP1n8WD0cJ3YUptGJ7vaAoZFep1WztbQM
an89qhhnA9zKfmdR3Wx3CVsVjC/tItLWHdLPkxKOFnvPEOmW6qdpvAvmXHav698OItbVJuN6nblJ
p2UvOhPLmuK2L3hzkcpnN12Zj714++9t2jgsglN2epVPsC5CNhAKvrAfhJscP66nQ8fTAKM/L41J
da0ltYVBEJ5dJnWhaE+5iqzyEcbL3U2YVH/4Gs997/4RputZGvOuWg7UW1q/+US0jP0j0K5iScrM
n8le42PGBlCtrCd5HNfKSgviO+T/TyUMbgcVX6SWM4ZRvrZP3CxO6vz0m8hjMuc6L1J8OBVAqm6h
1DEpDekMGMWXYrYOEv6iiflrGTdW+VuxZMqh+IsgCzPzvCRDfSqUrAxkyPEYwKCiIwnsJUI+/Shp
IqX5lfvZrVWcg0LvfYtqGdMXiXMNb3cvryfd802ytYyXf40/BnkXO+2LOt4xxxPxv7fExBBY2gcP
ov4Yu4pp7PV/Sk6X94T8i52JB4HS9Gchp5+wOOdSR/J1KFpbKvRVUtqytJ1e179eLkWHdUevS6/4
1eyBsGPjKs3f9la4Jliq+7W3zKTajAojwBOlfAk97LzNj6Eb0MqW7adGJWgFSaMQnCt93P0wpu8U
Uu9rsr4LS05Y6tRmwnKhn3xBjbcQ3Wx7VbMasIV+SxskSz1WStQjfgtY5UxstytBr98Ff74QATKT
Bu19AiiC/QW03t9IYEw78uCHpPh6CJuTckmkpaj4x4l435jcIiQY/ZRVPjvG/2OLv4EjNDmmedqr
kAaDw2KD/B0cOWjwzZWgxzSuztr2/sg7jGD7Zg93hBMrUWKGWvfc+oUB8RH7v1Rs9ibIBDAN65Fu
acSavF4Bud0w7z/oJKNZwWPMaCSYURhFI/sjWY1aZx32/LHElfZg5cnziAP2NmEf/n1WOvaIEM2Y
q5LTyKaMoag2p7tGu/v5hPj9N43MRBRPpzBHZ62LwoySgf0ME1/U8LHpIoCwMXQoJLqQLH8/N49E
1Y1uONJ0YAjoM0FxjYcxrQidgeLNfKljxJMOEUFJ13ZTk8icodexidqnmEd8CXNDDQkYUNCy3Ak0
LsvYGMWPwYAaUXRHFaws/8LusSqtLmKQWNOjtdvcEBmgZZ+6x+lxEMkNw5A09lzsshB/Jt4Hy5Ud
ryZJZZPa/BRz7A7HxsdSaKRooy/3/u7mxbRBmAG+XpbZkENNZ0TddcoFCpp+hpPcRCmlTUXdGoSA
2Nk0qzB2JM3qQMqtJ1aXre/g6k6GYYrhR7+WtNX4GZ3IIRN5pavjzFaXiiauurqnVg6sEFBzrbN1
3EJDESmcaZ8mRiHZbnCjeay1AsG7Ul66ZD9L8n9Ktrvpuqhr9IypsDGWFzP2N6yCk11gcfnOgHvf
dc8B8WMSuFHD8NwTSoGBhquuOPoVDwcVEf9J5GuhbOC/JmQeG2RzeVD8Qa+uohbzR2QxdpBJTu/O
iNCtcKVm20Y3Ubq6sIOVACnyqxYXoXmqUas1+5waKsj91kXiYQbGgR0PBwToy16slJeJW5P8ZStn
is4ORpTYYY933F/T3EGypfExpO1cZuJP3Tq0R7Y/hrG67XHwdKaSERjnNkagDVGKisxVESpqz3rL
QVI0fSyMo2UwWH6zWfVYrElOcb4gJ6e/YBA7SoO6PTE+/ycc9H+kSaamJXI3J+qJ/WclvHWbfGnP
vh8ivkoZMMB6fGj7ggfkXPWwbMFJzMADAGNcvlRgLQe3bQ0pICpC26Qm0NW6/oHr+OqWhk+1wI+K
LBZEcfBR2B47f43VF8MhFBgTmkAknTMe0//5rgkObOvm9DxtvAMYpIWO0LrTMXIrAJNSz/PFku8M
b4MzMUhick7IoLB03iqKfZkkDjgZxAJdmeIq6wS2xxrZs2tcOjM6ofcjxGEkZIO8rJqdGDhLzxbo
e2pbLyYR9l6l8M7xK3kE4fO9q3QNOAJUiE437uOOY1DbaVxQ4ZOY7swVr7uqGnPWVCBEyvKm0MQZ
b7Si9cZj7Aj4BmrwQBJ6LH3ydG/FmYt3FBAfo0u9MYAeBiNG60bdIveCyeEj0ERBYGlfQaHUC3Dv
GthRc3RtPINRhnDLu8mIAMh4b8AZFeB0K8b6ubtUdQGtJCa/AxF+8uHV0r6dRWf1sONvqZM9/800
RxrU6v3gxIDBs9lNSxWMSVpx0P25CtG2mWmsCxRwwXh2UnUICOOHhETBMZsD5R8U7yaoKXK1TKmC
eiMX6N1rVnbGVVF5V/WD4OcZVVQSsokn9zJdhBqxAGDU+mZ6AYI0Oed6dUaRHlhMMmfYnUwkQw21
aYjS1Pw4mAaQDpvq8m1hGHilLUpUlFkFnKFwtA2mviB+8xLhW7LcrPBHd9jGrD57SCxaOGRC0+sx
CWbHMxfxZqQ0P7l+cXxYmXvY9u11iQ2k3E5HQo6oIyYUqY4kP0ywqgcqE4gqbZf7P2aaK7mz96vO
O1Oe4Rofqmp0/rZtFVXatD21Fx9ZbSvRO0ETJPIGa2f1nyHKP0YDLHf5cIocxCERR6GVTBi6krCj
jjFXHPSAE0WG/jB1r+Z05DaIm1QjawLksWiMKR7hxRNEhMzBlXYxyIK/K85Z3VTCejqmYQqYLvTO
5nusKpQhSzejdDPVsSiDyVG8QuoppaYqUdPmgshtaJde2/bKnH2ZLDfxtfXPqiUtlHEegeZXnnks
3IFDJhFiryGTdv6ZgnhfsdpHpcPhk8jctcWhINyPYgEmu/AZpX2YKM3y6mRdvbQqjrr2jlZBKUFg
xIKX702+cAUr1EHW6h1RvTc7aIgDA6D68+GlxfRbaYPTWWCKVnXG1e0RHyiLTcpkLFlLLwl0V8QJ
7vpb0GQOUsgfrWtw4E9XtpnxlYpVM5HuEn554NZ5F/1etOKGouByDpD6f9OdWOD51iRWA975Rny+
vq57VkpfBUYMZcsDQfcz4SOzZcNJWWkHTCUyjbQuS3h3grMdDPcM12i5Ikg4+It7G84GkL66irX5
WjlfA1x2VcIur7R8lkyaAk9E2i5Wj/h/beyUVgI/y8bXasaXqDYCA0a5vXekMCMQq/kPlJAMt7i+
1bXFibeWZKX7mIRQxp0Rvp5Xuqg7I1//4ydGhbe9py48K1t+yn35dNUs2Npvo+TiU9gVAaGDqUdc
1pNPydCWS6rQ7jMro3I/Yc/p97EusovOfAlWJpeMxM8ma5xTQxhIHzZqCwR6tp9s8ILBZdzmCuCg
wByrJIlIM8jas6FdStrmJG4Yb+Je+OBU40PSIhiOKq26riWPhHLOc9r54MOvo/3ZkVIkSk9tdNk/
AqiFgZ3mdqkkc6m/LHkfJ4lapVcrJXkjy+cZYxOI8Dwtcd13ICLZP9u73ZsINCKT80t8zTHYfkV9
tkQFbcEPK+c8n0leSetFt8Ze6Z3aUnDU6Q5Focp+f8pA0U/C3TPLYLlfAlo/9Y0YkwM7rm3ZQ1/G
xSdepRVNNSFVz2uStQmzlBt+a+2lpou/fbhoSHi59zvCi2F560p4NLVqS4KkMeh40hEuvdFv5PG2
ykwaU2vbe695mh83m4usswRPjG/Z51wR9bLbDnMq/E1fI/7anxEkA7A53rJAOTW/Maj3nYM8nxwe
jdijPakoEp7PtbaEjOq+H6B8oaqTqcSL4z01G/E0ZuUDV9JJyiNAJMVcsHZLE3CjTmoGkEVQn0Qc
+mvupfL6SjzDtec4/mzD601b7s2/uOL2+MUQgbV/dzMiKJI4Bb08LbpacODJGeg0axf6x5M0eowv
fTQvvAV5rwLP5wFcFn5rVAUHtO8ptuyP1cjUUZfaM7tLueo9+afP/M/3ZjcgQF9BCWSlm7lEVhlq
/uhsRmhssgbCtO4YyO5AuWsmVB/qlyQ5Ai/C21uGzv5ggdy5htCZDlbkab3ENJ2u7BS2xZHVb+fl
uuIQmn3pZqNOLV8DlGgnpu6kfN6IbysjPsXlazZW4Kn3xWJtSJKSaI99tQgEwYOt8h3E8gSLLUfp
2VBPzkV/Hr6GG5UHHAJstKvn3GZjPO/q18VkPJILqDyvj3rYHnCjn36IDYEX8w/le8uWkTfS8rM7
6NavAJifO7AL7F7FUj+xHM15p6AT9GiEoVSUMr7HajRCA03Eug9pK+79v0Wi7u+RcsM4emZMNDHT
QzlLJxBU48dEXULDHFTq2+sGUX2Qab6XH8F8ZkaKoQ9H2YlHPchgrhpi+8ul1Se4HclsDdysCetU
vS6d4JrD7jVortCwLthbTIjD/AFgg4AeHEY3MS/aNkZdj6A1igEtQ9J9SMSjU6REb0lH4+b3lZNz
TtFTpMTATGKyawNZP0BriULpQEmraI20rvGoTuKZrrGa4M5gZ2O1rIn6d73mnccdZfqiyOpF/lZG
Fm07m8Dxb6gUr0Ga3vQS+QgN5aVeJqdf1nTDtfXA6uItIbuMy/BAsuNtEEjtFnBy9gPoW+RhOaZH
Kyr4OD+FnNpRhoMrZ5ExvmgJy8Dis5XK7epup2M08Ti9tMbkBamyzoVWBs3Ae2tXp8oyo7vvIUDY
oAGegrML2FMtOq/SKL+NA3yvVeaeR19A8JTVhE5yBnK+3XC3zZS8bNXM1O5+ZbsNj7hJodHQJIh2
uDkFnZEOLfgKavfTTu4rma4HpGrkTpyiH6cXcso6PK3HRlGzP+ICmz/Fkyt4uLPZeKXOQsE6aAey
TFH3oRjSMhsbud0d5bLauMmZgOiWqcVx+A/vfJwBhZ8GxC9M+E7KBKx/GgrDKIhpXU3UBJ/Lsgpz
0NOHYEcI/JN1hBSIP6FnYLC8SHOHW+Ob75uZDku+3m5iiQ76xBgsxL1SlhZ+gb6M7uv1mznisl4R
7V0XBN+HR6tB7J09u0mJ3So2ye+osRbxd8jMvF/tVoMmTTUhHAuKZ/g5ys6PptHYiuYVcD4eUeqP
rAgV0USl1NBbuqUffJgP1Q0yHRbLazGtVWoRyvdXE6XRJ/Od3QDtyZoM5/SSTuc85Yf3ZaJDk4A3
IrOMHfZHFQQtoGsZ+t2UDmqZdq0sdnhoijFAi0AJTzu2Zfjrv94HxBLxxjR7fJp8XjrWLXd9XNO4
FBprw/UAyH8ZARYspguRwFw2/WaD7blPnzrSN68oOgHsHLNwKMZgR5BvKDCpRxX9ec5riQBk8Rgi
lCmNxM5267KZ722vWJU8q/DToHmNBZ/qWmJgY14fKQRBnePiHN/sM9NiK8LnbuxnB5xIkrCprI6v
9xEeEE0CsPzRxUCGl/N8clrPVAWx1GRlXWCFJfeQy/qH8sOor23UkEoepska5uW62lxXx6/ylsOQ
H7zlDqRoxYtgPFTnyV79MuyaoFWw5K+988oTnhHjKZZww378RgfAahcw4nh28Lr0cOOU+v7m74+Q
hmH6fA+0J4yqSQ5G9mHVlB/APpw+YK3J+AxVTvHnR8UvbVmh+COw6iZPrP75ttjiEKw2azNjfnIi
m6m81QQjQTHsAXhtrZEj64ZlYJ944F73/ooHJtzRONS5cfn322G1w8txnFRGWGDkbnps35au4EgT
VFJcaSe99kPfpaxDzpXBW8LWUFG3UMd32+Zlkp48tKgWXyTho7VZ+elsWLAqUSYpn8WEFQbcyXh9
X9PWDRUq80dmOYqcvIl9EQfkS9SfCCDkBlV3MIY3CUKVMCs+0B+s/S932vE+sIn205cKIt3ThC2O
kJ7B9qP90mqU/wuBUuhU4k92HyB3szzwS6gCVfKwfX2ZmR/aHthysp2sKXNoZEC8MZgXO3mqOU9H
ivmgGA9G79pMpUHGZ74+RdMfTLx6CE9uyH/hug3tdD3wlOnSF3N1EJ/Qjk58lkFDPIilc+A6bLxP
6MGDiXdZ+CwrsYtcincOSvlDOefrBE3v1REJ7IPhAMPKUDqUpFv/scIa0y+miy4har+wONMQKnvY
+rz4iR+/Fs+8Tb8eNLUAp59rQ6QnLOeiRXbqpRoKYT9knaCYTieUORfJ+F1asSJCjzLEbfgDj8lO
HUKkWtzUmPdGF6XKls+OBQy+bWkdxPpLqqYRQ+qfPGKIon6qCbhg0Vyz5psnSnb6zN5PVyifNzHt
3TSqoTrgNs3R2Ygcy6BQg1EsqEX00D1d6C+mRoJMfdHx/4fpo49hgW8wAWMg7Ax9golLuh6/QsPc
J/QdXtsG8YVqnhivd1j0MKvElKICLIzN163qpM29v85sUczD2h7CBqJzR/kNSsWGDvHNYor64nYa
TnAom9iPoH2AxeL9OC3bd90ikjRnKSLEJc5dDfpgJA2sJ1rgf4e85XJFXwOCxDCERO9JgiJb9iiK
AJUALUsHse2u2px+JX4kjlhqR7Dx2yO9VhHlIXfzi3T/notI/JvdeLWUjYOd78fiXEEwIABWkZGz
UJWQPe+LeQKX1qvSXtrBm0LTUdCFDbWlSkdYZsIB/0oS8YpW45bzG5spxZUFLNiQcUGPe/lMke8U
rFzj2V6I9YBgppXMFGQrkiO1W9j6OPcIupcmk6oQyNr2agBtnAciBO1GQaj0G9tqoJMwGnj3gSWb
y57gtmCGHqDtyDnuMO7AVVLVqxZmR8hNNnN8w5WsmGHsYBaYFg2fP9Otcd30AWPwU4bPcwki2nrp
i9OEl2Wv5YdbDLfPNSUySxuNfk2VTmx6fVCRWqpceKrje+JTvzcUK/hd8V4Q9lU9XPbk813Oy6//
Mhh9gojfj8niZF0IIUT3QQB7cGxq4pE4T46SA28pg2SS3tHN3LgBs6OhaXN3pqQXHV/16/vTj8Bs
RFHD4OPg2uNRG8rJRgSoI5e3H05EQcUu5/jLi0WwHuGCwODabndelVfCbY78tO+FAqM6e8JkBRP5
Iejg27tbr792nt6HAAbgN57vc8HNOKQPUGRJBZTTbJ3EwHmMq02gzZPrUcYRCTUuHGzwHAHhe2X4
1Ad0+fHBJWwV0hwTabVPXuKfxFstopEeTz4Me/zWGKKWtA2VXj2SbuNj5c6nXRF6em5kOuvlLPWr
NI45o2r3mU9/gJcsriq6PmoNikcZF46Tt2EJXbQ0vKHizKW/kUqXE3uOTihCOECKC+f1eUldISDA
0cbl6DTS4Be7kf/EpC5JYfArRkzWL+obuseec0xV1PVZB68qiyIS14rO9w0+aKCl5bFjUxGg14H+
xuNj2IXfGKP/8h24wVs4T1VezfcjPaAumjaPUXfxHVHoDT4rZttH0K5kqFHHN0DDs1vH5uF8Pjd/
XRL2rOFioli0BPBhW7pqHzZ8Z1btnO3PJrKOXl/X3eqgV10MJBjRvo1NYw4w2O0nhUgQCwMRWp02
UJQt56GDqYYu8aANh8YNbIVQ53GNMdlrq4hIGF0RrPjCwMk94XMZXkUHmilDuzgXjK7kpmwVCNAo
lhg5AmsGxWIeVRBehLLe+KRS/9ZxPDOCPQnYHyxOJ8by1WLHZUuwLpgePH5dgdjyNUAp4UlP2W4l
23o+GybV3Ts1GR0uylt62iY+Uzsw8E4pSm/m8RQRb4Z2ldUvMRKx67EiA5BD/isbKalrakAPIH0S
megh5XY0vOf7BtGOKFUwnJvUnT6aHcxUY2SgUWVpZTCC9XrrDTKpFD++eBDfaGzfKvDK3uSstUSa
tp9tsCLxym2OAC4P2d/iSgTT8Xmrpt5dim3kaWEkb9GW01c+XhCHE7k9W1b+2xePaL1s4UBnbAOQ
HAGXJVEIY0sN8IAS6olb0zoohdtRQSIl076mo6pAJcqYQDfw4qJBTLvG0n2UZxHeA+XvfOeXbAaO
ZhRzZ4yVWZRgPefa3RINeUVUrOGUyevd+h95dS7u8+LdPMGtlZvuiCptNqCHCguqdZd/GYpCOpbI
rGB6CEGfukO7csamoZa1dsqnrjv3vOWJkL0ZwqaYGzo0ZANoOZJ+rLMShrSNQmo3GyZnhiqiaqfn
E853m+5muZE+md1E9WEmhqTErDjAnclP/W0otqmuFdQeVfVD8rx2P7VKrKlH2wdlKua3bKkPWBgh
7jR+gIvQHfdNsgXIIor14/k8FGBXzBlJ8UZ6bSTVmm5zki3xhYVrMrYUQB6W9FwKjlo5rmaSUak7
8OzNq4sDnzSHyjavQV/oDAHgLyDmCuqWRyHc9ymWOs8vn+6TonpK1BKB9zcxA7Hv/rIdfjKXC6lF
GCGkS1Y3w0+RA+OhsxhMHP9QD9HMNiMZo72MqXFGQ9K5Q3n8TERyPi5ZDHuoXJwTBd6IxadpvAT4
ZKtX6QBFrck7J5TNW5GS5Si4wuAeB6I7Y7f8E38WyiKdGteC8cJIdLHlMKZnGmILajBSUDJI6f8c
6nhV6WaZsWRtQl5cQ6CToRXUlQ66et6mC/TM2BYUWnXmTPB2HixFxzn7nICmDKe7LlVoi9fcPlGL
T5xLMb5v63NHWjRmc73ROQ+xgK71bg0WymAPoLYwltaC5dXudAxKkLxWS9NHHq7EVXvn4P1nBegm
DnRevE/ZJ6nd8Qj+KS5ODdac3YKGLPV0bXUXycgfsSjxslW26DkRgDs/TVAiYJ75w3BAX+MSR9y1
4Ih72N3CiR37T4bze6hA2C4exEg6JgVjHhyMSuhdp9CxJK+xnAaBCVeHMvVXmqN5GX+p4w7rcKXg
kTmOBj92Ifl1a/eAFNqO6hYheaXL4Fa22Sbjd48bfcqJH4+vESt4oyD142mApVHx9ot+2tiaZS0B
mZJogj1GmjlZqbA+u3gUZoX1IHw5mTridpCqGYSosg4oU9ALTYLoYzrncGnPLsWRfr+URCafBjY6
xhwPNKFIsRlYgf9D3MPQRDVLVYaNrFwjwtBd8PqA/ucwd5R+UMQAUGMorC7/Wk+q9k2vW0hIGxMj
mcXs1sLkzIBsU2KJP1EVcS6+gUs8UfWLRYYvozKzFQya0u0AKbFgZl5uD139jMRiOW+yix5ATuTH
uiCAepLkUthxw3A1Y+gHT5+eEd0/uanQbSDjfDQrQi+CzqPLOEcNMJmQvs00K9caebHlele2xGjW
StsNRyAFOEuNIdDdGgajj5t8m+oJ8rlF7BJkyQVmXv0mP/2iOfAXuJEaq5DNaYQ7DgpI7p4bBk+4
JBa7epNm10C11HK2kqKlxuqfhk/alCiG2eefhg8NR63rdarVluWMHE1CP6lXX5BiI7NRvVV31qog
L9vfQXglAQ1kvddfVlrUgSV8/zqN4Geq/uHeQ9ZhyXcWTylZn4n+CXOOK9EWoZgpgQnX2QmjgUHj
N3aNK0B8iRbNuZh5k12hvuN7Vf63WRe2WczUA3mcJqi/tYPogj3JAaf5ya0nJeK58C5WquaB1Wvb
MtUd5+qjFUtnfJNea5zJCPLaHkCXscy+bWWA3Qwyv3XO2INbHX3D9Q5RHiVll7WILprwG45OiqHy
8Jo0E3p7Pyb/e022+oWVd3f9iNRiOS481KzAYJuTY0lxh4RLtrPBj9VPTijySOmZSKGYgVKkZU4e
SXHjWu5kglpOD8STrYu7+yjtp0+SC+OMk55Ajw6HLzZWsv5gWsuTWz6JYivkE1D6PZDdlVoiDvNp
YGRTjta1shzc1vtCWqfUZh9vhF9gLAteAEHf9XJkUafNNdPEu0Qx7uy0wjqQ06q0mggYWGgRiIuc
LUt28YZufQOevkmzmcDYme3P5tHyc4zznbfKIFneY8wKCkBlv2+MSBrYpfrkvXSSAmroqJBOh/ZR
FACBBRzUiYie3Le9ah7q+Q/2JvP152b6Nssk6LN144YgIqOh0jJgRHROChbKkHhs7fIehSgG29/t
KbnaUFvE9ZbW18xRlxPz8OhgdwBCq8rIgW5bGQ76yKw9xBwFAn6nIRua9Wq39pJ5xRQY+eq6feYL
FW2ABiDMKvlAcZOZWUOJkf1hnhRCuoKqFC2fg7mKP5S13WLgZKiAoDsNcM+tlS1bDoi4NUGua9Fg
jRhpNEi6XJgxo5NRtIeCMZe3EzvCaiXP25JnK7R7ZzYZnoJgniao+KsSHpwLg1+LgDohYwsbr/8y
6KXej1UJuS+pzef/zIMrVm8RuLQ3DIYPUB6QI/rdrDmGzMGG1rmtryGzGb96+WsldhQG9slEv7vQ
W8olArFikTgWmZcOHg0JnvSVo+iJw/Sgdf//K+9WjO3JkBo3XOzy/lj175SgBwioVGaqpZNTh5Le
RqtvLVq1pMuBz0sCtX7PfV21fyu0N1XYFdgd1grtKotlsHxaYKrvvsxSUQ2WRgQgM/dHdhMCm3p2
FjnHbgDsLvNef5ANqIVR7EZT1okBxxQTgoQq4FRUEec0z4Cb4sxx2ikOWZ1KdzDEGxjRZxn/wHxc
NX8kcs2VrXm+f6z9u5GLS0IKs4Pm3rFJUY0o76Pwg8+Hj1YVXxITH/VVwdKWIyX3UBMG3uTKOra2
YBlmm48SXg9SE4ozrW7IampYlfYeQzDhI6UutV0Eh3g45IYNx3qDgV5PMwizvEMlHXPfMIgBLOY7
R3qKsXWmFxqezFL2gMJb8UYNnHyevhSN2gZlYMZy1LAxpKN4YI901QBKc4cEELNX283ZWHkZ1xpg
q+w5/zySC/j7YiqHlX/Zkyui8CrX2fPQeZBA5ZgMHzdtseyFilgaC4yHjlftxzuulKU5E83tr0ii
g7tO52qqt6xwxXxk3CSjkgK86uS6nPg1hk2LjUnFL5D9RNxIkTezRZLVijwHh2u2V0/fapuGpX8r
E4awvMo+cOwRC2ssPpmi6B+ktQfNtimEyfbd15t/2MCkbak7/uJFWTYUS9qjdtnLOxXfBvL+wLD2
z3Zi+QeLCeN187Hy0tJsI3vimlqf9FeJj0KCqOcYYKUOzjueDQp5FMWA8tyTuRDqGPcQt8GF1sYm
5gXK0qZMqAVPNyZtdku8BiLLjsro5uEoRayqcMGHjZurcKOkafyoKeRaCs1UAZOs4coTFiQWUm/G
T6JFeihd9H+T/KVHhn0/hPMbRmQ/sLOoQy5ROKwfMlZaHCKq5Rn8TSt9YjmQ/sLHoPryCLsO1+Cv
uvkGKQ3Fp0yjdmbjN4BzD+SxFQyqMfhJiY0CRoFz4ztcTHSKVIvRUhMXxMqtr4ZTwPYzT3rWCAmD
HM6xq+aSyRT5ntq+4vuIQEpc+ZBKoDRDOEkKytBvAndNbrP8uV4vZZsMed/Kn9e6eGBLxL5YA9FC
5zA99bF2ljn1S2KM/Wwfy+gUJE7k+aQrpMblBjM8M8iXvia8iIV/Ywc/Kzx+qBwX6zbCZ/NbfLfL
3j3n/EvqYEME3vdedfnnceBSpT4nsCDZJGpxxsn4AartRT48sRY8kiEegKhctbBft8kxS43K+QWz
vkBB8XkaLhDV6A57MCTT7HeDh0hDas9PF76VYb9Ecw94/NBIt7LaXzAwDIw8zwk3b9zxbygsyPD2
70cUNRqBkuuedaETt1cJG58DP4MraW58MQdHXADg8EkyHcjjn5GoTactTIj+mXGs0sE/YGrbG4Yf
c2NNe0foZI3H4zNy3oYaOEvTJtpFdvrXWepiaGBAt2xxEFmz2mquxsn8fPYRU6K/98//ziNkhHvE
atPbZJQbRACAlEpFxWjjO1G8Yn+VyUjOzs/Ojcvp4LA5UU0S9e+DUp8q5JDfcY3xw0Yj/jHc5tCu
AaiY0LIcoKHtYEbw6vVPqOb1KfGkwtDGDU00PzvPB5byedD+kG9Le7UAPrqg7QHC8+riwKYBoQPE
1TAYn24rxfJm3ATwxX+CIQ1lPU7og6617fl3JvLT9+FYO/4fCqp3UeKXy2a3GPHawpMhxN1/SPsT
SMJhxxlM6VTv5Q0HbMdq29OQtncpyl5lHtkwEyl0bbNPpLB4hMQq4vgj7bZNEGpMsZftkm9oLaPj
9CIMPm7lmvKxHNmKtjYK3hF5pZrbEoR2agp/8CBVRQ+oWJuCwgmwa0XsBWmvXph6xUxW1H350zod
S8FKWaUrdOSkjwiLjnq30yfwbZ2G1HpbbhSIIg47FPIoKzIbaF66hPao7p/qc/Dq9QkC+NVaH1H5
f1hExzmlBj+00AAzIgspaKRCKxTyc9siCP6QTOvQIRasuNW7t33hrt4Cfuv6NIqQieF/KZbOsjzb
153wBdEWCVvzXyivCAgfKmnedRpBCHIIPKY/M9C3NF5WgZ6RTZatqOK220lakjAaVw29iRAmy0WA
5bLAbTI8gMo/70FeJQwz873sgho5C/T+tyEoJBDLWoPbnIDXRznMNaoDH8PhvH+RkQfC85JIC16H
AMxL20p/DZx2p7XYX5QKGQx2L3GDLngIwMSD81woKdFYoWji5bGTWEicayMQvKWT6Ut8XVbzwdfG
GvtmKzfd4Gmf3KiaYPsqUK5PrGBMF9Y1CTBWdW6lS0EF87ZkaiGprhhuuBdz6DMy7OPHTgkmWkeu
mdz2+NJLnSL0jfZDzwoCi4xYpIYof+t53yc8cKupiCrZg2vlPqlDb5vXEckjhapkmvqQEv94Zlkf
ASuOYs2jPvzNlO1hPsAY6Hk6VSQqomRuqHpgiuRtIfjp5h6eYfdNQXHX1Hb3m6KWvzm6YlBO8/m4
vWa9Pn+/ExEjefHeTrLn09zbK1FWfC05QYrzRx7m0BxbXt+52yzEdvN445eCLWAQEtLalSzy+BF9
f+EPG1/5eqYYSOnm9v3UzWUnWlrQ1KyW1u9mk80hJSRQ5uui54/xYSDT/SgxNH9QXRAudBPL7F/h
g6phY4T+mf9YUKuXjn6WHBH4QrZzJqADI8uPKn/1ox8cGDiCmRolRRl+BWmZ8wgB505izJBLLLRK
lgjsjz0Yilw0qMcp4CNUkHQcktcnoF4iDQ0jNsqoo9AB3iFKfy7umNROdMKdl6+L3ci1tPsTfdxP
vNhkHLVEHSd4xDgdKXu3Fao8iBDdLegxzjNeozPvqVQrSNRXLTOtr0EndcRBdo28gMZ6dqKqF2Fy
/ZidT5pR5TZBcp+thzBo+II3spLufpV60WjNVag0RZOrBL5oNQa5WQFz2ZSqqzwK8jR0r44hadau
BgWsesmljqJEVbkBAYv4p9B1lzlWfVE+2KrGZlSr7gHJwTXfnmjchrCUcUeMKIhIkZCrj5E9oxqN
Hv/n4p6uylgCj4tAluxF1PMfPyI/NEVyOlOotzJb2hBZ+y6YquZvXio4F7UFB1vNPQq82dZzcQ7q
fwx1x5wB/m+O320Mzksk6hKM+X99j2rjsUebSHYxFSwYAS5J5kSVREfS9KtWFKel0Wp90bPJMK0U
6sDMMt/+fQ8pCQnr7kjBqEzLDZyXqYhQogCxtWgFEQjxuH3rKeNTFl8UQpeQKDtFHO5ey7teDPHL
UoTQeumaK7vBtu8D1QraQLCcWfawWW3Y885LGpDGMU6Qx0RWLMY0wh6PVs0vz70sGAVjb7fv3mbV
YvBRB3pqQxaPlv+wPqJs7ls4rGHVdWWVnIAQ760hIB0KAk0H/TK2X2QeErqJO6+uaKj3ouX76jKj
o/cq1jo8G6ej8La84v/Cp6Kwag6Nf+yzRLOxu8338GH7Jdf9GqJ4XdymVOU3rsutVjhXtx1WTPqS
E0acypGBoHBl61pG7Nl/OZ33uDdEXODSOx6DxcUkeqKHHjht8aR3QNJgoN6rCqM16C8YOATqz0Hy
fP2Jy04NuHCJx5IpuEQAYeMtc/BKj63gb7gYEuC7QB5JOoo/r69XAZnZjsYmN/jG87d9wH9uMLNW
oZXHSMdBpFSfA6G+JTtvQo46PtxV6GIokfD3iyQ8M6zt466abyk1/CLcNZ5PbJQpREiKWwPY2BSq
9ce0hRQnHxdNIX/+DbGV1P0rhCQUSIyurWQa8o0vLOk2Y7BIElqkfb5t5lEKfq3nWPIQqBsLGYv3
7GqIxexqzO/VXegeZxX2/fK6EGSSI5VOdynIPXCl60gR97y0Zbb+RGy2G/bv+xHmILFNuiQEwsj9
un+YXu8R8rbR4QOMhMOhpWxxm30PR3wJoE2raBmr8JxXoVZ2KV9hZx4qYiNqFaNt1TFl0P61/nnV
0lLl8vHMWt9xUP5mWyA5oLQ9DyNkH3k7Iu+3RNz45w65a4YBi0Yz3pxhrZLaLtrek5hlZSWo59xK
t0KteWbhHwhqe85wHM+gAJ9vdL45a9jDwqogLRdDKExEysYxmOaBKobRrXK4D5MKW70/4GN6U2xo
4OSfehBGQgeeeBKNwXZiWkuBs7yDjW5ffZouit4l2jtSZ46uIxqJQuyiAbw+qNQYRyI3daY1mFUA
gllHBNJaq9PuFWgck6wldbAdHW+xagf/7yninLyIceD/6C5Fy4YsA1Ba8zCoBgJLeRKlJ9nfaBqI
y13eqeR+FYJa4cIzVw8g4Q9BD9o3X7i8RHamoyZi4d+ksAAyMOUT7O5FitjFRvX4JdvbPdvX2EoX
dsrC/gSpjo7iAD+kR7kanjR9EXuGo0z84jTP3xKKUitMG/qkmihRMrjEvqmY1Nt46U6AQEai9f1y
7Yknu+fyP8aSwtviHuxMm9jrOBWT2+vsTEmfWQRbN026LaFs0aW492F7KQD4Tk+Ga7RKqh8U70uq
HPypxKMRG6S1Nxn+CK4lMhDvlNtNFD6psyBrDlMRQxmXlnzXPmehUyqZ6QlaBVe0lX0ONpLZcqDG
yGqJmFZ8dUnKiAYJrDqzQQoDD29SU5050AXs6x+lU4kpQYu6HSR4ZVzIHRYA2ah2s0R4VZFZjQ2/
I6HoeRifxla7cXSwUdnrd4oX12nYSawM1VKk31nvfEZt9dloe285A29cCpe4dKit9JfCPVj4Lzdr
EjsiDl9REOxxQ/SsDa/3PFmJ1DCb8E/ybqDKY6x3MBZV8xdk1gvxpubeWspwLFsMStHVl7ATA4VN
28XvtPzx5edp2+Rcg7ASOsqYV1n1hJGnOPAV6iRK9pg4NVhQRmK/C/iROvpBDRyeLttfzrH15ZNx
ZF7RFmE8Es83WpENO5t3vZWMaybF1n4U2sJ2UUiSyTBkvC8wQO4Q5VPxtz0EDMEFoUb2S4gsQ93c
dqxJ9GkFTe35C4+xTTFLByzMgtFjQRl/9AjwtWmtlwm8wmP85XgMg4nQFaIu1+CNtRXAbhtYaRIW
2Wq1eppiZyQ+EvoMWvot68LIH6D0SkIhD0DNoFER1/rLuZJro6dzlYbsCxzT3CFShtgvYbRlwpsh
DbUPTwNcF4wjPz3vvXzwm/FamCmyVvobcOPCL+e1ad2kULc2c7qRj0LbN1gGCtlM2ERZFwlroehz
L12JYif0rpcGtlkKCMum8HyGHA9DpHkRQYSIzDMZ3roO24fepU9fBV3pj5M4FC7g/LWqoRd70ij3
cPjQtIYm+Z9hu+0lVY0ETw3lTaEN91WHagWByTOpAuyexVsCG/+WlFFZrumZqWQTOr/amv+IB0oW
mW+pvGodTU0SHqQvahpTBMItGvl+cV4BApWwbiaD59l2rrKOY+69gC6eTVxV766ZKJ2CqU6Uipei
K0axZDKVs0JKdy1nVYGOyrGtRtzTyzN5HTXnv3Am4KHrbX/JqIPG8wituGFfBtXZMw7hCI+mgS52
B+5pZXh7QrfJDPyPbvrhBbzBA/GKfZuwkSfaNd8qwZZipe6NZ8P2OcNwJd2kFaL3+5raFr19evhG
xq64bocNK/Sn1CMGYAor7eXDZKqtS9/+RCCjviq7m1iT4xUI68eJ9c4Td/iKG01qbCyi8vPFLI5L
Vj7+ejzJoEi5g5uIBX8kS5fjFRtBfIzo3IgdMnNtMQvo1SjEE1fLsIoMKGNLph32uqHwIKONUv/4
6sYp5fTIifOrg5mlkeH7/qI/VLCR6de44iamtVBdHL/2VaW38/Ps53n7oBpxw9VtOWH2D2Co7i9M
6e279U//+nIhmtBMhqN7SXNQdcdFOGB9q5OKXBtONSbxYd9nTJhuAop6Qr2cG9E5P3kcI7E24HeC
BdeDPTHCj9v5A5S6czoCCFrTbIlVZbhi+0Nw/FzmyYt0VL0sNMC6bEq28vfEsbF2On0TMjVX855t
0dWL4Wab/gIoRUuHMTfnAO3dAhKVAHJCV5r4gPLe3GvHLT3eQgbyBNQFh7N4//cmZ2g2n/aQuQUS
NSL6f7Ifd2M9tvm4fn5Y9JkDcYy97LJEz4nghNYem6/PN103mzEK7TrLDqQCFX5yrZ1BTXX+qydm
/GWZdasHSBz6hOR+WUx9vgu4+zZzW4aSPXZjC/FU9It8pr2mHCNY+01ER3edM35xc06zS+/qovzB
0hyvWZoAVT+B/AaF+SVfDD3skI/o320OT7XvcQmENOOw7Znyq2zsMge8ikAFUXeFJQK0mZXXMgRT
8KSMcGMy3Y+ZmyWmJlfxw91qFeVDip2cmrQ9faxpJMCHQunKiQ2UOMtGS0bVWrYid4rKnZmltACG
mdD+CjPJcElNspr418Sex6TeDgGYVgxavrP2bRinNJWQ3sqV20WKjfEGDrXD1twu2Iiv4LRtm5js
7AuAffnmdYbESrDKnNR4y/zj9kdBWhPXg91k5uj4Y20BKIm8yxNfT2/QPYLnP0y7ji7r+uy0Vkyc
wm1fe5ISOYknzBRFzU7XP6ql85NqF9/JutAUxv30S/H/R/ng7fmIdcDT8z2O0a/goWoHcYjWQfyk
vt/rwhRtLX7IixO1t6Acrthelta7HfPV6qmI84NMllzC10FhIvcewc9lga7rGnXVwm9Y0DUXtQO6
cXGASfL/I0FgGO9uQrO4KLcf1iH18yFiCOr3L9722X2sdPj04r8n1MerytoxQU9zH1hEZzBcHqNV
Ul4i6G1psekH12KgJMYpjbAuzppf4TtBDGoCEoYNwqdLUFgUXaLCvLIta8EpZEB6jF+4zb0yj7XH
lYa0XVFj2+XU8a37NdG3cw1inA26YbT1SKzi3IhLfKMn2QcU7x3BcRxRGRp9HVpZTOOKm1RuxEWX
pDKpaZt+YIBB5E8nzrylCTRXRLWiXjuoxUYI+PH/FtLjKa2vfBAbkLpUxA1d70ktMH5FsXkfC5TV
VauFEZ5YB+MPVAncfWvPI/b1cOF9aq3+pcnQXW4hjLjMdaBC2NL/Gd24B8G7BJYHMxZAUS0PeDyu
i2ZGEGngCVFui8k+19q6pARcyGvU4Jlpg2tY0hb/Aqjyx1B/+fkbqIuJUryjyNE6j1Oe4F0zOIA3
u5ILMcXIPmRiZDo7jksi4A9ojDdU4+06+gkqjo0DGmrcyTh4oFvRaCzswmDBmol1BvWvTgizaxBa
Q9X0cE5+x7Xy7V3KAy6RTLSw2wnsYTUcbGmwVEUViDAWPNBAk8HDfmMRc6tRrnUlMPT5ZI9gwVBF
RAa/HE2CP49HEWlPySCDSH2WtxRZit7No1Jo77p7/73oGUcPo5ubtdNc1IdhiD5h9gIL/wXgKH39
L5yisboJT1evESYEmCKSAbPeAvaeNigl2etIb1CzTq2br+u41mT7x/Rf+P/rGZe8ZpzMVCsM1T+8
EBWSBCdz5i2eCVSHELz7M0AdfdHxgtdZpdZ9oaxLz+qGUTuU3poANEwXmGRIirz+qh2e8WD4W/tf
HYjTCnchlrrCq12HVypq9WVRyZ+8E6+kwEX/F/CC+VCAQwvrhb3LXqWtWNlS4e1i7VHrSV67GcU1
MTLlvcoN71ITF3jfZBj+/uaXAABrhWPyTSCNN5m6fasCkw5uEQytM0mgFKc1rxxG9zlxPevLBrGl
1hs8HGgTR1KbGVUr/V9g7qh/TcVdq8SFUN0vctzfiHM87UNCz+Idjr+HcJl08HEt8Jrt5PkyZv4L
Glik28DOqs0Sum1kYDvQWGoh+WV0ZlxGG2GhWv2IGYn0XhKJEFhJVM754Xwn3mmT9MiJkaAdDrnh
SwCpGJtLOn7gHroUyRMYFvPBYdbMxUXK/r1ehbChakwN3/TepE6eVdmXL2ol5mcLhDc8oamXFc7I
+7HhUWGiklNuc9rUaoJEY3FxEYO6B5nDjgrYxZpw8VDwLg4fkwiXCF3dgbwg/uNkAuOdqjoUJrax
p9nM+w1lH6p8gbCvhKJKCAQJ3MvUlyluZexX/r8qV1Cxl/O1or9JojbBAl6GblBYKuV/dXFFTnee
sDL2E7OSfkj0h9zhf0CVPjA4257MImxCwpFitnWdSXD6557rno9019Q2iW92DnOI7IZ75uqUJtGA
ZQnuCBTnT48u0YvCT8kfivdxHTWrHqyfgQIeNbqp8k+nKSdHiILubQTZh2kXdB7WQYVg850gP3dx
m5jyErrNq1lBn6Xp2Smjpgkpcav5BE1Dg2oJ/OIRKpj7hfJqdPNb40aBAxEJMVWrfxYa6GeL/4iE
MvdGLyfkw0b8LATQM9Tvh8CsALg39r3mFFyYGSxJakfkDqnY0OYj9H+huhj2Btg2WtUqvnfdMGMe
mKv58Wml7BUnWOMIbit6UteYhGYbFivMvq5CK6Od/07dU9GHLHJpVpknY2mmX633cuq9TZJV7GnF
pS4iQCBlthCx7tBSWhDgWxQf8CTjipLoXQxbM8UsvuQ+g6HrXlVS9SkuzC9Bgz+pouT9/O8K/YVx
KaY4BFiiO3B2EzoFDME4abWQFGyua9w7u86zhdKHW+yQ6CWPDNFPq0k6KooXL462nTpQpN5wrmMg
vukZOFQSzwEcQghbOVQ70jQsvKEwWsCsnp7uLqQOjyrWj8iz9vrP12IcuktAI+SN7eufKFVoS4rI
tmTMsTjDt8sYfgk+mfqczfyN4ceCjnAWvd5MqXR1K41s4MSl5VXdsBHmVpoKQ87F449ZiCb89M0g
xJVcfBWbir+I/wL9Dbnejwxd5t33uR7ASYYvts7wfPqtfT2Faet8Gpx/0cj/5zhlM1ykVB8QSoDU
U5CtEJYP7qEfkTM/GYUpjTGvu/hF47Hrsl7JwXnn9SAVH77D7539uTlx9cXXPe8oOkdeFpBUqM8B
biIdim9IjgTyo7pVRU0+TGe/P9nfGTWiu3d+4PrbQQltg8xL/poBreLFRL/7NhxlT74kOue/MVf4
nnNzB1McyX9CNMnKdKJGam6l9PNLaQqir9muCunNbvI/yQekcM5yt9lf5TQKfhawoqZid4OxptrD
S/YSd5pdS3Jp8IMcat1TQuL2hF0LDLG3RI4wpsZ65KOFwtWAthtikTvwVbcosNm+YflCZGW/e2sO
FBm9iNrp9sulPIKp/vuKnNWn2HFh/MTdkMR0yOumfM4ePy2BCI3TXSi7FID3Aext3Y5n3nGErAvX
2g7wdnoSy/oAsfn67AzcfhmgTwYfRp+F2UNZS3jCVo4lw5LpFekfwi0iVSzfcnmd33PUa1bJHu32
3E+364wWiCtGaYoQl8EmE9++nzBJbcr4YLn5PQd+hmaTBixRz8Y6qSSNXeaFIXQEGFFwr4PaDtfn
uqw2Mq8kgIEvMJIjNd1QBNX1YAgB5CtU3WkqYrneyOG4gIG8kZ0BG2HDmQQif2LjMuotv5cPpYJt
LJUolw8D9FOfk8ev5lDzp9UqEHmeO8ze5W/3x6C+AWW+r8j4A/Mj0ukzfqIq8dVVYJJlrwl9u6Kj
p3a/Ue0T/Hl6sWrHsaxa1KiD7WD2Agp+A7Sbx7zpWaqLuCQGGsRQlhr6Q7y2W0IxaibPRRKeAXX3
9f8VDAXlNCcW6RNU5h9wcri754O/DkqOjtsDQnqX7AVgxUWPSqyfk936yKYwlvVfaKlLbuBt65+K
p/0EbkBGeT4EffSriH+E/ZhQ8NchKnhrifsOud1Sce9leQa/rusuNBZ7McovLgdoMDQVtZRL5mIO
tvthxLqN70yLK9GMYHj9dwvdZ6y6iWTKy8g+AiyN4z54kkCVgWlPZl1JsyP+rnYqq2HKPPVXk4x/
XH38u1YsVAkSEg6i9Kqd0cl2v1S3hgMnohox0NEB1PJeHc3tdtU9JylR5MAerGRFc/FytbTzjwG5
oE97WmqN1CQ8VoHFht1lpSxvdR6oLMPYWKm6vazP6fRgAFVSUBkLyntkrDrESoPsGHE9rdJvsSqR
0EoBI+IaD7bYUs2wl0JHmtXVfaqMUeGDCdCGDK4ctV/7W3OQOebRG83/adqf3smBuAMQsW1CU9KM
HCb4nplMDcO3QEA0jXlIaWA6NUb7U2cewxEge2G7gx9pFI76jxODZugoNz8cGqerny3A6SLCA6qn
lkK3MI0bjboMvbAJ6iexVPwzPJJFP/O7Pb2GT5KrV87UkKFd4cFrdF7ScvZM63W2JAnBwVNKRH0K
v1DSAK1Ir30yw1roJPm01teNyCLBQrGGa3Ul9bESsI8PE1hQ4L5PlJI0RWCvvMgwi9COiENs6/wD
qmPxvg/EJCB05z4P8e684VZKnHh6INjAHZwkEHFtQkKTbqqW/G6Gc0TfkTRFJbSdJ0hzXiB+Rcnq
OzlX1ezK1NSkcw+qNUQ0U4/iQVoabhGDqLRqHZaNI0Y4BaglPDf9x0qd4FvSNnnfvqAe6i7OFFR4
lxJ0vtwQ/Fnys8ZtjJEEUPrziSc6tBzdi+jX9moyOZFicNqFTpn1XkXys8og8NuVvJuKKkmyuaxa
6kC03ckqQaLIWOZnj9rZ559EqgaUPuc1zvmegkxAUoces/J2avJ5igcNnkMImXGIe86xYEUj1fwc
csJ/K+Hlp3r6DHep2A7vfTee1xcKOhg/LdXXDYJ2Y9+FlK8wxDhcJXfyEV1RuM8A7DAePWOEU67Q
0eho+DB1FcTaxNPuUseOX0oov2lVU6OhviXt4rMH//2n40Qo3nh7/fsTP8ygxSuHkYvCoU/Ea76C
jd+oWNNinOQzn1xqKbJpZj/LXNSrmp9EkbC2ei/0EvMWfNMuWRZWlkK2CzGmCaj9WYHbT/9HTuPd
gOFr3s6XnUk34XZ58GHgSjvnbJFfcTqRq5Rs9ZLCGArapAwkEvoWSSlpkwF94WZzwXNnrNa5UBYS
wEL2p4k7jAmmZbPsaFEI4HOCUHqXSYs8QRRtSm3+WJOWQnlHoNb8cURTdiD/9rK55eTQ1zZdyPgQ
zbXAzMgdPtjH4iUaThXnXAtNQwJgFad50q5tqllJhhDapzAuKdxBF3gRaN8jFGJhnaXjzOmiFybi
pWtEcdN+qYu6tJ+VFwDNxDREDspWxlRTWyJuydNsLbn+2BdYbqHz/DxJ11HqYDWIYFeN6SeFEjeF
4x+f6kOk4q/V8BSXZXbBS5+s/XFC7V7A9IsKwY9gdU7TiyiwGhXkB1ukHWdAKuR2N7Iv1tNUqxsU
ZMs0E1nNjgijUIJ0kdhUQXexKio0fiautlr7isHDFi6zKoG1FWlXHAHsh2egkeNzupJnBIa38aJ+
QloiszancjvFwyYZOJfaAM88F2D0BN7LKkEV6OOSia1qJ4imiauOjn85zZypW7fZzavqAkwZ0K1S
TZ6gOScWNk0goyIrHzmh3smx0neJv/2SQ3B9lk/J+YMfSm2OmvswhdT1+0fpHzdD4MVRWTh4SwQb
nFAH5Y7jrdCyDPtjXhqZR7qSSKE3O3gPEowfjAvDnm3aGu6HHVl+uyIcDRpVVulZAyLtLHtY6Bed
cgU3GkdDCgWGder4dOXwUhMDUfFAZ5HFcLsF3H4FKYd74vg4lHfzOZ3J6tU6CnHT/I4Mkoxi46kb
6gKbuJ9aI/FHKOSu3oUU3a4TgAef8w3y2WlQYuRug86y2l4IBrUde/8HJ8Ut/zKsnviyFSXhF3Ij
LTg/fZofAnjBxBFBg6yjOhtIL7KFOiUxBQe0aDrit2GvIZ5OQG8+mHiV84nMqQyvwh/hfJzKBmxg
k5Futbqu3j6BkX82R0TCmtOY/cgKHm+bbZqLm5OqIPXsXpAjphal2E8ZDm3ItPTOS8CeuPdhQjYh
I241b6dPDwxyyM3rjtJIvtuSXYT1wRqR2vAB9/VvPnFE7cC+Yp7brJfJdGk7/JNvjVy5JaXnDGpA
/Gls00dHJ/d2QHCcMi/lPFfAll9WauwuNgt/KCDf6zYfov/ezUqBXwfTY8e5S0kBN3rkzukX2Npd
NgIGiUVGONddBWGYOtlSfoOewd8P4Sla463Kx9SVgTOgsWF+m+a81yL3UvGzYkOnflSvXiF0vgb1
QVqzRQVAwv1vh8YBEdwAvoqP3COGbjr8MOBUKKx302RmAYx+ykUPq5x/PrnLt6t0HcIgtmy8xr0P
OEQzk6vZ+otnmvmUHy4BLZlgDCFaoc4EMfGHH/+5F9TWh8HAV8GsMB97HOxZZFGeSHGu3XK4JD6s
igbEqpbp6FVNx6teDoy50ltUz0+QlUXr7LUg2Yrzf6zPHY8XK9tT4U0nqMOri6za9R048NGehJwN
wo31wKfLZnVII9st31uo/L/+363t76KRfg4hIgRliJsxMyE15uvRhisNzAP+JECYArc9IYnzNb4o
e2SlpCk1phD8Vs9W6u+7x67Sgyx15s/vdZHwpTSj84n9TSQeV729gGX6Om2GlDVgQDZ8tR2wphZ9
vpbVVL6NO8zaK6Sm5kb5rFz6l5z06mkfBihhxhtbymo36NoXLAJPqkUJfxSXDeuY8b0Ss4N78+NO
0urmXgCODHBv8dLVSVmI9OCQKUTyX9fncgXYfiZr0zgHjoCe+01ezPcLp7szYJYuWVp6Yh3QI1bE
D2jIMkNEUzlPsskUPCNOCR42HVVcH3PAon4CKvRxxdWvlnhaKO9CqwEv/jGiCq5nG73/rKPD7jRz
7XwFrOC7ftf00gnZShzB7we5mUY3PJJ5QXM5Xb58IoiM6KIths3J+0XsDpx+7FEVhe1k/8zLHF7/
mWrMw6dfUmUsnzob1HVfqK0cZHHBFDqCWeNNF9WOdGuPal5qU9TEIWZCGjJm7WnnuC6WJJVx3yYQ
fjdqpyDIK4LWob96Xb2Q7Ecb03jC+yldA3JCdTaxOVD75TrKzKMRIr1td9A+MsWkh1vp7K4WhX8N
R5Gfb049I+qAO/WxWYKzpNmhTjG3V10WXd9/ZkhOQHuxmpRhM2qj6y3SLcnc9yHfs8mVnJ9filv/
P/ZCTUybKhAsre1PO/TeKQH8tA6Utl7qRQD77jzmEs2POq+je2EhvBDJ5RZnUWB6iYv5AhT3aZ15
9S3UBhuFMqU3PuXtPQjcN9mJ0FYVP8o87r5Ehc/mU8o++2AAS6CenqN3gjKbDQATfnxiuaJizXqm
yE4M957fPKrrIiZMsNI8wzqdIOGdedBlCGPM9oeieJrDUnjPmFZnuvnW9AHtgBBmsD7+2Q84ftKW
XuVkgDw9heqa/pAW3Kk4xzUVu1VA3sRHvCUGyTDZdpKFgcE0jw8z4JaAgr5UEzgnUHP+0hnfNJav
bkDojLanpHnLN210aRkVynYmqigREKNaoZQvrRav8LUcEWHYdJ5iKi5iozqrF1paICe24vrh03rJ
FYSdKYXJXMtYXlXyx/C96RE+AURBRSBXnmY1IUItF6NRmVI9grY0DSUXzd1mxx9hLDB4xoRZrZde
KJc/QtuTR8QVeyqSFQIsISHwFopssZHrrFpMaDuIMocZLhc53omDwR832kL8INSC7F0Hqcj6p6b7
wMXHL8nJtunknT1iOt4/kqdELxxWY7NjDEhE2ZRIENBoF7qLGnvWCxOMXPqLS04QozzKeV4/kwP2
8h6db+W/bgf2iigiVcMYFwI3oq2QeexK05u/ncO44VIZGw2iepFfwxgDxPAMvjHfLpCj7yFqMiob
+zsEffUwkqfb0CYNXDqkxdhwiqO7rf5ttZf4N3FbilshnyJzVb1Lvd2ZnxGMfGLAiWcsTvrOSdVm
ZfhUib6Ef7T6VIWRo4+fyeiUxirf8F4ro5pjlTt80tgtor7FjNfSyT9IJVZ/iiM0SBo7hcXanMEW
wLXSPmKhu02N4ZfpMlvKVn8caWaI4cKdnpS/Z8h0Wxg0yjFe0l4RKERMnZe+2CTRiw0+feSA5Kzu
t/pjsc1ulq+hxhdjQH1l/zLVZhJ5q8QPS7eYBbHuzf/cbmmLi71+kREGWRFUcBlfrIhu2b5Ewmtt
sc5X/NdShvgo7DQ6V7zlwHw41MwKh0BDoQgqpvgklV+Yyp9QNDMEDEiDebZmV+qCjpUC+K9Gho2J
swtDdqBgFo+yv8VA6MSxxQ9WhNnWvJ3bXKnnx0UzGhuOZKQZpHR1NHKF4Put6QJ9gPqM6hL1tqm7
zWoSm6dFt8/YKgNsQwdF2OBmjzeL9b8kEZxmA7zplivCGoeVKmgeuMhVC8fGMAQxIWOpFrWUn7F5
/mgr09V0GhTzRr5RUB0iD6NlKEDHjPJA75Hzv0+e0ifylw3QpOJ/glmS7JBYSSzUHld8naUlHO8z
LQ2oGY0IAPhrahV2P42VFcwG4izSWxh6yErIxNSkogLGJy64x7AN+pM3YGSe7emYBzh/ElpUfcI/
tA5aE0h8/O7j08WEtiqtTTfknCWWAilYA3psHjym+wUIMwfGCe3CEX852kW0eszKNZRYIE6yLCnm
rTX/KAoqvTV05vcyuV9Dpl1KivqodJUxh8zdXVtG5IW+hAQEpAdApoVCWf8mvaN1yhInhSNdDfLM
ewoPDHBIYMtlallCHcMxwuR56kyOEsImfIUM8uWescPtAsXrjGP/Bc44suw/mQS3g0+iIQsScEaz
ziM+/JHU68x8hVIWWxhTjE+lVpfkdtDbtpQpGYtv9zma7KcETORPbWbcduiZw22LakP/PTlVlWXL
DI3qbj0eQnkF7XSOMurnArrkDPLPl7jmcoHDAANfX7xnbL5vIem/rB7WzgxDKdSHXWJErAjF+s5n
uFg06LwQormo21rQDVJch/548YmmyOLK2mw4Y3aaxlv1giPziTW36sV3gyw4yq1aBcYFfUISXZ19
S5uYl1CzJB6w11RCzgH3lgz/b80VBtQbUKi1fDwMirLIuIhWojqc/b1f+FClLmKLjgf6/zzIrnxN
vGf4CSPQGK9YJcWH18GIkqhRtfeMLmmc6BdW6pS0B83VhWo9HtkkyGaIDZEnKXcvzktlvddw6/Lk
ZHtj/ZJLgNTzuA3MczT/6rVSvKysQhaEoEXVnvem0dIjCeimV9AlF5QuDIZiW3PLhUlWmi5mM8cb
IcUTdTT+OoC1W+IObnnC+zOjOwn1PTJfzEBRqXXkF2tXZ+w4+dtThDwMtjwwTcKMzW4298ey2PUq
IbQE5vjRR8VrKRjM8VMhNgOc8b1lSxFqVt6loDrfVyAgLpUFKj80fOgrrWl99dSi2WfCGQf3M16C
hsw28LN6PNGarusoD2Lz1KmbDFTg7U4LQLOwlQBxRYr7d/OS+rAVRYZP28O1qF9ge1j/kaySI3mN
ec6+wlEwPilkVn8HYTRWKPcyOYvuqHxJys3ich7V0P7tttrC07ayZLDcjxF7H/VhHAlEniCVhPCF
QMb/K2Cqj0whQlPzNr46n7sXwEmXLdytLRJFDvrRtVwS9MWK/ZrY/Ss8X+tKG+L+xApTsGWoKW3x
2HDCu5nYXCZnwmZdwkKgaongMdw3uioHHZcvIioEk5h+VSl5rksJ6qvhlTmkgyrI+PBcGJYYCaOz
SNjrm3sqPqwUBpMXyrbX913kiRWAyOZO+LMEfgoUytCto+l4FNyZ3OyoVUVEMpN4ylODCGwV/r+A
5mNdGzEFDbs0siCV9GftSF8WNUMgLgjoGdslNOz9kVaFQ1k6U7iZzGlby0xyOydtrBuZ1YnCe33H
CbpoLCZSbjO/xiz50oOgVchoLl7xBj2dSloymcYs6gn0rmfAMVjLQYm4/Asx7o9K+7LNEfizyHRA
g5xXEjzLcstubrDIOxcdxD2INJMqjTbIW9WUIENi4L6kFuVp2C/AsFDdWTxUs9WJ4t4JJHj/OhdO
7eP44dgnnM5HOHQPxY1tO1BK6Ri27HVDpNONlhu1Lub8KAKNDhXRDBfRvWLwwshpICMB89om7obZ
jFlpRwdCvpXh6XVsZwYXA/vqy2+mt29XBtlapspiJjhdgc82fxhkQCdfTuo/rKwv4sJTUR8Qm0OF
sVJzTVb3tX+QJc0AtOH3Xf2gUjBKZYS8DR4xOI1Se6NH7VJbkEwrBKoO+ruTU36U5wtEX/zsh5ap
HEfYXuueQwMokM5dukYAjxhxuQS8vFXQPzmKSjF8uE4POxUAk3242JBsswXzfbBfX9pFlNnUvkkA
DaRDwbZQiahx6h36dHtrgHRS9MPZlYggvg4yu6MN+JBlJJVSFu7ZVWenIL5sU5WZJMz0Wgmk9vN3
I0gyCBPLGZzI2l3grXlvRJcGepjvZIcNe1PiEizplIjvYlcqBZRWC0swIT+gYj5S03oq9iQBsgw3
l89Ez3aRjx5Zp0ZZnDx2o9RFA9KA8EdOHM3fjkxO4Fskxt96PQi+IIdd+x/fFPy3XHgvAS9CAp4V
REe67HIfLLVb6rNasAX0u02ZpgsxrdqooTmcBPK7Zybo4F8/Rs2kRAsFBOaKhucKsZRXn5Sc2hNJ
DozLNbKwPNy4I53WHIm0cCtX7Ru2pyjJb+5rC+7UoNZOxgN5u0G122XAnixna/wem6oeA9wPZ4B4
dw+MqIKyjycAwF55FnMLzMkst0vtOPp8ZFN2EaSFraqFOUFVF3UlqrSgfHgoLdFl20Bo5QuMZBD7
ryLtANXMmKAUzbeA5A2sS0gMy6P3k1YcTyRvXQVVBwjeYCR9H9rDiq4xFhoqEaG+s/sNt0Uv5r0L
5p7nsB94AjMjwy4k0KHPPcOfU9z/BTyX0on+LFmNWGXbjkRcc263AjdyRVEpte/c6mQ9wBtCt9zG
YJdyWeMw4qvlUkGJd26UDNT2nVOdhYJprv7ajsCz3XFX5Ve5HjGAACuyjxQmhNfhlxcjnawUc1Dv
IsZthPxQ+nzyEXwSqggh4hwyQT1xEGjt4g/uaajy4tS/nk4QH8VoG++38MFxZOYk/puPA+yujkd0
z0J1KecekAFhcWIGljaO0LrwDwkPXVLztj4fjb41IcW3ZK9lq5YhMBe1p0OOYlbMdUDqNXiu7RGc
EbZBtUBM0Csefak7ekegQTRs2JHoy7F8G9loKXjQL+RvDjHyPm8uYtF5MLwGgVJ7TdnwqnrIZy9e
dsmyQ8qOukQsRez1JqCwNExzETrF6KMwPBnRmimynhn1N/qzvoMDK+og/3G3ZDf93m5epWjJAOHG
8N9zs55meq6HiR7MpwH7qdr2JDUwiy2FhD7oAcBBhs7dQbu96BQnbLhg0z87tBJVGuPjREiwdyha
gTVr21AtXjdfG1TmCdFfA2e1TPYE+qxKIpS+A9dgV4BRNvaNyG8ORzP9P3wpaK/PESuD9DPWNC98
GcSTS2zE9m/OOOpg9MO18a/tI/aVpKyCY8ivmVgW5CbnC4oDxaRezQKGD+5BNsePZIY4a02YY4dZ
MNvoC0dZS2ZBO2FoulBvM1juHVzjIYcRxOOllOlsfPy8QlW+NPDAyCIo0jD/TMybE4TywEqmwii3
wmbkkc6e1qlKgu9bAABfa5q63gFWU5hDdo/NEW16kqzk4Dl0e/1Ng9yevO4xUSrtRcTa0vYRFi6r
gHpTGUFF3v+QYgHQdNRyJy+Wz6YlGhJ/jeeijnTo5NNm8YxtpbSj2tqyilPsGy5pagV6l7BU+xdw
VSGBWq1v5vQnOTJAIr8z0ljNrg57d0WvFYMOGWlui84SFCSXIcD0pCrvthhqCjCN5bF96No1nA2v
gftk82xXR1TWaK8OVSTDFCtH3hXiKhEEH980hOwQcVR0UgPcNMSga+AUMUSvp7PHyN4YIMa1cBcH
c0aXemXg6CJqZsHw3O9xRA+pV8OG24EiLAKouI6cJH9CT8eWq+9nySaUYSBUBK+u8Codtlq1DI/z
tG22BJPOhxeLwYRlj+ItnJh9JKQ5erW0jdF08veY77qcFjfUQNFbAymb6inrgb2g5To3MNFcUly+
DXLMo4GhUQh8QZVzeg4FBM3wmVQGNlC+QfWP9rCv2BuTPGcTDehP+LNUmr6i/t1c0GpLJk0eoD0J
O7FByka17VXbxoFayvpsrYQNXpW+i9N7eW/45ngH8wBdOtVtg4oAUjTiKsglVHvAaM2AEDTeXGRG
hwZ3EzDDj1f0qAXqs2hfxNh13nAvPXF0jR3szrx+BcRy8cFpAw+bqjokDIO/aStgBXBQKqwOojK0
rpBws2BJtr0dRL0U7go+CklvzNA5d0pOSd3G3GOEiavZD4Q5MHEfG9nFsGKXdOfaWGJMbiRU8oPJ
4VX2Up5i0zCdCANhUOoPRS0GQZy2fpx4TaP6e1VTXwrrw8KNspJulPBVd8SHk++rEKOgoLTj5MJn
YjfzMwhE8gyaKNokIuyxmweR7qBUB6WlLrjxsdDreI2Ell8GQaNWnzAYl0bS8FpSv2MIDp5mHyBL
0ODOBTQIkswyjeGsfAp7QkTJFo80ommWKfyU/CTj8QK5l2OEi1i0UreVBLI2IY9uKab4cKRnMGcD
Jwww4eZq8fPr/t4N8OJ35sD4OhzJZwz7VNeXby6kjY79I3EvqYiE1iZTMvl0pTmVOSSMdq2Wm6dY
nKjv1bwTa4FCD5Tb2DZVfRhVacXfqlVsfirJ92Q5uUNIw+zCTD50aEG44AQClgwMPae5XOeK5b/l
9PtJvaanO/7ooXdWNmPypQsGmgxnYKWMM9CpHLnqympEfYIXBarEesr/ZLwHur2MeaK3gOeVErUJ
hc3pLHCyF/0rF17ZDqa35SA0kDFEpaJ+bZFLaACRCvMsnKIj2P8JCXodblrLL9Hx11KOqHi2WrQT
ogibu+m3oPmWb6oBSoFtx2vHYruJm7e3Uh/9jlc2I+0u3CngGIp1CdiZOcpiFk5OV9he73bsDblC
+EAwAZ0f/Cp6DO8ejqE/Pwtwvx34IiUoRF5kcunr5pVIeus2DhNn1fV1VjD2beDM5rl4xZulI+uJ
/XaUSGNUQE1oAGulWtidzzZ+L9UFIgg/u/XbJdicZ0zmFw2leKzlP83fV31HwboLRQr0UtI3g6lk
tMI8B/ZJJoI6Easr+F/pdQZz4uxwNZKWUPQyewncwzqxYJZWujK/Jm4Ze/3oTCGuvh8HRX48KbbX
gXkPG55Dku+4pv2IjFnHz9t914zva58Ikyr6OTfPXKdmHGuxmT9QYNK60ikmSF2Q11DiCmXDoxML
Wc/rvo0vbbRM9s4ZcDYI2MK4lXHB10xk+0EsOJE3WTXIASXJ00YvSw0jPZS5ihAkiGLu/R2flMcA
DtZ9pUE9y4UR7873eqU6VpasuqBpRh9BvxdxRCCP/JBKXaYje8LSRL3bbxu7Q+KmQDuk62Ah2mQE
32QpX7NTRer5WffDqnHNLqJL2lvk7txy5vho8pK6CdjAjhPhnJF+2gAM4lVI1z7Sf5sIFL7jefQm
2ljSIYTkuB4yT9HyMEmtL4rQGVnYvqtgeUzD74S08QCEYn4QUElTugzdaa8PsbJUk2TCIpFE9k3Q
dShDalYSkaPtaZenXxn8kDOaeoTGrTBU00YZO2+fJM/7G6KAhdOaIn7yrMS2U+Eu5O4I5jZuURPW
4p1es9tjIGCyylPurAJ103mjtqXB3LJ7uj1CLAudTXp988ZJQhHrKCKOqgFzhLw4JatJnHpW1rdm
JBDFAm4p/z/DHq0K2P6ff/Pu/DHxDWypUDLjpkpLKdcvsid8f/FuKQDrNurbn2Z07mdVIPEhjFjH
7xymipytrZ/eZgE9CU5Q7zObcv7bW4vVRmmLIAfa91IbKSGqojkXNzhxgoEWPYFVYN5Sk+shdpjo
kyJMx1V79FyskXGIUxJVH0oyovql5lfmqC4nchSMrR8YvA5pKh0aYTyBNa6LugJOZ4sSMSWOmbBv
tuRpDU2KTu0daFnFuvqf32X5+qUJVgNJgkdiExT9hM7UtAzM48CtjbuuxYbo47XZWjBPW6vZQeBP
fSyN2d0Xa7DXjLiGCw4jCz1hknGBBkxeT28SFR6z+lmb4YYRhUW+vmTsjM68PqLjD86HdHiV4j6V
SlT3lRXeW8Ciy1GSKWPTgC02mQSxPvlUbs7py/IpX4AYi9Yk0actuveIO135LZ+2Vd0ksU4kq3S+
Dx0giIHsvvDEieSLHqYBwAusLCwUuLuocqHzDW7zsj05RaT3uRy7OrypepdKECLwnu35E6f8zCPg
ljnZOwwotEo7TqyXnJ3VzipOEerIIu5Ig8k+eplImQdUuwHC7bmXRJarlBdn7e1Rxj1p4SNWg38o
FraTpcuu1vOLQyXhas3aROMpdq5pMdXNelzYbK0YTKLDVq3qhobSIFBkYO3b/is1o38Pae+DrqKu
4QuGsLahgEmJE0MHU61euYHrCYdVLHf32Dq/HWTHb9WuzfNyInNrkgfVpYC/M5jW9PRolzjMwn2r
DWJg5pGrFFN6fFAURjATqOKSHY6ZVTS6XliRDxxWv+kDxjma4Egh0qJP4Yr2cKYqVXjAkIjxkCcl
iSJnxIzpVoyui2XBA/GiSaK5Pjufi8jeT1Br35x7N81APzeNg9kxdXUOfMJAelJMpViKQq411F4h
Gl2ShGAAR9feCp9/g6hFiXmYu5cJDulJLxHzSaiy75TQwYX6d5H9a8/Np18A3Gs72llJyEhrdNBz
uZGqrfptZX3c6geXzOpfap9tbxEug5/5LOzNrHJ5XSflKpoPyT3VcUyoVjZ17a9nTvdnNmnxvNXa
v8NFdXOhdwUMNFDw046JnzOg9S7DxpsHuS2kP2xJrRX82fqYib+KEnu8DOIaW04YhyN6qHT63+qv
KJTAn/FPpg+UiAJTJ9Lm3tS6r6UMLjlJR7p1CVIlpLnGOIRBlA1S5Nl26FGfM4KfCSa3cn+BN3eF
LXNZruMYID7j9bO260XUt6G49axKqZ0Jgf3bWvdm4QIEKplmt3hlvs8sIBXjHa9Gdc3GAIMp7sR4
U1v4bsLYZ7eM2ifys3SCozbp7ge8GKw1MI5Q6aAPkrgAqcnBnmVQW+MUJqkCeWdpsbGquPlrwhu1
eAhqXTZoavdYnLeW1gXeLPNxPJCrYhx+KyFl+pM13N9ArgQxirKhS4BDRdWUHuH70SD8Qvq5MCNX
Rk+pg3w5ikW6qeSYtIH5TvBgZXKB2V9+Fn/zeQ2VkjoSob3+0yXZYcEls4oFGT/mI6FVasN+/LKR
g10TkSMtEXdIg7DhGIGfDnFxuA9FWAz29bxR298ibmpDg7QxSTUjCqWKqBimBTQwE+e9CUspX6w7
MyypnxnDKE0Un2k/Cz8dfVRbBF49nZ87V5xodHYJ3Prg66aTN1uxWb17/0VQnBa4biVSk5HmwMPF
VRO+2b+pIg37O9tzSX4QycG45JEmT/wbhzlzgcE4nmqjdhjxG90ECkfhjTE30EyS5dS5rCsucJTf
UcYA5HKDqIWSKd0+n8tgFfAnChrFqIXqnyFgKl1GuQl+YkEHS6EW0M1KWplrPKfK4+o+tJbP+J2/
dLYPq6r+GUbCX8PyhyGVXtagfbExUF5YiXhPXkqlo+dCtUpIIEByJifq06x5ulaftPFMeJrihkYJ
tPbCnEJl8BLi17RuhsUYdeZfC6N8x5BduKS8xg94RK5BCURT9rJM5hX58tJ2F4eLUeDgoWnsCfAF
4mK25EOjscy2sPoe1IBen+XVPzNZj/tke3nW6VKEdZtuI40pAy8dZZLiu12JJJ7oMloQAYUtPq84
TaT25wC28xCpkJtTARKkl8TBJSdPwciYTO8BJhIPJ9RVlnB/SwKVaRS+KSr10fxdIcW0/SwgB0Jh
BXwbdEHQ2qim9sq35sDf7eQ5Ycbordb9yHma8M+wSf6sAuW98PEHtSuXRb1jleedx5vXzAOdUREV
YRgUIg1bX2HRB6X4kUGhl9JjB0qRGf6f5QlZXpPibCn3O0Zuclu13HJht7u80rq91/5WbGZI1nHh
xrrPWNuAO7/kXfnhYvHuJffXEuhi+J0qLECrjZ8a8dW5GiqRS971SyRuM2Bxct67oKFqZjAuTyip
rtt8dbKCqemHHjcpZjVW7aAWGRJB1NB9P8kJu2PQV6b8D1KwbNdIK/Fmh8Xg/hWVpmZ57xj0oGCk
V71Mpuz8s+Ds9cXBi85p5NNdwPIc2itO3cBTzIOGDDk7BG+sJtgvCnjRB1OuFpbAQo0Qtq3gi0fV
eL1+j2rDC5RQPAudcurP6o1Rl7ZlFYkgIr1BMqfw/EbKupdwrnzdlbmDJsYxHGKpq9L4lMi0dx60
k+cWntu0u5ZAjRCkeaO3fzyCAcxn8V9ausNErlr9mtMO0GWPyhsqxhakktltpctq0p+JehjnRBKE
p6k4yKweeh50ngTJMrXYh7zALI+yxNYSWyf/pqGW+QdBGIJoTb7kGG8mgmGLq9xlH9RclqA4n1N8
DFQ7I5veFKXUu+LEfcV54YyEovOupm+wuEH5nCFbFInLTGBrmc1fpZS1qAN4CUJ7jUjr1gVLfmPN
x07SZP4bBFUKF+kessy/XRKiwvUG2tK5GiQA3X6ID/WxmdJuwh0x++i9z9uj5Gw+CKrBoWbn4A97
KXpHWQuWoAkwvTtHyW/dxFN6g97lyc4NPw5fwMoM2EL2ZjZD/XcHKPGASlgIFRXIFm9l/+PSYUEz
DLMZAmxGPyzGNX8/0ZNkc9KwehndQI89pEd8j7QbYHL4Xz5rOxeIZYN0HUqHlMQqUTUqc3C0JCKx
GmMqovyd/CPm2heT0RDakj42293LJF77QZImQzjmHOcDu104XMU+SzqJoJZ8wIJjrk3tM3G7wN4a
N+Ew6w/1jharJ1FKLwN2tcsMd7asJWniKfGXCufJzxAvLbzmJwA7zr51D1cc0D1kVEaFi/YVZD4k
GPOvNZAQel4MJ4i8dduDEB1JTAyVA1wAiHP4grg35jcMxY2mFQBX3tXRzdMpJYOZB3N2Vl9wUqVS
rR6L5RuJB9juUp+bVntmN1FQYMp56SAz8dXhzxjRUhymNc9aTXSVfz8FixsM+O84RLgDtTnIhM3M
uWkiKnIZOz1sR8F1LDuS2Jvwkv1Ey9eWJz83QTumduaAapT8zOZyDl69bHVPYslWSagoqhSg9Zl/
IQNWW7QpNIq5aPNCq8sjZRvSMSgs7LF123xvTayob4LcMJjZtqPibqW/eeQrswdbXK2CQvPVEyHM
Cz+pLah6HlCfmPb7bIemuExUQCDje++7AklRo8SzMZDEyxqdsEnt9TgJQeHBoWRBply5wLxqWCf5
9oh27tW1bD7AH5uDSRA9TGd/7Le7zqRY7BCmng7n2LkulQNyMjp2RKyTemzGh2YVjIVrZiIzO3qF
o4t/lylDN1PvodRPLjQB6gswpYb65k50MjSgYS7IgGLBYQZFNYuqGOcozqxyh1KkBPZ+CIF58FkV
n8B+uRmxTM5Au9mMhZr4aS0kaVva+Hic/ZPNPH0mDX/d0h+j/K6jUIkC87ixbnax5dBk2FVMPUkx
C2g/nIeTR9Hf7/2VVPeG14mHcHU7GwK+Rm4oZKiP+k3YlDdhSXA7w3nLjDdpzOdxiKjLJokkuYMn
7vFyZeEQDZ7M5Xp50BQlI/FBugMhqGmvog23azSQ4L/rpmjuR0ALb9ilPcHjBiGlsnZsL1s+9YH7
9XYoEUxu/uXdYKootXuf3rGRYDaqadf0cMnzOT57GVPFQdLmt72DpDvjybhGBhxnsEC69TAsOnyd
ipKw7qkAMIh+byJakM92fOyQhMLVYd96frRHooz/qwY3PEFjlh2h5Hz2+f7Io+efLk7iR8lQ9k+a
mlBEK1scGmymT/1zRjCM4j/Sf7ugiD9+SIM4pgBZ8Tj6dlc/8F03I1uO0tT0kGd7NPrg127C3SvX
tY9J9iSFyadwJYzGkRJaAiRtO73FcqQL4MuRcAkeyfVxVzjJSZbmp8ZvD6F4JMO0ArvyW5nFfKtO
pP+CVR02cIicxOkCLq7LVBkR5v9HYXTN5awWIsw6a7ZfbftMAd63UZEkz/aDBluSBE3Z+OYg0JOE
SuHtD0yPW1IYVUgCdVzeYaLfeiA/vkbl56YiVPefXRrWNfuH2ak8Yd5vJ9Wdt+1RUVSCY73l27nS
pSwIolxewz1EmTkUhsL7nQXJSLBC+TOheTJJeSlRNUhvTYD5fXxlNIZOjJaEpTxO7crQ8l7sVu/Q
w7TKfDiQmtcB9qoK0ZRy+khErC4uj/Jdfh4REfMBRQQoTGQTXTO/8Zkjqj4pZlO8jbe9HCcixXlz
zbkyLRra5KICAmeXWICx6JT0ox2TflC3cvNzj9YWdXiWGWkQ+XThhjJX9H51TeBjKA7l8mdVia64
Yg7dgH4fHhfm25W2joYVPvRj5/s3h6JDBINWi1gotVuv8qklayiFYNzG4fGjbTqTGYQLGNXok2MW
fvkWhkWPly458tU7CR1Svq8hDS+f+czV8ewut/KRqssBRIh9Ju7xY+LA6K1cDWLiCe3APtarcQgb
Ij0SDi7z/1zlIpwxSib9SXjs765a2e3uCJF6ThzEUN7hAiq5ruPnY0ihUmpye/g68Ms/tfI5ayl2
/j8hg7O1rnyA579pcy70Kh1YO/eDuoAj75hMCU5HmAJ+1tzWvbOoeU22fJhPzXmKsUIkhnjJQfGe
yqpcvmSAYDruHigmlXRKJVNuOXrtOiHYIT9y4LASxGXnmlE0vwbHMO9MuDdVbFsdcOseiWrNluzc
je0NsaNlokenMgKUZ9zp4V26izLVWgft/DPoHlMz0jnnIhEovV039lnFjFHUqnb5m2YxyPjDw4Eq
SknygkpzR4t9oDlw+uF0Ti7XPLys8qUobxf+uZtYGnNBGisLOujOGeREq2mQ6pW/gqtz9ybpThcU
cQ8z8AHD36mc5JFPjozfTExLyxmkSKcusux302wsC5Y5fX1IgZ7Lb3N1RTK4uRA2RQIZN4rvTMqg
vUizu66+6eZ/rjdkWFHa+aTCCcVM9yMjF4J37douB5VeWawKYqdIhv/HACd9hgjw/+5QBCwpjXUI
06QeWbxRRRGCRsQtNmjaijE67PVhgEoFuMn9olhH237qcp5LbZU+AuLVnztBDZ+bcgb/sN/Mo3rS
p9KDt6V0vr10vbLmXpyJWR66kbReufGrlgom60oB9RxOdf/7Ts5PCYEV9NTLTa6sIYIJJW5L4wXk
nCcZ8Xh4DZ53i0zZvde2FDLEXRQgL/Yi6n07Spr34YggbadNLKOgpUQuhi5HaUio+USdmQTGyg6V
UZWLeATAcITJCNLilOeYLj51LJ4ozAjpbIlSpxKh1d/M9UVhmxKn1GWuZNOMdm5qtVhVh4aCGVKG
u7NzVZrisS83U14pBtNzo4IvMS+vh+GcD0pbM5+MXrvihufY64fDIuJc6doqu1M9tWHSqPbLip6o
XM7YV18tu4/nYR13TBWgSKlwHQBJGkStTSOiSqS1kanKhzjpqJE44tSqkdakTUXW9X5kBlvkgKhp
fwnEDvRJjax2EyGyh8r2u6Mt1X9POpNM/1aNM8hLIHya/Rbpw+HxedZhizU3u9HYiLN5z7MJ3rNa
KsYZl298bDh7n+e30qURhatJP0oaXMF6QtbXq1q/W9azPWnd5Icov6BjpoyZAJW0VckNBVtvAwpj
Clxy+5f+Ed8Mq01nnK182nv13ZcZRMq28NsUicJKGRwAPvu3TCZ787Y9YExN7BNDSMgy5q5EFy3X
+SfAgP0PA0RKeBHpkmcnWTKsFiS4CTHHu1YGwDvVhKSJOPQB9auRIg+Jgmib0lIXulmtWk+thMKv
lH1dN7Rows1FHWUsfZZQN/geLAZ2qqOrH6Eoj7Xt3/0mSx+lfGPzQ5w1R9KCsRW37E6GTueMS2fZ
BfWVieuIfcDQvdhz5zpPohyr/tHJYdVcUN9XS2W+BYDgeXD2aUwLJhxLoxI18ElUjffBD8YQrrnc
Lqtal0AKQ6+W6OqtRTDDJ5v+92DsrczhGptzr3wk2Ov5AoniQylz7lPA8z6u08dOiB+WpBnlAz2k
QROZiwHQdy4jrqmrAMF2/F0WD3dQIpUc+1QPR5mKoKYq5OEkiKtPo3ZEi/6XFRNyokGeXkH5TjBf
Ahko3Phd8oRrt+BOLAI1dE5cZe2En3v6jACsh8IIQKyKAvDur831X4kSLfDQuK50U0ZQdIJT9/5u
bY06afCc+7rNwt18MIvoMhn1AMQJbrL+6TvQ4kd4swTH90E2rqKyiYtGwhuhYLtFIPiK4zeQ4L/N
dsA+tmmh/8erOtUuTpY6KJI6eA69xVjYZt/mCcXuofdwJfyC7c3LkXqQUUXqDT/GwvesvoSulW89
CLeDYzGREryAC454WYuGTZgj7v5xmtmfEwknqy0JDw8SxtzQoZ1fBytjesMYGt79MOtKj9kpzp24
ZB0vJUT6qiM1vXfMZ0deK26E4SjstLld49jRY4Po42syt3QfTW9S/+En9qKg050CKiEGyXlSXt0X
RzMDqcX6YIsOM9T5Jf15CNDKpQPqPZCDSMkKejam0y8Gtt789akrkFjYwTu1Q9K4Yb4bwQIhWAQs
3N9Wcju9E3lgwzlB56be7FrBv2QrLQWwmHIDFMZskP9uPtB3pXHKjkj8WufemGC06BCGH/ptBFFd
ynHBmISwJr5cH6ASPLF6vSTBw7jhOCP/8fhFSuoOpwBYuUR8WOJPjG010bfRh17LJKbQkzx4EDiK
2VUxq8klhZcWk+xSyf6IIMmiUG3hzxlrDvL38DxrrWaNsEuj4DytrdIFV9RSCXXTn/tsT8tGHyaI
BLwGBsVwDmLhmWhni0rh0juHgMyP6OkwTZtHDDJZ0JDOpKV4aSJbGdFPlYMcTnj5PPq0mJ5vVNXX
NHOCwt4839jaFc8BM5vKoXOPgH0rOWF85ReWuAp+TRgRv4vNzbJ1h0twBc4AnGDRlgrdl9WV3wf2
y+2b/s4nVf2iIa4PtjNUOdFHf7KplVym2lWvB8Y7gHYUqijceEpWVSnECQU4qwQQGC2A5yBIaUA2
rIMEdB2TNErWXmgiJf0SoYYx1V1gMY/JiILNSUVMF8F5AXIoj3/i9HvYCiO/XpqibpyS6tkhx4YV
4N3wRVpvH6zHmau+jYJBOeYJR7lfzZ0M+bpc9BWF0WP86apecQ0Aw8PXYywdeAFJksEe3gihEvIA
5GwuGmHU1bOckTac8tmVwt9oSxg82uyF3AvRSx00Pem+3jPMkV3utlMagait96e7bh0/os0mswiV
5Ws67TCTzoker12gUK7kbLuO44stG7jitnwn3NFjsbTeZKfVYAUi+3sxgtRgNRnHJ6P4nHDXU33T
HyyxeIMYKTaI0+Pi4cABXzyZZdf5QhelqXSuvximN1YM5bqoKXxhdgRTa38cOpod2nnrBbYTE7sC
T0yLrx41DE9QpECHUZZbsmU6vCZyMWy0v8tAtOddb32rfJQq7x/O3AX4UDAo7t5GhSHk7vUmuVJ1
+kDfWbxsZG/PlWZ4/2JM13HIeZF9z6ghRkjz52GEj2BDC20TVZcjLYSw5+TKIJ0BpFNvk+Go8Fls
/4D0iaXKcMj2mZ7HO3u0Qm6HB94NeQdHkfuQyE1hH3YR34WpplMq41609ky3+4Dkt/vh23mbt66B
yf6QApOC3jw99aw7VRR/LX7HdYh7PqBvyqvSbKgG/U1mqC6go3hilMoxFyHC90AvaRTJXH5UGH6D
hHZPHl2iZJE0kd6ZWoZvrsQgpkvms2x5IymM6Cs/0kl7PT/JGaPpDks88lhFS/S28v/gpbF8343h
BCduCSVv/gWLfYxoaA1mrU7lnQaXDmNMUPFYILn6REjGMAae6OQqHkRB/oaHWOfKvzL7m+92QBTm
nUZ8kCA9jFPcb0KihSvPSCU9nuPiJ/ejS1tPrKuoN5pHR3DtvF/x/0RTdeDrr4Bo3Fx0dBTDUmP3
2QdR8EaFyo+1hmg/iEaGA+ENUT8FaItMawPi/7EIr6mhB15nUFRGxs0mG98vN0x+f4gleU8H6Jxx
Sw7NbmSJB+FKkBg1dKI7kAeRYAC98llAw0Lxew0XbNkfcuk49PlKoiAcJ8Xbz77TZCa8Hqj2OsGo
+4PXxdLEZD9MUFH9+r1uhwAx3sMUtnvz9vhdgvHHxfvz6wFVmpsG1VmkZgVrh6T7C6vrqnoBU3RU
lYwI3pt+ofEh6Dv0ISWRtiBEJoVGs6IfgHGn6kEPa14nga4nyd1Pr328DmDSlfDxsec8E1NITCCt
6qeJfa4fqDGxEGGwY80cwmxj/fMjpLcl1DTbzW9sbwlLBvZEMy3zFdPJIw+7oX2dfEsJxWtHop/4
uXM80F8+ln2TUR0YkHD10eCtYsvbAJlnJy1J2LXTGtFqpQszW+y/tIZVOW2XgPHDWEPF1r6yZEeM
hufTqVnJqwPT39a/0EnuZeHOUPUZTCBxDohx2BRBuX4txDpvs3x1ZRfxP+koXA4dssY8HVlAfRyU
dTU/Mrznqu0togriUwgK89AKrrq4++eHw2Jczw8oF24Ah7+nK6nsbZ3N41XfQRiQEGfXjqIMtPA4
7Eh3OuLLLngkYXRkl9aIPkBSrsJMB+PdwSTeocUaWmpoLnf6RLMTvYHBDyMuUwzy2lMsIoMxvUCD
QrOKRXQDEVWPPzkw0wjbhCVdYvDMvqoEtNWXzzUlfcH6Hf9oCwezMY5Xg76tzCcCO0Wz0aKhJQ6S
5KJP6UrmPw0F5wwUc6KMXqyQjN5ppFjpRzZ7KCQBlJ+rFxo69zQ+eI1HxF3rdzIRqGzNofwW6CZU
ZDSYAIQ2w9NEOSPIIcSW2cPGrWeGSjffwmvO+mroJMVatSYaqBIqy6GVRVkLiYasntZ6VFud4ENd
4H24x8hBPJJT1YoK0RNKCn82MsG/rZddId/TeardNK8y0sayhrulgjwxRwpQFxzq/EkQorKjJA+I
ebBoGitYM3h7e9cUeqGSzyFTavznC34/L+sn0Vh55yATi1U9evAt/hUnYXni2RpSbk2G3iGBXGrt
MQAeRrrCzeqaK8lu/zRGh7YgtPPTu8lyn7nRV8AnEhVyr1K5XUwQ9BJCFR8IuoXMA60MoWfOX4oO
9ALIe9V99uUopi/12I8Q37m8Vb03q2r+ufVCYLva6z62iz4ky2m1TwOcMWOtfDXeY04pmbEwVjod
VNGMf7g1N/ICE9Kz4lpq1tg7zNILPLk0uBpI5AyE1aom8kfUWrvJmD5d849nyKWxT58Hvq5MPsdq
0lwPbIl1DdfaH4Iak9emytai9UC5pP1vpEMW7XQmMO5cs3KC3Eb4+YZ5PDRgvhK8JZ/zfY86Qw1w
CjKJCNmpjp8QCG5LNzahVcALSjhOG17+/UQOLi88TMxOM8CFFV5ac96bIHRrBb32ql3R0p2ttqlP
tVF2L8Pl27lHLWyQZjrq6Aarnd+HqCsv7o2+E7n+8Z0NzOagd1w4CB7wflKAcOMGAbEoAAUBrkmg
5lo3bmnWDVyg+Ao/gr4/CFhnVPrzY5vj0OPBZ86duQOiF3ftOc7YEd5WHUungsX9wa+otkgM3fV9
XCU1/6nOpi3nQg7mAkxpNlxQoMFRQjiPgK/XdUMgSZOnzjtmESEopbW+SxeXQSNpPdQDCI+ctxJq
4vDg6If3w+bBDjgDsGMTNSN/U0U52+wgkzIyl07XJ8fcIFcs4wqJs1KuguRAzVMaLn6tZVLeNFm/
KKRRKrcNSgycgxfCUNkkixeIRMLvfZl5Xk9nTVUt3KYj3GRWQXqYj7HR2QjS5yEU2nO+AEoANd9B
ExUvFeVhTepaDvgUAWDM4N8pfhK3IuoyDadwsuO5ZgiilbCA/NEdNbr+p74vKLAwtHN1DuvYKPTh
Apgzhc+zDW3lo7Cn6OjfDI427PwOUXNLB2XKF3mFaxBo2Gk+WhSSQlkHFEQdXWzxCWGXx4Hl8Cxd
4Gtnpv9T8HXPq9hL1UYQYPZFVqjh5Z5IDtyIUT7ZPXhA6q/fevE3qyF4pKq42b2sGemu2++M5vgX
GfIcdQhlAmrPNV0FryywhlXdHwdxb66RkFf5+uBubk1QQnebbG3KOV86k7kJpR4e7FndTypSgdG4
lbp0HjiWKL3ggQgmIMPnDJyEOBfcfPsDj+oT6vRqRhPED3TAY3d8Q+1HPbUwSED9bYhLSuTFAzQh
V2J9pRsX/JKUWWVKkviU5/KvRP0AJcnM0OuXgiwvzhaPGGoYBq0XUMmqCD3W1zOETWoK7sUZUehZ
vyqK2aVKzRBFSTRRPAeC5d6LaZFKTBQWNwrGtlmNiiqNGUHiyyckVwi0qcof0I7Tc03q7fKYyqMj
xpJXvs1X5bCqUkR0WmTAn9/KoxRaFm6+oPqrgst+LXl1zI/0aQT1hBOr2qfvSfsD0/g2xPTHltc9
JSMrHwf+I+SkHolfv/8jIW8jqyi0q/2Yd6pfhiQfunwGRdFJ13rUMjMx6OVAul1Sjr85j58klq0h
xnwHqJfx+/4SdrUIQ9j0xlHDdQk4/Z8CCDP4Erknp6gR0jLHCeewUXBK0SA1l8DVl5A1Uw9AnGe2
TpSHNPB/CFOvfhS+iy/5WdbQc7w681+UELiD4SJMoQVXPT49LJJecuvZMypgAFDlOoKObwUTkNtn
00jSxg2fq41duTkfH1Nhui3tm4FZGtE8GuFJMXH4uAIeuN3fG5N4+tMNbBFp87NVcEROQRiJXjvK
lZsOs/dzb/3gxgzLQY82PG7KD7APdyoIJemq3KON+BGlWF32Ax2/yUUWLMha5CMvE9nQHqGHL1Y1
1xJVsvHmnzIUWLINkE8r4nYu8PTk5VS1qldpgwf8YEnh5xDjMboDECDJxjBnET+qqxJEyaHAZMJt
4/S7Bmfrmyefs5MigC1ooqVxsenIzYTCids9Sm4i+wtSOUSFHhRIu+pj5KHh97IfQiJ6bJeEaZTS
T729S6Q9lXkK6+WWgb7vI9TPXr/vnkdwj0Mj5YNveQGQZ0WGvcKG0jZYyCvvO7BwLzz7lK4XxdNH
enyI2RcxkrkAizpg9UWGd7ldyyEctH0t98yashTHnAeQlTDNJWp1XCQU83UUOGFAOvIwkwOCPtAP
thd7QtUwITD3M3TmIGMig5OIMEnsZU8n/GF7GJOqtgPYGwBLw29X/qSd9W/EFexIT/6cR0MPCq7i
KzPWaDOVF5tgvYKIEUjpYn0vAolaWToPnCe6Ykeebr68kYJBbP8bG6JqfXf0+lksOlGw5v4DPpCs
q7gBXTLx2xZoKTQm7AjOs0oNArtRHNftSU4ho+Yw9ELyKy90+VcEt7hKycQw+yzhv15GpNzLGSZD
yzTjgePHl+snm2L1lOsd51X1sMnXuAUbqW7QLzyyAZAnFoVFx+mCi0kkh6F7N8yc7iBXVbuCWXYM
vQXDpOpCIs1iuI5OV5Gd5hxcn39LNmX7Ip7UKEY6ut4KXOann1PW5lIGN0yq9ieoJ5PyZy32wa/i
bCTChfT8G7acZAcwXfLQF74UOlCBREwEFTgwFQiMJ+fLlA2U/eLqbeg3QlwPjab9CMN9Rbuungwh
9DiCZT9HRsNoyyKgpvX+9zDJhSSzkGSwG+s/TsgUeJKcY3DZYqmYLIo127p358N90kMIDjdbTiEk
KVGcKazRoiJVNhAVRQ393fVWmYoNmQ1Y03HGfrlWP52dpv/gLsoPgcm7M8ZWwUWhGUNJJVQzvBLR
N9gyDiEQJTry6s9v4qXmNG4m4oWFiYu233g03M5Z2fbmpPaOQ9eTOsrf/q03HYJkfZJ4sIohGaqi
s1vWl2UuPuGSY30A4xdRic581RcIoa+fqvRF/mIqF+25SOP9qDY72npR+63iS78S4vE1qN4u0VwG
ynvrJr9a6tMBZY5PT16qlaELQapFib64HyGVoAkH8+ktSFtCA1WIhQw4tdB+O5hANBI4w6nDIYxF
urT3woFf8kHZjmey9PpGb5OG6SnY99Bu7EenPmUeximzgOrTNO2VgVCMFcsZiEY7bBuRu7Q2n7HL
QbKEn+DaL8RX1LU+8QQp8R8G0zb8LHyWsREJcQ7Yvy/7lasXNT8F1PW7wpk/WgqpYvladthrzQVu
mC9gSKQqRAqYtLTLxeb20lojm7+NLRduRaVu6BdNP1IStZH9iLFxscFLPQx/B4/e1/bGCg3Ie1/i
WP++/BKThmpcAWvs/MgKongMg7chPjJOgByqGnv/j/B/tdVDteAtkH0LTb4Qw31AcIqjWlfOLzAJ
FiHiAfcBPdgFAWwc9nFTTmbktyFuH/+oL3EZRPKr/oRmbYE+9Dy06sfGGMdEwyUDg8quKsx3WuTN
j9qh3++4M7h8dIcKyyem96SFqp779WoLEa39fzpss8/rmk9eYAdAx6YXkVDI2ScCPfcQeLFZl8iu
vW6gFd+plGS31V/f0KTPnHht9/eSvntAfrrfpP+4h425K0lFEWd5CpYsUeqObd3pkv6C5e6SB742
SCmj+R+cUq0aI1fGsJYb34weFr/vdQWZdwY0Q8sZ4XkaKdUF4DNk6EjInFu7o4ZUNp7WC95PgOYt
i5oPVOOXqcy0BwDmw5Ub6wBUqdvQIo1Ns9q0tRGWpc2u/WNKVQQUy0L7Mv2IXRuUb2eZ1rdcRi4C
dJIlftW6PccT50w9SQosrDKC1PNyTtOXVh1EInL058JMhM9zfMxNMXs3ABfTzbtZmYtoBTRI6x1h
POfy+0UVZFhdGhRm/COW3tYbOKME1ArTKqkssKt1CkQdN2h3NAY6snpgYI00kgEk9YjwSSLN16BQ
T1j9ZmE+kFOLKrX0J9PrmoEsJ/GXu/8IsUjVusm24zPv8KDUwcMUWoUUcvPxX3CgaRgYWrWls10H
VfrI8qpANPKQGwGoaH2e0+r5btHTbnkepHitOkbbZflvW9xrzr1BPaUWSO+cLKARjLJRZj2n5Nu8
q7zAQASQ24Gt6CXY+p2DHR8cE/57d+a3UGSwOvGbPqCY7s1nyxZzDyFfC7Rm2q3eNWNKn4q+gImz
P14k0QRDq/OngoPqCNRTzlXXS3mfl/SUBum8HagcLvYBforx9tI2DFUg/BBus7Yxye9YX4gHqEb6
hWKu8WbUnh0B+0KB1NBE4f9TXruVTI/4Y370Ccub3hsT1wEVuenlVmzNlHZx1sNj6prYVqnSMKXz
7ufKk5LYg2YMFw8lm4qrJ9GPsbX0dWcY075X5E5nXDLCbRMliEVsEnwNaMgtjOefnRw/tz4PwE/3
aQiJNlQA8k9eyZYRsFN7Lzm+B1qfDVRzhIyl8HAuWhrkLYe/qIjJaY05Lg4G9QDGS8mtl1Z5umUv
CudNt2mIfxeH83gZfA456zGHJ/qUi3HBIeaqp5GPbCm4+bD55hTOf0QxbNm7PGQtaQRPdhdnKFtk
ShQGguiP9AJairNxsdu4x2GuJQkMKAkyeQxSHcbMXFnUA1l82DLCRihwlIxZgYUhd2n6b+oLE3MH
fmbfdXXvHGpwPcrFLRRJNWWMBCEdfIePHkPH/hCPJX6GCiUH4lro2uvopWoPESs+3SMg70km0Zu5
E0B8YfYbdJBHxX2fVXfF8qU4Vvh30WmvsdmvTehdnng+/56t89rSFNJlCI/ZCUbxD7SKcxa0DEDl
iMJr4ee/KhiMavYTUEo0i4QMnNbvrcA3uRLMjFkOn2rqSQUnin3uL+SFzw85NNLhQ4vKkk8Gutm9
VJWlda6emkJXXHKqNjbOpnJVJvbZBsJpqp/HjzXY5p8rzIyMRB3NlEBJLVzXH+fiZ7L9nPW/u8B2
hGNis76b1WhRpdC9hp49d38tmnwRB09Xdowo6K4wGillkiHGvJl2qBf3DHvOkA9hH7fIXGJGmLbH
V5pikJ5Zyl6iyb0CWP+MIrZPhiE9Z2MI8IvMdGbEnlDLQzcNGZJNUW9e1KertVD6gSeXvARPF8Q3
vHjMctTthQQPkxOcsfL839zx33cKjNXPSyaWAIfAAlzASa6mza/5Xaru/bkKs/wx3+zXXPJ8uqeA
iOpOPAaYHA27+RY65UD2Jt0Ddy92o55tgBjXnuUQJDvufU6gBjcfJuZClRvu8NZ2XkaapVZaFXpJ
3+Mkck3S1lkCpfpkObfv94WmVC/HktL1IsNyZArdW5BZxPd5PXJUmxQasRvcRqvmM3d2YIQhoXEP
3JAUjmdcssGtcesxs7hc4JW051SNSSIBsVXoHvTovHNniMnxKp/Nx1wEKqb1VXFIDGiMFSSwouwU
XAUr5CqTzJ1JqY4dbS/HH/WkxnKhEZMvhCYr5aX0E4hz739scLaDJ+JwAND5K2586g0jZU00L+U9
zTlb902sbnpmvCQsxG7g7TkQzqJAPvcBToajan2mx+nZAjZKqRfSaZ1gl/eXtxuJD4/Sv78pp2gb
QmXlm8pfpOWovjfvD0CWQyHbgscoSYQABvKCqXH6My7nk98ADC+h2W9F+4bpZWPbnGXqkwMed1vb
SR/jm60M/iiiWq7zz/hQfWPp5492w6byJR+gr3qsy0tAYJemF0OCLvPewb1KY6aeofhh63CwesIB
fjaBM8y+cZ6TSbty646NJ0QlAx+r58/aH4F8c+4NPd2XVDRecHFHpuiNAY4H2ClS5W3W6/jCcJFl
/pJfVpMRlbuXlPmRj/Z+g2ZFkA1b63CkAqU9YUtyBRiqTmaqiFBICEJXroBymy0/ZEf15PPbYYy5
Xwz7wtChhzICzXgx7ehWH0TixsKOWGlomeZSEhE7N3vbjuv262WaxyTdSznzst0/endmRn7Comvp
cPdNS+3d2enqUnieEXtCjATP8zVuTLGaWWjRcWStXgfp/h5MTBwqWUHT6U3hkGeEzWl8OckB1a9b
+CRFMLhDBK0aleVuVex1/3f56xJspY4CvWKpqxo/ddWvAz3yyShpfkLIyMdnE7kowLlAk+ubN7sz
SSKLnjiuIwuwXqFVoYEpMos8jz3eLkubutvXVjzO0eq7G7deOOY5eB0GVcdjJGJ86SmlZ4r5s59o
Jw2se9lo2w87hx+iU1ct/01y88BAdpgh44FbLC2RIsqAoliOcdFNC5N8q7z4628/3RgxkYnUhNh8
xGPWHAQdmtPxEwb7K28h2F1II29Sq0H4FCML5EvUweEO34CBRqjnJ07lyfMRzQlyadsFExv5tJr9
QAbaIiTQMnnQKLMMISKoJZFMgBeP5VLKcrTwCF55maSQ6moavSnwC1ej8hh2OwAEcqe0yUrd2SvR
oGkibwg1ZlP2KdHZOu/j84JBH03CXEWOf0BYS6inJWl0gh9ZO6RR+mvpI1C8nZ/sIy/Gm41Ttx4L
z5w8EA9OVKlV76C/1qHLRMXXB9S7Pte6ltvig6LbaEfyLm2FRIrlsa7hXnbblIyexZPQwsUNyT9e
03edYfD8g5DcyRSq+HQhAKZJWoKP8hHv0VykiNX268iTKT4uwSVKzQqAylNJWG7p0lODRWSHJ/Nm
1oJ1ZiDZ1PRNeBmVqY+/loySE/WKFvaMHNA8+QuO4TFopUD4XHzCo7iNgu4w+TksfuFkEHpTzoZh
BSMbUPn3e/qzFui+6/tbTT3QM8HA7Vmxh8HsPxRJvFCfiqjhLzteAPc71m6ER/P+TOWBXhFWaGvF
qOYw+vIcs3WWxSBrkTOhMqEQXpvt/U50mVAtoERP81HlxUBqfJXpJQjtN3BWYR6jhVnQW//E2w/2
Cp3SY3Xc7i03BhBeMT94m3as4fG8YfLIC8tfeti6j4HbuNnuJ8uz09zwEE+kutRFd5pXlCMYcl05
OrBKnKep4PtmJy8P40nkJA79GwKd3x6HsGml6CbFGp5gvzAqUx7I546gP/fVGm8WNMwLjOLQYXSF
60UQhVH8qZVm9o/Cij76m5P22sGi9AVorBre7xx+Ue2lM82WXUQsS+oXPb/pRX9rK7iFQzQdeNFi
qETv3irCGFJ+TA5ZzmSIjs3Yw7gET2b9199/vCqdKkzb++uiIJt0QVquxgME8umqHrzvrjVwf4TM
dZgv+yQN214m3LvvFeqhE5gsBCks5loah5AnkbicV+xRJI/Ea/Ptzx1gxMNo6vzFSmtHeit5csUU
6s1yBu5FT90Dr/8cFeoGxmvUWqQKkJYn9rRuaBd8nXcO4XSyXQHMOBy5/SYTU0WdERc/KwpKOwnW
Bd7LrVDukvmlYMHrhyM5LqehCcqcfYg9fr/nBmeDcok+f/uORs7ae3n8WLZR23AzR8p5zVTSTE7t
zXigExV7Sr9j581bHnT+KQ0rUQbs+nmk+M9A7bs9zG63VHinVfYwmYLMllTtE0fM/b+6Pg9T1BMb
F5XsymnPePC/wGwrBvgKB3/MScjZswYXGDQsuCuAgLrcMaRa3Pav68StkSwBwqTNym/q2u1lEsb/
T2FLKSwKPU2+073/aDUy+Z/MrOcnty8bO/tFLh8IxlShcbKZMDZZS2gxubY0BoZ/ISuFQZ80nfEi
VR4O6+vWAeiCSvSr9dJenrhFxhKeCtD/1vxC6iO25svuxtTJ47Wi/RSCv1+PjX5bZctZ2EZArBmV
lpCmb+MPwcRjSCoYePKXCEbCgxHrGySNFquZNkCnBfEzsRHYxV0KtL0Da9MHta6UzwnkfCLfliwz
auiyWpzN/D6fmOZVKZxPdJYoluuKwRyJnZFCG+Fa/Zin1/WpNLFrvSDR6J/yz6sfJ3wjjjLxCVYk
BStknmkvYrJXweia3K2UM1mOpZ2v6PGD//1sR/rKbdakNm/RwdM+HDnLdY0XNAaMw8whsnmXNmSQ
noR0WhYWEsY/clylmR52RGyZAKkxPeVrhhhcwkxvNyXKDXF/UWJa+C0FYh6eCf79ye5I7ypvIZB7
AMk6qOsBY2CG1HRGAIwW8IaX4rN7xJp5YOoeAI1c+uUmMwHXht3j0XZg9JTyX7KnBS5X9qyDflu4
Up3hRw2yRfzkz0KcJ4/Wd4b5TPhuJx38SyADziZbZ9c1KHyTA6ZBWuaNNqe27aWYAXtwq0rYdDky
whru/Oy7LBpzD+wQxO8f/xjmRBCwCpnhbeHy3pSsAHmrjXTALSuBOamRGNFr2XO5HV81ZnDoZsjo
FF5xoNYP7axVIcPfMAZyDV/0n93vJIyFnHjynJ3TVvlK6v/DCyb3td7JjET6Fk/PE6+/tfBjfT6y
hp3MQKWgodBu1oVxumm86YN+1eZBv10rpZf0NDSC2yZRpgud9GjBesAJ1kfh+AiwA5EldrWBTRPD
U/7zeRqS/lZizHKfV+9XejrTet1keW2Behp1pUhFG3ayFW0jVudydwIaRGUg6HJhl5nmsPI6qn2K
Pc/RuP17mhmILgae/tXIYoyMtn/TOOx2TmR7Ze3Uv2UrniLOL5pEw+RW7wwAsfpJ92MBR3pWjmXB
PGpw2LlPrlSM+ZdZh5iULLQhPG9dD4tt3xabt+uT/Y/j8qEtUx5qvCW+vrrILDDyCIJvVRUxH827
HUdKaXD5jFiSC4ZRJEKKXwMWuUCBLEblMSwu/G7QknnoTGGiUCCl9TFQK3VhjlKJ3PXRwxvEvBAl
cj4f5XfRq/3QMjdFgRy8auSOfWzXBH+aHWbiz8wGZ7GGvK8B+dgrRevZX1/qOhjHLoS770xIe5d9
OaC4bZgDc86kSAI/P0vOsbUc6YIu/hQ8fh5DgV+aIeCBOIXrn56fI3YIN8ZH5bYnGdKG2A8ioIPY
9R7irWSCA+q8a/gf9Q8NUmuQaj99xRRHIlBqe6XDx71Ce1ELiSm7hVqJ/ka/ruFgWWVrcZv/3ntk
lcavvR/mkHEaO26yripbgmQhMEXXWz5oawwtuPX17SdHwE2eCn/t73CbbkqzwoaL3MeuUKMJZfAQ
SvhHj9tyPgXTJ6cUNEl2lytT8fIifv4F37SYAtzdqtaPYpAjnFALzw8IQNlZKjjbc5kW1/fGVfaN
FMpGV6jdlhKEnTNmxMe3LyuH8j6uNAWO34CrALSrCaPH2RHf41afFiqOcazXkA7JTNNdMZtTXVFC
ZLaCc4UufA5ifoXSWFBlgCzAk1h3Hxy91FST0IsjyDCzV2jV+HtUtQk/gYzs7yF2/bH2JjgJQHID
GdjWM3+8UuylZjttf/GjKtzJEtoh2HxqHBj+dZWSHAe1jIygc4kdNsrwc34UBR2UI2AXqMfmhtHg
K0VnmrpSYoMPLi/UWK0Ne1i52o3Rw88BE1nuNh56b6pKIxU0WRXlNcXZb0HQdKfgJKJRmdMlWsFv
GSX5XmT1AF2uelSQ569yzLruXfD/4FkjkQmzzMBA57V4B6C0idvQC/+1rbNp/Ky9zdbZtV07nXte
2jD7s3Akz7fhsLPooLwDrJiIsSTv+arf4jICsUSEBGRW+EDKK8GOQ6U04WjD+5A7V9trnd/aS/P1
zezvqsTpeofB+A/kk+deS/hCBv/tBPjAmFX65qV4pDxnUJsKieuN0lEmPSaQhhWOOMIOx4LegCpP
vo0Z1C+hbiTFUmydXDcVtLPIMMNAaervGYKBHMzBuuos35U1t9H1sqordIlJp4ReYEEujZjAlbqW
V0aT/zUKjn3U3i2zGuG3ocUpWK/tIh/D/VAwn4+NqVU6zO/qyZ1ikJAAedVW2DnfcTicI4CUa9X5
r7b5URiZ3vfn1V5qfUq6Sdb+eNlylbuPkNx2TZ5+0oiq5x7gP04fwazO3x5O0aTa+s5i4JbuOZ8F
fMpCXRXEri25tV2zbaJLhsmC63fRKdmzhzrb5CF6e489TRGdjRgn+OtBjraZOpwT+pPv+aF4YzTI
ynUDLOKCFcZuxijUQ+3co1O9pLh6nqL3V5FDxR4t6u/J5GPuV2Nc3RYTRPos4GVeJjsA7ZQf1uYp
3COCOBZ4BSGjvQLBnV7aCjNOjB8SDPLWcnnwqld5OCV98CT+YppWw9BYdIb99AzFODHgnhkGbHTP
PAPRTunotPlSZHw3LC/I7ctjxsJ2NBWxEHe7yz9s2zvXocVnZqSKGBG4m1Kj0uszNkIyNwSsykTQ
urDG/m49j1rhqlTpsmZs6iRhF9uXW/vx2nyznTOzcU+ymlnHJtzt4pv7Vwh0pyeWIJWz/O9j8KnG
Ve1ymXXFpthktRJTCJRlQarCJ1+XObuo9nAFxfk5Oc10ersE1gTddg6D08CEF+VLNFsBcR98IxNo
jMGZcjk8dDAt7PjK0BnqmcEcd3QLYVYSumgH/xOt+NU5VcfOISKTcKsZ0jyKts2WuSg4bSED2ALs
eLT+/yEHBKaCmvJomNnMBn8RA2cSFLnWLH6mzXtTJ6GG+jys5fv6ShuLaiMvvBpJPae6rgu0aE9S
kJiB+9xspxDKA568WjRkTLzu5ymYPquEy5vOQ8c7JoC0XmLgD+RUgWpcVyzoIE7lPphn0daKJHiY
I272rldfZ1L/YTh8Cqo2cgEAibG/ZTMab7LGHCezAxe1mq+gNWsUu+qUC4MghFmm0JrmaOK/NT6N
7bWMIuLiocLaEz485E0AreEZdTOHW8CzXh+4DAFyC1FOTfx9xi2BVSUQXih4eYt68VJdPrw2OAz/
dorbsS0hvZCV5uH3cH6d1N3xgyuEYPdu3IXfkpCfKBm+2jVsj7V3MX+m6ePFwhx9vc+XX2PNZcz7
a0c8mHxa1ezYDLCoDpZGH2t19BZaBYnj4cByiRo4eQsiqXUVFU50Hp9pJIzLiPlXwBgEIDuvJV9b
DOZCAxdYCuUXLeQJfvPyDlVbg9T3kRuqqqohbtM8cuUT+jhRPhpNg568kJ4E+lM6N07CY+p2ShEr
E7JUwkXGHULGpR1NKAylVb3opRIl0P0afwxryy10fcWbNHH9ONFRxLKKXjGRVF/+0KDxdTkH8TKa
4rpXiXcFj5zM7ieyM3YqdxTMFW1/+NNL6m63TTxxcQ9pSKkO2gU6LHivQIGOsBD1v0yWwlMigaNp
rREhwN3+VJXPg0W3c2fh5BYkoiBaVHPJet+Bq0ex0SnAP/8NYXfz4oYJwMjqszeTePqHwfLw2dD7
ngSu6K5Ocv/6Rzq2ZKxb6fypC+nCyeqTQOQqVNEpNhMq9b5ekHpnLD+4ZNcvImldcoG3Pqw2gqt/
qPVrZAA526BgvRaBWo8UASUEm+yAL9KpHRaB3T/G6UxBAUGm7VayQGKHwFWquGg90ZFxkdTMNbOC
JeCOTtWyitKc6YHBpFS1uWA8Oy//jGXLHcm05dHJEFDZPRlPbMJcIb5MV30AlZZLbtQCgOAmQCRJ
0+amtrMKNs/cPYMyMj4KkiLMncjmErhl8FOkakHE4i2ni+Y5yfQAO0eF+XAsJc4Hk0+XyAFiCIpM
jPFqS90MzhqyCq9o02GN4cEF+m8pLZHopf5ugDC46b/x490iQbzL5u7B/PsxhqhZlHAQWL9z8lRK
hCBfSuVGLJbZ1S7YywFEKc9pz0+ZO+kUjvg1idLjB/GphoHq3yyTTB8JGsiJRVGLTPMA1/zt26dn
rOIY2SHE9xzDfhnEYFwpGmAihd7bAgLCHQVea8gx2kLPvHq3JFpllqLAGfS+wqw/1zJ+Hgpkjigg
oaSuLGoPpZjFFYaRoDUgvpSkhbrJBJjbrQv0VrQPwoVMp+OPCSXBwRp6fcDGM4m1cy3IrtijYL5H
wZIzQmgQyk9LkPW7me1FdFAo2A0OelsJhScGZEPRd5SkQVtGwN9QSgBK27UB2dunE2UFCZBsKyAC
i9QMDjHjmBPvZKXWCUnCwcZTl+Ie6/+7/e3/WuHyVctOBkSGoVEyg1fkdaVPdQ1/l870Axugf/8t
zMRjttIA1PmmF0deBuiJ97oX2ZnDF4vzkh+gWWN5VLk2uJ3gmkzUR78W/M8/VVb7QFRMR7Y/LR0h
+fdIME1/iReRXGOvt8WPAN8NnIib18UGwqRsQsKnMbf8gAwItVKrbGVb6w7Sq1B5iY8yV88bjE5I
MA7Ogk2x/H6nTBVjmffH3HQ9+ZGCOEdLcZGIePtpfZmCS3m8rz6X7k5YNcfgzSw9HfLJQCw4Jm4K
+dj0i532XE+ybfKlRCfYLSoHme6JaGfMHcDHH8ykjAbv4xI3E83YKGz3aViWxoj1oAETDM195qYB
2UKm/4alQ/OpGYGgH54IFE2qsqD9Fw3SXrdRnlNqh7wUhiKnryq9ZV4a4h4/idOEmAqWLE4/LaMK
uBMf2OBEdjRTkygsA7BnhCOA1UuM9n1mNx58baYrGy+brphWDsmW08gWWuuDdFQRGmBUfNC3YGAk
RXuDluUIujfCb6inYIN3562+7bLAP0MZI9GEUsYkzg3m3f0EGME3ZMtPlcSNHlirMe1idzWNmZxA
wTeRkJXw6Ussct/qSXqZPoO9e2IzKiss/d1X8HlrI6rUoDpsim3QKkLfXuYmysGeUhS+gRqnrU5x
a2zS4z1aw1LpnrK3RNC4Tfkk12jHJtoXLVFUF8lxAIN5vRmgv0Eeod+zH+4Gpeu6WwQxDnunJHGR
JC65bN9nQC2C4wlNAggjDsYcsSbPDxME3cvvMBruff1gWhMIFNNCo1sLkWCISqTSSF30DKJlRos2
z86c1R1ArnG5arp/V2EKgniEC58YxahaU6H0HprzzCZ1T+bAqJV1jYtEa1qDuzpzL8dFLOhK52y9
+jkZDzK/BR+q8xz7zxmSNpNnD0DQuEg0+wNiF0uz7CO8Y/it2xPNrwca4OxzalUs/oHnR3kZs4pp
CmYs1aVvBuYobvcQRQr0AdT1JmbjaYlatqE/C6MmGC7ZEZNwCMNr+3JMaiHMDdDlgicg0u1qaicZ
S/8MgmpbJAEZXhFghJaVXwLdbgDEXAD7Bk7muFPu8VktcWiopzt0zTCd8/qymepm4EzN8Qhz0z7Q
BAUTru5B9EoFOIi6P9wuqSW5rOlVE7OqbDt5O7fjuin0/fnsdbzhN91W0VQ56JyRIhUMgqxUM1nh
YGe07CyVGOP3hzJ/Or9DtfA45wNO5gHYhNGc1S+F2yKtN0LOTcwysxpmg/VTb13yLtaauEvR8HDM
TBXUZT6HkCUWZ71QFI+8/gxYBNEoAbUOFrx1XmukP9+TW6/7mBYl9rapreUldEBFojR2Nz88lZf5
Nz23/ytLyqjHrFAcn6jepAXHJDLRS4oe0zdvzKZtvdHzudMZSfqOd8e0y/soP9Z6q8IpTEcx0cYQ
nwQMLemaHnaH6WHQZ8s6bsLFYSFBhANOkiNf9qVgHlLEIih377i6VTgr7o0j53YmvD+H7E7zpUGf
nwwVRW+KfLR3JKA+0lufwmZuJohfzxVV4lLrDH/t+Kj/Fn4EVEpOjfSfcGOoLWr2nLKJRPaOaD8Q
WSmg4yfCZ9/4kMBb85PyK559hYWrWxl/8VwmIL65gcsHBjUFhWQa0Ha0SuZnxtTmVaCqSZFQA2mN
M2kTqcXAIutQ5cn73m0/DAxnjnd4j4qCTXQC0htKuz8c54iGnFfUpaLqJrDXhbHxK/6AirzRV3C8
uuluJHXbTPepsxqTDej340+Q8DnPzzAz5uolb1s9Z0U4cXo8gYoYfDO0w+t1tonA8Zk9X+Eof2pH
3c2KIbUpfmRBOmyIAjGEjQmXrpDCzQEYIMGIcRxZCQXujY3zBAvTWNUvxX5/O03FuhoQW6+wDKGk
1/EUHMKT6c6dd6Xw/rT6uwnRZJEo8CDDybinJix7YM4fzP+ye+tkbB7Gm/7d5SF9H1kbuHqJCGkg
JUsyRzrROWTAu4x11OrJ4Cc7xbqjnaqFP/ADtnyb5O/9IKTNs8AxBt3bAhmEmH0XoOELZf9lst/4
7yR9jfkfKRNsZn6tF4FdCUZv7Kf4kP+3TbOKSpuBTxCGOaW7Jsj1OcLt6bNl9k4+0MpzQ1gF7SUU
P2S9VM0iWaaNc22Z0IkLS5Qgok0fshXfORqz+55+Je//hNRMKMgYWwg3AHLLanGu00P5XasbSWEn
ElyHSy7R58s6VZfJ8nei2zujmJS07EkFtJJuSUP5BXnTyJdgUWyMf+qIG4b+0Bz8y6mLo4V+Z15y
GOq2+51qIc6Z7BirmNs3VZrQoqqkb4Q4Yn0HdbC4OTEAX5mYz331auMTuQ0KiSG0UlH2vIM+LCai
eJxQomj2AV6jJCpd4YbH9qZPK9EbSCc2Q2N5Gx6Z45XEWTKROTukviRBrkdqroBEBpbbrsOttW+0
GYksdbMlIa3scwfQXFcSJFxtJf3sClLMvBc0NpmHYEw5dp5PnNGbKLHynWMWGJ87z3WVAkxw3oQ4
4OG7DI41DZoEFKT33NtZDpeMZY2LJAbVlvAOJsgbgNEjmkCykiGKoJrlFg+hzadrIayU1uMxmmXr
TsyYlPJxcAFEU1yhcbkAFlnQ6IZuS6PWEU+Kr4g3f6l2TWnhzaPnlMfQ0MnGcvx0C02qIER+WGae
Y08B4soOCmmeLcXHfxTzh/pNNulfsMiS525NU2vcTvM7CfNIjRUnKZF4CMd1zVphxA52kfeTq+d8
4X8z2NZiF4rPbGklLiU9rBHD0WF1bK9oVU5BnzSXkCK+aBy77PiSYFAr9vrEdNKyN0H2zdS2K6gz
c5BRsC2fgz4R5tM2LuTCfF50m+oYtl9zuGOcisaDprjwA9nFKzwIFxLOmrCdgIEHNroLG4hSM2Lp
hn6536tELpxl/yCCmcqDB4KAj55x2AG8/gDugkka2MM1p/XvA2kfvxsSt29d7UP+bjFQBdRskdhI
5sS3HgCgr0gL5/kx4kNmR+yrC7gXLnQ0hRxZj8ISIv5Uu0swImyzCvsj7rhIvfbjeRlPxYAgqEIP
5Bh6umhSEaRUDkMpGJUlBOH2PH7Gh6UdK0MMsaIq3163+vDn0VLqgEKMZiWxPbrshSQO5JWNMwrj
2jvuWY3IO1ETVEsEcKG32/cg4m+c3IE1pKBS+MmDWW0W59CNASDeJqNj27JlpT6R9hAOEucOInn+
wTgOXFQepVW2OFOsQ7OlkrxNebVVkcgYiiP3wtkNYyki606LnkYNEd2O71E0p8jDBFnbFiQ9Mukd
Sc9IAdc/hvhRqKuRgZBOTe3OncXRkRi1HxZcahnwQNPuxec8fYbbl9kZkVjS9FMY+IxPmnQBdZY7
KYxi1iJz3q4BAeyAxglkirL+ns+8HKam7SLQtkcC9XoRXClT/xD+YWnWGdJgBpsNfYg7iEBCu0Z/
PTNVfK9wDKEaunNGFtTSFW0Q8RMgW45MAOsSbQfhWVryNyoRa7YqJOpjrEHqx8cBGiPD1IzzpYsM
Ke2wAx7Dl2e2IFcPlMKOxzVpP+K4994dk2Wxpp8bDNCcPx6o6JPioxJztWRNBI/yB7g7bvFrpR7n
9lzscNc8TSP9T7iAowcL+uc+XefIpCToAQqiyJ7TUvuym+smNWbpL1jo+c7VuofF+MOhNS2guvUB
3A+t7LQKpvS4STKbBzyPwgHIrowFfJtOlaDn0ppA/9/iolBEhdvtQM4HvXnTiOP/587ktywOF5ll
VshMdmYZI+GgpHts7H4jTFqZ3JKIrWkvBLKdJ0RZSWJXomOaMgQwQxCcWic0GDtWR0BsdDI4lj+F
LDjvxG10yc69kXxqNp7IIonlYNHsqaeqhWf7j0dPCI8HUVJrkUsl1FiF6LgpO8X02Ufop5hTCevJ
FwgK5zHKFgbYiUYXtoQjG06T7l5uxaC7F9AulFQRUG/+ubRwWXl23Nt0y+K36nME6ps/E+KT2TDu
LFVIBRN9tPxhHlul1CXoNfq17S8wuPVFoR0OkuQg6qXH1QQqUEtrz4pVEtOsHNu2IvKAHz6vr2S8
skyGhtSKQln51al7pl+91syMMtRMtfvxCR6wTpBGFB11hciA4E1jFnPILnVTd5jNU3rz6JNbL/x7
wWdO50TFlckXKrGHmXXwnuxsOsBZw94nD0Ls5zNjlsiPPorD294+ka+ud/ps3sKr8wcnFuCjC4tI
870EwbHyzRDSGWUhb0AcRW3Yinb6PrtOZP781T+kVMOuRDVThNAF3zNwfDf7OYpees80vfhAb2xL
sAg2mIJ099dL6KAxrsWEHGikyBNm9SCx+6ER1/Ibw+CQJIiDZ8JNy8MLEmKFyqCLDmbsW0vUZ+AP
qsHe+SiMeAEfRz0JappzCjTtGb/JQBclSvuqAV+zdVyxIHiV0Ur4D41OgwkrCg57OKdqXywrnwTf
hWbFWjgNnuK9RhFfbR7rCvsiMUfrL5k8mkiX2zSkeU1mgb9BMPLmgZF0jJOgVMG+OKwV+kaxxIAZ
0N80fl4tiozvMwrLTJ9qEiSUHu1zBcgGx29VV4f/BN08aL8rOIg3ZoGt9qdl+N/CBKBLspoB/u+4
X2ydyA7ILFk6u+slUYVtbETVv//Q9ubYGclYyIRtnuDHqid7pHmDOGiWLTdwKq5DFjX9sk/whHNd
gmC2h12STV2kN9RXJpAc5OwK1P9Q02lBlwH4agzB8VmrVItA5t9+TAwLb9xuG6CkMH5KKHYhgAaF
4bkQqBQXcBlNlJWBPMGMQ4kLNdxxlyd6sRFIO9CAhK87KPbixuT0K/l6pdhW6OmyNl08Eyns2JBK
RfPLCydGKvyxmOLE5GU1ulisvORjOpT+HOv4td8F/Yve1ZGFr7nt9dglRUBJ0lT/bmrU93l+d/a1
7OjUGdaSG8RaQIfALygdXc2wUS7WhduaBA5hD3NiwHZaDY93HEaeFz0G9Tt8M07IdH7ir3ZMrUT5
kSdIOsbjw6Vnbqe5wq0t+4MenqQ+X82HHhd+65BEZJelAuIoyp+gEpTwq5sTEt/UmevEqExNDSie
5PpGdxuHtBMLyl/nhud29ZnZVxnzN6ri38CPuDSnkI059Z3wMP8ylyKYfXMawBnf0LEOnQfuYrPC
hdWgfBBio2BNFE51xdQK3taBQ4io7Codup64ruyvI0xk589hTltt9jXaPPD+0QUwVDmYa1j4+aD1
HuXsYpKKCzBsem9heX/zH++Sfp9nD3vzwK/z1WP7uiH+ZvIadvk+GjfMEslNUcEtE2tqk/ZzByIc
yKr9qmMeO9vkpCu9vCM5m+LP9rISydJ1uoTiJadpVDk08iDm0Fc4coLfBVPYUeR2pJrZ+fhekphy
/+3rKWjpvX0UuGc0362KKQrZTsDCT6mQCjYGkubSXwW9RWYgZa5zZ4IAj+aNK34lF77tCcx9IAgZ
NbnjNQ5CCUyzX/zvFDu27I9edZ7YZ5lYbtfhpurVrAMkLSCdAi6lFqVOqj0rOGUXO3N7Lpx19tH+
+hadlaaAjK0DoiFnga9hkgk/sQu8BCj42tWbm0HHV0hRuPDZT2fET1Z+nWqin59Yy9afdLM/7tQG
LfrjY3ge1psVxh5T57MtIrtVB5VwH74KY6g2wCljf+BF4WptqoX20KPByd465j1+a2A2+p4U0pOk
ZTjeZ3HSukbbvPq4bLZfNaqPkmcLiQ/mBqyfnjG3mqhHbxHA5kOXaMOu1noBNEpJay5EyXKesefF
1A4fT0MqfcJRc3z8u7XhLhj0aWy0UtMe9Zw0hOppuBcnW/mjI3CPYr80ovwtpJhBaROagPQsJpnT
ivdAHW69ihQ5qGNfyCn9YSKIGgoNJHYAMNV2iJCE6PXeyQref/bH29q24+NHRgY4Xw7VITypfIZ6
2tPVQl5hNTR3cCsam/bEBeIgmxg26+f6O7nP+tRyiSDOa+bKIGwhEDWBptekL/0lQUdwMfoU0gzo
AZL+Adhjl0Y6WXACMw8z5rUJEfmoKK8I+qJIrqfjS9DxqHtWQu6BOTRC6a1npcQcQQ2nifRL8OfZ
Y439Jfwx6LGOXsvU+hfo40A9zywZ1q/RhxRMSV1cPVpVgFtcnbd4dYXZbxg/HN7a30dVRYl7GQCW
pcOPf4eOYhwU8/NR2+0OxYWspYZtTHlziP0Y4RQNF3D36DzZPtWxBiyzz7G+EPP6N5XYAwy9ETBW
6bbDf0xtOvfWJwfFxrhI2wX688idmxyVUPM2UlFU4UAaINM4Gsl1/LOofMl974Pq7s2myMXEEtb8
DNoe2IrhexnYhrxXojMwNP/KA2+LRbRjLlsA5F2I1xQRkihGFvD56pO2S5srk3tGWGwkObxvUgBB
O4Qc62XIFNJoxZgv8/jSP+1vzSylAGsdf95p8H6D+j45F5mLr2BM+/kDfw82tHf70gr71EqROuHu
6lLCUjiv7c2sPlfa41bNw31oRbDA1Br0fDZAncCMHo8uvSdow3b2DpyIhZ5M5RWDWpckkntm7A+9
AT3/tXM76qib2MgPUE2lXFfLtC/GSog3p7yEPyEpKoFD3rbnFO4ksnPAAPHcgiGG9gUdbbCnuMVW
7QR2nq6tQBKkfh9rLQ+kf3ygTcWz7GxsdVnrEpEnFrJWjpANcLYuC82lQ0mgKavR661T5uROCdiS
yILJu1pRulMY40n4gThHBxMBCDW+lBZPphIxoXBSlHQfSV9oQ9/0D8t6Od884dH5YobZKbATIcPn
UkVJACAl7HyfbX1J8zBvxSW5ZZ7XC7Txr0rjXPu11/+qePiw2yyNiSfBejEUBW8GzZSGCOEMLmFs
R1ToOQGWfWPzAVBPoczaQoPR43FdYB9gOKzfAEkRXs1S4kpO4+jRXTYXAeljCX7Mp5wWfDAmKFIB
wkqYZGtwKynC2WXrDPb906J046hzkTUV8q9wQ9TDUvGy6QjXY///4GwHWbFRrP9xfmT3jUTRWhfY
eJMuAKN5bYiZuZ6XFACrE/nVDI32qn2lKB9t2B87VaiMQWked0YqkA6WzIcucJ9RAgaieospXYpq
v1m0m29PgHr04chWvAyPREcV3yYorucTCBm8WJyu52YMZHBFEUPlMBFm421reFWy2I/QMCVWamtr
xa65CU+Eoa/svtSimShv1dNYDhYbY0l2wGWz04S5Hy2XnCNZtKVnDyD9+HOeI/0SgTJC40OQ85Rb
b5Obj54ul/+shCw8Pwa/dAQxrlCYt22nkEZ0zePEma5w6wSWRsT2e07S8yM9gFfSiWXIYeV/SMx9
qJfrkIObCgyEZvTeU0/RmHjmPPWlmgByjEbggqAxxRzjGotpVMD0am+WNMrGS4S4Qxt9lH1K1x8W
fJMcugV0qbOFskKe08uZOtbgDGPS8lqwCTYCp3nMMR2QOsRq5PDNehy+c2GndspHYdJ34F3USfKt
/LyAFCSQ1zvq4/CA22CUTgkdb60gvAob22tnyr4mPeICotJYSDMqQi9H7p92r4SKqYcTIPI9sKxa
QOGFGgLwPfTZ7/sQ614ETutgNav2VLmu8EWGJKwoXeUwbgIOzm4DR38aOxCOVdKQokOyLdzq0owl
H8kS1L/PeF5IKtV4kn8E55X6hS+eiulbXMF3BSMwWkCpffnPrh/pXH1Ny5XPyW20G86oqkBudPZj
32tyd6jbsmhOHlBFvEMnY+C2xyRMmaD3jO2l0zG2CENPW6LXKxhH0k9gUOkpTknKe5CVMI5q7yLZ
46sIpiQbD98ENCzvPoIvuUoNqqjdz8zELWP7dXW1PPnhqdOEgYSH7yeQwM5ofSndAJlwi7urkuvm
PeX/cTsOVrZNfn7IIh82JbNEPDswx9qIi/tuhKLR4+LX9xySIraSGXzVOqYHt39oi0fB2ekgNtUX
G+lRZ8Y2qHvY5L0JdtfgYHOnpjSSUfp16/KSGei+pzJQGHFyIvIbKWRbnOfv6JtTujEI4FF+BxVV
qbTf1VhfbFfgRUM96VE3eHb0Qdtl82OIqnE48QYxmC+ZtWwhKZ5I+eKWRvmCMx2EC8e2al6pL+k8
NPuYBN4RNQrgqURnxnwMm80zHGYUU9v4UXqyXUdP7L0WMkfmFXUMyk3lNvdYPBMIqOVF6yfMZ0eu
qQFLjSrUmLTZuwk9zayQhRlAWcfMOkJ5rrRUW7tZ3YAk91K7+rLWUSRxaJkq5ftp6mjH8Wj9GltH
EbIqz4OBMbc3rLu/NupYy4SUQAXiv5qiLBeTD6/7TTsXVccVhx8G1kBEZOo217A012INJEx5YZ5k
/jUaxMMvfUQZWkEh7SEwsFXJ583dAJB60qWcz0GMRiezrs4LqfpYtXZPLZ9mb/r2AWmmT7k4WDB7
f9Kuh+J1n9lXNqUF7f/iBiobCoHC3d4LufGJ7tRXUfIQVvV277Mh8yxIYNeSnJWiuf9pYv9Q6n5V
+rHAG2K0Q7eGH8v+LT0wd4n9qtAoQEJLIQ6TA00HDekgywElwcrtKc4l2I8WU8pnE4OI4yaD1s44
0eAZWILAGAoSuCt8NmwNhpPGuW3y0D9MOa6ZHyOv1PsQ3z9pArYdVylgZmA1QSKYaqeDu4FClP1Y
ODIcQP7WdI9o+oroPnP9Rl9QcTemoan/XqFzRm6Tpeg7y8uChu+r1N6XAtE5QyvmaN2HFxh3ABMh
fYNElMxBpYmYjX9xXnLN2lUBPrF/V6VkoPBjeesYKW/o7exNKUM7S4AAOB8VRDoJIpmVr7qLs+Jt
4QSSZf08DFsIF/fogjKXajHVzPsp7zoG14a0o/Fr3rOKmKMv6Kwab6eQGD2bTZEMjylPjXXryNaQ
vfc1iJsH9tLUWJWf/NBbumLkwz6dovXJm9CbL2Vn8jX+/QoHF4eIdzF/iZhQ2mvvHo9jVsJhiquE
zltgC/Y6H2vUIyUdtckfkOOq3GX3UgXWlQGHBxrnfS3YjElXBt+/w8925ScjV5Im03pLf0Ef59so
9uGC7YyjHJpOS7SN+qkaI9JiQeEPwi5U2c5FUrKdT0Y8+o2ulDZQoQyCoYSQZEaOZWu7Wg1ONoxY
JBUuMhr/ZvrRjnE8SZWPfKnjN6BQ19DAQqu9z/h4S5r0sPIyQWDnglXnGWL6szUOhFUUAM+tC88H
Epjbs62TPfcVMCv95wL7t0qZ7ykaZV0s0U4IZ3vIHMHO9Dn3OiTdKhPFmvLUok0dgEpNTp3pDnCE
p4QtSUJOYpAKmRP55v7ZqCO8CPKHacWHAoxLXUASeDJniYdm9S6DPKszgarQ/fiJXnqYk1GovbMp
A3rRE5IIfTzuSpcTqM7rr/0dYQwjnNfNVLIzkz2BXnvReOk1hazhdnyNetwCsfIVABz6R88Jfcfv
bNb09JMy+I0JqzJu1yoWHmdvPfoF0yDEzd2rKESZtOaoo7pG1F9fUO4sBU4yRvbE+iI9m0VQJnbU
D8NSjuCkvqqYwJZpmXmWPn5PQWm6p87uF9oza9RM1z2kiRVICwVoCJVGKe7tUgnTCyocudPnYN4E
pVLEZUAK7UgsZAniHdU2nx0rLOmL3tsDupAId711pc2MalB6s3utABd+na1FC7hn6g6q7DX92Atg
5YzxLqzXPws40CRKak4K3xqV4JFX/MDYQIJGK9yR82GyWI3ugb5vFWD43SnHwS1kQtpP0Rw7O8sE
j7+jBE24JWgOtYDf4Gyl7MYYX8pD5FUgWuRTSQu4OJ7mAiH69gWDCwV3Dmd54Qjhway0/2y2rA7U
wpIeUKfkkkxkvLpWtNh4Lj3xUW4kPkigrc7JngDZkOjsZqEYKvLXBdEwy57QbxSFe0haxXVBdN6N
SSg2VtoPo8p9cWDkEFczFJKGI2tfr6FBrel0p7JjXmWO0zDrkZ1A9aLnnlLhbmVdk5oekQbQckgB
9y8EKeIHAn76x9Vhu4HJgrOFXeTqpP3zAH1CMXxBt9E/0/hzj0/rDgVZrOyNNnDBC4PodEplbLtU
BFcb3xRM/mYP/FdwnVohuEI4fwHbH7ygR2yEI+JAAcD8BeZAOvaYGwe3TGy0FI0WhbI9i8eVyS/x
LD7ixGNynfpgcms7mJi5N6nirSh9LwQOnuHzG5uup3FFMTcdN1OFc/RKHL0LHgUqUC0kHYOh4YaB
r2f37Cv4CV+VvWz6sL1T4oCijhTo6XF3OAiZpD5GtmrWdgOrhmymFpFlDRbokFfqdpPDuVwge8ob
gA9KpM+jJqqnZzTvgFypTXYBNsXTRpugkZTHAwO4eJlKZQNJdxlfwnDtJcaGNun//Ybv5I+E038O
gClH9naI2ec9hxwrprtbYZ8qQUwASK1cBj6/mv98av1yvPmdsx6el4HTZsnlOc920se9tq86IVIW
ErWOY4M2mfndylTCKO2OV0zrrORSBpGQV9Fo1v13Du6fmXTUVakQZjFfm2WDXjLvcSFAyZKFsSiL
HGIhH7wTVomvwnATsvCzGwrEy1j1lJWDYqrrzPHK3/QuRe7327reX5ok7KjLs9GPBIyV4dyAhEPQ
bw6l8HmBuuLpeO4hqOc3aWg/VgJj3qzbh53L6IxL8Flade1o6DWHL+yoJd4J42szxxL4xPd6Wkur
2foyf7EzJmvlN0MP4p8NcaMXDhLcjGL9LQtCDckFs1cdDaTSBTDt/9O/+RDAAyVVPGLYQ7b2FIXY
AzydvE9XSsGm0MsRO9wOWvx77tNmL0RUJIoYIGdtLVSSwBBqYeFF3aX1EKZ738MpeuDNQo0KZOqs
M9tjmOjosKlqeQxF23tfq/GjzwqQPvN0A29GDD00frRVpAwLfKjL4O05r2Hb4nqcv7r1QWQT7fK+
E7ePAph/cjC8ENwRRi1oscfcS7c9XPMl7wihzkvLc9VXTG92Qw78arOHkc6qBL3TVouhqR0qX48X
BfAyMSba2TfUUsGotH+dOtLRl4dk0ri4+4tym2rO2uGpy5bLgqi48IMiIvTC8T90fttReFX5cOJn
f1xv9ed820C6xBSTRC23HPVYXUf9MZoWA/QeY+4a3moGv4fW99MkY66+IOJlSiHNjeBey49bNto+
fcVJwsfH9mwmEsckWPyaZut5OuhvISx0hyiflAcFoh7r8zYQrwgua6yYl+zcCVhEeH1zqSQjyjKG
powLvlpyJpQJz1B7i0jKYPBa/M3XyESt50P1S+hILppRdViyDCwHFsfmJa4Bk4d1n0QA5MU+kCD8
/uIBOFF+OejA9JT5zJYqVfaycty7SrCGffKxRDMW8snOS3DoG5ZarJm8jPJjDpqNU13H93QBgOs1
GVfeyIz7rJ/WWjaoilq30mvUpQBF4/yarbGpgus+GiDYzhJRdLNSOyKy0h49CmOv6g9uz7p+lVbx
Gnd00XkXL6/obsOf4f4yI04L0q1bAIyuRWD9zNgU7fKtcLgtT4hfp9SHNA9xwGLMsvGnewqGS50G
z68dB7onq7gUuNxVZGzd+lCDAtKS/DM+PVXpNG9/0N8IfjTAftBlqgbkfDw9v5jLJ0dMsOskckl/
0RrotgD9zxw6Iq0/+YT9g2DRD4YA2P6w0WgHZQTV7OIJPluCwrFy3/h0C1nrOY7qn7LwLqJZMPhN
71vUQfQLwSn4GS7yCBGEg+UJo3/WcXRAPssv1zh3yldBbj1LaY8M001Eb/n9EsBDpKcZtLcDMBsW
htAS1MS6zMaEuGIcejoxcQNi3R6D8hOO6LNJJsfANw98OJOSWjq94S1OOxA8pEkZynY+bq5IYK1z
RsJ74K7Vu1s/Hl7Q8HjGDl82Zyu4V3Xam2wEeFYsfaGKWn0zEBe83LISozxhrMmZ6ivEoXCmYzli
WVefE23Pzzl5v+Jzka7Tnv7uLhvI586hWLQX/4F3fk94MWRHpT15lShA2o2GS6wvt3VC73Kkqjit
c46MR2xYt+2Uk5Uq+Lv97+nUL8d8161OpHDQ6587GGQagw6xGy/Nr2kPoGxmJGFEE1uyCE+PbQgk
jiaaaz0BzJ/SDD0AkJQnB/9BFTVJiU1PDt3agWuUMa/3ItULWjnY8NwEXndkN2rHAQ/hcj3ssZsM
e7WcQknRtpZ94wmDYwO8vM5WmVqIIov9ogtuEi6P6S4Wxw1FM9hrhzkzGF0jaXY1t7ICGxZkXvuk
YalYdXrk8yNvSKp4FMpOzrJXouBea24Rh/Mg2I1xXJ7xYTVJPmseHL5FdGU/fmkD4nkJ0oyi/7CP
Z5gJSklRcTuJls5sfYgL0/+ugM8wY9jyMEmXnsYrZNARlaSg1w3iilzPB/Rv73Vxkl35R9Siggcz
ql6E7HWuiwNpbBwhorXSfc51OUhkFASeF1J+UT9M6cFREKhdrVtNNqBlfRbdpZNKxZTQApPYTV5y
Wh0St0pV5cJp0aDEaKqx3MGEly9MtX4NroVj4w7nwEMCnynbdcRE9JO4mnjVccucGRWCbNaATVEm
/wTjUmeH68me+71U1ELSowVV+znvrV5SFt0yVRrWr+ne0or7Ziz5lRd3Cr/Uojg4kp6cV5SJXU14
gne4JHNSRfOPIkcSHV+SW4B469TbuN5MreIDdh9dMnCKoTlUBvsY7/on7i3xpx41LapEfkPPf8nN
Mdl23A2WRxboTg7fDbzMa1A7rt0Fo0G4yMljXC4b9M2jbdYvwwea3X5F9ypLgM5mV4Tq+rsZ/TYl
qv2nDx9VQ4LA1ky6gySgEAVo1YabEuMxijSdXgNAsW1XxH0dUM4H/as4P//wBzVbUKtI9l17T3GP
HkITiy4KFT0IfaSlthsYpUsSV5FKc1fRT4oJTjXY3Zt+zGVgu5dyq+zaMd+98zUGcKm4sIh9ksUq
LApHtNYFSnTB2UYAmxUcYBirmv02X4LDX1waT0Q3b9cO/UwlhS4yfJ7WLwfQVmiu+sO9xFWgXj0o
N2YCtllm6O+OVXTSVc2oHPXWNi43Eu5MArrXkXx0zovwC+aDTSypkYV+S8qKl4m+S/QvtKyoK8Rl
jrrZvIs3qgbGW7iJ2HQo+0bcEb6VUeYFlifFz+gkVMmHes0BJS6rOfY4kVttIUmPncfexYML6dHl
P4UAxCwQs+F3CJ3tImwlrsMUxfGyJQtNBwTMQ6frEMjM7vKRQEPP+2HhFy47sWa6KmurMZtgcUiK
Fnz9XWTrYOFMY1wK+WYGN4wNFBZv2qcxmTSHr9lc8m0SztNbM9gPYq1nCEycyKg9gCedDJ/MLnur
2d6l0l7piJ/D8PDA+MQzc163Qfvxz8XosaLEkzv6Wng88y+jAdsveSN0zcvoFQy7OBUHQKLVhv5T
5nwiLhHNXfa/B0aLSZQ8k8QeP0PDCgSU0+uvdCeiXWgVI7jAxNynSMUKwUqJPYmGvztwOA2MWWkZ
7/TLu/CbcWGMyRsspKmbPUOPhLbo2/vg2FtiViSICIdFIUYiUJICqAdvMgCq/iRGkqPaPtRzsU1G
Q+Xs4/6s7R1r0KndkOa9dubzTQaoRppuaEj0wh4EfNcwENTSISDEpNmcQXrso8esy905EK58c/rF
oUVI4QjZyWmrJc3cK4fXSZCuRpy3JDMlN4TiHPHv3Msprti1o95TS6tsZSja+AE8+NtnmkU7Daxc
+F3cbqGGL/CRNA7CKafghiB6XCuFKWh7HKISfU25UtlfYzRqG/CLu1LdNFPcFCLmWs5WGpRfjLbt
YBV0MtWtIDwxgDx2onlvE5mUZElGyODX87Qo1POz6abtyuMTQqlZ3PzWzDe4gGShGU4BGMXXvVj7
ym5SlT7LUEmDGwZCvb24/+oEj/RKkce37etDFwF56Y6tG4kJMW9GOowgUS/eMEK76hT9AhLRr8nt
eE3F7LY0ElOPjrR4nlXaO6JmAqeg+PLIJO03vLZe7etZv1SCyDxs80SMDFdMncwxfdrJS5KruHFD
wHQtp+xkv9/SBY7tuBoC/CxmcbgYyFrmyeiI9dwyAkwRx8HRNhkrGzYSzPNbq8rShNHgDAVZ4aRK
Sd3r3IaLSWlmEW6ZjUhfJQGgh6NL1DQEyS8Op3U38Z62SCAl+RFHZcazyXYbpc54JOMnWvklN3ep
82G9U5HEsPLQURdb/difGrygB+sjY7afPRu3mxariA17XSMZfJPusO3d1O3baHhITG89yp9N/9Y4
8mCRCsi14BHQL/P/bWHhMQBIdtK947aSqp4DKNGClBvvsHErA3uFFvp/pvhYFsQifidmZ7bzt7jX
6+POMqFqZe/5bIzK3UuUfTUS/RXzNVerLHeuNVocQwVVFj6gDe2HMYVJc8J66Rvc4IxvncjwHaRp
2Q76eg2uAYKcMssZx8DWpa4ikgXU1J3IVW0/N0ZjhCTwEgnx/OAdU3+psTOj1RBP0kbY3ZbttlxQ
Vmj/njnXBSX6QYOqzPWeoVpjq6lZCA53UjInYCC1j7ChSrDcVMBM58gRUqJdAw5l/I0jde7WzpT+
mOyYhnflWhp+baL0h/stFLQ3OIh6BhGVbFbXcqR2Pn2zWc6r1vN8OAa9k/by6UyCrhWkYDgd/1Pv
92QjRxAqBan2k2rFqjwn9wig7UZWmDnGIy7QusZ5v++0jrEFA9ybzc3oDcwMUg+OOcWYtUdMiwTR
JCo120EQVNzsoLIgcdaDp9RgDIgI8RVZ1JX3LijBD3aoE8hB3klY4M1Z2+JrsVm2pvLawZX3YtA4
Z9NLIo4ZqjCAi09pILOflsyCKKl5z01iA1DCof0+Q04BU/muPHoVH4l/vN7y2W26JCCCqj+JsZqB
hBo9DnVKA7eSNZHuRINuGC87AL3G1oP5WQYXrzfbYm65PV2OkzV6RfxaMQSzCnQX/UEK0hezWo9E
Ezzw78HJt/TZt+lgBWGeWpKkkLebEVYODHK0jSUnkH3yKS0MltEe0s2W5WEAkNOb7tONqTujq2Xe
P4L60gFK7yrt/xfjD+Q7aE609wF8GQDfoYcitm+t6niXzLrzBPWWJXlyKvZL02zwdz+rePEzca4D
75mleTWAJPB2TBsgExP/nB2aP0U5H6XpJpk9gXdzKo70mDdHD3L/LujJ/mBUESdTpjoTMl+MEDcD
tnRXqQrXQNrAyfwQgwSkwisPE3T66HybqiQeg5N6A6rHt7epGk5CiOtKDjAVtrAqdFuSnR/AHFMu
F/AyVfQb9Ts1c4+M4WA1mfzUgFimMEulNqfxmgvwfvd35xMywVuR5MmsexVXwRtRz81uMwxMUxXR
tDyVlJxAoEwOEPsjMelvAveuxFVBx8HQtVIUSGAoqvcqgOGxKE1IcjmgaoxB6XJik1UVZu33K2K1
B9jwmY6JDoft148+AouuXyOKYIj34WiFrTLN2yqqgYHDdwiNLp0DCjvwQWeJzjFVGw59gISGzcpW
qZRXGmr5EY6QAHt8vt4kKhM25F76A0Ol9juH4MabxQ9uQfWvfC6iR2NzL9f4wLsMEi1vqRsyRAIu
W/srMzE6Y9gYjxp5Jqjx8QrqIAVQhzrae8tkw8C85qhxE5vnXj6V7lCBI4NUz1xee3w1aJCdnjWx
iF9r1G2lVeu/QBvVVk4iyWqEWVoDioH+iTbIJyZZRR9t0X61cUE4ciwtqebL7BUZ4pL8sxAfrBZU
1gzFdUfbgSFWCHmrBCxxbalOUVoUrOSWSRRxt2Tph/pu0+BWeBfGRFsTyxOJ8D4BnPUnV9H6O+kj
vO+KT+yS2Pvw28HqEt3Taxrh2gXsHeT6QrNtLi+H6Tcyan9V26jrJdSVlgQsfq4pgWwCxRX/Bthb
UQtOrne/NzZh2ZiT1od1Q/pasXMSsHeYypqBri0xAPFITFTkQ9STTTX2yHisf3em95MBI2pfLoLO
zrEn+cQ0IlvML1Q/P3TDmZoc6V2Ma0jiXsat2HCvKAVh+O+rQzm/6BQHKpZW54JuFxLZs3cuzL7/
w+zDx3JpzzofB1GbLaXRXlKo3pqrdQ+g+ju7Pjs+Q9TccKF8b2SmaBj8oumvsAWWbF4f/S70QETs
Rs37uJr+J2g3HrEQXqD+Sql0KF1n7qggzFmGpEyWaLAdfuZDo9m5Xhc4j34cwXvQDB3+svr6tInw
tHII1i3iVqcnG6X4gn6jprhjpzBl9g+vXS8FZ2tNHNzwLP+Q/MKdJXvHPBQE+j4QFOBnbRFJouxf
331yAlIsDqvNyYW/a+er3bnLhkpPQl7lI7IIkb6rcl1AUM1oIY5efOJ+f2eC3UEdmSFYF/h/8bUQ
63O7e43I5t1vMUdnUvYwkGkmwoAPyT9fOfqooqMRPlcGjiKKGh5yyoYaK3YYmLHOmeMAzfXOH3Re
DtX7YeS6wi7IDdeRSYFzBGwL8dsX6lQdz/y2UnB2COtf5ZGUw248q4l1pKBlR3Ltj29YoiVQW0s6
4ZX3yR++3m6tW/xPvYmFwM0mwIB3OXfV4Py8qYbSvJZIDQj5oHQzevdUTgT7BZOyiR4LguOo77ab
a2lYSV31Hvf4Y7aGOYoNp/pHLR+4JmJyZH9oALtCyeXzeR6/vLsvrM+mAGpaRMjPfscGZzgs0VkY
FTI+K0+eitdEUjnFKa9+Ju6/rT3omV7d6R7sWwgRY8zTQASsc//euYz1QZX46KyansJ0YByJCrQ7
MLolgrQrlUeswP6AWxD/8rPq4Fm3grMIa7EW4EZUoevFChae74Sr8GP7kURJbZ6w+CYbX9INZx/u
N3sVpF5yJf9KuESAIH7HYajkaj+Jrj7JDEDugeo0RwP05mmOD0BEUDCAVo4wU7z5ZnJxtIDneJJY
l55WR/cnGui19H7XLbYlwvFTrgDmn9OVet35tFVm5a90zhpnVKyVsmPrPVEbb2maViRdJMeXG3hd
HV49UiMtHCjLXWUos+87itvt2rR7Cor//QXtD//I2Ng9a+Avib6D2Xtp9Nv262/tc53UU/JuSBYb
svbkZ0jHVMGqChws2sDP3DFcjthUdt7MJuGx1bcCRaR3iI8+XzODNxQn7XU6DiKA9O8YJHvdmRre
BXhvciub/GipVkiIRWQm3ugkuVRnra7yrxjF+PJUmbyBKAiEz1rw6DcvdYaWpBqoJ3bNvteinb7n
1yIxZVesbWjKxYBj6AK8hXVX7PszpEEQ8QS9GzreLtQEprU+wPnBhFr3PVulpoQXCqxWwjIZpu97
xmWB7E9vIKzDabya1skzKLCMfof+hcrn14pVQMLNDYhwtQyLFAhgTew535kiONy/I5LiGTLZtcKL
Hiic8c0Kl08Zqwv8zF4NBJVlwkzUu7waQk3WBlpUxTBqT1x9XjRzmRCNe6YVEOS6pFkU/GiuDbCw
kWPlw5NJzpjllQlXJlCoyfM3WQrIM6ViLDggTKOBiH9f10eh0QF+pO8oqW/ZA0Zcoe1L9u8kxMXh
iwOXvrq85KlisIwRxdJwf1Vj/WEzmApIEtbOuasuTBblAZyZhVxotBvywSSHVuEKQ31zhP5jddag
9beFGkAbezRbh7iV+stobZ8Ink3aPI7Ezn0xKT35I7Oe16FaZxzlYHRtOx3DTYtPSkKjgxOD5i3u
vdDq0b27jvxBU4Phz1HFm/Ki86wHdGVUOEjF8avivQNuMTrCZ7w+UO4SP6sshNsH6G1LrXQB2tdy
x/yaBibrBgdjKrjR4eQAUIhloF1YvoICRCyLW7Ti7UklqFC5u/OFoBZ5biOiF1IP6WdSqzDYSrsD
PnlHVqpzOE392XHc2AyC4O6C+9Nk8ZIW9cWVYB7OB1fwK6b9s3dSr1+nZuJWbvykW/3lhcvLq/UY
eHoHh76peyA2UyRVBP9zjur7WuqpjiCjjwr6y+VJIngHrkj8QaNNC5aoOuMLcz/IaxuyhyjBamcu
lI8SXwJol6vrbYnPmnatz+rAOpRUBaXYtyxXTCdEw6ThkMq/n85Ihdxxett5goXekmoxojLuLWtg
kh1whzZLx5TRie3pTxxsCr/2+BON9pk66+GC3z4NbTmJfQUSd0c6MZxN34pAHfyvkxOuGoHA8Z9F
M4A/1EItA1J0bK7y5GzFyT+d7X3hdanNrn1+BJNRY9nayVKU63E3swe7tPrNhs3S/Lmsq/3vgqg8
/gtmFVTC4yOVoQK4C1pvGICppYiHSON5WyvBPhSnJcbNXjSQhUZQ06qy7xrFwNEcwJxct6JojSlx
K1aSuKXJ9M7pep5yP4sFg6CYX7aWNR0xG+JD6RPG4fLWrvXi9FOhzBmwpzfecpMcVXWakhTlQrnB
CmxC0FLhnSBk3Oul1ANBMfWLqar4PurhVMkt8+fUeChzxn6yv0upRkXLPZzwWdQOId+PZuvfEHd1
djrdmQYpGZmSfbAEMA5tiYmDrtWylMMCvt/92J0tP/DvKL4FYNNULadhr85I20Fqx29GKm0Om8xu
JxuhCLgR1F8oV6BlQOIZURfOTn+OF/7pt/1MWxm28LotpVyj/avxdu+fQQMYKUuMa4VVXaVujis9
7mGCAnf9eHTyfwAZUIg4+elynAOR4pu3Soc7wBOSPIe5+ZLyBPCZrJbeEdAkNteQOZyW0fJe51KM
qWIeaEJDKPy0aFiJaud5EuPNz6bPUiwVwRHXwetfgl+dFw+eMmr49LP1KldjF5RQqIeHQqO0aAMB
S88iuz7ywUbFTP/mezlYJ9oqUsgPo4hq72gw0yjf5D8YQNGYwAijSzZkUTx8naIKPIqGBum0E6Av
9RoKFKMw4794hcVjULwBOQck8XB2yDsc1zjvwiWBeH3acnY2Cj49v8z6CkI4C5trbWkIFNwEs8RB
b70Z0SHmjDzDNUSmN9IbccrwtPcH5H+rcIrjV1MzdcyTdKEVsAdweOFCnys11nudaSrZjdpggPlW
aeWZ5ALnRS2X5hi75g3ZN0zoTWmmJ4vRrCmo8w7fDoyyexpfLmzEOEOSpYSLGixuUYRpvmPR2B1d
BY+ZWosB6SFj7ZWnVlwBvhB30Z+OZi35qhXnhqtC+pIe7vz0egYdWhJyWoms7UPvWU7H3CLz5tG5
zu9mt/ICzoo+nZ07lP2uTeZErrt4qrsadCcMH9ABKyrXHIs/0Bw/0pBW0/9G8+TmeJagpUfpbvQY
PLOP8+hZv7SByvyrKg/7tJUjQ+doy4+NfCucQtJ1Af9pOI/fwwfGUONyRt3VzUWoQNWNFoC6EKSU
B8eyu8OP1esAXzAVR00E2hQzZCasOIq4cm2/pGvAgpDIYFg3EYJkc6h3MOd8LnwX2WyflJJfVrll
abUOX2Ss1si3bjmqCI+hSDhIhe2RmC+MKfc7h5zo9ioMJogaC4GVpsc5xu1lY0iqvRPPcVhHxMUc
ddf3HDmXTqvMVtt/L+EiDNMU3c7Jgsn2McqQuQuBVtXIJ9mYsbI/vouS691mliVVumD/ehVG2FYh
pApoe2iWpRQheM0xfE9O9IkCg350K1Dykc7gJFXgU9E1qyJv3TBpE72KdKljP5SSDWaefAigNKs1
S9rC48ygO1gV7soU8FINNaWmSIk/2bwIQvrZ1gBuq38LdJV2Xzzl4kiU6rDjk+9bSeyZzzcsEHu9
C5GLvYaBTtH1hzpKLsANv8eMfzbsOrpKRsJJ2SkGEyo4zAoRVBTrZBAYl8ivx7NWFsncHtCu/6GU
ByVzOB68o8uytQ9UM00vdmbCkR4arIVpiuUWCWf+iSxhydgM1185qu3ym7wxEZSNj6RCElTy0y58
YMwCki6vXfTRFkCwY2n0Fw7gWqo//MTMwkC1ueGXPnB4hUzZ1ejj4r/Nhpqsc1L0rXrjazBzPvn3
DhkiC03MC/sxh1JGScfLlSZJRI39vSCX/j7OS0ypF1RUMAaq4YE4M9TGc2TBhLvsSxE98f8rWqZ1
xRaKfTmFka1zqZVGpQO9IzS8PCbW+5Dr6HR+enT/rwJFw4Lge1IsuDPZUuTnLRWAsFUZpO66tliq
3ZnN4oXSSO1yKCWAZOsUiAhDWXhYnjkafIkCsK6AqEdxbbdO7tO7YZjaFfaRBMgB0bcQdX0QgrpL
2iuEdxXgtQZmPdpOwdC6lgjJ6YVFMUfn8yM65be3pBh9Z3vPX73KLwWaX41YrM1wvoPLMM60+2QK
sFYOeCbGYcCXhfh3uB2/owocPk55O6V3GjIQ8p1qVF/2lfzwwRRozBZUZuOQgi5pM9riyqRRAQc0
mgvLSuU3r+3m5bhKjuQ4+LM6h9XkgB5r8suQsIFe94zUQPdSt5Y8EHjGrGIYZph45AuM6LUlIMfO
kCPRj+FGSW3GC4YifiesvWx/U7G6/uuGkJwksk82Wr26kVNjN/taEn/hc9xqstNhUZvQ9l5gZz3e
I8F8if7CGU30OANaH30UQs7KZikhvlkjie76RlfeeKrD4HWXSnMlLXCr0iz/TrC+JsI9L9hFESeX
a74AtXkLOubg/DP7+cA0uZugpzjphwiDtl17RBKsZd1pkfdgLZfk77t1CEsYIuhQxHLY8o/YQqrO
/rqsPtR+jMJQmteAgwJ68GaUan7Yc3PG+dOg61M2as5KK5WKbezPjqLCML98Z4ofGSLjBdvnfNtE
g22lfRYCwUE1o+CSwwOHkt/fioc+kX44byOaTfSmgZkJNcuyZ30LwO2EZz3voE1+f2ZM7+1knpKS
GTlX7lKInrJId7jCOdU1siyourT1dYxAkpp3CcXfot1DUlwm+POTh/9Ds6Pl0ptKHEntCIArrhr7
Tasg+w3Oo4Ci9YPYIz2vuUdcChOTnhQ/Hbm/xFrH4I7N8bTBHW+rvpybAAWJ9vp741Fa/QPPLsV9
RYOp4e+mXBEAFTVcnR1+54v9h168wS8xIUms2f2EQ+EHu20juelILmxkL7KKyT5X+cxeSXWRQfmF
KtbR+j5CXvHf3gT+BiLMZ4VHr1lrhrv/ydzmIzN2/KVFPxxIBAIU9F3ZYgSHq9tiZE8lxVhb0k1T
AoV+n//ZidJTHCsK6lrRhQWp4z0oQmtPqZ5Pnifj//Uyd/s8eOiHkxh0FCO3VW5ImG+6GhTn1x5i
f3timpec4Pe6TUYqAK+C63wQ7aMS1aZ+alj9JtTtEn5oOXmNVFqL5Z0C1rPoFfGUjeDfqAt+OH0s
obg1jn2p31K7/MWH+OhcMJihxExy5sIsiU0ERIStc2Qa5bESuqrS5aA5hl4YO123TTL3FSVr7tcb
L7c1Smpl5jezCHG0tZnl7nfThjsl7Yf1dgDDMvMOfv/ptZz4i+nGEeHVSBhdFwiSfTPgd4x+1yT5
arWbxtNrkxV0rGiS1D0tR7O2kRrO4Pe/UXFuxZlHZat4TjxSiXA+BJ/44A4Kdkt0c5ZxQ/Og9XXY
gzXLctu+7h+AJn6RxXVmtjucsKHak8PKTnewvawNHn0rJR1UaY4iXR2vT8kuRixySci39cT80DQ+
+NJmADJaVHqEmCjkv8jMbiBhUB4ARfwTUkxH4tAv+7fzciYZmyRcdfQqqhS43iMH3uYVLiqDmHN7
aRhMmU5R6KCRk3l1gwofcBLZN/8y7pOTwFg8xySCZFYSD+vXfCJ6dmJCMTe6QOTaOZcIMxMM4/bk
CpvqZG8ZLsXE+6JWnVsAvZ9gOU7kpchKeou6UUIckiSMRUw60X+dvD0u3JathIpaSPoaLErBLnX0
eP3DLyqrAsC11tSce09j23xCvGfaMVhdzScsjQJSiqTCbNGQNNvrCFUvt66rf89sahQoWs/2Mdog
uPozc75IAFrfKDrNvYk6HzwbdCRF0kpiWyuw6EwG8MwQW/i25MAhN90R6Le4MiXDaofJg0e9bqWb
5K0CRuPf9GU+tEEsUg8XGcugcXmSAkWVeBoMDlZxd3RDNICxwfzIoTF6WQsJBUrIh75HmetHn/VD
Hm5cy+qGFSkZfeaDpKNAe7+cpWgl4/3tp9OhkM+tU+gQeMBaKp7kJFY/P5M8WDfq8v6R59So6spn
4K0zBAGLkYL63OSJn8lHJ1noE/QAPJiOZq2cQKx0mUMvwN9OMDzjFH0acI37zJMGQukcdBp4P01S
4qc6O1MAJdsO/ymOkrKLOGWlxbopylSmSD8m++uMWiOlGHdTWvlROMTbTYn3kaUNRn0z41MJdFfO
nE+LgKv2pqqIsf2mYyLgiOU+skdaFH67/19XpwI+s1ttltTtJec3wd+9iRm8arNtlSVjVuedbbK4
bZ2Vp1TcTAVQLonZsSzqQQu/vBPt7+e/9+eACyzoRoJNl2NBcoog0t/yIIoRCEQFO1mP9NL+RUkD
Oer0WxBNWQ3HEWbE2AQAoQ2/y5dMQNnQhNZ9wb0mnoLGdNf/8hCV7yKICqzhUFat6aIa6DxVVoMe
qenoidHRpIOCnqZ06E4pevRRzN/56b70WHV2e3dHJZ5JwoR/sYeqw6k3IkoqYhanhi0joZbx4MuR
7x7s4kDpD1Rx8hrcdED7hhIQ8IyIw5wy07/A0+Ro9Udkxk1FKXLxfUTWiOZqPRBxQqXeFH3Secvb
PEBUwmBN6pZ7XrfQWjGlE6nJg0cHW0/wHf9z61/M6xjKZpYLYsV75MXLtoRss9/PNaH9fKhTX3OL
vLGx8zP7KBNq4popY4nD6W4qAvLULOwMmiIDgPp1f0xN+d0rGNhRRVpq2NHtrdVFJVvZyKJ0NuKp
S7mCO6T1snvQOJ6NrA2nkg3KzpwtXvVp9CpV2Yno8wPufGqFHD2xQKDupboEPIvU6l/rlnzf0pYv
oUda0OlhabdfAwac9iosiBYK4Rgw9vpnBPECEXFMDvhz14QQRXXxvyodEJ6nPTIzIAK0uegRTejY
jXchOjBj8RKh+Pjw0vlCDeeSb/pDitGrW/UqHJUTAZzE7gcdnM5WtrqjodKWRVhLehNsiyQFM1a7
/4QPMebcI7SwEO8flpuZkxuD8xLHL/ClJlITU02YMmlBroz8+P97MIYNPu2OxgJTkrR1gCwmiERX
3eNcHMoEwgp7da3iT8h0CLAsZdxZyHhbKCUf/JOdqMDKiKPP1aJBMbMjDlzPaswwHZMaRkhZ2kNZ
VNaXOtvSHUEPPXUBZKrr+p58VjmKlswPDfu6WZPEu3PwEFbu3XDn3TlGxWt/fsMkKzvZXTVzPt9d
gcInvn3AGmeUcnd5zD+qlTay1XBw+Pvi8oFEA1dy9ElZ+QYiUfMW84dKo2BBLlhryCBo8afTUtmP
ysW8CAodPco7d+SF1pRKRM77OWrlmmFH9beKizsY5YKYrR3/23S6K2VTsn1oXKNyQS6RR/wXfkkg
8GWTErsBDQFod+WrlGvAFEz191VLiIiwxN2l+yR19W5UsA3/PoD00JXgAYyZbvPeU3j7I79QH4HO
LPIRpKuA9OggalMhhDdfl1NywdV3pbStYAH0jqoDuc7St6ueOc3Z2az78MmnJ1w2pdgU1urcBJ3F
nWHn4OCJj8t/lPJy1F18lxvj+SSATftypwKxmk6iCEBuvHwxpN7WU4RIUZeItD1lO7gThYetpFb7
y2ekWEZmIC4Sbao7WfSv539ZPYFM3bfPoS0yYTvIJbgxMwEGOFqMGSkbwa65uXQp7M5WUucaTODk
WVK42fcmNjg2w8LAfULgtKpzte24TmlC/L1EuqH2BUUbHzaJlM5EYyTSnHK/wZ9/3c5dXKfxNtSO
4OZcJqqXehnWu5V7oCoELLQbLzsh6ToJ1XK95bY9jLdW7INvibIPdy82aa7PqZCMamwBj+j9DVHh
1of5rPB+8Go3mpTp2HUiLgt1NLU456+2mG8pn3AuSB3CeGP9muysn+7yr2QmkoOvARvrlmZ0Ofts
PtAjMO5gvzUJ0QgHRpJMjCwu2YsEBvd1mlXBBOqORO/wo1Bwb6RUehTdPSiYCXqQdxgGcfgsSCym
IPMZjFHNG/rpwqKPgyLh0EmyxBnND3/atIYeu7OlWCyV4v8BpsLL+eSrlJMcDlVUFxj20xS/hIhz
BHcmhtfYBpvckiLdLqE5VCMhSTD7sFcFPiUHYSb6GVMowC8H46U3GJ+7C70/793vcnEyWijV6BuD
2QN28Sh8ZRArpqnA1rodlqN+XzoE1GO7gMd7BJreLFO/ypsJpP9sqmcPC8i640wDn3cbjm000BuR
5ZG3alJe0RelkMJT9kbzrKZHYi3U69wpRWiDxL2sh+X43MuBM8u3uMoJC17BJqnHZNC04qcJdbW1
GKW4Yr+d5aqQ8Qsdo6eECNjoe+Yd1jq7xhIyId+TXx1zzn6gcNATn8zrmvq5Jb6B9BIqnN9RD5dZ
Sui0Fvg0neehbMlxC9FMRRMi+uGzzEOVL5SbOMd0Srzlp+rAyikV2CFdgbdMV1wR3nSJ+M+MBPy7
QBczGVs+VE5Gaxba/nevugWJmKUzG6Js15vcWZHTG8ew2EIlM7sQcZxf2qIxbf+tTn5FXJy0XwQH
R0n4N/bbxBuqbPlE26AVrTZYBhFkXvpxo3D2OgdjhvLzH2hcVor6MYA6HWFzcagps+vlC6OuglTv
Tev9LflErfxNGAgf/rmRONwRt3jnmGmXNpj53V6dkBg4R9/RAiNf/V8UHYBUSzdZg42cejduQf+u
Nj6RwaaftjIx48nrokoEIosf4nSax6yh3oRelTur5z8CuuNWAcr72VkSwAMMuVZH7f8k0d3Y05tR
6X9Do1MOsOWAgnea+GJtOajbNLOHpGVh8OmP1peFav4+GXhXbd4ZyLyPzWdfydI9UqBR5IRkqgzR
AmPaIeDv0cBqE8WXxW87mAYayyFEkWWIeCglRRvbUbZnAeJwU6B34mtgROF0BE6sUMZPSGlyD3jS
mTjDNa7vQjdXL4j4vNvhfvvprOitQU0ApqXH6wXgFX0YIU+jcpQiJhZcudaJRAkaEsZITcRUUepl
sSX7jDtPHOU8TCDI2JqXx/vhz6lkM754igj49HFJBx4prl6AKCWkvppzq5jGeSvvf7Dng6O2twHt
0FiXZyKdPDJmDGvruGlrjZ894ZsUJtKsXpQQnqKOqZG5C+YzWWhC/0mhb3bkr7rBT7zC0sfuAi7q
ShIwXqsBaos8HFT9G+Z2+3zkZzItmc39s/N0P2QJZ5E36cX3MAlLg31F6iTpEaRqxeHIbgqpSnR1
wbPXBIwFqh3Nw+5AqqsByxr2jJtlfj4FouXjC7bLdGG6it9+Mo83NFhj1xcFomtLOyDg9HWlK9Ro
Wh9Zrw2JBxmApq8N5rgxfmJAi0pj2loR73iqF8hBPoiDixIl6wW9ElJ8tFZind54BRynTWa+1SQi
lTWgKF7Pe4j6WTg4Ukx0NYuPnzhS66xCJnE0lAU0tM8LlSh6riMIOg3sGzOdTGKLn2V5pKxFT77S
/bx6OBdvTbJpQk/ARBRdRCIUYnHB8+mf4nSczY3tJoz+12ROZ08scuZH7hT2oaCxbtw1/PChJcUX
2ui5XOmQioF8BEYun9ZYxxUojXsk6/0i6+YDRXMAqGXhg1PRdrEBoKXiJ4JRu51Tq6iE7PNpvlnj
3TcVFWWYgfEO2TEoA1vFF3cDcVo1t0YL+0YANdqTYwP8ddqlrJEZzUWKfGGEOrM9H5pfMTYMupL0
A3tyt8XNBCtBj+GIb2eX3AKyTwQnajWHFdyLmseOB04UV+SyaCRc6j6/mNRydsyRRbGi62mkgLyl
yjFhvJdVGViMbUDz6145xFoR2lt/0o6ycpBWlc8MzoLlpfttIvZxJQP8NeqdkoAaYJ5PoeakksRb
tgw+IqmLZk772YHb4muVQmgwkq0bnvcbE+rO6TBIXmXuGBTBr5or7rvQibZBOrE+jAGlYn8DIg4u
CLrYoQGvNOVKc1SqiFRkOptrp6j4xwKkVBPXvFb2iJjkkxHve3EnUKH1DpJVrXFWOH+bC40VpQrO
E4aefVYzECd2dEouYaeujUPSkhgp2eEkmXNV2/MP+JYtX412AM81MIIOZK7gJrDqMS3SjGGeofM4
LbvVNzeWPI/wYiO6/CkVWLX46b5Efjo6sEoSw3ZS4cpHkP3Q1C0RqsxTsKmvtW/TbqijMARtSWp3
f4tj7F9ZFM2jW6lxPGP3osU/gn9H2ne+DQGADjrVJ1V/zybZPH0UFPK9wmGI0AmMjmHW1lfKCeQ8
jXlVGiBHX7QFQWztgvf4le/N749GGMmuyhdfILJKopn0hor1pmBc+tAQtd47XWmArN/CUm/2HXPb
T39Ea5OUdlpefUXdR91+uMB6ba4u4TdRORXOyxXDk8bNQc0MXe73ebdg/ZU+2M3pRPlgHa/ufB29
wNJHrU3vde8W30L1sqb01+mEYfZ0FTOFjIZfzX7rz3xLisOBTm7UgyrW/TTg14u9AjdCE/Ht4FVL
6BJ1H3IYO+mziSR6+iTaucKQO+2Z++R89LOpQAigbtGLT/8zBE9OfNTdgI4QY/nFRodxa/CCsmjs
60uxZNhhKmN4Ts+oJR0HzIQ8aAGN19rn+vnDAYBUORoIxDAwklJIAEZmkkms8kHGbFMYvuh29Aos
WMCP1VmETJL7RWp9ul4WNNIIFAuEewsUqmNCTEt+YX8zuAOzjfQyMWYf3Ze2Xo2E3+V0GDdAfa3B
mLu4rOGI/BwdRNXh0OQLZEiu9gavHNylHupsJsh040AiZZB91j1WCe13clPKhaQf9HXLA8Dzhayb
+D5DTz730ccoqoG1LeGWNnQIhfYgmcmpZ8sydb3To09bqPI4vVoWKQ8VNDjkXux/OAztP2TMbXvb
B5i35Twp5H1ICKtsqcTu/86xXMif+NngsAEwT2uppHP+sA+e+KP3qW/8sJ+AyJ0ngbSgBwBiaW9w
1H8FXDy93J+Ds5u2R2a07ajaoy9YhN9hMHToGzUv0pVgXq6D4PxgbE+MY6zui2TYEIXDFrV/fSog
I20Tyr8ecEuGIz8FyyM+wUsaqzztXHUplzR/uDcXbvATnCJGTKnJPG9kH3gdJkjq/Qjka3YfuZTW
WN3tTDcSlibK9K7UXI8NNutjD7DL8SusSwIexidvuLRkxbf5xdXPU5b/QfnwELO1b20TzyRs+8lP
tFHaE+8tdcDYE+Ui4kmtdKBbKvu4I77EfTtPrMD03/Dj4cNJmf5/WQGGHXcO6HOWOfMBCqwNzPdc
jFHnnsGhFNtYhSF5LrceM37fCs12egTCpDD0x7sD0oaT7MIuRS5RsSr61mJbwrQR2DOxN6pupSUN
dKSW55HPfpxOSxuvU5IAKi58FM+Ov82Vq4O6FGd0qeRTiCWtj+319uPYkrKQUvkd1USMEf84+pqG
GP/vC+xn5IOt/buiIECrdU5lnmGk2yBKyexCJtcDZ6xotN+l+SOW/rT0xzz4nPciV7xkB4OH81Dz
DX2Lvns2XUw78CdJ5VeDtw/aYjaK9zStK7+ywckzPQ0eBjYwx+V9qqmdeu7Czj+GNxgGLuqFXEkX
A/NG9nl2e/2uOaIrnqBhglX0fm4I9DkWqbzHKhXN9Nnx+NGBmnqgV1h6ddl01VPyTAfCRBymcAmV
Er449N8Fegt24GIqcu4f5+a1tDiQM4NhkmjYd1frgKn5EB/rilpBAEy1yFMMpjNLt6sSS1rWZWdN
j0GRZIPM9HEo2y5Jifv+cobXd4d/CJJgMiEA9Aj8YnlCveDmAjoLM8GOkdSYFubnymFzPQWvDPo6
ANzaC5D9L5/erk5JLLJlGkJ/rbKOSgwLMUDebRmgZOqXJN8UG0XPu2ndahVQ2Faem/tm9wxYp9Ar
jxB1n+aWpEXb3aR3Xh0SvmhibLVd4zg6kBPT3YLQKjpqWLdrpSfJ437dAZWGnZn65xnwH7tRIhkV
sDJLQm+wgCtPKsgWZSua9d3YI/Ue4TS4Keo+XyM+SZghQmclda6b9CVfazJtopWxNAzm+QXAfThd
wnVZcAg7wT71Qi/pv011kQPvplXqkh+G3lkTK1VmMe7oDr3Skd9nQUkOnB3i5QJKBMT/souoplr0
jvZIyd+6ZBtGZoFCxW0ybyL7ikZYyvwm+2ydjzGepKh9sCxpsZB0nMN5WBhoF3FZVRiF5u/a4MtZ
mSOorS4kdXq79wRzfC2vIXYkzSjKgSVmt8bcrHg3+2hVncDqBjgMeXILYYuwYySs9IcN/3+YbfQ7
RoyY6/OxHcoLm5d/6Ka97je+OZ4DHG5gQ6VCVKClOYBj6uSeoODU9ivSbYMwE2m9hDMk3UWXKZRX
jHxmFTtOncEuB01OR/Qa+5nbqyHdNDTM7qt5KvpJlZBP/ga3o/S3xxmce2iwHI2UwUjNfKONVZta
bUS85UVlzxh0j6dk1xF+are+2soJlx2nO9S16Hf+K2zvFuigxWlUP2vVM1FzIjCIc4eBC7WAvQZU
PJ9jSqFctfeFyIU80g38DYdkOWM4H6Ntei35HdUn4G3AWck237vFUR1ABxVJ5JlnEyxxlSmOtRXk
aDvnJQYvNMOXleYR/eYYrtrCjAHmY2ArSEVtZo3uIdj+IMdsxUY5KB93EHkReMMEsmOHT06w4C75
ybjXk9zDFkMP40Sp7at486Vga321KL0pz4rczgpRIMBwAESG+ohLIL2GNizhUqonxkJ6A9Fk7Vlt
lHAMMT6Rft+PCmi6zXRqbKIks8/PzoHWm/nF5AOgW8i/B6X1U2V+XZKAfy4sojaHBt33hxcuKCVv
8WhQVZtmuU4mZ6az68u004mOSjfTpKiwN3VSYcpQMSu+w3J4Fm0Sg1+TAxl4CBKUArQqtaRCRPJ5
zfsk0tm+oKr/92LdTrwoB1bjXrwGUSbT1z8MKvhBDsm5359eZGg0zddKDbCmakMivRqU3jC+wLVA
X+zUe8Xmp/b8GwvEfNDl0IFvo0v1A2aT02CXxoIXo3QAU03RaCA0a1jl2nvDhO7WjjGe/jiHzPds
Vtihil/PRkXZD9ihGpCjPGb11w0s+Sf/6yB723l9XcwHiaG9eWQPU6Dns5kIIfiNZfGulCOBSd2e
r1oNN+mxf+AsTYk8MCWEGXceDvSNuHLjSz0Hmv7aOEUFD1tGYz2lJ29g/f7i9h5NtY0by2N6STXS
yeNXA5pJp0ZoK0qU1OjZ9MsI/fBUjRG5aGOOxW9a11bkvbbkTWY1veuZbRbY6R07oOml1lAjYzgk
62uOErvguKJrhAi6cdWvbo7hrIlD+9X3R6R9c1kxdFTtrbqX4jdx7dNaCWTRQYL1lDbTNQbt++Na
SKdPJW4ziONVuSZrZQ2KyF/3OWBGSCUaptyrTtxG00Sk5xXpY5w+ehKTAkHSkwnSC/4AHp19Wvvy
yaqmp2qmHKk0tQ8dMWf6JDuxHd2Aym2ebGDvRfhm0UaX7QWlYHTDcAp8tHWC8IeLKicS9hwHh2FW
YzxPU245fSREGaVhj59BtWkRQYU96Rk23RMBOvEKuniWx8StlWTO951sPsR4MEpwBioxphrt/ed8
CT/joP03zOhJDYk0sNlyWfeJ57pyCJl0blfCR+bU9imRJHeJl57BO+oSxSRpRoZN9oiIW2SGFue+
btvYprMagtzexweKfS6ewi9BJJEvL6cmrmebbbeyvkcU/DUx2MFj9HIfLbAT2VNT20R/xXYeDbdc
nr7YJDwVlwhI7whtEC6yJJAoP6/gzDiZd8GCl3cJQSPTU1GsmGtL95HaTMBnlDIGVQhNCzFnDHQm
mNpvUg4YRcf2h6Fksf3/hFlIqKmIgtnSq7weNxMFTHll5fjXlmmckoyfVSUmsjFpKL+Bz/T15AvK
rAp14klEWd9oyWOubwPLm/qbAVjIrWdgeyOuP38xA2fh2eYDUZ6tqr1k9Sj20GJex/sM+v6uMXuH
Q7UB0wRvF2QyEeQEwMwDy1qh/f8VKCARWy2mWBE2TM7MfltEOdk5O8k6XWBmxZDUOUt+TNttxS4d
mlg1zd1QCeers24g5QvoNdZFRf8w7WkbjQBZytmmhFeCHSdipBWiI+NHSbeWXZNLxS5cvN3LLsaE
Gba41jJ55JsXp4hZgmws/D+MXS6AkLCMREaKDkZnCFXb7ubrb8lJK+Tuxjr3R9L9o+UEq0zFUI0B
1iejFAz2kQFLpIX7KRxUyZ2KW3TZnJ+vLIEEFu30I0gxfcC01WRY6wcjq4vMSjrbiBtWwaGpGEUG
/Df69BDN+4elNWyCtedZHgQUW5l6x5QsX9Ary8PsVWv0nK2dnL96fqpCqBVJ/Huu/GaLTB/Jja+A
z59aG66/vyTjZ7InA4nJoBZtibGliTAw5e8TOIB0F/PvKHB/fK51qBcUaMZyHzkOrbkbKqGAeUJ2
Bq2y7rtGW7AceoAzIO0yQk5IZXTKlv675Tcmti2Wl3lH2jbipQPVrHQqotxd0TNd5JwWmtuxzyNN
SdpxvpruzG5nehYEzr+f6Jj7SpPZ9ljiIwJR5CBNroZhHUxdc/ik7Cl5mYUNmmeH/cUZ5xrS2xAg
wc65WkJRm5ISoHHbTWT+joisbOfDGOxPrl0iy5bfy1Gw1ozsYWvyptt/kay77LxLe6YJs92MEu81
oQ+vWYGdnXJ3zM7lW5LJ69ziWOSp77+Ezj2asOfxLS9jt7n8LoY4m868MpV0V1Mvoxwddc1B1/7P
1xStwhwYOl5xJpebMIi3+z0PASf31waY/AeRIbpED31gf/QI6mSapEfByBMQdBT1BIpvFnLyhs5w
y68wrfK8ts7Da5TKnhZxaTNe6j//3fjI8/8lUuQMqINmqeYPR9GY1Uf1r6wIDWPisAO1ROW3MyO+
Q/PwwbK378DXPcvZ29PIezc+etQIZjFgKL3vt0+zcVB+o4x28ihANTHqHs7yeZ5Nn6gg2WkSsbFV
kR8Ibkiny1ZQYVLmz3KmDftqJz3xCpbKL0+LYX9/bl0ild/AVg7udbhxqsDsmisQM+GsqNu6qNSZ
7Kq3q6scHAcfv3PSIFvvGmrwZUdI1Or8EiEM1GZNo/X5YRZCcWRqO9K3Dxzu+2svECiA7d3tMbdg
xGlB+WWZid8+Fi9PW+xMy3wq2g3A5l/941FF5q5lkx6KMoAMUYYW2suwN0VIf62OciwfsSZ7RcJ/
j1foEWPqvj4OblGHCb5VLxgWDoogM8+c/5ushk3KmJfZnJ56cLSFQeKi4I39Xx1mK04d3fOT4Oeq
DCUJ7ORBwORd+ntvKzCYBvcqyO9txHg+PoyxIHGOoxpASU9pzftFII2iDX3jW1nQo+fzE9yffJ60
gFp60xhD8vDMgmFfho/hhPCRLz1owGrBRtuh8354pwlceL25pA2wPIpy3pIxs7jxFh1VvDYN0lEN
Q1bGp0NvLp/k1/u8jBAZf9X6GNIQl4HYG73udyL//uIUlETqk99lD0dJ062cyh9J05CwY0NdGS8C
ust5czR56T4E4gcaSJY3w5fxqKrzTEALZhFI+yg1r+qPWVaUJXZS//PNPWDvSoUoM8wd4t5nSXNd
ZzrFzBI0Ag/384AjmJEqSxvcxhZApBEE/XcDtnVXBGoO85onjBr6ZxRwewtk4NbccnSqR29q1wFE
9Ejy86K/+gBgjVStT/K5Zh3n4C1mr1GqNiGgeGybBtyUYt71fFv7MHr+PnaTBCPLvdbkj9Wm0/mj
elxvujqW7IvvlvJ2ZWrBpWxTzHnrzU4D0rq6uXhci+Y/tpk+ZH+pQOWCjpXKgFD47k+QR0eqECEx
K7mAA/NjPRw2ec6b64WAq480ye1KtNczx/yPUl//Bj/3SvRUItpsku/Yl0qWM2a6oMEy17PTdumw
HOAT4ZT74giFSe6UoL0X3BbF2tDj+jqR12M30i5qfTQlRCisv/n7H49V8+xPcUSxPRGcIi9rqY5u
ApoGqBL+8aBIVHGvCTwNOVCbheAeuT+XWIzAtwS+ZcPe+VHkFVbx+7f3l67RXClHSlOI/4I5RNdk
Qjhps6/t7ZgZCEKQWc1lgcmgdeZSKpEGdOtfTrzocWzXJRmpulRWEU+SAuTksQOg1Pmx2YX2DndK
hSVBcdmA+c3EHfICFlzFQm3qFGSxiDNv05G3WScduEHLEhy+4EXx4G6qCWrMh5YvL9tXcEf1vpGo
GlNnRyhY6DzYpkg9Ha9x3bxVxdQbfxi+8AyVdnHs32ZSiN18dnATlmwk1KDyP/rlUfxAsKHGLOVY
NqFL0u9xdJ3Wh/8v2yEKAkJ5fPabeXSmcSquOkfDB6joTOj4VVNBxtpj24WGKdfYjSU1i/NfdgHG
ASBnPvxgu927HE3Q7xlw3/TTky7GNYPLtn/QhFK8KBhFk/QnVp+xkixaYli6kvCn+O4wEA8zdtKH
Qn4Hvvb2o1UYRLBYlR55hGZEPUNq7t6S2Nk1PyQfVj8MdQjQ6Fhyhjds+/uNHxVwZumMuIIexxfd
oAJ+uJBTudMb7BcyK8c1b9/Ni6ErTIkwtds9uCK8C9yisH5Soo6UiIP3+yu2Zq3SHl5tq2uGc6eR
m+sOpzxgD1+mz7tk+JOgFN/MQXRiFFu1mJPBdThHJXBTZ55zuZT/lGaDr66Vt2BfI39DJfqTnD8m
gB2t7ykI+Di9O7Z0EfjZkVrKriU+0Vc2LJo8xNOA3hxWXu8fFXHG9tfoAainRbfjSRAPqJ+bIt8z
uFlShoqQ01SMT2qyJUEb89OMThmg8OYYHCCXDmQW4I9+uyI9Gn+vOwjeMJ6oKxM66+VGyMLxUY73
Y2Q6znrU0JU9K4aFiZg46DkPJw4/TBZoHpIuXCkOJ+WscVPwxxdOd8LguSJIHbjAgv2AAAAPAMOa
MVzka2IJvCvgZHwzEoz+SwIGONaTEyNFj3bxiw3poHU7bXZoAgd9AC2WwNfV6wE1QU/zUnmRBfCL
g+0XhJ93vby4ClQ14W0uoDAEDfOEqDlUfOc78tEEX6AgxlC8GldSqPILkbVfWb629zZjOhQvTSUX
PA6AbgjgBDLdvy0ei1WAVoeDjY1SLCGO0VjXCbpGg84wEpZx7AxxzWv/32A7saD111VGylw6Iejr
q+GXz3JJIwWmF4jDPzQzbgxEZaPiEiF/5BLzWtzR1G8W0XobsChsXtsE5mqqU3T7hcNbH0YSCup1
cWiRNMygV3wBI98svfX+XqYlQpfS+5Hb1R5SCSqsZnk7zngYBmKg9fee+d4rTqOv/5LLDaROoG7R
NfKSIXaHAx22wkOEmOAgS/4RCHUEeyYOInpqddX//wR6Wt6Lit70aXLHEOG62q+JrbPdABCcvLBK
/jzKZeCy+1YxBUq0gFKVaGUo07rYdIyUWBdmTh+H9ruUE35N9vblvaEGm/qAoaVkdSY/fi59qMAC
E4v8cQp4oPoW0hiZzaEv9thwdbyVCEftezeHZ0pO7asuHSP7iuwZCaC4WRPCrS++prM81OFgMfBQ
MeWIrDxS6w+SJrxkgvyJsIp/haDc4dmNtJsoBbP8c1h5uVlyGz/P6DsJEA/0w6XrjWOBrLHCSoXX
A1fRnU4eJe6/IRGqWQUdPOL+451M6PoJYdgaCYF+PUuFbubgV20aGbL8zyePfR/Hd+slppnzzrSB
EHYUSTy0nEVYTWcFJYydmKiXtObME8/2IunKE1kJ02EO1230AbWk6sHDm3/48edVmbTDhEkjuiop
pGbZzeXuc+0ChMnOjCpwXjRi4ET1n9L01hx21gpBREbDDC/1oMRcTLbWhjABYnxqxqK9vDcSvEAa
aXEUGtzWep13cA2xaPIRue+cawPtkOciEL8Bl1kFbxqUR0wMVgCh+ruT2Ok771wkfhuyS173ya8M
DEWsFp30/ElhJQ4MqHPMc686vznPlOsk2v9WdPSfHL54Ep9sKDziCm3QyXaQ3zAz8VQWN5+YVGMs
8hNfdb8gtgHp3MtWoTK/Yjn8ROX0PtiT441uuZXFzozyL4bWbfVGETpjyDzoMMcQdUF5CgI58d1s
qp/o+pGwUJZ0oTMUh9G6CMaCjhW/d3PzI970AYFW0Kc2EMv30vCO80GNEShShxNEQlGMBMmYgplS
afljZauzeosXw0OjRlzO1Dw8J9kemXUbA5NJag64DGYzAADuKBA3sZrAQzMc3q2VWg9+zoWXSJs0
qhhiQklsF0vXCfCMr2i60RUlyZOF9G0nmOddUO0QtYFLD7WKGvWTjkxXOhZOB6x2u+TJ1u2bDBrU
2cvEghKCaPYeq+tP+LtEFi4T5BQulvdeDZ9Cm5qVAQHIN84J3OSCUu+tYpjVZEY8KTFKzINTu2Vr
VbY8DMI7OW+tLVueYhtgnmwK//OD0mzIUtXGatnw11kVxVrhK7g2+7ibDSCWcvXsHRdFb4Ohh70S
RBEVWLAYim2expRA/J5vr/j6MJfCZc+Gug1c8dxDLzHYi9LHhUjHwU6IlnOsFXAIdifXmF/a/N7G
D3GtrXsYig1KdTkh08SFWiPRGPyhraGAUGoQJVkmQqOzbycxVvTkdAIWUuFgjGEbEMs+vDChOiN+
6F82YNdOaI6iJEP1nN9ZRky0AxsiUyOQwDt6hQxVQhWm8mULlq8WsVS8gsVDvP0Mvz1V+nRxgrie
H1sCVixpyPvCNP/y/uDy20VkmH5iRQU1h26mUYTxZZR+AAXA+zgm4p1WKMrb+nZK7xPGAv3GRI6R
lpv3mM02dRM8qDcZV79UJzbYqdQKgfRGeQeZj3pLCJOFXdYMRXPbNpAWouqqX9inhpGJQT8Y8gXY
b78ztC3n+i9f9QQgN3jc0zRuIKMgbFwKkT4EbAronAe/EzdD5/3pLAkJsaN1b9RzT4uu7QLmHVtM
KnZdFwV5pztUKtMs+rsrb20Yehp3vYxEoYeeLpPYeP3T4qvm24E7VZwIY4Gv9rciLm/mftjetKil
EiwaXwerNJjWOQM7eW/5EF/pZostCzjqISIs08Q/nr6obSeHSa1Zar/YCE5tURqYXMXnE7qxd7Zn
GOfGdrS1J61ZSWBB2HoHfak0rZiofcNH4Q3G8XEsRvwMPanTDcwknhaTjoJIjOYIe7bdie5pW7XS
+UxpwukaQP+80m65r/PiZ/q6zgbDrTlX3v73ZQ/PlDAZ6mJJqpvZn9SKHi9+eFWYidZEnrSsT//6
6p74d0UnT9WdG6B568xruMN5PyiTYM1eeACfaQHp/LERg5MamA/QjaLdELKJ/Ox14GpWVQlKn0QO
dEcb/R02tzxjEjYlHvtIVX7oUOfNGX6HAJ9wtCN89eOrh9XY48GWWkMdhfy5U8dUU+yalIHupcfw
SEuRrLPR/zRHHcsbg1RkviRSTEdqoMwLizaS3eMWpl8/YWZSk/8k+eTtyPhmOgWzYysaqAJGOeu+
+ic/G6YlE2lheBIBvTtGlFkMNZmEAC8IXpNf7tRYqKrwXnOBM+mSYF6ErSvWHPKqELPfbAQ0/368
lBc1jObdmETcphrKWp5Z1midzpwemiPfLyWI1CBG9MlODVaN8BMmhTiNgtgLzBK01uOzfGpMcBxZ
EwEE4CfRDvu+AWQlNttJ8jfXlLqDWvfCUYazGU5L7NMsZCEFRz+S8f5iG9gBRrjVBWeS/8gzW5Rr
Cr4rjxVv0xk/2AIss/6sZITuJ4+N47TYzR6v/4rFOqdXBHkO9mpbEfCLfz40qbPWssk1cw4qzPWg
1rATkZoI4oYxOTRStWMz3E/KFKYVViD5YqDLz5mqissURmy3qon83jOk/Y7/V3PiT++uOxduqWzv
vuL/0yvfTYRKk4KKVBl+WuIUSKPiY15OFitGwx/bTxFLngUlh1es1bCS/w66Enj/U4+g+O8XgJ1l
Dzc5Cd6F0sbHBTR5c75TCzmvRgsNz4zPfLVknZDjIlQutvrhjAet1bMA5t7z1J0sXgnhX8V5jAY3
YY1vLRPhsSc90ww14Q9FDTQgssP8L+fL3QnLcE7YCDDVWgCv2HmgAAUNfJTbHnc10kx7xA3TYJn3
G48Abs5kvwSXnWmCvfY0+Y3qqTHk8BT6O06+GsYTGsFsyfZ2q61dyZIrxyFhlHuvCJt4pfOgb7XM
/k/Cw7Ak7HN+Pc7mfCyOI380Q+ZqllWdf8bUEAo+X224fkf+aOz8O9dLwm8281klVNoO6QDlVzS3
pwKr9o/5q7xCP4/2C+RTQq4aIzG6tzzW9HBdOZRA1o1AolCHFcncWGG+rNuqV3O8GoAD2RDhKwRa
mBzcwHjFYOQvixhgDFqFJ5m9kCRmkHgZ4rlYZuINrA6j2GqrFzlrPEOL81+/iHk/30xEFNwSA8ff
YBl2AR0+cxEO6P6I1nk9zTTSO9oSe2yZ9DhzhFEtMDFaMWB5SLLM0Fya1MgjCyYV5fhKLmpz5Ayb
0uiKRaqdOzKr5j8yWaIw+khBx8FeTobsrUYuunxDsbAU5Y4WZNUkqfzMjxoRr2xM4jf461YUcD87
tQx2AqpbZl1r5SkmLmANNHdbnn9t6FW6zgcrciKe3ITs2uep85VmOVwtTen00+LZS7bQwPmGhASu
eU14JxGKEIlaOawgl1PGrbYFRhzsHkRWv+MSGFODSVKSrPMfbSXuO+38KSqryr5gWl5tKuvN8LW5
bSOkJCzNSTBZQTjN/82PA1oP3dFEtAGr+jnfSyncnilQumzNmL6j2s8iIQB20upbzWxqb36KJGMN
BOVE43qtzUlKbJwqQ6ZNNqHBmYZ+cSYjoHUjw+1mEu4+8tdEJmgsPz0vJSgEntuFjGnRKowTOoSG
zUww0fvhy/FnhKmnBux2Aig+sjawnX/++iGhej8hPFnkipgN9qLHRFKrUOUYIr7Fy59vFKJ/6LYo
OtziAamUe+pPpbuRNYZTQo9BqcIZRKmk1x0MzbsNhs362ADvFUUjF6IWcI8O9KnPt8dIjax19Aw2
yDNURhGaDdv1FgNrTTPTLfqkNWFBL9Ya7/IymiTn1HcwVt9gjsmnX6Pdmw4Um+WwtnEWjoARuhLT
6aRbYVqy2PMpYsukbnQD50xL4xo+LyKq3QSyBx5l9ior4j9KHE1TWOOvf8w9hITY2Q3EgGl5yGtz
eULXu0wkptkCbkLEvufc9+pFfTikRbalk6dKr2hf/ga4vKOFidrLbMams8UyYSElndlRc0e0+KKc
X7YZDMej540nftL0z226Rl3sFG9JgCq6YSil7kVWnvXCcSYGsUpT+tlac0vuqdOHUnCNKrc8gDwq
fDlA5MPtrA+A01OEwTKRGBaruZNCfMNZwZ6qenyzmn3SlTi2EQG23XWdchOdfRBx1T8ksI/wMmDW
XbB75s+xhcHdBacLj1Ssrk+Q3Bc3KcIfEjFdMO9dUzbK+PlsxafRu3MCgJTa1dfT3QQXp/zSBWxA
QUavH2FJkqAV+4/YmxUC1pLVYSwNOVAW36V69XNNbj+W14vV26Fx5eS7V2LiiLCg4cgQlLaxVRrl
mC8WjQ7OuvxXTl5Ehf+NJda/Ewo0UzhjBu1CTnr1EUAJJ9ViSTe5UHLpc1AV2dNuk8tgoeDc3/BS
VLS86agPKWTdPXOiwP48/13GpR+L5+IhsxKm6PUmbUISK+7NFkVh6ruTLQxvEpa9XjEe2JHWF4cP
/pvDBegoRJZ94tP815WKEqVvvNlqZS94ky6eT/22zoCzqTpN+5jjhYURBgC6auFSWyIg+z//Lxxk
1NB8wxRRC0Od6L7XF0hYvkJ5iBZ45zTZtcFOa6d1uLB1g5trMuYSLChaTen8bP0OKGqvi0a2zSlj
cQ1sjPmHDC/bWktFNM+6NebIiG+t+Mk0lGUOCRuQjg5dK5H0vcFl6yJPSiPJhHvWcQyUMYwEFREw
FIJ58Q6sqAzyzngOvENs1fuVz0Ojx+0a5JQY/tiZZCo3ERaUa8tEH5aDrsigWGveTCocvC+46ou0
8nNCjwVu+XiCQ5N0V192ign9u5mcQp+Rte/fNMFEqzBSK1I0O5AnUshLtrbhN4HmLX7sj5+F2aqM
Iqs7BTX/8wV3OdJna8e9O9lfzS3jyO7vBxzgGRMOOCI00oPIqFJlYlMVyYOlZ5T0HjNGJ9SXBiLg
dEOYxyc0Zjyojg+TV7C12T5ZCuWrgLDoBO61GM90tKwX0yfIsjcOGdmF4DEi5s5QjG7QDIwp7G5m
V1zOUBprF/42N8gRIZtvCCQbZbFQWu2EFT5A1Ep6Q0UyJG7602/LUb7BzNth1W8ULy9zByRK7kxX
82YNFCE+KDk6Xq9q+JixX6V3Uu+sg5Lwf56oR2M2MSqI+pao4VC0jnyfzt3c/g6nUcaE0F1rc56d
LaKRfQR1/1ANqdGLyBMZ32e0HDqHmnOpxp497anxsSl3JgDvbk/cGwYPmvASj4ZhxtEu94DVfADK
5vDQJDFUjl4n5a2LBVTJAnYgQEqYPP7MQmE3OC12yegoUjBMhHFdLBdiNvxq1tFIjo+BGdjyO0ac
mbzuGWcpLSkfZUtWs5DqXffcHa0a0VAepCQio99GE5HPXO+YIMSpmZi73W+MxZQ2THI4qcJM4HJ+
vGERL7e6qzZspSOXuKI+TL3i1MTM3qtiPd/Kvdq0tmFsJK59fC22dbWcRnYltXSyQcNWRaK2V3TV
xhEjffHrMx6a39SM5Enzu8LDAxCBAaG3djvJz7ARLLYfIqkOLceeC0gsBEAomVXgpYJ86awFqf7U
mNltJW6HvO7KFrHnF3cmSFRD4GrxSElEWM1hkISGBCHnvEj/Q1/7jCO6tkLxr3Y5lehRWot+N69G
ayyBBSqBHwI/xAodhbVw61d/aVqrVZ9y/wpnJRni6nqCHTcssIx8TzwdQQkz0WO67Q9mij0TOJ2v
BsYJ7GEMMF22h3TqMLY2IVUIfS15wjUm7dxMuzbF/fGCK2dfsxPGTBmMKoIG5odIsT//SnzyIUqr
filaUGEn7GZ5GXyJxAkTH6cfGL2JbyOS/Yf4o20kC+s5pOlfQzMBPtytWksfKwoNFuueWe8gl1Gy
nio47U8XfPmGF5bA98kL5c+ReM+xnH8sxIUdO5Y7JgnvuMCunh3Sb3tcyRZOKazQIRDTemwMdh+M
ttTllVduuid0vAybbdXr6VnFAp0k2mtiA4VUoV9UeKPxl6CISru1HfRnr+XBC4lBQsRF6mT2zTFB
0lyCUapjvFn5OGlzNU+mG2ws5/4OTyi9IJFOfyJh93lkXzY7xf4RrwzmgQxIDG53/+fW8yZdnQX+
fauVdNiUcfNQkFG9saXnbTmmZsg/aL8eOMa+9xK1dpxIq3YWozRuN/ty+9D34W9OXPWr+P4iriAy
VZjwYgD5LJIwfgffX8h6Ry5VXTRfZZiY1K0LHTp2t5LRRJte43t0Fh3LM1C4SscHaVda5y8TQAHr
OkxwPdi1SdH0I33Xdd4amNNE5sjGisDvYO+XuN3pAo3xosOzrnn7OeVy5k08iVh4GZD5larpyMku
vGGXnONPZNfPo/QiP5L6A9w1Lw8x3GcQw6ojLiUOmOBrzOGqrP1jWomsi7QkX0iu8r8b9z18YwO5
k2bOf23VFYCNTiJHaARgZ8XGL/6UaWikuAKAnJxEATjnUCPEDd9Ioiyad9vStBsO4sEVA+m1hPye
itV26iUORn8LhEf9FIIS5vAMzsuSZgRGALRTvk0p0MPQPJMfDx8Vn9xxIbji92oMXrvaQf0PPcnd
mGTCae+uaGfh0AkTuAcaLjaZKaCkBHYPDqASfcG8oqpg31Fk/k2HcdrRQPsZS/t7wtcR6DjOyD0c
9Ae7JNuFkFNXVe/DxM4mBv+wdtD/7WFacAvifBdelqWfkGWpujjbxv4FWPii2jOh4dITJg63dVW6
xcCsSOl70zQlSsesSlhoErIeWZ2ZUUxGDiBLmGRjKkPttiIf/CIjtIg+ny9dJnQrO0QuUSXTSufm
Bq+ls/6+L5ZNKutJLvEzy2kQYek+Tff5Q4mqATbBtvjMtjLqPJ4L55sIjQBDTt0COWwYhdGGnG2t
kcSGNz+55Lxdl2yGVXyPTrkiLKvfXHPRuAkmhEIz88c7+oXxnQvTP+bcHnOWm4QG5yDJiqpyZ3Ql
n7XPmQya7vK9rIRZzYqBRLgC9JMOX1pTWvtVFmlsgs9HuMtF+BkBHpXvuQ4qoptyST4a5yu8SELt
I8ofmVRil+bYY4C6fa0BZinWNQjzoPxFFh21iTXDKs1OlJLO+8bz6ct2FkMSX8V+BIH8I0SLuhI8
GJ/wu7YPo51VfuKH4I+xsPUo0YkP4pCjyn6hSaRDOLpMEHQhnwdW6MtrEkbDzl1YmfnZNsIZL2Vj
iVPAYTHBVxDxjf5v8NuthKOzumRbyssAMzvHQKmQj7KQdefswv5Y78UC/b85ZCHI9VU0Bqxv1pkx
WNdPdRYH2Ta+MUvivWaE1o92sIhYesKbWEVXgM8FMAndRXz7Dz28GncGGrPZ+7IroIDsYynJjRSw
Ycz9rfaKTiV1/5+Pz/AVjRZ47s6SclKSGQD2wKH5MOkwBkEKPfUN16ncfAsFBN3so4UfXHR/t+DD
2QgdMHpqvhJsORLJgjBRbHiFfdL5EL31ZzPejN5VjUbisdQTDN1jytyYaHc3KOvdl45P4Px0L8kc
3QBNctnCNhfwnROsms26sbOU1jhDOXIt0OZgLkd+FV0UAP/V0nHO6mLR4uLowwP6ZDETUrrEMOVT
xhxgkp/iqreLYGHCculPJzy3A9FW2GDgI0q4TBB9OXjQrtJY9oY8UmfTlgVEYkY8C+0uNbss23dg
gEXzokfve5ISUeR7R5nFm6ltzfgv9Z6wUiRTIFXo/9pFot0HuTgirqXVR4hX2TXeL+2cX1OT3mYj
CfT5iGHwqie8r1TnZJ1ONLrhfnvsLIJuqmjWjulrUZ9nZadTcs7xQIeyo08nYhhICqnqz8+nymuu
n5JCq1l2SDVrLrnDGZtNzmEZulGV2pT/0cc8PgQtZJyEraMqT4ZgGpvUD4ituOqY06EaHh+cJPbL
l6lriIAcAxOvkN6toU72fl16r7rprAJq4SQe1F63a7KKjwEQ9Dj97yHBXXzYT869BQBJN9fpTSec
knxzYd294g8DLn2E+6bT9EG2sAddWBgPWZtMfbeZQXfxn68M/0KxmGcCBFJWdsg5LezIkGK8MY29
KRRe0QcEdvI2/+Gj4VE89wzt4XoghInOA5R5MNtzU38Uz2kebSiiwO4fE9VbwdbYCTHNmc+2jQDt
RqlZ6ofrtUwTkAXnQVPoQEVQqtkjFWaJmzX9ZeV+Zsq7T4T1TiZEBOQRzFjxUxa+yyITStXKby9a
9ltgOwCfr5auo7rFR8A4PNQ4cjSLPCiyQwiplDqs9bVJ61KwULwEDqdhbho8JopoAtTZ/2ADE242
gbIVFtyTdf3RDf/UXcsiAQgKZZOEWGcKZIxFl82yiNIahQdLZgHJyUm+tqiBQKvEV+77bWZBG0CA
D80X6TKhltYGbBpHBZ8HBsQPpc4rlOHGTg8r66d3E+hMt/EkJVOMG0BzVqV1ETry9/7zFi021BUl
C+WICfr4VlByfFQqlAAO1xj2SocTd43WnhkxephtBAEpg34Ly3DRhoP8lKOhzqqDF9VIlzX3mkRj
iq68pF5BeBmKZUapkuW1sCoBFXk3b7EYqvp4yrhdooNNqACn2UOsGJUMI60Wi+YD78aw3UK9w9by
7ssTGZ5sa0x/QqW/Zex+sTqrQCtGabwUvpVh4rXfeQTgXb2mQcACBIsZ2BPoQOiQPRfR28wusP03
wYdRANLjhBt9QDfgedNVVBFhw4VsxYrQMqSLkKkJ+vscbX/UlIiH9hE8c+d5rapIfnRg54l8vYvb
imTzGO1Z3OYb5y1L+F5u0xlpY73AH0auVOU/aHjr3WPXZT7hyR0VC7H5lI1Ex+Dyl2hfFx9IYtON
n1W0ScYo1URoYQNrMoa3FOCMBUVWOoJ99KCFsNnhnM39jnYI7K5SyN9bfOo4FHeOYTkFPRreduwO
IBLkNftU5bRZsGmaMVpIRfyqDW8rfkam/JImZpjgKOwM1kSvXbx3ti+ioi9FDrZ8ePdtxzZu/tx4
Aif2lQ2HAoyidAy1geVyUK/TmBwxiruYg2Czq9Awvhc8uSwpeQpCPCEWMM07lEBl1pxkUqK2KhVC
oEyZaK6yLzccTGAxjG3TbVaj06LYr/7m2RyfhMJgpGGcP5UVQUAFLJiuRpUBmwFuWSSYSVgMJDMv
FXZMFVIEI1kE8WPENwcH4xDBjXWyR90ZljVMsTdCp3eYQm/HJ0+bgMkNVuNid0MzY6DeAFvqVnv3
3O6kUeq0eAQRnUSG/Jw34tw2QWmQMvPuf3oZgHR+hQd7YNh4e8ZWns05LwnVP4WO1nGYNXEu4pIw
ztG6dsEHYwoMrgz8ffeZ5Jwcw+lBsTtLzXTIj+nHHDJyhoVILtAdIbB51LVWf4jupKdF8ZNXlEAS
rKfvZWU+5Bm8b4FHNEcZKsY5/qQCtR6Fw/Q/YAxwN73pXIVxpqJ3QRaJB2GBYmqFGhaz8rhYIWTQ
cLAdfiH1OJXGz8pB1lj7eqNb0qGafWBxjLVi8TnYtrskG7Vh5cUUe8WBAtoObtFCNs2iQ9qPNDRK
aw5XHEiQRVVoj4fRtFZ7CmHS+DtrQkB4GQY2iFXu3jNWPmXBrfmEnnj6MNujK+0mKigcRRiera2z
/WyNz1XPwZWMV95HNzNqNqEilyICLUAQJjwthQScXA9jB9jFv5vw5eoAmi/snx2y6T6VDorXFmpj
cGSTSs+6nxtggQA0xlVNRT9rRDqgj/PHZmC4IGjJ4AlLGvw7C+GwZrPSjWhNDO0EPg71Fanj7p6o
VaPpy0DByi2jnftRyG+3aBOfmXLlMgjxGle+DfBt8Z+ZVheDjnZoSx97jKbPd8/izrVefanjW+jC
TVxrprq6adRh7JykEkIWm0w4h6RQCkdj50ZkFZb1RE4hL2zxYH590F+rn2zyYfgkW4GkRze9JR07
AVD25mMQyt517dEz73bIKHVoYqK7fgZrDB7sQ/TCaoLb1KDtWjviTkFtRXLDwYjAHKLPoYQxqwR0
+atgIC6i92rSIwkPkeuGu2r1/PHxLM86wk1kzCzdEqxA0x+h8+0HtyHG5JhVCHxY9F+Efp3YNwvt
1H/NaUOVszBqXdaE/muslBCA1M4S8Z0Brow4y7mXjiUL9dOLldujx4CFA1plyqkkO8bXAvasF9gO
AxhYZtPvU08Pl+O7GivbOIY0WvxT7I18MtXR6hlI8njOnDb6lebDz2FZbwo2fkjV/CrwpTk1DaMq
ciS6RRZRuWj29cpJqKIpKglNbjvdTWakqnu13YCuLuWyDXEhmRnnFU6nux0cly1g5kRqyEHQiZKD
nIievScEsfuFiaT/FrCLrfqlMUQZOXRRodNGhz58K85crRRZ555/hkseiVFJo+8ar4d43Vp9WMbI
hx2A5RoR4RS+AKt22k1Wzk8pPsvcluGbZOjFheQz9YBgYFFCMQRxpcbQ4euiuU4EotJQwRQa9wFD
e8aPgIbXvrf17oX7k1Ia97Z2vcE/+vBNPaoR3TdgBsWyEmLnb+tcC2qFgUSVzGhBpZn/gaDPK4Nc
3loaDtK9jSsUm9mfS24tVFo/YduT4/4+4lKjI4l3A3RRpXjQA8D6yA+X87UGRd61WRblax6JzEUi
LIlThdoBY7qWe9Zo3RENRz5XWUVsqDHTrqWKEu8UZJRPtWdVEtiZdVOgTi/Bwcz7tcoMySjTMYrn
QpXU3dDo5+W90DYpsRMAbll1xm0b+23VnzcCvzT3Hxm2Yjkhr1B6CgnOGQMvr8hsVXcvUxR5fAin
NZWMv7cnmKozaQXcACNcqkzAwKmObUrP3FF5Qtsu8eZjDZw1BvR/DnVdOP/k6c46N3U6Cl8caL5V
EVGNCNXKfqiiWocId93I9nERAN2mFYivO06OTS0F5vVfClQ7n7dFp8VhjY4tI2Gy0UryWPIoNbvG
Raa12SuCyVuaDRE2Yn9vBbUFAkt2RSPKi/cIPvZ8ZPyEZtnfEUCwB/tEMoOXvskud2gPvPAbR+LG
c134Pgxsy/Q8CMHScsLHYdRmHBpxiPq/mQGSYxjDLnmMiKpK9NkI7qO3sHjoFUOEiTjGDDaM56iE
3o5uXNDmYw3207QkWNlZJgfh3WDfkfti+SrrwloKlAHdTbu2o6aotxMoze9otL2/WBMcp8zqk1ns
AmR+YGXI0m34LCe6k3JfP9V3iEHVaYoeZkGySDwJLJBs+EAZRL1R5wx+cE7YW8vMxnhCbNeAykVx
NK9IP3R58X4d7l7oSQAT2832b9MfGOORkUGVeLc872AnLuyCUxFehyBfg8NIVwNDVSRTkDng/0gW
rbKpuL6M37Ow9dT7f2DXaUpvOQBqTbFupSXqvwXT7Yj8AApO0KFdVaEbuyokENuSuErLNoPvuIPi
oxoA8h2EPpluKaphN1V/Kabq1h1T87CVIgf3mDpiprM1IcQ5+yHQMqwspj8byCXMPkHh4BRaur+C
9XY6enJb3qA3IwYX6wubOCbXC2hERYle4uBuzF7IGEtSNlu2Sxk6423gkviqBP8Sfvc8CfL96rW2
0BkibBAx8hSjWEuwTakUtzzxxnLMfFrjXA6MdvVyRDxDitQsOzmlM6S/ITJS9htsk4P8SxOdikL7
9N2vSaVVAzaLqBKcnTD9MY17VuUbtQStMogV7H/xYra5x4+q0hwiRgJRK2z7pb0JU/A0JAb41TcU
CyR5tfODjiJS30GBCX64tLRmE6hHv+c516j+OHnLw2IJAnWG1pCofXbZGJ6K2MyMkkoEch1vtKdI
BIZIzCnYbjSDEPalCZuGf0bpxXSYCcD1upM6K48hqD2ZIAAdSxSho8CTt6TJ7Ghiq+aditKgPjC/
DypK3Yc/tgxgzvJhxzHG6zws0axXB3Aew/tERnhk2LGjuLtgZlywv+14zg/S6hFBsVyx+3bukBYx
IRAT9KMTKXgLLRhgJAJ/Z6y98waDxTGxtY3yTmCj/xfGQH84ByipISRQ40Rs00oZpkeFg3wyh18G
bG2Sxck7dPE9+Mu7d+Tr8EtJaOW09Dumn4b1Jc+ENwzovz+Z2pX94oM8sps0+MLZbgNAWN4qudNa
8UzgBiZQHE4pviCE0IcaTK1tqPXAATHES+qPpeEC6PLkiG1JzF3Mj9pyy8ywoBmtFddG6yYfxVyy
fV2Kbi9ZrSC8KxU0+gNxr9JyA/ohMlDSE8JiWi1DllyG4MPolOC+2TRSahkRYvRMBDtrLXesOIDv
3aAKIbKu8WUXlKpsqo+g/kEb5E05sXjGljbaaPypgyifZGXMyOJtPiDTPSaCeiv7MNOZ+6OZXuJn
xRvg3OI7yquVEnm7eJu6YHTnvZkLqqGJvrgCIEVN87kq9USaWRZ/7lWRJ0/9R1MdEdmjPC+RXuVE
QY3lrRNMAuCUI4KqSbzH/ucDT8uMhdOLLnBXXDs9rWA1NiP/9WLFqZkYajMWXoJv4dG3txD3G7bB
Mp6fSdyomVQoE61KxF+PvoripjFjQ3M8gpWg4VIPprCf51mmaK5TMIa/pujrIhIGlFsRKaEIDfTr
d7Ze+oSOVudCyMe5FhVv0PQYcaokg4ufuIBDSherafsdF58PDmWbV+XgGFLu7t/LXduebRBiHWdS
nPDSbdLJE72+N0L1/MJss+f6ttu2JfoyPE19P6nmTjFjSJ1/CcI79USO2LwdpLE7zV5WhVG/a2YP
HhhL/UOC8/BkdfHmsEH/TPxtrwHQJ4HonoInxyzpfpHnIaSuL1BVaDyjbsT2/MW9H957LchFkc9T
DkRoYOaJdX39MgHCjPQUu9KGiQK/G1X9cexKCeC/Ftx/chqq9ny9j6lJn+KzKdEHr63N4TdCcGNg
295gzskV3bTHCjAQDnq0eT/AluRvVJBxw+e0gGjnUi/h7LlC+t8qadtAx9OKxYAs2BI8MluLb53M
VvrwOKNSdQ3trObcoftjhqMEltON9q4qIg/2qFrUUlU+ycNuUbFHKQXdzHqM2T0qStUGriuCnPkt
2bj2t2RmgHtrHKF281NthF2x5IKm+YmaIMk9WS8EpPfpGSdTVy4fQjFd6nflnfC5ZBx09k+EdMZZ
wj5z9V20diaqphQuKuwQReTZDGZUofeiyKfuFQiH9Pe/h9Zby05cFnUqLPxQG1h3VCZ3SFLiD6tc
5WLM097SzA5BlZp8ZJMi2Ui0Ar1ikOUUsWNF71u6UWy9PvNOV6/0rXc7+Ryvrqd2EJm3NIqOa0Sy
hRxuSojH+KTNfIy55GiSHLzIG+M49RVwSdc4LD6ZOMpfOkl+zV/gXzZ1HLLLcURLBAt692TXLRSN
/pio5D4YK+PQVDMhNCAvsLwW/VdD9ZyPz4tWr0nDVRbZ/d9sBeiRud/c9d/nC6FRX0aT7LLmeRKE
N53Ae/HvWw5golZTbIX2hVuxhGUnnVVEjY4ppzWDvN7Uj6ePdsVoISrHCf7obSYODI53/AC7t7Nt
Qhe6qzDrA6xW563aBRWjAWsJqAnatg7fkBaMGXzb6GCqi0aU4PxZ401gFt3RFcvrOFF9QurVQUTy
qaq5A0fLKVPYJ90hQGHGGL4Cdi+IM/Bqle3DLU+ibDsCYbgDBdn+j/BXIkVPKMMBijmAa3cO6Ryt
elOQxSqHHPSBNHuWNx7cb4lHbjB/KWEhZBEkwTOApqcHQZ+E23TRGpnYzhFGRwVrGuuiJE8R6oSU
CcCA4Vqh9Y3UMtQwqNpNiXLdw0gvtGE/GJiO4Qo9MUN6uhjDyL0fr78jZsN8n6mjVay4E5ly6Iqa
NNVhAETqge0nTEWlE/rU7HMoCLKYC7RrCB3xejciFkA0xWpnRh0oNSRX2PjaoQc1drzHXJDKFi9T
O9MH85uwICJpjyZdy1mEdMhY24cpkx4C1yFmilDXSNYMNjidBF9Yo96g4EMc7aAstMOiTaNaSAMH
nMzZ5jmqFDI7caPCh2lacrCU+T1vrKPUlK3SxM7Zrl4KwhJhaJDyiJtGEvh9cswG2XDS9+ATcVrM
HRd/3x2LEcMT6a2dOrmFk9u1YY/dBYcRy6zukqPMIVXLvruaPe7Kunb3sNmDUQXuzU6yZD6dPu16
9G4gRyxh2P1WMrQQAHGNVawVOYtcLx1OGFT3etgGQTYlvBkiPrhXQZFEKDoiBsDeMpdOjmWj2IMq
OuoHl1ICYHIEWd6GtaF34zsOxMt0hXWajKv967jiSGh2XpEYfPZKIHnaraQ9S2MuKcmuqqP8L0Yx
FW+e8W74oigg5qsKLvRMiwHOmByQcN7VeZHv4XHJIrhrG89ablFgDtLpindl+dDPkQFWBFJfV/v6
1J9ik0MSkuFyTkf2GeFruBlkWOypH6njRg6HRONh7+1f0IL9kJn6YTAiOQrqL55m0kxBW3Ig4NWn
h/VHz1GLG2Kj1w+9kVHlVYe3L0NCjnJmSgVHV9MWrt8ApnwG1eLGAUOJ68sJIUO/0LghubR7yOMM
CLNhMXxzp6MAhcHLugCN8ru5p/ObA7+pRseZ5bJA0PYJlMH7VJzdAX84At8MExEcN/mLTdfVSWsL
DYV6fzAMgdGbNskWX50b0xeiDvHJ0IMh99fy0F3y2jeLhwiyTCym43l+9g8YRNePlljxpr0djs/2
MjKmq1b6sx2trY2u0WhL5BwEBfkOmgRlOBhkApoaB5LcZjg08au/RDDHCBRyHE2qj3c5/cADv12J
516XofcKPtbHa8rAeLThfbwDLS/QmDeCfbgleqbDJq6DZd6pvS4BncZcgKetT0dxRt7RVytZr4pg
1susFjv6mHpT1vj5+JgEtYzLx6wmvaHicvEblEhSW7qRq8o2ZB3eUhJ2b0Gd6BlTHWiRNeIQBwxk
zmq8bo3ztiu320R2fNkPfgmYZf03cdNihOiNa+satB52Bqft/8M9wh3jRzCBE7bijw6yf9GrVk31
QOkBW7xG8qhJn0T/ubtW/dJrGWjqBQx7vGK3lvmN0fqyJ9YJxO5Iz1NA11PdQ33BFxckYzSnb4zS
PEbiqXcaSms9nmE7VNmup9eCNJtciWiVLvSYTvpWF1pmDSCHfmwLidX1+KMC7+9oLloeK9uxhMRV
DprgquZwlbZMznfTIaOTZatJ14Cc8burDiLevd3xAIw46MX20aXoG5dMwXZ79PFwT1Da/++mU+b4
/ip06rPh/+M1cczCUZmbDX7GOq2qtMX8pl7QcXa7IVpdhr9ZsVTvT0Uu6cj9nDaqpCPy3NlJEjCt
TOUcwHRC4oWPPrVYqjY6zQgwhGNJg4FsXNKflpM5UNJmtmOgcdZJ0OZwwJE7apu94/2u3sET0a0h
BLJ22FDlvCjS7liaz2d1kYkpOsOcPu9xHHCUE1OdxpWasAHSBj+eVifvcLP29+hzrlPhkBL1OVF0
FIpQ//+gTgOyDmECYoF3JTEwcpufvcmaf9Exx8rd3AL4bqxwVGuiSX/cgpL9pvInmZzI2m5Z1rJo
QHM/W/Xv6LllNSZg0r5mjAQssq4KBysASRBxS0kiTYClN98H3Bcgk74rwNdaokVTNkF35u8AVFGc
VZ+hC//n6+knyVtTIMKbfG0lErSYwj0m3jBNp+4wF//sbXacgUgGRHr7dyMrWlmlURxa53LWC5kX
EgIU6JyCgij3rTzcd6c3BLpDLDS4nfiWZuU2Lap39q153NNIojRneVty4fkG86Kol9Brad82xito
NQKJC+0r1MZGpD0ExAT2sns8spGouQu1OAtRGpVm3JkqgDGK/jc22GU+D7zQdN9lkhvGbKhFVutE
vsgNVD2CqRqkM9C0kie05QgHKvG2whIISo7GhOSW8Nb8md+cYAMwAsv9SEtIW4AbzWGIQri956Vu
sawNZFWVnNh8/cX5aiAorjJbEfj253zz5WOsdgCGs7Q15MOEEAjOWTDqOd9uuWk5MNtS2AeOE7mM
jBn35xtFpkO1qyAzW7p9cCSDkZE8BdlFgC27bNmdTlz55jNHq3kJyAzuMRDgblP/Y2WHVKR9NzjB
K8hOXJKPJAC/4mMQaJVTkGE3B9rlEK/yEnGYbfw+k1iuFFOb5IWx0wR24pshh045nmSWmMJriWr7
7xDDWTkzaRf8NSfdy813r6QLmudaQLnkNxpleU68veEsVBdyOFN7FLtmEAM582T2EgxXdgNB6Ae2
OnsCEilY1p3Ou8efgoYqwMTtz8EE3b1gGefpUwArRl76x9iVEYWsNwOYKz2bkQnn9e6tGqgthOBA
f5W0uoxwAhPcfYVodQi4Xhg9yCoQ02F1j61oBmTIIqqNIM3Uw1s1P6kHZcnKN/t4XhLfb/D7BTRW
JX6GptzMFtk70vXztuQxVo2+hh/3AyK3I9WxiBzHKUVhOkDSGSqVpGPvfAWHmra07bO3oI8izG87
934ac2mKNwEyaUuHcrDiRLOO8hVF6p2acW+GOYl7Z3+aZt7gPDDhv9l2kBF6vtZdiFwJY2+0gQJ+
AZgvMX/s4sKLWKDlSyXx9liWWNLCg9zL4Q4CeCjukj1376YGSXNbpholUoCuVkE7EcxHJoE5Hqns
iwloysYuGpLZ+n6iSSMMhjUc4Say3f+SpY0lfREG2UKbqMR/mBFgcT0OQ55GJHzSXQfOhQ+Z/IJ0
9PP7E6mm+ZWl+sdpZQXNTngptfvf28qglkjtcLBUXQwi5oSSBKVvT8jTw4vm4jNFiPllYG9MlMZH
ZWwa6NY5YQr8VMCsuhs6rck0QywZ9L1i8pqyp1SLKrYN4lv+T2x/7LL60fntJCqUzmJLdwxbQ+Z9
aqCcZSpSYXMllakd1ETQfR0hpmy4MAmy8S9FLoAiARgqe6EZkPCXWw2dqwjJphH/xNQEy5szA1SY
5gqvgrb2Ai+l2B47YUhLwglsSBnVnpYI9F1prFXyCm236vwUCflCr0ebxdwNx61Ebt2J0Kq8ZS02
5L8Yg8eAJ53ecvha/h2GGh05DDuMJTkdEsB4Q2fmFbUeP1TGLjjIzXQOP56kqWpbzzFOAnW/63Q8
eyNdRQRAVoMvKJMeZKvcsjXVqx51jTEiVxXD11dHSJAktzC4v7EhkL6MVP/9N9GT6ALgaQk0i7Bd
aWHH9vGd/fpKi9j29sGyKDBilDoMN1OSxj1HMGf8LKuIwLtMZKC6D6wvHIKaqQR61/9UQqhR2ngA
dguGPIWdEKanbpMgPOlS/3DfdF6leVEHYXZJlEKtBapBB7l+EE8gZqI7p8Cu3QhpQV3wV7rzBVfd
sqTn0iU7KTyLYyWpVb1CMUUOlDIcOkwqlLb0bjrC2DsVYCS08WL40xomSJmkW19pnspTFZLEqnuy
+w9uucPNhM3RNn1/JALJMSBmxPfJuJVTnxGQTdhh21jRXqkYSfO2AhyZ77y8w7qd61UgOErSJ83T
JXE7S3ZLzDItTowauCoJRnhWduVtQEt9Ahag+C9Y67cmAPhPS3V8UXfcrBYVDGj3dsNKXmW6pXOk
RIbgBgQWs7cZv3TxYZoxfhVE/zLNvyguErkJTH6x4dVyspHE6TtIMLnhJFVk+BF/jHgRsTtCkPi4
gFvdhkYUjFsD3m7miQuswx92Rju6PGm8M84LnO1FXD8DiQbxUQ3/blymWF8k2rSba4mumnHb0esz
POCdRbwb2flyLKLKiPZnGHdfS1N5aT+x/+QgdjhlMPD0nP//Oi+/nH65uW9LASndPOgNS2vTzg1y
z9rJ6FKFO3CHcAQLf0b4Peu4NJNvfE6UmjU9S+VCeRCeBfBHUxp05DzWhP7TX83tUXHbKxQzqTIe
HE1WLi2uORS7ruo4aCqeFlJq7h7MQlzFhXu8InPvCTn5inzqL8+IFah8FqXKNnvphyzxoreGqVtY
mPyR2aaDgpeI4p94N7p0ycG6UU8UiEpiivDYafCPINuERm5eQ+pKq/OB5Vpq5LdU1ED8QYgZeN/h
Uj+sTkrKwUhUgrZlJUXaVt72pvW+ezyt9Dnw+bI+qRQcgV713k8WNFmC/l3f+UdGEkI8qs3MZudy
gFtkgwxyzTGD3hvnqwiWxBaCzlEnL0dGeGpuHrBBDCcOk9acceOmgMthXDhHzNzbnCurYUlnA7sW
D0WCtHkjOpF1NZOSHIWAC1l+TVShTliOUbUcRjlrIijxr4D7E+VOAbThZScsVlNovPiFfuFtGotX
XhwQN5iFLaKjP7X5UCtaNJ8yYc77bEAzZPY5mXJaaTAAf0piDCgXLTVxHvBBr7KhnfRGpmjNU4zv
3VwU3SL6p9O7dBInqTvJ6ZoLyLHde1BVq0czU/yuiOYUwNE5ps+SxWt05tTOW+sUw5+DTIdFOs7t
mF3ruraM9usVOEeZZ1VOv1bsTGHQXrpFW79JltmEI0pZzt+lc6e7pjdrIggtdHQAnF9rIY0+2c4b
clGEHk2Q/Y+ZiZnjqLPuBXn7sxcryXdjGVgSpT291it2laPCfNPUQIGPnnXaxeFEbEynPg6h+Iof
WX4HuOCe/gVzLxuCHQOH2vM4RrMAE37gPCcbQtSMVqkHHgYZk89CGTTyDPRHGiJ/jNMD+WZ7s+Tb
R4Bd+rqV28vZXPGqqI1zPhFcdWrk8O9gd7iwvwBe5SgrQCuYsF7jevqA3wrvptR8Z+ddXKVsSFuQ
sxvLrIm1p1OIfZyWq/1MQjgxH9/mA0wCCx43l6+gbGQI0zKg6ivgkwqWFURngLbCULmrBvFKrI9c
2YwiYbpz2Zk5810r5EUwZtR00AhxkuIyyE+HvwBpLGMkYChHwAMXG9FB/tiUK0oSxDcUrA0DNsXG
1MM9UScslHj2AL6IrUPHwXBuS0bD1s1Rq2qvOhzOHMyzCXu5gOlZGPEaa3pd4ATi532Iur22B9gJ
6D2TlX1/8zcNgHD6bQL71QZOY2LiBtn9w4DO1Z2llaOroGu5H4ETunOdlo4wkQQh7tuJ+edlxhmH
AHWh3OC8l2TJwv29WcixZdx/acO90H2Mv/kz4uxkr8Cc0IzvZBLXfLaBNqG/rM02GpJJT9Marg9p
AHG4z7MQ7/yWZCG+fW4V17V72CPxdem+DBcbZpDDrAKQfg3+EDGYApSZPXecPMhbGNb65kpoJN9/
VSm6wGUIv0AtMAsCoABSWTbN7Okugf3OgQj/YnGXA03uM0Md6sThua/mPQTIp+nE7Se+90/wS83T
ZKE8zm75BADSStXHDR12+ZvqfDsDsjrOp3DmxcX7KIK+xxo6oFb+kGG3vRTz0aVMdOQC+kF4CaQo
X1mHRBu9cZXGxl8BfR62jW+IklfCQI417Y850do7uFWqHyH2ei66VbPgc1t5YQmQ8UHu2z4oAKzM
+rXH45Tlze54VbxEJ2jbRIwCgCpdE97rTZm7zk1dFEgaVPjMt/2ZdGIq5asJQsRt80Jeax4346AI
ovqn7JVXmLMg9OxHBnGa6ABMjIoVMbc4qu/DYB+yKzU8crkN+GySm0cE7uWtX3m3x/xkLTLbKE3h
fWVWs5q9h+bmWSwItDwLiP6ZNc1TWjBk7plPG4DlWnLl0QxpIXBzHdyv40tF59poCHNAJSreCV0m
fyFZcg/Hlqz1fPUG9rSQvYO1nrpRyYCBszIsA4oLDROT48wap624zOua/ctF8juuXZe9UpgUWT9d
FIvkaNVw6nO0BX2Va1E9TgizrYlpG324TxYUvWYkQjjG5sN/f0uK0d6mIS+vfovvx1FHqjzOSGdV
QZO/Y1vKHQhOLdUDEsuxJElGlMWgOoSrKMR71XpugUV8J3yb6wxHeGqzGCnuEvX9jGuFZ55ysaA5
tDmlTMeM7hR9b+ocfN7WkcSX9KzI9fyTWGAAUmKpVnwrSOR6tePpeKupHXnmuszpPYljZ1xRewM4
p4/l+UIdQJf1+OlsZNXRkTgKIWTWOReNp5Z5c++mH/ZiZeTdrrBZGqJcv3WyMJ6xbQJhfxnjZOux
3FVpN19SbZ/CiTEdnB+NA27m8yXvnDeGLUFnwFV6vHVO03CkjSERwL4Y2Ym8jOzxMTRpTDfYRohp
xzAqJLkkuUKc0giYsp51bflI/F75OGrMVd2R6M2LCmK+g/cUU239YXEqB9eza8HE0cX7gTiLadYz
vk2pBhA1mgxHq/dbrxs2u73RAGRtr41e8NHwzh21tiy6zTpAbJ5luu+UzCTIR+JVLbSnU9jB6yfe
ra1OETjh82gVDAwIObr/uqtCXGpBhc9vuXSVZ676oCcjSEz5B45Vin+WptpxkLMnqmPrC1hFNip0
xj5uxCWlqJHTobX7ui30Z2Wk7HhgcsB0gANrveM61ZYgrZf+7g9Uhj9AJgvLvLJd6FE2z8dvGyDm
yMMt+oJS4/HkeNlLWRapPOS88lFeeetkRcbgNAcKqRwBIBnc0Hqb8Yuj6gtBLLo3vYr91zcgNHkn
wuUrQrL+I4IQIH/naQm2nFRxUVtzS5GPem5pzChJSBIJQgvFHQGgqPACc8ulmoKT1hBc7ZTP3uai
sobGKFBo5KxKv8o7pz7fVespAGurCmx6z5U0mUYLm28uORmZAFPYKN3AyPL6qfcZ2onTk6MVi6bJ
uvAygpC3tf3Jr9aWeF4HQWOULoSRQL1xuYt6UWkNsUjKBxSvG7gYdQE17iteLBxyBp7T3L1q3Vd9
n1/qvtMF31vHZLdeeM4vbiG/ceFd7xIyV1lA1fRkG7xuGtX/QFbCMacZsLXhu+iNUP9sxCqVFfnp
vX/0SLpB+4aPHeywQShhN8wuYidfhLQ2Csj1zEe7dUdCAWN6MELgWQh4RWtCLz07QximqK0B/Y7u
63H3B5OB5OMXrgd+x25Lx/CnretuxNMJiDL3xKXHbRx5Z/1un5Vn5vLOmHIYSC7+CpT/27OHdcBC
ns3+jhRpHhnukrw3k4thRKdxBeaNzcvIkqsTfavrFzgkUcE9EW4Z5e/M9CKhjoIVO7WoShpC0Q8w
hjLJonAlq2jO5DhXmK0HmNjj/iINVjr7bMg85CRBzzONBnlgnSE8rBfdkXhVZjgNE091u42DieWK
rd4iW+kfJbaapN9wklEUwj8bpSbxoh93iWUAz2tmjrsadizguLQNqWpXeSVI6QSkXJfSUuItgDfg
xSAkU7kVnXuJ7CfYW8N09lv8MI1VkwtnhzYSO57JMbxJY5qLFiRhTTvaDNSagPKQJyBpXTnmLvH5
jN+PozLbx/P8moRd2VVCLmkL2s+cuQn1jdqrbH9J4YrqKdXfiIDGkZt4xOrZlnIoEkZ5SYVyEi6D
UR1kqU1tj4ho6qjk7BKzUYoMHLgWz8441hiym+vxj+BZC+so5LB4ojQojpelqvbktXQLX6uNFD7P
u4EKpIu3rwLvr01KMyd7CYpcBg2PzqaZ/yU9ByrM5W2kcsGPYgrDWIL0EC2BYmdauiraaod7ZKar
56yy7KDZ/5nwVmU5BqVlce7ng6ATsZIMwYqFS8hPs/972tympWIerMl2tVANu+dIJamhZhIRJGpJ
m2bNvEnmUlYmAiqUoBWsnBbjp8kWaa/9TU9JAhcx2x9bo1vCMhsxgZUePeMY3GNixF6kmdNQwM4D
XdvXPZC8ssajo+EJ3hWbbAjJeQJZXX1nXZGkBCe0EXbARJey3GPrcA5NZIoY047H9mlLvj8ipCWm
A1YpcGn5HYq0e5KQ7moCLWKh3kRHEpODtupSGhDIWiPe1GDajvSXzuy+T3uaCcK1oDGhKEfBvaQi
AtaKn3pv/AdNipZdi2eqt5Ko1ACrKTA24fSJ4ePxzhzMxrBDcPehaOT7P5ykL0Gu8+F7z0DwJvUK
dsOAJ0gZaYxnylZpfPcqC51PJilS/aYnCWixJArHPThX6xndk4LBmleJBiFbPwBFfqJWA0Y/AIeG
t7dT6xpzQSbJGCTHYJKHuEMH08Ml0p4g4J2UsDwdxmrSgjyqqwNq+Cae4FjoA4JwAMfnQn3RAdxk
GACtnZZnL2gv/5fxdWfkyy4xJQQp3j/Qjpj0m+gPv3zNKghWNhLYmRl9V1bmsJL7QeScOPbGm9NA
S2Q9Jlf6YizdfaVDGfUFjwc7Kxgp6ViM4NSfK2sZ86EdtsaTTXm2ndPNm1gLJN2cESgjUnw+RykN
ylLcYFcaEYmbPRxF/az14g1gmX45dq9qOTMz5GdsUn8AMSXW73ww0qu4AKdQjIo4bw7PRBMoZCdX
8FV2x1GNSIiAaDB3S4s1+s/7Nex4xX4luLTRXvnmTbHNxdnywpq5jh4x/A5a3UQOm199yoKgopp6
TvYIlS8ot4wR4EkNQfIayaKxqHcSdDQP211rF3az61VbzQVNbVMqtNADzOooH1zVcyCDrF8ijf8b
7Tm8sZyavG317ZLc5mOZxGBrnIZ4mrfBwxPHmW58p67m1Qp/FEMgQKC5YbdTVE1LmwjjKuly6IqN
NUAMvjq295Azt3emRhLxftxpqQilGiYL0WdeTfKPpVX1fSl8EqLzP2I5ZX/d1ndCJ08/wHKR2kFq
vhT0rhkwf21HuNG7pBsa5z9eoPIZes6k/gRXI/6sPhjcQTbKVubCSEPFTYjNOfMErYpMxhaXKgh6
5JfPT7vTB7D/tUQE+M1lN7t9pfYqFihBd9SrhlY/q5Of0EBDOcWX/5iXFoaG9fKWa7OOqx77eEfH
lW7T3THmtrNuc9yQodLnKUqwB4L/IyAc+d0PPOaly5L0NSMq1IoyHN1z0qyggkdXo0hGXlyuOxz8
eNpJ4npagW8AAJJQsum6kkM3EY73/d12NrzBuQW4YFvHI8X3guERBCnu8f6zYmeFHwCbOR1F2a0k
ELo/kb/qOdmhQEgKdetxQifZb+53U1QO7MQKe1ixqv1sJYt2omUcx2ilUfUUbeXdT/OGdoTuqw6x
W2YiM1TWpUU8ws9U6mgQZ6VUtgHuEV8R26mFfzqYbX6cjcfL+TNjGUGJKv6akd2AC6eJNQI3NUcl
JnZNYCma+fNuEhZ3jxs2RyuaJMWhPI1RcaDB7y7VSePynKeP8CN1E1us+07yYfrLe7BYP7gOJD5U
un/3vH7PJ/BOtWusR8M/dgkKvH21d80hzoqJr5bVXRiYhNi0WD8IaCy/lFNKX1k3Gjnp/hBea4AZ
6kVKAGhFKv9vrstsmSucCPHnCV1yg5KSMpCp1cx5loJPz5iLgobQDg2UDFlVrqX4tgO6rRz0NC6z
UMjs7VG24iMXgNaQzTaRYfBF+QJoEsp14qeWx6cRn6amV+9sUjLZDzUlSdoAnT0Esgm6MBsBBVKb
yutDrz03WzZ1XBkQJpByxCi5JwuMwb8YPxYlCmkQe/LvyWdXQcPugcVzb4EaZeuZ29tjwVdo+bqi
HTOuf4SOTzo2aXcpQzP3LAYBcMf491zgB5sqIzcH+Juv6DzZZX9Fo3TkSOTMRY2/R0123ggwcPkg
k9HZvE11Yclu5KrJihFs5lNw9YuRyz2C9gMwzIqEJ2sSHDAu2tpvwKaT3JhuD9qBpMOK4NSG6Iap
8ynTG1Nt9doi/cy3D0xWn/Rd4yILvGFPwCjKPrd+uJ7drrZJC74BkRaxPTqMBqd6oiX2fTv5ZEDD
/sz5R9T5HHiqDoBMgyBrkyitdJVrCVYKqrbnVIWnTk6jYJGjyZwxO/RBvnRC9T+1ihKd59hRt49W
BKfs0l6soGGwN8uaDrFMs+J2ZlitS1BpYvGrE3ZaS2XSTD07Uxxxul87IVH6+rU/6wnVViwQ2kd+
544/QZX3L+gzjj6hLS5ugADb8t7VAaQ/yzrUPiZ/8cHRnZSfGHHsUS2WZD4YRljkYjt1NXYTJTjf
TLTTi1vfjJGCiZQHMWOtt8JiEC0uBZuEQYj+FVeiJSD5aEiXhCp4v6l/VEkZjgR3dykeo6K7nGgi
FCkE/Jl9eOEIiuG9GU6HFmnwIrbtA5GkA8NGsrMfTJ3TVtfFxCV4slWFe3Om3g+kku5EJX98XUW1
+HNnyPL5EWgfgtkfMLEb6vZhmv9gSYkGocT64tm0Dc9bK/TKpQozJycyyS+RpjXY9the0+bfC4TF
hwijJjTXw2j2L6ZXqHpDh8hIvJS20wQw4osS3Fl2lXmkHWojTBLfXxdgeK1Ny5+1zF4A/FFcHNyh
0PwNBuEHAzwvogZyn2V4Ep+EN3VPZyqfE18aNYc7VtbwTq4Z9sA46Q9EpHm8g6vBCeU5RBzzpYxh
uHU2vdc+LTrozmz/mKij2J1bN/T0OCGPQoJ42EdBTM3KJkd3/l/mvHCX2nsW7oWOSsOOlK1R5/BZ
JJ7Rniqb3L7HqxvTC87zkbjKQR2WhT/xU/KRtKFcyi8pkjyPKWFdc0omAM5lZK4I5Qyh8MEwEaqS
nV8VLK4v3wxx+0mEL5aYXpb16aLmBo7yrrTgPhs5SSlud2potqNne4oX06yp9LLDRaQrq47LwPCa
sXXZt4eEMXtFD9ETZPxbLV+zROXWTBftEeYJRK3O3B4fXBx28B5+Ms+RYQWmta/HGXYu4sxbUTSv
ZwW5tD3GXGeIr86tSDjdLR981eKpy1ooledPAdrdSF+rrz1omEuIzZcIB4BsA0xysQJi+GZmIsqW
hrjDXrn29rHyAZvtto/xlBp6rwFXPKu3r6rTo1s1TQWpn1CQS4aHF9+zUTIxKMQIjGjVfTK2PfjM
bM5Yewj0uqrAufLXsi8Q31jN5UaEkTTp+skkq2vMUeRmVgzyWWT26KOnGdx5qlF1B/sLyfKk4Tn3
qBseyX/OadmWpI0YGPKsPqmew+aUCTv/RVMToc5I7490g8KHtyLX+2wdPZB9SNsc7cQwu//J6+sO
6UTS13Cl0XnqEn9Cbf/74uPKYlYlzyxxAahyGd6s2TwouZ9RgzRo9htqohsQiz+ZZ70QR+LjjK3M
QFjmApkAQkifvf3TlaXQHZHnIlLtTcfLPgUOVSIPRb/hT9uv+UcaHkLxQtzLPhNz11aUiwsTQDvr
HnXVoLmzmSCp4fBjt64ttpMjT3AWdao9GHYaDIMqi6ZgJviphMYmZdfBqRFqMlKJTBxzWt7Uxhx9
NJNDtDBIu09MfLA4L1Idy/7gXTUhdmyBFc5uW/GUza3ZiWY0Q2HidV1oZVvzXelfKh7Hv21szVy5
A03DaI9bSDiEWlyCghJbV+ZlpzSbQmH3SLO0uQ3pfye+M9MoTAorUTC5fjTiPQtQGV2CnJpPDgsK
YvBFD1mxg6/MgY4hIPLE/2fDua6UggcxdY4rGrx2+n/6s33MX0NF1vef/G3BLI9LcFI8bX7CsLVN
6aGd85vXtXk0r3j5bHDMLEpsImS2uDsizusXb98afJ/4oemXp72Cwm/3WGCnX03h2Dfc9Mrduwcr
iF8WYV8V8Q1LK/kJx4t13rfdzcWbeKUgupri3DjJQjsAl9WhRhORegHgFrPbEiq9xFLYjLParVy4
+KMbOxGIlH0ExJIQB1sa4U39MEeSvMbZx30Z/U4zjjHOYgOIyE9psOZmC89T9VxhqtoyDMkAyv80
yk6C9XpHBElvaNuJzgfY0tPiA4VDN5Mxh5DAEdWUKfhA3AMmy4tVzF8SGNhtVVL/BIEf9ruzg98e
vyYPlTY3GQqGYdwsuDQ6zaNit5UN5Lzq5w0gR+0UXssPZNvOHgFIKtL1Pu4R+jFvV12Z4AR6qx2T
QhRzygEhYr9fquRO9R7lKERYUzeJmDlj+U5n6rgSVSzFafaLPbTuhENCYj7HFU+QpVynHtDspZOj
LZ1mkqgs7p5beQbgJIpRIWxz2Vw1Fz9cbQ+izbFbHEH1N6cD5kpqBAb7brTibKVQsBdjGjeTxhr/
AcaAe7AY8nKCyP1k+0zvfwNRN7/oUAo2Er8f3qghAfcltDVrCXlkkpIcUXVjbNrJceyyDGGtnjr+
OzR/pPxu+4+7tQ0ZPKYyh3yniND1Qr5dxHR/GlYv/xZQbR5qVo92MBvoTyzFIATOEG7yjlcMeX9W
EKZXQ6HmjeTZAPrvuRcyLRTJNqnHNB6434kDTooktgENad3jAjAbZnrtD/lndKFeafXJEPpuBxp0
w9/PPcPv7IbvcoRzRu+p++OzduigmTpnUFop2pjmDaxMsIM8weChfC79HTL8AzALrnfCsTp5mmDx
xN4Lo+DwUvEWWJagIbIV85eoWsOV9+s26FTzIXE21QvaRb6TEsElE9WWN3JvWLi4yqTMbgWaWjIN
FKnuaPPzyw7hIrW2I3aXooG1LfgVvgxzruhCTyyWFB73CBecIMT6CLdFEqN/PB0pEQn9UPVxtLhd
u7OAB6aknYnvYyYkL/t1MHHY6xOU4t/kzTc3ew03MLJ84JxAygtsrflmtfQKmH2ES7EyeK07jOnv
3IkA5La91zABwzNqn1+fPRgv0SV7M/6+5GnDs2L7Jbfurixa/xnGmIjSUjOHixNdnPlz00Jy/onF
n+9KVqufou4NkcaVUmP8Zazr+7mO6WR1A1WDGNnE93dH+F+tqMjjjhGn2pQa/m9wpZrEkxnn27YP
AbPz/sgsUKb9XE8/8YkvZWsP+T/cCwopJXL1aesQw7M5B9H/iSdPpQd1b3YYAD9QYYUCxFEMi85w
JFKdhW6umkYvLN5LpJ0Ru/KdchjpwLZD71nu/9foAHeJZMYYP/HwpziWzMLePrRBO5THAQz/1Xsg
Ko6pg8gZb4RHjrFtRVEM7HVZEAStxjtvMBfLei6/Uf9xFE/oLvD40Ppk51/wwpf9RyxT806CfHM1
2zImQYMDqQ5igz7keWpc90QS/TEZjjk7K3KlCvvw6jQDDMes4Nt25yPTQnhbq8hvPu/BFoR7umFN
bz/hteKBnRmhq98raRS3tX9AJf08fsa/p8t2SWDHNwx1KgT4XBRevAapb74jPhtjUUZNQAOzz79c
MgxCCDJnVRTx46FWKmImwwYwHgoIw5SEncERifnqxpc9Cyk+w36CaNRaA698MjQ4gvNzv7C14alw
eC/ncHFtLZ8vnz9CJLF4ktmoWeToOQ0wehNl80uuvsp+cDfaEfj2ZaKGMo6T2Fz9pSPT+hSWaeMT
JIki0LXFZaCGErYPdH4mx55jdhsWYGaxNBGFnyH7cHGicZm76/9QWghbWXzNQ0Y0DTCgs3TaqbCM
dbWJKBqJpR99FoG60hDmeZ9+dgTXVqkQ5e/EM6jZN4cG/fPo+WX76YOHkCdK/P1lYir+m6nqb4Ib
bR1621PrdkpBCOT6CgpxPug31tXFYOOkaL6il/Atdz9HPCQg5u4+JSCv4xZ0CpOPUhgKsU4KO9LV
HLLEkOcO4p0Znhsk3FH9EOmFvee9+I171volSpzfuvFSvCPvla/1PHRQ6p0XQthFhuYeR5WvBVBg
x9y0wDh4hBrJpcffhpUWwekz4QL+VldB92FAv6Cc1S3/DEK/pEv46q0w3nMdFBkREkMsdqiVNXR6
3CLHG0EPxOPwknN6fyyP+/LRb2HjQO8oowvQQ65ISEmpjnAENVk9uwuFI7alw3CUY3caR+/NqdaQ
t8UuEDoGndi+aq5oFBvzoO5xbMBcizm8pvLlEeUU5JI5L3xkh7fPfGbGLy8JTAaPfmZ5gLwt5Kht
nxVsfml6Rmhzp/0OeDB7UlX9hqnIn6RUseUPSoBSzDMZhAiG0VRoXP2S/3l28Ax/eIJaEaCbVDM+
o27zAWkacgaC5GfM+U921szsvyO6G6Tf88xV+9evuHKn4ogOqKBwAUnfmNSDJUDe97xAv0AvB1+B
iR2bdJtER24zo1wDF/t0uvfByqyQbVmPakn87n9WL0Rzm9xRwW9TthQL89jOlxv7Q7mBkbXD6dX8
mB98pMOky99ya/xxsk6tDSOH4Hxmegtj0YhKdg2nIb/5yNIh5J45o+XTDPGXDcWSZef/WSuh4pN5
8M7cFRcRiV/7Ebqo4qZgS7M7NOjrF2y4god/bqFhWYMIjgug+w9J+MII1upkV8m5CP7qwOCJGq3V
uhQRc57AWuAir9JdaxjmQESSwZu3Q4mqNzDhJ52f+mGeBDHgp9BQ6UEMtGJ6zcs8wZiKbUDpWxg6
BBae8Mrqr2LrQc9nSnEmOr1T8fXIuv2fLdZunuDZZ7I/bBUmGNLz7ag2AykcKfjobflA0xKnvR5U
l+4dIuSyUoi6vLG5OeLof0nc/JsKwnlwrQ+W6XcWCJ7DWqsOxOZz6N/MUJ8unRzdwa5/FC6jcSsE
ExOq9006DCp+cs1RbANUgIFtmFr/uEeC+ZkPmSqAlZgh/srieG+ee1KEkCNyoI8w09l1MddFoQ1c
DIg5eJzsxUzPrN9OnD420dO48/E0vo8Ab4BQ9l4sL8OhWUPioUSnk++O1eYZNwNOK5N7mXtj7jcZ
ns5PoVjbR85XlzwW/+Du2MpDC93zov68nLx9RO2K7fCBt6RJQi7vIf0IhpUny/6bWbPCVMBsvvsi
ybFXQnh0s/CCeQz0XKCU+VAz2JiPEGS0WdDItoCaPLx66GMu8ZWBzBxT3FYOvlx7jDNZtHbNWVzT
sjBwHmSYbfGasmrOabawAFtKku9ZIvOPY29MbKfl4ghrSBNjszy5N23RWk2rbaP8b6vGdIIitGfQ
2uYXvDOBrPFsSYnMCWSYj5XL8pVAbk9gDCYluVZawFMQkjm1e4ljBI1+QnoBqhYdeTrKKrJfEQxH
xFVKqwkHfwIkUQB/bc6BsCsShI3UIQOtvROic8p5gF1tl4FLxZUuxSqVuYNfPiMYzq5VYha4zAMb
ZN7Hp+SYB4JJkqzw2QDRf5MtzU2PHrlbua31CXB/yTQhd9LSIo7X1EZoa/FQTB2KOHXxO/fjQWy6
4WDzl/OXnpPftUeuvqCvTXMpiXYJxGNr+XFHn6qDalejvCDrG0lswPe/retdftfNy02ZLDBvWgVd
n8oaOGFVjmBZ8ap3BjGURsJxNSWgvpYQMoUC2ZuwofZI7LPL6Hd+W7BQtl+UXZNcix1yMSuwajTd
TDqfoJwBIwxKG+5YkN1YFh0Uq22HXBaeD4c7XsyLiGnL92PGXbPE9pIB+7fC7e9cT7OCyTO/QkzY
g38EL1EPupcUwVfjfaCvKe25o+VpQrLuqgxomKswoMuEc3CBDPHZntHbCRpeAf+uGzvcId+FHsP1
up0Wl0NiLzkRGonu0NXhwmQEKC+QmWT+hYDttvpndMzd6tJ8h9YK+nRp5/uUdad8yv0JTpaU+tXK
V9rYoGrPejZn1H6fSjLNCzgJLwe9YL7Qc43ZyC0cfLMvnLn7rQ5YnsXIJTJ+6018+Ssnboj99YzA
wGBscu3xDpx6dn3MNMHNq45QSHw21DV4cFyjMh6ZlGiOsTjoBR3rusQhhIsoFpje93BppZePem4q
yl+LE7ypgb5Zsq7eLu5ZS2HpOShgxomEmy3yStBqXHMFOz+cinQORP5y40BCyrjLjkw+n8ktB7cK
yGPt2KMhC+7mBf+bIXnvYbiMq+QAd+TKn2ttMS8EFKZZu6KazCsi8TNt6vzd/pxdTMJbRIB4Pjgp
+tNJStakjfG6zU1ONgUQEOD+06gHhgNSW49kdvbcR0qSKdUDiSSLDJGbyXwpIxVQl1qMJknnQKS1
fn5eEAz9j0/IyeukqkFpSIvP74qFw+8+7gkyeHYyetzam8UUNnmOot0ZvVibrehiyK/sw5GuzMKD
O9XmIM0phECAsS29qvQ/jUxKT/qzqt3k8CHPpXB/MnzQg/uhBh37mXC6nG2/vZ4QMfXLrYoJ6T+w
4OuHHolAIO7LsIft4ilGcteBUcPtLHGksJ3qE2ZcYFCCxIXlWVUF0FpZjJBCcwNtmhjJ8CV4kz2K
fSLUmX7qgggY3fipNVwuu+KaqwckjUMJT7j+mzh9hnJde9Xv+FY3QUvKd4Ti+EPcpCT13vNnx7sH
kBgeEnbMsbny+XUmQRp36b+WLqIIAq4A2GNMd3/ij54fL+xFo9gu/e10VzeBt4i1tB0VSOOxTnpC
/gTxifupK8Vt5q1uZALbbQsahn6PQLUjBj2IcMGdOtf6qV1+BXV2b6gA7vRTdAcnoBVoBAAM9cKX
6IjAIxuZhAuMZi+CrdV5bb6U+zKE9HkO0BdAVPfF8cgCuutxQOplPtrW2LmFFLI49eSN+mVtXNuV
FhHkdlHDz38zJxy8gebxODlVBGleB+gljASMS0QVRKXSKAVbfhydPQ03axpeYZZJw2ByqfUm4W2n
MrQ3npBOdnDaOFsMZCiGb+t31naq5pvQshaiDRyM0VCZJhaTRkK3+Q/LfgBhe2e3hgsSnStsv/Yn
o70gWX1OmBi1COyCiiHK+Gam1C93EsORNkudFAiX2k/bWqwZFE6yXwxEQ3S+a9tte2YeSGXbcqOT
7QwVOrCU6gr09hWbSSPoPSNrr1zqR0E/U/C5a0b2mWm4B/wYIfEpa3LJ2/a9rZSjtCx5m2WpZG5g
toWfHOBURUGJDc4fSbs5zI7jQ3NqyNUUamiOUZsAbZj5VvC+hRon7DPEUMG4IIP1fL1spKk8WjV0
NyB5TSHRaERa/XbgC+sfIYsLdFplt/HVs+fTf1cncVZsTKjHCPlpgsLEzZp8FlagJP2RIoSOplc+
1GgNOuR7j1Lk0oddXVIpe+dr2AmUpR26cAySVkVTo1aOFDUoR4Cwmq/n5OvAyCUWa1QcCTiF9fth
dY3DXWWxLBLLvvDq9OBgWr6mkS3/RdrADNEnXnuwzHSM9VvG+/I1mP7EDLu4wABKlUA7X9/NqJse
iRuth+RGrn0Q4FwGOJfpKzIVIrZI9B73VZA5eGPx8CIJSS2ozsK04CB7yLuVP4j4XK15h5zNN43Y
T2/Fon6b4KBSb7sfq6JSjvSiG6BHrbM7dpnl7fO3+6xzNBKBY3Dld3ke+zoL2/hW6Vt37ymKMY3U
S7X2US6iGcvJ9hD5Du1dr29KSOdIwuEcw8cN29DMx8KRo2PfRnLx3tYUnakPOUCgg07kP+eBLGm1
O970NQm/1uk3RzY2E9VW0o+uN9YzaFG3HHW+0Ga6KryTfP3rOWZm7c+MOcERVsyHDq4vgBA4O0Cb
iVxrsf0IPjj2Pt8MG/bfZlo91KgKVGipzEBrygoBUVI1dVDkwyYBdpYgPm0sQwSc/Qol55ZN0LHS
HcGak+Ci/1pjVvWPrFc8Ds2pKUHYkSUIxD33HD5AfVmCi3FVtgfaNj1zqHwLB2G49+kaUENyWYFK
t/VnvlFC02VlxuxMmcZHtkII8NVcPoQySMt7YG+HRp3rGpb6v/erceclKUVhH34XJq1iTSLe0E0m
vwn/t8mPOhclQrioIXXkg0Hmm+NGzGz67VKDtZ2bFOfPf13jom7Sanf1NzmlnlqOCTRz0/MsY0aZ
XPPyNaqO/Aw3oPXZQlPMdSeE32IdoPQcL8I518FbHkAe85g0JY+pMBstW8n5OZ6/MyuGF6t5akUq
R1AM5Axm2qvNpvhC5CjROYVLm+SIKzGnWxoRXg+GNNW3bO6XG4iUdx7tx7ilZUwRKxKVLPVORGHK
ZyJelZhzcAxsegfSLUDZxf7G6g145m30xdoGNY5LvNuyf2JAlL+SG9r97x2GKClkdrc6l6vMjOn5
46tEhfnZppKumo8cNge4HKQePQ2VKBKSdgb3Ct+t6NGaA9nN71uapgBtINF5p7CBUyNV+MBAqP4X
UWqVUDjBgF6b8f5PojOtvmGFh/gVPLRjWFulOqsutLbxRJWx9cDTLzekKQg1OHCQ7+0kPOhQXfko
uijURIs/q4v+QtU7SzkSv1U+XdPsQz29BxwD+8KS/UPrrLYzPjN+5XRQuTq7hEzcB+6xrlYUYQWI
0OCLnHCpCfJ8nceccPaOkCcyY8C2F9amSGONS5YeQQnSsLNHUyPrPCa7Q4fvxDB/X6yKCfacX5jr
avLCjPgKt9+iwqdcABw4bXnOx6TTbo2vQYRsDMWd9C/Zs8xDlIUReE1S6D9phOAs9kshLVDDoReo
wM8Q4Zy0CXZPeWbKb62XeB1CSt/AY7O9FIe+t5E4AyhwWew3+EfdH7n/2J2CullIPxPeuSPiw2qB
SGwwJf/Hvv10uWU7rV4g3wkjQWssSNou/uYJyPXv6UqXX78DyhVY9Ejk3nxwlyfR03mLe7uuJuM7
6cd0uKHCU4sN6nHnnIXM7+jezDgE/7fanMl4ECVYgnQSthn1HSfIwfGS7xOaPKELAVA0519p5c2k
lGLQcz7fgk8eoECVuNW7kl0nGFbhNJ8aeVvcWd+byRpJ48bf7a2/komq0dLZp0mUOXnTtSVO2RJJ
6Z2hzynLC+G9LfcUC9j9B8WfEqGXL/8jThLPWwFKVJhispfuvo/jlBk4SvyLvVXYc9uEDEsJEPSC
CTnWHJA9PMlyIafD7k9/Ux9c3Dyq3z2lnp3w0aRELUmy0oN5DTXGGILsz9nudHz+q/LRE8STmTSs
p4U5quKIiTkrKC9JyuJF6yMk0eh1PViyPI40y0WAd7V8s8odutAKYkqktFjlUjj5dSqArHPF6xot
XW4Vf5bnI+4+D8mNHVeFnJHbYI0aSeMh2LmgKDaQwW6bqqZFKBswLvCpFxTmUiaEvYQ4Wjcl1alJ
KOIMkiW2MQ6CY62qGF/BNrgfJFCs1uZKAZJC+/c3DnVZRlxyK2DcxS/SlwvRXgT0bTdIHwfqIJgv
uauC692SNIlYzX36zsZbHoBEQ0XDSdEpaSKNcKoIS3KLPSekZ7+OO4M32iF2gEkYnPMa9fG3Qbf8
aYugqFlxtr0NTKR6COsNZiDmGGhPE0TU33nvLVMW6PAXocMJ/NErLko1WzQt3Var8c5Uv1qtHvo9
2PRSUHXU0eXnV0GyMBdact55G+Ug8iOuN0bn9My6AYlYUfCShmjqzJueKpCsZiH47dsxzXhDrEz5
ISmZHG71DdIXyWJMYv1LMmQgpPIIZzlqmTSw0QMQ/fYfvltEJBxgz3CpUwXE3kjr376QspljL3ff
ImfCA49VIfkHjJumaqDs2R+ziNSMwLkgcuuWiZsHF57moiaX62o1uEn/3ubAQq0T7qub7oGdsG0T
czwazCjgb1ZU7wVoCmXupTa2a4FLj1UKLa4hMZnMuH7ZnjytpgUm7KjjWpjp2jhYniWFk95Mgxtf
mXaD/adLNexs6VgU4Kv9V734LwOLNHPdg44wWlm+TpF3zCgYzn1Tkfqx8SfkT6OKilNRbShq8dHQ
F2qdgTC8KJ93h69wqEquIEzpjxHjq0DuN9MifxqDB02gec0S0qK6T4Sg2SkZC6y1qj0+T1PMkqUK
oTCGQ/YvHrcUDsu96+XVQZpkEzU2B7xDs5y/4uE75fK1o23vfJPYQ6svXpspRwiN0IiUheq7pQk4
QvO0J3mhCLEqRY6JSV0MCCz/rs3avppzwStx3yQwnAsU3EUBZCWDAOOsvIjW/A8/9DcSgDexUoRF
qgjFeZjwv9zxYSwf/9u6T8xkicuIn7fpFFcz/5U26IYAps8aQoMXTRaCOIl/JO8HGFUDzaix67vi
Sjnk82AunKtg2I48VrXK3N7+3cpBrr4X5bFiQtGuRTgvXaSd8fjQH1OqdKSKY4irIMaaSumdV4ot
u51dUU4cLFdUF6sll5fmSTvYh/Bi5kTMQ91b9n/yKdK+J5UT7+Us3gMrl/QGq4PxU3dt+P1jQ7oG
cc9wOExgw4FzhHddpidlNq6lkr6sH2bxi2c4os55HGIZ9wbM7aC+KOvFok3C5uR3CTN3w1RcwSrF
LasnlOQX6kDQeN3+x8DXUq+c8w+tAiierD+HTQmdC6+z/7R5llw9Z9dF5AemvEKYp1oLiI9/BN1a
tjivNO6xAtY7rtxgSjqlqA6HL64BHnbmkt+BFdDwjBDIxdT2uq786xwzXGXmqnaxCX6zhwfL9x0n
tmgFvRaSa+BtkNyP9JpjjQI4oYSjHZsIdaEloK6vNU+Ia35/VtoeK8aacBJ2J31o9p2GuqOPXEsA
8IJRLY0LXYad2LTXd3KRTDTaxnppfzfOvuD89iYEeGF5p4Lg7kGJioBHPGnAQGECk2UafDdqPg+0
Q2G/tC0kCoY9A8OycNNLO5mlBIm6HtoXzn5+9a3wfiwafRryoPIvtV37Sj8ViU6L8eMNbag/nrNa
8bQGFR6eAXvN5o+I8giE0Fal20ZHtNH+uSRQDZN0OfWGX7H2QaFACl1xBMagQqLgoCy6iFvsjGxT
D/0JjDqEbg1pdtoLVur73vtOa+aomkxxreGVCt21ujGnpL2spSW2a3j5sOVwuWWEzTQPPB4m0HRL
+tORuYpDt265qcsKfBl7Z6qqxVVHAtuwk7RH02Xd6zkz9Gk+uhIlOjOhmxcb0fcQk25BsHbR400p
ImLK04SGyJlNwLypvzlq6S2L4EfDc/yxh3qxeprWFa13gZSopYdHhZ093T/6Qts94M5Dnv5FlzyH
DYlWNxPTG38c/cOZ5WA4+DIt7I6DV0sypRJb2ZKN6fN4xYgY8yPRAjq8COJWh0JKmbZ3JV3FGsUm
kKkMvn/JbJ7PPE137ORRnvnSG93TRuJiOHP+vATX6wZQvPxgI1MUhcnnUbGUROxxwHAoejSedoZR
OYKCOGu9eZ1OE41P6QpOxcNqUx+y1/1E9pjbrI4VH/Qle9KNBzIWZ3b26OPg60uMulunWVw2BVOs
QPFfTQZptdcC0SLpf8jFCGYTygh7aSdrqqosE/hKJfSLWsLH7nWDyC4MXDqeQJ0rCVlSQ3wb1/Eu
ZZhumOc0sDOKfPOT5ceL9ZO/fcjUiSVhIX3+mMrSd8TsLACDg36kQAGO7qncNB3PZpD94xmeHZIs
Riqb/mu3WIBnYo3FkdWexv+1CuSaWJ3AMWFHpkT6KcW1whHajSyVC989nhhoGYH7SgKWBvUdtFI3
64tMKTutuCLew7X3UWiGqXycJ03BjaP5+FkwlyZRfgxVuf3fapAIwcZic567UaoLhAwqq/JkT/qh
QFkA0Y3Bh0uzrNimFpm0SSI9VlvylrlFo9YmO8wg8EDot/6Q3REKLJBl7htNGbxreL6zZdHhaMBa
3Cb7O9Dg2kIO/WEE3Ce8dXnpejA45p0dhlcby7rDVDQgVQsvHupuWlmaAM7UGmNhln5Mu0yV1SMr
geEZHyqLXwPdf4CCGAV9ULfC4k+5WpgpSuv7IaA6OecWDn+9+AFHbVeySPcYttN/qr+0hmDPKR8L
QcEGrEJT+A7ov4Fk4PyXnUalW2BMMt+RaCV/NiuWiU0/+iVHblFmuuTFfvHP24YPfbB2luSe5HCN
5/0hnFkBp3OhqsO4Rqmqik2jYQBn71iHux80vcXGm6CCN8xHxT8URRHLL8OqpoljMi3jPq4dACKB
Oc+pyFTVyORoqpKzHnYdw6a4s7uLiD+OblQRhCIKaiofYtC+lFHQFM9UyFcZMaPbMojA0wUYKWav
uH31Az9cR+9/JXF0GSkdoqCv9paSJTIxj0gXmWwyEBxIFCGNZ/IsehIc79/IOu6TvOnI1kisa+zW
iRgTX8scRfbhBA/mG2GPhkBKDZpAUnTBgg8QUtuqtbcWGzVACPzNnNEsiGIrEzx9EnbR2O6RGVE/
r400/bMxj3xBoNjMnc+4tLriZ+7oebn13DiTw9L8aKmGCV1tRauGTiMp125J+5v3wH2+dYUsLT3V
qoB4KDlNjWHERM+rWzdCixp404vtb6/2/jausqLQlBqDmMALU1CUeJATqoBDou+eUBImMqHhuPDU
A/29eR4w2RPIHLIN4ne1LTbNVeDFXy45Ic+GN0DSj1oEEwNhBLKypSt2uf/hAgtzL4GyFut5dUnS
i9B6oipCl3iIPpIU3HbbVjL0D9/vjHhScOsC2vRqcplHOoRYPM59eXzKMjVEBZf0ES8KXFu7iySn
VmGL/iRGN5HSxPQoHOo2ncHyhEZ8CGBruMonUzFh70EFxn11znTKxStiwFlzRVAWKMZOpoqFZtvM
OOXTqknZZDHLZhx4P9gi/OVhElz/C/5v4NdedhmGdHI8nczA+V1CRUpbKaCNomGlPK28Xr8XEQQS
UKaGEZGAAkAlpYNUlze93NBAs2u6fqw884Ne9WLXaN1J7YsteoAIzfINK9RiN3aHsunwsW0Fj8yL
6J9GFptk+07V2lF11zyYvI09Jy8JKpAGWL2jMBpQrbHVtJ3G5SJ9+DZkmbZvSVuxnXKNAuwWmvvU
i5vvwC/E88BkWebz+bUFfdtbFIPR9PVCgSmDMerPczanDLncgKjNJ+/aiI/fhMy9Q48qdtsS91yT
TGJPY4vUfp8V9VT9/MWQLt95w/L17nGu/AXoCWR2d3jZudp6qld0EGD/K/+St4rL3DG+F/LRO4Dr
OcHPe40VleE5gVpoPl1WHq36azQIPjRgOKBgaV+8+afQ0gKbmf3oUtdsWG7qAvJKc/+rwzIAZKk6
cmgxO/oFOMXfDfwDJumXrp1D87d090B4wiCWaHAvyh292uV7P8cKmesMoqc3DDKKjT44bXo7C40E
a+0DxiAgQOOAV02of2ZoxZTuOSLXBhVgHNDHadz+595xqJcOGGrvrxtNMrblQnVXn1+wvh3wgr7p
epWuo8FLczQV+dhtUi3nFD19JqvDrkoXMYX+3SaG7+85T2BYCn2BHglN15ExVkxpnBCdrnBc7fTM
zZHojjVjgv15D3jNZ7Pm5XHV4SxAlkmt2zKXauJ2rl7zq5eEsunOICt47VXCmQ+rT2TPYldjBJDX
JpP9ujhiQb/xD8/5p2wPxpC98Ms7vY9lP1/k6z6dHCyLMXPN07J2wCVtpNdEjXWfauS2+KMm0cg9
d3bcGC5F0ogka/OGYX6hPG7M89DXhyK3RnW6fzhtpPk8OryDi81qn99gn4zdldHpmdiiWjpNIZSV
6HG3iboJsSPN5AWWRMTTWJcbTUoP7AVkXQeruQu793eeZcygp6sP7ZbtlFBduIa5c7UxgxKIw6PD
P5s+Yv7kmNm2ODmVWlUcsMVz+Eq9wsrooKPiPpugCMSertHpUmqqR8ctSUZtLQg0OGwTEampOtuA
TikXIfoKkfqQQEmUyRzynP3YQk2Yh1ZoseUWGJJ+3Gk68g2VTKzIXb9gj71NDcsOoSRDXPMZBhoe
5TZiQCqLqx84bB/3yfLVxnk+mmGakzC0+Z3xf+AglsvlSiICUj+3jOXR8vjLynZ0i3xpzk8z2hRz
Rz8iY21iLXGXkq0M4/MLG09WnBls88tmYFdPXCsqYMR6QwgtwQtQ0W1qVmTKi8QrLw4vqR+Ugcta
lTDbEGQirAr8AIU2JCxeLfV6ZhEGC2DYrqAYHOiUcvl23L0V8S+u3qtQyKrBVCiJTOLZ8ednvkoy
LHJ9Lpk2/1y/MFPhskFVt+clT1xpea+n7LoZ9pVV8K1Mw+nUJlYSsGQWqAWXuW8Dy0AIT8peW5LI
dbE0wVDOYSrNcnJELAbY/IDfidXcw0G+2V4YtyR8Hvg0aMQlXyyrRmY/8Ivp5KLyeSuJZRHVtBVV
hEiuA5MiUzOlBv9NIFPoBzZggBclQZFirp1GEi5g/xzvp896pMndMwP9HYIRRfRacvaENMD9ztoL
kjpn2iqFyfsZq/G4NifV3ZqTZ20YKjxykd819FBlI1Sg2R4cT4fRzfe7+UR+P99CAO+4mzd1LFsw
P+l/hBVErVPg11Qj+ZvXvF5UKJy2prCmH8Sf1Qw8sD90S7Clq59wsqrrTu8Dc6Hhz39Wvtgs3p7V
j05if+yV7ibm0bXEhffrSSRlGXdH0NDK7gJ7qjTcBAbLLC5lLX9GOZL/J/IUnWupWSMH1Rg+aSab
zbDgqTJPzKJdfLin+seNzf47GqEnZJLh2OgH61SI4FotJonV1bvdsWhcEWLzugdrVDLpNeonkOpS
6ZEMXW28yV3wbOS/TyZWTXNvbwPtbM3Do8K9u+zh2UZx0TFmCOydv7xP6iAY42ej2JP3jJD48Yl+
5nmyEXjTNSnQSsk6Lxpttm6nAqxtDA6BrrzULEDtpeF0FDx0YGPb8UmKrUmNZsK5aqqKRMVHnOYD
9oK3iNtxAJ79HiiPHpur4qtzMzdz0Nr68YelLlYUPZEGsxJFdBcut7G1dU31bmclZQanQUXCcnJ/
neXS5ftOldwbTkAjl5dqKAtcWOLi5duOg5fTcHTovWWvyhJOVWpT++UZLnYQgQWkaEjo6v45WoBS
W9lX8FgItSJ/8Y6xo7tet3jPEvSybQE/itCbEqgH3x6braVV/ikB5ZbrIfiz4dUCEtG/zplhlpZQ
HYLuj9PXRYi9ykF5EBTKjqWiXxW9dq0U2SwEw9/JdQIv1zwlKYX2+Yv3KfaOBb96TyfV1SltqwVP
UHdngUXkKdBoUiD/C8ICHMn+OL25/LwEQanML0TQdIo3Fw/hvj+3YspC3pZ1M09083n7JxJFWMl1
RPDKShxrAp9krcBAZponUQsSEIo3MPb4PRWgzJqMbU6Hhv+3wDHRvToXgEZ/ySzIs5fqmlXHaBtn
Evsi4alDaJ4DqlJFDZyWyZ1NdLb3LPhZ2GL61CXnDv/cNdB3C7+6SKO03laV2+90uBaamZVXN8eo
bpcfmhK+iOViCOPuo1ZVURPxHdpYJzlsGnYKlvMq9l+AM8v/sEnvvICR99DbA1HE9GsMUiC6rNeO
3LgOn/+NKtDQju4eOXVITF1NxsuEkCIlJUx0UY1dt4f+a9ixvwc5yVp/6dntoUIpUpEnHduqO1dR
Y8r8LSxSF0x75KHyk+x+FDQZ3mJJt0JYO7WdfdPRk29fdljyWoLsu7e0B71HOjQ1O57DuyV82qDc
n/x9Lrtw6q1TReCA74J+0hUzZxFFs8BrbnerA95YC55tnr8gAY9vq/+NzTqmZt7mYEZKeiqNKYE9
fabYqqPQW6scqZt3zXgRVQD7pHLddK/efUKcfBcF2x2we0uAu9xuyFSGcKE4RVEdfk1C3ggWebon
Ot1vY1kItiErtYQ27JE5ZbRlFdx1kKLu8BCWJcrPz0H3Kzw6MFQsRyZJc37rA39r5PYd/XzrDLef
GWClhYLE9hQpyPdnuHhDzTNK40zXftokGuFWH0JZ3Al9xX3iS/vqQHFR9afVgmhenrz+8mIGUoSj
rg7yYoF1NWaHnZYCveUKMfOz2enTsTn//dgUdTz8klTTSvHSe1ytOUjWME499Fs5Fz4sni4z95Mv
h3nyRlvJnCrR8ypa/Wh2Dh2C6ncwgGC7zST2hkb/LBaydbA2OjuMUwEQ0+22wUL+EFIA6Hu3M1Bf
lFdWyopIo6/3deWbQvyUUKXjdhez3bqyiAIxaiqoJFOVtxmCMAwPJzw95xizontuE6u8Xtavj7mj
/KGEc+nPunsRnBLVe3/i3i82dmzYuo6CZcFZdgkoFHzLWyn3UzOc0w62VRBn7HUIZ1tjifDTz+rW
UCB3Aa6hKJ6XOUUynKiGMhqKA/hRw5aXF0vJfnlzCQjtAXJisFsRQDL+cB4L9uJtCB7hq4mJfSfN
eJk36oGwJ1c/k/I6wDnP2ub+Nx72uhYnXIqA1rx5vyVitIBRREAZq0TjUXVC0q7Ku3hzIV3F5sxA
1Brfz/igmc3bEuNMEwCA5R2HQaiYP8OFeR20GecJm4VMo69XASAXI7G+bJ+eQrF7o62fJUmB3YPX
1RsWNyIWnEd77aMTaEpleki4PkaKdJjmSApAv7SZlDkHXNj+3IzH6lVfqcssQgtWzl7MFAHpElUb
Nfimz90RfqT1cTOx+vPlulSrO7a1H2QoFq4DWqRHDdcb8d5LAA6ShI5ke8ppOoOHjXC3lhFQFtP7
6p1LnqV1po2tbnFQ34hZR5K+gPrSISHZI3jAKbYzxtLcXSh+pBridzTf6R0ZRRltLcMI24kA2QUo
1Zn8CDCqWAhYAiIwFHa43zjRTS+/1zQmxgnUK4OBTLTKQ8jNuvZJVAWL3dZjb9Yz2LPZ3yykdfvN
XiRqM/QbGvSnrbwEHigMgwdBK89nLilgqXP6rbqrIJHvccnIBvvjJR69FtGseUKHsTUPsRN+yH8a
w3mdva5z0RTj4YdvzO7jap5wWIRkCcyt2H/qsbUj62MznJ4ENl1Fse3DAQVihdyyTv+WE4MfRojK
HvMQRVrRoAM9iz9URCJUey+qdnucqn7tWpHpzxAfRC9kuiVMU3O3J/RNoTC8jm+tK5zl+v483IXV
pgXdH9pCWiyeApwfvaQdqxGYSqYjYZuIKTBZ+4zwxY1g4KiU7NCKmBQLu6Cexh7T67dLzXYaoXDo
eKFK06FUFyVHDe4LotcMwkt9A29/7CSt8/S6ojS08IZkxcGSy9MQ33022bAde9G0xMBW7iPyi9ny
6qNiTW9IIog6kskc/IjXqiYAyKN+EvelgsnwLTLBwoGQLXUEjW0qYZiA6SnRjQ5Y/QutNDYJgRTR
liCM2PFJbOjC2CZ4kQoU+Dzz76z+nkjOPrKgitvbQmK51KiZ6rxlsj0Y8hR7aEgexmO3WGpewBf0
Lfs9wYBI21ELYZxcNwjIyuRt5Wz4yZBPbGeqWQAgAKBXgftVyTeiadQrx0mVcC9XBOmAbHV1SE9Z
giRAhLAFHA58iLe5cQwVPTRhRkRr176pZP4j33EEvORYXJMLj3X7DujFMoZjNnL9TApIkfZ78ZT/
7nOPJIG1Iu6fWjX1rSZ696/AAY6ybTMf/OfVlGloC6+Zm08feMSolLsGTZ1rGFSP+2cE3C7fcgoI
UcAD3Ue1naDRv3sg76Su+EVwkxNtUS8odpW11nAXHul8EZTtkl6onU4N+3bdw+gMNH5eIQFezMVp
b5CZSysVQJLT/QSEOdEoP7afj/8yUJXMnZmWg31gJCEHrlsnh+dAIj++KFdjx4LQvrxO8h8dkxWh
A88nyFDzqXFo3HCUuKp+dkcVxZnnouJzAKMaE7Hcteuo7tkP5F4pMCiqPQzTC18Y4s8ARc8/ZP/9
GnySiJCvyeQntR4Be1iIijsgZOgOmV3+jAdvQxZk0GAJKnweAflbji//wbtegH6vOP53X0Y8yI4s
JoQ2MvG8hhVao0nnTBX+zBP83Fb8Ac8SraF30P1vSimQovlqlTLI7x2Gpun7ew4Q0fTOmpHHNIyL
jslIOJVF84xLDjWc6d1rBx4B8o1Aci94SIswiQqtOeifXwkeA70x5njtZvHkaAaNYU+tMgOPfjKk
5Iq52mZlhYhLa1S9ZtmSyuslNlmd9L8DE63/WbwF0/ZIS2TE9BXWaOTOVHT31pNxwduBBJIABUjb
jiEYIrkky9Jw9s5NNd1i1PeMM0HY+CXALB/l6wbLoS4xCmeonNNvSfsJfX7t1BbW3deNNcXQQBqo
F1B4CPLYoJW+ea+KTzOBr6XGaw1iWQ0Ce7Ab3RfG6wyhw9Jpf+Z0iEODHE3IGpZhQCfd60Dbx0uY
cDO6GgXVLfZCEWj+djBMo+CGAgwJskSp84cj/P4sQXydqA7f4I/ftA+7MfHy2sLThFNTrLz7qRnY
vAAi2SZ5BCtgZCIxxcZu2BKfYqSK7KOusPbUkLa4WyyYsXJYnw7SlHmlzdbexZCEDHVzSI9d84EA
lt9jSf20Qq/Yfbat9R0RJcD4as8TCn+e0j+4PqqAoTFzFLmg9fbIbWRKoFe6jv8qk4MGSV9FsnzT
tO46EDbEH7WV01sVae134sDCQGXzSHOCkdCmq+Nhekt47HxYpPGF+O9A1SOxKICh1RJbK4q9PTj/
anKNLYR8Bqjoz9pmQnxGPb0tBZOYwtqcsjGTTyozk518EdrM+2NwNxYXImZYo6fm9XVlyxEKsGjA
tgg8AznX7YVwvJ5hZOHBEEWdjjoItdEDA8cb84znmmzamOg7w59zwdQTV2V9O4FbQqajOzps+a/2
rdjUAW0zh8NOtX+G49w9Z4ZB4mPVO1vRjbG2KMA9C0otQXT8VQdjVd/79cn2kqttARACs+TkaZxU
GJl6KJ+oMZf5aNwEh3z89L9Chs/R7uNMuEwAT8xpPtjoiqJR5/9He7PVujGXtyVhSfxUrcAsetdW
pB6zr6byOexbA7hGexCJONu4EZIW1C/Y+0YKbr+oNQdGzWnB68TO0flMIQAjI237EM+TZVfa17/I
3EJI8qrm7HmOJC8uLkOxEBacN5PLOACjJVa+Wlvp0yuAUEgRLW/XbdVmc6cX1z6rSQwE6+p3dSaY
nGEvA4YdIfatKctRv1s5bRhwZQSlst767BbKVFVKOhKKfXLcOf7wh9jQuN0sGDK/QSBW2ADkETjF
4NcFODWLsr1EqqboW89xsR66Iwllo0dGfpqvqPjcu2wZnguTfWbAHMQImvQyWAyK9xbdxJDvBRxp
ukpE9mn23ntRCURezNil1Pyfr2JFalUKGNPDMeu2eQjk6tc8C0KStXF4zHJMaMXFBswpdkW+viPv
Il0l3vfwDafEUAaKiOxEyBm0BhqIySdmCl+cO5SOdMzgn9dEJEPoCm2v3zl4mTHCYeVpKUlpxHNp
rBbLP3ELsPzMv89HADtzlBJnH1MhJE5I7VJVMBpstHE1ca99f7/NUb3FIxPjRjbBZT7NCVKOnlzI
nNUxDO/rlPiW5GOjFJaem+MGiVnsnt75JQsi5aARDIGquZHD5w8G4mIeJXPu4vK7VJhqauWhawjO
WXEKfHCgVTBYOTE5ktXJyquk5acpek7ot0xQycP0C2Pcr7/tqjAO4SgdbBIcpyM234pkwOHCnXtC
PAkvyroYRw84kvITlF1L4b5oO3W1bn+LworcqrW8Obe3ay3BMzvx/ot7Ym11vVX/oLmlneVkw54m
3qlvF5WezugiPcibqObOCSrKAEb805UEFS3XDNJF4Y5+H0HhztzLA5puPLe/L8J32+v4LRlGv/qg
a7cbtOFo/OwBKk5qspk/BPC2xtvsTxeFC5y0LgWffCAQ7AdM87qnxvHLg0mPGDO8Km1eX1YnGN86
bZVKH8L5pU+C99uLlyG0zgNHMjnDvel5btttNqn9TkxtRlvvxj1cRvYNdcu8oqfIg3uTVnaJtlgU
k2EMWam0Zhb1jRLSREU5cNJZJTuxbE82VC9qB84ytSPIv+dnWNAI5nM6UonwiJZClGtB5nidFDsQ
BT2XTN2oCyD5kmjCHMgZ1UlgmUmlYmRCPCbqeEiZWD8DWvGM0tHoRbpEFVdTh2GnhukuwD0lxaRe
4OYjbarLnmis4kAUbVQxn7BPLKOwOoPnVWRQJlrXMXV6peYxC4QeEz0ZAtvII7UWF+6qsZOypeUO
bpKwliFT7W8+kLoeL+o5IYslUGPaN2/T9Qm5tcsPhwaTcYHMfx+0TlzG4Rie1EyphWSJ2J80YgMe
CJSyMYJrk+1HdycGMSdKLOAOeX+rsXM7clZyTKIWM3hwxpGR5qky2t5Dn7qgIYuSPFEG8jskiMn5
PgPWpdeJqzfwShWDcNR9Rb+/5EFyZZRWBPavPczFAvqzvAmATc7HDpi47X92qNdogJH9fV7HNFXr
jesjxPYK/OzfNg0pPQPBEyrpPdyKLxs/GMvAa4aDWMhQsyBbYasdnfrAlW7n9hBoM/nQNpe/jVf0
6KrXsODBz6S7UmHEti6CC17IPxBjXoqTPe4KaIJevUiNE2DIgrY3+NOCWgh6ahgWOnzBhwgGyJLi
1tYhtac8cS0nwnx6vGweoapv1jeLwTjkupEqQw4sZrcH+EbbnrIKgMO4aIYPSbQ+nzRSbOvG9gSX
3PanBXpn9PBedKEfCvPOTJQzK7x3A9sCy/mx8V03jzbxm2qa8tBGnc3tcsDlHbtnh3XRZ+ecUMqE
XOhFdH+BLT/rDVSZ7thEesqf4c5hDGJBtG5lbsk4d7A5P2UCjj9DkL7WQUtL7MFLCqToj7Sa9GTd
DGJTutTRkL+hsS8NOZ5SOiGQHTfa7ibb7RSuBuKlMr8Y2AvvdhA8JGG1PnXDmPJoJtelZwu2knG9
3CYV6oeTEHD7t+gWgKjtdwu+WaIp/GJHYoxn9nKxQvH7Wxc301Ah/xRQzjtLQLKBUj4Fb/cLridJ
Ws+QEjyf2M+WipwL5wmJrkEoZ+x1ADi9cBg9/tYo5KxfpkSHPtTdwYssHs0aHiY9++A41JGpsIE7
cRzCBUiY2uxlhV9E1l58et6Gi8r21nDyqwiCZ/+O5xQ3Sp0+O1SUIcFw/ss+QXwZqOI4mGH/71+k
GoiBv8fXLewePYhcUTpH5Nt4nrnLQv1f8sZBzc4lbaQnJEeCPr+Cfw/yeiNWr+jm+TVVHge9lXtB
Pch7bmZ2K/gDxvWRTMlWWN5cN/+nf/hl8Jz86Hdg3qMUvHb4UgVfvCDfW4s5BiXgM+z+9Gon7adQ
wxnUdHA75/R9PAWGXnyOTxmP7Vix16+6IwkEwzZRYjOTnslHD4E5BabdHbWtb4WFbgM9UQnaaOBn
a4hp5gbUKrUT7dpw1/85XLIDX98UTVb+L0ag0layfGi3kK2raFPO9SHDQhe/JHnZGDQ1WPCPTjgj
1VPzm/a/eoIf5jJWhjDJ9T+hjTAbnAqQfqgoC8U820BLslNUkVEoTYNcvHwulIs7gHjIs2BBycJZ
6ND81/iiP085NsAZ9Oe00cSLbPj0J0B4SKUkQ2BGfmUmM13YmdBMGkyfQB7yokCRmnyBTGV1fOfs
/5EQKhbuz6NW34XqZVhMErJO+3BsJikHQsXfPCH2Fbg7Yd9Gq2QCmKH+1QNOc2j3QjavuRoKHZjw
t8gEtoSg22MWgMmB7JUBHuUzJVkKtRsvXkNM46oiBrq0LdqoPYjfUUlrv0LOjaurh0Vzic7sajEt
hW6EIYgCtg8jIpD2tP49o2IFP+/4oev3LeTcCL6lfFe4Aak9SIA/bZ2o1RBRNn2gj5zmoe8eLQPb
a2X+hes4F6Fr0+VKSGscHpJuYXJJWYmzyEuPoLs2khuNHEV25f1OvPnnWZEKCqjajyhNKX0+neZp
b4opZ88oMqXC66rO7rleBL3cHpybHcd2fdzF69HPvpsy88WQMqrG6PGVFbOklDfgqFSd/5iu0Ol1
JQqZmjMN5qUmR65DeTocViyaANnulkVSUcIcYAJjYXolGo89jYGCiDTfNFk0SPHWvDCvMhcVIWfH
KaEKY1EHtj7pV0LoImnPCV+MfPyLsn6Lq8Tizp53aR/vZR/oNQc+Ke5GGRmRIDrAOF/o5XLMGgLz
ZPCcEfDwZCJhQpm/JbpfaPa0kQ7g5bx6fQKx8DFYco71qeZmZ1F9O8EeqE0maYRRShKSu/p7oW55
wKfludhGhknpAeqpw3Zfd0GX+XPptOBBCMCehVz58pXg0GI02RxsxGzvju0dFHPSqW86U7lgH1ZC
gjD4Q1AGASQCVnVwLU/walOrZNJVRCRbPQ/N2cF1tCe9PlD4F9Ed/l3fbYYBqOE6eBlkHPg6psN+
W+q4dfV89ii0MXO2xjLuoWlrQoz8MdDo++vv6VTCcaC+nn72KvuByv6HB3XnBjwJ8Qtfg8JAgbWw
7YBrw6mU12HdPMadfDtC7XcVHXS66KEikCunxFsXtcV0EScicBllQxUEy53b5yQ40S0r9LFdOlHb
Ev+loO0L0+W+LzKewmr7AJcnBxv511nWzSQZV2ZHlsgvkfvwBMICMK3T6iUXtWoe/Z1lrS/+pwE0
pfa8QfV8YV7lx0KhmG7ig640e86cp4AQ2yaAmquR8sJDM51DBAPbUoMvJdGmi9aUBNY9XOtKLlvI
c8n3kpBDvK5VVFgJNG2PJXpmcHjkeuDNepOHkugQqugQsEYaxUe0S5z4TxtkKy+Q/iKnj00X/EK2
xxysnUQmpbyGO6X83jOOS0zzNdfgYCyKeCjnCM0iHdX9j/+UeylTdH3aJtOMum5WlGP8+VN0lMIM
VPuArOrpOOkGKlC+ptPYXCcXxFEkRIVHnDhETLOCx/Sqb7MzuYLR7mnFZQ49SmJ7q+MlTqFSfhQK
sINzQXNBO5VVB787T/NMm8HM4h4g9niyLFDJCXw7Lk/+oRulj9PaVhgQlA3GHx2eOXEIY1wJCRKL
PrBa7I7yliL9vzdPsIbzE6eE+tBxAW4mq+VmQZoQYSlLfbn+HriWUnlOQdY6m1F4VNnjcVrPQwtI
oHdf24FHdYfpwidUQ44GSYR6xtcHh6FCRnYfyhyD4ICXjSmz/JjO1gjJqP/ly9wN3O+hLEajNkub
zhabfRuTOoHJYqpdETSzWV8+d/Ccy6camRbRP/ecga/kyS3Vt6t+LspoGG6TzBPVi3TiZZHFE1wO
YmwD+YjWk3QAptvLMaYGST4lnRR+ShJuQfWsU7dSxPPYe4EH+qiuFCSFxIfM6IyAotYAYIl2lMgb
a80wFdN3oYKPlQR/Al0urMQ8iD523WkHEEvu06M1Ff4iWogrfDpvtLCSEiVLHO55jxPmautEOrj7
nmeQoObVkRj2D7/WwbAIVReYUML3XSjOI4TsCnSLsrp6YOBbxrfMHENVbM71qE7fd4DHNTPALqkt
hZ2lMTwB4WnqDwm1PGUqATVld8cMF3A9EGIqK0m8Jkahgq5KqK1q3aHkwWBvei1BDH1B5YdI6fsE
1oaCnUEqVBmPSXnNaLXE9l/VZn9mtjlu5Iz5nQcb4g++0TTurTGxWVJ0lLbRHLTT4C3Qxb+JbeNp
SETYi/XHVDQybBhgmMH6dniU25ev0DgU9GjanDmKRIAyT0dg9SulY9M86nVbXpuPGheohwrK/Jvj
BIjyYPk/i3YJBF4LSgFGXS4Zr+MnsTS0gV0wIQO0HhUlOqo7aqPKFIoY++BL2Y++xJr1BHjOT5Vl
yspQpi8lYwi3lSyGEOrVxTzRbNLEjjMNhRIWagRUlM7J5Y20Sw8xsVMJuVRhtr0EOekAAUOMbnFK
HABplkju1YHMrJXGDJPnLfzgGf8tpc6fJeqbagzk6ssd+sQiKY6gCvPjowjwHXF6sjQ24A8zartR
IuCKwRc0RnP1xqHBl/AFlKPYZo4eMuwwQsRrv31nXwXSot9SIilw0eOdC7NX9oBBczeXo6QCyZBh
d8ryWj8/o6MZWlxNFnMprni/l5ykOI5k5aNrC/P5tJ8wyJN/LbN6bvjNmXRT+DqDIN/FpabrTlyv
VcKQu930J6RzE0sUru3ahomU18/j/VBFu1hsic3vD+Kp7JAZWr/fRJH25LqMaGY6jCWBpASGp5rK
hGycfAax8pHIgZCo5ls20XwGpsn9iLkFVtwYx4CKy6ryWRCJjpFngbszEHOZoRYZRJHeq9jSdNMl
sc9vHHkgsWcTId0SzHwp+frR4V8EdRmIaW3e1DcdR9JhohM/P+qPD6A1Eu0kCuwxcwgBJC4+Y7xX
iyZmquZo8NK/nKCR7Jffa6kW4kR/IeryiiPMnjsDiXZBXk6BLvWUbApE09gBL9ZrDfitYC7Zd8SM
jVgJs1ayDdXc496hsk37InQfwOOy+wPWWGK7Bc9iy3wMp174iEHTw5gAV50mfErNu2fTNo66jNV5
pJhygsu1Z4z918UQrnLjSsdQuc3y39vxXYM/WEezK1iPAF7iONeVrA2L04ACvccP5az67xlsFb2j
FM9anivwR1wMPKmndYm+OK/Zc8n5Lr8w8qGgHT8VHCSijmfHZyetStqhxRB76/L5BB7ydjwEczXI
RrGYpviH52kAKPmFYF8dTzAeaPbmo6juV++/NWBSNP4RTlu2rV8gTl1Cu0YVN/4a2Z24F3dRFP8T
AC/E1cY0ulfMLcUqgFvvCFcQSwbTxkJp+FhvQVGFtEDZ5ravQlBTXGT9YdLoTKPB6WDbxR4AldQ/
Y1kaY97d0+V4BIrP07Tl8h8IVluGv0n14xy7Xd1dffbc30MW/7w2cJWBRrYCHdSCbf+OXkqpvdTS
AquIoy1ywTTN0PVK8fekT/g64wwv8ZcXM7O+noEK2NPceNReSK6AGPMDPtwZ8a8Tlkil/mX97dEr
pbDgtVNcb4/DHye6r0XEjqyP1StFFhP+uv8yOPCXOb67+nu+/J8zIlvLn/Mqdl2AL0jWD6uJqtXg
IlwuPPb5MMzmbblN7K/uWvkCfgkRAnOlnX+ZA5LE3xEAdhw+s6VlfQyvUEXDMvD7Gd9tS20pjfgi
H5NPuWzLXqFyUxMWMUQ/8haKWF2YnukoIX6GW/0bg6yi/uIAtnHPDg8jUIcBHNGwRNsE+nJBEl7i
0+cJL6OS98oMRhboIoo4JKj02ICs5GMoG/EOc4SCoQN16nXFFcUxgOvTLyK2MlsJzaZLgrbxtC6T
Kmexp4++04sCqedfFzslJ5qGs9u2Bg2DVEDNd13o8NN4LK5wLT1RR9T9j/DOU7/n1cB3dR5AD15l
tdN0OuDXP5q8l6bAaay2n1mOG707+U2gOql6YNaoa9E+oXEMy4NWZfWpmHUSaPh6D2dQiqBBVwIu
jKqqzSvgfPJO4xiTQZdwnk1+e4F2xbDNwNt6q+Z5QjUIsd7+0M7h7ekET2fAYFEh2A5ZE15X90H4
/iOyW0XOcAUMT9rD52nRj/6HqNA4D1w9zDISLvAg1NpPKJk46jY0jjLew1BFdNG7uArO2bg7A8qS
WkCMbdHTtgb3JHYwOggQP/jClSsEKOL+MlJ4Prp08teSRbsIlHJKNklUVYz6N4ns4+fCMr6ninxf
YfRlnp1zUuA5PKQ04DYy7GU03jqCUVATVQYwRSO5yNLdCtKCzqeJ+v/fUlvYHOxLaErXuSoUU5Er
7fqLmgsYWkLaNUYnuPayWq3Vv8H7f7LUDellsAkNq33FZGRcPMUSCO8oNdkqZp7UiihregfnmC6l
RRvWHgDrx2JWqLGMR5ops6BVX6IQuCDyFxcLX8GSgWBkp8lqyScYpPn6ar5yMkzVb6PedjoTyvJC
+6n0jN2/092XwAw07JDcpOtD6tekMMwjCdvb0g0zfPm4CtUpXCg7dyecZcP4o3yVPpEAUlJkMoiH
bxMc1H9qJfVR7hySP5vwqzYAY+QWrL7Svgzn0BvzlTtzkL61hvt0/AR7CKhknzbNxgeik9fu0WHS
uJdNQTCqMeW0ZI6QqK23Npga/qI3NzKTn4ctmKYF9Ad6KuOMo+Iul9tt9cQDJNvJNHKp0ohQtx7Y
VTii3vKE4DwWaLcLpROckbI6zlaEhVfdSmWnBhmtkIfuttWSG010/aZ5/mdXkdjC56xVE/g7RkDA
8H+ZdFAtgMMCPbegT9elLk6+AleW6o+INngkIl3Pv8pmt+nfXkvbLbFzWzOK3RMRG6TxWru6uc1o
nKrncHfWUR8lu/FDk5rJPmNzAqnK2Xz5o9WwMOP++ycVldqbO1xyub+ThxhVFgGyAbosQsCMlswc
REErW05foeE32U7Foqr2qLec3wrHXS8OhYGfE6GajbZuN595h+iDoiiE+EJGoZmfUtDQvsrKSmig
FG8r8ZZTJPm4YN19dwGCmwjDO1tkpNlnv6sapHv5MJlaG/yr1aeuhXxGkUistBjgObCDKbPMW71p
AjLThaDFbKJUuLUmg9rXpdZ3dO02r1nq0SKV7bMTpzVqHiqpaAdubBWZ7EncA5HaP/SsaStkMeNI
30MmfRW8SWFp63yNp4tfPWr1PfhO0wRYzo7OKYMMAUBWT55krO5nC3Xd1d4PWKeU/ZDoBkuwY0qz
XdV7RHaUhRlfWg/NY4e5O6Szt93TJL9AcHlro/bqAqbLpK2JpAyduhhLeHVC2Ir4lEdLDsjOJ6p/
qoyPrx4Zl7pDL6/Zh9W0g6N6tvCGKFG4lzw9LjTlFX6rP84NixQ/5lhOPB1GK3fBLGGQNNONVGzk
EP9hSpCZtDWci/23T3WAsfBijljjRpbQOzmTtq6K20QyjPUuZBdjSIZUobkvrEaqvkk4vwOWoTK+
zrmDYRarNK4v0rvL6pvou45/SEdaqcOPn3ljjQ9zPt0qvfpS6djm6yuBQewRkjfj+2y3iGHk4rLJ
CeXjn/P70CLKDNjTKzjkU2i8awRhsqUogd+tMpa3zDIzVCA/dr5SHA9RZUtYF9hwpXftGnlPI8DC
du9wvYFot2bDQMMPJ0cUGZo8OPY6v4bxmFlkR7VxJI+Ef99D11NLShvfYYhbf5kWxpggU8VLTApA
5PqwD8BFr5BZHfGSkDQxQnjyYBwQhAnn/BxYQL7/PNaTxzCaiEMUtzMRCpSd7bfjqNoqcHBZitU9
EnFesvALiCBSO+s9259N/iqd5FEcmfj+xuflfOKFQy+ylpBv5FND/g6lUARpWJeRW04CPYgynF5P
Fmkz97Tw66WCT7DE4/MsuOzYYqUTqPGDeTVYraEicrz3WsZCYO6iVklazWAOiyw9O9KkTj1ZBz9w
nx+ihAr3Ingk0gXRLEKmx/LSl8o9ZXCMrE3ciaHB0l8rhIyRccJaNkx6jN40EXQ5BrfjVvi8sSij
aJ+S7p6rrNZ4EYdOWthAmbu8NQW8gzQ1tLScK+YbJ1oS0uEy08C8MRQMr+qJilvmqSVdq/J9DHZy
J6EeD76c4DO03AZwI6kzUX7SQ2MBP5RUuvcgsybUGfM4PbQrGPS6CzSyug8lRMjotT0MgF3T+x16
hZMvqQLVuYAOWz5jGA2+a26HpT7CiS1AokmVdZlGU0X0cse60ADXNO6ADVo58HKB1SawOg64DL/Q
EffhMczWFJvNyxrXJMMi5rUo63v35YMpmwpypJ13H5nfQrdMpQ5FppmT9lgQ7urfSpcPiFoNpVje
WjTazxp+TfK/W63/lCyDwE8nZYBrp4pEC91GvNdgVHqo983HUTGq1SsCtBkJ4wXUdLsI5GG9VTT5
H8T7oKllpMtb4zfjZYyGUxtHclWhru8lFOGmK8li+ZlfabHB/BHMtwt6G+H0Sf1Veofk3tNPm9bR
mp5f3TzNYHaydFR/NWA+BdkCVolYnebjMl+5CuAYWVdRjYDNIBheG5Bg+vOTbobknhxCF7DtR2uf
LlrYd5wAjz3tJR0pXQZ25F0kNIWNp41zmpXAv3woR9jMhTSXJDzkrJqze17r2xzvAhRqjVCJYD5C
WQhEE9PfCMDWI6t1QNfOs1aeHVMHjHLVw9fNKtpDcwpSwU7kAP1o/GyNk5ugw5e3gmVLNLZSyEd9
CyJbCC+XwnpIaN+QnSndyUS3yeCJ2NdRPhmp76x6gLMYaBxzMxO/wF5oEcj4RBmfUvsEXa0fikMT
z840XgpPxQy05KHr1O83vx2acup/KzKofxxpL5fcwRoF2EoOdEVzGCQUEUwB9mozl97LQAKr+MQl
7Lbsi0vBMpZMef31dbDLaBLD2/4wSKdgEtJ4Wf9Go3ihfa3zXQoxvoCUlWyHy4+0c+ZuRmx6UpRz
Ini0IU3zLICDc6S4e/rRcW2HXhgYo+UlYvbf1g6hbEizsUl+j/cmHU8nD458byjSKZH+dMUV+fb1
OyaiUgFjGU4KlurY4Ov8VR63tWtgRo1jWBvQuQ4hALk9Z97gToDcUT/Lguvfy6MBCxKjqRQnzljO
noYjsNWHMBWibZiOqblAJ5Ij21SPFRq1cDUxcyosj7akCdojZK49XLYMUPCuw7W4Hwkd7ES7XTgV
ez5gDgrmHuKfMeKnIaUquOMqiaVhJACCEct5/OWsJGnqImCHH15Vw2cHVjOnjqvIhpooL4KrK3j5
3p70FPASTx8jIoxANEgM3aDC7QTGPusMBeU72/FGYVUk0S+gCW1lcgWlWgRbWkOqYaaunERF0tk4
vRudjlkHhzx/VEWy+I4Vcf5gUg+CpxBuwhHC5PPo4g62z+Jlf7nnZOtiKnifMdBb3Zlce5hO3gKz
6T2S67qTa10e8FjZNMVzxeYEfA3cuEUJLLrZ4VRqjRXQKYOtmOi98Cc1JVs/m9wKGsVpSaG7VPKW
7M+Ltw2RFulnHCtWM65zYdXS8PXQaP3WuBheeiVAFxWxMGa9yylspZ0BdCXdQ2jcOZ6+yKR+cpkj
TnYwPDcLVSTmEVDzsl7yXoKL8ASY4NCYFknjlLmaa97hij0vDrQ8umuaDH/I7Oj22IzLBTYBqcPN
pJsGoPHvBaRlXAG7GJarhG06C21aj18+iE7A97k7Xluk9FBn4jOHJnuvliK+BXa9rLdrKaQO0il1
+pe76jn2tETt5zC0PuR+dQxhr42ZTrygaPTrBZQMlGDcj9aX1qbJ6cuH3I44sv7eaSqMd0o1Rqqd
WkgzNQTEzyMQlpkB6/t70QI9X2UHyaELBphZthh86utuWC8Mph4/YyxdTSrPffbD/NhQVQ+LNMue
UdayU8mO9ijWJi9fVKK8Xjk3GIoiTdWJZAGfgtbAORx46ZohnOCWQyQGUTVLbvroK1MIygPeb4ZM
VViB79Gt+ujqecJlX7+H6YaomHKdwjEVtpX/nv5G13Rxw3/AJBGAQ6Ki31tmtRN5ubI9cXgZLXmC
Ylc22hPGjvLu+lYrB9cKErwbKnlH2W3dVjHyUs7KjKcDsJwavbfBuxXRTr6gcYjCsOpc9kQ2/5/c
OE5O5K2KaE6UyhKdmvFxRrSsG+Df1XDeWeoTBMZuow6EK7M8haek993iOygkn1epq/9UkfuOaADQ
N6jyYwTdRyiYvik3AaTT6+LgR17bfvlFBjmowAW2yBWOi/8+0ncE8DssLXVAcsrGj9EWlLMRmZ6T
mSSrf3vYFkelh5vyh6nB+61xCT1Lq+JrikP7JJW3/3ZE8gviq+jlR4pyBrcE9FmxSI0dJyPGx5w1
uP4tMvR/ccnL22acobjShUjMz/h9S6KIpk5zHbsoo9EbKiDcX7wR+l131rKf/zlT/JPvVoR6xy0g
3FgZKbKtNPPyNpzhKRBlPJrAfwLU95vAYpV7tFq5ofemMS/39RpWQTaJ4c4eSzDcK1JtJr4xZlIx
TVeaocxIhfs25yNvhua4hHnkBeFi/bCIPzsm5yPfRsa9l+B9HmTx9o9VZ5RoutJ70Ln+EK3WVEuA
Zn7JMjYWEwBNj2BGEEWxG0kNIctuR+ElquC/uOHi9l5xGyiA+3+Qi9mowApB9i9dU8OIjhoAlA3d
rYGw3l7XRef8+SqHaYckdW0dVORu2Mgv/ykRKTVgGrFn9Zb1sy68FaF5H1ikSQJzm7362FLXXtRZ
IR22wWDh5VIU5egddUtHBjY0anKn9LGQcizoc3OrK+9O0RIJVLGYr9WMDNVcp8NEjvQLWCEE4B9j
qzOaPCIXLKoUDnavfMENMsJoKTi8gzZzYsVkSkFbhPXFSTIq236rzEWeXTCraTS+Cir2UJaG5cUQ
rUmve1j4t7gbiz/NA8NO9nMYLQlNGCXlrs45e6/Ywrle8e5tfDZOLWbECsR46R82cUcuHUvNwOXd
FxQj3N1/46/IDFZz7uy4EQhkwChnmuzDtJ548QPpNEC9WN2XAlveAhN+NNLleg7Tdn11akpd55+G
+43gk/Y16QQ7UiuI9yJ1uR3+H5+IdBazHwrDAvulLrKjn4fa0EO0UZe00iGFluoiq/BMB6Kz0dSN
17EAsA7AjLKeOlTroshxZ34paoSdOseZRQEkcI2i+s9rNPwKYOrnNzB9Jjmu6+t+eWYp1nzIBVmJ
vDgxgg1s1Kv8hdGKJJvZQQidNFnI6rcOvUsnIG0cITawlW+9Zct1o8C5kizBdP+38lgKyPOcxA69
CuPK9BsfnnEh6kUttxMA2DdZQuNsM+Lf2EPnL9sd4xNwPj02Cp1xTf42GG2V/d1/gDeBN+rT2ku4
wiFxF86VOdeWLUgrJ8xLkKPAWnZvgeO7+RhGBAfNyfJpJ94lOlYYNr7t51hDo7euVpADMWU98K3y
jda1Yj/5L7pHdwBR9YEAi+R3V7R2FNkjicYPXvZeGWCnxNUZGhPKunjb28gU/RnqeDWCgHtjeHZo
ghOQoTGIFMb4Fgv5dp0kMJfOVddFS42vM2ISv98rey2wOsQxjTuxzcEY+Haz4m4tPw4kREkropqc
Ym3Zk21g86xKHccA842Wme5mEmiDx0aFezWGc1bIMxX8MQD+AExQBdSbTujMs3CT4yd5Pt5Isk1W
hIYCjGsFD52k2XJB7svwrq0zzDqS8FA71IfDjiIvJ6DXvOsvxzhzP50CKCfjWhgKYcsBrggn/Os/
LZNgHUj04g6q3ow8Vm3QBgomVjhqdj/JfGj5LDHyXCjU0RxuIbVJ0EPXpDy0AaJ54jINlqTVPIJm
pMRhDLXCO29QPXgFusj4c4jf1cqN/mrZzihQcGJ0DjGIMTcED7Ym1wdEr23tS674yM/FohtnsXjm
Aq7GIs96857kPISglcXsWvl18YgZBSNhVee9/JHKMkggsdpij1Z/HNqH0xhBHQBj+Po8MPpe4Mt6
6Cr3R8lUonQtHdjzWI25xY9hyPf9Yb9lVY1rom8/2GYTRmaKy7g85rkHl2Hzbz28nqb0iZ24ny+Z
T22ZQPU9CjjmJvBkIAUkMoVEsiouz2JM9tALsoIhb3UEgyKYoppHHBbK9+tel+SRaq2o9vd+IAoq
WevYMD+AlpDwuSiel7zcNKxg2qbL7FCNPpPp+YXEB+P6cFVLFyZkz7EaekUGVHnJcbTxLxBdGd5u
qTrhdijTf+KuSgS7I71WLIQqKm1oI6/U1Sb5T4he5w0bvnL/3xvIuo4Zc8mTgJx/frVSvXCI42Cg
M0HrNNAumEcdHkukTnnsX4TMFOXrZ2oK2uj/zrBvkcNQ8KUVbAviFCfz+dJljQ56Yn0Tu/CflNLN
C9HinrdzUPjM5wDZCPWg1I6Is8nEN8HB1KYtf+ft/W3uQOB2MInGeWkpZc6Xo/BJniuceqjY6iWO
zhvkClYr4zhl/QzT5OfLTnYgVtX4cYZH1wElL77T/PXz49XTmE3jQflk2MPLWnYVUcTnULNLqC+6
cYFaOihsvNZy1TUoSX3QnhvpqcyuaKPTPwf13v8uHHdpBcgmHOkUSkri+TuuDr0yaN4fWdIdeMzG
kJYqvBJKhHjCRPqHOOQsC1YUxFVqodTkNb2KJasRLg/oN0qUB2NDfkeNmJpqQtC06Ffe+fK72Qu2
XlWUjCUvpUam0YO6UPVzU2YXI5U6JwdXqdVm/jFQZiAWjnl4v0cmGoAytIDmZdqCl+fPLVLTYbav
JxXQXV2C5AV0JQRTHFHl9k5vrw3Jl1jVZiQzOo2taGzasuqW4dHqZk3bi4tqm30b1aDDCW9n8N6x
QKlj7ZDAzGSLp8xMwXmCn6xN0GKrT/8XNxzvYSKGg7NHk/kFjRFDhepjAB4RG9Tp8zTRxQ10MIjL
TezEwXxsRp9uEg9fbNHVCQ0RypY2exCYQ4Tv46hkvnrafZ+x+8vK+NC3gDgsiPSqBTd80cq11OdT
JzbIIbnuoQCANmJ3yN0pHAdyEUFfBu1J0M6y2gkQeXcc0g82RCPTTYhe74a3DFVwlvDAx7NALUhr
OIqNrkUfFaT+FHZXnNPb7j9hRauaZjdAdlvTTRYJxU95S3FHPmBVnAtztUi8yOuIz0Vd7I+X2CqK
xxebeJPgT9BQT5yWJqjE8lCXSZSsU3hFGnKAOZ5i5oG89vsT9UirSK8xPT1bsxZ3mwapvoS1qvDB
7nrPO1MM2NwhZfsrTE5RmHn/r3arZ/cPyg+Ss7Omr5betM+dmm5M1mBbMm7XYMN49V6qDmdj4PJm
sFe+fGIqv3367Oa46HAn+soeHOiUFprBcBuszlvIdlM8gQSs6e4Ue+nbdJ6cYzYg5DumhnOUM0MO
W5cAbx3cAxjBCZOZ2Aa/iKB7uJw/2fS8TYG5tblXb/Y3++fBPYTsTCd2PJOUOvFM6xKNvzBBgV2E
jtNxZXRebI34ERQPctp72QtsB4il2wRK7YpOooovCFh1hvX8clYupC5kdVgnJ4uL9SJUWS890KtX
tuUR7KvLAqmVrP8sqRVYv/Y1gp6MkAJzQWhRJaWU4gG9zjz7e3Kck7K8x0MBkqG/Bl1BjVMGf1Pi
7kgKiaJIwF2/VZT4OUXxxAcrn/nFUxotIgI3jOaugYlX4Fnwb6pPJRmQWn+veDTnzZhxP3nEauAR
r1J/lPocl5WNTLlPJ7ljGQ823CaPMo3rwvA1a3r++FKiLst5ZltFkuTh3gvqV9FWIcHv9a3235Zx
za5Mc6YJc6c2Om+4pqgrEvsZUM3wo36mq8op9KqoSSymwHpEtzTdvncLP6/CHbRaMcWYusmCxZaB
ZDKp50oGYRUI9wf8+9nEL6slwxMG7jV2Ut8KLLWt1Lcy6LI7GdKD3CuL1YILF2j7W3xCfF5p/86h
qeMQVmHup1eIkMogaPOP1Is7JMMYVQQro97y2H6tnjEVvuBWwwFIX1JVOAJMnoPY0zURBmQFUQoM
EWYR7lzWB6MznzOXgJWeOCJGbA4fTwLXVE5XugipD+ACkHFKUCglZW6hl/JZgYOubxB9Pc92phUg
8MEbWQdHzT9JwFto9OjmqJaC2suTS/tYg/xnVuI1HlYctnVKIc9qS+braTOkFyX8ht37KwELsqIS
tsd3XW9eqp9oRYFZ9+GPc8gwXXEK5n74X/2hhpYkWRbtBg6/1OYIFb11DVXzl8zNdRfCqoFUJYQh
Ron3OCdxOzRxCEPcaiTKnM2gAnqENxyAIAMdYu+pAk5l999/nYrmwQf49MIjEpNhHUhmautTB/tF
lGT9ek4gyvbKV62UXzoCYA0UVrZZvcAtIf0TmdQKJ2y3LgvLhd44+1a4U2fKkPzudmBhls76Q6zS
Yz4f4gzQrvDXox4+2bgPoE79uWL0Ev0My/AC3YegIWJBM1qrZbKEu7BOEjYd0rI/qQWRskqX0/g+
s+fLqQKiLH8NgGCwlpMLDLxCBaSxUr+P+fZr2BEhjUCLRl54eHzzJZF/3+G8zQKR20CptTQktXlu
hck03CHwXKBhSEEZfPawoaWRYb1Fblp0Ir45Na14pvyQgww30js+m4APUo1yzG8juXYJrfbKzVet
4cvied3WvswROlsDUoEn3Ui84SqvQONqw8sPHkX4YUNYZ/PODQxEyMdWKt+FxFAb55X6YZZwBkLJ
nVhq5CDOXe2Al3Bk5yJhnNOLDCqtLSLB/qxkAP1xYZLAGkfKn9pP9F/fCOvKXQ22u918vLZkF7Yi
sVTvxwTDQIz11virhoPytXmHUCvcMLNI8D/Dig93ZUhHydRQ6UVmxpDBx73EafVbm1asgWoPQ9y1
jDx3No9RTbb9ut2S/1tT/Im02cl5ZL7HxaoR2sL4+fyQySvmgRC0yjJW38EKZbRMAuacU+ARY3Mt
G5XhbH15ZoANdpf18z7yCXqmqEoyD045c13RnDQ80CH8bSTUC+zr0hvqPurhGrMsUoIsZtxlwEIV
Ap4N1NlNmdGdLIwb/5kXmjtUlsBrXHCGoisM58kUOu8CiTpZ35VnGfrhq6nfCgXNwAuJBdKx9OSy
UFkPk7npLEwHpEMbeDMUorjdaFQc18HneDN5K9dwgju9S8cSYljyZOwvQ9LItDZsa6Au/Ps4pZ9G
kpl7qQrNY6kjdWPTLVq4EU4gtmEcWYUHUUPeCZyl5mVoLGbZeLH0L6W0daCu8Ngi78MbWCY9lFXU
sx00QqgfL9o5x692tUnvqMuNpWN68oeEMoVSDgtgG24HTdZo3fFy1SZldAafKxyHt5adOBrJwJPl
Apj1VV+dD7oxu3/hjPX1dlcp9fBmId3dlaPekCTObAkjTWRMl/Lcua2zODzw512n1YGqdCMQV1wi
n3B2q/fqo7C+7RAW8zYKOTjEIAi182q5w7gKA2bc5ChbDtiR+oqfZhVF9EphCJZzfszoQQCaiyXu
aXEYTixtuZpyNywYtt11GUYDMTvTX+/EK9DIVWvvXSnbcZo6+SPKNrFlKZF+K4BnYSW0luO91gVn
V5fWshjdN/9gKtlF6CPfPIpZWN87f0gqMDQU8PqnqrnHlEe6qwM+pXRa7Y+rDg8OEpcOzSUDuYod
qLZUFzJNUFpA3GHhBrAJ8XBoiUcn1cMEaqbyQ45EL83Kisqs3Rieq6Q3Ubl9f/g2rgMY96u74U/E
PbqObyALotSxHfHk7G5J1+LM71sb4KxDHsTq7HPaJ1PoIUA/gQSgTNj0KUE8W7qRtwaEs+8ByGsv
AqtbVR22hl15+cOqk4oaYAqQo9WhDpg0CwootDyRXpCu29yj7Oc8git+awaP7mthcEj1PR4YQxX1
HU5VTpP/ENIp+b6WOx3B737EUiWnQGHRzD0Zq2G863iM673E+vhGUZd5KSagBvSGq7CettI5frLh
QaBDG3PwWLNN0BZ6kH64QAENbiE4S+h6WmYaZ/YGgVkG8Y6h87tV6Xf4oZiFF41J8IaqryE+SIEj
/LeIdgMTf8Iz232YEo95lqkAJvUiUhT4VprTNQJq0Qn1hzIuU5jGcEkkZ5u/r7d/oLyEFHj2f/7+
K23zB9W/ysOzCYGcGCcIGazn9Q1WpJxgEK0bCNSqwheLj29mG15OEK8qQz4H8oxBfb2ibL7pSNIM
DZmEYSDejmlxFmQG1RvJSqbAa/+ftjtFybaBnzABKWiygvwsdlyo239KWSscQMb5/ImY73NH5g9Y
bgwy8cRrYLMOEYDI43bB80cNww8UvlQEpwQeMLnZjzfBXMqLWw3v/ndu2QMl1pDYlx0i0HFCqzjW
M+RLiQn3501DyeOqJs6pVXF9+hsWhri6ArJc812kgOjXCcbP7FKtPZHxRPHJFoyQnswyNRYx2KYT
j2T2GyZzF3rxu7Fz2Bpz8xtDY+AYBwoo0F7UjLf8ap2LdMlWK+8jQw/AtnoTjchPIrozi52XA2dL
s+3tzFm1eEpU8MGCDhp9ZvG8DWGv/6FQXwbtZAMiO7Xz7KBkWm/C5F/gmKYR9tERF4lU7zhfmKjM
2IvjELYIQM3OEZZgSxUkhE/Cs2qIlakOVE92V7SeUR9I8l0/Fc8Ac/gRnuzI+LVy/bqbvqtR4GPe
GGaY0T3u4J/XPmhB63cCtUgrpVMXAt35vEdUOxiuOsXri6FuV9zQr7EXCorM9huCNNGzqTQ3T7Jw
DMjArfhjTU3HdIxfswltmbXawSv1GVPNj4ALCD30hhnKPN7Jg3mf+kyz8f2h+g9g6QxVy03c++dL
7RD4FmIVvVFxm7aNU0pWA6FIhn1CMPmQjyniAkNscU8WH4giem4KLV+k2kgNJK8sijBbR2bFaCvC
i2hAM4B0+r2hX1frDG5Vb58O9leFtNBKn98npf/13lms+JsmDtrK7sr3anNGKgHoaDkXkgezwkZp
++rD8h2iK3JzZFjRAG6VnyagKIeFSNIIAPNtblshis7o5xT+cUWBNul7vXEYzcyV8nPzXttUm45o
0IA8wQuVcp/czASLYykzJBygbZHPSqGLSY4zR4cHJr5/6U+fAHxwNt+V2di5DkqvPAENVEBG4shO
5t1E/BW4Rz6fYrx9kwEncSN/MOeN9aZdMZ8y/3erV+lGs6dFBXLmF/NRJaeU1dwxPcOvZhXRC4r/
rzk4OXIHuuuplUzORvMBXGNUQ+FUYYnkf68AsXrjnJ/sPy3fMGuWNsSL7pwgWS75c/GMhld7Qxc+
smTkoX5LN0PZrH4lU40o9FmP027AR1SkE2b6sRugZUvQMWs/nU3K2DqzrVR+UVY2cnnw9iBDNUrp
OIjszCuFtHOxxi7FmCFJAmaj80LXoGNAl22zVhPdqBTx8TL/5F7Qj0rU5ZSlKMaDToiq9+dx8ebX
dBJRUR/n+hUN5p+2blflXiGy6D4gmcL9+aDjCJjnCTCNCgKoFQYqWmGBUviCXI92GpIN1yrI3ahx
e7IggoU9ULyd6RMvBnOxo2nphkCzl3ypON0qEFB0ImBnG9yvdsZOJrR/Fa/ugDVoFCfBiaCltW/5
WLHU2fRxuEikXcDIQ0blPZ6fUqTZXVqrnNdNDj66w3e7Y8uKIJ/TelqkXeVq1794shqivDSKc1tV
SfXPOWcJLX28jeyZUtIoWlVwYIBD4J/SzqwXKPr9wtinDaub0j7Z8iqNtRIStZdTnAS2E0FANVhk
EJCPC2SCkZnZe6ENiOa69s4Th3X1wnJ3iM8Pu2FJc6agsR58CVN2OX/+IEFTA49cy3isZwiy1Srr
lBzO2J1HUJxOTLgu5QfiX4vQR4OrrZIffhcUl3DvfKuyij8PETsZNrfRdH9QyexOHdsopCk7/wZt
cjQxxS68m+oX1US/xT4JaINVo8KzTUAgA36/ABlHhmFsrblDtfG36aq9N1K4U+zZgkQ43YtV60pM
T5fj8byk/CDJHoAkl8vuZpDrLHxWZHP3vrbTuSbCXKbV9xjY/qFhMpROwK1lW3z/7yrfViTP1tyb
umEUKH8VaPyodsg5afiqwOdHjlS33Q8tq7el1/QCiMsLpNCy8N6MusfP5AzHt9gIK6Z6I3YAfpmK
JboRmnRaFumkYtDKDGfr6MBrIsJIBh30T3wkIOJGT7Q33eIfSVflCUTHdLBQo22k7WqlrgWT8Lw8
NLwKwhTL8nZVKZ+HkiuHuEcpIujrWnuJvu9DSEIdA03omQ0vlaHs+w/WNW4YLbKLO2Zj7aptWmYY
N0SyGBpxs0uTEDojrb6ICWJc2G5XivhMmAzkjqEEXKRhJRFH+PI7b1gYCsJRI176bODh9ixmP1hj
SmzsSP6KdwCQPtVlCx8xw/u64YZ88eLR81emkeBcn/KiqtygOqwAU8Jtv+pYgQaga6whbDwgt2iz
RM0LOXDq4S9JscB2qZkZpOY0qKVhWbZjlZ9JspxtBmS/Ce+xImQ8kDOx/W2O6RBK53BgCJBuw9ER
H6L85m+J9trU8+xAfbzcVdIUe+wL81FEQJGLZHGlioWMdYsCVeJ1SAWw7sL9kdQFP3HKUzLDP/xT
l60OcCsTzOhENJdOFCfZUO5cDdXbRsaCF0fQdZI+QBf1TM2BMYUXLjqruatKiSnKNWzaQfYhIEDm
0W36qMpr1OsTNN+VPQAmJjhXOMlRU+3nifYowEw8vzJhhsvYIlEHXZLm2jJFh4x5WHhvbLqhYIzq
q5TrEKRzI4Mg49bUxDQyejg0BeeBrT9sAg6dFMYwsu4wFbHpNl9OtfzgEbhkrzJs4YrvQMAsM66S
Aps9ZCYRrkWu9hceZKMJTGURxrmT0DI95tGFMHNOk4O+3t5VTH03+vqdVju593qynYQIinUEI2ka
AAa6X0Ar0QJfMpSGCx8Ve0tlwsOSPMafRD66eMctYIJ0N31yQOyrc2PegA/1PJNFi4o6XOREQhhS
YuxRtzHl77zdTJbx2vfcmhZ7tPLqNF/Gf5TWjy4qiMedxR7uhE1GeA/F8eh1iVpNQFH8X3V2CZJD
GGcra92/FspgZ16JhXcDdF61N5xP05HbtGcGprlhB1teF6UCa7aJXIsNDLHmJNU=
`protect end_protected

