-------------------------------------------------------------------------------
--                   PROPRIETARY NOTICE
-------------------------------------------------------------------------------
-- (c) Copyright 2014 Semco All rights reserved.
--
-- This file contains Semco proprietary information. It is the
-- property of Semco and shall not be used, disclosed to others or
-- reproduced without the express written consent of Semco,
-- including, but without limitation, it is not to be used in the creation,
-- manufacture, development, or derivation of any designs, or configuration.
--
-------------------------------------------------------------------------------
--
-- Company:     Semco
--
-- Module Name: DigitalCombiner_tb.vhd
-- Description:
--
-- Dependencies: Top level module
--
-------------------------------------------------------------------------------
--                                DETAILS
-------------------------------------------------------------------------------
--
-------------------------------------------------------------------------------
--                                HISTORY
-------------------------------------------------------------------------------
-- 4/17/15 Initial release FZ
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.fixed_pkg.all;

entity DigitalCombiner_tb is
end DigitalCombiner_tb;

architecture rtl of DigitalCombiner_tb is

  -- Define Components
   component DC_DemodTop IS
   GENERIC (
      PORTS       : natural := 5
      );
      PORT(
         adc0_overflow,
         adc0Clk,
         MonOvf,
         MonClk,
         BS_Ovf,
         BS_Clk,
         amAdcDataIn,
         spiCSn,
         spiDataOut,
         spiClk,
         pll0_OUT1,
         pll1_OUT1,
         FPGA_ID0,
         FPGA_ID1,
         BS_PllOut         : IN std_logic;
         PrevDataIO_p,
         PrevDataIO_n,
         NextDataIO_p,
         NextDataIO_n      : OUT std_logic_vector(PORTS-1 downto 0);
         NextClkIO_p,
         NextClkIO_n,
         PrevClkIO_p,
         PrevClkIO_n       : OUT std_logic;
         adc0,
         MonData,
         BS_Data           : IN  std_logic_vector(13 downto 0);
         video0InSelect,
         video1InSelect,
         video1OutSelect,
         video0OutSelect   : OUT std_logic_vector(1 downto 0);
         VidSel            : OUT std_logic_vector(2 downto 0);
         dac0_d,
         dac1_d            : OUT std_logic_vector(13 downto 0);
         ADC_Sync,
         ADC_SDIO,
         ADC_SClk,
         ADC_CS_n,
         ADC_OE_n,
         adc01_powerDown,
         BS_ADC_LowZ,
         BS_ADC_PwrDn,
         BS_ADC_SE,
         BS_ADC_SClk,
         BS_ADC_CS_n,
         BS_ADC_SDIO,
         BS_RefPll,
         BS_DAC_Sel_n,
         BS_DAC_SClk,
         BS_DAC_MOSI,
         amAdcClk,
         amAdcCSn,
         spiDataIn,
         lockLed0n,
         lockLed1n,
         Sw50_Ohm,
         pll0_REF,
         pll1_REF,
         ch0ClkOut,
         ch0DataOut,
         ch1ClkOut,
         ch1DataOut,
         ch2ClkOut,
         ch2DataOut,
         ch3ClkOut,
         ch3DataOut,
         DQM,
         sdiOut,
         amDacCSn,
         amDacClk,
         amDacDataOut,
         dac0_clk,
         dac1_clk,
         dac_rst,
         dac0_nCs,
         dac1_nCs,
         dac_sclk,
         dac_sdio          : OUT std_logic;
         BS_I2C_SCl,
         BS_I2C_SDa        : INOUT std_logic
      );
   END component DC_DemodTop;

   component DC_CombinerTop IS
      GENERIC (
         PORTS       : natural := 5
      );
      PORT(
         adc0_overflow,
         adc0Clk,
         MonOvf,
         MonClk,
         BS_Ovf,
         BS_Clk,
         amAdcDataIn,
         spiCSn,
         spiDataOut,
         spiClk,
         pll0_OUT1,
         pll1_OUT1,
         FPGA_ID0,
         FPGA_ID1,
         BS_PllOut         : IN std_logic;
         PrevDataIO_p,
         PrevDataIO_n,
         NextDataIO_p,
         NextDataIO_n      : IN std_logic_vector(PORTS-1 downto 0);
         NextClkIO_p,
         NextClkIO_n,
         PrevClkIO_p,
         PrevClkIO_n       : IN std_logic;
         adc0,
         MonData,
         BS_Data           : IN  std_logic_vector(13 downto 0);

         video0InSelect,
         video1InSelect,
         video1OutSelect,
         video0OutSelect   : OUT std_logic_vector(1 downto 0);
         VidSel            : OUT std_logic_vector(2 downto 0);
         dac0_d,
         dac1_d            : OUT std_logic_vector(13 downto 0);
         BS_I2C_SCl,
         BS_I2C_SDa        : INOUT std_logic;

         ADC_Sync,
         ADC_SDIO,
         ADC_SClk,
         ADC_CS_n,
         ADC_OE_n,
         adc01_powerDown,
         BS_ADC_LowZ,
         BS_ADC_PwrDn,
         BS_ADC_SE,
         BS_ADC_SClk,
         BS_ADC_CS_n,
         BS_ADC_SDIO,
         BS_RefPll,
         BS_DAC_Sel_n,
         BS_DAC_SClk,
         BS_DAC_MOSI,
         amAdcClk,
         amAdcCSn,
         spiDataIn,
         lockLed0n,
         lockLed1n,
         Sw50_Ohm,
         pll0_REF,
         pll1_REF,
         ch0ClkOut,
         ch0DataOut,
         ch1ClkOut,
         ch1DataOut,
         ch2ClkOut,
         ch2DataOut,
         ch3ClkOut,
         ch3DataOut,
         DQM,
         sdiOut,
         amDacCSn,
         amDacClk,
         amDacDataOut,
         dac0_clk,
         dac1_clk,
         dac_rst,
         dac0_nCs,
         dac1_nCs,
         dac_sclk,
         dac_sdio        : OUT std_logic
      );
   END component DC_CombinerTop;

   component LogToLin IS
      GENERIC(
         LEFT_IN   : natural := 6;
         RIGHT_IN  : natural := 4;
         LEFT_OUT  : natural := 6;
         RIGHT_OUT : natural := 4;
         LOG_RATIO : real    := 20.0
      );
      PORT(
         clk            : IN  std_logic;
         reset          : IN  std_logic;
         ce             : IN  std_logic;
         LogIn          : IN  sfixed(LEFT_IN downto -RIGHT_IN);
         LinearOut      : OUT ufixed(LEFT_OUT downto -RIGHT_OUT)
      );
   END component LogToLin;

   TYPE vector_of_slvs     IS ARRAY (NATURAL RANGE <>) OF std_logic_vector;
   constant PORTS       : integer := 5;
   constant CH1DELAY    : time := 800 ps;
   constant CH2DELAY    : time := 500 ps;

   signal   clk,
            reset,
            XX             : std_logic := '1';
   signal   Dac0,
            Dac1           : std_logic_vector(13 downto 0);
   signal   ChPrevDataIO_p,
            ChPrevDataIO_n,
            ChNextDataIO_p,
            ChNextDataIO_n,
            PcbDelayIn1_p,
            PcbDelayIn1_n,
            PcbDelayIn2_p,
            PcbDelayIn2_n,
            CmbDataIn1_p,
            CmbDataIn1_n,
            CmbDataIn2_p,
            CmbDataIn2_n      : std_logic_vector(PORTS-1 downto 0);
   signal   CmbClkIn1_p,
            CmbClkIn1_n,
            CmbClkIn2_p,
            CmbClkIn2_n,
            PrevClkIO_p,
            PrevClkIO_n,
            NextClkIO_p,
            NextClkIO_n       : std_logic;
   signal   IF_Data           : vector_of_slvs(3 downto 0)(13 downto 0) := (14x"1000", 14x"1000", 14x"3000", 14x"3000");
   signal   LogIn             : sfixed(4 downto -5);
   signal   LinearOut         : ufixed(3 downto -8);

begin

   process begin
      wait for 5.35 ns;
      clk <= not clk;
   end process;

   process begin
      wait for 0.17 ns;
      XX <= '0';
      wait for 0.90 ns;
      XX <= '0';
   end process;
/*
   process (clk)
   begin
      if (rising_edge(clk)) then
         IF_Data <= IF_Data(2 downto 0) & IF_Data(3);
         if (reset) then
            reset <= '0';
            LogIn <= to_sfixed(-10.0, LogIn);
         else
            LogIn <= resize(LogIn + 1.0/32.0, LogIn);
         end if;
      end if;
   end process;

   LogLin : LogToLin
      GENERIC MAP (
         LEFT_IN   => LogIn'left,
         RIGHT_IN  => -LogIn'right,
         LEFT_OUT  => LinearOut'left,
         RIGHT_OUT => -LinearOut'right,
         LOG_RATIO => 10.0
      )
   PORT MAP(
      clk         => clk,
      reset       => reset,
      ce          => '1',
      LogIn       => LogIn,
      LinearOut   => LinearOut
   );
*/

   Ch1K7 : DC_DemodTop
      GENERIC MAP (
         PORTS       => PORTS
      )
      PORT MAP(
         adc0_overflow		   => '0',
         adc0Clk              => '0',
         MonOvf               => '0',
         MonClk               => clk,
         BS_Ovf               => '0',
         BS_Clk               => '0',
         amAdcDataIn          => '0',
         spiCSn               => '0',
         spiDataOut           => '0',
         spiClk               => '0',
         pll0_OUT1            => '0',
         pll1_OUT1            => '0',
         FPGA_ID0             => '0',
         FPGA_ID1             => '0',
         BS_PllOut		      => '0',
         adc0                 => (others=>'0'),
         MonData              => (others=>'0'),
         BS_Data              => (others=>'0'),
         video0InSelect       => open,
         video1InSelect       => open,
         video1OutSelect      => open,
         video0OutSelect      => open,
         VidSel               => open,
         dac0_d               => open,
         dac1_d               => open,
         ADC_Sync             => open,
         ADC_SDIO             => open,
         ADC_SClk             => open,
         ADC_CS_n             => open,
         ADC_OE_n             => open,
         adc01_powerDown      => open,
         BS_ADC_LowZ          => open,
         BS_ADC_PwrDn         => open,
         BS_ADC_SE            => open,
         BS_ADC_SClk          => open,
         BS_ADC_CS_n          => open,
         BS_ADC_SDIO          => open,
         BS_RefPll            => open,
         BS_DAC_Sel_n         => open,
         BS_DAC_SClk          => open,
         BS_DAC_MOSI          => open,
         amAdcClk             => open,
         amAdcCSn             => open,
         spiDataIn            => open,
         lockLed0n            => open,
         lockLed1n            => open,
         Sw50_Ohm             => open,
         pll0_REF             => open,
         pll1_REF             => open,
         ch0ClkOut            => open,
         ch0DataOut           => open,
         ch1ClkOut            => open,
         ch1DataOut           => open,
         ch2ClkOut            => open,
         ch2DataOut           => open,
         ch3ClkOut            => open,
         ch3DataOut           => open,
         DQM                  => open,
         sdiOut               => open,
         amDacCSn             => open,
         amDacClk             => open,
         amDacDataOut         => open,
         dac0_clk             => open,
         dac1_clk             => open,
         dac_rst              => open,
         dac0_nCs             => open,
         dac1_nCs             => open,
         dac_sclk             => open,
         dac_sdio             => open,
         PrevDataIO_p         => ChPrevDataIO_p,
         PrevDataIO_n         => ChPrevDataIO_n,
         PrevClkIO_p          => PrevClkIO_p,
         PrevClkIO_n          => PrevClkIO_n,
         NextDataIO_p         => open,
         NextDataIO_n         => open,
         NextClkIO_p          => open,
         NextClkIO_n          => open
   );

   Ch2K7 : DC_DemodTop
      GENERIC MAP (
         PORTS       => PORTS
      )
      PORT MAP(
         adc0_overflow		   => '0',
         adc0Clk              => '0',
         MonOvf               => '0',
         MonClk               => clk,
         BS_Ovf               => '0',
         BS_Clk               => '0',
         amAdcDataIn          => '0',
         spiCSn               => '0',
         spiDataOut           => '0',
         spiClk               => '0',
         pll0_OUT1            => '0',
         pll1_OUT1            => '0',
         FPGA_ID0             => '1',
         FPGA_ID1             => '0',
         BS_PllOut		      => '0',
         adc0                 => (others=>'0'),
         MonData              => (others=>'0'),
         BS_Data              => (others=>'0'),
         video0InSelect       => open,
         video1InSelect       => open,
         video1OutSelect      => open,
         video0OutSelect      => open,
         VidSel               => open,
         dac0_d               => open,
         dac1_d               => open,
         ADC_Sync             => open,
         ADC_SDIO             => open,
         ADC_SClk             => open,
         ADC_CS_n             => open,
         ADC_OE_n             => open,
         adc01_powerDown      => open,
         BS_ADC_LowZ          => open,
         BS_ADC_PwrDn         => open,
         BS_ADC_SE            => open,
         BS_ADC_SClk          => open,
         BS_ADC_CS_n          => open,
         BS_ADC_SDIO          => open,
         BS_RefPll            => open,
         BS_DAC_Sel_n         => open,
         BS_DAC_SClk          => open,
         BS_DAC_MOSI          => open,
         amAdcClk             => open,
         amAdcCSn             => open,
         spiDataIn            => open,
         lockLed0n            => open,
         lockLed1n            => open,
         Sw50_Ohm             => open,
         pll0_REF             => open,
         pll1_REF             => open,
         ch0ClkOut            => open,
         ch0DataOut           => open,
         ch1ClkOut            => open,
         ch1DataOut           => open,
         ch2ClkOut            => open,
         ch2DataOut           => open,
         ch3ClkOut            => open,
         ch3DataOut           => open,
         DQM                  => open,
         sdiOut               => open,
         amDacCSn             => open,
         amDacClk             => open,
         amDacDataOut         => open,
         dac0_clk             => open,
         dac1_clk             => open,
         dac_rst              => open,
         dac0_nCs             => open,
         dac1_nCs             => open,
         dac_sclk             => open,
         dac_sdio             => open,
         PrevDataIO_p         => open,
         PrevDataIO_n         => open,
         PrevClkIO_p          => open,
         PrevClkIO_n          => open,
         NextDataIO_p         => ChNextDataIO_p,
         NextDataIO_n         => ChNextDataIO_n,
         NextClkIO_p          => NextClkIO_p,
         NextClkIO_n          => NextClkIO_n
   );

   CmbK7 : DC_CombinerTop
      GENERIC MAP (
         PORTS       => PORTS
      )
      PORT MAP(
         adc0_overflow		   => '0',
         adc0Clk              => '0',
         MonOvf               => '0',
         MonClk               => clk,
         BS_Ovf               => '0',
         BS_Clk               => '0',
         amAdcDataIn          => '0',
         spiCSn               => '0',
         spiDataOut           => '0',
         spiClk               => '0',
         pll0_OUT1            => '0',
         pll1_OUT1            => '0',
         FPGA_ID0             => '0',
         FPGA_ID1             => '1',
         BS_PllOut		      => '0',
         adc0                 => (others=>'0'),
         MonData              => (others=>'0'),
         BS_Data              => (others=>'0'),
         video0InSelect       => open,
         video1InSelect       => open,
         video1OutSelect      => open,
         video0OutSelect      => open,
         VidSel               => open,
         dac0_d               => open,
         dac1_d               => open,
         ADC_Sync             => open,
         ADC_SDIO             => open,
         ADC_SClk             => open,
         ADC_CS_n             => open,
         ADC_OE_n             => open,
         adc01_powerDown      => open,
         BS_ADC_LowZ          => open,
         BS_ADC_PwrDn         => open,
         BS_ADC_SE            => open,
         BS_ADC_SClk          => open,
         BS_ADC_CS_n          => open,
         BS_ADC_SDIO          => open,
         BS_RefPll            => open,
         BS_DAC_Sel_n         => open,
         BS_DAC_SClk          => open,
         BS_DAC_MOSI          => open,
         amAdcClk             => open,
         amAdcCSn             => open,
         spiDataIn            => open,
         lockLed0n            => open,
         lockLed1n            => open,
         Sw50_Ohm             => open,
         pll0_REF             => open,
         pll1_REF             => open,
         ch0ClkOut            => open,
         ch0DataOut           => open,
         ch1ClkOut            => open,
         ch1DataOut           => open,
         ch2ClkOut            => open,
         ch2DataOut           => open,
         ch3ClkOut            => open,
         ch3DataOut           => open,
         DQM                  => open,
         sdiOut               => open,
         amDacCSn             => open,
         amDacClk             => open,
         amDacDataOut         => open,
         dac0_clk             => open,
         dac1_clk             => open,
         dac_rst              => open,
         dac0_nCs             => open,
         dac1_nCs             => open,
         dac_sclk             => open,
         dac_sdio             => open,
         PrevDataIO_p         => CmbDataIn1_p,
         PrevDataIO_n         => CmbDataIn1_n,
         PrevClkIO_p          => CmbClkIn1_p,
         PrevClkIO_n          => CmbClkIn1_n,
         NextDataIO_p         => CmbDataIn2_p,
         NextDataIO_n         => CmbDataIn2_n,
         NextClkIO_p          => CmbClkIn2_p,
         NextClkIO_n          => CmbClkIn2_n
   );

PcbDelayIn1_p <= (others=>'X') when (XX = 'X') else ChPrevDataIO_p;
PcbDelayIn1_n <= (others=>'X') when (XX = 'X') else ChPrevDataIO_n;
PcbDelayIn2_p <= (others=>'X') when (XX = 'X') else ChNextDataIO_p;
PcbDelayIn2_n <= (others=>'X') when (XX = 'X') else ChNextDataIO_n;

CmbDataIn1_p <= (PcbDelayIn1_p) after CH1DELAY;
CmbDataIn1_n <= (PcbDelayIn1_n) after CH1DELAY;
CmbClkIn1_p  <= (PrevClkIO_p)   after CH1DELAY;
CmbClkIn1_n  <= (PrevClkIO_n)   after CH1DELAY;

CmbDataIn2_p <= (PcbDelayIn2_p) after CH2DELAY;
CmbDataIn2_n <= (PcbDelayIn2_n) after CH2DELAY;
CmbClkIn2_p  <= (NextClkIO_p)   after CH2DELAY;
CmbClkIn2_n  <= (NextClkIO_n)   after CH2DELAY;


end rtl;
