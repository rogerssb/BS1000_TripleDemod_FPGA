

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
jeN9kBVWeZmJ9XOrLt5doMZhfkNE0hibaag5IsZny7wcSCbHzHmCrccr3rYXU0YpvMF4Hh1BBxB4
qEjIsd8Qug==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LwFgAK9zAx2XBnmXZBbJMir0Ce+0RlPtWeodO23ubQTVvXh9vIIkmwXz2vZHwYBR36ttM0GnDJNI
gNKH5GdFTduCq7Ij5O7pD/bf1JGozotHDQiXdBT8okYbBbUMfiOYTK7DBhY/9m4BJVzzleNak+v2
7KY0iTRNNbAJppipwY4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
1A6R7yh4xVuKpZLi7FbnhpjcGtQzhrKHw5usVtsuh8w5wqraSqWIq4JdsNUwuJbdDVU9+iJ/XCxe
CmLvrILhqsFDMNzCMh/u0KSAuwHr5z2VlTLfiwobomEki5o1gpNcRSHiVdL8UAdLx8r+NFpZmTDW
oZUZVB2BTRZdAeK6ZaA=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FvgKmauwQ6gQmSHzCBPMYwkdBkEK9mNkHSLmBTD9+GioqizgHG8NC3d4JFMXKgujGOLfXViq7MTz
NtF1fxgnA7qnWbO+x3kiXjQoNTfv4Oj9v+6J5gws2FauLayTLBlxIthSpTRXE/uVhq/JHUBDD9tP
Y7i/+OO8PUzo8co4OpJhZ/GRtF/QyVO5kyKgyfwYBcWmefeS+u0amYvxbtMwazFbwIGYjuPiyYiy
9Ai8qPv3k5PQF+mLABkosQRseGZySnDYcP/BNMM5mS2+aLXHOc8q2V/tTEWCzchiyEUWoVhi5jKw
LwBg3j47HFzzaNQ4/4qrgU33vYFmgB4x35A4dw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MEh5lfgaayixZWnkLFgtpYfxyUgCkjB+PiTS+xnnvbarCN4QcJAU0RHvKrTHcpXBTFiYDiljwqL2
5SAlSCoH8rMhdDOnu0MaekySCSI03TlTapiHS2r6ERxbI9XHw/ttTWFfwmsYjIaSCfmd7ffLq4BC
1fsulyAzhY29sMXeVjR2A9x2/hwLHgzmDyULy43LV54MAk/SKeRoannrh0KU3pUw8A2lZYx8Z94o
c5B4//wV/TuJXubjEJeH0eSRhzSp7GqyjhARvpaSiejiz2HAjqdFo7TDBsIhgi/poN5PHVdyoSI6
zw5ouOkmYCThT7/ioybtgFYweTIsC0WWFtDdeQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rr6p8CbdDU+FXi5rG+oDWTUK8K6+hgThbFH8XWrq7DZIXLkN0H3iGOuutQ2/B8Dnnm/S/WvD90eX
hNZvjMvroenj9JfGyBVsjMUbQefjcGs61bkKiB5Hn09ua0krokb3UjfLBImpPSnARmaQScdOImvu
J3BRHM/8F9XTdHLsZ1hYZ8AI1tpBP/fPhmysNKN42ukKjxRqICWug/B1tF/sTzqFJQsCmoNu9I4P
g39F/06VR7uvliAc+0M9TGxi7fQSllRykt8/j4qHyWqaY8q3x59uC5M5aKmes5Gxexnqw9UG7JuK
+AkmfUUM5CaegDf7Jw5NgtOKXScxjVGKYbWXlQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214080)
`protect data_block
3ZV17ktu+MpTfii6w42ch9VC2VxPDia5WYgj2VRV5A705O84yWSJQHXSEO+FT67ablfktvBh0P3T
bJlJdMBxneiot1hFgrE/h2LLEKpmz71w513l6KW87dXQerj5gL3PWjxEQK1iYl+pUgz3JaDmOJax
MTvLnFh3YNpg6r29Gc8MvQKqHZpsylr4B1SOswlppJHJ9F8JVx9VRILX6GfOxHnCB6zLFm8ylaHS
R6CQvWmjVBC99tX2TS48k04+ZH3uDdnhM7F4L+v4MI4FIDYR6K5nd5pWYiKd/j3j0rGspH9/d+3m
XObowg/QyjqdeGwXFlZlJ7oXMaTWH9Zf1hBF6FeFXrZVo4zJc/ZxUJc+DjtYWeJ8UM4DnlAWTLm6
BQJqA4JE/nSXiwdHSpndU1jV05QPVWdXcjEE3IAisyCoH/4zh/OGHcEiZo0MkFzLJC/sh+gG0kbq
s/Cf+qNAS6XOsXpLm/cFq4yfq/dljrAA6Klemh65UXcOMjJ7G5Ip/I7xSoSApAuGX2z7SZ1sX1pO
FgMGLhZa2tJJGRsGyo9eTI14sqkK35AC3i0Y1B48YrKP4kMcKIxRMIRgqAbK+u7aWVT+ffUAPfsL
oESgZswhK4318+14dLJ9A4XKpLrUceFZUUL5uf265m/CKr6hLwtXCsE/pQy+lSWcRZ/WytPx8yNY
qy8kN18FZx4vnJDMdUz4ekq7R23MCtZwLwVBhPZhKTSQwhgSY6jzKVI2o4St3dSFl8OrgJHSp2tW
44NZD3bkxBneMjFEKGwRzPWP5EKyB30v0NXSzqaROKDoF5dHGHtJFqbi+8D9Go3CaTUrAZWbj41r
U8VaF85bkXBt7njmoS9TuPUIqcxCaw5M/I8ng+w+h3gslJg8HGCnUNhyySMMRFCSv9sxQO8YSBaD
IKAFXmg4NZRnpC8Vzw3CcZYc993ASJS57n2ZslY1dTBnK5nUK4QhymcgLxTDGOB+jlttTZiTXQXv
rddO4iS2p3+YNU9M+Nr/7DxtbUfJ1nf/ivPmIwrl05pDIHZyOEa27kVyjRChgNe5Wqmn5eE8Q0g4
+/C0F3Yd3Dj4QS6210w02zv5LGRN4PpbrKVcjFemS9ncL3x/M/N1jHpiqTt+W4Ok8VDUg9DF7kJ5
EB+rWNo8ljJFY0aAkIaz7C1LepB85ranEhcvBoNLrXNAP/5tPPfZcuqd4HHEbbHn4/3EvXqdYOgk
yta2n5L4F0gguw7bzGOjkrJ1Du9Hi41JfjfA7Tvyu0odXqJuoTlT/zxCuHhlI/JTbUxRUWmGNdsa
qW/FbRG5zLUCjws3fRPNIvewsw1vxVWQM83r5Nn1SEBVQbYVaLvZerauiQpYL9Lg0xkbR2AgVZTD
OF62EneahdJjav+CQHBvCm4wvDY1bMCaaN9j/naRNAxfDy/KZsWVDEQogY47vAKLthGDUYjs6dtr
oa0iKd71tThbLJULUl97aeq3fLxID7KRDCFbB/SmhMSpJNNJg7tecr7aYcWXI9VVvu2ExswLPtku
R4jZr1oE5PgmXBbV0SBdjYtbg2+z/U2vKq5h71kIjrfljMwgCeCJoOD4L5SCHbwBHYZlBsd0WVCJ
PELUCmKD3lNAfZo+ylHpk8KawoisOVLBUiKgjdNBO9BloyiXgWgLItPVTy3dCNyFiuT6VQ6w5Nc/
Gk8Uj4+v3p/uPcfqvsAidK5doS073w90MsPs5jgcohUTrQZa0zwnyOq8vkpU5tRsuBzVL1hjnytW
+90LeDBGYhbIGgCEGS6cdT6uxcAobzvObrdOqMuixRhQhPyk84AF8tm+tA1D98slN3TbCw0eC9IY
MVy/U4tPTDpN2kkoN76mYPs4+zfcgfg9p2IwQGyLvMoRiTBBe9Ry6fgbXvEmCsVsRnfPd+zCzo34
Z9u92GCBkTJ6X+14vfCtVazJb6nfwj+ZuADRW0tmLrwBRXG3KnNyW7ZN2nIZhVxuXv9nRdS7AmeI
OMpwL3ZA7TBBT9hddsZexPTH+bcKwjaIGQY4ITpKIU9ysogsZOqzzRgNCtuVqBNxuXpVNnFZy8SY
k02n5TsqjTmmVgVdnWrwIdKCHwLBkZ/QvreNu5kQs1IRmImrBpdVKmyPgJCVA3zBoC+vsoePixn9
aQWnUsBZgb4fZvVUm+bewCgqyBNw2fYwbbHBYJoalqM5arVzWC7PAKyArZmKcabqL+7x70LTeRy0
erCrP92Nz59CF/bmvc6uJhlNreCQUYAOx+oapFoznUpDyBGJX6ZxulhXZX5RCOudIdSnj9IdJBJT
I99L0opbFGhwLSErroWLQ7RfwKygi9NvGEgLop/LEKTxp+oW5AoSpTbax8tR31VHOKvJLlfmGH1H
OoPUlDoZIOsVKHXGh80jHMtQQGRjY5bZpB+OURzdvm55DxfTW9F9JpIYTWRZTweDaNtSeKNah1xy
+Jqe7GBXafuTUCYKy9ofkD2SRWsCKSuBEuES0Hi0MM0OV+XJz1acC9aS7AorW5zpRnZKt82nUJMG
tzkIdZW79pm+DlaF4cj+5W6joaqdkp73tmrxEl5SEL9EDffT6b68fJWKkZfVWmjDV2TDVxBUlbxc
Cms99L0Dqw38SFZPJl1JXkfFJl8IjbMTKezfg2uPsLDDHodkaANabFjg+sccGRWaKIAIjYpP4nHm
rKm1jMm8+/h2Z5cn/cEM00uX2gXxVyyliya9y7siWiyKxMs4eBqnkwr7/R6oTGgo7eEuCkeSSM+H
oABKQeVxHPcagGfzY2KILh6fcesUX7MPIOyihObswYjNIKfv6T7ZuCbCOX1cU1IAn/XWFxiMf1tu
Ib29ABOUoZIxdcH6oLTQk/ZSRobsVSqBJSyjHUxtO+BYxzjqYhMYLGWRDQV+axniAd722bAy1YX5
jYG+ptui5V7GY689lFu8k0yRCETcXlpurR0qDgXAh8VlnAJZ9hLXF06e3A3FEXrDnZFXeCy3bjdX
lr1zk2zfglojzO2nHSf+lMfNIrUoCrdwVw+fJrhUl0EG+/uuX0KaHIMsLhvEmUv7vzh9sUzCjzuG
seuZZjZ/kofQ7Rz+sMjoQ/FXysg64mkyq/copIq599fDgttqDl0qCOyNxJ2OQ0XIl8t32st5PC6F
at3K66JLJlICbFpZYtyBGC2yQ30obBbEacr/vy6eCuGieJrtGC1qGzh+HQTGj8mrBcSTxsLa0LZR
l9nvaLkl68/VNzwIPVxRZR9V8OCqIlM0fQNDU+0jxoUMGHzdHQeO+y/frd1g1YWKfcuuxdM8e7YG
A+A2RJBLRr/PKzQicJp2mPvoxSdU+Tqpvb3IoJe/Ce4zTYtMRA0+4r+c8t+R7mXSMUMyaS/0Sugs
FoCrLdhk8MheszMvO1SzJZCj5TP6vUgpNWaH11NXevzjNQRmW17HySEhh74HoOvKiciUAytkCLoz
gto9U6IqiFVC9x94AHQu46S9r+Hvx3l5TadTJAvNS3SWq+hhEuogSDn33r5dWCRKdyLl+SP8JuGa
RO4SwW3yDbusYZACbKVU8v5Yf8UyfzU5E4YlqQiPsK3ttYCGPUKdxKa7oJ1VUifJapuBLT0PNRZ1
UNJb74IGkgtruEwwWXxPPD3tb4AnTreHO+ndY2wnZQu46Cd/b7tWuB+MZcTnCoQv5c1Jjy5fPQcX
tBiqe8WcFsuMSkv3wswdyuTagio8OJyXZcIOtr3j7jheZEKblRSTvcbOc+o5UMWYFmzi+4a47jGp
j4z49a4kErYKu39p4mg6XrXMXXKSAAgRl1TBPWzx0WbpXvm/SBjfyWQzWrbHt3Xluejy8Goj7vHJ
jnzCwtZ3yzItrfg52CC7NPjhCbaCcn5zOtAwfFhPyCqn1frFvuOPPblwMoKXdsx5JC+1gabV5tuD
j2U9/oxDbMSnzIic1jf8/TpfQg5slXG0UGhhOWW/rzIqx3qxvkNzs3FG8bIg1Z0l2sSWJa9pdUkC
IXSVWdD5JfJW9ZSgJNnKdGfI0w/MhExucX1v1LzJx5Az/kUG9YjG8fjcSvgUjr/gos8JhW31ekBM
N3fb3wxdNVJFs/rTeuMkZDoGTDGKFcuJfs/Odrvdpjy73ZKTm3K5nD9Z5JlnWdUWV0B+IDUbeYNN
b80VbFp2NOWrQ+ODdq4PkjegGeC639BoFyq67yWi7Ba5fy1Is6iDqgL89cDSk+SwwPb1VasptWYc
emI61kjgj/IfaPeZ2mGbn7B6kpyDu8sdV+scUBK9XECARFQ+0CyngZcCBcUVvq0g6Z8c6o9KBAnW
CWG/DIRRZj26gg1aaUDKn5U/ygIY7RjcOo90w8ed+1SAfAid4Unk3nJzys1/T5tDLiTPcKVrGhFw
FbPuhXGice2kfd3n4lqz/sFEP1IMmRXN0EV9Ox2dWt3JwZY+ZtqYDdlueuk4+86vNIZi96SaX0G/
1JL+D5QyMaDhmryaG+kB7NkGdWuWWGkIgBHW4znThF3PqLEl2Wbq5bl+cbmdpSRkp8mJcZwz40eA
NL3qY4c0iOCQVYRfEniSDSo627d+CyOLnYFOpQ71sChbpsN8VX1bQlGLM6RQxp1cF/DLuvtjexaQ
A7ymmNw7VTR/Kq2Mg9+eNTq+L7o8DSn220M8owzILVM5ONrg4ZCthKuLXf0uNy7dRPeTcqAc8IbY
bSnCDYg17xhgggfhufw6UFtoDN5EqoxMKKlkgvC/9VauslL9phnx6DNBFq+GvyFK/SYXSo6jMCsB
XzECScEMzA/tQicPNBj0lFH2vx/On9qtmmmpjhSBJXDM/3N12fmzloyJpBi1crpd7HTCyhVIGb88
52s8IGu4lxphqaiYI/jcW6+uhYndpsY+EUVibeO//4iFpouKR0lA3dPNWufvafbIZVt4oe8ulHnE
FM1+qgM+AUQa7XXhFJMifGFtwxLVzYuctJ+5+GEuC4qRmGLFul1+BQ4n3frGASu9bQRNKp8j/vIB
IvpbOTWvScVMafotwmd+FsinFtKNqd+9Bxpv+SUnVJN3werO1ZEeZB4ouxWxrmOCgy7GTIpJ4Ms+
7ncJLsrVKfcT2xq5LHtGfoWZqq1rJUo+TMNiMninUTMpZtTMGcrugTllvHEooH4LHJnfYcKigM6f
L/K6VFqaBxYpBxXTqCBgxkXrFMfueg4WVbI22f2Nie/WzBEeHdH1TM+djnmT2zypKwTc5GfuW5qD
RvOTnoQ9L8d90nC7NdFnDOZSTHWTIP1cVGCsr4uP48fGsrYUERXUFPStdBRCJjDpIqqlqfo7xsrl
xBS6rKSYDJWUJtmx29Mg3/R08vJ8k/1OTYpb7VvbtD9sqWWK/oHQdPsvtQ9V327QKBr7XlexOTJQ
d0eboosQN3tuZd1/w0dz6KDezrC2VBe0CrsVaxNTOgS587nmg6w4qvwzS2JTbU0KLhqOpc28iK9J
Glbu6Jjzd0OIBz2L9HFbXR0CoNRO/As4/b8MzSG2KtHF/AxLP4p1konkeTOESpqxTfFI+0RnqIII
vGuMmiHs4QpAHlpf8a2l8I1QyLSQqdMtkS4/gGilooJ3veIqnpqT821clS3PLCRod09BKalF4MOc
ZCXOQQwFM7S9HoWd396yUmaGZBozKcIhngNH6HuRsxAjXB0N1OR7djPvMYQfVBEvu8IlWomxdQ6A
1uYBdji9n6U0ZoO/w6gu94y6fb5jrVGQLRHg1RbVcHC+Fm55kywQl7bgRGo4fDmFsSv2uuILZn1X
Co+ur/QBg38btoJHkTND1gH3JCwO2U+CDPx+uoGAMRLBw2T6yrf9E5MWfavTZWNYGVQz7Hu428hj
12dTaTgAL8zV/hF3Is2/xVSe0NRa454A2iyPOC3sACAghmN8LeKQuOlyrMUg5oBPBN9RSqOttzps
LKdWuoGrJYWvCHVP4iUv9ar/6x5QedqFjNAQKeLHKwQqeQbkcni+A1vBzzMmqz5iPu0/IqA2uI45
PAvvThWxa9MF7lchZnql2SIPI/Vh/W58DIhvO+1pBbTBwFabAFVVE7cEr5VCU7vVfo+TSMFkvyvO
E/OMYHvhR4isXNZzdip2lIM7yQjudLeZj3HlvJI9ZNoiK9fkj6PUVaQP7sT1hBq6FGwTcSnppSvu
1umksqVANUyKn87rVgymiX6zs4Ajw1o72iLVQNL4iZi4PaK4ffY1dvZqJz8Tm01IN2JlNR6YCtHD
AUDq0yh2jNXI1aYM6MJbcHJZjRt5c2QmSaqJxBz9GHt5npw9/x0Ze/pjAop9Knp80gwQYiGOz2of
uMGcVBqQitZajOIssOQzXsl0LYTYjCJD4dbu4pMT857JDr8+R4tG1jvBUvPLsG0z6NwUC6bN/3W2
NjWV9po9DpFRlXFRB9EmAZJ5HxYIYAMQ8tgoL8fx/evOuA4sjMxBlVLnvsiNALR0wh/1zH5HiWjW
Dywi8qBlZTHaePFpAxyOBWkRGqlDWKOLrqMyxHObHLugxFxez2W0liRS9qLlSCcovj+0YntAN91x
CCOrNuOs9XElR4arkMSk2j/+vEPyg7fGeZdtvc9ucpBiiJ4Pru82az/JfdnKd6mAQckb94hC06fm
SWqOv5ctkSJf7b5NOcq8e63mrirJ/rFEBGpnYncLyCUGpkSCj6XsAFVIDQbyZUGjYQSGWgfEBLxS
GaeYWoJSRve5ssisEThCn++wYlJFmQxtAdQUVLQQ4cOgM8wfWMEBoDk5fnaTzt71orfTftaGHnY4
uLFp3QrttSmPzl0ZLluYBKdro0TrXJabeNAQR0XJlxeuPBj7Czle9jsqZyUYU2075fBeXci+Kf5B
kPXbSJa4lxeGFDLsfegSyfhK4a1bkPF4VPxzz70y5n/oTHTcVKIsz8Vf1KTxFVpoumaFb5SWtM8l
YQz9QTUO4uR9iguCs4LLn9YcBELDxqI7V4XAu/SfgWi8bGPgcu/GzmiREW8IPahxc3FuPEXZ3e4A
M0Ap49jR/IcxFYYzyQ75/dr6JhGqkJsgdMOIqbvzbPCt96bW//AuU4/nvAprcK97b2R1KbhL7EUe
/TXqat5MM4u0+VpvcJgqsIzAyChGAjF81BWTFFSAl+b/tNcn6+jO/ZeOdsstN3xk4RmPmvqrQzZK
2QwIkxWrfe9NFQwqwA8swRels2svGMvrsTtdZPy6umonGvIpD6OFLlQSE1+AQkNZuABr6uN4icYt
nmzhMFZgZ0ZWl2BqY4Ju0btnhbWKnFfqWsF/mXr/5TS10Dy2wIB8++B/oclORy1/8lmY7XMVZ/pF
6RpumaN8NfzAZ6dZfhv79K3IRz779420R91RHSOn+Hj2hhU/HrsP2VvxLXKiZ6PBNh2hE0vZs7xg
8UrUrCVvzSYfsO3+7El/wmhQo/s4sGq4jCgn0ii0KMnHzC0NCjaduE1w4cy7xZP+ID7ci3zxyPHq
0T79Ls1+zQmC40ZKh1fpUBACvHyifZL7hpS8/7wKAYu8MR5/yFSoZb18DmWWCQ/nuBrUiYdDo6XR
jCV5FAeVvEkr1GvKhxkp6XIkLoYKg+Jj7lwU8kj7belC+Z9wqdXADYThl1fA8p6gvDMKHYpcr0Jq
LE5zAhxj1DVr6CcWUp/vFM9UZocf/8mIqjxHkHhQ4MdNlICHpztQ8VKhfk31Kxc8jt1KOV+P/oKS
tqgs0MnoWbHq5H1MVUeV8ERLKhUufRT3SSnFsM4HHhxzdkmPKiCc1JA8689MwbdlWrYPtOHxj9YK
S4n9nRiYzsFkig/jDcc7uTw8BlpNhzLd1SvN7dRocen4Fs7ge+BLeLoTPkrukiMmxwSanjkvoJN0
aBye4fZN9pz4Y66k8iQn6wqm+7mXBLTio8Lee8aqj93MXAMyNblaQheaFplq1de8GNcjPrCixf4b
SIgSv8be0c0fPnsoVRStCY/nDXTLxvM+lt4UgwJjz932oXC/114H2VxKQWCv7GoaWHYCyupqKGJt
nJF75UgTdmPP09lJS/1Ks2M/NoiZAqlQJgmqA6Y0Q+NyCzfnPoxbU4+JqBos0GBd4DHYj2lqRv4n
z4fGwflKvCuI/UXYkqhnpaDtxAHO7le9uFJkAsJL/MpCfnie5JI1hjkMTfYfWBAqgVW9rIJJcluh
0KG5EJDnjMb2omS/tCwqY3GMt0bBeJ76paYSoJHz/D1Tvg2lYrc10aDUORFUp4cemjyR0GAhxyNc
pR44cponxzaxoLbBY+oxEeb4/Zw17qNBUSQUM1GETj7aMncA0touYjn4qowDM/zm6rBdSNFggs4s
Eoh4cgkJNyAjQDFm0ZAWP3H8LSo7UMOPY2qATay/Gmu6W0bLLqf2aCIqtDu7+D0tex32aYkJZ2VS
kGtfJtU02hjJs9zCjZEwzqkgxMBeFYVo27iNyr5oLvyJVSEdbizapk3NuCoMVn9TrLEDRLRySmBh
4FtJsd7pPOe036YcJKSAAYH7zqhAYAsjEZrJao1eNn8BdA3OpgFhctQZSoB7GJmkMNSJAO6huF2p
vUE1wPdgyP9Oyq1vuwBzLTzPMKjyLd85MyL9sPVvhdxC3urs+WM/C2gPcFt8Mbk6RaqrAqlBSPX5
v8okKb0ON7I0HitlA4JCsGCogY0Dh+WnvmjjkCdgem6CZEe3KLRFG99vun46XJxufXZ50Iiu5ly7
slpfnc7TSJjWQ9C+c26T6l0etW4JrFo9tDJhBk+Ra9aJwot2XFRaz34Mu7bzsDIVpZUYHF0/WNoq
UP0WqJrMNslxcMMNbF9DPs9o1Os1o0FW3YdZQFGAnRKc/ThxThmC6MNevdgzTwT4TDP3+pBKIhBL
wQvmzkgwLnKz97T1lT9GCrErhxNQ077AWkfvqBxeenhIJbn94m1q40kEfyFuas73mk4UwzRAzaB4
OG1pJmbBKCftrux8AgkqSqewKw0MyXVy/QSdAI5y9QDQ6rSFcG7VJVF/8DTKYePoB9a84dQy7amH
5Ytdx82CGTe4r52zV2yxuRODLrrTjjrNoFgge+JA2GXTuaxUk6/tZLiVkvoteEbC+CBg0vOUuHig
78dr6pEFqGSFsro2JuuoxScZaonG+doG+1dUgnxlZGb7uwFnLWjnqt8gB5qYOG0Lq4ix7MJwYbTi
Z3TQyb0e1FllldAeS8gJx6vuifT/NHduMSnch835DYBWkcFDXI6i3Kv2MFf4nO6HzLKCbtXvcH6O
lSpS0TJDi3aQ2N8OleOo7P/fyqWa3B/gK0GOFrxTLIXP1mAA28evPAbrDWwgjrt2VqyN5vmYhcJ7
zNtcYoqqfxPn2aALr81bNXtUBV8cOe9o1I1eEDgBeyhIo/JFXTq7YGMAA0IQ+TFEgw4Y4yS/be+y
aA1saxcWzEIscwm8Syt3LHQkGJJO0RhUVjSQrir3dZAqENRJIw1NjJwhItNZOmMosJ3jvKSQFBy8
JhTkdSwNSJZ9w2x6n3WuQY6gBvu83kghih77iq1e2TGvjSGOUb0sOWbYbz3CEHmJQJ+9jMEQn3fI
+Afqp+UinBLpABOSTTaYwKeYtua567tE0HiH2YjFREo11ORfHO11sGBcxZKLFXxvH+FZjpsgv6He
auKLN3I5Lcvv3oKwZexIbn4v99DpGKpfC0XoxlOJgJJUeVmKFRRGxiWpP95xWLJnwqCphSp0vYIo
rB5MpGik+83mVvAbAdEs7FWconfOicM67bvkhkClNX6n9mbmsb3ttHiS7btIbBlWdqCRo8ur7zvS
ElAHPEqHU+O45Y6lTZywXu0Bpo1y/IIdAesh13SA90TkGP92vKCVETbO6J8nGelOXBALqwFgD2HC
XUZoagISKFfDO5r7/yG3i1RQ82uckJ4V52E6jiRi1Uj9uuLxVVc39lFygOYDT0W+fkSEXzL4SfoY
QQKuAOQFiignJ/kwdsFecWw3jaU7iom8f8HipYieXd0ku5Sob32b0g38mKxLGFJ3TUlOA9SfJkUO
C8ZNNHUVPuuBIEEPDa51Rm74xWfiAIx4YRDxQNkXIWCv4TI3End6Fu/g1Mx/moEVkI+jcb6vm6V4
Tn8tCYNF24ThefFz062hZcQ6k8Mq6jZA7b+hVt+JWaMpwOtAQ6VJOQG4ruYw0kUZynxLPgtWKksq
wvQuNgObdjcMmyK9u/YEY/pn2fzpFp0rwQ0f71GfYa9p5EGGlmkPocIPI9/yxzjCD87anTjAp/Nc
rRCPkYD2kcR5zF0y5VP795B2J11q9yxMaYfUO4LbNa1lpY60u/One4BrPbVNwTNAVjgPd2oouYtf
YTBcMT1Km/XJnmDyDZXY/O2C3579UwtBlugrnXjBL2/vI6b6KWlmxmkbSFli7FsYr/G2xPS10nsX
DF+N5oChqyTmZiCq0GYz3WNp6/TKrVKsyYDBxOvXdneIeqqGYXjSsot8zMUNty3hb+dP+obpaKuA
pIDpWNWdu3TMh91pqkHw6UbUfcNfGDkmEf9UAMb6UmVKNmmQtecaeOy3vz+CPX4vCg5CDDqTRZ6W
uPBNWnC8QZDgNYaN5pibSmzrz692RjG5xw1NR0gap8x4CRnBYnWvIDuidmEcB7Mz1HFMh6cHEOkT
zq4AOpeoPykUJvHGTD59fxeovM/T5Eo6cRv3p3OG6gT148xHQILclhEYpN7Xur38NJI0UFktD9Ed
QSt1Ajqm6zTN0fsvG1++v3xHjtT0AjSCpWVi9ffr7Ew7JaxFUBoJ7x/8Rum4RwwPicp/ZlMZtw6R
q5pauZk/NLXvfEH2iMW2UgUdCoeNGqqWcC9DCKy9Mx/+D8Zsui2bpXQ5br2sVMPDOUZga8ZWzb0V
RpuE0RRJApOmo6hyRiFwYj8O1OVDOhkl9VM3bt4NMSTS0OwDAvPGmaiIXnz10JgDfHbe78veqTD6
voYWY8w66o5QhHCi53+iYIY5+XTBuJ7mb2N71qa98GTMw4HBVNxvFPZPVSSkGeCjJhGxhGEo05UU
DEUSB6jS1XDbup3Q5zpe73EeWZpHPNMhrrb0S8rLk8B857J6hc9s4AqAEavKaN5TQhy1+qEiqLka
mY2tSDjE13okPppN+UlCSzTSq9JsQiT941N5J00fi/ltNBitT9ErBp6HC7Af587O6za31a42v4nx
pbsEwBBd23IoAqB1A44usWKBrAcXh1MfHBcMRvQadB9QK4N/uLTi3RYl7bAp+u3zH8MxgxZhsltC
bXaDyfGnXapv/mAAfDuSA7n7O1Ly9k3BDrd7uFUikzc0JgL0KEs4qjifJodG8aFHT0R5pXtcZ/Zy
qdEISJSRrJ95pec+40M9enAYDfZ4RWws3odIDCndtRKG/YO3NMZ3imm7IoaPCMo1Ab1I/Beg2Lck
pkqMsMiVnPNe7vLdSfxefi3hi/6EkkUDNIUOckQL/cSU+xJmPSUSJjdNXffah7EHp5pgahHJ+fqv
9f3s6zTM8tceKWEFpREhSYdVCbbv4cdi8sVcW8o1f7Ipt+EGBtfkCIRWqkOhpq0Sk4lzazWdz8lG
u823y6HjmbUw9gdYMvXamwY/0/ugcWb5d84/3tKMhSj8V6wh42AnS4XkqW6biyoezqrrs8IUQ24Z
f4YuTN1lvAnpzhsChdae6WLIGekD4pZheXEo2DuvxdDsxArtRU7MADZXrIIOAecESjOqk2E99QxO
UyRjb1F3L7fG1v1VkDmrWl6djKjXsSTmf7m1GwFyXNcKTX0CitnvUmdtebZVwWwEsNVKYgBn7s6v
STnBfopHSfiJuHPrzBgpzbaBkPLSplEHCzjqC/axPXUk5VWE4hN8E7vlo0nijBaHAGsg04rY0X7D
qBtGu2EhN08zho4SyLOqBXWIq9t8RMqB/WgZoSxFWDOC5TO06LA+E4+eyR3OZpBAo6x58JK24LYB
cMSv1jIazWoxblzopLJc/gd8U52vLjh7BywO11H1AcIvDZyosBnKAny6HDwU1YaSbeFVOep93Wwg
j5/Lj+AH+Nf3MldogDRVIUwcUCUotiCc7KYaxWmcV6tWgmUgZTaM2PRNVkBIApDnIrfWSnBW2js1
oLQV3Vz8gYirwFgYVF5ZzXP9l8T4RSv9g4TI5bEoPpxI/WJN0hjAsaAgAtWErS1lskh1GDSDlv/y
BkZliDu2sX4sSd7LC4v7NUPSsZmkemkJRLwZ81TkAra8Q6LBQl2yF/pF84X5OGFzeglKzFCL77fq
TEQiJa5Xc24+7UWKXqd1Fo8NuFFd0ZpAN0u55fAVHr1I7zHpg1Ls6zuMwnek+BXG6WHRtgIoncGn
0ODDWIa/OrVXx0AcpPz84ckMgCohcdYeK/Wp9UeK9g0c4jXN7h/all+xyIjojs/jGDnjytEls3Qm
MElkTI94GvnR7tZAEx4GVqnCOnqZVJhtHoJkKKtX/fc7xnQEzfVE/KeMOV84Wrq6SbHHY+4b9N8u
xRuQamvwbUOtCvpZWlnD4YAw3ScfJtDfJORzB2wRVFl4XqD5dcBN7gfwEtWyzFwAzlbTYtyX7C1b
W7JBAyERdzqREHT6NxEz8AjboBqnf6pc88EYt5J7qk+H+t1A/QUgWSuEGKBz7xu+eEtylBAtX/wU
q778yGUD8AnsWTlMIGzcm5LXzD8UhbdXnEkdAYtjQV91OtIDZf9gQCFDZ1vWTBWpVtZW5gvSUTGi
DsXeBMXwHOymZXugE+5ThNJlivN9uCMbMtFtmHddyHaZY7k8PvW3Td7KpnGlEToUGkUkO2ZOlim+
4ctf25010spfO9h/mmzqu93e8jQ0eWHM6ixxRQBTmD6aUjDg716ZvdSf1B/YuZ6TOigbylTm3QB6
WPKfa8/oXYl/oY4cgUudPSGRVeru30Me4AEKYN/JRNP5sAc7yfeVZIO20umb+xFQsNAm7eyzwpMW
FWv4YH4t6M8SYV0vfJq955NwlXQ+uqoVKbhaTjbQi28bGIlyCMdB1bjBuWGrc/9Le04XPNhkPrxi
JNwxEvMpp1kv/Fs4QfykyKq23NPOhSMKVFORmMWELX3EhvilQt196nCowO83o+yjbIvF5FlsbQu9
ICKzExqHTZfgJqgmPCJS0+czMTC9MPQVbvsPTho3UPtcorYoRlFcspA5Ej9Rklt38eXwD5N/Jijt
BqXBngs0WL26MRr0TbH83v99ayKRAre0StX/dIurzwYNJHm+0+zO7srSVwQUbCnlQUUXtMgyHwGZ
g5gFiwucUjp6IVOcAy3y81qHtKLPNaUcp93eJom+JsqjCzByZf36oWy8OxfX/kr8JvVXAr7APzPe
z9i9KJnK/zSREn1Pp1foDNbEeVKVDZNKVWiORgnUzlaueB0H1z5XoYOEDqZQIfZatAK1sCnd5RKf
Ne+Ln3LxVzO0atjoCR2aIQdKJ7ppwHAxqLaS7Kijv7uONW7fu8K+ZnR1tfn9LOUkaeyCxN0QCgIH
C9x6vzQIHn5jQMZKpTHxWeo8fS7vCjXp1AJpOMAYPMbo1kA7IiVpBzRp6dNHES/XnZ64g0OraRKx
idMZ2KlPC5UhhCcukUMTvWdmGikyeHYLoqMqn0yPy4eaaI4fIh0Q8LWg4769oMmlrWHshB34pT0W
4Lcm9rVU9bOAfd3aSSnMQl300nosuLHO1HJq1uSGi5/c63rD83eKjilxldI+gAly8UGfMt+kjF33
VbDH8DDclFmt6UtKQhRajjOMiAPja/s8i10rDfR+jLnonnuzbnWu/Us73OillOsw3S06UjR0pNjd
Wbo1mC0k9qcR0z+AJtn2miBALBGkNsvtaQWmDAynbbEC6FuoVUIhtL7wTdhMnhKjPDr2aV6cBCDL
9/TV5RcEhbe1UPJmC+LQS5hLbN1ztngUo7D9xPMH8AX1xj4PQSv0NtHejG1LXPLXZM9urQv01B8q
ZGOoZQGg2QjdN7uStELQ2Qkj/cRDA13Fo7wYKeb70v3FwheZPjP6cEevWn+vmv8XC8iV24HEyFDC
Y4tGnS8F0ApAaW0ET3X9u7br1ym+CDn77VPHNG4mJt0XhCMf1t97rjZwhkrw6Ias1fA+6axed6vq
/jnMqT5nZBU/aS1UaLqt7kdHk/H3sazBO0MDB+8MggDWVIs7KgxlDtIqhSc/3fBL/lOzfhtpKB8g
sbH1z6VjtecdziwdeG065l/9rs6NDuUmXjpqDUfuotnd4cvqrM21jlBKqh4ZuFQtlHAWdQ3UA/wx
/7CTe9di1pqPdE2ISupyNxG9NdC8lu94VRcRlBBrHcX9nq64mmpWDPo3woWE7/JvH4OIqvEgkepz
lXN8PRCiFXe2sKTGU7lRlG1KU0IuCzkZLtGTZZ65M7Sl6K785ovUSmvXrzY3omUpOhlNn5F29ZO9
lrHM3d75QmMEBEEn7MLrpV+GEwbYBLbCYR+1ukg6qfZdbYdKcrFSs688SYHbsHraTNbmQ4AR6b5j
C7AFXzj4kWynSRjGDOFCqRakzaVJC65SPnoYvAJ5Fj4OaYAeE9yEeeIFfp4MrrKKBLi6TkT3Jv7a
0Zvfz10VADVh3pByip0SP2tM1FcIdTP9m4Z8YYsugulmm4lPljtakkmN5NTXqBXM+azcDYJKR0ij
4VfvEOU82D0Jd+Ahpo+S4MbYToDZ5/Yld8s9GtL7eTn3jWorFqJcTV9nszOcnSmm3Kc+ZcU9Jq0l
UnkyPl7m9kM/6j5klSY0SHbmVY785j+WFNleObRkg2m4inJ3ohXpxQ0OQC/YohLa0smWokIOvkKt
HcLEyKgAKDvrlH9PP4zfRAbWLzew6wvUv4XV6S5XjXfXqKTuig1HcFbQ07f0pJEBceqTQ537nhBv
nIqkTvqjXXy3fBAG/1m3yJ+6VvOMKEg8Q1tq4GWJGRFgL/O9uPA5a9wnByvmFr7HWNCCNX7Q/OEy
h+FUEHlaHGwJv8BRkDa+/g/ssM6UkiellIFp3US3GfAHlOuKWFf2d4fUBUfIIuywrx/Ata4IyE+s
JWBke7uUhm5Pg0PfmYK2XUohmeJ9qhgSZsVejfn2vvNG2G8CsrZ/Bwgxk/VqxsIWr9cGDy7XOraX
kZlTtgwhx2iAG4xuhOPkr4TADLbP4tjZiSCc2vGRAeLNXI5h01yWuQSsxWA0n9sqJg2nAyG03juV
aY1DXp5hTlf/8yAh51/1FBXA7Z78P1ZD/QfGQEg63A9Zt9C46tSITY+eK5PIhqoQEhOrjUpH+zXt
Nd4I3tX/0qCw7Fn4TY+IOl882pKPJv8cLWYrMVjFI1f6XTdrn1CSQf7FAU28Kst/8tlQuMTZAmf1
T9OlmxGVatYT4LEoL3JfqCR2ujTJK/e57bPxI2sqQMz4bIG4zsfWS/yfl3Tn5fWi+8NYEicEjpd4
2Uj9qNmdpljZj5Q1HSkkVkm6cekMHEg1zJMdSLVjDjUbx70FqVAhGurp4pYQImrqhf4hE/R4/iun
murv5kkGpWLmK1QApYqxjYcUzSbTxMyZdTUbR1if96e6hLDjfjg8EqdmjDEy4yFcQ9q5TArcPTPa
GiJCkHa1ng83U80QhZZoRNa5argHTb+qK8QWk6ewJ4R55U07owVCdgiZWqWLA8V8Y1c7+rk75ubg
DL8UnJWM9gLVv8w0NM8ihsVwh+jeOFzb4Q6VzmLDhlc43WqH/jGDXQfK7/1D1v0vDOs9hUMqkDOT
9WDU6G5nEwFcQiIxdgFtkwf8pbBkCHEMZyJauDvjMpk6JyIr1/mq0UZTX9TMbc6VG1vN0suf+JwI
wwa8ptW8L6luysLuJOHaOvJKxmHg5YUXL/+12VIJMIfreBerZsONa+STRgapRhijoS3fe8Wc3Zx7
OEbzMJcIZtW8hE41LRfDjyzWtMHnm9Q7MGx7th5SA65rL8jvOU3dIyudQn+4CFpnbJiNfAo/dW9S
9Cu87xo43HCoQH8zbbp/Lipv8tXNmgVcQ5uKsF2AV3Cp0t5TUmwa4IDpfTqCRznqC+8300ytMEAA
lkDanzcw6TlwctWbkOpdFiilZ2ftQBrKdJ9OAdsDK271bEfcN41HEbwJ7MSq6E/RpuHxiXB7w3Rx
RgSMSID2+NSo74f3AcdAJL7eNG4Olpf7l1bLjyxLd3oOHbyQeaoxvy4OMA5i066kS2jvSzYGgBNz
YnjYV2EX9RCfvC2d0M3KxFRhESI4JEr8OZ01eolPMO/ankcJwZ5iBwMeD6whs8E5Xcrn3QEJws+Z
7Ks7D4OoOhjk32OB3a7J8AUwiF/ahtwPAokFUhBR/RLHcwcSEYEkhqyMZlls/WLpvjAEpdj1EnO2
zpxIaj74MqHEB5Fvt6yIcMC06MwgL6uEZscosjX1HhWuvDtsZgMpPKLlFamYJ4y7cOIg05Z+p9Vu
twUeSTc3enrG5BNazvNBi16BIk71XLUsqDV/fapoUv0Knz1Nlf5RiGoosG+q4779zkUa2iUAJoCQ
K6hsWiRdICMrr66ufzTFCjMUdMzk5uC7ih8ZyoSnLobEVGv6mZzz//Ioaf9eM93Bk6tZOQYg2S9k
XZW6NB0McnG9GpT4DrQO7eXg6hlfnjM0pyBiKX2YB+i2W6OCG11uDNo2tGHDodD9lw3HJCfaawYe
QLxqMn88vJlCZ4RX9uewGiBKleRiSypI08ArXXPLvVpO09sDtJYc6WAdiDVgFMqURXb7PX6Bfgnl
a1NXhtv2dpUGm6I0Bsw+KmaUVVOtzo+R1z9GpNE33rKoi+fEol9OgYoUGXoAY2hL56EOBOsTaTFa
/v1BZcM/Nb9bX7J1doQSNMiIjk2OrApl2MaGjMPmJnO9CUe/sX70vX0I2nh/D/CMDa+IGdQyA7yx
gl0HjgjHKZFxT6pNKOYt4RBaexgwHzZP1Fs3AEZSKpsFGgru+GDoklXKZ2BtE19DqIy61J36HCzV
xDMVU1gsQA4koUnKDkBMZjbxuzTjeNavPGK+VyP5wIgpH3ob2O3bHRXt3STX2wrm7J9PJM5bzNPh
2eAHGnPkliUN7c6MdG7FLuH59FDemiZ9S87r35xKuXE0KqTtsRJZnOm1k0S1JdLeponYqJiGXNOy
zOT5ycSSOIO13BdUT1myNcPvmRV++Dmba8YWBzwmmDVQN4gJvN4TlxPLyI2eAFvL4B78bOYVDgvb
F1z+LJAsDLk3fJAEpFmUCAqkEGCPsXuZYI1IAkxR+gVoTXAfg152g7+Lfi5v4KOw/3zmfuUl7gNW
B+tPmwkv5LEdUae0Y9wR7pyN3nJfC9vfYcYPEGZhxGsNoYdytueeIIKpunGLH4emzu2Jgox+oWxJ
txzpZ3/RYXFOgjWIOwRHeEloEweWUefXpqmXg/0JwKGXU55p87Ka4QAFUHkDwY2GHbeZ9YfzPFYd
EGrNup8+2zI3vlY2zN9+8kjRVe33DBx4liz9y1MJ6md7N0LbwjTIMS2/t7/gaW9rrQDpKcZjfn0Z
y8xHIDNTLjvINDkQJ3IiBCAvyigL7IPNaK0WxSK2AuvKdQsHcjLxBlUmDq32hD4WnkfKVbGQ/ACZ
mFZHpf7rFw/21tPNe0ymoSbLDA5KnanKxxibVCSo+9GF9rkBZo7JQxaqA4TKlM5mn5aegePZxcqr
o3sHZ697TQqSwsJBa5CUiSlyMiLC4Edhyh9a9ljyG3XlCIt9kZ/j8DhiX3QkE8jxsjW0hVq5KznC
AzvEjkq8G81m+jdfEbc1nmwX6d8yIZP6TkDr3IfXoHKQsIfUVhcvfzhA4azvSr4Zzb4cmfXUb4ZU
MDUcJVnA357GtegnoueQJ9w9gNNIb2wePZ+hHwGqO66TJ3z/moWEqYwzNIoU3n3iFXFzp+1R8DK4
e3ptEEw5YVSvPbrc0bVg3PY1U83u35J6UVswyYyfXhTCU1+M6fjpWsgDgk6YOY/rEfsiSUrn3Uo6
2thbA5soT9g3IlBJsfVFp+qUXjRr8i6w2ZLlHeRrDIiR/4A6HUvzLLIoOq+ulxpXgarChurWbBM3
k8sbXm4fu7oVp/3J76dppPZb0lVT/rBT7ZUDRXaOsO3b/Wld3XSRrxMhZ2eIGDTwaQkp+A32/Jr6
oBfWHl6p93BKYneWGOmIBD2p96Ts9OXQDFMR8UDvBFk5CRPS/GCrmTBz5H7U13qjm5rl1ewGoG/O
Ssd0kR9uJVEKxNDek/tTJ3HpUQPDUvCkpYtpGhMZJa/zc8vofNyzMphexNf/RcIkB5RpJaj385iL
uPnsL24YqWBsOJjGW5VarrKA7V5Rtjxxqb9oBYjYn4isp1hUcOsW5s/lWQ3kUEJmEHBLOOfbDLVG
CIgdxI2vX5qZ7e6XICe3YwxIa80vUBKj9Ud14BSE632rh+eXtI9jG3pXZ769uqE/aJCKZpQGy6wM
39KFOCkKjRPIsM7bLaGTfZqUiXyAydkutb72vRMbGz7hWm8IKXcTvF4hr7jloP3Ru3EqZjP/Kq3s
Tcs1cohjjyHYSZzKCofUMI+wXYxjtCySvOd+T6+zTBE1WbFKBMH4AmNrbhRaCefscKS7pmFQaw6e
kJj0rlx1iVbpJfRKoFkyGrpzqtDqQ/AwZxhIJH7gegDbvj83yBFeb7sJnzlyiqa9Z9iFVC5lmgkU
tvvKP09eBppIq9keS0lOCEG/JxxyDI7B9yPLIwAkwE0Vh+KsT1wT3whiEsTSQwCLzZ7oLK5iMrMX
labfXL33r9bY12Gt7tiOGVNRE625wWU+rCZPX4s/XnTm/BnVOsOaIBW7qAHkk/COYgGRCPUW1Pv3
F2upgbkA7dAP/l0ai+m5BOOoeLN2FduySdFnt1gfc8xXOdSbSWbcU2HsUUhqDO2weQrDZfdunmlN
DT8nypNbmL4KQu86Z+PGj9Hno38efSAZ/uhAdl1Kz7khgy+0/qvkM7oDZ5+L+M5P6ws+g9aDRWdF
1XNZzpnrvSwL2f4H+F1/iT/IBf+JZQ6UomvUaYcIiDfFHhGcvhLttNtsjma/zEa8dy9PWqErB9hv
RV5tbBc1fqRpzD8QjSFT5uA/N6CTTdoc2xIvvy+obhvRpxuIYWzbyjR46aHdN3awrKi4xzKdMMIH
+Ihj/zYrWwxVQgI3JABazmaJPUbI/HmLODBqbpSnN6hRvKl3TgM73+AEw9ICcvI9QLKciJIjR1F8
d8zLDzqfBaKjU1g6mNt/cIalTuQpUDE+oIPDEo9SLf9/vUMlIoEjHUmaQDwbCFZLzK4BJxBU5ixR
y6L6Q8poz8ygou/JaN8RAescuFOQl5ZR+cTIYLTAOWlkaq19Z4u2Ee5pM4NTq8EwZxeGS0SwT+oR
v9Xk4HhuNO+dRxgQG/husRBZRafvzw9JGuwxnVTf8v5Ss7tzySUD24ITJe3BQpjDauML9WaZyV7U
Tt2tz20dfSNR6yB0f+OdAEZSIhhugZy2pDmJP2SyAgZb//c4hCERvkGn5wBOGiV6EwW628d6muld
+TslorVlv+ZbrpE6d+ps0BfItWpxVqhUab9Khaysit1BxITmpIhNut1hi/LZ2CaWPY19HkXjXj8r
W5YcknJvTy1hZn7/CU9JLi7dkRKeOv52r63qOBpRGfIJsjdjU2kREO3PIa9Quye7PRYb6F3LgrD4
Equn63DHF6LA/2NkdMt7/qbcB7inaMkLr/7BzdZwzdGKIiGp4lAqWyDZeVRBq0ZFOSeDaTK9YNSQ
LxB4zu7INRNlMjrncwFuiqmIlgP2zf30si3n2OIzzchA/ELdXlNO/0f3V5dPAfZdwugvA2Wfvrr/
YzxHkq4uqQi1qirIdjoSvPKGkGx/6tot745Muf4wsHnooyrEXEXVIhv+BVzCSIkPZdTSldycYsFq
+yqRxkSy4QKT9h3lMNwqaYeF3u0Lonis9F/yZ5oB5rjKix8ZXj0o9EneQaoGkOg5ss7qQnkFlk4k
Qz1ZtLLGOB6Rh79P9oL7KTvvwJvQA1NzEZV+M1X5ujOnhUIpxbHBRImo/KnV5TmX9wlYSC6zjh71
dqhVcDvghidxDSTlf6CBqalgUtfftis0wbzgzt+Z1GbpxfgcPDAtWIJkYT1IEioE8dKQgQ+pm6xA
3wwJnlT48W00Cz15YGNCq1Yzf3arHsNUgHexGBGInspXoB+HRnwU2orjWicJkGBc+otZrp5ENjxy
FxamP1GuIsc9RqzcZhAwLcUealoLYZDFFtfU5FRotmKDUZlD6YLRc7tG3yY4HQEdzjnnBgduo0ga
a1TIbm2X7cPy2iqEGhqM8bENSHXkIL9ULdF/0fioJYddLyKR7ETxlMcOkTScxzFixIMI70kEIKcT
guTckTULkDSS4WAYqyQslLmueHKotjZmF21lpQvM595IQXuR5Ie30MRtJTYzMRYNJBwM/0N8aQYu
fZSbPqwfGX+3HwOAeoGLhrqT/IwrGKzvRXFXTmuZ6bYxn0vnJPQ6GNeYDMMUdvnlhCe/msjuvQR7
N/19YGzM4+kVc/UEcHuIg3D/Ip6Rl37zjdyeDTHcWO1B8lPK0+1pJ6nU1CnhNZoFfrlm8bFBeqWl
Dcp6GwJqTxVdN9MGEzSChEnFff7UO3bu+V/l6THrl/vvHroCpIwcCPI6rgcWaZE6YobYfFA1PmA6
9Gtq7TFNECM/mVCeSZ2wjcVUacpSE3CLB2Pq6Wtl06/JZRBwe+aDvksqVa+jXcGSC/CzL24eRNWY
djNYNPKQUwk+SvS7EJ3k5n6yNtQERt5o8CRTraxFHn3yWQTz9cQaF/hV7GkXBjWzSPCJNnpYx6pd
WBLklrCVqaKhobVsx8A2DEMLEu7uzenc6We9WSLNFT5SKpDhLaaKRrHbLs7AWvmhQzgAIF9nuX6E
2SfsvsC5UlaDBuFkNb/rXKvFYJz8Bp+YFKD1n1NKoyLMpm4aHv68mXxopwfAtNehiiR7T3CdupYB
Yqzdj7qBkbT0UiYXBzMIxD6nq4DjuEnwyYso1FMzVqJJn0Tg0zFfH27a3ctNchJFMl1pWybOAgVx
7O1guikVp/6PMLnW3shCb3n2B0nmYX5139iXbfZW7JLVOh/OhWCMbn9VMahUlu2AH2XpcvwNJ/nN
GcspQueLdGI+Br/3BLv/Gp89juwQB+DvXMWkU5uEq6LP0tonjoYbuhw09pNIbPUU72bdjTzHmBjh
AT4+wCKeV6GPj8jiJqIbTE/OzdvTT9N66MG8UW5XYpgzUncFA1AAr6c1eck24Ql5r/dW9nb0aWJ6
rG4p6qg6qXRF2sTVLhpWHfeSbs9RbyL99sQRCzSVoBze2YiEFMtzwqd9+m/zR8FA+uQasaCSJpqw
w0Yu6wUZmnwe3em0FukAqT67mEtxlLVPzrDA9LqMHdAHy9O00Boe0TaNFF6GjAvOO05ZCFP7DO5W
lqZNAK5rOQtRwqgCpG+OAhcIqtCqciTQcwA9zms0tH8tbhZrQRmt36QeWz0PZEAjguSErDHcFh4Y
wA+yJ5nQkkFPKqLpd4RL7XSJsDk0Jz9KD7ig2IDINWM64hMxohqkn2YSuanppkhcA5Z8QnCzAIOD
TnAbwYNbbpD26KOa38yxxs5yPqMBPdrQUx0gjfRPp83P1aeAoyZJaVau+6UBRS7zu+c+vOL8YIS8
SE+t0B1J1rvtfMgOACqwN1deTqcpfcn2JdefHvScawgwlh2i4+NNxCkpBTXepk7FGX7RVRDCbJ94
xZ8URp46mCGRBP9dYpNLNATojYXvARlxKggB49BEZECIvNjZbi5c4ohWJTVPWYTOpGauQV1UHjML
ZXcFOMgB4bvE2+Qrqd2r+5+UfPNbHxBf7jVTwmycaQeLZv2/SyoYDax5lTSqBsqrwp1bOktWNnlk
lWFu+jiZhw6tXrsHGoTB8rAj4bJqfG4qhW9Qvw+D/jGZv2wG2gCueRdLOntJsxQjvWdKm57lxDxD
ubwWAgtn+Ta+sj0ZPjJz0ndoRp1Z5AYE8z4SJrnt9CP48CUeQ1UCQnLXStlPHkRdUH3h9eXiK44P
epufaGGmH6gxxwzr5tJeKS7VoRWIGAQ22Ium/iCWRhi3td/UlLsfZ29mXXnVzaYrpHkoSdojPUiF
vbXdlpN/xX1xC1lZ8xWUCtGQNWheSzkcVqHEgYdDpFlQqK2eBci5VsKeyvKw76h3OmEG0Ln5W8Ei
g32eKfX6MSzWJyJlRxqAz1qafOv6ZSdKjpiqYByP3r720AxQc8LaLye1OosGecv/kQuEFMKxrfpR
ColugKfeXu4O8bYJFWkpSbSCVP0UM1jxBa1TaHm3hATu8Ou29dbQ49qscAukNVeouBTsJVaO9stZ
FI2bDOECChJsTASIFj9ekwllyYsRrKk8W1fM+ZAQ+xDAwCqLLkCfsvpjW0VSHrhfufhgpE1kDurj
kR0Y7M/95QOBAWKmAJKB8UDBEciMr9JVsp6mJZgMC+WYi/vaVUjTLDG6ImY2jeLT7nxCizEdXGCD
DXEchleSkQHwwhf/F55wUrUgiEygP7sKhLeBDOEjn284kmOzX6u5sAmn7r7yjLZ8w2BTNxsWAoD/
Cc+R3dT/kPA7YWEUL8ur0WIFesiTuXZbWaWo/0AJQTR3x3uVIoB0pKjit7+NRMXf81lgL0QQabSQ
A8RYQhu6HtpqMGHEYmXLtMdqTEW0apzgl2D6Wqa3xM3IucyL/h5kzwRdRMB/rFTwro+0ttsPAV8V
S5Il9Xa1yua1xNBcsS0MasSBym/QRY3cl2GHJ6b9khZeukQ0WmFUWeqlAApoxXnvZsQhZqS6iEHC
z/wD7MBASUWHxtD0YrA+YZs7Mp33tLgJUJF9Yg2fffIZTiwePO53rjYpEFADaK1Iu6rmwISddJLa
EvFpIzIbhJGRirJAWtLC3aDTfBCTQ4plFw6rPZDAmaEJW+h5qn3LF16wVsM1uXfCuUHoyPJg4gEc
k0/Yo3MJrXIaWTrFfIL80UT6O/iUEtOQGYtiVOD4OCCPKy1cf5c0TQ8BlyNiRS0Uno2GKQeTquYK
ugpqKEtT4FsJcd6xUn1w65O5nwxZt80TJrjB8KAhz7FvBgW7KlfBtjkgSVVRm1w2SD3JtJzbF2eV
WO7aqOl/Loz5BsWGUHziC4SmZ0cvEBELcHD4x0PQYlMHpBph2cHOAOMKgH2uqIpMfMXM9C56EyFc
MejLX8k9PTTC9Tmq1AMe1oXtkGx5LP2Y0f2jOpbcJaVk/rWmxvAhVAjM7g1MKuUVuTt5ZbapX5pg
A6znJB4viblgNC3wl3X0AkuZ57C49D7YTE0/nYoC5FVyjlWz3V7RPn5QrbC+Qax3w84YOmGgzr6g
DIVT65oBQmV6xxKI5p5DZX57/gwPnrdzy0dbvKlpfbDRLfALpkKHqXRcuKZgIiwjihvXpUcUBNdB
p8illvkcPx21v177dCyfnpsDB6b4DTV/0ELXZloZSkrsGhmSo3ewtOnVI9mJAuFfJTKyvq0Z9p3u
qNlNFIau/ZHomdrVyHGOuDqurV9DeRSRvxzy5yQpveS/eh9ZtX04XAQOK8shsFI9p2/TmyQ8bgPg
6dhNi8yF/LJGP5Ek5BtBey0HMiIZ74dgmfEXIKT2uJkLe1f6/rZdas8X4zyvhMKFIBLWNHUGz2WD
Hhlt0MN86NHfIlKT07lI7UR/PeB9KhdzMw5wX8qdb3U5cM5fIQyQ0D3AqikZG/fmNHNiYJTslyre
RhlXPAh9MAT3pMJoYQJh31wx9vKMh/osoqnIMZuzou8fU1TxQtHJOjkhek3XxF8GW+ypptNk7ryc
bsl0mDHRR12YD8aaZMgERIpJwFCdcAoVX2klCEupRm+NOiUjAXYlDlhGigLUGdbqLExIs0BcUkXh
+jB6VBA6y651UBhWv/dIdATnue/Iy3nPOHMLMkXEa136qPybAR4gvKmneobYAly9AVj/3GCqh9Ug
hITKDeABXDH/MSMKrdx3f9v7x1tuOeFIuQEeVIRFT0PzypOXetnTD+RQHpYfFwwmJWY9hBdVE7ed
9F3RHToUHb/KMM7zhTit803K7GtI+7ndhSjdn+Hv1xHcy1xitHemFQbh1akmUGGoFXVcYH78oZNr
zKBEDkm3AXMhgWZG9D9gZkb8Abkd+dvsWHKnkokLbVX9uBcIrLQMbM9hH8NH8pbS9slPlZ+p/N3b
PtFaBBs8u/tsOdJ7anAA+pB/aHrfHZSAbtPVVZX5WEnoQmHlmWAobhlkGoW2wJYwXuPam30js33/
K2FvI3o7Zc2vAKY3bRIE064SFnoNHlMZq4qOecSxmEiQH0/a//d1F3D7r7twB0xT4z00l6htBMd/
p2r1GBe51eDbycyvNUHbGMkoWbs6ZHeX3xKHxurYMd2Ob3rOARcKKmTKt4fWygncwXOXJacfg2B1
Xs/ydhl29Hl88zbM51bf8sTz88BuTsstfb2//snu9ZC4ZZRoEYxoMX9mXANDmlTx2DEXdsVHwXlv
e9w7n1ppLFR+bUWGb/D5FZ4u0KY6NdjiDq1bTWp2rv/DOgJrpm6wUchfvgQBOWQhP7zjJ6kh79Ov
3EaLoMVSxqGBQ29JYvbC/RAr/e8tDUmx8SgldpAqdKytuHVLnFMiMklKAZP+i88FLWnUvURPbu7n
28QfB+Z+JSY05f/W2fSPZ0kmUDcwgHVpyLv6E29RYfcG5TpBwWtMdGjX9rZGANeGNDz8F7RsUpCM
2EXvuWVjFToDKRwjuSIyYjgRhNaejlU1ZUaIAgP7UlOGJfUSZC3UfbY1Dm7k/yrN2Ng7tptrHw9Z
MiTdaibITSAkKZ/EW6FooQFrO4WYXxy/aYRvv2QYkZzugjqDvjUF4XVZRWOmoCKfeXX61cxoP4pN
SmeyjPTz8CZkDtg12BkIFoipq+/4Te9azsQ2ugbFD+V8iKNCd3pstiuOQc6E5ut3S+bD9D04+BNV
m+bSnI6Jx56swRvv9CI1FHpn89AO/mi/WFqZ0AMEMfMZBKR/nxlmbqmaf6nL1deH7YTPHWhjxjh/
Hs2JabyclVHL1hDt2WtS1vaYPBxJLRPknfRidANi6h46GLhmfLbGiS9EroXurpJB4k1c2IiJAgfY
STo1VEXAH1sToozD0c1NzLcGl1EP7Kvq/z/aDE3tgv5b0hXfbjPS445w5JYWsvZ+wI7hknfm8KTw
NOt+8sL2WTSZROFMvNXqF0kS2q6iF69zwdFC3Bizfu4MBUvU7QdV0+fAzblKFYMQeZz4RIHoJR6W
9TJDcSprFXDDXjS2GfKty96Uc6SQfELtbyl7/IN5ekHMAzyT1vI5Cr9HPZk6BT9zwQN5N9Z8mEhF
E3x7bNZ9cYnmWTFSWhP+WINsn86d532NJEtxytZ7/6sp1q0WLDYu01Qnk4R1a4Sf9iPHDpqZfWCI
F5kS/j/YSMMqpHwRRUqz+0P9hjYqohWaNrqVlDOn04w+8TB9q6nreO1XdFeCi5ET50eRhEcjYmtX
2EgrGBHve0hZoy58BRZxYjyAX130wbQY3ZVOM0VYTIspX9z2OMbXvqsupvANI3NApXGoG0d733UW
3qSZo9iulePk1lF6ZFuQYqZtsUh87aLKnSleA6d56fevYi+UfmEDh0FCZPl2xhmbf73zDiVi71o4
akxOCx4F1nTBvYBZ45nwSv08M/u1z2ZSoTC+goP+ZZtbZ7d3qV8u4qN/4O3ZWktgpis787TvKXNd
P8EiPl5LwjXBACcq2mUj4rICur4eoXhF1m6JkOAwN5aY/vLP/SSl5k9/SDyCFimNYYS8sgGS1Qcn
cdlCVXjGsR2ftiQpI4C7PifC3ijS6sq8uNOWRNtlt0XCQ2/1nbVYC4ojlUSJIuw8NAA4mA8MAGTz
f4ggeRVanT9Eq8iqGPt6A1VE1G7LiexYLr5OeP180X/nmc616aYRCDaSzwjf5qvvSE+QTlagMNoB
FQE86GcIYXzAGpIcKQp5jRpz/gSocvDmuBFTTYc0Aw8duRHOtQhgA3ajYXYCkAyNYyUSUNAOYjw9
nfE8IWeYTMWvqUyN6l9+6selBLcDYHE34G7WgSUQJ6yTQjgoIiF+qLiztCV28y8o4vOJg5nKJUZZ
Dwfm+/rAt+g6mW9m+81XzTqV9NSNsdtV4g0ulxNR/PBLvkj6c0sjBNsUrAosnOGKCMPw9fYzlOSg
Ts8De3wB9HaHzABYVyUv9mQsHw94RZYUcn8c/Me1OUZPnSdo1t0dbKwYmgpL1zvdGOg3TLgaRRWk
upv5YRbNVM5jdZDrMiRTlfBzqPZ4cMxPINBsgDDdYGj2pO+zBgtv+H0UoRMkCItT7cT8wzRvmdm9
92s+jtaT33b7GBWcsCeDuXcgrXrfZwYHiKUKaY2X7NV188qjkDjKzFODVWbOMX9oma3wxB/narjK
OsMz6MgcUpDLXm9tSGYJc3Hr9/2C9A4/opgMKBYmkH4jVhpEsLFUZOqeXvhLrgjEa3/+vYKtfcg8
tgVuiRJ+fZ5HqIragXsTW1KHl1l0GNHxysksrDQyM6kV/CIdjUOen8Ysgpx9pjT3ouWKCm0VlY7f
SNC58qOIjoVGM4q/OvnhSNKQ9gdUqgNER0B1D2a+xM1ouo8JGBpVXdZZ3z41RuZW2lYlcmqVIjBT
tWel0Ssh4FNyuK2F7mOwf8OTHZALVqqLYfeTtUiZFgka/F3juWTzRpW5CCCMv6NgK1E/MTFApzNc
ntSJeWnxSCcwvFxRuWjRfnWOKNNYcEGE6M7ea5BQyUngDE2UUOwW08ii6emZJUG5iBm69NLEDiNz
jTfqI+yzO/ImTr1XGM1PbMIEkzzKLjCKdeFXXzT7Ui8B9qUHP/c041eLulpbvl/RvN3Y+Z8pAucC
ddzR3QGFRNpLTbd18m2Upg6TL5gHtgUlgyHeX93JgEKNXR7hz9a0aZwnbhDF8EjT0SlTUFObANkR
1x55/+EhRXlrTa5pHYEc5RLaDCEfCB0lcPR/UCtDWWWI4RUac00XCxU+XRrCpHUB9fEqmrET0SEi
3/nC50LCJec0ez8D6qBthiJUfFJaniUWYS1zC9Ukj3TO47ZsPkBaq25rCesdVZ3gejtO5oKctyn9
BAt4/UFoxq0q1DQSeLN1oY4juQoB2YWu7rbGAU9wq41K/ecsC8vZo0dDsIAtq/WpLGVm7/7yq8/t
22VJOo62vQ5URB+UiQfIbelVgxF0Hslrow+Ccf/iLLrBItMVOCrtWmJkIW20W5falSAP2XBR381g
M106DT/bgGxRA3MamPsuVJOr0adAPXp0PIM1iNf6UxrdKX4xbTu4OmccMC07lP37SiFeiy49lHZU
AoU29VprBXP9WL0BF7Au79QrrYQjtiUU9mPyuNAAw9Vu6mTXf799ApcpG26A+vdh2IJay8sMEuqa
EUOOBZO+wMRYsoSEXVPXyFTLvgKPzrOzYlH8l3mkzoKcABAzHanHzFdBAhLb1zNvuxbavmvQ4iEP
4SDeSlkEepZ6SclZMs+8o4arTwusiBgf67UCxW33A4JVnjNw/hNFRPMXDfw5CoyNGzrUq2ci7z4s
09OXNzPCg/rL7uBQrJfPTDYxcz5nwsFkjS676SevJ3TeAgsvEzuExof4HFH7UENZwW1/5uMyL04X
PI/mKWztQ1BTrNa/cqwEDxqNW5lkvdZqUxjoHAEWsuMXetd8NiqFCJ+6rYTh11aDomNgvqA5ZkD/
Hev1HrnE7clz5PJn3mM2AQ6RxuWLGJCbPN4MqWxONVldXH4OvjUnV2G0LIGc3xt0yyPvgXj+lJJ6
ykcqM1qf0XuPtlKok9jVi89+uU6Ja3Hif5tQq9LT6ucZV6qhKf1dTTqn+5XfsJInIm8NY2YK9IDe
NeLoB88czW944c3pofvqj4qEJew6Jxgr/nNelWq7a6kx9Rnya/Z4EW6Qwlcv+lsALKKNTSm5M5AJ
0g8PZ+Dl5xQGKigNcHTvbw1v8+kChwce6dQDeOM2m3AOF1B1AinbOucLK2mpNIRCbTSztv+acJYx
XLoldSE92ZtaKdvHmqKFBks+7KQYqAMJcrvv/ptZWf5yXx3OmWx04RhESms8YWgCbD/WsM+EyJi3
1qGw4Zdmps7YYunildtLeXG+AhzvoisII9NsqUlW8wRZsGQ9d1cbi8IQfQHyNRwy8Wlp+jPQC5xk
fJK2IvvCZcEEkm8jVKpKqrwAA6bywD3cpmKQIp38U11PM3bU1JFM1HUv4Rb5M+Rn6c2ESTgtjT7U
wxNNJGteciMEwY7BrtiejihfTSahIfNK81j/YiYdtlaDNeydwpG0gx43YxzjYu0ZSsK/EGoySd/6
drViyukCa9fRCFQkyjpSj8H1693Wau5rB2/frwcf2KIUIujN+gz3G180aq9wGHcq5W9feo4vV/6z
aDZLD8yOloYc92FiIdPX9YVNrFkPmU5Fg7PaVL+IPdsCL26Ao2OhOwZATeDhP19AT21GjdAVRpuX
UkxE8xhGNmZkNm2M8AQeN8JoJWyjPWsuB/vWXA4Ayg8Q6hRBhZFSlT+yThXpZZLE5PJqkxTin7q0
8nay7bSIdRTHmdz4k24roHchSwXBFRDGpq7hQmxSNg/O8MfGJWSFW+rT7zzb2cQc4x+4wq8adX8g
6s1e0JaeP5I5PidWb8q4yB49mydItCFoCF0Kl2XGeco77xi0THRt67qfmX/1D64nL0OH/whtwy8W
FYd3Ne1+nFLELA3N3PHGH2Jz1jHllQkY347NJtY2lo7XwtuwpgrSwvbygf6NrqdwbjhQKl5WlgwR
RiVKjo5PWvlgGIl1rvoFF5mn+3uUg0mqG56GbxnLyhpRUnZS7B/3B390I7Rf0NCh2fvfu7WzeVhY
QK/Cdblgq2BvnTkuHTYuFSeclhukFyM1TZOb/izBeC5NUM1RXTWQle8oRIVo41j1yOHNwX/+K1We
aeDR7k/8RFzIwoB9zAnopIn2YJa0q8lWV1kNUVfkWZFjl/0XaGq7U+zpBq/zd6JRD3vL3aWIb9UN
3J5ZX2fIatSYRltm3e0jHCrjYQgtn3E7aETTQ/OevQd+gHtSKoKLcNcvuTUEjyn5rc9m6xTBEHmx
48g+Irhm1hp8i/0Y+uqmxTwaNkLxItUwFVFF3BnHh8OK7U81lLc7efw8E7nz0oYEmU37TwsDEGmn
ZJUiSeqhPUSUWsrYEoMF0s2LHclvbJkOt7fdLtkmtGkA0puq4FtsqnJhYi8YQnYzgK6Np0VHPDY1
A8vcfQGbMMMIUkji4enI0TwWhGOWsFIfKruV9V6ld8uhFm+fZGzHFmx6Ehx+XEX7+Fw9Ma4kJ/c1
03OexqyvKWcCVkGVRfI5ldgC3WlbWVhMLkF6qxvYU0qomEA/peOU5pSxd8KHdHzuiq+rpwEgKiv8
Dh+az1s15NtBaVf9J8dBnLK+ojs5r23sYcl6ccUl/4tfRwIYwF7jTk7kFdS8aTol1gXfFkYpbwau
YZqQebmGz+DNYYUU2jR44lQqFH+KChLv49sMksTvlXXMP5yGiZt5SfD8j3zR8Nvain8/gRrZ7g+c
osGIq5vYS2lYhg/yx4RMsZ4x95swP60ukNsCW4SdDWQfZlaWH5eG7G/HQm3g+otKXyJtnvmN+QQW
xXzrXRzHylCj0Bv1gEVMDXiZEru9oQG5yV7QC7J/rlIrDBHu3E7s35Ecy3opPKFxM+72XImCh1rU
yjy48xvFx8jyPhXZ8hFKl17JX/XXCogbG/l44RHMNSxpxcd6w3cWzZkI/5GVea2jRyJGvtG4R6T5
HVoda1BnPt7V5PRbiKnp3VswH5LRJ8Ytzvv0q3kdMHGp6J24mcUAjOfw+dnsq50Q7AT9ODlgTbn6
t14JnTHvNp1k7l+BG7VxsNE5H7Bbm6n45lb9r9zKlVuZZwQcUkesXK9mRGze7GVbv9ZfEKjde5y0
uXgSh+uQxlWkgWF5NSuEfvYI6cXCkR8h1fdbkFLXVsgI+JAjIlF3ULyJdMGrOuWlwM9qamzqUTF0
MGgCHGWBP/POH2PZlHLq3hJf2YmMKVyZDxdGsW4v8EvlcM5sLBOJTQzcqRF2gEysu5Z6yqdrvRIi
ntdEA34ocX5Gm2RmrfdyKYsP8NVyaACVOZ/fDrKzNmvUZxTpQR8kms6FCVloFaxuHL8xiYXU2+Yc
rHHb52DgH7jCLmHx9rvmiNC6verEJoLSlF26P7+78MuaFqZzb54+Tm2TVt1YSk8ibRZ30ngF4RW6
1Yn6c5KE4RzjmdHpWWzCyjeOUUjcRU0EjB4FRMsdx7Im6ykIXzFvLNJR8scrUzBGfaVikOn9PqLz
Q9SU0qTT6avEL8phBIjJHh3kW3P0o2XSQ61BO/25Po1lR69ZtrNZS08lOkUJK6Ypd20QBV/N2/Uu
PJznon+xH9Q0jCE10yC09OlqHXPI7BYJ45ok1EIR8uSNPq3YJCjuIekeaDqEQQb1WCjBRS3VY47R
7IptysCUmzVa2RXkLsQzak5wWx/qrzvPctMsV1YQn2x8WbSgPkja+6zsZqxRhBegHf91Imy/26wV
SNutTd4zXYFu9uFe00AYXmtAXHOGiCNAiA7byfy+02kAfVMw3+8Kj19kF1eduD1cKYeIfA8eGRPO
fkaK3rNrYMOUzhSjGRRFZkjvUTAd2/rvLby0WurWCFL1niE47Pv/P3uOUpC88PD54yDKuMQwlNXu
u79ip09LUkpn9aqMNq8J2agPm2/tLe7pyXSu7jVlN9y8x9N2RmMDU7bzRvPcJdFG7ao9oO9wK/9Q
WH3kny+IN2Cnfp7rVb56Zc9BHmggbaKimFi5lPVTxqhMKdDTn8awEvhr1jprbfwSDBIlK2lQtrtS
Rc+tOV3hnXPTIR+v3A84SFMbotIffmaDFtgbweFDCFzH+P6xY8R+YFggEd5+MFWY0b09QlZDWzcc
K6I8v4XiIHot/tagpLwESI3RMX4ycaZWeys2RTGPKagC+g/e6x0Zu7WaPzZxZAPlr4XFRavDYqP2
H00AxN14tPQY4bvbmWgKL4AgkkiAS2J3LJyGmCoDqEa4IEqwrYs2LK+nwh8JbQZn0ZoTisfBqBx0
js46D4++bKFq4qjpaofoBd3lE+LG8duyC3+JfSX8Hbp95DBx4nhvOBaaEM7Ixp7z9sWnKAsI1Iln
qEGD23UC2Ftc/5WCwu1jJWFEiMj4hgoNZ3SatgIDAixHwcUS8GNMranCJ6FAa7LDXuTz43UE4jq3
vgrLspV0b1GZox05oCsXmMtfw/pPty1T3LuBds0ri2eSqKDyj/wJAUh/yeRTNUIrwgPppCytHKt6
62GllxUEXAaL4jZZHujwBVGrzxZj+qaYfc9LyXjgUVhRPcq0v9EGA7uZN/yQuCLmTnmIO85vpSaC
6prCu49o2eNUCDB/B0UG/z5jWIdC+UFU08v5OLCaAVeFi1Hehpz78UX/OSfTe86mSjQjRAPn5ARY
ARB/T+ayhQCyEm/pZ1o+YHmlQAb7YJakTi8UTktcXCZiQB1cGRlJ7I+h5XU1QOJC1Kc27E9HGxtp
yqAQt1A+q60lyawsclB42LHhLPE/gh3OrktkjVoXSCMESavh59AapDOPSLRWYWiy+rGNyGXyZ7RG
ACSzhC2B+mkjNm/mtWDSoqLjGkVz06cZ/UxVmWNDFOWygUQ2njxW+jn547fw4qcN74aD3/UUcVIr
b3Y7bRg+rnThu5HVxlmLuw/XxVyRYRk1gAvRs132uGmnqJ9illbrUB8mdMBjdLU66XjTIMhn1ISA
w6uHaN1/A+bemYPb4BmJNHSsMm9vckWpNElMFp/T8YDmeSjZ+I6h70ltx7MOEZP2wooKdje2L5v2
c7OZ7kZReGaU6QRz1iQJx24+2VEBDE5ygSVJmqhJ1YM0Tb/cZYQA7aGh8edlCAMAPm0/SVbHDSy8
WW5XbxCRrPnbRe+WDordkaGGFKRGI9RORDKO0Yxq0FRFCpMWRbr4i8MRGGxURHw/ZesrtxcFEmVo
zwzxDRoqY5sj3E6/s6XDBoZ8m+e6bulioNolB5Hn/C66T8mrrHLhMakNzUjvEzFixs+dDuOfNcvb
OsYH3yc+abfXjTNh9591GyHWDSPKgtKBaT8aBKzns0p38nqsV2eNHxpnZQ/A0hJf7hL/Adwb8dHx
6T4QslLlrx9BG120H5W3vRKt/06D/dtQIyoWyL4Lh+ziBCB6iyaGz+qmAsEnhaHokGXJcdftXFTy
olJXBM1slF95Z7f9gjXk85QePYYtWuUIwwffYzJg03Nr2BBwM5NOsYNsrYBDYSBtTbFANLQMPdeB
EXvZh28rZpKVfO6NyMB0hWUyjpjm6VoC787K56LR4gGUyu6A3uQ+ekReopcLlRBWTKetOXGtyKny
8OmmLtrU2wz5skuoT3RKTlr98WIs+N1kynhJqnAxDd1lbWovRwIczrEpFrBZRnGC1N/YLXq3K+Y4
vhUWIaH/RcrxdXDRcDSrNErw+86dnO+QVddixavEobEBGqH+f9pVAe8WDdadrcDK9Hq04DRf8cFb
57jMeCJSSADghtmEUcOxRkY56rxj6sTfkdXjXmN0U5ypXf6yARrmAQGMm95fjeyYkPuMLNICPw0J
19QY+AJ9hKUJwMTl7SsH0JHFPDmOzlN4oGIAzOgGPlnQPyyVHs3evhixKTiFqiP6JBfGSWpw6Aw0
RXSnG9lOPZpJiu3eMiceXBVQurFHG8/UPh8eOz/L9PcPgttEhQi6KYxwq+Ohz84tsv9O1EJJxYrr
oBXYJEA/m7wTrPT5Ar+Ud4Nw4fIf1I2m5XMuBWko1oTfXnC2+BVrTls8MLzS5vfTei7hU5bkATYT
Li+/e8U9g0qsxzQGmEQEOtPFEH5gNZrcKIMksWyZQcDfUF/AhEaHQegncSSarC+q2gWqG262o/Vn
cKBZP4GQ2jZloeTY0xkwyce0jnRbpymF/o1Z9R17OJQOuX33EgRtNQJ9XisoKalcAot0iVqVO9ub
bnh4cpsq0wa9NpRctgP+m9yqKmkpc38AqPcgGyY5JWjhcUiNKKRazMjITPNiudvOe68fGze87KiI
JDKKIyHX5SsfyNzhnAiSLyHxn5Fz+VRq5qdZC70lhr7V40zzMTeY4n9cocJwav036fplqYBzsiS/
RqqU3wQqJjIpmYGq3ucNj4INbJ2GTwB4RFu96MHCF5XUvaoEzkAsdKcnAUbjtNeAa6CTJpvAF5M1
jdj6lKp1LQRxWXKSlPOx7ZdYk3+gQaqjh3MT98n0eMK3p3MCXSeh0dWKEeSvyNckKKwpf/PGMm1n
iR5c1ncMLJMKBUkTTEaRABZhSTHSPsZIbY7imL9DBWYlWDtD91S8wboKjB2ITRr05AEx6HR9q4JF
1J4ZSAs0QqUpJ15a5+YoUfQ1vxJ5I4tRFdwIvW0jDHsQ8jZf46fcAJwjrD2wm6JuuYYdmOPezGEX
hG1xZvKsXzTXzUV673qKKP9J5IcE/TMftiIIbkl5SrurHDEJNHXgWBjPNBKvz2esXMKlzbic2ne6
lNfnRfBMDW2PDswDP2wzjtTwGRxMLhQ5/2JNd6tMdFO2esH/D32WaBKxBjLMKY11jCV+ZFqRs0wW
ebTXDg2w9NY+UuvqMr1OWWOfJYAfcptDMxqykGtkJiEZH4qWaaWUL5m9XmeSMzBQXIHK+nfFo+V7
ASAeKQJcclO1UmXaykSOiejFSIC9yPQxWrqVBJP5U/fnZSH/4xq5QsR6C7MLyX/lVXqvrcwA4upz
SB349bQWCgWvjvXStOeUMEcuGoaw9JdQGFhg3mLrRVWDlXGpkzR2ydDbf2eZwcTpY2OgWSGWM23S
mSBg2OS7eHsMUo7DISSPrRSroYLZyCn8GHfDJD+nb4ktFctdueIdC89oyTCZvHV4YQTrVjKFP/hP
qpOWUwph25Pm13TE5Oi8Kd/asf9q/gNEp2/dtunejj8YuIE2tWSxy+uwkM8lUW2vuA9BytJt9euf
nmUV5SFfzTLwqKfQdisYq/7h/NOnRXVwYZF2XIeqEoEtHfTZNuoRvRoUPgd9MykqJgF/LZYwe/2V
VLwshyHeTP3bSHba0W0rlsWTMWXc+gJopLGWw72IiB1JfAtOVOY76D5YvAM16J1IrAEVKhAWokXx
otbPNropAE4VJxJsLGjxDVQIHA9a0ldCPoK99LmKmI1gSFGMCuQjNns2wF7pShcDSWLH91A19BMO
CmSLZUuWMxg0xaFiUT51ot6MapxJO8r4kDDUovz1fQEXz67DW93q6AGiJDiNgcVmJ4DK6mRW7c3F
Mxi6Qpb9D5ffzwctGUJXaboQ/tfZqJ6b8Xa5IUoDc4FeJMCxbFznk5U+7Gcl9aVdBXRrf+jphKrZ
LGnvRYAuEtwYwgQDjvOBU5cUvmhm2uCyX1wepMlj9W4dmD0TZr7J1T+Az3rps7JSpYXGtX5BR9JP
31/alwbASx3kcEdK+4hDsKr85SxqwODjm5Rcp80iqSKdpxo61XMKA5YlV+NQs2Gg80eBvUisagPN
EDxUmLdKOa5hfg7BaS/kqrU1SAmh4ko48kcShD7MMzSY6Nb8UPvWjwbkQbCODxY5zYqpH4J594J2
M/vL7dkoGq8gTnWvGVQ7DW3lPNHadixF755y9aIaL7SIXZW04i6EXf7yFFXkYJ+OiZh4UPJK8QkS
UO25xRCUikPFxLkU9lmXNOXHE6FAKvsAB5hxgRsetSmXracrq8qLHLa5WN6PJYZ2B+UFbMLmaovp
aR463jNkndWZlUq8smiiSKAoXCymq5ARPhMU2Yz60H3yFbBi1Lkt8UCyHx8gEg8yvJyNvSPJAY/W
hszaUzjfeoGTX+EUku5asBE9aDLxU4SjIPXxs+p2ZbR04YszSeEAwbMGZlF3E0gJ6CmDkHTssOnt
pKa26TD16VAB5QRpgGwE9/gvhSnoqJ8x3NyyMC/De5W0bgciHjDh236pMjCFVP9JzXsYLxuufQb8
+P+xwIdbWHnb9VxqaYIMVLRvF+IHIArOk9BOUWxAyqoCldJT09uwgP/ty8zIJyMb+0mEkNYm7Ybq
aQi2j2tcHsW6hKE59MHQFC+Fxs4KwN+sLcLekUwdgKHwN9l7ee2z6ihKsG4K5+ZtVuuxwN2vh+oP
TOblYuX54o0JWixdPSls9RkND2khn868xgz7J+3QygMMPV2Ou3gsmppV/I3FQ7VP0jU+/uZUU64H
E0Io7TUJ/y5CACdGbUkiAP9G4NOa27orYBen9agEV8sP0cGBUpY9AN2T08qtMiQYoaHW3gbFjpmG
QKZA3e7HSqNT5Nk6Xl9DvfgHInb69fupthnHSKZjPV49+HsNWCjBrpYYuO9IalXGo5Kz2jIfeH82
zh2U19Kez6gJPjLXG456Udbhc1RF4A/RLVa2BFVZ5dcLxvInb2CiN68NxjCUU3cM/fKnrGhQ04H1
KBC+LqHwz6z/5kr+5ozTnkWXjySldKdta0Ici/Ju9HF9nYQEmrNZJcQf9xqfoDGDv1uid/iWGHE3
vGaeu6NQOqqXfmn78HA/9JdR2Q2RPJByrQtfPvYRZfOswXUI2Ly/ndYmYjF9JGe9QjYO9vW+Cm0L
cL2Xk9XqOMmV7hoUTROyICvD8nUgnDcVo0z6dAeISTWTPBVU59sK9xl5ieK8y1vsHuhUzQn4w5Sv
kdxhhqLdRd8JPTCsQ36zrtzNUpWxUlonooQykQDQ440xvizjUvPLPsbidZ82cYbOYPRAIVFBV/jv
vOBvoJW+gcDHR5VhoFhNJu/zbopOI1zwACvwqbFzVtHwTRKrVgueDC9wAIKI4SWVd2TVJxP43bG/
J2phujra+VNppj9YtFUgSufddo37qLTgPeGZT2x+28Fz2yx94jBj7Gp5zxhQ7IvWKrm/V/zX/pmt
plgzM1wBrUvsRAEaxbPF4wCM4eJSevZigSlJJiLCBN44OrfH0TDugGDj86QHHYTl+5Rwdo9Kxcsn
FcaSBaPFS38qAdhDTPI1BMFgsBIihZVbdN634V7b8JT0P1gRd2JqCyXJQjPtevXzPVbKtdE0TDlC
ymqepnoc6Ey4CLMlw1D9tsGSVo77Q+UCk17A+03oFBimSvC0lIDPmGsHjCA1Z3n7+Re4DzQPpit7
M3w/dJmXtOHJ9sN+X0E2Or1sNdxd5X2uWQ3xVQzg6o6FCcuFMyEyP8sWHKr9Qd+cvgbDbQPnzM7Y
tF4lf1kdVhYaIRhvcWExRxcP/W4sgKMrWKfjNJnYQRINcLjlaBrplxn26T6RThrx/iU/iehS7G5m
HfHMvWI/U+bKGY0xRtri2OMsiEmluarxrIzGJoLjUaMKL58oQ2SVeCOLSN5awmy8U1YiyirmbZ3k
0BlIfQFtOZybZV4pt/rX1+jblCLrRydd/OQsvpBEOve818I9uAIfflx6FXqQYbMXIzLPsg4pMrT2
c7U6JOJZKHarkN2wF0bs6eJKSxxx3by5HQPI7YtBGRgULh6jwcH7dnpHdchWAhYKeEkXKXr9T5pW
slByKlgMTjw5eUpXrWtbO043JLOGlchwXIH328DDyAKwL2RST1pAVsf+Ri8L8tJ1jrLa0U5C2dWV
3BRh5umvBEC7jAE4f1ShlIejcrtTjmi2xFw85p5iz6GUqHIt65KPXvHn05bcAwaUscmZeJ5lrrL2
90zHmgJ2TyxCMlIP19wg7ImADJMTFBVYL9KbVbCFYe/9Ba+e+OdYa3Fyy65X3rNLLxEQEVi+wgHn
XVUR4pwUiZ98gPyHksVnwcKTznIKfRmwPJ7jGO+RaJhDVyc4X5wWv7xE91LateF6ifa16z3wsVAn
U1aw+KyiTIEFtCTAWIUWjnZgikt1nO/mMny17xHnZ32ZbvlTQnoG4BpXyu4VmwMy/IL5PIO83deX
Ar/JGK16m2hBOKEQoK35xwIQZjSwKh/Ihhq79ZHSfz1reJq2hDZAg7aNp0zxeK7eJHEMSYvBoXGh
O16Gv/cU1HVULQ8bc0XLT4xAMmtIbapmESEhE0vukx4DU6IPpxPqBjrhr+cJeKsiBj9s6Mcbiu5L
Y/LOW6PsI4BEHFgO29OAVCK43j7j5pCSwvp5BtkEvMBpit+eoVWZ0lw6igliLcfaXTsB/a8+EJhU
r2+Fach0jTzvRw/UNvNjpHNIjP4fKwi5f3ZBCgNqHwRmZ3x9WEyF6yHyErtUo2JE6FO4yT+BVEH7
DzYTakWfqMK5fnPNwtljXVWKza8lSb/AeHx6ccGJKKxNhnriICtKLe30MpTKZvBByKMSpt5j4sKK
Yp/OWZrkzvh9Kfb9+fYPSkSgvzg8aXPzIK86JSivOYClnmF7DaJTgkoEPkRQ2Tc8QvF9m+cUVNhc
toiG+fSU7C2cw1OS15L/QlaJ3xebE5AmwxJKSOYWetc6CogCBrc3vfL183G/kBYIYNAWCRNGehuO
fo5Buba2waCCekwpJQ3h9xkt6PquDBn53psGw8A/bVw+SZIC71+7hLbpAKIxltPdoeNkssP8n5pk
jOCkgnnMnmtpd/dXHIKsH8DLLmu+7OUVgKNRsbcp8Hy3ZhDtRzLpOu41g3rbP53BEZWPVp0WkdFf
k3nwiXQ2Wo0OcsYTCFppfFMdDvGTeHv5kCRhgfrOpJL5xI+M5NJZyuHzCtqccM49NIABKo4ZdwDS
IhCaQWPeCRcj0ty2xoZ9bZDutO/T54DSjpQwrS2CRWz8CGBXI53cTG5iwKcnpcVknjSFD34J9iH6
NufZrL4XYcB8JSLSSOjPpaf4Gpi0C9N9FbqyTev0GYIJTcrpR9LJL3aD9lnntETDX/e+hcqWBcBm
x4Q4WX27Xir2z/mAWE/ssYmPINvVktBfxe/A+2/dSw1k0CZW1FsUq/0Q7pKxYz8TvuQ4ncClVC5n
hB2xIuaLd9u4FsJdDaOLWK2+sUHdZB44oGkJdI4rrvtv8iqsQKEbf6BstPVavbChEhiLtqSinFf4
cUXgNc7yIszUleCbB3jrRBFa+JJWj1o3X4cBMmjpLluk7XXaP9KBuuB28Tb+zIFmFdJXy4HrguWL
izQQbVj2l5PrsJuHmV4iQdeoCoEIViR5LjXYdN/FLSiDcueTJT8u7V/juARaDi6+OAKzwsol8/ir
4MXfeTEjob5xGjL8CJgL0XxYRnzSIJELIwAGfAjguGm3wttaqhu5DXhrC7rnnyaiI8BzTYJhKqbg
0YWt8HpM9YgsqNzk89Sukqs4ZgSib8HiA+bILzVy3WMlY9roYQvdjgSJ7aCqGxcuA8fa+SzazYzO
xrG9QMdK8DmCq0PrrRH7hPpnrFEos5FB4rawJsElM+v4X20E9+E7FYlecmiFbFJMBSXZN6uoi8a6
9J1nh+fvAzXVGG5cVqpQLgOPXYTwPjCyah2gYFxaBTr4lYMBtdF9vH3HS06FFMFF+bHQ/OOjwJjO
9YXhr44Mjod/9ZXdmW2jHgd0RuxBtEBTvDVTESSMQa4pHBltX+3OTbSd1UH2yc/i+eb9oHyWfGjR
Pzm70BxQ5KiWYoDSPHZuiW3CqHm4jOZhYsmONYblU+n7g4AwA5ifHhQnBSUvHBCZmoWDrBC+CuhK
+G8jTgLw6f3UhEXVp64dsD8D02/w+jOukcehHUsX5BFA7//3BvHUPiDT3XuDqwuoJiGMZChFDbq5
aCU3YRCsW7XY16iWiUa+KshxsJtbcKU+/Yl1Lxv2qK8htep3s72egTaDcJykJ/5GzjyqwxsbTmpl
AXCneVovOrUaIx6dvHYDtQzEpCy0x9LRPvbw6kW5cvqLYNBySJN+Ed1ViDtedlXN9S09Brqqyk7u
coXv0qOQWTsfWaUJ+uZ63bzStc326e7w24mPTnmgRzKOdEYQPUkNYhGIOCF3FYpWMtgM32xRUR2O
DhXfJSfSuW97iec7EBmSDlhDAu9AAYEtn5rJIsu0xSfofBxmN7N7JfGX4DA4B6k0G6lgBGul/30B
hFRLkX5+xRlj1jEGcP4HR5td5sus+WXKX+lGnA1cBeIaUis85DbabutTbWVgkqhdH+RrEBApXee9
9WUFGdKBtEiuWyVPxNJvNKam6L/dy9xIycg/l46//C0ZwD9UgJ8JCLXUv24Wutw/qz9gamkAGFcI
XfuTaqqO/FPNHgqXr813vQFizmbr1Fwh25JJky5nlN55z4VvIQPSQadaKrTnd6dnQ3NmiDZGY4Fx
P4XiSqTm5/sfR1jKHPrdHB+AunwaLPSt98Y0FlovZpQl+57PrJE+leCZxcD4pc8h0mG+S0mtcNsD
G/g7PpxkIuRLqBW4hJ7MFrmFboHY3JuRrW9xsNgbmwLCtTXNYKG6I4896E3d/vyN4Gt823kHkMLA
zPTbiwO++pCKPWfKHQY91hac13tI5jmz+SvU1VKI0aZq4QCDejUmB8uzFVCHy5fvzUFZSVp4ccAY
9WhbPn7YAST9D5X2Pk0kl/eCMB+fKR0Delj6L2uFvZFCTQW7pgh4jdP8p0T548r9ycflr9qqshDv
xs95PO1xSsIC4P4/j7LfByIjrdONabPDorfXiWHaTVPN91U62J9Y6/rjoB5Sr12fM5jQYCyYo+/K
S3CoCfGbIuEPKGxDTy0CesrqLGjLEMRwnUb3x8Vj0RE2IBnPjwccVdVKi5tnuKgBv6PRaMwzv7aR
O38I5lFaq1sLHiYkWUmLcxkHDETF18jU6Ey+wJeVswE5wPLUux/PS9+ldmRaeqGV8nCQwPhQpmam
u317/VaqqmMuKI3i91FgWFVXpVqzMv0Y7ZIEpAy3IKLwwkXZzvUPyDsT9pwjfInhLEsbOT2OL9FZ
ORMUEGtuhYfdF30LT1BYeZzdSsbLfQGPdk70/Ga7w1XubpjAujsqzVm+WCfJ+duqcZvkxTiTVoXy
4CvJg/1zTFVBLm1epq0jdhu0ED8WK7sa+ziGT13y915Tx+S3vAKWLpEH7VsxtuFrOXoD8iCFycql
sBOHYa4PRDhWQ/+UPC2yC5QnevB4m+PMeQJgq9lcKojEKDFAn3ofOGT7ZPTJ3vVsDtEmGLe7xTb3
mYUBYBTw/1Qh4qajlHFmEnr/lYp1ca/8phRIhP7Aru5V0DXQ7e4wdsFTYqDyAjWga0cWwGhCF0AO
HQtgH4Owp/FAStUy8MHLHkMj7wRA0MdjUHYIH41zZ4kOQnInOjB9/IqeuDqV1cAtKbWzWTSlDKdR
VI0AknLBzyC+kRs/eo3um53eVKSOS2yhZYOY15c18KsY3CRan1jlwBi+hAmR3Obe233IQDOnN+Eh
KDQnFM8FJaLw7tUQMrZAuywu0T8+YED73CLj1xJOt0U/R4RWycT9kEsIACq0w26YdmahpjW3Ydld
vEmZU06DeUsUhvTi79NzMIRBbjAhd5W9TUxe9N+YjsB1AtsPo3i2/YZ3ZFu3azbEXxlVndmMWiNk
w0d1yLYHMbn1exi1Z7zI1lWaH8gYV8KHYLUX2LynUHDRih+S+EwYKFEE4iYaAJhA2CfkYILRJFte
e4bicJlv2gfV9ffqYV+gbZC9ovna9yDbo4p4FDxHyz8rlkcaUn04lf7WyFipYh8XcPRspp/dyeNe
UZFrTO8IipIrsjULAZQ3KC4Wt816+7EHWChVJQpO6eWHDCzeszjCwIlI3xYEqM+4UW4iv/5MxUUm
LiYWLQrQomvChmQSqk8SZXH13S5OpnCemjtuKFimPq/9lGXPpKBWFIVYrwGakXulPwi2i5V7MoJ1
z/9St5Ylo++IxroK7WQMU+S86wlhpWEa21gvUxFmV3iI81DK8wkXrmtQQxLeSejOJYlFgAumxjWU
RjWjytoaeh47PVJLIOZgIIOV0Jyipk1NaS34BUIk6wyKg+HUcHwjdb/yFVm/z9HBoPTwHS8Agz0A
oNubpmkLVpBOEvOjIieiX/gNWEtwJu30ikyF86n0+cZ0xrJ1ChiVH2VABe77WrtO0dSh36j19Mf0
5Hyu54J0hZyi3Ho3zy/Wrf/uzXueywB3IBKAKOniKVuwIguhcpTkKL13bs0XYHxAUen6HMv72YXq
MXAKOtsvHeN5xjioW8I8blD2FsjriATIFYic0O2NsJONC3zXheqTKLz/0A8NBL9fwfalN3fHoE/7
pMVHQKAEVNnI2cP14DVXGIsOmP2lJrUPnzFrK+CayTFB/u6pa+sZptro/6sp4Lkkiw844KLBfANn
oc8tiNQD03ViRUTElZ2LWh+f16VDh8ncKswv+oHYBunAEHtQ78ggnOVKGBQJkBrVWY4H+ENhz8Xs
6uWjf++z3KEbrC2zMYLgvpQgzTCE6w1iRgH7iZpnfd5tcVUSJ6ckowTm+INKz8B8f3HytGg4QRCq
xhfhpqTg6XUGzNCCBatOwJYj9ULceysO3IyVI9dDS+UrvbDyJ1njcln4+SodV9LCMMWeyDMg00rS
5ubzAKYaeuAXN0Yi/1GILqRgJNNpMnbkS+OKzr4vqe0NaGNKT5SZFffIvK0MqhvvGzs252t63ut+
pFGHYytjXkzgGrIePR2HTP/O4bsUyhLDf1imt8r7UIuDAmTzQVFOGecA+KlT8h16nK28OiFK99l9
avZexBIjizx4lvPj84M7Q37emgRIUAG7ct+7/wAg2z1sDUmaPeyBP89jVFXi7t7ccKA2u3qgQ341
Z0Algf5lkWMowdLEAd/ADjpybed3k0DWaGLsL9shGc8YQl3OxRA1OMNru3GwUxnLgFzJGGAV1if4
WGnEwZuvnv1xgk10YQldEBP3LXn0T89Ke71SwgYwPrsnXL5gur5G415MYGLrxssWY7o8kGYOBZyn
vtYT6lzrIuUWjrQP++jRlUn5Fsf0p6HINwKHVfZ0mUyv15/jq5F0kP7tKgomjFZLaYTlXCJafqYo
Q1MjNAv8Ms4qukM2rkWmMkWKKgtsUECbsEvAg/kKk4WtYjKuPZH91T1URlQB/kddGY7mf0eMtwoN
z3NaYYucbJq5hhBAfzaE5WWY5ks76c0Ipa6Pd5DdSjNuNmqGwEkbHLGH26M2NsbVrFxW+NnMdERS
SjtHk6a44h9kB/MSGlr1vbgoXMnS33UKHeveRTjGZVFYGxLUSj2rMTK5pDRBkYChv3ZOKZk+fe+c
kSCw06O2XR4wxmCf4OmMFhbbv8vuSLwnHXM+N3/coBpvvKKfYZ4YZeMNgcLRZATiH74nqOdKLn17
wRahejvayRxIxIB2d6oxVm4+krl6prJJ6kHe01tvXO6MOaRh2zGArkNY2JB3wvuVJvTuy5kKgo+8
qfQi7JKA8gTtflULLGRJ6WhN95z1jk45Ygvm34I7l4DenAiqY+SJcDAep2TNqu83RYqbL9IMokRD
o+YdUS5G7eiowuQTj9nWX2VmgGwbtYrFWxej3S46TO90NABmNeJ+kw0fEhZZFnuXpUaZvV/bR9za
CrYE4jCht7eljanhTUTIkschSDq9YjpI/gQTxMg192ZcMPt7m0PUsS6Ue75lfE43EOCUpbAIe/bn
7sXupKhiCQ+kwINR3cdMSVn0gG4pgVlTGdoSy5KCowhaKKqOkW36x6xOXRl+1zvWnYmmVnI0wWWE
SVKrFKpu5tKY8BI3RexuGOb550csdATCx6iVA7Xy7Ld//kZgyS6AeBHPiL6lvVAX2kL01/e6dlRP
U9toTwIJliDGUIYMzydJgOs/9WJW9TfPoTPOlNE21xZSTpIxFgRqEIhKVfhiDBjITZ3/Y0baCVP7
yFHqeUN5GbrxG/pbuNOA35RuYjdWpvf66YjaYMK6CPKZ87b9x+QAgzJp4sDmGfyyd8QL6XE1J4uF
nY0vMGWieIWf52Ksfy2hmtIHmsRIGPxzW9KsOoJURAS0mPF0G2bYVR/PMzL1wv814V0tZurPZG8b
ck+tU/WX8+HS9fHWpfj9fqVhjk9WZWQyNhrSI594jTAIltWbEhAQZ/SvECPEgKFe6bwrcYl/L6St
BF/tP9plBIley+sfxduiz9/hYdGY2+/Aw51FtlVK1kzywdgz6ihdgpRA6MnXixIIpVpW0qpRuwWU
lD7rQ4K3GgfXmk0RO1jciq5l0xxZe/Bf2t65ZdKyHAFLLbWT7tX1jSYKVtRM8fLxEijxwom3q0bJ
KjtSZCDUWd4EG7BnEV7u6O0r3GfwG8mEmV/4G8AaBjLEVkXd2dEHuPAUGeSYdz+xjG1ZHpYVjhki
8p6bDFI2GffuXGH9fnO2+9F9sC3EXSPgjkYph7Mzq13bQKxF5TF2VxVU80exDgpWUQLTR0m87bzq
ujzy+YZxRsuw8Igb+qht/mVz70xbAZpcqj5ky6VnP+lE1AmqigLr+yPbveQALy1xoWqXzvbXSq/7
CRRTq58Yk65t/uOUX/krw8ictqL6Ky32zQ2zda13HuSf0s360ahoWRPG7ZZHbpAp/iIxcaFtx1c9
Nfa4hxHZi1mzTg8z33gODEIRMdhR/RmL+PbPR0QmaYgUUhP9ZgXdY160erKfV6XQL21kB94VgayB
rV3gjLL9USCqMMDzRqFtgzwmxNTTmrniiJeHkHFP7xi5qThsdJxcrp7np4Vj2tDZJ7xpLRz2Hev2
hvaG8iLjGXypXtA2cLdokCDlhuRJwzG4Kj0unEAcw4u7NyIWxXWTBppyi/07ozL3k8QcUP5Xiy8Z
qoUMici0wnlByK1lgjuGwi5xuHFj5T29kCfxdl+4oCry6hLD6ndI9SszKWBXZlrAoZ/iq15rEuqO
kr2bfJ75EXNBh4EJ7x+23AmH+yqImJPv4P03wEluZeTbHqDyu9SigGJBdRtomtwQuoMG4Ya6NJgJ
+rcca94dQ35Pb5YuTkB4WTgpmToRt3NofdQsDHvQO31+MmdbQ3aoz47AUZq1ymL/FOwU9eR5cC4A
v4ETS9yUF+a0LcJtoX3nWImHlD+4BxIbMSnuvd9tmYsIa0nFVdCgbLZylo1Y2FA/k6GxtezUtVt9
pQA6Abfnz7ESfexeDGW++MME1EaeUqqLrhCbjiGYiNCmxRh8vJZk2vw7wEONgjHgVB8FOMdidtP8
guTjIRfOBRShJ4rCBLHiRnUo5qmcHdxlzVwy2TumHflIMgWe2ET8JxVZjCRBPI3qm5lQOrFFSa3A
1ic6t2DA3x81t5M3Rds4XRfHAvVMVpj9hDupFdMirqdcFiwF4TRIrRc6qRDBBfsBLr9f7HlHzz+J
i+m2A6W652sIqpMHXv0nPSYODQSMsHHnlsRFqnz1r9ZjTTuRldWaaJQcnSIfdF4es1LNyQuuIOAx
VB2ScXD88KtWqA7jpFwBSwmAVdgXftBkA7nrkgyURV3Eg/srQ/7AXQPuMkSjaF8TF31eqwuz9Md3
U93Ke5c3ovBaIs5gbs+hGKNZ7nV1bGcwJexgrBiXf43+HZ3E3oert+RXLxiXMTAd2Zhm6GjHrnTI
2B69iG0tuzMv52LkLYHXpaYGXrHeKUxjEdIWGIln9gyrrEwBNxw7lnT79r+0vEzQIvICqemZVven
C4flad9zn51CjF7pV7Cu2oql8eye72OPud7ZtPloSLDR0Hn6AX4anE82PlOhWKMowNoKvf0S74i/
X7HKJaIC57lkXAC5zmTv060Fsc+jP4+RUlv4GACUbYdrVUaRSZjE0YzdbxVmNPL0JyKC7UmWs/uQ
h79odPOYZu99YkJsHi67pgQG04VXXMEdBsNmzEw0W2hd7it7G7zBepLqQzdnIcghun8w14TPSWpQ
dg5vsCOyQ53AZ2HF+RwPUYcvh72SXtR01zCxrqlCp2mUhTVeuvvXoW9LYfJf22y+e9H959n0VJRG
aeSskxbINojpOMMQ/GTi/9y3rb1JKKqI0Ft7A1E4VCW3ocDKk4Jn7rdQkCZwXdgaFi5dRGoIFPDb
cGDJ1xsmQOFpgm6X2wfAZxCoYWiNTCZmkWPUVxz2SBV4n77lrc+YVoTd6/mDq1B+r5RKhwae4Hu0
Ie0ZXNeowGJ+i9C6jmAGBvC9bGRzQX5RxZ37YpmKvtdinXoKlOS9k32f5Xr5g4zK3o+sfohjrWHI
sthhX1CACs+YXcQs7hxbOGL+Lk9dSlZE99/fUuMqO+iQWigyJ2/0wo/dEFxPW8H9/9uDEBJ5DULy
PWFeahfeaT/gomGhfk2Qp4DfViCHgADymPQwN1c+VQqxVzOH1/S4nAJ7sQlyOl/1WbJO7n6oByaO
ovwod0q6kc+7CFGQXrXnNXzoQrSzjyQQe3VvQ7imhixyvTVutXhMXFyV6anSsf6vIjwNGRIKlFJS
1V93zIxyRmSyQnEBYkW3leIfzJH+iwtgo/fhOlA/RMUpozHy/2RLWySlc+AxctJe6mCv8oCJiY+U
AVC4dmXyHb97i2h1kodxy6WvZHcHXdrdsoBCIkJAhLbhpEiR9E+ScnBI1JqxsYUAPwsG6ycx8x46
2sftEfbBj0d8wfi1bfd2+SAX3c4FD4QVJK94bwZe2dPVS3l62G3P5DTzEj58xROZAXWO1seqb6Gi
NesxMxER+tySbrQXvu97vUGy4TjvE1+A2XFQ1BS2uP1gvZIWmonIOkTrpk6WRhQFNRc2jWqqXB6g
vOkULHs0xuvv7NxPSc9HpQerFH94tKeCCXXuLgNvaV+a/T05iRP7dkEVYeJOqo26ctfWpjkk5EtY
Bul/gnJXt7M99z1NqQf6ngfH0WlkJp4w1chXBwOoaO5ZwrfVsjNULHt/Ydp9UhNEgKmFSYys/uLE
rUeYpixF533AFXUoR9rKFtAEDG+kHnAEw8eLJ/N1zEjbCSekiVS0iK4RPh+ZKrsPPVz7qiVBqLpK
dWerXV7O9uLhMdYljUGwXpgWcX1tEBiA9iqUTMFdQaYKU2h/Y10jdF1aEEv6ANbcs5RgJxg2uyN1
NAEGfVevGyDSZ/XjjX1ExJG1pUtecdcSbhtWfYWnqIT1daliUIdlpXcDz2oMU8Tl3Mo7MA5aoWiR
C4Ds7dpBaP/PN/ZpZz6tsC4bmz6uTR3qWe2lsKjXhlnuIUPllpu22sA5KdUF3ic0EsEDQDChFk2y
1wKwvMFKeAyI7j/uS2OtcfYBGy1aSWd+R9pvRpRiYmFkv4PenNcZ7uC44YbEal2ghQStkTHDaEnl
T9jXez8e8Uj3GKaZX03KEIHPsqOK8/h4hU62Fy+jNFMX/JNYJV6P4l94h10WLqnfp1U/6o4IXm5f
XbbvZYaioZGhb3PAnrQM8RzwJy4b5Olhjk7HxyGg2j5JSXG3CVGkQUD1g5ucAlww1LHIcqXpzApo
or1DI/Hsgf6uFo2oDkJoOs+EqMqiiNe502mhDxjN0DHW9PIgFwOC9zOp64WNAjcj/vT++bjOaSzw
nM2AV5KP72cgHw9C7UmE/GDMef6SHjWjIzLThRHChcDQQLQzQ3i74aen/cGGYHv5ZpFDTTGuhb+e
nGFowIa3s3XYbTl1j/Mngbv3lj0PAW0Y0rHt0Lo8PDmLjWajYRYKvouwN7TTXtltes3qYUoTQYWT
p8hY1PPoqeCoEs851j1wnhk/7NwLRnGH5Lb3OyOHs6XaS2T+5j2VBPLpqHp1RM5mRjh3E/gfKMji
I2vUDlxin4L8gZBKwlNR5GpwZnHR+RBs08izuhS9OR+//H74Xmx9WYfYx+kTlTAdUrULGQpwNy1f
AUSQm/06mj4pRxOuTQeNnwPCvLN2nwg8U1EC3J3jCAIfn6gCWzJxTDsmOG9kc9XW+9qc2S62hBJo
vnOCMsx3xYAEgZofc7byZpBIyb/DDDCk39p1O/53MZziYmjvFWBRZi4CKsHh5/z4W79dXNk/yZ3f
O1gfX56sTcVvBpbpIfox2luFd8nkDsYXjrBYMBm6STWR32q5/op5wLQCe1zEOk5xdfpFWb1jKc8E
xCDVh8lcGnd0yq+TB8Evm+buOW1hY8nA0QTRwte6GF0QfSgSo0k51h+mnrYSfZGe5HEfxstOeb+j
8TryYnaspfxmcueImVPtI4E1CjjajEs6k9+TNuRPPtQUMcm8svjZDdgZz24Y0rVhOP07aRnMzOO1
Bt7bwz6/6O2RUXMENZ2ko8JtkAhaK3W2vCbzVgyNvqMbc+7xB1ptncWbJLl3EK/Sp8Zt8Yvdo3Mp
UuaaefzQBfOZsXF8iyxhfgCx4QUi03As4dXxExgupKWT365cf5mYROg3AnODs3QyaFxKpaLwu4wB
X6sJt3T5M1CKmTD4r5eRj/o/Mg3PjLcwK2ohhwEuWlCG8xW4u1sJl/00UENT7Fbrrf+eFuKvuURS
DJOwJ32QAXlG4PLavr9NkvqcJhTZ7WLzv26dVj51UvFT56wrQymo3PmiDR2NPjE4Qb1k6lqI2CoT
l5TFN6flKncNKglr8s6CGO74PTT3z2n/q1Cr39YSpueFTZH/X9NvHcHhifM0Ty95ClVlUVKNqLR1
u5wOqLb6EC5kKD9RZz5DWZRhC7qOx9nc/QOXTqnh9MeKB2wTlReOFoet25vl596jHdrwCEm1GJwQ
pUryTYisduRt+EAp/G+jsRjFAJVzia63VDy9b4OhjrYJS+Iw5mLJ7R3D3z8LLZA4drhab3LlkUmz
52E2zA0GrXdEwvCprGFgenrII6+l4Ss7+n0N//WDaE88G6tuasE3ufaliwd5uAfLRA47iC3NVPkz
PBUz0ygFEJ0d5bJ0Dll1FvcL6FqULJ9qMj8DTT7Z6w7QOBZEaBjc74wxfTMf8FL7p8u9RTLQqPR1
klR/zNkDPssoenJQ5QwSkLeIT0vuI825nMRq6vVr7x1jWmCxvaVj+GLdkB1RaWxBp4yXMKBjY3Zz
7duGGEteNQgSlElH8zHIwk+Oa3SzOyWAy93I8VD/04Isivy5hccJyRYFyxcH4SQnZ6cBTyi077hA
UYbHZ/AEOtVFg+7gPH23qrw85wuNs3OcBLzllx8IOo//RvBreGNz551cKozwbGkrzqxRTR+j5nFY
TPeJtqhegHEQjvi1xjrFkviMO0v3oE3oVRColJZU+36lQTxLTaE44kHeT8r3b/vqUUhBo2dclpC2
nZjdFb0aExcJt61wBfmw+BflOumqIRYJ9N0sB+G0JtRThk2ChOrA6tYWxBFXwetjkZo9sXUjq5Lg
hsmwVFZcK3oLLOlIYZaYMAdvXtZn1CfzPlYu0LeMZpS0+n+NxZdsFxkJKenLiOqm1rWPRH/WJvqs
IlqDrkvEkSjgCreD2QOAtS2hz5irj8OCvCTjQ9abB01IULkREOvAUfxBn3UvO1hdbpXPeeK3BySo
HwSCHTO/CBWcnSzzjH/AqhJPfxV6YwdOPbACgQ9v6zbQWdWtSFPkdPcmOhXZcfEi6jY5r85ipqN7
M7j/ywHwst6UFfWMFIvq+TOWdVxe/ijRT3nRtR3hfbuZs5NuM0vKdbkE/nHReTFzptGvD+xTt7Z0
YvVZLVdNCsw7hK8ESP2uNYU4dURWE4xc/+VrkozJcKpovDGw5BQhc2IlGAd9l6824pMdOaTi15gC
OZHX5aaBRD2aVbQSHg+hpW+lrc6Jpm7EEtsYSNzSy9AO7piHS8mbKPMdHAWd2oFiFcwbrwm12FwF
yMnYWJAgCplxdCS+3S0o32L2ETJNfpChe1oUaRNG6jFcv6m2u1VitPi58Lrtv7RuhS9t4HVUFFFI
EBsow6cClW/+wXDv3jZFLnxL91Kwaoh8s7f4JehVKKvU0X2KocZzTRF9GqvKKQfolzIRkSt96A51
WuyM8Zav+kwieVpbR0Ahz2+U/bw1UAnlRRIAybAVjbGmZrTyMCVcUVhLKRmy1kkHr2YWUl3tPJLN
oHMDoOa9QIFBMV5XqS58g91UGLLdaPqEDhRvPru5Fquxp5BRSrdzQjnULF3axHrG50PP1O4S5wBN
XFlDYy6DMiNqVNwjhw4cHu7V/o6o4po6U1GMVCQRsmgsYkOA5J7qvqRevrZV1xRrMxiiQzZYS7wX
zFQChumwPB1xyGVg45N+8XczhlMsc6Ttg25VY+XBm2JSSaXhMIVqoztCrX1U8nRvNKEglrh96LHB
GCgEVj8l5CtbCVqQ+ss4Z1JjfnrIkHcTzD4ESp7nxBj4kVHpgJxOZagS/ZIQcRRkpdkpLs61nd3O
wrNPnQHVXw5TV/PHRC35tBOE4am5Xzqp0pRbF5tcg3+wn2LSsG+SbCcy2TfUyz7F/h+MCfWTwhNY
pkSW1AQQwIcRZw/Ec596Cl8kfrUDPVZD7lzKEiTf0x3M2mtcdacZo6jSKV4+m0okco3FFpUXe1PE
aAOSCLOAnt5S60IdEANb+St69JGYWnEfI/1nFFIDQPfVvjOlDnrGeGwTTmsRll2AtpMmPxI+MvOe
Evt+CSnBNQlON00ND7u7RX5X5OlkAQZQ4IJKusX/iYYQjhqPSgiToALRj9hZmxK1ELufBihlbPxa
PSJq1BF8AbR0sZFpB6HMYRTkBkon5gW8bZk8vc9y67b46vN14z/ToGxVxaciHR4ZQCydTNVMnIaE
sxiW6zAqITAS0DjW1UpSY94EJGVxDt+CFz4Pwc1iC0Rsx6kFF6wzPrafx4dkyrsIrH88Pp2pFnzr
RNxkJt1AS98ChUuHIFSc0ad3RzYHVQU5Vrz3XCmJpFhRufV1Gnp+lHz9xmUJbAlh4isjxGfg+2pJ
myZ+5v/gTag8jUGiMyM05hFtcAUPLy9NQamkIt9gU9bTy6gSehh0AaZNqbjuuiYhabnnBU1gIz7h
BN6AVnbUkZA9voZYTYqITA+qyPp8eQ8lM2p+dMI0KovcMuwhBGwwqFLzaTj7k4JG9k0d62875bgX
/5Cqa36C6XLten4x0/veWah32l0OxCRWySiVsgTv6qE1vqurqC73UUdU3WSNK1Oy8m0NPYnIYEgQ
i7X6FEXjeU4tMPQ596ntnCSCknZczMgjyBYsOcSSw/gMLzrPQZgZGyTTYTWU8tEc5HJ4jEChy9L8
zXZh41292qqrYUBMAnjDnrcD+XlOSfWBB3Z3oDaVcqNBxoPXqBBVThXQvhUdlGvocOALYfmziaED
4hSPKj0FBrBaWLLlybK5BwGDDWriRxJu/hDKgQ+TnLmzck0EXLDISoDN1pTFKViSFvlEHLokNeWv
3QVEphY0whZY7ecAHL1O3s7n8XcUFMRvjfJAp5tNbMWn9c6ROmTkQIByI/j38QB5riwMc3yBiZ1u
4ROvr4OyUvFFEOh3GXO+4XByCkVzbXup+9f2pGL1oM8GckyT7/qJyyLnKpkrlRznGtCwucG2mbvX
PXyDtOF4Nr/YvInZVFoQWfLeWAQdugfBmBVrzUXrVihLEIYlL58T04F4PO4kBlBDkQmvNCHlVxNF
xo09DXGw41UOQsrlXWRTim59NLJwL3d41kFyN9W2a5yK7VsWvPzGhBlDT9A0snefInMduYm7FuSw
++9pssCx4NbpmSMq4ozTvV9+7dbSjJZXaJY3AkKE/JBx6Z4QWa5Xoh9oa9DmP6wippVoQya8Ej70
S1niTkY7E0AqSR++AYp1W12LQ82MBhf/7MmKVpZf0PWMbv9DpCDknTtmwEFH92B+ocwaoWzHqadM
HvJ9i4N24fYKyTfLf8Y/iOt14ib8iwx65DvNHAI7E3aCPib28Kfphrya4sE+rfTGyPJLnjhuKZUa
0En1QxjCHb6QxvTeLceUHYRmiO/4bbVbUnB9oVfK8iH8SYIcowb6FRrR7iCSGNjH2c0IaOGd1WMN
wYLrfcxf4sameKSp0+HgkFeMI5SbCRIfClR/wv8qMbl2NPFql/YKO9dEE5C2KSaxIqiFFmbKjodX
p23vdPp99RCCAK635JCPK4ZuSZi10aHZBnrczqjFpTx71LwBh0sa2WGki0ineoXEizmGknWsNuOM
2a4U0Of/NC6C2GKF/NXGso7FkhjJRR3fq2JjjMpFlEBdQFk33KU6sD/+RTBAplv9jtO9fcY42NMW
1ZSXcg0k8FpbeSXhythuGVs6cB648XRPb03wsFXfanXsuR6rNpX5/BUmdKz6NvFdGpbCrVkPun7Q
+WJURlb0LesctYSEvDGK0D/yZ8Pavj4TgwDYid+cEZqzCTEmGBNzzwiDGXC1+pstXu2ZcpJCaynt
KiTgf7PUDe7pNRnIu0bB33kE4OqKsZ+H78Ms2Y0RiPNH0mHRcuGwQdnvOW66zd4OCFOOoi2B/bWl
8eRlZuVrC+qdohVVPUR9pXPGljOHDRMbowyEfb8QZ7vRr2TVpqfnBWAP/QftpjFgS7XVkb9tmAH3
fLL0hSE7Y9OwKJjc1t1CKVGI8EAWUfNv+gUPh6fOaIc1e3qa9UvqLmnJididhAL1LEOmF3DYSE5+
gcAA+/l+o01g3gbY1WRQeujXivdUL9xIYPG99tu8Qz4amO5xtLWdTrYqsmgO0sbqd9uho5Bujo41
ifu291Y2jFV9pXJB8P0Rn8UltEF+OzVXnVsUNBcaoawQ7zzo4LPs3jA5KFe6HK1+l69lyIcvWMhG
iX/piX9+uN+y+FyQLILEDQ3Et7DJxR7dwhESmkkUnrbS623PsI31/CWX316sEEF+5qFiK5dACFaU
7uRvqg2k302g/8xLy8QszcQWdWQJUSLY++734o40QSmGzGo63ro2rRJKvms+0rC0pullW7XVx+PV
mVYWaiRr098gIXdlptCytbULtR97Yh/+bqPmMSKC6PIPP7ibl/23negON3CCsPpNSNQQyVNszLKh
T7k5uHODimtZRJWqa8W0oCRKYqIsUJwqxRwTQ+XTW4jnENRNh9RvkF8uMD1v8cdbxX43Wta5foi4
WFNa7jFIRd3CapaeRaORQ7A/AykmMbhvOUTXyFFyL1tRm6J7IThH00lyOe+EpkjY1rnmazR23RiG
abt+4PI4YJ5dysIo2/+4eHqmoU+k2STUYxxkp80/8+qOegTWQG27rD7o2Bz+0HiquTbK/hb4LxJK
1N/p1KY4aWbUNGpmGGlQxgoJnIbpDb2kO7YTZxCFOQpazjGIFgMPk0BxAxaT7ThqGjOt6CzGSRJ4
oi4S9pxVrqOV1pnKqZX+GUPeotNgmTkwLcItksrT6jF9Kr2JzxVsFKheR8QfIR11EPN+Fj9sivdH
ufYOeLIsnlCAgLph6pvV+C5w0vSMLTJe5gyD81LgRwgh4+uOrhbO+vqHkY1M6NHU0wyzTxXb4eAk
pbcvzCLiSeTXcaxW9lStTe2E1Mk5rVg8K/WFF6VZ61mAD32PqV7+CzspHPo/WknYVX1B3W4voT6r
0KiRCnMG/vuodchyxyqw0317Eow0WyExWx7xbkgD3G+s+Ppna8hScn5yi5y1lsRs546eCX0FyNsb
T+pcShfCrLCWLyv/oqHgsWYoaRxye9jyX65sjCL+fBT4tsRthHp3WNDQIsCrGYKYCPOgFONmhhr1
K7tPVFuDPEQGkKirdRHglaHv+nYi5EkMjXrAqM6orTRoZDf3OPOz/mIT3FzGrTYd7zr+75k+w5MO
+Oq37ltVrwl2ub9B6x7/a9uN8F62J3BEjIWWFTdd0ZzQ1HuAsH3NxcXwAHj16wLrdWRguzEAt7Xw
ixxA1z1rC8B2C9/6VqlSmU5dQNtw5zYVXFG7Tvr7Y2tptnwvY37koACy3DFHbAplrNQbhXMynWxY
7SMm0Fy6SqU1hNufCkRbHwyNnHBbME5BsTK7kz0mjwdZ0OJGYJp6tfEe9fpO7AMNTXKjJYpXpWGQ
qF6GFJnvrmcmEezk7pVHp53W1dEhQtDsV3k3sj8mZa5nHRrZOSfVa1HIFD+y1egi5WIiCTcWsoOg
vsHHBGcHyO+sjJNFuA+nts1aMF3EWT1yU2ETORY3sQQQKHWGTsO1BAAvo3YQOv5tGXYlmtsQukkI
dmGBBMbEm2QSOWLL7Yf50rxQRKhwENto8qAmD+jAODSehBJz3Aa+AXDVQ/OVDFv29T5C1UX98v7R
ctsYK5sTd8xUDL6fohJfxpC/sURmCbC9uZlx6XnNpCK5SsGsIwr/ckZNPtJrLqYqLQp3DmNDkoCA
3MY/HH/x5Lwx+pgjBmvI/sZhu4dKVcEhnJC8y0dRxHTQ3C/rmVHK6EK5ZtRRpxxMWt5n1CP+hItO
M5SPoCsYpVygjzNRp4oPoSjBFoyTKA+NIcZIBk54EAsh6wLdIeu+cRY2GS5W5lyPTAWtvbMarA24
krk3smNtkO6tZCXfxksddTg0Beut95v/PWaNbTHGO0rgJB1ObnqPB03ErgRKiVk01phpOBDSG6cN
qxLCUUPhbM7S8O2CavCVAFGncfn0k9LNQ7weRoNDXl5ZwSyKnYkUWRiiJ+gxJmahefCvHioQ6Opk
A9zJf8WghaXDRlU8PhRMRs9sIhsMT2vnjMJ6xaz4UWJu9goxixwcAZBGLNwnbmFdWiYG4TCX4LSW
eCJ5bZkdl6uK3Cni6JHVRdnBeSthKN7T4uBId0KMfSgjmhYenYxE8X7dfh1eqUVZwXvP2djXOiF8
u7NHgRyVHJroaNHGr/AfRcIyq7pXbJJoVQkan2hmld06osOOD4z/rYaKrVv2/6uFFQWVSZrCfnG1
NgPvCYmCS8OZRjKWHejhvJrW66hrO1/mtCXSthYjfMmuH7FhZ5HOf2Ay7BFC75f3dIwCNgVTnNiP
Zjfec474AAdtDn8quSHOTWOpTpnawUQjTnHPhHRz7Di2EWQoiNxljy0i9/wkYaKv8Wa9A/UC6Omk
5vWMPGRlQ4ggIial5pA1BiR3YaBYm9cBo0cB+L7VHcPqok27aQyw3genc4NMeen5KvKBXMyx1kmV
5i+WorXBGkRTGrB+cfkKwH9JIkAMdBOlJdHYuvSPCkqUwz+VS2Gw+96TAHSyMRXy/8nFiPV2/e2h
4zJDTwiL+nxgDIxH45lMNGlX2UWFraMSoSxxWH6ErBse7bBTKXkmivxOwoNWaAXn3Eqt+IW7uZCl
Tt1IeN4dx4DrRkIyNvwMAdjOoyXdwy4BvsAmC2gf1+8sagpINRIJm5tZV7V2zFJWXW1y5PalLG45
Ch3i4efWx8L/aq98aYJ0scA5kW1WeQf9q6I6B+dpP80gVZhfcZ338EfgVIZfxF2cmGTLkwfmWvId
wr2GKvJrPkIQYZ+tITkK6OCjIPoubkITJRwQwqCX9qRcehbHkIsf3WixP8hYBCWMuIuOMtQaR1UR
F6fi13u8Hu+YmROWLRXgnE2iBhzGozy5WmBMdrqadrOsHTCtESGbXufsBZx0kL0DKj3Fj//SxXIw
mKCmRg9iWaC+XcgGwL4fivUjJJEdcGjHxqC5HnYWPvm4Qnn3QbzP5h5JVPocCRAaB661Ny+oyUFu
UelgIsv+ut/+N9bevQ2rY0CzDflqT/XUHap/8qBPI1IYR1KwXf5Zg8H7ZAbgqbxe11ECa9ftDAF2
cmgUwZ9sQFOjA2W3b1gGz/owGhE07A1RcxkleoGb/mmGFY1FoaFcykpEVpd9BBwoiLdu36nEEI8z
9B1sC9NQz3jpkdwRdcT2by/uWJAQb5YNS5vXCPBIIhiuG9ECvlS00uKx0O145xp4yXnLsBfhPyJJ
/otJW790mGbFVelbTmtVW+r4DRhc46GdLkkcs1W5R7gFSYoP/KRZLDWI6L9OKr5fx2VyEUPjlYUl
9Gg/O1d4KJJqw2IPO/QEceD4SY3wtFh5bpXi6mta9Gqq9KhJqxjRNEAQrANK/PedP4xFQkbYLwnw
mQ1a/eOnwQ+0kA1G3jRVLN+Xni6WC2swpLshHK01YBNzJV7aTcybgv45PjwsBKRnfsZPIbV6qYSI
kmFTGmwwjhAVU+sRW4tvkbCyyfFTwa3iqyUcJkOiCUjWbTOiXhXLpV5Xu3BNw780Cp9uWPmpfkIQ
AHUzW/hnwt3GjPIP+Eg8DafZSWoqz3GweM+MOv4fP5tKiMq2o97oGI7CfJnW7KZqGiMbBBja1C9N
lPOtZ6VdT0Uv3n5yROzv0TtTq2m6TRq7umzdGnYwkhlgqAdJv9ZOLDIQMjbiwNEa5/lik9JYQXlm
TATzVmT5BYXbJLR3oXKk3mQ7AUrBe3t55JMzDBw0PNTYrGlGrqELafzqQgr8yCdngEv8JTrx8a9x
FpfmcKjdgAgTnPmBTUXO9XL5Gbjt7A4oowdgtzQPR4chKgQlEeLQQuA9GiSWj8NFUxnIFiEkWxG5
Oa8vZGrtRzylWuiicT18fQapqjK1y3xE3r5iIZFwnzrmEff+qgVVuMthwhl2yI5pGkYQXjAqb842
lI360Oozk7/8PVeVIqmfQx2CyGSWlDF4yAtXdJxOl+CyqeodF4aYXlfiYnTDT8b+fn0gKVoN1lZw
0AKmWgMb17vzvACG5dTvr0BvPawkRXdG1MHqbApZqUNwT/fBwGG0oze4XMlTWEIfJxmLDcmumZmH
VjNyJ9UHtR70a1u+16VUCP91J6EQfyMiPH5b3TtKDfclp6FDIs/XcTAzLJ9PcE42/4WacTfdW6yf
Tb+J3AmKTkMFK1/xejDses92iPH6Ydxc4oPxWw5iiu5vBL80GvOgIAfY1bmqog89L1KmGDmMfXNL
9XGfm0D/YOMgKvIz08yeI7HGZIAfnDmpPTpJrQJHOlGsDFDEROX44lhXvNXpqTb8KQbWIoRCJNHX
dNnmqiVY0H6YBeJnlkHG6dttOJAvrbv1S05e+3jHZxLD8IMwgCpz60RoohRSbceHB+q4/nAs8JWz
kiDLNOaCGCEH6M7ceoyb0cIi2+Gvpg+U7FasFGigZWGMyR7PMcE2RcVZWJpJkcgumCJdQslOEYxc
MtkCfQlC3B32XN6oGLFy0ymbkvu1NVmAeWNOaLxDOlPQ0j1R7ni8nrs3sOuZt83JbGvM90gBya6h
ARdPvUp6jlILh1sBOa+TEcZn+mjXxk8zwL7gY7nvW8KI+/Qk0Qqu5QZp9ouqPDcGk+JZDkoDED44
ahIFIFHukbU3qwlb5kcvfWkYSXQTN9BeNI1Sn/bNK76KsElOrz0N2zzHyBmWALq7GLhh011ahNjj
VDR6do+iIh3teOhMyJ29b3xGybUY/50k37/85atDFWBDVk0VMWDxJo8aBDAU02kr9zTbLmIga4Zh
5xzr49axx1DJP6Woiyc/3SIwZYc0m40WWbmrCbaXjm5Jz41xNYmPCOn1nY4i+4hpSPINwoM+x9iz
niz6rr6KWluvQj4U45WkB+NT51mBkL0ScuVMYdb/bO682PS0T1KSK2ViZ/it7DTYt5M0in4jiXGy
b61JZvJjoKTHZAsThXbgnuYFCFf2/WS4nH+ij8gh1GklX7c9drWFGm6IBv632ur7S7KARgrSuCUB
GZXGZeywp+bIAHt5Po+2BF9GI9jKuwhna6tZzmUHUfWMMb98oLOA47lT9x/C9eJ5LIYt+BFmwVQG
cIqVrkipDRlG59M165PiXuzA3bTnZPBriaHqn7PCQ1ZG4JiNfYLex9MJimQ1YNn5KuN2z1BuWK5S
fmRXcCwGrWmBe/xySrmsQk/FifvZloN5w+RYlEr4O5jqT78sX4f5z+z8Tmm6ofb7YpQjLAUbmF5v
NHDxUrGSHJCH2zCmmZ+/AKawcjSVEEMWchP+m7CIbJPFpopjkV6NqYBQhz+44RNRS5Qio+XF32Zf
8XXilWojJ8qxe6/igiAk2ElkaZPzvsvedXw/CFUS7PbwmfketI2qkvL4Mygl3la0mstHJZaLRJ8R
RsG/C+cM2xQtWIzqW6i+IpAWS9EOMupV/NTpXy4sTd0EoqDPrY8r9auJ3B7gDRzmYerA5hbHOMPo
dNtAzmCOh6uX4JbLYTkwx2v6rH8BsXEhImq6EbUvuEfPcntz7UiMs7wnF/7Y3opsXzC8GSjjxXxG
j8Kqx+3q0aBJUFO9+fr3HW7ZVaUZmmkHW9ffSfrbWAwX558KnW6y3bITZfDh2TJ0s04cv2CNjzaj
61ilOwoMvdtZUyoavGA6E3ktqyp3hi1LKYYEpoZ/0ae30ycFCXiqAcluyC5Yxv4vXMXTGgGo8QA2
85qyByJcnhrIuyTnjt3acla9hoHRnve6V+rB2331en0jk+FOOT4l5O+C+NW369xcGK29KMfJy6X1
G6tRjvG9xgPs4OSMxxp5G4QvFAEUVhz79VWbpll2jR1Ug7OAMYFYS50lKQT40J8QMSAGynk7z5pa
nq1agbr2Ao+xS1JcZrp8spAyNDFEuMkimOvg7poD74/MeepPFCnwmad4HjlidjsVIreKUOhMWEWQ
tEP2TqyM/l8hLNvI9hjaJ6cfh+hRtb34leBieXNjZxACHuWc0eg8eOn0gvugg4E8qysGuVlLIqMl
ftYGdyANRkV4y30t8Nm+9rdSztal34lnE6JJPAeBctN9BUkmg1zsyob1wAgDH3qHjJZXV5X6+1Wy
YjcyPwZl01obcI6NittjifVg6xW5GP/siD6cK7nTMV36K15re7BWgjbG26a56eOtZvAPvShBmgfS
tUxy7ef3IgTJwrx6Lf6aM5szVaQtHVQHiKMnlFAB4UFpmYXEAJxeKzHpCkpuXu0BPmxDxtck6NIC
NX+h+8sv4jTsbF9vaedbvW+rdCbori+yBfC+cgUxxShtDTc9DaZ3W/wakxGCeBTeUGYvQvB5iigb
ifJV9EG3oG/VjRFmd3ZHRiGbjDQ8R5wOcSDigM9WOMWhCVcWI1LM8XFc2E03cm3stEd79WL8leE9
YheSZGBZjkMmFkuro8Bf9L/8IPU0XWu9MxjFHNimg/IK+7C3+HcoIKet1iC8Tghq8lKbTO5w+s0H
rZmRqe8zP0c3sktIwTHksXfbfADCjpFRp0mlkSM10sf/QVngwkMpMHM3jrlvHypmIE+XcfWthdUo
yDGOCHz3H0HjfxTezUGi6tyZ1qhTz0UVRoNWlO/gkCEsPcf1XtdRGGcM7vwpgdfxJBt7QcFzpbjI
a7tOWMvs8sbp4sqAAn1DueYb2P2uutFA/tTWuwmAUysWageoqf05D19YQpm4ILsWwhCbHGHdes0t
yWgE2gtdtKBGiiU2xv40+MZxkRV/imtos6IBySq0Sl7V6VzPdoznDp/oXR84jkp/9YJCvw9cQ5+x
pDlI6TU9Hd86NtCj/rREZoKs588hSM6V+NtEFWP3jBeWsXi/0LUkXcgHJEsbEGVTfOLQWzohj6lu
4cy4uIhTS3oiVPhlgn4xV1SNp+J/+DfncnIbQe1CYmSDRiSo9k23drvHavscoZWbcCricjXiWb3A
4+Qp6qvoaa1By5eXDUPA1wMJFqJxotwzm48LfoTFqTSG61Rv+UWiI872zOgEK3jFdfYVCBVXVoJ+
EylwV8Bv2+9oOe6UJE3R989BRpvYva1zUImNllmzkFAaJhQj09pDTVK/nMoHZkqoOoFbjMtWrG/b
6NULdsXsHyfiSlMW1TZkOyxeKySW0JAYyJaWXb4QRevvJqJYrg1x1GyhGbdiIZt6cZxc9P9PyXCB
NNoGvAWXAn1JTF0/7XetQLNiAp+Fce128lCLOBagXccGl7lNZ8qkgDqXxrEyOEtrenwpLbNn1r5H
Wi2q76XBlx/pjYrE9P9eysiWs/2iKyTaRX83CYEVDacn3KntGvdPL74Zp05+ScQSHhd89Wv2loHz
yCKDF0nx4YcOd4IabRkT24Xxa3nOfxpmVPJD0lpaiEoIMphRR6WQ2lGBHyuEtK1PIb5uaVGkHjLO
1wI3/eGE7Ah3lPsQbg90AOWowns9qfyLxDEYvCsxIzvMCIO5tNmGiCQAKknWfh98orrDEyUjadUr
aAybjAuqYGk+GxDb0oSbixELZe5QTyBycM83YyNKYB73TydIxE5A+OybrnJh3d5u16ppzIpr+Uo6
znPz77Z5384ptIkY3rZMFgCNkqmduYPxgbaWWiiUFRItLbM4ELNHV48u8vXS3kV2nPb0pknFdZjw
fGmEeb8phuO+fIcWs1HlRx7p25cRFLB+tb2tLtZk5UPQ42yCe36ePwaHM8fX//utwoZcwXJrnjzv
ozmZ3KH11kM6yMwd+/oTV1ZXhbq2U3f43xTLtZPBlf8k9qWKGAyuIpd4/JxrwcoL4su2/y2cVq0T
v2MzdRvr78HuPhW9wlhlJ8Ml9cPDMjRHA8h72530DyFX5GDopveetZKhzlzYXUPVeGObQg+UFBk7
CfQPVql9QEJAucdGH3F6hjm3XtlozOQMnhTutSLyRHo//ZZf/f2MSqrNcYK4/wO1SU/g39eel6yh
fH/XmsFXA64nMjW4YmOyuXCq/+3OU2VjjzleTFVJd2/IjL49oCIjLoswq90A0lqucQ+o84hTS8HG
EEdYEx6jXx6A4MLnqwt9xltCy25UId6G2TjPWhBHde215BJGrqQ4anlQary2zwgEaJpgY/udcXMa
BvjBc39dKUcMjlr7wzJelSF/GxU7T22a5qmlwK3otl1qJqWxSW+OVKe46AOsqySoAuVBM342Edoq
12f4ENYTsu9NHxTQA1DADi2reAHU0S0KNFYjEoUnIxWz+Txp1CHwNJ2fDfABiP8wReFWCJviCnnI
zv+8A6pNWWHQ43zJSMYCXt5oQKLHmV4Y4gicvbIvmB3o8cgjbRrphyA6DVD6oqQO1qixR8QHYrzZ
i5z/RTnH9t0AhPKm2E07dhbRYxfytnydbClhkiyDfruPC9vLu4flPt8yze4rzBw5J40obtEuMZkC
IRDWZvIKVnH2wbkEHy/7DkmHxWdjz/juzlVbUEkCmopQ5UaUgKeZ2TOKLFBiRbfi55pRM+gqqirY
AQ5LSVpafl0MjNjhC+yyeI4ENTH1ffXqIP2TJuhe0OtNI1+JlbDMD3WDbvmoa5LtXyuMaZmM/J6S
XVWhUb66XA+PXKlzAn6RsUlsqCfZ3tb2H6XrkaSppSltOhLlhNmDwdYYAUemSAViJ7IOEWD5f7FZ
JE/m/fc+G4kCRxQtzTSXngVPAHOyVLM6n6UdP8DPzNTB/LnyLlQKdUtWhV7PPE7Vtky2OyP8gFuO
sqO9aEzc09aykqcg0HZpUzUBjGsW12oNl7FeeJzTQvOxhEEqf1RrQAUSDRx5qYPwEIJxvvLTnjNR
Pev2zZz7sWPTLaEW1WCKuZDIeY4Cg2SxZZQqV28UwLevYd8z3ZeVPhuczS2dm0igSWkqNu3bqiSc
3b+v0U6uhq1s9433ZQZ1Ih3H4QFfFwoU/uGCPEcc46dUDELIUKXOzUXXeM8zfEAPLUPo0g51R0qW
eWC69xvxhgM0Kc06p/zi7TJqQG4EjqvM0BkrBdFR0wHs3jR9YKzcAgqP04lREP9cnP0laBMMJc1t
OoAvnSSn/Gl/77FCFhpWvfI33o5gbLXMrdjIulx76LXWQTzBYJvr+vNP/u0mV+JM/dZhM4MTc4U/
eGpB4FGQ2JIrRECCUdORfHCzLCqakf/amDwDHio1jooQ5RcsQcnZhUmpw5c9S9Q9hH1Bggbemz+F
WlcAcp4mguaFJYdhTuAHG5eBcz0zRcTmjgB0qNWb8GqL5xMGpfmg2uIsX94T3oXZYkIa9aLZshdj
tTB+ySfuNI2wziA6HdSHk92WSx7Ph1DxkKmgbItWzLmCADiYZx2g7/SrYvwABYfj1BFgHWP55lnf
ork3Fuj+Jpsdez/k82c1VCJcE6BlDagEtg7pqybfpPfZNb/Ja5weNJCDiGcxmSWOIOzUxhzsos4q
W+rZN2UZ32LId47IRj1Gaf8+NjdIbX+odP6zwQw0rer4MJ00RePS5U0VrZGN+k2yTxug3YTnivy+
jjutV9kshVYoY1VZO2KJH1uwNrCWlo+oEm4poY7fADBWxIQHZJ0vPFCUSD864ZU8jlSiksgppJcR
GnPGqU4kBsLrTKACiyacLm1bihglNsbx+by1MMV3pToC+pl3QLmSmMhnYfox/Gh/F6FnAWNO5myp
1TF984V+YVJeNn2AEprCFr4cDIUejXmVDuzQLVTqBd02gtW72/Jj2NUPNsufIRAOviryTVNQXJmF
HwpNHlCONvpo5Aslv8b7jRea61x9YwfeZSBP5fB6k2YqybC0QssRHU0i5iI2SpYsiuCqcwQLftNk
CgOxaorf7zvEdKPXACtgXG4CSUuqNrg67l34BIUhoSPu5BQZNbvghWJoBrCbnQRHVYsyLIf2zS8B
STsXlYqkqXXOctpiLkvblEgB9qlemFtrcXsVhkjyvPzhGtcyK8+3P4Kzc1InA9NSl1B8VT1HIkmu
3gJLEVWFpMznUCP34HuAEmYvhRjo+cHOWSTiiNqYd4PRX5urWIr1525mxKjDVgSPJE1xI1qceUKv
6hGNrOdaE8XOadHFf5ImUrzpqoA4pSwHICJplWEngz6KP+guyTD3bKk8Z+QjMw6bq705LIajp7Zw
A7EOeTpkFMXOaanOHL2NCQhx60AtPWt6/05pOX6C8+nIeyf5RS4BwxgC3dsQDkF2XNmeXaL4+3l8
ZoHoCm/XslIjK+Ddx+sLxL2RofOvt1E9uG7bV7tpJNW8qB6PJRMZ9/CBPQAtByuEtbs+jrHCP4PW
ZET+y0OMIMYV9Li5p8u0LgRcsRQfUptPQgnLv/QhOgnxud7eRkKLZfHOHgqD+n4EDPvh6HY3EwuK
UPwe7+UzgELU7bT/71C2uhqgbmN7QYoX3CTii4ho349r2ZjDqDadTaSHelXviTM/6wMo9JFtX8bF
TulmH3mtgW23cnGwLWKdepdWmL3Q4eJ3SRJNiGo1j3yqJSWyHCuwQAK2IL8HUAZHx+eiWw6emxK3
EeOogEQMSIbCXqAXoNs9jEfuAGprEsoRaDvDeLmuzKKdXeqGggz+gKhYCdE+HADlyyKhUFNliZa3
f74DECSh0LtjZQtyC+ezRje3cIKus/WCAncW9ig1yZDHfbK+L1aDKCPTaeNIW8UTaeg24QCENaQt
pHD/cc5m+JHj47YMtEFsL7Kuj2HPIemlB4Ij0vMGLatqNl8sbQWwglfHBN/gA3iUYgN6clENGOam
T/oxhvWHdnPyWRGIM13n+eDh/ywVP7tGEiJKXqI1S/b3MJ+h21MsP6z4p0mChE9JnUTmHQ6BZM2x
NsX5ha++IkvfuUUqsuyfCx8o5bKiRexGn9Dje5zrM58NX16IoGv4gvXBCzNZB0+O+Cb6sFcuL+AG
nXsdojmoV4nrLJKSJG+DkQqd/LXijmUmI3GJF/cS76idprQ+GyM9zFH2Ef7NgbOHcD8ZwbkFRPoe
Qg/ZOq7+D6Eoie2N3r0RsfziV2MmRXspI/qOPDU6tz0buHZxcZmetT8tj0KU7GSuPymPcTVRBoIn
gtdg+4IygCxXf2ZBtTRvFEkjRRFQCzC/DFL8OG0h4Xg7SeRfqqdYm4dqnwTmnyepMpz+COEwGVeF
q1V0yLNXAOfVHVqNqMG9fXA5xugru5nE0w9233Q2mdA09rltPK1du32YDCERhXPPC/DpDba2EuzF
ALOrmIfIRheLYhgbsHiAEDI+RjR48nG6mr35WuN4oG6doh8x0UPQr94Tmay6ufUf/Mb/ZZDcclGm
B1H+ELudEBDwpSA9M6+fE4iLI2P5YchrWjkKCA3/bqBCxsz2TG3/MxXCPShDYQ5tNAqVKnyyD8nj
Fk0w7YdrJA/Q+Uq73roxwTz0GPAky8G/hsHUkAIv6UH91lR7nnms2L20i0B/RgklYZBYtn9TIXNx
GuW/FFAGszhPKoemngQiuSvpp3PucrMe2PeJ1kLSRxj2QqsocvWCIXzJcc+YJ60BF52eVAyc2q2P
mElECDhunby35B52BFK+sXRYeVRY8mMR/MZd0NYFmR09j3ru6CyiOAyMHQNogDrP4PNu0j5KgVMo
EF2HzbhZZF9o3W+juKKZ0mfqxGiF3yH7JXws1vfpC1BDrrcd2lEM7d1kY4nJAn+5y7sPSBWI2Lbm
uVNIAE6U+MtYrYZ6+wiiKvjqz0kzOJdxvoe+Y77DOWLichhDOCvoTvvQ8VpUv5NpWXw3GO+Rrg3s
pGqY98uPWX2EsoXcWY21Ys/y65PsXS75tlflL22Vsnm0sqLhD6x4HVFYkcNCv/eXY9b0vL+GdSVD
Rt96J+I4ucKZf++YL2WY8WDJi3Jkbd475MghyGWGsBStqjc0Z4xpcnYdw9xpy+7CbynF1tAYGXTq
SZfqPjwrMhb2FmRDSx4zcM6imWtWyWxfSM66uVHtI4df4LzPGGtpxSz4EnUqVe9hDGy0YFjKkjtJ
AUOzYiFnM2UldZ0lJ206QZDrlWNj8SxgVN2fLTrVYOQH6kGnUdxkpY+ZK2GPq/KfmHrzL8BqPbjO
3zY0pIXE1crXxfKf2kErN6XfXW8Y0+wbrIwPbcS4bwG1T/AtpqRvw/YyWOmqc9bYzOE6u69/lkke
c8nK2Z+r44SbHg7XJpsK+Ks2SPHX1M6peNCS+XQC0ZYuS5X70YDTCHJkl8rlMRLJ/E7zrYiIgkvb
DXGALuAQq7Su+br0eB0Nr3J7J6/SL4blDu8jLWXlXghww9Gm1henWBG9w3dNKz8tosS3D1S7cQlA
idyEH1fn9+O6Hxb8l0Ccm3uhWJasBt+NzBOwcO66uHNPtbyQI4TfmRyKEzTdzkdrp8Ni9Qbeqkoj
OM34De1CXZ19QOwMHsO2WMNjubAvVJcXAvdB39l4fq6xIF++AQ4lUnaCD0m/SeLu5ik4mwPou38G
q49ON9yXzkSAGitvrEeuLWuaYTn9J/95nTOYMJ5Sea0oILlUb4b1VwkuaK3cPocbXPW2B+fJDY7w
LmNLyJtQIQkMfpt44W+RIS4szFvdxNPFHBZp33skuyBiskHFY+y/caUl62KMOGRt2Rde11DVWXu9
IOPJYEiY+feRDoVaYZdfeU2jO3/B3a8dNGHt8Np7ye28v8ZMk4tOCkr+Na1IX3a6wm6GBPldx3MO
GVky1Ufa1fytW5Xm7acmJM8UNE+36krCAQcFRmE4Wjgp0zWkMkYiAg9KnuAE6FBQ7bqEmMha7xUg
by8dXtfZEVIJroRqHkV1UjwBEpHNolKfAW8E6FC4fBb5CfwhNPPjjXhPbL+0YcveGGiFjIVQmNN6
VneZWBgEL2r1+9+EF6qy5qlbAvhIhNJBRs+2ijh1dw2KdtTGVK92523GQntBEOLD/qbJj7ueZRhJ
MANQCC9Vb0UWFUpIXfiUbPZYGsO1ckOD1etZAfEewwe2BeubhdQa+AqU4H3lkikIBhZDnqGFpf0c
5aBKCqA6gUmGPiMmBCcu7s9DvWacqf//6KcGM90u3Nv4tiP4FCRB4F8abOPCe6+n3TDBH2H/MNhX
7Lg3JcV6R7x2q2ClrFpBi90b+0eKRFmpD1SC54W/dCpLGjj/nnZ/l22CTi34BwalVzwAAEYbVhIK
cvxpRB1pe6Sede2GG/gGnS9F1SlzMu9h8+CBfwfD5HYRGkXRGCGS1IzrBCDarnExuf68h7DzR1/1
wHy/pyScstd6+hDqTIwHxCTFPck9swlO1x47AWiuMzwSJqStvaCAqCDkfpqsnmdksQ7oR1kk1h/b
O3DrV+dFotsNT/iWAN50paf2w79CxsOHAduRWx2oFkthZZEMn4tGCrbWeNnitrVw/e4bB/glsSTY
nSR7Zeov/UjKavb8VfeW35WxVlzeKU1O56RS64BGSTzdtk6dKN7HPR11/8rBouH2CZdoRriBBXBi
YNVYwtGsCaeXmIYxwLaxv6sYDGNfx+cXdwWHxc1Sp4K01OcFKaKCiH05qM5YKMEcoSTOozGSvAkb
6B1V1aiMimJJ6Y+5Kq4xKhFR9Ok27rcFFYBibMV04vpUBoaVJ2JDskxZPjuBSu4jwjeYggUFJLje
utVdjkYc7M7CLSBojHT3X1/VMvEINElK7Q77KpwW6bJXdSkBJshUA/w1A9tO0Wq/xY1EWKtxY8z1
NMvXzLYpR6SiVPWQcVkOz3CCJjGncucxFTanCpbhw8rfBEmfyQqT9QUMjMyOkY54g8JqaELYrMLG
d3RTVkPpZwnoybUzZaKB+zgWSFo7PrsrInXnmTzKISy7hc/+nBgrTixxlEmFjYr+vVa5mkSIlJ+I
ZjgndG5NVc7Mzdzuw7g34vZXe8XyuTMkmGpHywBAGwKE+h2uYcRArZMDlr/034Pt9OGmM0ZGr0Ht
AvT+b5r6LyWpilbuHk2KGcAGniNtc3iSUxYhl0cpdMyr9QS904zVTmR1lUEk2tg6sPZeTiOW8nnE
zwUJiisG7239/GWNEKdjF/l7Ciyavd3/ibZ4NjJNQi86BRXE5rAH1cDL5AEMZbQ9dcRUFpde2KMe
BjWSky0TU6BTs69ArdqQT7ZlxAlWNaI5BlEaTbbwNBh9gbldo8sm+7sQuClTTbNm+5GkPnSXbZ0s
JKjshWts2yF8xMnDOA37y+wPj9JqBTX7SMQoLXdV1x5ZVpYy1DmFT4ZUnfdBckLH7i9/kX8uxxcS
gyoM2IfE1wxFopW4KNry9zxjko0hDX1Fivm6CdWzY42a4I6SBwRWBDU9tmYR72AEd7mHQ0rlf6qt
E388H+jPmd336MaLrggWLNjAXc0PlhBJ0qLR3sxE8pA+Oelp/IeMon7z2JNwQiNxaZXZtj9A1zRh
51zCkug0HHxRgr6+dS3qNcpsdTOT/dZL6XUOxjsXj3jatv71hGu2LB4S882fA4Jwt5PDv5hIxhsn
ybHGBljrcahJ4vAneEzn5eXQ1q67ZqvBrBNX9gV9FVR5CpDO0QWGZGeF2287mER0z0l5sOVwf4dN
488RLRPJV03dvlgVoS9lzrkUt5By81tm9lCvYPI829AantlHezsp0NyDoTGyZgrpD+Zyy+3z6SRw
aotOh2eHCtFd+Bm/OQStKEx0VutExL3nw4HnlteumrGSLIwS4QFO3QXSX284whZqR1cJbffiBOjp
8PEcEZDFBDJ9tv0+lMsKnWzjI5ZuMEUu+f0S0RMX5qKiCFTLwcS9oTnV758k0aIrUvVwTVrTsiW9
tSFnBdP94xdh5JFb5axmmLdsRPCv03C4sTxWZy0F5xoQ66r3djuWGUceU+d4FOgkruQilp+inB/H
3uNWAqEPqvjFh/KAUwBdyUKzRu1uRwKp0u1D9fdN23LW9kqfKq1pHrH5YEdjZEvStGkeNqUsxQC0
tF6K7fuzTIjilOaNC31NyqxUbawTyUceZGBcaCvCgZGMzgVIXlBFvlebRYze71lAgGziYE3FMlIx
DmDBwuMUU0YEkNtDoiILOx39Kg2iA4l7lkXZD7znIUGKltMoULVds8/zt6+dJlTVO+yB02pKT6xN
rscPQ2dhHkcAiYzBtXQRz8SjzX1emdkKgWnh4+DF3DKdksQ3kIV0nvDNR3oKDgkLkdkM7eg5ZnwA
69t98RNLAZoXD1FsvZJnhSZo6OPaludCdR7n3QBW4F7L39e+3aF2Qx+cXVfj8jDMW5AAJzuFlUyg
l1bErdUFLn3hhCMsEGniLus7ZhqzdHzSrUJyqxFpev9BGS3iEe48h56Tekqbas+giz4Q5epO0MAY
DWaxafO5DncHZVEWHsCjkvX9Ep9L7uPDh7qpYfaPop6XcDy8uPgvFm3U3E3W7kHgzYUy2VHe2Yyp
LUDAwpszqrYcpo54mFKSv16FXoWNCTDpAz972heTYIXbwxdTkg2ShoMvFDBr9vcQ/FHqMU0tbTQ2
Lw4uoE+/6rKtMv0buYgrYDeuyeNJfYBRtgMqJ1k2iaIILF+YLR99U3UWzmBs6f2FV7HCxYnvg33J
/3utncvEaJ6rM6WA+531HHD4XPEPmKhayJxch1bR1pQTvEA313cq7bE8KRg9vZSk/ua0S+mOpjh3
KiKg7IZn5mEZfhsXzKmaJu78xgB5dMC0sZDHx+EZPfbEwH8sDBIDb25EupHoRJVpAufcY55MAiYz
+0sc75D5QHQ7a9tCQTrcV2w19CAgjYugdn7VTs7cyUj5LD+D+qBamkS0DZ3ehGcfNpiiMybbuVsO
nXhlbzWlubzlgmEzPvQnl+j98HnPql1SvcieBaKYGQVB0jrgGOGZy5DPQAPuYL6HtucWsthWdr/+
qj37PiSrG7jJ8fxpQOh6lGcZh3mgE2uDJzikmG3t3lvgbcD98k4Ti1UX53NH9VHlrUUGd1Amoh/M
e4NBgGY3cIlQ2WkxGLUVLJVuWE8Q4OZ1CgucyV3tor6GS5NGMhgvyezeZ9sUDoSkpXYt1Z7qoq/A
RIG63JwvlJprodACz401j5Y6m2ngDnPsOAx1we28p1J0OgDayQNOIBdQocCWj3I86J/yx2sDJh/z
CTsllp+/yvS85BbU3lcmyywECetDyKh0Wdtu6N8HKXlBXahb7KqIKYhvCr78ImlgD1xeLfNwbn7i
+TvEg1eua59D4zP10sCklwfJ74Uiereamr5/PLaaisxAPUph/MS+rqauMZftm2vrLIngMVvFWkZu
3iqIaobls70bxJGBxiMQkzTJZtBfWTgZPLbecpscv8tx9UGWXjyGIPQmhmuBafgb9K8fSSe7czXT
IKbKT6mK8TiHRTNGpYJ2/IO2PL+9vj6yIt+vbFTsbWz5EcIKQbxSSrP1hBVCZhHc3aydo6LKbVEi
16m/YxdocXsJSbgf7Lv/o/rIsRH+s4PFqmCvw3XwMJr6Hksqikr9n/DqdspLfkN13yloQTjawgUO
cufS3dDBy8ImIloWM+U2b+Iw8v/VbEQKuyuJQ9EEKFK70jT2gNWjP6MQ2sUzK5ueSNEuiJORMND/
bKFfDKmUmQKnytv3o3gcDvSdrXfdy5YOpI67l/oOjTIW+IKeID1FYZ6D+PopsrXafMTZNtK/2OJB
OekBrmN6KHxDYHxeTG37+HiuJzPfBh4U1AABj+ne4SRuTmqbdm9mjZv2eanHu0PPyK7THXw96OzM
y1tqUUjvqX/p7MVFFOBTf/FQ8G9jySCP8sZxrE4oy46yFINYle224NW2s8Pv1GqNiN95KyKSkTmF
tML+5gLyfY4PlImiZrT0S4Yf/rYQf3U2R+O7buPKjSGDhm5qaTay2jVW2vgr0P1xYlZbG8LnxW20
mmJe5r4EVCKyvO0j3I7VLXzFaROTaYzB45DOb4XPqnGea09xdiDz+iUBvPTEY2K2mB7wDJSFrBF+
cZ6o3X+iqOrMUmUbtXI/UlclHIHWFcxgfLqHo4gKWpNCnJsMMIa50Gvju2artj80B67bDGBVnX8c
mOhoMsVWrmzOPVqhXPxcK2pqt0mrzDJIRtOuUC5Ac6YI2lIKvXrlp+J+z3O9rmBPUwfZ+7hkN5S7
7iLJQRQYGbgFEEUIeKjPp7Dj/Eoiom046/GPlU38an9HAbgAyoXgMs6eTUhihm54Y+zHUGS1Ft+C
i8vMbmxe0pwOVWcl7897qUDvBvI5uTU1japn6S8sBV9aSp+7t2nc4digpv/Tfq86lmhhCr4eLEwk
mggFSGQgyoNz+w83zNsv/kzuj1OvaaGDMeXku56Av/sIfCcl/6nUcaXbQPvno7gIPtKqhVbgKy5K
0eOpAhq471FC511Ui7+rbCKBkaZbL682XU/aiAQrHDdMJKrDjY0Yvo/UBK5d5ndEZ1pgbj3C4DG/
qv3h8141raWafFuzLC6pZ02zMa94p+8OMVU0Czr9nNRZylMfzd96DBJ9cIOzfdwL2pBJJIQ6hLB8
qPhfcAC5iasPiII407gQPR61O2G2vpG/yD67r1zsVILl3wjZSQEJmW6qvBL9xzsx0DbaKChFi7Nx
tpcvvqkbSaBJITzMAE8mg1/wKYV8ePTlafDJplOq4dPIv4PCvCFd6UnhimPiI98iIV7fQRpiDoML
GvQCOzWwzCfO2ITEFc3PBVZiaN3O89GQBqsqEqq+hDEQX3xbPRbZwYxht84wInNMEDWGydmXakFp
tyyro9XyUDtS07A7bJmxbkn9Nm9o5SguSkc8gVqo19dKl3btwBoIM7oe68tn7xvQH3DwwcidOnz3
ctSQAar97TfBJ60UUmCfu/6YZaRK8z0rkTFiBwBYoUEVBhZF8GNY5D1vqiedvQBIrlmmDI/z2eTE
PpLj29jXwvAjIBndPisCQMdRlODwqKBGa9gx6qxdEXq8iPMws+j9/sm7/u3q+efA6iBxlYV8MUZj
fKa82UGrpm9q+quCJXwa6mzxXUinnKWO+gER3QkPiwbPtkirdCUVWlOnh1F8oUuyWYlY/gMO4AYX
9GyDWXekF/OHj5HEFdnMXLfE6spM7kc2X2X5tUuOAI3xZZoRxey062yNvkCr4uE2IMoj8dJqR3MX
9TzsqXk35AptSTW269FBzoqyB9WwcGfek1E4C9O89DG1LeZXq1C4vraxz5HB/dn4/flDA4opioZV
GBC6Y+VzICEhoWiZBdSQ13Bnio+HItjiXkPhtl3/ODT+NQYLdCBsMCHqQErJghE6NbwXuQvrkc+v
23PrFPA/UmDydI4jppNr21UC9Ejz6J6uT0lDTUcimeTk+dzzb6If9IV/oLra2Typ2EaVEnce+ms/
LyXpulgd1nYvo2WbJ1DglM4dXb3gFZEoKr8Nk5pcVu9ENwRJmYWbSpE+y1MzsAsgBMJCrl3kbbXz
tmJe16k6xS6D0ucrqqTZuB+uSV4SRzs7FmPetufN7AD7j+lTa1qSIqbYcUknkVxjNU8HQ4pe2sLe
LN7suRRQYt9SM7kPkMSk/jIiipfJVwk8dXUIYAxQORG1jO5fopB/SCrNdSsx/xXmRziMFZRyrxWR
5KVnESJ2ZmpY9Wo2XLG8AoQ6XGwv9bxjCx93HEt9xYr+AgMatoblQzN9HFlZLukm5e2MuVz3/pCD
Bd2kynRmSh7VD5TWwKWoQM8ubEuU7UtxeoDIaOfDpHpBD/vx3mkzXNflb+8GZkIo2OUWNHbjQo7Y
sV2Zbk4y8H26tPxuGx9Dg+E7XClb+XKwoqYz1BVvuRS/8Mgku/vI+cPpGzVq2e0W2q3f0Zo+k6/7
R/YyqNGGINzL2VuDhfjymmK4OeAZ7vZYz+k/Jtwau/JuOUCWGz1X2Z2DwJwDZ9KDlls70JBhULt8
wnzd4Y5H3JE/ckm0BzC4E+gob1DG2AA2eKdAKxBUzBTtx1hGDLIrAjQ+l2wcT9qrf5x+LiyA2u4K
BmENvjMjB8SORtKP2hcqVkJ43HOX37C0lkNGjQ2Bntdh+8Cy+HFRv19m6qmXKjBxvVuR2J7b27jN
HJlGfdhcAKCX+LcpZft0UDMOZljE1dHmf3C1BhLHcSHZzcErx5tbw2puQZvPNxWwK4bof4aVGyKb
liDskK8GnL+lZ1rwyspU9frXWsmqO4g0hJkFdpxLy0Jkjnl+aeBESzMk6weqnf2De5vgLlcXZJhR
u3xmfqBkzBL4blbDRgCIKPsggwiUbQcWyyAh5zXusTmyVo0SQ89IOPZ7bTZH3wfMxrszJDW+szfE
sC1j5N6VsaQntg86GY5FReTMWO38L9aXjDrjfbGVZqY9gNFp8HO15zs8qhUvBWL4GCEpPr+IjupR
Gi5mO8c4+O2xLJkaMOW7Lxri6/wcZ1tmoaErS//bqJLCqxd0yrUKxuU5EGmvB3vR5m+unhZp6rEK
SnAMopxExqN7DIkN4cWTsGpzjK0yIAm+9MOwI8c7EEJXxKsCb3Dk2+jt7fVg/r+vFd324V1+EsKr
qdhmbmNy2zSg4IE40KFIYwVU13ff+5TWK4n6Xh2VjN7ciCr20WgUJsWOi/ijD2tPMq1Vw9aq+6jz
yJdOpxyAvaxT9e7oWdip+pA0i0v17uN1uAT111ZIFuCPySU+JCQXwsRiO90A/ZsyL+377pquae4I
0JOK+OKWpNFrmc8QEw0BkaWrCKFKHwSNGGgVJgr9wv3Phes9hn1Y5WuN8T1dVw0T0yti2CNfDddr
0848zX6zK3OimnBLOSBQvMRLP8AMBJWYay8HsHniAxOVqAj3HYgJ1yuPj+Kn+7LN5Q33YthwwnrZ
oPzrqYrpCWYrdHt/9GZ3Em/Hl1lr+BJxRz+38JhgjlYpIKPZkmpJyLZDDKmx7ayhdQdMBD0hTmY6
Yj1wmbC8DY16kVZ2AGD81LEMmw5aDpRbNLae5I5rAwkFZJMGR8lDAkby6Nk/e+AI4qkf7HtBQ099
RyoGkkihylS5Or755MNJUn1S2dZ8700hswKoPq7btsb3dLd7AcxxVh+/X0GyC2Kd/0rayB5YI8z2
hsFKGX7nQLSAfzoRFR2wGF3lXjn5Q+5eMRA944dAHYqCY2Vumc8e9AlFjAhUZcl/Tyqkxw/MyyxP
KKU905ZShgnsMiLRZYLLN1qrfo1qbAh0dowMgDA5LGnns5aF2XoNDmV6cDQrQadQxLrsp62iaI2d
hCaj37oV3nyE99SiKg/g50lz7PO1i1mgThwZ9+duuPOVZEQzeq/ACxd+EQTLx2Iy04EzyBSw6XYb
nBAYHOrebODTWipBphWGFXb0hqDEKfKvbmOvwWYGmS0WVHPVQA1XHPr8YpqPrJ+z35BxUWwwF6SI
pmx2hTcVL1tyQakMTsP8iT9kvgR0Xw3CLvvuQUmS0SMUzSm9HYBSbRoWuwc4wh7zSVQTTxiOOWIL
bnqY88aSQ688T22rVgkkg2nnes3zOu12wUgLV/+GqZT/lc2hEd73mp4/p8UYtl3wLTvKU48AtvkH
D3t2lAZCarCAOLEgE8owzUi3Wr1c805pZrx461N5ZDwRnMRpC6l/Yg83LLwc6VkhuxIu++Z60ovY
H+bAiNym0myO0RMhEtmofLFrH0PMa921mjPOmYesLUSLbV5KRR2lrRoCxpVVYC6lJ5goVISZxt4j
RVx9A3/DwipEXEM1Y9Lfb6ofEM62yept9TT8dkHlg8tf2K5H0xgF5Kg3wy7o3wfEYslV0vzZmBOu
ZtFxNBJU9DclRewqNvk3OcNnHtk9AlueAwwwGvEdbcs9aO1rW0sMntRXcwcDbdf47j86is3wmmhq
iG59M661YZ/wPMJfvPoa7wucRADrFBBR5t37NX73P7clcgJi9uUlcKW2W17PLAysz1M3WLgaPwtP
M6A85EwuUtlciznyD3z8ntmvk6o5qBBxaGe0MsEd2SfSSFamOG8zs4FwmLHJ6sJgUKKfvyUTooL/
LVzhrKJ4f2LoaaJEOTs4t3hxHacMwFz4nlY3U71qu4ub1dYgvucxd51nGXWbf1Dq8Sk6WXa/EuiQ
iS/Tg9nG5VVduWIFDwuUMipfwU/G4NnKyeodb+X5i8C4Owkg8io1WG4Oc3voY0vSyfcT/bjxJ5m/
Oo8+IGZQgYh2MJgJkiDfhbvowKP/e2muKHkE/vtj6aX92fyV6KA7aFx6AN4R8c0ww54z37xLZwRI
wsYAfpsGpKwbtWHNXjKByhCPNUvAgwIsGxg4aENwMqFGkkD7mUlRD5KQAZeiB7/SQ2Q7LVXImArN
HRc9oa42zWQXJ4x35ZH0nfRK5jW5B0qVyttzQ/v47X1wIRnh4/TqGSSdikkMIdwhUkf1buwOXAYW
J02vnlvSFXQFZram4wfzNR/u/8LY7Z9bWlGjwIUx/L7jgx0IOHLX2t5Dz9CTZCd31WQJwsEXEpHy
ISgKZ2Mo/Kd1QlwKxZ1Bd+STYSFdTU2MRWTtLDMg5Sw4RZ8ZOKRpO/XBo/xQVyoihLXSugyPaatq
tSfbBta91TGfnbNpfChiG8uIyiIyrqbNVZueqfyPggdxyUeCuJEopk6sHXUZjN9iQmBXBlGW8g5D
PLxkL7q5KijRLedEiLIwr/tpPycjtfK6uUxjJaG8/808B0N9JR7+QXbTmjCAuRRGk072StcRpVRB
76zmhkpY1hDKcMVdYA8Gz1Enfd4xXx5HNnOJuk9bmyO8pUYFNeZPSTEt+yRCLBfT887uxyWyyA2z
24S7Oq2KyIBaGYaAo+eCeN+loC8mpv8FGROmbky0P59Uq8XT5KWwbIrMnzViIHJrMN3gTe8qZVhq
tzDN5scuyI0Go2e9k48sCBNl80uQZbnsPZ0y1pGOjHcn+c8H1HEnGjo6B4WkTJ7HFq6ptIFx6IYz
qAwqtP4xopHXFMajtNqcGDwdrMDfpN6Txd3q8c4ffaGs5Ulpc4P594gjFGoT0RLZMFS55NbPj2a+
NJ/+Qx0uuac8nOR4lEem42esusQ2QngHDhQsuCNvXongms7KDXd8etux25XlCBzxFHC23M/PuDgX
m4YlA2MmHE8+QWswJ+5IZ5xZZTQkMWbY/Wj38z7ayjN55hEiIeoAGo151sXC9LlVgvBI0gkkFavm
Iz3Qp4/FIYpkCePTtqtAFyQRNrwrtn0HfXoGEaVXbvS295+ReHg1WlahgcfCGSOSR/2q0mG3bGUz
xnlW2ecKb7G2ZTiUoc4ia4x4rxSA4PWyzzCPcavPE9bRx1TQMxTC57/ZFPn4n9pGT5GBMaA5y/PX
75MGYZQ4aTWXojRc5G5ufDM6C1RdKz/8hPhS81VG/IZhwEi7aOAU26JSBJ9p5u7dYasigDCrxTcf
rKXDBWjb0ee41wueyw1F620Ko/Y6AalD6sJbYjbmxRvJ/djzQXU1zkT03/dEiCJe1pn66y3TATzE
z0lG48LpVVLQFKBrm5ZY8bnmIGhlGl0YwuHq8MgQbDWIVzyaZCR3pcFwX3ZsViammabeeCJ2b2Ul
2iImFjmejPznElS11cg8nlqOFzcJHK57grgKfJYjoHNuHA771/ZOfAzxakaGGxcJC4XdfWh0IubG
shp8UalH5Leros1omyF0EZ7gkIsdn4QudOyouAI0w8ojgGaSatxnsjiIScgejevO/3UUiw9o45MV
X7vDNPIDASsl4dsRTnOifz5zPRnxraRbjsGuhK9eE9cXNjpUyNc8qwIKer2jzKl9hgoRaYjGW9DK
ByEvkyj478lAGs3svjoiOY3H8FjS8tRRV+ZfohTmoeAt+GvzxEVuye+yNk+AwvXs2rpGYRGC2bB3
hdRsS2DFj23rwuPZbZE9RTo677MFG/+d0rUAK48gdE0fAyjYfoyfS2iSVdYnjyzT5cvBYHWfYq3f
glWTku2VLMk4ze9Ys3Cj7mvmJrQqXYu8YzC+11EZO+UKlXIzMT75Q3UgTamCQcZigQlmOXfdrK14
S8EbhyGXoXlQ/+oUib7sI15rzr4vsbokx6dyoVYEWYiNJJ9Nv6b/rZwUq5tnSUj1btNmnRQMt6Au
lQc4Uh6Ga/ktV2JG+YLLbolxq7I6pc6D/Idyddti04au39oW21Y7D41sZvqVoqffQ9DHZgvXylM9
0hXcflCoUGvrKLnSWKKl3QYtcv9BDGiEOnDm2yU4iJft4BVgBhdskeX8MEXnScc6ITfXTEg+0Dlt
coIHtcoOyqi+LDBZC6imjj0cnf5O2CgDamQU39APOI8xDFtLGFk+iUv+X3e/BfrGd9Wtdq1gnopk
+0rR7QFcbknuBAuFNR6Z2jphkg3rBcsens+MOdkWV98801RleJW+bgj7MHofUnJ/P/7hHpuWhdjW
V2oR1zoqEkjm2WG+Q57aU4AK9/oIs1koTmHq2SOeNi6EA6EBmXhyt7mOrbbmV+u4fNEmeZUfr7ap
JObNW0mvNiFfSPlDw8xefmaJ320ajUFGW8ohzdwlODxavi0aqsV7aoz1Sa/3rNAeTlbvHsFp2h+u
TTcg/Fc0s6YrRHQuR/7xIwZlVyODWS/CuL4c2oInaP0zeZevxxuF2AghTLMChktAmneVJ+vzHbpq
INPCbg/Jtu/xRPd4JQgqUSl2zbK22J4cQ0s1cecateB0oKKJdxHtaykyPX8ug9idwKdaB1siNGVh
oFZ3pq0IKMSOjRLjdPgxeKnzWrHZJ6fFeQGwlMFKJJWNVGDZCuaOc47hdwcPBwem4LRY+5W1INGm
344tyu35DBpKEzhsGzQzXGDOHl5zFhmK+6UAKrWAimOd4cgTA6PqJLxJM0RfDyyPboUO2IfKFGjf
tdA/06oW/dUlQ3ZRqb3lfxP1J1vIeKrYahEaal/a6W41yRO+M9AYAXvSECPrx7RLJc7BOfDVkPsI
do+sPrdBmAgKNxiePX8gcVHenjaJV/VSUjRo4uDCUfuTRtMhWRAhkyLK0knOMi4w84/N+z+HV0G1
IYqlKuYi/yUSI8eu6KLyZKj6Cer8c0QpGDLjOAjoGHitg7SM9lOCdt+7SJvYjgyh36znW2oVFocj
b0sNYHuD49n8V43V5/PfnEP9noGSodG+2lH7X+iIgp+MasEEs644l4slrOBg9KiN/Aw5OUh4hUbk
3NJL1sJYUO5OV5wIcBH/vEVNrb5K+MxQypTP7w+AvbLTcwLI7E7nBQPSuGUqymPygB1Go/bOgG7T
nYTFeguPS/uaV29XJ+zEke+QnXjF7yjm+mw/izAChL9csXUaicRYGKEn76DA0pYkMVPNttloMBBR
iOoQSltbhAhqCZFeAT4dTjnKRqes2WQj+yDLfS36pn1YVtiGZ4MN1JTewUgJnNOZtGE/VvyhuhoQ
sJLxL+99DPpcBvVgb89bBuaPIW8XNKtXuhFvk7qaCrphyh435yNQ6g87JvOEROdY9D9qZ4xtriNl
og8ktPYrkOPoap/265wyXDKbJonGWI/H2EJYiYlZLoxbFa/3gIs5Le8R+0yIAdKj3Zq/uafyML8u
lpTNeg7Xa3LOF64IWHfXmKD5f0pO9i/AzfgoMyqiIp8Sn2z6HDBqkiAD7EOcrNnM9KZgbeOU21Az
ed44dd1HWznNHr4knoQgOBipfa9DFHgT5MYT5+6SGhSmki55pqhq8samfsm1FP33nZo1wiT/saG7
H8YU97wJ5PeMuBVS8yxvEorxuqr/0wZX8GoysQkgF5HFMOy5F5lpw6Z7DuUeFfaTD+pGl60zY5kZ
bke0+gggXKzinjOe59cFT6nTwiQsQFpcCWnLXfwMM3aUW3tKv0GPEUAx7DrPj+lxVZkJIYe/zmo4
y5XNxSSc8eOcEug9MsT05c3umFuLEqrCetUjmb6zOKchnNl4MyANb67PfMjuDdXOt07mW/wdQ8ai
+11ls8QJN+l9TmFw5m8PmtcwnbjW0HAjMUyHUBHWCPFoHf/9LCjTrQZz49bI18qHrz98b/4xUYsG
r3aRifTDMjzXnU5K7cxK0nfO//1GO1PrCtt3UEYUrbKbJHAjbsXkHadQ+fZ+tExigYZa6q4X1pDj
8EWy7LbUoHb7syNCfBWzqd+HqCAoFhtKQvlA06MufqweUg3rCeQnIEbR+SoDh3bWIt7XaIUVzrAL
5hlwMBgPJI7dMNwZ0c78K4oO3hNPkguntyqdKJfbY/i1GwG80HdbAKw8Y0Zxyqndawq/TIp1JUrY
3/IBKfvKwnzVLGIqBq8btdAf47Folb4/7RQV56bwAyFdx0dczsVYFDEZRTtrcNSKkTegRPMSKi8B
mZiJIeJtYLxrUiFrDnX+hT3d4EI7257hxliNY0U8241I8fOG6n4fl1XpK5RXEwMqhMRhRsmbmfEx
9nwv5gtVsTQgdI2Tzdbp+BYORrEXt3WWO0U1hNer2ugYSdPIUzzCepUPRcvxXfVWYKaXp7ttuMmX
avtxYpl2apGUymKQx00xHSnEcCH4jXLTExPcPi7FT2Kqf1sPIrK7fQtuC9VVN56QHgghWK7VO/75
wz4MA0SWREC4FhJgSpG96RMR1rBrh1cqAqDEAxBXCdSk54fWaOZaSnJFXd+sK0l3rMBAbz0M5LOf
kkHhVoX4bPJkMTYzx2GbVTU+o5uWi2fzB4yYFeXcTgytQP06KgbSpdOg73wLQWzrzzjnfpegK2jJ
M5HeoKHtUj0dUhLqgqEGgYUrrJyiggCsjm8v4eL+7D2mJ6hb1zQ7U2qz5fx4oyS/ow2O3mmNtMvX
NHm/AHPhXZHVdDLlfajdW630WNhKN2MTODMSIIiH4a28Tz54MzSnWpXXMGb8tHwOf5ggV4uoxKah
Eudu5mYkPPD/V8pmSZ0TR0rnkOV7njUOjJ2pZzP9enjhdxeK9TBEBqfYSkPhC49oK9522s94JOfh
7MRWD/478gyBBMcDLNScxRtG7K2795QUVQy39gch+lX1XRCX8Xn7Z6+0m7+XqQb+NjljTXH6GJwg
HZa8/rwBzj7zsVm5tim0/G2283osB6zjKaUfX+ELVA13c2zS5roT1ACh1n4woRaddlCLFjeR6blv
ylfrVIDDY/krq4K0XHOMGW3qfye89J5XF+Hk6wSCOlVex20nCKSCBAZSo/wIWTMciLEnJTM57pvV
cYXYDuYxibZPWGuf6l2c7oth8LXy+yYWqx15w+Vfjl7mkS5G4DoLQsaFOssDkZhzYGR4/3VCCkkF
mSwnCaEcmanClwvgRLnQBX0mBN9ogukD2LsnjHnpRW8kIfZQfqaWrC0NdGBA1Cnv9rGMovWAqFDe
6oQyAv35YCk5CmSeqFHBhq+6/4mU9G07sb1rJzxFi2dlLUzuDvTMv9K9qnjBOIG1n5YlcWpHWPFP
VmhZzfw7dnDTWJfyesQaWtuHtsbivioT37EIvbtS6O0Ok8fvSv0yVjs37gHVZZ8bYxariGL53G0K
0kkBilJzo/QBIKiBKl7aRhyHS37jgdxslr9lA8PxaF2RO1g9Rx/LKC0ZW+2+e6jV7Fy6Vu1yuGLR
DECCofOe7p5RGXWDAf0Cxm4tI3z3zScOgecH8wxfJTMN350oFKKzox9XRwxBQjV9z9jqX6LY8VAR
EPMPx60dNWh8Vb91kjtRjRZ+ZuQlENyrUxDbc2yOi+jL2dSAf0BSDAsvEyKBJX1QULQHRYS6NqlS
owgwneNjfy7g/Wgea1KHY7k4m3Fd3d+b+7TEd4Z7qxsz93OQRIrUYF30UOj93mg82268kc1BD9xZ
fHtbgzuTLSdP9bJ3M6RQi5A5t2aJWJ2usP6pPznz+oJQHgK6SSnTicBY5I2lc8xGLkAaLUk9L0GW
Rs8rlUHWJBj+gfIuvd2kUiJHBFKJDS9nW0AKBpUv4j3ddm1WHOSlFWLOPwCuwryU5utCUeUuT+US
a0uP14CldodvPKA3ZCbOuoN3TerVvJSiqjXLjGxQJq/K+RxXOOzOVS032uZcXZzFxMfxHcF2bUo9
hmnrzRTDLwCCv3dq+P27TzWgtWMCqKl0CCuBA4HI/Tsf6i8xQsJDLIg/0HQFZdMb0oAxXpoP2QXj
//lgYSm2FeGocKRiFUgAPHLmfOUjqiiEdAqgR95sHDLGWYnQEGW4h49PvV9QM3MQvjp9htu/vjCU
Wauj/qNVfw1P4/zZda0OAR6Q2Jo+miJtTvXHGEZJSKQ7C7xcEC3hOL+/Loh2hfxn5m6QPRul+cVa
r4vWrFktOcWNTW63hARv5Ts37DY5CtOE9jqjosktkzweW1WzIMlDh6gRHytWemwj7RA6+BrHgP/X
1VJ4T6SqWFhR4SmIGNnkMtITmq9aHY/lStPkLSvK6hTWWGYp625Fjh5fcoHMH1pmcwU3rhiEuwxk
3y5GGH+E0C29tzyQvQDF6qw0VPzRrOHIEctBR2NVkaM4Fb1JT17J/ir8XhmxlWNJp1hqImHep+fx
3QgFn0WWR0LBN3Jg3tkzgNOCE+ge2rmdB126EFx5HuwgE4xj4wDYZXi+TT76rDDJZUGzlA8zTFsb
SlZ/RlzbrFkBGhjOpleFXQhDBp/+e4ZbAEwZ5OM0AZUJQofdnupKb3p+Wx9aPlRExW18EvXZ45/m
ohfgJKIxaSrGK9bdYW/KzOiq5isGD6tqpsB7MzuJDkUxIox8tIifPTzZWR2QXXS3QdnBn4OIMAzA
Dl9ja4m84ymU+dnCiGWh/sd+FPajkTlweRbo/HaYsr91OMCxamVVfJM9I32TfCME/f5UNDEHpBOC
bi0hOJ/y7cAg+GcSAIF9J02WUchjNhTvSDpFsMKqSEPhxCa+MWCIxbbhCJEhdFkXaPk/q1a5mtP8
dlvF4GKaExQuHdupsr5gosa7P9O/bAC0KS6dR7JPkSQFu0OaRC8TBRQhY40BG1C2PKyU8qm0cx06
cB4q89/V5KcnVO5VaoTq2dntysvCmQeRlOOE9mc/9xq+zgGZPoBgjUXOljF4caeuhUGUpQzapwbY
Poz90PeUOimHj0DBzbQ7FigK90EFLE9gNjFbvZ+oTx/IW5a3fgA9dVodWZ/SV982mDOwzYFdHWhY
AX/0ssEIGRxFehPy8FUhQFMwdFq+aPILGgxDtsRdh2HKE64Gkpz39/8vCtTv07nokofuVhRI99fC
crEJHJRKO1ht1R2mlQM/sEbfKfBS5nkxhFuVx0MDwIBGUZZ0xEZcEFrK7HFiBGw6xUWpT7d2eIRo
pu7rvXgQc/I3wu74vWw90wyOjVm1mwaB9QaMNkkKbpS1230YwkKF2hSfFEkgkt1+RTvcmJsOTGwc
h4G7T8F+2RGM3SXAAOyjK0PpucQzMzN+c75g4oFDcnTaWFZ2nIau95NjJzH4lSvbyg/D9yuohlS8
YMQa8IwDxU+E8fJ4SpZnfgEQjV92pXvpKgTNN3Vk88Z3A3wutUnHT1oOg6xqO3wmtnP3+QYAV57k
EIc0xMk74c6J8g7l6E2btG7s/L3e9J+FES5DNFPmjw2PAzy73aqIsWSUaxQ15+/KHF35OyZNUfnu
DxIJL6o/p4AxjDYbqvVeCa/oyLJg0EPzkyUhI5TvD90FIPfBRVQxMDfDyfKCOf1o59ehQ0G2wnyZ
cefEztvbw73qhp/bAdjc7kKb/o6aPaJn0sorktdvbh3nkMVBRlWq7jIx/y3YgooYiUyY7lPV3r9O
RUxPSdRC4XXOXxjCiSZlO8D8nc0y45gE44mGD08yr+DfpGrL7Srsj1orhaYiEjgOB2q29yxaSFgq
w3wj41Towtqq5wgRBcylQYphHcVOC33deCLjN22DgvcJjkwu8c5DnpfmvvDo/Jw2vy1hUA4XEo/V
8LPNdWD7yn3N0Pnw+KS7KMyuTG29lEvPOklIjPqvyTDpBoSuQXzO70xDY0NtmEGhvHT6/3RRGDY5
gdNp2W3UFVQFKgAHUO6mkEU6IGlW4fR7rIqSLk/t4M33hzeaCDbM2AacRwBDvHyt+dXvEIIcmuq+
lbZHXFG85pJFTHL6xRzCEmlBjn3Md5o+5O2juY5W7N62uiHkIlFvA4aqK6631OXjc+6NtNq1T/Lz
iMZcK2+l8r684hf9YJXLiDXauea88d3z7yuX7SD3L/eWCt/WOczaC7V9XMKzvGTrThSXr+yH19nF
RGbyjOvkfdkEfdCUBgHQevh2t8s9eclwwsq1yQ4hQptRFbz57Ovtn9UIUeXRpJR++HYSIAY+WTgf
m3vaDDj80OYHl3o/OtSygLVq54xf2iLD0Uq1zoqd+WI0Fxq0v9I8Oy/3Eb2CiARHWmUJ83ZuG28/
MsCOJ0ahM4S4z9zFziOc8OQzjfeiR1V/VUH3P5quAQdfuEMnzces+6sKIEL6SEADY97kXLrBBfGo
571QOAQx39z6dhzZFg+xFxAqGczpxPUuMldQq0+PfFAhMHBxT8ThBOtjQHGdGZ1lw8F5rdJOH+dk
LAL5BJ3oXJKt5CbtEUgqW0NEr+sHTZAkUROcRAVqx+CqAgLPlOCHPbEJdUOezXtWU0BWCCz7dqaN
4cjjFvh40QHtVqzz2ltAuMbb7Mn21UoooG1fmCjX79pN3qBYwXbnFr/vzPMn3tA0UIrRmmrDNAxk
OnNyFWFZN+gNhm6NTq4T1a1lxu7E3qB+7w5690+D2bt6+Fj0FN7AQjRCv0oJIRO5a7UNVUlqsuuB
hQMsIQC1HnMTDJsrG9vRSFIyN7hB5ic8/icoYApvWuT8duwfRRMi1F5md3H8enq49zVf6YwtLuB0
oitCLuyu8AXy8W4r6534lWxx4mqV63aNjlepE+hSsUkmhpgad/HUrZE/0Yiycr7fXwE5ErkeSn7b
sAwMpzjeLEaQECxi5kENxWpp1lu48o8IdBlaHoLb64VhmzVr39gRCwXMh2mju8ssdbzn5WN2a3Lp
oe7Tj69nw5MLasxX5Due9UW9guifYbNBptH875mMUBgCFKFgiwZDGRxu1J6BQwy3Poa95aAYhWhf
3FY5jdm5miZn1ERDlvnu0B/7x0UJFmy5pf02GpaNZXQdwF3OHsOVXIXOc50O69Yw4od8qtq2rrAG
NGm2JrpoqoJN8LGYPL5wJLAwHYxnOFetf4bXRquMQW71/EAr94LadUR/LqxtvBWhua9K1DyUdxG7
xTUsJi0PB241c8s4aOBcaCDsa7SWuqUQPDNqr2IHTWZ/uUZyQL3dz+PW7pX2uFjttJaIgYPL1nFI
WVcaEHujdz3FekraFjZZrzzGv0SSRQacvyQao65Pv242sQKjE5yacPxNeYq0Oh0RsGJWC98lbSxD
PymYLSib+CkliL/rJdQ0Rh42VDVioIaFggp+WOzyRDQ9gYN/nDvR1WMCW5g+i5rsgoRGFzuSgn5l
1ceomQnbzfOAuljSw1eNO9oT52MOXPE8RfITYzHJrpFsT3B+AcOr5A5s1DAGLzYea+JhhzHNANuC
4vic1w0YPGKjLVWKBQbSleGOvnv5Hp+v/QCB0mf/j1GmyuWxfMz6joSBYcVT+j474AA2nI1W0gF6
dC5ARUHN8ePJm1Ihkmrueufa/4mqB3oxdW3PR7zA3c7kw6ZoY3b6g8AVt5/jnYXdKYhgUUcpkgHv
qdQzDpNrh6CX/aOJbGqNvb0RTgi+qyB1zoXunnRB1zLoX0LYv8rhViC6wUr3Wn7Ej79qegjlaH6E
YFOL/xxxTKSFGAPt3hPXWpoY033LEK53iXB7tc7GGy+JZ/D+/pmFutFvmGTwpZ2xjrpGgzi7d2ak
zur4ZSFqKBIPvW/UwYEb7AsaoYD7R4Q8+Siv8uW+F4i21qKnHMs72nkJ1cMkeZ8LRAwuNmqs0RbD
gd1gSapRHu2ot8sjL7lXP2UOY6Juzm0gayeM6bmuQ09GMYVxyvKTsfGhFKAVx+StxFj1x//zGste
GdPhOUWQPWVaMwrkoOMnF7DcuRSDBtcVeQ6haDzdhtLO9uCnTY8ObfmTmoludk4N8UMbEd7IGe5j
eCN7U5RS1kiSeWQ/UwhmTGxfrG64E4yDkFwWhB57y7Ji3TQBmAd2WoU18ULNrwWwca44f2AfIfj6
3rrCnM+7rGJiSMLgdxIqsQRbxyKE/dKI1Lyue7VXuFsrQiMV7ooT0jqsKXJLy4rKnRVPoThPpgxg
xjvdDdxxYTdv8WEAytIEWT1D+wwC1W80KLhJrl7gYVLCSheEM+HglPS9MwL+1C561+pYAnmlH5ab
rRsKvOriz9qOhUtb14OHd5GgLtceri10y4XpAdem3u7loc29Uj7Ua3D0P04NP1kufCgzdg1v5b1e
uXtL1+zrjZquNs8R6ogmghEFJE3hWCbqNwjiyyR9hX2TiehBgsttcOjDfZ7it2wBaF/DAC0Z0gZ8
Osa1ogDFSCc8zz06M0j0RY28k0IovTLdExlWUF0/D+eQXFeYwDjOXBs+KFr+ccicMhJpmnUqaCYQ
nwv/b6lMjyan3dNBwDsvMug81fY55nR2oB4h1LZTlzV+8AB4ERQED+Cqhj3lqcgGqya7UFofolWc
3d9PsYaA09gKG9E7pB8aarpwstqTE0wwYUeoUoDlT0AQf4hgQTOA7RgNMtoa7ZmpDlvr9VRxOgE9
TeaF1rgrCQdpVfpIrb3MXDuI5onpEu6J3VNSu/CtzS8dul0BzoEYWzCnE2nqiTFdqKDez8rDQASr
VRW3DMga8DT/wN8NjABC+scyFUUARTLlHQyngMshWJv2+Zy3tw/6NBU2TdH92cEGEtKHix7F3luI
x9GS1B9zK1opdOh3MgxTzX37YjmYPXckrQMKYOoA3jWFPUi+QNAiooj9InuVp2csB08MbBxrGRR0
E2m62yaHAfi2clk5NMq0S/H0Fd2Cq7RzmMgW6AjxziIoS5NRm45NXyMeE2XLglILG1Bwo1oi5BFU
/p3VNCknk7qa+J9Z1mXhiOGfzSF+jqi2MQMRhiPwoOH5KeuaFiRsL4nb0ZKTQnHgS99Infy2vb5C
3ctxDeR3KhgOemM3/H7iIGVAfCHaTL/JlrSKId48/FSOW5CkpusqSMbJs7hMHS7wJnu83dq232xQ
x/Uv4rEDwkCIXEImjddH3fkDX9MlUyUsizfcKu0SiBtFMpYncgjOIFd6Hr3GODyFEPBJKntVSOQd
juAKB8DnTkmJJbmXwX1OnbqSAg8kx5Gt2qd8dstkMDzRqW+c3t71tnOM23xPsPihnAAspXt1ylB7
hCHq4PzOvEUnHYNQc9GkAjU/QbjyirnklyAEojfISJaN2xxFQpg+aVX94pSw4S878dK1Dhh7J3f+
ucckWTn8Gah3+e9Z2/waqYQrwU80+7KMAHxb6o2gLxOU6UELq018trmk9WehSl3p/9aBPQoI9jVK
KbWnUU0/HloaRi5aq4wrCWAmijqm7iQma6xGujSFc6RsEXHUlTlGmlxNtwLcWAW8SZwCpG7hEKNB
Odf9q3WDOXeB1qzfoFiYXfHZ3hcCIbiACPrGYt3W4ry6WvmB3UNS4ZeGtKp9zjG0KggWgqe9YRzG
b4GL8mubeDFZDw0hAZr/zVG4vvClgbpfdujnY1fMSLSTcOwAdbczIgkhQxU6XF5Bq0BUGlHM7Hn9
fltp1KthGN4oa4w21urnr/d0uwmdy3en3+mfyemVzje9W9IPd6+bfUTngHUgVYTuCDYnT8ModQkz
PMkbShVvj+5K+xfx8JHJdNeV+fGK0dh0IXO15oL0cCJESqsHSVPK0apVSnVhNw9NZHxTipcHVClJ
CmEgJYp1RbAyAU0ZDCDXK24+LP1krsTiRlNun7RJP1LTMcV6CHEp5Z5w8KeDopv4oNWIhQjBW2Hn
/cmlFzrRLNz6RKvZNcEhgttP+FaqQ6KLdsbsyDO3FQRhVoIKzP2OL4+r+HCNRU+oV96e2huT0uNA
s0pFn/sAvxQ8Gg1lbHVNIgyPlx2ygu/xPeYfqzy+Yg2MPwVIXOFV4i/r5iUA6fTRaXar85W+Gzq0
+mQjrQMZ9+j/sZa0ZoLcqz6ahpZozi6Bct8lgYPE7WfbRN2mNTQ8a07lCjglz1VY2I9pTrY2dW7T
iAzDwUXYj22eVDTz4nI2Gel8H5pPWn5gWY38kcAaYeF8V9TmzMlcwat33WrXpVkXTVzGUBIO7SkG
E4QnuAjvOyhfi2JDPCzZ4ATvQ3TUweiE8o+yQUVtRDNR8hUpQxWfLVF6vG2JtbUpYkOruOcUGwzp
CjQJsQEI5cPHdV0wzuhLUFKSnxyitJiJrByz19bbwSDa4P2mQChEXv/vhaRNzni0EPV1ZrXolzBN
nJ6SUJMf3P0nLvpzjUz6MO9osLOA77O+HMMjW7l4sjsSnGRcaHbmHrAmKileSXCo0hsLuzMi85Cc
XFDLqoxLbS8Yny/jgwe2wrwbJ9AcQYziDavqnKnSmSTSUaGtts85OjZJ4UbN1VRU7isGlZMrwa5T
NycSydLkSlf1BgFtX5juDA1J4gk2Rpg+GFkCukOQCRwUxLMwtr5wsVfht/Zs3cnG/zCU+ajhnXnV
AAAn5OVNnxbXNSP/NiPjpV/EZqRVoz8ndNfHrvh6JGIN61H0aI8SwgnBuiUuzHa1EGQeRUsVuBPK
3jR9D8fUFh2kIH9nj7CKWYcoBo3TR/InCbTW/1VKWR1cqO4zFRZ/1uJ8qn0pDXODgaRmR3jCWcFb
XzrBOdAu8fXzbc0eUjhU+4mQYYFaGH0QJZ+8uTWPXUvQYPEsd/w88KzGSavSWpRzE4oq3jPpj//4
DAJ36AxJGsw/CaxL0J4gmt6D7aRqVfo3pPPpvBzHVNHlCrz4h7wlYz7mOZ0YBb8wQwXKS4+uEDPN
gNmFvJwtJsk+avTBTTPd7zgzNUmSDwwwj16WV7Bi7eG7CMcdMg/gM2JTuxubuNzidXvk9l03yHFP
6Zpp3PBpIvUTYjUTgm+PVuzXsi1m354ScTt/TjiLUYx2U2/8yn/JX8Ihu/JSszq89o2mn+msVb+N
61p0zvGua5R/KwC5+b+DEdnvfQmYueembCt0ctsSLDR32FUKUltNje/oQ/0XVTtWsJHF6e3bon0b
gbQ2B8/820NENkVK+alKkLC2/V/TWFxmGvuQW6vtTjCK1dgY43bKlaO+f+MeNOBeNwB7ElCCP2Y9
cHsF8FLCXmGUoLFBwlr3U1++/U2E+jRLPmsNqwadTWdVpukvgUDh5WAtOTjVcoAPD4RWUl+37dI8
oog82j4mym8/N3GO6vDiugkLl4DVv2XNXM/Mn6Fh6enoNDloOb3Zfg/AazS7kTT0b8mBInWRCiiU
E1LWn4HqCRzkVWAM+z6GlLR6Gl0Zds+2odm/bmGN6z6A/e/Fqs1t4phpkIz0PgF4tSWii/xcidMP
GFg2SVKys7joOxBlHlqTOBs4vcoWn20yTS/8dt2M90oXF8XbdBrTHT75NQpapDSOcSPEJmLnq7r9
NycaR1FCbBvpAW8VAUpjdTiKa8Jp1CIzFYU2px7ayRiW96OQ6MAlhvdC2cmMpD4XUHJmotYiV0AR
faJD4qbJ748YNn2wYoODVGgN0p8ofIZmOAK9le1S/2ta8n0yfJzK9cheMhUoRqCXZrRLW+4rZWyg
Ol16HUW3Wm4SA2dUTZwhozPDfq7xT8Jxo9/60dWDZlDJZIFe8qnyQxPICqR8qA0aTp49HlLZ+8vj
2HWaKvIf1rlyvT7oxnKFyG/kEaXLPTe6kVE5UTiRUYkqmaCA6GF/kHHamI8gMlQuyBaloXvyg+gX
gooc1cvLPpcQkjZxS9xN2qmQqQ3isX4kFTGc9nzEfS09QwVl9ARRUzsbP1wxy1zEl7vX8fulT5pE
usOZp1C8HHjl5Br+fheuz5MHssvBvBot4zE3Gy8VKqa6MwqPMD+iDJscz0+OLPRFfj2+3IbZ3MZj
K6C4NvBuLUaaWFT6Gg0vrxEVRbeYnhrBhlU4Y5GfguBbINHHBMRBvLyYSAfe2iZcLgJl5Tq6G6UR
QBg0obVghRNr2iLW1mjYgSeITjWz/6uBnj83jwvPDHqWExssZhtCLaJBmUtTZOdXXhaLlT6dOPRj
5Pe5VDDkcUCA0rqc3rI0B8cWUCTkcZTMkmDOAgkahdMoTLVpfaHAzTFQxgV0XOWa6jYkidO73sYI
//JVJkhIs4Ylv0KvieyGzhcxFC82uGoGz1WRTWrq/hYiMEttVvLIEl08LcpHe4Nzvr0JhXWq6I8W
HCOAKVJjwAYx5LwXZqpqezO3hoEudjBay7TXxt7+Cx7munZBD5zFy4iDF7smbO7DPCTPbu6uGbtO
Zr2YknpMKnCYuqIS6kffVsdBfKfGCBeH+YgeJWDAJMkcC/cATFMVe++JTKOVundED3lkcHjs6t5n
nalwThUchDpghhzioNsW8xWOtkahCy6g7fl6DMAz+5os+k2w4JhWdwFoG2YY11Fy5HO7TPmFrEGu
5DUZmMzueN8K6RcmOFht3RK9CEfEyNZHcJCB0DHSv8BUZKPopwECBYCSdJ/1K2+ApxCAxv5bhvzR
WmOeR9BPLHVicuNAxkydDWEQ9fDhSdEdC5N3jxfgH6yq5aV1LxS4T9xcC+yqsMtB9vrek/Zja9s3
oc8RDDUZHoV5YefNfUVmnzV8gUvcfCI6YJ/gerSnBHgHnRPFrMloDJoJGL46ErgK30hBC5vbA97H
DhObJ0ZtlrP3OKtnBZlkK8b/3cjYhw0UXflaF7jF7TDmkUnqk6wKAepZGdtYEwvFvEQIjN5ES3xm
dmlHiQCxgHbUTqZmklMEfUMBEgexB3Q9/j64jkmN5bGkyn15DSmEZCc0+vd5dooPrnhEWduEalZt
G4EWHJ10V9Dif/5lSVQ/RtUYy5UemYS8eiUXzbh4dbWMvCAQuuSejT95B/wgN6LTGvF0XNTk0wgX
zBJbm11mtsC8a632qSVZccpxYjL3kDDErSfwj6/AO6IjfUTxdTI5t4G9zN52Tm+kvELA2f3PH2r8
QXMaSA8czlw04l7D8j8znz98c/u1F1C3/3vCsHciUMUeyQxhz/SYZ7QiNl0IecDwbJHRsgORLDBd
md11LbAai6r89f8q50lQenUM+ZJOOQ+47SrqAQXQDSASFtuLpiIBMJoRJfT3pygIoFaYsqSQNa+T
nM9gnN1/VH93HeMcIIMxXHAwWVUGZRDIJqMYm90rDoiasIRHjUzFWrq3auLQGkOTxPvkECNvk2Ty
zhS7zxmqZV32HjTYYWXH2XFRQKI4SqTQbR7QOke19hFwJXZxtxPdNqmP/dWG9r+O4zOiwlHkOfrJ
WjYWjPpi7J5Ej1lbxlU2RM8fnoHHyelt0ZBPg/1wMu2CRD5bkSHsITcEsCPV/Hitrg8lZ84cbJCI
gVbAWwSRoFqYLZjxapRCAu9BVQ0C1vPpH0WHJDossno9sTAe3xxQ77N4oAPN+UYjSZTJaRYrhLDU
k43+4HMiNGwXC8Cay8w4lVXDEaQ6YhwX9OO3hLzKlDU3Uw94LYd+X6A20I1z6puJrfJougmmZJEI
j69Uz4E7SkH1wy0Y5QCE5cfr6eTOp6V3N85Qgc9BhwlTvg0iorvRDSGUmxkYZAml2tca3xZAbHKT
VQ8BLv5N+tXjDDeqVIQhV7wJZNk5wXRWyugFNaw63QQCR2RKbpMzYmRQHuH2LpMLdqi9VAKWXX7A
F0MYZUx7CiflJfM3WfUErfnK5qVM6iSyVNS1SEWaIgC+XK/PgDZpniE8QjLEz0wgfxSdJXzfl2Rz
gIdk6aZW2Dd+GGQKHtV2qTjUQdMf+KBkCsz673yKV7i8EbNdOB49drqUuEXltpdsv6tuXGlfGZSB
o3FnSJF3uMnjmRsyaQFzhFaA9h8HadtUj5ycPZ9moPVktaPWFWIjfkQeM4JnJzLB0yxxNU1xadil
WF99e54+871NdR/IKW5y2ej/Lx6qJcX2M3B4wy1oVo0qaM2aFzIv0FHhEukdnhUAQ2VlIIk5WbLK
Hk9xTGqQICjrYX5JfgKiMZ77pMexzzYrgaIqn/9JZ7GLhKOCKCEsZ5FSv2fGK2tOU2VKXXQVtYRS
cQmm1XRdfmYy6/5KcvMUqBAk/aa1qTWzveJybfrqhUTv5O8udqHQrE4xpbub35nXW40Jvo0qdx5l
mXJZQACbCaKFj6ZYnmFY1Yoa2cj9u6zlmu0OjvTKWtih9KOMaRfnbM+wq0YislGC6NVqMU2Xe/6v
cVQQQOOAVXfVVYYfjFv54YFXh8VtmxMe74v9jgutfMke7qSnvr2Zvo5ebBidwjVOqcLyreyXxm1I
Zp0CU7CFVWi0Eoz8HOjGz9xIZHrq5WqxqABwBG6w/gqK9QluFjdzoOKO86FBB5T/TtjhhDTMbujV
e/+YOtqMCq2i90p7O/2wJvMiYsa4p0FtttOms37DgkTeRt7v0GoTGEeBcMqJgzxErZbWVM/HpTsj
bVIdvERy8qkgd+N9a1N9TenUqwmVvYKH7+2ZjKSGCwPJMrf8jbsE7sAvmZ8iU/ZuxxoysMdi28Th
mzi/8t1289YKde6N/Ws5lOrAo1AIUz6LwtkqxiGcEsCBEJ05KN1ptuPnnpo4fXX77zG35wd6SWbL
I/4/baLC4NOv4fXv7OPenOxo6H6dRPS9Bxie9ZndYoQkE8FY7j3ib/xdIy7WeDcQOHzjHGsc+f0O
OEVcAA/bUgamWMXlwDFGO1by7hv+rBM/RryZDRztbCLliJxERz4V5vZYF0XTtxMsceW+KBNZNAaD
XOuDEqitBUbEYUFkJOW70rOprstkte6FN0jX0hf805254A5AeoJKLd5hAdmTE/hy2IAofdfL4hEW
xKAIls1kRK+WhN8ape/hKyGqr01ypk9DTU9L48ubnvDNUBHKEvXPNb925SSdK5b5+e4uFW5g2s4B
6NeanNKWG4IdAGoW+AkTd8gvbUq5sPqohM8r67PGIXjSWB08YRP16ugrdp2+2QrluhT+hzBI5hU8
11j1QrrYNvz1i25Qbb55lJjtJwLiTRN7xnOClPguh8QJWbWJzP5wEnGw9wBax98Cz3+LKdXlX36t
pRz9CGiiJuQVpUoclCVegEV6cgl6JL3XaJNxutWrVHMeQoHbm3ojx1f5AQ0VpKdF5/d5EBhe5pkw
m/xU19BIqJwEck8NQWxm1DJrZxHZpNgdqdUu96X3LNejxs1ogHoUXWtY+kaCj8+x//0MNzFqayiT
lv8A5CCvoq/6pVkJ9acyEdkmUoaeRdvpJPZFdFRKPp8rUb2DHOpiXUJ4SUFDsfQVXqnQOF3OtnJs
1GPLpfkjkVmXwf5gvNXrH0/m6XLKtE3t/19acnTM6qBAsU6ZV4Aanp6gA1U0eHQsqUbj6mDCIi8W
JRfpLMgiPLJ3YiOvPY9z8aF2ttfPK1B/Ac3+3PuiOYYgxhKitH0Urac386o//i1hquNS8Bj2g3RT
9qvIN8OiYJ7j5ZrlZZKUBn9XXmYdPu/18nS8ezHPyx2SANMuz4YgDbIaMSKpturkyk5TbAZhDyKi
g+HKatC9874yxbmeBsN6J+QzDfcNCaLFULHb5p93nhUKhwZX8JIGikrPRg46T2NGZvFQ+/wkeS9L
xLjcKv/Qt8/RGc09zm8r7iE7PHhu3Q42Dyuu1YxPus+zRyzNZmPXR5AkTU6802Os3KkG/Bpbrn8N
BGyx5Nh9aR42ubaeI4dcPADSS3Vzx4eHxv2Eq2kMMEd3uOLrz3AUT+G2Bifh8RMTEv5VGhMgx7ov
Z2b3dnmfvPt9GoUwHNk1TWdwqNP/QCNrNjg/H9jgfcCu27Zi4KqluredtTivy1z5q3JFIe82Mbof
nU9dTFZru5dNuARE8YGmuAm0X9cODZ7NxPiH3m//nRwupKjyi7oUs3lSLy2r6zyvK4IKmq/TOCFX
fuuy6ZHsuEqadlJ0l85ZjrrVpkboTjA40KHsdYo66A2nChWs6TTxHmkvQAtpdofLmRYx62IOSJxO
PNVtBDG+2Osb8lc4+19x+SpHhmeSpHs/qx1oeHmFmxv2noaBBiowkNWC4r5LVqO74CzUzfWz5HE4
VTRTqyfv/51umdmQIei9IOfdGR6hg8RlzvnPAP8jDD6kXvseaK+GAyDuHdRGIdx2r9PqDoe0RwlG
GtKdOK4H/yYyPXuehvxKjEWvEirhiM/GPVMCZKewF00XPpsXswtnhfBGW6QvS0mSf3RAM+c5yK3T
AYJAo7xvRBqmaj70dgNC+2xVOjSWEazNuBXmAQljErPf0kZGFqRjTgrs6IRnPGWZlwk0qzBEWocG
afEkhBFM9b4xIejKGX7iIzJiVjIRBelNU+3a7JPO6oIkFQ6fe/obpbc0UVTU0lv0iETNJGAYo1yU
TbaDDy7bXTqMb7z/EKibW/3rrsAYH4ILdHBhZm7pS7u4MscYRoYeR7zmI5b5O5QcJhrAAtTIo2pt
5gk9U6Fx16XzThHqSwoP7ft+dVbak9hf9K7kKKH0fMqbYxIy9aY2w2RwbRS6VXTsyPDFx0WLSVKX
Qp+P93IOh4+KwOXNgl/09c4sCpTyLjFVN6ftbEL9mffFfZG+Cs3Nlw5a/427JWzXvYDWDqjxdHz5
XmecX09v7TJagFskJV4bkw380/1S54dzAa2JIZcjR3EscLaNHnvDqBI8a+7Zn/NoWqf742SZJREl
cJsWTjtiZb4t/c9WGs3Nv2N+qxtGifGJt6W5QCcxZDmhzwm9SuMIrwQv2II4IrE4682kq2gi0B7e
QfyxK5jY92xa4Yimi6JVU06jZsPEcOepCV+kITm09UTl11iH4QHDz/Nbw/+z4TRewV3VCCmbg2pY
kFyv6vplAOcIUjrD31WTzBX26FaCPiB5Nh8GtIg8tsSCIIMBgulsLjnJ4sm66V+YUI/7xAVpi7TP
90I+DPfOFPOw0pHomxBwNwCuuUZvG78yTlxd6y8ZcRk3Te7K+syfFkgKj2NljQfpMmJ3V6I6V9t+
WHe/0aoYL9daqfBhgkg4oiRFwWISTM1LePaCa6zMMkat+s3HjRprJoio35kZ2TKISVZOoI5/wKGj
3mTpxyR8+nN3r2ZoqqRgi9QJi3Z7llRoymiPl3/hquKrMxDWeK05rwbab9fRuAHqAqa9izU49tDy
N/bD2iVisVCPegbbKB9zgHzVM/r6zYeEinjkrcb1WduuoQUuqzF+OLe4sU+8/78+H2KU0Y8rFYh4
kdOm7GyvwuNrF2VOEa6dYAJ6DTS0zDK6nUMY5vuqoWpXhYoNoc4DBCHfJJ1hWBrk9OUww/p3zq6C
PispbU3xx3Fujqr1Q4QafyhlUffIrg6nRxD4JUX1UTBu6A9OPWLwySRCzcD9k7R7+0a3L46fXQyT
8zMUPOk0nRPN5LoISXE6niHc+zfkRSGTeGVt4AlY9nrxJ8TFIY6LpHjg2RcXuOSZmPCSCTk9M1Ex
PgofX9pKAuG367okyIIarcYhbreOnPa+KVeeJLtQOROvWDAzsMNVjfYZ7Ez2Phqqn0AEzJ/vzzhk
fu12f2J5nF57lt3jcetwz0d5x/8jDQvBpK07suteBusF/iIfCGcpZ8kGv4jldYMNAurVLu5SNbA6
l+/fmgKkSyGqvJAbax1ARfg9jcQ6Mz7crvfGhFpTqglWCdwUUiUV0eUxSkHYX1he9M8XgRbAfvFN
tiLt4+LzlHzmXDfgxKRTAHcJCwe1fZt7dNTNadmjzcntxMz4BZOh+xqwYHpj6PfKcV8bgpZ7kOKc
iP5V36umcUgTvtNIN6wmiOmeFWhbd8v1dNcswrrSwGcO4LLxAWGIg74uc0HrN2f7HbN1RH1BspPw
ofeB05IJev6OeuYwHFy0VBGXGbNVJLHr+/ejNEGtkbguUmaGXLikjc9CL3zjvyQmvHVTBN0iEbbH
2GIlos8mYeg0lsFAj1/86mnz2w0DBJv+e/+VDNYyPNQahaB+76I8f6haoMmSVBrJW43gikhfXVDp
+/aXOwV7v7JWUicT7v7CljRu3/f3H7bwJg1S7Ykd2OQyZTw0si8Q42gxKUF72uZCrxq3tDENQGLk
BKZZnKws/wv11Dbz4anLf19P7qkp/EJbpOW/YvvneqpSNWnrcVSu0XTYN1VFKz1Rb49YsU/k0o6h
1s2ofvAwqgbMwZVIRTjnTudUG1TX/SmolXmh23tjLDkqdWIuyUCDtkKCt7WRfK0uspzl72uDpIcg
DcJWzarQlQhAaNs1y0Xgf/VV8NsiAytDhvnqSl3f6GwLKP85q0xYJC2e8pMM5Ft3/r33yTy/RTAk
WYonxBMr2ySKoHVDG+P4Gcw5kfMXRdQD8xdoBO+V9qQfYuzk4lm9vE2lXaUheX/JP6jIttrDHhMQ
ltW+yV2gEyp21I2m1r4w6I5wxvuQYLYhe/XwCffxtethv2zUp5RXu8DzomLJq1L4gosBMjl5unim
LQzSZM25VGyvMtVQEqCRwK/LjigXc582BT5vK9+dbfM6mbkaIRNHGqf1VmeL2/2wvrPvURV0BxD5
1uLrpTKHjZVN67qNHy4zma9MKg28pYpE90/rWW51BOd0XNv1Vo4nosy1gvXNQsJrzUZRQs5L+SG4
ZjIjtJ0q5+cNwevq8GOjHQwc0rnsNHuIy6yKlMpQ+6uIhSYujY4H6C+1FT52WMXzSApIj31lPx9G
QJ7/pty6dh+a/jnSLmYMjHANAw353bwEzMUxgKojgmoLvrP5I4hzdHAi9aE0jrtnHfvgr2hRoJW8
zQmPQyYNK1peinY4gKfRDvNrxiExULpg5zUzicR2RzvvnBwhtyghqicUshh7n/P22swQxclmZJx8
S4EPXlT3EhiMLznfnTGG33RuEqNxWbzf208FoQctVtoTUQCJy3e6VahjqpH91g/7hC/y2TihGT1P
cEAWFp5c61bqcPboNN1I3sKg/XtzV0ve1t30O+fIkbYhEwO5CMmihc13e3rHIKi3FMZ6b6MeONmi
rvh+3hCcywnyFuuzyauEzZn/+V57ZpeEj9g/ENfLTFRt5Fh/xTybRNUvKyPMjEHgJr8Vf/4djPlP
asp83LpG61Yu+3eoHQCUV2x2JakmTtZZk8LLVZbodAiqHhb1A4YFDs3eM22LgqohA+STa44rzKch
n4eceLLV/ajgb51neGAT93zQ1Eypo3qFu5Pm1srLiYXVmSE0XkUDuXl1WAT8Gg7EeOciey3HC9Ua
ryjs7z4bwkHF4lrp92kGnaabeb799F0/50S7//UIyTYoIvvvZ46yybWapOxPhaCNW6MpCxXRR5VF
SLZQ+BMiDspcR6OG8JJHaG1FlP/5XFZCQkkJzUlEtB8i6qjZTRsUkmTwl2ck9uzDZihn01/5MKJD
jp6Om8EeSEtI7fkcw3QI1kd3XK5FbxWt5e43Prp63ardu5ERvA1L3Hwc/NWgFKV9GoicCpSdD+lc
GjfsnPWPzCYtlwau2ADp2Q4x365oT4clYIb9cltzIM736cU1unj3B+W0XpKqRFSrDSzyzbB384mn
yfiBCuKWewi2Pbnhkw5krYy3GMAiAI9FCDnvNz67ieFdE5Q3MK4nYvp+2sh5fJhmbLC2/+KopBX1
mcHcLXOTyLFighvkvfuOpuKlzBQhaiPPMxgBVE8xjCdwP+OYBzH23FDwMDea7ddFA/QDPm+pqwVa
LnXj00ibc1HIx0HB5ZlSQ7qKNeE+1ZIKW5Wwb2+G30ND00AnvJf/c+8jHM9uS/IKX6Zdh5S05uXw
GX1gFPr88rBUNjqYSqRnnuPDh6IKLMC5DTR7khDzNKrXjn6UmMIh4zuoz99DaYIZcrks0qaL1wJO
2xHmr87cEvzVaI9z3P6NoyQ7LBro4hLKyO8qZdUbZ4mFjF6nvx8XvNxKgEIeJvL79oxZ6vYGx9fV
qNDxgTt8/5GNCJnh6o+M9I5wrGthzkaTXzK+xh+ejlUW0AAY0G3289CrjaaKxKsQISfPyg3RTHo5
fz1LI9qnRFWoH06FtEZWlR2HKSCBr/6SgiBSVQ7AjLvF/fL5PC5jTCx/PeBfcylJdTik4ndsr411
RvJxaJD4mNpRqKOvgwS8pS3L1svZq9qPYeVjyPxp6nsIycG45HrjKYKIvLGvwU+aAQYuAEX0mBcn
p96f6IcCQbJL7N960uKaTCEDn2TxBY01kX551Rrbq124wNdbYMRwpluyZwAHzNG/6S5EjSaHMXHt
Qj19fphCAsULhKLy/oqlJZl3Jhug0scGbv8hpzZFqN1APgKun+5TNlcGCckT6LIv5Vy/lxjJIzoD
IKuUxydyCeA6MSZ1gjD2DrabZlCxtDIxrsNt8Vx9ZtYmEa37zLWAGVG8p3tl5PcUV0V9SinkaBiz
5cxuekSVFRgs+Vk49AvNagdoiueyg4WL4GN8uPAYotlb5+mo3tOTUd9648e00cDLB+JCKosZjHsM
kL+qfY87kpC755TJNLcyeQkgwceJdneA9nv7bGXimL1sL38f0aiKtXj8fAUUm3scNNGtpHvBQ2BL
9Lk7Rp0sHTa6+qIq3L3jtDRGNgwLSWsT+j5nwy1JzMfZl98Zl0E3VSXuuKZyJqj0fnOPk3YX5O05
czZdR2CD9+eUJSJ7fo4GTWxC2YmgsFUpch+PsXivgFDogizgC9ijpCZFItnDvfc+C7viMlWt+Kqu
W3mQyEcWmHeAiy/UOOqzy/scrZ1I1CT4BnbM7AOaQdMYyl2BOHHQlOUN3FFodwcxUt2r164KMDEX
1uTinuzVpyQA3YbF395zrSGD7iksivkfrwptbG7NTxCLjbly0n+sCAb8JVZnxuYIUNc6aGI1l9tx
zImmulpDMyOpsRy5Dhyo8cBl1be02WnLrSj5NC0M3+u4qikNmuMKnwmarZmhLcRQwXLURZdudUce
C1gphTePpHUpC3OwNTS/AiIq/lB+CwsXxZsy4vNdmFMUWRdIOSPJ+Z3jllOAqUnBsKyJ9yTh1gCW
1bG97EFZWdI+yoBsFtl/vyaGHL2vn9/PfIXVI/U045dpR8mgZzOkC+XVsPTHnqpg7voRYuB0D0y6
a+zfA3Doyvt9ir9ZFWo9WsWyNl7wacbG4/fwWczDhlJKAWHheMua7ckJN7yfW6L72SvTaSBhOiXZ
WV5yWQo03xITkIGka41xRRsi2Bylu+TzJMZnAj9CoXNPowDmptQfJ0+pIY6I9Oo4GFBJn3fO0jk5
pYmBJt6S1w/YPmwoLh+75IblNLRZcMfc6cgPcmSBJ3uDBgG3KzaAz/OBQVv3/eEEteFiKgzGeEbY
/liGspZojgdboo/kxuoYiIzNOsPAgHHbLzPBmVUw/Q++d8o7l9iSKoUYwMVUcWCHfsu7jlBkUSR2
BwtwXtLYm7hIh0J+XAj7dDdGpbbuw4czzuJ5ac6KxTiJ3CSVUMlBPaFU1450GvN7voaksPBtGXlK
QNj64Ot8oilB/JEHq2zlMeVPue+pw6e7zcW3Wlrh62q2fErTJrGRvhDblng9vQ7HBcFqt513wsMh
BjYqDb4UlPg40EAUXXqRvKbUr7MXxJAehf6ALA6v1UB6OgC1fo0hEUqbyeaSG3kdye1eAMHcw4ee
Cn7nA8mpUkad9iG7EpW18FRDx8OpSIIcMUS7TMyC1eT1L+HD7YQi6zdISQOECwV1JrjO5FxqZDaU
vwPVrCdGrgX3Kh69VJIfLXo1YPGSG7IfGSvw0TFStzpLn16IJeZeghoVr5uXtmVpZrw+VavRyltr
2MFhe+tnLhbFon5apLiY1cXDw5KmQc5HwvAxdFLSy2709FFT1YuKPULd9eUOEq4Y+9Or/JvA6Odk
yf44d35SMwNpZ6to6186xe45lINc2iPXFGjVO2xG4T8TxTrjb1hYVEwwPi1Ja9ka0Xk8YEPZ/qzo
Pc+umtaYP7SLsLFWzCf8AWKL0k6J6bTjuVkpXng/YYnokGaH6F4Kq/zGIKIvAQ6dgugbHDnOd/a2
cBdoCIhONNfbSV97bWwio6waA4Il7SObEMUTHT7ZJOtHeZj+1smHUhR/t2GZSnfyWL5q1fx/MZrO
+TJZ6kCQGyvUzSoMvszunM75gmKsCDfDkKCsyIwiUpSuiTnFTDzUssFvSKyzBJlSlRG+dfT2DycM
215ff/1/7l6BENpkxuQtA1UhzHN1f4nFJSpSqqASGOQ567QF/TKa0ECk84lXwnF/tQI4aYWhoKTl
mPuxhofv+o5Ljmswv0QdHjQgwOaILi1TdlQpQ5qHuDf0xP8btgosGianRQLpZVLJpOsV8rFQdWd/
8uHcp+Mc7Z1ncf28pVldJ7VultkY7TW/tSVzuG4t6g+mOwFGbOfu77paq8xnydarfKkQq+wdLZCy
One13wz+rzeUkfYC7XYNe2Gq7VXq2VvFuAr/eQKu8Wi32nw9iVV3llUnXAXl9WZ25sibjTXd/Kkr
Qh01EmQds5hZwcf61r2SqCp1Xf+biDikxidCgCqF5sGVlwiaUp024iBPBGe6wtzq1iSf4yHZDnJK
RtCjVSPPGCJSpXtiEhPc3ejMKHmuwioLZURzIERaOBgiK2FqPwmENQsdyGRAQOtKm6cX1bRBQAwn
YAehPs/JXlSBJ26Lr48svbNHoqfDz6PuXdkmFLi/BFx/9oNkIh4NluwDiwXPx+BkIn4pdabEnYoM
qkcik4p/+9qmaj2bEJm5SMslYI3+RnY5uWxAo8FP6M8D9n1Ffqj1QEcaB49UlxC01ECQ3G9rWKAr
7gzlKxJtkPBunE4n+L7PKENOwi35qO1qNfEeC7/UOeFOfDimgGkFQuTElGaMGeVtvpy3G5mBjy1L
8uVdYGjkRj0Ki7U9MAOXDLzDQPx4FXe3DonsGdyrLpfKXoHPPOWUmJbQp52CIFg+m1Red86PSOG6
suI2XvAZNLKsflq/iRXxRausXrLdG4aOYT/YhmcZv/p2fzQnfGlg7dTJcoqxcahCUIbdelWKKf//
03o3DPZoBF411jvXW37DF8uXyHp6QrKoWpP/1011Kwgf9pRV1Re3CVFTqrHc7KH3TWjpkoPupoZU
A9Tzs4cAFpix1AAAoVOPuA3SbZYJ6tdFURL4aOpGHjXhgwXMHahBVFNdqU6qsg3vuMyUxV0zW8op
IP7hpi7VVODGLmpIbjF0CzCFxAZat5VTcwjhgWH/aztXY98jfXoTveq+xN/Je3O6XUeYYTSce+2n
rZFl/W9bkV5+vtxGN5lfNu5ePmiJcYFwtCjxPmbk36bPQFyjo/3hWciXYehz+zYJ5Stm5GJyatbG
tt+9hco3F9TC+b7ArSKpLmU7iKWGKXsOYcpgRyS+uV+lmRW1N+XxU2ofRzw0E7SUrci/dySIU7Mh
LcfO0TuE+z3qHLVoKgjcIxQbwmNTBdC8UxWB2gt5ggevzAQe0wzZJTJK5dE50Uwv5STNft2KvnR3
nydO9e5a1zG2leqbVBpaQmTAhZECuclQ34iiSfUvtA53v0b31o9XkDQN30sSojqaNa2QCeBxPBGc
FOn6oKiqF9BqkgTDs4XPnleP+woYmTc4gE+a5C0x/WJ0fQsyvKu3vMU0VQ+wGYhNqL5Bn9PnSt4n
C/tI7PYu4nVAZLDfFfl22C6u0OGtmqol3bf/1gRsrNX/M6yE/ea14xJFhc8EWVFyKl2uSa53Al3F
4RdaZovmVQjGJyeq9f8yrkIVs2EKw2FLuGg6FrdzODA51wL1QqFCBBD4Y3RsiAhv1HizmO6CjM/8
ZnduRBmntaPG/a8b7L/xcaFu6gAmTLDzc36QbJ6hYHiZgo/cGufq1pVULqYzVsqh0KBjHh6KfZkN
11P/VJzxucW86CKdzQ3efrJ7h6f0VjSqAptNTOlRe74kIOjKNWTbAyxXxVJDqLde/2eLx6tHs6JX
UvjEZ/5jk7QtLBYV8h6F4BEkiLC/D0byiZ9h7L3/rhYGu2KwLbYJk3eAgtzCMFWb0DoEE2SlnW8e
JyBcL46k2W9j9UeIvZIoQXLfOybIdzelda3Au+htpP4tpdMAN6U7uBeAzLJBBfVKQX3bzBfzqEjA
GzXST1yi8z7Hvf8PSIm42PPiY232PLiD5Vkql+dfenQgN27ZImPxVGhce6LC3mAYcKMj7JW1Ldjm
DWcTrqj3zqpZ3zRMyeIaHpg16XXFf4ygDC+ZEgktWjOGam+Io2BUjuMcdNTjuo70ymdX/wdOati9
II8f4G8kpbXU8fVnSnvRWhkuXisECLsrmyE9j6VBF3f6J5y1AYQH6wIZp0EcEviKqbEzGhCKITl+
nRzKa73gukpI/MEz7M2RAWlT6qWPFsD1j87pQBOSWCbP1M9SMw0SZYIau33653r+oJEMUzFFnwIj
2a9GvjnWcRU39hS2FOtjN8/WPoInEMEh2BPiNeU6olVKMAiHbPsGkYpq22EIuhGkAXZg0OX8KJ9+
QyD/oq+RB/6dWj/9Kb9ZpyKR4IFzkcNLSXZ4PnZ1BQCVm/edQLVHYD1KXGxzNhlBSNjngE9LHUNa
i3hqd7m0M4NsAfaskvWThYZ8D722/zzLqe/vv7FtYHWEcRN2gnZevT53sLzizAipT9fqF4gcbpDR
Vugq9UV+tqO3JkflxHNHy7bLFsGmyakE45vmQIfIIhsh+ATvCx3elyhq0JtyJQuwfTsUHdMyOL/T
KDZLRrvgdrSoB/gwBydTOEbynahFRP6Jxg+HX8iB+w/ghywLEisKnQ6YXNIjuL6GhcEJc8XsYFVv
BUeggSGLBxQ9gPE2uVdEIImYDtKUltxp7yc2DgsdgEdAQkWekPCPrSzCmKZvN8V3B+ibg1c+fUSp
/5IN0kWGE4ngwVkoS7KxJUQ80/eALvGDjO+dePtcBLCemJBBUuD055+6YhsGN9O6Tw2Smd1fZSi0
9Fvwy4P15onVEn+PrTil1nWuknx+MvzGy+GByS5Um5luPJFc6W3ntjBPDyBA2rUSjJQfEBmY36xL
nxDsKnW3UQLfgPDgvmXWb0gFTYtYw2jwjgXzePKczPp2jYcLt79tWNTYN2QaLNgKc+uLRLmACT5M
lTRw0aPonLnAmjTdPgoqpL345sNxwkWurSHXOC0VVembD14AU32ojqpv+UyVx6E+2/tjNjURTrq4
6OYE0FyBamwHJQtfMYmQ0yZBZKAGOOfMzX4sVjz6YeSazqnpQj8ERgYPFoEMLA1y1e3EpdSVzoAt
sy2ja0BHxIMrzphYIDaxuZRWoASWtxBNYa+PN0aWSqg2juQo6XpCQ72a0QR3bpZcIaiu7UU+vBRJ
0voOUcjwhUjWZjGRGdRHapRYuhdRNLDzZgkgjNIJF3vwpSIKTZiB7VibGkLny7d5TH4/yVZlRaEd
fBe3CtLItGFTq+3uIe1IckucxLh7C7FfAzcmHFGSVhcPN+lnDZx49FMg7VqMjwSAy4UmdqeCsQg6
xC45QHbb5nThSqG6m6D95ptXDpubkG9YOIeR5N6BJ/8YxujgWix5RP6R6g1PwyRr5WxoPMrGbwV5
RgR7pnbTORfzogzrYdfmG7q2NTCpUYB7ZqdI5j6O4djbfcfTA9a9oDVfw1Sa9Ft+VDdtEagPIcNE
h4cWUIBs5fVFA6aBNYMl1cUFERnC1ctLI8ztAHa6GVzCPvuEBTSRPBPMtMdbJu5oRgQPjOQUYgxd
RGwtdJgIDpzSUTEYqtQD76Ic5rxdvxLDY0dOEBrSxHv4S3guDYn4wRMk0/EWzaHvbTbOVQ9aETd9
YVWF05aQ93uNeEwngdTeCVWJeRH/2vRa+1aZh6O2DtxaElXqqegcew19EVRyOmXDdILRJRkoAiMN
hDrhWB+6pl0Pa0HbRll5VbBTQn6Bm0TiQdTAIqr5kNYnOr5NeDGPUMvH28ZOkd9NSdh0QeuJFkTx
xixrjGFuZFsKF88pGUy7hDdGEHyfZV3hNB3IC613adtg1MTBHmTIfV1Ren6X8FduykFNdLHHiB8x
NrdTojUykH9uHyYUWNFOHvHPsdqzL4X90zRXvAigCkBlP7ZXDPOCvFpImRA535kUlnrA8aeiNN4h
HuIc0swiTnLDx3tJ2KLx/3jaxg0fftD4ujNg7eiTXeiIDk2W8ymOT9bxqgpxf3wBPznzx7WfYONG
FJLguoAAssf3tGcK5J7xd24yt3LFG+3kF4FV03fIwYYI3S2+M0bgUMtNofrtPPP5h0vQnPhFy2/9
tX1p8hIrz0n/1wSG8KK9ukrSXlTXuXB3n07RU8KeWYU9PMVYyYQHzR5jFvO+PiVB0s/TksaH5iAS
873bpUVT+tuEVzGGSHa6qFUZtLt80ZHMZ8If3Ta565z2eTVFNswJvO6aMm5f9j9zCCuZrorTC+sn
7gcJ6EA8WFFVCaESTx+qx+6dmhObOyFo/aJlxDGjxgpRjeOxYpUHCLm6MvMDrG3R+R2zBYfnMi7k
/pw5MeyyNQ9TKjxbXHv3EC2DxUuef25Q7aw32F35GzuufUUB+hT64WyiHFVd40zCyTBeZyEYR1FK
KmeuCuHdT7YUkfHJVIgnV1Be5s1oy9YbbHIwjNNOeyg/Q5yhDBkAlBuTaQJGGVpCNYmREooJISA0
0DI1oeJpxJuyJYhNXtu+aWzvU8Qm7pNQbWv4QS5BrVazrzlLdWmzEDoB07guSNmCMW9OJbk5zuy8
VJZ8pbx+edwy/s8DNY2OFCZ6LY/6ikVEFciMpmsJYHo9ObqXCsBKt7NJJqA/1Rxx1U9gVwINrcMj
I/KFUrz9o7/7XwUzXQn20I13+VcezxIQnvkkXz7UipzCeQe05f0JyAtARQ400WKgg9M3cvx1Mxv1
Y2fm9fFztg9zxgEX+dd1jpWdBs9lJrXCwHfq8Y3HFBWhTvAvZrJXMtJghQJZC9GbOP5NnJYWvG5y
TYN31ar/89PjI5GmNikFZ8PRtutLhXQEFCDvIwuWbOhy0M57qTDplx5lsXnHqImjc78UiDaf3uUW
yKBpnLNHWlvU0EUs5KmIZL27VVmGJ8EBlyyuFuqaPpDyfy7kPG6SL6CUzsLNCdr0HEV2d+jHG6yJ
mBCqs7I4z9WaUhFRI30hO1t7t4HDQ6Fo5oeMPWMVQb1Emz9vYZwZ6i5skEStWupVLc2JfblI+h/I
Wqu1/tssDcjDBO1rjeECr1JTHmL8opd4qKQ9LPAEsAxS/P/wGzmd7cxONZYGc01jjlOkXrqvJViX
IzX92eddimP9n+kVLk3TvHe2MOZ9fncnS/i6o5+JmzsJIT6k2dHIMLWx99njgbm8VGbcqU2h3r+/
LuBq7JLDUmUE+AW0+IIKuc/hGD4Qwe765O2hbJBhmTAMM74CmNBjLfPeEIxHZ14SCWkV9MOP8zHh
g7DEtQTWKlrF4iTpvXLg7H16umC72o5m12Atng40Wwd8v2MwPchOtNuWVVY3oiMcAqOZE+qVrAbk
Rg/u1E1xE2yAIRGAo44Zm1rmUhTjp6q1nt9FSepgX4EpIyc3y1oFvjCx1/UH37ZvY+biBGltRZB4
q7HIhrGJSX3ZSQKPLGwxx0qHIogFpwgf+Z1/tVK7Wu/o8nUcNnc32/4btWFvua/vUk37Cqa32f7D
OLOC9tBEaXxJpxxCC33jeV93F7y0qrqQ2kZnousQK0iwkU/gMKSBqPYqcYvKy7T8nklJTCtNXOMp
4ORdv5DjGxviVKTvNvJsMNrAHbE2i7+R1nP0/vnzi5vN08FwBo8MDpzCLrUmQBGcFUt/3g5OUZAb
uZy4FxHU91xiTiic5EuGH2TKCmjbVOfEzP5f9u+KyrWsWQDzt0RLrJw+1JOK5pKzmRxMoyWPU2iY
buHX2ZRqrphcdboNWPr8ud19Njox60sAaO8zaTvoSDNgFKgcJDSsMyT6uG6sx0SlgOf1UbGrcLT9
SMIYsNQX+PT1RStw4+kLZx9uKO9pRbHRbQjcZrofUu7h6+Wlz6P+PPT59djdcUEjEUcxLtxhFC9L
HUzVOzf7kKhGYjNbFkN7VArV0LLqeIwJPrDtek8MDmTTyDzbUuyJFcUUr1+gXbVLDSMTFSfeha/o
2A6v6Jif7Y6U0Mfr5jzPAfkJM6FMxHsZuughITOzKC7GegHt7HpViF2FZJ1EI91sgSNBtRv6Ad+g
qpfcmO8yfY4uRPjq+GYBeKR7Eo1eUeZACGoUycFNI4sbQsNEPrfV5kB5DQvK/Q85STgLMkQdkmSK
VgWp79gg0XvykTHy2VvIMnE03qWdeZCQbohGpaf/X8SiJ0cpqS2TnJNNi53KyIZfuUG6O8eLmuIl
XHqGfohxhMEYQKA1dLbC4DIbn3WUoAG5+wvrcWhdaplBj3cH2HdYiE+jV3+E7gChERTb9KDdLikk
MxgPqs8tV2hfrzUMwz2QXUEZdBsyj8jlAeaUYO1vBNnGyoUN+TknOM0tsO1qFUqy5PlU86kRsDoR
Ur5zzwPeu7WXnVmEVvM9CoUPNCEuBcPpkbBxicH6xd1zdIMfeftnVJyojbMGe5JryL+KasTTtR/K
4NeUGH56FLTagbekrLPYPXDVZQ4ReozMzmGvL5MdfJrKFgLUv6nyHMJXlFKjaPGd6OlLqCPwOkt0
RFxvU+6hbc0ISNzvtOPCnCNb10T6J4qleUdwJEYsWSTy34wiVWAYDoIs7f/cwoaXyNdNDY+wX1+8
HV2gj6CpPOtNqI30/jLCwhpvhnzlcHgkbnbAKQRa09OhwOIDE8Ukda5FZ/afyYD3MjEF79KoeCy4
TVISJg884AjWS5Sc57X9KFlQzWj4O0nQ+9KxrzmvUyFv3Nkyc+LGYWz80JyiGGGvAdC9Fwl+NfLU
H9nNiturGTaSwk6n/OFmi+Raei0Vs//B4aMsiMKAlbZjV8yUbR4+ZyUVt8cGh/zsw6ueyD2Dl5V3
1QqrDIUw/MMDFuK8aWXWAv/jH//AM6yxaV9iha51JrvWfYuvnvbtFxozK3LJMeSK1AnuLUO8oTJH
RtUL0FWxgBrA/eGfi3aD8w1FD78pvHkLNiytCb2I3dxhKV1NDceknA6dCx3gQFegtzMNlgbkmWdl
FG+sPL5DasGkmipb3ZTiozjmntTELrnW9dJvHlHwNwiNrOafwV1BgQrzdHM25bLEKSJ7FEMS/hPo
s3GdSQnnd8So7g4UJcEmTZhBc/vcBh1hTBx1ebCtYUd5M8xOS5vNzcSOUCGT1GUArG8ToYFp0gUb
vf80xTdKoioMiOBcWvsCbpoACm0jVqP8dPnDgOum5S0MywRNeMou1G9uu2UhJkmQ0GEd3qVqChtg
Nnowyo6YD0ABzaethW/Kypz7qSjbMCoFHuh0a/Sy1LDP1Vrejh2edNsEtsJ6Xr6Nvln+qgT+Zyur
4jLNNw93tIF68Kz04S/3e1BWNljrce9KxYJlVHyslOPSxTb+7CBWYB6Ny2syByni4n6z0ufFBRB4
zitdBBnPbUxQYMA3QOFMif5nXHpEJXs36HCVQV8GFvL7YTRGNEM/INpGx1XQoRKa6LJOkg65meJK
rP+B4fXBeOEs3aWW1B4Lz8QvUxEdRa/AHqMVBQticp/Rimrhw3LRPnuFX9tTeA+uzQjbx6fuM+73
iFmxx2ph5z1PYE9PCnkzViwIDv8d0uwyK6l+AexuCy9S/A8nlaP7K9hhsSS9RBzwAfxmzdb1Zz60
7MBdVxmt8HZmMtF+rPXmnYKY5AYXoqT09Az2kd2k/9m4YC7/m63b52//Xxc0tCuYyIDeU/4vWOgi
l5EPRYngvWEDWCNWOFySrQr3DyYKo3i5AcYgvEbN8LHqqEAp+3pM3+cJgdXVwzGpCLYw/CtwE+Ae
uVdxZuK3K2bY37OH/e+6QVVIWwJr09OMTIVKb9LErwM4vlOToR9PXYkeOI62bHSDyfMWuCnUU0B/
s7VZ+FNiUHskXs26p/kd9SxKqy/k61TX+LgYawwqhBpPSIMnCd2DivBNK9SAHSqj93crwBH112Ls
wsp+kEI4rb/AAVIq7DmraN+X0KoZdsQhKbJliEpsVoGjiyxg+hRm5TT6VSvVdcR88nf60QYCTYnP
B8AoL2Vw0QKvmrIsPPlKMb0AdSZ+LvqCSIVoQAD9hJnw7F9I0rKW1U+2MapzAMHsgK/+UxSBBLzO
+bYaTkosF/tgyNuzQ59SUo6lxw7zs83q1WpBMZssdIg1PWkWrMyndLq7sRQ3/l6ow7cxDIc3DlJf
twEQ9kPvH+TcrFnOfSqt9eZUtRwZML6+Qst+vGp/1s7VMISOiHlL04XNcZR4E/QseGrR7uOVkIGf
xPfRBaalwKrQQl3Qj7GHib+prYgywI777zwTDiJegbpqftWJvCkkFZ6ioQijNKEBOoMm+GaLZR3y
CqfYJIz7OVduQ8CUVsIlhwjhdd2VGEnOK32ruX3nGJuj4CzcAmfQpNmvC/vCdzSp1IddkXZwPwES
OT1NBHG2D/l+DSKiXvK8h4WjHRRm25X2faU6InGve0vaWP1HFGUEwZodzBe+m4IELDH2CDV6HT6Q
smrCHGVwCv/ZE8F5UHCEX8Cb/nSoWfwdno8Y0H4ww3VW4t39IafekQpuf5RwKfu4DeS2HPVLIVMF
XTZN9Vvo3AZGdx/9uoddwN7mLxDaN6s6b8e/rnHX8fEHqYubrKPUxnHo5hatTM/BnraShwNtoFIJ
JYn6F1uqS6kO6t4Uy7aHOMG9QbyBohX6cHm97Jj9f/heOB5lTryu0m7DZCILr842PvzDKM+hz8OK
YtnflbNJrMlHXJbPdzL1U6mW7VfFVTBLg4sTz0Z+TqF1crjh5dL9UGeJxjTTnZmtduPsYclxk9dL
WsaMFXB04M8NohY8C55mtiYOcPP0e4c3OgOpJdc4HhXyneSUbauvLIP02Odb3Yr1sHgm6tP69hR0
KHM1DM9jOb4fPOu2ksLsYXEIsVOz/JvI4VzeAUM3nKFz+Zo5+lSb2OLe5C2oTdNtKM53oFXP6F0e
IO1q3RNVQjeVycSWhzZNJPRdbZTfAuPoAmXf4nikcn1fCmO1OLSTSs8wiw42ASbAWAWdASx5dYip
3SEzm++/XVwvF5PCQGU/QyTUDSRPHG6o9rWBib3e2DMRMnjE5I++xBBg3cPg6gBHtY9X/XrnrHBm
jVPhdyq7O2nrJoJ2C6vEiVUdczQjz/pFBEWJFkUE7ukztydBZktqaYDdmvUQB2HJ4yFUBhyiZ1Oy
DC6Jpj466bzi0Y6INPJYnhCRrMxNU+meIsvPkxV+HQozksdUamrLxaHMTLQrpAB+hrZBS7Ae1CJ4
adBARg6Jf1kth1IIxfztXN6k0o0pNIpmrcEOTuJ6S0NwUJaPwsEA/CFOAFiOr6kimigt5Occ2fvb
ZbFSLR10+RCBIL//YCtP0IJXrqm3p7wDcUQ14ArGPLEzfeobm4R1JcALmyNNwf4kxGkgb38OW8mD
0HrUbWtJTSIfuaLm1AMl9mJCfRNonpq3ylRBdvlPTQPbn8a92CC/KL1a7aAuo4vDx5MdN0yaBnj6
sLz5heYm1vd7ZDz0PB9a3DWzGGhxHLSoBzRtDMoI4txmT+jnwJHM2I4cmbZeJ7jSDXRhGD7oZrPb
O27K9Ax+PHZl+63Oy06hnlKQlnwKR5JBVFFZcuQHBJvWkYIIBKA1LZx8+HBxtV/08rPDBKdChTc8
U46Xj+5/+pEEuP/fQuwm4j7cdDf1SnbZyLVwuu3T8bYyIXV4zF6jVZlF7FwibpZj6YEIXeME5ZQZ
Et9aXeCLCpH6GA0cmbkwKHkwmu3HCaot48wjUvFydBlG9vaKDZagn2AipZB/plBi3DZfGD3j7Mic
lL/dHJqNSzlgdM0tePxt7jJ99hJEVkSypZsoX38Ega5MWtEZKfSLIX7BaoQeyV4YL8yk9tSAwkDL
k00sbCsHM/X4gCh5HqM7EDFbSdDAqxWXvFXF8+KG/tBSNU9ZlJSZLTqpHphDyzLDLqnq49na0kDD
AD9DhDMXrF/Ez7jl9tyPUCn/ZX3BIINzk1ywvZb4x2nFUDtGZzLEOzn9qm4Dp07ZCQ6mRmF/7goZ
ybvwB3j4HfM7wlnM5qsocwc6A/Z98NnMZRH1voYlHXoQ6yGRIDIsZ0Yb1zHzWdurTM2eDvK61hGW
eZXUZqOO7Bqc7ezHLQktOvo+JUUVp9QxcHyX5Q8f8tzPq9gs8JEJk7m6CKoDCGzxvs9MQ4KSAebs
v0wW32Bu7ucow0+fIZ4W7Ox00Pjdo2HvjW0EioFH0ZGUtaxmxDpSL7zIhkMm/LXjStTvrhMOuiky
vxrClpyb+iFXcpT9vvhyLrLHGz8+L1n+AG29SWhmBZjenjnjQmHH1J+t2ytG2Z2dpkQAj/bhHK19
iwMZAuYiMmsKuJ753oprirI+UgUfd0VlERbj7mnog/XFHXoWJJ+eMCs1ODsDyBtAuHKfUyYQx+zR
NnM+UhuCFTSXDu6N6huLj/TsaNH4B0hmHOc3SlVh65IY/766WZxoUaUpAOu/xW8vS4JTux4+v12o
nEb88nTqsRcuKCe9BOKY7Rh7iILOUjUKS9yN1WJfy/vt+OW0UQFkg43v7t3Y56FPpShYMuWIufoA
lHokE6Q/ZqzE5aHnzVBHNCH7upNDVGVvBcqNo63oxbg6IFxdJR8kvLaoyXnteQnDNIxKbFjZIr9a
MIeXDIhTd6moqd/NF+P//g4qJBeQqV0zRPyu+SuS31AOAOXTLxpEZ2PAbhXP17+MJRSTd3FJXDUS
t3YCX2t6Xcjk5G8gLdl4pDNfE+97caTySK/Qfk/Y2jX0KPoTdLUZkM409Rs1wQj7nIEShnJSuhGg
xnYwa2uZzelIe2MWZJJgBJZrDRFSHt15zHr9YlPnfGQoMjxEkGGPCnher/1jZdirE376UGtx+K7p
HMTGBcsU+GXZSk/wPcJKgf4MsVpFAXETv977ptXUVNsbWK6DBcfLYuMix+0UbfkhZlObGev8etEb
9T5SouVbKbxp20TZFXWbdOKGxga7KkE335Yi0CF0GLeKBtH/LpJO9nDlJi7pdk/mQbP6kmLuv449
G1FZ4yMuzdPj6H6cvLyNL/ETMjqho0aexv61RrENpBppb3i8o4m1j0af+56rZN5s6B1IGhU8mCKc
/7/rCuIN+LJdv1BwK4pjsldPVRXCI+jsvElv4321h8MkTH8w/zlNmLr1Af8hDh6Wq15i9EQ/Dc1m
a9cLP8zxPLH31WYtK5L5165h/s7ii9+x8jmSrsNTLTk10F9am0Df3+vHCHFzS0dugavAKUhJvx2N
jagwxMvriOlevLEcUnM1mS64mwV8kqkUI7t3e78eHrjEQDmvmUPodxueKsALB3GFs1mDcMIipSGV
tllJ7kyNDk0KheRwpvfFTKsD6bcYDlE1FVVvDd6XZjF8utnla982yyRsQmX7CuC7Yw1vV31dfdgc
d+J9aFK4pCrCreJClcMl7B3F2AyY95jP/UtZinJ/JPaABBYr+xCkNpVycd0i0iZM9oXy3lniLUbU
xg/ljzcm79sTt5rtSb6BYLVdYYT75m16t3fGkjJkbSCnrd4N8NcVBhA0D7Ua5EcbiMJwJPqjxnq9
3pvwZkvngUHTkS9wYYsdlZvK7qnr7R2IfuMOOPZrqfzYs6wudACM0ZocYFXcQDV+ijZA3w1KH+Ps
8jSSroB+3KrZtXN0kMHH/Gu1xG/WeG1IIFYawOKChE5L16nwpkJUZOGK5cFmrpvITEfbp/O5MsSF
4RvDBPXCtYNm39aBXqLPi0p4wZmYhRkpD4/iB1p84B+w4T8LLBdizt6ERnZvsNTPyu431APGjon2
YJaf6FAjp59N4yYLrABeorq3wZqb02E4uALiruoaz0nE8JQm0iDki70yKnR2ZAM1K9Ocb+wDbYVd
xRjqk4oUccAddUfazpyOXYf711pXDY8M2lbaWo5SrKyxvbKs3gMNq3UqVB6rjeB0aKnER0/1e0Hb
o6AuegtJpkgSowfyHv+IuSxJNiaED36+yEO83nO0LsaqCnLYrB3PeNaydj9mXbFBfC75vScTItE1
AjmKRJ//phsZtkIwPIf7J2uB1e6Nm7sAZaefZkB3HzH/xYD121+9qzXmeBT2H+yy5I+sjveVSOST
b51tGhDPVcYWJX0Qx3xmBSxLj8c/nmb2nEjvmwQljfKNmOxYNorK7w6lUh/De5o/ZtQ/iv7/fLUc
BRIueMmDwDc1L4l83vkrMAwMo9KMlmkg65msH3Iqd7QRJwPq58mvUY1/WUnr4V5UPhHYUuR0lAk7
XBOy1N+RHGFo2xuRRUT1zAtmNG93bD85F5LF60lf/0gBBPJDlclwearwkLz0WV6NGdBMb9+RwKaw
RXOBvdR7Aa1ripXIshsaoX2aNTxWUw4ynv694ENqlivdGGmdusmc+1RM7fNnV7LxX1pvSo+i1hKY
mKTstGkKFAx3ENICMNG1yWabEIqC5IuSDO0vnirZUwyQWEj8HfgtaFgF5gqRWmeRYPq9l61FLrae
ksiA4rpkVtdmn9K51/V9NwIihyFc2rd2TrpvUImdiMqhuVodv1ZagcNh/6aGKv0fhoqLpfSA8+nA
E3lfLnJMK2sG/5TzcNuOOTKNUUP0n5UjIPGtxLtp3piX0ICNzFbvn7/07B/DQayRMP5bSCwD4Apj
iL6cc5fFADJHDdiN3yi+vvkb2ElXhlxCV8XNe6r2JLDNh58TXKzq7hWova5aztPOi6A21jhGdpXY
OgH9Pa1IlGIj7FmjZcU7g9QXq6EJw3AodB/jqCiOdFVQJYfCg5eu9Vvwv2zd7TA1oaQrlSIYGtLe
25IjxGGI78voz4fsLtgBD85jfOo8i34bQxBG+zSefKFRIqfiAfczGBzNSWxozfsSlL1tk3HQgiPg
fBHvMctT8YcKfIQEAjNJ7+iV+X0xTZGBSfMFiQ+Un+2QtfaAFoKnUSCOxH+t8aw3kvCheyJxnQ62
5MUE2kMqJEN8RwweWoRSi8rG/Nhwbnx7+niBUxTrypYw0b8gS/EZEM73FT6WlLrChPK3jYDzikK/
oJi3AnhDciFHNETTm7WGqvLaH8pSw2wnqdHjD+F7apsnspQRzcz90sYYHE5C4PyMGJOtIcMcwT/d
Ht1g73zXWA1xgzbcA2GFCUb3f2K2i6XC8rMkjYcXPlyIKeRfUE8N2mFdtRoizoYj3UFnmCwwi5SP
51rbxCqvgW2BDusaxgNV1xI6DWi9OxuJ4hjCABUSutz3Q4sw3xiFpaDA72ZFjZV0iqlhahA7dqEZ
ktw4OabyevMBbQShlI5jjI9UOT3DIv6q0OnQ/ACrE0dQ/mtfdY+AkpPaY+Ii1tRR2/rp4PVp1hAH
W6PmTegJ2B6mSoaScgtlHzm5Cbw/hV+1rbFK3tnwGGGijp15MrfwBcMYtm83AUNzBXIG8S+i37hq
5wb3k2S5/E6A3LluO3EbWEp/Mvf+10g2PI+eHqPe4zfQPcoy1RzXw0rVwgBXSGS713y9wKWPcFp+
F6gvIXyGo2EtpH2k593Xr4+y/NB4m7wB3IslMVvnUol9X7VMf4Rf6GssoAzZEjxrgCBipHx1cgTD
RF7uwe8g29ktQXgt3jVQhCMLvo9AKsAbHEyC3+m5LrXIZDW8W+LiBdUIX7JOHZKd89GRbCeQHV65
oD00A9FjsnccKniRTFxnqghgEUVP+Z84DGtFeOpqH3cYWnLGqJXglvvotz+GjbANiWUV2WMGwjNj
eZQbYciDesfcP9LOF98M2QGLm0eLLfyssyDQmC9cyuuQcOCbCQZufBe6Gmz2tY6qX33fUhrK2ihb
2z+JF1WVbfMGJRg32pO8Lgxrxl8utnsqM4bgT0HIW+6HhB0e0OpoBFYW43jzB9/RZnS0CB6x6ySu
veVk4jhpOY6D1FvnlRH7oI0FL3Ejq7iD8GTHWgkAekq7LzcoMDMG3p75xVYK7P45VSBiz1xAopGH
yGm1b1OVxWNvXZnxk3edFDXYS6Oi78eNRn01susYQnRNY11vEgTB+GwzpbSkdCx4xrAF3cyWwhiN
Qy7B4FVutp1eFiV4H5wiwduB0YkJzTwpZdoidcTU/FQ/bZpZ/6k5FrMWwMoklUdmVDyxF+YEn+uc
o+z5ZsHfL/dlqwuVPwzYNpta9DjDQRSkS3to1Bf8ono5UN0AcnkHR8DV8CrVuZEa3+KTHUiPMqVi
d/JNEtADgBDcns9fyPXxSA8a/XjpLMpT+FKyiSwlTgrOVQLO1iaFjX28diGAvVt1yrOFENp+7tWC
Bs1x7IlbCroelz+i33tBbBk/HdA/Ai5CBV5OYCxa5V4vAUF9EYcBggl9vbxK0THyQPm7u4jK4PSz
+Dj4U5URrvGGu/ETFcrL/4Vlgtt3N6HDa/N6wMS6ufxxBhKnVQxUhsS89PJ6hFcFhDyAYdmt6Iip
bljmCv1cJ5a4ckiKZALom9BBA0D3wVTBCfXpS50uFfa20kb1gmVa3gt1h/CGW/+clrzYSVztt0jn
tMRYp3sup04dUsMdaM1j/g9O029MtCDZUJsBs5IeWJOcy6amTDj6gmVlFzhbaXwoxWrFb7Hw5TUz
V9RBAvX3vj//iL3Yu7T6U0SuKHNv5Sl3a6ajkujki9OQ6ygfYKEMEaJbZqq7P6OnqbtSPqNaTAvH
zNiA8ar4XM4zPtp92qkARI1ZA8VyFZs/uFIuDkiT7El8Um1INsit72sfZWnVZFHiogWkJ22iN8OH
s3Jg6Ie6oFHoqf7HFxioRGIMHO2m37OUdnbYLRPNDyM5ufs+6W6WKRe9TTvllTG0JCWAMVuWZjDt
iOZWTx0h0Ctpm8aGuHgYRts0cvkMNp9quVlYW65CqK5MfPN8EwkuPU5IxvL2iKhy5RGJqGPn0Z5r
pEjwCzrdu/Ml2790Aiby+9YhifAHedRCJ9yMDJ0DdcEidkabTlSZhy4YlyxjLEOjNQ38MgvuaPGu
16gwTdshidMIl4aD4yQaWq2OJXgUwXExYvp0FO3ZUA4Gm8h756B3r3u7qGHdHJ0ay32tMjM5IXyo
fnnwSK2SSoHtV7sesLl53f2Ejb1Slp6kwE8Jz4VheUZrvOROtFJDVou1smR8yIwaLh2BSaqROtb8
QpTF9SI/rejw7DkwK5+kTLQfJsrRjmedboqWh4v09yTbHy53tz9PjLcp5fHJm0vWqgiIBPRevTd/
v5b6e14kkm9d3zPhTE+xcvdNWvmVEuzZEREvIBRV+Zhe0u6EON5GgTMz/HYywElmZdqOBUdK0BhS
odHUpORM3nuUi2RzA8KS/SOZEziK6t4/HqkgYpana1Td3kox50Rbc31pTy+b4oyUx+Ex3JDOEc1p
UsHMTZKH5vQTKncapjnJSd85/2gL6Ho6zqIIdiHB/HTXQOPQWwuuaqTjQ8Wv0RqvKA0l5oR18S8T
tF6f1iDNvcG0zmfapZwZqczs4Ar/eMyUJ8/5YFRL9ZxVBu0AZQ3R0KCAS4btN5+LG+uiVOYBhKwa
k/JKXGhMzdbDvI9t/Li9CjsG0+XJajXZWJVeT9HH2ggk5/j3dDY1sPPRicFoFh24lz3xHVJp/6uI
aLVeIGUI4jPoHld6z1DJxM7iDZJj7OOhSqOXRPP4Lhrfg5ps1Z8ud+MEmI7mChGYsfmc3ab8E1Xj
OB1gO1cGcv0IBqQ1DkZNPLIfAxcEQd1cqSWUYtWXGLficmAg48hzAjHetBK2AK3LId/zwF0oqxgh
HOkEsOBxP6I1WHu8nUKf/KmPUmQJdiDdLWWF+JTSDX8HpvqzvQvA2scdtyDAB8bIuORKGhYVqq2o
kMXyBzciUgMFnDwT2snMf4MeMsy/8LsK+wo/GfICZsg6eoTvi8hZPzro2a+TykV0TTue2ceuh8Rg
q0qkovJvld9PYCtO8kx1NFSMBxlukFKwThoBiw96heKg4CTmkI277RQpjVx0pycB3US9Ni60SNBI
yLEB+8lR167A+5bRjq5aXiEteyUQD1HvtSNpUseqxLgk7sPldEaT21Se3r7R5Ud4XlJxRRP7NhWP
Vs2ayWCnLgi+DoP0JIJn9KQZLG0EfqL6OzCvoUIaQA8kDyQ5u8k5+ooCuIVw/2604y/yEoKzs7jZ
4LgJG2+ysY/a7HAXHbPUE7W0iJdlqrQ4vdIuBqH3BDWJ3kg2Tl7Ei5OvpRqXIMKHCSH3+IQu/hJk
rI7SMlpPgfbnilGGRAtObCxJ3/syAuTff6cPe2sVVDZOWQBKyp87xSSdtLjIBB1tYyMlwj7OCQ1s
Y/AFH4OzGYZCpy/grum62sHAakhEaUMndPG93QrPCumG6xeix3qpRWMMfEz2lNNFXp6v6H/Oi9dQ
wasvpCBFj0kWiDoiLvmziHkvM7DoOGcLzuMJru1H0v/tcAJI5CHlvuDQ94yceJX83mcvuHbzUv/b
5KMuTvjtvbJQgZrt1C858kLxcqG4bB+zr7hSXtj5jNlBiPtiFz/GbNQafRufNKk6DlMwj+mbMiqD
gC7X0w7kaXRbhvz5agiBx61e+5Bu7nRsNkLnsGGfM04RPyf/gfrlKjET3gOP2Mb/RNy7dQPV5ttG
XTUXadYnp2NamImFl/3OgepCurEp5Yyl4rEiDya2tIC8S++arO062RYeaGOPdaQB74S/ElfFuAL+
Va9+F5y5AXcCdeQUrqzv6d7AuYI7PnpM+hkzJWmlYn0IH3/H3MaRzw2y/t0V3sJfWDr/B5/wVX53
Xs3xZPEVmnw3KlS49ZYl/9wMn8rBAnhYAjRX7uI/E7dDh2rGekfkez5Z0dbM+V4cET4jcyWUVumC
kJNqUCrcq7QsuwkIkQJ2jd9KsHBjgD2m3btRFeTQdeAMCaBLmfclojx3GwJpUsJvR5eG7LVFlc7i
/yuMXSN57DPGTA8lr/YTcs7uQG/xGokZQPhP1M1Pv5QD353M2Q5mkBWic4BCcxR6qnlX1rd60syp
hsigW35oRgm1xt0VzZJt27FLRVPshioMGYMAuhlI9N7RWnn6qsdj/sWDbOihKRTvNhKDKJ6XQviP
Y6NtM3yf4T1X0DnTUmAvSplYRNlndLDYDeR+fJvHBGR5lZCmKczBJmxXpl3neCGuyFv3zBbVkMv3
5TDbhm54Qc+r2JvHLY4JNliD2p2b+Xo3t89xnlZd7hjSjmMtT7saM5Co5gEVU8XEPIW6Ta9ZmjIk
0BQIfhRRrI0o7MZdeja2Da3PUWKa186+PEWBf1KLKFVUgTQjn+blX9IhpjXLKUGvHxaXpAevI3fF
MlYpUj/ZNwXJOFT5vi/fopqsVqqF/iyRKRopnT619dkKaWQBIURfp+e8BiZrGzh7IrY5xQAtYfly
dqxqQW8fOEMPqUB4HFl1gsud64BzPf+Fi1MJuEOiQ5tSIx0cQJ3GlFWLOQhJaeaL/s14IkpGocuw
VIZGPTICNiF3In+C9I9O7ggULEVSWkl5rXrqemIartMmuSaUN8AaYUWMGemE+3KJXbQSefaWvB1D
IEoH6XsEey5YKTp53X/dAGsHK+XG3QQiFejoF0gt19F5dIdgLFemqepKifzQQXr4SYoFrP5tI/aU
R7DDi5XN4xaYI1tSG06ZJjcHmANLsAZksaL4WpWthPDBaTr24AAV8oxeLtVaPpI3ZmjupUQAeWaD
5UPZqMVVDm7HXrwUfDTzPJFW6oplb1Dufqp4UzBvnt2TpS6CDBpWuM4JwajSzQDaUg0pvp/m45Yj
uZNS1guW4eDxKWfa9nDH4Yr7YTsmtA8ZONDg1Kbjky+Nh9+Z7CqGrdgbv1bMaMbc3g5FaagMadeU
kcmEmHDz3D30pbnB+8AOYHQsLdzS8br4rE/5StDatNh7+9TOQPNhMtfPcJLpTNBK+7PvIwA0IRM2
jRRHrGDP39Bvmf7oiIh/+ezZWetWhL2lg7Yo/kzwHg3/WRSVuTg5glW6vgP2pNQ15JJD7H2xUVed
VQHP5AbjHmMvsKvFBAx9mCea78582O+7Xeq1yI52OqTkjG1b1FxAweTXrfQfrAvS+MoNwBRko92N
Va1jlbKJj1fcV9/ZVMVHEeW/brniwyqEU7+63RfUbDOli0Ptye+89E3dA8Cys+u94jPhtkrVeTOF
BjVEytK2NesK+Og6KlJx7hKoOwxqSQNq0xrPLDRmtx/v+JDZgSm4X4D2EBOUit3eJP1ilsWpZl7h
ufrRSztmr47DwYghwz7FgTAFiYxSVRhYnxLfNdB3UDjY6DM/0RWZHNvUltNvNVajmNoFNpRP3Gsi
SXwTje4Oq/sIdY+j95DTJfzjFLeyYI1NuQLvY9yaRyLAPY1uYKXOnS8nRQFhIOb/KVyJber739cw
e07u5yyz6AYrR0kp9PNisHbcNkqBO4awXqmMjP4tUMWAC/LkHZJ3DTmz8Dym4jC529ATWIFTc3rX
hICovN8ykZ64Gervxb77ne5uID5thDBIMd5/TiWw08DKONhaFVsGcTkYr1b8vHXfrqVALKgWPmjL
bYXt7s7N0DniMiRa+0KN66Qa9JUk2R8E3C3nLWyCVA9V+6iLWrAp7nSDb6xZN2PyAmcJ63ZsRi7+
5VEjqIEgKfFXYHR7SklPdHDRkoifnoFHzxh+dxUqydzeN1DwYdydZie96h9EB8wEeSb0x05RDGF+
RNR7LCJB8qEI8+9RZg3KTKMngMDxgj9+IILKeWmro64o0jo+lBs9LM+8hER60GIq6kgp702PNsDM
jf3KM2og2V1tem8TY2AU91RNmo3Fle647JS0jxobL1mQoUkISt1M+1VeQBFLcl7d4k0Ava/wKK/Q
KnFzBPaKRZ4hG583RCLI7HL60K9bcbIYeF9l482igqn4Li74XfUc71XvhANBvRzfSTWwkKTMqzph
9Y1lPtx3e8N/xXJ619nXdFnxZMhL1Cc3sHzEZqfvDTFgrQKVkyErjfZO0ODEFyTvSdC/FxsbIG8U
Rz3/HI7xr7r067wYucnfQ4ThwMFYKBKkiK/U8JnS08HSk/NyKT8s74e2zscy7KB3JH6WeyX3nqXj
a1dFU8tCJhceXr7k/iYCBuz+nFL44aM1p1sq9n2zZaGgOSR71y4UhxHLK54TAA8MvBCpDdkGGKAW
5QnUjb6/RFlbup6xmARxzcRM63K4vF5lMUHgIl/Xxf1dndjO61zl/VCLE0HaiMFmfsdQqTYEhXPn
nqv1BHo1T6JSbAMbCddWfEGOAWCPxRMnA2rfaX6byZyVPehICzBYQfgA2pwBCsZY9Ort1o8TPw0Z
2rgahnPq0aBJKMuWUUqdcZaioNVD0fszt5nu+SAa888A391+UA3rbmph78t3RG333RMwVkj0k3XQ
P01QhDY+l4jCQ5iKGJ01NUSjkFT1Gh5v/Ng7USxtDB9zQ/E7Fvpo+8/3nUCxWOcHW3lQnYGoovQB
Da22EVuAQGBPg0NcmFIV0Q7BoP0vKf9p+RakRnayvDXFLtdnGdZmVrYPju4QONnutGdIj9KOmDC5
WK9FHgj81pMJ6BiY4tWNcDPpzYpBWAjHqboZoOe+xry+4msbXA4DIJQdyTl2PzU0yPrUxIkrC3PD
vNZDVxpCcr0tUZ59GGZWLi0WnGh+GlXDtQJWflZbuaw1lCQFtIEgHNcSj/6Pnfxg7oVT0YgC4oqQ
um9avaqzapTcQ0D8IGNh9daahqxQE3x3emZAv3pdaEt0zfdwMCYZ+CFAtFyrVUJXmwvdYHHoh1I9
+COlv92x3OW69PqkTtA5ZadMB0R7/vljtJCnfkHWee9a5tAHr4sGXRicyzBUzelh/nh4k5cuHa7N
fMAh3I4XHpY8/mAxGECUiZHLih1DqBKgxQx/1f3+XnoFug95maiIBIo19g8DnCyz0P38AKz31nZy
2UueN41Boo19FKluCSqfSagkorrwexo3+C2n5z5WPAJmgV7UZaq+HhSRz0HFIkkLkLMm6HJ80pUI
ERRf8eFiX18up82lOB0rzGZBBsSAgoa3CMazVbuwZSEOGx2YQQ0UDdPHoYAOo9lS8MvvUl/6WJFq
BVPLcn+d9GuJIwSDHJ8uwpfo3CJao4anlVM9SIsDrZWtSGa6lUFTawN/bxl6k6pALf74odPj2w+P
hQWftl+SAswvl5Q+fMy6+RQJkrTGeDuFskcwlQXYRtcsnXo8mHgaYPiNrj5dZwpFPzZBdZuoXc44
Nc3+jgXoDFFGU3IsKthkVXv69j5Yh7F+oxL5P90T6039cBoZfoL6/PIB74Elh51k0QuXMOeC/jpn
gVpZIr4VxBk8l807u09XiZEMVKTrbBqZcCCjLvYYD/eOgM1gDp8SyDfeALHMqFWPbmWSke4FxWdd
i1ZXeWnXrdq/xC0jYEnJmM4isdsTx6OU+HIZtDv3q3Rxaf9P44zQxcGmnxDd2uCrSMNv5HXPSzo6
fJGjh6/pjIyA0+0zDRaYYY1PMTfEuW5vtoXGBpOl/LJykgh/7TymLkuT7zGYq70SOvQNaTzEg48k
B1h+uPnj8JmC//jmYmQdEGt4KSv7VzCefk4RI45BOixmSJi42visJok3f53tBvikq6QDTez7d+hs
eTGNU5sQ7DK+rOscQkKIwYoOU2j8knGJBBzNQBNMPCmUub3ldRJ9iMDQtssxxL9p7Y3M4zEYUcxS
ZrKYoKpczhh4Tk2RI0rW7BOTktm3YwQy8vt+cYHVUUX4Y+x9VCbNRwJ/SAkHbn8dtpM2gROL6s6t
g9UBcTVS45vrNYFwJUnXNqGKCVpXmZJgIs03SdApm6kJNx1eE/rsDcfYeNH/dkT1+AGjeWKEJgbs
ViD1EdjGOchUNc8L3tUgOeabXNEmmaXe+9Zl8ANYwtb9A5lR6FvaiVhkOSR6V9Gr7EVSVzFhwfPR
xv9WXW9TXxLrJtMliJHQ7Qy8N/CScanpkXeEXEohbCgcjhBvXM9x3VZR4dY30Ugm7nxaO2VWRCFu
f5WLYJs+rHaM90L0VOwFdX3KW4ZVjepygKZBM1ah8IHQr9N86AZB5m8ccXfhP01DshrkHoY6Q4dl
XUCjZoIHVbQu6m8Z8WTXK94IUL+aNezPUEWHrW0kHZgCZJwJCYszTa45iCSzGufUmsm12N8vAau1
izQdS3dPCsBCCyg5cud/CIHtDnhfgD5vj95oSr/kpzRQMbu5iZgkqcOyx/4I4MVghGcjyk1W3qtR
EOGANSHSxGzIjuXBWeokbPPpUGBT4CZxqvMEpsmk15SFqZ/v4cYrka5htgpv+dtwYcXDIVrYY/BT
MLG5FfvTg+9cKYQ8kO554VLgzdWKTTt3hsQ17lTfjxzkCZZ1aINgHczn7FNxlT2LbZdaZg+O8C6j
nX9q7QSTyCtEqRsaQVJBya8uge5IwgePY+OtkdkNKNYXWUBgQXbqzu/p9od6l37MDFs88MqGB5+i
qAwi/Yf4/8tsvo2WTqcsUNPsHteEhDAtELO8JdRft+IMxy0bJulWZihxBO65Ep0uXFSI5a7a5vs9
2Jm+ONCDUf48ozylEoVt8fJoOzpm4zNXBuNQQ4qyHbK1wP/3e5+QK0AR6aI9PTyVkYw3833livNN
K9tg0muDUTEGo6QPFLkVNO8NV3RdEFDPbCimdBhPiv/rsG1nh2y+2Mf4W0j/3j6nadIwwQjwz4Rk
0uuDy4zJFQJ3NZHyCbT+GPWsgFUAO5s0Kw+s5+OYIoi9/RztfvV3Pvi+xsj69KPpAU6KAVk7RK0G
7bTLg3qRJXmRtzzrapUrP3A1ZTnFpwjpTdRIRR+rHDyDI2RIgy3C0Xu63eq10AWO6cNeYZv57Q1s
otqGvZE5WN3W0AgYqalSHSuiMatpIzH9+ZZagCLyRZFzSaxa/stuGs46rnxbfWbY0WwMQghzBnYy
WjTxQIVHi9KGD/sqDwT2vMMZUmaUILh3ysLVD+x9CMYcmLlrTqBr4tjApzQR2TJywRgXnb1O4iyC
smXKK8Z5WgHNkPDR6+u8H7cE7Sq4tjelyMz1UmmLB5NB3SKoDQ/sWRGFYLOkceFteBQC0ST6FqoW
/NQ3GTKH2oGbFk5IJTG0+Hu4qwwHLpC+B3sQJINua4Y7/oFJ2JoE5Wcm4fz+Ria6MoTARF/RTl65
1g7wvDz+AfDwuIdpWLpvUHigcxa8sdduGXa2Ys0WH6HW045CDv6YqfsaShU6jeOfc7EcT+QXEqmA
8AWFl6FjK7+gAWRFEEohz30Io27LQ4nlMBMng5zW2EmfI9HypjqNjNV/pbLr+fU6eAPLLQyztwUo
t0OMyjBcwXi3TobYS1YV4PbQGI1fCNHnUjg769fNuiVajkuIA5OxT6RGlfeLR4HWdGV3PGuhIjpv
yKssc3njNg4yFdwzpzlFKZi4Ql1UrZFxq8eM8dJea2czwP+XFqLofCesquUFAGXF1SYmoYzajeS5
rPiipvCHAa0HMJ3j1lM53F1ZvXGTb/QBuGphfPWiJbosP4INMcKubYUOPYCEarY0E5Q+3NN60K7b
a9XRZ7ez/iLL8U8tUcsuns0VQEOITt9ZGaUj9THW7Lg8Zb7nNlFXnly8jnkTBMGcIHWYb3O3r3PU
CMYGZinZW7vBnfOx9NQvYR3rb4EiiTRtAhIx4erPBz6ZsPdyVC2lsvL/tL4ERcpdYku8BEAEHwmg
KUwQBA9bEJ3jjvu73tPl9ArSztzMTUcUno2TAW7ZRsLPZs4nZZ0b8kVOvtuxY+aHgih9P4AxvDLi
o3mhfW8w3RbpVYg4o9Ivo93Yo+gr/FdCIQ/cWwi5FN0KAzv31zK662ednzqkhkkn5wWQt55l62sz
YOaJ9WlLDO2eXynleTFY7BlSa5Og4Tj3Ii8yd5enJC8aVfXrHL9K+BvENwfuU+8qulanWBehm0SA
/4hblLtoNroc9zOL2iUvh3+DFC6C9egn0xJBUQsvUSNR15I0xsVJxMXs9jYbEkFs1fEEgpgiunlR
J3+yMYT9ukYdjNpmyB3SSjtO7uAWFGyddWJsfLZF0pkVr4yddp8ArYlcncPy4snrGI5/54iwV0a3
2bnwSFBtl5DcquGDLOOgcQ8SPLZNM+TrDK89v21Bcvmkr4Nl7XMCy3LkxYsj7H1UNx2HBPusOOqx
L1cYGMwF2ejdgxfZlGwC3FobUadalZzRllE9hYE24dofOoDQAzQEcKPjXYdDEHTPdeEBwogA8159
iGYifVx1jNkxHVHNmWhyv6/MM/y0dG1oA+s6pVVec8YQrHOV5H5Bh6wqA6k4JH7kfcgP4C7IbKqn
cv+N7MuYmRrz0Z7Y6fT820Y//M6PogqnjwNz1fFQ95Q1q87/Fnl7Uy2jDMQYuema9vTMD2ayZ/Y3
TMWW85DBejhCu0WW+EDqW36BQY9H99YtGl4EOZ+93k1i2LtNoJLC3w6ZGBjuYiGXC6ys5CqhZQNO
vH3JvMzpsIZ7i7Z6JQDFg5/7Uuk76hLZ5kvnEOWl7ZDJqcqdGHIJzQRhtJvM+KH0e6W4rYhGtWjB
C+QyHsboX7GqsTly54Byl9MWTzmG3SyB0Xl+bCVKM46p2hs2JYhSfId0vfpqZvLae/R8+qwZrR9o
wpPp2u+ne6p27t1IH3xKYCSOxGyK7ga1h7ct1f0Vj7Ys0n4eUKSEBYvOuHvuPpIox+UlOZqGCXD8
NGmwX13SmmARA4t2mzhZ0HXp4aAyhDgk0rYOpOEi7HN5+Gk48GMkOmh0fTIFPh1D+oSGHbEVyWQv
srLV/aciVx7KF6hDn/UDxMgyO3JPI4qQ2zBchxT9d7QEQw2/nR8Z5e2n0CrIKAFNj/hX97AVhE8q
fZSJG0VqdJ+4hzceATV04TZ1MrHSNAIjm+d7Sk+3/lWRAAFs0BBAGC+7RsaUZ2uBtKhLKvA/KdKF
fROkwGcsQnPtbpOdoIQqFb0bypr+DVGPToWryIoOkSDOLwv68TaRrYPQgIe1WbUoTfD/EBKkSU9h
IrIgRnxV4ZOjwueYHvrHcrN2dsBq1XL5F97ApsQ/OpB8WVCGqIyTVlOVGw0AZSBsxKNraqyafgR8
owOOl1AdKSHh+rd2OY7aYJr8+bfQ5NJDBEO9C+KFNFEqssL1tKt+DzcQ+aWK+vy9UycCWWkGbMLc
EyJ+k05+uU9eaaEMHNhp3PVmM2zcLElInAlifOah2S+oib7FcQV8DgQ1CaoVhlvnWB6ahtNtpuE6
Qim5fD0TW1fUviyvwA1GuR2FZEqeUZjmyuXtJ1g2z0f1Q66FpJlbHckzFeHdufs3lr3UXZoWR6FW
00L+p5KBrHJx33jzBzyNPV9dG/LASGKltfLDu6Q1NuCxAYv8wxPItG8wvSmGnlqqAajQE6PdbjIq
Vvk+m4O5zdBhzmFy2ncwrUireqEK91xeLN0Z+jnvg/V857oAT9FvS54KB1voNCFg/3cvdW448iJ1
rDzvP7Ps0gyGLKVYXjKa+yiW5RKCP6AGsJqWwJwIrr/g8vmuBQdc+naMzA2SIN8sa9Ujy11bMVNL
Gjz9StVZSaB4OX4v+Tf2MJnUnVCvIFHtIwxCHFTOEUPGySUCScpoluLR1KcrRKK6bsvBxydfWEs4
oTA9TvDARVHsRIUyvxipJQ07udOWrAX/2vMu8eSo5yPA2fn1d5sx5P1MobSNk+HuRhMgghj/pVbq
wJRIa+FV2/U7qZGZyA7+cJuVik0K6HwgpCCS01kEUEjETJzGUPvU1fAwIcQF39cjPMTPveIec+8X
XAqN0XGzeOAJM3pjH9tJThs4OonryrZgeYtZuFC9ME2+cFPdXcFkLVfyehnwDp/2D8FqwRFH5EPB
/LTkilaKuFnXOTzEMV5rMeZLpZdE/rYj0Ll5Hdtk7oLYnS0GADj6TU7zUVrL5P1K7bDQiDjHRiyg
0MRevkbgVvWifwK+SaVMiOHdcR77D5Ct1v5IpU76jqwPLxI8srcFQKTOJgEJd5DvmAR+OWA8aaQr
i+XMN83ZrE3FwuysvPg5qKFaXjDBchF3REg6xs3kCMDm6GgCDJIioS0RnBfZLJHLQWGUiovnx0gw
O0/BYV+x2mj1RDUFnBz8Qrm6Z+V2QCR/bT+7jfIMMOevuLoZK8NyyQ3AA9eLIemqSJdSqc3Zm9WF
1NAyZpMISiilrQ14B8N2PwdYvQGycyq5J6jf9n3IA2B/W4MfLoMq0ILCeu8DJ/1u5mqA2Fxdq8/K
HJCwm1ED+VcIoMMfumYSnESHYmtv+R1/apjtaVbQWJqYLfCUayNRey5kqcV+V70YHTU1HoRd4Uir
HKqMJHyYGIArZYE9+Oib3NaN0tqWxuJdh4PGg9nt0O1tx8B9et0lKYV7WRie3aY4reyIJiuErXHf
1RJls855dtVRKKxxagw9WOD3k1O901vta8BIHoKCEzr1yRwJ7QilI3243a0+YhjajygogA6FLYME
eKbSKgAbxIgkdWwEKDl71MwD9OB91hrbiPZQeZX90c+0rppMpFmhXnfexzr5Zk9V9UfCcG6V4fqZ
S5TGKPdlmHf/i4XLQlwP7PC/Jk1PMJDcKf/KsFB5jBhDIRdyq0WK2efz5RsWHNXug63cDFvsYwMa
NAMXz4HDfbhRpIiMlKqbrGFWNfZPwEKoxigGA4BhQA0AJfRrnEO1NKDSJG22TSxzjaxTfZbAbmxu
xS/ttnSNCugpFdmwAdtHYv9iBjWdgp3O8327s/IgJKnmr1Yb72lwfkqcaHQ/fkDPbxccpMt4Tkri
9sSU6MIAkwbOdGKnjPBiUHwxc/f6ByqkcaEh3XFYCQ5bIYuQo2yFK50rYG2iVj017wVaFwr9xFT+
Iv589d2UFp+RktVsQqvQRkiqzKTw3jUpf/F+0n2QnoyTd3nQqryi9fCxEYLoIa6hAaEc5NuvOQlk
TPjXQXw4ujeviSuMqgX18SC1DT37wzwvDeWUeVQZChFM0mtUdso9a3OsrofuYVXwN61GbSUpeOLm
cv08KXuciPwYauYsmJCXZyFeE9H2LgEKxmgUVJEBmTNmSeBZQDlK8Yyw6fRO92+03twG6IibsW3a
XLmraa95beEbf90yTL3nmuBgZ4dEnUKyvtMASXyl7qQyOhi5lR7qq5u3fiqSyArYwnNb8Ro9JlS8
8gXy0ZJG2ssO4NQm8LssEJXQdGDP1DYtZRQxAIeQottX3QOMWDuHWIOvXzMWy3b+gl/lrW0B0yPN
/rHXC7/UACr+kDtYDNMUftFbdsG4c9W9YJJ2ox09IoPYF5xHmZ89i1hnnbPNrlypvnuRbFf67TeV
hk9zajEtvt/HeIL7l88cSSWc0Hk4FZymwVfkNdsuAqrTaQkQZKcI2KHcNuFFsQH8YtEEWIgPeftc
Bac2Bea5ElLxZwG9u+LQs1ud+P6oBYwLMPDXecbeJl6vWXCewcBuLcV0rAlKQ59omJGWMgeAcs36
en5FFd6Z6rCzyc275Eotd/VoXyomKF+ZUDdMAeuunQtXPMqDDLMTZc3PnJw+cVBtuXTBqR3+Gpqk
1JqKQf0e/0a7K8xvWQSI1efDf1Y0Iv4vohi8AEFt0d0KametVgpnFEFn+Wz9WYZZzirWwPuM8Fzi
vMNyo/ljrPuYdDI+Z3Dn0lipLvICTDfE2MJ67eDyY2igu3pzkAiTUM4qQxev9g6X9QahSr8jNDUQ
2ctTWpIxPfougy6k29sDiZPqOQwy2t+Q1/5e/fjFn/UhbTLBorbPap0OGUDw9zjY/7A6EvTdL5H/
uJuxhrQ3jeS6RThWwFP91OER96k31Rppgvma18gNU/fWeKzA2vibXGd5YQF5732sw5PsacC8YNkk
LVdZnkIWWTnaPCimWwYSw/WC1N7qFQpaBBs3fZZkIRtPeG4tKwJimQDVlGP2DyFZ5Xnrjc5Hl09O
FjujCEQlTounpvsaW9nwoCOEntFECkSqfndmvZ1GuxhpGpAV65M+YrTs046IdCmMTPVXz0eGEJev
zlivd/9/LAmaTKfWlnzG8eYStMzx2kqE6382n3J6xoKLmgfefLzt2AMn1g6Sb/tr2s/M15zdrZOC
ZZ94SCVtYx7NMqxUXDx7NV9gLfDKH6Ceb8a2f6+NHfUHLwvtOuGotTC41r9CJY6poka/qJMIrqiz
bvdFPe2RWtdJKTVDjJi0vQz3zDIG5BAx1/1n4Ev2LKrvdAnuhIESfTP1kSWrnkxBrF1BZ+3e8wAO
Y2XqdU9srZFsICvcX3cXNq5EuvjmXbac5QxWwYBP4W9cB77yDk24+sNpNsr8TWmcWk9A8mvFy0nJ
8PhKkDYRFUoO9Ggie7U6Nu8y7La6JOYo3JOZdDsiuHSyqFMKF/bXF5McNYS/71SyITNuLEk8FU3w
axBPY42WmYjoN4/1WtR2nPNHlRwQFzlz6aXni3SmmwRPxA72RhwffXpqpvNe+0gYXuNmhSMYtzV2
sx1t2kbXPnznu7ubXAkVW9k+lTY3rAdwtK7bqq38A3hBcmQX8yq9xAIO8ub1tWFFERO5EF5d/VDA
/DJLjeit3ICDXe/dloiXYm4Amfe1pTJURc82CxO7O5mMb5yAYRhHKdC3CNust+Ez8cyXWelXJnK8
H1saiSlgYQM0t6hFpwH3Xu8Xu1uDk2SthnfLjUZUWtcYmZVDfYTkvib1ThyytIGGxodmbgA951bf
elxjGZO8rmR0dOZA7mqqxUdPD7N5QZRyZ3MN5K1GUBZcE8kN9jM6446siOobap6LH+9zif+tubxQ
NfW/krc01M2tGYEDQmycxzhlGTZLFXj25U1cd/pgONW+XzXe5XvodElbmNi6rNqRs1l4YsrHU32b
U/+UHEMsfm3MBXnzWTwF/u8c5EdX0JPcEwQfuuq6ULGXA3KQr5Ar1noVn/1aZYwQ7WUnEZ4WSpB3
wCvfxUDfQN1/bCDpZ9p/K9wwS4dAKtLCuvj74IA3mLGVfM5yDnfaaD2UJCnqd52Kc6P5pxPw6Gqq
UhGtoW1pIOYwLUlIXO/1Ci5lDpoJ8vDKDykpam28s+mYpCnOf1p2iVwVclL72f0+o1XGcMIcP9So
9R6MeuCv31h84BEmqgUC/MQYX4+eFPbkCmVEwVIXbifkjx7H1E25UhGe5KdhaJaUHTPJyqMZ6qXw
i6XzqwcJbH3qge/Y/oucymqMnYBn/+FnCz8NgVpyJIMdXWQd93HJsm4KExB6Xp3RMjLVIgXdi1Ue
e9X11nT+94pyvnyO2oHtgFZF/NSRV+jJE1S0MdVeCMmwBjSfjVopUFVIfo4Ec8CvGFILQAistvc6
HIN9pEhdNZ6trypcfXDRBwiNbfZPR0XJj9niovgaJfdxCUAO+M1PbWGgM6F6jM4itTZulqCzb76g
J/7ld0fUP0Z2t/utepcRrfN+ZIKHa7T4TF88myGeKZhl6RbNtaVv73mVnlTGnwPaHyZlFHMsndzl
h9BNgGFv+snelq9V6hhlcuHaTdKmkqG6Xa3Oo7h4mWGNSZoX4QmOC6OHKpzEIhgpc13i5MKlvY3H
oG4wI8z8yamwl2hmTFmP5wu00EvKpytis2GaisFjAKxWJyIUmZqTvof6JunwZVSUzDdyvDjKfLi/
OLs+d/vqdiRGOy1VblY40E6WVn7DrREYtci/HqGq4r0TawNX+G73EXoBZwhnOru3g2txWY6QjHNg
A/Jh4wria01TC9sPGSBYTBBPRuRZctFERPS1FjoI2WfgQrbldJ1rpdOQVkEATULp3LcCPA5WXSj4
XDa07zFdrOsp8H3c/5Y01/jhjXyJFWbmAIW1V6+2ltrLFlfv9+PmpL8V/RiccwTVYj7dwOXGYIRB
X0Qvk4Ow/JGaxiMrq0FZkqjc70A6bAqm+w6oWq0d7a/kassp2tD0GD1aF31h3dmVGZR0TnaCpIol
sc0yt8yUXSgw97pkIp3mBzStWkSLrAESV+cU2y4f9WazLpNlNmPBdH3K2P8csjLN375itTWeKv/P
1ZPr6R17LY4Ju2JGTnJ8qhxb+BlahhB2gYW/AW3abUWpww5ti3ru8ggzvPfgctNAoSQrRcO+mr1w
WxpBgILiNjdlynvY7SukZSa+PjE+/j3Z/AmJ8XlIRCuJAnphmxt08bhFFQzA4pmXmzqU9hROVLRN
8303eSg743b+PxPHUNq6zlaE9HzVVk1URlkAPPOqrIeOGhlHTQgXX45Sgg/+KM13NBbiogoMOnuM
+23gOhaNtA5P4eEWZHDgGAAUVKuIssduoggQ/yRi4QtpvcHpmoEeXIACOjk1sZ0Kor16HiCe4j2p
2Uq5D7wdX5MZezZ6I3HpM1Zyq/5005uL5KTUWxGWVJuChZMV05YsfSXh9eI0AxHBYc5BuisM6+3w
TpHLY7IXZ40AGsDi3PBcmBaunXBRFYyQIIxYi9GGbz45wgEc4UyUsWNrwUGc4TubpklDSNs8vjqT
P3sqGMeRTVQhrFC4WfSxFmy614aUdy70EJ21qRFaK3YvSfepxy7KtZzhFnNRgAWkRMG2uC51i4gD
dQvtU7h1+4W1JOWhlHITDjVMg5K0+QoeNvhQ3FTIqVDVv/ke2Fz20UfreiLvhIsc8fzxYfEB/UB1
iTFQlz2UUr38D7Xx4hcrdegNNkB19aUxREuj3Z8DsezZPJL637/2GcKzfnGyVwGlyAmM5xwZd7Kb
II8m/yr6rWZjt777zqnDfybSNxteCUtMdcq3oMI617Y2O6rk1T3Hy4Awgq2/ctIBhMc2TLCCIXHG
XO3uqDWXYgr2U/cK4ZnA6HOaidv7pD2Iymc49AAMajP21PGKGXfQPZgScx1qjuimoVrmgCoz7MGe
lpG8+crJr6HGkPGszkwJ24v/+rPw1AsrbIntByO24VpI06ysYq1pL+P29NHXmrhQhAJmM8kuGWGL
HGCIUWuAdChrsFCywtyrAIeJeUN0rMUCUg+E/s6BTHnc0aYbGYc9wZNIP62rBjiIEhIvC+2PkTJ0
naWKeXGB4dpz7UqzMLzyAvvOsi3HJ+1ANyHHxLS4goiLg5gOt32IKCQ8YlD84NRQa8XYp3xVUpnX
ZTDve07/UIytGsiS5xjBh++kw2cKjvtG2jBA6oBa2PU7yxcCKvtGOtJSViAtsCjNTwI08s3PUNb/
urSb9x5lffVpAWUr0qsipGKWfdIyOJGfA23t+lJOuXMiyvTZ/chN/HWZzx+WZ3CHJWk2t9L+vcEV
i0jeB79qvcuQ6frIYIqEksG6B8wSI8INmY3newNvugqcfQkV9ynTU4lF9i74PfCXI3Iot5QBtJpD
mYCPpr61iDhVOag5R+NxjMh6dcAdvAEHafPyvHWRRutShtURsPmr351SEQ2/jGknOQGAUeaIPMeR
kgaZoEP6TCU6v7JYKON1VCR1Be06eDF+RDN60JKLDJX57Zokiq/RqFvjkTWfg03ifqlLFSPLyLw1
3oel7HE7UP/MbYZs7OUVgu/krCuEnaBJdV7BUXrJgsTi885atmTNrR5UoHtJRpfhTwrDQSyCdmkG
texYgO8J3/6PYIpaxltmi6dW0rNc5oqnfdhj1URWrwJN9ld9NZMUpfeSFm2oWlYIHccggbi79H3Z
FOYdQDQz+mKiBjBQDnkEJTNIbUVz1uHWTI+mDp6Z6Rcx8Ya0iZDJ+2fUU3B+hi5vqC2yrpEguicT
IYHUidcgIC+jCZDmAwhmVpUdCs4zuZ41CU1bH6WnAB+jOVTkqIjT8Y/O8wDkXPIFrWczBZsu39P1
JjRF+E50+Im53OFbnv5f88f0G/Y5lsXpmlPQKAZVlMP+1P5llCGNTHFqsEbU9NyY7TMFwCAQ6t/S
djAl3uRF7SEe1LWtSgx3WdzBpek6r1VmIhmsedkJTZyLfre1Sn996J4hTPuP28oW5iv5It7DRua5
JFvG7tDIRFh0TFm5AIbaFJrkAsrz+964LaR4bu6Wypcfb0eoLVLLZXA9CjAAwEyckaqXVFu64l9r
Iw9Q0SsRGQQ3honIOujSp+6jM35FMFrPvxsjLMsRzgycYbI/+kvcw8gj9SMdi20rbzHMg3m5m2LR
HgICKSdnQXt5Uj3ZNEfu7dP/JET9W2P/KnXfvCnlVAot149ju7JNZvPlVdheDjZktFICdTV+aH0V
6rHmz1Qd2xdgI5I4o8tnHCAEeJf6RNnQKB/loDKyBZB2Ys6n1QC6i7n8AOOF/8nnKTgDs7yjcVd4
m9sKdXlHkXThB5QajSzb/rbb4cIdIRxL+gxJNsCKpoj6v0KCbEDB6NnJJvpQqOnmg2xzywGtL7sa
tcLz6733E+Fb36+jsxG5IG2KcgFu6tJesrl56d62VIeYpTXM43tb8fn8irx2Y1BmUCFky+HnfPGM
UpuXNpyEA5D65cyb/YmHyy1qB38ADzIdh29Mzp2wjVVYmILualGqc3MKsTM5YSQKIuWEO26fEhI5
PleBfh/gxEXGj4kXVHKj9y85/M0gOk9C9GHdgPTH8ZlkhWrfwRZinnBPRcwwMZMSRq+wiod0KZZ2
uImrP9seb/HWf4CiDy24t0gi9sDdEbVC/JFcE4SAcRA+E6N87PYkrPLZFaUngc55oL7dPp9j5/L1
0z7tjrbCqUYThoF9UqESi3iO+9Ss+eK754nF+3wGGjXQB6aQwjO30iHsKCIcQ8/59GcF4q5UTtn/
TmC7Z13oNISD8XZL26iSgFRsMN4R/TgyCCAxaahD47uV7ZMI3UiMsv3frdTQknGFxNyCsKB225cf
zWZUt6uFLVkGzMNpJ0CPWH8cVHCNpRuTYmxgEeob0RJNikPqEfPk/e+wYr5CG80UET0BqDlod5MG
EO1Q/MqS7hpkCZoU9zAYs0pJfOyz3A/+unJaVoz0LgINIHuXo0fbIySIxGQJTFI7IezjO5Cwg+BN
j2Lh06ODSCY71K0kr7Bq3ZqjC/huY18HjK8qa2kzejO44WErjMhw02EsJokFzuL7MkxdFKMELLfy
XgQgY7WQPVuVRAucpy2b8JmE3f/9bBj/jytvYh8DMTpGXztMkKl+09BxNV23PJJ6A5t2VHAs6Q0z
DHCzeq9cqvirWPhzBakWbp6UbpEftR3dTYYJgdkKk+HBJXkdc+pXFwADvUu5jGjkBRm6dnD2PmJY
ZtvumCmQ41703bMYpG0VX6yqxpgBXij8USpW+SfSf7hX9+qWYHVZhQSDWdoOFdweBYhZQeeSyc9o
IvT4Zaj52iWg62hKUWOFyuIRIkTq7hnPIbzKUCvezYC+ncQMBeQhUTQ/3UX3QGH26ujSHRDqEFaN
kgiGQtXPqhCZyiIdY3KtKM5bYkhKqlJun4PtdSrH1GCYtZRrQex0UOJyjclEUOQx+yEkjwuZxQIy
OwXGWaYXgsDbW4iLjYalD50mQ3rh+S3bpwQEUE52pjEVC4Jplkir52ZT77pT1ZO/42HcGB9WXUbM
Dm4VWN0IWgdwzxqr0tEye2DXtark62REyMdSDY1IjOBnsORMHC0PAnvPsv4pltAIYXEypCU4YSYB
rb2lAbIK7EDBLNsohpmiFFz6FoiuOT8R1vW1tnxmXA9JxITRhB6lMhQQZSf3V0knLrFavsBTQeDj
cyVbz6QmFPGfPSh8t0bpb1ps8TAJZJVawCD5cNlT4w+UrnO66jcNxXaLHobmS1fzDAG17qcZJEED
WWQ1n+0rW6dDyYkgKyVEXEL8SckCQ+EJa+dCfBbuO6XNhO9MPzWbF+nHEz1eMFHv1GO4ouw3VSnI
ocuojqdJFK1yrLpvbmdUCITDl6AKOIvEMXxonXprBF3kM+HYbBWtOb3SI/En08CXvSXfoMA8pPd8
PzPqAv2gEqFHp0JKjdSImqxV4H8EygSJZdUyoVwD7hcyzyAtDcOhaI2NfhrktBTizWNVs3iP0i8Z
QprmKn+XO/mG9xJ8h5LTuWaqgRgDWuEkp5EcH1RUBuiWZ6ftHcwe+wZrL3KDCV4pcPxNHtDMYLrY
CShhoUg6u0VUf5hmM/RqNJCxFF88iNVM6GOuiILoSL3IGiuOqxdqLPr3xZ7IctRYYyyDsZFwVzWK
v0NcswQ/R+flblY0SsTu8Lk6EH864pC6dGV23ejB4UW6kac09u2LA84BDmrRWbPSpJB3kQpdaLXD
Q45QNWbrLiReGxFPJ1m7RtcaBONKPwdtEaPYEWfIv0hU0zglBD6EHCS5NyNc6sGB+USMbIa8TlU2
PITik7DP7QLtYSqR9zvuHls5JiD4DPDZsJcBu1sR1jh1OmJd634Q9Pnl1swZ72WbU37cczt/hQFm
zB0bNhQ5RfE1aG1b0f5UrAQyi6Bq+rg3gQdrQi5atjBPGtHmSydwOM8Mck5NNuumEKRqui7InQFi
MCFHVTV+gVKTJU2NmYrovDSob7u83AXU+9ie5sFPTe4B+6vd5G428ACHsjSNunqu9slw4PevK218
4jEgNJiKIyHN+dnE5GnnO2fbkqThK/tMwMeFDIWJCx5L3f022XhNLMECoZ9sGgPJ243DqVlTbgI5
jYKIeKNzJ98fWpTIQ7hzTYKwZkn5Es13nDnvetKlmGE3OhIEqXQhOJUU6gD+edHNOp0f/ydJk6iR
1yo/qkXM3LN9MHKUvgq8gjeO3StTiObFP+GcjzfH1pIN9ZbdgrjNtiNuXKnWuVIXsThWKf5hWn3t
nHWTmRRkOpWLcZyY40u42vJmuK7rRGLuEq66lsXF6Q8t6F0SfntOhy5rdmFB0fYt7dQkW43kmLDj
CTdO/LtttioFVDo856kfEFJxtyBz2oBs0V+4PqvWXueAdPAikrYoT77o8aCItc773xnZZz4DidrI
kgrQv9ooCWzg1fvvOh+287LZXLcKj6QzuMXh1YjUQyDzYoVKYkZzlu2SBQj48EoGdzgg6Xx4wQjL
ZVe2czmGBdSZ7ir1GfiBqEOa9SX3IEp+l+FH3sFbd0zwZo7pJGgeemmwSHZ8onoS3zwHR85nqBUF
sYvhVG6UVjOqt6hRM7HWLIHfvR3d6HI7W7as3knIFrlXEHvpsnMYNEeCCkUOxcMIZKZfO1UOeYYn
pEiT58c/UVt9JsBio2ZmYBBd+BASGoCvHL0phXlxxEYIWo0j0SjlsBoeTQwbWsxE0lmt8nSXBXS5
kkJa1rvstXfMevJ74JIc2VH3kNGOc7axM1f58ocDE8GUel5aJFZlM4hEM1GK/5+vBLJ8WEazvZ2C
s+590i4MadxV8zVy+krJow1nbfsJcIRsCCfM3lqo5rBbe2n81LhId9nJlMu8oKKBla/HvRaMSb/X
l3WCNyTYyRRKYbk9YpiE+P5cilAISmooxXjd7Ry03Sl3OCiqgatRK2bnLnCbInIOEDKw/JakklCO
c2AM5yr0qMOBCSyQPwPpzSrxyHo5Zxtt5i4SYuVzJz/5ydf2gcIJCLeNDz6yerThQqy9CeEpINhE
z+nVlyOES/bck1FQw7KbZuPlRWfMhT0xHrfBKHDs8jzgZ3uq54oQUQzzYK+NlpnTPzq2k49EDwGD
a0KVhUNEtxe50UCElpVFxaxwN1ZkhqeKJwm1vPDJjnrpguV58a3VSZy9yN+/hLVZM645RHOC6BIF
S1nHLG7+1Gh/cutqe5ZkjtutjR7bAf9nhm0DGNvJ2yed2R60kHef4kRXhdfGAX27LPuOXZB0nRD2
a1Pw7MaMagBy3/GitWWl7xulcpr4ikij5JSA6HOwlg1RGpFVFb+6nOCzu3NuqAU7sMT8GekI6oZ1
v0tc3B9OxjlUWmOoM60SbENWn3l9xb1zhRTfntKSJWraYh65UwVZK9PgvyjWpQWvisw/3+4Z7HIj
Nd3Ql50MJW0sYSOtYCul3NTxg41X3mwWG5fUMxD4rLtl13Jewp4T4uXvkmEu8yiUk5mo6d8zhT5r
IlTCKrSd372v0l+/RNsRPstbH4EdaxD3ocyntQRKhytA4HufrtTesDrWe08UyKUE/qWY/4RvkPI7
Wcs3ryY/j39F80oPlfO4U4jaGRz8kbj77Yc6MZfP/mvmnhowzxdDg+ufUntDcIb0cpl9TJgEN33f
U7KQsNawrB7xWHcIJ4rMVAawC7hZ+ixHurj/EYAkdks78zPLciqPE8z4OuCzWbclKELscVGaoDDQ
75gqh1LQeT6xHn09ZSLRcEL2B/GMrCuO1o05wC8ei21BvWZaTK2K/IJAtiVv+6zIQOJ8ytStY134
YwDWnkp3N3m76kXcJl65bz4PtQylOtMk+iJF7alQyvFFFgH9/3tlTH2Z/d7l/Clnox+q6xdGBvHp
ojZwe+cR+4yTp7zsAg6Ud9iz6bYQw0ub6YlTxI1G8kgloh8KWz4AhPbFY6iLGGShjtAdrpcjT4Bx
MRTA3vrzst3LiE2iaMv1flOUckCmjjSacaKMKM+g/SIZ1Dw+5aeBtN3tbM7LEdCrs57uJJmSEXXo
LTrC8RzUEuXw4MweL1gHOkvIUEE2TcdQO15NniK84pb+lvEMrSXRB8iCRdzeahWeBW1oZRu3LsPm
Sr9iasGk1IarVNDCFK1TpA6fgVBTh3w0+D1vTuhWllJow+nF8ZQHqaUT+izbQTmX1VFgpa7vYYKx
rQg3GusFzX02sm6FSzwM64Gw4VbFp1LAPbuL6q3T0d51EHqb9s8qRStFc6lLkbN070vmHyifBMH3
EgvUTLHCfe5WjSL+B7VEk534h+u/O0Lx8ZGbfHxk/a6R5aYn45/x0yu+RjuWnc5T91T5cq50/brw
e3cnWxphNA11J/rrLluV147hYh5LKpXR4GRjvK6lnRHU96j8L6jJaKcPiPosUJztzoe271MXXO21
R61SLh4Odrjaleh7XlAQoDl8pR7cmNCH3MFDg9/Ck+GV6KKh4dzyyui1Kj3L1j32o+WMXAX3hwBs
L6P+gpBCI9WXlyvWDTVcxBYeealO3tEuPu9ymB7G1HPzHdDRlntAyg5bWTweCWsEGsVYndiB874q
BcaMWPkbWNrZ40twd9GCtHZlNhBgTM0/zhfquqD74ovnW8GTBV8Su2HoHwWVkrtGsz1+AAhvR0+K
7vdgNW5hFfgGfnjCQxkrNGgUnywQBdx3N+tNJUQzBthMY5kn7/T1ouwAjgMNa6jTXMExE9rNvlOS
bkBMIq++R8Hu8kCfe426RWOTKqhHrvFTNcVKRK/Sktmfn1Dq+7ZLX7MatOpildR9bqAN/V/cjU3P
0Pbw2YsppOj5nw/lpt3Ps9PKxGWIrryXGZWFXOelyfOOxsH4YqbNEQPZCInr89cu/LDXXOkjkI1N
Ct2ZlSaU7dX41Z72b/IUZfvwssVitG5sHc+as/sOFy0QuahS/dULjul5DRL7qni/hrMnJDVnqJpi
VpUwHf1dRBuHuZjwmGOpkbAdS5FTXmUnHIg6zWHmssrP3FLsEyPS/td053ZR5GyxnzLHs6NZX7VP
MvCzhEbZLrU1opdy2vgtZLDCn++B/Ny1YVoIpWOJX/dXEBplFaYKEeUT/iWhqrO2yab0Ke0w/mG0
+u4AaojAYD5rIlRLifdMsPRjqKc+hfmZCHUXbYHFjGcqc9xvR9UwVd09fqNn5VGsSpI8sDu+ZnQC
6hKsxRGK4Hn8luGg9Pf4p2Eph5RMpdYLrTGKIz8KnhpdoNeUMJaO3GHiVlzU2dq0uMWmlOWfKG3b
3LGfQbNw+VtcVTA9gR56cBhDCRqir3f8iFwm07i9gCLl/OYIy9ifcEaI9JrxO70zJ0k/xrTuMfdQ
RneC9qppKHHdYBAp+4ki+UoPubCxQEk0vDivvHeZXYbvvJ4Dy9f2mvoCUmXGnMbAiT2qzL47zJBB
0F6R/ntcEn8hcQ4IGOxYhVNKhVGv2voYS8fEwWEijUW0wHxTP2LRGw4CA51Xh5Z/JZdzZsbmo+hg
9YRV1TuV2NRUCQkkj/Sb68C9Nvp5u38i8CIQNjUxR/um7YUhI8nWkGXYdYGlsYoN3KgaxT4k+uQX
IKXN09yHo0A0//Az6W0BBN1NCBNLtvbc7pQs1Qeb6SivrWqeCbW39ufGCiy4giBWEmev6/yi8z+K
hUKusvhNXol1AuPyygB/k57Kqj3fabdry6UNSTPug2ODckh/iXxrTvLfY9lZPRkWbKUK0/YQ9Exh
l0gzTECYDKrvpze8zv08u9Wrj96nBa3C+q/MEP4D89hK094AAl2ZaZeiDc7+TJi22gPMZw16iFhx
vKDkqz7h+BJVSszQP6sFy+uAyThn+UXgp+rXSw6cOaoqdGi6EwZr86hEr5q9viIz2Z8SJL+wzKTR
wJamq0IyvGoBWQOxvmvD6tW3Xiu425oTrltvlAbeFSMteqn82+TxhBqJYtcubtSscNJl3srFNnD6
IUKBf+IypsP5e52xUOJQk7fQDpP9+R+gfv2peGDGeR/ZxxrnC6ak6k8R1XCCNmZ/ZVvD23+w2+id
kZEjvyRzQK6S8lqCG7NlkO+2/cX8pfPSG3LVuPomGcZhZS0TseDMOIR6Fmj1Tr/v0XcMEJIt+2qD
vpWLMukSgcNUouIZLSYvXx3hNaE0yu4ehUb2ZRPVzuU2QeRNrKEHkv2C7/rOYmo1PZLEK+TBkoBT
AEKLGpKiThvyTUKUSYA8WeSZpUxtN9aRQEEyQ4vV/AqIxgb0S9YcU4eDd3SX6pq360Bdctx/LbYa
E1yjx1eLep0Kv3eZhKLEASGfj7C25xunHF59BkOjzNxo8GeGbhcxVjCY9ZZN2LcaUM+kcDLctw+C
wSM4xjzBumtdP56mqwlBPTYPhsdWV/TCg2UGC1meqZHzovIEFjkzubWTcEOWFlvQnWkIgiLGR6V0
BBSlUx/j/84te7dlad28NVKTIxMKAXKx6u2465DtWQ7eJoLCR8oTIa54S8mfNh2bgBNYJbkSwlIX
NSwi3wxNN84y+qcsyXa1zsYehJAzKpCHCGOpf25ncESgOQc0XD+yvvNY6hOysxQ2HcDHdGfRG2Iu
DrnrmpMbHxRNVqVe5ufhi5hS4hxABkcKYxm7LWHTnEU7KVpAU+DbFTiogzslc8Tdv2vH8izAemhq
iE9yc6NyOO5vuzKpVSuR42wam9xJc7XK3SV1eKYS8ReVaC1Y9VlfshpJooY8MXC4nQr51XKQsnX8
+IfSx/qxc97h2rqT+Kc/61lGqEo9+lbH2KYA3AdH7RSz0ReERD8/WcxDLImJAFJzQMysR5Zso7p+
DGsxe0gJRRUxp/5s/0JW1VDQWaukYsaODwgWyPrMb/EsbHrM3ns8JH+sVGKfZtly4OBuw5NWSPUB
4X1D3rngp9ZcjGaJzKw10uxk8OB3PgZseKcwjWpBNrrlkJHPulTOkyt5d/29OPu7+xJ7yksl5v9B
+BNR2fgVZV39UUFavjhIoW+twDe/tZiDqb2NJofEPK+pFL8czaZnm0GEDEgcUhtaGy/A65sBCRma
67VmmXvE5OYFT244M/qaHpl75EE0Odh48FPPyCQ7eKjhnQ7BMOfwS0c4bz21sWFNFHJxr0OhhTpz
UOmfskFk7RYA0C7T3hdPz2vl79oWes+aL2t1kHe8yGDRC30B6kcWmDJKi33rDp/+SpAf6ZFn6D7z
qGgru11LGPTpGK40vuV6Es2Z5fQNaGvYDiF4bnAj/kPCudQHGWlXsVLc81Byn3xqkStg2DXTteG+
1N3FftTsW6EG6l9av/h/CjjAZ7ro4WX1/ROsX/65HZyJz0OeEz3u8tWxjNk/ZByaoZL4KylfwQRN
NASwBxdIwmbEPy+LN2TjiEqD1C2Sdk0lXkFKlenQXZD7RQjwE/xgQW2ye4zgKAZrkq8yM7rZ30Zq
qA1oIh1y+HyvdD/Z84sDYRY+Xmq5bZM7vj6F1olH+KENd9qV1uGZ3fDPhzZwWKgWvS/2++rK0GS8
pUomRKrMU0OKL3K7sVZXfGQfpSOITZpE/Z5WxhYRwUCxvg/1GAUJdgJYClREUt2lLmIE078qo7C2
N0WVuWc38/fuMouPDj/BRoAE0sq4PiWo8Wf3Tb2XGTR7AcHyDk5c6AK8w32eN7WaCmd6Bs0OHpod
mhSMbox+xUJqf4tuMSoNxuMgbuY/B3AU8/dAZRUUqwSORrcDJhAk/nHQcNwNx0SxiFEa0GgZfxNU
BYHWpFVC5hhJOnGdRJYZiZFbuz/BzomKSrbVG5sxFUmbZ4zZrH3RSOi6RHGCVrwcO6MO8truYPEL
nRUpRkNsrTbI9VB5oCkG4gxq5WbHdq5LhP5ZGAi5B4fuBJ8/XAklJYhqhQs7lIQOKYAObwzvX4av
Qx5DT+s1gmon0ZQW55z8it+Ft0aOdLIbFvBOmeJl88ETgxWUdDItgYTdaZG37gEPPBybUHsKO4BT
gp4NfyM5PQVEgc+KqTiY6fcazmQXeG5RhesvmATIjK16V+DXL5WiAra0CCzu9dXr58wZSCw7AVS/
kBGUHe/Hy8Foow+2/DQ1xPuwqEkHnbURta8Ix3PBUFczKv7uitv+XecR8r5R2JtVjZ7jBcSC1nTa
1MRDdlWzpfAWpawQrKxD8SkuQVwYkZEDga1jUfW9RvaAaG8L6NgcgfvVvHwnnhYiNjd/6tPvHf7w
W3U+fHHhIlSxPeu7AL9mcZL9MAsLJIF6Pancsok07Mtf5iQgGzYfVf1SdqAEzzCrZcm7gpyv8qRh
q27f3NkN+kJW1+xxVyO5MPlUZQph8bxOYlsHHB7DEGOK1WeVbTFvVnKWHCIQ8YAM3r7XXBsicS7r
PXdATMR2eldZYnMcRtdGH+KSe1Ju6gTDt1PGjkYmAq/CnCv48Uh04ZeZoTwLkd9NpjpLZioMweXh
eoJaY4YnW49OcMxFhU6GHVnOLyBSqN0ErAg4UbbMmXILpK3Dm9vnokxwus101nF/sX+H+IonWAgk
o8HDViktF16J01/UvuWnyvmcc9B3Y3hP+tBKbOmb/2BNUWOMgBt20rL7BtqogIrMOULHsgaRg34S
HzbhhReC036Q5QGc5PwMP8uOTzlL5VKCu8SKWf6zDXMiN5XaW/7brmAmSyN32PloC0gdOZNTCTjE
Upb5zJ192wIxH46ukL1XeBR1K2BgKlpdU4ZracannDpEagtiTtqnkTT3+kpASvDJj9N0LXyvPT8M
REq6qC9Mz9cBYME0wO37K76QHSsCMD6lixNcaQ0YRIyu2a+I6xqN/TpQIkkg1Ldb+vitM6jciGaI
z4JkPuhNP7tyv9tKZx0YcqN6hHi5c9A/j7AS4wk6bj5vMwRROnCbCM6T0P3E8QR+7fMuK5/qNrGq
lCkTPYx15dwxRL7c+/Sn18pSy2DwIcH4HI8t/38m+PykU4W026lBWfVfsF0L8+ccld584dQGifPU
s100JPYcNppeffCqMsat4g90ABrFBGlz3AlghMfVML0Jr2OdEE4kwublLnwft/zdd7dbb07jaDZb
5mBMBiMAarPMJAt0WmiH+DV/Gjb8MfA7eQbYkSuxH+lvJiXdexHoZ9bnw7uQcDD0Bm24gLDoeKRM
f2gnYfZ87Oz85HibLJBBonvoDFdH36pvd+iIoYxpbfljFMl2GgoPayYDJBYkx0SqHU3IVyQNsR8v
iZibmF1QFFftcxdCSer5Uz/bAcmj3nN4yCfAPxteJUqKA2DNtlXYGfo9ODXwoMXHITpL3euNS1M4
JbqZ/UaC+eZA/5TPM2ujs96x/Qc4ljmL+fTGUujCPq1wuBtN5pzzot1NyWTPQqn9qnVi1QNlIW5K
nblFeoVEOuNe54eRsQe92gw4OcqI+nV7BHcy+kwOIpKlbyLAPEvTzRSAilrTQXbWgUanrNO+bshg
Yk/QhZsNEfgjBR24gUVcjQNOj9nUDo4PanfKNapH/mwZfTEvm1P7l77C9YQ8QDadhX/GCF5b9g0S
hdY+0EqNG0JnPi9e/LVJv0eh9NdYGlX60kHDe/0BnzK2OjeEYmqVgIrYGf4YCxb8qgQiZ0pwUbaV
ptCDqnG1ZfXobj2lpsU7vfX4qQZQDcRxoWWYRgkbK/OB4qhc3MhaMTFGDUBdvPd03q0Zx31wujt0
3+O7Aq0RiiNSSvQTukK3nrPB3VO1M3Ie2vmwy7GhXgMya/jG+93sjL3L+elYnPKopDOiaBHhpLtu
Dzsn85f2F+3eOwlR1ev0dFMNXx3AQQf/q0undLPetZtYt9dMSBOnJlcjuEqqd7jV7OD6YPzOaopd
KBiAxdzgV1L4KoOb+9rRdKUVrMUNW1ZKEbZRXSa5IkBTAywMyazkPaH9Ewth0C07EOvsakwUqJLk
/PR2XtNMI2LteAmlODrGUz+bfMQjZFSGd78IKjbPLE6thmoTkBzh48mX5BLP6NLEttGy9+CYeLVB
G7Ws/Rzh5AP6qASyqcO5DFlik4myfkv/k05qYmS77yyoxM1UMQrvhLAc8eEfWu/wVskTJBweSIJp
Lylyytbz/PqjMt5vdtt9jrNp5V6OejcSdOyM3AK4ptiomKSV+AZbqd0J0slfFzCeVkK655Hcqe7h
nWbGDe8Ps9B2PM1RY4LEihJvJJxRrseTWEYtfj3btfGloti6NK9cLQvX+egoJPfO5l86gyLEeRRM
pzG8GtcdnJrx9AEpDlYDVBdIpYZ/UlVJWqLi3Q8wmlMH4kawRm5MHkGjXvZGbY1M2IavZTietmv2
6DX25B5AmFc3xsexJW/o3jZMrTGf/PHAJ71OMBmgStee+Adu7ecqwrTzozHwb3gLqDt5QWxXRMvJ
/lZ8t40siN6hsrqeSY7B7qQbs003Ipbs9m6tHeh6W6Rb9Uobkmthul+UuEnBBQnd4hBxoVyfq4gv
OzYHg+HjmMKz8YJQbpLMpWrCZoU7ZZFGchnc7IbchHuKx+JrMj/fZUDFCWo1l1oU7+8EjFXYvxNe
GkT06zTYG2U2BehjR8pivPJVcc+vJHo1KZIfwh+32cA8cwH8QKl9atMA+BNcUgZiWZqrGMBkTWGT
bnNuavJYZCR+8IbdJC/Wi3qnBfCm/88n9LtUmFQJfGKjT32G4kgQHeJrilN/rAGEPwM91ULjivBs
0/GYdffG9ddLKsr1FhDJeKsJg/hXTxa4Je+6r60cPhvgEVkqL2rtzj4hHYpBdkMC03FOaqAqxU/B
07nGAAXS7cLT+54AwKzV7Ejg41YP2h5RaMmz1bhSX6b2KjqvPDnAZvmefpmTKQTNZ6+QrYJbXH6p
Mol/lw4hIFBRljsKD8oc+dFYiAYowVEA8qT+VG/DCmYtOfEy7nTPxkgDj6hqUSWth2lHcTOgtoeS
LOO9BcGY+0jp6JZcG2EhaphKetqsTgzh32tTF8q3GEoe/kc6FgPTijCmEY+YfEejmokWrl/Xf4Ht
vT0tzguvr8r5n3VaWCm1/QVznFRBVcbfeenwDfRSpL5aThM0kJFAdJPh1txThi1ZeXWDfiGUFtyA
Hys1odizewrgvF39Oa9YIEerM4oCrCKLNZv0/fPAFgTYwHA70g3aE0O6PxFZgWPQsX6bM45GL8xS
uvSNanImC3QJvDHIfijk6I+Eno+kTZ/gv6mOpI217NgGxKa28eV7ON1g7ZX1Y/Y2EjtHDmHSSWbv
jVJ+zx8jdgyIo6WTLt/aGhAzRl3+QBMpY1jHQs2DNy2zXqrVl+VyvVbGnlKu1WDeYjlIjyPhjhzU
RIK6vz6T4Sj5jielRqFzIJfb4ZgmzVIwf53ZdVbZKVoVzs0pCXB5KtuAluNMm0UtMVF1vWkG/31I
CRrvMhYsoFLGmRWlR94kEZrDrhjvnL/X110AZzWkAPbte6x7H38EG/MvSLsu2zXskX+9EKIppcMM
P4Nsxd8a9DDhdmlYaV4+phcajT7olWP4oBg+YMGDEadnhZ5jB1iInTZDi05TiWWLT4iuYZ5fIy+I
H/z4sYdSWdWar8KlTg9e0en9OFhq9nfbbbgn9TIjKPXtKAp4GEyE6QwYEPYS91tsDIVx5TZeFvBU
AT8g+PhSf2nrqazDYZQ/4wy0+FTPTjot2S+jG9ccYnp6h55jh6CPpOXck/9EXqzwnOdja6oM22md
igI5jGbpYwP7OSYgYJDRGQbuheAQwOfGMgodmCN1GdrVKrqxYD+FfRYhxo0G6HyQtL3Jq17p5S41
qVfWQQ9gV6GK50JWD/z3jgJZI16PZ/U4AYl1LprlwW7XFRPQAD6hVcPNuaxn1V6BUnaFteUvym7e
UpyO8jtPg1ZsdyuYpgaqZKM67V6HwR+Xh+BFDvf5oiZynpy+xoh0goAAxjY0HuVJ19/OFK1Bl5Gt
xvdTrlfAZsw1ZfzfY1VGW+ovfyP0qHUGpSsywGqC3Aknizze9xQMwACPeOLUIJVcM4QRVIwZSM6R
W4/CLrX4GBb6ytQLPrRPBTcFOIbgPTWZJbMcE9bB+L+FXUe+QoWtIJ70jySOnjUa0pCty0QjtavV
EuYYdX/Q/SHLFflhLZe9EPq6K3XC6iJ5WPty76V+aUGEH5/1rvJVM0cHvNsTNEeGt8YObHYw7dHt
Q5XX3Z2/an6ADDReyRTYfd+XQgy9qybA2j/mw+Vixyve7sY2VP/++KPaum8LIKpyQTh6MJlGf2Hy
7b6arNK9syZ/ikPYeX4mRTENBy8ztSkgdMqf1owhoD58fEYOuiCyEXcQcP90G9wlc70SH3D/u/5H
xYY9VhnCXZYvH241lUSqG8UMolbI+jCE4hQbO28r/L7mQ0oUZ6SYK5H0Vf2KL2M0yHqU8TS9d5Lv
3P9QxgBRIM8TGYmrlupfXWD4gs4tvfSClGs7Zy6DzkW3LG7ReQn9lJmJC7vUx6bJPi+fSG7k8xET
hBhZ1zjZsUjLKT9StIUdqoyQfDPMZq8IxOrahm4FDwG3OCDIpLp77RPVfCO4KOIXJ2nVdB+GFqyC
Yk9RF4oeoPG8xiudSzuzbIbl3SbZQ8mYhOQe1TJrIXz77OB5P95ZXzUDDCCbRBP/khbTpP/MF4O6
QMTUYyJETAuxki6jSQoCzVdUVuqjDZzxFgMof9XsrSn9dxuFIklcL5/ThT8eeqWeNLJRtjHkjiHN
pDlkL336CfFgW9FKEUSgraH1hWNGdUgfO12dbh2Vc7YkQW6WAKObNDzA8VJB23G/BDBA8aGVbSja
SyczcnZ3YsG9bOnDtzAWiFqhdhQpIrLbLea6CYRKjBtjGhJ7n47QW070m8BHzMhEcFiIg0cf3MRz
8wp4QmCvg+0pcOtP0QYs58v+jHNjGPEK9RTjaL/+zdWid0zh/f3frnEkngV9KvuGQkU4aqmrIC6h
4aRmGy2L7Bndxlrzgy8Hh22QB0wMqVkrGceqFAPh25x8iBLXxDP1PPpxTYd0qq4MTo2UXOSUJi94
cQZKp4T8kYVmpMFECMkZvwDyEgd4juNMmC6Wsys7AB7Vkr2vJIKqYysi/Dh5XLo6Wqd/36Fu8Z7a
znMY/pc+zAIV9/eIuN2PT8WMnI9isdVbjqqZla/Ab9sTXuAlbGl6Lacknxx2yKr+nOlqV5I0R0YH
WP2qgchp/c6SAOledJLZ6dtMHfkjnuWWfaAb7on9G/NxWIljAGlqol5Pqek0Rp4j+AVtdmhbSWkD
fq5ccJ95wfpVzBNwauhKRzvcV+RJJ8IF713KufPtMAzNLPWUYKKfidcnlUPh1yS5BXKoa4yHEp7z
OHsJNM5XgcUtKsrZ3vrov6Uf15bsbcnYvuobmlS2srg2WhNxFG2MLn0d8I4hOLYAz2Bz8yo1cE1C
aoVlinzRC/KqZGjzMRGiUvwVVPxQkp0343pHdJlj4l7vUVezToCzyDMQlSbFh5h+9uydTpSOGdBe
3Zhu9IbjPvWzMaEsiXMB1N5/nDHw2D2IZn6i6BKY6vgBGvZtdvgV2DIYgd8dLiTRjDIJhJ9XNR7K
q1CmLV1668wHl2q0h4qF2sZTCLY74Bq9cU9Cl/m+pm2XMzs/8MOzojlqPAnVqSVRuCSFbf8Q4/sC
F4ujIZYdNUvSuk6ZUU5i+eTzn3XzCHqDtS0L0R8JjcbnvQ9J1Hjf9aW+v7VcHODctKFgPlu/1uoc
B3m9NPdyKukzieTo2E+PEhK50nzPPY7iA6MbeCVj5/mZMZiEZjonL+21EqxvZLckC8hYR3uvPb17
wmcqgdy+KPSeLZ8O28EJH39SMHaHONqLDY9kN0GtgMt4/cOuPsKnwufCKk8Z+jO06+pYwM05+PWi
iDE9wyyn1tI7SbHEZJ7mD4/gE0Iro8KzzOt27SM3Yv7d9bPol9OkDZOXLD0Yj7SblzCEHgdJ8cBL
vXPLSdmg+G6/O795wN+MOFXOPGJAwq420LOJJ7grKAWrCagapZ2Qf/Xf9BgKpJtFqTQGobio1byq
usF4QISm1L1ONzgC0SmOa8DJsHiEkt98f75RMVwisyWW15vFo8UAFzYrkG4oLAslPgJSvEVB39Ry
MJ3XSP7e2UEnKbPySpicY+imCdxaofmMXIfW0CqcAppzRXfPnUZnHKkJSrKIxAZLGa5AiwRdHDMM
FZ/sGUEHLHrMStlXfnT6nMgHb+Jmv36Ppm+3fA1o4tsglVyJXAhDTrTWrKJyueRmmz7N5itwQn+l
+t3THdT8Pih2DgroX2rcaEKH1OG8X8CypZ/zKVZfVS+HBXT/fJycdVXOwl3lOiaQbcf2Aq/Ij/wH
r/zIFprHPhyoVBajfQERFC9vv4g2/P3wvzpE9yORjjm3GPqRjOLRabYysN55b9BwAu2998VbjyXa
g96h+Os4226XGlLbhdTdksr7gWPEqWaRmPK50NdeRVHLgh1rsnJRxK93M6K2ixd7lU1Ak/OSxFzc
wGanrXAzIp+dKugxiNw/O+oOLaP5fWwLOLCRK2No4IR15/uJPa8v0w18+alcQdXEVJGIjlUctcsv
42Z/APO1pQAkiqPYIBG7WSMmCkLfX83n7G5CoWBDndQegS2f0KI9BFNCf2Gy88nDDEv8XFrbKyu8
Hx0zOemTX22Y64jmM6RI1dnoCCtA8BOoR9AfB/0vWoFX7MV4Py8Hi1hZF4u1ga0OONWpj/dc7J3U
fHS3fuZGQHXm/0sCt4dlkQWmSVwwRXiPIfRtgPaAEomte15WIKyGnlGYEnAHlRWOuegL11HpszHa
t9ydojrSwXjo4ARooJdDRIjzmpr8ie8pAWhhnkVLPiKJuIzxU/FGuVIfpBlsEdjMcC+CKUjFhVuP
OhFUdufeMMMjpOt081a/fQzj5aZWuXslUHBBy83zTUyAW10bndhXyXbLrkeDEGZTMTMp5sK2WNvU
kKFdOqKjRkglxGxykMAJ4SwzZZi5fX/Q5QGy37RP0cKHoxjZgnNyfdDkkE4g9P0n3AKFPBp1UT0d
xNYxgGPPJz9hOLbV8l8iaj7xxXxmuEWgBuAmsvHthNQI/KRHC3Q7pICe730mgX+C8Wqp5qgLxBY0
IGnSZmEiXqD9xwurLMwH4sfHJSnsmIURfld37t3X1Sypp6gH9ahhPEFC/NnhXYCi+1UFmidXqdfb
LpXiWlXpjmvmekSXwXX9ffqdUg4ujNd3nkwnITDl4cXG7qz7bnH1kraUoIdGdiUY4K+7eqwFAQ2F
8SlBMPn2fL+HuH1YVIKE2UzeaT+kfUE/X1sHje4jXKA7C+ue0OqcWsY8q2IuVe66av6tXEvF3Np4
NGv/6dCJkxVmaOWkBusIbLngxhuF2roEpuD1TgLIz7yeO0zWjGqkSEwylfGIbyBuw1a+cExgIfJP
wKMxbFT0YOYztPxFmJCx203HJOwxN9n9mVVc82LszEqKVumfHZhwnN/rE8NFgFz13HHaKU1MTiSp
l27T2e68emsjmmjsyBOoW7EQnz7qXF9FLDK0k5PJmQJ24PvVdEZrWaMiYM1pBNETT84lLsKyWCl7
vvxXUsOWRVorEXiV1VxI/lEdQEUfLFK0xiwJsth3fH6unNj8438OzNTCnt4/Qa8mj4LM6FY3dBtz
KSSjCceLP4SroUuPcOpgb9lYvviVx1UVDs9JITryoYuZOiJkFpiKvb7VA0Z6oFvc1DcQvu0eewMz
Oj3i4hELNOOBFEzXPwBKVUwdpCILx0rob4/v7K61HZ8YB4MJfrDqkG6e8kGGjYSP/g75ijdV1iit
vgBJQJwi9K39bktNuJi3KadreJRG6uEmGZi2CB7kc+EPc1FG7eRiJj8eEH87pNwVNCOUrM3n8QIm
rc0ZRd6n7OgB8OUaQi7ectsL2cdr3n+oogh6MhTXmX18Q7/wlqBKD4m3i5RZKph4ZUvLbPFSMm/L
iTVqNOD0q11LktTj40jQwuso+BwEyA8UYk2Lw23zE+YAaEc+hShbvvsaKP4eZms98yZaRk269mCV
+MhWmyBB/HKyFn2RoEh/GtszjLpBTMJKMkUPlnyYmn1lfCUVosPQAHFyOd0BVppQf7Le7N1RrhbT
POd+1eKEuLlcWIMFuWCg58XspfNSZj3795emdxauAdg+/TD2NqsOvR2GKDjDJtR+U1Xirqp7p02u
Df126v7gb4+ij/F9v5lbp9mL8XfjkH53NnmuzLw7IkJ8vgJbmlWfZ6YR4kKWXJKAmVfPXdtZrsJk
NKuqt7GkvQIdyuW2MBVJ8Lhf97xTsVNW+hH2/LvqWxyWr4NPm4IjCp8W4sYRwmYL2OvAhyidlG7l
ZF7MHNQHBryqG+hEKdGQD0tV2JjffDuNvliN6R28owL/iI5eIJWzaOHxltHyY3yV/OsdYz9yqFlk
Gxm9Wv8QYB3rxDMAtGmAnGpPVmT8DGLmfZFNEnDS//+N3ehY5bt2/8dnRnRFt2/ZqJvU2ykyGx7X
VgAovcP21GDsCdaljDp1vWXciIyDIEwakL0CumztNwL6CDeCbxfJGzzG6XNT4tytaP8/xYarC48j
x2B3sfoq4vny2CcL9W4MqA7FN2MYiQtsJ8mUbIQQZhi+TCuLzGKq8uwoqT02zRE+3gN7QzwHDQ2y
7kEigNSGdttKHnHpOU9TsMYfpFFjbRXk5gQKjeATDPxerZkxTEZrLLEAMIYkIFtyHCVdDvhKqE3c
w0QjwFmGveJ2BKEbQrD75BE7sk7rPBwWXY7EsoXM8i7v7Oq17VK5WsEvn7En7TUwq0P5AgGovuet
FJ20CIKl5rWjOE8Awl88dafrw42Ye86esiu62Ql3AWnktIfoGafOFRm07TzxWMJ43NsSzudtSyzM
ZVCBI2SWZKTGxFlJGChsjT4Oynwrzqa9RdZJj76JjYaHLpdUfxrEYUO9fNpZGCdoxE4khen0H87k
izigjokfquRTGgjx6hopcprZ3gVvwPlgY6IK8jO6uGe4LcLIvhis2Ywi/7laKYMvfTXXmfJUKxPB
Me264DBR9tkyllzeD0JKAVTB3f5Ap9Nsx1Tq65puaSSotruy8mG1B5YwwA0YW36A3R+Uoq6yrAQA
46KpPsGhJY6LyseCNI75AFHQAM5Ml1IDxMSdoqut7ChFREz6Jl+yDS7U+LLWTTgZsSdotlBcYj5I
7z8bjMpZXB9eNubI1RyFWs/JX9n99M/AFE40/2XRWZ58yCwxEYsuEhXbD4RNKTtr4uvYNWHNKJjW
HUGDspBWe95UMS3I3Twkb+1UldZ10Mggg0UJqeugoIJjHdz+wEAv+yEZOtX2VOiDGnOvyPVcS+UD
+RFJjBLebtMpKxIcRooYZqiSRWvb+1sXb8whTjoSS6u6q0VqdE0hub2ouTmVH6PxmzIVGuzZ6YNz
uEkV6BW4oVhyU6Qu+neuZ0djH7I/LTotjB0jsceMz6pl0vLc+UG5vs6MDdg3JEOc9okwAfdUs8bO
xcKKnlhQd5CnuAoriYyzd9iR1s3EXCGAfMcYyow/oQnOlY6V3ykBQSAvYJJSzguKqjucqosG6Qep
l4JFI5/kRd6NVEIi4NvdjzgKDhDhXmAT1tvQRk82oAoBuln4qH54FyqJoKjNeQ9+EkrR2Qv5gEE6
fRqpeiQtRsTxU5lx7WqFops/7Gv9cEzVhVDi7kBPONEgh3RVPhfrX8165XjvGst4OX02zaX4mbEA
FwCUuei7Ztp6CON6qrTmso4e+gi6GhnFE/OubPVEkyFD7J1LIZoVZxrdSEmWUWjlXKlD/yu+X54b
ZP+aBXmvIRcj9kuyax14dUezq5LKTmBVSzQ84Rhml3fXA9gW1R2E5ChkJAenCtFlNYBuOB7gwvv2
vB7dhTE5/imzNjjFikG8VrrfEd4ZOsRlykyRLfbPDtJCgCE61tGoZY3F4/W+ILvj5/H+13bSMGBa
z/JsCdaMCZZ9eLXzE2gezJoWn7cQPyYSXovHX27UI2fC5ngceDhFaQI02xp0Wp9fDxLsI71aHBqK
GhMEEjjvFzFJTA+6oBoGwoY6t3jn7Bs2TMfvHOqbvYpUZMorXZv86JkoRHne7mwuJmo2eu2czo3/
4o1Mgg4G3xze8mtP5WHtj5SBiJkZWjnV2nhCfBhNE3FBxdvAiVdSzUhS8nDXhg2Mhul5rMb6ag1M
6CPMqcomjM1PILN3TPfLX5o29wS6GREmmTKdZNl3FkFNyTXykCr5ZzzS5KeLSzXivAQ2NwUF9TF7
Rne3YYcelki7wq5SeVQuubgGlrEJl20CAjEZf+6gzh2mibI2XI5ukWw5/7JA18Ya2E2IHUXw6wad
QArHiJcwWPsd5EXJ52pDrQdocCH87I5RWJib/Ok7Uz7dZYRQJp0qHHnI6mx+KCHff9oVIWhj0sJL
RAftkIhu7xsykclv1IhL46AdzSYUCz4a/9lhI9hTkq5+50WEYNTVw96I9BIXBNDK3KlafXOemY65
mVf+04SFvJsIM6Igh23LRyCmfIW0g0l5ayMSXtyUJ4V5SqE5VDMVEpIN7sXCvozbUjk1sB5DPodG
2JAt+4Nu344b1ETayK/wD3pCu6+V2JK9kgEwZV5vOYtVyZ0t3k9h1VJl9H1boHqfArsVLHliql5Z
J2r62vB4iaYj3fhsgHMXEi0eUiiojGCss4cJL/TC9dLoa/KDubKE8aBdGFac0Ce95ojTUJbWsI5q
jTETSBdnO108tSBLNWPzxfp4NZSM1MULC/ib91jpJ2ReL9rlVrPEDt1uM0uHZpB5GtrYIPsKePEQ
8KKCenO3Y0x2fA3YA933Bv7Gf3qYNzVFa1O6fvCamZ31QepOxxkNaD7PGHm0EUB66/XWu67RTP1b
BYGbcjuHm5VMtTxF4ERCEU/Cw3oEsj6CHxe7FisI0Vy9xKufFgrCQrFRiU9Zg5ynIFGp87n0N5TF
PqJb1k1LzrBhzfdJkDRVANfUR8GPlCk3Qjhvv05lI9CrYqSR0Yjr1sIg2XTKAdHknHcaohSpEoDD
MRBpUL6OlUw4gNVNqM7OBx4TDwB4vzcfv50wHnhhm9ac6Y/gjNxEjG7V7qWINSaKZWvIRLBcLNgA
lNJmkeRk73quvo02BeuCSFgFfP4lGm+ShlnYI+wjaKApiBQKGYjNjIukmn8/iGuYz/3Z3cqXD6kf
gqfl63l4/QjhmKaYwIgiKxzNtevA0tIEZKZXcQr4QozFRIhDv+CdDZzj8jRq2Jp+ckEHRxIRbafz
ddkcbyIlYyQVPtb6nYTZ+1Jgx6pUsqhuK7e0XXjfKghpyRE5xD8oHvnuNBz/P2s2y9e2PNAfS7g+
HUBFm+JriZb8UbOYxHaZ9l0k5LxhPnLxLshk+GTHtooUJJCIiYn6vaVexEJEuBiBl1OCfru9Tqwa
PEe/KKqEtOJkdWbICB4qDnJvetS+19IUL91/V/WCqecVr4QK3x5N8YByYf0dk+uW+M998UCNUoxi
Wcv9CM8halBRCAzdrDouND3YnG0R6aiXAhGgghkPms7T0I0o1TjRRF0AxeDyTyk4Egiik9i174H8
J4AU0ZlB0JV+YUUicow0F/zDSFyLjLi5AwqundV5An5TasR3ezREvJwkUO4okMjmdwH+PldNHFtC
KGcbozZTMyu1QEg0goA5R3L4XReDYREK6JTX7By0kbMNQMiEsaWfyFdDQxX1tpnahfqc9EzefpK5
7u7rrsdsIEnTsAV/pa4acIeHsknS8SNgVJyXGYuRydpS4PxKYI+ULHW14Tc9Fr2Kn6wy/Bb0aLiC
ex/bDQA9ui9JkgvavVIbvUgTMJrAuWtUc7fzvpp2R+PSwExkMteITdxNPQyXEEr9lUNC4Ll91WQq
EzMdxMPmNTrr4V3sDxclZB8iPVVynM0kKE6YGcoMTiNNO75koKZn8NBLA+j4X8JBKa9wvKsoNFIS
eN1pp8wL5N+OpVtiwXl9eFplbWxaA/Gv8Zm6XezsUwmMhjF7iSyobGaxs3CRiAu/PvUI/3MdKSF0
mYXlETcw9aDqXdM7iG11ims0vx7T6kZlHCt1+CDo2rpvOgTcuGN/SXUT1XiQu7Fk+PBYXFTphbDC
U2TySQgvq5fGe/C6JLmZC0HOD3kor30SN5AWyPCtChMcQId9S1KYM5vf4KD3y01SS0rgRHbVjJcf
fZgAl6LjvT0Wq0rK3AIOmMT7qHRr9q3Osq1PmHDOBTov5XTKRtf63AlOj2bnVAu/SXbEdecza5xB
xzbbrWE+O1LzKlqat6HZsZ2Wl40oImr9VCdA7lv/okhEJRl1QRenbiYvuQoAmvS5wJ5Egeex2l/9
nag4eeYYIIGOhwpzb51C3AQi1UtURmuKe6hGZw6uu7fkZIyCJj7l+NN4N0MeNrPzSnxX+7ir0jDW
3q0qpRlVtBu9l1Q4KXgwVlAwoWgXXznvvYztmG0drywBjM/3J9KZFsZ50JpzlbEZZll+tTU94MW9
1rvs43rQNTnHF0MAFheFEUQbeZy1F0nWY9Xn4kgr05+Wo4hxl6dY2SEJ+DuJJnOPS+TpWX7n4h/Y
hSxpcrzlIw4Ff7Xmi9L7pigNmKrcUh7n8n1BNY5kpnItO8/xvgNkZuMhphl84b0DyJBNURM8SBMa
oq+COivPyPC2pDinB8srlZQSszr7dtk+QtdBeh1Dk3l8TrtkcyQ3r74K07kA2Lugb3SAnETWZq6c
7a+zr4LhtwQ4fNLHRt8UwYGkgQ82URN96FdiwJSJQ7JEg+NIXaZwELc0APLzj2e1DoEDI574NWXU
F1pbDXr0bAcC0sNJ5shpeVUsWMwo+bWBEnuSNMufi3HvkY7D0j6xM35cOUKfG7MhbcF/tlEifD0B
Fqpe5Wx+qtbfgIGIzfTZTQsf64U1zVaZiNbxWGN24ExzL2V/lbuuMXi0StU7ARVpe40nA0MnOKqm
sVNlJzgeUoD8eriCyiutxC/0e2k9whe4RLjIhU3E9NnCFQYcI5PKNRRIjafp6D8zX2QXaTlnEfg+
WPdTgp/gtIZOlYRP6sAeIgORQPWmSl1tSjl5v0+szlQbhjFUPfa3X8QaRFxjzuStZlhXp2/BQizk
2S8ZXUuwlqNUD/p9S8Wn+md86Woa7Hkkgw4lb32AAK9F10ACBbUlEQYabiB83k3yBWa1TWd8jM6z
ppaFs+XZKGo63b0EwQhy44lFW5Sre9WQ87b4J4LL+OdqqOtVPkVekXbinHewhDJkOij4eaIdckYU
nrrr9nLNJt6MGbogc9M6iNy4ZbTk9Q1QjupTSnnwzmG6T5RrhTkeCnsX1htICW6QVzhC9qcpUP0C
wUlqXH3l8PHDiG37FeqSDFnVwQTinI4R0yAI/N3wIZzqpb0mI0Dq6bdYen/zTkzKDLHM/oXdnE79
Z3YOZ040Fc9qbBjZ65xIGk7eVRO+hIIyOgk+wxQ5cfVozq+MSYr4zLS1dLM50WsNJRgEWJDSshiw
CS2cKCpeFAkQ4e7tauUmcx6+NGTKnvj0cvd6cjr3hR4BG5XP7NBke0Mi9qTTzpn0sYM0QlCS3qyf
aIFukRDKGMDJGsAKxpvAtpRVtkX2XSbaUIk/IKCiqWtZMtZOXjqoYFB+Pi0Zd6rOuuECRcwJqHFI
s2btpehNRgayGQ8IB+nD9jmXkwS+dreNCM/e2+r8S7gYFnTAQl4KcCn9Tdr8SC1+GVa0K5/XHelM
5L60NlJ5qyJlTfLGFcXrHmL+Tb9KB+v4smjWd66MdTpEUNNX8V/3GDTyemn+RE/dk72QEMrZi2la
gSNjpip7OWPx1iX5Jxu1C3St4duMEPLQB5qnpLfvZVanOoL/8elEw9VWhPe5usI8QnHUzl7uNATQ
3EBN6TMbw/EMaKICFUtO9PMGw3MkxqeSLsnyC8WwVk5wii1Qj78VWv4E2klDT6FkIeQq7jWmb1i0
6TB1Wtf8x5SNqC8xQd0xl4NlfXWLcmhf0W4CNe50alTnqeFHYHWZn6fixsIqnVfOB6tvHujr11T5
esEhv68Dag0/iYA3jPXaUY2nQBoUFTe45GS/8rOQkyMeFmL+7KteA6gZw2XBE1eszbmMt7hoTof/
1Pk2yVQj3e6TPuNXKRT9ptbgqqjLGc64EB3d1wvAP2SCr7KCU2u5XUw8Gbb2oGI76kbOq8IEu3ky
fgsjoP9NxeL+1Qofw/GyOLFdVcANPtekEJAnLIPNaoekGaYzu5hdyfwWnnftDK2Vl8wf2UBkFjpe
8MVz2qhWddrcJCu+J+4Rn+5QU6oBWO6NSjQtt0Kem9hsDQBzmUnkgeYbwpSp29EPGSkATrAgR/Fj
cIixNaMM41K6QUYrI5p5ALU9ZCSJWx37Z6/vHgJG+VJYlU3i7tFWSEcGjjof+WHSlv1cYma8Rpmn
pQT7C4vmlpiHmXifsjlx7toGf5W6uPDSQrH+HZffLjl1o2IuGFtb27kwcjrbb9WlzSsaz1ih2BGt
LBejv+6ICeBvqTiYcvZihoKAYddSShjDnQI5lADhf78oZXPaVM9/PIJ1+0t7xW3KWieR5Ted8Kug
23m1E7r0C/nhRhGR/UL6LSgCBZisKu2DW8z45xLGR+hm5jLMi83in4Lapt1qCZ6k57azs2rCNOS5
M10sM0eWIiowvLH6dJYTIK4eEJKPKuhQmSUorUZVIbFdHvgRlz/VNRCysv2EGcyVFtb3Gmha/nTd
Ertj4k39Mi4F7wmzAry1fE5Nc3fGanu68q4mE6srb0pd1iY2Gkax2peuDBWlqQpm437dpw7zHoW9
Q0BzhsGS2OpIYbzUh3/1ObRr3TH8K3XuUhbt8VWr02w+qNc3NsvS/7eZYvOxlFMMLSGdCnf3cbnH
9d0HwXdMgyR4ie5CnddekYcxaiwbpUeuBNc45moN3BsDIfGlhVq2Y7Zz/rhxIMvX4eb2E1h0o6Pb
A7/Jx+IDiuFI3RtJTHtk34dZJTA5UxL+EWYOjDe3bGLG9+TBtGPZsqYeDJKjh4sKeKvvFD8mO51S
Rvvm8BXY3PjS8ssY8KDwyQza/m1lMLHeNw4/Keu14geCm42gm77R0EcgNz/tB1rcH1ELjmJpvvcK
Q7MKKi6iMV017lg+NWxlRUpDOQwHltDBkSI/asZqtk2AZp6b1iuQ9PWuqmm7i1n61Npu8XRdB9Nf
DeayJmDERGGbv75ePnCQkfgDwbwo9ShpY+NFjqy+wvc8jY/G5pPi2OBclBjccfq0PUoLbZbtxrmf
daIIQqnDg8Uug9WsBAuKySGiFUF+gNHWhmg6/Xr9Lx6XDgjk3IjRiGXWbxO4fDB65QOlCLbQsX4H
uqO9cfHucPW+a1KLI3xE1z1VXX+QsEVCmLsT0K+h8g8hHiqPVhrpLLPr87zIBMYpDdmM937Ti6R5
u1vAxTriyT/xqoapBQRiiiN6tdrs5J4o6dJZYNyaw3t0Vv+xPhz2evFfhFX/UKp0DtjSK+AzoLHo
kIQjsbCWor7uoBEEaNb8xNsqX+taHucqCklsFm5fJSnctJH8S0mUVG56E74vlYiAn/HGQsML6fom
TjgXzq1HJiRQ2hjiavEuf62YBQmPjdNpHplI3wfdQKNHy5ZMr5cKpqOaeA5QOxEKYrH0RQUUJcsI
bOX72kK/74V0PJKZnHrkpIDwUeC8J6Mzvia+lzF/IufQ61HkrmeVSRzjVNcYUyGWPRqhcK/sM2k7
28ovC/HjzUeGPQM+dtBj3sJdnC3F1M32kZT03SPJpMnjZMPyco+lg5cB56zt4vwSswv96y70wKAS
bKcYInsOHMzG6WmXbHTNSJy0PB6qJD9r2Mpd2Ooq274T2IlCND0tpzD3dQp4FHac9m81sePhxgxy
bsyI9PFb7dw4EUJY2kn3jCUk5nM50Qv81sg+RPW8yHOquQxSPTNtYoM10kIUFfcKXVK6R32D0Nr3
PiPoPyOOYbOpg04uQDkcX0B7aMW2ymooaTCFVDi/L7Hu+UbTUkCwBXMynl5czsVSKJ4Pw1SrhTEq
rzh8vyxXEF4xwaOxGwYjnmjf6sU/AYQFrT/XEiur2D67rVskcav5RRWfpEGspJIa8KcIH4U0st0Y
7cZnz7p0EUK+VKughV9qvDJPrW8UatPoyy2n6m8htUVj7daZQG8e1Cxr+nYWd9sA3n/WQkF+qIPY
1RwgAcz4sb8Ku2sO7UJRK/qHp9KF4mR2RJJeryf77Tu6zsO/aNOhnriKq8D5FSXM3EjmuDt3vGzV
jY1NC9ww1XM0ga5V3ttNNN/oI0XUFNgVCHMGwd+MpkqEenBFfgPtXOccO435C1HNiDuNa6HPL2II
JZyGvOaoQpOhWvotyNZ8n6ADepZy7kA0eLyLiCA+dJrL6y6Yg2OLsWcHvLYIEszBEzeZ58cQZMxj
6lIYWMiW8hLY5B0P/PzCrqIhq5akIN1Zv57Zlilz/xWS2qLJf8pLX8H0dHCmCWlRvEnops0NhWzk
MlQbPqubXoIgY5wek6k3pdbYmoFwXlzz2cICdMTFAGgv0UIphc/kTxm6C9C0CcQKrY9RDBHLIoz5
cj6DAwLPGtXh7wKynoDVvnmN/W95W+H97PKtk3H5QuoOHwgTk6MGqE0zZi8WGEeJ+kSW6Z2ldhpS
hefVScKbjktakYw4RGBZuYOycnIQAQI/0P6Vo079qNcmbDJjL8n4oyrkX/8iG4sdBkxj/7TAvuZp
oQBhQyLljKnOVRSSzNvraOzab7sCM15cjr5v0PGkVwhnJaCz1D709BPYdy7QdPXsp9QCzU8VgH2t
CGsMlhQV168Ylaq1Vla46YcksbleLJ/5f1Td+lOPeF/bv7wtepOVSbzcgA7xr1v8rQfxy7RgIcfD
ViOL7jeVZGZrXmL964rAhHn4Jpp3YVUmljWAcRpBf9uBCbReYNvwqetBF52c9zXKz8y/j5YWOVpn
dimr+ZB09Bujr0L9pzn4nHL46bDGwUEKwtD1PKNYTeCJj/tlq4vaxrP1yx0CL6jrfh94kPGhjyNB
bUiv+X4b3Pid3ACfEdqdzqcJ+U6WeTrw/hY09e63ljo/8hM4lu5hmyGk2cToaC2z54raXAVLKHz1
W7tEelNYK5myLn2psCKLdn9ZBKlfXXJWIYsYBY2A6q9ib08y3DhG5b3mTM++z+XYcFeHNpzNPCkj
wnLgbGrZS3GlB7qUowynUtNCVAs+mJxaFcwIv91RvBvd3Uj7KNp5838XzcG6k+/GSIu+9LbEjMvc
DgcBD31YEY6UV4ZSHqfFMq/9dgvGRaFGE0MRCmrQ1YbulHbVnWoTNOhAig/DOWThtckrO2FY3qPb
UVcW6idufc9wBm1sf7nRkRDRMF31Bh/Xje5KfnjwE+srOZsy9+js/RBg8p/bfVd2FAWGVCkTV5HD
9lNnYa6ph39xvgvLAC6Nr6aoWgV/ukuO+QDwQNSzumfMC7Q8l/4wS5gqrbIQ1+RM2YU3quZf3YI1
/M162uVgcLjKY9OBZsNmZBSFpGTEOebXh0I0Isxa+rg/je2PIO4m0mqupWohGzADSWDhLGCKBd+/
taTvHyM3DrNbswm5S78Jvi8DJplwtgdDLGBc/l7VKFBTJIXLobJaWpSlfgsPxg45HzQfkW5h58yq
2pyucwAMSD6FFnnYkVP25lGDVUtlnuEoHLNM0F3XuDemJ86wNlnxZ7N8DiWIBZkCLoHbkPUPNKWY
ToPEvaW+JSd+Q0HMNPwIKFivHcNaQJhpCC9Eck/369bqbGmjhvQnTBu3FTGBcEez9Ag7GBGx+Gw7
zzNCkA/ZTd5KmrEiN+3LUCHZaMQjPOiuIT0ApHoM3KrUghg0Hc3OpPTvzhTyq3QPelWRsWmThYS5
GSIaLxLyF24to7JfxzD98sV9Z13LO8l29OEVCrfcOqseCkkbWepi9vC781bkqQm/wCLlDn0GoNAj
LTJtUh6wb78Bfk17bs1Fgyw9c8G823BjA0xWxnZubDEHbdj7GSqGUL0Vut2WcnfqEQUJbVJSGhiJ
BMkRmV/gId1DBzZN6EU1HvfPoj9zvHg5tGL7nTeAYnq9CuK/WjBcTCUJU6YXBplRdhIEoqJJRl4V
CeCnapH7MxAbkpKMaF43vk9hDU25uPCpMUo+wXvjw3u11WLpZsnkc9tT8VLDSXKlcidRgD40TCy1
UVeBbfcv+Ls1oTwi0avEQ+nWjQCFjqMh5arXbcj1dlPSZAGwQb18iO+Dv/roSJAep2FJsJtAVLIh
qso/9ZPGDQYpMXVllh640jmjcsX/xcsl0mlK6yP4P7jHWDtppIj7XnFABdfLeQQmHeIjKK3rgTiy
eXAPNnDoDaeLZBKTY4sSlElQGVkc5GDnjAHwb/2tUZm8hyVJjULU/QOQpxVP+Q9E7R1AgRZI803i
i1rC9eKztb8fvebOC56p+n0FZ7LcYeNM1rJ7SvzAIYdxETb9hyarxQzk0uX+Rq8DIgmiqaqSr7NG
d4Aycsuo3yPetVBHI5TLmYm2xCi2iAh17l8I/tM2AfPRl1Grz4a4J3AHzm1trY+NGzZsxzKDo4tO
1mGam2oh880HfH5MfvzJjzvsY96kkcyhFstdt8EAcb1ULSiwFQRNaDT7QdA5PrlTW07od4RvorBp
EAqrGeCzJs/2xR2iErRJPXy5yZuTBOFKcHoYhq84t5k9pIJfZwm2AJKO5W1V5T/kjIVzBweBtP/9
eJ4ThdfFIzvNlUDpMH+9abCBvg499ZQHWGNnbPyBfVpY3e9TaZYgV/YV16wJYV38ebVAkAkP7Z4t
mmpFtrPeACPiwLLSX9EeewqjIg+RqLsCLFaRN3HOrWQwqNfgd7OzWkXfBUPm0gGmQletSaBgt0GV
wmWdNWkR+O7Shaqj9x9cFvIHHLKA7ng3b+zJxDUjHgkr2ckQ7v39vycIxL3CzQq77UWEUoPpK1ix
/6N9d97abmA6dJW0QBxOhyZHcjS2KArnGDE3vzoYJx2rHvwTUrOVkLWELkqG68qhuGu2RgKyaLkc
JCIEvdza8We8Y7536kh/+xLOV0IYkoNg63XimG4poA9WPcdVbW5bWJVdEMw70nvN8eEZhYk/VB0R
6AWalb8dURM7OgLpsMnFtlO6JLN2s6mCeUxajD6gDz8L8bh7rZqg/Dhm39cvc5KB9XmZ29dY8c9R
qCVlxTWvDrBZb5xLBkZ+Tf9M3eGdx+gTp/ocAqdpJPRegJpR/xLg+h/5ZTr4+NVAgA1NLB1AwKtG
KKvr5NgkSaefUyVHZi//et8J/ikUjzLJsnzpphnluP0E9fA1s0dqZh46qfIVwy9m7mT2qp5T3wwt
rF6ezQJogGWnFH4szxrkz9ydIxRdP6T1fJdJX3RgcvcbEzQ1fwwPiNk22BopHROMgw5rip8KkzEZ
K5XO/28893a1zRFVS+W8MPy+X6g1HWXEZ3M9aqwiZkQELwa4/eG9xeZe8X/d1TS9nwobgXaop4Lq
gJYJ3olFbJm+Zv8+2x5IOtPf1tI/DKWja6fy57yMiBhT4YIn6kAq9yYDshHvpm1O+DV/7PGJKm93
NlS//deIY2UzvDt3jQD+oghNCka4Rr4L/R5ZpculyQ1JHFz7JPv4xv7u1XNPRcUQqOIytl1OWapb
1Fm8kUh9zFghLzfv/PybLaCP9hnDiz3AKOgsJccd4aRzRdDhtzJ1CiFqq0nbXhwpkaqSe4jRPXES
5d2VbjgXDAUeEjwpVEW2gJTATfJQPswLuJNyI5Wm203Jm9U+geMmleNUGqD/DqECiHimSIMcqlKY
mC//+sT/dXgu4zMBqgQZvZ2QX5nAzuF8iCyfvuuGkJrKDzfmOowQ+IcqC/7JEZI5wFojDYIB8SFn
Yosvab5+i9rS+9WvMm0F+fHrisnYX/jKEuTuqheGrK3u8FDgLuwJkspGkhNxWTH2KpXTlvsuCd7G
2qsmCIUTi8m8LTKUZjCzcFr0XUnmncQ6wN0V2mVv8TkVomXXfPUa68OlIFUbEtZjsQ5TpKiELprh
sJ3zgdMaukmHzaH57RpGCbX+sqzMtZ4T2fgVw1kEFFhGvN6PA7giJXA82EnCslDT6Ml/OxqGU0tV
MOMPN5YAQId5EgD1GmJ4rtR09cH8T8Lm0YBvsLPv2BU1VFJSPIqAZZVggLkBUeBa6GRLf1cKh/AK
ASZOWaMjCcYMacmGW7hbz+/dzOI7zdyPcLOZeq4EY/enKYKRGeXIhhi5PbIHsUP9SdbdDE1sxKnb
xV74hTLSdHp1hNqjK27ID81GZhcUfgv8VZ+JV5n55RhDZ7gsXsFe9yj4wGc0ELbF/CL7285zUMq7
U88FkN4k6wAsMlujA1QnNcneNytn0MiQB2g7yL/+3pXluh9u1RKfFwCu1tSRlbNTllJHaJc0PZrc
rD7Tn1J80vAI6vtT5lz5eCQul5Sh/QZlltRTQSMDpoj1bCvDHYJ9xORiBBzseJV7gruq+2W0tv4K
YNuq/idLGxPwOgcv/gpqPlII7UfRmApLxucUdoiZbnjiBrZVh+UH0b6n6GqD2LpeYpba64DNElLM
HY9zPtfkuUE3Kw+4UqvAhEACvKHCvoqAeoxBAoZG5gf1PthnY/rSxMRGVoyzh77oIlut3E1bOPSO
sc9nNm1voV8bERnEcOoAaVezoziVkjg6nmueVpyeqEz0Mpc5Srl9+375+zsvnJ9WTYrFWhDmiIWk
oWDeP8eTNqqHgj+YFuZTqTy4IZt6MTHwwCHOvjz6I/+rwj6X5jg58okC6rR+aVPB8p5Da/pFPX4s
nQEVRhHjP3tjMpdCmVMZoj4/GDklpVJNbhkHgZYQTit2mIzD0lIxZyJOt2DCsjRhjen5kDDdQstY
73a6r/MeUxZSjKXocOPUTXS4yxTua+2u+eAhdBxpw14e47ksNUFFKfUCRwNHQG+M0Fek4D1riln1
Ng/WnsU5BhDFx6162kMsM9I9P4G7xjDbkdrrQizCnisxJXcLDoCEa14jlccmgcKpXlqkPbzQv92Y
IS5Dw3pT+LUOP9+1sj7+XBouQWGv6zxc0SgHATPe+xI3z+KYzxXoaFgEm4KxF5O5E5jaaf5Yqny6
c9+7fy7Ve0LwTktO/P1wPNvx4kFIvseWeiMkHZx7c6hmzZENGylBpKrfFav01741uTX+hXZmqqnX
GzU7zdW9okFFBikh5mv0etADk56ju+vWYtKaekGlTrqXPqrM7r+SoOjIuC2Mv0Rf5XLLQUkpQtjX
WvVMx6/ms8e9gQHBtk7tUiSlcR67uP+ereVZ073i5aNfXoWUglT9aoG3T+UWeTzUJb6GLumtte51
efJntd060ur9ixtSl6GnDFqTrZrkvmANbgQvfew0VlKv4QQGN+FkA/UXu7sgw5gzyAIu5INji+Jz
hwYgoTh6ASFsjUKQb7qsadbwbGhS6Ln1MUHJxUfF8Og3n9bu/8+dWP10D19nZIvsgPGttzFFH4Vb
FmgUTpND2QE0+PSNOTIvbzpUafhwhcR50pZ0VaqNgXEMTjsHm09RbjMtlSnrUtmBfzt+Zypu4bTF
l/WPfFfVWWu8pW6Ht2lsC90aXmnMSWsuOc12aKrsiSdKwBsjf5OwmfXclIKA1q+WA0DTkanh2cVD
yyEmxSn+njKHwEB60eKEhP2djSUBXGjrqDg3+8xhYcT252ijGbH3Hz1SAL3hvkgc93u/H1Bd39Jt
ccbgLn8cCp6JdM7pvfiOSQDahuWeJ+LH6rnrLtRkh714LzHlcmlXF0/SwYKb3oBpBZjMaG46eoim
04aokjU2F5+57uk3kInGbwwoa6ZfKLFMf3oImmuxauEF2eYGhyhsEhRlp3rXAIqRgP/80Lu9Teq7
AzjItax3YCtVdRkSWRPcU/20RlevI9oZIxRV69EWYlifZb7FXj4IQTQnwc/nuXFx/nip74BLXSeG
FVu8Su2qhBmXsFNCUNKFxsXcWUA8othdcsru0dXFerGhmmql6q53cuH/Xuwx3f+jVwjeaMxtKYn5
gotK3kKt8ta1zXRjCpJf7vnD4PAdumAwvsyXKPR2tNkw3wsysAX16Wf1KhAy0C9udcbtEJryGvzE
axrtqE6XuqMG3FegZAvIJwi8SMbX1Ci7fzwEN9n4kTs1Qkz5kaaDFRYyKLAlCykLcJ9H/juDwRwv
w1uQlVPbD2vxgBQpLXyMJKAsiA+z2ZHiJ9/UKZsPmVK906/13ekbTItfZviim1HzBNeeUGHn1uq4
yeET5fGOb6yHXeweHYKB+Ah3K4aBqdDZ96GQgJ+vrwZwTjMwJUguC6FRi6mVnXexM2XRZ3Zg0JmZ
p+jgOtHOrFc+skm7uld02vi1ITtDfn3S7eBA0NaGXdhnBxgbT8z35MV75KuepybmcZ9X8fj9+tU4
ATe/C08aZpy6JaatlbZD5IGqEiltXgjeU+AebmWRft0IMqvAAXZ40VfrOO9gMQhLuRmgMGTCiOxQ
oV/KixfFg+UeWVng277Po7giRII7qBM/hPe/Zx91oSC0KY/UOQyj1RM0sKXoIrR1VmoqMmQaGRCb
hyavRIBZ5GZhl7q+oRAbj6Jg2KlobFHhYZ8/L71+exQ5+HuwaWrJSyWrCukRbh3WYQik7L3V8TN0
48iHW11xDvNer5HTTMacn0RyZRGzq3rATx+aSFGnlMKqy08ZE/eRyeumTUgKjmYhqabZg8TFpsmE
re1DVnf5MbBVEXZxezWHt5ONXeIpRnPpbZZ99WiE6kIi+jwb/GVYO7quWRP+Vk+L2HPfHGnZPLnc
FVfTnhPWIy0zp7sdgt7gwSo3xD8ShTaDlepSUOXTGKL494G6k2TfKLdBDwM6FSWrSKHS/nZiMCGA
JUvXFC8yvB09N0jdwqaEUsZDYAktL2dMuNvuYecg5LqsEB0a1g6N1SyiYRB6VgGWXafF5ZgtGPtH
7wgdcZCRCkopsq/eCXr0zLcFCxaJmYi6L/y4JnKHQ7pjk0BWADCwStNmZggzbcMpCxr5Wr8UV282
OEhTPqVerkCLXP2LG85YvTk8nRk8QFVjVgsHvdChbLgy85vXqtRAVuAvafUmQLJljxKVWrXpMGUR
AwdbtnL1eqmCKPcbzLPTjnVwcBuztW3BOxfxOpCgT8HlY2AlAOG3QYfIj+Fh9mjKfSMhsczMaA3t
T79IGGAa/xMlKxfIk6rop8dl1yVpE+PlwplnqAmX8etVgPA8iSRqcdpn4YWK9/yjZkQ5f9cM0QRp
IQBlMmUeuMw4UN4+IbF+0uTpmbDphopH0wSr5iV85nQvA3XnhfK7CzNyarVKW2E+dd93ZSRLTXxf
hFFdt6nWEzYmTIsicHagsgpPP7/5UbHwOvQeuIyxjrwKMHFeXNdR/rG2WD7GjSRprsF/BHOOcHeJ
UjcZP8BmKXrfK7rNMXX0wIu+P+qb7jJItIVOLnsDhkC9f/fbh2JKlwkH/RU9H0JnRftssdlx9usG
NoGHAd07si++Hvlnlgy8nQVcWAJ1lW20eN200JSfyQUJDWuwuaTGzqVnyAga53Obw7x6zyThMvcS
qNyfK1r06ceQNrYEvVirzFPquaelEYUaiq21qYOH7p5XLpTeBdHxah0VhV0Dao5n4HjjXV98lenn
Ka0hQOt5RUpjA1PDu9oE8JaKG8zZZHExPwP7nQjJBFD/3gqyfG80biHN0CS82nM6aOIJfEovad0R
Y0H4wqgWTQSGcx8dVsrmHrWXeRh8WFOpou/YtjsZQTiJN68avWrfPcYtNsaxvJ85bO54qCPVAWaO
sDZmYgbi0R4Um2wSpViQ+hNRsFMXnQsI5yOtShB6SJSVE2HU6n5OFHE9EaHwuPHnOg91IcJikrp3
52AXgBaeD/Bt4KJLVTaRSICIZS8d6t1ag1F2CIjadhbqH441BcKXqAPnDOTvLEuIw3UhwgyA45aF
VfqIObavcBWJ8B5dcAUzn8Nt722tWgoHMrVRPaOuH0lhCCmjPHrnJzRPShRJMimiSF+OcJFgCQ9x
NRQSACgYEJxRuqqDtI/PVPQOM5BmJPdM0GGyfcnyIMUKMKrb/JiM5deh2jmk8KuAmXkyfnlu7D9P
Ank3IrQoJaxDlfPnyYDEk3i/c6ks4TuaqrRqU7DIpkUzZLv6FpDfm8+OGAjGkNPSSUE+Xdo9OGIB
YasMmmXea2Kk7q4MLD+m9ziBuQqpli4btNDwdV8qEHNFZv4s7G3Pp1mPmkYkxbFZFyXSXwS/J6YR
reJ5X0opQR/uFE5qTxsoaGt+hmBnXB3L2zmxs1/2LVw/tIa2qdJF3t41S7ca90Q5k7On+xrbmk5A
bEsUzxn21DsBlYHalEoTDEuvCKBuCcneXem2oy63zor2uRJX09ZQUPp1+p4NlsIp8635f11eiewW
V3ePjPY3aLfPix7P+iN/ydzNnMVdsqTEOM6iMTw0qOERcF2xLQ2XZWrBuR29GmvZ4n3S9GXGKgK1
W8c6GIaIiRoQzAATf8rttgE8PjCtQnhS565EiQ7dIoAu07TaDLo8HK0+H0iSQug8SYxo3/Jx5Kx7
kJNOqPshny8Ms6K57A1Yn9acFMJfU6AQdGjMM7X2rm5HbTLKhRX3pcVLQlRFRe/18qtx7SN0iWQ2
PG76VTHI+WhjxW1HeIAN6EddCaHdDfeHdKLYuhxm6ysHYl3sO9zC8KJc3J3t1S1INArQ5rUDJAwz
oJ3NPtvSJmQ+zUIBIGmz7PHTSNoEcO4ZcrwVyz+H0HkpduzE099FQwdgxIRFZsASyIrvcFU+reFg
1QyixSrY6XiMM39TiuELZjvKJf0dRNwliH57C+HRm0lRloTUyUv/UquJeJMrgGoNNtOhWk8tTZCc
wDvdqfBALPcjN2FymypVY3IJu/GZE3IFCo5eM+G8WrrKUi5vXdEu+BhiPO3UjT4gA7i5pAMK/1ab
eavToCpokj+oYXbc2Tt1UX+RB7JMl6G+BNnGE+Yij8CijuxM5OwjU+2pk8OVR/fVgiJKj+Dso4Di
svi0OGh3ihoMfdObp6lZ3C739y80KYBjWZdh8yizVuGk9cpUbxHIaiVmhsxHh9dI+7UWxdCR0wJs
ZPl6oHzCi7oLrb7XG91OprTA9DLUOPnGi//VvxLbS4vaOMTnTKtr7bgA6qj1IWI6Ku3zikjjmEhG
kKDZhXv7LmjqqCQiJvN80bEjVRXq5bZa5WsWYB75iXLmFuPa/4LjZbvCGlRVGkMImxb6Tfw+eKHY
9YyghA8WITLzR/BP53AJm7J/7w/67Sm2Miznt7Abf7M0evbRFrkx0lCbKFHPipOuvqfUrBIbbv9L
RWJzlq63Iz2U4SEYasNa3ZDbUSVAcTKpUyI4L0tByPnaNfsCuiGk0S2s4t++ICLpXhIyy5I8giqc
Ky9cjZ7fJkNXmLGfEIA9u39ZEhh4nGPAqUpZqaTkcAaJo8cwG7X2e2ZQXnJzp6AQlz9DwZvO/N7t
a7GXBibq0pplP4+LdxRyvXjMUm54KXnQYwvXlB6zq0A30W/Jip9lgRLjMkHZ6USN7rc7tUrVMMgk
tLoK7AWq6Uk91pUK76P+tTIbQgVZ3BeYjFEQ2hkkfM1BQecLm+WwKGdRlou7mMcuso4aGi2h09S1
SRhskJ/5mXWN0Zir5PPDkY48QXllJor5HPIFXg4aSzcKlb4mIUCC4Q8aSXjlWQBQmA7Me7eSmrN6
FnSR0BvzNBVVbTSjLf/DrNJWSONzbKf4Fr65CKUBvYMLWybwwvDChjc81/2wvnJ4PhnPC4ZFYsfe
740q23lK0ytGE+s4CkBSR3pOVxg6lGIuEqgoUnoIOOPvRQQbHwcQ6P5+qX18h6++vmnIcMiJJ8Gn
aDxHODFBYa+oc4LLQXKOARB/g0Al+XAp1qwa4UBpIGGSpYThYByeKKa810CSlZzgTHtrw24YFn0s
4xr6zA5fZUDitXn09eAXvHT7AhiwY3Pjab/Y8CHszbpQLw7RYo+lXI6LhRdpLAIPgRbetYhIsxJ/
utpDImBPPAVXSWKgTPF2PRrcQvUutEu0ixzFV/Miiu4edt8iHRY/caQTB3CtptlIofyA/dxz0qhf
CVCKZGqhXxlwBmyyUY4vrWQlMfQZ3zo7S+bNJLccTU8ZGlpPC3pnsc9JmN4HbJk5KmY3fKCfUbzq
gM7v3HL0LtCcrvd0JmOstz23Es5qwN8rtH/fZMeZ5BY/2mrjjsw8HWb57KacL6zRiYszeV4SrL/h
68sccY4zkpvobemkRg037AfmVbkAQ1kTfU0cG4j830FKv59Gb61aRmmMKQNV/HJM/MmtG6k2o4bn
MGVOUSsiDb0fv22XmFk7ks8z4LuuMSaPQv/AVkCq4Mq0EqHUe5GBhk8bvFJ+D+kyL900T2mOvN7e
zOcVcrQXefyrpucDbur+TJfsUhNkvvRBd4yK/AIsJtGBmpfjmVwXQPBKChzaKfpFyC5Jd4q4eIx8
hcmIsayVApmdp6ea3RJRpf5EzxfjAUlAvCISbtuFWs5mS9RAAshdnV0CJR8JhV1mZLERl6e8ybtc
ki835McdxfTecE9Y67nfe/FAn3XpskZZzO+PJTf3uV3AoUyJppvkeUfwsOpHAhLWDXhEhZdq3i6t
YQRfikveu3skXZXjs9YC/CD61lIIVr3xGRFl/137ud/sw1OGmv1m5ldcscSyladtWUbQQE9IA205
8nvTcIKZEixu6HngSK5UTl3YkFxd+1JYKdoAafTc5UatbovhNjwRHxv47SVJyUw5Fz48nlHIWzlJ
dT8DKmSJAYzPDPrRQnjXWL/iqX36yMYNv2ZbJRk1+swX4oR0C0pwyr5rBg6llj/no/+QLP+ylLJx
XxA/wjyLsdZZz38UDaQ4NAblxxQ0qFucII5SGNsC9Hp7UgqgABnS2s+y9vyCPyNuMeefQ9koKVT0
u9WWJ3LpiU+GSmCsFMsQ9bloutAH2l3HDGGSVi8LQ+szKrQCpSw20DmUWEL4or5PkcqXD8MJVK2z
9iwGDix5uWpx4DhIQt7O8+IEnkbib8/O/AXwJnzxlKjsXy91vsi3hWcyO2J89sMJMBan+L9yxHww
YDrawdp5rQrWlzWN274H1qNsEIXSsmSbkrfwVJeHhTriMQ/GB+WXdrsfQzowHkFP7yzbSmPUIKB/
skhZPSEQvcazum0m3eMyEXcA4YR6x9USaktC/ay+14SGhIzduO2lDs5jLbiszL9FcGKpjVFZseDC
u9cWkbEZ1eYMaGmdkiGnF1JaGKZg1YxsIBCx00hUUg8apW2iH3uZv1RZKff8nGsH8Yv5Aef+S7lw
Sxn9azu6YezXFpg+9s78a4euLrpQM7Q42J7sAtjrSHEgqEcBr+PNyw1/iA4Kai+ynVzRToi3N0Jj
gB9iRcPpBQte8tDSgkeCAjAf/bjllPAhFu7GMX1pJ2ClXNIHCTppcAUPSEiC5xG4jINxDQEVK6Jm
y33ulnexBwL0ZnHR6aAywqYBK1cIulQYgghS8oUlB1Va0SS7jJW6tNwVdhUI2Px6OfrxbMGmcllt
uo7yCx2tC7cqagOKiIHBM54FMSuZdjat+qt1sRxFB9G++WSIQCsNAujBVDk3GyqD9HFlEpl0YqYd
SjcdV+ebuUxDWfV02uq49qvhitvwgzlsA2zQ1hWBjrz1QUz1qvfqSmwoGqactDDui02bR6mHPL2t
Z/bSPUC7uz44E0GO3+S+hn3a6Yyw0CDzEI3NjYeKQeI8REnkxC78Z5TnDE8Cjb0eCstgzcWaTV+u
bcYRPjJZH/v48YdYH7aKkC5jlWSIyMRuk8Cthj93585H4tdHEOY3A/QdObABzxyFZGM1LTgcInwV
axVFLOqskBMjy/QNhk5JxNP89fdauQAbBqX4ex8uijL/L8mfld2A8leOs2VNJDGa3hKENiCyGZ0h
p6ZYGQc2AftMC8ABW+oBfl8EXdghpTwd/L607XHPxVH1tSrkUsktfdsks928zsDkOLf1xqcPecIV
Jy6WFuf0UI0oxKyujkUctOvaXJv62B6SmNU2+BEmQCS8mtYxxhYU6NewW1hAnJmnhsIRI0HJO9kq
aR54mZuj1VoC05Bh9Xh+jWmLoTkwo3AbdpfzILNFf3NzdvN36Ku9EsuJu9waUmHiRXN/QM7BpnIi
J1ZeNA75JwCzkhQantb2hejGzTE2FIn+DN9f6E3fFO6HTgZ/tdLtRvQLbVxPALFb2NSQAZzh2aHE
NNKRUr81CtEbpgijPjIy7y1i32KXhapTpXK+4eH/OHHliU/QESzcNOcvxpKqF7pdLbf0xic7pXJN
K8DbtJUirYvw6dneuO4h1p7K7J57aKHgewJ/PKzNxoe8RRfsCeqsjwradpc2KyTpmLtQqNwB4ncA
Ip7jpq/bb3yvvx+JPo+qJIbLAfKFkgjmBnAaSaKzcXNKC5EnfKhBiekaWhhuf1MLxZxZQiF9wL/1
x8ZDc5zJ5ZZMU/KqYKJ/64e4JlDGb2ifkPxcw3ZDW9TNdlG+8yvcwBarNTk2D0XuGOaduUjNDfOO
bmpf6c3h6RuwYTnLU4wTd8mj+z0zfg/u3tyyaowg4f+RVYJL6PDoqSY4fU05MNIHPS9OYzqXZbYA
/zzkBCsgu6Y/3tHsKBIVIspNJIn/VgAnZNKwQEVLKP4VQFUQV/zznGkK4UWQTUz403bpF1M+Mewl
J+9ao8Mo+bNN5A5YHJkuJGed17zGrphMKREY1EqJs82rkb1bKosc0R8t5ZDbwl4rtJ6k6D+uvWx+
D/hkfrasr+BDCbtW1JOtQGyQ03KhcArNCsWvwV2hJ30RkK5vDJ22YLYGFsgyuqz7Es+H4c6OUZoE
dqlj8C1cKhdRvzz4ZC9y+lcE5mDJaKFxwNFNuMO5afjxj5z5BDeS3bTL8siYNdogdSTw0fP8Jdh3
KxZO3+EOZV8LWVntmFAfvp9H8TrZp9Y20zTKjW5z5zqL3NFA3cTYd/vbhw/0W2YJrW4cDjJscpZO
3YGscn8yzPUrrGkJcxlqOFgtYUd9b4wU8nTjDMpi20cTGAausky4AZKKd0TGfawfShwRCHXDkUVt
QlLXClbOFGKrFWlwZhenIJfqvPU/y/brSObGK8caLV5gvoYAPq6VtwHb8tIXJKwt2tSEnUP2/v72
jV/eomNjwvTLkxAo8VGC+sKN7NiZ7fo4T5zY0PdQLv6uTIwkoCcTR1IFj33rVOUQMGqcN3JyKmp4
Grh8lvjAJ9OGl8wCfhxSc3Pdcql7OmKvsA1+n+e8w0jdS4GZ656wNIJ6EhQe2TpWoF+SfYpUJNDh
hm53Fwqvb9VkLlO/BJH05/qmOyjX55Se0UM7ZlRjd0G2qI8RLKm2eDld1uKfEXrCqiRgxTKwIsQ2
6wXlD7SVSiL0qhiUTlmaUWWMnV8rE/ZTlPxxOLYErueRunoumNmlhbdq4bGB31M7If7UdIQcvMpl
wMfsEaJqXv31e/YKlSSGnqfDs6TYGPh728GTPHbZRfayMZTjYg3hZ2GFJ/yg+fao20fH7ITHFfp0
g19kTe9i8z1uuNRghx6hNaxeIYrRm0cLw5+pCEYT884OvxEXNglL7Cj4gYEkb5nKKaDzzowhaE+P
9VEV+TJDM6z7B88DjaOdujnURfE5B1EsHWBzaOOVrUqkLa5JpXmywdpS87F0xU0tuMG+WBtWmyn3
07RW2QGdPFO/9J8IprVbWi1uU2dl/lJch2SybNuFhxnZQeErsUzMGg57PDyug5qHwUlN1dGKGqyk
jpnY9ClfqTYdLDxjf9EqCNEhGbpoQ/bFYJ6zJ6B78EAR6yKOH6oOSrdfvyFAqxDq0ZKVGu3syfS+
OWFpWMaBYbnvV6B+epTAvGYBIkyB7QUmjB7wfwFxiF+29LVbxn7GTRkwsmyceODQe//FQBMKNPOD
c9K0eRt7bBE0qsX9x6pPatHqabZj4Xal2FkiQuYeKb4ASFfW+r1m1N+HvsYlSnb8Ilb9kF7DKxkd
Nvpo+UW4PL/alVDXd3fFj8Ke/iuWVi7HHmOLW+jBh2jD16A2Vu1R7ZC96WnHZp+TWAByxCGsFfJR
/6azi8Z3FPGkJPRCjjDEkrYkp5beYDqxewlvLTQJoQ1qClF+KwuniVSaSuwhgmq8PqunqmDquC3A
CkWbYpniKOZn4fk8xadrCCHTrtrvXpwOpFml38CTX4dBI+O900TXcVEv6d5xgOkXaHcc0rBMFJWI
cH6J9SSCO/Hj7pnxLUcfusmzwj9yX/FCd9sAOsRfcTjF4k9TiapFUDyMk+NJV24WJwzm9WxHBT6q
0fhem+1uMn08fKPH0nGlW/0pSpFbxBRTTF7A85B5Jz4MJ+yB2DcK3lqPB7pVtlZQVGo+amWkjD14
PXzw8yOIp9P46isQ0tqXxb5krnbybv1BburJkOfpL151jxi3ZjWP1dVijpUqN39SscJSC18zoOGf
Fy6svxhPAcmCvbui6qYd0pPPDrHW3WRgtWN6AmVE2PmyASth+wEQf9BIrLUIBEO6XWdBdjbtE9Ag
25BATTL01FmidulvWWP5jwv9FDeW0wxTDmqdOgP3N37i27dbiOkeG8foOjZu9Cvj7fRu02n7WMMD
Co5fl2aU8k5abJpCmxCd7MHVdcKNNJQ1UFUcCXwscf5zGkOxyVZnm4/jGSIbYmwFaFLMIg2sAK2G
muJYzZDQmPHnjMS8s9evXkHU7/HMdyRIfEKK56oJZbLNVJ/dgxolSzJaYR0ZgxOCY51h9nmJ9S1y
ZsX7+5abfe5tObzCngqR2C5zfI2fHCP6C77cg/uCl2JHPbA1f07aRE1tLBxzwBFIegXTl80PMMkJ
j8/5fjv74kjkvoj/Iumesbh4dq3GOKLwiH+vC+kvO2K/hiNpS3qthbMW6m9S8kEro1VAvkb5frAw
yrQjQWDKMk66nT83Rp6wFADUFjNfiMDrH6HV1nEBueZCLBVSdXGgTrZ3KtiWc9sR8/6moZK17fFm
TRT1kehL3tBnMex544KnYDvWWn4rPu++WSh6zbQRMcqnld6JbGYsaixYz5h9F2saLgKUdLAmdqww
HHVAGlGdryN54SJwbt4Z93zX7UIuv3CkTcuoGAiRjTCN7XtDKQ+PfXFI1Xb1tmHbCpJce7tgkymj
NZ8mVLyjnbvIu6YXao9BKnOxriprHDaPoaQ9kTWPeWPi5y633NWf6fNyfRo+FV+C3SpmBhE/d63I
aFctMc5zhNyCI6JshO1nz8ooo19xwPoRFap/8y+Z+Mo6q0unxdaYVIwL13FmsVPPibvVK2f5uEjV
sU7BF76yDYumq145rqoWYZqtGgAvWWnY2YRJFqV11ORXFQSYrf74/x1agxE/EVFNWlb3zhR955d0
M5L51/6Hc2kcbESivOuq69nYfBmx51RywJtXdV2e+ejArBbuBqVTk28pKtpaqDiY6PM07h6wkJ8f
VmaMzIZlJFb0EyGo0lLukj9KbFw1bdDF7lbHdc6E9P8e6UgdukrBUfOtiA+bB0TN4aIt34paEIma
oeb5agkhKzYfXDTOPqYabVjbz54RPH3aI8f9CRW7xIwDa4fyQp4umaE3btCFp/hO8xicRrgx3+hE
Jmc6UuiVwCNU3a44xXxR5y38FK1a7d3uzxMBNajP96fA4ANNq3BWrNi9yO/0PXM1ohcaEGGz8XyG
Xm9+n9Ar94mB2nR+4o1ddATjh+LY7IRlmJ6ualuDeRLvDExc34nupttFNbvhyy7X5BQKU/CEZL2V
nPK5eHAlRluwT3mMq+9yYNDzmCCwBJKnwMW8b24jO0uQG2VE9DLFmWoBeeKdQ1bzOlNIJ8aQRdkh
Lk5I3kzG7AP8lA9oQeIJVWUYQNp12qVSax9MyF036EnmIxTPkDNQJ6A1T2pcxIv/j81aHzHE+Mg8
NRSiUuo81EnfrwXm8JnHQ3A8cO+IlpMr+X/0fkmhqSDWv3Y0iTn2S6Yk2OJ0kH9Fj1LObuOYK4MW
C+fuFrAVJd2+/ylFDt6yv08lp/GL753mNgCCCr9GF2N3WXjzqgR5M8ASbdHT+zv5mcBqzpQ4hwgm
xkYSKiUqtkQ3Lmy6tlekNJCBK7/7TYO16DdPEWRcV9hQmEnqQ+R6gNMhHQ6d0LaSg+jlYDUM2Dai
XbdYGOVM4XzcquR3x0bhJBdDnn8/nsACPXalrk8MyF+T/A2+gooW5iliMnOZpOVShx23CEKd8LR8
isVh/K6fubEGjf7r0Zd6Vt1tlk33/lRPyX03E1FbmNSwLs7TW+jjaEJfWjfw6i1krp0qCYsi17MY
MDxyfCVTgOMGRJW8IlFI7eqZ9KYg3UUhm9645+MxhvTyDgUxZ9x16rxBTr0qZr6PJAhFZaCrvbmO
l6WKdhpFjjNAQJfvVISNmrRouGRCoUWm6paJZhqCH7/Ys+Wf5xg+Sc5hURTH6NCQjLIWWk9fygkk
hYhDYkYSursqhI1wdPe2KYFl0kUKBAaJgzED0+TQdE6NwWs+Wnv19gOLUhUkp0EiN+O5tKTO4owB
lb+rTZ3Hlw3ZgkQFBO5Zp5HFqipcTkIg7QlhJO365EPfKCCr53MF3fHOZa7KVX7NSj57DE393w5e
SISmDD2kpfBCH0j7NES3Tjl+iDB/tp2Q4hvFjIqaN62QA2S/KI1dTTdPo3CDwypWL4pBYb5I/q0v
lyR2MdQTiIXlOR4ifhJYSM8giPEyYMcKGK9FCx4DgvFRni0Ow8guzDBXdfn2QLkQ/ut/WvS+xaDV
MyTIO0A/S+8VlJyIEYU2SGZcMVomLj09tqpAHJcu+PkCrvnaPqm8uu4njb3JV6Fe9fpcMr9ziEHN
hBpxsV/yQFCtGnKVxtZ58Ln9JzRzST5AwigqOOvGQwdBrLrlkc1OhhOjOJinz9HwqcRhgn0OH4W7
TrPwf8Zwe83KUueuUGn/bGZ8Sf7bSXVF9INhJmFi11cnhHPQvtZvqbNCDaceRX0S1dfOS9P50FP8
bJQQFhmPOve7R5a0tR2WjlDE3hq0ThcdId/CjYeYjGIZxV4TCiOUJwpCT3ueUN97c89YRL9J+GlL
KDSMcwThwvHc069ynfEk3mZDnZYCBo8BjzQRdcpX+wyF6walq1RbJ/Dr16Re3VHXlCTGP2J/6g5B
u34bJxi+GOqrnFgbZ2t4s6+UjByTlNRKcAdwFKnmX8C+yDw71S/0AKopLfIG52a6hTCgulGdCiSB
apLTwVZEUHIY1v2Xc4O21+6UpLSgr9QeN7vOXPyMYg/LeKtZLkXr1LsykmRhx+FxoyDrkTxld7z+
ONCpk5k1jHHc0YkivsEFk2rSVrV8qsE8kQT8AAs5OTZT5wPXI3+wUBxu97JKKCAOwLgq+1nl5hgc
CToBaUrG4cU3kxc5cKkvzgLHX6B5zsKsRbCtSI2brDLmRVZcYk5g9xnu23e/GocCc54BMG+Sek2v
sxN5NTsb7Xx1OPIeu4t/vRTEpX3ayOsvZ3TzrSFM/OawGwNvuV5IjBmDP5NT0fYD9umVsNrByoDd
sqs1kPyxVc9zLdv8E/rqrZ8CvjrMUsVqXp+i2LRNeEsFz6UGa0lqQxFhnJbMT5pPIi/OQgsC6rt2
V33u4ZLEAcwTxp5ZYWl9xHmGbyn7nMsilxbG1OtyHe7kX7YuiqGAibJSadyE0IM8JK32WQYfAbtT
fyVtEgdG/It/lEPR6cVPFJMLohZFMmz3LS1TXKC00wKOIbGbTE5rSfZL1iyt0s9ImEP0Zhsrk5vG
LHB+kplnmot2Y5Ajvimi1hFYQWQuBR/u9CjPuxe0L+WgtYdbv70ZORkwDz4IREGAvDnp57dBjGwn
fypAyzfCqxm2prJ+/hIyGODHxSvV7hjpO4Eo00Rr4oKxwZvWNOs5y5PapEVShoh7mUQbGAmPlYHf
rX2AenyM3KlKWcsZy3FxSDCG7PCg48ex2N6NzVh4965VdU1c4uW2LC+ZYKn3oFpZOCb6CZz9xLeU
nyPnVkMptbwNG0vFBxuM5dyHnBopUMxjj1b0g/QtArIsMS0No/Fr5xHIm3Wuig6fBfJukV4cXTR+
4QLHPDFkw5hHajtGm/y+Uu9rbgtNW0ghvsw60KZId5bmOH8oipGwOnpZVWlEZWKvHXyVyHz9Qydq
mdr79do8AKIPrnHlW8vR66ZqMZEeQH4Cxpq8/fELMfCUwxOiJadJ3B0YehVV/XJEdPVO6/bPaOQV
4skA6+NdelOFXJP2mb5I0ykdAk4jDraTA7s8fOGuw9QfX5bFVaTQKSf9VDs8qdI2vXZHY4Kd80dz
ctdXdwEOtSGUAMMp09LEFeXaZBqwJcYex7ct8GEKacLh/JfO1Llgn82WhOeW4G9HnEeK0E9EjElC
aaUgw5Xot0jEsU8Xb3x9sX8um0ia5Nh3QLcMwOZlpTbEHQXtFWyI8nwjSkFBijkH2KABmAVR9jZB
Xnu+eZLvoJKUk39OQoEMnZ8uLAYdbWciXzj2gkQUmXzH98f/+IhY1Ym7XwsdmrgMCyecuTL9Cc5Y
Qkiw/VO+gaevMX8fQsvpox3QVHfu0Thn9mb1aoD8TX/5XrKo2acuic5IopASve2xr4BrrjP+rDHn
fxZNwXSz/3RQCLiHSzop2egEBSgXKdBDBTWRuEy/SHcYyTtnITSPe8cbaxsMnVWeLL2bTnBduDTh
YsTTdXs4+u3FTajsYu4NKW+oRLvSB4LU6amZW9I/mzowTC8TZvt+UsIm2WIAUMuA7bBj2+SPGhoO
zx3++TP0P46qewPVPLcmiwuFMwxEDWyDxYPuR+2AusaY/B3B26IWoepavxXc8/iYPChnsqGQYoR6
NB7/Hn3VCvRf3xy+skp8z/Bi5XJlqkl5hn9q1HGqqavmAK4O49dqsbT4qnL3KVfs1wdRCt8RPsxv
vXiu66jnnDyStyTz6op+HIDClPmJtacIXk2j0SNr87kKG7ZHyMGnUcOux9xFNDToCbA8f6AgWXMX
nxwz15DOFbE7n2WmNEByeolAuY1PDGWvVY+7bkKaXuNq1njFs7GJ9poYFleQbc6x+x8grSlREP3S
Mn78M10li++iZYWbWnpCFy20JvoF0Y+hEzd3fGWAuZguzCMwX58QWKjiHnwygAG7JmNTH14wLDtL
QgvWRaMMwl5Oz2bzg8imzLDPjiXAz3ZrhFdTM2klrbdpy+geqn7Ev5bP43AEeD7ypYGtq3+gTdRF
FY1Q7GM1cSCoFfKoL6n9lyhtk4IgUu9vyx9nVd0g3d0UCyKA8a+E/9+sg4HD5MWNcGQfh1u7icZi
u737TgYYH1r/GbDjLZCsrsIsAfsco8qhUsyUYx2zPXRblZyRqpvWq2h3rz2824eqJq0/y/Hs2OJR
5brLOk6nfr/iCfZ6yP8g+xAboeGBvEVpoihT7kanrD+4cmYpVw16YevI7/Q21thHRAHXj8pEpFdK
Bl5zTcxA3PWPezOMgny1mzBfSVTniEDsP2K2GCIA7Bz5Mwt8zjgn9Tt5C3BtafR+w0FMx+R7vvTE
1oeuQPBgrRIyrfcuxnHM5uK2te24m++Ac2eb0L7//gRZR+ZXrOqXuzl2Wkl+14X4nR7cKVH/8Mj0
rshbWRiKR3OfYS7fdNi6kmSVsHu+B3U2mhNM1lJ7kJf2dBvb7ZKud9+Pp/IZkMxLP4455+qXnSSz
+aqbFCPJJg4Ty9HksGlv1p1Z6l7PA9NXzuiQxVYEOlxjWH9fEY4lwSmY8KKjQO+17mtx9trAiMom
dM9PCyiOIAv2wauvezuGNbdC1IjN62ji7goxcehGOEltv/C/NOwvagHey9s/Hjy41Co6/HP9JGs2
s6hLtyRnmoUGsrLz1KQWd/7v+Y4YxpgxMIaq3kFJqGUyQXZUrnjLq4wMfCfeIBwyUNXsENZVn1Zo
QdUiHj1IOespLtazwJ29SNrENkpW9rDTx4UZv5bomJ3gm0z0YRfXx4/jKM6lw6TwO8aEbs6Wk4nr
YPGjzMsFKlb3kuamBgqDsZkryEwKmMnCyqLjuKWDHujRfEeQEtbysSyq9OzZXRE0qWS12i21hqQX
FAwZZkHGiArkG4+AjdDUJVUx2MMQvxbdiCUm3NsUl37em/EciYKi1Avft+/39kamF3ckDBBmOfio
RcwLYZdPXPJw10m8eXCyqUSsKQiPpZwwBP34FK2PTOTRUSGa66ga0A7vc72BnW3H54NKnudAACWR
7AIVZ85bPx6pxtnqmN1B8qHN2jnbFZIHRye04xTPueiCCatrKHfAmguxYIKXmMe79Wc7dJHqpJ1N
KquxWTRBq3uquEu3RUjphvsaDhkbDD6XVX5Znz+iU67LiDSzjW4iCZMwMFP/qwXtbhpRtxDe/18T
wjPI5tSiLdsaPpQNqdCfCfVsJVLEibfgGCa4NWy9ZIz92Oeh306qiJ+omvVwR2r3jg1bl6+jYgxC
RJBFH/hkrTC+viDnUKlTE34mbbkBj+2rCESJ88+F30FD06Nkg6aO7cc7zV1YCuLLL8qL6AO8ssKG
K4IC4Dmcd1XsZVlYjwfhADp5hqF/p9SX29/qTa+kEJmhtpIxTmS77hpivJmN55ODLgfB9VyIjKw2
Ny+C2ZUq3Cj/jyQUNyNYc2yh4qjoCHwlSo9SxWZRuOKeFSq5gNW2WAfynT49SX0IYNQxDWxsl/7W
yCk+BBNNu06qfgu6iOSzcuHBZrCCTIges7B+HXigXu+vDyJxPmLoT5yc6cfQlHAeEwE8Mte76Gpl
GSwIxXR5tJ6ZPFZT/JVkyXN/9CGN5wNWOyNupqQufj9fGA7v1UuIsCe0GCa5sQV0OFqhOAtZpSys
1QBeiVnZa9/XAGqXK2w6M4ZDjI1DJXttkGCRdb0MI/Efh6pZNaK3p1V0Ev/dzIKDHsbFzfBtLv32
SkSCG3aWiT8zffPE7aUZoVvyXFaXJtluTkW9f34amEq5FNr63FHxEy50jkelXKr7LPSpLxuSSYR5
n3O7JkSXZBG6UxnfhZ4LxFxFXsc4TP5NRs3aJ3+dp4qIj3vSIHyzh0YPe4OBppIT4cO4R6qRMtGy
2nXjj7e2i7ixxiVxphtxSCJYx8gpZ4dRxlFeH1eBv8ocrXrP7JV/Y9M5FHH1gblWCCRuJs7pMDOP
ChrP1kqmejb2WjrjmluXGM1xoHXvxLfo8NffcmSb+DzRmwfnwzLe/0AkvgJfHEdeTziJXSKoDj48
MaSVYTpUuxl1M+SrmObOIX5Yw2X4/Q8b7FXCzcDQSlbK8hUZXkF0pye8jlcG+ToivfR3S2YwVrSk
QsaMh8WQ57Lj9ZHHC+J3FsQLU4hJmKE+yn0lrqpn2MRI8xKZYMnvutGX5OWKLPDW6ddiq20Ba5VK
IihfnMrg7t08oRRaffWTfLP9PlzwHqTIt3DFxB2oyGZ+sFnQS2EXGBpO05qJYp3iiKQYMSscT1Ot
HACThu8SobONhPVYSysFbzbmlPvT379MCUP3UWenkds8t4wuYcKZQu0lqZUyre9gxQrP78jRPtBn
Tsa27Y6Bwu+N/ZnHJbM7UBn6pJ2BLgjwue6NWoRDzsYkGcxlDfeR50D5kSPtDqFBRyJSJ704IU+f
XQ6VqZk5gOLYO4EY6BcJ+hYRvb1gxdqV+qNmuYSY7UtbuRUyT2IHn9WFRbJrES/TFwitrw5zNP4M
lOBUFSHX2+SU0l7dIn/Z2mWunfLW9NC6Rz4HtwAp8FruxKKg9fkDxteKc/eQ1bdR4yMx2MGwYzf1
X0mkeIYU/5WHqAjYRqVdqYQ6jMQvkH3IFyTZlLLSMymq0uQW567RhCuiSZV+YrhcPaKKYDA7/hWo
dReaOdPdGQ6WK9gxqI2fwNpQb1qZZE25yrbJXlTr1MgLgRrF13Q/3T+MPC+tiMjS9oHDFsUaEWWJ
V+P7/UXZpFAH4JJz1tnK/9bIIz3LrP+DFEVkrTD+gguAysarVdxgn5FKHiVKF+Hupx7ZvWMpSOtK
FIwEh32RfmPAudLFsbsAqlaDIURtq7WFAMvpBbbY2+LZJaBEg1FMUWn5aKt+4BIeC2ccCb3sE36Y
DvMIxgXuCudrzgLVt8D+n+tPlT8g8/sjZj7rpvyLVEVIlrUgpzuvJUMLFO+4SqEcRaJQ0nYov5en
Jxhig9l3euLtw1x+4NOwn4tPZfQ8mwTwkf4IwHFCyGjXWLeh40W7loejK2F2xjsiAR+4wILTvCEy
LLNNMxxwU3oP2+Q3utFMXSxaNygw01FCdHA1lAWIJf5/gKWteoL3G25i/DrmMQsent2ByxjgSw3t
+W/oHtbft9AVHPIcIakRwoMZS71pIVHGyOPvGT8aNyc9YE8Lb6Pz67dYtBwUz5sAqTmuAXvkanKF
uDF70aMKzzJQkE2prYNvGUeNFbEpR5F6NPZB4TmEDrSJ9s9v3SMLg2LpePMQ6Pj1+0KKVvOwdE8r
wruD/35eWlEk+JEPVxr9PCnvbADwJTuLTj0aPeX/r1wNrTUw4ljJ7ySQDg5samNOocq/gau9u5Q7
FEORAOyXpa/RXNSG2Xl0v/4wGPc9U7XXZOok0LzDzxJAtpdLVny/HT+oa+UCmJ9JmtaNVn6Mh7Ub
mUNGRj2yXAstziNJ25TENKCUCRHBi7jxB6Ja1+LUtiXoOkvOIyjXkgu3kEUIE3vHevs31eBY2uZ6
EAzFV0aiTDk8SiOEv+36wqx8YDlpwH+vH9ObmD1XckxelCp9Vm48hNxiLSpoWR7XWYy3CsXmOC9R
bcwlWSug7806zgU5QH/+2ChIb5f8Gw4n7vHUVs7hTh3xPyHtXrO+iy4O1KqYd0JDVm39B0kkxf6n
vH1E1Y55wIz7VNjkYtx6sqDeGLqhrjzJdcsDCczmn43dUvdnp4facSKY7hZf7/mdrzP3eMieQTt5
6GSj2jjxBaNgjpoefzskkp+G58jkCat5MpJM6Gjx/QbOq0v2IR3A8TKIXQekc2p8FHQrVa1ZQfNF
1WtRo29HuHEs9W7j+VQBLTKahNFFXQ/nfwprbKMzFJYiPYyTCCWJkKeaiNqjWLT3cy1/T9Ne6LAo
y4GxtwSHvX6vBMm3GxIE8EbRiVUjqqiBXhVBqNhR0hCbS8+MSHOdl/RNs/m0EehTJwJfx0Plr4Zf
Lok+EyKMzILkv93TwMgC2fwW/jCH42Ty9FD7Dgs405XDtHKT6CAecSUJrWGbsuOHIoDjrPg/9o5l
m1B3Kp9E+5ybwjRRFy8sK69SUH4IDusS9oDmqt9X2DOPCcXT/gAY+0dGzvGeM7cbFkwpyzCDBzx5
L1olz6XrPIiJZXarMb3xoCp1A3kW+OafQU+KSdpii9H2AFkKcqvJQa9bCCDw4i2VEcqy/8iQBPV2
/999B9rATLsEniIeSl6+Gd0GmZ9UxWdhyLnm3KWe0SA+gZlhNl7wtLkoz0TF9Uqvkk+tr+lS1tju
nNRKeGJsPoVMHj9WhZwrBp+/zoiYqMAyNZmOvBs/2veziw0UqcrnjVuA8Hatpg+9TCjleXakRtSM
WC9kQU66/xZMPNLPjiKYGEzvH5I/tOqOg8jJc0adjfNlS1BNO8KJ/MsS2Jg5QosgUVapRNXBqK9U
tDe4GaDiXwVkvCq7q7a3SwCrE+Ttchnxql8k1J17ueDZKOcYXyDeVmp+LRsmNUYbj1e3zaRrSX0f
N6boYB93vqhhQ6ShTgL1TSZcO4/NrJI53URx7Sls+KAhCvrvCvC8oBdU+43b4vFLF1if7DXnoy8d
P4MezJpZ8mXVlyxKVjkEwpQ98TiUJqEcMfOL80KeCpo7vpkQOtTAQmoBkwtdxdJRTeOIGcpbRug5
R43h1oMJQiDDQICkQ7Q4Oi8UFkbtm43u1c5PPllTi4SYrUtTJBl1i9SUVdc7H7ax2ovQcmss9X6c
3kFirO73FNzmE5TDr+daG5d2L5J1tLlocdvUqgEnE+4NEYoono0Yw3R1jAbrfua48tCkKdoV3gUR
vR5Zp9Tc+P8YiwKD64Qo4lGLbSEKE6unYwDoFq0MdNgUKEC88HNkAByaRGOl7nC8V1GmIbYVocAs
25mqVIMi1lirQOd/hmyr+OM4839Z7abJcuyqJkRNI+SgQu2YZ1RlCZ42xp1qJpZYc6f8Vg1W3GYq
Sj6py+ELgX5gPFHLO6h/iOeXlk8I1O43FQvNM+3i8JiG2iwnTTAGW7Sn5oJY0ejIQGimgmWLv6z8
6xx0QbRpXIhhn41Z+6PhzrN2tSMeVWn1RJ8x4xWTsFNx6Pdx6juFj4diYBbgou9DgcdXbDyCx5sB
tdyrxd+YDA4irs5jfZT/w93A2wYzuBlqbCFJbJzAeJWg45UFiGaIMNh7NzIQ1xAkuEMD6FtRev4o
rxp12kEhFPLV8+RV0rCYQVRMF5RAPhvY8jgiZ634dGr3iiCXYaa8bUUzmCskTLixezG3udnMBwYI
zHH19dkgEtQFoHsHsPq7jzDXqReQwF+ZznYluLrx5Hh5Z7700ZAwEYWBk3B6ovWpRkMR7p/SHorI
ZKCrLGXO9Mqo4eiGdqeQbGBaeFSF9Ec2yOEwa4zj83bnxtuf1y9XrGwSgyoo9WZfK0z+YzRnRSVW
ntd1PS+Vx7V9vKuICWqHRYhUyWafE2tMUVeJoejoEgEcGheQeJoEIJUy9i4WY+XHleQUIypa31uW
mR5HPXkXU6Mq2iTmcqtpgZnffCvc73y5Q6VYB2suo9659yEtYTDVkhco508z6Qtob4XjnLJQWkJk
j96h/0bcJV3IR5d8TCEZva1t504f6cSHgoYj9NMvOgQPundIBTIyGNUO9N77kdFktyI8GWy6jqL1
x+C1TjSUcBnHt97oObCfW9ord2bG8Pt8eDzzHwACbK9ukZOEXMBziwAtNe8sxzkVATz2LoFd34q4
QhAzzRnhggm0wfkFqnviVq2f0LLh4hxXKMFExy7z7uiZzDt1MhHUrWZhckr2ROsIPjAxyhy4ajCQ
n9XFnmPewY0zc3cYIfmgpgI5Lf64TXeREmfC11NxrqqOG5TgbNLVdqhMlsMLLQQC2W7k60XdUjAQ
Lec1YaH/Fgr58F4jI2cm1X6LgPIS+sX8+Q7a8z4q/eSUvUITuzMpq4iGxP27onaTATlDJfSkuX6M
KrmqgOxDrEyhnN5mX8fv49hA4pDg7ZhXwcyQDeOqIPa8JTUtrGoEQDw7yjruID8YCsoa1Z3d2gU+
/JSAuCOqjOxLB0AqlA/h25i+zgD/1eDia1m9U0pAMuknZKzddTKsYXrAoJd2jPVTXnU7MsGSZOO8
6I9kPwZvyJpSvgvzkWjxv7oIOq2CD4NpWnIxf+swJZxE6cAu9W/UC2MNyX00muEmEwKxggfWum6X
eB3NVOVb5iLuSVlIM7/7NGgJrw46YWfxshy3VDoicWLaW9WYGearR+m+mP6k65ogAigeNM6L7nET
YjpgpJsH5g+DShuLIHSmREaNBvFBPnfMinzTS7xUU5Z+pCuYoos++mM99Dh+nY50KvGOEqZRU/e3
j6dcWiuXzolgPdVMuCCptINA8YxeylKYkBPLxy2agOc8HwKe6Skdodk3PZ7kTzubUASbRKMnpHr3
Kt2PzLmFfGRkm90/W/zs4Xx9npJqvpeaonwKOgs9IjhTgao7g12ySUncOcJeZW5XLa5t90DUE82c
KNWmcxqwaET7zas+13LTKjOskyEsNu+niV5ktk4hS5eSKesY6hHA6oJqF1b7QkrupTgcJ71jgbEZ
kbvpKD2EGWrj0oFkO+y9GqRm2m2xUtjF+CWKFU7mJWfsmfECRSXs8rOJpYiE5xzmPNAteyVF5zJv
NVFwSK63u1JzeeaMfLxiABnziYy1r58y8N06Gsvl+WUH4acTa3weYYHkACxY0cNCpAjOkCy80h2M
wwoe7bWrYgCatf4x76Lgo0M6lg3neoNw4tZAQqB4+UgoNMhS7eIXg11lKR0clwCr860zkHzi2yAc
SKEsFHJ9MbDHKxmr5hb4r4sKWrh/d24pdFoxVv+Nl9IIHmo0RhyzxoZ0f2Yxqo3V1dJyuxrj5CUc
IRJuKCREF5+6Q6RM/dru7R2b4PrwRMD8ODbDcBRQkWB2TIjqj4LGs+bMyjaszsmRyOTsTdvNg6iR
KRnOO2q4pVA/VQ04uDcU5hT1QIJbGD3LDPLWDPUM0Rcouh6CJirclTWscARAfJmflLfzjRHGACxZ
ukoFJXeTKkrtrYVbjjdtaONSukgipb1NtJyQdzbzj3bnpfkJy9njrFxal0G/w9PKSarCQfTG5z2k
lDE2zMbmYDIswo9/NJuI6UwC8ZWa7OP46qnQruHhy7Tu/K1ZUOmsgIIhsCeyAaMk6S3ekqblC0YP
5oCwUIV4PC93MuyOEgy18eMJef5DQpsxZKPmjCfxUHkvYCuOoTA+k2sDRsJcZjAmWWSLpptXgFaR
DKe5vghQXyYo6L9Nw0KlTTxG2jLD6Ozod+JVgSmZRofdEEXmS5PPkBA0Z9dS/ts+JK7lZWM9D7aW
JiezdrTPmvzEAE22ZAXHkl3rEKDrOenGYzQi2UN2FdUxE935w1XVGubbAUuyYOJ5VKLzcAsFfYvx
LtZyVocN85tEPf5obUT4v/q8DyLN7Vn+rEljTOnsVNOOaMWSplnf1O3jGHA3gVPDWuj7cUz0v21w
v7Cvr6kl38yMeEoF4L3AeMcj7LTDOgvuzWVSKQF22xzd/IDNJB3TyfS/GMfmS/W9ZN6I6/4C0jlX
YMOEStTulHigVMgBgGGu6JVDfJRFXcc3Fc0M3Tih7smjyTPDpv1VJqA3AgvCpVTNxllgIgwoJXtx
PJA+4iawoi8nF/XRmJhRHdT4G+JSZoc/f2Z73V2EWyCtSzKZrkwVTYoA/xgMzuy7BZII1MfpJNQx
diQxoD+Z3de4hkdqiwGRQIluMGb02AAlDfQa4/i69vfo9q2O57MeO15A/axWLMMxQa6HolRC5VSE
h7TwzPj+0D7i69SjlnAOyEEgAAOW2pZEMGl/yLiZVrFU7swXm4nTEaJGRUC9t4C16m1BVrwuYMG8
eeLJYm9djepKk64yUiJ8lgFbIXnr9ponzaUEcgcjUm6AkEWYGHwSmfpRCv3o7g/j05l0o6klsom1
yI00skplgxLGbFW4KuJRziSLON/gU1CGfIF+DT8qxe+kDFL2B967mghm9hKivYrjocDd5Rfv4nKz
z27nBkGDWf6jZ8ICgkXFDR9i2uZ5Ibh3cGXx0eUjHYxzsCImHmyGFIMnSbXYKj/Lcd8LCBBX88wA
eqKG1suCa7VU0jubyZPFhLcHjrySmZkVnL4FAma7SBntX+lRNmepWH2hS9J1rfyx406oMjGi9I3A
uqaj+9cCvSnm0LFCPHnXbzq9SGmS1Gl2pFZd4ItPLPIzXUHIdZTAC7fXE5zBA5spKR+G+rGnB5cB
J5m113wniyz7+11nozPHDHNEgWU7J7Ij4xbOxldnMcrwh7Vddlp3O8hYxIBcaM8A0eYmc7smtwQP
SCxc6HE5ItIkFZJTsYIY7fDN3cLdiZNtyf/sH9zDR0E3W9msudp1ktx5G/7RoEWveV3BC0RRCdDw
AqRnWyeIkhRM3ecBjFffV60nDL/hGoIarJNx6S5Jp25GOKfMEgYxAGw3I1nlNUrpS6AIsCs/Yaqh
AmLhW3j+/6HIVLc7wDsJyBVSrZZPatzxxnwfeZS4h+MOED3feeY8EIwAwK1J/tW5Kt1R6TStfI/2
GmagTuA0vnNm1GpeU012SZihpXoaAv1ptjvHbFjya49QcUjh0KV6J+7hCL3boAbn8j9AFKkTroR9
cBVveB8ESmjNd/X9dh+WxgEZFd6odbjqGJl4TjENZDnC+s1OkYDPJ1+bq4vmwU58E44HDK9stUed
e6FBm20+N6ww7yCn2tXuljYLHpos7gg4AlQ+1TuLZMx+4bu6z4HbG/gAGzYXbi0H8sm+z01INS94
Ptg2kEP64RY4dGcC8wwk5cXiP1CajYRZLXcXODW5g53CXel5oL4yvN6yLHI+J5mQh4Rrq1vXmz/b
ZMhr+X6gorvYnA3AmiGWGD6C4etSiWjmGA2nZ3NiysOEYVigmEQ9zWn7oHX45SOZvgOfIGCwW5ST
VbyPVbQTJLdFaocsyY/Ebd1slDmlaSSMzkhyeqKh9h1LrqqI8ML6bgs2+GocqEHN0HhNf6EIvQ1E
HZ+CcuTHBF2yLQ59CAcBZPlnMWipawAesBMUeZGOhFm59T5EmSMaQbQGCcFSBvFY6SD5cRvFj8pk
qPoSnCNqNMJZ+yf/txzVTJtFBwbFQ1ZT9l1oMbs44V3DZZ1e2b9CNLfS/AuR3Maoj8ytVxL6itrx
5wSiW8k2kWhJ5M5THLtlw7D9yobR4S63/1uZ5Qz/Ta9CKMi/Mcw7TS9JwuWnDG5mJTL/P6s90O7B
nqkr3G+Dlisg1fefGPbWzFkNr2p49Rd2Pm2+ufddh/3ZnSM0EFTqAqdjHiBJ9VjCAwFwvkpPf6X2
dEEj1T+UBBebS3iWrsBSEvTbLoG0QH/1GS2dd7wxrEGhJlacJTaEEMUJCSYojIoMcRMRybTkyXIa
Z1mXJaqvkRwzr0EN9OVmexd12f6TVSNkw/FbD1U1afV6CfvPSaZEoQxFRK9B14c4WsEqpahQwHM3
/uCEhxrWu1dFb+8wXUd4fRu/mcMbmCrWgsxCVWEhRn69q9bFMvmTK93wHHYohHd3p9iM9qXVjwQi
28ViPOM93x7GrB+uJ9WV+ZRlGIPGuTyCiVXuNSo45CaUPqZTyUwjIYTRv4I2JeI1KIUMUBK/0zB7
kszPtbvpL68nkR7CUnr69vK+bAEDSP7F64Th/631Cb2vGUvx2Zb0YbEkXeonPL+gOyYzHX1qqKR5
PcwxM+GShGIUKUGLmZgfCNhKXNWerXyaAu55p5CkAX59r7W7/G3XyX04HtApb4d+mLh+WG3EyiLf
RtvpdinwhDtQfmbS2WfetsNEKEddt2QD4Dx6zo8uWQMujl5pRvYsvkDE8NJrRpAwiANXfELgscIo
BFyXYGufIccYJDgv2eNpOAAUy+xG4yrwyt1xaoWNX8Ep++gMJr3Rqp2XvHpl+jMhmhILWFIV+pCg
dhpe2uBmlOZNNFHRXOqFOYXIHpkZiGvdTuh5bWgQuMVQ6Md7pI5LH1CvdriXlkBplxWjIxwCmDAZ
6+su+8aq3rV9yPxF/lrBYV/s1SZxjbImZlhERLhapeSeCsWEipD/uLO8Fe6ZAX/t+qem0d0nblhX
b2N7sLZ9qHp3uoy2wAPfVhYsnIWzk2dfekivntYCHBQmZg3nM1whik1/sDdVhn4z793HUGlziK1U
tNgPhhr4vfCZhknlMku1bFbfTMS2GZqTWEymJfZnyqEKjK9uQ8ZEVwQ4o6GXiPTMIJXgwKi3v5/u
lZwWeDjGerk/3jG3wPYuqJu2G+2hOOuYF4AUGEeCCgNKWd06Yo6R6aM6iU9UWjNBhXMa23NdJMJo
RQvugtr4j8zrABT9H2XiWM9NUi9qEwOUFVnJujS7WSCYzn4VGDvWEudrnnVGZ59qty+DdePQ+6Do
KdC58GSfC+VUO4IWW1sOyZ7+Lm0YhbTU2xTtcBkNjkSo0A4vblL/7ncBn4iOH4luaIAkb9iVdX4V
edJBcWmM0ljd6A725du8dZ0ABFws4GO+oYynE4OE6Urzkl+8BlMBP1k4xUoXRcbDw9d8LKFFFPIf
81Q6WOs5bMZYfrl8QNtvu8qmd8fdQiV0p/PDYOIpziCWS4Ml2S/G8cpVwvGW7vuqaNvdY06GPEar
yTMFZxCSALOuF69bvyclx1D6GQHphVYrVJaNaXRIIsi/7rM09AxuJdw8LYwIRnb9F3AU97Lxt2Yz
ApVe4PGGj0EDz+NuB0r01yVLy+3Q7fyGblzCT5eqjRQu+wq766r+QG2yD4JIkFC+c4BNfnPYgEP2
OtHLeeR3lSYMri4zNQKbEPhg7oMqdGwyM3f26H2Saw2jzGjto4t56wESCFuWPX9BQSaedUT4ujFd
nRKnOJfCN4aStqrArJSrtiBv1lOdNOGdOjq04rnLz/rSvxzg6yEoOyFvsF9ulRboQRF7PkdDOsUC
ekFa11O7KlXHJ6/yjFx4uSyEqaYVPMY43x6ZTfxF7d5+p/+sXf0tqeE9a606KBcaQsFWhlYGYrRl
TibOsQ2xdwe2QPyS4Z1p2y4lh/Af4wBEiGeTUsAbeEjOa4PqRnBRIBg655NBRTZsPilVm53/HBE2
ZpKIhMVeV+Q+M35L/C0NvyVcPemL3+9Y7Gw9iMmhaqLezU2Amy6FR3wB0uFaVceK9TYZpBAF3fGy
Sn6NsGGyyJ5PsirmtZS9NE3G2CbSvpAO9gXg/0xB2HXf5sXAYfCoWfsH02Z+Lt/kMPLvexQi1D8P
RgErFkZ8Co0OvGJXB2iYzpfkpeXT/3DDh8UJJuleIJxlbYuqH03ZlG21fKeQpIQjBE2hPeuun59Q
BzBa9eEj3YOVSAyneavqHFNaEEyXYG83JptnQa3RLAP6qxkwbm6DN+0xjk0iKQpAfXaP0wyn6sBO
uca91JctC4Yyvb838U/YJtXFjdURsz1ExldBsTB0kkkaowmBbbXr6il0r4M78FDotLyuOGzPMrie
KfvZ1biAI4heNyXLY2L9t3XT9+81ULu0g3CvUI8gvnDy/ZfcnXxopDZPzNeVWF+vpZMcvZRmcEGY
3ChSDnS+E1d3KUQddyB0iyZ3x8zpzAuSDcc/kibe3YVQUipShTQXf5MLrH+JeL5Zsa/kDqhHSPFw
HvSrlUb/0FhepbUxXcDKLOiSqr/dvLoAnZi3RexTswfPKGpwhrlGjpwVGZ4wOmZpfiuxnb8b0RYh
64spe3+8peyawVL6WPArBOzvgSH5s6cv2yu150pMcRIhyK7LnPfIF6qCCKa7njya7wEHlISxFBeq
C/NwR6oNs99HpNOfMWjssPun+eTpq90JzWvaqqP7rIwdxuRbovmYbbo5WMiuKA9ukNQ7qXes3iFB
p+c3ghUcIdMbkBV++b/kO22FkMQlOAtTEqrlFZOUzdJrdlHynuvm42lpmovef4elztuqT22MCNZZ
I+HPluxr9KYBd2xYfX0csNakCiXm6q8BJEPZOsNIqW3b8Q/5yn/8752tqiJChlARpVVsLnERihIt
BjE/LPfNOaj4YB5mQlP5hHVKhVNDM1nE6+uYEZKNBvftwcfzbQ7znDL4sdShmmQ9ajMLAxMK2ejk
sX+KWccTWGc3owsxegAYbByMxiqxyAQSZuVjWrQdfM0+kReVpw2FtS0Ws/lQyHCQRAcFcZrqxoKh
6e9RZWy62TwEY4oyR3j+OPrI3w7UvI5x3TyEOy2tUxDfwy3t7sIJtKk1x2tauaZWMm53rZBgzbKA
rnEXaH4WCE9II0k4iV9ra0Iv2O/tIXhzaQglAInjOUU7PjhORhlrJ2Q4TAtR+KJwJPt5XinMy01f
QkXEw+p4KkgxxBE2kXksG61sPvVYQvDFw61x6HtIYzXSQZf4fFgShcJgjLvWiHX3UzB9mlWmhbac
D2KlkuV70WsZWR0KSpVWyUmPqfz8IL4ac1K9r4wDA4xuhRmDEFmgwS70HHgE6QYfP9aim1L18U/v
si8PSdkjpfFjfF+GTdrDRcxTpkme8h3WK2CHXQ7RZLyk2+PPd2la7NI5wW2za21b++qPTXoZoaHq
w8W1YsT4D5h4fT5mbQXpZPzk/QkS9wiieff3+6lRxlnsGD60MczJ/XSa8LyA64VH8A1UA6kZolW5
PQw8cvxk1nloJFsRwzG2a8/08qEGS7K13mbzUuBxVSTQmW0Ayw5XOLwRlr7ls/OvsK+lzGDD9RvT
GmUIyYnlPIaS/wDPdYp2f+ElCjn7LHqOccNsPdEmI8Tx8xnvmxDtQAndMAxGFEHQd9gSjDNkX4rn
v0QlaPIFHDGhKiCICKrh2kCbKJ12U/swwoEVHrnUaBfKzFXjrD0rDYdGTFW7tBBd5lYqC0zpzKmd
e1lPYmXujv1Qlzy9WMsiAjiIoV5Bt/XwX7L4vv2rO8+dYtelDvvd4WVeju/2X4yceL5C6VjbG/h9
niJv5tk244WLArd5vjAF+BKPhb2pIEfQ7N2naKROtSXKeRchqqiQdmB4XQmDXwUqQ81bo45wONmu
O6Hf4J6gy2hUV6nc2PvRbq/zyQ6YFdSQ3MdWBELpOL4AKKprTBbBRcNE7D9RIv6YUvZzENVXwvjT
RjeQV35m2BDz+6Xu1q2nSC9/7GkDIsI0ZtETbqSQJPjt5AbxivqUu7+YsS8cKl7DQs6ukE1fMLP3
Tk9o1ipLmBrmlOVMcG0aeMAOwGfPMncva1e6kl/blKg0NXdjvrCKxwzaB7inSTDiZPNotaNf8S8A
4vMGJpC9hLkftlsdk4s+MPbz6kLFccU5lyWVeZsHETjdOjRXntzx040qieBGnsU+4B7AEIAFNuGw
2kfs5e1U1a3zpvHtBruAc6q1er7RAzr/NYXdpQH0BuzJ8lMDGfsmEJ9BqLgMoM5xxlO8mevC7ONu
fS591EW9T/JDMyXi8/3XXiGipcLP2xmcEA0TRs5rZueOMSQk9do0bycDkB+67kT9mKxHhFeOICy2
5VhedPfM93pZbbixHw03toNKZFsss9ZTY+/Rj2f3a+ywFmplXEbR6JlYqu7STdirremUt2qgSoAb
o/l54Vfjvx1DT6MU2/D5Vpmo1wHrIkodrad6swUJErOk0Fcqsim9lGZP/cvN2a07+7OROKq72nOh
OfOvr1YUxjL04hv8/cucVFdNZ3pxZA+UN3tiaTQWyn/mXaq9N+dInsmHJiQCp91a71nZL4SjEJzc
k4cOs6J099arlfwqR1s2tAf0Db59JoYg3jm2uWV0y81MdqjxlJ7yym1gCUnzgkJazcD1CCA41KMP
oZVC6+ZNbz8sGZrR+QkuEHWqTzNp61XlPgPNvTdG1HXWDyr0Ym1eZKzFL0W/69ghaCmm1SgkMNFd
l+1P17+TkpEgD7cPSFf1+JyMv/65Xd9YvFxSiKMnpbpvn7hlK0ZTUVPsccuo5Mb3jpzPLdB3k9k2
JUd2RR841HomH7mTRn2qPy+rgoSUB1KV4wRP4LgSiY0OTAqin95gRdx8VmMae7YvQVLFxFq4yAaT
18dyJNC2GKAovQ9wMDK5QEzaxeXtlqh29qTk1GHqJkN3d6RgoGY1JU0oOKi91/+CU/mYw1pTw687
O8dXB4SMx5qwidaotilCOs6YsDHNBv0Fpf/TgqBS7kwesCaLMQnjtorzBBCPmzhSQ1qLlfP8+Mxg
Uzsp/2LJHmzLsVybdnyXKHhsOgpsmL9YiQZCEd1wJDD5oDSLQUAdR7rdq8Flu0FIod960Ey/Ins2
uoW7jD+AUBavT4Ga7iGiTIt3T67EVLjW7tY7J6PCJVCbR9oTG0RZcRZxHJjc+q58a8sMRXEtuBzU
h4SMXO72der2bgTZkr8LTw0fGk0jHZzKzt5iyUMMg0yOkuOA8JTFdUebRz3N+PHTcaLKd68GNm96
+Lx3M8xzDsS6E5WKFXA+cOCdpVfkJkDhFPK2sKfWwPlJUr5SNk/Hwpimiq6eFVfjfww7MrsDWm8o
0KlM89xANPhdybcTvTP9kbRHXNmMp/2Cx7J6aWHjlRdoFPwwji9KPzuCQe/R2/SgCH/wofQIVk8X
lcouSm+eZ5D0PFZYI1an4Kk4tJ+sYAZFQCQWezZ4sMLa7cbMa07wu7bya7v4dJNqAAJsS6sOehcE
eIz1rIwkE480cccRcvn62zVsRh1MmIWRFBIMDCmYkwf+c7V3X0lLNraGhpTq0ElXjiOC0JCSeCkc
aszR0cRhbHK3Q12r/EVsm8AF3uhZfHW4G7wHtO7XE7GMP1tZPEVqtVqBSl5Hv891C3BbaWsif5K/
WAayC+mKWfAHu91vsYmYMuxIoCPjEn2PesRTmqNujhaQO73eQEyNuqEoHzbnsyevKuXSGdZps+kr
YXjGG66ewcTrJYJaO/BJE9AGn/DfRqD6teHi5PrlTL/nk/u8BUCc9oRiqDBGOAP1nZ11L+Vs9wHQ
w706jlTnReoZbrx+x/N5JdxYkafltDJK0wOEpLxAHPIn9uRiIJCBkZZ0vuX39XPqWETTNxFEnSkd
b0l1cfMSsbLxdXAeCWnKYx1VPgAPHfekSmKLFBN+/JOSrSEQRZ/2KInfScjkRQ+QX+niQ5+sTonb
F31BIJ7PSqPhKI8HnQJSgQR1uviDRMcaBwiDC+6F5EDA3b22DSIHTsaHb22M42+cdBbZ5gwXoh4w
dhDwKOKO80rdr02zMDjgmW5dzJkzIYLc7cOLZ5WpO+SgkX8uWPSHHv3kIpzD3czMV3nH/jCN/iyD
NwNfyK8kXMo56/7j6uDhC3gIVNvAKihOtvBXU1f/o1h3lwa9LD8QkjNcKrqcwljJo62G4jxvvwlA
7Z0R6DA+hZuFL1AbpJwOBQe3dfST+RfEMCgbiJ2iJiIAaI/cc2ffa61VOo0388Jp85en11mVuYYr
6LoLshlcMXdzfLXE2Vjc9/rSeBVWGsalls4g5GTv75VyAkuNpRveplEgyvxLkjT4RMEWykixhG8k
4dDxPmhPRBBHYTYkPcHhVRyblximtx1tVUxK9k0Phpuixg35qPW818Ykm6/BmyXvU1PQpuQ/YUlZ
R1C0lMgmBtgDzyFWqU9Xp0xEz4z6ciP6t9R5wpILNQ1jJqpQg1xIfCZWr8vWloFUoxNehd4fBWla
35cVB6mSzrIquqmdwVNrr79c2LVntAtLQLap91npY7oasLKcUbrTxlEQVymqZmXE6751cmMwejDz
oCfUns5+SwnJ21LZkDwwfv1KhQ12IZ/FqUHpu4/o/O1Ut2j0xL5STkbHG90gZ1NwnEjXucio4lGc
X9tuOOaBg2CumjizlsTTxMDMmQkC0uJ+CBuaXjKWBwZshXYa5FezjTXTJq6KsgKbJeHpMJO+r2WZ
bOLxrqJlSqc9ECfyLIr8Sy/ljAFFy5MDgsI/ObkzWD8TCYNAZMTeER5R/EF3sAJrNwzMZk2JiZnE
6TzQyVPiml7EUqCWD9QSZd8eVWsu7eQCXDRZcoMp8yc4Aom9o3jICa5zVaby65u8YRqk5khN9lXH
sSPraGtA311pjtiowx8mdD7mkFY847qj3V34C1/9dGyBpV9VqS8A05UbCTKj3E92NEpn7AehQVR8
vKXIxdv3fr31NE8s+0Y72edg47oWm9nhpm0tMB3A5mXPMJfEGLjJU4tx+fsfsrl1P0j9J6FbCLlm
qJ1CpDH6RylndJL9q8KEZ47VQnRJnyef2r32kmcSNznYGNmnGOXuaYf+7Ij2YUuIS+h5ocOHNO0p
3QmcTOhpGmf9wzNTQjU9CGKWRl3+iivXL4+17W4atj5Gl3zRXcx1diFX7oFY8AHckq9DKJk00SlZ
xq5IrUVu0sOvBg4Tn04SNNegFkvRk7y1p+HfRBoelmLeffZKtBGocRWkOPBFfuu7NA4YsrG4Cl/4
kjXQiU+onYU5iLPa1+FA2dMA6vbfyhgF2QllywQpEIjF6+pL3YUcv5mauy9XvDkmzPqhDJDSZQZO
AwC0uRRefjsStO5W1BzpN2d5ffCfXv8UACUqSW3hs6xbT65dYD1PBGCtCp864OCuhYpVfMqaRtUy
QpsFpMlGHqTlcBNoAn6kZTxLyx8Y2CbcfOvCmtiP8KJV13NPl3IkpHCUv5TKRpAlQyNixWG7TOdl
oyABR8+z/G2kCeOn6zh316pMLv0Pr6ga9IYMdGrLaK9RMqkkc9e+YHTyw62olZyc++Gi9T+9m+zs
PJ/ZJCOd3DkQ+J1CnVxbGFSv4ADfW5f9v7CMCMWJJ18eclgoEKD0aB+h+6p9t4wxC8fsIGHXZqwv
UEe0b0l2ImSPdfNw2wgidnsFTQqtTUQk6aUoVlBPX7Svi+U1BxwshM8cdi/6EWiE2XKHSfeSdYSl
Kb7Yyk7oxzLOazrqJa6HBzr/IQ79NEZjWMrrnQtzyH8ECAIV3oDRJx8HqpSdyi0u2vMwNbY3/vvG
eeJZofyNm2Fib3QgihW0pUrKPuenEoaaD+9UO+WPvOT75wV1B2Unt986w2B+4hoXhELOjkDrsMif
ay49tvLBZizJQLqIK5sk9TTcY2ekOEbJb76bzh6Bbsx6LI+PX5Pl+mkaXcXh6WmVeeQ1BBzjtv13
uYnYhdaC9etQeM0tSXtrUL2wjilnv1dyy8QrdNmoRnKcZy/egvlidanYd/tC1rD7GkoWOK/UAKbu
+yf59a1QVG4mfMqZ40roDabcY7dKF9huq58iBBY3Rn3URV5hZCNkQa6GIrEyYO5KrzbzXhLDefcj
QgYNs8+BwmRxWxdXVlEyUUqo7dGcepViKgWxy6cPk+x86YYMnCE+hCsKMQMyHR5J4TX3KqvXiV8f
40hyeY6RU5+3L34x/Pgm0es9+RU8HF4tq1NfNbqvyg8uVKK6LZuH6q2kAvmuWIMmeTdR+zAEsZ1F
yETtGEdVqi63LTAkfuW14T5ZZkbAT9Hsj6dljK5ossAKAnymdGPBvoSXQMSgzhj990mr3k7Fu8CS
/ERVmD4fveaB3fQ/wdTMD5/8H5KLV2huWD3c0uBnM5HB1N7Qpo9CL2eWexPRjNJVQPizs4lA+MUo
grgvr7eLdeijjMDWBvMT8eEwo96s/UOStA4JhRG0QGVs4afThUEG0ypjk7Hbknr61Cn4nTOzT/+M
Vfq57UkugsGPwMu6qKCcQ0BKidCk2303UN6mBTFR2qz+X7nqSRVc4CRnADLR9w31zgZOMeM1uSKA
mUY2zxcO2ZLs0C8z4EA4fuASacS/3tuiKhOfs3saVBeHHC8NnPbcbqYen4LzLPmYuOD1cupEP+rP
OJUldLreb7VD2/VSB+qUz/cGDUCQzxvaRaUqNL/ki1qc7hdCHXiv72Cxb4N8RhMokf+sJ44shymC
CVZCE6+ZSqkOOGvQOpnmgjBHYUjrNHAAXzODqNcpKfKpAzlxv33xhEQu6XyQZ9BhJexBezyB5ZUB
RF+cSx0Hl1Cu4KQKPIMLcWioGqSRSYfYdk65djJTjzi1y0S4AD3jnqZAiQZ4wR6xEAcOAEYozsRV
9YjeQKKwKUyw7A+wOOpF2WZh5i0xogC5ZNpZIswm3l1nti2s2pGMA/nWuR9KQw6BRcXywTYDpddn
Id7gVrziA6BqB6uAgcieACWHWnawxX6iGqlM+WBqKWTdy8AVxl+3OnBIee7ikoB7taeCuDD+gH+k
N9GpIE0GAuTY2jN2UsagKVvlxvcXDvxMXFWP5E0gkchgY89XbrCU1JtPx7B065EPXK1m7kLGynf+
qzdfDjhDJNf4bzxyGzRh8AfDHwgw5aAgpFaXmGZPsreh0Osnf9wt2X64JTbi1O7Om0WGUsWkdK4+
45kz1i7IsaI7DYCc7d1viV/9FyFkoe5BNsq3Lj6diE1qdbFd7JueRl6xgb0hW1VIV0me3E8zasQj
cRJM451sPOyaxJQPRmxJtB/qy/5tBE+gmgzn7Zw6LvQZinD9Ym04QeFgJGMDQ+JYOmAvX0DXVAi0
yIocOKrAhdwxcwLbAjKYF+3fMrovuws5V2rVV1j9/D7ku45DZmXiug40qspqOoZsOLFUfHHHs2f2
knIZekal4W39G0R0UGwWOMyXbAPxbnINW2zcmpGR5hy4ofPRLkIKhXJtUOLQ+GoS3ddJZi5aBRTE
MIS/LwitgNgw9Ma5tt0FSiaq9VShoMSKOFWpvDyrVLhmHbYf3F/OHLa5+4KhPtqmLTYCtniRDXfl
bcxoQOupATiLantg93tMJG7AnzY2at6SKJqkGl9Q1uQ/XUvcmPvbxqI/Bn/NVZnNUVR9Ph1rO+nO
O7ybgcsAh+I6vZI6BjPTUNDM3m0gxTN0wEnH11cekdprP0m8ulzC35WR89PnYz3aYaU0Lf6euSyY
pA1XuqA8ah1rHzzVxaV7/SXBaIXtwy78p3nrdxBCuZtWhNu++k1ymjY7wJQjEMlvPK0d/AL/CTbg
BOhCrY+mfWnWG26TkrGcJK40jK3VAWfGN/+LcJDd+PqcE8c9VO1DoGMSuCOGZn0deNXMP9J2zXUw
64ECPcruZjGlvw/L0+47G2iqc0lUiTaYH6j1Hsjq96Pm6cDlV3Hq3ii/ZPM06ftvsLP65tZSKIOb
mGZnkYtx+A08ayC55mdGZtpDnUqA6J9Uvj0/SW+YSGqYNnsgk3jeI6yTxQHEYfqVdgJuMwRP1K3y
tJAQYyMrHthxFFDfIX+fTY+70NCptorUTgIjZEdaDZFUEf+ZqEMCej3toZrlYqqRibv4k15Uxswq
yOxXd4jSnX5pL0gJbxvsNqKhNq8BnvXwZwFMJYn9KbBSmPoEUPbDoalSSHjr/8YV8Y3Rxq+3F+HK
/L5wHXVDL7NRP4+0WG1NOurpbh2oU7d9lTwn+KbjapmvfnlqiAt1QduGAuPV66LKdg2wgHHo+mmd
sawxeMsog1nwyAWuRR4PlRlY1dieRO8h22NrPTOEw2kaamz6TdORWhG8isCUcxxj7QoJ/5/yEOXn
Heha04PkQ+QoBV7eb7iKxmtpV5/SxxZvoUeGbAQw+R3je1Hl+VqHvndn+JVl6iWhXaHr3CJR7XXd
oNBuX+H3oNATJz8MHSH1TE7rLRb4Q8pFmgzwTT0Ju8i9F5RCRA4sTEr52Q3V/tdExFCFhapP4Zrr
kUthJVbfAx8GMPDo25iMi8NlZdjShOhuaec3kWSJbSYV2ETxWJIR12eKOlpp7wGsXdXz6XJ8PEcj
aoVpHxciHdmT7Chmlhcm12BlmmjGs8mWBVd2/vNZ7kRq7IFX7jIMcjle+RBL75VadmlkE/EOZ+2U
lQlBehZ69BYF/RK8+x9lepa5E2BG0NbYTAlULPFG8FwrVD7Dr8QneBRli5gIB1kWj5yu64balMtz
M0X68IRCb5KqeHOA/prz4cDEa+lOPVvJxWQ8XDEM2tz/Cc2pBqh/uNfAYpvvb68KcIxs2UHtJ1HH
BwvSn6rtd6PG2e4//Pac34kZMpwOj8W0zR6DRXJTE9x2jt4dCRbhiI59n0mlpVdM7erAdR2j7a7W
zHinXODBpaOd62cVv17YU5h2BHYgRKxCEyLFdggNWvUM0SzKf96pdd55lhAo7Yjh/4IqFdtDiWBP
du5+hF7EEvi4264kr96XA1XI5PFnif1NJkJ3FEfLvAnYS8LbOjnfFzcS7Q19Wi6GNfwLrNeQjyZ2
Jsi5xWtOOp+dlEg0poPDlealoRl+yqQ/4jK1c7xOxaM+DoYRyM1/TideqxFLLVi9+KmD14b4jSlU
DXUk1SJwG0TWA7aK57rHVKfEW+i+8KLoAOLHdh1NdTiAlS3naaX+gbht2ArKxutt5cqt/Xesv45Q
LZOM1qvZnzfM/hVe1YTZoN/JNaUEyEg1mmQvycPr28EG3xP+ZbqcxQJfMSK1jJQJsl46vi5+Hyx4
xaul2EZ3JhZf4CrdJf1A/v259R+9V2uLl0f5iUP6WXdGx5n+Vb8meJp478cS4MOXvDLVsGtQkDoJ
zGJ5JcNOdnIWS4RHAaRgpozi74Z7QDp6D6BZq5bNtMjoD+Fy4V/CeF68hDPLJgxbpLAF6y8dV89X
sb5Qwt+N5wDh3r77ric4gWYbktIbyIF+lKrk78+SKDXa/tjOIp5dhi3iney5ntYn/qBnAyR6+USh
1zRVa9auJQvcaIQeYKSUHOvd6PfJfzw9Kl0JzeobfLd3Nu6s+E3Nhqw8juBliGc4obA44oxE6r8O
j72Q6GZh97ZGWpSdLIMXPoeDclBmAKK8roDHPtu+02zzs7NVNFm2HBs/hT6iHjCqLJ4KTz8FkIHc
UMSiwk4A2dfOYoca9jECYxO5Fpg9SaHEMsFP/y6Q5GVbuzisplNeh7kbtUlqfUdZS3jLPB+IjQFx
3kqRJ//pyS3pwVfHxiXP90GPHpcufX96nmzvsRkCH9etJD5pO8XxGQ/J4HuZcMc6gYDrCCHYXFWF
5G2AB3wC18tENz0P74OHyeFrlsC2xC/VQBqazmGsmxZS257tf4oqaRthP0QadtVWf2yMWt2zahFV
GKCeMbn6pMSLAolJEh8qLQqbY0z9jsBeLC1bZg0i160sqYb1PVnwgVQihRpBAMWvjXlkH+UooIA8
8TK7gLgngE0aCe8wnP51BtGRv0lk7ogHvqFFHz9Q1ywPTtO+b7cpEs1WMghrQvnSuB0Pa8+wDCL0
IwBCigXAbsnLzCg1f4+R+2pK3pkxpMY4YBMm77J1WYk7mrx6aZP5ZEFXElu2yqvi1Ge7bmifBPbo
4So0MH7sEJdCDQidEPytdy+x0FVJFEROUgbdAkeqOjYi9oo9NWMJj0Jyi8SF8eGiFy+xXBNEyP04
wdVuRIhi5rBaH1G1FO/RZsCvuhx8U4DcRQnpVjh8wcTPH3aNcU8ewYZsnIls6IaiKWhOYLMBOtS1
E4k1G8AqdfvspP9CoZIznOMCjbhGOwNs7mUcNtW5EE1Ou3eWb+6ZC0WbY+tDFmp7GROcKl3KSUkN
pXWUAIvumqRgSovtz4C6jodEmSb0hgVQmoaMEVksq11GYVmVvXVEZxlItArAZydJYYGMKO/yRP0y
InQAQ2xEJS/3Pma/bhltqS6IsXr+Zmubjoa41j8ldVPS+IAquTCZI04pDgMc5TS0S3i/jN0vHQm7
N3x9GnB/uAhAVpymRalZbvAE21JHyzaGIgxvKBEP7Yk2wZFJYdPGlUImksic7Shsmw0cPWZsxWzl
4AcfiLgDS3mkEMklrrRQ+zR65gr1P2NtG1ePHCzUn4+Vqul8rRu/sTH3d5K2pH3NVoQUrkR1JW5C
HF85+v5YgCp8Qw9aHuye130FwzvdHZP9scTwszcQlGaxioE6vgq9JrwbCixF1abuTgPieooOIpMJ
qInoSdAkymwZZjtoCBoNJr2//poNKobs5/80hRhhFIBiYHBJH6ovVzcaSE2sI0L00AIuOI/OEyHT
9PNbppPo/wgIq3FTLjvi96/gQ1yd1Z3+Wd6w5lykqNANEio0XO3ne4Xx8iAb4imPBP09Cl2P3D+S
36JXao3bNO+uQJMgVOkQkK3fblrMnZ/aWGobJUlSCeE0QLg6QH4TwoTQQjR6X8Lzh0z6zfJETMPY
jd3dmiyPy8BBZnb4L/lNd2lAWpDStK+lmXzU9vJwc9xs+afJMQAdWA1FczcaOdK1ifChCse4Yy0U
KGNrQ05YyekmEHNa1h0o9A7sw6YofyRb1iAMTJ3W0Zf2JaNJbtbQUkcsp3FK2v2fhq/nQDz/RWmZ
Ukc55oTKXflFi5Q07MXNOknvOI/aO+rF/3w7dOuq8UPU9OkzPLvJ8D9lBAYSlnahVQyW45VXxOcI
OeDonXalQRfvPBGGDsw5pO0W+zQKRP/732LLvZ1hXkcmyi/GCH/VYIMUw8vSZUEyMTsZCjCOI22K
XQcTayXITAh4yOwD4uGj/1OCIRQyDndoXtLtNJsbSsfkFs4+OS9VL46OShz99hhQPjKS17ayTTWh
4NwpMK3tw497IDftSpapuDfxuzgOjeEXgeMtHTofERkiyk0cWXhtWQVtkcNYmAyxAwL+BwD0Z3D6
ni6OeWnL3VE6crhe0DDpycOWSjlUalGQlO/dFTF797e17fX23NNnDj0Py73uiXAO+QAfSgaj+P3k
qY44FCVtnAFA91fo6OTiYUfNFy42/O0ZHsKamiolUuSK8Kw/Ja1mirCd3GeX+9aMs8F4fibI6IZN
FTXXQsNBbSW6rEa9ewlnxwl04pZsb5nA7QNZvGyxydpTSaKmwoG1WiIIU88RwH1SrBj72o7AM9HZ
sQk6ZX9U/KEdhBNrF3nJSQqrOHNG+VV1c5jmsoB6Y9VHSVbZpcWd5P6UwzNnzTh2IpUXOQe/3E5b
d+sd05BawpEmWhQy2TS87WV0UzPN+J4De6jWYZwuKhXZaZj9foRGiF4WYyX60q8MJh9MG9uEVzpD
f31IU60o1KF2r9Vh2GLQBxdasGSX3jKqZo/4dZsGe8zrhe9Xheirm2icj+VqVR4BFBWTaLojEMjT
iWimb4mfRFbggZ6LbFn9meqmOSaiFeQWZ7y9OxmE+AaM2N8VoeGr11DzVq/vXqjPZHy/okWy7mZi
RldZVNGfzxz8y+GDpdIlWjk6WmLPP3IpC4aODFx0fMBc3jsUkg0+R8N6Ek8V/kBp/j51bcTagdaE
a8RJOa1inddY72t/aWriTd0Tqp/Xrjw4ujyyNZMsCJ9ae0EwWw8MLtBe7n4i9MBE6l51mBpT6y4Y
IzWkN7e2S74SnKccu+WjwyZih1P2TXbHJrvhRhPBA8HrGMwXAytpUtoGnqG36i9zyd364sgXkbMQ
lO3hbO+ApkI/yjm5KtgeCPqwfaHGd0GQh05OEBYU73/hdh2DYiOXvym181ZFW90ItnHQ+DiV+gsh
hyHVvYjyTDuAZSmQqr527aomqjMMK0+WLZ/wlwxesn/NjftggulnZiCTn3rEBzGbrR7wzZDQInnv
4lXq79qFGHO1Rw6MLsZVzmaB2RZOZx8kbJCqVLphYjnjmb7VcryTUJ0y5pLR5R5t5x7l3TAuJ27h
gk/dZRY2/Beii9GfZPehPFZhs6tYaFaQwODkafmFN0tL3j0QmswQocZblzDO4+UjwIgoMWXcD+Er
UdaPRxKbqeUgn9BeGoFAqSjgD9Kp9XYKUE02mAb6mb2Zs8nnw/65Zz4wODWQOjvNObuti7OaLDwk
kVH0S37Z/bTVD2fNyJp6qO7/nTC5VOwA7uPvItvftvMnUaYGG6FVqFeSiWDtem7WJGtfQLbXrWZE
7XoXPnMmU1jN7PTnjZPBhWMCochXG639Eub8dvp66YIhPUtrGFgaAon1Gpx6ciYldxqM+8X8MS0U
GP5qNqlM5Vfz74ytGfR8EoQJnwOe1kPAGt8BsvrGnrtXjnW6AxUOPY+Q4t/30CMnb26CeFfKvzCE
iSXdg/DEabqMoV+C3gJMWj9ZrupQdOoddA3nMdwHxAA6AoAYvYp84VmbFj9dmHRil8gqJdESJPyz
VJIA3ebGM83lhBm+DDgDeXoJktWTOB4xwV5wYH0X8cafF2FRua5vo/jV2tmdFNPaTdcYnFITOCUQ
tSRu5picCPM+q9BChPpd6/2XZYO59cZpCy6/HOiJSb57YJL4q56hONcYeKS9+yhy6SUv21b06J8e
KkD4m1zWjqvM+7TzQhsRep+0qCRZBgG93ES8725JMND1tByU36JGDWJ6AY+Thvf+vkwH4Efzr43O
NwgXJnWGdEzATHkl3XWWp3TP+bhZTESGdqfJe19qTD8NxlAzT2/OO4LnyWDEhoUnwMQZBW2M2azO
+N2iDuuypxnzhSdNEz2sX/6AyPu8gWiaqhsAjvRpfiW/KuFBbbz/Lu/q5l19LRpNGm6vR4cwU2DG
eGy0yDP0mm7iaC9JsWWMJ9zozLYeUnQ8OwB9MUipi50X6JXM/coM5cpSV57s7TulnBuzGxDXVYDQ
YYuO2Ry4T65jjhRfjmjxISs/lonvNOi8YYsLvGnofu6QEOkYRXi8/ah9Avu5WgoVP/zlkYPoIol4
z6PAGp6DYmJzOYhG2byzeXzo6jI2o06pYmC8QZTDyeLlhevtgCdvO/Pa/TWuwi7JQZZR5AKuiUCu
uOk27xGYN0+vd3VX7AzJhCxw23dP0tG1//N0wbPsi4fcxxKUhvlULHrxdih39GOEFpuHI205Wn5W
NI2D0Xl68AgmwZQ2U8yJUCWJcaeRDl5IsJIGbINyjAFP21eKREAiftCXadU68MvKunywIH8kgg9h
OSB6dlcUZsebd70qIrkmoy1rRvlRBd9fM7cuZp7IMTSWwQ5GMRzPLf23pK5jalzs56zMJLhMnP39
xrCci885TFcxv3rfNHQRV9Q2z813BuVUGw9ARe0A7JG9vY0dyYJj47kkR/IvwgNS+4ltP0K6z4qL
YWQQoKTKd4Oi/Fyjjnug26uNNQSXEENLA/YwnLL80Lu2f7AKxLszFxN4EHUCRPPfv7YiojCBVlQ4
CIJb0DvkQgLtEV/bUHzSBvp4e8twXHD13I9n/SXsdbiBLH5HfMyn16j0nkydgkYSnZU/nKCfeYZn
UsLq0Hx5UUNXS+YHfRg1aEYqwy5KjUvYXhTNZE/S4w6n/bQEKLl4OI9oGnETglJD5qb7j7Wcu8V0
SNIxRE0UKWyftUmWyVcxo0Vtr4m5bDbYQcTLCpfKlI8c8GJ59Pzt18OuM9Bw9VWE+KxIEdmEf7sx
z3naxmUYFDvzs32Zg6TAxOim9qSeg3cCGAE5OxgJVrjbVqK/IA7yXo507Ay+7SPenwx/o0JgEAEY
gSQLWrMUXV/0nRhuzZHLtwNlIhtau7VWnx1zr1L3JuysVB+eirGXemoryBrxVaoW7u3L20bxKcoy
51N0Q0gBKzozG9ABt4YKbNf2W9HEVg5WcWuALy5YvfQmWGI3l4MSrPdKbP09e//P1C1bmzKVK3kA
AddYGttmgmeTyuVKk83598slOSo1EG0Jlwvx3XlhTLKFyp5zkwllAcPv6iVdBn8y4bzjkKiI3ru4
ZnC88Zng4gwvfhe2w1ntWebxtNJAFwovRKO+igNy3kLtr9/OI1EKJGoazzgqgEj65m/7xUqQTx0+
pm8XtQWyd5UJu+vTHKEwg5IX/J2r0QJ0fui1uB5FbkVWr8t97p0NG890BPqX8/LTf1ot5Es8EsqL
O+npn93AuyPNCqaIelHrL1tqji1sI9p/Qz6p1Ev3wO6LNq7pEbYeFfQjeFS4oy573PxDRSGB5dLJ
Km6yz2OIFe82FMhJW3CfL3y+VKuF4UY+kN4jvtsz5ozxH33MSKO9It/jmKaaUJHAhQ9Y38udxiKW
c12pzXRogD+DZ5ANcguFrdDoPcetbANW8lujhRp4wYfw1hb0KmSKrZnHm83fZUqIIYhb0Zo0GAmb
7fdO0DXPABnMBAnXDe5dthK7QZtxyceLCJxV8iejojRFUoGz4Cnz3Yn+nrBoMUPATY2HFKZ+/NjK
unRD8UKjMyaZtEAW2EhW6zUXisZa8v93wpk1dW2waGLL7sRLold9h7nRoGOeTaGd33aoseYDxfCp
kGGZwYPJQfMevPDZgWoX2ctVTJRNitdwuBb9+VpH/T0rwsoVcaAIQdzPK/Ho+ygeRnechJvkA51p
oyq8uKOixvhVry3u/FdLiXhd7FHgCjLlGkNWQoeMnviEDlweUKN8cCCX9sDVYcF/EWlqJXQhUm2g
FBxVcKZU/wV0S3rmIKhVbsKfKxczVAPSmvWW4dkZiXnJQEyvxgCvQVMH3Lg5S+FwNECJ7QSsnP8l
hNESaVMEGQSB5uMlx/Et/vsIs1n3eVzlxMVwFCbDIKEQwkgyRLE/mNhze1sCIdPq/Xm0nEqcroEb
bDbuGUSgbIEvJJIo8RgbGl1bpfj4jrDSxwsA337rVfBD6GCzEIter3jGqksb1gpRmfGA8kOgv7TJ
RA2tRxBNqpnHEZmB+MCHBxjgNylf2O/7sAqJqxFxhQ57EnQW7BHhQ4OSox0cI0X+MFInUz0T2r2H
Jm/fLLFGX2cag5eanUTj/nHIGBgxKcBchLg9gK6uXhHSaH6G3C7UPoGwcIbeG7kGET8J/JrIeNIX
/t65SLwSZrAgU+CbqQQHEtRqkvu64XwOPqTRibOwnwwPV9qEYB4uVITkg+rFxVxdLQollEP2X1aw
RtGfVzID/UerGewxQ805/RMV23Dfh8ikxHEDiAxR2n+lzfbL7/6Lp7YoExZEETj7sIZRg/jKmOjN
G+WPdDDmE5Nzv6fK5Ccwidbcf/YJWmaSiTOvUWiqAfFtjEDQSjtFoMdWH26I0N7IysEHVfONGb2s
v4YBU94dVwbi/AXKCT/J8QW3puESHdNqXS5yXynzzZz+qiV1FzCQid/RtogAZNWYNHDC1Vwr/0jY
iO3UGOTGYuH6jkHP3Xk4WIgPniMJpHzsbKUabPCFyhghfZihV33mNXqN4Yljcqql7qE8I523X6+O
H8x2KkGhaA9St20ogwPBY1XOXMEGWVTDl17/SaMOIpONX+p8HNWX7JGg/PrcE4Pp+xDy0z1hszUV
/FxGQUXjt1AQWLRq8S4G8W/0neTVZcNG116YHdK7jio+0j0wA9ixHq1qiyCS7GPMZHnp51p6q+vz
Zrl6uc3pAqqHGvkU0XFOdOofCqYDRIIJnDTTFOQGX+eQe9cP73agIfDttd2KZYtGZa9JjS2ARP8j
FruTaFt/XvExEBH2MK3BFAcT+PZvXktM2NBZzpRsmkq76cYjTIVDRNhtUPfS8iwqLNCuQINsiwp0
68LIdgw9KPP8yEDb0TUpxNJHR9q756JcKg5YmnyLarHjmZglkJp31SRrdtw0WSaKMLVb6yX1xtWj
2cGhZz45Bu1mWBpuFFaEwV5+QW8y1ErTg8kptk0TeBCzftXJK3QZ8Ylr2z7s9akUn5ReB+x01Wsq
KLOIllk3mpjQX0YskGJxrxlWmAm2Bc3YPOrzDo0cIr72V9r4+RDia9FS+hMPYi7s8/VZIrGeoBaV
uRpB84zpkaex82KTQ36L4vE0aPy1k/Y794bNzM6GkZEFMGQ0N4dU3CIQFEPfdouEmoUmZekXsgvk
kYlmzv3Yu2ZrIuTS43vSn9pH3rHkArqftYCIQH4uWRe4aFHIH1l8fqgDMtIOb6lhBPGSnqPc9tAc
2sHP6rP7eVk68qpneUDdNM4RLmPAz8EeRJfQZ1D+s1S7uA96PPbwezK3F5szukq/axzhXM2fKEG3
ntMzB85IGu3P8uczFupiqHK/rqzEcCMxR9D7nR28mA0MAoLXjD2hQ4fWEsm3vrtzbfY5hZ8JQ82W
+sgB17Rr40VaGY6+UFRGi2CAs0G4WKuutYaqMZChhuyzYxreQ8sT26goyKCt08QE5VJMp0sPUukW
6HezPyrDKoM0aRvuJFPFU69rcKLPJNbqt8RkJtQiU122Uvhbzcdwe8+UhGDtvz2rm2nhX9tVJXW+
mO91ZOBjSqYaPzx5mkgR00yCgtZmAqtKTSqSCrw+qnyRGkdcahbyYDpAprZ2YNERn4K5wx26PoMS
0ycLmUSHADVbvXKgbwck7MAfAJ7wxCIWDeUnf1PhHjRoEzcFnVRHREptrCMosbCEgmYqrrU7P9ot
Dp3Pe8L68wc0NFXXipKEUrGxPFa96SxP1HzozTYleT+pqNNoW1nWL0KuSPXKBFtQ2tuDMOCosm5b
Zm1qSESQ0fn2Ywryhcnv60wwT+r97JY6lFLE9nQpBqDwfXxaFUoA6Y8fClaJR1xb/LY+XnVz0CC5
K+qvXFu/KNq9CKsIyfvjopXn5DRHSChA5m8TxZKaqvKHr18r6OelLsmLA62Q04NyPROVbGZVB6Tu
jV33tcXMZ4z0iyqXLqltfVEFXGc+pwUsyrp1bquCecBbzXXyBrmfcUd3I7/rBNOprmS4JumzRh1F
NGJoxxSL5LAXLNFvomC8rsuEEViHzS3lowQTAD/yjnS7HOMjP9vEnZME/3zU3ulLa1u7migcUL+r
uBNWneUGodDINlpSrziCT1E4BsJhV3rBjqDKk6ixaV1sehLHglMebeianCfoz9Rxaw3nOun4sGYs
ex9SaLEbWgrSI6mlClwB7lntrwBBpjFAyUTWN9lf2ghrTXccaInZVbS/ggW6qaDtcM7v8yPkJRDM
5+1rk6WY27+TtCCqQFs2MMzDTC2N8sIq3RG/4OY5rADvMXzvtOz12XRxvxy/AN8m/xnlMgmRRCK6
ur4LwzaMZro45QGpvs04SmUI88hj4QKiMAE24TeusKVmwrVgB5ToJ3RiVZNT59aBjEyDxSZxamkP
cM4nLdO1+SG3F8W3Lu61WCUuLrLtRE0V9trLf8tNvlEX1s9MBERQDw/b661VQ3SR1MLF2zvOTrzj
2i31hmtjpOHwgr6nxOX25WXZigrE96hDvTQD6nMclm0MF47GJLYXVLA3BUoa3Ag8pqeJrof72Dnm
L+7A8I6/rhohYDZoB6CjSe78zL4TR4eKIM4Z9bqnZRH4rBtid4DWK8tQv8Akg9uBdN2og6t6YE2x
N2eQXcqyTByWJnnWztiJZ95uAdA355FIF76fgsKRRGfWcImU8xOgpXdjEW6lQ9gInDYc4rzU/Sce
i3d4oVlMJzFH5FRxMc7Bo5DG4iQZPC2N+iWm7b5NbhJnTa7Mf/i14wBZzqVWtVgfOZMig2nTspuX
kKBjxg2kwSkLvk4pc9Q8GmU+9rBc+63Gsg3wVHLQz5x7LrblSiBJpVKNl+y6mmZHlVE7mDi8KGzB
RcMDNYxtgJzPYi9xi+JWHFOh9KFYHr5CnjqLYHNphphQygMBpAl1sioSXJwtR/7YP0IJdIU5IFB+
5nCIrZcC9HlObXuDIPrhw6JZSxIfrM+3eJTR3pQTXUGNBH7MuM/UXvd3Votq+lQji+olaUlgtKK4
lTAQ3VJoUQAQsqEGMxYQ8lENUQPKjF/oFwo2rs4E9PAWHquZVQ0UdMoo6SjV/vB4mfob8ouOjqaE
pjdH+uiUqUcK2No5EeWOAfMrA/LjlaYwq7Umikw5KRTzz5xi0bCYUywIAovf82XZxPOEH1J8f0eP
Qvt0yyjujHXniSwOISEPndgfjZvUhdl31qnj21SQpN3qsdSNlYZV8njOy+sdHixaqgyQafDVGmzo
92SNWX+bqP6S6V3sSXERXfuQjN2sX4XocYB+o59qtDRBTp7k0mK/2lJxKnCHmk7sxvLVbMTF8nji
EFQJpyDAYsdBB1m9BT29ePfCo26ErQrEGbVLl90YofrrvrFTS3mQYMpfSN6WP5ebqeipzqx+oZMy
rtfWvhqx1gw212CjOvKJ5Meyc99zS2AccVNqmg6e4xTf2jHZGzAFkcz/cFEfF2rKFofZEFCh1qx1
uZrQYbFbuaqZCnvV7fhLHjBCoyQ/kdvtlXETCRtcEXvT6MPP/Q2h+X2tg3DmWUoLntOoIMoNk3Qi
QJdNw82EXgwaoXQHmkJEZSH+4rFmUpkgZ6p+wNEJNohq/8HbAcIu6eb6hBIf+c+WDWwZrZehvxw2
7Y9wX23I02MslQgiPJpsQyNDuFDfj3fVFIQRtUPHxEHAjOTgNcnWQ0rUyKiEbDoVhDd84NW1xBJc
wSfgSKHfL/9QP/c5xwrED+i/BUME40fd79suU73yBa0JlbkYZmORZE4QX2v04GjYK/ZsVn+DkHpZ
EeNJ0dtMSmJ10tANFyml+oUiGV24GImuLSHMfjSn/wPTfej7YPh3lUnDN8vdaEhY3y+CGJpXmBuq
tGDb7LT1+FeP8FYY7NpPXk0sTIgAdpTWWe6CLtutFicNDaRa6LR9bCpeCBPaRrn8x9NmcwfsuqDw
Q0sNxOdumzYj9hRjfxC3UPojhKpTJMqbTPQwqWDlKZsrtIOnh12Zl8gss5ORvGQNdc7EaoTYAvOk
Uc/lN2e1kXp8qTXK7wCYXOjaoxOTYdqBHp9SlAC2HC+/4FP3P9QVCjNDlt0CgwCDltq5goOOjEnf
auIds+1zflj/LIvcQehFk0/b5A40ZRPwRJCZDVloihOPwL5d6Q9n49fK0bnD/FOKNzff9he+ukqx
jr4lvRDmYmxBY0JXCozBDvj1goLQIxS5EWn9B8rwb455/bEG2J5mjVOOOIhvonAZ8tvWBVEolMsl
lAuI9BDmY3EqYcV2c0OO4mXXyBQ1BF4BrBXRSa8zSqtANNSXfNEsEQEmW7y462lHQ4kRvjwNl2eD
4PXKYwsgYgFxQ5IHntQK/b9plHSrfmhJ2G/ACIkPjpDv0SbY61oIrT5WXPT54KBWGvhZAAkkFs6i
iyXx1MADNohVGXvjdzIW7i4IAWOdg4GI+lzdg0QCIFl+RUvAJRLt0IOr5zDOC4T03qlGxGuCm3Ue
tCeOY4OEzsyRNYKVmhMNfAj1APFlD9umeux6o0hj2yR5Eu7zJOl9NzLVB42ienr4iYNZ0IYQ/G6G
bJK25/M3/OOxyAphGxlcbMPjr6CHUBV23dW2Lrz3NFeZz1NN+Lg7MiEdqTq+FEbEJEFfZZegDCEz
RJnCmg04GGadJZIegCGwtuYGV/gRPXDP+YYYY+6l0ias42cqAgGbOhqgbLx4OAK9hj73R/rJcXlQ
BqSLjYXnxGYSNkdvZRxG99CKRzNzvGAw9e4XrjXXewW+VlAEPBZuJft2MBUVDEsebluqKC2FtuG9
54LIlQLxMRpS0UuvfrZnSqD+hueLVF5RJOq7l1IMRNxyVlQkun8ISGYLNuPfI/Ae8aIHaRiRmhSN
j27Adw9pPJQPb5BL6S3tPi7ZrxJFU7Sf5cTcusEC92R+CFvZ78jpQpoRngVHqqPjGMaXuTYVxJRx
EFItUmFD3tkh4lPQ8FraXscx4EjaNOo5dFWMp7FiLiRZIghx+30luuFdDMTXLVGzCH6TdIOSPcnS
+IBI3XyEJo57Qv2Qy3pbKoYmdiepFIq+41pPdIXk9P0bPkVBh8jmzi3YkZG7LyA6+YoO3YmtPwgm
Crpw5jGlQHAr4ibMkLGk5RrMpl6LRjfHvw1fstRaCMP+1lLeh5INnaiGuS5FIdmlZuS8rc4hi8h/
GX7BJv/m6PtlB78ZQO5GJO1IaLJSvP3Vc3BPO1tPp0b544EdXz/7uu3qw2b59+/hvyOlu1mHyJUS
mjOrWIQK6A2GVjzDo/FdLbotagGSuB1L+8Wtav1fvyMWnVUGmnU7IsfInazTAj9GSaG9q99qKs+o
eq+QYJ8uwM41s+sUuqR32oUF8Tz+5d9Vy/CVkFicD/bBn/vWPJkFkgTNz9X5upaNPTz6RYRwvrDO
2bH4nqO6yYKbbCohAa0AzxY/skauLMbqKdHdGPXLswyJJpGvUl1w6hrZmSyco4vAhCn/TR9/KJRk
hNg8Y6ta27NkjhA7D1jMYXNJzuq51iubPZ8wE9X8azLBQhihFDH7EYP9aajkdpi0IfyljBuF9PoE
HkoIXDTiqBnl3FMBYjpp4NksnyTHvV10rla8io3VFwcYQIECZVduIYmj9nn6hKkkA0K3F1qJiRDi
5+xKFtLUqGk0Rg4umRIY38QUysnbwsqyBJR1hY4Mj3aFp1js+nq479H4TdO6Iafwu0rcnYZ/bwAx
pHuBV+tutxHqsqysxNO5IThe+/XhxArvhDv7rbURj4r3jj7ApninEK22U88eyeqZbTYkH7atiou7
/xxbzhQr5rUiJbujy1L4K4fFy2VS45WlUcRicNGZdjLGmCftk7kNJRVxmzM7Eaj+8KtHEkOhFafa
aKfaJQOLp2JJOYD81+dTlEo/h8ZSe7d7543RCSEFMOtihOdDPTAgY7o0Zdketw2fw8CFmElXCp57
HWPeOj02wAv/MQYejji5tsPCRldNoWf+ZVFwwMrsrWrywBH/4OsUngp/Hic2/4uxKE3wV9aR4UmN
cvnUumAqmBd5eCW27tG5yye+hT+8UqvA8t2yldgIgtbc2apZvN2XeqGAAKK+e8ISrVUA+LTmlp0m
uVdUE3RmnNQ8ObT/+rPFrB/FIucrKX8jdCS9rpZkd3FXzEeLKR0oxc96rC9oxuI5kZ0x7e82F9hj
adRfKqva/v8PrBNlIXuAe/XyTz+idLYHESj9DtsSwSTnEgXJN7YrQytY8DYWgRL0tVkkARzHnP89
JuiqKdcrvTGEQJIHlAWObt+F3m7/OCQ/fmRNM2XTOan/Zch/bortqv4gEVXXIjopofnWotojrWx/
qQTERue7XHoFP+pb+Rv/hO26xAfi/UMrqU7oh60eIXM1Z+Su0jLxqEKlA+7kpm6NXuiQ+Hig/5LP
+JFeKbHXyQglTz1TpnlmS5evVCZN++uLIccBk9j3GxspAR33vi51pOdJuvYjsRQp2pmqZanztEEk
PigMHGshg+09HtAKqHYrrs6GbRLy35a2TAFBnRb1H5bins2kN+uQ9ohyAN5Dc9NqUnbuD6RJ01m2
8xIYGC/7ouX0ydkFsyoHnn/HLuohsuYJKI1BXSoLGo00PdYAqQgbehvZows0Qd4jShwHYzIXlTlQ
DhzVZ/tYlSn10A3Apk1iAEjy+CqI+3W4nSlt0Rlw2rcIswaqpBVQuJwYOpXpItrxEuY5DG+Eyoci
hrZ6YDZb5pM+/Rq3HmrcexNQR0Lx2QcYEkHjBzfvYxseyrglF6dqxeYDkKItYug4vU4UI7vZQ/Wa
PeNyFkEiK5RXd2OVYKCAHcqEnqWFCJpuZxH/FK/cEcZh4VNok8MGwRDQ2w1BbMQwZ2uKmDkYUipA
GdtOxPY4GZsgU1oUyVC910bIVCwSR36CKDtGT7kYfJs7AZOa8GLdba7rdnAOk8OPIVS7BNRgNJeS
X69CrqUXT7Pf8YvIFHXtlMzXs19b2E0e8b/ROltqHv13/39QoV90XkrUlqYFluX0hQa/S7NYcpEu
y6frYR/T4x47sguLnT9UgvWBqFeDytlK/aFVfdBIXUwKcfctrU5V702X+fQYZAmwj34GLPWjzqtT
+o373749LT27eMp6g17oKMDeAJQCWWRyQxCD4jTibiACrHEw7cLw7F2RTvxvxeW9H2CxGAxmCqEo
03Q3sr0J4TTXhVXZLXeDk7DEcHxPn2X1heUG9n/PqjuDU8TR334bR/1nzlR4TMaZffhKe9E0qz9K
L+0X/TPNVUq4b/lDQ1TYAy0eAHDO/DRNExXQXo62gL5jnC/KyfpD1dg9qS+cD3SlN1ZHqXQT6O4k
Xeou6RBaCoiuUVXNDF7T24Y2ZTklEw8x1gtOojPH7h6TXo1rVtV0LcOpLYOVYA8SR48RZZQx30eF
+pxjeODZY01HtZIc3QYXVzy0E5Wf5NP1Ostc+6bMOfu6d27zGfxowhqzL1/zV1lYJDCGdOrPSdtv
TF16FLayjACi9Jbn+AjfBhHZIuN0rucH6N/VTDz8/igaHbogVd2kyAWyGQ2uI5N5j8VF8zx5+KGi
nTLL4OkNkg1Dad3+0G/asmSRwE+poqXGZuGN/qljNPZWKHb9EBIkKVD+XnOQB3SbRok/jk/HCHir
SCgV/ZxqVgOINKpezrj+om0wR3z+xte/AY0m5Ob3Xh4GrmAJFFliPVrxILLL+VhgKN1CuMR1zvhN
Ca1loCmzaAt/jASgX0b/wa4bdZIaQpslGsl5afu4BrkV0MWpuAhkF97nOg+fWdEhbzvCNxFDTAuf
f0KNomJgTj/AuaGyhEJKJRPAp/S/6C2nYbLDEBG8J2YJc/DguI0/029YXig1K2xFKJYzi6d70ECt
9JAiR/hHv0IXkAtk3UvxKUwCbzi4a3vkoW4oJGKMx/t86CFS8YU/fRbCUoNVOGxICVaDbcAHcbyJ
GPZh8wmVXy9+V3iuEarwa57pb4uSplZaARm4zi2lqOzbPyWOZHIDbsoRZJPbWhHfhThzqDSll1Vf
xVb5FT6ekpGupi7GraeO/3vV6Kw/po09ZtOVX2IN1793HvsDpmXq2GhgfCIE5A57R6sllPK8F0vx
cbqzLWglVjTphdBGIV9rrL0k5jKlwoGI/Uc4ZgwaAKFWTncZUO+hmXLp913LWPOzuSXh3AM/A/sB
ntnsMw+jeWprYTNQ50iB5+2WDjSJKwz6vb41SmSposliTUkwizKTjPb+MmPHEsboJbqXgHcSZfrz
QsMwuPsSEMEymldver3x2DwelDHpca7y4UFvBLIURJOxufsKg4RGDWJLrsOO3i6VXIUm4L7XTOdd
ZtzNqhK3EdJ6z/YEvIXFp3d6ZfB6cthm22CCdGCLNpjlFBRJDyQMrmaQ3fF6NvG7Ih+FdctVlrzP
m2oV9qzSetmdyJp0I/xC9FqyD9fY3KqJ/RJW2T8TgiPDQidVxkyaTkx8QT86CX4MzJ4X3LxMoB5N
Ei9GnyVGHOEp1nMung43TK2bFR3r8xSR+bU24ZjkiT94e1O4zomnb99Jr9fdbThTYVU69MO9aQw1
TUUuG8M4UtAPElIgyl0DeOOa+7asL62+/JgICLCnTqebHeZG445FiKJdqnV3cvxlpQyZHXyiInI/
GgiF/6eFXTjvEVEfMw0QNpIpXdNiEAf+/NaDXI64zMQndmIPh2PkDMX9dwsm195g2Y1Li0I1qj77
59uSfemiUOn5go/5tUFYqMTXSwXJRiglWMFOPQCd1lIpLFNP+Qe5TSBOqwND2/sKXFUgcVglOLy3
ugigKVqRmjzai9W14D7gu3Em+H69+99+WEBbrgJzkEwFA7vYq4ToV+XHXUNy/HPWvWzvilux4v/+
52rNmqujaVyJ/Z/g89ZEuG7E+uWO4SG+zdiSV9Thx2Ch1tDgcxygxsHsHdWYaoGtp7QrPL993h5O
0PEHCdzcHQH7E2ZH9BZE8ZiJ7qunSHr4hdKTKtNYkDr2grxvAwGkAxXQh7qm7n1KMpDIbHW5Zc5Z
zU8FHHfPC1PY43y7QlU44TQqn7M/7LtQbhjLizHvUUVQ99QgYTn2r+GF7TNIWuP8RwWh+sMfqp4U
TYKR88u8oCbTBdxdeoC98UyytNZ3tio+GEV2bJ5RKXSuoffNClH+6kThamdrlHprSO5RsV38nawZ
JygnkplUowHBxQ8/IuPoww8vvUmePzZ+LfaTkO4TO/rNrT4Qbs5W6oZwUjyhYh9AgEA5SddM5NL8
BgndG7QyJtJrD+a39Pdq2n0akMOvQ26/KwXl2Fmudj3R0ZUmIfJncR3EjCzEItMGwggEBadNcq6a
9SzVAbWkmxtegMKQ+i2Ptjpcv9ysg/Hum2BPlNwwBtxV6M6nYzuUitb9l6V8UjijmfrQ4JjDi0Z7
QEmwcmuPryRnUhDoRW0lm1R8X3MNtJ4M/rRY0WwXVtQqakJD2kHtvEsps7AZN1WdEO2q3jNITr9q
rR4f6XKVDUg20pjUrMJG9NYExlmyWH30p1JNi4l9jwZUFrQo98iCqBKfpHJDZCx2ccGRoIIfBKVb
wncMmmi97iiD0XARbnzVynYb5jBi5pT1ZOmg0SB+ouaRJIrxDUWVbTnJV3COWYKRuvDPsmhaCvPb
xZbdN9rbyQca63zRsoOcWDIqyAU5eDfD40w79hEaB4+vZYTyeI72+t58Z0+LBa1YYCbCYGqxmUpp
kxMTc3F4nb0ddFCUM0Vy3CxFa1qxHNp3U8piBAcX8U/pE+ccMeCdSTp9565RlYM441sjiH0qHyY4
E+u1KFw0n1mzSTleyvlLdk4++2iX5da6c5U0UCOeicswFNVy5Bs5dahxJN4ScKTxazL1fN4RXZ8K
x8slMMDnt7ORVBOhflHMDsXrCpo+hTUulxu7VNogBO2FHfDK2MLpbRkhPcEFmdYJ3XJ4yBB2JcSf
nZxjobOUfbgBQNNj3HFQ/2zPqza3QzQ81tqZ8mC8F4/HPehyUMwUCYvNmSXxg6nYY4ZRx/NZ9cJo
5V4rnuj4g84yRYu0Y6QPiU0b5n+nbEZ17o56VIhlklrLc5twf+rgYifOIFNFX3cNdNq4OV0SLqij
/Chl57b/DUhxUCNJJFFZd6710Zi5KM3k+YGV26FhYnK0/Ry3gPqxooEEbj+dK98cGvLDeHCdUk51
FR31/EUumi15Z+qQcRNCBisCWp1uf/Iraa+akd/4xmllThdsWmBt8vNkX1S0cGK5wHBJEf1olX85
IZwAFDQfNh3q85tN882HBme4UJrXx81SZB4GAapONefGkShP2PoKubO1oHtCvj0MxYfC5pZuiK7g
kk63HBTWfQfUxCSQ9w96jk55dZ8cuKwW35NQxeH7Xa4tE+htM4PS7JWgIyVDxclKkrGk7EvEzPZd
SWyzeX4/zOaX1EYn7XCEcEsqkNS/A9rcfEFhYZJZiBYdBDvCsHv65T8+q9azYwNB4yRcsrcrknH0
EOhEv6mINLhBNJGxybuCGwF3PQThr/ER8S9hxGevpyw9VODv1S4QfL3j6Hpo2mKlZtsrWby4u72J
7Nch1x5+ppVOwyOTPRz6uNuCCZ84pc7K/qd5p3Gs8UFLidwQaKKOx2LSaIXWbuLcCa0/E9drevIH
nqJkDK4JYaB4POvOlJOyorqg5ytsK1gYQAp4mHH/kk6mYKYOcKjKGGJ3PiRxOUAESy0/YS3KHyEQ
dQBZaqXvDCNNSRv0jCnYJXu1ihGAquhySD3aQsh3omZ4jCBTSHnChDdynWVd4yxQMAHgn8B2PzVH
prg4qLjT3kLnApVi0Mg3ky+0wFUDpubjHsS7JkNFVA0AXq7HElMoxeBz7Tm5SVqXCMB5DpcJgfDi
XlmtGdXDwdo7NnPWQfxcJJtp5FRekMC6stD3dmt3LqoqAOQpwq7dwBU7cXeIvS/eFwEfXOMhYtpW
dhGBHxLK4ckLk/GJ+0+FwivElbWrxbZzEbOXc71INoxcmGsCzUoQw6rTLHibqVMZp7P8YgYcEG0O
9dLBLj4mHjD9qKTqUpjiB6LECKIVP0TlRjo9HzSIxGp6B0FKDn6HNbbhHQsO4D7/aefXcE0sHPM0
21+nO1xwsdjvEJyQWvgrY+a0+lwM1mnnCMj/keEwiDzUw3yiA1SJzGkPmHgeGg8Bxremi0Lsk7aK
kQO5sjNb0C3MOTIqb8bV2CeChse/ahrXsURHPfK3ltkcXmz1PRkGofAIf8ehuFyskyAgjsM8tn9o
KufmRQaQ+SGdXMCZ0L1ExW1oF9FAkuNBmcirHrxxDwHU9otZRgHsU3nRwOxC0EfULJIQG8/c8U6H
19MXzZqHwDdELo3AgP5VcaeVkbHOZ1dUCvg1Y16rPPHDd7DW8HcWSljb2YHLHme9IqboWnkHAj53
V+BjLdyTn+2nChGJej5LjcGO6B2XW6DzWhTspW+lC4QJjppUqd1SKd/MF/Y683/o0sNE+C29Dge2
b9NvsdPte5ix+uW82avTRPv47+XokhFtc6tTF41aaD2NIg7pELi6OdLdRbxmFM2hNvdGqUuiKNB4
tV0wS0gquXsaXOPGrs7gGA/xxzAOHjyiWCCWnvUpMW2JBEMnpu3kxK3AZq9dl/h+uKh2uVDDFaIa
SjYwms7bw7swjYa1sE4NnMCQV9tmNiK8P2bg3qOG0WiEphHisBIsAeE+dRNvhdJBEWXTsRYvFa/A
sOyrbhxKPbM0Uc8aRGCGf6SWmZV8K7ScyYpPvYH4+tuY6KMfrceUXV01yrzSV+qnWNmdGNg8FPel
W+jgImeJo4gqiA3T/dfquRVIeFg8eJcdGPzcHaATLFHTyyWQfeABbeV1kyHRZxVl+1zc7wuVj1iN
xHzoH5HU2gewHm4PVnamMgURnQdZCzTHIQXBsW7NMbWwyTJg67TJ+u3AFXyDrSQvWjNOTSRv8oph
nnw4tYc5H5eXScHi1pobFqNn88q6lURk0dZqmqs4Fj4hOayOxgcz/GjSKD7k0qHWhHN54kG1Zxm3
nspEPLxOIHD5kFfyhnpE6D6rUi9sDBg3c4B1qvbMFQsLmKZxu8Y75jsGvv3ELLRCv+t0lc+8Rb92
Ji7ZCwJGC0BbHsbBdG+tzF4mhPi/4skT9Vqgey5lh37S62IuegMyCJrcJFj4qUyWm/sask3TvWJM
im4fyxqbqvyiWun+zS1rwXSMqcnDKwtWPKzdOGr/SqGO5jqzOr/7GCGnaBTnpWuqp0ZkxCuj5hCs
HTIvuX2kg7T4gMQouJ3JShcXN/z7X753ac7huqpY85hbcKS44c/UWDuzjFUe6UIA6CVTdnf+gQJW
DiyQsHdj+OAlkwfApq9VqTZ6SDytnB/Q6CrRLOd8BvYbumIk4UyA+gwmGUdX1fucGKOp1ropSJNw
KpdPG9Zuin33ocgKEEi5WI64+Z3Qf3SI6XWoaaddINx9Bn0SoZu3+jYVyKlm64hdPUP81gDskiyT
iBLQbV+fUHgOWMgrsGLZ22OjXFWMAOhxBsXAqFQw3mUVwI180opHtK833BYSly3xEvA1QpMpC0Tv
c665q13J/49lXx2c1VQbBeQ0jgRsHLWYp4OsZRiLqEkDNy8PcjyUfyVYFGIZmvCbIL1xQ08GiWmM
21DxgE015of7bScaohr2c3k3NbCMp+4Bu7jDhn/0td5w9r4SLNR3CFS1nQM+48C41TctuNZ7blW2
RqRhSm6WRKTTdaj+xkD9dZZn90MDcLz21prm5Yg6s/53wgh7wa0uLCQiWyHO1iepymN0GQCE9YER
GcrTC34ese3K2up6YZyzIx3p00ZO58+cnF6M+ipR1/4Semx3oA4mC319MbRaK0zUKhJxwFDDTyqs
2FUkddwpsoVsVVGlBnUKkEl+2OyahphlSFbQK+mzLkJ2XoQcvM/fDEJgAk7CziUkDRXUpS5Cs08Q
0YT6AevYpeAz6LpGcnpMHWAdnYXItI4qqn7pS8vIOCTXi4YxGyu2FWnXWAU1iJyj6xPo69eC9FFC
bO8Su+8lVDIxLsA354kIUxySVCxLf/XmliiwDbMw7u2Pkz1GromciwBtoa5nX13YWUB6+WZqcS4Q
DVJ6QtvlQ+NiFijfuYzHp1qXAwJ4xpX5jcmrbiQIoNEHqKyazt/v+LWGOIPSzqu4oMLEtUEjoMFb
AHl37jyvg/NZVhCcBP4maPdzslp1mTDZ8HCqmeWnhKUrKZqIo71BTOeKx1dyOC6XBUb02EZK1AV1
4deJN4+o2HgrXeT3LETWEA4XRuUltm+C8rWVo30kfELLM41nBpB874uwUF4yAnTUOGkdQ5eZeRhK
XJ1/8zgLKLb8okmGVcE1p32kSLflKI5qawJBSgj8ggEmS7TroTF+H3kdiGfDT2JhXdOqh5pEV//s
sXinquMy9hwFXpxapnbw+tWh3n99h1qUpVi/hBu43cSjUvSlfpfHFdUDLO/j/dGH92yWRdTF3E7F
eyVSUUSlV3FB7NjwicS7+5BhChGAT6M30yiD+tCCLKXKrDF//ykhi4YhOZxjgGEvz2xQxTArvBOr
uISH+t/8lwO1CvYyeO/OGyPE6tdimQT3YsJTHATHv4rxByoFqJ/HIPZn3TmE0p0eBoMaJLezx+Qm
VK8jkJLYbWqiWU6wbv3d32jofqUBqC+UJ6BDoO4kENi0CGSey314jLM000QSqCPyN1QHieDJxSVj
Hh5Z0OvoJaf1crHANG6dSwLwvhKnQQiETVM6W6nvw0IDCFbzCmDF6zDj8lp4S4j0DZ4pO36urA7i
hved0+9vgWJ/IWcoNINVmI1nj800XWSM6BTLiOXIFobnIPJgRnWbWcBQe9cnkON5ctqzcHpRfc7f
jaMzAKTfkEiG0eYrY89SeWUH8lEt4Em9CN76CV5spvwR7L5fzBjTnIE9ZLOQ4KzIilcpl/To+vBW
OGqPD0jEAPQqYHsBVDyCHwcd6St9e/xIVDsq1HVXVk3+uKjNd+/Xxl72GPfmSsNhi2QIOmZE8w8g
cWEQMjgXxl7FcLMxpiXYB2Jafk6IlIeuyJnYiL4FGTUKariX7FypQkErAQ5r+vg0w91ym5a6gkG0
PShyMZDmfEtRz2dpa1huYMNLspIxB+M9Idn8A2Fgo61cr4bmjH12kDUPAkKMr2nKIBWqgGX6ZGvj
batqeKtoPo72Sya//NRetVToNSAtIZRi4DucZbcUO5Ib5OyMFaTCLwgeEzScDaDXXeuY8i7hH1+V
kA7LCsA9dLpXdLdqMKXytOdtzZ7PIylweQrsyu7drObIsnqZ9LBu2e7F6HcFFhvryfBROriDZW3v
8Z78KCuuxnv/VuWzR4nrK1EYGwn8wf0sNWUosk8IbTILdcYKrNKMzh4AVzBqy8CVfEwgbvpBSfEw
9B3kQ8G43GyQqRx15tbBs22DpaaIqQv1DBtEVp5MHgSkeVa0rpniPo5fsAozCYWRQCx2RsHpan0N
spI3/L6sujhKT2gcdt2+TUvLDKjKbK37zEN5quT1c38tov7R4bA6JuKzNJsRCvVHETn3+Y/4vd7v
ULuxNirB3IzpSd1UA5du9IOsBygvtrLpk08cLev+GRAGiqY8P+PMKpGk2QJqUzrHVkI7X/k9EaSo
52uAw71jbGVM6BwOFGdPr48AXoDKYjVmDU8KZaGnKGdwOCb9eQsRyQmYJLYaa254l/eePIWx8RJl
kccS1wgfMKluuPDPYTeN9UGu2/BqMwefPW/J6l0CBHyEAOa4oTSlx19OlEMN7DUv4QQ4Fitaj9UD
kNLwWVUK4Q6IgOBnzaFSdlxUaXhyxyQ46XevJ7kFlpXZuJ0NF2+od3i4306eVsQIo+KROFHHh0FH
o23KHFMZG8LM0NdmhDJVUNOwKnL+SnkLWAuP0wiiKC6PnOfxUJdW2b5BfXcshbXQbH/08LimBlkU
5TL11NWqM71lx7Ez7/CmnKeiulEOxDGkphfT3GWoFmUvWSYuVxxuyKO8bdOxTENVnz9ou90ZtY2r
dx1lq+sOSdsDMjD5j+w79J1yPnCUe2DtZeFS0D3xSIWrP6yz6+IFwX/k1ORB/K24fAbCsNjOn2o4
5aslirjH4VI+ESXqBwZWnxIMwmfF9brdh3c1ctHyBDQRPe3hdaCXEanx7bYOQpyEkK5f0X4x6Nuo
NRs+uI646K1F8qo6y8G9UZB0FxfmXK9lE4n+9X9OoE5znbvaaP7N3peix1M1ontpJ5FJgIcwV/+r
9R5zjNESFv2JNfCvklvxzAjx5/7gDgbkOmjoWJKvivVhZbHTTT3Yy8fTlyAPOk+vu7hLPjjWRjKM
EOkRy4Ed+r0zVgobyo2cAXNlyMQtvrzfEy1xExzv3BXvEZmKUxL99NY/DkHO1C1XL6Jvu+zFS3Uz
EFUtq9v+SpFmBjVSBzN4qWnHNUlLpDOWsEm/GvlBq2HDBKNDwnuvw8NqyeyHxdGIGEXxjcswyMvP
Vh4hCeSVuzUNXdiXMJnML9RzD/i9yCfR8oZNYJm45TqZ+Mxj+Qitgat6hPRtjjGpjSBc3AbUhkLB
zEivpYVOF8HaHFLuivBzyhNxNIIx9QM+0N82TUH4dmXKCQRr8NwE9wc8bBPStQ4+7Dy29tQs6BOJ
y/ytBKaKdLNNVG5qW+44VM41b0/enS3jCQjMwe3Su8U12gFjB5u7/eHbMil1lgAuU7Vq5u2qiXq0
20k9aFgGosiUBvI4dLrykP5jf34kMt+CWTHOizIIhQxj1qbDWV0ejd4cj//q2K0a6EqBzc6XgfJi
Eh5W31c2bQukTKdd3BxKkoKELPw+wH2P1KWruk1C0XMqSl2T+AKozRKKb5Tmwb2ZUeoy3fyZMO6z
B5thBINEq6Ei8V7ViePm7k/u0TTtf1bA8/p0m9qIeaARjf5JcUlmd9QhVtbfukS+80J7DU6U96ZS
9TEvOKp7aoQVCdKpOwUpFchYNYxX0ppW5MYxHyW45T6CZh+TVh3UunF5uGF+OFnSjsDAhKSWssoi
hOzboeeCvoXbRFW2cyS6D9XvGfcW22qy5MiTaAhQlaDebx+6RNApybU8Vk7CpDC6fIkqh1nYc5Fl
ZITQyBXWOk8tSwJZDe2tZKRaBegL3MvRfVNOLP+Vz51HIGjivK2EHwsf1uYZ3EK77mr5dEgO0o9S
Nsk9Z6bxW/2fy9DmWxlKLY2iX4toDYoU8awE7wOuXRbf4orYfiLaq2/ODhSWdj3o29ddNdUmYnbZ
u0mfP5YPkLK16FfjA8vi2ir2/fosJbxD5Ok2UAJUjpAnWisD+NeqWsBA9pux0AsvgvaaF80WISh5
TFnKxoerWACHO675EnZdokpSy0pEm0AYgCj34Q1OuXpmLOwW7AiKtTu3UoKGTJeAyCqbp6Iu6it+
TfCEqecWWGW8JT8EYVoFYNK36X56KKiNmzoKKp882YDTmXdOZ49N/HYlC4iFhQPvlEoACt0sbUEN
0576HVH7gygSxIPsxIb6uEud8vIQLkGbHIXTTB846dVjt6r2IfICvHXY4sNaVP1nDyvJmXbQYKYD
VJg+u3RUpXwZ3suW+9Q0ibR+E5BNcZ8hPAaClSX5KqzHUFFmj7cJWRSZ4HzWbVETb91ybYTOeduz
jN25wOe5+VTZZ4RtJ5e0V3P0+22f3WHjs8GT29DIAr/cwY8FsCEIGglon6G4BG5qKmNZs7MLlw5A
ubq1XQrhMhIYh01QIm+d2PrRqPbnw+514QXL1t5acd0vFZkI4tW16KVPSyftGeVuntKmKAuZGfsl
nJTnnT+oOnBOIYa3qDsQX+cib7AH9PWeAZRMxM7sIgXC/qJzgxFBWZSN5tyMUmx8qkD8lfnRwGEc
WNFcC1gBeDefMMnCBjKmKwpvggNIijvp4J3bH1nA4nbmiaAecYlBi5SAOygRdNpedXrIVXn7fG5g
D9OsgltlJ5s18xRvwyI4T6o15sghzpBJXrDkPKoLFRnoykrkB9aDxXvmiGiuTcSSqXNoPLf0Gutm
98x+Zskofb9lVOynnMha9XRxAMV/+puIL0x8aG8tlmNnePWYefiogUI/Z5rNAP7QGf7zmgAmJd/Y
UnZGi0qMLgrWDtOVp390hBIOyQSR3ey36GmvLmcPcNe/bK4uQX3nelijRg8YbxYUz1oO6WB5PajY
sUscBffps2jSK4L12fD/bq/fZ+s5ZupqvIpp9SPUY9A0qjHdGJqVPaTlt1g3DhYR242QMsXVmgLL
ZCNrpbtLpwo9jsZhPMactpmpTmQPMNSbpPf/opwZalyfCAtDSWAA5gLlJmwmb4mmws+H/2HH4TWS
KlywwGDhOVrFJucHZ6CPkWQAYJ7LD9XEf8+UXw7+Uz31zAkc2mb1V0PL8xCSI5GMebf84o4K+nqi
WpCaUpZcmbJ+0e1DakU3jBw5zdqvfchYMcTG467tDHsXOuI3VinsCdYD0SXJ6Ldm65695rqoo1T2
4tP88iJusr4hndgfilVovadXkRxu1TDMgVDXy2dIK9+s2hYeOeEkTZAJ6XJj+lF1Ne3UbNSRd7rm
iAMfubwxii55y9FN0h6VudghrgJfJdqfWTXzqTOTv4PuY67+f16pjNSYof5r+kgMlCYT/aH7FkQt
AOyaDkS/SihBqKTn6pUL1aVfv1vLynu91CbqJRWczZm1pouq42yIkIULQtJ40s5gYRLUVioBaVjg
RENt/Muo1SZUz6dxXGzemYm3QlOvxZxG3fMwEmpU3fNfEgQhYnTXcvDQvKOFmOO32wC0o0s0Yo++
TLqZVjuPZzYxIOMYe0tsGz33dil7VDDp5ZQTuZs+oesjz5+XgQ3H4IodE7gGC2IjvkwzNbEcrHPm
CCOpVAFWXvxNuYKiYYGh5fcS1/ZkMpitCoiYJAu+VBohsfFtyYuvHKMt0gv4QNY8Y1ZCDNbq0iqj
ezBF24ew8boQUvfqWtkCKzmmnJiVwq6a6TRwEdCIDZa4PnSBeDoXoKt5hzHkRA89m+xzHQPXrq0S
0hdLf5axeCvJUgNv7wKgwzinw2BJYM62MY2wxucK/lWro+5orjNPaySm1aG5+KM5AFbBW5l/rbc4
oJV1AJrr+NMRLPk+1icmTIcHZd6vzdZsrViKwrs8+dF8ejg96OZLVo89KGHYkLls7LXLmO4+kmrZ
4gNjJDeDbff7nMSH2X8GLBtyP8uqEzEQ7r4ztn0ze2R5CsdK7pzL033VfGzmmaw0+oYV5NxqZmp7
dGMi8Ol3+3OSa9AooYQ65+dZInhZU2fM0ZMe2ObEh7Izq8Rmxr+i3qPahMT4YDaT+Y81+fpoQIS3
wjGjutmcT3atFp2sVwJi31MqGcqksCMtPALG6OqVOeopxQn3q0n7yiTwCUuVLeSSQARvCwVJFpWj
g+RhJOn+PiAp8d+jEDbk+iodMjqDQ9DWvRZjkukS3fkkdPTI0lbRvLJMQHi3ldnaiiDgIMeAZ3DN
KUpWx+nSTIb4eHd4rdwoTS0Du0bTjTm2RYlwF/+T2GO7mK4QOHfZggwEZdeUGakWYNQ63ouJKgCS
FVUAjOY2s+fzjBKbV5PcfqJD7FSQjaXMyHkTZlRK+ejCvR0taqqemRnNHtSjG7h2h6Wza8nAsN/Z
jMr23wzhCY8JHFWSBTWQem2twopIPD0V2+l2gKEhYr6IhMg4Ui02neDFymVSW+I6fdDn9O46hJ8T
Rc3saDH20NO3k9sOUDImv35EUwZDE5zo7FwotXs0imX1qoilEBbxIrgPQuwncVpIQoOFdxXCjUz/
aDa7p00XqFp2FsRSCT8WRZ54yqt6YpW287/q4WfZ8VNcVGNHrv4M4Fip40etWUE8GlN4OgFTyAp8
yZ0xxU00P/mVu84XpaNVqnZEBXu6eS6+qU9mx+P03qYK9nKhsVU9qX6SRyf3xHuGr02pXyxgdKnD
Fm4BUpwoko5xqydmrgK+wS15lBgRRa0tgsZH8zTLqEd+k9ZUS4JBmThjhwYWv5EJ5Dr4wORg+K8g
oQCZx7QicvlpR/8bLb7Dp/ubOe86AKtNdXdUkLyiKZBVsrxFdLhTI8lY1l4ZC19EgzL9aQ7KouVf
P2f0G++wvfVsrie9r6np8Yn3ry5j7RRA7TCh6b8IG70gJXnKn4BnOtoi+D9QYEbP0VxGUs+EJHq+
UKxOqXgr0Qjol/ueXf9KbK53Yc5n7orPRy5sbzrjIP7YrJDOvpptPbz8A+3ZMA0H7pn11PtrKnCy
UZn0sC6e8+TY1InNLM16UAYI/AvpYIKQiAz32IW2BoIrZ4eqM/cjeg4eBGIru8cZif9K79yovbBj
X8umXFG4lpMtsJeEn6x3NY6Ub9R6EbEq16Mrp31ZxHTN+qB3FkTx1J5t4we2UyxrDfV0TNSOOJBi
WaXmuMejzkzEBt7ziAzjtbDxDCdY9ILS+zDnDpLDLdYqzZq5/BZ2blvkcSeuKp7+6Am76ebIapca
auh+mbLmXHfKZu5W0iAyG+9U5wSlC7AcAUCsnrbSGiH1Ro4rld379HCQa71afrowPoVkL16K+tIa
fi3ZIqwosW5i2EQMBMDCY/ZrOgECh++5mwY34HWVG0Of1JDxgvu1Oz5WrINHqHr+B8BPibIFR9sH
sASD2ueL7oY64QSB7DjWlkhPWh5qGuG7PZlXcPhFGZ6z8L7Q/g5iLCSPwBXBLq0zByXBzA+7qQgy
ONDvcDSvIXIypvSe0VSXcLTxGZtAZy2BI2B4cWkSetQJGDA+CWAc5GA+ZFXOrxj6IzE6SH+R2jcp
bHPJdNNiBN1f/uhoCmBfY+1haqA2Qz13lJalxVcVq7EIzc8NyYhnWowWF7gvedaek/upgsmkRv7u
OX8zouvjlL4jugQwDQcIyO/c7qK/uh5tNQ/zyikr/H0PT6yVabsoRHxg3D+jGcki7cVmbhq2nBva
GVCFGhz5PV8hPQ7dmBPqPXU8BvS74LYX9RI55yczFdGWSVDOyoNzBwFpaGztUzWtGPEGjKhXdeqi
5P3xQYMQpNPd5BYDMAK2GFlvYVcNEqZfZ4HYIV4gHSolmWI2S5S+Oo3x3klEjutj2xIp6kQAda4A
HScIOgzbV3Ai5qeg3K8yuDB7WwslonMHMG6eaOTd4bK33J4Pv0jqlhnfdPvl/srkB4EIk/kwFAWW
/jhP7LfKo7Q16rixYjxxAtAgtmp5tpobRvn29xTRN737rv4YjeNAtejG4YpugRn52Tk+rKCNWs7x
CFtHwmfQU/eC3MjjkXZcCr1v4ItH9F4+y/tCdIfcRAiBFPcevEVo1An6liuRBNPDgEBUrPVyj49M
qbVOJcrlUY1DV36ZvYWphbkGJU1PVs6+w9Gl5Dwrta/6KqWdC22IfuSGVkgMq8TqvmLtd8Bm1nPL
IA93OWLKQLuRYkAMVbraG7DEB37AxAgoic4WdK7vtPT4tVnvlLHvUx4jqQ+s+wGWm9rYPouNza6W
3SLleTeLUliuAfW61XPscycmdQ3y0bTOoofy04FGKocsEYKoFu+TG/mFMA3ulwjQvsV5gl+inXNJ
u44RaHRs/kiAA0+6lxjy0RHMM92O12+WdvifJDhWKRHWE+NDyEj/5gocXzchTxlI7gyFLGTtEStY
6e28QickpYCtudItVNpH0JX0fAwsHqMtbFMawV7Ja5xEkm2i6S9Kprza9tlLlNN/CpGnuDBg7OGx
hupPKwNER77tDxgwyZq6BVaz62XqL++P6z5vPf7tPMDKSXrFe2wLqSJJ+ceg/ByGgaNeowFwuRNB
aOuLb8PGCoTaXYV+UGO4ahcQEh81IOR8nN0cKQP86p9B3frlYGpCzvKm7pqRAfxWuY/9HVj/sra7
Nq5cADUX89H8gyL9Okt90pnJSzZLy7DCfJm/89WdBIlHt2RJCdXA5qFR4ZGgqgaaLX8O5Zfc+6Kt
w/Eb8Nnyv8qL0By7fG6jkDwhoOp1qpvjJqunmMPLrtKZdDC3FLujavWLjYduH41IvIQDyQs6Q5AW
4EkX2hnweAFHoPc//Is20y+xaKNPXUfyEC7R18ow7fzH4xmH+jitqgqcVfri4H5t7KKbbbSvcwqm
GJDUAsBqyeQ0YxkBLKNORNFKkjG7uAGQdjU3tRcw9Ivm+zKbzasoChKFClMCj+g4MmycUu4SFHjd
MNU4hWwiCo5U8cAvcj91Fz+9yQtVTsni5aEtY59TyzKQczvUFhGNv0BivprPcJARDioyj4gvJxRL
moOHNfO2ckOIcx69ud/raKHbi4RhJMMCf6UnPR5rYaH9/04SRSEKiVsw95Qp6Q250MdkWDnUBtMM
rnId8dH4IhG+b8raSmjZzVMp3qfYYJ9c3tlTqPPkux8E/MGQz+3WomfWyTHo+vjha7tb10EWBz6I
JbpTf59ESIDv4k7NdZnVJwQI7dVfPaPRdNCJegQQxYR33Fd+q34frjp9xla4fRSFWeX6334SA6mJ
CkDhzvlyoPds7jUuWpz4qpZq7f6YJDAKoRQjG83xaEcPQeVhKtDGApCyiMTEEUFww1AvN9cBa4RJ
INnI1jxbXxs+D1aqY7KwD6ggUVhpn8OcJcTvHGq9GElaz1fW5vC1RYKmciBPxbIj8zlJ6SzEeAt3
SWljGVs+jivljIaiTnX7zMdL6qbTlI8Crs7BO56t72Ao8b3ZNTlLhiISMMZqE49Uyj6BQ6y1J76L
smZ4roN4LwPDGQaGE+ezC+hEpRdrfxL1o002X9RzetK/ySDXXp3nqdlWkolK0W4jq6Cj+otvsJHy
lmhJEc+Fxto4kr0x8kp+l4sjbFTS8ppkHuz4X4HSuRscCgVJLi/N1yPWozZs0+oeLBNhFBcS/2rp
a9h1IHVF+NvqdY82KgjmBDXfbH8a1qIEPoKHmG6UZctJQFGptu2ywcHKKcFgkKvKgvarR5FE7qJf
lmauDiUWd3/QIy9TESCbjYqeR9Vl2+AyRocFBy+eRf34Ym9F4j63X7sGn54AHj9WdI25DlAXyz+G
WAfgp/Je687/vn9x6yb2NREkiIpOM4sZc2aBEhqrKtAdXxI2WVLq3Jewam0JGkC2nd4WqV6e7xU9
XG7Hq6OwWbFFEu71SwErm5uTRez9VI9vyK9BWd/Xds6Y1yJHn/v72n8G/Eks7EVmwCeZpYysVWH8
NJbktw8upqlOVupbrMBSSkWsLVnGzzEp+QGyJWgXKivVZ/AqQwe8QUQH+csGYBaEyQribvObw0I0
1itVe9xXwoX7fKMog0+g1xlontXoNd2tnu7/1GZ8cdembUfCNW5lWYOy9tlrxP2HvBqE80mCKITu
L5DtULF/w22vjIi9Za8Y6RpeeKFd4Cwiyb8y8aYotD/qczfP764o9JHYt65ZO6X+dESqQ3DFSjRB
rh+Acg+gM/2pZATkyhCKncK4PS/A6sgg5O3xX9TN+jmEQrMeUJKz/KsMozJSWtG+a+A4HRc5lkv7
P5EdBeVLsPVd9FNqAg19ztXmF1xSTF2eY4iyeyp1sgMMC6OsXszshKpOr4T75PfM1TQBk2ol+j6F
u2ySIWEHrdQf2QWM3Mn+d+YfXjDN6tK+nG3b6311M6WSmnDNrLZmk19Ii/w7JjROmcY/zxmuuxDk
irHWCfYQZ+TJwIPz7oVVJR8VTpAW/B4X3PfLeWSdCV9cmgTFTRSNcFgZxDcC38TC15Nf5RsQwLrl
3Pw+C5DkoxJWPzZDlynu79PnPoEHsYyNXHyW1X2+P0ie2iGF3ZfBNSchY9wovMTAJT7VQ5sVHIu1
XyoptNx5kZDgoEpCAE3JZvTS+tzJEP0Qusx9c6Mwf0uzatPsMpxtq9gre+gnoaAvfHKYo5yyVeE0
+cpb9j/L4MwYypB2voCJ7+ARImUZeF1k/FAmZ2++mV0ru66R3rbHcV48eVYCoQLF0qMVLcfdmPWc
PWHwFxR0qR8Kzwq0TvdsWbpFm583qaFi2PDPSIXJJ/uKV/I0R5ruVtu63RJ2sUUMOwlrFunpiVly
qDcm6mfnH93hg16AFB5fUWEK5fcMowk1pcp5bdSPzwnypX9S/Rcu4r4Uy//rfutVe7j2CT93IGnD
iW+8Ko1EEZEWYagc6FVNBwGTr4vCm4R9HlCacFC5ZRdgEJBmOfj/DQlOE7wAtyLYN2pd2JxgYjlv
4D6ifPjFCgy2DShcdoA4LdKwFgxU6+LFyBNJmin+RrXDkcYZAA1N+O35/CDXEx+yRG/iLbClyate
vzPEO7WLxiopnN2tcIFSmlkIjBqfucOT1sUaW2If7hFTlatJntT7atKJttMUscNBOjSR/Z4c01rn
2CwkmqhPbg92v5gt0+l23ToiPj3jT/P3KK+debR+ZJuKUa9Q3qozeil9aEzDaYorfkB6LAIKzzTP
I0JIrqkZ26mktIMMAKyGFASPbBuH/W8agDrr3z9wZHJdqi7qaX4PkaHivlk2RBcF8F/l0i+Kwxwj
PmDujLeo/XZW5Ww5h6nxjfPEbDr8zgI9ssQB/i7Qt0X++VvIZwPw/V0sB/TNTjqN6idrNmui3SVm
+/IZEADLVUatH4PfYZj8EVYttPCfbyjr8/wGUAWCeOQYXb/kHiJsJlpZQLdMBLBavZbcatlHJqcw
cePEhkrNuGgodb4XBick4teGDUGerCjPatt6dSpOMzMx6IKFnI20014522/QfvpEBEoTJItriTgL
R7yBWXdBINkoCpzjJ33USwPXIJUCSk7930DYvxjFKam8aJkprlPcuMYdjQpDmx2bJI7ZcVOzYUeo
uFoj3noJEUn5d1hZgbldYJjDy1kgiaSbaDKrpvF1ogI7CF45bxGrGB5/nfDz1HJlC6nNatYOf0VV
kuzChHttFw09mA6YF4NnSGn6OBg2w4OvnJwnNmEpa16zDTdUX2TViPez3Cyz44Zu3YrYF7LTlRkY
MR1Ax8p9ylqTun7AZHkuiDV8ed3VM0IaVikNG6WIBDQQEkVK86oVSvXI6YatCF6SprUF6mkhOvHm
ItnTL8aYuGPeDLEEpCBkc+mKbnpDAISc5cQPhs3kHj+M9sZymFPCQMulv5ZIPHPl4OJKCgYiKZOe
Lc2EdX+Kp36bLlFCF5xKp0GrgEZ9B4EjB8g/FPYf7W7ujFKkuMTU6osrjGTxGo+4sKPOIju+ClOi
6wL60liAhzMTMeB4Z1KPxiqt/F5FLIh5ev2EQ2k5bsIzBdHuXeRD8PVTrqMjxjXzEUPt8m0n5UCQ
xh92p1rs8tXSyAnaB+UPWnLVeVRBo6by5niTeHoDtJAHR7zSIYXeDXWjlUUyHAX/E5NiZlKTwen4
3po7DCutOhVKFZPVv/NT/Q4RlWXFNsDGdsC0VsA6VRgDW3n80vcZimOuI80TOhq3Q1Xc+DsfVRLd
IQLzpwtL7pwb8T1UfMv8UBxNb8dbeGOC8orRuidAEj5JY+hN9Vxd8xjDBq8m7N1+plwt0KnTim/k
mGfsI6vDz9EGYdMxeOHmY8WA9pqavQohuPPBsezscyzusPx2i26Ah56XUf0vyBIcQ4EvNcHqCyZb
oFuyL+2jOBklp8M4tqzmlInZX1ge50+CQ2UX+RpiUM6Ug4l56Wuhtkn5BE8N9VFhQYG1G3m+Li7J
xHlnC+gMeV6szsODq5nIQxhI6G9QKS3B9WClr0TOxv/LPR4zQAzWT9OxUqWBtpqkpi9iPZZMyKI9
TRYcdbnjPAHeiFG5U+Xgsy5uaJL6FPgjIEMKYdDpXTsM0JKhF4hRfTFmk1yOHR4UjHkVmkpu/X2/
sBazpV+gR7WQmAZ1CQlfZX0AhAlDXSnzFK4TpP3a6PoWbjvNaKaSrAX7i2gP6KH0ZWgFq3GtavY0
36nsWl/j0m7O7cC2uk4uIsVSL6tdLoBe+sy9JhmNCI7ZpSoSHK7PIzx1rjy1hm/3Yg2XAX6SsGPo
FimEZLA7wlCRWnl/8/OowUixh2iwSJUIDIn4pQ603iQzEHchPJqVygciQ0AX6HYRdUqcFqj0xDp+
8qHEF4Ror732SidRrlJH5epBjfOiWJd+VqnFREhJhJBnXNm6HrpGCtCpH74johALfu3U3XfPMPnH
6rGSNV9cTRNk2IV7ESELlqWXHv8/Z0DtrHALfbD4ELD37C/be2Y31ogIJpi24rsTPhuV71XAWean
an6lARGH3IfAWOoiXYCTpufIUePmptUDWVHxqMetrsVkGPb3+GdKl17JC0sclmSWDn48dEaMrWN1
Tihrc4vKo2XnvsqjlYDjQw6d1oz93+ld1U5nUJ8wWxR2xl8EUmaOxZB86ELs/ZdWyu/YQUk0s7kK
dZ6SetGY6A5PfPyqsM2JenQ6pfN1N7XJj+08h2nXZ6mLT6d1qgMmnh87UCqBFulfan6NzbvFbK9k
ByGyZStDitm9TqPb9ag9Tm3NSQYoRL83mmSGZpiZ3idSagXsGLInlbG1Ymi/mSZfENDBBscwox9Q
jxqSVHaDmV5n+PXjTZv4eA9mkEuehBhmSh0OF4g/ivTqQ4bD8YdmwWOU6broW/zsCykT5xW3qL6x
3+LjE9f1CZYNcjsiKOo/DVFNX4H5uMgaVTuKWCoicdMc7Z1ARmyWZ16p9VEnjC5yaytS6SJq0PGF
so6xeNX+5wLQ7DmWh3ut1IvQ6ZidxcNkDjBaV6Jbn8JNz1XGCCiJVgc8eAvcpQTn+x2U8iDEufOF
loA4c3+cWBxaS7dA9KbwBwpdNF87k9aBbNiUcU5aFlfGoT0k34FX07S7DsCxwByGzSz5ZARihOFs
FNJotQpe2xWeraLa8WnielKnypS25Vlg+MyHY/+uGmR1/5jHdi603Zq+u4F6HAS5+hLmJ6jn7eV7
02/ebuT9lH4NXmAq5c9HiePoSooqJ2hcAFQQiA8q2UcFtfctXGlvMiuTj3jMi5jNcJHBpVwpoQdO
TWFqpMdJ8hAfqbb7PW636uilIg59HVdL9tpluSQ13HMZHJh+skfRT6sjbSXit54xV6quOWU3GA8+
73adt7R7VIg60DvWaVP+Acs3CLl1HcZDe8nxA3b9Juf0DkSYr+S82Bcu2QewemNIPVoElkpjri4/
YNc0368Zh76AsnEkYfUzRq4nkIVecOIiEfyCV3uCc+j4X9/RZHD1AWOZMxVdTgm+N6eUMBDur+OH
5omFUknqm8jHLxD/kMudQT8IRg8rMq30freox7hghW+wVtG/nNP+mPwf/Zf1tkK9IEGiMsFrkCpB
MTIlKNWOGgbqyuJoNfBSou1YcB/3VZi7MJRBMs6jvOgS3bF/vGEQ4YfVvuwTxZJNW/XcCtLuEHJl
y/haFJoQ8PoBMjSB4NKV2kLw1rJQnCSxY7OBQal4DSLMwI0v4NISPmuZ/EmBaF59a92H51lXe73i
NmF3kOq3ftzOuOKcr/S+3FwuTG582Bd+WM+yJIxerbvmb+WVYV22rVm4XJAG5mS3Isc514ULD8tS
4NUHCmjaIR76NhMZuQiJxZ0A0YWxPBnFpQ4i5zKUD+K4DDwUCihreIyHe6EX7XvMFKSdmhxv0ztZ
MdOLp/vGGvBWK4xLuDAsB2R1kLuvB238MLR2YtwiIC5JJoCwkOxczeH7hCNt53aaJK3qZqsr0bDC
a23oTCRCpO9QX/miBrDE0DF58FUATzFDglKKf4kKmoXZC3WQX1hC35VIYzKgWbZ5sufQK+ybCLkQ
F1WIhORMB8csG7xhSx4qq9jiJQt7WIXJtqMsKSwPojAvwGJjSgPhTuSS2Y4WBuQu+1bAvlPm+lV5
TPKZKTABJ8ZGioo9UEjokaEaRdlmUBcmT6bv8V/S5I8/YCQN8dAvq0yMxSUN5le+qdp9YEXR7ccR
+4qS5XoDjDnkf0kkTw8arHlSLx86o89ZXSJKeVxgqaO2BgGacgYOSKc+U7rzQkNU+FhPD04/Ptt/
UKkPG3dmBuHb+MJC8bBYehW9IQ92D7pPv3WcBgQ0vUlpGcoWnMCSlSKgVXFvIb73dzenztdT0MzH
hPKeZACpzco+FvE7yyaziNmto2zHh8jhA4I/6/635flgIndqofc6/KbPacMq50owY1/jJn1ly22y
NF8V+2lNWskrBoaT6ykPe6krFKGSbwMsohiz1XNweCT3r6BWdyokvrUYYGGDfiXJTg7p7WY+/BfO
QTZPDPKVa35TWDUuVGrBpeOAtCfDu46CsfDQOI4IsTp7aKFwjIwUqvxVOpKFBZY0Bc3/LDMy+Y8j
y3RcGcgPJlz/liZ9i67cvQ/+l2Vcmud2jvq6bSSo8ghYiK+u9A1g1NroKtvOgPWwGz1OWN+EywY7
m1yOYki401qmtbCYZG1zhO7d4R0VjOq7rjeo1GdNfnOl/GW2gPqzUF/FFqzKs8F35/euQ5SSQehz
bKdDvRZnFmTnZrXJFwjlWj8keP2gYaNa/ey4VZ/JYjQ22/XmP0xUO0y+xrkc1yqhC9P/XR2jL2cf
S6KZ+5YZ38ywqzwzZRP7uzvSCYdAgsTPpITnvnG/5rSfBq/lB5fpFCQKQr+H7dctDWI/9OpCz7Qa
5himPe40CoY68PX0gRdB7upsFpxq9SdYXGXcCFPJgLTsdM8XmcH+QX+1tBCfEhZNfJMvOoudlnLG
/NBJ4eIRD40lGKMfm319rf2rWNfHhY4KN0XYLOedtp+77kwYzX9477bq6m/E/8sIKqfdoCx932uk
KKDWKbAgKDKG2DikM6UnZqDsKfadzdIh140T5eeIaL4xOUrkTczfd2vpc0A+noYVT7wjUoUp4U3D
Wy95PxbztNWib8W/QXRcUY3KXIDl10qFXFarMKM2PkOmGNxMC2ydcaomPuDdyLjQTu6haZy5vOku
2Y8Q9CWsw6IZxLmb6ZDWNGXvQgbHEo7gl1rRz7WZjKMJauefcErOSubDaI54itxKVqWyhnTjtns5
vlmVKobQKi0gm2YPRSkGpmLWGSROyPgNz+8uQbb9tdi8QQ4ZUP3Kh+XCyn2PZ2tGr/NISzNkBTcy
IMhEO20oS/5aJ3rDK/3v/ezZcghbdRWcS4PzskRzy4GOTOBqPzz8rXUVkjnypDCeLKTNqrCeHaT5
fSUDO0Ovr/gPW25Yu7WVXzyfX1k4VojO3MjldUzXwFVKe0LAMBxChtnDAV8laaiCJNwz/7U+qtFY
ZjmRlo0pnpsPwfbTs5nllvWRJ03NMRmAhGeqqFAn6YJW0Ws3PtBkij2cx8e67TDr/SPP2E39MG0B
Vli2PfuJaiotjXqJhNUU0Pp/40fwLuL77D7SDKbM5J/W/yhyLP9uLXNq2xXlRv2SZMeojMgN/9VH
YCeTh8VoKg4MOI+LFBCW7lZPvPKkMFZ7QFipqTrGhFX0wMuJkcsPEZWO1e2SXvGlVPw05/3MrKzs
1b4hXGp5GEkwTYp9vtn+ApwJKGZNeVXvi/R3TRpB65yVl34l5BL41V9GPb21TCxd+0Uj75Z3xKS0
MBurAbWGx0IvdAD84gnGop2Ge0RGgaeTDgk2r2jtDMjGCf39fDmMBqkmxucweJWrAnTDYr/oLEv3
ZwTyqdr1ct9pZEKPrnW5lAtCeDpovKV+gmeW+rlrhwZNvxW1aw3f8c119GuXTSjTdMb4UXfrY0Pp
HbSQQnbnC5GV1hiHZt/kxbySEQTxqGL9vBBxXGBBp2TCFCbfMvkadfJLfhMokEwvka6hbxsIxO2i
qs4CD3V6kOqqoUQAKO35Y32WVi0xZR2RFNS7u5W0nK1I5dligqzlRLNs1C011wFl56uqY14YeEPK
m8TGgPCVEbw0s1ZSWzbIk7C8BncANaoLjMzdM6l7wb+ScD/8kDGVoLYkDAzGqtuJCcUINF1Hcks1
icOJYrm8FuuKZUW9kUbXFmLcXtRn+ia2F9ILVP5jA2YhA0KUdIXuyAvXrGr9gRxSHXwW+g2MYQ11
O49LJn6vt8B234Cq+eVITHyfalTzFahsBk3LBTNsDj9LjxjalwZyTAlzeaVGBlQZsOXso1x4Dt2M
YIjSMcgoAZfU5SwpcznD0bjoZCkMy5IkXkLqoXhU9+yDozb9AF8+3MIOXGRnhkF2DXGMTa71T6mk
vUu6PqCNbe2NrY2Ga/7YAqtaUpdgcrnsD6emqSNjOwEb0IegxQnP6DDtJvTReqFYqF51pJ6OHf8H
ERPF0yBoIBQvstFguWWGzUqv+prKF3fgs1yLF+82BOkTAUxwD9RpzrYvsRZUx4XaL6vk5VgxWBgK
80ZQ6NzSiNyHK7xJVHtFFsruPnXEEkXeA8+1HCV9XWJ2TEjds7Yug7Lkz++pZDwdE71kpnGqdye6
6bOXW26jGS4/LxtwlMQAvVPMcDS6HrBBknnj3sHXwvkBansrusCKb1lCzYGNszZUX294AuMqVmg+
osbXAi5QZLsDT/X/nANAgLHl5G93YTpa2TpL1aqWU5WF0sk7PkCIRbd8WFDkRfH+7WrgrvaNcaW0
vnrYti6oTyEsUi4BEKbcXBBJ+e8vg4BrX5qzSmvUWuuHpraXJNRNZOIMqRVz0c4lYC1c17Vp6Vbz
0bjZ+S1He8tQfE76HxkwKKmc5YJroD51zhX3if12QuaClguozZxpVDQP+Qn7FOkPGZ6m+YUPyRED
f0C4YH0crctJKmnif+GlejfHbIb+dqwulFyeQWdOZyRRZYaZQpAjD8GnaZFPg9GtiYFQiQitGJJR
A7JXjh6ZNa88R8bwkxEDTEXBLeqZz9FxAgnb1I9yZWf6pIicVUo27UvC/OIIxae+q6hJ2XSHJ202
mf3iV7RrnF/sLc0R5jixhBz7xiRlPxBvWfZjqW7DYBRG650scH7evQPgrwKEeawxxovKzYJrOglY
pE4v3dIuyIkUKaeQZldgcaU/oQFRcDlqLzzSUToFxilqz2eqIY1FG+BlBErFwcns5U119itMyo25
KUdxT0K6rm3om1/ZwEdIDoWoNwueFu0MurLFAAPS3KWagqctEID47UecAu5lTk7bjTEO3K+jYbY+
ZoGskivfahLRGLVKV5fah5DMf7psF1N3aT4f4j1Hpx6mM1IK32Rlr/8s2qUH/7l7lcBZ7wy4kkiP
l3l9Jl8LzTI3yZV/cAaCJ64TPMxcjA+/z/VQBGpraB34PZY+3TVu+5IeZsYe2YV0t0S4VkuPgT6c
CL84t58O3/GGtylvd17P+lX0nepZV0ebsik1FLorKVY1ytaaJ4u4wpUqRHKV2guegmZrv0IuFALI
c4QHbpqOfUq1wKbuimWhS5+TD98I4zfUrw9i9JCBwIc4lMD/h33VSs+eN/QZqWbpmNFKf7m3j/td
xzYhj6k6bFm44Ibj3+lTq6cGIYy4NoqSQsAmyfkihKC7smgQji3a65+4x9632jrOdT6GcN6zv+zf
loRrNwGGTwLtv9Zpo1yN6mFp+fjo4ScpkeNOyxuBPzGAhsJSCAHVwWCnj8Kheu/wpJzqeTK6RRHZ
fuebqrMJIDrKQ+roL9fkloxWDs2LoNy+8QUvER8OvaK8AvPSvPPXDoaGa/T0z9zgGzoLzeUxbPJA
zOa5mIEDHjdjP/VPrp7BWvnwFeDEznnjEqRkWL5HW8jmydOsRVKoTj6XAdAWJG1fChcVTBnnNJqw
ZaxfU37pSdVRSiDjZoc11TCk7bYNaiGMmPPtI6vb8Kg3OwG+GCO+2ymo9WWPRySyU02NYnRf1GTv
d6G12KmakwLuEbuIeXAldDxQ9H2SLLPkpKvLMEd1kGAl5r8pOZVkUvq1NspQ45c7oihE3/NeLnlU
vIsKoZpWq30uxz6BDXEcjyDzpItf6mnx0Oqjb6bDCF57ZNMMJDEhFroMl73qnyOjOUjuXNLHCxHz
LvABTpu3EeNKlXyklWmFx5sl79XTetQbkltXaecqcAi/4u54icnTuodGzmhSuCTaHo6gpZXzM6EU
wj470SJ3qX5i7piktPl1Yfl9iyfcq8XHSCE0lItncilpOggfQqYhFHNjIv91A34eT1fDQkLEbur5
K73Uhu8ChKcALbWrPdAsDCo86i+c0KngSWUg+aU/PtjxjFxxEOcsdISL1MozvQ/SF+oHL1Oz243J
Lp7enbNLIG7MoK3kNgZJx7BPAuNirfd7LYSRQeEnAt8ikvGjkgwmqnRq1qAClAqMRgbF0PC1mOQa
7LiIrpKBa/Z3/nXyA9VRfiCH+9+sSxriuwWt8eNH0W7z7D+IpQ+qy/Ah7w2ACZH224+hbq6c8U0J
lnRV4o/sO2jmblyXR92GRH03fp1HqHKyaWDm6siKQsRa+0kMb9kBObm/n5QcuIdt1MPZ0/NcSxeS
4gyFSIpzKJdectzF3PfvJnN36Y+xSSHGwj1fmQ1eM9kVDRiKFMo9ObCJUfn19916K2RLCmLkx5iE
cbxSGZIHzTE2QeJhO9NURrt9zNkG8URWDpBoIxMw9IBKXHo589zFvo2rDKNxJWT8lIQ/63zifzQ+
gAg47/NZAhfhMFO8jNr+kFaJ5/JXNj1knvBjBjlibWh3g+rRYX3MGTjcV+LGnIHJPVPc3pKyDley
jBtebv3YEbmMRn9BBBYp3hkTC6bdOCMc5brGanEBeqT++Z2eVSXrHLLitriK8EBA9Wdhm94Clpba
USbnGeRm7PldgwR7aY9lKGAEVhn5/gAGEuWME9qpdYfoH1TOKPOoZdIzqWWqXm5NwcRMHKNSFNW2
OL7mwYA989Kl7q6IFHKF4WeFVIoeEjOsOISokIEBHDRmg4jERvJR7sV3pFRO8/EBW5KzvCpqnrSe
lX4mr3yAV23WWdo6uL2sg1jOeYIyRyDgo4Hbj2rgoi9fvCiARlCyJ8iDuXcMB8+5LnksK/GbHXih
HKLzQVWzme7KeqxrAt5F6L4x8iWqAMz4vkZ3T+WYjqTGy1DzXSyTT1wCQ2a/+owOE8CAeCWUUfl7
j9WvFfDNW4UbsaBkmPrCqWhGOGRkQ10l/37mAK6xMpdbx34Vfhzs+yniE5gOfiLdYE6LlV584R2t
pbCPuehTsy775QSnJfWsr3sJWYHyDWrhF2xmxLi5x/PaBdlOuq+4YWf0TO4w4/EED8H/zczFHmrD
VpMqYhawkA0FfIhV5ZDaB04YF4JaAnMz+dGbbX7Imccpv/K9FWNS5T6WAjfLgzbBLb5cwFs+DJvz
1YLlMu4+XHqvdrrXrjVIJZBmEYMWP5lEm/UXWJXk6kpkIQGkNR9jvDOBuexBZcEN22L+CtXUyV0x
H3FS9ZGfRsqBhAlXWQBRg0vUS5juJv9R0ztMjSQMi+1ULSm4dPrPHBMBxVmMlL2sV77MKF9BWzKz
TH+fzvmfxeoePpgUyLXUU+LVA+/5UJ40Zpnnq/WgjaEQ8DLuNIlnASVIQDoR65CWuzJy90WKuq9T
36gSRIAjz9heEWhVkdeNg9le2+HNr8WkCeuVWWlWyBpUe1wAVYtjMCWFO/Jlk+32TkMOIq+l+O5l
9eUGFtXemDeIi8PEeeR4MvA1KWVxsTycG6nlWLsyX87/mhe/4Wwp6LRdbftaKaQ2KX9Yfo6AF8V5
OeX9tWMs/w+zDwyuoZsl2bCA+Kjbi4ilF0onfVmILxT6WCiyssGCOWmSSHss3JiaclyS1Ujgohea
SZW7vadlNp8dhNvkRgeOYtbE2ZthlBwIzbZSGEkz97CRXLF5UJKKADJwZQxtBua2eXTPaedmbAuw
/i2mtypAlsMSit5J3Ah7oolOL7cFp97BFk8oOYMNjkEF+TfmMv2Ubpz5t97vmP6LWHl8xKtB6ZYr
od0r8IMUI0UFuudq4RZcNoAK1PGV67u+tqXuOD7qA/Tb/NKus1I6n4ijOi9m2u75Es+62NxtCG7C
t2xBb/oRvYYru2If8mZxbXgMMbn301ibsPRWTqqrhUqbtxn0xclQbcQkQHNKjwDTM60ZjZbC9Nfj
nbdDzhRwStYQS9cqmWEQWmY5pQ8OD4PJIChs/zLLpe6UTmghwwMYVGA+/vYhdg9k/FJj/js28Bga
LeOYVZaCNg5q/t3rQt+5AlYZz6BZB0Y+BVMJLv4Cyr7GabMNog9LJgNXSvSCAij6zOvOKWIF0OSn
9nZYiF7lYg3CRIaPsB6pGCIX7CK5qg5ift9YemU2qUeFla7g6knO5YAtCK3Ciev6Uvf0NVtwqdbr
p5u4p8+sd9JGwKNmGgOmjY6atggqb5nD4vd9jBPEbaTpGksLvkWn2IjJLswtsejdc4gw8W6mERtj
SptZcEV0sRCf8SvBdJNEW0L53+aT0JkMp3ZM28C32FoN2XGBwzuUBKdn8G2w7gMOALqbJbnoYha2
ESlyXq2w/ftfwXIqoW6K9GBe6UYI3EQGnE0TyffAG+Ly9iJxT+2iRa0e0AthNMFdeAM4xFWSle/j
SKKCA2izRZj12/c2UexkGcDNm/6a/nPZX5jtMW5OO+IoTAlc56p693kU1UoVbm9GMJQbGUPc1bO8
jPRr/dMOhsJyS2xGjXwBRHCwMTTPDZVrNV9p46kYSIOPQsjaKPLQ/TcyUHGKgA0NYcTw5GbXyLI2
XCbloDlnOoMtBD2uPzSRJnYOynM8jENbA2UvTGVgC3kVTa09O/sndtcJzXYbWFVkrDFNSSjLuO9y
eDTfUdiAvqMatQwI89DWRg1Md3BYb75Q2xMvZQmf2ItXiis/gsJ1Or3CE7UY9A0VPoE+bSk/tqLj
oXEbYz7dfsFy8cIjuEpghNe4BTDUbCkLoDmF92CfVgPA1yC762paSUyBkAoAFbnaVeKIWv9BZHb2
sxZVwv98FeUuKNman4EB9RQ8Ov6xd9ACxtdPMs1Qvr8ElD5D1xW50ocTYcS4rkMF6FfCZ8tus4Xz
UxKYpib7j6nR8wYzfdLL81I82h6RBP3ZFpb0jigPAXMAiHRY34qtfSaJRfU6105lum73SAJx0jlE
MYnI9T/EOO74h8sUSmNaed1tD3pgmHOhlgHWrE5f+fvw+10D9IUq2dIJkztwOWBiRFtdcy/LyQxD
bWajP4/Piht5MmZjnDKh6KVzhnALPX3QgBh8HJrf3EUxPOrxn8VWSE4QBfV/gOXGgueJcldzNnQD
YK7Ht21McSXoIWt52r0bokRUk9Nlv48sYMBr0db1K7GOFyIJ+i+aVQBytX2TT4shQIMoAoxXr0/4
g3lNBvk4eEPMkZnkqVOdEaPjjRYXD7mHjpAQXbSrdfh1US4sE01/E3lpoIWya0mrYvpcd8cwTVTR
nNY/NysnrmqrATbjC54U1mFj0i8dXvSkajOxEGVf6C6I31aNtPFqf+wQHq+CYku7p75Pdmg6gx50
5mBgawno0BqzJhbN6Z3rUqHQF7tIRoqKgaBvaZ22J29rGAbqmvQx0VPnO6AXg6w7cgXs43BSLxYu
hOCDrpVy/dvJ0TS9To/LzX4fV4X8w8UCxymt6eEs38vMC01lBEfECdiVX8SX/sdoEoEMTcKKFzgr
JRx0Wq0WQb0EviPc/5Hag07UYjbb9bYp6VFzRofAK1/58mtl83IzpcIfHRYfVebGbQiwMmYmXJxy
CJRX8owI8DyATvj0dRXdoWSXiSbOqUHlJk9fTXXAB4zIYRE2LEHs1xpEf/iukxpfgkmSlH+6ZCjY
o+BXXgmKV6HLhF9q83U4jdOOyBoX9UJZH+Q4S4jh87xY9IcE8iEIm2jvM2eBa2019ABnaMp4cxbw
J0slvFbcwVfcvb5kdskkREqScQoHclY2ZcyjTiEIn0McZf26W2y0SO2PZ7ja7AVmEXDaIQ0jS8wU
JWL0wgrO7U6qz8jdbeexCUp88mzgPkPTjzvOtu3pIhqFZnbrKAM+4oNv+Ckn1FoUxYPZ+6KXjMpy
EVi0intVPKKtL7IybpL07O4k1wADhh+FdYlwV/0r4cAEcTpRYIxeKFPSC8QRL/3cTgoCRNywCHoA
a5bTJqYRBadvt6fnYBtllT9FkDtbDlScuu9robzw7MIS41q3oN/i504wDzfCyOYnYiVRkI08/CBU
2AGrLW+oEyyVXZcPuJJ3iiMI7pIRqj31UBDtJfWwYBDlptN2QVj7wdZmGEhvklyCTcF7+/umZI3h
32lKSFd8cUdVN6jrxi7B5RorLPnVRI34/WxBzJyisNV/Mr32X9uEZ2fxSLmW8Umr7QABnQ2fXoOY
USQXtxVGyHKPvSiSMOTuX1OgiG5UHPjvRxneq6NJIUvbUqgr7qiu6dHLp5yJO/Nl3CjvZdRN+tmE
gK/psh1ERcH+wXQtfkaCb/U1q8uA8lJpVtX2wAzASFNW1R7PEL8VTbc509og3USE36GeaJKkKogn
dCFjTvJj/7bkB6CSdvhXDakmxKLlILcZzD6ZvZw3dnlleaWPRQ7Vw7kEnuZF69BjZWCUbpkWfuqy
sPIVlQKyVgRT/Un5NQjHFZU+9p8dmOwq448DWG0QyZf2tkAGmGXdevMQVDHarseYNykI6TzmOQk7
DwEzB0oENnjxp2eJwICpopLWUECIr7dmQFmd2KhPhcPlVO4hIfH00qvfP8nfk1poc8Aw31osZbvU
WmV5/Z1aRSASLJznxorCa/n3APq5sNoAPb31+3t1S6/6Rm0BJDjnQPl3jM2CuFnHhDw1HWXpkK0G
rGEb9MqOEz3auEnCDPmnz2tD88ZweTOdBbclhCbSeupEaA5ng0IjM+D/R37hTVjLc7ZA7iHlns54
bxrAHQc/bKnKQ5EtvoE9CbW8fAAw2pegklsEqRpl0al3AUxvrnWZx01JFPdBtl2XNjyZsN6SXIYW
Lbg1NbRqiiTFo+SIMPrb9zQ75xGSluYccYgHnxPkMGmJZMJh+rZxbKjW53mvctZZBqYAN03PWqeJ
sxX4fHzPPvD9CxOHE37zkVKB4Hg8VSeY9OzckACp33M92hrKh6nOa3TXQouAs3pTa46C/EvFbIwC
A/n0GR3Y2Dlkwz4yeAY9f9/1N4zw3pwF/6eVxH0PQ0KtGv8+nzLCPLXtJWlLDDk5lx6470ifE9mp
+oQNXDRjNvqD7jl28dSJpUxZKbzmqbW4+1GDxA10cISuFDAAWinFuzceaVDmGqvQAUfAFS++hhUN
dmo1mAAg+PQ6NbF5eZIJKJqv/vFoa+AjpLkdObRo8ZUyof0i8zklyKKyOsZr5CK82T4AAm5w+elO
w0t5csKLR2+SI4p6dyEeWRHai5oRhbh/J0Nd4Zlmkret7lVxvDI7HXEik6wSMk0jRa4cJ0hS8D6c
wml411iEfNm/S5wroM/ljMLxL6c6FyCu+K1fHH8ug4dJtpqvg+lAr3lH/ytt8gvfS3aJuwzEnX1T
eVpUKb57TdtEw44pgTQGlvwJ7JLhjiir2JazWIcFESQ2DzRe2plK0SdWLqlGXXAGnQzUOWOnEOA6
lkFEe2LFZM0QNauelSCQgsI2v+uA3SxXOMGOSHp0wRzxb5RD8g8ndxEdFo0KEFWsnysuz+Eo/VuL
cDEXby8KR8LbufZoKSzHCQ0DokZ7Wnf+Mmfn+vqXXbzIuoLLAYrGWheO++XLzoN3H+vV0OvTMfvj
IvlIz4lMUY/gIWWq80lEWkR2PXKcUcQAXxsM3DiT3+HueGybAViIZiz70XQ1eIm4m8PuCLOJnP3S
nsuLjTMzjNKXKlaJxkJgByHIGQVHjvNcyNB6HD9GkwPKwMWRR9r5WH2sp5ICXSYqyOYzlRcoVkQI
ptvueEeQ7aAscKAO0nNTuig8wHzrMfc7zATgsyLjF5cqX3isn5ADC8yuQyq3zCt/FBYWDsSjK/I+
KQF4OWK4B9JGB9/CBTz+iHoUsKQUheAiTWlpdLDjM4UTFNHetmD5JC3gw4AaRjreeGStPC2U66ql
YyVQwSqfMGhI08OO5esvcs4qIENYWvgzj/z21CwM/MXMmtEh/0KK7Zrx3Bo3gRTASXNXYsZPZOvh
l4E6c0aClgaQ5YvNU0Ak5Gqu6A7zCvIdf55Y3m0gXIRtqWizfXeI91bK83mafkHJBttuX7ZHf8OQ
E0CE6oZLFQrBGpyup83aAl9oJyeUvhYRZmSwn6ncI/8TaLo5tVLYxV34/GorxYsdyqqore/j9slT
ZdrkhjSYHALfl/8TiQkAQ1AqbHh6423tIc664DamcBA46BFsNdtecG6f+L2lqhP2/x6/B2Pj21Y/
75oGbFNNggzTwOpE0SWcw4mefR4+OZF87YbL/GgHjkmsclf25FTefo9UW5eXonwmNUmPhxXXZkL9
EN4633yRy9WA6lqOIxoYUc0k0cInxR+a0/IbH/05Fvy6Ay1bj/spSAnmzd33NojqkkSD7Jo/B9za
vz7beX9+5+n/Ke+2oUaf9C1TcheO/QXKkkABuU+44isPL2o1phxCAS0aUM00xvZjW54vPw09VJv/
8e/18B2STyCBZ7POyN2VCjonhJJODlUdwltJvxvrA0OFMAUg040kBVZ96zT4VI5OzuigPxNhep12
Lj3XNp1pNP1RRLLhGKznnEFUTi/21T+UpQIrLSyCdQbhqB8bl0mhdP5mCoKNpy3ebwUV9Iwt3sPK
/qwRmcAEWxKUgnuFT9n5ZSMBvSY1wbPFXlL0xbG79SIA6dATh+mJwUHY+bPhFfd0ptN5Edj1hrj3
Zs2d6spzfYGlWoHsOfPDwjTno6w1APwXRq7FzgtEGSYibzo0D6F9WHDHRWTYEYEHlG12QMgdTrbI
qDiuY+NIPYe/UN8b4WQP6VnrTN+pLY3Crc6KepJN3sIN2pWp3/3zgE+7aXj7KmFtb8Af27B7joyv
CUFm1xwfW2Ki9MzgqtpKeIyEDUd74ZZXWWQPUpIxsRISbidG0jgExVisWgSXJvK6TLd5e/tIj81F
meA79pje02f8nO6t5Ed/JAJDSOxTBl2wW+r0bTxABqBtsYSx+mjce+Sc8Ph04CBTYnV55KJgjFYo
y7/GhySa76ZEdAdK6yuX0Yjfo47A9Miiu0R2fWOKUzJSuCtuOtf2kBPXRJAevInjYqJQEGT3KCx+
w166bqvXFrixG5GlUae66IPknXvJYZh3fdZhWYuBqagF0yomaE9zuMall5MdERmlqIdBS3vxBa66
M0FUcT3VwQEZzrtA1SoBfqce51KiiGszYcSc5/wD/iJOnb0FtpuI0gcTPz2yhQHaczVuy67u+KyZ
Knne4Luqif03q3WUNN4SL0EWhFqNjizlle1+9pBp83qPJucM+iVstU/V0CnllfEqZsvr4Y0m90nl
xORZaeyyp5HIt9BbHzqlO45syW/fO7DsvpXbcfLHwGbfkg4nDVNSJebmuME6YnTZTSWuzyini3Gh
jv6Mg1Cr+4jMw2W/NwUe6rqKfHFi9UI/u9rE8EwOvOQJBIpEslcApDPMWaFQx2Ptx40EIif1FbZV
UIg/n80xeFceHTgroHpXeNMxeNTaFw0iq9JBIDdMunRJ8FQJcm5MFEC8wDzigFJOKff9+/K/iofQ
8AIJwwHPZerPaBkK+IISAVwwcW/Un1NSDQ1KOEIObNbrWXSCGlLXRcki4Erb+WRKYW/WTgQiJ6r3
Kjh1eGqWpaG/EXX1vIOSmTej3Bny9Tz/pxIjYyk0qGxEbahBIFvzaPcrMPeKt9XJGH4bnxeT9+z+
3vG6kX5MsNADWX/HLzUCKZyyFkvzLaEZUvm+y4n1+mPoZrI2p5s4lGqXFS2ynP/w8sOJuAt3+dK7
sB0wCG0Xj85LqGD9yJ2LxnKtlGSqmvX7L6Lg98dZ4IngZePiUII6mBkLGyBVh1FjnITlSzLRNmUl
jkenm3afNG5FywTWvc7VCRSzMJtPVrh2lNJIZaU3QRm+jaMo9Qhu5g8Wc6hFk4UL3b9H7w4MRpMR
mIN/El75LyRNZdoG1vmQK1FgCz3KNfHKe3hB+DRYzTX5w2IFruWnLZ4+XDwErnGff/YD5zN2f8EM
BLmRyEDsj5asGmOCZ1XQ9moqmabh/ITI3OuBdDFKx82JBr43+2YFZKxchBBmJyw/9/FFJ9OwkFsu
zUvovNPF6kZOhESjpjTEuTYVzTjQkfUubtpaGES6cKewCLyscoJShTnCESu2xUZVX1RGIqWDwYk+
sA6/9EvZHKbM8Z32Lcgn5I4LoU7z3WUF427n85xExj+rWWf2ETqh79dOGEfytQFLlYLyXclt2ZFP
YicT0+KnKjhfFNJ+S/16MSG4BLSBR6HbI03A/57t5i4EwEYIc8aLqjKRRC78X2OC/TL/F+00flyP
Fxd4nZG5YSAa5zLmDOGuLNv+VmSASpjDCCjin6DVnEqiqLL1gm6dz2XrgdDxvsAEJ+/e5EUiPeJj
U7LbtmOZ9NNIjSxEX0fV3lVg4EKwjcJRMu7k8NhCFzCiwPWFpA2shDmB7LoP/JJrCfUMqj4PDvmc
CI3HFsamFy/zg1x6NUbw2dMsBv7YxNI9slXMLwMjU6l0WBEAvklT7Dl/CnKI1s/OXfNn0/GRP08y
KGKP/hqVgCMRRicW+SRPmueR6lKLZsknc+1vFOeixdFY5raHkW2JHrD0BMNIf61yZlBafP0SHaOw
F1jz5aLV6scB5h+nVkIhp/zIU0l+6RMVbA5NuZX7MiYzxtL/TfmEHNK33mmR/MTrf/hSiRVJLwzq
qHEj20gdU0hvlUZCVXcn34bUc0+cMX2ElWgtJlf3JPljGO2ZJU4QNE7X9o8RfVLi4q7dnPbMUNmw
ZkhfaoixutmPFu7xETzOQmSixapPNWOmdgcPCqliNJmFdOaCrb2iQHuGQQGQaIQjdRV7f1AF/M8R
oBh5Dij0plBzUotc2dy2HnuTJzcs47/aligrQsECJjD1hUnCBxvIjdzYgW/PaQCNXTGJ5CjZMSr6
VpH7UhZxhLdvwO8Xq9wqAVAmLjyBhbsjfAbpP+3xsyfAcNz2153Y9AZ2CVG1bwX3+4fmoHerluCa
UhpXvtIGgZZfXn+kdDX9wpY1ubxHY2DoIYvRVzY/Y1ufOQGQ87D0LKs8ZIIjk+7OxO/P4ok21eC5
yHCg9LuAwkJNIgmLTEiIdrCbZ+GBux0EGtLT7XS+oqyOP+cIyiv16tR/09Nf0KxrHnnJGOAWN07a
o8PWni+dDk7s+wmgBY40qTxVjMUF4zHv9fpKNWRLLmoMwrv0kwiOzT8I77xmua28tB0qJutoHh8C
xu80CgKFk6A4hM3gHzfGER0r/wtWRxkHEGpxzs6AMQKMhKMcBYDKhFFJHC72gC1lF4jvlRQU2Zmo
glwoQgIKqB0Vi8jwGqU2DjIUkZgLZ9cxoCn7ytAh/wuqe3mIwPk0JGz86J6LSmIVktOUYuOaCoJS
iW4ET1/NNiLlPzFOGm5PI9TK1x69PwqElO8IC1DVOiphM7QfhZ9D9JtGv1O0comz67QwHb4PiUgx
MF50YpRDfIywxtQuNoWWsKTFtIkPRyZNSL9nCz+8ucVy9a4fQ35HriuONWFXpKcKHqWOFfe62wfl
vrCw99Z7qJNov5TkvhsQlLZOZdtixLRclmcTrFJbic3guTjp8Osh475uTx7K6kUGkFVz6iGy1ZTP
xGWJYXLLlvfAcjOC3EgfcjgXnC1IK2695QhpggA30GH2nlOTd+614Gu4SprVkjRAk7fb4jgoAhAw
S8/gJO7m0whfl2WauVZT5prb0neahj/NP2g7CA9ufB+IPhUucLRaYeMVYsGXBvQvWCvyMGjLxgpB
mTd7HC+aco6g+5UcC8F5W/L72TRnnynV38CE1tH+TB67a6vR3B+M0MkD116e99N/Etp6Tq9SM5NH
uWBpw19emg0evtIgEJALIAK2DNXwTks6F+5T505sda84yLC7m7y+M8NJRH9XzX82lbEyTiUcCY5M
ODsy56XXFTKHRw5x1VCD1XsTcBqvk9Y8BBkPp75ky7fwyYxFTUroPMte/A6Sm74OcL1i/0AONHHs
XGhImu3e785sNZJY5dGaWPNqAefpDsoCDUvPBVHb+gM+PLZ3Yti4IjV0jI/zEQYeMXMo76XvZwmJ
RNNJnUDyUHgDKTFTlWCnYv5SxXDhivBhpRN5EK25dvJVvoGolmzfWZ1uGFFLxP+4lIEE1GBbK7r6
heiDUN5NBFZk+/PBO8F9UYzq9NZEhRnO8CWnIpxsB+4PNS94Iev7UZZPfji0zb5z8zwuFWSNFeW9
T5MvsB1fxutrYG07Y/BIuKaK0cOJPqex9RPr7fN9sQzVP5wkvAd40sElM86CZkldzvD+36xJWrJV
6f3wSm++9dVOGqSTMSrdWhkfXC/qdj9g4rz0QWYQ4zysGg0kuK9fBlI4VfNPsf3VZs4GngkMQu/C
Tx+eI660vH9KDz2XEriBSZtevODNoY2hVky4bNolu6B9YU+0vp80BRMBl2nzHavz7YyZrTmQAO/y
Yh5LWg6Cgnx3WPHUDe6wmPXena2/q8phUDNlWnTMhscKhiDf5MWxaHhwoDRPtnm267yOUrgB8ojZ
26T7SzdEQWavDDcv8buWit6pQUduyHVzhY/zXc5Ls8WoIMEMt94vTRYogD9dqrrlhUA6g5ZP2kO7
NAHRrNrQ5MQu+8sH8cBPuWnBtnW3XUNFXKu8x8chn+1wM+ytdLDWrjT4M6QoxNChy90PwdA6ktug
bX3MJu959Bi0zE1BfcH9hhrsVNukz1dxl21ex3FIew7dzRZ+XppuQP3bGNqsh8WdrULt7XjxdMjo
f19f+HIR/6ys8koX6RQeyc5157iT3455KHdg9CvGv4E6LI1NydjrIYncyKluHwoRAFpJrEveqZfq
MRRdNOIoN88Cq9ngWfpFcWeUHM7602G8LTml5h3k1cKEdjc2Kgdzy+Wl3xmivxkcUQAEEfT8K1SZ
fCkfbBNrHRVolDL496YF/0pCpSiFZ1+txgKPTwfCy/mHqYdSqZTWR2SrQWxpck9eKcxF/Lt12vUm
XCAKiqGRezKWUbiADtrbFsn4zIAHgm5Rjf55tVPtvH84wUTfR7hOhrnwz5DHfsbpnaAyke9IfqEz
p8esSo+1rGd0RD1SmxUa5mqcI4f/cn0BQpxHQcUOyipcN/JDyOhXsfO7WHAxR5prH72QeykTRkA5
VfgmeDGuzT/dUwWzogfdPFOmPSP5JfTa0+gPSAq/UUrAtAEogRky0rKx/WowVqW+flc5aqHaNORz
Ha3C3IpRh4M20v+rqNKYgASdH7MQJwd4t/lopin0QGQu9qeC380Am/8gSOm1K1jnknTeeOdriVKt
F5qkzFLIfyMUxEsC/+DHkXUGZiE+kA2c3QBRE3vr5l28XmBI7J2rBP/2uaZ9hOs00z7uREKcBOas
C1nfUAeRRUjW/oBA5613PyumC/y3dfr1UzjSR+UVeCLbPKRFuk548WcWKpbgoJ42ZM/pEeeZJYqp
xA3P7dK2GRdq+rk4bagBdKAqIw4U6Hz6CxmZNXyamSS7lyM7L8vTpf6UMCO2XLVgLfobPPiRSwCO
e2gV7ZzeCwnR7c7qxMYsjD3uLVhFsGkDbEkdkScN74ru8RQRMrJ6v7orTdcKyN7HfdgeT4CbOzPX
ctie5EXUKGqfphs19EGmoow5VN/jXNxa/tZmyscM6fE5zRmtIr1KZKwjJqhFchwy8oIx2/odn1gj
jlhkHeUCaljsDtey4RYWJM0B/+GaFeKak+Een24ABAsNvH79oGBNvN4T7bWmtkgM/KPkLxtQ7cr2
ILe5/juzR5EVqZQ2S3Wu4VQ9mCztBSoGsUrZeEd8d+mTSUaO6POuA9oZ+ZmA9oZLBL9iW4xy3Uau
0sECoFvTYZ3q8SY8fx6ZcFT0Dk51/x+sXOhLF1+rmNnGzhN/5MjQUahywlX63hZbrdPn8h2KpPeJ
yhkHYMigbcDTexi6FZZ6tq3wS0ie/6Ev3YJS+AGXM7hCKNBbpnnl4Va9djqHsnLKlOpG48I3VU+0
0XqkZQJj3j6nbyEGmA9tIGiGFB0xlQGsQtYJqv9Dkf1x8tdfneKi9GyLxPFSXqgPPhdP+dcWcAil
9qYebpbvGftF3Eegetr79B022DzuKat2Uihv3DdhFVOzBquAY8mS4SciT4ooYcwZPl7TY7FX+Af1
aX4UUMGu6uP5CIsurSs6R12g85aYagd0H4xgJPkXi1t/9I8O8I04MsbtthRFvAArzWT4FmnkBc9l
8I/1NALTqw2DxqTZgbK4bb/lpxLDGbwvla61tH/ZKgDnrt0GjObGZKT2xagkEf2z1bQXI/mO2pie
gJLXuPGYyUZoQyOKFQgNbVk5Lqny6pWv8s5zZjVa6KiFrEvDXFWSndGUIflnYTOsJIoqjUZs9WfZ
hYblgZrV2Zayo6EKpO8Z11NszuyFF4t5UFk4OCAkOwjJr09OwjOKp6Xu3Mb1IOb+5CXVtitkY5tB
FgxUZKCrkozcKdC3jvmMvS4hWEWKBEcarwbsm4WOm9ucj5r31TbAMRfYrsL+LUlCMFNdorkrYqur
ZWy0DvcsAXlCqulaoU6RR81FBg+wVou+5+hK+XC9MYbXASp5/aVaF+pXpHEcROtqXcdMYqqI7ROp
yPQrEDnGrEHDmp1vlHMo3++nJ5gDnMSBd+ZfNmdW1zSEf04dAgI4PDLBZ7r5pa3LGsp4ntNBKOUo
LeUIrRwC2CeBwtZgfHOd3PyCmQyzgz2ZjW1+jabDiNkoPaSF6TATNn91TvKvRlHa2yiDppqBzR+G
0D3NTMnIoklOcztqlMyDjxZMc5O1pSOwzd/OK3h4UiHdOSBtayJvu2o4imEcBSGa3j9xLxkw6nUh
1T0ev/IQD2bq1lNYYfKKHlMxed/TEYXdcFpGtgiG5Hdm13VAfhgJ+6mQHQJVLJj52ktGpuws/yzu
a23ylk7YR1M/tDJATPNCWMTeNscwW30iWsMzl1hMh1O7i2VGuJ3BfdBLEJBvKFPMi8Or6flqXNkY
NhG4AKkLSvEhmj+DWw/Fy0lb842wTr64R3VRdz1jNpdLsjheQpn+IwOCXPLk3kntJSNtrmEpVcMl
OMz/RldSzau/hKWGnWIPEmkCkofMrEeSmkAqv6DblvC/b+pQbp1EiHc63znro79TQyye2mfPnBhr
AhRCncTQVEoC2zxVMFl3S1/5MWkqSEBxzXYy1udQN2bt3Jc/nhn/RziK25gPViSmZ4pwjNWIHONY
JlUNFelz6jeEYbJBz0oMMagAd0CmiY9StfyAV7IQM3gHq9B3C7yNKEwuDnzwrjCNJTmmmbPPnmpY
VBRG09D4L6HU04pLsA+XDM91+TfwaUe8UWPfwXCkt19e46p0ophVPap7FvK+9LMCsrIgpAWO39BD
2zFPtlcsiJNsn3pTk/3UwV/KRgsBY3MTuavxXf4cQ748WavGcXEGSCqzwaU+yBJg3ailPlIxZZoC
PD+N1DSEeFNgYf048P0a283FXBPan84SzqD4K9P66uwYMtxHVRxYZSG0C1yCekRQCWR9aFCEimdt
2HA4Y5vn2c3PalehQSvvEwzyk8717tia8tIP/ueTWsX3E8zmddJftOryOIOyZntskMa1cHU4Qd0b
d+jJ54x3GMg8N5goAZWFEV3i0KLN++ldjxnJR3XYzJhyhhZckGJnmzC8L6mjRxBVsR2WE50YVJxy
gVGxMRyat+S4m8Scm3U6xnaa16INOxXZVDtdJdG50NiMU7om2P5HpzYEbdpMvfqbs1YlVis4BzsT
nFAFCaNP1QmPwq36Goq3SDihy1+2MPPxyBgv2+Xs7HEqcRcPM6l1AiB2Q4T1vzqEeD5ss6leDW7t
fErOhtP2KeCUU/HMKp4tLKwxieBmHUlQWnCr6zkqKpMGJe7+U4JgLUvH5YmjCMpTtiRzrVCIBNnR
/PkC1+uTaun12LgUX3ArP60cYsfyYsuvO3M7imwG+dbYXwB8RD7MsaWtnCQL+BGZHoWAvFGznIcH
7yghWRkHwEpvEm3E4XmuKQhIcn92lbPSBSPoNBgZtkDRFm4Jrd/KQRoP9fa9Ks5FKvzV6Q98T8wC
L0NuX4LHSXjsRFqe0b42wCmrQBfa7ITC1RO6cI6afbAVP7p2h0yjyKmqb2qbQF7QQMmzjcaYXVrF
zBSgCss4cXQXQkXTbAaU6hBSEsZ0cJH4A5MhX/VKNQjao5iSSaCeV08r9XloflQCLRAnXkn/GQ1y
EL1al2gqIA+agPb1KYZNk0PNZSAx9E9F+uuCe5efhatGsU7oaE5B0FYfrwGs3YCaZXtcy8zimJbb
Dz9GR0JJimMwLEMF4Vc9l82aKwPBJ0rG/CLGEO7zDRGtqDf/Cjk0qjs3p3N26+rH6Ih9BT1zHHTU
ypbWQqLRUFxIzr2DtcO0BkyRDQYwxMuOLV4sNsw2BHMzxKD1tq8USTVf69VHmbC2SYFZAHRtbDrc
UN7wdUU7UDYV+4YnfWN5TJmI/Dgxq/ceK4K10UAe0gNLOmyFhe6kxSNbCuXGbyjcvDJpS4AmB341
3NGHCVo8vu119Glfu3vWev0GTeuEf7LwGXnm3GmdMxNTKSOCQHaqMQlGajebI5wYVU56CZJftNWg
97Gu6fSGKR4/IQobw2LKwf0ja929J0txzPkQo831XF1hv4IAFFXzVXgL4cqBaRv+UtGWbtkFQTxO
dWHEqRqAJoGzMdB2OoC3fsgWwafTRIRYCC/m3K2IumeSozPLVylWRs1JSBRU2l7HFTvCQ12KRa52
LMg+w7Kpl3IVRWzn2yVJGZpJq+O5AE7gdqTxf/0r220y8++rWWr1HLDkdGt2sq2REA/AVf7cs2qT
p2XVbcr4hP2SeadNALJR6E/CkXYcXFsP3OwiRhPi9mw3ZqcrDwvYA9g6u0nfjwMAkW7QCpAa7Gzl
WPpBb1ScdT24bRemMbN7N4yqeGaW09LjlKIWXkcqpKL8+qem20tVAUMXYJ0/cV4cUuB1267mq9Kl
dfrK8TW/JNKlzpOS435mK9trEMzTnv/H87klW88ws6Wl/jOzFY4kbnztd/ysog02ZeJRzrQ9adOL
cAb5cJZoMsbFuYsYSIrQA8pM54s6fwzvyqANLzNZ4clWllwrkYTlgS5w1V3CpLUqnnxsyeYBqnAf
ju+PFgoZp3XNEHpz07QniIMcvd1C1TGPWt2HUmCrsmmlcbtWrYCVKcwVIdCeHuazRz/zCQvtAJXQ
4F/Hicfq7oYujFxGlgV3wtFE6eV/o0pwjuNifdYV+gY4kb9TRVPxzSgGNdWdM2Jy3AvjCqAVbnkn
NtqQ6VYDHVOYccoQaQkpUidsGjrlnYo9mIi3mexMg/G2KPaAu3nnaSsFEWmN7+g1ov0qbHhAERpg
gNQBvFy5QeDZDKcnkvoFcfN+d6zuzSF41M8NFWrIbyi0dJIXzuvicn6ypwtyvpN2dh8xxzdAR7kN
9xFCjGWeQIGi3PWCzhpV6m76TWnGT1vOPba0J5ACVay9/up+xZ9/2Oy9HxsJ8RJXem5Fwlc40IQU
IJXzOawWqdho1kVIP8HeybZzqBYqqYHJ7QTw3KBGU7e/5RmsTv2hdvrcinZ0aiUrazkqO2VikDoR
qe/UiujzOg2SyZnESgEwdhDH8Ivrwjp4J1Y567FHzCf42Wla5UL2fa6NG9awv1AkwBAmuGvLwaa9
YZAEpTLU0Z8z5l8brPWd+t9gfokVlVhQcl8TISnbh59cf55hMUzDRxMtvPjJ8cAyhtmM8Rsfx/+o
iLzUtzpNlqURJ5KavqeiVV86Xiy0BJ2qR7XAILwngkxV++Oie/fuBC6B9e/WTuLm1GeULyeWDizO
IlE6y2jM7Y+1sWTrwSQLzTeT8GS4B2bPtqINI+vM6xE11p/mLX+dcoYepClL+gmmdEvmNN01Biq/
vfdsxdX7oKpCeDXQTrNr1k6zEJjYTqSXUpSDFMttkOWzEveAUuM6hpOaCA7lF3I53Fae5yc7zEEQ
PGbpjKloQbSz34KF9Wh1gZjUd7Wo7KRbTfERMxDgHCSu1GQOQgbqzX638grjRuwDcxUgtoNk0PAC
QsVz1AlH9YbmjI/2daWpPP1DDoyFTFEAd/lfiA9/aCJspiM/7tJ0waicnb7k6ednIyITd3GUg0ED
DhlpUeJSQ9OAgb3sBKFzRcFgaM4crCLzCSHkbtMkumzqND2+v7udD3PXZpMV0T24OyCTv026/OqD
+YAaeGgvYjZ8WGGHcq+fUkY2/4qsaXTIKVoIauTb/bXwuQTA6z4Fb7oLLXLvs6iVhMSmlGHzGEmF
8xRPngiZwyr4EkHYM5bA70JEq0XJmYFz9cbSI/JAhTsf3581uSaCbEwZ2h4D7JVwam56AXJ7f05Y
Bc68/pJ9OaoyjfYp4EGzJwKSiK3XznRhsDF1o+Tw5A4sJpcgVmuzusOkOCp7qca+f0vNpz9ZrFyD
KnIBSXUMfNvl5n5ZGLWTfmc2WNTVl+i0HhCRWpKPqpfbpto+wyNWekAgi8GMiz6wDGwkbXZGx4eO
/W/3T1AUOaiaCjWQpfuhk5//RbA5MqbGB5gm6zacQIPX62WOHN+SWaYIQSuJdCSmL8kzoTbJepba
otU8vlqbd3q9XWwR3LS+LuhgqjDWnSHdPo8N+Q9i1vXi29VJ86srM7LOezATr7X31XSFNXv4ZVZC
wJu6skEhSREXDno0lukhHUA1RO6L55TU6UHsYkHQjU7BVuY27KmupqpLb+9iomGOBCUblGkUIUM3
1K2338hAOq0u7bFX7nGVkkohHSCPsOXbvGpb8hDLkD+iI8gKKqkcFqYTt8KkBWjo6ZRnfJqY2R6g
kJhwQiGzbcTWWJq1vIY2Fvhjo81h1sQJ9YR4b+9wbYy7yZx480lWnL4AIMzTxmZU+SPmPP2vF/5K
lDefiHaAjzHMbNEOPCvfmcEcoWDxMPRdisJf1j8SVS+ISuLqgJ7Q7+wBDv9XyQstNDdT2IWBUBIE
38rPfGmXW+HfHi8KGatkcVJniHl2x9JsyZcTSpj52qFDUZQB4rJVAWdUnd/yKWlzCo/itWqCSC7p
3/pbGrhcoNZZtxLIMcUf37BBo6aOMQG5SlCGEH1oexAqrP+AwRQPw7D6CgDsU0f5AgMKM1+TL17T
dYicMZXPQ0HfVTAio+jQGXOArunRo7yon6vV5UhyIfnJ9DIgwdCFKzs2034a3kgSBoNFpcXYnsNk
s0fCn/zUgx7QAS6uQZc4Cj38gaR4DvfTXo4Yq7Tooyx57qBUGKgOE2MCNPR+BIuJ3i+Rq4DMrYVX
sYLf9yMb0mUFzGUjQkpHqwEgLiJ2sh2pFGCBIzaMLUuG0qHs6kr1QkmQDFkCDTwzU3hZz/BPpErh
hphaJOBNa5uUGzO8q0X5KN/Hp8bYl1c9aY7JlDaPYxzP2BFU5a2ZSIKYr3VxE1BoTcsa5HN/AQI4
LkpAWDkVn5c8rrdWk9p7EEQiMRKSFhnmZUrczImSeRXacN5JzWPZ0/sdKKgu5ULsU5Sphvcrb4Ud
Cs2VsTieup2VKWbf4r5X6UICjGM6Wy0SF6kprEv3sBV2jeUOXlqXYBTMfHsUeahzVQikdjLnOuBg
5eUCnDc9DRdgHPHvecb7psm0ujsU5+X83tJ8C/MYkqIZwx05icvvbo66mfOWhRtkToklJlZK3nDK
qAk2G6ACJJ442mEpZmz9nhp9MosdaCpJxEV8CMkUl0VCCxtM/dQN6XPu52z9UJNO+/IJ0OyoUQSh
t6UxXZP99CNW+mQMSfeT8nAc3Enn+wyHvM3yIQFEy2ej7wqy4FUyhSD0uS0ynjcuSz3SaFx89fgR
yyW3CWWl05VOnz4qGG4UWimyPjicyeymomh04YsXzeLIMcyiMXIlZm9gHdsZzLMDfH2zYC6GI1Vt
WAlJmBH6P6ihLL38rr8BObTZlaQkbTxnOLO4ZsUfe0fuUmS72/91PyD2+ytY95RhEoq+ribL+Suw
dJPm2+vx17rwjC+TSpxxdyJDORssvWOhF5PPy3ezhCkxmg0WdW5VDMvTSJT6oFUzs61A8XkAgBG4
77W8mER48171eSaxO2XhbQVmjZ/eV08TWg4MDfDNaEz7f18qSPUsQldBGXwHKqmHeSdEoF0dVY6o
WYxgNhMFYaiPboBym0MC8w8QpfhJh+ShaPyEzBmsT/r0VPl40t3rW/7/UkQqkIkAmIE/JSsbmeat
rD8iPdq7Z+ycvXcX8Ww3Vx1cE/4rZKrnKp+XwG5w97SEKp/vlueRIL78eE8Kbr2ifFGEaHHzjvtO
mynUk7HOI8IsULQqX98+MidRwz8/TkiaZXv6jYZ0S4x1B2qRBxdeBc3osorVHtdGxtxLBltUp5Ae
6v2mipMI0daQotU4EvymkoJicwlZ/CppMePsZ7AzkvsGIq1D7nu09Huxr2WPs8YUJF3oXmGNpvhF
Dk1PSYB0w/7bfaiFt+ftkHD0Czjn28Arq/qkSYpQo6oUiz7tkXoXZR348w8TZVv7P0gqaL8yRDaW
W1YYUpVPEQhKPpanf6xb3L0kERieoU6WF+zhiJef/VskHMfOJ6QfXEJn7NFr27kYEDjtFUG0VIi5
l7DAJA4eOwx4m4nn1+q/nbcN8xaX2Goz4ufAKLPfa83DUFYDH8HHHaStsZDoc+XQpwI2tHv6hlHG
J7scqD+2LHiuiJZFlQPUIYvamXOjtQXpWe+fQQ0QxiHzhGNHW4YYaJIzVKD9V7pSWOwzylZycxmZ
CJm9M+CRK3YqePFCcYhiWVYqrZqF9uGJJbgSCNSI5m4Hu4SlelGnnL5X9r8EuWZu9d6fhSJ6zXWw
Xw9/fgXhLkeBaq2K2FsPFwN0A78oWCNujsRuM27k/Ueiur/0bfGfLA7VraRIMre8VqurUJOoubsE
+YtavV2V6FgX6sho+1j3sRjbRb4U0PYqRZWqlB3Ut1Bo0XCdPwHeEmHBZ5Z3Y+Zjmn0oh4DudzAy
O/w4oB6zLf0JV9+4rVrKFQC4iB1eJXhrgWwtkD5ajNkT3iHwnHC+kzQoeUkwTMOsyOe6s2inTZZN
S/n66Ro9CrEMCNQzGpBjfEXkjFKSKhAvjrvDKXrLur0IUTPJiOULQe/g5z8q2qHWfPxT3SJp7mlD
K/WSaSaOXlt5Zde0yBTdWwUcUOzHhK2JB/O+jVR4tvRvfDV/EWUFPAS7LFbbWxN8rJvRBUxTVhkP
AzpNoOgF0577BsVgbMKDcoY4MzFCFfHk+rA9DXYYpb7cVMCEDv7OkAL1VNaqUang9mUd3gFtcjvg
E1UAbR33QA6zhJs7LlQT+PgJJSjQf+zZQ99PilEdWDLOpz5D240dP2PyzChTv5CCBPaNEESLmLq8
IedHtB1K1q6AstVegXsn24uj6dn5282WTrmJ4QOA7iL4eIO97rJTryVDEJZhv6p7GIQ6x7gKhL8A
4uXYuI9ZRZpLM15nLKUHq/vyChOcgU53XCwXarKWpEw5k3DroujcAi8d5wnI97ExVuxr7zWuPv+r
kah0uLj4DoNvHpijSOZ0EETNHiv0bwgdfF9jEoMXfimKXnoTzGNKi1BIv0h+/rpfjLiXmQyrlOSX
107dzGILduax5EvzBHnwneDt3ghhoTEi0lKvm4MkHqcJHG3asvVW/4WPBSqolWu4Uuy59S0xRfU0
lzn7LoA/Gm10pbkIy2exwVBDew15j4oUt9B5RvQJAm7JRKJp9XiMKhAu/E2b025MRp7VKUtCMHTS
5pi6WF3YN0dtHtBrptpSMlH8pr/Oz7V50akoGDmeDkMexIqm6nWVOpQ8QsJP/BCzWGSWECAcAqNz
7IfvkALxtW9G7Wqf2mszUqvlkSifdMn9igkqJFCCL43p27Ly0fqMHeyPNUqTxMNCievTDLDOXPzT
DgSql2/Dy2u0e+70khVEVcGWQChb7N2Pw+v/cX/CAPcHsCTM8JXtoRep1NEKUd62AGDMlo/jCd+a
L7EelA0VoKMq4GDbJbGJX3ruol/JHpq1n1T9XUttiPRmpoRJWIq6ejHO0BB9gYJ0fhM39TpuLMhW
Q8QwC0pWCSwmiw4kIiXh5nBMlCuYsLyFm3m+vVj4LQUGzpnJy3VLgu5B3BdgB5bQnius9ODOTQVA
yCTcbcNxjy+GpASlKNMk+hT6Ceo3hZGq5ELs8/6pctvnuaq/cPTCQFBeQ6KDNFjqhr/Uij561qTi
acvL05uIS/vGZ9YW3TJW49Xt9+REjCwrH61u0RXhtYA8KyczslUFDy6xU0sNklg9zXZpM8VPSj0I
rMTNV6u9vuD/8nZdGE168liq2JFOrs43gMgXhak6DiXh5v/qljCNaXV1JPIOuIzpSxHycLLNFCG9
EiaiQKvuuaRz8wZyt3kcfH1riFUpSHiJmkf8vypt1F+CIMVzuP9fBzuKqxQflC3KEcxkNMHzrK2X
xvHtHBo3Q82UsYZE+Qi0lHU0mhgOggA6RXtyJhv684MHcZSf8UJBH+3RlT7FFl/zZG3vhnsxRCVd
yqKjou2Ao1SEQx4qWfOjrYo+/DIjPxkNcxEIHELoWlOAdAImNvkJUePHTavShguc04NoNJjVDl4D
3lm8tL44mw9wWPZVXBYjuQYqYiZvEoQXo+4yN8C2xo6uriBNqu0mQnzlB5wvy8f9Q7XVJ3gq1Ahy
z9EMxhD6x6sSUxlemI6jpo331AM7cNMjsCsvgKwhrv8oR/bADJRT90X1QP5NuYz6b6gxymcotruM
DeRUc+8Us7ltDDarnAOHJSc9MI9L/cQscmbsQn7b+6nSYaT1auLT5b6eWgkDVrRlsoBVm6UeT0Z9
CKsPIbXGRzNXLGVMrMdMpHQLd/v6QiUgy3VTKN0O/38uNDKNv8gjRTKMmoFRoRkPLdSJepTJp9Zs
IvRKGxN0sgvocBKJFr/xHpwvHbo8R80xBfHuXQ/1K8/s+YCy4WeXordUuerVMMJ+xThuLOzEMLxz
qC0yRa2TvUo33Be7o7JmPrWsR9Q3cCuu41i2eRQDvbNOTCwddVC0LwzoAt7lC9Rp2RBCQM0p73jj
kyb9MWiQizgw5CRsbtAKpxxmppw5XYL+C7L+FX+/r/hUBvSXNzxu4QUnilvkmfMfv/rcARJmmoBS
cTsbVcWuiItYgUOw5NxHxhZfTJkZVKFD0guypz6N2hJia1Qroe0nzO4fyUhrem+RDmda0/tD/QTg
y6/ZOxiFEKQ30tqjH8U3oULecUMSYSFG/FgN7ok1wQm6HYYr7eVV4JAo6xTjkNaZuZB7IDcfJzQM
d3FcItptNnaO6QVGmJeWW47WHu6Do3PHXExKG61yLleYQO/tXSPMAM6eSTIk4/wL6bdDLfaH/V2N
wImlDZ+EU/nyyBQazLlSoLJ2pzPyVa0SS+4ah/hA/URU7OmdeSigetxxUp1wNfnk5O1ZhxFgqOzG
OhUMDwZWAgVgEP4h/gp+3N996YK83t4hjd1l44gEAprQLRoFQdf9UXV+Ifo70QMuvk4voPcOfVr7
ZbKFtsTC+Ya76QFQmJZQualEWsYG7QW+KOHhHNs89bGX77aYWQWwUK8KIluf6SuiQ8NF/6YqPyQd
AWOM2ZBkKBEs9EFATi7e8qYbXd2eRMGJhWC0089buzXKiUNt+C7OrlViRzIFZclrmTX1IYztNbwN
Vd4puOjxow0cMHR2PGinaZq2TExgFP9Mq29WNfIT6S79ME81NhxHLj0bW4OJDvCAPzicLTzEnXxT
J7bTKl8y2TydX+3U0fDdcLt8sPFQw7RNTD45A/RFAslZBi720OGOZMklHKaW0m7uBSMqhuQShRgg
xiqZPo0KOJsioi1csFnmeWtqCnQHIsg0iJfeIszQ/b+WSLLxlVbywYeYbGdYJErImYivhfqKyiCS
oVaHT8v+ew+mVqT/WpUFM2Lw63lGDkUxPssH3Dt+hiTblHXF0RW5U714vzo4gIy00ICZzUCjN/17
HwRWalhPrb/u/V8a9xw2+bY2MemnSWZ7PSzftlDmUaMFY+MFksWbqVt/M+usyGg0NjuPwtYiNktN
Oi5hJU3YBRr2k91KJOOAWUGrEosPS/TTxZqqOIAy00OatJWKxsm55e7IMjkGa8Y5jn89ISk1QhvW
Yacy4fI/XR+2ro9rdIuq8Xd0gfPIhsJPwCO7gW/yNfLHcokbNJmYBbGouhPriaG843HYmVLTLQbB
aAyHGX8mlmVSjA0PM4rl45GYQE/QERW9x8eULELWhrWisbNPFEB3v1XdoyyFOUSxGMY5i8+zOgGO
udvqT1TkCaZKLTBSU6fTvPiGT4Kp1FwGdjh5fYDjrz4jTIikgk4IulSTWHKwP9jbDJwGkqZ2OGUt
iRVezF7B+zEEWjWxzOG6911le7TGoSOJmi9t5VS1q3IIlKdem4zTLrOexME2nCTXDjNYCOEa22E7
KZ2RcAb9mOTr0cQNsMEgCIQTdawa/S1S2YrAkeVtD8bhvBubOmWjMurMQSrZ+5KF2DwnVWxz578V
RYVlUo9crgysTLU1hJf+Gr7okJ3pS3hTR+B3QYN42N6jpP0ypaVNXP+1ZyK5ugKueW+QmVLfNOEM
nWvqTUcOc0p6o0GNa0iVEdmyV09Y92WS6kFtLzWyfjsF/dw3j5/2s7cJNLSCPQudKFHhFnNlxFZn
MpyJggmZ9e6BFEl9oHs44mCS+X7jQapNHR63gBzTj605WTq12H6uOON/kuHU3nIsdEGB/7XascXb
4YPOMHY6Ad1zNUYybkMCUV0SMgBK6BLLESVEzcoc84iepbG/idsxCLNGTN1eUH0oYIM+N+DbYh7L
Gg0VztC5DlsLdGzDEsEvl/q77QTlIeKlMoOzsXbFQu5dxNTNdutwKs9zWKOd3CLxPf3q+h15N24y
RLbi0SxOKH5qwMG6gvURea8czSRkGBM6jaw+JUV68LKfOxfJlNL83pBYh77jPI9yosQaO8y6CdSb
uZQcIKRPNG3c+F+WSeCUt6RrG/iXoS/AOR2EFCCrkDqDlSy68EyiTnhJy7ZkjKlqdDakiK4trsfI
fxKWjesQy4KYK4Iq6We4HvE8aGeYkqlSABRwtyyjl8f1QPONBoB0Qx+ca5yXCRr23MLCr6cnhVQi
Xudmzat/gIg1emqxcz6nvFO/3ZWbnYrYYUj+QDFA8/jvYUk1YPh8oW5nCoZzBlJmxJRb2bOf9LE5
xXqsgDM2DO6duS8bygSpfsmQDvTKN2be1PM0uBGqncVdICKe3eUcAKYYx2K7s6J91KHn7V6cNGe6
+kVRWCnjVUtWdgoS8q81lp828uYgt3qfYClfuDpwQ58JF+xfxFzWX+wH4vg6DSe6uyL+azxza/pW
GRep9KD0Mk7lacgcxe1OCp5Yc3MwcX7EqPMk8RFnmznxIp49H439SyS5efl6D3UF6/AG4PGp52ik
Eye/MAz44YDz2dJmDf7Q7pAdhyWFfJRR5QvClqWqrjR6TgixOwphYLcXuUApzSytAxQ12BqLlfaN
wvPgKgmcGDJO2j4Jk7QBrlUiJADUwyUM+xb+yLbgHp+4/9gaN9yu8rZWmWeEfzPRcsFM6BfMZfXk
gJjmHE2+P6+xmWlmvF0D5eECsn/eIHmr3tHl+prS1KSFiX3kz1KbvHaw3/+g+Zm1i+VFWBgCqjku
tBortG6336OnmE1VLkrvE0aM05xrChCUvTPeRRT86vI7F18/kzI5foxEJc6YC7KCSz07RjVqw1xN
vurB18QFk47yUqCZcSvS3djhrBuFd//vv1JEfk+LUyJb4iJQQEE+RzDIHLMQgqtCelRa0dWDCEyw
jcldAzKOU3d3oHNiaK4u0eZRBZMAAIKyT6knUKwL9VWjnsuNPyEd7JNc3gn02QJeS9Z4tJX7sp7b
G12OgKJ6lnslC2u9dArFmWOA2eOnir8tMRDdCBl75E0gBBEbKKyj9XZqaVvEtYDxdqpUK3R+CRYe
PU/YgCBkjX5QAjm4pRZxNECdVCyOYyjBHQcl5rDt73I3APx//U3hXqcJd/LQqO4c/ogx3RJBucLd
DTx4wFqjnfnFQcJG0Q0blpDmfPosWaIz+fVxvByw9sZLmCW199PvTV17JyD62b+m7KTmA2rHGEC9
ZAxDejMsHbQHkNDg9yAXEu9EySvi3apFl4zR6AHiWSJhkGAnZO/FH/w0ECsNwOG/MdQ280lezluP
INKjnl/+p3smywqKyAAMQ4fBJuwzoYZviabVJcMaDtxg+VjqI0xv3DmFF2/X641Mz1yXE3Xy21bp
aqghk9867NpptILoiSxnOCBZHAZzuM0yP4d8JiCQZdWovsW/cilwnei1FiOscW/z82HUaaYya3el
lpZbAW8EyQOPL4R66puZI7sP+i7m12Kn5xQe2NDB7DLvOvPTkgB8nIWUq21TVCgEX4PHS9W/b/6Q
TlF68EFczjNOcDSb/FIEIvtOpTe9h8CgnCFhmXinwfsOxuBFLMr0ecVG8T7fFtVtUzuvjdgaGIAB
orDKJal5sSbszrtAY+I50ctmifrrLmHbTCZU9znur5J18Lz9pF+tVr0ykF3+hGeQsxyJDqOes7yW
fqbXOlY0Hx2PZTNC3K0CfUvBuV+x7jcZvWI0kSmdxMqqRDvejpbapmusRg/GCDvwUGUWJwnLkYdx
F+WK+DjMGWOAIQepQIn0iN2JBxAztv2rgW/y7nSR4TffDSBbg1iyyopmgk9A9yVnvf5DIZLxY2+V
9hbmwlzDMKrele8KVEh1vN2lCbhfuDJoB5Pf/wwg0EQ5eOZAwRzIVMOrDiFA9L81n1r7DJIcd2La
p/1s+f0aHGub648H+S/N+Illgw1ZSkj3lNnDcK0rnVsX6kYt0a/fcTMhIVXDJZ1P85wY0/Ad/ub7
HIXkD8QJopVMyAF+q14eSDR9KR/Bst3yHJslqnXMx/0ylvfNqb+Rj684wQyWAValdVmkeqsbs/4W
qdW2ykGqJ18mhHUmnrAGtj3D+fMJOoAYpaI2ZP/3qSG0wgrUIGDoh6yCiRACYTKbIN1WCuujCrps
g9iMmI38qb6OO/+lSYZxlGVzIL75AFgjLOT+exhDV3/sPeX25U2CH5GoSUMM7x2y/sC1C8aVARIn
JFNKgMrJE/3jhedev8wW4U62O/izi35/1olDPfMTJenrNzcnEmGxWg89BMIjDeSuuhz+n36jZN5O
LvKdqRgV3pOLIWL1BMppWtvZzaicCHLw93ZGZfQLqsopl0gAz7eRKZpLupUNLwJN7eYMKC7ed7vR
MHVJTaEOG/IcOq2A+3RQf96AlPr9JxBurmnGr5djUwcMZvmyhInZxPeJnSkE7D90c1sAM0Xr+GsV
hfGfRW2+/hVX/q/E1lXroM5XVrTGXr07+TyO3kus3lT/VxINONc914w99T3I6cZnlFKSkxG2477/
uigSJmDOVit3cTINFAEgipebIPGdiqRhaTT3vPuHxFpqjkBuf6UlVDd4swkAj49JvbRoBuE6uXfi
ybjQCS4AR5l5CE7V9e8AV1nSRc/yQ1lGzrvnMpLpETQhqlw9/wlHCy6a8r/QMKjh8wFz177Uzqb5
JkSSTwMCaBDjCkT/yxDtqD7tC84OeBkaPDxe7AiUMTcq83gqmLF4aezRAfVdr97zFwg8O7euBA2x
CXseDHeNL7hTMLjnPAEHFvlLeNezzqVaxlzLNPAB7C+O5IIwSRvfwBEUrnQNN+ZwR1PQOuMnHixN
1fFKhQdKKLpu9wuqYPLarRwjlNQ5czNqmtbK9A6Nvm6UUSFXjoRvj6r6D067mGfjKj98MUzyIykO
oMqAXKz/oYaDfQxhHhr7TS0TZlj68/7DRMFhKI/NtPj8orHRoKpimZZWiMoO+XkP8/LNNd5FFEtJ
CNsX9NWfVfIduewg2XvsY6+bCXgtFuqDKVXXOEm30oAEn22uEgF6OOmPRnCj2v5yg1Yn4SvT2SXX
CUybWawpHSMIPDgvZ7EZgWnwkz5XroZqil6bw6mS4b+b0XBbv57XugXiP3lH6z8bXrfBCcud4tWm
8O11NLHtLF8Ea1+H7a63WocRQ2XO67wfdryl4SrgBY7kNG3wPw1EHbOdDs2B5a0SAKtbZQodvdNX
QsMLS9RvIGTmUCUg66ebsck+cwY+afpEc0MGBgABNtViXsB79K5N8yJylFvBuxzGaJhG8sljn2Z2
QI+8PAxxlF+yN7CkBV6QKE1UW1NImcYeiHhXvR7zfFtZOu6TZFdDa4lwXrsIg4XVXJnlL9x9yIKd
LzAEwmoypj7D+95kxhnvsnlkWBtSsiRv7odP3lmmLUJZwfGBgAlg/mcm9fb/XN6zEKLGxke55U3j
6jYoRcDEKXf4MgaYDLTqVUJsP592mFjKslsMG3cXLvL4yHlZMXo6Jdl28nQd0hqWosvdWB/vXwOA
VYjV/d/X82s7Hcw8PKerZaMQDSJE96C4Z6d88decvKj64BhnWU2fYdkXM7iEeonBywUE59cY1L14
pNGI3gp8A5yhG0z2RMhJDbtMbcM3EKia9T2ncD9soQUtmUrUPopw0YB5I3l875xlHn5qcOzK3QEG
zJQAtycwsvQapmC2SseoU6Wte6BYHlJSs+kyfELTZHGSJSV6SOSnBmA9dFTn+CefJFGGFiVLqaxq
sM8sGSdU1HwtqEmvLfxlHIv/CktDu24nbDpJgNqASCckFFXv5+egnDBdQwa+MtWz4+B6gMBVsc06
pP2xAtrfHvM6jlQNgdOFaz6xawdJJqBM+m378KVms6oe48pXl2+SaxFvSDTANNhcdwy1vW4Pzfju
kHwCeEpin4ZswkcHV5cXtT+DAFSd6szbBA1+jleatFZ0n1JyrNMIixv6g2BGekdrW2FLnoiWGphL
tyRIGnO0EbIdUUWcSKVb0BUi/sOaDgNB2fHs5BdAEyY5IcYackhkZR39RLVlwbVEDYH05jJ8obHn
IXYIC7PwYuiMWmmpSKOdQNWuEmwKOaZOCqFjMOzuZi7vf5E/MRyycssLRPY2kqPxdTgq5e7Q+tAa
ZwCkZGGtKtwK+6lMJWQOVZgPAgfsEE5F0khwmpyDdtjMR3dOIz2TTIduGOknqfEksuG0ohlaL7Do
kGCY01hDKJBDX0LjEHdr+BJx8EDgCQKkPuP7dR07ygYKGw/sOkRU9FgZhuWuaNav71ab0uNR+YAW
vTt5p1orHdmRa5WzprhuyuykwqfU0JapsFVWsXY2HgLGeZRht8EOnzJ1iJFUxuDYhc3BegPESoy1
78SraP3uBlGD+Os0jAPxSxRpPfsXWDeGdOC5MJE231OPNmHNe22jGJpCnP+IunDyldeVAwGKmGWT
8TWXXxYKkqMXWYmcRUTqzmgTjrFCVQTPF2SnXZc7qJrfW5rYpYrmX9dEVWJElkdpIHofk8nP9LoI
Jbj/k397R/RX4YAsnHEg1+oiRVw3AUM4i0p/yNAVSL+Z6bhOVHZIH+qFnKwsAWXtvpubQS4EqpFt
Ve3xw3x18ohUaLWQt7lguKqs/i5yhphJOygKCku1S58Dyk0/TVQ7xU/0ivUzTHugh77xLlvckl5x
3+s8sa/9j0tFb2zjuXSxlgf3HkeJj2Yhm14G3yiNCrGVmXn30ZK7fqhqsvOwDGE8fN/t+A0Hrzov
ckSUmzeJlqos/I2vaV/rfxiG+RhJBk01BWi/07jkKzr9XUqT3SeCSupb30udKZAtRr7/lsQzQC2V
RjcIwoPRgi//cQEsGzFrtRJtq7eDW1+vUfkPHlhwGMjgknK+s/iZkEYGxKWMA64mE1Z1lACYjCEp
QePvY2JcbO/U7xfvcZvs7lk2OMulWVQfxUUOlE9xulucGTcqjAtXBd6J+vJKETvij9IdthuRRuoA
Kc/q3h9Z0qdO0EYPhmEVTA04yld68mkSBjd21h6a5dXmGEVI5ohLaUWD+9siK9F3ge/geoATUW+f
ZMjWTJvSrESCn4QxTDFxkm5X1QeCSLAQxFyyu2T1RsuvUUjgeDHcWZ8fuJvN8dZfQF1cnuj+Bqlf
aOzcjDeO4pFWoj1vA+2Sqii6IKR2SscPEIINcTSgG4MF7xpcC1oH4WuCiGsOD4fb/eQoilxCYmUf
NcYSfuOeDDLfLR9bCnW4B0UGSBIfIw4rGuIbKMxiRtDvvxy2eqEQulNQ+n0yIjCBiBVkRdXqoidz
A01ekONGie3wOlaWPPdhIzK2fYBFFWyM8xQhm5wIh3fwNNJZx4YsOY6YulHvdlFmx05t+f9rYf/V
G681Np86s2aVy7CccaXC5sVcnxzvrT1wedhxX04y7VK4XbKzEn83kHqw74c1NQvXMGNXQxnpJUrq
UxSVeXNpgZo47aKAkyQRjpz2pPZWkiZUzhiqSUTjdrH6NYSccbQI2kDnLLvTo/u87JVsgHBpqqG9
/61s0z00PYJ6+HiwQd9nJUQZmL2Sv2Z08Of76EMX93itJdywRIrwYON00fkjWp/4pI6br/LpitEN
sv218DvIR8XNARU1c8WBCQcJ3uNbDD1DbBpgsOVh0rodWtbfM9bJL0v6FbOMVs3ccgjI3iOJa56Z
sXupZ8FipQw8zsB9lcGs8AL/3njJiWqGXUqYUtgIFk3gIFxLuvP23kRBqYFFXShIv9exziCNrLdq
k+tY3/1UkbkV1fvMYLR+BRowgdRfnoFIyJBpPcEvDX6r1pA3hwFGaK8faPaEpztkX4FW9WgkcVhv
sof10h51Iosnjj7ypU0mbbZwqHKgxHQl6F/4Fx8BrJuTKednCVG01fQhOB2HzkCaC+LT4cjPgqBp
bDZYOpGviiyHw/0u31EXG8bmQVwjHFZZnFt+fV9lTK4QwZzI353uby8GtTav1U3ltDhTmGySAomj
HScjIxNLbWgV81//6F7i2+sS5bOmd773K2VkX+bsblVJBSSYbWDejkqrwYeM+tktsSvj6iJFwiIn
UNiNJycpDWciZGbYYJEIqeCKpETqXfYGsfsZtPPjZLpDwtT00a9EW7GhkWFlk1WcONiQZBE4Hu6w
Xnr5h15187NQIFwkSba0IsZ6DdsqMd8nxM64EojmViyYm/BvVjaUla8zPbaGOHdO7uNJ9T8ns2k8
IkkVuhAo7s3TU5tmNLG0UJgr7yZf69ZkMihHUPDMqrPq8caLhodByHrBc915+vuCCj/6PaFAjM7h
cvIGckYoCO7AQ/xVpHkMui1/UQb4mTNf/bX5UrBdiBES6iGdpTl7HvuPHyqPSdqLzuxf1P3LVxuL
ifZCMj1Xa53gwcS0yZfX1qR4WAU9u0nLxrHXmpqsn5y1o2r4KpX5TVaIOu+uwzSjbTTW4KLrhyKY
27yWD2+D9DH8xd10JTrLyc+L+eBT0iYYVoM4g4ifaO57EGdWBvHwlnofemBQL6nAgAqfieO60M8U
dLeMB4pU0cK7TjfITagshKA/bqLwF5cy9mOoPWeZx1iaxmBILxWe7t9RR86bho6ZlEaGeG7gTQeb
YkAmewaumEgOAVynAqiI3YJwoJNI0KC/xYyafbTM1gcJSG7xQNq/Fg5Nax9ADcqCJRLLnqu3aQ2c
qckjrDzLpdpNGm6AvzvXPwJFkrX5NJkdQbREC43h7lGD8Dlirpc34hjl/x3bongZq0Tt0unFoEs0
9Dy5v0Burr1pnYtClwJQAXfL7x9MhVrZIJjkjzYd6dVtxm9ROgdfAc2R6KIDVYN1c80ZaDqIG24D
iHN3a5y10bkwrxcWJmMkSzFvCu8yaymwClIiESePbAk5ieTuPqDXKRSwf8ldPTV14rlJTkn4t76g
kI+mdBOgFtWidx3R7VSBgpQ5AO5BC8a9QJQVLdIrTMH+hRME5KPa0iTjVy4IMh23n1smtlO06TID
1x4mcbbK1MIL/Xkyl0W6K+V7s+3XZdD1xO0zCvoVku9e7H0onyW8hZmwiETB6oEbYePS8oz9yxuq
yT5I1SJwnLSG6VWabsMqAn+gbaRoKstjmqOVJQdgyxM1v4EORNSEiZjANu4xrdxOOggoNsEQetBn
AopeVsIoJ+m0plGQ5ZFY+jhZgTCwym86HNXdco5Nf/QO0Ok9xIiWwJV7vMakeR/fP5eraCM/U5G7
CZXcvfADzxWmiqfRlvCJuFOAuzNlrJnc+ncZRf4+AOaWvMtZthXUHDRH980er2M65buT5KIPKWg3
/Zl9FFVFr3mXaayzetal1G4IOQQU2HNWsXJSr0j2MOzU04/xWjSHtJEE7M1OZBzjlMbjog6yLtv5
jc0JEXMg84H58xCNhnwoVPw1XWTZUYTTEcFpBlHqSnt/KysKVlo5AfMRGF8JurnOpxBwanXaKQ5x
nTSWTYSLy4vcpYKenRIjeFTeGQgwQvB2tv+JBJzZi2k8LTwSDcTijon6/GGCRv5nGSY8dFsL3xur
7GIi2PllKSri4He/yduw/qvu6nOztNwVYQ+HWJzuuYOe4ijFYLnPePWN0dZMQI4c2yrQqx+rcy/R
cp7aDh2Y5cJl/FRddUEDpSnZzu6DQ3RmvBY1PsNymWU+Mj2BbAoSGyn062GlpeLrku6HsEpI0lze
fSnDRW99VEUSgUIUQxQPIP/vpHzfsCr/BAlSM8iVMBXLJVic2LEqNUssjV9FZXLi2RLbKZ0afXgv
OSL2v4kc9YtAWLovqw3RNfmZDUvokY6cxpkMvN9EuBRrTlH/AAswyP/OY7jOZuY4RZv/rhHgRjf9
pKbHX5FeaOjM8pMxaBbsQnA3TYP4+WPt/0aT0wzp6WERPg3z4jNQiAa2VvJ9hJfFiqRr91fjPn01
BD4f0zAv+b9DAag16GpFgE2OQjnpooT9HVDG4lB/hcSKFNE25/W8Msq/jiyQYt+46ysFZRDGVlZF
Y7oAQptkVl9KUyxW411Sntz2jXsifXGigJUggZDP2xoJf21VBEetDBuyCUg8XMplE7uhMaBhm+wb
wnxPW1bZwT/xq5oGyz93drh7LdrZBzbt+NahJZ3RHZVBXScl7E109KPRhrEOOfM9NiJbfUSeB/KB
/ES2gT6apUVrnTVpGb4KyZ8l5X3mu0ZbnSjnCNvJW76Wyc8p7aryTihr2cC9Fwq86VkxaUXhIunm
xwX4IK4xO9vz4Oqle7a6QYl7IGWM5v3xi5KMFbxKmcgPkVlZUhiw79UyYopmn0fvY4a2EqJDM6Gc
CxFw8+uEd25j2BRyvHX/Vket5ABQBmnZAj0xn2p05A212+rjkg3yw6feCcnOuoPB0F2OnA3xuUNJ
XVWkMNLL5FHGDkmESYmf7EI1Nwh9KMHJVhph4FDzmyg3YsQl4DvUZy3qbQd73qhnl4EWX/9P9Rtt
HpkZE6YNPdvpgU1yiHyjELXNCqz4eX0BtoPAZXNAHkZYWyezvW6XUhY9BW2uDbgMU0hIaC9CKMay
5P33+sb6Uq8XAUsJw4bEsfqMe3Fdh2N5xd5Q4FvTobjXlkSSd1lG4hOTmwvHf3G8VOUqA9R5v9no
tNWyOn+qnx7r88b+uyjCUTy3xWxA7ebpmaR2K+8fVWIsUVe7yf3onCfxsDlZzXPbOSo7RAefqil6
dhY7TTXzXL2DF9L7OY0ik/bDDqkVdowZrJ/WMEQx8yyMnf8FA6uCkUWgNdYD7xodYeL5Ax3cSDL0
LG/8OkZ2mCVO4kmU8b3kesLQzzYRfWxz1nDPaaFyht97oETfWd5SEpsURdZxE4l1hDm5Cw2LfxWr
BNWPBccdqK+MAWVpR417qNHPiOCMdwtF8DuXE/E6qhK7xIzSGue8n+7jYb81/JGyHI1MD9+/y0nW
GNZNHWaG71CKO/cU08eIctIoeLHGx/9kGeA1ooMsZuPtsS2+WmsRWCrinssMFuBj2HzmoS9CNJuH
UCf6K3zjPE6GuZpDeidaaL77bc9a1xQHxQ2MS0LCLTOsbsX9vJKXw15jZDRyEY0JHqtOdFg5wmAs
191WHh9B8DglRRGeh5pj8d1u9F+OKJBXiBw9Tpi+ZGe/Zf39JdT7HcFyrtMfeL8+hGgLVNbG02hY
btNNBWF9J6E/S/P2humUgp+thiMZ5YkI49bvqqssDKScjx2pjZ2J5hyAk5rpxXpEh6oTPz247jnO
vAuEl/zhKn+Zkis0aiit1g29CbLYarH6AtGxXH9fRU9L4p1fn++luqs8pbEVoy5OOlHp73wyCmPM
O52IrbfvRUfc6kvOgw6yQSqr4t6tq8bCaUMsb1QKQ5gtpYrDKW+nuzudZkjNdtDFIfiygmrslCva
qWNkWnIEgqXybEtEMromZhxCTR1Pcrtp0Kpwkcdch5lelPiIRyrMrHKUJwsom24NN/eIfqWh58rz
HvDu3x6Av/BEpEV3Z3TK++G93aNJUo+xCW0EWEnoTaxQ4BLdHGg0Sz9ykG3ozI7uFI9uZ+kzjvs0
x1Oxpeg/Xt+hE+Ve6LpJVW580YSWys4Z7kaj7aL/1WpPZcQ9GTgY2ejI+DItORibV5NyNoYq9O8s
cyKGCYxo5irorDlGN2t/at6/skjQrqkaGLc1YCSscT/RgqyIzQM6F9cjK8c0rEpq9VDpYa+1gSl0
sOFQFc9G27V7x0UC68taa+STXek6DvKnDDSGFeGrBRriwOtNjSWGXWnLfyMAEGFUy49J6ZLCQhHh
IbzVwU7TUTyIYBAdsWC8hp9fe3Ara/FHSyI1v/U3AQX7Kqj6Qd4SLhlywaRWySL4MGas2PPsZEzm
l+qweXT6dNlJP1nL9B3x2SIxrNegghoWJA3Jm7OD1wCB8pM+3JYLVJh6AB2gGDjOGYLKEGy5+7J9
AvNnsgo8F39JHXkdPoZ8BLgkTLHkrasllrXeQXvPuONJMJhA4QfMEeHv9yD0p/qyQVYpdPKrYc+6
87E9FtSqrYlijVMSRfO+ZAxBnZuphu3OVkWYSqI99jd8i/mFl8J8G9ALy97gL2g61y5k+gNx2yGo
/nBD6l9fNvAZwY+ZiLGHw/bCCU1DCT262YrGCp3Hk06UkWuEVCYDtYm/xBsczAq6G+wCC7T38eWD
nMxDKfJqC2YW9MIkKomb9Hhx41obJ/rDIJT4/lpaNjl5vPTzgjmkPu8LbJDq3QGIV36d2LF46hUA
gScJ/WCfYd/mIvnPcXRhVyqVT/qwU9Lmp6UZkgm0YFGHBkNxk/iPvYFuI3o83ilNOFg7Ofir5Ldr
5gbTAzSkgJiF5L/7mKvp0EFHfKZkRsxPT6+xJ2AGxwMron4C/HFsNcK6PoZgLofwoKq9gTlpnX5o
cKFrrLw1UH73JZFI6dw2qiXkZOBMZAgOzOeiOkj2QBLtUnql2rOuWFVdOGI31EHIoBmOYHW6QxKX
jj6A/E2YOQsGgrEuttX/vZMNOLrLDJyx0bmjDuaIlByoHXDtLySZOUp/XZNtb4f8rqDys/Syod6R
ulXR5xXhJ1AxSYwCp9Gn2Ar03O1Vccax72dZi7MGqzk4jOR8rfCTNbp61zz1O8omMLHpOIbEG2yv
M5S+KfplT2J6mzSyy0vRI9KMpDtG16gw7Hxb8h5l2vfxQEXUi0pwpY3GVAuB1kiYU3GpNdeUgUKr
fSA0WE5zq8EMMhOFLy2tl9siL8rCEZOVr08jvAZTgLDwZM2YM6jocMzjM3zQgtX9eiUkghpROt5t
b6CtWqyx998UPrx9lBsOgwwFgnUjwHrLw4n7hzMYNjyQ5xRzCj3nV+gC4AqDJvUIqW+UKk2zLM/U
rnSbP/aMF1sOunAM1zYcbhndrebSQV6ACIQVu0EreGTS8AUijltbVOD4YzHddN5lejSbP4FOeJMa
pZXRaPj8QK3RopzO8+V4aOxT30Y4vIiL9VCeIIqRiGQSfru1ctZ6QaUyf/BLqIV+8l+iA6c1K+Wg
Q8m1ii3mfV/fUykezX0iOdrnYMpRPsPzRVBrXdFs/O2/o23qdNE5Y4T0AvsOTyogETw31TEoo9yj
Qepk1zWcPrOZ9xyc6RVQ7H4xG6lNc8RJGGdFgXyZErPL87omKF2QJOP8xf/D3w1gtMX8iAYpK4Ff
ujhDOIfxx1QsZGtOuta5pdoxmb8uvBrGv294OQgltt3N82VduJJ2IEqLcUJqm5ehwp9BHhcrbFOR
/gxaAL4v0/jUNWUqPIv3ZHuYOcS3azeNpUhZEdjWODOMqcjqsGyaw/f/1EV2FfJqxVyvR/uFwYpW
ZNQCqNdZsvcOBmDO8fGgxkUuvfvpscSxItoB/XauF7oO3SCIIlLGRCPK1gicWANf+Uub7C99Rm9+
CLhZK+9lT4u6atHuLns5kd5LrFv52D58LV75C60r72LbdibI3+ookkbrohpp4K4WcHB//99SCbSN
lCxnOeEUGasqlsORPC0SibkkMCBgxw7pPpbea72aYXd6NKwGxVnn37NGXyAD2ICRIYWEttr3AID+
cn3nSFYNde8rZsiPpI3FVmMCI4vOQTAvl52upQuAWwW+Y4pWs4SimgPgvvUXVyML8idTZi+/l8Wr
wVCnfbAeMrOEj+osv9zKcTRNTPGyaEJ4XQnlgIQWrywUcLB87ZP7Zfiy69J0GpTpSgbHfn62Q6aQ
bZd5joSEuDXZTzuQFC5+wl37Mt1BicJO5hQuz3WWiCwVVNH93JqL6ej8dVVH0zz1sY3WcxtqzbJ1
dbT6AluGDf4SjD0VdM/yUYt78bFtP++uRt/wqSSuhVSVsD5fin/m3ujEeYJ9o7NTbqvwCXjjJzGc
wUFHHnyfGBwjmBQ9PaH2oo+ad6aJoNkdwDwt1yIxOc4H8KzWBR9JWSQhKY3pZdf69QfKKUBPxewO
sYFwiwf3Sbd1s36/ldc2v7qezmpUCbolT3XdkCn9lOpiNbuU/koJ7Lt0KWSJzfa+bKQ8QmepW7IJ
LpT5ERFrRIAIlLNF89bQg5/hDnmIQsDY2sFdxuqeUhckwk8t+reTYMrhB2l3pg+4uwDzFrw0AdjV
2Gx/0hqenwZLd4BX/IE9GI2JiZ+qWWce9pPSrOb0iUW/2feseIKpeco+t6hjiN4TH8NITYvQH42Q
KDVZgjTnPCaAWkCWBpZtukBbi9dG9MiHs/7lHWELHsmHs/QQjoApLphOupPReKdTeApZo2/0GwDA
o3e0INK4KOfF4MOBjHjt4ByhAQr0uCXeShmntqfwILhy2UllFgFYqbKtdjkMMco0woPRX9B/2j7l
oLZeNyHChUIH7AtsYcOAIczqgRTWfPLxFZTLoFcXgY73bwEEGBHOphM0xBTXtV7qaX9Q7qTqMXpf
twsS7bAGQlmkmRzXGDhCBhiirF3Ik0vO6IjElFzS47VYqZQt0Kh0VNOGjvlr0HnHN2Q8NZpaEESf
0alW7JU92iVie5UcTqk75BYl0k5pNLMmTawvmMT+yeA7MwANq2xuvNCC18hqJda/f3YiFerYNe0Q
Yfk8DR402fL3EEtwz6vkT/EpZYLm6SD/AcfJldWD2ls4Zis8bU7lxDj+C91jgNLBAWvJw4+VshNI
CDzymWt1DZfAJkTR5clHzrkw3+jxu2ZTak3LpK60h6hwfDeIpv3PDiOIxX0v3UnE+Xp0aah/cSJQ
lQo/alWmnq5vUdrhnNPx4bILErL3URP19HZjsy2piTSq+PFHO0XCzSWgzUL+WX/hVkxuB5UWK8Vl
Mgl1YEGb0DnNFH3isyuvr1LW+/zlF9xioCvEDkqMrM96/X0H0snXGwATsqDTx/Jbk5xmYVWZQ0jx
3TOTbBmAtgWk+92lrd96+Cs6RV/umcgUwEyod6mGP4we70hVs40rnwELJonTYUvUe1gtzDRlnPM6
JTyqRc/a+9ZtOfByakfGVjXrvYJpKmlT1ogvFtxl2YMMYiRnaWQgIA0A3MvWvVBWhuOO1G5iAPiX
COZ57Y65l49e7IzgIbTLq4fe5j4FqgqpZK3eQp/4Rt8qdtEzRlRRlwS1vBkET1HGT/+I6E9lOl/y
9aEvOHOnO/3ksbmUhGBcRwb0ndwagHREYY1GATO7x0FGoyjl5RWHA5TXwuNUy3Egs5U1AvvlJpl5
EAFcx3ttJ5LvrFm4165S8Zk4IQ91tccHBsDnL+VXp2VRLWwpCOtWw2+mfwi1IP7BF42L1pWn0fe6
s+vCC+lAfVkOw/S81TrDWto8LsEhTdrUKYnRxoQJaoERMd89rA5Pah02vBATJuofB2F0E/uym0oC
Z7iatYXdcFNv1wcIPDzjvV4DGiHR0ablvG1kUexCf77MOxVmZFv64IvhWfiBmL2PzlhxeFy/qnXy
qJ/ZuVAlkArmaTXfSXT3UPS7KGhBY9IZmstIB8KQ2tszVcqkW4ct8jB3fOHadv1YptyTNL4U+aju
zUZ7FzGBXy0zcenLi/trmCA5KqoQqrwu8GQiA0fCh07FTzahZhjWgVQOL49IXfrP5EyOqPuFH0QJ
4IG/AWcxps4MshR+RIUmZ7Tk3w5PBzG7cT1hLyp2qN9m9vw7Xe4gLyWytxrzHS5a5oxw6YMrdAsI
naXUocZmTNyEuTjsli4Sw1ji9g0TKqiW59vNBHM2Fq6/PVFrwSIG7wnwlvAPRRzKJ38jGSYYKyfi
dSH5kd/UI17euMnZAKwjUk15X3bI+5EOsp0+mpSz/b5tsqZSxl2HYJfv9ITKNnLn3/hldCZGuMnW
hzBsIuApXahqNUuVeIHIiMKWmuhw16w2zDnEzUGKcyWVilAy0cNJkMo7zQIU+dIma0xwqT8UX0q1
IA4X3w3ufGmx/glGQBUDP8JH+6qayMfstc7yyPfI9yFwic3byVnIG7LeWKg95uM/+yYNUtqPLpyf
w5op16IABGbbSiFyqXSu43DoprOv9ez7jg1UyYWeaDJKmwellfCY4ZHSNjQjxmC3QuvWXCR30TZT
f1xvX2jZ2sps4MBWtiuiqjro81IX8x1BtIrJVAKP/xbEOKXt6o6aoUkL2DhDSQrZz8d4AHn6GWEQ
q6vFUPuuMxfn+a6MfQtdWF3bwsi1VJ04sqUnsKet+7mZAP5y+trfXQBmBxgo6PLDftHBsve9a/ct
YWZQP73FoTPM1XDv4ajK7teI1E2+Aih+V079XaOaNdwge64pPgO57OtESiR93u53vZOjhteEE1mS
tOz+1zdtnQ02LTeOmvNIEOJS+nI/BVn0sWIofAISr6bEQW7HKyp9WGWhcxBTBA4w0ag8KtumT+Oz
36MO6EJJmA0+Dack6nGYH8kLdVPqZl0OWXOEsEgyPINfV9EuwFSoVvxeGW+oz2turwStaa47LvoV
lP1fybo+DOQj+B1pSgOuQGSgA0LvOaqNx8e4CWOe0W6QGOeSl1z/hFcqKeUyP2Dz6a1SoV16rTQ9
0nXWKrCKjvljU3pYCPBNKje4O9Sj7/K56Q1XlslNO/W242Zkof/Ksa6sK4nXR4xCdJH1qiuRRD8h
sQCYL2og39/fXtcQ1nxoAHyDSf9u6z0t20sFSvUJ8JepJ0DbAAm6Klbc/tizstSrzu/AGQ6kfBh7
qiTfcha37RnxAcfuXAmOuyHSokVG+JZ4fSoe0/sd1glNgQFRJO7rhfOSh2XPPq5p0rkMisfJV9R2
zCTmy58N/vStxcCch0hn+784cTUX8MeyVuZc2GOXTvGQHqCf74pa6Ws5fGrPYoPh44Ba7D0nGUrs
9YLroMKxG0+iA0An6JnBhkdF5Tb+y4dHS8Ig4ZJtg9uLechaRf+SerCq+Cy3UnHkWRO2hPfELOfa
h+4/hRGnj+UqRKzQb427zUvfG3tJPy2SWXaUPo6d8McSdrpaoxxkzpxxc2j/iRAiLqKf5fwnsuGu
Taza1iKd4PXW2Fbd4UoLDGJj/EFTVSuxIhKafb6F9Rs7xXly8GXO4vckhHhAiZNPagat/Z5nMxAm
EED9m0S3MZBTpLTUf9nqn6E/L4U3r8IXo6uaPWtVZjfQL027EJfSeXioZgtA1aTnICzZDrkT0oX0
uZVdWaQlLMr3IixF9gu3AWU4ksYqq9dxUWuaA9kqqaGgP8pjefrXUOqwYyIctkGASQk/U1Za1m4O
t9H9Wr4/UUZQ+mZA+ZO8PYb4+KtI5T59Jf9clCBjevrqsFpIOunIqYWhY/lvZMb43tCfywviFMjL
SrusqUHMxvSfQX6ynH44uPPNmaLO7WK8LQBeMzSQGpTK7xC0aWG/s1bfjcHvqfpMiuPqS5pEEDdi
LvS9xWvdkJhH05JFqxti6rL+8i+4+eUA8go93iPez0bJc7/Mv7kEwdyqRc0WFPeISZ8bqS/6PRip
BZchkl7j+U+n11R8Ah4i5yoO6ViMvTsFsqyfdEabsswBn/0kOYkvPIdsYmszrGJY0aQZ5/19003V
MJxrWmnoEb2m+AtFzQDkSxP+Zpfs2oKxmfw+1cxEjHe2RZaKD9kdgHQkJlu7phcWeY2zeEkNL9WJ
MsZgmjIW1+/FAMzIqqe2kiMFSvPclMWt0+CTl/ZEXaJhlwrP4yGINx0LOu7Di1l532UZ2+xbBXUd
VOtYOQVEE7p7LzYewnQdmhHm95j8Z/0bdFALfgPbtRUAZU3AOiSuZRqr/wUGa45bvYBTO1BQoPod
AuuiFi2hPTpWQGf1q/0oEm+UbjDbJ5MlcxXRN9d2P2CB3XshwhT5CVFu0zwXnyTft7BkqpTGpA1b
8tIiWk0w3EyTBMupN0VbU2JD5CIGmixCBfHRgTV6tW1pfTMPK/5HieN4S9J0nfcDpLruzJbrPj/d
AQ955A/rK/S1upK7iQMDHdvkzGuH0c+Q97LWlDGMOUwSCiXKePI+mdY3Ks4Z0Ud6YfLUe8tsE7+4
uVj6OSF5sTDWM4oMM2Z8fbmBwz/dJtRIz+kfgQiKz942wbmT73WyYM7NL9EM8nSjhf4e8JdzKOg4
CXyyj55zeJrVTEA9CnTPkT9sSUxsPNE1n2RTUMnuNQC1xu9xSjfS8d/Ia31i/mhiBIaYJBWrzYPU
r2R6YecTzisf4y+rVGfnZVixF0ZQVj1Fw8OhtG4TBEKnWcy3ct1Xxe1l/OW7TtgTY9JKAIRVqJqL
4mzAvViDNoO7xABCr4TPh1uuGU3z9qX2k20tVz1mM7nT6M6F37VtnUyhnrQQRGeDGHeqfKIR/Ptw
MDl3VwCZciQ+Ez7FjnbTvcL1qL578sL8shZSwvcIhrDokRAo8JIQ5gXcmGKdJ5RJj/aJ83QLfN/a
0Frd53bDcNfQ1gR57T2Jh6J2Y3ksBqs+6FD82kLNnoj3NYR81hZs7oM0XmInB0SNUzKANWMKIZ4h
HoQcBh76xZDRFhkjC/hX+7gr74CCTXV3V8kkb2bn6Yj1dlPBNRPxmwJWylXG3lASXeqgTHTsbcZT
6nlk0ChMytvBUtGO44I1R0Qw4O0AlocP9vxJqkwaAHq1BK7hvGb+qWcMYjNb56uWcujqCsn1IeEG
nVwReSvxfiz3g4x/I1gt2xbTX6KQVRWnNGGe4tAD1rUHOCjjycxmDqwvJYzzHyWmFCAney2s91Gs
NheIu/tdF0sDWAXDr/GgS6kokNdgIP7sdUVHROLuELpurxYe9hJxDEp0tksYMBnVmkByfxQrk9Ig
PBMTi6KHz8/aE2zbBqrpPHfu7p1ADe4xsQ3GOZUa6Z86EJwCzOI+MxZK0xDDGYugscvbkvuDOnI6
GPKWJhAQfdShkHkDTDwivleL7NnB6xrxFczmbJx9qWjVDzjnjJ4EgmZaBxifP1jnJyDe7HVeW38k
IhOSwbDiDNUdAoz9kCwHJMNHprH4fUzVMvlzxTSu16LDrwnaq3zc70sBX+4HcZ95BgKDnbfB5hMC
j3lN6zNQQ+p0ZI2WwFJ+6OLcqaOT3NFskpzLdAesbJRsE8ecGLOS9C1rJJsaRbRCfPzrOcT2JCv6
7Bdrh3UnPGM38ZmDVuXlEEoyeD2JPnWH9MEYWb6EJvjVAEEMKOP9CKMFD1nQfkwUV9y82Z+Cgdqh
8Ckt+Pg8Lsq7s1rfJ/CWCflqKWMs2JLCmtArUpGsLxal+6QQWU3izElTSyW+QHDjddyRvzJtljZ6
CUfI28bqpnvgTUb9QcMBI42vtakWnSLgMNiDau2MD2KzR7OCN/vl4a5TrgKDIod5PebobI1/YmaB
NAv3zSza3eCO3jP5YSNlZuGaAzjtsVS8q+nm6inDUP7wdQvFnAGo79lk2QfGEjdtQm3/+ohyQnYN
wiVFkjKsguHlDnEEwxsMbnh/rbdtyavJAmyDJ4qG0sPQOjJ1U26SEJURikONP0pqUhwhftmzbaa2
AYJtV68UmGmCPHJUxMgQEHx9Kb9gerTZh9LlRDiq0O1IKyn/sJDk7pk0eLNcNtGT+Zl1gD736T22
L4sNyVimUCCWo9mJv+NB32Dc16fPoSurgNMXqxMTTpBEFjHmPaQW6iMu5mY93NZTbL/8Mgm7Evy/
J+zma+e84caf6W7+8338+WtNZC3o72o2Xhgmd3iaaULwck/KhW3rORuXH3/Y06soQf9fzDY1Wjni
HtDtc96kJSG0Yd+sLxSX9sbvCMWCmnBI8ju4dvLkoHunKESnjJ023BMNXkvkGOjNhZUgJpF4cDor
jgfZgH7Qqq5SS6kFqo3HKyRKJsMyjMCMqId74TU9jbsUBMjKdRu/Vb+6ZdZg5Zl+DRjhR0hCp5Wz
JWKyXUteDC+93RTaHL7IiLBnvg+4+6a1wciL0pwzWTTLlGYNOn1WHhSJVQTSKTvvKmcng7utw980
Q/6de/oD3KqvXxMLHNSFHVDjje1ShxdLrpOaXMN7qdVc0UH1Kqlp1mjvxqRWIU5g5i9UTlX+S4S8
eVAanHRwMK39NfpoYhOQuV8VYsg+rgl95a02Pk7qi2QgzwAzumqmNdIbNSodyntvF53jMFPmjWg9
f2fh8IwJZfsWNt10hvZ+LJ4+oW1GZMN4F461RWe3mvzMQ50Iei4VmnpcwM3BAJnHiphNDqCzPjzC
OipmVUhoojD2EPA/fSHHZBCNa4CtGac255g87DjvlFJrlbZwLl3BfaPdp3OFpF4Ce9sPxKp0wYNQ
qjwl2oHPp8o25pez9o3RRPebxszT6Y9a5lpnVQBoyAchIyRJjo8Ox9w09Gwe5a2rLVZrZW+MZrgy
MNVDkqWWjDGET7FpQmlM+LDqDYtWLsDd2Wh5zIBs4skH2gVaS9dgKMGbb7fSJgxQN65SlTsayxzg
X6CVMiOcp0TVFBsv1r+YZjc5yy0x/Xf37ekJ3CLAfLSABMzC0B0jX/n87IQr2TGlhCA5KrJt2AWe
dWSCcsMtrbAUNdNrIRcuQ1/0Rtcnu03Vc//ecrIbTyqIwx/IwdvKfuOgVnccMLAQgf5cbJyNp0ju
84CPDyqkE/NlXuLg0b7gcmpHJhPGtESSBYhvWGJhFs7uG9xlV+E/qCWKp3YxgBCtuFX9e4YvCV5u
fiBOj9RveXIcxy1Gf8MWaPdaLDSyXV0J9+Pt7pHp4neghlOsMtJ0d0Z9F8gqDdlq5jBKP0KFNAOV
hK+D1DLk7twHED541pjdyq+uRTK8n3h8HYjjZtZ1lfFRWvMnq+iSYeKhCAQuKJcjL2VvGMwCnjZ/
G6NUbFaKZtL0MCKhfcK5uXHe2ndfbVSiuSW+SnDqHBNzGx21B7o4Rzu7A0wS+7Wl3CqSaJ/OVCyy
gus79EbhG2EcPQhleKG1a4kTz49d/x14azisIx9Zieuqskw26004hIgSUzvt63T5n9tbqGXUNiuF
6UkXtkS5VGWHLTZUT8MRn+DS8J9+fF+iYpQ9GVpT3Zcn3416xQXu39315W1xoz1wIWQax8vOnTlB
dq2VbNIx1Fq+O2hLPIljhpD1eFEux49Q0L935IjpLCJxZPnfySZ86AdK6Dh3EOLONVhMWWNBP9C7
jVIBuVY70zw222e0SNT/syLu/tcUh1CWUXRV1N3kYbFatGkK75RJWhaykOilcxnZ3AMNQJ7Bgq+1
ImJAmQKBGQOD3yvUAPfr526ghfrOmlPh2+0ACTo1Xzu6Y4J/tYrlbFn8TIbHQFNenR/qqChwCgrP
rlPdAffYcg7BmnwftwA5SPXHPSERZ8Up+6adHayVgkhDKOfrMTTzJRJ/1t4oJt2bavvpVIfanKRL
oZLPzcwb2o5PvEqW3Ig9tlLywIf4SS/OzUaHFCvgxRt6+g1Gtg7ImK2xYKsa7UhUobm9cv20g99m
EwVcpQwzeVJuAwui1biV1OAeBPmEZnq/OP4TVBhSEHDRURnAlEXEoVkbuFtFd6P261jAv6ZvUkFR
jFhKGf6VerrGjmoGFU+MLzSl20/7oo5/+QzCpJB3ioKP9jAmg86If38pdZj0MKX15CWn+g42Lwum
Wyraran+xTjLpFoOnkdHub0C5j4nANXI44PlKFGWeEBwbETdmTu42maFvufWLoIO1pifz/inV+yN
+CUkniJiC+jH6ibYQLMy0/OOFpF8P5x1YmNwflE/YwW+8jrRjWxu1A3kvFN7+/ht5Pnt49aKk5dq
qw2h+4glBp3s+mBpTr8mEpJqzsSNVFiW9f/mn32mmsLGSOOTzzCLnq3v6NDXmbq+x1ZqIMNljgII
oZRtOY0QfiPpGr9E9ttyVLpH/55t5NeCgEfR8ulu1Ki28hD2W+RA//hAJMREU56JaMgYo8EOS+cF
bFrqv7aDYQx06evUEggcBPhAWXhZbvVmbXCgujPydN8vn7/vtRq9MOjojaYl4WIu3ng4y1wotVxc
2tAhm27tKPjNXJc36wCOEGDYd3DAgoSZefm7kdBCNQEqhsQa3+T804mXK5I2XuVKB3T6nJY9ZgIF
TmFB1lcJL6XKz3uHuA6ssZ9zarzUBQYu/ZXAr09/wO4LXuNvxogP3vbwFVK1SSUJoizcriM//+xh
DiVleLIsLt6e2RxkVFqGBAqZ0KQBzMSrJ2g2juDi8Diz1OJFW0GCzYqGTHi2zcMfFWi3a9vCxrhd
VF31TVJgS/ZdSn1kw3XtrDuzNerVCIC7XafvN2pJt+BC5b4Lk5+CWDtm4EtVgoM73VDFwPhwb4AJ
MP0neL320FLtUN3QtVpfRMaoHajBu871XkBvp2YlEFxPd/fiXGhNmkQSsdJglKF9vqG870gij03F
4KXIOlvQBPICXX248zkXVTrNscsa18RJ9MUcFAsN6IiuGMe9PdQu95B1P7ADZhwNNidfQVkRD9Rq
5F2BfSC5Swy4f90FopaMUpCB/2AXLCw1V52U8Yi5gM4gwCxEfXXbf75hAESojHYnVmnstuhoSDDP
jEt7clFxU8nY3qLIdGb/j/4CRlAHA72UKAKoHKaxgQqWTF9Z2tljzcWZsa+MyN30dpuc22yNqyF2
xfCRXf8W2Ugs3eDcQOu9a7rv9yx1enE6o8CwLE/ulLfzv/1aq8bdMIonqwMh9c7YGjdNrLMd9Eyg
m3noBpWW4mIyIN6ZbtmvfhAe8U6YP7IV6yRD4i6S4usAYz8NLI7dGSpUWKGANLrg4+yr9Nno0+C9
BXyTFU6TKrPAD39ZLdc2mrh58JyciD3jR+ph9t4B9Nyv2mYA0VzF/m+h/5P6/DOQfUPDv/Bfw9CX
waRsEXlpAAvZBb4zbehUb7muFSWszseWEoiNwFwVdJ1QhFcaw282AoaqTZ3zOcJgELgeLPSi7Agw
NKguCbZl+yekOi17G1iC0XgZ2fn9XYI9QTtU0jt3FXUCMv06waxc/RhHL8SKxX19mynKC7kkCBAc
Laa4uhtiUouC0uRQ0JKGAQi3oKarjclaO4nWsERqlKeW66JyK/j/Jjp1aHXX9jJ1SDj/noVDWiCJ
b32CZ1cq3Iwe4sdZRsevekqBu1Q1tteaEIEwJYG9sBY8cyjAfyfZZAYnIeQbQqiGJCE4sniDd358
o6tZNZu0R430QZXybL7jjr90ARIQYD33NziLwlm6wSSCyHhV2Vh9Yb83a9F8yn5XiI+c4vY3yRcN
/xEV9axeIOHB02YXb2MCISmafDu/kLb2fvszS1O03LAlg8CrbCJETlpFxBPyACwrsjZyJxOEcXHG
B4h+PEI2trV77j7WIMDx3W8LqvLz55cMGdHgMJyT+jCTN3jKnXJtCTwx9THty9T4Yv98BMHkV13O
wqxRfauyF/srA0rAVdPIzFkW41zsBTR1W72uL5ycX9p60SjL2IkbZLwZ7T65k+HjBW5C8AOUNSoU
DqqpCDmG9l12sZDD5R+abf+IlkXCGTqjAxrgb+Uv+nOXywi/r1Bt8yj6VZoXRgeKsKnQ+2xtDWXn
WPow67N6TjuzPlmNXV3sdFFcycnTXlUsve12C2b+fnuNcwQ8otiPIUDlXtBcr1eAuqptL/blSnvm
EBqfecfnN+8d3EaRd7SuK5j8pq8IDfYp8y914pUNhcp/BCeeA1IOCRur9SGYoWfyK74s4LJvluIO
tJOZ6IvyKEB/r1XnZtO8DYqDGLDe2IRAqmSgql26v4r6qRUNFnfLYVKTKYdYjSNLM3oNeNFTAoLB
QroGzEyB/uo05z+22IQwaPcVN0zReHu5kpRrhbTORCOoLf36DHHNNROT+GtZxoN7xiI8n+gH05HX
/N49qoeD3+ChzNMQFXrVoRbTizygSZnQUotPKV4Z6c3g60jG4erqlqQ2GfrcmngqQuynHh1qqw+A
p54fYmSu3tpLyS1lYPLpCEA1J32DeFHg4ffYOMRRlAgr7ZF7PIH+YEBcxgBEksP+fSv37y5ny7AV
WzLjBI0tuxRmq1x6B1F2LkwXS3GPAZc1+Q6LZ27yvBxuro3rk5WRxVkhKd80Gfw+DMCUeJYzdXOq
ZIAHY8qe5VUumrMiBebFEn5JbDCQ/PzzrBiucPinDk89/pBHsBpvEg1XtWhi6LMFSNdzrJGKV7jJ
011zkyIwqBdE7vf6hY9Vobsu/QWHDmFZq+jxVJ1qBOEHdsPza3WEpFQRV1yOoyOhO4kykFnPeAuk
JenDskATBuxUY7izFZ8G94/Rk0zXkd1nK/xty+KCcYIIll35kaaqidlTjiIEQmx7ztAY+Nd8tcz+
b5/qvv7x2k1f4hXhImmhGLPChk8FM9TfXiXl1g2r8kEbh9hPGvmFpwTOsCdRyaprayKmcbpXKwOH
at1PCiD9vLOxjm52396jYR7ywi1VkMPlek90qJ9IVO6wXk2IHmroCzOQCCA306a4NagBJ1ZqeQq8
iel13pJshZfgwde9RCA5w0QEEj+SXZusxXe0hzaziDtESbJM8s5O/76u+GtKWp6gAl5uNBqz+Ymx
Dq7l+5f+2cpgsVb2Lxr3cj4r/9J+va9Fj6vvXGQcUnZcnK+xWelrR7hfITz5MRrgaulLESy7nqIM
9qeqsT2vajWYEp3PFUaN+L0Eyfi49+Cywpt5lWedGskQPZo4lNHzNli6iI5UciBLKgfnloR3z0Yc
tpVrQZEg7Stc83dzNA2HwcCkowhhJ8m8daU1x6NLnSTpLDVdJNBzAFQfqDW++H/OjZIHQz/7PymG
V9wTecnb0CEDIGY9WJpDJ6aW2I+6cf10h4iWZckv6wn5/I8SIaOIlbAabbTyiPWwN3xUM7k1jC7d
CTwhbGXUbC+pYKicumMsIrSQlNHr6snw9qq5ybvtj0Y5W1lLPi4kO6clcZYzeOvdwwDsgkPMQhOG
21tupMxy5K6kZuslopHtgAoLaC/D2AsKLOAeXaOQ50ybqc9FO/9dmoCy0k1QgCu+uqkdPcLG2hBc
h0b5YArjtTH0iPj/zY2OBhzrigJ78Fq7S9fmRUX+kTb6Hyk9cryY4G+dnaw025rQfE92ksGXn0Lk
hjI/mUNJbS8qB7pBVA9JJOo+IS09S/AbQ7ZtL2ADviUBdGu8FX0Zl3CSRnkwW7TijexTS5LWM22X
/1tMiJ04FnftXZ8/GyFCPtiVTKYCAobY0rXEFd7Uf0g1AI9KgsZstkjMdrmmffpkImfYBJ7bnS2/
wv442/llUqy9TdDdi84EUrtSN+EHFH+qWwsbLqFhBKYWrNqV6khOxZF8zYIfgDBAh+P4XxoiWDHk
YDx3Rce5LhoC9GtT+eaTtggu+s5uk9qTw1CylyKVCZTOjGwUR3a8FZZDXcpsnlTZisu301UqvGsS
b/SvHSsdFsNmzdiPAuIbaFQ6IcWZcLq9ztDspaAc106AI1KzZPBdS6WVuRebMGP6dAnWwdGja3Xt
IZ35a5tzJhXrVDhEPeZ0INABt+2zUK4IFIAUZX96YwrudFoSnR/ibdNFZ807P+Aq7gDHm588bESQ
ljqUhzpuR6s0rlWwFLLNf8FcytafO38mSGnWKeKdzalxnvGlGHNR0GtJOQWEC7muw49dOnnB/8xz
Cwd0OUSU0D7v1fRM1RPS6NIJ5gw/BM92QNOU92h+0RtTLvmNf/M+pPFGBHpljHHGsV5O7mGCB/Jb
PJboa8aO2hNKaPeiiPLZLOLJFIyD1iRHyICu9JegeA6X+ywfmg+T2mhl9YazvgY23PmG6s3HR/TC
7HncxjvMtjAZKdoZ3GJ5kITw6dzycusKUCxQHjq7Jq+Qn/l66ob05bTIKCHE3MnKZO3/C0gBhjN3
MKsL9u7xlHYxrrXIhzpeHHjLia5FlflVLKL6GayY8ABe46SJbq41ECDss9IihenQdrwSLLEpjOTN
b2pkI+sdjnd1ztwuWXNYWsGrXgputyPvJ0V+fXCpX3JMm8bZI1WJ2HTMjSRFhmA8PbhPGjdzWB5L
g/ZR3xI1qv+8hoi9VlYj5PsUFvi8/NPyWeh/xE44mReclyoVzqF8W5jaWco6FftoVOFrjWmdX7GN
JdNDt9gRgcMc62Y+yeFREzqQ4uki7M97y4drdHuY8oFzMj4LUNMsIOLiAHA1/vIaAhIz7b59k0q6
Bg94m96jpf4BoBKPBCL2nXZr2pZ+rcvtNbbHrNLJnnp1OtrT70xI4Fu4qAi/ZGjXSUql6SNEn5cw
nCzbgZQi4kMboCAe2QEHIF0R4C2Rm3p2bTId3ixzUgJuZWnQ4WkS7J0fZZgZxTxJbGT14GnodHaF
Klps0PhEmK6d92hGYr4zy3ao/9lCM8tgMnQP6L9sjpYIJ6z4Y0zR0XzGT0wxep6uHAeGNKIgxWTe
QEsFESEfCSTc979FbVjtEqWxuhhYMSmelQZ3sIhl4RRjJHydQPEOnYmSmNqTjBXw0HAZKblAu//7
P2pB3EsCh5bFjrn0s/iIgsl3h7lKStwr8mdFhd7ssHU4zwNQg2HTGEx6BpCl871o6bikQjYmP6lo
2wxZnWCS+tYUV1QpPesdClmPJZr7rqyx8CnLo2xsLPUW0bCizWMpUgezxVW5awOizL6OWHvHUYPF
4TJZxU52m/Vk7En3WlDVG8iQYuj1RHofiXikOy/Df0m6VJ0uCqkQJEkl075LWL68KwVtwYflLaiX
ouYGKVEOYsuUHOSaV6KUWKB6w95FIy78rm3FxD5T+GGfwsm05cczHbAjIlJmHDRElzWgUpFYh6MD
4r4jn8rqvijv6MqNcjezPtW8I1SnT/CmKOEW70PxgUFeTtwSn2gi8pN0tH3V35Yq3z3hDprMOPvy
oXme5IeLSmcn/OB0gsnVtIYzs+6nLNfgk8RNtYWBFu0sWVqPYgniHS93vsbsPxhEi6TgPa2008sU
4sTwIokN3z95j7YnHvRX5rA2CmmV4Izj7Deqq0kTDBb1P0Pwp3f1rwgje6QblzmGzYHUebVHUD98
UeaJQ044r92VgJhXP50bnpG0pC8NsiaAxyJUYcClUAXrZ9HWIc9aO/cCxy/WP9HB39ZKWFvK3NMU
379VoyMkftqQHWVdQmfaSYk3aRqVVvwm2gHu+e3ePiglHfcfwHLWo7+OR4nZLJyrBnUDd59Hg+y+
BFyMLD3iDKPGv6ijCn+AQU57V3THoIiXl3uV/4eN4Afq3gjQkASCmdaROOEnMRoSnA//sUCFuIid
7uTVu0nf3HSBkdq69b1v9yA8InEiOpeWgwe2fkEs8TlfxU4fZ710u4zaBUY3TYI4LT57uv3m79BF
Lk0Z7k1rs4lxkvy/huIgUS2mXFAEMuBS+I7qT0gm/VpkGSB/URgi6VROO3nUqzkl3K63Tr7o8odh
QWA5e2CcWpRVZWNDP05yP0/hDYPgQ0C2gScuCfmSNtx2yvhYh5cdNxVdDGTz1FILYYOIxQuTAj7s
jcxhS4azGaGNQxz6h5kA26NzDpPHKHVcQ+QKmSIPop/C6PBbK07Kt2xuTbO3rfmwLTKwepmAmXGh
RPDv0kT2JVoPxMCcmN41pD1bnZRp1QnBGoZccL0910br0nlrBWjfky5OcAP1ca8vmjR5D2fdgWnj
XNO/2GT/cII/bCNZJXtNXpYjNxVPzKGy0K9YfVmIH2HQ6hhWJMCM+9OgOHrBp6MPJi4qNtDANLQy
akmh6z5Y3sB4WCueJHnTZsnj0tOcmAmb2UrFAQiFPt80/sj1984QVdsT8gHLNNEE1ugRo/BE5+oA
cFs5Lp/Cya/d+2ocxLJkMA9KLIg7ibkiF47wm8t/7hwzzBgBmrIF9cLHRwkzKd6xhj4QZ9o9RFfq
NVU1GhzojI8SuL7Xl9nRWwaepffNAvImfGtOfv2u605dGkTa7aQ7iTbioUn8l4HO9oWlCHlR3Z8K
CzB3d08g429cSLhuIdcWy0e3ZP/hYgFRjDrNT2vGugtSjQo+yW06ct4qjZyiBHU9iojCZWq+8mCH
CsgFlVOpVpFvH70ACAfxAMf/j6phefTJvEMj+NkYAwEz9C7k669jiF+LmuFYAH+9upasHai3jNwf
QEWAWGWu9V5nNP289SLmoLDzbqzNvnouPzWFIIaR4ZBa+hqnkNYD3FUNIh/KUKmjx6jIGNQCBTa1
qwqHOYb3BAk6NqGtapVJdDcmxixX7v0pcZUyLM4WzrzPQOvTXNeG2fbF7CSA9I+NoOjXLvx7km33
k0wOl4XYuD9lHMB6JIRlZZoprYVsrSmf5q7OBEAkumQsrgTZyNMqOXe+8LGs32o6ymTw7q9P6QZp
YCL51g3Eb+0ZgXnS2mtxKaxHFu6HrWUYwHgpAG8dkoQUU6M1gHMKCeEShUyP80SqnuvS1Di/y8Ss
uaL+NrI12kpMjayId3Nf3NKfE/xV96KSvsonkI6TBxA2QhtYmTFSa3rtNC7Nt6fYjP1POvqA8Eee
7eOqE4E4JCInh0HNWz5gsUG2qvhWofodNJZbD+DS0FtHuavzR6j534F0ZpFyiK0c0z76MY2qlNeG
PuzV3R9omTbR07mJc5H/rRKTIc8XZHGdTS5zZRnElLcWxLatXiM257sK/P0+jVAt2ZmD4Tz5rRHO
rDQIwZM/yKi60QuywZyw7JC5hisLB40gaed0nifP0q+tvJVjs7q180z+vpySSZ0VO5iwegiIMe5Y
5ruYskHk5rsC1dUGvGIMub/XzBu3lX4ww5mu0qzBzPirQ1gwWz8pk04gGdwq/simGcH30tR0aKsr
coaddtVAlpPTBDsc5RcUmgCJVRZhja2r3d6GyOzf7CXJ3KEivwQ1tdioShmsHQC46gjcodH0PwBo
AQRS8WaFizVq9ftD8GnuAKXKkgm4W2ko0xI+2LU7H+hvJ+laUl2lFwqxiEanHYMa+CrHs8JArWSm
zOpgFhjxuVYTRzNJlJL3Yt/C3IVkS7ZVg1MGNpjLvwXkwAoEU827nT7KeXLan/UG/ypsJRmG7LYA
3K/eIsZd6RyB/YolJqq3kw9TP/681+s1HJN9UF8tOvtZ6RWywqB4KDraGqZF2vGHdvDgHNGxCVqT
e1bWLWKgfj0QGoBnN1g1teidBJrSy2v0Ttq0PV3eq9yis0BTa6rVhMoSxClEsklf2YYmHUpRZisO
+AEuAGa96VzY3OjC54b5K1qzGSf+lrwJC05oKpEQa1gOWLS53R1Ts9Kb+kZ/STUjx22+u2cwbq4X
Jp3La7zKXNUSWp+S+iopeqGWplrUAuEtFxTGk33mYQQYJf+vXL+3lNfwT8UiEv8blW3cEwrpEZb1
Ds3BAcDsQETw0yU7smMDn2Cm2SM4DBkLg0FbOkyiakUtHe0LUQefjoK/l+aHsNOwlz24kRPrxT2i
iIyUexC7HEXB0sCLVcDDyVnJCfk6iSHJjeVFiQuUFuIC585vOKKZ2WwTAOyFbuBVRAYcETdn031d
U3bj26euetY3klfojoeyvWseqBkkNa7WhW/p+RZTrquXba95SRphllZi+bpWWBN72M7SVaBo0GQe
ep418aY0UsMTaHeg/v94VjTaBEes0ZAcesQyaxVYPVE5LXpKPwYjWUWLNhuQ340BratU7VG09BTo
3OJTHmNVER7NbjunzN0hmEC3KvedRarfSjnvnnhP9cDGXIi8GeVGWcMyCiUQhxj1Z3yiTNlVMJ6O
hoL02sBvZXQN45SGW1wtC+6SD+o/0tINEPtgTkbo/LqB1lM+Odp4B0c5+JP3LFvKR5oM9Vo4YU0h
B48PwAy1eUlcv4nVf9X2XuzDxPZnoARnkzqir0521e9h4pNOdoLrFT/xvB6Ni35OO8635Tp/1+tK
NIrSNgM1qz0TX/9pUcmQLujtPgBuecOO7/X+caYpoAWj/uAforZJX31+sLgYrcoP8s0Is0F+tAbO
t1mNZMYsvatjc6F/P3Z/Hvk0uPiuOv2X2znJUzOujA8ElwAzRntXzpTQlfPDd8VGV7rexCw8UaTj
PHLQW1eLvOwJ7vgA9QRFCQYn4AKVyOg0hMjRyX7Z2UzehxcXpc1gCUUOx7hb6aYeIfyw5WnU1z4X
F1MiqdKapcR2nYaYe1Sy9owW1daNi9KDh92tQOOpNB2KPPSR1eCxeWmHv4nops3fC9KAnsPCWfbC
ikWHkObzIvlvhFWCHn9Ri6fmStS+njG6vCGnNqmUJN7aQDWiE7Knk2KsCwNM1B7q81JGA2hGll6u
cluxJjOSruLu3PpWdsA4teuONPyOHJb2uDi59LJ2zqgwWiGV5LCVSNVCxWerv3iPFZxR37yohQaD
IJ5T8ewBvMUMb+ZuSoktP17yK/ImrQzfNh7bVWpyEKHUVEAAsr9Z1tAMlciRnrRlhDUzyeDG+Vyg
CloSg8RwEq6H7YP0PlhzNsAsV+jGxVMPs11Nd7k1pHLsVf0nl0UIXooKiayi5hTNNJ7lXMMeAVjQ
rY/meH5Lr/NW39tjCA/DkuqCFxKgXaZBxdoAql7obzQHJzgSDitrnxXKPkACgXc9cNcgQ1/lEe1D
dGBbYqnI+l51QSfo6kBEpwuV6TQz12MwrtoeReSYdRNkXdUkkvyZYbJZ+6bu89w39pjR1EuMuRtr
emKgUYUEamiVYPprzskj7zZ79r8E2O/ePAPV5wyOD2cn3Lo4fyBMeZeT0GAbQArtBB0WY7UHNkpa
jdr60MdH8gyda7M2cmE3wVKRbNAbd3BJTQCfzOTbuJmcg/uFzlTqJdzp55Y/kUFq/ryk1MVaIp41
F8FdgZz/7O+mvzTQG8wsPxu5GQlKz/sVxQqkRTVkjubMR0wVGx2oOAACC0ecI0c07I9BAwEjih1f
H8A46Dhhtp2t+Xx+xsEf/DvpIOKDa+kgx/dfQ+d4yllA3ABORHd9OAwsKS1WrYiw62CNRO0U/bmM
OaU2c2H5Ijunt6M90Q1nh4bn+9/Px2afG/MsMMcYx7QNf1TXdS7TlOZaelNQC4KWr1c/elphZ/DF
TkC8Qz7C2qTL7FUwni2DAr7DNGUAVBPS8UVHHbiiEx8bbZ2VxjzR2VsiSCXJ6EeK/wYei2aWkePH
bUFyG0CwTyGWdI7tod0eBTrv5m2AZger73qdtJGw2nH0OTQD0ATa02p2DXaOEaETx/5NlBoTQThH
WV7dYYExUSyIOJspu9v5tumpNZz0dAijAbvjzRXE1B0fFr6YrflrQp9SCervcmE+U1jDD3NnNxPi
EnUqTcPhHNLHvn6WtA7Yiwh1ZCLl6+Kv1tO5RrDuOzDnTG0r1nW3CZ8Mzhr+fKO4rptaLt1o/D6f
O0kJWhcQ1GPPgw4IpHtmPQ5tND3yQLdRH9oJocbm67gKJFYWpcjVXkP0hUCerx1AuN18f5l8GQ5Q
teNI3CIDdiQ28Kt1xGNQLi2KwbAmMxOVw1erAcf6EGSKaMyr/fQJ9Owue7u92rMg1xo2kl5Eebbl
3YVXsGIbnqQJ9aOgNGnoEIG+Q3AnqMSaciH/EIYxxd3jgthAmKGKcpuvqMAYLp/Mm3X1YDIk8Hke
mGcK5VyM9baN+Obwx6eDPlKcNYDqt/ZQ2BtFsFPd1Xe5i6n5PZ88hg32ZNq/Cf+gT0jO0KFKl977
kwMkXrQLTj9fSXQN4Dcu1xWg7JYFthV/lECIpKiTKOgpu+u6wq8sJ8j3FBUNGqX+4CBrpAyqiCTA
IkkOY4neAlVtfNunIcpg8gha8TIaSlvuJhiFvWsGukno6sv55CeCeJNgZXobufqopllD4hqTbd5f
9wEOQWSA76npXYHP2LVlsz+0BNOdpXaZqpgvvjB5nSY/rB0GWcwZ5Hh+ybL8FVeXHaAV4g/4LdWX
qwqIZe8tQL9JHPhcDNq69BKyHJlo9juVbO4bWiCdLBtfS7Dbqi6JELIByK6B1ebsHrKUkV3v+2es
Nw04wA2xTya5FTCGlUdgXZ+56mpHEKDhiKpVJvupiF3t9y7kRwUQoM0RDlZhT7/LmSjQJgujOrSG
qcHwEEgOVRAqqKNveu/EfKNid+I0TMOCqaVS+abu0hLcA7eHhRPCb1XJ34gUSibiJ/OH/7inFGj0
sKdPSb5TUdCPToeMfshlk1uI2TnDvyaXS6OuBTJ80ryJFRl2Uxyzuj7wqHGtq2nrB8pGty7eEzoj
0a+ZjxNwWcM1HZWN3dLF4K2wHT2m+0udyFfOCEVm1FFpD3bpRTgz5ZlS9uQq5FqDVfdZWWiNAjd0
yMGyF+P0rmbSBQJvMQI0JbB86bSwGcmhD0FhRrzZoOsP4AS+3n+7+cZjiAvwEyT6g5y1JjmDK/D6
I3d4d7bECOidIJqLy/RMe8TcMlxrM9qbdSN3ZN5mwYDXOj8ensbYhYmwf0rILZPI2hnYHb7OYA7C
xFU2or2eXfsv30VZHtda/hvwZ9olpBkiB6QDmzHbOGYlEs5LJcIBeq50g06XGFEqEwO49nDbYWOS
8a7nksRcVHtqLDmnZLWECKztplU5zLrVQOyNmqRbesIwjHQpsIrBTyShgXCvoY7h6OyBOIzjqJpF
77lis7KCo8WnkBBu55bSa/D/0Xg6ug25eWAlKwlym/sVG3LYdOC0PEz+NLeXIS2Coavv319/YeD/
YMgpwHCI+dV58dO9o/1cJLpdnp9uutUDmzOrazQppb3B0e61C39YP9Xfaujc9ji5lA3hhUeKZ/QR
8wP+0E9nbk493+26ScDhlqIdgI3g5ENbWfNZnj5TWiOI4A41w4fcZ/1zO1XVS33NGDwQsWeUXxHR
Ntq/baz8ZRnyyVMiexUrYL+HkYY8VmBkO0JHRyXRZfhxnRAkMY9oCzTN7aJp7F4vLn3UJSZbfQFA
Xn5yx8mY6Zxi+t8/6TUPKenTeyM7th/k4cb2vTkc4n5EsYq7hx0JlRFK/8Zyw9h7QNeudVwW0cJo
zyO/1YeWrJnpE8BJ821CfAVgJ7Hd5gwGoH+Nr6CPzf3H5XyG+kWGoJRxVb4hMLFrxspYk7KTIAdr
+My6msrIUWRyvOJqi94wQ3xtbEzMns6gtvySKMSX/YBx0ZRazVIyB8sNHCvVYctbVa+ZH0eLRjBv
QFcfcOD0EDXd9cwScVh2igvMEpLPIApc5NsuK6KlB6CvoySc9Qmyo5l+menq1acWhVGlxY4EPviI
nUQZLSrCxWSPb9NutbT2j142CaBT5UbSDMNDguUpcZ9DqZJ8b+v5ME+k0LZLiEcU6w17Jsf4IrZe
nrJuaEXHlhiPzgBGKzhDjizctj+IAuMo+vTgapsP1xtJxhhmwlxhiqGNvFpGBIzN3HwhCqmVFxqN
xpsJ+gC50TykxqFh0j0t8OlIke2Azn5gJGdRtvOq2DJH1X8oDSR82LsYEH0JUy4C08q1yqGxSpEj
ARfcq2Z+jSxjAAWfdvBtkvcduHy/r5jQkdUHWl0coL1wAw0ZMzrU75Fz0M+t2BRwSHYM3mikPYtH
xZmtjkq2MfGrGh7qHk4vd1NOe4C0/uyBMbPYYZhOoMkVM/uGgHsxF4xNz92fmym2X+uAAhaiqUHT
vf7Jv5OAaUfr9THPG3VyzuHZtt8UOobi2gXJXsx+rm7rlAg7cl5IOGZmrAb+IdRXwx1j4jyhBkC7
WIMbJA6Z71/3wNv/9H9ByBa8dkaVkDbSbAwYkVBjHwuUMjzPZLk82LXeC7jAh7q2y3Pia7vHL6Ex
HbCdYHFQU87vqVQW1AV1E5+a2ITNPH8BP1mTHknctcM5nl39+JFopKnHN75hiGA1hmwZxJ7EOe3U
Lb1/pQln6nCrbKRcMqIcNB252GOh8uMEtkEChKmE4LZo7hul4zB8maxhMMaD02q3SkvGQKGat8rQ
BZYN3H9p0L1cHNYTyC5gZ8r4+Y2gsIjSkl5Felrl51hmKqrl9KopROy+j0BuvgTWoeRvtmbZnI/5
jbVDim3l0szFsWYoQ40VnCPmItcMUJ5ED65s3i9K+HJ2dFE8alXg77Kvo6nYFQ7lr5Ijv9OLObsK
Azug9ahdgLE4hKdZtkuWwp3/4EjtOuTajkoGoQ42KdCeeLHODMEQvCiECYa21oKSzqyJW8wc4+vD
wjSVInfQyHUXF8bWvPDdx0Lq3J/fyWPlzI9eLUYFuvbRUwXOrLExwTqyoyYv8umSMzjEkmznA+8N
UWFAxn/x9RqYeQcMHpR/RwJTVePQCMkxdUB1MWCJ4NcMTSbvd2KThkSa23G3gy6m7j4oFfSAIX63
gJXq8/Pyj1mqiv5jBUfTVVon+f8eD4lkgpYvgnHpbiFiPkfP2B+YDXU032SWDPdpgTxoqhgciKXc
E6lylFfVNbljxEkbxxbQOQVcv6Fu9metMn/Bb3t01DwFVAOyTLU3w4WeelV52BImi5jw6TCs98zP
sBwpWy7XgcNPmyaVJai9DQbw9Pn8jDTJlah2yuodE9Lq5q7W6JOqYZadP/LiOXzkuQ0pNFa8ouBe
O4egRGZ7CmxoygZy2lzeXxAO7dr/JcZlVRBsJ9kYavKr0H0zgwGNmb9coSH6VQJNvYUGVj6sb+K5
X91eljNy5CSwPVVPDGMhHDuixIl39Ywpfy8l1B9JjyZohUmagvUluV2Ir+ge6/SVCNRU5uaHYm8r
dmbylWJ1ztjLlGqnFIvHSZ29CD83vVMimzBM9xEt6V+oBp03mmrecFlSZs94PSTOWnUAowohOrIY
vvyKBXuceEXpSF4eiUpAE4ncGBGGa3bwraSnrestzHUAd/wKozCRKfPrveKGcN8pweXkYDvf6o/u
r0erYHpI1XpCQWQj+jv93MhGlECOM2F94a/ranTi86Sq/5WEJbSBt+PyPEi7b3SXtAn3lFKdsuHw
q+UP7cODQ9RPIzJw99LvxLAquTzdqsYYSXJi1DLxY6nIOT7v+viXI2S+M/LwrmLrPBbN4l5ZIuki
8jEI7H2x9sCCBkUQHR/3Ibi0kfLSlC96SrB5NA+PANW1DQ9+rfCP88oheiFzyo/fEDvz0jG2meze
2qfkvt1Y6qMx2tweJ+D9nV1jyota5x64WBC7tZwVyLGNVsCUoG5tx7p/BxMrHIOxh/w4iMKotwBj
inkZJPyX68h7zW3iX67IclIusqPamxuJzIWWUx5JZBv45zJGJGUPFQBqEyrxHf9TicLVOrRXk2rJ
+JwN25ub9s5ZQhMdaG4C7ofAlGv1xrUvvmNHKwcAiMvBbSvuOF8ItkWdGd45QJgv1zv9rToAxttz
/5pBeR5re3qdZf2DqCQn+IT+nPdo9s9hm3z7WAqddoqHKG4vVbEzlvBA0qOAMcnC+ZPsPJrYcIpx
7a+OGIfcRvdbN5wlEwFyEmEYDeVUCI6/vvRhABWZGcZeIXIRrWpMzYuzyDmRMbe3j8w05KAngjmT
l5qTf2XTg4O21G1n3iD8gUMrMdb0EhOrp15XXoZOWfPrv7uVFtwvJl7zsNvZpzT2RWQvNWc2BITU
OuAVHfU+/rF2iD7geAjg84GZjHQfjrYlh5mIJXlB2uiZIr2v+dWAAkLYXbOIfUQ6shRwSN/Eh6O0
OUEDhVzM34kWDmyHbVibjNJhzKA0WLYYH4rUSY3iDIQ/HVvceRH074zo5ZC9evOnQmKrD8Pr9+uD
nrOZQRyjKP4+CjhrmpqvQPtdSQ43H0dy+Ffu9qwQ6owVxQDmi+ip3WmXXGLN1dTPHMyL2wLghfDe
fH6N2MHMGZiSS4myDv+NjVZlhog6mxzRFE9KTcJBa6/Qh3+pjVxwQbk9ikxkv76LbKTSOuIeQrpz
/nNTTMZ9fUg+WApUbcqweSXEIVmIRZDUolpjXQCIWlOYW19QoQJDjO/OA8c/ZoHVFcTPj1mKDkDD
cNtF/uYJiteISUqkKjBI8gzNdRlFsSZXCC9fGFjHig2e3w01FMyCRiHqgCYNhAzqmfFqUtJ9h/8J
F6ISCIf2zL08DvQOtIiuRCnaXQwYa66sff3K70W8u21aqnCt7gysmi4wC8TUM/3/ZWxxCwvv5X8d
/WdjMegwdSkAfXfGoRKtZrLZ/YtKTGUUWTQW5TaOxZWNKGm1hnjXx37c3ECm1jvZzUAzoe5r1KAF
W/ymXHryFW+x7xhsfh6ptQs2po9cIgLLOu+ZPUkSH0A5bYqZt31bQq2WJ+AuxF+t+rU/d2q/IGdS
x0IXurumeu+5ImRVTfSWnEQMQIQKoI9R5VCuS5y6e9GN2Zt6rF1OyG+wTpT1H5ydoYqxTzTU1qp/
pPVcdKW2Vc9zQESGcu8jCsEAv20hKtZxosIf3FfsHr0UU40Wv2TRfQbO+Fzn/DNPQKP6ruVG2yGK
R3IJVkZi7SOclTucuk687bN3cNzLOIZdW4e3ib1F85H7yroVx//DWQm2muFDF5bL07wlp0sIt8mM
vuElXkJUzhxfTxqdK0UBPZ/5zDOcAzvIKx1St86axCq+Ve0IeNYF/2rjl6fzaDda+Sbi/2HRDIMb
1PlGUsFxaysqR2cvtTeALpJ38XwEJJe5v3vs3R0zft687Hf6IrbDBwLrubQbQO3fPmNSqAdtUG40
dr+8zYaNu+cJuJ3jLSCCJ+3h1ZAZpW/rA3QWE0wW6UtGaglGHIr6yd+Ni1Qb3w5QcT9ejSUP7/a9
/KgWSd97Bvk2j/921D2nsBaU3FEN+0PEZrz+R68P2W2d+TW4hebZIuTsj6+xfewFiUt2keNFeDof
MkYStfb9CqelNaJARLkbuAXFmJISn6RY2FbC1AU3uanAqSFZYnoyx6GiIcw6axkG37te5/4+/bFb
6PMbkbom4GikcxqI9tNQWPEcBwGTW9ghywEKS0jjnfCSFgpO/4p3BKWElkRApuNkjbUjfk8sh+/M
AlbHdw9dWvK8qDqUu6k5KXlW8pAs9yWGAgXxTPok7jjhIAX6aRJVdlfr6IjcDqEf8Nd+CXXJippe
cBgP7QNZpJqy/ruys4HfxE40fgZmpkzTOG+501qX7ZlfpJhoaNG/Rvsfrip+zGcSjVOLOemMkOdM
e/oqRi7Z/sRXEmo/97sVZW5N61nkml5aZmCTyYVWisSeVEul6L8nvOn2rXyeiCgXTePAqt7FNQGw
oAmpxGSYeUmGh43BxOGHdXv7Anf+/icbLYj5aNei3MN5wQE1IPCVxrLKjZfSSi04HGas2ZOexc0k
8gbm/M3ArVSbXwUcI5ULJwWw2pfU8T3XZUOQ+Ovqe2Q9jH9kwK3EywWLeyn2iWNoXijQVCfObJKT
szYHWaq8ieXDQCgbpbRkzhj5DHhkssGfUHdntEotSekCC4ASJkShUaMHC5h+0xWYr+qkts76NwNf
FxxMKYJQAcWtUbkB8/FVbjRd9LnoWeDpe7knpN4mnlwS3pq55eb6KExGQ+31c8g6a2D2QgIZw4Mf
xeqTU8xhbmKF49AVPhtC76aAx5LQh36skMWY0975niA4WzzV592uESXUa/mFZH5t3OXN2Vf7JqIh
IqRUNrmjfwvfnaav0Nd5of8FdE3Br8arOww2UYTb3tfFbWP/EQA4KLLSgsa6ouhbtPMTjl01zdxI
9Dns5cDWKjVqKFGQPfVfVGNPTfbI4ismvYJaP5CY4VaRSXa/RCLC8pvwGee8eO/vL3nvLmumzyYZ
KmVo/DRpLtjX4xUa7HB51b+JbHOZryM6250u5I2VbngmC+eoadabuhUWKSuwiB+U3b58IzSVWPmX
TK+qSYb4GDmX4+g3eBKWtH27pYJ9UtBNreQt3ZKry1gc7oueOB/ESbF8a/8VlmYMIbdSNKXyJcMB
0U7USwe6rfkLsJRuMGZo17Fo75gu2kWdASO5ShUKFYU+J5QJFjsF1X6u3Gfy6DBKxrd4iUq+pkl5
uVler6FHqQ2tNlAfNxqh39WWHs0xNSxvK7xW8RLvsFIAIdR268CnmVW9GnjR0iHNigRG7qjUtP/S
fC+/OI/x7YeA4z6zB/znP76w6sY5vNW8YjtY3cTrywSQ9jHrveEM4QwtbRgkiohXM/RC2SootLUo
0P30U3Dyq7zqmHcF8dKBF2cqfI8nOTcmKPgCRdh3eE4aJOOj3fWU6x2zuYXInaJHCRTKX51RS5UT
+VVY0Fji1AenFIl+XPnyFHq33Rf5WXxTPxl6J1fcdQN3tRiM0jsE95bxnFMTZ964EzV/0xiHKigq
da555kF1fLX9N6Oc14qd5iMaw0PS0RPdjuVGcnNnQ0PeOExc30Ce8Tf6LxaJpeyOJtUoUCx5lrdI
xV9+H4eP+o0bD32l0tmYSDJ7ERrn0+Du5+LjuV9DwXEdxCn0N1/TiNMZo76Ovi4ifCrrzl82UnTS
wU/nMgtO0FFSWYfa12hp2GhLVaHTt5HLH94N3wbPi9HOI1N50w9V7TmD32NGK2w294IqaxvqkmZz
a/ssi1pV+2gp3LeMdP7SQmOcxZfXTe2ShMORPvjWJXUgjMdNK6SGkHwZstlQcZGDKyKUcB7gUcUm
XZrQYdwOcUcuNTk4N+DLrlW+r+Ef7h3KtPpmKOczwejefSit+PYKRlydTAHCyNTAjoCXvthocYpB
BcWqtEP2FhmdVYZ4E4MCiXWNdilAeMAEkTH/gZFUvRWj1a/bLK/PQ2gQAkELuesDFUpw5CAf8Ua9
c2btuAXIPzOzhdcuzB6LmopdEvRTob49M7aWGv3DlUfg9q1SKjsmLyRVkeH8vSvvK4V5frAwTj+Q
C/6v43wNkjkrN4SUsxH8D9rqjAT/akQm1h756YSj2UyZjHwZCeGYUhrJWrlJdHj/7ekM35t2u0Ph
20h902OBIu6vPA8pJyVk5vor4057/TvZl0Fd5SiIy3PZaJIE6HnfwHKFIpYXrNvkQ/HvD5rzTaD8
hvgpCAraTQEJ/FzNoqhUTH0LcClTLzEJ3p3/UO3f5zjzUQULVYr5zWU4zvxyHp558IVnOwn6ahYr
+oo9F2BR2fyIk2jFOkczJANTGBl8Ed/eALUDHfu71pTBJjf7xcNygrBi2yeJLDGVLbqAy6Pdnqzz
YlfDVCZcKEzpnZjWRb9GIJ0lUD3lCI25b73B/MWomTwRDh5pQxfp0+kTsX0TK37o+1kvOLXyibOc
UHBy0VU7G70w3/Lt2q2MihcqM7T+xGv0nzC5a5cWGDOgOaYCsFBghLidUYUUbOf8n3P5SzvWNjxL
5g0rKOom9FiVLb1paZe3644wR72V4oWnqBltYFYzsbdwFDVPzabmToplZo9QGyFJNM3ZGi3DHOZO
kwaFN16I2PobgAgmFvcG+5gpZeWJUYsQtA+urQQOdSteiG+ulAJ2GoGsdM6zQX0YVU9/cbQpgKLE
1YAMVLGj9TC0G9SVtO416W3d+xxHmZJIG6aJNv3sU80z2NSaHwnfHjmxj12Dl2xlTWGEK1EEbma7
YSlSpm6gqwsjD4UgNKgmE+mkvlAWT7VidDxv/G+NxfPWZR3GDBmLQFiYSbLedDHsoq9E92K5tmtS
nhuU+1uxQqYRkKMufNNicTrqr6gyQRK9ugfusPNpBtc4xnndnGzqs7Le52DJnkQHJuG1wp1xEuug
Avzp26KidmDBcdmBr2uqr4OXya4HCniXlKdxQ2qh8oyCpo2CskQWFWtW2YkYDqqtDS0TX5jrE5cf
5MBaQ9wRrllmrbQZBBh8zw17aUQrG79flAioCJzP4xm6Y1o01W0ZXfJTRwrPKaTF3I9JhE/HQGr+
jN/Rua7ievcDGIicIc6MwhIlwR8UXm9ExahPQ4ssenhqgJdzptoUToUMWUf/Mn/zhYpaHIBxoQAn
Wq/E4PLiQgSQwSwv8nmzCZ1wujVBO2C+Le+eaMXCnob4HkJaV9YD/6cSHPjf9Vpk87FQHnSSRCbJ
WXEr+aFUZ3BooRfmdH9jdPTUngsxZc5GLJuZQqEEYxakJm9MBQha3G4pTz61
`protect end_protected

