`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hNWJoYUKCMS3NKBPDEqpUN3/tM5SHTzbnFf0cXlS9O8wG5bapAVhnYo7WCbi5bZGepFHKmhoartg
GTGuMOCv0g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o/7RDO4wbWYzMH7PuJvAeLWF4d2YldLw4LiwgRv2KwngM+dtzgPoDX6Xlc7+tNZk7wN5pm9HVSJU
e1Z5WHJKuMWIWDThlSkp7Wyzj8nsoprneMVnZYb/RuPiMnC4wphkU5WYbqi0EXs8zElrQiz+n4AW
bAJcAfLBkGs9PdsanqQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mH5ZLcJWPKlcP63Kztre2q+RcW6YrCSHi7ZKOAxBNtcD9c/y+BEUrzt+9ECzaV8J0LEv5w1RLRrn
/ZCtyu0HnM63iFGpCpDLPxjPgQ29f959Ju9/ISOpc9fReaL9c8zNHrQxPwX1fw6dUq78YDc6M7XN
sMc7qNW6RQ/BOCAdaGlOieEXIwAO/2Sax6zccyCbfXiXC4Xm6dWIRazbF5OyPRd2o2c/Gk7xPiBM
SJnvVh5RFDBFthXnT6jR1LmTQhTIYA/ozDqjsI2ZNz0XLDKPMjvsYEXcBz2/fW+B1jn4ETTeBiaE
2cLUC8Blxwb2noQVT2naHav1YCnWxrQv5Jc3VQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k7qEpRV7lVsvRo45xpEsAw27hSHrKfLOebKwKQnVNusN1g88wfmd4eyitfZX8dVjb3vd4o49h/PF
RRmgH9roiY8MPeV+zsFuiy2PeQ795sIAgaDBljM4Gcewzl7MaBmLgd0c/5VATTmq1ufnObHs88kC
mb8f8+4Fd5tDCb6XCVc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V0mxbyBT0xDddcX5XrI6T41qozITpFwgpZ3WqxRYSaEDZum2cGWMlqvYBeYiOts0Xsneo3+ATPEm
c3litnzywSdTeVoSWAt1ppn217g/wkAlZUzIAEiNGf9zxOpX7Gzp66vr/wRdBmyFruFS6+Vifpo2
WfnferF+WCG9nEsn1R34C9H81goFYOq2gRUYrpwgr+GfBZL8rh2zFLS8c2l0isEfciKctmmIn0Zv
BJOtitBfQyusNZmr2oQGDD9lCXnv0OVTvVQW7oP6+4qQADzHgtuz6c+PyBeY0x+jjI3FqtL9vhyo
0Ez/J4gMreBvZ2WbKSFuRq7XYLc4QZWkI+mauA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1540512)
`protect data_block
riRx+I8DqrZY3BtxICLWXghyDqVHkqkWBcx71aitNTunG6HnWcxIRFMls1/jeq8q5SXqXxwBbRzY
JsRqJMEekNHi2xcA0kNP6SHa7LXV2DjtPDJYe4EBKQu/ke5mfQzzPNpfYU/Vtd9U+/wV+g4SRwpT
1ZI3Sat+UkLbrAjSASGdF9MmnPzreZty6rFVqbVVcKr1AQZVhtSAR5pO77d8/HgZasG1HoWF9flp
/0HuWVP8ynqr0Bv+PLdRCDBkOIETgkZ3MaM8npuEtMVjxH+Qc2VCXoheRN6m/+SovtysohYrYVSh
6RxjdDAx160u6/QzRnwbMqJjb7ojdeHVcZ83qWeSvsmuWrBLSip6OWxVqH5yfPaf3ehpSnZD1eNx
aduWIHxbBFELX3qassDMTb7NYzEwRvGn5/5faSBBOLuh3snszzYayq3AyN1MqQuqEohffcyB4Ysg
WxTBmP/f0yX339Hn4L7/yXAWA/EznYnF5P3T/F+ICKHPNU391I7hipECjR/1VpXQLyz5D7KLHBEh
VwgaFIVpwnwE//MHzj9v6jFpiK5BMTvTDmDjF1tbsOOlPyoJhMGTGY1184f1tR2BwX5BrjG4C2hS
55GjvevHVCTn15O79mXMnfjNYZLtESB1c/9Cn0Y8HUD+Ts0YASUDkPw5OwrpLiLALWo7P5NBOcEg
YxX/puNgZmVsbVaF2GK4/W5XABkQh9FglX3Rc/eolyCfvT626cV5FkryRlJPs/H3F8Hn+/WNvuIC
Jho/zOf57y+QJ8Ew10V09qWZkGwtBnwemB4ELpAFX4HyH+UvLJwEzQD40tZtNxh4B3K5TZ/RE4BQ
ZN2MbEl+iWSIFzavwLRi6X0IEdD9WXQslIUmLhmq4eZWL4Aro6Gusbsc/sA9IcdLrBb0nFj5RHHE
vUmG48vGN+oc+HpAVUpFsO7bs3eIPNwTGrr2X5WiINrWJX4WG1VTMkfxmExqWJ8sCyiiAg/C5zNe
B2dvF1Eja6cIGSyq22hw1rmHdVFxdxuWTyjUrRYa2DuD11c/l914Z4skF/C9oyOU+MlaQXpz4kVx
BCZAh3Oy4qy/Xc7XeLezoTyBPaDhfiTZ1JSiFJRlTdN88Cw8NYN55dTLyolt31QK0Trab0Yyk0Nb
H+Bnnf4taSW9MjRhEW9wkHPypjZl0/AM6WIdfCFPAOs58GnF4hwVsGZ75enQqsBukSetO8zAj3eQ
sRyWTx5RxYgsOdhfavxC222u5vutsm9dPgwk0KX5Uqo6xFpHsZDui43ziE0k/V6uBbOw2MF6U3SC
J2U2Xa6qooelF16wK7kG1e8xYYgWKrj1Ba7ETYqJXYfekzoVn0dVNtcxDdWogln9Mua05Qei01ND
s4toBQlfGw2SVNNde5ajiAdtsfX38jJkQuSQhmOJI9a19tl7a8qn1wanLZGYblAfPKeJWR/4Ue9l
yFU85v8GqCwGRh+suGN5s2dNRE3G2GdiSKOK1hzDrTttbzonMWYPv8PtxRS0+rPEhkvpWRbxk9wE
kCfKk+4zKkoODwHFqVfjIDmRirb4Z5MNrgVDTIAbJ/JR9kElnSdT1y38uwAzFQHmZa9A1XJggowZ
pCamvPi7r4/7y276Pd2xgV+mCS/fEk8cZLeBbFgnGbxA5vcOQfHdBVcPIFQf0WBZRGnaktWrSY1a
coqwf7G19O5aLSxiJ27teKHS5FNeSFBadKYfMELoXttLcdZRTsrN9QeKAF3WHfYZKzLZ10iHOv4B
Td+RS24AFVYAm9QeKlsGocE93gRopl+VIh1n0pzSozBKtaSTVMucRznxWDv9BKh3FVeY+aQ0PxrB
BEPESlIDvyAoXtMQV2/fD2eWgbVkv/XyhvZ4Xc8Ng/8sh74UHRQS6nQwhHqEu+IKEHBiIbRR34Tj
9+wymFOaJTRpleM4oO+KoV/4CCUavWbxSRvCv/CMxlPcVBsc0VzaUHQ3wxaWaOir9P/r/SihULOU
9pg+TPaBLqMejUSy4PsrPS9mlvv8XvVNAykaWaZwrB8M9iAsbuti3hK2ZfIM5hdnZOZgd0Huu2xj
haQZJ40rhWrUMVFymibUrqg824sVWx8dpLse8Ho6LUSZENNvI3nScWwygEu3XJTXbqZXeITIutfq
39CBN4usjB4BwOJfrCPIwp2WhdCBcbYeaASjHA6R00WdjGMnxxKdUGHxgnQDUZWRHYNhzuVN+4c1
rPePpNCh3xDDtOkNGYg8UEI49E884xYG8s3jW2ARVSs2sW4S7xJ7Jk2FbGu2uv/ak8g7j1Ww7Yf1
4Qi13KBZBHH58viAl9cIvIcjLSYSYjXysXyCLtEi0ZHmVcO9Zz7Q2MvAvyhk7zPKcxpvJsWfIJdL
+EgQ91HW6NpY9G7BpNDFSXVANxXA0YKBgH+zqk+LaX5kqk2WMvy/YrNAjhbc2G2iawpSuUN7kdrk
jv3+FF13LNHWBopE+ADX7wXnnPcK6hY3QjiCfrV54CoVAUTzuzhNbIIKNLOnnQaIuuCDMXzpOwB6
3hulfFtzokU33SHA+q3q/13bRr3EAEbC+oX5OWxahc/bBsETtx4T2tjlEX24bRXEJ7PV4T906CxP
SJcZzRI8hjea4pARekNQdadUZttAIJoo+/gRtvbh4iCyL4aqbND/yWGIc15GWHidoI6C2xhbelqD
sIGCLqrKD4frM2jMW9yhLeiRfzX8MMo5/UtxfFP6yO55b3XCcmn1hNrieYBtTy1v7JF46+RhLwhj
cVTG56bgHnCwX0SUpG2duu4hpB32UPHBw/mzE9D30ZdeZJyOxniFL9izr7ASmMGJ0huVMkk/b/Ee
lLS4MjQoXn6CKpqDsMbPwwAiBfe5kcy7jd/SyZVWuJm2XdPwRGW4ryJPO4i8XYPDzDO2DlHEqi/X
0nZqag0iAHYuzloVHzW/Q7RcIr4JlivDDUbgph6fScHkmI7Xuc67zGIEuV0MomzM07p48rpL8Q+o
WdUSm3STP3F33FKfZm0cEWR8dbHb0xn4+PJKG4mZQFboFXcDZyVM2LTVs0gvX6qV5EUemtcTCDQM
nzE6jAgP6LckA0TnzgWj78TO+7OJLCinPqhC+i+CIuwZGyxVL1+S/sQsjxn48pxXDmZqCRlDI0yr
uiXbJzo2IuYehXUgdtBUsSQQRzmvUqMhgF60BQTEBZ44XWvqmysdcI9G69iKYf8XnE/UQ3hzs25X
ogHrgNPpxKmGyFLBCpUT5BGFGBwEpeSaAElpUjKagOvFd4U3jswfslbW4P07f+gndMlcPsA3MKDx
CrOKjtcvbrLrF8Hypg3WtvHFjZ19lli4PKqr3g/R6bU8V37rAd2igt3QO7UKGTCd5+KBByrSv5DC
EWsdueGEe9eKK2zbQe5g2JHt1ksqke4kUo2FrKJxRmOqalT2hOZWP3DuV+O+x1+LVA2Xjop0ozve
MPxUFHjWRO9V7Xx+rPDPfta6Iz6xrCAQYDvOJ/nRZ6mSNnoPwaQnhw/WUR8E2yF988feUmV0QSXC
QfxjwDalopX3OOoTRE/vF+Bz0IIJmUH1J/aSWFnF0DkCqLc2VNHRcTEjK/fYET+RTjCl18t1KJk3
MM3n3802x1Hr0YbzFDgmJIZK51nNFqOUFHoK6ndcNtE0EbuxmNtyVzE2RaVfncxOT0HhjCFevEhd
BgR4+x4t2JTImQ5b7zR7Wjy3boD4y/THpmQkwTtlgV/1+iS4vujeAjsJOUXc9LwF3eysPuU1pYuV
jT4cuu/GxmGikMXZEN4CPHv9uET6Wv20QKED8d6xGyxqF5EJqis9SyKHVbH6YuQrDQjAwPhgkXSz
SXP1S7JHWQT0GF6Ea+E1Hwa7mb2Qr2jdRey3oFj5dMRYi5YipXTeKHM1LLWOieNEr0Zr4AWC9a8S
LAvsjWgq1nb73u4J2yeXpx/egDL6d19QWRDykt10aGtrkksRdyZ7T7W8Mm0/1aGt57Kvi5lMN9KG
DnRiBFJb1AEPU2ZZVPM5zhpSUK9DGy1t3CHodc3Le0+mjm8v/sUevB5iKoFfqX7YiSMlc0moSJuQ
cDuvtkcC2ATnCKL728poajVbsjRuk3vVEh4Wyk/jl6kF9adz9NMh1zlUIvEbw+EXQNBsxzobcSQY
62lDA7H+IwOaNV8EFwjJkrGNOXWrZIISl98Gg3yIkHKdaJIEiUxYPqr1NTgGHKZWEBTj58gqIqfl
TTjTUrxwjBmCRWy6OXDQ0YX42R8jFzwVJ/jSR7myPqJcEudRe3ZBpAVT6VFk4GbxYthkEKdPvU96
eJw/IkMX/bndnxWhdrxGDHbZN0np6i5v12JGr/CdWf8rQSb6mK2Y4cFwqYT0s4bAv1+8+AJNZHF7
2UU+9awo2Amv5A/du0LfBirlP8Hna2BnfHKOwv6uzvAa0UAWVCLP8LPwhKIaodNH0sTTVByMxRnj
vMjrNcjA23MNqKI/ztAPpMRYj5EP2k0/7J4iuJyHa0AgPzVBxwP1jpZtfrlXP84q0t5olTeNt5OX
poUuPQqPTCxZYz3LVCRP2OJNaYn2+H7niIH3V/f374lP4kHIbFc5cSTl1mHJQZF2+LnNK6a+xTSA
+cgp706L42SY7xC7MrwLkaQ9eA0QqHdakLRYl2OOqoP/B1jOCbWndo8C1gCY8AixrOrXJhW2NzBr
sIuY1hKcq8Q0Th8JLiQnoyGDooprEjuNI1BiuhAaJt7HCj2Yr2xggZ4tuNYtYcI5POnLGh2wnruw
5PP2ZKE0+ULyK6hdPpMVdofga/RTTwmpdOkHnJGX2oewLmzDIkSc4ssLa3h/3e3R4i13Qmg6MuOp
k0YPjKQk0j6OIYJB4CCKTDYgPSOnDEME5xROvxQfpuZC3RcPA7oW96JntkfddSFqCCT4UyhugCE2
UpAD/3Mst3VjA+tyn12ikLfbZLHY2GFSj7ISNdARKF/g3Hr7m8RfVBQsa+Xzs6vEMFnWkS8lYx7y
kJnh3zWicYRSVIq5VY8eOBkSyO4zK8lEumHjOAIC5gKcqUdcoijCy8Pkeh7jvA0qTiGpz1xNmTJi
uHBhmp1HV5Rlfn/+6azTWQ0oWPG2IGsDpJqXYEaY8PvIKPgQAkv7M19Z4SmYlrF5miC3PFwLp0ff
ps+d3vw8+xyoEuylokeRzI2Utt5J68XTOhgUhK/rJZPTkgfgniRwCBx1VPMEDVOnwPRU+62HmMmi
xYKfFDSmLxJ/vfrsAAj2HNfkacZJOomGhAFwckwxvZd/rtL/dofLqke6g4RnUCXMdGlbYWfcbYPe
eiJj7dPPHe7XilOAWYKfmBwo4arPSVs9FOoJQRJi0UwlmMeFvRML6XmwfvrIWV6/tEeiT7tQLwVn
70ezRnJs4nyYwpQystHbg3RezDR5Q0FoKNKpbyARHfKYFCp0LFMBB/JP0/zdU1quw+MojHtA7GUb
w8KWJP3IypDTg2y7GeIhjyc5oVN8/2tHaKOZnRndpWJ4fxVB8uy4gBhwUp6ErtEx3qHcm3Zo9hjG
sW0zmaZWbBMl6jKFM3SY1dcQ4hm+bLvhi7WW1bfFTFQCAFzIG9Tn73Eq5VK38hIl9DbYvADfTA55
gDBB8IW3KNWAvR2LGuWZwF6tBrOJmHDbN9NJZyxeY+hylsULlWE6i98UTL3x5+bYgG9wWkWX8WKP
mc74GhYcsnCWbjkzEvtVGdYK9bPcAtRrjk8eLZaIzmrdmq0VbcUGrnmRU5rNMt0ut/s3AqHwXaYp
YPk2/JbUu2nfq0r9G+FmJjOZNonCmQz/GtJDjBZ1ajwzeakZ08w0wfsSGgGrAV5SrPGs+dJn/PhH
NNaUxw5EN+n3Dd6DzGugRKJzfBsdCfOAGkbOBrp7qlKVedljp+uaDtVLF6FXsTgot12Yf7sHiQbd
G5atuYNbBowy54DlqkKRp62+k5aF4qS3R3hrk2qW9FFp8lH8l/F4ybNcCMEe2xomFrPHA/Z+xls7
E1mP5IrOP3+RVgqmNNS0Oaa39t1va5XmvNDKAQTOniLRA8BJVImxOT3KzRSvoxFqoVYNVAYSw9IK
HSvSnoN1AH6TPRh4uZVLqAHz86a9Fu5hrwRAvd3MLWnzL601Cg7drgqQBd4QA8/0DVAlaLDqdvRM
Ro0b9nhQqBx+y8fOnhgjyAmCmocIBiQ/DX8jXEm+hU1yCubGDvmu47HvHthiTnnRielVXXjY9wTG
z4IHct9iebx0Nf/+cyIClCHdX5d/ei5iJwoW+reQH0HI/4vdfDV86rLlvARFS69NQn+yHYXvIuBP
2YUD95RKbrNZffpDk0lyWOSG2PiVy3PVacoRpPbHg8s4dYIUzV+eb5MMfkwpXlYafLaLiebhk9zl
LPqeet5efxyR3HKJyQuKjGlKqo5TqJJYm7Z2Pi6MMs3vliRua/VyZpf+2HRjBYQZwh48L6uG5Xkw
eBU6aaxkjBHbByhEFVL1MO32+hSSgw+nzlY+DBTFXuSU926Pyfj3QuDiAsP321YSpDI9G5FXCZb4
GDiCBi60p52oMOTBgvKW17JrsBcUOgytUjlyjPPGQY9LRjINRxAHbXjgAarjuTH8uvRKSZ+oJ9NC
/tTygihMFNmFiWyPYUNYiTDslcJsWYquznQzFPAYerivvgy0U3XjwDfG6QnGuTRjpzv/Y3nUuCsC
ElZwubN8tvTRUguJDiKM2Aouoo2FnJF87RPqKWE3yyYYE/S75KQY4eOxNYhl0xRehkqd5q/eECM0
oxQ6GfdhCgL7Qhy0JjcBvbly45/ZqmldPFTeFuIB7Y9FfTltHHg1He3dc4kdtJaONgzuREtmUGYI
XgukCL7M3DbcvFx6Tqx/6tZVQUb0F1jq07q8nYjxiLdonuuRjI7iKYZprLgtA9NIvgfbzs1Rtm5T
r+NP1eqCz2NhD4OFOlMSV8L9cDbyT4amG+gqDALdH/VO61F+jzsyhHQoyT++nRmlrOnv+O4ceHPu
3tR8xyE7vI/7ZuvyQeV5/x8atRIwJy3Hk7RT5Tt+6mfAZZ+ZVyoqxwGUR8InD9iCHMpnrwOrrk6G
E1sAAzbj94JQw0HrxTo0d5fd4W7zoY2gvZJyjkQXACJqBfqMRtg1Gi+yTkIHPzYiIjOaGehigkYf
dkBn7zQrqdp15SRFi2+XKKcHS9yZC5VjpSXMZ9+e7CH1isWyf6n2MRapQ/lxtUmWnVGUzl+w7QKJ
am9uK3Z14l/+FlhxbcwUQjxtien0Qb+QJRV4w2fFm1a1ZX5yJ3swgkkoxtTNy9WMV6Y2JaeeIavU
7bM5P09SEyc+bCygeCYeyM2R947/dKdI3nVr8UcRCQX7ExEwm4TBYZcBtcwK1hYGpXyIiZMnt1Br
l2jc20Tp1oDNlzAqjIFfIDSI9St1E0w7uXCv2aqISUUsOtYTg7d8PS1t088u40INAWsIEokJOhIp
QTtOGMdJIixmbwwEO13MEOy7rQO2T9LJZurRLL1EgPNByxkuLIoUn2p4kMyjUdPCg1Ui+hp+c5Z4
q6+kPj7nD0qpFwpsCW5qZ1uacs0FWtwlCBlwJkvlDv6JqQQUYcF/2y9Qj7SbJjvWKkx2R0w48kJh
C1pqLYlryc983GkORrZxqPh/aP6HB/o2h5b5eQ5r6cdeEgVkLsPeQT5F3KwgdwAnNZxwHNUqIc3F
zrHSwaxD4WrouiMgLzn9kBLgtjj77A4xSn/iDKRp9Yc8uuR7In7PDtfqjzDqiqukdm69WaN0n1t3
rbCuJar59TJJqTakeo+yuzej91xcxp5h2cVCtmfxpYvlcV0PDhONDiw/HjDmCga24arkRh8LsLXP
/Naypusy8bBBgNPy+3v7xFyTi7QzLsfeEkDi0yqF5oKpw2Moy9Xr9nWKjzXlcwf70UBAdulOC/ZO
emsziihlLcGQUkKoDpyFqzz5LOkrtYOVLQCAgta8RCTFP1R2KV1l4sa1BJDDD9Dg+swiM9B4yBHD
sBSm0fjJrnoDpXKcAcqllQqWJQMUS0/Z197aLRvduc52AfqmsHENo/EJlt2dcdpO2jKXbS3hro/8
qd5lukO7DsH62C+I/BXQLzmMCEsJ61x5NnSUN4Xds1oGq2ir+oSCxUI+W8afBS55f0siC9ew5lUj
xKdv8J5cmkNXRDbynLvyQu9WeD9gAwWxuLBLeTETtpmcrQ2Fj0MmIST/7sBxLwgIAHzsuXQCHCfJ
H2OMbAuH7WoAUW/JnUJPhYrCoV0mjWcG8ODmzYEXK3wTijvs+5qACg7qQBY+n1Hghjg2eUufpvL9
7UBxOziskwiyAQAmMyPULaKc8oSKX5K3+gh+5iUOIy3ugk9GbjCLJSfVpoy9X9RRnbqcqKacV2bx
gquPShTg7r3PH0PZNqkbiIKyoQiNapLsk2ql/rDPzuesc3yoRwlmpSKfW+1Q57Hc+a2h0OgPGU+m
T1Y8HI77mSWsyFMNSXOsLHKvKbfVcCv0+A9ePq0dDk9eNzbhqHST6CNthB1S3C2xcwqp0H/VmBqD
82dDkasKN4gy+7Zex9BC3bg13GgNU38+MBzskVIKgFsVrdViuM3cVChwa1qi765qTNsWvs/syIG/
ZNgOzwzOrXXEu/WsBgg98negBR5gp2KWyNH/TBQc/jep0PR1yF7ZIKo8tzvNitDRgCaS9YksRGuZ
eY9LzuzV8Z4ig+a/ivYOBFvUUrH9rHeaS1JaSxPKF51IyzgvgnmUeWwDQojI3jdv4XnsYBVClGkZ
rfGJYW3s+qvn3Fnfp/l2+No9bUFmGd5LF1liO0SQ0DutANuK9y3WmGi/cD1tFAnxwGzQC9o08Uc4
ax0qYlTBlmRfplaJ0DXoKxGVjYfNZNc8B0il6N8KFF+BLh8ynseqShGNB4cvddyXqgFU+GDWwO0m
WuBdbJzHVpMLO6jzWAxEcU8qQfgcV/EFe/9SxVeFKAZ6DvoKwaB0j7b4xZcp+aEuYuyfe8xDdQHx
r/Wy6PeWZ0eJIi1NWiDsz5teWvDhSIlipMERY+/zIW24bTIoRlYQuM6HpTTztBgOlep1F3M3TF2R
V+3P0IrYPWOdezWcNpStoMqyxpOG09YuMa4EewcjuEq4MEaA6LEi2/Ig9gpDG/FId9/PhCajFJug
Uty3WdckBKMD46alVL3+Uo20F1ASEgmZgn4K+r5+GrwzvWH6hn6a25kJIi+tLdtWzoMFiC4jbdIW
t7hgd7edks5Lz19xaJAoQ6uELy2kJ7jjsrsSJKulWA22msRJzcnQsmU/aMiujQaBEg3JvZ5nF+GN
AFRz42FzEDwomhpmAtcEn9Cycd3NcGgw2rWRoSz3Pfno6E8B+br9c6/bJhSh/IyejThy4YLsQeNh
BVNyIvSTzn2MpS50GuD5yBiUFlu+rtgUQGclSGGWLlMIMJTO+hD9igVGsTkU28uuKsMaxr+T6rza
Etc8A7ko451tIJY2NPof1ExhPqpOBIXr9+J0oREos2g0QVbM3R08KXPEUjpgwsi32eT0Ze9CZVgC
arbzlQQnQ9gRXOBuxpL+zmoTkVeQ2999ik0zHgH6OR2zEoAX0R3Sub8AkWKrUkyfW6xgzcWGoFCQ
/h+v3zjRr95amLwLw3UKYRVTgNmsKqMRThu/tfZ5g33VsexSYRerFFPtYUjCwTIreZSykE1l3t/H
AIJYArEKl14ufEaT4U5Kh/d7JAxIOQC3r35VGNcYw+PR9grvceN7qXYgOGa7iRhELJPuEWfGYw/q
d+7nWsxqpQsnl1qni5mmJWx3VrIDXtd2UX+aOLx//4zMUsmEJCFDoaPZDVOR3WJo3FxG5SIJLu9J
a9scJ3jHHPm6wdvPj/AW+gvks0oSvj6Fi3DWOQpP6YqIKORu05ZdITSYLGih7+8Dnqsyzj6DU/DB
i6BscMkQFm2Y2pM+LEnicdNlcTuYJjw8Dogvns1psVoXffbcY8Miy0fTn2WyIuAVFqCmOBWCH58u
hBccHLZtSxYhmqeqM+/ZC68atzvurbKlMf2WwojUby8VmRuVwT2Ev2/kBv/CRZQVyAI1G7j7I/zM
jLuGOk+GMYeoP0Ihc/xvc39dkb0t3YvttBaPEPCclkGMlLLiCyV3hM9CkmnmokZ0iNLJp4c4nNmd
6n2cUccMTq/TkpcP28D89OBs5WRJU6BWbkSwsmJi3soSkwpef6XFHMvGMTzkzEvqPqCzlWooMlGS
4yVLGfGwRQiEidpgIYMlxxbr1P1p9+KzUSlh+qsWhotRyIj0vzEZHxXtesC0OwvAsFQke7yuehIv
ORcp9XWP07Mfav1qui0CKJ5I/k11ixmcGcH1Ish+OSkMundLcXBVCiTi1XwvnuH0Ko3E8oqTSFsy
UFQlDDt5HB643K+bmjJj+piCuiuOODm9kMPiow3VsoaxuJh41/Vl2VJkaAwhcMgjf72xVvUoThYJ
gaKSvtdnDuw0Rha01QM9+07CV139V1cAVvZdIM+qfNyfGSbNJbVf+OIbPKx6g5UZ8L1Cv1kTqj4w
FKjkWCopv5RdLu7OMCwM8vvlxegiaiN9glNnCtooDok424KAwB+H3vnScOsfODFgWuLU7hd7h0zs
6efLgArkRSIy0emMhPBkHUiKXsTbdAj9jLlv7BOwOR89xtpEsAYjQtOuacvL2P7fX2khya0nAMkl
JLYnPTVTcB2V3u/5JVe9Qhj+wkaprnI/+e8cFAA+67AeZvRw2b5Mqap0fXgNNu/GuZHnoJjmYJ9t
v0zgpNTmQ04JA3tTV21Fd1z9lIXeq9X27TVKqmggkutUcD48ccv3YS5xAWGlO9ICuy+EGV+ug6c6
1IeKJ+EMems2XpzrvAUGJgHL6YwbkTYLRUsRfyPHqkxNTxjq1azxDSpj8MbbMtQ+YLC3RRCsuHvQ
8dZG4tYWVpsEAF7IUs34fF/t3S9YazdAfSrosfoqqHExQzZhkaBq/xLmxBoWLpFYY1pxh9M7A9hq
BWzpinJsLfV9OQlHhmOvi3Q3EmvT33lJOIleaVBmuu5KOfcGUGasTVoF/WXH0faBKjaaR/Sr2v64
u0TAuarNe6HW4DShnKWSv5Sb7audpvF0J59XUnBJ5u5trLhpQipv/VRP0QKH0PgtNLGzj0NU0kGJ
Kt6BROdMJMia8rkcmAhhb4z09CpcBXvjmBG+oXPFkVjvVwl2qj2LdG0CMqgr80xPEHaYRRN7cZDm
fxxD5HKQVODoIIDMtwPRx1qaJIXgwl4kmxDGss0KkBRO1SJ4030NColyCJ7lnk6qe2YHozuzt+DI
yjZKXvvcJJV4EIPTlUDgplAcTpuTfaUsjQd9Ht80KvE9L7C5oQ/B2QafAHyUbwONeOcN4SslYkBW
RBxmkCoaAYUSy8+TgONQNuGqLPn90uj/jWYaNNKrtT52I3Ccagv0Hbds5R9hLfQRoa/iyc5YwLX0
5+dZmBtBJRXte3yvOg0KD6a0/gPZM1DifP+2kZwqsSqFO+7Rd6XDpqNbgDitrcXcGbEVGZFl4C3r
uTPC+b30Q1kvkg9+P77EC1GgaqydCOmDUKittqSA5QxJNesmVjsr9CqvifU/pAdzkUY1mouqUwAu
MdkrHB94BlGvZYAShxk8Ceu4AjUsSuf89tHMaGlBtg+ema2pU5jY+rHV8AuLWynQxa/YRqq7zL9a
odzxN4kEbAzFyXfo1gexWVug0X5RCMyhl/5p7+f3XPJqYnDGIp9RSXXaoRmtueCntz/n+qnqldWP
OISdrvTRPHbxI3eMRzZSM1CkKgBSvhTXRV5HVBn1GcRw7LtjuTdZkjBAV4RPVaFF46sT8LooTjfZ
/6Mib8uYtoXMT5tqg4gmxxRA34qx+2cNgiOwTX4voi17VRMF0cc0stoT8iLLLYgYUfIdDxyJxzHu
alAFbd8Dqph57fwxQF9D2fa+zH2J9MYbKAEY2aVkB28LJ/2h0Ex323fmY4aNjBTFUMKSNXtd1/MK
E5vP3SLjMkjdUESde7yxZeKFuOfg/nuwfvU7I2TczX5X4aBpQ06sEkYtd0EKFtfNWhPyZVLzdItb
4DfH6Bm9EOXPc+hSTM0/YHjbynqcSFYBB3tMU1Xi2XOB9WRlGfMrN1itpsLI3QmV2edZwEKt1jNy
jbsOzTFqSQhuSjJpvumhEE69PIcfqOK6qFWPkj7SRBQIk1beDJBdL/rwgjzThGZs9Lw/5oh6YbGe
uLeOCxIHD74JoOEV7cbnQi/+er8thIRcLqbsTs8M9tlga7huLsEpMC+ivo/rnl32jzqiUwSLUkeg
hVv6CiC6OT+a7nSKp5PrY5ZC6Ipz1NA/JTF2uTManjIK+u+58BVM03Qm3OYv7ExK9Yp0L13GbOnh
M3/duTiWIU0zxx/Z/AboAS7v/HK4agJfX4jqC5LG3OJ6Y+UBprDW++r6Kptai8ajk8ucFvuJd8cA
K2Eh3UbG0N6c2rGpvbMMpzdYYDiO9e/mPuRkt9RBd8EE2KWlSb7iysABmmZA2jPWNmoQWcvrAseH
AHSVUweF2XrlHcKzQJiTlZrmnI7XYvpN5uAogZkDaCb+JXeMwbTe8q4e1W5iCOQjTEARQIrBcDaI
4TZeEuyMraNPHDqLCv0zNbsc9pewDJsK/9nJHu1XwGZTyNGYzR81FynXofihyC2xtYc1R7B5jKzo
RZwFHVwuZ671PxVwl113m8Y8qMAA8gjjgEEBAYCPWA+V9ZrMbc+uqSB4DyB8dQqO6YmeWpSitfgy
d7OIvoZsjtsr+wK19oYu40FUiTngn3ZnLAzPoYKWiic25fGpM8XedgeG8KYjPmLm4xy0lE81N6Je
cpyIUI0uyjktxNilOPYifH5budYA9AZOFcWVMhJAqCCc/Qp7spdh2ulW+THasBSSuegvGsVOU6EX
mCPtP88fGJlJhFRlRy3D5dIfrwdN79jn7DOs1nj6cInhhIWIe2FIikh7iyDP5/foW1kgLmnlKTPN
jb8FhrLWIBZhw/7OJLzs83/23AV7x6pjXIyZeKNnjpvj5duz2Y/dc/h3UQoXisCKC2Y4Ie+OpLYA
rZofrW+1EGy/noSjmp7MPm2JzBB1CyPXAbqw037En6TWJu4EO+Gz+Acg4xekfdlzyxBOka22H/Hw
XR90FCULY1RKHs0hXQcQtsO1/qo1rdECXvWdS1oyd9xh6P/7pEoVZlf/D5AncucCDbNiMEVgYkiC
Q9c/JUBdZjIOdWp+ekUwyfpsCmFL0VfGswIwMTwJWpUEn3mSlYp7qr8yylNkUdFGJEZOkYNyUXLf
QCdupg9GeHxoZqRQOjoJgwxVxLjfKrxxKtOaBDXTqXrKE0Ip8HV8K+oON0cmmil2rdeqDvtqk/mt
UcTzON2X0JkPMY+PuSCgcdkAo9QQ22S6z9A3s9tXcQMKgH4Q1APnHWnvf6ykSrQJ0/cezIGOia9I
H0GODzb8osHLU/LgVe3Lyo3+ftBPkesdb3bRRqQOUrohaOi3qPhc+8gz4W7k1/5wwPmEZAkm5TzN
xbeUm9MNjXL2j3ThgysWYRzXWhxDBmYREGc1QqE03jfnDZ0TNeH6Cg5bIayJIjpiCgDwKWzvlbWB
CMfiVcy5kx8IQvQGtPECDJRjjzsvcLaStYaBXDrAuBUREQbhwa0uxs2cK2Zt228WIs1uzn7qeBWF
vH767fF48NynjSFgHK9M/HiDcH22r9ihvCBKl/0rhJn6AWZKLnYqNMQsWQ1t7TIrk4fhB8BG5Iva
vrdjFP7jUqMn+7CknioeHfWdjTOOzP7jf1h/SPVabjbNz8j0AwwkTwhR5TuqAkrqKOBBwI8Vo1aY
cIe7I2xfB6GESgP40jcKoHKUHLn07Hkv9MKPaOM3cdTJnbeyArn9H7+vP+dk/VtNj0XOeHAr6tw7
Udm/WaL1c8pGBAYM7b9syZ5PuQjm8fLmix6sSyQmf+Sw5bVSrYuGhdsMXLRKiJ42Og5m3FjFNqhP
DSTgv4OV0S+NJlBRH/2zEITUM1YfWyelESRV6JOfvjN3db2KvNd9KmtSojUM1zqCV/KiKZ8DhAOf
MF3LiQ8dfhKnV+ITR/DnJhr91mQrJsn+L83bifyxsHwgmb3MXplBobt1LJmcpxzRoUkIadYLGRUw
91EmX9HbHfvLKgZz88IyqNaNsBjlSC4sNvqPsijl5Y1oB/B7G0t46ObB4j2BKH8HViEOB3F2XnQz
T3B081O937q1hvJLlesTw0K93w5WTsDdGYjpJJyTxXVQO6IojkINc5XlGWz1avaXX4kz8rm/HDZi
S155RetObf1AcI6NkQSjinbMiieT3QTARoFzW0AwhTlo+tBGVVcH/hiEcEKYsLz3mGg7hdFNH2rt
qNFc/E2e8krPdVORdrnMKghIGsgoxoux+pMDC0MjyjisvhTANCd6lGMDs1sQreWeoXzczxHSdh/Z
yHGlWptjlTrSXbsRZleZpc9Mkyk2vEZn2CwaUZENwy8LgkP3f2zwdDq//+9wHPwNonQZg9DlzCUp
OHmXLdrsIauq+Mjl7Dk5Q/WR0ies1b67K5lkw36tiXwO6KpUhDTHXinEg/Aonep1WaaDLsR3oHFU
bln67mjNq8u5KvNp9N+DEZSE0Oa3gEj2rfdqF6cn/TAK1wasY1WyJO1YdHDSJ49ANpdWqNSbGlnt
aisbQ8eF7ybvCD0VzRNdI/yF5TlJUq6GKNFzzf39YYSP1vEdLgtJU3jxgsJ17XxNendRriSohbrN
bGDKG/nibtrPnxbfzZDkLBIaO5L4HhYlZNZsgQZNY0qjKCJl7sl7cfKEfkltjRi9lKs79x9gohWs
xt4cEDxOda1EbtsS+PnNbvBfiCaZC8GwPeXma0sR+ueXw1Cr9cxswuISAPkGuDz3ylpbrKJME0Dy
zYClkZzv9T30ehPoE+F22F4BBgvy5J4P+2c4wC6JTs9AXEzNCk68+XbxG2/6bbSI+sfHzdDYrJSb
XK5snoym4xkTVGuYhUY8WvtLd+n+wCLwgqLLYmTSsM0ekcKL34hgcFv63BpdKeb4heRnn4AISWXT
VWmaYP5tLd075fQzU3TbASPV41kCq3TEX8o9mihmn+gvnfqBa9N2K+1hK8Wk7moeoI/O9ua79H7p
58rZgknY0oSWvWJsnwO3JC63HNA4cfIvTlv2mcAJCeG/Gpl/An5UB9N7g3dBQz0NTZf5p+NaErmO
+M9qbfiP3a8mBxZ104POdWN+Ptuu+ND/F1WUNHweDhrWlG+BCY5y4G1IBV9/ywfxaQ/JgtSuuL8i
H2o4qwtqG/wG9kDB9KAU+v6q6L83WlKeICLUR3gSn9sWNNHWbCiqhFneMN7FnjvOzUk3PQYrviUD
PYB67y5Lt8DIXRaoZI4PpmbV4JBrh96TsK7zAAI8g1SEbWPFMEJW5wv71pPMQJVrfQ22eYOTLhbE
47XAW0NjIbEX28IeTRQJRM6Un4vxbiNOPquf9jTnJRbUk7d7m7pjtR7/lEhmtTfaaSJNqttsEwtX
+h5chNzTuQhQkxqrD0NdKgdlYGwXHrbnAuxruqvGTIwY7IUDSDS+kM4HGHGd+kmBHBEBGJ83oweR
QUuZ3aJaxL8p4ULjjMejiVWQserkRw0+g0QUwvylNDrSWgeBa0TbSv4vj9a/HPPMBepgFdMPMSOE
nlXNhBsrDvj/8bjSoOyT7S/QT/zHljc3HHVlUupDKB13pDod4SZyzZ0LzB2G0+/iTWsKPE2bRTss
m31DlZg4aTKGRQtis2wfocciIqAz+bhph1aB4hQOT7DTyP7pod9uqVuICvmomYhNMPLfB87jxz/S
QmczbhlYGi7UVn6mXGc/PIc6V/JWBQOlPy11VJUSS+/zPRiom3fvQ626cW8ZU0K1BKm9NUEvDagi
z4wmIF59QgVTd6wrtw70BwPhi4rzwcTO6V6PZJ1YIEcd7pDl7sPVHOnQ0mZb9cx20RfcnCkaVsbL
utoc0DJq3WH45grRQzZLbq61rerEDrexAn/ekSsWvetfZxVyTO3MvEfAw+E+rRdC81yKeXH/kFBd
eVUxgTpnZeWn8XMeG6l+QcxrI7etqvHSlVe6dSGB/7kKMEjHHTwk6SkWjuCpQ3dfkl2+BpX/IjDW
mgRPSTaARud71KWJifMxvZ8F/BCsylHnCqAjICCjUdmDCWK6b0UYZJevqToizl7+yD4i2R+YhtPX
Kam6Nw+Xcm2TOqirgLiKJ/5cHCygVEWK6qqAzf2mCTB0xgucKJpTphi5bZqvZYzlrcy492pG2SFo
CPTID7thOYHnMg1rCENipYe/2D1X5K/KjejQWF3sOMxxOH3yX11Ji2YY0a7PalZb4mPQan9Xv+RL
Q7rRsP6j4gCTshJ54yKIXg8mI/8WOdh8PjvzJnn2et0BmerRMAo5G2vVqttjjn0A+FRP9G7+RDg0
xEwUPmtafkMiciJNtFxEKL3stPJuFfQ75b1hLH1+r5thDZJK+Inzd+qR0WiAOjzE5r20vmhYyLWj
YSb43N+/zc4tb/yOS1A5O3Zqh4bn1WhPqlueRzMyxv6DOhPp57SOCYNyo8G+25AjPGg89Vybwb75
lje7k6V9/z99YeOuqlNnGNpsg5uymm0aEMbhysaunR8mUlot0tyfmz1oTRNJPMCCJW3yyOMebuHN
ua22P9mRvZ3LFvT9H8yfSXii3H69Wp5JSxVyFa1fiBmefarh6Z6yX9d54RqVJdKERkvCrCICSYhH
kWQ5IvdgxMsgw3N2w4EC2XDDsVNiwhiH+UpXa7ZtcusW8RMh+o1ATItpmY0Fd55LU3Yr4wqHbpdP
hQmNamBflUVUBGWsj7rg6VtbOo3faFoFPQ0regcN9c01YQfQKqcEEK5g8TmxuD94QTvrPUNtbsG9
U+E2W4hFYVE+BvfwM7wGe9w7v1bkj0y6zqX9L3TRpN4bcr4Xj9OpxeTYjKyOWxOs5kJGC31NN00E
XdEruijrD256zcffoyYcn8FvZzunrVP5N1mx9wOuwxbr0hMMaHOpY6g6gcl/3PdW7zgC0HR9nYVo
JxEzMw9izjnat6nyIPpt1Gl20YtU7OoU79cNC/fl6IdtlcYHqUgNTjVetxVO5PSU7YNuBtduJ6A0
A7kI/YSzWgCITQMIBFMhy9nornhwhQEfaVCivRserEc+iYSeBiTPtsQnko6LZi6/01BGEedraGsW
N4j8E11gpqeRtCTouGLmv/F9eOii04SLT066L8q/GJ7kgv6GjpjezCAlKBpni/cB1KR4xynophWk
4zOhj1uTjFnD4kiChI3bDMTIG0MCi2mKXEP7q0gFohwFAG2acM+hjG/OBUS7B38M1KL4YuwChCTC
r0OKQTFSArcFf2aIBVaqJdsg7vtUj3D68rnCyp7em8GoC2i2S247YV/dwiPqvlqGK68eruirZZQ/
OwLKK4Pj0ymL67FFH0NNIBtxX4KIkyRgFgKAqN+J80lNJvh3N6NejdY0T6DlEH5VMYyCXVlqr4HI
MU4ZhXqhTVdyvbMprnVGPD19RNTYYjPOenxtC3Iva/k2h1ZMFNgpV3XxCN4fm6Cr0b6WstECtswX
eTPPQXMXL5GyXSLAKeTX6BVZQTDVimQIleoM+UP/3QpkkUuCGTCX8n8ZVtov8JOAQCQTRiUXQct2
yLD7RblKSdi7OMT2JuJqE90hBohdl42dbf9LrLz0YeMmPXf4MQXgtFJMZcNZd6miOAIK201EIsza
szQyPRNdSzG3w3WcfeQe5f7RyWjAEVEsw9ZNa588x39SviziaBXhsgT5PCemwfhl1QqhBATZj8D9
PRjyIg6tSc1BuL3WAWzBhhGZdmb338d27n7icFNTEViocuUJufHOFm6nO7HtTSAtWzvLV3pnKV4a
68trOpvPav5juSfBRn/Y8BR2BnkivqItLMzSDUzYyJPB3coL6aV7+JN+Vfm41Vqoxpels/VlwgLx
xom7FtTBJQDbrQrefomqwGSCAgN94F/WH9JgzYBQ1+H2XCAfmv7mL8CW3urY7fgtMPZNPQzvoiIp
2vfts4i/Ab8T5tLIntlDLqkWKyviy4kie9ZwdihxtDv1hO073ppzvB+rrxUE1XiEsnJlJLpWjWsK
gswPAnOUCHUjyhwx0n+sC2/ai1/wlMkP3j0srYB6PQsVDZgzTdNFZkcGmHNwGQBNqZm2v0Utcx16
ndQwrWtuHrkv1DOP7RNrb9V5sHstdZbDeLCWOyc9R7Gh//IapnuJpgLg+nbXurWWN1NYNpSRedyh
A3iiVgzBgcwJh9nZuAHyjjEXPYRo3XxZoVMhLx0jE0kImtIViwmTUIu44L/qj9Z/LyAwi4qBQKhX
940BKvxOqeFdtV6a4SOzttI7UJvO1d06NGnFn2Y9cxPOPaTt/cVED6EmmVdkzcW9w0S49GC2qzOb
Yy8nR0j3gq9bupbxv/Jw1kXFBGjVb7ylltJ5jrt+7cFslnsLZDfcOd5qxEde0QKk49fAOU19VVD5
hHYMWJZoU0AQuU6P/oMsxyJTrnrlZazDZYB1QllEJUgQGOy9phlczen4Vuq1qoay22/ByjPAVwbb
cfMJ3z2spyHQ/+JSz6XnyeK2pSIKnVYG07+jSLarDxAjF6mklBk1Dfi/fo+z9GRsDjHf9HbBCkiS
8niy+wda4AuJGSVPSk/zlGZN0BvNTWWdlqFKoq1aftTAXd0AAMATzPh011tLUr44ZouFAnwVHWSY
HuYtWEDLI5yjO5mKhypKlVa3jWcXCHxyuau/SvFXbchSbBRO2KfQK7SsPaY/doJMu1Cfi+Zs191Y
KfBZrKUeDMiytXheqGU/o4gHq4VF9lcxEmskaLtATRsUQRkTTXz2+Kuu9kum28qSfU0v+zkDmbfs
QQ7Fv9pGsJ7QmKUitoewvUWrhweddB0zjJOvKeVhE7M2Z5jXH9V4CirTvnP/2sHWv5tJsPyLNY50
3kCTJ1Gew6mpr2b6d7LEtH6Mqab+yIdVACHvsGSXBOvW5Nj6U2zwOY6E/Kv0fwhkYnjF6tEjMiVJ
/0yPO6U0dUsNpNy93JIndOnJZTjKy26CHbG38LvH81D9W3OB1dTqp7MLyaGKddVd9s+pJnCzmbnu
P4p/QG2T0WreKJK5hpO+VhqUPdWX0aH1/e+ZuZ2lJHlqPUrw+E55bxr0cG0at+Ze9R6qmDcBxhpt
djVJbtD44rn+ul7w10HfDxNCqizn8EpbVykC7Sx2qnUBL8wSNIXvMxFV7kEaIzVHx08GnnAoaaQP
GMp8ySljW4GTsoRPB1wQmHr4lU4tVnaezWCRo+Jg24wnMtslaIQizZaNz/zTZKiP7gYFglKpeY1C
wps+BCWLocYXfq0cASbPR0U12Ff9aJG3vh8S7qMOfIZngR9olcn81o1MmzdmuxN3wsKEbM1uII9M
P4bo0tLyjcbNrJMFICfVFM3aAWTiSzL7SYCF9fzRG8iJQEsQuYtnMKoTg3MvpVaUZw8CV8HQ7fof
XPBnMyETXNwFBjxvazGVfIhjOFE1BbvRGIqzDXMwR1lgYw8vO0YAqt213l/fYqIJnd31Z9es3aTv
uQ3/ktzGc5FQDR3eYwFdidbbRXB/q2fZB4W7bfw9whql4T9ASIM4nspedvZ6cXRiLQ7A+iT1gIVs
1b0fU6/w9jfEYkxWugVYuUioFDCBBCtN6ASphVTTXe0hoDPRNu0Bec7clYcGrGQY2uDkXfhuQIbR
ee7hITYGC1DVavBgmH4E4L+P6kp42wZ5aN7y/R5VOjY9IqSjU3jhhzkW/SLi4a0bVoXvAe2A2yJC
IRQURe8TLgycj3qgvnpstkCqQptr2VxVE/hhttlC3ay3abu4ek62GuxV0gOA3Db5+aEwaPnBv4Yo
TUSOyEdV4V8ZNlmwsxZUkQSfNcxUS4A4BuR0/oO/kBbYLrmketZ31i2Mo2V7wQ7eJo5zuSeJLNQX
bJDK21683619rl5I7cwTkI2UHufUHScI/ntzosU2HPhdO1FPpg7agXf5olCk7/Amp4Exnm13glyG
xA7Nd8z8U81NuLY6YbH5YWJYcXRlKwuspCm7GA8CdUThVRRGGnDFrMo6G9x48GsXu8yUP0jGRAjr
DzOfv8bSxQDmR2Nh7EULKP4WhdieqbC6LcbrvLnVem7gFLKoASp2DsJDwNmUQoaFvJtI+vjgKTi7
2QE9hkHsT1aMrpI+SD0dmk5HhOkWtvNe1+Xs7w+bvLe8359OCQmIwz4nK66pRotsiGUmPPgQw7Wn
95L7WYPKQBmWWf3L1aWfNPDCT+bxGYZp+RIHNHOpiUSH/CLj/oBLfLx/n1HqIEoFx3+ZhEenGjPn
6wUyfM1qQrcMeuxcmSFEI22mmKKqNirczEiQ+5mRi+xXFyVjvuAYS1G3kRoryUsWjJGxzlg1QqTW
lqILESw2vaRMEObvk3P2+Kh4o3gJSR/+N0zeAVlMRonKZ06JoZJM7EZ+yAt3b4C+kWvMO1hpdipe
mYrFnJdWtHeT/8okg3VFZCxvPzLgN/Bg2jYy8EYA+9mHCGXiryrb5UhcJvnRrq4hjXmYdmoGWf10
tkmLxTaRVUdgO36yJUxwEi8v0QlECSi5e8SOPJfydeHm8pGVhMcB7ZzoS47pEpsL/ur1at652Mxm
7JuNZaZQ7Zq2VN1xNHZWv7gKgy8WA/Eu4hUJVNAzWslsBgnYZaswyXrTosSlr6pXnFG/TtNY8O3H
hOQxMtdLkwqLQPh3+b4QJ5Nbf3LtLSeH4a3Ffq14bIDRcL9efI8SX6RuP2rww0ERSo1LU9YVqUof
X9rEasXojvpciqQAasjybBqWJKwoMkZTabtVnsaZe8azLNKlx1xsxYRhSfI72jqWdTVweIDl6VGY
uQdjyF5GAO9Ply71Xovt6GG5STqZAjqkBggXMjAp+6OWt/8vD+J04KRoaShmo7yK/eIBvG6mzJWS
Qnv4w2yGZsHIjHfHky/RwnrcsTA9u7ngFiK8c3dRlcovjDfVScZfi9QAAtDJbj4Xc0UhtYj904IU
XETCwshmrrRMBxXR1x1iZrs38QouBroEvdV1ZMzaNk+rJ1Ea8a3Fp1qpdI4yglpC33MrzD1JFTAZ
zQbFwEOMih4iUgIBKbZuPEQuqF4yp9VhKElxzUaooiIFxJr1DjdJW7UKPxC4LfpiKqzb22a16rms
rW0gCCsflpWDpn1HQBhibEsBnpV++verUlQfOoOSnmAw/1wq92WgUJPfole/gIfBkVqwIIbeY1ha
r/NnhM1AjJ/A4IAi1CgHbkF6ER0PXtF4E+y8ozNK2Anmc/RLBo+8lwNI/pg9fZ8v0YDB6CpeyHZd
8WiXAn1ZK/yzmaJSOlYMeRVsQQFM81m0xqaNyy8tZG+RWViQm6AoqOOddApS/j2fFE2GVDRUNqjK
VsxiuO2NMCSgdTkfpdMP9aTej3nQSvYEhd5dUbpr+ADgprbREoIdiFQlTXr5HV1tTnU1J/HHC7Ax
BxLjW2aSBEXty4UmAuNtjCbtfgWQBn8L0hXPSSunucm0g2xov9JFhnA33lmL+EIXZSfXywOvzHPe
+wW+HyYxpvLYA4dlWCj/KHyBWxzvyjtTszBLCewdBh+H3IkTyWxQ/KohVlSV9qNuSTLIBxE9FI/C
Uj7jX0ro471CJTVFo3vCc4FAfHhF+d9B7UXKEOjxRj8K+r5Rl174ihsnd91qirSLYh2h3/rhS19M
mxPvLFUkkQnWLmFQ+oN4NTjt4X5Cn7YC3NSU8b10DJxQHCKVfPqrVrFOZJolgTzWbZAIWj7bIYR6
2WcPlFGGJXUlXSjxZTzTW+v+jwGiklH6cay78NAFl4BhsVdzlvD4ipluxWpc4spmRhshL6HZrk+a
tsUBtYqVDaChu/Qz+ota4PcfrMxzi94geW4e5Gj/e8YNmyzfZtrVKYa/hxMfMhbhJYhSByEDAfkC
ju6PZD7MwA51m1h/iCedw0mknvD3IouvavKgSsJGpnsjrt21clvUAoC00RCAdg75bsL+HCIoZaTy
AtNV2ne7BOkKrKt+kVpH64lvnc3oQlqh0C/r3l1oPXlcByqD/EEfb9gz5oWNEQiWaXl5f1p0Kx+u
MXZst/Dck0QxJj9KB0iJaQLgdhRVGS7CRdyjoasP+hRRpn+cC3u/5jbkrBtvImqi3mIaogTVrkzu
91+Zb26HFhcFUwwQO/D4re/g3H/OY8XA1EtT4tMZ9i/dv3eWk6p6avu6ZEbVekek78MKHWKn+Lgn
UOCjj4d7SGCFn4LEmOQFq/gi9awWaA5ZOyifMclT1TSxP1gtYomF3T4geoMojxRPr5GAJKsUAgFV
sKJGcGJKxMM43fBFzJGZdlJ+rjy2uN+M3/b2WRSS+9V3SnwP3EKDLJNbexbD/aGk5BDUhxrUS5Hx
OeBmXukUWi0+9GERImbRoJ6jwA3jGnbMiEL5Xzf+VE2rHmJZYcvosupdvSp+6ez7Bh1r3sV0crgA
MGWVEBJ/Dg+YeYy97BaTMusHBZqn5HhOnH2wYC4HKDf0ErR8NrSqALaWEV8Hx9YdzXnrYc2l7SFU
Sc3Q2u0pNPfcKXeHVQcv293N2XNRDa6jtlh+S+03xhAAvZxL5qAr0PWd7XUupr2h4UhxjHzA8ys9
jniztCaLY4diPJvO5BhwlZonNRAsx2PHznAdXG/Br9L9w6yhlxePaEmaLbf1z/OH8YuUrqHc1BRI
Lf5U+hMrK5a8SDu4LBGrbT77HSvlBu9yPPzOQLD4mP0ulBtEHQxdM40M9EJW9Pc3+NmUAzYkXmJX
kNC0DCqFPUynNcM/LfPc8hs3RM52QadmgLGEyYuI1WMEJt4ZT/ISVyt9yBis9t79Wz3IkMP3rwCQ
RMt64eo/kC3bXaDLeKdyYjNNYn5lsYlgCMTxpLIcbiTxENHJjQQomqV+0oSrnpT9hb2ac69gDzv5
ZAhRAYS+Hu5wWL8//pyHu2cxUMxx8vOQ02y1isTROEeZzQWHKBevPI263eULyyllEDaI4LEZuwqv
hItFpoavZ+UVFJ01aLEDiIROiIVABKcvqSoBXHggF+895SfEJtr0DhRO/53gGIOTuDqAacXrXpSq
EqhJYpLB4R2/0Z4ZwC0DfLR/o5D0Vu9fdg0isaIeEw2N1C36QbJtQFmNFf8RndRZgbKdWC09aT10
smLMXvdE3jiiLESDyMt02rkz4+jPSMxbnM7b2CgkL7sU2F5CpGCtkCOltnqJ3zzaymYasKupUKWC
lnc+lrmGRDuIQkhDm0BIT6DdBoqMeDsXP3jxzgZ52Xb7PWG2riPyMh3ygoTBKWOU+3UbqTQT4AtE
nF3CqdyCT+KAaLhp+BcDniREYDuBC+yiCLEkCXPcdBq9dW//2p5Rs09sR3nu0xr5x4ejPd1XoXUq
/zP114Z5hnTBvkAMGew2KUZjqleAkqPbXCk93W1iAO+7UIakC97IOtAb1P+NRrEB8OAJyXaTN043
SE5woXl6M5bEQmd0anulhpqwlEMYb69BiPc8tg0FIDwBpsRbr17FYkmeGK4KrpRdmWxfjE36dIXe
i2c3Whoo3yKOUFdFZJffr1LiymsaA1d5J2uF84rqHEgQwOlNsiA2OoLRWr2mQpiu0prHKW5g7GOd
nquZtVBs/4NyOqxoui3V2nIpwzoLy+ntSyumhW/Ypn0KZDsTNfvts1l6M/jepioHFcSHnBi/7oeB
5Et45Q0gGaha961LYBAvWiVB0bjqJjG+dCdPfPkPgSNMJucrSAiMCBP2HyOfRRbMDBueSb2+elUx
Yo2CiHWK66hY3eEeY2pLDAWJi9BkI8wjrhN9ULvPfRete8JH1Nlgav4GJSGLV3+tWUtKi45LPbrU
HVFZYJvR0gG/iro7x85tOQ8rX19STSm2AqAug6/Hb9HVrc8IQ2bMqKbDVYr4ayFcmNL15lBnJCeW
zSkEkCENovm7LOxlD+Y6QEK6jTwFqkFmNP3KOPTnypSz2ytHyzbItsgVVgL3oD4tHtkHylq7fbat
RKehGIPqz4t3gFXnCkG7EoZWE/vio6RNDhxYtbNzipovhV9zoGcXFeYAGCJSKqrsfxmU1KUr8yNK
DPRmv5DSp5n0u/dJCp903EgYu3qz64SfnwqWifFrGuIZlkYeyQ9FyzkvF70Uq3G8jzR8+5AI0qC2
3a3x0L7p6K58NeRLo6wvRRS1XMHa8Wq5dqff//XTH0CBh3167BI7ptdleCpmucP0kJbye37bfW74
/9Mxk107aXSELA1YjHAiU3EaqXcDw4o/QS9ZaFd6N1nQXDoUUWKncAwQxy6a2WvXoptMJDTNvSIO
EMJG4b+Q4C8K9lB8SrO89yrqblc5Qkcm7oaZg5AOJaLmrrzBB1YRw/mi0lkaa6/+U661NyZur45C
QBdwl2dWpKqllcSWr7BqROSBH6kwJqEWW7gY2jH12xHh7r5s/7lMg9rmiZAZ1XgVTI4gn+BteCLn
mSQAhcNxRuo+2NaFDwM28ZNvBDyhs58As7ipFlWVvN1+NCdtAYDlubtvE1Kytp0+60wjJD3Lp4EA
vLzql4ERP2sjH0NMS/cEf3xtE2g1Q7lIf+tFPKQIgtk8QBosv4IyqSe0qrizFUaVDsohicvvQMk+
iWqr42pHXgcRDG7If8HhrFxUmpERo45Q+un6D0SGwEo8J0qKjdihX/bA0JrcKnBXSFmpNZvK65vt
TxALqZQ8yMIlb41AATvH9mQWj8rILpHdniQMbI9YrIGRjzGN7Cjx3pkfho56F/kZjkfFl/YDMlBj
y5nAVEjNyh/EaU+DRZKRPQN7rxS8VPaECbEqaEhXs7AQ2SG/V7ZMJEOIb/9367osxlrpOuy+8gqN
k7F/Q58E8upPTYgBFTtZQMqNA+Fv3zsItcAUPigCkhRc1dpYLUashFCwh6VbNZhOAhpbsP0zcEcS
mfCb40bP66F19EP6VjkAId7UR8Mj/96BZ+SYCcKvEu0g2QV1uStqPDAmlr5fE+EJxhyEw8utpA55
RF63vmMjg10E7HrnrDV/pqOzikcrhiw0Rr4YdpiQdlL67oUfGVKMkikDPFud0Uyn2TeMEUnNd7fu
fZd/PmJLhu93/mJT29MySpKj4ezIq+cgSLCO0lYcDu+twjghDRoM5OixW3QpOF50W9CPBrAQWwwL
p7OI811Lp9neV+Fwy6I/BWAnxRwgSByl6vt2qdcZmyhF9nwrtu3KyySqFNi7zVlIwGnHudWuFa8o
NqVzXKSItm+dE/YlGG6QrZ1xBoKBotIIoA3gvB6CZ1dIOojugwn6+UeXXmTmQbkTNka5tkT0PEFc
s0OxQaDUQES50mR2JiCHSBhYuMebBpG9CHK9mNNOug5p0jbPHyGBwLHoZlhWB8hVNTLWTdIzTH57
fOkKps5dGuD5DRa+SpI/bd8xdGfhYVuVq7LDnNyXtQfnAX7/X3Y4XmfsWCk7RUoN1wy3XctA9zNs
RHM/Tc+MZfayzTa26s8l3b3FprzeRiUmKiZ9eli84ecGgF4+DsMNMY1NM5pKsfBEbiRSRMz1sTgN
c2UB93O+mWBnDv6WvG6/8LZC6YE31WSzFVTK0sGUFV0mTEMMi8Lhl1vZHI+W5euechQQ4aJALb7i
qK30bzfzfh29CngXo2tbCIdxQEXITs/y+lP/lJncjP8j3tBBB2FVmb/BYK2bLyZLFZBnL80+d/92
FTLokoGlzgv4CYd/cMIMzcVnX1z7kT4j6N4aGNKz4Vm1b50pDR5SYLqw1PGXoBhCDBEOsrYy7Au2
Qrzqy9yaZSCghV2EhdPUx5WnghgkPODrf92oQFj0K0je+Zue8/1TBxTnYBHFfkEyG9aXEOYdMwD9
JfRDsrEQmzAGOORCC4+VsRgUVGYNz2DRoFDKKoHprHj9A/zzZRuo8fP2xpyIcGbCRae7y9R1n1nt
LCkGevrnX+R3Clqg2HZ9sfpZI1C6mj7hOoi4AUuSZXKa5M21gyd0YODC4wcDIkQwRSUADPSfVUjo
HJGacKwbwMzuOOUAul9ETQwP4L84geEFMM2upeQ0dHka4GoJl0dllE/p3MU5bUMus+HQ0Ua5tFUy
dzOXEkLfNhTdglvDxzTjf4XBYLtaoTdvWeDRTAJjDEcxSYJ1PNjx6wgqRD+M1sI59NG1wFpZxWAC
ljTaWuOy8YqJ9bjF7mr6mhTkMe67DAyIQCq9ClQOWVuIBjroyvkwVfXkIpp+QVeCkMe2S/ulmu7N
4sLANA4cc1J19/KbHFDCure8zpPWRHk2hGo1W2TXUkXHp6VDstUH3RXBJobXISDk9MrEBN4NL4wd
0+Ag8b/p2/0mulQLXPzo9wJAGm5DJibQayHYPuIwOny8UGk6r9eGlcD3B39fjm+1UZ/KAnt/MRBe
ewXh7385IzWIeF77QOA9SyjiGuoK5Z4gNoOUaZ1CNojWqqUx647RAoAN1MbE1zGKSl5R8ZT91u53
ZkNwIijXnJtPRL1SRTiagjyrqCM8PY4/78LMx5vzSwTYalIpniazvydr8d9A47EvI+rCL+odGyz+
szUpVTFuVuXVLwqLnLm0Ckb4swPtCymCp7IZ+6a3hjq/pHdi2ADpH1ng4QZ+8e7jQ0XMwP4s3hn1
p/cHcV2wGmPieM7wga3GfeXjVvXmnUgLeh11eQyqpO1sWXt4RwxUAmPrZnft7rbfPzLFjGvMtX2z
ufLitBR5QXVcaK/GewcYqp1YM6u7+bZXjNJa9Z1HvgcEXpoeTg2FDPZR8vBIpoe9UKS2MiZ/7LMc
xRXzfC/l3nFI0SsrpFbV7Xc3J3aOxkzfuavKna3P4gv4pi380P38njAIJ0FKfhm1rh5z+Qz/OtIw
AaH7GscElj22tzXuJekZbGEUHb1jrf/2EEWeQ2HPKyZQ63kZ0ZuZRckA0X5gsMfhYPmsedVDjV3U
rOo5+2EHbqhMOCxjO53YMsH/HP+UqVexN9QWnas0ILUWr28Eep2TdhaOQkOVZzTBHPJmyY7CKGha
Bpl4ZtbMedzjWDqwdEh2rl+yw1K/uWUEpJQVhCK9Rf2EUrgOKIuZyrQh4mjOVOTpcbhYQbu/yqVj
0+clEQyluskeL9lgN7Li1bxbBiZooeCAZklg2eFf9JhBuNUB8dDSxXQCaCdO2eUATX8TwhZk2CP3
hjofazyrL9d1NqrKZ+1GLNgpGXRLeE5ZvxjH+HlZWpyY4JqbikU0jOjnWzCZ9DJy+jUlqvO3OndG
M4UY6RgsFGE7nS0GR+UiLU5zRrI06KnBH+3+dF20fD1eVLsuUz4P1HCXOq2ddLVME9MBl0BzRTby
opjEttVvehUETnTRxdSFKJH3Bjq6FyghX0dmQtIm8zAm4ybjJABWobw71w4mxvAQLt6Ww6cXkF/Q
PFNNIjb+g+zr1AED/UWj8QM2B9v8rYfAezRqpqn0C3D10GUBDHddOgy84hfUIbdsm9nVK4309SWi
NSgmY2yfrMiAhKaSZl4cRlosNlXSMn5rKS36zeytWdiy8GipsW39vQcSBVVFoyUE+YlUNcC9L5oc
Wz73KAvlQp/LFNTZDsFwdQAUroNOaU+uEBcgvrpqUJ+A2692wfvANjw9HXVj7cpgbuHfpKMVY3hY
c4gdiCNlyktSir5iovEnAE4LgEHcBcPazVRKUin6P1TGEjLUGyjI/YOV0gfY/7up9WrlCCL42EwF
XF8ePVJjJSwMJ0z1hannHmlNJ3AfqY14qERy9lCRCIujgIqKt89LPTBvX8SDX5foameaR9QrO68d
IcYnfZB0mVO/CocGqOKy+HcP2r3JwOVpLuORJUuh3XFhmtgg7U4iKpVE1b9zdjCJQHQDS6GkOCec
2bUCWeQBUiabj20kHeU3BLw4ZWB9z7JJsDTQX7mZIKSV9FZbAoj0h8c33qEWpLuqKkOVsuit2+7P
IVXDu1oFBPvD6xn3t6BniGQ9EQ6M0QZimwqbp4IZYBpd2X76tFbFIM56iMfH+xQAycRa2mTnHECs
EiP2UTX88skJDdB1v85spIcWhl2VlH9p1S5fXWZ3ixjPTFeyj5Avl/XTsIE2veneNLz7Gh0+qZIq
07ZWAvcLwFtGZyj12WFc/7dSQZJRAb4aTdAzEoO6ES6vgPcIpKJdqvnaBANp6rqKZtIhDDFx2v5y
GI4+gYv8Z0wpDy5S6hPQFi7O96FdIon5QMFA8TYNe+PThKrAk6WAz5zw0qE1L9MGMj4RzJN+2edx
XYCWWoFiZNcWOo9ZvOh35OvjzWx7xKgZQ0Tn+z7NMaux7Fx+qEI7QpGwInd8Y71FUuWtNGn9nF64
fIjxk7RVyDi9xYRZFIUKAuK//7AybilKS9IBrQaUxXhl9vrEI470XgvKmwGMZfdUNCoQxrzfBPAv
IEM/jEAezc3D9uCVrOHswRtvI0sikJpo/NdaJ8jrK612Qjzfjw5ZycLJpfKbzPoy6DfvK4drKeGR
CfRk4kJwscPkOOJcIXhlLC9zhCeS+2rppMnHT7VxnHzPkqbr7BU4J+8rbfF9euJkBOvdLwCby2Kg
o/rfDQwjAA+HDRKkU7T25/jKOfxJTfc78h4qHR81UznxtGdh4Sad97ktTMXHxurnCeOCzm+sYYyT
zDToZZlnHHc9Gh+cueANRc3uj0/uU5lSseX6PVJvKNM/s01zDNipxek9BI3dgjkt4c42Brb5nGIX
usGkzXIqO9twsn68gMP7xjBNqmIkzGL1jzhzA7LSObzOli7g4TWaGiMhebvXoxu+NIoTb8/7J5FW
XcZKsXDe3aU+ohHAKjEwxYvsHeijNndeyeQBqYB71L8FFwWp5hkw+IPIfqcfjEhI22KUT6QGsMvm
Z0xyXmPFK2B//dURmsZDWtyBbitCx3eHDuqHZaH/Nopr69TLIj8nNaV2V2onS+cDqnComBpkPMZn
nikRZYI1Aww60to2rwC+32704fWfAoTGWUjC2WNPowjNkgFkcUVQY/iRW1bGg5CirqIzW8WDK3Ty
cfMEn3Sqrpskzk+xao1wYIX/EitaZIJilsp6A1EjmBJOqp2kvOU28ImK3OMa3/fHBJAZxJViR0LI
1VN1Y30mdRblWZf81KFTSpVG0tYtrVM5TRDeN7UZFcE+qEcjd4Nrqt/ksgCjrGaqSrpYw8p6FJs5
e1UYgpChc3pyjcnViLCu3RXmI340KscFiFkvBoVAMU1moFmikZcMhX1BJT/4cNMfV7bW+Ptnr8gS
pnjjYx8vEBiomh6xr8R7WMJsqTgKqKW60RZFEtRzlmx+2SKGMiBJERCopSM6M2+7mGQTowXshgyh
zmzoChHOYp1UwWYqrujaAUyUINTPJwRqszrxQBls4KXcolzX7Dd2IcNVM7tTRTc0eDsil1ULOB1H
JT/nTBYB+v/jiUNnrGDBLzADrQzsCGG+ts0HS1FKYFc5rpnq/K3u0AwMnAOHj4Pj2z8AKgvjwKaU
DV1VvvE4P3LlcSBc2mXUPilxHpWqJktwchX979YNElBEg+BtJTs92xRpwk89GzCgDWupO68YrXLF
ZuRfpeCTJBXT+nroC6y4haLL33fSs3oD1VaVdhfbzp8vtXtWu5lalZuT2WUy747TdEZdzAEOwT0r
BdKnVvJxX8rVkR74Pni6k+0aCgli0IvH5CebkC4mIRkvCEYkLs2ECPWAI1VimHY7UO+WBhCulBVF
WWAO58I1sXNSpEh/enxmQ8A6t2LS3t9kr0EXnyohSaP5bN+MkZyfEnQ02uH3p03MofSgvdEhD+N3
NAYXA0/grkbNxqPnJ2WPTVV/G5hVhrx8p4KNgJGyKJ7vh9pgNoLsBbkry8/t81+lwcl6vc4qADtR
KaLrRQgNxxaQYKNG4yy4OU7Gymb0Uf12DDD4JRgm6EBuIy1dHERJ+EYim5euQSQ1mEUdWjJ1RID0
15sB7cuhs/Je/mkITECwzHk4MgM0rdfolRRJmesvMRjFV9TEiTtei5FYO/SDSK6o3HCTfEvFnemt
zSKOQnNLKiOiCSXs+Y6vy7LYha9xVOlNf/N4ZmHhVyn3S3bDSd8SAH4daoOzkKIs2CibHS0FTqA9
2OUbHImrONIF8CNEL3Vh+BHo3OeDP8VGF5NLyZJfmoYnEl2EhW+wswL1tvBCejecn//sF1UHFUpM
pydg9sSXsv6npbUiIgx64mLUafDKpKgYsFqIXOrV/4KUVxE9b8P7eAxDfUZ3tezse7nQLDkC8QrZ
kQhaxpSDw0ubCH5SF9P1rWjS+94a3TrfHqpwF6s95bt5ZV3+SVI4wg/uUbsbLCbis4pqDGlQu9CP
x6RtCxMcn0lTWQxhNv0Fch7lM1CCXDj5WTQH1a3FVhuQm9WHfKY9KNdo1OT3LmojzzcDrB9F5MsF
9SVKg91f50AssypdkgMhkWGTcopoUDwrmBd4XzkNmJnJMxAkLWuPG9GHoNrEJc18LQiXMlbnRLum
kPyoRxe1rvM51QWstdG8RMpowtWi+JfAHTUh0JSdnOsRUlLHWpEK0oP1odLUncyAjY9KWNMfT4on
CP5B9V1jSUunKv3mLVb+Z668hVrHbv9kfiXKrDAYU2nJH05CAZaLfCj24ivPBwQWWgX6zmN84/Dh
piNsScVntrcgg2149KVsFmTen6C9DVusu5uOEP2bR9NZohO1ToXjkdmqLFo145BjmwxE/VNyBF7g
R+yu1ykPofhX5BliqugU1FIIAUrnOr9YCgswMkQ9VOm6nEWyXB5oop+sBCE+EJAc8ecRyjhrosS1
m61WYT8iq+zAUaxB/KF4XK7GJmRxKDCZcqNrOxDLb4eXqxAeNz1EBQJ8Mc36dlUVWeNWfk9McYgd
VnLAI8cdsyDlhC5sdON5OZ4lEggFnxyWBgp92tNjLv50rxprvMt1ws220AUe6qK9LrIYXnE2mmfW
hIymSD4LJ6j05Isrg/WDhBWF+P6/i/XchZaUe50ks5NkecaxzpqRA3ddgOVsGkC6SImW0VsWreW3
90qZGelvdoe30+24yIARx8OdOMRZKFbhwdQGkFrzULTTo454MiP7efawABSYKiPDWduXV9onjxbh
3ufYeianjDVIVHUpfCpG/qJiKl/Zaqqb0k0LWuWf0Wc1fKVNUqn7pSU6rDCWi+Zneap9fEcjf2KD
TiudyoBwXG6iegNTb2siWN06CGV5+SvSCDmWWcobRVJbUQdJpcAWgyQgPP9sf1MCsKbL4qZiWUIz
ROWPvADBp/KnhuP/RlyaoRs/iSdO+xK09qKuUZuaKfrUO1UZOV7zhvZS1Pctr5llYqpIRuWKdNw4
fJAZ2LjDrrHpsv97mnKAN7jiDpR+3JBxjNj3BQp8uKmryMCkuY6J12fDCc+jenQ0TnOPm/CraClt
XdiK0DWDi6lhE/wuxn16UIMieE6YIMBGKWYezcI3Wgj4FML440I4EX7Y900+yvpGGwYP2x19xy5x
jlCBiF1PAaKJBEBOFDjG4ehVs+g/CtfZMW73owolaKuk5fnID4BVLE05lfjNkKCIOZVGcxHLp3N+
CTv0eTm/M/U/fKYD1gMoV/dPIfLdlCkpGpgtux8DEiXL9VPJDlCgB2ylj7saygxGgQERrL6jwe9L
u8x5fv3K8PcGdqcTsYR1lHRv2+7eZosX6l7xfvYFw105GRKMDVqeAWTL9hLrHvCnrEGg/MGyr5G+
a88rWCjB5GMmV8x+DH4tfykdLm7M62liNzVuTetDfMtJCu1pDUxhTEClDwm850Ar9gAB8Q6rnT+K
xq34aK7JYi+9flAkSNQbscuomIbj6FJdIpH+DEhNPK5cxTOz3mHaVq3pXGYCO4D+twL+rhFSuLPE
7oj1W39ajfeLp6D7oNGu6Nk7Nmz8guQYJdVKjZn0Bq8H3iaPacCRUI9VjZNhD7GPXZohoQImkAHv
pOlL2giy6BPKRqF3K1SGbkIebdlPg00V3qPIJi6yCBxHQT6vlllwNNMxjfCsYkQxqIVwB2mEK4wc
3Rkk0XSoJTzAe4D3oNFnud36XlCJb7wRCCkskpedJKiM469rFGq7mhU3W0qoj6aUVzcD7K1t9CMH
vtJ6S4/PSNPghp1+pZSYh9ssT9c2sIm6uAreeSdBkdmRrojjhusokGcETCueoNyDJzaV0rwtdLtg
2jkDblAD56wPy6zZvVbJ90my9HeVTqznJqolpAyaW3pP29+XpQYMhZB0CylCpCMKVUs+mF1QR//i
Kzuh9x+HhXNqj+yjG5SPik2vYI/pV49b5KYD3wvt8uo2sDO8zOP3jwhFXTkjFOMiDd+Jcg1b4L1L
TlsC7VPWa/h+xs+HaKc6Hp/NinBrNYlST2ihSZqcIIUg1bkvh+yeGUiP11POCgF8OkQj3QfXCtYC
szmVUWbzd5iHybL0PJNob4DMo8ZX/Lya00kT1UNQDHo3uGZN231ln53uke4I8FZx2i8a+EdRwoyn
MHp5gCNDsB9wi7Xfm6dmHcquybYntvvPGh34/RSJhp0YzNyRmtg4eNOlfM/NX1kZA6LYQNena30D
qy8jkxI9n8nIBRcAF1PnrRXTFU2vyDUu0OZHnuNnl3/0FTrrm3XbYLELC3CsT1dF8SHIExMwD3q1
CXdrBXj7L7XQxhBcpHpMhavy+zqHM33nWX4I7XHfpGLqgGchlLiWU7LMZMHDqgOBIscxLiTk4Bzq
g0zYmZgUCIjOH4Wlouj/9m8ocwBG2MRGnhPNMizgBFfEZoi20b+YcvCxdnEnjnQdW3MuikvuBj/V
reF5hiFP65PIvgffJxuWZ/OSfUUEHzSQx0Vs8hRD4kjLZlVMDHzbvyUc9VBoV9SFG7nemgbz5+Fs
MfMUU5/KVStjEei9BjJaQB9zr/MVBdpm9beTeJbWP1ySjk8OFjflv31zWAvaGrVDFE+cCRbHWO20
LoHAgOwDPeBs0mF9mzXORwAg0NkjoXg4IzL7i3x6l3JSM3vIS7rcfkAQalFV9pLSdrUJto4aFuqJ
YXPsta2r2Kaxbbd2Ndn8grood6rmrwiCC/ly/42To/41e6//t7CMPJm3aKj9GlsDPjy6HK9vJosb
YVoeQL8eDGL4zF82/ma40yJNbl8AVA9vERNuxmh0dIkU0GJfCnzWCJH6A0jj01Jdmr7jU+aYkGsl
rLJWnguHg8DD+BHFMHgW/W8oOEolp6tPYVxvcpg3jvf1ex4QJjoR2w6k794OC5VXe+kAJofvGLky
aR9isLhuVa8z8AaftqiCluxerV2todo/XxC18bmXQitgD/98mfPmYnWSOLO+nCfXIvhT9pNntuds
LMWiU2HUzMssk+aoOxy4iIbyR7fggroyBjXLVLic02OmVjwct5YMlrzh31D6WdSrwdjMlbhX9K/4
CzCRsUDDf7lWp/Ww9qGnOPVGBliQyG7ywoBv4zXk/m85sgXisqzmtqr3ROcb6zWgcEflIonsi07U
Sm0Q/M5Q3bGlEEOg9ZEo1f3JTD64MyvRMML86qk9zlnmSI6OhqcAx6ZnohCJbeSeeqdO78sODfO8
n86ZqmdYp6ns/0VBx8ZTgP5wcRT9Mdl9Bo1sveTeVI3kdh+TgAke5ENGRgefzK47ukL+fYvUN+nf
Bdud6/Hiiblbp3ftpd+fyt+LMmeCT8pK4YBIF9dxIbd+NcTX/7Z4HgHLvjJVivZGz7C1S/k/luwt
PTnGoKE9LoAg9PRwtSIVKAWB3yqkp60M19mCtZhDP7s9Fc7WfV3I0rEhszbWySch3nJ/Z9pF1Hci
Bibgau30/aIE+DZ7PFe05lzupCfK9/VPm8orJVbNsX0zr6O97jzrUq8TUWOSvSur28IWb06DrR9m
0x6WQxqE30stdK07rCcCI8nkkMcrRhmpmkCk84nO/8EKJvGB1Am+Ib9MxsHFV4QQAXmY+LCCfxOf
M/+TKnMNZ3StOjVRImmemA4n5oy5OgdTKgsk3WIIU9BOFby6jtLfKjBrsKNMPJR38GiUjBlf5QF/
Shc3jKACpg1jqBfFK0mLb0zVp2K8Ug02+UEluVy8QBJa+pd3PLcsUNbE0ZtIQ5VXiYit40asBGjT
034Zd1VlG7zh4/gy/mttr/eLTBbimsNiSeYo31YLosw8VQNr90roTxO6P9oBENbNhGrh8z+Xg6lg
ZrBlgOtNKbggmQ8ktFNpI6JtJ0RKwll2coIocw1FYY0Qw5koZg/ZNeQmkMsHbdLTJGkSaVZxVjY5
NiOy9lqG8gArEy11f+2StI7SPu6oojdClhzoxUsDIkdt48WkTBNocfVoxY3XPUckMW5vsDSjWqsL
xqFRcS6Umh2+YtCMclbDyUHHdHMNiqPciH2aRz/sZ3L7orrdyTJ9zh2lllNpujmc1bCBp3XD2fRb
uAnXagpBh5/qEJ8HVAgTETUMT2stpkF9GST1wF22AZbHGWOKYaJLGxEgXCYxV41Le8QTpYyRwSem
5SaPoYzavYmOq/WVNBEC6N6RZb8oo24RIxN6Hrcr9lfbhXLx1UIOpuPw8y07brYUN5Y1l332Gs/Y
A+Q9D8UZ7poRB5LY9K1VLcfH66Td9E70Q2LtjvKqDV48FoU4ekeVvZwdoHw3aQC35TT5oXJ3juud
zqdLQpCfrCJ4gtRXscVtEOHyxGzVzJx4aNDhOhVpX6Sm20gzQ3d/lWx5hZg9aaY7NylPkGKDRW5+
9+9+fIHOg7+RYeF7yrops1lxDy5619KNg9n7zRgmtoWYh6RUYQ6I+uHJ1EGH2ZOkM9B8P4qKWNML
bYMcrwP/vAX0uzZXQtOSuuqcMOptWyJH/uUL9IOEcJj+Mywsa1h4UCk/ZFLSKESjkga+FpW0Fdq/
0QWyfSgWz5aQG1iCiMsjH5g0OrL6pepj5RfMoWvg8q57wCC9M63ivh+IJRdGPm4E4/hpzD6ivJfU
X526KvPFMnY8btvDTT98jFrHfgdjhIhNgoNlS7qi8NMTIX+KEfKqPYMw81mnRrczavcRTAj37jMP
HnbbskPFlrJuVnovDn6TA1AEaZ7sYi9IW6uvKSI80mi5dNtFnbgo3IiRYQsLRZ1vq3u9+j/UvvF7
oKrKS/7Sf+eL3DjLYZSpdtHob1Axg1jd2R92xmbB3PIywW5jEPymgp9KhdHIkTnFmdE2JsiA0ghr
jdPYDxDGgs24ufKoKkxUp2pguoX+tVYnw5bkt76u2LQBiuPPOL499AKwOacqzi0npSuE0HLi34k6
tGViJqXqI2/b9chGE8h0CFgPEE65M76TDVr4vX6FOC4/m/hKvUbHwRplFMfnNqR0A1m01NWOQV5y
b6uBsQUtzIYI5QKCcSs7Yg/Z4pXNcuimhZ2UqKV0fSGz5QJCzTxWeEHFGVDl+KHE+itE18Hbsq4L
sSB12ryWBASad4SdnvWH3Po/pPs2cqIlY003NRnzowqlMkpHbG2zXxZ0zQCd+3X4OTSZ58gy2Vzl
uyU7h4gCwZJO8796ASiCIHLDK6YiyrHS6wJs8knwY7UxHrCfRvHPKI5SpVj6bTYlGhyHyXLlTpTP
++dEXRiVrBHy6tCnUndyZMYhOHwSN5pjCGZ2Eh/vVWIoglY3+zSQ/gURTkexNfE7hfcgqZsy8XGL
BfCze0YsE2zkHO9LJoNF1uDv4aSkMOjb6ULzljxzIETCo7bRguJiVL87Dx62o3CxvluwTdbWOl8r
EYk0n8yMNP+Fz/Z59bowck1rjI5/kggNu28rWmbtdEakpu6aCYEHhSEEuq/edf3utYAnp0ewUmJ+
LCIX5y5vRGlDSQdio86AK8HFUnCawZROKrTum5VSS7h9JKfGC8Mndtrpotl2ic+sSTwwsdPB14Xh
uB+AN4UM5JS8nnMa/vPaPUMeoTsmUf9+0L6WAG8nW3iAPxrnUG72oJ+ja57gIX2SFJfWmmvzN7kz
5TeHJlfmHGDWSEQjbmlhUw1+gQSDfHH5hRBPsrsH3bypRYxOAPNwq5USwa2YWWcjSRK8i+Ip65Vx
KP0RJ+VdbhEs6p6ijR5FGtwX2LC01oWz2QszwvCZs9ecNcKwQyPz8fZbGBCsBkMrfQRG8T5cad98
1btwF9n7PiReCfkJUhiqSJSyr3LurvZqAw4x8CReGPmujcPca5fEuzTF7RysyJWAC1Y3OYgAY1EO
pIXfc3FxsTPZGAFQ6JNae5zsFFdIKTHalSRFVEcbVk/EmKkEXLGYkA8sECbrNiotdDZKDSHnJ6No
kTxg8vVHsXn96XIDRewJcy+1tnwEvDUf6gmyJ8if8lYPD9qE2JPdTgNoE+s10Kee9T8HgbK692rL
FXd6KZc23bByI6VOs4uQb5q9PdiUwisDmA1Rjk93JX7BsA52OfBL40vmhjIJRIgP7EZAl9glqd7R
y/N3b6uAfZJd0mE4cLnKj4+ouIZSmovYHQcCuVQ5qIZF1R7eciAECnUQFjK/MeOIv3T7zTQ7cXjf
a/kB5XuXVFdCDsKuMHHzdDfe5cTBNQpSUnO2ZmjXwpU9lam5uoewGZMfktKwY+dnzsRmn3S8Zmas
lQzV94w4wxyQFYWZ4LSOcgvkpF0vEhqZmBtwmn4Jz3sLmXsauY7Vjz6/05JSQAXco9FmLRWG3Fn3
Nb2tFFoPqak6Aiuz5dUFx+lROwkrU15MKs0afOZ22A4TVBcTjES7V/CbdD7xRw1XwICOls77qOXk
aaCd0SIc/avoKm7a24xrPCC8GtJI2YZlGTsAqAkIDCmPYT6SCGlyD+8lqPkSfOwau2dkA7Mfzv5d
PrrM5atfkaH3yTxs8Vy4yOk4St/t8+Lyjj8k8grurX57COwTzr9lASCrgqnJGs3W2FbvwawAGYRL
kaNFAOzL/Lj/3YqplrTjZcIRDHGBvkBYjybDy4Kn7vrdl2TkXPd+ajbkvpHt75Vi3akGk7X9Y5xC
FaQrCn770lnvDuugoA4Ek8QP5jaMU2jiT0XM5BcitnjIAYUOmYFrnqn0RJLh4gPWZiVfoxxdOFJh
/iSxrkaxhfEvVDpRdCMQKVZBsKuU46zXTAP/vP5ju2DPc/SJ1o9IZS3gtnmz2LNyZw8i0/uAhq6C
4n18GQevDPmMNCGTbH/o3804oROh1u8C/8lksMj1cDT5zBGPVlO9ksipxI6gpURb+RQGmNGziTbT
v/z/Fg+HuUmlfxPLASRKlL0LSwuDzgZY5Gfhj4PEgY4LRe/yCh8fJiyOUGlx45HHIHQ/vRA7njsr
CUSej0NUMP3PAPxvCyuNSIpOQNsgXIYxPHrgIsEQ+kiaH9n907UfcFEH7AU2pamuMruxbfBHutfx
mjP1DMhy+YXPeoE09Zi2Z3fFQO9tkLzvUg29AGzodeayPUE9JuMkRl25rrj4ZAoT+hL3x8IP+bCL
B+pto3nfDT0oo6zToFoYDCeT9HZeYH/uUe8sILv7CUnbHpbeLDoQNPNR5pX8GLMaQf+PWo4WzenB
ZkcRzWMuo1bzmbTm5Ac+PuU40+Xw8rSBv+sSfYoc6kIZcP3MXwCAFk5I6Vtslag2MA+KBEDN5UY2
p/qgqh/EB6NJhWGfuAPMqlaZlRSBfxWe5CpBz/XGcc9HOoUyg39KsFnnRagozJ4697QmFcCOcx5d
7immpdK60M3EsNF7X8F64gKJBJGq4x2N6GMduOmMm9H6mqn5GKdUMzzQDss7fC+u6TZKpsxhHKar
xtIpT2xezV8c7tqVf5NgZpj4Ea1snPD8SkW+JoPYvKxPfoIzwrI4+b5NEyvsPfKGVuPCgu1FX6lM
pHrqf1Qz0FVAfQfWfFMJvnr8G5L7wrSa6l1FhwYnZi9YfByDgvAM02xSaUEHkucgLm+zZ96N77gs
jF1kS/u0evRngWAdYtA5wodpAzchPQpk7MCc2Y6oSsX+GKXAmRtC2K8IIlK2jtxiRDPpyAbsY8Ht
69/EbNwRnbGG1sy3GJ8ot/9RtC4/ZfmkTQ9ZgHDjCAu79i071VCQmc/4tNqdh+u5E67evtPB8RKI
ieW8M4wXfVc6Y98Yp5PM4P7kWcyDyQ7fPMGAd81HPatgUt2zOlWKmpP+8l8TZv7OPQOVV3+s0I+S
FiIO0Ad1ySuTty2Gh6dDh68gZHRgDgg2dI1TR7vVoGAi0oAtYrOMXRCVfBk7WL1UVP592OtQJNkT
Kz9Rr8JgtN3wv36/vYDF5RuYdFChB6C5ppBk9FiMZj1TrnUDIXRHzrKR1vlR2h5KjGa96cBzLCR8
RnCyNTzR5ET+DIEoNO4ZSpvplAZF/P93dKV5ly618XVYYJ4HiP+B52Vd9wO/GIV8aYN4FceY7NKx
nyAP2FlI3LafflxLvW/j7C4La6SuQhExRSRmY4jQfc+GmClD4rVHB4fp7zXUk+LICSV2bWqik/2c
XmjaXR3SEHnyKV/wUoAEuggVMCrzdlGMzOT/Ak4h4VVoKYeY0v8uCTT/2uAksae/17KN1eozDE20
urxXIKqvjrrfYuMgfHRwe3fERX+tlngBfspmTZH6+5zeo/KbWBj61dkgGuCWHZv7dQuIl5Upkgoj
na88xCX8Y9lXBLR3GWT1eXPY14tjHxdL4RFF0ycrAMNIA7doQBEeE96V+H+AUJFtLbqtVhuLb3Fy
8GM6t2hy120x31X5g8rCWQm+EyCXlK8Vz9AlkBu2h9MKm2NO9hT0AKherjVJOPgzKaAS/mrQ8D2l
sirW6mzLp7a6WKaK5wPu08QgmzppBeCKHiYG6+TimPbkf+xjwYVDhXx/QUDYXRUBhi0RaPZvluha
mH8XdKiJyd14kpSZG3u4eswtY9Evai+15N5fliz5Kf7MWDGLPyCqYCBkIMVlvhLePfTqWcvHO5q9
ebXNGZxU57vGjrfPTBppAJy9IbuYTOXNEJIQhamqd3dQ9aeIdJhpf/yi01lva93L/K5zF7ndGSyk
yDQgAdgy5wQomqGCQEAc2gNX8OfOMjR9540JcjkVRAFwsCiaHhIC+KfDk+jKwxvG4uFNmYwnhCDw
UNzAiRZauxA4y07UY34oL5O/lHOE9iTpqsUZb8+miMNoKRuLvpre9SSjWnF63d7Q+5ZUemPJJG/u
RK9JeFfFhxZpVtTAuW0koraw0xGrVg4L5DZ2p5puvxSOXpvCF7cw1Wkhv3zvuqV/N0ZFb8WbPxKk
0O9Ml7OOXohmGWDOTz2VD4AS+vyVxOept5nltLPzNyUCH9URNapsmVd721SCbBm7PC/Efn13vJUO
bqcsn8SkWxiCn//tZ9ZiUzCbQANa+XQNULLWPDQCHjiXrZYClCYy1m2c5wjBHQLcxJji4QvgyoAH
JKeGs/rElTFo2SwK+FXMX9acZwLqLGHUmCsOHsOR9/V+juwEmq8l8Q0vWdnDZmkkgAPLIavwNXEK
r08a27eXs/EzUia9naLZ8IAJlxbN1SV5qbeZU8YbPczPKZBwTz5AqaouvgeubSdexWYjyKPWHoiV
x2gk17JZG7/mMSydM9T/ZNYNoJyBMxPWaP63Et3WldLJ6z04nSFnPZHcrA/TD/cXjkKFlOBPYC0l
EBjMML8fNyvXzXdPsr1SPrKLpS1U333qORnKGKURh+Wvz1b1UrVrkdoQKHE20ADRAAxf92VWxHiq
tPl0z5NhDOyq2lnmEyXRBVUDVFga/72Rn7REhOqsWUZqdGnON4KCTwFdQEkJ6R4AFOPsGPZXRxzS
bB04fUdOCf2WLbjLamSZ4tXMIxP9SShqnwWV4qrs2wN/SBYsdryfKeB92MqRpP9Wsokkv0R94SvB
ajT+OkJ0IiaGHYEr/ud6tOT+uxYOwqyEDGU+t0EnH9wi3kDDl4oDEDsXrQxWvA+GezPC+IJRBzxW
09rPGhRPXKI0hCBzRbIcf8KJz7JWcknXyTevFDflqZ4+2oBiH+P1IzsZjZWdL0EJ+RqK/Su1s5WZ
UY4DnGvOGukQV7PUadIm6GVd+FvxMRoN+3AXNSzf8YUlNAIkEp1w920lQScjwmRLsPhXOknMA2bk
eEKZX7QWA8Y+9scGrTSa2g4xnMD/nYq+km142WxjKIxHHhyhdCaxuzsX0kgxb1i9S4h0PP9fHEw0
WV3v+fj0ZOMMqLR6AVivKECDikb4uIarLwTAuRJBYHlKv7V+DumBcLiITxDdbGDfkEe8HYpBItl8
ML62sMz8URuP4C9wbRVaX8+Vb0ACovHMW7EVLEMJgqchwYeKl/AnGNBQESeTLyVJ0IVeuMTNGZjs
iATctbSUsIhJ0TVhUmZ4vssKyP61TXXMFDrszHThEBi5iFNYeVIiBUBMXNznH3uU1q+xJ6x+f46G
6VGy30Y1aLcK4Mdb7XLu6+DY+nUBWtvT2eKqe27fAgKJRBcDs7Ou3XjqYMdLw6ukvY7r8yIiyPPO
31jn2wc6V4LbpMUtO6Pof6BG7vG+bFo9sJkNKYVFgNyox8Nc7y/baMIZnR2QX2Ivpc5sPsSe2GaQ
Uk6Yqe+JRxzVU1iFYP76MSjQl4bPmpGIX9Bm0YuUJI4+OckRA0Mivq0EMlbsl/gEwWcbKs9lpFW3
kLot06Q1cWGT012QbcK15KEulQavp1zKi3586ZXq8Oej+QHOmY30Kz+Jc8KZrwi/l6rwTm3lfjlC
m7a2oaj7vRW/CWw3EjbifTGh1cD2fD8S5xUaJ0LhI6Ked6++9pCkyViFbCS8btOBaaPzN7YMEF1h
Sa8Klrg4P4DaF9V1nXo8b/zwpx7k5QNSt3rfnGmt0RXxq2YwCz7skG9Q9fdbkxS3tI62Z/Fh5hca
TSWT479YlUEBf0qaNJQHWVioaf5LO6Jz3eR3CXgPCPI7QrCeAY+5RIaoR/c7aqq/JXlVh602ZLUM
1Buye6zfD+EB1vlfl9fvFAU6Hf7RT7L0/jrcAmL7mA+1LTERwMYffrCmX0hi8AZasejfYux8MLZf
L2lMv0I5WpYidtWJqkiwqySAjUI5FP/4QmlIIRpqrDKgbYArhcyBbXiFVijgnJw6Uyn7GGx12orm
BlHCXKvDZnANNAvgq1R0JmstYE2GmAvqqH4ap93GeOFkhYY938SYqY5tyo4I1Xa7261JO9nOar7G
ZF3CLdd4kqpfswnOu8A+w6m2rhDGIbRJyKR1eEeVJkPnc/7c05io8nS9gzdgE4Q3/VioH8ylOyCG
D5fkhzTEHeEv/UVK1EUXjanQKchRZkQZdjzOKzBN1rCQLZKn27O3QzyjxcKcvvZJSqJw99kKRaEw
jQa6ezBX8Y7NZ6RcjFgZWHJjgs8CHNSGAqeshPM5iSsAWIn8u6fwB84caxLOJ8FLzQ7/PNk/6wbZ
s2ochNpqRUzwrll3SFw1wu7obMUEeyQTSH1EJETWGt8i4du1tdPIpKG7+LQGiLX3eYvQtYStq1jR
069ZLV39QuGzdvrLfmcHETSfo7cTRgo7xhhYMnPE/nQbsSPGsZjFjCLM3IJZH+jYBQFedrGMv9MY
rtgCoVcan5T/bjpROlalvYgPQPXeSVduZRk5Ia++QYc1NYNuOytvolXY/R9KA0STX1+Qh+WinjiI
3Rcf/AXmAnUUDjq+vUc3uqTqHB6adlKzno3kMY+iQuSLmVc9rj6ICaGuD1ColW08/nNs+VAAYlyy
mxzuD6bGk96Y/b9p8Ir5du+YzbPcyGMYnf1k/pzAdWMGgrhhGpEGahjnkDldpwhYUYLxpFyFiEm0
KjlBCi0k1RlHTacrFY2ittY0KthMVk6yhGkicQeX1dXR5/aqAN3ETkyS+Ylbo9d3YacNkQuhjSnJ
zqfiYFEQi1Hb4CZjW13Qb8AMy17qFTRrYQlC2h/NAFs8qZSzIKRM9QJ2Otzw9i7LQ2bjo0e8/WTg
6B6OysnuwH9+b7lKdAmv6q6AmwgxYvbmtn8fXPAKLzdcYxhmlLfoc2wvBL8tDGR8lGGHHKwDMoP3
my+ZrZ07xok0PgJawVRAy41xu+lGWo/p0ZRZCEGbEgZV15iVv2tK2KYUz/sTOQd9t2pYiMxWV4Tc
Xr7wlpMFUGOKVNTFp7AxfWohQAqfNwLCMDZXvzQzqKqAHkAVfF/wrtgnBHXEoR63ESfaSyg30CnR
KpIsafxXBUNCQZGNsJp+/GZnffezwS2L+QpaJjb6792BFyQb0PdTjlxdLB8O8kYHo5F9JiSQZKoX
XZ0ubqMJyOoK+yz0nRjIrVO61nzo5tlOFCfCmBtWMP4mjEVJ4UzwHMNDcg2b3Wt4pjVc5oBl4tfM
3Weu1I01+6tTlWvWfCsIzyc2RjgX8p+kHmjCMg1GHkxvEJV1sjzrpkZlL2tLG80h74TPty7LC+DS
J5Np90ZLiFh+DuVV3dO1LENL/89cMoDqf4+CAv7RLHoPnElTt2JTV+Aik5dA/xqU7IrRi23AGDXm
i0yW/9L+GZNNTRuTBHHg0mhurg3NQQKnvDndNuQbJuRbufUvFWKZ8cQ5ODo8hQmJhvby56L5HXuD
ULDJLrsRnzzhIYJGvsOQhTj7jDmZlCEmAAc4tXHYdNgk8G0lZvN5zk1gCHVYbT4IcNpVJQRbX5Zl
kVz5leZxDYkboKhgFIX9KNsd66O0je3+90yBwLidvJ3OXHiQgCdy+A7Wpt3h2iXcWN5YEaiwP+mx
0OuJw+WP8caxuLAWycGoPJQ3gOpq/ZW9Gdw9l1Lrd77AHHxeSjmpRyuH8J9iEuepORM4OnII9+mh
dGKK40ggfOQw1ajVhipt/qND97SFErNZpJhzPTmdSPs0DcfzNh2Jgnk6WCvc10+DXxhxMdgWFOT3
vFt4kUEUmFS2lG1PWO60A4Nh/ADbXBGLXl6kjStJwtpOTitFLo2B5jIaK57rUojJbc3umPhl/+uX
HM1KnokDomy6JeekSCIeE/dz8mS3IzjwFcd+kMB6KWesIDshaGUfOFCkV4sGc2VwGFY1PleLuTQl
iF8n4ulhhD8ZXa5p0j21TXj0DH9pA7z0wsmCGWs3494K/NcfR4napTZcT0gLZcMy8LNXTIJ/0zHZ
qkt2AErJTlgIcqJI4VlEIHeMt1kKTfZfOqiyKNTsiBMC1R4d/V/tAxpfbEh2pvq+Mg75R5lO6QNi
mgUX4KqIv+YtSvKs1xw38sWmBNWeG+661BwbTdmm05Ed3m4iUryEVW0fAKjIF15kv6S4sdSzkUnb
F5hi5KxolqR1n2tL5e5NgWmCxADkCsKwIyHaJrRtqn1/6La2JNGz717zFcM4yYgyccvdOcENbBRr
yplqi902T+guLtPkUcu8Se72L1QhdUwmGB/l++/TsuZom4qFidRJ3kQ/gtsHAYAM8uY6SvjBsm/B
DaFd7LePE8TyUb28b9S2cB+Aw5J72/BSALlW9GcGartT/mSfAUG7zrpUJV6xGS3FM1MgnJ/D+gFq
mbvAJ3R8HsEP5nZc+aBi9Mcg8cjWtoy5o2u17oW19Yne0SX0ORYzf3tWhcoGBMR9I4VupMjpYzRt
HGN1KZnQmYaKlJIypS+DrzpeI+7FQn94EWu2+3BdNKMKmzZYUBV29tnjj33PHBWXBm0k5oj9qUst
1x9GoWLvc/OXYCH/UcSSYc3hz1iNBSBMeI57w2zBriDpNqSvOk/Q4+I4IGJEuEd23OrwXPoCPbfw
ZJr9/gpcYFExi9KZiTZ/ChK0JwdPEJr1b5hv5RmuaKHUJqTs/fROUtCW9sksKEhWa2e7iiIlWwiX
kspaDxtX55ih5DiqSlNO2tDPFim9v4/msWV7aL3VYEvV0Xxr5dVoseG0DDqCACP/k39MZS2whIjH
2dkU9sjsuyLtKJwVMSnx2+db2aV7vhQ8HEacWqvD2rZ1BzXis/5kzFFegr+sDfMssPwpD9PilpCz
A/rLAi7Vj9NjwfhH0x7ROPnI+ZwkPCQ6FOmX9uVEW5ojDg1aFFXfcVx33g2F/k1NAVO2afmnfsSi
7cmuS6wHXig6iQbqy7Vi0/xPe/VsIwcB+A3VkKYkqHn1XUOrZfziiAh+7ZATr+jHO9xT7LKJZcbq
G9Y5SrTd7+ced1aGi4T3l+6urPD+Y/uljg0kqwuvIM6dk7O+qjoZCYmWg3mwoeKBTJa22ffxPIzB
hJPIgvMoMsF+tX5ni04RvFjk3/LBxRCLKkUwrni6KlgFrYrd/dKz9mw3HwKJt0+qxJtXnhMEFiah
4wZtf0yM6NytqItDlJRG5XBy6EcfljYPZeZmD1HJ8mzj9IsyL7X6Ju8oykZ0lH69AIVPqj1hlNSr
wUBq4EdX+7i+bkDX92k1xyULwJWpkUV78l+qgQ4ZJbvgGAoM6k8zu4wkV0vfHmSHuVNFRJt3FBBd
HdHyiIHi+h5tqwZS5vpoHqKgn6k6UKtwYnasVtVBmvIsqz1I8k4Ns2oIIpfViHxbaQCDNg2/wAP3
oHwJAna0vnaGtXlfDsxo+7Kg0OrJf7ymvXRrDPJkXsE9762s0YY6fe2YQkSho69BrD/hrhYtNr0Y
1mluH8/pBd1KZq/FwKEEJQpxOhBVSjniDH/9RSYHZiCv5oAjdWCR3IYog1l1FXiZaxs+LRjsFBHa
KOlb/RPiGmVvmKzYP1rXCcycP02vnXsw/rGnOXe5vjVA4zFjCaCLrqs5xsPd2mtdGH8iCtH9vG4p
70nbJGuGoosodk5WWvdShCl7M9loAJY2IBa6rYlCfF7q0O2urqwF3Vp4BJfGbMRMCQD7PRBrtEYY
EEGQD7bUhuZo/MbCoLRrht9TJ3/hRoQaKxJ/TLI0tUNwuCsM1FYAGPNBNK6rej86a+LdGe4LUHB7
4XQtI8e6akTFXKlVd5zzYpt3h7X67WkwvsAoTox5xxwbpWXpkDja69GrsVRUpMLzCD9sDzT2dGw7
3ub237JDvNn9hMgSXV9kGsuPZGHrPI4xfw0EbB1omh7woXfWoerfo2KqgxRDQoAhM9nSeAg4gSON
c59W8vPOxn5GGNmEXxWNMcWEWFJgRPVG/iFzXkb85nfeGC4VjMNm2LQg2RVFaof2HyiRXIbDVgws
xIOPuHDbmk5rTqVD47lpR+NCvtnvbVYkxXzQW508giP10AUw9yCH87j2oupNMJTCQF/zbKfTYz4I
mQkjLrRHJW5qBPUO0qEc91AJkHPkeUGoZ3SemDC8eSoIgGTwosqjnB7czp0GERFkAVJ6bUY4eZOe
yNnmrjscu7kGVB+M8ttKWUrr749Lk3XOE5pf2Y9BTjYQkb/2Iovfpa4rOI/xj2mCv53cK49lkvzR
McUYH2Fhk4OBRS+ixwPl97Hm38TZHB1fGVL0A1CQVqiVEWWj8YSyRTYshAnyHrqsVCeFmZpZ+4oG
IBRdRheygT8+58R5+vPPVPZllVBURX3F1TgbLF1hWS+y8Hll6PWhD/xojg1m11yfJ5rDxu0JJ8Bv
zLI2r+zNwVrpmmL5SgCyVPJanZrtXcCSFggPS92HIac9+G/jjKyESsVpnjVMwu2N2OIPOCgJWdNa
c/is9ZE+yP+dHuJrW9mIk67QkhbI2l2YWE2SJMbdIf3rul29f8DQVMhDnuPg534POwKCWUByFgbA
lMkq9pEw31QijIUVsRIxX4cFIsDLyTTJYwJtUBnTCoa3+kmBVUyGI/RGmair2gVSjlmVD1Cs1MOM
XW8p22KpNDhGMzNdDEfJ7jCuWXA5Os/xjpDL/ys9Y3YqB4xdHae0/FRUlVWlYOL9E5qlAgd9A/Qs
NJyOCJTwyGr+0mTisiSIQfZp7tYPhosmmUNT2v0nDWWwapyldhJyiQeLgnM7QblttsZ9PIEZsHnT
z3fo0krmPStkuc1D7ayub0ZgcgBEoC/6cMhAtN4C6khCbZ2ekFDSc2+d6ZlRis3gEaFeBNEhliAR
Y3al6fIzW+MO0CQOpb66QOBcHiFcwYMW4xCGBL3dtQsodZQY+/nwrP5zYJtEL16fzqA0SoMqA1XP
h8YnlRV21CRfLPbn+HXPTW5ma3Ojd95HiMXJ4G6JR1LO1pBSt6AxbNTSp1Hu42rSigrFWMcxtG/7
oqokmlUzcLGezGUnC4HKQ4luIgzbGlwzEMm9BPVEm056gnYi8yDWgVolQgerZPmv9XL6WSy4mJ+4
k+tniF23EzmV2TpasQzEo35xBXSr7Ff4hLl+dg9vxVTHuEm+oQe38IF7TZgFTioxAcZzDUv+aNFJ
Fy0HdXOK7rDNwrF2cwmTFIYafJT2gGTyFx/n9ciF+Ijpvl9OjeV+rIoT7w2Ljam6EWeNcZwLEgIt
HJSbFKGdAmXnOaQ1kDy7VVkwVfDyuj1pUTQN5a8qGIgKNStkbKgqYhurbGb2i9XKv9U03g7fUFpm
OqpgKknrw1PtDOIVyG7i9YnMN7GVwz4SknltfqQm5SxaOMSXI0x1GobSI2cb5Oq0y+dXbhhRl4Pn
YanFh/FPXYNUyYcWFMPrb3tWLb12Gru030PRJgsHStRQnwGZe/UVt3segrEUttJaTWCpvknTO1Ax
fym327XXz8FVdcaN2ZuzQBCSzpnfnjxdRLh1O2xSoajwK5FWDE5S47P0TjFW1YixHeZctDIYP4gp
AhbFNezbaS3zjY9NxJpeQucMp4//U/YbnnK9fBgjPxhYYQipL8aC29TqcVeEnPbD2S2g4/5lv3GY
J3n0OknYrCm5wbPmKHewXpE0Ix1Cqt+esl0j0B6yQUn3HQzLJhf8sm4vIx39cr/VsTOq7vgTVfgF
EXuNrU/R/BlWObW4kXHCIGYvvB++WdKJFiTBBh8M3WTZpsRw4fZddIX16lWWY9/Yjqd1k8jrquGH
hLtq8ykBsZeg83fd8WU9d2vD2xqhDAVFXrCahYVfXwTWtPaLySf5IwwafRnh5FOyHqbAuCKoPVsj
1I5W/RSZ0Fq8LKPbaCO+M2Wne5iM7VO1O/IV1ADNSS7FKcak7Dtqa5kUDm6aH9fdBR9ZwSD5MnC6
vsWtDfES+AuNcJFZlK+HgcYhD5fS+oQ6wjcjyZJ6yxdprZsOGf59i9XEGfrNNkWRm3cp/xoELLFI
I+iG8E+4VoP6ZHbc0IDLhn4N3O8O1Ao64LOE6sW5zx4g5iFpICkmGa8MsqEfBiP2+FvQqzCnr+CF
FCJoVi6Cvw+s6vrmYmvcTF0lHaZ1sbXH0XdmTUqg3pGPwLIAyExy8U8V2FvuueEjGmOmpH7lL2Ds
QPh+csdpri0hewHXMtZpLs1YNL+1Hc42/4NqtD0JFWDdgBZq/P2Qu6ytKYs4vJIg65DCjrdfifkx
dnGBqolLtXlePrv+sB3iY9oB/ZuiNp7jPtft2zxWLsTYujoPisUkKBb2p5vT+m7WfDbQhqTCcKtO
6JT2IWkMTHASxsOfm0DzuXKaRRsZfjaPS5JTjehmVMQX+K2Ly0L2LLFos/B2TdEn92/t9kjCQJeT
5UyRWICQltwFbVtMXpbZbioJGCdCh4fuy8XeIyVwElD1cA+H1Pzo8G7MmSCA+jmbTE3KJ5JptJ0x
8VlH9sO0AKyYk0oB0K3Lurn4XEJHs1zn3EJMHhGyUr55Ny5xNJ+S8I6g7+jkSzyZ6LoxxeV4bB7B
33XRBIvMQOZoLY1Gxtt20wrMgof6mX4hupVSsbqVHeZQxYW84hzriEkj61XpOWJJh65zJVXZ7ePp
Xp3/NdttDW5CqxuMk3HHyV4yu+kqMpFNy5T7DaZe8ShOUVGsK7nu51PFh3oO8pmZwmgjPtO07Upj
0LzMjGSgyIBN/n7EoJ3fxm67Vwq/3ZkcxtL5BY0jgBHs9ul8YOXATarVmBs/wDUo9mHUkxFrVw7B
521RLVyaZhOwxDBTsUohhU4Qw/nEJ3Hn632KTOUiy+jbfUnKoRzSqSzTb3SCX75wxclaaNCoZwtT
H9wzxc7wgI41iakIap0zyQQs5gytfhQyFaq1XevcRQWIbDwcAI2sMU2ALMtiUGmBTziI/VbmKKX1
S+8NGG+pL93Bbl8nNFiAhQ7llnwL1h+vJPkMPCVodWwgZAqi72ewpyj2j42IJdrFMUuq5ezXP2KF
G3mNtdnuKsikyAyNc5lzBJ/OR9HcQ2QIlrSBHl+UCuGhYqswYMJWLAMYRISiMjtncNmhRUliSesF
QrGAN1KSeTO7FEY2k/QqycvViw0Gi1RtTBMMWFL4/jLJ6lfoi8PmuqAMIX9np3h2sfhAPNLiPxFK
alVa1Pdc0cD7wvtvdTEEuzRQf3WnAr0Q78c0lyklW2GoLv8UHzHpgsuPz0+cazSyYHVvD3t/XMwK
sAXar0dp8L3IJpGYOsE6IgDq9LVKuQEnU7yE0J+TAg8ekdSQFu4E1Ut5p/00kibvfmNHImGGu+SS
c6HGDkutCAJU4Bg0iun9KJR7n8q2mHmr976EQNnUr5jHKNYZZGzWzVM0HEVXGvPittBHb1HLLm+g
nKY8C/s+QOUbXK7hOI22YRp4+XevrnKmdl9O4UtbvjCAb2LmGjRlGzA6WZm4/jI/jei6psDk6CWo
8G2GHd2B50C19Jp0coYiElvD/rJ6qCTVKOMMWyDf2JxiBDFdpm82im3oRax/7C0Q976roqfsp+MW
UFa8ryQ7UXJ08W2xSEi2r44f6sV1/4ItEjyo7lN0tirC/5ojVyfoofbrcwN9jF9kNXB/5zhnK9vx
qbc+q25d5aaHei7vTkTv+MGlFZhb1jsQ6L+HJAYr68Txfn3Znz2RJ7D1jV5BIpMnuyUh+2AwgkNH
nJtOAsCvrQ1FWuGQQ4SBfLNxV4zuk5RZcOGb1Bm/ul/9nxyyETc9cnJmHdH/db+cL5wZvCccIpUP
HK1mjlIm6+rUz0eLzZsvklOeRbJMFzNROJQWXRYLBtujijM1hSqjf0VjPq2vXTzixNLO2uMhazMv
+yUV0+1EKy0LtILJiSW3SdT3G4L8fN5ipNVdU4B6CTtz0fknZUXlFdHzktK45/ntBgTvxvOlvh6W
D2sFWE8Q3ZNKnPoDFqK6cdBx/co8ITuRK5uHgvDmUS9XgczP29RLmz0nTtWE0R7lD9OeDQYkCtkI
kSLZn4FtlkUDP1dp5qXp824do/r/7hr19HuU5CRspp0wU8haNWsnbJAgkyBGTLnALgR8PS4M/PkB
R4qIp+kdcZHAH+8bSu5i428Ur+r+/dpBt1UjmxYkTPA0HXau3syQCydkXryOBCcfvYimT2SiHv8Z
tS3B7Ao90KYKJwaSQH5IgEAJ7AM8/otXopIMbZZEvCZLmbNud1heb5sCspD9e60M3dg0jzNwO5jY
UDL9X6FM5pJhLBWOGABp0EFtrVmde4DCPKjq0oKQXludq0jOC/vbu8ISK95SYFbE9H0mFi5XTANY
oI9Ft/PwnmabwOvCC0fWL6G0mCJ8E6qMhtVbMQffr85V94pBC5zk/a0/bD73FylGgQav8WOXU8/k
ABV83ZPQVSpcSXgHYMBw45cm8krqfYuMTN4ciHAlK6TyyrpVmcsH+MD4MBT9c5ovk2/HOZZQ9zny
4xb8ic1hHdm1Prv/C8uBgdeZlyikhVr7g8RKfdrxCcTPBRwiUXKSM0pOSHGWRgSCM5hDMxS/a9rG
akqWpR8tfkK/6bllM/MKUH4HNxFuz5hmK5WLJLxJktTgeAH4UDCcxCgEbiieU66P0o33HQlNsT1z
KYJPmPhRhmLzenbM8bnJ1lmn+iCjnv+3kKpclZvh9nrq26X0w62V+YQ53cQ3174hSvSV0VnTGc9V
YADoyU/AI++Az6869m26bj1v/+1M6fHpfc1RB9rAhp+QVfabqpQsIybJcG0vdjF3b/tq6VgBZlmW
CrPLZS7g2HGmf82KN5U92DbfswCQ8QSZaX7X+VUIsmzZmsxm5luvBGca3lShDBsgEFjH6Nj7aJ+L
ZM3P0cOjl6gUNuRIBjtiI8yim3CnwwhZruZRlwhTOFG+A7aw/VYecmtrCDExjYk9M7NVuo32TTtd
ZodsUVI1VOwNg/hf/Zenh8QaC9a+Y5/xt3C0yrl5hcNdhxIxrboVAZlEpAJSSvnvWueAN/3MAq0z
ltbrOMEZUbCtsPXOyDmC4lbUBT9olNRHuVm874iyTjyPG26ioepvH8mByG+/XAxuBWecO7VxhLGB
bU4h5JNn/rwD27bYstEXyWyeHrlO1axDIPnJMJo/hwNTaems1l39UIG3JjRMdVV1u+Jbfr9OC03h
GrrXr2WsqNFb830X43J7qIsBKSCS8c9oO8GN0jXm3XwwBliHmix/eT7Wz6Mk+uq+XlxrdoQOln0I
aFU6yn+6y8XcYRQaavyFcANMK1pTVQ0kzEn2+Bb9m98kZIArZxXKv4zSOanEsIMXZBwZ9wQ/VRlk
xe9RIdaRmFVp9a2Ykm1BFCPvnlhSGj9P1BaIMNB3Hwkx1cZOvDf1wrdALRmIcsDhq0in5P8QDq4P
RSTXCIEi6Xbkr/rxhjaN08M21BIPLPyK+Xs8n7NniWkQzpYQ4JfYzXryVYvI20vmBaPb7d8eRmDX
eP0CVlZSd45FGYOnLW54hmMDVMbVWDIX5bld9h+KocskqrqisJ1vnetVHGlqhGpEdGQXcZ9qqcv/
jM0gj8XTQm/4gJOvrsAlGm2jp24nMq218qWINnYemXOBx6WGt0vVFKdpxf7kcfg4HEVJOTC1/PHE
MQg1LFidYIUXH5hgf1hOuIyOcjDtvh8pOkjjEwhdEz8UGvgNv27oEkafdq9WsLZSzQSPmslUwtcH
xtAa8o0I5tFIcVlk78v2svVx9uyTHXUbtSXdYMA66dbeMci04j2fgOvNAkmgkDjUX4njgBVnrxfD
nbonW66WwC5KstPN9KVpJRnAGhCgzQq0BdCV9PWU0J/Syjiza6jgZsCbCZdej6UDGLmo4XLbCi69
Ni/8rpC5lEtgRlAf7m5NXFy9lzMKtNdvPIoi0FQcaHH86vF2BoPFamcUsO9tPaGNqmnolgusRlNQ
v2ZcKyoWdcdCUvVL53XyRDdyM//mslXczFHNvBfpKhNyYx782xvXR4T1g7KikJsohLGatNHSs6Zd
3zQXwjEXXinJ1lt6QFF+m1dfJrSuDKzhS5Q3UZSp1hbaj4qg1EAGg6kWDyNOOoJv8XZb5fDNy4/X
Ku4U9/BoAla00l/pa1yZQSzXqA2APGnfR7xp79UyscgaWc5aGCULzVe7HUs7J+N6J08TDEnhFjsk
+4zZPwIdOUtPOCj4H/9fMwQvE/K0M0ihLWaFNBdb0SPjS/mDbB8nK2DToQnII7AmQqAooF/ritIv
q4LcJFmLkDI/UpOPKg7zTdeCRvrsrFHjivwqpfbYc5NxVh+gLfnDUieXvozypvhz75c4rC7KGYiZ
qNnYMKc+LqVBTdnlX8djzPd8PDzL38i7/zqWxcReN8BrtkdcIySuvv86TGGf/3wAd6q2PtZPvMlT
GDyrUJK7VZJBPCmB7fxySrT4sPA9NgzM7EdZ8YGnk9jYTSOU0ivHwafFFZEgmni1UjLwZEehyhWl
39rCm/Wm/72iZWZ9WYTsNXzXRjQoDSgmiqeRK3eyiG2c1xb6KA73G28UPoF8SBQpwF108oI89F+q
g11DqsHMOANFy+4n19y1xXvv2vn+l60anqeXfikOTzWHjPDeo9flns3f4T9WUW45ofOC+tm2kYOu
pvdbW6+d1+6AmWp7VCLx9NtLsyvLnhX7zfxEMKL/zc47+OUSzj5ljyFQlKcBFna6YzMfBDr+16Ih
t5ui4YElM0J8Cv8/eQweiljBS0+ynrshCzrvAaNYrWB28hRcYxPaN9bRoGrTw0WXDbTnQhMch2oG
BmPGLBosIX2hhqrhUdlBrOyMIQl1yFU2OCBUxSm8Z4kwqH14w2a+PMXDd82s5+v8uPxdZGs4NdlO
kCilnXCl8ba80OGE7mncX/Jum9A7jRaferuJw4fKIMJ1vH3H7GZuUDas5/HMHpXcpulvHpkGiA1b
Nfa8LDXPgRDKZOm5WGUo1G74tgzGt9ofxNKm9tLdrSLLzjSVRO11DoWuLnksbQUlL7pbBC1U/Ldu
KYv6GEqotkQWe4tyGfR0Ng75/4mr4vT9IU786CSVnG55DMXjWyhxh6DBGIMdq/IbYfZ/b8Gc18z+
wtSwzOvYFaDc/zdgf/prtyIl13iBkawMUzc4ORrP0KWUeNrc5fzkbKz6ZuJbxdZbQA7VtjoLBSDI
ibIF2akYkxHRkI4mLd+2Zpd4P59iakxL5qEDp2HC/lxA64HLLl9WTeOtVSZS441aSi2VbZGVI+9w
8yI357n3q7qE5SDa8c4c+E4obFc91WGk9NYvChFrs8ReFUJvxfoJiGqRsF8Pc1A+U+GnKDnqTAbi
X2WV2lt2THUQORUpXgVUAP2p3U6U/XpV7er6PDXxXV6b/yqcVSyNOx5xOZKaid+HFktpjK4E5JAY
AxHpWFnu+d0FYFi29sWgYG/ZFK8s2AYTDptA52ohIU/WvqdFmNMfJf7BJlzPhVB9KY1+3KtuWNmt
pO4YUrKDKvoA5e+IofMvt4PyaKHHDxQKY2RbopAx/orRPyLGYbQBLZKYsSHWk3U8TEKN6JbsxqM4
L6K773kTRi+LStUNdu+pAs2hQulRrTup+IG8b8ZXAD3bOcDG3UsZQSAQGHCQyYDcI29wPtAwbk0Q
C243uu2/+KQ27REgIVhCMYPRxnOpo2lxVB+3KY0Y14EdAM0SmK7it6aBajizxiaOvjVeViBISeep
mz9Il5befie0Gx1g0K2hCdikxeg3ZqZFwmX3Xm66VZn7Nqz5e3MhR83l+L/zUuX1fQcMgtAHJjJp
L/n4/OxJoSjobgooDWcxK84Es32ocppANite6OrGzPQdq46jnu9ctE3Lcp3nRapsSepC766uNsc7
ETd9GbCdJoJ3EreG5LkyJVY7B1yuW/c9OHpfRXwzVfQcay/A1kj7BITkLqLdd1wZIK/Mm6lbf2Zd
jEduouihYbmJFSU72Il6351cf4whO3798u0/J1gsl2CWlLegrtzsxX6q1oF7JyxkbSQLsaD1/TzG
fsF+FxwYKrbDXU67+CSKVuB/W4iA4ayKhbf3ra9Kr2qDSLhuk9dLRsAppWHZdIqlcrqImOGkVNJs
ZTHEwsa6pbonSRCI/MdvLKE4Jk5LnrsKSwpnEQdv8fzyhf8Wz06Yw4UC5Rc+TO8gaUs/ezcskWaU
GxuLCxG8AyqRNvUhOW6glJEulK7kdwoQw8IC+a5dFYbTzXwmib4YIqknwjw2esmbjxiZeFQXdaIQ
/l1tny2OmQgSKjV0w+AsT2z3NkymukuK+vY4sLornxud2M70PAdhnziwZa1bcv+VxYrkdVnFOKEc
G5ojBQIiopERTFSl15XRU/msxVzBnGlodtIgk6/5o3PuY3PkaBtT0noWHj8/ZZJBC7Ujjxgw9GOO
5MeHdEiMB8qpUTXTJkt7wmxe562uLipOqaV8vcCOuYgiimzSyJvHHYou57kJAhfeX0eaE+diU53o
6t0+0UzoCMTB1CZPoFX11B21umX4gyJBsjREI3vC6sF03B/xDUxeOtKOtyQViFxTPDw16iVhgUFG
wUT91ayTM2JQCBGJJ0owoyCbuurK81PlEdUB1zS5U756yl5pYZAqjgdhZxznZOwlNaJl7gWR8tg1
w8Huf1mJZhWWY09CGhPBzY371NOHuWv7SN345J+a3koesLGxrUHpFSs1FEzbOjY7PkaXFhoTEJ0S
++vIYDV1IOLvP+CBqNZE75xdgyZen5hRkynxvJ1v3pqUmJONuN5HpDz3gP2ygafwZPuGaLyf3zaX
3Pq46JURGjNr7aU12mYOdt/rOmux4OMRUNHSwqgptwLAACIgw9DctXqTNaZPeG+bR4VrfLOa3ayZ
ljk8Cyk+FPuTyMUNCcDUDHaeVJUkwH69Dk+cWQ0A9SAgTYQq3G96v2LADXdiSZzBKP2aa6wtkImo
QcFBUQm664kdFuytvg7J5LkyJ3p6JKsog9zsvQwNPdZOK1/HjQSsUJTl6pN/uvEHJkXGQIOk8f/X
rzvMTpMHkTQKTR0AdJ5hT7x2vyrgT1qnmPNZ+TBLFsDhDwqMZSbJRslrxFXWhO5WZ6JbTxrFaBxf
O0xydMHngG0QXUR/EFzKkeUnq9+aI+6sX1pYU9Q2YZYX5MvbjdLrLgMvVMUXDRAv+6q/8s1BMzwM
z+NBrhUbZ6AedkSnl0mZortCLNKRVHKBSVqH3CjQGlW45RevvUEoigM8aDn8BYFsuSJtggxONaWU
EbpsM5Ci7rDqanl5JtX7i1+lKzUny3iatLDyA/z780svnGpM27GQZBYebsSLlvhm8VOmnCpuhLmd
d3QQ/2+yieTMh5Ml490Pv+ZLGR7jjpiVl/Q0Q1e5h/Zu14ehJbu0LZ/K/HxQ5+TcwJZbyIgHpBV1
Qd4bwj58rBwD2wqT0yrViU5dUS/6oFlmhIn3xYfyRYyG3pi9n+Z5hXDsBeB3OiARv2iOE8Z6MQjA
uRfGYmngbEs4tUn4xlSjVNnEvw9MCBCeBH7kfVHgTe1CilbNEZkkKvMzqhk2+Pcc8/B5Hf39KTzW
nYd4IFpSfWMLKaxf9tH6S45WNNf8LnAS4AmmrXg2H0s9WXEXBpAWCl6OQyK83wWaxXQ0dJtqV+iD
YKbHMETDsbOYXA7AR9v1GV04HRU83atWNsc3yf5F+IoJRpuHw4bITPnR3+TUYDQC5ByECbcazGJU
3YmC3DO7g8tjkFpFsI/6irdrr/laFHIfBfs4Rd3+W6LAlyVjnf2k4WWSjJAfLWBt34WbRPhAAJ/b
Z0XsLxzXE3P4IpFJbgdxX0J74D0yy/c2bsde0UzSGQzTXxNe1zEGqJIcP4YnsrXEh9p88PCLoQW2
W5UOkdmwDnR5NIROi9K1u0jIM3I78qP+R5hWOc3g97dG4/vb+9PA0aNsEjVAaHzpYdFzxr6kLM0L
66JLASlOx6Z1cMH2KzqhY8nbMZlUzKM0mMZv1PjgZUlEcAOvcZBbP7cdbG0gjdfZP9Tw5ds8yWN2
D97Qep+fKl8KkJZioQizM9aGvTyr9hGJ1ms0IwNvWRfjIAuM4pdBBrkEnICslrkI/H9VjlODnrNT
3rg57xWoiNRA8OYp1M2VKAbsy8DpHPKHZBmT27X78f94MYT7P9D70kKi/ywdGDwHHN8MuBpwfQ15
GXwXL5QVfp7EvhHy0xyaLk/QhHbOTpdq6mADaMxcLIHQQIkwSFL4Xy4XtaLLS46QDgsLrcElKzDd
juAmA9VPX8lNWJ39KFiJb0YoGzsMnLvYaT3dM1SCVIWqLV+p897VL8WIz43oIi5HYHIWPQkJqCoc
n21rTMfBjhrXuXwm70buyVqYDz7oQViUNO34Fi9Cb1kBaKja/I0oKJxNOIILNMwnHa4beZDVbTv3
48uhZYYhiHTWnTIZ+GxtonSeg4au1udhFrxkAAND3g5zlFmSh3zV9zVE5kU63GACJTKl90IA3TMU
XCqalmKO2jLWHtcPPGq7mGXbyq2dpWTrJyM/RpNKyswbgwMeZzqpA3F+TG5LWiotvMhSb8tRkwRH
xXl9OyLg9cfpGouhAq7O4cLrFasBrMsWw96KtoWy+erAIuNC8eVA8W1s1Vb2/8RHSsjBiCkANEOt
5X2z87AaPxlrjfjPCHV2sASRroDTW9QWLPF2rCFLzZApAAGq/ezscuABZoGtjtzkp/pB8vO0HsPv
R3RFiiWmWk4a2RY8alpiYg4TnTptB1OLzhFvxozit0njE+vECFHm0Wv6rcKD1VHPxPcTIa8GIPZy
lil/M8QMJWExjIubvA9y0dUROWYKDsUuPtf+C5ZYF3tw6QwWquARkVROGqsLviZah1b10H9iVYJ3
9UfGnPNJOXrTKlMUsaJ+cu0iIC7fAQCLDW0pcqUka5JaSngynLMUASHMJ1l2yYXheCiXlvi8CYOF
nq6vl0/ziPU+8PvuwnRSk4K4HdghJN3Mg0rEf24s/pdMguop08QhRTLumtGIho71CyMeHChG3p3v
0NqGZyOGa+DeIPhb0RVaQnxSgTG2K4uqAGqlYxqQhShax07OaJaXGHKL1Wkp7PLfAuspFS606+3p
JjspImeDYdD7wZHvlINLYpyAfadBFnqGYduAdOZaxJZ0BFydNyg5ZPZQwgvK1y2myHRC2B2sLZn6
FuLvyjVrUe7JCgiqf+8DDtrY2kSSTZEqkIbIDKQ/M3Eyxdfwdn+L0i4xcWaZnDRbkUIx0FULm7zm
L5oPOoOrvpYQyORlMyuiD6HO+3GXREtQk76p1F59hskiIRI1Pylc9MU/kTUtY8o7PYyQM9mCtccN
ItkjYBAreGGBZ8yH8Yl2t0RiCUJENocpYloGqhrjt8QTJN03QbTIJaiJZRUH2TsedEUaz4doM6Jt
yJ5QtuvEsePC6GmmoijVFUUTfceulS3GMZtuta0emaZUNeaXwOy2x8OLhAGUWgqlGb7VK0VXE0xZ
nr4CHB45EnC9bQw0kn86ZWAm4Fbo0cnutiql0478Poh9llaHE4uhMdAmzOcBwSGfzxXTNWDT9xtq
fsWd97CuRdjzTGwC8mcgZOXJdcl73neGSg0TD9XmPsx0djpTkiBIcAFAau3dcoNzPLNNIWc/QvCR
zc836bkBgVov3Arnd7z5r15wH5A0/i/HZcgH4dGaB5IocChaSPxj/6qMOm3LuJX2Y4ZRHzVIlUfn
9qbcXA3XEdNxWxLGllz26lFjgeCL6ZlTXiurp+uukNBta1OO29DHjh9UYO8iaNwFpT8ng5IylGfQ
RuMQjnMyKEdESgjRpKmUQLkO6e47BFor4/HD4HxtLL8e2LXmBs2U0sHYObyTZ7O5OZHBgg7lQEbz
PiJ+sGRCbdTOWfoo4RVQOx8wBthspLnLObdaGCKiDmlk/7IQaRkrzphSkKfrPnZTkKSdb6NIy0Le
/XI7p2JxR1diDXHWQi1jCUFBB+Z8QEcEnSa//JKOUAYoi7JVEmSU4higHgMKoYRqdymCZ7XrAqrC
6m66G6LKh1WZJXPz9ub4dEr4wZawdg/IzkTugpie5dKNUO4GNvvdyDM5qoC4vXpQ+Lxc3yAccPGr
pphXFRxUYwvZTWsVhx8lHix4ozF4kQznMiv3XpEllE12iySuKa1JbAz2XTwCQC06Cr1HI05AEayE
zOQOntKMr49LkKpLMYvyXVV46dXgUFSAIlxQWD/nk6r0eX8Fte2OFL5OJi1JD+cGwoEQWIZwwsGO
fXxRv6TuMeJVp9XhCLAo6CtXRL7YIBmI45zsezArk/PeXUHVEvK1PknniwHmwjFkJCyib2JGZS/l
/kcy2cG6JlArrT5n0DjsAr0zhBzC0ocGZ/LFl0WlnXDWWnPTdef4BW1tj9xnAJfg2+0SSs5XR/L8
IEZFhNTqrz5Z1fcUxwql83Xxm/nSyT4HIk+QsD4YUYWTjM2hKwnO2TiNbz/oUh1PIWq1VnXqdcse
9F+8y9YicM+7StZsVilh7pIlQoWvLStXgKZFxDIbv16U9bUEU7gL+JEe3wrNJQ52F31YN2mbZsNt
bNNdHTAUcfvCeZytWK+F6i5EOy39C6W3dgUaeHYY8ONsypqRfGfOSRazzhL23tiTvbIiXjcZP9q2
mlqc/3T9wzfzxd7D9WwdGD4ZLx0DGXy8N/VdlXAVOgK+W8q00nDtNx6R9wE0DH7zUzDIMUEtx+GK
x3BA6LhaEdcNyzDZONvt4myIqMV6yPLgbSarXF5eZS0F2IgjIyMvq5uoVRRkPN9BG2UYaT0PftmK
Thg0+1cbxzTlM77nvb66f+oBKC0NrehfdmShYuxnWoN+95Q1PAu10O3GCYgb8HKZMRrJpqblP6ch
9wBkIIfK2A2NowzqjSyBIlJc78re9CsVb5faU1Xsnwd/of5r+WCNyfXN8PhnR1Z00nNIvUMBKfGx
tVijHKxuIagfU+Y2OaK3c6YKo6oUtVhGcykVLWeUdk5xq7S7EtnzeAjJU67VobCULtLZgL5Dne5T
6gbgcQJA2JLXsSAnZqfq6p36FwXPqkYrLsiKwD/LEaQXnJmklKwOblH8e46cXLxXIB17PiHTkHex
xO42eoM8j47nXmP/j+IsGHZ/neV2QGAfKeOJnHov6ad1uttOf0wn2s1phsxybdhwZPrfwchCneQ+
WG5ak+Ef3W2A6Ql6ZLA9PWeF2WIErdp/wRzqRYtKvF2Ot6tovzcOuHsgok7jf9HgDYVFXe8v3VoF
8l8sr34YKfgGayXjTdR1ThC7sM94iD0mSoszCBqE677Re7DS8Vm3ee99BDizdLhbuj4BRion+pr8
Sp7jw77wBjhvQsBE0l/W9qggJ6xULlF517GNiqH2mA3NSFmWTGXrMlpQx206vLN1ukL7v3e6z4h/
E2F3pgtv5OB7dgzs1dbsusV0KUipy901Pq50tL/NKUSQ24BUCqNnK6V/2R747kla4sHuv7Pe+Aan
uRLWwhGSkI6mfWKCAOc71bG7eFxClmtD2oY+FnnrjWu37wpWyXSIc2FMqyn58N/5H2fPfm30oXgW
B/h9X9W+ZdsMgGK4jf+GmImv/St8b51YgdmbET23RiRuMzZj5/eVSdse0ga27YGW51Yi/E/4wJdL
aabL3BZmbT4J2gSB3RUuXUQ6nZJNsC7caBu7e3Py8WSs6f50XbC+UanVKqxOdVVH8p5nWlOSVmzK
1RG8yFqlAsoe+L8/Ps9lJXdCMwp0ZBILj9jUi2BIKMqCb9Lb7u+JSN8NCwVPxCbMbaiXFMUwYLbQ
fvu1gs1XgfbCJ4yYU95+UDRJdRg78f/k9LvMUkX9PRdv3J+h9SslQ3fCuELjX7UJbO++pQAC/3f6
bC+w9Ux095AxEhMRPynPE+P5egAaI1574CQ9Xre07+Rst2WcniYcLVRe2xwJJ5Jn7M2oy6R2+dbV
igP6rkzH6pv7iXhjW/qrkEmIGKQZiL4M5KrX9D6MKV6QyJ+Z40XD/gxNsnk5PkIigt3cTA2VSbZv
X8Ktq1CEwRWHDXtEBENIn+ejIKHTzdajVsfWHYXcOeO9ol8s8yZ8vzuKnMMUpEjhK7vow6HcNWV4
oIYCQmO82xBh4e5K0tYSZ/UeqiyNvsUCxyAFTjkgYw3YXfbmojOWhM5KvgNAsdbr0xYD7T+ETX4a
dLsddWBm/3jmChe/8yIGg5Gy1pFpso36FmYdIpFuTX8bNqg/XE1ibWBr1djKjqVpgwNnROiMJNoA
y2BGy/Hwr3eCm+ycrSOXUqkZKUcpd0TBpAmAq8XjEvGZjTsEE8qVLLjyG/LHmhyz0/XbOpgnItGF
THzIuLJUvEABmIa6MqhSfl172BJYcPE+2YQ6rsKP+L3M956+GPiAT6a9QE9ZnXUGkv0sOPQBHZD5
t6/0osNVSqUVtzWIDuBVcpdcg2uIdMqbunLrrApCeuabyXgacx74dUDcKbPWfoEj4KyQTkZFb16g
Kca6xef4vJuPKtuOgD//2MZ2Yw8UGf918wrecfls70j0P5klo2n0pc6OCQA8N2avQ/8YQDFYr0Bh
yJYPG7L+PyMMP6vH2Jkk79GwwPVhB8HoQANd0cGmCMirvZ3/0opIytP9sOores2Oq/8EenTKuRBq
TqYZ7cZLuAOsbhN+HxFp8K424j4PdnCO9Dx7d9NgjK08WYCuo1O28Sj7fU9oH/K6E371r166L0rs
/3uAvcjT7UXh/TQBwwvwwbGt0iqHhGH2A/7beIc9qKE2HY96HXTwV0XascFPr9NVpzIoDLHN23VP
Cylu2b+qLIFvQeyCcoaSC4//3b/UVuGr/d23iYm3AvNXjY1sbmvJo9d8iCBX2Eowib9EIpbKNrRp
V7xI/qgZ767a24dgbR2s0BVP3ipo4ZD7U19vmfcaN8beQWJJ2zgtijD2fHkySJ+dhDk9dt2x8sN2
3CaQIrqlbYOmjZE1Rqscdu8AZrJ1w9N3X9LQW5n1JyjqlsjG3j6VdhTeBUu9DdsPH8pedMrDVuxL
yplstZx99FnrG8e3pwqfWJnIG5JCm4PPYEx6I30tTicunWyP0nwR+rYO73HYiKJEUMCg6amU+Ptl
Y9K1P5v9cp/lJeo+Cgb/GfikHLXIxTd93W6xgVbOLBp/Z56k0NJy6xJJWglPBo3PfEuX2DgrQ1cd
nGrPk6Og4PbP5GNWvGy781tUizg0qA8FDzCtDOVCF4XaQAcRsbNgDpApxTdqaBQea8JOxs+1iXf1
KkN2kEGTs351AiWqW4HMI9JH7rChlUgckvq9GoLz8MRKrr4Ro/ElDwyYkTa9HLmV1MaGZmWXl16O
k4KFrMQrNQYldBNpSzTn66Qnbw7i5Zqn7cK0INwou1QmtnzukKteIyo1gILj9v/kWtRXOv/MsJQ3
H4Js8w4GIsc6mgBsxkD02x+mn0M/hpMtsK0CGDgQ28OHEDhtqyAqdAflQBxTkCuiKVT+6ipP1oQb
FggPNM1o3VUb5ym2dDpZIw7EbIUR5eM7WAtd4iYr2EVvuwwREhjR9TsV3pSIKax45gRLiwQYlq0G
YHyA71Hr8szJ2f3Dh6dVmedVXXgQc2cPITBcR+mvAd2rmRtxwFEVIcf5FwM5RKS9ZEu2KhxhHY9q
WuavhwC4zy9ghApi6bSAuH7AyfiCotZDiOc7xK0JwDZ04SMYzE3zURgXYRHPP1SoKS1s/2fUZ2KM
4S/rIx1MI5MqcUfixdcxEF1EmVNSG3fgG4kMbinXEV0GZPZlnBPiU1ElI+TolyUzNlzCux8kCE5p
uUD+1myYVxoYjnmn6M+5LWj/e5M9gfOcWktcog1M5igZMsgR+xi7iUQq/3PoZe073MO6+LlMSVeG
gV3ecTLTRMFlX0YRSrCaZJwPvqul5YpuNJSG/9bF3xc88fgYJZnCOreUyUJWXCWPYMscnSrLUup6
krEB+YhWn9FmMWymEAbeNvz+sf5RBGJLaS3HpBBzVfxKrQEdPCNUn7+VMh7FzVygNLIGzcEUPh4M
QtjYTixNmj/sw21ZVXqNzAZ9WFR4I0pU8aMsdnwL9ilrKtQM3ddTl1iE0LZxZUgyfDhfEczET4U6
Ddk2e251sksq2zIWt7Y9KV9EaxRhZe57QdfwdghVjeWi2TSOSmd7YcmOc25k0ulZxu9sPp+QDRKG
dc8mREYkm0g40/LokNVq0t+tqOZt6Ye9MMIh6lLxrM629pCAotLcLMnk2ZqN+wgnJiNWM4+gmkGo
KM0yObTTiu4vBAzPfeWwmb0q7jB3vqzMWitulXGDORq1ApWwcSwGk5GOULZxiVQZo371rlAaOTFH
/+SgxY9crtGAcoK7vbXpq6ENz/cUsFw8DZoAyl/4qRKxJ1c3hlkMPSeZuVxyBGVR+sg19iRpiwye
zypwORJABFz/D0VWFvG5GkNaZb+UfOD3UhHMiTC0aZpnMeHzd9hj3k5s6sWuMRl9vWAkvd9or6QB
yUN7K2haWVAb4bM22I8TVPQmZ9pVyqQtHK1iVhAfE00EDqCAYmT0al6riMRIbdDXrEBAYXcv6VFo
MMJkidafMWk1CAQMAi2azJEFp59O44/m9AHvmb6sknRCU37luf/qsHj7m2qVtaq6AjgqVxjCnI35
UlCuMYgcxZJuz+ozX3k8yH0ltj1gcwqKFVzL6NTvgRpUGOmGUmai5emUp8rRBqtSiePJpbqNQs9s
qx2lor9gVRJIqwZItm2IaOsWLJZpRXy+/91e0GhSz9ZeJCWCVBYHALuZ5DNSmU0+czxI0MATkGWO
8NX9frk6nFINothnkqS3ymGXxFGwJqGOCpPvBXM8i8mWLOrlXNIMQb/yo8UhgnBaqW7kl7bddCgf
UYiRHaDKTbiyVaSfQIKs3deFaNckDF7T0sLY5X2PcTYDhdFOnBo0QV1soEU5TN3zjZ6HNrBn+3P1
25wOeGDqeqVwcTfTZ316NEic3eBqX9PiQ0/BZBhno5c06kUMfp3qVJg/g25TYosFfyuASOtsir4I
qTsv0+G5dRSfWQjgnWhPYJ/T0+wIS9JNZrjnQYP7kUgQLlmcwyvv7g+wDW83JLr4ReR8pFsguQuE
z3KjXXr402EbLgGpEBHmpGrw2rgFzyiDWg05dVxOje6wwC92VnG1tEHGSHzUR5tqLTanaJ2sbLYp
19g7kBg/2I/cowNSJPFrg/OGybB8fzDsTUnFgRAeXb33BlUIPq/YeMeJzZtj4oJU8+QtZcE0EN4z
V7m+zkdS4Dv1bIiIqjv0r0Y5tbZM9awIe45u//g/kzrKZkIoU3AZOYGv8nQo0LPjx28WPv+AGtt7
RiH2E7vlG6drJSsBMMqy5GO6Pk/urOimwCFqAGsveJpv8+8PbskGNsQoA7K52z3JsUz8mfSilt/M
cIBPAfgDuM5fbv9U4Szz7BHyCxtjQszXJ2dcRJho1Py6JPsQJTaHPzwuY2cYQXiotowPU/PGi9Mb
txZy8DOLt9imEs83xoRUfyLRzOXjhlmT5fwL7727QNAdUQN+Ekvk+AS4lUvupkzkkXGLunA4Lbl6
PNAbIqYl83f8voAExNlLgtbBNXw3cyq+z0Grf/m6w/lCYqaZuol6QcpkMKL7fi8dovpwf4VvQ7vV
UmriTYrYnBvStG1LHByRrA33kZTj9uXuzTVBPTithz2Rj5PpYpmYV9TAsajRNgL/GV/LJhgC0SwH
MxgVsrr8snsfTu3xBUk3Y0TF3sxKQGg8NFbmCdMxQR710MR4irK0sNxKv2pf2OesU/NC0giJU7zN
FEFas8BbNW1XYmkni8YieN2Rlz/QC6umHNJX0R93glXP4MEGLac8U/KqNPQq0Pn+UbCId5skXIx9
TEQ8NuxhitAIwteyBzW+aXtHARBhyxFZU/vKslgygoYAWTjzD0mhndZbRwCl4GLhxy14lNDsY0Vc
SCNdh4IeieRDCuBu/tiM4fM3f9m2rVtMT/uFzg0S0ANgM0Lu9TesGZEgiY19JbKgfcxQ11vV/h/3
6DmOOae5HLP73T1N3T9obZbmyhq22xiV2Q1nsLt14S0juVb420Hts8nhlciZjYh8BavQ1BMeJ9bk
gD/q/9myuO5ouUO9tDeRGteru9s/jXhX1sqWyN1deHB5W+/rwb9U6Y1fsgxx2v8DbW8fDBwogP0P
xQw21IfipKck5rDw9chZ1CI6RhXLMv70NQMTtDFsdmj13QIWMEzZJY+krm5cAG6obGoT5SKERboz
Hl6eXrZ68MXb6g/Sm/aYlSLCm/0qmHr9NdNOHYQdpm/FxdXuedlJvCkWP83d1DV4rEFJmc3va8F8
2v4hHhQMe3HGNFtDrVq8AZSzEXLMCMd92kGgW3bPasDHXsP+lgUvf3kyuJb3uURrZCFO86791IcF
cAzY3WU/JdHnupjw3yrkz0SyErXhKomAMMh7iYN4zX6KdJpvKHQFWhntAuKWWZaeePp7px9iMSb7
LuClIN2FTSdN2DnovaMcQlVzvKW5zENYaDIFB+cWNmt4EEJlXNay/3aSSXvRPOAgDPOst/6fg105
83z0DN8AS/RtDk7AEhyzG9hvRVH4FDFTU4MAWHqvVVWkORKYTCh6YVQTPxou5IxFzmxGTtaffSc+
8M945E98TT0HcosKEijBhMvJIZTDWcWeUwrEaLynY7u94rM1NVUUghu6g8Jvk8A2A1B9uHqxAZnK
2EbvqxMgBodY8OQxigBtdlrVLEPQYTUPDiJ+TFdfz6llLycQ0IuSIGZFJ30tLvT+amJzMRiHtBQF
+2wWY2PXRMtpC/P6idwRP08qgw77Pug88oVx1yF/Ckb2cMOLlsvpQHEfpN0GIfOyHba6xS5RAHCo
eGW5r1d79YhuxxGxkSNgA1ls5ruGgKYwLZhw0d//ZuHYm3E4ZE+z2ok9cBvT0jR+SMIgnwe4vMbh
rTLjpGHT3ut1Ye8+eBq8nIjTJwlRbGcKgvSJA1l9k9uZEi74v8hPIah/iBRihNR9LSHk+DCLI3Vy
yBl/5XmCJRhr7VUJHXoJGO/pYnqIkIRK/72mGik/HC1dD//BDSS0EdjTEMPhqNfZrl+WmpTokuJ7
Pzz+rWuSofek0MBFosuk/ZpcdMN2rBC2W/PCy0BOnvkUuG+qCAf7LWAOrLU4YdLKW7/GubaYCor2
zhIcaFDKj+R+2CoKNJWIx67KB0KdmBHlYOLc5FfXRW2qpOllLUz/ZKV2+EmjjkPR/Xe6hNOBfqbo
uJKCckmJdKvoqWHi6ibo3ta0G1mWdxU1wTplK3XK96ichqLF0Fy5fmZ+xo+h3+rnaS/Ivmh35ZQJ
SHkPu8eZw8/w4A8+bx351fHT/iyfWz1RfKwVLX+Pt14c8c8F9P/lVM52GIzTDC6+1ZVUxu+DPAgC
EUq0tTAt7YLwL6qgQNRQuzeAkF3Klw1ATvBs7CpB74Q7XcUdhBfgyVByFCEUZhRFAdGtft4amAWj
wdZ9u/qDqXmKd7SAkrI/DqDr/sO450kxSri7hYK5T7MCgbO2eqDNyaDzUwFuYUaoE3IKARh7WJwG
c5zBO8KFT9S6vExB2TcsmggYPWfDnZF+lCkpiorT9H2gfQ6U8EpsCY7Dd2xiot0QZDCJCoukF+zr
sbDcn3uRy+LqsAFNn/oDfQCErSg06GBuFw/sC4krNLbrxq5I/+4QlvhlfFwPzRFkIJGvFWg7hXoT
72FWKxNg4poSqKC9xcFDBeQ6+iRH6FyzzAUEP8Zxw3hhYGyBTGOczEblgQApmTD8vPUKaedlUqJU
I9iI40ZT+a6kDtvN3afv3eq0/eYseYLV4pCpW5r1mNG0bN2LJL2PR9zvfCex04sjsq4aGkwWZ+uC
8OYxy1NT/Y6sIERHsIPfwVO9yZkPAOZ/Ys2SR7NUUmnBi+REVOUxNokWswUerVXxZMTddOFbouXw
yEAArIv0a7+b/gBdNnvEeDdwRh+fgeUXXH4744J9RZk9+kdtYRFvdh//7Ehm4Tu+Asu7BFWJtvqJ
5N6bz7/pSC5lh1l3UysCXyB94VA6PzqmXQk1rj0PbhWWj9xtNH2S4u02emK989tQ5WquRoSCwSzP
adlbEG9cENUWtlT6Aczqh7D3MKmm5Q4KkbHP/GLxN2mXILba8F0vTwt76qNmXs1I1B5Gc18x0+iW
sON5VUR6RoRTUNUc6dSgTN8k3mY9AGlYcd0n8kDYewryjygfBIfi2HXHgsVXgVmTX7F2828FAiOQ
3pTtEIhr7bVDhZwNDXbWbpytD/8b5mzHOaCAYsLQJUJNeJ8+Aong5b0QO1YTsWKs/pcFbzjVO1vH
Eywg/uKBC1U/+GL8iOz66g1SjbQ5UqgQAb0RJ9ZrNocbeTCQhjmb7xDtMT/MXXGjPlJfiBRSEBLL
iJLZ3MzAlDigkhnl429m1vHJs/swBI1rimy+OWHnNTcyk4NQahdwCJFXNxUY+By2ryvkvlmD/Sd2
S4YIQ4SJJuF0twUawhr9pQLnf2E/ajPr7O6J0rf7bc6gwODcr1uZbRO3Xn8IhbR8q7UMs+z27R5T
gM9dpZ5RtCBqCkQWdmGUDK6XFpGLsqX4A7CWuCcBdkobhzQPgiF8o3erGx0HrbFj9qUBzoAGzCJM
y0MlQERXoeHjGW5FETYk3N3DMCPiSdo8foeukrEO9MR+j3W85HW/dxoXiaNMoum2Kvs/K5dWxsHL
3pXRSSuTkLInNYpZfPLElmcbrqBI+mdi14bHAdhKtieEiMOtpxOCZ7ZE0ml+YQwTyjyOC2UW9/Nz
Pdmb+ij8+toDhN+MZfzl9+gmVPqfXlaYZsJtQ0S71FscVOH7ddqer/uuVywGznJjY4+juBUVEG07
V+vqyQbbvv4BUSzt7RL0Tpx9vMN6HiIZN48jzrt6fC0jbrqxWKmOtgElvaN7VU1ZFjL1EkM9BQpJ
ROMkP9Nyr3tFYeXDifw94P9eye1tdb+njDiMVcdbwofkvpyJt1R+k06XcnirySvIzQm1X5dbliUL
xzwPqI8e2AsLLYPSJDfG48eEj8Npoi7gnj7/hp7s4bMDFCFFzY+OjYnryEcyukHcM6VRuVopTIzh
ynNGDCdqu9W8unxzJkJ4lD47WFgM86e3jOfIyikr2kCQ349BQwNv1X5558YmtI/445EmWIAoJdhM
9NPV0AEBC5/sII2CzDBFgqhpOkDi2HQynGeJkgr2rASdj+JVZehJzHE+rZCyuAP9iXtZW83O1fDu
W2cJQepDXt94TvPNnzO6GxQeHaULRVaaZr9m0Xmnivt+rG5TW5a+h77fiDTYYOSmPUmS3mluYVSy
2kr1MLczHZzxpVSBfyh1gh05X0npC5RAZA7kSxTaEr7oQ/BGsmMxTObb3qFalhkIZpZqhjJh0vyl
NlcNmEn5vX6FfF79bZ9Ae/OtL2bZa6YuI3w6jqKhQw76uxpc78tw+jvk8xT7wwBTfln/KRDF2dp+
IWd1xmcMk3Pxh9JJDAzicTnM5mXzjZ3/6L+iJPCHc/dSjgqQZLCde12CyBopJy7tjG/OAwhIfGnp
ZL9NbStDkdJj1iWWCB/nPxaLFSPG1/rPi8b23Nf4umKdluk+k+VITf3lN/5y+pry6YUdBqZgj07n
3Cw7DY+og2m8/D8p4DCVy1LdDLjW3knK0ve+V6fKU6p1rLXc/N4Mpn8ghX7LTDhNNYukPsyl5VM/
FgVdkGCG9s+eeJ6ID+FebFQrzTt1D/t3yyyW7dnJV1JFsUaY/GzB8MhktjaaMDmqwREFynqTNXj9
s6BM+P6t60ljKSRROr71Tldl5gZbqSalBWC0S8gh00SSGzHo39uSEtmRcx6d+Tlw4kxTOmhvrml3
AuScvoXCaOnGvfDSoL0GlTid0KFhpzKxXoXNaGhadGsjg0KDX9ErGSYLzHAXl6UjNu6oWkynIvn0
OvoG74c/HKXwgOhrcLxfqwwv1112tVd1BPnt888bUtPQ3PiD0hdxKEKXCJhBj2hg7i6YIDQMzp2U
TCugIEvCrsiY6eQ/jawWETp9NTLPiJwEfNTHHOFmiSYkgIZyWQViLi5RjpsIjsv01Vlpm5ONZMRA
FPGiWqdKrxGnv73rknYNjHxpddmn7EkofmKP0E/N/X856OMGTJnX3K6ta4+Nd8x8DTuReNcmCaUe
+V6UV5As9hG950vH/9ytpzy9exDOs/7hRC3TWhi9RLpxaYaivT5Q9SNGzZmmjs59Ti/hkrykovP5
R6P0mQaorSy9WhChskn8mRPmoeSG/xFDV9b4kHr5s2945cFO889cY9Pjf8Oc1Y0rmFPmVoV4M15m
1H4AjLh2p3wgPnFrCNH/ejunuHR7iMDNyhW/E1oTZ0pDL4yaPlyerbGPcU9qCYzQMMTqzvNFxBsJ
elVHczGqd4GNo1iMKQXKLgb6ImntCfXCURV8AnGXr0WoBHF2TkNcAXzFv5/yRr8DdwMukwe7iQu3
v7me5liN0n53kA6d1Ixkvp0A78ghkQn4DuR8+yjbbIcF4kLv1+A8JwWWMTT6LfBuixt9u6TBOqSz
fYJVMHUc/bc84Mms/u4T/WuDIFaY4e+s5p3Bry/5iRLoQJXRTimkc8f6gpdFK9rPSax/z9XiqWpq
RbCi6g3LtbVlOTBC17ehezNGk6t2BA/vD1NTnAuonywqGeVE+DbBaCz520wXjXu43KEdF/YCMowR
xU5KjPwSKQboLiwg9XGUMqbg9Y3npWoX0MTZX/qL4QNLOoPgkF14guX0+cjyDvfjlABsCgjxTp7b
AQyhZpPO7GfjY6gF4wNKu1oRy9lBB2E8tuAzy+G463s+yFsiB+i7jIfQ/4bB2e1QtmezAIh1dFdE
pxkh7valzl2EE9cjTq/FBJUn0zi923EGO23Gd9f/H6arO5Oh20+DTvt03tyQbEIur+HTPllz5eD/
KXaKi7mBD7kxECL/Y2ldNYtm9TIJRgQNSYkDfhUh1b36o5UTemSDTUFdild3lfSnyzpewOHTOY5R
k9guDSfARNdxa7Ct6GsJtndHNGi1HFaTwruLCVGXHmBTTStGDOQrafLqMx56GdrqhBp7nAJg79XQ
7NIVz59722rTCEHsU3KyXdb4QYuB7tUEUPNSaq9z8WFQ3sB3mO5Cmocw2mbTVhd+CQZRSjjdDdnn
nge9nr2xZHS3HY8a3GDWAnB1tQGcH/VazIhMpJeEr++EOmKiPvxRUII35uiwrDem9PgqEXzP5A/Z
DkUlgUoDYHnATs8sD2mnob1kDpwMAcZMfCSNIj8Iitp+qrtxvwR8Iz3A6UW4BnZFUnJwPYw1/JBh
kaSW89/GOzJV4moP+rA7Q8cwrLDNam9ZfJSi082V529HBdU4HF1szXL23kCgkN7iPmdzAzKsYQKl
2oT8xk5bE4X0tYu4gaVeg313Am2l7gxZFTzfK7DZPEsh3c3GojpFFqPP1PbQojtFkmSWJXdzA2rm
jBgm5+Ie2TBvMkRAnLtysOOZWYw79MvCBG2YibYVF9FkwOhH7Yf08UvvfFoBOjssTlczUwWc+eUj
tjciTRW7Y1cwv3qDu4lu2tWTXND2VhoyjmbdVzDbdiaLGDQ1INBu503WzT5QbMc0qIja1jH2Md/k
DebCuCV6XuO8M/MFlyGze3e1mdmTnFhXUsyFs4LQ/TZ+aITdmXP5j3kfX5ccaKaqF42ixWqTOG2t
6wgAadJ/DcNKEZhVHMwFVu6MIM5fN3BjJM0tEOpdJmmZqW2lEMlNpzyjcZzhBm2DRhIj0Loo5zc9
/FRRB5NqqK6QrNqYAusJCHudIFWCj2R1Uk+X6QwaAQLWd9Hwrn9NKocT0zGUrBCyvmRV7apNgVDT
0hiai0tAGb4cKUVs/7x+fbpPC4MoJQM+U9DYEcAU5rvVi1LUSvkJFM5tFCEG6zslxAhIkaWOFrIS
MNDU/iDBbsef3OFyGjnRt62Ila0mtem+ZxvxazlburxjzuneSJYNMtkn8VwqnBXOP8Fee9ckYOk3
be4fY1ck4jFsAGS1crSV9yn654KUJOeE8kRJFlHg9aCDEEwPDqVYLq8pbnV138JUK8I4sp2yXjRn
+kA/KJTyrHd5/gM6R270lk8k+eQDKyrtOV1p1MWCIu7yZqruITFMciu0EacqDgQiEwB1UdXfL56J
fZ+qgmYpMOFGAakwzf8FRsBjdmfUa3ZA53l3XUekD5kDHogp/95CQC9Tfr6QdefDFCl8l5HqDo+f
drtkCIkMV5J6VZ1Ir82wnPr223LS5/ykS9726KvT/zeLxnbFiaGPrTdsGBcuTfukw+x5qW03+31Q
Xq9VM9S/iWEkI0KZsNHXhId0YK/xGJYWqnWjuHGs+7TlcmKScBlp3TRjeZnaZwfzI7YnQOht1PMn
YU/XqPxAFHPRpzvwdLDv0JWjf1m8PD61rR85E4ta8OaBvEU5TSGU7IGMJ2AnWRubD0skMM/tctKj
txrhmCjsZ43xod0965P14O4dIF4ZVz/8hCXIw+sROuKwSVtBIFHhS3UUatwlGp2wLwpMDSQt9HKg
vSZCZjEwQx+ndbxay6Ml6K8WbsOWZTRERz51LnrDUSK/UBP0NHAK+5rzlYLd+SpkS7Ijq+TYMbDt
IP+7iID9gjeh0dbIdx9UZxThWVx1MjT872RMOUkOz9WmAJgK438FnqV9IltG3AFt019C/OqBhowz
osKi9O8ITxxQG1y4AjW2iKn3WSVKRT+zFxQb5cGRH+webuy50n5TRULG2ccXHVOA55sjqOuo8nqD
y6d2V9GYWPMphu3BN6cxyuNcQX/Hvd9lRm4X+FAVhUY3hUFpYY3nWoyCRTZBKaPg/Eg4nXZApXPK
NywJ3Xk9jQTVnisIhE/POroKRVo8sr8A3l8EUHeM++NgRB8SAyOuyOzlB9qVEoWc/yehINofsA7E
Xrkj4Yp+1hHuygdujwSfI7uayFnN1WbWAd6wUSP/hOdUHs19FEPKGajRD1FatEEMGubXfuz/tJxU
ZjE27VxdgdnVEwE6pwtMLva2205IC3rhAt9VXN60T48otn7F3x2umrGlhZ/mikL8E3OmssCn6fam
GzD0Pl34WM+G2Bo9/eThs6GLmj8bg97yTqBRy5iqoALJfZLywKtm1jxdlO0BEqxPtu3I1baQtcSF
LwRbrwqXQeotKBu3kQKCTo8H2c8cPKfKoTNu2f7qZ7wd2yq/m6Qm/vr0KWllZGRu4VzyJBhlP6Rh
5oWDDyi6QewNpKMHVwnGpNcK0gXqniTunveTR4SXSgV468j6qL9m8Y+dvsIVl91I49BIkyNNAJ3h
7LrXU6IAx3AeAqhlxIGfpp8Yd6ts1WsBSs7JnoqJ1ecvSyFHLPAV/a3/OhK/xNadIJDKoR0XMJCS
NpARo7aWo7R4cAOGLz5H6bIZI3vH68H6zPhYY4YivJfmKmYYGs3/fhbOZDAp7J35zh3nplT4LPSt
E36/sXB4CPwQ32F/ysRsavgJ4Xvngxzu+D33c21Z2qwtoV+25CWw7wr7100o0eA8w44lgd5PzPlC
DJK8YS5nbbRyj+OWJQN4L5Al8dZMDezDI1MH9o6QQIWBpvRDgErmmf2SBqUL4mG5JgjQt8Da9Jlg
TW5pLnojN8XbS/BOtmSzkIcuoEowebbjhlopfp4N1ojRP7xzAlMcYHMPiFWEaTCtbGUuqbASWP8r
7FsRvfAq7fAi2oDALdxkR9p2AsJjF/3pHoUTF22Ctrj3rjkc+A5/FAUkCCCDqE6qIgBF9mumi3ha
B/2AFBxW7mrCJOqRw/TZqWyhu/VbhafeVzziRgYvz/WqRPk61IWps1Qvj1CYr9BFZ5v+Bc1G0o03
KCsnmr+FImg0dT4Zs9QdArNw+NWqSWV5rxJRRZIYl6imru+qwv7FgmgVXXYbgAIhNtD/F0RWaVPq
LiztMrle+t24egJ6IuNiJxq7Q4M6tRcVJ4WPHHYB062DOhKzFeMo81gkMdlI2CiysxJiUUet17Nt
gSbDVrXYWoUmZF4ezzMWQxU1Zenl3pGJEKLoYWVztof2IBMEARq0bxclpVs2oQFe0yq8BbiZ+0c7
iSjkLUpBmJzpkiuqrlxzh/X0XkUYf3TB+2SQbeUW7PnRDHXl5YMuCG8Xy4vy7FejMSK8ZT0qP3ZA
AkkmHiOgivPID09hYrcbfMA48bcEwrjLhaDCGfscOmtDDOm4nJYbWEKT1IoIGK2pkah2cbj9WtT1
2sIt1cx+tgi3Xw6aAL6/QRCTUzURwJdn/ZlwTiGV4eQikFpanr3YEadMF0bp5LK+PkfN62s5+5iB
SaHts1CahpKCPh3oFICO23SN7JXWEsx2FdBrDeDpsinb6PMtYHTi6/WHoL9LxnKJQvTXqqaTFqrl
jl/lwP5QEpMwPt1lxC8jq/bpQu9xn3j3j9FZy3G6qayUZCUdWJ8lyiCDbf6RBnGQSxIYmwX3t7Po
kdGGSvUnWXJmUVkC2f6GAEk7FKNtvOqpyEeYRjAIRuD+Plrc8RegQd5AUmYZadhJq/dP6Mg3jOdh
QCv6bBaOTQ6S1R3iaT/aa5G1FH5iX5o41TeEcxBUARAx7Jq8FtGoDcRGi2FiZi4pd7lh/Xn3Yzz1
+bH1xcFhvHeUERg9VvbooOpCa4KtF/vv/KwZiW6mlTJK5ciJU9KKLTEQ43+quikYqa/pZVDZIAuP
GLofIrPnydcI8i8/PS00DPm1na0DtMShza6J4+6jT+iR5Nr6xDYJp6QHI7G6PWxUyRBFci5gG2J3
ksSoT+IF+WQZoTfnj05CUFSa++RTGRm1Sq8zGzg7q+u9uDU5uefsTf5ZPIOJk7lAJZDRC7Jv96Jy
UffBm78oe+7TpnIXvZWP33PQC8IpzYxblGeZkV/NNQKzvdSTB5/VWNdXo5JvC+jxewh2NR3qFy71
QALa5Y/YYVJfqZv/USpFQuHHv8dpZQ7jAL7BKqMfqJa3ATgs5nIptULczjVYTtsKFJBylUuuwiFZ
oH5fHzQrgy+KsV0zPCoFgiLlflW5mwZLhruSwLkslgJu5/0/6mGYyLOpxJxp64riIjkjnof3w2Kt
XxPBwAS9rWJB/H/3M3DyUGhwG7fqWjatCsFU4evt4/0w/kR2kCWwLEPA/7ZOF4HqP8GAftqPneqw
QtwzryEL5YJh+0XD908LTolUvV/M8KanLFRY8eZ50lHx2RJogMefhHobAFDTeNAncch9lISzDryh
iXwfpniNz8ycHMl9nIfFBH4AsPYRL/1L7szpKZSdZVGo9TJBNnvuf58zG9LSPzvwhI/lvvGq63th
eGUkR2a7C8r7eAv7ptU6EGzf5D8Stbc2L/X2sNUbzqsHc2Mt/MXCz88lEHHAbTOhA9zJGIZB16tX
rYVxhezlbxuUiubEbIa+XHDsez77Is2z1c2xPHxHGp5InKDHynekrs/Qq28nl+tu3skVhwcueq2c
mP9pBkPM1OMDQmq2TduZVVdyzTBm8uF/L+sLLUdwnPvqCVDDIeh8IHJ0VkMbLW08WU44S23b77FW
S5hePA8cBGPjTTY7PVPvPamw8o+kBnIG3SHGP7XUZAu6b4uak4tSre3+T33pThZK3/oi2680JoNo
uAF4mIdAlcmDDaKfIbZfBoiwrCj9gKhcLDy0M4b50h+c4xQE3+jKV1RpnihmhvxvadBeX/t6CzBK
0XqqWHl0vat/qXiWdG7ZoBc3IO60v6UC3gLSXucbqliBSoPKD18eJi1WyOxVzhoIBXc0My11zcZ2
zVLmkqcj/jG4evcLJEM5PTTBga7qmLRnn9qKcSBZcwGMOd4C7gZ+AqZxftBIYZSlBIAtPEZ48K43
W2+/ooQKe0Tj8vq8Fa3BuvnsUKap+he2IgEHTNVIfvwdx5zkaL/KRQvsKofYbPNDFLX4JrF1GXgO
bDE3CcxSxIh447IM1Os30U+T3OFOMdMjb9Ls6z/3jWVrBXKqmVFUVCDIMntGhjuYl1gr8bRS6Brf
gfFihXsfM3s/gk7SD8d47ZZCJ54ev0oH6fmiUp6WEnNpYKxbFZnIDgQsXqTR8ePvf4JK2C7uOT38
A96AdUhhaJUAIVqvs641ypmi2v8du1ZIPNUQXxvdxWfsyHGdFVwkR6vTSnlRfgQDAudTIV8vwvoK
XhHbjLljBpIL8rtU7w4P8FfkMZBDrvM+ehJl3+50MO8hds+nsOB4V1bj978JJhJwI4mraZ4w4oEm
ktbRCZZ/b8KRw+/DRxzreH5d0JUmbNoG93Tmfm91o16Wo3glGv12qlPlnbLzu2trZNjVQkHADqIi
qSloGAAj84GzweJo7rZBq11MuXGyr0N+b1nhsrzYm0atMT68dDhpvJM4nzU3grsWvZP3o3te+Pjg
vSs1lO4ZV6qnlXD+7VWH1j+w0ZAdaoDjHObneYjVMCHS7iXhRnyB+Z94dY75J67by5W4LGUpiARt
vadmvB0d1bRCvCyrXdplubWn3zuZuxdAJYHqnJD8jKhWooQqyJu8zQT9EP0wXn4vhBcRzxrBycAM
vlkmMlk+PgJFm7+lSKZdGxDkUyE8RfXV2MUHiXYnH4yXPm04MC2D3wzJW0R1PataQU0d1YYvM0Hy
U0WkfA2tGl6OPXWV+4I/IBiRhwiO/vH9OsRo6IUY7vSRyiJD4fd7mzRc+Srl1zbHIaIdc6Jllhiq
vbWKLIrjyv+hU++pthyi0+b1z727ujLdxFProndLU4mVwjO1pE2LZ+A1fn10JbloDESxD+H9ae1u
b1XN8mCSHsDDs5t7oXSAa5Q4bKhzWv6tkbaYu7HRzLOzm4BLsqaWdf11k9fwNiHdt+t8I7weVrO8
UA+ZaWKi7H5zHSdEcA6drtJAO1cc3Y73UM/UAtCDg43rSKlnOh4wUFoVj0KHKq9XtOqhtUJtG6ld
QuPGDG2q0pSqLNHX9x7ew17orGhhYCAZ/dGKbKQvm4Z2tbvlmAZFvMXMZNGHa8ZthM4tB1pal/Hg
J0XQU6FyWWzeRoeoq9ar2oIKCkrSahSk8aTKopdkp1dCM0gtWBz/+OgXcYZTRV6xQ6s78dVA0+Lj
P/Zp1MP/XrIQDvbiLtUEqtFm70cAOpMr8pHTlPQW4z3/YH4paqI1ULBIHo1YcVaF3djPOvXYEgYS
V52QffKEZKP/IfQVvAPuguYv5dr1RAb+SchpVwlh3Q68A/k6R00ov58n6UQo3kzQ4/pKJOkuyrCj
XKvHa/yW+WlnvmOgvLdxQECkmKF5QLi8XihlZDBwDdfv8EYFqAj6w5DGwm3wX4Sk7G0q4l3QuEfI
VsG+EmcPuKfUl90KigRDsv5nZ3VyPcryf463Pd2I14tIlWWTOHJoGmLA5OwCtiLtliJIH0r8PdRQ
w9cB1lMGpemuFA1JeQnjWwEHj4O2ksbER1sdbcA3ZPy/tDaUm+XHsQpZ3ihZzZQ/1gYFh6WeDTbi
4MqAyMo0sQldxU1/DPZOwfNo34ZjujyVPkTnQ3Nr6ZfO0aQ8CrF94FT6bko8n9o3WLsisH0MR8On
wuiQsTM0TBWjb6hAxKYmp71WTdkAFG56QR6oOvL4ePp5VQaCOqTMyOBfD7RIogAyKOiFlI2XXKDu
FPfa3eEAkD5flzCtAti5iwMxn9UE4hTY7Tc2EWP+UQFgUlgkvd15hrh6gNHPkEVTvge8zYglFfTs
e95zVQhelxwrYrXlCoeov5vxYgQgnOYDit6a0gBnOQVRz+VtpSQAN513THo226wC9hdvcB5yYqU1
MCuryS8N7lJEK0TmtWWQVoV2MPEPtdcEcQXuT57S5LJHSE4Hq8fUByHzDIwnTTJuhNWfgx/3Muts
cGvoDw7AlnhApQWmSsXRr1YO0mivD+WmSTBhrqsIEVDM4Q30qHYXCQB9b9khNurinBbyCtmNcN2B
s9aFVDB/G+d4ROccK4WeZ3FEGv+CqhQ2nel2x+4jzX9I7ehndj5Z+uigRx32DE+dP0yX+bLlGvpr
9Wtig9xvIIN7ilXKlf3Qw+xnEHfFrPeP0Ns4cDv/VFb7QCEgkszns/JMHndnq+H989RraMWHLQM2
Jmy/4MKLWIr6QEcUnXqTdLXy/epiD8N59OBkv5HMQ0HpXqRG8bLDBMcxd8VHqS2Xbp4ZwHy3FuxU
2TwkPcoalAUx2NJFZo0tBV0GeZt6B8hVpiQkaIkk88wgwMbiyEHPMgqXQc2QEbl43BEWAvGXkfps
d3+EfwBCV1qh8K6SA/t8TcSOp9gufg+GbxZOR38Sci5ValAqquW5iVLdXQZoEKUEzr3V8IU/b02o
q+xl80eBK9yMhHaPLGavJ6kgqvueGlRlO2INgVLdko4xGA6jUDb/BbYSVAYs4ebZzIB1iZQmFYzd
EqE0Iq4gd2ap3vsq+4T2DBPI2Sn+ZAeKvhBFjS3iKvRnAKzt1lYrM8BvFiZXLssAGFbD2GsUqLhM
yjqgmGtyMB5+BPRnDZnUu+wo5R1aOSrZ9d+UsT6vn/rkhcHFyEPEk7ev4eF/rh8dYI0iOVATmf34
mL5EqSbSc69unxJoImH5GKMTM2zX+XaXSG4v7BNQiUFmRmqhtVBZXWaTWe3BMfDlqLRsqNV10O1P
k0Iz9CAVcT3AELlEPmozFlEAud2YdH/iKjXf0HUU/WvYQ6ZPUCttTXl4KyEHoTRMRUN3J0pI+0Vz
dmCZTo7/EI3GXSzbXV8OQDl+Is1rDZYN9HYSk/v23YltEutjf2CMczFrpk4bdkfQD64N6sI45Ox7
huPH+CYhiMyZWwC86kIWQYG8KTl+hdtYdKp68hBNmsyvWps6Zvlf3i39nHV88dvp3XEUiXdm5QVX
zOsMMoF4/o6l+UNi1JN7ikqNwFyCgZmjp66SiI53a6h8XVzQTl/p/wo7GMydKOfOfo9EBqkGzNQ/
tbopENMTVAXK9y8insfS7EawHWVTjOgKKJGADK8JzNxZGP9dnv8/17hShIdF+pwz39sDb6RBK2aK
0iVgBO1LEha1QpE0yTgZ6uq6VRO/hbuKjx6QTJ9rkil5wFVkB299tCp1wUvk7CMr5QbuzA74hr94
aL4Bb+MlVXhTRxUxN1qw3Ns5/caXBosyQObEO/4vk5woD5Z9AXpXbPX72EAYO/91pixzPUHaUj6C
gGdRYXEz6NE18Fwwp0+9Ftw6ZTDG5/MOXNbz8SEAV13cJNLXD6EOCFaps5pRld8mp5dv3KbBb4I1
zwCmJSiDSpenai5GrugJVdzM97OmcJuLyTAvw//9G+CZF1qByTCiQphKxzjnMaJ1mrYYmzzEyQvz
vvjRmTtXkATAFk0QCxYtjHeRx6OpFnBvF/1gKZjjG+rbojK1IDTUPgxpOlZQkkBeVQobu9NCNnxq
AQ1UY0T7g02BGiTviOGopCV1u+pXQ7XmwUJfP6zgxGzIth1vE7r3E7C83OZnlspS/JbFmVHTpGsU
5fCnfx2Vd0HQRDkE4O3heB+7bdsiHGkl7ENnT1gStDGei8TpcXKvvZBo/9WDSkGPZ3iMUPuFIGs6
2oAbb5DFm3qZKxpaJmj/iQdHKnx9+SsYBUPSQuHjv6sPL8Aheq8ihouQhoHmjtW6R3q0FeoGXtUJ
dAgiM9fYMeppkr7Nq8EFaJpQ83TJt7Am+y9oX8UuH4LjCW8TcQdOT9jV0OJaFOByj5dLvk9LWewN
OOtABekuzUcqz8N83r5v2zBR7fuCo7x4rUDcAsMuZ8o17CL3Q+/fB18Cz9cGI6cmsTDBy8FlRC+R
qdg0L+S72GlqKQs9Yq/4YjUftpMzc4e0A2jmM4OM3ZFMfKL5Fi7o3O4VMlWcYsHkAcGhHdS9n9I4
/f/jq5IstmlTQeixkXYlWIPoxMjr508hHexOKZMwbsN+Vf8o44nQvG6ejMDY8SeCdeDIAeYLW2VQ
Zcht2t8XmJrSjHost0JvfNBaJfAnirNcX3njtuvKHI9qq7fxEoRIWPD3ikTE9sNAet6pTlhEpkGF
njPe3K2vjNXuwWPMWmXXOYE8zlFyMh+nTbUXkFePgB47dAq8XR75Tb+rJsSLg23Dr3qbq94c2HX9
tM/S+t/N0+IxUI8ooVhpK4/r2C8HpdKeTMUinzTzP4dWP+NSkzbK7ETuklrOHQxPjWB/ZDK9Z5eS
JIysAj2r3fYicuG5G7YfUoIXGetBponewj1vYbFbyygOvqhU2tdHzK/uGAbqThfU+lDUr6V1CqKs
Dx0UszaPAqcfx4V+sZcajQIwOw5RtZdtdt7nTpYF4bILoi9mINI2MTnntLhnmyVMnwi0/pXpVyUC
AReBpclNKC9acQumfuoO4IG+b1xAK/aAh9o0c1GYFBpheztXzaijMIF1s5HCseJkn9D1ZzOYIyxh
L4DYKFn7FbWGbhuYCN2rs0l8eeCp62O1DFEucXS+mksE+4qkiDv7oKAu0CqYdVmXftxq6Fat9Rq1
SNKiZ7hDW7df0PflXXFk/GlwQvofE/tz2PmnPnEqkcxDNkI2phhgy9B5EIZwjJBQ1pksV1wOiKQJ
Md2FiZo0JdB3DmUOArsrDuiD55iup27Bc7niNjdziCU6RGRMlcWXy5BDWD8OvNndkI6nifpmIMpK
BbldtFb4ieF9+IZE3EXlG76mCY4sZbj382D0gFeew8TzNYGLHdMpMlk0/NAxKBBfeqUXDAWoanNK
Rc0iu4kAIF3c1xQ39lpNDfX3C4aPYBDFCJFid0x/MIMN5l0P/MlUVHrD8UGT0Mb1UwLoQMnSBFzx
Ywc153h1MHgfeJMRNQle/Qkccwb0KGo6gz9rPmm8oUFp3eDAX8J/9f9k4Bnbyf01MldsvrZ2pRWD
HH9XTd4x/92t88cXrCS6zkpifMibMNb7ZYRd8DpculwbC+yBkJfFaaQXAilypFTha51bdmZ6w3eR
YXOODEAB3i+YYiUoS8MvYvC0ImVrqED3L9CsYLkb0sL8g756WwKjAg5GibnT+wRns/qvMGpLtJ/P
eiUA7YzLf8sgjfE7fTMThACEb4YgMZwzbDGKBRglFH/dQspV+UMHiC6YfMB4zyl6zBOUHY5yQPQU
kR14peRsh3TrtBUJhgCY897oi4NbRncp0LFtf9VmnvGNjh2g4uexhjM8fIcZfodHO07Z/o13RGfX
7IgJTYUIaKYTU7ghnlD4AgHOtxM0Fsu70F4N773KO16mC//cfjoLk/bQizOtahguQ8PafxI+u4Ys
cmufZ4Pe1rL6bHNrINciDF5/Yw4KKEHZ4L9+Yhe+GGgn7sfjSv6vR9jwEpUWKOBpRpv8TQWQ3vR/
i3Ey0eh6qdLgrtBtPHGPXwu/DTktl4BAzcvg4SWePBUUvaKQ4aldP7r+8feMu+vr7NP04DF9XDB1
G6y+ymy428scbDuFRvCuvhwcYpStRzWYhDhFGiisJjEM9UhEu8emLFbFE+Z0cTYyLCawIl0xvxrF
g3l7Q3DnIbnOmlbfo5GLVMezLCzicWWdAWmuNYWXOd6AGoBbMYvjApOQQdr7kxIn/1ZjpEuEaYYt
KvDPAcdVvKvg87COlSx+Twq2CEqtI1Iz87CreDCKHGQ3H1Gnke1gG61jx/HU/qNZRtin5RDgFMgK
p7ItlHz3EqJn04K3gL6LtCGEeGEVmSrSfeybSAZuPGRNSgzn3i7oM1+byl9uetUkBxGYug2gWMaJ
c4XSPYU46X2c3lqXFr/zKJ/mcqqVwPjVQH8GermlGUbxmCUMDe1WWwVPsVxqkUgey7sut3KolKJv
+6cyIUhI0p9xfzp0xNQqygMDKmTQn1qpv6w8x/lxuAmHsg8C64Onyj3eF7taen3r8ppE7KqggRFo
2G1ka0kek8lMq3hM0deAHaB/XTctl1JjUFYM4UJ8ucvaRffVPRtUeoEpAYR+JIRrQ/dgzDkUsIFk
cu2kIrwRBkxRKQzcXqxN9y29dqEaY1HbfACMlZim3bTSpoNM3PdCPxV57uDF6qoYYAsd/oz742lR
HOs5NtxmZYCrWeM7qMWswpCFuMjnteCstb3U1D+yTmBhC+DIrAmlfddil4vgv/CFURrPipj60pOf
tY1jP8mI7w2q04u6hoWDFGa1dvzLN7kx3VdEh3AC3XTc0QT83m9KY9KdMSWNcKNTkNKtip8SRVgg
DIfXZjsoW2/0NF9eRtTTWjuW+xQ78zMTr5kblT/eiyXxkeD6BJ6yZxGRoEMDlQHppkU/V6KFNr7H
YeU29WKvtsN+CbrJM1HIMLJq3ZJGRFD93mIikBjkfF6EtIb18LrvBLvKIGhdzM4lrTo2gpQVbQwS
qmS6VOR3bQTESm0mY7UOWvkgmiuMHYxMqSQACM+T0j/GoMpBGT633D+qNh2e0DBBYSzO90WzrRkE
YqfHXUOo9iPZ9Uz5OAsbGCpMm3YO4cB4vcpUWA8+UaQ+kbuvJqpQ5exzRAov55eMPXRZKNAREndH
N7klrBTjREES12LiBfDn4lzqzJ1M24SnRh5kPFtOOWlTLoRRa8hJP04swyH3iS0nAdLE7L/wm/ui
+uyByLOfng2vlGrQVMh6V0hkUh28yVQ3kdEe+phFGR3IH717TI9S7fbwzl0X5morXe/HxyuB+Uq0
Zn+01nkmcPO0hOc+FXlOeSKZzJZhieGeQH96lvxg27IqmBtAB7uz4eaDFZ6FWjLmWty6OcDsgAAs
5awQTalHqWnlYjiSwuU7QJwR2ww3+9BlXE7e8tz5wWpnWFFXHLQThE/WlxVeHSeCRszikj/ciXnG
3BvZIm4NB3TcMXSOcNb5WCQxrDXFbN9cbz7nYtZUZ+sBrkFobHcYybKr0QQPkWJDyfWv2Qbbye0i
9Brf5aVvUhgaFqph60WyJSFWyFoP1m+UTUNa/xfB2cFzoRLa5kD/a3Gw0TWztkPNWwfukucWgfHe
anfDYyXAn8O+yuIwCWDjh0KHBE5Xi8fe84CkGyZbbOIscWRrl8M/aOns3VIEjaznsR6GB9NEtCim
L6tmpcOHwz81Hf0IBIcly72iJFrgyLt72ra8jg2ML92C7vO9gcQKs/1F9qcoV7npHFlAIiNEYs49
Z8b1J75JrfWI2igu1T+M3py66w57m6dvJ2GXsZSUAkgyZqmtYBkxq20xrDvSfkIySJagZrEZL3Sn
EE8674KyboxOPuWAIQixXwEJWLNaQu015EWzlJh0mXDuaiC/xf423a2lH4C+PA0NLf3oV3SWK7Fl
J7sBSYIHavc0kdEAZUHQjPOMjlaxafIIMCbgI6EqhDX9WF9WeNoe1igPySGOP7cZjFWxGeWixjfA
RwSuxz5iA3uzRpF7CpEnHpXxvm2gO9Udg1k232bDUmH5Z5knodqcBqRNJg+CYuo/PkgQvgdEnlev
JiXdhyrlPvCGISrlG2Az0V1vB6mmIh21Hkn+SrmPQitJwvniZ6ZnU6MGcYiLXYq1/fE0FRaAER0Q
9rL7sHyXf6im7CnjB/T3XNYZTtJ+vDj9Yk103fquvxbqj31dP5q/WPL2Kq/P4mNpNeU38oeUgAzL
sQeBj8PJ3FQ8R3tsxR+P4+xGCt+FfsApvozl/rjsqC9YqRVChl7j5bARJ4HKwpw9B79l1QVbLGeN
0ZLoNE7zKvg222d/Pyr+ZCMv1kPCCD2GpkjMJb+2SFZhxxw1XdOyGmU2LEjtP1xPGCHhZoAWsiWg
bf6D76dc0q+6k8H9AnEbKcLADM7Rndr2mrBbFwPyKRUqOSVpNBm6qgVdElM/VNgritSEqhZrIp6w
NZfrIRzvQM5694VyE1hRbFMgG42EYv1FTYFNH8sgg435Ti5btUmNI/hRL5Dj0NvdbBz/C9A+ZR4e
hzYk0BsZeYdO+a8fNvzJoy6fWzMrL1Sy/rgULRYMjlVQrGSScyyOz6H+LP1qUrw5FwHs6JRBsile
McQRpln+n6S+I2bXSBP5I9uc/X5hE5JFrXGn1r9fnSS9PlHXOSv1pf1I0HOMWEtfeLPJZA2Uq4NI
mDdG31Eznm3C3XzFYPw+aJU/PZaURybpPmY1XomNArtsQ1PzQ+tMVPhTDw2tjH7nuOZDYrT5eQrU
qL6ahEjq9rXJ5aBkOfVbrb9R3tmeNRGnxHdSKcRaZArzUpWymsUcgyDoXJpX1y9zSS0vtZpUL1zd
UcA76BqftNY+d/yngB/eir6Ww3ofPJ0yMliVVKHyOv6N/VYPF0FpQAX76DNVuwCxE96XuepO9u7b
xq6k1vJxHFQqnEiDE1HN13N9ATeDVExzceg61URF/ZbSr5jPUX1Z6zTF8CFXILmh1/LToLBoSSGo
mpCSlJwTjuuoDT7v87C8XrZZi1r/IfBh9ZFj0W9DBvuzYIDRnmNdy/f/Zm8kWmlheropg4ZJ3zPI
WapFTndqHSyeyez484Gg7QDVB4hE90ZysIgnykZYW9otKvNMtsxQcG2rpJxRh5IQBKNibX418utp
i5ZspShmegSbDCIntqCOhDVdvodtH9CjO2mvikVMWEoDsQJgMbMDqLjBEhlGf9RrHSS90fsU3gQg
N0GyhiwVFp7oCjiEc7jo7xHEAlPyEOCpF4C1+FrTCpO+OXglhWH5TGOD10TxG13Wii36dUWvELvV
ys9C1shmucQw9CSRjG/Zw3LXh20mn8Vm+Qkym7rcG4n12eWIVC/wz3bvJyFPwYqsxVEpR8P5NncH
hfwNl5gUd9tjy39H2haPeyMCF9azYgBa31DfvwCgwB9S87AP9cEt+qUE18FodwQPLDK1xBzVsJ1/
gxPkb3DsHbPbWFTbC0SaeUY5HN2BxYabDIleTgln+u3/CQqoiTl59hS/Wf4x40YMpZR3UY2y4NFx
xQD1Dmp3KnucBlxbIoc6yRqG+PswviR0LojydiOuC3Zgo46Sz3F7eMDFgr6P7VVCugja7xMjkmAB
zXX1S2IuuRWp7i0GiB9LMjiZfR2EdUnAW53MkoSx8DAiDHAjyfosQ3TCgnKxXUwQXP8h6b53y4uI
wvye66BWRVKikmvbtUfkQJ+DzR4RD0/CCwxzIinw9m4P2E8lxOaiCbQqPexMXbX+aPqIG5L9LrkG
4W8yiJaUberonwf1GPnYnNLby+ukvOYcEcYI3f6GX51ZQzjFZkfAgNxMXhhpW5+FLjwsaa9Osipo
3AqaOBwZ9vYzIDjy1oMVFF8bKTZepsePivfKoe6iVJce009VQgvcIEcYMWsj0aojIyALZL1eKuF1
wgCX1QYAVLAVey/dgkWO0GtcEl245j934AQcwUjzA4AMPEDrRIe1QZbv9z4Jl4DZ7oGzWf5bJPI/
QwhO5KjAmJfJuPj9Up+8QMsm3BLXQslzMI7X2rVOW6k8SZpGp2MPVZItMpURZ5tacOnvihupr3Gp
Aov4Qlz2NhpL1kSSlHPd0EcdmK6JOd4GqnITbwKAr0MJMqOnOnRtjVAoOBUhv4JSrcqWu1a6IPlv
eonrniMbOigt7XLOpXVCKivm9uEHKCH6+vb6Uqqcp2WJ7XAo+3x3katqo/itHslIBREB0DGLcxqy
b+6onZMtuy+8WFbXf0iHT3FAgi6vwosQMVSJyKBkD/dBMPkeKbC5+w4oaVtu7VNdZnocD/oPD6EE
p6OiD2v88wLfJWVykhAScn5FvpFD60XCYIKaGDrJ41P0eGG234ser5U6HqNFCoBavAO1qVlesgTs
2r32KXxPgNwn4kNalVumbS1Bh+4hgF4GeibmPNvcr2MngaxSxx2X7WhpUbRHPJRTBrvc+frA36gf
LMiIDuBHT7YnTTwp5dsWgPmPNy4+qLeHpKHWbiFpJ8MVbZdaU1Zmx/zgqwSZiyRw0x2Bw/knKKcy
kfwrPdhTaoampqSchQ3GUpiLAiho5ntDVRPx7I3uLvoP28Bdg8Eklqs3zUpdAcQaKtN3Cye0hArq
pNbSVtsthUlwy7gcapRGsPjc6G8KK35hva0svOuK6WQB3sKOjXShPXWKEyHtWzGG6c01xJRzZ+HI
fZTNFOiHN8GGVwV6HYMtfLzR2AgfmOn4lyAVM7E+6vxouPFmxenBf3XeKnxXw1rThZNjvFEbpdD1
0e0tXhGD4CgJkqDZMm7KiaFZToKE8wvyrt5PFHodS9snOlkIFIoB2+JEDsG88hZXTr9f1ya2WUwg
S36IY2F1rUm9EoTK/4mzwkyiWwFoSPka1ewvnnQq0a8ozPg+fB8fal61V5JTLkm5wKXaSI798QCZ
x8DGJFMmPLmdDmJxT2qF0HHkuV+Mmnk8V4d2kuihuaQC4b+8/NHr2jcTInV3bPfIocGJy9I2mZpb
LM4a0ttcybtCza6ULsV5kTTTqwqEKaO902qmzBpZApqMjdJuYvajVsdS8AvFN6n4aGiiYcs0j3YV
HxBokyUIUVKbS1DjiwL/N80iTQ6HjGuC+Sr+skdWzcM5KFbylf2+rau2C0CZqVrd0LKfuKVFThqE
NnKFbybnU9Q/20dKTquHLcYWYY16vcTpzszv+oo9zKrh9orT3HYxk8WgtFpi6qvvIGw9Ozc3XCm3
pMW4ogrNlMBLUdCMlya55/FEJPWHYAlmaA2Hah8Y1bSK0IfaSC8ehdTpSE6NkmnjtCq2uazmfAF7
/9ajSaEsHQ9kSoNKf7fOB/96A/W/fW6sUMt3S7mo/3LzYIV3mp6TpV6Jv+XXu/20bxvgsk1cU8kO
Nw63qzzpC0++u9qSzFWvRzdmys+EXfGgzHD5m6+dYx+IK8Ju6GHqfg6kmilg4rrZvl+TM5k1sZDK
5I4Jk+zHkuK15mb5ElRjri5/QuLOpTH7rrFfDeYZSTfweVTTCA4JhLHlBg8WcBc/CEe8xH2MadsI
nonJM6QpwCwg0437JDpB2rfKhMH0ksgfsbvxS6rFD5JAV+ZgZUojl8nHp2lplxi/eujDmbjEAPSR
Qee5wvU3Dp/zuDIZrX/PtNd7GUGGJlzNGNAcK8LK73ROEKOTerZKK8bCVb0/q7rfXzH0xbCIEPf9
wmFStIaSAaOX10Mc7OhNL7iVPHg3WaNjiSnUKW+HbviZABoEA/xWge0pkYQEAGaQDLKh+xzFjyMo
RyBqRaRC0xcUvtj6QjKO3stL7FmOjq0SOGWWKP0zbSRDIJOlA81qFxTQtrJHwA0N2wqMObY10Ly/
mTYzCbOvmYGddzV6AGiUeDXknyQ6bSciT1PPPQ81ZJBZHc9+dIlD/jJZHPJ05i//CrO4Fg2emgBq
bP+kbJR2NMF0ZegfcrBeKqODcn32rRhb9Xf4dxXLWAfNbDLtpVVC+bKLiAHuWzvfPWvieC8d/v5q
sceTibKR/n7RLdPlsq4UsPbVEKWrNY6cN0Knz2Y/FljP6Y5UuB2NtZONs5IcIOUM5WKb2BO/fxXp
pDPDpKhHg5sVXYywrj+zIFnhP7Ke8nrDozwYM3K1ZLmD3xxQa/Wen+LnlvWLOUrUra8XGIAQ/Szj
99hyudtOb5s0Ij71+1RXpooraRza2I7/GY8NfIY7eH7M4n2l/iLTKw9sF7J0B9uHcPeok15upOX5
LwLtmndOGqxl8f6dJNm7b7gowy7YQ+pry90fiVCz7fBRnYx6c67Qc1YiTNOK67obWHDnl6Qg53vl
2tG/hUyrgn0/1AAeS+Xkh2UJ+TpvatKth5aLYg5C3oKBeQ1sD4piUwrETeJO40gCRXyzwZkLp6dM
jw42EN9ob/bYPfAXpyMEtXO4mrOhPRialJNnr0opXezyYbXWZcgdYu/YPL50R5Smx1kMflcNaFGy
Dnb4tGLGtnMHCxEmrvLlemp1SHvmadbl5h85Hpy4cIlYcO84QO/nfC0RxSojcJv7DWmm2JugoEQ+
RHIV05x9iwfV2qtmwntgHiGwDUm03ESldcvHla5LWEAogL6RmApFHRvkb2fDAXnPrpf7QDkDJe9r
5y+AVVyPNUbl/cKxBh2glCOk77WIQo7M/FJXu/DVmmoP8QLeVd/JD6M7RIV4UZSqVygEXT/ryUht
akj9sL7bCBaBKDi+QkOuN4MLhq8lLQxp3Xpuv52RrnldWBkDQVtCg083A36nQVsTTXVCXYFuFGA8
5IzaKdmXHpXweEvH6XXJlritOsTgyygi7+FpEQ0reIRVoiIHJbIJwysFK8oh2KG0nHkWFnSQopzh
QuoDdLmhy7/BagMHizraakGuu6jFd+/fSL3XWDVFUTpU3GpNJJLes30/Hvui9s6KUao1jkz931BG
06h1t9sG7ohMdXhrOEUJYlujG4h6OHVEBE2ntd9MkK6/Uo4BhAQVVGPYhMJnCgOUUYg3LVHF3cwU
VocQEu00I+ExXdtaFXqMdYbu/HMHaGOQN8ypGBdDigCCUaSk1gA/N3xLk3H1yQqxplLFwCuzSmBa
mMQZxPWIekA00iWf7SUax+pb4FlYawpugw5LZZwKcpKZVjst/oQlOsETI12Bja8ySbF2He8urbXL
zWCQ1Tg9D7Lr+Y53N0kNA41J/Us26Jd3uMH95dk4mmMrFHtGrauk+LuML+td9sfYv3bH3phYQlMU
DepmOZprWzL7sQy0REn2eaVHNcOR8TiabvQwmLKtjaFkTYiQoZnRjagN7mFYexy+qyQIymWuNgE4
XSg6Ixk7BRsPEK8WbPHbcM1+3CWpY0ws7j7dmYtW8h76U2htHflUBBxqhKcoGjhMOnzI+9vmHes5
14W91fT8kPZbYVJi8/QawpCUMPdHd9LfWeuWHJ4rto9/FzS5eJRei06PUC8Xs0e/0fOx+Uqi7Au9
wjHqtlRvEe4bNPd6/debI3bWs1vo5q1ma00HamYPm40ypjH5hDzBlrn02+3Rl7S7nkyld8f3LM5J
BHtHXEQnI4Ns3dz3Q/dnRjiFEIm/FV0uT4sHkHX7ykDK/P2WVmh85wqWtWgbw13G83CKCj0ZBt+u
lhfRVaBikH2UkmsJa+3N6ucTEa0yl5ZMpF/aWx45rocTPbqFqVey2zEukRSI6AmYffXex+PyxN/d
0a06XswRoJihbzgtnuLv5Fq5sY4wo2pidiUMj/Sc2fzl0AFFcNDBr6ezsFkaRFDyUSfFb0Dd6Xo4
A7J2HPHPNYDnTL7CoioPbRe/GMyJXcjWR2WKqNoZUxFvC5BzZheXWhcYQvYR6nFFMRkY2maJiTAG
2/Xbqrqm/eTZIPiBp0OQn+ATPxI56k5unBcNIWee+bY9A2JklEVGVn2Lhn53PK3iwnPm3LwwValn
ah9qoFmTQmwKpKnai9pGGzq85JMf6aWpH1mIIvd2p02mzqMae0i7i3cSFMoHssU3RTPV+pKjJdS1
RbLUkZsy10mA78W5wkZQZ+skuLiQdwyQollixrMH1u4gHEutA8OCToIXyxrTXqrSpB5H7VGh1LfW
b8yUFfDQfImwew4V3heTQeaUQpl/tb9fuudcVSJ7ljx7/tj02+hX24DTgwbDCvdt3M6iP9/oNFiO
pgNCYLHZxLKJIf3SnJl05jaY15Oq0W3VmaUZBznOl6TTZJFr7ReoFN9E/UTVugNQWwH8M1EBDOE6
X4+iPjj6AxGSxWykpt9BCdcUxeQYh/RUXg7CTry/z/l3esE+UlDKi/n9yqkNkkhYmlxYRPx5ynVN
LXyvA8jj189kHbgrTa/0/zzGImwDIWP8BQ/L1dfiQs3Ke+Y9Qzrlt5DM1YHAZws/LlUdLwg7jXHN
0x1U/FIsxMNjEC+QDzzv3AB6FvhMCRSBV/EKCYpVsVP1BsMIaqbCaEf2AfQ5a+PXfxWci5a8WIkK
Iz7xuxApCF6vye3eDqTMfQ3qxGyI/ip4Hl/nKDuh4GVb9uXNNYaBPLAlqFy4N+/nfJDcv5D1b1R8
Kjmh+Ol7/vj5i9BsXS1Glp1nqQmCRmtV+PHRPi0GndtkmNxPdlUNBDJI4WkVRPZzZUj76Jq1sX6Y
hAi+/bTGqcnPoC3JQW76lhFjWuCZM8wdjY+wqIgi5XEVJ3GSdAud2vMk7NKLrFbgDVE4YXXAyWvW
xKRLjISaKtRrMVD7Zdsfx7+tHw6C/loE3Zd7reTTX5LG3CJZ4mIP3mejnnMBgJGUvJRQKwfkmIdi
QvHdf1No8Jf7ju3pIu90C8ZsIHXxxfVJuNQL446DjahmPM3cjm/XBw5GW9ao2k7I6MwlNhbmkkd0
Busv09kzcvYNBZcFnRaO2uDXq0TIQrwFQyrGQw3frSRDFo/7hkwGS4ei753nvfETy8Yb91yoB4Bv
ZqquBO0YeFRr3hJJ0LALq/LTjEQ8uc7UZqcsSoL53fwoA/2qDXLWgfg4wd59dRa+v0MnVuwezdYc
A9xzowNhjPvLSzsdnWSRfIHkKZjjyZ6Ph1IsuDzLS5EujjMmDpNamtS86S5sPbNkIQPVYQv4MR49
y7SdeSRqFuZbYMUVKsc/mikNFjre7QQ7HQ6+P4+DNVhGah5pm6zURXm/NnUaZ4Rqiz+DphpIDqfY
8UCTMjTlQ4ASLVK6xrZRmUE0D1Bp9dda4iJ8vEqdyR+H9H129TLO3jXsxWBDPKp/Rd8H/8AP9YLV
cgzyYj/NXPj6I83O88MK/CGthjauFM6g6co9WtSzfMhdRWY4ED4DdVY+4mV+VNUY95wkBimUCC0C
eFo4+9OvirUxmC8aVUhUyAqmvE+cGD36GNgrr+a/VwYeCkX0JkDhYy5C8RN8WhZA7k+r7ijed5lp
xl4HsMrV9PN60QQYjz7BwWvzZid7Mxbr1CsFxxrzIGovJjtGml1LRiH/4mZSZnJwE65rhiAYLgN1
CV5exlxQc3LhlU23hlMEOj4WoTONKc68CGLMgw8xhBNSkQCvXJ+YsoSIU0Txmkh7PdcdwfO2g2D+
DkFESN0Z/10Mmb15ZhKzfxHtO/PJn941L+/Rf8TM//8ylhIuZglcQuNR/yq62d3/6a+gp5jwrshw
+ciiRJF2NVyykmNBam5ff1G5aJ20Xqhadvdt7OPTWcXEAYXaixqDPiMqnaL4jUhq3wnt3Bxb18Bo
BhqoPVZJa18M4nuYfK/JeCeVrPkmC7HZNRU41i3LwVJP5in98Jz2kWT8UTbpbJYR9rgUgTDcavdJ
ogeI2RrAxsUBKIDIZz26qtXYlLFKORt2Mq9icdxIizlA4GQBPQFsgvKTOw+x4wlxbPjNduoUUSpP
OTIIQcb4IkogfKxVEtOS4Kk0FXgAeMTBq6PyoqI5vXMwT/xO5WzyPxYVOU7QpSFzrlEZaDcfzfBb
VnlIH6qGd0/RZfP3+OEF2Bhz3m8ObCvuypDkdbQVpSEwBJpFb9pdpfURJOwXA2ZbO1ukJHNqpwHA
zjBBvoi4NK2B7i6Zu8rZ9MfnnQRMtm3voJrlU/di2LxxHwJJ0COsgiBXU+vTM5kylfsDAVyZIL7e
ksV2JtD4PlbFR88SZ7xa/PG/U578NDB2LvslEUkRqKt7pt5R4dwhC56g/DHwNJGHCV5fW0hoQztL
gXq9Mqpw6R9+iHwOZZpk5DX2A21MiGMZx5q16Ii+86H4T9+ZWIBY+aoPOZvt0OCpIAXLtUKnqT1a
nQ24fRAayU847rjKFP250H+x6yQnieUBi5rV7inFo1yW8e+/6VgFldZHavUkGkeOS8kL2XCK+FLv
dT9gbUy+76+NxVkSbTkaGVm1WsAtdtZV1m2DILGTz1cSMJLzuCb+cjuzXP7J4BOvUZuAufMePqfp
lq9OVB9SJ6XfbtCtB7CnsO+hN/zgxnW4ZaZIw3B/sIl9FAIxHXBxZ+/2H3leoFlQWdixIDYX62dp
0zdvn2Cz5tIJ2O6FknnSg6G1U4zrwUAkjcoOMHeAxc0VIfozjoSTfiB108xylM8lh93nGXvlmY2U
IhIaGMLEk8BUC8P1n0JdQYgAM4OAzSM+CBWzF6/KF9R6LAY0E1xquwKkes/ZtO/JyM0QSzX2NEdk
a37CjbuvHn+AUkdCw7ySpLUEyBk3DkIezZQgBA+29fP2DTouitxIUDkWm2PKQnfr34N7Yd+koky+
8oANiJh52SZ7mfvzBz6/+sW7xae8RkxhfB22dQdtuPA0ufwZ21DHRF3F2l3Y1s/Jo3Ds6XjuxEan
6IDx9Ih20ihhOyKbtscx1bZlBTfhh5K0W8D/F3cH7CBhinVa7sot320nLuL2rMcCacaxIjAEcHna
IViZdbEwvVCNc1KoCqNL4xB521Wa5+veW0M6RsxMBBQjakKByuHsIKJrTqXDfPYvsDXQ1weBLLUs
XKTWs0Zt/cAsLYwgJWR/5GsJsCq6Cu0aO//T6u1sfv83agQ+J+BpvmFKLIc7f2rDsgJgnReelh1L
tX0TAOVW3KtugQay8Jx7b6QQVDy8to269ExDZASBt3CY5jXMTnybnA5rGsp/urwxim7xB21Qa42g
58LBeHB8U1cnsiBWl4AKIxofvJY6M4/VPISjGrQ3rRD+dRo3jAkJkQpQjcF2mBItNIL3q5TTyvfA
zRpZ6BXuxyDfFeG6MZwW7hWSvJqROcDPlvg++hLWUjk8MjXmOdqLEjrtGiQ/ZkMcexbvTmUb94PT
7UF//z8FknyTcCk9Ibv9P70CJ8evBdBwNBscuAtxbqrbdpw76POv5hYquJI44ooJol+rYhhQfEHc
QzKVMWj/2oa/CitH8oVINMnBndY/9EG28bvykLlRDbjnzhMVBIfth4Xqb/Mz8W+PrvigS85g9bnR
RwskhZuWci6h12PczIdvC9IVJRTk5+FP84vjHmCdmNxGba3jmAF6IvKY8lxTbO8TURRvLywX5c3A
aBhdqNRI5+86wT/9RxMjWDrra4bC0Ms6DEoIkindVljvt/U1/v6wVIYbMnAWSnrtFkEEULsKohQa
0f9DH61xiK2BVrJ7OkBzjrLhsnnbpOd13F36iQmRwsu/FAx4xoP7ptlgilvKXvr/BpaqvifoIBnO
t0y0s6Gee1snhf0vuBJrDIcGmNTGa4GVLR1d3L4IAs1s9zAUajjJEtBHc/KLw6y2GiSlyf9swVrH
eyYcA7mX8PSIQvww6QLzbSVrrsDssoqByHV5wWZqAikGzZZhmBcdYfiJNKF5/3U0QZ3qzD3gpfk+
N1e3P6Ur6Xt3GGNzW+va2LUw8LkZEYr9hKgYKEjCInzHMrt/kSoPsGD2eUxCGpngfRNp/xjpR57o
/vt9gqruOEmV2bCxuwRMm4RwhlMK52jCZGNn9KfTWXd8BLlBorXhvslYhTsm44eRXsWo1q9SYmRH
opHvPOLQ1sLpOTg8aQ57XOzykHtNLSvMGADZJ6vRN5HeqTRJ6v+QupJImvS12Wb0phv9mjJI+N3b
UMoZXhw91CdyVaFd0Ugd3gjDG9iX2Q776yIinFQGZBHkueBFRlE7Idq1W3ToSxLilOrJ4+yZ+p/4
CECXRrD/Pp/ANF922o6LhQjeIxxjw4nxPn734C/PGFbgG9mKUddJ+XvUaTntkMCA4eG5NyQCRgGG
VbPGyGzENHxiJMHHv+7wgW0lduoUR5YAuSht2E8SsRxKB+7wzZL6lCSJU1mczYQP8hSsJOHfNcdS
jx2B4eyaVbxk/qc7s7jH+XqOxgkpRkeUiRKzodeyDJKmoQLJ6dMgoslYwgIj9xadz+TGsa2jSurD
q7yfZnlBGDfcYhkE1hQ8jYO2r1hqQdfWXE51XaONPhWKwyDc8Nw2D9f55LVNipNMTJTKcCe7Mj7H
0bJIbm/zVaXPfb4GetquszTxe/L2edEZEjRjnGQyaXhSAlBWfKqSYUmVphW4B9XzvtHxkLvbJK8o
ra4HNfanY3mTa0Oz3IGEGLLikXjXJBo9Iv9vQBeRoVvUiNMy9prjpeABOh3/VxxMKnWkuI7P61y/
aiMMff8jdyjBUM93xj5eyPGEN5pqepqrpVu5MWLPTgpOyQgiErYfBXuUHY1v9EUwo/8ZAgZczj1K
yYoJQZJV+6ZQVY41kYUbK2VIxkIXlxi63xM4zyogVMg3viU+RImm/DpqMBCx1Q5OOjUXdrONcQwn
o4yeu9g/YAlbGVJn201trlgmHJqlT0o38ZSD4HO0f8mR3Ts4LNljFNEoUDZwAB/0MWhENEnSXZEH
Ny75w1Lyz/O2rIl4gfVEcDJjkKJkCXHU9DMu2d6yNMyjYWnW++TUBrx4a2cfQ55Obn/C2oiQXJbk
6vySzHLOBWfnGGfz3kD07kpgT0RS796VVShU0hy/U0YdA6dMxF+RCTwc5EelCfCJTqioKkkaJha5
WlEL32T7l1inJ7lO38BMSr44bQ8Gm6LBPiwSKe3LZlJlkleLZPOeyMhDU9xeU8pgturfAhqGS2S7
2UBAp8DpC6hoYNhVLJJAdMQGf3RCjA5EvnRAQ0SGdPCX0TIENf0eGL2qg9PdGjzjAbSNhZ7tnv14
0OiDngOyKpUwx/7LQBVBCmkiAlXMR024tEQFa1YytEWvPBR/3FNxK562BYRph+OsTQlNnU3z/hML
YinNqTjuxVBMjGAzT/X5ge+6uNvXHrvvEfIBlfqDBdjIiRpLZyHE7dGt16xM4hAbpn+jUId3suYZ
K7VoboaCL5p4nDI9TceKxcEu5vmeS00rHo+N+VhiA89JUWgP0uaFJjfXbXhFkWOWVYfbIP4HM+32
eM+L25jMRUN65Jsz13w07mOq4oDAh2u/W1z2oiwZppej1D7ir//00qpxI7XHaiq9Fa1sjbyw0lwo
lD1Se/pq3V+Jh6ztG3vRxafR8hZNK3Zq3kaUj56S3ulzslrFn2XFa6Lxl7KHMa9xas8Y2KL66VBo
ZDfSRYzeoLvSQ2G9FOKKvF/LLG4WExdgQp+0PYOjVWg/ccpwN+rvzDxS+iww/jdFgmMXvO7LzFe5
2zEiFRJ5OrEvPR9odLQBa93VDeK+9VJjjw2d5K5VlY99CZjZOGo9WwM+k/VHa2okXk94N7yOZo15
JUSbnS6SUd+tO3MwK905aMN+QOyscXszt3lQlzQ+LgvK0s8iJMkkAIb754WlMv9HWy/k7dNvrRf0
X3O4B++dbaGCcH9e09yo32sZopo+9IlVLrjz9ikw0wgX9R/PgwiPcGw1Ub5WXxgPkmY2G7LFxpu5
bB6742HkfDqEY1K0cCs6ISZ7ECs1/sosCdh9ToVwT3izczVkM8g7dMgty/T61qxKgo7KvPtepyQX
vKSQZ2u7OKs+xYp+7rr5iyrlA1BoB+nXG5uet/H0JRt+sJF+Dxkjq5I3u5P3nz8ABCxH9Ef9nCDr
ihHfldbQ79Wtw5aHGIuwWzHdY1g44OxBpncuBjNt94VKCgeMdlexQrOD8j0YWtMm49ViXwS0HMG+
ZRVwYHTcTdzm083kmcyTDyQzcV8O3e6dB6eyfZPAq0s6zypOdNcqTdCvvCJo5WKanIaSlmZXgTZP
dKQ80g/LP3ZO9P3mvvXprkHhrKCOwznv4nozLurdgz8xlbZJZmFN1mYZA3K+qJ1LmefvMVwhi60H
J6nnqV8VadOBw6NowQYaRZd0q5mhfc8oFZM1SYQ+OPX8T3Hfi6DaT8PVRQGi6UpqwdXumEWnSYGT
0jqVn4W72sO3uY5IKXS8N8P6f+5VNvjERkuVUh+MgHcKuGmyAZsEsqT30kuvTCW18+LQAW+j924c
eFrZicXXEZ3emKLNzQBqpSY1BeIcyMnhJ2YHEPuYEWckBY+uQVv6En8jWg7tCjwF1LTxplHlMmdF
p/3QB0pRUGX8D8g8+zVagbx44WvcQnbmQFvikKfrclNCppzw+Djl/ItFnkMYCHy/dGV7T+itvMrz
NuAKkeosYS/XzO0RoxmTru6vJ4fCPqw9oTzUytjtTHqXAUuQK4WxzT7FaHYasBPBpjzsLE8bWgyX
WbA/tDvfCzDiqVWoq/rnBizniH+fOmvx3I0tWWpsuFSEGN50sz4Qqj4FXDmjMUcdtpNte2GLaDk5
iDq+eGHUGUjDREWs+PDAStVKX2n49U7CvC55UArr1deHgyUwL/99Vja2bbdoni6lQlafg7E+LwEH
DZK1iEd1SBok8PlfKCiixwIwXPpHIb71/iwOLah+aiiubUIRF3Q+G3fEuTnYz5lisrPnLvK2ril9
m5mVaQ6Z/spHS/tzw9QExnqToSA18uz/sdUr5nlzBFKX+bkfVT2E9+pgGFJbf9i16CzAxQfgR65p
WQ2/p8V7Eya0HKf1S4jDmlmITiXZj0wmP0ZsxdZBNd0NzIvoac8NONFLanvsv+7y1dCMycdUazHn
KCFK3wZB61Ql/yQi9ftnmVnfSX8HTTYIF/QbsUsopVRjZqF2gNazK45IODcuyKS3HDtVJ7Xs3LaI
iqhi+0655nq9oDRRcwPNEkrEQZ4dwYTO4skdkD6n80+U9eu5k7D6rBvXh6z3a01iVtPtU5fng4qN
FtvyvRFfOatqkfZtpSvpbHLUXzFQ3xNHqtDPdJZnCju63MPhARj4WYsTPQKbKKXFPqk+UVAMHbTq
H5hTwmwS56t9UPq4uqFUXuHDockR3y4T2Stvk4Oj6VnjpLt6nOtFlVhWmCmY8xgM9iBL2QOw4Zxj
NmejpRJJvPo94jyaNflbIqDmpp/zjD2ePJDHo6fN3q7tXc7926NpSfRCPtX9lAY3+9uM4xUKdUM1
nTaz04HxTXnH3Qcg/UaivjU3XttAlgGYMgkQlEb2FCkXt09INreA/ZvoEUzBpQoeNwJ0VnP2K+yW
Pnlni+Wo2/FsjY51g1turCY1Oe5cHZ9NATBcPvMu5p7HLNpqLLnjnM45y+QOtKnk76SHTddqd+iZ
mxh/T0BtQTP1FzLw9plrQMLhagc2+LqrSTrtUdKfWpqyhL66B4RoxhKk6l0arqO46JUpkGjMEJfP
/c0xq8Zxb6svHNmnUGBzZOBciD3LV3YX5a7dAjWbUMTBpRiATqcfiqqNO85OzJ5NhOQv2jDCUCNd
AcER+dOvNmPE8p7+aZJP+1uRVexx75ldP3dAp9VXjm7qMDGoghGwHoVzW02kIJbFwieMrzFMS856
pLzS90AJIGJ9g0nQFADq6jl5yt9OSj4hbN1/ogaqDsbdLH8CedZe9ZSkX7kt9cEr1/yC6hlPshgW
kMlkhADUeOdqbBCaCE52O5k2UCMnkaxb2An31YZehdrD0NlRcO5JUvu8BLvr0N1DyOcVMhylBkAW
L9S8IyXBV4nk7BmYfsTCnMkRDaa2PYtyIULg2kRCdXSWuuWQ40rqNRVGJfFKlNM1gbaOEv5tyVhR
o+63ZHzO1Vnj7GkRo9JVmmm11M1E5zASmNhuKNaqMprGsWN4TQ5FkGsbc//7k002Fyw9n+MxCviw
Xq238bXCiY5SkBGmKDX120mhnyp/26dBUDkiGJXQYFahb/DJ4xF1SyOqD1qIkoxoln6ojWyP0V79
enIdjD3mvRKR6trmylPaeaR3xsDXXy1e1LRM+Ao6DlQaT6ZJu+inbEfoiCe+vccYgrl6janwBpb0
3pi9Q9gC1jrz3xyLq/ljRSsHX9ScRS17ZP5LspS0UORqBV7K5jWTXLIYOdk1+Nu48gcpSlFv1alC
PBVbTl4NTyXyGYC1xDupegsigg7jp/JgvYu/crUNwM9nfk7ztLWLypQBJhUu2MEwOqdS9cH/Lmkc
2zBJwiTaxc8Xty23OTtwm+cmcOPNFJKLafvBQpeKxwK44Ws39zCclQ0Mc+zwmgwTRdUwFWdtx/+G
7pJiWOvSMztWNHbrZrF+9xKDyOyCmvUilvI/0NTG/2rYs7yCOrOrcrOWZe5RHxb5ARgJtW1srmZS
duEQGYD42lPkVjRfqa+QGepItWnA9w8z01qmWC71reRw1MKWzVzF/CsFrgvJBhpp2niKj2Sj67re
1ze0qXM1TYxkbt65/SopSb74kHMe6TGgK0OZ15iMNefj6WytjVxKh2pFXT5BBQEPCNEihaV886FI
2+I1Kc7133mIARlditJfYEVp54qC/RRplVOyZxkd5c68bBa64+URbET20L6H1m89/qBFAoOqG4CY
Ixi/ckvhr8SaWJyKvgcZuPQ6c/QFVc3OY19SyskDKY2vqc3tUURAEZ6HTYRHX2XQUKnDO56f9jVR
mJXs4ED9zrlXpjFn2ez6v3WYaww8dNzle7ccosHickEUJUz79Quxon3C03+agCZPLx/KpMsBlAki
xnO0yndXBVxDJJaSltDPbepBNAz4YUaDfdHAVNPh4L5TCR4mdnN5aHInTkknHNnlfvjPWSr8PWaH
EF/E8BcwDq4N9UruSKKuL+fVfRIHO3Vw2Wx0fdxMoP4BXAWhIl21/VAtVy0HHs96CtXelyjiOqsk
sutZcTPnzGohQQutiMqfpg/hLL+UHnAzDleDpfZQDZ0bzlYOvLbDz1vu+ei8zp9oWaDq+U+BRoIh
cxRhHq2KNDyJ8F+tBrwTH/HbTfOSCjAjkAK1aB5wcK/pEQkxE4qk82C1Q02ESb5z2ESbOTDOS7a/
alVKgS+3nzcU8R4W5b77v6d7YJLUoT7NeOAFu0w8SM/zhqePiQSedwa8owBnzNF7m28gmHEgp1iE
dvsE5HU9w6jP/CHjqZojsFbCA5Zqc5iBltj3UDum48mZKFfih/CKfkJ+iUIfs1oTjtz9gdlred6p
v4LDr60OE7kcAevWGZA5dVd1MMNjW5od1KnzEycRHyiM0N5C/g8KmYD1q5K+INozA6VhmoYO0QvZ
PPdjcJMaEGCXT/shf8bW/gVdvQRfrmQrVYAb0QFLxu7dRNjlZ65ZNikG4oeb0FkYhp1l5rR7V6MD
wQylDnRNuBGPU4dTRRki+KI5eyCEHkGgpIhJwncMm1hahUC2c7EshvVfik5DoFFjdmu45ap7Ib2S
LXuaKRiKNI5swvlgjreXm37Zh5/RsP3YhsHhbCOV/q9lJCtc5AxAcaqQX9BVjKNREkts5xzoW1d7
/C3cl2cIXZ6RdSY9AQL0MASyf3otSG5aovBTNQv/8+Y2wPoKTYquPf9B+lgrzMkOsFWzJtSK7jkD
L23QKlAg8lsRNdin/rNZzGTC8+Y6958fu7u72a5VKmGl7KkEfWikNjx9aVeUQhhKWhjA18oqE4rz
2qYmTdtyCHWm5NiczWfLYuuE4nt8587fUM0oNNwoknJRmmRglypMXFo5r4GkRsimvINxaPatRLAD
LORU7jeVuwlQtLW/gJj3mMVSWFeOBIgVVyDgYCuZEtQ+2c8Zi8+w6pwau9ZZBGPhOBEwsx/78X6l
yCclz0HpSAyY9coFAUSX3CFOIc9DnxDTkEyHazMmYfJqSWhSb5zVJS0lCLI8xF8YOSw4t9P+Cyr3
GfWHIMHAaTIEOD09tD54Nk3VUp4chTgA2NaKI4JzcQR35ik0nIuG2dJuyMvIMN5EAqBC/gHpkf+s
ggGmYdjFBjqfBc6tQWl6mYfWQm7015pnFABUCLUhouoCHmPjjZ2cZKGgaXu3nlcCfKLR4dUP2P8U
0TxC87JbxHhFBKvfi8xRwToDV5vNbgvFg69v/v7aeJXGFEgpjvbT5oMqSH2VegiWpu9hGQO9Bx4A
D0ql8wbcc/5Rd0AQyA91ut0px6Z5WFjuEEeLBWDpu3+MpBL1yxqM6xdSMMWN06zp/B98aAN89GLr
HI6qqZ5aykHWQE2H1LGVL0PFeXWNNSbWeCd+e3jAL2O/P0DhGhrjWO6nQGBQTrJVle0+kD+N+GjN
XlfFERLCX9FV0FuZ9lAwzq3sy4IIcrQftV9DtnyoUfH76jDK3MgCZlQbXI+VksLDTDUE4AXx6Pd2
c4eImqAyTDXGX0tPtmBMUY2QbLpvrfLSjeaTQjnlBXOrpodUKnzPwyPcWB8y9yq6IOV8hXFje8vs
quPW3TMQau7jGrJQB09zbaPMJs+UJ9B5vYtQn4kMR5I5e2zZCpCMU2khgxump/RK3zKPuDkeZdvs
EGgnCT9/HNogtbQlHavpS6aIS0eQ9gM7Xes1iUdaH+5M713kGTSOObXacB+DCLqBMjPqdDo+69jt
S16hnslFHWvKzp8fOF7ukxjU2F/iiHc1Q6tvKM6pbwTY48sBp6Qmc3Yt3F0n7gbbIuEC0DjWB6WZ
X6XtsbJGf8JtQtkyPN9Z0L5t6CSgMzOoaHkt+zyP+CAFoofLqI4mtbhZYevNnbqSLSbxhxInNju4
YYzucazvxmxxgItGMxl1QOBHdwc9B/46M0YWcklHYzqGDpHHJ8DzaJ9jCLL2dD22PrYOb9ZybVts
guhNNSymn1028ZfWaXOqC3mPyZWq/xtvWcWyFHQj/2+m3472mclif59On4Xw+EJL5JzgGkA71Ylo
4PrtmiW4ipJqGsOvSkP3CVjwNBGgyK+ddWxWfsAW3I/HwONwUB/1uNEj3o7BO5SXvLf0K1ZZ9ZtM
MNZ/hmS//EE5MMWeIqXwFjqmxgmtV/iqX328hWYz7vds/uew1YsaKCWPknJhM47guNnpIH8zzY6m
C4kwrp3EjLgEcTzItegcJY9kkNSKOfgIswwyPBZl5fZF2PTBLlnlJMuGVvSqCTEyfVBsCu5y/zGv
XmgynpiGlv7M6aG1tjk09FVl6B4VB2gEl/I1U5TUEp8KKG9ykwFueffMcKDSbSO1K21Rf2KIFxsF
09a8LmOMz0pW2xZTW2+HR7rS6A2ET2RKMTjP85Vu4hIHDb6AD522MbIzvxznCOEwoYYCwKjPLuJ2
AeMH8TnwlfdHTIzFUFedvBIz5MZ+fSgq1YpHCMsZHUv+40fRhgv7KOja9WIVzlFkrxspvpqphsmI
Bgm7O1YRsgVs7/bXExvYSSNY22s+aFYj3pR/RMClcdpwfArxWGpBGOTK37oLqSEaA6P5h8CJdO+4
9e6Z7EOU3MmYGNrpnWdjKiAcRRJCVDoEK60fMfBLn9pba3jmVstERf5psH9F960i7bT4ULCcKZKG
eRB5CkGr9ucoPdaq+OIQeQDY6vK55T+z1goZ6Vz13stgzM7RmEFA4U5dUw8AYWoLSUNDNuhgpccA
2RnIYF2/S9f5v6H/X+CEm1jwksWRk5/q5Y7WpRfcQsXdzstbBXapEki4vbO/ipNGC27znFHIAlD1
mo4GWLQiNwX+yzdgv0FxN8eE4/sA9194koGMt8uG3GAwUdu13ZYZeYWLaCwJuzKDWnY8FA1bnxRO
5B+RKLsg+Pv5DTTSNROgwERbtkey9RyDgTFe9yYUzT1+jsdenlVrnwyVD165vOIfAkmN9Azqi2hE
9zuAGmD0vetBSSs+rHj88XrXQgilF8jSYSCx4le+z+wuot11hxdZWf3XdLKZlHO72Z84Kpfyxdo6
VBogATgrnTRwAcnxtVhRDlDmBelo7etYYmJfCZfbCcKCBXH8qCIaBAPxi2RK8dIpmNMEy0gu00vL
HcMIIPxFdPjNiQYNWMHXW/dj+Du4QR0LTRe+WFblWvjow8w6T3nm3o4wJKr+31OAxIWYFcNsnXDI
5YyHkmgT8t+oegWvsYdl5BzlvhzxZsB1eeK1nx9gNZ+iO9/+w7wrU+ENg1GLlSA/FqNoOnh1OLzp
FgUHL/JeB+QL4LcvStsAh6Y2S7W09v/Xqg99+wYicZvFGeOpLmuh9UkI4Sx1B+SQreR6mkip/h3I
jHEvA2fOtO5KvJwO3qGTMa96pbfZh49Wja81FXdq3OorF4ORnWQv37tO4ihjm0sxOeO70AaFvWoY
TP7eetzZeRqKYU4QEQYH5FXNzo5Ih8bw8dqYpNr67O4HNk7RjuYzagfjlM5oQpl6C4YUY2IRZhuX
e2awB6MmA8wS9tvlCGX6W5haJF+rOrfP+goMEZlJjI4NHe/RwvEVJgiO0lDJgKLNnbansnSMsghZ
cGc6c9x+PH4GabsZJ2CjCSARDOv1NB1AKCtGpF9FVz3shSLHAjLYBPwD1NaDCBzCCt525YvIy0/G
DwU9CaGmmeGrSBdvm0VoBWJcueec9vCmJ8/Twn4aJ7cO+E3JSL4uMe2QA/mg72ciXARG2Qz+Btl6
W1bKDiNUp9UafbE0d4tEI4b2rovHoTzpvplGyoGO0x3jBntUheJ69W0NVDuB+C7zxi9ZYXhrwoLx
uYKiI92G/nFE75VvjaARpcYHnYeM6ovYxDtB/CwFmrwZzMVB0hXArRbXjR+tMrxDR6GJqzTy7QwF
qffBFwguhTZy7uyNQ3FZZK+sUaxE1aad0u5oNSAj+E5E5Rhz2OJp/1K9PE46Ov83wZ8U1Pyw2kbS
IZSXtSx/hTMSS0gz6xL3GDyc5UiUCB/DPDkmbBKbJ7Bl2LoXHtLoUmOB5BK6ur+u3XxDRFjkL7z1
AosxkvuOkJwluvgf8ttxrdiaDhSAIhufAZuRsJlpUC/NNRRGD4lfX68GuJO3luHygWgCdXrCfK7A
/j80pwVybI3GCjyge8q9Z64s4Gp+DsinigIfl25AO8OfqNFHAQ4ynv9TVLjdai9Bib/0l2aPQWJu
pLC5ubvALddPneNp6I6AkQDr6UD8MJuQdeWbYs/+g09ska9PQHWXQig8UHb5gJS6CW/xEeDFrTJi
J7jEuyix0240jCL34XU2S/zgg5dlG608xru+sbaWmSaxYGj8z7CS53ANfaLLu4SIxO79fcT5wR8T
HLgVpQ9QOleAsb/beY95gdVJgkGyPwHe/k6RllXC+8emP+6HQ1xlSb0vs+waKQnpk6hfei8AOkej
cPiMD1shPnd13lpamEnZL8rOeAlvv/iyQYZqCkJ2pO+T0alA+jTC5MjIda2dfOztmYzNKZf7CMwW
CwTbiP6x3YUyZKSn4Yuaw3M7F8DajargPiIq1tsy43EY9dxMs6KRhX4m3Md/oLs17KGQk3RKS/Qf
Xauj/6K/6N6nGSEkgcumuyBQi4neeCrSmRSWIHdMAsC+ZyDqfMmD9zbyqzSXKpBefn+dBL3IR8DJ
lsIlH6vQPG42D0DN74EwxRt0OnpXGyS/iw27ECZQC37KzBtgKlAzPZBeYYN4w670PlLEITMskaqD
87EVlxw7YwZbEzN42tBuPNmL+GBzlcDEU7sNywzdI2MQfcjEVUEadKZzobdv9rye/auJCUmG76Lz
pqj2RGzbt3o1yAa+/fP8yzSpQGsipWTUcbZTLYt42n5qqQ5whzknY//rKXFAjYgE6tDhC7KIgzF/
+57CGaCYiygukgr7FEbamgX0gMKvv2+l8zrc4YAx9Fjd4oJHfntbshqunrhNfZFeVFxhTQvHGLPi
c+1NWE2lj5KlZ8IfeXcvCl5UUjYGdFU0AIRO4Aavi504/wa2ER820NOg0jUYHVdMa60q5vc7i2Sn
PKX6mVzM59pN+NKPfXtN8qKIQUlO5akURKrvvoG7uT5fB/Y/TV8wdbVwKUxMvKCrKW3ICcJjsC7u
5KkFI4EukSNkb6fCQ7CdW7ut3+6DuobR7V3UMtRxHmTm7tqjZl9RRBKGdvNSfXsM9LeOH0fhbMbV
PpgAeytKsaxEUB9Om5YYC31o5HHV5Be9MIcUtD3NFDFlydyDZVWxyW8bCQayNIPL25nmBBvECSVu
IddyxgBOpE/RCH20GtWylmdQdOdFsHECcZvtGRYRcVqIR1vFGkwINVQtyxTT75iHtxsAja6oVoMw
kYaYowVqqFm0mMMKpOWCI8pSnYE8vN2OXU2WY+I1eN6sf046ftaEIpc90St8rKlawp0QJbQeb9Gp
8XYyxd5i1iUk3r4ml0Dv9Hk6iweJ5ODz/4FL8DOBECBD2dclDHOsoPUmE/XcAoygDwuSuMkm/8RC
L9/wJGSnBE5qYzIqvxXg77rhJPB1n3edtvXgX7dRffifB6Yt36x4LkEopRXQqJ+56K03yuKveaAt
uLFz8rwxWV7/VoJEbYTnk/tHc8j+iayy2L14DDBTEdaqvrSW3RIM63sYZamyiXmd7NEQBn2oraxS
oF0p4s7glnPbF6L+RFS1gWTDObPc1/cOZE358j27Z2dOviUgU+a101HQAqgKxB1VR9mLip9LoUoG
HJmD8NdPm+fXad97uWkaytEPVQFBUADo0f8ahnUHdUHu+4w3mkZUKZuiJCyRVdbahxtvNDjFJ1u/
v9Y4sNcl2jy3oTKx+FMfcWp2EreIU1WJcrbFP19ZaA0piYwrHVrIMa4Jkf2y0J0WE+EYVWj5nfdv
rJFteoSiJVVBakf6EgFRSjjG9Zb6C24tDMlwhfcEWcxabaTv9EgyRobiENvdxJ7qbCMO2frh7L8h
h0pi1UrU/9bnTHCUZBsLsc6q5QvBHU0LNjZoobEQubq/ZRirZ+Qo8hFPrUXXnnWZbk8ZPWSR44K/
qHTm+3oHTu3Yg5qZaBzP2PTgY8KbWE3w1uQ5M/MqNPs5gXTKgK/hnhid2qGWdvuJ4M5zSEutvrDl
tBUlJqidRFSzLAb0COvizMJqdMvXOdd1oSS83tPBTbbXs15iU38U0jCPPdaENx4kyZKdH1xTypMv
kF+EUAlI/SfL7p3M6DjfEcAhWApvprHkWTRHrkaEU/fiIg+4lDbXb0LjP1dap0HCyfHPp11Frgll
TWXpPSxfsuvsvvSjbTSlB0Gm8jnauY2rBgDfP/ZkWheYx8wLlohR9O4jSjWDGjpf881YHPDaijJ5
H9nvKyDY2rbFA/ueRQo5vKo2nLezOPNlVcfoP9FyE9+XQwo6k5Cu21ShwjjjniOwNfHmffoork6r
9J692ThDqcWAACRl0gi1SHti7kKvrh8GciEIPhgQ5hietCGwKUj4bLHO6Z/SCsTz3IYH61m1DYad
T2V9aLekEcfJXN271UF6XXF2MsAFDnKOZ7EsllEuH3YqOfC07Wo68s1VHbFEcGzH1aT8mJVQs3Dz
4hznu0KSEKZURS/o99RhSc4vF5hi6i2BZJrPSD+fQR5j0Ou8aWCnZj53+OwdVu/4nMLrX3AC5YEU
iTgiHnsDVcmdmI8Pf8kwHmEPq0oDbJJ6t/ydTnjIrEBaTKoFZevRArum6ekgIC50RxCyIhVjUfnS
fqC/u6XG5UoqxvN75SrlopkrlH1yPV3EuJ8U/ibfXD3rgGkYvp+/SWnPWstSNpMJzJ6fwKjzUrb7
+7PMecVZaCw5hOA6Axe9/W1sf4lmvDgjvY99VopZQ0iHHRGyo6ax8UQGN2DnTosqtfS3mFnMd43Z
t3MzlPASr77yxbzL4eb7yZEKJhgXBdO6SLVCS4hFrQmJV4yKMThMjov9YAHH1QpHMUxPmJ8oeh87
b4oIIZ8HyOpl9lIFK+NAuaFld0ZHTum5pDdZybLtGYd7kgeaF8PiS0vL6SE1hU86WbkI4de5dxLj
4FO6/Q5GK6IugZVPorSDfxg+sdxef+vXanuNTK2MGhJnmcJ+a0nEE0qkh2X7j10j58ATbQLxqk5D
NLabzM2QkapQFc5Mfg4Gtizr5QpiXW472fbAhFuWroAI7RVxwjwpN+oKEjHmR8s7JZwhf68EcLJE
rGiiqJNk+3Ah14yWUftrodM6i3FS4qS0x2HV/0BXfW2bjbwwz5NZG+3DoNUGIF6xKfuoJNtXwCls
O198tWjCihGoFj88tO7+ze2U28GjRWuCP4S7oqNfqOsO9RBDrVa+Lj70ErTZlO5Q/O5va2/gW9An
w4mBJ53kYyMqEA+YsZmu4AFSxE00Sd4LCrq87InN7flbMx8tpFd3cWKASAA5EMwEL47LL0TfQFGu
g5iqltthD4wxCBpeRAGl659YvcBMvLg3jh28K4YIlBoklUXGj3LJBK0tbAyw1ekwWCjfw3ZYQHUZ
tyI4MJ4WPkKLXrUqBa9dlTvPDyyT35jf11yt6muoK2weBVpTBZgVprB/WVZXZHV2Z4AizW5RPo/t
RMAYI2pK1PpiadUVovLM/VG8OGnj9zbjKdx9MyxWIWHxvD+jY5WYqUgbDS6vlUSbAueIiPPERmn5
yk7/cSwqCApoccDdEPv2nZL0Ik/7q5C5XMd6zF8qxHbR/2gjwkSq9LtMSvIgQpsQVyb7fbCixlib
1rlLGrtba+mhya/CVM0qkXyoZc6h8KjC7IXrv2k2zzdryp8BG4r5X7q2gmCbp2NHDCKr9nqEtpoM
41S8i0rZknXMRAHyElH+IQP7hkp/IuWXmDHlazsV1xjvJzKjUPRJejxMv4rCMIP4tN4Dj8V+Ishe
kvkrDXVcDUf7ZpXyEAWM0VIk5xHfasiI+CHvHJwnClAw3B+/5GaKE5RiZemKxO8XtY1SmV2YeZMZ
Vvlsh3j3J8oaBfPlzWLp/o3gguTWnT5GYQPUMWHP0suVm1DD9YoipjRD5kTqw1cC7MojRwgKql3X
nFOzCKF+y2ikkLnMPQKlIoxT2BmqslrzHezk9C6AkiFkRKgSU0KqF7h5ZQUd+qWDkD+uJb2efRu9
2hc7oDhWMK961RSdJu1uErUD1A1eaVCgy2rgzg7F9kmDpGmGgOAbp9+aKb109PE9PNsBsnYAgjD3
AcnU08A76LTmcpHdqF3fAEBAeqWxD8qjyPznJzq2bcEShZRHs4QvKE/Sx+8rjZn6pXPzFi2KVO61
670aV3G0+POlEJTSShIJCMDyYc1xxucXLU7MTFBrgU/S93jo5ZyEuONWMHvDSVFERRYrLpbI/Eep
+JZXC502iQycQZcw8zrOGoqYh0+JzMjy79q8ZKp9dIeHiyHj1q4IR9QtlBs3KHRp95RxxjJj9oa3
WyEIvQ9fblTE/8TJCgx2hUXzFhrWhpaxkOY4TU+sxFzsrcb+RgqyV7kKn8Qrlppv9cbUuGA/XNUA
Ugp6VjHqLd5aSJiyfPhYSqvtsGWSmAiZ+NIyLYo0jnhoR1CKA6QOtNBvbO4o+bXFU4oK/9u3gv4K
cMq+8cVjcM1S0DUisKfqJUCgxsZu45jkvxBTjVed2P8NkP9ZnHEQWJQCzRtRZrjFo9oBvRB77oFk
vyUm3uIaSKjp0PptXwrLZWCuylv7478PzQY9cpd45Su5quuEHq5ZWtmKVTfaIuAgSMg/ldKaGHPb
MWFv2p0VsnRaJmcI9axpsVvotU5vwJXNt6mU0A0126NMjrKUWmDXTh9J+8Uom3Zh9LyoEB/hMkJi
fK12drAmgV5Cds9/JNgAZZMp5q5tlSE+9b4d5o34HWzmsl8F/tkWQxFGn8iIKC21g0nKdOVcaSOc
IY1Rm1k02wvz9TVFM+5RqF0m2Ul2xpmSs5tWofV67ilNVeEbiWb+ZQ1qHW9IljcLaUyUNjFj8Lul
oURk2m9C8OxLMjcN2VkHddhko58dVlWDYDQUIpEsdcTIcB++t0GQFHv+gqyJTQS3snpFcWjMW/jW
ja/3pi4R3aAA5fi2lnReTmMzm3Z01nPrZZ8cLYbQb+QxrFr5On3h6sriFInB0ldNoPttv9jX1nSx
iXUrvdPrFgb2NE4/wZ4kxZ0zzkUvBgPiybjiD9fOLH/FKr4QLSZlqMxQ4Eoyeec/NVQ6uUGzeegD
noR27z0zvsCXLifhGbbO60zjaHyEOw/PhyYZHMfOcy8TQ9O2/HIBH4xktzaN61HVfPmMFlaWoaZe
nz2X14kaiIglY/ueZ+713AcAt6Oy4Po5xToeAC/+Xt5zWtt714UoZ4VifA/v59KuhQKHEMzHSO1h
gJs+brrrr9sg/KBZ/EiRz/enqFd31X+fWI4U8xb+CaQ3Pwr2efPCzKPzy58VzDbbKilNhnWlfsik
SjL+ny5M7YIrg2YHkHfs/KRWhZdBV7RV34qx2B4fma6eTG4XdoSvnZ/eATKNvlJNEiBsOZNxRHQE
cKlWQFpHe2ukhesNHuPr4ViOpQiHJZXGr8wleswd9HQ9lBfxD99UcIVKkAMmmw6n445oXiYSzCBs
fvTU+ULR3yq0zuxMewWSzLP/fvzlyb42RTZ0ns6R9fD/4cqBV3wZGsAx9GGIfLaE5ODaF6RbfpRo
2mQgQv4s9IdWrHqqb3REjg8WXBg6DQTaH1bsZ8+BIFo1e6rvEuru4U3cy7cHk96Nk6T9XvEJgr4Q
llxn82dazmcV2yIQQg7iPXimKskuD66Pu4aZdZuPVW3WnreHMrwRxxAgx20g/qSpBc5wZouEoDES
+fenYvc2Trt7Q0U6aAGEDIwSMnbjbhEGcJfg+16T6C65QwlqExU312hUq7d+UADiOUFzQ4S8v98w
9a82RMYa3MeaPTPdbZB/0QBzzKdrnIL9Y5JPNhR1BmfbuHzeDr4LqxOB6URFAoqtNTTV1OjLYStx
d52LEqw7ldd8npcs2rz8WlaEkdtHAor5IWKxQyJwI7FEm/9Zo75DAdVPBJvuy8VI4K+1BEcPXww2
fzDjV+GVhO4km5LsySYirOwjILneBGW86b+Im+W3sQF0qS69IIDtvm/LS5qDBwHEDu9lh9EIvwFh
wLjyza+HlvLp8mY+oDycCR4/ay3ybklQw4dibTasCs1hdMerQ+6gr3lcUuHBczIRCX/WWoJNu3CD
tCkqwz2F+WxwoEf2zktN6Vg1Ho8lzW9CXSMoYzzgBZb8sacAorYmIF4vF++a0eq9Z3eRspAe2ktp
5j9lkA1UJCHiQYGTIkGbZnP5Qp6NkvLX7dA7ZI/ebNMIxxB+RWczNx0Oq/OSlEI/TRPnPqFyxVp/
LKWDIczXbzKIi/VZPo4gkqZHwBfD1Gy5/xFZN/r1v+H7Uzc/FoxpoTAEscG7SJpbPhHuYOEAk2uh
K0aRD5jqj4QR9oowJ7AJ10n1+ziyDg8UA1B1sGyEMNC9XQ0aYMVPoxHGfuArVqlvwtbxJsM2k3qn
uG8OXPqVPqM2feiyS55boGt7Gk5tXS76Aavd3Uai7i8WPjyIuM6mvWqEdFpW4YlYimfeWn/0nr6Y
YZpRv+UBVBLsnjOjNVwHDwgCx9JFcQv8LHzxH+38nr2ekPKXnSIHJvZeRZ3Nso6olA4frNQrBL22
Arxr5PBt7ce1D22Nt02FggPXtYOkvitxVuOBaOksXRWbJ8yB4iVIjVW2DLDUl9sqJldNW3H262S9
bOgv0kllLV9V4x0dXQvczr2KEURNTLLIMReKWLREFPWrrd16lcrTfKWH0qB6Qxp1AdVw7R7sp7Gn
hf7PGbIT0TRrDAW3iVYKUKVWv0pwaD8ZTWIlpQGQIYN4/78vOcPv5Ti+r4vp9z1Ey0l7A9k7e9UO
kzgvNZUjVa06uXiXnW/HopEDGjJqGG6vkvSOeXjYwa0e6G8p4Q0ZyM0Z2BgqQEdj7yPTHxO15maU
TiqJgwgMN9DKfBYPbemA0aOH7n5NHM1JXNJYaBIXx7yADl1CGqm9JdGd00SaPuodO/kKxL9VXzCI
dZjutrQA+bJ1l4Tj+fbQFyxYK8BaDYWE/e4hfvLpvwpNY3W35DFQD8cuFuXdEMeKfdQ66F1kajhY
2ye+6J4CtLANAh3dhFueo0kdQ/uCZzjhEdY8lKfYRxUjx0DuRFovK2Z1Qj4EReUkDg0pWAfTiwlX
JST0GVcAr5QaTLpVqCTW3VNzwdhIvfVbNW8NJ0kY67Ar5R1sFh/6xh9iq6wjOyxiqQtnDx3D6E4M
Xt84/yEYDIZT30yBPgEhzHkYZ1jQsjmM+AJPbxIMhV03uqe7Xh4FXxUN9vIW3TbCWoWMxBRcqp4p
ePi2+dLuMuE5zaGGc0lkvHddj3L03Rnno1BXx5zlaOo2n4rFskqRjLn2iY9t+Wp8jU9RKY/hwGyc
QMXWQ59wBf8Zy1tkZVlir0yJUeUaLDrVtQD9jhiQvuIxTI5IvKS0OHbecmrJBDxUCoEGa4yUeadZ
6FI4AuRMEaKc2eT2FATR79NYNqBkaT1KQZyntYf0Adc8zzXr8tsl5dZmeuQB9G7fXVDdY7ao5zL7
rxuqY6eCDKH57TWsMElFz17og8w0rOAQ/8r2NlyyBSM7NzTyqboRE04xkJCdJU0qRRXPPSoIhy3m
qRdgvaHzFDCuatTJTSTpREvpsfETbCMiGKjnw1QMjMsUFdH6OUmf86X65wK9Vtvn+fGyDB7OQV+j
NUrCvb7zUHQgsemFXvxYOHc2XXfj/WwdsUB6LiMawFbFgbGOS1pXJJH+lNMWL94WurXlUTGYtqgK
aYGYbUdwlTfdIEMvS74EszXSFiZwB0155BjwHYhLr0Tn/stJwUjNIXoF5VxvfzqWLAUmqqNAomKy
khhb9VBKWQoZ7+neS2J47zbt48CtRt2wYl5+CH6HsMbfQoZ2NjuUYiKMDoXeeGvgAji0bD0UFed4
/M+6plkQ0Wzt5Imo9xojBhz5hhlicV06V7V3VRCXPp6tECHKwa8d+8wCP2dcP1pMCD3XMAMu+h8h
05MeRx/AGJtPpQDrXuli99zKoHo3cCBErN+0lNx0Y+rCyIrzcz3dXDxPElMh31zHz8DefhQMzMzY
3Y3+yHJDsTSnf9UW6R1bYOeDvHtnMRnYoPph22dkvru/7ru2Yjv/BJUk1jAZCWsovP3L824MiskX
fMIrMh3450m3/o8kFc9oqrh61tDrbYbGBgQh5aTgeMGu8j+laps7b8qSsYRR+SusSlc4DpTuXsmB
UHXwigGI54p0WslirBdCih8+nIgzYt4SLSBoLUfo5rfY/8JZqPFHm1XME0+viCJ30wUcAbdy0akk
czNyLLwoar6szl8f2rD4uGF0QAmxTSXhftNb1J80xmFpn7Sm5ZoArH2CSQ4UNtf50kb+RUcKxDT9
31CvEHYJ44p6ohnESGts2EPlKmbAD8tzhhWD5i1U0f1EDX4xp6M7fcFWHD0Gpuzqby9Gu3cnqrmK
WH03rMmOgtnUkGkd7AHp34jzftlo6uMgQnDE4cSbcd0OyX8JpmAFL9rZUndVjW9QoIniWJ0n+sU3
1mbqxfN3+u5I1DIsM+So9N8gDNBtgedrfcmVxUg/FYbkky0qgcnymlahVUxSKiHFdqEzjPTRVyFh
0+204F2NRi8GJwJFVeRtjXDw6jAJzDXZ3bFZ2okMu4jcKeetEm0ZkQTbPkkIo/T+tx+Gtfg2Vl9M
by3rcgOI9DtqsKRCWbCvNDk6o+6Z14te48kyRbAO0jYSz4QNzqO+YEflDoCbs+a+AzcMLOzsv/Pi
Yfvm2xrq07doNSR3ypP3TUfM7tvZF1cym63s3zxDAqucd5kI3DPOj8kocJ2RmC6iHSaKkLDZm8gW
Zrm9E7VoEf1fvGPngfKZzbO8DwxvlZJREHnSomTsWBATgKSflhijicAHRjaxJe2n7Q63lO0HFwLA
s5SNEiUkA0QHNUvOClwSJ9AfJJuGquM8AP4aNBL8F+TaM3odYWfwRnz+Cio092DrkjUgKYul8Q5d
AGyCCUXXLPswtR6Ox57ZxD8L8aLmwWnhXnt2DWCx2Y17YudTaapKa4a7ZZdYYDnDE2aGu6djxAdH
gP56fY3xL01/Wjkc4ZVk5+tXPNsfT/VCbXY1E4Oy7LCxGHlfmiej+jxDjtLiR4LYK1HqMMLJBbpd
iKefvtMOSYdjtVON6pEbl5SGWWv/wh5agmydKAv9qkhF2te30Mo/9VvU1KCBc0jyVfeSXfa7NWCO
lLTd1AvzXDif5JdYM+/pkXK4q0vg9241BZOvjxfp7jXW6j0CITd9ZIO+ihvU9JG7bX0YHixffVsp
yFiUbW7yduVc8r8jvsMt4R3aXSe5xgY5iW0y2OKbG052SKo47qiGkiUERjoNQS0zEWzU+LHwe2vR
KWTasZ2qh2/YhOYowLi6g1KzpBR5AsGARmBLY0u1NgsYdf+KTMHjtEDcSF/kTYYkUASsmIYwTi+r
hpe1Gs1EnbgFtjJ2/lT6qYk+i8xkFxg9vuUJYpu8OasBu52mTXa8FPZlL/VeFwE/5rWNdtfmcOd9
ufv7ONjMFHikz/SHYXFteTag6mRKoRstWPdGECd4A2E8XOIJ6mU8eFon+iMFItq39eTKoFdA7v61
s5AlfI0dljOhO8OPnOA/R69dzMzK94gDRASES5pLsKVUge4GE7e0y5lSiMoQQVZwRZyCZDCjdU1v
YnjuVv+Rus7E6wjBSNpMj81Km/pYdZlwyd9y/28zvVK/K41nsoUkAcoHtRy/5KUvecDSdJdTMziW
0rlLS1jQbx7OQxMLqGbqO5HPm79BTr5DgvB386Ls5viljIkpZ2AENHz0cKQAB+H/e8iO2WQZtCHo
ypqEcc9pmEedM7b00URpPeOjkMjmuCSCW/sTIGGxKMvwzgOWjQSeKlmUjJK2UdzjaT2SiZO66TXN
CKepyLc49WZd/NCKlFIUuN1mBUY3N7fm6LkeCAD22FTMAueI+EkDImlbqzaT8rtTsRlHPXmpOH0B
GFuZRcvXSk2QRs32kds78QqAQq72AkxNEEeFZRGbnUpzbqG2c5WtbOhLvAn/NfcZgxZAqJ+s7Lox
kVJKgLIM43OKhZAJWBbIYUOf0RbrZcI26dw6qsk5ClmDn94V8NPJFZ0DGLE26eG8UCtaGFCAJpox
Gxfd5OazMrh1DYPtW1No0m08QQP9iSb0xG5ybqLs//n/TvqXMXhtElzP/RM3B4gb4DAwLj/ppHqK
sDGuxUarIivnmnkZ6vOP1KoPltpNRvqs2soiUUC688Gli+AP3JXOhea8qryVToukF/FmQfIwLvB7
J5gdF8kC2lO2jpy8ax/T/RAb1j2RNPErYzQbIvGWFPrQ1c7Wb93iWyzM0YP7gH274eZrNh+jkueN
m7s0vMfV98N++KRsIi5TkxDCsTO9+zgs1eC8dlZXqz4DD/PTQ/4g15T2J6CM2sJJBsNswYZM3I8C
O7we589Me4yYB+aFkDSCBJzUnn2nyw+9pui9QjjUAmNluXmmAkaOA+RUtakKMQyuy0dl8pgBepc4
AU1ZDBXU7Qd1uXIh6hh/3fb6PkQOo6QyKy6rEDiOCCWGQs4//JyaaFUf1m/d53SVavieQZdSPqG1
TFssW+I6VTNa74VPGVGnFgjUQElaHRSj6bm9OzlfdTpFrKDj8+ppC0z6h94NTtCkjpi5Dwwodthp
qPClm/HTgLYMCsqCHniIzIOxPQxFdt25RNNc2r4fh7H0wXAQBlmvpqnM3JYJvRk+DR16zRTwksOY
ag/yi7B74UkBaUs954kLij1HgbUTGXGen7YyZDRDDdWoS04Dvp8RwmX+iDwxBeR6t+Q5YWghyUWC
H0ijvsmGpxqR4ovbwbSv+SceNVu2llQlKyDnloVfW7ojmVeP/Emte55ICIT7lCysD7kSHkp0O1FO
8hIV824vhHNlrt/Gg18cOPPtnnmfDXpiWdfeELfGDDuMWhaT/gBV8EzjVBJjiFMa8DzXfiAinHQ2
IMN5D7a7U9QEe//FOPOshM1yfDiAAGXAtirPEqnIMqYKMGsRwGi8WjQeyIMQ5dt2fmMEHl1+H6Vs
wFPljCJIKHm0gkc4OW1rpgzha3CPWM70uS68FAa7Mt+hFHm2lL53mqKJewyCgeqC5D31iXNRA22i
4/Bw9FBTKraBy3K7RlENx46c/gNs52OgmiBmWrWN7hSjiiMRFzz1Gri+uQ5Gtg6GM0Qo/L2D9FiJ
myKsXlfhYl2J4Q9ojMs8mr0Ax2Kr6hvYMpulQk4Cc73PwYoVNyLBo2g0H2HvoivnemvmhMu9E8vT
F68qVy0fDRahtBWQD/LwFVRJCMvV5HZujxmHlEWxMO2sBET28NyO1L13EKKfkzChHu03YQ9u1aOI
ZEtDGPWLt5OEqJLHlDU5usblZQ1HpyRqLuhQ36FbDp8n5YS0gK6ySbe4SL340rmZMz1DEmLSVwZv
KvCYF1bJ0fQ0VvCbKHsJN4BmKCovzDQH4mtBb42UvCVudqL/BK+iXCYGxCrPbqHDhwrqB0HTVjk2
CqmHaoM/vrwMNoh98GiJOLs4DKCU2VJztQJCL46hhkiPnyLBKE03vfKkZKf0Yg8o48iGrIEknDAx
LI60/9lTbtPLc2tB6Du+g7MDdAxd0l0ewXTacplmmJ9PlRcRJ4GDJh2f9IDb8xos6JfFVCXTKw/I
sYPLZbDNwvTgzXHRHP/eGDj0sTRmnrNxZX0fTm2mmOBwoQvH0LBLnZjorvZ0kn1o3U8Q1jcc4PwQ
cPgUqVQdesX3WNwhWGOiLczXDhU8ZX+TDPnGElXy/o2XVIiNepf5wXY66bgEOMDu6N0cTd3lZy65
4HdPhWex2NX1T8bXEN5eYwtaJ+Yy2P2QeuvQjeSE/+ibWlJnHOKnDOw6OEOiox+sLmtsLsBnuAIC
MHkMHys25i9DQuY88X0FBTUuuExAhoHis5EDUbU/uADnq1IT37xl9FglMYIzXZ2BOH15ZwWOewgP
01FwLaEvCqDwspLkfq5NrhgKRIuhvVmhp8J+BNEhblKIE2TcCNaOXLyvhLac8GARWvNAQEFyl8OC
MIkFBVVbCVnNEMIbVIAlFamOtvcZAfsQfGEkBUwdKQvs1B3b5MceQH8KDbWoG+Cda1EoK8eJz/Rn
bPuSXoPqwEwXHUmGrWB4BNPreJQyxLwNfnkADw5TZJkZm2I6mdVQVij2cDb7IlhgMIplgjjng3ng
wcVqbrAt2R26+4mk/o9O413zYBeeCld100fC4daDRglcJMTfhbBf54sZp+ryriIU5WlXNGfIOqyj
FP+r2crnSCm8ZFfifQOpJ09r54/WfE776v4LaggD5Dy7eOdJRkyXWsvaDyGnlUvMM5HU3zpqd1yr
ikIlO2ADUY6y9rfSwnMra/eQQ685F8BGLYNFEjwgAC89u8YNLjtzmIV/mlQftPVyZBQh/d6afQ1O
6aADWuH+q9E0YIpr/iIlip7ZhXRbfn6qBCU29KCbVI+fCwro5fitQFq2tG2kwPRpuqggj/yfQzIk
R79PJ6e6JzXz9LBULsvaRwf1rGsSeXdKKaQFuo1tc56goeXuoo0fBPq2Lm5cCSEKPbihMVADM7ig
eeBSi8a1Mn4q7w5+hO2OqTOaq30XV0OuRQceZ8WQYIm1c7UxKcQAAWF9WEuZNAvIbWZl6og8IOke
JveBCncZZL8uyILtvMYMD12Bx3BvMfN7MxE+vqZBYx4si8FQsYgDh9UpQ0t26dflnGa7yKU/U9Lr
AYcdkWRnFDfFgPpHcC7egWYXjEsUpORciMw+K6rxGHc8qDOUPyXnzN+jePwtKwWnuZxBEiiUrZbJ
JqhO333K+3IAuCP4z7kIegsr+e7UKgl8fmGLG85aoGqPePFICMy4IviXJ/weUzwO0P/2nmBVz6fR
2najgBiuq77Waf/naHdmtci6AjuS+tPcJgEOc98mOm3lwndXGP5QVtghj+DAtOanuG55TRC9hTq8
j+fEWyNiZVtw0LOVg31IiVGou6AaQufBF7WfIGpLHETKFLN+STADsp9h5r8lMHyoVxyPYnSgm9qM
1V/Td6LwMzaOSVE7dcAuTDCSwUviff3sry5jd9QRdkPIhxS8Z8VTsNYFGj13Y0zfcIqHhnLx4rZy
1Fx6GVx+6rFsseERyRSlWzODOnkR2jM5KHekhC9e32MI36gAI8fJ+SY+mn+FbGTyNK70FaHlHREv
m3YCrhv83/bGVEgzCnLBqNprL/Iz6E/IowR8Eabju8HetFcL/e+Ej2PSUrkGsR/wuNe2Uc9yFKml
jvVkOAr2d6GeBHAFGgVD4l7CrauYJOi2wo4miW5zH/LcMXwG7wmF40tHB+chgpIl9CWY/CutkNRD
WDE/ZeBYW7wfCbt1GH+9dzoLWybRmEQ9d+ZsPEaMYJu7kIUXsn3JhR7P8/piQa34xjYgbZ930C58
JlrUjp06w9ZjTVofs4HwqQGevPlA5JWZ01njJPAkX7gXOQ6ZdzFfX/LUcnUqVHTWmg8QCgYjjpbu
lkPmwFIOX7Os1PrtzNPzSCi0EjZuoT4LZ6A88cekLbCnHVs5gm4ZzXMJUGW5CC0DGJb8k+9tp71n
FcI7n/fG5yTqgNM8DZqVfDhUwfRLKZDkU8Dz1Lsro9glBhCzf9zMVtSjGyjm0+Zwv68bUf0hqCn1
oW5eMZ1Lex2vV7qV713OFHuNQoOeKK7ElQeh8WbyLt+VGwBJWeidO1Lmu+Geia6kfaaGgXn8/cHl
egO5VF9GWFBKsbOy0Eq+yy7TPMkte7nyrP7Y/JIXF6ptfZ9UIIOOs1rRJF2QOmw/qjLv7G6+yi9l
kPOihlMKCjJiKEeQ83+iB6pBjQIYzE9fgI1zNVVsQs56+186lmaZ57MNWhOZbj8dlmkTE5/jjERm
MTSRMoRmzR5zkfDdwI79YVhtDlEwFR/fXN89C1maSxm30HSpdPLTC2JBnK6gWe/xCUIGm9nwTgef
LA2UBiT2QAZeV+ADr4ap1ZbhAk4IKry18JcWIFHiTbL1UalUqJZnr11+FV6O4n+tTc7rMnRZVGCI
AesMj3rrErMxSc10zNmSJhywB2Q8N4U/5JzchkqUDDXXQCGBpeYQZjTePuv9E4EVUft6/xQrLdyX
PLXkIsv1jwWTiY5A4cNjFNBnF7gPhxBtoS9PPwhFh3btCv/xNBDj9VntPAWnfzACFVqYSHPY+lWI
+5oHCNqAJTVQhxb4d2KnJzvxG9kAAgRO3lffWOw4K9Ta+Yla2hFIoNLGtpE8G3gxUr3ut4fxeH9I
Ym73fkv9c9I46WeklE3/l3cmXMz/xayJGw9EIy161NwzsRNMM5Ab4djk6/mWlQGuRCzE4DSVJJmC
r+jPl3eUzvWCBDJbhWAFcJ+9Yw0r1FStfKQygqxlSmM3xmFF+aPwFx8lC54ACs+6akWnwlXn3c2Z
257kYE7inIVz2OibvvXfNgtAByoNOiJ7BWY8JqzyM+FB/2fsxLhcCdmXgriL7L3rG50OnFiTM6Z9
p6YZOhZv4vU/pdIsGSWESkPy+SBOwSSxaKlCMmWJzGcW7KBY2P7VVp5FjqAYxAQND4kDKAxSZkbc
rSMIBR7ivkv+ywbffD2B0b2lEXbSOAueE2sgINQYGGSyG3BZVL+MU4EKGm0IP7nIqCb+HKZO8OwK
sDt73L1lfgeyjUxmhv765WSjwCCGDpR6n+50bK+JWRXKJy5wixsgnhSHBoozCAiENc7KLJ1YPsHL
WiLEGIMBevqL9LnMxlOWTLT7hu233Zl0wg6r9+fBffLawIvUEr3TSE1sWAKOYsajXuJMdRoXaLLo
JKTifvaU41rfK5LdkQcRmoSQg0uGJ/YNOqufVA9BS+YzLgw2iqewAHWFTnz8edmiA/yltoUr3WLZ
23JiR6Ar0dNoNFfZrIq2DFRqiNhPBftQSQQVPpZ4OPpRRaQf0YGZkL/Srwa5JJCZN0D2Qc8D2V4+
QpbSZACacfFmCsS3N1daSzB0/UqAGbJl+qb76IcFkfsBERe8yLb7XfipfMrsKZa7HYmLOt38oe8E
pOu2oJyMgEiAFf4ten6xp6HOn5ogLiXxxBxAJmN8WBZsZwkcwhuoRO01K3DXRi62PzOZJHp5xWJY
D3Q/twd4aYbg9W3m948diPC8XEAppTqTKahGIii0rWRt6zmvlPj5p5ueBvDp+YHXRyWx5FQBNF/i
wqwnaFjPB7nq3yz9Wt0MXspsk2xoZvsR2vvaFm+nNGhgZoQbzyeEDeSuFh+fp3AOGixH8DADKfYl
vHvqYl1Zsb9iq7JslgPVMHAy9WdQ9o1cpmAncG5xYc8tWsFRUdyeQ5vdLM3f20MqNIc2vu5vbymQ
Klbj8GHhvnBBznMBq25lJPZt49HRY4/gJ5RQJ1mh02TPOzYrW1TgysLnysVsJYSY7Dyk5W+nBIZ6
/0sXW/Kw/gJYPRrpZdzpeYLmPuyypa9UES/EKZiLuyjo/AoLBAO25TGWgK6SpIPKhEoU/NRl2rOM
B0AXhAg8cA9iHf/LYi+fHwvkpPx7AZwUMss8Vp8Ulta1W6MypujMj92EtNIM5A9o1pYTETXRazQo
P07jehWG+AhNLVHsrnAD7/ZOyIDok7fFINCCMoI6uQZeyofZf9DBpMBuB8ybciSEmhC7LVVM/5ru
DqXwDyegZn9iyrSdgmtPcXYwQr5fi2oTGK8tiKXA4BKaH4v4j9D0N69tt875+uQkIS6itiN7GUP9
BAmSm1dHEpHZ5sCSwMKvxL/9qY6SbAQaMUpAoIewoL5lx/WgjcNIwRrmbW/oxuSXaGTM3Ff/SiHH
jrGBQrJyJY9oxZUeQzlgDy5ZQPotJFTXHqNSVpJvC18em0Z3z3S1KnSwSb9VjqpLfT+G62xl1nQw
88ygae/iGxWfCMQmMjH7bFk3E9xWDXT53VQoOFwbubDwLloX3OHdRZc/bJuO4q5BeK16qETUM8GZ
cISIoNXOBMHPOxbGF+0A1HJd3EM8fOyn9nfCHEYQJN7thS3SixSLjE+CoozmTiCDROoV3V1i36QL
4npgahM+WlkcJ8hlbNR0HbM77QomUrz0Xxzj06E2aFpAPRngtAtDB4Wm3QybioKLvlFfT/KwppSH
NTV1AftPVOiBuk/B+2zlNv5Hgl+mvaZxDKm/v9/wDwG+Ne2LSTJM6i+iR8AmsIfikBuPqs1rJ04f
bTQfUoAb4YyOx22OuMkaCAr7C4b1kZLPcbF02OJWyvttLcX3n+RmEhTuZhclWNC+Kpuc1e7CGHbr
HWiie4RBqDDUqIRwZcgDwO4R67rlx63JbFfgHtz8kfQvLh8ZDaTBMrdb0OZtimPEQ0XNcmpxYcmz
DzcA60p2sf/xBQ/6QoXBSNfUJrbCmYQZjk5xAtJ/G2iRIAxWKYI2aHMyLlPPyymF17SpPRxOS06E
/0lOSCAR1mVGpRNH2CFc3i3E91uKWZtWjXYolD7q6SH9SGLr3ayQkUxG1nQBSZOI0LuHVAJfOJFk
KaFwNZ47I5+49+c0EE0uRLS+kVXaLa4z18w/vCX7BTkQn9IL8JVCgbgVXg0G3bKegwjQNoGgjuMZ
OgdleMmX6vfIBlo5RjQ+zYyj8PkL1RDNyH9L+q0xbGmRujKEku3Wyw/eE969yUCwr9VDWSogDu8c
9WUeFxxN+MBkVV5q8ZHYvhcvb4TwwiMdH5+6r19htd9Q+Ku43ukA5tQOR8kZDTkcNqLbWoA5OWIz
XerevD80k6wAgvpSVfHm4uiczLaaxIUnhlrr5hjxEy0pL7RCc5q/vXRxDdXvJEyCrJOKVHjvXifp
M+p3H6+v83VQ+DWHIwtjL8CBWupXJCzIc5gTVcj4Wk8VmblG7xzNg2aaln1liSBEqwraL/cLcjgC
ZUotCAYO94ZD6GBY2PloLRTArI9PJRdqy2Bns+JvAGIPATUSQwhdOmMlwXCfwS3y7PQAhhxOHq5n
1w6Ad4utLOKF2j594I0FQuNdivH1CsLm0MnC3wgvdRG44z4eA12RfbOT0g8oYWFMsRG6nUctnv68
iubTQDSFALxPjE+KRW5PUMmR7n3Ie0WpV00FCAWr8Q8N9pkPtd6ozjkozy1ldPIuSiSTaxCqgvx4
EjBtPJ028OiAL+O72+cSNX2/TCFAOsNzh0DrAgJqb8OhjR6H9mHiZoCB14SGZDZ5BAY5asMV0iRx
pFsOuAbgOCuDMwhzivQ8NUQpNmRAr0D9KyW8SJ19n6zcH3q5n/2LpFwe0gSnPv23/nqAvYHUtBfy
IHScMR+HU1pwrgOPURRgxlL7GZAGtJ+SWfX1XuGPSAGeKgz4TUIWos4YhmOmDqvOJbWw9jE7MRM1
MOBAzthFJdx5U32pX+GXkL9hqMTDQ27DBnuonFobh3U08q6ZRO2PvH1rqGicro6Jhj/ZrQtLvco0
smvWRYXCEvKh28+Z6SvfUlzEShbBfzSFqyrFuubzyBNv/ODuotwfInUzM33AP3hVrODDggh3kJ1f
y8NEpOXMhtHrUD4RANbLbntpDmCSJAHka95x7GLSDOzmBZTSxWtap6GznMsI17GuOrn79eJRdjO0
u2LZMvu4jkPF666nlc0ZEM677hU2WbGRY2Ki2ZhDlXFWSf/Fsgv5YZgAB5aVFH6DVBKtpyjAGBDn
D7WUYXN631+En3AWZjBMXQWgsJj79r79e+znAJNSDN9Tr6n3k78S/nN2MKLRKXKf7pgG/bve2Xaz
U6HyoyHCi+IFUcjd8EAeMs6JszZ4iotG4NXZ6AulF0JtXUl6TcQq7ESKdDcV54uOI1DQ5oAjS5Py
vX5el/u1Bj+r/UQjG3kVpFRuVWT0RUHmlpJjEpezMf14qNjk0aWJg84+9p+8WfCTozsULHyrdvQi
k6s2Krt+zkYkx/2G/cUEg3P/qGZxbZ2XEAtwJnWh4rBDfE58D+5vloAkUcADFOGOHM1LOZRx/R2e
glRAiakX+Jd7Jsbq56snPBhFlx2GiRvSfOdZLwuBRRemEZ9SSdC+jwHbv6ftw428IIiAam5mjxbc
K/QlnI6dPMNuCGVS80ws3UMZSuCDpUCuTMoYl9WgUihk7mMDe/mHlfj9KuL6Tgy1n2FO5g3aUD8T
SlA5UaSjmLny9jhClOueboVIuxSCYmZvpvMU3jp4iX/Lb3tmWFs3FUAzYE3+3eb98NaQu2cieiXk
dEiXeCM5Z+Z2CzNx7uz2Yo1Aiz+ZWvtSyGkPltLl2V4RN0ga8wh3xbPlS4pLpnBChStwfldnauir
NvRobuDbjUVVGD1EiDcDguln1E28FxgjT/du7d8VYwsk19I4tLcbqSRa+Ia6yIo2rqTTg7FDW7XY
6CGgW2U+szjZYTJEXBEs2KX3gmsqeT+bELECuXXO4tRaeZJQpRoZDCmWJK3+Jay5fp5gSCL9FmZ7
H8FskOW12Ew+feyhkCq9+CDe5s+Dolw5vZj7iMn80FWUmrfTxngTGNJsV8WKqg7/0UMBgG1FYJ7b
n7cc+3H5tJtjauYW0dAMnxMpoiG2IirNQmbV6wCXzIxEI0apg9asjEIS0bYWnOtBeowB6nR5V/b9
oguJfc1/Cm5tlxL+IXUHUhukShSo2okfbOIpktf6C0JljdK6KSxwb6jGIy9271UtRRSU4YXwD9BA
HiN0/jRH9snfeJuZf5bMqm6pKRPok9gl6i5+YIXxowP1eXyfYX7nXvmbAwG10UzjZdLKSGWm6WzD
8BxwmPoQ4qAQ9QyioqBBmv0DBC+MFUL7z5zd/0EX5uVZEqPAT9ME4ci9ZRNOeLWXlFfIyjO9+0JQ
ZC4GB789x8XouwnavHZmGNxngUQaU+CHYVU9rNRRJWZkzEqxg7keIJkEoc9nfH/tBMUPFf9Gu5XO
1xA9p15RS6GjcJEYPCvMTM1nwQhjC52kGINbsDA9TIeSVk6gfVqtzPRlrDNy5u+xWKa09vC2aK5X
FLcrsS+zFidVQALAIIpLncR4YMoJjaiyNszn0knsyB1TVqcYbhT+1s8gq24sec1J9MNbuMP6net0
sNHFPZnI8mCgG6CHBvSVSWC8kHJZ60KdJWWZfmfI3wKbU8JYbBCn6RIUOBE0acj40AWHc3sp7U6e
LjRNhk9Lqi7vwxCLmMkgNWGVPVrHao1KsgkN7hlkFUi4v1Pb3geWM9redcjb5QqGGrpvyJPw5oKE
Joho8Iomhj7WL6Tc1nmRv3mv2n41BdxGvHFCjq+vqQ9jWGK1QvXcFgWSMrRBMWZndfPpKGEseeyf
JBMrK+rYmh+gUuQozlQA6zaiLE4/m6mak/Tl23yOpLThGRmGYHNYpA9gL3Iz27X39OL+JdfPkOtz
PKreXmEy3jgWCAw/lD4bud8KT9QCq3kr8842RxlMFFLKvjUMEmJKnMYh0DDIMEtNJT3p/vNG43Ub
qXqVH0FIL27gXYV9h6jieMS52ZaGMx5x1DwbweOq+8VE4RNEO3CHRcFVmStczCOtDFna8wIm0Rnk
8RKzhge2wSg7tfn9ZEH4zBIDqGcC8s2/akDSj8ks7yXaYsjMoP/F25m9L0Lfbylhizz2rLBZMjbw
4e5TeJh504+5tYqTyd8uCERoDBaJb7p3I2mmnMaIR78OifO3Zn3mmKRR5aQ4/CQs7Ppeb+CnQMG5
97Viq3XB3sIRQjllYqKVqso9RJfRJGxEd/jFDu/rz9vocLWsWdmVFe3ii2J+8UIsMTWkIBfMIsPq
+eR1HFYVku4wp2klzXFXSEAUCG5z1T+bbCPgWL0xQv/B+S+q2ziBhNcyGjL5IzhFHvZVs4Wt3O20
vulBl5+84vlylnZq3IEA52HdZdHa/b8PFsymu4t9mCyb/fxm8qHlol4wWEP0OMohOXTacEGe9VFE
Ku7L6Jh0JiN7wyknXyoskeWPX7n3VVhbGOYj4HzFgSXtqPAyiXIlK1uMwwb33AegMdqKmUl5gh92
sirF7Fn1tRWSpbI+bNrEA+5N+qmQAyE7bQWlOMMqMhPB7sqwK5TbyKcwGbVa782hh9PDsmJ2LrpP
GdE1LigZeHoIJ26SvyX0MP3ud5CtFxxShWbFanbrbZIu2l7w9Pb6ihbIx25G/M1O2Q/OXdkvs0TW
GlYd59OFy8C47OSFUKSFpLO7j63RYCJPn5cjR1ds5Wj4VcRVhnGhojvbu4jglR7NltoKEwDDsamx
2GFnbW+m4lqqRyX6zJvf/k7cj+u5uhwjofOnljOc/zqcL4XltH4qBLVd8PtLK4eP3gToZFFUWqJd
VkdJtVoaxcRVxJoPrnYvMG5nFRHxEyl24GVRe1FxkZIoai4Y1AzoNDd/ixhTMhg/EmCYnPpbfAAv
wpir5IVF0z7q1+UkkVEFveCmYvrDuiv7sphe+raRwPxDybdyALbdWZSoNLrA9/5pkRBI6NZnAAct
pQjneVKXj3SUC/Iz3peWKQMrM51NpXEHRMcMnM6aXDkmf9jsoszXW+vP1CHkyb4tGUyfhy6Y2Vlk
IkH3qk8oHmPoKBL61QROkcuts2wjQrzI4AondQDrS3K/cXRkH+Yr0DPAytRmGNWXSowXC2o1RBP6
YwmZMUyDtuP7upI4q1oxGBXsH418P/06P96R+38kmKVELHBD1o1RF6uX0hVPjzTn+fhOWEU41lob
LQ0sDjtj9vcOn+s6Mt5eTFPoEi28GRlAFKZGWD8XA1/1lWBC8dP/ACuZY1tzcxvSU/IYDfFx8zTE
PLlkofFx0HaqGz+fR21kg0eeqrSoF3es/P3yVcQGy+vo49sXoSBJF2UhqQ8QvOhqqG8JkJ8kRavc
MoGKIo4IkvnSkhuPGToQCYO/FSRkOt7bASSUUMUK8eWQYdf19aE3qKwT9/fLC7VqaqURXqivutcj
X3hVIWynO3YWxFUDA/pOao4JYs5RHIaJ8faEjqFKi39/IGjBhp6tAWEJxHcJSbG8qOKRDqbr3X8d
T1fGIuQw+Roo+qrc1S30/Y3SMKvm9i1VjstOOXWUHy7TP6KIqoz9lHibWSXyVp52wyg/+HCfaqD2
sKZ7hEKNGTXLWktNyGfQSGBCKSv9IFWzk4FleT9Uiw8DsDQUYk68lPDKV4HzvqiHZA0/y/TxjQvo
1ApCyX1q+bwelqJhAXjjUnahRj9kMCTZEdDJ8tRD2PSzEVEtj2PtKKdRvmSovWt0A8i1NzQm+YXC
vjIbIO2UR+GKBAcydjmSUlYbMRKefgB+siO1RUxR6DQ7xt4WoNefGDky1nDHl9LoKhemX8nz06ax
YIoKUefH/B7PRtWSl2Nt/OmxU1gSyQ09xsoAni/dCPG2iRZmju8rtD356t1kRU1skxUrwuqbR8vm
BuEZJUaQF/pFP2bD9wAyO+zcDmjiEjePnnVuH2VpZ8Jf0PXaW3QwFdauc8AvEaEluue61/cIsq0J
C/WwmMEWUS182SV3CSyGj47wLM0WV9jAMyxfEywzwgXyyq3ouEWvwFjOmm7O60wxD3trozs++VEj
0zBOlsEagXaxE32EopVdkqjulgGVaM+GJdmGKN3U2lDGIhcKW+2yZrCiGHPDK7Xnx0Hj678sJPiS
5DsBT4EIGTaZKD1rA6VoYIGoR8vMCQOMkfnqBJDtoVZ/cK1UcFVdCuc00OksP/vnODwtEjGFxgk1
64G36dHHyswTvzKLxTV//p6SfFMEv9Llv6hQjlQnD29H+90aCA0XPKUDCkCAIKnRgTXenvy6LJY2
tH0Q9ld+08tF18DWejfPBNNtCXPJkfA2YWCnjZp9K/Q97tO0KQik7/W0bHWkAiWOAOCLgEsnlF+n
9ZXrEEQZQxwIyIBVz5nGEHURdPdNvt3eIK0qHs4NDCl1JU65sDnSXt3Ih3VSPlUpVzYXxMdBJgcA
n/MB1TAYefLqiU6dr5evMYioNJJUrMc+8z7nGnKLBBycFYhipxPLcyVau5jx2cZk0DbyjCojg6GH
KqYhqzpO7kzct3HsskGpbr3T2Q/i3QHuCe/abS0PEHRVebQZiOY9xirAKO+cNspQ9yyQR3ngGHhM
tWqr8E8b0L2iGcjFz3/6RifjhecQWwtmHjdtxsZgWdjWsz+rWBBOD4iHPPN36+uwFbwJQGQGjVa7
AqfGPkPQyk0llEyT7mDYDtCHMt6pIAepfAPdiirgInrfRrXgQnC7MpAcFWMf91xORmGTOEWSw4HL
iJawmjepeUbyeKILG+xKKV5WJmC1cKPLkLxcnPqtzgbzLhc66j7J5dK0q3XS7QB0TWA8hZvtOubr
7y5dUyUVMub0KCAvm1wqhYusiLY05eKPT5GDNwsuNNaZtG/OgMK5wKrf/jd/NkCgul6dbU7c1QoU
XCxnpJGbHZBBlM2PzNcHkduIOPpxAV8TpnvgNhkJc65aUkxq7UJ6a6FXmhGaWdicdPNFErxM3qVI
npCtcRU4zqkCYk3OwCQesMtoaapsfAT7rtfDpYGdFO46/rK/Ik9o65f3kf9GQONKGm/ZQ+oWgCgK
6lSAC6PYaKMs3msuxwuz3wmPSBdxxOaSnpVMptXYUAfqlSMQCoWAYfxVaxnaT6q21RCxIbUOYb2f
bbXTnJnRK4CVFHutDJN8bbbom7JEhfuvu3bWvvkTKGZqPGZy/NJwqrMwPcygxLZsxwJcuoq8s1++
CslMYeUDpMLe7mMuMLuXyQF+xWyQ2YEeVVipL41jRw7NLvw6ivJyNbj8ks+eL54q03PpDRDJo0jf
abFrH0RsLn3XYvgKo140OsYOqm+QOWBldpk536RYLvsETeQEVaMl7yIRBlAuwWpq5CGUEs+qVv3H
9HNX63fP7wgPSNAIoxo0Dhj8RnNxo77VIZMj0hX5QIEsAxwoZT3je7/e3Tm7EzGxi+6AwG6UlECk
QSDYiZrv6TyrU5bd1pSjko/PP6vKwAj0M6pg9V7EhmCWuASEBUjsYLF6viwrFNstHCGIwSraeMWQ
hbZKwPoZBvtDh7o8FlY8GAK9Y36TgsVtrnwJu0GlqjyoNgYOsQnEuUCvXD/S/CbYpvht+kvqIWrp
jumL/y94EWtuAQ69/vs6Varu+AxSDrDI4az6qzuuKWyfom4qJe6v57WQpkm3TL8N4oxNHPoz+0lW
jwYaKf2jm9zjL6zNbA5xqV9CfR6+3AfRj925Xu0PclbUYw56o7gPdIMPIdos6DvPtDImDtAd3BMu
+k9h0xsPUltFl7KA9NaBVOxLgMMUHmvAVx5hzeiLej9hbQUQKtGEkQnLaeAKwc2sCKz6R6HG7D9X
wwtDFFeFH2VWT208yISn0IdoNBDmMVO5Dqf+JbVwgbt8i3/IC65Y3bGk3Zs9rGOzkueVftqszoZu
ECXcOIPFw00D7W2lY5oAQk4v1A57z04w7ON5O6xxnt4lft160Dn2KoNoyNoIKuunnVOxLg0AZWdQ
Ez38RCZUCu0BSf2ibYRBAfLYXnZhn8VHW/RowVA7Abd+MHvOEk1hsoWiAlOW747R2p8b3rA4ciJw
KrgcDk8YZ20L1q31gB6h4SMnKCYyF4oadEReNwdG94RSFDbkJHPoEYz5sGpPx+gfmdXbPOvcjO0Y
BTqSZgGHhjMXSl+y5DTuYXNXtad5YkiUfU8ka/r2S7gRXTc+QfIW7Zobi27NXumDe0CjggZTW9qp
cAaBo/iqJM2OUHuAebm8CCvboIXzWMDb8X01s6sg5xfyBXsStIvdPMeyYAQ/u3Og6aMJXT2A77K9
cGnDzypo160F+Kd8Kx/Aeu8U++kwmC3wm7QHQsQvy5xB3aMFoFHsBEM9Gnw4u8ig3qltfj8rV18g
EMKyOB4upU9xdBPE8LT9PJEOrmPTJucKt00HPl7ink84v+KCNKLVEUVzv+aDcSb8dF+ryOXJeYKR
zaUPOyhuSAaOp0rYrdCZqaGGJPIk5Bf8lvE2l6Rz7s6c0J5FQXzR0nl0MaT6+FF0bI2Tfbmvinj3
/VqMeJuKYyls9oTLmf48lRcqaMwXmZG7/7Jp0msrtUuPuWb9KJS7jXkDVe6Kxt38/qHoIgecGmh8
j/GichBwt4CbfSDNxzlNBDeNDMmfCUNFHbIKzddqkXbKwYioCupPqelgN2ktBnn3VpqQShyJiMtL
cgx0Z9dDeeCxfoXYqRSXx0qs2i5pCZ3toTXFSlpqG500UUjH/IoM03r4rwCyVcilQmwHPCNCLW20
MW0WO2irP4+4S6VSUGcBPfDpSG3B1MnujQti1ll24gEAnhTj8sqOb9emIcyu4kpknIZrYSOqhAqv
ldJZmbHuvSzQGiMass85KA+Y4DFc9mjh2fpqGw3bP+lIxbdsmdPaD9FzRqpF3M8B1CVxX2UAR+7Q
uyLULo+WfuDXCfcZwIQ+T36EPxqpuTKBXpt0Ske7z0jCA85mIpeWY9UZHCK5jjxk2G66xrUOZEns
YgEXdqm/pBVn8BI+qMjTddSCm+nnA6FYVhjnyF5ISRzWX7tBugeLY+VOftBrug13OvktyljoQgOQ
/HyqbmubNE9R6g0wi+itjchZesQ0x+2wm7MlMRBwe7JHq/3Zp5uWiv8SVJGPfNVczC/DRGHcvETp
sk6YS7XVlQYqhNRr6M4+7FWXmt7NhBAAlTEnNkTr5vLdFlbaHUESSTYDu3B6Zj4C/eQ3E6kFZE7A
N27GCXAUk1huh6SSuQUsVBB6fTMjrJgcv8F9SVCsoUeHGVBzHck/TcQiK2MJgA9j/CSTUryb35gK
9GfANkHKzmtKx8iNLJOSjSiN/CbmRIEOyL27pB8PEtnSiwrp825VjmN3RcIG1XyE/hJUel+o9Q5O
kW6t1qZOVYpn4xMat7z7OC23VhtGMFgtwYagbapXH2Ll9Bq047Jz+icC+7UqHoXzLAOH/T3QN5hD
dcJTBzZdycu4cDstB/hOCqtIoOnMkb+aSmNv71qnix/1H6BSxEcTfHo1e/ZrrPVlTrBN8v31g2ZE
bX/blBA/y8ZG7fY2/HIVz1iy6c6mysBR5spwANA+f/BmvMRm5+6vgAxYtZWe6UM1iAgYJp9ui8w5
up3JxwjCd2zueslbzhvFW56+oN/BxOj/yUxRXnd+8KFpyJFTrVEVUEji815HpkoIxWb0AAt/5af0
4PeVbfD/U6mzMxwgOZUeVg+JJcJUX9mibDFPC06gwQIcXpAK9dAcDYTrXbcBjJy+0DzKaS8oigF4
913n5zUos0MlTTYkRQXJ/QDB6mjtwtdSe5JivK/y4W7uHhj+jICHR6xfhOGeFGxadFaxgWSjQvpK
QfQCngRghhAMdZD2TvppTQwCh6rkNZjsMbBRbA1NDXMshlYkdiSHQ6sB4A7stMaO/a/8J47gcr+G
29pOOLgYg2C/JzUo9RFVemnOiOS+Kpn8ifr0CFGZ3age97LQgXMfcwB1iucOxIzqBBF7fXavXO36
xpEpv4AKoavnblUlfFgN2bRc0Cb7l3yAD03NLUXdbS+/H6BoydLsi92SeBl85iVbggBJOsWJ855L
cYG56h8nLD5Wl5CI0arf5qdiDA4YBr2H9FHuLBjwMXDU/yX1X5X0ZCdBZYGnLPXjxeRYkPY0qAAJ
I3sivzJVq7KzP6pdHxVrovgZ0DaPeB/nV1h/RA0Nnq7byqhApA6pmgyLKtK/XSYcpzKS289/culA
s/y4UDVQdBk8vLlLPgBqFVGIM6q3kWbeU5Hw4THmJohDCxqumKaZoclPdQLb9KA9PMqvnJ/bXCFY
IENBd8hL+vIwnUVJMQbtCHNNmuHPxuEcLI3KCArkM5W6+yZCr558lu8QZnhwPdQMN+Hg8XLUVwuD
MFEQVb/v7+pI06WRfuzxsCfjXVGioDMGmB6Vlf6ayBvkWux85k/feZ63TETFBcBLhkl58Ufjp7mR
T2+cIK2bP1u3bE1fuCSdmYCTEf2ppmiYWh/l/D5SvgM+isHBGW9LYGOBdNe/wGJsO2DCXcxpDIyn
qm14Wauk5af8CZp/OwIKte6byHq0O2Hm5uPzv8Qivf2oXUyP90qlE3FvrZMwHOS8TWpGbUxiL8pl
iTW5I/0Qvqpgg9Puz+26pWNEFVh3mqpRqFtitlK7N4ywFnB3gW9EjWlcWZPH/f0rF1X2y/kLGB70
uwaPGYrcqUx9TXL7guB4bWKvub6LGbT2MrvYw9/UmN+rqLI7CWYHLspALEYCg2yfZr08vzu6pClD
6zja7iFqjL02cSahupwl9mbysswzK2KvRx2YJ0Kv2EXmtGAO6oic3MDIKlDkWnp35o/KJYo+6mgL
4U7f2Oewm+2J7Z804UFidjOfUDEwcSxpIG9f9inFLXYPEGZz2KSngIi8OCjAWf5tVblhqtaO44Zq
cWEupjMIYQPNtbuXbkyl4g9gTTKCMCSj8ahsQXVYh1bIK0KlcM20Y2frvlnWKgd0C16Ba+BdwSEE
urxDIKHaK3FRYcACJtB1wXzEGbenm0TxWrAzZyrF06j9Uj+HcN7DwUjHQ0qyM3hIoO5zkOvcFeJE
JumPa/KyDndXyM/9EolY3+vVSYA74hjgubDIn64fI0/OVnJylbSbtRskXecDFPZoD3LSaumlkq6R
AyQUqOCAgcyC1MK59RJa2ubaHUXGOX9vzRsHTBYJc6a8AJ15DYFE3k282F3NlwgaGUSD9W0POC5q
mXmBpmb73Q0QyqHW8/Kr44c67k2v6+UeUaXxeRggOO0k+nQViDeTr/UUaJQbnAwcHmubWtWaGOvb
MQQDCGS7KmhkKPfTSoQhU+lo/luaCwWgMxROzcAgSuR/JMtrxnB+beKRVYCCgXRL3QnK0vuhrrau
gw02D0wmiWcHP3IbokmQayDJMWf6Ore4N7n1ZBlP5HLQ7wsJPVclbfSXTAwl4YSXF3Y6NsQervai
4abum/3AnKT2hr1ldj8Sw3DCUxfwpgfs4our+y9dYxUWZfOigA0MfUz/mzckJQwCYJxKBK79c0F/
aWknKxm5JJyPJPW3ZZ71IWyQiUBSY8eetV3Lb5KqDDGeadvHXURZ9xts+7OPp/b8WXR8ECYiPz07
PP0u76Yi0Ph/7wUUuiXxZt0f274lqa3I2Howb1NLbpL2tAy2IrBdsrUr62sgtT5P1vEFAzjbtFtH
+N/VTKYA/G+VR4uZI09CXeiecGNoKNQ4L81+oi8Jc8B39hYQkTVjmaq1YHAnfa22U3QL8yzXY7Y9
+FTshxI4Pnsj+08ATguhihzBTeuZ6Y/c0FBFdfm+02IGX/iJH8YDUM9WQXv1+i/KXtGLZwrTuY3a
lVvy46VbTgPbAmAWblQjj09B4l/m5Waqg2GWzLwFj4NvE3iOi0y4c0InbuPxsBxfaecD5HcG3tFw
xzDHDSnaAwJNkS25Z5qG5zDf3miZvsMKSvLN3WiRcFGHnOZO3HTK66MV+V7NbRB9SqeWYulFTu3q
PfdD0ZN+r0o7LW/knwBPXXZ5d/TSY/uvf8OjLJDSk5ekbhkLlRPxZ0z+5UBQMcw65cqWG6unUDt9
gaHOHEg+odq9QT/TZgkVLdWN5EPAuK8STU6ZrxJLdhDoixWbN0rieodZZHuxK+AmZyJzi88dM2vR
/x88ejj2FWWjKF6zRThlVhMOF4N2ORTjzpygqNCHoJKKaNyXff7OQ4Jn5pTP5XEV/TAeDpU+KvSb
GtXKOwtFAbq53KTDkWY87DrR4/SrXlI2qHRVFTfxvAdh8t8TtM8An1pwkHR8PI2KAS4zR9cuSuPf
omPUCAcqvYIoWdA8q20zOPkU1mQC4gR6shiuhV1QsaLRIOzulQ98xxY3LV/1p+YPoE09KvR/UyaM
8QDQ0xncaviMr8n25ikHdsvNbgOPtChnoe0WoztX/wO4CYee1O93KBBLJZhu88hfPUUWOt+KponT
v/0xQE9IrF8ejhi4my3c1rUT96NUleMwELjU4sNuUR6b4iGVRsnmYt8ml1fx+8rJ69Oit5XViQM/
WzY73syfyfvWkLwuySZHsZfUCVY0bfeKYQl6+v5jKow39NtuzNihhA+riYJ6QLx9Aw6hLtAXuDAT
yTFBSR92PZwXddMnMosF86IDz8Y1nZl/gS+5Urh15GiyCgCpATXr9LKfQnWXBcPgUxM0Ht2yyXMx
Xs30NDFcc7lqxB46U8r4Okpdcng2fFPrncwNRTbxWrxoeT5RKLYR6I9Pl6ROayOGelyqaLVmTeYh
6O71mhjYQRkpwvlufRdEf2J4Y+zH6ZsSrC5d3pu7J88Ju8QxI4mLpOHe8iB8qRVrTzYQGmaMHPbp
fVi7cHeBgHz9DLuBa/vths88qDj39SMVYu3kfLCtm2I0RX17gGlVyUo64wXpEcgNJ/pcshNaqt/H
dC9KUzk8aWN6Lyx0A587A0lJlQBAiasrz8MN5kNf58ltKlo6Ish4agmGwQUrBpVsbj2grVs5pKwf
C8qDPI9LzCkgzdgsnJFHz+wuRkuKNlBbLO/48/EwkyLU/WSWTtNW8VfZ8F7474sQdl3zAE8LxZ8s
Jv+YwOHlUn+RcEV3HxEt4bfDGcsYZy8SaxDhH7Up3n2dDVJZaO+5s4eB/cOKGcKvShcESqwAfENE
mfjsRFm3Gd9dHFpJR4CrTYySIHpIe1vbOiB4y0mlaZJ4hnPdDddYpDBN0vFWFVFwA3ENkune9/Os
e//arjQFRdbfwii2KuXO7TzE4lr/6808CZvLAhvtpuLe7lbyy6roESgiUc67GqBAhjYuEEYgETCZ
vNSqQNNseZ4CERjJJ5SxEN9t4BLKbtv77zR2c0Hy+E+t5kyN58S0rBywO0BTZ1jpZpteumH8OJkl
7UJB4OnEDdcA3SwXQJ/s1aXifqDzWvi0Mtwq34SB0v4VQmV/TTzy2FIZZ49oPyUo/pYE9q2JoJgs
nzvIn28c0mVRGSfusfwWCZ+KL2xfpsMeQihzYDNPyaewcUOhUo63RAvaU1nesdaUIhy1+eUDaqy6
0RyWHjvT+bNJ9XwM2rYPyBCvRG9IbLfcKYHJlHKScxngiZgcaCibV7dnHcsiUrrZgvbeO5zDr+Wm
ZXlSAptOshXp2gGCbhDqv6NiBv38VlkWDZV2rV3Rbf+j3blHdSIWRtHZfvvFJ5X5bUfW8G8iHOrc
fjsAhrMdl63kTp1DJFUQz5vhIKqmF/Fj9VZZxG6oKRPBTk81FT2JriEtXk/jY+OSCTQ1qN9ZzQzb
kyhokTudeN15UKyfYX/E8G/5cDH9wXA+XDkjtYERSODxFdcwkla/D/nqf/XmiR3zN+tfNlNgSwcd
3/G3boxMv+TTQ/XA7IoztHuGm5NZH/x1zKuAQ2NSyOkgbFblHjMHAOXpkrczLUmGWV+nAJkVg3oD
24Vskkoz1r8o9fBo5k/Bp5LLEi60PLGKMLO09kCUJ1tWCPHS7ABQd57V42o9mlURAETh9tKNr7wI
CWsnJtwReyFgfpNiVWc6wcyL2i5nmC1vK8pSTuBLVKBS4XXnfssGZ6Ne5VGC4L8TB+KxsmGPGyut
A9cxGA3fZQVx+6LlY9RKEuDiD7sfu8OjXq6K/ZM7g8qDGrGURuTOuwO1a4T3K+zUQQCv2BqTydur
KFLuLrftUkxHM4ggr2weyAufzt6jx2pL7e5NT67Z4yV+/2WJpa/R3Xl59VMbIlczUhpr9C+6lAA7
sOBw/OUjq5jR4AcYRFma/QYH+MQVZK0f26GcIEo5gJWwgvEy7VlcDMkRWF9fg5CYqGift2dZg+G1
42z24dhWKuQgTm3JABvTZC9A+Oq0txOy17qZxhysirGcn/kZSuQtF3bY5ly8fl84sBiKruyuuCbr
Vj5pRYJZ7/Wms9nl52yK0jD6JbQF0f5c0dC5nxQsT9eDygWE5dWMooWLURzydhlE7s1Y3ikDt1qp
6EMPJbwBtFwMKRabFG5V6GAL7wQW4T7j9C8sMPpYWvnlv3ny+/ZnrA+lkZ+6low548toXlKX6oww
uPLhIePn3XDGhvWlLJBNpuDlOiyaO75ezLWLx3uzu609mMctjsGljZQf48yPwRRKqI5KoZwPjOH4
8R8TULP6HF1WxXH+RDPaqc+9j4yXlIDk/DXl4hFzt3yLL0jDXJRb8SZYav92pcCGiwaRqJrfbG1T
SlycolNuc/azlO5fEryo08abdoVfdB/CNttLO2sAz23yO1DwAsVRH36U9q0ykNzK4QjO/SqQL4Vv
jop4ipM1h4GIJ18lkeaiZznO0RgQ5JZofZMN8OwLF5aCkdUJkHsA7oAoZtiE/1Nj+QQQMSK3r8Xc
tw/fE/SIhMqIB3UyX2EVHmj2AGq+qN4GJZy9uOJvdXPn04meZVHTdUXDtj1dJ/dhxA2QVEOJmu+C
EiBAPWObcZTLZSfUukaBIbxGJU755Lqo/CidmwCC3ZZUiqNxVwt5Pxz59Ulg3sL8vsk+QyjZAsGb
NLkG86r2BF1bdebet0HWqtvfItd3r0JB6S7WPTSSvsuA+VrldqourSgECgWU4uCZllfvP/NmQuVd
STNaYj65NZ++m5jtEsNF/pxF/0i9PQqALePm7RdGk3HmDwRLrx+kM0VYQ0GPfQmI34REiundx7ON
BQpOxtCtq13IFx1vJ93JBQfm8zyV8fPx4k50okdHQQyBvkjdFREnFx6g0j8fDOMWeA3d46tJrB1s
vTbdD7wSDfALbkhbow528TH/wHE5oG1ZDY63+jXJPT64SBdf7o9nAy1to7ikVobvzGW33l2cN7TZ
iOSD1duT/sVv7aQKCNdzuTageTe4kjGhDZTX8kKamHbDx8VE6OZkl9uWjr0S6rtCcjFU6PDx3KMv
l4Ci/JQWTVbpEMQnkFgoD5qxIm/oA8gwBG4fbAZQApsufapgDOCVKnf6plDBtdBILs2yhUL1RNIg
Yu1i+w+PmBwV/C7P3n7Q2/5dJgj+VsDc9TEwocidZpXPVT7AW+CpEOcm7YHm7uHX6mJZysXbWZ6d
YlLqHw+pt5GcxwZMD+6tHvwQdFW1YeZIZPl6s/pCd1v3Pqvnkw6J3hZNGeuVkZOOoquaaWX9I27f
iPHzOJOSS5cf7rbrRv6t4bc8/y6bDHHSbD7kEkpY5yoUX3Sqtk0m+YOqaYHRbazAl0tByREAcSuk
0NcPnbD/ICt58GY6BCOQwN819sVvTxdOtx1fKuk3qDHqSvMnCnA/hUQ7N00+P9zT6G7Q69EgOhKf
3Mg6s2Y+RLo2eEQdlnxvv1zsHsOC6bvruOeOFPLzvkfg1bp6izGsvhFh44MHtjmqtQFc3p5NNWnB
C3TbMtxEiNxCQys2am70iD5Yig5AZEencMTubP3yFA63gN4XegI2BLrnGYF7U6PDr8BSBAvRuC9S
Y51U+rGpZVLVN4KdcdBJYQnaFgI6CCLuJlRO11QksgHgHcpoDgzVZHiiCsjayOrFHQTGJDJ5igd3
rO98sJAMBBxHIzGzkf+BFivcaJO/xaxbG0o+AWZ7btx5jvVM/N4xe3xFLrfvZLidrqmoKq60vlJB
Fp5Yg69nAwc56zif7I8GVEeC/S4TxQ9gon+Vit6aVvjYDm0h/0NFdb+c5KK6p3yGdLTDzucdVdCK
Jcv/fXIldKS8Gj6RRt+f8e2Es+P9rmDeIZk+MLc12S+05LDvqbDipnRhFJfvmiGDq9xrM+uiYP0G
Zy3/56yRXQQE9j2wy/qxJCvZlQgEfuUoeQmVdAldKXs1C3krPiYMjntynSk2j6PRsS4tq1I7iGf/
ZZN6WeUKnBK3uIarrxu3ORwq3zSoZN78gU216J+w7+6MHVCYd6X1sN0jgq5Q2GUu0ujNiKFAxzLf
yFks1KvkMfRSKJrTahat5IxvyKARQZUBeXQq8xwOf8keb7UHeZr5brEG85fQ+SzQcZ82oUYw3PY/
KFBhi9HFbdU5n9K0BQU923hjp7O32iKQHEJecOpM3OvTgUNPatl354b6QuICCLQxJ3p7pFQhADQI
ux1AxweN7L5/u8ct/gRF2a4Z6oPttLB4bGKymVOUKHH/Zxd6YlJvF2f+gzin+qUO6F0Go0Jschrm
UuVnDOW1SxlebZgiYCRpU/lQbOqXMTTWsmWsT/HsuxZR0p7g/JSTXvDjZSPnbnwqtL1AwY6r4LTu
BzcdG39oTKxzUVEbG40vTHa505Ed6XyS1LkNdzu5+scApYqiL7qNNBYvXxEtiOtr8bua58BXIIQI
MB+AYgF4CBR5w9kSjPv83QdjsM2cC5S9Fps9ipdxC7w1u3XH306fqU/nNaiQRQUrHhJkzd/uN1MN
A1oeL9oUpuannYZftOTXRmg7dQp1HFU0trIXGfDBM+qSCkUY9QLX2slFm8UBVw+f3KQcyzEhocW0
V15RykBZVWyci/0OG34/BRAT9rlaE+5fBcqh9+AIEw/rWFp9rvUQ/YdNLTB3NXNoJmPiw/jVoTCh
k6vHALBNLYPmAzBP7YVtxDKgOBDrtHa4BPbe2CvWxRnWQjRLrLCmvZIxRfsTg5Tfw8CsfLyByCjS
k1EpZvV/L5sLr6D9eQWUc21iV75zx+ovV4ELueWkJH0FifoZ2cBsFpVbJL6SSuaJeMws8FTEEWV3
o/enXQjTL/K5Zd7LjipHKx6NHNqWotwu1R9h+vI2/4zKojUuxTtiJswSx0h6epekm2LFeMZbzaTF
G49WVHl8mBv0SXhsqyaEOp1yJiL35A6jlbRAvqgf6XFM2X3MnawHfdZhgxHnafMbtOIBe9tFdIzq
vqBvU6zOnXJcRJWVIJr8LBblwCFIRiwAcwhxF+YGmN1/wemmn3cn3tTJJslVG3njfg2Zp6MGoOZI
lMn2ji56thPTaNrmjzVY8XaYhTGxWJghqSP0ap+TtQienj9x3CcanCF0dmof2ke4OdAlbIspyBzX
Mv4pULL3Oa6Lr9HGQFr7mk9g4J+JYZZ8wCCCl2ii/ti1xhrxR6EVVcwazEcgqE34kRKS0WrQRPH4
0/8LkRRytwcGqg/HBcGtOolDqH38NKjBsmkZj83s3AEeSzGsvpALF0Z/FBQ3hmZTO77faEPOTRfB
L481dn8nrkjGBJ/2LLvyq1Fdu5Ou00lPRA0qzI7SZqeE0zd0jNwVJHAQJ/+laAlIGBERfJRmTYOj
Qp0Lgh8vhhwRT6TooFW1wMYFYLQLSI3TF2bRTCmBXwMmZpA3CM/OWillK9LhdfCfTG4TkIGUEEIl
rK172H0Ly4c5VgX4+esN6Lj3R5QSTVD8JviNtOENzUnEYzY/OK2/ffLmsHrBVRySDL1lyst/f9+c
+d/04V5JtAKHilYXTyLrWkgW/AQwxeLBRwhDZt7Slo7CdCpxO+g2eA31CBpw7AQLLb/aC7u6ODQU
H3i/4DmFlVfhGgM37UDfP99ey1Nml0G0nd3mhtCWsfw8LVgE/5Ctw0NhNqFa+aew8iqcJRVdX30J
AiuS9buTQA+oOFIZWDgRfXLqzSO+M74k+yeGxDBW4HZz0s8I7675ZUtxbBqhkBNMpEuDeKPQI57I
OwhReimzx69qE5nFh8DFu9Ept/GHI6T49XV+PnNtGtjyz2fKF58nlpDm4gKyZz81Jvh3ij5DFfA/
5UaiGV+hKpxmqs9QpkkCunhRBWXZzt/AtyH1nfta448zwGF6HhpmGrvdMiKX/hMPS6Jda9Dw4SkH
prstSUlVxiXSB43OkujgiqM1shkhmLfgm/19goH5mvvxdbEpyE+epsl7inwIRLbgiFmL3CG47o9b
lsvYDY42u5NkH9RxkqCDajUwqMJIqKZ7fUlHDqIl3GEemaMcQ3CHSiGvAWclL0G3K8iOedRCoAOy
1+W7gbKHoKTutzOmvO+ii41r5GKkS8sniEPmRquhe+AYYGbHLqmBC6GNNHeZbGIIZ2y8QmCohmKP
i3ClSRdyMe3VMGrbBY5oUeM6vE6Hkl89QbXtBQu8u6/O9txVlaz0/QkiXsb8uyue1CuVAB2pA6gr
7BJaNEMNDiS4EE2SQEADSpyal69T0Lg0lhrLpImh0PIwgpOBUIrTeP5YAh3RR4332Y6vYf2ei+PW
6lZ6E3mmqSnZgPOixrz5dv6ZznQ1W4bmfn2LLC2AHA1ye2f4zsXMhsE+0PM4aizw30+s73XzTywn
HHaFwz0oXs60ldqdxMfKUJdbBn+gDsIVMFjS8x1Hlj0phJZkQkXnCdzn2Q2sXcoLry/UjuL0pAZu
Nr6+1cAl5lvTklVzDKWZn2fUET+i4kUSN0YvLRgYPP05/LkebxmkfcEJIZwXJgN89CqdgnJgGJyf
GOhm6iplAE2aCZJtZnZxUGau/4imt9dVqe+81/DjndjagbxgHlR8J7+miuhmZ0qquCN7xD/ndak7
WCFoyaE353UKi873Nhyfrg33v2rawZEmascK7q2+165FbrIuoGv5kj4pvLAxIFyMBbBwmw5JYu8b
kgvEkDfYrAw4+wKdHbmCkZsNtTRkjRrwaSKz95p8AfbgElDbXl06FrlrYHfhM0LvcGwd4+Vh+d+9
lLJgpWsKp+elGQ6H1nwabMJf/ePFpusSEUgcQL9OZ/LMr1DNAZ4OjR1Clu4QcuB0VxRsZzzEZycM
Jzflx8wcPW/b3BolX3cwrbadKvv+6eWxU2sBVxAAiCCngxYe4dFJr74qCEKigmryQejAad5PKw7X
jJCpRtHAEMwQIKGbwowAGNWrulkOVH8Hbk37+Cws6caNEHuHRBsdMEdPoxEXIfZz5d9mt7S26K56
B8ALiwuvuiym7Ha1NTPcV+nMESmoEfVn2riv5sa2nvCtOVUy3H++qtWHfEqBg1X9UhQbaGSmcdRL
g6EFDMxmaeAr422Gbt0fSBAJXrLjQkbV3+LNEiFPzmseDw1YEfzRdz19v8rq2mwFi74VU7SjGTyi
XGnqx2x1VsuBSwHztJcDTXqS4CR4RPmkk5pAfJ39rLB38jbomFlyiJvfVQrjEA3YXB5i9PYCDKqk
8U0wVwBDwVZStLbKWVU6ykkPrRaOwfMMQE/dohvv0gzDJ41TZf72yPvJhizMohMrJImhrmkkSdKR
fsufBLlZwc+cm9MNcnVYikyTabjcaedJ+NBKlTGKS1uu4lQ46JJE/jWRS/356t3OQavV7C+Q6GwN
wRvgZWFhpz8rlMBCa13ngP18U51SXcm1NAfZTNNd3+A7EeOih8MplExoK5gkfaqUylCm/Iapl9dY
wEnbn5QTR14ZwztHghFIQLeA77Qtujgy9Pz7mdHng/GRhGYwG6JNx/WJfKqW09joyz0wxoEAwVxd
f1Rc6bBnabNusPF8/Gg30vbvuGvLdF17CAaitMLQaoDFMTm6Rkulltixc47rWBTZ7YzvaCM3vXQY
sw/nNIbW1oruLWkRSx9qatsNBc2yniENzSMavu+OOz58LY41ih3AKo+cBvoGTgZkhMvxAT3mVP77
ZaydnFIs/x7BJrzB5JOffVZbtSbBgqDiaKvU5tlLfyfAU02OBlStUKP+rZ2qlzN3RBmII7Ek0l2b
OUGwylk1KdZvlLHrVseiY22whn/e+Xq55bJ38EBrPSwF84+UamsB/NQHa2nHz9DSvjpOwnXuw+1F
rVn6a5FlfzL8r3gFnB+LlYaGgJ5s6g6fTaLti01p28xmpHmYC0HzgGbUgGa+9k3X07QwUIlbe90W
GPVEDJDKMchcRWFKrQRLtEJnWYU65L40aedAQYtUJmllaCDi2E+0RNPhCVwMicSaP7Yw5DSUMmNF
ql+0xnpQG1R9bPBhTmGsvPrwp53IqPrJ3JFVyqiEIaMl/yXDGTsy9tZ5VGyolU0OX9+bjFO+v53y
tzBuLMWKXPj/Pc4RzpTYJsOaXbDLw2d0QOvSJsWFc4Bq4TMXKTRdXPowY4UbOLSZpJwa4MVU1qCe
pDwnEnDLYby01eK7EZzuVLvn/cr0SDbaOz9RnHDL0pQxHse4jdgdl0PBckWO+ShWVSt3EaJQZ7j5
We4/LwiZ+ArK1d3JQoMcYLyZDUUkmU0wqtL5FBWcmDksL8s48iieOMdJ2AsFeyHVGo990g2o/oyR
ULxoaplnM3LDZm/n7iNWJCXDOtBTKVaGOLI4kJs2hh64QmC0lRgECgIdAer1YwEtbO57AgAZRCMS
BBtWT4WVIGWolIC1xy75P7fY/BK9iHfNAjmDbl6ji9H2WbtFQs8Vitdj56s+2vA2QOMgVeyehCao
MLkzeF9ZcZlXAB2eOZKcFroVA5xsGsa0PZVhmJgKs6CcecLt5tq2RXBDwnCnZpITOOn2mtXR2E7j
N0qFnu0v1Pk3LawQTRc/kLi7Wgz20B4N8BctUZv4PprAEjRXqrN9LktVhl7+7m5hZdl7zl2q60rK
QLoMqLI1Cf4fv6tMl3BZaF9mzS7CkCjM1NJumYf8mRed5UOsJIi3LX29ZQ+GEOw0VKAKC2DuXCSg
Wr/mkPTNOVIX7h5ORyqvm/7urPT4poom4Zf4eYAZJwBez+YvmTHIsKd0heaSY54qp0qsTdCnJ/4V
VGxqos4tMWEERvasF0lFDHLMu8lfFw+zYRoTbMvU9NQhOJAm9WM9GfEpP4pUsm2noFwBz0/ir8KV
wrfggU57O0xBLXExAV1Eg5pjqA1DhrUWkPDogHb92uuRE5K6tP4tY1u0Ph+3XNOjEeCNBtr2aW63
NcCbe+01TV2BuSc9jySy6FsU9NGrfLHTJK2c/Y/wa7O/MVGVzILcyd2Rl81jGzNSK2xWWoAWZWvU
55vmQ8OcDG1XvNHaNZmK0Zj+iTbOAKt3tEVGAddeRnnBITA6QjUfkDGOqXG1EdYOFo4ivHB8/IOJ
87Fof8HSvYyJy/AupR3fY4zjJNvChvXEkZcUcVUrcmXugrpHqOrP2QJUVPGYwdCjRGgpXJ62BWkl
sssujzmpQlwS1nx0zvsJuX3Hu4HaUh+xxTFFxHhryGc7QiBCMWuofQ8AnenaQxzn7gJjuj8RV+Pn
PIlBd7TO2QvLRSEntqaTkFEOjG7ubKTwl5XUvZjHIwK5ewfK5nZ4P4xdpv0olVsOErtTJEDV1u3D
OPYOiWddJBLCuL6W68Zc+SR3PzuQq3+SATC0j4lktrvSzSKJl1k75lGCo/owKOKKbY4pOWkiRy+z
gJ/0u5lebTg6idbCnD0SDHI2NVShFYNDMY1Jj6eoyf+OzzFyhM0q8hlaN3CIjaufsiNmPZzjYJvS
vrSnl94oZ69+NmFxernG1QJ5AT551DC3H3wH+/nAK/ZeMAKKBCwom9v7NQXqYTpg0GirDt3vAMGU
cxFA2qVCPX60y6hLT1CqwD20msYe2WERF3pBiUDgNlJ6NVUNy6+jSq8NWMWfwPFZoc/CtMS9o2LO
ouAEJmKb+noBrJdmjNE3WfTm/ChS8wTxXsYm8u2xG7vZWkvg2GQuibhZsvKEDaU0bMqvSVz+EiKV
BsZK5LqHI1M6B68zA4XrnjppphQ+w1vP5QqScRgzhF10uN1IufpanyuYcN93SoKCa4nEjHBA5jqq
Q9y3U4HHKoba/Uavbkx+LsorbOC90NNooN94OmNnrrt9wZkrhFgV/pV0/m5G80szodgglpsSUeSw
B7IdjXai0C0wXFK+PKTfMPYg+Pc02xvPEcJAA4onNI9DPzRG/rfQ56p9JZFtla0UKLeP2A0cSJAP
i4S8aEZdi0MoEE6rLfMkXSWzCGe2Yp96QhatZVqQlckiIZDL2iOQRaav0lGYUvo90DLGBMjBuiSk
whP2pQ2yV1tzxOWCzAAW8IZeqSrJdWhHA8fSWCOyXCDlwENfTRVMyjKecbmmNB6KBaijqXbMBjnS
zDoWGEj9A4SL6onKqozJdLWHkCEQa6RkWeV7mDPjtbT2+5p/8iJ1dxFP9uDchaiOusuT1fus5OkC
PdL+et3pf77rGCPRov/ympMFZlsT0hUo72IW24NfokQ11PH5GMPm1W7M4XPXi4WoOR9SjLtpPFD9
sXIDlz13Cp1P+oSH7GDpkMDJnBjmruOTofwee0nMOpYIQ7w+Iu8m9D7sIvoSrH8pLRw0rp/j44dA
hdkn4H61GjxDzfZ6uRqX5K/Y57IU3kiXqSg27OYgs1xV4XXIr6kwuPDn5IB0jPQN/jjfJaxW/PhG
s6A9U3y5t5+9wy0Sivq6WHekrxns1ykQ3DQkbpPoTsv+RDXnzdiH22GIVD1hKTdic8i999WODC3+
YP0K55OmPUZ6SM13QnnUxpYXyjx7UzShEMU9HScj/3sd9aCk3xJOMgcEAk9OaGM/nYNssswHdeR1
ag3lR8TPZ3dBagRs32HaZ3Vh4iUZ/MEXaIBl2hgbL6flRnYPuntwJKLMaLQrYZRBnAl09eVNw8he
Yt/i4auoqbk7A/ub7ijHv+aCOkcg0ByN+jIF71EgpNzdxorcVsAfvbt0dDhhn0Tv4jw0NDb8+chw
FB8X0Fx1ffowbztgthW01Xr8RE7RQJ0fevXjA4xMi6Pg0gUz9BIzEAFbK7EAv7s+1mbGazBsGjyn
78QT03AmtIeuaac9pZSRhSpOCgVdfRra1QMoJAx0cyMWy2e75eFMP9yJOJyDaM8BYxvoDdGA6J1g
Lh/SOnJHkCszOoNac+yFu5JxFeFbfkUN4WX+fO/kJQiVqFtI/GmjT1V8mEjkYrBTNWTFr342asiI
5tUa3TX5SaYYEC5PQlhgIVveQoWyUZYJ1N5kKr4wjiKMVAA/7KPxKCF3N4BZ0Ohm2bhSFRkasH2i
8UztTkzHFRDu6HSrsFntra8oCjdAKnE2eaH5tqI9O5ptOMcNcWNRmnnIRmYoGkYf+iiVwmqzveAa
BXlQXsbyxlTsSHkvgiGpmAg6KiCk09EiCobFmisP6ivRf1/ySfvCkE7fl8nM0kFeU6se70s6g1NC
Ywff1ZfwLfVcStkqYB1HJZ3p2jERaTL6b4VyEUyJkGOGuOgcTEkfyOf1Jw3DlFHgcdbjoBJ14zl0
sCjRHW+bsRj5ePIpoUHpECm7s2wv+o9HefAm6KzFek5shSR2PpV/qMusGb5qsJaHSWRI+CCRthoJ
dOaopq2+8yyK1gvWEx2AIdzr6kHl+cRqG31KCYo9qxJKNRe2VbEHCBQGC+wUNRUe9YAK69y/vxfH
c75bkFSvn3LXY4fGpfAC5h9ieXh+/2KciA9/GBiw10Ac54xkRNv2Nfp+Q96PryisbgxuMaePGctN
DIDQ3CNvvnyeEHIKcKYJcYXuHzmgvW2EeJunRtBrgRu9cS5GTtqvr1XyhhyErh8i0M0S0YMJetcP
qaQAYCp8VzqWfpUSh/C1Nx8FvISwBOoeUb8L/7fCJKEOKafOWY0eFB2cFYM2LHNmpUIebfrbGbcn
Uzzsl+aFc9DfLMjgAInSWmTxL2yFZ7XkuxJB3VPUKpyMmfL1MKVkVzN5f7MvvrP+Biq3Sub+HF8U
k/imxR+OW/Fj6A3lSZZ9mI4wa8FZVjbi6Y+87jiXdz1p2sRIMDF/JMY329+UoEPRbLTsDgr+4jxa
coydPtc6dnXNZn44bSNqtiEhAvWv3KqlU7VT4dUZPLydsKAr1G+3WUmV+HbfQzGCH07oQtIbdyd6
Tv9rFPa6aZyeXMg1oSEUjE+2uTmXDCCsHlLbVH+sW9lBHCpTQ7nCq9zLohBEljdZ6EaTpkQCeQuG
f5nD6PVdzTjsslxT6/iEiHQgqaqCZN30VrbUTjYzNKSBAEnA/EYwl67+sM2kz1dlAZgEtkX1z/Cx
pURAinhB9DAIeZVQ8UL1Ga0vQAzjpzLIC+sPUFRQCWc1V8gBx2kHMdNH9EdKkLf6pZ8vrtQ+anHt
ttl0hrDkDlByfUK5M4/PCVDXoGmfANR1F5kyJ/15aA/eJxYU5q2s/Ybh3FXMjzB6MF74DUR71tco
cotTsYYGIBdr8bqdvy442y8omCgri4OyTCOt8BslHNd9s874Tny3s6dVowCDIuzKaqr33n66ZCuu
6yqZ06SnZBazNn3J3Fhav24Uo6jdwc4LhtgwaP/+7ZvELqYtZa0pzaOQSPvUfV2bVaU8wR6WMOIS
SDh+ta1DZoNLtgDv2lU7sPVQT7bVCF29CT7w+MjBPgsplQeA075VEJVw2mtFeqDqQagYALjxNyhP
ZGZi+H2FW5B16MhiEDUk1H4yCjOBg8pObFDWySt9fUNgOetla2iLFRG4WV3BEbRNruOtlkVV0Crn
mRrgAXQuZMokUPw0+iyeq4/+S+IGiXKj8ce7uK52iKwI3R1DNw+35Z1EEJQbcf7+f6YzX5Wk5G+J
jYCHn2x+3W2zhQo6gzXp61JWbJehoXD8sNDXhmpCNxLbiCzka3NxUFOz2TY6Vq/bOdOov8dOM3Df
Mbt8h+hlwC2zFIt+t6Ncgo/5aPfl3hxUdWxZH8pcAbGvVI6ZPp1yrqR8b5rPuVtzn1Z1R1jp6SJr
26bMrF0M+UGqoLGAhnH6KWeGOoA62WU2qO5u/eMPJer/eAa9uSEVd4TFVz9FLSVly1hZS/GuyMEN
oUneiuEpAnRXgDS7pfL8xe8I68kvRaCBeoenIAc4reYCa6gkcd36tZyultNnWKfn9+Omv73EAM9i
204kGqRKIPlbaS8i0OHF+NYqEthxIpJGAmXeUagj/j2JLpndmJpqvaFRdE+SUVPxeRdDPiuvCDKq
vAIFcVp+gfipBOqi2kq0JbnBT6yvsHmZkM9/3HcEyH00E4d/p1Lo02h8JrF6aACK37dMlUN3mx5u
t5GHzNYMz6G5VGBfUidZiVeKcs1fJj7O728vFwfPC7UxCNVnhyfVxkkG3kvofSOohCqIBR6dFPo+
XJTIfWTVfjNh/ObAkGU7uO5wHFxyeqXo6+kWKLSpKTXlxIxqBKu71K9Mup4TvqEvoQhgghZv1iOp
3TXuNtm1oLexpyOeTIqxWEleoiPML/sV2Il9Xz9R05/7gxHnFHtd1lvKPJFRQJN5qV4RgQs/xo9u
1IWur9cF7SuGkxfFxZrM9vwsfUvyqQm+DUKxp+4mX5iflv2cuvYlpCTxB0hutqbdGBXnWOgreyeW
sLtS2U/3DnR1ES9YALGr7FIgNoL1AWyuAqVxrQuX275vdp5dgE+bkIrmuG04vnFMZHMDQckMfCCY
0zxzx8JRqKlrStQByAOsNPjrHQ/wPxWP8+rXaa7SzW3jIaZmIRcTYG4phF234dCN/qz02bxBa+kP
ah317dGQfGLhW88TyeCZU0Cfk/xVoWPFXHqQWWfxkj9ZO56Naaf4W5ZZVyx6Kpj4xb+QgbLNDGJl
li1egTT1Edx/cewAmqEDInPIIrCcuDC696+YnF+Y1tuc2u6fyWeFNcMhPFATe+HmOa2Cz1zbjheB
86sKr2vMmZr2t+hpgdt9zPKVmKzjqnGOHeCm1Ia1sQnqe8/AgEYXEGqT/cAsV6EOtKuOi8CKxiPi
vh9dnEw7bWKwSEZW1kFnm+p7LGVzarAokUUCoxZxjmNiagBw6c5f3ArxhHL6umcstJtU+onDOIB9
X29axZ9D3BfA4oTOhkWO0Dew1LlD9h8GyT5hCR4x0gzaBnkA2a/LV5JKUl0uUYmE9RGTJnNCo8kB
xXzRMneGKevtDoRr73SK/MIaL8r8WsJmxQyDeEyy5kvTuWZNitKmPi6rPDxw8lvc59nc7TwYSlyn
RIMEIfE2c5RiwDivz8pO6f59WlzFLEq8wqhal1cif/CixJhSHX/X36Dem9citqX15AGiSDsjjlSf
prnmmiBNI0iS5CH38mtj6D7gy+gp3NnrbLLIXOKD328BoQNGrbg5ZJReeODeKJhJvhHd4bmL/d4F
LrHW/diX4r6Z4YIE8/mW19j3LNSIzbafmBjmEam2YdWX+X++V3EX9U5xcOElblH7AwqqgciGh5nl
ba3Y3vygFczZomTh9OB2PAWr34m7qj1n0L2xV6TKLYgVMc+m36gSO5/107mb6Bc6mNl1yyj6bRjt
zLg2+ViVbT3pst/YiLVWACDSX1gWQ+UWuhU8aZk5jLs0SA+UCYZN/av5EYrfT1Z2J9i1Xp8WwjT/
v2VI4jJfohgJ0vTD8TyHQ94UsTd9H00uNri62/6dAQtOgyMI1/Y2NkzOuv7OfO7RTfTUUVH4ij6m
8/wm6igFZptuqfEfS7ZJPeuviPfQ4U+6syr1hcocNmtw4Iv1oHcjM46gBntkWkbcSMFkzCQnrwJ6
w8/nDzXzygBYUMNMG/LLQBzlyYa7OqAXDfQRKBHtU9bPmnmoYYk7CpD1aoDe6DZ6c4VwkCP9UJDw
wgpEHBO6QwvUpLOlSm3D3JXmQTSlILTjTEiddaksK4YYRX4rxuxSnLtyNIeSjzMa3EF+ZLB25Kam
wXOzebS2+Xaytdd3cIuFx9uPEwmqlmZiEdegp6aPOck72BhK+87YwKzg/aj4/+01oWTaXoaGL4fp
VMStSgc10gVyd9orbPoBcxSiIROPlMRd6yAoLeccRqUS1rlB5ZAqHHrXo9GKrS3mRnPWLTmnEJxz
5sMC17Z1XoX5ACpO973u1/NXIdzrrdxuxnm4DKzO/tQ5G0Y3JiY1NyBFpqC02fWpMBSMUdkDZnnH
zcmKofxjOD3hYwRFMWq2DDOaetyJkEl+61uIq63fe+aMozDy2jhAALT5xbgCYA71NvzWJbG5WJse
H5df0GX3B+XEHat2x3wQa8Mu2fih/GXD6vsezUW+InNMX1ajdIof9cwIKD9lnp8HtU4yZegDT9Uy
IB1Nd74oCSXslMHgK9Sslh3DdsSdIyH0jEVXeVVEYKVXcMimLVMcnVtq7WTVKUrLVq3U5NT7/aeT
YJ0WEBwix6UgjjKOJ55DM/OEgbymTY6NdtCmSZ58uOBsaJwhmB+9bMfSnJlONICu7jPJG+zF2/1A
td2uD9ooTWsYs4cD8MIx4UrWOPYxRwl2UVE+5YjYPJwkMRGJKDyg4F9ZnbZhqcVfA8TKIba06R+p
hqU3d+O6fY18bR05zMYY6y8W+2+DNslpA562l3iqJ49MsCJ/3MkgmUhoXQxgzaOvlP+POfDxCHV+
3KTko6ZnPJ49lSWJe05gKh2iBaoQC+jAkSpQJ0yw8cwPMaHgoiCwdV/Y1dW/OUSJp6DIAAO8TtZt
678WNTAEmxFr451AW/pZhOIpNTWjcQ8uhtYSu89f5TaLUg7KbKjfW7i4/XXJOkDmmsWstJCTlyQ4
hyw/FX3RrIYWpIbYcplx90iseIYTAoXE905/+LJp9X/V1AgPt/u0cV0EZJsgrrs7RLTb4DGLwxNJ
bb/KRU57Xg3TkruwpLFTHc/d0mjrXjP5eg8hf9g33YhBcch6q3fomKOElIwcckFf5UVPJ5RT3qBL
4/NSHpXKXseu2HoDLbvKcugyO7FLbaaDBsVnZqX1tH8KlQYTB+XmJXuCHBrsIBmzTuT5Gekcw408
I3PuAQNCK7yU/WITk6ItV16qCH73XycGLR7z1Xc/J6dbh3+stEUII5TeKuP0iXpGqj/+aVR5UvT8
LuhiQ+XoFocTLI+N9SdBvqtJH8RCGoRRWIAaCRZZHv742VDr4eMeoRgDfJoIKpIbBCN3S/XYWlah
AOam0pG8SDlX6Q+FBmWm82QuJeSoRxoNXl+q5UpoKpl0cJIuOsT0gGdUIdnRXE3iB2j9LIYzjrvh
1p9BEnYSAdxQ9K4XfJG8Qf77vOzq2vwvswmWYPRpdPxj/5lMg2Y8Ih0UN3ffYMPCC309RVDR77cw
C72bsWx3+wM1TkxwMsQx3LHXUy3CmdDk3wN+7SE3JI3hBtGehK2vHMXSPVOpA82IcL0aqyLIyQXZ
XZSzhsFs+78TqRO9J6355zahrhfsU2OKHq5oypHDLNyDlJ5FsMqPaU9TUUFXHhThR77MKaYLU0U7
aV+JDENBe9+lvUYH2whNOw9Kaml98W5kyK0WnXpLs7LF1P+MmMFnbDF5gM1D04e2JQWhWa3aDkSP
A7oPgt7mpc5NFcNQATIppklyRShmpuo87HJqOJji+8vFOOTzNmEGsIdTeLtM8rzdn2vjW05LiRIb
9wcWPVYycPSR9Qf1BHYHQhI1exr8O3GfhzQoddnKtkRT/A7tJMpY6kVdY8RFwdFvsheHewhEXdS6
4C/QfFSafHq6jZRikLZ2XuUPAXDAM8uUIHdCw7qjZcYUs88f8fLSi6uapDh+BxCD6zrZTe+D0mCB
p7ESfDk+uRmWimnZHXQo/OO2RQjfo+yGbEpPxs3fKJwYyQvr/2EnDofAISAU8CduHWdGy39+lDEM
ZY8f9kOIfHBDoWQFwhX38s+8RLvpI8Sas2kMgPPmrYOFIU02YH7PNSTl9g5ns4bFJaxbmgX2uezh
jvxzeuCr6EsjgNOqLHStDfL1pvzIC+/SZp8S/QTE270n7cTSajpqes88csvAZKCp3ENUXEAp+1yK
FMgUEVzeHrjNMazTmftB5T7fMBoWWA9xJMKVxKzdRF2scifOt/L47FwPtnO2t3F1dG7H+mll4n3B
rdNN3efAIXbdLzau67iwAVi9jY6tEAHEc0aj7Jo/J3ojvMnUWZUvZDVgSUv3dt3Du+bRvcakfRIj
6UlO2OtiD5KrYJE2rYP7qPAgY5Z7NlcS9/NHDBAr6nNhFLuW9guI8VugvAp0ln7GvKpaN+xTpuSw
OTNb9NZi38KC5WrDciVrfIDttPsG2J3wbkM5xPZ9Ve3mk30fBJw69HwFSWUZnrbYh80/xITHqPPg
SvyWGSNikvvKBeRiUfs4ai5PaCLz5U/yEoca7yNktQcImvr5uhrHrPTCFM2LezTJCJarn1k+PGpi
CIg+zktIMcWfxWObERUtzRVjd9VQoftgN26wYwoEMC1tSBlEyDZPmxrzrFzwqgKE3fKfnNNDczru
AJ/y+iNk0eYPOx3CJ8xqW1ewa/xEr2BXmXwy4xmOW7Y4PziY9rZirrDATJEcMUEUzZHLg1A0mJco
K1pPbw0d82W23Y/IblIySkMuNMmPMB0zs3hNfV+CBjBUI17zhFhNOZsJHLuPIy7UQvz2rxxf0qdN
44jC1wPydEVge30vaeBDHawSrmO4uxfVnvviUuq2wVmVr1v4j8BHRtwa3eNawduV7WHBcg5UuYRH
8Fi4BBG8rzbW0kx4ejepFqfZM9H78l9btRU97vdXxltSmxf0WXBi+ey/771miU79f2aaK2VCQOwo
Ol3noiz2stZFIujpT7v3PhZ6N364/S3Ub6/Lq10YOsn5drg20ELHijpujun3rxm68HHByqVYQrBY
c+2YVYpbotHQtfKfXaloDahwh6Y0mpF/hUE6SO2NM1DCr7ae2/TkcL+pC2OZYw66SidPm4Et/4+I
xvA5e24WBXd7D5rhjhsRPNjXvIIKWB7Vh7cKz2uagUdJrNeZuflEQz6t76V6daUDbcW20ju54vob
l8afVUQ080gCpifn4AnfsVzzpO2WhhZt1Hd+wAcfXh+ymSLOfbmisLhJQlyN556FtJk4Owm7kHnC
T4IEQ6jRV8/c+55tduSuNMNzjGk8xPIlk170t4KwZBkMBtrsHSf4vpBwVfZJkcadT4eE/t3vgCP1
0qMefN7a702j2ANTujfkpmj3wK/tsT7SSIDmi7IYGbnUHfEcdXK0xCqsmMlwvYgN2jkF3cseKPXi
SnF0SeGqqwwEywASSQxpb4iA72xIXhQ8ywbeCA2Ufy3Dp4+BaHrvXf2k2cphRZAE5Av9Sz2tZM1u
a8240EwzZPYyPhjKwBez51/JblIf5gYAH1GOi/+Oay6e+vt2E/yn1z1yY9WV8Oc9ZXm48OWNCMD0
xfxWxlcUa0hUF26sVzVhdoclzqD0MFQtVOObmKu+cF3RlGyx5vwS2DLFNAkRzMg/4SS7IF04FV1k
zM1uqgr1HqXnuRHiEjFFrDOu54n1gg2huMAACanfh9yZFwsHl+JgeSCQxNdO6qu0O0iC7bQDRfCa
HWDDBB2sN78sjREmR9qnzJ1iFgRBo/keqQe619ujaS0kmOVTPuLoTBm3MDiNXXmOR3O3BKpxjUCP
0hNKBUxlN4w6G8l12noopu7u4Uj+w2zs2eJAmiC0rbR6WAaLTEPqQIFZTT5k1UgrD4vseJRpp75a
MpoD1u61N3VM/6Ew3V+rDAyjltHUzaG/7PWuxhJLLhTPLcu/4lmKXcchdZubfo4jABatr4ZVec3k
KHLS5zm51y6kHQC/bGCI4as6j/wf55d0C4cdRZBYzSe5Q8W5M7Qcat9ep7ht+8SkgO/brD34haBC
mCzuEFQ7hKB4JY0jgFMObRZoXjGd1fOfEUgjiKazTSGcIJIE9hYOmzNkjD0zE/FU5EjAw2qoGIww
i57H5hYYTPkDTaYBtMg0Ra7N6T8GCsfh88zpwGYUx6of5+bcRaqo1ZNfSIk4KMyiSToGuZREXvZq
UJFYR1YqTAvcrANX9FO0R6NHo8yqJ4dxL9zVrFx4yf4FVw4BZM1hHQ01XhiMluRyD7peDyRqlrXr
adStO4xQcqz9iz3g2IqbBCzM1OohyOD/lUrieht7RCETPxCRn1oaA9nEKVvEKcTSYjAklAGMVkaw
NgFNJzSy+KxlEVzSS/5XNsxGZCpjICO+I8uWGy88Noc3BaRwn3SCj/+AeO4mQgIjpyFc/azJeKU2
8KW/EH2B2CgwbEOa7grxlUCtNpU0BkX+EId/2Jnd9bhOPYCqGdJqfbtZg6rwqvswXD+F1aBum/mV
t+m/AzWZ86wNc94dXKAYrygQCeWNpf7qnjH1Kh600KpfsuQE9vEpk1jXCqNp2ZXrApkv7JTAIE1X
+C0xgYdIF6J4FlzWBZxqWiS6znEMo7NcMzp3WeX8DUJRAQ/2WghKlNIuC0/fklNUiS+Bc50PQfzO
DeAUCqF8s7m0FMIxJagPAGJmftmc06GhUW88qswVyaa/6DG24O+8QM5sY+KBrLDT1MWuVVJOb4uK
S7juPdrQDjT+1gvxyo5okbYjnM/wp6N2BiaABmXDFmm/V8GPuav054inArhz7GlYrNOLWnZ5s8A2
KO5PEoh6yd50Y/lrSEHLn02lph9Rtq/vdJd1R37IJo9pWyclfHw3yGBFawn5QVHLDy1gkMPm7njI
TMejVQoJUiZNLsezm+jsSxefDMbMxJLPmnfqj9nWtbRJ6ExbpF4wYsaQzfNMDA4k6zsEN+gmNtWE
UYT8aBtZxza6sFgfwsdSlQSKBQ18yJ4eWh3U6SAyUzLSrLUARWNuQs4LIxWZNYtanjMkimAF8GnA
qL4sdEsRYeyRnsdmgpkqLg7ZpgEaqt5jxcxSWZo1fiLf3jZUoDPGaqJD0GD3K15ZsMn6VGYUtGJb
4DCLwFJLfqa1PyLAwpVon9Ki1pBjjY7NpZptOGlkzI9HslcSSIjKpUz4RdTTGXnW6jk9cqDAuDmE
NsDO2yeuaiplz/tFn84wFO+cMrlZJAQ/9AeLHyTOKT9s5N9UfekGYRu56/xTk2uguenkY8EYFmq0
skPHd9GMpRUoTSN7H4jKV3T3fto3AntpRIx9e/htd1AYor7wztbQvtD1JNbUGvEaSqczidHlyRa4
BKg9hXUHh7OvSUXcVGUglggWkO1UyRB0f4zrzYHnY0hmnpnRYQkl89Z7p1i+ydsWxFWR+BHECt+m
Ao0O5KfMIYDgyH1uH8kwVrVt9nk5wTxZzZe82QuuwBP2OppkuXmB5zc4ZbAmdAAmAswnI+ZpIR4+
Reuw1wMDWZmqeg4FdoMBxj5nRMFJ8Bvpb1pYIWm+kKI6VboiFc+qETy5EjgfX0l6EnOu1noztiLB
jlIorNX8ZP16+RF2JmZ79LqKfI6+QKLVDGbtYrenCaFU8w+LPOsbr9W/0K1cHAJJuKAh9HjIs0AW
Nq9Uv1VOedmfEwX62cX+b6nkpdauqHT8LBmw4Mpx+0mu3Wc1/A61xtvGTARyw+YVuQ4Q6YbrnqAT
rWWC4CzE3FURYIAedYZcZbaYirHNle4+5MhUmsjnHP4fItsQ1C1TXCByhdCyKAD6Slz0P2EuOWga
Fr8shXgzD7gCZtF54NF26hx2RpNvCsHB0MouG8pOCV4Jyqzxg9Kc1woGuNTfHPS91H0cyE9Od7ua
0pf3qiAm3dpnt5RCwtPlKWxdJi3QnaoxN0HKvfx9mBBOwYPUQ03GM/gjD3SChSadXkoUsV5YOh9O
kOx1ozpkZWks+Dpzt40XjgR3MLAJDr56jqWP+omVSyF8CNLQkQ9QQWxU4lbHU/KlyqAAftcSXfxu
K37lX2nlLfPRRsq+Pu3fJZycpoB/zkfKmg3JGCD3qzdLOdfFlP4Ci9oDj4I2OkQxb8pLwRqCoS+J
sGUJpdE43nnyafXJF2MITlI5IQSxPgFHbjHILeX0Df6jGAuawhrlAdmx2yKW79HcqZdZ/W9EWxjq
vMriAKLOjjWzWJUXTF5E5QBq02l1Qy+UreoAmQd3Rw7aXRYCbrAqwd0KOcspAdXcvKWIrd7BzFGf
X2hBUp+sPmO+jtJcpWwTd3uFo8MU84Wnlsy/i45qxXheMiOAyMQHdqAPlKhWJi12NyogdjkBoivr
/8r4Jvmh9rfyUZKMRdP7tc84RraOrkkLe7gJkvkXp+GG4WDV8XVaCV+imxHmc8H49Mj1YdVoflUs
b8CBdO3vkzR99kVC/XhkbyvjcqD0r3RmidZ0HTz+6chx/XOFwoYXouK+TRxn+1k+cCUDd4ZHhojL
Ef8W9GmJl408aW13GaFdzkgA4f43jKH+BbFqqqa2PprvOkGFi0wLL5gHaWiFTHmUYXeRhscCcj6v
1tY1mjLtmVPv6NtjrYSr5Mre4BbP8tAnJgZNT38gOwDTkYjpUA32EwkX0ZOTs+/u3H9QKs6ht4Lf
/cAGT8mv4Y/WtIwpJ4MbvRmUYvcxvfc5/U/INLEPmm72gO7Jg7KvZ7y4VtLkf66fv5+941N00J+q
hME9vzHdo3RT80aFszGkpVruEiCzYrTFKdYSXNF/OkGCQpdL7Ft00ImWwCCgHsVYa/wvroIfYC+U
14G3iNSKCK0IndabVm3ATVEPDGZ4udDE8dRii34K1EtD9t8AgQuFfGfgrvqsCL8HfUblYCOBnQbq
We5+IBRWfNTTv7aTnYG+nG05KAbocO/WTjkKoOXH4yIuSg6FyoqBO0KuWvXZ0YBQEiiwpV08F+jZ
McjJoecw5GgaN35knKWihYysEt+athP4kapWSzc0d/ZxYZlPYAs/Ut2ohQAaYulnJvvplqRjNGW2
gBPucipHAv/TCf57yrY2JrrahoKOC5i5x9JIb+vOfzrSCJngQd8R5QvoOUcwwN1Rt8r+DdaCngyU
QFj50L9TQTKBEgqDFmhxtwFKUPWYgnMZx1BRou6rX4WILopivZxvp+As4GWuUWznRsobjY3FQhj1
kUSgXlH6bKspZmmuJXxHcN40Gk1Zjo9Ou4YXcOh3dy/o1UY9yFMbFnSBeCXYj7JgF4tOjzo+6AZI
cce1XDe2tWAtTwkYaU1YmW1jsQa8mOeT11hgLi0VU13aYManwssXrGfCRuAsjHwnzvsB3BCTEBAm
pqUPMgvVm29YE29UOW8zL6n92XpH2qzfggCPVwhty5Ue8+znn4hWF8RRgNA3+wfMYP6s2TDQDd8x
a/VHajhnT7x4qh/5nOxGCDWancgZOnalCBM6h/uykMSinaPa4d1CHhs5O6f0YvpVgqIUg9J5Z7qq
ZcRzWUiJ1oq07yFAE7uDWiqwfMpSuGgN9raJEZ+FyaZejB3DQSvvUQdzV6h0MteHLx2r9R2HlNhK
Jb7g1ortLMX88Vd3lpe7h5HFsI6bwu6lJFmcS6m7seV/TMystIVux7vMAD64c9mEzdPzPgKtq2WX
lsS387xOl2+RbbrZuTew4T4dsnvDN5LsKsCZ0fHtfrWk9FJApgAdtgN4wZuBy88fuPTaZ7o/BCeV
h7ssdW7d2dtqVJam0ih5qsF8n6j+ySv18ewyPjFwe+Ht+LpeOl+o6ZA/1SPU/3ZDIa8UL77Xno/2
x2O+cJ7IAhCMWrP1bliPpoZH2qTo6j7sINhu/2jGeQd9pARu7jXowqQJq66sN7PBdOTWlEwt14Ur
Y4fZlSr/Z+ICDPuPu865ODz748PI/uoRkh0tVuApLQ3r/FUte/J31nDrvWvsB7in0KE6sc8TotQo
WBdnhyOOgvZHkRWV6Fy0FZR0Zvfaru4jf7/zZ0CJzcUcChvRXTyzOwMz24UCLV5/NeomSUJuEAjy
MGUPcxuVrKNfGVRfNetm+pstDj+lVJDoB3RGY9UsC71RN5KdcHrqofPVuFzJgUa7Gl+X6f8CaGbM
aCLA3wT3E+tLPUkOt4znnhUFZKOCXQJFmBISq2JaC+dmgOBBJEU72lFHv7YA4Fikt2JxLIsr+DST
Ph27Ek1rtla4q2jq/SFXAiD8WsCF2yum9l3M7TvKVaNeud/fGhAhByb+iYAEMtLgETbvw7NHyvuR
DCVWkumkWpljPuR51CUkChFSWPI0CKel8iGCAwo71aOS3Fw0e/0LjDTY5TX91gaGIW39DKI0aKTX
RrHWjptF0CvJpCg+YecEZri8WQybQp/04F4bZoQWozQ9E0ZZURyOO1L8QiMV8fGOMk4VimIJsNcm
Kd9n5eQ6NdMQ0a6qucT7tMiDl8MGpzCb8rZEmX6TuD3S5dDVDLmSSq+RM/E0oaz2jILhErFoWjWG
ojqOmLktGiXHrX/125hdNdlPF6mRF1BSIH+snCkj3J0V1uCFfxjte2So6tJ4o5AlN7bTmPkSeMh3
lkf2HVkBHgKnVu8VPx67NzO+mYiVZG0UZyrJNeuCeJ1+2f16WhM3Ss5vf0jV1w+mXsOwcXc1z6Ha
MVHpmkxVYMuflJFBuZ8UDB1iFxeVqA24I7qR7YNw1NXySAAr+QL+TaLJHCKVsjDumVA4dKmuS1xx
TX1yknWe12xaYsjqzRi2cpg1gmDzLrzdq9YlWgtxpktuLnBsc3gRnxOVT25p8tnP9tfq/tdWfaPA
Y+ZKihc/C7bmFhs9c7J16FTi+xWF2mFTMUUxi+5V8xv4I6Gi5k0xE6PSyxvLfLcav2JRf2mLK2KT
px4Pf6BOyXE0wuCb1zgOFLVnNi6PnJk+Wqp4os25nYRj3cOBpXp92xHUenRKb1cNznTWVk/Wl+K/
j+SQGPvgay1K2v3epK4Zr+OoOV8fttIGxKmT3P6Tu2KeznbhGPgxC2/zlteHspYsR90utlSHDIH3
XOf4MC0LKKs/138qhYFsfY7ZDbHOVjYiqCjbOJE2JI3HwIfdwGSdeQNFcg7bWl2syGumMZfQw8Kt
DNE5NgjhmnOOxH47NCFAfYYJr2h2rG9oc0o0zPK0yMoW7iXARvSFCPvqciqF4OMVsH3oybbD8LwT
CxolgZkPH8nuMDDEZHBRX9qV4TmmjwscFn3Ywvq0mpBPu5FRhkzoheTmsLrl+sTQH2Ja/GhZwE9T
wuzQX5uj82dKIXwhZD9zZqtNXJeUGpRvn/NGgoGZWWn+sooOYt7b/ysFZwX4O4u+NSqWDQaLwUWb
gVr39+HgY2RvnCvpgLvszEmXA3ecLK0v9s9JE279b9ND6coGB643cccxOsx7ADL1IkM7Q3KsOsgY
3oUzNtjgU+z38uTqyzXrOllaQbGJF1yCq9ueCNvcl9NyO7lXzuZ4qwIcAOzbRXi6RFjHVxniIS+W
TMtNv9iW2G+npLKBltBhKoLd6D7R6xZXJpRF3t6uNmst6ScJijuZ9sNsuWbMxZSj4CuZ9EM7H3LM
64k5HAMyN1Chp6SwxfHoWNDMS0w08QOPOeCTXueHYja0iEO7PkipZTWB+hGF+wgwEx+Xj//m5sEI
UZB+QjmDJUNuEEGrYzh1HveLemmZ0QDlNR961rdX/xc5g8ugaenl5sO8DGF8tAtMCHw0WYVfzQjR
+aJrwiskqg7AhmrTtRgunm5jSWzz1elkIXpkq8h8bXfxXP+AnlVn0LlAUWbSvdO8njp4b1CnAmkH
3yeJfIvUzzazvY9yVUMoOlyk/dFJcN0pAfT+hJ67EvLL/nokyRU5hJiZMr7WuWBbm/xXWFV0Oz1n
yS17YLnq5UCe2xX5QT9WL9at0jB/7knXTfoBTII7v6qJCZ51TTlr5Gam+hhtI3oxJJn7XSqPBc+D
K7pzWvg68gIsmZSrchjs5XqfLlPHyAmjR1NBOj1f2gfPvzNMCmDxSSZtw1n+FDHoUWCDk9NvbMhv
q0cm4V4Ko4U28U2B8Wt6Q3zoSVTdXWm6ZSkHJ1/0ci1BeNf/Fq7ekIlSNnrMW/9h4GSXb9H+aPIR
60EWjAjNrfX7UcOfmLuCzmxP/dW64FpUsshKuJEB0+oOroScki7aL/6tCVrhQ3MWnFb1xZp7P4rP
LhrY1wVo7v6TaRYL19CwbTAwCnHQaddUlaAPg5ueg4oyHXSG0SdPTLB33riRS4Y4SIV61OsTUKsu
pnQhxzvtr7adSnfBGXfNftx/WgS+zNMIkE+s/fvJt9lRZqnDGJsYrb4cRO7K5bpMyoHYIrW0J4Zh
w5CTBfNyAhG1fgi9bEcgOTFb9oM7R4KnWwTMx4/Yzd/wQbqa0RXOoPRf+LCZHgiCiL7Ix39tbiXC
U73kcYMiibNHVqiRfwxn23nwmuBYW4RUIMUnbWGlMmGxWm74d7tFkajCh04lkn1FzIJLfco0bpuy
Yv3+vmLEoI1l/Dtnv+Cywttue0bTUYYuaotGKBwVA8lKkpgR4sd3c7yTVp/VxeYmMib6Md+BTNJI
ysnQgHIDqz5f8ghoJS2RgR3v9VSKkzoV0IM4noNXBgeB9b3G0kE/OzTHvnUQYSpIvn44s6pvQM1j
r3EgQNPyIV9TD2MenH1+XAjfRcvh3ZV3J9ofvZxNf4byWhgmiLusz5NkOXMKGbz4uMNuzwqy8clj
uVUtGdrpHCae7lz0lyK18IzUwiaEnv1mDr7q27+174gxUUE39WUrRdi3aLiFfomc8DWF24XUaVtk
CYddgt1kCY3aFKnXFMGtI7weoQ/JcQ5Fns24+XYccgQaHyVZcndNcIm/lZPqpaQXqQ04Q4d3GCKw
Fx2aZrZZfXX3hxufrIWmtJ8L4BBri3adw5JexkjNw7dOkoptUdd/333+8xrBYw4ktYzeZqh07hHR
xVBQvvZ/nQK4O4pf41gDWioWKVxSfibDq6r1VYGhJLBhGtn00SukgFhhi9GH5K7z9JSfJwgoJ+52
Q4/9bPI29q5kDf+xmGcY9/roob43yPQmsNHVqehGcdIy02t+F+iMAob/hMFSF0cR87RFswl8dbsl
OrbbG2gGQY+2Ckc97z811Nb+ViUk2AEkpZHAz5NjlxK4S+mUhxiby3RuYCoB1kNk4LBgGe4Gp4kE
DV4zqGLgMgB3tUeLKC4hIbavljsalqHXue6Ai47o9Vn26aGqN+nTSr5YFe2cpe2Vc+B+qDkb01Km
iqfMGW3VueqkQKgIhwKGinaZa0t0fuozitNAN/US8SILAH1/Ogt+FjxR+GSdgNupt0oCPmNDW5DJ
51k0RlId3R7bYGZJqRgCLP4UKjVNeO+yzEq0FXp/bT/OzZxsZBMWYxboKRoZuJ+MVDFwmbegpB/i
5lDGglzhRJY/3eFG9YaU5q6f4ONvLg6h0UBNgYgQSCXp4dx/gqUkBSPFH/EkMu7woOeZMBC5usF7
AUGpUpoRL0Tr2Xsv4Saoldxvw+FBWCULzSWstqW/MMYN2NiMZnafF6X5uKAEgo4i8u22CiHIIVxU
pHQQPI/Q7n5A+qYq2+SZECr1frki6POMdk6FEY35o7r5NUYvfP2hwzeYgC54pQqoDaENkVN94uSi
6AeFkYv83pZVRUrr7AoFi0VXfIBRo0YSc58qZqBfjQItHeYywYpU4uG6XrTUTyVEQlq4VzWOto3/
pVPuqPWs8uf4iethv2X9Ji/VPga4sigpoMcyEhlfAsemTHosgOC2bWxTef60dtBZfGcO2jsxyAUP
r6XBFeRv+E+ycw+OFHOluBvkAPuH4f+MbgMyruXWoSg4yQxTd9VbE5AAGu+OllSMeWD0Dt1EFshS
B/MveHQ6cB+ziw1TGkcrkfAQ2l5PFR4LUsHpBiKN8AvWd4gMj1/i/QUoGE889fcHcnnGCUE1rDtT
BbK+oaQzGGljFKMfgMtavx81Er2MccJvxaAU8Nwxo7hMgC84RVWfRuG6XWlSMSD6MpfTKHRnhdLE
RBgfrlp41SYa1Ia5bRAKyKxI9ftqUSokt2ywnd0AMQwS7XjZXRxJ/RmQPawmj1knV21Wy9XSuV3Y
cD81mbmLj2vkBROghst61xF21WUTIoYP4+t2hXv4A40HE68jagKsRQ/2GKEsRkEH0f9mQ2dm/RlV
24oXnIpfZOQVlstyAo+wiftRqsqpiD3dr1a6sVm36C0rHeWzCwQBVQBG3p7gc7kgk//6s6/3k1ua
4z/M8uu7TxNkEu5efYxrRUHBLNjuD7ENXeyrUWuaVD5DSWMXlLh7MiaPO8ke3m6uP6kaJZ0hJ0zz
XTNzt5aNFsCxUXnAWW5pLoira8ygVnVcIQcunO3XsItnUuHbCTlPWOJafO6fw8kAGPn3svMAdA2q
izhDJWl+NTzXWKW9iH6oe3ArWnBpPTcJLbr+VPyzNodPHZOz7wG1SR2O+XJpDqmDm7tPA4RIgI30
QaNECvYmQy6zIEcSOYDFxBOmDRKuC81ObgqrNe9Ai/WpgzmgJYlsR0GneUfd5hytLTlwAxyDFgwe
D+h8iJcbyZvWhQlFvT72EEIhFu/qlPatmB4jGC3knLfMd8lHQ6o+YeRCeN0wxAeETD0iO6A8f9eK
2AtchioPVg0IwmPeAScm5Ogsoz5o6HDC2xQ/F8qcDgigJj3pi37stboeC2kJx61fB+7/yLJdCu4u
FLCVVkf9W3xkbNv0D0Jv7/lDBM7RV7MuOiDKhrHBlqRX/hX8fiDrlCSSG3ceuNLUPe4kpfpD/z+b
rRgcbzT+JZQyy4GsvL6z1BoEx1t6a30FpbmRUPzVW+60+rvmrPUGJnsphNefpuw0nc4rQrxrxSSi
XxQ72xh+FX3zWjnxNuLdNK5e7EyEaFkkpOpULMvBW8LmJmWetk1HIWSMEmetbhyWFXqD5xeuT6Hy
bQeeruvVny/djQK58OUIrHzE0rcI9fMSAOgswUcQZ7Df/0YNMeEowbAaCCA/h8aBJOQxthcGO4U8
L5c9hTmbhxCSZYsY1NCelZ/PnR3ScQluRI+SnNZk1c9kx/PX03rtylu4PlqwxaDSW8QiHAAuRLRp
Eo6NgLoDkXL63zrN8Vf8Tq+ybVT1Yo/i1NReSYgExIkHUn3N2iZZvuPA6MQ+hsEu91muke53vGJp
G3MNcisXLYOoHZIL1u1AsNLZy5TyBdpy778V0z1pRA1JelfkmQHpjkS8qgyFhEAZ8m1qN20QGtKy
FMmNwzxHbuzezRu5nHNASpUtjUSxGIaIObD94jhf5xEmgkoZQ4JDbGj6Uphw1T469vbLjn2nOl2v
Db7ZCTc2WxWXvh98ZvhiG4SHmuwbkireyTzobYh0sHbjLvTlOgN89gvznSybeKFJRDK68vAXL2Nb
msITteB44+b/fCfJZil08ndkescAYUkmg1U6OZ412vamNFXQUVXA6t3daGovSzBk6YWggWq7bMdj
HspyEpr7Ox/jdN6Jl2tyG2tR2PiFLo/NIq/sCLP4Nb4MM7lknOU7d/Z775GShOqEJDwMWZJg4UOK
MzTTqEx3eKK4ZWPpdUvMlEO5mS/f+JCb0ErVeeHvUyNMU9DsU6jvGmKl6F9ae9gnvZG6ylCuVJ/G
CO9b+msSP0oPRLrfFO7sUQ75GeIXWJJf20VqCi10ZmiZWGXmYBMHrK1RYp12/AsU3GESn9Ohotn8
MSRvfPRE1B3/pKrTxZ5OqxsVKEbXXHZ1+IiohiX+W4AA5KuLB9b3DwLW5p/LMUeZT2k236kPMKzM
DMwZbh65CdoRH1B+FQflmLbnshTLLrs5Jp8RQejruzmqTbR6EbyteoLBRQR8wqRPJmXMkmRnR+Ah
GXTVmgrgPUqOV1LNe8XnEG6sl+UovALW+mbvl9X6ZLE6GcByCyJcdif2n74RHHwEbT3jvjfmwcUl
nmIAV2lknjCpJQN05MUHhnemHk/plAEHxHqLC0/QhRlQx2uoBRyd3G22A2OQJ8ebDYYwxKjofPTO
aVCKvC2IZqF1yYvnTCBPhKrTeCxnlwPYaHc+n28UUFcRveqnoHDamyvcB171UhjFLJTaC/C9AtTv
JSIanmMHPYzF8VkXa6YHkkBLNv5T//4SFBrn7cDDFgijzfZki/ZfFzvdMFR8PhychQTUpYiE2+3r
ISC0pUiGzd+nT+xwakGOYcLYn45dmMTK7Nd02AfBCda5x0Tv2n/3lUjvyQ10z2yPCR7KDQWDk3b/
gNJ9FrcwwhExiex3janLFKti2Nq8eEjsGXAyqIcRqIzNqei0hfYoUJDV08t7MRWwrTh1z4alWpP6
Odpy+SpjkV0QZN2MoRpyksDPCWQkfFWgkBDCOcEHondGAo/AG32qJ7EhodLeSFebAy+YAUESzqIR
Lfl1NkR0a/6OHG1XmhT7ttRasj+XVuCECaHP/gTbxnbLPxRdR2uk3XdyILBY+0BEgZDnjX37C4B5
vN+18j54rXN8hjmnfxKSni26o1Dx6cLEWwjVLuNs1VyDIo48NwVAy8Y3SWNusffszwOcW92kAWA/
f9tpsSNRuBVY572dGHrvbE5pE4STn6Ft7SbBsKFpL2b2CUOLauiVaKFf+1aS1N8q5oWrgj1RPIo3
Y5F0666e6Xo/QpcYD8HSLsRs80rShvvCg42+0Lob1AJaxS0B4e2JIpwiSDe4rWBlpbHMeTOF0qXe
hy4ePn4vnGdRYdAvwpq5D+wHKEcNJE5igUMcIqDxiKJxpUu1cxTyIANNCgISaqgxu8mTwWKzITW3
zh9qaornyKJlKTS89XiVgssx3rFE0tn+vWpy34F4hYKTsEUdg3D4IbXu5RmgPGHFI2e1PGbUddG9
AoxczrR3ylimNI7RAlmMEgpFKC2Z/fY219Fm5juYQasXako6pWOQteCF++H5wnJ4+LIl1ALLGrRt
EaW0TrbRJc1lprZQvOBP70qDZ2k4DEIQ9xIbentAmdB6grMY/mWkrOzF/JJvrcfiRgjQGm7738Sq
IVBjPq9H1W1CC8fkOPwRcZya4qKMLR6eaaqserRsTV/nPTM+XeTP6DcDbhxiddmVWktOdb24XpZ2
xh1RmElTJH7t+TwjWKu3SaiQ0kqw+aCrUmbRr9KmMLpX/zp+VxH6/pS1QLJLGL3GHRvNzeJFn02N
0+JQ4nbo9pu3fRX3NF5UyB+DM/CIMXdohce2TrDtEts25ZHcYgZe4cCj/F/RcjPJ+gXbHv/zTYlh
PdBzxNZebNJ5BYmFw9Oy0juwlx1RvZr78iFRVl0CCQikHHhicT+f8+OgYrTSPaoPsDskXDW0V7gn
qL2gbGctLdwuC/It7/mSlcx/X8mScOBcP/PgBQChTvsH5/8oeJMF8h9ukCLbNeJ84JXe/IYPDmyK
ZVwbPwRKqYido7oygo3iou8OGiYp/8N1X6Ir+2GZGPhpWQBqLZ3EaX2YimAvrx9T8w6FuOLDQHPV
p7c8ijargmrt/1whvWAvE1mYSsPCs/ZVuaRZDzE+E0ETaSefVWaCuVyDnttdTVdT6ST+SyZT6/xe
Qx+GcQW95VF8WoqNx7qshDJqm/8qFNbwh+RCkcgHlB0imvy/a+mb0cBGx+D6UTAI7eWd23ts8dGS
YIQCL6O1hSsk83DluF9H5D8L7AB5cSNXd2T4ruwyDLqiGDmCiZ+tbuhn1O7apN9tqP9MFnvjYFhD
/kyfFF84gs/KvDsXHASzzP9HuZZTfoLiFlU6eH2by03X/bosUscI3Bq/Q0QQLJ/oQ3+s9iiH+18F
zz1XYCUEfEAfxv2iGYwBZDXgwmojObCFE83iCINrL9Y1DPNfquHqYf0564Kaz9b0ld/5bMWUsDyT
OD2ky++72zHe1TiY0lA/HzpCtscUGVvrfCBDfI4xeYMK1li2XiI40eRpSHiyTVFgfD1WciII4O+5
SDSfPC0wd814hyp3zPrEKDRAXnMWAsCsTkWu4rCBeyHkrZS7kq8JuUZX9oHR3SKZHbcTRt7XTu/T
bNdInEePyO8M5AB5HUrSS3nOBbKEX7LzhdLfoNxnB7+m7R+h7oQAxyqrHePLWxb0f1t38n54Vr/o
gvFPl0cYMXO0DabCjJngcIlPt/cAQaQsQp4FQtU6Tj84rxF5DqtFHe/XaFFduchAHLzNtSmGYJ6u
yGyusd9ZvYnw2mxeN4Gxg3nlt8vywfbIOgxKh3qRgpZV4v7MxeISjDWaqnMVrtNvg7Kx57s1Bwl3
WgBQQzqsecLsxo20q0JRgrSZIQ8C59LbdxesjNXjsZjE4nrisiR1cboInRmHDAnAnAhlADj6P1pK
Ohvx9P0JIKcNDL+bN+/DiA6X8EB09mKbKkToaQufIBxTHPllVQqjRTdrYDrwMuGgcSecb1ROzK1Q
//9wZ2t+MiNUcYpag1qXzeaQMGWO9Y8z2QOH9+LQd8ZUIqmlhg4BRffDYn1M8Of5wniRdMm+GRWn
zHtIkDaV5tM3Hg3lOIvDrNC23Mao31P6aPMASRY7Gjkq1HyUehJEE+QUjszVEZ/8QnXl8UCyWoIa
BkVyj7/+Adt44RRxe/L2sxtZzlwmet4E4NS0RrObimDm+SaDYTsl6k2yM16zcDBaXWiQIDoxLE8F
EYz8r5Qr++eKBWSl/38A58hG1pc5IMVmth2g0NiQN+p1JvyDCzWGd7cO8TBFYmQyUI8TGZFlTukq
Wn6L62TpMNOMrlTcRIsfV8rfY155NsoKvYNJ2brKB24aW0lvXCDizp6R+s8bceJgZ3lxDMqiE4sF
uH7mBu1EwiHm9sB0HI6GVJF1MkPjoj7eMHSA0gfiW32qBy34NdLv35fFYkLOTtcKKP5/ILCyd2bV
hLZJBrPAsE0uqwYJbJXoXkI0tqzBlKq6MOmVxfOz4+Gs0rwKNfKRADc6TfmHVqZkhavxW/EGZXW5
rqNypj9+MnCvu2mpHwRpgO1+u4/diwLhkAU+uD+XQ2f2PO1MECdrJfKS4k9aqATSxPF2qYDP8Utl
BwWW8pLrRNTtvRsaZ0Cb/gL2QYl+OFVgkIZIAvnDUD984RD0jOKQFYYJdEzKaHAuVDTD8vUzgq44
bhfUavHbX/vii50rfjPdwG44kUwRBLRIApswcdURtsE1iZ1dUsRmVuZr7fSqF6eHOi1XvGGL1iwt
V/mUYxcPDrHcnucjJ1jdY49JNamSd8+xD/BC+9X+zRHU5zzR/HZIkcS8RWITjnyANZVCirfh26jR
yKwtJsWqt3Yw5WEoogOQAMEmlobcRXzy6luOdfcBI6s+rb/ctgn6quXf9YmyeBB616cBd2BJKafJ
HKUi1r8wTKf11Z4Plh9fzFSLWtvMoUy612n/f4zxcsJeFiIhvpSmWfFez00LMDRtJd4+IZA7F6KT
WYUCPO9eYFndLq/gTC8Go5wUZYuzS4G8sNMzPvlsWrfGc1jED+pzsJyJE5D6FJWG3oF+hLWOsxJY
ZZx6MaVYFkyvkB0AsJO4Zm8Z4ENt6ghp+yPGUR1ArI8rvtTh3KOJj+frclAgrK23NBQvmJPYwJYk
Lq7CVu++/bB/he/yoxoHrUdg2nHqeQ1r1pnV0XTVbGPPGoW1cc/JzZTMuXEnZOQQb0RlabXX4cZ8
QIaEk8UMAatXEOaPlRFN4lLB6vMvZGhoS1w26kw5CF6eEpSuimYppHPihJVYQ6wGsXYlV1Tsn3ue
NSDuvkDXs+9LYMrlAmiZYN8UulMsogtBIyApVqgYlMqH5d+wYtbyN6KhCzoUhLJyMoIhhwKG5XtP
u/DrEspwijWvTX/MniF7pTb+lvMs4ACmpyqaB2dfNB+3CuFejDlnn2tPFZigfslnW0gboMcuyNxW
FfFge8QFnawyDAl+YuLfiGajpwoK6dLpnYDqP9wbcY5YnGOqDi0kU9kmeb6GWWb82/Pi8dQr4zoB
kXlMVWVzQT9/p3dqdMqW1M0b1S8F2bxGVX3ID6y7H+psVFDw68AWihzorfgbj6KIp6UgNfRcUObg
ElXnvPpz80cYk8eq8LIibjKgMKI3ts8FBemr11N+gTnqLjRbB/T1okerwIjytPwSiWrPSQx+zzYh
Rp47EYuFLomhdW3IrBo7hBuslwRiPM5qhZapiAmXxnwyhdJkqPSUbRd75Kjdz4rsxOi1OUpTKuzQ
pTFk9p1iTLxrdUgVEJcfMegdIjCwS5wjB2+y3TK4PtZFo3SPFsHIk8mHOHiHkp7WXKBAagJ9Hhw3
RMLh4nkh2Q2EozNJl1JPaTVUt3xWmLfdDczCrmQ/xko28dK7zACqcUltL4APcFy8F10oxUSwyobk
sfC1AjuNpBE18wvJXgGqucGzcgEdQ3tCx0Sw5o1dysbDEmA6xxhIKlvcRfMbS4FgsmGaRtv9846T
DQDFAtd+SIYhto3g2MwV3LegTwYFT1LynoUXeWAh5P492myQdQZNS53wIEd3RzKCIRGMjVkbSf51
Qp8P5Hyo2ztC3Ix0NimkaBBP4p3eRNgoqGIdhwilTjPMQtGTBs63xGzlpYvf/RvVW17lG7xjozVE
Dk39OHYP0bp+H7NKfpxIfh7eRwpWV0DnCMm8soTIkwb39Km3hMe5WLlEsbH7eCjZUvRTx23MOo1Q
IkDZP6gGWLHcRZJwcmZ5AyZNLWx88EeXZrI/cSv7bdSGdgalGw5mNmBbLZNI0eNipuse+HgKj3Kb
JrjE/9DJcK4PVVc0IlziLn7fMu6khrbn1vSd8zoNBHRKffJz5lbEDtg1IKLxa8NOjoDqTkOWtFW/
eEDEsSUQ53D1XNwcum0Z0Xk1oPAbDLlT+kGxUy2KPgYxhbRN3At3KwYO0F9FQamf3Etu9cqFJM4y
io7eCfa7ebXNskcHc+N2a/nWwNiyTbjP2i86StaMu5LJNLnzr3twD+U1V4H9HlnqfJ/GKYnbQDpr
/eUyM2j5StDT6XymZau4GPNcjZaA+GbJUZ8VIYnpv7DqfWO0cE0mOoG5IoEYeqUdmiDyHPcDqqlD
3ewuLgW3tphe5L051KiN4yp3xiMmaArz2+MfUvrpAQqHCIa5/bbU0nqym/fxTg4WkxMkDRsDmjTM
9Sv9QXdsssmHw/CG7MQDq8hdZEXPOPD7V5GmGnOWSiZSBVUvxbMFnZ8hgySbaMk2682q3G/OKtZS
55mtmjf2D7+tt2axFK+kTG7g62Ngli0/wtgFfLpVmx+nGezYmMpBxVUW6fmS1sU0It+2icOZ5nF9
A3BnHlZhigHa0c3DhI0plmo8DE0iQlTNVKyp4AbnYBb+kq1aqyb35GNA0KTW1o7SxacD8NE+vzqC
kvW1TC0iwNkEJkF1NCGSYRaCgr2iyFoSQy3NR6H8GjaV/LgWxzCGWNym/wUOrpRfyNoXH3TjIcvr
bL4f8G+98aqkeidbyMi4QCD/R9bb+XdUGxpJJpfcmXWhev6ryJhDZCwwfNSiJ2m4+QdwX4EwUQUS
/spEhqNMCvE0RIca6Ai3UlfuJN3GZ4VcqXKpcwYc6VC7K8U5DiQSxnyndViD/thbq6PFFD3g3E8/
bE2fSMjhQ/ngZmJEgqRXUq/RxaX1ynKNsxwSpK5RcrUczl1BpS+4h64h0rct21E83U2PXuRUImUF
qMyVXkiARC6MWe6Aa+tshusTORvZhToeQb0GiR8HCf0u/fixT18IqPIcwwWltnz8A4qu9QKFEHaC
rGWHlUvQ0/jPDM+1p02OpogjqPAODeOYboqJUYSXVT/xTqV+b7erIkVr8rPyK5EZfejZ6h00p0qr
iPBnaeb6n7YXQ8RX6HUXQr7Xy1M2TZrEdc9lFLlCqc05rEpTN5g9I3TVENNQ89H2bG7U9EC4WBGg
tmHNVGgZi69tLyntxMwOb178F2grMegBkOY0+nmKaAoRuTa/J80oQoaEmqYkbnIjZAC4cT2+auOm
6valvXkAWOMhpCQd7Kq7VUPBYmPWUaihDy2Gjj1cqZQaI8FKhsuUQ2OMwJNoHvCZnpOPHffsZ7gM
o7HnDMT996QCJN3XyA+fitOHgOp7FS+HhIo3o01kYGRyRAIvu6xlo7KbR5Goltn27DHr5FbwZyKf
bms9M+xoAl159zIlIL6dAEbsPxiuNzfSKFS7F5jiFnxjxRHu+7zdFHBihFyKYq4r6LfyTGC9mwxp
0W475u8DOcs1fEj7SDogOM0L7pnTioEo0pZoXRWm82ESdDs47zXZu1btZGYJ1uprJ1+RGExPGrB8
G+VSnukL5MheA6uUh9EFCnjNFJuhorvqlkLKjxmv0C7QZabY0/MXsOk6JVOYOiwdPu+7LnM1/8vb
Ac2hWvIWFv5854W8Ju3TfKqjZCLEMJ6jryYeLlUh6F3utMeLTCX3NPrvYJ6PxlXqmbxRZZmu++CT
b1Sg7lVYteEXrxHCRzPUzRRhFCi3Xi2Y4c110NWP6Fq5prglXvlh6LpR7VbjMlPr5j5jS/x/RqFN
PHkT/jbKd94a8NAkIc224hJjYuHFmxMtnLFzJtxeKCTvRrMR8GUGg+liWmJ6ZooBL8QDHLg/nfmI
13UFT6agOhXKvRU9t+hV4GbDkC2Kn9JX9jkBHYJ/kZBQc/ZGUOMpxdv/aQiDK32IWKnd1vNkLm/P
6DZ/q2GrV/KcOiHyw3lBQLtvcbQwRjfACjMe7Tm21yflK9/0iz/2A4oxG9LcadP0PAxMOw7+Rigx
LDZlF9qlZWeuqyPpOVYzOWtRpRF58rAIH/YW55dCQkThjyehygQ/ZBhUQXhQDJx0n46elk4htOkL
P5GVKfwG59phNS3rvgZ4psTvpbIlL0ZUVJcTzF7ygL9FHAFskAJM1gg5liNagtXn/c0ajs7rmmVt
sAUTOKMb8UeE1K0WfrJ0ePSfzrHQX+GU2mBCSfKwk2Eft1bo+9y2l9PEqxsG+jJgIilqDLTyr9jE
KuzRViWsD5tg6+3rHZtxsnp6kUM0KWRmWFbuQtRl4JT550v9+wbkrWoQGq66VMzqEj7Vt/7+y0+r
6Y5EMyYtSZ04Vf3VFCICbmFQEP0797bKweVVpLkStAHfyLVSTcMCLGY0U8y1N9y/lR4vd9kX9OWO
frvr8FwbFHe2JknQsuqM/TB1BC7phfPy1WRVVUf1ZkumxgS976xOb1AEbb5pWPOXH8ELC/vAEPHk
5r0BiBPM3cS9RHhSBksMARZExMvSdGoaTVFxDpydXySUeKz4uMFXHQQyFFI38Rm/V4525hDsvocE
JJM6PcL2MhHiPJt9Van6EUqzqh0YcUE80rvTPvQGjEohaKYVrN8dB7pZRb/V5WcE1K+M9uVyFOQ1
5NoD8GhfdeiARY9Cts89pCQMjOumf5lb+aDtjiMRBvyjqnpdc/WGSmhpFSr4emPoog4qlk3Aj3NS
xfiszvI20qIpDlrtAt9nAfkxfl6eC7KLhl3yEJ5CzXjlmHurMbUNber7O2ddRI95EKPCMnwldvfm
vjkmu+po8FGtkN7pbf6lqRg33bACAVaBd+LGiy16L504lHFSyXWK0ttL/Z/GRXCqgBbdiAuv9P1Y
a0boTcgIY2b3i3dFW1B4Sy5Wc7uk/nt/WmdMwynNbSn7eNOHXaGyIi1imVRGI9qkCv4EBLXEEWdt
q0Oni+1P+VBkAJ4CT1IG9pbJHhuzTSH8I1kPScjkE+zcHnM3xDhqVst07lg0KaTU6jzo2Hm2qsB0
4UHl2QEbBVuOpFyPAwwkxvUs+2M7y1CM+xJO5BKiFjkwOfA/baDfWn5dS1gIlFU19+SFEAzi4h6u
0N1HbUaffNKiTMVggEnSMSppqJ2HrXxgSHMFUtVN0WLv+O7GQYzWxDD9TJn0Lod6HUjW0dHu5VJY
A0ltie0Wew0n+NY0GkEUntHENm/5da61j/aAmfU8izEWMDNxW1tIY8KeCbpw5weUGXeVVxuwDNvg
8HImBqOIONWzMWl54+3Pn0Vbu9afovXzg/QYDI9TgjGwkWei9LD53ZElvjoJJY4hxDTiK+3qfXFt
QqyE6/+hPKrP3X4ZJ4bH5tjkUnksVMCb581tj4KhLO+8DiuYLGGVvo2ha4P+ApmY1428QoMd6cWo
Zm4eo2Ea/nmbUnxPXmmyDj7HXqBZFvssEBahX3xx6MDq0m4Y99ajNfXax89v90D4zJGtGLORDt0Q
1YqkJr5nmZScQXyPvWKiZDH1VqLlZEZjrYuHYsKI1G0GI3elJPqBdmMGV6sOnTz8roLR42a61U8y
CSXUESNZeo1JR8sFsrBArzEEwX/nSgiaZpTtBckNti2VveZy/Gd4fYrlSBCmxEzlKZQ2SON32GJv
RI5ZLoBGChg7H8ao245bsl9lw8PerhDCc1IvQzkG3uCFlE6om4yuQGXI4jOuESBZ4WtxClfr2BVm
HZZiFgeoF9Wo/Cn5mTClisG0BdsdnaAu2tSNeKnUlVBLDkS3CltKqHPUD1W1plMrtZLAYVUFrwn1
2G42rKBjrlwetcAdUXkrAZq1d8iO9d177byoLyuTP8sgHhukNMtXYyPTd8KmM48fwG+GoCYe69/a
KdyB5ksd6ET1t3g05HGYBKyEJYUEL3SwNOdF/yAPgB7YvAIf+AybCXW9DmM/3An1w3lc9sCjulx3
JKntF1A1/UDW2otz7RQ2xX+D8m73Cjik9IacqxI+6nw//XdDO6nCgS6laVBnNY21fp9+7ocCcltl
CW7yuZNYBoj29T0ZnIsFS9V3+SmKvUFxDG5l/BUZPzo5vKidD7viNMxaEyQVwsx1iIWw65iFhuoD
0l2UojpQZEs+hMNO8a58dF7gHS3Zf9qjUHMS97YDVCEg4KJ4lPHLCiVIoJZ2p753CUs1K7dLzIVz
cHkD90InH5PNmoOfETbd3DlwpmwPxT/cm4if+g+uLybFj967fFpRm4HIAKymiVPFlsrDsBrY3RwG
4IVS2XnHAeUYU9CRnSZBueZn91StOJKc3otlihFxxznQs3d1FZLkvLSG1f5V9eTsv2scSQZ3mR/C
F5TdqFdPKtUcuBBVOPyk716s7YzZxjhxWdEjMncV+fT3wnD40ZQHHR1xX9Vi9cWPYwYw/WYY4Jh+
c0rWH+kyxbw3PLgWeNxwySgTA7tCONNOy7QF6DcHWVtFPUZtK3HTChg3RmClkYzOMfoly9JQgDR1
ot3XcduJhTUWOhw1uf1QtyjK9vt9x76YncQfwAMTag1gRS6qzmHKd6EzbmxmcIArZ/XJq+rp8BiY
KRRlZZBtjqyoyi//2bWY6jWTlCQ3VfI5bH2p8bPqJVTUS+8KVnJfnQaxuh9Tvo02goHmDXqMDeP5
1pKUldWbQITnZnxsUe0W1/g23vmIy9KATDBR85mVQ5QZWpIQKWwElETV4HBeQBcbkTxM/dVI13Ff
DWnv9KXt0z+YljiUgnk7bTWOIG3T+d4aE8ujNCtfMxrWURhJW8aZ8hWKZTkDKj+WmPbE+JAKHQfv
MraYfXZFGjSFqVIu6TTDKcIzGUtUZG73ttTVVkj5Gfv+NHW7D0oJ0E3vPQRkmzREGaVmZ/84Nxej
XB5nCnvQKdNKjYoRZcCJwaUpQQWI7NV3+ZmMG/ucKj9jFqOgHIIbYj6lIq+tduKIjyxRIzZyu7+p
tRcgSaSPAkiUWP6XNz1tXYzKyB3Lmp203oDZodp3zyM1nuLeEKbiTewpHkBSg2v3VBL9h7JTmR8/
2+hnGapvbgR8zZi08pY9SP4+Py0NjmjmC35mR9ohgi9Rf+bUvTTuNFvD8zybEgq6PgTp7J623VYg
d7JYxdWRnM796q16LzioLDikxAjYOJIJddLZu0f/gT6dCra0NorkJHbdC/D7HalHAC2IsXf36Fjj
XLN1CftVk3TvKNcJqMs285kZj+3krxprd7+TW39WHtTuobzS6FXgPp20TpHYkZqq+YIVj2w9O7Ao
A6ZpxGdxeMnFXc8Qu7Za/dyqSKvhaClwabHE8RBzUMnxqR6B7fCfnJea6N1jpV7SFkYBv2yxtz0C
LnUMhDrVWs9w4GLRatBBnN5OwWZ3sIO6da5RgHteIPQE/iOiQIZIOD/3tfzokp22UIEx+FMyDsBZ
KENwe5ho47CiBeRhrw4I+S0IUj2Hsu8a5Bzb5CCR56kQTVSGnrOewlNxM7Y7+gWUSN+cRLJT2m1Y
+F+2bd8lvyQ4zB2BPFmkBNUO5is64LamEZzkw3BwAydIv0i8crGoD0LK5qS3ViOacu9jfWAExMug
RK2n4PkALAHgD7KGq7/Lks4/Gd3GVqSoKYJRb8GDJ63FJ2YT/Gksx5/xncb6w4TRizHU4iyEnyOE
zBZ5rrGASmtGYeXu3/54iURX4OEXvaIPs7Qm4oHZ59Y9FvYPmavfZjlH0rIsHTqqs3JypHc4LqY7
A8Pvai3s44p0Jp83Hs5Wy84Mdu/DHOYgYLqjQiZE7XVW13fkj7RHVtvgbULsSEpiaI4c2yOJ9EeB
2NHmK5csub7ISSsdKteYCXvnRSJThNrTBaS/0Pyw14xYcIrtbtT4tKJPi0gnU1nZDEcj8BSriu0z
EDV+BKqsckb3nwYEl8g08NGmWjPIuKbS0wX+fGaT/VUTHH8hAntNH4iYYoBzWsQ6B7cysdtquwmm
uKolORS4cEMz4C1X9c0xuOKAaTFXYxJailtlLZeRLtACXPCyYOH7RXu6wZXvbAHG178u+mkrhqK4
c2CROKMHM8KQmRK23j0yjkHwBmf0HT4IB+3zvmYDe7qQeu71r/MbS+cvoDzGnW/nxGlbCpkLMsfL
QBXme0/vi4+HaFIArl/wH95MskjD75h/mZpF2jvime7vjTTM+UAviRgBlvVdXhdlMz73XPBSDhHq
Sb7LqxrGqLecyowQYlrF8e3R+gspbEUDEeVbviTZIBZ90JNnV5/k6lQwyDV5oP4myikqyH+V8ip+
cVp6lfG9CxNQ4hlc3/rtKg1p9/kmIhklxej50J/lDEB4bXqOKOhZ0S5NwubgYPWFoSl97BktM0AX
1Mvwtf2JFceYHmMyifcTkbYQmCRSg5gdMC2EzABQjwEAWS0kExLraujy/5DN/3yZWbnotmvIJS5Q
BV2D8oEhoQbV3GwAtAPADv7kRuKUp3/Hn/l8Jy2+M9dA0Kc59qZDEbCYTF64QYtAG26QsTwEeH7H
NyNGi5h8c6j/8+HZhc7rYqOakos4vWnQXmg7sLsaAeA9LLQwuDbKL+2VBWaximtOUdDVFBe2gzYq
sJApuUW/8DDxcJICrMzzgNEIoKdyU636TttHSOixCYyQj1/+a00dtHoNWASBFjzWLlUZP/ABd3K9
zZgMKYsP2Szs25vMcZOoDHXxfSoONli1td45xPNu78+uMF0Vt2nl9f7exNKqbHkicNb582AqGxuk
0yN07shVRbL5u5xXedMUClZ3CKsM9r9Y3JB/6pVXGHDN/tO+aGYv7A/Ih6W5ob8kBuRn1xUkqR/F
AE5ZdBbYT3DBot5S+9tcgdShZbCZo4PdZTXSyyxCMF2yrXXAvGGGNxUuAFieydipCj1D6EP/hScG
rxQ/gzqYDqm3N+g2HnCYcN5pii1MHEQN6m/Xcw6WwvEHySD/Cal4dEwtpII89qmBEVOK0VfCDnll
PJ4avj09qLoBsteURsI2zV04ZCTGxPsiaCAbQ7hSy/oP7DValX50+X0hWurl16Ho7qu3BXo+YyAz
wR9Dzpv94VtQO1GQ7Nu2REr9ZarEs4f9rVDMQnVidN+zL26s8Bkjt2Z0ZB5MoEOacjB8xk0oeNwd
Qt+f1wwQrHIEQvLN5ge+CPBvBAP2FVk+e/QgJLKB4mkO5Elx60frpjL5pbAj1b8yaWF/MBdmSqhe
ufxb2hYL0vHZe5jeVUQdSZvzuy0V6qf9OPB6q6UEzqVHd5f9jMg1cPyaiTrOz80gWbR0ThTHSOfp
clye3J8XhgDVdIeVKTAgbDtcLLoSD1KCkfssz+QGCXZO5GJZ8ZeW8/z8HLU5JKNg14VtMquZOSrD
83vG5Z3mcA7Po2krFW5AlypDHjlTArnIQhMye6MJ8pVUwFIiTiHC9Rw0nuTKDZwg/Sx4eKRZu1pN
rIQH5CqWe8Fcz0Tpy7vaG2iBV9PkgrN9B9s/KcQ/ypSJvJPBkLzG1NNTynEncpoC9eVeLfjMxBb4
XJuku1zwo+mcoo5ikcIIoZ2J1nGG+IHrYU7f/mci5zGg9W2FELRu0VaTihf1Z5WbjahZzxP1Nfs0
ZMULlKBaX/jRMIYRJU9F4kk93R0F8dK/k+1c+lYYkxwGaWRMHQY89gHfIcb1aES6JR4zopQHihQC
y72dfeQu/+4enrusSdIZPF3KJ46CGGxi5RWLQDIS48Jd24J4hKxsKNGiAaUc7cguAQRjgGBbXqeH
VsBvX1m+EbntTkF8PpOd9cF/wO/DR9rkJ1u6w/4E2vjME1B5TdTpDOG87wCfxqsnxDINeuJS0Y/h
471tnCkcYBbpAAtdro3MM23RJwy7NdFemZwGdiUPOEvEaqvSp2cD1yZ5uKWkxClJLUt05bwb535F
Ffu8xtiZ2pMaD59bbzw4PgkUSTwy//Usf5VIE2Q3nqUj1L5XSPeUbpGAPMJW/ozbzm3VwOmYWgFp
i/TK/18RFA1oTVdeoDrtho5NxNF+v04X+xzeE5eJVQy8C0aWoZoc/WEBTGKaSEeG/9nRoo2NSstg
RZbc+AWw72zvzc6Tc4XnqbOOUrTymVlq5jtFGtKy4v3Z/gHicUkVpUhDr7d8fSCscwIUNgg7bxuQ
vqrzm9KWzRCkYK2If8UP9Rd7HBT2+mDprZDVrdjRpZsJXOkIQGvuTP35AahQBnqgQP8khcTwAqgj
9beDp6aKa2iSWE5eDn1iQ7CkNjDfYSnr1W5dpmyRK87kh6DqrNSAFwgHn5cAjPJLKEFQLy+uvC2w
I/CeS5Q4a2q920SWuu2uz4ywvyWkHrPWHCd95hB6zSvYY/aQjpAiTdYKzRTTrb5cv9V0DDekzzAO
s8kgRtVH9RmIQig9IhMRlkFaNhBw9yvAQlx54Pm2KZErZ8/bZWUtMePdjhzZXpK4rBaYdVjWT3kC
f/6g82pR29CqlRvBdnIfjIahBUX8mXLF2G1cONCJcOzu4SzrT8FZCn8DPqIindOxt1kKnY03C0IN
P4A3xsVQHynZxIJiboReCLq88CBTqfB6Bn69bnRuXBP62NcYKD7bgIxp3kDPFsDvrdjad4Yd74BP
bjvyqAnJR2NXaoaqxuaEhfJvmuuRQbVt3kL21raj1LlTJXLx/FJ4uevqnWZ2/BoG85DlxEMYmktE
xN0c9fUUzcmVD6WGmsSG3nak9ItUK8frseDro/2Q8CgHPJHMeDGIyUntlVUfilt5yAGdXwh82mM8
uM55IHJsZejXoCpy5orEcVdwvCEmTgnr5WM1xMP74TOj5xS7dXvur+uFu5Ib+83BlborwuMgM7hm
CcQrFiLDbAsyYgK1iOgWzvDznnaPavhk8hXFDVaD6jYW1KA8qGHdZBYRSl13XJjd5tDiRE+/+iVC
seO+zAP4R1Ql4vQ8k/p+/SD6wk9cZK90n/XF/mzrEzkhVvCqwGdWqqTm9T9Sf01WR/SHUX6p2USv
YkRbU5Uh5iifKqV3cdup97PbRmpDojnVIi4WEhhcX9Q/Wj2AqFzIlkPlYmARh57NQXAIUSK3MHdI
LUB9HYSrupXGW3zu3Igqp3gptoPI57miLIqu975pYang+BaUoikHc8UBH3eEDcAYoYPTF+g3g+1g
Pd8kdtfnzviT6xL9wiASWdx8nXBjtzK6703XOJV7RwO4KFQ/tjHFi7hSTGRbCyiSTE45lblmZmRv
eXoeNidOexfGuSuWFMckvfa9RMn97mlWTTn7XsqfWTBLQ/bmsDURuuoK5I/mfP/5khhw+zF+uQdV
76b/OyPPBRoGkKBmh/qSK4hevaHLfiZcix8xO3Z6Cqy9WDVXPJ4tNTisfxkuywXXWsrO9Jpf+6KE
WKS1s+F9wii8rhYRnGGcb4Lm+XGrTNBHYL98GKCkoZF8T3S/PcJGu6yNJLbi9zj3MEJfIKuAJ4vM
L7K6D3N4PNhTpnF/FLK7PUHyujtRmnQGqG7Mh1ox54YEZ/P9y+sxCbs3aXzGYBdZBBOwXL3NPLN2
4cHfz4+atFzr92tlfrvGPPXw2DxIIThtfDjSyJXLiQSFFsdfRYHcacm3FNE2wcfeaL1O2qnulKTE
ERjYbOUSwhrT79LRvCSJOMedUmCgfC6vShlmtdhVEkFk9H9wvMWC1gVF/7WXW5HnAxh7droaRcUv
hVl+fKMTZ2ccOFHjcdPnfkrb3Wab39PUPVvEXAEbmHBv3IEwGT278XolfH2in/SgLru18cajeiqF
Zo4apsJxbtnL18QrBzHWzLoid5ChgNi1wd8r7OcO8QVTP962WVNMJuIKbVazf1pr5oQVh5/+KPQM
CqKtCdqPFY6stg8NTXPREs3233jz4mQI1Dt5XPSHCoxv8PIPs+fVmMiJAzDV//u5/dbnR/KxgZYh
qwpLqfOzKk/RGgXlvqFjH4mo10rGev3n81II/xm/uaPNJeLMqPgkSvgOoH1cQK2oPnvSz4SEpO55
SHzgSZ79gftDJknKfLgfDyQzz0ouDtxKEH/a2r4eNHRzuClCoATDqigKadH6TxD/2iD4WAXeF4Bq
tkfWDCkAssL7sSyHPEZ080x2GloTKw3yUcBxEEBVZknwSFnYN8l0gh4lXNK6xp92yf/o4ozNWTi+
mx/+FLGggfUbFk3t974UAWjZHY/2KZ2x7N+WkOtuBGwREGXJdo6m4lvXA/v60Ta4Y+hCjv7oksSw
J96ffHLVSOYRAfshw2Dj5gCTVKKLa6a9UxhqLgxwmti/8JZ2iCIlqt0jfniGT4WdMDuk/thsCHGE
JrUqVO+ufxXy/k1FV7mxib2XqRYBGX/QLX/CW+6Uyfq5SvnYn/CUziSO8fAY7fbbs3CzfBWonF6k
Zf4F44NmTBerrcY4gNBeQueEjPkVoqlaAfAs47ZdZhwuOgj9mJ870oLn8FGOnwgW/sxwB0DKo7Rf
MDLgESwVfJMNuuppqX0tdzqA7K+qnP6O75ePCjc7qBWHJ9iSi6hwJiH97VShN3dBJI3nP8HjZn/3
INRtPr2X2KkF42mT4Vy9HT0lmfXc7kULorcM2v36qtCn3p1qczlvX6sZkYvyKpxwjbIqt08tv4l8
0/LMVGsCN11H123j/xPqFyv8PddM29I/SfnaqqQBbyMXz2Et/QBjsytGClmqhd34BmL3oynDKVl8
c2SKRBJjMAzIMucLL+/oaTGXHOwgvxbcHdt/Zctc4yD/p6HlXbhTHe37lf7y1fYgOw4KunZ2oRwF
+FAj6NsQtCbAMTm5oUxog9CgeXzcHlimdci5fHey5BOevEC2rBFG9h0FSYW7c3Y+BdvUlj6uNp7p
VJBsKOWQG9HsbFbxLevwYAMwho5HxW74BBT5790thZzUz+nkkcds/e6F/5rxUfIUxChiM+DvLv73
zjige3MIguV9bVqjBjh/ej5J0MpOOSjp0Abd+y1mSA1VpBWARcDBGGpFkORU3P+IJ9JT3FIawigC
KwW8LZSLhgwU1wwWFUHwAmUtaXsU1jbbSZ1B57lHHuvA+Ml4JtlNtapJ6VS/bbhZKSmMZHXDGBDP
1qjRosbzciYq41Jp0id+uzgnDbKtFFDH7/t9gvpknZXYW4nye19qNE+YZBhTMRYPz/PvSOeIgBc3
nWtdnVYyE+RcRllqdtBtN86w/a4v2W8NI4XFG8eDTn9FdSL49luVsWqld1RDoI4qHZH0aByWxmAH
mYdP+pn3JIGgzjbrRf41wRCpve8jBdzwRKmTgcjP+aru2rMuhG+m2m1Bi/M2CIawNB78TxpMhAar
cEob8gE057AW5FsOr357n8887RwYMIg4VqPoq+o/I2yGrew9+to7/FxE0zoQh16ZNYiY9OuaZM8F
GyHNF2uOfQ8+xE7wel8hn42VzW0dSTHSfpODgvnOxF5LA6tOGAtOF/iMkVepT8xjfLD7sWKp1JWJ
GrflVLnXn/C3Qxrp+SB56NXh/fof6KqJnAAXQSqFM6VqOvb8NiNpNwJfsF++gqY3govGfEXxWFLR
lhO2vb/n6/j58LtkTZqKkjBJM1sYJapU7j4NvXRE+Mv63vzm+tL9B4yAx9yI+Z6onIYF7/rBNDj9
2rgasb9wMa8/oxa2xv2LDzU8cqxJvUStxyKzhxzRd7sZjqmaGQdxmn8dL3CQSmVFUaDCVcT7wO23
rG89TICkiX4+KSTWmiqdlW/dgP3xjIO3uyRaOrsNQxwgdzP+Ya1RCVynUneqlpO0qpCtOXRC/cQp
+Fog8BsUvyTYYVDRjMSj1ctc9hzi5V0juNtFT73WZ+SQQ5gdg/9fX8Ec1BVXAnAsWDcD/1Zdr7Jj
HRYvh6soh1JCamQ9kP+1PxI0G9ZnaaKgEGNOQImPzSmgwCcxQoaHt7wQmc8Bfi3MW3nr1jLQWJjs
CGPLy2Eeb0znV1yv4dhN/ceOpYM8xNmf4/oreaO0pIWoi42TSe7V01tcTzXN7icVBvpQn7QeJ4WD
tBjpsUYweGYRwLaUxZArb9kH9AwU3SXLqqL36fb9fnnu+H1SzFi6vJcwbLn+hWcGuPD/XRLxRZhV
UEUaj1SKqXjx3c+9ZoKmXOC4skmbXzl31l6uFJuLaRVcQgbgWFq9vFNp248yHLRazFtVjpH3Pd9r
aCBYB0iXIIy3rFbLL5W9+1fGdb+Irab+UyfVvRzX+IrjLXgVPGDHAL82uqEhln6e56mLg9j6VU/V
w7oiXZuZ08K/k7Fb3jze0yZduhttuqtRJN679rCRPJ02vZBqCJrjbedyTIuvPOg69BpWbcVezu1b
lR5O3KxiYPnxAQoharebyiSL8pzAaPbSSewCNz8x8dNcx0KX3H2bzObrHjx1ejoOhpK9Qfj/7HYh
3bUfx8WC+FpQkiAAM7Cu08LfT59X6aLvIPQ4XZgC6xro66rpc80bKtSefgimYCcUVj2Rva9cC67v
aHcFOi/g3mLPB1CG8Ob9WSzG8u3sdXiqChdAf7Qjn44yJQ7Ya60U1rGaUOKryn8qRblLWZpSTh53
qaiiWimr50Caq5JUG/9B6ySmzABhAchPxqheg+WxngxREL9C2luHWk8Acr0X84nC0vnkrxtg78pV
2jP3CF10X4uVz57/EB+5L3WOKEK2KljZSJQdczeFDRM/qPWGBZttMyuM9C11/zvObpZP38JRm3zf
WBjGjKd1kLTS+58kM32oDRnAxlAD4wtU0I+7fXD6kE0ybR3BXZu6Q4g3v/PS79WvX+YfrfA6T+BM
hwiI9HqOQLsgo6iaX8+1EY5bkjFdySdL9j3xXchQ6nA6x8mvKISsnFo9QaAcFUh+kBStNxeaebJH
g5vGTfdzx1RTICRR9YWTrTqk3ujexC6d+MQDfzAuMXVlEqM6OFI7243gtzFIBk92jpJj3yVN7kzT
Rg96zWpK6UIRKp+icDSRy6X2hj4XjrUL0LSWBYW/ph0lIi7tYHurvolvu0gOgQQWbr8l/kX+FQ/q
23W4Bp30z9wyWtzeJpjoKe5pzQ2xIHYPY4jMpLZxpu/yysvV3sWIMd7U0ZMlLyRoBcKxkrUZogLa
72GaGaosW4rAYFinUPQf5ci+WzMnKyrCqIGIbfsNzO0WzoeHHpz3ckCaaE3j8rixDU701YUE6GbR
ZoWBiP3faZ+DtR4o8hXnuf21uePi+EkgHBHbicsd5HVwW7A8IYti891hdjNbXKFkK+/T9NhoW868
Nq9SbUU5xhjAWk3ANLZjX2I04gDoX/hSSlAuufNcQuU3ct0G3TFud+T5ew6WgG1iVOLkqDJgwR9k
kzZJN4CTUbmlMp4Du5UA2blX1+/dmZosZzK1TetTsLeHjeO0EYPfUtb1BlbJ1dpg+394p/XhyCSb
M9wF3iEU+bNxIPnucC4h/bWeH085HV8a4F1cItk81Oqg63B/K9oIEh/c6z72fqLfoBggS3a4aE3U
napUjLzIU1fnyar23W3gbQL89MkFvK0ekSth71rRdyph21xp3J36mo3cYZaeKKnZFFyFtsLOOZ7Z
7CxUC+Jc0+ss5b78J9g3V69TL9LtjxcbYqFh0jNtFlH4XuLrG55fbCmrTZGmqw1uYl7GohOJR36K
vRf9poscQaOSmnWXh6fhm/FFey84eA4VgEj299GfmJm143DNvAzcbmoE/dSe88a1By2WS9Dm2eyH
hGI/dwKa0X2m/lcY9nFFn++OOlDhBGnLBaVc74FYhn0flho/96Lb3tLw5G2s215rcM436F5jKOIO
ZicV4YDQmE82R7Hy4r15VMJit5Ci77TLgMgIoZsIRLtIwOS3a2HSkHCqk9M6fVTOa3CXMTfuqIHc
XwbfnBNM+nhQD4J1iIlgYTfMXGkzmMuXnNGH+fTkpB8OD2c1ttQY4LzMRdJna+n1FaTATvVanB9N
lHEwe6dj1rBWeqYiim5x4nKzTPNOxfICMAdgqUlRw741fCro15rwHhAmdFEktmhlICxhMZSjalmF
ocAkByWsrgNXPUEVRt7Q9PdvxQJhxrx5lRa1IcC+anTGxEt5+hkuktvrgJUJ8+fkazxFrjr7Er1p
IPxeqHBStRqgLCgqWfYLJNctvzNFHkkQiHrfSb14Fh3PBdXOd62KKDjuOyEYIPCNIK+FgFmGvI+h
RJyfC1NtMz1yVInBkrLyWgCb/vEP4+COw36pS3Ig5bLsn9ezhzjXkdJCr6wNvpGXyonCjRzNyo55
rXhdo7S/y4u4UWDM/+I3TvdiEUCUbyWjra1KXixOVzU6GVBPcYUE3HAlMvCnuytfp3znVEIivp1E
ZB7rtnMHM3Lg22e2IkdVBWowb7uLHzuCswBoAVz4GzVOaG0fGlVdhoeIC767twvW8Qldf7TOKAcu
JXK9GXbGbFVLfXo/fYUsjsiEWk9pSf1bS5KegxDlJPFE6jVZy04NWQiz5oDcXH/qwWYj/HDSnCis
yIBFmx9OKBzEUZdAK3kr0bKiySuyIPSOfWLD7WD6AwtNN/OWS6XHHaxsnmsLjDoIX8/erFdIQTIq
3QdMkUMsXKa40QjyPSHQbiLdEq7dCbwqkOhA1L0Cab3PnztH4OOe3BuKMnKtZaxBbVkUfoKXRAfv
2yVGQTt1soKPJJv/Z7nwOsaSUk8qFzUQepsGmBJAn3CykLFi61plDgV1scHksibr5+rvQ1jEllw9
+rORZm8xOvG5vY/Z1JHbiqiSUEDk0288bXbjaMZXYw8eZY5rTN2bkTSpxgy0TarS1kues6hjBMDo
sW9ttbAgCtQYQtvlaSxd4qrwQb7G5cc/yUUWipE+soy9tfnsXrj6Mka46mHqOpx7gBghKeUgw6Vg
t2EWgaambIFIWkRvN67XVyUiVs8PMS6nIE9iuLp5ZBPf/VZwVeuyvFzchjB6nf73NYMrmib90A6k
RWbmW7+9oxqtCRygc13NPtvWkTc7kkIJ80mmJsKqoC8XhfYeW88m/lOTcbhxoc2t8RgcNusibJmJ
POk+hl8LLQRD21u7dzeIdV/iqYmgsEkjo8IrgFEj/CXyA0diF8VLtOW3HkuulhR+YwlpflYVLQ1u
Jqb+C0FhmUbOQ2VQNFHHMgzGo9XRlEJNxkK2+bNyoFF7FaANDPACjGspZ8yrd1rMV+kzwwF608ST
Y6eee46neCfKmQ3I1ce8G19Ljm8rYp+7ZaLqLwCGfAtICJM7v0VokoSkYxdXX3eY5Nx0uQPzHwjm
zFFXyzf//7UbHbgyQyvpf4G1QjPmnTg6nCKFX4boblcbvFdk+bjRJmJfOir3jrx3K+Kh6S4TvE5J
NH5DFb4ytrwkkTwGr0UdXRUNqQQP3KX/FrUF0DIoavmNyjZ31vFe8S3dvNo0wgWPCoTa39goF5P/
hCCESTMAlyoUNmTHrdwGs74G/quNJCcOAZ6MaBtnZyCIEhxou5HGjuz1PKBBaKCs26rP9REH78GN
MgRawT01aXVcFHMvwvxA9GlPCZIr/Ug70rPg6ypn/kknPeWYgMNT7cYeiaFbdRl/B16lDel/J1qS
gLOhwRosNnBdQjlveqJl2IqDfL9IBIPrdR2qj3VBA7bgJXKYv53nwtGa0JqJ1wisR2jIU4d2T/eO
GsVkKc54Z6RfHlMMrnsrqZ6Q4ahkApKT+EtrkAZNiboW/CMs4G2DghgZ6PeA7cI+eL06trziz9QQ
BZfChYwt9FLskDEzBFHLoSi2iHG/g97GINOS5HSl1QIxxrK6M/sqcbNc2gZMWFhsXf50jibt3y+T
1Wj2uZ7B6KH3Z7Ud7Qj/6wB+bG/mw3tKPQO+J5nIK4m0Nd0nIr/Q7vASgbfw1fefhxBjgdrqvIH3
819WldEUUVY1pbwnmQtu+UwRno9CGHrwlkhz/qUMqDKddFvXpcIdI910z6N+p3XuNMm4vHx9mOoi
PaoICAHQRbg1V4y+N0pcSclLXMl3YVZV1FsdrXSWX3PHLC+UoXDbUQOw4hlMTGoaIjOiRUx8djtU
fWYykuNcaf72OTnUdX6YMcND993BTgoL3OeLNVwPSQs01Hp8pVMchwiNHvV7a5avCg+7qDhZsy1u
XHEI+xsQ+uAPwmGbbeyNp2VeIKqr/mNnNqJqdYStwO+yj43KQpIegeTnn7vM2iQtwk+7+7/oLxrG
LxP0z8NR6bfCtCKpMYjHdDJmmt6aL3gaewP/h4v/jkZsbzpxJGKrwiuCHVE7Qr2m2OPeuZSpfDDb
YHRDLWZxr1Yqjz8lvxf/JRsuwJHX4o1rXJsCh3pKndiYvfjsdByRI7LmwThXb3GfAFO80w/vzsLz
ya3tM5CnYIk7TZzuB+B7YwwKkux/ROLCy6V66XAm+OPBqQoQpXuR9jbiQ1I1GEP0e1q+QzbORjo0
uYelYJXm21iRGr10afb1k/h/XXWoY9IZ0NAPaIoIjr1N5KhjkkluMuNIxE5Txv/mqTRURP7CcBo0
whXIAN83mobOEQ/tM09shbHwDrcwmsBTGXRdM2Ynrym+m3Q5iN0ynNU7/QbPxQXi0F2KGBrJ/c9I
Umfnf17/0FXunMKzCqOsTDBFLHX2+RkI7uGHmTU5etnL7LisbqnLAmEVrhye5cvCv1HwNnNhjNmJ
EdTjqLO0xkh/M4tJ5wwjhNWPwgVv3u1REBrssUeGJfAdpa0dYui/37J3wxcVZ1qlrMMJjDQ5qU5Z
28HNvIGqAKS5a0Cv6dNHuufVn+Ef5lTIFzR2eMjyo7bVnjF/VYnWn6w0HJEcmxdqaCPOXgM7akhR
RGyizhSQ5xNhLQriOF0b6WIUcHNqahqjTUYGb/OlbY6a/Ok0HW0ZTuhEKZtc0mPRIeaa/ClrNAz4
tzcivB8RwgXzyKZNaQXs6iEOXyyzHScaXW+4tp2LxWn0q440xo7Xjo8KWmbNxE05j1OYSfHBUHQk
U2G/sxzWG6UF2btxUYzQ+41b5Tj/ChgaWEsv8dmI0LZ0bXAmPCcMxt83Oq9MCPf5Zrem/DBmkxMH
sNxRYYF57cPWjJepsz8D3B0weXFoN9axfC8s3wyHLsbVetZbmWY++5oGmPRPEn4oAHtDZ/cGeVTC
9xr9OYyMvCA37CtrahpokDAnPhCeDVW54jn4nMlCjVeA+jIqOepPqjq6UxPaUlurMYxRmbZ3O09u
b0+t0skjuK5vZxQKHBgzQNFMi6K9A50Bpqv3oLL9BHXLYj7YVViTz+s/SwDGoOJ4alJozWl3Qg43
SPX2S3uwiB4gQv/NQ6SfFGIGV6HfH5GoiJNQ5GQORqNkx+apIIKf5BwXtelTNfKvYUIDBScceT1E
qb6D1/3TUGDCwZvdzLjoSPcPm0mun+R5luc2yUMn0A5wUs3klMhodPLo52/MiU/ESi+BW8oWDzmt
PCM2mi5dstWu5zt5e3yFyrpcALQh5Jm3eRj+oyoliHVF87Q8nRUn+l3YCLN3liKwUxgArXy/C4aD
KwN/zkGRLnxsENivxCOrcqa5IREpr+xIsI52F4aIOdsbKWlOt6P99ekbiVm84W8mrJXwgZGaKept
aV61e3SjWqODqoCa5seSNaZTZP6h6s9o3O80cHwcEfTloyhGQHRBb1LzLVLHhAtGxK42biOHrC1H
qqafHzpOnH9foTWAG0k0hkpWzR8yAqGLEuenRsotltVPm9KsmKhWcbiTEbFZocFh3nRCBUyhC55P
cKVLXESkyliWj8FbbOyGrFEPkaf6WH/zAXvm097J6RHqgBsol5upJmE2PzPYokbLlkVxOadZDV6J
rKCQkUJ2eNRCHi4nzpwZPZfs3Uxl9i/t6yqskA2ZCRbQXsa0p0lzNOx5UNTAYivyeqROMAvwBncf
dDeDlhcSg9XLZdNmbeyM2K8sv3EtABei7P6dSzwuPAOh9nZfYvXFJxeh51czJVb9rfkDyp8N/A7G
vhmKwE6N28rMnoL0Q48QIftKnyq/4K8EbTR6VfK3nlDBaEvpHbauUtx8fdy5e9drrEcZ79LHbFTe
oz2oM+nAx7zG2m6AyO6pw25O+1veTwBIHJ7CRcDQhLdQt8aPtWjcIooRkaJCTXmOrgJfjnbNnUb4
81+8ibh0q0UC0de8gQ7PWch6GCzSyQL3MkQHI9wJnMDgvMqkWdVkPqxRYYIkGNcdQCfsORcRmn97
CEaTCktGz1Uh8ybvbqSpcY1sO8J0SpFBG4qZILrXdVFBFcT7sNTeNluirdMSdYZfPxMLF8sqWHAX
aO7OnmFtKiibJu4ihI1obieXqOK/0FsyHfxWTEcefdLrxgmePTr0dGPPxTHzntdql4onpR6LvboD
8S6LNtx4iXU2B/1d9eGezrJFyl98vYffYJEltNmt9QxxXEXI34/iE3txyufeqR8yGdshfYyHEtYv
hyXUdKOvt4CD2QfmMUjGkfept30o2MaoaKRtaHTK3n/SLazu0nIUPaXVFc4TmA+qkXzh57M5i7lx
+sKZ+8FgkT/tPplbZMwRhOxX0avQpy/dM0vFVTAj4flc96E2GndGrmX5ELCWwD4dp21zm66FyEWw
8S0bHxeEKGGCzYpNq81e6KsQhfnKjZy4O8qB7ZJGkE6Evp+AbHkYTK3XqznXbg5Esx1aMp1mgBc7
XQdvqT3cRdVPHv9gBfs2A3wzaR5zrvMP3PP8dp4pUC+oZQcC+gC7b/4zqZfK5Pjc6Olu89ycl5r8
00lpq2e8IDASso5dCLI1b7WEvPYnIqu+XRYE9GgvE1yXTxm62ZxMmF5Vt8GHIadAo/BYGHF+L9Nh
d8MrYAs0GnRt5MQXj9VeNZPUkCu7KrNP1OSENSn/RlhgzVBqM0ab/Kr8pjhwefnWWBFTJg9S2nG7
nzUKFUr1S6eA9fVE++7LD0u2pOxzT4I2why6B+3eJOPxyni4ji/HpPYY9fjrYr9/JLSPFgl5BRqB
8RzuuE4soW3sZILmENTlqO+56hGOm3cKfvGGiAAUZ/VWP4T+4CH7ToB1pbw/EzaVkRToKQynpHd9
73q+axIU5fNYc2Njf3zCf6dtvDdKgz6dkbMtMYwO6N+y35T+NpVHAwxcdi7ATGT/OsA5iSXjTdlW
gGWSaKGP0rFHRFu/jmPHW6O2IzmcT2QmsBupxL6HCKnE4svvIkYQeuXpea599c9aX7jGr4ui9KHO
HUlbXLFozbjDhjYBzPfQBeA/gyoOpwq5Vo9bVKUfI++WX/3R0znGZ849oYIuywqRBLzHAwH1WKUt
GguLXeAuxXGKNFnhL8/NkBqrE7dpS7tkblwP6PeTyChRxiRkmxzn104OSoEB3OnLDkJr5P9Y48XH
fZwC253Dw3vYTpk627gvWAChicrVSqQ+wDVsv1uH8OgzqACaW3fZF7LMxreJMU/hfdhNJzvIlIZ4
W4QmGg7yTNegGa1N6U4WHodTojn8wZCErkkOMzUPOfUxm3byWVA0jo3QNIWHSiGG5QfzYorMqpgR
3zLinPR5qfvkGAAD9XTa1I8ppOTb6vVwq5uUOKK/yEP3DmL1Esl847nfFa4uRTT/Cq6yfINUdLbC
UkvvOxgC5/NXVqw6pBKpMQv75NANKoA4cE6KU+U5vjLH6XBMiEi3jd8EUqDB5smNeLm3uHHW7DmJ
wArhVDGWiT9LYv6e6jPFVVfS6mhETFdvySVr3DMKahms1kyE1mwwXsjJhwUcGaJLPbtmm8X8wKKV
as/iMvn2GYSE9afr8w7zXao8f1njf6WNFjGddthAF089YiI61L6JoHxljQkeJJZCIBA/OWDoiws4
FevHu56MZDQNuPhcCShd99TfR6SEQCxydtE4FBrshsspt9uvp0tHZ8ZlO1GrDXTZaYnsc4SjDxTT
TUB9W0IplLyO5n7hC7pFbH32aoW+LW97fXOjheH7QUQKQDQK3cL8fdV+SZMwkJg+FDKsGKCTLIt6
H6zIUGIwIWDckaNtvRmkJGJxAtEtm5ooPDSy1/N8FowXogaUNiunMcoaH4ZOxy2Gr3bKHzryd5Tp
pEiTmCrNKMQyI1N2ai3XRmg1NDcpt91YcvHyC2eLKs40VhLSbfutUheEFnGkm/DmRz+Mc5rVf+UF
g2a5W/b5cnJY47WK7ic5vV+ExMh8qHxb8mZxgv8QRL9zoMrtiOJWERM/ngALS5buay0qfLgTDvyh
mujsHLg2/iGRUXdSmcXSzahpWWjrJ7ZSYNy72evs884VyalNhTH+ItcuoFTk15fT/9SXcsRVQvCD
jKQ+xwD89rMfnqV+VHufPI52hbGcFnnmMcJW2dPK0HfdiyK4oQT3DSO2rSA2gZTkuqvu+hOAAqQy
aylPUzplBYa0P7khdtz8k0708yBsnLXl6++90jPodmLvwEtEh/2IT/I1wEmLGqXr/P6hxgnT+BUF
fZjVqXV4joqYZJoKWwG6LZ/ktOrT+b4poxXmgF4ak7kkXZaUvkZfuWwEFy2RYO6kWqEog5GaFNpV
YE+GGjbiP0DIxzk88SZww6cTJZKk98XESnJpabWZQFCbm3nhrnuMM0Ggigh1AVFZmTCKPSSEN7A/
yG1yaxZOXmYRjxfYNMgKgRhAi4nLYtvRE4ziK67/GYUPqvQsCz9Jytcg2o7EhDyvVU1d1/eHKiwz
bqWKaZnpPShbAb1QP4z61ZXenyVfL61dFgPWIvpDJt3TrXWcf5BN+FTMcT+QxN/OGUmbmuCSwI7A
Rn1caJ+1oDXgYlCrtIMJl2msJd67L79UW1nguTJ/H8iRtItDHxXvr7lXvzeLBWMjltCAwhflgiLr
hZsIXzyidiTz3l5zIunWnw8kHfn5WKM44rG0br58sqTLlYb20cBekcTkNHVdB0tSasUKlKVqFgXk
hwWwYEp1QBKPPrg/0hZCYG78abQrqQWTj8SbNtNE2h5NbqfyPhOLMUPW7DIEm5pJsvAS4Ie2AslC
P9CT0nCwmdjhS+AEVyG3Ib4KajVFMeETJ6wkLoCSfbvi+eKWBuf91cwDPPRYECoFUFbYeSNg6hbn
akeeYNBMkyg74bTWshc2D/+5m7xkHcLqQc2hJAdYATlZsvGiZ+4j0QeGt5UMXKtIdbnYDyJI5z/I
ydH9L23fCloUjYE2rr3v9dr5+8q/pRI9aQRm4lhlKSDS+1LS+gDIdJros2wAZlvrbK3Dd8Aq8ba/
DN4iTBGCxguYEQvmohAvgnc82bfc4ZBmPZ9ex2jC1nM7MI72nkGxjtWN9SNmyLGRjnbiDLZ4zCzU
BYeYJ5jLPwgoBY8HEI6n5HK3VbWmY0l9T74uxsv4XrQ2aOhRg2NPNwgb2iWfRImq1fNzzEDaRbDR
96W8D2Wdp2ZNR9ah9CfV4YoT92DEDzs5kXa8gkbni1ntigdKKlHas4od3iUsJ5EOJ10YiHyUWetx
ZIBgMWYFEa5sgUhRcxG+I2W3cg9NgTZQYa19plzByQ+na0UeNVYOQUNxJAmgsF4ekQE8s+wEohNF
cNGYi/kQ32hmkSIcf8jzVSTwGBrvJ9HHjz5Sz3ax91gTGKEruoZpwDvYARBeAkgc1SuvVoOXj5Tn
1ucxDL0Zr3XOtIIgSYnRuIO61kKx1axk+Ud34gY5MTJuZEYFaM/jDRo2Al6Jxbg05jY6GNsnN2AK
Ws/58z8DZDqOw5Mwxlz6qqu/rSElxYne4QeA0tN5eLTumhFTwiBeQlJMPsVJuFQ4sae28/cXJaR+
LVAfQUEcacPg17QJK5nQhjpzFlYCBwGOq+16rHm01Nrn4fDSFu8EHSMEe5Xm2l08x5SHTdYyU1aI
uSPN2++vBYMPWhr9sTw/Ao4WW5SLzHxVKe66a2y5XhMljtxfE1zOuOxWxgVyiJ+QcbqjNMiDxGzL
oaf6chnzfVFFl3tRh7exK0kxTKz2REnu19frb2/WIcrQdWA+4CipRvmkKUhAqno0iqRqvfba4mD/
5EB5sSDtFkAJFEJ6AbbgG2srs0yaKRgGhkbLVwsyOAs02uawbfncmbHjqr2w/xHk776PU6jKCCRX
1XnBMtJ/7ASgFzxIvRzt66yGVp5KpHVCGvKwlOgBL4Mx9n3xfORg9+6JmtK5Cc0FxLIsu7AaUsKF
lDV49edgfDWIhaYeq3sJWfQrYcm8Gwv85hsurrOyfNt+WQjB/tcjRCh7KFgjGt7lv2kdyBVvRWvT
TzfJocu6mZF3tKhFhQiShpPKDl4xC3dmcNI5oSjI5vYqYyXCmwYDS/Zo2pmJaCncCd5Ywq/RhbPF
4EHdrzgO4Afh7mbWPCxfsrgaXeP+AXI0l75Z9N9pjHvq/eybtY6m/uIcnJVIBYzhw2LW5xhZEwQt
Q1ECwp29KpqnhIqBfLY/O2to/Jp5V2C0/b76/7nTVdFwyYFT1Brg05FxVZdzu0FXhVZvHBIpiXVZ
2r8+onFcK13X+UK4Hdepmed+mbde8CNCFJvXdLdiPB5pk3pK69bd8hggx8XRoo20jMzdFdkA6yXf
iaDftHaT3wQzPojIdKpoj79YIWS9q1b54jLRVHdaaY70dfMvHdqupwq3wh6QtMlUPmevJu7/AKmq
H5dz+BhCBf+WH801LYWZwNynfFpAbmD4UV6mmQYHo/TMCQw9BGxey4givl6YUUOLwCJu2oPJWd5p
UDdNNCQtmAJjGK5mBG6hzGqQvvs2MUOhZ3eeu3eeRo4X58KegsvFCHf7Xd2SRjxQYrigVPSRrWcd
/AA9G0fWYGSBnv3CxS1nw5hk59lE8prgE8tkOqneE21mz/dGT1Qe3qjqCf7VhpHe2XlKU67jbbRC
nOn4WdZm900/EonyWyUtEEy/4GXsLjhN0u09z1jadEQk8d2oAWhMFnMUaNS+2wI06wAnt0uF1j1N
kE1G6f42ojANIGPSCC/0q2unrzJh7ngGRZkCR+e/z4ZfcAr28GCIGY4IcvnNZ+PCiATM3nWBodJ9
7HHqdp+cCgtiIQjJ5PtiY824SPu/lkEWCTPnu4sKvnI+QzzjnXx4HqovYahIZ2KjK8sqKzpsnMZm
swZqQaeF8KTVKKBgxFrVyGi5J7jK2uliFaj5NMPvq64rSLkU94Cdfdup+4kYQMpELEOhFw4dGlOw
VUfvSOGuhNfDsK3I5idl8YHRb+MwSQ+xhbjjwB94ogYAqOR6G+WJ5pQ1TFP7dMnFf5bJB2TTFtcO
GcUBOlK43cJcFVo7qJaJR0IBbWoHS9DB8xU7O2rlhV/trNiwUItriCVHs0SQgQDU0U6uoYO+bu5l
HUwtvbu4RriAORv8egvUHv+Uqjt/JKKrAIT4mtbqFCWOmJQZfsW/rK8ptjvjxF+3lS8quN6EBMxo
QrlU43h1qq+g58OOPexGgG18+y2tErGEhbTiCLb1L22Y0AyzZYRypTi5eMCjfDUgEstDY8HtJJYb
qwG/QXR63HNoJGShafpgOte1O8g41H77Pruuq4Jzhgm4A8ZsrooSrGnY9mrgl0zNCmK/1BgH49Rk
KVhwnWUjquP9o8mB2nsxV2qdrcRu5gBrY5Gj9oGZ7cYeTiSvASoFgvEHoTNBbY1b+TBUWfA7KBOT
S8pXfTTSOX5L3FJXLHqW/+er4ppeM7QFrmJoyYcn3FiXp3RUbjt8FDj3lRkWK/F0KLmwQ26paidX
U+UYj+cQ2KGF+CPDQZolT1fUSaEcNDhEaY4rXyKgtNo4tceVVynuZTj7xNi1QMczQZSSjHhVcE0y
pAz9d6Syy6yK+pXkr0Yb6Hue36hdFvPeo1cZOP0mSfjKUuqSrGCpdmRJuso4F33qDfo6bEW43lQ2
DWEjr2MzczD/m7wyna36SAarvSUg+4QMJILbZLCNOADlXONtd+qE5v0Xj1Pny/hmlYzitNfaKX7k
/Mgt/edSgCiXz9O8ylvaDc8amqrmBcIwS9xIpE2vVd7YJXhUzVf0fV4UwQ8brbLNyR7MSChfvXBV
q4ULOe3Cr7c/4yJS4/lWjD5d3JW4tgwkVuPA5yyww76hG0Baxt3W6wYlfFcRIKhxQtbKtlRqpWcD
OECUXBdLvND8wVscn0/OCVwMK4FNzkTK92GgIuEOiF1uXzYjJ06izPSsiHwq70719WdOQNnTM0LE
AuvXLX1Gvwr2aSQ4SNrpkeZcb23MPOWDeB4lY2wyhYvGGZqqgm/EAGThcagIIIxs4XMXy6P2YH4R
7F9jxw+O/YS1s42RXBEgQb0XVmGADFwRWJSARoXdGdLIRUkwHslcIfMMHr02Pzssl0G53dbLXBHx
S3S47bB6Yd23V+Oq9eED63egeLbuAcBWXhdbFNX7e1noB5458NfHrGPwN61+U4GeJw4yC6v+eh0i
SIg4ahZqFAARN9XxrR0bMAhnccmBEIgMnXi7GGVv8mti3bE4/SiZnDOAlA6LYLbuzm7uRCe6d8Rk
k6I5dYJsvAleZHVR00xZyDUUMIRtOAQIvTMeyNJnA+QUSrKUEA78IqykH9dPNgcJRHy07Y4GuV3O
haXJ9nevmoq4oorRTy0N0vcvBhgRWbqOcComrZk+anA+mxfCnHzaGms/7lwMm7QoxEcIxN8uPTrO
/fH7ciCjllWjcZawAsIfzV7Ki8li3/7+o+6PF7v8SyX1vzJvFPQHZ2l+oi1x5Qc/HKaVcvJ7aBrL
wZrXxy8UdtKTIl2yrFZdin/E/N/RXKwA3bMJSrEW6JRHogYoU1J7WoX+3bSUD3n8000upNtdb1nh
xOR6I3hR21VZV3+tIfgJm+dd8TioWI52moiIkEDGV4iSKTKN3oPEwhWgJyPRzR53AjL468rImSW3
LZi6IeK37Ku6cVA7Y+43fNhE0xgbH7StXiy8TC6BDFyFoVxSMjUY+A+/NPKt18oADgXV0CEWBRc9
3xAORE3hxrXtTRQ1jVnSV9dRBxIKDO1VPydeL+tAmssB2aVfZObMZsEhTpBQSnTHsEA9MZvEiAZ8
AwGKSEFn1RwL+E9CJfLzfLz6g9agJQQgb8QY1roQABAcaSPrqGv3K0AR3yqnbxKROZQ/SYXBqZi5
mnoNnmq6SXMpSi591kH7ZiYr84wfuJrusZrlh0mgBBe28X0EeSeaxdwvQXWMX0FzVHNYUs0jIaqy
UQj+BoVq/23QYxJotSBerf0thLO/xLmpRgFNhEa1nUw4H0UZsyxYjzhiQNIbx5yK8ZLMJW0VLYWx
kltmO9CkHR5RNk+CRjGRrGGvrOUFr/S/h97VyoXZlnOlxPdOUQOuFe4LAC5+tjHLMCQtUImsg1VN
duPoBbJaEpWlt1IQObUGYdX1lcnKiUy2uTMu+kRQFLVexs1sio0TZloUJSbCd+CSU+uB3C5J7B2M
ogpBkieFj9pnAX/xKibUtdWRRvLJcrE4GCTifeeGgJHEwiGROAl1ylxnqVA/n6Qd16HddT5ZAt90
FGFjYB3EwIn8bssIMVS4m95pil8q4+Qhpf6C3x59jqGIIM3W1uqISzMddqXWN+EE9uNEAM3gtsXI
N9K82nQfe4k5fiSYkUPH5cUJALxjMu84+V5jG5JQWu5jGI2LbO3zzNjsx9pPVhgz2iDww7dwMaDW
Vyld+eW46pRlU6pKbTPfoCoyY5hO0KuJPXxbh0XY9Z/bJH45OUfFjTnAvx0V6abCBxGtGUIR+OZI
2ThtFaYyMOYwlFqLoCvpRETzKg0ufDqx4UyQXgXUxBFGc1Xp7Q8JPzFDf0ZwE0Qb3fPttnk72mBp
Umz0a1pb0gAUtseEVFJCPZYLbEWKDqaxUUwghghXg4UlNHaOaAdMtKgEKgiDNikfaI8bq4Ahuj3V
ypvP5K+NiNqPR2F+T2S72xC6Hedt2XLxzu3EEwJUnp89J20973x4cMzieDykIwM9te8/++psnbCn
vA1fMBb+SxkqfcPXJXM4pWWc9OgStRkKI//SEs3YkrUgs/GOrT/uI9WP6LdFOma0ChNwToSCz3Mn
EISA3uNoNVfnXmti2aEapDY9oeL8hCDFm41NRsIPFB2/+t6aSCNkgWdh2eHc8P/e5qbJ1o+61LY1
4hEWm/T3mVhj7q3UOmMaxAQ7BUy2FhVLcQ4wVqXpXbULbTq+xZihILrJYaL/+GmTWIsMxs5/uBgH
os/ICxEQsVcmIUP69aOQ17Euh/8MzcRv+VsFsflOwI+J/Z8bhGSc2InsCrAqNh+gHasvi9/K60cX
W3pU1w+71xR7BkYgjAgvdv0Q2YpCQ1oFYuvcvzcCGGjtU6hSofG0wfzp3WxghPbZn5wzA5tC/Asa
/TBuwUTf0rFQE6ubQ2+Gf8N/zEEjTSOH7bIfaPA2zTJRwlUhjwsCbhm8DKgnJFLlsIfbO9McTJV/
1S3sJfdzhXMY0Ey4oBxwcT0SFoYtcJiJQe2F6nKcvdq4LXzfNKBw/3VONAKOsNOgUD0SwbPxJl3/
qQELchpn7Z1rceoHmIbF/k1eQCgzAFQQvVJZKpIQ5QN0NTdxbrrHvB6FSG5XAQlOXHtn6mrtI04i
9hq+TEsdOa7IiwtPyFStBnyqFlMTtjH1J802/M/uaQ0VQjYF07IuL9nQaoe/UAyO0tAdq/rH3hWa
1wDibeElMpaDTbi4ytG7ynCW9jqmtSk64X/Kn+v3yP0CxyI2/xkbmYucNuR1eWReqAiYUZkQDXGo
kN0k3oGrX6qtg9xwes9v8OuzseD2BT/Lqe5qIFiLfW7JG9/D5FKEeQK54jacjUQsWDbpngKJ2udg
jBWTTzwAzau5uqrFWoZkI5yR/4E5wXTcV7Y5EMWUoj99kkJ8Kcaxcn0PXcyK/U/R/Ogeib3ojr+D
WGL6ybc3flKqsf6vMUSE/LxED3yCjvRUxCuk/1h1ZJ7xRvV20rC1DeFJUV0rzwIYCUpxJ3Nog50r
kmL0fQtw/leBSnTujp9ox/WoTL7wQ8RHhdsL+5RNrq2QRE+vbbZCVlf5QWC80B9ejK8Ao8FnwkvZ
6wDAMwVeIyIdGkpgLkLdDcaVltVN21NnxG2ofpNMt6juoms62sTW+JhAhYLfUxAHkxHe2IIDKnq0
NBhtYja10Ht8YpZcw2WbiJLtjKv4zvE47K4TYYywLYD+WPwFIVzAFPV25wXR/zT09x6IBtZmETGq
NC/qZwRnyRMObmMYESOg70e4dxgH850382nxPy2cd9oLeO8Bd/eypORdb1JrMh9vOB1zpTj5JOBe
gaOAx/zNSlCe0f14O0EIQW+0P9AEIwsETQVAoUoOl9WR+mLrtO2VLedGrgOBTkbXxsb6arABoNB4
SGDApHd+Cj5PWCCe0YFHUTQC0BDzrF5ZE9tm2aJVtBELUxt4ndRCtKZwcviJe7lvA56+7lC6RSFC
cMTDhjkEfjIZqlH6JwRSCSIl9onYHPa2N2WxofT7rZ6sBV0l7VCIZ69AvmgN9iW8RyD/L0SY1BAv
x93FOo5Nfn2tiZ3o4w0HCI0oOr6Yg+a/HvHn70xx5Z36t9CUHsuMfAGyPX3s8DnoQHLcHAuAK4L2
yS2EQZO3Qqigvjkg8fGOV6dNQvSMCvXUeNgWv1Gg7cN4CsrXJ9Nl9gRwWyS2HB4lAfQGuHqh60u2
MuCT6rhtVXSpqm+JvilO/Cd0zwLhECoYuUGV8wVwOdr8m4BAlWDtE0FFKNerrja1BAsfW6+Wmfsa
/WrgJX+Oq7n6W45UZeqyVpuPEJNeQIQ0jTeQ/oOS/JquRbYFdHc9V/UKKgFMMoiVLNjDtV2FWx58
JsVn38426VUC9fggROba9VNdO7NkOryS7eFo+1CPiilh3ioAE5N7uuOiOg/Ht8pkE2pAbMVtKMoc
Qud0ZdUXCfHPnTgwWDZhMjJO6UyZNN7fx/WumAEaQpm3PHFpoQlNYpCIilZf189xuKoxt5OlpwgI
ljWMMmQs+ahx4xPvf2aIet2GzhXO8qlKQZt0y+5qe5/ah7T2zVwHylE6xeml50sc9fjynRrArwC0
S1cxc3WzYvIbwEb9E5TKPHeeUyovu40SJl6DCpyU4Djo5o23EqOAUljiALKpiA6zFlW4yYj5G5vr
JoIj+vlZb/XD/qolg4Ux3ld1BcP2RRMpl/SAr6O91Tp7dgLMEK5M6D9jXndaLariH80SL/77Z5vr
1yIwaGMb2QVR0OqtiB2jH7SEovliw5b1uzaxOMwZOsptvgD0tq1itTg8peNxNkOZp4IZDfvDGyzW
A6g+U1sn+Jh3Kwc4vFxIrxV2oLnsipq0ySw7vsP+ag7NacXE5RPxgNlhzJGNfVBtmrRmIlrmrdqi
ldUV3TbwJCJht4fWZQVnB9SVgUZst2WJS2yQvYPf9pW2n83wML90fqOkE3FZBlBVM7jmarInqqTJ
LY1HVFwZALEk0kMXu/rsRu7S56lgaIczzF+hXn4j/bwDxiJ+7jcEhMIVXOwQauWOrndJsMfkELi5
wKsLZgMKOxoLXcHn/J22usLwMJgX1y/2QXJI4WiK9JZNY2Schop6HisnpU/FaCLvaS6hrrXFvH3p
J5b8kgNtaqGTd0Q3bErBDzcFnKXHJAFlcY7+ZpkHZjbIxpKMU8iLjON2OEQEb0PV0k7HGX349clG
/7T5CZuPntxN01rtx/W8gtDe4xSZhwsWkZiCz0jnUxYMItOk3IUTyPktmNikexK8jJ8s+W/ukZQY
K6Yyil7xALWEXV8ISudsxoHPCqdCMENQoBBpPG7V7J+oU2z9vtzMRsl3/9O37NMVkYMTXcNwfKhM
KpD8T6URao/ysZyDRjvZNOTxFM+Y3/KqBwTUoywfD+8x/jadZyVjKIM9wPXRNrvk5fD7yXP3MM8/
4cJW2VMLEZcFhkEzQmTVDh/zDAGK9MS5gAGUU0qQ62JHgKL6pnIz+neUk00n+C/QpkIwOxFzKwsN
Hp7XNAsKsccYFk/ZWDV+OPe+BgSqelBJIBbruAtX+FrfI9KYIfW9k2/wcmKZyux3rTzaGzhtaMcU
tN2MNqOVTcwDPkS8GSN51jhXPCqo67J/f+c+KIqeQjG4qN3HJ16l2rz7v3rFMXETtliv7sB5FTkw
QyX7zOSHybvzFqwqyO5cKAMp+yUBoxbcwH5PVGeiVmzPOXomPVZykZ0u45j5PBVRD9yfHQKEZEO4
ymZGhGO9mKcxEZl4qSk23F88k1He/Ecrg6nWDgORt/At1UaPTWIIjwZNNpBOdrzBvQBCgravp7d8
OTOtvdGGxWLUw1dtGdpWR+aMq3UqKyA0yJzhM2aHx9wHcacj68Rmo6zY3qn/9mY0TQmjd4igClrA
1NaeBS/sbp+x6LF2tBbT69HmQlxuS3PmxXtLx+JmSCrho6hxpoFdhBsMOjJBLgxoOmcGfzPDmjcn
woSLYJFEzOg4c1GAGNxHuJtjMoGNk7D4mIPuy8SVsMs3q3aPKYE9xt9vuJFhc+QlTlxiZyKU/Kpl
nfACzBV27cY2b/RaX6wBPMyqGVyelCN0xzNdrovlaPbvPF+kRXD1S0xFeKk6pvvKvssUkvOgFJ2V
3bxLgBJNW4KilI7TZF5IJW5AbIazmzorivzqw/CIk1na7uErslqFmSH77hLwZ9y2hUzpJUx+JQxk
a/GkICUTqGJrzzTIfzqTHkePssHpDHGX/tbIV2XLLZZ2Blo6CNBFq5chaboF87TrNG4sDp5gFFN+
u742MAdjTRgxBLUvXj0Xq4EYvShfT6kcXq3d9oeNeUFVU6928BfnqUVMaS/vH7ju48WJ69nFLAc4
ALO+M35qPCpmirJk+HZ/pHXbnUonCRvTz2a9+uecePn7JMKfBsWN4x8FwMfJUR/HtQOnWZQ+rNHL
moQGhOuOErKJ2Wy2J8jskOBHuUhZIuz+HMa0bMy8f6vhVl0YSMsGpioNyaQcWuYqj7Phys0PSpo6
+zEP3hNxFmUELe/FUHJPVsAbkGdiG/staPvgUOxGClALuIhr9JYv9GaWf/qWk/ZKG/cHXPx/ck9n
KpRodbQKymmqS0fbCNpYroA5LhsTAZS+r6iVmggaiInVrydxshYHoXb6069vFZ+AdC03zr+DEOAJ
zWHdZbYxENaRCOFD2hKf72QE5H5o9MWymQt0+TK8vswqK4Jexhz5QZ8oNQs8j/w8P2z9XAqBR+tO
D4f5ISXOtDfUnBLo4IVWvcwCvkAgyeZ04KDPgMJ44H96grCZ9xFtX6hz6mp5cM2i1VRt/Zo0FPUF
dGD0d223CZmrNLtGno+FW4JL/U6fo6HiRnlCHR632opuDYEfQI6OH+9/L4jsQL+Ateiy8kU08u+R
2JO8uO9g5o8i1yMJlLHRuQwLTCJDdMVwUoXXRJ8kRSacHDNzbr9QqT5h+aq3lBOrSuHW0RCdNzoo
gaN/hQi29MkEZEmn4XE4lZqWKFrj1oQMwlPiucpwOa/PCdf9yAU0nHuWO+jCQjRgAWVSqImJgt7T
aQBNV6n1m0jPZD9h2hYpb2TMt0bTxY8T6ftxZNkULksnHhj3okCIx7o+uJA6Hsfse8X45+QXHLZ+
3uhSZ3NowEXpwjhzH+2ysC8bUrfMZCn+Pnn8dPDPW5I1YJ6qFkeqJ0VKRh6Di9I3Mrvwc49hHQLu
1qMuywfvq7QabQG+pMpVamqUMQBl+38Cpa81Z1tDXtWXrbWgUUgxKjO6wuMqqB4dvELmbJ2fvBIY
NWnbzqq6ZwZT3CgSdnALArWUvoV+jPftFOtUnkOEHHWrRUM2oDomEnz0D59l2hqiuDNEvntKCWoU
u1/DUMXbNO384v7dmKXz0r4/mZumY6QbqY86+stdVUyFiIuX2L+XZsXm97h877bHWVgbX7SOKeF/
dKFxOEC148PxkZvx+Iu7RJGnkup/6RdBfOXHf4mtHWMH0GjvbuylH4Xy5asungaC7IBaGxHVLoZ9
CHdXSIS2LJJ0K8PEgEV6iUUlmYw+T4j8lTjJAQvkjfSRwkRTnB9B9HckGoFsNPu5v5axIt/Nop3P
yOsCQq7lytG8e/JLS8D+21FADg82J7A9Mi/dlDtz3T+xbzKManbmMgL2vkf9hsqole6WDYpGzcnb
Vv0pVj78HLhTVTBDH8Ls3Cp57SBr3WBtNRx8vpCHgjpFXaQPl1aB1WsrzV9sVCmX6aROpcMqKh92
nKaBZj/wHV1hudFXfut1/zgztqCLNIjtSRPGAROnlM5ODXZkV44oTGPXdza+OnjCuwn4E2Y/fww+
JSNErJTOGp6YU3nQp+gklJFM5ZdeEJ6L7uMeqaGRbg3HRPeBV8+lIVlsmNdxy3xrfPpcDclj4ssN
VST0+omZnD4QINEoWtk0N5w3G3aFPC6J8YfZycXSHLovxchjKiTaPrl6LxWyyta+GYi2YwA+crT9
Zb5aHgrS8OxAV3YcQYwqAGjTC8xsV5uPA1EAz9GUlXqvirWBwblJUxEHW6w/V8GTYHHoeVkCLOfs
fOEGF7WXw5C/SPMvTH8WPKpTpyvfdpDWYi9GQ6/1m6VgjYtSnpTJvgFbEfAmXRB4aEUL31bUWZvL
mCj6Y32T31zyA/cF9/MYefsguYd0ivQSuNaxwJwBq5iOfXRwp5HEVz5IcbvgtOd+a3ZMnXzZDUB8
KRyks24twsUAlqdsK9WCGpZhs03+wbnq5bnlPgFR0W4Liz749ytdP0gSlsqMAce++1ZJEBUQ+2BS
DRq2IpqtISBQCPLFcnqYRhEQwixtthUnkarYhwLHtvCWlbpWay2fXgspBVtETGEnArWEDq52biI3
keGJ1Hf1e2e8zp6jLpRg75ucXMlfi0OBW/506iE52iutrQzPHSG6a1iJoq6i/IYVCuuM95bkik+6
l3fivcJk6gng9SmKvlb5qeKkH79R+cW7RrfCGn895tezRYzqfUjXSFbBIw04mclbDifieV1+3YDv
9WgTJmqkLuMH1dMDRe/Vmp9NqisfXqvAQ48Gw+zB7+/E3wdGC6RrsqdUKUUw+jR56yonsXEGzrj4
T6ArFulo9F96T4UtNQmTU1rKlF21cvzEhS5tPisPIqwmNr8DfUZWoAs1u6J9eEqlE8jKb2aEdOuC
x1AKUzGbole40lvJ1nncDcg8W+8VL3j27OLMI4yw0cOri5EEfSBkN9mJiRPzX/0Ys7T1M/D8ISJT
ZrN5nBgCJKxw9U7OHA+/gdnhjLneex5h+bUZtUfTnVkgMz4tNYtLlAnkvklvCt0JAv7Miu0v7Py4
9WlEF/vHcFcMOAaUCWV5zfnE4TggShLDgM+nTt5Tw84nt9NDTJ6eO2LAUS5+82zczuyjUxKSMmrW
VFfyzPPuMgGAb5GaXgEib+87H32udh6QcDLWXNl6yB4IZQdJdz1mxxQXVaIjRfO6SLjOhXKG+IVf
1FNzfDqr5Ges/MbWR7WhAOmuThyZS2M/s3BhnizE4+O+1wk5LTz/tt0KmPKGbUEsJ9wIwnRWo6Zw
+mzBQyr8TpJEn9v/FiKIJErhErapklffXTlKYaswYijXLsHbgbVy0RnrjAdLAOcg9PkJRsCvba5O
a8OfRfl6cuwC3VGci69ayjUDVZA6nsBXTDbUK0iFk4VvEVLgy7kIyUw/siCRQ22PpyomEQFJqSmQ
D2fG9I6EPXbuoA3HzaODB6NnREG8tevJwkIaIIZITNzOv1/LJeb1ev1UuwKKEbzA5/8T27cZkuZ8
CawJI88pRJz8SPP3pM+mFFd2zHqeTrnzkyRFfmitE+U+g1C3u9DLX3i5pod5cBRkJmJXRFUnZLtT
hAJI3Cupva4JeGxV3b8oLyLSXttrSbw2NA9O9+zHFK4CBaEYjeQcOVcQTb9qszKhXNyC9QB1dT+L
HqCJk9rBYhiUUimhGY/+KURW2pwG36KtcsYp3JPtiR3zCcwnGmzq+0ergqPtuNrEW8eFzxkqBkGr
6+QN7n+fhjHc4jNJqaBaRX2bDAYqCBiw28d+6+LSiOESLd+5KrU8oNHN0gssqMU95lTJf/Vw5jm1
Je046yL8t2I0V007pK/KBa3hrA1qjxbsnW6nnxFFANb3iMyxKcay+9mHLjPfbM0jydt3/YP70fEo
DeQWB4J6w0s7yc7AIxNaOabVY7N5ztHTEXmoNisXZeTkPuVcyU5rmr4z5Du6meD+BeqxFNTvV+mG
JzYbwV3B1yDJTRrgHKyQSZJn53Y3uxhy1ZOouKY0VKMXHPZMJulzhsnvMyF5vG+mF7/0q/RjhIlO
4Qu5LlJsy4LZiIxr7wu6rEfXHK+g0i6VbifIKcyBSG3vxhN3ml+3UGnzjl2iLntvdvr7LEftEIev
N8W+7ivOtw5KAfjVVkj3YvVOebjwB6XFJhKe//O7PrmOOLTnGPvXYCwcBQ5FWfHrFaSsEwJvrz7k
ZNj37tBlPrxXooLQoEzJ7zqkRppc4RofoAlilUWcg5+y0Avy7NexrOJ6/WFDPY+IeI5LQWXadh3u
KIR1Lo93vC1XklFegj2Pvun9SCzJaQRpB/IfqPTYAjGe9HQPyHZK3dIPhPxMs+dV1bgru2RlCqLo
CvPe5d+E7xdnMP9A5HlXV0KdjMbQQvmjP9PJJLRs4AV/PtHbHQnvX4hSWc9nahBlBtaLDZylgOeT
/YhJcNghvpU4A+PS+u7OOq672Sm2WaUyIlvgN4qO7D13+up3YFvRHZI/n6I6ZKEPvrtM4E5McUcm
vBZRaZQixNCf0e90sD8xKCXEoe1jjRf0gtEdn3pu060PrtB9Ju07jb8TLjc63M3H7U7KBLFir6U7
NprPQPNVzr862u10WMtYeUw24jE082JZzvkex//xDp/EV4xQOBXyM+EoiUvW6pq6lLh/RDaSrX64
q/Bf/HYIy16+W07Di5CpqAVsC5IfCQA7DlymCVE5iDZLj0pYO59TlOL+/rIRvNKtW5cRJ9sJEL2I
4HBOuJI7bmmYH/PDprgXk98kXYvp4nYjh++3pJCsA+ihyu/f/u1zffn1faq3l6mTTkXHa3MvCtw5
K66XfCCFnYoWSo6TVaL3nsP1UoUPoWuWYPq1ISQJNNpjEq6Cb5LmPbmR8xq98qWUef9deJEAlxm4
vp0pHUXyFd8+D6+P+0AjNI3AZ1i6Hy61GdazrsZu6ImMFMkZXpiPPAEqeEtGuKQWJcljWHf5YCA4
Gcw+vTTjaiV7cNltHowoIYdRRrOLKGtl+tCl808sgYSfm+eftvlbDBaxYoeUQkcxhcOglCQTyIAw
SSKzs7QsxExmGH2BIGSdJ0KUMCEu4+hlF8YVW/hTV6x4kcyrhjHHSaQV1mGt3iIvs9lXl8LukSeR
K5opSEBNCKUKeePGSm3vV0ytur5+R3fobdV2dtzb55OX4mlcZP2YtKEi8ztnpXTQ9ZK2Sy9celK/
E5fZK+Z0TnQmK2CXw1ODqis2CVe6vQidvElPYqFwpKXkEyWPneEj1H4rh/IvrRN4CkpbYTuEDk1B
jNxOjUFgR3l8Ep8z0qQcJNVq4lyuhQNi3JL5zGWQvqyYwpOGnYXaUz8Oz04EmjCJjQqySvR9wfAM
6l2Mk1ZwLsc94L8BLuZb+Maie2rvZovfARsgMD2zvW6zpcFC3nd5M9vcltQSMyjRbUobZg7Q3c1G
Uu6n/dual+9GDjiN9LAEioxOle1IvMxJi9is7SDMt+LvkzzsFsg5ZEVmfg80lhbDvoNQdl/U8SHZ
q9uxqb98U74YN80mroHuVPOc77BDW3KqnO5JBeUsf4cdxVc1cLgvDm7xuWLQb7d0hLGcCzYcHpDk
NDbQKUknOvXP6ZrGkQjaudctDP2KU15lxlC9AWQtlkog9NeOcFf9B/+KrpzJCryuZOanjJTsfMFa
eNb8eWz481mDxnF8iYvQJjUzYa+HVdALfpDXp/LTP02Li1+pnM/VU4pt8a4UeCvAQ3xTbWsJEtQn
1wMeA7X2CVY1pTw13lZFEBwjJOYXQ1773/6O1cHRKv7Qb5tFyXHu0ntEPIJBwWGMeAtqBWq4JcAD
sLKEphljTF1J8rT1+sfZiy2q3e0NsVPMeLHkQpcqREVmQKetmN/SoZnIrtmpaC363cZWzmQjIROa
qHpyukVogu9yCIwaXtjRBKEGsv/kXl/aRoJrtDGVj3Qn3zT33VyFoY+N0VpnGzEAop8Y0nUTLisl
4LAboXVvRvVJJtRvPvgKqC9lANyvYeNPLTIU5MTMfxUmPtoltCwnWUU+YkikvVFIM7fpdBbNqpc4
sGjwYDe2os9/2v1PrgjP/xyKtF3rVNJPQ3tW0EBwzziXZFkE5LItS/m+/AwdXUxCd46PnnB1klEb
neqfPwdZudCP8oNVajg0CvNd6KnyBDLWb3qBjMw6A/Sl1mmZUg3LPIFW2O9E0IniB09wxDvyDcxX
psRxS7a0Qw2QC9yUroLuvOkwmIgnQ7ld3WAAPk1MvJh115txjhmPyN3WhCXDWxCrRduEHqS0WvIH
gwbyrRCYGRhuEutZ8w78lwf1ZjGoyxED/iWbxb1mpTZ30lhvNcrrYOpXjtq3aWAHh20fyZyVvTGn
oPkAh2vp0ZedeyMf3evpvUAhixLkoszF61N/5md3Xp4ZLcMumgknzj9f+Rg7I9ukJ/30NDn6NG1v
ITltv5lDeOCpK1HJAWfw7w1K3XVQzEwksyaaxOQ41Kdp/pm2tXGS1Ndbme10cT2e1cK7W1I5u/1b
yzk9VQSVE2SYCf0l0s0P3iauBxqWdFYftna9xtuMNLQ+ZD1Gag6eQ1/LmYQ5wVzUYhLDIo5pglWl
nf0Ej7WKWvp+NVrSBEJx+RG0A+qVPVh4fIQuHCO7zJ4X1VHrrUrgcGvhyt4G4FjuiBaCzUB88k6J
ghFbwS1ze2fWNgcCdaSvXByn6SgpHiE/nfjvaU6pLJze1urb+Dbltt4Nwt8bhfRxWtogmjd64NOc
yKHfr5079WWnLvknWmtkXXFEEwuGGySrKnA0KOq96sRy0uMFnXuGrnZNEs4ZtqRNitOHTl7ivcuA
FG7NP6Beth+Cl1lhrNhknUQQB3WT9MCQoUhuG5GfK2p2PMv0AMh0SqRm5tCBZTkKdvkIcneq86ZZ
p9vqsg/mkvXnDR38J+mrfltTiIU9HoOz7/3uQY8PiHsni+ugGaD+ra0eo6TvN0M+JjeVrGtVmJ3H
s0D5QuNQOf1N2l5EQQM8uQ10u8m6D7KCWhypur9e7QDiHT+DRGDEv7Tpx3wO8Z/WswFIACPFMx/K
oPWrxhx3p3JAEXpAV5MUP6JWwkn3efzCvZAN21AN9nH6IDXhJO4w2902P6jGkZPUSl83PnIG/Vmp
RyxEzKVPz1yEaZOXskIgMp12q1uZO7q8jQFtGotWs8ExlVIeEsbNLbC1L9o2Cn3TK6PivMh7eRPI
f4pXv/6QwxPtwt4gf7cbQRrQzwx42tk9dCk6PKjVa3bizpHujG7/vpOezJMszoPgji+w5q1ROEfX
i+CWQQOAYQcBf8VVFTiSPgKlmu11MR1Xm6bqNgASz69WEzUlyS3GOqdDoRQliAS4bTH+Qj06PPTu
oUTR4+JqivNbOgMgHlDwl2hs0PTlMOKTMvCjFp6a4+JV8nNldrB/d6xmc9TJejmbWnuKJrQbOqat
cblR4GuqkQ6QGYuGlCn3MymEBRkzHDxRcSuknU3nT/gvUfrPIXN+WJg+tZETulfASY6QlrKcvsgD
uIIE5GDerhmfc0zPIzUTA7SptYmWkUwCoKGUyGecJeC+a4xMHt+e4UACnZvtRHVqJftQSY0qlrBk
SLQjL9OLBEeeWEhRW3CyU1g5Hp/biEsjlBz0rTUw6bLMvd6N88iA+hcdLqxju/GLaQPyBN+tm9GX
qDyCmahvY+iILAj6x2Lc4uMP8/YLWc0rU/zozHw1Nf9YOX+eopyKJbnz37uvICIscD/5CRyqM3fm
gIE5AzVABcgdz5D7XVD5b1q0S3mOT2odO9/XqHD/2sMVtMDF23rtCPPBUx7O7Sg7mpQA/e8U6Qmc
r4BG3jWimvimHXy0/spspdySrUHVqDgpQnYupSaJj/072PGJv8jlYOQCwuaaY24XE5cG2xFD27CO
KBzFa+hSplixFxsV5w33HxVueTiB7y59ypI0w0pwxyG1BbmkrNWqrcJDOcSyI52QuseKeUUna0e4
qK78f1rAhDZsb+LCCGVVq7R+OjLOERnjefCzXGOrG+wRjcFhEW7NP8aBW8ANLonxiC38oC541GsZ
DqMQOMwmi/I4xVum29A55BbCZbrtImRJbYKopIINtwwLq87LcF7WjzgEE7DcpuhFs5yq5x0zftYa
FcXCcGLwp7NOShEYhYkiQhBz+xWBtUTBX6eUn+UNnCp6kjvemeJYbjQMuwct2/HsN5p5dYB7teGW
4g47Zo12UZtsPPWrmplUdZFuAIMvHKHjWj2DZJvkVBIQ1UvZ254bTlhPnU7Fr2gost0+eSa8+IiV
szp2BeIVn+okK1S4BznW/8wuX/EqaijDw9fsnadFhqic0NkyDhERf/ecDF1vgpO8v0mvKCKTtJXN
czOTy0LZ3pWBikB8lxlloPQFfOlT0jXIzd77UrfjCxxY9qgs6LQKwtvocEfUyGeyQt6HyjPfyZiJ
w1VOJSQhRerRI/MlAjTlH+NxkEDe2pDVHw+gJMBvYU4Ka8EeJ8ngKc/tuh9stE9KGbvZTAjmSD96
AZnkS8RvNg1PqSiRX+VCxvgXLVPEHvhUqklXYPYEr24NthrFdvDkwcVog/VnWZ+70mHpG0t2B/jR
0En9Uc08XEUGNF28vLaj5l0UjDdUVNqJMr0RiQlpU/oV7XloFcbW8TVg8+bDUbQ+J6jnarhQbCVx
1cf7racXukrnIcSS4/s5PYIxmzgdRhB9REvt6rIwdxacQRiY6IZIGA3KGxjBVnHNZC93Fc+e7NGZ
kRqaRYysbhh6nmKj3UHv+zSScFefwE4/hrpOb6OW7FbAr6RbzxshsTHfvhSv2TLbRK/CATNzglTi
PGieXrddwm5lvRxhU3aqOZpmqJasZQ+L7xzdxYc0KGoppoKQOFt+zWcokBVE8WlLWxM9OXWpb6Eo
dSW11/sKyMAdcuZvQNf7/qmBaOM7EBwiui6oROTiGrSOP9aVZW9CVxDNyQS1bn7R+VV+gzzobF0x
jZZ/zxwRVh7zqPtVDN5LNB4/kZGX3atxAcE6JhveNqk0pnlZ5rQkuNLvvGkzV+ECrb9QoCnlSIXU
ujECeIAcfr15FDEPyMhkHyOUhQ4sbVVNNObs+Kpbj+5jocSzjkiJ4oqGzrx3dqpul2Idqq4w+YuL
nbL6R5nOb9e472at/2gdKCwzgxlypiN7GOTVTTOUSZKszI0Pkm6S//akV/bRpGn4s/EJpMpkgNtV
VsvoxgPE2WV58VomDxpRCPHp5xqHLKV5PzbLKbPwtI16hVeaj3E3HwLOsUxyeLdKtCNHpEKASoKD
D9Qj91uJkteEvWqIsBs9UwmdWjVdmVmaeWDjM4PtYi9jWcq5ifXB+ZE1hEDeiT5WiUGClnZqx8T6
4dUM86E2qWMHFy9UCt1LGtANffRMr+GPdkH2tURL3yCm3QJGtJwWuM/7dQ7RmeT0GFl2bM8vYYjY
MfERjvLuXLfsSQRC7J8c0z7t9KlwbK7G+woEMdARORh4Fo0d8nY6qvCxOsghlbEhPIQQ/GTjTLsa
ZAe225wUU2K/GLZRpxPG1Za60BDCtF5bwkskEHZvgcpk8VzAwncf8l0LMiTfZVAJqqFDlZFTIKQL
89hI9JBTbdFkhQCU1L5MMZHVlhnIrqhjYU6xBl2ZWZYGg8JUgLlqbPFW+vaOCsjJyV+0g6vWg9JK
COqOstFhFoLqP2T4iV41X/Gu8h5+IIUBDoxBSXSvLoXICCZPRdQSiygRnAXSSfvq6Okx/CzaiVB2
4In2VAC5s7HGEJKbYrb69rvr5VER7O1I/qPlqv+p5gvNrnWnUBc57VjKbyfyqUtvMZQJ+dMfJxkS
HWhwuHtIcNT+pEfJ1hBFacLiFmKzzWZXl5Ompc9MBBR82TNY7eK+0FlWXno8oe68xAXBRRUF7rU1
FLRHuahrDUX75/FHi3Up083E4ktlXhzEpVHJLo2SRQ1ziUBrObPeHDFgLbbaliZ+8Pry7MHeD1nB
h2X7kCkyFP2/A7U/dEan9xe1fZhJAb/TOr3i7qdRED/f2oMHldD6BG+ruAdMFweFABeZf8HREp5b
Cat21T3V+H5PuMASfq9Iz0NX13f0/6QlY1DTBzQ5Jl7P95+Hz4AefWtcJ8rouDildrUG+lhzNAgg
ZMprAZdjD4lRgfLvl6E1ah/cKbQTb3MVNaw4jUPPmbgpf6vDUU11wkvaLQZXQRMVEvnW9B2BBjFV
Dt/FugQAmMdlXp842//vFkTaxuvKSHf3ecUFjaaSAZdBumbzrazOKLDb1hT8lIHVdLnB99wsgP/Y
ZhrHDRCVcP4slfStlGHeMBzxxNG8YoPejiwhkDYZbBRt+iTJsMQXuu0uqLNkTQWyMEPlhzqqY+XM
N61TEDmY3T4C9mEqlQVden3Qp0GzIBkx/OiAxsF2CWIj0ta2NwhTsmUJMYYTHGynIIkwn3CElACs
mfxOAN8rtY9M3t99bpFQYPf95Y/Fz0Sm38If57cRGVZ0mcUVRRICar3vMR7aOauD8BOvR7wCOwa/
ogHZVdHx8CKhgDkphCOJVBNtcFcPbQGlk4Hj6JUSFmHUXK/yd4WiNxpWx92MpdL6Sld4/J72+N+u
Un8mtbD5t4XrvNGNopCKGAhIuz6C0Z/t1geuwVEodF9qUA38xegk5Fcu0WaRspzO053ETazHgw/F
m+QhS0mPm3oMKk3CCn7FycrPFSvFKWBGofHD5KtvDsOM21na5jvf3zx6dd1PNAgIEAOiQJmcLedv
7eER4iLM45cHkf7br4DpJKZyZpw35JcPH/NzRyynA9YD+n48q6YnmDG5TWmbBNUSCLkC4bT552x9
sKhRRc3devRM6uQdn8mB2K8DlUsLA9MR8CkyeBc+GOH9p2JiThCYcbRiiVRQLncAENQu4Zn2JdJ6
yQpMps/OBCNQ1TtrdlYG6O/FDzgjKjRBuAmvNZ1MnabuOloElkFR6RrzYOCXkonAXK56PV75/Ll1
saezkJ+7TZzZibSsxBNq8p7DE0uqlgQo4J7a1e5s3RW1ofpHW0aUno0JqRYhlE+/b2idAuDpGSFr
RZ7OzeNKWeFSsDl+fs7nZaoYfhzUt3sbQ9NzD3KiquNN0BAvY2nUNE1G1rB5JWiddVUXwPLMSiAf
Z73k+jnwvztdAfg8FaMjG1yRMcfn0IP0ro4SsJTCcmSCsnS62d/wW6MQIf5kgqOA933dFXaMKNhA
wF1RWr7AiQebYpDHQhNb3/jxEgYD8eN+z+esMdq/IZkSdgZgyoQwZjEsWOwnSokJVEIubTyTjTg2
57CkS8nd3SxkIiSf4WaHCkdnlu5K5c4DQZK94bEtSWNW/0duzYin9WXY24VUR8Rfahh75oaBokvz
2t2i8so5hJc81CG/fJiPLKqLoX5WN75KRWV5yNdYLTq4NPWTPGjW0psdTUgHN8l2/nw/mH9fxy7M
6llXKex01KlsulFbNZx4GX/xe5a9CZ8UlsLSLeg2DgxP1IC/tBT2TBi4ftTC6YJfKcG72tXRHLme
eYKqEw7gOmJRXHCVxQ63ha9AnGeyrBoW1thKjU+bWloUoP8jLx0Qnmda260h4akcZ4ifV2iq7E9g
siRZSwy66x9y3rB8LgwuRqiBPJ7xf4ueajTL+MywBIofmKBt0Xc+yzlkZGbG5J0LDIz0qNMq5gA9
wORDlzfJY20//lBOXUX45dPrB11bPFJHlPMh0MNvicR5ITNfVVy+wGJi0FZnRTIAo5327kB8h/RV
a6I/d81zmzLScNn89Epf1hVkJadzAW+LdDCoXFZ+O4a5ADdxlpN8CUAfu5plJa3yqNgx1lgyPsQl
d749C6eysBjMOQdAk2ZsA+RFLVsTAPWRYarrWwSOrRuoaZaZBP8Ct7Z+iX30ehA53h/GpROYXYSh
m49OOFLLLXsiOgXRqwRqGmxJmqukjsvHLPNhluQrYDZUibGFdrxMPs+sTrKzwx/nFlG6rfQre+PF
yGhqbpjcc/Fa4jHCYjDOFSvCjMkmtfwkMdpTTa3ZWqKIJYNUkdoKMU0RBHYgnl5TlxtmE10lDULJ
t9tjeV5Jl3Lm9qqWd6bUJfe3zo041onlFo9NbHtAF4ZMgygxJsnpFEBGvNGCg1sPE2hROxhkThhU
iFkyovoXv2OrfPTbQF3Fjfvyc5eteOv4Ssm2MA68GyLH1qpEErr1dEU9PGLzDl3+sd/S06FRMxve
/8hpBljUadeGnrjqsGxzU70ELyVKOFFF/lDtIRBVf38TYZioedX5z3O7jyMofSQmE8OnnQaVC3+K
Ha3QBXrbN9RtlPBNxjpMUyso6chLKa/ZYGQ/Pp1b6V32tiadNY60VjRwyI7BRTdEjuZupkMKMjTZ
E9j7rNiXBm7pnJ7WXd/yTxpEY16azgEBukK6q74XuYSU1K+2UIb7Jr8m9e+PF9fnICUSMQc6nJ0W
wBD8k7EqZvAKXeQ370Bt1eeYwuf92nCi8uyJQA60JMgBqhKV9r4t3WPTNFrUMHo+vZH+PJBC6rn3
+sffJ7zgVBL7NSE29vGweMVmVJYrZuOXYegt1kdDu/yM5evo03atuvSHbyiIfAvBBHa+e04nKtEH
4EufCp+GuKnUSnAmEyWdvM63Ae7SYCYAY2JwqXrcfRBgXyT2C8gLNz1zV5uFQ5WvJluzVDpxipIQ
z/StmyUmn8eFpAoJuxrtM2dxUvB2ut83fcrAvhhJa6v9jn9EdWPUAOOqyIWnRNySYk2+p/1G4ctc
0q+Tq40V2gdWL57lYGCDvNig5r141d2z9/81gMXlsR9NxvY8lEMW6BSect/dR14n9R36ZShl/A2Z
wbChitNeGhXp9ol3JPcyPvIrwD8Vr11z4iqN868ihOUazX+XngW4E3NmrTZYGnYdvhI7lSXdzayf
PrYjalYytVMRKwFA/3hPvSgETg6mRSCEPodp3g6idoXue76jQqqF8mgDhYGcO8mr/KcXmyN985tf
0xpd/1M+fzjehPa+/oBCRd+IvM834LdqCK+aIUmnkxF7RALxFynpvmxk65XjD+IMIDBjarw3bHD4
lbZalVkEhiWuagDjncxaMjWdlIrQRL2h0r5OU0XsXsxoG8zohtsiJWJNkUJDW96To5X1xOfUzwVw
HSDggItuCzr3pnrtUSKLCxnWRiADS5pjDb3HayihNPqH4800FmmczJR+6fMKXT2v9xLlQn/4i1ci
Ot6/ca9k+s1kDYE1CPKhWpyb2uR1KNVC2DRUBbSQGa0Iob3DQFVEZZE3+Edrq7KF8EmkIHfSAF3z
49PlSs2c1cNPlYhUk8v6uJwVC5U2iXCOrAh2pAz3UbAPB0Vg4Xl7eGaztKYWqeqwgdlHWDhmQPN1
dzIEkanTB8V+qKhpy1Qv3xW0apGt3Y97pmiQ7DI5pLL/kOxe713fwXg3kocfv9l/bykLyIn7XkRZ
ZWkmngcRFd/zLcXLsSN8T7luw8G5E689pHcpJsl2IYB16YlQxBOny9EryUTcqRZqq6JqNGM3F/0o
7gNvLqwea5AyHAEZIJPNihRVFJOH5c3NRiuEzIuMKHfBHTwSl5Cw8FiYPCekoLUPqQonxierJlMR
QcEkWZPs2GjEUMaIpjFId06X2f7E33pSzwdYh3z/zznkNLeWwBWmLg9LSDr6ttCJ5oqpzg5BUDcK
F9JLgFcNDaKaCe1kcG3SwzMwXurV8c/mi4a4u44tMbbHVZv4M29LYwvLJ6uDTLNFXcfxbEHZOOJS
QIXo06CWSq8/acirceJZVYZkNMGEFqCKh0jD4k3oucDoKUf6qDJTtdwS+QYmiP946NK4iy3E0wxZ
gMScQWFJUEnNILFhjbOjO9PkNrzP7Wqk2MWcohZ+U1nYKqwBL82GzUkZa2sn4JeW5rMR9v0NEx+v
WqHXnwvf6H27NT9/VUst2lRUFT6x6rvw7UUSFnuqj3fdvCPMVfOOMymk2BU6BxtdWO8y0NNgwQuV
CzB1RL4N1vHJP1KSuXipbtsgeU/iHeMwmn2VvZ4EjYJovNn1FGscpAVd3PJd/9mAj7r5pXShoB8x
eoUl4t7yszn+Oa5KDOh/x+2DGNLbDrLcxYNiewD8u/NMFV1Z3CWiM+ES69QfkmhCKX1HfmZJbfeC
rEalEgWWyu2oHR5uZPMArC23ExCfVEnA52ZMjcXz4oslJMdTRawg4UhfeHd2HMaMI1BXLaUkdfZW
UsqsX7HPUdanoBdtCGmRS/BNvTz6o225DeE0eU6nAyD2S9euJ2R7MuywaEThSYwa/OrdvOAaotHY
cJwuiwxErZOmuaiGV+ACD2lNOaXrfE7wYMvSeV7h1ZkXkVqeC4pgdu7x9WYSYzZvoB0W0LhMDh3S
QwbQH0W5sxTFmKF1m1L8saFim1fcRajWdCQ9sgYbDg3FgEj+0yhLb2ZR52sbPqZaNxga0/AZgqUw
zccWibzxmTjKiq950vyFojp9W1gOKUVJniAL0BbHD7hMqmw1UTULPEtzznq81MxXL7Fv50dZPa6L
bYC22enuJRhAM8pO9RKF7ytQcdv5hMUNMua1oqO2VwScxGk6jC4bLiAkInKmuC/QVZAsTVu5+un0
ct5R6k8Hkk1Mu9woy+I7373Lg3SkBzBZTWle1vnFvFvWfmp9sBdVnyBbNG1GumWzZ0QxYLIztJs7
JT8Lg+Bg8QJbWIzQw9st8fWa+oRCeYf19ypga/yLy7RqL3qzBK7p9BXddhDWoEBI+/Hfs5ebByLm
+HNuRYMvi951qdPRNqVxuprVeJhWQLIEGT8ZbaVSRsFbpNLxF65/oSGjx5WJcNOzRoGw/iKeg5iU
IUWCg8QTCKFQX/pbqin6dAhbjTJzn03OzeOMx5cuDGdL7mKPojdD//Oyc2af1AVOnMHPaornEY6H
H0b/EgO4T+u1jxlsW4dwD83d0Xwb2p30Vtlbp1EswcCdPPDRMxUrmWLJPlTMW6QXXBHBquMznMH1
tT0y+HLOHPM16MmnaozIFvqPhOzBZXXZ3fI9qZJRBIUb/SHdO4ZDvcvB7+VQlQZX5DbHBc65thAt
PQ1GWtfecPI+UJNQHbBbHeGtMQEUoBzd2V5cSFcCv7ITgoTVaoYAukQj81+J78R/6piwdKR8I9vJ
cBbD2ah1IBGL31pH1ogJorhSQGS2onhJ4QSrztQQLSQjZ0u/aKTrzz9x8AF9SKhlUpa5LAjbr6PZ
mJz8x+fyLUtOCrfjdFjNcavexTv/Rhv9ArKrIosykZRkYAANOYMszQTmInBKwcrBaJrT6a7aV5lt
npTAhMXuAczX+VoKipUQ3vGVH4fSY7Zuso2AKxCisdb+Y6Q1BZqhi3otk8VSZyYAJ4P8uKjAbofI
11o6cmLpS+3NEzYBtygXcQ0Kge1yj0YELTNAYjMhD3YIh3BCPkI0f88EEnBXm8/vfx14cARe9ejL
5koS/zvu3aZlEUhfy2aWDEo4Eh47FpDACsz8MbzCKb5wpYlHV5P19t3kxzjUBjat2PAaXbUAPeDi
SIhpH09L8VVM3MF9854O/n3NbkNeIgQ9qsYEbTjocfvR8NhLpbEClwHO783vGWhN1Kq8da1APkxP
6aB9O8Lg7x0AwoFvhvZ1K1YyP7TjsofsulhYInZv2hsnHY2s6GDloBEwxiqJX3RY3QOMgeFOy3Ka
kSdtkLt8BRxpTY7XtoF3qGeyox+x7csTRNrYemt722blw4CR23dGvAaAtkEHv9klq6NieFN7wfSo
b/a722fPSEjnInoYoc5r3tIUhc0h8zqlAy8vE3aNpz2GRXcdZOp0JRWTdL278tfJD7IzcTjbbVpZ
aa/LQiKV21zKwP1C3rWVZs++VXLBdK92EDfT6L58vAHSqtmfV7iabwFp/ktX/A0Rc5zHTeleVTE9
LGWr1GLDJRSBqpn1XyL8aj3q2dLVkIE1uNj0+lipCH9b4A78bHU2NTsSAjAozS1Xi37fGGZT0uPA
lx9CyPzYYbPNHaUdyzLqkfO01Q3rnE/VjYF7XpUNdn7nj5o31DuXpixfR/eVZUI2LuYNDkgWENNT
Wn3xjIlszDVX82ADdPHPsEb7sWW093Qaz5/uOyik8GGs1yheL4qdmOVBiElrWTbfzXFk27rY9F87
TKembg1JVJO7KnAcGycl4V6jr4NADIdsekcR5G0cZglj6QAu3ATLHYZLPW8COuSZtnb/0AJ2cXho
BJ9bPlJ9p908T98q/iZ1fzMV8xbCnFesor1Ii+wW4B/KuvAUoICm9wLKQiH43T0I3aMCd3Ow/HVB
lBy5kLJvQCTtBPzxVAPZAPL4qhW9QIPZC8BfISaQ24nRULff2yI7amRpsDYWdnqFMFgpNqRQzmho
UNNxEYcziCrv59hWsgYzGIgy5qBpBCYjfIfhMPiwv5JoBjXS/IYnyGdxi3J6tUkNizeCqQeg/TJg
qLi/tOg3JZ4iiuKG3R1Fc+SIzz7HS/Ltex3qwmS5PbJzraV4baAk9c+7itGE50xKLzKepkkAAQUd
zT19Gclt467GpJlyu6TqrgtMDURoagU/WLupieAorkBNtILd5ROYxOR2/LwTO8rm5s7kRQcUvZah
j6ayqVQgv1ZGv7s2HXTEMWgj/FJKDhBlfOqLiPTaIyOhc7RxWhDnNxTHj7h5pxLwSVD/JEbuHGwM
1xTib7dxWXPu0W+PqAH7ulQwb21QAAvze6pgJ1iNZ3+YeUlOcfDBbFt3pG0op+pUTvrAUUaKjSfD
E9mmhP0Z4rUnwnOuSWl6dfSXoVW6m7smTmaLjSrmuB+JZy/yL4wR0jJxPeYV1UaIphbyjQT0gt7K
75VFbAsLNjnXZgbIAyTFPIDYdtOKeaf0tl+um46WxSF/kDCYKEPzyLRMcuHXVHCUZTOsj+t+JEMN
YRQJC945lYv+5yjZuoyuuu3CqHcOpJCgaYZeV7Neszld/nNV1BMQXVW1bEbNDen1AII+jAylPtpV
XDc3o6g+G9Xi3DLgZirnX8PLC/1L92U70s9QXU3iSLJ28VSy1Wra3iv/IU77lftW48L7429KqyUs
ojpKjP/ZTLECrv3jIq2UDvfCNA4dmM8yBZdyvokhrnfxgfU5c1CkrG0WTT9V+LbIjk91CVv7jKx1
k2JeurFRzsM0qOnVMYdtoLRO4D7iewJdU7sgZak9Err1Nqft4t79mpxtt2uxYFlpIvCmW+YDsM9w
ZejqZOchAq9QC7rmCpbbnEyYtXTbYxlqEzm3wcpS/hbj8/tnbEaYAzMRWebvYX+BToMFwF9cymxe
+Qnju7+6OAO9CZCTAtMQttyJEwU8KqKnsy29JnWIIwwbPiSuewDuJCQ9fI0R9OM5xTnTiZR+DsEL
+c2xDQpUu0OCKIwKEpiebywDsFUrln9yTVFx756IrrjzOCPgf8ZoNRU3LD2E1vWwZT8LEKsdOAQD
MU87DhbQSF/6Rj/mcdVnOnPdXKpi6hAjpyPA/Kh4VFAc6zzcLr1N0vKG7GuhlEeUEAZTNcbIPEDl
TlMTxMN1u91jiT2+UBzFY6HKboTXweUiKzZsEIxVVGDVrjqrW3sREWnGm7Uv1tbNMnk+io8NF+rI
It6l85FX76d/CpsRabYhmO37ZykmK9wQT7/YgzOU8JVq/hP1wEx/z+AOCCaX6QkVROyCjcDT/qnD
39l76eSQi/sfk0Y1hVQkTCJCBGGtG3x4aNED8Fn+Nyxd7d+HL8bWkuDh3fIdHlC58fRLJ9ZEUJk1
oPDqOIFdK9DFJ78atNX0qy+aSzHNJMrdwltlFp32/FC3O6m7BoIALj2e1BrhNj6yaZ4Wd1Wo/mZT
0YcXnyJzXYDov4i1kmpThXlajxgP/fUq1SMV37aCUTeVYp7Ykag0nBVL/KDt3nY3xTl33bcWH3YO
hvRTky7KKdalnbDYAnsbACGnG9qNTI6WYICMrru44WmibaaRelQ9K8CG29uznf6m3dPjqitbQlN7
DJVvkk5BqGnr5FILshYuyK1wPl7kqD6gs6Z+JXzo8n+r0WRbw5k63YX7vfvlURm7QmrsDuiKQVYx
m8kjQKR/IIGmAYcAAfzdWm/xXnb7gL9JW4mImM2Mskn2EYELtg1oyh4rUg/F/fjyf/i6bQ/sKuIn
KqX34Gkr6pxAfiPcQKx3oxNF96OlNUoksnZ8JT7xsHL6qQPYm94xTodOXdCHFtQNpXQ1f+VedhtD
6zRuRIIK3tRYPPWo1hbi7rQNNYZYVY/Zpsl/YKcRU8JJAj1rgC7piCYxhAZGuIa2q7S9jYhfPFQ8
WquBErWLlF3VQ+Ox+OcrWRdQ9HlTp320uEHCucpgAXK8ZysST381bb37Q5yD1KDaeCOAkskc3O3Y
iO+ofRH6EdBbWhh+ZFB9ApJg/wN+MRU4cLSpLIJvwmFq1qoZkdvg28x856LVsi1Xq0R17k2cIpGY
CP4X4JTTYp/sOaVedUF4n5vcCDOQPkieIVwKXJyraDoTP/RAwVj0ogx+YU0Zr05DTMVvNWe3UxKk
pM2M5xR1qYrDU+nBDTzrT/5LX7daYJfVcs3VgAJTIamyikTYH1iQBlHpkUqCj7UqCdLbMCFL36h2
lHFj4WO5aPLppnCngMAE4bPSyOWPAoPcr6zANjF/28mdT9teKxQsRwBmtEGnTjDdfqcaSxV5J1ZU
CuUn+Un6qLyUkWLKKb/klOQaDcH8kHH4L0l6tf764H95Ex2v1qCw2+L64bcyQB4DUZM2OxNwPkjR
4jGvPkWmdUKT/nSJL4SsN21tuSX0UvLTM49RGIGaBPx7Sa/JSQWeM1LsRKw8QX2D7zwg6f1zkqKo
Ye1OLI3+nFe62BCi+uZcmXLYYTZwdIcnrC6or8Ulq6iL7v2jKFQ97igob0s20eV8TNz1AgRRtzZ7
UvU0Gu1L4ibv1JyVXOnplqkm699og/7AnvNugz2LltWMKNjEMSIbGNd55u4sSwXfaV4R/ja/2blz
aNdnU82X5kqeHSh8G+++4TnoIdqWDbexKxoRq2kFPN1yibsxMlmDaqaoehw0JtOeh+5L8dajpCJL
655bFcI9p416KcFq/ONigbFbu0dsdkjqKsGe48lRq1Ys7/0SncnOV7nFvsbDsxY8+mgiPXKETuA4
QrCBqqt8DLwHMn34qGtbwuKjS8M8zdSlh5TCUFilR/8wXohCqxsG+H4CloY+N2gN/4+8/rCTrsqa
nq9yJw1Yhf3GV6GfMdquDkBK6XcR4PoHiPbEWsvhIStz3EHFPfGBeptwo2vxbmtMQyHSw7PbIdvV
b+dS9TtuYxNMHSuINqvRYLViNrm/J5/RF/uuni+ZlF8csisFJeyvM/4lxWdG45f4ZC6qqYGY0YBO
dts0b3xbA7C2MYBjsC5iqoKuFUR0q8isMd6GXUox12v9XYepNiqIe4/ZIxFQK93zQFTu6raUUnBI
gkifkGJ0Q/AM6pC3KmL1N71k26ThPzoxBP+06tQncEZuztrRoFVjO7vHJd3bv371bsANCRZWnk+g
y6hppO85XgsZfVLkH04TOWN0y2q2oKr8EjcNr1+p8Q+JjH9JtPdY3+hWThyB98izVkyToVpp4yJz
dB5YRn5AZeBUgoUMHj5tswR28NBPgy097ewZRYhCy6PS6eoFIFzMFix9z/vuV2puGS4qt9ICB7LA
QvBtFoUOpQRVFrC+PM/qfwS14CNg9CN2XmScqywHNmd0ek5rvNNHW8vaaxzSE7/hzF9D1D9JJcaH
3hDdFTgc4Db+skrqwGvzRRVzXDsfKJTeSRVB2eqAPiPt2k/Q1A0xW605GE9x2j0Lyy4PFpMx7+q6
y2vMDQRG0eVYWlGcTRaaGBKsDluAzihLvkCtes7u37vrHHIDsNS9/wX9rbLOjsrrepGbFyjToFPK
3pico5DOPSQgShE0QAkmLKNG3F7WsdfMALAlUj+qGFpKV44CBPYtNprVTy4mJtKrQ6KXsdIQf7om
xX6J/8e7Sv9cSHOktxRxFAqHapnAOEC4SXCer2FYjME+d62/BI4ajZjvg7It0MdLeEZ0ojaWWchK
mLrSTawvNVp62g7hSiIpVF8SAsJyVYc+vUhqu3V0IJI9xcDz0uxS3MbLKYS0vY6jG2dCEGUCW6L1
ODJEZ11WAObY7IHffOqRovA4Wu30EraOtNAL+dWz6Wf0P1ICGBQpWxTCnNvJOY1bCPnL+tbfRhYt
yDwtwlI6785fu2Gq2zhUnlrsPS0ZjKs+sUFdi3444/NIfX8pK+te/mSqdPKm+bPOWbsVFtNoDeDg
va526ptNypSByCHgSBVTKhDWhYQ6r+tzm1dwi7PFKxYx2S2Bc4eBlmGAXaAn7uuaH4rE4FFzgIjT
50hMSDeJ9ni8U8PD9YyAXp+C7Znx3i2z/12jbPOnprp00FCuqTmO4AA9Ze1in38qYYLuj4E5WQ/2
oKN/MjMw4Gz4Dastt6HgsQBWGRnXGBw4gHBOcLQjZmMJoi9L6EsR0dwWBZKziY2Lb82AsyJY7Opy
Mq/kmtpsRXTa8HDqEz8RH+wI5dhgJjr1S7MDyWy7Yav21gM3yoIJBi+O0WUcnjOAAEnp0BFAfzUu
iSwif80O3O4CpKzUj9EK9fz/aMsWTrUyLeM4EdEiYeX4eROJS9DcudjKBSLhyJbLIvAQIiqIPWjd
oyOT9PpZm0R/h+iKlcEqHIhH7SiFVMwh6lJKODfD/YFEU6sW+BkN25ZgqZpHAPTDjYoWvzBHVqwr
ogpr9ybB28Eq+bA1TI/zZ3kBh8972TrkkRqnz9cUlfk6Cn6nwwP6CjmN9pob/R2Z8agclEQq3HEv
6A8S2UUpTasVR32GoIj9LnPI5e80NYzpPvLFkcXsMeT4GrpTP3d9+RIJfEsoDdUIDdF+b+68cWjQ
wXeegATHruvaB8YDOq+sGZDNM+DDKDfYLdIWVMHfJRloTmOf+XyUoEF4mPnuChDY51MRX2zR/syB
ppBrnTtAYy6cmKZnh/pTkCH2yz5dozCYM/Dd1MxvPFGE5G9e5USR45BJy7O8w0RnMsu34eY1e0D0
J3gEdVjWQwYmUYrmgKHj7yTWHpkAvVia/lBM7xjJZaTBMakkHLiT68EolGp9XDvOwX9tsEFYz278
ZxY4MVwZPUQf4zF1YtL4lazTEhPbV3Ny3JmsVich+IBJGNOB667KDEh+lRmy5oUdlPoIOB4hdUj+
hwp1DyvWiPhaSkr+Y0BhC17XdeGBhd6vuqaeW6N5xRjeYzKNXDZftcUqbP8JzybL4wZD5ig/XbgQ
ATJuJ5oQDiXp7XYpU869O2tEnsg4ulvB8f16+2gq79lltXJOEHjRNCrXYNjpn2fX0X0VOL9Lwu4w
Y6aXaU9QV4TJvYROS2lBitnQFWztni87yOK/uwi2HULjWWTo0gVCHYCe3S0E+qmUnh8Somc3+Ptm
UQBjTPoPsxRAgu5jlXfR2qL225tyNmgORTsTK+3Y8R9jel7bALGXCnFzrD5wsjH2/qctcHzrkVJV
LIj6Ga0HMMfLVZwmcNwRTWW2Ib1PDOmZxTEle6ax4o1xbGWNLyNCSKrn3frR6MbNeAcU6NksOWe4
gF8BPT5dXCnWax5I2DmvixfD5fx57HNFr/2JEB15vGiy5dKq/Y7zsN4WDqHsRhPnsWnTB3vIBycE
Z70qt8aflsVVD2Y51TbdGBB9R3ZON2UFADlqZUFS2vqf6B3+oyPe3lgooF07Ruy2xoZ9YB8eMY0P
jpPZIyco7ogiiZ2o/ED0jzK7SxlHuBbniPfuqnLLy13uiAtmr8C/vkhV+WBnqiPZ6cK+bAoJGHH5
Icc+NmEO4sZ8SkGlRj9SIPGh3+5MCYx3fzg3Gkk2Nwx9qPW+k0pmNVsdfWOJVU8rI1GCutKtH0lY
METPEjyjzYxkDHXl+keZN86AaTLgagZWDWbZQKLOBtbpXOK1wmkL4ZhTn+aIKN7smVQMwUxX8Dsx
QtUvTXkngx42HgjWwsC/O0ND5FO8CjPLg8Cj++uMlc13R9CC0zEh54ee1xOeMHq7Sx/lg2Qsee9H
3g8I2FhuOG1HLLUhu/RZiEp+as4vvhej/pZnKlDGfqTOZuZ4DhbPhATpj2/r9IM+nmsW5/UQ8/oz
hw8ZybiW3oITnBgE4sCBVm83+AvoMinGMSmZD5fcMQILS1Hma35DSELErXhOpIgjdBwf6oxC5gDg
AQvQo9Hz9plMDkNo3APsRVuCIdtHue7dQ+VOSpzFIicC4SXZWyTOitHfHCkrV1vqThsTI4ZM1Ctj
1FU+MwNrebjzPbLePbGkIMR3FjLh+XgJt6sy0PMNlSTJQISsCTgw7X8k4ETSI/hOkOUuz0p5yRz5
ceyBnd6tPgU9nDGVMbGZgeLHVD6jyrIzAl/YYgCbEQdokG/qe/OpcpmocEkTEP2lZ8PvaIbh4+9R
SHHHvfQ3Xb/qhI2COZwCsUIoQCah7t9HKgPofLD8auzhrQag9Noukr6eeLzywycAi5bfSgBFOamH
fPyt2oA/DY6lOntETiZrR7c/RE7j5Udqv2Ov2ol8CJehAaVgdfemo4qIJBMUPOHjzmwCuI6YGlne
aU7sCPGZOoCutSPi+vUVIPS2fKuj6lg5I6+EGkhDBqfZPSMJ6ExxzcO2p/A40AwYCrW8/2YbJjlp
uwmYduePr/WzvP542iB5usbNPJbU0RH0bdc71QP+tTuPppxcnOjsWW1eLZMN1B21BS9c1uKitfqD
UNWS357hN7LwQL0QuiS0tqtECjZ2fm6Od/pxUdVLkcrqBhoaSgxsPIgchzrm+cZRhWHS6NjG0Fn5
q8VIT3yu2TJL2UJxEIFZVuVt1Lj2uc/L4jJZmJwJ1GHMyqInhqzPKhq0CslMlPgwCcLM3rHbHDLS
OJiX3xQZRmUhZ/0/OUDRxBXlpAtY+qYLo+iKKLP53O7/XtNu3QQELvabjeJj+1Qsj820dVkyHU8+
XLSoYDsp7Dcr99uSeHAh3VZf2kRNNRPjxWpSQJbUunaFRmz4kDzMZXmKJrjRUG7XmT+aS7YDQB++
nPtzmKki/oe7E1xSC8uhl79cz45YkjDmtqbBEKFpDOV/9S6Rl6H1sTeueFoMhDmHdzRuDKpqkfl/
ajjB/LTH6TpXU5B4rSCY3abhnVcwnxoAQFXc1E4URADo5SOyKQzS0OkmJ3zLxw3IVNVppuafHE9t
cBENABJfn6j8+YnBNsfbZCclekQ46D75vVrtfMnphs4VnT9tW8/YH+fp2YWUZHKEOj5O2VrxZOm9
HyNEuzYXocuR+aCWGPQhwLgDQFE/6cCl4Z6d6JwTtxxx5+1lm2r9T60WusPRtVGBl2qQeFtZGryD
WNCKmq7IapE7TVz7gq0qfKsH1XkH7+/tfCCRHUUjajhaj9rx4Ybf64FJ5aAbe0+65tasjBvjznYS
hEVSSo6kPiLK5sz90YK7G7IJw5oMpZId4G09N8ZSKjB59KWfPPc9LRtSt66Z46pBRJZ5Sx+BgbKP
vhJgVEvB7d36c9skoCmbJBa2gdg6+MRhMXjnpGbHeQs4zatmh/mZbnl6+TtkUyqmlLcVzK7odHcq
pIyZs/vYI8QGPERWiVZinzjJmNDrayBPFvYnIx7ZLCSfKyxSxjdv+R0t4OIAsbruIdbJVExQK4q2
Xu7OXPHm3+p8isBLcJVVzrPCSfPY5ziLvxTxKOHd5L8dcFf/2hbdfLIk895zbx2cunFpHJGD11g4
ZHYwzvAoMsjd9hT+r2wDPZj9S26cZZALwXL8aIr8gH/SLjWoXKzNYd54+JndfD6F1RicSqVzSnBy
Mukkh4sS0HeEFS5K1sqpPifrmCVR5jyfGg7kVbiuD/tCYIA3Uenw5KSMUjH69UpOOpBHhvqGYLWH
FoHAgvozb1HVtz8jLXQnwV7RbiOD3K76B+d3PdqWWRQZR/dtbaDsXsxPR2I9AxOuhp0RiB24Zqdw
v519zvJ74I4BeUnhiEkHSOvEc5SeqIJ3eaq0TRCe9vAQqUeZjOywps448N5ywEeFXGcSSpe/SUKH
PAjxQkVwwBONhj9Tb8PnlPrEe4m715U79Zc7hLfJIyaGX8+OUhNKJqlKfrf1QqFOhNZ4r9ddRSF0
veP0iFMB6wdVcrY0K09/qx7srIRAT3jLouURiFvr50e8PAqja7ymA5CMuVnsl+Imxa1ZsfKQpJeQ
kK7gB0wZfJVznbwUq5Htf+WTczoTvy2tbnU/IzjVZCiVI+THhkNc/yXh47hX4Hp7QCEbWpQw8/Uc
n0sMVbqhPHS0eHSLF5E2c3zudAGWamIZUXGOsBdglXZUp/MAVl0Cm7tHR8Krkq0vBb+gGCjLxYSZ
NhtzjWMFFI5T3LowXHo9FxWsESA6ZtyhjA0xvzm1DMA8IlVDhqPPFNi95VOeNDniBOGbj+rmq4v0
4y+y0YGoueKwNX3j5Ge+M8zPSmDQ6rbn5DGTFQJ4OFRW1pt5aHpeCsui1+PuLZ5tTA9Z4VycXtYZ
XI/nFTrGkwkfuWudKsrB1tdTF1RtXfO2AtRiyTthqQs1rDxY8euQHyS2i0wHwJ0E+dxwtgXMkxJ+
dvYsZfofqY9D7k3HIK3LzZmLHE/NQuoPSSW+hAE2b0Y8Jbhu7fVZ6Hj/FzE4OcGr9bsohx1ASYDF
wamblJ0B0CCuyDXtcW4FsXjYMSnCYcSoDQCbxGve0KlivhUXW3s/lSWGBgv41WvwVlTI74FoX4Gb
5c0QpYQq9i7UqOl+DhdfipnYwGXetXYRaXAqLLRODGyO0nWRPeCeRlABQ7MQg9e1TTBp0h5K68Zu
s3NWhzpdJOldOBacvLPRBWNN0ruB1qqB/r0wCLY9lrl9NLJT/2MLY6Rn4LBB/Bvh9+dwos4gbVOL
1MFtl9vnbGWucSVUs7Z1YI5iDjJoVACA4XyDFGAJble5vNV/zOU5H59xynOnoz0zvSykcQGPUU2q
+HI9zZdTS8V1T2OrV24Agem5fg5ChzGRrAogBDWWKPkgk6la2FQPwOX51UbF11+cTOJFem4zcB0z
j/tG7TiuZ/A0tFrQffeJq8tst9TicKbX9J/3ebT3kD1Ol/sPh2gLPv0H8h+MBw7/n8cOVUeqNbvv
x+CN5wD2ps29dr9rU3Mjr9R1dNkAUYfo0Rw3RDogvtpcZFtqbiSsZsj2X3ZUsWC6bniX64mHDIJs
S/LP0S7Qc+SmSTdn5UOOADVfslPOv/urBW25VYkXISHj5+u7KlRzTLnBERVONIOKxFUFcpdHBwwP
8/JfXF0AkM/KVEyiV573VqiGZbBBOei88P4jD5TxVTFX/FLH5F2DSuzftq+CZmhz45lyvO0vjJ0s
GVzbtNHkeeMwQNZ7YuBrsnS2cbP4k9mCuvPQySWiQJ1ukJ0p9cUfa1W3xbz+uIVVrNqlujo1l5cW
kqXiGm8+2ie2hH9FJaGKMuilY+IndJZnza3CIKO4A2CMcm9blXOd5DrdSBlvoc26Al4dFo6a6Wy9
GB8xwbdSRr/RZqwGdhe0mTWIMxp37lt+qVLejKTDVQYCcbg4GjIswAnUeOCnQkWJCOdFUakrFolV
R7BIm8mqhn8TuGTIJWgXFPPrFhTyemXMjaOghyRq98KbTloBjoSPfRmqqENMv4wZuEwsTiTfgev9
cJ8y3KdevHvFT6G9wWrHg6Av1/L4AhC7TctC0g+9NN5YwHjNLSRa4kJ1ALh+IuVQD77rE5a1o/Pl
1/+N73GZUwVwjji3xQTgNQgIROEkDj+9Iy1q2sF9mLFQ1oYYdenaX0wX9Plw+PSE+vc684Wolxsw
Px/eTrMCdmpjNmv8G89Fo/2D6IeapVnIL5ZNdBOx4mJ975iICTdvqPs+6oS3ioQWazxdpHt9z6Xf
o44Cb92cMkgAlluetvtnjwLnvJtFdjYl4KIjSHyPW/yiM6HfGa6gMfexTm5g4bd3wYCQJXlWJvGp
Ks90/xmFIe457FeqYrJa9LR5MSKNtRCtLU51FTf4bBvp2Iv9x75mO6GALXI+d3pn6OsWrWT5vBhq
m517LVXkNqD5yY+GODw8fSpMtFvJygTtl5JGFWGRwrO+PkkfTu1ohaDU9uUyxSIM4v4GHhzHuF4T
iUoasBft+0lVwy6ooX7zNLtr3icVaxJDY2nYQ4enD4NXeGQbY7KXO72Q0CafmpBSRRnXgY7EsFed
a5tXWIkn658ZaqGeoZF/09UQzynyukc34723bHeEQIms36yxg3aPPjhzZYaumyr7BCRawuzNo2Ok
2wHvqdzvluL7WzDZTd2hym0sMQ/4HgrWuGVluTKZI7SYMv+/LGrOQ2r8DM0SU2O128HxO8GstkV8
dUEogBG0E0IxNnNunlt4Hd174Cy6ULnysp7EHVSq6QzNH/frG2MRw/w6vLsQh8smex0qia1ZriBe
cid5f3Zp4gM7/YhtqnhmfNa16HPwTAgaQGVecg7LLrvMGBkVoRfm0HdtQxhEwv9BN2f2uPR2ToF+
w6S4XemT+9KhT+a2e0gyi/PZFgV/h8zEnGSC6AaSd+zpWAEE5zfBwb+P3Enw3TSg7JrQpwFagNtq
rFkTXUdtOgWhJcbMJq6CMy+kFLueu4Fp0ypGFJHdJm2utLIx/l23VORVbf+Js7sS6Kl1xe47RRCg
KO/xXv+1lCPwLMmLA/qYQfiXBRnqa0Qztfh3WP35q7CA0yMSIE6+8hGSBa48X3UTBWUolaXI3c9n
TSrH34J3Ksn/a69JevtEbZ8taKm0kRhR+xIhm1gwElRLbCktJoJpfCAzia7tee2vVMHXnQqD6PYl
5wEPbiRrJSxgo84YSlCHw0WoGFOBQ837rBrnpSBKsD8FvgOExAHwSNtyrgiZZThR7TOghr6mj0Ut
/UF9HDo00ZaxVQ4xay+hLRckQ3VNI/GcloRCq9u8zzQte1ujAmyTJrp1SMZCf2r1db2N1dRfBx3h
SWZmST6C486iwqX/+jqaFmlKeWkdnlTPlyoyG7lEjQKo/0PWDj4WreCQw50oVocJSgLtJi+5z+Ig
rS6E9mweDsYv9rMlaPgsZGFkalUFlrd8jg5ZTVVC+wfdbKtMZU5uIGGt9DLeOdDrj3wA65lK+aLi
LAo+gzNTWyogI/VzzuHLkNapmPc7xqauAk8PKSJPTs130L0mKA49gdqSj5YWQ7yqNqj+5hAp6WwT
+WtvINGqgMn0RZlKdahmfN0eqrXs9j4kdEOKyXGndwD7mwFRLT/7uW+3k7oRS+C+J6EXttp/M5Eu
8SDU6peGYPPSYaXuXb9tRoHb1prrijx2lP9+tMED3d9n0IgqkYdd0AIpzv9I840nVTKP8ntE+EjA
dr1IN5iC3Fo+y5YHSLL+5t5Md8kQnuIRvizMWC86yQNcyzswmr1djZ9BYkJdk42H+ccX4TdUHBrX
oVFTRpd0ht6Z6S4IDKKJMSDTAhY2n29UrduQmLzpMHPYuqQ9srt75M4OD08W6jWSrhW26Q/DJDB3
TeQQBRqNnrrc9z0G6aCbg1o5KlGeiDPO6lc4p23mx6fyA+fvbsj7Mrnb/dVH0aTYoyO0/lfI9ttz
/FLnmkWULbcsMiAEOEmPCIe3icUyArOlQEWqgGdujp1FGrY2mKGcNVyF0u65m+472V+izOoUNqkE
ymUhcsJVm8/mN7rEFyr3e2F6X5+QnR9JUYrY6xpBv75ErGOY2YOlltanl2eU4dyFievtKq0k6eUt
/A964Y5si4e2S19G0w0ke38qYGK2A6Nmkt65fKCVXFPx12AD3mHafoF85bHJRjwX29UycT9KNMPS
ZeVUWAkVjd0X6anrVRwwWrrbhG4SxD4IzdFuCI6zKpA5HIfmnfensjna09nQ084uzg8kB/bTc/8p
ecK6gOItczCLT1zhK58DBKGjgKjVmVOYrNnE9j/rG00hl4or3ZKs/B+XURFwdjZQNaLi481zwed9
CQNGr2BZT1dQHAeUZQL7ii4QDmuVZ9tylEpQ/KGwCIb3cru+oXTc7zew5fcsmMttRBLzSnTgLUE9
tHyxca6jGU+xVqrq+fzWd37jDHuhEwQcCJ1It7YRfaXw+lNhl+J49czoKPS+yNR88wwV954dGmG7
YOw2zp1fYBsYkWz4AJd0hFI58QxdPUZ52XVa8hfDG2kn25LTspPyQklRzlVuMbuuJmViENnkcv9e
rBdiBK0BI4wH6lovtSqjAh3XHoXxLIwF1AGTAu/M5+s4GOY+9uE9SpfRRv5T93JfZlP6xJPqBWzN
1xKLiqAeLFzRGKs1Lu8sX/CRgxB83pzpAeKBH7nI0UZ5HmRMn67CRWKv01DH25zI03wgeClPB4M+
q0/Qc1+9h8m4X0+7fWEX1J6jWFb8yFj6GwYPUqQRExhWYmb8eui2cNZgQDYzF4UjFM5y4BH/0jlg
P890+cWLMSQ5LYw/fTzTNwQ3T/UiSAqbRi6kuYraYoYvOj7bhwVXG1y8PwnXac7rCErfPrndfleb
a39J14RezRsCI3NXPq4yxKXB6/3MwmxFPfyO8EQhMRKAS+oTR6JpGHZ3F4AuGNSveaAOLbdWNVUf
S4+F69byH317YRT9uyl5ZwhYPW75UAtXcI/bPltqSQWTpW/N6eTDXOkCJtudcyCzuo0JMqnH4teW
MsdqFufk+cGtxnr+1IoAFfgEyfKOB8kefmtJnZQyYBPBX4t6ftkegaHq4gZ01SNuClJdAvOxkYAM
yLc+lNLcRdIsUzms0GD1hz02TFQ12yrvo5u/mMeN9w0r2XNtbib+uR93dQYaJVe5jskfZTZ4p+MG
0OUs23rMYHGX/UCQVdGmqf6prA4EQayxJp0XnYDTsBFfvPljOGObae2ysdPh/uTdYZNPsW8A7/QU
gh+bHPsHkTXrWTvFlPe50JVEpWHbxZak/idE34Opm1Von5S8YJUSBk7Be/6yNsP9m37zcKocTNa0
Mrg9kPXJ4T/OWDOrV5UnV9tq9JriCzV0YFPQ1WTZxBH9NF1zJ+huhvMkPy/TNzKeJu/67ihxARYR
oBqrtjcGe2kvhUNYKofqGdxGk2eyTILlDFfT/T0pK/tsT9bilziUr2Cf6OkTbZQqK5ETvYdA+CD+
cAdmmwG5SPrs8/wOqC+rkwEKmQARm4RJNhHx1jwxO5c7TQSgE3TxH+HLMBGfjrF8zGupgZt5I+Rr
SMs5Ai+fHOH2pzGPjwQeMKXS5W0JHKz6H3tS5vapFWRQT5caj6IkMCYSMhockBYhpORFlSZMZd4x
4JiMKl0fz6BumG0DsN2kn9WDRaip3CgMR63Hq8kXddMht+PQi87GFAmF/zR+NCC7rSI93++RyQOK
vb4nCb7Vl1qjXrprMyP6GHu6gPVpcq8RRjF9C7id8TCD1V3Xjv+sujSCZ/SivphkBaaVEtFA5eKd
XU3t6E6oLkz5ZNSIT3PqPghKe6rQi9bnTxOUEkAQ+UHcz7Jsa+6PEWAnOexGm6s43Pwkc3SKub+w
knbVNdpPvQMYaPA/W3MYIkF9QaAlfOvotgMgrsyViyvA32FkEUlY7Igg2OC9WrTiTthCqxTyDU6F
3I0jWj8AIIK9cVc09YIw5SBYy29H1iZ579xSpFWximjA0i1EselqpT2rtn1zTDN4ugHJ9hwZUKLn
QK7js2hBRw7gCltwOD/4pnTnQ/JTX2zr/XJKHzYnnHSOZo/ZG0ZE80Ph2iq0O6b4+u8N8DM+VVRA
X9w7HfqyvhMxXiV7XYNmXN3RwVFcKA4LDpTgIOnjXP0IR/lAyGji8oNH6GjgZq0jjjGzFdeQEuzO
Pie8SUjsgMLyNT6YxKX875AOev+BNArKx+pCaDEl3fq1qKi4u7evQE6jNotJrV+PRta/LXjgpvCP
mQF/dc8Be4vy5L5nA0UX4o7RfLioteL7lWoJNHYTpMaR6Wvd8Q7672H2dUvcuIcxLC8Co/kTb1zo
vzcJafhrmo1CJKuJWEEJyzheKl/7Itu/uAONh4CC8rtoQvOFlrWSJpIW0Rh1JKToJYqah4j41fUT
E9JH4nrCBi3eqKZ/rxutSi5bYpoqlni+3/VhzK5MuGxuoW8qJDMFKzo9utTSjWnhLKqrs2drxuZi
kCISxOixkezxZ9b+cVbjYB+pOVSC5UaLJw2SI9uxC5WIVLdBeP5tZ8qELQPqgcVxXM192XzHja8N
gHPxLXRc40l9dOQ+q8dDU3fFhKjhg8NMvmKY5HduCps+TNN1tB0nO6UJoQgWi/jGl3QpDB5S5hh9
/egPSpdXEx+VXp+IaEXDNa+YNm20KR/w3OTEwCU0BbcpxSVnV4puRI2ZNBs4EFHS5M1dpDnU/ZQD
DAJkuY8TvaAxo7pf/DMvUHUa2TY2yhUuYOMbpgVv9cL7roHCu2xAeLJ7tFqGBRti9AxvLFOWuwe/
u+Qi9oPy9baev9OKPfhvem863mMXlpmhv1BJEw+frvGgT7dmJVtTuMhebO6jnbT59UMcYW+/LfHu
3gaYdFx2E7ynoGH8FY11WWoU8/YrFMp4omA0FKXCxkyyBt80oq2ukJufWUpuSAvKCbxtU/iPZlPP
h7XGsoYCX6YyzewJjNSMpzyVSpTWH7hDa+NAJF5S1i93LL9ihYkplvWuZ4jGZ0e7K3qngxB/p4k+
P3NASzcPG5U1EghtVq8PhIdu2/IWvSPUZWiBB1pmFy8wTT0WqvoqgFFyU5HTV2RaYQdc+yhAdEQv
o31ZwArDpaAtVBJ9eJ2f5AuYBTCE76sBg1XqFjwKLeSISPqCjilY3B4zmWbEG4xeNmEZlk7kGK96
ypvcxFIWpyiX5+34k/PgDOb01EyXsIh0O1idx0fV/Q/ozokTNeenNEnOGaYGALhdb9wmRhK7CfnC
Udes/Wp+kwUT3If0J/ObSKg3GEv1yXSM6W4fFFAmoOtSapn5etA1ut2CmcjRLKF5o6F+H7DVjDPd
YdooYW4n6N3AXZgwionNhbHAOJbUPkRlo/wQQC7pZXVHfKuRssLivlAG20wXyqCWFgzeZ26TivYL
kQdUhaFDn2YtREx/5Rq6drBS0irkUTEq+4KbrcB1KRBxFkXZrq8sEykPP4Vj/id4QuFBqwOuApek
K5pjDGvkfico71QJHhOCFQGuKVcmUvnrjJTTl3u4Q9Xv40EIcxJFNRlGJ4ndvaciB9O7QZH0z9W1
CvdVzNraVCU3u8/Cmhu4J6+qZhyd3uek3thKWi+jw8LkCTr2ZYWablt1FeaRttlD+9DaDMS7tRJ3
3TIGIyaCPwtkqic8Tq+yazKtV8CkDosGANP6NYjwzAkd/ol74GcW74jxaJq4pYSYxRfxcYhCbiXR
WX+PNXelZxWKVUr6uCkFSFdHDz283mE6LRzfaXwrsL4A5ZtJSVzF1f4IXJBYayPHbMpesnQiuqIv
Stq4LPzJKvJ92KeCLsCVsHWz9voD6J4nPTuVrWzicbKUfMAALTUd6DANpTohsq2p2YciGv7UKbKE
wg27FrvyTTBJZy2aOOY0y5Iyy75IRPGRw3yFLChUz/cesa10BPSOubpwie5pUK7f0g8jQAuJAVfB
VhqALAj/d9xWv1i8gm1fwk/rxzJ6qKZaqeSI+tExjfovNwvca2h6b6iukRIanKsaq2gvU+7FZShs
4A0eWyD8U7DhoQWPpmbo3jgFew5DdVjt1Erv8EEtsCUB6VZFARSD4TgWDOIvl2Qr+4P/DvxnXJHQ
1Af+P8D5Ne8tBpfHWMy3ez9yYsb0Iz0g6u3coBdwmIhHVfVNaD6G/Vz1gCX5ruzuRIsnUtQSx5GW
bE2PSm9VijJstTTqGDdPj1sH6TJwA0CRidzPy6TOdBHy9DQMI41pKHHlaRd48z3rSXDbox+hV5bK
xYJI24B0xcyJOoycCjv02afpi8rFiQhqnE6k58f4nQx6cVwK9dQxA+Uz2ah7zCX+zGrN5TB+ffsw
2DYYQza9Hz+HfkmOL44jGEOFpVTwotkIOXGEHI+KZ1liirzlRKlVzfCWaFEpYmbpHamnvijllhLx
EBvJJwrzljMd5wGIhjAc5FTsio74n+F33bIuzAspoJfh4xfCcdVqP0h/dFXjZO2RXz9gtgJ/xnpm
gpq7PrNV4QJnXtmnIC9U9AS1AygLeB4uQ873PB+xebMGNrO9kHpoWZGgTLnB7xqlfgL1Te8gw56n
AuIpd8+ZwzzKQPiwUT9/vzwldKrR/R+uyO4Y4znZKdFEiU8oiD4Vs+h0kwQ3x1AiouuKUGhIA/H+
e3NGU+wRK3C4qhzIbEKop1zzAvnJq3LNN2gYItqmhFifgOszMgvzSp0TaXvwfa13ye0fFfWT3hjW
1P3f/92WB+pwPc8bz4GJkOFGqVNQBNdhBkdf4dlJCQ+TyLhtgTQ0+Fdkx+mTD5dQlls+WdWvNTae
6JxjGKOOB+YnhX7YpK4dD0k254g5/ZT+TZK7gO6stnHhrEezxgy3/MKOWsWmM0NbrOTq+8twAmHV
pRhEd9Ek1RhWpjigNv4hdYZFnu9EupE8B9l8WZfh8lCk0NXIpQKDvJUCtF3VXncO3y0iHRSlu5pZ
CkjOfLpu9vnbHhxj0ChTYuqUjcBmv9/qPMqd4XV2b6LaLSJ+6+OCrVk8pOmpRjQFuScHRiAF5kEx
aYxwsqVM27rMccWr2WyIkb0ZHAJXRkuwsqCfkeGlFoDzzkcRVvCruvBizFNyRfJA47ogb7bZqbZN
70ayTqWfI6YhFXvGRSyv1s5z6Pzaj8Ef3RLKr3F6sPF6q/alxZTOguzPIE0y6dDQDkgOIMwCs69+
/lA9jy1tdQPFovKzv2WIsVxAW5UWrX7mOoHOe/D0tuSvK9JshmPcd40UCE3WaVTIfcQKB2rXgmVC
ng+e8KOZ7On3v0OCP9ctcqhFsBc+HWKMx+AjMhEI9V0hqUped2KHhwWNm0gj0MCDnFp79WqCpusG
zi66lAowkSD4tSzgmnUbDgV03B+QoKNa99v7UGDP929QCG+jE0nGvZUgQwtdKRUgelFfboIv0JuL
b9OqVjZgxmU0ZTEPx1jS/9Qn61zU8Ss/wS0JIWKMhsFs3DHP4WXVPoVAjAstrVw+lsmkpCXlu3sE
7cabeNINSkI8b+MIBKb7vnr2/AeRh3CoGa4Pzgqj5inkeszi18LaKVSegnaRWaCIxX1SiIqmpKsS
D4tpJidjXDFq0fKZIzuIxJp7vqJWNsg/X3bVwMgY4n9gQFe9ybGlchd3TcIMv8MOaeWixHSPB+HZ
kN8MiFLRqxO+5haLUxxPgAp0CPfM5C7G2THabatv4tWk6EmiDlCNiKzIq9q/ZVpFyoZs9zIb9PYH
R3LOULeWZZ5cGn7574ei39+PuSPIaRLo56xgNlnPvN/7e5t1ntLvIOxaOppiUObByIZMAWRz/ZV8
/d5uHzDyu3mY1tKM+gpsjWEhCIMHy8FvBBPb0VoFnbr+3axhEKF5zG86Rxdj/xZUX+a9u3Yi7THl
aJ+GrlDOpDp0u1EM36wgJ/mQTJ6ot6e0VEyey7kt+7dNaBuWVtwMShtWLNtE+QHn0DP4cBL0uN+x
rtqJE1u14OtFB/S3h7PFkPQr7iMA7yIoj1+WSMbHQql6jXM0+Tlq/cFErfuet76gL//9UB1sRkaU
meftJ647+3Gv5YbgaeE0mI1QIFGZNs09fGlXWkHCXgCdRCTIC3rm6SOrwSv8PQRVh/uR/EKpDS9w
tU37I9GbVAArb5f853DE6SfDobeE4O6Q99NjintA0tZHQSRQCYtDjlrGDjxl5bZGHslvIcLX9Y/x
1rcjFfBlA1m98BVVEHQCUB1rJF2vFU8lvJGyWq/iZCsXBZsnhfjBBE4mbrWDfsjUxm1/UzWi0Znx
giZthmsARJH1OFqW8eyqlvDdZ5lk8WJUCX6YGJVqJuI5DD0DKgPw04jfDN94TUNgzBo1IOozXJdl
nH917evOv+lbdh66RHTddcr9c37ulq6GG6Y82TSCjSDxpzrPLUpiiqQfSCNwnYFf9neaPuctftEj
s2u7eG+NF9AE3hNJ4m7Dod11bVuZQr4M6unFtmNi1MZycK5HT1Ooh5Xyp6tR10KUJtADJ7H65pIr
8MBsY8HFfcsJ/wMxx/KXbHk8eULDqat/z5jvZh9aqD2esq3Py1sggjjeh3J+fOR1h0FnUJUuVgcT
epoS2cwrQL1EhEYemV6bu33DzywZN295j8aJuJBGLA8ViRBoJnvgxyu84not6OqbQ+xkOiKhYn0P
FKn9gTv7oWeFBUCAQYhgAcAoap7qSV1+F7nTDCQVhai9vk+hCiB4Z7JXBJYMwDulZrTVnL35BlAC
8sTPNnFW7GR25lVU6Vs2rY3utn2Ban8NSlW5H59XR8pfL7/wGToBRpbvtZyGtVY90K197QFe1nTU
R9jmsfuEYG+ldC60zTxmiVt5OQE8KqxFaLredDIwEnXXZB0XWFDgvZkTAAHXt1/hQtr0phS2ASJb
g/N+QSYIJgDpRiiwXYkUsOOL3W2Az0Lmdzg4Mwtyj3ONn4rDQ5X4Ta3VMJ75HdIeVVadfHyV3/Ts
y/kvPxSnPFbWND658cCYr6do5A40hL5mlBwMT6OPqSS+pTxzyDJJt1cV+/hHDErrQXNTTfEPU0up
jkz0RvOBBINZgufd1cj8l/b0nn6zlsWVhY0jGUCa8aiO/b2MmPN6Gde5Usb0+u9gyFqyBbjsXtj4
HmNftcDlkJgZmW1+gs9xUKu+FEXfVLX3tDfVPMuzipzCtyNORJ8cbtrwN8MpJ4UDvNJ1cSxDKPpw
PQt24eMgYFGwxq60XgJJJ4lJyrrmUKDIvu96VrME6EOMFxR78as7p/KtzTxnjcDByRwhQ8q5zUpz
TvRgSfmWau+JGExWZ5GEda7XPX4JxlZxXUZXV5BAoY9+fsnd7giPBPMNEWUDoluwHxhuUEByDXR0
08yXEJE5ERKtkQMLzu8IUPuSJH8vBBRw/lbLaO9zHfT8sfaMeP8DAlTMGOyTJuIFv0HZ6FSD0yn0
XkpfEff4NpGWuxLz4G4u8fJdxTcc44LYVTJolDZBObJrfYu6EgmiB34VXAS6abZ8s/ihHmuhr52U
liUUraj3TcLDiWvMyJtgTBjQsE3PANFRygajl2snVGYz4I+SCRbJwA9Myeyt8ntHZU0w1Lp384HZ
Xu43LLcW4pAHfv32j+VgF+1dXn+qW7K/LqjC2PklaeWR5wMCCv/n36rSpmpRYwsPDRudRDYnjqWl
XE+lnF0oDjMQvgHsXMBc7wyfmYlDNCcht9uLl8xftks8X1UrMgQClZButEJu2dmf61SfFtBpjIM+
G/PpG6ixeYlysDgYkzmfV5KlLky3/RUJGJzHp24j5aoni1J+KdNBsncnmbYGTkx5ST556N8rapx0
+l1s4e1KKgRQQvhoGpMjnkj887mGJxTFTjj/govEkTG06QY+jGQxwnWbIWtKhSxARQMMssQVzIaG
OO6zuYnMeDcm7cWPTSv035dtvDtQer0hirVTZLIBNMLlsu8fBcRK2iNDWDWkSC1gPch4yfH8LKcA
e8rTKd+tqk1ao5J/DZb5dSdbJmv8PtrCoZj7NHzT2wrYS3zhrBWM4xYkJBCAKauPetmTioacwI18
pbRclUZjdUeruTDuHF+k5dPC9pP2nVDQ1ia4giXHqp1gwaEsxEvOkOQnweGJQJycD+lqwUArCJrO
lnUFjLaHGYnsjJPuPpt6L5I5yK78eDB+xce56YrwVWLZht7LOg65kY94Es8fL+XR6K2k6DicqmUk
yzzpko0x9iLCIlye8mgCuvOHO2FNgMCClCsf1b8k2r0rnj/ZvU5pKqvE5BAFf9Jv6OPNuQg2qgAw
UZHucqK3PYDBhjYJfLd90F4tCQO3yWFKi2tl+iq6q9eFwia22+EkgKFn/duLQA0fHx4Qfv1VfdrT
eOeXELgHb8OtiIf13DkGt4c8ec/9ONCcg4woc9UNpHIbJr8kj2YoAePuoPvXGZVN9f2zQJcLEtQp
JQa8hFJzA+AVhQtbjx8ub4zpB9wvJKfqVSEdxljwcxXfRJFgwbaSVgeTCeC409JdNUpcAJAM2Ndg
ZhiRyw+M7y2Z36cm7sxnFwDFo6cNmWpUIY+QpEK/S35yyd93sQgvf8upbLaTsiIggYk2vpSTGchS
meJoeINMgBIec/OMxIT2SSkeIW9NY0eB+OvkpCWEp4RgjzrZYOr4FFU/IjUNzSPLPTnkNVaM2IuK
fscQWqNep7jIrMWmelwchVDjODCBcl7B4Rgmeoy7YaGILO9QRjlDB6uA2KzFYytRW5nziiISmBRk
SNg8+3MvtddULW1md94NktgIp7jH+u/NBDQgRnGL2rXXRRPVA6K4AeznOzge9rvKC4O+vD+iMm/m
ZMUxvOZX3BEb4+ZrzyqTsZb5KoJfD7hfftoht4ivfETFDb9Sc32hIRDqNLvUrZUBqE86SUe8oLba
6Hx+kYpMEky2Lbi37oGWgHms5aFtH7C9R4IRS270uTrqsCVdM+7VkpL+XAy/XF3W4k0KXlqpeIPQ
JvvGi9YK9KKjyNdS3E9Ja9HyT9NIak3PQV62swe8aR78UcdX7tDes8WExcxj1Lo6KmhEkBA6VLKN
CtbgmOoPwSlEEClpSVTfebDDOwR0zA2fgiLU4bzotNUSQPb19oqk1Sa0qH6Oba/Y6QBpj53kKQq0
JKfKrd5FaEibp15W2fCZE/2hktU119LRuJ+wDmRpixjR6doq8MJNUYVdeQfAk31ve4svsWX+T0z/
r0p1W9gB9u/qj50OC+afNKudVR75z0pggAM8vPBP55qBCp18Bln/M+/ZSSR7xQxeQgkbs1IZWH1G
nJPTOLLZjQ7e6uTxgcYzvC9dDLSYnPvJh5o/2vtNN4OWwElBIur0x0kQDs/a69u3pgOSqG6K8ULc
EeG4OeNn+24SJeMaYhzFn+1ZUx5xDEyl8HXZNZAZHVQDBcWwNXeLJ9dfPMkkxhTzclS0mlBJe5aG
STZ3M0NnMYCOivJLf++ESDlEXP4v1w8HX089nBWmTFOHNuZ9+PNp79zUT67Pw1TmjatqkiDHPqb8
Yiy4ZKd9gfTq7ITquDCCz/u/yojJwuYC9VOdHWPRX9vZ7BO9dOX9PbILan6g7eLB9QuURqiWLFsH
RarqwiQameOeGceacLQVxEP6Qdc0O5jkN1XS9kd6a4gYM8tty37fOiV8nuP878H2Ox2jJpOgCS+s
RwgoyIZnLq6cNTVQ2yAVYqy3brGIwL5/shF4q1KPKIFF6+KcVi4lsNjUmvoBAD8BtoSy9hkJtu9+
AJCZuY/ya6bCgBDY6RzEJnSYChjh/UpYDAOzc8jLTHCGX4zDmM9iSZx+IaRH2v4tHi7ydFC4pc3p
ZH5tkCmT3qrcnT0P4y7hiumscJe2RuwtjZ7wuegqoGGOFu6+iHuals1hmLnU+0NIlzGZmuYzRUPI
2MXsowsJ0KbtPwELBlJ9vN5upExK0Zul5SuNi3Fk+nnqPJE/LK6XhnsE/UTRORIeLu/QZvwX8sz3
kWl4AdoADmJJpmItFmcJgaCNV0+wEnaJoPkrGjFF7ufgZg8gSnbLatH8Oi9bJXeRgOkgFXSAtFvk
Z+OVxYJ0xhpQc0RnwQG4AA1iFJ5hANLfI4s9tWubR5e3xMXroyCBKezCe6nAXCMgVVPEdwCVrrix
t+43g6pgO8rBN0p6nfAxLq6beC9oTDnGRYZyASdAGZOZqjEfBezjuFAwgRRQukZm6ikYcYbliJw4
4huDNOkSzM7Q8Cwiz+RxpAmUgXzOb9LDD7IuEoUwJgoGapmusrktk6einNX/nLsIvUMQnnXwfsLT
Tj+8Egf0hvyyyqn8K1vf1FwMgpHN6+2eblCgjjiHOgKAK+rGVJanabNe0xZTuB13EQgniD4QuXac
NIsvWw13T8sJbpXpyVHjx/mKXi/ztesrpq7JTaUS+JVhQktTOMVE8zMnIpMn3bhH1kO0sbL0mkZb
wR5Vi5jDmaNk7sZ3bDHUPdkJYGtArhSMj1VtSqPAB01Z+33fjkKxBsrT0BGl8JYhcg0XDx30Ln4q
7czgjditkFvTD5akl3h1UxOEg5u0D0A92cRRsf7DGN0zoDMlzE5Np8ln8k+/Ar4v0pSD3hwpMFYB
78mU9xCLM1SjLTYx2VvfMlpfDfluGNFKYMlxSF2Q1Xa5gPv48D9dw/xuEMkD0N92YpfcH/tMlYv8
6jqJxRJZQK4MW262k2EVY3fu6IOZzRUxGBGQKdSzH3uQ488wgCksRiRkNfcQ9ruK0/kLi/GDc4d3
01FCYl6GK3q/oJYutqEB5HmL6Yt258fOJ3D4GoaeJQSHkPGFS9z7LJRXpUgw7pDBAbf2l/pSuFiQ
geS2ObhaSx+F0ak89ILChEIBGBwdtLe0RWECBlhBBl35AEG2B+SEL1UJNIy4PIYEHcexbCl2FtVm
of23/5YRKAvpJ3oZ341t617eei6LADeO6wM+vYNIryWJsACwV0ooR876RRwgMrS4U94rCiE9omLS
OEfF6UPYa047/SxMxsn3hXnAJ74YHuj4wxzL/x57P8uuRDY8nYUTlQVDXmJCl/AWQRac+V5LRdt6
sNb2IB9XR4ONHL3Yi9uRaGWFWew/Bo4zry7SDMRlq14bcjLjgQN/gnjHioJ6hw0sjD/sn8nG4VAH
bF+tKbF2E65YSDzgDCBSS84vVd8ej9kfIsMmLr84tuz4KtuEkWHv+Z6pFbgLzrHsYFlkxqmXu7sK
q1YUvuhMr4erew4wU07VyjaZcIdwjr650TztjxQY/okjTxbeSB9VMdMgoSvXwQRfiCItj99M+ABQ
mq78doeGu7bcygOsUqrckBrMTnZJTUmWnUzSfD0fgC3NKTphCXTJ0heR/l+kSXXatZK0fLlwtrWE
XYXhsSyddmrLc2nTj8LbUNrno42vET5VHA6IWCiFlxcTEhnMH7tLSiDI9aPfeSSRQHbbFepv/hqE
Kc2grFdjrHe9k7Yho+MV2fonrBidufpGzjwg2AdCu+ahlOpG+zaZMmC2Nr9vHh3Qa93c8WzM0/N4
HWAKv/HTIkDUi5Jl0YTRFNOL1j5qG8vMBw/ft3lThFB9YaB/g/nFGQKDmtPmxXTsZynteIXot0Pz
7yww+gW7RCjLmLCedY5opcTLiSz8qxyAgACdHz1qx3xvUwUauyp5IrD1Ix7+J+DoK7iUX/oMddfp
hHygG3afvf+c0hEYgqUhuGdWs0heqUZq+XlbBDgv2+sRhTibUUsW0hLtdrX3rfddOIkodHreTRPN
BTVtHKOmv5bP5Ku7Rprh/ahKw6+zRUkjWgJZkMmmbcvI5tSLvZGsNA8vLSi8z3udyQBMOPQG/+rY
wjA5OHJLW2lbW0uMmbKBMHm8fVcHZaFphbWLL6ipMQfCG09CYU1ClT5RC9Vs5r4vZF5EaxbRxE4i
3gX4SoOPrcKIa3Uc2evtrvbvgdYRco7a657Bw4oVp3mgm8OisatW4AD0oakQHwLv+CshmD/lrOTg
IpQEEsK0LkN/mhp3darexSLQKs/BzEibgcO84k5CFKnItfAMiZdPNr4zANmkQJ2jPi6aFP4rz1FA
euztvPbqOCSxa+ahF3w9S+Kre4KkLr0UzzFafstA+8KuBAojARfWGZ37Wmns841BRC/5tHC60BEN
OouPP1uXUYRjdo7oRJ9CBnKFp39tMvKxAnBMcCnJNprULHFxIBXLbUyewawr2OhuIomF+2BF4K8x
zZ3zDE4N48+UviClyLyknM9yQJtB4ZTeHdtqKFiE7VC40Y/aTD2E3dB4DyKdFtGaqRbG3NdjNrHv
hvC29j6id6Z7bHT1qFdcZfP7XV7B5uHIhLKrXAXTuBleFPQm4BIDSKAVl61rtvfS7giNixyUKnUQ
TSEIUUOswSgoURiWNaaVLln0I/5zya3m+vjqLEIWcniDvQi5LpfdgHh0563dl5I+7B5HPY7QH/EV
8ayPunknjF1O2TEi+7GPMw5hRAwZfdC9NTkROvDih8z91cRJX72jRfYaRAbM8Q5Ekp6i93UHpxhG
8atrfTbEnvtlEHuaWsKK54GDu+UIz6zUtaMrvJK1eAxdE5QLc2UE8HRAvqR8hoAepnsdsOaMobSj
k/NQqIahjjjcmCSiWxQ3ECU8FpfD+dsC9bPIZ9JODlK4t8pkg56Y52vhQCpCJWspYFCCbWp+y4RS
IJp/kHQQOWZ5qlBjp56kINI+QkJlyEWMsRYiDSmclMzT/S3HF+MRvUYoOoATfAG7tMBOfWX/0FMp
T23nT5w3935GctGIwkXoFeBROuaITnb5Qml8CGa4DytOye0Fo9UNkf0vL7aAYODr1fQdEbzeqRBt
/6S1vVXRrj+ChaTBAAN6S0w0c0+c8hpQU3lDxYOTgtQLmWvYFSvNoF6uew1mhTljVNbNos5bON2i
lKBafhYR7yCoBCD9ECgK/qE3nF/qxyzt5Mq3Z4lpbGjq9K1cphvxa61gliZ+GjW/cPfmVnJs1RwY
KPtNAWkuytEp64fgvv2t8SDIaknWJ3ef3bKo5gWzh9KsxA+hbzd7q7BLxhJqGguidxmpd9MciFoh
3T0zpS34RSkcGkK7AJA1LoQXPxIvNP8FXawy9fCPqJWtC+9zzunCI7kBoeA70ZUemDIRtqURk5TT
Bm8nipuHt18BAj7J81YnqBRBRBm/tH5X8+JNNW8TNrbQX9HGpx4kzj0otgTtmGGEWVIpaLbZHrtf
vNKsLlzFZU41D00D5KDeoK5QkXoHXQtrqy4Oaaz2GdkagcPD6c84GzScCCnHdPqi39cVwMu+9tNc
2rWkgZ8zsGvJpBz9LdWx1BIk+VaO6ipfY2Gp8bsQzyf9arG5XPq0hfRS/gAfWcyV1WRX1Uz3Xl/h
CwqOmam9vKElfzBDAbAFhG7T8X21qBZNMt+/YtfljI8BjvJT76iF1Mp6jzkRtc1MQkVDL65vTJbE
flJfen5JYj11cuIKjv+mrhHI5T7zga5HdLvVb52gILyxEiCk9eHoNAwwYn9NDMBEJ2wNeO6wLzv4
eiAe+0hy3sSd3dVZ38Zs3rSOBIMGt/SZvpV0tZuvdb9n6+sy60dFPdU8o+4GIWH4Oi3M7E15AjE6
sutdo+wwav397QqaX6N5cOnLPBA8NKOnIrFcYLvNvmhYpn/8vbXeEmzmFnsSLYKxmUZ3h+/549sx
FMcZsSYBZAOFfxJbR3OKqCz5nYHRUlGA2WWAU8V0ucsbiEQuL1TNwRM8CDbnNYcoOzWFk0b58gfP
D+OyEjVAFyAPZan/dcQdrEl+GO1Ev6xzEASXN6NsJDNm7bYU+gRiBU9/rTSpay42R24jNgC3v7Id
jxDG8Bkta1PObnUKviPAr/RdapSEpRElXr4KbBFWM2yKXoazvKoePAzXjV/k1QyO8xw43BG0f891
qZQfoilQqzNzXjD1nbhZGsoRTWoyuT/bSGynGYwE3x+YPGn7+1CAdpV63kvYS7PNs/tq79gru2KC
6NEHtAsw5A35GlK2zYP0rLOhsVa+CtjEuMhzPSs3xzhb1Agliw7mQEiuJ1huxPZny9dz9GQItA8u
exSzOVp7IfaeenrU2bwy7+BpzpdA9YwHO5MKLq/4D4yi14/0rcc/tqEmppgk0ybRdaoVrJZD223V
wRi3SpX47yX67T6s+4Ve1vUazwf7G9mTMxNblq0FApH4910OqKqfmN6uD0IE0FB8dC0ttNYLDqDL
+Cg4qyN4Aluz+9Nl0AE9l913UR4oZmMePM0kSKr3ajI6UKX/x50lCa8YPiolbtwextDmUgLcpVYu
u1IJ739gTH0JTKjhaRvSbqvzwR6tVNM+p5ph89QOPcOUSO3u+7vLFtspUju/OA6TVPWH2dAL/Ded
7Hre4KlxMcDQzKOBrDZOWFipaVCyJr7moEJb3pHa7V6gOZNGK6zCitxVW9UPTlLaoHB6pJJzNcyU
xDbNB9SsYA1k7Q2Mw9PCQSlKsL6hnHma+os6C9zsgnqSChN1l3nL5tAsFimBiyc/4gKpSEuVxXl6
YMemvuLHQgDNCAFDWnZeVz1ttXHDzdHG6R8PYpxo0CJCEvkPIMz8aDRPVG7qIOgUvx65NqFBamno
QzLTF2vrmUlrHXeincItYyC+0/0n+9U0sBWozhGhsIEwjKrX3VVZY63I2FXxOV2mMObc1GKtMZeM
YQ3YpdIPtYGloTuk/oMXh8VBTkWYmgorrkLfyQuDGXzqSgqS55RaP8NYCtiMeGPrri7/buTz+i8x
KRPGIah7s559DINqM0qt6ALAYNaBrqoMbI4bFmwA79fw7z/UNPZcvs/6yFj7uJmsbt3/ED+vAM8Q
zYg1f5YlUgzSNe4tIqOriNLb4b/gwle50DZDwMvhf/xaaMNLDhEnHW8G486gR3DXnoUqjPqCYz7L
zdii8M6/wEXVetHhWP1taX+hxQbIsND4LsDU8QrMu2PCr2jKfOLgtY1PjuZvk0Us0bTFWbDqD5+2
FYcMxNzw1zFnqpicNVexKSxwO3iNO3GiyJ0lDPSaivqC4pbHMGyZHcFe8JY3AKFNyRaa3qukKCdC
/QCaehsqrk2VH0LwTUfK8OV+vYRyhj0qNPqc7KQl8Ci2lay89IdoMqnX6/GqWson5nTXXsWfA1oS
qPifmDz13xm8c7HePtX7ryyQVAK5FIaT9QywHho8B1TEGRd1MRTtQLL7YSe27SYoZ512d83EqBo3
qmHNANktO89xwfa4SpUs+Lc3rmmwTevTmxsDdwerCvnr2bWOUZL3nhxfQql9US980Srr+Edvu6qK
aJzEuP5gSAqERWal0Yt/deKJ2A91w9vSBGTbLx0N4pdqVjDXfgUdInT9qdZZ50JStRchFJeb7g15
BIZ/kvw3RKmjYpvtOfXkGU/iNELu+AXV0+3welGVAs2vZItU+uWPlwhnQMkXcl6PnfIyHMxJR4/f
rOiaJXSwwGkamLMuOxYQwt5vLBAfNnBhSL+85roYfumrc29iqZZ79nNjX+R5ft7S1m/8OOaeZZss
A7TpSAZhyFrcZsfccIpjbhY/RT//epqjFog0KFLCirHQ+Irr7TUVCzejZ9ECkE62ipALeGqoFYGY
LuF992a5t9wtL6uOrT8wBJKg0Zv0o8xxBuR2rXr/6ewDs4VHuyucjKBRNxHzInmADOVaR0DSipbu
bEUNGAhxNTYSZDC+2AetuX54DBZ9bBf7fNN807gUC7c9itGaCvE0YsVgPzaUbnwOp07wBJF4QeJv
YQIbRaTXFjewoHYpz+pmVGfaqFvKLZJ4IdL7XTBIFQRxjwtB/Cjy5UcnrR0owJBXGo5I5O9YaiBk
W4rxryVnBgL936ofaNZzJ02ryw1uLvsnMv1bTDwc2KbMUoMD5cVXrM/DBsrQ61tCXgtFJU0shgyQ
CuQ2e1qOdjQ4QEgXVv+kpd/8ekRlr/rp2QfsqfM84t54zFZgGhAK12LL+TQEb4h8P5EPE/MiM/Jl
NGVVG+zdX0ihQ+GLrWMqL1lyu7DlVgW01exL7ROADU3QkxqBMy/iFF/sGOwu8kbMRX6jojgE3ZxA
d9RtSQ3CvuKMR8RcSfhBpRxBvvSIGeDyABKODc84e00hzmTCjfbhTY80AW4DEu3jJmm5KbZLTFRF
SteDlag1To45QphSvugnZ7YdsZYmiJrtgIQ+l1n0ALiVEv2Y12rssCJEglx4eaHMZStyGlHZeRHd
NsxKhiHK8tdfYpY3LQMKiFuasyApj2kdEmPJeZVxZXKeA7Zt0rV0mrTwCvaLlgJWT1RH1xWem4WP
6lDiSk3lqXcK9jwjpVWNDut3nmcrUnaMjJziaary90JnyM/wzNr1XEP+1ukCXnEJaCwQDHbB575p
aWS2d2PcgxqNnfbQpL736mb8sIXp2LhhjqPB1re20AcZia5ErQ3US3PEBrdzIfK7B2y3NyUh8vk1
5ruv6vYW02SqwSuyEPjD36590qRzRS6ZjPykZmRRHryMPNmH4u0WcL+LFJ/9EGSKC41NkLEKp/lI
sICnRTaBiWhSoJsFDFX6jp4QNPK9SNbRqngx2cSvWBFN9bsYaUi+Fer8vIS4OrFvbu7qw75ZZpvN
MCaiw6pNDmgSEnKrh9hMOBykWrxcSlg/vouVE/SaW/r45RoO9r6WOLnNEeUMKAoLqvuceTcOIOty
znHkLKHZ0h1F/duKZD1EJz5pUJUg1NSxCYoyVv0PWNFS8XAiRDbYXMKLQ5VdHP8Wx0wq8fz33uHh
63fcVwluAAt3D34uRyJJzaeACOBCQWQTUaIi7hLe/2vNXjtz5evA/Q1M6fXNYbQtoJ5lp9XR0LGW
WkkBCOD+wdM3i8Gv+4q80umdtcM+fJnd+RPpRmi8ynF7VTQ0ubirSnVKO6bqYrgpUcXvMfXWbSlz
2Dr0hfSsFEjbq+ET7aEKq/JP+43rSOFIlSyADEBPdLOfvO28yexTTzV7nBKlLAsX7zQNoKd19UyD
y5RK4oUDbwESS1xvNb0/7bdkJuHGmhGf7/lQKrChtMrpMNkLH9qazVM3w/EEptnI1FFIBGmv6XFi
cWqbl43t/Lx2SvPO8WIdKVkQktWqkY4ckgh3k18IwclwNFzce9Js+JXwOW4oivAk/XcEnS55E60/
6Z/iZNQJSnKWtNBMUfkpKX8jsCLy9pQGC9A7wxgckAT2awipQK6R4kOtsOJKCM04e+aMaD8U8Cb6
gTyfluwQNu9I2taRmDETIrHQ2AISbxcJJxF4d5QV9cuREhJtRT4dRZlcqdKZi09lSzcDTW9sHoVg
83QgJ8PCH2uGwlpdC9q9dz7FHrJVUorVZBIAI1mvWdDOhu5D1J3k4w+W/A+Ya9I2OXQi5RmbkX67
8OV81/WKo+NoXNPFhKeH/+4gv3oAVFXveOsavtYYA0br8qjluGajZY+59MMFKMGyecqXsTLJw9k/
iARnebAoJbG42STdvy7LWn7zxJtY8ia/MolVneEEmm5uC3+hOmUjeisaEnCeXT3F6wKO06k0UAY0
j/7SOVdUk1SpbcmxYh91DQ/Zn8Iaex/UOmIo7zUSkznQ8Ol0z3pVeJAVV3BvkfePRM3SKQsdQrZ/
zsAT0mD8dPY552jd3Vyg6namwtH1ZLUxv4swyH63mBireiqMxXbSlbak9kFuhbILLO1ypTQpSuxQ
d56jwMaG1GYNBNijaUxYmpeuiIdbdme0s0nmIMkjL1A8cWVTDnCVme474DwoNj/2O+JkTRUZbkCf
dfWO/ugbjC5lSgptyYGW/qRK3ozy0dBodg9+y7NpOJaHZ+6u+JslN7ulC1EZdELI164QIFg4yPAv
7kKw4DdryhgH1NitrU4EDYh/h1zQ6sYA5Ua9/9NNO1my6f7ykGUwsBO8iPMKvaDx9fqX0IFdTrAH
+l4Jzjvh9jG9N9cMHDuRAljPNxWjhHj9euBBKZWufaHyQ74U0HhjU+GeYxJm592Dxg6QZiUnA3V/
+nHvtIyGBsDmAUN4bLiT2l0ATpEvzG7hIz1lNLXzr043ifCIv1g0ntwD8kbOrq9Xea9pxxO6mzlR
+g8/xOm/P2eeXzikD3j125oBsvNaGzxFKgd9AZ4caYlPlkEpCB0UrwPr1GI06CJhXjQ56ghsK5o/
bpthaP290GfY7rYl7M2BocW49GoUcSH3oEaDUYZuxFfbFAKgFBKeCTfIbxhus2oXAvbtRjORZqzC
1g5cN5PK5yhaZbpqwcVQWF0cSgRbMyH0dE2mn6N7YO9VOV7gcgUadtgS7Er8o/C+rdtTO+HLk5gN
TSagCWUwnuIh3UjFvWL24HTcs5eWfKNJU6pta0eM2h2oLV4nC51JK1f/6STcjBTuWScOfzqWp4G/
bovrkrU9YuxV96NGhOZO0zC/ZRfA0amL4WOaLfuJWeDvtsuODds/8w9ZvzTFNhQoJmDwqBKVDrCF
LjdwJoZjYG70eDrqFQ1UidH+3Iy+8qMYf4FjWLXjoGr4VwKWR9rFEnRP8APmJd/R4tcAF6bHwU3X
B8yrSdkpaxjoyZ7lgHEfi2jNQ8j+r77fS8HDXerqELGypUVrAllU4Bp6Q+TQ/KeSm2FuHusgSCqr
hYfW5YFaXQW5+Veytn+K6v+OuI9DjEhm9AtqRt1ZDP20gnqcgXexVPHOSLEXjIlNlX0LdgIKXsWf
vFZIsdAjcvWceXwtoe6WAKRi6I2hAqUiGZcUb1U9lTTChw4AvKyjy4LDhRR/Tt2deN1zZwyaDrHw
0b41kBnaK2GghgM3ltA1ZenHvor070QzKp9llYRhW75ODYqO4fzl+AfAITwz3R6zB6c59eljppYA
6f4Ncz5xy7F64ciAYIHkKitXfBQVccX735DGZAOEiu+h0j6xlryNC7x+KflH7kGCMktoRqg2uWv2
mezHKGhH82BxGAtr/12gErQ2rgOWoQfch+oCu3kT2ILvHslMJwbZ0V7OdgRoVSiuI3SI5NPnUDP/
z0pyZw7dK6vDzCjQ4li2ToJWRoKns+G0wi06A27o49MoUCR3qr2CoCTyUYubalLZSDXBFQBQ8u4Z
pQZtU1HnLaR0cbf9eCkcHOgF40C8i5jGE/8XS7qe5vBjIcu3v4i65KCM6ARf53FIXCU42oRRlDAM
gW41OhTLc0LgHIDUI40TdPNq/IROxAlufiKMVkxmLmpIP50UbjaLYKrbWBvkfH614iVQm6aILPsY
xgPD4uI11ZXBeGpp9aWZ+tlSumau13bC5GmoalJ1HG4zYLSeBKwwLHWNBhFDMEiPHBwpeTfBZoU4
CrLqEXSnqBJCXdLvYeSPDOO94Lnp4YST5vzus4W8ph2C2Z3nARv2Azy2HpfLTFEssg0+lHkwiEaG
SvntLbsb7HIQYI8hh3UcNzo4XqIFcdE5IfKRK/1CjRnAOk3MXs9HI1gbEA+TiJqZMPSogh3sKeKO
qM3sP4chwi68etY7agpt2z0D+WroBZdzkFAemKgu24zzLRpsKUhNB403PcpNZc5DDZFzQROA2BE1
DYCIXmVXewxKtKm7eiTwgoxg+mDXyNpf4/j1W8MxVTZ9hDlTwf43Lf7vi/cC788jRNRD46t9oj/K
ERLABczW8VM13dajJOD3Xetux23uCpOP+JyuzE+qTH6EhhIPSCFQkVbFXb4VyXSyWoGP1V/Igxqa
fXARBOkUSrRe0VUHKD6OoYPUcEyCsMXhF7sxstCaesNbhz+sG9gkdkaI2tZ1fpAbF6YUH6knkiTA
qbnCub0ZRLFapx8O4l6ncEjTCX8yN7AkddWJEUIqqxI5jF+N++3bOvVaVdowJSV9kKf8NoqFBYmM
bQ3wwh5dbD/Bn7LijB7WdFzVEoBIeqLmBYsMcK+ur4mtaX0WG7sGMOel5RsunDLpKKgaGvAtM4kX
V2ctm8rL06ALzrtWO600roI0bg5/Ggc/CPNHFgBt4hSPtpaV6EmQRX1G+UaZk2g10cQ334MIULc/
zKJWm8H+8+xhmrZNN8OAIZPhgk/X8HfoFxyPxoUVzowMjwiYV5Ime1bNjXP5sOYVgGp6xJ551oLp
USprMP/0j3tutLx5b3jAHk2eZF7alS0so7gErPDFxz2tiTozvaKv/S4pRj9DAEbP+tMapsrHPtj5
yE3xW4MlM0A+/qb503vlM5tXOQFzyb9PJzt/wsykI+qjvU6Odvgj0BR37BnPkbvNzUXiLB69QSKM
urv1ar8DQEi35qeeqaAhTQvAaJlVOUsuIjwMuVN0YYrS/njbsBEgR4EyjGqWvsG5B1nEfAOu1ZG4
BwnCtJrFxBq+ytZqlMaod6E9N0BZLOEKJCeInmkFnoQrs4if4qhbeYXGFr/N7f5Qx3cMLkud5h0B
Gh83PH7XxIeZt235FKbiCnrl1LN/+HsaQ1jeXED0xmjb2XFLf5Q4+5tMjx4bFLwNRATfYPVo98+I
8TfSdsDVLeLPkoGe1OXm6NOiUUu0Tw83eQmnxnZqSYj4egx7U6MRDXiSt4C7/i8mM6LlrBLJuWNo
b3/DGJgSj05x35t1F6Y7Z2sJMcx75W6U2vFQj4LH3iz6BXpIj6X/E7mO67DZAwo2AiZmT8r6PEAd
5HLJIuDGY7mgj6a2P2Nnl3vXRtRxWZAX/cJEAZAwIEyQOrm4iqVivX4MF0fOwQEi4wuKUrEJ9JhB
kEicFsw0+7VaPVCpzfNadfxcMcmful26xy/2rTmoW50ZVaajKjM1vwMXHVbkxviSKGwTPskJE4IW
WaN5Og6pC2Od17FBv3HzPjCRa24560tDo2nVYP8GigwDbpfXBWspoAkwjyNHrHqAT34F4AXOiKzL
k1JQ6jF/QbpmI09dge3VLNrYEu3VINXgU4wOie/c0pNDPS0C+GD0HRD4dcO1R69q57yzLTJzVjfL
sfl86x/HPV6U7RxEy1yKjec95rUC3xqIut9JGmJzo9IoZf4v47QphILDV9rA5vNmDl0IllrP36ZE
Vd/yqeIVZtlJ0Vd7yEotK+tlUvrG6b0VPTy3wtjewsnWRG5qdkr+Ppwm5Q71ArfJfCGN7L6EV28V
nue2+2korZo0hvrcM48mk6zooao/kUg2IKsJkoYnf4f5+zcWjlGd+UH8FZWzQ8/+cziMoGrNUwLa
EEt+3AJMVBAra278+Sq+Uy9GSOdtqfkjvjyRvNChfnl3kyWZETaYKsNO5yPX+POf8J+bzfwLb0FX
J8xksT1HzdoSOukcYX16THdgtjJA6k+Qkl7Gk/arg4/GYk2e8EiNJO38ILEJn2rp25iJh1LddsoI
SeEn5q/jxByh3D5afIxcnQLtZpxpY0FnCCzoQNypVBI/9FMLZzOPtky+8nvS+B30uut/4P2BIXSY
rN2ZpvY9IdPbaPrwY7uml0FUuv/+mcdnUqKQ+xRBqi8zOv8hQpM7IGjJHoMfB+tVs8fxL3fNCbie
C6dxapqvV9CuyQ6I+rrGsWxJgJtfFbw8U+mfavEZLUUHL0JHZ+IQVOKFFy/kjQcK+/XfElg0N1OT
FgSlq95Ml79H7rHoALG0pugVH94ZlmjtskHbGc8BwnToFzyZ4KTKDzHivr3MZw3p4Py2tzYPdO/5
gVsi617XCcm1LwbN1NjgNCSXuFZ+HtT68uhFQJ7jMn2lIxmF3z9r9yKF8ILmI7tqC/EAbYi88Bcp
mR0aV/Q+V0u7Z/KDR0z5iUG7WRumr87JytxeIWYjLiCiIaSGcgqAXYw8MDHI9fF4ZdW+GBUQdiwK
sukQasZF5GyvKLG85noRvNrYFs35V3wu8Qi1WR2lNAD3rRBjSMtXPmzVmBImwoI8P0qs8C81fNk9
gTl7ja/ArNDWZPPEkHnGRnZlG+rcTIhXvEcl+rVR+gDFoHg/7V8HI03x+Qd+SGuflP4iuLnmTDJH
lou7U4+Vkc6+v+qNaw3NsOA1dwlV7azxhsTYelC0Eg4jfHUYLPgqzezhSFK4NsV+w1lVB4Si4wD1
pZwV2YeUQY9pRa701Mar9lpsqtn1kRTn6zSUvPD01dHHG3haoqEOEfYxQbnn76g8xRvGEE9hNriH
8wDtWSZnvyVh3JNzltH1DKuXnPdsk48i+RqYNs9rvsM7ttSqgEgz/coBS6642eosnVf/HuNmkEFk
W4T28Zjw0aHlylZieskSGwGrNTHueSEKSqkwAHjXlS/7L5DE8NmRYqTTQZ3KepyXNYBenKNazL6P
6ov4sGXdsp6+boxmnLlltdrns7qQtsJ/3uF74kAUeWhtJuFUEMAsxfR0OQh0FjVSEmZ/engCMdVA
Ih6OonsK2GJ4MjHp6lQP5Pge5831Cn5XgvdiWsl3KJNLwdqGKgcxF2ebQ+WUGE+2Wb1SS5Gwk882
eUv8Cuw2w9s0J6bMolEs0LnBFBE39ORiXm6Rao7D7MbcAA6Qz7Xs/bcQxO26IhmrWRvXnSRdl1uH
4fdf4t2U1xI215afDkrD9zlyb63hZrdl6viCMFzh2NLHaJXPcyTlfNRFXz2oyZEOeTdTGoPY2MAt
12zVf83wXvNfTLm8Jf1FOmEjWiEIR18mH6xqz8rgNC8B/VYFzIccqCJfdpse53ZcAblYV5JRclQb
1TeumBsBB7ZfCHu5i5BdrgNvfISTGWPI6kVqg62Bfh6bmGP97ZmyDnDLAqkQVxGo3YWblTYLMXNi
w+lmvrgItNVp01IthxanH31al5nZoeMDocOVZ2UCSYwb86eyTNsJsExDQi7jy1tZWCHRuNDDVNIx
cy37Cn9InUYyVvBibYhzrsZrlKQ8n6J97Uva8bhbusMb5gBkZMiUqQ+az4IXvcZYDA6JWGIXGdXp
AofyqXgsoofC362K3oulB397CX9+WogdXTPpv+mNr1Wos2+WADsqs7cUfIk9sLRdy42XHYmPjaCy
YvAedevvf0oPcgirU6u8p9DFDvsE/SReYTP+1DXHgUC6NtUQ/BUuBz3M9nYyVoZa3Hl0+veWixH+
MYHV9VxOpy8rhwlGGXGfaOQ4y5lrZBiBoH5Mjl+vB+GuC8GTN3Xmd5kvunmPEhk2ULskVl2GQpqK
EOu8lhp+NJM7YepvsrMWq/LbCO+TKTxDa1s3T0QAl39iqYPNv4sCt/5WW3HHyCLpR+AWVThc2kAg
ynzvgdzZa+RaXF0MN2NloiX7DTwY0Fb91b76I8PzDpxPJYcnlOfxKouZeT5phyAYN+TnWDObAyDs
EM8lGObZ2+IFleF+YKUJssx3VHf1eJa0zIb08jnubMSnNBvUeeBi/hN/wVFu9yimO59uDjaV/Hy1
VLbFkQ3t9UpHrnCdci5gg745N+QEa4M5j4qhoIT13pqVlRUtSQFrobsk1vehCiNzw7o57FLypWG9
F9Kn22xucbvTDkBysA0Tc2dbbcgYp3E3fDz8zWS5JPE6NsuwF2oYUpWw/STiGWaQgFYRzmC6Nr92
Kz6qmUNvks1F4W1B0jSxo9mRqQZVQA6IRG3vZbwFr3cAWg+iUEpVRHuhNUg1f1hDZwvg/qEyfY4z
BrFWO2WvfcRxRvCIDzrSxW1f+jKNfKaic+QbLlUroIHe9BS/MRrCed9scsMc1xL5AgfLhaUBZc7Q
EPbm10T6xFV/LltOv2iCyPDeGGoD6wraH/dr8xuzNGbz8Tg4PrM6MzQcefe+lh0mvyMzfM8PtKdq
eVQvhI69ab65+Z/JG2rrn1qK0LHnqPbAw1FVLw+9zgZ6aofVBj96WQ70byhBjRgJ/ab7Idz0LA33
vQJTon6iuMLR7kw6PdwiKA/UmngIY8XkyE2xrfjRHU2hlm6/Bj83bYK3s6RGyLW4OWKZDfmGO0Yl
cPSGyNXJqiTUDWsPWp+YVyk+Hr1xylSucTV+JEu/JYdWjgHgq+xJ8je/n9f3zHGAbMmfDkOZxr85
2yeZ2fXPh6Xe5WReMNu6WIzzLe4ytVTiBJAQovmnzeECKMHp1/sL0yOI41LzFTkZoa79NAX1G7fx
JFXvni3dxI74+MN8SFbD4Xfuz/El7t+977M466CEuyOKB4JOGMEWbA9dkSS3VyxLRnwtZQcRlXi7
6zoYUyiaSwelRQK6un+6l27SvblufQla03D2WH3y6jyQrrb5r/WMkSCofY7AlMx8GcYQNAGN13RQ
XemGl45QUsQes/kXZxjodii3qm7Gzf7b5AvCEHTsJK9nsTvUf2h+pdBEKMiEurQoeDpRc3/jy1W5
EJEGGTUkUW9LA/B3T8tJCLlHZANeYXFTyHIdPPiZps7kK1GZA8C3tZR0lHUIuKzUJvP+nRizNgh2
RQ8jlopxI4MUaCH+gzCxqRa/GGKYgNaOsYR1q/FlTiLeiy+YTQ6zyaG2P9jPvGqdCx0+gxv1Mq+W
eg6BWNg9a3VGXpzS1n5eCP+Xf+h/vbRymqw3pq316/kNYTgSaOI7ATCefPgzgCgZqzvcFjs4wDc8
vfZGIKYXntoBzKaYxcGglmryf2NwqWvW/DFNUqletY7iAUTMsYCDFnoAKZE5D3zTL+3N0Myge2lD
CuVsa7jgIHlk+YA8zIY643maT6KXS25TE1n/2FmpUkAx4Ya2g0ifkke31aNKuyuuk1Q/xiyeKO1o
WRW4vC04NfJMxyUEfkadH7fMdoDW20QgCJXxPiiugXiLJd5SwlXuQu/6/N2vvTPw9oQpGurAfpTE
jbxc//wGcKcyvmh9EPP5tiGNNx6agDKArK0y3HZLT9KTsodsAcva5XwK7eeLwznhfC34ONNsvPCG
yHfENELXdyVgtMUSFYzZvp+EbZo9IEfKSX+X6nD/U1YVdvDpZiBEHPkDVGjJUF1sPnH+o/t86h/U
lChF0O/ncmdT3q5u0Sr1ucBSOuVlaMLfIRMOwQoXv9FhHmX5joD0Xy2umscnW4htcxM5z3tC5IKS
S+Cse3NTXkNt6u7tUtHFYHHBwuVqHcgAjuCaPEg+XdDWrYH9Aeh8E/BgzkN8kHnvDvjU64NVqwkO
LJQvlCSOWHBvTpGHveY/HSje4ZUEVdUrK0IYFb0lagatZgxInxPKdNheqxih7+eda3MAQ1J5oEnS
FAT1LrBx9w82TjWZylYqOgTKrh3BUof3uzsIddnjyFMSsA3sAMC6MKshg/cItdKnGAcLL5Sos6fQ
oLM5iMcMCuVERXAraUTdvywGsPy+zrgFgufFmcUgEdw9bS7KpraqbKspj49DXxJFU9M682414+Rr
I2BImILAxfZIxOPAlv6cNBcXyrEYF71cUXJORh1knt34jJPVHu4WJHYReURFtz17uYWZyXLFChYv
MFvHEiP7HstCytrlLzS8SbZ5B/5YcoYdkWAUU9VftJ0taHMHwFs0PwTTYl4fyfsZs3KIk09Wbx6H
P8hCmO1OednaSPvfTagU6OdUaPvMV7K+37JVzg6zUTQqRtNF14FlV3thiA5Sjpxq70BV9NICfxaP
GSDf1OjeOkbRfZgXQamtUSuTvsulkFi+W4sI74FflEztWf/nk075qSLXpoeXKRXanSTtJMWsszIx
HRZpFmZnOO6YSoDzFQzZkwDTToUO5m5KVDJL2zLNJsSoeomd/zCfUAuRO2VQqzU3QEAs9qj4gfVJ
AAu9Oz47rykBE8+Yat03fAb82BQforHDX18c5MwM+pqcj+ucV2feytThlVB/DqW8jQXFIC6/NLZO
4+ewTYr9cuyrx7lFZBSFInR0PBuIbKguKshKQ5KDsR7unloaUS5WHCIX/kfHxK/IqliNV5B5z7hv
jQpZQGRop7azZN+fYBT8y8k0TJ2ZHNXXw5peN6uj4TYDPTZ3TMXelx+e5HXAYD3ExlWf+/Pfcijh
ZstyyozBWQ4Js6aYtxETW+ikA+uYD8ZbKG/I3VWb9S7KtLXaWXGs/8M7kkQKxn4gQKdZHBQoREOT
+Rxe/U70K+MxSgn/9RYlfPkISP3A1fYRATwes9YycAaItsBruZyMeuDZK79b1pYU8dH8FLhpWr2K
UkBQzxH6wkn24tHYpH6/h4msSrFpgrTz+QEeqhlIPUtcHsE82YHC6i8gy69q425C+zOvvxz4XXoM
xwNWB0GVtQQV2XoCBkHqQQmo0ry62cCU8R6Zh40gw/zFZNun2n+qUPig7WX4jMP2CjvoXSkTDGI3
OP/69yIWZsA7em0ZSiI30H/25roRE4qPvO3LWX1gkV1HepSqc0gshd7aJl5n/ORpOyb30H8lML7T
p2FvYKr+V6GnyPLNug6ANLYiR5N7whJQ0XAoHk9Uxcu//Y9gNWz7FgkRYbp8HlXwetE12Dp4QzF1
1noKljNUDo5ELtMOf/2tbTlthFNK+77QDIiVHnUbMAZk0mAJaE8A1UpLeTOSe3RiJu0p1CTrTTuf
rnrPjPHQKwDa7iB6QeMjZIsAwx7LYCQeUNHm8AOH7BMGrIfm7fFR11gYIoqCOYh5ZFSqiN1NpHdE
Wu42fgpZQDNsVmoiaM1jTiYWrbi1vjcb6S44mTyTQ/lg5bfUtiwckNLIwi5BcYjv+VfHsTUpTH+z
MhlyjrHgUDrgvEHsrJD/Z3QY3pBOKauIB+Goin45NLDuZT+Uva+Yk24TrYX+jxq24IMw4ZQHD6Gn
XGQRxq2W7BNiB+EER6lNwN+96gW8Sht4ikbIoIdLYy4g/BPfUBaKJkiiCZusIfysUFONZZdYSVqV
dpUkDSVcRdVRLgEUNLBbzepO+sgcrzgb+i/qA0QeYXf4IA99CU1MbiqE23VH5qKGK/IMf+RVqNv8
d9NK67Iw0jWE6yWWCvpCUYUnFRp1QWR4f1rpZ2L5hYy93qyJqEcL6pfRdnb9LlxHBUO2u7/uD2RZ
B736MJp74DxHW5nvXGF2nPupkba3T4nMm4YlxO6QSqmPT8jGlFy/IudJUR0y51jPKOosBdQc1DOv
PGLv8yyLNaRsFUjnmFY8zC/ms91omTxX2PCV//9vn1VoNFAg3z7tJ10OpxmLwqhoZRwyaiQUyFLf
Z4dBiLRgILftdFHTi8pjPeCGR+6HeK0Kqk5l032jk4G/jJXyO0/oLr2RwRukn/L8YGvI/MlNnT1J
97kC/Qr5A6M5nJQDOavouhwPQdgt0f2wltYt69HbkSKa70YU9gOQRLzE93AHdRaCYtH4qcqghYx4
83yULGnZqXDTI4KOvXw2rUwtqiEAMwXgFWzqHCDtAK+UWIxj7JIcUeK6vO7oy1/ADT9vCs/7rC/U
Szt7vs1Gdpxoh0ow02kpj3v/zJKs06pNxSmec6S54ErFlhxT1xPmwJHRl/L7nlbplR2aT/qQA6u0
eQPAPx4qbyiwEF5k5KNyzKw7nOX+zOCGdgAYlkg18zunR2i1nyQIylA8TW8wLiCYD0cKl4U/KFTf
OwqrTuxiftqvn0vjDs8Xv4ayaVb9k1i9Eq4sfYSM9n8QuSNlmgF1cm7cX9SfU0LLKiusXTkUWEiP
nKmOm5lEd35BEYWGPiPtI1RFHzxGgcosslM12ysK/fs/PycAQr3lS11A6OhuWvwk76uk1CYe+04F
ZglH3oNtRBb/c1NdV0ydEL339+NV8v1lEwOZjCPeN2g81ZyDKtdgBA16L71FoSnX7ZbykFehm/hS
kY5Xn6c4a/FnaGayZGMhRDJvI69R4yOdyHTu58/FacHmcEL0bSRTRd7ZCKGx3Oa9nHKEdg1h1K6J
uT27wxi+fNf1enpjy+W9z8rULWTbS4BWrvCcE9fcJyj0THX1PnOl4erHaWW70Euf+cOhcUgTcCcH
bnqUW3K3rYqJEf9BPijF4SMPcFqnatr72uYzC1PpT8l0WzC6MierEX7aQbNmH43/Zh1a5zkXo+Tn
zqdGx9sKYjflWCJaK6WwUO239JLr+tylRkB2XC90tbdS1gXB40GUQi4mnwWhxrGQ17yte9kdyPnv
lZ8Vx/lW55gpacNSMaJgBMnhZlWEQc3BfxJ9zGLLEUNuSeomm/BfjG2MLJwNqntflHnMB5Xu/Do7
hwaG5VYluI1jpoisJtAVJFXFqMi5A10tjb0Q6AVmBoimGrrlYFQLDghWMGSoTJeJiyTLe1RYJ26w
8szzvaMVdN5mPBxbd+2Ykr4NsFUsbk+9TMcbBIKCwbRqVgE5Khwpyc4gIyUczZAAljo+bwvpW+gi
XtZfMXa+Lsx0ZBQnc7pm35+CI61g3PzR+8TaEqf1dEmMk11vFIgL2Y+hbFhcCTT8zXoQtHFuaOrZ
1cabqoKzAIQjMKkxaLmG+jXv92DQVZaMImFYftlxlR++rWrJrWC1KbSYMFhl8lKRjsrPWRo6z+au
MYFfwm8EsmOK0e4WEm0aSbNQDCEabsE3Prhsw2qtx4EKd+FkI+Q20CavNf9xm5co/gZPhsDOZDGX
OKITxjjw2UNJmWp+9Z8JtM+/pAdLglXvBx2q97aMHORmutK6y5lZw6kap9n5FlmjkhbCDnZZINNc
agzVqA6ILW1lsGVEfgKH9EeRIcinq7sW3TAiNM1OEcv1km54sn1Pyg8MV1TyWq2+2SJZ/ZOybSur
5XNOTaw6iePCRjGsqZ/znJUQj5IbhU41JhJTlM6wsF384l09Nsf8mWx25Pr8dn26fCKkuBGGnDx5
KXswo9DNdjv3JCR7nECuM5jXOGLG27pwSUaXsuKExfPqwzoGn5mXO7k2d4JjdDPpCtdwaKIoqNKe
4UWNlDEHnou7+fuz2w/OlzQ82N69jLu0m+lmRQsAIQ+9CrU97RsSaPekp4yUwXmkoIvZp6kLDOVj
/Am/Y/CWgwQEIyscc6sH/6qdNA7lnKa3oaSATO9kinvHHgZsYTggZZO4RepWwg/twQkwWRsW2h90
70VT5u2nUEcVle/xK+DmwcfPy0FWjn+5VX3/P/BfPvRp0FS0LiDrWsiuLzRm5guI5BX5BVtgc44x
oXbexRX41zRed1FGKB7GjKTWcFelXtDpUb2G0FA4HwhHpsGkb+dB846Gtdlu70guDkiDWk+zXQim
rH6QeaqyLqBpJixAcb1dGLy8sD//b8960wGI8kbK97vjUpW238AiMY8Uccl53LHQwELPB3bsfcRa
0DDy57AiM0t8bsG2+R0svCH4yVW7zk7o6xAfADYWr6gE+7FtWGgrnh2Bgrgew1kMLlkSinQMHQrL
7+K4grQf37FYtNk2hlez5wFoRFtheuORyS8S3sq6h9m1IAKRzQ+kS0IybT0Lul9tORMKRJhtkvCw
Y+dNZRLc5UCqrPZQISf1BN4PvRUHb+/H07l3cmMMANo6+5ADb0MPr3+JM7kFQt+xgjz/BhIBchtI
THtMK+harOt7hDDNUOolhfQ5XD7KVg9KEvPrqo0ggsFO8VuY2tLi9ZfzO1vUZ1ah2OmRYl9baPIA
zuUBbrGFuWV5tUAHFZ7tMW03WKCjSg69cF7Zmy3Lehj8lHPLaWA34CMoBBHNNJoWjfhd3zAOOJdH
i7qSJAStbg1t1CNIKSp78W92KzWtVAXJ9yDk33aUQZhMwUjsDJ10YL+zabaOBcw90K+eKAium20y
GYmoCZiLxA4Re31iTBrXGug5MNwuNVkApG/yr5Y4AVeG6nx6z9JIU4698r+ri2xI15lEWaQH3FN2
KMbsuFTmAKsFFGY26GBEx6Vgf2u2sKkoBxvLBd775yLefSGoDWjhGcSOcfJt9LkwxWXwCZiBpnWd
FC2DHzKViVEdjomcDOUcBvskx1C5kzXkVML+J8IhFCZwv9onr8bF/uew0vQq+7xWkiKtUO29lrBw
YwTI1XTtiXABAsM0GsIy9qu9NIK7xpsvd2EieXXt9hqIFZIm/Ht7QXIizy8r9xSNz1bVWFt6E+Y+
V2h6NSncaEmxNnr1n72pTYNXLQaQWGv4iA09HNNOlCWSpENvn/jDewZc/wpoEFm0Y+/l+yzbkOVc
lIGtSqZmMvDH8xrTUdR/R7VvmAqf7u36tBrmY/MOB3lsukVNbKkEp8ngm+qqAxemtpd3RIfmM5YJ
IsYI5tNoR1at5TtPGDDH2csTCcsaE5tcApPremSRzBThW0iASAbqpsdeEe3NdNhTbvXAejydM7qA
O/PqT0zStjn8WXG+3ch7Q+Fw7cS/7FzA2lzLNuMWXd7C2PIdE6BTky9wALSMsGhfDqtG1Z43Y9be
hhEOakqLPvZ0KriKiXHKWnF8neMKJXFevI09QOBQEtkwNoHA0H5ZG2H2cEgWzdRFavNU0+Mo+Iw+
tiFina1OIZLbzMLjbHXgez5juvzh6eeeouKOrPRCF68e/2MN1eKM2DZ+ecbsVHnp7FpVCg99+oct
i2EP2jC6Nxzbi3eP/x3fexyrgBrf0BLauQmP+2BdPby8c4HfOpIPOO6g++PQpaCm+UpQH8zNmitq
b1bhvUj4HrHYCAhpgRhP/BrgDNPcLhgrVM3pqXYYpD7J6pB5RJuEntgFbVngX/rmGq+RIXBweUOG
ZIa7f7txGjX39FHJXLdQ3phYlJbn4rANuL5uSQOy1InnqFXukLDO4k/ZmwGnOMy0lBNGC0pk8JG5
jf8N7hkIX5JlbnLdFvmODkkJD8yCldjnJ0QrSBRQo0uqivnvZzCJQnNMFEmkl0PRyQRYy5BzRN2I
BKBNsQq9F0m+2N4GsWv174F1Qcx4VZHMGbzxnZSAM/NbE6rO8rk3vG+Db/2zsBxFAzasCuzY/ach
j+cHLIYJlsZzH14MpxvaIzhqhEqVKcv3LML+POSXpW/0HXIRkJ9d6g1iqPNfYIHXK4IefZ8Ur/QE
UEsFp6nMwOR2HxhKcXNJWtwp63pXQW6U7h04mi3hNJaPwuD3XhBvx0V1i7Yjig7SLkjba4LoxULb
9fmfIPqq4EvG95ZTrkIU5eYCai2FMp8iNTnujSniv+2aHO8/GDSKQNUad0xs4iUOekE+w4zwLF6H
Zf0mIaQDls8oPEiXqap8pl5tOERa00jl0LOnqImMxAtYaaJ4fdcsjhCvToJw60Uc2mwtBelunSy/
m5YzZtTmEOCKqi7XM6zoU+j9b/BP+Fa6OOCtF/wPBXUx6qCAxOuUahK/Fw5R5OkLbwFJXJ6Eh727
e69feV7xzggPQic7Yf/01fhnV3G1gIIIf2V4CszA9ehoAu5Gv+yuVXGKtcUfAElS02U19b2+OazF
nvfalkXFW1RlVEnTLF/sKNWfd2yClazEkNzgbw6KwF6iiy/Bs/iFHcIOlQTyxa58ovpOeR9ypiLh
Izwd2V9i29HyFJuCIRxUIPOkR8qEgi+NKuVvttW6Mv8082W0byzKMfINzpP94uK/Nvnua5GMzUjV
weapLfSHHOvVoIdzGPzUYMJhX0QaXMON6xzmM4AwQwz5hXMzzJ1rLOmXPUev+m33p3frj1uN9lKB
A/wZ+yWICM8HtbEPrc0WamERlPyNzz2W6Tk6eY07f6sD2w5uqHMyC76yMkWQ+BA571xyN1Ck81yJ
gIQ8h71Xqt7VKz0Wh6KkxweRiYvoJTopyGTNSHke6RvVP+BYB2HZ3KxqmMGTfWSN0UOallVhDwq/
0lPpS8o7XH1D550cA5QnUtDmDJx4iLX4CpYWRZTlq80hVWNbPI8a79Dfg9hQqRTJmodX3HH7kFOx
SzLZCtm8BY1QIjFBzUk0xFnErwshDAn/6Db4KFGiYZVrvlwR57I3t1unavibiEAs0l3jtGEUZTNl
sPl51enrK5nPOzdJQP0+i1eSGhZFbzWfmrq+C8XZ4A+V4UElS+DFo0m5QvEjIMG5JGGGZAb/bhXA
pJqVGIu7rgQgqUrwY9167EAUBlwHDLa11hyp+5EJIPYlXfNQTG4tQfEVLNi+nzJ+mvlh5tT8fGxs
3qyKCLZ9mp5wAuBqMywhVZZ+h6EJuZo8QUJzoo3AWZG30FAB5aWNXFfxNgD18jomdjXCOLcIFuG8
06IGqLsbYlvzxeHH7GTvyw2LWBjvy8OC5uDbbKW9WHd3gwQfNRNErdoeyzLUMlPeL7RhXCpPHTje
S4ERrmhVM7Vz+TdhawFdYWeSAbUc9Hot09f/lUV4cOIqI/Cbwzedc4LNy1IKjpA2RU3ts0xoErqb
WcppE1nRNn6EhP5yb4B2J/UEjpz6qNHtTkw355OieFf3EC14ZTfsdIEBYvZRxBPhf4UBSFcRtP/7
KAgrqjZ/u1y8Ji6rIDQ/91WBl2Ye+257UNE/Pk1Upy9IaFFjKHJhhqr8B/oDM2dj/d1Q1iN0mWIW
v/grQAAnO8CQzq8nHoBsqUyJTdRtOCNzpDGut5pITGbWTv/u88NEreFais1GKBZTa2iS02FrZEUh
YyWCml29mj99fVeu1pGDwy4F/ZR69FEjgwv0pj6KFHGT3BgKTbQiaLmhEVvku3mQyqPGWOvmRqZR
R11y61WDLgzFpGzrn3CeLBItZC+EvDUSKmgwqagw6fd/50lrWoNCwpf7pls8+hcIVFwmLVt3JPUP
i5jMjjSqyBgnlETaGmgAAXcVIqZF4leRFLfI7j/Z5IrCT5leizpZ8M6+rF+XWVh9ny8CmFrZyFIJ
gJXji3NMGkf0EH7PfiigMypw56YMfJJYejk6wxR2Kw8AnMhoCifQ54nlu9/+5cUngMtMSlZtlyuf
AjHamUJXy6VEBCKqDJc3Un4cKqAJpagI681j4ZNE6q+JY97u9a/eUMDOCOx14t2O9rqiRcJcWcYB
jJgPmzUUuX7M49i5K2Gwwwm0ymE5yMAY4DTqS6ydqvlkUtJsVisjXUubggsB5AThw7e93dy36QPt
AvqNkfUOnvTXHFT6mw5fFTCvJroq3cWVNCkxU2MkIwYDIcfd4Ai3s/Vq3PYXOTVO5YCCINil5aZZ
vESC+85dskXrZkPzhJTp3Y/zAB7z5zUCRd4K3K+/k9JywPizvo5VyhZr5TYbYhtYp7qtKn9bhyUv
n31vqxN0Szj0Zy4vOmHRXXbtCyDbS8fDHbxdadNchffZjdt0XKAM5s/LaRhTWftj502gEPDWXD3P
Pjdtmr9keibRhWIqmusW0w3MUwJRVqcs/b7gblWvFoKZZoSWtRV1+bq1aeT+Rhmb6ZCSXrKC0lwh
oW9V5T2k0JYHn1ryH3uoMV251JE79escZerYOBM+VRhfhELtRomJbXmmifRDKnTQmN3NGHV8bOgw
CZriYHAX/cqywSsD07Rpob29B/GLACBXa8Zx8FrWs7374lglBaNcf+A1X1ZnJmY/ht/lXp91rD3C
SYhtAjBF4c6aj5WAKzSwC5Hds1N4w9FTBw+hZJUHUntliCYvL2q4Ktv5IPP6KvMnrolowKD72zrr
Woe2AT/80c3RT+e05soYxOsE2cP62y8QDM8LCAizv065Js5cK8zfbHc5zE2usj87af7eZTSgKKO7
YmEWRf9ZznmeXcpaaJrYBUJH5oeLl6JRrBM/wnA28Rur82bUG960XVwvBhqnXanSQkAJuoy4ShRB
x+NcGmILr1JhCPXblPZPybGtBv9y3POB67AefgaEzLRhMiwE8zkuC6u2ucn9oUbAuUP1AkOMbEW8
ED7Q+q0DWUw55oGnQ2lue0hYWMg9Esps2tVmlokxtPj8rZe2owt5ie+q9vex0wfmlfjcVopyfa0u
9eMFlFTxA/93INZ/RZIsn7H6t7gGfEoTqbTJpJ3SacYGQyddmhiSAVt1Y2xNsvErOcLztu03Dmwv
dxUkU/Rv3whxScV/UZgj1mZDyy0pywZIG14aFigBv48cI0gtVAH87AnAzmcooe0CD/13ARWuHnML
aohBMH1bLdUNhsoay/3QpHz5mXUBbBCBIaUyYvqQGXMvSUD7oS5Y6b5TtNwIBGqlr/ZoocMiVrUH
79lWh4wxDmlteowev4g7OBGWyX5ovi/CQfWCQnafBObNVaZM8KnN8wUsXGQ98kKUbdaRRP+wCvxe
skNIoRWmkUsJbL9x+Vwcic8f5ha5zej+H/VxIErdRjhCDsjezrtWWjV95eGtTAkEkkZmuL6U1gBX
mMmX1lPF3zTn5lF3nniKpGyN2JxsBAz2iAstozbO/nny8jdjo3HSkHc2d2fkNxE0ckYV+A9FzpZF
jvbXiztcmv2b1wBGfabnGNC4iWxeqGRzqjLdRvMOKjXh3RYnCs4sTW7xNpZwiCcAGqwOvpUJv6HM
S9kgzLF6NLj3jBs1cxRX0CVsGl4/gRqbvk4x/sFXBIXGJktOzv7kShS6VDPk9r4emn6BHD97CDuB
3FJ9UgMujb5edWxzUlZE5+FJJM0hviv7PUgAEiCb9cysZdKKtZnHi3+o1OBLF+9u9Q3TqjdrKD3J
7MZSMuCs3+j7sPN+x2N7cpVxmtw8L6rRzIJXjeBU12lnAQQKYFWEXi2GMhIrc3CJptzjtVxp304i
R7rna6Nt0yPGHjho1nIy8cpbgE3GO+/s7ck7SS3S70TVMweF4j8ZbpGincDaabcCrA8GEN78F7tp
ybUzKeG27JARHW3wHQsypoWUl3YQJiZ7r6b3JIaXy5oDpQWT7SPlF5vye6USv6RD3MC5yiz+SwxQ
3AwT1DXklmLGZx9fqvZyaVLqCXyvwzYLbsTcpboWp0vILQPLBTzvKzdKtIp2uvCVdTKYfZQryyG8
2ExcDuDKWMsafiQHfbffnwP/obTsHNiAo9vi69Th+TTiFNnu+jWaFlIna10eiVutSaxP8lHsJcF0
7SiC156mMmg1eSAHpBmx707UTUFPB91wfflwDl0k5tO9N5nO0NqXPpr1ltz4A3B+VcEVfIe6Zu6E
KPNj/KyFRG2xzu3JSIyO038zaXqyGH6NFe6R6rNUVFgM83fvo2RLRpagSAZ5pjA1sXpedw2plzZ2
FNIzKbYGOfV5QAsK5bzDO2TEd4pZA8HTTErbAyfDS10sbLeyNFHS8woBwV8CuhxiP00rw0QYjQUJ
fTBCCQBbTRmzyCCcx7QtMarCzO66cflbt/84tCCPC5UqWE+w7KBpAtUXXR8ilHBVh7BWuCDH90Pu
na+AS7q3C1E5BS5oGMjlKMHxST4VxBtxzWiReMmtB2U2tIm6YAyahFuqM1KfOft82v36WQzmn5zb
L2cOUd0dIqZyqdrKqUZla+q8WSVaQA9bMbhTMWwfe/N6GoWfq4BmTRe80G4yXaDSCmbv7Uy9/ATw
uahT1nUOEq8x7EhjcouvN7qFbd47cDbCh0BOpd8gkyPlZ6GtHugnQj9wBkd1vtPG7Zglw+eiV4YL
Da4FPe3k4PFMgPoZn4hzgNPsZ3PzjvYTSe/hP5mgMpuLQ82r38gZHNnqlSkx+Yl6E6b8UB/zTRRe
e2tKxgFgb53NznnNawjNDsO35A2Wmj/gTmfdOFUdusgTjYLjzZgc8w5T9kB3Tc7CrE1RN4QWZV1d
DUEeXX7CYNP00sFdQdv6wCxc9njJbh68Bu28ZibOiuBARrpD6c50fR7ospyprJLjHtkgmOXynFEO
SGKz44JK8nyJSHjJB9Pg+GYFRBAvqM+McyDn5S5lhTS/O5oj1r7UqUkJ5Jklr/3Ffq8PgjFc67lS
IIefziqNhnIHz10P6qOyuY2hdZpx0Fj/11Ssx2z4xn8r0lqsPm/ix/X6ivz5Aewikzh+IONFFtuV
TJS68yWHpy2PYlOnCi2HEKiXlqsdP/P+biolX5oDQYIX4s9Naq0xYnDrfv06GNZJzb6NAVsXAWGP
kGR+H6pFE7Y39bMrzXlXRD6VOLjwz09MmajE8oHQSSGtcdesdyT4W6EHox5dlFNqapfzi4nEevhX
f9gk3XUtSXyLK0fSE6vjrP21AR16KtxPQ5qwpuAnnZxpLI89wyFN136dHqwFWdNNNxWqGY/++D4J
rHoI126pUNDPaQyhvi61cCNjaNW98BqD0s1l/r9EdMOWxh1fOlkAjurV91WASDyiN9xFG0iD0yCe
jzwHGOXdqCEoUTayu9kanzO7YRugJ3xesmOhkCONeumYZFvdWXOE3r1n6NfWyoL6cccG0EnT3B0W
G1ZJY0OzXLxhqzA+tAt12iyZtFJwFfPS/myu8D5ClDDxWCpOp4YgJwi20xU6aszYo58u4LrkJhhi
1ilUG22foZxJ0inm9/vEJVgsfFCH0nW25gZXx8Zy26sX+e9zxyGDZqiV20dIq18yEFTR9yZAdwcP
GKRDtf+7MyDgKXA3p9HiCYJNDIqJIAHvW7kbI42/cRPl1ACOTiZD2Y0JMQfr0ZR1dJDjwyhd1xnQ
gt+WFzoz68TGSz1pFdD9wTm7lX6Pms1AyuPpug8PiF/xhVpYsb0AmDHYwd/sN1qQsokAmOp1oDxV
0OIhVMXNUGdQBAB3ahMuv9SvbumbMNZZwLLX+UiaXODUa3cTu58wWToJL7m1bYlNxJIEyKueKxac
NcrtWusSoNlmE/q/CxedhR5DMt/qlr9J2FgxgPoXWE4KSAQwN0PDoZKp49b6JIiOZD4PZ2VtNYiN
p/OWgx/Xnrn+Vw4KpZ51p65NLvnGePq0XNWel0YL8/Idmsttm0o0eMBlXzq3+SII2XzPpSU8j4ZW
+FvkgMWgJse8d8mPLFvXGxc6W4TWUZQ+tblJhY17zedquCRsaKGUhYiYxJJRqV0f/xkQq7hZ4nYC
PaT2eNoCR4/kI4b7w0tmqxU1S/fGgq0f7mR05u/yXQFkUWnUWAQPpauAOydNAozcWftJvB4DcJJh
LgW7ZT/BJLkJX+SrnEJoQ4s6Clz+jJk5HWlvdoG7l7jtEycCalCvcjs3UhiR+VIOfrBPbyD+E+QY
ddjAaNyyj/uAMrGdFwmG5Akox+hoEucTyQk0gmgf21UCEl4gLpJzJWELriw1ES7YZ5u2m/I7thY9
MWd/Tjin+MXvuY3Hn3m8klbJJyQHNWnKvr1ifCcJKiO3THhCnQjfqrx9SSdFf4zjYzvkWv1oI+8b
U9oLxs4r++qS+v3/K1XztNJsX7eLPH1dayM6MF2eMMH4EJy/RtvJkJvq1K5rUYevO/7hYT/lO5W1
lPgzcKEQKdKQGRwHVbymJTSyjsh5w9mSO6Hh0qtKfv7o3bvYJHYoqrADszIDiqSeQSOHgSyOISso
cg80BTupx7BlsHAo1IOlmfPJuA3S1C8xrfE2DCd87X0ChPVXetO+O0kZsluBH7nxFcm6AmeCiQ0y
tnb9cIUFVLsOTaxrBhyfTvyBxHsS/F2lLL3fvtuJ/bnA9D/Z66Slme1T4kQFegHW0tAiTcxbRBVh
HfnDf03HiDYfwo/XXlPcgfqaWC/nuMRc36ODNiDZHWq1NYOwFSlhkw+brLc8Ymz20wSHGsTbYneI
Chy4qaCRLnAzpByml7/yTr3p4xhe/Bsyn9d9G1y1VRJvPJuf4hg+WcBYJh2Ng/15Q/VfmJcbVKvm
Z6gd+DuqNEVCH3CQW/A57a8MMN35PMnZZG8KnD/mgTE4G3cJhl731DQ4M4jBCdT2l2pIqC3XiZM2
9J6JzOl1h19yZT6LK1OS2kLl/z/vtLaE30bP8hxyneggFzv+rDZOmT+F/rPJe00Hz4Yaqbw3wFWN
f7icSFgs77Zspoj5ignVl1s6YHN2GG34uG+6IdkGjR7cPOZ8g1gW+G8WSZr+OE9EdPGBCHa2Rqha
jdbkVIRGOBk7rmfNfxALdBihS9mdKRPBVr6mGBUNSRx1jlnnRI49TIlFijiLVhQi/l7ht/hoZlHr
9K3xMRuw/mLPlDCX/4Ig+m/PfaGeh102nJ2SfmhArR1P8w5lz2Er7Ut4P8FzK+Wr2VlAv1gPllxR
EmdvXqbz7pKhm/1F05ZTkiZiNvnAs5MQr0bLr9WmGEcgrvnGTz/2lIH7T3MWv6TqaoyPrPgfMVFT
pshmRW/dXkmn1hE4G4xQ9Z7IymZkCRNvL/u15xt7cu4PKIWbEKSB0dZf38UU6mR5POcLmY9lyHaK
OZkDMnB60RLz6GpbjEax9irn7qi9fLgUoRRRpGZz94OkN+G8QHiR1S5wr/187O7qLNPTXA5YGGtp
YYDDGrwgaDryAIwdU5vuadGe/0Dr3OV5kkSQmsbaX1/32FiNhyx3RYupLEm08BocJD490oORWl1u
RmWtLWBB2Xx+mxL5rNI6/5gDEuMtIIMAuRENfrEwrZPrW5GIau7WJDUtVSizXroT2MrYQnXSyYAw
86nQ9drh0bprS2mUme1kZKU4y1xOEMM8kl739ndQcuz2c2BnAwTWfA3xVpOqWW9bjYrb0tx0P3qK
zR7/xgTLmt+xN10GMazKVbKYe8CThZ4TetWL0whULAR/qYa6Rf7gpHKCodSvC8S1lc4HvFSt5Y88
66tDshReb3Zlqu74vxevfF1Vveqt1wZtyab6p1T/HHdPEe6bLThV94DWk6wCeyg1JVj9nT2RzC6Q
R7E5FuYzj6FE73+cATCX5UifQ+QEtHx8GCLj6+MVFeaU/nU9oiJ03AlkxRYW0PNHRcxRtzyZubnn
Y5Myzuxo3UNOAu193VsEZPXmlyVQWSB8FVcFoZFcOwskiyMRVCbaTfftur5Owy2hhA4jyckgRsoW
p4mOb/Sdc+osBbQg+wahM6Dq/0VOBsXRPUCgBcLpPEMy6kGOihhLGCUa2iPLxRsOPynowEnea4Sk
bX/wLaaP8hyfXiTOrfD/mQRpH3vV+nXNpsVwKyDPMgme58zG1M69bZJE9m3/ygD1wstxg9y34NR3
JEBfUL4pu8t4LUc9Rv4RwuTnPmmiik7kR0ufKdO7AcJuRzCMNVI/NZtGHUyzpV8HFm5n13usnUnt
TvgEM7d365qguQjf0vl8cVIgKKa/LhpmxpQoLeetj8ch3m5IKijdA3HYmHbK4e5tHHSKpahxk/dB
/lbi4KD8SYkRYK0CcDR0+GYbiRkE7N+ywp6Gv4y/D3hyxHJJUzg1W4aZ/qjaBmL/rWQ/eR855JdD
kGz/0Lpe8LDkK6UqACPV1olUXDuHMkgm15ZVVQjGGpzKdXzhR/NYAmtmdYZBBo1FNpMvs24QdkKe
fItpiI7FRatOYaYHOzHakylDHaf2Z++70NA5KnioT8a39pf0mncBzA+cjcSg4NTltGJvc/b97bHm
q7+Ekj48agPSBZwifKbYqUucspRO1TZp+gojc4pEQS4ktrn7veep/ZD3DffTiPQ6gp7BiHW6Mak2
gotYu6W+dvYLcZrhBnQqVpNRMDBDfSoNHme2pLEXCVxp6mpuAKL+yHUCoENrbhz7xa1sOOikEBcT
t3mcXO/8Y+HjH0zMdqEdfhvi6aczUl1mEGxo/Gz7U3OxPy7LzdVXpf3JgmQSJRp3JJ7mfPM/ojsG
zj1S7ore7XfiLdZbWlgRSUPZemxTkAg82MMenOvXsFs1WjVpohJHjQfe0/ZoU8gVkWsVQpPbeAGo
UHFfI6j0t8gH5I77Dap2rs4y3ROPXk8ePMXlUq6BBsclc11V/dpgUwZch94IZtHQlbCe5j2T70eF
27HVoem5wbKIYOyL3zp1J2tX4jZ+LgpyBlq6MXFYqxEkD8/Ha2uWbWh1jPEI6NWwq4KofaF8/r2c
L35jQHYg0eebJPxjDKfoaN92wQvzOy3IH5VfaICqPUc0cy/fX2HzMQMXCJ1pkP4Jh+6x4QVJKTdH
qnGDmqxSB+gzMWNX/5+pJrzNy5TLUterMxQGzFprQrlGdPWhvAF9nf+8N8yZsY3Kc63yJEWfNFRJ
wMsxyMqObhIO+ek1ZH6iUPtYONQ5gdSc1dzJnyO/3VlrrOw6rdVzbg8fossLFXOY0JGVUV3mGn4s
D/67yBBD/76+BJa1Nf/cZmRRGU539KewiYgSAh4CM0WK0UEn8eAiddRDubJiUQWt/7WKwhs69JLL
TG5QMyHiKD/TOouE79/PRCgNAFOoLqvz9cRxTF1fPuEV6XvIlIygBBF/lVWizN5g6lKxUw+9fdkn
9WYhiLUVV0W209h2I/Pwr6N73VEoN1yDmedRui1MTyZZcExX7UJPdXJNci7tw6ayuksKqZZqIiFp
kLJ0Dk7xC1LAb6y4+TWGh/r2cET083OufW8/JxxieGlaYUcSTfIEOjQBSERQjOKrwmsa/tTyOSzD
hGOBbzf1izeVh82GF6KXw1BewBRZNbfxbKcK5nMbEBrO8PeUGv1yI6mfBqJk7C4QdNe7OIox2pTz
akQWzBhhEv4g/bNVyutUICkWVN+xvQFmWOjzlnKEvAZAFfEFL4RTZdDlIXUCN9wAIXwhdNheDtKu
oCybfruP6Q/SI5xeGADidStoyvKwGyb3OPp+ApyfD+sgdL+wvpXns9nRTRVDR632rmlxCFeecihU
qZDLnwJBR1NQwasHBmdoQWnAKuATr2pgFLtOYqxhL7n5KEspvJqSlPxa3Yhq0KKdjQH4VBlCI6MU
2vibdBIC3DZrcijC58uEkbFOLmG0z9dqn1VyjfvQYRoOnVmASgHljqfmltHrRLwPZgIRC6tZBYXM
UJeGZdx+Y01PdfBhZ/qDTUwZqdAaC1YfAuDq27Y6reA6XtbwaZK7nbTrKOsK7XjJMYZ+Uq1PfAXE
9o6fk1kmxnhGKOKBphVRlYMhHlcAXb5hFyru9NKolt8WNYiSBJhQPn3UfoNdiGDgM1k/QPccxfQs
iShQQLiyj2f7JyPQSTtDMryMfzAE402EblqXNOAlFI9lxCqg+nO/15dfQPnXGpEeVU+PyL6NzmZa
DOz6IGqyWSPsAaXKFJ8aAACxxr3dWYqBIqb1rlUOLZJ1Wj2p8tfoZJsFL1/P3ISw9P/1p/YxPgW+
1W9/3JGMZ+EOym/WPeqgF5iqHx9GG4qqPtaVDvyaGh/BVKfuMTUwYQL+5CUwEobYkeoBPfowMR7F
8gHQ0zD/ckyS894CEwnzspfTv4WdVfrdb5e1NvkKpPit+9rriCu47p/MV1p+KokEKVys3Z8jNZj3
3VQ9Ui4UH0Ro56DKthNwVtyr/lYgRl0hTuRE26JF0szPE3ngaIQ01UhQA5l/O+2iPO4T66hZ+Y49
xpvZtFgwTkHWN9VvF+0tvY4WkLhhGWx4xveMHXRGuC0I3tZI8OrJRmOcoUeeWZP7IvIKA/IdyTSy
2+Z7gyvPWTe2k3nci5tnekxT5bw7a0jQj2j/O1gVzGKcZOI/5ovYAqf7d5hP6F/YYc2YRyCOqRVT
C1N6fl8uckY8qJ3TuR6xKT+YUM0Kec1iiE2KtvKPF1ccVTsTY7CUpzYMJ7AEV0GPlJqVIs2knPSj
dQslEVhaOve/nLaFcn4Qh5Wr8AJeRkMIMfxd3wlgcKa4woq3ehCkBz0e7tD2LZFXDqZnzcvQ0jlN
s8OpLdk69Iscw176vOeuM3YNbIwqw1S/AZeDQaEi6+p0fWNzWo7xRhWYEzZaZWtUlzsqWHpnbCwP
sgmupj9sfptC9mHQyaeumIL1irogx3Kr1WbG12/EZUv6yyMBb6MZFYU7ZhfbPkkypGwLpxK4WH0D
HiBIuDkEeqS4KRty0DBabf1zAFVrbIYxW3S97rJ3jupP62YBw9ChM/9K4go9VoNZKqP7JXQayqKl
Qo0xs84dsFo8zZ9hfb5K/qUDaKDOuh3uk4VTQrgGjyQB2X49v0vNkV3UpoXM5f6VP5b6S1XNX2yE
vRlSD+WthDGeJ2152WeGmdEQY3eXsINm5CbPYUuvpAGdmSYRALBD4Eghb8mUr9MHQrxxNd4hTAeB
t0DvVC3kpT8m4bBL06IQDU4KU9LcLERcgbF9q+6IabJziE9GlddlEie1VUmBKjwO388tZxeaiWrf
PZb82FP57ETEcdpccuG7oZrxrjPrwjrVawkcdL2riOwbBGJXWI6JMiaejmO2rIFeJgJRLsCOdohe
VaIB7lSqwxDXrVXP4T1ikROcdxK/l9C0pyy6HFur/4aUzeNYdVjd8i9i/T/4Q4crrsFCD6NE3a00
XrNjY6ZlMwBqd/0gOepyYNnwLUuCrOxlLCXCiThNAh8jBV9Jejiqlt23sZtNHj2FSR5nDFwu+ISS
wkwQdtTxNGEBh1N5yiKkAbuIsfEhx+nPiEe3nX5HcE5NNDYbNuOzz/anwP0StrOeYI4OnJ8uz493
qMMY8vE6qjSogPGJUiobT2WxyehZIKwjq61Hqv+xrND3QSAzdWZatJzB3fmZ00Tf1up4jP6WV0Jp
PYc6ZdSv3abELMUbZ2Mf2RoLJV5Zo0O5ENjzY39juUH8HY8r4EXUsVaiQea2/KCm5Fy6EHoBH9eh
hBQAJ6JZWjrDG2jH/erPpft5EqW9tJQC6EqX7cK3ybbLyZS/9LggSwSFVyDftPZyVY/9j+xyje5i
PpHmkRjH+/JL07VBeVex0IfIpnaevHu+YToU9tgGhKc9YyRnCdSoSNlCD3TgEI4RJup0SzMYo108
VeQJqHN9XS/G/RWwPAC3Vz1Osutr4svLtzXzeY0VcVfyaXBrIW9Klxs5SiEMl3WhgDfoYovePKjq
31EUwxZJTYAYmMDeY353CfVmEkrLHLIdjVR4uV8YOFo0c6Wc9dKjyn1o2W8sHQGW897bVDpvwJ63
Nky+uttQ4kz86f/npfqMj4Sk+0hxUM0n19aGoFVayzSGjci9x8E4F7v/2YWge18SRVv+bhZvZNn9
C4F8iD38VmiAQ7FRTuR/ngjJSAXqz9Ybpic0U0jNeVgMudRZgXQgw0DapJZx2C3lznEjQrXWab/E
iBDkyXmeJTfmNNo07ZwU5lyGZKSt+8TYOASpNZIx077QW2bedLStxiozN8q/IT+Ov1uFyHvfThjh
czKwMrponMCebq/WiIk4km19OV8m9yuNHXbyaf3K13/Ur0vRmqGs65c/e+W36VeuPztUp14s3NWG
oExFbNy4kQr5fpg7KFWyq3ToYplboR75JNADfDDLdwXoCZ5AtclTyI9xl2S1jUJIDjwdcy5U3qck
9y8yH5PoVlNXc0adJHklv0RU/X3/5JlHdjXYIpsZUQil+50hXKxie/XBg/3HhwNfW84X7xXexH39
pY8vCGj6eoyMEWPIpoWAdPKCaRh4559c6E6nyRJv/I6YoA0x+AaqecLlh/Rwyfj39tS96izDpTcD
cpka8GM/45F4x2EMkbQBjFrLr0zQYCGOS8kI6AXYXhCiUQmeC+942GJYvf7U53ruy+tqLH2qL3Pu
NkO3SG4W0KNVJMYphnfG7CWR6YtHBUtmqKVpdBmA7Yx4yhMQYkmBUBDD7WgJItJyxKShGaVHtz7r
tYdGtZ/BI1zULNoJfdjGXPNbv6ktMug+pRhA3L/hfqSCa95GKV7FcW5RfZMzAcwPPaMD9WQgpEKs
X4ebNUmNBfbSFdMayEo+xuBmGXEbmR8UHslge3lHCdrYQXn7tj44/ZCWQfW2B9rscrCu63Z5pG24
fsMwnsPCcYG1qx1cvZExcfYS0EUY9WEY/Lf1yKnYqw56Hee0i6L08KxrFQN9CV7oyIWxsPj4/wE/
GYdEH3iPskwZR1sUOAbe+NQmWziYTcmQxbv3H6bM4vduBoYT8d5ydjJfql9eOCgm+MFf0OQdCHN3
dAdJClDlwEh1dk6y/WA6c3fHvmGN5cf1hnV8IXZF7Vzb0PgiICzBOD+rJC+kBeoUAz0IPVFHMq1W
0ZbRAS+FI6gD/TaCIbb6Ne/EtCbfM88QcrzWG6q65lpM/bh4nneEFFJxXclCWFJZuk3WtJ3zkBT8
1PY2w74N/rw026gC/S/mIDv9lBNGC4FMc4oxM3yOCMH7NMyso0/+gX0Ub3zMg4PPqh83VV6gN9St
63P4XLplgJSKzdMfGhbrOvyQaTDFsbIM5u0pBP8I+l8LOIAf1nAlib+CaLtH8P3cPf4C4dYEsDCN
+c/32GBRWaCjyzaJP6RymBf5OSxial0pDbsd+ky9IkOLwjPnywNBvW1xFhUcvd0znaaRsU4CW8/H
E1dLNdU7GXwxXqkqFwE3NVsUJKPrHmOa39joIA49VrDHFmUvdmVZcsmJEMcxGNyel4Nq0vkKJXfU
ER8alid1u1Gkl3nF/Y/0RRvvX5MFwT4YrK04jyoI5tKzIFzTHgV9axQkse31sL4i6+uouvz9NYtd
5v4M28JHVJ3K6qkhL1OdbGxsdOXyqDzevr8Qg8fONr2834wescJz1EQJuZUfIMuom8dj72esWPv7
rGPl1UH1AO0pjUEWumpgvvQaydsFDfW/+dkWIvwOpF6SFutMIZg5naK7p3HV3sViECwdOPHeGiDl
v+x/zVJ2V2BmpqpDPgCmmi+AHXv69AdFGiQYwtpxDpBRjrPeNVVRTuqYMEwd1PRWoNvdrdzgCs6D
3+GJvLEGLrN6T7YCpEvRTMU5nH8mYi4Sbkw1dp0R6+CCSv6D72EGrSx0CQyBNGFMQBcSichRzI0B
nZ6MxcRqnO73NZ4q175c5NXuWPgFUGDo6rsczGSyDgN0YGk0VZkRH9ll/IWw+bH5axCfB61Y8JHv
TPYeLd0kAwWK+DRdDmG6cvt/5iNeLJekR8dyuhfYpfZEMDwiaiiWjsm314EHLO8zXwPUUayGB+LP
0gjYnGHIcP9vOOCiMJbZTsWHBAmQAhfqDX6Hy5l/4KT+0u81vKzL1HlFOLmKPNZUD9JqmtUYCOWP
3A3pjALBOg8P5kEsYTi4gdUvHfDgKTCnGrNXaK6MbiLRxSlrhUakHfqorAbVLqwG8x5k0Lo7HEku
pZTB2IWo+K4PgeR5huH195d4paNyhk/oX5lbib8uUsP0VLnHkBkENHiSCN0xc71Q9oOCnjMXQNMn
gTDIaTcEUd/Tf53BXjRDI0fD/bWLc+jVZqaM7UsH86ml3UO/gHjxIm8xdyEfs01ql3tkPegn+v7P
tsXSw+xy1QJjBpdn0Jloafkzcd20YEeHZjwNwjxnKTP9WHN1WTJ64V/AqPxY+6yCOHgHm7wJH0eA
ovkPau8KRqL6Ifh5JaLw0IaEO6k901bLDOh9P9gIIoaEDFx1pBqrMi2MEAb7vR6S1Z5p7FuqgaqN
KA0UXHeTg754fgfNxY52iTx+p+8uexLQynobWAxm1ku7VZMNJOqeYIXMJND0LX1flw08eFBGaahA
Hld/VNg/5zf4gDm2IoXhJVgCw17PCPmQlgn74M0vH0I0rgGu5OsByYUBrq8hho6FUGaLqnZTqO4f
U10nr4dgiYBGOTDTJ8v+HyXhW7kYGdvZ17GG3QZyhI7thoO1A9Ssg5QPBfYMIgn6HPQVFOrJ0S81
cLKwkAiKb2nfRn8dWdVV3OdBISihWeQZAfyM4Lmn7Mk0hVivXOLP34/I6gLPFcqyGPJ9/Y7Mn1yd
jGpBh710x1Art1ugpmP7OEez+08rzYkqvscZxWRmHaC2EWaUWVKM05xHES/Uoj7u7GUQwE6zXivo
gdF1zRachnZIflGne6VpjSXPeVdgjg25YulzsYdlpP8oO3LKQ2jlwetn3QUnKg7ed0SnCY/BhKo+
clz/iVrvzN4WbmadWfFA5ImPemJLV925SVBB2wrGUoi6sEOwK1XaOAGunkO0S33E/M88149eZuI0
KMRGUdRcMO5cC4NbnwKMfWzYYs2nzgYdrjvcwI8KWXXNVBpJ9FMwp40I2Plts3e3pmNofLaWaack
1Rq4sI2MVgDHx3oGUqozttUN4FHdt7/0TAMHsvt2wQ1tlbQxbocO830eCJEYcvWSPyRA+svDdpUe
XyfLMb7yrOxYh5KQDp3y039qe3BO2KLZYxrNTulLPS56S0SuEfUqR+xKZlxvIwCVkoi6MqqkemEO
s5IikXBsqYKjKlmByxY57kZz2d0sHqteVj3pcF+8La3JZyYYYCxpW262RhY/EQxyjVoyCn9e7gbs
dQBlSOAl0gZBIhHDcTsHTA2NEbBT9lwDf1mN+r7jnzR/XuDZ9s0NoPElEpvj/KnmY77G5fvW7rcY
7pG4Bc71rK/DjvjBldogWd/oZGN+ieJ6nzU9YQIJ2eVa+S1qYZemz9M5GYklcB05sAWbQFi+4B+s
cAl7X+tn0jkOTmyiZjftl+uVh1o2e4jxQ7VzWk9KVManrhybF+PATZ6ZJcq1XznvvfvvocNry6cA
XJJu/jwcrh2a1xrSCzsRrPsS8pic/fP91fgoWsT8OzmYwQbt611rY0fNgwMxdqvz4iADRKmXBq6Q
VKwAvEzn5rOUPI7f62Ma37CM0/SHKr+fGXr6tb40jV9xz2PFBIYXACX8RqRbT+ZFbb0Bt/sLXdzC
PcwXbuDhukcs3cGU6nhh6DWsA0kAh1vQ+AY+sYblcCMhkiy1fg9MGBCsyjocJf3I/gyqjp4lSmyF
fiV0pHRq9Qh+7KRvC47eM8Y3oQyguTijlNLfHrpCcwFmOFcE1Q1jjKlzP4Pt2G17NPaVYlBSpUJa
lz7ssXeWqvh9yTWKWVUYTUhcp5f7zWdBa20qqVTLUMmfeXeZ8re7kcUN/FhD/+vI8+/1PfW5g0xP
5ZEg+OTzxJy/AQNDFjalhm/mwGGVUKPM1udJzUBRf/05AQCvginWETGR6qp8SREWWAwN3xcGiCyE
OEc3LlAXo0j3JFXMsSb7xei/3x6NsEdGu6Po0bzVwfIFkBmQtwlguTC+2KxQkKzABRD658Qrn45M
bq2QJfPlm6TIsXuvgHDkNsDiyYrBhUAUVys/VKQNHvJw4+6z4QZ955FZjFSI2Bwi3BtasGixgbEN
QuCzntIIQKKE61Hc4Ha6tIMYwoNgEp2Xp3YM4BXuASRgwIMnDVXiEAS4x6r72+eBqS0hzTceg6pm
bqpmM93KH1FxAvwZW2QFVUs2v1g0pfHYyBzPIeLPvNVYoXxMyXPDo0l9fQtSb6OjI4yQt4oR0MiQ
wiTf1V6cKsl/0joNwGydwaMJvFEOVDvWEDqtrNEuk3xSbTKf0Q3h87fBvuL1ntJUaEpEIe7dSaxo
hzepE3BoxeoLe8j26NzSTu5LnGeeJCKmANqjXrlm+vLoBkWIJn7PdwCFZf/aqOlA1Q2Dj/IyYO+Z
EfHl4j4nPQx9zEt8+du0/kAoXrJmGt8CY4wY6tr18wmqyzHrQT5MlqRSXeNlhfIXCNlicxheCFMO
kjo9X6asqxDU5cPMY3PzeO413LB80WaX7By1zxi0vqgPuG8AJ0DIF7sCRlbkM6cYnijQlQ2Tn5LP
iGBsiWbttCd/WQhYfbfatE4T5Dfz1/z9nlYNv2gjQRsImlkqyf2JYyTT9/bPajRi8UTzfSZhPTgY
9vjjImz0ZpInR3P6VCooGVCaj7KJm82oERmnUu3AAUMv79uYzjz1Av456M2djPjcFE9Ggc0b/54/
PI5NjAUdpQA3RXCsDacvTK4VGyqoG8DbEdCOm6rhHYY82Hc2f642srs22LuDQqyhNtYT+MPdt+E+
MqTjB/Cl+t4NbbKOHKXXASsFH/b0f7uoNNnA2v72QM/U7ofLHtRTvPv+t7p9LIL5PbFOeixiKnDX
pOKEkm6IaI4FJ//3OQXSK3NhyJg2uOqqHjExiyGlxa1MpieCUIgja6emkCku9q+D+ky/2khvcVH7
k/GwTyiE+t3EIN5Es0MIWM47Pa8ZYNN16QtZLQug7FUCBvtnSRiAMFvvBgXzgFaX+o6+HJwcESLU
QXn0enUtYhLmUkUywt/f+Yb4UsZj29UazxZ0Iu1O2/L9Z5r+GTrrwhNcjBzWFAmIReul0uSw4kJj
rV6KQuMqiH3fBkxIo3jH0jb8vHw8JFTnFgRyxOBaiOk87eXWpTrAB0n8W8WjGDr1KwKB8ZoJ9H2m
kUY+UCn1dFAqjqcKu6fcKWQH1oz3DDnNKti8koNQYaIHNizzaoHvRkyMcARCoU3dsh81em8FDe+O
RqmJ0lxXqw/p1O2kJftDPc3vNiQlySfXPl7J21BtNJRW03rBNhBNuToApsijjbft2Wk7FhkSvMjR
oR2p49CzT7nMTEzU1iY6JC2sXNhRFhmJKd33hakrkgi4+RqMkKZtG3SkDv8YdnD4GSBQaW23PLhF
Xmkqz2Ui2BI/TdAeTEG5irhGivd9XKVdKfRHVLatrnqvEKYFmuXPE0u6pmop1R2RG3L2PJL5ya0N
xaSeYISab+3Yfhjv/W63VSMCnFBeB3t3mY3pdR2cqWEQtuYCu3Dq7N0opCgWwUBeQ6o959OQ9Yo7
CZXlS2ELasw9AfOJyQbvIOkWs/MXRJTeSd/ReZluKw2ruvxabugmTwlOLjxLhV+sr/JrL8WBXyJb
16wqswTo/oV01RYMkpYS0JWB1z6WNneJBQj0EPjhKIb8AYnatjenSx10wT/dfgyyIEKWmJZxhFyJ
Tu5DDM+SyeyMlBrfza/dqacxCqU+nBoj4GTSj97fcl4MabX8Ua7RP62eHACOHfilLhgBWoHw0SZR
6Ff0dQ+KWQ0jydZpo2vasArg+FCETT2GwOwfB/3q3j8GaSSupZFm6gD9KBn2PnARfLoyj0fCJH4r
4fiYR/czkoi3dY3gMvjo52u7+6b1z9w3yL9Ugj7HZJef3XKZYKbB+lZl0UUzD6VybP6t9ZiUIclu
FwIRwUAz5qcWznCWXi4r6HdhZJcU3StYssm4X5GV3KGD81BDoaTYKY2I9FYJdTWlpo8HcBAn5IEo
P2sPdlyD1fhMQQICHZ1e9chgHrwfqSRYEUhfjhZdi2IABbpi3iGD8TxJJZXkIOHqzqjZiYw1SlMQ
af4YAse3Nk2DQANZwC6MAz6NglskOICMPJCKSYOHsL+Woj6Pbo9KvbdUKYcXVrR5kudlilw/SJag
GC5YpUPxUE98b6S0j6SLDhE0Koy4xjqdk7mwvPcuRNvTrFBRM7Rg2QF2S6Dr96aHhZ1GVsRmooRB
yEF+OsEinb38AbNSXKmcIREE85gg2MM0MlpqtqMyAxAbeeF9VHmURIBZrIdwnICZsS3puh2AL49M
zbq8UapBRTEdSwcf5fV4G52xXjnYtEYJksorCDXrS/zp09OQrXPOSQW6TyiqM4F2ckGapIreXx9W
NFwz4DVtM/3bKt3Zo9S72RVIm/Q9ZrBY2nt0qH9SaY8jpFgCNW1jfUKT6DlvyziwuxNKWdocYCxk
ye4mfgyDapdiCZgRyOsXiPuZ5Zc476DBONeje7qlWHTVWNAY6Afhqp8hr0YTKm7w/0gQ98aYgjxx
AvpOjQan4xmfo2tZsfxOEzjzlue6D/Gwza10CjTc+K3J959xILt6fwBpIkTPq6VFGrjgMScqTI3c
PDx2Z+od/DRuAhJRHCMgJLPZwJuMwDGm9SJJjhJ2eZ7ZMnDMM+KE2Wm7cLlGYnSGHeTrkuElPEEd
Nseli/huSSq3/a2x0ESTXrsIuZCU8Ga0fkbkq4sznc94TGZASZVqBA2BrIgW1oTb9aU++7atMk8X
dwiukHllZTrIHfthIzVl6WzVdCTgdhv0Q1aB6kh9lKDE9aXsmpA8ZBXIQNTjZYgplC/9Lc6tjdy/
ghFdhDuOdPkfduOpHyPEOA7LIDx42SA5sj24OS6tSEXFi+BR1gzOngT4ymCOtPB1an0htYhtaOLi
rI6TDabKxS1nP97x1QiWYgQ1ckgn0R2EYkJTjw/DOJ1fcyAcRd4SG2bFNZAXg/0A5u+G3RsSqWhA
+DGMs2dqc8jN49O6yRt/nf5KcJEZ6Yk9WPsyfowm+kpGcdK3jM8jVabGAWZkGo5LMNOx36JnaH+l
TtZKSgxG1n1iDKSte7L7xap+QGCvEWQx0xyYdRAOBMcv5wmso3ImGraxZzeLtwYM0Cfb5Ly1YEeq
njzn+giz+ss879m+QAXUTTvK2/qjLRKO8N0zS1mBNmmDaCs8oyX+PpJSA3UKjvdT/CYs1YNL3eQ4
PfsplqqllMPhgZMSRqdk1ZtlWdEukFJOFc2CP6HY1rtBtBWGYAck8TTAbtCxscl880KrqzkqblZU
d9Y29wIu6VYHRGxmh6qCyzwk+ZYkJ74KRyq4gS6OC9J3EWS76AU1i5Auh1UjdvVmRrYa/rVtlVDn
HhfvOEZk4Y4MC6qaZnXKEv5bXI8BoTnGTsCU2byzFOPZdxQ+SKDylVzzlagAMWCXbunfZXIjT1eq
DdD4e1a8cMcnD2+gMqyaLaxxT5zRPTe4Ry8IjaX/WgS984kqpbEJlt9PK0Qgtrr17UgBpTs1TcQH
Mw8cFA4PyCdD6rII1NvcA8fioLHy5U801JTrV3rZYUvtuTha3nleGjunFxy5LfioSxooe2bmG5Q3
HKpCmUzwstWbV/FqFEZYc5XdYvDAN08NljvVW5axlUE5r6p0/eVVVo4Dq7//5y8gHt+kt1Xs4kFQ
oj9SK9NpKJ4pHWSVcTLO8Wqq39LKdlxCQ51qokzmPOqorNbtetEVbsRHYcYqIQA9lzc83ttWH9M7
xoPN5gtqJXOlPhdSGFrlII/l7wzn6Io6oWxjrwhwH5l3aulEFQfZz96qyaCNwr8gTWPvQH6fFzd6
nHN1S+tavjHXteDxE50ajl13B6sex8qWzVbl6m9CFxQbunjeudq2BpqxhVR7vZjPxLzdWwAX7F71
A7AQfEGmcOEnW9wSx1MufMWyrsm1gZDKT10Wa5LkbbIzIxXiFmiAxYvO4Xeclzd81/89eO0cuew4
N37kCMIkUAg8D3mcpUQoaXmlxvitpWyjlp/58FjZUuMEF94QaLj9dxbuosEjQ5rPBoxEzDiQsicJ
DhgSYKl1eyVW0nNyGZusoTMDwZrb8bNLRLqkyAUrX3O2CpP3DlJk/U1ideHFFOSMJt4JaRDixYT6
BAXUARKO1cag02A/mdZ6az8KE9tKy/XHZykXDRB4ZvreZUVuC6+PtyA84Ind9553gDsq92tUVNi3
qsnZqTQgsnAjyOksR9YRBj99F3CRQl13N1onq9Ys0Co44g8zXGZDV2zaP0/ePdVvsMkOmLIVmCF4
hldxl2Acz1R7HUj05rYrnCAWI5fR/JEycUJKiVtM5VoB6WLZ2iEzG6loSkj/mKdFZ1xv8P/+4om8
6A2ZWqlORr9qRFqiEoi0U9gRCvOMM6t8Bz0zwq4Eo4kXsFCvSAcxpLP3jhJInVq0zW97U8FTGHqp
z37WKZeVhPTWxG1Rmptm1juzLiEa6jNJKbxWbj+/hYGBZK7SyR44NL/qGZqk6eLzSz3Bw7bM8zhU
qzF8L5KbOoxl6kqwBYG5NE36L4efi1ohBQyoDK7XYvQX//BsytAZ/3p4SbFXQRyaN1RaEmlgqbgs
5jRXH7bfO93mZY5a2mSbkLtTwwkKNdkYOJS4sgtQHtD+G0Q9ChTXpIPq30v6kS4WJLLu063Y3/m2
fEpqnn3Ffp3QS0lioZZ/A+ZmB7paQfIJWCMb5K2Nd2UjWxyiHNas4dT2VwUCDXur2TPQJrSxzmVZ
q5nwChV/MekQxRP3fvk7RW6iFfG/OAk7UFhfx3zXEXfHHbttDn2zp5v4TF2Tpww6aFDZnfb+C6aB
7qn1e+86DIlypHsp68KCKVucHMiUSZDuKaKwlcNldW6fZLvrrrszaS/bE4Fi9bzlSYjcL0NgvVOs
QhXZqvjItDEJj+ooYtJoEHWl2H0/410vb0Uy+K4tcb1eY1gXAqWj5RVzVNhm6YpjWzorN6l1a8+F
56lGtyVVBS8CaanZ8ZzA6/EXILS/P5z9CmP/nMhFM58+2HjrfzkfbxWcQ4qRZjTUvI8lrgNWZxkh
ChL/HfJ/G5Qnb7BalE84dH+O5xc/KX18BSxdrqMbyLjYKgYLR8VSGQCFKVNveeCBgYgMhiZ8R1xC
c+deNTHKOFrX8ZcHxd8O/tWvLMdiJpA5RL7uabDHOyLry4a0hPLhyw9BUlV0UnN19typiBSVm9F9
Us7w5xYdlk0VGR9OAOyilJNbtaKIMUppfTptZf7R9zRP8cCL+J91J9nS90Ah0IcJNq2WB77ECHKQ
KI9JpFEL6OzhwqJJzX4MKo9gLUHyjTsrV4UnvGmjy45m1xaEnmaIAoy9RIGM9llcxQ9KlhgXCSdH
jEUUELUtC5eJt//431PigS9kn5aPs7+OiwQ/q8OMCZzfqcRTiObb7JqHO9S/72s8pq3FUq7JSPwO
AajZ6V39vtG6eI2DKu94DYIIg68ZtaE59k5xSqsNpgw/UIl9+mku41yPw8hEBGOv3cXRc1NSizQ0
AjRCZQfhy3QZhq0SVKO9l6ijd47Vfv/fMVBxElpa8Tg8s0epl0RoYrJBQVWJ7tqWIBc0FkNrLbuu
/OgW18Y6XW8QGm0oWVRyzmFldIjP9JhiqfsxvAsNTKNSQuI8Fpoo/FIu9jc6tGNz80SiKw5VmVj+
uSfa+8ZeI+cabjg0T/9AFqgXBlkVqySQA4AHiubTu96p04aLnOGTx0oPt5a2Be2a0vTo7YpVJeDe
hp1yqsUla7GLplW9JqTyVzK6kLQCr6QOEhGZ3vXA6apsoQKInLZnqdWZZgfgY5R8ECt9brsJUIrU
ZtEe3mM52kMqtKtuvR1gNgJbHSOLRzRodZLWMJWqkSFyfqMF97OFXoDySs8OWfhtP6svL0xpCmoI
ZLeo8GE34ZIIByqaId4kyrxPUWWIgCZ+jXsWpnadV84qVSFCPS8Pstt2IBLgZMTqKdtL9FgcjO+T
V8tMEgWdKtOFBiUfCiuA0WMNb22OQ0I+BNe5iGjWSpCruvaNlG+t/2wPriToKFh1rCaFfm7kyBJ2
hE+JcpqeXGRJfJBq/8kHngHg+0hADcYuVjZdJggSc5AjqIqqDxtWQQUVEwkfuHaAZqVRMEICjfbP
4HPUuxJEAvJy7yBLAHvwQ+44U+AxQK5bJbgoGwC3dLfECk5LTmEZ9ZurWHCtoT/G+i9CP6nHbS6z
cKKKR1g9LUhwA6Ae0UIMPWDw9/bMRcAJJ80+wBzMQeZyEQyU5plB48Fo4tVIbctfSbZCKTX+WfaU
QRId9cRkEm9r/3DfLiwk/OgEMwdWooQcnzm+z04ZKiG5JpamNxM2wo/XVefcp9VRA1t4kpU4bUde
NG8+YmuGveufPhxy5phNqwBOjFF278+FOPb1Ixr6ulDMcLtTTFCXn39vhfbnyP0M9TF5blBsl1l/
VmyS7HS/+fQlXJbv81dJQGGZNYpjayBXLRWirYii6hWsGjWTEhAusGHkZhK1/Qs6MPayHI1RgpRl
8Z6rqRRu5Da/V6RQkxd65GgnD/PA4DAbDK0rtmWD/iiyHRpC22GoIwkmxc3TLBRoDNMNOw3GGFTx
mYBjcFTrFvoMCtE/Dn1y4k8ntAvpSLovgTyXQxOVGt0aq9XdYPyaSWG8IuRzRUJ5blPo6twT39Iz
BgEVHw0mnBHGzuKGCcF4npK3FqkejRTDVUe/zJNzKCj49foS++9xwh5mHL/ivqlhMW67JdBU3cPe
HFxgUXV0fzOd/Kc0Z24gzM7dfbmD8XflZ1zS+1Q7zFEbV4cBUsRbCuhO2Um10HdBojzDM/uvX9qJ
VucVvAOjoe0SMhoCjqcmyo2Osks1o9XTxNtYeVWdezVYU+6A6ym72gKouCBkK3BHSQMFERQ40CiJ
qc7yRzR8d72XxIqbJUjhA/BSXZXGLAiF7+KQ8zhAWKERUW1fWaJCYGmhtlE/5/G7vmZ4UbTvrwwp
IuhP9z47ddtJPm4ok0Z5PY1RZMVQX3Yl3J9vC72TtAq6XnGdlnY7jbpWn1P6Gu5F+xA8T22M2QNg
sc86ubGtnKU5BSZg9gU4yg7FC8PRRNQBpYq4JEBr7z6JQnK0x9k0w9913KJG3w7HawBy3BA9rWvc
+wadT9C4lMRq2u0InVw+wLnAj53oKrCoREfrViAsmmkovCAKulfv10r+y8TyYmNdLNfi2q6QgqU4
WYuZo59/P1B9zNP9Erf7HAhDxj4wC/Ymh7pV4o+fU2HXG2ep6dxZboYBAM3hxtGrDBnUXdh+27l6
yUevZVQB5AHQiSNu1RmGNXn0LE39MlV7ZCWkN9McGb2v8+aq+j6x1mLifUM7F3Rq0UMksqp7yaO6
BfdqJtAKVD6XgO6DHRoluhou37fal9Gxe9XpYU/3SqkJzR42myhZSl76SHvCeStUcpAaH7PfJyjg
keB0oxrNbqigjL+yWlRKkFUYyuLX1jVKGkbzAah8wMNg/QrFVAiap+KPjNF0AKCUbEWHlel3EIuL
rqLh8+UFIhjKlly01iQXtkrzWtuI8rQnA6D/+LtI8GFVkjbEpC62sIu3wOBtkR9JJxuNbPJJyCn/
ilVMVQDOKe+p418HavfXNsCFWa+oMNZWuDTJAuMWCOsfnXJXDM2cQ3j7fBB9CkwODRbLf8cnFIir
mBA/GhXhech+cNvOnwyqxjrEV51LXmzw5r9njWd5MGCuIzy5al626MOS7LIbqgEJXh9ej+6fq+Xv
BZWyB9KnQmMMcUqqtjTWe3TBIyyFmXLxQwWg1De08imo+Q+VZGroMJxRSRRbrQXlwXE6QJZ0PSwy
ZK/erOG0wAa/v/wZrfe3+RkOce0AftGY8jPcOiVOLZl8nuA5xyQ41saZ8osWU/tZ2iEGWaZi1kBf
pKZ69ses6fJfatZqAAZ5YH5a5pNfr53xrGGwR/WlbzA3HeJONIpN4sR0Cht5VOof2+Coanq/Qn4/
exmrUUmYgFR7MFxW6F460+CAIV/fBTI930kMJr5cLgSW4N1QpitPjWBNwVNDYev3nJqZLHYZ1ujF
ZSMwobADkwvXIBXaBgmIrXRzuDq05bD+9R9JaXZK2cOO/HMRvWdKRiaCCW6VeTeQLhu4WWbIbjBQ
l6TZpT8Ez1R1IlAhhAlp4II7yrlduFiP/s02ztpc7wiA0DBMMdC9nu5M1gNfklsx3IbWGxIrGduN
wO1tiJPdrh7jhLoxqmiFKPISI1BKrM3sey8KiTkkbRcabMg4jrZUrMvuO2DmzWBXffmBRVtJRsvA
0Qtz8XRkHefSmq2pwDThuorFrQhAMl80D/QAkr+1jH5+wkFWMDlbQQMJwSpMgO6WbZIny3+efFhE
NYAGOFG/nd6kFMeV54XsHJ5Oz9tiIJgA3frzOEr1/V1H3w24M7pphLO5a+33pQaCXnpqw1/H+u4F
bkDaOqTlBxOiG1FLSV9nFFSPCf/o+yE4om6ryIPR7kZng2cmPyAJW5Fpm32yfwkpeWmTa2xL66BE
CNzoO7ryfrr3vq7IYneBi/QsC3Rk8GCsLtQPyMnDgdiaLorg45v3mq7O+xy7UJrZuTbkfLRrsyq+
TeSoAXeuJGbEkAaMhjZmjprQTMv2/ZxKtcFxgfhx1sFubcdqXTs+PedIFtVUN01f4m/rObZYSlhc
RJQ+9P16+qgIWGAa919Feg4p+3pd9Npl9qe6qexa+KGL1xdpb3JWjvosa/DeoShehpPMz+Ksf2/9
gQKFRIx5Tz0LzeUCUlyh1WjJmDavplBOyMwHdKKbEauMs4YNwyUmUlyPyeNTJ0LjI2EclUSqNDG3
ksfpDMmPlTxrV9SPAfWncIwF6zMzbmJwLTnaIC9626doVFJg8gfZEO8v3btyAxmmLJ1xS7k3UeYo
W6AfpV4PaXIEYswKQgQXZR5r3IIVcRfrOWVFG0JJpSv2PZSZI7FY6mZ/DEbmaRpJ8KeHHUzSVG0o
Bpc+DtOACDbogLCCcPCNKiqYw83PLZJVrRlYKCLIQ+nLCWVpeRxdrvQxl83dYg+Ra9oG8P5pkuvq
3iJ2gefyGw6m6pTbddpiYNYkg6dbeeK1SwCLBimHyJPK27M57v7oOb0THVW3dd8gGZaeFoVemuOg
6BvfbGCzK5K+hjZnkwhZleWL+3ZHaZKbD5gIcg8q9jbsuttQ4NTlWRSEgpsWcOrQ+OI2tZqIMEzp
ru+nayHlfkPW2r7AY1WhhaewKZVWf1zyfZrgN95TyXuIsKkBUK2BSUMheWgWztjVb4tyJBSDFzp8
4xF+jWM2ATAmWLwv1aB/W5v18zXStyqksOeYyc3XBOD7SaWgILqDd5nxqexr3by8W5XjCQk5VElW
8EeSt7+vq/MKF3tvTzrw2FaZQ58EIzq5v6xmCGDknco9z7jAX/RKEesb3jI//x/gJteWMq3O9dKt
zbVHb8VcMgNy84cG41qhPeAGFnJ6gZfHpMbi1Wkyq+Ip+lmreihtS7lYz4g/HiVKUt8ajEPBtYEu
T6rMQBUUDtOuhWffNIlTGmnhPLHTyM/arovAJA/joLbJu8e/+Nwt16GXIA8RZ7xDW82fRQi1Fpns
mtq5SsLu64qYdlORGq8xbU9FK5HQzmfSPwKLCMX403iItrIILhPuRilLUH0UxIuGqd+3T8LCyYuk
Bq0/kFelezBCpxxHKUJ8Q7QPOc6q0ZfjpU9ypyxWTh2qF9A8E7C/sM0wRhftIEWY8qmCXvlC3u02
AAXk5+adHUXHnjZkIdDjUDL4cBsil4HB/g323LS9FkXXnbONUUnyi3LHt7Cq1P2UUJGTRPLdggyl
JcnTTYe2hjrqDE4K5SQ8Op2oaaY940yqbWlEZh/ikmALZcaiDxhMIwrXRFpe1wF3ybeN0Xd5005g
RkJr/Vmtq+ebyZTRErXS4GTgYRd9HUyHn4v1jaqej29ZPWVUw/zK5IpUrRhfL7XCYQj19btKG5r8
HoEbVdezcOfcyjRUnoZIl5cKajYnT+Sus9ddppMNwBGM8XTElDqrmf/duF0ZxZyA9bDhB3+ozROd
cXAJHoMkQX8lftDG14aK2uszDIViXFQsYzYdiYaBgshnWeY7T75BpQt4yBBl+5cfY5yxmDpKmcUE
i+wr0aVDIcP5W3lJ+J7npt/EM1xeuP42eCoMHtYOwgRZTqjNz7TSmPqZgDYZKEx56UCDDGnq800S
9cOOjn8DqhkLEW4PduQAlRM4UVF+NqQcyBu5Z+xY3jFwTtrCWnOvVOgosbSs9RtSHB8gvDIZR4hb
gg+K/54BehueKiKaKP1U0+BYudV2Wai7kjdohiAsP2LJPN9NZjJdET7coTuVa5JkzyIWXUZ5fr5+
SFzH0fxEXovUZ7C8zp/NaYN0S+WR89kJFtJKbqC77VBMZGXcy2mUjWK3vXua3ilegJxPVpZ562uV
TxxgsBbv2fib/QeTU/6qB7mF4G9K2vDqqeLbCzluksFN9NsqLbQjyIfGyeVLXIFptRU5L3rN9uUl
Ikw5jg35OZymWLeBQCa/houzAqpajL4QLtJYLOAqoj/8C//siyjL7sD0D9Zo8WHVu+YHTGFHp5k6
nluDtQDZa+h18YSVm6KAMbjdMfRISy7iMjPxSvirpxWkFAtun6MuH7AclnHF83TKFBjH9YUZumFG
yAlI/m7PHEkwBv1L3KK7SAwIAO1G6p4oK76aQ+lrr0jrU+yrG0VVG5EUCwiHaUwBmnTl837NLkyN
1cmbi2270KQP3/17o5/rdHJoTCJdLRAip99noQantgasPZl/u3A/rlSTzjX4T/37xBjU0dcURZ/I
L+DnbuDicGNgjJZcLzW9h33IrxJVDUEGyjJZaJZwZDFReSecqePC+9bSteQFM8epoOGbcAO8lnGI
uBkv3hk5hSFy/BVI0vXYWD1GmuE+IUXVBdOG9AkoqXKGPT4lZRGDdOCY6HMDY2j0cLB+T6QkVum6
i9lQASfUcHFm+HsdwksYQ91YKG3fDGDZJytHJfNZt53U1DM4O+VhAyxYQyi7wcGZ9KG/AcyTrJvD
dW7xv5v1RSkuEifdZhdqhWEhddLmHc+Ercm/5XlBRay64qfKIw4gJat6N2OFXNSjDkzIon6wfiNC
1E4+s9I1nmA0AdkVTtklmQgoDmD8uLqJbeARIiJvEC2unX48tc/KDejOVz6RiX7tKVV1Bo5C7b/t
ylIYD86AN8vBINKtPeUyfHIfF8q3JhYPjwEkhkpfXg3tyJrhPY73Q3xk9RFuf+X/UQCUVhkmfM58
TVDORNc3j+8aDNM/lIq1B76JDlFpyVcbFwVG/SIJfoLJVgTm3IO9vyQdPalx1IoOVIe62pmGvPHI
Wf6XEnKdHsGGE+iuoB3W1kLxV7G3ugKOeNhHUVrE6+ZJ2NHNi+DriVxVufYLGytnjTgiKZ1y6f4j
/aponFd+uPPFP2sWHLo3BJK3TkH9UIrxKMu3PPUhKMo+fj4TQZeqY///h4T2G2asqPPoGEN2ijWM
8Uu8Uc72hzNiBYU5DUgN52DclUnC2cdfUqyQMaf2iA3wCyiKHEfki0XWqulIXU0ZxzQLiIEZsePV
q1qwipezcTZ69gYG2zcce+Q44rNIvBHgilGS8It02F2aCKrIk/g3KZwAA/BcXluXpFE00zf6n/Pk
QX9AQAmkJIMFCiO9nSFU5+29WZ3BFAyb0pyCR0N9pD4M38tCXgY+HuQJpWJaAd5Bk9Cc/Rdx8Iz7
wF25RjvQTDA0TrOvbkzpabngGG92Da5SEt+LtKOlWt8Qcqf+XYfB/2frj72dHzPT0I6IYl6YN90x
YvEWABeshDJIWKft+XZfxGCAPkURrFLJUfUiMdWcGAfDZyDZabgLJ96wPbvg9gqzORRnF+PAQ9zf
3fFIBkm8eoEm9k0NXjqPnINhWku/IvUf/SHtbv6Gzo6GUNgQkaOfgQpjJVP+cnGCIdnXez4DqCU7
SeNH637nbDdXhrU6oooDhLOVZFxiGGQh1ER3LSViGE6A5owlV6/8SUYqe4giexoFalOPk70sRq97
9hmYqwhmCoeVzQAflekuAoBr5aCvIxQKtlmJtK5PKTSbUNxstLRc3l+ysCwN6WtyG5Z8zLaBPG+I
ywI2/zVpzEin5Hdgtxzo7hlxy9hEWoDWsXpCgGbPkiOxTPXY1jO6mY0X601hZx17YJ9aCD9unKYL
uBuSdBsxYYWM0HTFaXDEaJ/nUwJCjnZjBXQIuU7vnYtARw/lgek7xMOVq51QIgNWltyX5YxeC1UH
es2dDmZDwOStsikgB7tDqbYEA1CTbpcR/PpI+Xl7+OrbgUzZf/DvSlN6GbzDhgMZhXvn+ZlzNq0q
JXJ17VhLYvIbDGhz/RSCAEim7ISxky0IqE97PqDI17zmVAwgEQQywLaUYz+YWJuccZX779uvIjVO
7W/52e8A6hx6SVqF9l7KP8TP8pNhuCRYljWGTrFXBkgS8UCL1GhTLIoYqm2oIIVUtjYk9ddGsG9S
QD8rae3SIybV9mPWLK2uZdh292e4C+xmuS8FFjs3RSjjKgAWQY+HREYYQVRnZgZB5/hK/5zdWF8+
ECICVrLPRihmDoY1AFne/i9ASDb5rksOjTLIxugozj2jwoK2XPNC09MzLn9QU8QJtzBxkFSbisv8
LNMYOUUjC8CT2ly7l9+mS/3txaMwK7nOARv/tj3czftn49vE/cocM+H0l82XMr7W3Ky2fRNvExJS
mrrDx82MsIjiZnSEVpUAHeIUgxTrmb/tKpWb5s1IMWlhX2/SZaIxu52b7UAF68OihY8U+X4MhtZm
cP2AtFEDKojRdxXZfhMEp09UaB1z7Rnfv7SDpIWL2j6nY+etOqfEb0L2nyjHG+bP4DT0L2qGcK5Y
Y/OHTz5ZItjewMdxYa6VLLWQn05Zab9hOGoUnk64Cka+xsjQaK5NVsFQZ7wafjw8ocY+vWA6Sa7q
6/bfp6RG8DoqAP8qy24xnTH5tstQt4C6LsF1cRuTDwDXw1DGdW/87MDVdVkzEvH2Y6Oguqm1C6Q7
IQcdT7bS2TBgcMBk5hELTVTok5ILIt03BXhtuovHmWpWyJh3GDPnGgmFTJK428vy2K5vcoOwfX8E
UAWuQFdinHW92Gh2TacGqJDj33G08zRx2/VtccD5IV6VqGLiKPmN043IysJAEC6Ivn0juWuFyd7o
8/jtyPIrs4N/piSvTS+m1hvBNQYDcyZf1mvqU0pajOG+XKm9EqXagLFbyc974XJ2LYEt55ulvisN
FPE2U5oCC9/Z+uDybGWubtiZ3Ks2iFcq0eJlznCwQy8XT67a0YYJSr6J4LhETWmUB4IU3o8l6Ifh
kCnMB8bhdmTa5zPBiWG/qh/nDYREJLwPqcD5R0tsnnQn9N5fRAxUtY5UGgGLTLdhbY6AhcOIilOl
4azviHGFd9qErID9dU7yxndkqsg3Sfo/ThphWNr312Y2LeBEqS+MWgvE1wAcYmVlMt24lV1Dzwa/
KtM9WPDqtqQz6Rjja1j/ZAvmaq+BG57QAhfILnCs4qA+QDTWn+qZPEzqEOvEC40TVYVwGxQZxBQo
N2uJF+HpgED/7wLEPc+92nr/ACjfuWwvFXje1RE/XDLBncO23TuaJ6CI+oL7K6MdplnMQUr/Gpzx
TDv5tMHP+OgORv3oU90Mda9Sm2S9Q+Hp4AmU/kpDKIEgm9yaoxUeRpZz9fr04XZKE6oWUlkVZ0v5
2TSBmUjLxPgYzgOdQbs0s7E6sGfYCiVpW0S2LXqAk3GzUwHixLBESvD3UrdAp7bb2Oj4WG6pMk4m
3rqshKpn8p3lh63iRp1pIjSE+3CAIXFkNNu4P58cUP0OX4MFFZ4kVL20cQsSwHjYzq1WLBvbLMwf
r42vt5Ss7U9/En8IGjFFKB1wFIeGrVxFn6ZrV1kpQkdAuTIs+CFw4j985OS5/CG5C8xCdIki60sJ
sbdy5DFmoa+1iX8LY0ARtRB4oDtV3UR8z1qrmC34f9hAI8fwjOxh5lgB5fjBVapOFbLoRrsZGUpY
4C76dX1ne47X6PA8mNfL2fKkZZKerwWfuA1uNNBXcziBJGqn3WyRWh8kLdv5AxcQ2AZSCTKB75Tb
hBnu3AtEv7aNbgEGp/LJpuhBhX7LmeK6VXQQSHrKhjoSNu1hmGVn48f0II/4JU7WZwDWitMspQpd
wc969a3GkD6II0R36ufk2b0GKYCEviG/YPI9tvvNUHBiqXQLmZDvBHquJFojOd6W3IH3foEx6zXP
PMQDO0+KZQJParH+of4qgm/yVi4Wa2qkO7A0qukm7SClo3MJEpzQUmftSumJ/EH4Lm7c4oSNFyNZ
0MOYrg2uFngirvRe4D8CwnWxeIMg2c2LhFU3yk7Ewytb0bsGvsx8EHCeGI9kNo19nbBoQApAZbax
YwfmdFREH+0uXSOl0DHcqiQN0pLnOzsX60ppoXxcu7sHvFJCmbELkgdSSl9Er31bQAajqkH+IkWF
SU3NHVs8L7hU2MF2FcAQbmDQSvsS9Spr+NmDjpSsq6sMQzQmkqJoDDa6RD8gtdloygyUBulukdSu
H0nmJzO+s/STEH2Jr282bqhyJ5Wps8kVOUySqlpwPiNjs41x5nrekF5uSN9HiVW38PwYeoSbguav
VHKBvZOFA5k7ITCAsxIEmsGcbXDJ3VrOjVNW6PyXKZwnFl2kF7RLywr7hMmV5RFkWJFa+e4r0b83
BWBiqd1O7CyXotcOSMJrBGWo76H9JQrTZZA8i91bEZjKHr6mTbdhRRUJ4Efas0u5EkwUlHtHTJZJ
opfHY3aOakGuTgcemVw0Yq3YjM1xo2MSrPCCmzyamdDSRn176/ESIGYyLBWNSJNU1masL/k0M+Yj
pxU+wO2+Qrm/oS6ynvqlVkyiZZWEQYwoPHucFk7LS1uio5Ut8B4ziP78Uh+60j3kOXCsUC/wUVFt
ha9fQ1Hoa9/Wo1FLgKZmJ4Nczidx8S7tvTooqEH+zp6/2xUuiUYzfuPhSIxddwj5u1j4OQIVgjJq
7fvLR/Mcto29T8DsQ+izddNYWMbtamKtUEK9PYOWPjpIUVrv+OpEWLos1kl9wOybauiMgwNy99ly
06FAQ4g4tPFpWb+NGxUfIDRQwGpjIR80zaIMYkiImPm2lmvgURs+t+VNqlMna5w2EVlMJVqY8jAl
/tqcX/uy4ism8/+MEyqBvfXCp6AjEGB8UFBgW0BlRuZySolFVSgAfRUK3jUpfn2FAV3ZX8QvIpzX
S/cd4k4MjX0Ov2yX39D/SOulCWrA7gNWydUSylAbMUCrzRMUEInLpTUF6ud+cHAkoAPqkoXp1thO
2a4Iam55vEZ2q+v3h1ebAI7tr6HlB1rlUgZB4sFxK8jwyLsjBfVdAM/HfcyPw3LjZcH4vHcFxkRQ
zlf16jtBJlT+xwvY9anydjjuQVaeTAgBq/zUlAPU3OkXXp1WiPsYZJhcRXs3JKS+8fbdZ4wUESDp
Pc067KNJcwSc+52V+qUW/q7JMmcXoQ2CmEVqAG4LBeR2zf9N1aDl+l5ZTTzMOP2KUAHUbSisDICz
RjYcRrP4EJ50dT4LHij9qxmF1PqOimY7dBC68WtX+DRxnM6nyqjt63dslZll46xCfOLyQEXhzFAm
3PhuPLsMX0u5WZKUxiijIYDJkDjhpIAqL9xXoBjoDyYyKTANV7Mf5xI9vj7uBOH/d0FHFl5nL1m3
bshBJMXvbnuh8HV/sT2F/TGve+JhEdZ4SY1E/zuOcD29Jvfoz0gELYvbBR77cMwECKpXw0vSd1CT
jqh6tZ3an13urPoAclMmg2MfpdLefaXKeAfLZFF8pm+vbHioghdWx/+05c0T7HirLFyF4yZfVtm9
FUWvOmVKLpVuDeStSJ8v1Xqr/ZJppjzJaRVtVcYF/Jz/9FBDiN8SH0CH7p44hWszzdo/3Sd5oaK/
sSJX2ETtDN/atugjuavseUDyXf6moLHd2LXAO6GDIRKQ5llQOJrs6wa3cJDKtKNo0A+JL/RKS6wY
DW0BO8wBqHnrZqmaD5cTTiRyyPYuejV6A4NvT3RRf5IZI54WIjMgc9xs+sPmUY0a2kY9iaM+AHTv
xuUZBO7PNqMmsk8DZE1u+LBt9oSDlWnLL9+bDJ3kG0xDGVkG3rLsBXXXg3wUNKIII775pQX8PcC1
m7uxqVewQ8Fc6chlSeY7Qm/U49DT5KgFxY57jCf6cTg5Ss/TjrsVPiguM9zNqf9kLPH57tNyq/UA
ljYp+z2Z6xeVg1aq8x/sNTj0YY8H7KhhaE5Uu06ny41CGFpGscCB9eSSM9clc7Lk9i5hCCEAdnD6
/VuhbYLs84FQ3vVvWvc8iMLiLDo+RSB4Jkl4KoZFai3E+hTJ0RFNShihqoqoMa/Z/y20gAimrYKr
55csBY1E+U4DxSNoZzD/LzFdR2BjvVo0u2TbQOeVHnE0TZRzomO160D1HuwCou7OULQE24F2me3j
s0Xx3/9zaGCkZWxJgHXFBdEjAYpYedIHKL3kr94orLAT8uJ49GM40PiMYqkAGxmoUQurRhgyAWyO
6rJYCy1fnxv+jdMP5WWpMgoF8OgCBB1QZiONklFtaSCg21j0QExdVa/FrveYy20J2+7aPWn6IiKf
VqWvJ+Yv66pSL9ag/C9SVc7reYs8uT5vd/nUKqYwHSjwa4ua7AHyjOukCIMscHAtKQO6YRw83qPg
2+Kcd0sXAwcXfp+dSbHqqseG5LHD8xY8CfJYTbdQas7nTEuTII1adljl/9Xnt8pKUie7sp18rKQi
7Z1EXJAEjX/fgYZSesNp1xKmihVkpoXeq9jDoSRnUx38OGFQJkMsDSm0pKpOQhc7VQWpALIcXQeV
UPNGCenoiunQqbSrvkPAWDEZmFbwujqqIqS9PZct7FkmdrdcZ/bu5cKB7UzdrfmSd/4ZdG1seYkR
wwfUQOBjRNMNt2hl1QSK+UZd2HG1Oaf1LyatCVVZgEeNjBTHPPLA//YbDjJRjRx2w1mZqdUXI5U3
mAiiTsHIbBh7h3cjbmJgn5aDkK3/UDVaFwNtIowzduyfx2ZOZCJrrWjeArTLL5hdrHyMmbJcLCCX
qiNYZcF06kdWfUSR/eaWAzRBTih+x4G8TGc0VXckKLEP4xto+KwHPDAuI+HAAm61RTY1dIqChxJ4
sdMdWLUFeOPDQce9H0Rn20vSuN1mwRkOCl/v4F0XSh4+78Mv6VqpV79DgPjMn9uSf+/dfcCdGlGv
AiovFFVHwOzSSUxCoeO5A8oPP8q9Xh1Y6KMXTbrSy5aNPt6ACSFjsphCNHOLieC+xHmob1xwtekr
nBQE8eZAe9HUNVxuUyhRGTgxl8REfZGnXThrEq+wZdEylK4/R749dSBT25xaZL4FcdD9Z/AC5qpT
ZnC3bImWr0NjQOqLGEdEVO3CEN9SvNPxtCF6THaILNXW1t7mhNfR/rxH19kjC/YH90yuBCP2VTjk
0b26MqA5NdYOyUxaAl+9B9vOXBovbbsJjQl1SSMh3ABjLYG21RWRMtE1gWR1ieCyhAQ6t6k8FZ5F
Vu8eR7+lzWprmVlxsHJyw1uFCUojO2eJhf6lBEVffwN0eKqJ8qgOcIzcaZhx1wFJBZ8qlS62CikA
WOKdUrd70q6QVs7wBreKvk5b072W5oB8oMi0GgmphYPUcLGkrxqUVLKbI/Jemf8K26k5nQmWhQLH
PUilllWX3XGJA+RN1HW61bDGQ4fSoplZICZO64yd7KEYJrNyjJpCfc7LsbbkKljfkwGiibc8TqWW
1AtmhWwgWdoYC95uwNCNwNoMn5md2IhtXSU6f83KBFfIzM0HND8vVlQWH3m4PUQmd2n565KovIPB
MTVV3ijP5aOth18SttLf2o6Tyu13OzsXFCS1QyFn4PEBIwV1KWos38Fx9owXDvpAZGpMdogVYcM9
x75fpS3FtbbbbaByW/ZDudDKGtruSsCz/tiw7c/RcEKK0hq11VC6/AEyYNN21m3pFZ9qPa2JtiFl
9FJlgHzjzUtrFJONKFL+4rG3qHI33n0GRG5aZ722DqnqaEzexT49NKLd8YZPkLfNiKTA1DkTXIHc
qjFmWlA4iCk2rAvUWlNANh2VP7kRiz24qoDVBoiVtHBOruTbWfnsmkoa+qrbW7hzYZsxjGW6nRzk
XEr3uh+9XsQUUaMQNtbxkFR2fTgckojPNj2RQgq2MPjoOw6fW1HPvpn54HViXFOFesTR/l+Ugy5R
bQkJTS5j0WbvKTEFZQgQn1EU6qFDwO8OCQganLAI6caaV8/OjcUBXlxcUGeVQknqQ4Z9aZUvlSXu
In/oRcW5xrqENX6wwaa4ldT7MePhcjPQH588nCERu0Tv+kglUJ3gKxpenZ17TK1E2SaA6ndx0WTf
ReRBnY7jv98u9esFTxJ81+oUlCYKhjyVe3LKrro44rjR71p/8xUmMmy8iGI2QAmI5LoMzNl6+BUw
/0ljXMq8no2z4+x8Fa6NkmOiyVWylh/RuGGXI8en/VyC0KrpHFv+ocK6/QIZw55yy3RHgU8oIqcd
z21/q7MtAoo8lAqYzHxlcpIFczpm/X76wsNtNWZhLZsZJFRaI2EjTKOiTm8nIbWnrvvegI9Y5Lws
qZG9azvw2Uc5Y/qFlTbz38M8GbwiPFlu1pxHhyKu06r7DfSEJK9qn1sDRvgC5ZrRNkfkfTtKIl9l
O3dzY9nx8tzo4YDa4b8o7yJfp1D/CPUfoHgObk6OqVuIQ5rnVGpRbhNKKZtk5fBFAW8AltGCXwNC
zd2PqB0OoQRFqdstNHuoCxcnJ05s5VDBzovu3Lcag7SFGcnxPYUAd5nycXPCrlPGi1b+3wW+0RT4
U0AMj+9YIBRrqb4h9CQ17AjBhKvxsowEmFDUIpelDF/AD5Bs/t/w1r91Flb+oBSjPBRo+pL4YQs5
jH2rBzGnBGh3p2yMelCm2vWQiDqEBhJC5IlNsGadCQEKc6DWZ0GYKxJfaLcZsBTkm9xPA2dVEHjJ
dMIWJ+LovzonO5kdPArDCDx0or5aP44KX5Bhq4mYXkHCYiv/jbwKRKg+n9n+YK/MMT2QdZLSmYhb
MnxbWo88aXOyIhTbdZ/MpdPRFw8zSRm71yBt8i3O/XhRTDEAZ1Xy/J/qK0uWRS1/WnuyKSjDpyDO
0tr4NoeRy15N3YE6k7zwny8rtnUX19n0k6exxAR1rDInS9QGy+VovY4tXITTVczz/C6Oecl2eJeX
ksZ3RcjVMGkdcmsGOwbNqjNbOrxpmA7rwReshuHJeH6eUM43PZJH2dm29s7Iv3wbAgRgZSvIp3Lq
fyyz99uUP7wZ3BjikG2jtUswarOiLFDtWaEZAoLZyLzhX40e1izZucYl5SnITqWmpS38LKD6Efc+
i7PPsnV4nzSARVKhhaL2kn/xPvdEm8DqfCEkqEBLPPErrS3VDS8ADNrOaPEHxwaEAacpGowL3cbZ
bQOoge3X7V75gHUAugKmQz2iWIbOUUsVlR0uHh1izHufWwt86UDp9NlQkLZ5IlkSZZiJYS+VV+fy
WER85xxzjHi6XWDTmpfOzPTztVIhUXCpo0YKy2c2X3mHNA04MmCy9bCSKVwlitIB5748VYWpggDu
fo7/+a/CibQhAUVsIh9/Zi7UBFPrplBbkOlhQ1JWzzddXU0cDtDjnbrFSmGoATjmtcsQbAdG7lgb
EI2uqYFdb8MDTUzpRaJm/SY7yw7ov4ySpaVF0StG6suSib9LQ0YFRm5Nyt4EBE6K1oRFIOug+uKo
XLzKu6+R9mwMN43KaNpZEwAutRYXhQYsd7ut01EkxKQ9O9ZFLiaOjAHw4/5T43mCoGsV02WXMZW2
d6jIwObMbYgrVyKg47UTZfM8BrzXy5zk3L3j4Jqgpgbh0IOfsiSFrPwtoa0YQjXPMZekBnqg+PLq
rrK7fT6KF8hr8PeuYXN5Gg1D4LJo2xzofKtP9Rt/e+ybwJFlFuXssBiM3Vz5lCQGjjoH1hh2sVXk
j7Nxwl6fw6pK/alAB8oQQ42b9biUvSTVoQvPX+YBDzREllkonKYtX+uKqhE4FdS9BJNAJW20f5fq
UiZEN+5ezEUeuR2+RsXJeOmYWmWWWOyittc1VNVOn7VmESja5T/ZhLk3z1O8/09J8dqKz91dvN/e
CYQ+8hYv4D9x91SOlDEvpST2a6Wj2ErYD0mvVA3SeqStIa2AdH5O9zItxjEcoLuSZKtAZggvP2Mk
DRblJeSKynD+rhVSDxotwywR1ZuJ3YGug1O93gEp+KKD02YCVZVv83EFZYzsgP1DR4oAzZGfZVeh
TvQDF3uOtm4F0LTgRs+YXuVF0eScaOle4wrR0pntjs21oiH91vPvW/w7ADY2LJ/cc8reT2hRRZO9
2dVNNnU1EMrQ8ipG7uuROu5Sba7awd06BkgwgBq7SEUDzXaaxxFFZTWw5KUQtpI1l7D8Kmh8RmR3
35Mol99LHQnaOxw3SkBXPq8nDTtaeZqpqE4/xh5KjMuvyR5xGM1/01c37lwKm+2XRK8ALgSfLwVz
KF++0fHo3F3vecpSn38H8bwGynbFIOF1PJnsWAHXtNy7nzgmtmalrsPftPQflOg94+QCSdRQp4KS
PJt3YKXJJ2dgqxVPB88G35+uuMKn/kJmQ+8y9Dlh9nJfpHE0QXsnhMHtdSznc5lVRM5VxL3HPFE3
nbct93msAeG0Gr3FKY4D7pSm5jWYMK/LcSH8P7UOYOTJC5RddXILsTsjT4w80b7sfxQoFzLipBZj
Q2G3LbU5jmV/X0ZSZUN03wArgsigr6rC55QjArpaIFIjCOV6I57Kuqe2JVKYAwn7JpCjgrFvdnuj
dPNbWEg96MDt0xLmt2oNQP+n6Iig8Fyv4Bi9iE6s/bGAwLGNm9oB6KW8AD5rANl91AzpREcnova0
9dr2QD4mFQHIkNb0SGDCoe7UlwQ0W8Nlar0ayChNuDKrTawt+aeJizu0/fYrLO8yh0otZ7gYtzAh
YkmcCIkLUE7v/lB1hsWbW64DgkVk9BG9111It+yMQKpPOj06nOAwiAQRAyxpEKvdyPdsrSiKY3k+
VcU9WDqQyJFK/QOOZZqz91fbCCSkyGDt888VHW4HZLZhEL2zI2Pf0DyGuf2orB+c6sZOwzYSdnJJ
jJtc51nclVKSXCR98CFA3oIXiespHMX/iS/XYOXon83eUcgO1C81BDT2Jnbr11beJqQXZLuZNrqa
JTnp9eZAIipEiWanvJtGX2lduivG4V6SnwLl6d8EuGlw5fDxPrdH6nz3u5N3wSSsov+iXufcz+Pv
7BY5G2/SzXA/QS9SNcQZ5oWwnchz+5wf44I7I9Ucpe9v+eL0pJ0PijGn8X5OMByAXJ65Dhu1IqT4
3BEGcuWgPDoFhtI1W1v2MOxADqcxsJ9pPPFtpkY/xlrQDbNSka1JrAuXoqyxQyHYvyqnBSUKAUrH
3JCtZQRMOyKW9pwRuCMBdlS5ZheoObuQlT7dtxzKwW00cH/XgOkIdy2gDgvRdOh7XLhMJLgO33tc
fVI9cXWtFDCjrjgI/A3jKeY3TUbolFAgoX1MvrXDRI1Cd47zPr6iOMvScJlGG7yEpspDeoodYKLS
MWISpZ0a+O7ggU7YkpixKraNZfv/cZB+JP4uMqJKdQz8okojs3mP7VdxwkVDBxVvax75CvDEV+6W
wveIQ5wQ+zl6NrvLr29E3ISkXexICpauatp3bpbkSUF11/3HQBAUw1hdP/sV7mHxT808K2ZZIr1j
ceN0dSrs0HJgtpJM/erR8s4THC+ggh8K/+/oCrNU0Mn5mZ/jkgSlCycaPDE/1E2KvS8TcuM515nQ
lzf6Xjhvk7BCD/P7W7qCH4boWjhn1zPIC7IsIFfKIR0r2xKZKFxZnqh7dJ0OsK2B45TQVzGbKUbu
V9rBQMam3eo92IiYLpddpU9lXeHwDlZhI8otO+EQW171U52fnKonSUEFVCYLg7oO96BuFnyr5SHE
mPhkvEaS7Kl9s6hMnj7zOHSn3JnL6lkccYabm5DYD8pTbzUKvEfEqHlUu8HmMiUrh82DjuZlO3Ry
/4Sm32sy7v+5jDQG38EJx5cZd58RQH9SM0+MT/n9YZVoUq0p4I5/0XbPuuMtWidDU9L4l1cu4U94
Our/v711Od58Nge8AFkRqhXxh3l7WaVqBZL+OihaAi1YpmYrBZO07OuJC2Zmb9BWLMrPK9p3Qey6
KMnQu6wRuZPDZseYs5ou/yZek9M9sqw6Fi/h7yje4m509nRYE/KHhGhbrvdQAZta5W2L6JPpfujh
twW4bXXoTd4u4OunA1IWcloz5YisoCqwSj6pVd7F2/TV8/l81o+y5bXH62l95uadRHB/YISRIKYD
gd/krYPgS9q5iJRENBZbsle8gFLATdk9RN2Aw/sIIxdTJBjU2bU9LLZtTtNvo4poZC3pEJotrL4M
bPfNd5bEO2D32bdz250bSEnBdHeFevm0Etstbo53bO9zpRn9AkB2XdltO++WoW6nOlkisY4xHgja
4tbNmzkUA0z/Y0oRfArY+s7JEWQUWgFIDyuGkWCnraWHGxxm4vOxsORPrMvNl89Ct68hGi7JINb8
ImPM5nLMNM0rSZt7BXOvpHgN4n1vLdqDT33qwCWmKslJvRYrwS3klVkkRPg32p6aeTJGaynCDBif
xeVjGySpagZqRfIGP8o43Ed4WGt2MTsc5VVZe1//Y069IKoyK7ozXUnw4Iw0BQbgf7d7N1vsIQqS
Nljv8aZlLDPUwSxf2MOAcaJEUZO3GMGrJsjzppfuuFoZ4XE/Kzd7pYKsAdMT9Iwxm8E3b/pH0iEf
1GipSo+drctfCwSKcP5hE7aqB6m6AoAT/56FWArerEPreX+4FDET4pSauJtqpiDPGQCbOdtDwMlR
9BAlrJ0ELOb7XMf3BozIe4OojrIFh4zsS/rZnaOjqBW4CUMF5BwvortoSCd89z6bkNb1A7IFN+fW
yakRz4rldt/qWGeWffYSxj2IO5mvaJiYiv1iKWesRtIsxumFMebY6+wLeHSbLbbCCcKasg9aGApw
S/JSvGD/1ngXmP7m0F+wM/LQ6AhypzApqBvCAt4W3w+qyiHJM6TBMQEh1vK7AYfgashPXZbNW+UG
9Ca+opFVgXqFRL9lK+9wOHIPeb+Bs/WaLaHYbqLolv9F99eT1xpzCVBgFNAOAOu8ixyn/abrF7rD
BIavUj2UiuomIzs6MFE6AMf2I+Ls7Qf0M8dA+11tT5AD7dZrXE5ocVQBEFouU06HJEMraUyImcA6
2TehcHZ69WrguYuSK7RFtlVBfyJ+OXOVIBjw/MwLNdCU25e6pfhOwFwfFHMRP0OmYJzwXxirDBuO
LiivUbNd3CcUhpxc8b0j8RyfOUIruXqN5m2boHQSxj03pTAqDSUrIgEv1V1Ojceex7IqA8d4oRVJ
XI42WYw8DHymHnruc98aEOCvTL0qOuE2JwwJR26qXtNl3pIAKMder+LO7XpTqJwlYISaVlVqKa9x
B1FSFYFAzBVXPicL01YB3s7gSjDxOAzEx9yJSQ92BaZ/M40u+E80/mT3O6Puv3bHZL6QjbXJqexa
eBfc7nM2n7r+3nktTzwEu1g4UjSO2KB2KNkxJN7Gd/PoKllladvs48m0+XfMZiyC58+y6VLRzOwg
ASqzUZD70YytobqJvFFGEU2kddlNZ04S/wtphnn5DzAahw9KNUtmoKNkZqurGPxpY/Nk2Ylx322E
hIjy8xzTDVgtavL02/FrUngTb5pxvFfKwtGZLTNiaGbakoDOaW+PtbSlvKeVnQqglBxOnMDxlI61
FafTKAoLkUv3fK0p+jSjTl0N33UrOEAe95mOr8y19IvAWQBQ+usSrp4u2cekbmSQaKbnxIbLZzI6
/SJoJ6H93QJBDAKixeP2BNSWtDZCUJlEntB3wjBSrAqm0gEWj+vEIyPjl+p6fB2oCrRzW6PUyk4q
j0zDhqhfDldSBk+hWYzMgkfdP3kcUiAU49k6JwLP796PAFvZs62TICMgy9Yvk4Qs6Kj8XmaowG3f
w62w3GvCcNPvus7pn4Vl8Ci5fnADWYMudPEo+BysFdqgHykWiGwBfOQnFgER6AbyDrVNqSCKe4Xx
Uj2ME/Z0p5ILksKIZ+cApLnOVCy46ppSl7KyeTWz2w/AKvVQxaKVHPUOgVveDq0mK+pIMh2wBVwE
Zzn2IIqgKCmQ0EOjlCXmadHqOyE39MRUL63/l/r3tyn8SqNe+Gk7xclsND2cAIPjeEFFk92c+FGX
ypc/I1gW21EH8WfJn902A4V2jp1l098jZVB7sf7BiIV2hj5C8jNX5jwhQMpMRj6d44aoACBM2d2V
Ixci+XXzhpbMZH/UIsoQ11CBSe1GgHvtSFQYKBosMFqETGeBfaM+ICb7aQF26aWkugL8dG71gu/C
bMQfgASF1e83bvSuJAqqxkVub9zfR72CGt/RHzed4GnlUVY5SLJm90yk7z24W4Gz2bXik9sDLkyQ
nqNGX+FyJUhTadL64SxaupMLcvmfE4ygbr0cw7Z5svFTX64qnzpWfS/yKa+Yu0aJUvyYdiFddlFk
f2aaSWt1c2PbdnsPjbA/DQaYox+3Ucm9XWIHGVWPBhZe8qoAh6IG0IxZ2vbpOkyHHAvu0YbbxtR2
Lx+fsd3o7Nqj95wN5v3Uvm20Pl/JaKObEHYVCQCLMBjSy1QP1k+eMTHck/D+sbbbG1Jq+BeOlFXi
tVFBIwTbcPDDX3hem1cxzY2W+mGj76rI3swjTU5tqoAeiSaFMNp8L7OmVlC6MRTVfRbVLeITbn2R
KooHSx1DYHMwPj7rl+YDkywjoe29G5a4zqC3G68vvFv6YY9P2bteiVcDGWFXe7KH8FPKraktMahJ
9k9D6orz1C9Si4N1PbDtOWhGghUYNUmdZSV07GXEAei7J2yXST7uqpHWAPf0y+oBmwEd4QvDevRi
k6wfGDqJR9amd9qOi1cguzDAnmYs9OmXCTsjjlagTF+XORCIhG9noL/PgaQNyPlSICMRXG12G4Ju
k+yMe10NB0dg7qDIb3nzLO8jyroEdf3Qb+9MnTTi4jMwhgdyRS50MsrjeWOCDXY2mxkOPp+OdfVn
U75Bo0U3FH6JO673J7nSAkPm+Hxi0A2a7rFWnFcRY8fbMekreJvXqiI+Phipw4OKkawwLKduvbMc
CfBxYiJPLWJlrjpEE+kfzlJj7l7DhwYtiP6AyMHT+kTd+MFAQLVUxETPOqOlMF6F4ytgccTKvIj3
tKQsV62rD9eWb7BVpotW+cB33/RH9Ckpza93WoDH3pVMiWVZMjolqKi+9zUMYgTtEQllJmgasc1p
1T693CWhxAl7rIUwnGqIKMwG90k/zIDRPtDFLQb99ekATTlpkP8jVVFNUZwahi8xBy1W9cWG3M+v
njPLXeYcoAcAUUc3pcxkBMBNtfKaBtu64pspKfoLlHCIchIzrTT0MdCCeOy1ohrbxI3R8uF/xz87
+HGsx9Jzp3s24SCx30pcb5eVGXmg0xP7IWrT6hSRQcx0DB3ulnVFcp2zpPFQQun7PCDEGE7tgw2N
j3AFiwAn3p5RhZi0ucJu8X8d879PM8T+IBVLhhqjDZHN+6xQFGUX+J+HlcLKxBX9K3KCMPwcklGo
B0t+Mxw2NJ+sbaLm42N2jjx9tN1Iyo/JzjpbFChkJtiZPaCNLNy4ixCC66f2xJ04XWUpoXoFJ+cw
U+nFapUVVv5lMeJRaimp1ZiY+BejSVlJZ+Os05L0PYqYQL6gzZaDPmPjsV49+Sz/LXGgQBQcGelp
ce3PA/C41qj5sTDdFu15EImU0FH9/Nj2dICmITQKB2OmYJkSqGY9r/iLY/r8mXsnU9VtV/vvQSQu
eZMrY5SK+cvCmSUMloxuABiGXForVnmJU61Zjds12BAI3swUDSGyj7WsmqHbO9pmB9lBnTKpku4b
1MW1y4ChdwSAMUts8NIzf2rCcttNb2v13PutTe05vHRen8XM8vCvFN4QV5bDvtAVw8iTZULt42bR
v+C2YnEXXdHBcQba66IOm6obKsYWs3WYUt+0cb7EGgATx0LVnSk4OBycAXEGlZ3qAFI3PJz1Z69S
UK8VplULI1vvXCrLVJhY8ZFctrhKkm0qgoDPX6p2bOHljw5bIrilEuo9KXMkaDIeniXDcVu0PW0u
XmfFX9UDS3gtRZ3B6bLuwFtKs+BLsb84bVH9e9fThbaiBw+TqBUGzOSxdxYIZzueg3nXx5u7dYLE
S+xPpBNIh0oKkpX+7xYMVkKbxxt3AG9AwfHdCAg+RPqXtAbDk+SsxzzlLHbT0Zc9lo6LhTWuFDNk
0O1khWA+q0Kgxs7gK6wg2CdQa2/tyEK97Tq0/JrV8ndM7vwbuXS42DFt6EPzxHzFWw8k0jDCc98Y
IFcN++44dxKVmkql346TK5jINhE6qji2rgjTb+EuY9pRQ1S015noB/DBhx8Ef+cGPM5jpNyfpyHU
cEoras/yCYg6nlYQKdrvJlOYZkLUxgPzD/KulmzN9tHo7lfsug+CGBx+Pth72f2PRwBLfMekrQ4E
osKUy6L+TO2nv2QkPcRTw+uMWAVLL3hgXuwoRuhEzveSkc3CIJKaI99XotiG1PwxP3xX24C68p68
zFKlddQQrtMsf61swQ1oKq/5IVpd+AMfdCQoSbdZkET0eH7u6y+s/BMosIKQS4iSN85KokMe4iOP
DN1HhLaIl0neSIiBopLw9tDrS9k5VoVwDtCMAdCPxmbnwTimfhuhNqNLOLgQdTr+Xw3lpTYoQ7Ec
fWILQntQv+w68wrS/dmls28pU0q3fqgyI6c/YHxsu5Iaq2tQxmdWoR/1/kgeZIVZt835yxitdKug
FCD7q5N3ahl2rx4BUx09p0NAhCkl6k0xSoftNQw2Yzr9jEpkB7vvoMBKJHY+JPdPznB65KtKQbK1
2nt4I3nUJxsRaFvBzCjQbbuvV6RZRC2IpD3H15JYXvb/A9CqNDST22E4jzUiwojCpquBZiT+U5vt
hXNsvDB5dMv2NHagwkJ+cevnJYY/Gh+6LlCMCKpGomaNM1QrDNMlo8gsjBvJ9J6XhrbNlc2OhtM4
TFnxmCDfuVXwBKkZVR96XaxsUgFq3cKaJP9cvx0o+YWhVBvtZAm/YsV2NJ0GyMjNMbzWGUUNB+CD
QaVQkOvRy2Wg5QDqX0y+XRwpW7lCtqHEZtPT/JBH1VvB/v46OFvBABjmjMpc6IKgT9BRPemlVZyj
MW4HxSe+If1GJ5ptoh24QNl0WtGWY22lusof5oz19Ts/8rVHNZtT8vgYtnPYjfMiPPVgAo8/K8Cp
IkM2rL4wVj6lJYujo5iGQKoLUWH2AO+uQQfbEyNpLe/5TBcqVEcLaxPX41/ITlz+ZIq4pGXfykwS
M3osCzvTqbczNlFIL1RVDYNj+P9UNvWYNpmx1ms/tdIH8j2WYQYcPFwNba3g+JYjNswiTHHJw6BO
Wz1LBNPP7wR2E8hwte9k6SLGRq80rKbFD1oRaGG6V8F4QpVWf7SqCgsWm3qXv11RonhrEaQVWjuN
Kuvd5iv/Cfe2znCkZFY2yj74jSun+cP3iFRSD+Ad/f0+30zkvsRNByZfm3SK51iwAmR+Fs4Rkpxc
O9g5dtji/N5EGVn8zS7YCh4ra+kqwF9JEMd0shZsvHA66mFe2VTPHYhV46E4zpUp6/kqq8N0gCQr
8z/M5coougTYmmkRg0Oau4X+ZONKtUJzAQHhSnbO8wuqouEigLrqtbTLJAr4bcsaVlHVyHn1v0p9
XqFHkLQl8Scsrzi8lrCpjnCbRzwnPD52COIDvjBG8Lh6f87o0EVnxR4DR1on6rvjqRLZ1xBiIn3d
g+BXOkvYgxuSldLDk0fMrmML5V328CNU9dXBqtfh4Vr9Cn72lkj97D/H0lSV5qHlR/DascIL+Krk
zOAbO2DBmXJ7rZg7O5BbKzNY3iT8GoVVx7KomDux/9j3bMJkdUU1gqFWAQzSo2NYXQtxCqpjs9Ha
l7FRtEK62DN7GAtbJUE+xx9+CnYD/9hdRm7mVJ6d20DdSfWF/O+RCtkuUNxht17zY+6Rxb7IMPa7
N7MMyioBTBiN4QKDef5b28w/fZJ8i4aRGe9QUZquGH1g2oCcTywolBNzDXoLrMG4IfCf0vN++xQZ
BbX6PF2l2OozSnjEJJx0ZDwStDJEOkmqZjvQP5DL3wJn60rF1hqSnmmJaKaChHejiQLwOltklpwy
qgRV9DA5MohsqQLkWt77mX4NlhuFogK8oM232/ij61GN5YE+bXxxmxAlTqYyEgj4MTP79kMEmgwR
1ANCKGiHX8KZI2iXUwJ8BDTH/toVoWP1wSsf2d29UfKj9yuAcWV2O6AgqawT/cSF/VGXIS3NX72k
4IDKsT2Mxn55xxCwLmXz3nozFc6G3aIJSZRMfwhYPOjzPr+2pI5K6DkH5ZM01usitcELwlEOapg/
O3NOlIpn/ZT72wUylGyuUMGGcaYNT1AA1GWFUb20M5ULHqySuvzodotb+o6ASJdTCBR2HIcoamhT
e/VSIG/5d/+CVg7KCkqQaKWQmDYgp5vy+WOaYLiEQpRUZdkYHtV9Lp7xaMZ8ZuPDzt/i4lULcFH2
IQuz5KmldOToVLO3RzW92uydaCSWTDyvlBmGl1u7Z7XJubFKE+lfL+W5V21QkSA9ZtEUG3AO+Kbl
6IqXIAVJF4CCRptqpEADRjJMkW9KzwdM/YmzmkGhF7Ismqcl2YpA2TsZnYa4I8v3aHcO+okfEIf6
Sbtm1bIKY3FUksU5P0L5c589aXb2dFLDVYO7V8bA9ne6NFJWuXTlyX7fXRYraj3FoK9mm8ajUlHc
uPuuo1/O3s0kN2WHNbkGn6aziYwz/dM7q3H6Sw7zO8vKCg8Uo2gqCfOMhLRHH0zA/1YkYQKjB1d6
VYFlPu0eCM3h5EuJ284bvcNaVnjE7EO3UMxhdsocCQefBcHxU0+ifBDcTXirq3IISVGpB2i8rYEC
a+KrUXY4csH8h8xFLgmJ83zDTG2od/J6qz138XI4YrvqAm16gRuq3K4RsXdENBKiolMpHdIUKaG4
8OtkctAHiqwikkmSuqsPaz25GYcesf3q+/rDo0d+IPJa1sJ3MuGHymCLUQtc0JRtaRV4SrAdoNP4
hzldK7b+WAD/EzgJJ7DQqGmUql6veoYxgHwpWm9CjGuO938hhiJC4hhBbXqZQTl60W+0As407awU
GKxlLF+oHMGqBPsMEluUZEwfrnyL8cLLzFt9Gx/oflgHO5oWTIKY+KHnajNzcOV/JKnPGN22K1ym
jnGE5j/gAvVCrjHpzoo2/pdHv56Vf5fWg5thuw0cSfuVU5Q0X6WVaJhmWRphWkCNL8d+l4tHaO3C
j5CvZoHqfAcWez14kgCOSoDCoTT5TOCX7BihfmwAkHfIhWyzI4sAVzmgfvDGbzzH+0mbgofQAGrW
uIJ1h6ZlBkDTCKm+mGcjFFsHchkJumRsO206dPoVdoOULurLnHOKh/lx1AXzkTyAOMFnaMSJ6D6i
HQq8BDTRS7IQ4bCnRJcytmsbHNWet7DF6yd3XEAsrjG19QpP50LkkuwGp7Jx5P9Io2ckHAJnbyMo
T4ygUu+qJ5dgi+v+QSD7avtk2hRl97nSWdZhmlOqDVDVpkHikw7Ga8uNQZZEmuRe0OtDMaAwCF6P
NTkLz1FWtiGKgLTv36UJFkCe+31O8TrYEWm21Vr3PnDw06yH09GHkclwwgOG54b4EvupgmZ4jVeM
KUkvacCamcwIN+oZIT++AmlrL3ItlIEoE/5ermzjrUwevDE0hkMaisbORZJ/TruJyR4Pj4eJWrBO
WZD+PBPP+YTkIptZ2P2eMBJ//Va2JCrJp8QyLsmVvO1Aa6OpSKGBmxh1DWUi0TXUkjphcMCwWOW3
lm4eGbfd3gqwdTGGWIAj54g55kj/28tlOfOFTge59w3vInhYWmmY8sIPWPDdaWH4tVo0zloiB3/O
RRS+dcqrdBAWfGeKy9WJcKt57a4d7fyuREDbdgGeIZRUeGre/zghlfM8hB4qdbdQ30IVeIHh48w5
iRHsEa4W0n87lQ3qO3L8rrFGcznYCUTM5B/nbV5E7vtJu0wPIhrB+v9fAakZLEpKpfxg8anEjsy4
B6o0f0u40UhBmTManprlD/B+L7ji7tctWDoH955EkqDSGyeMeR+8jXUEXiQobhOicgzyaCjqxd90
2CECHP0cTKEloUPC1Wm2Ids44uhrypFZbHwCD9FdJfFI4Hazv+aW91fjz6CcttTw0QzxmSTffjor
F++vPkJWTTsFdxa0e02N8ZHoCAs5/nc5nYRicdX3PyxEm35crtDnbGo3aewNIRL8pVADm6E+lTjv
3g4FkoHV7cyTlEBKKzphsJt1X6sAibaJFSjJZZZO7sJZbF5dJLqfOEjPCOopBVChnkGKA4ycWqq0
tDSKkYaq+YA/I+bqJgvZcHfx7c5rhnwe7upxcY+7b/7QqllXFaNI75cYAJ4j7wd85q3PjbBMv48t
I7ydUyfEgbDSWNkm8+MwgvD8PsKOlNQjaNQ57ZZ3/1yPpgu5VKy26Ze8+eicwlJm1qbmmbBXyaXA
914gq8oRByp8G0n/+gZWuFC8mEY6dqqPskFX4XV7+TNP7MJoVJ5YYJvondZAWUSBlD+zcakdYbI/
gO1qi7/2c36481UyLMpSBfTMgXLFHLEZ7XrsUoxI/0RMPylqQ/6NXrdyCKDG34t5E0bkvnRizLJP
z4Vg5marG0PrzobxbJ0OVtrIopJywKFu8tjp2vY9Zd3bS3LDd1dbzYQxwUtRdJoyyizo6ukm7p2R
s+Z187bqhY9ENnoSRmEVPO8GoEMAIowsuRZoQTz3TL2D6o/lApk6JCw32PBfCfe3x+u65AQRY4KG
Ws9r3JhMcurMaWwKDoBOY4ncXWOHFWPeBmsaKSzd2LDBy+i5KmgT4hC7kPL5c9sSkKTm7NHq7LLN
MqifvJEsu7WvWrYDWOqpeF+anWhfmTsWPXb67o2YRVmio98GhwfwrUrYOhzw9ntckuYPPcI//ppQ
C8m27qHD2lntoLA0jA+ivfj+Oku45Ky35SFZ1FuS85arf7HC/UFUn57JFV+coF3R1XDuAekd3KnS
8ws/YnP9oanL7Tjjq6YM48sPfyBHS7WeFE7EUJmBV+Um67hyMrbpiM6vVFCX113ueCqjyR8JSjW4
BDaV1YvE96JedN4LjuW5uWH31aNCbECV0FZKRY770cANBkPM+LF9QQ6JOYsJBcZBYxV5skYyijPa
szMswQqpEoTLVlj1w813LrF9aaFrWR9KjW/tLOH2cfZIAK3urLuajJIlnj2ZJtEJrSinWCvB/uvd
Nk/oDs3JR6ZpglTvaxRl67e8OfX0SiYhKzJJ9Rhr9mLBBhv7tvRtGqwlERnnZn6Wn4+Nx7Ap6Vlt
j+ZqN4lKL1clUH5rY4OiaoldmbU9+RZRwi6h1r1A8m9weimnq3R3zSz68lx5R9fsV9/+JOxnx9Ei
ionZsYNOZnxK3u/b9n556UTdEVBnhWbEqgIt0BQT4gsDuivAzU52iCsj70tinaCoh9QAxr7RSCWf
0LjzwltYaumtPlUQZvdWXYt00rAwoZOEsXqeAco3g0tHL8XsVExED1mOecvX+NcxjMlkM+zisc1I
Xfw7xC+M5gN5AGQiN7oexElxevLBc1V8N1/aaG0M8Nb4x/eV7by0dXe/Ru+Z9a1fGr4mVmIBmNTr
6c1nYCR/U7YC0xKScL/nkpVpVV6fv/kl+63WbN4sU7vOcMLdp3xluKcqPr74VbzKmTPJDirsX6pf
ooktpjGbJretggfQmEL0MPUZvoDHfVHDonsJuJBs/vlen0LqOVRdTPqvT3adYch/35X2lb6cTmNU
AwIAYpKtGQU1DiZZyEFqyDYJnVmPehUTxi34SYKhwLd0frvjgSGazpWWuzUVLx2REB7noC71LZ6/
GVd3QMjxupfHi7VB/nzbWuqWa/aE6Z8LZlY0llpx5GstRNhYcjcyUFgs6J05UgMTHT5TCIxUs0wG
LL16c+i7nQUHqj8fJ6WMZCUSsA1ujxIFgQXr79/7iWoCSEGCh1JPbmu47Lz0I12b53MbBJzJh9kV
v5WEEHd0efYVsfRXJBD2/vu+7qHZvqJmIg9hRrKYcbgDyArYYeGx4mnFfAqTkeTbeWsxG38HJsid
UV4wP8Jh4tRvEK6TYDRvj+6+fQAd6k2U3YZdiheIp4kXDAfasKmE829kyRg/0cfOsvNZX/1SL3bY
5nWysgW9HX055Y0YElJmnDNzoFEy6o4DtUqKfmN+Tb2n6Y18pbrwWEirCYXTI30k2Fjv1jWgfM//
e3lnclyNzB/jObvaidb8UnjcugepXXvMkRIu7XzSk1lVZt7vZhcz+sVrnaWl+9y4aavRV/O1CYuS
Ns0/6mUoGS1vqmxcUP55btHSp6ktIeQWMZnOL1J2jwn15j27ywvkgWAGXeqNiZX14NWcuOgf/VCR
MoP5oLPBh0oPjCnafkBUj0KOkT/CCwoCoQ/7IRxxcmN4Spwpm6IPlHo16OKqo3Gu1H0Wv09/6cC+
7i6ukYY0v2Y2etZsKchvTTuTOYHyOqgaMP7IYKrCscgeWuMTQ5DN8lvbS1/gjRRgNwyipBDN1P+D
qe1NraZURY2iPt8riD5OcpoAHpYlqsymBQAdEpENlTaCScYL7my6eGC/kWcDUZ+R5nvu2gJ4ZIYM
7K5PkjBq3C159OR+9CZC8EqRvmy1pXvVhP5ieR8KxMLadip7EYcmv9gMwAEE8k6kBRBwBSSeK9w/
B9K0ZA/t4eqSxT4XU/aFjUmnR4jDa4pjfS/O72y1I7AakgS94yJVWBmadTFmVAybW75fWin2wL7P
UkdyqvG06HTlQ8ZmuH+CkoTt2hax0JJRt4slaJdlx8eqQBpriBsRswGDoqD2pNQW5OvpuJ/vx0iv
qUaxKfrmxATxYT169nG6gdz5VFzSyrZYg+tXVkmuGTshh4/Q2dDOx+WYFJeV6B4FezyVy8Y4qi0U
XnJdKDLupyjpwK6q5jhy82ZpDz5bILfr6M7TibPPA0IU3Z0DwPD3dFDRMULo8PyUUFWR+YqEbOoj
vauBuNA1P60upfdcJ0CdmelyKahMr/U9gIlFmiNIsRrqZ0shcaHKGRroKBQX61Lja+Bi7/zhg/kJ
PrR5BRZZ/uef0m7tmWwvzr5ECkw/MzlaRX4bdMaZ2M+T5m0JvFSsufHockAbPSmvgZbUxDoPFKDX
AvU85NT4tj1Dp/gffVEmsYEXzqdvVn/hXTnrz6IbGxCfmRmnas8gxTqIb1tYkhoaWFcdkoVM8MFB
eO4JdYl1TkwxldAU1XE6tnaWoD9lTQFZAbCbhOp+QquV2Y8iQ5mTOQDX1pxj5qhKY6g6iFMrUFOu
l/yrvGXEIeU49kaBaB499859VD5tfJJdnovq+htsRAE4YRfXOoEJ1zyt75mBCHbuEkE0SLKIvGgt
jcZpUTpfAz/8czv7Sy3lowrf4uwnm24zABrkkMa9tgCbEBELTqUJzyW5HqTOqFGR6aytfN8Elhkv
SCI+m2JnfpSh1G6YjzAOyQGxJKQ/4O2Z+YlUyLnRZOccpDB/qni0IseDXzEzhiVs+Hm86fmHuUnX
asRKbQTPft3YjOXeVSnbIHS8ZZBMOF06M05LbP7ClUoZXsI5TWi/BSTWbtVPbiDJvWnIDxoSxMp+
XJoEN+OmYAfeyPkWE71zDy5m6h3HOZvdcgbk7O2EYqcZdzxyYsyVhRGETncsd4PuSJiBFCOvvtTW
7o/GcShfhHPjvH3PAUEIojXXHWiba92R4sH8AR9PSygI3vpqCri/qYm7DjoUo1Gw6XOviHBWN9ii
QciGPs4xNcbgALAg2zF7xajzCD8ZdzSZL+dl1iVYXWoiAY7Q7olHCMhiJdnP5I5VTEszok533LOg
Mq00ob6ZqgMRgmz9Ta0RlDl8jmOpJujwOJyC9RDBJcCe3PCgbwxQeztti8F2LFyyhn2CDpfH2D/u
D45eBgr53ct+jCxAKCUnQu75k2/LjhK/kG+qEi6juN+dY6D/cqA3A92cTKAJSndyRUNuuaicFDX8
nwY9Ib1yH824PW576Ro0ofxlb2jTPuaykn0bulflVtHpJ818bYfaItI2YM36cVePMbkD0QPP2xnk
51PWx8TTKlo6wGStIjmli1LA3Ud43bjI+cUw4L57gDgfZn6uD6DtD6jS34aUeHif/3ETCaZmlx75
y+nlrTa2eVDSJURHFO6pfl2M4ZYPRHhsgQVm/bpN9BPby1+FlVexN81NSc5FOzHZ6hDghkj+z5UH
xzFzOksHS08c08N6PF1xqYYGc6UphUcJA+4WLAHvwlK4femQGXGfsRkb0/caiJ2VmM3ppvV4f7iZ
Zc6mIoUfAH5Zel5tCnDHnRe1VxTKWQ2zR0TOYPk6qXEVJB7tYP2EbmCpufDML9BmYRR6Bf0Ma23Z
nMFBnHjBJ182NbvOQHWGL+Fw+DKK5fyOfh1hXPxWfZ70oPOPTxeHfT7dPDF8cQ8UHgimtD0f8laP
aOdNFZ88enZtfVNQjtiif6wbhAGrcvHlg7nGx8Rq+ncFy8H1TWlgMlSV54FySz19mHvbE83shHgw
k7cEA5Kcv6QKZnH771WTQWQfTibOnJz6ccA3unEbH9USsbxmsMNMdPBQUhunxZtzIMosE6gXJTKY
aYKSMvR2Fnd0TINXsZp9284jzf1/pgB+ryGnLVlMj0R14Y5D4hm3MyFdl3CTq2XlnLdC7ZYZSxxZ
XDuGCRolH6vHU7gINObvqYDzPGaqqQLqUchPHQt+tnPKKNYX0/2ZegcYlifQcODQ0EAkAs1tV6/B
jkcZygy1xfw9x6h8nljXqBc2+eCAlJ/Okxv113WUhf0l9WA2jyTERjUmHqtaGbhNM9b5saaQ8Mhg
7Ysca2FDHb9LuUUFyvzyWolhjqpLax+VD64OzMWA4Vu4NVO7G2oQaADSFSMFYblPeaDYEP9rCIoa
MypwS3OwJjr4yxyFE4eBRJQrZYYX1JJEMTdNM6sHzTAr4tRszIVe5fs4cTCYZVYwGPmWsecie1TF
uE8L0kPuGg7o9b2XWuoja4r0WpQ38b8Ws6FkwOzu4Ske2il2aV68CmuXIgrww7SsmBFSM0ltivEK
KUfRMvgsFOaSpiQsA5sy4V02KgX4cJLFvPMAqS6yGqJtuxH41dnmmgAyYeTh3a/r5NL7lZ+W9i/G
EHdk2IVgRV1dYD/PzndB1tr1E3eHK4Odd0HPQuiIPtKkWE+TgM57M/AoSuwD8iypN5REx5/kIosM
Eyne7xuxIYIXq6w30WYg4z/o0i2Xy6M0Ah263sIKuUUBGZhtqs2ZWgK5YqwGiy1Zsvxlv9VVcERl
/D+ABiVYI+ijexUb56l3rXEttfrb4UVn0Nex+IBQNKQuXp1MmJcxbT/pQqjW2SC2ttx5K18aVCSZ
KoZBEHkbACmkqD3KRy8ZfO4zdhnyFFUVEURo2tctr3yY5ujiVnbtI7zcI8ul+P0ee14fpawl7tNl
zhET6Kers3tL96SOVpihU+Av/e4MSYMbnASilEAk8tms2kT4iE0y4eg4yMHHztTFQ4sZ3o0kLqBF
XL6uofcyVB1cIljwf2Ae9c6Tq1lIYD/QKzThiTK8cVE7xnI8/wX8X2vwinq1KYcqvW02nY5LkLKT
Jz95ctbcdigXJ9mibF+gpJdbuvhpiEDjcF3AzlegBkIPHZyIpZQMvWTuTYSmzPA4peW7BB2qeUpZ
Xvne81KTndXYxJlYGjsoOYJzbjt5Rqu2EWqIMOkZ+z5q1OZQNlxM851WmxOepLFrWolPFmLRYvPH
oICsQ0y9DsR7kceTl1gxGA0+y3GfKYcsCxJBeaO8ROxZxDEoH8O25oSkIeBPUAW5ur4xS8BbnkOn
chhSqqchJpC/hcp9FMt6hrJfcc9DHkR0kE5HMJeeXuqffWxmWgm3h54X0orjsdmtYZ4mAgBISKsM
i5cLpCBnkJ/WN+95NymyiYda3p8Eku3jo6+mshfYEDNXo3N4BR3lAJTdZIJKBKT7seR2CqYoLQXJ
7Yk4uZa7PlFd9P/34YZTPGwEz4/NFumGdYAC//h4GsOdL6fsQEHy9GlKfKCcYV/q31vqChoJBiT3
TarXjfxBptUc8zEwHBC++gESTb1SIoa7aYUNVSa6ND7R1lpuSXPE6J0807NVTljioHDq3HK/Y4A2
WX18SvBx8wUdehwYUvzv8G3wApjYilmqfZUq/uNGn0aNy4W76BjTM7nLDFsGZXWN2jqCkHqo7edv
WhrVGqiTgChRJgGKv6H7kAbQPCA3I0BYMxZQ/zdFhD6iLVuIIaDfYvUrGGhHKu6Ci/vXztTvX46r
KY/WY2QJ6C/i7098z3AlC8I6WnXsQiAQZFTpxw+mGPD4PEruBeSjSZ4Jw3Po4/uISWjuRebPeJiX
MAXQ2hrMVCW9Q64lgNfxxaXfx7SxAkjAT8AGEO1Io35HlDJxULPg8Wi9t05Gm/AoJtmruv/YfeZn
ItF9Bs2EA3taxJePuOFxPedNd5rO/r/64dcemaPx6hFDg9hMWoIij3eL4fvvKMw9IMKurU+iBl/T
3RSfWDZobzBFqyDkFPRi6E/wPjG/BZh8cvBf6nYPz66JDpLhzrP2mjLJK5YeAjsPo/g9EuWl4Vt1
DfTYoQjXkk/Oa8Y+LYqEvgv1NgA9XAjDKyPFfqDdInsR2PerHsIalg7rm+mcqPTIcGPYtXyn0Cda
LktR/d6XqBv5mB6dUNDR7u6TycxdJRXQOLQWlZ/XO26LAB8HMBIY4H1bLApDqi5Xjk9YrOfku07T
P+JX7PTyxuYXFuX0ag87F21EYF15nlJ54AKAg8j7TJ6wchyikIhbRTlBoQLe6LQyBYHaI4F0oqpr
ObPqL5YEldy6EFXe24LmEpr1YIKJqXMdAau+eZmDN72zUPMV/SG/Ezeq89bwpmmwY82jx2V62nms
bmd2fD3l5EatZ6jo6UoArY/CQRtCG5l0SzimCFSKLPw3SjzBDoHSFa+v14m2a4wr6KQuO3odolri
QK5gUN37cUMZSGaNKGo3CqFnnQuDkVOxaQbW+DVCxRDG7AwS7Bd2ymvxXNZQnT6nMZv11cZ/U+Wv
TDmE6zYK4sR1EREnBYei6vRWBg6Fc0Eu5dgO9mdQVlQwcLVvfBIvfcJ3Pf/QZN26pfBDMggnu8LF
m5dZOvXt3BBPqiv1AkP3UPx1RLcK/rBRWw2b1NPS6d7zYIPPvFVcJqHxPu9P5PKbn5A+iMFxzhJ+
3IOjkC0+2VtNXHa2SQ2ZJfe42zmH9m9pQd/Ye2WHsE5ImsojuwI1tOoQydHia4ce0n/6SgeaM3G5
cjYPryycurLjewkCrL2wCS1nu9f9WyuKeOMsZeyQlT72R3OMN0YUAUAcl8YYlRqdgHFsE+o0Vn7q
O+S1vJCNsdVFmKHdQzOMD3Ethqd3ddHnUe3jXADm0ZBVbQxHQrnoolC26unxfvGtqdH0AsLiWHls
Yc4UNp7nrh5odTFKOHOTlrRVTVWstRbDFmKPJbi+vJdm+75VMxurBBswTLkhxbqMB5rfs5XZKF4U
vYG3bwMX8yH3lvfiFrFslBPcSgRqgqd4HMvKoSyKWNy7fTNUUoYyPvAoifapbN351095pkqHPf59
m16nfgeihjz6rWr1Slpkx2ffk/p4CwQTCyAat92RaWHhPoNv50YXm38v+vrQZYctYe2tLInU6kmu
HlanjwiPtbb+h5EOASilGQlz2tpjAqBYEQ/1pAh7sv+JMiqSqSXV3+WbIpG37pHQDyC5T2p9+zuu
m+gQQcZqRXv4CV8KMaufmtrxUYuqtCgZQyLiqreOPELJEnxEPWCY44KP9NmXYxMvrhJzT02Uq7NH
Z9St+VBgDKe6vpMivjJRmLpSu86BLwyZbDKPwZSaZZaGnDPO9iDG+ynUc3D856SztHWM3d5EbMZv
Y2G1Jh2lVtBbg81ulwhItng0C6b3KCy9HWc3jLKQK8Y71KmkEaO/VvtKPYI2QyMeQ7SA88kMy3HX
m+Z+1+O+HEboGQdsvZtN1zK3hgdM4t01OAh3Iln5AwWnNXKN+Y2vQuJuqU6LHn78HTOLM3PNTKs7
8qiz7OjqRTItq00vyDTezMadS/epCSqJJ4HP7+weCpImt7mjSp6m0lOs4PLvp7WtJHVoSO4WBeyj
DzthkwwG/sY0JyI2A7FAIaI6FVqnpBuIfCtscJr2olCX1vfRQhwINLy3uH7is8V74YFDVV3cW3I/
OwsA+1C/4PnQLpjRS4JaSjwtQ8/0FauWhTSAQDraHcURq7ry814Oia1aVrSasf2tvvQvX5Ih5Ill
dnDH5szqkbbaKGfSqa7HgZcXDd7ztCXQ/Nc2qEvmbmbIXxwBzOP/lx2ywMSlW/Vc/Ak7FOylGbpO
KXLUV8+aUiMFq6NnjmoCe3hykFD298YPMRpRFEiAgKfmR33sR8b7bUOh8xGFnLestGljJYMPNORN
FWV+Gde5ADx7zzmS69lZOZO2dl7VqSrrq+CZy5ukD4GBMDIE9f94BkrIzgCPhCwL6NacnrtAJiQR
uKLaalZGN63+KWRb9AJ8vmNKpT9x7BETRgRZqM2sA3FyECN11BhX9fo801HOqCYHw8paa8WOXZGZ
hsT2Va/i1xsoS7hGlo9fOBYuOEPJbnuDMJpxiKM0A9TfWljZHe5mP3XW1KE1+n76fLn37bBG1cpI
eKa+4Yy1JKbmT81LmHpCqhTB8zoCF1UjgMkAjTOwdTnfBPurxR7QUSXPz18q5AKmHPIsMYu/hb43
mRSdPDlXQXGG1ZT8Uh/O6VtAYvAvAbG/xmSSczRhUL6oA75HUkomR6VyFMDyd/1nmr8CcJL+8Aon
YAjnACKwqFAeDhY1+jptkAiKyEdwnqDb8tMIVJYQ4yTfdEI+faX3L3woloztR63Fjm2TciYIDNo2
N1Tk+PWng0n55OyZxNd1d/Y8kKO4R1+pGKX1A15cz8v8C0Jndo2mazU8YR0IX6PUWjNWJS+Ccw4W
J1xOeTfJ8auhqPpEMyyoFDx9jznfruA50cNlTZ6uMwrbeVheUSIZ5LJOO148dFckR1+psURwfrbZ
AUXapeC8R0LMpPLDKapOFIPeceAtSI3u/hLH2GsXLcW0GgRd83C1pO5c5fxdEVVKCjxDpyB3Nc0z
LjQxQvegPY5m6iFNW3uyRYOg/3N1t0obmOkLG5qcGAyQ9CQOrPMGTRCn0CcO5xFqWUBHQb6lKSMx
5xlYWD+MwOabh3Rnbwc/dBeyH1VhF3pa3yGp7K9BnJ7pOlElfhR3VDfpLfI3Z8UgLL7a2/LVTF+d
+W8dVYlt5mx91Ksst8/QgKF5RjygOvNZQxchSX2IIqNrNmzKc9GOZoniVaYc+l0JfkaVys9W8DUh
MYy+A3EBIGZzH192aaFH8B5vzbxuV+njKqlxaa/JVnpGlmRIcQsnYBDwp4aEzrVtYEwVk3u45Hwj
WIH9WxWLJnewupWfVvZnu2Vy8s5JAAxX0D0RumArn38+Qg4j5wbILWl4cJpV53dgKIZFChKWZSVP
OttASbtG5AMOYLNlMoEKZ2VeTviooOur7ZzvxH9jYfNyqb3S4y0XLekr97CRjA5LJE/ASRZ/WTKS
pwf9AO9Is2AfJvxGV61Ct7IjfhZVJfi+MVv7Bn2SOvdLCUK/Ge3NMgrcejOCfbTe20rNWXg4WYXP
9/lTBjihdLFtr1G93oiERAunl9/MuAMLFTyAMjqHuUFTCempRNO3UWVvDoLkxKKHNDRXOREpdm7k
WK5B6rty5vI5N1U19adUztFXA6NFXH9EK9hxo1pa4R5V7eW415MBzvgmWBQ3TzOolzn2POa8+hNM
z14bs9DEombhFPlYgTilanp+HfXvjiWoj7Ku6FssGQ1TTiuHDUfSpUjiGIfJeeH/A7P5nW4hUHAo
3AYmQ1mWB3O134Q2CiYIxA2pxfIo7EfEdtlY4hpxkg4SuMX1o+e9r1P3XG9gMZZpr03A4VhrVwsd
VlTuMkOIjty5sNyn1cdXvOanP5U6fsYxVgvTNdxawriIUUD5kFTto2okHb9LDpgd9j4TWtCjhMlp
Z1Vua7ynw0jsmZcrrN8wTUlo49N/VkiZZm3Q1bMDzU8YhgfAuQJkbQBpxrDYsBlNuBHNUIZYBKSF
mhHKmQyh65/YYqo8CF14hbwDWlkLhEJC0gyTyOs/7R1jB9Dxqug++AE8kd3ITN/5ZMW20Qe7zd5O
AAXIJac8ADVd8CkCXOyeTDiXCQpcT1Amcb1Ka+3Z9z1UW+gTJwp+4N2Bu5GSQ1Eq3oNv2NfW2VY0
9/ZN0bOtpzni0rkm/sDRww66R7PVb/cJplLSEMx6H7c2UWKlPZat4bebDbPaPRpLUl4fiYaJ6iPR
wn/UF41fI8x3gPKjybjwTs/hGOtXG+V66ea+yhOtja95lY21lVOn1M51kBGpoC4ZQlwYlvcGQAZp
l7aU0l4+wcYoJYpw0o45Cni4WD1yIRVq2SSROk6Ah/wb79XHdgSg6p/hFtt83a8kzSKfOgO++wWp
MMIjO1Z7mbc/aMaI7pa/LqD5gXdTSutW7wTOhBB8c2jb/mgYmNtqhKZLN0TgdP/7jO8O3tNI7wNh
+v6MloPMSY+2zBJ9vZWPXOt5hwAbSZA1VMXX869vl5VG6USXb9lES0PwG6Wexi7tRJ9XeWJK3kNn
hvY6XbXp21bQSFzwx3W5aa2NJIwdJWpe9VZdcYnIisKguV4wEKVq9h1bzdP018AWapaZeH6inq+d
2mdsHErdjLR2mkLyOtdjTkX3vELu9CPzMGGAghz9CvAuRpL9rx80fyEhLJcWb7SYmaM/OiBUXSq1
KmqWBzonMyDSdoX1VYYZzAxF8FQjMeTc6LmV6cvH9UYT9ZX32bC98AIgR52VKmHn7Th2QiU+73wR
FhZnyn8Hm17Roodp8jdbJPkbRq9fSkC/U2nkR6jxBwEoa30DTiklT4zDwDx1G9c/LvnyRInQBDp5
qUl5RFFRUroTbaB4W6EjROproVQBYan9sWRkB/acslwgamxGwf2+64m4fOGYTR2SYzVC21E/YubZ
kveQ7QiNPqe+QnR+nIU6mbPykUkYdi0Sr2QHgx+G9CXDWpUr7f6zagpvfhv2peukdVNHbJsYF52m
mMYTsj1nIQe7zgvBerUptzKsuCxDctnMXQSrokf3aPseP0co0QoleLOuSTwH6E92lPP06lMy+Crl
eyGD772D5b9nzhxUgsKEDM4JVSrS0KCKV9HC4Ylb7yZa1immMgHBL5zQf1gtkZyAy/9S7VyEC6oH
Jv80CzUfUgxbXGAADB1hFE/Wlz8u/a2ztiruZTeelYY5aT9ubWyG5VVZZc7uirtiUH621NKF0lSu
9H3AjWY2ZZXf6wxVnMjKb7+1ySZvn/Ibc3MdOpzhctkfEdvjauW5y40bKk0CfVjqW6usIgklWTt3
GonYwqS00q2xSICbJw+z9n/ua5YGTWQg/nIB/9R4RytnXoiQrcGr3PePkWtVHsjV0Wm5s/mW9Sdp
JW7OHhZPewh6qEkUkO3BBKV8sOmwtk0D1zK2MZba/S4RzXVQZjg6aIsszuDYuwKqvNIGKgKPMfWY
1tcpQxQ35Rpl3FjVvDhae7egAA60/YIp5J7ihgRiXo+ItVbHBuvFGQbjGAAuHTBibMX8VoZQXE8C
4J2T9kmmAXE6OHKfDY/AweV4TSyvnjGnA6PHkIf4hUg5AAdnePhvck6BE0X4al5a49jNe0WOxN2I
aAKGrdqBisRuxq3l/rjH7wggroNSwK0hG9H4BGiXmE/lNGCEcj9iJBElOjIIkqWxD5y4CgZzr4I0
NAEEFnY9SfGhMush5qIY9Z/Lg7QPX4qIAtX6v0V5ZUEuUwZlHvUdT1pxWz6F3es6s4EszYELIcWJ
IDyBljDL5x7vT18OeJjhZA4CxS2c5kU3xyHhwNW8LPzgBO7/CgiwLIWvswh197AnykqFNK9Nug4h
13s7HA4jhGzjBr27YDCTWUiZKyjskmyXKt70C3EuOAXmW8zY3mXyWHYO+Zpfzfj/EfjXxoaMg2qd
0L3KSs1pszD3e2CSM9KG7kziDiafSXIskt88oBRXYRdIPDdySveKmRSYuuOZVd0oh54LKLptf/72
28SPabyfzabKsb/WNoQ0bPICORrr5B17lGtbyBfmQuktV1ULR9oKHoZb2wADaQmfbzaugeb6gZLO
LwPT+PwQXfTycVRLQu/ZOn++PC8g4GwTkDCHwbMN/r0EVIKZ+LptPfn/CsmS+n+eh53Bsplx5ZQb
RXJ4eGPOeBN3vEJyYHNe4/g0aQmu7VGtQnF0LJxNXtvb+hG2D9JoA6hX0/rYpjAROtmHYVjpA00d
3WCFjrF4Js13ck/F43gNydDvdiXgjmZIrwFWt54qN1lArMQsoj9wQCMGsdBvx9jMVfhZ+rc/et5+
c1fMut1JdvHH6pyJAWscEjtK0awcpFooQz+HV/sr9A1v9lzPP1XI40fLm3cLCt3GOKGeeM3B37WG
ACEuL7AdDY+i89CwAulPkYJql9RMvu3f2Ap0w46XW6APLwwuMapSc0qMFxsDMTIwInwd9yWZuaV1
To2IvEa9sMsvzBcR+5DqGL8nJ01OCtJok0fxfOMmklDzjyG/k44K9eIKfNbdHHrIaRiUEQXiH5Vz
1u3cExkgZjlQGbvVN1HGQwm9xZsPqvPQ/TFcLGbQr0bmPEJSpgTL4sE7unyDKrrD0P0L28gGMrRe
aTQ49W511R7tDU71uyvU/bZcRWbYmPJ8DFx7j/znqEhndjeLK6KOBK7JSDLh5TQIUNz4skEuYBAd
0uMysKODG2dVY9CtP+7DQDJMS4YF1mgmPSJMVD3iw6nwA40v7pOsag4BmitMB3kBMwj2rVzJCZqE
Z3Q022aXzqAUkLIUlN3QxJN/TekYv08/Ud6Tlwg277JEaO3fi8FO8JQvJz1vNy/yGTDhBoh0Thw0
6HGngdMIVdEBh6NQUWZRFDFikVZO3wBDJv6GIMBP6vd0WDwKP5XPC8MvJnzioAqMw+IEtkPt6Lun
0Y8iICxF53VbUErV3sOh85nRk5z7ilja9gPzMKa4931CJ2dml30zc6clN+xubcS2eqSBa+GuWcWX
+fghn1vuS7IgiasJyfr2SAjVESwWcxZHu49gmOdwxOc6bmG2+PJ/KMWGPxua8VunE25bCgreX/FL
Ftfi6BJ8cFgCRBQHg5S+Vq2TQuUK5R5/yuvEp2YnKasj8vHrsl6KTHzkc6cLnImOoUGHnmQwdbj4
YgfI97DwWxES871Hs8kyMwKsncMPOASu8+GnfG+GQSnPQe90uFOLF2rfcN6ClmEB1+lJzM199Ljc
8wMr5racuBi7KZ8Jpf1sn8FMSFUJwIfYACukTMAa6NtAbXxrEai4BbDrNX9mh7UZfnehQRB8t6cF
qK1EzE28X5nK75oJv9qTowTd8A3cZt+HZSuKml+a4O1HGcNI3KnogH5BDRvinXS+GlIyTou6uMTU
xLULneQVpIWv51tFjvF88V4w8hSGiE4iqFcKR7r48WQZqJsE30JNdBVfamxDeULgfJ52JcolsmFT
ySW9CaxT4nefiC+Luz3FURT/ODL7K4/iWVjRzAbn7HwiFMQVDZoRzJHlS82XW+eR7XlpKu2HIqJA
T4GsS2wB2S1YLW2b5IHrqnt7WcfYoBD8SdjGaHhvFJWh1JFJaynT0hf9zNS+VT7kO2LmqPX2jRfW
NdLlNxK2BuitehOP2Z0abxG/VPO2cQZWKtkIYTHb/QuX3iY/ZdK+xPGfNJBtvAbyy49Ll7B/Flxk
JW6S16FNy5oH4GyVu1GglByuBgOUjn26FWVY40koQVAlQnDCr3UjH4lzyDRSlXe71RxmQptGJZI7
OPWk8vfPpv67f6OuhaSn/1bPjFYZZhjjoxn9BFQ7IE+MF3/VMC8Izaw2sYDMQTepHLAt0vjb7pm4
K34Ohs55SKme5bEktYCSJhq8+DgWK/Cn152W621t6WTXVu1ULKzOY06eNXFElakvU/G2x0ARjZJr
+QYwzWA0O1oezuNeuI2tVPVfBpYZc9p7wqxH7toDQWHemali8OocQJKKG+MLw+U2Kxi05hgAK52c
fr/Wp8qfO9UFgMTFuHYHUk6C1tOlC6YNC08HbzfTuWozgTA9Q7whDF6HutjYHbgKKqB2H2XeDH1K
9bYDriskPqMkK4JPEonHlvKma0uHTyMhPHrkHvESxMQLcsXrvTCD1F99gtk2/xD3kiZIIIu8h7iP
+5OtqzsZ3jhPlEjsgLQX3iJJT3l9vlC2h9tWP+tDs7F8sCbBHq80ydDoeOYQ1pqPjNftqUMWlPj+
BHKvifkkZoi+i/jGLVslH8V53+l0IndhLFgj2b8D9C6srkxshUMpf9YYWYoG/FXXng9CKkpl/mIS
eQ2lTYHMk8MmRENfk0eJ4I4dU2brerwcdcVhpgaFEwQfJiHJdkg7+Ra25Cvoz0TRXJSYc/DwTOMg
/mw6cpa3yBkt2cPastojtWBCHLLhpA/O6Bg0daKSGQBwJZU04dD5EmXbLPxpkvM8267Vdr+R8P5x
JUTKMsx0QXDGBj10PHsl0XQuapli1lqFRFI6cQMa6MSAJxNelbOa+RQQDfCoWVjxB9KutLwG1TPD
zne23jKEaeCWFPvFIdryH8OfrdbitYjfs0Kr0+AM5IjOM4YjzFWWJMayHDgOYDVkdTu2AjSUI/xj
C80TG+h7xIc5BPmkwWWGAjJitjZIzuFjh07Cjg+cQtzC1pp3L5E8pzvLP4FB82/fxhY6/2lq2QGj
3IIrmoCFxydji3UZJ+gLM5qgEKigctgGK61qaa6lmoYeNVhcR8F2WzCLGXG1CBL3zVoDtKO1tJUV
7yl1Ny276raHPxYs4lAAV0Iw4SsJq3EisR+v0AJklNEy1rWfhbe6CalGWoIKhrkRRsw8QBZY7d7g
ep/S0TWKC17uP1Hmk/3u3SgwjGPXCq7MQbCK9yEmxx8Vqp9Ft2lvZcfoessT+DXUNNsWnYCLA2aL
qAqIHyQJX4fywsCMZvfDZ2avfv104k0gnqZGYmMIVeyrNx24IPC9/VbABnAK/3cvnlz93PRsXzRE
LOTAE99I11PNssyUbaa9pHYzq8WauvYbqkeeVw1f40HK4OEyKzl3X4ZoL7WuqWF5PLG1cpdb7dWm
5afF2jAHl/W2uVBilhfsTEv0IZH+cnqW3iSuxXkQf4E0yucziEJVowYQcYHi5SOv1b1Rt5mdmaI0
2uc5jV+ut6JqG/6cGS+VzZ/6/R7Xfa+Jvx8D/fDBKSkfwSpvs/fNCB4hjwWXPb3pJG423K+waxhb
TrDbl44iReYmueyXbYRNq07R5VIorrcSwS0l0A3QoGIOIjQwxbwzDpbFoSWbGKPeVTfIO38sCCej
eJ0m/mnNvdTdTjmI3Ltt2s6elhzx100/E70DjSACqcErQ6UtZmHIPgnYkI+xY2TJp0VTWtnVT61W
eLQFO5BOr65WyMkMbJfhPHQzZDVGZbmYspaDUeS0BdTFE1YNrcoaEKVTY7BJ7CEe8LBvTwCS2Q18
M7HFKCRLBHrxMATZrrc/xjLysLH/QpMjfRYlFsAsoF5nvWCsAFZHXQ0+WaI8yCdTtBjnaoCs46oF
1Wdg5UDibTnOqumkfeBHjaLY21gfaNqmcz7oybpQC32v8JwvCziqKi9LDUycLpUxm+Vrh/DLZ2HC
GgTWLNnk0BgaZPwOEdxPcR/NP1a4YEAVlABLV+WHMuzxs8P6qoSYaI8aYJVYnXdluXXbK2m4D72c
yX055+S7OcdK+Cfi7bF2kcjTpNbKduH8KZ8k7lS/IWxSEHDVoaiUpHscmCL0mwsOjNtn66fNw89w
u+A1asWJgfrB7W5vO3wyThkTyuei1s9UZ9peWCocCa7OoAbPx9TxJLJ116uUpMZiNv0z+EHksKUW
NPvBZfT4pxfxrI86kEzPf9fEXZYxLSmQ+tFN8NhlW8f81snYjiuYUV6aALLxf4bbpJEl94zzYPIN
b46QmRd8OaJPUGdQRA03mVEJOiPOuYomxfOmu4EnrBdfuOYGu2wFaemDmDuJYgjxBuWMO+Lf0+nr
V+ohuMwi09X99KVAclvanWBqUNeUVNpaQmVSXxEeoSBmBGsNTl9iE6lAZ1TLLxNV8/iZHv76Ea3F
3I3IylenIuN7IkJ1m2KZjDkuAg3s3hDRHdMNdtE/lC75iWza8zVEqGP6hxoyU3/72Er5oewVEHcx
M1z8ojpve2xEZ1W8z1HdNIiicDidcPGAA6BlXnlUqVHR2vpxs7D2yyWY+esziGFBqHlK2hPftQY+
ZgGFydIwVRMJOO3Aa7xIhym2WkfyajE8xi8mRy+BvnF1f1l2BXcNj1Aao5kK9exF/q3uc6D1k8wJ
+CDwDVGbClD696r6Iig28QvPQSI6KMrtuvrPCFxMzXNmLO2YEb4x6rYibHUVRHdbAH4nm4sBoHsa
39hCBAaw7o6K6q1diiDWHMjOcJwfoufp3JhHYTnCWDUbSiL0F6uIoS8c+KpK7ukDx/A5ui8Yw9kt
ij7lgXxSejotb5gqbdUL9A0hrL18hqWk6V1nmuNVCkTGLW3StBNia1krVx3AeIl5UhsTo+89ud+S
0v3kRRxVouDVCou4bJ6u7mRCUXKKUeKwlV7K/PluQZFCeaTLBXLzXgUIDR7rMWjT1NQ77X+P+Y27
1sLbNGUjn24UIje4tTxlVBxosuYXF+jynI1XlQpGokSqiCLtQJFP93JE4zjGbsiV8XlxjEmG602B
TAEB9KeqFNwaM4/fYL22l4EeP/n8nvdnY2DR1lqae/vzKNPumFXojNRiI56ZXOz7wK8qix86mA5b
jhep/KZQp5loHwW/iIR+Ru2ogNR5++Pzjua7HWE6tLLd9TPhgX8OT6pWDdXCn4cpUEe7Z8e7iQX2
EN6r+4TBa0jvCYpWxVYoeyNq0dDShxkqSVkPsYooIM0trO+IexoBNGNAiLRFiwpdkB98jPzW2fe9
WLVTSSewlxsOJ7hMe/MlIPsfEDRYha1zAJ9vs1Xy+5ebcs9pLScWesd07DXoFTWEJnmDhNYqR2EZ
usBmw3/tjlURJrifLarUzzifBJLsAHY6phhW7Es5+SneCAw5MKxn2ettlMlhjmzwo/LJwjWgorqF
nMH4G9fl6jYXaA4l0/lUocqtn6Is52GP8eQ0O/ZHeB6g+/jDnP9xvjh13rIQ7NGpCy7+MpVFCyyb
hBtABvKH89nbYELwrhvqCcjuKfYDHiw8XStNZbkRfewLOfQDE2j3fip1E/dLBDzAT05oZSuF/RJh
vqBPNQKuCgDH7C2yNzCuuZ1SXJLP47SrNa8vypfmJPKrF1IveKzD6lRH/bf0UNbAIhGGCyRtuNgP
qkdlItFNPr1mgW0dIlkeeAXYlJP+Ocw0ZCFWTQ5LPYX7LxyPbx+cc6Of62hKxnbo1CycdWInO+20
++zqLbyiN+IudWz9ymzSCB4tl1cozZ5oFX593BFIy6955wXv29+ogi8BZrvAvgkem+i0Jz/o2MIs
rek4ixdg0ptt0MQOItyrv72hdJX+ZmqXyv+Pat4kaqd7LBOIqO5R0fZaduDiQhm/GiaOHBIO7LTy
FZ/+3PeprqiyFUMiRANoUUXiDbSIVgeR/6L7MeGv0P2vsG6L43tkMcMQJrdloAIZ1+G/RmcM7wM5
cuLBOFlXNfZ5g2cRCK1Hl/XQRBtJk09nT2n/MU+krPohJ3xuZ8jGGPUQYDSYJ4e9/CpeowL2xNmX
9rxlB4laEK0wnbX2DQMELPF8PRZPhXDyVD5oTb33GAtr+iieNB9z+vL3bElI4Ei0y1emaE5/qBxX
3PywXiXX8tLHJTJSFtleCXt5IIEYoUTpCoIgSx+y9b+LSVZEpIwh4IJmRXKenCJZv8qY8L+ru8qm
+JphaAYxSllz39ZcQOZP8XqkAqw/wVjTHzKfg5VthsaAZupBRN4uW6Dv1hNYiqZC97i5bUucO/hS
JhglqdlUd59/THhMuvRC7XBrh+Fmoxix3Ra6JopbLUYm2Nw3/FXcjoyZ01ERZFyUAL2muUg758nY
BJf6K6IwPufcwmVimn/ilphJ5wwudYEXUztZ8MtS8NHPH9aFCWofGUXW626GkMoLNTKjFjEsfMNk
GCCtwXi8SNaRNPgUOUGdkeJyb3FYEos6Ww2GeVYRruwJ/1juG0OjRQTTGWiQKBx0YtiTIxNHNWni
hQm5qcYvDlGrA4Rq8oHILga9K26bXnJKRFXVUndQ4iLZ9IfCaE+xL0fzgdGTpHSIbXpHgZ3BQjwc
+hBPmv7tYMJ/5W/ZuS9+bRLLs+UtHixLRA7nMmj8zidqGX6BW1W1wZDJk1u0YKCItjoJb2bKw4zL
sjG2gXtm57y8c2UZ41OYkoGnzUj1sObS7fS4Hp5ZCjOzh1S+wunXm+7x+8hG8Asd2ABVq70kR2g1
Sj+XZ306Oru7k23vHe4YKojbUCM00LHWmx8RfW21etmOkjDLgcdNRnzH486UFNncHbi+ty7lH2wm
3EDGMlFZHJCMQjkGSbu5+5ysS/tefNtZUO7NwjPMMFxpqyp9TjpwoVjkd8vdvDZacLRZ/32l2zoQ
/NqRqUjSdkkDRfD+Fuo6AEE+aNxCFvQb51yk5JyD5/BAmX4Ui9VZDQEhKwnhVGqXEHozbnM24fQV
uyfcVJ2Y5KVAxRTDP/z2Z/BYXUTfGvvN90/7cJsRyu5ahZ63T2kue4eve+OC9nUGxekkQfLOjnx2
hyWVOUfv6WAORGuIvYsIjsI6h9KIsGbqEKuVqRaSleoUpFFQAR+tjXGR9eFyQNw66EeDl9NI3q5W
eb90Q4Q1u9fWm0O3rvp8YrYP3OvfBNluiypVzQmvaKlGIj3Ufo/okPEuy6woQsyNq0mC5mVHj0nD
uslzg0wna/vvitMpSwdnHvuUSv11w5RMXpkmHEE7IT9X9p6fK5WbxpHdpwixAsTwwUWiq9e6TDok
aPtiBzu42BGx+5JbFZH/ctO6/VXCsCDVmPqlyCSyVGguugLI1nF9q1udLkKcbo5vgS8RWdJBOkOz
E2zQuI5UXZXNkB8YOpL2mdK/Kowb+hz44yq5gMM5+A5AcljOCHdTHvEuUjA+/E02fJRNrfrFHnhv
IKry5+8PBbRepLwKo3ExLBt6mlvyf7RFGkgaw3MzFnTHT6fHgdbt2RA1KQyuwqLJeneq2DHWhktK
6GqsoiVg8tBEjklLLURxAwfL/nI9E/NwcgBvFUvmozdEwQ5h9Kr8GV0Yyr74JF2JXsgH6btufr+Q
VR3shytSUMkyVpmaZmqAK2+7WvT6K4Gf7C3IJJNq0L61hXGwUQq6vLOR+5vX2Ib0K72+ZXPdRaDP
lvYMli6DIwqQ1zlPPijj0cN32l67DCjGrpRExYPOnsh+mo1FZ9GYEQjLzdAsWAJeARi/yw5BncNv
g5rRWNCtwDkvIyLOx15m08j7MacBPKie3IcbpDw8C3IYv74L5ONv54tAxhZLmSX60KR/Z+Xg3ZV6
p98bbxaTkFJ5cGv2o14luTbpm/mj8EwDFlSwEV8aKd6eMrzHFaG452O51VaiV98T5q6whEo2YpPu
UW+D+tJRLnLqGiX4svGKUfJbI0IKIfNMzpI13y53PhwPTZer+HCBmZDXXq2eZ/r6X0O09Ca7pvAO
Vd8V0RMlxe8kdULxJ6uJIgusS83fFk5Yv8EuUUlZl2SvIrcwxtGrqkDG3io6nJkAs9ca2cQJrGKx
x1/jlYp9Ikrnenv1xxXmMrVF0EsEmCULCSnWfv8RVr67KG4aP1JYFD7xYlNgHAjTBzV+K1b3Enz0
Nt42Zbn/2MaxCeThqidmUcbFyA1e64yaBq5oL10Mp7IvzO0w3wueVZ+WWhU/EgcbKnVsLi7eTSG6
Z/+xcBj8E6ShSiEfQh7ur7fnMtxQlLi7n4KzlTSTeDaApnBdmUty/bHd7GMIx2ardQmc4Ttj94bM
76He2NkcculuguaHI80Yeuony4TbLcPTkcYg6cSS8ZP973UdZiGSlv6/oRS8iYSiTjHZhuph1G4M
Dt8e1zm4FE0MmOpvqF1yj8kRywQjYAEziPjH9sk+mm1H1o85Mnt+d3nz9GAVcHCr2CvrMsCUJHTP
GkUH4J0zHI9yHa15Er58k8dzyX1Ctnkg7kEJtnGLEHAc2AP7rQNzIa72AigGuGWVHAD74XvAAWl1
ovzv1hHWqoOojIZVrRRgSu57wgdtb/iOOrIULYIiSNFLbC6RhJp+JGoPMENd//6PdNMYUcShVxs7
9FIj6JE3Z3uLub4cVp0JPojLluvUqg/RhUQk112yAsOLtBbU2J1vwP+J2E7zvTdsAydy7LbtXQI/
Bq0qax6dqT97E508EUyVq3lGVGi1x8KGWD2IjQNMe2Xg4jNvzw0f2eVemJEt4Y7XzG8bi0dpVYkM
qHsDWC3GIXRUDU4wdM5QD9747Xp9v0mnc+0hpuA/a85mdPYVutyw131DQ6mJN+kFO4GUeeVYlArw
HDc0SF48s1BelFdnKh0rU3vHn4eantJEwDzlVBJJPJ1JrumW8R5xUMFcWdgEa9hs2StVuxkmhQxu
d6NISi4iJ09JRB6xeRtEZbgMhAKvbL1FFqgF9dijVtj4ZaVnYpYPocbjxrtsfCniAmdi9uYsISBi
ecZNGZgpaPVmGTep9XDq2KcRvpBIwzdYx2WgqEU8IN1LwedUKmJEDXROOww2Nvi8DzM5qmqS+iHb
JmOfzTUP+NiHoEz2zcQeBZ0X9CtJXEmO8Z/jDuoF0NwjtbGBfGYY4BNPotXtR/JptrOuDrsObVLI
YSNZqd0AI+ROheDJDTl6rQyGK/CzauhbzVbLVzRPLrJ/GD50Z+54BjUH2l88E4lhvEw7ATueeeU8
1uuc4VvRxhsufbJV2ercqL3sobQA2A+1Q5s8G7/GDIuD0sE0GmIATp+lyfnuBFWgl7R8XJdqtD7c
sAyI95egHqQF1XCAEQmZMpAUsHwPBOCDnjFwnsIba71pDzIvTXZ5tX6fOkJumI5k6ncX04AXcYIM
a52gODcZcb2f+ZQe03ANJVBC4aX7eDJTtL1RRSxAdvvTdKY958F5He07ok6a0R18O0DkLsAbRkJE
vpl2907KCOvbWNgtXOv916RiXr7w7khWAQrxiBCk4UYlpB2lkkexubGfk+Otfb1eUVZnlXi+HjA7
/MVbw5+ipcccT2FaBzvc3g/rEeg4qDEWWnGOvTp7Qxlo3soZndz3pThazTjq7WIiSy1uxASWRVWR
6Vdr1cerwAaf+VxBTV/zBj3SHO10qzeYuzCJkZ6QoSOTtANp43bwrgJI9HceYHEO4TiFVHfC5EY2
fUsxXVLkIvaAZ15ttf8dz7XMdrN/TL32L8bMNEM8GnnPSQY11NFnLnpu+NNGkTRgQp/ehJE5LSlq
Ry9H8Skkahsp+f8qdcuwFCY9bMAkKt5N54F4YAtfc62OAAAi5zACG5dpkncHR2Tn5VA83qQtzmj7
HquFwtMV4U5da3XEO27+COLAIqMWn6Axb/Bz39fRnwQzjLhT9THaU4cZ9fVlBsoNk5qEuxq1QSRl
c4PlYUL0EkCvf6AkTJZnD98RoGt95CRC145sc5PE2j1ZRvO3N1kQkw4JXiBtIXOUWAJYKbT7vnOU
EGbwj0tFjjRy4BwqfMGlhB60ajMqyWS7S1z1qZN6v/elIW6jfwEJfXMiuJsErfmIW9HILQWnZrQ3
mVSkv9kvlZBne+ZDCDu3LTgANYw+xBIsyRMvs7VLdKSTWsisqR7mLqV6OJdj1pKSLkUK/7tO121q
xBIva/2hV92OZwa5ko9ZcFfIALyMuwv0UQdUK6RVDEyHSNvA/K+Vo2yeMsrE6h1LDk/8GdY2JcN3
1dQFHiJeiLMbABMluG3ogVRe5v0kTm9QMP+GGF4VLrG3zVwkRhuhhJlyBbWH2SYrQQrF1CsMBbAr
uhcuLbsihgTN++kpZX89QIoCpWTUs4CkYVAIAvzo2R+1d4xcRKLwyiCDKHhsJj34Wf/oe1VHezS+
pVewSLLLLp+FTcwFKDV+tuMn5TgyDPhtPT2cQqDR7Om2nlQHnPXCZzAK+CiFYTjI3u3QquHNxecU
IQ3Seg0fjUQTV8GWRe3jn4FAafTLCDqzuezl7sGC9yYOYTGAnpy9tPqGfGecRR00ngCC8QAKMq/B
zcagnLNKVrB/BYoAZ+0djxyOi5demSt89a3KOPZLjlpf31ZiQBW3QB+EHae4rjf7diVTsxkvdENI
9FO7joR5CGxKTnhbcBV1XsYLYNKoc5DPS0Cjx2UjHE3fv+u866+g3JIQ5MpK5VxxL+6ircvUnqJK
ebd15NcO9yWVJZlHPtLTO2LVUlfZ4VhIru3xSlRxn79woLJNVoAybmnH/IAHz1ODE1f++IvtmiJC
riaaC0SZ/T7vgO7rubVKNoOMvuIcyanbv3e5eeLa3KuUc1HXTIOWMZGlklKMn6dzWQu3dT/qK+wt
isDgvDcqTgUHiW9lWKOar75otW0yTgoK3p9tpm3YOjuG/DcUl5w+SCY4e40DQXdb2u49F4u+7O5L
4yJHcSj5ZMFg4PMRLWQE8P5P7BpPHcexGC4BmZr3eVKA6G//CRn3nPy1wvQ5gyGGX5adQ0bi+dRY
eo/8vGPBEdgPwdjpdC5xuKuPBz5b+Wl0QI3Jf22vpApTGFB57mAi8fSpRkxnFVjmTf2X9+y/ll34
OFHuNQMgqOmv/ph999vmxMQjsVLAHBdmRM2ApYA+2FXLkGFS1phvzkaxkL92RPO/L/YhHf/Z8mUi
sP+k5t/rYVJLCgceiwKVFXexG2AupudmxyvqDWGh6PaPlbS/qjjyHDfQ8VppEhnUoszUHT8Q3iZJ
AjS/v2NEfjhScatxsCKUoCJpUX4fhq/2KMc5zZ9NIsWMJx3snGm7xk0taBGDCzMbyx/tlpWv6IAy
kUDUHLsiIMq8Ay1GPINsXHKc0GKkHBKmMQKQR68sZF28oz7GHkmOWQWqaUKKutVzrQ9gu1Pzkihm
u1G4MZKP4uBHY053RnTteOvC7I3nJ/GvYLfe/CSzBzeITX/ttI0yb/08ik+tBiuVgT6Ezd5DEd2w
x2Y0fW638DE9rbpxQtRq030QS5z2LUuinxVL6uvF8eIqU+XqOBJFi9aspjSsu5mBYHTR+wJYs7kr
Et0UKv32gzmgkCngmgNXt8JDdcYL6LNGaEOXjboIgAs3oPtLhC9Lr+yzc2VNBUIvQTGZ7M/GHjAF
Frngy/9NNf97vARWC724bD43K42ieq0DVjn3Zu9hiLO2WLS53aZcZ88m/uPlJHUA9Q0TqJ//JKFV
Izbbyp7tT4zvEh3A4we4UwC4aZHYVh2fQ1UcqLISi4bCjITYsr6BPGwzcSvciNsfHZhHmWDIbO+z
oJrNU5hMjy5KmeoogfTlWR6HYI9VsSyP4AZSy/aqnx+l484WnEljUx6d2E0yzAo7+44Zymk2lsMk
w5Z7vkQ87QXPi3W7adf+K5kJxz2SS5/mbczSm1HP/6q7GEraz2xJoc+0THc2IlFpzt9PiEfK3Zs3
8SOW+xq6PfUrzuKrRRiWovLW+mkzig2siCmnyy5TTZhUdd97uX0k0aA8pQYZOgoCh0Rf8xU45qmO
Ir2mY6OFbVyQUYlxXJJRgeYVIl6ZnIRW5wDR1feOBG4MRDa9XH0R9Yxpco0sx8RFzf43MJxe4mWE
ZjQtKPMMYCvKvHPrNZr/aJg3YkSLH1W2umDQP/PhJFtJ1mqS2cQmTe6KqegTV3TnAzoQCrVTPanB
hB5cyPCZxI5uQJbXpl9H7Gyn7eEyVfsWD5pVTUYRm6BxNv5vbzlI0w+/cIm3sae5NYhAtPyhuX24
62JAju25EVL079bUjTu1JqKuLP3CKLFXq7/Zl6qoeBqmHnx+nQPrORimM76v/2NyzpGR/FRkrx97
xmoR/+BryLDfchlCZRAOuePl/UJg55neJmly94jts2hnYe5QNEJP+fOgF38qZ9YYFxJt7CuHGCEZ
+Y5Z9zMKPl1Hsul9kosKjkKq2uNSnq1yk1qx3riMn324YJIitmFtGoJfiCFKPsI+NHSHExce12YK
hq62RotOtZ3AMElfg3AM4Nxbn4goS6qpNWCUBwFYzedquKx7YY3MrFd4W0Fwm98apBTkB++5C5wX
AfrYHQ7y3axknXD/14l8yQ1faSafmm/7ET/8rpcJ49OAuBQmJyBd/WElXxhOgEzzqqBqZ399Bul1
DFjmPOCLOmUR4BGBWoCz6OoGIAW08ou1TEdftQP1G2hdCBNFqKoyUjKU3EZSlmI9/vD9Qlusf5zI
IwVa78GxKqqoij488vXe7Fg+fTBE0BoCidntfIhKaGdGrGhZ28+CoW9UrsdU3ZjbF2gwR3QGlraj
t3UlzJypnoPuUKL2+iriZtEbGvRxYN0RyziKhjYhe9VpTP0f3SXHgOlSLLblyFJmrl03mZfTz6uW
zg8NG4zxh3tnj/YUzdI9h52Wwlw8P6vvDo5pgODfeLCUXeMP0uarYONlSGl/AVt0cLc6Mh7yGWVc
GyD4yg9XCvQ9u4T0Ephu8wtNRMudZu7msq9PexI1p1dfQhO8m1SLBIWGVqv+x7Giy/qR1x0EL6fV
82n7D6KCgf02nH2BMIu3HmK4UnjO2wOjmhZ3tZvUfd6tLKSsTWRMRJcGHYKJG5BMFU7rfQtFYaAa
tWNA7AIJvBIzJJw+aGB/Va1s1Z7DvJRdOQb5Rb/oxGsavOHXL60YBx/JLFq0KWq/s+Q7brYBiSs3
kwqFw+YO1cVvKIheSXQK1S9g9pGrKYhsDFZePtKp9008QDE22pZMs8RWS8NhVtUn1LG4CNpGPJzL
hIEMvpgkPqCcIJ1kI6j+DL0qiXs1J7Ynw8G182A7dU0bib0OV/bkmA34Z/va6wtiIBWbezvenWFf
NipLOa79ss/lw4bwq4wjFSRWZtmjiXpSVgAFFQBZ1Fui0vO2F4iw0OhFBPujeMIbM/v/C3Y0Lg2H
sEgJTTH/qYsAliESrWRVP8cbEfYzc9TBfNeSlyA9nZXyF78Vwtails2QrXmnlr2Olaluy10bTP+/
B7UbmlXFZw2uDmMeVUS3LYfxPmHsfaBp4GhgOp+u3NJa30bfywM1kDt2ydqRvTuDVU1H+DEdMjde
B/X6KcDc3awXi9ofZ4lc4sAWv7d0ri1m3Thgmv9J1z9oXmHXyqGrsDysC/9L7IvYQKQT7ZgAt7vV
cC7aiCw+zlipaCNhKEFtidN5dPEttgSukB/RgbUozWaHWsBCmH8A3rWBKivJFmEkh6lh2HP7arhU
l+zwkIIWtwj1BTqxRVL7yDjkgpkWtpaMdk4UNVxGqV8EjhLzPPndZc5b+QN1OMKoGud/H8UFe0No
ti3YwNsCiQHIQi4iDv5GUOB3LEFrJQQYzNUrYeticKSYZvr+sIgishaI2SO3Bu6NRsfIH7r5yZ8F
vzIPbd9cYc8jpx+6Aq5EF4ALSr0JWAKkaSIJVz/SnhSS+CtYaCQTYNXaoO9Rh2PaldRZ0RaqtXZg
oIKToBDzvANpgqjV3mWo8cFwHuCkGgd2JhaW6aRNGNqRqlYcwcBUef0ekRu9EsoWgO3IEJV9stbR
ZvCp4D2YO897uciNClhNIobx5uFFA84E07L7ct+Gyv80C0P8ltW8DEz4/X4AiV5/R6a5fEdWxCtm
o/KiWwZonwv2jVGabtG2MbHUVBi5c4cxmDoBrvMivtb8cbtB2pzXlDPi43b/Z4ga0fUWL7wwYcoV
kwW4w1yol9w+n4ScDohJyNVtMhuSZ4BN9YiVe58r4enhynI57GGsNm+5GQqEEVlZG0HRDs55n4KR
Rrb0Nx3cjbzChI/hhsGTILT7M/7p5ccw2GlmQblW4Lj36E+I4LgQqgcn1B2AxXeELfcifMJYYOi8
EiKVWnF/sdPx01tw61EsxzVznRjcP0M+KW4x5Fd/AdYh4Ha3jIJjLhbWu2PG3zdWk8VZVvjBHkNe
fLBu+4wugZJT0rjT4amPJCQaBiXNc+o/2GGd0ZuzgrW0TwUIWH67jwP1hRFOXOaTz161lMR3oSRt
n7zd2DblL8HDZX3vPM4GrtZEE4JHj7JbS3DfCYrTWBVYBlTHoEMiW50cIoq5QC1/W1Ii1re5D3ZG
dbXutFfYmok7yeIrPw1FyPo5W0TMttA0+164zLIoe9tvz14oZiF47nNgznqpCBarmMorglw9CPQO
ZOZuuZs3xMMFLVln7h+5TCGczruHAr94sJtw2IgAK1SY5CuRSa0bWjrX474DQ/o8NNSaRn7bV2p5
J3S3elJAQ9Sxt5XQelcP5lV9EzzHOytWGXCqbGTHw0CEsLyZsZeoAVsPeQqsOgazkQYHtk6id7wG
MlNKJOGGHlc4+6//VmPI3s7STfFuXelR7st2T3jx1nB/Lp2edGdySy6iQ1iSBGEbeWDkjSxYBhad
d2e23hHroAzMh0qcwArwgmnVyzSGBYstnNn79wnkb9J5GsylakLsrI3m2uAxlgX3M5MrrG1I2FDD
58u7ZhZlNVr21DN/VWSRJTZ7NpYmkLlkBxnc4uHOut2v0KbHjSN/lqasUN2J/y5rxr0pQqNy9dzp
s4LG28IsMGWfcj6bXSBSQLWaw/ADJd5A9DfITCL/v6B4ep5AS7tPEO3Q6ZhonXIack/YRhU83Pcl
RYsv88Yzv/tuEKvoZrUeMgMvuaoH9aCZSxdxVAIkUSLzhX5AeE168fPLMLkw/+LPzSLH8rdhd/7C
LjvpYlqCiJu2MY8Mfr9mfl7KXH0eMC8xDdfyhHoZeTPgRGqA8xyR7aZySqFPFMhAFj8sKdbySEHB
sF+u/SBJDWjtVjx3L3oVBoaymeQKvX5nLMD4aSKX63qJyyriCigdSdzI4anKg5xPrttI6EWzNzIM
zBDoKNUGTD4QjKlMTFtVRNev7ysfMBSxHoCLqwQpsjpj2NR7wLP2XrSqS0s3tNll+ue60Yp0aJ4o
KF/aYumX9Yz4ojrN/sp3L2LwMDdi1/AgoUUzgZxtDSU3KTG5knh2PQ++uNVMYJMcAP3w1e8v775C
U3QiQUiRNPo5yF3DKN1KJWraWfdwKRIvx6bycEuCraZ3NkvqcneJG8SoV/zlJQMcm9hxfkssX1++
aOOjEtGG3fq2I+u6DDtZF/etST/VsNb2RWukkAEI0Whbq5OWS5wgje/yXvKatF1O4yl+K+gNmBxp
Pbn9Ow9hXUbjo4oC3kJLFbeda9opv76Lkr7VStEaokAD0J3TSio/71/DsewIzuvTnts5oYbSct92
0zQ1s8aomeaRwjPxuB3u5Om6qb6prkPSkNPsUsFi/zEt+jDVrMGHBoUgbk9kA8Offi5KLhoidE0a
L121rk0XuRTF1R0EL1aqN6FZcrsq6JCVacC9pSxSixJi+Y+p508NZYguleaenGwXCevoxgNXcef1
zWoOZBA/TPize8RmTJ20KBQmm/nfVLd1Tlag7shaAeXFYdPfbyPFwuT3tMW2VsW5c4rqEM4jL3Ob
4yaILEs5ByunoCmDxsNsdHmwko22R0GEpVyxmPaq1XdLlT4Nly2C1GGjRLl8X+wnxN2BUH6COiww
ZVpKUjvfxh1f5jKAPShdmXw9FRdp9UKD3CPnd3hR39bLJFgT5Me1OiP6Kx/Q6lA263qfTYTj34zj
qH5fVXO3cKMBchfXBuZsMHgcPkytwj8QWFtIRlUyQno6vYnRtPAeSLUiv4oS19z9ro8Ss7uAqgIR
uoWdrIL7GJzaw/iHWhc872yFzw4c9J9TZcvG+WmPTAZP4zEihmQkC738KADPrTjvD3KXIWZ1q6Je
Y5vEFvrjCWGnBA+aF9XK4PXBUy3c3poMes3tg9iuvPN/ySJXinuE94nnlWY5VfmuOnbZ+agMM1HQ
/G+q8pQlbU154HKRIJNHmuQBVQ8c2hP4dNBCd3/CM6JvtbCCppQ6bS2E/u8bwaNfTx7sPu5BztNN
YkZvkqt0Rzr+14AqSFwaBzThA23g1H4ie1CcS8AchC0LBMNaTCGAyLkNUxhHPgEjDD6y6w/mIpGz
5Pf0dd/S+cwa4eT+o0k7yH5WgLmqUDqVX/oh3tw4fW58ngo4cYISBZNcvV/dRv1WgipnyYE/arK7
zSbvWoKXCGjndez66E+RxTZB1sCwxtN5U11bfONA8WWFIpb/nCFokX+FKK6kf9/eN73qlaSFhB/B
DrPGc0I3Fwxau60rKh4XR29A+FXRdWHb/4jzHvVCnxh9hMNl1dJgKCy42TR1+oxuvK6mhcrk7nRT
WteeNGQjSjPe7ZYo0S2R7PlG0GfzEXS47K9CmLFRsy6TCwv2X7oPPs5wFKiMNRT+pA6K/3WF1aCb
/2POKTF1MwVdrrCGIH9NTXuK0xW1ADp+p99UdmdSoQL1CGo4LelQ7Q5w8xa2OFs5vnOTii15IQ/k
IGbATz9VGtjrEIUY8g45LlTv2uD5n3Lff9Y8vV6lT69orEtbTl3TyXH6nnsw3gQaz98z8UXmGUZs
kbb2IUgxWOTKDklUDXNO0wBOp3MkGY4Wt8KWm1OgQ/yeOsA1rdm3xBtqk8gR8OOIIVScusFpCqZb
jwNAGUEcJ9PotHqoRha18jgONTWe+X+zsPquDUJELor348RTX+1JFh35y/p9ukUWkfQG682xh9vG
2Qra80LU6rUbzRWtL8TwuKWqTqO1GjcV3zLBDSL1DrMIuTkKS5JM/Ve8ccXTnY3R4ru8GLewRvV8
ghmqu24bbae0EVQMF/V+Yo1a2ouiR2ABkNrtGP2reG3RyipO25fhLteSu/AXkR/QUXnDNQNXczlA
efYiCiDs5vu5k/V+Nf6rXN7e6gywMcOrwsIZSI9iOB+vbBDfcVxL60WtkSVDKIFrlha168nEJPPu
sBHlXlQDezgB0VFh/U26+kMI3sw39/aPAbTNeFtSPWDxJ5Ol5ZhvpLRVfkb5dK17yCZ0TRAMYlII
c9erzpRvl5W02yUtNU3oUHTbA1QpXr4jOR7lS5IbfGEWmX4FbFzjRBnDqkpDIwz01+YYKstJP6aG
8p7R2N5j4hFOSwHgiQoD0Sa6nDy+5ywFszKzVSTCLCHxOh6ef6N59EZzw9tIzHqX5PMcibr3vSmR
551oEe/WTuXErpua6lMmG3MoOUtYubQqCLfWZ082jSHKzN2y2WmhfbdrmE3+P9WMRzF01LQGwk+K
/d03ZsxCUIOPgf+nKRQfTVLn7ZDH0Ym1DzgX50QnQ4gosOToyCRyQM38N8EObbXJe/lKFslv+gt+
z4pTPa97ft/CPZ8r3cL7EWlHcQqaOBOTlrOD6DaOEQ4DryWwyU92JGG3ScMC3kvu2mmBq2TRIzSl
wL1Zlb6+BRwU2i+J5jeFUhQ3owtftT5MjGOTQ29q3evD58nS/XJmfYRktElALzEdBjzCMVogtw8Y
MWdxmIblEsw46JSbMMKiWTTcHJBBtHSUdYEpEwdvv4RE6TfSVX958dYune6sv0Zw+DQ3VzgOLsZv
Mi/IfJt3zzfdPuwu731EVyvxpDTEswN4+Ugi+US+DXH3qZ7ZY/3klqScK+/FLeVQwUL9Drho1fJc
z7Fv76EdEcNnaAcoc60vZTtK26OJMi8r8zHOay9KqjfUssJma8AhdOeM7b/nq5s88gPu9PIwtlKp
mT1mf7PghDGbHWB47kBY5Y5lDvBicFc55vnFfCabRTkGfDvWMvO75dwny0aWhYnT0ofSxOCaApJA
M6FwsYo7+hXxGCjefDajMVav22me/l1gTMksjGVrTz+OxBaQpch3S+doLHFjbvujh7VS6NGe4Rwr
kzoJUAKeWCKTcRqwNCOMop5O8yvmhyNHWhpTNa3iLfKPx2VXI4CnvIBeC1amqKABhzlYPqneHUeI
4HH4M91rIK6lc6uNXmvmat1M3Js5OSpSwHRh34iG7Reb1YykAI8LQedJ4iDcScJJ86ZkAXFpteE9
J7TKLzT0eal84HOxnTCbsGYY/r9Sgvz7nx1XOdlveu3tz5zrvJav8x7caUZF8A1UmE8blegabxDF
LRB1qSHQ55YJg6AAKyybMathSrwG5pMACDFABP+fbOH7ymgrz6WyXKgxxZng3AkhIHi3R5DWzyWC
Q/VuUw9MlS3hzZN1FT4faI6dDNmmNB5GNgaKdydXlJqEpQDF647KA3Qmxbz7w0k+07i1GlVz3yt+
rXgqmIuEPBehnO3AQuOmaNcE4QYlE3WJaojWj2PpwMATxctemhgJsuJdPb2Vt5e+Z9yybBwUNtCf
W2cgnmiTtuD4YIJQkhDPNz167H674J6KwStI/hBprrr3tpFGpRsnPa1P2yGJ24/bqLySoEo9g2jb
9Yg8/L5uVBSUEQYW9npLKeiRjPz7Ie0eX0K+IcCEl8/hldJdyiNWgTPxahr1ZgIFKSSrswvhETNM
aB2YP/Gqi8MhpocPhzFjOWutRtk5Y9P5Y/ahDSXNsOy8UuguXT9G6cynFsDTed3d4joQHn50DrmX
z7hBILZRcT3NnTQaFSoZ/eewIwa0vsmUM4cJ3H7tmTmXXVNR+/yxy5tKS2mybSsn2aYuc4V0p+/V
Ej8W0+2VwhiWMCk/9gMvu9/oQc0L3RJKMyxGul7XFULdpS0E7NYvKypnLJM7Qln7teFUjmc8gA42
OrhDGqfp7MHbF8T8XY+6rFSIS7lIAelBZIjJ0B+9qr1rGhTracl41amaNVcJBck73mJoGaIXRbbc
lUvk+VWHQdtmMWSxBpbx1UnVjVhOxmLHV+XzBu29uAMO3PisEwXLzRegWP/UfWiscwIo/Y/7THQd
ynS6hHRcp3JO4IRQHP103sdFNJ8er+gsrtezPml491ePHAkUKNiMUpaULb8W5lrUaFbNX/b+sAGj
00rGq6hdf9JLdJUJXVE0/4LZzS1bUdv2mizViTsxTcnuLT+X8FnJhemlPCuWttGnIGeYSuWC6VgQ
JwkONaIvF386jOiDYj2QcCGEDxZhsEUapfNuOXy3ms/IBR7CCpNiAnb6uokpvwL99XDtp11v3Zyd
E/sDt/87skck0wSUCyic3JtvpC8dTODrwUyqMW5vZUv5Uk9VTnX45zNK7jbJebWlIQFNdX7r/4uJ
mediyQ38vEYh4C8hP9fa+BA+2SUybqGfwBhM6K96xYJw6QvAN61mzig8h/cB23PeYzN6ncawUKjr
IKUzl79nM6TqV1fUWteoEvrs8dGbLCfnpKADQPXogPkG8wAiEQ9b/DGmUX23PPXS43YmvWL2hqyk
nZ1BOYlDoj1YNUwtl9LMMOHsTmZyqBY14A13BXCl4r5lSLVTCSDTbhj7VOmqLmg7RiHC7RnsBOgz
zPRFcSDWKf09GygoJIdYUSn+liPZTWp7ntfp7KqHCW2jE959epcBSpw0cmdW3yVYK2xjGo6/vUUy
GJVZJATAiaJ76+TnQ9Jm+M0luK+9NZadaBhiDXICWcB0VndZNLlfMNpnRQoebqSRCFvKHDlxmOKK
Puu3xhv2ZOWI+6FLiNwQbP6TaETqELWiTKsISfIQPlQprbl4pXaWqKqkDhuN1qUXtFI9jD1p6mVo
xLL2yzCbF2w9B0s5zALaAEBwEZ9GkUWv+At20nxd95Fr1sjqurbgCLABlKTU82vMVoP3RazYCmHb
7DZGsbl5X3Qx/eliilRqSyC2S8buaX83hS5fgVB6oE41YccIwADvyWo1BrUsKyDfDCHit0uDx1mx
yiw+1QWywwAdui1D5Uh+gUE3YTJRwPrEf/X8pKwWZ7p18v9BjiOXN9YHBrtwkR0GWBJjsmi4Ei/X
wwAxg+Ysd3pmxq28ZFkWFQNuGmvRdOqF1Jc8w2fWbYmgGT6f64X7+uZVeZMcDm6wvJ5P0Vsrh7e2
sLCoCyTNsMoz0wb07OGnnBkGUHaiTF62jxfVxj7a8Lol7tO6ewb7B2LqUdjJeUjK16LSy3l4Fiev
E73WpxOUccqdujsrFStye4r0HZKGcCJFeYQoKtqdqctTslkld7wijsECgFpWdWiJbEdZbCh+sjX3
W3xIf1lSj7R/umeGhc35bXGtpPpLzRpAH6huWL3eR/ZLioQYgqGDn1KrPwkqY3tEwVKILFZU1xk4
/Z9YDApJkDymbN9KP9wZHETRv4PaqBxmKhXVFJjG62DYY2o+bLUUGcZEF/Cx5Iz1tmEPs/BgAZuq
NGuER0b1WDsmrumPLYoRcUSC2/CvQnvs7eby+min19PuH2uvChqSJObzkVRDMBk/kitYIgjfrNnO
3A7pWH2o7HDozPldTHHAFwXcdzo5YJrDDaFokH9m1vU+gNXxYauEM/+kwJwqoH0NHPWPwIs4AjRm
vb1yqFPlgjb++vXQXwHI+Txewfx3jRBKYUf8Z0L8OaAO6LjC8abkiQAXT+Ts4l8zMBYU1WwUhbRe
d6Lt2Hx8Lwm3o0ISsc7L94kWsYrNeLOLmfjBokQMUeiseTba16W7nzNylmg453tVWuoMRcMaquco
GPqiFLdWaTlQOha0qrf69p7hL4pSpPraDnC3glO0dDS3iBMeoWae4ZYJ21YVI6YdJTbf6QqSDPKX
dQ59wuciEJdLzwstkaXTPkJLFoAcB2XZYUO5rVLl1rEO90+l9HRZTrzZdsJO6nmN5gSKMlaCODHM
OjDpbOgYPYjpAl3go2kk1MN4+ioXrYTOVmB/MKiN77uMsgoFemWMGszLS9brqsicUCjV5G+FVQFs
RJE3pOrirBUitwXLPext61ggZiZsEP1NUcksxTILqKJ9VFPW9z902QAyQ1Bvmwb2kqlpWGayHTNu
RuPb7FskgARdG/2EYu3PtX7/GE2farCaLzHdUEVp/Rs10sky6drsDdZmLJc3aqcVIGFPw9bPOv+X
cPRcEiX2XB2rXMH/cwoATQ2q0yD/Toxox86ZiIXS5SrvgmWxNb1TP9Tz+UsZTfQqoGEQXy62ccjm
gJbCeByeeAu6IYB0ZG/GFR51W7TRVAnROjtANV0TbM71AhHTFryfRewE2swHc36D4m0x7pa6MynB
Kr7frqs5V7/xOz3DS4cgUrosbauUdBTcc5oAAc0CQkI5qgpUv+Ysb5Cyws5S0KGK51R5mbvnMCzn
k6JC5Y2Hi7wO1IquvgBY2amYh3Bcu62WaiRpULpFDOyBKrdqRZ2u01qtyg3k8yVZvkwYuHv6uesj
ND5vuMP2yCm9SpOCXE5eXb/8FlOxpPdx3/i3YurmaEODxfmIpht+9TG0xXrdO8BBVT7gifLt2OtV
CGGsKJhXmJ0xU5aMc5znhNFtFqKN7Qv7hshKnUkCFUWgKEFqrguE6rXynrQIvfd4is5Yy2g4Bo0a
cIzNOWwvQKK6ymC6s+HQi/x8q2Dz3IvfnGCJOtlnAv9c7ozC3P+oAUlPOAnztZQgxW3L16fUcm1n
4yA3rWyGSolibZdd2FIkFL/0L/p4YXUKoejc1YRzoQ6ynVFIwKMvGbDYW/nHCVA5WWYfCsT6TWeI
ra3Y4BfA3L1zHo4forjWnBntgLtBXyhksuLWnWy2/53cq29uFDxS3LKJ+LQxvdhAWeuo9Mu6xwCq
m+lzQYY1tQCkeff1esvJ3st3i7lMy3TaL3Ic3hxLgQa2OU+6dJbIUk2BhDKVYw0IFGjCoJximShl
UVmKgsKhsyU7v8Yx8Z+scl0Ax1nwNtmcDTtLhOZktvg3HRX9iwkfHzNaCIclSbeZUD1e9hvbGW4G
J/sJ3Ocx129ONHpKoNzfiurrvKjkolSex90XTum38ojkenQUfA7IsGK8FQ+fm6Wa6F24W4i6tVxn
CEnXt2hUPEd5A/ShzJDIHguonykotYpAoKa8hY/tJ2Msi4jQyu0mc+wJ6G7arTMf1AaDFvBDC3Xq
0ap5+oJPhSbMBT+aOMM0h1OOguSsR/uEUiNQWQrx1B/IoPF+LGH31SD95eUzotnqJnimbpe4KNB4
TE1F1WHkesqOEk9oHAYlskuDrMxDHH8/PAKpUeGdINtKsWI8BiFrgjlOJn6EtubFlE1smKGHO9CS
KnLOnv1XcpUiL0Z0YDyYjeanSH7rOO8iZ7v09G0E4tjo8PuZ/I/bpRFvnhlc90ZkN6zsC+nYpUQD
/wUekO04XU90zyqJFirUeeLZTHfjcX0INA17X9gwRVW53xrCy0e463ExZa1Vbg0BkMo3GGnlAAxr
H7fKBE5AGK0Zkrqsbn+CH+HL6UPVQyw+rlf108vhGKN/KBUQo+7fpZtftNnUvaCsKYSewk75BMvR
C7YfPOUtkA668qv9GPDp8RsIGzkwN3NqQF/NKqiCtxfEg4ZqeoFqjW8ysng47wzP6cLVxKfCyzs5
Qkp8r1fvMFKY8nhhLvnfaQnfIUbcAET68Rqy6/oYKqSQ9dzIay4v2sn1qOr4f438Ga30SZRv6C5g
jVRInA8fPuh8c+fDVihkdYS4YdJRAnDk2R4HRkwDjMC1Dbe4MOkV0r/0sP/ykWNee+IlB2RxkEEb
xEUhCPSmnjfRli3dPUEvpTWUZ1jqXaNqZ1CxXKfzL/skzlvQ/l4bJBb2mKlyDLd3AJXJDUxxtCqI
2oP8WIhKQqHyfJdtGhcZSVmkmY83WEQX4Ww9gPGyuJlH55FjH95qCGw5V9EEUB14v2bdl2fpxp4L
p6D6WgR5pKjiWBFu3O6HemEcrH8ZPIRc0iy7hwX695f3RI2eTD3BL0JSkQd2d3uWNYmxevyv+zf3
EwC2XTMa+CUkRIogJ4rUqVrZtQqDXfIuG8Ku7oYZ9iZP0uY1AfZnES76/kwA6q8NeZajRge8o5B9
BWLzugcY/BO51J4nYv3q8EVwRFuun++o6OoY5nUSJNfJDM2c9/jkv9OP55p/Z42f5ai4ObYyCtZp
0pQHNP0OG9AOSQ63FVUoCRuKF+5P3nQFiKoOTAfYpisUjDZZpyWlEUIDT7zU0Py5DOWeeGubYXOW
7N5M7oFHswa0Q+74d0m7QPW2frVpxGOfDi0h6Yw6pMCcGq5loJ6PsANKBWvRFBVhgEbOmIELfXyk
zrxcpy5+TgNBsHS17ghTf2R2hULA0F2B1zapqs99o3P3WVj74ijGDVC0XuYXI3Ebzrn+T8ApDiow
FE6nwv9ICPLJW13PMIZlNkcRt92X4Cq2JopFQwyHC3JY086Txm7DxJ0J3X95XtYilmrV65EeniL2
/5Juvd4zGguNI0g/rU+NanqgwC9O1UYR1+CGFYxzh5wYhb64TmPImeJKkFAsJLevg9BatVPe6wjw
wnSfxR09DGxC94evAJmC3vEHxvLuy1Z+g1EKUVmyYPZPmU1q4JItXXlHXBxhBsVKX3AtVaS9aC54
Cm7aHV9jCGu+qD9Fc2lkzcsg+xPbNPVJAvbx04HEvjoGXlZ2bj/6YYBMMeM33AwxeFWnMq1Q6hwr
bMY1TXvVDjvsuEMMZKk05cmKdof0jsrcK+9ZSST/H6IyVJ0RDoTPbyiA16iJH3GlrVqGIU58GK/S
9eBmrzpuACm3q0cmQPna2nWd4L/1fxqJXKH9Zh1hgHtEkISslkoXxlH0uh1f+FKAIKCcIHICpP/w
y0qkl+5q6EecjHCyDRNkDBRmwqesc73FbBdZ3tPfMGvjStXUELcxgmw2N/9eXEM96j263Up7OsWL
0eMZDiauKd+qHF/EfibjsNE83VD/mocAhSGd7QVaBsexgcdnQPoJNnq1TRCxQouC4WGdcqt7zMKc
/EBfKgqdI/uyA4wQ1ZXCMsluyxaQrgjZzGo3X3Kgo1QviTa8vUzaARHZa/suX37O7ZWonNSd9Rio
/jlAfXRs43M0okfy92m/LlBoGdQ5tQjVdu5iHbtl15hoYb/6ggJrnj6a7CbYb9dp7Ml+GXVYbmIk
jvuiuLU/2lyWM3jIkKzPdrj0J4zOQZfcpC7wJlCBKoxiPNeAbBetx7/BQoxiWHd3SSBkc4w5ZBdD
semqOo3u6hnaWw/kP1BMSrnPuZRFz5g9dMTDccsb+IwphP9g770WZjI0e7tdig5ZdbYCWFIoUIPB
5Nhao9M5cw4jwDFBBlQGdm2U1/N3kLU9e4nLVheW+HuPUIZppV57X3eX8fUzwIc4ho53oHpPBtEA
wjp2lEEExQZAHwFfux7XaWMc3Z+J0UFN9prWgocvcyMrvuQo5g1JGSH/lC4fnOHnZOpthR/6gTPn
JkbuCgxteCzBC7rb2oVnN1bgU+yFYW+/oP3GeaWJYa8vz5WmAoWR/4CczP3s9FQhlCILg4jBAsPq
L78PZUMpoFkJtKCCKqGhOdS3uCxmrtTD+6obVw8v4R52whxMp9vhW8tQ/egKowG5n3sBDqS1DfS9
s1eClFT+eHxh+xeubwK8nQlNkzErAPHcSrFOq2BmPVD0X9eSpVfOvS7D6gcwXXWgRMX9gZLqV1bd
uFCLthZwPg+wE9rHZbIrvSQxsvvLf4FKVnaMMQ+5y8VpQf22aJ1fpYtrYG0oBjQLSpYZUTkKow0b
sSSu9so9rZH6vAjO4WSa0PRPmIRAVMDlI9fcNZKpqlg+rt1w1XbLaIgcnm0z5fY/+MJIT6ygVeaE
XpvjKwnVwvWtVBGK17nQluc+ZBs+0/muWWvV3svMxl+rxrspPZv8b26cJfEXhHQx8wiLxZs7oLIF
UxwiEI7v92c5z+kJ4SZoEfunisqjEIP9ibqHVMLiuGnpvPYJoQWr/kcj7jgxBPgGYsDeELvadBKn
CHuTwG8fuB5hzxj6OCgpRDsxAEafUUG5gu2ycu5XXC1UmwsXwnYf6cdL/2YCn1lYCOeuU7toG44O
PqZpCiMqDHzNVurZnSa7ruPq/6H1AgO8ZOi3qe+A9n2fAv5tlUs5FPnER9rEG3rsGNG4LGRCfZ0H
zpX0MeoJjPEni72QRV1M6LGtDV7Fn2UqdYzVcSAdnOtjiwgvP6slV73CGHeMXQ0nTREIPAigWns9
mmZqmOYHhcOCzx7mZTSTytMJi/byOcDb97IRnIk1Zw1gvj6+ehzFDcSl2k1fQ93eUsxp2JFUED38
zJ1rFUJNlG9g08OuBvnb9UfEpZ1KyWTFbxzUgxYIzuJ9zXo6P+P3/4qrZJmRD2CcPNUSjpCSIq/j
DC3N+luoRpzZvEaX0a6sLL+OdKCKV6Cz/Kw6UEeSSKXVmnuEyfqQ1rh1YFJipk23w1wNBHR0Sl8u
t8jiBbE33L5/USMB4fjiY1G31/COO2Qch4CJybcxfHd2Pi7R2ATa5EomtXt2L/h5aqQi/Ev0oSgx
lG+++g7eG8SefqvOayCq1UHI4JDL+U/rHrHn83Uq9MYuY8+cJcQY3bijAeSPZ8RniwzP5ttPkUtr
5eZ5SL54YXAdq0dRY65rF567TNaoy3/aURZ7xYNoe4i2RJd1zeQCHpKS1yM3L8DlevoH0oWhD1bd
W9A40WxM4hjKBrLxCp/sOlrm7QKMjDXiFlTJvDuPx2tcXg+j5jQqY5/nultzyjgt7D2/nvnQKuQc
r7xGAAke4J8RQ3MUmfTpV0PeB1zKOQTGGgGp4ntnY+WpeLt/R0onNV/eHkgLu8hptft/RdwZOt8T
HVccG3/zoRH76zceuW6rLyvIhk9ENPOO8NjohdozhaHYOGEHfq9tTZHCzb5bxrBiULxUfUoZr1x8
clnvXs0beKRUblBwcK2qgVC8cluR/D6bCuat5EFDsoKT+3gu+/aH+qYr1wcuPODl3UUeg9yx2Zk9
1ce/QXeUAKB4GXQVw7WegjWwgzyepfkyoE8xIKbnGtWVopZ9wfFkt2nmxil4AJjBAOnNxUwPnVPS
TZlbdTajKoUKt4iqzr0dsXU2LJgByIWxNIv2rzs6hTEljpwkfxXegCJYQuRteIfbwxh9InvjH0Bi
xhlOSHHut5nbucDiGt9G0Q30FoOAxGNt0VvOF275Ovrk6iq8IfV0noeeJXeBil795y78kWl5dNPZ
BUpn2DP3E7DQw2pTLqqj7fQ4n1sTj94SkEmsYU60fHGs1wlXFBdXIyOzY0AZw/Bcp9KPWxIQUu+C
7a35aa9OjtHnUV8IkxbciviCB6SF06Diu89ez4uIEWrP8nmQ5yIN2rI0DrzAZnENIIYfdZVYFzIn
ZSfRZQ9sHd0MWC+Rl2RRKNvmZV0egEm1ivdpdTucfmQCgHcZIjdBUrzyKZx0nhi5atBH+Qf6CZOL
iWOUt2R1Kmb8ZfOiJUvcMkPw5TUMD7r0LnQc53ChiTbWnp197v8WqIQW7oQm1RKoAQniuH0ua3LR
F4k9Yfj5DwII9J9qDfgSU/B8aYlUDYeMu1Kz7JTppBV+GvUGxmM2VwxnaPyK0VkBidYUFc0gV7Hw
PLG2CxuAZthJOL/GKnibI+azoqCUW8vwkHMDlNEfuSD1QCNuYqLBZRYH7XID/3FRQGsxgEtZMg7B
0/UMhv8U49puNDaUdZFHYy+++YGzl1NYiNkvocuMoG5jKCtwnW3Bx60q5p7IRBSatZQ3E/hd09Xp
hGGQTEKInQpXT40lC+8cXx2eRhj7SI0LpwxB7v/4C141+StTtXxHk75TTkuUs1+40dzB+DFpZ46W
OO0lrfo1P1MiYBSoPSfhWov4i1CTzDPkWtpmN13Yzln5vvny3EBDkUxlhY54tqVqLmmTIonDh+Xn
Q8i/uKJhxjdGIz3lxOG4COtDGAECZOomFOdctGSl7GoxletJYV7dSY8ftBKTVkL01SolDRjsNy2P
0U3ilX6hq6ImVDP1cPgt6P05rnDUyoZ5Riwd7Gkt0kVzC8gBbyi3/Q58n5XgO0DzUmIRb2xeM8vP
6pLXrsQTIci96FfeUV6jHiGU2eyQzieZQ9tbLijdkBXVhJ9u6E27Cy8slnTzGsK2RVSHJNcyTWCZ
KP4OIUEVdbtc7POJoxDUIJ5SK5v1JMzhwMwrL8vNb+dnIZOx11n6ELHpHnQuoIPuBxQg2oj2oqjQ
iN0JLu2yGnjb7gDgDN6mIW9V7bZY5nzy6hRG+195zpJybq8Zi1LIXdjSoOTA77zntk+YvEiOP/WM
Um0f+HNaGkLpl7m0EEcZVVhiPTNAXUZh+380SBLbdzpPO4MmFxvx64cjYVA3TQaVGrUnHokfi6hN
OcelsPlYCLEQ9ZoGTGNcvWtDN9EF/VPAe5Q4vYhAj2T2Orc9OG+D7kenFQXG+MTArX69Kz3kGt6X
FvpolRuCjl4NiXigl9p4IjgFEM6sWCEC5TFWPyRx5vcVNzAFkUHRXHJUCOmsxPSt2N6BtXosqHBK
TC2onbYkLZzoj5MjrGXA5KcrFkpRNWILujlHXxPz40FOHWmvrBqkhFOc2L3wC9LQLiL3vYHz8fQX
BUzHwYFwLWBqt2fmQkfzTc25gQqTZGw0rVPYgEnnj8cK2spxb+yBh6U6A+bTVzksDgb5t33vS8yo
zZJ5JcpDT8eHup81lwz0U/sdy7PqriE9dYvYDoeKZZ3gk18RfUx2AlKHhml1Z/HrY5QCp7FQ0LLB
xJWuPbV0bfkcMNnugq6LM21bzUheL846ty5t7BEmPqxepcLdRYOyZ6I03MJdJjrg8KwM21czeBCY
yrPQgygWz8sEaEezZ2AxBPq1oSs5oaTVs7vAg0zlzNY49D4QqapMI+Iw1P6GyPgskmXLAwG66Bn3
84U0MXK6sq/fT6CFK0b9sWDQO0EmzarI2GQuJCJfU2xoGuOKplO+w+bGWSb9xLCnp/X1Tmre2ayM
ufIiJ1zpgVRNJ5oFXFKdWwwsyJ5JbmZlh47uDh5aoRPAoxs/JjE89MJwvUJPtQFndQdH7RPrZRtW
1/F+M0tNvoAWQDiWRyh4I3VmELhfiwPBjzvJfwbFCsrfu/optWU/buh0zueEzXXB9jpPOEmDAd/h
xiqG4lxfm38CQoYPdr/MGSOBZI83TcT/1L07sjb5O0HJw0niggY3M0fQf6qyRBt84SG6HQQ+wM8j
qFzfOG7qwwnxa80cAB4h8tdXtaz7/flL1oajMlpa8cHDrMZ0y0INzdq4WsYgBkuULLt+DLJ5xKnN
IgxTA8xQvH3DN5dEgyrB4m0EBaAB0SsuIcTP4/jFlC8OpFWUcEVTVGxokfXpn+wVpHjgDBmXLSZa
2Aa9fCi8Z7ofNvOUhrIU1FNldFYBO6jBBOshSlaxSxPj6BqlWNOy1nD5fObJKPzr7G4Acha2IobV
H0QoxXMBzrqnS55m77ctwK13hOi9mReEBpORSinUJN/02aZ9xHh1ALoAd1kLI9XuLQxaoBOVSreL
l5skv/QtkQ2QLNhPv70PoA9DEc+xsiQxIkr2OBdVghDQF0qs6lZZtt/0IYnpy39v2T+ODcrsWNR4
KoGMwzhVry8r7byI4Dk/rjalFmzroLTgyQH+voOM3s/OfY4whCAGjC/5kOJJGrgN/SQ7ubfg7oYg
zE60okFN1YGyV8qRsDQrugBdDb8CAXRq4dbUN3y68imXN5iXA/QUYDlS90cNF7XsDy9tWnV2HDaB
bBHjaXjARJQoIdhmkH1pCvP61buM+sxLAU2+v6ftTgiAuBxXlo++d5oHL9djEcqgpqp3jgQ1w7bv
YiIIlEp3rjnN3a3Jlj4+kCibrOJLKbvBL/7DMQMTtkrFEO/WvkfKYcRTivUoJXDqcYfmyKaY3B2d
kA2wxbl4OqhRU7BSYi2H+ZH1EJ99ErzpI7TKZ5B/v6S+JqiBlOFYJSOe+lrCtewQlb1Wbb69/eok
ZzX9844SHC+tKQrsBx1WltVOdKRRN6d7rXeYva1IqbHPhjv+J41kueuAz5aYLPRpO6UGWm7m/Dxp
PcdQJs25UCpiSP8O/DehXoQLb6l6eIi9x0cmOANvB/lB0+h/Epz+Y0bjfrSFnuBi5KXuiAeFS4bU
w02gfExj3iTwmbhXZKxiR5LpvoafyXVzXzkrGEaY8ccrR+FBygM9Nyxgqyzhc6KY4DCE+PVifjPU
uW7NPYDv+4OVtgxzYwEosAeZRyPfXnHPRQ7nYcVisIU/ZW6JnT3W5sEg/punkWMlF/GY221KD7qe
ckUqt/0Rau+2Ne4sHv9l/u3qrwXfhfXklJNUgZRuJeaxlCKgbn0+GgU+y+HfCbAj3HNSIOtFWyJ+
jLCTqtvU/JbivYbKRE+QSkNhscCyXaTLopGoSsgut+zG+5yQA8i60R4G78aLfeC6W4IE61s++iG1
ULvMHBDGh/YfzxG7DjqyjxDQzQVmXB22iKxlaXMXmEimlHmUHV1elijHJ2MONDG1GpVPhdebpDH7
gPUcdKcT1yVkegZaBSGw6WxOIcu+PPq99w2Bj5UH2LakHsdkIdfZ+9yBlh22JeDD3vYAdQRRgU+0
EzgGLd6LYFsSQZRm34Jp3fjuAEfJstMxvkWE+jkKb754auSv/eGMGc0a8l9E2+RRK5c1hzh+FyXq
H7Zq4nI7wdcNKnDF5mGll/Bvg1img0VPfgr69pjO8l5AYsnJzM3jHDOMsBYp8tB81lhO5TRWxRow
7NOieS+QMlTTXQ9yRUzLah1VuaSpZ6odKhnUALcDi1Aphso9fVsP37UjAQ29HMh27ev9i9A+QOvB
YP7wlufvuRgr0yfhrv+0czBV0xQNONydLPMzGygfIGyQ+jNlGZKU4tU+OsfZNEbOJor5o4xXl2OX
NyhhdyI1unEVkOS+SsLlmBGPOe/8pwoCSvsxXkLQUJucKmn6mzUBRXTaMPJI9PLp1Re9hB15Y1aw
WZBQ5LG1z4B4LpDMrzj8ksCuj63FVdVfYY4Nla2l2NMhbgqOSqRDw/Mx+rAnn5CQOiQn9kOWU63v
rgypLsZJCnSHxZVu3PMq5IcYuGKY1V6Z1j3I7bCrTM9UrASwX7WibtGY5wMKH6o7hLF5EWNbYj1V
vgL8QGTiwmrfDA8sU4qy76y2gEs1Z1AJCKE4ndpCdBt3BHwwRlGkgstY0v+7ZFo1XOQBJC2NplsK
lasdDkh4hRDwEJWmiAOitJBqGidmdG0htwmjjNYlXsnOSqlVgWP245PYqe+UawgSWumqekK8jzk7
2Y405g+DEWqtCfut2mNLnK8V4ACkTFi1MbesEf66HBDkYZPZg+m4Q6uglj00gN9f5ceIFEsBaYsJ
/rK1QgrcpuLWvZ46s/iuH4tDZSAsi11SQnrSskh8fpriJbNV1f2TsfR0vC5QYXetkNXwYt1uyNJV
iRM8OQSJ5bIFD1tCUtkDtwyWmLV06eYX8RxDUS66VZk741ECxvw7p3YuvJjwrwzd85PemTkqX2Dy
aMnPM2cdi0D2nIldMniSHt8w/014rA6HigURI5QwjFmKqJTrrCJVzxPglNc34tpUY2RFsZ2CW8gm
1uqtvM16nhE1hsRIPXu1BjdVFRGFif/sVLVd2BFxc09q7G+DJo9ybuLTYhxCt4whP4iGUWKNI1Bt
WehZDwO9taI+j4SOHwbn/wnJqKyWoVhOfLqvouZL+Svxqsao5VCSdFjY5EMtWFAhg787k164tj3j
sk+jo39bxN6xImpVNEiaI6zTrg41Q6ojBC3oXnth2dFYIaYwQS+4XdvdyOFwtoPDFNnGLlKJJYHu
y77VNxJ+nWlzvTAmlW9mgqoVAyBZl98p8tpeEcq2+cEUUAvrhYa2d1yVWBSd860hYd3ZvGAw6mWK
gpOHgy19Y3STyobXCCP0x96JBzRx+MPQsgBsu6ZQ7ncwD4SgIe00VDEPlLVxhVDgdWkwlo3x8Hu/
qFjHUmwsAlgLj1AZHSoH3TlPgIfhLY7ymYECWfxkPvJmDoFigTnGu1HbvHN4xme1YCTZ5qeFvpb+
0TihTC6wyVFHhSIAkY+44/+w5MJgYwrT4MUP1gXWhPglmcknt0AXCewMjFUCi6+Koo+OGOg15sVB
hhbc/vLLNdJv/zyhVy/vYfSMCXiABpLNB2vNalfKD4RgqkYS9eaTF6xojE9U6dJ1f1HVYVYDXOs9
gzlmyfgquylpIwH+TapQuL1q5XrFzIC5SKBbzLbUx+v5hx/rKWr/VjwYlBnUvLxOj15xLeRGdYEE
v/b+etK8SPSujHQPdVtLiY4Auw8bI2uo0TtmIb4ZQqxOJHazusZqpVIs5CS7sXEerqRHpJp09Qbi
Fih5H5mTyWy8IOg/s+44Kjikxdr7bj1dAE6RUWkBNrA6uZz7eXkdkfq8QWbYG/K5OuAi894WJutJ
bXFk5JQDcHT7fD33ppwNi1OCPgFtjEjGQDdc8cyQze4fLN/XC9yK1pMkPpiq+BvuNwxoWFfdBMYW
oMg6hp+8Sd0g0ZH4O4n9NInWlLQ6UZujAAutcqieXGQENVU20gEV7nuJ4vzWgLgymDpSeJ56p+lP
kP1apzojXeakJc9XHxHLe8Jl+CG3sLUHEBDxOAgm8cTpok7pe+KTfn4vnGJPeh8kN5To89bpvi3P
w5iRPsH6j3zkhWR0QgylomZsEgweBg3ebNMZzbL8Dof2L7/CcsVg4RrZs4aYFccCtTp7PHs7m0bH
G3uXTBmifBSgoTb1BiS+u25gevKWFUGDAWAAS16BEC/x2kipfXbY/A/eMuLqU4Cc9ydxoFf+RE9P
SqSiWZgs0AdNMHQ065JXLJ+sAZkBdT6L+MGfelqnnLQWj2GR0Mh90GixJUZQjXQBn1Djr4RH0ZLk
HmjUk0gGk17s3BzZ+Bq1TlRN/LBOEYLxSQOCQ8zuME4luy+RNQqiMG278OPO1oVA/aghR7LVcOEq
YSWHHNLEWXJScOE6yXi7w+CFUMQlJQpbHlwrJ0rLtUk7zcCD67lnDj1BYnKUnwP0Y8Otlf4T/4K0
FPHVEh0ph/oUcwFkgMu+Oxb4ln4W7l2ZxRmU4qkcMwNgQVilW7HqX74WQjPE5nNOkjN4P4Wd7Qs8
PQ78FKjm52zLLbNghWQAQOdlZHG/BGbRVZNzu6njQwXA5p8ewjAKETKKctPCbPqto6QklDg1/Z3R
YjIIFIy+kkCnQos/8a1SINl7WRK1Aur/dXrTh3TlDnkJFdGf713HuC8l+2S/TpWBEfR37LiAJqdO
lA81j9W+kVp1El8BPwDWt2neGXEvpqgYHgCGW4rfkDid0/UMAqjx2V1mUS4qdnefxVwgonO/VZcj
XEW0NBCufHHaf2gslyjtaQwRY+kyz1apdAML16uE7Ii3hwI8923rrHbDpHPuHxSJhhn7j56aXNM7
OH/sKfpE8Vx8+lD2jIzYF2OYhTSqVhGyHoUkIYdlGRA0cgBi2MdQp2AtOSEDbmsjWeZ7aOMabYHa
Ba1LBkHd9Nj3od2+4r+8HUv36/GY5xytODaIOfP5OxIXqvyUCjzsnz91Ckw1o3+hJw5H3t6stylv
r3kHwUFImaFrkMbe2egr06iRm4XlPpmKFea7PdzzToVL9q6LZ7Rkm+sBWnTNusmmaGWPU+h92PBD
wfg7U/qI5hUtw3gqW/hR2LAYS3B8nextzHR+KHzidLxMV9M4F9UodxKOiw+kCyAVw0/SksTvN4CU
pE5QSOxJRLxfiyTUkbVE3EP89swSDuRqQUlf3GlY6BE+Y2rs4HHx2rFP3juMAgbAxWPHG089CYM8
a+7H83B43Vg1LM6FvwOaThlB9rHGh8mqUcOqqqwuULuKFHW+cipMKGZoATCy8Hf6dlZ1BBc6FJlr
LJuArecdlbZY+hEf1s1c0eRswE2lC1ASimR4T/HBfvuKxVqBeT2upMlbw6ZstDGFfa2dKQl/Dygr
Cvb0Z9/pyuetN2EyxhfTpj4r7e0zqzLeDV8GR7Cf2xaxhNKI2Sp7hmKgG2XtRN0gcYNGAxDcRJ3U
5ADwISQZyHM/pWPIJLY0+z4zsaJUCg9VtLzPIvCVANNLogH2vv8QdslennGvkXK01XA3d6XFqnEC
WYlhXzWKxIcHuKnZvDWGpjP1hzeaapEZDf8x5uN2WUPhsAqNffbTS2AMsSjUTgU46oLMgBtgo+wq
Wi7Uk2qRXR1Tgi7f5DeN59t/AJE8/V+zGNA6EBwXeSZcyDYbEnIVTcithTe6p75NzIKOIkE0wLJ6
5ydV4Mglcp0zIG/bbtXA/ndRJMlyz0CfOn46fwyfbMf2WeNJCMzP3PkyMyWXK83bHJoniQS2EBjg
joNH2rlTWwro5q8Odm5CWj987mvKpMyNnIV/xwCy+zrscF1IBzMCc3JI8671npM6bBWANsSwcRs9
W7uCZ1sNgmR5Zsra58MxRvv7f2Efjz/P7KDFR3/MdG0p5kxbMFoW6fATgxixPBvOMVVZwbILpymp
BHAiXVOiPqF+GdaAwoI435iBTBybUr9VGPEpy2C+emGd/9UpfQD+OgD5l2W0WiQ1/jaK0trE3O8m
3MO5Tl6Bkgkpdr/ey+dQOdLDA1fMtygIcqe2BB66w8D9aUgIts7/iQ6Heem9sZbhnAlXxErCynkV
z+kytB2KFGJmOqiek4yVlPfNoOOs/2ei/jDCnMUHA3e+/u7Lz4ljnSuPjgpaFNs/y7BYESc3oEiT
yuK+4zn5RyvnC669CA/n+vYjTrb/+5tKiUrSajK8Mwj/fjbbJOqrG/8XKXQDlKsQUNsbKhe4A8ZN
Jhu1FUMQrY5K/8DiQ5dhV6xcPNmrlSivb1pV4aGeY6aewsxmKBwaJzcq8OmF8+44M06Z13GMsVvj
3HgBTC85aWo1FBgI/DvL5gsvA0I6+gZpFzvfllcEs1NcnLiD2jv1uiuVe4sT21Lvz5oyX+vvxgHP
tbtEpBVJ7f7d4FWgQYfXK+GzolAq3GUw4wrgXt7KUBNnQGYAOMgZc9sNuLUEdAYSgc2Y5sgUPN8T
BEo9dEHkcHy9IFk4GE8SjQwexOKmUBzfHIEEgOlPl9f38dnsDad6Srd+osyLjOhHJ2s7s9M/+Lux
GtJJbyTeYi0wWW+sSGNJmEMljb5JfUYK8S2WGGnHyEPD60e68ayyeZKHlSpX4hALfYTe2k8a+8u5
OFuCD09NNpzQdw0W4y1TaedK9yUkGr1Ed6IliPXgTY1WuHIrFKsjOVOIU76VUvsPZTAneeQ9oA9m
pZVuutiAsmUoKVVbPtBJAeSCVdeqZc44CYwsGl5HGGlgD2FU6k8AiVmJ4C9f3Xi7JjNgFiWppjzl
KBCaf5l+v8jA1tpBP0Pv9F0qZZC2ZCVho2xXVnQ4U6QAgZccYxm1byMaQfrF4IAGGRNoSuMQR0jN
CrXYmSSWdPLTrt7EZNa6Cp1XAKTUCEv2gYB+fMEqeXIQtmUzALYaBPXXC4iq1/RpeO5q52etZw5G
kI1FyX5abN/siiPHxOavwYarbskPOCx2hVVTOAN3r+CH1HXGGOJHT2KVn8K3icke+rPydJRM3Oub
Z2BgHPdc5pOe2JZ9A8rBH2ijcganrRT2/Kx6Z0K8tjiguJacOFQ7Z5zF+DdF+CU2sHQh1+6+vB4R
/puN4gnKoljzJU7PJpqG570G1G65Aah8DDrst8NwOAECHgb3pLyyR/CEI6U04nqTFBjeBQQAieEs
CW/DYng/Ye1fTfH6r9dHoun+NEsceoALq53GzQiJI0Gw60PamR3xDB87JaRjK+N9bfEpZhUJTF3w
/o+ukYB1fVDfAbU5nrfrVn8azaC7Z4h68hJXV9S0JFZ9iGu5TxuiCXbC2K6BXSOBijRmYE734KBL
QuaDjexbpwfpQOc3qk25j3wfus1NYdC3Sf/h3obM/gtsNMRJZh62Lno48ncjWYh7+4opcWqJQUTf
K2US+Cx9YKBtWuRXgzBjUhl5239+Lt1DGpLozP4hwFdmMLGYwsjKqlwwnysGouDZLTBxDH2KAk1q
7AxVLj/w0sW1JNb39SwskfmtpNIL7WDOUmm1NwKgszudFHg3d+q57uwA0M9RLN6pEnO94L93E7bA
+eJFkwsiJXQG9TNlgGp8S3kuuG9isV6m65EDHrtM/8a4m7mpxYdI1vMOsJVAZwJniSL4lSF634sd
eHp+1ywSnMqU094Rk3ZRKZNxhaesBy+2RvUlLEFYbL0bd/IWTGI/yiq1ksQr1MRs1kNjC4sB8q1+
5eKyAfnerypZHG2gFNWg+lFKQcHS+k8n3jjo2HJijuhndiyJ13bNY44sI8ArOuzGEu9x1617L4UI
0XC5YfYOEE9iegDECS2XiHVxZCWuT/Qsn4ZQ4xEkYo8v9YNwhdlaQCZmM3+bVxeiPvCAGhiQglnO
iQWz2SKF8LHHwdvHw1LF0lrw3N9uMQXh2haY57jnd0D5+voKYSExSq3TpwXNx5ZNAmrFI/9Vi9qv
rND8zv32LlEebWmLD1gVnw0caNL/u1GVTwtGwDBtmdndD2nA8mlNuju0LzczidTP08F7mYh2v/8I
BQgCazzVNgOSOvjs00/r+HnKdE2ENuLr6WXsH35eWceScf1jK7EpNhu/BqThf0pNG4/mrNFe7v7f
pPnLsH6ZfJ+Oy+T14vCjmi1MR9Yp7KlXjEZWeuSzcftMhNUdjNzRGdetCmOO41z6B6ekxLsQQOin
OCKBhVEBRy8GbHBsk5RfED+6J/S7DoLunLzIGGsGVChdzFXa2oUj5qlAMW1S59blpJPNZ8xh+xzN
ip15LYTWSF2IPCZVoNiWBoBuur1wapCoYxGmYRfeghofDFA5ZKt2Tqziz6sZJFoJZqwwri6tIySp
3DMip3XgXVTsHM/vtznDCPlXjzNnOIgjdElGGqiiKUzgzztHoddvFJVcPuLACDC4f/8S6OreIV9E
ust7AwUcQphXSxKM9H1dfIViylO9RWGKiURBvP12DxDk3+nmMHp/3vlsBsK6O9oqNTvjHQXhnHJ2
2iUbqUdiL5UrUNocmpzK+zNbsai/seT2imHhbvh9qDEZJe35L7ZqylPimvtX4hF3I9mC5jLzu6TF
4TF9gEQDEDfdzE7+7UHIdc75srjk8YlQt1L1H4GjGpBaqhuiK+ba5frM5MMHl26/8HVwKBL56bme
6UUoZPrPVu2drHOw6j1hfWvgrN70XZvgIC7UjmVKu9la1HRS/6k+Xhy0Jlc3mb9JpdJFIQjEoApP
DXsywn3eyFiPE/EpeW3k1kHvHeo73VmAuCChwtW4ddyg0PFAI8FeORsmEBV7ERavoIds3NzjbW4c
QyEBCJZ80x1dUCBxJRiAuku3pLsUg0w5TsAUvHjSTaeE6b1rvaP36y/p7yjPvonHcXzVldZ3STr6
9tdOtqaYtdmzzUDO2w5CqeGFoJTpvc3mbwLK83STDz7JXJta758IcGjKhEU5PIRc1iM0AJkNcdqK
zjJm0LZjACjOTZkIU+zfUqEWz+thagV+Ogp5Tu+eo2VINKJp1qZdB/UE1uEbkyrMMLz5Wq24DB/2
xbKOdZ+jp/nRHR/wm79uzloge5vzbRJgipwjBPAM3sBIQEK2VZNLyYHDidYO3KrM35m3N3J54YW/
pxCfnRilqqy1B8/P2ExbHkTDtc866o42L9vbzY7vK0MQzlcnvbEyMnJJtSyvuGXdMBJMtFOwFaRd
TMN8kxJqqAXWfWnbQ5+J2doO6DeC6G9ZwQ5FUEDijvO5eqFvzP1N2Y2/oTjITkaE7Yhcf2d1/L49
Nk6wXZxaV7Bs0Ea/GesNSu4NFGyRcWr9/EiLB3rq8YQF2qCfmxungixBt5/isVBU2HiaxlAZLoyt
pJ5lNw5pd/e7LxVgeDAMdi5/yPzSH4MI5G5w8FULQs8QFmIK/clBP85C+Ze5/uaC7UH7kNRYzfBE
hVXc8QSZfuR844ojpnQ/bIH3N41ghd01IGSXb/uoDItPqsthDTjfR2VxExRh9PsLNh1auXTfC84R
MiSGglin65IaKTYHe5H+IhbsEJuVGnNAbRG1V1YcbY/aCJ/6XVvNY3pAKpX5EuVae/BjFi+bxa5M
/u/Xbu8NXLDrU3no4Isc1QJwRfAAhFs3JhvdxA5pSVu4NKqn2cWqPI9rlrwineAWbGyJCvbbL6/c
Nva6rkH8kVSWCdI9zngbFNpHHiK0TUqroWJuXjJw78VnW4Lan1RNXA4JMrSth48/ObWtT1OgHseW
/kxmnwXL0xMOsgZ9ZTLAWdJFzDSP+48WgdE8xY7UUsgINw3Sqed6it9jBErKFd2ks4kC1LnaZJOj
JJrijwki1yy90NBGl814ODTneimP6fKSoxhJgayZItfrb7x5SJlxiGFL/g97sxGgTpQjZcviEhLs
ipyRFAZbZsGWul6lzrg/Aoxuju7pVmAJaMBw4dfazIhSJFE7wRbyZy54BKV64g7F3ziBAKQHrcZp
9ZbPLNc2zWrL4YUCYiWccuZx3HGwAYQLtvh9J+3S5UhX/u+2Ed88ePj5qY7gs1SyiKzRWg69Jv3d
YnxVhLyEQorsDOWAri0UK4rMi6L7347nsz+26seZ//CCBBqo/lcLSOYbTpd9yKKR37tD4DFNqDos
1zt8U5YbxGvfJhOPqNbiXAZYCTCzt48d7Bfmh2cIG+IMPN/MIxNvSUa7GccXD8VOHVsWiMKmgRhf
lvNYwgHLg1F30BXUYd5I0r2OglyP7gCxQ89qzDeyvBZcIxhwAvkoSCskc9srTenEQ8xkNYd6wP3R
fiLlAWf91EGQqNlU/akCFFkNOn8kcFAaqPHkAljsN4W46G5NExSHissPbki6AoFUYJ5WTMVfW0Oe
dnwylhDU36kULxhkb2dOdLiVJi895kOVkXCaLqfr3m/1AgQY1qM97nR5gaoKAc91bAtUUJeHkijw
pKzmYN3ARoLSCB/PadpWLiTaCGKd2aYSXqFk/jY6QmAe0GAgViaGmVjaZNqW6YEaM812bpBVbVC7
dvUpVUbpZEoiFpiRfg8nvtrJgO6c2G3y/0PZv9BLoZNFkQIFDRfZGJ4cOwTa6svZr198J3Fq26lw
16APR+Ob03mRgK45sHJSkNBNU+52Tjac1biEyO1EigSUiGYmVFcfOvVOI7cNnsCX2Be4/nARx9lk
akOtuHzzhcppeD7rvO7n6wOFPaIwLEyIMi152vF64dKjqdAdFuW+k7galQoSYI1+ATKxcxzAVhjQ
L7EQobY7f7+vUTjooJOqqg0LX//wbyFHPOKrWGg9Exi5UIcrhjJJ7AHwoB5eeseT6HtiwmuVurgq
Q8hG2T7lOCQoMIFSV4zE2kN8a3gri7kLueyl6cky/3+V0DpwosdQEVf+DOC00sLfylqQAC//Gt22
KRuf7p6HlvQ5r9OibUzquVShROMLB6LPz6sRpBn0UvgtT6yU2nvuzoHPq84EytiYQ2ROB/WJb61C
rUhJlwAkjkh/hitUx8ghTHByDasOJnPFEpa8k9QCXN4r44lNGMQMM9JEYEV53xk/wVm9u0drYplR
MzHdaykIG55GjuIJJrg562GQWDh8oFKnzlNbvWyn0hmEsLAmFG14xKROcuXRKgk2BSBqm7wJafvY
uDegeY85ubWq5hgfi981sG3pDn8zz7NRimhD1/fXME7N6IKhtvkMCEzs7GH4KfZTmiS4jhHGCIW0
PzWZhUkIBWp55d1817/BOhkN4okSV4Zv2i4ppugLEUSh4gNHEquitkHj6O9Sb2IczsmdYTkDoOvJ
3GhV2PVQyFMPFk06iHlcozzyE7ZedOqRXy3h3oNZGKPMQ+neJxQfMi3MPIGr+Dt63mzxjQSqsTKr
up4Jv8y3nI0PVU/dkPiwO9PTqWj1xp6f65HwTIK6IPigcFZQnBtA/H7GiEWM2FmP73d3fH1/8sXO
98rYyi4Fqoa2VkROTLUt1IHjHQVBbuyaENwrs7pZS3kV9+u+fdrEwpSBZeTYi6y7ibBA+d/Fbfey
dSusXCSfdH99Bg8SLcYhsveO8coIslGr3bbEq42xxlj9QLloqmDmLB/KXcI1skfAaL4FLAm7Pec5
4ILAq+Ofyd/Jp/zvbuELCCHZQJEG2J7VQlLmLjPn5MbPUTRQfUm+QcW+aSKhXUHpO96ZOczPLPd9
77WI5bABlgANs/NRQMY3GgMfsXew67Bz9NvR77u7E4lNoX0FbM3GGM3TiFH7NuWqqCVpXjTonXBR
aBIUu04Gc2JE7Disr4zHzto+w2ii7uk7Wxj4TvvouyBurkz33hAAEtbTCJLv1FaKDXLThjekZjah
4zvj1AqXUM+Rrundouza+eLYexUnYAL1YSwkEAwQgQQjH5+UtVlgdZsaGFDvkeBfO8CUquAt66WY
WsVQkCxdkcGEMOZxlJxjwxsr1HyGEtXeenxD/84lA+BZUlhJlObe5CxKmBbjFGvxvivpjFeJpVpa
mlRzCOPKFcR+QHP0p7bdWU02eCyXUEAaeRova8toB70Kqi3tQJE71/pCtiWoJgmivZBeTaPHQPAn
JmhVq0cvqdZGh8uFrtgs37FmQ+YxLTom33RZB+gQp5jzSPPUmkdQEJXihvQCidJELaCN6vzPw2/m
xe5C6ArpM9KBMGeOmDlOq4QC/0r31iYtrh2NUYwgoRc9FgNDTet7n5aTxF1ri0+XjynVebVdOJq/
aS1Dy8db6HGTlTv1KHowNRXpqS6WjFthjAKFDzFMDOKcRkeP19GywGdgjwrU0sN+YLbn3ct5uVrT
4HY+PEenBJOgSF4B1Jmhe5C3hM3nXpgp5wPH5MBjpweHBcactsLc70h+lqfgc080p6kraOloh3jP
6CCTFfvRBfuRO3SUDCXpgf1T3NV82nRkrnwk4XFKn0oYf8nR6+4I6YCn+gdGGA1RMKwsFUEmdX3S
zyM13X8U0DxlLpqr92FbtXvLYH6uqCISV2ATmWUCjJfh0BRK1M93yQ1D4f9wiv8epGybYF5jfHah
PSw+GaXqJ39OucDJPtTtMrf3yXbYMhm4bL5lUR5GnQ0U2MtbJD68C4iv7uRXNk/QIdW9G8rzd7er
LEB6kBiklvZX3wCbFhlmybJZZjFaTRQz/8Corl7WATcpQtVnaVIiKZUT3jL8ZmIreV7dl+T2HqUb
BJmA6GqcHKR9PZ5cF/wJQ6cETFgHn2lmx3wKpRQhmmUGzmrqLP6h/+JH/2qJ7FH3HnQVfvD2CI0l
IAFFNArUq5aDxBjdxmN+sxXd9oZbAAzfcAjkAwoRQiDlLenulYnVvmlj5FSvrnzAhxKWtYPrcQL1
yiPvu83bLz/fjlK7ufYfYXilWNWjgKf2IcwQ5C+TYX8Nz+pWLvDzMRa8sQxQ7AZJIyC0FFRxhe2+
RZU/QY2HOQl/CnrT3EmemJPCr7oMiTy9mI1V2coXLtGo9u9cGxfhddmYORFnwrxqOsSgbEehpf0m
PH2If3RPMSYSIG4WTIWE0xIqDdCRzXNCnq+wBKgt+AUK7+mQDkQaLjbLPwozdQvmnJZWDqmf6+E8
TdF/tIwtp59zvAkN2hIbwdDuaPWouwV6R5O+d/bEsYY6RjokZ3rwevbIprniP6UXmpb/a1i84mwu
a3K1S1SmqDrl3IDHXhfmI1LElEsGVZSGFof2e+tT06O128LisvNj2dhMMl1Vd4BLNu/UrrEwNCSp
n6bB73kLNepnFyIlzXFLZc9g5EtB1YjEaVvXhW5bg3KaJqwm3K6GvnnjJFmxdNnieM5aluK8bj2+
UFWBRSpGHfk1lxqTzuJXG2YdZut6+J+mmclpyMEt3VvPcwX1pc7wodIa3U3c3pbEQM4TBFZOmK1G
F3zobIKMZRs8NF39VmSPuPxZ/GcGBb9Cn7ewijc6rksONQsgulFsIzuPYGoG4YGQ7lIrFro4Rs0E
9KLAfs6Z9Tyuu1/VDu9Dgw7f+xHpdRf7CbjTuOmNE8UQsFQi66QPwadU61aaViNCzvm3gQkVeYfM
ANbfqN4niEiY9aXddQMBIUQm4AfEb6LmIGv5TZa2nrq75MWWkJEINqXwDP63gcSU6I+bEi05oU8V
zyPpgzxiCMr1XXiLqvP61zpkHX9qymoLgCYxMXdMSXeW850XwBxBGLeYXdfff21y1/y488iqawOS
T4oVWSzzVjwSW3wC3CPd48BsLzN4hgai3af1RMfSuetI/wA/Ka48qerqsTFqaymGYGMsr1YN3Chl
lNlhZSzXyIrL6zgaBlLO88bSrvCU0KzDiqXT47/7oSoqRYwNiqlMPrHJ+l4VCYB3NKvaCqiLtXUy
Nnl6Y7ZEykpqxvec5/y3j5wFXE6Df2OdztamNGk8jY+Ci/l9gfeEmLs1d2jrFJJst98UMK7T4aqC
MTO4CYXc8MvJ2IHvm/uOmvi1nr/5b/pfDzF2YwGXBa4xYB+I40qQXmvVu2r/HrEMrnCYdkjajdXJ
9KN0ujhBC+b8X1C2NuJfuLqfFYsnzA8Bvn4escMS/4/NYIX25XA/gAdyOiXLuLJbdt97eGnBmkd8
VGNmH/Ftqxg3Gu95tmwLJmTZ9RX3rZz63RtcVgtErAQ/p20h55VPvQawywJAceNzQKucAfknohsL
K8Tv0WondHQgdEMOhqZdvgC6afuwEenVgp3DlUwYJ1/L5+K9znRauJPBvcw3Jnh/dpjt5W4QdI9f
GDE4oXrlpcNm3okyttWyRV3osTHovoNAMjJ6rNWYEtMadGRgdFLDvIM3xC4gB/LnkFgilpLDby4m
DGZ2qC6miC75qsleYELgzMCJQ7/gF4OIFJg9IJMO3NlvG812KkOFL4jZQfqB7xLU2UMfiw+gr8+N
O8kJjTmVtoNk1/m5K/hv71Zy27ndFZsYMo5togQ05vXLXqe7itDKzBKrN8maETNt7xUVG8xe28A6
4tl+LbHH8oGC3woL8FCj+yPUnxjUu7Vf/BN9l6JBAY7ZB0CYZKFy5WzlbEmY9KhsSD9jZbb4uFvm
27onuBm7pyfY0rTQY1EcPWzoe9Xt/k9GUgnD5yddpY2Kz4fo/7ui07TqRzbiK2rAsf8tSt8wjDA1
2qycVBvwRaMa9zyAsVhxaEUCWV2PqY3cdTahss2OpEmRjK6qJXYlx/dnq2mVnQ+2FqKRAWVb4zMs
j+tt8O8s5fHeqI19YNBZLlWCqy5YgKs7jVHKi0OFWLJjPlPc6CycTB7ilyGbJgSp0Y9t/m/Yy9/Y
xz8wgrDfKv3WZquT0dcr1i3fQ1GMTFBflHCjfqMdmQrfmewGvbJZ/hF6HCAT9RhqsQ8lZqaoazsR
o1CQ1FjaNQc7ah6IKlgjwNz7vGLZ/RySH5FkP5zSjol5sQqG6HNTaQnpJLmLtQ1OJOew0CPR3zyD
3AYfl6IjZg/6pXmL+FN6i0ZPFSN+sBMVGwwOumTToolGrHzDxuBoF9+sXI/wVUjjo0Sb4Lkh4A0c
hQZyvE+pIK0VCO4lQeBvQRYeNqmCjraA6bRaHPm3c4APdsz6Twe2D7X6q31vQTUwL3U+p7QZewDm
PfxIQWWmkzmJneUmMn9qfopKfPhRe/gsi+FqlqS5QwxibzLYUxbl86rNC5jjdi1adEivOxqMy+s4
4/J1/ZmuzOmpjE0LpBK9wMVn+shfTh8/iDLU6WMB6huuv0x3JM0fnDI1aF2I1L7kAnZee2WJr+Cz
jg6grZdcClkRDxePCuk8PTzx5gbirhEpIDp7P+ZbTqPRGcVWeAWJ4MiPVBQZbsSMgYOD/ZOC6ReK
FHFGUuki0IaHWJwQPKhnKOaYeLOaOketrSHnNq91hIrOROvLffhBa08PjoT7xyh8qI8cRkWe/UOt
WvcitsHH8OlUYrvs2ReTGKDJeOVS4uHxsWLJbfawDg52+mQEa+3g77TWm+4tlYegkzedDJ/M35vz
kRVqB7rADGba4x3upiHFUDpOt0APSJB/BFl3Vr7hMP5EbdM/5pGMXwRr4dzDY+WOop5WxTF84h89
L3q9D4Yqu5zVMa2IifcLwbOpzsCsI5JI1bx3lT29vc0vhuHGAjGdCbaeI7Hh4LxAs6xV1hJ1H9ZB
YXE+DOz4wKkIQFx9+3DrUvHzgjm3475K5iYq+DxlnMutIG3t4RL/Pni3HXwETPcwQBn8DzWxUqpU
K8p2o5GhtLf251w+qQchaiMsZHld6+CsWRwmqaV0YM349e+LIbsW/zemb8Ox3ClZju14QWGA1/3h
a0IFNnLaCOvTNW8sALWZEr9gGh8kkCU1KvL5imAGj5hB5CgMVzNQW3Nw5Dt99Ur2IlQNOofMrq1/
/Q+eEWQOyLfa2BctgXsWL+P7gDjcA0un/vf6jr/ZRyyKJN6pkyh5GPOTrQ8cqMACDviXDEm27nWf
EvDYW7pOMw/6CRI4RYYZaD2UvZmo5T/f6J14Vqsz8Fy/2rz88/QAAoymulS379HJaTdGql+EAwe8
bzrdEPisWmWrkQ7cEpc74dUfhorr2Z5K064Ym4stobGIBb0o8hGh0Cv2CK+7KUpq38k8vlsvayEl
2yYWleog3N8rcZajv62V3YZqWpggBC/5XAXb+A7UIbrLu5NA/UopkTmHX3eV7LGAm79ChBkfPNhc
kpO1OfVSPl2MGjO45KRQd+G3E3YimMJfGmGr3mEPZIB8Xl64AGwtnW1t4VV1Yc79YVKQne9iEOjU
S9+ag3wwUQlwyzNC886hNbABoL/724mwEund83hA55s3BxZKBe1O3A361spTEFAfAdygvaiwEw0t
0Igj9bzZVkbyQ82cdqN5/t0naMTaSCkOkxv77hdtM9G5qgEX0n9+nX4j5VWKtDPNf1HFtn7knV0Q
fZ/Kxm0pDviNvfK9Y3N0pqdRB+JYHTmZ+q/9iU9eepCtlGsfvRVpwxR4SoAStaxnCPWozax5I8SQ
bI4gGzUua9F3NKPCceBDLTcQk4DiA3OVUBS3ZrCQubQzROrBIJwBAt5S+JYwjGyORlPzsgvg61VB
ris3430WYcfNclqjDBI5y/hz+Rzy9j61XA6IssD2Fxw154Y8W74zv3xSAC90Wu81SDrTHdmGG+fg
9+jSU8TQo4rSQgd682tiq1Ob7BcZ0xAykrLlZFIsOzU/d5tovi9BapWxxniF4A2br1IRRWumpprz
Cob9d9qfYQOjLJZ7VouhO/JSUGv2XZ0fXCM99CA8VZ1rvHWk5pGqEDCjJJfQ6xZvgJidlI8d1DCn
YvdrP6JIiCg57L8Ro6OzypmCy325eca/5P52sC6hXCeqi0PZ2YoPPJKqtBuYgRyICmFgQrE5ia4Z
HGFreHdL6dmJfK62QFVkn+Wg7SfEvUbpbbnWfzPDCXeNvc7VZ0+2sVL64YRShPMXJcFU5LSFc3ra
AY6GVZo5wFkQRHilPbp/lSiHAhXXJLn+iq/cFaHfful5MY2PoGdUXnbmYrQPZ+zVTTsDM3kki5Yp
0qBlw30lxHLu1xajCdqlrW5055GBUXw5akKbtU1wxu8t//gD6Ez6IG76brQUrnOHVREapQhpS/CH
nnDSbmIlJGlCsBsfrY86xGwizZL2OZFinuwji6CxXQCVi1zQsC2Kk7hSXH29t80+61dCtKOVR7rZ
fnC/WshHecLIkpwj94BqYsnef0fNTEAtmB1ZhOJJOGslXkdQYviEIOWu4DZLL6bD++KPxQZxxjok
x1ey4uO6JEqKlrH5tKxB8kveD3jjhgaDhjrEk5bkTWjLnDNUrEBjMND/uaDKqTaGFSMEjTJKOZ5v
0s/OnpUNpx/zTc/K/fazgGwWdl8nW+JjyLS100PIs+FgzQTS+h3DhJ/7jpow8UAIiYKCkdF2lVSJ
bFjtR/QSoRZAi6R0zlykgtXN7V1cvbIhjs8RS5wXkT1iZrb+SRaYE3BUGRtMf0JG2+dGNtJcoxeH
47HAW/lsVMPqBTdPTSIiBkHsDocYiBTATv7aIAb8N2790OcHZz1pD7+b5jOYsB5MtBLwyhw4EWVd
8qgY59TNnrg9Zr1Vc0h1brttnqij7EAcihht70PVQ9yDS1n2C8UuWC72+HU58obsgcPo+ZTj0I88
XxB3iLGO6lqYF9XjIqrTyzSZI5eKTrvA8a2nRrB8+TrYbf63ILL8gFzC28rFH7dDDTeFIeBYm/kO
Iw/528jaXDmV79E177vsNH6qARLzg+2U4lmjmPBEH7hHm8f/RRDZrNWfg7iJC0xbBZdr/V35x13B
emwkmBStDTT5Bmg9B/KHmmvtZbm0m1M5rZwqMosG+AeTSSVXnis5JDCpg3gcT7ls7bLK05zRbCj5
H6fKO0EkHjlgQWZgaI771BlOHjSXYCVbV9+OiIW7J0HXJ/dBNLYfdY8SuPmTsHIZDsQpMqHfB1y8
PGdo1icG2Lg4aTaXWQbCJecAQ2tU5fU89FhmJgCYz7QtTJ6SKW4Nfh4KTF85n4BFsJ6ZSkb9enlC
kA5xC0OYtbqbvX4cSjhXDGyw1ml94bBWskfUBDPYEI4R83ldKV0DoD1oTwy6/DgHbgzyGDYV2YQP
8A/jL/9vrLKc+x8E1W3b57ojDOmkDxfpCevew7WAii6JsO+Dlzhk7/llN247lfMIKW9wJ2x6X2S1
mc9QwYCYwdN9MgV6xcniiMpQcw2p6fHJPtrD3Ef6fGFOS8bolZThwiBLL4u39ITvrmT2AgaifkWg
3KF2MkIr/ZWe5WKP1IIOKp0vrxz43fF2l4xeZGNxKnc/Sp0RnJOf/ojUPQtehrDCKU31MVkQVBB4
OSiaAgpE0EfLgYR1xuCOI0Hw9ZmfYxj4DRVvT+FqmTP4YXOyMMdO3mvRicnkdp7j9IO8803MJeV9
wZiOwHyefMs/gWZD6c9KsIW+nKud5KERNbvl4VE4n+Pr1q2EQLHy5ZvAceU0Mjc3K7cICW6neANj
z1pyUmvs2eRr50Vc35r13SuvtanuOuc0Jb4Jvmmn6E0Bh6YUqf6twkVho+y8/gUurEAHBBRIK8X3
hrqSQgobQEs3EU2sVRVN+/efsrIB1vwNuW4GmS1NfYmTHz9WV+d0OkNgOThKCrB9ZSSYQlG+2KTL
oThXIaWgqOVK54y8BTZRH21XS+PK/qc2nkzwy0RbvgjU0Kwckbxz5vx9qeRENelRMiwOHFRgyDiJ
gxh7k3xvayoUiQ2H0ucCDW2cEfONc4hYzdUhTS/TR4qvW7igGOh6iUvXlWE6ki4zThCX9MQWubzT
w/FcbDL8cZsWHTVhhYYJpX4+tg9zHHqRp3hr71/3RqsSqauinzOfHYuDEgVVo7XAZJDj143mrBMZ
ixjir3TrUOCYdOD9KlGr3KaAVUVrWjigHvIYww01rHb9WgKfbYaW8F3qMWHuTBPeJg8MmhNS0066
4QxWZLGAj3xSqqpNUkDODKQ+nZ3QOKVZBr/QSqyrcP1kxHu51JBCdNqqbmfBvUadULGaja1hdmol
Wopqt7QYNWxTlBR2vt6qW6Gau8kjRwXSYqGKg4H8W4xFv6fscuBIlNVjMt0YrAP1f/KFHl1q65z1
usfxtv6QgtXkID8bOZZ0aLCrg10BeglSLDeKaDfGYBbObsBmotv0yBqa/ycED/KDSB24FMJP1kKX
DQ49X3mT86ktbjMhlokZXqUjSSWovwbgtrDwkzo8ER3Du8g+idsofsMK6ljO/5s8DLlmxVVsv9sO
bdSmwX91crNQIEoFjlt8UjcGG6JW2mbGmYP6g7B2P9LNIrHxe3T9AnawpGLYiK05ocAFJZ2xW/fr
7qjsil1qh+vYRYFZtH7muOPoI6dbrENstHuU/QnwUCIzs/bdOpCLPY1RGmTo2hwln16H/DwHtjQI
7jxL5ZsbrhB1RUdP+JJKM/+CIjeU+m7TEpRpvDVGIOUB8jegf/cWxIMIw0+DNLbl+eEM7FYghdnY
KXLwFPWc/nga4O1vgZX25rBu3e4WFQPd3+lik+1EhQzJRCaJUni5oSYXwK/nw+cLNQvdy40QEjxv
0P0vFCsHk0HeLByE6f8DkAsuc32VXwrHj8UYx/+b/h5BGC9wk7n3QXuZocPQdv/D45naOczRYxbF
ekrfBtJOGCRd3ARL3CeBD5gCsFfnugL9sK2XDDF6F5BwNvOjeWAFR8RgQl/ZaN0qcj8063YesI1S
IBL0IFynuSjqFaZ2++ldW9QNO7P6SsqEbDvBpXL2mcAu/5mIOQJbF2gTahCnpQcfHR46RBZ6rbtJ
7Mu32Ew8cIpkEoZllow+NX2Hdd6Y/NgAMBtW6W0Wls1JGV2Cl/PO5z8EdQSW7ffwuEOG/COz2jId
8o+vnU+HmvlG9CgQv1lhBq8vcYvqmg8tb4VR/XOtS7hEO+Vht5n0h7HXcPyF9v7u2MXmpWf16pAU
U8tdztb90E1y6S/lTOIxzSsqG5oFSd/dSBJ76B0AFMganxPpqwQij0o/EJTPn0bYjrs26yqi0yU0
tEMiQhR0eAeayk3odajvfk1P6eP2blf+vPu3XD8IEzfkiZUK8NRQGsOcvuM9CEaG2/4RAZkdx1EI
rkWJQIkBJR49nasQllo5Rzvuxafp0IXZVcTP4XVQ7ZpArTjjFf5GElIJchJnf7gKmAa9chKtidNn
YE+E5oG6qqfnrh4vhFWvxSGdQNHFRiKLtUdusvjDbcK3nWk+5SB9qOhOZn7IkyUj0hJl7Fyy9MrO
NJQoHgVjkrXgU9BEiBicvA+ftSkYUriQSDPpshFxXR9sMNLqea+WNzPwgq+dCLvlZHIYyV55hTPW
/3pcf7z4oNxVI251SnzeloocTtSh79L06OVE2Om5OUV2xTPqNN38qnWL2GsnT2A27z7XL9eQn8cr
2own+uvs2LjUrUuL/Ey4L44QWKznvRnM08juwrcIiGUrWQQA1S0vza6wfjHyl4CAw1vs3j/Jz0Ti
moy2V9Kcv6oAfkzNXEaSFw0/Zcq28/rkRkZIctnA12qx+uO7GRLmGv1RWZdpb3TpF+qZSM8pAH6u
PgK4rl9cs2qNu3M32CUShKW6u8/WFaYt6kG8o9XiRPh2uahBHFrb7n6fEGxwmTTVEVLBZmFkiHkh
KzAwUDOXFLeBYHf0iXQ8GLm81Q0Gp13W+N9TEULUCKpMJqadSrDNBEjLrl6G1AI5bMcnnSUOR0nK
xfuB6PMudgQ1dMbmnt2XDH1Qd6JTQN4bV3cFAopO70t9s7C7Xsey0+FGUCfLMWyPRpsQIMeN0hl6
mbVxTShsXvljTwfyr++boWXwFs4dgR+cYa373pnrkZjJ9P7WlDNhXHbyN/oBxsRtINiiWuRzyw+p
bLQpMUICeehn63G/I/gSpPtjEKKkuUbvVpxDR/G1YkirWmc4UrZVdiSjVmOf8HZPi8eWptkOlSyx
jt5IKH3e+gk0hqOyJZygdwix35LdoT3/UW0IfW+CzOG4tJvqzMMafkdKvUv3Ki3LdQOa3B0zKvrV
LH6asdr4yZu8EYlVXTf1gGpDo/p7NiscU8tzLWvLVDvpKCgQGcIJCLmp2R0PbQhrSzHevWfGdAEj
a7nOi+sKUrLdEmh3eYawqgnDNCbW4/XxAvhNGoM066hst/DjQjU2l7rZuRYEmujJSZFZZWcDaYKj
EcfsRq0ApCE3Q/wgRz/KP7QbZDxCjD/f+7VaPEdHhkN/OXZ3FNMVsL/v76IqGyfmWBadyzgXRzyz
1YlE0jp0BhwK4xQJlY8osJ/3cLZRSx6xW3Zz+I0VDorMq04VaU8rlNhRLy83upQwUxCuWkrrfl0p
9s/htnncadgFUgiQDRJs/xSuYAolFDmpocAyOb+UMyqP/a74aN/FjVSyflfN3TyeDUGwC4nH5z7D
k0LiL7awKRUAVA9m2z+sR/g7qMJpqHaWmznzznd/V06iDdwW4kFWRKJDGkXPMPbBSvENle6uGBEN
7Kn5VeqeTPkEm0srFovm4kD9yaDOMDV+Nebwu7zOj/5hrkTGwBt2Cm7yvqLyPYvqO0tt/zT/WjOU
EHAetXTUe9GVvhtUfNScksm+M2+IS6kniuE+bDJH2zEm/GDMUO2DKYxS0iWLWuLkDBtDqFXC86GK
6qwF2Vhb7qGwaB/zfiLPgWEnvjtJJ/1KxfGyGY4F5VgJqCPk5SYwrviZ+6w9XCiwPKOHtlodsQCk
kQJ9LoC2CNjferqhLXw3b4NU67/cp98TfpPPNOwio5nSBQg2GouZO325YqWvAqfK0FiryytjKTWk
ev9KAxmWF7MjAcQI3CW4EJFO3kEIZ27JgDbJVEwTQ+nmKAVQlGqQn3gwFTHdH23yjZoWfMvKGU5g
MDsGuvghBsxzuTIFW84avTRHutQBIAP1HDOnGv0FdFf8lKe+FK0Ia45gp7ABXOsKWq7Z0RcPrJ6A
jPiqmtKJ8EYQrcW4SKjL3MtOmgNGhBrYAz+KK/Wx1GB237UHZkrQGPR0TcQlBrxPd0xvIRfB7Teq
UB4G8UqAf6EmthGEhzbKqwMB/8OgHJivOxhdQ1yv9mMDZKVXfKJouIOacL7MZ74xUD6GV05/VUSZ
Rc8L1QY0SKaZ+1IjVctOKjiBZ3sJN9ELJjUye0pScI3LMFJC0acDFmctP5fIg+qi2kPm1JQ/EbC1
eHvUtChcyQCTJvYA1CKKmpSIWXRe0P+TMNH6qDo2YkmyPEAGemEDYKl/GXbp/Qwty1D0sffKweXr
uYwjVoaFlb5CXYouuBjeQXEnI0VFN+91FSV98GTZAv5qKNUpxbGSMMIfcK1UuefVitvrTy0Bcp94
O9h5j4CkgBbng69rrTsaRLs5odGTFr0EuL8rYMRgRCAJ13Wrb1FLZyI+sD4gq6sUFMTPXIrEx0yq
Verd6MUiAICvqQwly4+0fTufL/+JK0lVIV6JzWfeaXFIM9Ywn3RYCAPuOSjaNZxv3hlja496s5Pl
vaA5ui20RjppsIaeuMS5qPw3+bB3r7tjMp3/hoCL38uR4Ch+Rcde5Y3+HTFk2sdjoPQMAeKUcF1f
nCjx55dem1etvZQFGM/At4UgCnnGuxQvc1Y0t3oNdQQHDRGRGE4tsswrWevnk15TyN7A/esMLVPZ
3mU5Jo3jkrXJKcahM7LPor1el0gmUqwoyRG2XUKoA0BkVKA+FghmhNenuqHtSwqLYBvkj/zdNMUG
1V5AUoZm/eiWFYJ+vClML/gWe99hUJuod3bLY9gqkwD5Tgd+Qs/1yjNinMVQkFC/gnNJuQuI6olq
kWGtYzrmvL9UrluevACoYKZzzMNIktjjsPm9IvhOLWPLXf6JaaaL37MwnmUvjY9uPfOlrT/uj54c
XTpJG2Q9/CSihBy11anhWso75BweS5Eos8D8CVw6utmxsj2aeh6Jdra/QMhnohJiUAsjucpQeItM
aP5aWscZUgZQZ0uHXsL3x1uHs1J/q7zhKxoznqtvM9zX4Slx09uMznK+dy5vrGXUOkhkKcXGwSu/
gS14uEgsfO8z3/KpBeV8OL1u0MPf4vxmPSYJ5zLqJ5U2rTCk6dW5bOdRIBdt1pIppfgdAIATTvzC
D+P5Xv8w3rO+jjA07JNCC036s31IVABUnzw917E5YPItUYzQXQ/wD8q5ktwyu7xgHtPXf0adhZk5
c+FBbEvY/GtRu7/ebq2wC1zn67AJFEYTpbpsB62BdnxKBYRMWN/KmRLjqeJfBrTokPOJhgJib4QH
FWqDRlmBp1Ih9cJBENxMuHyoEGX+w/MQdDxRC/4IZomh2OaDMnIpr34NFEyQS1Ufwq14dyuypxwJ
Cl0gOJHfvZqqQ0gRkywMxNFyXtHSFCW4PvPZQU3Fekb/XO/LaIyeiGWnwiAJAVFNqoz8o96jHwhw
iQhorQGfvyrU+HDF9RYpdW7X4qkBee1/7JeWPskDctwv8yke+h6yxkzAcHjiBPJGmWUHyjGls3RX
MrRjz/X06Osui0nXO5IT+0uuwKxK/BbWFEwbC/HYG7SGXZyRzvmS3oXvydKK3dvINaHvsLDSHGxQ
bSGJTtvuo/XvqItj7ghlZbZdMn080dCrXOXvXLs6BuPSELZFiagqERWfjY81qnPNR/xqUg45qSjJ
il2Z2d8lMS5re4JcBoxUxI93vweJFVBpVTa/gYczEZ24yWOZrmJKngXWIPYDaNxYfDyRGczYVvcm
+jsWT96zfzQk5jMOnUC10jhMH/iwW8aGuw7FnZSYhoSrBuY33WMVXWFhSqdZuHDOHceM7pChU2dQ
JFMmEFLe/HI4XS2FHs10jhWf3taGKk48IGEEhAQEdJAx3+B0MxXjzKPCxNG+KZy3JduVNOk2u4Bb
tA9o8GTxFJbVL39mwqm07J5sSHdt/yeiys5AFQEgKmiLN0lipk/MGMAzf/4zg3x71Rmyuege0bKN
mJ63SNJUxQHCMCkIFHesbh4LcM2dYj2OHi0rSFXz/0/73unHuGwLSSmnsu6/IdBwsig4yO3eDEq4
XjGEvKnupNKUQ6IJSFN0TKJ1rduK1DcjR+bweYXwp+Aol8GUwVND6Uz9Ucj8IsnK3N0K/qTKxCV5
VXTJAE94aLnciTyKS7tvpwr9N/vKjF0BMk/Y9CXbkraUlnhacwqRgTxoIcVXM3mjBXcjbTLTUxlT
olePRTNf5itPMuBqqLDSmgqgcupASsVyK43kAz/3EOfgDbeQmOfPuZSC1q2QOuGf1csUzePaeM0R
rQBACwhMjsHsZeyq3W5JaUanCDWUrOVKY4IDbmbEPbda/wTJXu7L2vCG5RddofhwFqa2QB9cLf2Y
NF2WpAj8Lr9nITOujzni4rdHNiDmL9BOSgKplH5heVeo52Au9vUMUcXoAlK0E0IrxBhznWU36bpL
OvAZepEoA4LNHbeQkit1B573/ftPr74n+MYViqefGb9+oKTv+muN+XvZVx8pMWVZM4+7sunfHeit
fpm62W7nkyh3SjuhmeZf0aNy8y7jYHp89J+XhSOVV9kPu1xOLca+qdoUiUIMVlIcn9lx5ZmVXoNA
pXYqNcvI+ySzRA68ev/kAeCU9a1SbMbL+Cc772TCtHj/mAKF5t/s5MhiNsd2L/pIRz/bquDq8I8X
UmqB3+wQC2g1l0Wy4iEyGbka1vu+xmkeQW7xLj5MU3kjGfztZG3dnmy7odXe10SNu+17minPQB8s
fWiuLqqYC7zGTeqhrOK/AEeRJXh4nshTrETTNxd1eFVn/t5iZwJ8WCa6zFQc2CMHCwVdA2n+u1AP
5IDEzS7vTxMgS+Md/mc9tcuyQUzyvRUx/XcnQ+Hy7MdnFIlRPeORZ0kmoy2ZlGNpkWST+OhcSGhd
eIR8ZVs/kqiZ/x90zOC4cNLVIU7qUwJ0Hpy+fPS3EO5pbVf7d1e5Gf0ZXIF/YHvevV83fH/pym3Y
y9ZXWdpUk8gzRDQ0Ow7HGyw3sC9JswATWTXy3nbYnTZ8ed11zk9GbqVuxotQbqugfGDJeo/0kDba
IHo/wYB8zssvkWq4vy0qWkOMQzDvnw1pnlfyAr53SBrBQVkW2SZEWMasURGtKgFTJJ4dbqmZiNnr
egnzRP2Wfw6p8TR0QJ5NME5nNlTtxL0Ng7GheGCiisAEyCmXgeCDqyPTUnzicaGw1y0h6nObUQiE
Fx1/9beRRL2m7K6D+KvHm1zzPZW1X3A8RAHbeJk02hoD/DQSs0H+qn9b0PGu+tmZiL/Ic0iODTXa
IHHJoMu3aae7wT1osbe88F3KT4TwuUBCQ3MplwFyoreLavc4Qaqj8wdMVQEO2pzjlNjRWpOOpaha
japTATydcWMGrfeLZag8BGJgAkQO/UHpuruyQap+hPBMkIPkLtjdE5ob3yP1NOdfsTDx968xHvfR
THuaSXE8W/5NAen+q+Hh7fdDjoIBF/nZMpXRvdI97X8pINQ0NZsZnqUsqf+YuBOt0G7mhrVZx7sD
SDkMJTHJjsQCTWt86gI/VUZabnYihMoqTIGZz4WRIrfmZ5Qcz4UEzNBCloAnHcG6iMJOmuD24Fmz
7+RO8Av35TRcAyUvvdrsF10+ymeV+39KV0Wv0EC2/ZVc67tMZprK5k86gMaISh/KFnqQKZi4vSfg
cc+aLWxvQPiziRxYIbo3Skqj2wH7O1mWGnX4FNci2vNMZoHaNB14DBPSpQa+tz1XRIEOC2QrZ3ce
4NChqUeOmQaGf2W24W3u3AGWbis8Tw+Ln2UYzZ2SB/3xp4Tz5oI5BIvkjgplS6ts2bfgFqsfxTUs
NdFHsfgZmufKF0Jgp2S/556gylMd9joW1rgsW+sBglni9NEWRPT0NAIvTEtGq1aS5kXCnbcWfUX7
vOsHySfwp07atUwcm+vOF4SVF/OyYlZowUc06NaqfKkUuG9mWc9/HRi3gzpzF9f1OwopGU6q956y
ZvCfGf+sTi9Ub3dxmQhMYKsgfU+vWqU2Ougn5B/nP2+8cg655hCXSYLToDhRWNu7oSTY4Yuh0zxF
H636Lr9w0ZLb9q2uuyYGZGeJ/JjRC4EXD574UduyUj/bk4GC4LJXkhsM0v+p1QLLHTIa1yk7RsvO
KPRe1FTTyU2sOXXW7Hk/cUc26P6mEP9WJ3ewDRaDUJSRVdw21QzlCd1tnW6ragL7ewLsR4iwexrY
FtY9ufhYhO5SDHcuyW6Abmu+M5Iu+jqg8sqRtrcpncJ4wPc8/l+EMTGywC71RG2RuEcQeKj14siB
yepUWFEtOs+irSTNhrPSy+xBWTZCviFMemmp0nJJhpGHGi3KxGBT7relnMctu6P9nyr+/22AqPq6
9oekDVob4CxhB5peFioXrVsiOoIJ8SdYQfkXePsKuZoRoxG0NZ7+Ly51rb+cBekTodeNF1TH/bi5
Hyi0H+w+guFjF84weeBMm42DLmeigZG+ztJTrLWukqL9T1QnhmhnvuwBvZ/PoA0Bhb8MX9uKrfLr
7k9n4XF77VflcgK3U68Rvy6e6ygSnupLozA9564ZIFxweXNH/DnxRI7G9urxE9Eoj8JreMICBDlc
nGzhJHS2jGRH5uQPAtuIBQaGypH2/CWZCIVXBw6WKJzI23pysesBxCYnmcwkKk1QnleyzeCYHylT
5+1z32+l/94mKCUX0Z9GLfcbqPDBb4Hcy2Nu4inHgADWcsIC0XDpXVIJahIHmjzFIYDcF9q0zOb8
bPXhe8L96CuKSBYoG2Zb6l0T9TLJf+geMdknhJaUyMguVpn0ktHT56YdiotVNpKkUfoeHcMpeTjP
qyDTRPe3o8d9n//BR6HgV2SnMuteT355lc7aLRZy2UJ8NT+5NtlbF6JZvADi7oT0vvjQWaN0q6AW
cahJa25mB414rZBYyOzRotrM7BCO0bmCI48wrkziIQcO8+DUO8Kd99KAAd/6fVoTGCA+lnK78DH7
NQrI0MbLS3erHx6keJxQ/wESnTxFp/tjzVbIq3XGQx46KKjIm0lYTOeoVmlBHZABww0TLGgCkpTy
KQp4q2iQLYvA3/qPbTRTt43CXWjIBGSEdUcsD0BHuD01kingWZCwYn7X9IomQtRdoyU1Cn0QBgbP
9hxwIxGhVB6vKKShiaESOCUDM9PeGXXaihJRq0lwrnh2ZLT6BocRV5aQIVLzMycbWJUarG+vVAu7
EjjwrNAZaqFosUM4NKRKiMRg1zYGBXEor1yIr4Pb7/Q8Bt0DsaqwYxunP/At/h3RB6qEZHBMvvNY
uBStay7tImS8w3UYD6diBxJW3KKSF3iVVB/ckF58zOSNXhkxVNpVXoDcLEpZ9PHAsyJk3vHdZHfy
McYPe/dQlgiL4KLOC05j1HOmBA+/fgNxClPmlcCzk5Ma8zf/AD1LacxEB1eVjFkzZHeU7u8m1435
HsqRVaL4KVXztgr5ThxLbRtjckjRLmwPoRMHuYuoM7sZ4ucJ3q167KgAfK9niMa4YrA2hySGxvhR
+AfnsT1F3JQJacHwqAtwmLdM/ImSq3YyJ1/1G8yWNx7I0UjNL3Ldhp8RtdnUMBdXGOr52L4sHcm7
HC9zuEq8RnoEo1VhWt5/wEhvLV+rq8kbJXYmWXRi6/P7JGmzLv7uwRY0rJsTiFu/HkiTwtiYjYsI
UheCUVnh8CzhMUf4sJBvllU4/hqYfZfXixGEFGsBF7k3ebBcWtkYb1lS1c00/b22wnYB0c+jShSC
vd7+aHSLKFHZ38ZnnZ2hnRfvV29vRc9xHKcIY04d+1ha6rU0yg2+EO1ETYwerZILNPckNNpocK2x
bnAl5THCtiHEkD8Y5DGgskEAUoOmzqcQhxe4+8jYpwneNur6zxrTYtWGJF8JwWkicMlB7oGtIWrC
xcxfOVDD0qlGyYJxQxe7pkLynlOt76U54nA7UBSgxTWFiVPbuNZ4W8ABkXMTq1/s566na6fgkIeb
HuODwmyOjARCEgNPrOQeEqPLSIf38mWGqcPtq7rhLtU4Bg1nV1HC40kcUqu7nSCsrREuWHwS3ad3
D4yuRf6RBnR9IIk/KhczCxup7qB1LpwoFmMxqyAGYvFX47Xn/wwP+pdb6te1/1Z61APguTxPIaE2
sRKawWbbcTNZuJtXK9gUF1LjCPpPmym4W8bdJ/7mvi+9eqwA/h0zwk/ZtEhj9yXaFsYZUrqHPRRG
X2/ZdckAvPOiFpcMB7xVmIy0XCID4NopbFxEy+UNaeaGYa+2at0P8TkW3PrQlfFwSlT75tjhiEib
lK9XZkYiKQ9VAYIMr3bq6wNmK6TzYzfop44nEcWSsl4GYx2VmM8kBaOTf5ftQPleXVaXVLPgXSmm
L1wtkT26PkRlhVC+ZuYBo6QPCtOpFu08AeJoUtQJGuQcKIYqgy/zkBMh5fbSgKvisqNrj3ApWxvI
M32VaQ1eUGhO72CvIg6FFTCz4zkgHvQi9Ks0KaSwtVbjPWJhVO9T1YmDHv6EnEO9OuqnFQkmip/b
k4/Xqr5VekdFmYtKnYWLbiqiRlBSH9gsYtTCVNjaf95+8T5ATXtJlh9ey+sM1XNbI4GsFYJDxu4O
CV8+H4lBx58Icad7gYNlUFrk5K3nnEYdh026691n396ZN/cFwaKXZSpTaOFUif2n7a6C7ePmsEqT
J4qkm3dToCDuk2Py4KtsLI7OPzhW3HgGcyosPIAdrzNH5FsZDNYrrcJ3VReu88LZLcJJmi3Q4LW/
PdnEsmarmNBYOn20qESOgRj04MThNvQqhCPgayEdEX5XvgCvylP0K4ejpSlx/PYBc3fusvYMpgtg
fQXc2L+BTIcSOKTjuqFFMssJZayyILnoknLniVO0JLOQhK22+h7G83/vo7fbUviUgZ9S8sj+G7CJ
DlLL/o6SQc/ux53oZJz9zj+EgmO+HqV51pWXTGNq9hBDBnF0R/0jXxgPE6fLSPByIe2JyoUbZzsC
q6U3B2eKav6If5Sxr4Zpq4g01DPVFfF1VnudcVn4cEPkjdyZVRvbKRhAfpgyfsyQuXEK9AuOaFlI
HVfV6buvhMt16umhbD3UcBU3Ol4SanPvTapyGIZ3IzbWIhGRf6P/liPHIFhtYPIYVtiFwa0Dmk/b
xnHCIfkeaCaTwR5ML6XtxhccuvzC+Ho0tEbuSmBH8hkuui78DwwiYmu++32DAwTkrW+FAE9Xdocm
mwon8nyIlhTeVQyszuytfHNt9LBorlmHwPabc7jAmfiTgLQDahELtd8TwGbXLTFIYfvwukWOOqnD
v/RnkT6Ho5eMuZYVz2eNfH6TTegUzWCmehJ9+OBDafTyvP1EH7gFbxwTcShrHkbIA6CocVcmn8Ov
nVU90hEFMi6k1xXvejDQmYGWOsjuZaSDqEtZmNF/6dCIDAgdWgol+GDaZrrmIZnwijruCODecssp
OFEAWXFHNSxih1g2P4VuvLQ5HCLa6Sopfhmsg9OaY42MOs1I8obnJyJcWfBfqMkfs1zI0cZrhdVa
hmYGMvyCwL4c+l6+Ma1i89KHr5ndOje4wj9kWvdlO3gDKIXh0+LY9TN4XPbMxuBI56BkHfby5Vmq
PD38F5wkeSTPxb+jkM69hWd/QfBvpx+T7k5n3IEQlmaRh3WifBvCPTik0DQgUuT6OIhrJeN1lH/E
psqf1s94eTXIId7NzHjWS8BMS5bC4hIWUa2cBFRRRBiorGCXevm3mR/BM99BnXC/SsJjSFZIH+Qk
HmcTZXQ1/UkOU1WTbdiU/R1FE5vLF0eDbLvcGVXCkvGADVl4T4ize37WQfTuEk88bTyGt3IlX6kR
8mmf+86lBWuonEtSlzvPyuXE+i7GjoQHbHHFZ2f7rLwjs5lmsAOWib4ySIHx6Rtf5/qZm8p1SCCv
ZVr/2RQsYBmkSc8Q5ZDe5Dh54FgrWjgNMTjXg+TmZ/32tU76vnif0U72EvbIYV7PI4/4Uu1udD3A
bDYO6MHe5iEYaX51XomsSwLzOCAYt7sZMWxac31tsKdJoXSq0G1YrUDtXW+fLN6cDLrNZS3b69BL
Xgt45p9O6U7qS+c3Ww5BTzcZx6+Ts1Wep3J0FO1igUqG7BHIJTBnJ/oSng4meuqt+orOO0lWnUEo
U/YV+3KNtFJXEpf5L32BDa4uJ/I0wGtAalrd/lI2R1f+g5Ih9RL/zIj2h3Kym4xUIXg0sBwta/Af
NYdzantrzwqggGO4Foe0nMKaZs4j0XiNn2E9iwE0Enr5CloWPv2pln53FBVhgYtU7mv8L1gMv1Qp
d2FrciWY9xWI7xYnVc7g4G00q4CVdxLUnoLVa4O/ZhzaIz7ViR2zyQrmllZMvYUIHMXZgNmbONox
U7pAmAxo3bmdopmChWEdwVZu6+FhF2fYQ7qqsQGSRTUhugmK5odjpQs/4qtnnajm4d1PQBKFqIM3
h8GXKpdgfWySPL3zOF37CIFGjppI3bKRGdYijM5x4SRTkQI2RFdTyKjn6QPs6nBWTzfAP6M2qC+i
260cyUtWiGPyHFOoU+6OvRAsRjijckFe1SZHXI4ks58R5lDiQ7kAR1pnStjrzg5e9hYSeJfm8fjX
1MuIbyfT1Bfiu74ZhgdqlDDPDWOAhs1DAufp+lXfDhO5lImw4a8HAniC9wVjMouDecXEsNxPmj7Z
cItOPpdJklpMcL6WBAy3PgpFiqkYQb1rJLl9poVDLwm3yHhMCyOfGWJHEylflcF+ZQ1TAdpBAFmG
lGQZsjbk4LOoJFGiBO+0eYAx2hzufZhM+ZLKNzFbKqlYdNcFBz9eLSuRbWu/LDQ1LGfzu67fECTK
x4v1/dQE2fuyU54xJ290zFABX/E6+QERQVY/5dUJLYbhzSYyMrCesA/7BrM9k/H5HXZj9BruLcbc
3xR1gOnYDV5tZgszpDzkO61MwoD6XPM6wqU/5iakiNsoGRgOs/w/YtBr1ApycJapB6J+A535Nl0d
PooO/gKhgIriz/YfJrR7iFHf1+FFRZkC9Mi0W5SV/9WAFKvu6yeQd2mouHYQwH7m+ix5eBZbrSWA
/HYIape9fzNX+AVW+TFdXVXKrqlqAdGGG4je0VVaO57m+7yP3+UTio70LOleZglG1XdN6jqrYa4W
GJYbKry6CaJNiLSdfWyoDO1wTAV1Ascav8n7Otn5VOMrGZ3Qh2z/1CSajZBnsQwgLCnaJvxWB+kn
5yNdDM4SSGHyuz15FlynaEeeYX6sMcAY6/oCAAe/g/e+VgG1+0PM1DraXKku7IkWFvMQmOVzeQvk
GrM0YA2jJKF81besbtNvvFmjZazWfOl/esh5EfQT4jt62CdjDEunBW01gDAae2slPWT3VhcPLiYp
oQ+88roiMCVM+Q7+0LjUH3CAmimz/WcPaB7EwHwZBvA5cixddRUBnttFMdIsCF641ao0Hp/Sj4Kc
5709jhq23AUAhKSffgZw9GAqjd3IDAWdWpFh4pQX/NMPeUm1Y5a4GcxzJN5pbnVdsIVFeM1O6g2O
jfFMmcI0xFKVfgZSiDbK5fgnj2O4ofrUMZTR768Oh3Vvka1kUooywpeH+pc8Djna57TujkSGqW+O
xAie0SomMR1p3mc85aTDImb8B/ecZAgWKpwTuOqv4LTmEBATF1Prv7a/Sf7ZT2ImoGeqeKeKMI/F
puoDk7BNjPtr4EEGALeDeQPVQJ9gujG0y5BO/J0PcmKukwm0FDS6IA7iahmhZ9e9WQK9o+aif/7I
l7VlQtx25yaOXz1Ila3/cwUc9IwDudXKwT42xnM6gBi1kz8dSV3Kv3esEXjqGQQs7GyRt4tJPRfn
dSSJ2t4zR5+8IccLrzi/q5mdBxHIA+pdgeiSTc/kViCGYm+7flSdtIHizB3NV47lzyG2Vn0xJGoO
5r1gbd7PqF0uE6+nv9HmC1a5/1Ootsi0kRJsXkrxQWlp3CGDs/Xq33fcYPv+QUyj5Crrc16fVwUB
RyVIhWel9VkwUZeX602EZMnxFAgVMZzED50EubyQ91q9c2iIFcb62F0wvM14qAkp79KUIfAJ7sqg
MQICDpdtm0iTLKtEQNwEhIFO8m3F4uIRdo0HhYV/vbOoMWL6r7xWBt3kqKpz98fIoGL/mC+C15D/
3tEJngOUPEjl80SwtnxnTVGKqeUqukTQJtH3629PE0sIYER03H5xskSynuibmOIZsbhSJDcGsvKD
gNIKALm1CygwryPssglJAYKVS2GNWYEHWCzQfISIPiSvaJNsEXEyMKq2NBYS17DZ0nDPyqOKderw
1y67xCUaGgSnBk9YqBSJmFOMlljbV53FRTUtvoQbyO74BDQiBnn9trHk4kmIXNXqEMdIgJBjpevG
cJbitMv0X6aYwpUK1A3V/UP8I6eYh9p3OsTXkH3OXqWvB2/ftboV0foKsVEWvnnsoqLXyE4OD16E
K+V2vYr8Zr3rIF3m++iKiabcUZEgfA8HgRaE1fPo4wmDDalZ25lssgFQmRtmJMJj8lfcDDfLQyxF
qo5CoK9lA9RoIEP3MD6iQR2HufxHcjjlhztHKHdE2uIWL4qW05ZisEUY6uQnffbtujQwQogZUzX7
qZZGCrRRx/Nze3dYqA3ssApbXixsYr5+0ajS1QhvZ+NxigwgTcoAFUKkZyh5jtpJe5a3j/RWvh5L
38UZJB29EIm5kDbIrsnbVKXwCVH993DhULlkY2/wW/ZpF92GaZLp11APpIRwaVHeWB5aKoarwxo3
osol9jOWP4PyRIU1jzP5xMDL+P183qNSJzHyPNqfA8lMUqjrDBikTpkkUr9DgBHCwU/0QMAIaLYU
kQAbzOqR7XRA49H5OTkyyaTDH5KgBgKKXdbwejsJFJGn0n/QjZfO/bBV2cmgusEMbWP8Rtt4SWXu
AK3bGwLGPQ/+oLMt5O1QKyBXG821Fpv1UIOk/+89pBbf31RgT0j7WM3vM6lwVk0VWE47yPfKvD5J
S98wPKVEqZ58NdY8p/faxOyiFhPCdnJkMxF4MUiQ71/PpATbXoCZN0AdOwal1ETycnUPKY2nSIj5
toNKw3Xuo4XVOExOY341JWT7AgxxEMVcLrwVhzu2rx6MN7QaTRp0aGzKz5orl/Or8fYf48VgQjQW
cRtAar9/XRmdj8LXWQoRBRLyU679UaFEihdMRIhTfboUIv1zZgtqtBq7cKx1KFeRO+ZpO1RGJfTP
bot00TWxOJ3BA+0m2ANCTOYhCKxju/Gpy1SZHgocVNYa6TpdjWbmAf8RoQdvc+yBk8EVbjRQPNlM
slbbgPE6+Y7SZXZwuK5wu5qGE6KVg7kVmrl6zpA1gCZ3V8i16qeZr4QKA5dmXvGOHhdUVYbyvmTk
XT32bU2Ycx841LzutNUetIYb8xkp6lwkA9+CyfSBzqYCXGC9NzvEgJRQzZCF+moj++mftc8NXED+
WSSyQNCTgXzWvlma1DJTd0hlvpRvAu4H6sQd9jiO1MGBrqHTDOyZgDjqE7J6Du/Z85UiiKacjDD/
jQkUEgUyM/ze07vGfNdcLQPzTP/f2LQkkdex6FMQaPUPneRMxR69F4xnFzE7kC9wCzO9rE+otk2d
9p5KQ077Qde2hHOmEfV03sQPqKbenK5LfO1xm3itzm5odTvY+zE8tKoXOa5g12yx9wG6+tFXnPk4
UGNPSuONroZRsBbIr9vYCsQIOZ9UbvVTUmPsPs13JYxpCZwKciUpeRq8NPYr3rFHdq62Sr+TrbfP
r4dEHIc7ycIpruPzy2+uN++z3H/K99Tz5kHAGWg5PgyNGob/BF2pf9lNXpNYB2lPeZzxtSaDLjju
cCRrA1FX92VZfo65zvK7RXDQgd99aQRsiFelaOdtcj5VkkjVTWh2IAhL3qip6l1Q/7NuXGxjWjpH
fD9lzrbU1mwJwCrCI5sbjjh7tZzXvE0UAt64nT9dwAZAe5t+uA7oBDuPu6YEVVi0bcziMb57m3yv
i6F3DuEKXTnFSNKwPUJRVH1aFWrfnfdDGJdkvhhOOkgdcwSt3Ois9IokSoO5NKkTC+AcGSoQzFwl
9k9WGHQ40Y6jg8fVb+Acs8afbvNKsj61Sc4Cbjcky3oEN69MbBEjnESYnfUpRkZn99hcFty6AaW8
dDib8Duz3ImQdoHejnKUZBUpj42GZ8J10PNtDFwrHR3xpqvZ6bYgu7F4QjXbRuL9gt6euA9TL6ef
ixhTIlN2XpV7D1ucLJFWma8o4ApIqq/9YgsgXH3HvfX0Ylyu7YFGDE4sJUrDPbhR+Gi4vBXNo5h2
71i+EDpwKrWu6m/ajDAyYS12BYidfQs4asBQ6sr+xTj2H+qSJPhZE9E7sBfk8XhgkmrEn4UOU5xk
deAAwnEKnUgfzpPW4gabUPXlTtAY+NIaWVD/G7aoadG0tQrE3Sj0sSrOfdZ1XoCGH6pvGNzrA7/2
1yLric5w3uOUw2wGlJ1vu1BEaRS9FA/5k+SK/qtNW43Hsf1bHBphc4OCZ/+ZoJV2sCO1c5ax3Kj9
uA0d8hcjqSAWldmxv2OptyEEuRouvpUN61ifiQ5lSFRFeUaOLs2Z5R0uD2NLhrmMfn0MIusBCbK4
LCh1DC8TyGd6JuewEznPxfQPOmiWU1wio5WfF/z1Ci7ieA3WWjPCNLv2soWJguePztObB6QC9A31
Rji94yuDAKYVbK0+PqVfWvkiCTYirF42yN4FELLumi7RrazQA+ONB02jKAUPFiDeHPgdQRD3rqoQ
rqSXe2yiRiEaXYFZ97AerUocEyP6OdM3NfG9j19QiKjrozCGiT8vt2pwJMUtAuiR3zy8gq0VIHSN
AqSUi0TIZDKt9AG1QjlfLyE4hxqEnazbdgZVpc6jjD7fYjjb6gyK8GV+1XRlajAiVqMCme1WAaKX
KOSGXjA2pYtgG855W7zvKGD1FKX/zwwU1K0iYpfme/bH07IgU7qSjK18leytm56ztqCPVvA+fHS6
JVkkX8yXxNRN+5ACzqria09jFp0BLNQIPOQ37ZbOP1BYKTMleFDDuZFw5k98SN64ZZdSWQwb63dg
3RwEApN3yqYulbJ3mrd8/1D8+4rleE89J9FUD2r0oBAggCsTt5DgtSIcXLy+StnwnInVsmFt/KNw
COAge69tP0DcrxF7X2o0xSMoL48zLPsGTOYA8yBwwpTObV4GEDz414ZlHPvvHKDnwji4J0D3AicQ
VUOq9N/xsJwvJZ4VvyvkmP6/35FzV62se6GFDEdp0Es9LkQZki3KRm6HKgLd9x43Pt8bFrjspWu+
84PkhOgeaPPwG6JCLUb4vTJUSgSTjR7cnfbteEVeeYFqB3EihPnJ3nMR3VMkDnwD2r5rDZlaNfL/
psO0uxBVMgS74Sk9Klh3zWaSjoVGbv+qsXf8MEmSpU011Stp/dE82wS5wRoN9/Ve7XaYBJrRZbEp
ihAG1VFeU0qe1hQbomWcD8N5ArawgMhcrhsOcKG09O/iHqs3ErBa08MU5XQG9CjY1XND0e7bG2rJ
iKWP9EWgzUS+KXlbfdTvcNBHAe6n3e8TCdi8uexC6dISUHisZDY23qFT4+m2ekg26t5GWNKouQeI
qZp4qSMeI5I+k1kzvNYiqQrqnj725W7T+ukcKl1eLgcw0CTGubS+MKc9suYDpFq6bLAxzfQlm/g+
mvr9JA+f1ml+17pewME36LLpvhKi9zSSHypgZg1zv+jZ3B22t+nurPsQYdR9GUMGz9WZX/CrpmbD
yTh8LOlrcXLyJm+7Pm8q89GXYW7w9FEstFfyzvqEYzALSQZN/JAtCogAliYfk/TA2Uo5ToSMFGGn
IE46r0lJYevx/mKRUjppYajuy04YYH5avGQcUyJyr/koMFl0HyIOhK+qVuN/T5WSJmD0WrWRt3pT
chmJA0uwcYfglnqHIutOT1k9VNsuNhdeSk93QsAIVvu5pWdKS5qRe1ZoxTQktLLxiBj+noN+JgLt
pnJ03kMR6uQmMxrnxnlwoqmjn+EEAx5WmW+X+KaGhlwN+HdxP9OVQHVFqmC2U/rKe+bIdZ/eTzy6
OAwCN197am+pJxfaqbxLmpdRBfggQbbk3YdG7FkTyjAz1hkGLwri2nA/Gbxw0YIN+2TMIrdcQhXP
m4X7beb/8pT6Iiwygo7nRr1M1lrJaZVEGfBXyAkOQr8oFwamWf4EZq+cnvrCTqQvHEZxGzLTAHzn
/OLQLnysQGEoGo7LjQSMMUwBXas9uGqfP6WZk7DwD+reNUuvazM5eFGxlQT2fCfocGKyUkFD3VFe
gjgELQxQ5qSHwp0zAMdtg5nu+bL4sht6Ppm5GphCE2vXFM0q2IrRWkb7MGM4Dr1VACVHLnzFqppK
Hp74SUFne5DEtiGJuU1SKcTjbHNczuJABMKzhjXlrdHMQwAFL4Ck19hxpOOQmqHE32A6eJfQ0yQG
RmV3jgL5LEa9ya3tEeVEnnkCwJc6rBFjFoCIzHIpoRHY/DOZC2RfB+ANFfPaiGs5OCE8iq3toN5S
7lXTz/FRcYMIqt/q8I9Sny5yx+oS2VENEQPx7MXoIaAKeSkg5Qp8b9Qwuz5GJC+lVE2zmaz6dgYB
jFuBmD5aSMAvv3tx1wQ7TJr+zwN7gZvePuS1JajlackQJqw4oTCJWcd8GW1KRgV7T3tDCRwjMGGE
zi3d8MX297Bh+94H1F66zPeWWv7jJwORQ3HZcQYoL9ZS2nHfcm8nQb7KhaggOL3jIeBdvE0OmRhr
J5TYzi63QOzqcfvmnGtCx3kXLNP46IoAAmwhyXQNxccf4YHUBwHvlpm2pQkAwl6frmeJAIHm7Nph
RGISgvo6Ypupkks0djS2mC1Y0Kwg+FpAeiwgBKXeXp5hw7/YuVWIyJNby5cYqONxcVTMvHN4VezQ
qKxLCf85+IbWMVcfX7dY7OgytYq8SDzNh1S1Ty+tpv2geDEqV/IuKlg5F+4UMQ5XIdfk0u5NsJ3L
hx+hQl6upcLhoBekKDbiKebYYjWVmwr5I1YHCyEis4mopNJ/6c3yD9qKFpnoc5TvGm5SddnoMqoi
MmViLMhNldzZreUPXbFiGJwUEx8IlOgT4N7clwaxpu6JSZ0IUm25jHbNm/9Y6TxzfqYASzlMcU92
c4kzvPMX41QRey+GJHeycXMyM24R1Ch+ybnHJfnKnWY1IELgSkT1VlUeNnJQWAJjlFcXvs4Ua4aD
KfFWiWI0VlvtV5QlWjFaZml5yarOiAqByLG/lwugpEBpimHIZ2ScvRjz3BGxYzTSmnhSGFoTW+F+
ATx+w5j7GbPoCj7ThuuOW21cb3HIFmh6hnwbArT7LRg5DFksW7jS8cvMWCPaKq46Ufes+EVdAE4/
uL7b1ag58zPw3O70KNhKBkoaRi8cYMBy/uMh/n8ukfjgH2rUJlpwIol6pQForNyLH38Cc0ug0PMU
xmbfjQSjaLfVs5yJmiGQt2+4zz7FAyhYpFYJYM6bMd2wxEocqCaPHvoCrA8VJMlMfZ9s2VM/zQbG
8sOgwc49o8vK/1nsA5GN2ffBmzHluumeUZE7vAy+XecSB+CLmDwcU9rQ/MteFL0gwAj0V2LcCP6R
PBG2J5yzGiutqe9kxHhKDIhURO13A8iNgbVeSg6VDd5L1tV/K15M+XMmuYynQRpyLtKxSEqaBIB6
XRSKiFbf8tSxjSeyhPZRqAOxr9NSp99LTIiC6kM0mQm7RcZCsjhOe1NEcOSfO/IArfdTO05/CYAQ
03lSfJQ+8lWbDNIZaVLKJgmmBnb+sG4g60BBcmRHBWzHWj4NNW7a8Azbg9RJSpjzyBexgO+FV1Td
ESjqPhKdv/A9/2osN4av4DuvUDo16DxgtVv/Pq/oB+wd2YwZy9kBYRToa12tHnr84QGhx4NvXK9B
ptN6+nGoww/zezlIIRKMs9x3y6eYnjNrXOBKrC/j5dCp1UlFJU4CJguCXy8Wq6LorUBKz3z8NwEs
Y/FdtZ/jR3OGpEWmPiunsqUnPAT69sPO3Cuy22ij8O+1K9tICHi7FcSAmkFTuJMlhvx3L6QWb3dg
Fib40icEVp5mqT+vY/xbJSiUL1GqvzmBGVA1eJcPsZc7tqF1lCZqeq+F2bYA9QzVo/tbE3i64Nkb
SkMnL6jiDDUuT4zUcDmnQ2G6bdqUD1AAFsBjU+7o2AigorTc9krlRSu0Kh/BsgMPf6FzjawP8dT0
e54XVg6D2ZH5aKIEYuwC6UxenbcvirWwGNpfvZNug3dCbUV1g5ghDeqeMtn7xJU19/IrDP/+1C77
UJ//VIGinAA4hlQz6C06dP/MYTPeRln/wLU9RceHwOvX7mKpH+9UM/6q4qG9W24aNF/hpwDKftHB
p0x9ABLXhFz+MuBLMkTJULtBK7Ovo1GLtqnSgF+2gB5kc1eA7znCAcOLqIgvcwgDv9mJoED5p1Lq
czDZ/RKuIQAO22BNjwzQC68TvecqV9PVF3vjqf01lTglAMk5Xp0zX0JvuJt7KjHAkXulHDeZpXvr
anQajdlfRRz+C2ZqytPfCQV9j2yQpqj5OfUvkOucOyVUn2gUuHsdaaQQSKEiIYqlPBgYZz1P0zOb
6CKI79o/uBUDcmOFRMmZhR8Swn6uzDfUcqP7aTUpOWipqNRMaoQvoxEJGA4il2zKB2fXpLscn1Sz
IyiHChtOhRXcS0UOznreQ2pptHulzPxHxK7U7P6hODAwfmT/F+rdj9YylhD33CjgvL0KeuwgjawL
4ILrKjly/KRdpmg5Y2bQDCFfjlvOe60nmS8ApJgPy7Ym3/XLHq29gOMzjl4LBC1rSVpK2dTy2Psx
G4hbEDLNinTqDOjnOwlIsBeYz/TuEkon4KtaBz46gj8mbDPlgQULhQtsigmPFshhoFnoiDPTeuGv
xe3juxmM7j/fx/ak0gFOEoNZ/xjFfn88VodwaP/UmKEwWS2Kkeq+/mZcSPKzgrrN5XhnbvZtPuB8
5HaKDQeLv1AjYIRMxKWvklUe2IHi2YmY8Wqwag1J9iQQ7BoVpUvRC62yGge3z/063+M5qut1CNrA
5FN6a6X5CTxHFdQv27cjCdolOhGGD4UwMjum0Ns6SPYnHbOX9p3SVrTNRghFCMkxaApz1JJZ41Qa
891n6+XRPMDWT9Z3PXKMrJFTg2na6J5l0mboXGkRsHfQNtawE2Bw3cmDjemEpTPn3u/eRAZtmkDQ
HG55HqwmRrHP1Q2ISPdGF1UF1ZqnrwAp4yLCV7tTk3whSfd+M91379uPBTXeEUGiQHhgDj5hZ1Fq
+DDK8UUkDI3ska7e0j09aEuTlt0jjnUKzle8kl3RZB6sC3KWU9EKF7PLf0NeI8NQWdCcm6Orp8DB
eWt478ow9A4g5FrymetL/8wyGCq1NX58YKmgf9KhxSurjcnri1odj4ekCvwGi5ucZf7KsFGwObzA
RqJw+ZTPBpWXXkgiAk0N5QZ15Ig17UX6bx7/PpknnexA5ia7peD9LJHHOwqGMA20bbG9ZU1+kprV
/4xS+yS0XUI1HqSbNMHx4p5m9L7x97AvNgLJ4gCek7FtZ72TYCt03TrRixQVycQN3MGMld9sYEB3
jLyRC0n8Du5+M5Jm2LHPuYSROZfdX10ezTXC/wM3f+t36z/XoZupRRC7YW5widfVCPi01E8M8vVZ
Qi1LrgPcOA/aMzIFdAN/DFV3zZIJHc8K+XWqE0P2hO6d1PzsW4D/nklY9tzQ01AP8FGO4QouuyPw
4MznOpVaRcNjMfWP+MNcil7HWmb7CxDrxsPwBT/azAqxhttmHgwT+UUjFkL60uC6alEhlmQO74Jg
pfkTtisRjAdq6gXv1TpFBadkcnGaFv8gGxXw3zojpoAhq6YgKLRB53uNLSFJx4UjpYVvBvlkUmfk
/FK+el5WjKaPiOvhUCTy7Xb1zLp1A/UOeP6bWfEaBHMM/aY7jaVA8gMjP8Tmrd0O02WRppwiwNSU
aZX3ESB8FtugmrWkxn9qLFc6k8ocUXrYP54fSEF0SxdbOyZUlL5E32bQ04lAkCO6ojkSZY9GV8sL
hfyjn6plxiMtpPFWwqLWHD6m0jesZuNfuzmOKewNh0/wqCK2/G3msQEpJvh/0eHoY9hLTcRiQ6UJ
5dcPTDtALKg7bNq02Ktnl5zWZhvd6YtgALP8u0tn96jqBhnTnb6gidD6ACVI1UmGenV/YtXz//QN
gp3bYjLpKVoqsryXx9QxXXMlr2eZP0xo8FkZTvHyG7hF4gDj8X0zgN7O7CeJwsG5qCBgBRr0P66A
Lhxy7kSEg3RhV87LGEPaDSdW3VF8nhx2qAbfyC8RrZPCJdw/D1GUZgWQ2wszuhoMPGK8QIlR5isI
zv1qO2agoK10PKWtWdDrgRrSHYs+JECQgGbuKUfNQZXHvXaZU2+OnKduERIrY+nM1A0w1cskX54I
MFjN//i/qMCKpCyEfnboI37YQEJIlw0/Q6v/6TzLxV91sJw1FJ8Z60Nbzsl06GuFlnHFmJ52n+hE
9Ss8V8LME5KEXzoZAY/nwUneXIZxSlMrhHheTz+P4+Tz1F3Wcht4HJK1d45RNntm6EXUel5OkbAb
mBv2XOCt+RYFxZtFM9iyRYX/mSg/MZP7/PU2Yv4fJD8YKsYUvXtUH3woQPHxpfBm/BO5b+O1kL0g
3ubewRj6KdAp/ebCM7R+MqA2yRrFc0ISONcgxNxr6KwI/9JkeOwJWdR9PwFTytOZ47uO3gLYKTCP
8mi5P6RQDGoLP/tTre0llF7f84Ewd/JRXxs7NrjsSEHU94CgHjcArmP6kjP6XFwzYHFLVOLE3UqY
+L+9/CsEbM6kP8dj8/oavq6qWCciIeKKB8yRVM3huP6HQ2hjiud3ILqG/OybAk2emQyZm7F488Sr
WBdEuUYZsiY4k1pjpppWtBGWFo3JS0gPwx3paqQ40mSPT6o6mSR+0xeKcwmN0WCI9vYwuh+TSCi0
6RPkGJLcgrj8XPCLsfdUdkwevxT/8Xwbz5wZQcJoCl6HRyjDT2C1lKrZYph5KJPnYJCfRJ/XFQ1E
08usSvamq8WB1A8QW+yOF8HNiU+LRkF5inOPN7NjXPFB6qK5/5pY4Qy8E6cs3fdezYFeGKDRZEW6
mjGpx6TUi3t3IRGtVXLpD0P33xWIQoVrwBMgcRk/UU15/l2vmR1dxUw8zSBFinTrrltxyvmbPGwJ
XUjvxvN/9OXlMO1gI+GaqL/h2+KmYCL6Zcby0dUhwDa8Oz6KNU2m4SUOuK+3xmgLMZAP8dvJWg7i
jtEXiZK/R8qlixeJEmNAx0HTLvlBPPSww2WRJ1zV4lsW4p/Z7DqC5U+JjFQX8iPgs7GXAO86W9zU
sQydHn23d0JBi8IzEo6oqAGwYNey9VeenrWmtuGr8sNZwaBm3aJdgiUkU+YVITPqZQgoJHOPPo3N
7zXN5BfNnzzP7zEB2q9DoR0yKD7LBHNn/fKkVjfHzfXK6oee5COUzhe6ME/Jc6xSLu8RmkvGBiwK
Ghdu0JV8FcCwTQ1XWqptnbzSq7nfBHeoD51iNcQztC3u/r3WROQwqifpOHhwrzIbfUzE8wzew5OO
L1El7op50MYPAoAHpRMjyTvKuA6AtIql6dU5ad0Po2aW7eYexCPGuxAOFwEOX61sKrN49MbC2IpX
AgTgTHktyUJ9XfcghGoSJz9aTNbKC3ns08akIwRHMTWNf+ydcpb3p98bN42IlXRgbIY1KAUUaZM5
tfxY6EuOcmkUdrv5bD9+DCmySfttxXZZRUicD5UJkTHglBhDFRb1YIP/Ww6zGrCL4t85q/JlayTA
5COZdbWAS5/J/iFC2HBUyqiiHz7XrAAbBtf5EkBwxaJbC7iz0Wi1ZfUUTnHqjD5/6jBLJLuxfk6N
vFM9MfivVkiQHxVQ0ls6FGOKw65aW8MHXDDPFeNP5Htbp5bHVqW3Jzbuq+BIvVA1dcfgsulupMS/
kEkAsk8VPmnhl2AasQIWfHn90VRXmjrH5NDDW3Y/KM59IfV7yTytgpP2JzZd6F/K7SG0rnmvL0/N
un89nWgJ8Mzrs01Hu3U1+gxpJpQC++sUQLfxuq2vez8yR3MEDGlzf+wWJ+ICb/LVd7n1M6YdZb35
8JzbtScAjrINahu3QJFWNf5jGvkZonl+/nRHtcF0bIxPrbE3ZMMDIWQT0UtTE0DzBQL1fWgot6k/
stchC+w5ExxYgexu4DmkB88ZJaGblw1FE74uXIbuSUsVFnk67FVa3CuanZKbE0FD5icYeCn45sOF
ZtaW8nZp58Y1w5Nb91O57Rw2S97pGKFtqQeQVdwrYtzm4MUn4inhso6e28JuUcm8k6Y0h8Krdp7A
K4z9CzoP+MtR9Clp2Hw/Ch+I+ngsCOmNgOMRRVQ7tXGePsy2TksaYFybKVvZkRIM3bfAlZD9BwNP
EkfDd8FeAlIHugNxDY9uKsWOVeNARdwOdOHWNkyrw9rXv0xOyVjE8Q/tTFftCJP8Qfo71kOY7teW
PuzMOCasX/CNAT5FnGyrifE3Rpu2wmc+wMXQ27vlnF5ZH8rCmMngKoKPSapA97zeVr0q4ZiqOho0
g4JBCz5qi9UvBk+WybySdpgRRdIGcLL6ZDd6xjw1uESfa9FecEd0DXlG5Dm/B1YVopiwCiFykAlo
4Jz9BgiD9oMGPOh289MAnmoDKdi5KfhPPjw6gU66/btIWMZhDptxyx8Qh/ff/bt+2JTRntXHRNvR
9fZuq5ay4G4x69i5rMH5ur2/K4D1djPuwkgapzAg78serhBxV1YR2gfXAhRvgnZ6m71hfMtCj4hO
Pe9KitnurOb+y8GCWu4JYEsJnlvYncfD6WhYQf3UAkOCtv1q7k/TGOeR3k/LT4U74cnL6HXEVaUo
hjzK2c8RJRvIoTdJMESOHouI48iUXpIBKRdajNSxeGBo5li1MJIXpA0j6uwyiWgTXJKiB3IkyFYO
E8LXWGFGf4X28JjqjJdKx/ESF+SHgk3YhuB1DSm8NbO3RfjnHrcE0JyQ5lcjaoUge6fbpRFPCXQd
48nxbenroOSB/74bT870B5Z81pFSnBTvtTlFsIiZLYgiWRHQHdQdeGHwEuIk9+Z4RbI4FZm5Mx71
RdI10qUCRB8HNd+4KO2x+OrS4kBvU31wv3vUilu+JJKT1O8Xuv5hWWSOqYS9T51jXWZByb5iRZz1
HfvRwnRzpGAkvEUSORmQV0PWU6aF6EUP/V1H61grdMmO5zYmp+2cpHhAckd5HMfUCukBNADPWajS
ZkEEpsEEmzZBHpy1ZA9EtEl3sbS6L4gmtcZrAwjOzU7ceSwiOHX4Ursvgpff4uqP6ZZGE1k33AV7
Z+Z7gXjbKiPSwkheYqmpaadiWxCXAcfRuEaLz3dPEDjtwP+TvdiCwxygYz/K294+5E7kkXaTiw3L
p2X/6AGHmgNndBkbZ/ZWTtBnbxYFSHOVK9s9z5IENhbfXwmJzJnWYLsrG+9MDJb28BLzVRNOeEqS
0d1m24VOzCgRDwg8IXPhG+mirhkaIdze2avxknaudYZWuGjT68D5tOX6NRG1KOhoI/SQ6gp+GtTD
bbesTM4YUwrl/NE87T+ZFfNna/20eCOa9yoiKWDw7+8dVw9CnmwCEROkgbPqK3W04Y18WsZgyckg
nVGg5Oa/XaS9+u+nWx666KicpYITrUW9wp1rtf4G06K9JFBw10k5/DLXc4ThrurEQT0owIxoeBBF
ucz68WEdCbafFFULgCNUN/vzlA2ei/H6ldSlx1vry9fRamr+K2jzReaATt4OFA+5asIgiWa/3M5t
AjTKYLSfmuwaTQuXmIwNGn0VOKoPXzmn8ABuzEKxQpXVAnxoQO7S7h/z7xdpYx5mRvFZ5dKK6r03
BA6Pj096rczB4dG2xczKdEIRgQ84oOvBzQ/gjVtw23uxrkv4Jsm07xPto02Wnv5VAlzMbeyhdOP0
7VStbMqqU5YWKxtUx+TgvrXnF/ouaILJOhe8GIAbvU2ISbjrLqcN5kYfUjK2U/ouPAEak1H+2pN6
xbSC9MP42kYw+HjkdFU6ems2fWBbGDCtnwmuM29+jRi2etiCBLFevAqioD9BYfXRD3BgjHmIDpua
xykEZDT0oiMDk3UUoRdoBZgYIO1SxVSv6EewYfPcJDwK4g3Zg08xznbleeis9dXelLRzTMeHPXOP
J0r8OIyrdpfkcupcTby6fjcthVwrNE+6vUr1ayO1gjC6Q45oG3U/e/mIrPllPXHAPaLYfQkzZR9S
bOu4h9ziOdvPF7G8uu/XRN+QbGBqAK2fgfrkyD9iKHkuVYyxTJ/1vdQQsyyPGGJGlzLqO1ucFgbf
vPI1vSmxE6JFxuWN0tTyZ94kH5a4kMMHnUuyIAJo7FlYjaT8dHo45BGjoNxfdze3xUobIO2VPHql
bEbvGuF8IP4wFEtNz96p6LePJ0gvFBU1p7bsaTBM8g9nqyMCQ2QdUZfUm7aBNOMl9mkgRrkGTplM
+DrczdDOp6J6ao+H1peMlsaJR3djZkzcdI+11E4XPZsfRqYBFDms1KDXu/U98yiiu6absYtnv19R
E4eejufLor8jPu+Cf3U2WsoodcW/vj+5l7VvAPn9sPNx8n6qHMUZw72Ma4Nz4d72QJO47utHyC0s
i8o5N/UGD/5yoFm7kVb2v42Qivk1xDE2MM7jJucOrHOxg5oUX2KHMaMPH6w3KzdNUGCYkinjrR4s
bJYRj2YizfC3TnjC0qzcxf2rRJLXdkKwamPcUbpNpub2xrYWKqdH6rjlImw8P+FTpwWRungli2XF
R5xy9/cP3fXgkcQ3Uo1GFqjZjMQcHZ5sepW9IaSgpYhMoCUYdoB3xu/d+lHsMr+S2ZE7bM0ddH0c
JddIoxjoXh/VXJXk0EdEFfHpFLqZiECDKKL/rTM7IDpKz9c7jzJjQAH9ozTQk+q0OOd8oEWh8rgG
FaaCVFFtPWE/GOiu+bM1AP5I2Eq2ok8SUToirYBlSiYez9Hf9arAqOjxqxrZ8Kko7PBy+a0NAb/6
j6QwlUFVcAwLJop1dyOaaRtmU7Ig/9JRt8W+oskJanDImiyrV2PXTg+SXKpUebn0CR4UlpI1Tkak
b5c0ipWFDT1XBUEvcPwDanIlPkzCKsXdI+GZSoWD9yLnicqhqKpWTKxw4C3P/PKGREalYhMMUE9z
er9zZKeuUDZJjDx45SM3g7CWorwMakh3XUoOL3Klv7fxdCJxGGMuPBjc3LPNvY1btw/lq+sw77Wq
C2QN4TbxuSGMqMT3wN99tnRCiftKN0A3MqINXuDPsj1JieCIty2zlkG3osuCtV+P0QjI/P+SxLbh
nxAx4ML/e+8aiReyRYsWMaPwmvWpzApyNGZCXfUxpsv2a5v+eSgukRP46DEnbMt6AIQQxqS72/Lc
c/6Y369DyV18IsBUwPoDE1qHazK7wu3Tl2sEmLo3d2M5kfH7mug/rGz09k37u/+B5hTDA72KcO0e
K/qR7xZsHgV759y0iaLzmVmup/20uvSNi6KCrLfuaSwpvm5WcUwj2TAk2qK+gJLK9J9oFfHt49p1
H4eYhnIrpfyP/BN1ExM6MVkFmDmd7S9m4X5jfu8yHKw3DrZEFqCYhXbc7VJHwIUFI7Qzf2sxG7y3
bLE9zm3OHLxFUdO1FbREA4aiq2M+nhKpEpa2LvFr9uy/RywQ+vZlG4mhRjZLuaChsVUvTTzPAVwn
Ac1zq9dZcAnqoFll/PAvgJqwM3AoOchdxaWVFp5AzBkc90W+Lapntp0cAOfkDrp/Yf9huOkwssvW
0ecuK8NTB8TpITU1mNUQ2F3bTr5WeFnJYaumTxS4sztljK7Mmw/VQWlg3H1KqLf7Cjat5Vxck21H
Yc/zXc5rBWjY4C93Fp4ghYF+2rkPwV4Yxk70zcCfrHMmgOclKtGsjSP0chiqouhGDQDSqEzta6sl
txFIgz6SqO4aRVbZVY+wq3KJkWXKoGD3U8B+vbtL6q0y3V2BsFbp5Ew4x/hmi1RpnaIO2U062Clc
nSv/ZAKdaawLe/EFM7F6/VTg+4LfEXRcIF7R3I69Ms3MLX+NjXG/ucrMFBHAMgMqBPw/oFFKAwQ6
9l4hfZwlLcnLKViGcC08s3Uexk+mB/gLWF+vtbpypMo9CcjuVdL3+Xyq5JN1AwI7ExdqB/INRYGM
ZRHd0X5Qe0xqvXdVutBRvWwFRjS2S8Vq++kKiFiS85kABFPxN4m7F+LruTdisqcWHkyWlXKkB/4r
2ngRAmCdNwbGX3sz9KBY8LT0BMzipV6O9/jozAPwHXp4Vk115hCG85rHzCvkjhqO9nlkcJDQB53H
kPkK/wbT72Q7keWlm37s/ZUZdtiyJrHphNR4oApWER43wv8NRE0iy4BxAf1m7L6biEEnH4cZXzTE
+u6+ekXbyB0+oQcPpv+zA/IL3AFuDl2M4bapuVJidKa/drG6sdZnC81D7Voc5q5BG8dOpNG+8WY1
z+U0y/X66hpXy3UT0hJL76eh4KNflXOc42L70KnL67Wmhfo/sRXcVZYsoGM/Rn2MbaqYDDjYWqQT
ebglSJb7PtHLFkqJ/YQr0rl2uoMAoCOGgErIRTBXV8+jPbvTilpuTVkZI9b2yFptnpx6XeeC+TEj
HMkCPR3wgauPoF4xt9EDN0pAUGRFzl7yXxvG0psYPdFgQrWhQKroDJU0Efoy5/K0IdIOQwQ+zCJZ
BW7EWJRsz0ZM+04YhR5EgUtwzgz3dzWElTXhu7sKwGdrnPUR0K4xWNQxi+/DEjBy9XEljZDWO9TU
jcTH3ktzT6DHOm3CR4ETpB84uivuml3slY1Pz4MG3FRx/T/7UW8jgHZAiTJvqpjYDe7gji1gRcwt
lv8cRjQs29+0pIe4XNecWMiFbdmEHu+UsEceZHQ+5+KmsFgqGZud31cFWNc+RKMHIfjatVHoMlQr
PugPjtaDuU+J2LTHzzr2gn1v9Xq7ox/Zumi2gLJCUXWGp7xQJc06iKb2A54SS3U3ekd65IJPGYJR
YpqQqyGGvGmF+8eUpcr8VVFnK3jy01ZCdgSdmHXgxYeEdlIX5Yl23emaNFkIli5MtZCB5mGHavAG
73wW1n1bAfd3vEkK8SVCoYyX2sR0sqF/pcFpz4T3FLlJrlEVouYibf4sWV6Km4Xqta3oFPiYZMZ+
quf78nCFHZlw9VX3SvYLN90MCjG0rQsSo9x/FhrHaONLCukdnu6l47N/64cNiuG8I2jcE/lXCJg4
IlhERaVDJLjIAl5S3VY4M8IyG5bEWVpDErqtld7Qs1RRmNin3OlDMGzfevZ5rMtv0W4q7mX0tmn1
yAvuOLa3QO1FqUbLG26tygOThbQalVMgvZxUudhl9HGkg3HICw5ulZvo7pm7hBXDXQOBI7sqRWpF
9Q+hWDZFymuUfw2OggNKkvS2qD0wl65mKg74JrkLBreUaNgAZrj9lthRRH6h5gyjgcAR+3js03Cb
lMG6ENN+0HoTYxALG4NzTHEsJmKkF9soUkjhyLNNFtuoSK7oNgc6XI9rIgiDy1Y7T89aUXH1x3+D
yMjXijZrjHSNrCT0xiC3yndrUqDTHivu3YZZCA/Mw/+mkvB8oL4O1VIzsDZhyf6Z+LLzvGdr25C8
KlvL82qOgD8onEKcDzpAZU5tgOCVtYiBp74jx/yyPcCd33uS1j5ycxNYvL87U3CGQ8f41l9RVIQc
yimv5NouWKEM3r3ZZpcCMe23xP6k3a22S545lApLgjPe+y2GWtBttOwdsBfq+MWkJ7ZB/z7Iz3I8
sNWg5Uw7iY1cK3G22B35nGOl/LEPh6i7EuJZbYI8b9VNAZM/OaoMfof52CaF6j1FO3WruZB+SMJq
a7ITfuU2EWBVOdbEJYHtfLT2xdU7Ct1SbRUVJNIWx64uWwQwbXeXdOAx/IHTZgs5OZ0G/McQkzsc
am1F3Rr2uncV1jgwdXZlWMkUft26aPjj2y+DAsuxs67ySdrRkSXLtt5RogRCceynCG14dWWklILR
+nKLvfqX99OXgI8W9lwwrKkf8VE/x/mmb7QzVSblSqBwfGqCLtYDdyS3HAuxdBZ591Nds4cqj2Wy
Ojb1dss/3EMIJF0Nvxg8ye7WiS5FDlSX1RELFgdvWh6OuGQlpd7aE/Z4LrL3UtjaNOYO5wOALEX2
k53tUfyP+SKLt25Z8PfRfq94fTgZZ9ecVRQm0LexZ8OBVhU6vGi48p2LyxLwXcui6xiK+6z5oFl1
K7x2c6u7iZel58xgim1gEWvK1ppeE76rKOR+OOh8GaXIt2bAaEtu96fsMBfuBQb3N9BrIbtIT2Fp
g0hDg/LBWR5+LmgnMnTs/Fdk5ep7FlklTaRg60FrngaIvK61IZ5xrsezo8H/6c51TAp7RyVK8hfz
8KuwpW4ePJXp4iNpQwmQf/afbOsCGfh/s5aPQpJgZUUxGpPANox0kVP/swKubh/n7YSZ0qfi/hBE
sDublxBhT324f7kyWCGmVjupHu2pT1bBc+W8Duc010KjpcDHOjGBRbx5AW8c2Vv9XhWtB04PUXzY
SwyDNtu53T0FhZYU8iB2AilUmepRk4JOxIYaYC+EAh+5/1mcXOuSFjDAZ53cKuB15ICINb39Sq0y
p50Ei1zm8eyMck4N+QANf9DTszNK+164liLhE4Co7RWO/HS0BDCnw9wspR9bRBoimZ+Y1/MLSIpK
N3X6uO6HijF5laEDf7b2T+sTmi2+6NWaWjeAodm3uPxtK3NZ08ytl+yaCJnaJT6thRdR8hcYwHKf
RUSM6BYMACXnC5sPC52PP0YtIPy8TnPdrVClh1PscKGozmZ0EcD3aZtQuuTzoPsIvgRCcknqZynW
XcQhE03KyBk+0pZd/NFPB7fo00QACG0nAR6xsy3T4F8U86mCRXarl+Yci48vpJ0dwfoD1fu7R3fX
FKJNAp7pB4F7D5lcYTj1JcMvW2ikr2xUqNdUE9bYKyA9QCLYsVGgjoW5KqpiWJe5/MQum7kWjNjV
vf27xJ9Q/oeI/QOjAw64tSCn+DDzEu8JxZJmnOEe9VFAdS854y11kLtywIJ60Rw+BKhgaAu/ef05
P8nF6saQMg+ghECgAkzGDjK+BJFu+pYGdACxjH75z4bN42+tsIfOEEJJnbglHRvNJHE13V/R7B8t
/6P3/l1WiPpq3uv0ni6yb9toPOJU9g2r7UbEdty2zEmE6HqMDEyc0ogh0GLKRN9F6nmlY+ledo5V
qcDbopY2vOOsS8SdJlo2iZIWilD7wVwIsfAQhfT9X3WzI/Do8mX/GrZQOmXtxMt0BEgul9ombelF
Ld8vUaKnthqjTiLIq06D4BE3BHz0ivQAKPIsAu6xh7lWOYH5xcJV4CUZIjSz7t6a1M9twb5wkRzf
9hc0KdOEseV//s5yMR8XxrVgBUSgSWElbkXrH/3rANVKc1kqLOHsDhhJ+mqThSl4/paTd81wfUSt
+hCJWHZQEFTYHxO/QXKkXu4ker+++P9dywxPSmzAWULv2fCfPEODIYBWW/8XiKWNsBFcW8XNFD0l
6HkCGwuaCYMxykpRbie2NwKBrUMvfEYiCM1XFWAM+ppSOqTAQ7ZFZUygUFs8jsDfseIm/CKfRYfT
LqFfPL3uJldVw0LMe6DQ0B4Av0bBLcpMWXB+kz1AI0bXSFBJoGTOshWIJsifyoWrN/hRnGWVqnb2
JYnJiZbnAt2UXafW99KCeRKi7CKNU8aglghI2DcmFPcSEdmwXSpF+fshTP9+HFwB6wr0u3/hLnto
4cOB57ZHSuec7D+5aLbganMz6P5NEZrbVToR2VBQxYLEttS7xGgL2BwUECBfvIcULOXzCLGNiX4G
DtzsW9UTguPdZDShpC5oTzCg8N/zalW3CUSj4NfwlwaFjPSRq17EqMjMsfFqrpQAXoZAasrOPWu0
tEZMQTMBllR0pVsvlH303slNkzKYjiS8dZMflRARrZ7Em0rnY7uj1zyfIfROtBKYbDG33bN3Hog1
ZqpEu0dtpG3xTeMRmwX42qrtqoF8M69KDqq/pCqygVaWepI+ZCFtcPiPeGbzq/lei9c2VlJ/OSzd
pFIoKLP433r/IW4oVtnrKgY0G4+sLDPASgbTGfHlGU62HHAKmquG97yJ23OZY6Z0HKkmsmETvi04
aAKjZV2cAnpgix6DjW7mGNr8bvqAjE9P/4AWUDCzluso6RgH8tt27+BcATu/D0S4m42TfwDx0Naq
B2agE+jMbxS+70jPHChGhRXMByxc3R4Eh3s9D+98vjUGUaxR6s/rDcf52hdKnGH2lhnjrQO+u/3/
CEAqYicUUeD8PqpBXhi4cy66rICjU+eaK5e3/NoLBPGWagNXWSd7SfCYeXqkSBQJU9AwXCLWLM21
USjPeGjrIQG4No6ByK/2vXM3d8BoxperT7jGGqITb9Nupt/tkoO9O/TaYMGeVqHcEa/xko90KZrS
87Dbtwu6aBhFiFgcLX8Z7srDV/t4FDb+dTe0iLSThtiDrb8BTdjtAgPxh9HjjzgoKyVaExrhPeRB
XIBE2E6asODalndxlrMXm/oV7m+rQ1tSGFtxjF8YSkuq85svjKnJHujxM8hveOzLpnuqTZifIQyA
P/D92da8FLbqxcYg0U+KM8/zIuRp5RGlnxHx1NGurh2jv6iPfZRGV702OIcBXQwCtgFx6qB9pJZ7
pZs/dkkSHstyc+dvtYQPeXatHQbzm/WF09k6zeQxIlEDbwCVVnxNvrmueYxuXw8ZVtgdren8MyOg
BixTRIAYqybIGF79D+Int2VilxB4ED4iFFErT/ZyBg4E+9iEMgk3WuhFoyAJYrP3/Xr1S+YRHNie
tv+PG8SLkQ8F/+k1sWHrpBk6ycYU0Jr29V2zjMJ2m1SkbJyfQeNOHjAQIQH8ZKvFEdqwTiM5VPGe
UfGLe4u43/n3HKLL21GV0ZwY+ocT52+08hLNQlM5t7oEXbQnPGsSaMYAd6Fs9CVCvRSdJxXj6wJM
m4SrQRw+ot035BgDtlHs/atyloCNcClWlzaAR6/qeXNTqRwoo7I6xfDOHGDM1x4TtKMWPCwaIimC
9e8FFnoKFSDnAMSB5/EVZWFSEtH+0RbUEIsJ/I1mxZtw0NfHE1lUEJXW1KD2KXxTTQj0jCbVx2r2
dUWHTGDqng4UsjN3LzoitWx+57X78D51vIhWOEeoJSAHux6m0Ca5pEQeMM5UHhgcM75sCAzoO6w3
eP1YLZT2DBOyEc1ZuA5bDZWVjEgFi0IcwRPUTKqQDmUqWXU2acL+n64vGIoYhzj4LwPKg9ouOlS+
6sg6O0FnZI+goPyBjM7ZWCKBHLello5d048MQyrAXtYSBv6rTikYwjipYRXPLBQdIkmGO0a3QTcI
+YsKLROnwNgRR1H4zxqbyFkKeDWjti+mtC7le9xpRr+a8H1sqLtPM3B4BHyRd26AZmYmLci1fcZ4
D68fhAZfVZ7Y+FZNQNh0jwl+3vnE4/LTakim6UVZoIyz+pUv6gFXg+kto0wmlWJVFVa2sd7f/tC7
Fu+8vyAPPMMrXa+gtXwCi3OJGnXm8Mi/XaYrQPKlj3XJzM81cMaKp+3emnE6/1ac/CTlaeQl923c
GnNUOoJmtxMcahKBwqBbdRqWMaiSrwY5ePXKyUnXGPHos+lgwQmnKhc/2JaLxiH7cce11NVwF8u7
5VRtzRrhoIeE9EJPJHcd2oUa5L0yDpOuwbfFg30+sBXv2Wib2n8yLvpZYwlN0F9z7EFGFFZE5oDm
fwfLxVoc8WZSyOXhew9+91cHHCwWvqf4CFF8s9RUf6bUlEckeldDzeHVt5ZpvgOQQd/ViuxZriX+
FfgGozDUNpb5CGs2AvDfJI9HOU6Xs+exabiK+BH8tz24Rzxyb/Cn/GvNwDn5IfdUJZ8IPq4PMRbd
cpX1gdu9ewuZCLV59E9kjygZU6VVBfJoUniF2L2nbX75rvfVJDIInHmayKbO68H3lttUqSfwQDiY
DlTM7ZH0PcWyfuMFc8wk2K+buC/X3UrsazSQPdXy+Rce7M895iVfKac41RO3oHUoMu8gk9aJg6ig
sK5NfkHc9ALyBvGTb1ANnH6K3mqVYi2O4+tMhrJLiKR5pzURdMp1WuVbIDK4mnsZlpt5pN8hj4zT
LvSXDz+caqXtmaXl718J+pSNMUpIY7gxbPh3IqoZcku7klvWVDAK+2aONRHjbnbZjGU13QwAnIVx
A827dFVIyl2trXgLufJguQtUtrtW2F3jzdJwSoNSCwOhgYEt69T8ReN1LqAqAciqjoHjpp74iTwU
Dl3QCEy2sS2QGJBQoSQqXfefwHnD8fYOjw/em4HAqWLDFKYuput5A5OSWcFsBahqCOKUSbeWMQt4
W+dUKOlFjMyi0OJ8evhULTiBkhqRpPJiBbPFAqCkeOyw0lm26Ws2i2fq1bdFN45rgttq29yiEq0K
7ZjR6IgkFy+nKAR5H6rdvI+nMkzfAZSCWQazptwGY4zCzlgBChq6myhnoKc2EWYsoe15veb+M3EV
VlIr1ZGn1eDBBJZEq3gppm1nh3bQBiKDrZI2UqOBa2wuxSgXotOUM3e0ft+OdUjH8u3Vug7H63Br
xzcb4ESL75XoDvPmSoj+peTShmojvjKBxHbnjo1ZHb4ovjXXVkNJTcro0NbEGg50TWFB+yggHq5k
bEN4yC1rd9a4tsw5Hnh79Wa9k1DytszFRE3Lki2s5oTaj193wb0LN3/u30jlhNBhe58tXp/ofLQS
g1u+aNa9umgW4/nnRg1TkI9IXguuX8BT8ju5mVT1FvdiwfX8mvFiXNOb7WL2WQ2iWSjhmSgFW5L6
zBxF8njgEwt9isNLJFmwen4CgH3T4f4pImeWIMU5mgDUTx5GyRzIFJyS3WH0qbKcMGNwPTo3aMsm
g/23LVrZL5Zrb1B9y80wYl/B6ETbNYCuAoj26DyKi1VeKOnOlkglyOK5dyCIbH1ciu0H8L5yNF2n
wNA0yjwzuBdrPRo5PS1nviczgdEwp7lWGSR5nHSsq/cDQOi+Dw/g38KT28Qh7LAQt13UCBBjuWLh
e4WIsqRWTT0fW0+X44KCOZWAm57QWuxjtmnpoZ7eh+Vqw7OVR1XsDhfMv76vR/HF57D6+ToOU0se
Ix1+rY8vTCHV17n35Cgt8JcDw2oJ/Gu4nBqyaCrryJM2hQpLPujndLNf/62G34RypH/zozGepVmV
9vQUsp/GgQ63SiOA5iu0PQ0AoSNVxFW21yMR+Xhc3FY8iYsRA9mcrJsK/YzmP1q8vv4izyL8GHxK
tGfGLWRL3u9pYOj6/4LJNqG2nIeDstNHQpuMEYb8LsrKsy7ZxePFqfAuLtyBu3LTcaKKQIXGXhtP
QtiUaYXZHE/dp5hBgHGOceWbpMKFfQnR3gFSBt2WzGPZgZfdrRO/N9GFtP9bBKmXBoppW0XpDFNR
Ug+K50qmI6ooIAILC0AsMCyTvVHtWouIwR2JgwC0JG2mmQdyO2GGLrbXMZNXe2cjPAYNMc7OEef0
ZZRrUwfW3paQBH3/U16u6+EBaihsJ2G6JZ8ym0RVfr8ZRro0fgDdgy+9u4Igd8CqiNLWX/tC+/oa
8zWoYUcs62gPQ+q3sMM+QLdSJZBFTviBNh/w/fbtkyVP6xeWF1BXkZ2FAk+MoNfTY2IwQsGWMW/Z
61k/+cW3kKWatMSNQOyMCkqEL9ZY5xQ1Sp0zIhQbO6/iCXuxfY5HHdkCeDg01lYUL30EqTOm2t2H
l0eS/HBmVTPDMd6QEDQE5bV6Sy59XtHJt+rxAKHSPDPQzM0ikmDz2rb1k/q9DlNHE4RNfI/YCX1N
H0sBgvJyeF7zofdpQqskRlBAxAfqhwU6+kqnuvHIk0Ke+Ca+9iwstHacm+T+yZWEvriRquB4r5z3
9tz5cH2MBeeLwtGBlfwqVWOPdOPLBPEgu8y8AzrfOl06nvtqCmaAdYDN719IeZ6hXbUBFbM0XTfq
MO9arCGfwNJrusQKlfmu5tR8OYBp0TQVvAP5+N9Bb9X0Ta4mlHQjGt+VXwmUx6J+RHTHklDd50Sm
sUQfNre+X/EdZYpsLQ0ziMLEvB/X4ffcFuOsvzAQe4EhiZMmwni/Jv4ZkJaHLIQr3Ynj/3hlbvKB
4ZmAcUYju/fFdkqRj/dtj/sg+0BxNC6wP19iZe+UitPonIT+BYBPEdPO4PTHNmEKj7vsGg5dEcF8
vcCMMcj7zPyaxk7eW1Tk/CvtQf80CuEahC511LRikZiEFzAq7I97EI9cj6KGlZSiCtPHeQBFjPZ9
/7N7APwxsPDMd0J2knVDdeNFA/cCwQOODnacJG2SqONDxDzX+avZGGy7Z2vuG02X1Rnss9pakU5d
l8u9qVo4sY1NweScqXc+KWO9ts5npiDcoEIu39BnJqb3dsShK0J6SvQrSzIFhmxBtmovkmyA2tPt
tQAutjULirF7gSiF8K6IMjBycniMR2ensA0zjvLxMl7m+CRvrkMfv8eRXvXhJBgmWW5C+zMI1IAO
3r9D3Ei7Zz1Xo3tEtE63eRFuBUXwp08pkFJQ0kk3GakDJGD+Jwqln7KCsVhZA64e4Te65Rm9kCzm
hJJWPRVrBHmurGSEzcBuuGTplD/cBG9QIRTxxkFyU03ACAdG/ulXB4STSry3cASodDGpP/L31iMb
kg8B/M1xkl3PhjMWXVcqzIDX68KUPUSKX50YTUFgEUUSK7XmtMRxIo+dHn6uRbg7pLSk4zV5O2K8
JxW2DREN31Kc0A+sWP0avGzte/8dae1uamyyGxKM6RP8Gsue9GjjtIyVzdfHLuZ0vVpW6Iqqp4TS
jPVP7zbbCHV8N4UM4bCqAk5Bldn4rZ0+yDhR6Ffog+SQzNj7Jm7VmAGithIwsSASPr+GAtC1S9Xr
/pbWzs3yr26PtGjn9K2FDqAyVmGj2AXZ0L4uyh65w6jvKR+lQaYgn/8T0NsNdBLxBjyF0I3dulxG
aDPFoMWgSp5GSiNwYzlqjKr2mzubJh/67aY6NWIo1YWX+r/25fGzR5qteZnxJazO9MJloBkktlDE
BE2nWp/jNN1ms49t8DUMaqLGYrycVO+JpcGYeAqWtKlx8ftDp3DxNBSpJ0/xRI/6ax60qn6n/yhg
e/qvozXJ/ZqX+lfmKBFd6BqkhNkzqcRorUCBN6kDG0sA+9XHNm0fg0e5JKsABThFPojmeJn7cFkM
cRzArqFDPnTeGKUrZSRLkaXXH6sWh+btqJHzEixXNgEkemhUsqj4tl79gZKDDgmKTifj8vGy0Bm7
89snNqWGx5wFFqApldQMbusU14ShSqP45wVBNvfqV1NffAyD16n3z3WCHHqfX0LV1JLzKIgiBQS5
Qk5PoR2nIG9PBbKYTZSZA0Zr6w6yJWDDz1SwRr3pWptKVjj5JuFrOHG/nD/U4f4xdo2mChSh99m2
VN7kyyou5J8UgDZuLSwV83jXDprgW2MyAgANqXEQXUdNFAgHMx1o6EPFQwvyTkekRnZ0VNBAD7oW
64Mc8x8dsUBEEHwQuq4ioppw7IcQN5J3Hb6Nay6KbyGMK64tkektAd/4lXGvfDepUO2VAJ5Jn988
CegCLh0XZN6mTv6oO/JKdipj9fVGU+sxM1fOwZLqPIhRXcioionXGsNKHRHOX2VcwvCYNGjxXxeu
vZU8KMcUQ2j4Ys56SfguY+zSnSdBw3SQS6tCTgINtJ+gICUm7qkznFXEGRlq0tQHg6qJ1SZDFxJc
eutLxgwo97n/p8tXS2K/AUGwPwkLWpnD+pTyYwa4w3/i+tafw4jxIGCisXmaP3hp2RM+nCWe+WKF
v0fLr5siY6di/wOkvJ/uRpfAf3nqOXf4KxoiCKTxozreSUXthgDGl1+VJCjEL0Xxk73yeWkGSPiy
P3vFwoJQh9nZ6bXpYHU4CZK3aU7PeRJ/PGlQRLdXKSUO7tYgV7muS2yp/d4VV+AmUaKRVJNCHtBG
ZUjjMJfng87BbnvjhFzWEvnhKcZni6trWOsQtLY4Rh3O7Sz2Au3zbA9KIKWV82WeEGD0rqkbBXey
3wOXObPA3iFSZsRFmfLPshjZ/fqi3pAeNJz/CJSKrVgrD42yLuP9xBqIjiZlfrubd4lkBhHkk7Y6
Mf0K8/CdAkaYryUPzyVUk2IC38AzjSlzhxX7NerKyrL1D3gDKLqIYCksfAZLdBCj9URSWGNdM2Hh
tiait5lErVQr0ckxbv303nsbzAmYXmXjnAmSZiUVW+WX6uRW0vMNqs/fNNgQOX0TynU6X4VqZEUi
6p+OQANVSRQo64XvL/8I/MvdMi/UTfeWQK61ucm/oGLcimYP4BTCB7whE3Op/UVa1ne0hDEdGx2J
FjcC4b40RVbvbwSWc6XMzE/JV2EiQWy0kG/jqhV3TIc13lGys1BrPfivDQRrH5NHT9IsjTa8a2u9
cyVONO/ctYd/mJbyJucnlOPDGTaY0yiM/IRvs3ezH/QG2GAdCgD7gCUJyUQgX6t4DIww42h/wDSL
p8siz7+YWoO9rALxqUVGrd6G/x5yIWwfyEZF6dXsv3/z5jvWE6hUs1vlcTDIY3AKb9RCJdv+lKjv
MDViXPV0Gb+GppELie6bQhRPF7nR30y5UfpNwdD1KhCEopWQxWaOcZBH9+ARMW2v1X6oihMbVX/C
G5Bc1+chcuVjLkBifMug1qk01VkTGdtVrgB4jazezakdoigmFs5hvh8GPBqcJvXIq0QHHQm8/t4D
YSDwrNG9vUGZVha/MgAi55xC2ZK9bmeyF0qWewLG4uLwG8WA8+YApjiJ2kReP42TwVllCRY3Co6p
ue2vovV4ttDTodNW4hPyrCY0It1p6Ydrj0TiImDMswCK94GELpXzZe4OJk+796Za2tW1QCHqednr
FInarIxWzlARpH3u3keZxdb+gR76emwD9uzH+8oCikKGVFqH+4ivCTNFHyPFBGkrjUodVEqNR9YI
Ol6l5coaxLOrZrrjCdJfUUv5e6HpOgEak7RZi0yaaBop5V3jFwo7sTGFpG0oW096aTPZIjXfHzAC
LCCFrFOfjeqhx195Yiik3necSxrfmPEpTA2kMd6Jol2KyUDfcH9+kBvYc6vPQw2TsZLO0Z9JzjkD
CzL4lJ4JO/tYtXvW0RoR3wNQdljtDE5xw8ZKr3Xe+Oqqn1lwY0hjO+t7BiKpU/bcSBu0UxrMNT4v
opABAB6mrYRUWGuS97gX8zfc4H5lqSP8T+CtdEX1Y12gh0vcs6vhfxGcvucpKznINJjRApQy6ovb
g7kJMKXcASHbGBAIFr9wssiSse8E2wAkYVGYHA3JS/0F2aFvaIwgAOc1kpynxJ0HM7d1BA/BAPPw
+ILQ3TYbz1fp4NjD2y+0MdTwbAm2iEEVcLQHqmUCABtemjSBKZ95pH6b0YbgExnATG4iTR8XyaX9
MSrTccGPc/rDjbGXDeA1aTFXUSGYShUBGxMpJ/0JC5A1lGCB36acJAh69oOItPge4LxxWKO6aEli
RwXaNYeXfUYDITZGaahf/k9p7uFARmRHnPHIj3lgtAT72/ZRfkxudIpTn25X3ysI3BLYv7Vg7YW3
Dp3/122YZRkdwdG59f1hG228yhWp6ptaTVB8sUQ+hgxdgNgPcqTvYwJaZobg3A1rdtOBGgXuISmX
87LqPgCnM7qpL6ltnGBI+lS5ikcpwW0Rlq8Xk0AOteFWvR+VVb/4j8KMQlB2KnSgmWg7pF7XZ8k5
2ZgNW2I5igOvCHVIYG9A5JmQhnTV9gqSnHHLcDf+hp8aFJkMUTdjwBmtQ2fogcreClC1mmLav3J6
i1LJWNsl5Iw4kNRwsFX+gqP7I8lhqGqeNMY4oDl0dWUzI2uJuc5hMRv7gcyjCv35qKD78tkT/ds3
/tU9a8Y8m5ag05R1j+30xNPjBJ8IWwkaaBx/1qaRp6OYJh6HqJYki7PPjLLMu6o/pfiy6QPbdnWo
VBDzADJV17ulWKuZR5AGW988exeXYjRGc1DRWPxtEQ5j5oWeI61i+qjvqZPXTOxcLRZLXH/tLwc7
muNFQog9SHw7a9lvTud7/1bGACVOHcFO+prZXnmKldzS9R/COYsRftmo5jPp5QZt9d8O9mUA158p
V+p7LjzF6swDPgoDlSPGumKTBVJQWIG9F/NFHseg8SCCZJCdLZdk98Hta5eCZoSb+Vg/CdWI46lx
1+ELmn2bCIUHLkpSQsmsNIMXcG9pwnG9YSQ9aE+7YUXthjjC+uEb8dPgCVlKK0epchnBGcNZ+6hN
jWxlQqCXBtu8lXWxC3PP6cJ5kGua2vRWafNrUljwfEJ25kX9t+mvxBshtanS9F2IcbbyqOXo4/T0
ZWcXJzZr9r3TM3uAcXV7dOYZ30C42J8dq3WEy7toilH0qGx9tAnuIXPNLIRYvKH5MZBRqCElMtQK
4UIi/FuD8EBLqrgC9fa4/1QY5Ze4jYFKzclY3z88rH2zxwbRcnMXHok56ZJ1iu548myGDBKpPBsN
UthNXAkUcMAJrnWhDx/fax7fghDBLqRDl8tjOhxds1ozu22f7iGI+SszPU/NIiTiMEApKwavZzMt
iLnwqVYmwMM6cGc86N1UsnndEXOWvTC2tW56YZHkME+HFl7MuIsNSfEonURyXN+y/Ga+2CJoia6n
a4EgF1QZM0TlPERyYBtmpZr1WXG77iQ36dnyBGRUZLOALCx2JXLSvl4AlGEBFTuMmm4rUoCm8do5
qlSYK97WvxdHQiDd2Y8VFBIu5J1iJ4C6E62EnQNKNpGAVCwxuX9khGkBREC5LQqb9Q2InH1LxD8N
oxcbXh91o3ljJtA1foH0Kpp2upKdtWtDe2Rf+EwnfSF30wYqMoK73jE0Rc9FQuBiiBouJIYHDVsL
3qwZ/HHZQeX0J3o+Tws9JT/rJ4EDSB3tju8SpZyFLGvy9OnKjdEv02vbk4zZd3/4SmbjtraMcfiQ
w6EzNV9HWysNCIAGknMaCvx+XCOh5wSRbN+qOaEvHPsVg4q4OTvYoRZ/BS5BvflCW0VtixNB/nzE
jWm1aji+/FcKYIw7zwVVTWV3z45WABXtG/1NYHs6M7lOcchbgrCbM9Vkdw/DsqTWP0jCMBBWC3qH
CNhiqv0lkPXZxinr2Iw/ox9kkZDgKAjkDPnldHEFBebVV2kt4VPXmsOb7d4/cSG0b+hhGus/YBhZ
r1SuHAR5Q+mYR1noD72l4b1m2fQG/OrdHqQEi2dzb7mCV7pKDJq8lgbJwKuPHJ2Qbtduha+34xem
cBVKmma8b+8Xvq5X+zQ7q/WDl1i9rhzkjxjI8KMPCx6b6cb50msGAg7DPWrZF6isHQAS9f2XurA8
GwaQXL6jyarNkvClmrtc/A4p8+1eql8/qpCcXDUS9aSe4RvCtuaOmhzLL0SUwwmCiFXr+vjZdBtf
ULhSYxIXTUnb1/LIkVMH3elccul7BQWUV+o3/qtnwPIftoPziB4bxkpZK1XQoQ0VyZ1QqSVgcc0i
Njhqsrt2Ywg5fW2Ig7YGkFd5vOZqGB6CAUR+BMJoz+yOIGq5aiFFmYjmCa+9Fc9TPBQhm0UV4Nop
oLJRLpe+ETV01iYBWa+6ns7D96Gze+Ts8hizyFSJuON4CtCVVU3RcVeR8WrFiHzK0NxuSwBHFkcq
OC3luKC4Kr9BR5LsvnsSJlIHRDaUkYv+/QxvSVhkCB4rXX0hVfiHYP3r/d7Po5wiBf8QY44qTvAY
/ABUsKoYDG2xWKSavw8o3fJRd8quma6zgX5kbFZ+BNucq0bGrlnk7EY407u8IAjkfKf7H8NQJULT
TxvhHbpcd4/hRKShzIbKPCnu+R9KfUeZvToLFNo8y9DxY9XPwCq2Rr6ucsG7Cyb8uyvdcyyS7Y9Z
ou+oaQ0T5XuVkpyaqYitJRIQHtcYCq4Oxw/WAFKhcFTp8N6UXWEdHoLDmwZP6s2VJHHXfraw13PI
660dFqiSHeWs4Qr9CExmGJBNq9LJbcygC8tQkp6AsFxzii3aDeFWoAF/iXQb8P6Nckf0yTDCDeyl
wftyFvPi4ghAzKKWfH4nTyfT2GsRs63ouy5RCuj+hp7KXre9DId5LaEmxLLzsQPdODoREiJhhMov
l/+/E2FVqhzjm0M75wWaDIvsGXnLdYP0UmkqCoUSTlcBscyBRnkQsoHx/qXUyyu2CVaOitZK/1st
3O1YwwluInU2iGcHKlD9nM3WjhE4dqyBBfO8CZlmWy3L11D/TWdA+Ft+j9A3Lctr4uFxc8CH9mGK
BooMOy7m9u613+e4sZw967rm84obkqjqDA7xBvvLq66RQydMZ+SyQI3BHQoxsZaLa/2q1WqwBqai
ep6KLTLoNaCetaI8R/JIAfv9KjsmhrGi/9dxH7XnfvudxdWEpECUaH4FZ3CGrPUz29B23m9rbp1i
P3u78E4+wcGJAU3LtwvWIabIOdgRq6ijl7d+p+cIL6xVK+pQ7mzPdELsykEIdT6AT5w90yOxV564
ZN0IQNH0SMXatW4rm2zyrcoM21HO6A7kI2GKclyw90D9oHFr+sRxTTdRE9JKLCJQhtCMJO5NdQxQ
qGdKsBqQuAdOA+76dN8aBBjROtq++sfNI0hH4+69lJW0wH6m9bydMlXSl1DNT8Ai+21PM6Og1eRE
CSGKeMFaMPUXzJjRYWnbRObFAIlmBOeeROP6HpH9Nz8OZHRmyydK5EFOLrdesngRHsN0a40f4zqT
EpOCcOdAJnmbn1WuOTwoA8V1xFYp2CihJtntc4jL2OXdu1IBUs7FyZ81KKoiw768Z+lHNq+HtdtW
zduXZsx5oM3t2gEX/4FQ8mpnxubU53Jv+uEgAgAsRw0sdLpyM9sd2uqUqfsAEUnthSJvy/hxz451
sByNHxZyphEPeke7P4tjza/OvLls14WPJJAA6KTjXd/aapITurMKztPSCEwXx7zABMjlIugWk31V
nStZcTH5xjsaUIG3Zo/xmnR6TKyOqn9k5FUQSS/CyEyjAGt/2Jwe+e24BkeQLt6Y8xdlMq5NEYhR
6tFe53I1vp8TUZVC4uVdNTj0my/WVKMuPwA1GBLTEmWnseIgKXKPtdVHa8teV9t75L7M1LknqS2G
5e/fxsySU1Wn7kIHI0yhLc7jnRh5WmR+izNeS54EtjEDb4g34bY/IpbAdbKiKWDaEHo7Zx6Tbo/f
ZoNQu9itMafoVJcWqe/d5NmIvNPguxA7rnJdHh5+YcLBez1LYoAyy+o6Ky9lsuHMNehO5l2N/Kh0
+bv4k4xYsfAbRTBKslQrFC4JqwPTW3DXLWt7s2hNnqML5+40scsIRtN8U+Gptg/qrr8westv8Dpa
ROUp4F3PlOBmLrqmmbrNaRvWGJ2DZnUTdTio5q9AWHAul+Ew3B5IvHgKQWCkvIJVtrYwcW/Y2iuM
RNVHdKpicu9lv3moCNSuM921oOxGHaP2OiJpRg54QrOE6INDdGeYjWjufLko3fxYs3Ylj+TKmcgc
9AFVPAv/b7LcPoR2c/Kigfhec6ZKGyusWARcuUes+JDsnS7chV6K8935SKaajiu0/FeVwYGrbn1Q
bzRpo47DPheK7e8zIEpEd0u9/aDDyxikQMrSFWAnHQKNCLhA6zyRLpbXI2xb9XAPpBSYY5otL06i
NjmRHYCRWXigKBiEFLoHjjwjMfLnvpf1HtSgolCnFrVH2Hgc94cwtdeQVoNFvP5H3GtHJ1Ivs71A
JLrQd5/0VHsmK42Y71+o3UYe3NgSEmF2+FPbdtvE+ePIY+UTZhZECN4AaQ4hZbroq20V0erKFY2X
1QS+20W53l3t5UhZNYpqeOn7N4+s9Ft3Iccp6X8+bXz+K7QME8vbaFkmailHP8MQatmd48FWV39Z
CeYZWliHRu1+WjKzNMjlGn3iXUTarQNi5twCmFc1Okty/awaMdGrPHM8gXxYJ3Dy+hDAY8OzymeD
0K7xUyrMaEu+0Hs8L62E9FHJsVUWq2cjr5+p5JERnBfMQbJRDqT2dyz7DYsqXkduTgXRtKtG7xvO
cXuUcJBBPVHoPjyJKJhY9GoIhwbaytdn5IoGXHM00psGbl77JbHBD9PGvZA+F8PC51h4EAeGbDfl
+/1drTiv8faIEX8XTx5FOJ7LrtYL+4LREds409Rr4CduLeZedYgWfwhj0HwNc3Pz5bgdbTXQ7cWl
VBaf47qj9Z5qYhpVJC1NSUqYZXjZbIb+xqdy1qZMJatv7zmlTCkYdlMiZDoopikLI1izuqmIkvGe
foaDJYXUr8uonn1L9lUM8fgeSaavo0iEDI5i+GlL8f6oaVUkqIriCVfNpzD0Kd1y8qdmF9vgPuoM
L+zpeDAcNEsIfoLn5d+gtuM8SH9tGsH/jNqHxWvShue7F+UMszzKMGPOSs76eXS4BhCrgkLyvvPW
JYA19hWAw8kd8b84KyKF61YMr3Gnlj95E0uM1QPlLVzL74JEHVXNXCkPPL/BPkVpVEz7F2ZsaK09
0KC+cm9N9utDtOf3j8HeOlttiHz3TIuRKV4v6qe4pNnE9FCpgWgKPA+W21/f712uV4dY9TDWq7sK
GtT06/dAf9S2GMolARqjTMz2IGUUpzPwCOOGGUHNTXIKWn1elw3MCP+Oog7K58LmJ1xuFmEMW6NO
T60hFczaK8bdMnvneCuuaMrho+fWsOjaiJQaUSpoMVlx5lJnqpKHeZfzMQ0CSkcFmXBpjXcEkmZp
nonPUOrByMkr5ApmPBxpLFftxZRsf7mEmk5lx++9R/Tl3ansrvKzJhkJPHZr5H1sUXzIrehvfbLp
5JCjSii4TC5Rwf32RRlqcJg+xrtv3VO52hGQR0T9OKeMKyIioBiegcr5XfMqOYLN/WOWh6DzMvCc
8QAK9hq3YqaKEFAzZzzYFvRxfP7Odyfx5A2nRPDPwcCLkPtw+NeYpX07PAxdj3wQrmSte1X3lx80
YlkayJ01ZmIqVlxgMY2NhIOXjtPl/SyhYBndVfpry93bx6hcBDoNWlmPdqGPw+jeIZtyWWLKJ5IZ
CsZSM5Q/9sWYmqDpIRLKyHG65ylnZaLwujBQ7HgL2sRlZT4iIQczIfV8yaa0rvjDH0eFgtC3Tsuh
ayNZSyAMf80PK6DT+5kLDbLczHMD8+Z85SmNj/Xr52rgysKs8OZk6+f9zNoJWfn8Tc+kfD3QP2Z1
wGGO7Y4t46TRF4vuroE8I/de/FaaTvshdyNq9ifD21m7hR54tCZHiMp7x1c0m0XturCDPhohH5Yy
NbETYGY3LwMKk1yAFPhhYCXI318eHknI4xSXZUDvUaSmdyZ2311JRWrUbqXT35waE+2/fsrG/3ht
lSdtzolrxEGqFE//MTQkeL+vcl82e3jO/HOODfelymLe16g5LuVROsG0dYaxd3zVEkvJZKtsa5v8
i8BF1p46Beww4QmP7Xe3E8VdOiNBtisjwQ6fDMxYjK+yvdEm9/EGdpt5CfaBKLyzo+9T3y985VDi
OTyubUKpskYbe1FwwT9dbOnHvdKbsU4r1Acv5Fa0hgzzHnnpHkjeaesVZ0yG3bpMSOCkh/ZGjv/s
HOxLhFdknlwpBrn8J1IF0QgX9D3TQDLoCAXCpJ7gXVF/SdhP9BUfTIVkzvqTMpzxOqRcvJXUkSWP
c3N5xUtR2bKvOT2WuADbum2KKjQaoCgUtfTGrIxG/q3+ZHpJzPdHafVkN4n3RJlxYC7Fn0XU6Wus
I+r8viPh6z1J50pJvOs+cw0XY/QrMUHHpAswXF9iRXZqQvcgmUFL6zX0bIhTqidVP5LS6gu2gYiG
8uA1xLxlfnwwCzlocblZ72lXMxMSuYz0/Bnf5ggxuiQenNlnx2/ItBJowXDQZKC7LnzgM4lbLMwc
3gzKEqIiusehQHXF0HfZWJLtKolmxox422UwYKfdAaCOlP2+tcxXe87+pSHNMIi/jkMUhgFIdQEL
ON3Ck0VNUhBuJeYX+gtVVg/k5myuFEN5TlruLIXPyMxdCvNxcvxkCN4PAL9VeVnWrFpw9RNAmLBW
YUQ4XvCJxkanpb3O7N+12Um7b2E5ZHeo9vVhPY5SqbzRu6nGUh7U4PPvl7lNRwTTsMLJprQ17aVT
4XyN7PKCwtaf0RHjX9YFOeT1TejFk/U868MhqGxo9RH1YcGF8f6MbswVvjbLEmwy0KLdmusOQSz7
ReM4BeBe8pIlyrSc/QoJifxYu1UgO/byTdIEpcyS+kKPAMPiFbWeViluzW4th6c9dFPy9hBf3hXa
stkfbvzp8fvN2PGR4p1vM+vRGZOse99MFgqJDrK4Fb6T5lVBtI4iYLLEWxHeldpN6GNQYUCbxfcE
FlcuXVVfi94U6GKxqJLSyaF4ZFMlJrXMJTmBl0dUfNQcPfNjQJXjSxugMC0Mu5+dmgld3dJw82mJ
uIkOAsL+txOfFlVGhuoW1AeIfRuVN4N5fxGTrcVz6efypNu22muVOGQNjvMBaWyVJv3xGZiZ9XMF
ID9bi2oqb0P41P0MzdhE126yEonwPEcBM65Gl49M9pdIPTIjv+/Jm7FqRl1Na9oliOvLV/TfBUvA
oZ5hkY4AjQEhl1k+zkaYuU5e4TgYC0ExINDosR126cFr75hQR0q4J0iBK/Yl23GlHVw9nLmcyYoa
pM1M+KFG2ZxEWcHG+7yP3IOwFoQt9ShtV5hOZR7BcRjQfo2FgexqiwbVOv9QHateGfpmpfX+krXj
acwbFAfaHs5m173qvzs45LB1ZkNrllfG4Q6lDmiUlp2JYG33Z3ho7NEFci1MggUc3zosvLHnHC0t
z8JxxF0tCtesQEG/BB3xVS2JQstrtWnPuBZZGroCW7tL+mPWr2qgqbBFUM4tt75vdgMX0WBWp/YN
eNHTiZUtT6YY4ygPxPuNtjYXVtVheapVK4qaDMMPdaOeFaI7fdL272g6dD03PFHsKPZ93zzB7/An
qU7ns26HQTYs8cf4ctSQORTvWGQS9tEfECwH/lnC1rh+1kikRNWG6RaOL/GOTGmnLuU/eomQ/Kzj
eL8j09xGouWJu5XWXbY0o+L6wuADmEmjrrg99j8WkZ1rjyO8iGZKsoY8T2kopjgEL3/LF+wQJd9I
oZAEt+0dlePb0d5n6d8nZz9u7QJVGqhe4gCSABCsgfID5iFwsIQnyTHh/YV+dL69DoUlSzBXOBEL
o0jF1Co9VsQSbWh2a57HnqCu0vZvBzIR7FHyEB3PxkjquUHaPEXLwGnoOWRCxIJ3Sg41Klp4zT8n
GgcwPzck9YJ39/urEYcHu0MtbzxsHC1zGiE1exW9HgDxQT2l7iAqDCnKjKHFoO6WUQluX6RwMiec
PcYZ7wRJm9l19Ry/4RW7oOPP8CdUfEEIjqcV07WX6CCFk2/EMLxaMiv/LQy8D8qseCctFNVnJNQh
c72t5CG3zeSlFiR2WxSMg0Sf5gqwkebbu+4nQRxWrguV0NTdKYKX1R8G9ByShqOAUXT/vanIn3pt
fBg09Anrzj62NwlzKHyd5HtFaRIQ/4fqPDZ5Y533b9X4NHpND8/3MpHk+85y+F1igsudJH71pe3b
tG+mi1lsd23eBz5FDaH5EJx0zMLcXHnp7cxmJpnnvCMTZHzgDnRNjF10Lvyz8VnoNx/y/RgoEqiD
Wc8JwzE/S0pponcuZWlE6uE3ADp7TyrwsnPBSrqOeElEDYZ1+CU0espjT6nygUv3oUvHC2JvzvTq
IJOWpmb5ZbYo3g1DCPMCGinH2y6LowTEJhw05lXpL0vptNoPlYy7iVd6rGxazGlsnoxrBtrZKYew
Qzx+PulDIy/Ph+G/Bz9yfHbXSjgjIndEur1L0LFnVsqBhEkUjj5YD9Ck1WkEJHdPVUQuUwZjA3iv
q1//3qDrA/UfzKUdqZLPD0nRt+Cd1sBotuwwRZxPbYrer3dwkoLBf/0l2RvIOPUljl5ZDnxLApsy
DUY64dQGUVefcSVAmO7JSK6PvLhmpo8lrYa5vPbChafjvMO16PDz8SlQOz5OCn+Rv49zPnegFJGa
0Pcf2V3MJ0aVpBwjGdOwXS1SsNrp0aAvN3jZkWcC7NdMh0Mif1JT3R2mdYtQQFQc8ygVciawoupu
KXLEDW+NZ0X7at8w+9585Ht6fugeyNjHTEZfkKs2HaVZgIRrev5kW99GA986XgW8rFxdgQ1r4OfZ
NuDTcvIMJwm7pKQ++xpiOoiBRUHZgpgAzFloxPfusS34TUJiId0IrgriqlsDPKKTpGEFlvO93eQx
X7w30zLTylYxt3Ae95qA3nXlSNpeyqe3qrLy6RdWzXlMJR/BQHsnLahyf+GGC5IHbcXsOvrT2d6w
C6cIctYAPf0AHOlviwvZVyo0PkoSD/wbWWqjVTTCHwAO3FQlYcCTb1FKNmdIKsL07/LrtGmd0SiT
Sk5EcYCuDOOOttFWRQ+24o3G8WJ5aKkN8J4O152QfvrrsCK3Xge1hiA5UoNH/XpMchNT4dgNwtvK
S1pG/HBFMWuKXlaQDUf80f150bVdFQx0lnP1lflXrdpJPpxw0RoDLtq86Ak9EnPmJXGpe3DEYygd
lKH+LjvUluOXoOXrsHUZm9ptNGcaaDbm+eA/+oEqLQ81JpVCmWEYAAmQYhy5QuYrc+3TBErWhvki
ikBx7yM5JSM3xGbKFsjhHAgji6JhFHdvh30LQO6uthG82LikARSxoMa6EDRbeSl7uA3nuhyxOOUJ
ChpyKKSavcz+D2gi2XbZJB46Qa5WET0sgmS+woZRRM5Ji7dba5tIQxFbg6qZnvvTM4mIbdZu/HLt
uXgcquiDVmtjyuTf9p0TnzI2PlFflzCfKrZGjBqfZQgaRbdaQWUIQcvQpGsuNQqCur+Y7uPvhydp
DN3NJu0BsUoiTqeUi1xrySMekYR2ieKCHtmJLc1qDMIfr9MkkgkbRkOEjXSSpXnKTUwvfOxcNGRN
Eu/WrAZ0ZJ753iSUHSlnkJcSeMnLSSqhT1ka8m5kedSUnw9N66Lfd6a6+LNkCOqjWGYzTIBsSMno
D1EQX0xMBUeFjVq8Isi2CNyJ24AKJ2F0Dr/QFD5ZhOWePTqvJtgRZS4SvWCCqOo/BXWMIzQWuvqF
NwnW/7fROSwv/CYZZCxJYtmYgdOz6hRFhMDFP4DGyzL1QthK/aFv9wUdvyQzWmL2Cfa0FVsUuCoh
JJj4+sQ0xjqc5gEB21E3F1C9YDGp7UJvIVpa7ouRdVL7dZ+5xXQ5n+9TN/nEYnS8QYuMFhg6baqq
p5WBJQ9x0jn/yzQtBw68MaP9MfouyoY8YGbkNlgqy9np+NG7OP3xc5wtdIugiqh8qj0j0n76FCpA
rNt9nsTvA32/Z5pHDb1qUaJbg7+SlM8xcI/U2IZ82iN8nidRrulxBoLFDEpD0CJ4PgnFb0WwpJm+
AjNuXNJkFrcop8/sC55mciSCkivDQ8M+BKsgl1tsahNJnbFB1Le17SMn1e5Orym16x8to8BzZ98U
IgH8kE0shfOaWq0ZkrlHBQFUEbdXWvu1R2lfPifSS7lLGBuk346OFhHqIQ/LmYeoVEQz5s8c0EAd
ZhDJFmkJ2ZiWEOPrQLdsfGrid9oxwqaVKv4nHeXhQz2+CeWiia/Tq2/GQMfQ8gEQ3JloHv5PClV6
68nVe3GPBfQ2AXfEqlhoekJzhvx5409Piqn7uCOGpGeuo9zx7sLLBi+nxEHAUDEWiGTXPxE4pgPL
xJ43WzDXYtuuoaBeB7zWgf0qBlAUOd5Qc5uhAOMXgSOIHpLAFsDLnzf9HaYhZOCujNoYy48eJBue
pQMRx6rOUCcIebCFGSOWO09NeuFoZAelUVZWbXvduXWqEACACynTwn547Qv9SZ4ezDH+2W58NeK6
yTZjAmOl37AwBirxGY6MbkDCJDLnLa9SjMlvRQ+eKNw4esPx5h10Nhfjs7QVjZRK32FarbOVWFYr
GFBm+ims58OVa/7eGev2wG9eKvgy0HfY3K5juJ8fjUW0/ACqLhawbkwQh91q6yZXsDUkPeZeP+pV
F3HiD5c/EbyMYPvQagRm4QeGGQFyysVJcnt0qI4eMzIuMoyvSQIKc0iYUYzoI5p3j7q7Q0EYeWS8
e0CYxHWKo/31qzvkNFnP8Po8//kbvCrs4amA+G4PkCYMegnqWdZzMAVXCs6ovT7W9zHJOU7T1+Bm
0rVWI0fs2V+4Tt38mwH71hPNhHcqhn1aLYlzfoMwq+iusqfT0k3UXbSAT4Em0jCSqrEpWsyrWRlq
LGYudhBFhyPUtfgjUneW8tfEHkteIiZ9ZWa9tfIgrnMsm9b6I2tPDy7iB57O2tmBZHJIS/kqGxWf
dbAthflJUz7Co/jBelr6Z1aBY1dx7UpKkrd2suQpl0nvRbzkTsLCDyGFL8+J4NKneGkNMcnd4B0d
6EmoWIepaHOs1NPXbhYYn70QJnuzGFlu5FYtfC5nofOHHQhR9k/hT1gNOf+KdJxdzIeAXa9AKiUY
c/M2OEmeEgRk/oZUtA00ngdUKPvyop84lHrdnUYOvptRw8hQqPJENopELdR/pnj7ykkWWVn8YxnS
cBbF6SF4q1kWm4DLsTPKE7MEEZE2YGzXZH0iFJbInGT8RjsyeSJ05AH2gsw9CKvGXiWElx4vpKxF
Ep+2KUCz74kqIitFV1YWu/DsprCZYozY3ojFjCviHEqr3+xFFP2mQjmbL/CAbUDDFkUAJYikTMmh
QVyT+4bJSllNyf3C2xxs6CqzH2RY33bWu5V6lB10ThrZjBErovZ7f0V0PvH/wfg1IMH30vPYORfU
9tHFN2S7d/aPdUYQNx8sL1NuJbBSB6pXYJdRhpyQO4mOqr083QMzDVI158QQkY4sMkxkdi0aZKNh
rAHzgfHJbJvzuli8dWULU3XS92ARADaR/HB0QF4xSEzDFGchx3u1bYoJ0fGQx8j3vPCGMqbTaAEZ
OCAwSRXoj0osIafiOfJ8K1CIFR3hPeUUmi7isJsbAq8qYyGdFpkrcdRjSD5QwDqNZMdeIt7Mn9TK
BS/3ndwLNlWDnOD3prB2GDAKRVKU73huUYdEfX2cNishiUtvEw/XseHmQfwau2SIAcIxQ9E+9GCy
XnU+x3jPeT1I83Jjn8wNXvuZ6xKPMCy8QZPdhu1K3PBGdotBiTvpr0ivkiJyXSqEm4emqvOiYzCy
AFR8sUOjiAZ5Azaw6VaZq6wi8etCPkXgvO5XdrKxJ8rGtpzSS6PvjRvGgf315zY7n7Lsr/VprgAS
+kIcLFQopcpEg4LEphbOiEMGDHHqM/fHOxQkVtXDh6jU/G5K+yyMEvZ8ebqXF2g34VHpp36zLQl4
4dq9SZ8XHZLI4ttJnfAWb7QaLCs0utK9AfWlWkb8GRIRrxtjRiZY2xiahP10RXaubZYED49YNJMR
w9Sbnge+j7cRHkFrbjlIhgI4MFYQoM05m5lV4gopR6xVtZSpQmgcSjP9S+ySkBFOW8hjMh4rQwv4
/lUPY2MGpRTR570dI23RkbX6TAQbfWFNof5+hhjKIoq3PrfVrfnnzRMvRpJZWIf2JPZCr2r6gWwQ
6JbhKQZnvgmzWum8RJY1yOPPAWSK0bFCWkKMBpea0+SQtmJRALvzeY7k9+unD4OGSEBU/1kPgieX
zgQWZKWkXokGSn37vXqjWxHnWuEh9iycTtkUOUIYBC3Sb3bveLgRLpQ1Zdj1BfIpUkpgnh7weBhz
1BoF4Z3BnNxSZjxIywCggYYp/buoYvDh/HDAVrQ0/ZjHbNpJSOa8mxZVwdQpLvMaxYP1CgMepUIh
/13GEwMwuHqbu5PuqEFM9Aze+2j7RnhFlQw54eWBqvpp8PH1mdPNcZfW2HtkJwv0hxMi08DLWmxl
+we1XgwnSSCDVlY/xnDhDnLn+mwVrEe30jjPOKglUk8pRrhcGGerdT9Rfpl+vC1NJ/vZ9RhnnjXH
JcAUK6TNMW97v/6QitIAIb157N2ELIMt+oD4Lp/Wej8CJ++CqgVk6suPXdcFAeWwsrIuXGS3eTw4
MeA/PACCJcmeII1aoWh3QemN4/kxzxnjaEVQtgw916ka9tJR4rlG4Ke86eO+PBGxl33k6pQ4uLja
X8JWQ/Fv27O6wld8yljN1cqaje1BPPxdMTbIjWFszjdFX4drj2Isp5ieFJcUKhd354shrFpI68Xq
/Z+aX+grm1owGHH6MAhHaCLgFv4t/V4U/8/j2l9oGzCnk6Dei5e+N2kgChnk9cZJ3Dbws8S5keLt
Rnhqbgq9aolx7u6OpsKiRKHcVTKy7t3wpt71FhLCudI/f0XTVxM2P5OhU1VwdwMIX4BQVyo3RSWI
AKxydqpPPRd+lXelqr0RQq4GTycntpM8dpECTA57OGbSjmRQhPeaKCyAZV+oP6lfKZTNS+2ovlMl
Ez/+AYZDpq34BIJOS/ToIpG+w4yDCPKgOYFHTrece56f0ORW/bcjzLrYqU3zhJcP2LCpOhsrOyTt
zxl0MjfpQ/PbAdKeytOA17EhpR2ibDR0JnG6Wt3gx8Ss6tsKXfc/Ni5mheN4G+DckbAj/Le4CWLw
lUlfc4rFLGE/f0crIuw6WwtG6a6Kqauv7ATnPJEfWH321n+/UNt+RnXr+zsuoSuJrlc11Ojz/gp5
CTf3VpDwyeJxtGSIcUAZobPS71fsy2LpD0U+nZWdhtj+/wN2RLIKOH2Qkqj8CzREuFqddmvRCbkz
V4/CuBImSED/149AP6cPYYJChNdW0yF9egA7es8jqn1m9hmvoi5pmNn7xNLbadJPttgBlWmXRo0e
afhhmjfWG9WlTZuFjVEJaC/QwzcDGrCEoC9qZYwGsuiBUVCher6G9oSS1w1cbFXwHmx0QspNZUNU
isEvovP9M09vrhnn9zPDyp+jHr+d9ZXs2T71URf3Ak2/M0oITCsE2SkN6Sj4ij3AwnDlPzuAx5Pf
YFIrlDssq4ipIXtOmaAl1lFTO5xKMO2mSM0uE4E4ZzbOqD2B79OmVYe539zmjDTazdVLwj45Rjg3
u+5Ij7hks88zRPGUTNh4zM8zSQyVamCJIPoRbHX/zC2LZZ6aPxZ9giUTNjL9bSijUbojmfGRf1Fz
O5WGPXv+POyOnJSkDihqsFwYvLezgl0gBwhp7Iz2R3QhNEWGHJnDHG4pa17K97h6jqRMxeZTLmTS
QUikiP2Hpxkd+OzoQylIq7/pvraP3hy+DsokPyKAKUTAw+Y5OwQvykijGdkLKtuBTX/g3evitIfF
rA3DZ5u6PDEdowp6yO+zHZ+hmhw+k/43MuA3cgT8pfnk8xS6OqyDXvRloJ4enGN6unCb+qjRR3fu
jbA5VosgmaxywdvFLeVUQSFbGgPrlFm+95hO1i/G2ADWdvvoucSHaQ2377QK6gHOQz7635wwy7KW
gXatfNNMentf+RvuC+1OnM6RvjWaZ+jtiwd55uzvYfC51kpQRsw5N5K1da6ZALX5r7z/PebX1L1B
q8T6wdMgZsotkCtZH6czH7Bh0XJxy2VcNq6CYlXmpsFUS5b3Ka5VCtln8asfNzcFNjqQx4OBW8rZ
DeuXAQrpuJGMYjRhm+oGjGXAaiRL2zMKzTSELOaoguBOlynMu/WSuEyIFAMWvgndZhrbPBDFPPIw
tdDl9wBeMtEHOTM8oAxcrQncNKKUhR76qJNw77ktGKfXnuFBIsv5iNzQl1IH83UijiFS0f6KsMym
5pkqKKTf8xqcvXHUyX+h0asrUEBkyUE+8UHZVPmS/f5j8LrW7SQipNwVyNJM3tQwqMgFHXnZok45
7beToQBnvwCavq8zXCrbem5+pe4K3eWP7ekcvg5ZeZ0ar3cuwHnKg8i3/GHNwBa77vuU4GwoUaLA
UjPfIU4/T0Mp75Rr2Rne7ngUdyXJGR+fGosXRn9IO449gFDF1Eqdjz1Bf+oSCQ6gRrjvgkVzo5NU
zgH0hfsS048SygfkQHGL70N4wsACiasTbQomaRUpoFVVzB/OfMvzTQm/bfI7fkHclf6rbLRs6/cI
ozvAnGbGnnlMF7xul5L1H3hNYTuKf/5+hWxzCVWy3AEzvZfyfGgLE20HoWLJhtQD0FN7Ggr3lN+1
+pJxzuJtiq5KNSNaggzwmhg5ZU07gmyfHNh9aVMmhto6Z9/CePjMtArV3HsrQ7aAheAwYCy1bb+t
m2Bs65VLRYP1e0hwGKnLSquOzMRLichTdQFxwHi/jty22EqMxPfAVoVgrINGJJkounZB2IfDnB0v
7x/7hfSFr7X+DVaPn1RdhhV+gEeuJXkNCPgFnPGPiv6/rnJd/OJr4RXeFj3HP6zP3cadFHOon3jM
e+LSI8C+zCwlRu0VZJa7Rb08POgXc5QzckSok0vFbe68CfEa6ukZQo0Px2lh/lM0mfblx62BbEds
UkDGs2YLMt844Ly10qPOLNibJlozEaNo989JT73q2BRAgkJWi1lmSpRoTzMyaMO/6IGEpXHkkwY8
hV+EN2FkE3GFQBMuBFL+9kIpYaDSOZZyAVfmMbAB64sq2iNNZkXj4iKHkwKHih2JpdxXwVB1TAe/
9o959/USk19Z+wwUmcBLRuWd3q0q5whhqE+DvMsZ0wCGhpe+Mdlof+GkD27XvjgeDNfUzz4zCjcg
jlVSLAwXPacVupTOw+r2bYSry+Z9M+DOkGhbe1DcqDr/S1j04KtDDWZ6MAERc+La4N4/dzHN3tFM
LcgXVL5ObGrgimXhx7RnAHICT/LVxIN7Y3mQTwLbd48Oh17wuDr3Pao/QtNQtVHfmbjgGvRMNRUr
hqGOjW+Mpm56p9nk8sEF3u6228QUStaAArdpUSRaATvgxjOUXjgy11a+aplyXYpO0nRkhTnZ1lTp
pDQBLvBMgLZ4wbWflcI6B4GSVWIHcezF2NMSPQHKVotglz9+TyRq/oKfuBs3W0zj7F6GPYiM9rQj
b/RGYn/uwmx2HrHtGYix3JchHMaXQvmJHpowc+ysOONFN9LH2zymEaCkJI856sX5dQItltF91fJ/
ytJBLiMivd/g52Q4pdXUhvC8XSysJqqDaea+Quok4rn2zod72Uoj1pJhGKH6vreqWm5Y9ZMBsBsg
Bw6qf09qgizVfT9SylB09uKT4pyFvw69A0c9btFt3vi1YpqlmnoRdJ98dMAovMo5jD18CaJt4j2V
vDuEsNjwALyp7+LqoxhJBUpvc4g54ZIrARAKSfOlKijVPyU7UmYLVQ4+80fyAoNgBDebzaBjB99c
Mu2oqOmmixX/l2Ni3Nl3bzlnkL1PaVu7jTPMsjRLxsGbR1LeEBc31uSpN/6gR4nMJ6FhAcPE98fA
792AKQlU9DoWf6j1lFH1fYmv7pmTBhicgdFfV/xmZ+8DrcRa1F06NjOSpg6XI4N4GwsGn/fpbYC3
79IiabyrDck/YjeqXH5uCXbtgF3OegN57XPqsfgs2bLkyDZRxbRs7lOJBJijnF6OoFP7tGk3vqx6
pEd8oCUAlrdiqCyw1RcwU2trNzIf+bXu3EkVMGRS6/tTxFZ5YkUQ1OvYF61i4vAMyPMxpU66LIkX
gVmuyFR/tjsAyzmFIvMTG5fGXZRcIk/KP+Mj0Rk0vWZCE/FlGEGT6VwKnrxyFqe3dR0AV6BV+9UP
2g6j5J8Iu6QFn90p4ft5mK1RV+OlpzdBW5/3sZlOm+I1Hs7K1GKv2HN5+OYtDD7Z0V7llSjMnyjf
PRdrh89JzyBusPk58aUK7+MbGs+yIf7SCzIYPRD9wDjiV8tIAEuVXlYTL7O0fwe0WpOWsIDliA4a
JL2lt/5ZFSNYDpHgrCL6p4Sxaa7vP6rvTR27NkSmV5lA5DMHt9SEQDZG42yFzV+oTu1brQ37v1+C
82N3WKmU+HMbz+bf0gTx7uBuwBa8nn2P6FbcEO1Gd6PyfIn6WIcTF+I+JaMBwPdyToRxfH9W861x
o133USPWfTr9Gg6zocaLuYz2tBoZul8OHoGof4eqq+flTyjDtSwz2wronIbUZ3yVxHRmHLWcKqGG
cQTzaimFGm1ASPwJQEfKzT7eQ3Bjch828p9u0H0Mlx0fUfTq4+MeTsKnjbAGQbb3qPo4xMdKosZv
Bc0cot/uGZZvnWu+aw1InJA2n1n8B8TRanU8odEriH5SAn0gtXy/Q2DnkGUkweqYC2PViqEbNh7m
Sm2GSISWOI6qCew8uS76c0URSe1LxOBYReU3UFZzZn0wt36xTbkHNvWFhWRp5msiZ8LXECzSLdrn
hFHrt72VJ4VvdiBDL+GYKSwXBCPrkd+KlDEu3PsHxl7qwgJLq0xOUf9BGapA7yFVMLCiut26weSp
ZYki/6lbfB/ZJeP7z6qD774wTL7aQ6LY8/Lik5bGkekXb2S/W4MhCIsFxKUGmvqSli/gcSE6ZaHG
hPDIQZpFY4kZov7k+elsafMzJ16oM4yvmrhdLR2i8u1o5hLWax0K9YeMPoS+evMVBB+MZfodxSM7
oelYXPCshoniRDsSiCbHDaMwvOwoKBiw2V0o3eEdIpvhkeaCSFY1l5BSui0RPNebGSIVPwchyNW2
Al2RVT/UR0CENeS+04kBJ4gLFoQZCJvo7ZhEDksVBWlnvN/2j4P4YB/Q5i73J/J4VGweCPp92JJL
+0GWbrBpCbmUiV8oZFUOr8eLm8hxQDlbidBChf8MndzJegFQNq4fbmI8QTtNaowHcVN+2cjrwDQr
VOgJxzKvi/+fnablTLWNwXuDHw/T8ExKg4yjlDy6wtIDZoxBMIoxlRW/fHA0+CnOX0t44tsyhlxs
bC2rf80dk1VyOXWWBAPqWib7N1TeNEj0kmZdyrQHumZ+XCm7mvg1TPW7D40/LIi8Y96fHEOaHnjo
2J0V3wMnGHM8Trf8VY7OqFAlGwirSkbQdOachKGL5asyMytu0YUzFv4vuS2QSGC+0bqiWAUSDnnG
mO793e0pYn7A6FIMBnEXxF9L2pdbzLWPB4HF+E+I1EUZqMy8JGaDyC/9wTD4hZ6razFseb7R9j/h
Z2yawGeIvR/oCrrNDq+kk9ke3YFtxtLDP0gLZ0Rc/h7QH1oHLNpbJWTU+UBkLu4bbo/6C6FLTNtK
az93qVSR8SgddRBJscjWgi86bs7eku1YxkA9DcRopVaduvf3laR1l8293UkoTuwQjDGgu8yRMH1W
kfiD3ziu3pliq7XrDwCe5OWpA+M/ecFP0EiDzFw+vRJGCfb+CxyNC5dOuEa70ABn716F3V9/zpgL
2RyaWFYg3M9KBdWw7Z9URcX2Z42rVTA/uHFW3VRHmveua/FfKUiPjxwUWTPHuVyWSThzAAHugfGh
Z2yh/fxQzlcMVYKm8KhRjR2FRpQ4drGtk0Dv262K00KmwZuQaWpUckIRIr6Pi/qrQeKA8ibDAmhV
LoouGulVvGgHAwZjGo2So5DyTScD91nfghboh2L/nh0OXzrf3TU7IeDh3Ih5oDGFXYYJqtAkVtLH
mG4mwktJo93z7UGpp0eATxQG7+8p9xXxFsJfZiBLh94nzoM9ZK+QZMdOxojPrZXUueC76L4m47DD
LbpQ6a19K1DLLY/qK2qcLj/KD1BvvaqNmFmgKBN847F8bVGzbdNy/HgAx3eTqPjo9BTWhypK2iGb
Si3lzQmocLz3UIBBINZsYFQrUkGuCjewlksa2WEomDNOT67FUjoonAgPZ82C3kmb1gN8y7+IBvXs
SyU0IHjW0d3LQbQy5cFrpOflTa/hYNDa9JRXKd5UlF8RodHpLr4oM94JTSTiSmLBlHjoFQR2ohh4
UxDzyD+vY8cIRvFce5RwPQIi3oa+c4RSEXhpqL7cu2617wVnGHqSpjP8QvJJa3Jylh5EP4T6s7Qy
I2/30sR0cw+AV4NwKb7yYTu5I9RuU2USeuDJtIeju/uV/hZEOy/3FLYI5U3Wksjm2nh2G1GwwTdK
2wd+ms4PLXSwYS5RO1QGxS7YetiVQG7SStY839SOp1J6BNC17XFDiYGVgwRN2GPWJ+wjJoA4/dPP
XxAGqk2l8KDLSWQPklgkfwvdaRjixKwW1h4eke7RnNGRSXyoN6kibW3PZQNh5vl9J2N6Sd/tAZNT
7E6UBucZ0HRP/L/8+cdTngplt6bMoC5mhJB6hoivkTv7SbLljPt8iKHmKtrKhfCWYKC3bS+tDzRs
5M5KmJTYLBkaaEVNOeeSTNSrZXKNFbKGSzzqxH/2BEx+bsL+G6XY9S0sM5NU/F0LoE6ivC1vx41g
xbjd1tLGLhrFl9u06WHgaHoMtfyrZugeIcxlfMf7ZBWE0EUXQTJW9NTKCDRVlANfBPI92Eq4mpam
P41XTWmhZdpDHuyUQFRT8M0Rrq3tEU+KEW00pK8u8a9O0fC2yxrcioV4QHOd+n5AznBJyfdohvLn
pVPGidonO7REX4WVspVw+XtJemV0aeKoQTwPqJtHPfnm5AiyaPyjdXXsyYz/vncbvt7f4fqtMO6T
x6hnUlGunPo8M7nwMbKoHOTU+49qjWVWISoEAHdFtDNs+xnGt+N2XxxembZq4SfqlHkjuR4O8Vcn
3oNOIvoKPdCCZ9dM2kA2s7RYy4cVvNhDndKZldJe0OcPPfMoWO9lPP5D0R/XqPAPRaOQQt5NH9YK
56McFLokVzJ4EcmMqqFfbOa2CnrYh7qU4rl5Z3spaytiFpwzbKOnPDw8eNB0Rvcv6yFP3aQxEHf8
hM4qGsNglAKP6W0Ermr5mXC9c1Al5pS9emM4lhQ9tSn9gYV3XBS/gdknZr4h2cx7HxNlKtioSCHF
SkKp3BzMFOlMigPo+e0JR4gkJFmZkXUkC2SozGtldVLnm+Q5Rj/5lITpHtNMNumauLs9Hu8Ygz9u
g6C+fbdNYvVKiaqMbmHeJbGiEmtP+9ew+WmGOhYu6DOwo3z5rg1RisIdkXCdOmGyPbtDkQqDS2kr
3RwWE/3LVyuOkAqtUatuBCmsGgqxOtXlDzxEf3thQIprVELoc+W1/FGKNSKBuX7v3TpKEbnp9LiJ
58YuXdHPtkKa3nKk9cf7SeFjuj63QQhaLoATtRuQmrAa8rHALxFKZX3woEGnAOL40dIatesgLgDl
++VfOZitzLUcBaPSTWxOkFXxDQHoCpb0lm78olzEMoN/w1cY0pC95VsmDvt1jLu5z0rVldUaRknq
rCjmBVXfVQ2q0mno7epg3cw/p4AuDG608Mkl1U1RdRotdXPioaGEj8eiwAk801bt/Vydeuhfsf26
H+v2P2QLWHxyDhJV8M//5C1Hz769kQCzH5Z1cwvPzVM1bRk5ITZkiWct/zkpgs39+eJeILB7r5tW
BGWRM7ZO4VXkJvJoCeTN4+d2TXKkOlWvNYqhUJ/CqPGVrDqk15ycVPkFdZKHGVGTPt/wDHuUTxMG
zjAClO7Unb9IbeaJahe/KVXq3AQcgzwU1iByjQMAFMRNOFnMxZCHg/yUwjJpIxXB6rIRKMck4RFB
JPs5YNJnh3tZhDZr8va+iogyYZrfFt75ApWVizG/SFWvsGhGxxJ23POP8zFsOmUsk+KawjqtYhpx
Jr/cizoLJ73V5DCftJxWQ40n0BKUy7sVviqLHIChy5EIiMjMlrC8zw/d5HNe44OKl2xcatufB6rB
nWZqvInYhbqnfmaecuS6npzX75n9AzVL0byHlJaWR7C2OokcpvXRgaN/QM7zpjvMuKLWkPaaE+hh
ZddzVYqbxV8iV5TQ7wsU+iCIVoUi+rVFFXLG3rW6NZM1oUm29zWQfw8kf9l3LP19H1x2uHLXYmqe
Mey8Kuhen8KH46v5Gw6JGJUL/fjXxxI13/zsZGEI3eb/DRMRf9Id10VtMIW8UFirI4CRVZUrFkEa
eOYoNnnxkXYfCtpaivRg53rKkm2N0208HV+4kCz7OCmxJ4GHfD9MSrWlQavSj0MaaEncdKhRQYwh
SZ7UKuS1y1M8rCUJrI0Anvh3vN4R7aEb8dpuEMSdpN5EJ1r+art9UwgxYY6bmkC9Shd2Jn/8R0CU
eNRDuiVfKQK+AhZIMvV3uPo1uNx8gX+ih4rmQOE2fpZijrcQ+rN6EWvrtta6k9cJAydPAxetU+XR
7UF01WGG80ezXD8GBtDOEw/RUL1LsBxdRqzaO/+78yrpEKxqXDKEXS7jZ4aYhaJpYgs2sxNObQKC
AI5eOOkPynFRzX4N63UGqO/i47GzCzf/ZRllfPLV0PiMtuC9L3WqmRqIw1TuzpJDVzJzK6gfcH3d
WX0sKQE+/EMwvyzzigXU0p9VAvjqgx5TSkwmq+oqsr46ddNMCIVJ5c/LPXdRYAwRK/zoUBH1Xz8a
gnQgVqq6TPM33DnjmiS9w9NnfhTkj5okCYgTUyRZMZ6kUJGJptuHvU2uWfA+tbeXeRdxp0uCwPk4
47deQdiuqO2l+tiHBjTauDzoIlmyqg048nyoEunL6vjnbh8P9wRs3pGF4UB2ENmYEZlYCR351gh2
H2pxDcr6RlWyhAsEkzLD+QOMtw9DzThLCOZ5/tYFrgg5A1Ky6p9cMZAm6ju1XLPgeWWuZsoIDzGP
B1SQpSHvoP/N5PBnJx0uDE8HSDCXPAlABIXo52Xp5zk8XHunU0+FTtG0AVHA1RMKSMGgVlvS4id+
spoDWfl14TPucyNV+osOgMqX7CrG+E+GyUInmZWFTEDUOLYlvMARkSqlNwLmBIMowSL92W5ZAmJK
iWNyB3ps8zSfIJ04qDPmP8MVpwmmiING7d7PWXdA8lXxx2UcVcRnWF6BxEquot3Cd1desiR9eLU6
jSN83JHYvuqRIZiUh3a/yrJt72xqwpnVwmyIIdkTUISljbzRdy//4qBRGmwwRxmbY/7FeZ5ORS3j
OXBJQPDKl+BTKctzrojmwyw6esc3PA9mmaGiXN5q46vmUQHYdH+StJPal9SXkHBmhf3DI6xoaOAM
/wfywmV2siwjNdSyJvgERJFxqr6UirOjSYRq68qZwT1NIYCUa3QUcvUA9vitcaqNudXr+cV5UHsA
a/moTnrCyhmDIFk+1CxZUuuy7XhRw6NffzcD2b6Ni7VoJGB0m8oC7ygHbetvaIkp3pqqxTkL2L3O
OZyDnHy25N2AJXd6NsocY1kwiVEoMuRwYYnOOTKGN1KPY+Xqwc3ipWcakVvmb2gjyQNpHtFW2KqR
0azJbWCfNwvqYiOrxoDcZKC8tunBitmj32XacemN3+39dKP+wk3hBLaBWxQZC4OrvzW4B29ENokm
OKGnX5K1uE/xG4YaA0/6iRtztdvUS49d1y79Kq7gNNvUKdc3PXhSqkFKg4RZJfqT5Rvr7Sd6nZaa
uw7pMHAgJpfNizP/tGyFgsi9UFKeXQwEeWzYr3g97kKmGi59e0j4FzFyh7SBbPdycNsUaKE5eYeC
scLNVGF29ExQMQrmUeDYT3gEUoZuS7wbKw/iMepzh/DFt2mKlj7mTpRDfd43T0WXIl94tj/eqRn9
UEKEGvetm0qloq1YGjAch+KFaA3Axh5vIAV3/BTsW5bLCSzJ3H5jJQFDYTOnx6kAj/FXXqlyoaxR
AzMArDpCgzgMAGYRLLwLVS8De12eWo2OlFj6UNVVqqAKfKESmgd1a1kmtb7J5EcflJDhfZvqA3IV
HCAsgyaIkm4RHS/9Vm5+kxByiUv5MNFdrVxhxseY7ATtRrZdqF+M4CMcK/rMuWX15f3pykyKwCvT
02Kqnsvt44cMYfhTnyqVaNs+L7zUZ7TSqePKnp/w/USO3fsj2CVdo+9QiRbPUrv5MwwuuKYD8rus
teOciqXrilLa+HAhI2+qPk4mv4Jm0G3Lcjpsqz6nuLozp58BktK4y/1VMBwX6vkbOGF7XkM8S9yE
LKbz2zeJmM0c+CHti/nLAHMzSh06oPGzgF7Iyq9lIRsRGtIt78Hxq3+MaOCxy9UBVlMF1IjU48M4
g1haz7wVZZjBEiJF/LUIJ5E9rqKMkZjHOv5P62IL5R4BnwEATi4QQM+b0MHikLhciTX61LKIaEeB
BL9J1Q6PRVDoBs2Q17Ls2QIYLf4i2+bUEJQWtHG+5T8oBPa/rLHUs+4ngya/QZnhPQ1ghuOUX/7X
vGZraXZdRynPJDLCSN9IhnvmSzu06HIp0Eqmjt/H9c+mIeOH0Objn5tSI+PDGxV2yHV5VUBcBhtS
LcsFJSWfys0CbkfyjCb5bLhJHaYhqItLmE7JwJ7xUFbUIwC8fZdHVW5qkl9yMzHQeyOnaZmu5tft
jJP8pCVSJ32mkKsd3Pvo/8m/ZmuE50PCl+n/VuL2AbaT4JYnezAyQzyDGHi15Tsd5duMXvleV62s
urRITcCLedLOEIlii5uOnFLh9vuXQbUvJu6FQb1edHCd63hDengkTA1dkiQa9C3JjbWUbzwe9mHX
aUWgx0m/XJpzNppvWkfn2Vc7yiicxmC27VtHZRH0Rso/tWhyaGHjI4krscm1o7nKuJz05yiTC2gk
jpoMLwKT3pb6nCBTVuEHFLTb5bHhCprP4KFFXeyicbbzm6iqIKGgcVEi7zT6jEFKcKL6cW//TUNs
8kjIlASu+zBp5Fg/L2PrncTlTeTk1bWm4e8XvPSZ0zTBCC1M1pH/1N5M1U4tGNs36j6VL29FcaWc
COqyuYeYNnmiKx8p/jLCJVlMMOLi3FWLiayUCYl2Hqq8TGr3wnMA9NeidrO/yEkcrCtOBxWRahYT
JbTG299Y3efw4jiqzL0LL8sjhRW/ZF82UG2SQYzYG1yoHp83eWnl6YAFWUEyW4iELcYrqOBwbyft
+i36bD9o8g0q0GRl0XgRZgOGi2UyDUdFT2JCcPZVF7rUNhN4k3ZkUmpBMt5Kzn1SwW4VudlIoDhL
sUbZtv54GdBJp4e9N8dbPfXK+jpzU5Ii3QODUgucEki+mm0xGQlY6uUhRXzpcm3s9bXhlpmvS1t9
NKN7MET+Ky8rfqQLNmEOxST8hhGiUjUcyBNl4Pd2niLcYBOhYPNN1ZWKgRd/eOVy4QhI/CxrGse9
RJWRrNncENxxjIkt8lTvL1OpylDR3HH1mahpFkG/sXisQfmGpI3jfr6XWtDJa4sOml+utW+wOUIA
Y7wpEXRRtJ+u0tqvXamIuJcoRUy58Rv3EtGZ5edVHa1oBHSCx4IjBlXiwvvI09LRiiEWqjQ4lQru
fXnAI9Q7i5MaHeP8Wk3hzrbVfRS17ho0yAnyKbCD9i1ajucnEx2aK9UemrH/mXIYNxducodj3+HD
OuSlWhHuPXrAEslMhK0JegvWYUKouyae7qImn9IF2vfohxFH5MO2bm+y//8p9CGCKdNBV8C5kVBC
9EwWo7mS7/5LMhB8poa3PqNhnWnNTpEMvshYFpiwGnJLGSBezKT+okqI1R4nfZ1+4DeS/dSyynIB
iPApt1j6LguD90MS15xm/XA3Ud0o3/WcBUXcz51Kb0KODoDAwDVb0a//J3NS5eC8SYc8Be5+TMbv
E96GqkKfSvVWKeAvR+TZmv30X+UiXjNGxJ9+oPJzUQ738LxYrJgfbtg/6OwzEDNs+cRz0QdcsY05
7bqLYdvUfCm/IrdQ+naQUQ8ayPitHI6NbiQ7PWZTFHF+V3+5T2UuWXgZw2UPdlJ5+jJkUEojumnO
P0JLJqZ7F37IqQznRHzUOWmTjDCEgPaEPsG2N8aK2fipQUrM7OgChWrjjhMxfjoVPPFPvRKIeiec
wNdf8E/w0JOSlsr0J1+hwCxEEL44+HSfqKy9YJVL2DSOiVnzBbKyvMlbHaE6yABSv7xYh+Y37kEr
akvYMIw3hlm926paFBNPBA/sBn5EvrBb5359wp0HfSKrQMCDpIsWLgeUwICs7pjVzRedroMAXEbB
/NgamL8C0sJ1S3SNfLntxX2+A9XLasHV2k8En+wKXTRpzob4Um+bM+Zv3K2ylGhZtHXjP92EgtLH
TZtoadN2h/ho+sYYAsOrZPldEDXHMSFhbAY1lan4c9UambWi8jn7jh/2bDR6AbFf9T7SkiiYWtcL
3k2US1QjFC9nbrQZ77/B39GAS9GJiD4hYjsDG3QZhTESU0ZziNqo2i/ZxiBOFoHjZm1eKZa4DVNi
K/jiW8XYBS8kB2cAJR0vmX3BXjxCGNwKKOyQyvhkmP4GUSo8aLT0PiFyxlKuRGzS8P5jknFTm+2u
WdDpPQMx49/06vWkQyAqp/zGjaCGWpXvToWvtmuXVWoj3qFNI9fWhEOmRgTGd1DfUbtWw9vRETNg
/RgXHN5yZxWMSpOAU2qRQYcZNhy5dfmP/vuYlpyr2er0gR6Rx7owatazDed+1Qs8Mess6bgv5wlV
CUlSGKhO2Gupm/9r9AQ/hnqpJfGFG3zic3NKXxhXk6MBQjbQmzOFO4K+tS2/p234uO+e8ZNwOkOv
p6o+WkPL6T5sqkhLovPcwFoqDaRNxe22tg11RSnpHJMdmsqixCESr40PxqF/imTZqdtSszdzAscx
U60Vpx8exdGh44gJKk25T2XUkIg4SOw/Zgk7//kXWiEKEW11igyVC5tXIHTGGu4thV5Lfpi0f0Ri
/fMEaJv/FT0yxyCTZMcahQH/tq9vDdo6blPLDcEpLMbtZT3zEM7wSonHmKG1tGc/WB0uSeBHnt/i
En5GK6d5D1povejk33AX8wZ6wu6zs6dN10x54kN0wv51IfOJlo+/AWohyvdF42pjszuc3pPoHyQ0
ketY/+Eetjz/3GDl7WhvRa3knnQrvOX+n8BLNAqosb+WDGPWHg2DavlR/HMVU+4Anu7jIKLlRi7P
2xA9sr4Ki2ySiIdSqEP40h//wG2qKC434DxwAdIWPauRe1WiF/ygvLwvyqrcNdYtbkWI36yL9Bj4
hwlRF+hQxghwVbjhDit18PSkPRw2SxOFHTD8cQZrIHWI/rknS4uME9DI4Kqd2mo0mTCNpnRL44Vv
X3WC0EO/XJ/mWYvZULpRFK9N9rIRytnWEdC1asA0Ipmn9uVyEVjMhpsn0yKGyfPi/kzONJBG+UpP
IaYFuMa3rK7a3qOwJyoNck6QtE7UAE9cGbVI1PQoezuv1Mvx/zYbLqK26ab8/O0h2dQlbo8Mq8Me
w1P80O4rsbrmTS0ny/DHbjcZbfbPtAmoLjU63qCKOzz8Nj7W/eGhkqaIRsNlXH5ew/aFfvWpvACK
HqMwmZnLHzSRTxiXbFqY0c0xX1tq/x3mh75JFrkgycrfvpN+SA1n0oDMx29xB5emuzuxtpuSOJkg
a8y9ts69Usy1B2/ASO4RmQrOYyHC6ew3UO6E5e6SkBsLpO7WWCZp8oq8dCpxnWpTGa4FFw+27bPo
yKguWadoUSykIKhfB3G55RDb3nShL5dzVj7zY5bqu3owYVhE6Hh8FQYY/yeGC7M/HB23J5aot2ao
pjOkx1slG1ur0Hi8yvEABATZh8t2ac4ePkY7qVg7oiF3YkeqTk94uOLWAkNgPKPXVNu9jSKLAxmo
xvqX3TweWTiVcDrCdrR2a7xpAzj/YAjWM6PW1UJ1wwi7i2In9m9DDBFiE+DOdzh0aM1F9kZ1caHF
J6laMqjIOYMmBezwXuC8mm+rrbWraFlQLkhl6ImU/Qa8zX8UdE8FGGzAgFgWA3n0G+FzzTlHdQ2Z
/bXYusBXFmYmQBzpY29xpJuMnNE5RlWYKDlgHmlHSuPGGmkOWSxz6gAteCyGJVLrk5jC188YnKDS
PX0Btju3Nb1vOQemSTTvPyaBReQsreMQUOdzERzNVYcL2T4Nuf/LlLUaW7H8zGVmUGxYbeDQKBU3
g+Vrj2d6mResBBsvfAvBGocVzmgBu47MeoZ+LwPImSk42nf0xvx2ZPM0RTWBsgkesp6f4tskgJuI
MhozWWYL9KO5n16yL3zboNrC5Fja/oA3sqPecjkxGKLdFj45TtJwPwtAkSYIIJLqJTp37crITBRI
0BNTHRpksmNU6BlcIv3xYs7jRfMbg37qQ1X4JwdzSJYhHZAYquOIWr8tktMb0mrBYvKaF2huSstA
mJUE3E8Ph2z4fMLUIejrpscIy2HlLjHqW9/eC1zn4rCKVrla2ivl2rvtPZsW6KP002S3oq/k9Bc4
Sr5DZNZZMNqyfWNGkom+0miwnBuITeIMpQWgQnhbGajeH060eJyZ+M7g7GrlzddRjMFnkLGKiDRe
an3YPK02vrf44/wWmr6d0nk1DbLcKR3dFrvrC4ddPkxlP6Uc6dVEVIHcN4p9cv16LUvFPA9BzwJ8
NioQuJ24j1zZVAHBQAo6Nd/uqRVvKEm+J3J2GkLZb6z/duDN9fu7ffopLjiDaxtAmCZAk2bHxCpd
FeYOM3wP3TbYrbnu/nYdfIY5pc+9SPkkzThDe/xltdiGu3IodZvcErbMIh51ACemVh3y6vQ1mZJ4
eShXHCF5joAVhMbEqE9Y93o2SUC8xs5Za9EWl268/9cikjnQoqzmK3D+ie3+4+arw6ZjMVJ4AwrQ
xM7+EhislfLOt3d/WMg8dYEL3f5kVDE9vCjMUGnetvUYC2NchgODivn2uOid0rR7/6W8lG+umA4g
ushNHoqB+/p93UebfiYO6m2VHiEORe0SGpHyYhXV9jRnNwRwhf+tgV7y6eGNjPls5WQmsJU3wPol
x/V2HKGJKmb0BS+BI813mOJ0H3XL3e/gBxjeuQXoiWOnc6GkyG7mFSB+K5c8L2Tnr4s3xhZUfzjP
DSaAJv2VyYjJ2wtzno/8/LNPO8Hc8yvy8jTPEZB27pUtVUA6ug8klWB6Tvn/9JZLZzoyA2Y0K4Xk
5fabmXt5Jk9Hiz43WrvpNsqzT4+TlqiS0iuscjTyiSlx6bGYcmNQty/3QHYP8SsdKHr0+igeNmUX
kJExp4lCfUTLVdB8dE4aGJMlyY0/tMT5DNvlx7qAAREN+bR9/yU7stXkTQWOCE5d5SFca6m7LjX6
yJ6pSH8i791MCbMileHd8LSdYXA/gvvz0siUYWumIV4T9N53tFmsYnI/U9KV4k2JLcrnE5h1P5rU
YHha/1VLEuTNMY11O1JmTbZhzqZSFwGzyCVjpamtnixrQD7w2ZwBpcaaR+dGTvEE6Cw2Zy9NrEsC
TYW5Lf48M0xq5jocRKjTOE7NZ9J/bNK0hyzck2apM/yoi1nNn09RZlXz3QsRMYoyA43msZwTJAgV
ydBsPT5oD9FarwHsnJntyHuEPBj+dzQYUmYaRCWoLtxQZHjI0DOKMpQ/MTYjPsi+XbjxBzvV3glx
pQJcnrwCoQJLmgpfVq7uyWtb47KhTldGHVlDCPs5hAw0xoR9MjLdQWg4c37XPYcS+v6VpwInJohk
Ov+P0LwNDTeYOZFY3CDi+zTTBCkCGNM9dQNk6OqRvvTmYAadHmcp0zerh8Em525Zk23pT42UlQqv
FVl4fNO3ozMBXlXBz/IZPXt2seiJ1hJ436fVUwp/ThnTpGXXc9YHhhun70MSqtfIpQmpW9rsHiQj
NSbeM7sPWbP77y9x2NFpaiAlCmZMHJPGTKiNSp1OnIYxP+BQIOGDaXg3FBuVcKbJihQ+DKBb/jED
KeeMdGzUmVphyjcV2e9zV/NaE9v9lsGJzXh32Y7NwBqE8CEyh7vbOOW73G1McmQXZy7eoAPcQ3BL
mkZRx1+Q3pp776+0ZQBxmWiSylt9nYj/Xl7VlxVBtiLLYOEOpJ1cHj95uHDQJPO4Ho+GVFGJMnfL
KLu2MuC+hUYWbksz/wdbKVSszcpPYxwsK0gmuLf2kGQBt97BYxiRp7U3tZSZXx9WS21z7XlMoNzC
WrPITRgrY7Cndog9u90e7b+4gm2BVv7F3AnZKZwxHPIQDyi85h/6UPvn2T8J63KhQJPEOT05H2Z/
dCOZGM80qbmhV2ra8QK6dihajRpRpcxHUyN9KFwgvaJJ/oRaXfrViJwdK3fDqFguZETo41tBTTUV
HHmLkaueDt7O3UWXwrasYdjAThOjL0Q25WsjUG+oN5XP9lROS94K33/+AzTIiIPa70Bnq3ecC/hn
2LvJlwi6du4gVORTfKsrmxtc04IscfZwDkAFodNgWO0K0sKEQC6K14S8ZeE+LNFgd6+/IT7rWgTr
Wq85boZ8mLzS48Fe119qVTNe2eUqruit1c8OjNGp6gNwnqIEwx7IQdBVXcfF9vZHXIKk/BFWrg6K
oasi/B6UMlQ/QW1U0GmkOe+VJf2xMcTEHY04vzRCAS9XRnWicVicmMIn/WCkcX92KLWPgfu4J1rv
xPLGygLgG1IEPtwoxdCLQa+AEf0lTPV2IkPCnJlZpvnksjdN70v3hrQE+/EWJih7d3HfRV/8lB21
0MRUByamftyVtIRixFshHQErHeHcCjedH8FDNF3XVL1USktVPVsc4+proO1o4v/iqhSenjyq73PR
n4G/fVHviyCvMmMC8kxc1sy9drnSW773E4PpuybSdWhx13Ae0So0zzqRmMlW1gliYIUOQCwN45bt
WZmLhjFGbm59AeNVSF9FDWC/+7/k6TTGPBD7s6OMSWukgjFG1O2D63fEdC/gs5np1uNCTwVvCNH1
YhsngX3GUSthouzd3xLk48ngrRRDzCxnCi7Pet9at/eN6MPqKf9oiNb9mP77L7W+UMNPSqF3pPmD
P6OfG1ozJ2KGqHxF+nbkA7V0hMw9rfutUIZfz2im1JQabK05d083BQIChCCbj28fIOuEJ7a97v73
JkCYP5axE3VzJR3VNPs6eZZYgMJ3MgtFPfvS5D+SoACvhRPzlq1fmdm7qW7/A79torRbAa5a/RnZ
RHz8joPQwsqVVSGI+vItOCYwtku8F3BUFoaDycHvc9icFqoOnHIKwaVtHfoqn6ltH/DMW7wGpakx
1aLWdNVpSjplcNurAgp5dJ9ln4LMSi30bma+GCoj7ax1BBHZCI3Qbt56L9mmgNU5RLvW8YgpYP6N
eiuFZHB9h81fvwwUWLG+NdpJYCBJLNN+8Ys7xLkwqT4eZkkERRfvR3SOzrfOAKSDkaPI4VbJRgep
P6djnhH6XojCylEj8wkxAr9LksMtoPpFMaEgMGAqKT01CZnpAqwm4e2ooIH8wVXrvTQPJ3xXRhVW
Ne3O9YtzZR+7FhYujEi3oSmVz8UsyHn/+sRY+ecYM90vmTYaLpuh1ZXXGej6x5ww3Mi7u0zupjlU
jRTsHT+F/7Q6Bnf5MT7c/73VhPdn89ExDb4bFKzJghoHk37SEGTc+pQ71mnlsKiXolPRbyqq1yPK
oij85Ab1K4U8KGFcXZP6nlz73TzcCSNJfxR5eM1x/obgeaBp7XNG+l/MAoO5dGQzSdkeJBRRV9/R
BG3gsGWRx6MfWRB4A/wxQq3D8nEEVRl8Q0u8AJE3v93YuoUEwMV/uR87SToQjj2zl1llJF+VLlYy
9oYf0QlOLHAOeBbkiyciFPEcct8fD5zGGqmxXYIecO3rNbY6PBuy4wFJL0SUeJFShJpEah5N+WzR
KPgZMaG4rbqkMYYRpik2eROhfihfwKvQnx5S1dQ+fweGlH4jP4xu82I43e3ooKNmRHSHZbgeZXs2
WVF9Ho64yGenyA1rPSNTMq27ijRsTLQy8xXTndyrYysan2R0PGLu31cy0zn1h3kbkiy0WgnYQC8h
7Yy0IiLaBLmz1TrNB85EErSvcwfbzRkIOUU5XL8+NkfSphPLGxOTZURtbcOwtHAe1Rm5vAW0EhQ3
aBGcoWMRK6ahmmV+IyHFfhLxmmCYSfwl3jq2Fvi0tlxlltrZoTauqjdSOV5DWT++1AH5eAaaxixm
d9tjGv5tomw03MpnEiDjYmb3uTFn966b/Ble6zYH7NGuGb/62rpVPkWGlSQX21C59l/tiEP8Rz+U
KByXxUTVi+Gr3xWfsfPEZ57U0QBZR89ps8SodklSIDCm1XjyJkjih3w1UaBY5jttaQTwpU7T9oTk
J1T0a5L2TqsLyvaujS7Adg4zDBPpxAhH67VyG7qBzm1byU6wWppD09OTiWVAolycir8aY3cTl5a/
jg2RdCkJma3KhLzG2Vh4VNZ8xFRhtjkzTgGFdqu8VSliIRL5qh2Aozf9Tzi2f+OD2f/PBqfxnFoj
QyQL9rvy0k4yLpQo8jUKYmhpf2w+UGw5+sutbF3+oEEzmM+P1nev7FDErJ1iX244vEoX+wFk4er9
Um83vQLa/jy8uIrj6hPgnlG31m+RX1HOfoPJGfb46zanzxjTn5/Xzu07yaygd5/nTRZXelufncIO
iRDdBujrQGCKUej/plZdCdPWt8Oeh852lEDfqgSWQDt13O+1CAu/HtjWqHVkNRAoPqVORzrGfg5o
qqQFpIHoYJ5L+AZGCxjD/Bh3dVj6YOAZScSCNDDLa/gZg1eOIz63BAEyishkcVM5BDIIq9We7Jeo
+9qn3iedNMK/Bzo2w6WJzAZD77cvwJaj+Zo97KCyOSsGnAJxOk9x/pKSJ58ZJtBwrzNbaa3wL4KF
/mOALqZu8++fdnK/JTnHapP8LRsoiDKKCRbK2NEFm0bmq4VnFnYdF9q6JWrGtZEmy0D9jfiXNcvV
XANdQncDX+vy+eXzy/03sVmZ+rfLWn6SBG5H2SvQPXlJ0+PqyxRu7J+4XhOaofDc6wkGMwrPCRBv
aiJoygUY+H+2ayobHLQWUQone6ARAOIDQEchLYF9vKw/R6zkb3NGq8MLH7CzQ24guyuUtBQ1HJTc
QU/BF1VWX28Di0udXSBivzAdaVraVJ6dBOTTOhGDNVdp3s31VThKZHVHy1kt5ke4Ej8ljN8SGL9D
o0DU0zid2T0AZLXhECgEIdtO6EO3nn7C0BSuwrtl+OypwgkUOyAEbTXkmkd7FLpV4LbFTH0GfIdc
l/Ae3dGUiL8SE9lxOxLdxXsmT5zyR7f/Q7S8fpq9FHuKEbz9s71nQ/3O5VDI4jjO0kxUDLPM4n/V
8xJJZQEwjkaepwK2bCBZ3bnRXE3lDWHNT2FJHgpYtcZpw3+GjfM1mRYSgINfmaHuAZ7gYQe+MeyU
ruY4vUXcdWWrXcd2SpaUsVCiXfwEsFSNBMzG9n4nFJ2netAGwFRBix65S2rca6M9k0xob/GYfYIY
xS/7OrVYMe3sJy9A5ZoYGYuKcHEAQ/Tyog5MxcTgx+8879yC5BIYoDSrw6hwV1hPddLzwv22Nf7i
OykBl5I+fMVR6ShCONeOw+IPsWOQ4kNs9Mbhvy65VU1gvKGPg5XQLEDCk8UgcFQt7zkbXYJi/bk2
kNOQEIltp5p8p+rY36l/2VMPJ5jQEFPHr+EYgdMV1DhQi+464lCUZ6EzOljhXKbHJvQ96ZzadPh/
sR12yugbi+tXWgksD+giH6Z5hMYZ/t86kguot1DXuPsib/58M9o1ehbVQbV/58LElteXS0lCmzGc
T5akQv5DQFOajJ8hUHoDzMMIQam4LLlbgPc8HPyX0fy1gltnInkwpYCirfDAYd4+6LCOoZaXgnz/
u/GlhAgYeAeFi52JgTA7Y3oFSzyd24RwXcMmOGyrXFCao+34WqnpcLPu1FDVSCZhyzBqKtV1WfZC
CBvF/KBj+/PU1O8iJxK51mFto1BjZgJcS9RxiH39lq0Oe/kbAho57VpWib6sTamCuXscM6hw36tS
JImn/jL7rD160IaIUACgUmCJktB7HsDupdPWsQhi36DOUcX0Db9PAAboPZaXa2ANbW1tVclV4RhK
RlPTywqzmLunNM0zyjBIrVf1dYR6Mi3EQMc4JFi5QOryc7eQuGRsWX0KwLMlOqcHbZYsDn4gwHOf
vavOt32HUY574eq68aq1t5DlsMJmUrweEyixbk/VyaeOrnWvA+C3Bycsefawfj5L/s7zuDhx4NOI
8Ho2nVunXTVtRvyoJGnarLsv8muFXiXgoOoxRzT76twWR+pYNGbJmK4y4A+6z6s9DnimKzoetivW
RDPMQa3XSBJ/nVbPtfE8jxM/3Z4O7tnv6NfKllffZpuWGux1qHwhuuIvmx/6A27fubq4g4QCnuiL
YyHX5d/FYbpW49p4jC7+y041iDQjRPEZjywZqXy6UkcY+T/kaTEmyzAXssp7cEnIDwwje3DSvPze
9fYnyIx5uu0QeQXzKqvwmeibFZ1OAXG/L8U8NihKWxSSLgVnYB8ELf2MuJfACkdHx1xOtdmkb9nO
MN7y4N7f7eLpFPx4F0PMRzMKn/nwsjQvyzKsQ3Wit9vDI/seKvviQEh0TqZQKJsn+D86XYMoV9ei
IXFISghjMAY/SwPy6J9cWv33UbrRIm6d40eHNgixf+UK3nPQ9ypbpRY17vMaeMb/qDNhahtE6GMw
Hravig29hPh4UcpQaT0MuP9aY+zEzbkPOD1ksaOA5OWd/pvCUp8AUoDxAqUwP7ZXiMABTSMe1JJ1
GTHyDYwGQrdH1NYAPEbTtZZfFT3JiaEGf/xe6BkkkMkIJdQbLW2SvsXxrm0SZPMIyjUUZKYunQrz
vPUfO0HwLr79PvmHrjZz3eIecQRzVkbM3rVHPUUJ15j3od3r9+6s6iH3Wbxg/duP3n9RoHa+UkKz
4qR2YXsTcjEldlMTZ+fV85sUj6n2aJMbljzvHWwpobZ+S24WO4QljC75CRZRUghxQltfeliJqTwe
G0+iAOS8pB1+wxX6XC9L68KP27l42h1j2t1G83KyI4zkkN4LH9r6nVEgAQTfMbgJ4eONJuHTmhgU
CPFfPzk1iKjvSZoLUy+u+z9JUzZA3qeA0qfBtZeUfcy53NnauC33itr1krxMz1poFXtUxqQHp4F9
pUiUGDilF12fsFtVCg0AUj++KNZsDWc6kDc9H1beRuNysR7i/h3oWD2yEg3/1/jJw3GpQ+raXjEn
ZClrzTxHcwiwUR2SeObwkVC/y9LnLqg76A+jpF8Tp+cRCuHvC3cXsN3r6ObF64aFmHhvmlYPFW7j
xLh0t7GAMdhIgcLikrnkIonE+Fd+D9BVvSZMMFny5t5gncz3eCzFI4RHoZ741o1kG49HQxjgcMCj
VFZXptapVHQmASvppPgwBxzObQWS4A+CPLclYgK8JJqKdOhmdyae4l//xomqQjQr+rCI+D5grO1/
9PvvhMJ3qt6GnwosAnex3mypreMJjmTmojNwW4+PozXThtpTSOcgskepLazzhnkkVFU7Vt1xlOxy
1H54eZJb41Jint04dr9+Yc2ZhnaaDUL2kzjE5mne6ZbPKPt/5sBY3gyzkQmkby2QrI4zWHz4RQlm
rV0FyUIinMGgB1B/Nv0vcwe8OQW66qnoVGK+qPi2kS7vj73PtvqeBy/YQmXzFKyAyga/JpjP7i3E
tDrmJUP5euTIgyFjHBX+9G8gaGx6YEX0+vUqr7Pj+wfB+0qLI7xO+AoPEkH78Lj/9Pm0eVMVhvpX
bXHwzBpu09lmBy5V0D0yLHoCtOg5U588F84WZaJHFGAFv8fpTplvBNsuj2oYTgHwufFmxE0dt9dJ
NU9DyV08SF19GyQ49FVPfxUa2eMZsh4o1OmzQksP5sVRHmdMZTxEYI79deOwU+V1AdUCFOrA7P2z
JbgYDk0QbwRdDkCEQ9xJ5h43kR3UmaCgVHBpWBD19gbVEGlFmUQ9LqSyfkQ76+0gPuDsTP472c5p
ktfSrGPZn/JVuYFDFVob5HsPtpB9FMxfPnz9Rr/a3jLocthymV0R91yZz+JNbc+TiTxOzqEIeHso
XOET0F5ZTrnSQr7fkUQgI+uZ+t1qkaJGgxfJ3o4tW1yzSpEl4xTdg8+f+t6frFbRkCdxb2+gtgG7
85l82gc23OEfCZA5hypkDe95dBkgeC8qSLsUIgfLgkxO2KCzvD7fJSImbfw4qaUb70pNadbD8kUG
fco5MMJz0Ka1gHhEG2mjif3nVKoXyrsU8siwqgpgk1402xc8jL6evNNRemEMD9RZIFqlNeQwLejl
PX1z6Si9FRAdD97PIgpCMOCLcWW7Uyg8D/6+dSV4qrHQepcfDWzE3AMM7WON2vN6lwIqoL8kTWGz
oKVVhlSvEun2R5QBR+XvJn3BSQfZJ1DjIj4ydQHytwD0FbtUOZLCKlSG6nLWVLsN5nwFNJfl0axC
bf/KaiLkZ7T9ktVT4WAhnkgBR+7o+8hVYPe8drol/PhnGbyLDfpAvvUQbSmALxr1gxqRdDiP0tvV
N2byVL3Z2WriulpVZEkEbiBWeLFKmaesJ+kYEVzlvqGbfekrmBD78utiHuhricLfsh0U3O2FfqYk
p7J88ksUZKzecqNcAsL8jzJLoNpiK55FppPqAbsYoW0omFY5LtfxMm8dAJxW05/YCNN7GXks2FoI
4lQXxAtU078PrjkltiiOC0RcUUefroc1gwNr8sCV3/JILegpvEq7YAeJ7mRV9+MmCwy4AcXsX9cU
zii83kVvHmpUKH97KHD5vG73LSpa0y4VPMlqGQLdbFKODVpJztIAB31SbtCYOYo1MPUb6N3pRyH7
O1AU47z0+0lwOmZk/q/1Lpmx06I4xjF3uXkSzcbkFvikOAixIs3YOBHPxARFT0noIYGAlKBFHN5E
HD/PZYlDkt6DrI7E7pM7EsJqN2WSFPc8rwdRk/HC4x29gVXyrFRX+pXh3V84xk3i2VyjZDAvXcJc
JNcNUih18k2BHKxqWuz0HDEA7z3nI++SBfU5P0W2UjfgBPSlHWCHVqbzc0hXaqx/pV1y3jVJrswF
J+PiJcnfxDj4yCZVWEEpiyOuZ0YwN9owCihSEUWK9Rg5jnwD/zFItlhBtsqKXV1X7zMokMqSwHnt
3bG9E7F1G2k5SW0G8KyxVQmxC0hGe+1QcpGi86SAV3puQ7S/r2r6JHG/l9BGbbGpupsCiQXN5EpB
bb7dLSUIxQi1m46dRpXbmEru+w18HeZasfB6rxBdSSlPq9qKWJT7x0g1VGJReUtWXk1QAZDiO8KZ
vrLdZQR9PiaXPsY7UNnbMI95OMUiG/+5Azzu2L6r2zvXYsqExplgBK4+aPhXr6CzZdnFMpWDNYKT
2dYYYQ/CO3F/CeNH3+um7ZBBHyq6NGchc74zQN735/geKUs9mMPG0Ypbx55fxVDMjGmE/2nqP7v+
JSN5iZ1Ue/r6/klmc1v1AHYhoCFGC7ONM5UWx6InMhq2UszDUOIVD0BpAI2k0c2X/kEDQM3OUqx7
EX/MPkDd/PRHcrkEr/asBjfET26L70VpHnOQxSuqtwVluP5O7mgQro4AtLeUekrTC/foiAGP5Zfb
J0rGHUqXaGjsaLcsH+hdS8jtHqGL+/utuAfLAu6chNLxuGsUNF2sS2XZo5VVAiih33ubQ/uwn4ny
DDZKNi24mOzowWFyD/mLOXhsJl7dBxDeJL6JAPVX6heQ/7wpGpzVQycwN1U6S4rEXflEITgrvmmQ
Ynw6uU08emf0ASx8StVsHuMVaeyfV9pUFO/23/d0FsgUrwjdLLIuEnV+T0ubUBBOXjkYbDHTVGlp
AIwlggWT94lXZ6ObBjQ+A7wwciLwwhmj9e1iHWvYhh21MytKNqhE1XXMVnv1owPqPIOcUb54k9gE
Gmtry+t6mAP8kb9yr9UmaS0+rKSTYTvycMP6o0r0UQdruHPGKshWfRPqQWPfKOzndWd6Mvyxypda
G/DhxvIZHS8JCV72artu5F8Bd2yRvXNHn9DOR8DZ+xxB7dJ1vQkEbxXInpwbMTWKou+aWEHc/W+o
IJGVkeLNlhzpU27QWKY3U+HJMG7ng15NBqxG801oxRCHxo2orp8O+3y81dBlf46Yg634buOG5Zfg
UUN2KJEF428KpadVXcrFbnrkh7J3U1PaHNF3ak5oubvQL6HvK5RijHJmJYBQ2RDTJckqb9g+7ZN9
USiYCbtgvSKpTmtkxcy++uYZZrseSGIbx+d7hwqmUhmOpXJ10ZJwYG+51oMZxnUwSAJUyQFb9f+T
aDFR09JOGPzYcI7/mJg+mYNYm1hZ2/Rn6xaAdskGo7CSKSxpw/3b9rOAO4tOz5KC30awnXLXyAJF
ncq1pDULJgMxPSPxoCx34dNMEgsv/fHdq3OJW1bjXMFyM8sSLUhZok8fYdW1x66DG4Q/f/NQNm2U
ToXSt58VdarEmWb/ADOh8ZwHRhyo6dmjuyPoZQVrYKV8ZRdG6hJeHUui2WLe9riWrgHwuO0HD8AU
XmwK6bJzQZogz/oK2Fh1qLIGFk/taD9+mnU5UBOlu6n1+KQaAXsqfkT9f5V7QD6yQRVSH5Rd3LMp
6AG5Sv0ssvsUuNUExRBUSjzY612oJhq5ZdoUE+4b15qSKsmYaIBGT952j+T4MFWQUk3v79o2/WfS
AngMS3rLWVuX/ruzNdRNvu5uq+jO+UaH2bLKOoj6egkTwTIbklb4fNjYEInv/R0kgRmw0pkyXhwx
pDOg5IGZ55+ijgta8O1RE0ABWINn0VejD/HTHoFzTFIpv+hntyOkd5pnc4azjGSAPgjp82y8huCk
n1kuzRA9mI5A2G6IZIdm4/y+bhuq/jVDlIzVShtnyGz14WqvcUMf8tFiziDG6cuxYDPsrmRDRhAW
V6akFZ0Jh79vtDJCw0NVLzQTisbJKEnxI6Ni1O3eRV70EyXe8QQ/wFereBaSitvjl9rUzCCUIGpQ
Kp1c9/MQcgBeKPVp3p8pvWcR02IcaucFsPRAmeApRsapRMHKIOeKNTwXqXrPwEncJsgbSmhw/a9+
Tf6C1A47N4JgHajYC0CO/6DwE96rYb4eJ9o8CiIt0G+GWfxByMr8Bgoby0aZPrqHcudgAd8VlFf+
zOqXO5lJzebrC5SioUpw9GXAmzDhVceU8bAnwxH7CQ4mOE7HV7jelNbd+UoAwbUdFA79JEk2xJWC
ZEuCMzd2C3hdAF+7HlVaSgdiwRUOMkWHrwwYJTt/1zPx9NrRxDCY1BCq3XBhtCAaaXX+4RZQBlVL
oCBfRQzDPekQZHBZDQwBsd9RGVBNszBcFY7SW6A1JDjt1XbbYBHngGAJsxihuYYX2VLgSTj1wGl6
ayz/GeyV8g6N9Ap9vdE6yeMNves894duHixxBY3HbQ3h85fM9MHX6s9Jqgu/UOhvCzrS+SF7OHch
yMwlvZdjp2kakCkjuhIZAJpKb605pFJgOYIjhgR5jr1/a++LG1uiPPfBEVEQAL0gVc0rolnRd1nn
TLaJQiOHZiASVVUwAETyNawljh2lguw0+jECb3SS+xG2cmSzz8HqLk6YyMNNZ2afVHzUBKbMQvQK
11LCmgInCwt1THPjB7ojjM9H+LBMZ3TlzC9bRlIcIXS6hZ2MInHTJY+2mym70SImDf3enWcMgVCf
tGexju87xcJJEkKPYKEdJ7SVoyXuLM1KQtUrqA9WJDAjQUroMe2kZOnCHYxrIqJFEEvDd9ICxfXD
PwXZ+AJatMl881jdKlywVBZW6porsm2Ow8LuftWCCmN7R3/lrxTPbYlHVZAH1IBPC0o4Ufo2jLSJ
GLLqGwDnmLbBbv9wqC64LEsIXAED3uFe9lggF6z+qW19q6aisfrhU1R8+Sgvsc66Bw5WfN7lUZQ6
9xhUSrehhIAzyNMEG/holw0ymKFL+Ys1y/n4btxIUpRSDBAXlRZwiJmEg/JjSq5g3uH+54lTzqCW
zTHzkFcHbFbrmCwWNS6xu9odJ/abc8b6qhzWVHBX+IvmBtx/h2ers07cHRZr1U608sYtlvUSQtBx
QdPtRVbHzd1hII6Nk3cdgLOqhMY61t7+M8Z+xynwrMbvAKc2W8Ii9Mcjw6XUEPCAWTyLoejk2Nov
qkMY4A16nExoUw65oeHourLjftFmAAl2+Z5F4pKt4HD+Q9qZW+9CiiXynIjFi3h1tFVdd7Twmee2
Wzs9ppXVdwIwvG4F4JHYMJL5eZXbap5j++VZWMpVaXOf1dRvln4n+cwyGNBmAk9brkTKbM4FW1Y/
JX7opUhEYFU0FvEI++bB5mGHPF3KhcE4dbl8cMASSNsxWISkfZVglf2VeWvZ0W2mg0TYsxhhbmG4
1ooRWWguNT57wv98QJxLUHmnvTJc6jO1jYjAJKMHZ1LaKeCx1SxTJhisQrwDeQW88rWujqiKHZQB
PoTEn9ZoLarj2S/AeGM9jEhv0tXHbObOp0pTjDCQTjL3JOtEgRnHVG8wcbblRCXvl3JY30K+DJCR
d4mABMrRSDMWrXmNVpInrjEXfeWtpGblGqd5WouYIQXv1HJiM+kwJ5DVUmvnELsKnnr4Jq/ABKsN
YRlWmqOyi+IU+pyuFc1Fep+wTno35lzzwoa1lbg97bjXj51d7STt0Ek2IIB7Jn/eZ9TqNHcTaiMJ
c8aW1akxM7vYKHjcCi2ANnE6kDrB0WjZlYgpKx6Do4BvCQd8TdZz5OgqS3frQFeQ8vhndS5H2Ikq
tS6ZH8jk9lEOG2Hdd0Svxs1cIFByzpVzI3eV8Bdh9gDN2Y1rgPUhPQMOgJ4ofqUJx0E75A4cyUqi
ACrnV75eMWVKnAJuWAdT3ZIjGjBnL7ej0rrN+w95im3e1sWb6eholtxQPFAjrpYY2Tx/x3DV65yQ
SaDYTCY8Z1zmwo8AT9pUZebQGHKSMyDLzqmDkZykESi7rKUSjM4KIZNSCUtI7k09beFtwI07yG+4
XReVIjHlBxL7aZyQnAQNbDv6R9z5g54fyNIZzQFxk0qdMNYaRRq9guSD2f6Rl2DTn+54fSBMrKgf
BZOtTcDp+MBktFtsv7J+GbF1N2dQ9FWopZMnr6Pl6FL1HYkEc84R+49C5+B71nNVO9d8JY8qgKSH
/uMLmHtQPU1r09XcICgZNTh/a1vdRiKvmFaeYulk3gGtASQG4lTlbonvty7K1oewBGUmO8WlnlAM
I/dRuwIty1tSo8qxhuAur23fbOPhNrcDb/GkhIxi/hLkoCbqkDrHF39ORdrexuCKPbvtw/fuaFHZ
CpmIY1Igjm0IatO+M/psN1cGsmbepzuUD1GK3LvD7HlztjWUAlKfwhpCRRpUcWOKb2Zy+K8RVnu3
ANKH9SmZy1wdev+ZgRR7SaUnJ4ybAS7Y5KTVdQVJs+Uht5SibqNkuHKXwYeVM0o95aB0VFYZKOjH
4vxWV4N4iF6DcLkFovRoc1Y0SEIldbKhe+I4I8hNAwZTULWz+PcpvTsVr9ypfICHI30hL1Vq8NAR
nbDeI/MB4giS6JIKcK7H6YPx93DLHLiLeYjENQcn2Xd3teCHPICtuxybV+bWp9T6DKpnEJcQBzfn
VZbbpmmvMI3l3jB4slOJ63OgxX5O5hE2VTOxTTSv3OAM5VaoC2rTChFysTmvqUS3zL0QY2zz94ve
hvKGb1Jz+mpqcYi33RmyFYzHTK3joWZ5G1Z8ssaXR5SUuGk5tZEtyN+ajQ3oLHCgzcwy2HY8ZpuZ
ZhQJJTyrUt1tBn9mAmeQQcBb/neAvBhnbq5feUD4fLDBPCxojzbtl1V7hK8GMzqkHxFZAJLIJoww
K+lxD1wmehBumJvy984SZrdhywVTvCSNA31Eye9vIdQFKlz6Ul3LrbpdNy7qaNlgp9vpvgooy+wR
XfkCV6boVcG4jvlzmLhrjGcoPxaPS+K0U4/CLKSIAQnyb+RFGYF/n81G7LQzTLPZKNSSbAQkwBN/
iHS0GQjfk2myjpYlQ0CUFh0678B3CnAJaEZIFsAwESBS0MzKLHmhjQOR6FzXtT3OZyamfbGoUOx9
n7bZA6X/+/Nfa9llOLJxESwfqjTh6oD5A5zxx254+yS6GykGpJykxITZkJnhO4saXrvAs/GmByyK
0QRXw9MQIDL/wfzVgvfDsHctfZGuE/VMfWm/XC7Bx7ZbNNtEm7t9vc+GI3dKIJFkBLtiyDlJBOiX
zXRoU82sK3bMFXSog6evDAF7cDqMLhfKqH3dD8DvqGSohcnrXbQwPaW6UHFpEUOqueBBuEHE5Lyf
5EfeGrpVPR6PhmOSKfxqKB/DF5mHYOdqondFqkML/0zUbzytlwaREbEkYRmQRUo0H+2O8VyTFKId
3ubrS1ihR4/M6i/88OnWBret1Wf4rOBGB67XrXTDy8gwpt8AAN2domJ4MqO5eao2ZXyCmOP2JBVN
6ZRgm3UWioeBeXKec0O2/aHVHbaC+vXv6Tla21mQ62cRZLQTsPgdmJjCEyj13sE6uNlfWjzKOrPX
P8r+9PVfy5qgTDBD2lmDVMmaA7a3Y+wnFH0+n9R7EgX3yF5LkdRoTC9Rm54A63CvQ8OOU1bR6j6s
Isf6yU3Jd0c7i90GrNcx+f0sd6qX/R8rtMnKzNONY4DewlFj5UzOpkzsOCE+2gXcm1pmFIVb3vDl
f0FeeXnw63OGnRQEZZlvckf0MxxuAhPhY370r+J9MLceEpPbAXAJqK/ZA4M0Fa8rvmaN2Cp83en3
KBTG5kve6oio0EiuyL/7neHLoDWGetbIeUjmebXjcg+5AARy4m/KN3SQIJ40m6RPR5dC36G2ameG
olohhjaL9INzZkH7P/1LZJEUWVxeJsqHoQXMer7f3qD0V9UQdRpT135tDyW7pmW7Dy93Rce9Bk8Y
YDjQzzg7d7vZkorATIl8e+hmTL+qaYs3wqPwInNnLiigadDVVqsZ8Iifqoh2gsD7lvWFiism6jjn
nDGOiQKQeT+7AcWGneLjrIETVvgfsyBc3FLjIkMOy9T3QqAVvb45xfa+s1N7YGMVUUnVNl1lLS6g
YnS7pjjE2/NVjEHAl9AfdCK6Rlqe/NHiO7w/L3VDUpTWscGKmU+MWqnIQeUPY5gKDTeFRbRVqq7w
ZpWvw3o9fZlg3gp5xGuJh3bhxXY7V3m0FOi+/iqEqRigDeNUPwNIHHmfoZDVaTQtFkBIpxV4lFXL
4selYdJJtweuhW1tKClmZUKwrPY0tLaB0D2d2yCKd6hTeMtxc+AkbfmCNjIhf2EIeZCFL+bobbpw
QdrFRqDYd8byP750CVvI4NZ3YXqKAdLD2nK86akrlbk+0l6xKznTNO5jg7Xl1QVJIDNlHhvJVny5
Gfu20amwgeK4o4blZpSR8P8Q+RmPeJDQPPN3iOQv2KKJoZlCyEZPFh+1wLmWhjedAq7V9UIug8/U
T40VM0+qqMbIrVORAG0QZTrMGcWzWvOFdARtwXiKCMu5rZFbgJ8+s/JVrFqIgqA1TMNkMlrG86oq
96iyUGTwjXWDE04WM7i/s0htX9YRty0tseyyV0Twjeuo77l/nw/oiGg8aVQyNW66uS2g48qJ6YD5
yHvNMaRvy4ejOcLeNgU+PLmMMCfl4ggBVRpSeWG5y0mQT7nOXXld3m1jGxalO8jVLQu+qsDibFON
RjHTWYJD63U7cTU5xWg+N2rUPfkKrfDg5fiKRIy3Z4+ICIVWBq201ZnSXWC3migdGjHCOekUb8IA
Jc7BWtoqAnrDTQebmGvKhDtAV0qhsb9nZwGT2cTCF7KcVtc2JSN9lRjfFQr6O2RAwanBCi9RWVtJ
QwWimyCwnu3hsyDemGxYJGcW4SNoBtOUFXe0j2NBOV73W629oWgnnLpX5pwPgcdSQlxx4UtI9Gw0
ToIgkgTQH7tJiaTuAQ8JBsOYPX+ZSjr7TP9masHrLJMUixoGWXNPDmSaIixBIP/kMMOjvNNo3pKe
k1PsFMU0HIhG46Kv47USg9UHyVjvEgYNMBUNoVz8/M3PTz3Ej/a2qbzB7l9JbrcJr82VgnyIDjow
CZrF9ntAL6ZZgcLtiDZg7LkIx2YA9qGuL5BYtM4zRqrEGVXDV8MlmGvNT+G30x21d55udB39RR8A
q029KduixuK0X/cOoOzzabpQnFAlR2JWNb1OK+EelWhjsB/So3hvobmkXcmtwCE63PN+nPmQgfu0
AD6sdD/5Smnpax7/wvc8p0rNXJThfbSyLduR8Nq0BDK0o3UUgkxyZAp3xjoEWpJ8l2OQDSMR+CAj
g/yngusvqEhvNlEOUtxYYoiRIfB7mjmC6rh7nnxrmzbVNvEFC2eAWXJXVvcOYaVhUvvqXUg/K8CV
rrnOdrNttbb77lEh7385LhlM6jGr2/mwnMCK3ISlumTY2hAN8HGY+dPHzeEYr3Qz3sfWGYgkW5BD
XZkNltse4s0BBvsv+XsaXOHSvONkSNTCGc99QhWcyLMtv/cQwNzrJMUY70I2IJ0Ts+HNvtD0fZtR
jhmsBTdYOXKTkVt7VapgTqLHunhowS/pglBBkEln6edXZ3Uei7710dqm0xru69pKBNqIAalhcvCl
GAioR7WqCBBqDM6V/VMXvyFq+L4mVpmFLIkdXjQE/7zPcjG9WByVyvGEMI1W/eYlP3b3LX0PonQ0
GN7GqsyU92Mrc4xyCZUlAOfVKOzjAbadFPXX6I2lo61Cuk7pcM065yPHpeNsTzo1rg0Vd8pcUKRC
6GMjYhVfCO8V9/vhNHKiW9S30AyQkKNkK/gE9C9gOyucRJJjabu1qENCWOGIpd9eeAa/CH+wdji9
JaSxizcIiTw3lw1JLr3qj9KEmJIs85bHtBgIbDoWaQcfOfSqJCrb1cmSqKn7T+1sdMNS8cTPacjj
peDM5B0HuDGJvtt97taxaOEudn2ZuKi6aFrT24JnazfJ52RWCcvsOhr2MQd8kJyycGWEjgEEVJP9
Rfr1NyvspnGTZhWDP8UIjb7b7hjBbhckCZJunV2A2o/Jm32SqHCiAFlJrX400qWUSEfTH37nlCiK
+bZUIJcmMcU+R3m2zExDWyke6TxJ0PBtVxfouMLiCT8Vl0HbXeM/g6wcLFIyDPTAWkl+P4HmCqKX
4DT7NSOJIvSU6+ngPvoa6fpO9mCiv7HROiq7XuScw2N7oVPh2vJFArrqe5noT2/5UC5bPefehNAO
UGcLgoT7zTjz1XK08gp8AjZwDvZayuESXRhGHK/ZFmrVsTHpUQ5z2BH0LBcLkMsZuYoqQ+u/yb2t
UeXXxIduAb9wk6xpS58eNw+OEH61lsSk5ZjzWrcjuNB2SjyXhFm8s+FDmMa/B5O9JMQNQ679oyb6
A+9KjihBrrXvW4mXZwnxHuf7eELYEBZ77hV8E1IFVbKUp+/6eyGVEiOpZnfDf5MdFpD5RR0KooNw
yzd5VS4VpRFCN1xHCZBkl9vwxiA3QimGrg0o3u4M6QiLhQrkDDMV9IfmD0PQ6goglO+7uYuFxV3J
T2zXVSywOsxaNPwgN9W9tu1Rutym1n+VZ9nGIirY2yU/TI1xZbzbU8Tq9+n6In3lqlyCQDVIzS/J
k8fJ0FEnRYTtWcHw8MYrr8OOIAUJBevaBZmjVg1Ez+t9l60C+pOGNq8MNcZSO9of89EiaP1NUdmC
QI8aI+dYk4ZfNICBKJkYr20pFw6QdAvlACKbnY6BKpLSuDDC7YuuBrC6bVm1J9+uUT2RELc6UQaU
tIh8CXE1CIiS0YRM9092EqS79uO7cQ3Epw44XtHA14mS9Km4IAg9fDVDVGkWDetp+JxztdqX0vmK
+A8T4kuaX1Bzzbn9o07EC21KODLk3HZz+MUznrseWIH5OseQzTmh074ypzbxuTvfEFy3/2b7FU9h
TDBwEq16ySXx4mpoUqrsw7Hxo3X1hRPjfhz2UMk0+S0by5UgacBmO9ZkL3gT0ZHEomP5HwYJQ6Il
EwjP6eDZGQeorDBBKEise4++8Crf5/gj1vJM7jPGM37hQCl4aujA/4Jm854GjT0Zn3iUUkjah6B+
dvODYWCRKK23VTNffodoxabIRX5MwyNDIFclT8yo8nsG/dsgSQp6osaBkIMm3MFrO+lg3f/taaF5
ynEqNSvCbIXQHVPGp2NaFIlhgsIqXC59zrsp7PushUohbVLHX6l+dkjQ2XXu4KzoEPgfsEDGNzTr
pm7hNA7DLymiqRnlCYmF3JSeBdRySVBiU7wTkUlTyNLCXxvESjTCPY2xx9jqVhj1uKkKZxM1L3JB
scjPx59TBrQY+ihVwce0ww2rHTywO3Ny+fWctrAyVjgSxxx55ez+KOnioTHoduZzsDIYaf5x9Ca0
TKUm4H7WKAdiUyLOa+5hQonpd01AoFBgVjfH/Ro/2ITaDjDHW904KQ1TCsv19++R5x8iMKRbHThd
bTxoVvZrbR9z45VEbTlan9sIhe5gqQ8+UR4hMj9UcyMc6N/IjGp4/cOqLFaQrxE+Xh1qKEpSGlI1
Wq1q0sTZ6VL6GtDyxV7nhlhM6k3uPhVL8tLqwLmHtaRAVkAElVilgGmSne495nAIETsG2/G574/U
j5TiozNzBXvymaMvdx6sqWgloGTQpodp/bQFu7bQUvM/4bMolOOrtkUtojlUlbvw14ZTtM5jyueQ
dU0RcDyIsUhkMH2+GyyacQ7p3dU6cEQXoCcAhNH0W07Rr9KSHF3D2Jp8xgcl5SH4DPxgNcF1zNeU
HXOtycR95/Tx4n3fp82uB51fLd6NkmVgykkr3RSqU4BISK2wpXKzhMRiiyaPYcfgBdRwEfPg2gAh
w7aSRh6+dy7f08zLGwlhSv5n1c9ExqPaKWr3YuBzHaPpxPus8ZxLpnuAWxFxhoUWDRx466Y51sc+
dGoJ5KlCl5Gek3tKIYEqx+MuyUNzAx4BnXL0dptTVOq6NoyAeC52+xoxC697ETufQdAD/f2nj+pJ
6KwWMXXekh5fxRROeFRNVq2MDlDxf1iQ9IMbe7dpZGtV89zmeFpgjKqdz0jMlG7A1fAkhs8yYtq7
JrMyCO0l0gfvc8yVkTPuR8LLdsFzj8Hk8r36yHCXlz5UDDU9bjR7FMqwKWkSDQL5Yyx004AO8VBy
RWqT65Fm3TuiaKz+1LIbjW39v616/3Cd5G2+D63qcrMkgyoyzHBzw+60rTKDRAEBygFWWEfbDglo
LhA3i4bsingqtEdE1OIXZWk7CNm7EZTOCISsRYoXWbtLI7yhkFPAy3zXH+/q+qiGxVchdeerm1bI
LjbRB9Te4T1oRqrDzyekNXjI++npnzz3VBhP2oOBnryS5V9WmSwXLSz+7s0HucWBu/TF+bHgxgqt
EOgGSxjyUFbEo4h7ojvZX+9qlKSFvDmottgIqhnSMa6DifwbPn9lNjiG62z17MMTgUMO9YNC9MsA
e4bacYUik9Op33Q8vVD5RuLdi8M7IiQQt6F0j1js0oDnPJ+c6p8GWcnM46JjtjAHM41HiDiT7JAw
ZlJM2sZ0+iN/mqD7D94+JkFVdYuailfS4H1BhtPywumJiq+CVu8uOj8XjhbUFWMfjUh1iHUw6VYE
cAO46QsAQv4NrbzJLK4o7FCfhzRXE3uY03b+u12qmYvVYvqJColoJdr60EeQKRRK1hEF5F9SDjes
hnbKlniBI9MgVWU0/sZj5tLv/kQnYnRmyRvBydPOy0kncHOSc/xybrZapjl14K4iVCMtVPWXZZTR
i80E9j0FCYRmcuF4po/aqJ9F8kD+ENXmfu+WKYIZiqzQqQI5VrUlB7E6IOK3BMDckOVCnhsTjHvj
wkgw+js2NKg3X0GJeUMuee3s+SmdoVZir2r3WAD4XEKAPNdK1K+2AxyUssXT8dA0jhDTzlbSG77q
rBVBkRG+oV8bHvgsuSt7KJ6rqas+I6/qusonUTvtHqRtRictc+UVMd9ZlbCpuWHQnSFIdF84MI75
poLtqPunN6IKP+2cEhhKiUvFQJ6xGQOh2hWXEkoO1BdMP9XoG02D5LOFxKYYXxdM10BLIT3PflAw
vBdB6l7HDsR+MhRxsQWrGj430tN/DfKwr2RVgh92kC14gDv0ruG2mFVAMxCFcCtYqEg4bsQJJYR4
Wl4nR303dCyxmotCHamKLAf8Jx5e/xHRgaBTSDU0T330Ov9IYUPR2Lk8+SZeS0VDVcvKvIcLK5jT
lkTE22KhDWchluQm8sj7CLfMaNYRpkMYVhmf+ntYOHUmowOgBsZuxNZXXnLeynMvn6zGbIfVUZE/
1PDy4+cAuyQXzJQJ/0a6425Av9pH8iNqqw1z+8eBBkwwpNhz8u0dELjlxzWd/lKjF1H4bG4B43Nk
ryCvBNgvY6u8xYnQRcCBak+/R6dajYeBP2SB2ExzQcZ6EI8gA+OsAaFHT8xl2mw3O1Xt6HETmRQh
/kTSlOZna54P3D7M6JlGIGlp92+cTAvMRffScnw6thl7cDKTuig1mwJdhXEktzjegqbJOGrldh/a
8ga4SX8UAwxSgP2l5Lsxq2GsKYcxSBif2sANZgM2DXBEc4/y17OwF6jd3M4U/BFyKkjOoQpBQBCW
L1s4z6jn1Do6eW8dXaaou26Gr5sLoUXLvzDVEQoeujUQ+xWpmqKRlgy1Gk5H7P9x6JceL9z9Roze
79jkQ0sc29xtG5QBVKEFBCnvNuzLVSVwSk8V4+ehhjygwVEdUsWt7o7LRaH3VqHaZPXywuLlx8ku
jogdbZUjPBld/UARAgiR+VS4FuaylMvNVN5wwJUnIeVIWio/WAOzN/S2gJcJCEC8rhM2a6to0ZTI
xM4zamdx84fz7eLl2j7sQ1H192bwLYwi2xNRhgfMCacV3IrprJ0eIePbcqyYQzrXALR3K1WQmCQc
QT4LZDadBL/VOP5NNXiO+/c/N4g6FCDAZdH+Rf0zrzpjKR2pYw2jcydxB+MEFfE+hQ4kcje+i3pE
snukVjJpfQDOpXobW97tE/KvIPxaS6rhfvw4zsBTKk5SNx2lWviWnqKEkso5SLK898pcVxgEFFAs
igEvO1QXxk5YzCqD6YA+f1eYv7y+w11F7eNcsgYYAxz7/tI0H3i8bqsFH4iGBW5jzvxx2k3U42GE
ZjZdFwqeWBljygjp7fdta+jj+stWQjHR1OzcV+BjjUJjOSWxYKa4l7vw6XKWiLFRFKaQ5GTbemhf
GHJrZKEtQpMVla5fYHHkh7hQprJICRmWWKDS1tbHhX5nUD+jnFkbaEdicxzUIlTCTeBOzuTDG2O3
76ojiULhzVDLFoHHoYvdwNGleGh3HFuKrGT1oVI39pRvIYReDLUeI/ClPI2bPKNcr1Nczxehn8To
mvFNTbFa0dre0kvmBB8EDWdkcitmR6o6yxT6NtxQmpdcg4r5M2wGSUR0JhHTIS6FSDOozyZvywS0
pSBmZMcR6Nti7ci3M/sn7fkdKJ1n+VF1kWN5knSzzocCszzIoL4skeAzZiv5TylkItv8naFsItHm
dSnlG5KiJdBNFoPclaGpm1C52DGLcEoDd50IJysALTbKFTVVQqxV7zNQHAwgeYjVW4dBJhGbqdFG
OeuPGFR19WrRhW2bh9sT9iYXqTqnmTUSbxH52cIYiTWa7xyU2LAO+lAz4dulgwM0VLaK0HAzHcYV
clz4msLN3vq1UL/BSVw0cYJZAgCYwVBpodfKIyiAAO4LmtNSKI6ej8sKVxX9mtI1TBHRycohOOk0
U+INFDCFsOlxynvSKpBDG4yq+e+A8nuQgJ68Y7xvHqpEpsXYv++GPBaMySEmYDZq3RZX9P/Kp15x
janMOBZZDAFzleicVRa2B8IjizdcFAWPuNbitc6jf9afIlYIf3SXCqXGHalPFdRffmq6yxO9xywf
GchUxr/S1n0hUILgLE5ZfBeJI3Ab3rjWLWXi65MkZTaxA/3Sfv7uZ5/t8mseBUp5ueNtQvzKQZFb
kzwXwRSqeCAHYX8e2eO64EiJtoZxi54rNo08bgSaXEVvkDpoEdhQ/b+mJJVCp5Dfa8GppVPCJ31f
xChp8CZK8v1GQWHv4UDVWD+ErMAqGjU8mw17qbSS8osE5eO9TtvcmhDa20F5qLqkpZiZaWR4JAUd
Jjiml7VeFFy9LxDnZBhvvheHUPqKESk3tngzFwAR91iNu/Jr7YLIeaL98e+fLDMhDfKcfvTaDgRU
ddJnSioacbpkmC58IKEnTNn3ufMhw00XiNw56pPn1E2/LWxVSPokhUAGxUkv00iNUaiqJshdzNlR
YPjhSkqTcpjdvKxrW677pygiteNXbmtIX/b2RdCnM74pAOolEHN2PZxKqvbqj/ZVjFVOEVcZhVYP
dU+JzSxtsBiB683gK9BYqNfLwNxX9GinxgKVvcwqT0lf2bZCrdV/AhE7h/81ADRpESgfUq3oY/mb
eIBCRpC+C2PQwhrQuZOH3DWijU+QNaGvWIA5Yo+tDf/64bhHMu8t0ymHmWfiLBV8fJ42HKtPoaRD
LdjNiHI+fSSKK3FUDg2dFhQ+kOQUXBpYGf76y3froIKqjWzkSzwczMwTIrdXM1PB76OQs7/XdIw/
IOjXpDowPtNn/XXe7j+OzeYo7OOAxhxZKvzkt2s7III4aBUWJCvi2FDTktQMEBbPu4cFCOa1NlsT
oOguSIQ6yv1d49X7vf8OoRZukEDCDzo8k31eGToPg05RKD7DlW46DSFi5BwrYSzBwN/SfdggumFZ
bgTlrmnqosWsg3D4FAGB6IsODRAdTvhpzYjbiR0gS9AqEpNA24ScNRoyEbOjSmD9OV1a1Lkd4viE
SeRsibtX0WPpLBo2C9vHVRzSYgV5OBX9BvsKX4nc5c2Wi2xZMZd4gnZliSf3ngDE0gM4qGGJsrPt
aLuG7ukgipF5tioX7vLWEejr8eSlMVcwroo1fkBCpJp0aXZnXPT+ayeWlAjvNxuAREbqd9KOoMbI
6J5P/FpFbMFWgFwwYGcQpmG7IKx7mCHFRw56I4QA04j4l8yWzKixNK0JPnhuA76JtT6IeYAdEh8X
cADqKKRgdfJsi5irO7c8iaLGtC8ICvPM3QaWn43qHrwIU4jm3vHq/MqYvOBPnyVNiiX4fHRnCrho
XctVS3Xzc6qQ+iziGsFjGUuVk7EbtayDj8nKbRF2uQ5TqUi2RPuTyVJOuWWuClpaI5JLGL8x+EzI
w085BNphS93x+p4kGAGcRrMLNYgLHN03sx9H4mpuM/eNIdapQ/7rw8hjFISPRo5tuZRdPjRhr6VE
LkO9JWV2g18mWgQLnuHzlamF5W1KpaPLW6s9yNMhc3bVtYQ76rlMqX8QYg4GCld4wkPnHQcdHchg
/JdAmfNvU7kYJYq3F4Z7dhdsv/lSTlXqSSRaXvVAywFeZoJU3lSiE9z4IkA4YKr4+rLmcB3YyybR
qNKEV9HrYADs+ElE0aM6vZXI5xZTvd3XOShG9jPdQqF+9mippYhXeiUl9fW2IItC7cP/gIWzKfdn
PLZbwG3GX/KznrmN5SY+/Fwfvre7Sv8hNnJW4IqYMvRoqwv5n+uPCfEUkyE9JKLWb5TGbbFAPrSt
pxYdVx3ziJe8hX3Nz3Nnh/ONOywts4owiB69aY/d9dFnfMf55qa0rn5S5kWwP9Y+pGY/LTOSpoB2
uzNmdnu0C+hDf6nopgEndU6aiC5lpoYdrAZy+zMkdYSA0SF9SfPcl0Lch8ge/5rUE8gWMH0piwrm
NDhRsyxBbUyxRih4iEPmdkmRU6TlOfXFes2N3OhEZcmYshbbNOGRtdx2r8fY4TF9l+ZStTBLWuEz
fGvn37EK3woldDTzl62WobW8oCxkeDm+Z8vaNNEYaf1fJl8Qsr8XBiU3Br/Hv5AjFD6tibPTuLHI
t5AFfQEGk+BcsXy6J1MZR0ykVFT65gLNm8pngcuLDZpY9da43vSkf8TAJ/RgXxHiCGL8MYMDF+iA
55FloFZv8AgBQr7khJExOPh9RR1GgAfFTyCF3VLv+6dFGeXISC5DlKkn73m30E/YqbbILz1pj5EW
ohvg/dzh92Eb8FQECHnEW0FaD0EdDz95lS446J5qY2w18hfPxsyRJ57YegFEhjBCBhUogcfkAUGh
WPLgbcN03s+eEXN2C7yG8xD3tPWDEUv7w9hAUwwrz4xnwNMsj5lNlTRsZuVgNOyikyXXC6stOEAN
p0KMldxMvdnwNb97f5/5sIVYMVuMFAMaaqqox87W5Ep3F23prypdbghiffZyLQXcbinwhIgbG0yA
vqT8SrPSzIzo4hKI13tzNVL1vLCxxPxnPuc8TYElI2K3N95k4SyWJ3UYCQ3wGA+DuUXNzenJYfFO
40f98EXCbwsZ8cPT53NVLZ+v+kiFGzSVuglSz/r/RWRka3Z2lF/x8I4Uun+q77/vWoQJ0TGja9SR
PWmwfJffJDLD06MFfdsP7wXsU2MsJDHmJMOxHDbPfZJPnlgfzw55y2Qk4vuJlAtCmfT4//DQtLNi
zkbUu6UAeW/v/XVUVs1Ktt7ROhuN7k2s/SF9H9Bqa/v347lW7EfgRg+kHdA7Ai8ARoKv/ZO4go8W
iIhzCCahW6oacakcRyx4ULcKZFNbOzdlTnE2uoinXBH5pPwVRvK3oBW3zPtsM6T16Swv0/IdK9Iu
YT2tX+fxAXb+ucSy1Ec8le105DZl4nyLKxG5nVmDiN0G1+qBDYRVikum7x918RadJWU6CAzc28lf
A4+/Rs80OjR+u67nvxVfqcG9mckTjCXD0noGCkKXnLpUs6GzJwXFet5IdPP2ciwjiBWYfNq+lvh8
VIYuYhvR7wAHywEF/8Ay731Y67ECdV4s4lqeNoGLe3aiuDtqJEMru8w4CQwfkzIi/NsUmOD4suOQ
gpJrGKnb9xrJakS9sxN43G2YJG6r0DLCdq2gmdiZNG6qBaHQZXCP6tvE6lxqyH43r318Gc7GIPy1
oHDU6HuWCkaGevKYksrv8P2AtBESJzJxLAC9lLAeeumqh2v7YlqfenGieN4ae2Xm8dWtVq49wXK0
tEyBxghoKfLTlwfr9QviY+wJRq+p7jzb6sJ/sPmeMl8X5q2urgbf1wlLiDgs1UHM4Pxoj55AoGwG
Jgb7Zq7FYNO4+39d1bOH0nFkhXXKKh9Gs1TYgt2tGv9PujzW4veAC6qU4Oijh6V/oPBo4J0+uM1y
qzVyfyAhWctC7gTYQWbVBhyHefEHa6nKcmAj/iKIc0e1ZYqzmMu6+GtpJbsVcjRyHjF9h5xILY1n
t5bsaVCiPXcpidzy/D7inTPdz/6LuALOg66CmVCYrLenE1xtIFLmWluLQId9z3gEopCt229dufoI
LuiYzo8LPe61FO4QOlptUMncJvlJLWTQce38d49s7sbZI/Wuj9bidBZOqrbkFNc5ndK8Y1/ThLiI
3PWbw/bOmduRDIqSTNd6jjo9VVOsMnALOL32nmvVY1D+4xOQcvo1wkHiAZXsVo3qIjW4uVvgyPTC
N+PfAXo6G5KzihqDi7GrW81aiS3Jh+sA+mmYGz8NBhBrp+1IluTaaa87jxRhOwUqwvhQ0C7Ri+gx
mTvPYS980wVHny+HZLTX9UHDqJuPaXplq+BSwi4VkzAfljR1J/R4te1Dtp1uuXIV12l9F+G+opt7
/iQ6OalbRVEKYnV2ndvufRBpbJpV8JY/J3BhJFzb5RmeAtvWDwVImVJD+GX1XMfyZw/0FmHkSTTi
a8M32x4WcMynags8ifompOzpBZEQtOr74Gw0sK119K4TRiWgzvyL6Dg+Kv2uuAWuT0m4hMu6gANJ
eFlPxykgrDib0nAJwgTnlpDy90fnjjTvSzXgS3FPmiwDoaxsU+Vftqa42XejO+pBwL97P7iHssZT
F17tVuSvYZpOmwg/wUiSQ1QH9TZwWDtAfouXOt3MczoK9gqb/UB525Meu/wz0D0Uji5FTTfiwjwx
iQbm9BImKJi3qAzNrigoqq/70BXFFP25h/27ssNH4K6fX4Lt8FYyjArVWj0QPYn9jLgjoN58u8K6
ndHVVyXQ99lEV3haLZVw0Qg60w0x0FjLEdxJXbPWveCEajrq45OMJJO4kgtMkY8F5MGjbUWaaD+S
pDBhXGFEDklXpfAZTJVGVe4W0lzUoEZHQNHVmjbwNdg+e1Sw7YnrSbRVsczNLYEsI+ie0PCiHqu8
TK6vv58yX6hx1qfac14u6E8BNBtMRxKtb97V0aGeMMLmc6rVTDErz0nRPgMK2kuo583sEbhuADJ9
f8j2b0JkGytfcFBZRwS3LDdJT7LlfqvK7+9E61eRAfOFuu2+zpeD32L9gaS87co8hS1bWn8HDS1S
FF6+8rqYYCffMiWd3IAc0vvlKop9te+40psyIIB6eElvCvMKuFSH6a5LD+0xmmWABJ6tavD/+OE5
bkza+e4A93SljeLFR1CN3i/uu5xpOS/m+IDq7JyxVZEHbmrvKZKoYhMbaZEcvrclV01GdOgd23qy
nhC1jIssMcJ7ZlsO0DxSVpxo/nR1W5yzJ0/aUVI7+yklAWi5sqArMiCdEvehw+mxfjnjGy8NleQA
mHPtSrv6tTKXYeBUCjburUhgMGoNJQRh6rMktvbiiS5eE0KfPxU9QEI3xtM76t1ooBV8UyDO79Lu
kevwMi08bTDe21GTS9fwgux8fLL2QGyeIQjBIvFjX9Cl5k7UZruP0k+LvuMVNp8WUXlQo+yHxQQC
ZnBPUSpMGb2NIUuK/NyDbXQpX87BP3gL/y63QxeMOOKDngMxsuxFga3kijAHbqy14rKaAJnDGbUo
O1pzOx8e0Vh4UNQdwZbMR0kAed+Rd2u4tNgy/+bD940cyoYlOk6MNNDqF8uQiqx4ubBg6sgUuomK
xSYjhDJ+FmdJ4Wrarhx+EVYNwmOfT4MtOb4zFpA8mwb5ddymipj+nHHW/J0YJHEcYC7QdNmjkayt
TnNu78QDYjKFYnUJlU0Od7ZsVt3LDcTT2cxVwSu8jCt5wKLqFRg98/RnVzUSbq25xyTX/5xelflj
59gxj496Gj5ucQm/fJXynMOff5zXe+R3lwbLOqRrM54q3U6Zu1SWVTxmHs9IDhg9ombPcRnydKW3
e1UZRUJ2/2O6MCRgQApnUaSTWUYrPaRO8sbvoWAwsd/kz5mDqZdCVzIOtoSmRyf7sO+/jCCv0fQj
RxqPAqjBIxc3MaA5vUPyaeyZ6R8BeQSw2cBKOBmvnEs6zPMaGgqsvn07GmQzLqEp2WonDLYM12U9
rXlraxFqUFFFOSUwVPfB1+MWfvw1AtfqnOaNbdeK26zmhTD41GDZrRGd984rh6QKyoUZWPb+Rck8
m8iiNNrYTN42+DR/AOOSAwkJ3GKQzpS3dJ0PuGDGAwiLybJ1MucFIlGPksUvYIFwX2uVwXysMbUk
sG8jZf+/I7Xe4XUOr7tQ6uq4HoshU1t6eAx0eXiXbloxLM5VEKRg7THwdkgx7l2qr7kjkazOvOoq
10be2fh1uKkw2YPXQqAnPFoOIYgUTOHw5VU2YvchknWBM698+0urVVvmvpwNonqQL7ubD3LERR7q
G/c3YugGEYWYkL+i0TsLSP+Y7Al5SRhRTeF5pGSACglQk2hDTVtaoIrAl5ghRISumADzQHtCt9Ex
w7TRt6dlqBu3EJgkh3nu+pNhRtr4eQgkosEb2i5Jn4dwLYoXOyBlsXuf0Ry1QwXlSKKAPuciopMu
RkPmNqV9jdF3C+dHUdDZffIvliMsuEhDA2dX6A3UuhFgJLI6fLd7Dr1J2K6Sf9VVXxCVBgSSTOco
GRjAy8jZnVnoaE1+1g7SgOJINLVDsWb04Q+vTjBGsj9w+ZcZzzlb0NpvO2ihX22r/krelT/LjWTH
6WkOGa/4MtrmCgokR5dLRrxI9VU96otySgMHnqqnSEJY7QGtk/OF0yNnVMUrg1PLdYQjMy7y7h9p
b1JgcIM6bImt0UgOpN0smu6do2kM0AbRBZGkGLJpPPinC4LeGuhcTZKqAIcJPBTN7xF6Lqahx92J
lA3jYLHTX6HGl8+ypBW8+jrAjgtdWu0RwgbIszCEzm0pdHGwwXXAl1YP8B8j0dcpc5IslDOjaQDl
ID/Q9clmZUzahARjEmHRcax5EGkTY0N4swAotpV5TFF2Is+AaGKzC9qneiRO+JBkY5ZC2v8a5BOn
Y6pDEpbNTH2Ax4K8e8MJeuDlwkTShdxcAsx+JiB+qcJsBdjYjp8T5JLHA04CnfAr8mqzbuy3vxIt
/eJQgq1H190Wc27HFZR1Vn0lN6x3GllQkclhUJNTtrv46jEK2WT6HIR9GT7oajJSdZZ1L4pnTAS9
7PG7I35yy8V/+NAQ26XVO3lPAhjOWRd7vMMdUlEzMr+Jw/X2VJCcj65w6rNUo0KfsPGcAoloGYGa
9prhZMOfW2FVcx8pj9YXl5iFWmTW9FAcDHJ1cDg2+CSvOJjJ1E/gpKEvbMBbj1hJPXH9HqMGWFbB
XfJj5Lt8xF5y2Ayvj7sGBJRtFxdEZvDu9SBh2JL3+cpfW3PzBc6y5X+7OK9wMYtfV3NDu5n3tYDQ
5fMz5DhrOuIlyZVTnJWd17mfYQJ4nT+FYpxopUuffdbzIOPam3PDrFKS9iOOx7tRcyFVkKtpfBC4
g6oLGP0Er4C923v/h1Rfb6wEqfHGgkqLahdww32SWE5SCMiNXxvLNB2S2H71fGq+oWhqZTalprn8
QOQ9eIXefUUxq+YjVRqIeXRWJpBDrLMlNtVEu6r0KLpI0z29MZvPcD33csydhYscPbO+yNUM8B5W
GI6bqTHNdjWBKa2Afn7EzT+RzxqiYcN+Fwo2ojmeqc8niKGeZ8ZxEy9BUZz+YHMiYYVry25PzA59
jgI2sYCMPKRKYuendJoxyCQrv7+lcoMDO9w2q9gkuMRupaR7jaOTXJuxmPrO4eV7yOGfIT78rldJ
f0gd6iiSRKoFjbw794HEbaCv5jAS0nVyRAUwrAk5O6iQLMn1spEfBw2V6BB22mk+CjVyWEKtVre7
WI7EnO6KdwTSiKoVyK4A4i7zLoEFBn6rneCx/verpftdwPYS2fZYyEJ9iLqyotOXdANovF/cRWPi
AqoTor+GR53xvw8R20RSa6slAnu3Iy2xLQUIMBu4NaHFjX0tmBgJU9/1FcvGAxJOjEOjoMHrgD1n
JUNiPsB6WEL8wyzpQlcN+RzEMnhQQE4borUkD6WLoWh7LkoGr30MX5irelshil4FdP7aJYJDI1JP
Ii+9seXBFrVNYOPuiJ2PM2BRiGAQsNu26KQs7LTz8pJ5eixS2VVEiA56jf0/lRoepeLHt0BeFWgc
GiiH5ZnfkWvEXb8tvB0TsXIPC+gDws8kKPTE9KDQgsOp9YHLHADFr7lRevSqy67EhZ9d3LHuhY3U
ZgUZhjadUo/XBVCnXdT+ZN99EBb9+fyU9bYIsw3TWuyisFje6gOw/8swxcc4YZmPndHAO7GlArTX
XaQAFTwQqO+9b1vQgdGPjTX9g0TYbutUlyAjEBSeR52TMGGHYht3bIMuKradFEcKptEitUEcnPQD
eUQRGPfebkx9fQxcHnILYeOUCkKVCNXPIaWVib1fynKFPXAOz8gQNfiwv9fwgRbVreLTTyCqE+OW
pBXmHOsXtw4hD42LfUSZZCCZwQJhRNAcl82y/QV7AxZrtuMfvRHFhAiABU06KO9ZvqEbBcSGVWVS
tJ6RvNdxqJAlbZxe2DINFS/Ho0csYRu2QtePmF2/Ql/VOo4AI+syfJinZKf9hx9uaB8N7c1U2NSO
sHqgI5BLiBsjDVI95NllFMjjE61epns1vsf18Bog86EJtF27dfdBs1Z2oVIi2eextrl5A6n4EA9o
ChNyGLG06NvtDgiBjNMRRanMFX1ta5xKEFZEGrqylPeneqPTQYShPfPVnPJuhWMi7ZToV5aOEqNU
QoGMEoxtfhqg+ruSZ3wQrPA5O5oq7oM6oKD85k0GyVRKV49OvOzdDCUKWYQ/Dsq+McH+hby7so0h
Uu6KsLRDodba55qON53zy/WvVhb6EFO0eY5oHuQTQH4XntT5oGdKaTW26Q17EiReibNfRdVSLDSA
Kcn7DaUEas2aj6GJaKsv0eT7V9uNvV1dvUC2A1YJbG87jIgm98PTq2+iep6Z1ukqFuREvGwOsA/F
JeGqCJjZuB2hOjuwTpF5vrImSIPhtT9pK+UR6uAX+rZEH/XiaNjc2wPI5cFmiTR+iuUjHjjY0zHH
wTn3m1koIR0vydIirgphCuzakqdkR1DyAd7fXeFRmoeCA2vdRa9b2DQyPLeCkIZyHkQpU0WcfH4H
eAuikmMnkj6lkXseGF4Kh8f+AAKyMmjci8/1Ts6AuqtryvAU2sXHuSlb3cXKR0NMIN7bS+Fml1MF
hVga8Q9OhZ89QVpp/fkdpYj5BVgs41OHCspcNEl3sgSwrzYQXKNBndZGmJsDX48F3Wznba9Py/gu
NrdlLrs5cLvp3cBwwZe5wCT/fLtNVZXjKwdhF6BKGW3BcWcBvDzGIJKrBS2bSQ+N3FzJpKjvdTEk
y2Dn2v1OK+t76lqsKegWbXDPn+OYCZ8lIIun4J/gVd54w0gMcGvdeWdUK0XAMeRr3AS+bdYfoRtr
+G1YRh99QLogu0RHGyAv40rJ3JmeOXNALNvs8MtKEU8j7OhjpDzPEDuxYhTU6whgxISoJq0M3lPb
gKsklI01oix19M/VuQYkzucuIJh8HeXOxKSHG6x2skiEWfRMnbFGZKF/TGENqpdha7z3RA2SFNQ9
HSP7nOB3GbMyEQF7IaTy7Scl1Xp1rV/sfRWNUO42HsQJtSn5IZ6vJwlAHL4uKBITu+zBEO5B0/qp
GxHQAiIIsBoojiEgBJZ88Fag5BEFav0+civ3tDu7DNbQAQk8SVitbp9+skHVnqrEPAAlRuJxC8lJ
0ri5zgwphaTn1fGA0CSrSlkzIBqFBeYZE9USDDSg4gaaBwx8J0Vks2o9Ztc542QVrxk2h9kKRVtx
3xaTWA7rgnyE3XRQLk7VkoXIhiJBqdGhQwq0DTWEQQW21UY6LAvnIXqezCXjkEHk7ypf1/+HW/fp
3wIgKR33l4eyPyhl1va0cEwQTxxgXAQHESLIXhVzC/0MVtpyaRL+Ki/RHQkqOR7GNb+5788yz4Y8
kUEarx5xdJLwecqy9hTcGWZ/JEuDR0oGkIhaipKkLLhWsQtS03W00GfI5B+e6buF9m+vaKQQ2sVJ
sl0Q50bWysSB6+X1aZW2pB25DayLmIZK6wDXlIi0wjCPq2MHbarmwtizuzwS5Y1EcZAssKWo/rdN
WFcXLBP8q3D3X63uCUVqhfnfMCbx1mosz2+r9ZHXie45wsdIv2SWrAXwbU8xpUxl6IDmryM6U+AI
uLNRl5AH6N7w5smwH57Z9leZG6sPZ+psooLG6iJhogFQ/9Wj+tReFAiZMzhwCalXyXGJBZxEXcjc
+E9rzh8FOfL19BTx5eANYOpZENA966ZOW+B1E72W6yjJhwxaJKLzj6vD9RPMAvsglVvpb5w4kB/+
xjhiInqOfTFOTl5TIkHERyvibDGLQxRtIg8r1d97eNHvkkseLAKUrdb6fSikyhWJKUfMyqEXIwjk
zbCiYB6CHnW8DYpv/JfpeKZm7TdpqdTPMd0qHeePMs2InyRE/ajIcLlExDt/fEjC0p7fjf6XwKb4
9RjEtiXeu/xeftS1q4D3z51huO9FnqsISgBC96jLbCQ8z9RGFYZDq82QRPTfitclVcQtx32qH/hQ
NPW5Dv5yaqVbom2NlizLBUge6ZuzjZfiWgHxgHyvLyfsvE2luuNFDidRnaEyfVuBuL2qD06n1NKo
6rReFbQGgnRx0Z2nPEeTOkOiWHd0pN3R84RckhMRuzD7d287Y6KPtnHDmoOlbjD6C7fZIgLAZqRf
kuC7PmDIyZ28lPU8v58ITZc1Q/RTzhMzkvvAJENCBg+aXuHKteXT5mpyOEuLv8f7FwiWqIOXYogW
oYsbfVvERm83I6TEvFegKKv9QkDpIDRj5W6Y85X6ju/j4UpwiWfUyX+ILYdiev7LVcxBTdcHXaJh
XOd3jCa/3QwArS5I37SPI5Rwt93lwulk0ZNzZXsKSxVMBkdtAOG4Ac0DrIaI/vemrElUbdQiiaAi
jfdsso/HTuEGBJ6dIBM8C8UWPKRRxJo5TtQhGbdg33jyoMLpEcNz8a2a4XfOs2X/TtDke1iHlgsi
nx5HGQiMSNJkuf6lFzNMZH455ozItizR8UeFpkNlmVMaj23BkFyTnC9soO7872og4lRZSKVloPWN
gqCa5gCjMX+8efGyTibv0oJGwWNXaiLS9GT6I+Yjon3GprkGft84zKP0aTkIp4NgwEoUP8XGjusm
Y3yUe/mFWBJ8yTKUha1ob0tzahc4uIGHC6PXIlbIp8n0ajehz9ChceK/6GsK/ooghIWWg2Txc1Is
p2WYJrcFqekcS4NdrmK4fkbcPjbbnGy4qwa29oVs56NHiAjmfCBgoaL2oztdHjNYULHfM588ugNO
B4FPNf1Kgv63gLMh53M0E6INVb/CmM9mDYK6P4APRnnskGN6SLlovJZeIKNeUe3nn5vI8WCuNT2F
2hZSnV7aU0x5PydT8X6hqcIT/KS8DXL6HpAYe68C6HreSb+u0NMHBDPQ2dY0df8LoeaF7gJgLNWl
C0g9d7rjS2aTZT20ORR851+v6dmaiF6WcCSejJn9TyRtFVVFJzaL3liq0LEf83xD+QKQvqnbYoQX
VCU8Ydfu9RP9/2WZ9v5rMUUWt4f1U16mFVSxdRksHake1v3/lSAlqmyCLDXva+yBiLfuf9OdtJl7
Dko6+W1ksvr2KYrRyvASDV60BI/0jlwFlltLbMDZvenflGtigwiynd7jgTl5JH99lRmUgu+vOwT1
O6KZx9O6jOgx0HeXTWg2wWbkPD3dQewVzc9qse4BZ43j+ALkANowB3GDfhL6b/EdtfdCr9jApqif
ThVw1z4xfcaGcAWw2q8voh0jqdgQkJGArXN8aEcKIQGXxa4IyjCGEDHLVB1OGh1KTRVTafAPFmR0
X52BLwWVXavDf1Lt9RmMGfN4kQb+oKLHj84uWMz2HraUREd7uSblmBuQvt/lEutA9QWRushobcXe
ZD4uLHjZlFMP0A6A6sPZsx+CQ5Sh5zrscPn9/ueBex21NOuCFgLt1kpg4/RBt6cgRjLm0npF5C8X
vHAouE3aiGRiWRRCsDyBmTUxuufCHZ1kAkPvvSodnrIvmWu1ZT/dOfHyQaFNn4mjcw7Vrri8C2zt
cbbAUpJR1AbHYiUKJidLbEoaemDy0optgchVC2B0wvltbetpyw5Vf6tlsdYsf+1i48Qx51qplsby
CP3xSsBlgrDtXg7U9ULFd3YAA+vNTFAwfmmh/5N8Nrw/9EX6INlCQmDFVLGr9Ygo5zojtGI0prxr
LBX68uY+ByApmPHIWpzRO0gcOdNvZrbAtbjDWXJHSUiD8Tl2RacuerWe42ag8OZmxG8d41n13x6x
Lgc9H3jRA34CVr3r0I2rAtNA4uBD4Qe/A/RTwCXaLPqGJ96XVTr/3H4ZtpuL5EePyLufBve+Bjw2
zVrVG0SNG7hpPUlmo75J4y0Yj34qPCwpNi9NDP2OFr7rtS548Af/LBRVBRV9mQbduzczZmXPhtRv
hotTPM9Dx2E49Jp6WGTovS9oMnWG7ADTuNbDj7JwEJS6i34ZrosMN1Bf5rPzasVbYGO8VTyCbBxm
qfXE1y0DraNErs4eGDBb/AJW4rSsEPcN2TEOQXI81p04SjXnK3sauruW/K5nIJImgmUK8h8IVbgX
3614I5M/u2u3uZqr15byBbsd02fE0Y5PlVN2c5GJaFhTiMSXngtZ0nTghgDl5H1ftiDKnWuMoYGn
WilqlnM6w50+OzqZdQBh2J9mUal7P8u2bqFwY0elGRBiS/eRZXH6eFgrMHxZNsJ2JZoo0N0qR98f
h3bjcYS3flG9e2afPh6pyfKoHzxhnn1LMfZFim43U0xyM9lPEPjSJBgHo7cDm0qPXzT/IL4egctA
Lrz9nKvvxTFgVK9mcPTekguuV/YrMt1H2ds6BSAWYOo8Nnh6DrqFNWfibavDj1MOP7bdhn95ti0d
cmlKNPUEp+EMJRzU9guo0BSBx9ErJTWT6f97wgqQDYXXFWtrKvtD14UNc9qpFuV2/t7K+Sx4e8Qa
sA45dsemZ46VHyzI//g/UYBIVCJcXYcJr9ibGaTlZwRpWSldFGLALrbTq2mirSt5u6lFeEgMic3v
8UTAwNSVMMFUly9k8pBFjV+2W1c/7DvmR0tHF4PHZ2fD4NbQaXEq8mYuuMUY2WfmzKqTQ1LXMBt4
HLJGnm2BjzgVuYvNkGW8HouHX0AITCmzk5hDSa26CseV+WNM12ogNBm+6KRnNiS/8CBmyVQCO7Lh
J9VFgJkn9agz99hexdtKwiMOV9xOY3rRQa5J8NGMiVO93ydKGOPA8h4kxEobAtMm6Ow46HMM8vQT
RXG1Va16cS+XBkyyINwpZzJ/JLM50wzX1vxsfMY5Bfdt07Zj0Wu5/PwQ7EyDNwTFY12mPs4TAgIR
VbX3aTT7re8Z/T8mQONspIz7ns897Kp+yYfaXBDZ+xJ/QpOtWvQTCi9RWoiOxKi6UsCEazlnZquL
304ZZGnwUd/Qa71zUAYevHMgFqjrrMIl0AHPV6kLo4PTfG8XPy0kPyojzgz/xiXDqdgnMt00yGsr
thgXKi4ZLYXCHkgvGisXAQu84XPgxZQZO+hksZlkAAzaMU0ycWKzSBuwePX6tm5yITPteDIMeVxA
99GPro3ZytevgjV1GqQbr1Usf1NWqdMlFiIzV6LHjIqElXF4d0qQUPaya+Lm6s7mkFxaM35fPuUG
acaF/ps88WzgqidP5wBn9C94O0DSjHjyj0rDlRzbNC+c3XgwNcibaX4tK/xnUMYgg90a8L+hRT5e
a7lg2WbVWoQzUneiNHLzcPedc3Vst91B9RQu/8Qx5LbiSiK7NfnTi6ATuomjRi+SVvhMVPXl+Jdy
TzcgEgL4maYu7hG3YMDiAISXZHpaaixcpq2twUsvlv1CksGArUVJX57r07Lm9Mdzbv9TEuSHn3uE
C2foCoFJl4wBOMYJB65JBjhYRwoIdHe1ehKulCsu/K4tUJb6thmzOlzDpWX4OLPEUpiu/vwm0sQ3
ppaEcX6kkVyVis+uoqBq8mikgM5BTh0BL3b2wHfglxjgy+iNRi4Sj6V6q7JSLYxMcBcw743I0Zb3
ObvpM4Bpn5dN4B3FOApnT37P/VLe0xRWn3McZAXWB2ukyiklNuM4Z3NsBCHCgogdOx8MAHeGbZuI
KPt7fM563s3ENaLVVl2G4lNSRNnFLHaIPbZyUwoCkW8Lp88G8tnCRTFmsuqq+yNRMPeM15iw7Ar/
iR390LOXfJqCAeInWUfw7sWebrAuJRcVI0oAzxxxENccPaVcJwphdNq1Al2tV6lucKtcwwbAZaDV
U5s8RFpdGTi9qW/tNXKgJz9wE9KGZQSopX+rrHKye98jOlsDGlenR51+r77coQ5dk9KBfQOdNHGA
QkZltx/sDH2Od1bluuhk1PupxPG1IPZ0tizq7pCsbR+dVUixGiK6aZ4dEd3ALj5QtEshjxEFOqhH
mcybDX+g+RSKLLD/Hep0YMPfk1StBN+L5LFSa+giOn6/btskfUt3Xoiab3iGWReUg2PbaBFsadKN
1/m989nbxmA+aBks9FwoeRw4ic7wTUm6mwa4deomqfvEVL4yyQNYxCB2/Lu2H/eyZGtMqLcbTPLE
1JQ0NN93oWYi7X+9KVaYp31Bp7hWc2L77rdq1/zMbBbyjxzAAVj8ijB+gfRwHjXAPAIbIt2zw7Gq
DhNRm0uk/uuzk9AP3wyM8KyMPQaxENhW0oGMQYBgycexVUZQpE3Ue0YSiXfFMRHx8Cf8GwzzkfYH
eI83P00jMJwj3OEQRNZM7G/MR31cRTSiI6RYJx+aCwzXYBAWav3Q7ozaSfqXn3Vpd6Qm7rM8AZHq
c2oN+gKvC0mqkzymiuvemHaaX9glx2iXYIGDQW+dIQ0ktHKWq9yPoY1Ai+WGOQ4zQ+VwEi6HnJjb
5cqdM+DJMIXUjlo1NTGUVPQ+zjQnQ3HSYnt+gTia6NbeEGexYyHd8IobyrCtZ4reKsoz/JnNhrqk
CpSZcJTSLJE/ojqqcti0Yf7b8uCmOj2CfKSZbRCEDbKP9AeWjDTNdTcGPMdn7lp5J55qFxzAxzbY
7oY82cCAQ0h77y85iMpdOLQfrNqpH3ZbYgSaCG4n3/kYhceapHBE3d5s0Omvi1ALhXnY+pbPTqqY
KTyS9G/ezMt5rlGhT/U2kQCisar90kpDLIeEjAQx2lCdMlLKBA07vhCYdkpBnqi3ryGzivCfZk5X
p167MzPA9124Q0rNcdtOeAI6c9AFLq7QEtd4xX9dWrfyJnxTwCyv/NRb4+H7Xov5GZbBV0r9XqIX
wzJtFxX+2nqoTHkF1GHaplPF7WtIpVb4j+NKQd9QHPP1vZFh9W9+qLKzsS1Ey4MzlpHk883wACLs
3Bq9Xg1FXoeZ6vIwtYoKcnvfDXO+TcSSJ5WFfJ5HVbjNEE/KTSz3D4/SFdYp21cHQKOSMuIVwt8S
zCBIcA4ejcZPZKJJ0GaSNBhvKxuN+1r4S4onvxmgLU+f49WaYSoD4/VHwZUZwEWfkI+/ZUy2pPdq
KwxRcWK7Gfr8LZ5hE0pulsA9/1fLGieoHGxrsaAqYm/OSKnY3497iT4SRiOm2wJr7aX2dF7ODWOu
WEk/CLlMsEu2EnS0bA8nopEXfkI8Ywjgn18s29zQQMBR4w8IFIhXGmvj5WMuiqx6+PaXAKJE9sRC
huZK+5wozrazK32QQejDiS/AA2lkZn3zPMI2+X8LqBKssLKcrM7bkj7pfOZ8FpPxGKc4ceTJRLJg
NvJ2Bc+FxXNYD48T9mKlpyLIhVfkMYmo9j4Wo/Ry0w6IblvuHVk/WKtKMX/cFUvZ/r7VgzHExjzR
cMjS2boTcd+OwgldCJSv0b+O+zikTo0n/maaaPJFj/AYwibg+n6jMKWdS42UEfKgXvPASlNhIiJR
vTY6Ef/8yg0FeUljJb7Y5GqUehpr0Cyfkle0UQZU/DOlirDMbcKTNFRTFMBrgoy4xKkHm8AsNB9D
LV8hDrUNRz+GbsU27uQcCw3HGomO07ImkS+7OBRn8UFpEyxf8Y+IxGCPF/g0gKSV67M/OHYFbQwx
8bvtjmW2uEReT3k5bdPDkiqT2S514tCBq586tRoP9Q1gO1bkgcAZXuo/SKgWaEPPaAZE5MwzJpok
MXn4SAAvrUPohMVZpj7C+An+btuc+CLyT6RmnT6l8LwH/qsHdVlGNwmwCA9V84Q3UVK6otGqMPxG
jG1JxVgAqqL4s1zs/u0l30oMoKcqd1zHFG/PIek2s62UdiKu6O/o6jd6adV4z4YM/a68+Zq7TStK
LX+Oy/IaKmt8OJ0QzeuA0xe+eA3n7LWA/NBeaZH/dw4RgV59ZmT4C/aciGiEDdcc0BAI3AznsPuW
i7232YUQZaqv1DD6R5XDtEkbjnbHmx6XRg+5tRA8jpkZBJXpji8NqZXatBJZtywBqUYBMGGNJm68
8w3j37ApeFwxX1dDQvpZWG9XXBm0UADMNq9eVWWAjpbYq7H+ZNmnhfvhr7C/yWtndBfCroQbEwhv
kKzJi0zgoislE+dQZbrA4PRoyG4N0tV4g1ZzcY1J4yH8ZSySofDwlWgomEicsNAEf+EDPq7JrRue
O29dVsTFggCTvIXj4c4ZaRERBRdKkWBtdy71FXuOPa596gkNerZNtPpYRz0Wz4e30QY1iXHBhclg
xplnMT9dJJTQ3W6fzaP2xKInZv6MH46US+VuPEK279we7W6OL8VGnlv956uhjwFSEUWsAmqLjST5
D2NHjFSPub4b71n0z9OBqDBUVknHeXYk9/1/yDnI+X06dcTFLX+6up1xdI98AtVfUzS3viAA7qqY
ZuK1vt0N8jit5SLc/t549xUZr9EOzOZ9PIN4l4FCl12aowpxpe0JanSipdgV93f4KR+njM9o0uTW
2EKfqYQX/GZX3K8kMtYQE+RfhYgqR4YW26rAQE8FetBLRVHuVwWrKhELarZu0KG6dnCnweYbpNLQ
gFNoITFS+Z8/GoXJYMOLcOG68D1LcGSTiEWnQCz6rIRHFgGhhc+MXh1IuQEISPk2EMN8ixvzweJa
u0LUlbTThirF58bWzKfRfgKCgfHWvaC9TM43zkn5ZPcsy1Nn+h8kbnm5HY47gLqqeHb586jkFK/2
zkxSVX4USmu9bQzTj27ALs+Vr6zCOB5heodQv2qMB2p4ap/fhSXGFsAC7kkyzds/onwWMSxKBXfC
WYTwMqmPnuTi+nCEYQ4Z97xyw0PgYMvjfQ2znNI3+5A0nEeQ1Cyj8kx3ZiWFDi4kzbMLMSP2l80H
9slx0Iqn5mm6KWJvSS6TOHdjkx71VBv9ahN1I6S/Hmn8onrprQDOLxfsti7YYoTNvGXhx3CI0IVs
+qjFRjDt+E13uNbg4dLTScD9WZdlVzTU39Sf4hrIcvW2qQWZI81TfwJIkrk9aY7XpdrWnxmhevjm
a8sSz88zJb1EAYa3mUxqRW35nGkISD6HikIjCw5PtHiEKzkIaRudfTlzb4g0LqhzwGWNLpVojwP6
diqbPGih/82vHTykpAAtkp9wkuCV66I+YEEet9fgPP2SKGYpV5Zb/2U5PdV+ZryAJXOXaI90y639
N619X36lae97SngtsW2HSq36s1q0szg02dRlhNwr5DO+GLjn98lK8xKUFOR5cVsBD5nPAT4IcnlG
aZp75H9spSeOoP8D8BV+XGizIX1sImlf7VuK0bWdLVb7FDEHUNdoxtdfIPOWblK2WGVgztaYF/5O
NIXVECsRmkHzrR//Z1MB3L5Z0yoMigEUnl174mhv3JlSgKJF/NQSC93Chn3nT+4lbWZoTvvipApR
MMqO6wmJlrTWO2qm09JoGMUTHv81eKssJDqPK9TKy/rzeuWG6OUAPDIkrL8DGPkNUJyMIhCVpgkY
nqYSczB9JToYssanuHmORmHVrd2fTj/jIC/HTD84Hp0zoiDJJtwpipi50xfdQDqw28jRik8yB5s+
TkpJKvj43DaKv49bpQlIV2vzOOMu1EPXWo6gKGg6gO7DTmHuYkwnkk+2qPKeE1pZN7Qz+LrT9fSK
r+3hyooZoBDKV82ypijWbBw1P0U5Oan6dWme8GEXOBHPGVM3uAgb5SP9tGGPEXBGNhAxKpJbjz0w
gEjxDEd1JpoYArWfjdO6qmw+U7kCHrmXLEWjmbgFDHWaJdCRomp9rA+EdU7sD+TfSshLW8BCKHmt
H3Uf2sFSvAq8cuq2NJAdwLMqxOJlVLliSln3fzto8aG5y3d/yvzs9si6kCzAbbWYqq3hJXfL1+wS
hfVHmePjuZqNUCZxn59zNXRMuC2L6Pn9X4M1tmz5Y3te0kjRkUt0FkzWAUeeXowAbp47x4ubEmDI
N9gqY2Je713pJLo9VSbY/aSFlXrHQqtZ1lg/LlfMXxwFyOktouA6nrIUNPLGeLbawRvR18S0wVSr
MgTYP8HbD1o3CuBBCbMtJhm1qJsr6Zg2ldwfUX63iy0y6qyOi3PVttDdP7mcU5ekmObVJDHfPzSa
Ra+YeM6liuPDuijizsYuaA72d/52jLoddZDKksI4vk6UJk1mrJ00ej1asgY+Q8zMk2QWJE2SXZDQ
kDXnTvJ27z90WCiGALxx1G2vOPmMl5JLh1slUleRz4d7I1alfFgTKON0NmyGvoIVcCbsecQ+VeS4
gelqJvpctCD3Po5xZsqW6KbiYUD581IVMHT1Fm5UriZATy109/ouWhCTxXN+RKKMLQrKdXGyBhIJ
TmhLMFOinAQ06IK0VA49TssV3nV6eEeNappx1mHeYUkDWDJbqOspC5mBpF3yaRgQaI4GNFVawDZd
yo2auTu2VXdWlReJpL85RuT8GSYaBEuK4tnTtZTQ7ABXbg4EtkYzvzx+3nNJwcp5Ngx0jlLGeFTR
2PX7C1uo30j9KtqEqFCQYlyFA/g6wbGfihPxxq+VmLKckMpHYkNNfn2X5cfbjpeImCdWJlBVhjUp
3iuzXkuLanXIZe1FHXk71kMUmaAMxMkqk7RSJWwQ9ktCNIdB6uBK7cLjc2LkN0n24icIQh3v04cN
gBhAKTziHOn8CdAambJLofkjuwVmJBOPRunLdGCQ7GwMqgnODQ8c7SMt5PlkZtGq8OSz4Ph6LFIF
FxnCvoUY+VBx7iLIu+t3X6Nd/Zlm36OB98cIKk/O1eRwlhQ9+yeHRKe3EdyS0dHOZSAsNFkOKvpF
0a3awS6OQllOZfKqXGT5yuLq82IzfEIKH8xftDu2sF/QsnoD03ntlXKeiws2vDN8varrgHT/asIV
dgtVfY1iZkCObAtG/7FV1AccHvChxIMHnSZzwGxejE1W190V+TEnSoyO3Vl7mOab99t3dxXyKcCP
JgjIupg6P9Lmwe6TbZ0R6DfiHIkXZc7Ovq8EisjmJHmCtREfbxxaRktOWxEK36kPvknz0Y65vVkY
PDiieKJhGo3HCyEjIBX58DoKL+K2uA+AS3lyi4ZZF7M4RyLH3hmduk1hKUVNw+P0o5whF+Tef8KF
Nzj6tmGtlkEeYEFwQvFQ+g2mSV6q9UESLouZ1kEgT+hDNIH3F9wqzWK0chhMHjq1Vco1ems3BeHD
rPutGV7pXqEY440SQpGUdj73HVxXT+qg41yG3KF6HHci4u99sN2I/4Cf7ob5hEBTVfLDdkmvmYwi
+3k0Zx/pfsNX892XGaAoVKCMsl/5XO4ZnNJK8bfLILalYOboljH3In9+hkvAqih9CWiPRCMuYcsV
M/Ffs1OZ7c3L8UWODhj3xzvjTv3DaothR56sqE95xKrZfyB3uyETK9mktDKchD9QunZAzn6oLKvZ
Wo6yazIcS/0nz1S8ftTiiG0kO3iWZu7a8OF3ePAY1XffeBNDaKETBKX0rvhFoyMbSxGutpwpnHf/
qkp5Oljt7nbJ8ZmL8m6SFb5dFH7X7oM+3JBX1OTG0PFV0pDnTc1gNmd0f9dq157FAvphfYezTr/K
I4/3HGfAX/LqrLMYFyhfOrzgGHUMO4mjB4yhWrWXyan5GSuzxaP+//6rCa+/2wwlDH56UndSH6MX
HOd1CBagzV6YdbCIB8tWB82At+hTjLzorgzyGRpo63wK+PwVosLg6wPKSmSDrIaolAOYkhHbz9Ce
/ZAqVMOy8VjAdbbmgYJNtbhBOMB5ff74W2Ime4BweTVu7y6HBgDzHjcj4sij02YA8HVcMlx6NK8h
ELdfjyMeWrOmACQmZN7o4LMURq0rLiZk1rXmvgO3GMrl3+K7zsSHIs+PaURwBmC4FcdKSGX6xoV3
PkubHoTGGA88fcDq+jqZoFNhrTGnr37Ymty7Mpef68V66qMze/leD93We4KBRXBlmleMPzPlQQhy
/g2lISWd6gqzpkta16gQTlALNwXfuWgvIVyWgB36HPBndbGWHSY1jFEyU0tJXMIie1gg558mcqS7
1F/ckTBvrYrD749Ko6LR7ILbhNSCs7FhQkzYbMZowMghxeNoUpZbvK8kVHJ95jv/eBpMpddmIUf0
wGw+Hfvfm3vlSSldqgTKyLhlb5GfptN8BNwnEyb3vGIvHSyDlSY9l2saBBPK1++Og4e9FUmk/pVX
55lxTruqAtmzuwZXhRtzrp6u9lWjteyTebjI6CabipcrMEWQuIx5HZmpuX05DFwcVQy7kO8HpUtK
BxGVrgA5aWRWbxqoYB5wjhQIyntdlZFdWQOOpH1QpEzzYgylqWexmlomEBGj/wzKL2YhFnppsmQc
MBZvrJ27DifGa/WNCYUDIr1wWSAe6HIVnk1/++WleMb+rBWPDkEnY7L9sPaBxxW5Di0qludsaScW
DPxqa3hoxud1HnY4/r9zIN7WT3UUPrVpjyEAJ6EPmugIv+6xJqJ8faFFu32wmf5vafYAow7Dwi8H
wBtOVt585PyiterzU/DNHZDfeFkp2bb1eRYs4AVb7xPr9hFUMB44G7AUSbluiwai6kVgNxtZtDVt
fNfEO+bwdHoozDhBCZmIidcVDwGCxp6rK/KnP9+kd5LrktKyphYKds1CiNfHTNNUcUX7nJHQakp3
Qt3jcxfI9vWZVhi/xmHDzrsqCJk79nC5iGeP2JgDgobZTUk7EYsVZTzt43sCEj2i1AsRaFBkX2lq
1xJwiCN9BcwoSgdD2qz9IrxwHSEZPWcbUU/vMG2kDA1HEO83k/5ouNCMBL0BKWsVd1KzLN1RC3yG
YetLcqsin6y/V71Laa9HLMrBY8lrK8lIeF9kztUKU4a/HVXmmMDU2QcbwCX8uApskDSDsjUGivUz
9ShA/59hQbOf24mA/d82UxeildlKEdeMQCGePm1awe0FNDnz8r+N1S+LsddJhjoAWXS9qJnWexgD
nmyofOCB1VG5eH8MvdETIdvE9bzx+pEcdYbhX65M7I7KRhDtU73FY6XYfPPmVOqheo0TC6Ns7uJJ
DpfOm9PWCca5reFrFgUHwFhFMW7Ul0/7gBfVEc0lYHTh20EoMSSId0L3sEjjTz/YVrdx9ZwG+7JR
u3OuTX7snsSML62Rg8yAueZ3kSK0gYWa5RausipYXq9SRln1KGCTMFNtZRRtMBIKzeaUzzf9D/bs
K4jJxNodP1owgb80VC5b7edbPJr00Iwu+WB8WXL0oRwv7QEKhac5HjasbhjpU175o23LZZYAJFVP
M1RU9qNC2glqLGaX1GBj7MmG9ZSsx68ze2VVS690sEuAPHKGqyQHXxOMJw/yNL5IJorX+jk3USZh
6Bc54DqLPtxFiDI02jfhnFGSOeiMCm+HWJXfkclWjR0nuEg0zFytPUIi1nfsH8V1dKb6USj36zX3
KLYGlizMghDtQesw0z3wUck7dwmh8/pnqYNPxqw0rlI7+YodGPFCQWR8Cya9xQNVMvmpZ4OvmZgI
+VxfTwiD5sTqhdPz5IBUPsgDuOoe5jKKCtaD+s35ziY9bviap+qIoe5y/LK68Rm7wvG6bB85JcG+
Tw/hh7aj1riNyIjZ8tesFz5M9BKti+pWWvgL0uq4tz+iaItTb1RuZnnpGJ3M2u2cCz0lvsoX4TOJ
Tr+ISaEBYMvsYjQ4pp6pvaA4V7AUl2gCoSrMNqrnH02UpA4DKnFp5Msa7bvujSavlkgPuAZlKzoc
HJ4jwGmt4TMvQIX6oz3YvxzDa3sarra99i2vkrc7APCl+v1rWQ/7mug+LYhE6DvsiAA4fFB3lCV/
XEbj3DN2FY/Sd/XzduNVs1QaDdJZ6ojnjEbwnCRI4u0bVfqdlaFpcJQClfWPKe1l7wNeuNk+/J5n
u1sDdxOQ5Mpu6UKiaNM9sDGJEEemZPOzKdzEl6fstWRGtGsDedATY8X9QIcX2nbHpcNdFyAz2t8k
D6XAbOtxQPpGUpVIO/KnZwYeER2/GVXWPHvqrU6OQ7sFbWHSLW/+ynxZmb+fMHwMmmFcMqS2kMVm
lyqzleNm5TL6n8aC+wLmutsMeVi2OILQu8KkhfOgU2IRBXgYfnqmWyQxLibi/Nd4BveC8Dnx9B81
H0ltghbYuj+RRH+XS0MZHWmAjcZT8TzX+GLJAhroLla5HFJD49Vb238BXaAcbigWuntALft9pvFI
DilsArWjIOE4Y199Py9j7jFW8fvKBWJRZqHFJY+1oKPS7/8Ru1t3r7aNw//hejU2eyytrqNSbdlN
pqf8YRFvxvrMhOA0sN6TNaMH5W7XCEXA2YV1PB9ntOHxMe8eDaNHLEb9HbhMQ3rzFlpCb4PYaMX5
iNLjjVz+2FaYF1EJRasvI1LkerjddxuihqfIzUeAAEfXQkN3ZX1+yrUsSC3BISjU+EUJ39yPIeMo
6vbqPLsSBfRUVlvpwCa2Td469aa8WbHNQwkR0IV16G7Hg+UKGza3CSNDkxiJhv16WHcRCLvsU5gM
XK0bQ7R+7zPbeFFo+NaBrCE7RCANSlXinVxbY7EEtTze/yuarM1Yaq0Nx1l0wsYM54nhCoS+HSu+
UoIx3w88xQGaYi4TOauh78ZwFifuA/9tY7u05/W/gz4ziKr/2alsrRPK/M9lLgye1pc4bT8mhZb6
s+WZadBf49gJtY7xqJW0exlK/suhns9T6dVMO7RkK4DggMGSVmHaC/qEsoHJSujG1RMr3ro/dqnD
PhvqfBIP0u3MmCVSoHh8fV0aZdD+7dV2zRYY4Xx4QSq1IA/1KdJ5YepstwbYH9XJBw2h0mevqapx
O0aX6jG2igPB9ATvw+Oq36bRrYC6QqOstvT78t6Gsde6cTaqggM7mPJZzEwmKtt6oX6JET0GUPv2
4pMeWB5jJgvUpoCL0Kvd67RIQy/Ths0+8p6nIi3T5cPgsspyPezes0sysvk6bsLrdVmQURrLwD78
j8P+i50sFcvE68H2fgl2Mv32Eda6FApyUhxeknaj7EnzsH4CghmxepV17loej6JfF+O4Vg6ZxQDZ
Ybk9K7NFwIBByrY2g7s30Vc+ZD5152CxTpI5Qi3lui3lWYqn2bqbSEYNo+SxZGMr7RYGtO614XWM
Va0N9LE6rDn/jdQ4fLNyluh2aFQdu4utXHrNc7a8qjOaIuyfMtmlw8Hj69eIBCdkDMvum7Vj1H7+
oS/DrlK+VngcMacRvHo4+ia0eBUFb+NSGazl/KSxkbwOI0JBdaxJaFUGLhRl0IDmAgPqIN1jD60D
W/75NzX9V8tLLgyLM81QLSETHCxE7cP6spOJpsHWSxLhuzWDDA6nxCOSjxnFfqqxMjpCuH7cpLJ8
nDm+XZX6uNY0t4zZn+M/RF3YfDKqnPN9c6mHYxQ7pRz9tDG7u4cAnWynxBw762w+50VjpnrH/+1B
jQHdvxeNHCddExxZtYUcYDbtkTWj47oB6OWdOGWOPKyJfiarEutdthKh0RnNkMma00uVnDWC+JE2
P2xg325kpkN++3AKt7EU72sevKKeNxt+5oCUGRpxRoORSrZqIiQB2RM1zyC1U8U0+L4gWpgVENp9
6nhVapTNBQ8j0dOMwqh1WbQZ1usTYPaR9TyWPaEXaoFDdWvKaqKHuOAh+0POvuiOQxDCVQeYIcrO
xEQAxQ7ZSK886q/Ob1UEXfXd/ig9o7UnKu8eL7ANrs7+lBoYmDxCTPKEA3pxuNcV/ycJndVyYcno
NlDitHVNJngZf5kR3FgIv8D9JWOpYEKYq9ethU4ZN11xa7gCSu9+TxzuyE3jfnFaMNZP10rD2QU3
MnzTfKvptLSmIPjAHY6Hr4nrLvAzncG/Yzjby9t8aIWPVQsRKQsFhTb8fX2bjlCedWRoioDdY4y+
GVtI3cboBB6Z8dlPBK8rrVw2oLfe5FHH2qfVvqQnBMza/NZ9tP3CCHMUNOPYZyKrGKPDlM/uIOJR
CFtbIyWFpDYCHptaY+Xn62YtveqtBVkeFYW37WdQERzD8g3NE1YBBq3/DxflJAWe5+ULrwujK3KR
lnFGsM4/SvE34i3ETvcWHVmDGyvcNADD50CzxM+oP9OpdSrP2Wv1n99DA4OTYcoGxbTNUv9RYQkL
rRyh+sl0AU7oPOKwbEcmN8x9/R779HV1YLyX0Ryx+TGbP9IDh2G8YriYiPUevyd8mmFMrGDpOybW
A/lVp5agfIx4cwJattfS+Gn6/Soad7phd+Rrkk0I+9Ef+Ob5LYJvUyX3+4pa/nUXBTc6kXQ8o+6u
20WQRt/vOLboD4bNHJA7ZQqBTOOAGLELaNK6ZD6ixxdh6MCzI+Otbv/l3F0UBfPxHq+kG6Qpj2TP
BJsIQlVjSMMx7efFJm5ZgqMTA0PvGf6svQXVbY8PDs7/8XB/Jno0x957S1UjwWiSltKiltawx4cV
Tg1+4G4ZbBNlLbZ2UZT90b52MEKwFs7rW6+HrpbhtfWPazXsZ2MgsAirJgMlkAlJDF00wnTsiyDi
RGeC1MhItNRH7HmKlmfepZH9FM76qRz7CQweARRRiedRjZyPEZ2Noeq0GKjRmKZ12deJjOCt7n5q
vop2jGuu57crg56kcMz1dp+6iY6Zl6CfrWwSXsIRZGyG6Szom0++u7urzNgIJAFW13t929uftEFc
3TcQqoVh5ra/BKtKiPEgq0bmIxntvXboF7LKgamnI42p+HGXH1Tg8ccW7kUENej46aQIRYwlLB+K
LoXF3fleYvdtSkBHCK6O/MOLJxRaAG9YfA3OzxEzydoi5R4qP+RK+Kq8ic9DwTXmpLPSqI5U6z8d
MmWR5YWhfFikOwN/SaRbzYYs22saO1czT9luV/4eIBCN/sBBmVAjbUrwmWMXjV2WUd2766rXrPij
45xqfz7duRbgvH3g1WhQwOxfWC4gIxpmYrixvB8ynD1kKFQ8xXF6IfviYruqaaM/OyP/oE+wDqY+
rnNbVJocasp88y5Gu+tnqIk197pzbjdTPdhnny9qNaXZFkS8AdDjLMlr6gxrtd40os2Ctw+AjGHu
zWed/yDiW8Rt7GRV7FhKJTuxl5BnAQu/+AozU/OXTWbJ9qFdzdUi8JMUwuZqJzBE6YOZjNuztr+d
GrvbVY7/NeGQLvOMGAmZC5R0L4jIs6RrNRg0A3wMgqhjcqmQFyoWqahTAtdN+FUO02jRjp8WIVdR
LaIRHvg7gtjpJ0Qnz7RaphFPFV3e3pEhXysrywy23CzXySnzMLHbGyaolNY3NsabAHUbyQkPUOJp
KEUncW2KvgTeSevkeUBazmEh7w82HlIY2zmLxx6EjOHTKjxTlDAFsGOju5fykD5FMuwDxM5zEVAx
GFZhTvIrbWFzB2UyVsN9EhtbSmrdbBJirMJVwe/nbghBwHQ8z4125N/tv4uARPjfZawYgs1Y2UEY
AkmMz9d64CYCedBWtobvkWiu0EcV2hJy9GpaNwK9lhKdzBKxnCPpgbdV2Wd1QEJFTgf8p2GWa0bW
Ke9Pfanptc+X6TeKWQTp3hXTusoofNB9qofPko8nCEFJQYqLJ+cAhieiRFaeioKBzvEK622z/YBz
CisxZWQ6hurxCmADw526MwOq+TEHELhfT9FbH1MTvAalYYxaqeZ4bAG5bMCLZ8d2Eju7gcYRpe4Y
OJI3v0mDQhNSF9Bfq7MnAlafEf3uLWmPjqLWlZCBpN4qt+2dy49NBvrhMbUNq2YItOIh/z0wT1lB
8l6EuQeoDZ8zLXSymmORjYUmK6LH7sun2MiHBMsIhgToTjNVGwf074r8wgl2qkkzAJMbj4QPxFDe
Lol10Xp8iYijsJy0gpaKDnP1CepXoVWOHSlCtHJlsOOiQVH6yDkrO1UH2POyqlJ9FwbTh5h0/buk
4hIGtebfWMTm/wPfUVJh3gOEK6cPCDIDBqNutNEy0sFCpLpjYf4ycLXI6f1U3AfM4c7UNfPaPxim
QwpXC7d4hn4FMz6MGH9buXXLi4R/GP1isalxFIvDrBzjsUjdwjmLBnwJWvDLfa1xcsCwJf+wm3HY
rguG51VxyDRiJ0lG+2jMivpPKxeFp5jv+WQQKeWWLzCgwi4AjAGMpjGbNjYQiJ6XrRzXzs0sxGdn
9nRfCqZxMRD3IwJ0tTbwyT8XrW3F45J6zOrqWMj6LP+I7cVAKEYuwovQ6Dra4IQGR55oPpO+tQ12
goQxiXB01wQg+wDBrJusIKXHTgtXCaKEIk9E91nYS/4QJFI4DmdPMLudqlXLmwSn0HYvoEXes3d4
VKj6dyNL8rMu0V9sk8aR12z9LLhtBpdgCz7dyy659vY3Nn9hbAz+gnn3pRHlBsmOYd4n2Qd8N0lt
hg2Q4ZK3Sx3zRz8DwkR92LDTl74d+zg3Efb49unczJzSe81C7wZvGAuyISnK6dX37Zk9ddtomNgN
0lbTd7MugGlbpfwqMnBT3kkjVJTGPPxm4dm8swQmD9PsDdy2HYSEsyLcbs2KzGHwEawuZ7Z9X8qN
PZCpY5yPStWdzuI/c7dqa4lPKOAc3VNFZOGffeGaETGnyCP84wG7DAr1S9hA1wbEPTZldrnmhGc4
BDq7NwDsWpG+IwuXvyNMWY8K/DRh/+85Dt/WQv4yas1PoS6zJzOTEUWUGCxld+19yYyFdnqW8P6C
U/RPD+OG30BHiVOrMulQsegw7VrE1a2bBrwiuEvrRR1KZCe1UjFfiROt/CjwrAsxoO+Er2x3uRFw
syEYn7ivijck9v2iWwpMY30IPMUNwkXciccTVLkaNBpi0ZeiMXwz8ay5r2ZJic/8p6rHip2IBaQo
icKFIPtMdm+9oc/+SJQDniT6+05D19kTqssgeMn0X9rgjfYj2P+mO94ERUpKieFeLNu9cLDaJxb+
smHzGPFPR4U/QQaD37FetXldrYpQSY6llUPk0mhD6XhNbfZZWsRbV+e2UYZEa2gRwrlvFJ7qZFLo
+zEfrqlm2/Il3GDfmhO0R4UdUTaxd08+qEm9ItWWSb8N6gESaxk/I7fQv02KhUVBpF2ewatZn7qV
HpncW5d5PYSqNOtIGPSvRewLn2fa1E/DsUIqlYf8rPu/wPferjY7pXlxQMjpPzYHMOBE1woSeGzQ
JTL2ecoJdkypGKQuH/uAQqCP7yUqtc9j8uGMGfV13YPMETZ+rD9FV2XWaMrYZI6rLkKqtR6D8lJu
am8zuyrNSX4RCMSkYakA7EHHGvISYtTh7wWpxhqKsPgkyANrNjQbmehH9CBY06XmYhMQmpoZ1iG2
v0SIROML2zXKVRAKtgM3SJSqBALHtyBIqb59sHLJaSoe3kWwHkusoeQg14R3TCdtCNxxhNWZx1d9
JtESiblqnE/0iAbAmbxcITcHknpTdLeYfad7XJoWSwcXpOr5CrJvhlwbU8ERT2Z9yCOkWoBdTUeP
IV0hYPJ4cdINiV1t/ssVBIVx8z13LqEjWU5AarVV3hoxF+pqb5uAVHA9Bg48dEyavDZK7KVmGiHp
BJRSxPJuB5cEwnW0GvRX0vv9V0pCIGNPqCeEYSpA/pr4Jf/clU/+Jr4POlDaq+p/W5WO8JydSy4p
DeuTYoTmmBZWSCT4IKWwWxVU79dGmjVE9b34I/k5U/NqxfBbBD9vsQ/P4Bn+P2zQ/NALsdgVUuwY
uesbaeRt5sl3xp8IzPg33iuo2hwTH0BMNUhMro8jHQGzFhKPWVUxDLICMfz0V9UxoTKPNPcoQUBP
QBKgdzNfvasrxUJ7v92xuL9wGN3g7rYf9KCV+qH/+sKQ1dGRapOIwt98gzk+JDYA6gAm64Uzy+Z8
NxGT0sjG0v//cIa4A67c/bc5kg5gDg9CthE0EFQR7a9iJSabIGagv+DwFAp0OPLz7aU3v/JW2lOn
mGmTKYFc4lNAfnnhsFSzgakep6BIRCcsiyWAW+pxIY6xPF52zGcMixlsRNfhx/laEW20wUYIlV/6
T+Vt6pOCqPrRQxjR89Old6uJhT46Xr/PNRqim2+ji2hz3OUOlYCc7JoiZs+3XQT4OQ2GpQVfsUjU
ZGjBwlVQw9dLV5DnkyoKzFKG7H21bNNhnaj8OdgaBExOCtrmXeYSzgjw3EQKV/Z7hSPXn0FuTPDO
WT278noHsyjqoqTCw87OUHCneTJ9FfFi/zOCeWRV6GpPrPFzXx8CUSGd8Y5+phHa/85S7u4Txckb
dg6iZV+3suEl/c16y/TJsS6ydpWRTKxaUvZf2rHAvCYzCxqEa68Ag8rDFyLdfKRipePn6uah8Z7s
sw6DAfmcdELIsK49saIVuLRH2fg94RnpfkSiOiZA2tSC5in07r21wgmR45NtK6OytiFQ4tRp5fik
Lc/v1muFWkkt+lXEvuwyMGbv7MZcWeYnMJfme9SO91IMvmxNUqFRogCnHW8MHofMijb8bSg7k4aE
REYuxQ6oWRQICLT/psMGBtGOrtPsWnRyz5L+AZztFfmPWCaXnn9lmqoHaZVFkMLqLWDr/bnY+k6P
kWiW1mDo+oF7ISL3nKb4xqjFeZwD4SHHw2R0uWS/2SLk43C2zfo9P/w1Vb6K3lfY0JpfcxGD516b
AAzOY8jju73uN4q2DoUuvh1rxIvMTPD8W5ql4Szk1/m8jTjx5ZlzAeCUrLgcBXEhnwL/iG6ZY2oq
iSEp1LY+Xba7gKz+hrj6g+/sgXD9dNWQFpHms1lvwTuXkDhSUNB3At5ENVtRU0of9z85FIq4Vr05
aiMZ7hci3WKCE4zCboMe8KajhtYfSwanLdblxRpg5XvlZPVajVkANiM6aorj6bs96W90OZOh5izi
DArGhjd25/m+3aktRrNcwkFY1gZACyFtb3h152d9CyxhFFXat+P3M/NP+omVBridEOIEOA5LNK1n
n1s5uMa/aRUUxpP4OzvyaQBUsNNvTZ4lzi1qb74lm7erzusUwObeSi+tb3epcq2eu6rId1ilQ+u7
wgLGapWpZkBYdVtG6sLsQryxG69QV686NTz2z5Bsh0vly4wlqFilMQ9h8HNjKUcSWkHM+EkA8DHB
LeXTMC6EabnT1jE8h8gWNUhwPZ9sES//GHArxudF1189OuMe+hIau24IuNZrAUihh/24oU+J+e37
XLMzT7g7H5ZPEkRLKQqFf/1PN/XHdhQNAFvVOJgrk8D0Dbsc0txkD62duptEQKSyS62ASmpWZVFB
WPKhwElTC/5b9W+UMKfHtbYujUG3Xmdaq7/EXFk70tnvxKT2ufir5rhBKu+rU7KrKXZeX04g1JSY
iJGRB9ai1SsesZxd4MdySGEjij5miKffBfeWpQRRSpwznQSPojU5/Bk48mPC9s091LeILLF2OKiS
oG9+nRPn2XWEWsIXr4e3KwlU14UxOF3/5wLxfZzISq7aBXi3lGeV2xTcuh9ikz50X8nhwZ0OJEeg
hrAO8AD0SuocKJup5cxFm4rzAaPFPz0lSbh27xn8pIZx6WIV/1EKSavWFijtdRdBl9VjGW9dpOdF
oz3gGthQURJmBbOFAbYX/fK36M7ozbf/55EKnug+fW2Hdv1sIj3XuUCTgcxSc9MC0de2H7lC1bIy
bciS0K9mULPDLWT45e7jf9Yim1JjE4DFXyF4OeYI50VOOC+IeQ7wa1g8mnjhU4gZrqqsj11PPopG
tQKeuv0G1y+ThLmFcaX4jruPlAD/olc9+moeoB/j4MiMfLeuHozvCYvuRB/7JPEdFESlFGiR5fgL
tAoAiWo2JwXr+HJiafDd/mnrh1TdXXUHe1hDxT5DaHpMBx0TNlm4r1xILder/euuyVqGODlMeF45
mQx/DXQ6zfng1DcnxXStwxsUlrMKdXrOLuccEZ3QfNyZSinW9SAklt1AcKeDp3kN+fA0iWUED4OK
rwfwFGxzXt/Za2wv/0MNjKHNWpxhCPr+uFkxhNbW4sofS07haLvgTDBq/mHZc71GONDRQTLk+3c2
lglNzbtnl9JJsnRTFHIW5gt8r02JdbbSbGBpy5mIz2lKfMKVBMih2TPH/63HU9vIPW9TklmHKg7l
ilsxgEv2WX/XS6yoIQYGpHww8N/FC2v1DjTQnc+17jrDm0UNrmK1DmlOeZP3dg01X8e4QGiYR6CZ
j5Tt5CdkqrXcEp7SfRcRfvXC3iW57fYQPmz2DqfXeQvXfN3/Ecsj7rW05V6GZquF0h5AU/31FLcg
H5rTfBlh2lP887+BKKZehu1fKxvHuyYh8ohB2xjbqghyc0OhyLQZFGsEcCv8Itf9cTjRdwF9dqAu
wEUizE6x1RNGWi/xvq3fYx4pHhcnZkXwchW/87KVQFCV40am3A4VBGNMAqJFTq6dbkEMUkKAzTkO
KEJw8GulhS30aSE1XODOe3BUHvIG9dbPRLxD/zTnFiyl26rdOOmm+vQOz+aazIQ2/WmYT2fdBgah
LOYT3hX2riku3NcEq8BRbEVWn64L4DI4g34pAp8SCHqidNlxkWun3hZTKQY/SiztG/46XWimH2m6
HzpE84kFBJVEp0xpmwr8+HQrx23yUygKbDAsahOPGZVpvvRW5VieBD5PKaUDILgL0iSZIdQY/mI4
uXj6tSCa/Sxl7WwfgC+rZzoPf9MxQmx/MNsbvRGxtRIl/C0pGjEpkdNy0gp/Woh8lfEV+Hi9qlXT
sB9DYgRNUMi00vnL5uarwS84J5DYMrVgGifijpu8LO8dESBu0dajTak1KFs+u+DrgdvX///W778o
GvKrtyHGSWOY9bh4vDXTAvwlzbeF8fxtxSDwPffZul0b2R1GMBFZ7ImKG8eeEeK1w46FTI1wTlr/
v8L/XX0BUHNQD9MFcEZh0viLt8aE6vY4RnSEkNpLmobtM98JXhwHGbaCD1T1/FtfvPTLFwBClTxc
BBk3VEr0Nb29BhKLTy905smm0yBKpSaOfX+ti26LZ8JWqQ4FdTfPB0q88ip2qmVetWa/uV23+771
ZG0d7TIxsq+ueu0LBlD7ubRpU/If2YOc52Vvb4PwlQckpfQgWDWMu682YQkDfvVDVIydmKW4o+Cn
6udBQyN31G4p1e3sut6uzWlI3kAuaf0J8dXgdRjW+TS85exaR2c/wPq9lCwG3WwxoTCs1ReUzS8Q
E2znbInKSX723Vdra7cVd+4wSHWpWwWYE6sqXGm0oPGXOMIT+CgKNyDQ5RgC3fyslrD9BDKYubLc
yXkGZpVhEsUHjj9DkGC34XMj8qe4NfBpxnkaWesZHF2BWwysa9gWKD9qt6t68RMDP+jESAKkUEGf
oc9aygphD6rrJF7yUz2LfnPgF7PZO10SFIT3jqZUCzFAUals2REx18gZCN08Y5dfDZ/+r3Fvps4B
E142CBckEOmk7L3a3KLYRVAwJVY3fdG/XJEiDCnPwkCkrXUIqBSYl5ZcPPo8Tshii9UbRHPHAjU+
rJdo+AV4C5pXbfQF2IRkAEWLI7lmr3RbAeUIKc+gs8nV6orUzRrFzezQ95UNp+1tRKMt5zEzHGx9
h88mbTTU0VdBVX05ZjnR9bVWcM+Lrm1AocveH45bumASn41EYiQ53ba5MV5K75v3JyMo4xzOAlVb
HG+IS6AcclZCynNdrCBOtoZQUW0xFpBfPjQHgmRluUJc0vbGkloj5W6budPBDtlag4r6nv4lLAjJ
VLNv6VbnlmiyX28hbZfEx6KXTH0tHtg8oEpL+ek7MIwLYY4rObKOAKk1atZrn5CaKr4lIz4Gt+1O
31rLXG88RA7Z7LKu1QunR8PQ8qb/qMV6JFQx0PwWIPv8+XCvJJ+/ZR1gzmrA5/HNRVF1SPKs627Y
6WC+2alpwEGYEEZej3zmm5SCuCKKGEuNqnSx5wthBkD+RT3TuxuMy1opvuArCMIKGS2AFYh46lhV
gCOzkBGhHwpVJOfiBxqy4d09Dpe6/DklZUbZ04zFS3tDgXgy7oMD+mYQbAW8ZaISA9dbBvi89XtQ
iUf70yGbdp6yP9gh+bdpe9fF8XdW739fbkLqykwQNy2C93bgJ1pxMZOY1x1aLZp6NYFLHz2CMT6x
8R9fRaQ1WQ9mSsxI4i6K84fHJqktBRauLo2TfjhjMIOuPT35xP1P/w67cqYZBIHNLjiVkXJE1IsH
iagkJFWd48hh3W7RGG6E7j/MdBPmlVXrLCXUUAeWHAx92a5DvKkqrbXK9ZvrwxzGiDZyTPZzuMjP
obwtQumB5+qarn4UGEHy03dZsqYnuaYsanIigGOYK5eqzgNPEj2Ppj5uLXPlOUytaCrGzVazpKyp
djv9qQc1192s1LIgjY0Kw/5b8KpZ6/bRiJBCSf93lvWvmcPrubkxV/rn+/ok5yq69PJSpSBIvBCG
QYnN/e6eBexVEfYLkGtGrQ3eoJvsU9vEGcn6GkHjNMgE/G+++3oM5NWtaLsbPFrh0IvpOI+ls/Ci
eLFoWrk/loTYwJqXmO29e8Y05AiC87vdHSSWkw0iVHxeT7Ahz6wzLMqoxvUvPAQ1mqcCYFWBTgxC
u4WKMe0/h1LAAqag8HfCpHpINcq00ZZpWqbJu9SQQKcwi6+rPIYby8YlkV6bp5w8rLZNBGL7Fxor
qrkz7Dd7+HsGy3cEtBVZtcUWY8hRCIuxEQtss5Pw7DdKGpMXgSgJkK3efYPdOQKSCqu5usWSKy1s
50YK/4Tj4trICqPSp88nEY84BskH5EEtaAZeJG2l6Gkh+ij/OhMeIyjBKtWUH+cymrt2gQfPWjuL
oelUqO2woK3T1fp0TbGbCvp6/NCRfvTGd++PDt1F4gUu8Dv/yJH1cjeDxF4JV4a8nSzUQtUaBYeU
mTxBfBcy+DsVb/FU49Wru0hanpVZN+ds85M/Qkt2g8GK30b3G8Nf/iwCdTIxB39A7UAL+f8R+ERP
tq5rOi4A1P62M/xMZCx+4+k1B6Q+2oZhyH02zfEMYUhUwQTbV8xij4yQd/inOasXlRorREcinXXI
RRwKExJOKtLm3trzS8f34qgs2ZexHDz7zWeqtQ6vbnQv/0IDbpYVYRx5Ml763mljqJYwbZiH0Io/
5qhDH9ioFErC4Hlfcd+E+qR4KSm8wzcvbDxcitvw0mxpYMJgEHfb2Giz/VDdXjVvC7QvbcJYQtne
A4ePz17hpUmYsZTIzP6RoM95kGpRukX6UHSDdViYdntlhcd3yXqxP7IACTgv3I+cUnyZ6v7NKTQj
h/nL4DwzF3Uw08xyC4ThtkoGCSakLZGC+LrG1YnmrKLEHpLsrCmF+kOqxq1OSbsgaGtlqe9jIqA/
QgFriTE/n9eQnJSGGkd7EAsocyRFiLRfIV3JTrs2znHlB1Gg/kEQduHN608Xi2JfAuCWIm4k596M
UZ7/cTWe4joooTvTG6/UXdxBJUL/jlhMrKgbVYACKipTqmZsOncdM9ijQEx0VEc7t4KKKb+fMfly
c9PZEZICN9kEDjhzt4pt/pXeOu2OwfKRP7selQ/fDjl8qWpzwGaIb90LWmiOTKQdC+7sb16L99k8
3Z7Lh2v56bCzoJ/Z+NXC8oUO21MpBXAlKF2Nsg3ceYl3xl4cxYBP3SnX4OJL8P03qAIJCSRPslb7
znnGQgiOOULuNQeFDM7Qe612BoLKW8tGLKNtZthdlSl7WVLJrr9h2X0hFlNbHuok3/peSXMVCdRX
Db4uGX/Z6GIhIEk3IIvriRwm035xQc2XNJZW6nbiyBwS+p9TY5xYrCMImaSWw6LcEP6ZdvLm89Gh
7WZABdDA4VcTh1VyT669uD+iASW+Gi+byBvexqUYC85vkt5cuFPinFlAbZ/jXtIUFgdPyRsxXAjT
VxHxZLSF+FrY9TzO2Hd6ivyPBr0B4Dqig9fYwAFOJ6bux9ObCQs+IVxIfdvwlZ+JS7rV02UMKrDu
2qkvp1cryy22IEbQqPUIasXzKes5xk8TqnoG9Uw743gu/O7gtI9n8GsUR8LgPs+1RdR+V0zq91vg
1FsCMiGG+cTKROvedcn1nPTN6F+zwe82uQXHHymsLFpMoczajbgoFtpX4HuIEhqeyVyfx5UIhWOY
LKtq90eA5epmMSOnnMIpdGtdLq5ZV7wFjv3p1alXRntiaaI+LmwtWhE3n9fpr+TPkhaKProXQ/1u
2AVBhxbrp3YlMEU4nFdVuODdWH829Zhn60GATybOt9dCOYpsKGDpCNa0n01/qj0tewItNDMaeDvT
Zw29SuW/Ghgjjs7EcDhxEo/eVNj6Lt+wXAbHgeOFt7VheIWjnBw9nb984PqYbX/dh/7Dn9NCXZ5A
YoPCseElSpwLWNEP4fp6KdbNLVOgovqSuanN8rPi6b0UbzXSTxAyxwF+DSZJneMb8X6XUPc/S481
8CQjyLgJ2PwJBDl/A+GptqIusl9SIZacRdGNB23p/y0QWwvK/ADCvpkuCxrImncUjwrL+Wy+KqHC
26pguTv4f3RI9re5ugPSRYAAM4jr319ppnkRtgV9zG4SiLXi/SJd772ncrWRWJTqezKJxqlh7F49
u/3IwiqsjBW0pcIOXxGu+oKPy5u4KOTdZ++29Wm8UDp/+XdVlxaAEs7fKRwKHUQfGQhBsg5oaDjk
hRTh0xyK8LupyIN8Bi11eod+4CbqNvkSXpEoXqsqeI7hFyabd+eay/o4S+AzaUZrSjSmiofDn++p
JRDlpK0r74/k73rjfyVZ229TKB7QgR+j3vS28TfrtbOKrxjSRMwHzksBmiToxTqXKtzxG5KXsvOK
hZWu9YEKESicC8CLFmiTSKGF69bmcEw1TgykR2Y6rClnhCsCGnWmtOnD/oaUjVNhvxlAqc2Jn+1i
sl8rgY1kDnnaNYaUCnMOfs5QIm77aRjLBp/2Z18LDKBrwO9GsPJTFwWPste1u7Z1tUspaTnoN7ax
kXp3ZRXnIjGlmMsLpvITnlkOD62kTpc8bUl25XL0v8zvZBrGZU4SDJEIF/DcXNDnAqo9aPkUIyPs
/Dj0WjhvXxdaD16KwNT/zSpt/Lzukhz8Zdn8MqCOp11d/m0WC18iEMvOKKYCr56mPFtNWn0feqcf
hbPYnBc7ttcussUuXdCoHt2vJO0f7P4w7o+Fa80F3zOuOSDW3E2lNU9WQgYDzL07xsJwu8bCx2tb
d88Hio+c4bXxvREWRud973n9eZ/y+V4huiCacT/Gy/3thex3j5Pg79/3w8LwyO5h9bdt29zuf0zA
S0ltu8TKWdrNyVula+8MTl85h4bHYgZIP6k7ph5Xa6q4ZPBa+U1/0wBVYxhL97REDS7HnG9ErvCP
kt+QLtL4ixSvOYxHuiVFiiqnNZc9ydOFGptDx+1BqTKGj5GQBakcNBMiuDYHt6bSD3FubwR5iY8R
lJ+QN91IDHP6TJ6MFT65oSMvQz9X0h4eDvr6psfQcSiNArASz2gapjJzhAV1zTSC9AKrj4d8O26/
6NsXO2ECR0Lx+BIiSHEiEF6RlVIqS0DOBX48eckC/LKmFAYKn4ZcSHw+71bozjXZtEOq58PM8r26
PJZooT8FCcx3ZRpha7N2WKAX9j8wUmS64OdpSCIKfeqRWURuFM0Q6qOSm0tboj0f6f6jqbwgR0n0
18R1TMY3WhPtGaUJvKl1fLzn50Y3gn/et3PPLfCcNzW7LZncmr+nyGPGiAs+dh1l8iJpTm3SJ4M3
FRXjUplTla1EC4gHTyszyRUZCz0KCFDqi9sfX2fXg7lYjZ+Mp2S+9PGei81/H6bQvU2b7xLi/ZJ4
mp+xoSiYAzbmYBXsxZB3F3PdXqvsV47zqxfrvilQn4sk1po+E9rpmxML1+RaMesyINSl1xhtxxbF
2RI26HtpjVVXwQz0cPP278pvWTBCe27ugndNtS4uJSO4M7B6HHg8XtzCMB3+/f//P/PxqQDsj7u8
tXXMSXB6l+HPFbVL9SMMNBrYW4DK/On23uzS1bvah3iwGMWJcIElecoSxOpfWcVxTFCSqgQPnl8u
OfcgQdoALxHJCteiWMDeJSwedEj6fNJP5mkaopKmZIopdIXy3YDiAo9k0aU4IB0G7sL0xMkROyTk
STA5AkP9Js6p3v2djWtXQ8k0vIJDA3liXD0LHju6+3MAEtAbX45/IGe7xVI9xby1PSqH/4cPPPir
2R1zuubdvNrz0C0ZhDK2uAjyggt5ro6XkxNBfVFgqnmHmo2pWTNLdDEODZwxjQyOMz+INc1boVdv
1tG9sBAc/uFBVb/EaL79wJ5jPIzUMv9sRJK7bAqQYXgxC2quvHX3hp5+1cvB8oSfUGgYsAfeZNi2
VWClYiLSomp+lplyPi96useCPt3VNllWZdcFQLBCrFqpaY4km2VYS0/7PYhyZpH3yIiV7wd3d0hY
a39JaRxhzurrzBsUJTNWmvrI6kva8v1I8JyS0q9UovNiN1pERVIhs9QCg0SlS6nNzfTDAoi3P2MS
3ucWHodJ6eEW2VnFRdKSZiCuv1c/cLyUlWYwyFn+WhHGIuQofePiJ63qDPmnb+ZKCeR2IrMzdS2u
rIi3rdNa88yC8lqrmxGjTrihfFW5J8epsUVWFoXXa/MB9rXP1NHyeCwn+qQRSPuWJ8OaZXF7uPpZ
Yu8q2v8pWM7NnCATtJLjXgln4vhgLtXsyJw/dc9stX/GWxBQ6jIog7pKlW2WfvDb1DQW/TNiFa79
M6k5PHkFyxgGbG+fmyWKQZnTYmu5bt4sDfiNatigD0OhZ09tAtPNmRMUmCjGoqZvxQGTA5nTJE5P
GFV5mjcyPZwdEWvthmvVYjmG/I14Stp3/u1g3MGYkaUqc1aTPfRutLQNdcgFrNIupureh0mSvMnH
Aw0uMo+RKSvYxXrxeovgyAv3PsRYQ31ui06NpEsx3Nes3zUAQN25UTCf/ZFwEW0balL5x3U0gHpK
dPUBJdsNSU6WHPNw3qklzr5R58fHU9hVTPC+QGjqm7zTmCUpE1MGdxe+whh1ync9m7fKFCXAnvxn
5H8A4CqXyppEpZ2+/Qo9I+bDsI2OpK1BjnFOMV3SXQSBBcF0rSaZb5mvzdrvUII+YMgkM/a/5OP0
GgmU+iLEJbv2OwGv4SoUnhMFo6YPUynK55Flo+zoK1X89g7RTHAUw/MDZvdtxpmaiIdSRkDcMA/w
3d87cA6eHsUUkGYYgAaipe8rUTTozj6Bzo/fbux5QLFoiUCEEOtKhbc2d01T4DG8bBsPOavyS7GA
12FZeVlO/D4d96alD8tXdesOTn++RROFuI9Cfc1mrN29aARpNsJBX9rVGguJMi3zTyhMM4jUZZmd
o0kEHxXq4GI26yeqTbJ/OxonS1B2P8Q9dD3rkb0Iqt2WxCGSeeBTOGn7d3MQhMq28uUjq6nqHJ2i
k+hw+xhvKvFYMT/JTu3WIJfLMBi3wo1C35e1r8XKX1dAbcRK+YadjTqni4Sj/OcHYkuzmjg+YNuj
35Mufq4JE0m6B40pIXWtFhhULH6T3eW/AEF8tyJZKQm3f7a+fPZmr7UZoTMVj4PC55olh1mO9QFz
H9Ypw4T91RdMfPi/aPMaPNvYVJNcp13dYJra/nC63yKeBdH5fOGESUXKdhCiudByqOiXzR6E8yTA
deTfcNALKhwb4JEM5TrDohrHd69tC7UZevDozTNAe9Jd4T8rayHqcsDdV2lNJHRo+PwdcBLA+nFM
RmxR1XpNRs75PGhBSJbjY2migITccrv1M0nGyRgVHnQrQKNLpVU9HSOBHF5aTV85eJj1gvro/KT5
IqTMyFf1gK+07mN7qHIYoOrlba242gws1OZjjpu2Lch5w20TuLk8tLRT5buh/TAatwVEn4ucKLvV
fI4scP6wHwIKQc7sRAc/uLFV6aHFILOPeqvfFf6nbdFlmr4CqUJV8XdKKHTq6xE5PVviPbT5oT5/
tX28t9QzSVBZ3VeMxaB6Lv9RjhcxD1rtw39lg2BVm3TjvxU3k8qTIwfEN4fjKSHiCE7t/u735wez
EdSbR2joYlnmsaBprTVE+uRcW1DI4nK6/juIHGYMtwAT5n7hwjMt/ERrR3NFXCpuvGvewyo/guqn
/rhFg/YV7AkSAfs3ctk68tTzcr1e7GGf02Nf+xI30bVPKph13gA2gjRkthP3a6VZEth2Y6oEbwzO
wSt9yHF8h0fhxKqkvmgANw2okAMCNsb+TrNmuDzkCti6pZAd2SwKHUMVth1DBaahElXARCzVuutY
99+tfP+LDy/iyPyCM1CYLcfJygpj4Tcmy0IjZNtsWokZ5I0qHB3UPuV9YKcGsGa13g4oA4DtQw06
qaBzvzurCw9sEEHKOUMhy7schAl80T3sUD+rEwZVFzpD32sdHM9bk/MY44uDWdtUgEt2sG+7x7zR
YTypYpEzo7c2+t1OznESHHd8OO+hQltapfdYZYPhLKV2LapJ8QxX8lxsARZTciO2cc3JOeJrCb62
NM34062ZhDkHnHVzRHdSY1qN/SROCNTY/MRnmdlipDRWmn+AN990vix/FPVY7kVTr19KiR1nLzvP
Z+PwudMI4bRWM0Yto6+9nO6MrqA4CijdmsXMtF+bUe/9v6RPLDYjwGUlbKjU9sOblu5Ogm5pf5fM
I+OmgaDuX1npj7WuVFMva4fxKhbKLbVldRVC3nR+3EbeYY5jMoR/LKH4flXhT5XaCgZwDwnpDrf3
YEK24Zwqs4f7zIaIm48p/5SPLccGM8Uy8r1wQJvK5VexDBtvNt/PUfbaLWygos4jr1DQqsrsIrLa
VLRysDK2ejr6VidwilmC1lw3kS4Pqst1Ru3NWSwXfD1sqkJa1b+axtiw3hTzqLSh1C3LENdPR/km
f37brMVUpgLzjDHtmYOp4aN/MX12p19ar3yy27vZzL2FXJtMzRysbJ9v8Vq2eguUvGrHzxYUEVdQ
KFjJaNF8uDDx0hd0HVOpGgFlieRFJ97qRH4vbkxYPUQ5QZZgkXAW4GP32uD45pfEXs2LtymNOnV+
B1B50Rezmr607011jTAcqSPyJsRJHzL3kYw0SRPup83gUh7quUo9dUPj+7rlENsMCH7a7yUTWsCz
u7cnUXRCyq0d8fZl44zdGZGjoNhzaIHJO8UTDewpZPpTPqA3WQM44EUNUTC0aaenUOIY0RdEAbIr
7ZFe6JDXWazbPpOgCf4BtCQzav4Ano7RDqoGhxAZuwO28D4/BApRORU8XJ5GWE4CEj3yqtUxVQ8W
r9E+aTTWcbV5Of+j6zP/3LXFbdKxnPoLNPeffR5JmwAx9RaXF2tVBr6a8wA7/dERk/L+AqQKCydH
F0RDT1Gfi1OXiLs1WWAeTzZex5dNO2InhnSCjSMJykmAWPDTEtYUEOFmwA6Y9lsqSh/0NDG6TRO7
Sy2KkT3Sw3iuY3ZFB80mxmd2SwX4xq9d2ZfMRPFAjZLWYZBmX1/Zv2wZlPiopDJrWzQUCXlfcla/
JZXWRYzL0E7m8IMFqcN7AEyfLJAmoAubXBTSHOhIdnuZyrc8GNclmjYgshmHgbDEcDJT4PUlsNbL
I/baltkepPAYcB2QxPl1d1zdahzjGPAibzxU+wkmmpZLGL2BFZYIFmexyXC83mJxzWA/CN2o39wL
quj63Ri9jnqCEguWeIyziy1LBEQqGHXLJvGAmqFMjVvMHBLasl/KaHtlz4t5M3VrCLpZ1dY+mMAO
rrf8D/Rw1ZXe/K2CVGXJUIfjAoBZaBLYPhDfDhFNTyE2ZPiIcsu2viq26cgVPnCJstJ7UuTP2geN
z1Hq6bHPsr7u6l6PLSo7TtUgQQBtjq/E5L/+zJQ0eh92kyix32+px8orBjjoW1EpB6T3f3UfMrqR
c/1SAeJMYiVygkhX61LXg9TveiOuB48NtKNwE6NmAi8aMxFZvY8uByyjYS9ANPFJNUJGRKBp1UMA
sEmAqEWnm0/4Ne9BHgqCh5GMohcwTlWug4ZovsrnjE/t2ylRjWCv1WQcFi7TDUNQblii4fNT1u7P
Lt9ZO3oZNKvOcCG+FOevPyTCUmKN5Fe57efWCWu/BFauLEgfMda0A+XEBKHj2GEcFhDat/nb+nqO
+f+aMdIo1JRJbSCPL+j5sqf7dbVSI0VoppbjhWjPNT3tIc8YudxI0P0ruscvlrQuUbc83ofKVKJC
D69l6bcHZlk9ZRU/tsF3zZzHZUKOCUyqBZK/go9Cv9YF2XsuraQLx8Ftnh4hmLCvjaMekzRrUk5u
7/kO9V6XHEFM3/j+33hAt92RAvew9gVvYzhjfhfz7dv2Om21xHg+ZheIwLs7wVTo4LHPXJ4PaJ56
7tv3kYQIm5hTHtRMAE21U6H3/GJXorE1qzvyQLLqvFwG41/BXUyCRQf29ISdfUQJqgDr8iR/2GOS
89wXowsLuryh0miXmnOh0SSXLBH37kPoRAZcJV3m8Zlu1E9z65ZuSD881H7i0T3CpEJXX5LOfjtc
14QbvY+BWC8APY3FvB8jPZ3El69GgsICBfEJsi/ug+SMBOlNRZ+VVK1TPd4QuHT9qW2jSci8/RDy
qqxSR5PfWpmlXKoTMYS+YAii9cz2ghVIu7wfbTCncIt+sRFeBTpYMqDTFgu/YgmwBDsJD87UTOQx
K+2OvUmhMBPzk2zX+QxYBs6v9c5mKhsOBxrhevWh/zWS3BjS18zghatdQq8c99ATnQkhb3G9tf9s
X1XmCEfrfjykmg2G/ZfvG0omWc46Qc1lZ8dSojHgxMA99RToqeJwO1Evw/Bsb69tP96svjcIcHEX
fOhOsFQ1k5j5n5qVa+WdYjhzPPO+hp4G44pE4HvWnxumvga+Wxd6AVXIDOrzRj9VPXsyaBxhl2T2
EaC1gzK4d6Bc5sT6pjBfQgTVCP+M+XklUgMynDY5ezcLTkNpGPrE6hCSYbSFiwlsYwVNvdkacQAB
SJNfgvvQwvAiYIjkDS9seHMVWojAqar8v0CwP55FoFvRJEWNqTLI1kqgL64yufOZR5KL9aXX4uW/
UFGoHGoCF1bmX5oZ5L86aa+v2vMR6x6xZF8j9L5iS4xytvoR2I8TcdtbHQLZYCeXyLOJEFuR/3Dh
t1NnFaENs6vnk/FPTxE8MERdmMkAZjU8CvWa7rbi17kQt5wGrLUhqA9NoPr6z9KyNd1a/ZoAasDt
8BEU9fCRc6fCL6xEIUPzxcBjTpiw6dmCb7q1Wu5QaVAA2QlejxRKVCS1pv5fHpI8Uch55E6FWCZw
yaYDuVFDiKIgTVgrBv5WvFss3J4Tg9YURTqaiMTqH+iTIndGv6ErPUZ7F7jzPYz7ErRxbLxnvrqI
Q3qi7x9Nwlk0rSJqFd7Fg0WB7/8YrNgsrv5KRqsJOXb1bN4qzR/61zldOoswDQGpkFryp7xRGzMq
gfwIPtX3QtS3T0gR6phgtdT/s8C8HRSieccp2vMf6mTrSgYsb6Q1C5Z1463lTSPTQYLxKDV9tHcI
7sTcKIGe5QWc4s1RlKB9rA1Fus9qvQHbBfUVM93yPu2D4Ku4x6xQQt8HBC/7wogGcx9uGNzVqlGh
xdPI9vmyMgHMUj+lL0C1QB36G6IuaRLgGJZjk2Cnja3/crPoxXlCcfU8vOqPzzmWZHHOsZ/dj438
aUZfs8nKpUd+BldxI7Az65DCCT6kVcQTMi2gtDtb6Xneo8BZUqAvMN+FniBkHCTFkt/D0L4kgtX/
Jj2tZ8cvsE6YN68Uyh841sGBi9zyomXWPQWL29qkLkUnGJKztkcHy0SiH0IHkKLco3vdqXFQ31o+
eozcfENEMmYsjI/qlLc2xvzxGdbwzpIjKyB+7nhzzW9NKIoUWLtRp58rDedSjOzCGlsCyQA3nQw/
fL4dvWRsHZedXIu5nOOpIdqnE+sFrzCsqsUJAjJDkHB7w2HW6AkfBvVeaAwOJPMUYL48SbLS3SF6
sXTWjv8AdpbsZICObYAClN1myj++Z4UV7J/9MzX39EeqasHaTeJi/TWbCghYOa1Nysh2LpOyH79L
02qR7yLwJwEzECwdtYDyMkCHzvyfTuh+ucqeEAEPjWtpqnpM2UqznsfRJy6emfWNGt7tv5mZcFfy
8zEWrx4Nl6ySsx8GLjHvVizzbq7ubV+1XtN3UC9Y2HEZ9UqpV+09hJ60u/FCNsht+ZSsHRwXL4R9
aWEX0hoDcFDdMbpdORGvj8rC7Ucto2Qe6FbBsVnwq9CSk53el6ri7SIp5a6mY4Nb6W/FXpxGqjto
UtSE5xq+xwk0O5P/RJYBRWv5iTfRwYF4y3T5SbPw+IsH6uTcx6nCvsHENCcvNs7nmvUG2Xi/L4g4
8z2Jq9j6xn3Rzm2zo7TO+4BPWV1dwh6PyGOiCzF3ofRzZsu1iOLqDCCQHyj1C61X/wyXiuezX1Qg
A13CetJffb/jt2vn5K2fD8z846i48ulF+rrl96yi2Ss8kaHaMNFri0pFMy4mtBXkjzD/2ed7lKZp
bS+4yE44bhJUgaBuDTPDJrO0f3/CavuaKGoYCtU/NQzgNGbr/apt4jsdu0EVndu+96w+/KEwJ1Cu
ly0jXRxys/LDBVkXyILpWX1JqTCVQXUsf8Ykf7+9QkAb700omA4hbgZvixErc/5LNwKKPKE9e+8J
YFKKr2mVIf2lkmKbBy77aPpC62sRaVq/MG6ap8lFtQGe0fIiYwmRGh9m1gFl+Am0/OnSHVQnO/6M
hpMTHuNA4FmuTmBP3Hzofp0LKc+lIjEVjSMdCrnfutrV/p1Hm+MCxrb/gqMv/S2Qm5Q2X1bP7WgG
hDG+7BanTx6X2iEtZadqhnqvLVtg0zJvj11GvwmIIPUXNwM+WDAFzM85Z8HqsivNN7U11fHqKd4J
IPtFPbGBiqJeeW5Izm2RN3EISf4Rc2bqcgts2cRGUxaepfLkPelJ+jFtVot/tdYeayH4YhaDvWZJ
iGrm9W1qkdKBMxw++ITg6w41Z0e5k2zVEkwLz4c83vJh/riJcTIwc3EJGUqTyPXorw21jZgoM8lB
B4FvKZkvu/LfIe3c0o9ovOR7Aps7eWIm/MIu9u/mt35EBcmHFabxGy5TiaoKrkUPX0caAAd31zZQ
7WjKvPvMRfv39d5t7KR1iQeSaeevNN3Bo+2pFoCS3jBNl2LfHb3pjWaNqAgvCpbYhIF37v745H8F
05qSQ/t2s2hmCh44r69a/ZchNWSs4tyMLuAzrebsQv4aXKE6k27GYQhK8uph/HLUZQft35ckYJEs
m7fYNKVLRqZYoVrhQZw1AbWDftFRSCstQb6wUAn7pI9EaQSw2edkBhMWLBgT2LJUK07blTb9eyW9
hZFDSxgJOFMrnth63cKsHxn0BorJRg5TbzzhuapcbpoIKhB3gN88RAGiHe4oyVk4wzE5L3xafS0t
E9NgoEVQVbEhT9eKfDcr6Ojhqh/tk6aa9Fg+X1FNtm22N7mgqCG/8OuoEfupICIq4dPqvVz4ILDp
My9ZGybm4nvWxPmWCZFj9+jq6BzEIwXLvplXj4JckarhccrXaxsPkjCh31xYZKJV5Ni/QdcFu0RB
Kb1PXMgsA8848r2GbAbHJtWD1LTbRCyGbPAoK8C+kCHjLcks486thPIYNdqwozvlUx2smGFnLyo3
qNrzju+hgTJ3Eu0sp4ZJi3/TZwBpvXC5dBmaxOR650tgGJmgD89EcrtJfVAKePIjNQjvkd+o5011
44dHPDHffrd5OcycdmfpdNEIZ7M2b08K8SrKRGZumxiEQhR9mOxPHGh360cipUUmbz4SxoHVTYXL
Jc8eRivEG5spAUSD0D09FPep4c3KAG8OpYrQjWtP3cu0kpOXxHX0aF4JU14wnOI1M4KXfzFmu+OV
hBq6IOifS2R737inqiIYEbmEWBaabVpJ9XeBY8Gcbq4FDfhInb8dZ0hSSmKJSKV374IVRYPczFht
/FuqXrZZ8x0pXWupevbzuoPf5kJffnnuuwzIcrjdupLG2WR2MaarYlauBDuZVzM6sWfzXOWGAV6D
5Mcl45HGavf3owtjzfVAv1oYNfhHnU8pwAJxuDi7II2i6UdUVQhrR6SrOaGupiO9MmN1TSKoyV26
tZODuR1JCi7n9ptBHAu+j9cZ4iEtFzVfvbODRhLUFKrbgUl7ZxFAd7OmCp32FPD4Us6XUPtH1PZm
lomc6hNDqUQXvTtfvyBqJsY8rRWIzKNWvrLYt6Kqn8rJO5P7exsdYyVGxIfF8gyvKP9oTQcMtqdI
rP8wZ7Jqp+INnvK5ByFHbNPQXFnGcSxKcHM5j++WUOu28oRJ4OKhTA/CNi7f02uZ0/W088wFbwAO
e4sVV9M4LU8Vm9MCNZKlt7EcCcMKz0v0Md8ZakTJ/wAgjjBn4i9HrtmZ0KQJBBo2x4ceKSArIFEK
kzqLydPN8sXFjUibW7M8rwNXtTktjKBk4vc26eZcBsP8PHiQJ2xfRItR+/vzMtgKzBX9rSlNIMGc
SGAau+TJUBWWWe3KnrhXgfA/c+2/tSmmtFWN7H7ctsbR5/q4uYWxc2kc6LauEKBR51acmsS3pXr9
xRXpcpdljsNlhEye32UOH2o4bfaF9xQwH2dpxu8RCmjGrldZ77dRA+w6z69V+NKS5Ehj62Ef+a2Z
czGbQEVugGcLfF0prUUmoUsaigYqVkRnEkp7Xfdl0UMQQWfoWtF2oYtL/HRmbfqfuozOhbbdYm2w
3UAFiDIwzjdN0OeYFzn6vikTaufCwTOF3EvQtMCJVOIf0yfgc9s9ULMOScTbBwkktp2tJRpqUO6O
wYLevXckYtPjzscxvBx5B/ujYRSCM80UdLrfvxD/2oJ3dNFl2LwaJDDpClhKhY6i8nZCAMWoVKOc
1wPuovjeb2WBWrS5McD74jHDrqWxiC+1ARyCT6DAf1pHIpnAkahDNiWE/tnOkA6HPHrPV4lILuT0
KFGQ/7CyUei73Nx9Vm+DydLsQSxxRZ1FucJe6d5fwSWmCIWAnjt2cMc2+8ViHTOIbhbbvsM6nj5Y
ZSNR6pZXq74q+abKEvyOWz7+jkV0JdtSqtqsQzvP45V8mx5C9r4FUXS+M8Q4b3n0td65FYGQa0H/
B6Dukvp+x9YRHGWVbD7dnSdgQWXjGyzyacFRZzd5wBosmBRk4bBeKpUX4fozZVp7BLpbtLWBxCax
tHGv7idXmW9Fa+bQ1u11Op2ZlZ0qZnZgJQNAYFCO3YJhnFLEgATpBYHoOX6OUPtLknNL1i+ZaGEm
sh5WLrUHso0LKWjHewYWWW+xCzQlk7RkeKQJILcuYpx+/me4nJgGefSC80OYhLC4kL3WeZdiQHdU
cHmZflkuX7pE6B4avIVBMqjzRTgjdGGFvvnXKawfELV3+6hiTEMn4kCWb3HfdtYdYgEwJuvmDruk
VsUF9utBLizbesrsZBDErRX4Gf4UIG3h1uCasVB5iD2i7wq2eRsTjKvh8VMcVnk+NzXvolb0zqlT
QvaHNkNkkJjtlN3Ew6DvEudNL89H1myYolbn28p1CtzrsmFMDgQlesVAb5iw9QxO4t9iFamNDmuJ
Zz9A1CKCipsCMc+gvGnlkRQWMi8n3uhH5VswE4H+E66KE6cHYkzEJav72O+YTrJt4YfNZTXd6tNS
g2WdryasU1iviCg6nMykkXGnGHc6o+skuXt6q5Kkr4Nembajuoj3iflccsxzJMrHXiPz7t6/rww5
fKjh/NC6nCKo7bwwgbOWJ85+upSAPXepOZdZltvJdL+p0sv3UZSOfEHM+Qv2u5w+n8bVPWR9w9cC
r3cKmtLe7oSNOmPxmfz2JVCVoXBY/C8eVyVUDSuTcTkETG+QLJGieT6vX246aAKwSHwCMZxFtsGT
ZH26lng3b8VeED+msaTo+rvwgQIwNodGZaJHb4gB7/tSFw3VigZJ7iXhW/RAqVeynfO5QS7DxMAz
QV+FqQvkcAaa0gKdZTaG1Nry/8sCvTRu1UN8KCMwXwXcKSKg1YiMaIqnrnVWywVqE3L9e8sZRXYA
qNWDzCTH/xS8dB+p+hTKFYQLZ07kFPW2FK1jrF+7wEMHn8UGzXq9vpJgCZR1gGZ3zapHgydhUbEQ
fKBD2W49zPDff883SqT3DT8kd4Jgfmdk/MARU7JyI7vIgZZ320LpgIHHOStUmjluM99+Q+DxNEmA
HM5Encgq70/aptdE6vGzjdr8mfA3QYD+pZA/USGKkqJqDGWv6h5gV7FdYkdpiYiDPL8ExuXX2e3S
1/dLeBnvoYH3dD50pyhgW/A7qixH7N9+MKNgseOcoWWFPVPK8SB59MKZ2lOHudETFPsdVd6qQG/Z
YXneWBBb9nVA3ueHD8wxCDo3NUi3MTQUdOrQJeYgVrUSraqdJ75Uh1bXSLY1gjynpvbr5r7kz8Gp
tovZ1FlQZxFVCRdHsQ2JRuD41goD1oUH+OEwTxaycdVU0NCkENhObQDxn85vw/Tstl9SMKoJvcyJ
Mknz39ZcbVc0Z2/VogGRDwBR5nlo3VWCdlRonjfCKFdIeopDFLxHCGNSEtJpkmiQc5Ld75ddL022
qoSIu7FsfBNEaadJ6KOUwhSFpjb9/PnfCqBBGvfAf2Lj6YzIUnXLyDTh5QRyIQcV1+1cYR+1v/yX
umpCXNIagtQBdyLruIuQZHhLuEXMcMdniBhj1ralz+C4I36bNE+N2jbz2HTURPwawMFl0LWzn2OQ
4aDl8FF6W4D3Z2yyCvLNHxEt2xc1AMn6DDl3BPS1PJRTt8o4NNxZ+fT1CtUVfIracoFtGlK1Rc2G
Mn+uJRjRp9lu61tGYbot0YgYhxH/qQYCVkjvahTPLiQUhTb+/wosbXJlsHmPva5JYlS0g9htD61g
ebpd3eBMoFRLORyFI68E4L/J9E1F8I5nf1XKIxlw7cm7Xt4CqwSGHv0QrCpPOwV/aQuBn39Zh+5d
qV7o8gq4aKoBY7cLqZEADDnMn3KiSzTPbw4I6vPNrmWMyghdK5Mi05h2TX5vveCgYi1G1cvRy2Nb
CPwbNau1+IDaHYvM821kQZ1TsYo6ttKeUDmS67GmD1t6scjF0ZzUlWmR82wNGo0J2zqMeV5sGGBd
L/wmXEP9H2ACMA3KI/AEd+/n1o6IB7eYsFbzYhqynQF2lBAB1EQDOdOu7KJMgSJMNpuA1cr1ucI0
wON0UEVWCSqosfHctUwtGos86o8VOkfA7AIJX3mGexmGufBkpY/knrG68/K0nQ+kdtrUig2alKSw
phdaWrSOnloLnU8K5QaGmlorwlYtSpQLGix8WqdgMO7BajbDR2nLEHvSj1sgV9Oo+ylZpUzM3Ddg
zBDX3BpYjIdF9fpUCAfWHCqOWfBrfURg1i1vUSIEaWHXzIOcK7Qa/1kpvtN9+x0MHDhvgJXH/txg
8UK0NnMRaxkqdmQrcAyh2HsjKOJSfjJtPBnzCQ1NGokZ8VfC2aLlPVraPIz/50eyw9dybLqZWpaU
TbJ6WTrUWsFqgd2J6oYT8A3ZbYzlsrHUM2KSZ3JqAGf547nOczo9jf9pPTWyotdg/IKf6CK2cIam
2oIkoxIq+tX4RbvMjyuzoPcj3pG1aJbgUTrBJtWz2toQ4qq7JOkU108wKj5sUK1AR7ztv/w1nj4T
HeqPSyX8NpHuZUXw3vVfSFX1lu2nPNRI6Umuixfrt76YnKRPEcFRvPx8HzMQ8l77cefSUrEUvYBG
PaXCfOuMODHvPxsdapGFC+/rmXbyFRrIrQzAHZfS4WhPYiZWpzfzlPbB1EGJ7yDVLIm4kNV1Ix83
Wzx3aB3pyTzu3UZ/+EbHr0iSPE/UUj+2GI9b6OqPU2MgccRrNBzmdEDhHCUex4+vAWATqthCi6ND
4wFe46jvUHtWJyxma3nZqA9t33QSMw/LENrnrdy2kkqJdjF8wD0etrpT5vKpLOFvyxtEA8yL7X2G
/fBJ2CrC4jBF8GbJ7vPHT6KOp3MArs26pTFRShkihyNSJTCBw6+Nn9SGyWBomXUOCW2Ws5+ylgS6
Lqu3RyeLBFxuyNR1IKVxmvfKYTEKtRr+9LyB7hF3sWiPxrwFtTH+zDTM6uMZv2yV1uVQeImrlEU+
8IkG0Q9xruENDxuIKHY7Euj7RqsnLbB5mMhVX5WUyW5Y7wFG4oYR2dQiJVjx9RyfgOm26Ht0lUyV
Jmh0uFGJ9vORtzqU3fshCj7ig+w2jmAZCfCJWem/imNfaq2qAWuO9mPWt0o5fwkZAXY0UqtH30yK
Omhm6Wu2vVHKpi7KkfYRF9PbDs8XeyryUu8iyBLToSPfFgZWorwqksQKt33PwtV9g610aVu/Ab3c
RNHYGZUj2KjKVWk8lbLBGLgZJ/yo3ujFCqBNs0kUPWcBsqGL06XuVTKFen8mS3AdVQOJL+qKjRu9
uz8d6xUufEeU/rcqSsD+20GDQlWYz6rYFp7ODZA7YiIhtgiS24S/fdaXFlZ1X+P3+cy0ShfhChuj
VdTVTiR4mAq6syQ42MMXAvH+TInNbGf9AHylNosvnsHsO+T0KbJU38Ey8O2Bcs6VBy5ylaZlQlUu
h7YzVho+yyh3g4wdhWU4S85Sk8aUiE4AlOtxPu4t34YNt0R/wZUbo+QSf2YhP7VhDDPgx5g9Crsp
j1/my0iMSbaalcJUb3kIrxz/7tmiw3llEmfrLRZwOZc1i2ndZQ1EUr4mI5IETklwlHV+9pPskrh6
tzuaMTk0i0D1fnDc3pOw2tne84/We8u9sbwTYoQokGgHluJhiUL/1LyywmDHByKbh7ki9M7iwUkq
Bxq7eUhcDRQN7485BxHB7NCrp+l5vinhLbf//uthraIGPX41SEQSWCPSdpi179/3kOuoS4c/45/4
4U5fzUeGxvg9TBwXiY0CZGouP08koemmcwfeRnim1InIel6Siixe8WSikSVhTm2a41zHCUzynO3+
Caia293b/CDf/QuCEIVKlZClQdG0aZyHFD1E4qorjIAXfojUwMyBPwX5y7pgOmMEQE736awo4iDR
VvKJnIb1hZrqbxbgCjJSYvydCTwJV4XOhzm0XusOX9RtpvsxrSIe+ToPQHuLYGqV656GgvE3vAbf
0TqWmIJfmGZ6xEcOtFliwIgzx9SjOT838JnncaWkC7WoaXJXfFNtRgyethe7fBcIMDogEKFKlMaF
8cbfQzw9m1OffqmLTfxP65zoAGre5gnheyIR9FHeiGljQVLiBzFZLQxnyW7DaCQ3xSTOxUjiRdUE
4gD/P+uh/EZf1zsTTmfhuYBUZLiIiBh/dHD8Fy1OmR1ijGS9k+JJTQNOsaF3jxuFMfGnWxO3EZcC
Dhkav4fvY2mQy9Du/W6AlepfO0/vYgwsG2/0Gq2T321Xjg+IXxwQ2W7NTHAKj6LUH51XNF4MtZUu
cXesnkSFI6vuo5hdlZVZS+CPEMsQ0RwsQUhBsxkZNpMb1SRDBrQR9raVBddMshZwZ+7XsnZVfKzY
0Vo4WrAiuGQWKDdnE1ZngwnQL5NmlDEky2fwpJY1CDpxf78eQc1D3eAtzpeLzpaubLqtV5i+5mSK
aFdwiy9NvynjPQvYajYBP+wx2to48lbQ3HZa2I6ned7QkSYapD7EGIlDtRZpOnqPbjQqn33QinXK
DuOOodcwJAWLLjelTzS9Xpt+UIFGyadbmy2F3a2aHcioJ14OSIKYwAKZNycltYlu8TRgyFmGasMQ
hLp47qgD6HOzFBVRcDFFybJezmQnSAR+qNXzEMPvwhSNsPkadkUxnHEUKe7CLFtW6/+f/NMyjkhv
okqU0VhOA+p7+vPb8dD/xKy51sXV5J8iudyy0pfX4IMndTyyBmYwcOiFyfB1dtpwl/kVBwDVVd8g
eKEZwIz8fqxpXNjH94lcxkoOI2pHkxvGzR3GT0bH+bGFBW/2Hw/AP+LSBJ8aQLSODIWhWT2Iqw1G
XDUuw6yOwfwyNK1VtIVKp4ZDsoPRdxjjVzHpUQHuq9qmxmv1xTMB/hwsv49dsv9GZI6+0I7oOmeN
N7KtOrAPnB59nw3FGc2MJpjmkxo/CjlRn/SrsCUZD2ol3t7UhCedV88Pd4p/c1Z2r14Kh13FXQMY
DnSjZtyzHl0xQxOc2kfZ3q8T9/SVUGQsY4pluXTwH89pX543oMGxgfiQIgqD62yuM2YSPqwOqIcB
k2gtadplZqJ0Zg07HxDnNMFgXnkfgnG+rotjjZEDWRl/7BXzmmwdVVeSF/CYGQZlil9RmsA12gSp
AsV5KeSdwQZvPfUSjKvLbZZOVF61mtFxoOHkn8B/XjsuvU8DqkMm26P0KNBEah+Zj21WUr33T+Mg
mxrddbmhIaSkEiklpUjsv/zIbGsyN17BAK/P47aHNwFVY5bqwq6pxFDET7Tt+zV+yqp7O50iPxpn
ibqKCXNhRx/R5CST3XmspYhuwySdE2Z2cT1fqXYItw+lOz5XYOamia/MSng8MyyLIDY3wWOe6D0n
v9zKDXnFmTbwPlPSFNfd4p1sUnTl3YW+e352UzFDn7tkqSGVh3Z+6Y9Vq9d8KhSsLcyUq6sEZyAj
9W/J0H5dt3M/Wf56R+afOSahLJIJhYWXl+atwRsioDNb7BYcHoquqOmqblCc3eizHM2e3mrH1PW3
bXfieQIwWBSUm7ccgR1DtS2Z5T3mRWD/Bz7KNR8acrfQBGOyVa3B9sKbaHZudkSHAseAGXBbrz5m
7iae+RRWCHpiLGoHzgJQC1T25eenz5eCSFXse1mSHMWZtCJWijgWauh6aRJ6axRHnbqfbQVX6HEV
mzkEnPFF/UB2WJrxcJLv9lh8Fmk6XOvZgri+IgdXlU1jcbdluhf5dXp7yqtUjMis4mqENNWw0xki
vQbu4f244c7CvVWWhG/ONcBHNzwXT5GrmR6M2lX9LPLlHGeKdZe6m2sAMvAx+RGp+EdlEn5iiWCK
8Z/mThM9Y0AZamudKrf4DUdNvyqnlYZ3S4Dmj6GUOC//xBbQn9I71WnS6i7c7EVHVxSNKEIColA6
qiFDfd6AFnvy1lVMha5bQ3R07aqjJKmq5AQB4/cI8r7IbYQGJgfuxmneTiLRPj2fSNjipzMqUj+P
u3plepmwRSnSHg2MrrARS9QNL5KcwCPbxZce/lktlT9u46u/UiMO5lDCmQI+GCxVPjsLXC9eh0jz
8hTG1SGUuuZpscLt43yRmvKNLXIiKYsX702RvvfvVBIC80MviJKuTE5exAyWx2IXUuH1aEQvLcH8
eOwOsfh0Z5JA6dqoaWamQbQtGqvP3i30mgVSLV4BjUqK9X2LFErrm1iiHaF92gEUU6UpLV4QnmWF
CskZ2Rr8ItUhma+nRdq1Wig+C/ed4L/+xz3peve8umlohNKOyTZQ8j2dNZlnyykm8UypA6c8TBml
6WSl+zSZjhsRPTD4gr4IhpqW/guGJNO3aAZNPvLar3LdXd3pe1ef59O5ab6BNekeObIsJ4uJWyZa
BpwcRoTC38Sj6R1ukhh2LtfNnPPeBByWpong5X4wnBg1YSPCCv5ZgyzE1BsSvlbgSQyyZvyDB3i2
68iYacxuGlOW5+DMp0iCkW7tp+BrOT8heHTLYOjIsOCk+fg/mY3gXRpdqYWJ2NT6Jrbkd1GacXPB
MhAk1fDuHjgeOzwsZBUU5IfrbJyqGFhlPi4Fy7Ij2442JR9tk8n2NuuH8jrOvVv9kAfehoqtCjIk
H/V14y0vNlU1RLspxuR9UDi1dLpqRDzfg5Smm+DTnOuZrK2ApVsZdTsHPEwsKw9JHmi2ocsTCOrS
ziEkCDaiPlBQzpWV9BLG+2j6CkDUHBVFRvLl0puR8KqMgl6Y+G6rZ9vU/bOdTUJX4rAv6D2Z/OUz
sV4jRPZNJ7gumENDVAdYPVbCw4jiBCX2dJErCRjqjdCtq+s0E450SurVtQh8lXLgyV1r43q6faaz
KfMwkMYXXGBjdaUEaw/q/iRjUvA0qLEv/iobA4FCRBVLrUKBacgjneWMwRovqL55VqyRrh+dKWzl
AgBptOBY/w72n6t7nSiw8C8v509Q8poTt3xluw8V+vTI9mLawasbHgTVpu/i/alI6XRsKw8ZRbGD
UarHurOjDK2eLEpVyDEzq92IFTcaaQuAde/yMfG30irJKj9lysxp+20g4qwAZ1cn/daQ6SHOpH80
47eNrZ9BEQzE/TnPsJ5uuiTRoxydLf6r2/inmPhF2arAQlpFbfFda9+UqhDCViaNqeb9z7aDNJLR
xWQ0NangaJtloiMZsTWh3xBQpHKSqiM4HP0MXYg+E/fkGDBcWUrDe5ezZo27xh6mPX2KGsXm9L0o
x6orA4nlyhwdvJeKjSYDQLy2tFc2Wk9+piyj3YpiX7HSLeR/ZHdcgALLzKcssPfGQPjl+r2/cccV
HflVl9u7gvp36Eyo57yFUt/7HK1A/jN0rDbVILdHS35H/bvOwJGfjYytk3aPx2XBijhKnn+YRoj3
yzkfSmUENV37FxWFwgThcZSh/31GDYLle0BwgJ57oFXNvWAYQDdv4sPGTeBJhGSlX8OBvjdtINW/
uPUsbhoBOyWmthW5I8lqc8P7NylGIi5JfckLpgU4MZCWkojOUUEbNBIG1BoucuGrQbeO0NGYY72Z
4faHwZRZ5S8ir4+fK/zy7kdxxXU+6GotzRLu/lHlGRFRmnLpE+2g+emHWTi5QUSWS19jvd9pcdlc
EEHcEuXrsVJQXS7+AEvH+KOy9gZMW4P1ApAYsMSG+twyqUhOV4/EdIkzoU6Qfbk8dsC3ePu1MadB
gt4cXhGIfkiAN5BQXlAt+/F5M6DKjX1ye2N9MpxFiAxJZiwIv71oMj84ZbjIXEs3E8q6UU+0BdbH
T7uElOTSF10J3yKFsFa6+1idX4ww3BPclaVlzMgTfrmvGiMNRmzB1/iGJSKLlRzOBvcfTzxw08J3
dygcwYyvZlmnY3lt6rTTvsw0bhn1mXxhlJJaT/wG8kiXwwZCAp183KnqAzz5dPQlr7qYqyM7eK3M
Ee4J7NwkVND4Nmrjxs17gW/sT8ihwwHOu3yjpEn4zOqqkls19b2iKe4Fbo7EiIvAvtsPbbwu/hxt
/i2Lg70M5xzXKBJvQEx+Ol51s12gFOv2Jgo3YKhnuo97JYgkO7r+3Vd4VyOkTkk6ZcMuwp4ZKJJN
AWT7doZ9+PkrkSTAU1cTQ4kmAfOCsCJ8NbuMKkUW1k1NODxoZpA4Qw/RY9BbNoxIUBepc3BnhYfH
6ToReF3UtrO4geI9kX+GDOFg3PmJES1l52Q1X5fgd21FXh4XRT7UcLjNqpAwmCHdnOAbGfzkK2RH
Ih3W5T8GGDphOcat/CWP1WTRFNLW7t6fS1DYNbfyNoZ1UOMQPgDsE0eAnagWQoVSvu/bBbZRTzwZ
wjZeI6E15yuWD/WjE4Hx6XfHjlZc2+3Wy+RZyuwj3n392E5dxZ3Hcc6dA79o6e5gIuGc1Peo71D2
Otx1sfx6iWMIjLI20CO5OziyDHVvFaLL2FNdrhbp2u9MwqsBcIt2O48NG2NZHxkkCqu+lduA6aVQ
m/DeVdoBqk7gkK0WT8eYPOPo4+KCvQdGdYcBMaU5Myio3eUZU1IUdKqi37NSq1OYe6N8GKIn2Q9l
nZKs+cb0pKojLvkZJ4Fbxhw8uEGnwq2E7vS/xJTCz9uzVAgCKmNDNn2mqhWPGynpu1zsFnNH828e
TkfalUbmnYc/w5xCNEMKAS5tegs9aBKGBKXnDglYWMqDENkqW+74xz9oPRWxFRQ7f4b50lATwkSh
G5kMur7qc+lfZ9fYFcVr9vJuGoi9BRzb2o9P/URIaIdAk4YaNgNQxgSu9AV1/C2MiUozcbWRBVul
FcMtm+LX0ETMwliQrerXut/jiKVPPFkXRcDgLMvEf6izeS6NCkh3obGcukcg5ZSILaDtXEvnex2j
6t19c5PaxzeILb4LtKaQyiAekvEDtCbe9bTffOSviiWd4JPwLMHbm4EqeDcyPrQEaWOLyxO7pSRP
CtOrr59v0ppqUMkkXP5d5cqKrBlXaWmOOAFJYRNEyCkoNt6tgGuXKmj82ufQ8HtCyatQ3E3v6d5u
i1rclStVcDvSDNMVkCRbmtyBtRYj5v8rk3gyqRgVZtY2tTqKhoDu0L2HExBgHaiEcq7tJ6cbu00E
UpUcKURSDbLqMLuz8lTxkdWfS85cfhABwWNqzU8/FrG20jhV+O12ggrsyHNJYmoxBof17oKA7YdI
k+1KMr+eAeHnlSynHUBnb9fni5dOHw5h7hYRDYlo18pvLbN1eyYfCJz6/Teig4WHM5YAnpS7Cqnm
KkCaUL1AwYs/+JGw+oqrKeJ93t/ihPNAgxdNN84rPtOuNpm/ZfYC1YQKT4HwExBf3YlcRI4fRknA
rUlB7iYnpNqcLd491zSU1156CvipZFTH+AmGYtanuVOsCdB/DUOp8gO9KKJJ6nclJDu5g1Emd2dH
/Ux4/X8fvdnUyZKqSShfWgZ3fZu0dHKoKNTgF4ENqwQ00GxArQs5ulDo9thfrNe7jc+3NhzrnPrK
dRBiZofDDrTfM49GypPMVGZVksvuaLBRjLij4vtkbX3YCzmc5enihcCAhLpMqPsfvI4tNVwB0uQZ
cSHsg/gvBIqnepyOR9aQcih2P63zFAs+y4ZGU0KB/wO2PGIstktMco7JGwMEj3J7UlLW4hvqPo1C
gKYPqvMf/+gCFHBjUNzDB4b5rQfFIeYYdt2W/vPTRFUWphLh0jYcYIQXyKuKl1u964izLXAp8qMC
9mxsdBGYIlFwpaK4o9usdODXiPkhmchbVh/Bf9IZnYkxa6eadsdlgtWsav3CRjocKi9a3USpWMHJ
0sj5pEuNtPqQk3O5WGSpM2WH/Yro3bcXhFL9SLRhdd/Q0Frj1s43R3XNWdn2hiriBWYw9uWOYZNZ
2jlo71U0W9AsbZYDOTDyCKtIBLxo/pO8vW7PW827zJMBDa+TaBJ1ga7NPqp52XKklL+bx7Gur03H
fMXFJg9oFHbYvAup6F57BF7tAfrilCgva+czqi6plVI01B8Rp3iSF9iWj2dgmxMOVupMBAetj5fr
xfQiDKTEQ7cJk4wDu5zeqzJ964RsmdqTuUclW9vDWqrL+zPlccgzLruCEAwST+jmTOst3uk5Ia/t
alhoUe945pOD75XpdM2+itdA8kXSbD4psjIkb3NxmO18/3mSV85Y2+md3IPhf0D6QPvhd0sEul7v
+HbGccy91Uhl/GcPoJwysC1kWdEyqzT6o95gnuS6VEJPaXxwzJdc/TI4RTDdNoKBqDYy23zj7NNN
jy0WgkuZdrLr6Ce4IQ+3kcclKt0QCPmXvOZ29aX4X8x+KcCcp3cy6+jMQb8rXoewbpO3emk1eXcB
s3h/l2i0aDN+Vs7fat7W/8bJAfT4S/dAKx6usjjbaJt0lNwZkpwKPajt/puoeMI6JIcxwCMnItbU
wLQbWTqmPfcE2zOFIpAj7G+zDcC8It1zczzESQ07xoPh7ltsJlfxxKjOe/masAhu57/N3OyiJt9C
S2jmguOGcshPwt0QspN5D/rL/MN/FKmXZdXpmraIY5U3DldGCnhAh6NN9udUxLOASlGZKWin9QXW
ZvTy043LXFKVVW/YKcz3o2/pjI/9dr21BXBMONWnfqaJYKzK32tHMth0Y+Wv0KBgcUQoKEQ2xgvq
2FsZifLsyUxcDrFMP2GadHlW2QiH6bYC5PpLwflnPXcGbvZMqJ8LBTJUnTKtMbuzvxcxARv5c/P9
Ct0/6mtUNWrWG/mCzhx4cDj48nJXTKHXJ8kigQBS4SB+7qnMbpMn4H7AmA3jgeW0CeNq/psspk2G
BJISOpDiblaWsIaFFsk5kCE1sfmfWtC/r2tWdvdaplWplfDJ0SIlxAkiCW4nXcdE1NBOQtXA31Ts
mViF+jF6vIdBGxQVIHp7L0exvNqqCbsrQjpcr7wGmPoTjRMPwrg4L736YDE7uLc51PJOdmY4dWxR
5Z1b+8GvWXF9YIDnQE/4gAm94eHsVc/CVcbkechuxfHCXNdqJ5TWUjl9FQuTsEJPPIKMoqWWGzC7
7ejEhPpfpDCo1Cr1z/Gbo6uRXHITn42J4nL+Utpsd8gu0ngbtghVYMSKhfT5gPDMIY3UDiFqorB5
4Nq9dSUXE2RnfWOm9raI02znYXCaG5bPu5evgg+gncOspYf+NJyIV0L3CAG8G9rfbc17g0dbPvQh
/ubGUFUqWcBWrhj+yR9lL9hiHSRH+saWQOqOmzaxMNL/+VQPWO6W2JCYo2JXaoW9crORRWDu5Afn
SIVcSad6oJ2f2kBNuoMdycZ2GPtLVQQvsRRdjRXR+v5jZaNPEVLXMPCr8lsNLzylD/X6QZF0IKS9
r3AyLiWIVhBp0COhteUZKAFAClASJfcf6WiKQhmW8AF67xGNrgr1uqZl+9a5HIsbcscpmtgtwCTR
VRqWbGpyqBCIOuDP9TyDEHdiTWcSoKRs54U4AN0dkRZUKLIoINOWRP3lkQim5Paxhs0vROqwJL6C
eVnljxwH9UUGnJexBRD63oF5g1D58DZTJepKXP8FmU+PuLZbuexkEAF7Tup32WjMn7TulZnQXp/e
6mM7zg9wbyoAQVP5M0HvH9+4xXMK3PoVy4gSeiOQm2nNsCpFcJHY9Gj1ckAm7HF2HG7brht08+b3
z+O2Hnhe8jo0Ry8jua/MNmGcF5NJE6hI+o5J0t+yLRCALE2/DPdJzevzEmmp3YIRl1T6CIt5tN0j
7X9g4Xl4aIm+O0Dsl8eUZuRpVKjcivA1BSORQ2/UpFRglDjqsWPyeQ/6EU1ED/rNPnQuh0tXxJkm
7WMmgqdCYbuvh1oI2JiPgoa8bpuQPTe9e0M8HexktoNGeoJuw2vrXn/gSGxG7pRsICBAG1pXzoB2
NvJCMVQY7Dfj2xSY9YrZbOiYv4ELCo2YdKr/hCwbzj0DWr8HBUF+bsEa9jtjWGJlxZ3xxqCsT5Oj
RRzhAXmeE/B32x+jTXXEu1O+s2BqFMDa0w5Prh+L2fgjDS+yAzVl2M9nQc/8y5JibIjGfB6NVRkT
kJbvvPd+tM17tvJumarJRcOWpuPQvhpi63VR3yvA4bxGxKDV6Io1uq2ApLIvSF1Fl826ev3aoJ6Z
pLRbS55qv0qDNdjJck9Ylmc06j2TlE3NZnCYp9PR3tecxZbpPltun987xtFe9jU5Ijd/Pz77KDhA
kqcbORmgx5ki093DfR+o8ndw2iawqvSyaK2lLHi3kpEK38iQElkzBTuBoMwFfz1ml3oXjdt4yxri
KlEOjxwExZmIyZdf3QiPna6TxQs6zt0WYtomoFIpkNTNYXPEPGnag/yixwwDvy+sABKeZhik0zie
lfAquCDIn1WYItR4ZNRJxR4xBz0cJbLSCcR7A3VrViDLrrTzUkT1CElZQEqSupIK1QwmnVlBO43r
WEPpXM+hFNSJnInxi0Dnt6fZbRz+SJTLlafxB8JxBtUsL716Zbc8c+2YjE5QUy+bDaYXyh15V0Mk
jj6W/0HnEqyUuv/BztWEimp3U2GnH4egml/3wSv2YOmoQU/C/eoXEK2sUFeiAXmaQ3d819xHPu5K
5ZNv12d2/y00xvz7ADvSclSadG5qJ6W/Qqab7K6auxAZQF7dYfi0zJwltZGiUUdss5SAL6q2FmPi
ytZQ5xvMnVIg9r2W8XY1r7BePQEQ6KVkhn0AcReIpv287/UDuxp2sl0x0YzmnHTnRDjf+pQNKJ6L
WvkvToP6NFv/9Q+Efo6fmtpMcCDWipkAlSzMOVr1TzUOO2jEz3rPsjFm+PjWk3OfUV2rtaWPWIFx
/yTca9dpThMLRR+cwOr//T4F5ZQ1xctE6Ez/PprYXLa+CgdFuWZ8XSOuesuQSEZiH6B7rIfqb558
oVdAKpPQ6xwTQEOLXnEDGE08LJ5n9I6N6qZOI/peC6cQF178QhGOXMiSVr7r+cAiOk4gpCFIA6u6
IsSMgI90O/eOfuh7GIk2LNdMbDk4uJ3biXLdGuI4ME4kRdXzyB9V4Q1Jiku/reyZvCxPCmhPs+5l
qhCcrtZJkB+6Dj+L9gTPn+NeQhpvpPs+rSIdeuYZVqoLUx1OX1YLAvzgpmCxEDWkzg1jXEAtw7s+
sTDuS6oj/QsmDULJBnwa0tyO4AhYGXAK9jqtPReSOTmyRjd9YBU28Zr2Q80kmiZI2J3Rv6JH5Nlj
9s6LMgVZmENCyUpEckkVx8mtGhxbZtc58bCGCak2k7tm60AFElUHJVpDQG3tCrQd+D37dQ+XKXxN
klxXuZgUZQSqtTGa9SJjpQda/46DYXJYBms9qe0AhGWPmJ7WBr+pmTVsjt1zUaZAEtibTFD0dwVK
u7NA7Z6ibaR1VbUCfZgvShlPYdE/4mKwBT7pIVeUdDd/92LBpQNAV+WlrOvTo5QSSnxIfq4qUk/N
Xo1bCcUqRgj8kkWfuSLbWoiBUcQLWA7qyhDOksODRAfJB6JGhGiUKxXFCWPWjIxvQcqVSNM4LqLb
1HJcwIDYWdB8ryL8/gGGm2hQtRod4Rd3MBd90lTGSOBQMXMHbTe+npjm67PL3RVXRsAjjxm/Rvgd
OjA5AA8N6nZNetb728tdEH+ZKefQInLpqt6BrZsFUwsdUIPSKHb69ojGDkNCB23d8bM6SOvV2wHN
RZG6eloxrO5buyCsP2/DV38c+SAY0YUTimmil8TunASf9izCMVY/FqFtYwE6VPU2coEjT1PjDZDw
x2SbRncJeOHRyV1CxYAKk0J2f5T1Qr/eb3capicDBWN+dQgpW7UKkvwJLA9EGbMTrt5/Z3hA+maQ
HCCPnr7WCNtifNdF89StD/XjwU0ABgCNFpXB+f4bTS/ASdqPj1IWl33fngtTCGMzbl6WjBkqfdEP
AXxXfxp4dMuXHJ65qb/48j4BgMQnQOtMAc3a4+6nyzytAwQMUyrRP6vo/2rC5zwSVK75MxhtDFXA
3AH6vJjcI4bgEYRKMNWLlt8mhBUkULjfvHGevuhfGGBMHRo8gGu5WXo+GzKqJZGH3uFUqGw93qRd
bq5S2THQ0iOOpooH3zncl+HDkeI4361P1NtsEKbifWz0nDMVEI5/eFSoj0Co/qPMeHpArWj2K3Nv
/w1BlYoNPP2WqHrpehXWhXw0ZncMSoam1qXwkp/vhmZdet0kQelemqXE79IReu/4RjlWdU5HJne+
BANx+9yKd+rNG27obu68K0zzG8booUP/ZL0mtWEp6Y+kQ4Ny77L34Xty3/qqZA163ZJA/jgN5ms8
XXY6ki51AoHXtO1UYWI07HCVM3u9h3EdsSEKpo1AT/dM0DCWgCAkprnIljGnvafKgaESzBf4KaVY
C0Rg+79JR2T66VbB2OZYnWZbIs6LNYh5nG2o2K1/SaiRR6x02fCEZRxuwr4o0t+/0aNdPzIR6ZkK
8UE6rphVewc/wGe8EQHu0QpzGXcVfBKbCtsIlGBNGin7dz2bR2LpuwVXWcNDlSVl9sxLnX1nlSJm
pwXTI8OkJ58hjPjD2G5UxWeKaoihmIMOZoU17E9xxTtDAPUiHojP9F0Hhhv0Ew7v3kkM6jGAQKvl
lF7bgAR0N1i8wOtc3H1k6Vh6umQrUxklBaXJ1YzsDO5u4LhX1+ZlAiosSvu3+rWU/aS5nb81gdKz
4Yj/f7jcj/n3bgbpx4k1PHbQzTxV/TcNty9oCr+7bgF+XqW83EjGFLsbbzeckHsdzzzQ7n5y4mi/
Rh9NTXXlh92Me/D4HIWS1ZF4a/ZdL/E7JAYRBzYq+E1BiCUes/AHulYic/pGAi/N/sC+P2SZhEmp
wWd5cO9wiOzJUAftme0LBQi+qac5N8rZg9jjSRSElMqJMdG7b8j+eP7zGt8ARHEQM2nb7S0FcRWu
014GPVyPeuzklWbb+37LoKCLg7PyAwvpcFK/JiObWkX1nyKMvQ6it4TI4d7PHPeF/MsmTjCFaI8t
rRjquZvNgfuGzggK3QRfLAVFt4DPbwIyTUjk0wi2rt4SxG+PXJ2HnttKZifBTZPgL/POo8Tyj38g
ad/74IQf9NzVq/A8X2jEskSLXIphRwUPl1/ZJso1qy1ZhlG7cfQ8cV7UypQcEnVyFW1eLn4xaVOb
qtNDWsJDj1jEQgsSgYgcjJtrettgnhI+oaG7IkW/a0ZbWrPJc/YFdsIELag2IqkFrLz2h41ZswmJ
YuKcKEXyv+SF590vJm8gquOw2VmutyJ3sgtRF+TCuOIrKWfqFDVpUVOfAEkOBmMRbeENoHgrSjht
RNlVmiqT2wVbpdj9lL2QnpnHGxbS+TWxw4+3WM7ll3D5awGhgDAkeqcClok6pFgsm66Z5tHLUn0K
EAzL74RqE8pbirHni/2yh4A7L2xQ9do4H+wiiPg/Uh7VSYOg/eMr1zumzid3HJaJ9ZHd+n6z/uky
ub1s2pr/GVeaiC4PL3F+DcfxqwAY809bYQtD/QW+wVRPZ+I9edsvxMfo10K/p/yKhqMQCkJdRjdj
R6u8go9w5Po2mqmX0KbQEmBI34o0x0XTMn+3GAOkIo0Ve37Gnfg1dApMl28qo4z1499oHJ3/ueVx
d0nv91mvAHmtgUi+owlmwAP/jSEqnOpq+0AP5tUwt/j/W76LZCKe8+CSl193gL7uO90epGpmKwZM
PgiAU+LdooRU8SWbdfuD8ZbssxJKV3v2CITBz39sD9vz5Elx+n+/kIRFG0Po4mdKb1ZpJ6ZhNUjT
Wr43QuWQB2SK4I4DgsoMUu7w1zn0SiiM/dlLxy96uzflyKxbYlcRVtE+oNL8tHyAZTSRvvmUr084
3W4WGQxGJX9U4p/Bostdbq6o3bnfwp6UJqtqUT227kmY8CI5rIURfLRGXuN5jEAqiEDuM48S4VRh
DzViKQ61cpQNwtmxZEPHtg2Ej+lU8Av8GoTU5GhrOiTN3RNgDYuqBSNKnqcUW13l/lTnJgkjzbQr
sQFnZDQMj286mkxEuo+V0CNdrs3ccwie9bC9gm/q1UayfC2QKdtVFNF/k+L05rzLr5PJyienhe8o
O1ccWtg4kml4t8E5RQKgUwUJCYSfANZcfT4Oq0bzxDUEEZyRhm+AJv4+ARsIM4dL8WioD/ULGrGh
wYlRenTA/HIRgTHSdkDdDWtmKg00CC4LXjNEHeGqSKpvX6SsXe9W0jfP5Ln0Zr7TD9eHYiNCt12Y
i7+ZpZtqqfhHkdyiagz1+1X2t+MS0iVFKx2tnMmj+n3/U/R9qLtJpnC8RkoLjeV5A8yqVpu8K9xN
TavTaNLnk8OETI5aY5Ne4otQk3TcdvPO55HuKRUmrMzNoNTK5PjeQwhJdTTcNGu3nS2llWi6gzwv
WSmmByQ2rAVNhJpnCjzoNfog0sBRBVoRzuiqohsabgkV/5G2zJ/mL8lx56RdY6VSG+jveoLOokpv
B4ShW/HrZ99BMXxVg2UllGIU/ZaXqa6NLF8E3cjkxSgvQeLG3SRcVNboeJl04ktSmVTl/+qZABIX
A0stCXOA2cINUGYz5WfesOi2XaBInhOLn/CoNLjQ38XqFRp18pAEejpu4Is0kOqx4R9eL/iSGKhA
Ig/5SwEMYbQCAfACSBSgvyYQ5s7zJeA8aqMSQ2/G/5ocPDGbizfaem7yznql9MhcW5GmCHYfxSie
fwrfpG1v8oEDW5G96BHo8boOJPHBrz8RFbIEy4IeA73p26vgVMn1PSoRXIxVT7rAuC0soKW3Yq4/
S9o/7QLPB5cxi49f7FyXtzoVaRWRq8Nw/GmBbnqP9jNxc1lqp0BWtmwzW6/rVBqdLXr2mKlyVdCd
MZC2mnPaEr5T+8PhgtL7REF3FesTfICuWgnqHgmdPTDdaXUkAMfV63h+Kd/wln4sZ+k2t5k5u2bj
+Q0HMk5NWRTPbelzbqsLwWQC/BYSY+jA+MWd2x/ncRamjc4E/o+Z+QBdq4B6Vf0a3AhCPRh2NG0i
l4SSe/GGqkSad84SMR1AC6aEY7rqY/OXO/uxf2b7X48BslDL2bXhaQdIM75gUv+ZW9MjtPx5OlTd
d6e0n7lx6kSyrDaUoxpJwnBDWopoEC1byOWotVTBSTx6RHZ7F3zKpY26UzUaQkXjRoy8F84eLLkz
nMLJIghNm2Ht2ynNeloWB1AXjDsZ4JWu4MHxS0ZUSzeUN3qWhvkS69+5s99HfW/AW3tbaLANCHbo
glPtckXdEJqgkjWwSNulGvais1Nstx/lcTqjjEwsoB0BbvSJ5y4Y+XSrobEUd11YbOOKVcxJTu2/
p1931wOu2FYDYg/Dj9NVyt6/Gfx4B4A5NXvJ9r5JajJ/n2ZoIDEjFd6F9LbmSLN8UJWSjUHaG8qZ
BuejFcIQ/CH2T52JI86vyXtIQCOwtybKI4fV5bq+oivqAyIO2ZupX5X/KzmTNMSL5Q1hsl0uAa9h
SP0AUIZ+4xCFqMkUgvfj5N+08sGe2XRvUKDT0iFa5JxBte5k3SOA2nQBlXUNT6Fmu0V2mt7q1Nes
WJ5Y4LZBBxENxRHVws0oGj5KABDmnjidWquWTi5+I3+DFzEfKb+s3AgHBvaG1A6E7rjFJeaB4NVy
9BYSvNEQcrYHKeLrAu6NYc2gS0N+3FPEjB+f/yWHp5dMiuMFNmGyfI7H4QItRxIruOcn85/BPbz5
PlJYQoH0CVO/D+IWPHRCYvOc4Dm4twL9Xt0uarCfSfhAbhPIqmePOYXhCcbdfeSOPtPbwYrEkEDf
TWD6Pug7DDj+ikWYCu12j4Lnmnv+lLPBKzu8QUXYdPVZqlHSzVf8Z/Gyhxyop7IlMpmHL8VQJ1BU
dsXFknfojHomzagDyRHQDEQkT3i/7S0tnaLEOAsaOTuGGugUOo8yjfRs+Ykf7a0wuQpwE1I9JoFD
7Z7bJyiT5IdfF1yMoZJV731ZnuRXX+qBOBm9tl/Cf1HEkb7SHcIOtVAMrn0bon0ztsw8DU59p7Ho
GmSZUxGbL7XWcdUCE6Zj/KIufGqhguBKn5/BtSePeJbrjCe1RqwzW4MVopKUrEKOEYU/33h6D2Qx
UjkRROVKaVqK5MBzusahpoixeiAQWVP8ePgXC5IqNOoG4v6W8CTE6LINe0Q21/6p/LbmlKI+DtvZ
cWXlOWB+XAkbskDxKm80/hUN2ciFhAHMKZ+rP3p8kTwvsKS0fKr1jHkeTCD5MoiPExNr3nPPO01l
kUZ07lpMZECyVMqOK/c5vlssZiQbaw+eVT2+AVkbJJCkUEkihTkLyye9Fb03RAm9guT5OghBmGj9
zUvcACv2bEOvtaB6ZWMb8rsNmHo1wGqIckCUdBccBJ+5tOznACL4X6fX/jg/HcHm0ULEw4GPPTGn
QgK+R2u5tDCuYwjUmV6ei0B43TqA+gBeuNfcZtp5s4NlYknNcL0IrijxYZP7cEzAoBhToKUjwKHG
NdA5cME91xPeYksCGmVkfNdbUc6z8j+8hKEzcyT3L05eedbRcuhnYfyCIGLXtTsPbIkpntak0PtF
VdouE2e1dQdiNAeVXhcficofJuj4g73Ac+Nm0d0eSfVCokt3Nhj6M4og17cKGD2J5YnAkeaZs2y1
IzPpVvfFmUGbRzBMUj+qXNudpADAPUWvOc8X5hEBZO+fXVgB/NS7LazQM3ob5arEitpv/JHy33vj
TaJQwzQNfGiwehKppPJO+PHu4pNKAzEnCzYHZN9RgcHF1POh/BQko3wJ/GifgcMZYmpVlBR0ui0E
Rc93PlBnViXoo2rU1lvbx7AMaVmLQXxAB1owq2CfB0vcBWPlwIJg/hER1aRgJbsh0kWZUhfsEcpA
R/JLYmRxJPrRYtVVOKLWNq9wLV6r6+tuYQuotSvjd0gbYiCeXsITHhCxFLoECKW/JePl2rkABZPQ
unAF+IghV820eU1sOq3FB3St5Gm1vqY5PnaztTiCXYqcCyq2aiJxHzKRzym6aaPSvErDZfKRlaaF
x4hkb3QWoK2W3W4otGrqkLtHDb0fFw6YUn5Lr3Dd8gTim1CQ073ky2efW4Tc6ipKbMKt811EHOpO
Q0Dn8iYPV4/DoiKDwdcz+GqBYLF6SXhsccdbGX4/E1sWJPJPlOvGS2iC9pHoPW789L6HNK7gDYpE
Hvoo/oph4lhWZEHMxP0wCym79cToqKrUx4AgOAEJLUB7psGmKwJ7QN7tvPjlxbTHK+U+TzsjGF6c
MIIOHPMYwN2SqA/CIlPbv2sJ5fwmB+7Y8PBwbZFYveEv9LDZHl3CokBRGKM0bvoOBYGOd/x0h9mW
VyDU/gPKC3dRDM/RNqZd+ibp4wWP5QnaCX/jwYHuNmlj/UVB3e+ApwH7OkSg5KxSpnneXbwMPk5U
Imr71nBcQjLe8A6Qr2gRteTFSWFk6KVEdFtgvkze1ol8lTYqxR2mxXHim1iziuUI5GwDKUcmmubb
dHXuR1hWajgW8yDTqrTQTEkC5SzodB33ZaJBg7pSD8GiKrro/0gGlhkzgOMBYrzlnzk0t1pIumDY
3sB4IbeDXA30Ls+/g5krPwe8ysa42ZR+YOfUne9nrqX4on77t/MA54W0OABrXsHEkPK+rLN9fLjd
cl2iCe3i18N8KMfNEdMNW9uLyDR/8r6bGVaMtIXlxYnf9Atp3snxFlqGfHWppSnO/U64G519Q4k3
IQew/BZnHxH2x7zv2kPDBRGCIY3W26Iua7dM0UBJWabOXQCO9Q6jR7xfUzj5d6Bkpx1ZYuT+qkq1
C4WrA6p86v5XHxh9AkU1MsIn/+Q0ty/gU5S9JIkYwnAMdJHKl3zL3iVVGlYef4b51Kc8W7KdqQ1F
77XZIq8IwRbGDu3QCJ4C6Z2PMg9j8j7S1pw6zOlBAebkvLG3b9FBChPHJpLOJ2USMKCyNvFnINOK
A2y3Th0CtCINZheg1E6n68NVjU41Js3lYV2nhOkp73eFYnclxQ0/H1YXxukQKuPKKfbSddrE5yTg
J1vwoFIjekYo6+KgJOD9PNEDctNKGn+Tdo4VNBShp9VN7RiDyUQnfm3suizxrrP/qvWxhEzWQkrx
0b7Dtmx6R1Js+rFHBJB84ZxQr6HU+saUTsHkIMRaVY32GeffYxhIUL8aXQo2oNtaFc/QC5mLQgxL
lfelkQm9C4vYCOk2OQMAU5Bhrk4ehFWLwD5TEdfnW4zPP/JmIvfq6R9ip1Jp5/s+5TT/TjypWCNQ
qldQGmKAUkLwTc5AEiBs3diqQE4TKnI5G6cwqajF07fFYUOowfgHk7Yo5d3TM04DqaaiXhaRRG3Q
W+WjXB4Ei1wZF6Z0ZIammZYPiB0SAAHbe6r3/qVs2zRxLLSdY7SglAGlRDPkvBQ8cTyGnorT9uu7
qfhPjBADXJzEZk5OUQsJdwva9iSP9EM7VHlrjg6rKu47LxAZ2GGapdwdnD7GA/T2yPsovyxhe7qw
fOvPAbFEwW+noac9hcwVzSHW3VE4UVISejeNQSv50sFUBayiV2ZGfkupBErJxa5WrspLuGZRx6UQ
6/aGYqNg0P/sc9V6BobTC2RCiO4egOEDB1ZeS6hTocn+fJbEX6PoCzK1auBI5ehBofv3yadu8k1l
68jCPHwO69t5tH6DBJ8P7y7Lir8GugWpHq3kYa/UwQHKZZjPqtm4r1RKEtTfnXaCs/0qUqZ3AOIQ
OWYSWY/AGVuMBbWQmzdXlE2EamX2/riLgwqsDBVxXgwUDGx96InLcgB34qK+CyQVN0PwnUwBpocy
ldLURBZ/KlpZB3TTkUy0YyHbc5r6X4caAVdqxB3TisHkRkkw5gPNX98QcV49csE2FhJjeRlyj0O+
PheiPowitL9bqB1SJe5cO1dNwsfbgp9QJ86g5Q1SCpohLqkR5tIn6IaCUYFNXos8WdxAG/Ul8Qoc
5R4jL9QL/+MvgXiYP+M2sVmnDZ8y98jeXfvU1TSqY1UVhHBChFzrUJ47f9GQVnuG6tIAzcsBx9B9
VLIMstYpEyclHAhD0XSkZHN3ISnUZhNeWYuY7KPQgXiGX0jG3XQ0Rb5W2Z7pbkOY0tBN1O56V7Z5
8LC3I+Jkp8188F5RR6ho/d4Ic8pzxsH2udRRoxAwfEorj0vAYKtFrAuZpAXlWmikp4Fn6iZrgHln
EGwm6eiv5+W6+KJljXRI6dxqluh1xmZzhLOD95P79uGy0ElWn5mWLTQ4uJ1pCZCU+D+3TEXpkEWh
m9WjaiIiOdpCiKMjX5g9a8BgvflK+kLuwpAcvR3Zqs9v1EOeTKAG7sGR2HyZLWiOSHsbAJin5Oif
JEnhx6VSEFEqZ2r7UpObP234QlWksNHAep18PEorPt+v4KMCZKhgsaLNlEhlRCwQuNCgmA/Dg8O0
N0eTNlFtjNSi2OP0c1fPGwzPMvlllSjmhXPOvqiJjd8CzxsqGSvplyY49KMJQv9ryts5usXZ6NVj
8hDwPiOBo6n1Lf8UTaa6fbuI8vELPTU/s7ss8vv+DrCjo0FYfA2QTh01yjBw51nV0D6a69RH15D7
oPjGY0m9Z45eYSttcl6kYLMCNmduKvsZzCxgTcTfJi6hyPhjJoeq+HkWIg2/AC0SZiNZae6XHTYl
SKSQn+DgMjk9MhbeOBDbATWTwhDEyjPnuwjTtk93JRFGH8X7TxnMmOdRGo2BDToyMVDK/AVVNPrq
AT0z95tSLclLVQzPvuQLrVPMECkyduj9bv0Fu7QeXFZvgHENtRnclOTZp/4R+iqQqxnhbOB6nTfY
4IBbiY+yWc97TA+BKstR3IcP9bbtFoh1eW7PzMVnU7LByR+lEpxbDMV537BdJdHnJFMP9Ky6+K/q
uI5zz5slL2SYRYuYH2WkK9aPMsQ1m6L4QwvzlIXVjlYFIADeqY8ctllkaave0+cwR3RkKX1YMK1F
K8g5c7omBvFYbXJHzG81qAhGMeSYL57fwJgCDd4YcYX94wHmvYHsBClBfrdFEuRuJS++4kfvARBz
WG/92wvKMOBztldJ2dUxeB+vDyrI7MLYiYI/CrcxnyX+Hu+eaoYKHMWg4DnukZGnTFpffmftDUbL
nuLEx2pK6DUtPweB9Jz7IETWrDz6ND4s7wrIoMerj+1KDIWwo6FkzfCymLt6MSl/pfQ9uTz2NWsm
fWZaTp4bg/ZTuOihrs0vcRp2Ude4DajBCxjd/mXAHUJekFy+wbHmK3ZZwCUObU+yy87TzaB3GKWs
vWPg+FKyZChQHsWLDdZ6VSp0IV8bu9hRtANigJ9KOKCREc92vwvBAR1SF1iW5rOaAs2ETx1oNIGq
9ml1sKyXbBftO1d8+ehrodnSUyBfxslbqNwJqnrrh9U1ehzGQf37IG4nWmv1xuAsyCLDQ2iEKe4Z
bvz4NDdBRFCT4/jwb+AF7JX534hJljEd3Dj/IX1/cFeZaAoGoULL0LkRgeWEtKrs4yLSZZKvFD4N
3pPN2sIPIIEFAWfFrYJBANfoQJ/GqEOUGhqDTiSzrDGtz4uUNfGUN6UAbnS0tTF9SxM/ftYGx+dJ
QGQQaTERvJ00cnhPVZnsv4N/0QvwRJKKC19o0XtcMgSTfWET2TLqT/JzDXoJbpUfXVcNXrAeS+2x
DGDlelJUKlkejKFwx24zL3HIFYKhH6J3s6I1Rg/savSXc2fUo4tCqOjpvO9H2I6KXuYzsRbTDYaO
hmUyVb5IRK79GxNSDdz0f/Rmv+UTFKlYvuUsjPjfASyKKXvEI0kZNhziPAZuRNMonCrOb/YGfDXq
EJkdR/33ryAXt1Zpvg7Rt2+TperKvZXaDKxq3Eo07yW5vFf8Nay5cQVCDTI59EbEonhQ66KcyNl/
Y9uiSg12kgeUseYp585udC1MZLXzpqSl6/ncYs7c6HNz56x17rC5Nq5dbmZPTLTmIqDtKu5d54Kv
kJeq4pw5jBM8U2QFViblkRFkWJ2dHbfeY+BOLP3WZ+fiwki5qjLAt2u1jTIb9u316mh0MKm6/q+/
3JGzjU+kOM6vk/pHVooKTKJzkDoMEx6UBkRkGKa/6OgjJMoqN1wNsbbEYtoyV1bfqMwFE9ELpixi
ovdScO9QpBQrl3LfMwj5kde2zGiEoHF77m5PlR7vfmO19o0Phu9CMe1jLlOOTUsnEGG50X89bBKi
HZlAkiFvVF5ezBZpAL+Ry9JCtx5LCZja4aGFX+RIiImzonQUzuDGmwaqEtT4BNq749cV8zEeE0i6
PDoXQfv4os9+D0+M/tY64DiYTbt28KWeSzdsdPcJ/G3XKSla5MGUeiT7sqzKu0//DklEO7hOOf4g
anXjjcY4F0LXiQJAaNGqOJaGpEaEgNGExcneg4u7k4B6wNGOlifWN3y6YUx+zLv/zS/mGaVTeIRd
2hnXcd7MVV0AE9RW+M1ckJAyk64Z1pFGzs5sz5JOYuwlUZGx5rnXDILHmYy/HZ23cftvJ6G7tMtj
onZCLUVjZ2yJI4oefFa9i+gb5QFsnxUMdNb/yD3J1HQvEvQ0dyge1jPWeJxio/1OSNGtcx0bKpgm
muRXTZ/wnca1zb2G7GPBrxFg4QKA5huV9gxBAmGhoQ87isJrkkx0u8E9OOWe8SDYNJpwzaDr/GbR
+noGd6AHPfRVgpSV8C5zuGVKKfneZCAECLuRb2r6IaAJaaqBbH5yPsJij8MAgXVycdCvd33+o7PB
fILxkx/punuEYOcyAuAacvt0lgCpHOEPLWdWXS0qhDeHzCXADSHO6k0x59Cp79f9s5tXwgbu+i5X
LUmkFoARAbOcs4C0YfHaJa39hvlwg+rFrrDFiX3vojqF/qF8SlD30hJTwUzFdXAu7L+y/ZttJK01
uP0+WYTCxDGpjzSHFhPDTx0GB9EMZgCH0alOCd6YkNBYg/aVJvn3ivCDWdQ07NKlPQuk8yRp0Q8T
U6Tq3BoA1iGuCO9hPYRHJpgIVcarWwuqygQAGtUN9GumybOh2P5XbrhA95Lr6B5EGL/x4/xr/YmJ
MT0CEZ8VlsWem2ao5y4tu4ibR870aWb5XEIP7j1/cLumBeNRrIbUfd0qSExhUVDk9PQRxodkTs85
mu5fE+uwnbGrbsZ28/49dmedRA/LdLcW3BKQfOcJYSftL5bPWLKhHPPFuLjli2T1PTrLrFbefcSB
Idp7tvje9s3LeGJTvUWTgd4VfC4yFs6jKTB9zRsrj3ZbQjoaGuehE9oJuLh6sNxFLyloQTB+AdHk
pSPM6iIYQVHFOvVIdFBxKZnTFsBd3XjvpQeozZK6Y0ft70TasaJ9yulyI8oeAPnrxE4CSKKdj4e7
EiHzkct99CmxuvrSsJCwKk9J5QDRk8SKKD7xqqvfWonWg8XMFOMat3d7pezkKViOfj+y016D42wV
dABIItkQYBOShN3nc3GWiGpz2BKP8IU6sg7t+FkUb7TXcx14fZ+snxt8ATj4BavKe1RKDsnfNkaY
tQlZy+xg9jBVPXk3q5lg1yT937f2nJbLbuKMYxSgjyJ6alMH3BI1EyR0nSe5r0Ow+/oifA/HybnP
ugJrNBeo7lQqYjA7T8xz9DVc95C/dDoqYraKjTVLu9vrk5zfscfenZy+Q20VMRCQN7UgDlmb0D3e
lu4e6KbBRqjY54zmLsBNAeweAs9IXLLdSnk1yeUs1LpQ+yUuW77mgODgkeVFiKmbxegvUGMNfY1H
5+DI7ZZzjcapjK5fh3ZOJkte6qZ0ATw9ZhnVBQ9S2tilwoQOO2QM7HjwS8S1l5B8Q2eDmlWbZlgL
mkg2rneRGUUIZtyc446HdXME/aZ7iBj0yz7NmU4SB0QdXjHzAgWJXAqjWqW5V9Z0MDbOn+WkDuoe
3ANn67yfa4wdwjs/UtRrMciuCoWynHB0KlOsro8UnF4NZCxk6ERZXR4toWKdJDu9fOjno7sA26nR
8txwe+dmtPLjdXV8sfkNdk5Yz1/9QugEwrRi7ZHNbVMyuC4/25s7qpsStW8CpUR3pNxs7yOR+Bg0
j0V0yteiHbeXSPz2CLkqB8UdVRV8Ic5hgNE45H0/y4ne4c3pAc/gJpmfTDVtUtN4LNBi9VWI2bqV
Miq+oP9mGz2MMtwL33piN2Ay0xhjJOIk9/EZwQhPBoVXdo3FY/pjetyUxdVTM5ogOsfhtouS7rvf
z8EUFvBV1tY4UZD8NWSYk5vKJBqNibfIFKmMthm3U3zGjB/aY5t5scF+3j6rSlHR8odu8f55TMqf
6TzQOPcuZy2rw/tbC6mdy13MCBXEa7/Odye0urNpJ4OMyb8cA+q6msPKz/1Mhvwg5h3SL4TFjSG2
2SAIun6aLVv6hVDk2XQGetgyTBhk8FLqjq8yC0JT/V71uLweXvbqvk85r8JSeF5nvpbkoqLRXofP
EkQU+2b/EAGipxZDOPICjIv0b1HUHkMNzvG8ENePrjUXR/U4fKaRix8Lxcq3BsvlFMy7qVY3T2nR
hby26LKg49/37uPiw1FrUWf/U4eDNGWBHPiOCsHA3KlcaaJS4cebiIneSKtEOEAAizOn4zbT3uh0
LWFv0yMdI4TLcYAT330MhJCqgED5QzYRTpHph5zYB4WP9vkSlZTIEQz9tNXlpWJzVcX0BuxJMeiO
7jsP8dQLvtsbVwlZudabS5X0CGlWJk9aLW/Q40wk/lmTdcy6F+sERulHi1jvR1Pxf56lKtPIKM/C
oCkX6JZHOlWFp2MdEH/2LGORNuiQc5ht8bcNi94OysUawVIVjNOgekn/QqNQ6rfUx0OhlyfG0Sws
3xHZhSCRRTPDhbwsGA/d4oJvTJJ7AQKWe6qSYcOaAy9wx33cqeWaEG16B/CsdXCoSPZhobqWS+QB
X96/HzLf0Ahlkc9ARVk1pNYESUUZFOpewqWYFzgog70iF2LWQTPz+PDXcKjbHR3IHUT8JtvwbHEv
PHe9z/xDH2RXWmJELFBdnkia2mbemzw9RDempNp6iVtzAgeBzaGX6Cy387+y0g5v6/zSuLw0zRoZ
0iO2A7q5GI35+ukjT1LejUBftmqILGaf0zihy/e2+ZJWTi8CaR7iz0zAEnYfbATTJWTMBMkgHv3w
SIm2FQRC0/etMmlAuyBwAX7F8l8WgNQHbeCW/olkK2Zv+iNBgnDk0EN0JlcpJ6S9lCxIGT0MIA55
XchPw5IXf0Adx/70/o/L/DZ3pK1+dqbEqY9euj8XwFjaZ8duI0HsvhE0gnuNOZKvTD6f/JCqyldK
qZNJ9QzNBQggNVoBuOXOQBUYudYMcIouAs/DSd2qOyltK88A+qmsduRuo9xTxm0M74j+iL1NIcEN
+6ph+skE9nUvEGuDeQEs4m+YZmsZ5iVaLkVE08mdFkRWH9ZhZhgbZf/hCQwqcg1m1csCuzyU2vLc
VH22Wcwtu419cdWnnfF3TyVKdTR3gFostT0xFDA4zT3G6dzDBRaVCLCL/Ojbe//e9gP+Ie/M0Owc
TdlJcXLoZcBn5CqU8yyCv6iexW1UCaPefWsGlR0F/Rth4Z4RxwGKP1YcZXOGQZrQifc1qEOgry1x
7p0tnCEiAxna059ED7YrYOZGnd6bi5kiOVMzMw061wGYpQrwUtX4WLFUeIGDq2BxC7ScCDtz+TpD
zZLC5SYpKMRcdD6fjV3EMHGGv9xZ7hFzhee46cJE3H7cb5U8Fy+Vx+Oxrlk1z+XcXO4boL2LmlfH
9BTqAkX4aCCrnApMaLgxBiVkLbuLAkyVOS95AEy3KY69joZQCe4/KhKLDbJKwZ9fjgqSSnV9Z7F7
h6mXrdWXOc8APOmHXwFudOISG5UR9M/89dvTcL0Jcewc9KELPa2EOXhIGbej9pfEIaP8xNA/PA5l
AFoMWCJ40cTnxgRTA46bxGWbx7nz412X8vpEJt6/lAlvt2ZCAODAXSSw1YdoEELsfMJ1dRVbXj21
To/I5NUb1+z4yuwBWvZZegHMV0a58vWCahYr0/SP91nW36RQP76GFDKqm4IyT6aPhvjND57IC6kO
eFT7v++gq/v8/Ut0AH1WagXprKnfWndT8XxJn9EJxWOlZmXQKBZqnyI1XjH50jSqm4xsaHE2L3if
bPpVYmN4pQ1Mhh8m4YsaI9/LhL3Wj5SG0U3j2Q8lMeX9Af781b0j//4FHE2/sZU+HoF8FDmWWZlU
2UBo2cQ37fhgJlGip/gZhPC5TwY1W75HPqJwfMPv5fXv0r5v7suEt9G90XflJcoWQRCuj/6P1Yd/
dC0CbQIhJl0eFzC5Jy89j/NlHiKSj0+QD74aWGN+xFPhq8g4t8H+kBTHbgQNmlIfuVq1XKmHyJtd
nTwLRqijcWu+vingxoxRf9wWSWUDQWMswfiQxbjox/Unq5csIt7IsVz+rUqs2NvfB3syx7jifVbT
FLzLw/wn11IPzhfRX2bTvp2ZNNz9leLTMfEH1LL5CayyBs4Z7MDrJGw/DqgbEHUS3aVgUTUCPIRt
WbaGz74iUWcf0pSdlWM0ZDEPCIHoFaZmauzurNln2XdGGMB7XvABnQxShvT5/FOkKn5zKAIIUYHM
6QO8R2RaDmqX2J823xHLqAv/BRgmYbyKbKzVy2C3nOSC8+6S0JNHN1XJifHf4E7DDX9yMI19zEgT
lsKBG+rwumhCXlIuiCKAEdYGZ7MZidEhuFFAAxSNT3a2Yg6/nU9X8DvSBWHjDuSeBwr/0VXiv/Nw
Wpn15qtV4mMUQoL2cttXaVYIZShhx8cp7PYH8ZmOm5ZCgRRyd+NKjYUzIMrqRorgfzpjckl0QNAk
FWNkGqLBXG+11joF4uQ6Y58BRaF4t2yUd+UpxqkI3FVE8719oEo7OBLS85WwaDGqDg+R0mDHPkCe
Uq5RTUo6BGliSEv49xSlV0xP5yc+z2IgzEVpQt1MMuE64A/YhSENt3HwERjskIlECb36mpgNydVC
BEwhlUyuS/m7wbBxmO2CKhZgTeh2I2xoZnNavoWxa87szcPKj0jgnI3oJM4aKXLTyAClRfVbKDXG
bV0iSK9wZApKlgzE0PBZbhbAG3maNskzUxULiVHJ3kD6Q9AS35TPrCOGl5GAKY7GjebqOvGc2ajY
AQElH4Vp2BFQeshIsJuT0nMJaRmDyUVUfcFDrR+IIoUoSjZrhaoVDlIOJfHKaePReAK4t1stGfRO
T9tBZWWYph4Y5RQxlVl+miP08Tu8CZLiMY42PC9Yc8MluPbh7MIwvKNLUOQw6qz49LORQumc+XO3
fGBuYCJ/qoggXKkSDRso6f+e5JGn4qo74VJkGt9MK1gmpFyVGYShflKo1iRumEznY+SLHAO0lEdX
R2zCyLrlHicnY5CjND3BWikjUa/XhycN9W4XGvGUMLEAnw3MjTCzgATryx7OA9+9iDdRqnvmE1CF
hSMeFCB543jpcFkkLtwqCDpRULiaVdG1DWjxXfZkUywuku75DaHUaJI68tVYRlDPGZrJQQ0+cZ/g
DhvOHAgLW5PXAFxvQ4qeVIDGoyawzIm0NwwGRqhBy0AyHIfcBPtRiJ0MQGSwRMPKvxtfjnTywqL7
AKU37Kmj8lzjykQdTPldeokRmZsPvGw3OEMqCO77jdiEgf/6opJbsWejZlpjx1uBDa8LdP6BL+Cd
SCV2IAKLtVFVf9ZAY86MCXwhlnUanbs+2e4WX9LuQRdQ7NAkZS+cZwHjM8a+tWicS+oG05KOdt/Q
Agl/w1mH7jPZGgfOQN1Oy1GiRyGfDKfO0VqVR/6kTyBscVqHpAiFwa0wOoC8SrcBkzzfyJq2PwVC
oHQgfJ9jS2q+vu0PQGLfMbDp4F9w5OPlKav9/bSo2ct1y+BpXOLbsLiaK3xL4EA58H1mlv/SetDF
B4C+V0K74e2j71MCMExfoLPW+/1rneh6tImmiWkNO1r1lJV+X5NAoHIRuaFhYqSr/yhlkGVTwHCu
QtCzVG1C+xnxnoC1f3itz7ihIiUxBnZfAuWx0rfs64zv+lpI8eqVCZikI55jWgvN8T5scSm6cqYw
ZnvlJC/Jebkva7DmvyFvFv9Cgarv8SMBL3a4xR7/7zFV+nJ04KiF5jGd9HxliIy7MZVt1olcQrYE
6OPcSnF/eI5r1S/ZbjUuXx/mbJBvfHlbs6IR5nnu9HeMee0YFNNYbBUDD3faWXmmGLPyjLRpV3I5
3oHaUbEGDQVFKu2VbquygIByuNvctJyJUVapufxM0ohn38fD1sxGZsMmVOgyB2WSfzd9oEKzJrea
rfMcMnXIUnEsy5F5TJ6M1rksLIhQJmhaf6Ur3Od1ajaUNQEGf76I93nbMX4g0dourJg5OPz5kZTM
pcGwShOAbCIZYqc8F9u6/YDvHwFcnsj3yhbxxwLfGyU/EeTOn6dIPpppqyF3AeAcgV3SD1GOy6H5
b/MUZeoGgVnMYhLUXdE+4y3VA1l8eU7YS96DMAB+a0ZjBWb0vY3qcLFNvp3eYxuIv9uFsQE+xSey
1ZhLNoSwtxbnKwq1MOtNX98XXa8a3N2IiGKw5noXzzVZmBHLef8+fcZqdkf9sFi+Xp00aQr8FQ5G
d202mOq5K8zJkTWVDxBSrS5/G0dat9sE5iT9jA+1UIRcN1WfQ2vOnl/a4CknHwK+MkyfUD1AKc63
0ZcGW75uVByPC+KWyxirYu5Czh1ptHS/o6wOiUAJCzhbNEWo4Q67VTz+e5IjtB0PZpkohKnpjdag
y0ejkjLVnwNAr1kgkOqGOjDTBB2iQQNw9XdXV5t8sqxZQRYNAuBWcEMvuMU/pkYHaw15BaXaJ7io
LhlYD2g8r3HV1SIpy/Klpmbu4COff+Br/jPR1QNVDh27NTgiBI805b01x8utBzIUHUSQsCRfdLes
yb1q09JJllJCJkRZteyEWhD2NyMO7OtbiF0SNCzs3M8PehJs3R549uItdNHunKj9GOZKELRVT9qk
iTfXpbrp16h2tnM2AK0V2CwZtsKf6UVHNya0Is+uOn/tLxscrbzHO9ir/buwWJyIr0ejfFk8YAEq
taFBeC7Gdy1U4j2kjgkvz9tQsCODArD/0wJo3VHpzoG9SSDLBcvEhI3XEto1s7EC4EhYFXHVPb+A
hfCJ0oXma3aoZl6oRo216KKiOHPTd1uOUlUL7VZFCrnBfdfQvBcL/UufWslUkGfGtEYa0OGcAqJX
wY+JE0xs37n4qfJt2sH4uCbiCiFathgyBGmpIeZUmNQaJtht8dVyH6sIHlecl1K8wIu3Wj29CEHX
OhrYo/EkdtYFDHrEGbli7SgYa+/ALnq765GSdvpgcGxxHMhFJ+KFVBU8JOCppcIxrPQjNXo2bQkJ
kUy3lQvHYsDPPOiW/RIq2ujaUWluGxoT+QFcU94YOWM9tRmii7opwerWrLa6bFpUp8zmtxhKSEpM
FGB+AQlDOXNA8youlPmyZrmTWLo1fqkTC9EPJGvGTnvew3mcJ0jeTRdfJbsMaq3vVboLIBL96xVE
i61QEMuqwNcDjqtkSZhCDGG7becNIL5bCwZlvUK7idBLFAEIukP+ckQuEyuQWc3S3ufINrXZPFhp
idin9LLOTS145YTiD7KztwjCbWo+xEDmaNQosHf4w8UxxdH7pQOeghTp3FiImM9FLWMo29WRk7tE
j+m1Ezj6R1mKSWjhwkrXoX9h4zuqY98Kw883bdS2ElMm8RUe3DoQeBj5ttIkTqa1tPG4IltDoU3a
cWwFKQNu6n1jCUWPCKumKUJBcbkkkLcVM8K1x2OTNt4F8Vpavk96b/lLXogNaG/hEMseuMaCYoen
vXshrlIEi6REJOKgJ9d3iO20OILhIC+k1TZnsB1SWDgsjqzM53FpFCIYB6LuWnUseGkjUGHH62Yv
TPPnQfw3u2cX89R5pF1cMcz3+Lj+2CrjwK0DDE7p+6TCg65IH1V9yigFvaMhUDfxjf6CBrHgKZHt
vqGm39N/42m99YxU6OVusSP4py1sNsBtXXlCrbCA18vX5rjonzFzxr1jwpBg28W9IKbkQn9Crs+g
XRZbvTiKC0Nt6X0t3X+BKRpq0B6CQzVXxWe1c87dbAzs3aBWROwkEl+Xv/ceIbTlJcZpPSOC7onq
K+lZLXbax9UfwehyNJjZGd7GPjUJteeK0gxZWS1H6qBBogyG1SZkf4n0on/fuqsqyOIT0N5bI6fk
qtg6yorLSb3MzH3WgRACXwx35ZJvyrygH5gGZ6ZMgqpUqJuSyrdTw2uqg4L8KFwasDE06dXDyQMO
jzJKymJAo+2YqhG1xl9R3NHH/sdwz8x5dRTPFV+1fmeCaNHyw2UccrCdR9WsNCcnfIhI7NMgLLP9
EwnTq3qNL7qT64QLYo7ukFYzp/Qf5DXuALecStsZOkmEDo2kU1yyUe2eXmOuh7IPRZeE0NCEKXot
jK9RGAJ59f0ubwaPHHD7kXjpIslBCk1mGrZSEZrvr+LxyN99ihS9Hk0HKHIB7Suyh89xp8IzuylA
I4qmghRrhtiKOXR243CNDTFSvmqQGBovw2FIPYPXer78E3n6vCb8g6VXMCmPWJrdMsDPf6eR5xQR
RNsmWOr1fceEzrzDNsHQ0kUxa0gV7Q0ohC5z0iotyKiU4f4TFoz1lvL1NC8dQtUHWL1UeuMFexeq
Dtz3ojYGMOJCzq1qyeyYpiDfuM5LS27BYsT3lnkQG6eaLGU7fmROklp9/Ir9pKYGK4KZHMzpXvdF
ND2wePwDGGH9W+vHhL9JFqL7xH3OXGgOPcVLT9YFU3THfajmv5QBnlgjDQugFX/Sj3Sz1frHMPvK
empqPfk3A+Ple2tTGXgO/iJu+2SzUauESNEXvWaSHBAVmTY93qxt2P9ztMjLQZmXtZBBMHQqyTkn
WCcy9hWJW117iZTfn8LwQXflL7k8sXFiia1d6TYUb0PCbVNjqFDRe1m+ikczD9d/nYDJd0IcKrBK
0pKTYSTCM3ctCbv3wUS0iK9xl0OQh9KNeoHf/bH+mYoWwcmwTuwQLsphwfB/ky09QICiI+sPomPR
PPyfaSbrP+CfOn1gPAPJfE1L41p65kV/ZvlDfancKoqwScsdRvuFKn8LzHU8o+77073Oq4joeJkH
qFM/G0J/wYQWgtdJNME6NnPRF3J+uIOW3iHqBQQEwMmUvjjvvPhqa2Bh0IdmXsT5yY0LZruRzxPr
gvxpdoRqTJn+jp8VJxufLIva+RcXZeCXI8SKAFydq4Y6sC2XQFHRm7mkJ5kXrL/7gmyDPaeIyWoH
ibmtz+LhRfppxYw5olSVN6SU55TQoOg9xbIWEeQJMJ7G+o8HtMxW1l4oQ/eYxEbQ9SNj9PcsCx5g
f+Qk7WY6LuGpcLmGVTu92jL3GuzJZfELnvzmdDTLKMflS5f68o7RwHG1bEEdWk3c2JMZZfKfQ9eh
xm2qLUXWm7SLNVvU+bxFzYQchKgQRTubTrv+YaQ/lyv4YyovXZSJ++lw2MI8qD5Y5D4BnyhlZUK9
RXb0NtRI3C9O6zRcL+pc2P2jPMYlS/oxPpF298nCaxR/Tj3/CP0Nn5oJtg9CuyiA9BRMID8ZX9Ah
TB2Qkl1sGlJZ00SzlCXqz+RaPCJCJtV47k/IG+ww/rizctY+mfoVoLqbUwYkFKgQgwUlOOv6mt1y
w+A/QlvnAz8HaSyayxqBfKzA9e601lrazLhEwIeNL1vBxGpLyUePMpvTlN/p4atU+xYeHC9UvFqp
//457iqLs0Qf8e4keKeLE9qQJpKyOiL+gPR6u5mNdTk7k1c6uSJk9n9otvfPj4XoxPBnddTmhTcN
F+Bks0lZXqz2mPRli0aYjfXHIg1fKg5zVd459YvJDBaPl7HLZnTOXSVHUaR0dqEEC8O1h/aOOThw
hrqIUrUJKWJsR9jNGrejWFKKBmxLkrClviBmWCLEODsz7k7whCKFkDXN3LAJZqTg/oDucJuS1YSk
Hp5D6WyYFgkQB2qTf+lnDHhfT0oB5D0oTOt62h3/DYtN2AqMUz/zWZ2IpAcceG18Vfp7fu0ScSC5
SEuAqT688KXNiRaoksljbGBAKdnTqWL4tEtrh5X5e9OCERFQK7wWekbv8BxTO8LVVflQshebYHy5
lw/VNjH0A4QMS71PDMIUGc80eHR4ud3d7WavvD422o9N4E1vcolkFVQJjN6q/UgsOEgkDVpIEakS
eI1VTGvyOz8pW3F3rShXoyOjvs++MV8fzsunX/eK3gkwPOXk8f3i+Q6WDGvyhbDk+BrOcB6ymRlJ
BR4sfh+bwJN+jqODJVbC2jYcpuSTeWEHDd4vqNnly0idF9Hb2uvd9wDoA3OuNMIR6g80WlVqiPeG
496ReG4pBSaSoAlupJzrBf44S7eQexVd3h6hcjsKEreT6LjDll8A/3iAusG1QR7S8gRccXy1v65n
jpuXyl/ok9pqw87Hj07Otp+yP/cUXCAPoB0C6fChHVVnEggcmExrWgiaHeuYwn5hCJN9fiNv+LAg
gNXEYSrYuX6fUtmD80wDFkZWxDGY6sXHqIaCdyuWnb0jP1zVQNM162obw1tYC4p786yoJQX/7SCs
Ao+uzRIof08xCU4NNiMZk7qVuyZJDGVIKOaM9T8+0z6qkDtRtqHFf7q1gxIkk7Cr4ARchHJWs4ok
RYGi6L/aRGPVIyWzSif5JOfcHfR+eJ2z5opTQ5B+0ZPVbvWS/nQ2CD/dm9b4DtcWS7yvoMXVMenR
wdtVDqwTegJ2wyBfi3iz1E/DAWzqsniFq1Rz1lmu+DlylKY9p9OVEwZ9/aXRrCmKSa8CHy5MUV7B
y+70666l/c9f4RQ9GYbEdltOc14UElWzUfRFqpI2M/Wgo2w0iQto82UKTsuvq5t72pqbt41CJOjS
6C6V8lv2vntQFStL0d+C+UJCBVJhj5QKvmiMhPzggxAHgCCyx1m/uog8eIJmFAVAFmJwnHzq9mB3
KPQlu8TsWPr3qsyNwMkq6DJN3zgXokVVmkdk+tovnCqTwDORGKCZlJfO0mihSoRpzsRyAskwHucZ
vVc6BrPtja/GbW8YHBBXlk2KeSHJPK6+nO0k2QUQeUkQ2vZbqWZL4Kb7vcCsCU5XF4u3QdymrxH/
j/IHjRGYYeYrhwAPDOCAq1iMf6KDcNpcBBHjkp6tbczvpOsDkAB+toxXfwdJCV3Tq9FTUSjYSATL
cghi5UBejzpH4OLQAuoL85x5OluFeU1qMB9Ghcx53UjezSe2Vj+5V58Mg3N3qu9HCTLw61Sio8Qi
90ycIeKO4T7HOOyWDp3pvL/qLOPSxaoVyn5AqP00w8o1nYh0RJvdcRrhykqpvB8Oxm24EslGPGpl
dkhkWdMJhXk+jc7hAsULaFMzojxE0bgHFOVITQYulFWRt4UC5jCSosnYFy00Z3G+ZTZZMYHppiBI
S2BxT5raX90teZqXbzGa/hvZV6vMkVgG69kkw3noyk1U73OYBj2Yg1oyJZTrap1q7/5QDmd1TPJc
zYdMHzAfjuM1wD00znYC25cqR8nrwFQ4v7FDSypSoAXvf+g2Sv5oafSjLc697Duw3CqlI7VNv6IM
SrWbfxLmo3yG3Vr8YjlfD5bwQMzTPcIojndaMO4QjvPL3yug7jkE71AA/CLGAnc15YeuUeaKtoQJ
p2fBka1cfrfU3zd6f2JIACu4QzZO+5jRISvl0oxAsmaHBSqVNBMaSZcncMfNn/K7b8Qn2nGIdYHW
UqjebRZmbIAZUfnh7sbTFCiEisevQEt4qC3AoS+X5j+dRc78SjP4h5qCIh6N1c6h67Um88+5Fdf0
TYJvM+3RcYJaQjiE5QmbTnuxt+A/AdxHUrvU9o/mhs4tPj9kK/GqS/5+UGaAUZHoVwlgl95KF8za
QRrkyrT+HHUAOEDbwCGX7++gCfAmmnzSEWIwkbxMiJA7bftlN46MTzUD1HaSPcMpuDaxHIGOi/DI
qdcK6CsORqcN02bWh/PuvFzcfP5f8fb7gZ4x7gmiyiak2FHI26ozOW84sXifuwse0rSEwPois15+
19pddZ4Y/62X3oQ7Q7qjCWrAweArmeG5JbuMBkHTVjV7v8jIlbiptEuLM2qhszloOK80fWsac9Th
hsJY6eHIHQ7sMJ+OydnbArEBCFtG9YaJe9Gw6GKFL/C+i8nbXiJ1yJpJQhYgzUnytb2vSP1EYUrB
jB+fc7wH1kZuyoAJxXbMEe6kXfy2cfMYkYrmvG1qLBQOE9p2BkvT8WSJxwetRh7lHYhlq+meHwPn
DxxRsiWctu5e7qHl862wTYOw/pV4sJHNDhxXoZLKkB5lh+7W071sRsRQ9dUAQ+AArQ5Ap7UTZYYr
TpbBuYLjhAt2EH1Y6yLwemyOlkswPPo6c3Jvpm3KuAKWnjG5BpImhe6NDDomLaVkO2O5gm9HJBiW
o+QCJt1vkglWaoop3GwPSk3DmMwQFiyJHUstCmMwrk4YwhDTatOb2o8+cMVaQIQjVhN6XGJDmHOZ
lKdxZa0YO6M1CPuH8m+yZXGgS5oJPvVdjFhYR7Jhhj8Uh1DMgS3kU+dHsaZ4Zc1c3vafNbon0wy9
l42gK7PMpRXbrw7tbuXF15qUD1UruCtZP3knye5dZ0khlveCmUCloA107ta9Sv3ktgIP725tncW5
sP8opMajsJJjAHkq9WEePtvR2L6GGeJSudSIK9LvAeBzj6pL231tbIW0fHOZrW8xmTKX+h5FZ6YF
Zyp7mr4KTDaXauGzTLJOHzBp949s2c5jTwwpz1reBnddA1UQaNbEO6i2e4JtIKuL7gWJRV7y1mzT
jIsP2D//JmR+uP4ROQSUhx/2Z5G7FGTI8ID3qbNAxdsq6VhHH9knIeruQannzrNuDyqge6mDjYRo
3WGbjijbT0MgIONJfnSKPe50Xj9/0/E11QvyCoXRvTMh1Q0rM/qbZLySCHkmwDbSoyIbPf0nW6ts
mrppcRYoy+LNy3WGPNIFNUk7v0S64jd7SAKYBXfPUGWY0bZwUUrznmhv+VyEn8Pj8zkPg2TLsfzR
FtxKsXMhaam6UyRrWZ7YdQWjVWbu3l+6WnS9XSfq8YijVYlrh3XRMCFjDEchN+7Epenkn9cRMhkz
g8Hi3doSVJWakyTmJuJXfFEP77wZZVAiJuPVDw92Pt+D98sA5KHXX/U7wjsILKWkxZ4AOnriYe/n
sQLB2nxm0ZbpWxLUZ+fXLiPyAk35LdIIvcIcDzEkCTfj1yjE+4SwXfPEIAZJ4nc5mBy75FjIRJXP
wFeugdPJWxfH7FTWoManWhQRUYwb8i2IO3AmgW5uLdBezUtGuLFxEwleFog4wVLSAyxuB/0kLJ0A
6cM6aR7RiGgg7z4g8Ene5W9yGlk9GyglFwEikuL+W+Sw05HhBVAP8jC+SYE9D5q7ehnVR9ivr3/3
NqFB6vuJ2eU7aRsmo41v61JibyQADTLVY/OfDsZ+KjZg0nCDW+STG9aqirM1YOs8ZHGUTtBaxTaD
NMgFAy66XVP4LzneoBp6YotA9B6jxIYX6PhwF+BaUXGTEfKgb/fO0oQE3XVDxSP7iv/I34uh/YWd
Sjp6AJfXaCjMS+a72+EFbUnBG/7FcZ/27nIgXQDSwa4JO9ilB//x6PQlnwmCwne909c0ZVRCUlT9
TeK9sUq4zZiwxOe2de0RmGlzoPVA73fXHepjY9qIyCQto9STIJ5j+eOjE+lX9mZ4Oe0Jo9WRihEx
AZeHkgmTiI3cOloLOBOXDeAfHDTcxzmlBhRvpyq/hXcMKdhM7IThoSm7dKltXvizmX2m2mwl18qF
Xkg6M2G+2ZhxyP8a/Kjq/BcjrPFaqaWFoPrWCJo4suWOCi6LmZO2uwbZntIa4imiuaq8HlgVFEDC
gcTQ28A49EX442fKavtbZX4xtF+fS2z6lrKYVVdHxmxyU8OBmNE9wlUPiew3Tfvize08l1ssC66r
g8RQJbX6H+1tb2KhyvE2nLTQD+S9GIe3a623VgwPrEhZJheNHAB6rspKBLvaK/Hhg7NWecwvZR1F
ihlTsYsgcfKK53r5XBbf66hsMt1CpLlNqZVSwneYd2LFsApD42IIXqjcgjc2dCFVncDAnDMXR/W3
0E6FvGVo6o+CzZQ/ZYRNERYqrmi+WBszdDI6bi4fjMaCfgkloJNcuJ6CpOVNmqhWQ4baV6ERVYOd
VlTsqwVpGlfdyzE+0N9QkgBdNLnV21E192KoTsvLBIheIjX56mhfKP1L6dLewQ+nxNoOQVbaw2II
wvvXpie0S53itn79XC0EmpWlooR+dQEipsRRSTZ8rw5VFhni2/rAQh+8MGIJqD4J6ayAoQ3G8fJH
xwwqgrYl81lVuaQGiNasfCGxeIyE5qnzKztvPgi/6BOiOq/NCMvokY6dE63ZxfKkCZC0nN9CUA+8
aeb0+t+O7mtXToZVbgtSlKQJp3hcVSl4nm4dC7uEbFK/qBGO4QRjT/tlIIYg7xRcPEJZc7cz94iM
h8/gYluoSCJS9cZ9imdduByVj/ETgQmmggWK0tyNXk5JEntaCRmsYujv/9UbjVTeBs1KVprUEPw3
mj/ACDal5n5j4n2Q9rsTJY7txDqzmY3YCPNFCuLOZwXVLqkz3Jm5HpmDYNfojnkjrrrVynsFmXlT
Exe7EOEXA+WCWAZ36VkbaSVw6WPNgnerrDn0vkLaGViR8Wo3vuMq9SJSmbpjVT5vyPzRXSxbVk7/
Vvu1oFcv5FmcPnF1N+PJeUpF3/865FJ0eW2qyGKduRKHWuBUmE1qvJU2u+fI8SHLn1PMVzmdSPBv
NI8M8l/ICDJ4A9uecAohH/NZ5raLbuiRJnxXHBovo7MeJSxOGWm2GidhbCtoCkuKCKoT0mao2Fwz
CgocPtk+ijfTnh0knJYtN2ssnkA9u36v/0ESciD39Q1ooiPLNNvJYh5G1ipqR27m4G5BH5SHAMbx
pXQk30g0mlCisQG6XeMKQ6n9GshNz9y4Q4YO35s1AdfRul/opi2r9e+rM7xPjW7IXtAPC2q4ltvm
vSbYkoXIq8XvuRbvJ39srP3zCSZUyTSY1MrpGHWsjecA6ZQQL1UQoAbq88JyszUKz0SIjySY7Nrh
tZGR21pFOz5SbCwWZbvM3n+LV5AOcSagZ3RSIHVPpqltSI6gKluN0xH7rj5Q8K/Sujp5vJtLVoMN
R+FI3T2cGyiGHAF7skeGAABlzJg636YtFB6HJ1I81kmndsZEmWn61bGCXpHIYBnoF5meapcpTc9Y
NKfngg0fwDX2cus/t7yUDGamhyEsU9U1oyJmKE2/ReGM9mpPGSKAE+bi5xqGtAa3vWftzl6GGdo3
fP+WWPpzT4hTFspnffKDa1q9e/742BtuyOlTMDjFw9DAVzzEVS4apAfSs/Dzecx2nU8Hh+raRPfM
JYNMim8RUDVVC440UBQKGvHkgF1l2y/C65cAQwujJvhDgDwCAs+FMKMsnxSDe5c1jN0JEy8z5BeJ
yiv9EU0rJvTDX5CjxM1gGnfLvUVhEYvB9XqL/80TMq9IKJ9czb4x8Mx0E42hr+eGRtEQUrtIVeRY
vh6hAuw5aPSpm04msCUPb8XVIKLYHsht1Xs/XSz8OVM6NIbc34fZsWKQv5oZS98Eg7/1emHofwL3
4SXh+7fMBJg10ewLMcTTWGatMvri4S2V6Cju0QT+1AyR1R/mcVQJr4FvDS/TXRpIqRC+/tm19oZv
kBRf+x/0LJGWlPCkKt9n3pVoelO0yFMg+k8O87N6H5wHt/GZlqAgwOY3g0a6PeoE+ZzOVoJB22Cm
/ozV/afLE9yFLwCgmwXbW3G9yg46wWODCzB0ahiWO65Y8ITwBEHIfQjHPFJid704b0qnrd1Mb4hW
gNgOf34xebWRnHNb/EqErjKAH3hyfpbpAL1oZx2a2Ch0nzIuNnPG14UFx46YA+0Anwlvwj10YL6T
UA+FJECVlBE7XGoVSIwAIGm+fv9HZe2K7SUzunRnGJ8Jtl6q+7Ti1B0Eo04AIWe5c6W7ckp7dqFd
3wllsbzaJVcJcPiwP51dz1BzwdqK18RMkQWDaVgwto6661atfsEuY+tvnbkBqQ7NiFaMxHdlEVK0
C2eZgBxd6NHAEKESxnYuJvrpHumCsNrV1Tbh+AJ3Yd7/1gI6ffKXA8ic1krZtJlFT7asqYUxNVeX
EbNCX8i8rCP3MJYd8S0dZ87pYJsJMgG/Fz50YGjFfOPiqLJ8j1vEto0jHkCZ+VHzqbVark4hTes1
uUKgQC7rBBF2vrHfnkIzPLJmYQnU+nMpO8XC+zReE267nBaxu7PGhmWH08yI2KmHB5Yz6SbCDLUv
RuzBcT489iAKbETerpqTj3l3tCsvYmm/EicpIkdoPiyoNnK2hBBpJvpGfZEROYxg5zHFjmcYGp/k
7YTKDXWjPc2xVYGQAefiXBlU9vNBGmaqHZ/oblhJeaHEN1EiOXp6F2aDIUkAuh3s0T9SIvUdl+8G
cwes4rkbh7BN9iaLT/hJ1ZjhwCDmsPmk7P75C1/wY2ZKKnOVAekPsfafFtiUM0F+CvlsidkYom/f
WbQjf08LOU12BYWfvqOkDFvM3Go5k7vrthQddkjUBLcTPXUVwL2jztqqYsQ5UPGAx1V/6gajkEp+
RqRA/BeAIaisBPIhIRHFAGQLqnmkf/r8DPFdxWpigpe4XmMMHd2lPPUsDzNwatpEG7ldR1UOgsQ3
S5uJdo3oFb2M+g5G/RHWoVX5hMwSgoacE5oScRhfAFS35sw6/M0LtMOlOjm6BBp/Er9Ev+U2gjCe
yeSRTiUaujsNlgD4A6I9XZWbFZYjUHnSGrYKd41Tml8dsjcBUBo195yNt+1HTmLCcfmHN2qFxm/a
TjZkuXLpTP/9K6lE+xQu0/ycnidkCaNnNLb/fCDzEmTAtbw7Qx+4M8DIJLE2phwyy8ngfO+hHEzs
9Gzm0w/0BwS1jOdWH2yZOYLqHKqz2lfg7/icZVX3woCtMd/7AiS4GHLewuKPRcwuIkDOmwqHQkoo
i9emT9hCj0WYXSlHk/A8VD25QqBcjgZIttHxHnJBT3kpxi6W44s3XO+dsAzUvdrYtp0tZUEuDX4d
EaN2aaVqozhQy10VLdZa7pH2eCZ99UZw6+bBTjVFrkCACwhXCx10tPnHTSs+cADtKTm2ypn8bgZ+
pIpUI4y+yapPekdhr38+SJxap1ukP66/WDZvn2SLyEFZhY+RRtmXbzh8Z5cQcnqP9szSdKlHteDN
5Mqh9UwzCSnIi0MAwJszGazCNEhvRSpHurb0MocfGGxumtjGBrXeMknURFR10eKlb0c5cA3ArgP6
Yqdxkh0WIhBnJFzvaxWG5T2ds0reSYptaPLr7zA35gQ5jtKXjDlKmBcLRihtFyHrV3JN0CM+CyM8
BdrxgYAotP/o3VKHwNdYjIYAMECcFi3SV+iZl/Gr3M+E6VW9Wf2dHULnP0jnT6CpSMnaHtrboVBH
/7473MIZuju9wixWQfMa73fux7mIYd5VXYnLcs2q18uFrAgobzTv8TjX+dcH5ke3jd8au0rfttPv
1pswEfML87X8Ga08XohvYpJEMzS2l7XdX5sxZD/1HzLZApj+FYjY3NVEgn6E5d5Gt9alhdWeNoOQ
ULGRKMbWq1sHb6Xb6/0JVdahWkcTtBqqeum20jkos4J6RIV/1xqkecLciQcxFmEuImeDr/+RAZAa
OGhlOmfGAqNkvHzIM+uCfR3Zv/4eeUGBhAUBp5qW2lmFm30x7NbIZOrW6CHLkiTh6XLkp9puJNtx
ki02siDXFSPu/v1EvEAw8Yh54Ze5htZWrPI0SZsBf4WeWm5sLKO+zmPLvwP9B/h4YEz/0L2HycIJ
snszqHVUlAVNUBQFJF3YoMOVu2Nkb/GpvdLIOFkuYKRqrpeM4sEn3T+mjTYdUrGqRu8Sh+3y6h6P
q4Y+xlCRNQP0lgdMH/UTsS1F1NixPsPzk9tPl/3oCZj8kxq/+DxstRRQ/xEkukTRUVrF7f2hPHgU
HJ2rNdvePFVJjCSfecWDOPiF/SANu8qUUuandqsdz73GyBttCXHQucGlYBFtK/4caUk64nwxmquX
4yLAMYV33XmRrf7F/O4XztM1tyjwrSY7XEl2ORVDDI9BnLGI1reOpWnbEXIAUfeeEUDO342gnKIr
AJwxF2vy6i3d6WydUmHbDHX1S6sgu3nGVjHgzsbYDQIauchw41BMH3seZCrWRIeKgzztSixji1Tt
mCcHh5lZFvKLGBjMNuA75tWgMhiCscIgCbtz699NKdXn/nTqse9UKc6niur27X3XAs/wWnEq+niJ
iePKT4QztcR5XJlBNcG3zd3iCPx9ekhcGiyt531n/XajSI6vKDEmH4LrRYtv+NgPN9ixOhxRcFCK
23NJN+Tz6mOHU3ilD2wAA+W1H4SPSSd6AdcUy99qPBWH9/7r9/ijc4+rd4ab69vbP7bzYum6POGj
RuThm1g40sRxEfn8g5xscmC+TBH97naGC4+l32AUrbHLnMoooPp3FgFkDBCfwQMojDk17o+AvJZl
2fpbqqeUDQg03pEQgxynofrv//qdCxfaAc1lgbqJIJVipJu6+avkL/+LSFKlGCpRVYbGSX3o59DB
KxFJCHdUGDLj2+zSIwaTDrSoJVpiKssU5Po27WYw8nXdZCMboxADytS96QtMm1wCYyaWOIs8peu7
pkLcOWGBTVy8DqVqx1Egpq7GWBQ1atUH9Vr4M1AI6TXJBift2cPjAnBrNEztYkuBo84PoFrMSCXE
Q9M2NGLMDb3ohVZ3A22+IN+jK6pz2S+UzrVf0+BWWDzEjW8KEYXnQy6nOjhLReivsNlrRkxSSV8o
hZF22ASbJD5d1pBHLFQp++chXCAYVBelgJqXvQ5YE0lzXDQNO+aT6SkzdXqVGfugZZz9O6G1qlqa
DnYVqqLxS5vJV5yhdWYrr4pFaWte7yfd7RBXKBGD+189IAdfXO3iAJ/MMWfkTQkZDen2WIe58qf9
mGUfL34r43/cXvIElMPxZ/koIaNXVa1XRXy/pt5z9iuLJcPSieEdq4wUVosLrXXyUV9HNNQch0/n
GUXD/hMsRPodRSo2fEMYoqhnljZZoDQcID4PZ8qERI/mQXrV4gIbvB2WYDus6HpQ8JZzKs0sdz/a
YjIvAZWeAM2Z3K3nuk665XM4sJA3y+L5LU/BH+ytHtuEEAgmWavd+1LIigzTI8U3aBrveJ5Ej2Vm
OS9pW8m3D5jKPi+xRntfIrnJdfUJwHVXtU+K9jrXcLJXT+IwqVu51QbuFwKn5prcrhsBaC6oPR82
SeNJJhYFnpgE7p78uHhCMM2AyYADPPuIelwDP3TmdwpBkT3uTjgKJejYd2AB1Kcv/A5aKosVdbUd
UIpQmjjDtK1IzqsQlYXF5ifhqexSsR++A2DZDX34uC6MVl2MSolTvOfHQxBv+ao0VisLzZdkukZm
8hp6616ZZIc4FmHeEtpYXTw8/HsOXpNfC+qeLXBuzQoZ901L9UtouVfYtaxzVGNogCMS2g/1It2T
rBloiXhVRuUPnc5Fe7fCs4UsqRyEnO09Nwxkcj7R6lV88VrJBEKLLxUaBSfJtImRbNXMjbAVMN+C
HU7FORvU12ZoJdydnKBjEgg1A2q2iwtpi+eITBQ7SyDG++UTugnHhe2FTj/ytYNxOmbBg5e9fmrP
vFP7Ria+gCnKowyAGeYD0RIG3I+vqbWKAwojc0YwMPfn/xroa5ZDMU5+RCE53a9NcBmr/ivWzqWv
cv25SJ+W65ip53fix693Ie3HAQO90hOIW69c7gN+sOhOGqibHUmoFOj6E0ykdkPmMyiVr/yh4VbJ
PeX06TQonDV8gPWZWjUnWeYFbsr7/bKhH2wSMsyXFr2XbjQiX1EdGaJdVyfwrW8A836md6DS9SJf
NACuoMaj8PK3ITpwt5FfIOH7yULMpxSJhHRvpeEWgoEbOr5ioPEGjPkkMySc8yqGxfxsA/i7kxgU
6AkvA1AHoJOCFy6ShTqO7UFOcSWBZMNPH6hUuKQ2BWbIt3bhWSDU7s957AItfkVHIa5bmRaFUQbw
7P5GuBeiwwzwHXwbbJYba11kja+5BpzIXe48FuSMxZ46cSf77g11mEFxorWcYtYHxNXy1GKK7JES
roeExNqtQ2V+zg1jTtP0yDFkfeqTXHjzIccRxTReCi6NPPZXpL2QeJvnboYsLqFYAVNV+pgxDew0
n+u8I5pJedlOgELFhiYmJTKlX8TRhVm31IK533QmdYnuvk5lBdBe+hjDKYowwoMdPTh4rc7C1DR1
4OsenMJk8Thg7ifmDO60Tu0uCYhCkmzYpI7rkanSvOCRmkGccY9Q1WRgLwMg7JNOJAPVZLy9zcx/
FyyBWAuP2uufibgM5U4jPl33wZOx/ieTEgbMIyQst0mKb08e48QDdVTxGxLXDOLrv6vubxj17qMF
DBKYU64qvvEKb/4/zzgJTjh5fQQ2JcBOJmborP/+Q20JXpx2XBimr7r6lZk57TwyJzZoxwkgrmra
UgJVREgr5krR7sxE2sTWJ/0coPYHrV9kDbeCXyrq2BPEmiNdHWePqrxZY5CgZ/66O9r2cZWH/0PJ
WrTtKJWbbSPbifrDsmUVh2qWx16K+4gZeXFWI5jIFfKUex4jCQ6GbcNAqGaxRzvs/6etjhig5/aR
zt9bBiG2Kcm9QAKr2Ogn2IM+aGlMCWoSr1IB4CutgtA8yb48EVWoOWLz3RGFtl/Tgx9Q1iMI2fJn
YqcrtvLUg+97ifW72pHzZn13In8234ZRskTIZmCp5R+B4VT0gvvhiooMW6ceYn4jkPOak75gY6pZ
038xD3nRhkTv1YfTDTw6FHPlCcZAkyDF/H8yf53RTNg+wn/megEI+nzxHyGPSY0giKE8nrtcfmqc
yo7oBDCd0jfzmysTdESmusrno76kicLRpS6yaweoNMWuTEerUpo7tDikxOcNFqdIrvuMha0ckFr2
O6o2lHsdO9d/3ls39e7hZtDJJRTYaZTsQlPmsXQJShZlSyvuNlT08cWLeFBcYU04l68wJbpnaJPc
nOv9MYDNqxeF/k91AJrl2HiCxh5ntTipMjKfnhJRTRnNrAO0aKU8bQRw2zzy1dx0rWkKBZoxAuD3
oOdOp0BNxEIR/3ObyLVAkiZC4EUJArs63X1jviUkgmwVJFJgYRXlyLn9mZCarGoYwIkVI29JJvuE
VP/OBF/1AvgeZaW+3OBhT7zROUBGGDf3Hu83P+5MJaB2ipmcS9f72FWxAljkPrLL7wyk+cwK3gQP
ZOTtZQqJE95pfJRb1RInCX88R5P4OIaTyn1ZctcPoknj0pNdQVJIEAVT/2el6I8MJUyKyjBfhz/3
xiBjgQ8s9YnDommlYuhY4gnUXibMO2z9GfEAUvnzi0dwGC0wYJ8aaLxiwEplpXGzORa4CQGAb0Vs
hq49uYiMACyv1P49DcBNwX7HCkKe7utXWhifh809W2et4nsGpZiKvFVgb0+WaxMAL2E+QRh+TEXD
aMReLr6SW7O8MInEufEuugMZ+s4ZB9dafdIvbf/CP1IKSOgolby4Qyj7oFZGKA4KaRngh5i+3Tm1
/i/DAIR0u4+bYWbc5lETHL4fxjBG/KJMlaTx/a7g16rmzQ4of8IfPwGipVQ7fuU5N34l+IMZSSPN
HhXSRykHKMWui6IUBHJbT8rpvtVjG4PM+H7RaYUm26LSSiMVDqF57qnfooQalPVGIUzaKTi/qvhN
1qLar9ZhEk8WbAofYkEPoaeiY+nWOy7VP/N1AAzoadfT3GVhgB5pLF54s6s+SpaRfyCK/+8HSzx6
UUGQvrFgyzNVQF8Qxh0NB6kKGUuCOI7ChzW8mu4Sdgjr5GUqwDIkRNjKe+9zvNmfH2akByDeqxrJ
ZC3W0dLPBvchNHkUcFzj+s3v+IQ3OuBYwkoGARBQUc92DG7jFVPpZrxdcRnb3UsZSKTOvWmnLAKn
KJlBDEK9dvxJ8jbxwMFv9vi6YdlGXCAg+J98bokiuLrh1yhB2NL9eAbT09ajS3t09swhN48rGSC0
r143/Wtbiz3EdRtT+Trgyj/qg5lq/wXeyKE/uqaijEg7kBURty95RLhvB3gTRoh1TeiVvVZYxITm
jP8cS6q9OsTQtyFd/gOggj7tDKbLi8BB0BwxhZX/gWEfC6h8irBOR8k94LvafIpwFrAYNCUkEerp
lSVnVuQC9b7EJ8TFIUMs5MLSdq2xMKZV1TW6A/s3l6RNJfRhmlCKUjHcixcy+WDYrxChuRyrDc9K
uCNsXmntiIP0QtpqsKhDe+bUmk+xXOzrXMfcaMSj8YSTlRPGkKvQe+zR5qITIbTmoyxsgmGEixiY
kM+smYFDlO+Mvu3qkut+O1oGveWV1WZO6JcVHo/JrYufWon7XxEuSXqymSKkRDPlcJ8Vqfux/XMb
4bEUGGIFlLt/f9wVkLnvDyMcrbfxDXV/5kq6Wl4yU0B9rznQWgzP6tEldS9K6I/p3zw0BIPW1juJ
ikBvCfFcYq/3hr2yMUq3MjiEi0u8tpfMgatIoc9kd6PR51HqXITM5rfqFG/amJZg2oRzeTRVp2Js
0vp9PH9sDmsbfRcQ5jR7v8CVqsRmmy5iA/j2YyTN/15W7wxt9DQQPel0RUZy0Sw6MXJQrkK6fJRU
WCm3Yu/c8nxZ4gtTyxSD3FW7nVoOdVsJHc2jQSOuPWpJXxWRBSndquaTjaNH6TPDRFKGTydm5DIi
aSRfkFJRFlz+yzXRoDpEqOZPnLzP5CdHuFTgJT0RIPvIT2SrPoNf5gxOEo/4ZR+uKCHA2F/y9OgF
sCKliuLYiid7G3gldlxF5aCh4EP2C1LnYfzmqdj9KEI6sqq9m7JLXILtFPtEjybmgCibibUvJ+IH
yXY9KBHJxjVkGSidnPX4WXd7UaKddCaU09hCGIn1og8J2waPCK3ncaPNeOlEHbXlvKxSRxrFM04r
RsNStLlFKXobJqhZd4oJj21T8YFXj/gFvKP+kiODFQnZM89tZWHh9vhOSgLt2J3lWAEzuimzqFnQ
Oq6r6d13ANSeEooY3nzeFsW9JvAgElY7mBD3+ZnaoARuOibE/T6HHbs3cIHcXjiS17sn85s11rve
NmXdK30oCOt/sit8BO8J4iU0DVlPhp6hA5ybrO4jgxDAsmpXcyxm6Y4Lva5wE90n6dfF03AbfzhW
nddaOQGEyirif5ua71Ktz/Bo8IDTFJ8Oy5c+00F/I4Ykk/O8S6whJ/mmvcGqNNu9RjDyDb2LY5Xr
0kNyz1eACBdTybJqYEdjfQfB8EDfxodoPnlFe6RJhq1bEpH91gf3eACsTszBvpeF5TGmIGAZ1EC/
M7vxBlXi9GfH6jfZD7EbqLOriQWQzyyjpX7ISceNqts6MtwaQ2+pR4jq43dtDOZmAzmZeTdqEC3s
kdMLfisG7Ifw+x+8ciF1vn/c5e3xuV1hfypDvt+SVAgMdKf+ZqLnGij4s/eia99WdXjqVJ/jSgr3
iJTYbhl6NESll3TQ9DZLw0Ya8dZdmS5N33+Joey/oHaqHxI2IRvgSiwH4NLtMQunl9P5NHOc+7cE
JJkJgeaRvU22hSM3M1CReeABZIUH4I/8CJXIaMQ33B3qJJnDMw9KZTzSYp+71qsQdrJpO76ChQ2X
V+ZzseX+2Nk27qxbaag7P/O05r0rQooFZZVDB3t/jUeTu5SxKSQyTTPBXCa3iOOcU1JD44SZ1ELu
5lCEn5y9ignpLRPDq9xau7cPlglhmz+rkILa6cthjkYNr3trqhl7fllvjlSRxp0vMuqVL0wRiqXs
DlBILO3dibYHdLzyZTzrA2B3WXFQoGDU/Oh93ZmqluNcMFdAPFQPLJfnGB7232trxtcYPfseaxEk
J+a2wFKe0SUVsMCsf6CCcXrb6RzwfzemSQ3YwajCgOytckCY5m3FTopeKWlE1lmm3LEmc7T413ZN
oT2GnHSmFXl8LezLlBTuqYiJnIElw22taWAfVzizecVBiSuoApojBVblyabmYA+ww5TUJjZSm1RA
UJdTmpBdvHx1Mk/fEzYqTy1D+t6BWNObIDonFmCKp5e38f3Pnj9oQZpiE+cyWhmYWAuhT9kikSkb
GC2O+iEJ0QRfQ2Ad8po4f/pXQz56u9evj7jQk0qodivTEHGVWv6KpZX4NWGuaFKnyf6MnTRUYdu/
2oG5YsI94+yC6KDFe/A/hGmNel3ir6RU9+UgTM3dXaHOcC74XK2LSUFy1Az8MA5L7H972ewI+uzT
hzkM18kxzLW7EN3eR9VT9mf4xLqIQYg1rWsadUUhikmGbxRnI3IoZ3C+Xkvmh40NY9SvxV9Kvls+
oWxexJqrFsr7yZ8I6KQNSp0L8ecEojzUlLOSiXNpamYfo19aFhQqkrhfTSTkZASGv00fP7RMLWMG
Vmd0zoYVSwD3RVzWcvbU8vFG1gCvFq+jmq8w06ITYxa8aLooqgMBPxoEO68+7GgJKJ2Yyp2l8PD3
OJasSpyNScI7NH12HSs424ZNLgCJX6D32pCZ2T7NxDon2Vfd3E1REHFygXIlkuGNDXJwmVcxBW8K
KD2BvN9MT+Wz4HXrCaWV5lsPoydb9wXYw0/LJFRNx0YeCHq6RCOl07AAyVIgucV8F9H7UyzCKIDN
OYoo8yz58jL+bjxXs9o0uOhBiIHKzE7FPs0UGlTxrtQT3/IdlHpAu33680kyfnfk0FiranrgTETD
ZbeJoke0+/Kprhnby9NJ/UQ2lxw7pJf+zznujnBOX3dTGoPy1CqpVS4hu2bSW/yYtkk/cUSeHGzm
sy6jbTtLmIPuDdd5nm7Ltcr25lXNiTd/zVAhRdFMgKjxrjIgtN+oIrAIgIDHeGc49CxT66wBuOWl
6jH+lMcrafiMlQEXSLM7EsydoIjct16APpGBbRngY7fvPNBpMcKigf5/Oxo5LbQWeDtDNt6I0kG7
YrRZCjg+NRJRSIeL8fIn3M/bV5H2IN9Nbry9Ce9yhbSUkPuZvWuaLnVukbqMMKkjNQN/HJXKPkOV
MQMl4FuR2J3KjMAqZOxfptfsQloXAP268124vWxCMcM5gL7DyQfyqtbS4/uBanB9FiTRo7ZdD3bT
X6EKspD6Fi1COU+yv1sXkh23rV06eJd65oaCNNE6tYafsbK8yFW1EJgg624kSkNpwHd86OkpigoX
MJ81lLSpjncjf2zT9BmGYz8QVeAC8dVVTdSFAAAPK2lq0H4ToUmKrSp6UR8PhmRI9decs5KsIy7b
83q/HysG7CpnHrbviD6vHaTNugO5Gc1aoNzq0RI9XHfQNzML2QfRhVK196Hua3x3oJMfClEr0HMa
F43DDXiyaMiVgQz3Ksnm+3X71qo7koTSd9Xo1L1honEv7GRHXMCGtmEJ6LBIQE1itWwE86gRYYf9
5MeJvxSXXZRqd6XYcRgb2dAsAGynyV3yhNc9o2g+V3K1JegV+ZnBs0TNcJ3bLjlag1vfJgw6vOFW
ehfoK1HLAliPTQEXbWd+P0XIZGYeG3AtsBHgHwUx7j4rWO9rLqbRSHsUNnJSwiZZqGqPNcXTO/vx
iuD/yXO9OPM6TPo5zYlLppgLD+vYI8URFvagqA081h44hnEUayMmDnfsomt8/0sPD4yoPfkWaSz5
FvGzkvzUXw55AWY6/RHR1SKaSBIZWMzIXIxQVQfE43tecvczYWwR8JJLElGd7pGCMVhsNgwbfHGZ
4lKs/qH/PvPtFGy9em2PYS5Ir0YOOshRKAEPf0cgDuTCtpmBopDFxMNyHBzM2t0zKeZdj/anlZLQ
N3MCzkO8182qIL09ue1FVTfasnnwp0uEFooD0sHSzeLa3iixILRUobAseYzUYNzk2CU95fMZ5QTA
Zcp+7Mbiy/en3qrfUyaIAihCFSd7b8rF9GMwlnFjO3vnLBcv4zvlt3nuei66HWb01yWbZZFZUKhI
FRnj3URd8Ary3czd8DrFWTKLOBGNMQR1frT4sgBlC1ZPiRYVSV0AoaZNFgG8K1iDE78GwV8jYJ8M
fUpz9q0FzQTjTdoXt94Ppg2qO5dE/hBAzIFYc3xFlOXvTjYxLZhxC9IBtYXPCob/UmP62Uff5SEY
DIpppyDxpUfY+drdU6lyQWcjBprQ4MEfizn3tUDJt9rCn/Lkf+AOHlHFq4bqHt/KjaLUYsFbUbJ4
vV83VYjErzVAMq8DwzACZVdGn62e2tdQrdMpTX6uFCdIezTAmrsak7DfozQBBAZAyXnreMhyaUmX
AcxJ9lACDAhjc4ZjSIa1CIqdpFcIW7io/8SCw+GobdwHvBNPNSmm7JtRvnfilncwq4rEhJJQrFZH
oxnnrkw+0gWlpC6d95k/6nVPZcLIMTAZ8be7TTAvGURipB5dkGivXXDKkPuBcApdx12hbdF02vwN
n334pgjI0DRsBJz4cQK8SFPC671bE7f8lgIUxGmj76gXFgcbMrP6sFHbdNYRedOMuTTYw+NCYHrg
0EtLRD3/fm4YSkjWKjGpvsGHEZLxpo4lO5Uvriwlia6zWg0qd1mbLchCgzh0c8R58X03wB1hnZ/p
3FtjGzH6qa66Z/HwQUSHQJkt/oc5vpd7Ld/W7srSmsQGqjhoy2kxafIwsuGVKuyCceC3k6nYb+GP
+RH8wVJr6WXi9+Y/LaSEyw/NFh+SHMr7ic2ibTx4QOBLbhZ4Y1PO1qXiWuJDkCN2TA1dYS7FNp6A
o2ZCfcD0gD3+zTMfCMoZpqmFKFPwTE2Fzz6N5kFbohxCVVS5YFN+91juynkD0i1cbhw5ViGZU7e4
z4FOdJOvmHVDRmq9KzjDx8kKsve+ub75JopThFUxYZx0VYxZKVp1Z8adi2MggP/texc/uLP35DqQ
6W637XPRkaEfSm4j67X5fAy9s3hFsmeWJj8oGujSHtryUDNsh+wdvPHNJP7ahExTZeuy/XYas3Kb
2zZ+MJMiB435cFa74PHYpuj6+pxXPssJFf+q5lUX1m6PWawb0ewwG6roYjwg/FqYDm26o74Yw0bi
9H2R0wn/FbGphLuldOem0I84hjlin988ifBcJvyyw30I1H5Ru0boVXxQU1FqQc4JN23urSMYTxjj
N+5rZkiK2p6L8njMToldfvzekV0X1Q48k9xYxNdhpCZ6nh+yEF2phOIoz94PYDG8Ljk/cRhHTAW8
i7acYaMq2lNOeYjGGUdz2adwAAeARiaea3EGJjlnlDLPscNH3rxiDK1yCVz0jBkiK9o5vDsafzXQ
SZW2P9W3SbImB73vHB5ZugECcI83CiGOmKXeJZLdrH0OHScyMBmQ1JsJ9KCUAtK/5gOEUxqDElkY
ph839rz3RSKNf81f6n+OFHCUPNuqv99jd1tkmZm8RoUZzhnsyFP65K0bgqlBHeO7zDcQ/j8ziIK9
y+qUk8M8XbfiwIvBNdGG0IA9K6dMz/gLrSJBfqskTKIkHHxqtG/S6vNwWKLxtSBLV6CJeTyEbNHz
EbJXrq0ijL8DdUwuYe44BM3paOFT8SSTlkHLV0gAQNQng2aksnULTHfN6Yp2/dwyNzpRhqDXByQC
bU5+aZeJqSYF8bGfBbUj3Cm6kCSxsmm3Cu+yBdjrApS1baXNs1+o45KFi1ivm66jwBYYgumoiX67
ATEjCim8P7SZ7PjHgImHkQhDvMGrSdYEjZNm/VL7DIa1CJ0Wqp7F2mHHVtcwbJBRlVhGpds0wmDS
Rar8lbfGyznGQNPOtEznkugG/D5A5r/U+HO5pXoGPljJYx1NqljOVrfKjPzUfyVoYm86+XFXr/rU
QgkCFGA2TxghOPtPyi/ZzLCbkFf/IEapEsivoWhgUzjJr8iUi6NZQZqXyT6UG5rXHtR5cv1wdLJO
wZM5wOA15cKervnJo90b4eFUj/e6FMLGSAN7WWKmP1kMQpOuVPOyWASb7EAj1dSpDxXxrm9G7gVp
dSjUA5gzc6cIfA5VDO0rJl1p/Nan0LMrAcEVoUN+daewwAW3iZj7DolYYIi73RIqIpWUgjjRFZPo
SGMh5woPf6Che5ar2IS390Mz6ZukXGvFVieIdqqf7jvEyYs2haXEogSgJD1X6D08vUND3Jl4wafu
PkQ6iA5FFXHUz1QEHLC5kC04cVwSAsXAy/ENh1LBq2i2R9XH2VNs9Xx59Bd05P7S5zb1gYyOtK+e
utxpMFLx+Iqvnu4hNKtHyR4mlvBrWuCaA0tRgT290KeniWNRMZXzVuVs/JvIy+mmFc93PNbnepdY
Hxbq3BNfO50Zz+JMd2CI5tRqeRI8+tvOhx+y8v2N+aqPokx3WWAgDfZFd4WUcN4v3y8aS1HRzMN0
NRdSp6LCHQ0y53rp6J4RtP+7gqZ8OPM3Eak6Xj9ssWKDVCMiE2HCkDoCIGd6sQPlF5ESAhqnhQzp
ZDMGi8EOjmGgmyWguqzEpFQZTARHbVmVUm4tJfq91h3ZEg0+S9IEDgna7SaKIVrikXmgCJ/mbH7l
7H5Xe+4sXYY4pynz5rVuhuvO54CWHv3vxVD9TUWKS6NNeTWtmQPOFjlkhDB+2aA0IbcJwDPvfIVj
B5OfAU0dwYwD1y/qPl2GFLk4LxgFU//21t/TNUAjCLprKVkEq7ioqdT03NYR2fL+LDZYHSC3a209
6FWE8NhsVKvW+D15tdq+AKqShj3L8NzblgLEWMPQZevS3/9gZBLZxJ+o965/vnEXIH7aVBnFLZF8
+Yd04oX1xXDuDuR1lPNNmJ66tm8irEfRqFX0/YmGx3jc2fOhK10BVdOSaGUc8sXA89wb02/mNz/L
Mw0CyOA8xuaeAZ9IJvT2E8gNb6ETZ6mlRzyMX4lsasUR9HdlryHN8HHfabTeXqNrtqd2lk0rq55O
glYyIkfQDSezsKa3KjVR9vqgi0IQhjhIOMHs111md9W7/BWt6cChOOV+D1XhAFcyPeeaSiNNANTV
vVo8v9pdEdxW90PtkBaGrAoVn01bxVDmCmC3qkutJ2D+QDCdmM39Ku2CTQicHv6lmGydoNVAXv4D
qEAJ3TyNfOrLrk+Ua95YrlLgaYYkuDwizsFloIYKOqAWzI2/RY7D61C8iiJn8gqCpK57Oub8eszv
AckaC0viExncmwe/CJyrUPV+sW1h1JcntYDejdVQA95tWZFwv/6iVlbec0mUhDqP5dVdicGsFHFc
PTKJ+5fsNe8iGnRh3pp0oSPEl6dTRAt8JvBnZtO0Bhk2HvepNWIv/9iE2vqeiVDxfcBq4ghqXYyV
JO17bEXNi+CqFNcyxKucSE8MSI0GTC1WGFITvZK8h/f6zUCoYfbrMdYFPTR+1XZkWsvUIV4nRBJ/
NsP2gUBv6o8RASYuzTcQCg7FR515y0OoQCZNv7hLETLoT7aT1k4dUco3gHAJn9SX78hfWXSG5luK
Ek8UuuoF/vVo0676dNPq1XUSmBP6bico6CsSsrvtVTjKFlbPItC4/+CR1BZJwc/PV7xUK9k5UIMQ
tF96ltJ874uvvNhItcZWJQFlLNRKWgQCq+VX4XVJtbQZfz6/J5pTTDI5W4nnA2NItdW1LNgdQJz+
v8TrU+r+GSHj96cSH4dMaT8WEP2JJWp06slI2hEkgvd3GYmJqQ8MHIxyIGKGN9eqqbiTyTPXiwsq
2PfNAwW+yrALOSStMVlqiUr5miuWZ7ZiivcpbwioQHNUHCSj/Oh47SL2zOJb/CA2l43SM+kkcHtd
+hWjTXEYQYlPWP7MVE5YuXO3mld9Zj717RgCK5+bqKHCuGWVACVnA3e/zCAayuxsLN8Sz1VrHbN3
T56I63FfHJcP5VHP5XOswBJe9ZbcekEF1o321bFZqVCVkhNQHD9654JFiMVvR9vFYuNUemHQT5hc
K7cFxS2gNxolvZiT4jHZBK9gs+9WeiMlVyuyyGswzcG0nNQFjN5glwdJOmPIGqGoZqBiaBJBvg8Q
Tk0QBj9Fq+Bg/WA0fXAqzLhWnXqvv9k8W3OGSZdZ0xiECdkl+MetxT2ZlLj2v0+TLFtOY3vwS+aA
CmmWFV5tKwylYoDWJLAriiGAGBnJ6wbYEfsholQNt6+bWILrPfOEzx4BJKN7H96xlvMh/MyStMiw
8fK/APuc8F01hKrGe4/0TsRFANLI8MyvhnWpVZyrZAyJWDvbkQZQjz5zb1Ul45i2AXIRtTKocBzR
+A9XO5J1FLYB9d2W44fBI1o2po9od0c86wMmkcJsldwIeoI75P3gAQeNLVCd3iiSXOAtu8VQsaO6
pBOzD2CJw2+BD73wTQmt5jJ/sUiBctmY07xcT5olpLHK6dsH0QmaSPW/9xeb/eEth/87xEP8gAKm
im0ByyEMAJbKzwcqRmiKM+JK/CTDr5wd9OTCSaf6W82H0W53/9JI1fNOi7wKTZFbKZd3HSBuiEdq
s6kqK+KejjpRLcNYEADDz85i2uT7FManP/bse1uvNlmkBNKbtHf0/lOJARPQ3oJEXQ0o6yeZvGT0
9YYbTKp6kmfKhU0mc2vLO0wRe9aWL7CUWAwuhF9hXY//eRy1EQONgRF4KpaReIP5dZq1o1qvU7MP
7vIOrcEqjyjsm6TnY7qKPoSUc12wj4gKjsyc2k4hrPoaGuL52RTmMLhoBlUtPwFv68VflvMsNtep
6AqlFKEgDitghyuCy1PNoBfRODDQQvhLYjDSEzDfhtnuCNgfvGCLnUdTlfy/fsnF4aZUKg1nY1mz
pMCfeMVBDb5pGrwFVUJJ52zIHNqLlXLPH70ko2yFngBi8q93VFGkc3CLjsEvt8jKxEw+bx4hqcoa
hNv0pyFiG46O0FNurWl51NqiKQd36MBf8rolmIa0TeCZm4P0KJoI2nb9Ma+0EjDxIc8uKInFaLS2
DkO/JvCv23TGwUucqRThTeZYQcwLzdOfZVhOUogY2wOU/FIFyYYkD4M8xuuRMs5E27i5G+M4qUAB
Jen4oBzTVfyjN6uhIGAqk+6n6+aV3Lh3+3MjZO7FfO0HMUY4+nkr5S2LJwiNhRpRRpJYp+vOGnHy
km/7ISo8NUgBU4BQJScBd7qNQigeG3OOnm/LGT9X55F+UuqaJdBWWTJIp+AEHVsQG1aBdyFF3NAv
cgUgyHG+WUvEgoP1vdEHTLblr6AG5p7+JR0w92fj74bvm+pjWwX4+7UZ+UAzpNRcmaCaJb1J3DNF
F4mW5ovhwqRSjBHVJXv7LIpfEiZ70xOPFSQRpKxJzc3DWachF0s2YazmXuFRrxzyqN7kbnnhbMYK
VACjRqK8ew0ZqDXee3KTxifRGpzoLmirYN3GwE20Q/YDxQ6y6/9oEDlZZ8TGn2C3wB49KMVzKMhZ
lC69NRvojW2+yH8IZGV/ltRW87L6ZGx1jdqJMYTZcbdxEv6Va4rO4Y9J0Xh8sYodhtXXHjMrAflc
9gtxkgL6IGAfnr9WbWGLKhO4Lxsx9Qbm+FubnEvhBDh71dty6fK3GM7tSBRGNlxRQTP1PMfFwO8x
3ba6KrFfajLgnjniabXRV57vN2XCRVym3rblwrCXPQu+DwfvUsiOMrgrevgrX5evBl7KACb/U5J1
zAJv65vzBFpvoveNb+y/m6LjjwEj1bbjaKIGimj+cOm0c/U0mkmi4BkfxkZ4m6kcqZks5SCNecH5
4qNcffnqqOV/kwoRW0wxIW9I52e0UiSPChd04nqIsMBfZr9SZi8tvVnDYxDR7lsJj7IGHc/Mh19y
KgBEuGgCiUX6pGwCN+f8eGgomUuoW0Gjbm2ZQr17joAcLIU0plf3lSvxfRyY3YBxXuLJgzLYXxPw
2+ClPhIIvUzv+NffDcocnw4Th1YBnaNhIPSPyoDug58W9Lj3k93mrDUG2tY7IfXW1IywJiQPB4aZ
/eB5RnhYu+uJx9E+MqHn3K+TEPAyORCFkHkwAdsIfF5UxTR1cfjjskQVZLz+Ftr6b/9O6pN0YpNn
mFOlDgFk2KmThrqpw5W9MOjOSDKT9UuH1vxHe7OGfPldCIRR80C3L1suWJHfxE3FoBhp6x5inL92
6xCRuSgyLndw19GHIVmzQtqTgT2GHifFIc2LrKnc36asApfOS4aSlrGNVJufHKWzaVOc0768C2R1
FRfm/dWJBjnZm9DLoaCwpqyu4NQo+MFJK/jIKyr5yVCEyCv9SrXk/Bycu3xypYKr/67XOB0Zuh75
WqUyybHYgNadUt+/8i21yi2wEp3hzVwNgC4sJ2nRRJuFfVgZX14yWEAQL9EluLrj9OMswPaKieS7
clBHMw/yTaL9MyDj1mDy//ZTPjvDRJsb5uO/YmLhp/S4u8W97rRMH2MkKY7hK+jf0+FjrNEuxPhT
6iMYI2PeGl6vsIdtLrVIqSRjqQ6Wf+BeqCZRgVJ67JCnvhr3DNJ3vH+74oLz+5DQ9STZJcgnEA8c
IweosIhAcZjRC5OLmmAa8dQ0napWmOLv6RwCKDelNKCLcnXP7cdqVS2cC9gLylwiTTOGZdAnob00
QL3yQxBDiJELuRCyjYQeYAqzLAqaYrZe1S+McdSWP2Yptt4f67ZoJZjf6peGEGmLnj7uz+J5N9Qc
YYHzqI+RxPcKuy2qK6MKVrdQUxRd2nVIqbjPwOAO+hbj3VNFEBV2BVnF5IKV16v8joE05EEqmQsJ
aMmwPLKDoAZGTh5f54KYeEgPGrORRVEo1UtXTTXTZckU5roCLo3/9FGqgVKGt6FqrSarMSH/fqz6
BUrYb1nTQOqlCyzWYrdvXdoQuGqsRDun75xRtVzVvriEOTQt3ZcLkql0KRzil5pHSvToHEK8F0Nq
uzg5bUEdPnhqWtWXduS9A32poDl6TeXjWM4TuhcusDouYFyIHt+SbjQ8QMxQI6xCVlTpsmZSjyT6
36AvCXoTr9KdPH1fR/+eAoM6pKcmwhOs17mI3NWt8D9jkHxpDvRXChPcpw0cABf7gtZDS26+g2Yf
hXQvvy5dF1bsJlMLIV6E6pbsjRqLa3946rpuIX2HHXiaim0X76r68hH51+89PYaNyDJkdu9PkNOg
+WC5rmKefzLdDpiWj80MACUKOl6HFb97oj0WvJF3qeXs8SEwUXwC4U7szc0pi/AuDo4bUP2mAmam
OP8gAW5fpg0xou4yjSzAfl4PCA2oo3aYlc3e40GgTGsQHKzr9ndUQCkI7/4jodwOedHm+U+NzDs+
KAMM9fVzLyylWgbLSkFZ/nYy6aP+Z0PbTpXHVwG/AlMkv9M1tN9MUvoGEEZwG4jcUR8f9RFBRU31
cbjv2XuFEs+2WSRsgi0O02HKj6aC0UdauHGPW6masidkAnUP6yY3oufy3Z92PY08N7AjJTo0GSxl
aD9V6qrAixTtKAHwQhsL4tpwxgm48HFriVPsPh8ktTl1sd7v10qbJNS8jnoTbzSry8E7G2tS383e
QCWGTgQAe/+IH1+ofJJNdXS9PECYzfP+geKSHJIdBH0kMXkdyhF25ZiwkbaQUGPBxKij/K/Se10w
foncIW80cT1buBU95TMs9Gpaz4o5zNUUB4CPnTOaPzlTpln3bdtZrwXX2cuLPoG+xrvcu4U0od0q
hiB41FoTi4oggXtC30t0r++zglHyXA+rpTgUWIJepnQQcVa6JLzrZVTIk76fswuasnF2XZCtDoUM
rmczeeQSYmNl8QGu00zLDJp6NpoffxBWhmJ4GO9IWiqiYVcgll1woV8RWXAkOTorqa/TagPz1qoX
UeJlgGsbbyiFQXPRuoty0HDVmmE9a1rE8BgPM4KuSoatCGLgTTF2BTT8eXbZ/swLncuPm7T0mWiL
90INkv6A4rWrQK8h1wtHAsY67nQudP2AzPkvG9Ligl9N/6bONTIDBigBjVan7zY2MC4shQIg2irU
aKQumegifLoGfi3QszLk1uW5fCF+zU4ZSkwrCBPgLteF9eoTJCDDLnj5KxWy4dvOqINfS7+7XHm9
4XBByYQ+EPf7Fb3XY9MsgqarOfo77t3ZQzooWLZg733+456FaNahlpjUlMGCxj9p9BIDCb3q8Dvs
8xmGRObEbS1LA/X+FBviDbsd3LCzsXJHTp1LCmTopuIBZObAfcTIKnYo9XOjyVWWXyZztYKfYTnL
hnOGCUXGyIsZ/lds+oML53yFWO2uQ71EmVxcRoa1lP+LdzWQuxvPf63WQOjoc5Eb7316V49gFZeF
aR4vUlUD8tCnLYaV63lR0Pwv2beIMxOF/6P8omAXUq8C3euin6F4PkKa4+2r7STipQNeiwMvDoLC
XUG3q/R+VHuLLaydM4uhT8blDKzc2hRL6939SCI2CDKSeoTs7XCo1wyK7eKu+w05BCR6eH0o6YOS
CxY8NZeUuHg5PlunR+P39mhJla/nGvkltBUfidXAocph09Ekzep14jal58jTSprjpK8R+wJHCmdh
SLpZMBaKktwdK+c/DnLR46ao9yv+nvDk7w30iRj7nf2BMvhyMbFWsd0BHOGtKU7nDKNsHdka0eDC
I4b+C0/exndA0LkMUy+JRxvdq5NU+ixQY9PvWj8xkXCf5DOuM1qRNtplXQhh3qy4ruidqez2IVlC
TlDFgXNO+QfMfIeMa9g1m+5EczlmpfCQQjjKdB5nVev2pjPoNLOVh+Xgmr3zbECCIK2EkwtVABdH
k7cLeucNSxxL5G5ejgAgSGyfrWMMyXsGyT1tOpO30anXiqyIVnVB+5sbAayscJtkHFr53/DcLKv5
u3Kreh7vGdSKvll0x+w8GSvnzNaNiv80tvrmW81sG2mLDxfq7yPJ9WMrV36pKS6C5EbyxGK91vI+
0g15r5fISFbC2sQ5bOoQBD+W3XAF9cx4SqOtUmwP9mO5H9qKM6EvfiAPVt+QpzfuG+/Knp8xNUPr
k6Vjx0KMvzFyMYpolLb4cTl4lq7ri5oAvjmaT4ajE0+ISUUCrj4n4Cp5tWm0z2d6833X1GyXgDmf
z1wJtoAmNkObau3KGj9kILmlbPDI1g65mNVW/tY0O/qflGATMqwNah0P61KQc4+vxmoonaiFwVLg
r7O+q9RljD9oCUO55GLPEbYSpQh074hKDC5cwrZjeMZdrWqRQhZnx12Ny5N+yUjVBI/QWhR6Bwtk
iENvFWST0XzOAhzA6pIwiWZXdks4dgDFnI8f1gDbPocy6gklwijpc7PIgMSOt78kvCWRBaknO6Wm
tVS8uXZdZtOAbqqudWrnfbZ+ByysS+oioxdfl4E0mgkhfuvmSsR/vmZxTMaGmufeQmb0KLQAdmjx
yefKH77z07MYPI3D3XtGs+NAy95aouCAHswvSJpR0NfaQrT7w5E0ourjfjaF4KdhNBOTEOE0vp/7
HDA5+ljAIF2IYSzYOHyfAOXkiEtnAgOk20zRH7KQw4427FKilkPrmV5bEskcwj2WHcP+92MKrqcC
O3pGgcEk4UwzMkzHoITTYwD4BUWDvWKkAaBCAPyn/duMQmUSlPx9zK/FSGEz42rHUtxr10REkXRV
RFoLBVr4aNAkoNtG5iqiGHmwm1xUlMxsxLG0SPBSHQZRsQEUfVB1gjlCc7T3er00aMYIO4H8PjPN
w9xUCp0mNhAtRa2UM75C8hDXei1vJuZq2EWL+c344YMnSB4KUd6YI95e1uVOrXg9iMqtsBO+3QLL
zJQjZRRMIAxRvU5CxK9vYV1CTkNu2AzEgL3i7WYJy8FE2q63TgChDeWGUiOGoGm7F8nPLk5OtA4n
aN0mnPGR8akSBwyTaFT/wdK5Mqg9oWI8Pbke+hW9Y0Xf1xMj/Mj1XJSqd3uSjlWgacbv8eya0lZa
7iDK4scVwfC3ppp+b2ZoC13hLAH98O+ovTVH5oh9Tp4Gu644rBiisEqeiI18eaPBokEz3n1XyeRB
4Txm2gp7QY0Mkhz4cXNOWVIFqHDj+MRBpBoOoojh5/lykY6qnaw4Hibbd6uJ++/n11pI6U4Twv2X
xuueAt5PSeEo9WC9tD1JqNqoplin1nLVqLH2nuHnYZ4obu2cZuXLqALrQbEhbwQBGNeOKhZNvQ0c
iy32R9Fg19I6DcVZ/rc8iYjsqLnaeJZcZMrgUSyA6sUqzW2eMHRqDobaRhSGaOgSq7Gapcd2hcGp
uDskmG4m26eTwqNTqIuk7cPaFfJtJ7QxezMvq3jebaDymel8Ww6LdU4n7gCgLTt9Etwh77Qvvo/P
fqsryli4kMUXyIkdarqET8Isv853fEU33qBK5rAawEGQtAa2T+FLyUiVPBul4tGiUrNTe1Ix3bZk
4k9sOiLB80NabogwescTnZAp9qTuutPmqesiL2/Z9Uc50p0Uk0kwZkseSut36WZob0JGXpln8bQu
EHZAzPvHgnsVxVFTNHHA8b9t5wCWeZLUpM7dd8V7Mg511MzfeBg18vjzvSTis7gh1fq1XDijR6Ss
ad45mLCuiPX9vYDkrPDY8UAyUxwY/W0v92gEAT8+oDXGAtXtXCAA8fFZL78yO1O1Ny/b10Vxl3SC
8jdB31+S+Xuezzz5rnKIHzx8lc4Do+osGsoQ7x2MYFkE03DM6okwjpsH3uSrjFB4+l6TW7b5mWJs
MRTyo3mgplbpM8Gc5iNT51OpoDa8y+lRZpQZDbg5CkMXrLXyQtUMkz2AdifBqbOfTkf4Mgmd+HwJ
1MKWkIWcpQf0LUAXZsFIdLY9rAoz6FheFMMu0MDAN4OshxLCkALngD36WwBGK5SPXNeb+90yOeCJ
rB7hmD/YP4s4uY9rLUwHwI+lNZ60R7TnfneLtTfobrPE2wSSaJUfYZZYoMlnT5FRZewLk+UBY4Uu
//FZcafDOUq1MPCHfPdV1ENCbzK1z/HPMTtBz+nLO3JlSE0qaVjN5gSsaZtEJQScVZSeRmBFJ269
743058Jmy8t9S9heF6Xpn244cGeUc/+Usv0LGkU2bcwo+22xFPrc8B6DEL2ihtUoNY2u2sljL84v
8T7rIJCzNEjwcEzQwtGWeI928ourAxMlOfO0WFowwoyKTQEpJOlhXW/w5QB4xu6iUhvzuZ8aqfyb
4s5t+F+TQSUou4sT+EnzTHF6qEQJtCfq92UVlrhUObK4Vmp27FLz6WfdD+r9uDWllFH68QD9sS5x
z2kSf9zq7/nCtQVGw/KPg/wGO1diwlE2xzkpiP4zlX8M2+yD1FJtuZOFDodJ3WBlOdx2Zk45UAy0
PKId8hca0978+QeYbv3vQmRyXwOcKlIqGvChYFHBovUUeaDIsV0gq+W8DwnfoQgHxESBcHKMz7dV
rSaNaLorAl8qz3v3PhjzYnvlHN/xtd2/4Jyd57eCpD1Ocb/kUUWwtIVCUdt7DHv7nWkDK6PTiUa2
h8VwDfQDE0nWtPo7pWiOlJ1YUyFXZKBiYXocJuc8j8OLKnbeECUMA13e5nE33L26w+7fYAoZURoK
/SrhDBZmTTd2wbX//gDi6Wc4ZwVOLTV0jFBcACKoLMwowV7VTqtoyw7HZH04zma/nDClDK9KrcAu
fqzv+M7mPPaUyqdibLzlqJ23mbx39HXE/LXCen/z6Bt6kYqS4QJiNCtjhA5oFRcyZplpeYBPR0En
pxKvS2Da90X6ts4BNX+T44dqPD37G0pUyXt0DZS066mY31ReZ0lUVy58+hzhCsA3c/nHWn40poyO
hMzVprlIZNT8mKB4ysuF5LOKZWM0EgzhVOCSzmnNAcDSWvNVYJtMbQwJtzmOy9zxlvuT1QBWcqre
ZzaaiqBp+RwQzefK6axAdqAk1ehl20a9o2oRmELpT9D9fP7hN6T+9RHINtXwjv2T2GzqX4gMotK1
rX43F7zZLjTZFylzzAfpPRTkPxdEj+OeYTATJwb42BHV05V2rqZ8+JcT+1QyPs5aKz01rzXqHgY+
DkSoF6FoQPy8MohZrjXMyQ5HlkfUNelvsVTZlgV3MlkusETOHrBAqE2yEm0tBxC0sFWlC2sxKq5k
aqnqXysv+B+e/bWoFhX8ktBJFyTpcsigkQ4SUM4cFOSS88VwImA8MivgLjX/FxLAhjyaEr/JY1wY
93mA+xNZD0Ff6poUWlo9xuAKumlEcjg71yyz8fd1ALOmAfMVv9fJc7Phz+P0ytr0kJTWyE2uuT/x
bvf510kt3TqQNXXJsM1JWvy9+/3H3XMXX/uogvnH4/akT5G8bV1jmZl7QNChpgeXZq/syooTc1DI
hhPoYsqrjjTlxcacvY62qzm13LkwDkPXNwQpudg6Y6dG0OPR1xQKT7jAdg5+74Q9H7lCxMyuimrI
XPjsGPKzCJ6tvt/LyQrQoUOS7klwtQkldkQvrDLHd/6AcVXLZN1O4gxbkY+IDxfs2ySjaLRlMjKo
pI8TlhxeTHYtAgRCjtg6gzC4g0rhrtwMP5jOfQB/6vijS5RQ/KDzKx/RB7H12APvYohI54L9pKba
fAtMeAuzH8We2/TnXQL9cc3ERjmkE/85XRG+Wc5T6DZ3ZjueTUJFe+k8eRGwUcd13IOucGAXDPyu
YqxUyX85x92lgrO48CXB4okAYXSHHn47+m4lACIL2EfcmKLjw4INuZunbY4WdKbHt8hymiMzR0ae
Vr/8q37ZFEoT9LQ/So6bLLvZ4fhsOuBc2L4v5oyFVZfSBDp+YO4U9f02il3SsNISkXfgwLHrN8+4
okBYY1QlRHRE+4d17lNu4WUiKB7oxHYLZwQs1xhkOnCm3xPPU9GNQ9+PMjX+YjsUXdT3E65QVCbK
lcKNJxmr8Ad52LxV14zM4oSaLbSf8lmTICurGJfIs5NpOWAKF32KnmOWI4ElBw7G5pU+h2Klj94X
LnGFN/b+1QXt98ZXfD5MCFlVistvjU91Yi+k6UDltFaeOQ/OACtIAPOuPII/eilRzQ1pTtRd+gA7
VRQGIVTLoGNmEFr4whvr1grI2uV8XhraREAeUqD/gMDjcuh8/7jPLRturgcGWTqeC/vFirmu16vR
A/dOc9fQ7pxJah0IlsJEBoUodsIIsnF/8h79sq52yNOVfD8tCmDgdKh+jrVsHy7kFQyRVFcupCMX
FR+rMh2SmMpTjZYFFQXRk1dArMcX4hJGmZqeiNzLfQIC8aNTiX/EoEB3CoYUBvx3kLdgatp7o2f9
WcPpeMv0KJyBJLVWmKHfdHXX5RCdn8HQfqV8KEzSXCsleL4OzhyD/oDRrAN2ES2RexMLOgnxmq+A
MSCknpF+zHu0yDH5xMsfXoU1ok1HIU4VYqL2jRVG+B6KTzJ7jJTyq+rK/6aedoLKDHsKHqgiY+YI
49uVJyCwxrM++0F0w6/gYdbnoMw/kWnq9P0guIUF3srQhV7QQ3tPeqvhGLyiAZX5do3JdJ91jGUp
gPRwfXaEcG3DjdO08rC1sv3FpOaLE3LnTECUji9V0+v+YOuxKkvoqJwEAztnWLoVxwPq2xiEYyi0
GM8XCd6fQgVn5jiXdpxO1IfKOkAbKjn3Tt7fZF23Ujd53Aok1CTy7EnL7nNFwZYgGCGdBs9a+Ho2
LRrZtELO3MQBOxfxiwhGm6Q5dGtZeMbLbDaq44ZDh0NcvDVCj2DNWc37bT3G+TNw2NKb2ssCvZhV
+BO8vYftI1kQTQ2lPdph1yzgOx/32OxI91dzDqsdaAijsYrokVYgunFEko1dfC1pL6Zju0YAXdwG
iB6YFVDnvK13Ep7Fq0+b0YnW+MRryEbQKE19st3mopPgeEaKsgt7wPbRLXhWDrwp6KsOGUyYoJfo
5AFcH3EYhV2yr6eUOW/rYsqgerwgdBur1C9okxDAVLP8zFHjv2nva75QGK8WIdP28pGhnro9ZxjM
hkEiTmNky7wqrKm5OwuQbJMwb1ZDS+zHpp4odU2FxXaxOm+gxzICZx9M2R04O1XgRNRKw9MjVPbm
g1fQ6xxRq3+q1/Tls+xlTkmwNF2yZu7xuWl7QHP44ZxL80934wD8cxt8oMr0cJLRu/LhugnoZnXo
6/x73ruVeZedDujmc5WPiguUsdUF/WmJdwI6Avdi9NdBt+KMMf+Qh9bI/N9jW8egYEJnBI4w2BDm
16AhMII90PufDJMdgBvK732kQB7e1eYiNcCyD7Mr/lB94d2gGkt+to1bQ5quJqhwc/0SmfiVFCES
b9+Tppu8eacxcPI0fG9jlpN4L48R+TkYkIAdG8OTuAeKAF+nvafU5gqNzaOxYST5PzeROFkV2Ych
YremkjHH3PDXtqNdKZCY8kLGAacjAI8vxFA2w8gvkrJzdgTw+Uxka3wE1Cc0CpaPeZiEOC+G/8e3
au1M5Y11PE6VAl4XNndtGKfRvNCftV9Z9eILE+6r6WCPmTt4AJBINA+S6Tg9YJfkYE7Bg+sQb2sB
WahrDuQDnJ3MjeYzpBoINneWukYgUYSGbIZ1257+638iW6c5ypixg6oakVxIj2p1HD93VFP9CajL
1QZuUXmn3a7hxRd9UoC+iNYpG/asy2qC22EeU24r0PRyUqCnD1UwHGJqVny178LFg6ziCY4HTHLY
aCRMd7UMGD/2Hhds+MHq/q2Nvdwv3hrRvX5JDUQBGhOOQW9ZuqcOFQVftcsL0PtFVrS8kLR7TiyR
nuzG0EzNF6j+Fpx6/zAzA4r/FuomNvgM7+VliORWxiXoR996V7JnRjBgJBZ+gXl+z8g3geVy7Y0T
26lzndzyKdYynkfLNp/GxgLQ0KigvaSGY26HWWpYWOo3RcV64D0Zftowix5EODA1uBrDLGR24JXT
2SxyU4eM16lbrStsdgz9CWxaR6L3V6NHUBabiuSWAeURdibBW1VrrkdYCUrPlUCL+wyaJgFVQ9bo
XxyheIQ/qDuqju4L5nVVEFPnPSaAd0BLKGTVQ1va5yx8TBtoVMCXOp9b8motFnLb1T2eTkmEknMy
u+mmfK0y5dPO9ja0R9/YRWjfhJo8SmWKJWhJO3hnarucECxCcGepSwNbi0Jqx3JxIo5OEkkR0h9Y
oCMbnTI7xYO8CUnxEoIo/qjFmyzJsaa8x1irhYVvvLPjHQzTEXoz3PgSOxocXosC5EM0B98cpvpy
/K67w+PT+3UY7zF1EJFEFEd39LriovkpsRTIl5FAmRhSNik7+yGytK6BbhdqFgzg2sXixi14/d5l
JtKKlAvqE811WUaJPrkAUYWt5pJfc4RX/Wontv7aW0HyPA7hwbiQpyFwC8tD+8j4raUf9QJ3YX9a
dVNTiT99Bp6UnKXHAwwLcmuRTFgAdlv276IEs9itTSL4d8Y077wcHMQAV1/4qV0z8xapA58AAisd
Oy/iUUZdettCwN7L/XY1vGely8pYnXWlFFtFQBOtVRntUAoffAKTmy1qd6Hmqghp5f5EwCc/Qx4P
mnavUn9mKCcehqFcJeutPPeCI1Xsz4AanhT8pdfj78sIeKNDi1AxeIw4ORCZIiGaAl7N6vaImLbt
pAWKn0YrRqSASa7iRKNIZeZ0f3yRtzG5zeeBbhQSeqQC3MeGdj6B9vWZDB514XtnFiGna4Whh118
K5E47an83SZopll9gSPZd1JopnXtEDcOpAE/iSTHGG5NDN7bvZW80vvTfQmR8hfFVy5/tO+SRn5V
BKpoLuD3G+HcB87kJVrQyzkwE1WM3o3iB81xX9gav0EO8hfThCAw/4b4aNL/ror5Ws/ZBuWl91si
bmEyKzTICcjtg4Ai3mwNf959fUoS9KSao/wfGmMInuFRYSYo6hQDlw3iVJ5uvi+Y8HLP2ru0i6NB
nzwdhBHBgEfoQi1pCSZHGc6Vx0CNJWyb6hQohuAOvUPS4x4nvwLPv3u8ro+LBnfqDWNyG4a45C+Q
7LXqom/yA+epMQWFC0zra69090rqkYcmFxN7rd19ppjVPzNlDin2K1A4Azbp0OEk3QKOn1rgNbIx
OJQXkj8uhNIu6l5B2tiI1D5DQo4qZchlSFmLbYUPoYBZTsUoEd5iKL1yJg3ssGGyAUeMuG8/UTQS
eVrKJmPzraUAwg48qOKxwWOYE0+d0Or0eqZg4Fx5AqhyFojIVxzgMdr8cPmPDaJiMfY8STX26+8s
dFAwohttkrS/KGyQuHoHHEhmJSCF1/CAFD8ymIQgVgrrR+ZgXhgb+VBa5HPEPY9TVCzcAYWujH9E
xgqRPpNZ7ffH7jwkI/zvTuYbal6ozlJJYC6kkByD/1ffUD4qyOAr91EZa6Qeb0Cg5VNKzFOG9TJM
f0x+xi/3CWbVlwSfIivNzaF5PRpXNobMHDTCGQwUnmkn6Rbc9gXMMahTTJP1EbNi2Z7KcN2Bh7B9
q3yUTW5eauVg8rHHaeNSY3GOnP9oNJUkM4/O3bBmVJ2TPwh91QHuSSofiIQgcrm2ggasDTtgMepm
cqAjIqKFEkok/kTNRFDUKdDsOt6Kj1RsWHlr7Zf6c+aQ97r7IWGtncir6dqYKISyxiS6JGF4K9aL
vqISJ/lVuvHX2lCdotcjq2P0EJiOjZlcKjHWvxlIQ9vy1NtaPTTRUCatxF2lMobIo4dw5n8IeOJs
cKscB7WPpkIA3eN45mtrAyffGEMtgKK4Ysq4pEOT1McMVh3q5QZgP29596+z85LcEg1OT0lUnIuy
zr2qTgk5/nmM3tc+BXTQ1tFF9NC/ZJb/8oXNzOuXkUDxc/k+/IU9HXwrXnNyK9aK1VOfLFNgib2+
LNfMtndDmh1/zohvvi5lXA4P2b324/e31rwS6S6gV0D6HnorY7/boYzWIu4sZTisE/R3AT4pyzA2
KXUgFYayzVxKPkKGiiNIHOsnFo9LP88f4cC1e6l2tCRrX41nVJZ0OY8VM+ZQqjEY4hx4UEQBUfKw
8YtkPJ8RehmemkZ11LZmiPm6nUzFRMpxvKHd+/p+OWe4eeJ4ZB+F2BmO/NqvxlDo5MgeR8oBorxX
u0fvuwsZYX5we91/o9DLIp8z7+3lpLgw8H4BB78QPEz2gRn+NCL1ah79VnQpzTWZLtfe6Ce1cTAg
w6gUa2JTnQjoCLZ5jPdE3VfgD6QttCxBRMSSQEVKB3Yney3P8CI2Ff4RlFK7WaAqqMViD58WWarn
gR+ztsvDORo6BSqmndRD94gM7cwdarasxYrh95wqwqIxTNWf2LUJG73ohwD9fd79tvyO/lQf84it
ZLi4m4LnGCNu9djzboM0PN/SkgABjJHaDZrrGYjCwsgEp/XsS8UcHFLaUQYY/WCbbLxKFwhJwSob
zit4C22pwb7qZFcYo1qwFlApAr1fDjlvba2YEG96aroOe76hIdtPfp4zPT9bQmtugtVfxcbIVrhi
9eohBolnwHEMWf8VG+Cfak9BxWtXheEkyhl6zJ/HR8LCwvFipRDyxWPXLZqxlDy/qsz7K1RshC8p
8ceAKUOeXr5VSe/+v3m2i4XrGZGxIqf5CK4lOxA3e3YfT/XlWl3U2g0jPbB0dndHEBKHRcuRZHgm
1D/JFkxFGL98CrrMpXxN7ZF1p6d05eGjgQyHryiEp6AG/4fXACuiGcFOIX8YxlmT2aEAxebin940
VUnpOPJw+4TmeluywKF9tYLCLmYfeabSDzIEZTSclvcopR2gSSXIC9G6xI6CQNbD/iOGjD2WJ7sV
zTXdrRi3UcXTM3VD0sDPZE9YcXQbsYcR0GOF44nrN3+FWaQSBwQma7uAZFHjLsWqn22JfoOSTDNP
9GncVk2KUmMY9GyMxyIzi1ZBVu/qU9LxtSg6GkLW5i8c7a3E1hAo0IaxugI0Ve1K026ThYl6jofY
6ETPfISx/xZ13m8jDZnCpuc8ktoAY9eKHUwFVONN9RDqz6lf0bgpfyYEPcK7RxuDfMm320hGX+HZ
2JKY1QoMYqk0IY5QOsRZ06A2oc/preiU2CBizEBIXqXMb8HY2ab8pa8Th5tFyvKlAgDRL4lbLDdm
L3DJRjpPpYgerK7ow8iuDM7QXPRJFm7x5ZJXnFn0plonKNT0hXBoMI95sjWw4L29+W439VFY7Eh2
X35LX26Dwzm8ouCJJSah6uUwTn0aiN9GGAkNqO8eSPXAN42JL63QTXHXsmkmBXUA7JdhHZimRM3F
jDRWGTcpBwa9cX1RGlXuxPL6M+GUDZeMQYGpXBHZD5KXOJgLHox9fvMeF6r0mdtqxjGET65PuF8G
9xVQ0jp4Kdue5w00TU/cd4mA1N5V4eiAuF44y//B2r2vCYfvzJxcBayuLLlhs3fKwhoKaL5vlIsS
Jma2pGUd0d7xCmU/mMumHHhAwzJqFCQi3Uy/uI+NnHBnkWd8d7l+1yIlzJdnwgKtxDpcs60nH8DL
ZV01gjNGtUf1YBC2Cy3tCVF6chQ5TLKUqfSKmm0jbzeKO/3saPPZYLhdueH7CkHe9YcCf6nsnOT9
dOuAsWN3/AUeVdq4V7UPNzX9rukLsl1q4nUClE78m2iGYjNMoT/Ucz17ytNc4imu9P2YFGmzE+ZX
eu5dzb7c0epjj7iPJ39RoRQRXeqtCooB/yoFvr/c9Vf4rldQXeZ/s/js1YcHqt1pcM4W/c7ph2qa
/VwAtKycHdCLjIn8wEXkfXxJX3lsqYcavtlqDQnmquzH1HZhITT/ry9VnULpXww5PTImHKqvM6Aj
cCe3AP3RIw3nMbvy9O98hGRqxz21tPx1pWsl3iAn2AUuxJspCh4TjivLTacIp1Ld7QGcMmQQBjL2
MB3degQ5xZVAyKccnIIpBwAm2A4oCN0s5/uHLUJ7XBmgAAWom1mg1TmCVbsxYpPBpfH4qQM01Tl4
yjN274tgu6nMdH03vQ40Wp0Jv7ZsBhUC16BYcXS2f6bEcWG+WCjHnO8cdHiysoHUrd7VJw3GBied
Kj6wFnrBCiCX+oB1DrXLEv/Y6Gnzzf0cGq0PM5K33LaDL4ktT3SYw7nb+8OWnHJFNU7Krj164pPT
TIt83cUyOSipXYaHwtYB2Lp/GK/PMbxXImO/igBL52ReXXLL7G5NjY/NtkDWK5n7agELgmrkCsr3
PhLmQMgnXeiYTw6kivBJgzhhWSwvYo+JFUsC/a+8Nud+Dd4ht2Bu12kayGIbbFxVHkuTlmp/vnpn
Vhosk4lTRTkNSsEtMXXlMxOub/P5dRwYGXzyvi1soNQkxzuqdxmp5zbZcUlLUugwdX8hsSTzNgTD
o5Ib40sGh0ZtIwJMV1TUSqke5973asJ4p+eLornj+FWWDyx5hw+SMTdPo9klcVReMdG9G+FQoKec
m3/3y6ZgtOyeBpzqQBTE6sanrJ+FukalkkepUnWkJCDsMwsBq9xpMRZXySV9ZgaI8PzHDbuzjoYL
ALnAXkKwo1tji7lOjfenwqbsGwJjx0sxwQQfzUM4jQ675B02lspnGHflvUq8g9o6p5Kv7jlh4eik
DNCKpkke090Mmlkb/hGOduEhEhAu5fANAKRVkLfAJlgyi7Lb/gsVRO/GjMSq2DBe2VSaTo44Rn7D
v7BvqOI/I8itvjAPxc5cPQRD1jOSyuiAmzpTp7fR+DnluBoQ/Tb+xUtzo+QHrKG758XQdmfCCxfB
HEZQvAnqsieYMbdRE6gWdx9T2RvyLPCpDSP5uylOjZu4hW9I85neBdly453OXMIkUBPnW0gwfctg
m1cf2NjLg2876dLHxU3KwdmWB3zrzU/QoEUYul+gDdq+MPZfJ2LuY2WetuwXiuVPJRG9I9KUN/8L
jd2XJFOwsFzY3IXN787aybtd2a+x+ZKe6vgl2w4Rbj01AgzjSI5iNxWeTIHoRz1pYkFwB7mCu62T
pGlOOI5FRsZVZYJEeieOd556eA0XX2mahZRpSWvHj/aJzJP6La0eqyN+asMqaR7v3gAxX4Sy66Il
7kFKwtfGS3jpVaUStLIUD79QwSiHrMGv510rI6u5Kpc00teZEub5Pn57n+xd8MinKtFxWU2PIGIj
RX/tptzR1nj7XZgEDfbQCF407kzojVcyzDzRtKAELIPm36+VGLsLXSFMK7ybNL/8sPEF+cnon0X/
QvywxPRGTY89KMgKDWfTQeWkHWwA8AkmAfvF64p22pMWxNioGfSghPeS8jqLT4fPQOYzXJSEwqpU
5Izo/KwJN21y0ceMr6qQgJNqJbksok35DIkWcbRpswGACm1UntpmP+m/xSTzefNEpBjqRrOgFG1C
EYSviXjdocLNptqzBcKxqDrZXEx+aRgPIIOrbtEjmJNmodpvA3gIfDBDDtItzHiJLHL3YJAsKpeD
oRvHSQiIibUgr3JA33UkbpYiPLVA74Tx69gw1rGH9oZAlMPVuGtRyyrYgSGYO8+52Q+ANqJkn7TT
SzJbKNpRdZK+lvn4kf7tQwVxGgRv7jpKt0jYreieQ8koNsjwBzpijZf8IZ9OMpNmgiJrdfpCWuNz
yqiDB+xFLEQ5JnWeYNW+4+J+oyPjjk8iW1TOUTb7T1DJpWbixjf9byseuo7IzPHtcMvWRSD1BjeD
RdkNXOsE9xC6Y85Rjvu1ePMxWzoF+2JFZRG6OcNgvZiHbHvezfubKB/dTh5LMF7gxPav7pu5qF+r
8LIUwNwBMTigvpDTlbesRkReS1y3a5HG2d0R2krfzwdQJ+A0qn8RBv6RcnJJ5YhbGaPVXfLDRHaj
BgabbaTteFhWyN1VArGnc5VChrx5N/TJyBzp/3S8tYM65jK2Uk8pMnwCwuxAfpc5WOCwkWHFcbTF
TCMv66VVCaR0v+NCLBmgLKFArIoN2Bt0yGEfbH9Q+dTgn9czZfkn+QXaqRClTc1WL+kx3yr+tVZD
aKtzjoHvQm1l7ko3BqlwM8rHX8Kd3PGYUt0WXwBTXFqjdWm8K1tYh99omleZph3rdoYqfJPxmlBK
S5VkZyuF9bwpsA800tukP7n0g2Gl67b6ptSiRgIyc/nXK6swJ6UfLoue1Jq1gjXBkibHEXvfNobF
55+kutP4ld2HzSt/vY645mgAQ0euh5ZCxz5GV+xA+oXMy0S3cI9LtKHoNbDqQ2OflGD7XT9H1Nuj
ZrZeCcJEHZZ1QYbaJmjjZuuGQLzgOVNTtCAp0wOO0gGkVF4ccEU2nozjvA57k9tzG3ZQ2g+bzUYr
J5iQcPr8cEvhVNtUh3qOt1PH5K0PMWwBZvZDWaaN0sZz4vdmJ69qc+3Ofw51iH7QZEZ7K4FYrLwr
u4CQ9Ws1QtLoeFFXnPNe8HPwuzpZhLE+mRKx0WN2CLibc7yNWsEuJofdDbBoSbFOi+NtBqw8m9K5
7RWbHsKtWU/LWcSXmCPOZGoG1MZWsPV86KF27jcCiZqjdLlh/ZRJSomWHua+nx1Caetnrud3s2F/
st4dzqAkMKEsKJM+CM3HWFXoMHU9bv3PfMUEyXZ8TrDITTPWBJI8V8wqx9SLcGwHneSZe+71W9DS
f4hOkElpFcFKA0u0s9BjpRmh0zj8T18VhiL94VoK4n2m+M6olBlKcN8Bikmc/nOCxsT1j+md89gY
56mvJLtCQBeKNF8Tp9Jd89wavBNQHHmF3S/tLg4/HtncR1vbaUsb40nhvQqpk37PlMsrgruIV/VY
tzDzRXJ6aLGSoys9+dy3h5QEUaGkTVFISwUnNMBfdQadLh1ES7xf681PlohcSqmQUUkfQ/p9Epld
OuLVPcV1KocHZThw/Fpt+9JQDQltHa/BDxZJoL2FWgQAE+VBT3+YMORlshGDVV2CU1djNj5CJicV
BsBnIUzBka3uuUq8md5SO5uMi8Y+N2TkvXrpK46RKWE0IdJ3aaeDkhYTYjQ7yZHf62T17gtfdeBL
Fvo+Ha1+FoSGw4h9m2Jd241zmWS9uuX/0vmteFG/ns/vdlJpkmOdzcNC9L21bZly5jdeKK6vZztO
V7tWMCONwepZ1kFJsfTjiKzH7zBgajk6MgMYD4bGtjfFGWgG9K8w+SCtJ3RM5pp4ig902SGPEC8D
pven4jvGb7jjEoKBrL/FmfcJMym/PrkhWlHNb4y8mwLBNTOi0A/PVxi0Vnym+l2Jza/HgL5RwqiG
aqoAyiqKtv5Nb7Rk6E1xIJLYJ4f01kuH+N6dkT5GVUv376Zi9QzgdRo0c8iSyxVWuzk46uvzWOlY
LZ1vIIRa3nonP8CrXk3KWj5H9kyWj44DwNrYSpwU/O4iaHVqfDP9BAXXbei+5/8Hk7hskWyhWKDA
OBUtWVhFrxE835Ve3E8pbfZ/Qc6b3UscO+0XFOlybJX+e7TpuxbLp9oVa+qEgGPmU2eIVCAGEKyW
C0ZMZXw1aDhtcM/tswphoVmVEmBbh2OPv7m1sUwISkrH8vrM0PU02hw96sjVnLdK8JqyNwGUyQkC
fLDe7TqO6BG4nLqEixFYhz4ECSynuKDUwKagCHEm6jhH1or8E6ZMA2BN/VtWdmOyBmZLFWnIfe5X
kTgDEqP/OVFvKp01wGH9PV/CvrZSsGrULT06UDeU7atwxlSMkTq4HzsmobOIzihB/h6jPf3YWdI7
jYguFFQQaVSwq3Ae/UO6QnVjAX5QUmT3xbBs2BR4TX5Xo1hmFGr4JHsqSKSYWbSPcvNaD6J14205
nJzCSUldPyUw5nqHfToxOfuOOP/1qI/7vjMf3HnGJyBnS1nxkn+TITyf67qYMI94wT9IqjljKTI2
aPvSH4HWeyj1/Eq3179HtrvWsFgnrpwGA9Mn+FkAoRkEvTc3dFPqqahGjMYDB5geiEr4AHNZh5hb
JvtkDOy2yEQPNiPiqNCTtOqxpT6ZI583wpioq0d8Cm5k6yk6S1P14B1xOQHXEV8qZ6hrumdn5TKr
dEt6Imuinp0S7/7kiGe6PTxYpkgFAu+ryVGYmQpwurfnpB/W8CqfZdFJtKDhWpZS6mcGk0X+INr+
eIkWN/yPKzekFs21Z5U+lsB/YYCjy+47rBsHGRx8Ht/hfqJZ9WEd5L7qchMdFv8Ti/KtTZM9wwua
yYI49TZUxBwaznyzmtoaybUqz/HZRYTgtVzl46okoW2pJT8pmTu862QTEGUYFo2aRayQ9NqJDp0r
nqfbzp+GeUK0E4umdkzzuEBCxrMJGObKmmJdxNEHzUa2dHdpL6jwQMV0ju9TNGtHov1Gdp8c+JFI
6CLLK5/2rG/+IrAg29yfOEAWDyCIWCAdeL7XjnO0I+rqymMPdltp4MIHb+YLdYKevao7PNZyTjzz
WeS3c5kX29R6oLbUseLcq7niX50tiNGVP5OWSEd5fEqVsb+nLIdxY29QPGULN9RFYwb8qbCN4wDc
RGDyH21HkFNiYnT/RP+OySf5nCskUjebW/PnGAo+AObQo9lQjOFRxF27QXCikjd5rOOq5B3bOtk9
aacLx9W/H2Ybl6/Nsm9Do3gWkbdSplGPVgYsY/edOvDUFJh0MAsjswTRGfLB3XboO17pYsove67G
Gnoq5bmHwAOn78t7P4SK9veCoMIJ1fqFIayA2TnJcPi2+6Wo4vvus4+oS4WsY8JR2Yw7lN6Z3AUb
0PLX7T0G+JJEVr6z9CAtyK8JG+Twcc6UhOhEBDQi+M4Bf6Bw1GhTSaifJjjHmvfpnxguLhsHvUhK
k8CSAGB8zDb/7yHqRIJQCo5P9WSDvquueFbJOmSPwLAYODGs48gzECqedvK28lIy6/xwXJTaWX67
FSOp889QRAZOaZVdm9Oko4IJjl9DFTFj8RGW8Ugmav4HwYlwrpLuQN2JkIqyE8vh9FozzUcuaIb2
s5bR3yCQElNAz/JBa73ZtsKSx5kjbPxIbW1spGHpEnSRVp9DVqc8Mfwiacgc9hKQSq6Uv++wRQgS
OHfVwaUV7hUKz+Q+zGnr0Fhndk5W5OFDjYdq7oA+5BsdF8ypyhd6cZZVuRqzmUUVQvfJqr1oEXpU
X5qgxhqvtiLTi5Y/LSPp+MeHzqPgx88GQ36eyj6HhbuEyXaBUphGma1iXxNOj7DREmzi+lt++YxK
Vpq92EU9rHTuELsoJ3a2cTN7QB6jFQuLgltJH9kJmjdnFhiBEdyFDzxA2oI2FTA4Gx8nvdcPUMdo
GJCUnzZHBYSIA9xrbayQO94ot2RmlJKcySuSwxvi9El91GJBqh6mYnLNSxFL6mRkLy8GGcb//ITH
rkcGPgGBeToKf99nXuiA6/K67gzamF9tj8Max/DsS3bA4De3dn7xHDZLUW+kEe4NGogQJy7MPnzf
XBMfvyB0u2I5Qcat8JcE4kHI4mDgQ6eh1Akp0y7bV4VLxdZxTnGHEaymE0utyKAzi6KlOGKXB8iH
KxQXUQFFEWY0GRrIRd+zRYYhyP3pGSl246G5nYAR7XaT9KW/C3GgQoBCR3+hOb8zoxQHMCmTE5Yl
IcyXi8RGUnkWPfLv+zNqeykcQyp9BHHoQdn67/uY2x60rwynZ7HC6n2NTqWYVo6HY44CVA5/CIOU
d2kg14QxrLZzOjJWNEviP0gTezLvSjXCsixagAKEk54V9WY0NE2/cQS7Q3dB022SjCb9ASrJcjgS
vPcWeD3fD9CJc5IgeaGkrQh3V43iUZdQNbV1Qn0Tl33rUezpoXHDAI5eS4L9H8GLwrGpcr+6lVUU
4nt/5J1DTdrquHN6ld/UA5YFPUwg5HMss75zdffpMRSYV2svVeNklUAkUahmnlal/ei72HVpm8mq
HvnlsZh8qE7glcfgCaPo+sFeFixmEp2dnGot9zWcbD4qKm3sf9FC7zHqaEPOwgCx5qr+RMgPJmJc
etR75BHeWxItDFwCtcDe8axecbhPe0Khj0GXX32cZz2duwqhYK/ynWkclz+DbXBTILWQ1XVWF7my
LbIPqmIHrmyibvjdb98wzlVBbPFOaP1bZjO65uc0Plh48vltU3q1ih0Yrtx0/NGpT4IiZ1dzyxSB
MWFaU+cRG23Thih/pvIjjYdP0J408iKclb+XkvYX8nI8BdKoGF/Usegsoshbn4pj2pSJhVidjZII
+OBJoVSzbf9kv5FuqSx79KTbX2CfHMgYl7QXgQgeQaFxkgk41TynoDv4+jqbV8T+SOM4zO0rKhlV
G0I/7OpNadDDcNRDisfy24HYDwVHg9wHGZnYX0E/mdchoCi2Iv4C4oWKGO91KeTGOrv/ssrk6q/p
jJrbDPoEvvLbXdiaum5qdyn9VXzUXKWHDwPaNJQSNGnSQ+9q+EkswZcrhmIN/iUJi5opQ9mS/ki8
EdIEnwtWQ/ekigR5KPYoJHtYRrWmmnAl4FMUkVjt++H/QKYhbeAo5ClPCbsNa4yHWiYtej+drglP
WFRn+P7pvHL1MzZDH7kkn/OOcY2ATJH5uejV530f0wEHz+nPuesA93vV0w8JRZz/367+MDIZRAqL
dPMgHLyec11mokZAvrszNaL9CCZTDJ9vV1kaCXMVI5kIxaKua+PUi8B7nGi+ZlTJneNDLUaUDjPa
CT/cK57ju3Ru9ksNkDTcTEkqPZNupUDnHqzSq1i0gHEQOqcATvo+bIBmdjxugMFnYzAMoWUhdfaV
GzfCUCOguJAjlLDrYmZ2igJFJtUkazyVPJWY1rQaKhrGaf1aVmCS+hzrPyVhVTarhH6CiuvrnX87
Q31bgK90qCtYAZ5fkxDHiBcngAJzeN5XcaoOBlCYdNgsfosB7vUo00mSktMFDyU8yvaipxAguZ/z
dQeuTsk2g/jQjjpU2K9DlnEx4DnlCiPYVKSi+Ye7tBrcta796esAMiJ/yW0W/GvBJyigvwibG8yz
WiOrpMqLuBaHfvW7nYt4ZV8Fk9bUYAH00EWlUfWRpcJeae/Hjt1wKwGpnxAo9mKFtWSyO5h8Cr+I
XM/lNWSu3kZ7YkJlwVyyluUYcTexGu+hAtYal9b3HOa6vobfwyG93mg42Ha88YH6/9PLHK0wbMdq
EFRninbNUrRWBXf6zSI/+fpp7+N7GoSPBS/faSe92WY9FmcgHjbQ65RKq6EhCm2+R8BJdnpMOiuA
imFERFZB2Djfs9HfJzXIALWXgT9inhXxyka6z6wOnISNJ1repF1fAAOIscmsKEuSTnyIXJ2IeobN
XMks3GoQAbg3xjl5OlOo0747+JY/GoLq8/1m6/2qtDmRmluaa1Tg7PYyUt8NJfatMfBCSfjdR4Jn
sdT13Ff8P6KvrDtcMf7NsVcF6PM6MfiKsoTnNdElyhhtOGsHFcF3M9X3nbaEc1KKCqa4ux9yXY1v
LQXKHHyINWS/Q+HJB1kRJB8i7WAXalht1aXA1twgp/0WhtKfTVDCsSxjbd+p+TavAelKgR0jvJK9
6DrxzxD1/fXhryfIahtADmYZnfvZoIJqBmx4xQRsMyM6ZM6uZ8PJAj+GtIpLsCweHhncn+XkafHN
yyL8bldJNLnHBS5Nvx/7HZ6DLUCQ+c1IYUUV1mtNeBZL1yjpFYFPsIa43EZE8bzKVrRDkdndRK9i
SXcA1z51vXxh7VRYrJjiTlIGB5olsxQamF2t9VqGrEMbLOJwmdiGEAMU0PmtJhwoL647brgzRF68
gbI+JfyR4T+NhrXCDo3DgFgxpRPnVKNiUk+d7R/CYNY4Dyo36uqjfK204sEO3/TwklatdC06VKZD
MfHO1TzGQN2IsLB1+v/r5d/r/BoWh4Csbhqsm5Pq3JKQzY4EH5yJTTnpTy0wRt9O8pxWQnLoLJ2z
1aD5ua2f2GRJRAf8ljRKOqJ3WATd8OkPDk+PfV2rEjRf4WZLr7z0saKQfChdCz0/r8XE6X8o2q5d
U+y5a0vAVXwD56LhnRBmvYkUUcWIfh/LNnftUbXu3QPxjz2dx4oo9icpw5wGCP35HvWSzCPYmeSV
hKpCwFGelDg3uuJx13N4mxXkpv+Y3ksvQKpL4yWMOxijAEtH4P2pM5z9OEJmL9pdje+NCn7gLpe3
FjNrNW7OBv+EJFviUQmh/byTE0oUsC1RZYuCzY1xZNpDkyv1SSNgRZZgTUl5QP9aKV1LI6JxxbCZ
dJkvp7TOzlszuCbvXqBxZcnaPbUpjq8XYKl94G2apajfQorW/3Xwrwvb16JLWGr9jsBPTJH2czd8
96wmv00whjvhNDouszKNW1ViFh1iBhdwqesmdHrzWwQO0fKS05KLAZvgWsGCY3oYHVPUWexjIUAE
SXmPCd5HhVL0PeOVoVKELLESuxTj9MVLoqE7uGcwN66in4gp4Mgr16fo5aOFkjtXMpSNxZLz6oVV
F0S7VqNnPpKK1CBeA5tIgUbmUsS6NXz2RsV55XlZOb0EJF2NA4VoJYeG3up/u5h5dK/4Gd+nFrBk
lGNUsJ7hIIX4JykhroOzb2JlZc56AjBRVHQiZ6tkk6GlSGkB+KARKDzuIL8f7NNzac7xVD3pACVH
1qTLPdVZ3aA6fTfJhvBaXpLDma+hioELk4G+I0gOvwCSMSC9Ooj31dRXGpGkhmECxjVzPKzGZUhi
aC24XGy58/rZOufjfNCvMRpUOD6E5oeF92EvmnlmcfOxMe4DulLyQGuSoDk6gsHT8IuSbBcWeHg7
UckxBrFGLIBPJYskUGuBHc71dx48wfQJuRkYDneiaAU73J8L/cAIDWajOX1vNPEz4tZksOIFobaC
UcqRzJfx/AHI/XfZdR8MNhl14w//9S7yK7dvWQsqxkuwQ84cfbGUKm9vtHuURxcVWiaZiExWkbCt
OG1rMoLhTPaS/LCpbYvisRmbCW8COdzIkkpcPD0ZTFKVDflV4qVRKObv3CymEc625UylJ6aU1uzS
Urcgu+W3kEDye/KgMuToHVk3pqB6WDJJb+g0jjxi277lGSqCDD4odyBraj9vXU7s6/cS+61UURDr
F/VvQiOLq/3CI5TAMK2B/x1d8aM88eyy3S7+eqC9S2UogTjTWtMnFFcfSWG6iBus1XbHMg6tGpsI
TNbBDLRqbss37xOrtRFv5soowoxS762Gme41rFTf8e5IOYMhRXTJX19ooll62qMdmMWF1qu2VhAg
Fu5XoKWNSaOO3QP1wLIiv0kqaEsnQBkUKsl8rOW70kCLch/5x9qJBShrRf04z6pAWG88Z7WnON8x
6/4iLiPAe9q2TLp8F1UtdPGJW0gzjY9/ocJafdvWk38r6Gr1xPIsLcRjzSo/p4oQ0KVel35IS53i
MpUMav6oqbddGem0pKOXLDJOAxUeV/9dRdh6sNmMNZvwCUZR8+YxXW5Kv3vXQqqiYw5Qe285mj6z
X6p9JrE8f/8jmR4YxPGaQFb+UZ3pDPO88C0PDdKYFjpBmwuE1fTzFULOPdxubYWWaKulgh4ycX6f
sBLZi2/W7qOe6aDkcgJ7Rf+JHemN+bJNd842pWCs2Tu18jfhoMUR+cqQbSa5zRG1GgO0YIqm5Zm/
dcgT66Xz3AecK27wc9hpvxVwnSnvQqAqZ5P2sYdg2NX3L0tpTR0BFHfSHazhN7n35m6OK4vx9uu1
4gzzx0P7of8eQOSJMFjhC1ezwjp+3K2v1iwx/3AfT8F5XLMkOEDJNQS2/Qj2nxe0CJ9TLYlJhFuS
DTKFkJgjkAjXWdeS84PjFWcotHFqjrp894mhCekUHkHtG9yJyGMVU+/9O+ZaDhgq0QFMEFS981cl
vyrbFsZO/5K1KdV18Kt/XKObRDAm+IjBPSRxPXj0wkOc5CWhd3owxgdRhUxcCQY+hmM80F5WEAiA
myMaXayKCAppVqe8Ui0FYt936wkpiJfVF+lzs0cdDKB5q38UYHJpjBi36/Yv28JT+mFS84CLdcL5
/T3WmYdS/FBP3QDExw1ldk++/ohy6nAcz4/z7poKyByj9nuPUGCcVdsWvCAJbwgMXKuTzm0n82wk
XL2mlCnCMxv3KGxKuDhJMd1JPhCxyBHa4JjN8ngM0PsNmWrrjZh4EeeXPFZx3jhN8nFyyH+982m9
aMI/MBiteYI6BzNKYNHB0p8tqO8hMbAVjAC1F0dk/ObZWoc5y+Il3Sqs5/V4rfxtjSY4EUyR/ydD
Pwo/0o/QjhWzRGIVdnjSdUYgK5quePoCjBPh8/WOYyhsqNxh3VDJ+Ze08pMRUGo/XmB1t6iF78q8
s6Tal+1omLoD2AhYEi0ruvYxYQdL3D9Qqg47nZKsAYF9cOdiSq6XPX6d5oP4ACYS+2QUTtP2bxFh
iFSnHLfKLIi8VMnJTCL+GZGHoOgvRZE5XvHeEJL11yA1vX6gIRGdOFHQLnBbdhY6FCR0n2svDySF
FlACmY4Fa1GVWbxWhriRUeV1jWBOLiV+GvpbiCn8OZ1/gMrlOy4KvG6ViseP4dPNGj5DkbQV5hSv
eISZuvKSmQMLBqS7/QFAcyNFWrgvZY0AZxgC2Q/N/+gHD4VvFDZTY/RVWZt/6ioNcnlDoIxLtBzI
qNJIuC1oxwN7ESiwgarJYyHfYYfdx5tVv45Ysjuwa5kov3KThaHa9xYrD9Qua6DfCsVxfHNNY9lo
aWy+DnVCcN0tribvlT9LjB/sJivEoH2BbY5dowUnipoBasBktLKOG2n1xwLQzFwcXMTSzTQUHm8D
7ZtPPkQjgJ5epY22EQxO2o6l383CpayPNNWh0KVhA9umi9bm2zNkyvfZ/mG5jgToV0/jYxUK4PZX
lloF7j/39rNZggBgqT12GQatRLcHkDTHSHs66xbYnMem1DsXH72uTo39znaLT+Njc2yxP+My8jXs
SsnWtcQEOY625MI7uEf7kmo2Ze4c/3OJdu9GAlnp1bKtwDJ0dlH3znARG9PJOMOQCaAp7mSHT4fk
Spo2AKVGqs7DZLiK92U7yPU7gsE3M6hwfI19MGJRTXhLLEPgCHqfhXwvVWxe4smSr/9hhCMuFMIv
IoVBlQapob9QMjAfRJREz6S2B/9FYe2st8kXH9s7BocUNwcEKdaVqyXAPWFKNk7eH7wgxjw6q0P4
7i1qYSobagKNbdQYYzn26600uk8sKnSb7FGdg4gHoR8C9MjFhso4QH9no4ZoiBiMKL40Axu7fKoF
wFRvzKx4+bwdNIbjq7e+D/Rp9ilShDErvFKW6YjMM0VLfvBaiCAqOhSgA0XqCLpU3xw9yi2Oem0/
MVNZDklfoDgPkqEAWL7IJHJFClwKo0Lrt1e4iLQQHMaMAbS/vYNQk50GVwXli6eQ3QbJk8amG98b
c4TYt86RRkbfILp2q3bE3x9I6RueFv1pqOl4e6e8o8cgQAY+UBQulERx/jww7jMVU6sD9TOGP/tX
XX1YOHwT+AxZ8sGty8nRmqMox4b1OOK5xu+OK6igPYfCnUWrCDEDcKdSDGsndi4NE3bXNv7YEuF+
7cWFrlo681JSUJKKOZ+BMWkgRwHzXjhPm1TF6WqVefhX2+yS8lNodT7Ie3rsEzAzVdys8sEDAJz/
BNvZ4rP+8DtO6vOWNRkXUwhGkZvlzvL0bCCQnhglusKyTmaihoCTx0rBGKv7OpuElUSvNAn+QJIw
YsrLkQk4rzBN4CnUICeqYfj9Au7+wgDrO2HJYo5LeyPTpxo3zk13zAh8rZir3KqOcFGeG7Ttri7r
YpvP5xZ3nNxkZOuqaGUfhqjmECXq0IFZMlEOL6Jx1KqMEKy2ShQ2u1+wxfZ6jM9Bm/AY4ApaWbZu
w1LQMQgnyhcftnctLIHJjPMoWD3T3pX5WnHZBQHTE0L1+M/OJm1LI9JPFe4pxrqaiY7uCxWayaoD
0jDO7k0KuLIoaI0FCDW2BkNX1hbEl8VCx3/aqts8ITMaCOaiaDzDYV+idqQ/wKTwZyNSJYwSBS1C
cSO4tVGM5AKyiegv+AvDvOvTLM20ns3NlFgny297uGXH41jUP9hoBk9dYREqNRXPF47VOi4bQr6P
WdT9wQEIfXil5fp1aoO+hXzXP6Vui7jiMgBZUgnm+0QrsTLaaAymxmcUeoCOVCLUgkhnUHYAivcr
x5+AKEosaO3onCRJH3CEUKcFsGhkxt7L6ZZrcjNz3/x8jLENxLY8bAJyDEVVzVhSZl/lC0JYYLYN
R1zDPkzwOHC/oz9+dhC/pJwvd5dtASB/NcYiuLabE2+He9lihCB81gqqEJTovGMoq1MoGdMz8Nq8
IjA9ERtJP0lF/c7cnXZJSQXzi/8Ktr2h/hcv4fB4BvXgughD3p69zcp4QLrbezDwYwwSXG1j/oR5
aj84O/nBNunSYW/J2el0e6ETX9bry7P5Klip0o+kjjIWkrLkKJTBcpkYHAKQgdOvbOagYK5EZjIT
aBbClqMKB1R+EoNnSHLW5iTJlvwiq00HUbKRK4K7NCxVZzbKHUrzP2VljXf3YLaR95n++e1PfxuI
/2J7WnVGjHQ742p6j3kuCMb93ghg7/LUgSlEIDerbEt2fU4zwDm/QqWMj359/A5/hOs0wm3YqYDL
+6hXfbq2eH07Ndd9z+xeY/rv//TA6zjsBn99f2qGlfVFFdvpjL1ao1aSuQO9cbvd3JLlm49atDNx
7EvamDt3Ij1JMMwMP5+nifGrIppxeYxPvN/DYkiPaqMwgJQsLKw5+d42otCEWttGJxN04JWHtrly
GTGsMk11yKijEnFUUzYIVmitPQkgCWkIfuzohOxe+qeUjGF/crw7oB3V7HrcXsFPkFcD0Xm0w4rq
t6Ge/7wG+3mEJXDDy6VRP9uYTGoZTsBve3LLnlGxwcsTg3ScSpcsoN9/FKToscXmPCew8xbKGriX
YYx8B5JppwoYjUA/4czwZjw8bGAJY5IKpZaZ0me0i2zDSl+EeQKBLO8SfThc+czd19QEHf7iUf2G
9kS3B58dQemgQrBGy5KFb5NVzn2q/QGcJiKikHNv8NjCqtdqP7B/S0sSMJcHkif4FRyHyTJvo+Sx
XQE/GdyQdT7vSR7cnFRNcZb1+mrlKRSD41rq6ueduSevmZb64HJX1XzYvH/FrpDiCWgCpPJP3ym5
sSc4knLc9oiKJ0GXhBHUo5952UahNSky0GgEEcKXyRgyn5eO1vUCXy3qonCOOKj3EWPmoeLqEbNK
znMpNCHOtFck/1QOEiWMitPhxmTQUrdWy+WdqgJ01K0PaeA1q7qY9VcUjGJV70rxn+SQibPJBm34
2erW5yWD7TJ2JvgeEbiMhDOWJqRVk6ZGH7ToGHlySGpkyoyzmb2roFqzeAda9pgEfhDiWaDXw8QK
J1c5JnftOn59pcof4g/b8Ac5/kR2BSwhwjKPavhNL6HDAR00IAV/iasmvMXHAjPUGAXOn2hDpOWa
uVi5YMEPyeJpDuiWbFEJoUroPphZhqoqjRXqYGIvsZWobyrmEHddE9TRoD3bpzuGYGNyLGDpgM5u
BULgb7x1vfBlE6qF8KsigiOXPYQiQsaU/DutXoWBGGOwrkYCE/z10RWIHGhkxY1/04rraiqVqX4N
ooFVjqKebonCmikpt5OnNjSEgya+CQuh3iVFTnAMwlZmPIVI8KqmEGKxt+Zy82q4532huTMoAhN7
N9t3LhI8GvdNqbULU74rHjsigtbMnZv6H2RI6BzFDQx/VoUS2CBrTW55AbMxTiLRnZA9Szl1GfMY
v41i4zKGNNDiG1miNAr1SwLl+7sED9i8Uz8Qy9e6kKDFrXxdU/Ivv4CqRjUYtb/h+B4Lp1HHCGWl
9bPBwkNI4l7tOsVK3JOSp9qjVmly8mq5HkMPMz5Cb4z/x8+J8GFqehlFdWiTZ3PSlefSfhuXa+2a
wi8x3VrjxzWWTwo5PWAmvdwfAcVMwZYTIM9c6aOKKZjMztkFFy4SWfK/h6pbJuL8cftdcID6aYX+
dtrumUlvmrt1nkdAZfdmQk/idkElHRdacuhyHzMDQl5gWQmT75PLM0qsM5pW3tYMnlP5dKNTFJOa
IYFnYxe7S+81R7bBlKb02qDFAmaF0uQliohDpkrI0kt9c0vCZhEuk1UxYWsa+zds/PSO8z/GRrga
649NPB4BtnQHL5yU7pwSA+vW28it0e2uuyntByMMPSUpQXsKv9haScQCBVPlOQTKWjHlMuJtYQ0D
jonHgE4kOdattwac1BqQSrtpvnXd+kgL7JnDlD6DP65NBbajNRxtf+LP/gooNb0r4Kaez1SwzC7+
RXIScU18BVWxCwZ8iFpSL+AKHNOpR3UyRpAukA4IM+sEQK+flFfVdsiPCXWgslbPO3RkvYx3Q4jf
2kx8H22BK7xlIMuMJEp1nIbFeYeiGbjfx/T+ax0j/jWSZM6BEgVAhUHJ2di4KbkoEhxqGBeWg6SL
fQkIADFQvnEoJnuO4CQVsTrWm69r/0Wl4RlPbIp5blRc5VtS3npxVbNEMRwKvd4b6Kza8o0TMJ21
5iBRoJVN9FmTrPI85gYFX8R4tf6O5k0iO73VrJSL4BsRRS33Tn2GGYdSFeLlzB36xHSZsMeK7ZmB
IFOS+Ow4qI2iNquAbY2/KdePE4Pz6Ava7YBMqcMfE0P1I4wNP5dcNfdw/7dlrbEfruUGHPYuGwPv
FbWFuSTSBFXColxTz6VbMPW2SLkK7b03Pom/IL7pkWjG4vco7425hZ1SfTobtAWb/mRXXC3di+v8
021x8WcOP6wkAjQu6Jg2LVsAayZYzyUWLblnA4qNWjSzWZqrEOqG4ZgWbNc5yLsQdsrK/TMi/2jp
gBOQCnjQMb7fB9kal8k5ASYSxvMiGoVe42fe6cBO1H/lfwttA7VeoZLvlZSGWkss8SJcRKPCNicO
ulWVmqHI7pV1/NnuR4KWjRZsX+jhkJ0lVYi78zxmytQc5tnTn+XaWVrYk2hv5EmuqZiCu/uFp/ek
RF7SW333FooucDCJR8rtjT0RWarSgqOgGd6zdivMW1FAE4B0tSzkrPXJYH26dcRoqjCibylvZc3y
/mGv5dIp10KjrHnfn0bYvCO2kYYK7NtIdNXuOwq9wt+wxRJPHGDTmw/zmWLH/xOKpB18s09xkU20
sKqNNY20Ocjm0r0DFZdGOwz8Wz8GcWj+BZVcbdYe25iOhF5R74pLEFCh9z/KXt/BfVQdAf1+6fya
j9Te1VyRKfkXthr5KmmqQlnUqgIxJMeI2qPmlv4FQAKT+m00dVzF0OHeBt/G9JpIfECsTeZehyrQ
tfFWdtlfLVtS3ehr+yqsCKnBotMYMJdjt0sqtNva5ByLyQtZgajhHpUFadl6MqCV2QsO0JaVgDJF
hA8am4EzU5PgtEWS0dtX6S1vuO1SAXlgOgGzbOO5B/JUgX5RSfbpwiuqLX1C0cCm2EEs03Xzi4ac
Dx8Nu3svDms21T2l0cZQNp4bJvCtBZx9ajb/JmT2iQgI0Gdyvsqi9C8rmvKrddJcbf5O2CxbkgQY
jzsRQFrlcDj7DJjqTbfpMjUJZoPNvhSVgZ8q44WmzQYfyUPOJeo6amTLusGN9Re2nThXhNIsH3nb
ZCD01KGvwmk+X4ZNDxFMhnsLiCQiWYqtKPOdKJ4sgBrr03XBkhLPgoe07CjUkAEV9NTGzJc6CmxA
VE4J5JZ7OTpwtH3TI/yVrh2iRuM1IqPHMmWa7a4I4CSedoU0y1+fdnSRcQeaNiQGKa3Pldkv8iEp
3fIVXbv6d5/KEbIl26sYn2ycw8gyUQDfr8ruNQMRUAtEFqBlu5qrudr1DmA7EhtPYLxlcORf2h/p
k2pWHD8qOL3XN5Z9gSFB8u1kF6+H4yFy4cLpik6pq0JI/iWVUfgPDkBuN6vWRQ7f8gSYsaC+t5EQ
AC4duxFmxSSCnwDxcnLFlsXGy6nvnR0e2A8QoO9iUIFV5uVm7LDUoDLgQTVwhBt09Z+eiwVH/rHY
NlTL50985tH7alkdtkzZ4huPk5L2AtMOR75D5ilExvMuduQHDNxh775BCGbwl4zkdt0EF3CF0As6
6SFVLjjl7t77vQKtP2urkQRvysOG+dFh8FukwHzhBPH4llr8busKy157p6UUzKQyWNn56PN/ccrU
fW0R5a/dPq8m5MIO9lRUffDI8qA7+RZZJ3QIMR/waKUlrWnijULGbbF6ICoB/eZ6uKYn+jYz8jBb
iDHFtX5MEHZMxpC1BNlbQAuI1MJO1gnQbybg2JsUQJygfnWhvoy7UP+HFC9WNOyhC0dAyF+SHW0T
Zucxqe7pIxcKDYarGxu0YZmc+/sM1fvF6+Njdn068Uvr9+iw0EUOPNYFORe5w9naWStsUSSWaY5A
Aln5X9INUGSFEsMcF2bbHsX5Bj/JsJW6mjOtuDZqI6a3KnE2gpok+iKUCNfAA+dss7IKBdpum8ZV
eBXz9MxhAuDscSJkVslGvP3Hv7MJqx52wyFQnRjyQIZOeYInHn7oVCJj3OoaK06EE2X2ZyJ8zAV8
zf43W6v9AH4LJpLWyRu1rG5m/QwKyTFqqIRwdtP/yeM90Eub61sITLR1ghDVECzkVzpHygv6WhsJ
afQYovpiTQqOZyiZ6mNT4y2V3fdqiLZJd2t14SgzGE2oN0dNaDA6Jl43UfI0VmaqdfWVPvmNaChr
VSrZ4a895Rpcppsp3SDawSfhfjiWhGxsqFl5r4eEnBFEoDe9+baOgnbj6FmdvsSxaCJPeBlhR1YB
M4S6y+6XF94GMQI9UZEykL2EonHmcdfmFAYwt5SjGo4w9bCqZTtXg5JzDsTZIV+qzzWiRmMDswGT
QSuYQaEJmKc6/7ZYXJ0ZntKde3+MpZz4YlvUk7Pyx+8HTGWh3QuSiU5OxtjNkEGwCuOIz0UFJp4/
adp24OTQVFxpIRKwBYSVdYZQKShir2FD1tqfxvrWnzNyGBf+SYlj5TYBiHh07OouOkXmlQSGXuuq
rWfqXbLo9h1L/nj8MoziSLyQkddnejt1h1HPvnNjo6FEuFYGHml5sChxZWCYdhd2oO7f6eFmz3Nl
9cDnG+fHThimNNswTQuZ+pSV54cou0yK67WpHzdX1f00JbgU446NIEwZOF5Q7TeHN+9CQOv7kMri
OA1l/oRHffdnElS8yTlgmuATM3YmNy+E78mssgrn45+eeXYrIU2eyunu2UpdNwHpFC0PVvPBhn9G
LAuqBsmt4p8JJ/WKDarMjFyKd1A+swF+q4m6H8kFKjPqGgwOAE3v0ZSC+foWbUa1yyZT9S0AHx+f
N5yVs1DpufZl3hhUH38hjlwgeUsZvQ25vikMxJXfOEznV8YSenypsuP00xsr6uON+tIqoBUkaot1
wYghKCmPKznolSutzUa14prRqNjj0WdbdZSolNCyty7zgUdIqE7tZDj2I9DP/QXHFhqmWhbkd1uS
9FugL5rbU0cdsoV3Y8RhJ2G2KW7ccdtUk4KhsVgI1jfHK4ukwPPWOtzFs3fhNOyO2JlTJY4QIKrR
P6RTBtGzsCjG4OUvDYcLNhsnaQMqoakUOumkq5i96H4Dn/qSgJZ21CmSeAg3oFUggMGcjljNDYTf
BouvhDWnTcvRvcMn6fB6zSxuic+hUJkcydoCyqwFUXtPgkhxvrWz5dLgF3qOCqZE8gPo3jOMK7j8
afMlc+n8zJ6vTYEVh0C3uEDPSoBd+hbnh67WUqhLCS3Fqk/b3a0qdB8RYBNzocxOCkfz/4tlVWZh
iJnzC3zD3KegjeOR8AADHo1oDpbD0qsnAkTZIaONC7UKIL/9RmTGbDvNLMY26+rV5VG2eR0SN5Fg
bGf2cyhtu9uy7VowU9DjBJ2HPjWmNH0DBd6ZhSTI3x2pMkrn0AmmmYJeR2XUOV/qKX/jlNhF/jhj
EQaimr5fm4kwbUpwmjofcoy1bPvYQ6zDWS5sfnijAJ9pM8Fju8KZmOthBpgvGWwGsT0vpr2lj+Zx
/3PzmB3GpHbf/Wc1hio+xYPY3JD3VIEBnorNqN0aJgLIG/IZld/VJWszteVidtw7wKZTGxcW8Z0I
retp/7lplcVtLkjfECVFmm1nvVcpePJXrkkW4rqn93Y+q1i6P1+h19zEo1f8Ziv6eFi+SREgKP8G
ioRUCKPVsHzr9YXgdaRTnfYlux/e9NRj8T/qUXQ1mtEaRB9GfvqdiQdiz+UFrgZejYoOma07/xd4
/GFC/NiVgtUWxzUjTcyeFYDCxN9mD6UNuWAA8E7BeheDYbTtuRnwKClTUr7UEc5LbyJfnpmAWNhW
cgz7JR9O6jm1xeZI0WWkhGtFYE2CYOCGCCkoUdr1jmgX0oyO9ESniBfBjLpJFKSokZXMHW+CfX8R
kNXjL3woBUHwAR2NIK/ZlmRis3/1paL8DbeauKoVUtrHO4NQd5vUJVCEqRAkDElxhecjiSGVZtJT
edB0nPC83fvM4zgvXPk7Fzc/0Mh2riRE8XIVO/tEg2l757UXy02ML3P0xKjF40+zHKT5WtE6pypv
0yaqoGLu2hcS/Hh9Y3yADth2YuIMC4uHNFAPlFGVmH5pnFdn8WQzLkFXWicqQNgHhfEHujVNUnfi
ZDL/HhyrJxC5nAeUVMq6CfofFtBKAy5OxaZdyiYG1ubPRPQKxn9A7xwsrUER52MZRWZ0w+eQCthw
1OB+wxqS/v8z2yjosFodM3VYoAPmyHHDjnYIb/1pwek+czB7vToldNfZEPaORDbJQDxQQzeBNY3D
zd9GHhMS7BLRFQrBMjxFtnXtjuyj3rXdOi5q0X9koFR2iDsUnkZQxXRySuIot3Wycf12DkAX8A7r
yigEvKvaD7uJ/aHG2jXCYSW/ys2Slry6j2DW1UFeYccL/ixcLZJTqV8Uw6edTyw+AT3+WVr0gMs4
6sIJ47gvmkk0JXbzLvPcSu074VoM3T3w3jamYxRQDmS9Wie0qrZx0Zv71bUoE+FVDIBlyO2fiZ5j
YsYHP3XNDCuybIuzFmJxJepIMJnqsOL6uQ2XKL2jBbsstTwz9nXl2sUGJaFLJ9qFbqe/wqcvlOt3
LEtfACBkQi3zw/xgNklFs394EE+ZPbD7cF4gaxjC0BaGYQydjONTJHYLNBX+9fGEGHj4WdbYf054
Wt0NUhvQgHGwxqMEIogFJ3P/hZJ7obhjG9E6jxS3iYAz2S7gnfEQUihIjMtQKO5lraeEzrM1ZaXB
fvDlaTulzlF3/ful8qNMIY9Aia8METF2Jym6EOovPA+Ulvd44pdOKX7/5rkOLuj5IYK+TZOi78X+
9tVfK7tPf2STRayIhQfNfn9Omb81SVopmiFBVb05QwliPSwFFVDWuE7r0HJbIEoTX9zi4oy/jnjo
7/wA2N96FiX8+kk7pT/LLTC5/lu5iU5R0HOjMRaqaOiYmEEIURG7YC877fDaNrj8xtpIWYye6USG
AWpYZaDjmGIxVGfU2isUkfBxtnC6+rTXb53SnwD9xtrZO3jPouC2HEMjNTUSVJUZZHYlU5nm5TFI
FiVMy6EbzToyvP7RAB2MhmHnxIYl9k7fvqcgli7gVz2LorxY6kbw5byGTX+oD0x3ftYm6eUa/xSr
330wv2r0btE9dAMVPh/vEyRly14TnJNckqfYc2It+DDlt4MQmGPkl6RS6lwI8pxdVsjWLfiOPuV4
VzdoaAHXqixT1x3pe96wZqqe2oPsTnfIvyB4ngN9T7CRK3f7ekWxPt4tu2oM8ocBtlBO1+wiDOvP
XmB5yhmOy8r0BgtuF92HArdvaSvoEa5rlmbMr/gNEuI5LxxshU8DjRCv0ZxQjNrYvUICyJKkGD7/
oRUv9MJBzCGkbGUpDUG0Rr4FhJtm+sLg6tX8GbZZwZcgkE9ccDwmpT3EU7UO0LUH+KcirZ/1BvIg
qLY7sgXa0w51DDjIPnRrqWbhpE/fKeDA0m0wj4ET84uRsUCbp+y6mQP5HIgCpz2QrSuOe3riU+Qw
iEzzmalmb7Ed83JerCiBJxd6V+v4/wQCy4gpZ85SKty4dkILtJtc/UXdiBIWRIkAZ5I5ILFGkPzV
8tvEtTX3XBqi38c/ijmCVSrOW2lArzMFTZLVpjCm+eDkZK5aqAdDC90P9lWAwenw5W+4vmZkDN3P
Pveq4BOeybQcmw5jt73cHtfd6LLpwf09yuGR7lpSBdz705oesOfnxS2nFd3Y9P8+XVK2bcZ8nKcS
zDihbxXXD6OQ0089tg0W04IVvr7oCubNpUy2ot5Rx+AUXxXfdoQHh8EeHi6TTkxAPl8RXQTxfVpY
nli0mPeyJKzfRVsM9GOgY8Py6PNw1hD0FbXs5aFXjQWd3lDuWGvnSAvfL73Ss0VIA7M/wLE5x8U1
HYDJgVoRxYFooeiJcljInxgYOzDH3Hmj1oryVFyTuTrmWNXoeSl7XThRWL52QvX27Evbxw/G6lMr
UQAnmvKbN9HD3LvjJo8nEyluiK36goNOUYkyBZ2nKc4Y/w43qAuV5iRQnib8FHJSZvEqojIg7q20
k6UC+TjOfZwufNhNvkL6jCZBnF7wZODEFdvEy4tETyZHFLbDn/+7oYhxHeIJQPWC/UBytx4pg0IK
7sKGlZpHcDTARavsYTRCwLXe0ykZmqZ8d3rNe8eGAenwYp+ksHxagMzNNk5a433kUrdfYqyu+RZw
18bS/BROxmN/ZQQUnsoPwiyudiGLXnMDAVj1ICKX3+zHFc7hI8VEwDlUZNcEljcG8ZwZd+jaO0eI
quW0cxx0hOg/kLY+foMySdSFm3U/5esDz6+BJQzZ3QFitaP5mxOVqtc9pQ1kEYwfW9T7cK5w61jh
nwUMQQ5IPluth33o4QSwkDC0m4ItFp2CNwKBIl1HRcDMaeXGELbIQfyaFKeyUeF/wxLdhgpThHRy
iWDU0XrnbOVa6ZPPdUrZ9aSuhtQ3IlErn5kbz2t6srenWR/lZ/kxopAAFisLHGEHJK69hUrVKHgy
dDROQ74kNLzpnfpiV1IYZkBnHlJW1vW9MGsDn7KSrFElof53mBEaCtTfe1JwEMxA0K1d5wwkxj2j
rzTlChxNy4r3UjqHWr9GWwmrsH5xgf4mYa+8ToT9ELkFsk9eWDT0XGIcZhIQ+nPxDVIhAVpAIv9e
2PZe6+eksGzfky7BR3CWxVH5azmKYKW7rBiWtm5BSDgIdyX7O9xqGIcx3zLopw9zzx84TUsMeZ6j
EsAH+HwiIpkpGZ9JMW1t8oohX3tPuON/+/12eMEl6PCyA6H9BhHedh/keJNYm+EiD9BEyU2uKL5N
08T2nIhaDoRNhO6tzUBtoHIe1Ltw+TgBRqvuVEhJ/cxVWhsGLiG9LXnDVf4f1V09WlER/Y/0ZrkX
5GKfaa8KnzD6oMzm/y/mOjLlcfbugHz3nuXViIGM+eYSvqFH/sj72A+9Li76OFIAHudg7VZH52EV
2qeI1BKb2LQXTs0hrlZoTd2hj/hgrBeJyBdhAeWl8Ljdte+jJGmE0BdH1aFhKNPNdpnSoCrSE4pQ
qhZ0OKnY8huYCn5F/AWGB0e0VCtcBtlDwHivduhb7Dm1rc9l3/QPFTI6GJStvs3rXH0uSjUT26UH
YRFH35FqMHe9KXCVcDQY8sOZLGgOhHPg21EHv0Zk4NcZ1nC4LoG7qc8pTg0bKVESYdjaELlItK2M
cTmWXi1VJcrYayq7rdsDnLfVL/lFwmZ5Y7HTXvKi63jvrZ+IZFKHCzzAtaT0QZWltzY7ddGd+If5
AKCqOCulM/TGZathjpEdzGE+BpVwkeKUaP/iJWyW5REUlUQkmzuj4yborSheht+PadpD7r3ZEp5m
50IfmN/mPJM97raZG47z3cvcYXesRDycf70/7+w0XzV/2P7j/KEQQxmyCEpX52wYguv8YZy3+3pg
SwSyaIMIKLlwZYLWc5UMcvQDQXm2VHt0XHDfu3xOxtIZLp+/Mo1w/FNMN4Mw06OM0YmOlpXEUrP8
cVZ6smqbQaYtyeXKnLQfk6ou6Uwg9BPKwtPKGJ+PF70lO4Whe+ALQJ3VMf/lRjEmq30cc9EdyyPr
9lIa3b239ydXwJW5GU/MubbPsSbC9S16OG6Eb5ou3asebfxkybq7hAnjBxfuYmzGjUjWJ40UB/iP
xcwjOyspK9q4FlCSYuH5OF4KlJJBJEmRWTNUeWKC02Cco65a/4ONsPMNfFOChGniOVQqxYUKj/jB
2Wl97ceHkLY8PTx3CbHee272VJhz4v4ssN5+GzzLINK3jLUw7U3lIfBIiJP5eyxRHGHd3y7gvnQK
Le3ydikISHBUYp7FBrU/UNSNKdfxH350EYcwD+8jTnZrjuOPy+mqkwqlb5dKKvWq+YiSJXjNe5SD
5Gc8tWBUgYOsXebNa1QPAMwVU4BwpFWUwhHRyzFk3jWZv+34WhvUTDTPIQ5g8zuCCjGpDKizCHBb
d2x+ZZi3Mp12vLOvharHmcRuUUj9Zf3xOxQxSkIl4DdgBf90EpQyu9b6bw175n7xjSYmuFnq6rbn
QzYzAv27R0LK3vImC11rEykiHKQIkEiLPYZ4QZoJ/lw8+oWHfibSPYSKsVS9WJsvkq35YtQLEpOo
oaHW6yprf9+/bcIDzCbHvQDsItDuL8hyRLwsDK/iV55tLCrnpV0RCKfZO1O/0cMh4DU7Zgn69093
vGUY/gfXQn0iufNrUvzx2d7QogX5n4sjCBDFVQaJ82v2uC+tKAALDPPrDwjwJJi2fd/wZsqUMJ0k
qjQfJnGCqwsAHyws49ICsp47p8VDCPcpCZWRQ8ORw+rWV9G76qz9bezX9fEy9OEM3JHnjfrCjU8w
WVvPR4RKIBQMv0DEJwui05Z8XuqWieVtgpRjit6m1xURjGvbbEkBMgz74nrQFwWaotWjETP81Lyu
HOkWSX6nh9Pl0eooJn8KNtUN8W8bMYn4nS9khL+VQCqeVjzpyE9nLZDWyJhqJrDgRGdbHSbwEstz
yiXKRkKWwmp0D6Em65KsccXu2RJgJaL1gT5w+9wFKXvqKYn2xM7zYdMZnglIA/DCnZOVLiKBoNis
rMa9XEaFLUnTGJ9pbJ5KRjNZg0ZwCrXxuR4a2d26w1RoCVRObbz3WY7g/EGfzWnST6S5GdiBuL9p
BmZ88e6BFA9g4Q30sZwp9uioqoIh6V6SptJmWZgvaFWQL19EcvjD7Rwsl7AZtulCtB971yeRV9lE
l5ZiBss0rAT6u+HbGs/jGyZGJjYo5DsZX3+QXajCLJXnXBWpih8KRSmoBb0QB/rRe7LVHnGRja5W
SqPEZozW+hIuUMy97mPEs1aEt4KmpA26Oej4Rj1UoIkjKIviV+vwEg+CzFavS1wjsNwqA0xthzNO
c+rnVmJHvSmD0W8nAgXmd95DQIqWK7oj6gaznl0Bpu8v2uv/0RNM/A+kx/L3f6V70fq038L6+hWM
39GzZsZt7EKEV5sgLQlP5gfugVDI1mLf/oLeMW1ej6mchJoZdi652k9mC9XDxf9v73Mbum53oJVZ
pADB0Dy02OxPtBuYd+wcjXrYB5FsL/nB1ivYLOhTOVZUXclKsHYeiI0mBKXrWK4sB0s/x19uWtrW
lTxVSo9gtL0jHAG6QciyUDFbsrEjtn3ebduL4K7z21vXcIaHDbXXwLfu0B/rztplVRB9R06Ks7+a
FEdkyBWioMkWNzKZJBFu415t1JSEcahCtgXFoeDL4XTW0LisbljpEHI4bgSzGLOHZ0KJIt9Ha0gf
TtF/blShxau7KRR3i1by9qvqwBAbFIx9xv9KVvqcFgj8Yw5gcCshg4o8QevjxKgY7BHhvoLrO6fZ
j3mw1jlqxZ488XgzJnf6tXHTP6Vj/T7rHiGc/LWEdfqpioCZw1LqIQ/CxLV6zR291+v+XAAOqrlP
6lyQIURssG9Q4qJ8cYxNOyQPwauVpppz51Jng/zrY/R37qIHcPiemdxPTtKvtesvTbf3B6MDTKHg
wZY0m8i3jE6M+vX3eVYcyWeXR4NRZCmGRnMWXHGoUb4Nz4uHeeq8lRUmqLuSaxum48uchjruCn6a
u42u/skUmAngIHvlw+kNryiEzjysM4HpaBtNFXZi7Cwg0kbqCWVt5MvU7tyGvyOklKzviO6HVfrh
pwHRm6Ofco+NDSN63IobSrUvdFQ+vTOqfMPejCss6Y/XiKKoNFsxiEPmWfVUcAYVyxhHW/njYlsG
vCW43U756hrEBS1MEFijicfQB3cAlKY/ow7a6MucCHyHdUWLDEoXfgnNvJB3ug1ZceJ2bXV0w3mY
pBSVy/bMHlVlW7XtMJMfN9YYhLjbOH2bprQNx75FkfQSbtv04meRpxHLJvEZIpyeNbJ9yt/3Jn8G
wKS3dp3DMzOFX1c+Ee/VvmBgpUuh2x779s13lBtWU4pN/ZjOqcqp0NvuRuHs0SzwoAwCPbCx6fb8
+P3HN4U51rneIONkAOn0oEd6k/yaeBl2qAbPE9yJi2DZ5WOq6HQG3Rs1gQSwo5nfMNSWUGQPkM9i
ssZel0UceRPtQKkhpbOpcSOAhNRfYvqClaLoE8TTmbSHV8o1qQT2FpzPQfSGHm380+vS4n+0SfW2
sRmGDZ9kYzx531DckCBzIhAbHH8VNquqiLWW2I4wd6UBpXEFgrl7FzmqcGQ0pQe2IVSR5gzjsxAY
Obv2arU/nz0T3L2tA1k5Ir119vbkZx4G30BRw+awqfKfonOPpTU7OUlWFjC3WKxzTANs2LFjHkgC
Ldd3TFgjA5nZVnhUBBLzR2wyNt8HwW95K95ogIu2veCKGil/s1Hdn1wFwRDokt6MTCwmBJ6gQK1W
Bdg2OJG+Fd4urZ9AvsbUPbG7tixcwzpfb3OAWlTUz6XnW55Jkp9ZOWzyx4nuKYONBv8lNB7obTUn
Q+/eWKd6RDij6Dhu/1QD80vPTnftbD5fdKol0sYK4dn+FnhjLYZpzj9OMjIu0CcPeD1THc9juL+U
Gy7a5Jj8ffzyr1jLfKzq7j72kpgZG0ftfAmsZSFkFE+EgUQhsR383IqEwU+Z5CGgHYFMn2ZqR/E5
gNknPjTnQgw5amg65nxW44P4nCorb5PXHxJT0IoDCG+6g44WcrcvQcu1iZ3Pt7P2583AwYlsu6j2
nXJWtH0TDPT4I1X+zmlHfhiOZRz3kvGCQUv3VQHlTCWQm2p4g0tAlNApPvk3WsOpY3TJhVR5BWUh
H/JTOgnwCQST899qKQ192bJWfXQIdE3qObaIiHwJe60ND022m5o8p0W5VgifdA4SqnHP1CwPWTtz
i+zDwJmwBR/btaWGWWcvEj0BfLTa0eAD7OYLZjeYsUQfQaS2/uGd/iYr5WaPT1vKIqCyyaAtz36N
LjnLZju+PTSDy8Uj7KGUuQ/082/KJYB1ob+XPb7DI3WWr7zJQc/T0m19sqx/vdy70fdOPXx+gWwE
N+oW/vRdv5ShENQBNyBPNdcLUu8EHON1meDpoYUfyhJP7iFBniQUoDrUouZj3/GDKb4vTiLKXmQk
VN9rbU82/GAE8+I1ZYtiQoToXlJlpJwqmI22SfJTOctM1Rb46u9P2Ui2gDPv0Q6wSkT8V0nC/qW8
4GNieI5F1f9XEPUQ8/kgBhyWSSgGE7aKeS5yznDM9cZ9o0gI+MGVKL26fCQb5ynGU+RBpIjrcl6I
t5qpJaxCj5PPdqSGwKhdnegCALH9jlwYr4z+kqDnkiwsWkomSQGPt828Pr+DMycSoWKFXUAhY0gG
M0SdcSUE+Mw+1BLaNK7WpJ3MKTvCi+jPugfIj5x+KgYonaADA+Vxy8d52WVURlDIyi7T3HRwIHTf
5laSpPl9kQCvZIdZzJJmqUshrDz2XPEKZMfgemxkcMO4M5pR10adA572NaPuaXJTyc0NqX/ivSDo
1Z/luJDfmhrkaCUTG8zCDNymhTw9anhcjDlmcuILCBTxXiJPTHWR2FYjojpUZ2xf7Y8I9ym6FzsA
LlfLOrWhXzVw+oeWoxJ3804gJebNQQokEIiiXfFQxXBCoWtXp/R+3YsPVwFixLmUbdjxNB6vd4Tt
ComeWezkloqHNLdltsYe9XVgsdHDwSMlWwgV0nWN3VYjyjvevbF3ojFQEIdvqAgf+DGNLfqXL6lL
JmGR2vIlPBUw0RUslHMB8wzdcpIReQXiZjg8Y/sNjIxjxXHA7jwy9t62FOa7uRTXdWtuBz0UPwJ0
WgTkP4x7Il7KSJviEipRSciZBk4jJNdXx5BIILtzFbieYszzkDfr6QFoowlgBxpkobBse+nLP9Fg
FLL2UOYrU4E75AKHbQRbLLn7CE2GDD2vLhGC+DMwRg2Q6AQ7bkDfm+VLr5sjY8DBLyObhTTmJCkk
VcRcholHskjN66ufKTbCLfYdHdh+TtkoZBxo1QDqK54/67Nd7lJ6tnbLHahXEil45FWJLIe9EDmj
WDziYyt2KMPi4yWI9OZ3iHGdAbadxz2Dh/s3Qk6TyADJirNRUa1yzqaGmXDsGuWiMgXJusUnRWLe
JWXcu/CqgFQH3v6n/koXSl0v23Q5cFhQHgrXx3K6gmUoN2H23sos7v4TinKhyGzI4zcgGOWTsS4+
QWLTqCawTBOP0q/cse6lz+GIbJyg4iSq4U85rPVqXKJFZLnFVK0qVysrrDfVhQujxKjFeP5C49YF
WziBmgnT766j6BZEC3PiYDZqEzkZ2NBpdpR2uf3gs9Wk4pmRTceP05+JfNv0UCkoi2IHy8YbfWM9
b2E19xJQ9GAYdgQhRf0z0FgVnUFpNzQgaDD7AYCIf1EKFacLrzDqmxk9yE+Vn8a8X6gPuQLUifOF
hPyASd/blsOgb4NiTzI937vv/sYi2v/CTFiEJh6yiq+n4OEjdaWPrq6ELM/3FnspXuihCJXMGI1T
u2xIbbJ8NW4F2gDLHcGVeWRANwBInaCvMWmIIA92MDFY1Stiwxsy1CmftgwN3h8sDROuh9TFHdBU
I1PJaDY8qqbKlf6BhOKeiKM/QukEcRuW/ISB3gXqZdIoS9i4I8NTQ0lMI2OUnOhV6etsfQ2MC+Hl
LsZLZ+6eThb7vxKsdnpZ4tukXpmAyCdb2gl+zYhUWYZXU8s4wJo+8wHMaD9hsJ9NsAn84m1VujiA
smH9Q7157z1zQyL4uWcLYETtLEzlBqdl3lEjmcJkFCRXjW7JktIi6tbuFJ51gXND7V+dq+xiDp4s
tDaHFJ1XPAw1UUop3+8ambxpaZ3ZBnDT1CenepenmgqC7eIDjmJmAh+IIlpGtQSMubTQARhCdspw
p7kSMm/zuA0Q3lsyMYv7ym7C6tyj/WUfaQbFtsd9PuRsF1wDW9JFuiR0djweOOxryvAVD3pzdOfv
qbwIP0p9Wxu46rWbu5xvVtj5NkqD8SGKl+qbCRJ2STzSAH4gsOre3BeCuR7Rn5c0FYfONhRd/JZ6
d5PE2ykWI/V8UhQNPnowfIgWAfaZgHHnLqmEqMs1OZGXRPmVDIwCzM1dwPWJyHKOzeyxsZ0P6OZh
xvVrXqQpjOIzIfcm1lMip9CW8kG1oLamX5h1qdvNs3z/YmiawGKD6N0nVhW7Yi3OnooIz431kVbB
/KF6HBDqfhE8aO5bQyVLpDOrIGho/O1pNdR/N4VzpRG09NGpqduATquTAP90lgIZ9JcyxNPksf1+
1IkNmrVjvpYOlCV9bMMAX+mYae48iQp18Pik7ez86qhnD4jedzC5tZ2yxnVWHCuU8EH04i8zO/wx
M+20/WCqxbCRY9olbqWAbRRHOUWxPtBUDFtcKhku7HYDciEWCqS5EqA3eEoozZiXmKmgjXnQ3LvN
aNxp2nEJB0KDbluEeHewOTCHcUYP+3ZbBbJxRVbTX7n6AAGzELSlvWfNmaZp4G2rsHOZPhNZun0F
HE2OFaGSbFkr8QqdQXGrz2dO7dIbbrl8wysBZw21kyetT7r73alNrBwFoA+LnLR8jHESLjXaqs7/
pCC9C0moJm6DxDbv7XJEtlZ1EXW0gaetra7sTo5joLWy9K8SOPDRWXQjixhkpcYLSMYNJBATwz7T
nJ2Y5ZNXAX+OsRQUmq+E99ErKNqYrgx7kj5p9GBD8/fJjYJcO6uwfdCceoKNHwV7eFOg9CwpNipL
QZONsU+uARINI/g615GZ8644wKPSQND66ty3Dopx0aNqLJf2ee7Eb9xGwUkNyAWlouASW5NLOyKF
uNKf5/yVdjSG6uRH3inoEs8JEsSTaI9mYWDGeLodbZyKYWiGkjuRottY9TLycGFRyWesWetRJ6/W
QpSV2euqEI1RMhvA3c6LgIrb1rPB7pZW1OVVklG7k/ZZSV8usBz3mdLqiD0cCYxDXiKrmzgCIsmp
k41rdjaFVyBWAZSu5njgd/1FtCbETCwNFF/7rFLwe4cXTimEoWubt2NxsephJGTw3A3wM/9qYzvT
0fUcxkquujENJKKvfC8tU/MMhKtWg5oHkpBOM/xfUdL8/XAJgJ5f6rVIw+KBU0IqXXcHIoMNqbaf
/qxOdSWP1I9ykkhq/b7ta86deQMvfC7s6Egy29OM77g62oPSEtvZnCxvthxKoIIVHJUaV0QoiM4F
WNvNwEyRsbqc0W7k5v+QRY6ME1pkk35k5QhxfxQNfKZUSNEZZCtmtLMB8uIvku1Ckn0a+2qu2E9F
TA6VcSAjlcTnssEUdWzRbk+x3UrvC92gU5YQmbUh1VX8OkF3d+6zirZcnMfTie/7yhVJ1o6FqLYA
ioEfUf6FjVq0LrfucplizZkdhvU0YaapM25M5+QqpM89M+f6R2Yh5tR7dqjjVia12kO/RTZ7bfg0
kOxco7EccYeCjY9imJJrDQYKdOS3ZldLYK7ANEZ5pDqsvq2hXHWUvoDs3uOMAYf2xAXklCq/BQcO
yLVEdDEHYv4jlmKKk/68Bz0/81or4/ySPDnK+ldlqgapa6Gue8+kc3u3qSgZKSV+1fAquYmPMF+B
8eqb7BdNZx45NSTBRDpFF9NMlQ5S3OIvkCB+J/9jy4FBeDxb6Tuxf2shSN+SYhklthxHjAiVBvdq
9ymFfLBtSePCYMcmd8SYLxXZg8yVNn17L+5BsR5x/7PARXIZ+o7CakFITUaOkkZlWBoP8Elbwtjr
mHCmqK7pcFwQBpdBI346rjhwEpZemISFU23deSqRZSfG7gI6kitmJi3NJok9oLnZQ6BQypdlIxSj
1I6Wz1IfWutIiItUSqB+Dr97mZeTdUVQ6RGRMrd3+B3ggkZJDkWR4BjLjiltde93E5KPdJM5t//S
cPl8PkAT44JS7LgddnlqANLIgci2FPLrasf1wagPV1EMltsMOiuv60CQwLo/XvtLCSWMiTFQuqwP
xvVy6FWHw0khO8rFZuRdjtQnU3+xpOuGoNbWJScZa2rfE8qgBwov0GAPfVZ4Ohkz34L4Rj+WQvWV
+1r2y08Fmvt+Q5OMynzxWPqKGUzW7FKP5I6hVcYpg9aFijpmZv9U3YPEUWnc8KCthFizmGhDS1DV
Ght7Gitoy6RPHWIJmES4u2gYuA0iyucUbN97XlemMA3lf+je8SGX7QKrbRR4CR0qs2xRHsw8D6yc
o0GzYcR6V42zaIzfiOjk81FRhkMFISD0cTEe0Nl/rzVxBY6/J0MI6cXVR9eeOEYwcCLktTxwtX81
wpDvALHE/0zFH3Mt+KGncRpa9tGZB5Ik5BVrLz8pzoO5kZfdMS32oPiBX5NZ5viLOP6nL4l0TxBG
2qyblADIHZjNuCNw811LBn+Ej1RjvRhymTAxVKbFlBCL33tS5uTgVh0CukXa2UR8YqFDfkxcUjES
ilM7Bq1OCXEvBMfvaZGi3vCkEajbyYdHUcjLCA2fHQerxM3ruAX7ep8G0mN8EHIdr66RS3EEc77w
14xMhviQ952WT225DodONLyIGHukPGnVeV08XuM3uy+yQi2P8uGw1zGyl2hqD0qi17WTsNB8fFPH
r6MhQMOfm/eppjErz3jig9ptAiCIwxwJFHEoKuF/iid7F3UwYljdCuI/U5371CtgzV/maR/u2IqK
gzsC5HR/Fy6IbTKOTJDEOmRkX8Ju/q6pJ/vTRrZ/gvAowVrkL9b0HRqYk3XlQLA/773d/N4xJOpy
cJKwtYSiaoi/eKrrqeCwhM+MYPJKGR54E21SSbUyX4hHwO2Kn+z9Y9ndHcMwSyMRxsCokyGfuQKd
/GSXHOru+M68p4quRGhsGEjdPaIpz0hw1bkdemctNzXWQAceL8OzKgi3eBdiOlBGadTbtywdG2Tb
iW3DCE0RyFVPUPPnjf0xGiTFMgdLvq0xlx/DdVzuHzZVYuPp/gpTaAoTbBpczmxJX4YVodoMQPdv
oOwoLhTri+NmCevCzq/924OCSDE2MfDP7C1fWwngdRQSq0z00kCCYxMI1ZDsRc+iQXdY22p4GsP5
wg9dxkjc7C+pokw9SuswwBe4AIRfErVSI5dAKke4YVMeT9xhqoL35VJPY5i4lRIxIU+0CvvQj1FW
uIbxbnkyj5tdsaH0gj/hz2CnlP6dkGMhmDUboxPykpEqaT2dAERd/YnOEDGcUK5XiAxlXd7NpWgm
rFqKvcDZgbVQRH7H2u29YRFBZVMVbRH8dsE989mXiwGG5CfwcDwl1OrxeSGQA2ScFmjMfyKE2I46
zkoPYbAfY/9Iv+gAo9uI8wdzkMpTQzKAQWfXJXrZXUBCpMYzeu6dgUX8cjhuuuNND4ruWxw7d0UG
jaXPxvS3Uw9LL2pE3Tu4jj1FHGEQgnAcoZpJ+fSRm0jYda/6UySe0h8PiYXMRTVzyem+ZLC2e55Y
L8vZGEVx9MmsAosqYTLYvJiRXoWfUCCykphfwu7vXiSIxPeRi/sGLq4Pm4GNgTPI4RpXu1+8d7vZ
8Ljc+IqTF79x9UZX1taEjd4UkKopgQJt8aWXWWZVl8o7f6S7Kt2AAstAshr3GKU9MF4MiJWhc9Eq
73VKnaQHrapTX7+6vn6NVj+E3++yCQtc8dKNOkGIoKMe9I37LhoRU4VE+TxmfqqnNVIB95TDf6Cn
9iuFqQkwijkYN58L/7r8XkAbGuYgf6W57RhBxIvBfk2Q0Jtn9h9GmucJ2OuyfZ1DzvSzwYmw3IKC
S+KxbuQUlxkz94YoXBLTtimGrDBZWSkBbTObUP/Oq1fLS6Aq/nJzUyRS8eKAivChC2t5jYkpjdq/
uihysfwjMJYIfINxs8KHArZ6CleI6JaTbausdeZGbK8NYikJemVTKkL0p01eTJlDKEUiZbDtiVQ9
I3u601j2dU+43VxC0eJaytH8yc33hBRgNTikXLfU4TEdOp7Y3radnsIgOcDFdlpDEOKozfAd+ZJe
YwxS/nxn00//l1TO4sa9dFN0cHt407z0ekpmtDQEHmag4Nqkdw743Z2NT4NR9oG4WMuCSkDCQgOK
uTb391gXY5fJywAoWS6Dgpe3Pk4iSiXn9Um5BO3npD6jW7idq3851B9ExmmtCNiG6j8rwaZDIYe7
lEwfJLcWvp7SsR+1sZUiN6Rf7eBVyfohGM4VdR9+VhorxIrS6QORCyiWdg2q5ucC4E2/RPCYlOj9
0U4V20KHlsWb6EntXUXAKhaFKo6XFw95xpi7sO4OZpKVL+C+uNz0KPab2zC1mvaY2g4atHlWsJuQ
NrAyVGV4KOlIyu/AvL0RjEt21GPm8yR/76WAyeXnH6E85QqhXqgQBKIB9O3vErZSavlwMUSp0a75
QD+6MRq1v5SpIc/We5tc+aYQ+VetVQnmpGX4wBI7f+SyBkO2NPyHp1YZtR+ZTGjLgxZHB/hSC4tp
SWAPQWwcZCGE9Ss6E6G0m2mhn4q3xqbndYV519z8KiismmUo3Dx0jfWtY/IKuu4ifHCqhdonKC6g
pm1TRlDoKgUQNmQgNRbiSJdoPhajD9fUBULr4bKychfYv47xyg8XW6vXQVMdRBp43TDlJX+P03yo
y9X5mAfTOLqaZQuXDfSqQ38RlmjszaLx/yD2AE9nwNYcKGewU/GlgM1k4qhBRRSRbtbHPur39LAp
pSDSov/GKQjbJLQbVoCIOccan7gAbrBH7LbkolfRUhQcdWMRQOSETdTAYHgytRAMdtg29yA8WrtJ
3dH/MC6HdqUem9+t/WZtlzcpO5LBmhTgFVjyP8YyckJNuvtloDKeeKAyzIIHcRjQtgI/UFR520zF
IpIwo3ZLf5CUOyGMuE1zFH6DeKGGZlkkYUzDgBzX5Nfmqnh0h8y/f6Bi+tJTvF9QSDkNOvg/pGrC
GPzBcFqnPe9N33wP/k95iw1XSnzlhPGzMFgJgti6Fs7VzWC3qiliSNWtqQYhXcRJyH0MqKIPWE5Z
avxIeSEyNOyB1lvD259N06ExzAVY+DKiPwu3OB+qqs15YaqhhXg3Ienral7JyzOxsLFaH1wVTDjJ
WlzagdUhClhxqycouQdYSRVrhsnplbCl1qB1I+cPcwOPLWw7O1/QA9FN9B8XsitfOQI3XDHu37Kh
ieSzfMPCxjjS3/yjlprbHFOIcAiEKpA1op6ekUUteElJ6eAavsO17orSw5xe0o58Ob5CEBJKc4yz
7WIDphTJBUfdlviKOCIwpBvesPoIII0G7PkNkPaRUgTOA7gd2lACVzhA8+T+cJ3VO32ec3TyjvPF
rxqmda43Rpa3xwVVI1DeM6SqBVljq+0QPxVz4Svbxizfzc6fRqORVBM83E2SVUExtAH+Y58UvGaL
GwONH9M+kI6biYPizqJkj/GG0eCa5ug1+9j6dJ5H9BP7v3xbZlgi8HRrFJhNWCHmpIJVwh9GFT9N
Pc0PJNH36k93dHW5IFuKX1WtaDw6KIYz5p6c0Mq82JVeMHvvG7Qq+xuT9CnbOO3K0rxdKfeOXQ8c
bFx15BYIPvuYwafm4+wEWd10PHB2slQN+dUV1UNQ44oX6M7OyQQNFcYHJt9t6ZTA8yvHTUVWaHwX
Q0h7HoQ/xptA/gBTdToxGznL962dTaTHuqarGwl7vTwQ3ieKOLGymqv0HUT4MjQIgaX8EfG/hp5s
SKyxB6yPNACCUWjNHaj4xRBQB0Qyg6Vf7TCwORMprozPtLpkWqMSHqVGOidN4i8o1TdQJkknkBt7
xHKS4vtjvh12sD29QQkFemoTKMeh7mWxgXnUJs6fFSbzyZCwbffC/IFzhEhLFRhSK6hfzjVtDtUw
N5rn7mea+ZJeh+dBlmwvpOdp+g2IoUPyYqEqlCfhpuNENNSBsEolTNFDI5Ybhxor8spUlI9tU0Mf
d6Q8HFt3Sq5qXddxm7Dpa9dXX9BoNGHGDUYzaugvKmAH/tiB2vy8UabI/LZULLWANoijC2T5UQwI
qWVy0//vKT7h9n44IoGysjzEUTr8iJCuloKYDKs1/61PDv8z2o6dhDIG1V8CZJnnf0NCp688qSrn
pmJMD0dNsVVXbMLADUTbJKZ8RSHDTXItShuNMSkdmXriavfLyrxRQTspWRsTFIvLKDD4msUBubEQ
ktlaa/w3oqzXwdQROqW3AZMOQ2KCxRC17vpgRjOM2bzj1HpUv/04usoEqcfi8276FkIj+dCuE3P1
TrdvhtEsG6MgZQuEniYE11giakuF6X7YwKPszm3GTLwVFgRjOJTnPKS0ILadlC0PGlQ0Vh7WMyE3
J4i2Cj30/huwz4sgF+38CDRrMEHFVDrcObiuIDPtQR763pCYF7NEpwUz0LXCZD1SP0oTvnvQBDfN
tNHGCsaGosbH8O1N9NGzSE3vTNXq0xH7QQrjbDaCekOu+m3fNEOO/6YhFaoUBPT25vwmXCq3PoWN
qVgPUsFtwIANXXgdBVRQTA2k1PSnu836NoRgRh52F7RHQoseEX/62tZcAQrxFoQo4v8Ag6Kpdduf
NFnlgFJuahF07CV0K0ncYG6Td/i7CIZ8QZzhHkxjYPwm4RzJiaTb1bVCT0Cebd63H848jcR5x4vy
41FbMLCy4B3oRn35vJiYG+rNLCixWl+F0HfnA4e335LZRRbAajGpjq2GjfPus2UTCSxnUjHrUNVr
N/loRHSFY2YaYum9EiI/AAHAuGD4Rx0z0kihxv1hzZlLlauP1Eo2duHi/0r+G/e5bkHckFhU9VNg
7i9WeqIu4UZl0OncrB6O/HBz8sTYQSA6zRYIykKitjo1qKIfr/fbt9phHSxwDwUaj4XRpVrq8CGI
zVqVgTqePxdNS53l7w7S+MOPnBnnHRw2LuyLk6G7nFj3h8eTsl8mX+Yes7Pgn4rgejENUlSlHm1J
XRyCHzliR8SaKSHbbeIFtSnoinfAY0Yr2rXgAO9VKUltDcA7QTqVH3Y0pvPTv6EYAD5kFdU17aXy
VjqWJ7c99f2O1TQqoE5vLMFqJTgLNHIUSl3OgaY1u/VzzaCtoNqAffXDE6OFspotaG/OA6LRNNAR
mE8AVK5hAe+RZ5Wg/aP1MyrAzceFp2ejpDzLiOYseCN3bdCENo2Eas5gqgHPIvHweIiybCuRuRKF
AdroQgVl8UoUmssjQUT3oxL+hnA3cULP9AUCxOh9i3waucW1pGiJmbM4q20/k/B/hxrYOjZN77BO
mdsaV8GLOP8B6gVqfLjGSaYF+I2iwjnrtujdX+3Nx1/N//W+VCo2Iuevi7ecJbMT8E4bJViUzowq
oB3BeoPg4pxQRADb7e/vRh1fcVflAbtiN4pwb0cXNZ3u9rwg8OhXBIZ8kJWrK3rNOc4r4OJKs9Zk
YxxZsaEbmNBsQ+MhxtIlHFd5vTUdqB/jma7PbLppVMZyavcQAkLnSgs5oIEAl+D5TR1euh+WQF1m
AbxLN0DMMmr5Ot7Es4VjM9mCV21JxVD5OmnCh7ngyZed5sPaApz/SBaBTtXoSeQtacYBv7rTrUhr
YWWRL+/hxFP/UbpT75gk8OJ+jfK+LzeSmG27ebuVg3snw3S15Yq2tP4lg74oYAA238ATfsak9HK9
da8sJGtEiYZZuGoWaa2UOojRLl6XBebmo4jMAVulDvCxqv+RGumjspmFGGY8J21SgGhgnt4K+GPc
uHHUqkETHwtW7il3DPg7VnPJ5rICAst+SLzeiKRUkv5eOZQnJuPTiDVAB8OTGWrMTr7wsdHVpsIE
rjpa4wu5DwUnBhxfFvA0xPza2Y1wIYgGVEPo2U6cf3zgx7Tu9o7Egq43evcadzd9f7yY8WUcZUdk
Nofxt9tYEN53GJCU+4J/PfGEaPu2bOTyc4qnfd8N8cZfcThxcOen+Vrb2Nhs9L4ZG44VP5PrTBow
1rlf+HrouaU05QcsdRRqq/4SGFSU/pTBAJaM+JYJQj0QsigqIsw33PotL/o+wikie7vEAijsuJNz
P4KPMDdMyx0RlEZ9KOdUZTZMIQZzmf5zDPXmJNlQyDdU8iUJL122YDfrGZU1IVw8FeQah8SkfcBE
AfhgfKSU7YQD9TfQdhJ+hmU0eHnmCLdW1MCoMByfz5LGx9Hsk62cj2vTVuRz+VkCE4FmWvtGmunY
6sdOs7JMrIVLHMeMWwHaAX30V25i2Ai89bgVV5HLi3IzTV7Qh7ONTfa8aGRxEtLgJKjaZbcZ8+l4
8QiSh2TMeT5SxWAsaoA6OWJMx132vVYljHOrHz+z3uu0AgEsn9QAYxagzWBXntD7dlDAo9MY1k6l
RzVOx5mG+Mzd+AxKVjRoTE0H7j19j+HJgcrN1HAQP4s0BqNVWWwYyflf3pp5Qaum5R1lNmhHerHY
QBqhOYo3kpq2BWBxRxAHbtimGUM9nd+WIi3QNMzAdPU7iF02ZWyawv6KlksZyrQCpYlQ5R8G/QIt
Ef3lH3StFDB1C+/BpKCH5xuzKyzCScniEtdedZK8DE+jcJmy+UDNLTt8qCqUNnT5QF3xuMqkWq+i
IAh2N1ViIwH7RYKb3QK54cRq123nZKZwXElnBjP2FWP441yORGZG+NNMkNFfVUpenH9krsnkhBpj
vvRGpWTGR0bWVrLoKE/aKIzcMiYhgs7eA1WxT5bJQq/BB/mbZd6ellKmbqqH54nTwYmQwFpSPlqt
xwKrAaiqMobW+Gku6JtDQWnY2qtbIq6mh1LYrzcgcdOplmW70FZ0nbmrNmqNL3VmTo6wTxxXo/01
d6MUeRE36/LVdkgIUh+Mqb9IhaTYo7T4nyjGUwSDbNxu3SrKAixROoA6MDrA0aeGktDfISFvVHBR
tsMPKIgML3XRa2iM87cTq94zpUwp2SesPngE3Qxi+koi2cJE8kvgmGPPI3sl139uLriemeE3X+r9
WB6y15a8wA4DWTAQa0mdinzPysFKzKsDUSxJ2oGUNDqJ7N4qnP93P11m7Pak7lmzSxkXBK0MjfMh
nRA2P0je7UlHSJf3IDJHdRpBqeCknRe/hYY2UfdZxOzl/QDFsbcO/KjBdtNfVc/vqc2OdZ2i4FvM
tZMnxO4DLTuB2i4ZLhvsAX0pfJEz5EjXcHAlASUFxV14wWNwC195ZMPgXps52nb9dSHxlv3U1DOJ
XNQEk9crQItG31oRd9gi6UnloO5jbN114cG97LPjNJRSs98T2/htRqgxU2KbR2sKSctQTKmhejrG
OCfs2KPvRe68v3B9sXijxgoTSJiruf0Q3xxfTXoEZn05/aKk3ZbRx1uJ+bj61lK5UgbgFxPftm9C
CUcd9yTAV5NR/PtHo3VFUjaOYvXHTixyD4lwtkgkNnWjdMjcwHuqTc6EqjODKdXPOd6NjhTd7ezH
F4eGOt/LGJ/rEA7piwExrnEhZj8PruXPQM0iOeGrsDxIAj2O4q5EHUfVQtFZ+1bfaa/bEh7uaje4
dSVXLn8urrXpoNbVcu8tnenp+yibU4nDTOPVGi0Iix3ORxOUkb0lLa7Fjxg6jwPX0eHdWTpuKm0g
OmlN5UKRiuMe91SZg1zWGz4slg/kfj9drpCQrs7sWITho6DFJo3TaH940IPGEwihfzMkNIxltLC8
ymqXfikJFsmGRJ9i38XfKohGGUASdxrz/MaOY8bDDdHy5++fEfVb0hAb+5nk+Yx7xHRP61pE3rod
BlLKw5fLNKrVaKqVCg3+zGRxPVsBV9iOR83VHr2Co2n7eNAuwIQU+YektMUfNXW9RunUaw9UjNSD
b9q8q4XpiQyUTQ/SYseEEK1DhUlLck/Cpg57mrtbh63A0gtigfmI5k1NWRv2pS6pKP2wdRxFIH/6
ZyjdATSVWl8sVVv+rkiPyoZ7t1WtAqkf7E1zXR6yy35Qp9WftFXvpTypULzjhD6ugLU11gg9PQrN
G+5y3F2D4ZNnynHQNuheo7SF/3EVB9qPxRFyAB5bdnZ63sd9XWJOXNXR0/pRp+DMBM8QjrN/0sTV
RxLoxc0Ov4CP/IX9EZUyoQW0i6Le5/DadcCgXuySCUgSK7HXI+hMk4ZXvnyke4D95pC2DX5PRTXI
prKiIFsKkzaXL/+srkDsucjwwj6BLa33svjAr5CmYNZKa28BLFM/25MSbGK0mi4wYY0XHSUcaPx8
SUFljmO7K/Ul4rrZw9yWD0gnqxt+3P4pd3S+ES3LyD9hlhUcIUnnMnptflJpvgMj5LsCCP9B13FX
IN5ei0y4DH6ADjhm2wfgoMgX8JlCtEVshVCfOjWxREX8/90I7Juz62jK5ilvXkMflTKuAfCMzIDN
KB0yjxrkOd2sJhaCtjMvGVGQiENjVyuCPfsaeIMME7Gk5LNbPNY9f2R7i6FTBXBl03/H7mU31B80
J/5oVcT1qh0h25c4IoiUMoydU0apPGTBLUI2yF3VjkkDrPz0lqsZutDF2z0D2mMfhalEKyNeNhto
t8ghtXD3vXlPyMPXiDni/lEm64Eh9vje5MQh2rCfcVXbqPEX8dE9ODf2n+5dLWIBwUz84aDfcH/r
qFxNA0C5E4A5YDJyDQxJJj7yCj8cfm7j70MLpeUG5Q/8eYYaFuUMrdBNeIRj7k8jMnM5nCRrc9r2
0IDWg95f1WzCwKrp6D6yuvlRHrccFlxpo+uap4jqkvCwDXchDi81r/RrrNIo9aUM1dWDxXc26nc9
deLzhjrWuUbQS5QVwJNvRHWe3bpJx+314kC4zzm9FlMEV5gRdiTYJXacYiVWkIdeLcPJUU3Vczn4
vMW6x8DGyFoHMaR8ASkoO4uMpepauFXU4b7Ds1/rbdmMT997niRszJWGMlZlvIqI4ZOANWGDTf2T
1RhF2zZa6iZXpi8/xhsvFTwtr4gt2EJ0A7MCqiALtIuMKnBd51V6Nvcz+cg6626Ivq3TweqkEwhB
0WL1co4FYPJuLsh2FlzGsoZm2xIg0cnyqJB2UPHFmcT+x5Tm9iGHUCikekXEdHLAIGFqCGoUMMzL
uNMi1pfph9TOteyc6oYMmYGKUebBC9ROa8eWxX+3TcMivIzbTakeuacT1xkltCEg6Ox9gItMSQF4
IKtrvW/0H3RRyGazdQaWbUuuugVrLG2gZfdk+vrgLlUsFi3KQsbc5tN0qsYGTsjaazX/DqXTWl3+
9liz1GX7LU5KwglCOHuF0gP7GqZ+nqr83yH0XhTF55qGssmLtKacvQneQW5ZEQy9l+3YC17M95aO
qAxt7Y5VfL2knFteDJWLKnv5oo8DjQW19ZnJs3k0V4c+Z5i2oLfX5rbOH33cEGJ+bz7PWbitH/hj
On3VU05LINRGADCR33w5NSIBcV7ezKDgGUClVb29N+ke+U78uUce3CNusnKQROYpLCzfnyZfnF6f
QMVOrEpTocKbuW13TdpFIqOaBjcCZ15fT8HKAwCxPBHEcdauHgO1MdfpwRI9oMdy/EnMcfOsoTgx
c9ggrg9t1rS5VxNzY6JmyuujFzcrrXI3o38v1X9R5lnyrFUX1tpL+i7yBrCzLXc6Ksbl3QaLUCaf
PCoegMKxEF4I6eemxE2I+ASv+V16Q0kwLoWsT8ecpvxcQrmGa9Ez+yfiIWkThxWQi6X5H18WUCdy
YKHs6TlFK9HG+O/+pBNgIKzUvHYWwD9SDMCtrAf2F26bFtHj/iYSIqH2pNPLROpP46vpY3i7qjCY
bXv3mEGl8a/TOzSYm6jft4Rn+17Ob0UR3zRazo4j/8MJ7X73OoYve0t7vyoaTnE7kudhTP+enoFm
nUQs5Jpdjf0hC5ahP+RdgjLh60O80NYmal3dMH0ABIrzIjIWBRqAzn+rLAanIW7cZlInf4f3VONk
Mru0O0eMNaxuC91+vTtvHFSH6SkaQfICrAtjooDiIq4las34Ql1TUiSVYP9NyuL20+NlFm2AnWTW
qtclYlDiLN/wIdr28CMMWEMaHDLYmrMzRNJRL6qXy/bRXC98a8GDmNTprilJAxh1/d4rJvQiOnoM
GEwdtHJ8H2Yszlo8UjSoVrXN3ahWKS6Hi5Hm8k/3p9ljdN0UsTaDD92AbSp8/pL2QnotI55psFdx
Mfuvu1q0WSCSyvUZNvruNCNMx8q1F1JTrDl8W+207bXD1bWNVTHCVi93Ql8lQkJaAzoreIXSwTRf
2RdfyZbHAlSJ6apd+18n1wBgJ4t0baQP7ryR31JL4FoJocmFpHmy4vcifulayPBz9zGYl0CBcaas
yw4LvrcytUFGSE8n2ExXV0OnTZdsL6pRXoEnUQnsbnpue6TSpq9IEiLGbSHuyKtyxpf/1Zc8azk+
kgpsJEGnuhs2ZWL55YgndapQeAm+bp9XereA7hHz8MoB3EDiwlVefJKWKfvfxJ3Mn2Fm6DmEdzez
RRMLepzVNugMMTrK2T6AL3INTe5ui57WzRyASXgsjfxj+Uwg/qGd3gqJzgZGiOtk3xJKqNqUl1js
RXhW5w44nGLv/vQujMRBN011CVJusMY7z3Afh9/SFk4Hj7180LXJwXfMBUAqn4iX+RXwby727Yty
RfAmtZ5pYVXAq3V2/27xjWXKOQ0MG9zescXHrYCK2B6I6tSTfe3sQ+1FQDM7DfBnnHCNTDFzYHzg
hQvbK3HfXrwEy7h2H7dIsGUjr9M/OeDPgAW+F2/yeeMZp5OEbb6usuhiuHxR7nfR2wb8TWUMyArR
du+8li4LFzazdtAjOfSnOIGm3MRP9UtdF+a/p+B8Vd6q1TRK2iNzPTxcwH34vv6c7keG1XT+acb0
1XBQBVZY0tcPk17ft/kkf1XR497rxYqTkD0bSmruWY4RxXyV58t1y/ZT2HWj6KaC8pqJSpTVyk3N
NEmGy7o9jHU29JGCAR7RPj5lV7tK3gMLXTUhvNXEPMzawot61JZYTdxjY077sqyqMnmDaI9AHer3
eSmHXbOZCxsD3eEgJcdJenJoNyTf+3EFslToc39FJ8p9kKn4K9FClvbt3zceZpXcRWJo6raEzMkY
wLyUCkTT1wH12kMJcVFsntIziJUOgSDCp76q+sN5RFLcz7HxRFimfIrSgVn3o21wvu8+KoNGr0w4
CsODzCoTN5lC1SR0QmBLqly8rK6CaVf/+bmyy0uzYarRe4Bp/SRedD2idY5fh5+ESe0GxR49ppDW
RiorgUnjOjLXNm5mRmh1oIkFcAkSDk8l4qvDntTpGx+KsXIbLJpf1C8k0GD6ueNh8YfgBeAkggAH
EgK+FQd3BnVbJWSnjvILLoduR1U+vEdlc95AoiE5pm8VXEgGTrE5wbpjBGfdSXJHeB3AQ1eCLJEo
uEmCZkmfv6vF9LaR6+mE0JGrdoKhEMU+FBpEsepu33xBdH4uMBYRvApMmTQaUFfAQGuUNlWC9dPK
C3ki7DQZAHqPwdiZz05OvftoM/OPGA1fTcbfXY5QHEyB7+81fB8EFv2KgZu6s4u7hlElre9KSNSF
gOAh3exokPlt67P6Lb95mefYE2YNa/3SY86Il6QeaL5qMkuqDBT9sBTZXibCUQvF5zU67/Uoe8ds
7uOAqPcMnEaHtIHH2Bsbw2RRbEsG9oLNwWi486D6do/T73b9mFRXqcGWr/S89ms7smfAfzwIaFTt
nRnH4XJGLjkf/PB1B1MhYkgyrPuRM++oNMmH6IrTATfo1qIcGbmrUdGMElR3/CehJMFOHf7hNiaA
9xadDKY7uoB5+fxEdZrfDW3e4Y4Cd7S3NQ6HSWll9HZkF7JYbxqIglL1gpII9AVcgvjIXVDtAByG
XgPBTTADSV6sot5RU2sc5YA9NIFTiKfQVi3BLkQJzdPWcU1GBQWEPH2cU4Hx6mL2UUZeL/3Vt4ER
MYDv0JR7uPEhI4omocaQH0liBV7R+RU0derJOch/jnrx4WDug2m6SkoZMUQaw21YiFf9wgekliPv
fJJQU8zR84M6Q8x4rh/GMlyaHVM0vrCwy5nfgQKBl+vsTontPXzVHr5mafk0b5JMO42xG99dtKzc
K0QCRHafKkyi4iUZxbEy3ylzn+5WiNTzdmgOZjgL339N1S8x5lpmYsLf0a0i56Ul/qadDuI7912i
LZ4+ZS5X5MycN/18bIQzMUWkCsVn3O4R/Iq4WoX3mSVfHN1jiUral8FuQX9+T7udA08s5od/Ybo8
PCWzm9xEDl91ipgauimp22M3QAryLuGTzQAYEBMSZzvPTnKtqra5AZslhANhQmvdwaxljQSd3G5y
uJiXPqd+SS/qLPtWnYP4knx5GjzCk/LfBuEfAZZAX0c+3UW3F5UMiUuU+KoL+5uNb7QKdEHmGPU/
5IBokjB0JUmgJJQ1fyV0li3YuOt8gIAkKLJPSzeQDrFPz7hKwjRZjmSymFjLG/W+I3veBwQW7QdZ
8REUKJrI8cUOdg1AoqJqX4k8Fw9g3PaNZtV5bGaV27Pguc636JaVLjMyXqMFU9m3tLZALpJ2L3fn
3hvBMmkVtIyrRwVc4bGgLNBHGOGilrVsGDsLcq+QJOLZXlGWyh9orbrWeNlWv+gP8qH0VvrfSZKp
ia7sSq7ABMp0/QNNqF3ecbjAWntro+gAk8uF0uStPa5hcY98Ov8+xD//NiX60W2x6yax9PDc0DEm
D6rPHODd7UpcEHqSvoWeqSvpW8SSOvO5+uxakwKkFKgIITDvKETasNDHUj8T+XI1LQ0v5/rrTsvb
5CZMam19zpUcbzTqbm8fnr17HYOtm8wj9zSoUu8PJKsGdVX9tRy71h4Dv9ZFmruk2mj5utVotcWX
ZtQTy0xHMWnV32DUp25tObwiy4XxG7sUAM3Yug94BPkgizysqbNbHpkhdLfNMaucN6JbjRcmOAj9
jozSWvP//qroOknCJpzbJPQB4CdB2TSePFePnGw3+2dlS1U62fWPvZbPEG0LDBBvG9Nr/X/73Rjc
HNEBD4o1O+4xv2b0Fy1CFO28f1XkldZvzmkSWszMYguQKZD0zd/AQHSNU6pOZwTml6kL2rdOmJMg
YWgMNq82mrq4mk57aChA9dWgMHaxCwjShqnX/zSvOHfhQVtvMqCgW7TLEzw3vZwQJbmyRuOpgMX7
Y9hnjN9tQi81hI5zaar0kON4jYi9ox+24dDTLdHXcJTer00gCZCvs5mCEDG5aatisAY3bCet881Y
d7XCR3C4cZGJnrd4icdOZCF0oixQHKrclcBw0KoKfLuXhjfB+0xtSngitYTvZrK7PtbbxjWn/rci
HjUa/06OGy5A93kTBPP1z/PwRAadMJbL6WccULj7pAqb2eVtzzEMFctVdDTk4BCMd+bNnjmnqCpr
Cj0CrVED6GsuOEhLjgPveeMvnyUf9w1TShZECVLYXqNGqHlkpUnpaYprSM1xHuDjHd4/Y+mCzion
lTPqzb0sVmozl/0p46IMosZvivBPuB3OiuVXPdsHR2Qc6ZIOQFhgTMVPXosqMmvuNt5U+PcunFSf
mccXk0RLy2xdPeOfCqcUaH9CzCQgBJzc2QpuTobOqQ2njjq1jQbGjk354mcFpEjHjFCIP7TEAH/y
SqW5/XrRKCG+UGlrPUKuTxlLpVQOvhYxNO5eslIp6uqtynikW6IYbO/lgavwjp23jiUW49KDCRF8
EEl+k2Z2QyXFXvh9LEE5OI7r4yDVf3I8WhAEDCxCHFhvpqyGP9CLbRwmBXDzaTU0YqDPuOS2FM0S
cJN8Blf74SL54wqv75GT+nrthWoo6rcUIWIS0a+JT4QaUvsMEEVW296pde4KtLSjbkKxd8O++u8A
YF41ehE0/5ZkKowd5L2tIqmXxTsu64MNpxR1ygA7RbxtrrW1h13+pGk68G+cGWDVu0jz2hEZeW3i
cSf4BAdizMWOIYlmQlxEHb+X4ZGHtIXpCF0yg0LYVbEjMlBsJHKpI14MQKmDHb6CMJai+8AsHHmM
ndVabVQEHZZ85vVpX6P+mME0TjUxfk3ambKF+S0qYdJhlOD9cpmi950C15so0sMgvq/JSqyRGTRL
rC4Ph5bo0ey7DWaFoh8csvsH6oV4C2R+3wHc6xmE6n+A1jMry4g2eg5YKKHB5fuBPMh1jkrA6og7
5aZJd8nVnBMWXF/TqurFle4zvMDYKAVkCMjtcbGc3kWRi6vgegM5lJYfMrqSYnRHAeJY0kPT7IG8
BKP7fsn7K+gGedlnHk2v6APiFsi2nKOYWE2PTT05JjzyKZHDizZpaUmIvgSeI2tTOLFULIculf6v
H2oWA+wAxSlVR85w917RfXS6hVkR8ax6bLwyM4+gdwXzcz6UUHKMIvg+cXrpd4TEtm82CapXFnqv
+NZS6qYkkJQCQbuDgO0NADV6AvsI+raRtI0wcLxNXN7LzLzeqfHbuJaUYDp9G73d1s1XyfJQJysX
6QlqibBiHvekmtWeYRGssc+TI/k045S17uakFR4rCMg9LK0nZ3lLepjjjeAEm1YlSYd3e+738fci
5ZRDsw/fX0HpIaHn+eD1r5zPBosEBrl2VQXICs5OoQzaB+XSy54dbexsI2YggDYTDMEkc2ASiqUX
wgL0RDpBhLLqw2KeQdWCH/2HZG0wIkl92Yq40mguFxDHKzfHXk80LgyWbgmoXDbHJppmzboE0TeC
6tu0+qymyZLVb7Re+7uOAOrXq/441OS1kNZyi6Qh+gyZrM/91iLyBd1O6yPSrpz8jG7vgUaTG20e
nF/pmAptzcjAnJremAv7zvMf/42SPMGSqxYiqa8u5E23jhyrFnZuwj4PHbCyb/E1LJk8bFHdV4rk
Q13xnTrukJkmnF/q7v9MhAxXeo/w1sHmR4/1ek3M4yDUMG+mFzF6kNAX5+1vxaCjcQNP5N+Pfbpm
CJ/K4yxlIcxSGt/R6xkI/yzplWikX0nxoPV6+grQR4529GI4u1+W+0QEyJedlWuPPEzzM4cxp9Ch
dR56YEU+//kA2UbpNIlVl3K+51C748nwFDRYady17If5yVzm4ice8dwZXD0HT2G5r5OLSZWQTkIw
x2XGzRLbTsLCLZIQpVH8FK84OvBNQAlYluqFljYVT1xRB346frQHzeJLcBNkvnw+xaMYVBLo2xVX
l9tlu1BYt7cxpAU3ul+Ayhc0wcORs7XH6aoITiFXVg/TBofxANEvJYXRVVQncCMSVhmHooA2F+e+
RqTnOQ9Klfp+3RpRtz3XSIjGm64m8bsN5az6CGSBTBij2bO3zgbYOqKRn6njxpAw4jFC8q8o7gT/
HZiBPltj54fJPaD/TdIy9ssQYas5Pf64iZVAHkyFrm3xB8itMRclzacR9Eh+IrH0BNjHzHT1uB5I
d9827fDiBSWK9ypSRjjQRtW5qMjRCbCpb7Qlz9SRlMjn6tPHeXgcE/YWvoOZA3zCNS+OHmycAe12
kFPXO5KXrV2TIzcqLeS1UPEx33cOQ6urhOSth2s47cdMgkLyXmlHUnEGPSva6/tNoZ5xPVmaWkes
nUhcNj0zmbYHK2ENhQZr38POrFAvZ+EvZc6c1FLGA/TCoNYb95yxo/GmRr29PVbj1We8JNimgr46
4M01QQZ7+PsH59yuW0I0BbynxbB8xy1zyQ1F6ispaKo5Lcq+ishq0Aa91A8NoLU4dvOxZ6quI5mm
rK6BmVkiQnVbYm1RV5vudQNgcxIZjI0crWCUe08hFLJZGcZrH97P51oj2yXIaX5S5o5dNHJ2SDE6
LyaXzIk9CSJXibOfCrqtJqONHVa9gjrtGKOjSHWDjsE7UOHyO+cXOKyeSsL7yDmUUKvnkmGgEK8X
qcBfgmDGvj/61m1HFAbIuoIiX7X/YKoxIRJpOrHsJVYb1dYpA00IIj9FQj5Bl2cMWv/50f6uIwMT
uE+qaMpfZo8wbb8KAFPJK7tY8zRba3Rjrz2ZXdg6jRgUX5KG7Hsw9tggflUCJFn7YHojfVWstiDM
TS71YSErmaj33MFuE4XtcurxhqOdtajyTf3dhloq3ljN//2KOBZyrhTmAf5/HgdjZvsSjcMw9S4E
8wdwNkcdJJg2FOJn0rW7KDOPXWZasC8O8C14fOC9GEg1SeLF11HfvWjQcGBjJ4B2MD3XI74O7qzI
iE/I8ov0rTJ/2CqruPXgrNoUB0by4B1G94exuYhWd34iBPw7dg83Gc0a/yBgj7Wgmf/F2gFvbqiM
wwKY/B+ID3fjO8J01X75KWIEcC3hvMWEZRfVBVAjmAmt5kobKuMuiy9YMcJZCtL5MbIS7HfehsBS
rIh6GmhfartGqps2n+ihFCB7MytwQHX2MaU7wY0ITipchqDDTGt6pKVf0C0ssgmQfCYNEf7S2L2W
pJm1ZxPxvtM+n9V0YpH6G3e6m1V3gALsctEtiras8NvcIAIK/VNVvrBvt/TbslSaeNrCncR5sG1F
s+FeOoXcNR8jypAEkYEl9ygkoxo/le7t3Fc2UEXsL7Ks854ABRDlnq6LyPDLqIVKBCYPSVxFYYjo
FUhk3ptxhyqx9Y6pSurSeXDXLRktqpTP6LhBv6ltIk8JsoRyvYVXcnocU3vNwGQS6wwle0BNIMZp
OQUjm2sXpvcnapyOL7oN1A7QnL/SyafJipm7Z1z0o8HO3+HyA9lgcKqnlXuI9QmFm+/If7Wb0N4Z
crTwCU7jfSTkkOhyPWi5s4PaQAFVdPB19fr6tbri55n7GsuBA093kpTBrrcvX89yt+4Z3IFsLcq3
wLsLjHlqmy5NZ1sqHeE1TL2tuTe175CpuxxKVPdu+u0/0YwVN4XS751bdqWzHm7jZTBUSf7KXsHy
aj4u5KAzu/1GhPa/RrZn6N36LEaWjAaRqbk0yduDewI35Bm3XjxYio//PwtD0zcR07cqgjQwRW14
S/7fSgzn9ZIFkNwCX47Y80PmdGK37kbm8cHwzRvVkMe0/D2peSvZlFBsWauB8VhB+Oolr2AfmDIP
Lzj7m+zeoJ43EYOkIiDgjtokRFqlccenOOyB1u5VHja/c/u9grTl3FYxnVZZ0Ln5kiJZznu39LHc
p+B/YF6Nv5+2+nIf5c4Sv0C1ru3XsBf8nwImLyZA2kccFgR6pteJpJAkA04Lx9K/4sdQ+uTQsmOt
Zi8P3hByPMy65YCksI2z83SPfRq1P1Cpyz7ecNud3gqWo1nMRU8gJGf2a6uKKXU43+OZWPerxs4A
+eH8FMWC9URR2yREiNTSm0q6YtsgGpk8lwSYxmE92TLYMpZhjy24M1A43nncFyqi6OeDiK0fl9qc
SCyUkgjLnvJscZQivCoFWWtwjrB/B3rHNvX10L3rbOSQzfM/WsJ7fc1RyQIkyba2qgfKPSlhgtLD
J2zyLmHboAbKaY3uHlm5OIDAzbaNSDCkmVJMwZTFWhX1BJtkwupCFOyScLghSB0caM1z8SmXgEy3
QNPWkHLf/glG2rfy/nXgREKn94g0Lh2RzaPveqWh4jhIgDVzRe2NNgRwSFmxFkmBLSayTLfVSRdF
RCx1FEMj6xZveMFpOwB3Ya13wnQWzH7YbKo6o7w4UiKheshgOdpN+7Z4hjkH0B237ySDhaMrS1Ro
aIPeeu3L4/Ld+4erqzwHPC02V7JHAm4qa3y67k6qWsvcg+o6jYuwgtgABtt6rcVdY00cL4B029oZ
9WgeG7jsqAKc9JgUf0W8URr/wITHZZEGvw3Qbxn5khX4q0qpXfRFAZhAPxgtEcmAxTgGZAj2cX3Q
b8ux157zOTtA4hkRy5fyG2ZpRxxiuIb3oWs4SAjs7zyRIYMIvE56S15OYL7da13a6PdsnZDdNQiy
+nQJZ1Otp1mEvfoVMGOQYGf1WW2B9SnFWLYxBXmv/doMUGdIK5S6Y3dGamTkgPVhgcRcBn0WY3a6
eqqIAUPhifeV8NJ+5iN/At/sjuVb15wK9nlnH1oEdXLnjQwmi6rHoB22U+sLiEDTWxUVXgZdZKe8
SMvJac42pd3KW++Ri5+eQ9i9d2gw8Vhfi/0rK2/zVUGFbKRtGHZBg1ffwaqiuyBfehSb1WLcyAnL
KS42yGdJl193KlqIqOa7NjnB8cvKv4mi236G7c/XQURGe/NBgZS/lbPrpBEkv8I8raIAK01cQFkP
GC5qqQX4tw5VObHjTb4hVtPjlTw8MppxRi3d8b4DCNDZ/SkNQQgg7y1OEMjRiXlm5z/IyMHX+ZoY
ajr8mCaKyPMo0s4Ph+Rwa3W5yGCCEn2TpryXwji8iDiiPTaCvXX84rkFWH7gukGIj4CPnIGB3xvR
jBopNfOeKJBI+WMTeQLt9nNdDxOBoPsRcgxFfw2wdCIIAm5oJP87CBw8tHu2K0ALf4lY7YDD6bX0
dt1dS441jtqQEKSHtWfdd0CTwdafKqwW6WEWUYZJkhCxgEX3vFCpHIdfp1EYFsojCdXz/hpRB2mF
yZbo+dGi7iMGjcM/w8gEmkjDbpAkYVG2otaT4ESQuW0MJI3gsMyoPOZLIoUMgTpcjj1pnye8ZCCm
uZc+fFLx5t/h2FHS+zbpNM1gh96nXtRoVK2Fd9BpCN1/XxIxaGijf5KT5ZWixx/enzoqad2SjATJ
PGrwFMt44s4zSXHzvw08zGSqvfcPAiLpAJot84PUVL9agn1JyTHGjcWHhB+2P+dON04yJY2W9hIW
xMgKGyLEmu4OvG+LYJ5Ffe2P797aZyqsQ6SYFccoh54cWjjb52GcoqvKbAf0n1Z7zAdxsDKzSqTO
+yilrJXOI3Zwl5hOqu2OZknt/fA59X1IAxDykIa3kvnh0VCOFbHGjI/et86eaZG+xK28DeFqPt6H
4ZI7q32Fh1OMt0RVOEAnck7jAIOXXRQIWPvD2l63P8D9WZfFuzxcEy8YRorMY5rNDeJZH3xD+vAd
6WyjroZMGPCk0PY1b5Pn3STpjVt7HpUEn9K9PVibv3h3oqOHqB3Wu/e9EoET4MSp9FqwY73K9SBF
0791lM9zgcACQP/RPezy6A3x9r4NHOe1+VTLxM+FH6iBvjNq8WvP9raUuyCo5CN1mVI9JUL4TcGl
fdGIm+FMoZleN7Lxa2wla5edmyYjmjEcUzjEWK8ODCLEug0M9mFiUei1kby08Bq47RDdAZ2/fU6x
DztxLY1G/Dm6/5inRXSc+joZOTEPAmlEWOchjLo3I2Mx5aopXJ69tKLnUDeCxz0kopEvXoP/RB7O
U28555CyMPv5eQ477Kl0ADc6/WnwS0JCx3pkwtFJRz0hEjyyI4+EKcAX2eD4Nc+xZdoqWBOuS60I
4U75rizEXIJ4FBL5UxLCavX/2a3p1d5MH0yFkvW42ypR4hA+V7fFZheCbICmOSlYCJn/2kchXwBo
kuuTSVd5gvZZDlmxI32RWZ2c45m3nVkQZGDfuQGDjYqZe96TnJ95N4HPtjkj2ydxFHOXaDYrzmkD
xB6hNrq8d9bO4jqMpO0imHfv+FMbbE1cZmJ/uiDm11XJcVo7O0/2gzqSjHVBlM5jUQHdYnVualXO
QSzPBbzYEJoieXdNPlV+8ahauMyB66yGDAPLCa17l+EpsPvdTOHQpGG1ubV8tSkr65ll3cvumYnX
OfNIXxidC8/j0U5HfcwJLxr1S05KmGE5tEGEl58wKn7X7UoKWrk0fYVbyLUBBbpqNXZ0hSUfmA1y
aKehxTce8S/T8PhdHd95jH9/vTVNOoRQPX69oLZamgI9UCT45q0EH+8ztoApWzvShz4IftJYkbum
IURj/iolucuMdYRmmscxwGGRz+r3KdAittn4AOcElzD8vB3oGWpfZ2BJSdItLaG6G6yDCA74UDPA
IGOEtZIRe4WEDzWmt+Ou+hEt1ThEVYy/BQd2sASK8SUm7LOSpFaoLbnKRJ4vZqcn9qtBEXlH/Nwn
Vtq4+Tb6hiJmX8TPFfvOkKjNp/LXl+RTJmwh52PqJScCfgr4YmBAYAQ1eZvYWcO3vk+LHUeM1klE
4LgpGTfJskI/RLFbRwdj00o0F4xx/zT26tvUg7cXxuFg72jOJJe90U71ZbrV1uzHS+Ym2nT3O7bB
X4lACRJhhSBKRdjbuDohpX3gL8E+jvGI+xdy+BWLisyazx0xmfQpCS1FUKLBJNEuxgbUo74S2srW
9bAAqIsZ2tYwztsGaI15p3leRo2Y6vYtEQW73uHhh6bQSsvdb9v9hN7OuRdXtzHwPcOuS2vVpg03
xiH4DewjBcPB9tC89IlmzPFINJOZTAm+UdaDzV+A7KUfvx/IECIB/GwIfjBcUQ/EWUiUOj9gG/ad
49ClYlprL5kbH7dzbR1dmeN50jRL9J3Y75xRN8f1sO1I8Xl163ZARNYQck/3kBaqBNqFvkpaHf1F
pqrGciM6U11yt6n6sWRMTnU1gnway3ibpwDhVMsACotr/DsepjtTMrPp8LwVl9qd7bpyI3uZUMB7
GKCO8+CtPQqFmpqZ6ZPt81QzNVJCUmli8C8Gw2iYv+Un9CKTHqseC9VdZLrgczcIyZ/qGLE0Vy8x
VyqogAN0U54gW22pESmD7GqDkcTJIB4U+88wZXJdRYS2zs50aOGVsaE3MoPUCs603v8rHA0XEPtT
Z8qkd/n4eigtRb+PVsSbPNuCaVZ+0AFG87Q/DVXbjzsyTMrh8t5ejJU4OPI9oVUpItY2rZOHGYqB
1D7mggeTDFfewDCtuar9k0AxJu7nROJaT0QVxiJ3WocdE5kWDBNqH9tIFSbidALd7GrVwNSIuhpo
w3nuD+240pUbGCisW1UepDwFyMoq9NTZXS/zCqqMKVwa/2msIoQmVRjOWoTHASxw9qWoxWa0BGvy
151icDeu3qz2THyX4G3IpoR91X3CFP051MsNxP+1IfjVJOQBy620qrF/ceuCq+HkCtcxNf80UCj/
Os0VvaO6Qh7hFFyDoJCuiT8unG9YJDoY/4oFPWpD9itW25r8My2MWcSZLDrVP3Byd/txGZ0fnRQI
j4OP4isyM9f86/mcZDu/QeulPP/PGf3frRlUHLOELMhfsVDA5IvXnvnbh27v1+Npz0rgV6MpXUYe
nxPAh2jpM2gVS6jvhJdxS6k6lrQmuOZysmjygg5TdDZe+/gp5zFSQ8rlvTrHpGDxSXB8T/DQgCmf
aPphST97xNYx0qivy4HD1SfnP2rjknR9KbYR1o4WufM/bL0Fwke4Y5mWq/v6xmknOuVPbNsBhuIt
V8UDSu6YJgqVdSeOqSVvX7ChtojQuw8SjnbQnYLKLZ4r/eiOUqbJ51NidKtWSJZZwVPlEWfkVQ3v
SXJFx78aPCZy9rSBWsj1zRNSY5HRi1Y491+tF6trZGbshh07DP76FMu/lUQRc9d4/madgWrUvz/M
+3pQYWLEo6D4D63uIsa4sVHaaAPW9vkHx9PDUwPwPp5g4YitTcO1UFbdpgMI1tBy9ksp1szVKV0n
Jn1i0SwGndZNx4swVoBG72UdvQdqkkR2yJWvtR5CRIvMastlvWgwUCgbg/HYtN6annbrmWz5pi38
cYGkS18+ffs8OkhZ4DWsZH+r/8Qd6Xe2bbASHFhwu0c2fncD2u3H6bl+wNsPmiJXIRLVIa2+WQ0u
WTfx1D/Inr+pVwtcH7YFbCqVtxj0vHCDRb8Rs2ViCtR5i9Chf61m9xOSfMZuGXXRrQmE3eON2fE4
On9xRTaQPQFDPoyrSTLrYupdINknyjqtsm+UQf/zoN8Fpf8CujOLyjYbr1gSOfkBSgzdUUgdATiw
2yRQuF2WFG4ftnyepLBFPFMiBCyoaJ4waxkk21ezFDr4oEIwpa3dxOK0u6uwSzNXMBL18wduSZ0A
L1jOqghAQhZS2kJDSOmQ5LqqGWnovXMbABdCWPPVQ7CwceE/yUGHvgTh2/MB53ztnq/kvWYWheEX
n5EZZScXaQqIVC/7f+u2H/kgAI4I0hu44I7V3Bmq/2f5K6UsSd8tMA9nKGDJQ/lEFsq9waqDvapu
5lFfwCWYZ/AZvzQJuG0eztL0ziRbibQV6FgW5ZvDgLmBKVsZFjPafZKD1BxSbOODJb4zFsIegMGm
XniTLTQSdN0QB7u4MSn+1EegKsyHqOGm8YGTGmnoh55dJBt81/b9iYogKnoOdNYwhmyQBPwKmLJF
6O/GFIBNHHP6Q+dUgg5ivZttK7V+3AC1MT6aOTNAtDMw6C0B2+le79wVPDVHZNqJBUTXuFADt4mr
Hu1elRND80NJS5JtMXB7/LAZeVAK9SRmRVOKVTsiD7ErpmzIXdm13wI3jhol5+8jist+XhG5i14Q
vin6PBFCKeBKBbJNydSvvSj/OMbQF+sMNFjVP0qtn/BiX6w7quJ1Utf430VrdnkDyvY2t6qoGzks
Rpn1f9FFkfAU1usd6BF+VFNuKOYTDHQmiYyZn0zaFNuFzcFOxkRRA8/P9CXwaFxkE8TXYxytpVvD
lJpOWmpFoW3b7EToQJ9V/z+eWjQHm1ChMm3gwz3APAZQuaTtyTyDQz1bg8JF3hKfjRMqPHtycyv4
hPbAmmhXyVQzxsWKu8Z0HiWErM1qswu/z2ktgP/0VS/e3YAjYFLLJPuRVHEvSISFNGH/lzUVinf1
EVQZOKgeeiDGxkHTQXiH+nI8JcLa0r6S01zEBTOrqt1uQs9lkRzWSYHXDiZBlbVb+WQqSJm5i+aD
WYdJenndVf+OnkGsqgp3cJiz7CtZsOTPpIXZwarqjYXg4MTtJDX/mqpRKRfGfZoS/hYmGvsK+lcK
ehB7cv5dvNlrWF7Pq4+vdZzwBm05cVXD16Sza+fa38novRqZSRb2oUQkOfKPu5IcHBvT1lIr2SzY
8We8zV0RvlzNRMEI4h0TyAadiONLHG5iNsmnoQZ5GmKjS27UIWcHUYAVG29h7NrNcwrhIxntUe3q
smVLgmU6oA52/r389Zd2QPldGsz27jgrYPiX3R8TUFDGGxkp0kCblaUONt5KI05GtfsdfPsCg865
LFHw85NRkVAnXoSd24NCIbQP5qpbNhff//yo1LHeXOVIG4yLWrRZDUcTFMmNiUT6HpM4+oxgdyRo
C8l8RyQCoYSSbifjwGX55MRKVnLUBrFctNBQn2axxUcCokrh7DmzbZ8S4PQ/8JLjsFskI7dedwOa
1bDpQrXRZ8GUBAVCxJmIraYCG4rQcTTRrXFF9VJXc9sYvhHy3L0geNGd4Ljg9X2jVknDJfIj+yKX
2+zG2D+37H11ehqnhnI4k9lnNIaZP+brDNdItjtKNZ9MVbeuQ7Q0X5NG9bO79wie6+sTvQ/wBoer
bqOJUq3uF04ea36Fopphuznz2crt/qtjzf/4954OaQxHHdW+xMhyKNrkxRMES2rhRanEDrfZsPn/
pOjYgMZyFLo+S/zE5g4VGYQkZ0BAIWTJywPT+tgAws4HR4VztwXd0RGI+fK2+DalXzjwxpOxHBJE
mWYUD5GmYerrDbwjNKTYUNW/DC1iffESPiMntOps5e3QV96n3gmzt9FwnDdSLmOEdhwCSmo/vm4r
LoRn2I4ByrMdykQge4Wt1lHae0Jsa0/DKrJ2EryG60y83VAJ8rAwv9bUyW608kNUWJbW0ko65LiT
dr99gIVIPmYllHDCDblxtwVeZTILqsRLJNqolC965BIVhDimAPgJmGUqVSfRJrRTuT/KLh52ZsQ+
Ld2Zpa6wwfYw+UjehcvEQ714mxTr7XSHWL+h9u+ifaRUZ2jXACGMPxANQYQMut87czL3wG1S5NH4
69SvrBkSVoV34jLInPzsUcVvD03pdkbIY9tjCBSGgRxDiHTQ305VIfUZrD1WKbO/2dUtm6r2bVPr
UNVJ43cm8Kb6ifPCk9aLdU0eeRMdI6hbbrVBbIS+SnKluLHsmJ+v3F5DUIQcFAX8zOVC8uoDat5e
5KbJfDp7V9TdYNB3sl69CsZRA6PMAPph6LcO5RCXqiP2qHM9qQTASclJRCOOR73u0/st0NOpFrk3
t+6X5XyfMLlDGbhj8UCtgbcrsC9K6rVBuHhTnN5k6CxCrNTChadijKd02fmGjz8FqsKLTWrDJXWr
MTwUc9Gzx3EP7tBENYBiU0jwF8Sx4pXRRZuWQR7CLcwUxfNT5StFQTr1PQvGKZNiAW1ZXCoz5WMY
7qQubjgdvLvVapyaanWJ2nelwyV4448NSt5P2mDWqRXMhTACz4Xe8J7bFFcIYiw3ezebYIXUyY4Z
dPbqj7pG2la66WrRn4HJH3xbASAlvNHdsWz5P4hLHhlttTadvBibB7/6X0V9t3tV5g/WOGdaZMJU
5jaocHL0FKwmVCmQFuESVrA9p3vPJIoEpUEl5AbzefkJy7ILJFdFnL23XP2p9eDGCa+PTnXYVQkg
xjUXd2zW0ySF0fbAPKHJwzpAsX1LdWQNAR0aNOYxdM7da0lVGcNC/FBHi9eCVLivGTJ0ppMD4jiz
gnFtXYXsYzQQJ98GxZBbLecn5vwK2PQHLLSp0CpCdHL59U68GIMPdPXqiM/lFo3qwKvMcQn6vuZb
+fq1M6oDHj2amOIW+y+9NlpCz7yugogSglr5p2lYTED/j2y2pbzxnc0ZkyqdK8K1P4zlH+Dk5iUz
Gubv3BXo1KSdYtisUA8GxaYruwy+rbq3FmUpq6U5Ng9LfYxsOhiOJxNSxEDYKan6ALtXfM5mT87h
9QYd8MbP5KCQ3JxKrkK1ovNqOthhkeItaA2H79Hp6UoQMX/ZDrt3xA9/LWIpvVECX+Pw0qGQGG25
OJe8udsITXQGiqhBRJcfXARX4gSqFFwR9j+6HgmQVWfcFa0L15kpKBWs9K3XSyF6idx0G+2nAMhD
N6wwY6hYiEPC0huaV4jwo/941WwY6Lg2E44/XaiUH1iT2Cbe4kcWKjQ6pYqt4BrSSL6/28qatQAA
w8Y5EF/hIxZJtsg4P2Ew2KULzkwDgyAykpnQww1JVor/23tEu9VoOxpRqHm6HMZv5mwztnnir0Mp
qWBOBlpBnNTp0SmIiItLLnX1ntDEIu1WxpLpzV+n/dNbesvlaDADViBjpqXOmH2LTcH+gwc9Pbzc
a/m0eDF/jdS5894FSxlEMhf+kEIWyX5b8flxA5RAu6kQv1t8R8cpsQ9Vv82VXtOApL0HIQijJQR9
JStIrS8butTJI10iy3D07T+CaUyJTSMPwXiphqVI5Oex2S2PvIw2Ye9kn1n6kJIBNKhrcm9bIDrL
Xv2ui8Cot3+UDNxRq15V5ZgFaJ14VpBQueTJFhnNQDwiz/tyWCH3haH/wKjDMiHKWvuhzkO2WxyP
2fCocy7vqYQmORUsugfvJUCN8XbYFt35FwdebwfgsDHyAAt3CTr9cG0zYcqVrUJ5g72YelFi9srA
AUbXTMgLcFOAvSOCU8LHLs8ZGv82wpLRAgNSOYdL3RJPIr8nq5aTEUXqptzptaZgAGPz88ZG0lEo
878iYlo/slHB6kbSAG5UguDDfWRXJc1l/Sf+Hr8FT4nojDU3sATY2MA8+ZjJdYfbfgGyK9hpbtKL
hTayD80BEV6dj5Fq765QjdQU/ujealHDaZzbVp9wzppQQ3jS/PAQ152y3ccQKmOkH7IGSCVl8ccJ
ufslyyzTc4iRClSJ12lc8jBuQCiJcEmMrKkjxzg/qYqI93orzlBGiG0jhzqFeP3vSPgvo2Y2ZxXg
iPyB9Vn6z3cqjc2PhCHTl39Qab5qqMSvqefq9rcrpBvEDt2VpgRviS14c+CHLwidCnh+qnrR8/6Q
nNUKGgSlnWw6JFZn/RMxyFT66dxaGZVZ4Lo12jyk2Q7udz3WDzvpqEy1rIatO5Ar8j9AEaHfxnrB
VBEpiAGvkCUp6oG2ZuVljVqObsbBkHVlrGTEjZZ0l+i3uwzxNKkjLc+UMROsdB0DArxtmSoGyX3d
UhGW9D5GO6693iQEwZdwwG9XI8R+zYRozYgbDYWiyCTFmhcppB2MrWnrJY5iPnpbRHRd/R9pqL0s
ZVoT9ZYFkD0iJec+npIKMBmDcOoDQvN+hDXmcv2R5eAlWF8bW5yPCT2iF73upMvg6KlTmgAvanFX
xgDCxpC9c1MJQbYkB1frYFyY9YG0EwNyhNscMSsDC0y75tolrizx2chB/UZvmC3foypVQuEq6Cwj
CZSOvqzcUOgx0WiHq6Lni7CHF5yokKPW2S+dhY5ndQ/nOouStksALbUYt+0EXg5ilEe5dEmcIp7k
b5UINaFOgWl5ulgZJRYuwCLI3qqaqVHNXyVC9il0CZgKwcN8kmPM1VLIf+5NgKTfvmPl60tAK7CB
Cb69tKKPPJ/GMJ7sOYCmFg2eEi3EjC2kSUwnYXAEIORVjHhx9dQ+599wm3L5ZKgUyL0j+QM2G8gM
H1eYlhTbISTefUJpSXAnxUyRgomej3/uFk8GdGAqLAkGJBpy8ySv5hm6D/mJrloYPGD0IfD0edZ5
uf739kwpVFsNbesSXO7cDFQqfebLGmzhv76Ioc/Tpvs7xsPN53kWzStke4+UGLWSWeBt8VzRT7QQ
tBIhrBZP6l5181xgv+6IwE9mCRrRZaIGp97sOp5PMoaJYfOlED1pdKnkxsrEithV4aTZ5hyHsgLO
oqJkCvaVJaqH+7i3ysJwoVq+kg0H/e9ccCwEs9mGIXygu09CH7NFL/2Yvu0qSB6ulWMYXS+lKYmb
jRZjvOz65YIdpxoMGbSd+SVmTydBDDcpmZV5v3oJwnVn4wTV+iuk0Dk/L4IyfLIjk0CPMEW8fKpg
zOJNikzgTfONl4hnLTh12+mSYzxWTiximoejqEdKNtgIhoUpkXYjK56GEsqFMYLbBLRxfCyLEO4o
F9Cvm7zuDXjolZti4Kb20u1e3qXgH+adM6Kt++5hRALnOXEcTfhGJgICRwcljUL5f6G2T98oebwl
GMNM4xBpBNzuIAniDiChbBPzJmmqoddT9UyV7Kjw/HszOdsn6B4oNa9xtmTWLJunU6HGAcJ9rHmj
WJ8NvMOUMYUL81e9zqp2gwSWKy8LEqLXabI/Aa/fvFSY5FY9gi384+jZjWm7ODJs8DRitrF8vrj9
YmJ0AfnXjvphhaOLlAkrTHH7XP6vBk6u15lUnlOjyg57yL0CdaHLvQO7Giz0xjQ59gMiuFMTGMNs
SWOnltHTBcRroyWdM3G7LMXlZS5L18ruCBMU9GRLPeqM5rTeDF3Ry7nv8na0iLkIJuP1y2Xqpcu6
OgkE3fzE57wG/Zij7quWDLnJ5ejDk+9TO6yPhTfjNWBIiQmL3OeBkPWmD2Z9g9GxKHTZJJVmWwEX
JyOeeecnYE6B67mngquXCR7+fjZE2hhgj/EXZfgoGn3ghueGAeYzMY4LSviWpadwIywBeH+AF/EN
zLg5+MmfF0gyMn5XZR2iY/icKbfQDuh/f0k5vz/MJQH0AQiVjW3ovx5P6J9qQVs4ZH+m7VXVl1cP
18ogHx6EWiWx70EcRIntNdQpcd6g69tLJHn82GtIlbYqsf9X1VKWOOIyYu0FApbxCyEagw1BqSFV
TfWTwQ6rjFy/8q3KK8Di229Zg0P2uiUTr5kVTAVVwuwvH16OUs0do464O8n2SuOua9OL4Fnd7HIF
9YnZj9ZNBgxXV8vCA/BgFEI/AMnOf4SnBxbTlW9wCJin578zs17f0Dfg5jdA99IdFAO24wLaZta4
AO5g1mAq0lC/cay2FgTcmn5ixWiDLphmldbOfWnsRGir5TFgNdzVqGC9+Vf0bINEsG6MlEO5IxB4
eyvZgLiHaVauRm3FIypEtY4IPzbPvcnTHufeSwxf1QnfF7OmxSqDQEhie6Bab+yQGnjJk0tMxtkx
VOG0KLLctOHEzI4n2BtAvIhbdKZLPLZoOegT2JVJ0I5/YXQPMX3MkKb4xmpwQBeSkSOYYXdsZxH0
nBKKWBxEI01eSYFTwD7hElbAqYJ4rd9C3X7+JbkEYZqljIdXhCsEud0OdaGQDqi1OnTP/QXY7FyW
RgAmBs5qEccpSPX/Qc0r6tfAfxPNjmkfcM/kBeWDg0hW6ZLoEHRBNHgLsDCozNNzFWez57rgUc93
StwvMBk5+ynD2GcEKrmETYo+vOXAx3taDPy3oBQVyAo6pFUJy7hKKfT2YnB4kd39yNq0ZfIsLy8A
N9MuZMCN0LD5nw/4V1XwvKZfINE8s4XTuPlRbRdJifCwQWB9BAHj3pknbX0zHWneAJk8yqpyV7WN
z51jscAfU6mYfhQPizjb3QPVvCJ/HpOSKZJjuczuyOE8He+NBjSMd5JZKFWAS9Jpm+rbfE7kxinM
wU8GFt1NlqIysxirSO/J/rGYlbry67+n7iJmuLip3uqz+1tTRigjN+3GL6vxYh1pp4VZZCDiRzNg
BYFx/TbRkB/ApkkTA2bu3TJUzh3kpT8j4tNsrf5ip6AIvjoKZxKnK6iiCy08ZbOFDigAzmZZXFg3
J0LwJImjQLvL2+STaur+yIN6kXrj6Z7xVJxpOOhNE+RsCcNS/vsY6k89vDSOX6qftfhwrX4bUcdW
285qb90DCSVC6Rw1c2LHli8CmrlnN25jzKTCQDNsKUSuwqR2CdCN2PTxSZdqYWRyndtuGCgCb+j4
UUdApvTVxLo30+8AJI6A97drv7VdljIjkoldcIR+H9+Esb4k6kSDizhge6jAin3swmtAeO+m1+2E
W50Up+q7OXqOWFERVe7rSuvDbn4mebI70urdK68pI03uR11JHYakVJCjNsttw7XCBounjEBRt+fE
cpBX4nvfj1x6TV3Nm5vRQkF5S6zhQyZ2Nbp88JKi6uitfqhCzfI5K/S/gFZ1Hd2i3m/Z8A1D7WgM
XkY/EiZzQ0oIhf/kXdLAGgCF6EUTzkaVv+BIi8V8YHhXt5ZuYQ1aAlDNi4Cstfv5VzVjHmw6PBSI
oK4ShNYPVGlwsL+oVGwtbd5WFjy2/ylsN3FbHqYtFtU2EHR8VvN5Fqsvp34ZlS4rPrPjsPFTdo6t
mXk6hEepsIIWjRbiQGwXm2JMYzdo6JlRBgrS2dET/JWmnJLiljJSQHJclwxGHGpeMnUwWEuQJKKX
Mi8y9CHa1frIibEcpjjOQi2tReMXeWaa5bdwVNighGdv178UTQm9Y7edVW1QTH0ZpZ4/7lt+CeJa
oPr6PXJtdE9ol+SWHAeFXs1m7JT6/Jpz3Vi1HN4Veyxv2lTyBHZ35ZoBGh04GDJevIUXr9L/cqVg
vFcjKQUreyYpOGvyn63LKCQIZOdh4Yl9M1RQDbB045WDWy8fxOAVYt6IvRWUieazfoJA7gY4RU6y
3lno7OcWkopOoMJe2L147wyRWqIveZh6LhhcZ3DnR6LW2/vKGDzd23LKY5jbSG5mcLucAGoed2HX
Dw0MMODWcyc//ljPJVYgFWxRFeK9K5Q7v0V+czQaBG/K9q1lAjAvry/5ckTn6rSLIP3IWxerjNdw
4BfD43suTBzVFAk1WM43nUXmj2awugjykZnIFfuM30LCZMM8DycRuday95Sq3W1NdfERi0bCstjh
8Z2hmLKR+afMjo6UmDYJfySEGNv6xD8L1qZQ+5WHcrzMzYYEuJGEJAJ6RWZ3MZ1n3bGmRzMH1VZA
Xgo/KECuM2Fjc/Lcg05x8OdFYnO8+gDwFMIx3BscgBUQmSuMO6ZA9pkAObpPYvCdR67iYrKhlbxB
agfBvLJmR18mtYQ7XNb8TXMQtOijKLBgDs30l5V5Irmb4m2Q8CgL1faVJP1Xc2H1lls9nmooPk5Y
YJyya8CqoP5g2km947MiGdS1tNX1wfMR2aTbbJSq9BpEqIJurzkQrRybOeMerXqH7aF7tgjQHY3y
ZxDrl7RoaoaDwDHTvJkOqd+jfdHu0cBHqz33Ttllo+qfIov6MdoZhkgX/2eFjMQn9EPCxuvTac9c
tgTINf4/j2VY65c/3rkvPRmHk4mLDDyQpKBTxoCZdAe7kxQ3BqctSQ2jr4CfhMEMuskiouBB/XMV
J2PE6ECO+9h7DIn6SuVMFn1d257pxgPw53M6dCu3nFJJfq7UGG0buq8BRdqs8H+CKOBaj7nFVEt2
HZD7rVSTPdgdmC1aMrBOTKvjDrmoWaluCzglGXY4IhsoNivZelNjoqty/xSRwq+U/TI2OQ9Hcdr4
ADRNh9F/xgNZMa0tJ85pYEpgV5HOgig8w7JtxOUF8IMve2OU6g1cSvJmXY+ahvs7beRYjtK8pBSX
sv/Bg3LrZDMtzPoV9qxnsGBGbBnuIQdBPTOrartvRqvw9tX+o7+piZ1AnGWI2HI6iFwQQ+IUFxy/
pG28aGbVLr87lFeRkc8K8jh4zhI2OITqqGM5Shx4kJ/igo+0xEsczpXuRVXbMN1fYZ5AYVlh3U3E
g+b/8fqNKeWwdRrMDRJnRtv0oWINLuIb23Ek87151zxM+4Nv4wIOmxwOsX6AwhPsUh6duj4LXl3z
Kln5XsLNg15NMA7/y9V+ryxtT1mSFY556T7Giw027rbAJflpdcwAVF0L1aay+KqbA5s2N50BSjR2
u2hWMvQfXL686uWddNSgXxCxq6/BRHEdFUJWny8Uf/m88u8/1rWnFn1S1sy8nsNl7aXJaBe4jlDr
QmSLmtkwj++tL23IQTq4m1WUF0sTc144x+WBtMLXq+yWpioLyXAnYV44eiQcrS0ca35cvYeIKlzJ
Q87L2297jNsXgIuo+XbgTMKPzF8fAjbhoOcAxakK8wiZVBafBDrrmxajdg6f6+Toh8EUv84USG85
Gw2uZcqYkh+vD6aZLzjgMp/2hGAPldueWM+fKVArcPrYktEVucGqyesAyjATa/dlw46mQg/GPQ9z
L/V+YlCMa6Nu/shX8tc9wQB6XSIrSYVtgRdYAPZnWWdTGS8Ij9T9kXtYOUaCAEbv+Gr25RKMRgzs
oxLrsd11JEV1wcTh6pYRDenrfhD04HRF3xULQDVlAtqMU8sRCfUQKmhFGXAEnM5QGXz0n6r0ayaL
kC6suO23/p7Q0JyCIr+XF4RRCbOv4sHdsqoKadzSt6ohBzVZj8JII5FS86ckC817+L/lDOWRz6Zn
2TMVuIKzfmf7ALoCS4jc9rKL3sSw/lAi0x0vlYZ4Vf9Qfveid9/nttRPpvmnVEGs/aSUCyxfnL+q
DD/cTdV/KOZy2FaTFgzyMxVRQpcS+Ki2ZqApZzjQtdbt3ASoIykYihe/jOUpwMHd4nG9gMIB1QOI
qWWUZm3AMV2CaC1OiNDQJNjqvphcUNIHZ6PH6gwxOQErBxhHcGGynw2V5wgynptF7ZWK2fJQbDk7
pIqVelAhKU+PM1yb+TAdm02ywWBJKyviSeYYuU5BIpplnZ7gPXj5KwyQQ3M5Kphxo252aPp3toj1
9dpE5fW7im7AFiSxBPK5Wb2WGIbCLvmQcV5mlazKl/9iQ1opNhFgpKx8a3AUPPhJz+S6lZDxddRq
lTXF/EHvfRN7ValibYYEmAQKMOWk+ofyhPwA71t97gG8dU5/FJ5Ag1ROW87+Oi6uJ+PoogHMtwK9
+ErszbghEH34o8GeqgKpYXWj9kyhhbxZ9E7WgpIXueS3V7tRAmAeKMYdF1SMASLkvcb+pvJQIlYt
/ZWstzc7gquTqEV38X4Na4Ra9ZeWh1fmAeBbnYBmh7ucHKFBRsjoumJukGq+8Fk4e6UMIhNxySYl
l43JQG9xG3MuTS+RRKNAA4n6/9BuSKUNByr0ImNQ59E8CjpR0kSvhZ5PbgU5im383HoE1fpPqB8Y
8qjEBFnzlf82P3utUOET3C5URMoJCFMekRa2ag+BmhGBh4YQBEbF0hdtFB26Tt8bvfjcw2yeebWP
L2Fso5aYA1iTXj1bZv4vy5n8QbcP0nPW7VG7ZopdHm2jHgX7tJULH3E88KsLl3QBBiM74/teIvf5
CeHyaQlBNryHXskZ14sCtzBibaRRaHas5yzsZusglrSK4TH+p1CU6HC+cXTjjD0hpBb6B73QG9p8
tZijmOxvO1sYGny1zi2XsmySUVDySi+YHQCaXvY2Lq0ACrgZJWtS4bQkSh5gnh+7bFaHhQW5gOVQ
84HTlhwwCXntAqZdAspk/OCfB37z92lJ65EYa/MzPh9kA+093SiRP17Szc/38bwG5HEq1OPHVLwb
YgDplnS+A0YIg4eZYV50CGObcUHLv2xAvZjCEbeCLUCKZpEDPnekpURg/dZ8MmwBBHW+Gnk0675/
07mRpR6/za2VRqsWM93fCHEP4NY7nvpG1eooaAqzEONBilZfi0Zz4oXWA1ytU2uhDN8UW2yot6sP
GgnIOhBe1VcDHooCopC6CzY+IBWKvI1BGJAYeJ6jOEPS21So/SWDjk7M+k6odCzKQn12HzyVnhzh
4VOZx9hHl2sb1EDqjJaMBLkhS75pAzcX/Jm9dLrMd69mQVDgmTRJOZHNaAdP3k7+Fed4BYMex3fm
RCn/GttVktIte5lt4LxHG+mYDtugnDKQ5ANtFK/cuQgt68lnleDWURE07ad+xbpWWkLDSdikwFP6
uC6XBRYp8NAMSJ0T6gohYmoi77owga9VgliLBgoiCoWE7uxTNSTh5gL9a8dU/aNadcTqxSx2TB7j
aNr1ltfQfV1wrWRxO7DBF+mfblrKZSgNMBvw88CnziuLZdloAlHsk6BonAsTT3C0bb5GHxsSAJ6i
cPC2fD56y3VwYXx4yhm48oqwrBUg9NEPg8o5T4H70HsOtAZPBDb6cVxTrZOupFokVkRX5UZ6Auu4
QEcrw4pEA29QsCoNxhmvy8A8CRFn9tr+IDOz3olGqZcSb3Dwr3EDNgVGi4JXC3kTArCwF74Rccln
R079TkoYv70Rn2IJvmO2k/f7b+Rg5EOtcsv9wtLvw+K3fdD7U92gERRyOWMdmraXkKdMDpoQPPG9
iCUMEClIx4iMM8CYVTaqfbq7zKjkWbQWP7IzD3c9roqKb71ppem14+pzolICjFnt1Eh7SDUdYTIt
JBAlSpI09P3WNf0aCehJAsjDfFsJWd/F/sbZOLL4VjuCH6Yx8G8kvNjgvkI8cYEqF0s4PfbaNaGq
JYeHJ+8tHncyiGapM7wavW60j9iXGUwgZc6TcChiAvc8xjfFq5Wc4xVvtZSIbD8hQSuYoP32344Z
n4AkPzJh5kAD9NCXVzgvTzW8XdvMrQm78HJYjZTpqK74QW2EVn1T7acZST+uAhozYTw0ZPaFo587
xrGfgy2vhrDmjCkDfG+quy7i/dHzXMdIRDXM1ejl4CalfnZJ5bWjCNA9kV9u79/k6VDd4CTMg2C5
CaISnWT48rgOBypv0Xo8kiHF/rd0oifuLZNRlZvPDJGNXRo7D8ElrSwEznx0vFQRHKLRzm1rgExV
mLLIjjB8Irof8iNV4gys3kerKvCVedCTKxDLxxs8ICdz0Lu7BshII5qyTJ+Vg+CEkzfOelETBKbq
ubjmZYQ3alxYsoNKXCwDmJcTk2QSNJZGzk7maINM0eYz4Y/eWReU5aJOAfP2IR/RWv/YH21su71F
F4xY6XLLAVJ+Y6paPk6MhHdrCWIbkX3Lr2kAXJitv431yZdxA2XC0M76irr2lcpEeFFizqZaS1BX
3z00arOUSgMt75CXzBpQAqdYIUm4wRvP2HzL31sV/NjHnuil40jgctpCJt494buyDZUGsMYQB6j3
y7GiVIELk93maY6rM3uzgx0gB8eLB3r0HMvGMjTpj+2qP0X+sXSSx+E1M5+b2q/1yk3qhSSW2oh9
d9KAK3q8LRcBCGDonuZW1mqasrOM1AIqRq4NbhTKcQnatu8oMIAVaCFlUuCrhiBkjU1CsZwth6Aj
Ly9j/iBOrKGSh+xfx0QxBWCDxnh3q1j6nuup8HIKvhc2aG4LAg+gjg24my/KnastWFK86SzgVzVA
7hTuG27EHobWC6PMD9OSsVpg47pktaOA3KQawFiA1/XUL81PerKeS3OCd/MozB9c2FtyC6dgHsxI
uCDoVeAFBmteHeIYLCG5YcRnuoN57YsRdVdOelieuE8HzPBHofnPVf/XL8BlLWFYBMkXjpdNMJ5g
PHmcDorSQ4dsM9luzuIRiAqxQu+/y/slB7rcu467ewf91sZZgp5dBWCUTJhoJmLa4TpMkAbCkGBh
Fu705/Yhfc6YW3kReOMZwj4oye7TJqH8k2RsmgU1zJTopnQnLAUXG5FN1qyF+91QzdBIcISjmhRD
t9VNz2w4Ud/+IiinylQMcyjtIGU+hCB6gXaZQRDvgK2bRS+5kr0w4oYuCOmHQvNrPeZtWnV7y2av
5c6fjC/m0AsqV5Ln0ddcKBGDEZAxPgZ9bbUC/irMn0jGKLTlB2/i6IC7DE0GLAY9eJY/kmPGeQ42
QJFqbKCel+/ar8ZeHQ0CAM0rPjTZZmKg9Fkj9QArF47UYdPBOgzEFveylkRHXyYMsd9yCRSm4wuD
UmBQVT3deh5p79+vhLlLNx7HXcL5iEMlwTkRyAanwAfj9UTA5/eCZf8jkur2FC7oFaMfFjz7j1zz
f49TWhcm4y1zgK6JwRQrLJfBkz4Z77np0uZcwvjnvArqsSVEIxbr2bUSm3LrmWJRlHTdgZ6LPgez
xjFxLsDtpXNWPz3TwY3p6jfdFkB2/8MY1RY37VZQfL0cpfNmRGugCPvFjRRPHxrCfVQOMcLytNPO
4nDeq08k+ejGnu7Whwa+XgPR+jvaNuoXrX57yx3txF7ZK0NJg/rCFHV7TOv9g0/8tsI28OiAen3s
IbuIyIKmRhToP3hV3QEJk2vrXyt+hpOBkWJlO5jZwurvdxKAFDlu5VrYtZW/HOpdCvTm7+RC8Gy0
FZUu+NZAEtdNKzyKDbahnSbxvXmYSfN4PTP+RuthSyLshSRQMIinZVM3Fe9r6gEfJvNsiehxNbB2
hUfO61+r0/+2CelTJtu59hDwB1/Y3naoIzKGe73QjCXl4p/XQIo3PdGJaVJ318Hp/HL95LXVNv8d
7PFHlclE+vfRGsSXzgs2AgsDV2uk81vOYhrkDxpJ7riJ6wZp9cwBjr8Bcty+rw/H1rOq9Pb9TWa5
xDswcpfEttnymhhzrz9s0cWjAnViZYSi37995rJi7J+bN+VyPYCU7Le4hAtyRsbr+v0aE3FzIvm9
vg6MUUypypleKk7rd1B55GJwkd0vua19kU6janj+4w4WdLcU8+8p8e9IxEAFP1omJmDmm8WqaenD
5wLDUzs23d69qMoyZx+LQ/UYZ1i4o5yTJ1YjChUSI+AIibPlnBsLW/JxsQdW5f8s2UjV45c/q+5o
kCxpWCJwVdhMtMXVgXFvihto1SpylU730ak+F1wEc9CI4PxdXS49xe6dv7SBPjulHdik44OpmqAN
gHuf/TET3nr9xDmiZrOmg3oqK0m4SUOg/MIoY4OqyqW/F3tBw91ZjjtUYjqOvy6vpT1oooBBck6c
ffbkNskpYsNnAxqeBQImW5VkWwsJ5fYJFw0Scnr1WgcjL+OtghLbydYtATUfqVzE7euPUF/4NRWn
4nglusZSoGoRsp4nFl6vXYlKjA/1uC8QSMW1rq5vqazEK66d76x2kkytV3CiqLcR4xOmIVFKYXoE
W2PH8C2rfFs0qRRR7VcdUVlehb6tqXDPNyYV+PskJB4RlCMCPvWh/QAUdmVbMUKuHNGmw7qQ7ZFr
nDMM4RoBc3MP++uOjBhEPIlJq5iin7xv6keGgzD5GFHj5e9k59AvB/cUaR98CgsLG6WE1DkW0ZZn
FRBH/lbeTFXRmOKg4vGFCHhmcHPlBIqDEDO6VT4u7FgKamhC2jnpyvQ/ssCsNkke44HQMXFX3sv6
Na2IpNcqRw9aftVKjff6L/qGrbDLhms3A2n0TJdGv/3b5aOYPKn1xcc7akipWkUNMno6ujG7H8Lt
pw8U2J5Z8NljGLPU79jqwMsTZAvok7ImnkAZdiRbaMAEehFb/lRmqafsZLBUzJMq253kmeXWTjNh
zoOGJFw1MTI1TS4lFUg2DSDgFXq2SsaILU7Ihnm5x0oaTLKs3QpTiyQ1e4Gm0NkIvGtygiPjJQRn
4vABQurFh+g3c1TW99/2bQg2Pu1qYZVyAnb4eDPSnR6OQguip8a9+g2w3cMbIKRA71NtNsWDmDFg
0C5yK4U8fq8jLf2azkyOMp9PBl8baBwOXgC72LS7JyQ97PzLG6t828XeMEIUOR7Aj8xSvVI7zWVU
TcmxjW3AwEF2mewY4wQ7zowyLech//BsqjLsMByYwkH7GLWAQaMM2ZhphRymrGpdAd6AeMULBMW+
s9ubig5u1f805wDDqEmf9I/iagweBvL/1tZFskw7JgZ0VTomQcZgy2Lnb4OBeLBfVdVz1vpwISFx
W6WOP2thgvdrEJrtKTrttnpd577TgacungiT9EQfYS5Ww1zfkysiJK0iRji1OE6dPY6BSKqMu2XI
ZLeWlfOdLgRmyPfRHQAwXQeSN83bI55aDfXgh3U4GXF6P8+eE9NN4slJDIl+9O0TIF/veK2Tp4hd
hfV9gOTpmamb91azd3KcQLEL4FgVukmrQdjmO87q0EoLejV8HBFys032wxl+EAvfo/ghnqQ34eHF
ua8iTRARtLoqdC1LSegDQBrRfYk1s+B6qTr/6GWDr34gfrHyWNoxSRHn7Cpdyi+05YHpnB7sgtq2
kSwAI4N2XVu9cbQ4dIMjNB/Ris/pdZePX1rfrB06oI8V21XaaqT9ubv7TlSjnzy9Dx1D6amkawMb
XHBZOIy0vKR+XATqXLo7A8xj3H+OYaNVwi7OuFSfrt/QT0vdwwd4jkzGeyAdPYUkOVgC5KS0NQoD
hyORRsv6fnQX33Gv8bA2PT9o2cen1fHeyuaI4yecxlI3uAhhYjuTubf2n3hG2hW2VFgyEiFcaJVH
7rvng40uUGzwep4TAfoo3S6Vq123MW7RnyDwGLpttbRZY5P2UfksdpxwQPxON9AOZ8N7LpnioDF1
Bml/1GNxr9apLkUqxzyDHfxNhIGvDkTeuEPChT4awekGEeNX7aqTkeurQeUHt4NX3rf6uvnGtGgB
cHeNYHJkuRt9EaiEIAZD3Lma2JU3NdXIWxtOdpgRmktInfmvmvq28c8GzsT2v4go2I2sOfSU3XxK
o6UUv4tbyn8yfBpwH7YLydhLtunsA1T0jE8lAH/umaUe7FZHunCss2wkpIwaYLXDtyHTVLYP10jL
8EO0cnXHZhxqp/qS6H+w3l0UpSfITBziZ+UbtL9Qrjc1hv3pT9d3pdJFkBUJmgK+BRzVU8HR9iq+
H8QOOeEqkbdM+3lkA2o2vOVOd/aHKUh4XBXy/E7HUYUhASMSdx5zjr9Jtzb7fUCv3tfytGxN9M2u
P/0hjW5Iu8aCA+HRckxOeaC71uepSiqq2inTCTAcm/HUqgkQXPWB4tOVB68wnadPCx029DMx0IW0
c+quoX2BRngTAN7lOQotJH9zFEza2KJVxUkkC7j7ZOyFodPFfHxr543G/8mw6Vm7Fadbm7xhuBZv
xJnbaj3SJjH2lIKMIi2ZvhDtqHzr51k0cRnhmXcmc8xqACRatWjB4w+F7JTgbvnDbyuPO1X/uhRA
8UIIqCGJy/vv7zVq2myAuBNuO8HuYmUwLXycyVWO0UKYJYe9q+axVsU9+whYqFhCoi0E5gAP8i73
swnKPr1fKfNZPwgbVJQSh0w8msp4MwGBFbvXuEvpIOxqkwIS9c/nmJdQ0R1O02JwfKq1y4O3iue2
W+H+ufSwWTNJltn7jv8q1td+JTNlGYkvjIV3/Y9jZ9iSJQxhEhAMWFC176R3dT3lsxb6+1cq9mFk
ovtI+43n3AKIVaO9Rh/PXW1iCAZYDOrm8InajsF+PV+nAF5vZo4uxqfAlN9RryNEVDFtudyM7rZy
RKSar+RZHvT3AvZCgywjY3sEpvUKLe7Ld/pXi+Aibu+7i2vBmnHVuHGegJ1dhzpqUceMzSMSMvxl
aFdDkA94Cu/kWnxsIBRrfKtOeJaAXhwt/EE5eLFH7V10UMOWF2j5pIcVGDXerU95i2HZfdNbgLws
L63HJ1t8PknKS1WOjoCU3Mxm0/RlxkmqZVhnRCd27wjmo7VaPxzHoIuwaDtpIujr7F92PLxwCuuL
NGm9PnA6GDaoiydigsC2r1XFJ0Fsy7k9tJo3+k99QuhbJyF050CgNhIhJRZR8U00fRCWGypt0XtK
VqexiKcBOrw/0z/v85CQLE7XgNllAjI1C6YX2edcvfOGelzo0l1jvwrHYtGo7LjQ8VuhAysZXYce
2rTtYxEVG/CAyNvcjuU5ZmiEQ6eEFkDUHr6MH7Dt4NWTaqhDgXv3SPY5A5JeqNFBo53ZjBeoaVrW
BdhW4vLWfO8VwdUHZCYTCEIuCCJ9zxWnJnbUPfk0gkGg0o9uaClJTBVXRmkDujodXEAFkJo8fGzH
YrcpoB692fJOLapsDbvjoXNBKYEMalD901Mt1wfburfyxcDDy15QKRIw/drEdfG0v3KdXUaGq9eo
I2rrBeqQNZV/57FDsNt+L/5Vt304DGultrpnhw62RpfT1oNdZODWWEBMBrProqnBUvom/RXM2N3Z
tfhWPiDmCDUxiHOV3Yt0BwF82JGR3/KjySWejfVju91oLQBff7DqgUiqh/W4sOO7MoXy4EOsbRMB
w3Y5M32tIwIQ8qRX6H4vrzsERVkM+cDKWbzuM8jG617M3smV7HL970Zw9BBKzrjZkQxDEMrfVO7Q
j6imVjmVnRFQ+mg5wUD3tdv7NkSgOc1jYOf1SnBago1xjaQj6xiCYIFh/EYKd7Cb5AVHLsyKOU/J
BjGEUPYz1lYipKJb42nW00GA0xBrJn1S+bJu1RhoVGmgh6MNIDAYBWBdy5uIjTIRdI4ic4rL3Kh3
IYXW7TP0CvJsrprr6ryMZm60Df6EufKygKvq9aQDktUo16elLCKozpBvlT+pS2oh4+UlkrklRVBs
V9s5AUUJRGnvU0XVLm+KkHWcasMQauOFiGn8EdD42FtiJNVaEo/GzssylMMHXkZdWMTvvnoTDNQp
IPe6PP33h2yVtnrB0CCZA9ZlB165HVTlxvYTeomow7j7wWcliVTh9EZaSwKVVVpGsTBtnDFOBZo9
5j+if/9nT3fa+SFf1UfDfJY/ZS1T0Z1DAn6fDN8eBcQwl2ltBPn5iTNZ4giR3Dkm8UcS/3cB9M/0
BDOY3EA6nEHCoKM9rvqY0CUXpaq02HKtaeePWD8KrsXkKtEtnLncESkiazEFHrT1/WXu7aww2orC
83+riJy4S4S4eJlx5Yrdz8y2I52tFTLtKgTb0vClpfOOYzgYWl7FW5DRy8V49FTxcP6/3SwT2CMN
jMl1VX4JUTMXKhvvCXC8FgMU35ogvnLeZQ7wgPvOVr1A0G68qqkFFvaoHInhhN0bHaGnvtEKWssC
7i05Ykd7jqyyUSn5y4ogzWHbKFRnGGfU4zabhU+54qYzFRVUNz0IqeoWiP2n3ZU7Hzq11lEFqAxk
yCRyzZ6YKxBmnx6xRD1uMk0VHzv55JnWPkM2Mbtqp/NjNEV0+3G6XK7czw6m+jXgy87/+DtxYPXo
40xRgSE3a5nUupBNBHPdo5NpCue6em3cDWUs0dFGT5q1oNYAVzjqCxmlSin3I8wyxRcUp9DW84Cm
D6Vr4MEM6tVGdl8ni1p8b+wSJjUlIcjFP8+76Tlg2PUkDm138IM6aTauPvS16mNyl4JoMooNbPbw
/VSGL61ylaS3Gn0hlbkxV2QH0NyCf4HIjbHmOdS8atFyXebZlIPYSr3RCwcDkYevF8btT+xSVkQq
RZvLbaNvIidKRWLBc2l3YvQJjaeZH5+dnpq0Y+wHaxu7R/zofVLWkvIzlWqnrgJEHuZfoF6mxf56
Zm6/P3wAqngedufKPY58kw0/1c/ZYAsyEKqdw6kFlEZ42T418ctmS555Eue3qG2qZuqBrloFoYhY
1FLxdxv9SkNxrofGHb+kcNt9+q3OAAgOZIxaBOyY2yIa/1xmYtQEOlTBasAXRmtrVwwmMs6ZSoLv
KukfxzWYu7SmB95gb/0phppgLZ2l2etsBGr2oDQV2vN9mmLYhjCUmSjWqsfoEeKQ1vrfK/t79QvC
K4sXhqK93vItNHwVXmXdz8LCjlJhBdB6DijiRWjL67uMveadiTPsSM/1ye/GapjarBpkqT/TCd7V
oWsIWCAqNMcpR2mytEDHzQO3WZ+ZCKQP/cl5cRSrpZAlYnKxfj2R03IBbXn6apRhq0jgoEOEIrFE
zY6kUinjukNkxOVVb3X+YZLMbsFJ1ofyEdmOUNDNHN35tDngqBI4yM6uig5rt1kBuk7asWqB0MAs
Na8N1xNCPiph7IfUWAThYMdttXH6xv/VOftEi3sMdhfqIhXl2pPcGDQYpX8TXQuUW0bAwaJPANL2
BKxUAo7f1zfrvRPN9P8WuF9yMVhNpSlaNKHwygBht9eoJ0xw2WrXqX+pdpnrnASKFmQK6qDIAa2I
PqkB1dyiAKNaaNMFGwxTcSUC8nM97SsEtT4/YfHw8vCgWQr7OBUxwr9aPKPSsTjbXIqhcjZpdtk+
SFbbfddd2SHoebXG/pqJFcmRZMQffpBSRKMbPjo5iWDq0cdCopJJ1olyDPJawrgpDEzPggS4SLyj
sd2CVMyNNckfGENBsDftl1CCfMc42PdR7bbuUoHrmrdg9E0jltMMqvJ/iGAz1bDqzSwE8w9cUQLi
8edeh8e8iExl+Zjip0EJyJ0JA4q6Ez8yvGZRv8Y3PFJmwOuFczxGEbKBtX30AOdcFOs2epCuzc6j
Kr4Yo9RlTKmRAhnlznxcm4Y3FKY5lLpP6EMkq/R1TAIEwuGWYTr2XuYThWdhAddmNhFj1blJ9USu
TfsQSBicyBnapwOXJTmAt2r3NucFVMGe8RbBKSMv4E/DRl3t6kIJkeXsYZEhwF09KL+MI+Eu5x+/
MDwZc5tq1SaGiZg53rrC/Vo9DL+AuD7IJZhku56nXvwaNawxlMaH1wDfBOF8usE9TKFa4P7GJh24
FOJgBbBMbjF3bgs1UXzRj5y2r2+pbFOWeTWoi0ZCxOh8qj5DdXBnHpmiuaogvPjUq2kvRhRyqivf
IPrWqGCiP3D7bUO/WfIgSLCDpqVqi4H9VHAEezse7dNgiXoa83lWRrux1is+Fu0eDkPAGrURUPMm
SiNs1OGfCQqSGwOOc1HX/Auz9lw4lucXXIZ99lELK1Y5SseGVPO6OimV9kxpKUptWooWkypGqg0Z
97AWn46MztVn3l4vhXjDkJlAU02vLarRFK79NwsggmRWItfBLS9F+k5e5w3tMifBze3orsZHez/1
mxYldDqRJWKvjFgygwUTIANlL4yxRaBt/qQqyHYRthThVh+Ps30umDDKBwI21wH42SPj2UFB2iuB
W0oWEwmTtbCJpFRfePl95L9tpD6NgCWWC4l+yk5kN4gf/JNl5FNO0QvTyncutFyVy6NahXuJnvIm
jMX1P5yPj8uURNA1KFzid2aa84BQzA39ohXF/Iv+Fm9TEI9aGUjubEWgn9JvjfByl0ktXSXJzgFG
u0pstP6sraVIa6ZCVNWQolvYOAaSjfhxLE/5bqlHlO83Dn3t90GMw+ZNTu7f3p/rH0Cwbk6dPDPm
03zdwmdkjsdp7tftb2gDfyE0FHmsZpfaURC5BXRTz4RpEOXQqPoUd4dsSaLFGhxGXURxpFz+Jzcj
c4ahnhlVO8AZ2rMEnsumkCyOTtTOMNoCarzdRwxu3/hb95hb6gkigOz59F9ASuMrA0mc9KrcwANU
UKSbkLu8deTe4nk4NemMoPmnD3CBEIay19HFBd+o+GYkWrdJyewSgB5FbllFlnRf4REwxfBOpNO7
iLHt+ykN4uJbrYapsofSR6o3BO/sKGpt8D0qGgROWejxBVUMDPYkhCLi3kDC8WZpRDs1uwuxXvLU
EUe7Rtl3ELAumtYLAk9oZPodtkCwDBNbOwYitai0f2jK2XvE946Wjo+UeE9M6nULyk6BOiMR06mn
mQU+J9ANsPSPp/z7/BLe+qmSDtnDbGTfd9OMnxeFzbxzVqO04oIU6n8PzG5+BeE13xIG3wCbVTvV
316h5r3HuEWTpObRPVsw9vDugtOXwKkOjsLbpgI6UL21eq5azT7MBb8SLUwJuy6CfFjPqzymf3D4
+Ht1+Vb1q7uw/5qPvj2uV2wCBtov1ox1QrP41bluJWTo/e8K8SwQxM2vWuFRiNmAeitatSreDOQ4
r49rVhm6THc1NKW/34c1khpYqXVpEBxbxZaENg27EDGISwKYbE0O/gi2swPfI+EiEBrxnu8GE75k
aBq2/zECC8HOFfazD57uPRZ/+RVkDd/PUbSNdEeorIHtmF4JfAf85OgaL3mKd7bzA00E7oDg+0IH
YQ+4kE5VExzV+QXXeXQhzX3a8Ov/FjdYRJCoycW8/C55ffml3+VXLYDYhxDP23V3+L00ftu8lEgU
iQJDhhl0ZhlHSb6wsAeiZwZdyP61Ho3TGj5brLLqS8WkY+VxANHgICBBfYl3oIy0e/75UB9VXveu
QuHA+4Ks8wAw7G6HcKB0S2U7e6MlgWF0lFrLJN43QlpZJHnkfMl99lTfhv7hNILZXiMwnOsiXY+8
HMx/TrfuHFR5dIFGI9PLbTsPEjthQvjCRo46BrxQmfI0V4Z4xb7klVcJrpXj3iW4mvE3EwS8jf26
QEYxYh+JoSzQJdyQnh98ACQkS7grtRmMI9rO16p9AG1wZHJo6dU+f/1zTw1TRFdwqe50dTJuEOPh
bbZn1Q+gRM2RF+bS9aZdl4E9UacgmWSLxir+FvKQXLNws79Xz+R/6FSJeSIVGdcK0voRhgJX0bV4
qO3kmmqB1a88YlvF+oS+bJZKky/f9I7MfJ+E8iFY2lQ7G1ILvgFwAh/UX9YQbCHedRvIOlDGEUzv
/yYntyPtel31zSNEMTN/N76S2DFMQA6S87ibhg3mHuneiGFoPfGUDE6H4n1AFwzLYpVYpG4zdvza
41gH/OIz5c4uiPufUDc5ChfEcIkOLOnIrrKS3pGehJ1cAG4b7jukYpuiKs6gdFcTAZusWr3uoRfT
udnGg25Gp25oKiI3X2BdykOC4g3Z6q7/yUyBNriyj1pGjg3X0UMlwwC1H3ffbEtlw3g6mX567adu
Wl54pYJuE3N+F+DzKQTOoZZkNAqGpP+qMlEscNSQo/5C/YATeICtMmVc5T+7pE/FHCY/CcjGDsLU
VqkHwN1fAquQI6lFPxxIin/UZqKGTCMrrqK2/p/u/Ju/Ef1pA3hCgXtc5Fh8XhmyWe/12rFQ0Ejx
yb4bduafeQ8Pq4BFAyhk5AZSoet9gKdTLmt53gow3Leg/ZHF2CRRrZzqGNm0zbm/70PXe5dgCw+Y
5YiIBQLcO8Tuv/bcofi+Cvar4rHma0M2I2PpwglMJ43AoCABZmWH+QLyLalJqroysRpUs/o6yVJb
TfbWTIvjPjSPEimb6tsjcIyeN0w1pL4B2oXDtVVK3cMMxjMybCajEAm7bG6GBOPK8noh4fGroWW8
6HXO5s6LfN/jZuwjtuE5SAlHtamVgYHBVnCN9F5dWj6ldgdEHxlVPpGjqWIrOlXvG7zAoHIOri1Z
TCCj/FNhHmZvYpDjwlvmlqVQhKTMijMhGDqp7gOKW3/Y25l06t+I4LLTUhZGOLNWb5SGb12zB4l7
trSyhhquAaZKz/FZjhic1qOLMbzkn7hmDR0HAzCYbDaWdL/10ObEAH0oB4iEt89MhCQEKdydbsYr
WTBrN9SPxjm2yWHqiUNEKq3n00A9DobDwkxUlYl7LTc1LKWDYPV5Op89sYMHUgqqMMSQJMEUJS6M
1CGLYHjwhjKRgFlAGdwUrK4Z1q6LVd0WbjEGFCpNbyP+sCGjdJywWuZfyMscB1rjcrEbrOrjFcBT
JlDTJiI/R5Uk0ESwIuDmUc6dZMFPejQezAr+zcXiBvkdkfbCqWRCWX6MfqnWkL6tZD7SlBaRa+31
eKVOh3DysGCZ+5OSM3No6wegyyafHfsgtxk4f02CF61OuqcoTeQnt9aBPwMpqORZQ1H+rg1HulBN
6OQCnIp9wJQxZ+4IbjdcZ7aBpxbowZMmsH1mq2upTvXNoAQW2FyUQwwQwQZOM9c5UQjgn00HY5PI
uRO0grKya5nlj9iYVkxPjbiBMIQ5C8PLu/A5OsXnsiFNZZtMFmiscyk9HAvD002iVH9hlp4NijSj
q9i5IC+SZ/4TUEIZDEjmhuhokN0/7r6O9ziquLhf4K24XGHLKIWAeFamVk1fPbHDnORHQjf+kc0s
Ldea3U3EYOGBXEwcxV6U8Jv50Z1pBBi6ZYVnYmG3kkyHxoB1q04OP+qpViYzCkx91lvyHpS5v6ly
f+DAD27bvrYV9K0GPtYxNDkR3HKNbVRj4AVLQWxI2NbjntJLV7svFIinYdQ2Kllk1n4lb4TRxVm4
2zlgoNPP7N/Z5lAavg2jWHgT88TqO/7cqjDgRI1xods8/TWRaAdg8o9NKYwGmHqka1eg94/GY1Ts
k5C312EY2kfqXIPF/C+4DarImb2Ajw1hTJ3ByaFS6nsrvz4XpdyqgWUfvu2AHEMOsW5scDNkzVsh
Z9Y4kXonhnNh8M8mwZSPENCPz0kkt2nlubY9czpZ5Nt+5aMFwfZaErKNCLVeXJIwPRVoyTeg9tT8
EK2yKNxMgoWaaPxGncOAhF7Zj407xlwWeIGr0SjnnN5kxqq4W++O+sCn/OMQz6747XHcEaKY61Gb
g/GvCRN44m0HmIW6EUfJn8cKqjnz3eoLOQUBmngUV2mBFfhfd5c9oc2UCv0RZ04hr1PopGT7mvl4
DF+uMXtOecOuVcD8JOtgjciPXwOJbIbA978HbMgxkpjjZZ23askmnoZ14DEW/EPauabh4SG3qt9S
BSIoRPJtI02dKlzTpLdbM/hpudH5+YRTGSNfPKJVuDoHEmNOyzehVHX/WxKUjVYP2G8J5csbe1fV
AwmrOvm1yVU5v7UlSFX4pg9LkRoKksAtPrKx4Xf/7OcGl4LZcohgbmarffHvQOGBpvA+a6umHTic
eIz6WB0JYl56LgDVsRwaiHEOhW05XosaT3vwcELwl/Gqg78LSNd7kVXSrLThpwClNNyxXgE4KBfj
/j52PxkrIzVh3D9l3Rm9DZCwHyHsIlRvOwx53dXZdh8K//D9JMc3q3s+fXEnpbPEPuBDYS90wojE
rjqR2pPFc0pZTBRQNRtXWyo0dUa2qcqymGarOlOgdtc8HQN3dylmC9+UrPV0YqhAb+g0FoM9UMaW
YLbvFQyfngsx7BeKv6Hgu7U8924p8JFir+0SRHAzW3bRQYDfb7deLvbUguKNOfE6WktkCawH/Cb6
KH+eIa7/JpAda1QiWcCPCRMwZsAcXrFdLWnG2PsLbkbTJRKUTqjOcNGvKrsXdD9E8muvf+HOrZni
jBZPauXi/qVo4S5GJDdakDTaakONExgcnck8veLJYwYX2Q4HIPKe5kQrwuBIYIXjyME2ZY5liZ/u
eNJZlqDKYM8sdp0EiH05o4cwbg1VRM8EPCBq14eA6LKaDRQqHy5lBlf6bUq5hP0tL/ddUOA2Vh7X
g4NliEx9Chs2TVxEPzXB6sC7VagnRGOe+qFA7wvCXje1Ft6CHJEYHN22GJlR9SkTltXkdbEY5vUc
787QIPLqPcHen6Ah6f+4wYfYK5y9Sw0QNdybZw4mmwFPKmeM2BykJHkPWYUoMiDk0ii3hbYYdv9r
A+1x5jYVMwMNdrxETiuTrmBjMT6qsZ0qDi936d4Rvs5EfZY4aZ26O6U42BInZ4vBAo6BJwBx04qy
ECwzMC2/fFbe0LhQrZTOk/wnVCvPuuSRlB8K6x6gV8fcof4WNQsRcuCPotBCcX7XDAWEYeL+h57j
rrg7zu1HGtz4kPf2SR4APUaqDbje++CT2PHhajuiC7641sHmXkKFU83q/dy5t+hAiXh/qaUWDpT4
/j6+CuZSUShczpXMnhsGFx6VRI4SXfFaIMirHGKG4HUDbwLdhkQqKiAalBSvsIC+tpKCMM297NGx
xz589FCDTG1Z6hEb1H6fotrNIeuXaOWvbw9mXR5eaQrUXPzKXyWw3M0MMHeHQJ8wU3/Dhm9ybooe
CkW0LKwyPjAUWok7rxNk8GxB6OdM74vaQHi9wYL98IAcvaecMwdjEXXZbZOXA9pSIjJOq66kPUZc
n62eL/hSFODNs/D9DlyrkpEGdgH2PALU+GTEexVqCsp8Y9EXoFFHTj8JtHEc8JOP/AmZ+X5JNGeW
Jpu/X7LAqDF0LBYQZxvwkeRxF4OMaVJBRkMgY4P+C47WIFyeWK2n54XWdoeHQqx2doKb3F8V32VZ
aAukjPi1uIhSUOgEe++MKlVAeKqY69lUgzRQj4iC2VaiZRjXaK4SiNnjporHcLfF3LsNeHyFb4RU
8spGjA5q5xc9YFeOX3GQuXfRccO4OSP+mI61T2t23Zd58qNiSD7hUvUDx+DRKBVTp779L/G2ojJj
5USz3l0ZhZHnUvprtWjrt1tuelg17dRLQoVJUu5CMzei0o8zR9XEGj88dQf81Cj3TAFhHBsOLC6E
5sTaXqvVJJKX0ElsuYjlZKERSBNbvWxYDxmrFV3LBR++kpKGtRBs3J0lIMTPWYVB+eT4lkNoOXyD
ckOqtJBGA9rGSKJV1Y0AGgngr0zuPuxHgLx/COJLbd+HRr1wEu5IrJK7RkVtigHw5dj7iEwKHY+U
nPEmLk3B4r9KKfJo7WLbyJosF+MME34fs7LlgJNPydugcW2+H3Nky8zgLPWSYZFdf2Gw29P99s7s
+QmDQFJTU1h1CbyOl3FpP3fSo6oO5lo/x3LtwE/VPll0ZCB0KJvsXIyT3AIFamJ6sL2vDn7rhVG2
PxFJ6fygVhhKEmCyAE/39g2BsQjzxBsfkxIUp/sfW3W1mm+l+VzwWM+gjJR16P7ktLIxdaZn8Efq
xuBR+neQ+P8RBXilLD6ikXPodpYpUnm6Kl9qFzBFe5gYtblRG6A13R8UeZFd5WuWYNDqso/kfaUA
mi2ThE3glSdWvDOUKH9PJ7sbGDXLliOK9MmQUjJ6F1cN1N++5Mc/uyrmfKbFKJzMPVZzHHwFgL24
Ce7ViTegGlq4HKJE2RXgY+1kwYdp6gLugbTyuT/y88fF+UkcZPmGtqGe5wmv3LsVP/u04+9n9jhM
rw0dS3UmnsWJE/ZKotv991qdgkPsgboJbU9WnpVgDRxGplHAfH81VUlLgVnh9IRVTokmJNRc6gbV
EyKe6NmqCqxgwm/AsOl/bDBkJDHx/E1WMA7F4i7pJhRnFtARwVycXkfc9zvdgKj6OYXv7CDkA2E/
fobTaRxOEX8Qf9PqFDcMfkVGxNr9mIo9lgT7yeDO1VU+gTlsSxp4aBAzPGf3Dv0WFG7E6uHYQtws
Ntlg+skT/PsUqK6MeAKsAqdyaEVpydAMM+w+2CQvemHrTOKxNJE+qlqWq+LIV5HytMruDs7vW6Ly
x5Nupk4Pys+JwYWqMAzM+tcKfYg4ObfodblwAV1dSB75+I9GIkMEDJ40JYzjfz3TWgLrACwAJupX
M2ArlnBm7UiYSxnObMvIFq3kd4Sz73LjTLZZPby+c8KDVG4vIFrmhAf1x3H4VPkdhVi/x7l2tMZx
P5US76hDm3/V56eVtnLAIvM3mFV1Lh28gpkiMqZCySfC9bnzOQuXs7ESSrvphPCi/OpSgmuNOIwP
ypB55FCdK32ABeOMVZBvm+qEkQq9tr8hMH6ISZKrpEE+dSKtZP1HHnEF7tk9jTWh18tjG+wNkkWJ
b/8nflIJQHjmP0tZ28Bxmog4WXMOJ90raOJl/8RZI/w+kCIFC8w/zd+jMuaW0zcPpDcEYUESQhM1
/MbcLyUu6td3tKH5kGqSHDVQXIT1NcYTvRVLsbPXx2EZPFiIqrbTAQ8EuLQ27gjVDX8cIz5a1xa8
mtJGdjB234K0UCVGwoYzhRdp2hGuEQed7PT8OUwVKzowHhF3gembl6KJutPPQOS+LL5U08yb1uYW
Kxloqd/vWa6AWo60bj3CeOSTpWXZkBO+4r1C4bvvGpfoDy+Uwz3mt29Htn3OfILOGi4iTviMQgDV
aN01Xl8f7m78aHVe1xiKFV6MQ0GBUvSTgf3sstel2pdCtKtM1eu/sJwUBlB8HbJPNvNa+dBLBiCV
7Zh9Q0P4JT24Z401CxLCsJCQo2tZQE+RPRe4Ku8PrxfCeiiStJ/iV8rhb+rdX5I8tWJv2pI+Q2Pe
8z3YT6pTauTMaXGCKNuJeDVGDlVsKvX/cnCVSxUY8/d6vSxf2DOOiJmp7Ln99SimN1W+4ThXREv8
UJv+PVNRZy0OaxqQDfclVm814i3HuXmZqDVpZ754ZrlESOoNOkZj+7xRIo308InP5NOR0112FUAn
nAZfYDSD5Ovws/Npj7Xiw0ZTwqizjPzkMhNjvX6G5M6Sg6cx9l1iParxYY8myCkU5koqSXHcPUBc
XmSOpxMv1gCDqCGa50CkKq7+ZMXdwzICAW78s5NBmYSIPlM+T1CHnXGq+Uu2WIiZR9owxZRgL6gm
PeCKWULqpBxFRUU+mXEoNjfuWj78zVEqFTiQ79PDLT+xG63y27YUWjUQL4GrmuAvMvDNQO235eaw
JppdtFCpa4qrDSwHZ2VCvtci03GR9cbcqz0SNkokC80lvjoKfCmwz7VneKDFEfRlc0C7ctdqn6Oz
9ezETsQxz+709tm21H8W3/AdK4Dxh7+gTvva9lPGRM/CgQs2I1BDqOCvBUg5h04sHhwNti10vsJe
NUUIMNKVXN3theXRx52jrkre89oEfQOoOXMo242GDGtC1jNApYHj7t3wlq89+iXWwEZGDfQrGfT9
93NbMLaB2Rn4juqDgInmp/yWsbQ3uD7HZ5Z8DSDGy/td6MAAmBXVxOc8C8TxU77a8BYqWph1sWXd
XAbPATbl+ua6bhUPS38ttbONMkEo1BldfwinVy54jZ3q+zM1YhBw1WQYj+qcuHu9J/SyOMIV2X3U
pqoXqNaN+gMIFljNsyPuAgJn3rAReCcPH6GWNYVnGN+BJU+VsMOHJHNM7SPNPqQFavU9dAvzjjhd
h4Z3oaOnmkPfl91ll6k5h9Sbi+AqYs2iFBKD1dc3QpKiATjovNP8HO+/VKcztGZDNUgmfu0x/AvG
00H6meFylbGF6gd6DE3rh5nDE5cpvD9H66kIvXF188pllXyhix6jmf3ygRHfOSJwpeplIjfOVVtQ
Dr9nX6SBt/9Ml9LwKlRVg2T8Z6rsl29pkzrnVMv+40ZrbojKEAFXvZbZdaRzu3z7e9QdC9WZ8YGq
zWTOwIwP/A38rbUGTBXzxQJCOj2ssYwJ2//zyfbJqBoQpJJuuP1itEntf42SY7G0iZr9E5FxyCV9
IMGAIdMgid3JqpU61GDHTDrmS1mrc/rfZH8YH083DTAV44Fb0YTbrTEiqtmFpWCbC1VE2BkqGDaE
viYE3dF1XlQVW+UiWXbIXpaNr+q3a85yxVrttrbnLJH27bhtav/J8qpsgs19XRuQCURBw0TpYCNF
YP78JS5ck7zY6DxmES8L+dSVtdU2wwNUQZGKqErDJR/8Svmo9sT8dIFes+5/chuE0qoJrgxkOenD
bb/x5QnOYdb6m/rIjFnq63Llhv8g6A3Ll3j9i2tyciqsx+pG/X7Z7dXVIXDkeDy7FbvImXkj+E1a
I+46JKvzef+LE1pfXQahpLWLIbpAMO9XdFutmZsIbpT8XoS7DzZYdBIJE8FzmmBZaGTZGkR3/BO7
cmHGBJgnTHKIWiTWI6DkOS+9bVhrcpeG9J+1rE4qQPPuZi5Kl1rVBYPY+ZMfHE+Tmtvru7Ob58Aj
dexZeo3rgdIOzn+N9jLoMp2YkE7kMKqU2YO65RcgIVWy4Uu9j/QjlwNxPjSotwRnjyTtmTQKNSah
q9vyPJ62r/Ip8gkqD+LdeYihgS7ymYPspuMr7DJKW+qeTUnj7ONUcCtEoIuECOG8G5dFnKu0VCuC
9KMhI4OOwwf+iZ5xg8KXV8kgiONdFmwAfN05LJb3RVayESJw4Tb9TLE6oneFj7RBI91WSHyBo4hd
zbjwLzjKBBvoJQgTaauXpcX5gpHPAWKQqNOJmWo3Jli9zo8lbwou/GDyeEsqu7UrKzuB92F2qXU1
uszWhwAUH4qGx+O7acSRCuyKrPcoV3VHXNYv9ox4YyAjGI6sdmSq1KLsyTBcFFw7YJTDtHytn7DH
lSNcpIIh5Ov9fv5+XsF+7ch/EBx46chzPnhAwIUTzLr4/qCyQLA7cbMOqBXfMSSXZKRVZWtd4SXA
rkorjNfTXk4QZy74IktIGr5kugiTeH0tQgLlN3T/b1rmXEihhLjHKVfZ98erNFTLGN7euUfvyQJM
AHkRrMnajcOT5BaaxA0G3CAARlqRbz3YDv7AuEshYWG2y/gVTKutEPuJInHR0dcx2ZmfQQIrIIaX
6KZHuW33ozj/J18100kXSFj7ud0sp0NnETN7al0PxjkVTqWi7NSW/XZ04+mVZ7Nn03lwkpft9lw4
Hg5w59pptiuCjUmd0xZCYVLauJgTRmaPNFkFDAO7fmzTt5YDaLZEO519rskIIDxHwn4nBGG9J4+a
+1HyPOmoxrEqEZkzL52aZg4fAKM+dgfvpImKiGVaHSB8U+HeQNHIDuG1z4dkAduljCSUpKFLWfs0
rNcG1102PdSzeGkVRAbfP5kIjykzSw5lSAwCkrlTqR7Yml4vjSPM+NwibMlbbRO9skQSgc5tPeR0
RJgUHVPuR07z1lih2R51S95QD/jRska6zgZ4eKkFq6QDrHotvghB8cGrd+DZSRHkQq/5OAxXVHb4
uG/fitKwyOkVEUQ8IyQ0flAzxspx9sv9dDQqlJaTfkScZsLL6Sh73Q5l3msHid2JyfyHKR6oPm2K
cCxW9mObPJ+IYQ6YWklq0Ep2bdX75eFIyMjHKIssuISewF6EmD865joV9Ll9Tx30ZS2HF0uVqPi8
upd36YqcO6jFWXW/UdSrrpWYM38bpv+2/LUp7ukJ/fkWvA26WD/LQxrmLi0DsgGLemb0e4nrJXLu
BoAUxRRGaK6derwAN2wBUlDq8eBA1IE5+M2dWGS9gwIKuws5tlsKOM4InmGfcU15icWEmUViNHAM
WjjWxI64Oj0gAigoe6lfrIb09Lj5vReWYw5zkUXGuneheyHeNIkpsacB8s4SZra9jwZTVPGW35cV
XtUd4G+P2Q/nnwkL8SEqzm7LyMR8PnY2/EOqolmBfKgpi23mvgl2NSxw9k4aEmNcOaxUJnK/UYu1
kic0W7gaOmKpaaepV/HewlvIZKBWPIJzYrxCPNk3sRvtP1D+7DE3ijF6kb7FKu1QWZvu44oQFfvc
jYHyq+l0KltbKqakjRj2DnSpozWX9XqkBVBbRYYoG+Hn73GyEz7ga667ovaPd55unHuDkRA+l8SX
w2oMGemZc2gRmedIjq+/3rtMAWhyW8Aj06DvwZiDDDHDEae3uU8hOjSxosUMe++ZsiBI2e+Gd2MX
jrL6FIIjTbezu1r0f8kPR8MzLQ/82fdUT4VAwAG6ydeBt12ohbM9yjPkHnOCKkM+KeUbBUMgoCIG
QyySQeNezAyjzd2fPVowfS57HPt0wevLVOcxb8snE/9EY9po/JkijusAB/7komPCjQ8uBiz8FTrd
wlakakD/TYHweUKIQxB1Dt+wutytaUlMfqO7IVcrsMbvVJiTSd+hWUl25IF9NcZo2hUdDoBHDQzR
3QUzTeQ9mhxmi8l8J4cWiKGtRV7kDnrvO1tyOFtX7K/8o+q1vL+XNlOeqIZu9Ai7c17PwJgdS1v7
3CYKGFXMVzBE+V4iLRW/xzBVVTyMT0PjHw9w4Wu3FbmK3h/gdFfE9CJ40nCJHZojX9dZUOzx3gpt
sm3OzUMjuCTGy7OlUaSjtJiPyv4+hqFXXwqx7ORbiMfmA0LOou5OnG9TEBUolWIgeCSqOP4SWlEQ
mMTLoTtHT/IPjSDyp2gtcydg5fyaSzvlGb2SFBbkpfqNPgQW3usq4QL0wTFY3PwXPNwsHRmAVr74
NXkaArISQLLjB1vsUrCEUxz58Dj5/kZVZlg5Mgug0AUwbzr+qkCnNJc6XxXBvTgPUAJFUFV4VGcT
mzMZRMIDk/PfB5cOZnbD/xGULmiumtiwpIlC4tlXkv9ZiUvwZbvmDVlFYxDMhffCrj3j0k/YzJ3Q
aw9s1qsgvz8XsKWdCXc8oZMmk5jLYgxVrCiC9tavFvMCD1xnVMqIsrrZ+9yGr0ZHA2qaa2gTtZBO
X5O1VQ6OA7o160iKv7hkQV+49dOqrDOgt0788rECms5LS3HsQ54SJmFOZLQXTBNYtoEWL181vrCO
3Y0s8iQAibAQrT0v2dVIU8FeoTLIb8iarjrNDhlRM8piLC+o4lbiqBK7liF7dJKOERhc2+HDbqz+
XCghwWu51Im7gdTK7YqsY8HTRoBzT8R7b5n+N8RHHYEwY1Yg5iFLzE20z9E1KYJM8I16BqJ+FghX
aW4CXUExzlgOzUl5R12ByT6BuTpjVm6/onB0yAdKrcbUSkSkEo7rpr0wceqOjzyCW7WpYrq9rzX1
1T+/du1fLaJdk/+GpIr7rs5uTkT8yu3UUsxfO6LjSJ8lWZty4wBu5zjtREXJlCx/hCBw0DE0QqdB
//jlQUMRBfTOGe0Cdj8Kd/Ln7Vl8QWs1Eoqf4R8sZ5vQspBuKaWnI2mEF1+6PvJWps+702+J/Wcb
eKySlYFFrIQ22qNytO64/CNjsskYp9mlTe6cIQ5ztqttFdVdZIv2v/8FO9upYiqfFFnfZ6tm2yYE
xaNg1GSxWObw0qyVstg5/oWxAkLNk/FlNs2p1iyfdpREnrnJLxRpnPh5KCVpoc8kTN/oWLvIypDA
wrUyPhaBHsdpCuajEiKZSeWHpIRNihKh4lxs/2IHo0bLmGZrvxRGLbqPUKtp4XmuXxhFTWjsiC3G
CzGzLpd883MHhGVyUI8nOBb6j2/hELjyENFHTfEm5ayksyWT3lnVUOn9ViSeUpOVAacN1RIbmWdt
/qCu9Zgcg7yjK8845Ox0rfPkoe6qbSqaugG7l2R3pgtgyVuNuVqZ9R6AjOA+bVnWCtAUQ+6cegXu
kXqLd+aYmYDgoXqka97NxJFGbGcv0Rpwc5IUWcCuaaeZUA3X6GK5YWqOTF1dSyUF6fiTNjHvim2a
J5ctzPmFqI0D/K8w4ac9T1gM3xlkDzvfz+YAbamoiY5m3g7XTZMee2aNeIKimAhEj+w6+Pd21tq0
nDf+gbfO7lxCcQTo1Klqmo9UhJvUMgllO6zbYlzJoCUq5TKRf3RbxAzp26lhslJyx9hpDmcfsPQt
BmUfGZ91/j0IFqjCvlTzcdAk1pz1YN0agxB/znAqLKwx586eDEqFlDGiqYVDkQnevW9bLUePqohq
/uQL3Jst+/btXTvfZ/xNLhpT7SVqPXus1Qtl1RfFODKCshE/YBfhv4Mz+Sc/QRGVFdNLgWE7VD+R
ogSGMlRYZh60jsrFjeJoDwqGSIV80WXbig4bLIlO7BJDt1Dio2jqG1XnOGruf9qSnfR5lnzHs69u
xLRrKGqkvShCBQVQCzWW2AFtRf7aaxSW3l3dkyq9ccUpsRoKic9LAGNfUQ+bzaxmhU54oiPFusy7
z94v4ZP47Ma/7XpqfbuBp+m5Kqfc4a40j45AcUX/4CVO+GN4bZSpC0+CfHKgrmaFLR6eTJMzcKya
BaiELNlwKVDTawV4tdQK73IT8W13Nc061AFhiaxIwjt57m7WpDahuxNUfiekELaleOVyHs88gjSR
2Lt95pIWi5JKlG/+QgT3G/o6tnzTuwG/1p6Zha+hA15HiFQJ/hKwrkIx9iNdMv8vtgzLb8n4cHBH
KuF+Na60oKQGh+MdUvzZ5YYjb3H9XKS6ni2PPoOQbQGecgubMIWwvy1sGh4lT4LHkMQQUD2Ltxtr
wG/yzaKmGEAJVc77//WZkDCHvKnKv1yoWEbdAAEWHnGtnbZNOaVkk6kSDWKxxa5MhwIDcbtkuggt
kkbnZOW54KQocHY+ARv1S0NrWHlvaWjUv478QdFjFOUT+1UfrbRZD+0FmzfST/mIsauF+B0No0ni
bT4nbjY9Bce1aga6/zFOta+gSZrE3CVvPAp0AiAf0kzBZQ5Cj2VeFesPUiZxY55nwHjX6unia7R7
y+9DyyWMw3AIyVnhB13P+bdGKW6PwpDXMMbXEVytD/kUMPHm2avT8czpAtcJxZYmo/9usM/VYcDj
f/HAzYnz5P9IlsT8rGUFs+nHWA7KKCgtWoIbYWBIfy6Vj4OBmzujMKuwljC3qYwxKXRKRILDtcjg
Ffphguhv+YWKII5tLIHlig+c+Z3Rz9xMixJGVo4nIHlj40MgmGt0mYIubC+8CuIoPDphqk7zeucP
8q1yTTNWtI6LfxYtqmEB4XatqHm38tokU+txxaYr9IZo5xUw/a9a01NeEyALLxFlHdFH6fEKNQ6T
jlqIIGiNdaql64B6w9Bq2LKxrp3VwkCHqdfHlA8iEzRbkGYsI0jIS2y2BulSM4/tpO8xh1VCZw5y
kn0G17BAUUSpT2MyeXrit2b/WwrEdUQ5WExhhkfhyyzoP+roK9yhaM2f2B5+nJ8VwVRJzOGOc3G7
fPfl+PJQ3EfFX/pLmlE38+XU1DYtgexAiJlG5lkeW0ySO1ZGBn5jIj4frrXtBdWAxpbKefscYY7V
t/gk3fPfOs4Zp/Rt332xbJe1tuPf+rmR/ybJcF8VYpuTtcMjxncdueinJfy64xXDcPp7q/4fRfve
JclZeOPmrFULlQkzhQbznAwctP46VXXoBMO2SbtTvb0xCMEvZ8kbSMYFgVaBOdQp0NfacqbvTCub
Zh81HKPna6/7g2eJBKkgjFaOksSVXY1Pf2Dbkqb8C57tsH9w9tLoaXgFBpRdMh2ieJHEcE6AXLCd
hm4HBmFRL4eFzk8UoOwAkD4JFTjojOasX+2+VtKbxQVNyBI23yL/zc0N14VBB1SowQq0JRyEFijB
FyQUdUoGj8MK52PhAkVkIOYx2E2M888RKKmmk1llHr6Z/ppiNY1AxI1Xh49CySVq3A6ebL+wDjvG
2GVrdsmpp8dg+Wkh1X9yu6AkarfRVcdPaYB8mY7hraLKvhE7HvdAJJPKTzKLGrXfcNS+oN73Mmun
VvCwtSrEo9nwYNtTzQpQ+X/lgysVEiu2ecMSc4R/Ok9a8+6mwRPbJIWex4wPdFEurn4Zu2MnJJro
YP1+32sYBlSP5CnKBPWzd88TdA57LmIU4CyyTaKo5GjLa2KXs60egGLLM6p0IlzrwDG9noUhGvsE
9prDkq2b+i2Y7xcuVb96MNYkgtTkoyPzXzwTa/xfoEwqdxr25+J1zxMjde1erSCxY5MeKjDUpW8w
do7GzgdcIbvdwPC50AgrfJykdSd9oYY8h/E5sD7IrY6St44KWscvYPJi5t2zKdfmarY0HJTFNoU4
d1FpmpNDJVfRp0uf6g1RGWdRoUa1zZaT7TYNyyXw2vsrex4NpLuh2I5fVi45pO44Lcg01DULfOSQ
S3tR4K2o96KrVnZlPIZ3yzhJDCqRwGVGAfupIU+46D2yQ4HTYRgSwxuWhNk78ot6S33FHzW1tmGe
cGFppzEYyPGFOeKKtyvCW13Q/84+l0K+ZN16cpFOfb/3FftB/a+NQ/8Rc4DP6DJ/f7asbSEH9G0Q
emh7VocZ9qDOmNEPvrMlCfFtVMjT4w0+MVNzDkMUnN4SAuiSjFclmPFzkAR1hghR9hHBja36cxOB
GXzvkw8kijFMDnDyxSQMRMNOrPJFI50pO0QKuXY90TYWquZVLAdrsztohGqfbAdHDW+aerrrq+k9
PxP2Ikn2k3cK595/CvhejNJabjFubkS+JuA3peNEB3yvjBsXDGH0+2WcHO++52y0ADDO+zikmdxL
uPNdk9ZhEh8k0TcNa5Ia0B4SxYeZFQPjyhi9aWjVtSUDdgfifXnJOMD/DEMXlsLnrJB3KtyW4Oej
4a6493W45CW3RJ0KLtDR+/iX5xfcGmSgN6V0JhAuxyO+ofzer7a66uu1VDPUAnic03iICikJm+gZ
AEOMF75e2UG+IYpk53Ovm4HD380IYHfRAMkkghffuS+u4Zfwk9Mbon+F0rNg4NY3lrerJHRw77bz
diXtvqeEOHG1LbSHRTxW90tvCgWGInXo3dBmgKPi6mpJtm2zjpxHzyW7bZE8hWiZb47deBU04HUL
nENudr8UJkLxrp+XVn9WD2alMuLbSZ4oL3p5+O0rPXLxeZwjqRfjHRE1TUpCYtA9Lm9K4OEVH7aW
8wC8VPoWbxh1OXrEpPdtYDpF/DT1+LMoPfGuUQS7Fn0UqdbU19XWM15tK43+yjjRugWErT0FG5mU
bviMYCUyMWVzgy7gxZCuFnAcr7B0fNQZoC59Z/U0juX2hnS1CuW6ExkyQpVa7Uvk/xBr6KaYgBG0
Bc6iiChEOsyiueiE4xDHjDR4AnjyD4gFUFvHQcWsFJcGCUB7zeIeWSGb1GFxyxI27n9P+G/anyhL
uWpeMIr+q4wsVVa7MXeO6gqHXR6Vu7pF2IvOYgKFPxgkAqbONlTujCu6RBHHSfNQD6GNb3dL5sLX
exL5LMx6gllH2w55bgLp10IJfZBbHFpTJayz1o2vPPU8fUndNODNLkchn/VrdVmDuzlnaxA06BDc
LP0Ed2RgnnSR+H2ulz3id+w5cj88izLUk+PnNfVS3Efe7uVWGxy7xN/OUMdA6KDJKJmxfsZPDq+X
iqjfeCcClSXacMlMk2gmVXCYg65PLSWaNQO1A0EfooXwcTvRnqgaPFFiFmVs9jOdwdqXmrH9Y39I
s5ZiUEvNbIX+Nq95EY/z1jZJm5aIJ/NeH024nJtjeFPJaAI1dPoCuCPc8DozB+epYur0NBLtloGT
YK0f08+L8i/Dg13ALVJrXA64hfP9QqMW4fzT3vJ6agL7oDtmX4M70kwzNuPJSp2eazW7e+KM5XU3
F2zLv8LxGjVDUoBCABOoKHG5Bwr1tGcw18/fHK+Q0QqgFTHIqzgwKxAxnyAcR3WXWEVEGkrKwg+L
1jI5Zo4Xm7sT4ADRAq0K5WeTOdr5w7GPCx/LyRNHVF6DfuCYo5+xGP4v50q21OqfEzx/tBTxJGdm
Ow+b8lu1Zke+bBZQpqoq1y+luJOto7fDoa+CoQRne+ZwsLGoFRJ3eMUDBK3jEk/CwA/vHExZQdol
pxcxcrTV01E35TTTewieVWfRAzPcIGbZ6HCsgrcnZ3BWwiktNthDYx6qVy4HhMNGksf6v7o5xDKw
pSLfTWxVpv3cJC/anYaQJjRdlodEC3UaTi1XZMk3o5ZUDPbJgOZZ6bcJh9BoT16B/PRbjz8nNbeH
guHA6RZMoEWpEY9d+LFN9CNIkP7toILR+NnAYhzKQmOkwuuEHPE6GKpnYzamWvMxH9/bjd/7lnF1
dajq0TiqtHmgvgyFKCw6P22bLuzIz2ZbcWNQPXwJXCKEqYFaDimS7ZQotcc4P1OmkL9tmP6VYPFm
rqbGpo9YSSb4fckvBzyfkwmfQqYg+O/4J/f/ZAwWVfFtIVqAqmDw6hd3xw7fpt60pOrhUoIdxy2K
c7L4g7TFXeBekXby/uXF8aa3/rGrTtecfGu/ZTv1g0bECkj/MqaZFx8w78PlSyKxyQMrEe+hbwyh
GVywx7w7abkKe66lO7AQg+6bie3s7PjFOtTC9F0cfrdLoP5FpaOVrVao2XRGjH3XojxSDRaQ9izg
FkJ4aHN3y+Cxui91rGV40ahJn1w15QiwO81UbVjnqPRolFwW3J6Jvqlr37sLT6E6YJ3mXV5cVibQ
LFDXyMuwUZLc/AH9FPv6DSpTdXO9zCA9/zb/hJO8l5Y7WcTVf3ZANnhRkLnSqT/E1huVkDcQQ3ni
UYouPY5+pTAeu/ArDYnyDvsSQaOVqu6EapI2vBRSxTgz+pv84H80A8h3ZUY+GIwXb7+B0XRtYoHy
UFyRAAks6lkCqD4LDocwd1Aq3imKZDGQgrNok8R/kpG+gtPTsq7OCCATHlZPMckiJdn+MRyiyGZb
bnEa+wwubl0OdYtHHzR1Bg3qo+HTkUMztgdGjLMClhRRiiiGtOP/E/g/JTPod4zlHmBdHYKovT0Y
Mg5s2l7hHPVfdMALwBPasaylqui1hXArJ61r5GR1kmAP3F9sRIDDH3vmxJ4ERus3VQfsmbCQtCaz
eChCxxtFp+a2dngDd+8pmd4Si6in+SkVWV0TU7nj8DkNhOrgDhekV8fHY3JiFusNRk9+pugr5R0w
IhuekH223fwlMLtnWAuC7/Re4i5x7xIqFIePVzkh1iOh3gbcvFsUM+ogT40NAO7venEhtXKizSNt
GmhfV0HTlbqjThHUcR+joWltK5DdlE/xuxJHqZ/YgukfBDYtxjecGsR9Pl0fuyumlAFVCLfj+FLc
G4dNyhDX2XYTx+WvDFHqwOA10cYL41pDlLgCZxJMmtbvm3Tpmm0f2G+t2bZYTTQ29KeTmY81+9uL
t5fdOVRleDxA6nIPQzddeST0kH3A/FLJipdlDA6C+XsRmuAiCyZZqnR/dI0UyFjoVYmcyFtJ0HCE
ftSprpB21x2ZSSxhkRsHAvfHpTmVSQQsCW3VjNPwh9O6U+IbL2+a9WthdlS8GN5o+4kttKUyBS9s
eFh6u9+o/QvAHqZuhn3LMNMSdVdVt2Pdegzguy6Z0eXygEcSVlzf0EicwMoNS6k2o5luzAlYAdtT
jSO/wg9BYBlIHtxJcOsI/6qrZyxejgO/M4Z0HTxPbBYk0jQcY9T0W1toIH2LSsRjHtImMacWJ1rY
EtmMicIcPf1pSYFlDHgaLyAv9+PUeOdyTzGgsiuwVkoL4tl6VQOR0fiUKLnezIZr88X/smVJp3ba
AUZMiSzQRg6YM2xp+fGkSFhjWPp29E37qT7wP67be94dqE+354pjig+IpQyeR5WP/0RI2f/ywPh1
6UW3FaFz6ETi/Paki/JBErl7jU6Be/mSPj4b1LKNPwxZ3PFlA36FhKxc2vdWEixMApEpkkW9N+9j
dlOO3kEctd21ShX4o+35SwSTexH1wFOYZlKOMBa/tww/2nCe041R6vRL2UuSHAaVzCpPz8/xTB/N
U77WV9GIPSDM500VsWKUa+DG6rrxpYhb7O0wtPFgul/+r5Un5La29zpCav+uLI5PHlvKoHwC6TYN
j+wkEnLn5vXvF4v5pLzMLb6GTXqE/VTFplwlv+h4OQdazpYWAYrDKDzBKh3iHtsc3YYJNJiXm+TO
jl+BhMYnh54C8PYCK9oDcgH8Tyf9kJgISpsrcJdNWBj1Muikvyq1b7RS6J4TOl8CJQTQrFlkcsuj
smfeVlabuaQm5U3KRfu3IHY5TsZlHHMzJuUEFoNKz61TuV7Vb0LExLulnQZljasMK5iMcBIWlkNF
egWIpzJkqlVOsvNyUgN5+crB4hsMEwUMDjADbmWavbi9l/oDLzHX41+GUcQDM51RbS6cf03PFyh7
nm8eEPYYCMBfVxE5+ttXtf8vWga1+kJCIJTN6IpybSz9T+98p0W+OGTTEKqDG53caUepjYsu0OSl
/IEjgk6RpOa/aXm9T2RZDLgh1fJzdB19Nex5bnr/nW7rpcryvF7jl0lcOPQBMzYwsW9gfX+DCFEh
KQ2ZxLb5PeMl5ir//ag9azMqtsS5d70fsMcBhDy497aiyYmdI0kUMU+3JoUIiovjjVstJgh63JTr
6Ig+OBtzrhuw8mzGiaROlbSoeB8RCoSiBR0kxdVwx15Md7eXbRVPMDCyOmoPRqndb5XgxsnI18tF
tfyg/TiGa1P9f+Ujnc4Z9uWqnGogl3jYKr4gMSuOoCFNUwJ7LIGz9joR/EfFkDH2ftLU3uTrKUao
QPQet9YxhrnppoTcIk9VtBvlJ9L2SmJPKAN1jO7sAODzQB2OTibtZO9PJUuVPuJhRVhhGj1dGK8Y
WA89+8rVUetJod1dodHyW6mUafgotyu2camafCw+ASiS3lLBO0XN6744Klqu9ikfyB7Trv69Qbwn
msM0WTGXhnBpyRbtKLw960Y4rrcktYMY3OQan2warMepo4iHiCIFa14OIYj2Ha04DejFNCDbJU2r
A42CBlGSPHdOBjfbQYNBBASHDSIqIBjTdVVS7b1pFMg4qYAYV9XKO8mCFUWSJ9yZ31F/UuN/COfc
4BTbndqGURJ0Etm+CeIOkZ7Oo264mrWwGh3gQpWCnDXS2mbMlzdhutgjQA7SkMvh/hxePK7m/6dO
GKJzQ5jkollcD17PF4snQZQXOePR8q0ydBJV2yTUotzRz9izLXCtAdUcrC+5GThqNt3IGFJM2crI
wFT6TrJvCocKhYyXgC4gAgeNk3T9xLuHaKg7Z+cLk0mu4rdbV2VqZD2/fe/aIenRpy2ToFkBa01x
p7Lz5wIyhOxGOJZKhkdL08gYP29fZ1to/Mzyla/vh4zv3BJ4Mj37o5CwS+cYmNpGk0FOT45NlCXs
mZbg4mNiTwbcBV0jLK4Aa16pP5A5W81dOjEEw5BOVmAF4BtzXCpjjmyohAD4WSAsEOJQyyYPeaXg
oKwiKxf2Syv4PQkdD3ClPE5OqWc/WXVltTMalsLj68UrQ0VOkZcJP0Y+CUqT0oZYhHXZMA7uw5KY
3wxeF17y5HAbX0TP9EVbEnWVVEoXOYlgrNBPaad+LcLY4j1evArkobplrTv2nQOi0tjF33KliWoo
XZ9OsZlWHK6aTCBnTZlQLisVPzADs6r7hGXmVs2trzluzEf25BEKCUeI5zB9yFyWZwPnO4Yofk3o
7/y790lZ8x9nyJIf1YmYr60WKbppfhfqhjNQ6PAL3vHzc2+BilIU8d0BoCHJ/OhInuJ+mn1CERC7
U/PTevjfbCnVyu/fuUZnwyhDMUah4WyFjKEPakhQMEzjaaO+4GLIe9GJUI8aS86LXWPlP5fOmhZ/
r6RiaTSRf76bVF06zFsud76WbOfVX26tWyhMbk5J3qWS3/gmVSc4H9mu/gwxHp4jIF97oLYK7wst
H+R+mGgz4IzqfRdIxyN4T0T+hmeJjsxQNlrQ4eHsXNdyuVQT4YlxiQbQ17X2NFQG8Sa0I86mNRwz
gzgEd/RUffg3UDTJC8EWysLwZcjCSmIhtdoBIi8pILPJ70YnM7FTHed11YUSGsCboCR+HrgIY3xI
fL6GPwBeoF0rhmczgZxeiwWX3iFQOGytZWl+PYB/ClREwooebuAPRopV0zdoNXItAJCi2FzgZD6N
EFFnDqJ41ULGEDA085aDPYHcgM6a53Fr6hJXlYraCWqR/P4j9GC+JYiOgId9TU3uIFMqzqgZSqL7
w3CgVBCBAF3YuS6ASWYHGaPLXScNb4ODk3TYMmT3LQGqHKAR7qADO8bt54j7va3HAZD9UvBYf42P
fa0/H1yVMjoc9tt5jJdZqLvMeNOS6kqBe1nLPs1ZvbFUE84SbBobk/uC1DcLK6ezI1H5uU2KyeZA
CihhIBna2mQCtQrIirmtYWU3Lh6XqrNnTbac3/URXmzQXbmOIh5x2KWdvGUPiR4jMJSZCR+iFuBl
HHSx3iIiAHBWr/DnPJARfuGmV07m/gePaxjyG75VlKl/ZhCBpl7KYJmaOD53z99QsQhz0JbBAVhP
rvgtD890aiSqHEAOwJKREEadZN+tVJWk/LaFrh3tlo7t2IXpbSLQqmRly/uhMY3yvpQcBW8mkD6z
lfHrvEzhikGxDobDU37fwQYcImHRq7ZiYkpA9nErPjr+kUfG7JdisfpknveCqdVDLkA1QMSY9a4K
Z1BvwcQSAdpgJQx6H44XwLJABTsIW+Xfz38AT2RQvL5tFgD3q4msnwaXaw6PBezRv4Hn+a+AlOVG
Sm+C/ModcM/bJ20MlZUuGjtd3kvlu7F6cpGIGtodxCi1TT3ATka7evb8VzzNicp5YXRzrE5uyx2d
o5xj6FrkBQgPcOUkjxLcfiCOro6blUrnrHQ1iVDNBR44B34e09QjR+khwK2vRNsYrkyQXIWQnoaP
+v8fPFvQMgBo/LYvF+mSqsop5LmeN7RxCgcI7UVRqdfEhVT+2HQ9aCYwIgYJCOOMTr+gdPJApIri
T6MMzd/v0SA8fEM740zzHeaJ3EvwCv/LLBaJ2sfLgfz9PlqcMgRegUe7CFAATO/bkbHsyKvYijbH
Iwo3CETTYvetMk0O/7dIYwwQh+PtuGCGTL8D5glz8UyNBZk8ae7IAIKV8bDdpjdJUWjYUPHxeEko
v6YSyvp/bRLu/1JaeH7bpUc4rIAY9NDL/3+3Ts8rzaLWFF9Ew8fNpwzQgzhooqu71FkWt51efQS7
JTGbMkHznj3PDrnGakBhdFMBMTI1fNdZpxJz6cKYK12ewjEF4Wyv1BKGacwPEYt1OJXD1enCJ9jn
ypydUAN1xzLosAeM78qaX5D0YsxcKB2LlzGgAlI/RKbQ3S1fvpizYjPXBKSpBjCTwvg/lrCcI9uu
feJZqlzNBWOESyHcMjNcx3mw2WD5OzUQzzb0JqDyIc8NE2SgQz+6dqVgAVvLJhCmuCnk9dUxAlGh
JB8IRIW4Yb470VEJQ1MXGPNWdoBonxMGIN6gljHSs4qOaU8m35+6IHYfT+UdIHJnFhdSeSp0vHqD
vglODSVcTaPPI/6tDCeLwsO3Z2mEmF4xETsDlde7IgII9ai42PxZVSmj7e+z9wMY5sTanmclm/S5
bfAvibOUmyev205Q4SptU42q1x6zxnZv50qUn2lMG4xAoay54FzcgZngAr7EX6rRL9SC6WTqtSL0
7G6JsbliSdeFWyhAKNlEnj+aE4va3g/48F5vT5q1+0ghCrWR5rwqPFLcEfw3DtNrfasJz9qD9LYd
rqWWV5DEE0lca9/a7qmxLs7aqdPx/HnS1WbyR+//7hu7Q3LV7/6+5C1CWB5zkl4RufeohMmaeXE/
w4cNmPLwNCwtqhy8S2/wYtychOhWjYf7+vh91uDc2Rvo3kh4xokXG8ScQEafnCZtXGUBOWmnGzo3
zJTktMVhhOQta7C1I4mFTBbqo4TvMYQwnm4jUMJy62uJE/t5KYmnwduVLE8KktANCmnovwVBJy3s
DoqgFlYOvFt0gdWc9WplqZP490D/JKuYhK6/R+zLqiC1TmEPceogqqcjg/LFFkXvtpTbrpBX/Wsg
0biZERDHXcZriNaB2xM9EH+Cb7tCTpw0yXQGtbupdFOuTDcoSqOhckqz0SdxqzXHJU4Iueds5AlF
XSCNuBvlBunRaDa/Pe0b2A70O7tzc68sxew3mdXl+K8QyldP7DI3vQN6srPXZSsLZc2zsMkxVSZW
nuu/fj0XzdN5aTGedY2OqJFgmPTtESQXDbh7CT1B89PjF6MUGkavc+XflYpowzb7NXVpiuv0RrZM
YniEaeJNBQBzgucs1bAN++QyJWN0VpRnpoRvsMpka/1eGGB+xcZoZRrCehGSPuDnSW4GYsKaPrh7
RWFEvfVi7iwJUKLm7M7GwyOz+fOMrCCNRsPTT5+qPT56NmWoDLUBOH5B02sq+2bbmimYBxC6sVgo
aqPhaE3VAu9UW0+kRrrCkIdBC3LUbRVIQNyxZLhJEHF3i9l8rZGWI20qoSSRMTqRaAo7MCKUZfK4
hpIFCFLxM1T0yw9+OSpTVIpjMmxm+WeL48rZwfWQi9Xg6mrlHrlVUncx6d+CFabFjVtiSZlfREgB
lJgS26irJ7VnW/1eLwFFaApKIdW8XfnJPQsqhFbru+7aTs36Pb8l00GPp7l/TrE3tHaI7hG1F/V3
9B41zmR3eOlrMewsAIoDV+0rMM5J8rJxIwcUSKFtWmRdKbVF0OPuXD57W4XoO8pk9iuhajUazjo9
nOiU25/mhK7ybjyu6SsMvN5ThjT6+iNARiQEhofNIx+Am6mmRQ2zpkPOLyaf7YeIrjS5vr95DF7L
Kfe8eRlsagXvD0z1kLzMcnh+FyG0whBTfAqw91NCjbFElt3+wNYR77DlCNgA6KVMv3CMxpRXfMN9
o0IxWXRZ08V0m8KTlbAiPpFcqhiJfi3wThsIcYMjj+ibJo3v3x7nf7IrvmiRq5oZOPOY32KeVDnu
6JbCZRaXuL7vvjHCVMHEgDd+Ehst82q9t3IcMMzAX4RAkq5sEu0jSc2D1DbMc+RA80XYVuei8wZZ
cKgbkATgKmII1YFh96SRClLreVj0TT2oOUQTQFJwq9T2R2CfQyHlDezyO3rQKBobVZ53mQCInxdB
dDhIcmG5gM+8RWIwX0kL5GrWXGDSLC4c1lcrMCobfHt32ULlj9HIPrVtXsrc6XUC6XiO7oKW0sCY
nLH/jwwYtGyxFUTXwL18+x/v0YA5ooWRX7cbJYxr3bYQN8GXhthe87J4F7gvgxR/y9iPVMDBi3DQ
E8lUJZ/s+Js+mPjOtP0W3gUcA9j35VUbwFzC2IGnaNR+zACp9QuvrL/+hn27wfJ8Bm1tka9k2ZYI
nxYb8G6qs+codl7RMCqOavX62SzC5/auQEg0qgvKpm2oU0pgxiJN8+24O3R5ozbaDPYNoPS5TNj/
36mfRB2QzhltbbMMKTMtV9Z3pLgJd+n088btawhs0m3ZZec/ZnL74pWHTzszCbRN71ayrXYDC/jz
+Ucd8+xFht+5XexsmW5sFhO7ZJ3rooVae3Z1Joom2bBiCt+2PojJC2DSZZzcjy2J7mSVn3Ydg5xN
2MXJuyG1K4zfXppCinvJrSl3n38jSltM1Vi/UmeYlMkC7R5hWdLsGxObrXWBxjBtz3rw+BDxOAsh
XdWzLnThfqhuzXJkaeT3ztCHbECDyfEQyll47MLBdvbdb7fzjWf+WWzpVnFYtISqkKwqKaHUgI25
eRmKJVSvVOJQVS2CZZwI+nax6OON5VPAdC8ZMV5fTpXF0axCKWM46oAuUKPzHJusDnfnvsuzFx91
qO6UNs8iVDidUvyzrBR++C5GvM+IBsf191zeFIJWXDiY9dxgqNpbbFePbgtJPx30PtXwomZxk0KA
gC2pwzSK66ynCQBzxD78RsRQtgC3lmWeU+3M2mlteUZXyGf/kI6nfDpP0X1WVfuNF9lFkXRdSvcI
uigIh28tksdDdrYbsadbdC3gY/qEHqnd57tmsujMO3+dLKKe6lhMykL0Q7OJo7qJ165NWZ3TW6ME
iZpbJCXxo0A+G3lTY/nCms02rIZ8EMARTP3XFsxOuQ1NqyntA/foOENUzLUzwC8R2ENuIzl/mJPm
z1yh0rFI8WMvrAd7D7Lb/i7qSyvWcbgmmrlyISmaE2IA6jnPwcEFloAuWMHU564O2bvtdZ2yGIE5
EfRSFXVYtSS910fJTY0sVGcqTYmFrZGuTxVkILmLeud9ZfpZkb0qerIDlRhrsKfkAyHt1uqcr02s
iVwN1Cy5NA4sbPiqINEvbHghM9yZFUaqGFgezwdyJDOeNEA9hFtAEI/fqYJhxJYX9RYneigw2fNy
eu1FmcmbL6wtRMFg5s9a0g4Cjt0GQnr+idwFF6oq9oHPxGvdPCibdDGr9qFjMnjSIsSoA4m0ZhOQ
BUGi+WyEBwqp2ZABxthF8CKUDrkWIcYwQ2ZiQOysaN1jQv/Z2U06ued6uD8/eEuUetIUrTfM4ywy
js7ctDBnps/hDNI6nJWIM3RtaFjZKr9aI7Tj17P5XD9k/+uPTn/qQS53/RFTC85LNBNcpXVkh1kp
wFFXjYk8uOSB2RtAOy7AOKmuo7SA35sLM8GHINt1X+7F2s4xL9LZEtoTZiHj7yt2LLZJPE/1Oe6i
Eu2p5Ih8VxNKPKWOMKGKPBi9/0hxRyKuYiU/gwFAXqQ0eQhp97YoyKWQbHOwf0+nrEABB+4Jtl5W
Wi2lOTk5ge4BMhnIC4KlyZKi5bYrO2fuyXl8sM1CdaIsFqp0C9BBYW6+iGNOwgYwbGE6alWCcCOF
d5tp4pOlYMBRQgzVitDV+d9XyCyoFP83t0Qe/8TRcU/oCS2rmjPrv70jQJu2qskWSmOMvySakURW
Rlqo7ENXmJkqIQOjTXIyue5nBFHJnR4FCKTKQlKyskv1NfdvjqtXA33O90KS8zMJH1NW35qDbkx2
bqlVPFmNWgw+rfbLtoRewyA6/oQU8YN+Vp44PRaNWfPVeGig78sMvJ5RhWqzDwIGqaP5DsKC3AUu
HFlAi/mQ3efn8yn/QjPBRfYqHXJdGiUvpuehznzoOVy9U40p3QnxfdttBxdFG1+nVp4y0cfGNGgk
wSyLCBp6L1mBPzTce5qSsda2K816BjsFmENa4L1BHh8Q9TIjbMsF0cW5+NznMKPk7AWRJjOi238N
YZI68m7CMCQ4anEXmkaL8oXrt8vHrA8f+BH4bU7rsafWZpM2e3dQ98UHxIlCxNYX2X0jPXD22L4A
j3GWZrb0KOS4m0SIJ2lmmIwR5lvdlH1iIfqtX6o4TwmOhS9rQBORVe8g7gIB0J2Im9U71Bzf3KGj
q9P+WUpJs4mA9tKFogiQ6DiGPYixUa8gi6x+E5Ovh6qrrwxDb/hI38RBMFBbGtsNOqSBR5cRMQz3
C+SjfEUrk16NvBnwv9pKWFpz4pOGv8kxU9kGDBATl6B9qtl0B2ca0wubJQHPGCihSwN1ci9QSt3+
j5omwmL1wYRS9u7uSMF75kZjJRDFaIdQpjv9j3NTDzec2FgdwAf6pUEhkDcv7p7+1rAOsLLCPUoi
2sdkD4vSZMddlu4u4ZNecu4hSKVrBDtwnlJv04pCOgutqNLj9QDSAxrp08vxz7IsO7nKZkMHtHzj
Y9brDfEQMGp0kXP8Pa44QHNT/FH83Hao0ifu7E+Ty5jQo6E3BLpyLI7Tonla2aSqfRD5qaIw+Bl4
i0M6hWNuJiIQ2umLwTg61vNn69xueFLPyy0sBZsAnPa5sl8JFXc3ZwpEvXCyS3MJTF4HV0FlCAXg
6M9zPxbB2MEdWVD6njjI5uSfyS+Gz5+gs+tioGyG0UBItK5f7rvstsEch2fjfQq73/ur+Y1IeoyO
F3viGA74DvP2e0Zl3Ht2lEFTbvZS53buciqW+f53Vsk4NA2I5z5FsvVlanEaVcKJPzW0ScxyZhob
+gGai7ZL3hOjYVKziq8yixTPbbirwRlzYw9tP0AjN1KXj0P9aNjJNf9d8eEWAuVxNw39RVJeICA9
7K3Dx9rE7oGbhMWby5mYGh+Z18hnmU7dGn6qhvQjM17Y5tSfnTnKkMr30bqaXwqRdrKa+lQMr/S2
HfsgYUwRP1iIPUC6ENr5XcgN+XrA2e7/eX9hG1aRQSKDo+K4h90tBDgO58sKHxcoqpcPl0Jd8XKB
z9cBQfolAfo83tL75eIdOVi69C5s3pxu7pOmKVOMcitfw69vqpn22y8YYziTvzjrX3YtExLkb+hB
uahNcXZoJkV0xT9PtVc5n4qBihLhUrXhyWDS9dUFbdv7TlRu2QeluskQiinZtd0/WpzsRdymqsuK
hIgUAhXhARh4qiot0oFZTulXhk2/RPP4hAWTxo+rl0OKQGo+oA/bh+xJI+dEh1uE5l+HqzwweoAK
JJUgBrg60Mt9ifGBuvztta4L7l6181fUiyaJynjPJ0gGIKrw6HSVlEoQUEtC1+QcVfrTT3QjNjHn
Vy6tfzjRI0YFXb1MwNqVXetBrf5Qyj5uKmOMW2sEiAXiIJLWo9LJuBpEhcpApPt6JYuLxwZL1XkZ
v0B9TVVks7coAh6zP6M1Wa4Wymri8NSm5kVvJqrLt4vvps6R3YBtbg5P/St2F/sYvP6t0GVVum3J
cgqR4mR7Qkc0P+y7I26lec4aWLeiiVbiZ8910NcqPVWqsd2SxQJ5ictoO/xsOI1BnhMu1+RGRUq4
tIJuJwCQLxlqw+hoWxcFf/cvzvUzMzeqJpZZ2DU4TZJrPrINvjNLLwGfw9RLOeHxkky8POdfCI4i
KaZ4jfsG11VBY3tE3eiWI3OLFVL3h+O40lICXKP9eEHRurOoXbgqUdrsJN/5yXCuVoGfXFJ07a3Z
N8ZgKKaLmcQhTIOg9K4ER/YGHlQqxwxAOIUp6cUNY+PZpf10h3yaTVGnTM0RC3Yzce2J4JUfJm2Y
Ct2KVqu9j/6uFuAjXH6J8mZwMMmxPukLqK/C4DW75DF65cnz6nCEvbHPqED6aOfzB9OVujUAuqZx
9X1pyVDGycGpn/PZF29Cry6fYk0bdUqD8v10+WjLXhVzMu9LgkUsFRWbTGNakDBLdXvnomcUHDWg
K9DbyHUbOs9Y50LiT80A5gJAiFlUoNgOHnVAJ7HTGFqhJ/CJPCE5qbBf0gA13Wktp/5J+4jnPtV6
POtdi92yRLuC4Dir+Nb9Am8vajHEYsCI8pnxmW17/e6vQjnX8ujc2q41CQKlBYysNC9np9i3eAIz
Sw7p9y6RmPEyWGLTVr2/473HvPROPo+LOEidiRUNomGrUCSDxlYqI8VR3/E46cZQIlsheSvhosXr
D73ASk5vFLw/hnOOp2GMMPyJnvACUO3LyFGQ770AC8B27s7f4LUFSkot2Akejs+V+KSGGL/dq1Rn
/Kh+ntWQ4nec0fMsFiCIVQnuKqLpdnQyuCzFgMNlVpFWprYr6prYq0FyWpQlGZEZx9C917UsJ8xI
eQc4eMiuLcFoTwaosilzQ0gGl6M2iI/WCxGmWbta0FApAluo77ovJ0IFWl+oALiVaQHxeG9wYGsq
Ly7gky+Y0BzrXiH/bOzBv6mRXeb6IcIgT8jhYZe/iwpl2tsvPaFA7qn9qkduep9OcFBny613CPqx
9OxaenSa6WMd4yKv0o4As0uf9nqgENEyGuUubs04IE0kY07Vh4IRPyvp/IHscEzFWI4mwS7x2T4P
Jmr6q8vDCFGS6elJueNTGkZfq+8VohYEJgN5V9gwZHst5NDppe3eegZr3icPiBm0TNIIGwv0DVxI
b1hjTy06fonZFJCm9INzoraZEkp9HKVooRUCMz5GvRFzUHzMWhKgQtvk8/dZU7NIAv0/OGpwTXax
0D3l1uYtjyqRhVeijSEemU9Uskf8AWdgcAM1ZwCnGbfyuJHwbvgHoZODThRVHHgjLONpOhgglxSO
5K/Ykv9ZzwXbk59fGxM6K9FdMNojrtEqvebS/dlZk06ClcT7CSiXPRXrZZP/1vh1dyNzc8OWAkWT
fUNkkaviFUWNch9VHVkWLHDOQaVlsqdqSCvzx0UqSPtvRcWSMZQTDNenjltzm6QHPmVPFyVgOOFX
UDe7Es+04IPLlzm+mt34w6m2l7SsbQeRA+oWMCs1Bvbe90WitP0gt/TFdaK4ZNG2ZHdd/gF7fzxz
WPtu3WLYnGesFC62Pl/4DWuytK3F3IN67kTjbwCXETcAqIrlmCDHWexT7pSLmzotgy4uU9tGrqA8
H5CB9UYaos1pn7FWLaTQodbPY3xLTCpx3++teGRbPt8edUu5yzy+46QQsL81wuwMA2+KkzaIIINX
n/ddQs5I/XhIlQiJAUNFxMJcNZ3RY88HgE+jhPCmkF6UxInsOYKNX60YWot5Yjp5QX4U28VZn6Z8
PFOetjQAXXN3VKPU4r+fqupWbxcYBAbZO1SqYmi2TwYl8invxm0KvFhQpilIu0h7ZPT6cvqs0W4w
ncwlXBNxtQGgCU39TgtEmqZxNClMYDPbCgCxhd0D9QLjEf5cUHrKr5T4/e4cqUx/mmKjTxfgZoar
mS4/PjzWsGXHFBNXBABKdQ6elh7q6FhWJ/lWZkac/tgbiL2h9siB6vQdbjcwXINF7Ijs8vkDl9lY
lD1odtrOLV2pr5knthZSsFaOmtHPktJcdBMPD51kCp7jnOsj4G+myZW1Dsdr8ZEf+EmgbXAg3z0n
wLPsv13ChhxQGpn6lXOryJXBE7qf8R8p5YpRCBpw+SwJbsxkCDh2lNiXESpaYDx6CM6ZzFPqDvxp
R4VfCSFjTg8TL2bwrqw9qQJS52jKLHrAX51IvHJNftEhakZbMEjjswYBZJifrAa/aLsvgrTvf1fz
frpYTY6iatwEUKFOtZujaGgLHqtlKK9EuEOCsmdXshYofWMEM/aKZSzh/+jWWdD5myVIB1rGlJj7
O361I0dZwFQZ+T1uj/cj4ObxlLmf7CUt/cHF4QEeNzM5s3Eydcy2Avz+rsV+5ZdzSaJydoWfqbRH
JzNUMm5JHaA26mEvrS4tTXUbkNRfRDxA0SXfQYw/SuySxhIkig4ECLBwN10PRrYYghkSpCzDoPms
0sXFjh6wFZ0FngQl+H3UGsDma4N4KiN6tIa6vGzTS0pS4qehqCpEeecdSn46EgHFMOASTvUwCnT2
09S93W2Pq3/BCdlJhW/0f/U+gqfbvbx4fm0sBewQmnzR3gRZjMIhPPGQ/fF9kCYe9eL0anfevdUG
wm3Xb9KWMeSMFC2d7dLyF/c8cSXLO9bbdAa5OernApxjMiuwf4obEDt9T94ljDDf3Qp2CDYPVVP4
ezDHYN7oRG59lER0GqjyVb02scJ9xYzl5TGpCKK32n/vTF950f0XwqlGil8rn3Vms+tzHgtXwaNC
QyId9UnqyW6t6nlXYkdpf6XthyKcrLoakL3eS0bY3EJV2R6ALi+oWiWLzSkisC7sVB4a6dRdyR0S
IJfNGl4duvHi5hwwWrRQXOe3m945YZBePeTv8MiT2qFIuSRHnZAW46nY3H5iYXXmYr6RsSYS4hp9
E9cJEI2eTL8+8LdXGo4dlKQTjzO0NeFmLdwFh4nSjBwBu8tGLT4XoTDwNxu4mks5HnWLqzS2LWw6
xmDA/KaH4xIFr1u+b0XognojuNr1UdQgrSRglwIUObEFOo2mTcVJCjXOIgD0QDZu3eRYJ17OkWcY
d8pFLPK/h90D9vJDbiH+e0mUGUkXh8IA0GdAeXlLyXdEqE+hSkSdOw+7ztkDItrkXecegD/b97hD
tjwgsjtoiUElK5Ofkb0lXvSVqhCZOIoM43mYzyFLxtQnAS1LYPh5Q29KQt1+5+cTNg6lB0kdskav
P4bFaLocnjFLWRe4s0nhyZfItUHs6QUIuzn8x2IWwtGprndN6IP9XzxVUTSWRvTFRsf6MuZ+OWdm
9mDPdTVH2yf2JEeBEr3qDP8UOJIpypQVVyJfC8rpNpm7HLhARw9QG8IHMYnvwyb5Fy+5T5q9EguM
R7gYGldPy80ZC+wApimmU2trigkgbJa2i0IGYBK9VW4L/Rb80YKLWeHqRj6xi+evQ+b3nbX4kzlF
srpjKLkHXRaJ2HDenaASgS6EFkM5uHGhRPNCe+YQDz0SEzzxfrDCSH3p/+EeLOmIpVkIF30j7YvF
oQNL5XIf/JyXi94uiVB79iVEmULvHissRkXimT6w9sfHt9SuJSncOXFMeySOfoKVi54JtYiefh+o
NfdxSOo0cASInqX2KoHlaNrcubpPZ+f6Mh7ynTFAtmggxBUPSYOWHiEbuC6jYToZTNCwtfScUXjm
v4K9NjnNcbp19LGX/nllnoSyBlsdyr2zloh8pDNdhr+eTPqzJFk3+jgTc77S9wUg1z8iQf2rT1KX
APUnItzGhwa8aEtjvddiSbRXXUVCbtdLT2UQUv6gpR2HHf+Ve8HMOVf+jsr5j9GWoymTPBCXwb8I
l5wOY4UpoB88iD3Uji5th7jrUS4OVFFxDC9U3KM5e6M/01a5BBUjPspIdouv9d/YuSu7rEPwIS7/
MJNpt1XCpkxn4viYRpQK7UH6DcrJ5SvyeXZvKH5JKBCV03dQvUqGiOlyAxnXrNmZR4lB6Jb51gFG
H418pdhQ75xYQKdOLEFilQOCZ9GozpGNA85aXoyfR+dTYm0vLxD2IIqYiyIOEWVfujJEdNv/rYtZ
Lgia4z5FDm/REKQv2oWn3oNOYJ6dWoxslHApwGqsEe8FnQypDjaa+QD8tXalXJLiIR4iZ6yd7EDc
uxEfLoudYzgnPhzDWnoEvNp0okRAWG6xUuEekix6hiND0Y2daqM2Mj4mtBdGcsCUTuXXdtBOkQ5K
aB1OscwtKX39lSf1UdK0tEzZo8NAq0cUscflBzeMpyHKIm0vonPqP4cy5dOFhpUuNp7Q1p4E0GIG
NwIyXTFK3rQWc1fcCTRGtVu+Q+EUtQFXC2M0HeEBl0le2iTjdOlxWInwwQxeKgNq74IycTPYTH6W
0mBFV+6rWkASdhoua/7mwyL9itx5JXTMuPolPLG541UWzOuVFI8Z69ppNQidr2uZQ4ulUm2D7WXQ
/eHcFsEkRo4EM46iB3NCTYATIxYNKFFWwN4Ln2f2ZPfMl6YG2zYQSLgNftoIHFuxnAO1YDGaeo9P
4lyRnj9RnvKRNKk0p7joJvIHm9jV0kvF5gncXjDl5SIeaYAc41fVFMRgj4fJKsg39Lj/vDfP/QDJ
8JfT0r1ZBmgEED7xM3/II37ogEXVNwIbGgS1sdT5idaITktxq63qhPCX2RZi7dX5UQWiTenZ62+z
nf1QjZI2Oo2W7eKPyx+aImHYc4lFxBYNv1WlnSVNQ1Qsjc1r07E6MhM/ZoLIrBnyPTX8fQ4xnK1U
MDPVf4SerCP/U2JkeK25to7gYVcFkQKzFDGLi4iB4+2obgjPdAQZB6IUlIlnKVpW9EQejlD5OktT
AqymmLIaBN7x5cn0lQYzslHWa4w5oiH2FZobrbYztv7XqWfY+cxw4X84FVuwHutbElWN5GaxKfCX
Jbm+6Wn0hsQO2b0rxYal30U5vIg/o3kYBZdQbUSfRBmQ1PA2myfpJikVvWSJJO95+BmVU0RIkcXq
Ah0Gou7jCSWlz3NnoNIZIW3Cxzq/sGQLshlc5IogKHlr3Kl9TkDyxYX+ToN12vGAG96gRnSPhPXW
5BO4KhL4J4SrhYNiTevoqcR8EerGT5Vh3GzKdeW4+YyX4cmj1XtoC7kMofAkJOIz/Rivpy74AlMs
GlwO4QlrLAAp5tkPYJUuH27F3vYNoQ8JMmWoL4+mfHjPdUxJ3Q0BPkJyG8Diz53vnzeRrB4yyFDK
EkVegFoXgoBuIE8qKjh9K+DAFg56t6oz1ci9Ooi/r6YM+8/4+UAf1Fc9LwHnIzPufXQj76Bw5nav
bsNR41hhNjT45/zzD4iYTFRnvd+BPG6d4G4pteYXKHGIHifrBMC1ohNVRLR1yuHJoHI0Vhtppn8Y
5GrC9ByJoE1tR/6m+V9/HdwwSNUsTO4aTruumGgwH5EKBgReelsxKxDbCAl51xwgA3dgFes49Gze
2HHZ7OrpOVJ+RCjdoSVOTkUAm2Q70KocnBS0e8rQyvClIStk2+1FaUKEbAYlY+GwfwgyNl/f8Jl2
q3ukp5sap984LNUE3bNqxPv9cM/v2Pmhm5r3IWzJeMOrzIsx+/dr3IbjBapkQlspQtFTbUuptNe9
u81xZZ1jBchafysivWdv0fPIohURp2WGWbGTPFlODm0GkusdkopP/acISCvbhqONCi790SLE8Hx5
8hRoUN9nDoTXmtH0R66J9c269Wo8SV2V/yz67Zyt9L4LA2/4xQyZI1ImY+htsngy2tvmDW3HjxcC
48ZvHVFQ32k+qosgmlHt06dnJk0LCp4X1dS8z6vwdZhHgpg/zOmIcjUTnWyw7ZDiBWzMWgPwLPGP
IRFLZlGW5mVlreHJE8uDVnpYojEpDCn6PefVdmP1TR23HypVAG3AhhqOwUaAZyY1CuNAAwXDYByT
ddY4GLDGqABHzkeVT9xr3Aa9dXiaBnBdkpBZZ/0HkBq5Oa4trI//1s/JgbjIBZ5b0k6SGnJg2zJh
0TNz2GcNkQhTneacMj83mqQR/Pf9B/uHZUG/IZFQA2Y6fcD8GqHO0psE9T68xp815bpS+jlO+nrU
9cYgHFo7svjmarkJ4TLIJFysycK816UySM/DWNQOKEhJIFGXzYn05jmpLyFDN8cbDuaEBsY/qnrr
iJzpbR9yhfUuoJI7mL1gRy9vkULcvXVEZhAlL0pKVynPavTsG40MzmqKs2rgpD+ghyE+mbEm3v5o
DQipg7m0BscHNDNRgZQtFJoUxi8MUQ3w0Xg7/XJHx/qIoo3xzt1kqKGj9bFjDUC54iLB3OANR5bE
MtAZWilleervulMoH7aSKmo0HNKPsIGCkssItZ+lCHmezRZLww0/L+UBaPtULkxn0ZZw/G2aZiCI
2hvV+LdMa1hVEYw8cd306Vmi84+U40lC31XH7UMPj+w2Osf+sUjtnc2lU57qP3k5YNOHzogN09ac
dSLVbyTpm/VP6Gj7WqSnB6F3n1X0YjqNqx+o8rGkJXRw8T7P3LyD5HKt1i+8kfgI7JLUaFwtZmIu
mlKKfBIZ20pWWkUya4jmmrwC9mcfYM/QFQkK6/DzLoOLmPzfZmWE5yD+kC5fO7kS1TALF/i9M0c2
bR6SptYrGc4k/UrZSX/F+RZCxNxq41u4y91nMqlP19HPrWg6wxTH2P45cWEr8yVNPjsaW2BdO6AF
Ftjafhi2FVADyklP0J+9gSF+7V3cyIOG9Lh+tPvWr95xOozUf2egY9zIEv+MzDFSJ6jYARG0pb1n
sQj/U1OTW/J26GqRfd0wRuI7rK9MJo2R4bUkCp+i1p2Ya/3BhLzY20mwUQTwS3BNjzexgKzcfCsQ
0x6m/vSuC0ps/uTSzAho68AaPOO5Mlrfd9cTUK9Gw7Sm183Mt6aQkdKN/Y//U2buPNJb1LghBmhI
KV/dG2+BMdTUXq031XqmSK9ljlwQTUeGidvtc0hAg/Ju2OwP46cDST99b2DFEjo/XpMRVGGhe7O+
dRvYR9RWSihaB6u4/NM7YuKfk1dMbEJY2WUipi/exxaXZ2IhB/zIgexqxc9Ye2m+ruO97Ri7pTr0
JoRwCxsjJNzrNMEgv1hjI1BfxjCD5J67n0zH3GGf3+kGYM72/CufufSlPqQQyZHTImeFF/dRUadw
iTowvzEJBFFPWfANytW656MFsUi8ex/yqUFU8/Q5eM7DwLKafJVi/jTv8qJ0LhqTZvOpRSiAMdwm
or883KS2WRkpeHYo6DT2m9RvLKu8p3DtCsdXmrjoKFt150B6YOQLp/DyS9tnWKTMOA5vGjADnI6y
UNywCI1O7lgrCfNQxYKgULR280UxI/CC1qak2M0ht+acfPRYE3lNEYkAfTDr2ys8aTh2E+Wd3xel
OFjlvhJXJwh4MaOu+NHa8rzSEFXpIHt+OqnwWOm6sTFQ59WQ6ZcBtYgB/T164ojq3LBOs8gzTaZJ
Sh0NNxOlUo6TBZP8/LBrRtV2SGBKrV4feoWtzXOsjdkdoDyFRac6kENFHH5UTiz6vaHeGubUfO6L
i6WWXqzsEBDDaoZ049aFULApzo1tZW1tGWjefSyj9EUfI3TcUv9LkzKF1l2kCghqNwNcBALdLgwR
qftgxV8sUYt3DGIX8BFYgTlQEhJKJBTQgMpBMMiADQhifd3A3cJcGJt0PBiKgsMHNUgSO2MRwm/P
ZB75LJwc2+1wOV9iFTHJutyXMtWD8QrNruDMQRZV2OL1yAV403hOlvwrTU3CRPDN5otVkqHj5AIa
JqKPzGBMcQi6/CXy7qVQOj3GWUTKvIY3zjWCNzwkXwk/oHUMgwCHpjoOYPAbFHAVQ1lYrkagAjU3
lAxzjOesh+j1rSRC4Tni+4mBmRL0AnDNgZCZwUy8ZtDEthg9XZqk8+27MsMbDKjajXSlxfA6GS9u
TvAKppgP1GQTnleondK15RqlL8j5AVFSxXLcXaPwkxyfgdM65IwerSZZn/CBg3QiTx3ZKYpqW8LJ
hiFcsv1HmAlYVsBuUwsmGCG4Rx6Z372euu8vz2XB78Nsm3d6CnM6/+m2sPzHpcb5uNQF/LQS34nd
hZLXUqEOdjPcnGmrXVZIIHM3XR3f4m+yiWcN73GUqEwUUynR+H+/mWb+6koPfFtNdKUveWhnWWuY
9+rE5q1M8Zqwm36cEqpXbkgeYcIUD+6w+4c4bPKoJi0FAFZbUVFWu43ZT5AVsls2HpG9bW8zauUJ
kVy/igwNEw1CsohTCDZ9U0yPEQh27I4Y1d1Jsa2LhJocYjriYdY4fkkZ5/h3JU32Dy/XYmjDIXZI
xY166+ORNoPHIttgK2AJG6Dnu717gFrVENdEGHJTs9x11IhL8RQJkMNvLv3otAEg+/6BQF6+7oRN
8/rEgoo3hHS63dd7VTIAOOkLT2bji450SxelGD4yPQTKQZAux0zfpxuMeTiEI3IVScS01z/Rh8bw
W1ooWpMTCv6BlHVX9IPfEndgAFxhIO+aPuNV27mrp0mm4chmUV0yOQ1Sp1i1rBGSOmvbMrMqmfZb
NiReOE9GyK3GxhmPAgtimUh4UHF24mnheKdRJKTT7ciUvI6C1T0Uaj1g79jfxMLroRPhe63l//UB
GcX19/gwNS14eMWXR3tKLdzHIRsNxrs7iIkmt13hy1u8Eda8bg/L8/gviAzS7HhjWMbEVzBt8vhe
mjOv6i9/6NcpMG3fDEpqeOb3RXtSrEt8rb1FU6H03LwqXcIH8u3xBu2BoLy5jyGKc3HBniMjyxwb
Es/Tup7gzOsE2E3vS4tIiM6Nzd6kFazC/qY/3TyxgQ0pLLkBk/J33H8b4P/Jq677H4k/Ih7cF4Qu
wPNxrESc476GgS7vVZyLL72vEf625Zu+Xy/m1oy11rg6ZkNtQuDh1aIMuBWMV1MYzR35a2n8DsZT
shDr0X1XNwrzqCnG55mD75xWKNIHHPVewNsWcHjcvwMkk3VsNjuEIH/dF2HzbKaw1VnrbpJzDGt3
/bgd+WaQd0DkLZkZdg8FA7hnivsRl2LAnY76mBEJ72tERcFKpcVyUxMXihVlHTSs7pWJnxJQa1PV
M4j5VjwOP8eri5uvD0ehbCiagVHZDe59/JGaQmpueT2VUYBCMn9rcFIBCsu3PO115AH0Qd/Q61JX
lVMEBMN3cwPQRBwF2lv3QZuzFkmd1aUvkKCxnmqesttXqs+joz7m/hUjdrwzMRYysNmjUFeZDzRv
FNjaNkxi9vy0p0PLWBb4oYjMHaETnGSHtgMZK0Z0A0F3yvxmXokZtLNT7L2dGXj8ibpcRy6hEcdZ
lolKNEd/5IvWv2IArd0W5M9OArTDSQVdf8UYM+Yp01qb9hLvqTB97m2WputslN6ZrSLeCm56awa9
Tnsp+aZ8vOoQqGfqQ9EidZPH+S7Ivm7a5e3yAPRvb+vwBczsQsfwSsXQT3J5yZ2qsXCeLmIWW7/f
6+ij3woGoaOBfEGga44rmMIQC1LF7BX8f7RSw6vFZWbkX0i0wRboeZPZ2wyrxRfjfnQKm37fO7AX
Qxo7hTPLuRL0X3u9YR/AFLaPW3ejfzp3hP/mf05WCC2P5+XJZLGqxnMLblu3moRTItkUkLspa6Ke
Q2WFK9YAMiBaSyy4/jRaAqnwmSzSn405vRNWBjPoRedMRXQyJ+fZngC3pKBi0syazuWEkKZLuNXv
GZ61JRTnvp8sD1Cj/FcXsxGFe6QN47PWHOlS59iG8KDGcI5B05TeLa2iiG/vnbaVUDQftZxOg0mV
Rz3hH7/ViZO6w4K2rPKNp4r6B7NrvyBzc/rQDKWXwgd8VWUX3xpAbix3ue6trDIFJEo7PBKMcixy
YkcW3+rWx16lUtSgUFF3Xnqh8tzpt9bzVpoLAf2W2icw3gEj68oMW0ZY+4kvoKRuhcWXhIbrbFpd
H+toCO52TYSwEKAbQIlgxOCFqUlxbYMyP+AGawvhqRYRkGENUWvZovXdiYPgWoVmELyPX7Nf5zMU
ldkqQ77s8ocrGp6kMsXnFEd4L5nGLnQcV9nnGOY491/1A/7Uu2qIyiV+FJnnXEFz/rUOKUI5Qn7p
qeiCS0tADXk3kG3ijYTpp0U0whI5KavMq0PS2T64N9JJ2ydAZe9Y4etURzNxbR95GQ4Ohg5vaXDb
qreDZ1841hROM09DM9orhoQgubIenGq9DIAsVUKibJzg+Q4jRaBPPizucEASS6SkQZUthWgJVeam
a7IszdsUrgp86MO1WC735iQ5Fxux8plaRqVqtiJGAsIk9W/RTggtPSNfYSnLxfDITXtwxttAkOiZ
93jRme41I+vrQI8iTimprkWihHRiE4lHhgzG0/x98hsl1j6c0D/8dDJZkysW+HbyBPubBx/Bbv6u
GEQJZAo3abSYOGJT5wlB+fjTdvT5H1skCuSkITdSnWznPyjh6DD9vmPVAaDNjV18nNGQIUOYWWwI
SAYvjQXZjDemH8bhL5hlZJuXEkmx2AkV5hgCiRNUEB2qFfjQvBNgpRtYWkc35FYoKyZoZQEH+d61
eT5JKWQyh2HQ3xCmXT0kHE3XbR/vM3lo0/sBEKQ/AkehT5PqPzfyrXAXpuYuzPMTYdvG5FWVwQgp
Qc7t8BOjBqT5PzcKAdDmgkoWkS3dIew6MrzXm5LofDrM8xaolx7agOM9xK/CeBtzsQSMkk2xEpdQ
qsOa+BFHUKTEI298JWrzNXvmYUZQKwd04/BqDiQGyw/SV31LkR0NAbVlKYCvcUH/afWqkBY1ooSk
s/XJ6ak8Wc2Dx8OmSOkFUw5Tiy0YTdCw7kh5RN7XxyrmpxqjiL72Yy6SIadbEcTxJsmr3CNrvMpf
LfZQyDA0sHGn72DDHFz8YawH7SggMi57oC6aOZowQG4JkiZIyiBQlLq55UZK5xQk+8+4ZOeg0Mbk
9swXv4CTwJM15cb0eBZS3Wi5sAg0DI2e6ka9maCN3s82CEWAOKb22SLlQuN6xZLEyA45xo02UL0P
HywkMaBGPyuzQBHuJFqy59J2lqdYVFmNgnN4Q3OYqjDd4QKeaM8bJlg3pS6y5TlR+nbFyO8AUNLK
cZ2R98bHLLYKYktq/cMYrbQCzbCgAUcPZNwWk2MhnNZDi8lmMzOjtPOWNZw7vOHum6Enqn+xaCWg
kpSxAXDBaEJ6ZD+Um2u8mnzisU2kv7ROt276mkELFZZD0pRiiH9fuh4JsZZvGY9dVLibkyg5ObH6
hj2NpVNnNGLMwgxHITgzjvz/C9yS1wp53xlsn8qJvFdKLqA7wDztz63u2LXScAxcZZu8psJrNP5P
2DQtPPGiJnvHb0CDslpK4tVXxY9kq2gFzoIty4ERDZbwJblQWx0f0MBFHAHYIRXdNUt5GjsGcsNE
S6e7CXDTmKex5nhpbyj7qVLpaADzdMPvx1gJq/gxh1Pmbsv7IGZdsZ1uH3Jmc04ru3EUqev3sAyT
o6E+2faU9qfysllxLKAahJthD3OOooj8OCWrRrL4K3o7tZMhQY9FkLnJ3VYf8Af6kqyvjnPIMlrF
8d9xXEBqRPnisPQv3WbZ6O4Qm9mYv4tnrsBj0p7FFWRF7vAH91CJo7xhf2ZUM2p07y/rGQhoZ17s
UooWTsu/oHihvywUMqSdGOrXJYlvEM8oD/QzuMulc6pVOaz+tLQ8DnDoOrAj2Q5Z+AsCRHX4d/HI
F2pMQYMmlCSjhRk5VAdLmovdnKoyhlvvGC6vPTtdIatlob1Mjtzw+fTkCOJqaIgD3AnarNfQ8oC9
p9NocfTIwHjJ0EYqB5wVMhdzRdx7LrMhYKrxCGlkHFDyNIRAcvNRvtZAHj3A/NSp4J0TuRI7255x
QaGiNL9Rl+bBqDV4vIsN3v1NYNFuvBhAYBSRnqMn3fd66c5cQgFBatGoqwlkQFp3+xpbKz9956gx
80eXFJcURkJooRBjj8hq0AVdX7OVDbMLc9YlZVTA5Pr8Lfsl5IfTsh3ncd/+b+xU1hGgWI/VZDS4
2YmlUz5x6xoI4yWcRt7Z7oBr4s5Q0Z8jVgghvPkftkqqHZPIZeG26jwnfJAximEqcxJd+drn/Cw5
NNKDByIxyfLSBnGNnkZtc6+9M015BlbTP8ARNB5DRB7Hjaps1gWjQVXNbxkn53O44+RbsAvtg2/N
SUsCxfW4OqG2ndlYTSNB8QNlYB3ih6EYrJXS5wbojabzdIH6b6ieTCOQBYHMZ74BhdXTivDnYcH/
Q5cBY3IAhrNnBV+Y92VW4I8M/FH0zABAMZ0xk9jNwg8cMbUmkAV0QjJcQCe495mqXWDtXdBOjPy1
/3YhNH7cGN7xsxPLAsHPyWcMq41BdoFX46KFMRG4j9jJdQXyzuqa+NgfsFltNg6B/s8J8h1c7HKY
nD02d0Cn540odElpGl8l1YonycD3/ChRCigU3BhQ31RCEKa9DkqEtcjKavcJhcBKt83/+/FKtDnX
KVK1yH2k5TqQh+gdzK/s3HXReyQqh2TLTFGEaQKx+xQl00sz5E/MwdLLvkL/QVi5hxkeT9DAwBm0
JjleY8/TDfolg33NpH9+Magzn7G7WhXInVDkR5O7e/yyh24wpflPvqPcHSO1WTqrO7p2FAi0kwy9
Dx+iDT+06AhL3bcWfBf/IW/xWDiX2TACZbRGpZgWis9pKsi4JkAN44gOMzyJO/DAkFVbqrZt7neT
1MTU9DZ1w33HCA6sgxT4PUhesfqkKjFMMBxYnQyT00fHF1W4mSj54KxHZpjLZuPhoQreD4skVbXW
8pl7An9pbXMQ8fhcXp2BL6WCWfUoXd2LxheTuwyzrFj1YIzZeFwjQmpOxiurEcmG/M4BW3J4gg/c
QaLGcizBDMpUDvE0U4Mu+CZV7j0L/Hcaz0EfxN9+0bRfboCK2kYXvA/mkV6fb+C3dTXtPnsXBdPI
YgRLPUlb43ZRLv7q0aflMkPhNDKk7fP827oi7RFUPv//1q1+lvZ2ino6vPvbbIhByPcwJVYR4irt
JY0iDsEmjtAh3DiDxoFC+ItRCGBank93bgectFrAzRC6HbHJnoH7BKxcSvjBsTdPSQHAfRbuGOX5
uKZMjbvenzv15i+3tzrRlj3fhJxblEKYVkG+qk/S7eBQ5LSL6Gqtv4VejwgK7hZHr0b86Wwn34hf
uzZOcnXYfm6Pme6p06oN+uwCGvPvYUVwx7UT4Q0JrmjNjZYp1RJTgw/KRqLmfZtWSb/DlbNx76oZ
INmpXQXqhXCHv0z8pFASJ5K98seclOJ0y0PK/jym/8Tzb77Kw90JItnzmNMUd1CJzdFC7++u0jI0
VHA3y0v2/sLTl/FrFGSKUojVKnI3xdtw04lNRKofj1oQXDfmszsHTu0o/6QgRrT6laM2DaLKUYAk
KHyuKY/WjzeskLwer2NYal2CA5/TRnE+GmYWBvupbMgtkqB8ZsL5SJAxUrVeRttJNC6gLs4pnd9W
492bpRI9A3gkd0KO28o5BB/HvB9FquDMwXm/oybMybCjbaYmSpXBKFWN5bFaa8hIk1JFyJ+e+sQP
LL7wtJ8Xh6iQ3WOusxkhjsb5VJYLCOmk93DkeWrY5fyAGG+aTyJQnWZ7+q1LY9Ae1LLzK2HgeKGa
fEHlPybP6MV72T+bd/Ikn2F10+v0h3MhQORk//fsomlvJLQyZ7cD/dRwT12Y5flPOXMA2XS4+yei
8rMKowsWUo2tvHFTXUXhGJz/vvSQ7CYsUEtvrOV1ebfex7oD30HUy4magHQDaJrJlqAsxVeGt/sz
9Gr8ZWDpoMrtSkKv5GgRVwEAfIKiPzadUXzfTo3oUWDMNEExOOKoUhqM1hYQTLKE2e3OU1igkuzv
hbDMSt2Ju0XlA483E1LiZFOMUk7CQEDmoFDmNPpBmJ13VOVTovJu0wkIk7OMK8nQhVjonjgMizsw
f0v3Y+Oqsgiwg+ILTFz0O6ROk/2DLQQ6CisiNjxL80eJ4XIUK/3NCytg01n8TDk9E/sN28UgQGEG
0ivm+dJ/l1OMxXNDuk4uHlB79GGJ7PmLobzfzeDLxY5w+1NZ28qEMxRQ6mYTWCy99K9vvXGTf6Nm
/Or8QXvHND0c0tw8LQTrUvItVGLHpo3mAa7cnZmxS/bXuMrlm3ivc9Ew7OkU80ClnKzCW3StDkkP
lTOtmh8wb3byG/FDc+0srEviVuI4R69onveoDVNscMzAup9eYPIbw3C822aygu+ZT1bcNKxNEjsx
TRVUWfV8Xv1hLxjnERrZjkLYZLF1ZuFsblDHVw8CaHIQ5TNd0kGLhF2OFW1gad7u/bGeVoRl57A0
tkzEgHcjZLunZjQ+ogRJQBeGFXYa+KZhfdqeuzCVRMFuclnS/hHdf5EjFjEQlzXl6aAg3CjwjvZP
abK3+2wcHyfOKEgnkyefvuxwlnEPppV5low4hQyCOgzYAoqp7QrWF/TFulPHktI955sAIIqloa35
G8yQuqSNYHtp9B/MJLXpBYJWiMHjK5PiMak4Oa0xG8dXUpWSY9V0oKWeJqjwSFYHfx6EqFY33MTn
zqgPhQNdAEyi12l3q3dziXZb/VAIaO1Tbv3nX1sx4/N+y7g6Axy6vZ3I0KHTZULG/MEoh6rhgMK4
DUOvIEz4y0q+ZxYbisx3EhYJ1URyBSaJxO46yfzJH4IFpdSZp7xorexEdcfz691b86Q2IJabAx/c
uqQT32qFtakHqqh5OEZrJqY9SH/1uGiZzatPWpLWpBWQcqC5ORLrVkZB2dubwnt1qlQTYRgZkvaT
BT8irFz9hXqCpITE0hu1FfI9pETKgRxF8645skx5VLMT6mo0eq//xgHt2sandtd7KjGFpxzk3Z3q
hjn/xllS8VipuVg9ASUX/kv4qPOzr6ckH/XMdFrbg7gH6/wFCg08BHUDbHnZ07qQqdIOh35ZZ0ZW
mlPoarNy96kTcSdc8+6Ggy7eNxCY4olOjOwHU0BKiWjz/ywEnvBUh7xncm37jzux4ZeNVL3hyw4x
lDxx5Ilq/h4X1M+W+jfNrmkyvG5Fjrulw3NdGnj5pWAXFjzg/nYA/Pf5q5h0QXBHUFAJTG0md1UJ
Qukujh2+k8m+G37XIGxKENKlQgiTm4M5oIcocczhdG6qbnuoLQe28StLuBHAdzg0tTTFLWgpVxsj
DUlYm7C31lTE1isQngUEZHgtR2qGwhI6XH4bXmPm7g1j2diYDGkWdz4VDno+8i8bF1Nf4stfH0Qc
NZEQbP+CE9n6T7DCkwliiIbToqmw5wGjvE0wfjZRXEtEMJJ8MZVEztTG8DfRTOEZ6e2gk5z75wsr
tOUcUCzXP7NlZ9l639uiZpCYhGhJbN2lv2G6pfOQvflRMOidy2+6aQwRBJNb+g/CNeI3KCZcHz20
RdVMPxzJdw8drRLwyi3IESJs6yiu3BTM3t4Md0YfxDvjv7XJ76WLUfPbRpM1japeRWKlUI3w13+q
eI//2CW3Vv6vrmXPMwf9NL1dWC5slH1JJfGZpvWlRPKO1Bv8Bam1gpCk0CnfTavh7Q3oAg+6JS/h
azbblGFwCAiKS6TrsBcqHnBkYtNyo3TVMnbKBmCq4X5O8y0zhSsfxwnSON5UUju4S77wx2wJxnJ9
PFlhrTOnRa8OCVS4fkOU9+eQ7JTu8FNnWFIyKBBIkExq++ohNEGeVCXCJtEOWs3rB5kU0vZQyLGM
UUUHhY6qVH2gXHCSLxrZlANRo96UBAqIqb4DmHcxv+56fJR4wSCh0hmYJOa5s7RaBePf5K3odvNx
LrfmWglggCv0b/6ZAO6VAgoaGait5k89kKm1tqOxUC9SDEz1E3CvrJinb1N2CP3vOykmUf7GLT9H
VkpMq7bfR3xdk/DlDjuRMobqMZiVbmj0Vfy3n8vtGOiFHazOvGT4fCkirVbE7ibY3guYe0RaBDbX
txtXR0b2TjKitXduB1AzjlwmUkB4czUwkItA5g+y9x4qCpgXCbnp+z4Cbx3K4rjZaDyX2ezF8260
lNlYAMHRTbi2ydnS/2tnCAO6xZIhLqbMtDHMfH1MBn9d7LwLVQ7M6ijUbrGZOH7m2apJ025mg80A
9hHpZ63qCqBeEkwEBPcWNB/1lybG2cj2y9UfFB+N6Tnbvj6J1jXbDHMuuAeJezqXAhtF7f/Hx0Bp
900jl7ZunjEdz4Q4PuxFWo12NFzA/YrWtEp/HrPwmlNZZK/fN0Qr8AKqdV/1a8UeQwpYAM6HMLhT
vyKDFybDHARE9LxcC1ELtJxog2iGJUt9X9sDRuOVPoeA64WMSrsto107kmrsTYZEDgJ3kTjK8Uq/
fo53PADMI4vYwUg+Dz+KekjzhyrPrsqKkqAkzOVD1Oj7w1UDqrTWYTMCEmpHsViLyVUK6vn6Y4SZ
6GKrD1+fhwCovIsn0uHoky7TAPaLjziqXzlgd4mMvQ+o6oErtYyrOWsQpIsE4yrEkaQTpilZHo49
gve1kUoq6R80kF8VRTqVnmYP5VX3paimIki78cMeIGIzjJZioy74M1L8A3dOZgMxkwd6w5m9zkql
B2/RAiwWw7Uz0D4mz6EM+KNlezKzPxy05g1SS2YKMr26bdnGoXZXACs2GSAfyFGc5tQScGeb2pp/
T7tAyUNLfIzfPajntWVHG6K8E2Eos7JEUHaixipwsTDnVJPvnAV3XwkE/ht/N7BwYMn78qmweXwa
dHJphA9pkYRBp0g6xIX6s73/r15ki1jdTsV9si0hZw+Q3IrbuHfGANbHmsfKj+KEyRqHthPVG7AR
s4dox4KamB4EUeehykMda6S0lIIfpRcuE+XroN2cdMUPtqmfTF270QlmrYyaVFFCy5cGsGkkqiHh
42DoPFsxcJMN6zSEb+lmWzzAyyQ/rV09bQU7mG1B2ROZhDsVuZC3VQq5uXYmYiPI+b/MSO7mkjrM
RFFMfRv7FFxHk2lzK3t8O7hMD4rg+vvOXplUDYBOkLuO84I57gpyEGQnU4hWtfL0h9TTzLTjSEPZ
322xTr2FgbiUMn8TAXupbdWp6icZrzFRIuhwIheHeLYdNKjCydraPvFv1QNi4O5U8Kcf8Y0jZFbE
TxeMSmQtWmjZOdVvVzHlKcgmEsx+F2c8jjijABip9caGA7deslzGP1UCdbuh2CmbkVjAEPAQNbbb
Cg1/KSIGZF82IByRENjyCgwmhnfSJ5aSbjmQDw/en4LnZ7S7xS6oSo9vxZloKrwwKibmYbHASmnm
iSXez8+FdDLirpnk+CovbLwybXDHM3y4CXq5HUYmc63XRo8ZLmxkhcrxcw7joGAdISci5acVWsNC
6L8ZwPZ7VSCkFaHodBloEyA+yJ32rjCGoPG5R0z/CLg1BNJJeYMuzDJbjOlNXVvh0Cu4PAXuYOK7
abfepFNSCXkzqH1oEknjMW4zEMrD5X7HwlQ/VuN0YrAh1MMICvDwWdWs3IEZU0BcKG80kYTgTMHw
aWmeXxaLBYr4S+HDyZCIF3uxp4aLEf9C33y3/hFSnFk8fhzZcjvC9G12OyuNecsGtAXnN7AQ3NES
tZM3Gu575AGKBvUdr78qfb2T7cUS6ArxNUyXiZX6rQCFxzVBzbmykplVtELFyut4nCibDRBzEZPS
zsepEFLvi0vBBk/fUNc2OUGllSVEuXdHJqCouUbu7UOWt8iyhfXmGbAi/XAXnCZrnqXRfYWiH9uZ
2x4gPE9BV56xn9l20ivHslQbZm+tOkSE804Afa1fIKln0bgoqagHNMf4Sk4C66xBcsoJjuczqFuz
MLzGh5CHAGcZ+P9DGUfPvHIv5m/YSB4k77jS5eLgo+rM//1ASFqrVLPzB96iA0Exs+Zol75MYV43
kPG9jUTg1023Pz8MlhkuAM0RqB/u3GW8RNLRBMY7zn6WnJxMEffU8tcRDoH+5qSqwLIIlt6Kwf6F
S5k7pFwPpPzsMU2/i28QFtndRYJ+4wFkeIgAdStofItg7m7rpemzWPbbSEnoNNp5OioofO9n0l5S
gFLuwuG7xnfrSZQ6vFP5cJ7GsYn/kHHNfICxLZ6epYHM3ZYq2jpNrnFirNtKTUX5l8fG31dnb2AF
bYUmlMFbFhdb+mRUJ1bVDtqSQwIA4JiKHOSyqN27DNtrDF2JOtV+w7q8XHMHqv24e+E9dU3UhlXC
lLWNE68lg/TT5JWL7HebC5ZtjSGBzpOuylKhFVDa/8ZoQ6mmGMxDztAEDMHuA1dokcBs5couD0xH
Sxd5Lg3CNBhunQy7+un4W/PDv5IThtJhD2ePyZkrSk7IhqIKR6uNvKm6u/av4EZVFsVC97dQGwUY
JxEZVHbcOeQrlCtOyyxqKbue7ijcVdX7W9d9USb6RkbufhHDq6bV2n2D5GUYyKvrzzbn5eRhAGQ0
3/bZZ+ycMKcMu0O7LrXSSUgi6XZnveP9j7qCojjU62Nz/DAoZvgOwK1EzVR4aP2PRGdtrvyFRah1
d6/j1bdHCzZJxmDnlw5y1+iGGZnCChsutC52zVhLodcioiK8t/uaAzXMnYL4cSDc8E+O3K9aV9XB
IEGjYAIc/1958SYb+7Y5GPibHCx34egUS5Hwwm+eJ/fGuJ105NzCU2IV1ifICjW8Nx+5GQhMOX+L
tfOCJ8ReoQXkyH3965jU+GXCM6Y07Z+8KmvueI8+RyN9yRD5Bp6v//m0NbbK3RK/K3bJteyaY1Z1
OfOP2QOlXiaeO1MxjA+QHEcSBZNtYSQkjZFD50s7lQ4sWWNDcVYJpK4aR37iVK9yVwkjaAieUXXU
NPQyrXpkoItcLwnQB1bbuCmx/fjlpMirDswvlQcHIpCrmMDQ+OqYd7XFaYZpeLsPfxHXr0jJn82v
DzytWp/IveX59sLcF3DmR4HaeI8L6gVoD4CW97C3hsktifJOfhNyTeRty78tRsua6tqOklh4lXwc
g8tlBo2wonWlWfXHwdeAyfHUvZmdQfOs5eqoZcNFWj38eGi1UEkzQj+U4HhxVIj+bhkLaFy4DZLa
c3KqOsaQJYDgeX0RdX3gdCFceD/JGn5IAk40UdiEhCR1sv34thLMMwXxMV/UlzdfQEDjZrhp75Tw
XtQ3VCmwlzVXUIIi3InASOEbrMGQQK1JBgvh57W3JXkZWwoNxaNAlT5tN04ryfAUUYPoy0fN289z
d7aZnja19MRBNzGBM5oPmLlb9quEaeF05Zi5eHqrHsiLcO+p0SpNm0wMUyEe+N3IHM2cLnClnohC
WPD0I9bNxnZI2WRGaov194LXW6ybNt2NrB/Ez7QrxVYQyqhLhrtXGUqVqiXSS/ZrenWw/O0bVkmi
f1iiXZxIcRpI4zotcR+TwpfnDQCxsD9ITEJ/G5yXOJ9IE2sfzZDKBtGy5pSH/wen65T/CHhx2VLa
jeTwt3wYodtde8cN9NTBO8FRy6VC6ntiZnfpv1l103zYaYwZPG8CuqZXfIMBoiYw1goF/FWBjd/D
TKPGBUKXfOF+Gc3rEfA5HcotgSf0G/wBf4NwFyRFeKlDv8uDA52LiWqN9BnYBYGipqgwt6Q5/gZy
n/n54A7Km5HbWQTNWxQJVCjZTfqbyqlVngCUMIQTujZrwmS73WRhllv0bu/ojsTTTULN94o9bQPB
khxZHbTyOyB3whLB/GmYrbcCUP/fOW4gmMuEdHQOUaafPH5d057C1uvwhPBPtEPqCPosGblU4762
PnFh4oo/4NCvuZlG+gBNw/zcKEBN4xpjQQvGhVb04dbiuHK0MGcu6sx1o3AE6Sex0QDKqt6Q/sru
/KZlN/hOzOqraWFCH+ZXaIsgBVR1XcTj1dOFuv3WjVJvpTb08SWY8H8KRyuo2qgRPLXRIFOmlUy2
uA29OyFHGRtrTGFCJcB6NJtRMuGvRqFtCBkzWos0N7NdZHiUVorkmnDWkUKaEEF0H2hGE+w6MQDa
9pPPF1fP6VpCxlZW/IR5wj2fOfItUPYZW2zPFxNn2Ypw1b73v2calQdYCg1dWvmIjVhswKT57UJx
9enEuf6eiL7rfMbfgNvcWjpsz7WnqHjA0aEZgfViz4E8hDmKBmZ/JUsnUEjUO++dPq/M6fA6v1th
a62vvM5vSbLVjZuw44nk4El62MjazA+VoyS8qVBREmElMQZWK54MSNTuEhUwf6J6oKO0EoL0lLpn
OV/SXOoWHAnk/SJ7xUXoNQpjechO+hFCTYu1L1X2/vkEYhMXi4D8o0eMIoi2Bf/nuGveYT7li/jI
YYhBPAIhGBV/xxEI85bhgNvmXGy/l7BVc+5mqH12RYX+o3j3q0xyQ/uu4p53KWLEgikEItrrqBFX
iFVuVKJTV6YAkjTUuhwAaBxwqVOmRpVELhp1a0Ve1t8zB7c+bGLcAjkp2gnyLO2QSS8oFWsZyQkE
Nn+CtevYP6ZsaDiyO+YejCn0JB+/a8kIE6grkP80yQMlADL6as2bNLKkuHaXSGhGVOn6d6xPHpJn
fz1O6P5TkGxQBq3QlS4ta8itpkgjuHbLutEQFRqIQbeiEPRxJ90kCgPZWqimDMnrSs6cdabipC3k
UYO6oOagH34WcfcSsm7Xvttzh8BhnQjKxkzETjrCgrB1tKLSOHxIVhW9oeHOz6Z2ZT+QoxwEQ9oT
VgQW9l+1ln4f8c8TCHTnYzFRgALd2sqLDOE/AU8oJ85sykuK9tEbYkKwElWcMLEW+Vfowd8k7tBS
M0r7C9cC/MbG25e90WR0+Ns/du8EiSb6XN6RcNopOSqcRET1R5yCgJJwDWQLgycjNfKbR2l6eCLT
U6BuUl1A9cB0RyvhnZafP0z7d7Ib6ZGTwKNrKYKJkU/SvViqWr4/Aq3iyHkLOF51Dnqe1W5c6p0c
etSCtnLWPwwD5ncJavHcX5eXU3IC+cp/xXneTtjgXovYnPxozIlc6ns9OjmIX8yowwHlA7eefgiM
erQqGVM4LypXl6W5P66bWSw77TwRYrNeZ42Pg/bhtdwhNPDQXqJru8wZ3S/O6g3p0/0Dfk8Rjbmm
MICKvxAmAmoxqFd37bEP7WvhiYgD+ohGyy15+QoBwoV6nVUS9Bq5M7z2gTz6Kcu0GftSc2vxUqw/
ddWO27zgy2HqfQgrawpSTtFjtpm1jRJ7QKCYk2H23Yb/Xb12u/vj8dxwpZMs5bwwvGo3L/+B0JiJ
U4wIV1ns3Am4H+lZniadEcHVL/NuCeiWS7PVwK/nKXj37accYTzT9A8+vzIF+dvR8zNLar6WLZls
3ebgRUPkURXLebv4kIC0vDxmHJAcpwUHk2E6RlE7nlLlK+EPpMncnM+lE5L2QR7PMgCep3tvZJtB
qEJETOkQb4vNfnpCD/pH3pzwtioup3T0G87YCvXMG1VxM4QPrXlSWRH2w+k0/FB+EOmdMzvVRic3
RBcUwbB2ntALZs+Ii27xmStpK4R8zlsmaYVstS/lMH7Ruv1Oo2Gb7GEyYmtKqzEHG/s6bHavkKmc
64ZOc8FPdOVb9+P7ENXc0ycUcJfK9vPPJpGpLsBhDbumvwP0TyWDx7adMgxh89RbvWh2ROwoXVQ9
vRPM3JUu6pv0YLmHTC+EYYBD0wYjrZrv88SyQJGOTp+GrEJsgBQatGVa6oTV4KV+T9SgnWW/WCii
+Jg1g6EzaSnXRKudJF3J3uQtsByS2fhqJgdJVXJrXvyV2FiWmauicBsTvhbI9+CKvc0drw6b+vMO
EsET1+ZTKtD6fF5IPFAwlx5OOv3eefc+QFCvv5ReOL9UZCIhlfg4hAcBnBpDSAlOoY4hGeo9kr+s
IHZUsCscSGY5ksQEjdlEnS8JsZyl484rpNpakb4GNCnHpWcvVOdOsy5AGtCdOnQQ3fSHmdB9g+W7
vf5Cji7PxGQf1p+Ppi8cJ8e/mci/+dsPQy++MWzBb4dKHj5H4UDeKZ68ZmZ3YxvSwhILRjKqt00X
ucgZfSc4/77shCleypztYExwAAREeZIzYwZFvcNhd273eivF2A2wPtz/3Pgpd+r0QlQyGFbA8fim
OnXzCzdvgE+1iWlBK7+JUR/2hRsU1JoUdnbN6ZF852FexJSNBn1+0WexjpH8NJ76FPHDee/tBery
aMbOi34fcD4E7AasAj9RC/8iKfXZmp6XaTF7cM1HAOI3jZxJEuuC4burYe3PIoiRjByVA5VHvv5h
5f/8dFjlSyoNsyOtL/7PFiMsB4C7B/DAr6HZ6CtJQaYlo1ug985V3w46IqXX+/oa4OGyzwi7H8st
il0EB2pNwrttyuIJfag3LBdBWTHSnEA71yaaitgBLRYjE8Ew0/LN+MssrU9O2mrzCeeaXNjWC7YW
2PHI/fUg0bdGwPrvf76mUwPkUZdYXbYbERX26uv9DWqiVfygxIqH/fDJeV27xy58+qaod6PHKKtX
j+3QCHYSh/SOiAUYefoFovO3rTrHm0QGxK3DuCorrN/xJPwR8bvcEGeRiiFCWZljd6mok66dwZhj
UraVxYU1KCIywSdCZveAMef0eaxgIOi5x0rcEURPYTVYvIpXZnhzPuxPeBUUZ+DXjMyW8L1QkHMI
Jh8alKjzwBV7rENqFIcKutgKfjjxRbyQehpZFg20YAMvPefas+WtOGDt+um3em9LyEbGChJorSIl
drMbLfcqwHeqQI7Uei8n/OeUGuuFsBaMhtADwwxZIWmMggmSEsuWBIAz6h/g3bFykTdlYUGYFk2u
b/a/B4ehYzaFd5STmvIAtX36R4z2h4QHxB2vabbrQfgu04fx9qV/1/Dx7U13z+FoaY/gXsBHhcvG
iA5dqVdhifEatpRn1AxSP9gSmXUGroqpRoODLMHbQwCb+FT98gwTg73Z9QnazwfKOlQkQoFPRp9a
Y1APPzOpjIege1jFRZP2+ymxC9ylhn21bTOxyxgpJkAR2Y5l6F/DizOzbYzj11Nf8f5i28tzRQLz
kIr4Vhtz7fx9N8mLaxqQG9IdV79A9HtqXPE08dVG+B1YDaODOj3ry7MGyBRGJ3dZsFjLI/e2u6vK
hYk1YkiGnImVWvxziTYfL6YNVnGxqHyf5CO7OIwHUC43VnwWGaw3EjZPMW6B2jXvu/oVo2v9udzI
5zLQMm54JD52RWWyM/mmRvGv1+IgFYglC5uoArNU2ykVnZbya4E45m/9vrJ1Q/q0l3i7Rw6jwP0S
/zri31Udysg2L10TH+9Zt1Qw7Fv/jDSjWP1Uqr95AJ4zfLRE3oOT3mS4eR4hzPC80qtey6wcQUPw
7ZoxrWmJ9ULzNb91f6ysr2y3yFF4OjsYK4tqTGKnzVWPwXb655cox/3U/fbw43aO19Q4tJ6VU3zo
Ofc600ym8KCOrX0pEvxULcL6TLetFdQPdWEPdCTt2Ryb3Fsf+OJI5ZBwpVMA/8gJD5E+4KIr8CJM
G7HO6eyEutMR2j+tNrKTA0MGgU9eo/y8U7Z0n+aOu+QIema8iYjlTCEKcjWguD0pvu9fZtt1oiPF
eq/iBqkbPKZe58QiTlmTQvFqcsiCSZ/sPf3kPP1cdjSDFZtA/DEv7IQfuF4tNTzsktZmECPGmPlg
ioPj/l6gchgAfngDhIkunTfM3RTOJnnFRMWsOD5sqsoynIIS98bwGGRHadFDsmw3uXjug9GNsdGk
ung9BCYkTDcXTAhkayFXjuSzE1ALYcdhhTVks2P+q/U8Tm15oUyFEphXgIJENu+bVXtrbCqygh0V
n24LD9P6lhtbIV2GmMNs9x2wkgXoaIm7I+DLFAXZBmOAayIDl9dOUdy6l1gxje225qPFGhtjXPQ8
9D/yTwlGL3rIdJzhXuXNYmCjI6sLbE1ID43VcpUSbvqocsrRjVE0h7gSbtHEM+Hd4zDCqaVs5M72
Dd7DREB67jVk7q6oCFreKXX4G1BYg6q1zWm8XP729G7+4q5zrrlGpHZ92clUF5O/u1tQ5YNmBWVg
iX++/2Yg20VMi3ktZTKnGJqv3JClsGDt4raLbHafIrFHZixy0YH3+yuPYwWlhnufcSx508qRzXhO
z//rDEvRnKQdE1ZP2apvPDd389HE0UicH8cM7e3/QPhOSOsDppYXyKLxcw9l17x5oszvPJirAjIw
Wk97qlER5zzJn6jw4T7YtDBSL4kCsB+nOkh/iyYIay1D4NX/CVrlapne/M6ejpqiFqukuLEq1qf/
hmA2orPVnVO8cMquIIdnabaZTrxe3iSh9cTrLLyMw3bzh3HQCGw3rahjbOaJ0pfOVfTfdG6ds9Z1
Cg8dQgPMiAK6xLy145TEQDRW6ONG74CWGVZIYKm3qpLlYA9iQEZQExXFRNwlbt+WNrzsK1ia0Rft
nh+MUDANOJaPpzm/1R+vKN0NYU/iPE3xs+z3ArTPaVOI8qkszZwtW/SWFdkKVPlo+3ZbiBCvZYE7
yTW2z8epFOedt0Q7JMKHA7ED7QTygDC3n6nyALzL3J0FII1oFc1NGsKoco4Sfpg0S9j8ajeJQ+jH
cK0+IhHrU1ojqWQHAIvdReBr9n5sIMGW8Y2xDQ+kNol66QLskU/VDUQwlJTx6EImJmR+PCNJcf74
ywxNeneSYWKU13R5u+ZzjgyHmNZRPmcwvGhDp+cHbe/4EjbIaMQ+7neVsV4MHzGqeEDJDRtsK/uZ
6VfnTgXzNz5Y/ITicWRdbg1kSUYlGtdzgjMOvjQNihQx36vW1ZSLx+LkZbA9LT7KP5gGE/aaFsWr
dOriFbM3nHOL1QEp+Gdj4Aeuq3qkAKTzQXsTB6tkxIke0xITVhsxDP5Pwvt9VMK5dKkZmIb+SLHj
ygl20hGFa7WWlw0385wo5rwwEDkRBwZBFW7R6/RAgCMfqRtw//FyCZSL7ZusTGIP0qolD0933zWF
Zjlbjp7v8pTxvkbjYhlf636ohRdZ28sljflmXYBkeGNOLpjGKUqydCZNepuTQgVApF3JUyqWy44t
I2+E15kyQUrpNjiRlp3t5Z5xi1QhU65Ao6rkrQOCkOTrWAP0NLzzu+smUyL4UPVXyAuTg28y4Va2
UoVAo9Rru20/inT918b5BmUFDeaMZd1tNANypMIZesrXJplZoJzNwAGCcOL6go+Gx3QdQw/GlEr5
Jz3VbnOHKIXl5BR76gtIfW4d9/+2fLyGxT2DQT+nbaQkuHLUCnPVF1EMybqt94wnW2Ob3z7Cd4cp
h7j6rqNcmB1F4Y0gPexDRM568lqoxKYxK60306lC6FBM36JYUE0gMQAjGPoH2PD5LnNrcJ0QjXEp
GG8vg11c/LhCSoj2MUyULxZJrgpBuMVH7w/Ak/4JvIBg0XPKqxpnbmNQCsX8F1AjbfQ304+VKOIx
uh6hDCB3WmwWXXRU4DvK2Bi9W7L6N39PUBvNftzYeqlUEHJJmFE5HfC/90HuM8DVPYRedyBiacM7
/SSx8stxE66p7WplthT/DyZy7JBpqpB5T4yHrs1eMCMgP3MNpT74jN1q885BMP12s2A3QWPBwTqI
eRHC4gS4ymwhodmyrmmsghb8r59MpaQXzmI5V/blqpFvjLbpTjo60v2WXzjuyhoC3YgUkEcToVSs
viV9hg9lMGWoma/4CQSnfSiFZEdyC53Nt84YIIswNgRmCHhju42WyjMrrgfj2MxFzFWexVmmz3ZH
DmLR2nbCKsC9zU+aWv+UtFPkGoKMG/pXMnYmwNGoL9NbsMj+kCJOBq12Xkrq+az30G8AGHWCOwyX
LD5QkSacQ+JdS2/rW2ZjFijF/GhMn9J03TFbvfrO/eJ0RGc5PrmykgXn8i5t3+28uuS3W257qw+c
jL/7/Jn+cBQwgdeUN2nf4x9dJM/ndSFMHVdwtjfi8t8BZlXq/VCQ3YJfTfZ0YAWM3r9DQy8UxC1y
vAF+3cN1DRRc22aRrV51u06mYSfT8V7HWcDClKXbBN3Ez9DqZdQ+/qZ5w6dIhr8PssPBeRvjlFzn
FrdLtKg23qGWROhLQueZ8WNycajF7n97boPNqYdD/StCGSofM305/l8DzyizWVbBCmb3/QatkQpk
4q8yE2rr/+HX7qz6E3yOuq0mPcFU+BpAa6SLSCw1xs69SiNTqlcIz+c2WHm28T0hcOVMIi+gkgCr
y6lUNtn4pJxRWj/+yGGa7n5ddcYOr5hhFb8yTkJbRAHl/IaGF+LQSDaGDNEfXfQYuDI9bnUO0/+G
seJIiojdopU7YqEqLOL7d+hV8Gus8+05wjAtrwjuqHlUpNuurPki9P7hjhICz2NK71itXg0H5OkT
FOG7/125MmR/9GvF1/+QbpaB/1UT61fiRhdJ3nfPT1pWp4o9yF4wPm0M4pLvUDqSvaTkO+qhcdKW
KH9TLpSfVYnAeT5cHmNASUC0Hl7apGh8Q03tNrcnjE1KkiIr5EB8JTml5/p17O2JP6FRzOYBx87U
kJCph9bSkJLYDYhFMorFByxqDb1iOxrUT6o8h4b7wd0MKsu66eBiab5I4u8lwPu3cRQ+xGs5z9QM
kRfGPrNLM1Z2avp84vY2bfAB2QYharPGshZl/7c8NwKRfIpc1kMbjoz0Qq6wHCbWIbrjh0HhNKTg
yDGnZeR256bpTXJvCYo45lpgLV/iT1fvXwLOJfGbg+dYhVdGePinUtwsWRXC9j6yhhhSlwAagGj9
hu1aQ2kUh1slkDYWPd4yUZXebJk6L5ZPDHZgDAQqGcG8WC3xSMov/0vhQWX9xSdroKZVUHyQbd1t
KJqG7lwhsnxkP9ur601nwInC8Hn5Dw3pA9ccxr8+W1+vULY6p+UZwW50UBXu8mRiZorrW6K6gzrK
XusfyVTfrX+3Ly6CvGSZYyFsk7kBjSeIDmet3uflzhXpzLSVDf31tZZLW0HRgtRxdtQIAQIn/ORf
MmN801fn/hPieVZ0f5Lg42EhLiKMk6mKZHNNczcOGpxwYn0W7QmAFcIEXLpwi8J1V85wLdcdxCAz
PPMfrgZsp1Sd0n34GyTzQCknzsEUX9zB2awqbSbCP2XTOFe9qsiJWWooeLLfhPEiTI9itxJaCP/9
7eol40Hka+bzJMncH7G+TFcTIO+3S0mA94CQC3D2UvAJwph2Jatz6AEx3GfRu47oMEkc5fDtOmFg
DjVtMLCvZKAk322cvxhCHxrktnONwUv3neWFIZ6xq3oP/CCc9R+PW65DcpZz5Dfcv7lPIgGLFjdR
lfn6VD4lGOly9vN4y4MZiUsPuJwSRnEw8o2cYKu7Y8pxETQ0Daymiicnt0jAZef/HNnXLHR/WHRf
IU4/QiCV0/izbyzeeBpXsPWXPrjUYEVBwzTh3gNCBA4+8+YKAMtAvcvLkDkjYHy6z4CZmcSh0kpC
Pqf9mZjyjNkx3CO40pQBhUuqegplhIoMXe9lraOU4JQFpmYejjOjt072EJACL/Yr24EEzYh9DUYb
pjkrFH6duP4amTqw64oqSnN0JVy1xi4/nQXrKaBaGuRBCftgXUW899mrq3bP0y+m6+ConxnxkFpU
/CnV645ZMIpFYaz+RI++4EMLZmnWZ9X+SaA1KapBd/tuVw9rCS3P1X/5ZsUN0SNuxTLxxHI40Ko4
Uz41RjiMxgq8QoDFwT9pmquJZOqvcPaKdhG5zOUj3shNgku0+4z5pvh+/m4NdlH7uioHg89Oy1Ui
u/idapdVZSV4HzoAcAjOoLl2ssmtem0QYMfVOqb0Usavq4yU9DtNQPI0hpKVGrVvTKokUoOBV2wN
+YOaBbW/TuDIHSXtjAhEqkPQ4q+dhwcCy9CYv8Ns2TsnW4kYOjSsLidfNP3AKCuZtvL2LNn5hgxa
FwJ4kmEfGqSKvMJDw6zc/fpSplbVs8D43LChT8Oz5f9UUwjxfSJXXryXvBFWncQQzSCR2j33SFvi
5EnXwVyD7Wei9yKyMl/LfiUyItZzkgQ016TkPLImfxvJyQ8zgpngc7Fj4qVOI4drjOGFwLH4wSU+
ZBvIl7J1efePHSjnKLAO9IgYFIw0WCl81BoJzu+qtytDyaFRfNUoBRQVCiD5YgN36szdQfizem0s
ZIoeHZDnm2eYe/wDR4Nw+omeHr/UcizJiDAUntC8CT49oiMII/aWzYSoPd89YNBJNJUCRnx7oWII
1dE0YPyxcKn1X20kHbtCwOFc/DvaAkB4xvzUoT+frAWScihOrSwDJSSpZ8gh0lIaBgkLHpG0Wuy/
wQ8gSjaZfob8BlRRP0aHkcBHP8xVAf5g/td18E6S3HBMNgSPgM7OvsKtAfI9eLqYHtmM07zrPq2j
iVgHDIsYMPzMShxhN3Xy8DusyVIluCR9K9CNGSiooHGMXlJ0VFp22dWR1HTftE7TbkEs09t7BsP/
6wM0lMqxCkHg14TWAY/sRF0pO8Y8uFvbIqrdBtbqXaC+dGd/opjU2ssRdRZ1C1GhjUtWWQQ76spE
XFpZkUfXUBChb2JE1k6hrrZui3TEpi2vrZY0xu6KgxVHMhI8qlgU5v6gv5hQm6LnAVwawml3DWAh
Je02W6q+WnwiLUh+LACGO2s+YkB6+SuKJoo70BVS2BE4hCbCw98jurAcrIY05Vird6IK+oIe/jV7
vBPBSZHeXyq5EcxjqAji61scQqvb2pwId7JC6zcql0BlG0ovfEHLGlzLwBWaYNfV1lkqy2OLSZfP
ec9kvU4s+3Lbiy4x5SLy//lKGkW2auD1pdlQA67fUU6Jr1+VSG2YGT12f5oIwNUPMMTfsT1ulSSg
rkEAFdhYiCv94/igDef3k/pETbN/cIv/YMzU+ZVrY69VwGzhE/NSl3fJltw8a/CmXdk25yzuT6x+
Gyss1hM/7Z/gZVKO/09BeUMmg5FruXowJnZiLJ2TvVG/ldfizYwszZjw86Ly/9aI+4AggBwYZapd
bZY91rXD8+Ofx9yfgnlD+tBEva7VwuOzFbC3ngls/6b1APFv3pbtftmY6P6HIpXp9D8GPpi2SyTG
xBzMncFVjFQk/qpfKzcaYIHlJVrx5Cjcf0bWagzi5eeU93o7/z4Bow4QWkPwED+13+8Ew5kqJwXV
WIwj6H4C+YT3tfmTyVKfkxAZN4RWfLsHZrlFrbBCEEfXBuJDz4INUf92FN1RRmUWEqIVROXcNWEt
ddAnL3Ep4dT5nfOFoS+M3FBvOJdwoMbo1PML2wfICAYyR5gq/V3LZK9xhypag0XSPutLMOnQXd+v
MXBOZ8HW4PNLL2nNVYAIIZtAwrxvEu0o25cyi3+CyQ41+OEA3tGLhAid0djEi0Iz8lKNKp2IQaQB
KE2HzMBVIJfqtgK4sJ18VKxZKlXMTOBcX2j3K0mPOct+VpmnWV1nE7srp7kjj4c0ns70pCBwEAjj
E3tKa5qSzQtbhEsFI1XMyg3bznCVMW1AKJEbnxlp8QRDckJcDC/Jrcl4lPgZ/D5+Vn0tr5Y+VXjN
cUDKPNamTH4UnrJV4hT1/dOmAqxXGH8pxruZvLHxjTjWEKXrnS/5PuQLTBVlFLEBaMUZRpj0efep
vc5mPcdL8387JQN8U/artMCcTlxxClih/tNbYaEioLeD87osNsja13VxbWAwnK5aEebbHv1TtryV
xXa7Lrt2n0nY2eMARk2IC+fqh5rlND3reNU7nSVA5a+vRHWcd1IULPVrf0U6UF25vetkK3YmwVc6
ZlS3xuwklg8wQf5JuhDTNSWb8h4PJN+8PT6ZtOPK542/QOPE6a/aKhwgvzR+H2CaqwrPe0gpuadW
VCINfhJCZPkZsqJLiBLxBLJQyzoZOdLCZUlVLdcvMt7qGugJoRDfOVsAZSsr0VwHRfqr/nuYv/HL
WBxhOdigsxpAewaLQd74OOzhMAwg/EnMJdrSslR+7hOyMY1MWE6C+12ec37VnLzMYEGkVqR1W+tO
+jSOVGfPY1I1HfbBMZlOcJAu0D8H1QreW03akkSPSny5Bu5PPslNmxMRe3twTvFBipdxque+Ix4Q
kGcPfkZnbEw/PUh4F7jQDmz4yUCzi5nTnfZAaH2pyAAzfcuNX6zW75dCDaigegsxCRzr3aL8++mD
M6Q4oUY2Jv4x7PkQ/iW1Ox09yBTylhSKhqxHkUeGwOaFZKbXUhgU/7sMBs5WoUgBMOG0ez8em/Si
N3yYVOpy6C57nUP2agVmKNiiw8jZgLq0qQD0Z9+sOPoYXZ06BCz/zmiIwWsIbZGsEEjuYeoxcVI1
bPykeRLIUdSL8SHBBUd1VY1gfVyPlNTYUG4WObDrTCn4nkFVum/qSyx6Xu/JE/3OfssDkYQQ17bn
vrBFYQ4jozvd3pBtB7A1rmhWBVxpTF6T+F0RS2/1sOZjR/2c9gd5wU1PbtGnTLrq+04sJUbqq3XB
YjVPU92TA6SCAkEruR+KZVMOwEvXQrXHuYnWAtLlnShS1SWi41i0OoYwAUrSjAyx0UT7PiLIC+BW
gtpWI48zPAULneQ19P+uGOrNLTR3MqFpMgohkZ6b4uPa24CmJOtUNHtYvfxORpB4UaUrRtiOfiZN
r0SnhxNXXqzn5s2YeMM3dzOcZ76O+lI5Lh2VncnF75HRam9rtaFa4wibE6KxAsp5P3Y5LgAD6h50
HTlIc0eAVU2cf0xezA1bGpy0Co9m/Le8ogvReMQzKuuK1r+/HxVHbKeCoRH6w3aSNUaggL1VtIEv
wOIVyRikwt5eazHczNvvwHPDzWzvu7Q0M41JQ+OJfiKBNjA6eAeGC3LR91duszFuDeuGuhMtbN3n
n8cPnWstVCZp3g4UU1h5bJxMeASF5mFjq9WB5ufsPeRHWLbBIPgXAPWNx4m8FVcjKr39Z4P7UgSH
HqRyHyTUzUmmswt7W6Zrnb7Fhb4p7g9hMMCgLxJhc9sc9j0TaEMQYy+cYVz1rKcQArzdCiW+E6BB
3CoRPyqV6CLdvaaDcpellft/qIf3xynxr9MKdc1+egyw8bHlcl4nSxoVcUNUUMQ0EU6ctuQgAWvo
9khcQ67+ZmzMmGV1V0KDpTZreBnwxHmD0F1/ODq9gQOqu5lClyE5EU/JpMHJI9y6oN64FU43721K
YVNfJmD6YwO8kmPm22AhvDPsEdGX3t/LDLdD/UhVyzTL/xE/4XGU8Tg7VlqPLJLEfsBrqQTsjP2m
ytkoiJmYXE4o1rt8qQBud0S6FKlkj9+SYhx3qkrt8VK7wnSNSRs9kzxAY2dGkT1rtVIlj3SRQEHK
dQqb77tv33MXPzK4NXC1QsjCevZRJHpyqodUMunlZyxx2+DZn2mDRXrM4Ci9UKoqT73TPjx6xp7v
atTiHLuOx5/oAKv5PWZpqcgkYqjuRs6S4nYTTsHq8HtO98P4SOlfoZl//dWy+shS8LoQ13VOHRPc
I1cInMYDy30U0EtgYYUGFW/7vsMJOfbVnKfzRuJZy2WSNrW8CFEvJCfIZJAJQVu3zKNylmzsMTkk
5OgXndAVSTzrAxzhMIBnzNa7oxE7NCPBzyaMCmfAH2V1t4cT2+qhe0KhV2iynnV5imApEtWE6hZc
LQH31Bb9HGyDS1kucr2AF+nUtS/Pf0p0LPqUl0Uup5zbI0N9+qbgac8VCnHlWHe1cFCtKagNx1UB
InC0LNFOM6FUlk9qsNddUJyZ3mciumUjOziAdo4zg/rHQ41OOvuJmBLt1gpPEJ5yeY1umt7jQ9/+
B6zrHcFMRSb2uyWzFsPhln/CKJfqMfDPoGr5gDlvG6TETwSxoKYvnq2j96DmK7vW5NxC1ZnZz9mV
HkjAScEbSZOdIJ3tB8katsxYZw7f06hED5+1qbE1ovn/4Tz3tbYovv3+Tgf5c4LPHsyDXyvEJJwP
n0mRof/DckggE7z+MK6YNiX2vtWp9IO4dGU/Lqdoi7j6SqdC18U/JJtxaNi5upnrxB6xdHx8/DeY
gketwmnEs27V6O9OtxmJvKiab2+RkfxuoAt/jtj5sXr7R8SnuWhUfxADC1U64BOfnNgB8Xlpgar+
Iizl6HDaDEcdov0h72pc/IGtUlGjJ4az1X3lAeSwXPZUK0mzx9xwvUHpc/BuQMI/xqhL8C2f8KKT
nyqdhmf81oJDAAzYwnIAI0aUVi+ThQoSSr1ypuI6TT+8xEo1AhoSyJC7Nd+/s6bbA1cTvtnyPT9+
e4a3HMmkbCvGphkS6OLY7Za5G89Gt+f6HYsydZ0jtXG7JPEh/V2YRgWjucL6woib0E28UdEBav7v
RppIqGS3BK9fd1Kqtw2u8VBa78aA79khPLFEDPjIx/Rt/s5tXgSZhP9ho2QgGecN8CFOlu76SKpF
Nhd7V5QAivtVdhr4Qs6QhRPetU/OxHJ2YGzxG+SkejboDdvKBQVtiUM66TDAFhiuOY6E/eyqVJ2t
jPE2bMJzCUEdKxuzb5Log/wC9lYTrduVeZAO82wLSyatMiMBtNsStO9QKqiOTIseSBSjmyIbwbjM
+IJzYwD24t3oQ8xibQZacTtlgXqQ11AYpIVuMKvv7Phaqzg/8IGytfJNFXX/KF05g9JlFqNCExHJ
Wponx5Rrk7mTINXYWzq7O4uZCVdhX01eTH+mzDqaXix5dyIn+Y74RYvTC5vn1jcHesOB5kucKEsk
LI+mrG1/kY9H+CjPP2e/wskmXCPkwAxk/kRpBeV2qOEFQO+MRM6VNXTOHcde9f2uEOztXxVSgY6I
l2Itu1cqNrwOvOsNYMpjztrx3qhoqjWC9f+kvt9hUYnXyTdDoqsvsZl2yBOLCbdPZnphwhq1g/u3
rD7QWkxWPIy9bIQ7tNAlvHigXbpkBd8kxurrCZ+FwQhQqXu5LlAiZ8Ri+BWaVSD1OF2+czEgVK44
BuiAchChDz9YLVySzW/Ymp+PGhxWrQi3v1lUIKX3OE/QQEdihUZEiDtYaigkAKexoKxMLcs5aXfh
BiKm6ftAsTL81O+V2n0czejJT8aM5EAZuOFiRgsZ4qpGNXtuiv1NzfxWLJsA516X931jsC0Qkk1X
PMpuEE1IF/to6+JXfRo5pfvQxUQOrA097YywvJ/xTk0rTdtqMzGh1G/BNniAmr+0duxqkBeGuVs0
1tIA+8aADwFZloZRnL7emMmccuizdaQOjfzdLxv9WEC3uZ348mUZMdqxRwwuvf272agoC0vmXZpX
PJMXIBG/5XTqLK2EK4ep1/4j/XcSg/V5jwQNzPyQyI/hSG7AP4gdEeOKoPFOotQCWmjWnTNWbpzr
vaoHr6VLdCkaGpOtxJT7o/XuyJUeU52tqOFvgvZORxI+uywZpKQJw3vWgzQq6BCdeuysSJkGOZnb
b9wfwRNUxJIppGBDoYYWpn+uImXUPduOfqU4YKndWA3of8ADRx4kHDNEntA98uI8u/qIt1FpI+h6
L2r9N9ci7/X51TcWxGBCXeCmwK49XFcjd02LQt3ObC+ly7auoossdECaYdxiyaJ46g/m4i7c+a2k
s0ijgesrhTUWL6x8QR85pXxgCaG5AN/+PHPzOXqt5Ri8o48mU/5KofKhmG+hQ9GSqh/QsXNCmHt6
8AVrE76mlB3ALIa35sz15Jd/6OJdfZ1rP4duqYnRXRoH7eXDantAccjkEWg6696Qpmyaw/oxwDGZ
QldKP/nwMK795kZ4ycylzskcCQaCTKbWV0PlllNV+agBBT6XU2Xvf7A1UGKDt7ak7IF/CZ2OCpDU
iFoFNJwuq7H8On+p/PpPWe53zPH+AThUneWZoS8MvkfRMYwKYQuz05VMkv7A1ulaWREKyUiqNPoG
+rQLNl+XOI5GiTbTScDL2W1yuNZAOPcIOgOhqbPMDoNUo9+XpdkpgLz95Z00lr+/xLJ3iPNxFt2B
mDq0f4QZ8ilLBhtN2OsQvO5y7piwcBYLrQp8hN5h2VPg45rKqasnpJkBnnbZldxzLYmxbHbeYV0Y
3YW1XDL5E6RVnZiW6saEhKA64amCkWX2a/TZWPy7/unG7PFDao5tjeO1rlsj/a3BsZhbYXLY+7wo
s24q4pg2TlzUeQhqheAaPuK0Lq59KbwVQU1WhMThFBHkZi5e9z8hoU5c6/BfKTCtGhueVVh4Izdn
gtzysTq+5Sm0Q4cOeOoXbePSGPTsWC9gJi1tvQfvJjE3EvIb2ZpemKDdomJeqKY165C+wWBVCMva
wL/MkLAFDFfuDAkPCb+37GWEL9cGlcwvEkCxYNjT8xxvzLZdq5865RA8dZbD8kDW9Cg8tdgsZ8T8
WzmLKCwgzakHTMGoh4AFePnJvwET0Pq9u+qWpy1/FTmeRkWpzsB1/L5pVnWVQja+yzc9REZCXnXy
tg5zZYKUpL6BPLRtVulgi3mpsvwqWMJ1vwRMTqGzxwFDhG7X+bSDujYqqFxPxy0XtQO8Uh5QiT46
8zb7cC9N3xAs50/w5P8qOVoBo3jTbP0qH5t5MBv1LJVboeLao2ScW6hjoHn/zXeU8kUKIJHxr2mt
inZpI6E+sT0Q4qwIUEDfeT++y8I1o/bGxf4QzYedQPiD3XbllZSD70txJmLWOVhN+s0ZSrQVZeJ/
4LXvc+sm4w8In6lMyoyF0EqW9gRgSTA9M/10WMGf2I7I0QqSDK0kazUugIRlB4WpMclS41txr7x4
FWHDJ2GQDY3zw6m+1+BDBASaGQ91Hfmuuoew3H6PrfAcALWPsqc81CgOJt3l3dJw9CFUJDbxZDUG
d+xatVQRg0EbSNeTLh+6dResNfwRIQwS4mp+up+pyYa9dVcjxcTtILhIowTY0sQF7B3yn7cBY5Tw
o2JL7lCTBBcZ6EKwUVEZ1gCPdqkScOlTHRBpMJRIIjXJVDxjrxDwT+Aak3lWYbnyewB2AeMge6on
ykba5+hg+eIeBFWCjWwy8t6PejltTXZWHC8cjfbgjFl5y1dgFpzKeEpnbMvqErAh91IjHC8FlhHH
5d7xyaQSm8tgSdeW2bOxcuu957uU6bcCrdHuDGqo07KgzsNidmeYpBeq+O7DX0l8uxrUWxtpPSX8
o6yiUBBB4PnZt+8x/C93Q7F3Y81aw74U2io80fyZkfMcQvejcpMjw/31oOhNjxupb6Rx/FgK3Kwi
ZuvY0hFS+DYyzDPFB+ZGh+GnJSzU5dzes1/gu3PSkw+r7UXPBvv1oXcDTmtU3AXlML8CjVL2oADA
mzuaaMUChu5mQmuxrUTwUCho+VQGwJbTVzkys1u3wXkg677QmerZzCT+32v3vjxW40KaVMLIZE7C
ukjf5FTTSK/j10X24ePYnlnq9OMEBYEp0GPPWzFPNR20oEELGoa06g8AZcVYDAmlEpxeRO6ekrsu
LNeTCSN0sC1Wwulxg2uTf7YlPyV0G7xU4KIugNUIMHci0sD8Qok8SznntVSRLbeHczVXtg+7+rxz
hWhrOS0X5L8VT4RomWAAVi2nfbOLNXECnW+9OULt71db9LmTJOlSUPGrOwgZJwO967J7Vmlwniec
RDmQr0jjytw6H6bwKts+TfQrRsTcxgxNPB8w9GD47JrF+zuhSVxgqXH5+0Kvsq8tB2jMPMKqkQsv
Xp+G9JSkT77Ej0FeuWxtqZcAALIS+P7B6ON0hQtGfo+NYejQ1F65HrLUK7yXPKYTmoK4sj7ml1/E
f14G5U8awkqwdY+gYvEz9PmTEvy2rIpgD0QcOlWn22VbNu2OdvC6ESRHicZal5W/TyPjb97ExF5i
r98pjXuojJaF4kuDvFA/UFYWAXw7hatjso8QKoXg5xbsY95q5IDM4Lm7ojH3dYa1Ad2uwg2VVBEu
AIPHUgSFcXgG5X+MSCjKOHqAl1formLh5ecaJcJrVWyhnTEk7sRszpDpQtCwOvp9bxavjHkdQD72
BXj+HsQ7O218p0URbmI0Pecu8anrcY7pn7s85lFbXkhD0j/fjzSUMr0DRydORY46KyCADMiOdb+w
PrGPaz76r35yD2pLyzodGGHRuFg/MY8hOju6r0iUfLWY3GXW6eV8yqTeEHEXJqYwGa/GW1hCZFmI
+UEC3Cs1yOML/obCyjn8bE3dR2WMhLJzw5jz0vSBRW/wJBej1ttrMB8Ky6DRj7cBXtWrl2sn2QGj
UWGESkPvKXj2fLBG0ts1a6DlLp0ZjTYutYNsy10Wz0MOaOoVpaTjcxDgQ+kja3YMxuA9C9M9R6is
9v1UIrCmLXMCPYTqcuBWrT2kA0xWGOggEvJzOGkEE8fkt/ksF+wfkks7NMDz8cplRysBlnHLvkiH
0X1EWAAYry+08ZVN3tG/UYIQBA8tEpxqsu5o2xIt/etgWICO0vTMo3mxNXbKpLvzB+pwrrmLU70o
LOYXEaNo7QUbaH8wtGsfmDyq5ZoYmb1RXddpLJtBVO5Azv3c/C1D0F5Zh+14R9xx5im19JrTRxYR
0KHj7M+EtJm/VewugVnIP687aKIbAfqRU6UlVdQD/6K3pPYh5SLN3olO8QpXfhl6h4o78LWd6mho
VyCzCIudIc7Mtr3XTR92csc7yxcR0g98tlnnM7PES/srAB2zPrLsXubqhugXJvqG1+Mn4qxKmF4T
d+KjOd8xef87rxgLR2tLkvljg6rwZVtFRfc+5ekpX7co5HOy8TGT4rO92FwKOfwdDwD4IRwN/OCQ
2jhmZIZb88VhinRcTUNlpYVNVmVhZDobzP1s4kcBLjhkXyudNSVdSrHxKIzhPAxhjRStYFQTuIqi
pKtRZLz8Wc0oVwV6vzkmpgu6Yb81lLLOQKprwSOKkifLhKD2sQ42Gz6hmS2YPxd+vuxNhIqfYKSr
602hRnKQ0Cf2dgSNIBzbFawBffF1PPgOZdaIjwPrR/kIqx/QQRfKbE28EbaHty1HcuOiROrm5sXR
4+vz5aQjAdE9G9vW5zk/fK5tcDDpq1tH3bnfWEQl57qM/DjUiQNbqfQzgGFvOg7ayqQSE24f7FQF
TIHd+U2zRDDHbro44wcUqe5HOFgo3B8h+UzW1YaK2rz++5me0+mSXJ8wksYrNfzx70408qOHiC7U
VrKw6wpHyl4QvmjQ2M09TiUiaesTh5T1xds8iRl7U629caNK5xf7/PTgjangziTyi8r09VeVKmg6
9QNvHumghVeNB5eRPgL1U/5QPCpYs+ma67C2RZLEQMWmp3NZakV6vDTczkeXf/kwz2/wcASm+sap
WjM9+WsUyVlRneH3wNdl7ft11BastAVIv+AqJJWlE4fXEOAVcg05p3Jtenza+4JTU4Luc/+xu2Kf
IE0bBGwS3UYszcAHSUpAZjic8vJ3AFekvoLr2wg6RegV1CGdHecFSnSf9GCOyhcpGoRirAJVqmdo
NyhQdSkV98lkxe2iIUtlRRbTQPOqiOgEYCA5W89uS2fzl8WRsL3IqmoLO1Vlm9/usRhiBZLcCE7L
2k5j+1e57xzUD+XGWurG4CfzQfupzbF4+KXaAWMIpHUW262GmmUjEruUh5JY4l2frFuctWP4HcmT
0Pnd4Z1HtIeOwLibAef7qrJd7T/5sev6UYzflLFPOsBSL+cyzc324o6j4X0UWHgdTYHib+2C8fPJ
WMKVxfj4qTWUA8J1C7boPkw+FqsmO3MqbsbPvKQIiNIvbP4viPgxWWdk3KvsIersKFuFjf/Jt6w4
n2NmXXHhzFR5bTFUGbDWtuI/Ylu/DeYuAFNdbw1i62CPOgbJn1G0SFDxmAMganZDN8xW2FV7jENT
Zk16VF9edAn3e0RWePPYyCvUvuYPkxCRelIkBDdOaSnPRLsqU4jGdxRZOgsOxAWJsL9XOp2eqa9l
NfSAujq/Z5GnVf+M7mgZyI5QE0Jvbw5cAcTGOOeIhV9v5Vj4BR2QeUyY2aKyKL0FCoEdlj0JMdki
VUx18BegVUCdfSbS6dPjoKYifkCcd6kTF8V5ZDJ1OelAtLAxH01GjNftFFUzt4UDiqbZodMwqEK8
3IEDfI1W1vycqQ1Zm7PxddfjRFcCgifNdDD14nHT1JyPNDYdOuO2ViPniupIbgVx5JKTDwghHqYR
VZb+ik2MZnT62v6dhX9I8BdzTSMMSNCiB4wVPug9CHc72WgDqQXi6HBg94u/UeRXaV5y74Wl6p5y
ZXmCVCpDMFsKAiBpE6A1Y898Ud9KMDOcI22ZoPtiz68HXtWk3YDN4eHnIU+nsazoemjrDS3dSwNi
mnmHvS/ei3O47xroO5I4UyxZohZ9IEaYMhdEyBHke1d3v1YOMGFgBgozoWw2s3/Gq5yYdcUTdCDy
6l+65KSxNz+dS5wPp0bJOpaUz9VsB18wWH/gnWLLyzyOd+6XMXv90OOry1/baQ2GlwqpONE3EVDG
LVDxa7HZwnin64I5AkFPao5+naurqwjPm+jGYHNqEk+wppk2nfLukPPiFTRYkE85RO6ZCOOYpIfX
U7rZB84R74JWclDR1AoP9scCquW3r4yEAEtmgbsNx89TWbjLfJhpxwa3cj4JCP41QmpopapCALA3
HYGeHa6CXshKVL0YZDoLuPPcsBbGDVI3DGCXxSk9AS3yEGfknWgIbWy09Sxo1pOXIamF5FW3YzJ3
dn+vDtX0uaLljWVvbMLLmEyNNiyESh0tsc5H+Qq60/7Hp/QyJ7YrCz0+r4miZoeo+MWkOWWFDKfM
rlljBntjkJtETBP7G3GlZ2HuhpGEBJDVb82GEoKrT4oxjiKljVD1MMYI0ZpBxEg+ZA1svYDOW1fO
OeLlsnxCrUz8Ei4c9ml2EwVbBPtCl2LsbWrbf0EWfUH5BwsMmH/WtJUgwYH4CPCF8WFbHwkZUV6l
3tN9dS4cqHTLFqQr6qZLuLAjDRxWYRmMpClA5q8Zh895eYjTehedO2JxA1+Lw8mZWvdy3Z3WJnou
91NFeR39RudSRZjALffBfdguCZESG7fqeto1HlRXjRmtDLSmEnNV/0SKSJ/O1giDg81YALhbXY9b
bdDkVe4tleY0bV0bz+rwS+owrNk4dwEnSp+7njIWNmJ3ASBQiq3rI2CK84ceF8X36jMxyf/CvAV6
T1qMLoTIg7r/qGE/zgql4S6bfKzYrF2UIBRHejrz8V01UmPh/mbhBButanpVrPVATdEJL3oelKOm
wi98NijHGvIc7bFNE9qE8RofKsYQRtyX6HO9YOREkdbvS/inTJHP6cYJPzwovOI1HLYixhpyL6W/
Lldkde/T1wmzWXcfpy7VlS3oAV/OKn4b5cb7BW10Tusoazy4JtDpp+CCl130Jr+T2I60UPbvVxVw
hSSZGRQIrjDNcwFUtwfmatWI7HKZLX3nCOaH5KaJAeZulcvY+R8SGjl8/nCw4He1vcaQwOjm5enR
RK8nMRjx8i+XbA6geBkwOfhAYl1uqJ3jLpH6aj0ieWd0iAqL5K3s05lYemZsbYlMvNbcDAPThdUU
ju9sX/qQTytFhBErnQzuAVQOSdT9mR9nD6bJtrCvLv6yPtHG4XeNnFGeKQH1PTMECDO1AwnYwbVc
Lbfwe8Tj8ex/4z0PYVVWyw8Mh6LB/bZKWo8AC3B/a4KgtJQjngVcvdv7PZVD2jQKZuXC96FnDYNe
sLHNvz630YaE16r90cLy94Y1Fbyi/bLi5dyUKupTiYVlpWm0QapxlAovoy5I+pQt/zUXHqyJyEjA
CYuDqF7qP3FPAX15zUAJKQglaqZjhmS69rXcOwfehi0DWKtgK9sTP0f/h4uCVByqUAoKMO7Lh9KY
pUPlVc6TIB506lRDocqJTvk9v6nMTKF0rmHJnEYYGqgYCPqMLT+BLGLsYUbWqJ4YLVLBAxP42vuI
PyrVPcDG6vl3nUYoESqCzSmWM549W2bKUWLJv1mGd8Y+5vgicoxjH1UcqWTRqz/fu1pIZvVBhTTv
woLK2rUlZt3fru2ypaWkNXm4BuoFhTJ2vxGNH/p4duUVCcen3Ju3JcwbvOsHSDYxO3shXoOy1JGo
N0dpSSuPycVpBsha5daEoxxJzLCnzbC+W7zzyx+lr47K+RmyW1ZO1X+qILtobmcu2Uc4UrPCNM/m
misbh3NDZa3YIMW3ggxSSUwp2sUXYdH1WtIWizPp3v/P3h+a56QWx+LaPq6rycuu7LlUoXnmVLSS
8hebKgbl3HTu1IrX1X0cAa0RgUhkxmyWJxjroJYVQtVW6Yj5Qz/4X+VeDtwgPOetxVQRz2X75c4v
TwwPhUvVMhKakBz4CfYMd+8QwkzEunjxRN6W3xrKzYD56oAAPMoGmFtTjMo3P5r9KKf5LcUT3/VU
rQpO488Pc//YxAtHpF8dUrbfxUD0W9SgLQHs4HDNpeo7oSaAhHWTUBNjHxMd2Atz7L4c1k2MB9eb
yL4c+wU0icUbSkoZvy77WU5j7OTinLyKO6cqwwJo+u68hTDMqGRJ4ZYbjIQJ2vyR4W+d3PKoLNUu
4gKvkg4EFXcz2/ShSD5UfkYt5J4U++VorUkPwp/O+VYr81Dc51aPYCieBdvZZZV5juXB+iDo3HCA
9rm6sgHokXxU/5HGHdfgFHpXIKTONSUGSUSXtcEwox+dHsXLKXqDy73r2ro7nghXmBsr/kjztcAn
umrXk1hkPHq8umaajKDaC7Lbg41PIRm9LGp2NBxC/6aCJgAiQAuFVDV/DuU51562YrMk9hSDm03m
aCYXFlrGOaHmkntWC5wY/KhvxaNq8BqB1j5Ez3c5TdEYLiZeYlp67t37udcCnU3fj8EFHWSxCEXc
bpF3vVwUGakeJkBj8N+3b7q9LOM88VEgbvuPGzdbVU7XaWw5obvbcWCb1YxQbuCVh1wML6T7BBQu
jrHQMvP2S4lFM2wbbTX0LybA7Jg69hDSt/ELodA15vb7UWDoaWupFNowPqXeWyaVqR7tuK2XLXZm
ErTcCIWPn5GGb10b1VL0PYhqRGG8PXrs4kgBG7rf58aYDIwbtKOu/KpQ1rAiZAN3ntadV5TC+eib
HX6y3MykYB0zeHAODMcrGmN5J+nbCtR72W7Cd/wuc7sU+49JSunG2WCRXxdkm4KuUwZWhXD5VM1L
Fmn4U2AugXR96qDnUMYQZRTzn2Y2ASBc5B5d6gwLn421AnnDRcvLXEb/LAMRk5RUdKxtpuvIz+IJ
xxY/sJvB4NNz308mp19iaU5ELuMXriGIVfzdiG0onHUiC/qVSeoSKgO3+bYP2C4TdBLPZxdMSfLU
LKeai/hTQycUvw1m+xsqWXYNWfEyqZ5LMzw926LAT1Vs34k2FV+v/G68GbzV4g5cRFzDWmSX1lez
0LNnuujLASiJeUtRMIZ56EYTvEBVtQlWafcIxsYtTAwmOatYVzxW7WP7bPFQn1/YR8nTjN4P5VbY
DyK6K06Vm1MWiZ9hJkvcKbvnv4/ddfQs7ZLq4zA5Wer7aRatDWwk9Kv3s6Q0eH/vpa7RXRxo7ad3
46c2beEURUjcp44nwCrLR3YYWpIwYWKYh5E91375OPB90FoKOCxSOAN6iwonrXvsxRmktv5REtk9
Qr5BF9WylqYaklDzfCnPuagYlxP2GKXwZ5JPDJ21XmTqnavTBpYAmKzOZmpdmfKMYXvj3hNNS1Uf
WXoBoSDLb9LVIKCLc6h+7mp8wAluTVP/NVifHKwu98TcuW9gWpOyNmgokHT71OkHnCg0F6N7WCr8
pFnLO61uLZ66UMgcyWWpYp4KYx057M9SVFFByB8lQ/zyWJWus7C6TXBUbtpju5OEYdbXzEhEmxEH
Xhd/K1hqKzltOCQiPgviPHtCPTTH40wRNn4AUeKBmVrb2k7ver5Ll0LlCX6mM+6lxTtArK0N/ErL
CWUbH11ez7PHGg0JwFE1+z0IW6yw8CBaCW54xJ8iV8Q8mCCzJuRjuUOAqUg5WVA4DQOzU0zYXZ3F
8LRw14TWNJdebYYC1zFw41kNlkog8vLHzElH/F0YmvVXR+QvDiFpn1FQBF+4GnOpLfmycXnkzz7w
PB/S0OBaW/gqou0ZbwA5+Jr+NIGOXcLPbaZlR8mPo6UoYrLd0drF1rXQGcTNLtywPJ5G4DEJDSOP
c3D7SQFw067on1Rm+2/DCRmn0in2Pd7TrJwvg9KI77Vzp4dmkfu9YlB9/QLQjhXekzn4kpZ8cxjp
pUNRJaiFEwJEK0zKjpUyBtIgqjazGbn0MWv4GgfLvqGMjwD9VgydjoLmM2oRnVfM2YdDHQB5KFKM
qAwfASagLkdm6MbCFiaQeK2FXqvd5ARbd2e6lQ1OkdCvy+TEqhG8qK5KWQyJjix/B0YrVmpzOG13
rP8SS1pDd0Y7vQvQeHnJ7cHdLf9nHf7Tmy2zQbKmCxf0oWumDzXlWLJl49SW9QOXYpTprOsVvuKH
ZpfOqqo05FJ6zAa/K511MqsOajDIciC07XrEjOTPO9RaTY5O9VjJ/TxIatxB1Y/9TGKrtXju5jHj
4iPZec7CoyIwIzxfsl58+l+fbido0KzLk6WIwoyqFyMulvdU7ptui04awg8+HuKI57wWAn6p2Bja
cBxlTIr9oBIwWKm75R9jKn4lBn3HNuPyHEwcXnScsQRyBonC39JEXWJDqtN0T/H6LFzGcJPNYJGS
T37pNGoLZAUeW0KK0jJpp3kxzBjUTZhUjnyUm6hMuQ9wzAeS10byJMEiEKdYHMmQmQ921tVXPWw3
ZnsVhz+NY4HxuLdWRGSieRA6t/UBUEy2Y66N85YSUjIrhzXgfv5oyejdu/Tet2Xxb04xCi+C9l06
ZPk6+AvP+9NJp8niFHcoZ3JsyU7rPvBVmqjZ7WxkkpUk9ypsSa+ul0ItJzz+450JrWSdv5IasCJG
sJ9XNNV2An5MJ/Ojec1hd7Tjsjuq6SxQNA2z+rX1mohiXD/1AWT6PBjZ/Mrzez3b4xcKcDpDfSAG
LNBeZmlqo8T189kP4gPh2yDI8iGDbkmXVGPOzr6yqZAbn8DceF+HTzlKDqfhxL+MXH2L/8Lg1qUW
ltVgcp9cWmFUlHqOxJutSx5hL+YUc6HK/aF4L/L13P279uVKDTm7x2HhGfo3O8+jQXpJj2k9YdKc
ljDBO+wykSTcQbPZe13gFkyx6cbGMD1Z42/857wLRPPaHmnvf25H+M+JLnAHEqy5nwzS7wYgRSsd
9SQ0+3naGLC58M1ZXxa0aKhRBh8WJB6tewIrJLWVm2JU5VYZeg7HgkVSj2Pody1DfBOomIBAdcI4
5t1iAdWH+VS8rnVkpoCxvINOzoJrCLVPBiXIGlS89eWjTDaw5RXRkv8wzveq6OZegT9nfHaUgZS8
JNum09BFyyJXF8eDR4C3O6amIXfDfsRo8221P8aKYCafpiONB4FY311pLL5oKN8+LR4VVjW1qvg6
Q04DLPkEKdouGkyOuCfCkLURsS2hb7lS8xx2yMJsgtszblo4WeVd0abcVDtGCjmgC4TFm4Ssz8PI
X1hjtLYD5lngBKtKZf3qmBbBGrVdAzK+hcVUxxgsC4nfYozonmgbRzdBLVVsHSwxSBIIn+YhCv3x
vRXLuovNhwEcvm/0HRFGTFrIYE72ncCBM5954AMkMYuImnKK3BOE9va99be5YgMoo29vQzI6k4gt
YfIzjAhlOSzQ3nDH6vfvpmVP88EaeuH8zWT/FjnpWXklgjr+m4TJRa3z9GJw1FApKMzgd2/1Numg
K99qcxGXpelzodrv4t1hFZ8rJOj/JwSL3k9mfJ4mZCX9K4q99bcIL5nDfc3JIpGHDqdgN+DQ+nk3
wbVph0j/LQ3k3DrO1Tjj423fiMoz18yHhGVzLeIgycpGc3SxwoSiNuVbNzzSZhkM4kC3MtVevw12
K4MdS35ljmepOIo3ZoEtXPLrOAgvFJwVGilgDoSB+VarA8lp1wwbg7pRzjhjcnAXIQRzwURYAjXF
DxSrEaMjLNB6LsGFyaYAQnWaDjLwsGGDOhTWC58I8Lgq1qtrU9gxThmfPGnzZiRE3SeLA88duJUg
RpFY4YHVPPiJ+f6D1RZmR9RXexVIthQItAqz0TBqmgu1du65bZ0XLrmZHqqEgSR9opCi7VAw9KAs
DMiLUR3MMgk5HCvJheODVtELRHTZr71DLcOjr3d0oo23YDAXmN9rpsNRpWfZrtI30imHR+9Ee3Oz
oBkSiySppdKhXtNfaznoVV5DTN7wSACZTewxfq51wKy8Rk6Z989/0EpxrDicDkgNjxun6C6E4nZZ
HDIq5PBOzIrF3T+ERQ/xzT3CVkIIy20C724vIXFjhJtKWtirhMuo99ZHd6NwVX6yQFGzUStGaYtg
KJlNvUiSR8/hG4yiUEe4JuR84YI8WtGr5Y1T5fOAL88n3PkLScCx9rc/7TBnJjx/59X740DY9bnT
e8qgBHPaLTpdAg6oEbQmsYC03Y1VVGi+ESGkeuJuRkTK9A/KSroIh1IJyAcytZ4vM6aaYEQlsyqp
i0Q+sv03Kru0G4+32SQlu5H7v7jLH8rE99JXlayiLEDFk1mLyUS8wtqbWUYg9bdmjJWyOdOYrF84
jDMmR9CQYHoIVIKTHjb9Z4MvE6X6i3aC3QpiEMWTAvtxOpnit7Bm5BOMZdc9FQcPK5BTVQv3rdkP
9psZptuacrJzvbG4xA1wGGzV8V4Ni+OoOE6RbHHiO/PO9phROiBeJbg/Oyh6RIWuBoRxVq57d65s
ixVpRxdryhL6y3w0hXQk/U3RP3NQKodhOmCEzmHA2ucHRqAVl/ztmFQOPYDi7KxZrB/RM6r09dIG
TKCfDk6/D07+iWdPEzFDW88oAo9Y7rQLkXOjVTkpUpbbGgiHN/qFOcX2MPgfhjuHM05MrGVB5N6D
rPudezOacgHpzdqUTEGtKv/fpPUrKdf3IZCNu2uqxfifzRlj+CDZ98sNwyaHEhF9eTIZcsnXg0He
vbf4NRr6zULCaDnK8utXcvbBwE/jLwV3M7L536JUJcU88Bl7GiXaSCPQ/4rs9SXiheCFFH99D7JK
GAO8tLnabQ2S4WXwBDtrwWg/pOjph3zHuTSUiryZY/A1FVmex8MBGF3a8Iw9OTYplIH20XqDtLL8
TwMmWXqg2eJqp0Yiism55rwU8IjWBBEiItYnDS5m5g8vklfHAulidVIcoEb0KKjap4gbqasNldaE
scS7SW6LdBBQBOTGDouZh8WFFgTV6/JajpEdyymmrpPADIMNiH4OjYFkiH4SeHjBuli9t1184NLi
98JhzrrmFtXXQe5BFYXSjj+28kaUIimTbrZ++DXyU484htc0BZVrj4DWW7pBqkZjp1fbyPiOTmGf
ZQOUOPm0DfU9M5Bb87CH+kfXUT39KvPYDud4MzD1339Qpye23tGYi0y9AanNeTQi5CZ8JxCP1W58
bu+dvvRzCY1UZXqFHzwBLINpQ/Xxx+uTw9w6qMGAAP/w7z7g9zfkbxvrJZCY0vcZwunmyX+NB3K2
xKSsDZ85WLcy7aqHUlWWjSWdjs3DCk4KZi1HkuB/FhPO8YiHLi41ib5zW583Z63Tjn5WxMV2JdYM
AoHImI6D2ZL5MGpu7JOzFI2NlPYk0qk/B69wqCuoZOWwaMVpUerS59F/RV9f8LTziEWPcRDAD1Ik
5cjn06/QSBdELFVZPHmOqLm1ITM+QrSyFHEbnJDivrMhEEq/7rc3LNhllxQigZkL6YewQr8SOz6x
b2XvY4HyeCkgLrhsTWorsk0sQws94Z9jBMq4FoAO3ABh5m6ZVKJ/XUFEZC+IuLLcoyzcJTZl5Lwt
Qxmaw7BNmZImoeTYh28fc9bywhAAQ5mJO3OQue9Tiswye4nDWXlnARR9HIwMIHFDUU83mzcda0WS
Zq1QGZcOzyc/e73G+6sjuYP1J1pQZ+JTWl3xpLJSz/07KrKiK/DZT8bdXCd4rPDYQZDdZRe3RPH/
aTdG28OwskljH7sI5NUEdYPCT1Xr3fCtvBnlALYMTPnTmyUKhmEx/SqcIWP7AQLQD8A/H8hSOqI9
Fl60xRRo5bUfhxkoCmifXABmKMHHSzMrWvYImzYtybcUrchLgL1FoKhGFpMZ0eNWOm+X2gsNmcSJ
R4y/XSFxAmuwxvAAVemVBtW1jQP9ppkVSbAgw/uv0iPMRMrGCN9tKP7RSSmcEVSZRWqItOZvH6di
iejqWMmY7XX15Ug6C4L2xOUWlaL3+qvnfL3jVBVzL1SOaHzYjys3ME9q/LSgcQM+nzK+01J0Rg3a
/xuItTOJzlf8RhwykSrloEu5x25B/kg4Vf9d839C7tdSfC7vT6KJfhG1UM1SxDR45MsMUPEKzuSS
XKNUitKK3bDifNqUjIvfLb4KYvpe8xB3UhFnfz+yPEeaefWHpCMVcifY7eRgYRIFZc5UAm2BBWGI
VkdXWuyZVmr/n9J2Hd+WWsJq59nRsvdLTyO6XAOXDHZ25zuBKR5/ETIMhIGYJ6b7vO7AMuampHDA
pPx3nyTLwXRR3JaG03jxsr/E6fTNKwOn7S5vRtdp9/jH9ann70DIFCrg9H6GeIdgGQ+KGb8p0T9A
UjeW/7pl9Jw2/s8FwBFbL9mCB/XsTsfv1nUWgvlmIqYNf+oetFEsiAEQqE5szQ4Y9VzMI/5qCjJp
q2E8+A8FXxashXi3NtH7sCaLZhBRMUMwVAZsEuRcR/LqjuBgEMEvRdhIqjfyIcJL8HH916Yi1xeF
qenOXd2ab3pJraid5GHk0bseGqaCqzgGf66EIKjvGbKaedpe02LATczfge8ARVVhCG49HuSICvCS
Pnh74g4GyeqVHDzL0mHzukEKgnIoe9q3z2JuNUKk1W1Tc+wnhJfHBpXo7FZBuFMH4ymJ5ziDQL3s
zp4SLVtdh81knlxjy65VXaofcgWdU26t+1Z+X8YMMjuZ+kkbNx/lYra6BkaoElNZ802E8cULE4RN
t6gdou2nX7M1iYDUSpSWzaIhFMjhvDt+rk9r4AQLK3zqL8txlZ92KTTAWK4nsO/NaU5NInc7KSkS
6J96O5KVUtPLCbYehNcHbsdkGaIwF62fnNu1LGq8WivoJPBRU99vZ+L2j61PyoBFBC9rUIecRoym
JioO1k6lmmSN8jVMickLwNuhs6WcsOcQyEII1x0UQc6xiSkgafnpl5rzII+Ha48Nrcsck6p4Fnbf
K61g4Bhy1XB5tesWxZsmjEPW7PzHfyPULVdN3bR/LXX013klbvclp7QCV1MA9Upip+B7CakYtBr6
juTCY1ZjrcXJ522KX9p0nWWPUccF8PTTLAeBeXVM+teR63r/Y9lmnASTv/EIr6o6T6NUSOACSoeH
Q9hbjNmdtMWqmDVzr5myhlpBK8NYZHqdkY6Du/+pUm8jsx1wshhaLX5Z/yXB4Av5InuvXLBEMpQb
nGfx2x0QRxv0s94EZCXTR+jGm7Raej3WgnNWMHU4CnKVvv7gs65b3wK1+da16YqOkrXC/ukZTUTU
Stgp4OpUfpgEsf8PFH0oopTd8cQEfkakJQ+F7lmKSkUOQOI8Cte84UO34tMJlYwvYiMobA9YomDm
jeWM4PI9kt6Fv+OCOyWbfjzEvdECi10ygTlC8RlCGitAfQoNG1JhRzalCgsBJvIJEvwosKsuVejw
+0/NsEg0TPDpzEZWyiSWPcUEWEM5Ghth0DPApwze/1ifXC84Ym3oXjGUvM+3O6pU0Tr0yMyTcHzG
SSHJsrHp19/Gr5Yn9dZLMoonoY5mUFljdW/gddmA1Vl82+ZY/sDHOYmjECz/Tox7Igd0ir0ofWmW
eVAFQFAIutTaH4ZOUqKq5PEwZRZTjylPBT3rd5IAb/zdRyWguMBqpupAUMfyVhkFjquBLcy1l2wt
JZTP4czDbHeF91ZessVG6YsRaGqB2mjE5qHI8uAI1KQ9x0zbCAlOZkgV5wo3v9xQnlZ7qjRdiI0G
wNGGH2x7IIzHBuPguMoNfmQYEKanu3Wd9IYOF4piL+3rYBLpiyT5jNMdApkBiqLvFU3ASXhEOvGN
XMeTMeqGz+0zAe1PsjAha9oJArz0YTLCKR7OaAyfqqBzr4IdwoQjbOinThuvl3+6jqLVLEYesshg
U+mIm0o/rZ5fQTbYDKeuNaLDlGb54ANjPE4UFM30AYMnCNKS2TxvzCDqw1ZLNSsb3DOAgf2ZBy9B
unYb9aMT8JhxLd37qFFGYWnN0uWnwZ2NbrKbbR1dVrV54mX8kb9ZU/8SvLTv0rTKwZovQCdNNjXv
OpTL/SACwKcxTjHuZaY1cshL+jD77G6eGnXXjrcoj3QimzM0j69sLPVE3cD3Ow8ZV6ezhvELzn+3
Dz9CD7x+57nRHE4EiHEIhyuGs8BYo8NP6omuqrONG342DaMPNMjoLgiIye38NRktzuuAFtlv9Ytp
Q2UFcH7vizxdSQAZVMJutjjbrG2XAQvN4usyIBFC+fXm3qSRME6gFNtgcprZWuIPxvO2nLbjlChI
QSZRrtW0IAkJKc+raED/NOFA+/Gr6GZL3c13xBJXwRYpdmro4Th6o/ocX/XKGT4Rr5YqTJ+eEqeB
mMbhaghb8VHsJetSmc5zzWx8JLInSA23G35WMz6eQTKrwYNidKT3ahSuBm2Jssc0z3YJGk5xBYiw
EJmE8SxBMTrpsZadIzxdVtGmqbg++W84uKaAo7/t5DwflZ+qRv9eXGNCdu1rgHZA6ys1ZMJL7c7o
fdSavH2XQDlMCL+ddThtuz/61fZH/77dbKeV+e2it23dNYe7gelJf6+a1ENo3BAVFnWcxOrKWBq+
d+lZ1JoG1IIGSZTpUFo8LelRXjCGHFRQ70ddfDNbcruIAN6gTqWp92aKZQUvA/DNLCv80oOj3KQB
n1pihaw30jhee+HwYSjRxoDtaG09WfCqwbfEIuKmIJ8OphoPWB864XM4S8l/puAXtEgFrGl4K5tJ
Sf7atr7vSLI+v9NTLr+fcN27YjCF7gK0Uq4KQQlboSFVCJBa6nUm4PtKndMOHcZzuNUEhEZhbAWy
+4dlo/r+DSFJy8gVLhHPiDH8fmNywc97G0v8gSoLiEpuiAE4C6PAMKEBujRQqcwtz0PZ/af1m86r
pvj/6/xfT6fmfehqPqH4p2HBuW/tLyZx1YDfDvFncHzuuH77qHqqF89U4ji6MWhkXDjFoTBlpDn7
/TWuHZbXDndxBQgm2AjMhOH+JyjYfr1sP600SBkA9D2iJEc5RIPTENX0aIFJtEMnH2FnTcC093i0
3xTGm2Hyq8wvfryLTe92JZuIMKTp1bwe0eh7yzXsrS1buCxN9KUn5RHSDIvZPRhqqtT/wEV1tOsS
jFozEAkfjsA15XBHYzbh+MjpAMoZTSffj9u3kfmUV16cps6kOBnJVqYIbmN6t0kpjTyxkB413lnl
YHKVu7fF+K8Eb5PR4cTCGl5L9dIxfGm3qWRSwkJuFqqzARlXh0KiURB+tQzoQ7Kdb8CQHvslKcg5
J8dLF/SqFA8mJMP9jfzMtV28I4OMnymuY8A6dvXOkbQ142NLuxsypNqpi0jM+eg0/Qixe1w6LdO+
KEvd1m+803z0mfdGqmqOuS9kQDd/AgUaTOTveH7mfMN1njEjQ0ZnYxI4DJc6bomJTwLYatXBrvoB
G7QL8Px99LoKud+tbE07c83vXoSZsLcwUrZq3egIJEnIFk0LKE4dpk+eVOSQ/j3bx7Eo4H4kTm7W
4oaFugZYGYQfjkttYRbleLJq83Nt1AbN3otqWxDcsLHOSUHjXOqx3Ye1TJCLWObyzN0I0auzsUjw
daALODgw7aEYlGMxKpKPrZjsOfOO5pkpK5fzDxmGQJNHUS8KqZlmXTilbEmO1cV16b35lY0coc/w
GHZ8QtT+J9KYbiuKNzSbFCb7JWO2NiJSAz9hZ/uXu2VsBnrFm6AMWBf7ww/NZ80mpm4oifh6dWQv
Pvt4ESh3PC3q7Hm0wRY4T18gCYhZJd/uISj4G+N3UnFvM5ejqJIrovSlzcGbd9uS8lhsm5bAuqNs
KCsZDmTKmGE5oqaHcEDOjsnIFp6Hjz2TVoacMiyVqUemKPZmAr8o0NVW3o2FSOmrBAlddA1XzmwT
Z7SeUyExuSQ90MRKbM3cVKejnWMneUY7Q/2pWzjNBrJPijktvrDEQXTx9gdSArZZ+IBvmyMpFcdt
jfZTpiAHGXoO6hS14vE3ocVkjC9FLpEJqOX2RtOY/bC/ovGJz0TT1sxSzXoIP1hMQJjp9tRwQ7tA
9/dCG+CklZAjSV+Q6a9Gh4uXwzZenTu75+viL5DhRucpnI9saKxn7YF5TtJVpb5Ivc3VGsZGoYlL
e2qJqp3DIVuLI/IGMFQi6ZE9ObubkOxJ2kRGOrlWpSriGSA7eu28P2plUGEPJyEOS4pOm52ijL2T
GAoCFrgA1BYd6ZcU4IdhgHVuKs2aldbhAvc2L8M9M/msjw982ertCAX8AQ8IHz9GU2CmUggsbQcn
xGoYUb6eX5mNiQ8RomMSouLb8pSP+i9xNWptGo7jRDmuptUgBKtI5n9lspG1/Gvh/Tvuwcv9H6Kj
SkqOKmNlXGIltCCOuD4+3qQ18BJPc3+9cy172X3BIUjrTiiuN5PSs3Z8xh7bgRbvtwvKB1tqRslA
tM+S+9+tyaPSF+CxQ2hLYgpKk6GVLmWC/IDsNTDSGX3mGfSKRT4TE+CA5MmObFWnxM1WI0b49Sy8
CrFw1BbmPQn156NpaKKa5P8pKad/IhuuiP8chWTzrcsoxH+ZyCLOlE5ZhFwwcUVvD5pHQ3Ly6NaM
ohTPe1UjMBF4pqsSNAR3+I/vBnGGMvx2SowHZJDqtp5QIzcDoSg6ZMxMY09YpJh7URIRITLAjhHd
MSECb8P+Va1HB9Iy7rwGDpOisMXHtwnAYlElmPG9+lko1qwKXGhuQVTeFLLPMf0N77BBlutDqV2x
tLiZvZTPKB8jFtT0UIciWiXfZ/aV82fxm857t6amfJxBdmf5uNoYBEvEdcZaGMwn3YquzuhaFhb7
W6v6CFroPbr8V7CvnsbA8aEhTT+day0DcrMAq7vnvEpNM2oP1RrCwJbHBnZDvAq/FuT+fRJ6+XkQ
itUmbu+6w6XjsmXXevsnbjmCCqS3bczT9eGj2Yni8JR7dk9jHSe2oVPct0XUTC4XjT1NOx0tBBbx
9ABBH4TVgMdJGCi2Vx3w7Hj3wU87iYUMJLsWYWveij7m2wZ695pd2evZVxMwvKcNDYz0CfKv4eVN
FMZY1+Gh8fitFA7TvmmCgxfgoYkv+5Y6Ryb2Up5pMDk1ChmtXR8VgFVIcnDNwiRkRf6aTn5WAqDY
bRQSPVbCn8xv5sx3+r8a4GKk5HgysA6OBxoAZ8rXNLxH24RTg0QoSku02wS8z1JvQHAwp/ZcWk0D
DpAIlmwDBlYB+HfykzAI/WNg+cN0hvAo/8YnYwtp1KnTS7UqppAhJTbGwwvX5Lw2Ki6pDZEj2T7g
E3R7z6zVaA6CHay6tI6zXefBRs6ZYTOz2MXig9p7AKmTRfug4FSHvw1t4LW+ZXGWrwt09BZYkJYH
sg5NIZEerD3vaGibOvbxKT2k50MhYuyhQMZQcPowU+bsH4NcfUPopb1XE//ICxbbv4Gn9aCRBr8F
sgK8n3lq927FoqRpomwOzypVi8tcme2pWvaV6CO1bmtwVNLaWvi8I/6v/q6WMRn0DnhX+DZeQ/Jk
JkSNYlyDvb2UH2vkQdFeUjV1/Qn0ds2vsn9VeAlyKT6QBVaE9c0eIK3hahK0KEzc0WB+QjxLgJLK
5Tn3eqyHVL9C0qFnNTG7NazBtwCtPssj9Ky+651bHUYhA+j9nwnTIh+nY6UldrJeXISBQbPiw4dZ
C06IkC5jWHMoFl9dmUL/lCBKYcAXuW2zaUGs5bRYES7IsvdaCVvBpbxovAO0Z90F5QvYCI+Bm1fo
hR3uPV2aeZAXm7bcBFGYq3IjLuJzf9EX6Gc2eO6wnHN3R+Ccwsb9bvL6tav/JBmR2kRhZPAGVrbR
MfVJLzCdP7nt/dRt+cvCb2VkEKOlBQWlYFz6HrxQLoeFGNeaHHvxwWULzhOaVy2YHkNfQwcOXn7E
bSs8rweHf9pTX+xOrn+CShQ85NA1QdHM/auqi2SC6ngmUWcpHbxH/Hx6V3LiE7jwaPT4m4/geRy3
OoBtjNcmnJRTySIDaVOeG2vaTbtiZaXeoIbJh273/wBSfqrnvvs6BR+0hj1KE8jrAr0QYot7ETdG
eBEV3vKO8wFOCkYfXklVUMxm+57Ve1oUqTHhf40s6u7CpiXptnGcd/fyLV6uWdrcg+totfOWi3rN
JJxqHom1dx4KDRb7PownJd+Pp6zmYbfc3D4tK2/QyWe5Q5SZTFuSmw3QoxusKJDOWR05X5CsaXlk
1DjaSOx9yVbKhqtaHSjcUgrSMkGVmO6YciVHPC+/Bv3adQOq8zFwKmTSVJoYfJkarkUreY+WjMz/
Lq5hNyLjFkwgFdPNzLJSO2YuyLjntl7SfO/l7G07c5NgAGBue0gEWobpHHMlwRqYaLeUe3ygKzQU
pAwyf7oU7vawQjigNHpobdTXv0JCGnZNtWLnwyaWNb5ISGAmVBJE0cs6LxwUNewyev3UK/meipVa
9JUiv+UcxKqrWnt4N/6NiONNz+dXvMsrTHR9An0QgzeFvGfVZfRta4QCiJYzmCI0zQBmtzScWPyE
+Dbz09N8YiNdrjgOdNJ9Z837OJzKPee/6dyx67spn1rEHj9mOtf31ECkKQhnP0GYD9d2vK+Sc4dv
vzXo+2lKix78kC2/RhQfqxTrGfTAB9a9JFW7trG5izl4KEyM1ItfGPui6E95r7xVgeTNi90Oy41y
JWqV+Ds6JPoLl0VDRaBZFaWPG04flybhGXMlzFKy+cCffmYxGIBe4s0Hf8lB7a+YNirUkY2Df+Hk
dEgdXrwBlvOknTf05n7WnOoeTFTh8bP3MqrgjAb+JPeOcmdfzeNMu+B6POfk2jAj21IjSkB5GRyX
YufySwzZOoBT6GBQZ2FEdN4WG1PeIdhXNWSKDiMs164AARHi0QjwV9xw5w5Vgcz7Drd5pbRJlS8M
HBb0AR607+iJNGXmx5Fzj6iqqQ264DX6b6Kga3KH0l6+E3f2ovSNStAZAbrsYtA3zqY/2mh1l5i4
2TZ4hZGInURABOMj6o7VcJQ4A9RSvfuPi7TRFth5g9EUG+zVhSMGnPT0ChDqk7NmfCspnQ1t8uhq
Iv+rYKnZ1zQsl+4GO0hOdhVlQCGoudVg4cQialgTBs06CsjwGiibx/0hB8zIaNxSekuCfm+XwQ0W
fzDFrnHD8tXyqKESumDc4ze7yq9iWxT+jCs9md90+h06G7lF6g6vX+D/UsofqKjA41JMm9PYR9k/
m9oG8qIY2jgp83qL2I/esdn5mZGns+dBH5u+ZJwhu0x0dukjZbTrvjDSFOw435ZnZJhw5uXZoRnJ
R7uXPj7ODDRR2IdDXPHrjlMCp0r0mfVoGfalspiIAQZE7YSAsLrwx34OajwU6j9OuQSjyVPRuL4K
SSRpQvZ4bt5LXYBwKduiEcWFHsDGbuUwFVGtBsBMMeOxNHX0wkAqBWnFjrpYUHYdR0NqugYUwG2u
ylJsJV3YC3M80JlgVEDjdLq/b1Er6Ydb5kryRJ24J+qt4vnv1HxeEsXfAlt61SshiuCN6Fk0cjdf
wULvolwgWGxMTp3fc0c+HRj/98gR4V2oaWzgSoHhzi6u/1F3fEENuoTpRdH3/QdwUDPgYiihBCTX
bNmqr3mkIO7WMZE7ubrfhlVoCfddB9RPjuMyroaff4KaYDrKK+BiBjCUIB1PZzo7SMYhIVmDU7XI
SDqzl0QTbb95VxGht79x49/pwsAx6hm+ttgxQGdNamh/LiSCe3m3BUnBxNZWoIPttR2r2KO9sPnQ
HFPL4f1eIsDrjSoDP2cXGUtMA6HLL02ZWUsLTNJ01V7n1Ox1PDXxNHEqT2PfnWQm0Ek2WgqPJILA
MSEZ3OIhdgFLC7jpXX39ages2t3W5JHDg1KZ3MMtZ2dxeZCRDpV77qxdQzoMabvxeW8YVJYmVodK
QRxV1O6+xz2XsKdkzsM5HCxUhMLKBZQ+bXspbN5dYl0dNmATirCvTEAVUuMb+cHibi4lk/Ye2LM6
c39iVq89/E1jQW5j0iDVQOWW0YBBzVKKVcBS/wOFCm8nR+qYzZd6PZ5zvAeciNngOoW/nHqRsbku
33kHmGt9GTjfj51eDu2JgS8nXawKfGKZstU7FnoXk+UnYv4e7JAN8yfB5NHIp9D0CX7XhZNpACM7
F2OVnnTyPf1H+EtDEdLe/VP4Wp2FNgZZFofDfPdrvjHgH0p/T8Gz4+XeDDA9VN5yBJBnuSxtTrm8
hw4bmemBK9J4lRJcs+96Jnv5+/UJHBJyFc8ReJS2dH55D2VqYwguehWWU9Alb1DNxrCHdDEpmhvJ
DJjWyCbdYChzqFA4rlmNIopAIvJhrA89WXLdGN7q6fGoo0bAcWRaylKsshjjILzjZkFUN5F9QZOQ
AIBiGBR3+cAUOIz+7DOu7TaxJ73oRx0aQXSfBezM8V5EyeXVvTD1RcW1WMZ47MZ4244zE7R7c9XP
rWZpHOSS0XEy9g1XB6Ya0Y6vHa9QDY8MNkvMZE66NJT5+dee5E7ayIl2roVfjxXJhgneNkifdZfa
6pyOlznbXg1yIjHEkgl2bU7v8I3Dzkc3EC2yOz2yF8QKrbqEQS7H/tmTeK7q80twA67fqm9fOSbh
MqgPpH6E2CfeyFL10dcHgHQ0jyBxB2qYJcwzk3pcfu2XerAJUyIBf3p0qzzjrK+g9vLH0qMOxJJR
/ZcIDE5j2ezLDOvIIesRDGDqSAN0ZiJ+aEO1n3F95/5vEaVUpVa7q69G4l5XpFMu+pE8E3xCftdm
DPFTIeE3mSr7LtsyEpuwB+pFtK7+RZuJH+wZv/iBYM2Xputawta80hfHN/rteA8Mxrgv3+ZacPBx
z2LMLdDY3/5CmuxvOavios8X7m06JmX+VF6iQoSM5UN1vKut4RrYQR9D3b622aXAvRrFBZERy/4M
Xu+fUrkudgqtsGB/qOheoBdHVWfEevMO9+RbZRACpjjudLurWOzUgsJMUyZZfmw4Orz69uLfgM3o
B06ywLpErXHYmmleT37xV+8QIr4PPdpYlV7mtMsGgzSpYe1gfSXivdo3lqIuu5Q+u6wn24Af0Cl8
q1BEyy9TECI22Ec0qx+ba/1v2+NJOaoT2OeSoB3ko4wdzQ0nHzIBJPZpV4Ryo1GQikDsv1fqFfY6
URWeFjHPWrCg5lZ/3JP/v8NNpjxl69EJJ1xaKL6/nnVEAWca+Qip+mwjMZ5aUbqle/NaURvNVZim
9+V2eY0iBReTca4AS8RdfMaq1txqUg7xO70BlZxbyx0LQCFxj0tWRMKm5QCMXU477epcqRdx7Cmu
2pmG6NanG0dczzQABwDi10R75maFHF4pGG9tVdOYwfKGN3utQ6Q4hkp/cRqiCpp8qc8ZLlqkL2pd
e29OiFlq4FP3ghhtGgHtdwKEmtksUa9314cM4/mV+EbLOKZTZoCZxjhU8d2FnDD31X/07aizASuE
iFOaWHur8HPKIaIdQDio8P88OjzfYTnfxjOePgq/o2CsvV9Av89UTXw3elL1HcgIjXjeGHmoCfoF
pOiCfZBz4w/WF4PlpNc8004ngBFDIJfaO1lt4lKuupV69gy137Pqr3bqA/lVdrYTA1vecv1sW7lv
nLhV/7Vs6RGeLs956RF6r7jUIe/2NigsljfT+EF5H4YQ2/6nVwgUTo5JXSbnrG9W2v4nz6Hvfic0
I0m2LNjzwHBxaFcinSoccqa8AP3I5XLark4gluTOiZQPS+AUtkHOPl0UxN0FodfP4tFwaSmEAviO
mfPnTHQvm8XZtcenulbyTn5BCG9wMegt9QCUkbAZ6GFX1Va8zXqQl14JzwkU+xwnOWDjePtouvI1
wo21VlC7Lwh7iYk7DLNElBoCjLOyILZ1H138/VHAH/Ft79vy2r/79Gwgf/MS1i2NiwLDq1bwnH9S
G7/Nv6Z88MATVMok2hYaSIJ/uWF2ygzAXZ0gdtnRIxwsBNMwHdEhn/7OYUPgfdUc/hsXISjDWMb5
16C1LmHj0UdPz4CjgG9q3ReYDTUmwZEkLw29uOzIRLKJeeeJYU97K3UAdipwa4Vui8rCrx6j1FSY
zVfFEjZ4dfRcxd4hxp7nTIPb6uaKhoWo/ne3lBueqLNZZDHWGu1S0z3lpHmhLWYYbSvLh1ShvafJ
N89c64AtCsdgYPRhWkuMgcZdS047gzPzo8R1E7wmFe95AOyMTFDSK65k7qMy+p12vXxV05BHH6k0
2qjpQ/SlVWNeiKZlKQ8a3dZ7i9n51Xh/FnPn4I5uHCD9Gi2r12tUnHt7vYQ1oZtoGytQZoRpnqpG
HnV0j1YAzy1ixGVkSW276dZzgF+hg7E9RxCcGxY4RI/fMR/TiAzH2xEJsqcSLiV4mVuQtIRqGX/b
9NXnqzPlG7/1rL2Sgs1gaUx0FhpwuotM3RWT2KMOD774efyhKi0fT1HEQyxWhuCi9U+7EwaY7GcF
4P63r486uytbNxcCeoD8AUvGZFcN4ls07cx3sw+Lk2t98J37ZMKaKb24Fl8xuSkT2nTLms/8koIs
HFaEUV2uc46duaoDCckPgONGlnOu3Z399BU9r3Y+0oZLmbjXU6ij7LYQ/irw38gpz0bGGQ0/gHKf
fmAW0TUeKhlYSJ7GlYWFd6PhJ7mxua+XYbFGTotA+y+Twht6Y5gL+/Fr9zyRZuNtlRRND2cf/Etc
gpP/S6ieWzvqel7sTvqAeTXe6WZr5P8Pp5A3p3VExC6hFNknMaUsUk0sg1iTm2cZYKjh4voUbL0s
vDSc//taqoX3ovsVdV8eW8kG1t5CBgLLa5Tshc7F8nsGM5I6U+aznrwPADuzUCDyLJeFVCKeTS/U
BL9gjL3LTwQtDoCOOURjcQZWRGTKhmFcy/64tEduDLS2hmb3Qr3anG75SkjLJawPGzS2l4Cx46PT
EIGetnzvYI2zEBodefOYymxHho82K2eL6xhCvCkH3av+Qj7NSS9zt2DTtswx+yckicptUO1SC/zq
ie4iIox4PeuwBnZSwDoaxt3bj2EdA9BJQ4lgkeK5zNWLyOjE/Q9GnPwnivnLaIGaJJDlXEbflLXY
LXyjkGqvItaCsE5uOFXtQub6eGj6daEivr0a/V+aZpE2Ptv33BM80zPSTHWIq24bkTOhOQbTZPdk
GXrhKg0HOevNPy6HMHL8TE9SdGUc5FsWh0naqBgPr712z/C472XSgRB4q0SFb2mI25A3zKIzlQqr
GzfnZo1Z88uEF5PdO0Ike2FIpoAjrIciRDNF0Ch/ex42X6vp5fvS3+4YGsc7iQqzFdov31GgRPZL
PD9Qjk4fqZzsp687/3eIM1LD7DokF0ZNjCp/OBrlC2dBHeh4SJTXPTvomAKk5isKrQQQ2fMNhYUp
9FMWi3lD3mDZykDl7YgtbXT9Dlx0cRFQJSgJweK1kxfOTq8dRKYT8j0i6K5Q10HQ11Y0k8Hcrsw+
j74eNQrt4Gu2u/CadEqmFhhJI+2jDmZvyLSE58/H5IUTlmiKbPAGYO0TvvxRkq2Mora48SDCZIDp
zIar8C7KrR16NaqtesIgh7IndyzXJJxPxSe30Y4ielsC2OCKVj4d7RG4IqcY041IaT3z+1C1o2ME
3tqVQ3tBjVQMnoBFnnczWlVqgupewv2mlvS6W6i6gYIYfiCs8AjqLN7r+Eqi4oVthJ3GNea72Tvv
z9L1VKEFivdoBcSa5BZps7qJaxf4QjmqwSwY10C/j6Um0yTQzeEKhwn59QUXOPQJHyJT3EAQTBbl
9q6kR/S9J82F4x8qWcPHa6FlTRXJuTFsR8/eOKYJWjt33p+ccqJsGZTCn9DYh3Dl8wsFEQ2JXwsD
2nboU1ZuyIJ66WMVTKLaS7pdC3A2z9GWPvQR8J8YSBm95fz2dNEcx1N/+VcDeaCXD9KPYdLmitHO
5Dmi6mQOE4VBnBWqPZTVRk3F/QS6KlJr5X0I6HhDQdPGnMjqg2KlEU2XzqZx2yL3IA494H+H/9ZR
9dm66zNMVHG5w9eR/7igWN2aO/5J/FhQdiO08zwkYhq7NLwQzc0Pn1GgkiOGV+FMofzty/wGME94
AAmofu/5D/Y3RDUElTYRL2Ts7IgIS7PnlsiBhWNsDDNoLs/VCesu9cuQC+PsokiXknCD/nYf//tE
Cqt7DKnwO8QNxFJwFC1py3dv8IGatfGaaU4y0pGrWOpmbWvca8UJQMCnhmrKX0gZWM2Ds0GnfOv8
Fp6XQ6iPjrG/6qZ2N6ZmMRD19fjioxgjzD9EqX4zoTrc4r7d/wEXzylGD+9IhKEoq05lZ2eAKHnu
E8gOs7nOngrTW+2VB9myQbqvl5lD02m0poAdYLk9OFTaBvLRbo65lFhiQIDZT5h5e0zw/j7wfJ0W
CC71r/Rj4acU/PXHq8ZI9NuCPcjoBtCRdrX3ui2aacUJ6Uo5NKyiAi9IzDu0CdCm6VMPwZz8+tbj
SX4PdMXnQ3JQWn2xag8YCnM5QTsnYjILrgCPK4L7getg7t92y59j1nN/4y1CmV9trHS+LSh/N/tj
VYVY6469WcS4wTv2/po9bNmAD2aTWyCoL3AkY0E45yB/ftkqhMTIC+h0MtdJvMgqRoaBsE+9mYbP
HjgrXJ+YgTrAbndllWVJ7dJpjJbctQR5ljqxhI7WI4hPBICW4lgbom55agTASzGrS2pg4CEXqF7F
wXe7uEY88UWb1wMQpL8tmaBQKeZ/TldEUFFL1rP6aoJ4I1/IsFZZ3ULH21dxG0njbhYBn7vVO1Mf
plqTWOMRh0ZrDzWOEdnUMIxXW4hHtyYn2lV43NCl+EF7B468mDDnGKf3fw1EV6Ng9z23PF3xSJ8J
xQe+iQztsPMTyppnvAQXjgCWYWQBYB/88wex+wQA6vbI1wOzjjKDVuJwP4pGRAxXSrkXJPp+Ly7K
M6flGLdlko6/8nsUXfP0FiL/g0KuGAcPsdM93jVR5+kbgwHDidwWHuZXD9l0SoPpxr2zf23gh/Fg
Vk4uinTD2O3R+oBVO3cbmzXFZBirHWscSTz2Izgw8Zmd6WCD6H5LCmAsyqgFn6lzVjaYH5QYOewm
UXMBAqCs7U2YEZ+yBhkZWVkb+nf5ggLhH8NpW6wuvp4Jb+yQQC2ptxfUHePc67aTx24V9iHl4k/t
30D8Dyu0ovd2N5q6WnRfivF9Tp2XMVsnnte2Nyvjc2ZFn4Td8ksIcSmepE9L6CSEVhZICFiiI2YH
R3bCFmYpgeS9JUX+t8QYP7LmR5uyyNXq07fIh3iN8ps23/qP3dXhGU5qNWY1THKJsb86I03sMLFA
ExcniT9KgpqgGvnJ8T+vPefPtHn/k3c3uqW1E3KPBdq/Ql0UVnstIuDmV2JjQGBPjKDpZM9fcE60
YGA+rwmU60acBiL8iCusJt4v0u0O9RCeLYYvhd/76MrLe6iS3wzgfMcnXxVCo1d5mC7VrTqlIfJl
xVNkXH++7rXn9ov5UoIvxn7BdNsM0pnAsVy6FSdELsfdAYaE0LIN/khy6CnZyiblooXBwmc/ztKw
rh44QXr6SuLCeedwYpJcd6TXdbvVfxBOGroS8cZa0cFOxl6Z56HmtqIA8/zqWJDAoH69mjR9bos6
wXAe2efQAC5Sjm7Boc+vj0RCBShCMYVJV0fHirC7p+QKeICRrJzWspicI99pPr0Eg7slky51hYOS
8hBFPrpHGldEeFk+Jz13lC/F8EJMN8OjYygGATnIRbwPVfwi2sDZJD/a6IBOzBXze5znLqwNpIUW
6b1UO1/ju53uva+kWWvk/xnqV2IvDmIzEmdzNe8Ovqqc0eKn09l0Ej2j3oV7dDMVlp94vwUGesl/
ut+9fUYHd5nReeffbdD8+apQwPZl/Md3+1Y4pYKvswcsXHUeV2d16knX7NS0ZKE+NulO45qK6PVk
llYLrX1m/6WJ40v57CR+aTQgZPwmyEU+BTuXl+H8TZ4LxhjA8IoFvG13YQ9sSBCS3rHt2GAy78FK
wvudEkj1mY89Lhj65xbiCVo3k/CecvjqMRhNXyn5WEgwm63K4+QwX7+oQOgZXkmhRJrl9UiGPeuy
0cfFgfDXygZ4X0K5wobe5DRKgHWjrlL6CRaMgvZxV5t+MvzDKKdKeSrw6T2SnVJyohn+y8PMySYO
GFtuTuzg87P8xdlpmULM/dnez9cbxlFTIDfYweOKpd4Eium6Xt3B64UvT1enNYXbFLAhPh50n0FK
3CUcQA29cet49/La+wIxHMa3T4LKYoOGKmi3zCzzAF7y5nJU7h2dA7G5Qi/yTzZSJZxuEH/kS+s2
fvkoAYJt0Mjzk++VJGGf0qjm8tAr5DrfkPdfrmUyqPESKDRfzLfhSVcuwmb1061OIFPCXxqbTQWw
zYTIMrODDFeLRaHWNhPsgQBAOcK9XdZDmeycz6gYcpi2cWtOEH1RBz17M189R1GyR77fAxvcID25
OB4kL2THYG4t549jEpfa9Y0JcRX1uw9qG2M42DL53XrJlHBzvxshEzni3PBrm5IB2eR6vXuJji5H
uS/L4OywvfIUp0iY5KKdncb0WgJaFGl/CIUPJZDJjwNx3LsiHq9WdOxd5EfLn5oZs6sOD1Oa70V3
NvOJn1Mb0QHp8zzd5hHtOVLLWIL/Y2+prbiCNvW1et0Q3WGLboDcsGHwuu8JQjRUj/dYFENdpH0E
J6WhG346JaXlCKF0ZrLnPyo6WIWmYyyIq+xV76ASrL1xlf5jcd491ZNglCaB4Pp/mWs4edxqRVLg
B1D2yAg2j6mU0kFiq4G7fJ+BT3ShHl1wQms9EHkzv7+5TGpOhzMq+VlIL9u7rmYECzT1J03NOIbE
/fA84o9lW/kj4hYmMuq4LS1tzgzllACkHl9DuZRr53smgnJh0sv6i9Ty756QvelGLPPqnMqndWWd
jZenw05NbYFToCPYmvgms4pqwTBEHTFZQL6hnCWG7ADOMhYeC+Kn7v1IIfZGAO8VX0ZLpN/gPOJn
ydMopJRGhSPpgdHKjf3IOsoe7+EQr6iD3jSBJ04t2hJb+73sYo8f8jojZNX2gP0shNoOB6mE3EhW
clmO+ucxOicE090n9k0yhwwXxYKl9XxaP0S7nlQDFIWOjZbRcIEyVGwJTvL9iOLOc3d77VVibmwt
FyQ+UZps37UtpkYaPvkMoTdFbAVEni7TvOjTeG+P2ZDYF7ldbplNcdBgffzwnfCpVgYxcrigVYlF
xqfux/HnxDEkuoFZGxJXp7yD/QFzajvAS6z7iA4qcG1QRYwskuK9lCrH8/dRt3Z4QuABBFhg4CCK
+S/xyh04ANKvhd9wiLOPWSQ+noFKY0HZdBn4gBlrH/SBlENQoqFWGnhWEVVmWes3LzW+YhiGF5Ii
qA/2D7wGpjRLLqNT7vEX+Neq4JRrroiCca3BWi98Sk/j7oVD/fBfYKPu7dukmATFR98DgB+4fKP4
8Z5UpEc4kBHoGZHVS/xvv2OjooeT3FAQ2wSRlp1TlRWZ95hfe6IMeA6UNPy5mBGXV7g2VXLbUzx/
yFgbowQitpZKrD4LSyTEw66LUQDEOqB9Iui3a/65eXFFyxmjC4YwNMKHvBYW4eGAknn1mollos1e
waALypz03SYU8duWCA5Ebuv70b9LGD6AJ4V0EAoA5DZQN9sbpA9HKkDtYDRcl9reYwpRE7I/R89X
2/337x2KUGNgkwgeSwEG6izXUVgb22faaK3Ar0OC81STGXylhOy1oxDMU0MxM41pj8d7KWLlH5pD
MnOJzJp8/2evt8LZueydvC1ttbjOB/cENb/5PbxqaxO4vcuW9UBU87QRyK6TC5NiWRT1ak/Kp3v4
iLpVfNgSup6lKyml/lpPXsAyCEZChAm9updFGu4VDq3F+0oisl2O2CI7Bl6ejxEdh2T3lzGbjcJM
I+T4oD99w6BhIoz6ZHYaNKqvT+7PKa2tTctrv2nhO1dkjy6POoz/HZWAj7WDo0ku986IXZnGTSfS
HcER0W/fpus3AQBN3fbigMAcPTlwIaRMTcSu1OYvQBTCYMmQKzVwarlpbRWd/PyEedp/xMpkPwdP
f7Wp91MapA1oBloD3SYemNTKeMnYAHYI+1hCRLh7kGWpmSC0tTeYev47ZXWM5MjiVBA0WLnCmRVr
vPK1mzBLvU+32q5len/EOqnBxKsOe18V7AJ62UCeGvNpfGmnmulOFb4n3te1QA+UG4sHWoIeHVUs
HyjT3XDVKrIi5OAXSy66RquxFr0nHjV3Ma62ZdJdmyVtDBmm23w0C/xjh79s+djQEwxIqd7ggyri
cO2d26UOYkmyu+4kRK2ggXL2Ld57jM34QJMQ6nkHA/+uNacPJacZeE9BYBP0E+/yfQG24Vacb9gh
n+mxeWKgT7J5AcPGwZh5AY+HWKVpkU/QAUucLgbhePJrXlpEnsd5EJknOb4exFCPCHB09S+kZPG0
SkmXlBfvCuWIxCsi3HLNZz5P1m8hfK81egO4M1xKNEyBCz9IyeNI1bf+EGFgLxTmZ/lj+/qixZiD
HOWE5AYVKsWp3qVEYEIKR8fjLLN/ZZL4J5cCQ2icynYfgBqWhiMvI29ESN0vLMP2fnMsrmY0AdKS
zS2huRCQZ9YYoLPCs4J/jTgwXyhbIxPHx3E+MP6efb6pVOogmiSMrJgX/xLiz4Nb00VIepj3ZmH9
nSwU6DDBfgc5Zpk8wrlTpnXhvyFS+pAHe0v9Q6vlqVGHXQlaKFRYLHQJqq+bTMsA0Y+OSrlgmlOh
OlOmBMWEyVlWTwIEy+o4DfNQDsH4JXotgUajgBFYg34SYHKQ0xM8b9QzTaanePgv6E3Jz++q7ijj
Tru2QXRmd4BrS0tDC+T0mNPZIx4jqAbs7OAEPRe/DpH79G9CEBEA7khM7LblrEMTluvmw2rjBAl+
8CEcdBY8S1975BhFvIYTdIFiwKYwTpKhfNABwU8lipe6ikKcK+121IEzWB6bJWn6mtrLBfYsKXmL
ASAcRorLWFjxfzngtWZCGrvgoXPMakE2OUsV2ra7fdyeouf4OIweEPtoZEiJIX4HYDhiARNWKrb6
lSY2D+WuRSa/mk+acUVRKF45y9ULffwQKAph6jYgYsboBx7+oMwB9VzPKJHV4eo5XXPtko5VEP1M
6JB/1kgGeVpFeG7WQEBXG/SPT51WDnRkfRixczpQJ+n7jzQly7UKOla4C2nMOFEi+jsZ1A82Glj8
Y4qZZmasRazSPyJ/VIeO7mooHo/u3gokkeFCBcD9Rvilvya1f8V7tH3cGuKijjwQ/ov233KwwOzu
4VPoHZvx81dsAlOpPcqYD+XPcK2xKmVRnyh+penqkosuwqK5E4Vd6YB6n+rYwPUuZzS3424ao60y
ag/9lAm5MgQwmYSLQH7rUixPtHofWJBrVEdxCMWPocTJB2vI0LBHj3J6rzV5Ttuen8tFoTj0Nabu
qVUwz3B6UDJzuJKXKeguG6lqM/iByg8POc4RfPiB7enQjZ4LJADf7GdVEGSLkxI5EY3qg9upWS+D
KWmaWDL+6Uk0RJWRuOT9Briz3bWncufD4VxPEnukSSCi5KIJX25TN339rxpDin2Od/46gc3b0QXZ
faKypdVEO1rjq20b0cMgrgb4joEPJL2APOz8pmvIlT0tjRuE+X3DJmLY/X5QANzSCo6/64sqkvrw
If/jgOp1z04bVAxOHf4m3V7VZ8NsSw0YL4u/udC3UoFtxnHPVGWTA5MnEiHmsGeTMwzf1oZq68bN
zwJ3H0r37HmLWLlMWDaJdc4Mcn1KHpctk9vjgtbOgCBTUpOqzXZ3IIFxw5N9RXhy4X7c0RM+C5UN
BtvKONa0kYqi3nXwAtgTu0XwUlx6IWApfwNZ2tvqHxTl7bDpeEwk6sg9Gtay8FX4Qpp9WizK+y82
KTdbK84RsM3YPeX8iJFXIdzfEsAKjPBSRfvqYORxgisf0ZbTzRLr1n8qYwnRgtGUK5jA+uj0K6dK
t388MKCjB4/x1c6KgN/NUDllnNFChslG25zFHEurNaVvv1GBp4HbF56GLWjEfViHhuEsNKp3NKek
30BGKf7bThSnq3tf2jdJPMTGtNz2+nxd6VnTGE5sOc4AclG1w4Uw4UcCfMEHq9v2rmegv+WTO/wh
JJ2QQai+fuE1LfkTUsBDUOebC+oOfhva9QtqZfoTJ1fypLcQv5SpswkmZhIFrw+9OPAd3OiT969w
wciNvTyiHEKEhuGmuWITpyi4eOYa50EwPfzI4Hif9ZX+fTC+wgFqFZ8ipL0A7PHu7TErb3/GhI2a
hY8X/po9RwFsk/uyCcqX31wROG/eTBs+8udKWWduY61EfbOhFR5ijM0emszaq27HeOGDMxjg6a5U
kVXkqp+UrBRet1mTkTyvX29muewxI5rbqVdAiVwUjpIuP3m2F+iTzUuQUwHDr0UUJAnPYH+l1ela
knRgCWnHl3PwUnC8WE+LQwpXmNnWPxXeN1kNH5uFh2WQS6pkMlv4y81eHTmozl+NfvruvTCnBN1Y
9gdVRrFrGAtoEEor71Afz49rmUV60fuW+dajaVqxS7qYFlEYJ0OOVhWvUcjsiJuoN2SkwhIxWj8a
wCzCm92D3M9DnJPwAjNZ06apdGVVacneBfYUYSGZHbJpfb77O/fGx+DMG5bdrtSRxBG8b12Dpuax
qadzQc3UC3Zx4s+ZvI3RuFzqsFjef6dOuPwsXeUxqty7T5STurZEUE7ALshs0QpZPEjoyJzcuQUA
gU2t+wi4EG/EfDJdpxqmuH0jiiDy88i04Sd0nUvvx8pKuA70DXBh1hMD2Z9NksTbuW6KnlxFjxug
f/2VR96jSauPXKvAc39DSyQhqqv88aD82i07mWfApw9DMHWQYuEmwL3un6FhXzYatTOMei8TtnPg
84h85ygLoA3akRIaDGXhdHDSkjPUi1o4rrndn7LBfzEz15aVH5AbE6uy8ga4qBJIrQ7EkcBEPiC3
hr2yfJIuMFQOcOD4W2aPuR+73+VwNY7Kl4Diy3PnH7ElSsf3jkVdAmIcWLAENLTDbJuHJZAG3Geg
DoGfKhYrTSAEB4XdSjWqTJCJnClmbPB4/rYg10YwAF+CG05/9L4f0qQ8qP9/wW55nfiEp/B8EIkr
fPup9msUPk1IrlUrq5Kes/I0KIgW0mXICYqy1e9Y7OyK4a3g6FECBvyKK5I1XMzkoI6JmICxSkFy
opENHV7DH9iTaDiesFPcwmHmNaLG1lNiwR+EXu/0LWXrFvON5pI9+MaamIGh0galUZmFja8I6Ka1
LEG47su/+IjfMHVsnFzahy/VxL1HbS99oQPz2PVOD8I/us/W76FuGy5O2Ed+MXUL2entL6ZWLoGP
qDtgNzyfQnEniEq7x0wiCQV/zGq8US8/fdYpH1MxMYyHY4J6zyLn/kd5Wl8suECqkYvLjXU7FKWU
gZtpkYixPFqqtAh+YWED7Ioapx5gYoY1C/osQSepZAeIXhUH1aRfmDHJpoeOoZt7fI5aSJtXqQ3Y
8W4lHABehk6+JMaFcPVmy4CcVCaXMhRQN9HKfF8TZq5nssub/DLZrn9SRy2wkEZ+fP9VOQYpHw/M
yMz66sadi57PtqNJGcXq/HuGAwsglPi2qXiUq+6E1CUa+UKjpm9+7l70xbmk0L3Iwx0VYAel3X99
rAjiBKlM78ImOrmxqoREfn7qpQk2rf2y9deLjOEsXFIlfBu1SaOOczguSPNBLKWn3tnNtI+5hQn3
sp6Kl12cwB6f3WnxidunVK2wcHZk+oJNgAAkwFFbZRD2MSn3LTgYcPK/t395eL21Tu2IpLKZTnVf
CuvntqilLHr22LaF3861mGsYPztzwmeWwvIj9preh0HdgvBrKI77UN5nm4853L4jReQuGGpEdbmu
xcy6ATm1/12x7R6ir0ExnEQeO/LAYHK9F5rl2pUn6SaI9N++ONNYYaZM+k5TXW+gLvlocwHqVbjj
oWmFl0lMtf4QsYFnK3AaGvm09cH4FBemDrUFixmo70A3IWg+i16iVXLRdZ0Uy2lH9rvGjSC24IT6
bv/ZzCUXUYebpgA8/TGNw9431WzGW4eUeTqli2uwC8ZgkLPKVz2XobWP4kTX2tDzmOSL5O9BPj6K
w5cmrBfhoJEYkXTf+DLoXk2p/1o4XrkfvvnjEWMyAJAUNsZEF9LRJD8mNOuNZ0QgUlAldrlhMZBq
BV3zgxdmWCbpGOzb/ihh+XOO1vP3jhdk6MNLy52pZml12hoA7xdDh6VcIUK0A2i+HCI9CwjpWlYA
mmTQejt/9ytfHpOe9WJrklI9F4q3an5l+EZslx7KbuhsqaO1ed5nf6QkY6BIoCOCknp5qPMJj6j5
o36BEt18gwRP/9vXoQrauBaLZZFT3QQlX7NgBaCTveHm0vQ91XiKaam0CQ+W8YKNlmYRTlvqXVQC
yG2KY5MdNt7C5HTtv011oDJs5igLd0HaL5GvUsJIcHz0RHAjkE42qG/3ikVaPyXRXK7dAj+80XUb
KB+b+AnCgOK4Jcj+OgBxPcP2YajNYzsp17SsYYxkPcYRH+bK/PqTdA4iX0dHSdjws503ysBg6fg0
6MdhI6gbSnhvFb25MJPExkc3jqQWmucnkTmKvigfHLo2YSOEj1GjGSKG7dm1tWQyhH3dWC2FYbH/
uH8xlI+s84aPfqyusNjxtxL2ee21U+/g7Z7og3pwAy3cIGuFwlShA8jhwIniefkXcwEWcQbpKHjK
qBGMZoxB769v8rh64iG+ZYh2NHTCJpX6iB3jNdg860sqPmy02NguYbTE1s9l6OTRA+V2wPurgT3i
eMdqsLc3vYujWJwFQBwpJcOuhh/UUC4tkqjP+H+hFhmNafOJNTmSJpSth4hgtfytcL2ZsgNvwRZV
0Pnef+pGH8s0mCMtzBSWiqz0uJEpNLX7p4NO49o/8zPOOD5fnQyxcjqMByCaE0iQYdoDHnQzNKZx
5dZf+XRSGaf0qLr+NLVHhzhkJu8DPSvbr0ptxvYpERhSPlTIMF5ILjI6P0pyBVzFmND5C1lzY73A
HfDezc4eYpaljMV4d6ivPosKybyjM14HZCpiVcfFiotg3NNcfIVzPJUicDqyGUIoYa0nTyZxcFCo
iFkqbk9OgmK/wquHHwvJBmreKOtFhAVPb+hFDW6lcwbDF3U9TNfPviijr0VfQyyy0BJ9xRSWTEPa
7vhrONcTZ0X2cX+ErSKSueHFAoJxx+dRawxGZnDqctrFQESGP1G5KSOflap3vT2l6WO72fLU//yD
FO7ZoIBxIWc5kXWoFqYspHL3hViP9+pWA/JACd/id2urX2rcihM1HN9U4XO9SGVVgJfrSh+DbudW
WLTfM6WU1rNz+0REzfZHD0QKBaCZYwskzr5E+2JUa11YO8z6ZfpEIAtSP/gvIwshQeL/Z0y1ZRJ5
PpIbzxgaILDdpntl4XnzIWgUH/PPZ1YFLrcyo7Cg0sAbOr5lYjt5iqqDiGx1X5wpujeOhkmk4B7+
hK+n1xnT+Nh8X4PAGmulZEo7RvWA9l4zFDSHiEFZLVP3UxuGeWy+jfS1Kr9OATl9Fpt19T8GIpOr
rEYjG76+Q9Hpv8hJewLlk8fdSa4G8Gd+ispd/IiOD1kgEZ5B98DzNgQ70KRepLGUWNuPw64G4Ojo
UPfa5d4ItVD9MjevUR4gkBfLZS+MkjbiQBPrGgsCYgeKjbxuBKHbnTTZgcMSrAx1F+Xr0vmZaVk4
MDdTKSD3SjyuLGCXx5N2wY/rVRUPy/JKD0VsahmoN+n3+uXZXymoLyudBDbvzI63phMzs7EeTlIm
Nd+3m+jtidjCjqotybeOKP4jortHu3JZessNjXabK/c8pQBpzE3TSatzQvVjP+fc2cY8X0a1vObU
30dIABxCqu+e4JLEEbxBQUnvh57OCGZLJ9VNlD2OplV7Q83w9IQ4V1aQGfAVa+194muYyLIWbR83
7MeWSN4D0qrA8ShGrrN349ksKi9o0V85r3kfUOWJYh3gRdPKJrjAz4IrB25g51Vc7SfzdWKgKSCn
cZirN3oJL/HRsR1PK69fLRwVaIFFUbBE1k04sB0uNTs4PGNfROt/op9Yg0x3l5FOXrZHo/Xulyea
xQAT6OJrg23AqLU05Vg+F4V76VCSEhEOkzwLdxCN3oDn1IZIna6zTSp1GKGyO5I/GOkt9tAj/J1r
wqFdjrZIuLMVwrd4G6xTS7Rj8zaCqMd3GdbC4xhvVLXkAddNuO8/t5x3BCquR8NiEmyxxhaL8WYm
04On168bGKCM+JTABpQYyHSHLlf4zObIz7TAWqSLKky2H+BXE8RJjSxq0B8c953rf0deUbNr+IVQ
tI3FeITdmIhp6xb3sw63Axj2nZbaQ792j8RhCUXq1K7Xuu17LVZSUA7E6hjl9PjWbDx/Zfv1qV9p
7YNwvB+4u2muXWKzJT7d35vcd448fIggH0FtfopAizXkt1+F3vn1JXXgQ5ARef/q+U5lfu4CoQ+w
LE9PQj5cXuH/mFqPMByXObQG/klOIlQp2mBRjj2udvkYUr9ZooL1FbTBFoUCl48SYYPB+azRGcWK
Pd8UMAqo5n52IJJP8178eAcLmRmfyo8xKmf1fjn9i4KJSgO9GPwwMIacDer57Mdn6TSu/jIHLunE
jOuQBbeXVZ19Z3Qz567Cv5cYvtI6xtCh/GYbdXtbT+e2H1PseOrBgBCXXDgLg/hdBeICHz81d/rw
NRDfMBIQ+Ju95gLuS6TRG40MwqvW1UlCshUVDNzbX+KVd4i8YpBSSuG7rKKwVM1kY+XE/6uNhWTW
fsYhmCrIkMygMjjF1DyFPU4JmkwEeP2+8qrx/hSMeaYQzvqX5pys4JUkBrZ35SbE4CI+37wy+yMc
ZvJTYeU4QapwuxZ1VwgF7ArYgsxs7/i6LqVX/ANak3KUpzieom9Zg9F3Xy3a+oesLCfXA+e9S/0A
vSQVRNvApibQg+w67HBcmYEBxU/bsUUrid0XRt1uofFUoeh32Dr2jCd9OwlMGv7f/c56A8q4u55i
XXeflC5iGKS4ucY5yExe/3PUWVKbLtgZvfI05dpkSfYEy2EZc2qy/6zyawOD99D42jy/hPbdBhp/
Lk703U/vALiCC7r39sDsXP/k/hTFpToNY5ps5xtksTmWxZghBRATiPkxqH2zZwVQf565P7kMFlZF
/JweHIzzLhSt8UFexZE4WumzxPGMJ3AJ7heH0zYY0NXhmOXmKUICgSjrQJ4/WYwj5ykTdoEID4lP
3lkpwRN8MvNuXkmwUqOesGr6x/tsY7ipRtdXNIbONzpct0Gk1pJ3rleEfyfmvdy3mf352JAkHMqJ
hdVE4SjO+lXudTipKedoywFARNLEnQPm2H43ZOXG9KH30MB439CdrNMq6x5RxFyzy1yTa6kHG7Fe
LwGztMW/6uerCQlLUbDd0LTQdLj0zZPy++hzKB8nWpmHz2HcIZOH2E/TrK1KCWwU5TssBYzP9jKA
Z6DJr7B2STPhomclyRl1RvSEOoOdpSMISyEMoDhSPaQ4CjPTYeOkZ5YjCJpRi/otqvKG8AaeGNWm
6EGn2u4GhsbrcpCA5iAqiM4w9+G/NmjgVO/W7Mtq8HTr62yxBkYX5aHGoaFCOLIaCpLBYbZNTNAi
7b1SPc0b4rrmKEr/piraYEja67kOHJ/YqmS1ovx5sZqr4cCZK0WX6xPg5LK1r1moj5vv/050BXIz
j3C1LYuQgJyL4yhsGKPGgx2kYqz9lNCkb0Cl8mQCYyXDrbkFKe838hDqJ+OOEX9TXXA72KedU6rK
wgNSx5MrSSUbWagb9tZpuE0Yk/8bfJmcwPjegKZIaNp9WJAYJomGViexo108MhAZXldzMVCmVKFq
UyybLNwZ/GPGql/GplMyDindCBXm7i0k59vd85JirdnapAEU0pANszVtsQOCKwaR6YEyexF0UYZt
d8DNESMf+hfdCnwCuMeHnunCFe8wWBJE0M2tq1TP26RRfUeCAD8GwpxxSXWrEqB1AU/xdSfanozH
ZvqAlkNRuclIdhb3hSDBBzBD/lEIjGJJGR9d855HlXXAl7I4bEs4y6oTieHCc47W/FOxw+OhT07Z
93v3VtcVnzChoE4Km/B1/5GhTCQfCKDx71q+GK1a14M/z0MlLugSKu8IREGdwMjO5QNY2b0yedIu
vzOPvP8qbUxLsUhkJ+zyLTxi4gIKqFSnG0WtAgsuyvjfGv4Kt5EF8DKMs34wmhYDdlfaERv33TDk
1UmJuP8OLezjYu/t9D6rUUkbALoUOGgjNSm1bMEFHwJVag+o8un2bNgpVbWzPcMSXUvLug7UbEgm
eqnYUwA6Wf49UOF2WKvhqr1zqXq3CH/qSqPDTGDST69p7I9fuivYnJwMDK/2LPSnqoOyHIk7osBo
HmPF+j3ZmIEOP9EnnMeQkjL2nX+pjvlaGR9vKLLRjrYiCnUJZOnBzJSCs1UxVgPvqETj9b7ApjW1
kArzVwr68YKKRPNE7seGsV5aLh8nCx66+mgazZXkop42KvrnbYtyGP8/uf3hOu8PqFnGrTKs14w0
VXdMXO+7FItS1/NvQV2DBcavIA8JfoaoNVL45B9QZa+HsX7y7sDT2sF1P8pB1D+IdWPpt9W8W2+T
Vs+RjnkmKq8fkAdgIwj65j1k+W5e+w0U2lplG/BdEJa6gIn83epscsC8ABsmArt7YSQADl3pYr3U
wMAJ1tDcYoecx1aMQg3A14DnmFzA/RbE67XsRchG7poWiM9/cuSHQ/DzhUFSmXJvezlqTQOaTH6d
EV7XZgjkeVvII4lA3Tm1wQmnNgWwDYcC9sMchZulJsWPudwdLW6JOrMKzcT4cjqm2ai8LTtVkwQR
qy5zISPJuUZuUmyOkePlgnUpcDnB8bUoVKoaGcgeD0iH4J72Jg9A7XADqt0He2TpAkav0lWiZdOZ
maB5wucf0PFv7WfjJkwMF6FOJ6TZrkD4WM1K7VDFy7rQV/Z5SdW+NY1fnMC6X9QRIjohPYj3CC0/
Npi6XDCcWabEPho6o1C7L2cAVBM5MGNK2AS2+ufT2NdxbmPNqTUgkp67wCevO/GL/+OpcRbuqRGU
mjOBX2Qp+0MT7/IOIIpNB5a3pXmcLI83HuRv6HLrYNKsoUTAAIypd5nmDV0H/KAlwuIV98iq714x
+Nx6UCnOJ4LzdhGkaSj0UiCbF4Rmb6HTuaISdfglE3F3sAKaFuFty00S5DdWC8srtJBrEnCEvOId
dah0pqap5movaQRMFm84KfY/qfsX4oWhv9P+hvGm5dh8NFMkrRRi9NlGxUoQ4N+L8q5dgTmT69oh
ru1pJJkUxFoNzGgBhNzLKmgGjbo6XdRbh2Kcyu1PxI2rxbBjQcVc/6GOPLwQwiYcT9dqLP19eLEX
2P9l9XvkYzOTI40srEkEpmU9X9T2pyJ/wbnQbRSKtvocOo6JJX6/bPGB/xmoxjWP8sw+f4VXBlC2
hB+tZazchMlSD6GwOU1zsUuefPyaxc7H+R9YmvUwTTVuMWgXNVW2JNyqlKVhDQBq4N9pE+FWo5CT
gaVu5MqYlx/td67TAvHjGTjJHuW3X7PPK7l7Lc1dujGM4xZGBpGs1oWEtXqz1Ux5xC7c/Roy/P8x
/BRRGbwnFzw14NJ/UuxcdZrJ/H+pBPdYJVpB29e/YEimobv5EWh+op2iQMZDXkSXQytyPtcBaIMY
4qRbwaCGoIdENHaUUixgRXmlzIfVDtD2F71dJy+eIJKTp7lfGBSFKPiLiIaa0x+UnpfuYuhlOzoB
7vPh8BoPAYDGURh8XJbJceQPDeyDnwsiI1Hd5muUa017/fvDV4GoLmRWlOXJ9Wr6C+GuI0uWVxWK
m7E38x+r9w+efQtw2zN6TL4Zj1uyIH+Y4JLF22WPCrpMyXPsr/RP1G0C7oOu6uRzW6ZVL9UNzgTG
cWp7si39s2Jw4EPlebnEsaMLyXVeIPcurwuhyBMMdFwL3Z5E5ACSR4e9zH2Csn4l5kI2230ZXF7F
FS+bvHm7CktVCmYkHOZxZ0HxIrx1BK/O/W7rsBXKYI3/7GJBg1bi2V7lN5WQgg2MdhiCgkwQ095j
lzQxOnMHAujBSc1seeYPbAEMHXWnK271GV1OpsDqSMf2zeQPgw9ZwCVBvXIkuHxlsEo9TVKO30BN
XFhByYQuvyGW4LNnYgwK7OupSqrhowcm9YMruWWxDpBa7pWMdHitGa+gcGKeNGVEHzDPp0BFMVtR
t96iuRdugWRs2R5qloDC/OJ/UA0P0fRJ6kf+TeIVjBPDSCE8Mb4CfNV65LRw1RlJINUhfMd507h8
F60DEmrYiysEUTnA9u3PUN578TAF+YG4Y1kAPfkk7mKeQCdREaaqv0SljilJ00Wt7CKI1L3j2yFV
8LxtAxN1zJwQI8c/jfU01qPnfUCzl+RLVfBnjW9eZONskDt2m7kjvy2cRfEpXdYvjEAIDN7OMNjT
ql/GMQ3BqWL5Axt8RPtlkv3nx4rjD06+0YD+FB5L6pdtQH75aDEg1VxSelTObLG1fAJOrHQ53r7n
ss0hyZBcb5e04zuwczjVr4tHbc6k7BNsOTOsEg3JiKuBO7u4HqK53IKpDQSnFWbtRHZjfezQqL9p
t/dNFCUeRC5AcDBR7cZOnZOC9ma9iO30nHs4IKSeFWiySUa2xFaHdWmKCJ1qGK2tjtMEYxeb05yI
GMwP3u8a5/khdG1yCDHDrglcBV3hE8HcZl4KWu1pveWNQDFvpm9xYw4bSeZ6EscaL8n9LafqF0rT
KMoKgRpP5PdDqAfC/GQrpkBruJshQbca3G9DEQuV9ugjvLQRvdZT/R+TFzSCDrvyKsgsdaR9BFex
76/61J2VM4tVc6fymMD7t8iX8RaXr9dgb28MmML8bH/Xr06GT0R4GKjebJjSVhk0fccQn9xKTXTw
xvx4zlAuFhRua+rHBAxd+dg19Z6LTu3E2a/p9+KGYuzqCdf8kjVcymO2K6UXoq3Hfqb6ji6C4jLU
5f1WSG03bGbh/vB8f1IUzIxzM4Wltwan2ohBb+8iyR1mfKgTRH6Iz7HDXV/4F4XmRWgksZr85zJa
///URsg+6v5fppkrwDtzJMy1lkNIXXdIgJ9KTTKgIYvrxYFjJ1r8gtQ0e7zKZ/ybEbH335bnQ0r5
Uep+KBuXiLMhnGfEj6y9wVJc1IU4SHTI6tc/SqFE/7EIsBPsb4SAwlFGa4W23KoDShdKxyc41SEk
uSWRylWxtGK01mFHgrAEZ6qMaG51yFkUbW42HcIZ175L/f9WzuvWQ9gPpGcLTzWM6DAjsuXoZDXI
1XPtj2sg3NWkg4IvFmAzfhIOX5WPDjBeQ6a8axoYpaBkqM5uG+HLvle0q2juknP4DE0YqNqLFf7D
/1WBN7FHUDOKtaBs9N8Bk8CCJXc3iKTJ90NUGv5fyL2FZ/1U63EW9VpQ1U1RpmzCLOSlLH33X5Tw
DqTbs73+ivGLCWarLWuF/536MOnUZ3tbZ+pGckDWdEf6ijpdUeSLRfjlvylJQkFGmKq+nls2l2/+
QERm6GPipgyuV4X649Gb+0zSE2ZFWGuWAHatNFeyufd+cThhsqw+vyc0nFHA+bCIVKihRLtW0Foj
z/7J/ezqK97a1uZO3oOSXwGjO9qBCP7VknCLRRWQvn2XSFukHTNIXnOA0v+DmxliwOS4xKCE+rFp
FijgmxGfwxveERyWWATWk6tvqwJudKCuFIZBoD3VdRuoOCyPmcB67Qmi6Zh2xMVFjJvNIcbVYRxh
Zu1QdJHQNccJSvTJijHbuQ6QLX1Hr5JELbrTAL/af3IulxANcfPWL48Z/c0cH0iR0moZ9Macfx9k
gzChe9tFSWRjWSZmSzbf/1j50xvzc4OR/RBGDuoDcwFURceGluxSHrVr4Oj7NTjoP3IkmuzuD47W
/rNaazPmI3YkGe4POkYEP+LkecGRnw+hNxuPDnLqbGLgLJuLm5hJ4RI0AYTh9gaFX9hfQlAluKyS
sPsOm6FSeLmKLBaJ7Cl/uSuFxvR92lTCnuohdmO8mK2ek0NfA/IDfVHFBIlI6BP3ycpeBQHhQMOS
eEqq7mJaLlAifGIgRkJL23j2OWry7xVH1AAbljaup3d8jKsyQlIEWXBpPAWA7JXF6rw9CxHgzGK7
2scJJ3jM2WNlf/fXH90IcaBU7hoUfHw0jw5i7io1Lmo3PxoKMwf+urDOPER2FXTlz3QX0FcKa0Kk
1EocfJihWytUGwbBoe/FEGshCh+TpZVnFoHL2+k49q04ySmmdlRDAvTvXf5E7ZNwc7NaeeebMXES
fI2m+RjFIGCgfZ0WSQY0GW6rp+FBbM/UlHFpMz549t4XGTS1GrO0C5muzYoubhE8KvTPd0LQllMu
6fi8kpNb+vUtYf8MD4tdQlX72Eu7WHK/NY3YPURTgpqerkObFaGE8Xf7yO7FtkJjhhkYKgX0Bf+e
pgBMgL3C01wdJQnozyR0PDbXtjqA4ANleQRekKFIzGcYPQujgmna9cZZts7+w/gNIxwbdQ/Becls
MSkUxqaWO8quuI3hg1miJ4ivYT4XHESbTOd6jjntTMAwF5Nf8jToSZq3XEJCngDTMprsih2srMTy
ilzQ9VuzcbzXjw6A5GjbVhg/kzfO3KkU0uMdiuAeiQebpKPvNLi3iCiYLEZSmB1M/Vpiikriij3C
bh7lvrAhSbyusvzELcFRRmxVrpVcm9ZGYve1KJWPYdB37T5Qut5jazcYMSiQQdjxF5PQZwtiN26L
TLFUY7snJpPOBBMVy7KhGeLp0Q+Vof/9O6y/ilDri5/kT95BeqRRMV5WfS0qweXpxop2dnt3ARjj
UXufM4iw5nwDTwtIKB5g/2nHAZY6oSWbXR+d9Esi6SFqpgDyrRR5P+iKOeumtWZ7oV+c7tPUQIgD
cKMb8XyaoLn3r6q/I73m4tASAVScVlAzoarFcVbUpJlCR2Ex/ralBYDHUtoPUYbuKRPiH71d/Mwn
P+y5PO5Bx9bSdfHzZ7348A0oDrKrguDrighE5mx/e7MIO2Nnx5JjSafFEZf8uPrcgmO/nSi/heDm
+iK5I+4fXnV4LT8EU6azwzYOQpfwlgG43mEO+r/Kffgmo8YUgZilT1oI3FCMBIs/dDK3+vZLnFIL
veqxl/U1OenLl6dfw5JpxON72vdsvtuWpntiHFKhREdZKXQchYvNwJx6mHwLTVVNgndQSDVbMkVR
zjQiVyjMI+pDZKOJCnQt9JjGDNuUy9V+sc2LE8miWplG31RWHCZ9ln6CxZGaecF7zCKgS7ZAQm8b
C0HK69Q4+ROUiWWF2gBW3dnje/6+P2qANdEDsHMzZRS5vJ/8GcFiDLRhjdHJhqRCgiXGEE/2Bf8E
xojP0SAE1/dyEEKBJtCUUcrNujuYP420ucBQjIuUAXJmBv1D6HOyrQ3qmyh8Sd6U5cWOyUlM5l+G
4nCPBCENemaJjmYljKn1wOqKZpNdEKyEjClJIaYq+o/+pT90Iwj6QHHM+f3GDE5je0ldDE2PSkG5
ll9ZyCckJqi/bMQg40LOmWmcsQFXfYjS7vP5Drf5APXDSYx2anNHEMaHPx+PZaMClrvQ+RDAMfRy
wgi6EHNkhpKhevamdLbFwdM98ALU1H/KrlGlKTEqj/x4ZcKBy8UDDgz9wOhTgN8w5BF2yWHN51p3
nC5xKsqLwek6eY45F3WdYNobOnzJaXWjQnj2qTOjt9ROrDJYjOY/a+Ql2KFHq7nDYrLfte0wvoxU
ZxT4qTXZ3ir3+TBtYd9I/C9p4+Ht9Q6HfYB1cfvHl4PraKsMbPkn4zO5wwG5LSU8GWbzxeZR/xdc
k2VeZgyTYRPR6IiibOfvW7CfIhR/fB+MyU5zbvz5kbw/LHbno8VVYp5Z7cTdCzefECqL+3IFuMWO
VHyOj1RGxuYLVbKOEBq1Zf/EVzD+jXSHg8b/4KUT+sgtRERp2S4YmaAv9tjQdbTj+zX7ibrDJY2H
Isb/jJDJJyWSBYZIeZ/NOJSmT1JjvoG41Jj6P9CH61hn6oQduOxVystsK9qTZpnHC47JfD1BST9U
8je4k4d/C3SRlFoyOWAsHdmx3O3DG+eLpryRGzNyuHK31pzPfsRpx1+DoirBhUkWzUBKIaVxF8qV
4FcsOOEEVZQeLK8uBc2AKwKMB2EVXRPJm/5kTeJLJycNd1Z+w75KiDSLx4dG7O3eZfReg7AV9v30
KT+o2hL7qyYx0eYaLTw98lLZZacNbDszlUe/R8SF0IkDjGQykDSLZQozpoAZJkNecsqyfG6SZ1Ih
lecxX1Bj/tLW4oXYMF2f9uaCopAiKu0AAugTx2eBlGW4N36x0MPao4pSz54hLpamPjrLL3W8Ot6k
3crtZpdazZN2fgvehAojc3ywXlWM5JxzWGpr324Hy86+LIY+/ytIs7KZxuj7uvF5rt616E6exkcA
dBDGNJbVzJciUhQhPq2G4WuyYLkMJO9lRIpGFTVjXx3us3E3KanUv1ZsXEueX8tnAWNZyscabC8Q
Kb8cG/VJ8nn6EHt96yrniaLZLYvVSt3nbzaZJGly5HdfM9qKG2tASv3q4n3NI47uZu+ClTWrOb4U
YwAruTO/or95GZN8plHrD6SGxIWRIqOvCePCxky46HXSVI1M3T+xiaS9DWhf7uDTvcfAxpexPbZJ
ijoRu55nF5372tDy/XaXerXtuEO/Xj3N69nD/iU6lYybU+94pt2y4Pgwe96EQbYL6eT2mZmNefX/
mWcwu67BSjDQwRCVvwC6zrQMXMfEW69lWeAaVftGdgWfrKW1l+zcxBnWvdVeB3lxeKtkvx72V46r
gY7cLPC39YZHN1zMFCdRmfEoZCSzVqB11IvFZKyryJRz0L3fMWbUwfRsSVDaW+jw/ifKCZnwwmzj
UFImmNhNTLnnSVFcAQSCz4ApEty71hpjiA6vyZ/i6jq3ClXAleHbgK5cPJdR03jspkGv3moaFwZx
PADV46ToiCvpOylyPhgxiZ4Dj0ZrRI/bs2JPmweSVu9pdXhodUuWMK/Vs9+2GyXux2uwZALTGcg/
PLQ2Y347XC9xXeKN5vwOlVe0J3lcqErdMA/qo131LzQmzngG2Xk6WkbFCJe0fXA9F9LLaE6RbECr
Zyxrm9/wJLszVtxHjfsHr/NZSKLulgOKwlsr7oNavytiWjmoZjnjvQmI94MDNPRyx5CCQF6u9W3c
+Nh2Djhj3F8NRbgnGGIxiR5vCmWnbJsc/74zeBjDKkJfgSx+VRPUgNPEY+JTGCUn2XOpd+5f7kdn
rpXhkvmbAPWdFfpS72A97nvkHYkIrAYv2QSpBITMDa6RiNVd85Rv+rjH2BTeUEvEDqH2f+2R2tyJ
7YXu1Ter7heHCp2KA/5nrfl+iTPmCdhKaOGqsRBPp697i7qs7OQ5ZinK6fXQJTeKmupDU+5W86pF
gEf5AJBdxzVe/wQMdq1Vui/fXzuOHwxaCNi6n/shgVWiZ8/1MN7UngGRu3uqpTosZG0z9cIQcZne
ZImHkaEuNlWjTajI3vhBg6uwJEl3DGg3Vl+/tZi6m0NgnCtPZos13jVYgfb7UJwCjYKNdnl494Na
ZMObn0xd8NyKu4ISgcp+3FiNXAw99C7sAab0bul9EDMHB+l8cJp1ukAb/yNlafRfBs1ONk3JOQtH
CmoNAjMUacrTZDY+AaOInra+V5b7KVQvXtDk6cnfN1D3PWJ/JpIAEFSuuW5yYXF73DUGAghsBO1j
r0++n8vmUpV5w5s5pehcQ9tQwmHNBL51+bwB5nZ4JV2p60qRMrejS1xsGVcWXI9NwIuT+Z3bfMT7
Wsg7wPgpF5rU3b78lQM7JkGvAaQVLQFhd3rhRQ27M33iTKo0YpH7AXZ5Q6UUXswJ/HffBpEHbb5u
8pTfPUWcFY1Egu8zomQ/m91m4gxWJFW0Hg3kuUxJyANUOlkYaC0b/TKLeDUMDGsRi1aa2mYcqe2z
bsIlJ0xR69ihnYxgMDYyiXIWFRdUnhv0CjR7wtySI18z0ED9TUMsX4JWqT9COXBzCPVo0g7zaj01
Dkdyx52+2XoDJph63sILdvwurnVaHScMCei+EavijN5XaXZ/gUvHG3RmQFgwGVOCcOhzsRx5MCdy
Z1965fJ2aZ+EJpoPMV5+/kXcQGmvxQ8LDzZuPKSCH33h+wn2ZtP4mQMnIvQWE0plgi+Y0sahBuW7
6zJeZ+KGbXPhjAnCy52/i8GpUWXlZ35aYGvPR6DLXNsQDaklOuJgA6BIEDPHCLT0BHpCeyB24zp/
XKz9K68JNKD1Cbfe7OcE8fHG7igGtAKggtDHHo5YDcxe+Mkv7c5+FZ1W+aDGUGo7XDO8aa+Jtis+
YnLcnC+x1glEI8k//5mss0LBVJNacdgNLH5nQ65/Rj/03UVpZd1AajlpO2TrabBjYRrz1//6+Lwd
XzKarwlE7FyUXiaaPqYlAj6+OFDGIXREPHmspoCjacFRLhPYyfKjZtzw/WvL58MLFIkteoVjs4Ak
rlW0TMikYFI/xuE+U0kgChn5T7fep1HkHDBsf1SB+euDpfXqfGNB0CQhyW0Ga6gwwaYdy/fsTlDR
C9nCGL5GxfOr7UCWXVj0Mit1qjwOuMnEC+itzN5QDDHqrp5I0w1s/WW3lnz530/sYEm78jAru4RK
trnuSO2w/Up5Py1OBoFnanAf27+XQbZh/fYGUavotLJfN98tLI96Sv7Pshqt5JkCZHigClE06J+j
lQH0Rwjn2Qk+i26ULjj3bjiulWQ4YiYCCbDOd9pO04zkQDWToXZF+RgzBT8p1Us+OAeqpiMVBH4V
E1myahA9o0y8Pt7W6DPNlK7wHAC8JjAZy2ZmrIyA2i5oQG1cPIpw67wqVOuU6/AQor/NUkHmMj0D
jjEpgdLEqBCG+NoAFYN8TrnDQFSrNyvhyEslpXuJr8Y/MhJLAwo4NGLzwxphWDhBaW4dvBpXMzvd
yQ5u6a70H1rnkj3ClHlfhrlMWe3DlH0VljpbDVZBf2UBVbT7X9YzRDJBN/t33qLCUpmO863fZ8KE
mko2N/+qlNsEwOoMPNDc+wIJc+jO3+M+7r6+9eEStpjkfmd77zc11mkavmaZtl3LeIT07AlCaQtY
eL0INQzPK54+nQ1xPGTXesWCFDleLhWz2wMC/PAs9Ai3TNo6UHS1Th0BGVxETFIRXSZWEJwjkZSE
0NlgO2BQlBjQL72YP4OFgkhY/QQtevMLwT6PRd8B/A9Phe6fxhN5um6azlaMzYRq5LjveWjTR27t
m/XsXfDBztihUaGDfxxwuK5yKKHeiorLjljzEDO3XpLMQGB65lkK18zpXDNDksU7sIOcBVZ6/hWk
oW1z+Fk2MWbVLpW6w3m/XLlYbZep/avt1LZh2EwC1cNioShY74dTU13RBBIPIe9wNVa23ZVr4+CU
anbPyI7btHGrsZic+s00IEegufo/nJz7c6tToxd4I4oU4ja7muPIUOEq8UOvqg9TOXv4M9QfhDR4
6RtsSRYf/Pxuz1WwWSdrRtu63V9IigVWYzuUFWBrDbgjG79oLGGcaDCjnTYAGzOrQ+wlgxU7gZ+q
eiYuKzVZR9LTuFpjsxbQ4h2z2zya2RyVcS9Ir1yvrH807NjcMuA1f9XFaD9bCGq0OHUTMCOsr2Bc
aTYgEv6Op+O4YXxewPCOqZ6RemU/U4CLINbSQzNfe+bcLOaUnyHP7+cyWMV5lT1oMkjnJVsvlMPL
mDYUdjf820FqMbFP8IPhcwbuqzYt1pPQvUm6GY3QwBeXti1PthXQbKEBoAaesRFLS6EW85sRy9qq
L1dzbAtWGV06HzWLHBkjk1dbC02zgm2CCEvs68iFRKJdlxTGwSsOvmBQ5GPFRtLs7pzoEMV7XlE+
OhI35puzhBrr1D1VpRJBQulFX+EivDMWwzPiphZpURZufbQiX2DvgHI3HEqsrKzBv17ObxL1RVQn
Qpo4YQotHd775OJL8MT4wH9b8bGDfSeOTC5bpDtjhVvUNQAnK19YbyNoUS3NJRMRj7MwXyn51GX3
1tmzTHPZPuJGVqZDm8e5D8wxv1kiZuxSs/EjyWWeFT+O0MdeOkumFH2YipbELGc34T2XQA85JEGn
xEOFqIz8TBPMCyu3/TR288lyOu09DllZ8yzbcuSUCxpY9sfuIxFflWgZoKy/YfIK8uzNiB95CXIw
q5WWkDqec6vPCb2VUWJiPhkqhHozi0t7cqN9NSUT7dKZExzxS3C0/ndgrAIq81lH8jN/ENnAYN3p
Me8UPVr04qn910D3HEpCZLNAJK884UecyO0s0PF2pzxAMdj1Ui88/NGVZknJdu30/+ZkBO3eDGqm
naePMfc51vbU2c6fYvNkzlk/8kJTSlfNt9To9CusMC5GxTfkAiizjfbxb5/u+p95i1uHExxfHF7N
P3n6VwliMi9ZBvFuEVZ6pt9MhMnJPkw0IZfeTTotJhkWkNQZdDAGTtgiDaAqYL1GZRsO8MFlnjL/
H8ydxrxywykGaMsIpRhBqzUF02elOBRzYo2Q5hxy32JLplq5M+DStggeO/DMNqqb50Ye1/PA4Qb3
19Pu/H5zm5Zlf/eJe+1071svfRx6QHBSJ/WxYGoIMyPnDL4J5GBmT46qEq+0BTaqBlUcp1Nmb3KA
B0yk99ZZEIAsY7zwFID9kbScYVxNk0WR1iHvxoRGNdjIA5xw1yj0nR6xdZdX/9H7vP/XwwcZwvqu
2tipkejAeKP06JBg1KfohsTJAOMQcq8wyII7DUmZ6Lm8ldZTHpCLUfQfmsjaSerXnp4W8eSAOomG
EX1uiMCGBLNxu8yH/rhdDlhvece/ZieKaOjF2rwPNs9mQu459q31Ce4HHXYcrdYv3Jlr2PW7fhaR
6W85l+z+jVK2yez3l/UttPA8IltortINZ12cpJDY04qwr6bef3opU1bU93dfVGMigGTbATXX61wE
vtrR7roRx3XcQ+rXz16C58rq6NNvoeiiETSx4eX1ciCMm7EjCRmmYn1S13NCU1JTqNdjHIB8WR1E
GL41hPqTr4eVRF5WIKxhVLeZ4D4B/bd4FTwUqOXFqE3R0zeABwRl3xOHzgLmlS0Uz0SRDY6apHBH
RAcafEqR30PZHMdF5k57aWi+Sz8MvQIPuPxZaJkC3XyrgX59+BGvIhYY346vuKAH0HREEtNMAvID
RbbVXseRbe4rLJxqKEEGsR0flg7qpq+rovKGmjBWHuh9cnKSbG59Oj0V0jTRV4HZUmOlk9mWhBN9
Pp9LpgidO63mWaxcPq3F3MVNcFf0FQf9dXzjJAwwY7o7FtMeu7Mks+dOt+pYzkOjVemxBbWs2yMF
hpNQfoZw+UdiTfFnrSVs7a7qqS8qhu/Eqev8+0M76rX7yfR7zq/SNuCa1jGDFoZgXt4Pmqe91Pha
ZwN/7JbztgIJBUfQ0qlIxu0a84KueX5xC7IzgWmstAZz4eySqorplm+FI4OceCuseCWMURfbaL7y
IsfLgCCqFEO/ij10e4UnDsNgpgpazlrCeWwmvLWwi3i0LjfGZ4w0pAV89VYDY5SgH5nkSbBDD2GA
tCBY9waGrrQdE48jEpNYDEguHm/Cp8EW9beRM3B2qu/OlrwzcZKVLKa0VEQoGiUyIOQ7PATVZeoE
sCmzhlpVnk2uKoATa5Kv15a7bRIyzGOxe4s2mZOLVAJeryF59lyhooKENcV30miRiuCgozw39P/X
KA76n/YB2L0dVhCncABGpQ66aZopaITksm1RE9NFF8qTzzQj6zyoYjgVTP8xWvWuhH3rAUidUQg4
YjPQDhXjOKi9JLPVCzDE+l8UR6VOml7n925/ZS3q2LYlnG5tnTFoZ0IrcJsev3NLi6jV/4ZxhWUJ
/+GEux2Pcpfv6AUukXGYxr8rHhiDLnYcQmX5cH1vGcmI1xAD3ieMZsZp+uPIaQiFDaiOgmLPzxQX
KDn/0Y3e+dRdAEUQXh9r9w9JsRgOllZVOKcpfUbt+wQtyJNoxTkG8S66yQLyiCcxnhk7UwYzL7o/
K9lG5qAS3FqgveeyilimrmUyWA80vsRxXJv39RPps9qqnEfvQf8594K4Vs/PDbGhbqBaBHnT9Mbw
MpJrI9+SE5NprIUJxLU4MpPFRox6clIrzB1HNTFwlIFvlW65sk6IBKykqZDr2rW/gRkvpZAvU6qu
XeP9wOnHZVhM/eX5JWXafb/8BiUPSE7wO6x4ljSU7lo32zq++kEldcfmaaDu3kFEJAiqFS8kHvXp
TiyosfcakXAzDxsTcDsFoAeRpgvvEoRH57cnF98Bicw9LewmnXk8gwAJn8BCslHKVKkD5RKNHKrs
Wpf1aMj71JzMAK6J3vdSAaVMH67pcGW1W+Mde2HKXwQwHyq9BJMYYu0/xDpjkUeLecYlza+iWazb
I0qRxsw6qXJu3hyZs8s/piGD1eTXjxXCnvBD9Std9hgTG8p8CVGrrfEtgdUBNhDlun/dWyTX0o6n
07ehDhvZlw0dpZwEufcs8U6+ihSirhbabaysPMCmUNLTyL+wneYWNuEABmfA6RJn6FCWNpa9mnJW
D3XPJelxNTxj27wLbT3dWkFdcskq5dMp145TQ2xdCWke+oooFQQXg+ETHRACiILiJo2Fffa8e5bJ
PmtNggFedSd5o3/1KXyQdS3a71N8oxUHWmQ2aeu7KmnSijNTDvobxfnQXPFMPqxEOqJGktH0okYZ
ySADAf+Ek0V2g4J5reH1zUmmbSD/pAZM/SA7Kw/wnqOlKaCo3Yg2GNCg11iaYQ1TAWP4ep6XMW/E
S9reeQugs3AltuleIO0UhJQYMkBINK+dzsyH29WoHOplhioui4+afV6+FK4NorUVps2Vz6ribrSL
V8vD4eOHcUw+jd1lRf1IcIVnU10JPfwvnQNbf4o/Z2wojN5IjcUXoM04ioI31CdYLo2N5kcI9pnO
y7C0zrLUE+rb9OznBPyj3MmrtAUPFvr78xrWjFiQqRyigJp+mBBPp1CBlOTNsRIHUM3G0e2g19DG
F2CKBAnq29T4Pheu+FPI0tgJXnjn+M834WcK05+sEklbqAlMy3ZiDV7ZUG0uOkoS4L5IEWi63lHk
YPe5ssl6/houtadcwqkqeZQRmuOhaA7M47R7qAP5OPst5iGmUwUXvyJV0mjZkfiE2ft8Rbvuq8TB
0e55Otd9UGFNhQ9MLUeE0jN1HBRyhlqUtwhDfdrFvGSkI94hGVwpZJb9moN27v8K5IZWm1sBp84R
4xqt8GrO+ANI1V/+92gLGJfGSWoOYp0hVfmuovl8bqr6m3qTdkTcdd3xaNg6nnu8cVF3QiwtSmKL
B5IJaG0drNiQ5zh+4p8bvZsHpVOLne1rCbtA6zWvbXnNHoy3U7ZgK9G13jaOZzYdzf1lgYLTRQnL
HlTcN9f6wdruu6pkHbwvAt3LUaxmkvK8LNpXoykYdE4wHzVdplb4OwJ3lcJo0LvMhMHs8ST/HvVm
iOCEhooM0q7tkLEd8gRdxJCI4BgbBaXrD/+c7v6N4+xRXRhJuUcgVElWiGW0vAO7uywNcCeSAe1F
9NnfjEwS10V5mcdSaTw1BsRWpRVewX3tRmkQ1ZiOEogDgtAiJWqh37xKdxcuZmGOvfSyCjYk3Y+S
vDUtX4Rdq27gh4Pl2QJchgLCnqkKfTwhRVVI+CHtbqn/HFk1Qt/4HsGA9I4fMsDO4WTdLSdOaQG2
/+9KJqAyxCFepk65N+jjue1br6HvipjyiRvTjGMU7HAgTbpbRpYlNYR3UiqkDtWutCjb4BVKKkxq
Q4bHTaoQ29BbX8l6PzQ9q3oaDWN2lK1a59RoliQBmm6pDYNH2qfkfbwFmwISbehvPCfN0fzMqB+N
JMqMPrAsupOe9mpu60iicjQO1+Qc7d+4YgqabjS5oAsKBkydnW42ZctqXR7IipQxHjFGY/tHgPsr
AOVz9Bj+BVVJWnp1I/9ajZ4CAn6vmcsGaqJikZbWRaaggrihwn1rCrasOn0DZPoxNadHIcFJgCDl
9i2usq99A9tkk7cOWu5xauYiJbgJoCrifPw2T4qmhQNjXMRi62Qtp8FyJs3adfqdsi1XZFnNhLbD
v6O+Qj1uuuWuXQWH5jAXWs/z6lHWwLyla2HbWWrsTlTx8OKdD+rU0IHzvmeWEJtxQuxpUrZWFU6X
I4WuBf8OUpiRfCGT8NSvJSs77j4xDcf6Qr0LilRK+DIB64qAz16bBjprbs8kKeABJvQLIuPD2hse
GViH8pYXs7pepoX7imECpoYjICoGAsIGbctCUSuuMwL5j3naBh75A8KdFjuoqUjkPXu3Ao2gK9X8
mZzwE2uERufcIH+h+/Tvq4c9XkyPHxiRzDoXsvrxXeT5Fnjf1GjrpMxzycv9SvjIKo8K1tC0cCC9
m7bZNnlR9hnnOv/bODHWHQnc+UCDhVT4o8dMwyS7bqi5QKaZBKvMWdy6V4XX0NwahCa05fBuZUZr
nIndLwOAvBw91k7m9VgIXrbghwawZo1lRBtMzsMgipAR6b6PGq4aHLRfgG+dp9Hz/KvgLT6h7JYM
J6NReJk4Ae1dRXkX1wipSp89kfF04IIBa1kf9DGESWn52TZLeFgrjlVr3tNijADZr1X+zmNtatBY
98lJQCBiIamkmf+ON6uyJ4LpfGwn4ogqgeUWjkcp8j6ApCRXKUpZDWqcrVnXOoZKp3bcIMcz/vhU
8X0ibW5MGtGr+3hj/p/gZzAL4uB4mr9COG/DEFJvpFJKhD8df9q+p7UuYFCD+c05++0Z7mAovNcm
T1VnMK5zeKaHl1zfGZPqO/G9+5eHBTDjwyCowZCvLNEdLJEFWVR+t0xKEsJ5PansC8OaJkVgvqZT
W7GYyaE2QffPjLhqEMJMbS9ZCYr2Yruiy8aHgMHCc6+Vln5VrU4nOo1Gmyf/WJjtvaJRsIODuZup
Z88HvErGM0EODAeqx0vMauofAiPbLipOSNf35Ld65nGHtxpCmR2zTmBXII1qSqM1xQ317wZ77V7I
uJfwLFRsu9Vn8CmUzmF1In5N/nn2jYA7BRG7xnXJe2cwJ0WdUMdBiwe8xthqW+fg2K8VmirJc/Yg
sSoiJJ+zDBQo4DK06IcIOe2zUlvzyORmN3thoMQF7hXRiK22aYX36fWTBI/KTIFRcy4m4c9d3q9N
T861JZ4cUQzQe+vzznAYHQ9boY5v5QGyYdHBxDE7dabgJHgdLxWbd348CtF8uWsNxaW4yqOTVUYH
OwxX4U7xQyj+3JjDIfI7UegoknKmydAcaS4xjaC3J7bPHbt0H2v6eayYrJQwF+cqIb6dXTMoYRHJ
SZ5Ok3ymJOPImq/gDtQd6TYrTBnMl7b8PSE6DdSCpvAFmc3cj57LDzWqVtb3hSM5mowiwFTlAa78
2TpJRCZlLWou7mFm8Qg8bJsHVwB2+vOXWFIf9ZGP7GDVRFY2AAwGtcMI0bCr5XgrVTdHVW1H9auc
7IlC5eyCm+hat5sDiix8VG/653QpTst5qXsM7F8Try8vZ27LzRYHrZLoAhWE9cBgcqWeHlSPG4A7
angCtnKf1Q+kIewJkHCHN41UK5S7lPx2gvggrxCYB0QAPnCH32mUGCqEiHjNRMrw861Uo5XbI5qk
Zm82wHGa/a+oN7GOYCjTY1uHtCVyuLNJ2NJtzCtV+Y04ExQszWT/9WpPRPJ4zTvUxi7oaHiKyoSC
FuxcF41PBR9/KpGs12hz7AFRptwwurnc7xscMFQ+5p9sMJFmkXFenBe9NHq9bRZvh7+t+EIWslb4
Op0PoRfG6oqxtEFvAlRJQe9v+WiN7c9zImafj0671eX5Z8b+iPrvB+QWwwopEFjK0vFfMrQQA1Wg
FdzmL0u295KBhaBGuTVQz4PfY2s07c+H8+/Slns6dgFUPu5l33XQCmGxjGAR3/cHCTikivnLydFw
gl1e15CqX6Vd5PvFuTXsg0LHBYJttn8PHW2ArM0YKb33IEJwj0tepPUakD4b2AXYZ4TZ3kTKf4jI
q1uFSR5PvFmUvAhigC8j37SN7UdidgD1AMEeSIfpgFzy+ZQ9+GYjHRp+NP5RiW9mDTh9aB+AoWG2
9Dic/bQvZFbDg3z5JWKkV2oIQ5s9k4TkvdEorCbOWLcANPqH00eUAXYfLp0/44tkrnzv4EEQuEv+
8TXtMVo6E97zpihWpXcCYl5Jti1BhsJios7t7MTVyZZO2jZkCiEc3iv5FZdRlJ/kK2TCQV2ur0Zn
Bly0aeXeIWua2WaxB88NdhktB/X0EJB6Kve6OO6Ae/1l+oJUMaesSAkpp+/iqdIcqnWdKXyXiLyQ
94Vv889rqG58gx5BYv4Zx4kumpiPKlHBnaA/pLeKZmHiPIYLVeTZ5AILrCdlW9pZs/kJE0btj80V
WnlX5Mp36bfPTB6o8db5VzoRyu2Hic4i0XK6v+WUI6H784yhSFd1sahsyjctqx9E48yKpDRdUYWs
yUI2rhPEovrqpwrVBSKUfMpzZ1R/jSsqWpf6OsaDCRRMShnWR1faaPzflxkeVLbyqo6T0fHqtmdp
XzUpwOyQpfoWDfMelxe2Wpg0pxsoA2vvslsKfeFZH9ztSUURCjEd6kSp19y69kdjnsqrAqvjMG8A
r6TNdvvKqGQGF3mQrVLb6sP8z+oXPxqSYg+W8osRrJd0mQyzqxb+kSA/Evc461Ha6TNFNS64sUjb
0gbA52fmlrc/Fyh4HxvWXMpNUPe2Btx4n6bOyliSMurqj6kUA2fs1cEr2FV8xcpuWIzGLVMtK6QE
MWqdLBuzImp9weeUVmCnisKWMj7T1kEqSBM/ZWogPGbqxb0SzFfvls9zBVULTDu6mdx0BYZI/ySw
nKQY6tthSNpwfvTO3UMYqHlohDnwTx4LhnDOZ/qfFB0DjiOk6cD6uTJZSlhCmUFaH7xg8GYV8Pld
Da4ZF8mfCHTVm9LYtdfgli1hVm4MahsufojfM2jv4enMtPIJsDiWHqSgpRIEv1uDwx7Cq6PfIJkn
K0a5uJ+EveM7evBZzapOX/pVOXO0N4J7EvSp50O03AryTp3vSBFLF3066JmZVa92sqpVD6BeZ7x9
+GZQ0vZ9EmeLI4VTNhm2ioRqLYTXHHh1IsRL/N2CWd7umtsNAKQ3tDGHFmql/JiCkEFLW60pIk4W
F7PZmCq6kLsIZvk/pZL4sbqiMU6iDCExwSSPDWIasVJOG9YOiiek8wy926f7RPOkSGPGjzSCOYnm
MQw2r7NOZ1/x+PsNXNDGtNzc4uXD0DmZKkBMtvyL7EIDLYgGeczQKwH4FJzg/ExcZ1H6ksw1Hwms
Af/LTTnrYfkH7DMimO2iQ1+LxJTbRRkB+OO2t+XGrFwRd81xF3mVc3DePyUWZ5zxgeY80DrCGGHE
GK7RblmeOVELXPU+dZhG3fCcoW8ShKVlqT+wwHn1Zn4swO8v9rtv42/MM8MFOrs2FzbutZa+4PST
BaQj9doPcXAHYqvNBRfxr3M21gnPiwh2f60mcxNLGA82F1JV69VLs96WqbJeKrJSFrQDcAVigIXW
YeCh0kWTT28Cx7BH40XoEFLvEbrtI0iZH6biAGcPy1FY0pE3NZEzcm7ZScCM/0wWaRLotDiVX0BU
68yMk3tmImd+VukMftKQO0Mq6j6PzMlJ3oVuOn3exUWWfS4cCGfTVzzXE1ygfqJ6YJmyod4a9sl8
k+cpxKcPCXwpp9VZM2boF2lUMVxCuciHVLMZnPadEgkMVLrTuTsUVshC0qJVBwibNzixuuFen2Mq
k9SxUwW6AV0U8S06T9uVv5EdduS3ohUYxrxWOgJRVzsJstkavHNqQSTew0rv7Twe8es0xfDalN2d
tWdLAJOKO2gy7wp+bb6PeTAW1poLJncrm0zh3EQdgn0/t6P6NpPGBWN3qgESim3UpXQsh1bGdd/r
Vs2DnvPucZf5fQ2k4UeyaHCnVAcKjr4+fqGQzvfY0D7hgficQPwwGWE3aq8g4UR8kiVawCFpzvLh
ogK7q680xY0PgDSl4TS+n2q6EHLGIJU7e5kPgheMkUVJQGfSGW0ClCRTcPs+DNO3arfBbwHvtLc1
E73dV17owyXRb0ji2dI8qi+3RNiq/gGkbViNKh1H848juGtO21l2dqNQwtJG0nmoS7xnKCoLlCVT
ZJDU5ZL+bzBD0TMRqmKJz2IAM1U6QF7pwNOGnykSuGPMhBPFZ6UwwHnmIGnmdr6T6JRTcKtpelav
rjERXbd7EAkrUtypZt/P4X9Z7vFQHvrqWfUlZQoDHLSjT3nr2kjFSwG30HoKkCeaMKq+iYbrxa+A
3dNT2PrXReRoLLomA0jrYk7gVS3pBRro/cP2KBLgZuaL+KMgXxYSDyQ1bE1hrFtvPtNno3aG9Vtq
dmDAZ9wWLP5FnrqbBIHvziuRyOvHEJouEztBWrdcnUJY/Qx5mwKm53YtqMgnJE1nHAIjtNBHzmyX
Ibc4acH1ex5sFz/0mCFe/RbCpGHIxjz2XnvpDQtXcsd6UqRlQLFPHuNhAbvLyhnA9eIjpw+L6aK9
XyqD3bleycbmZdorwpeIS3mARO7C3KMQ7gNlynaVs4NajX/XY68Pky8F1G8IJuISpbt3Zhb9YWJF
OM8NsP8m9Z2rwFWpnIBXN68woNRJuTa+hexNBCVzBs8BrQG94M2EZaij9uAT/FMV1Se3eJF1pee+
BR4lTIA/ARFeB3EMvhTHRq2oPeewdww2ZFRC9JcN7ciPFONMJBwiRkxYUiKZK+nZFY4TLdR/gc9U
ghh1WOEd/gHYLy8kW5dcE3tUW3l1rR2yp1YcafpRLTCl0eyOX5th9n1V5ejRrUZW4axiv8FBUzH6
U7m/NulXB7cr6Qlt6rl92mC8aLFe/Jjuy7w5TqSOQkhuWPsf6CTe2ZVRVUYnMa+wCBiUyoriZTI1
3UzUbaGzWSPf+NBZcC7YYseVUKQf2yeLUm5waHEJwbJNvBWzcWWTPFXAhpxXanOdUV+ob2zAeYA0
ZYWibaujImfUJGad1gZwb6Khb5DqS9D013h2BYv8CSR1vSquL0KLbKsOGD4zmvySTuWxEQ60H73P
gNb7BFj/JSBm8cjoOMFJacyCZc/mIHsXX5ucLjYxMAD/zpVadJdS+n017b4r4YXA+P+rt/m9ZUxp
nKEuf8T59QEHTbBog2HADOSqD6vnDm2yE8xIEXSrUccaeRvzJRPLtdLpND504KKbDLgrlL3g+nGZ
ZDjgsVdunqI/qqW0MDv/lKdr7EjcGQ979Zi5WwYoxlY+sy/eutS74bDtz5+gh1DV6/a07ej/lbpB
X9KGsv8ttPiaaWPvPar0uGlUUaTuXLuddYXnxDjVS6yc14pk3rEW+rU6AUe4RC5xg5zQKFzdVM7d
kGMeVGC1nPJ6A/16TYVJ1h6gSPPEwPA251xpy2LehnQ6/Xsz0Pi7UVyUQcCOS5hy59qmFOk9wyZ2
7qTM4hZOsOdro0SYsGuV2/U9CwLMYnN+/a3gEdkZKmfwQbnBv0ajTuNKOORxqZT1u6zcbRN2lNp7
SiC+tGFjw+OGX2NtJriGh19bXoPEjKO1WXAB2VWXrTRMqiDc5nfwmV6TBeAYosLh8Ls8GaP82M01
qK2n0nhBEXWszD/Edjgm1r4p40Ltndk4evNQgDHRydPYMBa1vJB1nMM3j/siZItLsoOVTUt64zAq
5M3/AwqBT59nkVufxb9QhrfqnvPUqZ17d40RgWhMpm1c/8LiKFJicnwkIWHyIyW77vfY0A3OhkaS
uSk2n2ryMWA3AvruBqs3pLC9GICo/OFzXUUXGN9PLdsrEwmXuH+K1oCIMTNp7XG3l5zC1xkW4YUO
VTv3w4bP/vpTnrBAPk03vv/OmVQgCHd9hdrmExsNrKE1TuGe4eTNmurXqz9FyYrTKlVvBIz0Frl4
om0uK0Q13Mt1fcySocWP5nCOaC1sjxFRO1WspHst1UaFc3biFrGIGMZ2z5V6rOwxuU0qT0mHY2EV
R6GnsZLB/xIZa97qo8+3bCetb2Sk+lJyK6++LbO0+0KL6pEsJAB4zkacDiXJk6Y58Q0JnfYGb6AK
tyALixJKODWtU//JdMcbquX1lohR6JbIN/GiglOcHMZ2qm4yMjTMYmUSDG3VpTYhZFwxOsR8couM
BJushKxZhWZJJkdMyxBD+auDwSmLm3kcwY4hRgmU7gcYd9zcAIm0btRSxzJzaABa5T89cL9WXL/F
hvWzCXyU0Da4fkvQqvkqzLEgC+pwjYqzB+u8mLV4ZUGFSR0ZXEXDu3WY6q4VNKw3K8LjDB0+2T5U
ispul9Ov/qavOTKNZOb133YcOFH0vfXclSf/BKkiuZT56JUW5d5tD0BJ2MFXyTwGjd00bjEWZReJ
XQaHfwE4y/6mLvxg7ACSfFRWitVljSue3ujGQ/fZT1c3IbB9+JWIju0sHcJH4X0XMe73WxiFSy72
bmNs/Wbf703BRF741M7r4eQeP+kVBFMSdsooCzVuOhSGN24C0f2tbMsEKEkheuBRlxRQiOuarNCh
6YSrQPjk+aW+GO76kJH884aNCFk5OuqqzABgl+W8gugKkJVgfM6jxWEqBuNztoBmW8UsWoxhPg6v
d+9FdXJRG4MGqp/j8Yw3dgygbDQ3vVHUasi+nQqm93Izq5IPNNxFraDuCEzSMH4DUu3hxZIG+8jU
2hQPDWFM+adBpk1nT5PSvv7e+kNFeFdYWGdidczbJdc14aWkXn+pawnnLpY4ZZErJuTM30pF/Or6
C6EOVQaAOa4dP4JYOGCfygUuuVxAzE+XGGDvyMonXF9EYGbJURW6nwE512h+kGhUogqeRMxo2Y2V
hkyDr1yh/MRsFsBwgDL9ZK2lvxzGxkaWA3ebL+8F+LPRufjyZF6Iga2z9gpR8FYrGwy4ORryd+kk
IjfMl+JeiBP/w4lH+hsW7P7W2Wfc2gJIbXjDGTmgIOVKZLcI1v1FONWmB2+BcNRgVfoUkI4Wtp9g
N8uFZlwuCTasvtduGR6Mt2irIQSNI+vSczDrogcW5OuDpxkRR1Zer5YOHkMyRMnxqUzqBgbgltMZ
fXLthksRGSi0136giwESuQpX7CY9vDZWJZXlSuWoBnzs70+phYAjFvOjbVhH29g1Et5StAtpU1t4
BW/6bBheIYT9w5z2WqhskdWO0G18ky/WgK/4gqLFO9sl72rJtaP4vhuP1XvDBeAXGZEqVvuP9HUV
htKtNkakg38tMTIpSXyG+B6Tr++rfDTLGvs5dEik1mFm32FWYfNiydr3oUsjbj40oU+FA/EuSmiD
WSmXF7+epqrZJADWELdfXkwQE/F/5JAQYgDgGV0KsyGGB5AJGWzYO53uzQ+zFeLTVqgGYrTtp2oV
iGWqO5DW0IiXfVZnwHqFMkEi/Pv0WzMuavI04BBI9yUUU1MpCo6YOTSSBGiuR7h0QY10r6ss3Sfg
I8tg5JsgEGlpmjTpXviQeHo1goY+36ub+0t1AYIl9+B8nzurKTNOW0YEp1dlD/7gradpMocsmOFm
O1Wvn3w70vpgbPfiQwJj/ekJyp3qggcNA10HZX4QlUme/qub9u6Vfq7LTbJvH/RThZ8GKAbjv84m
0aqdglcNF4kmf04woZTJiWAhBMlvaKUAxbuBat5OTrSWR570ldk3At5tOaZhCCjByU/dvIrq9Mme
vIuf9UIf4voKFu/Oxd4GSKSUXunFGI1dI4iom8nr/utJN4/kUQ1enmn1fvdOFp6fUofFR+7ChxQ+
020J6IWLFzRw4YcdOiFgfO/R1VRKte+TzVnMY1MpVymN3toQMiOWrMMb4P01XJqx5x/lh6xFOivL
XEdoJ+GNjgp8GrZ7OBCq8xtFC/kWVVogyHt3bebrYMGpIRLZxHzQWdMfNBJJYtGTqoL7R2xfvO73
wYrpGDr3W0sxv4ITVhxTZS3ltXA4Zs4yVebsAey6U6U9hhjLCqH7JORyT6kTb+LdnFzXgXaysUaE
8z4F1l5SRODay3nA2d5sByrF19ltuvuGwM01Ae4VbESX+vkUZxqE64bS75dz5K6vcN0FWQZXAtxM
dyTfjL2a9+uLXVtJu3LCH6RBiHg0O7gAv3kNTvTBM1nHveSeJDL+XXpiCWoNiOO2hcR5VHNOTgDc
CHMvyZaXr9w9JMJ6WgilN+rkMCmGszELWQrhd8ZsJW9z9+v16x7ULVrSAfbJtixB3GP5egdTwp0/
4KsmIpnXGbtXMIh0RYXNGw6dTkN753Ey/+GEBKsxukmbO3uVJs+3wVcMHTw10xBk/2GZaLINVSoY
FQ2dZ3pRz84LINcI1yoTTbhxOTVjxX5JSBPmmsEb0rEtx8tgpYau9OHmzabb9lGIi3qLTTuTdsFb
WUgaysBQGoSkfw8s8gDZEzyecDGmt1E0ZkyxdLakIxM+NKSLeeaoYmCnsynlipbaUffFySplWbHk
BN74KjDBkUpYSFQy8WK0nW8RDYG8WUgtaX9IziE6X320ArxmeJL/dgWCZRZ3yiy48e7SZ60xaLuB
+KRac09lO8aleWKvp7QGYJUlM40qrHsKszdcQQ7lN8jWbIE7hbg0Npih1TSlRh2JMvdSnweP+HDO
0JFEVE39/vs67lkABmjJ1LPeKXAG33T7WF4Dz22xuUFIreH6K4v6C22AWQFHM4NfK8AmYLKA/zP0
bzM/bXy2eeearns4hvk1WlrI+1OM/B/MK8QNatk6tP/Ek7DcvpTD82oZ81tUqeCcik7Q1BMGQrCa
JA9haehtpjtFy73eLp6DpK+UAahzQU/ivCSLg00wYZNGxTdT9jsxw/AwTzyECI1pFJCNFR3j34Vz
qjopEYjCY1vsEoVb4e+0SvteTLNDLz4T3ekgZShxWNYDOanjBSj6FaJhM4/Z0LxZKukZyWTFC00e
0O46r/OvAAUoVnzq8oX/PCW+0uKJrcg2kYzmybVBeaZU1boysSBdS+/OHWMOK86l2AqURo+opLbO
r7NGa09Szs8pa8Srw7eogK14Gu7NRFaUvNIejRuO9l/uzNz3gdVccqFgXbw46mymCBPQ81Bf7uxB
AS6z8inDc/U9Rp5u8ayxwW4DNBHRqoawz7H8D5YeZ5DcxdAJGErLwskqkRLVFG+1/kxVRisGEZQt
WI6rIQa55HccoqlMfk5SAHIFtQNlsAQ5WQeg+c9SmXS6Nz+qpHInoTFj+glL1KkuQkzhO89pOcxx
cf4O9bcSWt3YZkrb8gWkAKLbxCSIdToaLVUz3UurxdP1axUzOyaYT+Ee7if3bwWUINZAUE1iNP5V
9YMzXtjf4gMxY5MXumGoAAYC/MOcs8OJvviJI5UMJcP/wCZA3YLCHbpsdWiADSAdMPGYh9AI7vKV
HCGrGZf7tI/AoxRgyCaCk8olhAvG1Oxqfrx253MFMyIhx8YFWSitee/n2JgdoMGwKhMJRPZAo7xv
fTA8DCWqu6QtUa9yvcoJEpvkFmxJrRm1+M8u2dnfKQxxLINXRulemiFBYK6VwQMz5rd0hClqfHwa
8vISSMyV2G+1lSiH7+aBiG7EF4EC5YKpZelrzYLOLUeazpVIxYlGlMOPZtJ6HsC3toVq4fGIRqz4
OYvvQTiBAYRBz4qoWfbAwrVl8+Ohe42uQ1GOnZ42ZoKouOdDGqvFOHOl6RwRkGRfdPomuiVGmYpT
dm3qf4N+2EqZRA0bLwXwaL5Yt2iuOY1XLOXsknmXE8K17zVAFm18QhLvk6JUEhMLptww41Qwcpk9
yInJXwa6MoUU2Cuf0Zm51+Z/32DQxf5RVXeutdM4WY6PzAhHNg6YN9ZJw3OGtIDDueOg//SHYhDX
LlyV+N66Qk2WnUUbofj1Og9bE11l4KGgCDZUc9EVCVcFm0udOjOsHhFsXMnhj+ONOng/0C7G2m5f
yeomiazX3ptd+x85nqpP603Aob++szRxOXq5W76fp1WOVTbDQned+yAjoQ0Ggp0El2u95Vto7tcl
GoJW3XHRDMS7WXJaDFkIDSqBi+yB7NgMxvx3HEfbB4SwVASc9UwCIYKcJm4GtghWyp6i2hKs/SuI
1hSBqt8ZkX8jo5MZP+UTt/I/Bn/p3xRB2xwMR1Y5O46GE4Dww5XSXMRu9rvbSZ7n5PBjJPcyhQTw
xzS+Hi05z5eionbsb+vCJgV1uwt/zFqhJtXU/DFe65XekjJR1Quai2KGi3E90Ko2EwYlWe5M1Z03
kMgDa7vi0lJl7FQeKMYuUi5SJrxqwpGbQTlo+bryDRyMPwiDoo80ll6luFknM2s5Amma/sdWEyp0
NoFE1DxKaM1kAjcgd7Bf/nVt4fBv8pQm0OwAEzeefcdCEj3BTfCBykao1ltYCmujPemLdSb6MkHp
SVsph+xJQ3TRPi15j5t22mY9bZ+rh9a5IpeJqt3k6kSDyWT3NvcsiyExPC4slTwhh4727cvt8eAN
i7mbFobgUjKiKghyytnfV64C1v4KjkKIZloElboKR+fRf+7aMDUn4uWHY0JvKdNFsN022rYdrYPS
uF7ga/uJ3D6ElfZSKObckMB2jwj0NBlcabo2YfVdPBotVzOG4k4CSFbvKBsL+to4/tW6iaULYcE3
4AzB+QnRRCzgMxBe6PqfTQpnKYGvN/wVYvoXHAoxv/1BZ0fGk7KIR/uah+qInWtV5kq/ajE15m9G
68XJ/vEGZrNLNW0yICsI8o6/s2BahsIpIexRLJwLQISlM9Io5uUOLJcrkmnclZ0IFNAuUZymXK9S
27gTKF1hiWO/Ts+5aLIvfR948Um7F83Htaeq0fiCiSZit1AZvGZu4XcMJaVZ/hhXwh5WSJCqCH7H
D3NhN0IQakq3shl04X3DNtmOzq8ciBEwZHCHi97287VZGrc4J2HYp9lm2lwRG2vINVi1Ed+DqqHk
e7mbIHScmJcukD37X0GMS2hH2+dKDm1RWJE4yvNfyu1FDZPDkqmz0s1w2js1HadrZnUw18fQYhbf
r6aFSt8QoCAMmVhmV/C9TuaQObCZGbV6PgXT+O4pRW8qwkqjV5AZHEDCVO5Z8TFVyBwt+R03CHEu
LXsscIGjO4l8L3Cr4Fjl5H1bEqhY15n/dZUepTtx89891sjSSBd8PlHxbkDkCPFIDkb2ftOVYx+O
dPdoBFcbWjp29sKqJP3MA7+OldrASvkSgNKHC3LXxZZkLDm2JPi9vxzsHm5uIjxWTff/6ecUEXkE
i1YFpOYHzx8UEpbDP7ThMMD4VKuZ8y31APo7ERGGV3t0M0FYZk3Wx9ZJkym9iLfL/St250scGIip
p1eXKBml4Au5eJkkNx37a7m/vwEBc2VzGOolIC9zvpsHDaklnlR7xC2FYw2UUXywXO8bpVXwdtd7
rbKloUQbGqOIj+mDai7jFrNZ8M8lzXJfAJIWhOM+fiKFwRvqCrK9SQAT/XY2HQUP8Ql3Msm+7JqA
lkhoE7ewcC195K2AIbwXzpPFYPCjWfAYCht3537KIPYfa+mfOMRb+Svt9FtZJdHBszPayndMLJxC
fXLi05Pyxlboea8j0TRwXR0198c15xVGnXCoXtdcppxbmVaoU/Ba69oD/9t+zT/bHWlDEbSH8mLc
K3Q4ZkbjH0KGJvKlv/NFmkMYjRoDkj40K7gKQKQLVli8IjoRTpjQYzLUQTjFQsEBihRh1raaol20
xOvI1w2ydzHhl/B4S0AwFvsLf5NWRVNEjUFXyw736CUZZKX9iGFtmRNrGs10AcaRb7pIrGZ43/3h
+j5QPbG8NpqrHm1tEEtGEePf1wxCdItRauT1cymznZqXQU5lZ6C1BcaAt38bfyuzYfzqYWNvOa3b
2mWfh8shWMtm73R+T9ww3iofPXmDnVV7Qz8tf1U0QL8e4sAh7SG3dYQPZduC0yQvNhg4bge9PgCI
ZHQeUdChxa+lmPDtl0sM3sYfMBpwk1tXb4qvRp3Nwx8I+tChM994rlPj2AvF24SUfKDfOtVCdn1O
NaN6xE7LEP2RP05RcNvWw9s0cinR8w4gRzUJi4sdmJSkKAc1nLng6VobpfARuxLJoiL1ql+6kuYa
Qh/tONZM6ary/mm7jXRjtunZ1U6QZaDfR4++/lNf0SIi/Xho2yyjeyZtKQu9LgBt9EXIRkxiBhIX
HwBVSSpLDQXS0fk2kwDSjdJEBouphspiJH37B8DV1gRvcwgvqJmf4FAeJcPSPx3mYFcE+LYH3+Re
YlDMMdM4su6HphBuBjnyH+0+Yb6hG/g/rhrMT5PkoP8gNTwuDYNVvSdjzeP9ltSAB7eJehNQGIjZ
5un10KCeLyPW4zxRlEEHcLau7f3wQE2vJD9nGZB1Xr71ElGZ41JfKNJZyLeNnXYxKCCiq5zaRWoP
uWbJrurRI1Zmup9fOmYBLHDyVBeNA8/ZT/81gOb52fSLRNXEfSE6JYyXOv3dh7Fgw5+FYfkyDJDq
FXnM08o50EycA2dDT3BqDSH7Qr81G2sJb25nPC/T721tg/A3zB0L7egN74Uli8hg14BTiJEWzBZg
Clfxkas0xt75Ek8twN9LwDkxV14U1Os1U2FDMqyhXuVqBnq7B3Odj3Ox/nMuRqWpIBMJ1HV+ekl2
k+D3MB1HGZX84OP5wNmhZf3Tm3hvi2y9tNpFowRY9i24y5NgygSwMqXW7M9z8DonYG0AoXC1AUUK
4ExBnYxLX/DWa4i7j6eD83p8T2m+1GW3eB2VESS7xt5DKxHqfgRCgjx21EeTsPqEX1BVs41x6Ftv
fKyBLASF6Nb907ZBlRZ8jKGeaZZJf+CVmnkaZCi+X2gor6WS0vYbovH9nJVJcms25nw1x21Eots6
MG1pCZY+j/btZtD8FOjAt9XaHHDX/0fMuxaQHFOCot5w0UtrEjYMLiigpq2HNiE4QqE5akB9sEoC
GATC0LWiAnFtDQ9aKmn+6tkBMk/Gw1vsc63S8p+i4zoZN+16/wzM1uIjd3T7nQFny4mU0rw0xXi0
E3G6cevz7ncNMxRDs7K97Sij1TCa2sUJsw3easpbIibhmSzcQ6ITAZP5HxkgBvrgu9ZCvaWSTZf7
6oBfF/WtSjD4S1+zZnSFxJrJBOHK/tMpm0pNNdfGAovg0kDotXbifqMK40aaomlvpSZhPSmDxRvX
ejuc3Kk5nT/jYh8IP8WCtKj+yrf9LNe5TkCKcM50shsxSjAi6p+95I7ujYoZqIbZ6EFoP6jhqQpI
7XxrPjNo1V0j34xpKD3H0c55uTaSfoYmkWdjNur3mE2SyBL0p4+0BC9w6w3nGonvveBQroslpZlR
rmYFY6dfky2emsj6cPFMcQ16sLC9xpR6VZOLR9Ss9f+fzEz2togfHBUgO4RMf3m0U17WGcSgwzRA
hUczNUCzS0ZG1FpdoXb+AwnzfuGHjGED2+C7ER4NUdXjOsXLVZtqduBo6xKERhqPJ3ylSB7wBH+f
B1IZH4UaozJ9rBggr4EuovJ2xCrsLjjN6MXWaPLvJDgog8btZP4VWOa0UMDGsD/vRjjCe02TVTb4
BfVkKKm/sMm0zAcrK60ezEFytfHaHDfVIHemyjVdSBUofn4NjhmNlmdHg8XtnoDwnpJ0LdYEyhLn
WW31yWyxix1vWy3UJtSTotCQ7jF06cgZTZXoy3DWtpPhDBM2eGUTfIMOppuG6oFwDLIcalHeKKRX
inCRF5Lsmvy4WRumoo0zac6khKhj4KcVzHlU3hDD0bLctCh1ABduP1xl3DxHeR1+H4TpfNTIdcKu
KJ1iI0HLaUrMnNS06bYolX93SlyyQ0qPWLUcQtKyX/ZIh3w3PewfvHlJacOe1CAY3kpuXrV+TmTm
g7xvvrNc1L4BWmJXCAXhfqWE7m49MYeuYn+6vQQa/4QYIi8KFt8MTtaR/WIFYae0K4K1w9zSh6U6
IOqk1YyadBa7Lvb1WMgHcqmFyCDDGLddBiahPqseZytDfIbZpbJd6o85Wgd+l+bRf1neztMf5HHv
9D4bZVaEEOvEa7TJ/ni+T/sokFgPZvylJ9PSSgBsXkxaTMOEyYCC+K3AscUE/2V4AqsJKKG0rRNT
jGOLxMnMrjnt6W8xJfdbheRrCZBAurJiOV8rD6GpC6EyFoRgHye8UyDEJUh5iz4iNTjWvk9R9vCx
vrAoCS4KMNzhWLTHTaYzyWypjZOsrgTMJsKp+VVG1ionYLpHhJHsE20OMr62dDlKz2mhpjXsU8we
Lra3/HsVfBTYWC1harbakWBok4OWIRZh1Av+FfcCeQ6iYPMpTndz4Qd3qZzY31w5fkzGxcArxbFl
sVfA6JFqsZhuw1zh25/AHU4nraWzXtxqSlg4p4ll1CtTBMoMGMNkewcPNOUoj/uxR+qdwccgeaBP
XExFKVZ1JaRV009yQNdR54HXb6DiS8oftODmKLxjUUt4JCfdIMBsCmJSmx8o6aAIbCq2j6DWCCyp
w5L/Dx1mDuDnwJVQL89HWlOyjgpkfh4KLbgNIHPpUWleKGhk4h2pbCBdo0SoK7Orwnolf8VF7f3Q
OzBKPqC9eGW+XZAqanvvgSTPCcHwETopd42RYOd4t83loVUMJUFGafHrdjJSLp+nf6WPGB2UvTU2
7d43JWogh5G2ADM6rC7pKm3BZElzgvxWtCtxNYA8lHzNflpjqIa+dzeBXVvYzyTYF7KyxXiAH5WS
fKoAeBcU5OhHKXLny0r287/TIKeyTCqWxuPFUCuSOJTPZ++IcydXc0Tc/5RBBP9tnM0yt4pqE0YQ
xUiV+Xix6K7ccnBsbb+G2KlQ6N98MALPa6jFmw400taXVryEPYNpsvjC7oICOEWazxX8Fgwry1lc
7hCDp3wH/xe4WEOn983sQZ3ETnJ7J0O0uB7vtcIZRPPa+D+qmIIbHdtl1/0is2d2EFobapJ+LMfI
Axqm+LfWP2qwTqb+seUUB+0WHLAU+/PgY/MR2+GYfnTMueOV6njyEvnk5dHi2GZfr0xa2La4XXIp
l48E7HW2ym2Tr+j5vKQWfPGZ+JzZvm0ZnU52vqB+Kif3yTKUOdkTm0QJv0VGb0FAMr6QhM2LuQF/
5CSez2+LYcAAa9mwrIt6jAR50UVdPrDw2ofux7EaZTZwkCDq9tyInw17BuvtAIZup+ICUQdq5/TA
PYoXSAOazUrKlkO0bJnLzOuO5ztaKGmUa85RIfn+i+I5rdr4IS1APsnm5IdC1UsMWBJsw8lr7eAH
RQpq7KVTErsH2+RAaeYLhkKBOsK9EnjRHBjJHg6+qWAvf75kl8BMKreNG/5hsgIl3yMFhoqsZNy0
iQEgClwwnBtSP5jJdmmuy1ISiM8zUwuWWOr26SAPVrDNp2LjGziPF4thOTtQ8lMnpLHsidsNrfVp
1hBd/vaLLNW64tIAWyDnCjXyzMy4OVdCN7xapvRcRPyJU8clXroyQwsF1URoQH6DsJL6K4Yc/V21
pl/0gLD4fokt/vEYRClLASmHAR10C+xUt6h4BfRNTBC7PiMdp72/zr7wgs61sfaJ0Saulb4+ZXGZ
QAbesGflwgonb7V//fyRtOFlnxjr7/Dh2enzAzxgGoRTum+nyPe3r83v9aVotVi1A7RhbHogx/TY
tWNi/m5gQvC+qfUtOv0oKZEQ1qswn7qK1Qu2uwoOA4c070WZkjvrarlzqX9Iel+oabJXClg0e1vt
NksrN9J340+RWB4+b0uulzWn/io+wWFEyLwkud/TMjCZgR9l0RTZCTbSpAxzo62ELbpOKt4BaErh
lVXtyednJwgqvm/FDHXO/tX9iejUTWBkM4/lo7R1qRx9g9cErtrO+CegFZYh09Kpxjwu2VXFg3MW
Ac3W9I3iRpS6SWuCrzITrkSZutRdjLGebGi5t6djQINeP7bPtrJGeoHoUw/STm8KQg7VTL0fPi6z
QlzGvzPxKrBghEAZ+p9SPJfMTY3JRyJO7Ga1RLkgjITIamegeqbKnn9dlgS+wIx1M70ua1QnPc7G
0bkS5O+eR6c5f4Bf2e1bULjEusDKvlC2C2OUvu7BPpbmnmBfD09qUbHPa3N4eXEOecnz8hwnDqzT
KUoRJBpqk+X6cYhJN3vezVLgmByko4genWiKAvSrb0V4/F5UCb/YC71F3Qn341ipincCHIePWKp2
erfxN9Anko/rtShHyM5OtCeDdKdau2lc94w1CsoWmL3ozD+NwunU/XFXmd5ki8VEORoubbtT5zkj
h/5XNumPSanRn9CLjiNt/BTdlkRXBqDh0b+LY8oD7l0MZP2QzfqsDzTsMcMRMcUPRRg+1A8ZTy4+
dkXC01mGqC1LGCDSGFdyIkGavaoHOmL2uuUqIZFEMihVR8CSS83XWigcZpBQlohM4TmcRa3vPPt1
Am7ilm+4UBXpO8CBIgVHpKv2Al+yuP2FnZaSJCgHPIfHyyW8qEwh9GDJFAMVGpknB/1WuSmwZyQ2
ASJKl2LKwhtRghPiRzDxTbufl5jKUpCyyaghOX9X9HxE0O4iwl8UIyJPOvnh36P+mV9CR7QAKSz/
exHCpb6KKHKD9NBrhu9ynFH/th4KSMgcEvXLB27e2yt9WzklE6Jumwft68Ps80bj9FAIw0zFN4Bb
KzsbCbFCBFCpjjBeYU2dGiNAKMru8VAhY0/LlIN24x2oRNNvwvtv3sNIaRU/pmZ/aWMttqKKZGek
T0aQVI8HZFwClm9T3WwTYzZTC2o8K2waaU5QFbbpMvcRYDlsypA5f2aUjYp3UMs5JoSUnUKdiHKQ
QokgEzOFbDkXS6ZpalWx42lfGfnbtIMCZxKQVIe+4f8sHp/+ndaiG1qBOlRzgX3Hxn+I6SfJduB4
o/xW2gRfCfSFkub00DKD3wlbpDJ2lPZxjT7rr7UruWhsArsGAkCogdq/fpunSJzxB6WskPNf/+B/
m30BwFi1NZBxQ03UrWjCujXIkSEXHB0HFram+nHbnnIXUMavv5Ltu5lr9IsRZnm8UVbAVVIO891j
+opgGn2y/pAIvTULdrIyOM1Iz0TjutIel5A/nMp+6hGl+JFXToegAGjjjyTDhAihQkwguPyMpPig
bK1U4h5+bwzsuVX9SgnmLWfSYGcgdmqhC6SRVPIrNW9rmJ9xWzEJ/z+DzgWaur583WmREK8rvxm0
VfTemfu5Suoe2JrakDt/95QkjOAtx7J6H5pKP9wYEaMzwpZ8U0VU8DXYCHHhr44Lq6rUgZlAhkjh
DS6aA/pFUC1PCy7C9aWVsbYliyEYbsESR7wzbQmfWARb1u5wEedXJPr7FwQiwrn3hXv4iJmXvyNY
jDT95fHFqyUHoTi+eb5WR/10w4bI5K91W5l5m+z5QqEXNeYtLYgM+qeUpT+DcJfQvfXxKhhhPPwf
b6bACZJrh51rdxEHuYSKlE9bA5fyf91qsZBWyhfm1an3zdG2eX39FMMZsQ95ujYwBZNIxd3Mcx9R
/MG2Pr98VI0yWdHmrCYTCCNIcZWDW+b4bWlnJIEScZYkrQvSpd2a49VZnc1e+etknm7TNCJvRAOg
+E0NRj37ths9f9lTPPfywluVvWxqWmhK5ebdFqBKsi2oxfszueO4XlCDqnpzvg800ZX/QgPzr0zH
5CJ5KZiCAeDxwGulfduuWGNdRXqSsYbNPCUw3EKc1nMhKwKkrcqWHlLHZo6rBhzdFAg3eKfSd1VY
ROxF1niP2Zf8zsKhBWJL++mTotuczLkgoOiq4wJqEr+4PoDkRM11CBW8k4ePiEY+hS8dHJLRZJlX
u+IFBobb1v9fUrzsOUSMlJNOOl/yDNtn5byGiWfFOjIom8WnhlquyF6dX+f2zJ0M1ISzbLsAwwX0
jDbBy/UvKRBX8gSwPz39UVEdRl6gytWZxSs6XTqm7641dDqLsbl5dDTsbsIyugeXQH8c4v7VQKCI
f8w7mG2L3IiSp9F/FcrfHydoC6U+K3iMcMJpD2v0rcmy93PjkTXG8Bttm3SbkTorMYAds1YJnyO8
vwR9S479CEqU3x72btRfxi6kpJvN6yZDfVZYpNJWUgpD9c4qscmZlJ8gkZd0j+U2SohyGbWxdnAe
27yukvkhSY5sH1F3+ObKlZo0lcXrTx1Mptor7bTpI+EBiYuOXAle0lHonkciFyx2T3k/qboPqJxW
Oe+rI6B498AxblKuhvVvUfxGCb+4QIiDpBmNsRAmZve4dorZLoVTnpM3bvf58Czr4oRr/IP3/5vT
HAFw7qX0ej/ClomS5CRynY4VFvPzYRX+67XBcE9Fz5gzrCpVFRz7ZKMChc3iwXH6ONviKEXSFOz5
JK1H5YTqZ5DOlMbIKev8N8VEIdxWOGWxtdhXsBgfq2AtsZ83ne6Y9soNti1JrJqz63+zN6A7gD5i
HP9y8A89pVW7GQWbGfttnC3D7hqTj3Tv/vbpRS+vM+17DqcKjT6/rE3NFTc1hYqxrWy9yB0xsBG5
HuWuHBE9L5T9jJhmSO+z5ta1BqYJqwirLkHEu1D+82kVoSVhL9erRycrK5Q2sy/7FETt9tr1PSRP
gHmJdLZBJ5jtgOCyNV2IoAA0MFbWYUTgFOvlSdiKjDKMmGoMd/2pjZUmR0JJZR1dTooo04F1NHZY
4PSQJ3U5od6jI83Q4HMT/FQ5UdiJYUswIwcnhRiZARGjAy/uZqAhUfiU3MTtPc85gljVd3JbqBop
Fkw6hvoKNjgyFmfog2NPTLjW97ZBOK/hLci2BF0PRFrWRJY4w9VfPZ3q2j8bqev0eexldGmhZahl
ZJVY6VaL2OgRX/SUkS/K3cfXPW/cMWtnu8oCoGuXYycPzt0iD0XVsCvksK4pxpzw18viSAazowiw
fk2bDvbVutbn1ehpWkbTiSo7QobfHAJcA+PhIYCfaaUAEOQAQNFUG7KuaDNiopJBR7DuIv/qx/R6
O6n1nii8l0JVpj3dtNfojYeoFYxihBMje+fl5GEAy+304RuWAHuiAPwz2aPJ1G4G9jsQfJnhvxPs
f/xFt8Kgy16OaWsx1FY3cNem5+FJQuHow8fZT1oKzd/YDgMj7rdqbAb0qBFaeLq/WbiYwWF/NkZq
qIxPf7Q8e+yZyw1hLVHN8ta7eMqJbwqdQvnoPm4y7BYZx9YsbDDgcHD5Y6YoAXONLl7AhdbHy2ZJ
zLOxBjZkCF7usnpMCgRkJj/qjXyK6mk8Wv480j6RBImMkjIu6b8+eV4P9UyXVnPUwt4ow3mvVHC0
dJMQO5r6QqH+6Q17kGv+ej5Ww/jSV7MW+ZdSQSw1lqSuvgzAsesELnejUZeigVGuG7Yxycu/Tk4n
ZRbxvDqxhCBp/DMQ9+EY5PtfRbnrcNFT8NpnoJLkVscTCcWNT96DhwAKs1gLmVfy8YAxConP3FMC
ra/1HVf8BEb/PjmLdCFDJrtavZi6Uled5Q71eGYhO9GKAhaXBak6zffnUcaKPCpV08Vb+ox10Dzn
Z9MeM/pN19GKfnPdL/vDZtZz0BGFjQNNYigt54IZzAkiK6rkoD3xAebRjUTH9jVX+lDLUnz7CX/p
URkNTeTC1/22cnTafxU3/O5iffD2m/CbIhkrySPQDp16yMv16ujJu4PbGvApgXOuK82eysc2ZM1T
Jo6V3QXTKlmk0cCGi9+d3E/Joux53uxvoQpl9NKnQViKajb1Ewcr2W0sf9KUDVCqo+c+1JNajGt0
tYsAwn8UKU0q38BlAt0ROhIytR5vuPpynbthuzszCyfBdgZ+kmvdpVDCTM1Xvr5CQnM2jyi9s3sM
js9ms4bJpcrKxZ7oa7igET1oWyK7sINu3mUxQDFWr3rvUYT2BSpSPe9Y+d84CUKAslO3PT/mVzG2
o6+FpRxxdRDl8960z7g9BnbqddpFo8/KxgJg4TSAW8bdgz1Od1yNF3FPTvnnGTJiBXlHA9eWSE1a
g+l73mTGGMw5oS7xZ7Pj9nZbsG/KR5Ko0GYH2jAHy6G6oTS14O0h0tDnAfKj7u1lWQmQYFinN63b
BICYm/jzZW+5ETNtI+ZR4xfL9n+dcMh/oTC53AG0MugVr8Z1Mt+YMucHZ442rnRX2RmrY3QSxulO
Sn51zpyhCdWcFrhP5mK2TxfU8MS7Te4Oipt1JGYHqPDHZrN6hITJiGXpwFRay1K2V3X+SfL5qQaS
x+XpQ8zbaFJDRF7Gi0IHkuPg3wOtYk0ta7274PW4f8rNnQNkx3dR2Ur7DK7CT2jff+NZ2i8/wbEM
KqHEGvm5tnUBqor6DmmLnedAqKFtvfaxkbH+zCn6G4RcFVO71gc4e2TLRovgcImX8OgpWg5tXJJO
IdRnE+qbzOhM8ZkUBYgGYPINfZEAYqgU0khS4QEl4ITSori2HSX15AfNB6yMfaqEklygou91S6cW
teun1iAjq5PPOIkeg3AVoSObTZFi/g76zdnuX/0EwcGryl0Cwyf8BsvGq2CZuh62OFAbpxCzxsCC
oOfznOexZljGFm2GQ/F1UeQ7F37PjkIpUxt5zWaCwfgvEAGXGMdrUjV6W70MMrbpBLw9GMLOQbNt
7jpPekVu2/B7Npc2wP0JDgiPFZp4tEzABnQr1slMCGUsBhi7Qmhsv5OU+T6FpT46XpGnc35XFyEA
ZEEP+hgoK+kFM1dbUzEDzYm2MORUFFFec7rO5um+s3RYn2Hx2/KB5wEQdG+3cZdiMaHGmaABT+zi
fJ+uvkN4Cpbj0jlHMPVaA9VnG4HUlU7cm7su5j4or84wjVzwsIZ42FrXjxrKfbeUAwfc2nTpFt0J
PmpuxiVrdK2HE4Ab6oiYKwNcx2kGWXCZTmd5UB/D+DN/0e3OeqFNMX48IviJjNq27BLcRTdN0Np3
1iheVjQjISZ6lQzOaBuVBCX7PD1FR0jGQ+i/FdNPwzjDwKoxeFzzPXg9GOxn8oltJerGa4j+W9TP
q98DBd7glIC3lxOZigwu7cl0t0QnHF2ncujlo2YjkTtWWkDZzrCuGc8tJMJRaIlhzw2+bTtvIDao
WLDe1v9GpoT/0rw05kmZphDyuuuJZMDfotzbzRSsXw4QMPiMjYoKqD7zjXt7q8RNZ+pHJfKXAGry
MPtNMzfotO9RwhjEgQcK9M1MtgaR7ixcVgqdf9IOar3toy6og68Ys8rH4Qb5ajrzvzwvSJYZOvwR
UWRSuU1BHbV56mbZrsOEsmxBEEd3eqGaCFmu0yn9HBiwhd4h/U6+mC2ke+GS99Nl+pX97UcLzfA1
wi7ET97iyqOotroPugY2bPfaQaZsOsDfF3HrKSsOyInhRX95+fWflPDE+yYBavZeuhrDMt7XD/ua
DVLRWoryi4Ir8LWmFqOA1/uJjAf9qeg6X3Lhdnd24fPW9YLRXp1jx0Ss4xglc5yxhwP2cbSUmeQw
UE/HNRR3Izsfxw+ilpKq2akqVAlgIlZQmZ6a6xB6J9numqBG5M26CxYAdsnknbgckGNyu+HubLYS
9FrtltJo5mEvbpEhsb66dR/4pb6G7ksJsEhAtuRP1OlyDkU0+MHlPsX4g47nqYnWD02nvf8ych+B
8w2jmkGAkid97LthlY0muUzvpA6UpsN0l261fz0venDh+MObwRhKzkcsJMF9s4HzL2IhiZU/os8R
SH5skE/Bjt5+0LKmEyY8mDssa3WZcZBjxd1ueUYBhg01s/DJV2I4+4Mu1kCjf+uENyXpa74m9woy
EAFKi/Q3bO1EWSF5lgg3Gsquyu1PmfdgTBWRra6Npv325l7LwHhmcBZEQjVruTLRxDy3smbactTi
y9d95tq/RoScRiVJ1J2xntdBksOCpN/n7WOBoSwKsMdDPmyPRE6fqRM3Uzn99zKS7mOciJtplZlq
8kr9YtAKzVyiMHA1VENMVaqzZ1AHYXgDtrcCjKffvcR5TuRyNaGAJiwRZBOOJKtRevksnJrMl0rY
IiYdhg68TBBXmuRc466c5OUIjH5uXragRODgNgVl7A+iNjoosdlq7SYeu5TZgZwY4JyAwOJjzi2A
/uP9PR5Klq5FCh2+ZKo4xcBXQlxDWUVrL5+TshB6ZCnquY/fht7Eqy3ki2uZv9XHM9edsWevsfFz
ddHgbruoidBEgjOc+ZtM6VdvClLOyAJRK8DNYpm59p5iWQ/rwlvGRfS/b2KHP9O0Saj9E0a/DGpk
51uiWOhG+IeaZ3E6MHC5QN/X71E+ynC57Y33Cn23DODiz+giMdN7YzH2mw7R/wdXwLWLl73929tQ
O2h27BHK+fvGjpAW0ibnVeuQkwJfWUyHpcTf94SQb+1AUVsV1gWRSnKk2G7mu25TSXweFW1rrrP0
qEhJlINRsBo/bK5+IqSSaJezryNU8SyAJIYvRe4SkYSzKeMM1haxQGarVuELkIdCGKr2rrMHfP0E
SgM94a8bbAUsTDl/p1TocfZxxX0Dwdpne+c3BxJtgALRJ1EFramn3Mu/HJVQo4reTysfNE/khNPt
kwD0kynzsLrcseYxvooLjbPRj6BiBcENjzZx/PwLkFQP7z6mRwLpL1sP4Gt5H4ehJrp88jv0xGJE
/Ax3ZMWAavwAIAaODdvglX7d8UX7Dmv4f3q7VrT2PwzTGx2yhLVnvPypJ1CRspH4fE6awMoOIVAP
AFb9YpkI7BhAEg5oYkQnoH2KxEHZ5im1lP6Eq2g/TP/316WMTgWZlSzhHbfLxfL7JFGqdSEF8RJH
1xkuCP8i6Us7u8CZuqxskfE8+ZtwiBBBXc6Dgt06vwQXa/jkijgPv0F62G9KXUESaxsnG7Bbrg7F
qiv+1CZwGdjlNmjNBoaL0+/4keaV0CzTX9Ze+Kz7wnG1n6ZQNTuPzLgDU6jaS1nrpXTVZuj/1tqQ
YZmNAYyETCx0cfjKpptYvBVpRPKBBixTMmYC3BzSZvxaBE3cJ8THK+GQOR8wBPcwjuWbSCeF56OR
S2BBBONGn8YJNSU/CMQgPtFH5h+mLbT3Q0hr7yfsiHlJODwnccAfAlEbtZjXf5QDgc4idkWFZlJ9
2vNKv4ElwY3Oc2gLIz+JYj+9kwmNp2Bq8d0GlG+7yNR/JG764Jn1w8+rWSQfSt6nJ3FIYX1LXUS1
2P4khcdxSdrL/vEuXdWyHgNbXy6R/S6dYUNKC2n+0BmWyeLaPxHfB/HB4qWKz1gtEmK5IFcU/XaA
WbA3e0inGjUebUOh8+Ae9G0GjOIwxIK5iy+JMKmXeDza5bUZEMKuNtlZ/37RY7lL4iX1MF9NSC08
hrcsIl8T+8VC1T/+p+ehpJ1xii2UiFjHXDe3wYcj7ZeGhdgT/rwB7FJ/+M4jJT2FC+zJ6U7E1eBP
7lP8ii0ZBUpn0+MKxCTZW0XCyEPDt/Q53zyRUSKTN3WFmEoAiniZ/mRZtMnnvpUAN+tsllaHAXkQ
TtZtsAtALzB7V+pOyln8mNyAR7u/P63Ryw5unB7NMlawN3qHwHMLZg89VaWmoN4qOFISVbxS0kdx
sk/ORxZbplqx9AOVjEwlX0Tu5Jkch4gyoMYibZxG+mcHQuq6bTHlNh5AxJkQ2dKonfj5+T9pKyhR
+HevFauOa9QNbUT4MLq1EGfDY/1J2u/FTKVuYqbetblQc50gLVTJa//aONXPV2PIE5sgwXyWWbsU
FLYnRjLbhBuTrmr4Z9S21wpLYdvi6livUCF7twx1WXypbmtKH+w7iLWVg8Lqk3VO3OslAze8miYp
mVZx5j+EP6z6IDyGRnHXXG4bPCM32uqKgoWDdxEByREEEjAwKa0pu3c1iiXP5ol3tU79nIqvKZF+
EAHRf8cKHemcjYAzGOTz4DIOWTUyL8P+nT8Kj9a9yV81JGg/VHeAPBSVoyoUrUozNmTChjEjvcpK
s23kWcIGjAgaJLh6jjWlEmNYlC/LD+9VvbQ4SN3s36H/3EcETIlOf4pRLDQcUzhPl19Bkol7AzKP
JqbukQ6PDFZn/zuVs76WtbhdJHR6N8ygUE8zi1uzrLiSPi1OIb51aT02ranFCpG3pZmpCZXs1G0g
IbbhftYwAG1C0PW+stHQb20m1yv8qAuLalYUPhW7j2Bci2IXcWvVgC7m9zdo/n/aKDndBADwoFxF
9oEdqgJ++bdeHU89qqxhSfHbIRB6ooIbAeD5XkmCyVYlCghQ8Y4Vtv6TZ0kKhiHiN3f4s04VVFmi
5rHBNjo0kxZEv/tp0nlGbGnA7KY9otg9OVEEak1/+gFgAhW0VOq0udRlc8F34cuxya8haJWPyKCf
LNNMmLHVwkVc7xhr/Aog37Xe+hx2M6wrlmvMUx1QzktOnXyF19OgjSlIcgqCyLl2SzwKsrcNZIRt
GiwUMOVDBXKjz3pz+CHMCWSdfQ8vH0z4SvoX+raHS39dcDU0OSvP6/GFcZMia4Tiiy+B+ubNbV/i
AOoW0DnJQQFKa8eKrTmcW1Cmr7VnsS1Bdh3uZi+dyILCAjQ5iBVj1BV98z4LD5R/7trleI2MdyVz
KUIEIlYwqXOFiKEbkzLzxxKDJ9eHdGf35wmwWykZ6bDFnyzv+3sjYOCAT3529qmmk5PQzwVYEbwT
Ju0rG8hcqNlf/FckQ9MigpVf3HjXqrdpbGPKVcWCJfKu6Iv/bRg9iT5j/mBpNDnqMaejpMv5K7cm
kQis4BvEYtQEdWndpwf2nayOBaqN+oeGVNEiTUbLfC1bvLX5t8vU3gZ6LgtAfu3/wHLRLU5wHlSn
bpHruxwosfZ9YfMl3Qakyq8SLqe0A/qt49Dm3/Yl2NmGZT9MhgsRmi9MFruH0KyFpb/rpwis5v36
pTRIzBUsIPENtKswhGyiqjvNezurjFGnU3EqUGfCxOTyAtAbgTo363hqGPDNqbWporrCp/SSq/wI
pXLB3WI0L19/yQEYZR0BP2YhzIDPKnMNMRR1FOAqG2m8q/mFQXIJZv2Y+72lVxs01XuoOBhv/y0/
NhzJZcdEk4irpRCb+n9NrsXu8bkF++i3gqU3i8W7QW0DicDYNWsNT190PEptxXvlYAqfQviLDVE9
WG5WEhrESVVoTCN3d6NoaQLafD/Gov/s40L124Bb/BSyQ1Mgn1jbL8EHvMZWMZisKpifQo9q6pdm
KUXcbvovoYU0byU9KCAzIZ8RNi+kM4f45IkrAFa7oiHqfGt8NgKjWDXQMSdNSgJQjYB6KwFG0EIq
t3hYsioBOB0axARw3bL87fS7+9Z1zFCEetEPK9/1OwKuFreSsNyCUyAHcGZ+JKmHWNkr7KfaFFku
H8nQlwX93rxNwdMQly4OG+CVLvk0V+F2DNhNlSxxJO6zzrwXj72uLFY6HCBL9+8De/eyw35iFkVy
QUJN39eJNumVkXXIEeOEr4kPCaSiJ6eIAE+wEGplgQOPrO3MoNdie9L/IbbXoNiAgn/nhetc+eGk
tNfsu3dtW3GlOcCCwN2H2o0/zXMh/HKfPH3HqRXO9935WP54Hn8MdxY9+9hOqrQjJgEgebcGg/e1
KalfGKE9LiVhb8HFKXJyhZQlqee92AP7y0bwCfChdtWI7vHkKOMRp/dL/ezAps6G+2tCSb8YkdZk
SPIC5pdvskCJWRNF8NRThnAc/AEWwAslsZXt6Kyu5IneqEDSnuNbKu6710eqkjv87MEStC91k5Vo
xnR+4c9pM6YtbRvgdkTNCkcrYb96v8f07Q6kIp1BlbR1mxZupMIDJxaKGPm34CW0o6L5fyjQN20p
e8jVwXLURVVU8davGd6PthieVWHF6AlV4zkJDMqbRdbBx0ymOFDryYyjPQTNum/YuJRp+8RaKFz+
tEUgHlNVEE6NNeCcRFp3aKAsDmQcnLgG7N+efaAh7j5OoqSHBywZxkh9yu1VYU7TogphHRr2yEwq
R/lMALw2e/SB+FLaWNKDli9EiWnrSLTpbFDOTivWziHFzVysaMXnYhX44oF4JJshUMS3zlbiniAk
IFPUQBe+vU4ZRESMASEkZ9mS7dyfddffsHg4SwE3S6mSP/t+oOUbgznHSf1/o6sGEfXE8FFebihd
rAZsP+8BmpPYRjQZzYyqHOmnSzawSJpVn7eGpSp9N/E6XvtVo1C36A2VzlrUOPwlnZXB5w6wPbl0
mbA8YMzx9gqPipucw+Mw+VQaqWnzilFYB1rwUcc9O5cczv7137OzNNuxLILMSo59jvkqTHkGSr1p
d+SUW8lFIsP5AYTVfjm2r/7ky0gVD0M3Ds5CwauBT4IQbv+YzdhPaMmwlFyUrK7y0/H4BxT2hdFk
pGPkJwgea3N1bQDRe+NY2lkgXikJXJdYMwExQ23b0wsaXNP1iAGrIOHdw27uEKEus2VBjin12Gch
kNIh8wt5aF+W/Hp301k1aA4JzOWXNr0jzRVqds8uh77QoSzG7peC7dkyOWtvRkx1RX2SfMOqga1j
AH3FxgI/Czk0AHiQm4Wn/K1LnP+eIIwSiSxFXPgZsuC40dmVQTTl3xBR+J+8lGKlFlI3vzP+U4je
hScKKaYOSFAYlKOys2XCHu/HkrTSGjXDd8CFF+09TIFCy1p8vaz/ehlZ/yNu9WTURdSyX1SZvGU4
pc7SpcuRxogH8sZYQ7wLg2poHR4P3FYY2pMhFF2ZeDGzzZVDv/ngzHoi+afEN/Xrsdvmo99dcio0
YysZB94L4/OZLtfCgjtx0XJ3Uakw+HXHKxkDI+MVaIgtMwN4vvKonVm3HgNoss2NvFKmkBq/iApP
iSj1xdXtveZY6Ll2E2giijJVQTEOc/YDldcBJ3G32ff7fAydMVoIc/NomPd1/dMlZthWM2C/oiB9
nPSyVJ71hzRLk9Ik54DKWmIkHudTmkxYHUlXlC9sANRt3xXuzPELQziYCcVEM5kqN9Y65FXARNSQ
lGlwbtCUxV+erMyi1cC3mppd0kMOiUwbYCstpiK7QaEKNck8mvXFn6aPAEA7xE3p2E/CkAIwDhb1
d+NeUMs5nOudqBkROzwUX+sPO8F9RA0qR+bDMHbqn84yGyDALb18MRYiq0mFcCBeNjzuotvMAKMO
PTIQvLJ5uog/810fPDFQWzNJ8M0Q5cqL3++fs48yL4RLHLh3TTmiNfd9I8tBMqSCyFxx3k1b6Uwe
TMHgIUocRhwoeHQPFqwRKl43ZV0fveEzOwn0KeyT6vgV2oz445Hz57NoJm/Y0lhip+vBR6JDKzo/
A0z07QQGDuWwvqp69MSEYJZOhEmhsX1rmGIHyJY4yIAxgkFmfv1I9PEdhE/iOSwmJLFPBUeNtwFn
QKkemLxhpU2yLr2XaJxSpekaA30/1mspToQxh+9N88ylnAkWXbBiHnYnykwDydgesrO1nAFXZRrf
sRnH2PbkNTihDIgH+HI6wR8ZltQHN3unAjOCTm8E042FbIL+DB+4MIWtMUG3/rZsnPxwesoxHcUH
PBKBKGQSIfEDt4MvM0zLDupN2tWUXY0LxS7Grh7gWnujDx6rYN5hdJUgYo+ELjI3cqYlTSJ7MQcF
zb2+1AL6OMsu/FKHCnt5VFwVH/k48I0XltpNx12U5FmaQHF89/pweYEvSA5DnzMiQtG/pYpv+V33
6niJnP62uNu68+CZgKWiXtYRCdojbbE45TyZQBz/KbK/CHwCdTTCP+974mXUDAnzGrpK0gyvzHrb
tvk5CBqXohJhGwiUhJUuf7paaxHI6X+q54cuu2eShoGXC/pD5f+Mtk7OseNUAhdz788LiXoL0Taq
QyJKZO5P8judzxJ8dga1Jb8mEtTYNA55c3n3pgUQanW28gJ4wHD7YRKmKWZNxGBCM8XDfdK871jQ
rIkQFAEwz1uwnUdN3zL9SxfEAWGMlI//mSrE9jg+SMs/nD0FCYlvhSlk/e/JQxmdTFFafPPMb+kU
5gOk4Zh1JjxFZwQ9Ruv9k0v4rBmrCb14kGkMp8yOJZZtsjmF80ayZWz8cJmaRcM7zPQ0rGbysQUa
7aOA7R/fsXbSlkedV4C1HeGFG2CtEf/kOyfHRTaKOBN3uEJQ0jAXVmp3zFB+PuXt2eOfuwUDA8GT
Ldv5iRSAzW+mXI3VZ/nl+vpBOvBlf7oXcPEpxauOB8zlFhd9Ya/1PAY/Gk1zOA7cffXWR9sI24oh
lC55f1E2qHIkVUdwkHOP8htfqz6t54edrKww4powYc0gUd94ju/V1eD9cmsCT5lC3C3RZ7VAIklH
jyaKRBLIQ+s5tHIajU2Jw07mwBIIVkR0cOPLHhePnyFAdOu5rZ9FF/YWhUe7uBRRvxBhKcG8UxEk
/Fs0TKuyKmvZQCkXHQIXfsu5TUJ+5cCqS6WSbLU4+7cyLtAv2b0hpDpynBSXup7Q6o7fluihxjVN
YUeP71xy4KYJqrvKisL0RtR0RhBxjRsS2BJAT9kOo4Zy2qaGgR/DIMF4o2a+oCwZQFF/Ql4DGoAY
WF+g4/P3eKnbmCH3xQ0NDtEPQuzmteGVLEzakxAuQeeqwrE0kuuTDh8gfn/uvqEUHUk+4OA9xs+Y
BhpisJh0FfLR7yw6CWLm0CufnHxoPfj/7fVsg6v9N2ASgbIXbngzeF7j38mTY6N3GnGl8Zn17sDK
62R54/c8ivYLKijtc2K8BO9ckAGJ5hJAEiXVBd0zLiv/KcnWKjLoXkIRoGMm6FWApEPuxeD4T6Wf
sLpiE1difNcgqWKpB0U8csIt6KIleny7StyDbWALQBjlywwEPeeiHv0HMAydOZHl/Vv1PPlS8RVF
et+8EyepH/Zj4cuKqHWb16EJqpBaP0cyOuvnqs5lzAGzTcQv5aup43WcDrjfqXPQvxc30OCH8f1u
nc+oDiHXHta5fGDyT2a755TMLrPGExIhLbKLzxS8gxCdN9nhLd4bJf8/WOlOizbKJaMmQLZbfwxM
7HBEPiQdr1j5jaUWolwvAxR02Ld37Kl+k32vNE8jfJcO2iCOcSYrMHYmg7VunjD+mlwc7kJ7EqWB
ip9+1msM6uGD+Me6x6JSeccTsNa65aswyjWPyOr8vjuHr1C3mgwJ63NQLba6aj5+5ULYtKcO8720
TZBtgU11IbvtICqUbXe7RB35Q13jaoEi2c2WNtuhpDvCzpArlSxvBNJNFT5Bcgwjd5uSvxWa1IDi
CMkF+UHKH32fQKdh5CLVI6Zq/3qMVKUNuWtZ2vMQXtzYUSrCugs4+L9oCfeN/NyhuvEzhFOl6Fd5
JHAn2KrUBHQA+2g1vCjVZYDDwyC8EhwFkANQdyYTwbmFlqCdok/2i+1GNYSp5oqa8lHONW/vWYqD
FBBnrzSU+jCsqHeL/Y8Pw9RsiV4TBPLkG+bEOwz85UCQjo3tXm8gQ203lZ1db9YxCKTGQRCgVpD8
tEPCQyP+Y2k+1IG8niSeEtdr9UmlnQ5g4A6qQiQ9DmNdNtQzCxy9ynUOqdsXNiPxlyrGCnvfIGAg
IzOuO/ilNDtfq2jac1pEphh4vBHK8p6iqhqwArtSKC3CIcf5ShHsj0fDqvIelNE9xYbEvyzccqL1
eAZ/ma57G/AmIF26JedysU2QK4KxOUcgTgs0pg2oECnzs16kXvG2UCom/9qWGhR3PVS8Q7+DswU3
uXjtmv3SPFwqrPy5W0ZAWPlEfC3YRLJKmJdyoCWX89pSlxTqYBM5AUp4nHfHKmdNfTnLZ3XAtdxO
w71ttydHdSPZVA6gpNw/mAsh91rpYB8rXfD7n8KswdpG+RWeqpE/OKZBAhg4aU9In3v+1ZaEnCS+
l40X7TUVFOdPJOVjw97ulq5mQ29yA2dzBKU//aDliiwLcpzKSGG/BaGOzzHmPI4no4shHrg2cd+U
V7JwifxYNtf0E9NkkWaqVamJAhwKLlqHEi5Dl8G9ivWnOi1pg7UMQPFPnksc2Uod5MRmSIIOmzz+
TncSDVM4UCvvCjyYcWrjeu8myCTyENBKszvhK7wu0HSQVLluhgI/fBu3gRxqj8ec31XxWkzd69UW
LL/6Mmm/JRc99QFqf1nDLvtEUAKmVWCRCjra/35QyzCytqJi2DVuZ1A2lXYMQpI7G4it21ZxpRqS
SmGz+H000JEKx5W+P/eJyuzZzW1hHxLRAmXrEW89tNZzlAE/RBjllGz9M8s5rpgQNHDkE59CpSti
bq4O4VsGwoc38WwWel7BtOwad9GzKT/w0UT/dpk/ZRMw2M8KAvWEmJpNnuWFIXe5VJmpCFSrikU7
1JpVrEmwYT8Caeehsxo5sVhMBsXkc+1B76Du78zENkcj8dQBoc3Jb0cWi8nGcW4TKTKcGf1yPIrW
xx7nyYP2Y+x8BdVhMow8Fmo07sVXVRcT7Izha6iJLfA5z6/PsK0GHPTLJai8RCQw1IxvCkvMW6WQ
h4uctTubkxGKVhlNh55ZQ7lzByJwPsnm5nu755Iiz+rVNqzp47d2MFIRjcn8gbLeII7O1WW8fWAo
j0SIE+O58DmfJ2X4iht2z/glhuqgVXXqIcuFlLY175HX6DjmKIVeFia0YQn+qRaUmFBVDsnxLydC
lrXHBadf9hpQx2btIh1Mf3vPV+Dp+VS7m6ertnTkB9RNLQ5+lmFGVqKuG1ucrJbWZ9Xzab1apoWQ
qjzYGpJ+XvPxbv8dAF4l8hKXWzwWbI16mlxcy7lspMm8u3RbjyxcpDC8XEvU5q5ZK4V8/4ndp7et
+Y4835JB6+ESrIhbolf8N+1AAqHNU4qwfIRTSRj6s9XpMFun9BhggOfu+2S7GVBf3kKT4Ln1ohgd
x1oOCs/ibg3OuSd05nvA5qIqBKvjL/P/IIDtzFuEdhKvbcfW4RDfb/2niwgTDBJ4BAjUHMnUiT04
Qc+TQ5D539lZV8aEKbi7hz8tMZqbdc8W6DtjAc5PwrHJKKvQ5RWD5a4ez9JJY0URHH+jVtCMmTN4
i7HvPc9kT2ovQ1iuACi9El5VcsuNnP7cXbQdT/mb0Q1+ihiCEgPOlFvyVmcrySmWKAEoeHS8dt1D
RjgFrG1hbIUDoPPPqtOls45TwIuW0XsPLYBh0MGRo2fgTK9uMuQC7hd7Ie6rn9CB4z1qfoHI9XKX
eO7cmPSOrGGxVS2OWgTFjxLzMe3oy3Iz6gvTQAyjrwhDAx6Zjr2plcsr8C/pyK2nEo1X3tpRcj1m
FVgQZtd46ZUxuvXz2TMGybq/488MRoOBi5jUEl5kcixyoJzwZZToS40NY+MzzLQ6O492C7HAt3AS
OVPAlLDXeSv7WUVWV0j4GRjQWYf1/q4IzqLwDzS/W6VDtHT+hDy7wxAcfW/GLnnQbvW9KVOrSxji
E039EEWWbkj4tB6Gg+VV0rGh7aHEvnOMMLRPNpgfn1TpMyyezm75dbAgn4AWdiYx+mUdNHr+2tJU
IrxSAlGDVV9VxsKsRtkymJGIJI6H3yiSDYEbPCyo7klRH48B1r3rRSogOOKIC+WJpL64CBIctl7i
8Phqnam9KkA7Hy0s/68FL482rt58DsDo8TRYIO0G9DypVPxzTYKfwZPE2x0wJVXDVGn7+5kysN0O
Sm7fwIw9RSgT/b5a6M6xjkwuIrh/oYIeS1jpbfiGY/3Z34QIVN3mswAAGmJ47NAfujMyCbLuoQLF
QLveaJBwLErwFRMp1vttCTJ2C9tVjHI+AT7T3CfNUEbCbBcRGlkG5ccZbadUmJiqFVK6WSYDwl48
1ppl2Xs7CQbhrBubVmkWSF5rE/nGGKMid5eariTPeTL4PGrcTs3iIDIp9+ESyEh3WT6NMyYQBKcB
UOsyz05mKA2JZQxQv5AiNBHJ+MKLJTd1D8wqnNMDZ6lNycIfdQC1ecvk117KB2gvE76dAXw1bIPP
svyLVbXzRryPOopqhbgavmDOdEaEKpuDgPoNEHcS407S4Ht2L8GhkS8I0rv7HTFv27NuB/qfbjRk
IsVwUuR76VJ0u4RNCVQTsOavM9OPxnoL5RFraw64/9YeZzDipeAweHAI/pkjWlajaRbIDRIH52MH
4Nrdk4lw7xbfg211VcmFw6eWNLg9sQw/qVLKxTiImRboP+IZNe412rwIRr0+si6olhnYoiYYrn6v
oZBnYqPd1fvK7ZFIlqn5H7dbp6fXf9uZDCCQgyl8hcC7a3tVoxnrxwCochWVrWOFVzq8OfhFX1J0
jEEh0oJ1tyIfCO+CPufQjdsEA3HBcECgiqSruZzjPJk1glo1OE/fdP5FbnNqyuYzVk/jvr+v4nYz
kBXiMScFmccV1Dg9pYroQJUl7LIZxo0mAUpvRsjwqyGfpxecZMc1l0WjkYDZZsRPIy7Gda7KDwHt
Lc2WXRe5BwENE1ypLK7ErIIALLu+sBJxGksT+7Y72SfdLihsu8Qt4XIF5FHj8/Uw5t8qPl7WMd93
c+9sx59eYwDuviFy14wgPvMm+h48zPN6yASDA7JajLVvcwYN03EeUOw9RjTGgbl4PoRbiw3QqNxI
OYja8qm/LFntZTsO11m5K2juJt3Ww/M1muxlbzy/h/pNuvd5pj/ZnLatuvRHsOYSIvURRWrm+xZO
m7EL1oWqYooQ5y2b3j22490geKO5OnCDg3nwXL/E0Bsvp32pcuyfEvkj6pBk0JoL/VVuq7sIcbyy
Yso/7TSBpGf4o6HeHvq/frktDWPx1Zf0XaYiYjalSFrCBicHC/dD0KiGkgmP7AnpVIbC200JYj0u
cm9BWqLCGfpflzLDwIRCRJ176ZcwNQKy9bqIc4UoqNs1oi0tJND83QazKctY51ueuoktfBbYoBEx
zanBmGZ6fZR56lWDOdC98dy33eRRGyS5o5n0FMag/rmNzPv02LaxXQ2dtM0gmFhzpmwdgmgY6LjG
m0qoP3mIC2ELWhCUM+VL1NySVBDKkbkWNGhCA2YwrUrNALy/z1kmKGq6SSkKVPxnfXIVBFigT/f4
xN0NKWQ7wVGqHuOJiXIMpWTcKlNfgG4t12Vi8brM43WdeFiRE7ZGAOo1jhY4jzRVQAhsIl1qGfz+
F4ecZK0/HwIsxYfOz1m/N+2zdTbTidBZqQOY9L3s1osOsnEVXuxm8PM5mFifu/womT+gg8CncjPn
U7pZYEnXJqomhoFJL89vegcHKgs1SYvdMEkWDEDtrF0+k2b0BdkYx9jmEx03eb5bmKc5BIYNvumY
TPUvJJRl58F7FsOpdUAmgN/OCxMdj6JPfY0YBBWG4g0JtbBzHQElAYXUx5vESzZX6whMzB9PbVI5
/O1LBmgX+pdPONn5H+3xDWMkHhakbF94YWUwif+F0H3xNmcvZl7WKSSDKAYuFqdr+PnY6idjDH+T
+15Qtjd33CruHfsWLo50OXt3zm3m5J37Tjf2bzGEaaZeWweXVmdh4NY0dcMcwslb/cLXFRo5/akh
nOAfxBtbD7JErYJAoBBdzn06D1AhrL5bEd54w27kPEun3+ub6AzGgOFsqfD5V6e5YslQbwa546jv
Ar2cozQ8lIVIWO1tBuTDNLSB8LX9xDm12Zy/yXf+RFfuZlo9Hq9BJajhI0d2zZzMlXMR+roCklAi
ij61QSaIwJLHd6TpsxWQBdQuv5dR1sw3diXqYtmEXavhIrZSTFAIzL4OW3ky2DcxJTMsIJRxnH98
iw3EA3Frozhfp+lllTiklEG1cp7pG6vlKabPr5DOLpDg368iCkL7F8OKdFuFKT8GIOfhlILOmst7
6NDIAtoyXDEGl5IXI6bwyxwfYtFgbxwgpE/rWJasP9y7TZ0dS68MdR+rmjo39FJJu26al64G4otR
iymq+TbJSL0SjRej/7xXqg8ZqwB4EpWfQ5bYZSKFou68bs1bg6XrFOI6HMai/Jyp67M/OHYalXCB
XPA0dLjXNshmZAP8EVyzAtXCWBoDhOVs9FPbGXihErFD8rzZzBt7vu5l60AqFSSaMRV5wWm7r0VB
WaI8q0benKvTw/aI51uF8++xu0Rqoqi5Juz3oACbGXTqy62mU2uJjPXcgWsgC/XM8WeytAtplglh
+mlZpUYaFuKZItchqrEpnWoC1GTZVFGjh9VQR2He2Xvzseu4J4oZdJqpeohuohsXpznawRDtla63
0d9Oc7/homWroKxSu7C9LU/IbPezn8CSjgQ4E0HftX6O2MsGPJK0vVAECnhb5ixFHJs0ycw7vMdc
5qvtP1RrVmSj5GCsc0DCfqp2F19I0g8VwS9qH2Aj9KiH4leTvHnRzm+uhdGsO25f9+A7enL1y0BK
wMpDYl2QXr8pjgmpevrD/kN6i5ooBb9bUd5sm86tePdRFIKY6deqpzJQTrEp/HY6jPhTrcOq8v6K
dC6xAatKSIH4SdamafmihLdT9/6WZKpczC4N8ZH9tnf7D0CVUuxXXC4l/gjuT+GeDb9ks84Cm+yT
OYwz0rySrsbSYAThcxekawR5KVUHq67ExauQexyc/iCEhqcQDF1fbozVOVLJrbuYotOzPa4fqeKy
sQTvWmS1K3NvlgQiFEvILngABy56yCGXdId4JhhY4MuzWwDfm7kKUwgbETbe9bdpPj3m5B2MPlwY
Uw/t57i2Yo5UnKMx83ljV35rvUpe9urN/Q7QNGB5JGZDE1ENJEJEzT/wSFgb5JEGdgstWwbAqMRW
3cFPcF4J3i4grckZvEB/oGJC7/b7SK67sKzyXR7+9surKR2THRU4xB0M8J19cc/kRONcO/qvp4px
+XIgI4rDbOKHHR8j+q/nRuxyCVH86geRKRmxRJZ5ehBLDMg09JgnzIVI3UJRkFYbO82qqwayw6KS
WRiTsmXgMnUF78JgO7CjBQjb4+hMKNO0VyxWfDm4YSI78vzyKOIbaFhc0w5tdoqH4CtM4cFgICCt
IR4WwalCqAR7rBQ6509c6OrIpI8uLy2TyI8fq0wSGD3nJ0fht4D/8OuKtqbFSPZ6VYcsv25z8PiC
0vSklIggfYOUoeLc5Llfi0SenJP1Ygb2qc7JjBuCu2r5DKQ/x7qdgA1zm0LyEJOENnVAPM234Qpk
QEBeEPq9RfClCCBpqyZya3DkmuODelw5DGnV3T4PmXdr/JFD0dBtTp4fxCQUtjk1W7JMu695wqDU
J6JQ0aaq9W+RLTZHv4ZMTi8yVy1mPTnMKgrPYkz/NSMFSejslccdzhRsAYWecwJiv3IJ385bJfnH
knjFAUwHKCDTTtzQlIPr64PEyQ7XWxjrzbzZu5ygBXrJ0tfYtncr0WQ6iz46njKtimbRG+tFW/PM
OYs9NaGvdHKg9tBtxYYOAap91xZVTPd8kz0AO4VjTlfBHkDtocStlMzKrsR4Q7mTdcf7K+yDf036
P53MuiH0YHzZI3lFU3KCs4hZQSpp+GsFfs4XlWmjjBjdLVFwb7bGuc0WiwpAeJshZuui0/soHHWR
KeXTPlCUHEvjecDA3CDFhOO3I4444J7sNecAF2OuqTaunDA7SKLEInhNOGUkcPL9yCetgjPXb88a
mz29cL4PCdYsjxGPXzNEQ+EX6hVI6g+r9CF2VYFMz85aO6t1H6/HJk1Zc40xz83SeRa299xECdNy
dsCSt2PIB6WBiQI42ORGTGWIucSYrZFhV70jI/HWM9f/BUUuD27HGj3bYZlGZAdKex+AjLW1Q113
wPrQIaMdQzus6kEE7gdnwm+RIjqobdV0OpOFLxkBmLaYaLegMhjeIVlmNj/+vrjPDjFDLMLOZ40F
qk2tBhFAiVg2dD5Ny0Fa5mZ6C3f4Hsbgj0nqy1AO9lA9qORs4Utgc87GGA9/GfIvem0rttxGoqzX
T74JlPSD9WltRugQKNMXSh5qiLXbv3Op4j97pU1VpBwwpXAoPqObPUe08LreT47kzFJnAFGs5Q0D
pquvtWp+tb4TLxPmrZGoYPfkwjwA+UB2cCFrxFMZovztCxmkCszDd6jqhs719MZmpkH/c4CcdB+i
ANtGi6IB0Iy6+rOyIoGXkGHOShH8kS504Q1sJ3Ywd+v5vwDNHaRMuiMXPFXnKkBqR+h2Qb56Ku8N
jnbgJL4QaqPFi/xKd7QvjuSR2JiwBfpnuPnT+T0ICjOHiH7Sar3jXmgyjUVZP5C8YsRVMGVqfFS9
iV/9euyYSAoW7VwnM7CTM+p7rlolSXZG/6ITZvtpsVWp9U47AqdBwDZmhByvQ3nx2skQ/uWxr9vx
aeOOGBUuBqtqLcNYyqQVvGQJvR5DJoZDML8u0u9UXDwKscOKmrUYaCd1DGOUQCAjqBs+W91A5dOr
RNlFIs7z7FJPienXQwVaXoCWwFksXYxpejEWmLYWxuZShoHLkEFJyvyPuLSDpK4rv8S1P7mYyYih
nc+/4B3tNWRvsulBqvM5f2lvD7h04Gj4OcwZaTkuF7wl4VjL3DpYVP57qSSZB9rUtzIxTkddWrhn
O+4p5DfrYpir2wK0krQaPlDNUTlTtFpuJUV+g2ya1TdZZApHreaALHIBu/p4YM0QqOeFMKSf1RDr
xl4T9fNP5HdFZ+WE6SekgTv+u0qJ4rxCeOm8KlJUP7r39o/3l6SPmuDihyh9qj9ALfwY/nGg+llE
RKF5BQOoUQU91/GYSEGvTl4d2o3GS+zh55ldt1EQDhjenjx7WtIx1BYK1ErsVrJhRccWFXfgwgqf
zVKyc/bxAyXwOm+JrX9oepA9bcgqW4JsTg7HEK057PnYO4fTINRyV6PjBp1sz4bXB+evbwcGFGMF
aSH1iXz93p2wZNPb5T3cTPSH85HN7HJYfl1L10XFKvx5PkYPhI1XnfKNbQDtXo4tdhSOWgU7uKP/
Jm0zKDPKUvEo/HnSpTPEYURYuzaL0p1odYdQuScdYClzvi53pST6jXzGJDPdqS5BLghHwaYpnA5M
5bWrfjhbivYVYjx3Cn5XbPmCyMMJWD2s5TeMlyMqVGfBJqAfN9d1poWEstOO9gPMCLfVaiSPB7Iw
SpVS4UWfOAdh6DjnxVgT629DcFJiyPXyLdQN/MtzBBAOQ9r7v6ummPGSV5xUT9sUDfln6etBXsTl
xgM9hdO6CLcCVyPAMpFlJ7DbZwz33zNpqBxLq1xqSwCqCJ9kQv2KdvIGBjENq6Ez5zUOvLDy1J5L
HrEXJHJvVEnBBo4lNTQCODcWeT2/dYNem+8kM7SuLzkx42BpfVgPU6uQ9oJK6ciUEyH2F3la337U
hghIJiOf1N7scoCiceYF1A0uv4DdeS2X/mROkSRdabCiS+K1ETtuAwXE/JSnq0Vfi8F2aLsHzTJu
/wouKXrwb22SOvMKq+ivcastnbHzW0LR7lgEbZ1aOst1NBBk7F9QFSo3dPS+tcTpMZqrfHRYlx5J
MROKpYMDCkiWaZ57qsUObIM4ksJUwPJH69biU8o9jMFg/qVV8PWF/ufLISbht714PlDT3rBcjjj0
zRCgDTLyKTw2zCJBkJ/5/noe8EsfNzhEQdik3OSwk3y2lmOaKsFVuwEB55mYFgM7lhcmxVD4i/qQ
VpMfaN9vcdFWT6rm6D15neSR+Wh4bDRRF1TN2lQRcgCZ9RvxwiPSm184mClkOaxRbLlvhKisiD1Z
jqNyKwPB0SC/XpUEhF2P1TAGKlCLihhtyLC0VQW/W4barKeu2+9a4axxUuMckjYhNLT+6GY/S9Li
wpby5evuXJ1eDu6bO+0mwGT2Dqz7BXnvkCVtKs9kDLjjsOJ1HQB4SFItfmekHkEILQ8BPQLdMd3S
CO9xvWExRDvpMzb5yi3gjE8V4yd/tddG8RDhI9VEe1dlsoZaoMu9BeIbboeS1YkKX/KRoOQMyyKh
D/q9XLn86Zy1kNIBhNCD2OFwzIZLtAWSnRBaFLMW6Dbto3+ZutZEg3GnGeMS/p4TQgEFyTcP6o7l
pQcjJqVUyopUfSPTO3HpeZ4ErQb4XUYtJD7vTd9Gqkx/Hcx0CBgwTafb5aAqKjgbXPua811Twp/4
tcD0VqO6CYcEH3Av6isCJAW2oJNzaX3tt339zUi7pGrjDItI5EpXINgbyWWYPXsYI4pRpQN8ZDnw
O5elyq1hg423Vce5f/OrJB6xgF86ssL+NyCQ0nZ7ou2bCVK6W9gXxFd+bKyq9NoHlC0bFNh2SVLk
kPYatajmZkkRkxBfeCR6wMhD446qXhf9YzG9QgVH2ZLMcIH2GuIgOOs69mFeYO2A7gb9xa1Hxc0n
MambN/0Q5mSYE+EpB6FhoUPAIfPgCZMfyadPMB24zEdI02GbB9iwGRhmX9mxz4QBIla0CNnFtGR4
u56layr8xX/a+5LW8Zvj56wWCDLAfF9S0z97iNiQE6W96p19HtX56jQeFwLtiF1nHv9/v/PAdeCJ
NaIPhX0dpeYvos35N313sBOQpBrmFPG4XxT4GLyZsJLUZtJedRWscJHuk98HyZqAyEVpV0xbP0/e
y4teXzUNNWiJ9Ei9gVX1q5aYJzf81izrMXfs8E2kUVsRf4MPkTZD5ZU/D1VGKRkCxthWzAhgAFrw
dG5l46ybgcRZk3h1QXAKL4douwwlX+oVeEftjnQq4t2pMpnSbbIFgTGHyIA3ZwpPtHf2xH0XywyI
vL7IMCQ7DKYfEBWKXgtayzkqjx06cxMDwA1VwodUOiTgTiCMKYQ1bkRzZSWA4iRtwrdBFHwyC37W
C9W8AQkBIpfPi8INYBzFXOZJnpF6OawTPt3TouOKq65XmNOD/lpq45kch0kfz0jVsy3LRxf+jzdA
78F3Soi0rGWu2C6+v5AXPwWvG+GaG+fJCGYQ5KqLNeYO+Q5k3z6LzgSKJYUh66a2egawwTjiYncY
gYuqwRxOTHBdgA1jE3eJZT9+t83T2aS35kdPGK77pfh0I5X4qY0RXIgNJy80Tb1PxBmpCm3fSXDr
Lhdtx9JXT+hE6B4yJJ79tCWrai1gIe2Q/SIfbK83ZGlIpyz/zWBX7fBPF4YzqCLQ3u9bJN/LwSx0
GCyAI/GpxfKeP4/8WgXSIV/RjE+a7y5hMrOq2jxU1kMRyXjl+6tIYfLYm4YffsO+6e2FL8G0Hy8e
76efa890ZDf8vglerkPgkK5dbn7clZe9jYv7TusbfuOBQcQWT+5n9XzI+6lrToPUWSkaZea80nzw
XLpC2zPY9QX2X3liV/0kRZ9/T9HMYmD6d7NtWSVRHK1FeC2zDo68LGSZkQzNb3vUX/A6qIVdKHcg
ySFLBT4c/TGP4bfr7E4OFeOiWg94pVevzfH390YMisenXE07iBqBqogv0ZCV4PhyevO/b67IO9vS
nxWX7rJdWDaPbp5uWpw0bU+7HUKgSYy50zmz1Y8fkMmH14uX+L0rnoEnk7iQZuapf859+6rm3NZg
u8WO1Sl93jaiIovd33G+YbAMsbCfk0vILeCILbZ2vW73UQ/QbPpw+bfzFlIJY8VR1Jc7+VAQ2ueL
uKwKgo9FOi3sOadHae7X37BrEuST4QCoYN5p7rWOnLz+phNwRjonB/p6ctbT0eWUgwJ75gg5QZVS
CS6QQBlpASKDslMXgs3naZezYDNqfMiCIrpCtZN1cALLt7RgVjtNz40P4tZx8cgOzi3sjjqWK2jM
Q1lnrPlCN1zB51bD83MZb4IdCS3XGfsgKsCnphLlPFh+bhJNHQ8aIVWjFke0lCqQEzedn7ODcQ8x
p8yL9pZZ7rNM8J3ZEZgUAjSDkGQ+3Aj7ZWJ8//ALEzzuDCuPruq6Rt6qO9ewOXixc8+zz9kHCfo0
ytUdMqW928aBOlLfkQvpAzakR7uDJLWgFRmNkIO+o64lv9j3hFsHk0K3ZMvWivpc5ot9JPS0RtqE
IplbdeOZyqC+TuAP4EU5KEvmEAybYjtRvuUjCk8KkQCoQWrACTYED24mahQOylxFHVtcX9nQ7ySD
M6m345ajJ8i5mdGfJ6i9arr2yFDORrOwZksPP2RMv+oPbGrbHa1WO19kIpeuSLXlzTwSkQwJKLl8
nye+Tzmmc/IzMlxRzfDU2itd2wUmHoQzy4VU+lbGAfnDLrfcrleux4RJf/ItNRyRuB2J8J3Aa5Yh
rdLjivTAeOlLWOu42dqcHrIMx3aKYtnQJbdDNg4TFMYeFqD4NZkrU+Z5DuCuFHlSY9/+oZZxlv8T
KZzR7dXxb7C47NJuOnkoeblh2i8VTOvguIdgrJ/2QXKaKB4tezB9o1UQp31Do8aOqLDKwTrbDRVR
kKib8d+dhHOaii7k6TNaHnB0Jyl1IyxrDgrYAGjZ6vyxX62S6AEFqJZ/V4aUWZhxFpq8vfIXeG1H
o/C3b2W9O/wtcT4BcPsoTZMC86aVfd/gb467splrO+Kywrv7kWFCg73qI/x2YfErOEQudj+xcoF0
Ru1uREW/sUsrv7vrRiZjmuomDvhS8EOTuMiFrd4KtqX7iJC9JEKrezqSl8czqkSyvM+jIuW2k78F
Nmq7BHHz4cT3i2f/uIJ79fAszUxSzi5r3qXPF4EfBrAHgShLRk+VxpPnLBbNsXAt9BeMvUY+YdgU
nSclRSD/qDh5YSRNl6jJjfBAe96WVi6AhfbWP9IpyqZcLTFK+a/Hfdy5TsZ4VkxIa83dTvcSnbye
EGkIFzihPE1NTdpK2oQCMOnsV0dfxzWvrEQWKTWubSzszwfwQNDVq1e+VyhR8tdiYl7xYY1uPCW5
f8Kw7nY5s3Es1pOF0aHqYJWo7BlrFIsBEL0du1iDW5l5eLuqgPHTE9IxpXWMDeYZFJGiEerjoYVi
PNQYcd3JC7TiR6mOivTPzT3LH45Y1kb6rMYNcXq8vLXMX0QkyAgPovl2RhROmg0VSj5bJbiPELtn
215R0z0rrrQoLELG96jZZe1m13qPu+pd4y9NDDQDzPZiHfkNuOClxgjcVbe1xfKAWbPDb0Oo+ZcC
xsF7WpDBpp4X4VX1bzu2GBYdBkP8+BjvXYCZvrMtaTVKhjsBTEh96iF/ijk34GZdIxuPE5G/zxA+
9nf9zukkaw42hQdxOz3W60pFt3auvMPyDM5mAsBaO2CBCZdRHAKLCFyLD28pg5y/NuS+Jx4DJvRj
V89aV8A1bb7lg2NJGNiyhGaoQFG3d3OxScg1n7Uz336Tt0lhSzWPE2pOlSAgWWfh4hdbCp18yhIV
vjiKIgHFPPlP53ywbGDM46aSqdcl0vlYkEI7tSyAsPWKKZG1H9blgBXvwngucGWF1+go1XW1ySIn
a4fyDG40pueLq7kDJFx96TevmsuZdI712cNYplD5UFSE/E9uDxUOKmnFcoCLm3bjXMPC63GO+Vpj
A0MTnj0qADkuMNy6pSrOFqi+ZHzn5z5fiKeWCiwtzzKKW2S4nXt7PbBPr46EIjgyblpQtkWrxN45
mDjbAEN3Yk6nfpBZTDAfjy+/RZ95yX3QLjoLOSscQ8J2LmtJFzRLBPTNUlulL2bgSSe4X17l/Y1T
MClniiNL+OulPi5AZFPMyftmTE5Fq+wPDQhMSQyuMhNlsQh8k/gy12m03u068snAUcYT+1XEHGnU
zyelFoIRVj2Iqs9eJ5ps/Ixz+16QguX5Kt7uA1DG+gnCzLmVvJPqcwJYWyzg2c+ORzmB8+TtuI2U
Dy5c8CFuj+CdbOgo4Xcs7AdzZ8bL4x3fu1BhkI0j8OfseYVNPyO97Nver9vXH4eAmiG5+lCdb4ek
EaXHXYzDziaptAO5YRB/IJYf2vQfTyY/RUPB3vhE/HmRLlcqMK3PbX72AtPutKWJ6mwTyMABpv8O
415OQpglVYlkwBW6L3vjuF+XXBOjvyx+TUDrulGe076IxobRhhyaD5JMVXPY7Bb9P475mN5vggjg
H5wVaXNE+TymzXp0wY0moeRHjb9uDtFNFE9DowA/FzpOMk+2WgMMP5UMSZMrFkQGWXgjH8AobRDT
2ukQaia2mzk4HCos7BsHPrR1pQSon705Nh+rbtcjJARz8qdLSIXJc8IoxqfX8GHMOvL0jL8VEdVh
v6MztufiSR4/dlImPh+w1klbwEKrtzKzMtwp809A/YhfKRQwxfyP3SSfklqV3eGlcKr+jJhJWj3i
QaWwfQqLhMpUM3gWkomCKEB305lQKdcm7OwRsjrAZZK1zoV9xRCCux53DAl9VB/ZrzIepuYB3Eub
7P6VjmznO8vFGxBDgQ1I6JRTh/IBi6ml8ntl5wWqXUZ2DDnEbCvztS6LQ6Qs0A/SPYE+SItVNHQ3
uEzQa4f0sN3+mtuQ/uO7IA3nGS5aIkwq6ylbGYSgLwdiehbumiim+DNnAXQjUznSGhjOI6QEQscr
IPASw45LHryK30oc4vykobAKneD/pbW0gMCffOwapVkT7X/iegdxlYOhGDEGJZ0BVgiyks1an/yV
m2AFkHjfzSOTRiOGpV7fxYQneaAEijkCfxi1+d25CYYLSkmqVYI2HMVgIEtbrl8dmv1Gw5M4B+Q9
NMK9IQrG4YkUNqKHpMvxxUZKCeYxKlzypH58WcYk1YzJG69LZF3QBaCAR4/TTXjK/dkZWPqSd9t8
IkQidFpRcYNtDq1y/LrVg7txOqk3NMmggA+qtkwgPp4QFe2P0L/hdlg9pXfIsrhv4OAPiDaqCFdA
igkYoTb4GYIl/K7hygT4keQ7Exu/R9vmy4dpwTVaOkr4vzmc6bJADv3tBtuwp53lHEbImgcY1B11
XsI8hfLl3tSI9/fX71w3jGLtLaWWBRqydGbknys2mgP6Y689hz2mLhWj/cy+ZNYwLsLVl8J4+GXj
SD3iDyO+SJxDMCoyzu8Rb7ch3SZlcHpPvAEfYvKWcsiZKq1ypgGGW+i7cwZfCfXPBcyndjoMRyqH
Wpy5yaWwtRLR+l/HVrhjp7SQawDaz/dMLyAfqlYCueXjReN2XzHWatFt6CeKRlLp7iZuKlDbGzsO
cul/8GglIXnOmmfw5rml0HVgJWmqTmr6nIFNXcJ4s/iRoks8OFtLhT3NKRMz94YvklsBoBXbQYbm
qpmd+4E+2yIZ5HXPV+VUJtJu/T8qND56zYlQuCF60bokFICMPp9/z7TNCxP+KY8bi303IqCOfA1L
CTdsqmN4CNtlqcB2KwdeGBrrNaPfdpos9UaXjAN03hAIKmRCp01KCWVDaixOW/7oVQvWn+hCnIui
wkJWiaADclHnjQEDmF01NQ0UAQdL3BUrPNMhdMFUPN7DBGdsnMe/f0G54el2EWVhDa9jCJG+KN6i
6D8EZUMOFO/ZPz5HfntyqR6ZWVeON7tFjKp/cWkBNBsu4cAL0oBIbRgj8kEwwM3BJfRygnFflPsa
SjjxG7gPMpQ9iMEUpj/nRc4KFfS0q61k3uuAXHeSj04pymorEYWO8TqPpXFTlUKFGgHBoj5mucou
RCh/uhOH0MkhGWf+G1/0BcU4QOlKx19m96+mFxTYiX7cG53iBczxCS3fmnD5N4YzTE/CJ+nYUL5j
Q2+9h7RoWR19Bw1oeFiJmrT+w32r96x4Nytn3B+3Heke4HIwncNCh7bi8njGPhWqVKF+qMTCa7E7
sbr/IDBDgSWOTD/OqdSQ3Cf0tBASfxh4BOHoPHRojN/7Lvsy+J3/kBbLWxB75LRJ+e7Xri9gUtfv
xsjOgx/4YPAvkzz58S2uTVrk+4lNEaVL3dz78fQd7oyRbJXOB4seixKuCLwMZ8J0c2/b8iNkRw3F
ePmwtUA36hIxGI+eM0AWU0RXeNY9eAKs2/Dz5akTj0fkNSS1CCbtzsaTpCWOG7G1rtD+jin6rUaq
BxN+3I2rN6ISoo/SL4/GqN8zIU69dUxtzCnjVL++Cw9siG1pfkJHgbiKqBqTMHH+Qze+X49lygcq
G+059QoAjnfy0s/WDT6WQUsgpxVQZW8ZqptXmYVU3gFFM1oR1eP5ssJUBLKmbiYh+8xTLHyYQ6Ud
Q9JQPV6wNBnBNokz6MvYIF56VIbA+bQE0DVj+/qBi18xLMj4fKs6NM68LxmyE/0ayfwnK35XjcbC
RYpy+kkQDMIrc39q9R0KNmmTrtnmllkf5Q4lr+TRRqB5e3sGUzbq9+tZJpmBAiVwutyZF0cTeeRO
iSbzEx/NMy0fUhV/DWNBLR342pPMF8FjRD0n9gTdvojZVQOfvaIWNYJiUeC8JZwQ1qIp7l3U9W4K
FONP0lQvQU1v+FIB1zmK2+1UusiBBJNU7lsnL0lA4eSkHYTq9Gs6KNwvslk+XS0M1J7NO4SSnjhC
W2mDIaKVmh1shumcU0qvglW4lAh/9POO2yaBzfOUGDLh9XFNKHlEMX8kjqoLaWKvKpsHw++0Bv6e
7GvToV3n1vCfk74MEtiZ6cfAsDlzIOCxhWxvRnsspk2UXvPt+7JmpAcSmRBVfWusZcRMoGGBnOow
YKBmgxMvsRMsCb8amUgwpis8PNt/CagD/N7vcZuxCGpYCLraq23t9PGXGJ+/UNfMRFI+xaWmCIFl
XpxJiVK8rKzVIkjNoQWXAbnrbjYoGVRuf4G5phYdnRHUZo/4CRkFuqUSE3kwToAeOiC5DhPwIo6I
KSgR3KUmmkw05dIAo5rSoQoMCxu7QLUApOmokqpV1lOd5WzcNSYPoL/n4kUNqwi0R9DRXnjl6aMT
yWpcyGnZC4cPOjrdil0X+bszk6W5OwIfaaANpr15rOpdaUVriBCTLOFRJT+zbIUxawqbb0jdWNuA
nPaVSDip5ROMWHZ5udsm3XMddRTvrGbMpXCyizY2YH3Fb3hlmrb1D3QLGf7FSXyeUof3wNZHO+eH
BjfnY5NnC/eqFFJJ7QNoHgXiCuuOTXwr81OSTWbcaWntZJJLq0JCWWlPAJ5UuXBeTXc0wONvpXcg
1T+8ZMPGkCDsk6pkPeNkD/M0QW/y1+yHXjMdyjCS599PXsQi3PMlLgw0p/P5yeFeeK3OfoSePxdn
jXAPZ7tobovPOM0tOMWkG2UqP5TutEBbGozB4dV8wb1J94rfVpOYkcKmwZQ4G4o6UThyupXv5Rqp
vMP+TYxy8mtU+jJC8Udl9a5gJDte5Kodc8sobpmrPPU1Zwz97+w/SEWLtQzVymDctZ0U2C3ZCdRL
B6La6Maydq+C1SJB0aAaahTbkPq5vKhcU0H+PZRA67IGg7ujaVrilflvWYhE9F6EiTTzDqO07Oau
V6fgEf5g5iU3ESeNyh5u2bnCKLdl1XNp6F/lHqIWCsLjI4M2yQxDpeKhFEwoaAdKxO+zL44u35Eh
I0V6w9QyLYM3ZTQVY+TbPeak41SgY2N5GuUqEXoi5Uf0QOEvG8OYl+BugV/+nt+EgQntbtEFym/V
J0Jc+1MQstoIyJ2AcYAXQWZKma5lQhAz6biiIbXzDRF/XDZG+dKjzuweYZuzV0x628A21Kn09Gm+
0coFfyplth6ONJU+FChKlGtbL2LjH6aIH1tDMG+mgrlV+Gx1AuEc/gFFh4bbHbiluiWHO1BlKNjN
e7UE75T/mZzJDCNJ6GH8S2ZxvpSYVmQL7eVGy2K14FT2xfUSW4h46IicwetB9QJEr3qOaGMFe8BY
+VzoyuPLXW5M5/sNkbWsxuDHPXDLxxUKy/w2llpucb6mK4jCI9XHDUbd6EJZhEfPYAcmnWqJPmXB
dkNVbfqWbyLIPk8VS4CMQJLr9o/yP3a0K8lpYkd0PQm91kX5gfn0L7gW6mbrwrWsdYaisTpqKHRM
Bvx0/joR0CnfuL3qnDODEs6r9QMUndZa8I06L191brZw3XDK+cY+VeCh9IyybYOSpG7dvmyBF/ro
YCisgy/b0le1YPlDihyANzUAA+4uXpAO8pVlkNpiZfmyi4P6kMc1plNoF6StOSPwvlGSME804HAK
GHHubpu7ybTvyIgnUWM1w57j3+qUjI+n12p+GKrWJIovofMlufVf0R/OFe825gd4SOqCJu0hyNl8
s/cUcztVDJ4DH5caJ46GOJnYanoJDdWeK35RJ2nFkSFzs3NzUaqctcCvS2OXF+RkoQu/YiVMBXbv
ZJDevLmqtti3Kgf1WtN83ICXgGyvb2n/jhVMdM2ItNcROBTtQ+9mQtKjdWyY7DgQYs4f2gNXcst3
VIe4DEd9pWPxtSARkq6PYjkaHexzVIMI0kEICOyTS40Lhuibku4pb+QZ5Md9y0+0UJLcpchBiXTX
0TnLCmY97W4hA7HMdIVsK0u3AVdr95rpxYwoKq/d+SxOu+UW22G0mBj0PiYwCmGTRCCrAMxXe4lf
p5rh5VcYCIkBCG2tUlMiM9juKaSln07hD7DVr+K2O9/wNyZHb5EpuOlDPF4QOZdwsCT24CMdIqgW
z1Ww+owMLI0yCTAnEKCTKd/t38GNQoSziroDOTNbmPo8GndpAV/3kK3AB4phYDrfh2V7gymfBR+H
9G6kKiNd1GG5HvR9QWdE+VGB3cSyH5+NgunR10XBuhlBSG69W1QaEPd2z3bumthgSlcufgY9fKgS
CVZhVXdvTnSy+31o1gaFXgcKviv3f+z+lRO2G7P8Jhj35lMFVZ/le/lV0e9OWALL93VLyfGnNoOZ
F/4/ADPSWf/5UHXU1UMAnjCb++sppnIQ0Mx5+n8jRXtsiY17dnNP5GY7jFY/7zhQXJ06xGW77lPU
5R4NJ49mayJZ3X3uPsKrg+AMoLuk4kQKqWo6Xfm87SUnNhF3gIIA5iYUdwSlc66YGGCDR3aE5QZt
hgEtJrGynZ0FlK4OqFq/2+oTqiB1bJIkPTWXdZ9l057lvquoLtm3iAJD8hd0n6EfWrb67EmzPos1
L8GVhaX34KiGosYjXYVCEMs1jlu+g0MC4UHO99wMnx9oUclZV14+BUPDBJ6Hchhr/AL9SyE41tv2
sg61RrN4ON3Nwl4Uz1/KYuRXOLEGyNs4bvP/XhAYZihJ7RBt2FB/ZC9BCrtrSJg/APXEenOmW0NV
qeMTEXrYzTxkORTDB58PO56+PEStSqq6afqZKfDbW6Uy8L5OlepaPIgQ6IGbEuANUnJ4VTF1TopO
sZTBSNRsDuZef1jK2sjLnayf4Gmj2Y9dGOGp3sy+/X0Fvfx3IBfagXtTslKfKWPrzmy6zVtW7YS1
BAWHNUvCQWCyUvQuAvbcMjasEqBr6oC3Mq4A9OaOCi9rE59qlQ6kUiH10WvR8Yk3UmkAKLPSGtJg
QNEx4SJLzjwe5F9R+Hnf+WWQuD9QE/WyvsU+YRJ1lR+NKDfdR6mPB7xj1d6YR9butyIAttHG4A5H
qLci9QXDerFbgQaR4LH+DpOPMu7HGjOq6GRHwv86vADBqkAKoY9Ci9XbY80Uj5/BAdBlhm16fyrw
Kq75gPRSJIY4c9J8HyeW2WJD05Z9H4b8T6Af5+98s9zMBRGtFfxtqPUriqEHJN/q65q5kx4rvY2z
7RxY/Dxuo6tcXzsihoAV+gDuCGeeL0Q0Qu1bG8nXmKiMY406D0dVHnALfqpZ63pIZdnQ43/NHsU4
gaueW2hiYBYmhiEdzRs9ePdvLv3H8JSqlwpzAF8hAhF8h1T+HU7CVb2Nj/qHLsOYIVgfLSMeR1yZ
MnjwWDcK/xYpCzovK1oBkVf+XFrqKcqci+EjoEqB4RmDcn5tNMGiN85F4ayZ+TDDEZIKnomM2kec
S088QQLabQAhHrut4osE1R5WfsDcL2benIBmNOLHqYSkhbgCdlv3RXPRE2unOkF15a6uEHi+eArN
cQ7sRv6PBYK7D/Kp9k0pfVolEygpRDYzeGjSMZGdm0U7EepLENVTBmCsJy6cHt+ZxFED8YIoAEAD
rbiFPy26Ij6xkTCDtPmIT9wdLx2USA+Xa61Ru2XI1EriOCLgs4q5kOpMJjm2398KlFw5WintFt+1
eK1JRd4GlR0x0tWRvCOA5Gliu6VS0YEBuiZW3CBME/+xnGuuWGLP3TIvaLWPzHMiPaTXiE15nv90
xvEly694bAPBQhN2POybtg/OV/TjrcdpjlTjoQzcVpQIs8bZKLp3dzgyUunFvXaqn0LneKAE2h7w
+mlrwaB7e/W82OvdiUD72my3NkbmQ39380e8c9TCLMx9PeskrbIYGwCpFPW71XNqcB9nWpjFvV0O
0tabKQLLuKF6qYJbtP84mO3XOKj+G8w4Xy951notjrcX2FL1gVBteiX3uYdjCYXjUruRxOecpX6Q
d9UadtnapXMRXeaSNTZhgDgXh8k9SfAoAqoz0la0OPemehnQjT48T9d0CVGrEU01dKh6BsSATmhs
0AD+JYq3jnIJ8Wv8zgb5jtWbgO0zwvpfqEnPyCDWEjxO4Op3JTYKl7JM2QfaupGLgmwWj3HFYEwo
j8tAS1//YUxG8jtoBzxe10AxYnXS6ZYohuqoB9XD+PoT5lGNyt39V282lICawp01sbDaOeG2EKOT
X9AVxBhMn4kekoSn8WA640NFdnpXsSWSqN4kaqzN2lbbI+EA76wbmfCPhC+gZrEnPWG0Gs4L28DJ
Gy8cdQO712Fwq9ZpdVuiBstltTj1XR6vp+QmOA0JGi/FIwns5oJUkIG3tDqNLypUZ5OnD/W8CkZ3
91E+r7oVH7jaNp6u4sSYAidVtC+pg4AMFYrE5oI7plSXjsfeCPuGdHY4exnl7s5wgstfSXCow4Ue
aogACofS/SLpaOUtdS6XR3psrls8c9kgJggsDOuiwzki8hhuE7qmNClzRhLU+wcCP08xVhIUHhZt
aHpCWonekCZ/+uXVjoXHkT/MQXO6tG1brfrp6ry1AmOXQBdANiFqR37N8exzCaV/YWTqXyhmJcGR
p45PHuI8NrNG0nJOOURZX6tbCwWACfueUBp5AlRnh743QVLPTdfvKwBZEBnL7Ty0IP0pJV2wGKKf
/gxAKKFnsPeoC8icDOXtgaS6pMTRn1IZdC09VpnSDFTol45HlRdkmgRu4x+q6Jw5D+lU3V7B0lFc
BeWNKaTZHXsUUcVDWQrEaaJsayMI2JwC8v0ogTTfwxa3uNRyu0lZFAYUiNNDpr9oRMSOp94hswBp
bZHPoAGCgm2zSUmL2anoNx4+WZVD2JjdJWaAlJSQ6PFxRO/EBcFH8mLSszWzDk+OxmmyhXaQCB99
uAK7wSzzL/aHxpUwk1PPg5rh5qAnEN7MYxH/zNkzByvHULBNMNKypDglg0ORnIWwG50GP/v0QQAy
pKLlFKSU8RHA4HbHGvW6WcdT/SvVuoxreaDa0oGv5yIWHrsk+r1KxiQCI3NoAc8thH3aTlO2tJfA
ePGsZaYhJ/eJYflkz1hAIdqhUMrPkjfZzYoligvew3wDgMueHuh13rUrYf1s206NltXcB1YKS1I6
HYhui/IeRQ+8hETZlaw4S/VX4GymkGqu1JI8L2MFbMGi1cbJKWsZdl7sHKLnNxvPLyJZAf1xmSjW
VXaUCLr/gDnRYItx5s1dvkyOg6p5G9K1yTkysnwF0X0CdDBuiXx2cWWTfeosQTO+FU0pzjd4+ujD
XKDpdWNZqhLt1XbScENeLB5gXJueLPArhlGYhhw8bm0a4/dC0fUT8vSOldYM5lkrv38aLugjKEoX
C7qdTJtfOG/toRr+SOpIupNluQEvTbUK/CO6fyd8IVggHz6uOVX+9cxA8k1v5iKYheTc0AlYztFd
tLqFaIrzZfquELFmeQGryaO/SoxnL2qHDFS0iVTTN2f1ytPghUrIHhBSkrcc0h5B2r7HGUmKyBv5
YCmzP2sS5JNqGdHQ6KEtkzeJvbdtVOliJu2mC7JWTUTkZb0oMo0I1vOtlm+86Rk50GNtfcJCBwgX
iq0uGxuZoLzO8cjbv0uXz8wTQkoiG5pxKG1fTdh/KEO2CzAJHFDRyclmGnrzyQX9Dngn7qFe6N+D
Xc7aZM4qKZ8AqKe+JeK0VMH40yYseRJKZaOYk9UybueaLxMweBlxBtXNOusJ8UyKTYq0cuKbgqrj
ZU/Ygl6ctiRfeSJHNda1/znvZyObyuzU4czvGs6mpYAhydjmqCd8ks3ABKIqjO3GA1O09tdONiLW
p4t14CwvQSWxTa+M2EhyRJlgDDb45MabdMwNhryXfbY2Hz1jDxKyoKER2lC7KzxvpgaatUIw9V4f
70HF2l9Len1r7livVoZH92D5NsdeE/5ujBX/i43NCo9KEUVMwvjKU1fFdcKnyynFX81p42e8BWMx
NrhqxdnvhkEN3c72aKXGNwNJUD+FAGTkmW1XetgeOd7cC2z6puJ3ixdtptdRYovdgHJ1lMqSASiy
D63uLeUa/nG/xBMLWOUcworALqO4sYOqBrKOxGhDaeSxgK43O08YUTgLrFWmduxE+DyfI+ciZrfc
4aBLJ2P2XFOqRHyJBIueBYzLHCeG9E1mgnCGtidLcimkpnSW6RdHfsW+oE4dvlRpwUsM3EhJHQn2
Elpc4A4XduHj4notWkjfRUBS5FczdTZ5pcJ5+oyRChxtgKrTK4yRXKy+WqnQnv9fIEVKCF0dNDlp
2eV+TPHJiDljXFegq+hcq/ZtwyaIJ5mbJOa/ZmjWC85CTOUKGE9FE14eA6r6S/CwJ8Tqb2q/yM3T
w+s1p6cCg+mSy9UT6z/ROJX0Zb+Cez36rhDqgH9M9OjVBB5KgKnbE9TAGB5qoZJXMkkjXwlQXSmw
aa2rztytEoiGBU0I2f3TetKTpuUDF+gEJShB2lIr2GSIt3T73AZURmmytKCb/2hXYC49xOz0Oleu
DM+aH1gFg2//QL5HxKd8x2TTbYeUEGMObx9UGSHvUSc35H6IN8RJHjirIG6K8JTANC1dvLO70FCd
Biz9I6Lu1Nqqf8hgUOviRkpTaJcyRXG/+B0bqIEpjJxeSiiYsy5YrwodDYlBSOMjdken1nuXsXHM
KCdgqJxv6jJQPFNHslye7OFhZbNU9qsnS5ESKqj+C+hYRHyvT/Bth1WM5FP8FyI5TSt4jxwcDfKh
Ul/JsV/nqwoPst3OSeO7i/6ivGtaX1zpywGnVeflBst0oQfCmngZ4xXJk96lynOYxmID0pRmmv5Y
+ZI3jhnBwlSkFjPrR/vNn38su/0q2L8BnB9ih3/jz94y39q6qdbds9cgXIy0X2RHhqpLQROVyHdC
n+pFt20NVpqumahW3px/p4fsWyrG8a8fkGxteNQcOu99D/v42NtTd0TfwwD9GFkJ8WbDh6bb6r6c
Qe9AEvZ7L+cuda8cY42Y1Oga5Bjil1xJ5+mp6atpZqWt7O4504DM+jOtV21/IeoVmKVYml5jvmqx
I55aGb6gUdmkQm/lMAVSYAmQl5Bcfxn5uxalqlekc537DWEkMo4TiobPEQ0rLu7YZyiVEbVZ/bVo
yRef1pze38SUgpeN+t1EvU6qpRWl/3kKyerbIKqh72l+2YUT8UpJX/yh8xAIVw6sE7DgvgFA0EYg
Q45IENNycUTuWfoR9RHj+i8lUEt/3Zktx9BWJtKIG/3cZEBHpOLZRDe5b0Y7k8xcrZIN8ZKtS83x
KgbHO2kwRahyU/0F5xtEdNrQdhfzk92Q4lAwbBTx0cMbAK7b0GJshVoZryc2Pukq5p5hQA0b/Jeo
bJLNAgNvX7VNhzq5OKhuejgXr48yq72UOwFjqWbj7ojQSchvUBnQjj8buXaW3bmL+W/++MB7y8tL
xebPpb6FC6IpGMs23YD3DTKCSUjlOdHYOaIAPg1rxKtoO8TBVq+Ea5sfNQb2pQLL+BIc0N5vE9c0
/8SGH+w6jNvF1tJR+2k3MAHowH+MQxMeFRnx0NgSe6CXU41NozRO/bSGb3Q1iP1Mre8j1BBCmhvI
pTfCQBWK4xgjfLheCXgcrkhGSgHIomMeeggilQ7IqS8LSfSi5ayfwE5UY+eck1Rh7/ZPzVyZXD5w
n3KxlTRVBULN0jpqHPPw8x+CwsdHXJOPxvSpxtlnuBMfN69vm7en8U+wAJ0yDzeLle5QJz9pQGzN
boww0j45H14nubDI5s+Q8B6EIerGijba8dhNRVsor9YlQkvoU1rE+flxe2OF1GBs5qpDBoord4Dg
L/w/Gvtho8OmxWzXozvaM6OCMH4BZ+IK/0+FMDRl3wp7qs+BiKRZtSWcPTCQj2zocAPrrGTpScfo
APnKpd7rWkTCJD4wWBa6R6fSv+iBuPbP6v0cOClUPPEhkHPrPMR4jF4GIXzLOKgoRTyA/ExDqy52
12xXWZdx0ZTOlUSQjWzkLHhC8clxpugBSapjRbzkGItjWlGgjAnXSIUcDXTe6BM9H1qd/mHR6/fM
CvD5cjwQovtqcYoKFVQw5msmvq4zttB8uJ0hp8iPUAblcck/zpxJ2b26B5El6J/xFyMz95zUS4rk
mJ8uXBgk0JwDSsQOJscY41n9okEUW/TiuVj6rad6Y0sNmOxnAnX/GTUv/vdg12ipiSNCZ5yLNM8B
dXhFyrHlhvJsHKkCs41Zntqdqc0Q+to7rRweYjV5D+BiSR0JBWKqpYY0RnvppzLVNgrg/DVsL6kP
WZvpNJ7OeOw6D5plQ/u6OouoSL9VscZYTyyP70zY5UzUnkIUvKEfBv3d1ohTzyinDVehI0Jfesyh
jqQeV8gqVp2PKzd6eUF449CqSaD92WwdrL/dAo+HNfstdSYbSAG8mUu7YJ0a9jMqoNd5hlpdiHLM
ZE48tMk/RoaWyY7r79zeD3/WoF0lzTYFXjIbwKYcd/gaYWumn/DOCizwMykyirrAnzptEm3WDWWw
t3pkmRONwjcY1ubgYGMh9S9OLdYObYGg82azd80eTwtihhM8W/btE1+JwWbuIXUJgtMjrfQVFOjw
VStpSR5rriKluCnn/+IcE2XXVX8cSHVQD2Gj1Rj3+ncMqyWis32+LAXvukwhofeyhSXJ/0ci4hTs
LyjZBUn4MJ4jZ+Lo4aMEalVc3dO5I7YmuTm47KuJ2sSM1Fxc1gBaWja5NJKiznQhcnB6mpaqySME
TgMH/VDLotjH7HcU0MFzdwdrY5coMRfJFSsClEcN2m3lAFpIYbT1NzmVq7B+II5Hs02mVIQE2O36
jYsg63kAh2MGurR71C2CBMusan+jFNuSTJ740fN4ok+4dBAVOQoyya08LBolN65umyAPEe+qwE+f
CUR7yxaJ18vfkvRIw9XfX5LthOi0PePJFr8Hmus2KURejTn1E7Q+UU2gN3sE6J5rKrtywsNoZiNH
sr5ZRTl3GhOvjTt4czH/+j6f2kIBn/08Cb9greqU8vSXSbVuM3kV2uLNhh9u2btSnA90LL3RIYQv
FsuzjDUH0mr12/CnUE/KSc/15x+td+DLAQrBDDhTUdVeWCDcqVUR+8mTjm7fkrDpu/fThb0LCQyH
MBGhyOfqwT+iNFp7JMl6zzCXZfYw7gUUwyNW04QMjEb8TsSnJo/oC0nVpw1PhzE5U+KnknCmGN5Q
+FZ7OiabzA6ebE3Tq2WCFt3N+YSORxzKP5ruXUgPWG3fvUnBfdXcqQCFbYy4XeJZhQJVdM9CY76l
7KICiNx0DoCGua6nUaBduwWGSmG54aRPOv06Pw28/jtigVbzetrJePKMKJpVFzTTaqIb4efZgmZW
3HDJPBEv+2Yunp+5heWQb7LGw3HI+/FKIiKSOnCqLGmtneEWEYA6Qcw3bTU8hZS6BSJrPm5n2gVr
0khAOOrKmkhR2F1XAQfXOVCfi5W9sUMQJcJ9jPbZfQ9TC0SqApaoyMIgeiQHMHzMcRHnk1xNUYxb
MlAPcY2EhafBQt2+3zHSiQjrTSzx5nGRqOiCARCpFvybJZOc0/celndepAox9kCkI8BAyzuazGxT
onOtIYlY1Glp8f8bDAlHTPEQUhKDlW5K86hUvfILc03Fvo+GvyfAUqViP5GQWyAbOSmcavtgvhd4
WJakfgALdr6XmBx7/H4S4LbU21EXENqpdChXFjcYZHujTtrEv7jPr3dP7BnsmS4rgZXeJyjQYigX
2bZE7/gkopd0o9Vs/EC0d2FMGETb/52HADARLg11CJCXXZkgJBZUqruY1jIE8gQX/5uB8tJ1/05O
r7KIgyEInXfDDydfX8cVkjnn1XOUcxNPi2Y16Bm1qFN9fVOg+YMKPP2IzndmybdeYZ/xsmC1MkC0
gRzzx3mmTfJnPsxXdVZiYcH6ohvTxRem+FiiPtVUekQCeo/FaNS6d7tM7MV6lQLYtCJCo49NInWG
lN1C1RHSKLScnQCAOk6xjsuS45IwWVMUyj+DQ6z3CeqnimgUJrOLb355lh3st2oOp5IDDnaQtgEl
H7WyzDmtvzQkhQo2kMXfMSGlCr88plihKHX3X733Oqq+FASFwAnFU5BKSDRz7SgrsyZN3+4kM+II
GjnwICbtsx7+VQ1m//5g0LNXKM42Eufk8mYi4QsUbfvaJCr+xTvL/+oFV15D6pCE13s1LXOJIbuS
qeFEMKKY+gLwguN28RFLOsYjTBeSQeBySplxT1zDyETQhBJq6ruc1KIhFNmaF+fySERXorFTlII3
fuN28R8Qq211E2qZ4AWdpm66Kzi4j4R/pElWLKEud5+0DvqUTqG51qLZmIaOOavU3Xg0uTsg7ags
ItAg7c7KzxV/LfShe7uo5PQauqNvv3By4xGV3+QQtal3HWxhLcllmlBm9s8JYptrVrYIMzTwswO0
Iq5QChbNViQxtx/DzeIDty7nRFmcWWA7zSOeVf0Mh4hBUBw0at7bUdKpxe+FG2XkJG+fsCCZ4E85
8eTSVdMvyFz1CeIqw8fGdQ4nzag6BKFPKA6RvV6iocOa2WimI0ARCCvt8sdAwbS09+/H+Zg/AIc+
982WvoqUMV4qupQQ0Cc4VbMxdlnld6vMztV7lgIC4rS94geUOA94Ba4XcvkNGuNOU4S4QQwku9WC
mS4W2A0TbE9ohgumrF+emTagx/PzvfT/i00qBjmiRMG67BXG9wEQ3JbUDqJnDEJieohr/saIgOjc
Fghj3mbehzS+TvXqYa97oo0V1kjyJYXeAx1DOW08hX7xumAxt2op41U6qbI3iKx7PONNPp0b+JJH
6prtu06KFVno/OVkfc6ZhCAVY73WdfR5BKkeWk6kmDCgTOFNtzyGjaYi417OLeXrQjs6yh516xeL
I4vevvHxQzyHGJZqUZKV1Dr5MGkPJu5gLO5w+ORp3HIhLdN6ZKe/h2kn2cPXsugMqFiA7TCRO2SY
fytuqZ32JiuFovOTO3/+K1gGNjf1wtWffbMdkpDpL/mGSGZTUavNYXNsEzAdDtU0dei8UmNhEz/9
lPlbLDyzoZXS0QC/pwkNW8MEzmUNGbJI7s61oog1eXUOs6AKJ+NESPdIC6bGXV5DM+0b8DjYFTd5
jNY1usgqZWVn/kGQVdhzKpbRz7jl1FWQOyaWqw0jkjj4jtr0zOpAj6FCH1TuUbRlfRK8WPN6k+fq
uIjPgfolwoRkWalyTLYsHu1FGZ/76Mg42xG9yZ4L5rBxnZfFPQPPxc3TzCkG17ccTrIpKDPS3P4J
Sp3g9bTN3Rl/+Mw0ZqNLpJ/jSGTjCz5AVjOcfojM+uuoKcT7ssDM4fTpHLEJfpwVoOVVrqURP0QB
Dzz9kAoUEaK35eNjEyhuOsD47ri1FYPhCrX+rezQdAv2JjaHtcLsF23u/FnmLzT6lVBrP3xX+GQ2
Yxc8fsn77R/kn/1BUActZ5ZbjQez7qW7rW6Q84KMah7Szbd6KxVHkXjfuVr7hJyuYKTKLCvEGLp8
u4IvV1LBIJQVdvNXV7yXuZZDBmx8OriOPsIdRd9eAPgerU11qQjj71m3K40XZxNEtnokNwi0dnDG
+l7VSE02mGj4STD0UGQVrPE+nhLJCXNBszXO7nFumCcMnTva5XMJEmcChhVvdh2Ay3KMrSCdqGwr
6FWaUG9uBeV3YRT7AzeBPGisqPDss1rjZmRIlH9MSQxB9IX0x0qYaovNOrMTn0KVrj1GpHWhCkBA
p2OK2qLSBHyycQyocnapgdSkusMGhw7uI0dGj020Ee8YD7QfvNpxM645lXiUTZdSj/SoaHMUgOal
4aggmEi5MYYAnXhA5LQjfP2rp6fpFwzBkvX4NR6r6XzfhN+RV3tCKq1ClHh76p6jK/xMnZUg8SHI
HIzpQPzQfvUVZcxcp9Iub3SqW0b7+a3kpHmaqBP1AJe5SjSO+co6nTVY5C/dvK6tWf+bZNevR/so
JVGbkOPYyNOcDycvv7YriwCrYtE4G8P8vhetAiydTQ2T4cToUQykBa30txTUMT8H4pko8KfNwAgR
8zqU/+oLw9iR89C2vCo121b8eP2mmDM9b0SaASvIGktXHgIPsWObxV9pU8AhSy0kzli/jr89rIT/
/4llA5EHCqrfDlEINiHWoVGXXtuCGGzQIWEuI3z0kp/VfJXsAkzGHUbc+hm4iACv7FvZ1AeaJeRu
45mCa9XdHQdvEhqrJaWLJ/Om4kwRrOZv3kGXofBxYGZ2NHDqnQjLIMBVYyOB6Aoz1ehGAnlccoSP
rKbZSkLrRewFYxOrPLfbzLukzYIwz1u99lfOGs4nfiymH9u67nAoSdofo2w2XqEEAfwK9z4EXsi+
RR3QvnGGFCcbSYTGZEWb5EaGaaz9htBV1YbPBoTWJpj7qnJmlP1imG/6m2DGMHigBNrMQ6Sf0H/A
sT1oA8FIEO9wEk3sxeP4pyhpYPRQ0QL7MH7THM5RSJuCfi1q3fN7YsSjQUPvPrQNYBWbYgEgPjoh
9sP+Hfdt9YV4soDLoCOe1QirdfEQBPX9R9n+UiPkJQFNN5HBbwHT3YKen/YqRcfZJkTNIUsDkXGq
rWoPP+JkzNRwXqB81+f8GBaHzyRZjwQhX3/H0I7EJbBu9CDp/h4+byKomScQNCF0EMSJb5nM0yp/
1R+FpjNUq75JJ5vzi50qycPzIASaHcHgK7uNS/rRtbl606lNPUP2MDIpkywDfwVSa+RyMgb5BR/5
NBaac2nRG/3Kxj8NiIsbw+bBowEzENHIroL0fwfSay40gwB9SOCErvf0RTAkh/+os0vk6EtjqbYH
9giwqR6SkN9A4aIa+l0ThtmmkFpmWrLhYkOYYVdBx9D5su/m/J/i/fq9oJ4f0AiJkqtHN06EXklz
PxKAbhnq5+/0tSyc1QUiZV7NsFyQO7vL8vT2+F+DcdJJu3wY7LdKQ5P3uOff2KL1P1QZ5t9QtscI
o04Ikefk+p1E3//XglrZe0fyymk8CpJTZNtRWBqF/BZoYGiH/HMmXvuvCoMxFHVHKyaboYDH4wXs
BoC2gzRRlzkNvT2v6tMlXltWfc/NjViRq2zRZ7nSDOLcHFlO7tBQs9gjcyN3rS3l9hsLAYXqTERT
mT3+XaFM3CaQFlh0L3I255tZcvf/98h9fuJoDGV/xTs4dvErii7FecrzX/zUPDKXC1LW3vZxUIUq
Y7Z4Ep29SdaB8Si36AHIHNvQOvBi9FMHGyZLCtDMA750AK6rxL33i9+Rklsjl/j9dZ8EmMDZzUn9
PMsCc3PAoP+G0Tc8waCoX3vimObopAtO8Qp6DkNk6BU38UmbTROAJ4cS8uw7lnWx72+cZECTQLVg
MfrGGiKzJokmLRdGM/zmMM0/n3JvQqS4oayTRfy2V38NOjOsP/ya6Gk3Z4fMzrVjgnIIqjArwN1j
ljBPpe2IyZGxjNMql9DSAY5vahFrC/+5cz3VPQ8aAA6KjwXIw0r60FPuP4fODIysniRv96K6DFtw
KbQNpEqJEo4MQsD99Z5nrM7mgYOXzMoqS9PugD8SQ/IFxlwyW19f39RsiD1RZiYDDWy6psWAjZR3
LV8+Ps8SoWcDCQv1Ioc1Q5p8Uk8ZU+M/Y3Hrn921Fkuum9A0ylr5TNWG6QRmzbYjD+T0np3FOXZ5
5KIKekWZalMHaKy/YnpgNepQttBjMPMzyHQ8iwbQtWfgvXn3bjrPvT5a0lru2JvanOKubnP1w84R
z4A5zAtXBU5UROLgk7zyytD356N+sWCMJFRQtCBqe3Ga+wuS4aXkGHVy2jCF5kKqVCaQv2IBl8Rx
RTWykVMnFGnVBvJ0Do+3p5UnuipyPyC0CBEd6SIXvn1LPQhq3fcVjGtz6Giylbt6GnGGH6ClM6Ek
GoIRcISrcr9J2L2BLCgJpDRir8X52Ko67SbbosLfsD/rqaOVaRbOdTcPNYc6mS3n7uJ+eiFZ+Ip5
5gIIoUAWItfXws1xeBoCHk0IXGOGvlFVLi/zmEoH+UR2YrId8yMmQSXVVjxxHvZ4dxK9qmLW8BkJ
ioU2cOw1vaeBUmFGgY5gEiAlvsNEMUfQNVXe4rl3sRvP1m8yar8+H7NngvBEMYSO8KWNYEjULNun
pE/CfOfk3/YtkriwdjpaPa7iyKA0qeksXDgb7nT5+/BtOsSQESZZNb+r5xIPc34Qbh6hXZ6rrq+N
B9HvZIBQU7fhLdnVrSacR9itW6llbPBBSKoJFB5cOO1KDDde3S7FZZJZUPWiVJoXcqPC6OcOC4br
X6xxYq3CQNFrwOt2PHBSxuCI6PWH6hcTzsKcYTzDVQTg2vUgZlgtpwqqnb015jxe9Q0R6FQ4LQ+X
IOm4OHPvbP6IYtylb6OPphyilrvIDZ4Ic2SBta+93FdP36THDfKtRLvN6LTl1CdEds4DKUxPwhCA
Kg0ELAqn5Ca488xgqf7L2cUBUgHWRACmY7k8qtWEh1rxxo2MbFDnDuWsHS4TzrzCxbINLwyxDqBY
4DJQSBrNs8IGs6JYc8vEg/fQUQsqa2ML5scSphvSikRuv+ESr4ttIZWpjcdtiljNt4LGT3XLDiYZ
9nY33KjtKLeg8xeHOmCDR6Ue5yd6sLud0rdMawWxvcCFGU6skgdi4wPeK1gu3G8x6mp76tM1mhT+
xDuHIZZFmmVDRlHt7CM51UTORl7Sieruo3Gem7jyjyDBJfYRr9otmivx3g1lNjE4H3krX/xiNhbE
Xes+MI0kmPZQuHvP/YDwl5dLsGegwicdwpIQ6Dt4E6qoyCZviKUs3FFb5Y4CCQ+Nk7sKhH0DI9D+
Pp+/IkJXgtQDjXSHqbkAA9ZANR79EGl0ZM/wKjQ/ShFqpiFw5fyCBBK/NCs9NwlTuGmiIDf1DJ5v
CPrDcXgFNRlDG3Ci8FLx3mpngUeNecOvTFPWjeOd+1ZjsrQC1UC93OznUp/6QakqcrTLiFB+bWgu
COl2PwtK31oD0sIGnYsBnr8h/GZtxh6MIvknkZhuHLvSPJ97oi+/o5Fx+axZdgvG/LJNaY4E1kaD
x24e9bgZWDolGcaOaV5CPZRFrFJm/hy9IfBh+RzwFemkspLw4TYuxvL4zQ9XU1ioYccy27R/0q4u
0IBuF6fu+BoxWwgAIHlXXtielAyuh38duFRKULGzWaLeP9dDHM8jPpbx6/Fhl6dbwGVOF1trSBZu
qax3T1pe27Hk1AJ1YwjbkzjHzSS7Xpq6nl7iytQMDCENqZzkeLB+5xLfnkqPddCFQ4LZBYdTmDqh
lbLSHsceTjyYB6O7BCOhqeN19eBk7RVx3sKBT/Pk8GI+nJzlS8qDnLUlLfR0EruXKpX/MC8xGFAO
IMmcmvwF7kdDz73ibb2psGPbTPT0e7lJCgV3/pfkuCSsAC4+Atqu0yB3MUFPI3kMzYsbrnz9ua6t
djOBxDyNhD9psViIlkLCOfq3PFVwK+BImgFa0mPsvru37YteaFVKUV8Zlzm+eEdCA8fBajUrsg/8
D/2K0kpaA6oYFPgNzQ7Da9odOzcD111x4ELqshLkA6/LM5hUbPqKMNyKY9x4QPWxg7MI4UYibRrF
I77uUCg0+wYJcSL7jCgb3sAivzpuE1EDOJeaTjEE2UIbkTAHlBTc/rikGJceB0Px+Rcd76tgrlo7
4wt8eJlQbIBP9tEguURLCEx5fo+Z6BF2/R8Ro8g8EJcGzlt11UdpLrPiiCKgKuodHyTs8VT6If0X
apjXk/MNOwiiwxwK1kBFHv0m0Q/atMFZinLtXt9LyJqkPnK4cY6JOkOcjMFdWLOBF1XYnqvMMgwh
muQ/ijBE5QXzTtWVRFRd0c8sodax4fcuKN+Cs7B20Mtd0OoMlPhupqea6l7zsixB3T2yJg1J9O4o
5bPRR5+tqxsmCup2PRPSYUyv6hXqrk0Y1iw8qavhJgc31ckCVaI2V6fWYFpRLZIKEdfn9qQ2Uovr
UGyt0CRtJDG+qNFI339VRf5ZWogmZOjsGCQW3w8SFepzPL0jhJ+vEaiNZhIp6wowIf/gd8JSeMbI
/AROLTVUcwdV+8p8w5QcuhvwhADlgYV+6xqHLznKKfZXz+6Un5qRl1u7+x5kl1OFnZ489H67z6A+
xw/bBat9EU3jizl2EP4hY4cm1R06aSJGpRp2zMESpK5di9+txm8dwhaGvgYdcatuE7OJxVLxrWQN
FeeGHfX+uth9FEk+k11jEXd1XQwxvJ708AYHZz1HbTCZgDnx5HrADkyWGvYOt3KB1ActaISHJibu
fQslixZnqxFCxl5izhGnalykPAP62OC/i19mrLbfsSIBgEggfkzMOZZ+nw2gNFWrrGbqqUv35jgX
wwAvwA9jDbIU67BwmesECYpFiTPyjYPDcWGfBlnfFffm5z+3Dff/xkfPmaUq5ne1koA1H3TQt7gY
VPLCYmlaUkgumF8MgZv7xRfa/Yy6taWNDJT6s/fHsgHZPpebG9asJyrNSLDF7tFwDkiUtXJXaSUA
ue5+Hx2HMod+sGtC7I8DzCSH6c8hq3K2gyF4kOV9WvYQqgoi15AppKcoUIHnULS/E+k0Fltw9r/K
nOEjmMfAAtM2GvfxYCYasujovrqjH5eO4G9AW4VgVIyfWq4vA34XjZedbIBJRfYu8EurL8SK+l5H
xJuqe4otx5KGY8bX0JKyBW9R1VXx9vx2BZ8EEevJTnCdlbCOMCzzirFkRUPMlgk+yhzvaVb56qAS
uryTsXK7y2wvsVlukg6IGc94FRig0VINyO9o90N6NUiz11WemCWLN6z62abDofMWXr5VTNMIUyZQ
nqcs+giWIh0yo0/nwpjOoNtxLu1Ph4cLoy5uEctBPT7Tdlx45IVsW7+Gwyl7Fj41ZQw9OLgd8+Rh
9KLPb9cysYIeCeYzoGfp/kJ8oyiPPPcjgTF/dpz+eI/ModdXgqyJHGGBLLvVfohdzUY2qvG71wZZ
eoKChLCN13dM/a0HJ2OM2MIUix8K9ZqXInnKEo5G7F3a6PMm1gRBoXP/NpWiD7CjEsS4oUHneslC
4ZmaWoU273xAxr4fUNjdy+yS71zWsnhu8pnfJexTA50aJk8ZLsZc7rpEd2eKf/3Zi9rTkWv9udIP
x0dmiL1z/XpenT6hkbV/dEXR6r7ZpyfqKjsKPxBY2yScLIOioZJrvMMe8hAhrClqJrxVjjTAWz+b
5P5fJyJB0D714mykiE7dmaYtK93PduwGDiY7FjXxDj2fTtCqCcvbAarV5J5yLPPb/rUkzVkTkbkw
1PYxieej+v/elEoR6WgDca8K7ncNyi61czisU1XJvgm6Fgve8QOcYa9KW+k9qNqf9uDd2o+TDO4P
xT38lhRf12YU5myW7j1Z3OsXdPPzy51LryFqgmwqOAk/JO8Ft6tHLpHXfyPZDfaRh+qLlTBMr9bI
3ZBjBae4EpxRA5i+ncDomZPqcJzqRbjGvXXR8RmCE7f6vIPYBbP5MMUfBUql5oPIAIWpQ85O4T6+
9/SVB8uwJ7eIH3XYl1u7+VSb1Yy4U3cQGfF4pFYok5RtiviFaKv7A0ta7D6slzS1CFgC1Eh4f2Ez
qcvWZ73kkJy1Y8tH4wfYg648mJD7EzquRqn5+PDzgyY8S+9jBNrMsNSW4rsEiC7WuySwa+ehDybK
6321h3/EhVJ2QstRBZY2V4CEqmHFrQOYYOW7+DXI7yXmqdQiWUb2eN0o4nWmp1SbPMlBOao9Y23E
+FMP9VOXHs1iMlpGWgbjJRIvmyL6SoabZEO/3n9Sg7aSoQmRMJad8O+lXrgsRZPEHXBW+FlYn0kj
CJ8r/rQhw/ddPh5Hm0bOT+ZRvKjntbxH4ta42GSt4uxHOQL5Nia0OG1AbWn6Oe2fVQqVkpTVoZIM
BNH6jd3BwQA4H1i66gw+YanbSLei/qbqI5CFVrQPtqviGjY4RKM2mK54Z3pjh9wuZfuatbSV8dno
ezZNH5Y2mRo2qIg0sSDdIms+ffW3en4BGUspw130N6k1tv1Rl6P6RDlY/6pJX81fG7tVPShMY1ic
giZp6goy9Ob3tk2cycgE052GJ2sSPsOTXj5kWnJAWUs1TcdCHohHirg8lge6ljpE8IAXHUUkxDdE
/glufFHZkdfPGzk+uOOTrw+CLQlsS/IdBpBJrh6bYwheaa2zXcNJ4W1QiqN7ooEuFvd5ee1v1wL8
bz4xJRlkjh7ikYJ9FbOPRMz4LQuQX/hMtoFXgFiLf+D0s2wyeBKVA5qFXT+7mOW6cklxPCaUHbtj
bQHBJ9R3Q6wEbIzAt8s2uaeVJA3AsYrdKTbfxQyVeuEzWOsURBBw9RtHXxL3MGhKBkINkXtF4APv
lkppy6Db/P4T3hYjWSdzvHzr6L8SobtTS1bblVpHGqnAzwOrlBKxwXDr39hkegokmJlg89F51L63
CWHUdNY9963JUcdK4GW5DklM+vOCuqR2yoI9/BODjoa9IYm2LS4/2prGbyDfmL7VlVqgbnkXfIdo
WNqJf8UdRef6g7YSyAk+b1r0H7OP9IncsL61wGN7hMeXq4R1ehkGBypsLGxhJq+6ypCs5T54dezj
If64RBcecAieyQkpTO1rD7AsoI5+vb6GjOJcqczxqz7QYdtv8NfsT4FtnTaj/5io8B+u3TXtzqX3
GwKcZyEcR1xTIkkOpcLEP3V75h7HpvO2W8lR3q/2fiBpbrrR77WMWLFtmfkgdkAzYIHdqfWmp4FZ
nmKHwqSAvjiZdpWzxZipLyu7ABrrD2LXooB6lodnPH4j7xuCyu0xSGXoxt2MxUvtSjVzlviFNhlU
n6Rj64bLGNY+nFra/lAJ699FWJ70DWaPrJcGNUSWz2ex+m5S1c5TVo5TAbV5fcZ7O2+eNpPU8l1T
xZ/muzY9ZlHE8fNfdKUc9waJMCDj0DRNlZpfC/VLkjAtPIQU32JqmbtR35RsXll7pFRky5epok57
6m5XAncpsQ7Faftlo29v+GCIMan6HczavWwBClHfEAhQrrN3SbEwUXLdPdVYpeXKhsC2R/aCU4O4
pyc6Oquk5/kPCCI8QxXYxzwwjP19njHTlVQvb7DXncHWJYLwbKG9YkYL+jQXfk4MXTXD5oEefo+H
PjhCLk82GoP/6+7ecbnOcI+HAzTUZWXeMjj5mea8JpV4HU2eox1g1iQBEEq3yjZ5f6cpxVVAVISA
obyWXCGFsuaj9I8gM0X0Jzj3LcCFXvKSxwyc3gYU9qzG5C26ubA51Oo4sKGuaygrP4Y2QSCq62bu
nYx0iSFyIpkrLWggDdRaYUpjFpCbuu0XVepPSWnRhq8AwFl8EBcEj6Nz+4n0IIZShuopaBrb9Cfs
35kR96TlCYzcuRlmzMa4/iK4FAHx57ul8hqnNM2VaAJ1W2FqnhyZhuuFxNdBGD8aR94a6LTktpBI
4rHUQm9KC99N+56iWudXV8Vxj68ls/ODgUnYOjn5uUFrzF1V0TanvMTyI52DCi+CDW25dmoHjn8t
Fh4mnNfeIwYxOc+7jgjCkc0Hdx7i+5M20McbPnR7xVhrIQswfiBjvPd/+mGnqn2GPzqVt21diJzB
jLVDKuOq0GUSv1roGwP13y63AnnR++MNMeJlYbod4Lmm9oa31BEjonGq/NuFTkoE0cpY9eeT93K/
GbPjh5UZdwAB7qKAsZX5GPvgFPlM3TGkLnzpT2FU367o2Q7Oy6ndPKC54NB5G2dSBOrswQXMa1m7
yM5Oa//nmLjnl1lcDeyDYlGNSQUXKG2qLws1g4BdHWUEFQreVDh9x9Tg98WIHsvsOV+JtKV2qUKZ
zDoAG7m1pRn3rjHoakZomrW1vzeKtvau8ro1TQajkBBotRpATeQrz4C+blrXtwcEKuNldjRrM2wu
KKGYvCfpGwdDihAC3eRTB3eoMu0+4IcBoAV96HsQyDD2lGJWa7/28QkESupBxeO2HNAyUsinj8Q1
+vh245GxzucKYkLUATl4VvoMASqPN3633YFUX04y1yG/JhSwucfccMIe5/Gj3YbkxbZFiWvuvxwQ
O8oEnXQoq8gPbQPWZrF5uLNWUfMhfEhkaw6s7pd9cBEguvM0IE0TCSc0V81t+S0ZgJdCb4xK2hQ4
WZIBE63yq0QOsQtFcXAAlL2wVt8e7jyU5EPuby3/56wC22ZlPm67nhWsmeLpRcMyuRIxfmyReyim
759KM9a7Bo4HHidgWTMEJNwKUOrbrT+okY8dE4UHr60bGNYhcF2fwUCuuB8s7YSDfidMGOWPy9uA
ejmYNtdmNBhTOx1+Ye+xqT+Du779q6CKgHw7GUsk2zTa0PyRffRJlRNgm0UnKbKQ1GQpfIJ55E/e
DL5i+no16rcxXByzO1P8lKX8EUNrgpLDs8NQHS1RzbTLptKAik2gd3kW/ok9nVXw9SQMZg5nP8Ij
ISlhXjJS9dhDzrpwZxfxELjUbvqSD12UuxS/wPDaFu4E+GlTZWJ2vMoitztDQLTlkfeRqO4Z4If3
5jQIqLicJYE5iX/D2OfQof0L0vKp9L5vZ8XxiGXGEhhaJ+EaTzSMZzIAzYG/NQShpZnr0/9ub57G
75hnRb+iSq7xN8v64amNRUqXZJRk/03USxqhTDflmDc1ounM3s2HxSC5WK+Y8atWZZon4ALrOwEZ
RQkXOPSNJKIX4bmeIdxeHmgJj7n0tgyZeLop9aFEPiwGk4Fg2bMBg8fLinQQ6NpZw2/WZ72Sz0PM
tR3jWtvV5YabFNONh0NJeKqw3UuP36iFE9+DhV5TCLGtcGcwEDIhGXNw37jQw+3/L5L2IhSOLN7Q
rDWfYarR4E5TJaB7P8PyRwvDqoDBRQ4RyGJIVApj/nJI47HXJ7TpqTOEeoEivfXSCFUSSxxGayTn
/uEc08srAu/jSABw27fpae4KIuj5jtxiHi6KEVRlJCKH2MwK4mH9S57v057iAt1JsyBc/hIARqof
hVGWebfE5Mh1DLvJfEjorlJQavw0creRxG/Pfy569SWgBfYMBFfMMsjxWBHWTe4J8ONhGH30gzLA
TFCDJegih4Q7v3/wEmJhiQuCO+yc33EGypi6cvmOJu3oaeKZ1iwwHdX9uuLEDlBilIFNhzc4BTFJ
liPEQl+YMgMwL3YlqqaHkjqHUOraBMyGMrbFsicE1fCN1LG8KAK77olXdmXMt7+ndPco3KXRBYgV
Fn6B73BndUcaKorpPr5EeyKYyv+c2y47lGtp6WYeyArEtNwCAkB7/DQR0cjyR0sOyihBt18RDerS
QpMLrbsKJtKe9Hi6Z1hG89Eu9+hYKKq10nsNbrrLWaJQAlEAKM2iWKznellNbBPnWaVblC2GPESb
TMFYEnaTqg0i+L5oTDRoy2Ssumr+qMXBdvkMZ3WnNgQOLGkuJoG1emEu+X7MTYlkiwv5/nR+JGSH
V++gVwQC4PFKe9i9ysXOZ86e9B+mTGQZTsY3lSAEbdz6rYrvjHTkDv8cCM4EziC6kPeRqTAKIyL2
Lk9VBKy76MbfKD7Hhmb0OzpRoG7bqDMZKnRWcLWLNhvZzNwbLo9+U70I6HEGufRBtRnSB/5F0Rmd
dICpCU3DJzKRk/kMI/Xcw6gdvx5rK3vA9VvxvfEMtP+Ir/eumMb2D2kw1HrYql91B6ofK2CRG78d
4MSRJoCK55jvO4pHYph7K/lWO21UsiJWhoPr2NBvXI7cJqranCOEa1weVhPcpcCXtZanSkDVmGHG
U/2llAbopkDAy1IFXNycZyuL/2/klgJI6YogcSxDrvG1IseQNH5l9RKI2ZqhZ/1cMwOzrb0rR/dJ
VAQCeyMBVpiK+nmXIMspAjxsKqp7tk5gruWf2v7dAQlxeDI9MURFxor7l9iMJh90mXmSUDRStct9
xpLL9y9UVrwqDT7rVG6g0V4azJ66Nwg7KDRSciHqVihN89CtkozrP9uwbAX4hrKnMUBFmyeW2GX0
bfYu/hjYqFcg9MJdDdo51lQBkiPNKIJqT3PxkgJFRhIgH3r0aCyW5ldhX0/J7hadD/rxinEqAONu
/vsmsqEkKanjC3BCxMKmsemDLCWToLp3N/e4HbR1eLJecLBUMN6gvPJlcxZvkEPTnoKoZz+cVaNL
knwfqqkCynqctu3yxOg5OANIuQVUpN5SzgqzwD0IYsBqw4ufn2lT1M9pQd6s7gBJ5tYiuqFGgx7A
Qc5CkVsfVpsekQJkNvOkSoDXcXwymE4d+j1kcDdmHTpnP1ywX0OM06ns9/5jDyDOIy1cWcjg7hzt
kuLLg8C3vY9gD3IYWnkmoxsn7kQTwn5Z7FmgI73Ho757MiwY5MiZf3z1BjMZ3OaKFS0pwpu/zPBB
aYe7Ps3r8MLo9hPEOKZUQ+PSlBCP9vCAWOkdN4+3/K2EEjNy5VQiif0l36vn2cihTfdKGS2lr2u8
6tQ0+di+z4kMFdf7UwAyt9Tyf1VLW41h4yzW5czMvp6Sr359F4jgggUr5Yh8WTiL8CABG/8nJa6x
CbBXgtASx6H4gE1FWGjb+00564EsqtryRt3QUVzScG8v3xVAvYfBMpQP3PgeaBobaqfKKgdiAoI4
ggENjGSiA0LblhVQYVrn4Tw0s/96gR6c4896d8WaQm2KORVYKzdREmkqvH5t+PvOEfHpBvJ1oGAh
JgIBdrlktzFdx+RINizDOwRNNMSwHS+I+pzQ9tD7NDqDIG0Eb5ZsVV9Abbr8W+zMNSEDQ774yO6l
54mhsdAFIxY/u5KTneLDpkTuNodvHcIdytFXBpbz7qqTLnir6+9ewpyQgV/AUwPq4fd5zYM3j+pd
q/NXrPYB3ej5jt7liZpq6LmnyaD35T+02S+Q8FWjXAbHrDvx8bOlVyHJu3AIjjNSrvqx8L0dD3hN
S5ezzM5HIldUB1ss2c/tQXSxr3y5JquadPrM0kEHp2kWrHxpyVHKZ6E6DUjzF7VgpWFejwkqevit
1d+jA2CgTUIA0mcgQYhq9M3CYBHC3miMeq5U6hyoqMUQbscqlVLXctiLp45MAledo8Vjv4jCEDpS
9IxtXGKBKy/+Fi20ozMBVdz9QR4InBpZ/W2MM989tfTSaVj5blwAIJdCQKcvsdZz14QjWcoG7vHi
WBxmC+lTw4cRyVjvCVE23GvQEO9G0GXMI/8ELBq15Wy23kGFopdHcAMOos1icGJmUdKjC4PSEFyD
eqhrMTT8QMCq5uHoELVbeYfxBXwz+i1vdDhplsedsAe8zuDidu4cESysTo4rLP3rsy+d6qKeMCUk
MLnLSzTrK5Ma7u9v+ZQG3GF/3YHnYs0dtfuVl5bA2zaLcG6kSjsbzyxJ8pVcxQnVtwY7nk1TEBo5
6qTGfLaXNIzziI7wGm8uKwM3uisu+B+97n3ld+QXPl0psKQHQgEx27Qx33GAbx+vn7ItGIv13fNt
rMyoALjZC7uygKCx6gOdkTTryyggsabwbFTV5YcTtDHqY4iXovVBjo5FAVEXMdZKMAVIXbk5L3eq
586pzS8fWXIBZjhtYW6dSmKkMeLj8C88OPyuZI49IBqU5qwKwteuHP4SWKN7NPvI+3OUttptL5wq
xVZsB2YN4ZbiddXgaQEKi+UtRTxrTdZPiu4Swd8/s2DyXIk071Y3yqCIpb3rWkq4YTbb67F8ilCM
ZcQQ9ZGz3jI3q5jC0zB5t/xHZTgdN9Shart85rgMKF07vQ/2Rhfgchoj925Kb2N2A8hAUaApaqr8
mha5Ir3AgWz+1NW9R5i6Ei/8vOW5oqXgJE42QxUT9SGu5r6HZWYXmmEdUa0vExSMXZBPCHPCzl+U
Nbl0cMPkHssXB5rXYyiQG9N2y4hy67zU7Lup7FxlWsp+v6o046XkJ5+HhGgZ8IAxWXk95XP9ru71
I57wVBxkt8ioD1qIchuiOLjWedUc8ij327rlEyWcwajJjmsS5kGfHAv2LYy5EJv0TTE4IA3D+tQD
Ep1AubUi9Lzb9il2N/Rscre1uO5OXKYFZ8Tp5AGR9fBdWW8mxh2yMxJrKOzaYqQa8RSNc3x49oiQ
yezvmL4qK4WtOI/LIKQrdOhmLmBcBq/PynqCJsIfybwOBOkrFQtV4gbuUtmwa+sxVfdXC4U2MK3Z
ZXq5LsJ5GKUWqWigztwvRE2dzMbQod9zcVcgc9GZxWoCs21IxK0NUO3QME/RDoo3SW4ivwlcBWzd
Xd4kgejMTHwWMOkTMK7eR1SDHO7S1/2Az+DTwqB2/dSH1d6Zx/uy3sIee/1MnKb2KOSWtoIFlEza
ZjCtIQlflukSnINm2VTIWcwFozxd+o3MFwWLPtb2FzibQCMq1ytQPKeSmjcy+wUNdM0l9VOZ857O
16ytoblaGlMm4WO3YESmbEWD4btCcdt2BH/5q1E2o4WWCZS5QQpnwex/4vwAYCxUpeU/0rqM/kav
vd+Ppw8F6ZajYdsFdnUjU7D28oKC/LSOpDhxr4OLIY7qqwZywMT2uPrFSXJ0McaSx2JWwHnbl3IW
eAP0rJ3b42+zjGZi39HRj5OpS5Lj69XC3tYo004Rgj4EWrnNu3BqT7/iWS+/U60QMozHImFS4Ame
a7ltY6b2raoSaWW/3z7HAaiSkASKknxIdaR0ypZ5oLirgQcPOs58yFKwQttw0Z3FODSpeQvxb0ac
VJmoqWm/4cCvZgwJwUHg6gk9YTdGk5sCFQk3PuL8MFtGlmkQ56Ho73qDgdhnKKWWPVmBuRRs5tQN
XPt5hAZs0w6Rt6VguwY24po02lSiAoGtdfaBoGFF2jmvawKI8SsqkO7wJJ0HKR4QzViFjLaAujQe
miG5OlP1CZHHx7iWizGGSSbe506Vu3Eqssi0pzen45bPSFewttZxzajsFzoDN4kJV00fLIEVLC3m
jKVkWVXllNqwXF64eDhCDruG1n1XMrOzpv+SVx7wtdm7K8kovEZDuXnupfYUSVKjkRGUg1ot3pAd
tCl5FoEe9UMJjHfhvmjHjwc/fWylWzFwSEmrcqS9ssKNsI5CE6ZOU7iEXtz/4aNPpH58TjRzrsXL
ZOizk6hrVB1rVPOlYafM4iNlXTuVB8lZqTR8XOes6zeizMGeho2DrKWSB6EIqnBLD2F+3ajvD8Gu
X3K0y1P5b15Zx0EjLyHWCQez3h5QHQ879Q7ME2gcO3N2+8kX2ec4VjyikKj4HwXtGEydkXa4h11e
vFg04DfU2XlzLzQB42tmYBLPNE5uMTr5JQuZeEpUg6lJeDv73I9u/FPeNfeq3WBGDhG9MUCJXHaH
88SgeDAdc0y0F7jRqwIXkPeYaR+OYilhxsJ/oXljn/iWk1/cSACNZoHDJKsvf7+hVo9hwXEsfJBY
GMNh5U7tO8eALcKZAsa/2R+ni3ZgpvvSM4Ov0HKzECUdZexJg/EagC3mopc5hP1ZJfunkvdOSJGP
cO1aBMh8FVyysq39QEXHciDP0lGHAwIIPmDBptG24yZz3vWyqqHJBFoqADs2Kewhbp3pxqO1/UHy
8sXdSZfx3oonVabCetWRybHau7G0HxwUBiNuB5UAS/AsqRJ0e+Oo+iACtWDznu7ORrOmgNAPWfln
cRaSUoiZoCa6tu3X7Px7cZJaEOiYSvupSD51snG++25u/4gsJWAF9pGwJsydrisdRH58Kixv14y6
B9mYdWyg8r9GZl2bn0tEnPZQHRIUMkmBh8+reue7R4n9YRVfhfXZP/9jAmaRzOpFGmjjkh05PZCD
+SBfFQRNVvNUF3c/gm0Hnjygrw5OKFMlMmiV6a3uhkBqAgMAwK1R2wlBbeWSBtfODPIvJ/UV1IOy
BgifdsNF5Dt3KTg+k3JmbNaQRffsG8rEAM8n5SqkI7ZOgLQN7nhWAN4pl5+3rx4LKajLPB4Q1Sn5
CF2ZkSNT+u4vXdbInJPRP0/doFTTY1bBln/xwkNcY+m/vxJFK+DoLQR6bMNLD6IIuxgpfKVGTCDQ
eQXpxhbWNRY/wlDjubkI5KGcxxdCm/WsHlQe3y5qMDO/zFMmItF3KBzKqIE8riw3wO1Vl6MrEzM9
Qav3dEKqYkdmk7wkwt7h0ammkUkVR0pW4l75CSpR2vU9iFsgX3obDiLn3lpzV87JT/fAzLIHLEg1
mb9RSK82KBfxZoqhBj3ax2XTyZVIlIsQUHwEF6x4EEVijoGjS+swRJprNbpaOQU2A4QwP0ODim0S
g2h0OTxbNr7ca4RorOnh2l/td0n1m/UunhFJVjSS7elsBL/4+MsOWklhNGNiiqaSn0/y5A5tHbL2
u9Uij5AjcEEEeMcsgRi74YgDmhXogazKJ5g8XQElhM/esTRi7jMGAVSO5eX/k7S6bu/XGpncmT5M
2AqiiwA9zMCiDoueRb7DgwCHR0ZH3gnfLfj+VlBtvDWkIScK8TBxl3QGPBHaESb1udC9PtwxWPHS
HPFxLLFO3SJN88NrJvYT/sEMcG0eBFfWOlJABTRSHZdE7BRwdPOXYmTq5KNJ3mYfSXP6p7NxKkxL
lOqYDkQKGsXtQAtnK2EBoZJEl+Va69bpxWQYS68MAUdrwrk2I02THTrL8OAhblZR/TQYCy2Snd85
6aMCSIy3kXnSDaN4eoWoVT0LR37CuGjDsB66CMFI5J2OICYUO0tkQ4SLyvjM4Y/JfyVHvI2vyyXR
ajKS6/nz+PBqz8T5bRUV1r1d7uNr6P0ni1jgd4GOe+78ECIBX2QNe7AmUmQsALzvmbFAVkiELxFd
QeqcEB+uhpq6HUX41E5rlEV0r7I2Nr/lbtFZuiy19q/Qyxm7K0gbKH4dT3NKVUGDUmZDIbV6JUpD
vzTTky/PKU3KrVge0tArRxbWfvhmVGoP1iKA0gAjyLdQbp7+dZmq8o3Qqv0fbhiSvX2hIl3lefn8
8Bp7t2UfMO5tyo/h1eIOLuJPx/wZ5pB86Li13UgsXFhYa3F5cVsLBgTN0VOzoQ8n7vM9wRDeqXaN
yrqXavP5+O799/euGMutlc5Ws3534HrmsFPJaGjYo4r8lik/1gpD9fdtx7Yis7v8j6ccNXnmR7dO
wh6V3VeHuwOpkDQOjZEDq9FPFhdkI4oUdt8GzXTcXLgdBL7CT8UDYRZ1SaNiDHZncD/y++d/YGFR
Mrudie5vm7HGNpqXYBMHe484teFnKCcT5gbZO9Jh5M/97kviOmYdiq8Nm8SG2d6eGS+JGGugzipz
iJHSBQyy20d9WaHum4bO2OjZ9SBjjktEEK5ll8RHo8+QfLkTOigOUMAZz7rAFyzxik3iKxqd+i+x
QL0cOIT4OqjasdChscuXo8b2ldriWkzTo0NA2qXmhpiTeqC3nFHNqW9bg4FfON46Lgn221DMN+mc
ieOpIX4m2lx0o45Tb5U7NY+ghsXFvbp3yr5s+6Hn8pED61rZnVZi5w+3bKIDdWhmxZeTl325g48l
QL9ATc8sZzWFOWcqGrwbhF8uDQyM7WOy2WyuWr/TyhpjUWDrw90zGtTjHPuZ/nYBP6KxhQkCviw/
0hBnPyjLT8v5+4PWJ6avLApXjLsa3CkRSpo3Np2wuqzq1ct1iSO5FIDnece7sG2yvEK2s0r6E2Xk
cc7YlUZ3BmyQgNkARibKULlpzcMHcMFTk1plZmchfv119eyc8cyN+pfGEexjVNkwOb9wUDonxMmJ
+KsbCFQ7yZtKI2gxwcTZ0gGKSu7COEzLT4SdrbnO4Mwe/mit37ziN35BbOqXpALPRED4d21+lUHN
XjfmPnKv1nugjJj4GB7bqMQFersfAHilEGCzx2iUpdExP8OKed6HveXc9fteMrvjazQKjPF7mZgM
BGc/5aEzc5puwh20UAz9AdoZg1Qe7yp+fCPycXCqJaLIN7zdxldyZO1iDUcW6Mz7P8ikZ4nKrbb1
eGlGxi58JDJB2OHEYbEyfGVjco2IQaYUtbH6j9rSKXXOjok97bJIxcv0PDJ5SUG/IQU7BfbldP0O
R5IeXFyLRoBXFa0tmpxYN9x50hP3qU3QGoTTlrUrcTHoggSnaP8mK1COMQEoh6pzErwduG/DUNRE
bBUMj2I7CcKHuE7z8Xugo++dTWZbIEgkN0nvo+PmRRNGpkB5ELHH5D0Qrf6yT2qxAvetivMZX2+R
WO4oPgMcuHGHnbrkE2qTakpAk2zUTC9hPRbsak6/LPQ/rs+cwvR5lVoTa9K/6LMaO89hOCtZS/Z7
tkkwIO0mtVidNj+m3Hnz3tjsNnEQja7viZBy5SndH34lSpNyRu4R/HJRCjsrfNV7La4bsb4o+ucr
5XmJzi4nzIoE5lfv8Who14AV9rbBeUGTXIM+Hjf0DKSeAeY4sUHLGZXJVlo6bbV2jLP+qpmeclxm
WPqGIvUhEkBiYXE+7m4GYU30zEDzK4szWkYeOu7DcrK4bcdM449nP1Gp9kmXDhrm5WqeZGapU2GN
tiNtnzv+ZCKLYWUu0XQysblIPlc65IpIqDPzYfAXjT0Gjt8i/oF181zXmrfJ3CVz5Rk1/9KjmGJw
C3878K0lHtDXdu12qA05EqmNWkaAeluClJaWRyVdsvSftJw6EkOCA7PxnjLuoslfC5kkwT9Gs3Nh
t+Iqg9x8m3arer2Mkr+8NTZuPkxmHMfo5/t5xHMB0QY1DW/qSQtJdct3wJsVG6O+UNuWH+wLcAO5
ESChOBS/1ub+cJdOG28msi7q88DFkG0F9wEb/7EI7tPPgvWhICmNEKPRgt/ezpQJUvmdbvHEdlGN
m2y8enZdc89yby0W4luotCdki/cKhc01JsMe3nLlouRorhyzXfW+53tw1wnAttTs4+5fEY4Lle3p
Ym3XIPWZS8DOWKLsNgIBQFWD24/C6UyICt4Sue3zONN9igbLjoKUjHWWnwFGzgc5YMNAOF2MAkDA
poGiV1PijiBlQsMQActHuZce6Y2BdF6pH95q/xppQmzyZ7y3CdOArZjsi3TmmfuLzZ9R0CxCtq1N
jjnwnO2CsRJvEMhcbr81HwjeL3u6HxSiZrxM3jMN+ffOc4HWL6feYghvhmlFBvYWWxiw/rkMRfv/
LVBS9CRPJz/x+6ERcrjwvOSTYYX8/TvwzT/ZQcHrww+v7hZSLYJndhwMmlzSF5ytPNAGHegBycru
Mee8IIAPEILM093kCw8lO78j+eKPEiuOFdRN9PWOqMXuiOfA8udP8xgK2IxjpgmlfXlJ14DJ6uKk
TOptIVf2CsfONew0ASYqB13CKqPHPgvcGjSqv6EeU+zD8z75SnYbqrYPtfCaX+eVpNe1mx8wRdpa
3z78UPituduMk9cDva0TuIigoXNY1fuH3aRYkoTl4e3yZZhqlN6OFJ0JrfOn34s0eux2ojfyPSPA
AkekzMIdOXjcVVEZb8WVFM/GC0a2FDVWvB7Uv063GN+TsHlRSYQ1BZLpXBAb4KsvQyBwgwXPZ2hB
o/ameKxylFwxPUBJqih7GbQQ0NeuDOzgXOfh8A4t9n3/70nh5Rzc8iM+FOgGBtvRIaZB0mnJ0yXE
fXcpCK4SltoXz0p5okvnCCmc1Ya0gapfuR8nTyBewdapq8cMpwxLLVZUkqeB/FW9uHy67WamySHb
TaYzwN/Kiwdl6pS2Ju53b7l09efL/oK0J1w1elGZsM52p6CMsJlg+UbVPziVJIqEdSycVQRgXxfC
m1OvqwVIRrzg0QwkdUo98qdy4JYtPL+M5kgb3jEnQSzgg2DLemalySymZyE2SFxRhfFETt5tl+lL
wpUfGEavpPt1JusELqEtyrBlYbGktjaXWGRYwCEn6XEY3w38PqMZYR80y7ePI6bxt3sRmcLMGskU
nCW9Q0iexeLEkeaL+cEIG+VGWYJ+XHTnb3syM19F9ovGPrc/YAcjkI4CYsssZkQYfOEDhlVZYzNp
dP0GRzPdPBEgKasbMAUr9LdyBLRZbten8nFpXuvzVnko+QHOOVQY7kSu5mzdRcroYyejtWBTRvuM
xTCLZvTH0FFRDRKD4vBk9UtuIOJaocK/FfY9KdUG+WH1MEOHkN9Qngmx4SYx65abqHX/aWP1wRAb
cGqdm5eFLjXkfKqGHSoVIwRrjlrtpnmqYj/BPynWfdIZG9Z6ClNtf3v2g3/34K3R2uIA5BoPHa2p
JHVpJu1LxrvxupMAygaly7zfEZC9ABHbqCD0FfTUwC343g5OG+WuI+/u1SjOWDIb8yUvnynDQfNt
gnr5VwEHgQPLwlZVK/24thj7Z/KfCU3T0foN9iTBDnEqjhsWw7NQcdMqWCFdxqoKqv6Eouw0XG84
opxkIoSALILxneilDBg/TDfR/pnZitQWFzUKWAi2hTKHV3tj7xrOZrGalgVB/Ma3LzsvAykGC9Bw
DkHzYNOU13hEpLdhHllYvg9QERhmk3XcDtm22u7q/Nvxgv2TWUPYPVoMrf+EkixZ+ctpAhlzF0o2
ALJu2q8/J8y0CEmqrtpmPgfquJ57rOe+78ciAchjH7hnQGDEAnBI7NvuyXVTB18raXUACyDHgQ+f
winLFEWTa6KTIUMfBoESuXkQerKp+re20/aZ3P7D6gnRm2Zicx4zikAQC5DBM2KNaD+U+hxFmjd3
MMMe1jbgoIZ4MlR8dNNqxFo3zjeD3Kp4u7l2VSigoX813IrN/pUc5BORkcZv0nUss75dgzUYMGqT
Zc+oupZYX43mhJLNJwYam/WWdKu5zOVZqk9696ApG/fhfpIaEVuVQ6PtyxRhgyC+mSSFZeao8FCm
FIB/8vwOik0MZt7/oeWYAyxUEexXJM7fKtKXnaWbd3SIxvoXXAqRikMxB8IViutuviudAU2B/pHm
pFPuSxg6F/S/iXATwRNycB3b3khVbd32OVfkEUS2oe3bjA/vyN51lHV+89DVwaz8eQ5rKuej012k
PU8aO6VOM/eHXuRfAmqHqpT7DznodLJ3sqdaVTxU2gztazXabVhUa2+VNPoYTvAxThaJzF8O0Ej6
DTymOeleNK95UC/ZRxgsdMK3lddY0m82528fJmmD07Vnaki7hYmLqTd8/0tAgcmz0/a5pMXFDy6o
bSt8KwhWdy9jTnS9pJV8hKe9KZ93pP8gU0vVb7Y5WhM0jtc8rQK0XnDttfS6WKZ2R9Rw9xxh/0b+
6TyvmrpwDuSJ/o1ejO+t+X+aREoe9QMg4ZMokNJNC0iXEgnmD2IFhmoqUALrJmJnOon3J0v47m+z
qYkSEbBRyq85nYnEFlya5u/Ah33dWkUSYd/KkQH3duERAwGwGABT2aMx7p5SUtBw4BGJsup9X93E
sPJYp5iraAqIfq/k7pwfPn8mgyUKY/tNmj/KhssefWGga2DYzoTuGqTPIt1sJC7Gsn0+7eNitbBc
hOoBZGE77LdqbMYNfVvOfN0tyb0Fx19SSTtEz+BBQ3AjreS3sanfHkqrfzcMhZ5QyIX1AQhFj4F1
Byh0bFTaPAa2GY8BIKj8bkR7F/XyfzK00CsNWMsxGYLj/Fsr549ebbuw9H5FBaPLL0Fv4gCm/nbN
GVy803ObCSl08O+hck2z1+m1RkWoLVJZ4ohLfh7IXbQDUcR2G9iewsaz52PA9erqzuF8a3yE0pPS
mEsIbfUk2ivH3e9PPcU2ym6vqQwpnz4EDBr3fqYsGv/jEDCVxatBXg8CS8WIZ151XGAV0+DyAIXa
uCIviSAAoFqI91gK1iACQXFYyexf52Z5k4p1vdTJg5GFuOrqKRzfKEKEq5+yOkiAG/oMAXf5UjLG
HyvLZLr1a42yZr/Z9xNv4InmemCToFzbdnRj0WPGbCXLu7YHWE6zQrqijLvf9W8Ovm57xGTqidN9
8Ls/rnZAW2zlWCapc8axjWHWV/iw5YuYFY2FUFuXsbDtBnfO+QtMpc3oAEl+8+6C/YEulKZKaQ5z
UpJdXzF1Tx6hWVbIxUdKknfR1GySf8sozGcTpkv6NtPhHIIM2aFKSXPb99cl9CoeGG1fUGkaw+ZL
+EkTgUicuBrzMd6SL73287f8hhirpW5mCy4drOrpybY+iEpnaIGbiwvHaHTv6ax+hJqfJNWz+/6o
eMO55ViORO7U8HK/P7vI/WeCpMMhvzwfDfpuHK17ADdiq8JJw6+f1l5ysPsgmbc01/F1s0tN6TmJ
/UCA0NTsk0rxqeEd3M2T5zDmj9kk5gqVhmyqDPyAmT4tKN969ITHD4ZAhC68U6pO0CrfA5gR87QM
5e++6CSvo5LiEfCQFhFCan+siPQ7LaW0TtqJ1dOPUfTw7NeVvPNn5bH92Ksejz0Mj8NB3i6/QmAc
LeoOWFDhIUxqPFTtbi4oUyR225Y60NzDF9HN6CWnw0bemiDVmmToY75Bq5HwAR3AmJWOWU5W64z9
hb3Xw+yTF+AMuYx1Agd7uXwZDaUIAQAzzAC9cv1XODd807AChNUCBEK++QjzUMw82jgXq8ao3EH0
dA3dLxPPiSjWO3AShRT3me/NscCJWWdf5j7+GNDY5cdP+72A+g15DW6byWRH+GT3ywAiSMSJYV8t
Vf3KfpUgZCNRCMvWiNGQI4ckFZipic46ibEOgPb/t37Z2UbBSD9by5SP+JCYVKs7Ch87PlzP27Hm
fbCpsxAvA4qUZ6FDRZwFYpx8ZiV/L+RViDC4wRbRdd4C3f1vHqzujQVsx04cUDspdO0cp81bnaFC
bagsRP0NlEp2kpdXzzu3pb/6jcNqyJhLWGYraXKtnTZNtChX5TLFWaBYBXAggCuTaIv3Jq7UAIxs
kDisyCdiMiDKFCYZYAzmSGen0NIXWCvU8/+6lvrF0Z/ZNTO3V3rG01oyyquY/1FwzO3W9CarKLKc
IOsJiCO2q04UglE8ZoIF71yfRCVABxT2r5W+yiScukOHR6gztEzZB9XxP8liIaw9rwFx/fDFaOE/
o3icGQY6JDMz7SxJZY1UK3p99FEtbTfpjLyvds0veUYFxp+NCBtyPMvC0EPEBPbHBzVyMOokLKAZ
dGXXUuzIDFjpqqtAEdMj5W/aoSstn1/J621PNDRElk1lj+VqPGhoMRr4WQdE8UIekw5/o5C5pvmB
5YgXyDJ3fQ+0WgUaB1CVqWAs800SMi24tGRSB8QnPSkCcWdAknp+/6Rs1DJiQfDk5qOKfECsQXrU
xT9CzaqPwgjZw+43q+gZ864g/Pp1omOVOkCD0C0OS8F9rdKOzTVC/xPO7ugMAA7CpR16/fMuo2ZH
eJRed3hbZX05tuUx/9yc92G2TiDXywW+dsg45Ko7E6LqiQ/zdt11jFyiFseTRgIDSPmN46yVHodk
/ZrY/k/9kulayO/W274hTgv+iqSMMm916HsR0V8FA7XElq/92/IxLsfhghmMKsUH68QY3d+6koZx
caTA1yuH16ixUzQvxztgefqpc41G+mQCpcfxyyE4Nebmi8F662FZyZJtyX62ihUA+hd1jbz9RGzF
poFxFZZn6FS8XFCwsfUBLL7Ot1o5GV7Gzm0F+RbSpMP7ldkG/gB2qfIqr+oqozPFLskZLBX2Ljv2
YsFKYsA+IdH8Phdh5vlsXVCwoLg+tSj8Vl5rS5J3Ne8ApwuFWqZhGUNdg5eYeKOsSCpo+WHOS0nn
yvUGVBJSobHEgB+LSrNWAvWxnwOm+HywntfXoKPuEMMyYN46luiFSwF/l0Gt6YVzeJrpCbfJrKHW
xcYxm2zk8g3hHRenby7qj/XscUwVeHYNbfH6wfHWXHQTrUllZu7VvLUosZpGKd8/LEjwZojNgE0q
ZiPRXuIY3ujMu43ZSjZm95BX+F7BoBKYhWMKFd+fhFSTb9+LdmrvZ5RBVqVM+uS+P7aByHP58WJ2
kWV2rbmWNVIU3NtIIaCuldUsBgHjdEcqQAHqSZba5uVJzKsLReNsh0Sc40AGtKA1n7WPqYW61jLP
OPkLRm1aW5TLOCM3qc+nVx3ho3imDWcrNPY1k013pW9q7J0uIDcBHpZVymbQA6fKGPlV5xTEtVaZ
txlLJ0YH1VXIbS5bf35YxYBeteFaGP5dJI8h3ryQSj47MTxibiVrQ5qrhbPh9euvgqCc+Uh6unCN
AYb/FaE7Frh+Q085TOBoMKThzqG5SOyeuJkgfiGosAgYajR2ttucne20qmiKOn95sx3U6cQFBh8T
nU7oL7sLwb3Lj1GyEgFu5cw9JVvjDCzrBT71MbEOlcHTfhkhh7ciPvKLOp9KbKRCV6dHfPvSnRCZ
W4COo7DWFyLywAODoHofzb0E0NttTyysMohWnHs1wk0l19aWT61jhBsTLq0LSLmDoOtAfzsT7xXx
JmSIUWyvMqC8NM/7hjMp7KWHNZ35l5+Gg+KlSX0wlup9M13g+YHg7LhFfCghHfmQWqKXzCGu+5cW
23qSelJQS+blIlAZrRb3R0A0+SfcuEqrkuHbNEzJVl/iFg+I+6wAiFKD3yiDxCNOwKlLsxMAJ7sX
JZu75Kblnpmzdr3RLN3k+HyCm0SsNB2C1DGgLujhPet2UA27TuAEHuNKsNePy3r5aI33tqpY7VPH
xhViXv43ivGx9R5jiijT7lJh7gCZ6jxl7MkMNn63CM7YRUEMpOsojALSs2yJXH4M2iEXt7yLp2No
cYf+tbN0wogmCCMjiwM7rhpzcw5T+SW/nZH3HcYSeKZZoqigAImIIXx1tyTv5ALnSq5lR46Nh7wY
au2Bz7peqPBSUsV2596/zPxnLqa51LV6m13qkhs9MiCBAxw50YW3bLqARNZ94AwTVVvm8NJpTvIE
t2tbZRnZ6mYc3PkiN3/DNiSIBu9Q8YNEr76a+sDSELKuPvCVUMyABCokvF8v7d2hPxqrBbo+o23w
nR8SpoMNHH7c8H7DPraFKkso4ZZZZySTApko05q1oNeGqzI8BaWI7NmJk3pa1VH2xXa5bG18YFkw
UvzuwcyHFhQhcmvp4O34P1YAp7mgXHo6CaOxJlNytxKUBYytucdV41k4U79LYODEF9EZJRQhjivj
Ongm9sLdt8Ci6jGIxkaorDCD45rEbtt9McGDWIH6ItoRjIcC8MNtXwWPWY++ui25MKhODfc65P8b
9PsJWzPl7lNvL3IQpsA0p8YYr632n2DVN4xQL3gP8o//oojGmzWiwkb8nmhpnVsKKO7SpkvJQErK
hVmCdjA72Uc84TX0Yjtv/dIgE69h35w/2d2uELnfAmaeiPqP+JIGkfXK94XPiEaVRh/0E4izEfX6
4OriaQ99c8KtgzKwBDg7eOQ3ABm+9bHatKnpi2S89kLT0cvWtm4+zeGAaPu2TemRBoDjNS735Ko6
s4eKA5xn7IvxRye4gYtwiYFzq/I6sTK3OtyXRI6GtaDbgorNrweqqXwwdv9p37o7AojbNI5ddnpa
tJpDK6ecpMeSG8YPAyet75gpNHIUb6AOtsth/79TvoZ02p7NA8p8YhueAM4sRXTs3Iqnz8DzM0M5
Yt/ftEliSmDGltQjGNA+2oPKU5HbubSyIWWHchFBqqZg/1UPMIaarDN/bpGLC3jOQtVtV6AmAUv4
0K01FxvmHLQ0YnfRmCv7HlxJ1d+oqHwvfzKegh137XRNrnaS/nXK0T341x6azVaVfrQZSq0p3maz
hK5Ft1fkY+QoMr8GL5gn3TD7z8c5FzjVxDgeJWc/obO1bO7Es1OQlkiz2OueSJr8PVQju9Cjak05
YbviETlCBTNfmvs9nqxmcCWKAvXCmdmq0NJGgWG2wfMAjFnF2QsEikFKTrFxzTKn+ySbgIb4ysTr
1h5vgfYsdHwXGKntzy6NEDRnMo/S+Hhvis5fpcTxzYVzFI8XoOuQxdursmZvW4fhV6xkg/dekAox
EObHOquW1CkkRvEWrpXpiKOVG/wTE4rlBD0rmbwN437C5+eS5Q5dxF/xs3zJWJAeHBCdt1/NQ8gS
Ky4yaZ43jy/5UhCjYs09aK9/niSCy3qbKpD3R9sSR2KMVVVuAipbFwwc/HEXl2QbTXf9mDF1TZTh
LSOuZ0Siu2+SV1UrjaaTMeX2RFq9fAxDfzgXnuuyMtf6WhzURF+02raINHj7IB3D7aqRSgWrqk9J
7PT3jZc0qJsgGVkU+x5HcOAvQqP+/loSSyECoaQtmmFjocXmqWFoKKhNJFTPvqeCpVOCrfs+5wm9
wZ/xHyCH4FVwu3G+aI/EPbcijyoxtNW3A64m/ygHLlHnQ4Bb1UGs635AeSOA0fhC8Wo84SEHnTP5
ktr8ZQqkzzYptNdYKtArH8hGPk0SfPmlkTui6vZ6ykltTw7JmWDr0lpmUKr9SN7ecPsTfL8rQHYF
WOSbTRZr4agdGjj8abgvyy5oLMqsVNtSiYIEyFwaPLUy2gMK8ei8CQQmlyEQmfit9F0YZ9kgL12m
/4Z743P8CM0jK11Lx2fJ4c1rlFWAnnon/qghlQHE8yoV9r32Ob1DfgjTTtBcgHPCboIqCYTUClon
7W13xnf+VOUAPkJOV4CStBYBhlArz9c/wfrV9F03x7u3oRHm6999m81kfPc40Yqh/TSsbKv4qquB
HX8XndhN+iO9YxvO3xZJFDnUeYtCcbKYvX2IhJkCh/DLcuBblnb0eIukW2om5QNBjssfcfn6akJ8
OjbKcIeH6RkGs6BzVJd6qjjVdfQpeZcjvRxZxln+Z2bgQPxH2EJt+fc73B/Nu2gOFRlHiJ2OMNpV
14qWLllSMV/08TJTyIwIuhtCeNSifYd5jqdsIykVrYj5JDNF5nBsP0PrDKUubAOmKMsCxQoYy8sH
0Mrjw9El9jAogPW6eJr9+CU1K9IVmnH6mL0KXL/s4OnSGO2AlFxihzMhlt74WHTug+PZQbf9+xXM
u+DG0dI/PYE4fDlafgGAHkShYoAcyiX4bAQzZcvK97JBWfOWQGZ0g/jlQqdmadQoHrSzHnMCd3JK
PeOzC2Y5NtQLBVXwFOBkF+jl7fRPDNPt4zhHc3qFHPvWFMPDXBkUfXdiQh2RdCTfb1fqF0PCxdSg
jXv+yun/ISvu1/Upx1mT5A0eDgolxCa9Ssc5WNm6IXv0caiKiQUFqlcmXInk1eg00N5Msf9yTa1P
9WTMyAsYjr43y4sAZW9JVwazleP1JUgebRG8RgzG6MfOavvRlacf1ZQDqRpsR/j10V+a9l0dj4y4
aopfCZC3GvsE/qaaalB6v8yMSljLfXcIAFIowGoMHI5oCsOBwbHF7P58ovvc1MDyiTP+XEkJuKlq
7RKTmye/hFeL6x7ZQxHYQvPntwxM+WrU4KdIFgdEnw7TU7sN7O8sOwsiu+PCi5yelSNLTNiXD1mm
3udB1hBlZLvfrLORudBIQzJ+IcpXWdrzsDJdG8XYI+grGJSatP9gHMyZEl59gyU2bVJF8YtdpwoD
kIx1VQTNglQA2ueTDS7/HfHs25eBoV3Vt5EVYjDqf705o1FzmgVjChsT6O6yVFTIwL7lpDEOW8Mj
K5oqq9342VHGXVz5nXuWDU7YN9rP0CkN+7u0FKWRC7kug6uKlFV0GFfai1+iGtag2709ADzZ/ZBl
4fHbYFR0EhY6ZOvoRtnaejedqhGLbx3lqJVL8VKkDIT8iMjMAHsG1dy7v49id2TZaQZXPABstitM
F3CxtxeOgAPgg3qXTEYGM1jG9Q/+yDUltGsMeJEhK+ESd5Qtg0/T+lrykCoj2pmIYYTD5YCkR8ma
U74rufXW6TNAfKLnyyS6APsdSewFv5TxfeBe11rCxRF99COzSqmeFsnzB8koBxGLlihFe38BqUDU
wyNz1UPR8HV7FeCJ401gcMJHCXXd8V8y5NEn12eWogs7OUcGhRe63qFbk4JOhRnX1hXoDYidVO0p
39AoB4mbrR0AvltQDWziZZHFyUXkRGI+98p5Hfr9JnOjxa97aGDBJerdTXJ7kdkrafPXQp4m0DR3
SFOAUmApSp6DKMaTAKpin9pCkBiURkzdd1pF+RgVyeZ0desv4C3hUcKVmOfD3BiZjuqzGTWHiLDc
tsIZqDAtgUNxelPmYy3r96x+OaCAR0apnURWciXjnRFPjEFWE9lRaPC1LYaOsWQAP2AkOv3DfAhb
wwzxmmEclipXBGEnyiZxZnu11ipxsl5y4tt50OoR59MvWVN/5Sddr67t3ZptacSGVFmyPf+b4MHt
ZgBGAfqYsLq2hY5m4qLDUhAA3jHo+V5CQU0FhPpGDnQpzf8BfEU8vejRPxGeHn6KBXZRJJghqhvp
Jkb1QSB2IoO/SD7FivgXk6G5Hn0DvouvJDya5cIH9Q8AgohRHiWiuIcEoC5Tx02y207R331LMW1v
h3NVBkMTVbG8Gr+jdTUoiVyBSWl3BgVIM4e2j9nkp/iDRCtaZAu6/LoiGHUHNi2tizqNztQ6COkM
nCPoACQ9aXI/jdrfBdycsFWxseXGAWSBZpdBOyIQBxw8J/Wzx42WOP1dwNbWYpZsJXuNvWFDZcLg
eTzyWty8IvGKb+avNYbWR2BBCKgtWDbPP2eXolOdBzV6DtG/BdXYsukVKsanyjn8VS/t6ty78DH6
8rkO5MmHNiABbKMXOobfZ6Nj2Z0yzB3nR1WBGXdM6/aIk+om9Ml6lergWW1stcf/Gg8c9fMdzk9r
Rcc8L3QnQQx73C964VLq0VeWbHpX0yvjsGly6W8bG1HbV9gW6DQQikxYXvi0S1+SvVdadg36wAUw
E5OGb9FkFgeQrlN1DklyReczpmFrHYitPuRT9MrX62aFS9j2EMvi486wrnC/hbCFpc3Pbt1YFZ3f
SVNXfEr8WIDZ0qlrl4OdxOrhk1fckR/j3de3iwpEN3P4d5EniIvmwHGRiNadEt3aiGl7hNO8Bh9i
MM5rMq7k6jm3C1dJ3x8yOoLHSFHE3TpX6YvUl7/Vlo1hhKMHlwas81cNOlpu0tTapJ8uTxJr6Azt
dFD2jTMAqnTy8Ym5bo+qRKTy6PyzGQmf5Zd6z+BJ6t2uFmN1Mmo+UaNPUCJ0XQZZKnIwjSZ5h/h0
mOujv7YjKE4FIPU+2JB+nEn2Dlhwp8QJiJJfQZ7aGT6AEGuZ0n5b6Q+ZIta3ZbjyX1DyP/Y2bYmt
8SpMElbde+2wfxyrChANC0CZReHIXs5SF1EMQlIngokGVDqRB2ctekfNWs4frtBJfF7vXKh7HD5X
8N9TcOUEHiId+gmFTqH9AvXvpc0e5a1eCOan6vkK0nzCoDG4+sQMWRkbbRGNixQfrWJW/fb7RxVa
5oLQym0cyVShbD2ikPEXr/qsRwb5O/tn9E22HlA/vWq9ETbCWqGxFYv6SbC8//nMo9ti2gayROZo
GdKD5nWWvDmvZ3cuwtvFdCmcaMIohG+cBRWo8NVx3i+1wftqR5jpV8B8En1ORBkjlYoxTtb0yhqi
xtdvTGec4Ckr0184LHf3kdzZJmBlgxF3NcwaCqGxZJ7rKzzU20IqnyrQ5iKekrjXK1u1KzpfKfLQ
zU49BdgB/soUdNjIIyAyBHud3i8mV+ANyEUcUwOD40p3rhUR2GTtvGg0c2oYcF5qoqjzsKhGo0Lr
AnHyxY0ze80UEnGpGMm+PYha2NI1mdrZEOisGXpp8vqurR7qLpwF2ZdLM36XRN/RG6j6Ly6a/ABw
O/7QjIY3uJRmrMGg7l4BKwlH6M8XOc+EHDL8q7TMx+FRwKlxSbfConmy2IIqTC0WHlsPw8rF5TTH
tLnp9d2cVu0FnKzHQLupTNPF9pxGpiEt6g2cjSfTS/ptvAWf54iuVL0FIlTHXE8BTG0C4bnLjs6X
U5SZ1gD/tp1DkYvPB0VKfcNpkG5/fzbKGn268zW5soWV2HxEe6r/hCKiJsaj2z5O0NDUCpBQSLEo
/VEMzK8hzApvSOs6xxf6J4dRPygwcw8NU1ksAsjhB0/7suwmT+UHl7pH7Z8LA5l5+fJExwmKoADb
kzR3rIJNZmtOABM/SqjwEytjROM3QpuNedHDnGuN7dQxvhUJwv20p3i63hhzy8oibYqPysX/Wim8
IfwyKK0CvNLy2M774VP4VRISnOvdp/jXu91aLD2RNCUnTKvkzqkmE7n64AeOhfuJFyyhQNFSdl5h
T1q2H+swQS2bWxXOtfPJ86SfbuSjHk0JAn8D8/hIPrDtaDQgQGozKW2cs3PIF4n/nQQ7uxdYBBtI
yZjBZ+2HMNi2/VDzJbNcznVUIpflSiYrcb+fNQIaaSZEBApGhxEygwfQYf5XcUhsKSGLNzI24sz+
PRniGUMf8OqO4f+wPiB7Mgje/8p8KDNEIxga4mJdSkdLKgPh8q/+5fqz9yz+9qma30OD/fBm+Eni
NBR7ON2YpTBYcfA590bqD3gCTdW04AYRiaEEQmWrgNI6SbTc8B6CS6KQpMs4nCNpYzMAhcILRrJm
UU1cghYpL9/RFa4y1ZIqh4Xep9K1VHGarJ89kTAMh9jBQ9xEhAoe+X3cabbkDMNkM+XNyoXWti7Z
BPw+lyO03GnYnUZwkqDMOAAqYVALwJxytXBxhztQ5smBDSrZNaRqjj2zMR4TCvOo0UzcMlYroXP7
fsuAeXfWOUsM308+8ZdbqjjNz0RNSTyHJXPleUoVLi2XDC52d99RBbBVUbDbL93by2bw2maNi3/u
1cqqeQaVm3cN78THAy/tLYxpZiM+0zZO+bGnv9X6jn2Um1Q1T9DeiknHPq54C/YA7dyitsqCpJa6
UEXbepxx74ax5F4Mo/CbTcdn2hJG+MsmGTU+BshJr+R+kKhJ7OIxlbeUp3dP0m4LWjxduFrJmYsz
1VgkfPQ3VVulP+5QvyeTO9KBt3LbA9gJaLMGHbaqtuV4yON+EoRhDOgdvmfrdx1MFL3Bw1ZDE09b
X3eURIrV3+efCOGacI/BMtPL+YpXvnckx3/cDKg+/EB8Hnni+34814PpnD8EScGkr102/8wVVU3j
nIF1iKNDXiFKCSkrbwANo3q9btadwBjcy1nq74EE1t3OVc4uJo0Yfg/KVzYHeo9iC10lGzuXfjMk
Xx/nlqg8B3PKW7zkZMJo6o4JgLoWue2Ky3YLu0DBkL9tqis++HozGU7Pi83B6QffMn5MsTIziHU8
tVqU7oqzm2/4vbm476j1RZAYqSRDgJ1TSABJ7v6Ash8XMzgllo6VS4TVIv5g8FBZLKvkCtsJBNp1
KYhhzgKK725WWT95O6Wsm6IET7JXtLYTU9F64evfTbtr5uj7Y88TLrYQ/CVhFd0mm/TOOVsooIF1
u2LIijf8qXpZ+XWOWbQnn0+bD6UScDTVfTszU/Ri3otjqu/6+YXgKJ2mRTl2sHI2qt96VHt0eFwQ
tP9sa9wfSgIG5B/Qwfs0PSKbC1+nbxwfeUPkBNeC7Uur9+nwawl1oBg9myTd8yLFzEl+qux6VcB3
EhJqBa3Aj3u9J97r/ceWk0Jerl49nPNpYKY16ZJ/bndVtkly3Xyzg733kervx2r7524lxcqefKVv
6Y3iEkBzXwakfUNG6GB9wig+I3J5yRrfN+onrtMbe6IQCP9qjFS+g1OU/hN9DS6XAUPTZWdpuZaE
dBr4u+Sgxxxe31p2GtGTcg3Fiz4mdwbaQ2++ZE7Rxn9zWLuYx3VyHO+ZCvwbWaLNe93M8r8zlzrC
ocK/z5Ch4WXk0P/kl7E8YCe5e9kig2fZirPdAzLooPCKMAFHJoORTWDwOU3U+H+01Y94rn1zVqqt
3KMWkGGCQbTlSLn3BSkd500EzEHsch4Kwjn/JONbHfCNdWaGR//WKvgJbdp++wE0mSOQsvYoML5R
UZRlXQLRHpbvIFILgn0a6b0NYuzh7qSwnYzc9taYL/54E1Y5CqTTkpXuCM5Q/usFAQg0fVG4RisN
26MZlhGCpPi5keTnh5Hhh/gcukn2dDI+K7uD8iTI6KtHybVaC62hHNHzdxwM6JAjl7cnH5/6RBrK
6+HpIu0G5uqwV1GlY36pj8XCe8U0Stk7ZTr+qL1IKkoiFXrEH9WmG/2R62WsqZQADlnNmr2417B0
tp2oKzCAhnrFN6tg6zwdvFIfB4Vo/3N8fdu2vyXSrNupCCDyCtWXlXLiXlwQM82stP0+2OQMHEG9
f4268ek74BWEt4MCiX4m3roODHm+9kFmR1Qh29T2ioa15RsnXXTjtFokDjvP69xWwYVjBg7WRLMQ
CiNT1+jRm8Kkp7M9J3e3pAda+lflzNDQljAXrzm374jLryNLR4qOOCAmJ6E+p1Q1EMYA8avN4qvp
qZ488ekwkWeZsZDUWrCfGSaVVR3xizTUtluebu9j5asIyr/LXDdoMgK/LT/zysvSOAugr9gKNqLm
FsuwxQeF2RSX8hxEshfnuaVB9uJI4sDmU3CZ0W5Xyg534EhW46Iswk0saVXPSfTcXbg26zqDX/l3
jc1kuZyitG69IYVNP7rf2J+ouoUurD66pliwd0van+8T8vhKQGPZrUPJ4aPWsf9KGYFGXN2ZwT/2
DtakzmqV+WoOZUFOY3pdIxNeUU3HYs7yXz1kawyIsGFQMF35bq1tjrpXdQOseGlBiZlFJhh9V0D5
318mizG2RdXm4WXdj+WqbLbze352bJajxeFoATs1GtdoMJTUF/BUzXDnq8aHQPoHzupJ34pmCzFe
gAJcwD8L66+hQ8F7X0SAox90xsDgWF8IfI6glADL8qm8nROCpWrXdOKdagQymdoyJB5erd1kvaTZ
hyjtM9UI4ZYdEOTyHoQBVK8FJHFvcB4tIolbc+HzGCs04cKfMcWGJ8rVwokG/nlnaKuuNx2TuY9m
iVDxEZepSapqdDoJ1BEDvl2wOMWMrtH8MS/l5yxOD3XnIZ52ec7MXmeMtgcnfxAk8220MrA88V+Q
CYwM1/h7mBGzaCQUNPJj7oUqJZZeL7D39JHs/BOeHFEi/TQPtdFMzaQ7756I0qG+Pfqvx+B4FJK+
BRLFvvV64PBsKwFTACGwbHTJfrJhNUZEnyDYSeA3KOXoABbwOzeTEjdce8DJw8actgbmdUvtcLyE
U/oXhtyENheZLfkssXURKLpEjmwb8DSxdDik5CYwXkUXKper+YI+v+dcYJMgiNVFyMZUM1UlLeiK
zR9aoW45XXX+AHNMFQDQSXb3W4CL6lMzGNWcUKruGRzUqDFSfX15SR6KAIE7gFnjdhGXEPDAUxuH
2r3/nKa+M0reH8UH9INovyQwLm2dx/gabRDveqvZNUS18gZU+0MKHCH3bAiCzZzZyV64rTXhQ0CT
auNcymtKgwTFHMq/me7JIEm/G9ARFdDVnONXuYaApLbXTHCCSOiuVWs1ERdDPJT9w6NMefzPfKvv
MNy4nNevRxTUwWypT7/Ib1O0V1ABQfQf6gfqbbrwpzcgc1o+UgeMDjW9zQKlTZKUs5BGwMzx9aEV
HbYZ/GWgBF638qH+EJVzERhvJdrAzadx9wtLJiBKNTi2EakxTZTMUU7sc4ay/jkIZOgnZZSnWtOm
yYzFdHD5yTv7nsj2q2/faGfNhuHHaMBFoHBAVJ0WPBDNyshHjIKxFn85tS1flz2+OrvLs6mBd7UG
4RK6Cik2aOMaSaXIeIWYfyi6SzIGyx4bOx8rXkMU+q5mNIHbf9/JaGJ41qdceTv13l8VMtZxIF7o
aubapt1TYZSv7W8mIh+op0AClqq5AapYqAxN9FOorYDwUUuODd6IBiR4NLa44lOOtdeMJwbR1EDc
2tPcwiQDD9JxUTLTkk4mUR+hfFtNy8hL4yc1L126KstV335omIpD8bw2kFbeNRPx0K0Zbfnd6XHW
Vj0lUemIQkMnVmppe8b+Yh3CUetiQNWRZzS7s58VJSPMQqmq0hrpet53PZTDAuVc/1Z+BOtbH80X
mi5zUasWnJakbi6BgG2TSkBVOjACl0pxNHUNkESQas2nS7PEZYIUcsagMDGewPOGr1CnAaXu0FCc
PKhrGqGW4B3gcmk0nxzS3LMWZ6HfQVRjfvi2gTjCxCDM8XjUouvHvIQKSGQCSsTaAOnBcUbpHFxP
QbwWlX/IwUkMEEPSkwIq9nDYPCsptgJTaWwvVCFUKOXKAibALgwC9a4J0GL9um2xVIzi0OEX0Mwv
ptPr4YPUovcArx7VGKk2sOGX6w4e2VFAuW5m7GgBX3MdNSBJ9s37nuOBclnHS7A/GLIc0ryappkC
xekPBBD8p8qhWesynUG2xvhhtT7PyBxFKPptqQFjZHoZmC1zrsGJtmfUJbST+MAI9qALA9PaPTkh
LGDGr8GOCz+Nzgyxg8hpLod/58DgNvwGeBV7dsaUxZVOz6HG0VA8ZqsREoRBEIM25BvFR7B1KTP/
3KS8pqgZcHp5zyZXipLUK0MBmJ438HR9Kf7hwzi6ZBHVykp6Uv/q0rv7ZJMKDLeOJIau0LAe3v6p
sOt85dqDRV8jxeCqbSvl32qVTx9LcQ+EGRHTZiUbAoRXoRrj8Sn9SJqgITrVCwsGAquNAoYkX54I
tej2aOL/+YoPY4EP+apodsfm+plonl0XyhwECArZOyUdQ6d0r3PsTPJj/6OzvQ1EcJpGZgEVrDa6
/lx6ble9ACa0G0vG+rvB2WqyjCo6lFNQWDCsRzO2h/thVonwW0YxE6ZrgoXiJOque/6ivABVaxOB
jIRxVghnekLMu6pqMfn9cex30syAlmyBSxEuzasnaMDZ7xpyjqS1NXJzIDWskB0l3PRXfWZMy789
A27lTJoBpPxRFv4ylhrdkl6jbXc4nGiSKpEAqlme+Br7vmrrb+ie2hUrQk1QqXHqw8TI/W8ySIZg
Wk9ciDqbVZduMA9WzaKOR49h6ZMuNEgczgAG9j/2hf0seB6/pGS5S+NZzXOh5qgByscwA7/8d9Kc
Bf3WJ7IDStGADJTlaIqW9DXUWKVotFNuwIg4Hh42OlzmCJpX7axbmehoa9iLQ5PfJ02Nn2rEsmG2
BAImQeosso8ewDTexQJyhWiHNkC7YUuHb0Y5AOQ7un+NOM+Ns+HjwXmpvGb1AoqUQvccaixDeL/k
pPn/VRJCCZ6KI2H6BFeIXAhAJ64vziIBi4lfYon4bKFblmleduXxhoLsJOQPBKe7T4OgAtJx06d9
XYoq3vi/tsX6v+Rq5jEAVSxiKxcZneY448qeWT6MV4bMRVwZqk7cXpBo80LHgx2xKOdakCPlgrGo
xBP20I18eQQajeKcwCDerPNxs4uyHaBonRZlcQToT1X5RlNMKswetST4MCikTRFg6iMhSR4JwNA1
I69bAHeZ9MdxtFiplVvMRADzsBqQQFH+bFdEJhyML/5fTtqh2aj2UA9csyjvqtUbTmnFjJHO05ZJ
Hvohbwxvhw9exNAABoGLKyQ6DrNxKPnAEZ9WX20sVLuqJuGoWXFQt1Myai2IYbryem4WjH8QgztB
trM8DiGDTQAMXzo+r+FkNZMawG/UPc+bVXb7Rrmd7+oWroRBh2eKBzx4gKowg2LfZZrjkUtCQbED
7KMSZxNeNPAfo9B0tyWWorP16lfjMTHjKTzuwEgMjH8yFPTMx1EWp0FQB7f6LEIIvu6wnEe19NB8
9fYKqn/rgCykV4mdXgmV+7CzAtg9vKHWuEnjsAIXP1bET1qKhBIRRtvMeJyvlUO6Yddaenb5dvIs
HmgQe2hsbGXtu8c6B7jBBeI72LFmmxkKXSomt5LYMWdYHW/0ehCUoImpzlo4yGmCof2lwdrzb75F
hqKjYC1r5roB1sp1VlKN+9b4eomWQkdOu0rijfwfF3a2kdwP8xRImBPf4X6IxcMKMuFJ/LkSRTzV
bLf8L2H9YfhLWDVMCdcZ9Pna8DemhfsXkVvdR3s24uHzT3bSOS6cfCCHZ23ML2Cy18RQKmKYCeKJ
EjMQcBPsw8sndg12oXcw4qeHD6dtB+0rFAZsQSlozMnxEYym4W2dvH+Kcw+8nZMQTyHG4PHqE6a3
MGIkEfaXIiB0UM4nd0C+rUwhM9hq9uYz9cRwmDPYoQngy09GySc9pH435ofWSUc1Y3oaNs3hByPD
2GnWIh00xB4Bgc+jDVP2b20PU5stwYMtUjX5Ydh0uoM2ekTI6tP++XXpjgZaLjHMBxvQSmG9olWP
GZ3mTpl6NwbA5Cuw/hJKLKowz+eVTEtUGiCCOcsLKec71Aqa0yqCmusNeAFtOX1dOALyXaGg5cwF
JAR3DmWMju6Si0C7X3NGLuZ9V/Qx9jxehqZaEX78t2dszT+HDaWWPTBsFFB6O6xQUpvqOxUcg23s
Ishhh1dXzY7prlqQX57VB3zGDygn2zOioLajOPcwoPWyJIu/B05dp90FmgbhezP2Pee3HwX18KIW
jJi9uOCaubHdKVjm44i0YmtcJhzzvMFnwmraaN4OpiDfcPH/qCfMqcTI5pe3W6zkozQKnarR4HCY
+5/eBPvrPs0seWmAg+dt9EIiMDFkmH0uxUfmPBPFb3aVFpR9+nK/dVxp44AwtLlkjB+/CRvYrSYQ
xCsPGA0MDfuRWl6XlxoZzmUHQk+EKi2BOtP6+P7JLTFjMZ7ZL6KO/Qcj43c5XjguLRIvd0jgmtwu
nRhrVW58Xt6FZq87x1VW4N7rDAp7to1ZobETBCPQwaDdj1H3BrQg8uPxkrKT5HkvX31bVq92EhnC
DLjvU2yj3j0RVW8tkLzrrsFTb8ZkG0HOprIL5veZt8VvAp/PEjIxLyPGJu4HqesNm7SRydsz8WgB
RFPJ7xx0le0pAeY7ffCwMM8tWFNQkhPdfOWoSVu/Ye7+5eIE2R6CVu3a2k2CObOTdeOzmRLsoeLO
x/YXSvr/xMDqtvOZeMra5uTu1q2dbty4aHx8kY9ImBuSmN59dVpgXR7E72rYlJKk5oDg77VfzE7o
ql4BHiW+Uf/c6iazrenFfrSFfhmh47sLnkh+T2+ed5oItMPa7DCSR6xiikFzoPdxPskYpWUx5GaL
By9ZwduqRFoLcr+LCh8O2ZjMnuXE2eY20w9YxdCh8uLXJDeqqv1CSmTfY/8qjR1eGn/w+lJdp4gh
iYRGRkjwSoBX42Wf/RKDFLJeXFU7QwVwwgCWVq6xjw2oxIZDh0z3oU6v9EIcrsU+3EbHsFzZdWSO
RuufoJvwBMtJQY+h8FO1jn4X8YinAByBwrIyJEbQctyEjMv46nXayHpjFE2lnOEQFJNQHz5K8LcW
DhqcjMdxMSxVcEqze50o0ScTOZutrQ6aIyS04y68XQpaarOJhczhScAkGkd+uHYTPThYTG6Q9m0q
SvpvxN0Xa2eeY5GD3rw+Vlite/SIqY7eoqx9ZjsRrZXqjM0kTgS487rPu+t2zMQrLFQJVfiyNV3L
N0EwbzX5cgdfA5gSy90ffa6FRQ1WXOTcrsW1zn+Hxx8xjes9VwS3OdhvotaWlpEnotC9JKRBUs7c
mFvnjLRxv88lHRTV85rQM2GdHSxjkrztdrYDmWGtz5H+wWSmafKCpv6WlvYPBYuf7GXGJzd9ZkYZ
EVN0BKM+pWO4FpWJVfnF0+aSoIm50kWS8yjPPfulx9UXGDM/5Bu8wKGj3XIBODU99QSFUKavI46s
JM5V/OcfPCBh9c1IxX9NrSHRu6lTkCSeFGHbi9wLq48Qx3Xukt5J+CpIRVdp+2+XtC+S85P5uH6H
dWxZI9VSmn1azS2ppBn8rVgPRY5IXiSBcHh/NfeS+jwLGVvPsWNbri6kGY4hCR0cv5idlb+cdcLR
qWRIfDiqWEgejqfkKRkw2Xj2EOUUJNBPVszNTQt2qFYk/petwm5uaEr3CKHM09lUZ+csqrJseLf0
uASWobVl9n1cbVaE1ujbeVf1rLhdD+wdbE5Wy8WV6ZSgQ4MdFN+5UY/NIlJwTnD4oFXGSpj8hMGq
YPqNosup0BysC/r/6ZYIzvIiKZ8htc+9P/VRn2+LMl6SwMIock6VH6BGhb0HFoe7w7LaPaNWzJr6
BvNe20UW2DfzZcHvOE0bqbJxVhjXoKpWvMWSErEaoIZsFT1ml2gElijNFUrA/3JB181XNmGxAWi4
r6JjmnMkMwaca/hjhNv8hAaH5biI8uyV1b+k90gs7KSLKQi2jteDFy9F53b07VexBS+TRc/gmh/O
l3BfsDWTiw5GYmEhgFXjaGCDNzf+hIyblkpOcMK1S3x//vVskFx9lbtd2fO222WjIwy8rmk7MlY4
r/kbQMRdbydySYPKRQ+yKL+OR7nvvZfTYhmUi0/Ig1kVrRe8uKIEEcidCbdvNv+gji3qxBJuOZzu
f6eDeHjeASeNsM8KgH0XXyb49OqR02TJo462MAQPBdOdBdjxEJ2uKeRvh2nXa3Hc5GCUF6M861YE
nHQHuBKTDVypnrbY2BKMECny7OmH+wcnym1aoB4vvJiP/Uz3jONbPpPV+VRkMzDsDK+ZZ83ZqSBc
cvp2z6JdHfMY8XgsczAzwyrwBHQfYyQs9Zo2CZfyRvXvATaN1Dyzl3ESbNQ99ifFxF2mNK1fBIhA
0rKdMZT+gb2RW2lk1xU5xar73/OsJ2T1HpVFIbz9FVPX5uK1BdIsat7CqKstCwmCxwpg+dbWCfx4
amllvlF2kTY5IZVYtsgWExN7u7HJX48m4cFULL0HTzBXzm63C40YMPZDAE9ToyqHw0+zfCruheuU
4gT4YWBCXbvxXG9Vql+PXOgkfIhRpyyoAkTYkXY8pA8HShlnRfzR1fyaFUQd5/CmCMyjQIp92+Fm
kTKiVDntXigosQu528kwcRpb7gBZmK6aNMcyY46IUCh80/lapmBy0444pPKicJa86O84RT8/48/f
dcVTLnDzpttDz1RSJjEqIYxi8VQT9ll2fU5BZlsp7Tam92l5cGzgD+pPflep/4OUZ27/jQfiyNvV
wLVk5ncvmywaS32LArLHcumgPQtOGjteGZi7IhdkRTqQqNfYd2kpxxVunhKNc6HKxBQlwkq0X1zz
cgEZ4igXFlusPGLNhR7ymt6zrWfcPsVmw/5NuV5EI3QDB2NeF9R2znA5TKOOOunzIb7pvSmdESfT
b5+87NnXGuJSF+n4TKKF9GQ6L05nje8iZtxgIXytaZWl22ywv3wOwAqnwN75l63gu0X28hlw1c/K
XnD3vqFg2xgGqA2bdVv7qcX1aZV9atG7UXIkLHqwDnQ5Vr5ckxevEe1Wg2ql1rThUKp+OoSohkYK
0Sh7ttfjY6SNRljF+X+pxiNEuaUuXpiSiAvz97wA2T4oMmKfUAN3zWVaQhT+FqIm9VGyOFIXYMfY
Vy+XJ7Gj/MmG3ShTUFIrTM94J26Wriw/Dflpb6yYw/j+16kW0ZVVICAFnGtSpegmJo1vRqn/Lp1u
aqG2IZAqs/CvmB7gpHnfePlRJf0HJq5kAjBLEg7bDMhjc0H58sxfUsuGC3BzJNwBiieINOzlI76/
9UO7FBE1gKhF3rdfQ+DVcnj8AGdgervU5apeW0KoCz5BKsW+nVqETv8bITx13O44NDUqhI+u/0nu
gK3pKphLG/ZB9aEJk7Bz7YEtqz7VcESmZNhaaQ/w71Rk7lI3+Tfo3MkLds5YNMZ0NYzH/uKlrUKP
oP8Hx0TMAMEM+v4QNn8K82FpOoSafuNOQFE+JPJf+9bxkIn8sMbIO5GJg6U9HWzjjoLYe3XC+ork
D1jGXhZABMRL6Vqbw6ZUTMyB4sgF1esB9BNTeANqX9znZdRwuzPIk0W3E+uKN+7uh/E/X25yaQvB
1CPhdbLF8zsZaj9Xg20YJ4HCPlF3F7HHXr5DMoGw1jafos5KqNAEUOupnjjngWN0tq3RPn3KVQJ6
jTRSEs7csfKpBGvdFmwLAMIiJra0Pwiu6Q/kD3eKiREY14PTNrEa6CX9hMpKDqqGJ1rFLbg4vLET
86mM9GKk+KQ8t3g+5wTi2kXjU01mBpKb0YGKUFydVbYdbWfI9PIUA0dLBmg3NHLclSSY1j1nq7Do
go5R0Qs5Lm+GbfMaRZXzF7GUNdGDrmBRb+1bolv5OwjbJ0zdbA/put+n0OICLaZKmKLTs9Ht9Whe
XLwYqXncYbd2NYuFoXJG4LjgIvUhZf3YcWbXi9H0NW1Pb9/EUySYZD3uJwsJS/2l61jT1mXL1lZm
n01rEArrmifS+mjYKG9+zRqmKm3w/KzLAEuem60a+Pgcr77twapmHGdowv9q+P5TvRFNTghVamxl
FCVM6Mx6x6E1qUOj0ihQkbkSU1vsUNLgg5dp1MYkjgy+d4ocWe/wMK9MbjKHAg1L/a86WVkGMFz1
icV8T6TAYdN3nBPEaps1ngP2tspGHYk0RZFcGcM0yuHSpOLsnqaZfNXSi89o11d+ZdEO1kvwB1DE
PILk6yroxSBDE7z/YyPBNvqkXz/6SMUB0MmyrObKieMGDGfP7xZAEPtY6UoPICuxYlzgRoVhniIb
U8w0aiOtiKxOuxPsZtr7kVP0PoXBEEYG0Fz27plLhjLCGwVNXfdNbEzCBYGcmMfgTRcyy9FfOdTR
Oc+JYR+9A+IJPeycXyTdEosrovfu6uhgdDNS6vXh29puECRZ6MkTS4Qc+VHzWBNQJjzP58sqe+U6
fzKDgsOLrdLF4D/t1/71j0LyhpYu+d7oqNifbpXJ+ksbN5I2zrtWRKA5MpeyZ/f4r7QRCFEVy2DZ
rJd9tQMN+HAUut9FC/h5bVxQE9LX7BNqTIppGKtipJNHOW9dfuePbAffdGx+vjvFb3Yx9TAjx0Bj
ev8y1F9qH7XSJEhBFfYbbWIXoup2kjdOtGTgAaQUZ+wRzWgXITvS0HJBLELS3eUF0NCj2sZ4s7FN
q151fu0kNctszmwarEfMtghm40j4Ls/+lautQr+vUZnP3W8zpt+MAMMgzhrpO/92tqkE606ryX+G
p6WR6fiKQ81a1nI3sHCAq4Zv10MV9RQZgY40Na3a2I9qp8Gu8ULyo8STD0HvzEJjRVioH0BNegzS
YgzhrglzBxXaEkF6auUxtVmtossgyHtsVQFg32JHWd6pwY4MUDidzhXJAjkcgy00wu+39kG0j4QD
/M45MuwxHiP5gAUADibG0erefJe+NGT0pRNC7tvv5fMXt/2b6tdD9DcDXGfs1JN5oR7Bqdpans+W
THV2HgusGay9BZ//Dw+sNhMZm+QPDKE/YnysZmWqQhWd+p4qD5d73+vn/Zorwz7P8uj44wB5t1HA
pXT26qmHF3H3IKAFuK3Xr5rbN74C9vsfWfzq/NRVNsDqcgvepyTF2gNjdjPn6SS+p0F2rXFbANcp
kJqgLobg5AjqBcHhagdZ3Be/zYCp/s0xMwOZMPQRt3rbbGhP9nLzTXUQGiRQ9UVSU3id85TZJfd2
o6/QavpXuEHrnCufS555aVIxauHkqCBtvfKLYaQLerDbfFVX/gNocBwaY/okf+dKZw97ncW7DEqi
BUfl4a/N/qJzQI9uA0wDU87sgPAFd8d0KG5opEfsTnKgoFgCRAaDkx9KnPcMQITDbo30y3i0GTSL
UY2CV7f2VfVTOvG6650g9LfIpzoAo/BlWsaweIz3mExKHDvsXNA0KT6D1ZS1x0owhcLqH6PExSLI
pWg1bH/wqqbEds1qK9HJA490aHs6vLce8CUTP8sx8wNZDDThCpuqBWqdyFq1mXNcJqwFIA+3pHOI
6gIm0VrFRDcXybV7fZI9UKvh6vdts3Z/OZi2+aL8+rJ9kCo5eC7pVOaLnZmajnHDpjTDZrngL4Hg
Mgiow1PEtw1D1lhmOtmN58k/4MyimGaSNeFznBkfO7LIf7fWgEY5tVERzJklt3xPX8gOZMakN3K+
bu24+SoPwDwhKwV7E/JEKUIyso2PTdwcvqEuxsaeVKxvoT18v/STfX8/zIfArjIvO0fTaMxM11JL
r1VDA6KZUOaQ2knz/K0lk0eHuyuXKCIHiQG6Top0mcBu/s1xcEHfLY5ZvLty7aYqxVh9uc/LVsKl
uNe9VM/U4lNRvavgoIasYprHKIAcumnzgoOEZIcpd9/aJpSNs8Zb7PCRNiZaFblmqRrFP9yTgedl
ujpOqIDEqwRbHJns/LXLVLUfCjiYFeZUXfQVrKuyDiFEgEoeskmd5qZ59KqeSEpoKbs5e00tmBiH
7F39QEaAAP4e9iB+Wsq8wUIHp6FaevERKM6uB26G5l0FWTYEENKOhjXJtliTAPH6XccNoRcc0WC7
F5e3YFHtC8jR+vFxQzXl4jeqdwde5LOntIoUIa/99rNhPO6DWT6yhrTpuZlSl+CPmFdHlfDLdzFm
Evsami0VsqzmbKLCdNfxHaWOgaYOxquhJd1AgsP7YGkZ2ifDRLPC2i8vYEjjgESBrwG0H4Xvhh0f
n5spcSrYTB49OacQtbJfh27UOyTkSSsmn6EvuZC3f5cjHaVkdEjbJua0Lnm61uHOawTfO68ZfYkM
X6mX+jQ9S//ut+d4oPKmjE6qonv0eOJaUIfHB6NyHDninNspTFR3r+lWhOnyIt4i+rBLyuaQNsi/
rW7mrsZiK7P/ExH3A2gImiDzGz6n1GlNzC3JwvTZ3qgoJZpwuq61Z8VfavQJIWQJ+e/H1fLK2Bj/
hdZSy005Q7PdmKr8AJexKt3m5nj5Ar+L8MRdgToJqiJRVZvkhNna5KHeQdNlc6Ym/bHiHU1CAixn
WVq2VnUZlfo7A8X+50a9QLVV6o29G/FFydLq1ippi5Du8wHLZqyzW90e4G0LNT7yscfxUsCJY/dx
UvNyqzG1UYhyflh728abtPellAsiagZamy10Q1juanTskOQNXjVi3qIvX6TNShX7CQMyA3i+A/mK
+WK++BJfXkuM0B9alUefjVW+Bz6/t5U15+CV7t5oeuCqJzgb41m4Cjw2L7KME8cAIG/a+J2nNjjX
FdEJwR11Mwh0664XOFp35c1jUE5yHPYs2E3JzbJxoUXWDBa6pHxhh4R1juiRpXJ/uBamBeFGbaTo
dh3Y8X82WMKMfRiAykQLxPE5ZIdQC5DLaK1xZZKg3F/5LHeft6+yMnvNhqUK0J/fYMHWoaJOsR43
4lMbtr0tNVjuzPHgYAo0K05hJqMK0Skx//nP56C9yeoHZUfRCFdih4qovlqiAdEEWddSqrYV/2RS
4Nu0MzaQwenEU8ST5gh0DVB5a8Bk+NKMteY3Sm6q8qdu9PjPNjc2HcfnTjluBqXRPdArkxciDspC
TlG3++HKFyxUvFFs6LPlrQrPwyFB76XnncQu40vwKW6KsO8o9J1aWcIa7LoIMoyXqLlotH4BlLfM
IgGx4CzbhpGiIiliwdKwV92OLLK71R1dOgrCv5H71HkmdRtIqLlJlE8EVcbLpdVHQb2ahF0hZEY7
z8CI1iK4nFIgYLrWyDSUQUqgC40CvSAO6NjDzE+AORhG1i4L4iUaZuenl+NDCc4JIPEeUCVMiqS5
DAlRNeWIg5G4spC/uycA8i7lBxwMCN//wIhK/0q5qdhUKBVMa8Gu+bpIBULZalbM0UT4e3bRI8z3
64+vnHpAPrup1TEQ/mYji0Xq/19xK4VI6hG8wSK3jtDE8qGHEqbeQAEHiqGNc0YOMUiGqLK4kCvY
csZJl/k8ysZs0n/9cOXnLCvEOgMUmm9IHfzIQFV886HjyNVrGoSp/QTatkgbqs24CHG0Z5xiAqUh
3tcIyUCNtEf7QseOfOxJPvZ7NaSQ3c87A5TPbUMNAdg769/jtRyz5AMNtlQQgaHocHqjx5zyacuL
B4+P2eAC23wX86JBVpqObgEHMCXDvyIyuxBUhnFFz8zHvtT6GfI283NASa+oZ9ws8UYpIQMAV/Gq
YnpNiQDJEn6Di6TSsQfqaojpwvFly0f+GVa4dNJJOEyGoO7Qxng/oD1hlwfkad2Xmocx86bNiZ/D
hree+aaw/jZY1PPUsTHyqFHzPdAqLl3Bcwb+c4O0z3T5z4qvAFWery3W0cpOJtEqzovbVqutjnQE
UnVvYMCVFebbttY+y5qItV6CA93G5GcmVX/esDb2h4Hwz8vSlr4avcXeM91j6kNfnjHDvIZ+Mn2J
xgdNafOteeUwVSa6xYevICxJ0k8Pvpu0SjWofkLUcVgRRH/LGjuQEZDhNjiovSz+5PiD0vexbmO4
uY9ZugkAg9gknnFJKKWgAd8fzrCiX/XuO4fIozKVpORptMsG8P9+CPKVZr79mW+SqF7i0zJfX6mf
oa0Djuey0MK4nD18Kng4y87gwCGyTB+UVNEnQebjbPIwgdf2k+WMm9jBPOyHE37tGiQBs53/YAXj
eXN/aFyAS9fsbRfon+syu8XzdK5GaAmmwaq8nBGrqHN21D4dEk69nVBhJKnDVkVfo7bU6m2wYH/4
LDOKOUZbu8H8S3Gnw89T1iBCexG1x6IsxIVSuE/KuFnupfbjeQODNHH7nJdbE9q2xX2tg88YLDOH
HQ2SZDTjkI0hM7BcSifjvXSDbS2R3C7UbPqodsMZSD6l4Lx7KoZ4MdnufYk/K1Fin/vRfjqGlV/a
AwlW/t92UFU/5D0hkpJhfem1SZA/efFpP2m8PumQNSRQ5pfYQBhz1/nsMyJnIfUixmbJbaAVVOlr
Fvw5vc7KTji3b9lYMvEEcU6CA4BlNHKIGQBvO0523SIpVGDwcJkryreAA5/ebxI5DaxIPIWEf3BP
gxOVEor5ZDiAqH3z2RUUajC9GOipXbjL8X6fJG0KLausWbyY07y2veE3biPJgD3QPT8IuQNUbV7K
z9coytdeOjtVxtrHsbvJXT1UmrUqEp4C8dAZC2OjWfi72qQUImv9XZoaH+ea73I4P07F0Fi/Bl5G
SgBZVnGWAOQOeFn5gMqIfWb/ujn/Ab6F3U19FtziPLbzeH9PRrP9vESowWvYuYHDAb4462lhZVow
8QqeB6cF5KCdIhCA755oXFtey/KKx8wFlarSE+0JgvzQQPfBKQeMlSRUYogmROAoMVkOH2In+VSh
yBnwrKSMZcjRqBpVX2tQJyp6ckMwUqz/CDwx77jA3dSEVbn1a/oAF376T+w/pB91odeXWzwrEyrg
YLYM7sm6OqpybPaQBvJfYBxUgvfn82mdKlut3EkC8/DZXMXoprgG6WNoOkqTNQyjy341wqF0YmUb
JA4in37AcI4UWwSXMtkE9LBcN9MIngtz8NAJl7z/VaziFMwrYE8RH0pWsxQQPNiMLHUCzRmSg2Xf
rXfO5rVEWsYefTBB+e5fCWKb9CahmANuT1b139I0g9KwoElc7KBl1bPP11NV+G5NbRjdIZoA+ayw
7+0Nt/V8mkyENr0QfDUJncGovDPcDZCkOh26hsTkHN3S2m2IIZjY8uD4Se+HwgiYmKTlL49MDbMN
WGoUbkY5ZVvtNQmjFbBudMRW53wL1glHgWre1c0WMIvHowu2xLmoJvnTZy7QfSHafmFJdy8LkDe8
Hv2El3/Ibf7aX8aZ1kWlRp834SEDIdQC54F9+vDQIWzBaS51ZW2BV93G5Kp64ZRBHO0eNk89+g/9
2GjaHv1Uv8K5sCH0YMmNh/lmNnIij05DyWraFCFs96+URL9lSoe0mcvQa5OLoA+cwpGE4TEiL2xl
GGK+56RlKLr9gYS7i9aESD7KwUVcnGUMRexNlt6v/EWgfwVx0Ek5E01IxxEKjeS7Up+iB2uS3wj6
VChdiY442eD1V7V8A95d8liEr8Fhu9DW5YlDkv9975XcttEQiCVZ3KHmwrWP9DDJJsZvw0p10rcm
wggwq50gCqHcBgVQKamicha/CO5tnc6nJwqsyyJEOM1UoMmilc/U2gWOWC0XYdepGj3agHN1E8iv
7GMaAFG9acuaboVtuXD745kwzVSX1sDjRvD4L/7cMZFgiRM81/bL7Dlz1NnMEYLYDZninCYwyjwb
L77GFO6HuEscvbbt3vmWMX8q4p3DJY8Kl2UkMaZi4gIKkJgapQ5RLJQ53EJPU9qfhbHaHtw2yDYG
V0SG1MwjbwSoJi+OaFCjsJhmFKPJbIe81Bl9CQbb0oDAlByp4ypN7AARpgdngh1IwPDt0ywReB4a
A5lAizAFkRM4qjwuLqF4FJdY8gPWhNd4jw834EUsadGoSeHVbboLS4S6190BQxCmW9+oMfGAXtj1
e0L417yna21pYHIHULGKhYB+x8MtbGDiOLgexhVP4JbYv9vtLmWzxtOKYI7kuMLnAak6XO16ZkFz
4W64b4igJ5wdmgQ7a7FIBPO0UEfs1TsmNArhiuz+aoTGYVxanyM8NKDcq+dacDxy0wINExNGGBDC
UT4ZVu2GOQyOSGXgKqc0izTMUV8GOT4EUGMZkXbYZ2aHdCEd53a+Z3FYlQm69i/SHOSocKSVxMD3
2fvGx/vqJKmGzuERGllwChEgPtCJOcz2P9P4UHlpwR3Ty/bJk6h3q18SNr1zJhOhU2lztsa8n8Mi
hnms8pmgQIueOhSrU2DbInjd9XJa/K6x7ioNwz4hghll+yJBDAoJvGtiXcz0otIrTVcKARNO0yXO
CPLw3ykvlkt7wLuQsN38lUVDiy64DIj341BoTQnh3D18PAdr5b+mOV6zciu0ubeRDE03wEqxXMkZ
ux+xrgLRG67KFLp/+CS7/1FbHE1K9lQ4YCMTGf9Rv18Q8HNi6NX/v90URAVHUagremiF9KoCeXsj
cKNvHha4W2MweHwXE8ye8tuNdDr5B1nI2o36cA5a7UYxQYShUYooie+y9OdD+KNxuy1aW4bcWcY0
YiZpgDcAR/+7CegQjxpzQ/FGiWli+LXAVuddT5GtxkW/XagH1grnXM893/qoW2g3m8ZKaCZQbdkY
DW6EA4dY9JSZsoyOYBoBLNxMxqu/o/sb3gkPPjYnxuYTnhMfSO5UsbOdeE1JO5oapW/Rr95yHfui
UzTvNj0GmIRyiH7Ek4zGTnsiTnmd35eMxp+1tQYTfX3/Jku3ioc4eUYD0Fn+i3TbNEpS3wdnRXvJ
65laVOcS06jP554jvohGfvsNBJ14ZMeNQPNMSGxJToPuED4ysKrWd4u+ohs+MWJN6Ck9+gY8fski
m++4duo5kodoHxV5DdCcBlkr9GL/SsNx/+IaDkFXDbDREfU3YHQyveZ6RKWvqRWexaSzxTxS262V
rEm9yiJvxp7Awlr+0WkyPXBwsWbVdDEhB6NuDICtMlEpTK1Oa19nX2HyUJ87INHmUcZok9LKAgcR
jmuMujSwDESGYfdRvhGIV8bEcxontDe68qFHnRrF90Cv4RUk0Jmfm7vPNUpnGCTTfnwA2A5zF0Ei
qR3XWMSPk6FIRtPuq08EhkMwRZHLm8VoIjfOddEvvqTEpvZAtGpX8dPoTeqSKq4rjgzQ5KxAumts
Vvt9GGKyg+r6XgCTK13LYA4pDCt5UCDmvxd1aZudpkqrJNC9toiBhAf1x9shQRNvCFlqCZhPS9/q
+G/Vq/Nv2Ib7LM9oTmzrmd72nUY11/3BfhgPDDMLH/yGSTalnWadTsKBxGV8S0KygILKCrS1Du+0
qgvvP/JVes6wse5yPXmJtpdZV3ofaIEhWgEBgL5fA6q0bicoUWtrdNvM/v1dvZfzRdxkUZNdOBmT
H4PDQZofqTSgPaTPP82pW92IeyYMEJvzSf6eDw+ETy3n9Is/EuLybKEl5aPJ3wFWkzKkmliGM/Dt
C3u8PT6DB/NUhVO6KkZibZIHOOMHZ2XIlmIo5hjqVPFfaCcUq9WNFTmowXzlYpNLBsHFpJcNVVRf
i6zmMJQQ54fmjCuFO4RPzD+cj7xFxcPh0QxzziVIPxB0Gf9RaXGZcfs8FQk+Hi5xmLDa2map90i6
GCQxg40SXbTwrWNpL+bqFOHG52lvHRM1d+QH3X4d8/ryBSmtQN6hhMxz88XxKKPbEAnKE9vQYzAu
RNwHe5aeWiCR9ncHVOSCeB4B1+K8rg3Sl8ertojwmzbwwCTbNVuWPv9fKgz3dXKwxLC9FKOfMAWH
H4JRxuYAcdpBYZyDpob68GY3OeOF91nKSVoeyk2n949V99sE+FIoJeEmgqiuWVuLQUBEB6rpRyxS
mT18A9YT+ZJJkFpKF/HP+3fokriHpFaF6M2C7w+NBPxdNIp7Bb15mTkpvRiVPI4NVeAoBLdcAWrg
JXLnEpucP27eL7u7YLA8RFhVTq1nrzRDmyP01IhFAC0ER9xZ0fGViMbAJ0ooPKMPVRiUeWxckIzx
bSskc3FCBMHiOH2vA3Spb95MNRSoMdcfRSxLuV77vYqybJafI6DIOmqo1mINlnRru+0U1qNsbuiK
OOWHiXFTXLzoyEcFEIMN/OU9dtNRkdN+wz8qnohWvgvnYYjOPf983pdLIJ7xY6rwRU7eon5kGuS7
BbldKTnaNNP7Fo2XGEl9S+AkaaEHev8IL9VDAXKxLCkugD0S6yajZHlbCjHknbSFzK/RnQDliqL8
vp+1PvjKxdaL6A80o8jyxLxpZ5p0H/45s+7YaypkyiMQZ1XwDBtE31XHHyER9Ufk7EJTdxxoOpNm
muwysIheOD1DmY8y5iFXusW4fzZW2v4qWevzZ2M3iQwIJxaYp1bXDqvodI6G+fdnrdsgTsbvTBLN
XIcUkrUjhpK+gdOsUOsQk9flpJAph64ClZ5ZzcYS37lgyNB2Di87R12sORn1J2nUC3oPL2/lsA8S
oBiB0Zw6ucJslR7RE07Ox/To748nWkNSCzKWOeNVynr+7rQsHn00ErHSq/S3RMAJQNOoxG1oayxE
HNR0sG0pm+F6DOUFaKv57LfcCWvWAhgwbqHRaGoWMP1uENgTF/wTuAOQ37xfw/wV7WcE65jSjnK4
eUFqdq3ywlxOKSN1BC920MGZyBWwxXkHfisagH+7yo4koEXAXzWUy5Ex+C0V9BXka5ApvwYjwbDO
RmFNhrN8LYZDqBQ++CCJGfVQc5auQ9ltTklVYN/V00VnOVSimHpKQQWD51++qHATVSwRzcmB5nA6
WILh8KTGl1JndZ/N4k2YzGJmwQc6/+UbL4b1iZZbw184lFNmiiMqE8zq/XnLEq/NRAO4o7TqNLL/
vMpn37fxLjlJXic6HbSpFHEjNu14y2npMW+zdRABx3PnJvwAUhJsmVpNR8jEt7Ff+cfX0D8buBpm
MolFb7tnWQ4fyBaSD7WT8eL4iwBOyEzRIswlCan+xspdEdoToRA+aAhw0BbVMn+z1/oUBf1P9t4Z
eIfOH6DNVLhmrZKWXLJNfv1PjnVyRWJipv6cWxBb4y7jh84QcMJNeqLJR6Gvr1cbBgsv0JQOVckU
5lE6fixvBuJFqZG26YuMlWUSzRYK7XKnDkc7ZwGVVS82jSaSdakB+8UthZUDMKD95dbieLfS4iLN
Id6NSmVjnQ5g8FrCE61z+y3ojig5eC03lA08l9xW8XX/75qJumCUZuPNnF+RbnBGr220dzxzafkL
KabFGxIV4kKdZ2vWTj3oj+oj7r98dZu+RCPCcMV3Q+0P18TPazF7vDQLliSgIswu101tI0Kb+6Gb
QFud/H6Yz3DwOM7jiK+4jlz8IQ66uCDHVSY8H6AnQYtFMsTiySho/5VoHk1wvorqQsXPpJFbakux
eWJouCgFL3sF57TJiIRfbFacQjjSj12sTejngSZl+B6fPAs8+mocZQ3pwUhNr7q4H4+Ey63Y9Ga3
ym2yPyFyg5ov8tuvVAolUUoyTHfpp6gr7c+nBN/vs1hOK5i9B029f92y3beyaZ2Lwv4fypHLv/k8
FnMhfYroTIXImV/BP5jbcYiiTp+Jed+8PGXdaHvV3EjIsI6ZoIaturrJ1XJ00YA3DxCQ2DjBuerP
hiaqKGLbGUgLKZD22kIyh67vmp+BaUK4X9UjlEUmyuRUfJK4RaASdcJfb/e1dP4sATRduMRed3ZF
ZQSiTT0PpJyI3OXg5dGHmoWRixe+yQFqc3Lk5cmi8ocM+pdRXfBHhaFLye8HQBJDkBg6ideM3CAi
I5wxqe20VOB6KCzY95IDRYJDMqn7ktA0onc+yWJReYV6VyKS5XGJlspdv8uQKAYwvMWXNTKm0sdF
Ik2u9+J5bN+1fr3JiX/WxY6EsfjJ6ft8XgPX/ENvL5ab4wBZFKTxchkOWhd2MsEtbx6dBf4eXOnz
8fTgCMhM4dfv0rQxh+ebhIQ1LNaCDCJlPfYYqMtGtLam+Z+eXxPH22AcAnS047pdpXIcdaZuBOI4
RmB3xREK58YhWu+T8l3xhuBdC+MI2jis420I164p6ukHYWqn1ophdL3nYWq7he2lTLk0QmyESgWb
bKHI2EWR5t8YoCyogbgGbe2xGqROBw7qJ9u5PrJUUxNskrHKq6HbzxdQsfkcaSzzl94whrCmG1Vq
l02vIevKH/KDR2vBQDp/c51dCQdnIw7BkQz6Qki5U3oeZQKaMa/6S+/Ucqc9JzyZIu6Z0NSWZ7zw
y3zLsKaXjP1I5qALm03IBSDw4Uz+ZxXTCJwY5vXsyrGKmaAJpXZHqJ+sMeyzNbtmggfKoIGzYYfq
GKpCjg/ePVKcUYWIMWn9a5u2QlwhtCePElg+6UUrCiwjKjxWQVUsI6+WLXn67DB9xjL31epQK1Hu
GYkfZA6X+LSiR1+THju8/A0MCPSD66hPcYmRO4hYP0XqGeA3AduiYon405OF0I7UnuFiz4STImjV
Qd3xjFvmRWlZBxa4j2B71gcG0jIZ0BnmZZ0akKYalp/oxPIpLsU7iKkC129lNwWG+q2caZNhSgKx
+Vo1KuRlKGU/R7yPrFfHd05L+e0J6m03FDce+fstsPv4+yhyKSNrRsT10OxYED+kwDiRwd/cZ0tH
0+6QZsmFcF3z97yNWiaYu21igPFJFDr/Y4GtYVjASHzVHXJ8YqphA1G83Xz4um3+X/HOUqTuzuQ2
PShucgPqxdY6euxQELseXd715of8TcUetiZSpLcqmONoGIn4/lnG3wC22ctw3UDxiCtAR9YRrPNG
jjsdyItknBbEgvPuBth1ArPQor3AAYaVnIukvW3TpNwce4+wi2cKhRhDp1pmcIsML/5flIagC+yL
/QjgYIKvGjaoYFoXlb4P8j5fAZEeuJkyep8OBXMoYjsonh7bjtuzUaPAoCcDprL+aQl86NJ1IhbU
hTiCFfh5MTAPKiHyc6sP6OwfJxoSKOMj+z/GoxqdBbIrUGqT8acyPJe22qGLyikJ1apOW408mws9
xl7cBhgKyUCM4Jt3idrPehc07R40fDpXjcPtAg+kelrZaKSjeDakYsAnKu2n9yxPGOmytrTcgH/1
tXiTWRGe/DLrlTvlnFEo6d8mof2PBBT4357x7OYFhu69nOjKFjFJVyquA2kK9UuqGUU6CR1hh6RX
8yw2lQqlvTeJCD7zjbO0ow6Jm+PUYYOGkq/RY2T77EwKcqmqhwN2kT4aH9pndoaSzCRs7OI4gqpQ
2UX1syuaPGwdUOYS1Z2YJM6W1ZuhAr2LWWoaNBXanKBMOpOMK4rlKDZWGwgWSMqQb3iweAbuI2ls
3oFLzotkk/yEEJcUL8TCFTaOQHH4L6VdrvrOxx2QTe4JbK0I285BXylvApEN7OIxc3RIKLvTPz3k
xnOTQ5BNhTAbY6n9LNMJJOXinHcZ6m1/5P+eQcivByg7gSGA+0OjqI1vGg+UQrL+S+yLNZAg5e5E
bEZtATq+R2bzBXb/qgdTWe9njPi+DrY1hxsmOg2bDt9vLqYgwLNSZ66Wnq6bVR2CSNbel8AgMd33
HGveUx6Tlyg6igl5q4X4fwhjIcOHM3Wjg7wVUQQs7GGl2OAiTKD8F9IGnOLLF8CUwwu8JKGNxxiD
X8LDTGH90qgD4k5ORGcYNv+d62hugE2loz59vKcAYLdEUA2/ZYUOviZWPKif/ifb48q+zuS9j+hE
9A7MoWyYqaPPtYqYdoDNoV8tXeNNlGZhfRcaxg7HUP3KABv3toLEzTFIFJI1DYkqDKu614q8HWza
HGcDtbkCuDl7+2/Q+XeZZUpNxAc/uaLYoK+b5+SORLC6rFI9RoeLllmTlxOxmDWvW/2/VqDF9qiE
C1/guG5U0h30C7GRmNnPHdHmDNq6qMxEIsx7wwn6Fl5hWOlutCAQ81R52DN7dbJgK4i+NCHhnJAs
1l4Fa5Fv/6CTAU7VOBPtIKA9usvHV8AwvBe1izWuRJHtqGb6lWx4f8LP6yyPvA5q4eWIw4/iNaHD
a65dDpMxZUNzyYQT8Xf5Bb1h+73AhA3TgL3KWUQffo9FiC2bOpx/YvOEqwYqX0K8Iy3BPwCsJLcw
9iY6tuusXDI94Ci6yby3yxlvUDfRyTi6Q/QW+UjgPLaUeMjuXWU7aJSn3tiVQSKHFhZ2i96T7Sow
wp7e8drFsHgJxYDYqZXwDE8VgKM2gYq1lGSQmmsONhjX/PAy/3Q03dePI70AVN01kWGwC12BjWVA
bjdid09A5AuFg6ubuQ21k8xTRVOF1ECY5L3xh37bea5dX4UN/h3V9+740drXa9oaxmv9V/N9+btz
kmAL7xySQmH8WFlwxXCGfOny72C5016ebdTIMYIOJQnJX7wHugp1dm5Wse3fe2aOZqAx0Jd3RNMv
AUnWA2TZ2+ZbRjx8hFbwmnomXRg7qLmtnNZo/CoRMtCYM+IqxhR9LMD3mPgPjAvbWNb3nWXPvYzI
xyUVIrS2f3umi1vIP62k8F6ua97Fmx98/WSCWLUumEExi8lmXUnjx8aDX+3BhQMZcRf5PyqYr9Pn
04H6IPJTop1wnPxntR51HmIKVjcVTG6pIwJTNMcXXE5cgtyTYRWgZF/Zlg78g9ctlNASKLbxz7vE
Auv5wotDQd1A2y+HI5amcnWW4cKKo3oWfoTNwl9uqn9kQQ6ocAYC+z/Vc5cEqeRCnXXGPMJvf5JP
ftClDL1ckirT2ycYaHgOfmynbXsN1BCQlnBeaDe0+1mQQGqn752APl2XcgyCyCYmUjcMa+wy4Jmk
sjM2NOS7VCKSezv3uqgQ9dAr4DY8HMAWohAKvt08ZmQ8zXehAs0qqzrc464QGXwQiXt+t9CafGq9
XuCSQ2+PZiLptiDPTc33eMdCvkgDbV5iWLTb3/k0PeAKs+i5cOB8pBxCQKFYwa/Yu/gQscngQIvb
ZEoE2/n6VB8FcsvPR3xGA/YSzeUpawFMJzai/20vvcXAGx1fVYH3f4JK8llhYd54rjhIV8EyHus1
7KdxoWYw7GIY0ybK/vBVVDlbwi2mGS4oA6+jmWZMhHpHgkh/sV2h+IVFzRTra1iT4Moj5RjLM9Mw
9yDlCtL53KJxGwmULeMDmVhEnh6cjoKwJom3lNj6QAqDXa8oLQ4HiOA0yF99nORY07ktpI3N70hQ
EHSrttKCnLBtBsRQBO5SOoEWLH1H98Lw9ovXbs//kBn30p+mNLeAWLAeXZhc4jV+tgnGQ8FN/S9H
yDFFebG7htP+xt+JJTaMTVJCeYn6Y3ypA6hchSFZIy6OZWvKa/Qb53xz9E1D1z7hoNnsAjcFe8O8
yB+SC1K0NJRnf87YcVhlVEH1PTPe/A8EKDSjmwDe+10Vt/8eu5rJUVPfxaJB6+BnEqK4wK9h1vD+
zgHCJGG5P1QA3zjDqazagioW+xWZKvctuf9wm/eEe/KnAYt0qQBQMQAszZBI07PPwhS4cRP3vHZs
Fd0Wb1ZJ2nVLjS/mwB9kzVoDzzB9Lpyk8Wgul6/ujudTxYUFStXI91OI2PiZxfR3RRmhvciTUslH
i4pEdigp/ppLXx82FzZvK67oKbrsFE3M0dC9eu2T6V5D4pXCHc0Wp21fCDjCbT9EpZ/SwKLXYZ5b
tXYWoqqkNPTuFIGBOukxGyTqg4+aJOO+G7WixOA0iuijjJatd11eDojJJuCs0reNjAXjgk1G7oiW
nJAPlWIfGZE64RT1J1dFQ/psa429tlrPuUNEjwh9+Cw+/F+qlGeCx2S9ctQNan0Wky3HU9aaATRI
387SHUqKlNunVweTKpixrq2BqWJuTG/7JiT2VEUp5AiHWjzF1or97eJvSAgo8Z9CR4O7Ew4ZKZ7t
DB1vwk+dnOP8s95xc2FOCBYDXeXWHNC6j6O3knj65JqJK7ip782EED5u2iQVeTzkAUMLTnBievLs
Cp/ANmteGs8STLWQNtNluUGJj0svWc4myxO+bcaKyF17S96yDwk39LDmXXiLJAVtMQKlq4BOahXg
4UuRqp3zyBCi2Z7DFbO2RgCQj6iHGprS3xZQeGXixaFRzsQueDBCufxWMlLnE1m8aW0MHuddVIXu
q6tizZDozWGUHvqAUWus5qxsta59QJ/kpk2auvhbXo+n+FndbesROYQ3obG6yXjci3SZmCl8HU5V
e/Y/sR/mnkqG9drsi4GL/Bd6SQbdSJH/+WiQ5UiL5ej6DF+S+KaNW6JDTwGO/43Xr9aShAPiab7t
wZLNfc1bOqz6Cm6saMUOSKJFn6xhMMz9/mm5Iv0dL5kUYYEpVtdTbZaFcO8I8zpqw2WVEUrSQg13
r6MrHw9JzzUEWyq1hoA8UwtokVpkI/KhFUmeuLG0Vy/kiKzmqIbH9crX+m0/1UCsiISTiKFJiQb0
6neheW5+NC5lkT/Hmc3IReEpNcyaTdyHKZXrGdkMy2El5Nv+lHcoKQLt0gC50QqwGCDwMVCvBCN6
oRlV4z1fRJ0psWBhgo/hHKXt3stCOJPB+Ah2Z8xxejedHr/PEck4VKege16UPwtHa0NmI/mKPeEc
2PIeMm6vx68RRSqRppwXMpJVZgf3CIKAeOyCv9X8oCN7mdnlJSUCM3eWg4qmv68Jk6r+zRXOk2zy
F2yOpu4WWxl7TP7ETReCOB0xOqDVjvQXzpZFCCpKe0yCfghxES5Z8nWu+tTepHxAXLmJWeC+fnIW
ISGiBM4eUNu2wgb8jgVA9tx3myoY7m4A56sfdv/XYq98/ey1NsXrziq/Oiiz2FY9/ZigCSk7KpRe
0wW+kK4kc23pKWQ5Sr40PokNjBp7PNs7sCzDBrA37N43O49dFKiWXQSXRUdJ2qDFAE5Z9eCWY2Oz
1cpG6tYO98k475WOuMQQcv7TlDZA1ch+KlV0yL/q7a45pEwMXXW5H4qFFZ4YEHYgIO+v3ALc5zPy
w7O6hYb6paebYt8KGKfe8UQNBhcWUbi0tQOaAxVx0SUWWM+2yLThjTwm+uT1GnxPXByVdBwHuliH
+tER3fPhf5xPLwPa4dy0a21upUp6btTqgeiILjfv4pf44JhbpY3MSDv9X38xXIkJOkZNYoEvVQeB
8O5MoWtjOu4qe98CkxePiSk/IjmdPLphyCbbLRMSK15sgDq1DhTwBuUd+ai4zarLQyr+C5m8Tsf+
8wzzR6ZNlFPs5cavuy335qvC3egvwsMCqVVk1B6+XauWG4Bpopuqcr04ylI7xg0/eG8SUsToS3fV
pd1PP5Pmtx5iWQ13yH7H5DyUCfrUfu8PKXnMI4MHlx5XTAsNUci3iy8efwwXqtPIJK+JkhOfOPYa
yS5XLRBU+1FZAE9xX8ygMhC7l6KGld59eozgw5IzoPqC94DW0Wqot5r5GC5SQZTv76B0rIfpHRj/
Shg5GLa22BD8pANV3Mkn1MdWhJxSLDX7VN8RSnDJ600fbM1RADAfdvXnK8sybGXNvLPmQ5inysMg
jCyIsfe2lzs+sAJN2qbAN9icxjKq1rOCSl2x+QMFLsU2Ztse2c+E84kHrd90iwLKbP3UqskfX6NO
dbHITedwmy35iiSot2+KX7BC6ymm+KIDEvAL6neRjGVOhZT5O/NhdLQFZh2PkwLOX00jXx9jVG3q
AHO/Zwv7jd3CjkEKYUMj9Dbxxd5k3nzD1g/GFrwTzjG3u3X9qkqkNnoGLIiTHQlStkebzH/cGnhy
aDeN/oO7FLiodENmIGV04cR2Z5XnokbFXYTyJgorWPqpehCAxO2Vq1cZDS5JqY7HO44NPwVJgrEU
q1JdkgQTZxQtvGSgl+vT0dG7Jm9LuMuDYxHFNqYtzXINfcisCw/ZrB9AOP1BB+N4Nm10Wog/9A38
9hf5S98vBPjKxjFA3npVkDyFbLeQBGntCWcA+AX+qUn+u85h7Kzg0s+s4wF+G6dZjMY0Tl8Wl+yI
s/tSiBUeV7cS1skV6VGS6ps3UDee/GkkKhCjCWR/ssQOe46DDxcLG+XrJhuh94loOsyZqk/G6MkJ
Vzsk8JFxxHLch+qf5Nr/T9MQoyb3klAqZUH/GcC9xpbMAw6+8+jOOajSfkN9uOrepviK0al2vnyJ
tB93Whba7FulRFRCRghRTgq/clowLoK85HH5OAnJreqLPgI9RcxjxBuP6/mUXr/wakmwoIpcdyBS
rcf5m3hYJ8HJ4zcNnUSjyDQxbH5l2PGRPA5pMr2dWzZffn0Cv9LwOr2Gp1goMYZROr9S5uD67Sma
1w72leJTdFqLq4H88caHVRlh0/tAutv83Kfb19i7q8zNGB7WldOHCyT9Jir0SaXjrVnS40yErLNy
gJFChIyVsx/QUfrMGTG1/i6VQ9lskkv4jMzN2XsMQZUIOJIQ5qQLPfcEdQGltVrpjhX3DO0SqrZ6
Jc0TpaXS0TSnmQtpIwaXAuYTd/+xgKwZUTETbj1iuaYg/+DUOgnXrE4N6oJbJGXCcvbnnbgPGIbS
xRyOJO8HgyicP6nvv9Dbyxny70v3q7r3JS6fUFW+GWABxRfbcB6c0bLG4/VMVJkP+6bxwjk0FEif
1xxKUcg/edGwh5l0euRfeSP/Ni2U/O3LBocgZ/yliSZCe1E7r2kwPecSHNY/II4xGrJakPk2+PlY
JpPv9L01b3sshhUr4AmpepReWSNdw+in/xa9KqqqRD0ToNrPeEqwO7dkPJx6VnC8GsAYNR+amEah
1OEpITnHm7h7XqpKrDA/N+HwJCb47twcz4Z8G78W4zYaJH8QoZjHWHaQyZlHOzk6EcAbBnfc8joW
nO+WI5P4RODumL/cBga0/yk98+Wyr46fDdezOy1RswTGp4HLsxIJk52Klu7vi+2cfUmvm2T7bPJv
7LB7Q9QLcnMnM48xaJSKJq4/rtv5p6IlSV1GyAw4P4x2hHxJDzNAmQ494m6+QtOXirZrr5moKQA6
DyddnTP00O/RIVRiR7xRLWzNCVlPNkvq0doxe6kurJHfqp34AOPYdi94d33XbL5pzI5noU3Z6AxC
2tPPTObggJTphof6fxlq5Knh87CJ0lHk2d1ot2efzPmtRf+CGWc+415pynArx/5E2mr6QW1YGg3z
d54Un4SgEMQowFB0EBYDoLUi27LW+tuk+1Y98UyQfBypwd9ZuVPFtbBM9A8fW6gtM71r25cXOI1T
Z0K2lm0IagNT9pR7ewacFOfVv4vcyZ/yqA27BFCKFxbBj7NnASYO+fho0PIOHwuAfbOdicplHQBW
+dDj9yoP2t6CGolw025KP2AfeQW8BcLlKgX5mhyaX1EbNFDIkzqhK97flPw9u2DI07ClB8UPU08Q
4HqXrQ6v+PMI3wYs649+edspv1asORQorE3zjsbsxmJc78lcDdMmSoNr5WMqVyMPtvei3BAmiVvM
FkkGxDZBSVsUHrnd4ql6oQmb1ulzgX6C1s8IG6ifGmy80Mf0ZHazHc9WPCbMRQWEFhnTFzMLSoQx
rJaiiSeZ+Tu3Z1UeOFymqNgwLe20v7kfUQVGNGXROM4hnLYa1yo2Blm2xnstM1Gd/yRu4G++1AJG
XdZbmSa+0LH9lT3wpYPA5rznpJ1plzjGSgAeoshFqEWdsHXT2NcqzKk6373VVNd125CTz97Y2kda
YPTkUg4LgkGaXCNt6mb/0VuTjzX+OvbvI8Kfg0LsdEVjUpWqyco6QgvAUxmZRBVSeutRy/o+9pFU
f6nWEjdmMtEkeFspPEPoKVjtupvgjtTC0nDD9BfkGn09ctFMj2fOFSBP3MAwzCA8Wrh3vqkYLUpX
DJMlYJdCW9FpI/44Q001U5LH0bT0M608dUULBvR+F69fPZhVJ++xjZrw4V5QIwNzE0rbmDSS2YSG
FwroQyvJeAkWhb+ThYrqIRUt4ORUtLwSVkrf3eReU6T0iyHysgL/RjEJG6JWPgGyfzQP+srAL0AS
1CKNCeXxnbKN4GGemCIa/SsrcSr+R/oJ1uwP8PYmZQPNWVWRmzC5l9snqVzaY6BkxbJzHTwWZX2L
lPBc/zZemiWCIkS/5qrw+1LKHqBP69LHF2px0CwZ2bY5QLQeehRzCEzOME4xhnHMuL+/7OU3FuzN
pBF/dn+e7sXDzxeRCnQBPjwi1gQr/7tYIfcbaOaDqutPUQEJv+pXwjXQRDkrTXBfgAHtS8Bmgvdm
/oNdVzuQ1cET4RIBTpa0elyWlYURfkv7LyOATmq7ikfTw5sMXI4Ju8bqL4Uf77zDyQAOxbEV5OTN
PfT8noQcuyJVHZCvwVZw0KOvgY8WO7s17GShMOnJqQVv9dDCBYzbxZfzfZ1LwYQxqg93aSsGvoL1
plS4HTh/UdKcDmaUoVUhAAjDiBI2n0xc4dw7jI+VE5aNTU8DjDO5oih9IIxwmWIU9n+F3e62xy+Z
Kf66tg8sA8FCHs7jYYxeqLGNXGYmjLkJz99eAXWNFS+Uq3rTjXPBucCQbe139UXjytXaWK2Ho0bl
0IB11M/zODHgRl4HrHBNhB9ehQGaa4d+BsLUsYayAyDEnmcTLBe5tY+ISUGXwe9GAncQzcL5AcFN
FSsiTgHEQ+3vqOWg4MPDGnKcRc4OAqVnqppv/7R/LXNOwvwmO53SuVCrKOr1jkcz/eGEzojFnOYy
emNoWxSIPJhi4xFyFodQoMrHI9l1aj9cXFfHeJMAz1AVmqD61o10h7Go0wp0ZJwvj5zX6ykKdpek
k3ucAq9fdadN3bI7VB9uYBzGiMwkBvE/AbqzTgD9VRtvmb30SrW3FooYLuXocmd8I8J7mjVCyiDS
GrugFm58GOwb/5yiQcXal3gOjd7VBm58KXopGYNESKis5c2mlSmk86UUzIvtlRYmBvhS2p774LZs
ux3JEPSr3dIbn+KcCMLIBlgJvYkLlh8fVQnOGltGMmZSmCCxbpt0R3tTibH3TuT0uWPlmVFJcu0M
l55j9WdWa2fqrZSl19pY8YHOajYFywhdWOrGtCK0ME/AI5zzqNlLk66KGglsLYJKSpOI4A4HJ6wM
JrFKxRtlPnFhGNkMCQgEQWY7aaah7YnBJTWblitKE4Qr25m/UGC0cKgRhBp+H/UQKIDz75PbvfjW
7/DL/fyy/F2w2oF15IFrXASlpXAzIoeRnvQAiyfW3gOcK96ZFY+z7ZUn9aLwazSO2A05hNkcJ1M4
4ggQG5eGNrM6YFavmj2UYemrSTqdCn14BB8Cym74X7cyGLfacDk6Vxtzqe2bZfBBxj2vEBJMwxPL
SexUuYgTMN1itsfQn70mUK7tdD74rdf6j9LU76dPeJdSI3/QG+/Mfjsm85b+HKVnj5wb+i6NBi6L
J/S3kcWsL8d18FX5fXEgKJDy0KZPsz7pK8d81eE0FWIYuPTVvdbrM8z3EzT3m1uBhpk591ufXdFk
/wtvcdxR34vg4oB3dDXs9pZVm3+p8ggsPMnPi3Wznp57/dg3tBcZMtw7rtT1WMigNnsbULclHQtU
1lzhroKpSoI4WZaW12UKzujLHHKCbyL+WfDTcHSwESDmKWU9BV/zlRDyVpjkc2kBnfiMoWjaRSR/
5hEyhV6fDarMpXjhufcHsTZyuAa+NGpiXp6Nx61869A7XgHt9Ub56ObUK+9MUMLiCX+wVopgu+Jm
G+CpjiW87Q9Lyzo/pl/kjoUu3ic6rcmMCJRfZ0LTiovcWZI8IH0Q+i+/Owe3QETSukC2K8X2fSFx
Fn8s6pFOuKLUi7bo2QZuoNN6IJvM9p9y2l7DJUvH5ZeDB3bxwSCFHIDlK304wDDKOpTjOCc4YPqK
NO5FfqaRyqyXVER5cK5YolusLhS2kUY1C2RUzYZQo/Rs8ZaRkz+vYd//+RHzcuGFOmv4c5qtUqHe
iFKCSBuJRNhQec4vT/A5LzvaCCftYl4e+UqHzrBSNK6aCCJLo8/g7FI/5tM9DCTWAL6Qs3q6umNe
KJ6Lch/NuKEbvSWn7lLTVJNvsEWqEIsrWwDcrISaYe9ae1hBwcErkDpe/4UgFXdOLM0QsdgTHM3x
QiJxVAB+lViz3pAqoyun9JWhbLRju4W/N4d+HGt8cFzbsVhRmB9rlz52LndaPsrYFbtiUUK8f8ff
+IjD3x5Ou6YcRQUNXiqzqtpZxA6iIt6rWpvtrSqviu3V4QkRCqncQo7Ydn+S28A9WD5i8j7KU/fU
c3TNg7pLzuopwFk3g1Uib6HCwAJm46v73eq9z6+4bQZj1etIOVc9ns0L/Y9FUwgMMAJJM2Kgsin0
mi+jdgTEMFzQyvdzJ9C/udb2mHvDCRB4K1Fjms0svcOC5mZv4en/Avkc9GSohoZ5KXwB6bAcsWtm
isKIyDUJFuiL57+rYuru6EAHKnSmWmL3fEurVaXpXxLxX4mjFCpAnBA6K4T/397iPoYdfsd5OtYi
GvjyQFEb6yebXi68Ghvpxle4Vna2g9hKjL+EL2vPLsAv90YZaJAck2x41J9PAJoLwSq+x6e74iVu
SFSPNdcebXRbwKQvcJ3S9rSQrM7xgsf+pOzBJeOMHIt3Sq7D+00arW/FhmZJvQdx5UzWcOEe9d/e
Oj7rQkm+MRecRahnxTyJlSJSVIgSAB5QKUuVvJGCKnR+/wSyewQlbikWf1EJqdGkmIzcJAqg4Ru4
bgabK/Hscv5ViH8exdmK8D09tpfFreiU5LC/DbN8kMQT+CamZ1YIwR+PUB7CFJ3cviLVS+0E9qS0
87PLYt+z9x5+R/5dc8xjm8SzW3OCzl4LTSf+lXY+Or9M1+Io7VaiZwgHSTj5cTPxi468MOeYj2kz
lyTim7lD2LleaSS7pGCJjh25xi9ENpYfJl/SxDtjREaH4JoH0aEDWArQzpAL7E6CnyIMHGqrbn7j
Gt37p8LHppL86pDDGSKg+qmxqDoG3euhko7Ew8QR9YXiWpeNuPq5I7DUZkNDAOhpKI66qJxH4iG6
Y+yj/cucgPd6J5ii1oakwW/Nl6LppPsfeuvPVseogXa3WCPfAJbXM+zXNLmXIrVG0E6jybfxrdIQ
IzdQnHZEzPzHPc3nPHWWgBYFaLJH0FmZLpmYO8Z94qkNUh2dIrjUk8GtFHdcvJ8xOlWrSy/nxJPr
pfpV1Cvb0bFKTbtcEUXhEnQh96PX1E2pH0L+7PEjV4J0th23zUoIcGw7WzH/1GA8V1Xg9n2GOSZ6
XyFwcEMhosrFuLnMRTW51p5sSmymKP4j7gN9azlPh9jJgtoaxSMKDKTJWcXu66+ZhZXP/hXkTs/Y
VCy4o1j6yBzHW+CUhgtPA4XhqC1NadmPRb2Ch/WWjtfiCgQLnEvm5NhzEHRu/J+kE7AVD7cw0dRz
f+UCGTBVgeics/qQ1N2GzoKE2ACgoFP2wmXVDCkdNpSwiaYDSkGlKSAi3yTBnHk9LenZXKe1EeBb
RI5VZfKALsdjJCEnpv9rEw9zGPAyV1/6ccYJRreVGpORsR6LFl/K5/QDyZoFO7+ja8RChnGI5H9w
OzT83VkbzmMmWiP39dlvaJ0Zu9UwOu88w4FGX5IlzgrSOBh53DqvZnkzRUwPl5pvZiFJ/egn5B0v
ORu3+orlAkw+u8TAb/UG8rhjTK/xucYBIB2ThJyYs+61fb7eV+xBRT68dafcQn252BOYXUZxqn5m
1TMNy1NM4oHhCj859sB8vnUYF0mUiveM8BFkkdEz8OsERRg68ApqpeiXD7LDjEjokW8Sxqx58t0U
rvo+xgkp8R3oLjmdeJJGSRTE/Jw1pU/wxTvLF6Hahf6oWQU+HMhNw02dQKX6Vi842OD+HjyqF0RA
HYTZ2WU9Rr5g8Ma6EXF8ywR2B6y2U1udkgErNr5uXRI7a+M+mhOEw0J2VaHBIv7x9TaDsVU9fQWx
xLQGlVg9QQQFe4jLVrrFLOm5X8bUpmIkA4bOOQHCrvkNN8jtrCBNX2WHXWKNoLuinJe5fs3j6gCE
LQGK1+C/vDjc1jKuEtP8d2NcXPhYQ4MDRatdeDaCay4YiBEphc57wqaqley6J+WnTX8/1sXyiPtp
Z8PlpurpHxGKgJ0L601RoILlGPJ5p4fMFQcPyyfRPUrhIxDzXeAglsF8jQMgl+cIuiT2gRqM4teh
FZ1tyr8vK64V9fGH4IN6iDs8uSxh8PROgrKFXFLFbKTYfDZ4Xm8LswqIPGcwiu0zbXfrrDDB3s+P
el3EKviedKrN3bEqYxQbmfjHUb4L/CdjYS6T/qPuZTUO3pMKe4oNsB4L6eq5XEHiMtEZ6/yKVNRw
XKd1R93vz9RtqjQMptal3hYYYOsBE9Qo5+nxKXY/NFE2jaLhoPtdabhCymAolxbYlmTqRNQs0onQ
tjumFDFvPtXPDeaJQB/EPuhCOMhJIkAEpry0gaxkDA/nD3cGXfIpe2wAe8WwzKVItbLUaRDm6HqG
L4TvCt4WEP6PyFlvA4UJm4axVWImY4R0QYCp8aobzM4pb2I5i59AvFc4Lx1wDKSRBaq/MuamGWgN
sh6QbhqmtpOt9LTQfbPgS3YBj9W74MGwQI9D6v2ezbFUb1PLjm6y25FkuFWUFQLgpLDaAPUwT1L2
asMfwknljLuioHFvc2uBjIUbJRoriEvVVX+Leu8PebSaQqZgXm90dEP1gJh7Q5F3WPraKsdr5+nH
Unt/kLlqxyxTeM1LlpJJeiL6tMutvQpGevE2IpuBDTQnlDZPkpJ+eqpubOwqh+DkSZg/YNFa2ymV
NlCJ5tfU59CyC8V3D4kmkzicVn7QsZrAgNQoRZfTkpzoJHmt0EiawmWLcTXXizKpfjv+1nY5Vn8b
YNC9gAccX5HAX7/RSS303dQVgUwYAQoV/g5qjc2WuEQ3sj+LG+uKI4HrV7IZO/XBXZjJeo0sqNPs
KkhYz6DdHkZlRwgSv7qv5S5x2mqyt3Zm7caIKrx53cz2R5yJumJH4A7i76UvVEx/LtXntr8zUChd
rN+DsX8i5K56jGe6hh3UHc7942stV9Zm4WN2nYNKZ0kqK/3sXE6ZReTRFxzCEJXdoBtOGlgrDcXg
3wmTOd62xcHVzF/CWif/mhYd3utrywfXvbKdjklgjV/rlEpmwkS9HfiIIeqgdV9BDBREv/2sSyay
udVuxIA6FciTqWG7JcDC5hTsRsvagQ7HO2rW2GAzOquuqIEbOernhfh7ZObz08uD79CazaoQCanU
Gah9Q4SsgqL5sfQEbUX6QN/WsOtxgX02uVQGxvQIx7Pmi2iLbL4m3Ygh7z1wCKWfnMg9rlxul8Id
xXerFbqGqXWiEEyVaJkoLGdpLJwuL+vAy7LEw0irhrjtv0Qb/G12M66rJPQmzTcCEAucE7ZDCDcY
idtjJyHT9/0xRV7uOCv/LRXyXeJCeUjvJoIHHlBNiecpf/BG4Lnx2aOntx7JLGmaV458Ad5rb/Gg
rDpS9IZFLdj3geFQbVY53RMyEnMYrC68zpv5VYXnsnhZ8/AZJnw3JDYhOaEH1ThXyDgqdDDpqt2s
wb7qBo0vGDVW/0dwWVwC7cHbn2WrI8rUfJivqRItN+J7zSmgcmrBGPtMrSD4ycmuiffWLwlyGgRY
rTPhhRbVApfFRqoBEL3Ua1NjRlsMlHCwwivVfZAz9TnK4vEnX/YZG8r+x4gwPlobcOD1ErDpqePV
6QY0H1KjagS2NCf44Cb3K5bpj9KITOtvsqGo510ZAeFJ0D2ldYlAM/wOlZ9g2TTr9st+VHxBY7n4
9MzQHtPCBXmB/ggX6O3l/60CsAakjAEeWj7Tg1qcnzu8JMKManP1wqeoR5lQ5Yp59MNgw9DcOiX0
QV774VL7DgrPQiXKrFFg5dvOHueIDacRs5hz5SOE9xTUQtP0yxkZ67KuOKdRfoa3Kawb3d5/guVN
CQCV68rOKR2Ug+twznbOZmezuRedZf+jBiUeAxCt+wg+5z0228vDJ+sj13gP0vrp8lVglVDrw+Zg
TdCvf6FvTfWqbgWJE4wiQgvDb0ERUPOcBJcYaH7Mv41FDC1SdQ9Zgfm7JnePg9jJ0GOvq53URysD
s4ApPmJhrXLi6s9PTEzToOMFGi8Zz/+q4FsK0U9gqlRR0PFFfaxxA1h9+ZSIqpjzVE4e4JCPoBHa
lo+OyW44SqfcW+eObNg0rIMPBBPi5o/hTZ/opeMBgKYjTOA2eaUH5wy2j0GnN7DRrFm9xRT4lT2D
VL0/L1AeLlMDRdb6mdB00UjiHQBgncp5zlMAs1Z65I2seIT7NJl93sx87BoQb34wlXC16gId6B2+
qg5RZ+WtLcYCFDjW1bycbHzNb9UOaprAEtwo43HDFNWkZZdsHavcEH6B7Zjs1QHhnk2IEZMqZmu3
2j/QBt88PWvWoh7nEEZmAq2/4M4LH5qVp9zE7uK+tW938/Izb5I128pLvDUDnt9ouCZXtgC8ipm1
UtqMaqZFKqrzd2r57NDijsRaGwniGdYYhM7Ckrurh93Ohh5ox1eKr4THGcw//7cgcj0Vwmq+lktj
zsnRPq7vXE4W6K+f56v58qn9gipxlCAmMCyVoVSaeqruUm+pwGE/AaYGYcuKOOTNEAUOkX6Surkm
qZw9cMJ4kaKEhYr5LjcJYqhMrsEghIfYU/JXk2AFlndJ6Bip6L8Yw3P7xx0Gq70BxtsP6iPtHFFU
pww60Y04o81X3fldzLdiSOmQh6YIEr8QamR6a9Z8NECIb0x+3KEpxDqDLUWAQe1jsrYCGMlnSF2x
KOE9yWOmdi6NfAYE/r5UwFD7xVFTwflCS5lEWNaMLa1IUJ92Dra1DdkYznm97+aVdjPXadXvF6gx
ykcVIRbX8C4LW/3vIu+ZfCqHIgpA+q9Ldgcv/I5qSTfXUZRyvpzORoIylkc346HH0towWHVabDv6
xgH0fx26FmbwRsbJyeJ0LU4i1pOtCBUwG6Ka/eCm3jGMdGKQYGEaX9P19lPyCfrjZI4FrcoFLkq9
PChXyIN7h9aVvml2y7N/+hjuMz4qA9RM3BuQzp0muzrcO5lCcyargpy7sM3lYnX8mV658C0NAJ/F
auAmcBwUy+kRnaCjYmi2yNbPQp1Gi0OTTDMWIxWBj8hWx4LtiNvU5KYccrb5heSaE2SbS5vn2lbr
gXUOj3WdsTt446F9I//nbaYdvvJUU3EZkkC9O8x8vhEgTGyh6odyYB6w2LYZHVSX2R0w0UeWMAbg
x09fCVh8fGqUFUwQCOXcXJ2Tw9Xiy1NVvqDrU3UEuGyv2CL59obVQnGWZbUskmR8U79FRZRU0Dm+
e2eD9uu/d82O4mPUrdTV5mXRf3I1c9D7q75y7d7aiTMOTBn2qmLAcx3EBNEM3Xuo1J4087uOoFkj
ruS0nbxZyla+4C4+tmsYOE7h58ZfPd9Stclo0SFmDQwoijjEsdak5TfPYEydRDshJDcvEVJxmbVJ
qx8HqvvScm70q7IIGvQda7vKMrerP5j3iIFyLyp3W1fjRuyBnYtDEovoqPsq4UQb/9t381CnRy3O
YGxVmWl/S5hBAWPLQefdvejgCIGpA/NmYzvkJuKBNOLBnQuUEgQer7aAzPGRpTmEgrNqZWtx9tUr
3M/ML4MYgmcMiRetkfWj4tDM9izVCwATpZWnNa+gvEDM3tEIZDMhu2uT+Zlj8iyp4AN18WEpYv2C
mnPWRhnUKvZRNz53AMOke53uVtHUuMatiBXLuS8Q6H7Y5/vFY/qhuMNqdKW1s08HDnSb1cMXgdzQ
hVkoThUsChYrbaMoAavSM9CDCteKFnKieu5GNGqrV5VxcV4Y0/KqKuCjOdmF8nOvKZddwNkuybui
efAawRVOJhykMGSX7WKeihR1Db2nNoc7X6ufNLZ8uGI15T4/TOTRL0Xgy5sbnNBpk5je9Qlp49/y
rOHkCc6FP/xRu7/qaYRWhu1fCw54rXowF4S6SRFoaNHT0k+6euDfh8vF5ENUDWZna91wylwF8ru5
5wsrtjbr5jhhso7BRJAHF2vR05wwLe3iwo4114iXqkyFBqQSIf2tipKJeoiwBUbrqtCVan35EOD8
o1mbWvThB0CHyzUzEpIrltGNqHGfO3kaatZABnL/lnulrZrCcQ9WDjYsKocxL3nkpzaL5kkC3hlG
dfitB5eTKrwpPKzk0dzDxZQcVTSMwyrmR/fKZ9FFoPiDoNqHL9srvveJhlEE3o2bP9VCOnplSZ4S
TCU8pi4oyDFGf/u9fS7Q+V7ghj0bK/dyFKSTCK2FACj5aFIJ+Tb0oCc16J81H0P8WoLkLRkAbN3D
GNDerGg97GXCu191BpbhIQ7jzGJRa6VCHKGK4w7WgGRYlmPjkBEKCSps+fDxriqWJK/1hth08u5k
ACdTVCTtojlXyi/T28WXZF5SjnHtbpV9tyUrjiEJ30tOq29LKEl8kctNZ6znCB8+p8+FAErgvPp/
AXN3kRCwH9A4jU+eGRguywgIK3WEI8aSrFqBt3mBWq79cED0eE+ByujLuInlYSx63BchoywFdllA
6zh8+3Ljn6fmwzbFgdl4nvQk7AvfXThz+ZPYC8/NI9JHzMQd7hNguxJG1kuyvn1TXiobvxsLD/jR
S/ll9fI24y9Z6a6vtjGtAhg5nXG2S6DsollME6pthWZGYJqEeVwwevCjcbtiDzCV11IOZS6/FZR0
hqcsln09m6bmCGPhfI3gMMGLvQ1gFgg9HOTq6sRMpIgSQr1NiR2ol2AFlPdTqRzEJGEmbv4VAJrZ
J00D+CwtrIpzmfZoeAhPUPoLvxcVnbNjAqskHpZv1EB3U9hR/wlSeEC2gCba+SExu4A7GPiqkLmK
wT3MKBGZD3dDwL3Y7KTUneBr7M9ZgemL7kmnc2ONawq+njuNDU9m6D7xdygL/1W0un8ehzFxKNF3
Amzz9K+xmfRUmBuFMUASxP1TfFvpRLDBk3kv6BxVXFs4+IA6sljHNOSEq/8bH5twLGxB08pJFoLW
QdVs9xCeSKIYQxZ9on1Qq0X7W0Gu+Ii0jjrVTqek04gxz38ujuWMf0qLpNbwOHOC564LvOdan3Y/
FsNKOmp4HtGy/u5Tgj1FEmwf2RAeXtAox8eeUfZmfEGxZiZPvjaqghHfyn4+iPU8j87We1W7RVBC
Lfm52+N9z2hMYF2xdLJn5/nO3qaznFEs+DBNLaaaKbOepDfKjZwwZseSRnTkFlijZ/TozxWLqwBW
aIc7DZTidA8guFJSZaTC51HF4APfM5jy1epBL/i0i/I5yiBhhUeSD7JVt6KsJMI7iGeqNpJHWfFN
7Dwlw6d9mgOGVR2T6XsEnVnDI3slGOnghQLNKDmqIY5DRu6UVth4aTmLk8TkOuvCqTt9OIdT8XDD
gUFWsrMnt+xsnsqnbtMd1sObNOaa6AidcnjEctycqnxqxEd3WrajyySKkyscyhMI2q93wMD6Qrbp
aVvoHNTNR9gZOuR4AvtvXbO8LppHGvdFDIt72oD0wC4893tNvKruekie0j4gmOrVsM1WL3VoAlJs
3/xg4SEAwMUVm3Kov7pCdmhZE0yuzLjaZCRq7v2eHiF57WF88/GqPrWDKkXJRUtgWgJWJ/MSnXqi
1OyQmrpyvsI0KSpmkAmv6+LewbdPym/mANaXm8UokLMgqxjSA9w2sgv4IYcQY0BKddXe6WMWmebO
r88it2gaKlYdqt7lcDWZqeeSoN7jbmpFXqhfz6ByOO7DLnxJQQam7Zf5fLFpXE7Ng1Y8XkPSo9x1
O8RuCDg9db79Wkm2T/MKnQTKr5hhWD2BOIZ/8hWoJ7UUc2zqAW9ZvxCithqkEyt7w9kcsDXWq4xD
IeC8MeejNdpvV8gf3W83V79btbosF93H2Esbz8wYMBN0ChxDiHOFQEdDTmkiK7yT1j2BY/uO8rLe
lm0knjHPSMiFTkDC7rXYx4V/txZYEnFZE45KQ9IMym0sg+DxB23zn+oYuupStz5Ov6ZKmQm0asIp
NLfnoyCamX+mge7TPcRhY44UJgQxF7tEJRYcP04LD+GXOSaijjnWohdWaNMqSvqZwd6SazBDZPgk
ovUxwuf++IWTdS7UCxisX1YmJovaIJjPx5yKA1lthcC7xpTkMV4FXrRDg8i+lFhIflwjCg4sKHFO
FzdWblwI3UQDNayGu+EnLcjuOGJM6uEw2CdRIv2nHx921IiYhGlwYIB8mTzx/rlhPRsfNgzI3TCs
axNoYJiARA6G0Nia3Upta8PU41Mo7vCgvJS6Aw/A/tYLo44SQ55I1m0EYcxTICk2bg2mFYNvOueo
pCekKOKLnlT+14qD4QwcIPhbPpKRmygLUbIMH2m4en/yiz2VYUmFFrRL2g9Lk05kIYQu8d1kaAPT
+BcHiczj6Xz7kN3wg+xirh8WkL+P/wSj/oE96B6mk40YuKZIt0Z1cERuOrcCXjxImiEotRgR2DBU
lkgfj7s+msfYHpI8c2aBrv8paCkqECoiqgb4dWht0YncUeLSwZ5fLaLP4bxGd3FOSLKWxNA/h9cU
YOSS3qUD6yXNvqc+9gLpakiMpY2Q6wQPp1B9J1qrHGb0E9ssTEiTVmO+nx6dP+E63iosOxazdWA0
aTn3b4U7VLL5VDCxflIKtmoTfmbfOIoIkz/VtrptGajkafwh2rk0+hNRPApOBgXby3V0DwfQQk6x
eeZK4HUKbVV1LoPhWiWjqr0kzjHzGg/S8Krb17ENk87IORtH/5TAJNEyYc9jWJWHgtpK3ZAAp6qI
fsfmJD+gYQUX6ii0S4Vxq0sjxaJ/aE0iCTFirxEdH9b8umraN5wnZYgnp90NS6YsK4qAiwSScpuv
rNLzo001VhXMrswpRu/3yziaqE014BnsLG7SOvW0k1GhehC7rFHwQsgVmgBR3r53gA5aCpwTCJZ1
cdfj2us+hAwHJl2BS9HiQgFOAZ/E2q/dJhrHW9sRrx2o7xBuh8OV6286fFJDL278g160ZwMPNZP/
JH2CVmweP8CNqOZHpbsX8kc3QkmlFhCyNoFfmbDtmMfCaO3nblrrnkTXQ78Hk4SPKMEt/tq86Ahl
REwfMVZDAx5HrbOoltaI3Iq+tD+KBi0VGoSwznSOqr3tG4Tl4XG4uI2z0XQRF4Z02F72rpH/c0+D
siIqGP0FLGeNv33e1Tm5cHtfBMtBQF7chdEdVPyZ3cKGe+5EtS7GDjAL5Llq6egrO3A1fd8CrBj9
56oazhSQZalh5PSIFkxJNMJLwnVO2FuPnzHO5iJ152zK9su0tHwhSoRXi7WCoe+yFFzWzerhkOQF
IqvD/51+20Ch6skAAM6lOoFxKA2aa7roQ0acE1ZQ4EAOeok12glQAPmRy9/wBM9lkdGIVyXLbLry
+w+nsNvVRnA9V1CJi8lSWNE0FPFoxIN0nTH2tzKhGZUwLhMJairyhW8hIQ371MUCnjwV1E2p/pP3
R4VLlgRjtdxyLD2te24v48VR+W9h/RXT58lCUHUFy73G4c8TxeaeiFMDvvIm8oN2SA9CaArgwSqh
4IPgQG6ajKwSsmd4HfObKtcLUUb0rI2D47zfFPVmnO4+yrJ6w3HmUB5JSa8Z6EuC+35KXeG004MS
V763BeSJ70Yq3a16R+XIxiD1P8G4XUXauRpske4mJAArCzsabS9o3dBFvjBMKbsoLkr6GGzXxK89
je5OY1wwQPXDGjK0y5GIVojsSa9N7YgsKCEDx1hmtcCJ3gtdmRk4l2NlDUmiw4W+MG8NTP3dM5MI
aa4HPR8mUz6xS/slhIkZbJjz1wlsdg3XnOSt90AVYYC+2tllfxS7L6xsfhrQbxplILy9XPdq6/dQ
JdsZ1FME6G8L/NuoTUvHFYBhEdkSqQviAbFSgVWooEbPV1hIMR/ziWQQ57g1MrMUKzXHyLryoAY1
eJ+C/Z62fEldZmyE7kl9d8pYRFDJypdkT48cAw+EeJ6QLM4auyENC3Nw8XaGyny6rtsk2I7KYi1Y
XV3QjmpYNOv13IX1RnwKk95hRGyWBm0ytfBR3pu1eJvCvqjqa1FCjwCyzaR7BLPwsjQBrhqZAiEr
VqaIKwS0dxRRuxDJ6czdnorpxOHDnSsecd5K5jv4RhK/syPYf1iON8Xzlz/a2rf/FgfpiXz71TuJ
p5My/Tgdz9mQjwxeVIN4XH9LhyOCyDxdGeeWzZZ84jKRTCrBmS0GZN8f0qQs0fJyQtagjg86F+Ag
ZFR9flNJSomPIHHCgKr4i0ZqLmqgxgisV5EuCYnIIfjFLBkhi2hW2dVgZ+bDzHVjK/TbkY6joBO1
bdw2HAP6Tj3noludWytCJJeNt2T1DUIFsUNV+q6ALPaE9HgVaS9xnt9HEbSbQq7obc3hYUtPIxeX
7l74Rvi8WqK5dpqhTT1Bp7Im69AOP9nIMw4nRHMv1Fja+bsFz+0Ub+yWM4eNKfEchGMXB0dlzR72
/xGP2O4Iv5OHAdjennwIHgcB4t1vt+Bo+kj+3UUUdmdBVUZ3BuNsiOZRlfj7hc/PyGVV2mGmCcSW
oGFx4YCWbJZAUF4gl2X1d6gDawZ4nMeML+BCl0icHHsbJXtgz91ifr7D9hvGfwTt7tK7DqgWBVTB
eyXiaBMVUBvngiZGs/14hpzgbsKSxS0PD8eELhPpA3vxKd84rv3qPs/PP+oKXxrnupJBxSxefi3F
qOgX7drVIDtCjaSoWtuuemS8Duo7wx5tHqb3HlvuXBGFwAzg0T/T1/t7mp7cYTpnMMeqIj1mcVTN
bcpqI6E87A3ulycWoAHJmkgOyREOxRfIzwzYh6lIlY3C8sRMmokHylZP6Gg9Dn1PxRqpbU5FFDb8
7+n3hEKC4eAY51AX1J9B9hogyIZVQcTNii3hCeO1cLr54OIyMMGhWoSP77S8Pw9vS8yzRHMncMnp
UguprwljAbJEl6i6iar5TzG+VQq0awBqBuyQU8IUj7gzNwdzgMhaj0yltZ0tvdUi4DY+8/QVKKSx
a2uOQUMF0+rDdbN8mckeY3i4eKDF8R716vWhGRR3/SXW7Gchx1raa2CrJ/zyCD1rI+YFCKmMSyPa
RpJfll8rdbB9Sa4YgUIC7rivmstAcusQwScKtGKO6rE1NJmyw11H9frXorI0YkZZqhUf2L+b+uUm
UkU1X6EhjmYt0O8aADL8pz4jJ6ouSvgTvrm213WPZVDUODHjhl2jcEj2jssGGbINHfqsyQqPG0v/
i7rC+bcSiO/3Hgx/3YZfy5As9qjn6g19cYwFPVzIwR+HhcEr1kWM3vFpi4xLMB3pEKs885GbU9TX
o+M16UjruNmKkoA4V1nbgTEarSLO74QqHf3ZXZ9QckKaaKt4Scc5LaY52BAeGCaacrNDc0dVmx7t
5Df/zBTHgugX6UNew4fnzZh0piKL5JRZ9wi6fwfpKlXy8cYWDOaRflNS6FCm6g3xSzNjOuNEEouU
ocwtqpKquzrPk+AuxiNE+RY+bjQP1uaQIDAVYHLgN0ouaj9s38y6vUBTAAImeFcRNShP/Q5Sci0r
zdDGhRMgl7QxxPFbw+A3r/az+x3qWKAlrPK5lgWEOLfQCNulTh/jtuqzFmzgw11eREdaJlKRzZSK
OHgKx+/wQ+CSIbl2MDGSqT4h3Me9qfPcN/Wrf+49DdozYq31yZ3sDcEASMeJApzWGKzlCOhLMLpl
LSHQDibLJdwrDICk+PeMMZP/ueKK8MU5OhzxH0g1ZAD87v9kn98+Dna2S5Y31v+Pv7RKrf2nkKwV
YYe4Aed0qXLdSFhi8Rnn4A4/mYzEWGnbUC894JgE5NJ9z0IM0tuYWnxaef6R68QCIHoh3exDJEmc
3qRhl+oNRj01eIGvO2BQpaPjk0PyYKG23WK2/kGlekUuzmIVQQh9GRAkexT7AaWZJYboeixsPtHi
K/hOT019kBPO5GgLJ7VrfV2fqcDkmX2aI61aaqzY0FR2g1YXtfzFUUbI5D8kWd5jOwxou7czei4d
hz+RBcXIT+2grnkf9TLEvJaHe+KKaMOsbxuJL+awwvZZ7335c/yBsJ5p4savHiv+v0RPgnFL8pdv
opSnR9ztquyVnaED1y/MBvv67pK5oETYnRyFAYqcmLxNOrlZgJHwyqhsaC9HeTjWSXrDOD7nLDyW
sPrnVpppEzNOcolvbRsPRsCmis6JMfXzARnnZGizswvrdoNgW32lMVNdipIDLQveS7byLTTT2R28
O0D1U3Cr/Tb8BBbuS82+1QLagK9QlesFhrShAubbaLG/HYHayZ7q5RjxGgWEWTT9JUCl7FRQcIq3
o6rJhtrZhVr6uL0baUI9HBfRW+1aMFKf5D2qvCmTLLsE66kCKBynM98HanwWMFax2xhdoMbT6up0
yBHbJ0I4iNi5hVkVP2RRo5X9CkA7o45Qp9cEonWXbp2Z6dDFZ8a0TUK6YkzFcM6X/7VP+AFMB222
6tq8bKrd+qJDIwbz3i1yA2XEPPpgWWk7iDrW5H4j4SBKJYNbjNrZek28BBVOxCvyvRCtKJQMhEB5
bhcP34OhKcX5qP3T+Cwuk0m3IiW2V/Do3Tt8famnXN3/sgz3oiyH+gsyiMoFI5DMA+xG8VXMkOTJ
AlMq47HBAVYaaJ/xrDJdoTTuTkvsr+I/dE3v892q0669O8ZPH+2SotS9RJhvW8ji5VUnz2zSTPBQ
CQBuazsWb6EUTP4EIZqgusWSMkmMvBlpUAtmywn0vE5b+QL1n4CDXPWi6WHNN9lcaaO6AlGcQD94
YYguaopLUev9JKG9bVVaOuGDPAiPWV3JfAY3Xsbs2ps02opZf9wp+JzertIOQur1NgxkTz3NQpUN
pkE7EmlM0fOFW6GfBUGGsbTgm6ScNbY6RUY3L268zJwOduEhp74yFfHAv0PAmHNRqv1E4D6BLQdh
hRGTpW7pbTaOjDmCFzW2hYvyRVhxzCsUUTC1TjlcR256mXzypTxwQ+Xaz/z7eThnX1Y5PcIkSWLN
XORae/WmypQf4sG2MQPapgtG0O+vRNGelil81eXHaVxY492xf7uwJnDNKcwmBMlxUzBcG3svyN8j
FN0yHMIclnfgzR5OvYi5mHBBFW61rKfD4Zq+RqsU+I+oYjr3uZsV3qBhuRgoUpRXQJgiWCpnQUDe
t/XJdlebGbENQD/fi+x7Wf6qF1Hqb6WqkiatVOtOfBhsdVE0jknJmMAl2/hMvy0PnO2ZwoCtUL0x
tAThVcTUgA6+Ejw2fzpxYyLAHb5dYVJiskEZ7GxEsRtE08solQLHmx6xYH3XuhBfAg+Adt8ZWN+9
uDhhDtvlQQFtzofo/r1Q9YdNUid5rPy2TVi2Nlpu8yS5tO3JeyGFd33WjjrjnNxIHYzoaRazbOsv
inF9VnFKy78zTyP0bOcJhctFKfum4vVX/SIT/QNllqhvk8/N5SqQUDSrTMLQUcV0H/OL3grTW8J2
ekVOJVkqPOVarZb9zDznm1DTAK1VjoKTBKPisJ9UXEQq4Ic9hig9O9X2I8jh62Wav7DQv3AfW76K
DXQYmEhqlG81sVwAv6loCP3uP0kSSWzeWj3hMNFMFzLuEG2S4A3Pvczg1u9sn3ZmZYwyt0qVnyiT
oTzB2i7iozE+gTX+YFQ6vK9wZHL2huD8EszWv1Lf0BKGr/b9qCVTwHAXu93Y3b1iex0AccjwSltn
Kvw/Z/XLQFL2smulI9B2lE3eoD7IturOMmsnNZCGL3UDAZfSJkrY0mZ4LtXERoGW0ZHzHKUFU+It
qjldKGleDblZPbv7ghzoXxJThBaIAXDEL453WR3ZhX/xzGD/T8Y9+1eCJ7XA/lNJRUW2JNwzJwO1
rzpLumU8QUM8r+5yBeoHHZDP7OwGA/Ctaumf+LNO5FlnHWfm6LXWuH8JVEOl5JcJTw1tS/M/diTc
5qiLdJ8IndqXTYRsUbuMBBn1Bi319aDYQZ5kbwXVU3CuvbgdzHqhXbnrPknjJxZTSRF6iqJoYLwV
Vk1p+Klc5yB+/dKWdrg/HrGnYJlLjbvEkOg99flMQbM1oH+CG/QNifIZylTpZsjQkuMkPkBC3Sjy
e0a9BGvsDbfB/Pjwl1S2uRmItw5nPsA+QW4RFpol3qoxt+QOZPk7ZOFhrPDM8jTIJBpGwgyvvSW2
2MJX2SMz/3mmfl51gj1/OGEvn6147Vo/nQltmzexRxAQakylC/S8qWcO/AO7fbRIYwcIPCKIpEjv
MXNgA2Njy7bSooLTX09joMC/3HDB0v1TKKCuRi3rIroyz76S2hD49PwsWKrTf7As/1Wtl9AJc2LX
6oQseq7uJJvBMKbiCuJq94Xbi61rQh9oqPaEZ/EPUNTxSWRaQoDD57aKwOauGGaHQGNQUYTvbk1e
Y2GaMrj3fGi4lBZITXd+fcYNM0kNnKbvEmFMKZBAJvSt4Hgcan2FEM78VPtT0QMiNR4XugVJs+YZ
IVmZyO4Dp5gYSBoYxJLF5x74NDFWanTuLSxrl56t70CZB+QAcCMWOomJ1yw5oOScAImlgp0JRURj
DoSO08p/jrdBUeytX/OafJSegD9LEc8k0R+XqQREQJNO+joFKWZqAelES8kB6aIM1UlYRt656T61
HooaGVBe0fywJbK/e7hBCJzEPywrOwZkA7zg1N7TxUjndq1bqRbYAIApFYr+0qHWfBUmJ5XHjFJm
gi0LyhcugWP0vTIO6bIuIbZWL79J0ENUHCVotHgWsu44xNqG8n9UIAZEUukUEOUE0Yi4XoWykBDV
DG6V17xnbYQ7doCOkaiME2VPnqfwoJ114N4stLVyi7XXm4sfkSQtP9FTmRR3mLyDYUo7Oz3SutaT
Q75xZ27jGxD6cz5PqTBArkvcwOBWLAXQ5ISomCUrcwfrWA1m6nB0cHd4r9lIwKdxJ+pDftqkKPph
xhhljUg9d3IUoUIQvslaVoyYbq9goAwnYnowzg69cqFF3KNnful3AYV5lDOtaLL80YPu3CsOL2q+
11JwJCVgR+aqUiYcnk4fq9Ge2qJ7Glv7YiccXTbHKUTXIXe3fbyEsRqIWLOPXYD6ufaolYs1erhH
hYVThHiO9WJTyy8ElrHVK187kgfPjxZpf/kQOKpo7FgiEv3AGevRsPaR4kMrWvI8xcig1gNdeePW
cL8/TLndROEgr08+vwHGMYFvBiDsTyqVNFSXkvw6mKa7/MmR7JZMLz1bUACYW89k64/Jm6Ja33U+
nkZpOhWltXj9+Cfpy/I4rqfbKejQsg03YOaBoQ14SZO00e/PsU8WPZFofWle8FwrqQ8S4N1LNGLh
k+xu7q5yy41wLHAiRFDYabRoiv7ma9IYgJaujSzAEFQy4mDZ2/d5h41w5007Ef+K+7jh4fIpTiSL
tv1ImFAsmVfrfTp/O28hTmSScjkc6KHmIyyUzF33x/Jjr9UXzxpP+gFLEfPD7NS416kKCyQsmMa7
sQcqrw85T0CHu7c1KJY6WI7JW+3RBF9EkgX8qsTTXwqgFX3TB28tcqtBwPsTPOL09Coj/7TOdzDI
ncRkEPFpyQehAocsApvBwCPGNwLLBbIr+CkAugcLhcwT0yjZBppPjJ+WGael3iEGAwk87Syr/VQN
MBU8JNzFO0hhDmUL/VGb1nOoVLCMdu34l6KhwKoRKnDa+KJvhhv4qd7jO9UJzEE0rENnVCWteelP
j/SzMcGznqeeD0vGCZT8ptl5144vYvUJbkBMlBheGFxMYEJhNRgtwa4hS1Mh83suWNO10H92ehVS
aRbPC/+lJibqejbhSKOKCIp+J4zFQkloQd2mh22r4Y7vOstZ5Bdh/CfmAhHlupifDtXV+yIbFSDT
iy0tVxJ3/DvYCqVp5GNFv7xb2feP1l1LpUxqY0pT16/J4tOBnde0NfT8Nacgudzuk4ymkCvza+jX
3euepG4MSc8SzrMirf3uPY/cyHjEtHrkPu46H/5PIVavJx6BoE4a7gBJvBIPbb15DG6mFuHlesjv
w3ZQDdOIfGlVSZpL0hpDztqTZHCUpouYE+KMT2KCymbRjrvWlZ35LaB76UoukpgtVF6fZhMKy+vX
x9SdvL6SLD904M9oph3yw04zoVW6zI1nav+/Lvzsd2ZJyyvmm3TdktyeNCsz1HCAA+YJWv6TkFjX
CywSNCpzVvHgbOJhdksEHDA/j4dIXeXMWyGbVE3NF/i2K/o6SY2Hy8B7apMkS2xy8PVmWBoFuhR4
6XXu/Ysn5ilmjUGm5Hu+b6Grz7PCfpFSgZDbkzj7KWEcNuTQTPAuH1NC/BFqbcJ2/VdaBuRUfjzE
GgBzC39HfSJ69jJQIbUQKLjKg1ZI/a2RKYVEk49EbMkgZwxgAlru300LON9n3/inZurK+QZIPqaU
kSJ1KUQSxWMjW4W2GToy9vzS0qjz6XhBFJd11jc8X7eByvIjbxNurwk8QyNM7fzGltrI3c6FAX29
SSHf6AVlbT6+wBSxYO14RHAnnOND0oJw7mGxBj86OnRlsXb4jqUVJ6OZtYlGhLllfwV01lWueNdm
Si8t/cwRywfvxWsdaFHSNDlDmhehkpzQ/HGZZRaxQRtrlS4Vg5BFZWXyTk8y7WoObTWyUvwq32hP
iCEupE+QpH51jA4TU/biZTSDN5zC+OLkj61g0L201SCN0kE8FluDHYNet8/1IrUjuv3afWCBVP3W
OacFn4ONx2l3bBayA3dzNNpiYPgOjyFSMWek5aPNPmrmflMqimrK85WttT3v8hZUKduX5uRalZE0
aXMdNAmz0OFGB0n6UkF/qn8zJ3yoatHhzLoQ6zeuop7l8FQ+6qV5nE5OuLpPtkOj+VxTaC2wvXZX
Hk9kspEVNQGCZ9nvv9KtHQHu4tFeUWDMGkwOaAOzzBvU9Njxj4SPfSXKFh1j4SF1NIsJuG1qm7KK
FgHw7lDZU2v+7f40CKKkrGfzZ2NWtV2hLXSl7xrOQvtjiFxH93EDBKp6i08hrW1efAlZ1RnulopV
vh0yLQ5rdpIOfaYNImeJI4HEErW1QOnAfSawE/zshfsAYHoBC8Xn0uwpJ2k1nrv5PlgMZBlpJh+1
xSxzs1ZIAFv8v33CAnc+Nn/OK/XxWD964q8SyTWJVZBHabx9dzKiaimHNnNmGZ2veoXmuTlscyDY
bS4twMCBw1f9D0C+MCOxb6KwceSUulsfSeugYqs6lBeHDaDuedfcTpFPZOZADHiMEGcgZCYGzyJg
eOoadISlQAICMlixKJzrTl+BNXAgJiVPprlpVRh/q35llkG4D+8/FjJtaZqkYMmrUps9SaqA3qZW
SsXOZ/xyen3veKWiC8RCodrPCTLOhi1WyoEIrAtKlxf0e8NcPYmRX+9TZ68jh58GVdy7KfZLpN+3
iavREP6o3AAKdjCO0PKtJIunheFueHxnyzOarUgG7plEXgohdJWxedTpCytEXWyIwXe5BYzf+5tb
kKM/h3LzrHxfvSlgtQC9jRkHHo2nFQhkayyCdUD+5eFx1Gxvd1603eGCKtAFlK8pSWuslY3PQ1Qx
9pFx41yRDRs6c22OT9SCsvwHyWGmvxWTVsAe+mFXbvFYxM5xjh5PG1hq/FJUxjA5fbz/HeXRQXJA
vtlAXccfRMla75hNGWWy98+4Ji/k6wdsmzMsGS40G1apMucd4b7i734Mpkl279NYQjl1WAX4HCoe
aQUCYcUnfmGM2QYYjrByR5OdrFtBKNGKEcEk/Ul7xDuxyAiLzVuA53nTQ9fVXYtcOavopHa1dItz
LGcDAPZnJy2dffEg666cL7AsnXjITV5nBsOZyxejv+Zc37dFZHMwFXeIkwVXiCDCmkBDcszPRI80
HBgt6ABhK6mlP+WU7ZDSeuBc400P3zMpUyUCxVQ0yE7sag77NcbhvjCBE8gvZDczSeEIHMSPC9wF
vNK2IZYuQstxyPjQTFmXFb4+SKGkYEF+3PcAYRJoFJYM+Y1tfy7od66paEnlU90rC+c/eRdH3bfg
TtNO8glIq+TDkTsbxFWK0o4ooAveztiAsDz+zCu0C+dDhU5O3c1pjYOS0yj7oLbuIrN/CA+K0Ixz
Q7llwLSkDRcfyThavpGl+8f28eowM3ffh24nX2iJIxOHVB/jb3kaDooEHYi3ztmd2VRfHPiYLJjY
oeUT9N8MZXYnippZjIPTp2ATP2Dd80D7DON3dNFE1MAAeWEV89gekYvHpuB2HgQki5Cvs3pn/P62
p2sieNjdn84iXre+kcTj9lqKcGDDVZrQDhcxJ7Y2VFfUP4HRr1DHik9nCSe1dyjiWuIud3DVrSYO
Tx2WnDfHrFS7W50xcJvSshtkzK53opTPbEc48koGCE88WZLa5AWmVViNLybVUv6fsHo3waufIOBM
OLAMkSJO7zWsTpR+nGljjUuq10vUNfa57A5RZqFISG9yBJF0b51uAU8ZTPCK6YnivCrmE/V9+TvX
vDXi4y514ajLRVmmzxFRx1oo8GwJjp+qB7qssXTaB+Z33EEdFkXILdhgj/hzhK1p4nT6JwaaoMO1
kKdoUsc7hdW3ABhLKo7ZQTviWb+LHeRVKewrcGt0pb1Ol8Uik7eSQUhz3rsWHh46gyAyvSpS2eMX
5dR4LB6o2Ygh8rBfO/gGrK9Y1Z+9Hq0Pa893HkHuACL9xYQB8y2bqWmqLzKmVs79S2Sc1lUkXdde
y9Me3yxmsL1mOumN5SHdF0F+JSzfnr0iPnUZZljm4PaMBlux+qZW0p9bmNYn7bX5fOOt1gZKk2dP
OzbOuSXzDsNxoPwC05LlKDJosZ6qPYUE8rRcsTU44jx8WVhDHh6YEjvhjYMhRTx+YKq2LQe1wltc
3tibK6uB/oVlkom/TMN3CaVJgn+60ORQTcar1OCeuH36uuryFoTT2gF/2/l54G8Uu0hWMCNOwM/D
E7kYz4SXUkWTRmmLi+9FyfTi8IaQU+zqSXtBFkfkUjdthgdW4XN2YyklUjBYbMdfDFQAYw3zAozD
i4JtUlqh09sazA/53LyhGPW4eEHIClCkd7NiRPsl+MEHR4LhjEGdyOqmPpWNgb23yg38eSh76y+c
Z8SqRv+RwJhLRnFxMyzGm/eGOWaG50arRIHGmKhUqHdVN4kGkqoiCrnLt3ZyhCaG1hfA4cMmVj3J
CR0nr6dqgyd9i1ALWU2tXWJgcGOszuzCM1/mOtbDamxI9rf+1k/7Z6FKGVeGbMx09B+10TDCS+Hw
8a3sWMfNeBdhrg/oKQ7B9t4B85PlxufPzzTN5W4P+74vo2mmMxia5hGoqBFZyeMaf1pWuQyg5HT9
JJ84gWwxdYyOdYcXlhuoPwkRojuxhOVV5TTO6baOdtWnsjpfywLzZQHBeP+4Kq3yljF3+bWgKpiY
0ms1nMWBky9aCgmHgD6usFrCroPSE6oBHRoccpLwjl4BeXB1mSb0cw9ohqg6TT12d/CbLjRDEy1Q
DMmS4bsgXlY8U+jIyaQMs3BCOdC98xaVeXTVZBiHV09mUysIi47AA8gMdIx50odMMssnosy1/h0s
SDkdvPR5D5qfet3e4dxRDHbI6/Q7g/TLaQLKSXPtzuvk5B4zsoKxIZ0b0IjNFWqniR1qyb2Yv+Dr
EM3u7+ZlsMF53f8JvMEQMWlrR4hloN2aA+BLNazQX+4udwIh2nMq5iRuFAyplIH94rL0E6f46E+B
ig2vnL+rWSXYoJx/JNmC8D6zP1BpyxNTN17RiIw72FFlmY1UXIRYAgUcFBpLYfBbswbabmwfjZmE
P+Csrq7HHQvXzB+vjO/xViX8fHu7egR97/N4gieSn0fJGv37Nn0CYVoi/Z01mWtvULGxyKI2xsZZ
05NglMq5mSJGyHscu/bu0IxXM2ttjjwQyX1XA+lcMCu1l71rwN8T+CYTrX596HideGI83DaoxjCY
RBZ4n6p1FgVUHG/U1Lh0sXGx+JVbgGQCI3cTxXVSEHW/c0KLl7u0vrS09Acce64NLZZGKWaWmfcL
4JuUUzQLfKuVl3ZJzwNiaSHIpkwNKh2RV8hlM8SVXo7gVAZqREtT/LzGD4Lkg/f1+I26Zx6cUKwf
hPjavpWVJIIkCalmfu/eKdG8HqI6nxpyxPi0MlxS3agvTB2IVMCDdw5HKhDeqX5o6ib5J8OrAoXq
nvDZPolrEPciiuKk9ZTAVfIMqf3oVeg33wO4x3v2oiGigAXePaqXifOpEAC1FcFFebnr3cdTwjAf
flWIEo99qZnTLZbLo/vPF2GB1E7K8otSrnT22ugWuP/rZFP6U5AnJAGTriVjtu8eU3UQq87zka4P
p0onf6IOiszLWzLHcq57t21+B906KYeiw3Ut4bbLHrRbESze7dG21APyYDz0WPRNNvCkQmI27yQ4
XbHG6x9c+RPM99TzBnrenhLX8Od6nX1icraQTmSF0UMJq/zpRd225meeUZ17v0G5Ui/KSDh7qFhw
hetV+7txMoGJF/DkK0tlAHOWZO/1lf41GxChHPtsrV9NhlRQbKPhCcuiAjrpYSpWedZAeMuXl0/2
qFpj+57wlMhhltrcaAL2wxiHO2p6ED1JJECaWaf4WtElvanknKX9HTP/pXNvYijiztgNIgZ7aZK4
wsbxJKipgZuc2+cN5z6eWeqe0CEH9+MRx1XvftwSedCGP+MqIUsrmsMU3QiWZygrYN3uSs41U2jq
u4sqMJySS1eNxpGQ2uswy2liMEF1NbJX6uOTzP9fp5iIaeCGsjYNP1UaHuP/1TJ2hyVS4N5sXYkH
iwgeWvCwlo4sOK+0eTxQKQN9s3q9PuFES3BJKgwoV0HXmyb3Dl1bUnvCHAOQ3hVctirQtl2QsU5v
EONEfbAHnfVAsC9XqKxtd64glDZ1iXGDxZKEOF2UkEDMcEm0SVCGIsOLe7tdYXfFn+pm6Yln/NnU
8H5MZJtWhZbhP/T2d5YTB0zFQbasfUFQYe8Afq25O763r9QwOSz0fhbjSBWWOir6ip2zkLDhDmc4
YZ0kvXNAqLehPA3ymGyvWbsNBaNjxiMdKCMXgAtjBRJxlEIRD8WL6bxJ9oBRkRQvcV0u5MeoQUeL
5fFN6/Im8iQA2y2xj5+UFBwl5EgL+ENxyx/U0zVWl+eYIRs9owhTrnA3gLu9o6VRryn0WtgQE1K9
dlEYzp/gV25bgqcX7a2l2PH3+ESOsOmdL6d0Zwenq+Qov66gVN2Fgi2j/IVKzMdvnMFbHDSFpXTw
gTo/kfgoj6NyElDZDSdOq+cmTHmhbcD2ExOIERzrUtnaLLG2nSGKqC8I/8rsHw9AaMUBJ1h9YBNy
on9jqO7PdY3aUkedeeUrv7VUXiGVsAOBCuhWDeiNllYfPdVjS0f5s84tycfusX2oO31aYL/3bVrV
BI19QPoEOeajssqSwFePbfNaKoEhaMb5/y4av+UGZ5Ey43FEBu3yVSV/WnXtPAMxOQE8ZVVD2KW1
tSvvgYlXR8oV8uLLrA2vDkrZdq+mEcS1/u5rkNTfbtL0XM7rS+VkgbDJyMvNn4VXFUZUFTYWqqVp
HF3HtymZgyIqIAb3AhuCA8b1kl+e6MiSq8CuYMDgza1RbQmkIG4c108WhDuadDhcffixgk1N6171
bOSEm5B4r1pv7Wj1LXZuD7xSP1dnpjEhSR7ckCU/NT0yqCJXQcrE2dVt5ZCYsMiK2aQ59LSpbEz3
tnGLFioTn7kBt/BFITFQSe4sL6GiEGPvEtdfx9epVCU0mGDek6sNbwxrjzaXbVqSmXkUY6Nb8ujA
7PLJr2DN8QzqwiePaOJcsHVOSusZJlEu4jiKrskxXfUiEor0W37EKpVbzgFYLuc7l6TvTrYZT5CT
gW7ShXr0RaxbrNU6sy9xGvZSm0PtFzZpQ0z2xG0+Tmtg80skZNxc7A4KZZFDFgS8lvFeiUae5nuE
FYpPHgRdY7kVu2HLqjm8U7oWnG+27nm6H8fr6Ywoh1+vMFmzo8xr4J9+DAEsHsvWkSnGRSLWJmZI
EAfelsA2YYb1kegbsQrK5YpdvILrvG6E/2AxoQ6ecKVxK08bSnUmTOYXd8g/+2sXdWR43Ry/XYCs
GUv0h7LYse7U4Y6v5L2tnHfnPu2qCFElsRpPWKhYrbU/Bq1f/AoO9V0t0Q5t7GRxct2Q+5hMLird
iPFQW7UFELvW+KIrJtpKjhekCW2brN7CWKtbLl4+chWWL5t6hYYgkzIfnM6qph8NH2iG05wnE/+9
ZGVzsHdnTYryKiZzH+U4w+EjtvgIe/9hAfJaPqN6mX+9eSuqotcuE1NmPNgB6k8HaNlk1+hjuJ71
b3jKzykne6HmITKVlS3m8EjmTtzF7dvUjnCV+fCOrCS69ur48f1TbP1stAKNg1vjbPlXyruMYDg4
YMNxad/siqyFvdvq6fCF4nznya1K/85vebMOyY7iU4CQeXVE4qgixoh5kyNtiVUzNIoIWLnx3QkK
X/x0dRT++7D5/dY6O7I+oLsFMEWRX5dVYyycov78AMw8X/Xei8DCzbCoGr5CYhL4j7X3bWp5Xk5z
rcHJC8wwdkkjCe+ZMZlrhQ+LwgEkSFD+KsRTy52ENhwl+XAFJ6uYd9WykRGEcvvMpmN+/HXpFwH6
5ogzD0tZLbCFjl77wTUtIBZ7cIVuYWCYb5nXSsSyVT04U4pnd+0xxb2jPbx2/BJ4kdG7hHFyxaND
xUZ3e7EDzHPNQ0IZhAWYgK0FHPxcOiAUARbL6VhFzzddDQeHq0vRaJQ/0mNaBqLMlHg/PDWAvTf0
+y11RtBKmXSVQ0OZJERD/qWkZQnV8J/6c9cBqVQaoUQymSxFDxhiGImJzeI77TbwQuxWlMBCH2Fo
3fD2Ejxj/o/hlytkk6qeGoQ0SKdYKhgoK+5s2JsoLIo/Ah4am4DnMXlGUOT/Z5YBf3ko3ZUaROXg
eapOD45T1rKRwX0wNxod37DRsZZ6mF9C5IZOAopXuseuejWCkk0fnkev5ukjta8H0YjiIQMchc10
1NE5SsKnrQ2o1d6zVhDCqwtYzjOpa5ojg/nhnYvVcvoYn9Q7mc2sUt+lYzpYFVTSPWeGQTSjyT0y
eiliAuMNXs+lvBUVGB9biZdh28S/LG2QdPZZLN7tyeFH8kQ9bctF1g359oKyaLynsvm0Vh5VnAqk
t7/C8X5uqryFjlu2ulaJC3JzZ8Y8eOHhP082QKRY/NoG6vrYo2Rrdd0ZFckqjeNNreI+R/Tml6rl
Ney7Sb2/3cR4hQr2gRAMqiGKf55GX0VVM2x/HUcJaaqei6xlUUchzVUMWojzrujJyfc3HStA3ZmW
tluMdy5MEs+xZ3LnQ/lToCWxqBRd5JesBVsh+lYyP1c+f9KbMIVQn+/1YNruzBM9ldghE27F7+Uf
0Z6IseTl9Y6o51kyTzB3lbZ7JCdwr4bf8Z97ofl6OCsWPB0xTKIil1mHodtOdma0zsNZyyoSUljW
NZBfw/pdxZiSdR3TJgiIZVFPybvAYyUSDpioihLCY1CcFXbxtZg216ZcGlUoAJWTZ5F0nB5mX+CZ
izHfQMgQAzdZS9rUGFE+1XjryzCHisLKwZfsOOCuvn7uS4SGyBuATCy0oqxAoQyLYJH6YLdJA18J
pZlLtnjQN96T7n3ErLhE0aFIJ1t6+mwnj2Wchxb+qas3TNBrlZJHspkYvV/jsFnDBS+Xc6SdtgEx
pLjQmLgGIzg4LgK6jfFjvY1W15AzNHMsLp37/Lwh7VDrcBRCBNBAU1wC2mCi32w8q+f0aM9pL2kH
3YtaGFfbsA0kDHpY+gLSS0zE018XzVwnO148O7+et/V6UVjT1fMAcdRx3w9K/9a1IBWjLzTZjWNz
vfH0SfWfUKNWgIdQ2TMsF806RlKWccGyJSMTUV5UEEBImvggHjY5zMCfjasY9hYcRZNXm3Oe9+aD
EonwqnGWkgxTyCidW65o71DWPtWiaVRRkU5agO7u9O3XBdeg4kMKOEQOGxHZvOsHW8nx3+0U/isE
nZgcmaLyp5Uh38t20Hzl7bOT70sOOdQmlgOjZRtc/zMOPkw7cwSQtA1wLodmaGPxauDPEc8Cft+e
PEQlxo78EbFY2Bn+4Yq9OR/78Fy0GruOh3gmZuvYRu2BmqFJv5DFyqL2GtlqqaS3sNhKhDycympn
fdq7cjkZmK0gHxZx7mC/zXT0uC6MFY+3ke4cGcHYJevi5nUk+awtRXLWtr1dd3BBQQn/3+QRjVpb
cZ/Mh0+clbrNwgl/QiOthAATkq4WnbJaexUT0wIbxmmJx9TF6/wYiI2pHQXQqUFsYCySdL24hLXP
6Xtky97vqUTGur+NauMQpT6/fm37b5a0r5Ev4H1knzE1SNfp/SwPolR4X58SJrcF7Yy+eczlYyeW
+xyQvKU1gsVpC1HGdnBqxuqXlqPCna3UHMmXAo83N7gP48FfCrGqu6rTNymj9aFuobfnNUsDQe8K
Tgnnb5bGCeIBNDEFGuUbpWkbOMRvdUM+U/YF6ndrlXF2myNRnwxUU/aa8O8nXM7yzXVmL9l6FsHC
CEnlhdVUQ5oFTakMGOZNJmulmBEPqVeK1G/2n1XQYM73l3SvovEMz+vjf2HU0sgfqOIPmJ9HqnDv
bsGtfg0ByVz0BShuimXitzoITf3GsNVqynSRCu5o7cXpi23C8ahD94AWW6IpvPqwUnNXnfLidCvS
/q4XBFtWnYwTH4UkFqSIkbKw6Y3vUbVH+Z1EVGUFAV91Owpzh14MDeyzTE4ostK2b7b7QmpdvPjU
vIDgK9rS6KvU78xW1WNBWby3VqO4S6n2hijxKVSP7EVwag3lKzkXEBAvhvtH6h8pSRHABrPsLWMd
YJTM2HPv3mf4R9WyYHfHOaw5wpL3aDik7KUzlB/DYRiAdlrhf2a4DHqSLd/rkw/qRlG00kLQRu7J
aRP9NfpEOiOgqQ5Q+w0WwKiN9M66PoLnwoD1ix7oSsdzjZKtoQowHSE9Vigj2avMGMdiUCPXbk22
d6XbKkBvnYrn8aLOdtSeRt19vlKbGnK2yHfTy0ySkKwoN3FpD/SooON2J+hEnl7o9LkSV4GVI4Gj
fCGx0j6YHq7KhD88msxqdSf6qfiFs0LLV+1JjKwimHgNNbnwqUX6fzUp56S9AoBGeE91KLb5h7Vs
kAGmzP12DMVNI9qWIHhRV8NXumXKeeU5gRNoylBs6hz9YeNiOC2yFYVDvtZLHWiTvyiJ/8mMIuVR
v6tzuMpwFCMjY8P9BgYoAjGRw82do6WAIb8QCTOI8Rqv0ALLVxPuYf2iZVrNVgkc3OSGsZ3Jct3o
SiFdYgxsyomj/8mseL/N9Pjah4NYMBR3zHVfKkVk4mURH+0TRojjSrJrE2lVWhidY53w7am/ZNrG
gt/Z3J6NvBqBIH70y21lTVYZ+FBQf+/yOqyQX4M+lvrX5EtnNA9MiIltD1bgUj3mVQMd68kWsZVd
0/YQb/7H71uEhyS0rzlLgZLSoqtPCX8Q4hX1fpsqL46zpaGtb11+OGYCo2VsSs5C3E7j8dL7kHVH
UmDV65DUgRvijISI4BHcNiHpEYp2k5POjr1dY5xv0cjrJ1IOevKbIKda3U3zcEUXHESAAeCCYLX4
zcqXkdctgl6lcz72b10lEi54AcMqM9PbNpVuaXuwu7ZXeLyYy8I940fyuFCWgtxDyjblUJARA12x
FKdVkjWElLUXvAe+z4klUwzlcehVF7Ha1/EigreXcy3MgYt5Fh1Kqiei0kgITIWe00jerjnVoKQ3
0NB56+FqqeJPRiACr7mUWakuYjQqZ0p2V3nbGjVc02lkNkyertTanlM1gnrL1RcJc2dn2Ja3CO/d
XUtXUWy3cXOMN+6//6iOLsCP4G+BLo+y0N5cj2eF1ROoheSocHCXmEG6Mp4uH66c2Qz/utz4enVJ
yLCapZZ8Ew27HnkbEbjHFGPe+0P/G08m+8osxPJMzc7ifef9FDug6xpGPmMPVl4bP7G064yejeMq
hCLg0OvTh6M2+Zbw20cgdc0Pfaox9/XtSLU/m7IvT5clsCezg4NvscJWRCRGU6ZXQ4G1aF/z93CQ
hqVF7tkakyIR2UADDkVtJNB0HGyldysnR7drWzrcELuCJ1rvWIrS/VpPNyVfnHUx9vNeduLXbzuR
40Jrp8y1BCgflfuuoNwo/x7b2Qd4IFPRkaxb/M7oncWOXoCohylthVhWFeOyxnh+T2LsCpr3hmqX
SzkzHwE0Nc2LzCzrqqYPxceEd3IgcyY793bM7nEfCGXJnwuTJtMqUWUazrUfJaYADNdsY16vv5ac
KfYKJ/fxHedblq6ETu7Q2V+ZiS4J4uAr4lojOYagipy0GgzVwuiYCgvLUhyL8KcfN5f6546if437
FuThxO9BG1zZAoO/10NNF8/oOj9MWsCcUY8NbRFWqS16ZexgRfqmv7VDcRLd+tuARkkMxuUZ1QcZ
Ga5wIUZKqe4qwEbLlUCYhDgOFvX6eX034tZbBTpJro12wS0VkWlhC5dhGObIEuYlpVkGMWIzVv5S
iyewJF6fgkf2qSztvA/2X/NTv4kv740RUvhNFMF4bNIXyiWmIq6hBAoRjK9jHc4YOjV1CbMo5nwp
4AUCPgzH+zCceko53a7zgo02NVUwl2Euf+fhIycbwAyXPyMZCqNQHP0l/LvyMKxOgMwI4kIVaoDd
Ca1LbCxufs2a01jeTxp8eWHE4NYOVh1gjxhKsljzLQd9c0xjRdnYV43ymW+nJ1Zw2QS2yY3L4nW1
jz3Rec90zi4CogPIY8kXC42FFqap1dwdU7TU6E7ZxpaJOCumo1PgLCgnuLgjL3uaFxeaCns/C4Lq
R1q1FZAZYkSnfs79H6fsGOovUNuEIe0CSOE4REHzZzinnDK3G1cLyXbgLH35DQAGgKbqIJXbMKOR
dAUV/YfFFenO9FTnbQk7WKopC0wqCMh9KBjqmBi9tVEBjckN6Lw2VtjCDJUBbDryFc/Zk/rDkTDa
HqYIvLrlCCkBS3kda9g+uqNQrPh+NlCvy+jerE0TibXmJvWXiedEzu4tbaAA9mMFIWnz36Hvol6V
Rz7xu0a9vsYYOFTY6fFeZeaf4y6SrjPrlN5l4NY46Omvrdab6EuA867sVL4KmUA0Ek0J8s1610HY
jSkmW3nEEhnoepIH3pD2vJfAYja0CHDb+Qt2lT/TyM2a7l4zR8EY4me9Eklph+8zC3xDUzUyQs7v
02DveinIQL2NOql3uqF14195zedf8Q8S+w0ueZMBlH8160nZ37pfwnuzwACVQnyAkeCp5I7BOyPz
nTao7IBcYkCNKaZVCHoE9D3W4cH1TTybgVu8FNceME/H3UVJUBI6J5XBOaQq4kXqaWxwqCdpuSsN
W2TWGJlajDp/jzSfITo7dpmSNPjGnCX6fCvolXTowZin7y5OreGuqTcYZSF9DDKCfinkQFLSHz6Z
mT50OobEmLpyjlLCeTWL1t7h/4gKbiWMLZZHAcMnCP7hptCrslJ8G70bjWA6RtF/kPXHDiVV43FJ
lwCfGGBtpZel9cecw7LtOwmAjpJBmvDl2sdwqb8sC6fnTbIFlOpzhX9N9vEww5AfWKaxmQB0s7cJ
7ACafompI9u9Q6pK4yKly7m2mV5Ydepf84NtZ+rbrSPGLUZuCp8MrCCjNqP39cAeV+ngwticZd4r
iFWmiMluWewdotJNN+t0WNFCcPo5a4Rske79nVdgxrd1pncEhwDihhKbkWWO9vNMdDZHfIr/0Xmf
xyUWe00gIYKtIwSIknEcTQRKbG34y7MsmeaySzLxYxtOoCo5pBHJktD+lMQHiNrf3HWG59nQK5y5
4xBHYtLVW8TOOFMmedBvle8//IzjSUK5IB2oMb8/0onbTCYQtxp6kJHWD7xlxqN96V3LLbOL/Pwj
Q5itZ/ct8TrWDxj95t44PVQtqse+wlENDivDJfa/jqg04zU6IZ5p0cZUkGsrrpqYRbIz63Dhnn84
eyhPwT6ALtiPtpiMbDO/MFQrM+p/hwSUyisGCR4IrVYHfx7AGbXMVWYeXCVsX547fM1sRtgcjYaE
kq18bXMTeMc2ZdiCfLpLS5d8jPhADK4uPrbKdSh4XFJ0GnLxHkfUoOlDWvwSeUpmgjTd7Kd5TG9D
NvoCB3qSprmguSS0lrpkANwFGgjWrx28gMUezCiK31KW5gyWP7ra/zDMCwVyq3WeeNJJjAQsHh9E
WNEBTM2kTPefXabwXukuEjZNFj0c7wDdRxnm9lv/Be6tL620RiUO7PXsBQ4nwCg9IJ42Xu75m6wG
Up/RVJKgJM6JHBOdrVEGtXnQHffHxbZsXW5l62k5euJ+58MZXn8JPTwNs+PNEr9f/xM6SykiTFZG
T/vOQFkjViJLhxiElskdLkndt+zTDwO5Z+Pr39hB7AQLOTUzLx/LRe6JZmp45q3Ijftd33GpteOZ
UQz7vJ+rtpiSDHxdpe4XlNipjvoQ2LmqCjnbtqS39UcauKeplEsQ4JeXqFbzgTdZ8Loq09OQAFrG
ScKFdpe40jXBSAjavHhx6sRyWXIh5dG9COTjZxFEqqpBePffB4NrMC9KC+NyVt5nCuVRgJLP1BQR
6kOJm6lYgiBqyfSGE8Qh6JUm5A/FyB3wpbVxjCu91gIpGnX6v4qjpP0zoOyo4Ln9A3aebPox0AU9
idWTLbMaNDq6yPaj8iWu31vR+x7Et8sO/u/RJCxuJyxs4sjNrDfNSgZ0x7UJP2kEaeKQFozQY4gc
QhtzZ0NimJ4i4h+iV9a+f+uII2jHBrlkj0xh5gpZkXsjOLUTX2ziIlji3XvBTtdw8mT+BPI8TKcV
9FOHDSpcwkA5WRO9bZXP3S4RYOEEZVUO1BgUnhcK3qgQjEuaJAoobcR2THWPKxQAg+Jfi+lx9VCo
vJ/mda6ne7rJ2FVd9MGxfaNOO4oxVxEUoMuFy4fVf9pm8VPSxleOVQhHzxMOoUmmYdv9vbdZw7V6
E+6F9esTJfE5lduuFx4Fwdn4a+LmR/+8rEonQ4wRmnw/2Beq2yfe5Cel0+iFKRymIeRFk7tGIdgA
nmmAQ3JSvuIKL9KkkVaycma1zmt0YSyb9XBUvX+VNQ7c8u6RDMdXU9vhLcIfgH5LkbjJUvikc41Z
g6vWDc5jANuLtnulPvbzgGOlC/yTwMQoonFPl88f9SOZX4y8ZMmrQNVVUGG3gfPHmKdHMS/EIAyX
WvHx9a9jJ4/v1idRW1OqCXfzEH3J6+6TbagX7+Ufaahobh6mtt+Z6wU3McoHTRAcTplzFE/qOA8h
T3nZYIAEOvur2UQWbs2qM2Y6hyMOpTbYuXj8xI3JX7mciLBluDMm3btFCs+35JTciy0PfwGjJSac
HGM01CkDORdXqGtcf8a7zIrEkuiH314Yq729oqSYXZr3fPQhsICzXtD+hXG8bLKVgNnfIgr57kHh
JZwV3/FrU/a1Ew3E/UUC1OBrtG3mPvkEaUJ4NyIGf9DDqu0bAYyLmnzJ2wey8InS5K/0FQk7lvd6
6rsTpow0yfwd3LnN4U0EEVcBdawa9YE7YXi6T2MZdEIiOANebpa106So5LfJqngCKNGP/kfMrzP4
ELUntyQqCojs+WgUfKmH7tSoGHXJNbAZvCWNJKWj8GX/bantVUz9MZfAW9qgp3l0kzbIqdyDDATG
gpaA09q1mBKe228K8aY23uNK1X1pojOOacFw4DelAsjZFfXXcnFH+BgqwMvZRAwG9Z0+70JmKvWo
GdKbXYfMwTu3FTcgrM3DVi8ACpYrA57lCzuLXWluxzjq7i5Ia/V1SY7zLZCyRwYOxJHApqkWtuOF
Aqed1i0f1rrNBySWXbFFzaBrlPnm/yKHMLP9Eny526QXZ+LQqPf9eHp2MYZ12Dqnr7qYV5/Th3Wd
m8gH1LoZkwHJyDDGW/CvIEKb5/GeptdfRS3TNQn+RwFqlJdzD1VjGc/EiMPIxYGlPp6ckVnvFfRr
31AyRx20CHOtNdwIqeu050LS9XwhJdfxvvMS+iJKA8wJak5OyMqIcvrzXFfnWLHmheR9Q/Q6rWmI
E1KCOOyDmg6s5KTjLLo9uXDupsC+aQ7NS2Lo+V7A0SEsJz3kL75QkPS1RyKN2Uw8yHuLUJ10YIrK
QUIyW2oAuURTgBT7dt50iybOM4SRU/hfzUWhpMGGsFOOlDlJjrH8jYUvgR/+B/LKOBh7+FevqnH1
wbKeP1CiwbMSpVvsqa52eqfbFXcZX94RJ5GS3E4vemwSR1wnthG2FV2XKaZDOLCBg8qjax+FnY8D
8NEPkufGUeaxaPTtXTu9PGa0E78skMj0Pj+HhKMhBYdO3WX6t4sx061d+GjR2UssHx3C+D1A7NVG
dzwa3qnfJ8AkxVSPbah5HvZw4Ag2ORyjglXciKaAKBnk5dmSbQU7M18CN5ktuvNmfpGMfPQVrgVY
hqvj7H3YkrIGLw4LQjwApqxpL5p9T1bOdfuogq5Wh/rh5qgRzEp3d/9MpE/kctktp8GS6zQ9Q/ih
38h5x6ITjd7UOIK8Yz0CG7qiDIv8qZU6eONRzF8RsMmLua9OxoE2k+356QE7mDTy/9q0HT3T6Smm
NQCDbJYfC7QQjY/E7p7aRyv7+j17CcLONJWJuhcMY0Btrq+Xb/pDpAshfnUAK9Abc7Ekhh41oOE6
gXZ0hbZ8tJc0gwtHefBPOzbjNyX3LufD69eClndU1mBJbWXQrSH6C/qaDcTonhfOxmcEFSEfuwOv
mj52FsUIFNRQpAErKm+WKUqRVp5sJGA5QE0nbekMR/Hmj16DWLDrg3leX5mTiKxVbIVbCtHCW+x5
5DX7WYBbOZ1UDSuw0zGFZYaQ6RKm2EJr6kKis3FySP4TofLZOpX83/0OTbXgWguABDJv7gxxGTh3
VMc6o1Vinpkt+Q1fHhQQZK5rhAi8014Bm7kdNrRPa25pU6y9CVFrVXcrZFhbUd9TvhIlJQKXa0Gt
VT8f2OV1noiaetbgzqOWGljvp/I3DAza4RN5t22pNJcWu6ReRfM9HbDYisOMFivzrHjJOtlkDgqp
wGZB7caAUE1CrhS8LrT0P0aLfl4FgXBLkHCl5Z/vQIXzmxMnNGya0fZGSp6GLrn2oIsNo/UuVOqM
uhVGNn4j3a3G1eFHGp40+41W6Wdf6F6jGnD3MBoPxJS7rZmZ2UaEmEpf91+glDro9QQ0pm2BBDoR
cRxRo0p8YGa+MESh1CjawQsKdi+X9pI9zEC/CnQJeG0I27rSbhwJ1UfV1aku8HwQwIYdnBU3TSOr
8G1jfFYdQgqUuw+A5zFbdeuhlKJoGwf7xJL/OQv3itNHcU3oExwiLCv7vl9GF5sXNOE28+txbiVB
Bm3DWCZFHzLt3f4GJOxfpx/hrzK5O/xbPxnv1NtPuye6FLC7NH8T/yB6HALnvoD2KGZ5JTKum6c/
KoYwKASXW2FlmnQJqJTGqqHbLEDqBAMTh+fvgJ5GELF4KOv7mq6ftmXOiBMk8HmDhSZqTOrzSY7A
r0w33cUQIAaldUcNTIzaXK5rthXWuRSgrtvHhSacuy469ugU+yljcQWOgvAOlgvQz0g5tSPCLDN5
pqPf18jPGzwCgpr2TIy12fsAHGw2hFy7Zbc2uh0XrTUE06NF4M8XB3Dn71Tpv5oKyOu9OHvQ/1MT
7cHfkiBs4BbtKTwKbXWzu4Fa7B0u4OrL1YGF70sIQrBx005qLKGN1zqTycVzDhLDVTrcvQ/Hgk6T
pxMLcyUTMb8HdDg7Fv0w523IKBkRqKd3dEDCdjftusgHbRnjxuV7yL+tCHtdZU6hfD2O708SUHjf
3jMTR0W2gd/1xj3MJfBLANX97Ik5EXMPIAp8br2rra/KS2EqFN78bzr3JvO1aKnPEUHlTfBj/GYn
o6wMoLFti38ohnkDx2LGPlWxFOQHUIMoOuAUefAzvF5moTDHTqojbcqtaS0O9nhi2AEd/GqV7sW/
5UQrtjHxWQTlfVfrzdCXRBaBMt2IbjAPa+qOxHJXIJ6cmsOfRlb79rXZaSYZQlZjQG2f41RLAH5X
VgKjZc2a5zl3CcBPLYrrfRQ6LRwWvVqKg0EfZDbg/OHGn60rgfFbFv9TU8dNhEERO7QiyPC23bJA
VeOZSKBFZWCNdsLWLr1P/fop4Aat9NpYQRXfZ4YHtbOakSK07Qaikznh9kLtcGGKwr00q1y02YGE
pbs69vSLXprrkb6mgtP1tJOlYCHva372Q94H0XlulU16vLh8WGxlAlOMekffGOHGD0yhOi5GHq2y
hqUlGgTbSEDuwdWjsHStHOHPkLeekX4m7e3AuNa6EU1BOTrKK0FTyPp0fpZ72lmiAFFFH96qWt9q
8aw+F+UxvPn1WA+wbwjsdboMfSVdfvz6aiD50ULo8+Lwf+HcIMdZSj9GfdlZAWMqLbr/Mj+LfcwF
hzzAJZzGS/qS+Lj36He93Fbbb5xn6wS5nYNu7XNLdhFHWkv8MkME9J2gpxueLTB+EEe/00JTryUw
oXNg2U/8ts8B5tVys5isgOjMABE/l2dtj8P6JGwHu7SA0o4oLo3VD6qCyfIkbSAWo9aOCcwywRaq
Ya9dlgPLHaCiyeipbcaaHVVnpQqSUAEtJg9c5DGr8PElWxRJZB5WvqJ1GfZA+e3zxQE40dQmymHm
9M5Oy8l8EzgM6WoepLnVZ4+YQab3JTwdsat5s8HjFhOSUufVFrbj2MZR7VV3+NV8f2TBUeerh/qF
tVMgRE0o54xIvshs1uLB/FYo1V7h0/nBKfyQD4KPRH85bPsyRNonnELzUDkO2YT/Fp6NIvfjTBLc
8pPH+hPUbdROhIf+0VuV0zVojTVrFmDw/J0/JLBjwi1Rmge4nnT00kjAA1FtQ1Cfy6WlfQ/7H+01
fLiyT9VHwOyQeJ+wapRYx0ofyAV96EhCuoJB5U+kJYLLX0AXvE1zUakFahzlUMgSD5Gcfc673Bvo
IeUSwkqmOytIRR3eRklsIekW1qA8U4RQ/QYh6gt3zGBmLLFIKUUkylYPwDL1yhVbygBuauVS8zOz
Gi/MtkYoB0qTAk8eb2b6w1nmTcA5AmADtfHw0FJ4XOhXnNykx7KC1nnP9uI2UBI/3u/LXHkhtN1o
orM/dxRnpM8F+s8iXB1aAz039eqJXTRKqSJ4OuiohstIJ/nyrif/N5bo0EIaJ2JdbH/148QL7xg3
GWBZ0Nox/kHwg9ZAMcrKdd2ADzXPHWKeiSpZbCoI9/O0J41Ojn3K5hZr0mfHV3wVbXUCSKBt+pf5
h0qDtUAEwMbaJs2o+LVS5+U70gL7hk1XJ1qwvMvlorWtCJHMWJK/+V23vqHpkZnhCpeGgvTtHVqZ
xCFs4mqcCGYE85W+ArvcaNmrWJrKh8TV4NlcXZjZmOyCE73xIelyM5nKf88qdAEV6oZQiDr+vN5w
FB/Gcp3jgd9OyhnW9B3xmYHURuui3faIquFba8Z/lLhx3DYm1nM7sLrMui9Uws8UGVGI2c2t/cW6
KPJmYdFhHig16z47L7pkqTIPuZI+D0BeI3w+VBcuYKt12F8sxXgCUNs/0sqLlmdds05MvzTXzt7y
9E0n2UofXSe54hR/k4zHZ0R00K8M5bn/up4nPi9TAO9RyOK88DzX2BaZbfJfNn9tQNW0XuUpJ6ci
Zx68FObr4Df91BEPF2R80EPMUo1yD7IAPMLukQv4CvzJJDAWmYDAA1a4aISazMvuvV+u32XVyNDi
8d5Bt41dW9E/cf3wn5lrLeRdMXEyYFsrOTscH78kL4fPUNzvf4ZH/vJoPhi227YG9e1MFDiwtPU+
nwqwEsMcKV9IjuqS2+3q015HASlVyBOIYmCqndX8qGzl9GPqi2V08H+O9g6EZcYlJtvGBVTWkKZO
AxI3TyjBKy4goFhJL2ZUsb5TBzJK0QmcYTuEA7WXYlOA1N39imB4OzyX57ryv0jhFIgcMfo7LKTN
Ij4tucvydCYCuVTvY+BgG3k0m6ITxDHtlVMzdG1qrVcAfRP0doCIf6nw7EFCt+zP1yq/xRvFuD0x
6jUFNNJ1o0Uj7bZdtxOJYz76brwuF2U27RmxesBa6Xx5AphB71l0jhZ+HzkVE5yBHNsdPBu0TZHk
+0uACyY95rDhp9I+QcA+aSTyGMfVITvMtR+3ek5z9TzQZk3xYYYo6YQHxyK4J5/CI4s/CWu0eLPe
g+X0zIN/obeGPw0gz3yo6BzrlgAWwGcoYBzH6sv0X75uEhMVOfy3DUDzv3TxsRH/LXbJt1T1n70Y
+GKr17NsZ7eUQ3Slod4iQidHA79kuLth2XZiBrgvRiZ8KhzZiYtQbsOmApfQOjEdfglm7huOi6c1
VALVMVWHWMwykLUrCsL8SMQjvVSrl/rGQiE4gmNTKAA77506/SXYyAlR3gFowAa8fxle+e18ker4
7box1nFG3fYW9zC6svgjZtt1PPFEfI1dFSONMlubkKOmdzoLaAP2Wom7fTrPRtDaDd9FH3Kz0pP/
b4zVz42eD8nw4MAKLxKH8WV1P04gTpIy4PyjIzVwjDFgmpGvRdeGKNrUCUjwHjv6fw5oiM1LM1Ky
1pNHYi3ZWFkRgWqZGahF014WbnV0aWvQJTM6vMNat+enQNHxzONdzGh/K6JPW/U2w3znlzPTEBY2
xS1wXvObqDkNkK9QG5PezVIk5gs6Nb57Y+tVyMNWAHEA0ba72eck6XYHSTIgChFXg4RxeJq+hc3W
2WDTmmmFtpaYExGU/pZ/5mfYIFbTcdQSX2HuIMQhMSR8F8i2Ntiapw6RzTqOpTrkxUtqFPCpxFxu
VY9M5zsFBybkMBY78GbHNxTwMnuz2xxaiuOA0WlZdYNhJqzMhf9kBkvl1S+xzRQxWb20CqfsEaoQ
VWmlIT1Zff8SaflPPUeylceryQcQOPIUAvyooZkExIS6OChZXuYk34NEX/wsEhaYWVZxSLhE2f4q
02QWHAC6r1ThNqCakpuQLZ2BNMaYp9wXcb/q6vfOuDbEXjKyK743buIvAYjRuSXsfQ/hEhtwUWO9
uQQyPqjnd4CWy7D3GP1HktPsPHj9rNopt+yO2XP8KUyVRZFStFJv6DEDW0JACwl5xLUD2lkTaTm2
VzPDesnsn+A+Jsn9Xr90Vkgh+27h69BTtL2IqcUwfbj/3l7uB0Xgc4+whCAHTpt4HXg+vUgIx8fT
uGIW4SnU/7fZz5Ktu22n7QYjKhvynpvd86dmArUQlMW+k87qHShoXtzYtWvusVgWTJ61cBhlimzW
sLLd/zGoW9mp2+ZgRL5/kyWt56EFod6GIAcPQiZC9OmZxh8DNtzR7J+z95Dj51oEEl+NzCSlaGED
+v7sKeNdavETArsmFuzrEE9Vy+IiXwIWGs78t2XnL7K6cfp9VgA6+PoVIrFaKUQn1FJ55Dfc5ds+
ElMCdzL+55zsqtY1iJNGEN7HsdmlUGyWoWedZAp+lU0hLJP/3LIbqlNUjtCSFZliMrKEffPk5RPF
a1rwaNYhUSqbNP0RsPTPvfeaDOFNb9lzAttB657Oj9GjDzRdi2j6+cai5FuO9ycCKrGsaKXXnAHR
YTfSL/BemF9zagtchs97fp4zSoJmhr42gLXXqbJ3R6k1/07wBnv/P626yQxHCtKXnXBA25RDYf3b
JVGSIAJkdI5qXrK+oOnOlDuHb7YmAELIBBIEKSh1dlm/sk35h8npO8muNTd9stGGUuMOWFPdqK7A
TcjSpJuJcVBg78l2EZhI+EGW6dEGxwt/JvLhHm1974HaLfrXuFGMppUGBuek21p6PnMhDuY2Sfwy
00HaM0yQirrYYOC/TRc0ZSSEVcBilva62hSIzwD6kvXRZLKFYs/u4iMO6ZbfwzXBNinvZEh8L4RB
3Qoc6630N+LlFnvuBG60K87IlBp7sNFs9z5RaETxa8/DcWIFbJP02yJR3qianBYBrhEp99j2luXW
mo5LUbwe0tstKiSHEJA/NTGjpm4ba5nbNKOnbC7yqwhtZy6zZXSIAsGB7yERv1BsENhtci0VekRT
V4Trft+sshmD8oXdXQXonWkEHSjSu5E23q0rmIz2bpwfSvpZunToVkpJaja5417Rd+crJfdtP/Ts
WuUVKRIInKYHHsoVUoPv+aR+baeVFYENtvNVvXahFLPV68SiHzjG/9/V0pzesNadh3+DIJj75VUZ
UiftgZ34vI+nfk51nDH5QoE8eP8pXFVEYVKX8yX2ZbmcoxUYbMuzKuIawXYmS7aVAu5RlaqX7eOo
a43S2DSrgwdiEYDw9xqW3moqGJPCHJ9p6aSwFalsUi739k9GUf2JtbMF6orEbbQbnhzmnXOwhROX
8kxrW8hYcL+bSKXBzD2apOztA46ltp872v87Ls2b+wnJ1KOdvHrUAzFA4Baxn2NQHyQOH+zLSk4V
SMXJKL0m7xLsVQT284fQ6c957sMz77AfAV/0DWlmfBdVoPWDfPfsEi8oFtaCc052X8Lv/gAQCK3U
wz9iaeMaGiK9Xtes6QiFBBnm7/gEOnttheWK5YKzMIrb5G64DpmlLPGm3m+BhJyPvsMPeW1DKT6h
1FWuFc+gru73gXSOta9Dx3fhpwtXJi+6lTONU596sstrwI7FNcsblO6X07e6ycLrtXVY75NNy0QS
fgbNzXrlY34TmmaLsKp/dzADS3mvOrvMV7ydEHeUl5QWwQi01OF7vBdLN7HuHR4bf+Nt1tWTEoiA
hou+eFXKoVBZLwvuXQ8Uu2sP0YdFSmdqmpsu7mPtAbLpOuZN+NIM+CYpAzTxGHxfh5pw+pXrXcS0
Cq7+uKHDXzNOcw9mChypQfa9msJrRH2t4Eb1kzUjlctQW99um4KLZE4IhLZHqTLusa5KzHnj0IXK
jbNz1iGURniftUvUDFHhcDB4AoxX5P7IaTwFKRppVA2Nc+okLmAb6nTDrXqvIYgraf3dRyzdGXBK
XdxS0/aKxKWZixWGfI506t/kE5mhuo5vXneh+lcfFYwjJ/vL63qN/2KAq8GjQiNXEORX9INzqOyb
gc8Rg0UDjC6YfEFfC/3wqzZvyyKU1S4PJaI5LUZmmS+6BBuYotgAr55wAq0z8p1Vd2BNpK9lzRh2
OdkmleNsaueuUXMp9x6p/TknvqeI4x2gMD/0SZLbF7KMMDYId+fjkORALP3dhvOaVIBFMPGowma4
UVMXqJC4v/oDMNl3xJFNc2ynA2ZzsFTPoRrNhEyF66xKP1w5yrbj4KO1rtDIjpYfhGEvZcQQzvvG
zVVu0TzYZI2oAxCKef0vV0uoanliXA7PM6DMftAKrGLdLtrST5zeOPSB2PB/Tyryn9nV+YaYiFJz
roxcDx3nxCYcAzDRShLSZg7NK3jRPKcMnOPkDsn5GhrqpJSM4CRWF304hWFKYqaWN1fvPgifZWUf
PEMNabQ4Lz5q3qU26StGYjd07qbqHgmwa57B7oKBH0lD2Yy7QB0xbVyIHD+yO41WWjiVEFgJ31vd
kzl3Nq3xZvb+o9nu2huK/B9w/Rs2wn2nvC0E2ZzwhGjjnDhP7PYRTIwhTWzFo38898c7HkKLTk8f
foEVxICVGcqftGgciz5i5vP+G1FkyQDCrTGPin0cq3+sqHYk8j46CysKezyCMSFlzGd1YmQKGI8k
7bCkK1diTH4ytrE4cFvOuAhxqApWd3lxLF5B7IV3i9PUMk0ZH8SGBN3dUOjE5AhBmSD/IGMM89Mk
KDsXN1IjtEbhuWaWtod2TISnnFfGYbQxVxAiMY/LaMyQrQwWYaas1Cs7Rpmb2N6vT7PKHV3i8z6h
DIiLfUqK1viLXldCmtUKA4qlsRDjgZa6UtNvFOS7xLEBT211X3EyqdXqVbNSfX9eyoKnL4vOBu/S
DyxnLYBBFu7ucDHsw74IfszzA9DW6OkCyd1MrC34C+Wv79QHE1jawQaOnQlOHdMYn/tPiWpiO6en
/XXUaeemOBiS5Xng3TAqTagZLkw5fN3azCxg0GD6lOCExMwpQl0uUkWOdlr90jN67GAN/SA2WGo3
NWCBhhFcSUE5eon/C/fNAApDSt6OLaGOzgCLR5CDTJPNsHk4sYYuv2ylPJ0IeK4gyeUYQj9P7f0G
GorlPSbGBpf8kUb85bWX5wLdgMzsGHR2IhpuP45IF9GNkgLuFkL2+k7Bl7bRjmj8AUoXCSulYilr
ohnqrtJZfjKE2K6HO45pZTYdw/9vBib9/0qBS77h7/KlprHRbI4JnxmMbkzdlbracIfCqVYGR5YC
MB9pKQx/NgpslmrZUWpQnxG7L2hzb+nxltPCYG9dKGhv1/o5y1x/sfCO2uezdWbpdHmLyE9+Prw7
plMUAfLAr1S4I/hT7FBmXDamN50GrOtq0fc1LtqGzoiJMOweKziOTyIBNH+e9qZSehRIAyfJpLoN
a/VJ7lXnVek4hF/Zz/igro821rFpWJPtEy/gh/AGW4qv17dgD9Hx5ac1hDiSkEA4KpPxUNFW9K7T
1eQpyTyAlzoYQkm967tnI9lRZ5pqW5pDJ0Ut7077FxpXWylex9DosZ0jUGjAhjY+hy681if1jntQ
ffexIQ8DvDF6rdCqzY3K2549EjxFDsyHDx8EcKGTa2VIHs3ICVlJyAgQrnWX2mYrg0WYbtj/+gik
cB+lLixLiB6yJ6xgXGnMvBlSt5kj1MeefjBxH/RYupE46UR1VAE8jPs+hwrZ/JO3Fgr4F9AggcyO
u5v9Wf52MEguNK096u8xXzlhp4fsUQ2SVSlT1ImpNmt9cdbR6Wlo6EjDE35hlCaVW1FT3cGEUxEe
1Lufv6TvBIeNlzUNUToBEGw3VmsqV49cZtEo4ztGEl8Pk8hP4ebQdPAgBsKPVYZ0Ws7Em+Y9z/DR
VjTL5qKuovjuqR+0w5B+nAjqssYrlCsmzwNuom/x6hGzWjEi2F3M8IxcNi87NJorOYGPt5w4cbaL
CB836ycVhum7LzRoGsmg4vBYC1Ea9iEScfiRFz/2AKX9fCYvHdY63hslJAU0ujKp1OrhMJfuWrfl
HNMDtgE/+Sexe1EKdcykOvumMizQP57bc8XmSfTCuZvwL83BoARZbSCKhsNgQHSdBo7H7ZIJytz7
D3OyfJ3LyzSOj2t/XX0hd7Shdfmuotx+JRB8t7He9KQtvXdRq9xHjQDJWlwstbJbzzrC+vE4siIY
tGZ46Rrt+gfa/vzghocQL0U4iFIQCFwW6pen/YTb7Dr5dSRDaNOs7+iQyaaJOXnj+0MH4m0KZceC
x6T28rQkjn2nKV+D7litA2SiKJxNuBzwya/OwANjeF0qT8UWPeVp39kBJaS3lQdqjmuIDTf4JxgY
FrBZYD1BS2UwvlYy7KsKuj5M75Nl4vYbyGcuMFRD42TCTT6SlD7yJKK2WNusxFjYc2NhygxwpHox
cn0ySwDpUbQTGVniu4dMSRvAE5y2+mUNj2BGea/AokiFq/NGj9Zz91uM8RFPRhKLoj0YMAcK879V
wZm46514FhX8tcofLOkdcWkjWX0tmHAZQEizBuIfQjMo5sjek84jBST8BfrjEPowJPdBk0GSnXoq
YqfkEZbxtfKMe6seaxnk8dqtHmhqSO/2H37KpjX1GTMwDXyl3TxE+l/pra8A6vTbdrhKGiTyk8iz
1IPshEsUUqKPVR9bQu90rpGMsdEGEhYZilu8tkMi7unqq81afo5AG06H9WumwUqxk66jNwSI64EV
IWouSlDrWLMHA3oMo1KGagvdwF8BJ5y+nCFYMod0bTMg7512zlSjQJKASO4WoJBSWqiRWpECSp3l
8DDugycisrdtzQLsLuPvzQu2xfM93nsD+HgRH/TUFEWTq7sUPJMDtNGacHgX5XBuoVyevuH4JM3x
ERnRQ8O5/mF4ad6JhURclDdH8Ta27jHSI009qLsoXIVqFtY/BS9wFRCW/dyijCMs+KL8hrtnXfik
AFsTsNkS6445RFxGOc14JVj8xUhmi4D8ipXVINgiltOAYzBxlYIZ8DTEV0n5RljyTHIDg/q+Va94
6gMYumgM/ri2uAh+dUf+gODjAFKdfaLqNZAAzUw7hquvMbKFn353YSvUSd7O66BryxkbRsZ8gbdz
PMssjO2O8CekkJKErre0Hn6Kf+INKYD9YTCNAw/yhPfb+Ks250iJL8rzE0RIAsrkPnDNezGnVG+i
1faFwl3FXfJdITaDKlpBhehFDODsqr3hNqIxHHANLKFI7D6eYtgi0/YCvAuV0qRFKNQDIHWF425/
Na4g5HAei59Yninx5AdYv8ytHq17gBiPfJGPmus3SH97qlInr4WkG6vHSlqMi6qCi0vmWaAAZR1C
WauUqrOzC5DbspTEMkrTSa/vHym1NXzytJG/vxZiw8wHluDkr0iOKwQ2cxBB2gv1lUZMAvwYn9b+
njET7nd1gsAU9YCOHB1yBoOiF0iTxfk4zKO7Ev9kfsy7Z2lUTMYF9NOq34eAPLzOH1orQOGj+vrl
I+G5zONGQ6RFAneb7z4l1EpfbZrt/NlQErNfVYAu5bQywyVh58ZY2Qxa1ocS2pGNBoQPYHD26CF3
UpanREBOk674gUPlBPj/x79+oVRCAffx3Sjg2hMUPBUAoczLq+tuG8BsHEmKRuIFS4YpXCAfgWNO
cuofets7g+rD5I9xqcoFWnrpWXB6IYAAfTIbX3z+sKV1LKpFETnw8Bt8vAQryX+wSROhkaG+57HS
UtDlhJzjH7x1vNYYamMN0QmDsYwDKV9yVHW9hoOu98Ht3dtutLggeFnCjIpgQ/YriKryj3CSP9tz
68xTR8bXE3P0J0Oe4MAI4TS1oE5Il6WP/WJL10ive/b80O3xKj/E16dg/GDtgfjMmcT73dyggi6R
7ljM/Ai3rzTwwnI3/rDth+VmDDgQ+H2oYFjiINtxu0Qurko8k8n/cTuIGYmII1RbNl/wBsEDsnYL
4XdF8aFIf3Wm2556bzWYkp1e7+Qgal8Yow77F5aYwkwzudYTbEksGKrLhyqX5vpHIbsHja0WZplL
IYe8cQU46R0DDS7SOMQdBUwigdFXpoSX34wA5Zv4tx6VJQjI3tEvXFXMZo99/5ELSYNyvy2IumcD
ncPUvBsD+nPjPSWvVMMX2swXAmh71vSQS2CpfEn91up1WATTebw6/vbF5Fc8Sr04Xo4HMHZZ/PXZ
xTZKlbX6Z0E58hEdi5bb24gWR9VrF8l4qjdcx4JBvfkC5kpjWuELw6httAXWHQq+s3BE+A4RTSre
taRKSjbROHA5Ztah0zMJxOIBOQpujVPunHPLZpI515IFxTkH84+ADBIuvV9f+hIDfvLyKkzXx/5X
RmViBjFo+lqJKhKojPZ8YsIrOuxHHpJQZGselhbRqhILJnysjdgaRTUAl43IiK1lKpCvLVJrqCUk
apiYNllQP5oTG0rBiAfbN4h+A2VMRb+YdtkyhwtalKL2tW1Qonq40Gitb65wjs2IEtfCXZSy8FWQ
QIpI+bk0VCSCVObC3YJhQlwWA3UpNoZmeTY2/cxkxj7VIKx+bV526ydbtZfzy6vajJMhiBjKMtH4
1Fe8qqYrPRyzKEFQ3DPjiMWyTO+Q4tCkIJh7YpMZau+sV9Z72++mABNw8WjLL7wfhm6GfQaP+2YN
kTW0MtTNt7dUUwDn1L5iP6NxL5uBC/+14eVq9m3Gd/q7XGd8d6TFi5NMyugAzvtkShyfYEgWKGzX
GFKe0R2spBqh7HtxODpVPwRUpNXB2hEcqN9irnF4PmXuz60HJLXUYHoIm2s0BT4OXrHI+/x596OI
eslBDT94OI1KpgY3jCCiwz096Ppz8PAxgYRVRLkkfzrIHkPNukb7LrOop6Cz1mJTwjv8Adn0fgfW
BJIEp8TBf9eiR/N6whWalh67oYFhI+7Dt7TTP4uCzDtBxmV9ghMpq5dE22TnbQEOxnZta+7Ez1Mq
Zeh2we97+jIkTpdCCavmDFIdu7dRVr6cHLpYINw9j0LDcsXOBf+w4V49CodYUiQxDJVFfNcZUkzD
dNJyaoIXhvmzBNJWEd6PaTNRn4seel8Pm7n3PiPvPjCmyk1gVZ/dyEzKrOFLxBmoHt5DNarOBePH
uhmDD5vk9FWFQcg8KChvVnRDltnKmvMWCs6flTIhjskG3zqnDf2e+CwicVms+cpEYInZkpAA4PDK
CkxlM4n5K88ATIudoh2TW3Co1qmbm2fKvOEIo8zqiHWheP2n/1S8Md5iqzPWCGV3pL+nfDdJPWF7
77Vc+V2URIyg83SHAJHH+flB48uL3loX82XffDpFY1OHc7cMcoPlbo1XC4b4By3HoeOKuUszI0xi
92R7jOPSkpTOito2yseUUQ0wQozaHzMnqBTNs7+ZUFidVEBmbWwcOpY3p9XC5pMl1RLpJ+M6LhJL
pP38PhYnNDsxYKpFE7g3oS3mGMLdldEiHN/beYDR9NeiBLRyVkPMLQAS1kDH/6RB8cGKdUIE2cTU
sg/6fl5r6JI0Je6MybLcckdIJLMIKJg+ZyQrWmrRZRh3NryPRCIk6moImm05Kt6f1rvRpgnwXxKm
miFVEkeRIEwKf5uQiaFQN5yMWdK9NePBdJQx+8XqApuKzu0hi5g2SaXuc9JJsGZiuId+3wVVu0ij
NYZsKxdKkTuubTlOKtul/y4CWB1lR7jt1DlBT0EIJrvi302+aYEnaUs6v2Iu6hnPP5OquENTFfIZ
xoEYUBBLIOs9YP1UjcOU2v5aHlDYJHqB/vHLTk8JbFmNe5ZW347D67zaErkG1lR8WidF8V8ywXso
l4TGc1AX9XKgxF589SpKYYyefo76ybHxg4dbVKo9G6AH7ADxtZ6AhcyPadksNblAywsQ7/+S9S8U
ktkKSHVJX86uLLrtU7aJ/01o2IS9ui0QB+twknzS93YYqdymJF2Ya/wBhgw9tv69L9H7lXG9/lkh
leG+Uh3Ib4oSjWo6C+AAxBjJlCPoPJtmTmWWlQIwe6D+E8785ezYbegaxDZdltv1/FQznfGDmz0M
zElobdRDpdLSfzqLBp6EVnL13VcfSKwlsRjlAR+P5XD910qYxjM5+mfkAJ4icoAhxhzQvNOJaNk9
GlcWCVv2nF4K/xfmcNKkH4pq1PUxUXXBbTpBuQx2DB8rXXuwwkLKDAqKz5k9aHHnHHTgIVo7H5IL
IJi6ZMVcA9898IDYxw0wfu8jwbwTCUWkngAu/8s7Oq+8cryM1eb14nwy85Q8iWjcoUnF0L4pBnxs
ZIdhGlemMFIpPMiNADBjqT3f6GiFk4x+OjROzAqFry8e1QbCWELlz9tFAvlfEf+us+PVsmRjScKG
xBj0dJVA6JfioAnlqKaTDozIUCrTFejW4ng8i35NyRHGw+FK1jIS5+JZKF/GMBWQAm5wMuJVbgu3
MaQWnbM5U/RXTD1+pWNKObHX5fmlVKZx5Q/02VsNFOrrodnWFY14U6LDMGGtSm3MsxVsbsp+zGW3
F4IZN8iYfvITNJZZ8lzVxa5HQl+PI2/MvB8Yu2ipoaU0aMMteQI6zJOBrxfePRLRTDZXoenk9cI5
N1AObsIk3LHqbytkTpR0okly27YZMUpBhX/r54EW7POh4ymwz9jolPdtXuQ4Ers1DXESj6HKuOYm
OjEntr5laKIGkwR7uzRjG+GWTa+9QFW0ssxLE1ftguyGtEqLUZgoQ4YOhGHcrJ2o2E51kuyylKzw
0T6jPlwywWMCkbQAS0kAbnhPt1MrfywZd7TbnWgOZf8xKyQiNER2Pa7Q76EfH3XvEzB84KUHxRuM
KSk3yLLNsJMiPa3Xs++9DJX5MDX1E7JK//k5vc9YrzLa/GNhl6HM6QsqRPEqSKlKrcNidYhbq0XR
UGqqndX9IX+8HhQbdWcBlJ5WKID6zSpEWcySf2MCSMZT4EUEsGGKuvpOlFHcnWpCcGpDMGQVuMQ8
oJpGTwbVYArDqVi2xdltPwXVy+oGvFSusMaSKwSXITDFWCiIZW2yIPMYCexlQL2GVfHf1eXHvtbp
f2R4KjU7wFZBqK6iZiq68CMuVkfXaqAgtbR0bvQatX+gl9//5h5ls+sUBEPpGTMOAK7FXhS/sBw6
kBQG4HwFyIFVe06vs0ZLOHG87SNdljA80mQG5mC0PvBJ9daeveXR+3zOY+iz0T2K9GDGdTpxqE7V
e4ao/lkCz4Sjln8shJTe4ADpAUt8ID8JeDsnDznt26YEuhFS9cY7f5eqFbntgRtc0qEhd4EmJVUU
ctts6fMF8qg64xOs7HBonfO90w7lOog68USlRtF5vLNezQmMgifz8UDyj09y0soaumg3vPm+7YGV
hUS9Y5UGyBRCQyQTfeMsLaQN566XiKzWv3UD2Yd1vZ4N9d7vG5bq9+9Ts+ZZP+j0T1u3gphZrhz4
AHyasmpGGqdgOLUBVrivltOU06aBFluzn53CJcnUw0C4KT3dqo+p5Akf8WdkhD/QyMGa/hwfV5eu
lgz2z6xBYtH7Sk/NG0JGP7o0UhFlDybIb20NNA6NlHvWJo1KAdF5i+TwPcpdBkcn9zsvWINOhR6d
5En+yVucYv88H4KVsPH2A4Y0GdhXJIDQcP4NMGehbcoVTLnBwkq0nNT1rhIuDAxd6jCZ5F+8jzUm
EPFvgKkCYaIBSC+nGwqkYodXF5yLu4GApqFI02FYOIDpKc/YfkALI1PIju/+969CDFhCDIcdpJ4/
M4ADAB0z+kZF3OmVi2J9MfbThZAlBfrSqZKhlknxIDPq2Ez3h/p/xHPYb1TpVJYFPSC89Hfw0Tsc
942nrFZjutcAd9DyAcWg3ve3md6iXEE7Qit4jGb8LSQ2yIkS0Z+LZw0bVtj4G8Pc6EG+HqmLaawV
jlI6Py7EoGRwNlrrY35mwjjJFNiAdn2X/nbM9XMyvnvwp1qad6xoVK7Dz0x+xag8L/8Dpi6ModvC
vmF0rZyz0Kxphgrv9JjETkT2tQqLU71T0wt9UQb8iEg7v+b2i3pnE6Gn1oG2AE4+3FDTPEMs0EDl
HkGSndXYO2iLgUXjIQioUJxw/HhU5GoQTMi7NXmUAZydpyPHrgmFNQAgRW45Z63ZEm1/z0TlO8tX
czXY0UOuvFBpgshIbQko1kkZpphp9UzneL8ClXt7aK6RhodX6xILxB+S6oz/ZET2RAevuwnkUFrx
ZAw3nNZ8qpfBs2LqWJIx495wXSdoCi6w+z37Ll9pH/AGw7xNhW6n1Azsg3f80XP/1M8w79XK7JG3
LP7VAERxFCh0w6p28PXgNwCkP8C2+qy4X1EQHDVet9VmniDEhUHCBflUc58ESp+/R1uBUpJ73a8x
IeZjmVb7z90JCXjWA+001aLE4GE09HUXGRy0M+cJxSY30RliwqXZq/JD9EJYJjAmq8F1rJtNKDpC
B9xKUKQx4qxa5+Nm5comCeNBh2KYpTjf3AAvvjoTdp3RXUh1pM6Ft1P6sHj40FjzYws3GHArZE1r
UTXLUEYbpMSAr7UcHct3URqR40n70fDsXHDEfDajmvTAQ/Wy8H3+DN4h/2xU2a6ZszHcN0wnXwcJ
BPOXh+B8lwpZyI7CijmowdR6pA+/6nN1fNQyo0F/5hbhJiQ35FCy8oNwUfJZV8T7QBMf3Iym9/9Q
yleAG1plc3Wg/6UhcRyMqb1Zjdz5OObssk17vOPCKpzzNJ6ltzrnrm5zC+7i48nRFrb4dd1cwfje
8dLjv0YifcLqJ2omDARFuHigr1FRsNo5TKr7qt3rDzCiVD2KrsiEuMwtSLUmJtHO5YBO4uJ98cYo
boBvyAAxfkgXbOOBU243cOiKaeluv1MnZXvAT/269F5PhVLcV4QVuzFTwkPomXFNyX/OKEiSSnKq
WvzBT2k4reou1GTr6LN1vnk4MQY6J5U9l/OweNwMmT+7ByM7CjpC9A/hptq0KezTFQ6AQFZzk3xE
3uj60M7feLJf9JWY2SwUNiuquCxLmyPIJ38Pm/rKXq5v0PMx0IbjXwtlTiIVvtx3xuTfeqyyb4YC
i+uSHcy7JbIxg78QsZv4PY3bfJJ0TfySVdFu3Nknkz03vway5wZngz044YA56xIFFeEkQTllkHyN
mv2fwP7OYIKA0f9FrL1O3CjlLgbWQBtfHFln2OoryyKa/wGBNMGcktYHbnr3n6P1ChDFWjuiP1c2
BZpnlObs1JdozxhMLcbogiFD1vhkFH6o/cx4y1R3X0AZZ5Tuu6rsKKdL8g5JCgVRnwSxT2NY+wGX
2MFJgDY6TcCCZ/RFHtH+VXccr5alDDKnWKSAvNkEXLJ+eZ/MmlHYfrTFo2lGI9cUaE8SqGmGjCGx
zsWF5QXKt47tRctFZYPoo9erRCyYRBzIKqJHB6HQfUPwPqsXh4QyjS3Sa/mrrCTxVf6cd5yxA2U5
Gzlhm5IvQs8DIZCH4g0MHNXm7pxGUJ/ZTnsyMKP0wjYBwRWZ8vGY8TDqJcTegRNRxANPGBLE+jCU
2VjDIDEFhHbVgs5AiTSxmbHF3Rpmsom93vgDTNDKs8n9LJcCDPrCEP7BIwZuvvEpPb9HtRjdHoFs
FDEmZ44v5sqRc0EM6eufTEpZbS4uiR5SzbFU0dz4VL25fQGfyiovWEYxQraU37EiT7rbDGLRM8Rg
PbI5dO7cS03VObDx4seuAm7BhJM8DNFBbRI0bweARg7QK0k7gLU5s/LUqbThN/TsrdhD8w8GA3ua
8wTJCQ/tMXBLvxAsWvVC3wvPLLqxIzxS8aUTS4HVAjaSUjITy0D39vL/ie+130t4UVUj4VXT7w10
E+TntOJ5yQ6r1opR7LMEHoLgkvHOKmSmBFMaqsdorlh6PRpzalVaZafSKC+EkHEwpohVUHoJbLrd
TQoBYiPbtMA3GEgPggLvgVg4seiz+mcHci41ksx5dXzxOHYK2/Cl8wroB0BrSeXKoOf70+nBL/of
Ljc3VnfHlXLMcMoM7eA+A9nPVXaI1D3gr8TA3gKHuBlMQ5IxpJjIGyqOwRyGH4rhk4WVbRh+jehC
LM09aWTtc/O2m90al5jAiz8mcmFMEofVcJl1fZkwnwcx5WjD7iw5hOU70zb1E0mREonAdUD546p5
dP71pDZq13AvIt5QpUZ/tVXHc8L7W+rLBBqTpg0chlMdBO0ViCC1TKggNfH8oANRKiZUL1GB5RMw
j/7PqcO7GqRghA6UylZZgIjFl2sLwv9cVijCKN9Dl4XJnjTwZ5XLdJKHYEGTd/XKiAfvQWg76/+u
9qlN4fSUHdNXaxsE7WAwoiRZg8zrd4IHEl6Seg8sfiM6yaJr5dA2FEN9hpftZ1FTEFryOWVOp4ZK
vw+6rGKv7GhZaCRZs7kME9UnbZ8UswLcKQukusHjFsbWsVhixAW0zcZ4JjS7L9ZDFu/rRS81cHDF
l51YCThp8vKIkfVH9ryHLWbAisPfMmcNOR4Jpc/T2c835OrZ0KoQSPSDd6xU3042VfjGCDTq+lwC
uwAqNG1LxoGF6iVwsCNMfnmL9sYHweJD4BgC24UJit2sh5n+PmvWd+XwabpaoPz1XiTnr+L+jKj/
2KutG9/eW/XgA6IX301+AKXo4amkNvMdzLQEApJRLlraucqQrLqrvUOM9hr7ZOCu+ZXMcGzuTf7E
n+mG6zGECZMxAqaXGeaOl1tGppk8ZwSTDet2gj6pUGF2E6zAxF3d0s6P/Ou2JQaio3GZQFHg72lq
Hh2mmGfQv3/L6ligvsLLlWdfghWBsc/76/k4MqToUP89g9ljHU/gJMYt4Q/OJ4hkbTju8yS+l1a8
uvvihE3McxtNB4gllJGk3vs4fsrW3B87eLxHLfi6Her2YV7do+imMeiuhxNePjPxZCtyNTzs/4VN
7L7f6ff44qjxxKEUjaL9uGoWAjgZ1mmIHnoKl6AuEnN2fIvfqgZ59OW855/5c2Ad0ST7/BZd0i+N
LbgoPs/8pAA3+Xu948xyKxT98P3PD+g/tTIuGiZ6utTwmrJ5KyjhRWGZMYaMgtfjB9OH3Q9TgCNg
0wwVeEQ4adw/PxZ4JEMTDGIdoXEeYNAt6NZgnpfsMUh55RkI835At1uUQX2VoXIglBadHDEGcMBH
kE8ZqLY7kOazLnqqbKBdreVwuktfsu7fazvzr8SDEARpAbGMTZoPdP1vtxS+EjLGynxHOaTNakUC
GHjpbTmTdd1GSyDzdct4UWfdUOJAJHxOsUQnOu2vHEwldOaJ8vwpB/s3gZS68/HODDmwpec9I6kA
yso2X44ulN1/EVcNFnLaFzS+BGNAOKHab9TPqSW7G+hv+m5fV4DfrWbF/eV3GIYq2kkETgHegQpN
oSkkS6VQ9WftkN19L4c8tU4NkK3fiJaDZb58KefWD7NTEtdqqUPstbsmWnoMtiizdkN488KQMGuy
n05koMKkv0PblHtec/Bg8AggPb94LxD4OF6Jd3nrx/bB1oXBIJdVMwLyHJ6YVXDbIAix9MBw+Q4N
vfgs+QNtHHlCuQt5XFKmDnOZD5B6AY9a+o5AjiyDJRuffkJeVEQYtwLGLcGsibLex2CYqoyXmW/u
622LzWTG6UqNN9uu/3BP2ZoWm7jPuT7JqL9p0394eT6TN00/sKsCha22Jm7SKebjF27HtH1KEaYU
JWFQFwbtqqLeAwU+yhLNsp2XHPbBUO3VKxZNHj4Jpcv/D+l5BO8TjExLWxaaBmR4sRfs7mq4bAHt
E3K35iHc1ibuWQL3KOuFX7soRUFPD7J+KVkr2NfkgdV9AffncNJ1WQar09LbPRJdZYZFDnxVcV7f
GmNDWtJE9q3sVkbJLOxM//cSmYVI9ZEzr2x2S7thx6Mb3/oRFZmF/rEaU/Pod/xDWEYYqKibhXrQ
zYa9PvYj1lE4KvBvZTfDYQArZuzNN2kCmHp1pQ7aP7eG3Yl/O8RR5Q1dcuRYfU9yGG/yjYDs0MTT
6YQFmuZmrCUtRxV3mnB3DgoQwnnjM8MttRYCV1jfngnSBGgCtyHl9HzUFBl4FS7tg7jvcdQ2uyZ+
HndRWLYdBzM2PHN71rTIaUQqr5TbIZhbzAtGd6Q83ZpkAuwysdPTkIhd0ibD7H2hVKgE+Mmaphbo
QFw6E8VsPkfnQiDnIPXzT8LN8CvzgCgUUucSeUzTOdvLWCypJyJuWmf4pImvJJmsiYRPMHXxNubX
Q7/wY8JMdiBt9V3STmyT05gjdAo90Jgz9Nh0d5BlVSZ07ej9UweunzopCTtaFpZqHmKQ0SZz3Ofg
1b08EVvLgFZe6xuSK7mx12d4wZt0ZWa7XFZm4VALsnfBz0C8bQkwfIYMr2bazngXcmTxVEocM+sQ
vY5CzEFwlGZNvmkcB/5x9A+V5kDeIDE32nie6EQbSdHjl2z4pMABnXDfdOd/0ANPeNfRJDQRp5tx
cysHWZR72k1PqFKcY3DkR5bIiut5nAvgmPuTrY5WNdUpG7YQ6UnolEPE0omVeFKg7VYYs+AFqpt/
zVHxTQyu5+dJTd96Hn9Mc8IXgL8UPQCpVUFboENih2mrNiIBqdzsDWoMxyh5tIRqmbVA0/vDu9GH
jtrGS0Tm3szhfgVZdb0MTqQeo66WqsSg483gpEqqThChQFSKW7gm/icpvquFnFYeiuTmIEgm1ISZ
fUM5umfEI+PiYBFfUPfA+UPFe8Z5XZ6EBpJn7kWLRPCHzTV1EWpHiqkKN7ZlmFBv5rNuV7c22/Df
btaYi2qiZUc/5Q7vt8PQoUD5vdyxAlfVvVv/gO3ePmnjnjUjI0VZPGsPCnXeRZ4Fkm5L7aMI0SbJ
0rh4tUWEy2VB5Y5m8rm/TrcleAyyLuKERGdSBxr63GRZO3lZ4rASRNkuLqrpSHMp0nEI8tZ3QKx0
kyhbK7/MGCkSEcQ0yOvI5iueJtnSsLo5QHm+GQ0vsN8aXaoAcnEFG8LiZrQUIThxRmBMx6Ju/kl5
5yJsZa6NuY6lTU8acw0cDMaI762F4LB6/R2tfUZsk6bjaKVQwm3iMA7/mDQlY2zLJL2WDnPinWdq
I3FN8IQfnmmo7sdxwHSFKdvfAd4UvWVN/CKcNlbyOpFx0oISd4Zy3QXIBTH43rTs6o2RVbdomGj7
LUHjJ92THG8p3LLNETql4BZ/BySIhz2P/9PF6WpBRSRAu1gCWXMjkQy4zcMDc8U+sGzbEmwrups9
/2Q3YB+kxFlY7hhFRXHcs3xKwPr1D8h0xRUi8mwdwlzwIMdwsmkrl837Dh16Pd7gqIDdf2p32k++
Aftf0xNstY1deK773z1LGPh2zpp/gjDPZ/1nwKj1YjneciMVGuDEGojvuuCuxh8gaDkPJEy3pJ+F
SbdPklw+DyDwdixpRmqsha+BCVuEIoDMtLRw+euc0rgJB/qI5Gzc+8X8V6tL3+7bMf2zqLoAQceE
9hPduxYwODfBqRQK73McKPzD+dM44p15yE8HeKE6k2Rw/F/KGjd/ESTEHQZJxflB+jOatk/Dqg7j
M7A0dXL7+wiVSk2yDqNfo8sbVDMMW4LhQPzAhx4gAG5nO/t/qRAN+aA/Ky7ZW+nyP+T2eXhdK6IR
6fgLPt+beDBFBPeKFYrDxcuMDd+Rh2a+UVnHCCmotobnD0T/VcmOtbnRBWrIO3KiCNJCC55Jfqtg
cJdmaZBlxQO1VdrSmA/Dckrjeycx21AmuqhJsfeEM5nMlVqLGba5JlD4dlS0lwaBi6wJ3C2HTXsZ
iPeOJnroPmChImBFpmlsRv9oWGavCpoZsRJF8vh8l56ApLcBUO7p2wskSHJad7l/NJNOXlhsaprl
Pn46JchsMnJNVdINRnNTgqXhEaeooS1yhGpXtOK7UGIZcaGBLQWrkq3Nc4R3Ke+9tGqgU1Mu7Ke8
3M2Q5Ne1yBYvc+X4aS0snjU/xF+nD8FEcsvgtzRQPhULoGwjD28cGUY22pYRDtl5IxtiVJ9SGOXX
GCC66YL8DQjs/aZxs5eqoboP4WDGi84gCM0zsqGnSPFwGVVpFxOFwL9njMeBbxRxWZR55sUszRBH
qUEQouG/9X0ef7tqCNFfmTNyuCcUlWCUHrAxJifXS2BuCi85Wy5nFOF7Wmg8vCNYp5r6ioiWrUdd
pyqOQ7IPcfB0K1ikFYWBZQvtiD+P1YglO+rxKKuN3EQM23JFT/E9mEDKdVd186dkbOq+tOam4V1X
dY0OGFZbwXd6jgCjk4NULzp8ntEpdn4onl8DykezeZWM2RSJZZfN4Jmsr2kYoT7tSODcG5yNnGFj
QGNBYD2BVNa3PdbqCRsDxyspKkqBL0lGgHCa3gR4D5NTPmcfXq/Xr00QVdNmOox3twuXTRuDtCiE
icRXg1kz98YEutJNmGQOCUWcnS8wDTjPWdD/Mg6VmPKKbwfh5oycULSCpcuuOllgs8OOQc9b0Myo
Ym67jTIPX9Kbruww2s4Bfm/i9P8VAcsmtUIaveAA1clBIYLFoM0E6EqUSSFp7k04dtpUMU++LBJr
xNTaDfyglXtY4qyYpRj9VMegAEngW/DO9+t7s/cM7e240ZzkD+NVRn37nxWgYIyjC3dRfzFNf0ym
n5Wq/75vyEL9ClNrksVlJ/skKbsbswuZJpSm8suUTHoP1SXLkM8S3O8IjoDpTPjJHdV1alsLkZ85
RODVlY09a1LZ3PnEGjmYc2JqzfFurjv5sLfmUpWGPnKD5TqhAJkK3eOCP3IROoYL5hLn7l9Hhus5
qJZTuxycE/k9mNvXWwkIoo2kehXZqHR/VUoFfpekZPk9STMGasxaipjnh29tD1UWvVimIl537HtR
c/5hRqerJPv6n7PMF8biMI35bCBUjGz8KeJ1/nlNtstYj/T+Ri0CWoufqlFZLzT2J7LtNrEGn48C
LZosEtWBctMVDPr3BxrBXjpreyMBUAwDr1Kw1vR5Tz+zDU41IWJgsKnvTVdPhq1viFuIwY1PS4Sh
N2neu00hYYFhVtRsmsLRoL7CG9xXFK7F4Kf8nz9A7OoEbNmyCgeAfdq+eOW1ePBvTAawPT2/iigX
iIaIBrP74cGaK4rzh9HdqSwtU2FQV5989ZBmjdVfLlZbEi+CH/OVwv7+xBlrSZENULWYEoz6mbjm
TE+rqscksKp6JXUS++XmnyQy8fjHXAPSmvOuQ8pnKw2ZIlR3jG0y7rFB3xS10T/qxWhb/A5iDs3H
9OkAW/1GyV2Ajlv4NLZnaidbx6/vglKsw0b5anbON175qcm0DcWe5BVrMmk/h8AVyOpiQ2Qy259e
R8N8tiLITm8icBpEfWNedHlf56Xy8hM1snH2laK5PlqYrdG0de0LHimkxgfTLqjvawfNRCKAnB0U
NDEB5z4/TPrU/N7w0uAF3BvNLrn6/ZdODPxDQiETvTpqN3GGPw/tbJSikik5UjgLKa4elhBPFcgg
9FP5z9Ryxiq6Xnd9/ySrYB/5eef/GXK9jw0Y8nzKSxuxFlLzq8651/LK5HsUNUdf+4ij5E84RUvq
3lyQp36NhHnOvBYUrzKxXEfHf7ZIar4+bNDyILMBL1zgrt4VexZTuTonutlmNjrnZH+aiVPk7Zoc
iqPzeJGJpeVYWOpfK/5C/ql06byeKO8myvJMtCuQSbHC1MpC9dbe/+drtYn4KSCLAeWkU4wOvwyb
lFRVpsnoch5/N5bb+Dp+vl5DzkUOe+43S0zzDU9K/jxUB9TtoYvgB8svPPviuDS5p3YJaxpiWFiU
b4BzUh4WWArSg0ML/nPXRg6Z7MSR5Omto7E9Uw/o1vw5eY1DjSa1Yv6ojXccjKVXyzEMQfqZi2U8
w2xziTROMW502qtnUGszfe8S8SN3OMepb3ejaASr/fy/2dmwu2OG+QN5P8/N15lIha4ll6/PYOwI
78IBTw/fZ+RTWFNB/In8vZtZo1Hmx7UZiSMCnT4v6pS7mbBXPZJ9wQRAHC1Dq7NLrBa/Fh7T1O8i
7W9s535QAsZavcnFJ3frv+hz8b9VUUpeeR6D6ekXJ2ZeIfzyMhsUPk7w3ezu0gdLBbV8SUZxstxA
J0wRPggVu7vwc63Gk7gVocDDAjOsiffBorEbWGUM+LCyQ9MKET+UNHF5k5FpiAtNwEUnD3lFKFOb
4g9LOgpKEzWTkoFDR4eZyFnkMSY1+dqM6A/kUfDYl+oWDAJfQgRDfwdZwRIVhtBjLM+9ElXHH0Mi
asyvI/j79Y+/KmWsQe+yTT0k7XMHCOiRHGJ1EMRv3yQEVvL3L1mb/8/4+/evbSuQjGU2tOjBa05l
zVRrekOSRgQ13iQxF8mEPFv54LHRRlI8Nf+Vtq4yvAxTmJVoRkvfkV82cPVHtLqTkVEkgNtuXq3k
bmslo1spbM5JgIe4w6GhGSCwJ40ETpeb+AZY6OapYlW5QNSO2K5pvaLUXPH1aRzibZRcSDw10JGz
esFJRfdJT1Bv4Z7wBJNIdSP3ZagtQQIH+et/gkZN7JHNptwULaYpzQtD6ESerbQq2thNNTDMFIxK
ausVGq85bEKX+tj893Ag/6An5DO61OgwMl8YTMFHC4jVI3rC/dmbIK4dN6gWQNsypZsY2jXjZsLA
xLM4Wygo07osp82POqgn2puKsrjLvZWl74K1fum/71IfAepVvg3xpDdO+7+yKUSWLwxvZDmmLjwQ
KZX97Lp4WIlpk4FshVnZnq8SB4Mvg6ilDRqnALGiP7t4dqr3DvAaF+dKVXd7ZzfVh+/WyVAjFVrF
wuZ88HVtEzdiCNFVYALaXoIgAbX6XYHxXgeX6O1d+qGm+a3kQ3uvk5puQAhEEeyGRa2vGBB/qH4d
0ShOOvJRxfejaAfDCaMYWs8bQVBwixqJOVG3quQvlx+8KvdAc4w5LLeDrpQm1f3g4HVNiPCnLUwX
y5zHWbxQ4P1G6IEQh1+eJmEwobE3EQ+F221fEVTJwjVNqSktsjZs+2yyc0dFuEzofFfjGBIJHGx8
sr+4ufI0htkbaXYzNxH7mDNUIsdl1esnLVD3LTqrE6N/CpHYkFMCpW0H45C7xgAbERoiPk5mrrEn
Y/6ZQZRYcbLjce9j9Mg5i7yhXPIC4QQKMeVNyAtor1pFXvomuBv/QCKISDTaqoYNJI7FbtELShl3
/bIpuaHHs3TphPYNJTrmEMwn/NJJMwAA4qzso2EuvRGUVClbyBWW7xoxG3Dwatqt+tjPyQ3P3y2s
DbBevT4+ruLkXQRGsEDBcbZHt4nXz7Rn+7lZ3sLlktb5zdf9M4MEjz7jU5bHfeWZM8iTKRbIxzA/
mPpNSr7KS8KEAzwgJUdOFSCtW0Kk0NaQI3quYYF5CkFxXEh3F7L+3+T6dIxnkkoufb5uBdCZi/KQ
3PFMMdromXWBJNgUQh9Q3TPkeunCRXRAqAs1LFK0C6UApiEIMx8Jn1R0Oro86EVkpvKCixq+iKvv
L4LnH2JSYfaRf0j2fXZx6aTIdjEm6+iwr9SFBuEE2hp12qYyxouEgwKicntcKyLhunkdN4LBcsmq
2TkBYzeP+6oV5dYA7X1sREtEyfKqMHEY8IOmmDJzWwwDQ95u9RuiHe35dAuvx+hJFo+vGXX3iHES
mAzhaTMrXebX7rG6BRrRg3IWJEreUfEQEfecdkszTj4fIYWaWWga09aFktDuFAREoygl2rXY2CVL
OZyhjisDCzr88W3kbBk987qO6i1hqhgNdW/YkukFkoHI7dnzoYHzRJR3GuExeG/HmM4an2gV9cDa
ucuEO8oXg73GombjcPwr4hJZv5U78PxKeBuU6NqQCfliUeMrTtpKPrdDFkkHbrTU9mXdSgpUCGLF
UIuh6ejWPs23CxR4LK1xWL+2r4qqjpan/P9HhzIlwlWHEGlU2vgNVYiHrjyqMmW5kpTzzdbLYJst
2sPv9nrXJTAZhvgwsgkC9gXeUTKdoeUV8g7vnENFhMHIz6eq8E8q0B2WKrEgiDEgg1nV6ksAIcXC
/P0fbDpSZhzrMOvPAvvB4C17MEo+GZyiL9104BU9eYQrmLq4Ddvijw7vUfMz+NNHvL/hpZDRv62h
ZZVw1l9FqxH/m8KcK1DPgWzQyFLlex5ugzcpNhLeHsBmjnmzdIz2/UxcPMLATmJhPIoStXSNgnEM
4VHNJqTQoypP3bqtdU6T/3Odz3rOTunjnOmihJsn7056JqVTi1ARS8cM/w2FoQuRMAUkl6FRRUla
9APrOEe897HU+kGuROuQ9p8pd5KNuw5NyQeWWvqTvSxgfIzGRyCCwY6ZcOYEsBaIiSm4pAZDXyjx
x/HRMdm4uzCpWGmjTC8XQJmGwCrYqk+ZzuvaX7oRRI11eHP1F//flHg6BtFVShagmZ8qyF4H4xow
ulJYtxEqj8UqSYMu3nnvctWSjNVr+id8jeRjzRc7q231DilQhEOXd8y5hCCinMMoNbQsoh2p/0s7
JQaoFZ6unViaApryS+bdliw+t0124smRXHCvtBUoV+x+hsTNUG2jIxlHTeNJDC5YctojuHb0XbRz
tp5zBu5pFVm3dzcDffo2mFLdadFg9/sS3V6cjeYtVbRWPwfY9PwwWRgmQqPP60oV6JbN9139LgS3
sMbFMJTwEia5h+Qf2FVG0zqbAoO3aFWchz6NQr8HBOuX3XP0xbh9G0/j17rNucbBaMTxEg5iLsYR
u5e4tbRqSv9Ibt7L4OQJA3rl2hGzkmqH+9Sa0EaQO2MbPiy61sMiDyo49NE5prshsFaEMfIK5cgt
HkwTyxTGjgTni+59hWHgjfdt++xhocXK/nRPCcOzGh9HTX9QFGFcqFQw6FXFiF5fmcmA9X1NFZ6N
VZbU5wLx+6G3PyMaqcHqimD7ia7SkcXQjW3pwS4pipyyDzDZgVXLIwmiGO12shB5b1J5CPk7L8E4
Av+QmC4la3+LOgWwr7Lo3DaCmFJZ3EMTjCfZbq2ouFmO7/O7H8jaTGQgur1DPdxhnM+JgsBMEVv8
6I2pH6TzDeld7cnMYSXv4N3fgHHMKmoGL0Trssmy7tXLL3Myb6HHu3kysz//kGwxaItOv4OVFAAP
hABvgL5kLuzsI9YHrcWZ7uVdmXktfm2/Q/xpYyq7qftP6CBSgCjaGVMO0mik07fC9x0hANbksdQO
ERhcd71mWi5P4/Y0fO2qKxCM1/Z41ZxHQaD54biAFYw4DYT6GOuYwkamycnYYy9WAkZHulPQc49k
FTFNJaEcw7Bb9uuBinoGBsAqx8zlak5xA40tFLGAqPIF/IQmj4lQe2igTBW5E9VlqDoOy2AWWol9
8qPt2SVYxnyo5WS9nqbVUbjLOF+qwL/0DDtp8/ZI13xCrufykGpS1sFPnS/TL67eHIRw/+2RRQg0
gAnlsNLRko7bxcQLLkudmlI6fU+DlbfdYDL5u2pgRm7NOyiVJsAPoOH2DKJXGu7y1UkDm9/OQ/nR
nwbxeFH//5B09CnxQT9Hm7+jikkmCz10bafzor6jEHTxSmS43WzN9jUlipmj8mo+9Wr7D4Dfn9LC
QECQkUgZFZIY8Hs3uTmVvkpNgQbYcW4IiOoZq6T3JziZZB0Ypz0rRaXE6XSXWtkIPKZWF1rjK8tD
VEOrcqkQVWDLPBAzWVoagNoDTZjSdxkwLAxA3zubwfuneeWoZZtIPmZOEvx/Cj3pZjniWl66mTW5
EJBUIfMZkipq84c0SWPvkxJjbns9OMLzsGhC6r/7X1FCtf3CT+aDko/fhOB6infV7fNgAE3ME5NP
eQLxsNPBQg0EWIWLXT6GHg20yHoOGCYLqB98H5/GLRQBs6bc8WIpk0VU62nmk6sA5sS3mWLAuO+f
AJ2P+RwbOs5L14YAzIaRIAGF+zAQk1XkgltErTE0AANSDf9GrF9fZXssUQSs6kxI9ni/ZeWUqqR+
JBwcX3IRdS6qYf+zt5a9PqZmM+t649xlMZtbZ76ITVriHBn/fv7lhtCrdb+d7EEBlY/8kK6XUjds
DxsmjiM+vOIP2Twf/7DcBbIY/jpdIxyzdkzIS/jouBxZ9RB/Q57LfEl1B3lSXhz8P/oo5zyJw3ia
O7nB7IBYU0BmHYtHq9kMV/aVrExgEEAAm11YJXv03JNlVGK8k68efnqQ56mT+Z4FPgqHQyDL/d/B
n+eEfx+Zz9sUCup4jIniCzZ2FJwcYB4i/7ndQ4e1AfTA0TYuqwSk0L/egJ1Wk82vlgj67O0RcktT
BZTpzsZlgtsy7CB3ubyJu1NpdPi/MZ4OeOwmk2aUQeyoKis/WjuUCbIjzY90ZAhSsXx7o+1X1edS
hDdVkP5Tge8RL7M8BCoHeoRdw0f9TTbxE+C4ERxUxNmoxONnc/yPYBisLUJeG4zEuX6KjmaVhCOl
e9J2/nmtjQRaCwBxpkYb0/KfPaW7OuM1591pQDwnDEc9WO2tHrM9ernKahd0ZCHBx4ATIKaoim2c
P0a53Ixh1A5D4EY6gVjJi7mkR8ByzvcO6AjksuXUsL94+ZIE3oPZughumGfm4yaXtkTRSyotKhqF
gtVL0xft/opwI4JVTVgKb+v3mj/VTNSGwj8xjX4vEWPYW3pSeHz+y+mbP6OqNJsnyb+t2jY8prNv
E9AAQzQs3PGvenjLbZBzxc9/GdwxUQx10qESClodoHmrwfrMAMv7a5OXxkH6bghhKny6vCoSq0Gg
GscD7qXJnQVbyYH+moh/S4iKRaaPWbOpjFVsWVNPl1lxXKNOi+qviEOi5mtG01CmTf2vtP+z1GzM
w+3p11JCf/mMhtjKmL+PulIzuFxIBpJsfWANLOedP+7WxmYtimQbtkrZvTmiIo6G8k7W7nqchbql
Y38hoLaPFZpxv/V1NASKwVSdxqYnj8rFIXMjSFGZzvLamLJts6MV9h6FYiZjcmQICOrOKBJUpjCn
BAssxV5F5Zqw9ojKQaEFWnM2PRwYKIQFMQ/cVyjekU74CUzvIGt6Dh3bcG//PjJYMEJFbYLGJj6g
pYl45HuiZb/D45ev3oelLqOO3B2+gQoreyqI/gIpXhpzst3Ro/hl4Oni3fZtYy/HQ6VTA9T53dgC
ikk6OQH79KpoZ4k5/P46phOldVf30rX/BMDX9MU/qdaaasp72DiuCeiy8zZQ7pJyZ/Gdmnn9hlDx
zCraiE/irvV6Hriocna02w47hppU1/PJLm8UH9FfIm4zirEM1E2MiwqaXj56rp3eoaH/6r8HBY+D
SNmD7Zi3Zvsal9rtA1bN8htAHPGZPCOpTDxQa8icMIJjpJAe5SxchyHhYChIIXbnfUFpq33uIUMu
jDIFD1ZhGuk+Cc2y5GR+BzUb5Y98+mXXjEJE/xvnuXtBZHVFDJBG79ZI1NhGjJDmJvG0TIddaQ/d
pNwo/+Ts0l6jyZtSjNTf8zaJVp3+tkbvHrBKV63uAT8oxbZ1CdpIU9G0NCQYn2xTcn676a2p4K7u
na3He9Rp1C1ffY/prDgu9tMwxhCc9jHPhBNmdjjoctbXkX2RBGVB+IoqNK4SREWK56qGJ5W1KZ8f
vuaEYIkoOFFDnArTihQlZQNof7BOiUhCGMkhtdadYiBdv4JmW01g3go/OI562k2QFlICusEt3D83
Sv5zyinR75ZpSPK3MuKJf7BjGnFDot9Mg1PMTTUsFJnFqlfxVA8xd1scL1tv6brGiX8oyjOA7gsc
qAgQdKe+BtLLQTsoNLCBCp7A50Vt2VSFPxzzuiL0luZImtq2N/6my8lW+zuuATXotPMlaFp67/GX
DmOppaifKhsduP5Py4YrIywb4174Wv8qe8RyQc5AHl+g6yWlT2kTejzGg3IWIfJQLyf/jEGWn3ko
AWjPPSFG9os/K91fYBl07FKDWbRD9pG/kcy6YiXQIkaEXo0OAd2PxYNdK1ZxeOlnd+OXPYhkQJyZ
zcugNJ3HNAJK1FKWkwt8M0fXskFC5Ti924TSQkJW6fXbZD7oGtKXNUA6kYVHYHlWjYe3S+n27eNR
db2lf1UIqWiUJYBNZ5AFm+1/T8HspYM9W1F57XdT8vV6AUhw/G+igpMI40WyWVTIc1RX2UxXxxu6
MOXGTml9Qzytw+OOGxqczH2g1GS2xQHJdUXT2R+pMos0jiX+5ed37wgmbVnBe7D7yNGlkO/VJ8QO
rE9mwwCCMYwYjVbvLn24HI5vNPUsPwxjRde2+hWpFdmJt1nUYgWD/Gpox04P3mIZ+IIY6d0jnDin
zP5Oqfe9U80/wShJfZIo5QQD/S2ucu+H+6QgpJc/VVKaFpzy/W5SKpiDSyh7TvOfDTc0+Uht4x1Z
N9YuX0qzIwdZPycfYcabZSmqKNZxwZRgK/iPUvbdMGx4MtZ5Mfr0b6R+G0jL/YqqnrRvlJCoD0Sx
OBU/iC8d9rELP916jqxfgzKTx2u9ya5aQ+eejrhW6p+QkQ9YA5MvhXsF7kSNpcehlU0s19531bmW
2XxgqCwpWZ0AdBNvJs/whCqyUShgRUh+tFczV8ii5XsJ31m4EUZnfJpkxMXzCNPmU67Wqh8Jcpjq
QcXLo33fCzRZKTKth6D6Blp6au1LD+vsAAVWtYMlWIqLLu8PRAasvSk//gY9jx1WjQq1htMJRK3C
YtKNHPrroh4smPHXuwCILpdiNe9Q/l96uZRKZnDaKzDj1hb4c70LI0jLbnSknKQUQWePvkE4bwE+
9ERAsg7Rsw1+PiktEkcVTquRxAsy0YfkwPzOAQKy08wPPABDNj0dALDhq8bO9Zo384TGYXzinb++
UnMcpjPC8JtQWlMGPFQXEittwJO0keFDLUHucBWbZ7xotri011v6dQfLpJGOfUM8MtMMQn5b0p4o
8wsD3d/oOj/7Ood16VmpnrCszoFzd5u2A24y7vIZ8CxcNiJLgIPZSwLSYSvjMD7yiQMfHz59JlRe
G1crcFY0BtgBOIi5H5FEqEVqa6qlDVNgTcFYTmY3YkgRwyCfjYGOBD1lUuvuYBPZwedZOLavUTja
BYyxowJdHHHT3wrdWGZTpRodHzo0aya6kmyRpeVa8KkiHrPnYqcvPYHZyDTYmx/T7XFhp8Vf5Jur
fQ+d4nRr0Vw++mPgEEjxHQkz9E2J8ten21UVcCsQVqUGFAYqfdK++2twnVi3H6eXV3Fj+2PyWE6a
Cwn97KM2HOaOdqxlXJwEcAfTI5FTAIsJNv77WiQpMkpDhMWwE3iI8IFDyyVWTr8lEea2yDXj/5/O
NhZ6nNzhVK4dHFBXsa5VGYmj9uVGSfAHdHRhpU927NXMBeemoghuqGFAmX61WFsei/Z0STiCKHh9
gjXGZEcx21yfNAmliHtGOO2FQ2BTiYmbKCUih8cM8npnGi4cs5+jS+XmFFhIaJ3U/bx7VxfCyIkW
oOKhVVYn9sBUI/buVAbVh7kY98bgDhazCjpAKaGANoWZWZZ1uvHOhG2eXEgAkVAEI21yyXYQCwYI
xmOSXRbKL6faCTZZXBt3ttDGBRr9LFjz1DNFPGMy+VFIrzzwCqnj/hf49uXd9hoFA/ladi1tgshj
4TEMspjAQ9yu+6w0VLH0ASowZSqHh7/lFS9Uy8UDF+3Nn4FF4dqYLrNhs/l6nZfPujvJ1CktxgTj
koM95NEEP7d2p4IHqv7FLDOno6CzKogcV5Q7yNiWeY69MUaKVFlZfNF4Ih31Ufgp+ZX8wGB/lRsI
b4hIK6qG73axhUKRxwuC/RJ73PzCdva/rg2NgCWWJA6CFbGCBRgQf8V4712prbY/K/Hhag7bLkZH
bN6C/Nf7sooGwDJaM1gT5W68ypMgF7fLjx1tKv4vXl32v7eD6iaUgUtkRi0hnPM9eUIMhs+Wf8W+
Cf+/NIzK9jwLpoGed82uOIXskKXk92MCNcE69UdLy/VX3y3T3ATvlzvMHDg3sVlfL71cmrZm/x5T
y3874gSRYayCt+Q95e/bk6nhGefHKnaXBgvxj+/M9HtWUtOYSqhV6RtubKN+NF8tSCZVVHXFEsyx
vSp7rpPxl/ftkg/P3aa81pj3p8lDsbml2wktXVqZj9S8tQnVTCfiPQ/RfHyRAf/KVcCN0og1rpEy
djQoL8QgTAa6tFjGBY7n9kwnq6DzjXZ95KbViSoV9KL4mPuFSlwORd86AoEp4alP26qKBVEckPlE
qhqOeGaniOAES+KdXYFraAriSvXHJKeMHbhVfh7ns0DFi4QU32nOgFLzpodtalvXa33vF0Y05IdT
P3byDhdg6yfOCHgepb1EAnmxKq3IeR7gHlTeTxZdafJixGAEnJXGAwUE3jx8oSOVaa09vL9ZKdik
7E1CCjsHuYT622IETP3s46iZlq0Jfb2h9F0mDPnQH+OKFpSrflXwZYDBKcSal6Ty5TGFHoJ/R6Td
FlDJo2s7OUjPpZTObS9lj5XfH0cyduv8hwOD4Jh0ftgIj4IO+p7RGwrW3NPjw6eHyr0kqA/0YE8L
4HmkTtDqPCI160n5lWwdsjRxiEe8srufZ0c4tBhHmTlj061Rhe2lhvFQYMvmydIXKklGt9Oju6Im
1N7CDN/xuPopXWQiccWPVJEbCQqcc1QUxpI415zAtFM/nRuiFJziiQ6K2mTCh/u0HXYGDJweu0Dw
n5M4UVZfWNBc3ZUR2tdzULgaWchX5xyPycqMIk6rt/Qa5GZJOE1COeXk0aMV5D5mJTmyf+oKoLBR
1Q8OQ7P25Pobqbq/XI4OPZT0Y64f8qj82GJkud66UdUHNMoVaktVcskNsS1UQ0dH6x3Ziew46oHn
IzVUyB01QQ+8hiIE1eanU/uZlEiDjM4BmxJrmWkASCc+NC8510fNDbpyK4Yn6cgL/3tAdAivJt61
a9Ax4DskPqQC74dwdrrL+w8Hj7fhcgJhSCO/ulujWN6/Dy9lAukDn67nwOQ9vMaxZfoY9tfuxtzz
j605sAlbnQYC9WoH48nMxFCyVKTsQW+uAJo2vx6hHlTyNTo3LG7mcFBvntDZjjzHs4Dfwe+TEkXo
hcLge0oUiBhhmT+g/wBLPkB8rcSfpLykOphh1foT2IF3rYVp+JBlG6Jh+lQM0p6n3wY6pEZoLt4K
Fe9ncdPaJyFai1Yjef7oY1HL2baSy2yG5Su7DVmDsQLyGJHVO5fjVOLiOU5N0RXz2a+9m2OUD3U2
+E3drTM12pgew+zCOSZv36E3uRB/8zamN/k2yDYaeEUfk8NpDRfeYYlu7tz0bey2ocf9b0+y5E0U
0cKcYsoXv9iZiZ0y+5VsGl2p0DRjISTPD8mjiGnCqnMwyrw36ktK6cjbgTXaxAuCWxYBzYKzRl2F
h3+aFS7oJysvQfKsbyCj8gYoA8QL0Eu8UJysdTzUOVeNq7LRvGAPN4AZFLZhE+HcaY37FYiujWsz
iQpTP1ldlJk6JdKNiRqbRgH6melAz09oKsQINNSGKmN/xVH9zVM0fFUAksp7bkxEJ+YEPlpcajCY
eZzxnSqcAW27M560DBHEqMLbd8x1q02zJOz+0dh4cfs1pqyq9Vl64wMjN9Ia6bBjV8i/imGRwflQ
PXtzWEB12u92n46x2b3FGQGggYKPk8Ni4n8AGfU+wWtV831VnY7T43SkUTHBMsHpniR027uU6y9N
1EHWy0f3SVLlY8W3IY2Uk8/AbYgEdZ57N09yVsfjJGIQOkuol3WoF+a8q4azVPvvzYV9+CaO9hiy
AK835sRd/4dXVGmkURiMoOMz99u6MvFliZhrLHMknWwIM+INay08C6KK7X8QEW95ahBWywI8NBjK
HuFnhLWFzd6zFCALp+Q+VdwXHmW+WIGVT2UTlsCjnhfffhLCDAPLlK1LN/O/Y8SNPBId8kQsms2/
DkHpR7OPILkh3L9j/oPaT/yTogtMyaoxS1+NhWoNzpfSJD3waip/Q8LQQyc9HuCy3k3vDO0Rjw6l
Zn6nXDJCtTQ5YTbk7INzxtvaJ1V0edLDHbPDHi6PZjdyxI4iy3vJC/Yee7IX/yT9ZF9T+YBjgYwZ
YYCbKfZCEktrZkKFypdRvCIiPHLATh5UKhb6ZOei1qA0UkuQILyktZjxIcTVBgtTmI/Fjhxk2PO3
cazcRFblzxYvBdxIF4lM8Drcm5K6JS0lhXWAFjx0uDSgytgfEmEiAIrwQCDzs5u821CQL/3evShw
isECTAqtvH0Gv1mZHEZGmIfaqYY/VelMyrAXzE2RLb0a+vAJeUVq03AcbAVHyUlnz9tWSoFI297h
8UFEhCNwOLiavE1HzkF1dtWXdWbEmoH/0fmPlHK9iq4AC4R3EuJNtruAxN7IiMk+hk5mvsVMLlHu
9HYYoYY9ZR4osbs4+16FDxx+iBWnvOgxhRtLqCyGtklJHiO9uq1eWCoG7TwPwMyFQ+BJBDJJkbv9
KR9tLzbTdyquDaAgYFQwDACcBv8XpH8hBxZodx4qgYZqZsnOzS8unqGd7YyNJMJ4IUw6JHQ0sXXE
gKhSwGBIHNc4u8JMuni/rG4ObHUxiSpJeyRafi30mxYhfyXpyOChDo+rnbxZ0DtEwOUj8aCkrgsj
u9mE303dOugTtLP1XIQ1lvZ37fCDWy/MoROEzaiKiJPX8qfI0FAL7NaLTANkEjKA1NC/+jP4dEK1
IXgyy2WLjgABc4s7sQ0cJiNg7WPA2aPb2WUEq7eMxhmJrW2EB4wdli9DQpXt5Ekr79ePfeiXqBRl
9q3N9L1G8Ix6APcL/oWD7ccvswgY5ZogvyCZPeo7PF+rwnNTfzmxk2InB0+eAvxaXP+MpjvjXgUv
vEil50RX8SMDT189rUStzsV8yL5xkZvfhRA43EXs5cksRqTkWtl5wlzDLraIBPL4n6l2IgX3WQ/h
eSwdtqnrpbcZBhhVVDOQ+D4VB/LBQ2HqGaPGqcxJ5PAQU2PmicdOxwRH4SlWbA7SVDA5sNxiI/q2
qWemc5CkIR1kSq0bTSvE9uxpqTkcJI88uU/1j6Tswncdm5FpD2+aW5MJdcb7ZlrkQpxSpy6nwv3H
uuf4tmPfH7EIsRgewvB9pjJQ/TJtB1652ynmvZFpPJkkGeHC0apO45XEv8NESgB1VyeUnJGGdFky
afsGgzrmt7FlB4c6QmDcDWixpG82hMT1QoXHJc1LvMmZAU42bnwX5+MspwsFFZg2/dgMWl4Q5Hpy
o3eMtfpB4m+GVFgbabZ30+nvuUdK0fSf6txUFcaHI4O890+epF9CXKnnS8+SRCLCUP3Cyywf0ETY
QDTu5ZLjDLIqnbjtWt2hlVY6XwiuYbck33Ym44tD3WVSfgy2TDSe5RXUNjpf0eiB8BCpnFnwX6Pn
0e4XZQWKwJmh4sb/zf2h6pBJ5SahyODaaAPj8sCIPh7CoG5YillZxJOuHUEb3cFCNLEQ5qWrrucK
VdPqk1RWnEqMVArvmrlU5TmibmklC3bv9jTQhKW9ATMiRrrCAq2Fqr6ZLuqY+hTlvfnVyTphLKq0
XJ7VdNVZKUe7fK3PEMvh/phnqU2U8kHb/n+j1UoKNMqPMuF3WeuSFy8Bs3Xms4DvR6/iQ/aLxPhp
KvyphNtD+FDwoIs1xSdKjwZRn9KXvDR2nA/fw5Z8Kd4MkTbPF09orFokihR14hwkXdRspIO1PcdB
udzdJhNjnJfgN+WXsqJqLvjzZp7SrJOQO2Rkk0w1TST2XM7+jFQ4rirQL24eL4cf8HFpqCkDxgT0
U2YsISD7Tems6LN4tq89Zsp5newHkx34EargdBRoFegSbNCQWcVkPHSTUl8h7YfRa8qZzZJYjl7Z
skzQMuJDM2Jvdr4hv00QKI8PBq+l6SbviKu27cqAGJTpWPzMdBQz1CdnCr5kx+nGyr7hbTnrxEWy
v+Fy1FPWiEJiV89fJTy5HzPOl9bQRTMpAjZBZa47ebZFMNXAU4vNAKNAY6Hoe4ydaHbp3D4hv6O+
HL/qr8oJ0W1Zs7ivRntj0n3FAHGTTf0wGBckHJzdoA7hrHvSi6VLqEYDX7849o3RIoUHAATXcrRu
oznc49w+lzcfu9dGfk0y6Zk838r8vWCMjHrLGT2nrUtqBZrVYQf4ROKJm+G15giskyO1TMGeERE1
7Gg5WOi0f532ypGM/WrUrur5lUzEPTJ22ClZhfTnykpeQKgru6Xad3nM7Yf4RSsaXxLwAIZj2fjr
2M364nY2oxF2pALwY28ZET74ZDImYDwgxYhjedYFep2rF6tq8hjSaKUQhn0rjJqCB9Ip69fQYrVT
xcnUiTSBgE5yp9bFe9Ga/+nDu24AbQESVt0a6MwUgl8o0i0UE72ObaDZKe5yBMg3FiFnrBs2rI8t
5pB26LiMtFXJFV89l1rClVvLeLlor1X35KySo5oUhyQYLV56Q2GYQB/ZkWHNE9CnJFDwjk8kr1MG
huci0fTqjpUhIp0yeLmQhlfIrRYpeSzIHnUO3h8cTUemo1HrZavE0inebMKmsrgF605x8EbZurxB
cWzX5RQr6n4euGFlWyYMDrZGQSVYqz3JT8tTVuLE3jez5dXBDP1i5UsS0kxXRj373sGedaREyNiW
D6fGZpFyZiLoS8oyxxz+3gzBXCokoe7Dcs87VlhyN4cWmqHXJmHP1J0183U/m+UPSZo6UMIkDnUR
uRcqqGZMn21tmMxE83n7SyyVno80pwfQoVObakVh8ihCYgAYa9a7rbmiY0MMNupqIe61dZeAfvj2
zqKwSWJiRW+5Q/zuUgea7hP5jn3bHc+7TzAUaB6pTGkREdKP6hBjC5mZxZwPCh547+278yvF7P44
BC/is3tjr3iTq2pt0tQgCxUVEabYJOTRkeMQDyuvFXrXh5/Ej4Dct4FT2Yx/OqvX+XP93f53dp1c
G2khTZJe9q/R6KekdTurWagiWnBKBp4rbFCMp35GnQ4e1hXGGoMqiKWzpQkEVehFKh3b74eLeKLu
XoLtNftlzNCOl3r8qiFjOa1eQZJwp1708gySAVYweJOElhVMCZu+3pkmoLwuOl5LJ4hRpbBS5K+M
CycHD5xaDLTHQLpQiPQqMT7aqo26bEVkCWWTtJRZrJ4vBo582/WgWEa7ryg5FntqQ1wAmk9iFoPa
ceXGUfZTT3uHVDICYOWIuMjGzRhUvm2Ovmt5y/C6aMz2YBuSEViPoV6PvitX3AISKPQdVjk7QqyL
ZWBoMk8g2Kb7ztnT0kMa7rT3SqqpUe2WuUY4uRoynLiBQiT4tV/r7LkW9t/VOUHdp1143pym5qjw
PKyHgrxpdEg6kG/xLgd+oCX2TTMBgSW4TXy9Ugc8j0GumhgfrzTjC9Io4GKnL/UpIpF8I1JGoTJw
1X1ZIZfNdRdKEMh+PxjGCR/HYgNvIZlluEDcnhA8WZfn7kgyR/3lchs48HWYsHcRDVa7OSMNrOEn
VFe0nRLk9oq/Rz0g57Hg/OkF+kIv6Jg4iSNU6XsiPmGOnDhpHpakM7VWDiqvpjSooYg04DBsgd5W
+owdfgiVmti70krZC81G+WTW288aXUDpIz4nAYra8CC5FIDlB5A9NyIwdz20Iwf09t46w9pizuhw
y3f48/gRJhwJbvRaoe7HXCX+WTw7W6EjRwBAR1Uns9vZrr7FQJ0mqIvKhRCFYveYJ7qTj5h9rrG3
hiNYwKui4Fn1XEFNsYabtl6qjLogolTSHQ3WQlXK9wKXowwt9eKsp/bmmaSgTh6zFju1iD8QpbTB
pHUt8/Nj+MDKa4Bfd25ehiXItRaO3SFjoZp4zsXl1GunXX8/FmGBESdsi2YgsV2F9MbDnSpKl11h
zztK8f6THmP4PwI7nBXV02ac9Ue3wRjRZqSwUi6hQ0GTgiwJNLgNrJXRAezqv7FOc/uo05k9xe8N
GBpIdLHVAhKzozX0zL8+oeyMCeI9/jjCFTrdRRr1vBwKv1Um1w7QPOw8d7CM2t4dQFlmKMk5jSO7
0pDyKjDWfBpMlozSpVCN3723WcfMYBzHhpS73c51tam54ypQbU+97ckYJNettrEKQurQ5h1kyze/
2xbAx4EQHnivGvwNYieVFZeRoSgj+Q6w8Xnh5BlEnTgiH01clpEJFezWK++mvqK1+JJCCFnP6udF
jPx4ThoGRHbdpeNtfovz8gLpqzcmSdUMKXQjv4YyUmZ7LQCcln+nkNrMp29ag6RTx0dkKpxtFWnU
pcKNmUmIjnoTYnvm2B9OCZP9xbJfFuczaHBx2T352PNfoIj2xCILxEp0J9thBZIrhp53pfxQsZSl
bgC2D1Hf3OLm078QSIcRf5kI5OpdlWXzSPV0ecxwQxxGqlGzABg977oT/A9LQcIzWjvIX4nF/yvT
m9yc0wwpJXNHq9ZJEEYR1D30rsiNTTkWvpli58/xSVTorH2JRo7CklTie7mQ0yD9OFJJlINr0MtF
zRkLrx8yGeP+oKZ5tLLckk6S4cjEkSmfSZZ9Yp0DAOEzwBm1WZoTUOlljidrNR9x9oNjeXQl8CYu
WrWpLjOWSdKsoqCekdzAXzvAjnquiOh7EdiMeq5caNhmzBZaNv9NA8SFxQtA5qkqXIOIARnO8qZ7
r1LgN8JkCQprL2J/eUteTixG0ETnz9C9G0k6spq22pOsUuo0mYUspXgECmsHZzMlaMJLLVVyYfqu
42QE4nR85++48FQcNlXJPekHVzyjaDZofPkZgMF6KolNEmSPlPndR7ojf5qbAcuRbz+f7GDWSZ6X
JDaJxNWR/rncX9Fg+u/zi7txaPJ8MR4CPGedoQzl/tM+XUT9X0t0LLOWqgDy0F+V0COOfMrHmw6T
I0xaPEVj4e6K5Gsnh1v3S2ckpW7aOm4lGC3F3ajA+WMxCLansVv6R2oSJccaN4fZD9yDBqt6CEZr
/9AZTEdPx+b+Fb6Io17nungetiZT1a3IttTD6zCMHjukn+fA13aCLvdYFopCt/7QqbNzohqqbt+Q
EM5LtVDXsZ3ytMDuJFylZi9IxL2bBLgqsHri93LiQek+UoZ9oIS3TY2Hb1hdViCG2zswIGvMw1Qs
Ornl3sT3nHcGZJoamZrtoGdnVHoH0st7ZTT8rJH+BSVWydcIN25TxozT5J8D/XfcF2w91g7a1ZI9
igp72O9FD+NPXvFDOTTHERF/uwfDvUzVOAXpAIYaccYJNysJlOWZugqCwq7kfzDXGnm0mHp+PDTM
323hbBew7Nh+r+W4OFG9NlkM6u+PEryY8vEGBQ7lsV2Hc/A8GsL7y+rDG21dxFp5nV7mS+mIAGT9
+QKG9F/nBx11hakjm0uQvYDhO6RqfjoxVIHB0xuSmKb1t9CaTWgHTdHIiAM0X317/dvzGeYU04Ma
IeUgpXZUEli1kJFCjjx+e5ea1fRmEKBjJy52/VGO7qInqHvwyHWS/93TXGDDHJmzGmGu+8z9y8rD
xP0KnuudTh0hjY+lSmMLmtnmVgutPFdv9HIwI6ztTRqLkUwUx5ClH0vKy6ZggpMpsEmcZKRA73Rr
2QBcYgSMip8WxdRIWxiEfEbPtL6r9rxs5wJIHybGr6a5eF2b6O2eXIxM0azC3NkfZ0RLTenG1lxm
NikZXs7vJbYI4nzOJcKQfRGcW2hmdqfLVgvBfVjBlsXzF7w1lUrcB13mbiphrx+ySF/p51eqZqAv
Mx0XE5uYfuecURp4HcofchUXk+DofCW5wdmAr7cfEFbqnhguQactulpc3zfTkoBBHZ8vcUuKMOl5
VlVjMciPq0Ps/aL0hgEZxcn5WxTxOsgWJ82muuQl9jJYSDOV+ySKGmsKuZevwHuXhhFaePAgO6Z7
3E3SdF5Lt5mCrY6jIs3SqOY4SRDIrZvVHv5KNs75POXv12TVNMdd8Zn0PJqmUcK2hXwuPkLcml6s
bwBanQiS9DdSi/w0sQNYYItEQ/TSusjkYIg2UHib2t5ZGPo7nnhij8md6PinSqTroRVADKfjwfHx
uReWUImNMtdGo6Maep9JW8AsCnOZj1yhK+c4ChtO5RJ427zSajVDqq99OXAFiz5A2SDeS/6w4Yis
kG4Mr4zt9Lpvd3l2W559S28vG/scbsrgcmoKzKXfxgdIwjUcqkplPjXFILdBCbLBbaDB2WKOpn2s
1PI9KRCrCkjarr6yZdA0TK9TcaBh6TxViOBFCqlThoOKoSRDWz4ZLeIZXahYu/GMYMm44DcxjErG
I/35S8jho3pe+MTjGiVVey4+oejcwE4AhFlAoVD/uCozv7EGGHqv4gTY+CRdXzOQp6Yy4c45CgLg
xEKRbZ9HkubHHs/7K3P9c7lg8Oz3GvjoiJ8AibxX2brPQF9DVoCPrEQPvco8KaJmigztq4lGGfeQ
JPmnasu5axTOvWcqoe6tSYZSQZWi7fImICH8PPurbI50ro3Yt4ApFei7n+OPb1eH3Vz6wNDJB2Vq
nQYVBAM/RCRv4LglBdeuPByt3GXX+oARWTl52Zb2u9FnhMEi/ZaXya32udhSNf5MhQTdsVoKm4kN
TXMIwTVg6IkdYxKtJVJMEmZP8V1R4gkPFoz+vLtcbHb6t/Cor/qLirPMH1q8ARbCpiHrzZWknMOn
r4PyV1f81lEIvzOgk3sV4bqzcJNZrhSESkbJauuLL6H4CKHXBvbq+qX66ZHh1YYoflX5Rfho/cn/
iR78dxWXfc850HwTqhaStXp304XAC6lb8q0vph2K5RgkTSSLdb/YMMWGFJcBBq/5DFCi9cqnknzP
m0U+axqWSLtsYQa9N6nqJbCMsc51LKUDplR6F1oX9bmLxr7dnax2IjT8neBowmxXIpcMbAWWVC6F
LJpUS5bFnkgM+905Y1L0EWyXDtYJ7Hz1hamfevkXNfjRhJAipuS7DbxhM9W1/2Sprdbm10c2XA7e
mSx0kZPRZawKsdbIcBzzihzbu8th4CkhrfjpGmUONVXOsv6mQNIlsdzJXameVFW8d/hbOQqL14+u
/QUtjJI4ZwxO/zFizhrn874xjeX4K2KcFryvK6WzRS/eE+Q7sJ65Rqzh/g6rHc/cxvhk53aG0eH+
sUgTJgwc3CAOf6ZZH9Z/FXOpcReufWrpxE64GWNbIe413fLNoC46NpcLX/4j1bX/rLfS3Gdj2TeP
W1TDBczR/lTatbvg7zb/kOdJkAOQBH4crn0rSYoIyzBO17QV3VUiVoyKhd9OqebuDlFkNjgQU8wO
Ljv+uVBXe1yAm9CAtbWJ4UelAi+UWUJiVzsYHVlGkhapLYrB1QYHrfUc0DUr0PejRyYQxGpy4+0c
8g5I/ECT75sE4n9qJWLClSCL+48LUDKEaJypMRO2zFcb+tKEd8iYkLrP2iE4s1lO6rK1HAdCYUF/
bOBq87uEADjDsT1v7NLt/1c9uJ4cdGFjeci0YMFWdvFzE2EgCp19nvKaduoo25uvzCvenzNw14Zs
Dm+7DORJXiBjxBpfH6bsvr90TGhr7OfOsRyhx9DE1rU/Re3yE8dt8xPB40EQ5/LzqYeZpEixEGkU
RnXyoCvmcllMqDBJ+HgoGRZQZJjGO8yvj77UsuoEwDvwrbJ/ZQUui8f2XrNfuTvRCu2GL5YnKyCx
5qiJ88L5BMle4zqWAST7Ss3aAXVl0QcYOzs37oebG39YTidJzX9uVuNxx8SNDlApwQgH+HCbG+7G
5RAOadZB3QP8Tsag2MHpkErWgCbpJqzwITTwMd/wi1bfPM4SGRjMU0LKFNZzXGvQtjgwQyIRz3cc
OEqSkKnFbQaJz+VlYMPNp+qS/aQKQiuSlct46vdRdvrRIllfkOZ3EHUrp/BoO81A6RjtBY6waHWk
irVld/Ym5x9ChVs4xec2JsOJuBYUyLSLs49Xh1WGJohMZcwFcyMmi+88LP4dVEoaTvai2mCY6Ckx
tyQH+nlPy5Q7IBAFYXMMwimabiTaZEuhqMOQNzMLM3zAvpEyXZwjOpOUFt6AHzykSoIPIghzPkiz
KE+XLpXRarOPYXurMIlY6mWNtpH/Og5eSYnmKAJ4cKUUNfI9OVG9Yoqz5O5IzC30qA2aWvZvitOK
sIRi44ynqcielId96aKpvWuySC96Ix85RI0DL1oZtDOfT1XexDr2ABOk4XPnvOsfLI1lg4cscjdh
I5Tb2opJ7JDib/th9EaXffHFpwAE0Z8o3noB+ntD2Nl+hgQeTBCNIZTt4LwdM8stSIk8wp4ddbUT
XfbAf+UBtf4Eaq/F2EhhkcXiMS2yvWKjNwdg+7PuPwGLIpD7YPv/neJxf22Rf5ROFUJvC975l+hV
qvO9fdAtPenYv82+Y7WFvKcQbvLRu8suH4Y6vwm5indVCge32GdxOx0CjzoolIONXL6doTmWbDXx
BbW+Zdd2pDkBIGoydvWBzCKKRirRkSBPrpI4KcftmybsH5jbK/nTY9R2Gdoj5OjO6LdqsPxiS/MC
76Gs+Ua6tA/DtOFrVZxs9LUhDBFBA7S1G1V2pRcjg+2Ibe79Jn35zfbtO56bX7X0TGrvKXDTiP17
LrO8Z23358c5IStFwKwE5Zx+SDkLJQpDlXrDc2tgyqXqkZg5SqKnnMgNABnKr/rvFNtqLBUGBpJ+
FV2MYlboo1FENuDWrDbfoYX/0umMi+XFK77pulmwUuBxZlZwsfXgJztXhPzxBBk7C18T4amJw2G/
5pmT99ltQdKUQEpSvFMrmtWnLOMbCsFqvjNpZe5sUIZxASGwAn9cJOXyPqrQv09aZH733E9cBeOJ
zdQZKYGxUXiqBhGr74yrMtJEkWnMLLEyPgBLi/MgaOQWohkXXSjyzorQd7chKAM3xqjHze8M47TD
imOR4EbkzaV9Rl5NSezJCV7+1oAWTrrVxPuPCTebh4NsL2HMKjiNznQZvZWw59jFXSH6ekVA3l1P
c8uzxFUrg1E1r0poxfeGOSX0jTPcXb7iBUNJPxkFeRLNoOjYqwHOlXfEA0HiF2rgdXkool7cfhCe
HFa//nIeBiOpIchfhRW/v1SFTPR3zkzKg4xIDfzo85gP2aLUeFNtk063MN36t7hWFdHg7Q6E4ZoD
ky7JwqmZYZuugK0NwavSnEyT2Xxq4u0SMbB+1QMy9mt9k/kGHOTKsl3NiZEJiUVFqopuIE5pfH98
HtqYvsz5VzONTcrLqIaj1is/CCaHt6QSvU1hFuvV1V1G0H4OPxoDBy+ZMysawvnc+r7kC8eb2aDE
myV8TzDHfK5z3hGA6AxfQZXVXATVenwQFDtH92arvYyKWoAV9jd8JvoMhkNEEY3FsYVbW/xNEKnM
kAByFlIwlRpNAvVIHD8VJMW0SCc5IyVJh+WOmg/nZ126Z4jRHdkT6Q3uk1QVkdf97Ua+TMNK5VmI
7aCQmMB96lCJwOAorNB6x2pOu9+khUBoH7x+As8rEMKoQDiRalwvnqCqsIWkX7fKW/YGBGN4tWPX
y0c5V0sjbzMm3TtokNRBWW2fhFRKM7PLwEmzZzNQB7c+xrpCBebPGBNUIDypfYJr5il6hcPMYKVw
qpbtMK+GG4QLp/YR8Vu5reiWQ4z2ImfIqYtlfBihIw/0eJ5FaxDOLVJ3NGpJfmSe7TUxFUQhthSf
sxaBzYZoash2kxnBYIGirh/yLeKqIq365zfHvy3P8H5licbsyNI/0VAGS462Ohbpw3Ep8ic9Z6wg
4XycYDGyDcDAPgIaZVlk8A4+LdLP562P4x4K1mXnv8Pf2WO8iQUSOPxEPDCngU7sV0F7vhRm2GJv
qsb6bjjJuck9ChUh9kLpm/kjgn2GBBbzXQOLYDTVdixILVCCXEkqiZXpaj0VbnPSagbIzJ1Z1vB8
rCN0d/JivcXHKiMstSsyf2HRvckuJWQ3h1lQIM3NVCm7TbB5QAA7tLLDvrAkJrmKUwOGxKg7CbHs
QW3ESfNZug7eNwkgZuoRVw5pSEtrxx/ZioO9/bczTkBHcgXswicI+xsQJ8k/RXwPXne0OyzFA8oe
lB1tV+A3+knqBom0w6GfS+T+J5xrZYuTeU6GJ9nL+z+eWPRskF4rwdyzD2juMRq94UptELpH6kOu
0BLA5j2Jl6uUUnqUvUfU4sg+G7f1hnyujH6SGvQqdf1IF5RvsWJuGbCEVeEXqjG2pjBdqDAUCASr
9ml5TU5zpD4APzMRdCt2viRafrKQ6sgYspCQg8ReorI8wB7i+fF1UD1KCJx4hPyb0prIzCXq/q6J
t+d7EYYt8T1deckBWNSZiRnzYzbCURx8KO6c7exjay59hL3oWkzJcKQZ1F2aeKxYgH2E0mzvvCrK
jt12/1g+irxseEw4+p5tOx9nEfR/Gf9s1DA3/EG2tth3nkqLCA4FzNuyvl76EX2WAMD0rBxDPxNJ
noiiNBZLbRpmnhJGmEZfVn/bnMyeNy5ZfUukgko36mXAPWaqccC1spmuQ/pA0trxLL/EvkqUUHzE
hijjU4AdeqZXTcFHsoHbSBZzyoOSpyv5lgBZusXVXtlxooUDlRqImwwRk0EhmoPdEBiEy2elUhi6
CoPZWt2PXhLVFYLkQRI+YKwLdmHhlOELhNqwSe5iBCvplmOckpkvrwkMNgv6343JDEo6gD2OJ2N8
NUCwzrvKYb1WmkX3L5+nwwBjkfuQgCNaHQaIO2JI3y5t7L5DKrPo70UuSpfcFo2Q+cgAx72zDy79
aRwWwaoKA1cOgDuUx21aGySxYJ7vm2G9ZGxVXZ4sLzTG1YdMJCgqHFUbBo0DlqiW8gSY9GEkyM44
BzvOH4afl0HG6z+XJaMNzR7RRH+QAxp2AYonhPFO6lIgf4uJ2LXIcn+E3s2MPXJPpwL3yUInlCZg
xhQwwOOwbaAiQ1Of7OxZqTEgjJLjTerCLj5UV/KM9IP9NERCXl7KzAD+/Ya/LZ4D1iumFehpX5v4
ZLkH0A7khhOpbrn8iq5wg95TT8uQmIGsuAY7tvZM+2DXuqHJGKWJBqvUEGmRrDjHIRhsoSc+KUGT
uJarvnYt6lmP46BpJd0Ab2sEG6tW+VPJBkOMbfSZt4xmDfLj/rzELiXF3kP0js3cigVP2YBxsOPD
o/O8ws4UK86jM0EkjMYbDvJdrwc8IILiEDluXyYiBrMnbZ5R0m1YtWhmmeXdK4NASYM3eOXjrAqw
gq42qEIrzNJNaVx8k1zmLZ/LJLnOuFDzRhOHTbIiqf4erH6S8f9c1yhXWchA8lIhJk+orQ0kJWW+
mCwTbNVfkwmelG9kq2EAKhfBwVKxtuqR6TQuI+4GBNX+/mivtg6uwn288SPqOCXrvnkEGXdBefAl
toiRoUOc3xOd+4N4Q4GyareZAvqviRvgtWpQu2TaSInZPN6gQh/3OFSVW3kHKGf1ZkIxfvvCh37v
IwUJ2imKEoCQCJebUfyT8X9qtOlaJU2CkaF1TNhCrvbag0Ga9V7Fm/rckOfbRwC+Y3OB+kirW21P
GD4AyVRQ9/bK5SYtZB7Tqx+IHyaPonr2JvbNaLq9ILlw8WFA52L/0mL2MrgmCfc9k+LpJzp4uX0e
dvrEKFyGQTbb1vP4oMdMvhZ1hAYNx2H77fx7e045FgEOI8d5L0i8ikQ3XEFd3mWVJj9VRzMp1Fmp
qny8oK4xFfzMWLht6LhbX9KPYsWnA3jW9CbsgiKq19E4IVrANEON+YmgHyCtg5YHwEZrQyEyPnFQ
w39j6raQvvYEJkzrcBIcxoMcE3BHjt1gvz2wK84zzcOL/spzp6B4iXwbM5pKTS81SkkfOXHc/avP
M7250pYmczrmMME0+l2f900ChPj7/Oi0lqr+zlNKCZ+wpU05vZqYLToezB1uaD0N8DANNK+6ODGq
chIxuuKYK9xhhivIJOmYy+NYV70qTc28EKOuIJh7rurURlHY82BHvPtQLkTGZLMKFw3VvPKvwnmy
TT2w5gN1fU7XtrhwUZwYEF0YyksnXemiZ0BHZrzvQQ0LCR2ZderC08SB+9RTKOeiPAmOO3/EAv4q
BNZ9TgpkGRMO03MnURCnRo3s0qmOZ0K2lePDSlU2S5tVhRdGbm7oK17Fh3UlQ/72an7IaAhAVend
5AXwD1H67AlqjLrbvd6aam7viQ2khZ7HXbGT3a8GghZqTP468+drRlNQ0AQbwE0j1SzqYzRZ3MfV
SindsqN8fO90GjbgkxRNeU+55znH+FyhlldOoxKUzMiv5peLW5XPGEd0TL8XbOz3T4MGKH12V57P
cQkO7AayaI7ftKb6I/KPDFJ5/WBK31ewDDlZRda5amtEi7amHwQd9weDX6VXqJuJi7lyUGebGHkn
mz5ynClSy+zWhEXbii9+vOSEMk7zoLgVPTd+Tfr6c9o2p3WXeAAn3RejiAplUirOj8J4F4dwV2mk
IIpn+wqOxvB9cpgTb2BvLMe40qdqD51QR9ADZwo1wNxo7lOrh4xhb10rAmrqEf6lIMGO1omVxgej
Iha0XrqNWzcehFXxw6WqJdx4zjvXho1s9Dfpik+0dVrTMe9+9GuqqOAXbjjMP7Tt0IyVtpRRO6Tw
inycVXaH8YpgvdsABUaw2+T0B4KiQG5Hl/WanlM9H2hLFS6xtG1/GyRouXbhzJ9eFpkGUDlTrWhV
UntnxYHguqQLiNy1OTsvzv424EiqTcKVs36PXSE5vwib7qjEYPrPCRnGbBTu7QhJ3+jNCRAGc4s3
rjpCqGqOfgrawgaYfzhAiGoYSgvO8TXaiszzOkdFVLxVPgL2+i/WgDoEZ5rj1u2UngclVVW8Z4yM
SWslDmDsqs2mKvN1981XAF1RTnu5EjiN3TpGfTFljkaVp8YFbYNyHAOQ+D9XhirJph/w9yHCRFpA
XuYrs2WfCjQQXSmdDvdWGqVyA5/R6/gvGdrAK/jEFFO4McqirGJQrZxCN+Xm1l+JszP8iV/VTsR+
JQI9o1o07Go9RW6KPGRILv4+dk8fvR57vvywsrd6sYjPhtTCLGikUH+bX7f1Zec/7/Rg1Hd3w9dc
hS4BZXeDJHSA2W5Qw3IpOpBYFDOIyXz5Fo/yIYmD/qewYKjjxW2LMmLMtB1c1+xpZpzVngtYUZBI
Yda/Z7C7FR7wWIadOt97qXVerCUqZEW/8wnRrjddnVMrr3snjBSe49dSVNKoFV4n8nbo1IpDWJan
+tEC7i67b6wSc9/lMTizgxsW3K4lqkfUDS7lmGRVLzd1z0atu/mR4ipbVhbT/gvZTIAwDnmR6m9V
/Gcj9ANy6BqX01mLJA2EW018o8JfeRCvO6Si4zfH/WihCe0J3fvkaWFEzb5TUAuPysPCIJ3pp5FM
9d4c/4JtTGdUj2LbaaAPVgFJ9Vv/m08vVtRwbpd0dH620SXygDEjicoNhEHnWs7dMkqljZNvMn9N
kZv/klh9HUkAIRTlBKBRA7UuRWDqK3UqdrhO2oQb3ytU70OP4I4O0Lw0e9Z0wNmwIjLwLJM2m5TY
lv2ssiQOuyYM56bWCnNWkW4UxDiVIoSicaJ34KkncQK6EkWDHLiwYJnqh15kVk1zpwsbeB5YRvXP
HkZgoAdvM8ih0Xo8D+X4V0c5g2L6NLs8aovugnnle9S/7De1CuA+kDumAdOvynmYF1hkmUc39T1b
a4reTA8n59IiFj66sxI17SnT/iPr8+bKw2I7ymKR7ar1txSkfBRlg6SIk+DNCEdbMCK0AX92qVjm
wexTzGrhrSUY6CmePVouDE5qQvguk2uMqXy1K4rKv0RarMOxAVMUEpB2W4GdeV6i/AMT9gjG6EEf
yuwh7E7oZOt0ry3xqT26BfCCRFda88MlDLNl3OU7CAKAVnNOahsJ1Y8tKfuXLgXC16qjx5Up1EZ0
xr5SMIozZFbdeLh7DOCSwadVLZB+9pcAvq309kYa9fIPR+sVQKueaIK0+rnSvpgLpPL7A/LI3S+5
LnKk0DD8Kuuz3lzYJA/XwV9w1xbgi53dGzhqaswUehYV0yu+oelfc2szxxa4RDsCKEriacnj9aul
gTjrz6B5E9ve03YQL1/tkEVhmiRICJBloQmASkyQfzKQPHVA7D6Xas3ydo1k8v1Dact3ROc1zuI1
J5AYDZ/OD3bYWCop67ipfIL6jW4yEUglIBkLGu/8DnMsGwSBLxwaOZcVdOU7xChXr5P+odL2Gd+j
B7Tj4tfm8rfShFlhwfCCCEpVILnTqS/tIjXenFUPvSw03eEXichGp5AG9RNfwEs+QXtc3Pue/5PE
azopRvOj5K1ls9tcDX7PrA24PPQwPT5GWY8+Yzx5AhplIAKjvG5FvE1OZ9/UI8FT1v3pfMkm3fkG
V6iT+UjtWg1re6fUsbx2L38GmCpWMhENYqW/6Zq/Ip5PIlFo5m7PUguJaUPy9/+XrcdJXMW/5QfN
XSSRnwtfHwu8CGKduaMK16iBUA+jv0yj/AmeDIVsD3VFv/+cdEmQecm/RanFAzN84l9eQATbnp8+
Qp/6GUHdO/KcU+a9bDlulX/X7kAtVkb5N8LGp3N7fULkiOqBKBvFL0oq5WV1XjBdVcD0jbQJyG7Z
jAv6zrHNtUn8w48CcVdRWXOw3i5iQEHbqkRUH7HulBu0+UVehk/FfNUkKY70itW3ucv2ud5VCMgp
7fBVerpvu3SsfLHHc4XC6s8f95C2yAWjFlte2GGKfaY67RYRMMTc9nYO1wNBAc62beoS5KBFISKU
iEaSPRvdY2FF5j0vdMYKP5r0RSGFgx+AlrSFzZuBGS6bAGXPeZi1UaC9NZdd+geCg74HUTYK+jpC
MEOzNEjifLE54ALCHfB2Ff5tSpm98F4KFOgqeM9ZhMNZv4suml/BQZ9A389wNNwcwj59WYPYEBb1
01OFJO3egIjKkSWXJ9JGVLZ3f+BF/6FMxllkOStwobOv6fPobwEXvhR2XX/3FAe6VzK5NGdG8fpX
0eWay9oa4Z6sDReSe4zubCZ2Vmw5F60Xo5X9vxy2lIUFpjRcr/mOnGqQ3ztZaK2t1rQSkxOs058o
0yMM0IUocghMd4kQJze1QDfQsAxg+N4mh0zluZDTRcAFl6t3s4JoT2Xg9flDz1+p5+AEUuTlr0ZN
trjA2+5YHbJiSdSgW3Zf05VTymE+ds47ulzsTBJxE3vTSG7bUPtxrC672uZs11SmkavnDj6TzFGg
j5uuGvtyRYUgw1XnQ9nyDJ83yJB4EE22uz+yASGBVCqxBwhSSc2LweW+ebMsTKE0cXnzB/YUPWOf
H36oty2ykOCnVRbwTcwlelLE31WtN6S6y0Gsr7tYzXVWc/29xz8vjl/Gbm2rcm+FCdRFtvsGJpYC
Ui+3dBfkooFJ7sPyHiinC2jgdamRL8P9naMG+ySwOuZFO5ga+MDYPlRWEcp9ny93PTQ7zwheYzus
Er6tGgPX+LmNsnZq8FaxIC3cECZS4/AxeLMkgl6kt+cSIZ/sTZkzKIs38OFp8l80+jpaROzSTH7K
6F/ewhWm9MvN05lQ3IbVXK72ZQKvI9ll4hVKBabxmob4xYkBj49wTYbyAoftkINO6nNFzWp04HfJ
a8/jZx1DbrTCWyWaGgtxakXLTgDLVMVYhAT6dLWLPxX+H/gZGHPhXy9eD7xXIL9pBsi7WejnaJfk
q8PIAsaSlZZB0OXLEh9VqYcTJ3CrjBxMPno06ufASlxFGwJohl7y9kfJaJaNp8lN0VVgREHgoOcT
CJmPc8JRWLr0uAFe2gFfxL18jWw0R1QY49fSqeoI8A0rx7ZG5Yn4d+7lLWyP/LcrtZZG+m5WJWT7
6UpuAB4FRwDBNNm9961HUbZprHpSXOxhQEz+Vcd0lgTkhkzzjJvuYFSxAYkjMQHPFBWd7Qr5e/wT
GfQAU3kSgXt0QoUcca4MqyLFOheQxlFyywPMlPROkFaHyL98qnkAuecN6jYep8EfmY8Z0jF1xUip
ctNeGCZt0Li9bGMp4ug0NnviLnqRaC3V0+4OTtrofX3RwvvTS3kOSZjDkn6SQiVtqx3yIJ84GL37
VDRKT0lWaRvuS+TMlV+lqByyCJuVY2tgdOBHWTBB4tYDtTgQtnFEsqIYbMUR2GRcZ+aI0Mn3ajhE
H8NirlRqKZO3drbFNsUeBuM8gHsdZaUio1G8BJda6x1qrPy/23Hy0hzJX0tDRrNZupo8YWOJONQP
Ho+PvwaujB81DyOGh2h1xI3TEc+7vcz9jspFRg34sTlg/3Ln+RALwwLUyfhfFDNHLahsytFDBoks
ONKZW0CMfuOeovGVFKw1VF5VcXSghwIwxGiFGAD4Jq0STb9XOic+8yT7bS8pUlyw8DhzmBIr9HFO
A0C5dj2mZSNp0iTNgeTO+g2+6173Bq/7PzEirykfwaX7wedQNENyuWEWbDL/7Ng+HmRWp6a+NgxW
eMO+CM+LrfCxLLK1pfoLpaa+nSWtN1kBA3nf0WBgBxNsAbtQUtri3rNHaMqwmxDAQJDssyDs9PqY
kv6HPcZGL0DVkUSDjxKKkpbjvYDjTGs9tb3Ur7d4fSpFCeqsfGR+KNwYMsSVxZ4ilAvTNyZVWd9f
eDKFiBS/lXzPR/3Sn0QdFKuT8wTbQ9GtKToHzPlQ2e0uR/Y9E6lj+zZvvVw7qyXRbJi6/Ww3QbS1
q9aynUygHGbI8HFtxv0duVr6cZndtUR1WTRawNTf2TqG1lD4DYZ28MtXO5qOAdbCc9WnQ2QwFrwS
R51I9eCx+FjpFQARLNh1XnlipzUYzDf/K/3vCdLovNmg1g2jRe6haCO86DoenpILPTPdRyNC0TfL
PkMXxk1Dtaz1BN0K2sfGNR5FL2OViLhMdOJCpGhwkXxiHqXLP7evDsq/bgL9eTWrRNOaB9+ShYwu
0R7rFyiaB4odNX3mNlYAagYGC8BlC8lusiU7jquBHe01Va5wJ0TDxkeQP3lPZCLGPAsrA0tIVviS
TlZSdEag2XmRtOUArzi+XwvwDPNUSPOoNcmorbhlIIj04JiVu8EqkrQACwkJtpVGWhVo7OubcZpg
S5rHC7ZjgV57PXVzKEaZSgSoq6iv8yXdegQbmAoUCHHfOex2dsOR8JU4i/84Y5g0lcqBBVbZNY6S
Ue3x9XYaC7NWwTMYNKBRg7nrynp0TfYTwf69JvuxMQLotN4emYFQNpvNbJ3RcAmwzZV+xyXn7f+b
ojKmf0/1yoHYc3XXd9h8X1kRKd2RV9Ta6cdwEDweXWHbei68SHyyJ7zapQAAtQ9e6vljyAuAUluH
QvXkQDbgAF/PSBf3k1RgxlWJ4Z2YC3iy+FMkgqrj1JTeoT2Nv8hHA6XKwP0ePf290FNl59pA++3K
POasn6XMzrawCxfzkVu725RrreEAvTKXsu4b4tlIcgaS2JmNS74RyXtmtp5ZxCJuBPSaYYMgxq6r
chNgw4PNPVyM6OIuLNhI8vGNHY4QtjrWazHVIPW2hqX67dM3gX62eBFoCvVN74tJSgTAaLEWhwzg
TfJiLM6X64c1ka53SCSTJwemlnIgFXRCAwpRsUaGspUxnyP7oNXCishVIFKvo2Zd9+LYj25kMz+h
+TppdYYrWSxEwFkthrD8tg+YIsIrdPnkQD9HaGPS3pHFwSxOxWGn4Pgkxx6pK04JhVKL4uTbDvf4
L4AVzBI6MVfb66M+wgpXokmpYA+0nnDNixbjiYkml3MLJ0aIdKAwnDPLAAMwc5bf/FpDjBw2TPxS
PLGyhI2ZgsPReGKaP4eHF8ExQI9EBXULZ72fpeZKLuiTT39w3D7V5+2L2+ulFsROZld/eFDdLdDc
ZmyX4Snm89pzH6MrbBjaO7YRzkjLkOZwo/3c/EpaTL7RXpbBpxcnSyv0MWmOLb4tdOmzIzQRxNQC
izwa5XooiG9ktpuNV9ZAR/XiVZ7EV+FLYSQdFfpsjhb5YibudDZPDh+96QTAgdCLWX9jWFOWPv1e
yVcHD/Zm+9LJsVmZi+w9XXAnRbAiTGjYupaVtypuhAWC1/uoEk4MC9b2bQH9RB792drOwmxv6t1t
dUpQc+hoTjVHW+a2jMFLPm1PHQi7g+cfAr2hx4w/DSpzXV3Kio1Wl61uNcNzSYkp+Pvx3aAsPhX+
ECm4Mw93taHZXgv7IouxJdw6irtEkCLTw7fLOJxrqtseUMM++wstVOTg5UpoAFmWNemEnQ/Du0wD
uk0UaA06eyruShzhDx1BMNU8XvJlIIezhE/gDYoFfdgU2puvQkvO5Jl7R5By8gU+YHenIeV0J4ve
TZnUYixisVO/JdQQuNe3oANW/L76cKO6BM5j64zxb7kd9tpakJK3gsOKqihNQifE/+1xvqn4Gldn
JKlg5km5+OWBVkn08Ci6FjHi7UnGMwLYsCgKtHRvquLW7fRr9Jeow+e+fMurJmuGFGKCMzvoeGwR
aYyeKqs3uuBsgwiWdG64m5nY8rFQc11sQQ8t0rA9I3idyNU6VztyvgIr8Ye00aSTRNcVN960oCTk
YHj8DEUfcORAYK/ZOeBPIqOgqx+jCE+d5gRHAl8oYtND9oKk+FFhrBl6+ERlFtNQNUDlygb7gcQl
3I2+bbQU146aR4qK+EAoCVwQFHS/hKqELZQqmQkVinb/m1taai4+jfOUN3LaMhw50525fsOF5chl
V15RVMIwZBLaOtMfh/xY1/p7g5rXqZSJHbe0Y3A2FyX9LtIE6gxfK+AqVPDte6j0yMKNwZUuHjsF
anNyhyb/yo7/F3pjIyDgboIF7IKpRqk1MEvgt3/No1sFe/O5UIhghRBYUUQWHELWwnAGfIBUs8ur
yL+yMhsbwwwcOOGboSJyYzjk6+XatWTTkpoNBlK/JCEAzjPjUkLsXxBWy6DDPY4DWb+XFdh80jlC
s6Ch6OnSDiuTuUChgWXzceqnOUtWDdxZ0iCYbJcTRhHmzdLG2RCffEASI3leekuX/UsPXNIXrXHw
0OclgFQ419Ba/Yg1NHriSqnJ1DdKStN6V9v83qd9NzPCdmZ4dfxpoD223bFDQGGJE+jJc3EF4qw3
ZvcnoC/PwM3NCbBdVUCoFdVlEh3G2C+539SwR3e/t86xIRVnZg4E3QF9bRhkIvahS8t7m2kaJVMS
ayxZBaiZtqIiUIiOT5BolEujMvWdcTqi1/FZrJRDgkwT6fS2oOzjncR8jZdFIArfnLniGhRFcFKl
BMMFeuRV+c6Mql9vY2xQlIcNqUvrmTp77PFrKbS8zNG4R51bNt7SxIN8QaGFKLMPrHfu2gW+V9c5
vcFRKjII2gTvLYZf64xPmdDze91SDHD5bPuhcGMGBwpr8xu4chPkkfA1KyYITOLkBD/kGLd/xC2P
tFnnj75PNi6V6e+ntCQmFMTxTP94AziNdWSeeisesNLn4LcWuQDCIamKcPwiqB1+4HmTUv2YDxZF
IaQ8+olOQ5dvsL0yBMLgmIp99Iw1+RpthnUj1KP6eKXcSa1XOlpt/WJwaUL1WWcMP0M8W3Mg4LcV
fkrR1IJdnqQg6rqGidJh5mz3p0izti60K/5m3y4cVKwdWzq1C9BNVUFSJdqYDH2FWAdS1URc1Rws
INJ+t1l5p8A575cmskp+wp4tHBi+Sn74VhdmbDZjRwLzMNoVbc0KaqjdI8f8on5cInk8WDr0Fg+N
c0TuJTUbbL5sla8S3dIsT16Zm1uem16BH3fn94kmF6JYLuun8ZSAuQskvTFgr7SR5OMC5kOkCLIk
6Ae2diQbeDoLZhfQOzasLK8ftX78111WL42NkLnbWBYj67WblSD/2oOwxStnVTdyYdEZ1OMo7+ye
8AEyMZBOkshPoMpdoG9VnwDi/54qkNzP31p5LE4t9sGUB2njc2EnQpy27HLxCSUKWj1czDIZGCt5
NfI5tvyuYj5c9yl1/cUrrMTNylxomVtjB0Rkp3fEFGEdYu/0Gz0nkKyO8H+o0mn0s7WWxLdh4Ha1
no/AgijNF968LmAbizV04a+bP5Bfqugd1++PXxSYqezsKosHIroZqN8qRbSKdZKLFXwDe3mdY1Qq
96OToOAtly6DBCgLZP+u5c+hz3FpkVFsP8/0LEf/7KzSpO2Iv1nruBYKs4b8BsEI/Sdvv9dhtUwd
+z2TEYQAfa0lI4JAXUBnOnyKfIVk8rEt4X/8CjK+W5C+lc7RamwMCOACz9bEP/g2T0bDvYgaybkR
gFu+pUMQtAG3MIm7m/JVHOOTVHDRDyrPnv/DcIev11POdx/Cw7ECNh+1asMF0GHWtjGFVPNCIjvk
FaCs+0gxd2qwdRLd+cbNFUYew2n6leA+HuhZaxaJ8QVYa9dtrd4+3K/UjpQ/YidZUJVHEX+SxIOx
ye3yU0SGP/UEOPYMXHWPBRlvO2ubhwupltQVBsaSjj+0vFHfz+pwaOg9pREwo2O+PDe9ZyqiD9DA
6dIjO0il63ndOx8oGkCtgkl8Oxhmx4K83rLvdZM3BwC4ryFZnAomf2JpTC+sAKxlbQivKUg+xw46
9uB77LpkdZ6PzG7eNX0O4THlRtzpbSV2L9WDU9o37uuTkWJVhj1fmGX4XMuVi1/MJoLvLx/wjF5V
H0bfVZciJsUVO6gogN/sqhF67izpovNL0IDueVeHcsTAF92FbyJefcLlnJKgnIeoK+VvWmD/P4Xm
Vyf8LvDz7ld8l1UOyk+aX65y4u5W50WVcE3jtjhfRPnr9RESYp+BxPA/nk1C+kwwoDK+feggLw8V
leMtveFOPLz0SOd3ybFtQc7+zbIIOr9UT8KJYVnyyk48i8pCFrycoPSfzrPIKCKjM5UxUqK+mKbv
JhTvPgFcjBV5vo4ignk5FxPHNMpH/QHtVfFLhSdcPmY7i1SHqp8/PGPSYScEJeLlvgohLwaJ6kVr
EnTUj0q0KxjbXFjnTq1Wb9ekTyrqQrZP/nbnFudD5wHctGzr7ehUZ2jXH7MwykTYHpxSItg3XjcE
Lceab4cBnT0T4aZFYPuFXpIcnL/BufwtQX2A3kLPyA/sYoaf/QViqJRUBUm2YLY1xtfkahz3CLRM
HT8x7JdW8AAgmz5DqCBtWmvI8Hsk9ZlPKXb9zuGLfn8yxEp/Qp6b4ploRkOjYMYHxUvyKsKRfiNO
1etTBbkCbLRFX/5vRkEud1yyinKbBZQ42tAaz4AmOXjb+g9zGeoKd7zUOlgPp8ro3v7P+DqMTISi
8K9Q6RRYTnyaxHuppf5lVZp2aST51TyicxDKGfGdEeaa4Xv4ZCmYqEPVczxYwVsPC8D2KlHDYEQm
SeUG2wgiuP/OI2m7O4F2Qc31B/RlGmRVUujoqxLPLi++8K1jiAf6CicP3WmfQCGGRWkXtbFP8POD
2UILS7jhDZNVV3wA63vlkMIAYtbd7zT9Fhyk8E92TRbTRlry2fDFmbQE3fZ+7jRaxOEbn5Mpep4u
xw50FWLyrSw8t6wdKdgA9K3MHnZczFiuYaSf1XlJhrtuu6buJJ9VXktE6/6AWAc35kDHJ+8KrGKE
b4cq1kU8GXRR0rtb7gjSpHBex6UhwysO4i9B6iT4WmiaF/fjr8QR/OW6q4QyqqK15FO/pG0j9lPa
shOWz/Q4y0wgGkc6izQQYKKoy+LCW3bQW6b0HWVsH546WFxJCAABIF9a8oo4WNS3w/YgTVcnWNCc
yiyU3A+atMgWmFhBX8SkrKVvsQ9Gs0ow9CuFoP0WMOkIzpScsSpnNRqK2tFLplDezExmIqImQKh6
+ABToi5QnnQbk7enibhRj7Z+wUcjWK5y0cjhBoFzRtWPaBQWiBL6Q2lwfCK4k7SUk3qMzVMEtQmW
hzlcvDszqKb1FULWTqwAMtijNS1p+r/3VgQNCw/7YVJHcbNDGJ/K03uBILBuf/HSLDlZM2js5NQI
vwAaKr1DCAldP/9gMi7iJQDDCdJuwVIRdA8qOQJCfCBoF9woOW03B0PP6mNBNcG47c2y/xefbh6x
cRwXmQujed4swvWrXjjb2sbZN8C4Sfa1HxereM7x3Je2qiP6qHPdx9OdzdrN0whEqwK4Pg5308XA
BF+obsjtYfABq8KPGPikHeMSoE81Lyzr+ZodiG1Iy7bdTFWC4rD/m0RjBWhqMGMxBnA60aeDLGZA
LszBy6U3kKdyW2T7SR+ykqfFr458Op0WcUmsrB+apyy7FvS5OiH7JTHUKkZVkyafFVJTYbwNKYpF
DXt0SWjUiQ2m9pLlDmp8jvHkR9vI48unPqgju5q/6BC0hXbU7ZoDIXc/wU6KLEV7Ey7ZdQ1bIdiK
gWIDjPZNkU4rkQGRs2GP9E0fBz0Ohc474NZel5SCgEJaYLV+Vg7tdzOmzfJw5yXGqpFUH5G5Tufd
X3nlydLSLvBc7mBKSrK06YpbT65fqKVKomp3+k8gZn+5OHg57bwnyRd9q4UQvdltdVEdbds3WpsD
0fFf1I3SZ0WpG/Q+AlfwM6qYyVNulsdwM6cgX31QtbcwNSqDFtvLEKbOujngQ2h/A6w9LyfKxZ9M
H/Izpoeq6zGC3T+8UI74Pa2V1mT55aWEfNJE+nBi6thL36tJMWG7ZKGxstO30LvYtsugRJzmjiEt
pGUcP9SwfSqF4lNof022/Rpbl9lMvUNcwunUVXznPVPekB2xiXTvglevoi7qU9q1SML/tVG/uGxB
V1gXIKf78ulgcjmycy1s+tZWSOcRFTHMobc+Yqv0DYUBgMrV4uW/KTTogTK25q38UWemqQGo+qk7
amPKOIdrMHHUPB1lIs6LOzmbGorRKuiXkfbQmWkWpU64NRj3GRQ5FsNfFgmPXBrVDQwaRZHByHzG
pdpt1ucc00A1Eg1QVLdaqz3KkEkYtt/akSwWiJbkT1NDUVsCX5d4McTLWc1bWE1YFt7xxMMRO9BP
Vr6BXxdgh6NugIqfNSt3BDeLuYnuyh6Fk4fR0Rg2Ev0qBeEUWIN5O7VRGzso88V/0YT6XOTbErHI
e5AFt5Rj4a6UTI2t+f3Jpa/QYVljEPYuGaZ3QfE8i47n9Bffz72p172kkuL7mT7ZMzYybrpAGmjR
2oVX5D8OsMMnRjKIaBs3x6yHZIRxPti54k4LkBD/K2//sDNkuQhfx+A6bW0icUjcWAnnR9Md3WYf
DxZQd9gQFBElIRKygoT+jDJIr+fGkMqowtMuibgqOiobYO+QeS/YjdPZjNjnEl0p8PZdCmKV8QFR
7WVx0uMonsgUBVqDdlRlwOKqE/NpeI5uo7qL3f0B7Cf8/3eqmIfkiJq1dyBWQTSM6mGTk8y765Qm
5I7+BYMzNvJwjMAD1aR6f1P2BUSvTtPs6qQ4HdKYtUSkzwQU9fN+b8wvwy32HlkYx6vb5MaAoyKW
J5pk7rrMR0hoh+3Xs0K4qIV5aH6BVjWBgk2KrCZQ1cz0Nq326iqs04xqCwgkazuQkZKtZjrqKNuR
c3Hn1IollJNtNVktNSSB/ietvewrpatAwr4E15xjEuEshS/ToW+v29kZm56uvYOfsBvUJIYsUIdL
eTk3VxgCkd9aLqOMJz97PSajVtsMaruATktZ0lEAFVULCw1NMVMiIZI6KrAXn7wHSCcYyECD0Hq6
9JdYRDKuAkpPELvRyucz+oPxPGc/yDvNOPULH0U4+lQMNSqvynT0m59oIgq9xIqxQFiIphhUjfTc
LQscf8C/KYhCQot+wyeXpcWrWc6OyNncSXyQtFncMHF2GrlNuXhpdurv5JxyfVdFBdOgU6Rz1l1R
mcpp829YbbC23KtT0Stluoi2q8BpsVPTLXNdh0iMQCeyw8u2CiOxRnsW0TnFIhjCwnoitewxpDGT
kr5CSngbT0cT2lkrzSPD8afyKw+/IiPAZRUhzbH6pDpAsUxXpL/KvuCYuoTQoXgt5uPqC7friLaY
cHVQjP2WvojWgbKD12JJ6nNI1mas1VqVwzm+zV4YKg0pi/ZrzBhXt7Z+Vw0Cn7suawZjzoAxOncN
DLtJkeejXDJ/EiiG3dkQUSa2ZyWEaO9P9MxkOEYEVuMIG8Vy1bjS/fwLa1FxS1t30HyHpA6LvSVD
vHKJcJXw1He93T0RfgyoQGyVcEJRGq1K27Ifd/DrQj6PlCr7EdvvRCL6otlPlyIoIR4baBL4nLtc
7Ow0spMyLxdKfPTOIjeUyqFnrqXnnoXP/5Asg+lPlHsjeCUVc2uuhavaMd0qjFZIBnHvZc5GhuLq
c6oSDNsMe4qdAOrHtc5enJMF75j7rRNdnQt/byRBNLu2Baja+yMebOOXy+hIpaQAiqRp8DJhJ9nE
bQSHlzeZoWJCuJjol7B1b7Vs6wbJtU1+9lMx6a6cDcESsxJGyJTxxqRuB3jmHshv7z5m9iKIqOZK
qQ70qG/K8K1VM9HdHlCQkj9gA6i1bQQE3lbFVOQ1AZA4FoPznVrjB/zvYDfUUDZjtvGxtpAL73iy
Z3ARN/VHQuCqJSf/9ch0p5H+gGY9gVIR+Uskrg64DhIXP9diOTg8Zw8vK7YXI1kj9EZ521xIiPLf
HmJ2sS+RJBiE0Tok0Q5QWM0TXbFISiouAd9TaYUjHzRwy0AW4Z+C6RSZxet6W6gaDLhv5Z02TjbD
PbdueL/LSbGtaXFCrB9I6dm2WuypJ83HecsQhnVTsZF8wug8g2NHXcdWtVtZLQiN/iYtuageGgD1
YgQXEmDKUzF+G3K6jpEyOGTjeDThD1dj4E6K08iYD9TzKUEaSu+fieaw8MGH9VaDakO7fqmKZkts
FbZJRyWVGZc/A/xhqMRAe8CYQup2aN9cCDcc5AO1rXHf2FYfeKzLMVf/OumW5UDp5BeGJoRnWPlx
zKx3KlHiO1KbMH6Cad6psuw14yA87NghT9apSheDKy0t21q3QO/azrL16SPsIxshU5WqadR2b4KQ
Ya/Is/odQUtxJuI15tUnsA9nKN4XUcEcA5iEbKuEAFFUbIv2S6BbjGQg2It1hcdev3ZW4y9Q6iaD
i0dpADkVkaGMqFx2KcXFpsFu/4I1kOsceoZcD2mALweVj1SSCfp+B2V1Jjs4TjJdU3O9WYiRk82G
OTRhBc81FtDXWqBMyw/oIz0SUaMZvjyRhApqTVRg4394Tzza2q5e81prbjC8RrchN1X7cmjgGN2k
1gDSVj4QGvyIq/BpUf2x3jl/hfY8pOuiE9rgc8vfVmHzsmYYjosdhYRLyfLbjRWMNsYht1A+IObQ
lw9YzTJYqZ2ndql8/fqCwZMY2RysctmmsoiNUkvOJmTW2cytBWuxasXPAnQQk7/9PAQZGcSrtPMM
BK7rGBmVa4LDufsn0aC8XCew/+v9mqRGKt0kbP/ANuVzR9zofSDbaf4TWMtQV9XCDT27Jvea8Url
AtRfoiAauw8fZJ1+UsZwlPseSSUq4Xlb0iPjhephe+CzKteLCKY6gQg1cd5lK5ssl8bvaugig4F9
6UC4BtSUgxnJM7KBbbcZP7uJ5YteXVjEJAAnbCMGzjB6XxsPGMfbnCQ5R8fDHNljDWPOOApQ5Bb5
kqXiVNMYYrgjwPSUrwSPSRHWvWd1WcknleI2s1TegxhUIJpZbWvfg+IabAUfYnPOAKh2EBsIUP7B
Q+6zMfabr4V6gXaukgPRSdXkeGKqCbTYxOfGyv1lwVlYL1TxZxSsVeb7eR4XT0MEIfcyfD6uqh+j
sBLuoDNUuap/l70BxqocsLhtGriyzKBmZDfP5R61D5D8liQEvZunt7GWBMiO75ZzV3sWPMX1tEgb
WAX8RJ/rZtWsXtiKxpQC/NFdaNjy9Mg6PVA8cZ+m+SDPaC3qTWW/nJ6zJBDxKx+hcBHSl1R0p24H
5iVBSceGZM2Nm+eX/YP+YhiTJchQyAyu4y/R3rrCEvYwLzfsHN/EgZ5wnfnLs5CXPprjTw6gIR1O
EVbSIqt0+0apbu1IXXVNuQiMtR510kOqt+5v8Uy2HmEfQQWuBARIHkuOQ+tXXAk9uPtx4+oEdC1R
Q2dXUtUqeOLLQW3rASAWoLDiXBZhA889yo0aYAArRQnbe7zsgzzbxGmDCuo7gBOmgUIoqKHXbjwQ
jXEp+grKbJ/MFexFoKxPy1Bvasnnz4LlVcwO1ifDkidtES5KaGumSiIrp6NV61Ibbt6iBxF/v3ge
wSrtStqxMR7y2NSpybhNjV3uM0dkI6A9P6EXxRnqFkkBDisreb8zKxC2ZRau/vV/C7Tlg/zhJisS
DnXkYsMkqbkfpx2mL/+6Va370c49yxOctY21BAiAS+g4YLw5YR00TS6ajr6zLrMqH4hxajYNK3PT
AfpNPV5GN4MFpkWk4AmXiPUFfNBVO8xv5mymUQVESv+DD0+GTPR0ouSdWB2dx+oQiVuS0WA1nDRv
6ZRC6J3gkgFgFvKroFQyaisSEnJ8hweLecCZrwjrnp9s6Qh1qS7A8uX1/yCw+cDylFHwlf1t43D4
DElVbAUp61fMLWE4Frfx8YdRHIBKTxXfcmGLW5a4Jie4T0fGJNNfjdUJiAZwKB7L6idz1gzoFV6o
O4u7NQosDaXqbp0OhIrAfs/aKnwTqoNTjqNc9QxqdxRgDMnauHvT7WLARnbd98VAu7miuajeUfxi
ioqHiIZJQinYPUL7busGarPNTR8dhEWdC2i2MmOWyyFb/CVYt0TF4y+T/RLqJPXYWB/yWu///ukb
4qCdHRk7fGE7LalE87IuB2il7Hz/GErFoGy28k1woSH1FuHlk5KC86DGV78JkQQWZ/P23SHSXchS
NT1D5opYq2GNaZwkNTbFKcJl/iE1pKrIbZF9SWtheKHqHvPnqnqfUrcY49V0OGLHKeM547i+Cvma
g4ckKUC4LObyh1xKo6c0d5gSMrfx12AraPWhQ9gysNrwC3+wz2/R6crIvmOhvFegq6xNT6t6K9K3
DcFPxrqYyuMdZeWq3GMskuw9B0qosLK+UgFBI+JMiBPymwIjTgrEciuI2A8quuYlbXBnq2RKyHza
k7XjdaMSKR7cIiLxsvXZ4sxIuQ8xuNZHnUH+90x6D+RkJE6nHhZGRYsAEwrptCc0CAxIKgwVvzeT
Pbw2ye/833k+qHIhirQKpF1gt0th/SYdIDv0rWkcAT2mbFlEnlKnuscqK/53pA/lRGgoTe/EEjkq
FhA64YehbhIP3IC0vl8DoBuuGgNevRf/RWLXM66jQjZRsNMou9VAAxtWj3RVGkOELbu1KliWXdMW
Es1kVZ7aVnWp4C9BMuKs2PMqS0sYtWrV3JbIPlewZSsvvxP8pnqkHQ7NL2MpBXfKljPQhYeWrdby
/DllQabe4o+YC4VKXezywTq3ArNzZdsUt7b7cqivlqjnJkHwCL9O45OogTbvalmFXtwpvcyGjWPP
bHgqfbNpn1yvBwsDKcfeX0Sl01CX7YzJHYSJ4CSne0PXvSJrs1S5SnAMuYbvhnL/7SRWM2xDm/TK
sedvLnN409gY/4TF06g2gpedX9PUz7OlWNyrAs3EypvGRP68VPdTOL0+b/MbtzUg1bCYrvNDtO0z
6DHJJDDnIz5fBZtSbxdWb2QA/rSG0WBCbYmlBluKujzAu/A0bYVJ+iZuAmI9N30XoJSIEPWOOb4C
SCjzIYbjvg021+u1IP9A2fC+73xrmHFnDNQqga/SdubaOStYOggV1HcMcP9EuyJ9hyh32/wyXQ7Z
k9ArXVRmvF/K8Idv4UZKPAELGL3L+wTdOejvKQbSkJVYjMXjIDRyAKPTJT3iA7vqooE+Wc9p3Ug0
0FcVafR5GmW8yaJ3yerJIWAmYKh9rCH/xJTupGW2lHHYCZ2PI43Ne6cvgoMq4l+ERB+2GcSqVUgp
iOWbP05GXUKnNwDzDjxdYGiVDliqyorKKTmMpDKW85ZiU8hAJsnwIqHd3mXFLrWl6EZYq9lpqaXQ
C4/YkMgCfkAawLpN6r1sZ/HbwjXuTxp7L940StzZ2xISNULA9UUgIsZXFhJQskvFzZGjceoAsP25
D6fPxcfP88Rm2N195KGw4C62m5QHFXIkyiHwdZ3EE6oQSkTSzTVfNHRX5RSIC5Rmf6/sCjcOUBWJ
+B1Qjx81cTQv9qyr5ijQghdRlRJlSpGcEpkkmGswplWrjcWAZ5/VRpa8AwGJ12FYD3ia+vyzu3LG
FkPNb4uFEFng6nhkP5Ae5oaSdyxkEuQ9POSbuitUNGhcn2makgcp1jH7Y0qaA8+PIFEBCA3T70FU
XVdWCkHE5qG4c4sZ8kpetGsYp+Yr1lJjoUiYQ0zDCt+usJwHm8H6DK3B98AUhyg9xME3gicMvS8A
iANpJZsixiUE1S3mdXoICXfa5DL2s0fHL2gTCK7VJZ3oWS+MP1HNhBNdJ0eE5jf5cOW8T9vQszC6
POSKDuywQHKAHcg+pd7NbLtzHuBbRavRoFKgB4pm2AtgNIOTy4ApfCgmOrlLamTmzHeKUufeBEth
H+0PJjD/Je17r7jrZid20IMeQ8FUDuzfYLoGn3lks2CGpNPT9zbAh9EwSYJp97TTG5M270fZWRt0
pShgdnN7Tag9a9EXp8OABbRXq409pHW4WZVn5f4f/yjPT2s4Q33tw+lmhy7foIDIpM48eBavcVPg
bvk3TacUOIYkBhLaY8ye3o9qXhcvqIk0RXCD4A6/mWuQV9L4Xey8S9LeCIJ4v97tMjM74pB1xbVk
iQKyVEj1a7geHf8DRNxvfXWIq9hTh8FVHBmWJYL8IgdyDvSoZGp9phGhE8aeJUmLN1iOd/M+mAaN
QynTXOaurxUF3Opy45DY6KvAZDvVw8WZ6q9ISSlbMQSu3HaEItPh1MvaPbvakRQYytTF2HGTmfpx
0V3SAf2sOP2rEnw3G5BP/vUrG8CxfJYsXQEiap5sqNcKprx8GAYAMeirYK2EoFEyyDQzNDZ/tC1p
pyqItn1jwIA/yXS+fkcXxR36RQXXSo2AiZwio2xJNqDn6zIxnFPBnq2uyiNXdnZFJl2Enc8RmiNZ
nHCSWUb7MlnqfcBY129pCRvr1EDwNZXi9k0LF+cyxj11KaS5RUVCjFiQOi/M4GQvjy2zOiI94wpF
uv4wBNdREP0EM0mxW8w9l6HmmciPwBzb1TbiR7e2jg7oK1YLoVlkyze34rszfUmDSznO6x2EuNed
tWOzbflTnXqCAiOn05nQV+zzve0BIb72aPw16JIUgNCKUJDkRKyY8vBPnTZUnXDj+k4da00dzjqW
IlHnZBvcDAtcelbhRGZKiXPk+vF1uEcW+cZGvrdnhS1PTWrMyrIDTTiwS8Pvo8zOs7U1NKFoZ5Pf
veqVD9NNBghb9x44T7fMmp7zQripfnoPnF2IozUj2kVW8ShMIfx0/7Gu2wkFGY9Er54YKumaJAAP
d52suVKloPohPLHXi5yDI5tSFEpIRoRzVyatM0KTD2zepvNsqHjDwDqIs5oz0IFzKJaOTQpAE8lo
cAeTevX8bzWKlHl4qTBA+fuPlNlNO7iO35SnAZLRMQJQvnWp1B/FLsS1QwTQHlWFGvw1fLQJFrJ7
V8Y9dx704RHe6itK6vIKscczPDbW7goCiEkWhvFe5m7U+jut+eEPl+KeZY1ntOa9RD+BLzsonbKv
mCvkzp5SYi6uykJ4NyoNB79hnt5GXlJq3i7Preq+rtnHHt86rnvo7g/RtIrFTuX1LMSYDd60g559
P0eK1tdUV17jg1eyQ7p3d5kv/R2tysD+0Mk7pXYq1AZeWTFTGomofkCfY8wLFZPHdQ70ydhTXkip
++ZOpvuyoZn5WrT0HInYmOYpDq1Ok840W2d+mxjiAsCkPMGq5Lkwb3Lss+1xtvhtxefTPW+vWtCZ
sJunjaAU3/HCbYBLBicKG9wKIu0LhQiNyXbD1E40LrxD33VGIMmmx3mo0Hzyy1c6Avd1nm56rk0f
aKAyXFwkTBlsu4K6IE0p3W3PPycjFaltqILHBrIVIN1K87mobR0RaE0vh/52/xODWWH8M7Cg59F9
W0KgYoYGW6EDJas3ih9aann28QP5Ph+M6EO01/UWcxQRjRP5bLKjNgPdNTtztlrqfRDUh+1TZMuK
w09kZK7Bt0rSFvTGsp8bjcjaFMPC5wwxZYSzWCVgqZRD9fKOxzfni0k2tQ3lfv6fIXBSEEGFz/Eq
jCqa2rRmIm9eo6NO4+DNq4ELJMV4LpwBB5iLbfo8H4UV6kkdj+a8GeqjAy2+O70x8dy5Qr6UO3V7
+Y5226zrI/xAvRHfc9hanEYun2U8VXGCcvpk3A6GqLHYIJbn8l12sye8DEqFK2Mst9XRKd8Ddcgi
86TEWAFH/f7zSSVHzdZOG0n4cpAnc7D1d7NAurhkbsDX53lcCUc9YUEiAIqWh1wTm+5lUheSNIjS
pe5SPtOiKtN7d/OBGtLMUA+xCv4OGuXVtQcW5jtpjLQfEixqla1/3+5OtYtByxf0bT9l0Q9jCZgi
1aoGagzXNBwz1ilELzNjq2uYGCvM2bnaCUM2dqo3GRJHu6dMWB0PlTskKKbdAgHfuDWEomovYN/S
Dn2C/JmTJXrqa1kfngZX5BtPkxP+2+zvJTvG0H7wNk+nGBzTeJIEPEudCSOEQSBNvXz+jv1H/eXd
3cIky2/nWyWcdB4iErvrqt8+iWLXPwbsk7a1jtUnO64QQoUiZ582G2PZCqjz+i+4Jt+L2gPdOtZP
b1mY0LO+pPTbYX/FMU/X1h0lCKik7nCEcM7QSvv/NENy8WJtbh6rTIOCb3hDiis9SBfyToTKr6I5
pY3MpEgS+VghcVDpcJ7wCY3rMxOr+4zOn0GJq1wuDl4M5hlETb/2pQ2vsjEWlvg5hH8dZ0KNF5Ea
LdEcTS8pOOxcXxo6iIC7vdLN3ALN8cIluGna6zNcl6pbTOl1Vx2oojHUgX1NZdCcSQrpDbWj79r+
bMEvEH4cMgtQzuJ1MkYOZJGRdQRvEQfmFFPA+YMCeGv6rqOOXHZGJXq8pM/itmyJxkAHZjDbTTPf
+pJpiXPl0PcMTk6VNWxx42o/2duX+oaZGBp5jEN3SCaeC+wf0U+TETJCLDHfHVYMT4D/52ofS0cO
0a2wv7fsY+sbJV9wlTPm9LVXbmq9EcPJtHStLn/0Wxnoabfdrh/YXgReOysMSHU0G/e+dpSCD3iJ
qGkwztWCwvYAXDoANXJXjIYXE1Qo3hrlA/PIIeFl7LoEaAMqJGTYs5H7QLNhoi6ZO41hHpC76vSm
IHJyHliPiSx7Z/K0lNrp2x8augajat2WKPrzoGkSuBWYmAa1O9kXaEkD737VB9s0wlDzaiQjRFpL
fV/ei+3DidMEVwFXSPe6xtLDa9J0SA4Uk5kNkdZLC1uN2DsAnTu4RTPt94pLx9NWgP3SrK+d/UUw
2XirvZ4w7mUhueZeWhtU83Mt8sKsi7zxUXDx5J/8w8eJoq8e8ohjfGlW1CJosMZfcCWnilHFr+47
+EyEWT4871GIcZ2bPJAhpWeQyh6CNtlhU+fdBZjvSNQ6XX7dmmTX98P9p0/qVdoTPOjptE4jMLwW
Iy5aFXt6gysm9Hrec505KinWFlc2UDF1xyYB8o5Chxi4As1uQfUWi6/36MxxnRMYRrFQ0gSN8cXz
kGY5e0CHG8LiOHDDJZZHm6KXX+gHUIkXTAMK7ItzKsoLNE/IbbCAzRrZh0Lo5pWa2ZOVyVzNsp86
RQFyweSELy7RhMPR4pVn1VRtFVQ+p1EEx2lAPF5KJ541izYwHsVJVz8gyUqH/hpTMUz8wVQIommv
N/Lw/hjT8EdaGUCbEIOWFnkoEckSlr6Zv9hDJsR/1MKCy3K1lyJgR7JyQ5oZuC47Z2UjPPWrRNYU
CFCfNVSSBu4r2ad/aN3CyPNSjxUFmd6ihrjwSmoiLvUpdkeJm/qdluF8KjbySIYDNqUj65yfXaTW
xkVYoajRHXM2HpSlxvb6vuK6+R6D4bbPISq2mwNLttc8tXbkVITJXxlEQ7pMy9v3QLmj7XlYnKA3
poz1lUlvuflwD9Ge6TRaVKEqQNsWxgvy84DMe92q31L8L3W3B5gh2ycJOsXCktChqrZYbN8RkIeY
oWmAn3GJluyPQgngizo3Suzqa6La0imPK/Mey4mTjicsDS1OwQBKP3ulBzYweKCIQk3fvc9zOnsL
ji6Ca4wO6l6/+BxzP1EvTmcgyjaF3X0Jl3t7UCdPupBhN4ejcGFKO3Kih5WE9wdIATX5dZsaXgY9
huw0UwwSs5qrF8/41p7HfggsTa3rAQFM75cXuQmwo44GI9Ck6eGon8AdtEDpvm8U1dbhXAm7Tm7h
gwdkutvK0i3SXE6CRtpIa7yrRys1WfbPFmSrjyhz37dhUhBCGORkzCIXofFNL2MtzyBsPO+S+pOa
YzQl/ZaN9SCjYx13G2B2d/qsBvOiL1jUq7VN8GmKHqj/Uu0AIpxVHAnXi2TVSrrtNIp6j4G4Q5Xr
KTkH7tRkOKCWSu9KeLSpwDzwy1dUIBn9eHGF0GX1ZmwPxXglcexHHu26ifYwRDvsmWj1zfz3lkOV
a6O9z0ejuxH+/MTiGHFwW5JU1IcOVXkfDmEi216NqAkjbqkxr6GcSQ5wkLG0z1wx9XhqFwwEw4rQ
5nhgSBNMbEoOrVa5GQsAXR4HMpj6LtEw8XG8uVlifXnPcHsb/NuFAiaJEg/HnnMvvgElu/WfHiTT
IsqrrEBZbVoUUdrUyGY60X8BZPKqt3FVUFVlncRlh5eswKk+KsDYEj79apiJWDb01Ole989kMFgx
3IsLdr1s7pl9svogGsZq28ZaMXw4yVQ18N5waGMEugPwv6IboN9h8MliG4gwMnVUL3PxfEw7j+/k
3TD+xTPmnIQ+Vspl7gRdazfnHGBf3xIhDEJ5Js42SeufhFMfIkKR65uYYcTgs5uF1ZBoiGpUICkt
vOGC59M+YBoWJvRQitcxruyQ5IndtLG0Ucx6/Ad0xkxXVTyHQgISDJsrqXfxB2A+i+c1+UbdZSiG
lWqsuyhZbGutBkHykAGp4dvjTdB2SV3ttL8Q3myy567VocEkDhJorCQt+1rCu6zeZk8bwwZetUYj
pbz9lBSYvNcMkcJjv61nnnMSCQOIUXS0ZdB7oC80tLW/x3yHuSaMtVkzmA64vHMb8cskpK7mXV4P
7pIOr+I/VR1mVKHHtO1effXgN6+A/QoqZf+e+m+KRMQYLo5t5Ow7T/MOGvuiMk110C6eBoAFDf2V
iaZsLVbp4xfDXWUZghmtuVui/T2eqwvYSfqXi0uc9EjS/2x16pupBQDwGR9ZDecDK7G+PDQibAEh
oFJrKGrAEjS/xSExuLXroKmiOnDgAZWSUIIKYb+mqnJy2TdAMwi37KuewmCfXR3eu4v0bh9Smwr4
RY59aTFXLuNrzr8dweIjVKmfTN85MwyrY4miK2evZeInhPRYJdMDqjPpx0Mq35Mfxs3BkLxmyXt/
tJVFHbhzemFI4Csjxe411ww+ZCg0uCPwbSQRVD7xhkROOjrUqm5Pd93HRiLDihLIC67n/4V2Rg4H
tEaFZMSWApob6DkBUXNfDndol+TwpYceUWomdT+0pJtgKdwnnQ7DgwFVZSvCqAI4TlPa9jrcRhOB
WUKoQSzvpCEMvq+yBmVErYICW1K6rR/dlyhgpO4W/x3tnrxI2rc0mswvBwIjCuOmc2YnyC0GaOB1
k8Rxa164zefjOvDgyFz+bX1sGWl681fznTz1HrtHlhB4ZYvSYpE69GigA8V3vdi//CpvfMhPf7tc
2o5TFTiqoZgINTjX777xiNZA03tPoZithzQeqDRdJCpiTVY840FnGhIC/mHlbSSE5sVGAnqT7GGp
sdoio4sMsRjeQWQoon5zo8InWikhzHiXqvQ1g1S/CCovQYawAlj1APhvkvtJRSUnqLL2ZE4pQ3xm
3NHdMqU4B1bwetILhdxT2FP7ZsiZixZg9ZbfsDVuT2ilpPNz3AOoXqwdH+NvuJGrCXknh3XM6XG8
I3GRnfMvQbOBpQ31Kfdx00bBHhibP9owkxXsz/4NwdlZt29ugJ6L1FG2coRRwI8fdRRMDmyi7V4C
9Zb1ssN4woZMgSB5JDBpIPIR9WhxFsqFKj9xZ9LRalF0oNOR9cxlxad73a8jc1WeYMZ4CzuM3qyC
2hFBTg73+Dn7+On/OSoCzD6lHdLMyWdueHWKPUS9M8Nn1BzNsM4t3Am9GtO+fjIcFVRcPIDQeIc5
NbM2gizEfm+Ys6ZhXNhrYDlaOMGmXaqD4aZE9ndYfVm3jQcHhUpVOgDZaRPKcoK05iI2ztVPCYqs
llanBp8W4wfUxPVkN0xfn5M24IybQYNWt8A3+6juOmrPb0AIVrqLFRhb0LogyeNfkDwFihX5t+dz
kYA4jvpBwnxAtrgZKnzEsj/01Coc9aq2j/NwU0eY9dnwu+KnD8FFccujGTm4C4HOteswegVPNojn
WKUZxldjFDt8/n9jXmxtrCh3/s3f3Yu64czn0E2JRF47wSOjuvs5+i5p1TbdDJ+WSEumzvXYF1U4
iGg8+rkELZr9vFEOuQErkpDvbaPtf0YERN/veAEXaUQ06m65A4zYQf4gmJ1QkAVmlZ0fw6w8zhGy
GFn25NLMBsWWRkSZFgdpZXnevhmMo5UZzeJS2TY17QmYde2qNjOg63VUG+XvqzEj4Lx20I0aAuy8
KkS/d6O//cdZ7XCSWKuNZ21aRLh6T8eoXqkK05p6zWRN56gnkJmchHk/C4Uz3KWuNj/9YWHs5rsO
N2/d7Ja9GM3KkUhJpGThxyok3Qq4e1p/ZwWDU1JNj7ibG9+nfyuVl0f6XADYZihQWcVFNI/aCGCL
X55hn5jpZ/wCdlAR0rSdPdWCpogIqkLsJ5MRUx2r66cdMEsNWCoG8wEZr/Q2j0q7R3GL+Wybfzaz
er6E+cyzf9j1uqR4K3YIah3V/qLqiu1VSLYohyqvEIVkNo/JFy3NdcTZL4OVgLE9Re1KnvGPaIQg
HNSuj0wY7O4hiEyY1h/CPJiwrjI9WKUwcLx2QJKUD+dAwmr6bggo2hnr/hVK5zmG7nc4P9A3zjvm
LwU4ZUZ/Y3arSXy31gxn4Uok6pMyS4DQEReUJZRJaqDJQyPmNdH6HfO20DlrLJv/4wDCUlb0t7Xb
cE/BvJAdhfga8EpTU2OJ/hInbI8UZWV4Ecalfs7IzGk2CJ7vxMy+mjRrN39qUwL9uGMps8yr5d0j
D8qP49o5SFo6aaNHoW04kDQqZa7pqxBP3+nF3rC8cPF4i30md0XSz5UE7WYao5Cpx8YUEudQd/i6
faBItX+dA59GAuE12WORigAg5rqLuMvFNwPih9kow44OaiByoTg8yVokzQdWEZY118bbqpgmC1jK
BZjiui/0Nxc7aOLWQqmRXZ50zOQlzvNjDKFebTVP5i6FhaHZiRU7EYxwl0c8YwSMHux6s+CWl5Q0
UcqYHTnj4TsM0lY71iFcpaw6sgyohw8BHVGNuOXLduZp7e7DeESv+mrjjY8SYzbDecMLzAldiAd2
5nZFp+BHJbw9+QlHBDj/2kVUCsY9RevVMzzSwAsoDcxBNCbTLMLYfLJj3D1ssN9wROaCx9E1cBnj
Aj2dLAnnY1CBo19KGey0gzrQeRci6NlBJyZznMh5ava6biji2n0XE1TQ6u4uML2FXBY3T4VFYBWB
5/Z7ANett0pLh5GQtNc2GYrqD7hDAn9zIbRuE2PiJ8MwJkEb3GFMXYarvhylcbrbfMQV8OXM/+F4
zP+OHv9GMMN+H5ubAHN774LkSLJ5M+8+kwMYHLM6VsMP9rXHNsLt8XEJChV6r+fRByBN9gCfDhZT
wrOoPUwGBG4PUEJHO5NoNMJLsX0RCRCFxUTVb9QH4zHycKO/6itTl6MjDZhfQRl1Bnrna06Z+xvy
XXQmjCqAIcskp7E+2feC3eXCfmJvhwhydc6dA7HmPzlvwfzKg8oNaKDJgQbnJ+Wm5+wCEym7s0qB
TxX7RWokTtt5FX/4h6GyZqxG5ifEZbRum2n0LoTUk4pkPY7C7kpX8l9bx/DetaF6qQOHP76w8zt3
OW5rDDBZGYR6DIFwS9x8GURrBS3ke9rQNyhgvES27gJXUqF66osesJmhUzH5z0745epA2SP1IPUx
0noNIC8Jbmc9os48pzh7dx+4qvIxI/3aRZztdXczzAzQnG/cYyHzA/f2haXuYYOcS9hmjyu8bGIT
FaizUqMIMdg7nmIc4tFDcq7pQsdeEdW0ROo3ooqfqiDx6aw23A36D0mxzhgqTf7nHmxSLaM/kDvS
XrH2XCOV2/LlHf4mK5LXlcxFfot+0Ct5VPX+0IvdB7n8CxSdKwCrdWBQYmYCLZVxoYdeX0dcS/aZ
oZWMVqdhw1nP0xfJLBB6jgn7Qx11FYcHRrgt5b4rfxDexT7gYfSW5kRi5eUplGOQdQ/4hxNxxAPi
5VrtwVSqMuoTTV0OJ598MYAzbORD3LkrFBCaxtoLZiNnLxEH3ducJ5F+rV3UvaKFQZlC6fhz/Jfj
uqRGman4z5bMvY46tJ23lTSpSLSaAudvgOz0NDvegPGOhyogw4W/ZrgHZbiA8PGhmSXn33hTWujy
MarcNHj6dZWaK4k/ek/RmNvOtLig8ZhcOhjWuj/p/zdaCduiuQlJ5P6jLN7hsdFQnzmPDeSiBjnG
si+JMySZNppGDKcyW3aFqi5qiJUNTMDlgfia2qWNPiTIwtzuABEb4AMyDRjutev52Dl320U1qXtd
9MBv7mONnpiscHECxeaOhMqDfUmiN9qO6dy9n0rPL9RcueWWrZ6Hp8/AhIxAcmjhTV5nW0kUhQvs
/XKRdCoNakJWuJBkTpFQfd4giBglIKtW/zACyO8hsGljoC25be1lqplbVUSS/97eJUz2T/mtpLuj
2Ojo/1+M5ApzAo9Wzd8A60UR8oWpheIaeznu22c6BKUYuQju6Az7Gf+ymJuzL1H0WjRG+brJYSTX
QdAhe2ooVoBYIglZsz4mEkojhpmoEMT0+V1RC/4K5E9S4T1wGYEEhiupoLfjDc4OdKui6QmgJBdc
TAj6UOYjjK0SFg3wVT5+lZRjlP8qeASSO8YTDfKMWvWGIT72KykkJPjXtsykjBf38zVYp4LPK7lz
3hvNFVODk/7tDN1+6EMd68Z+wZKqrLDPsOV7F4lt+OxN7eBVOz63lBsrh3UXC+IQmqJuHSuBbuZM
saV3IJw3KG8ExCOyoLmEk5gXqIkDhD6MQqJzyy852n5RyhSDpyEKyGwyW4rwekynOVkDBUGaQ2gG
7apYiwa+ex78TBIekcKMXCju7FTmfRDigH4CVTosIUaFjtqaB1KZEjz7DhdzZP/OJVyePKoU/fm3
FCBrVP1yXgL999RxwZKExxuV7hZu/daSdZ/ZWCdmTjiB2CoupJA4u4Z7wlOf/YV/uw48oceINK3K
d+Z53c+tBmsa8Qzj4/2NI89bXC+h/p7bU+gvyaF48URQP2KdyxC8WxtXJ7VIdENeM3jN/s5/VnO3
U1NecumWGuFWn/dI0kYzoJFswyuiM02zFI4bayS2HWtdVNxB//rNM1qtCupEucNZqw5a8HlNEXNG
saLsQwokVSh4ztEC1bS24aOHOX8/OlO91B34PEleHAhwpDDN7Vxqsm3mOeStUViZB8egQIFjiDSP
iiyloCHBMvCSpL3T5CuGw0E7YGmit8rzlNxCgcWYWbcsBwpRmkKyxWzZdQaEaYOCzBv63bdCOCBm
ASXt1jpUr3PF2kER+wonggVZx9V9vkiJJNPnXiehSpLqQNKdWNRa9TLCm3ABGtXkfBIyXj6Rgo1H
IN939wVQ+L20X1eZA/G63SBFgtu3GebOY3C41ec6ZAuaJb252bflKRD0Ktr4q3EYCHqHZ4cv6B9L
h1BayriDSHFGTJGkF7NZY7Z21ck8lelsZ8/ZrRgy+dizFj7wK4waQUsbnCcgubUGz5OV4CS2LrC4
43WBGbynpv+ZLC7Oxs1oP/3inFmoofDaJtwazujt053xg6kcsqUMgqnqcnf789aLgvRltIjH0FyA
6saUc1WaW1fHY9fwOZnI9+IjuDG6wo8bdJxKN80/O6skWWDguLmi4vLj0VOguFH7J9Ul1KErJ8xd
PkeJVWoQQ/0tnfKoT2JSXLkCMCujVws5HA8ei9irblE2p5nrKZu6UoU2BawdF52I3vaC1eirltmH
Med6T1fD4WpXmZ43ZQGmXAxtyYCnaSbyUfT3vk2iEEx6RRlrfELZInJi6mIeqnidZ8AoOayex29b
PV/Qu+bNUdljfaVD32KVc3bE/PO5cqgO8Hc8siFktSM1sgitiE6kx+4ldo5YZxA3KmXegfcb74lB
CMJQj96CYaVg/WSQQURebp1GATVIM3yZMR7YbK+sKROPuk7ElBpT/fuALF46glPAySDufEpkxRAG
YopeJDo5XhMdeN9e7Hz+sMAAz8LqUJR9+334tYBifcKFC1c6nUBwMxTK2Oe0X827yNwTnRWc56Oc
Alhilz1yxtKwuNxGtfv5RgWiaCYQBF2H4etH/RmCbphjhdILkhKZqPq7IcJEVcpYuJNE9Aag0I6e
GNDk1dLCLZq5BeiEgVf3NOV/uYsArJv/pvpxo4txspKLRLdoUAl2ydAMornljt18/Xid656m+ONT
U8Wbg+X8CZDd5mqUXJSV51AH8CTTaQuElGiZ+46KGpcGzEPFDxRm/uH9GqIa+13zOGYUhVlnOmsg
jq2/ncexA6ZBCuokOrdWf53xAhLeJGxPr8yAABeUDoPEAKbknt+kfnMpCyYK5cOgSeK9ViidXCkH
AdwXd4EQkG9+pMg5L4uOyzwlQv1Ux5pM3n236s2fLeeGqYapjbvOJrH8JU2YKuVnoFAHhZiO/D6O
Cf3ShrhCTrLqknE9D5qMHMkqbfcv9dSYxHjIFSIL9gHxh94z3H73EgcxP8wVxkAAuIm3ZgkSzlFk
FS7AKBHBQnUm57zdHlx2zbIvHCfPiWNbEuy8rdsKtILzickDDQDbc3cTFuYs/T5OyKyJODWcHTVQ
gceKxovFYNn8pOGN9/rb6Oe82LpWBTBlVLOWRDx8oPC3HIS8pPFBkv380MsrdAPtvhX0LHtsmZzC
FmbIuAk7ULUDSs2VRmDnOVktAopYtM16l2q7VZ8nhtmvTcEK7vDc9zfSfb38/x0d2wXkiruFzxWC
TlqtQlJo66uTEteW3Hfj/vWvxR3d7ACRSmzcSaev/6inMJHIEUQ+SJ41I8Sy+QZtpS+JIBw4zVNg
j27304hOzowEPTQstntM+JTWMfI0648YkK+pYwD01x4q2vktuc/wVwIUcAewdwfkpPUjrFhHGU3m
l32jSXu5QipF/XJGb0uEOTtb/x0ebZt9GpYOTrPDlIjtgcZYrNAesf9v5MXhr2elvUkzqhn258n9
1G6d4nGfYLxlTZKadO86PlJX3q5oP84xJf7TTKsrPTsGujU6HqOtWT7zd4JUZx1YST5gJO0gL1CS
WPjh4hFowk7joJ+voxj1x5ppz8xwSwgu3AHxQCClnRuchKcJP9fYGF5rpcvQBQshHLo4zi/7u8WJ
mbM/Ji5uQ7/8/h3dpFbAFODsMi5U9OnK2NHwey76d+hTgtDja7lK/583T/B87yKgHOv4+b0t/gRz
IeqD5bBzzqifWC5vlTtl2rcE34Ak5lR8UWFfmATGF7G9g83oGEdxtGPgX79UncvQWcuBgS7M7mKL
EihGu4dj8I82xmXMITUqbGhUPQKFWaKqsYR6I/pjAMLvkdcrKuPKbJNT4Ue5tyoegObiZHZVVXua
j7yQgxLkDWM0kZoB0skUo8UjZnN81nOgXwN81NbNDuZx1k8/btFrqcXDUUiTFZqFIhNJjEGzOKFx
fiIN63fsd9bnGDljCHvvmxMAoNMj9Np0FdRgLaVLE+Gj9p+UmR8RzbehbX7kbK216A4POLgDgIn5
LI7gwFXku+lHD4YybGqLa3juQNjtjgSwuj+fgjblbfa5XypjvzEYFLdWf+n4dTdqNq5lzHx/af3H
YVpoeY+zoD9IiRhp+9HyxNC6/eQr+gogrz2mGMpGkzGmpKE5chagwC23Z7ptVyPXQ4zCnXMtoYAF
Mo7sr+pKqOUMNanjcUQQJbgsSHk99zc4VEvEBN+gsroKgtnRgnBIg4VD/t/kc0TIyiqzKPHJ45iP
Ch8KjtLg1/592pbcxufHxP8TiKvtylVm3CTx+FkWJDLGe37xWxUHpVCKsPtzyI9WsuOQVUrtH7Df
WwWCU/p3KMvp29vyU4vzk/1Vuk80OoM1lHWQXjdIsguYF3v7+XCyVdcAEvTqK6dlyG4slGqVmRnJ
QSkGPUI6vXmP2FgEN29X2Eh0t1C+/beCwwqvXewQMt/KbA+MefzCKhZ3uG8PzjF6RhAdcIFUMLgO
OvvOLdcLQI5qwFFmDycaNe+m5FBouaPXFzUKKMewPxclxx3RopfJUW2FEH+Mj5WCptEuCOg4F3P+
sQC78JCa1hDCM9MEZxsDdMXDp6ThJDNbU33dvws+kSDi/CkaSkvmh+ANUMEWUjsB96G3DNA1+oXx
N0IScwz+tRMvp+eJIx+ubZeeqjoGjRyXd2VmmbO/cBGj0eqclOQmX+wCCi8k6MxmOeQmMw23Y+KO
7FP0mFlf4aQWS7d07b4kVMHNyHjPMBSCaC7X10zlTCQoD+EGrzToZ8s3jQ30eFUEmmkIYT3IqWUZ
7gpvAMPfvZjvTgq6Qc+llantb7HPgBV61SmXiBV/BCVCRiaE9tY4zscGiDTFXxBLQjK1UFP7hM8F
kCtKD8QYRWWhFTOZbhn/T4xmNERoAYqCaKDlfppr88QCUbMufrbbqIF9VThankQYCpZM82DxuYCc
Nx2zi5vSLcLHlcx9HlGI00XvDmRxG2SJu09LW7Y25mxmJQa55A4qMwia50XJXj6DKNfSA/tPSpS3
H1AlpouYuFLas6dvHJK0VVCQZio0W8GMedfIbOFBGtJPuI4WMCKWKnhuXsG/br3VQ1s2DS1HKteC
Y3VJrdjUcN0V+gwBenS1ko1KA23TN/XVMX2ZwmOrkcsiNrlppcI7idF22Ri+vbQPUdeDHoEqpuaV
+PxHBMRo19bZB5YdHTzESG/wLpDhd0YbjbtftC3ZdhSbWe0MYPuAd/tfVyzGlhTOVnKTr/bC3CQS
l8iiphwHa8LdvDPog1wrMVsszXo26M+M+Hddp5GZrfCFotn+vISMUFNRD/WabaWjIJ1NhYxRgPUg
O3XnOoa71q7Ok4Inf5lc4ScZEszf2fQsu+VZqoavr2b7LG9Rs9tOXVFMnWIaog1UMUe+N6z8OxLE
gv1Cpy01hNxVegJ6xasfuT4HoWPSBQ7DkpbU80uHsbS8P/GP9LuQ71d7M6zpyn1WRt/CTcXP/FWl
jHundYP8UbrQQIIrENiDFu2C087Jb2lSOQaIp5YdHlFVUhUrZOouUi5ANC68nBqv2gMewLnPUHsM
yhegwhxdFuE7tIf/PKc+x2mbmJztcpZ5lSSbm7KIABcD44MZCP8p7IBkr3A560RiphA8JM1Q+NNa
HYez+C3aYau677NBr2yvEkMQFKbUMubeO05J3CjJZCcsPuwAGr1x9+hOnbLWyzt16GzNBb2z/xjk
ms4kZylISnD6D/Q0QVFGoO2tUDvja9NJbLTICs4nIcR3XClCTKuXCzr4q+CyAAwU2Pk5ls22eIIP
raqxSTt90LrkXl6Jko9nyCZ4HK6vTtCEF2asLF86lczJZ0/Y1gw3hKuwEre6C6MQXnTMf9bnSBpy
mpz+m957SgnciuutRvlBzYomslY+3et3Qbi0gDz8gzeu6I0wuIk7x7qo1Bz4tBkjrodRWyh0JnKK
KtUbB5Keh5cFSUn4zG0ONfTyZQm/b1Be++hBZTK547yskxni0r+cydOmU2zWTw46B51jjBdT9pCx
yZBTn6wWVGwJyTRdNBpVHWSt8EQ7WfOUDyT46JxLkbEU4vqHNU9ML10xSrWxhKn8LrFgW2I5QSqT
Sa2SPkgVJO+6EJv4tGS9DJ5Hp/TDlgQrbXpbbjmKwqb38lj3tSUn/J8IB1damVVNVRF8c3DtiahX
PXL6ey60RinIf6GjGHF/2XP+ma2Hu/bNNOzN5a3zLrVEeC6eSDfqKTga4rrDEJxvGpUkIKfBvCY7
PlPp2Je49Il5VuxKZHlNls55FFvAm4U+H3se+DgisEqTEHUcYgTmmseaiy5wgzUUEB34BHvfmW+5
m2S1zTCDrbq+cBR0NYYrfRqC9yN6BJQifTzyfW7TpOiP4Ux7q61gJCDW9atcGuFSTsPDIvkNYtZx
t0ZBjhPnIxXxuWFrzNHR2Atk78j36JtjACG7FXJuy3ZE4UlPGLuLu2UVPcVroXPFzpyUjjxR0j4G
kwYp3uGnFhHtJf3T+7tgzGhnyPyxJpkVncVRuOhxh2KHQ6Qmpkz02uYRj4OI1GGIwV78afIF8n+6
hV8ARIIQQT7kFMEdoC1MICjLjSN/gK8Pr5RpYqtFqSsLo3X9jithXv4HRwBgh+4Wrhb5iWtv+BQP
Ohvulx9C+dPlwsw/kptNrhu8SAjdrIkpiaU8bV6xlG/YZukXwSXxndpGyYXgFICFnYKF2y8yYKqI
8xN0S5cf1Dl953fYPPhel/w/FloSyvhRvPlpgS5E0IWXg/XW90MferrMvGnLEj3J7v5RGeqV+XgB
tDy23N/KdqumDSRvTs8bnlxZdUCQ5xjoc2WtMUzPEDbCC7XQg7klJxLDVVcYDvmKZFYdbzFV+wOl
Hlsh1eSOSLRA5oGqfYitatWitZ572O4OPs9+VBHIHo5Wv3FoR5JAO7Cit1/1TEfgmEZW6UUDMHfl
f2bxjlV31+7FVlpoQwciQDFj/CeUd0VGrxtlqEIPtIVv4r1S6q9QkuC4qTS4WxVIcEwPLG6zNtGJ
pYkHr8kuYoOnkXlWrtphaW7Fl0X9HyXkianUwFZYQdWUbmBr3nYzs/ugJI9cChuaX6Q5l91bZ0i9
eZCMdccL12zJnUrq46/vy1JMt5t0FFxLyifRPcJc+eKUKZ27HjOMnc067T3M2ZazpkPGLLkjND43
0le2XdJo5vESG3b+iwxMAmb8TrRGEVHdsxP7RF9QnEH53De6putYO+CCOWh8zgt3kmIlsm3mYoZG
jKzyLiabYnjBMcWtkCm8of4yQWj+2SfWDqLyUJ5tPYNuPmZ9o9s9FNjxZ7RhZp/jSHXWSGuKzTj0
F0mZ8Dq2KCjROlYwC2OIqYwCFn0qU4+xwQuw8GQLF1MARgxs4ZGZHTYSAwYOR7217RDryFktTqK1
rKA4JXUHQd9GC93rGFx6u58RjqqKmmEFRu2dunYhnqXpq0qCN5k3obPxyvsRExLGVZf+0+AMgr9F
yPrmBTzeABrXD1R2ywnV+QZu40hlb6XF6z66SQlNFBcHm6rxHb8+yufh9dD7EJgpLaMwGc+GYWsJ
NwJZM2IBG/5ru1FJ3PLUxJdNWkTjDtb7eSr5OPQSlrHQjUs60lxlyQafyhqv+aGBbfKSrhH6qg45
Of5uEF2jKbYBUcIxg4Sx4ta5+bXETKavbISgjAVClvkciPLg79rxr6mUbhFFDuL7LMfVnJH803dY
s+jM6tw1hQ6zMVf174fs/iyd0XF0fwOpO8HKs4I1lqIMn+svgZd1U88HWZR4/RwHtzju4v1uz29a
oaORJ+m8MIM5645/9Yd2Ll0CvxSfLLgja3FFYjIzYFN6rKBp7ex9war04sf1dTgOD7j2fV5wRllw
0Kc8WTaPIP570znL+HUh9uTnV1xx1yfZUDxZoLZzEGiK1I2y6s+z64Oz3J/052s/3qq2atGWWpDP
izt7IIr2mIGumHjNiZ4YSv9e6gqu0kyTB4zd4qXONiE8yyFGcewk56cLk87dennPknROPOSStX9A
gggKA1URLy8T7Xf+jZTsbP/ZmAmCTOKCE0C2kl+x54516bWAM0XXWZa4J2uFG1N2NaunuEoOpuNc
dkHrT0tKPcWtdKmLnKWaXhE3jYpI0+djebPzNrWjS+yhg4HXGbQBX42XMsuO03rEZZY8RzWoQMBK
rbF+75uIsQyCdiNPDtMNsI/3nXaudZ7P315GeQ6QZgqUCb6cju+mFDPOTbs8uWVTIuTQqzXmKCiS
GqbIf6gC4QxdTTQo8e5glxSPzggototLdtTZeEghiUlX81egkxvHWInHMGEUopUkM8ufeQk1RMh5
jg77oa52U/U9HvH9Qphq66BLHVll7Xf0tEkHMzVNw3fBtnXx46SHIur0/hi6oFxXTbjus7vcsGvE
Ah2nRhmlm33iTk3ard0yqVfOs6GqGmww0yUlOmfoOyz2ShCqe/pn54CjFP2u6ahgONIsvyJDIK0i
01t7bnndRDYGWuEDqPw1JrFfeSYLvmKbwLadlDSNCKgIhBupq+RIzu+xL2JQKCrIiO3hjv7P77or
15DJQj6eLJOFlsvaa1ogBNEZRfLobVkfQ0iSaW+4dqj21YgW4R/HYLiWrjCe79nN12mDTLoU+vks
aPbTFeZmDDwDKwgG7c22hyy9BiBcz4MDoinnCpDGxM8BmMTQzsQkoJ6fkz+WcMMjwl+QFAj3TByG
cSbiPw7UCcAbhQcNrK9mekna5aXfeHuSCxeIjFft3A7Kw7ts5wACmq+V9RO7aMTkhJMMjNnZWMLX
KjQ3Ga98wd9ipJkAVkoHK5qXsysD1OM5NIEmHKitKajYuwPApee+TC47AKKwLJmeE8SMwj50OmXs
KrPqzqlqB5Pzmh4Nj8rIyWaTiTJeGUfIVhZm/YMhqc/SelpA+9ZZp7dh/DGBkDGbUYe3r0TWxa7D
/Nw1dz0RCuI1YM7MNGlWg2In2f6iUV0ykJB+Fw4+IStD13w7+zgx/gwIwAfKPxpTlwQetEV13F6L
PyushYaCWG08BUpLvpj2T0/5DM2oQLYZBGWT41/f5Z6yNXz4mixTPQCkHCCEEnUnms0Z8udqawtR
WICgPUG8z0yJnFwhfPkAUaw9UKeuKDL9bn5yy8YJuSNVt4pm5olZzp9IUViN5GOJ5Su8bgSbfqPe
xcXoY3Z4a9L/6PQUKXo+1+FGrFjR3alcLfDsbLCFTQaUinkCcynRoVHpDA944a7gv3rqKLfT3DIe
4XikyGkjj/DGBVKd3p9LscS8drA0Q6ujjbR76I8UZ7YGbzvun06GlM+oIC8SHg6qxpbXharN40S0
i655rnjrgIbe2uR1x1afacYRGamPeEZvlYaBqlC6dwMFuK/wiPqiw/XZGp5HCr745cBgzqSNJZst
EJ+I7Qd3xBk7pe0K8FpwzPUxQlCCj5oK/+0DQZOI5A+cfcDy2O61p1SqzP7fLnRn4ZbvGuZ57SmZ
ryv1FW0c1FVgf4q5k7IgZsjSqclkdG3gMxFAABY4XKBnA93wNJpJpgOdXgy6Nd3MITIWhk7NbtC3
CLALpP/FI2XIoCiWTVFMIQbr8JUgUYNUM1FQW5bNfFOiL8fxp+MNDMVKL9ZLYD1x7TbSrFHXyQe4
Jl4MD4y4NYYvZZ91ZhEWCSPKcGH/e/ZUSAPjLZAbbNZU60aIsN8iKVAWQX5evAu9/ZNFOJYYWoE3
DZViNONTk9iJ3JmThWDV97e4zCXW57rDjLi2544Moc+a61wQ2XfE6z7W4NiSwjHD282TxQSVrM9w
3Gtz7AO2yF2k7jWZHFhH+/aK68ziKsM4pSamoETvPk3BpIhg5JYNWDQBPuRrMsBe82g8FrtJeAI9
PfbIs0GZMU+/EG2Szql//cUzJMi+HmtgxzqWObOD49tsKZI1mSnfEsQD0qrK2r93jYR+5+DjtNVx
AJb375g/vGPXjGDDih1uxPy6mT9DVJcnniUwPUhZ2qobBTmjPhkvAU5n92blK6nQBez4sTBdbLUu
bWIDSw0ELMzBnxVSG77FAeyR5SDJvaYROPWsmrq+SCABZ+OLT/+d8HorD4bS7bxohpO5R1QeccHh
5TBjPztk4nlw1iS9gHa/PdYkgu+HDBdRN1NUtoAiYJpFcDogcXs8S0+IMb4xQRSgphQMyKRMDNOd
x619mEaj2PusxKZprUtzIaCLqPEuB59Hx+LjKlUsB57ZGWopJnxRzGn2I8yH2GE72thrshNInooc
4actg44ipGC6iQgbLizm6GxLnvW8fD1Q7avtPJhcGDXuYOv3X9hr8tBP+6EU9PsX8Rrij+bok5/h
qbcDu8tOUY8j+0P1fBsagfOUjWlcKy8TiK6Qj7fPcbGnnrdhO6yyN9dssxoPkuZfZr70xd1Q3Cck
Oni6M7sazW6zddrIJpKeFk7oJjUN3QGU4k5uEq3+ahU2WmvVpjVOXj2GRZkVHYpcksWz5BHKNg3N
N9QY3kfu9RdLWEFzzktGziOf/QKZSkv0plIoxQzD9sbxi3dLBE4Qib31CAMWqbWOedsrkMumX1Zy
tlInOkZSMlg4lJ49SP09MmOuUTSVCYs3hh9+tA6o45n7jQS92UQ3JVmIqAt96aBcc+52rtde7ecN
zw7/PqKeJ1KY4gLZMT1Q1d3DBTRlEoFzMXtozgyyOgoXlEH61YqILaQCJ7QPqSbDMTGY1ToHkx6B
HjjBKDQDvB+4V3NB7t/TD4+u0RO0o7Dur9Iq8PKA+AanUETb7uixA4BdcqchDBjOaA4hMHUxmQI0
4sYq8Q/Y2lj6dFyYVz6JVaD3idT31Sw1+zkGB0C28hvvbC4Je7Xe1vhSBpODZllom+gtveRNRtCA
fm69d0jEBcL1f7ET0W/lqJBr7pRjdUxcJeQUj6jGSSwza2mEWUC5fEMPBIEPhDaiNNlQo+mpB/PZ
0Db7LFPw+nw2HBEy6ptbbqhSJ9FrXFIhB7yBYH2+A+RZKENUgf10xBANDAmHTZDDuPaR7AUA3c0T
lFMFyrK4ZBdD/SYIyZBkcbQCBh+kATaCvFo5v6iRZSGKIQbbAhl41xpxkiLv8mkOeG1l/aksZ4Q6
4qdz+6MXtPoYMx81TDZ6ZmlzaGX3DBOlWmJjmmps7RL6LFArF+BvOIHE1Cjc0h0XUiN6i+JDH2yG
d4ZpQso9us4WbJQwXcuFrWS4np3xJx0fTsqdflH7qedLgI089a9JgL55wHcf9KProqGPw9u9AlAO
HdkGcFp49g/ddqMkgUYUYyAGh7yu1bDtH1ZAuf5/p4vLN5hxBaqhSERBO7zqugKTFEEYY6lFRr7A
JHVzi2VGjOBoFLda4tYb45ejeScluanzeGavNFdnxPtim+NP7yJ4d6ZgGNMIpav246f6DusRbxLE
X9BBeX0oHPcKzPAzMRBYXBd2l8L4UadiI1NJMEzm58K3vCsg9Unuq+xB54Pow3EFIVUrsPj90dCO
WjNsWyVACJ9K2YWclEqTqfphyPoKXxjQ8X5GNkgH1hRAnQxAF2r0hogB9Tuwu6nBrPTtUH1LXynM
yFVwziAb7CZj9GAvEqFhe6wmlb73739ZrAt2UQ0Kj0quC2Rkv7lTFdcTd6Qvu0AnpnYPSAUVFiQv
IuNdEX06o4AbdTAANj26BLxyYylFKPRF3xG6X1UP1TLPlN37p6xOS/ri3cy7VnFRo6bj7+N6JcHe
t4H7oCV3ZUUOGaWvjgGgJEGKtJ2lMi2sQZHBwSihj1DjNpsjT53RS4SRRxUMH6YLzqYKmnYSkayu
dOxgoi8/DcDwhKxLxXflJKaQN5Jq4BWMYxrlGS0BiPv8yFxgkm+GyCUWCeU4iTqOItfHt5CacT9l
awZVntcrr0Nohy7QjCpupCxKzkVelYliy4SX4fQVb78qd73l34ZFUIcO4yW41W8gL88kelQUTMFN
/CvUiAV5KJstUWSfz0Lighuwnn85bJZPqzzytKYnvGTzxLnCKRHjhoffpsUH6gLf9RrSLwTpoHWk
i4gCrTQ708jui/WjLzhJNshzsOQ6i8WRmKw9e77s7E+alw8lr2q52O/fCFoPxLOu3hKNncBbAmqo
NDkjwUJb0yxF51dUStG5ooa/8s4teuPt9V2QtrvZ2hz+XyX+P4ZNdVrRZ9Qy7mNqGJWlxywUsUJE
SRkpioIhoErGOpDrERYbnPtsMSKhxX/JVgLbrtV+MRWbK/w5Tj3K8NlE7CN8H5CeXdn0PsusliCN
W9ZwsMNYoKc4kgiuCbNWZzyGo48IpQSg6CSLNdjg6Tr2YzJlGU2MxZukviJt5Totr7R4hugBSMtl
D3mcSh482dn2+BaqnjhpgNmlGSSZhgd74uS5Qac1f+2PDRrBlxQ8zxnM7ZHsBpSW7A3sN2R5+1Wq
P7bFCTUxvTze+E7zDIjrLbLCOd89Qm+zeuILPlXT4FhXoY7yCDDyF8+m8QumIOa39LXY5S75ZP6+
WuHP8DHuV714BSTEn1UH6BmR5yXlX8mJCJnfsGPF7AwKSX2Bc+kty/1Glwo0bsHK+b/t/bjKUMIB
8VrqJMyI8WCOPCsGko3vdHlcwy4Mk1I3a6zo7x0qeEnA99nKE58vIsYaInZVPKO03Fh712JUBxTc
FW+ywhWN4s8LBBnZzy3WZ2NbDRznqiv+sA2jG3GRFHsJXfKJg5/Wn2bMTLTvqJ0d/Anq9U09mTXw
wdHy4XLfUY/ZggfY7Aw4Lu3fFx5xEedFQ+GxinUbewHUq3uNUVSw74+h0qCL+XjPUFh1ReWimrJo
tSuBD1gWlExkSpnMCDDHiIFNwkjrSyjxYgWI/rSQ2fBFwOdHhiCqPBXo16XG8Jv94m3K/86yx+YJ
PmZAG2rnexq0glC5w3NXoy7i2u2z1pq4PbybdWSTnOXl+Px8j5WhuHjGC255zKemqOH70l7x6qqf
gVYqIJuHnv0u7VeG8qz7Vo4V2yQGJcgypiY35DPTnnBtQbCYkbFFyeWnTXwNckDoyb5miPVW6tRE
33/AK0zVTbY1X859BG7Wr1UVzBvFOSRBiJ6Xcw9vXaTziTepHWKpoHN7y2zlz8IHZ1RWJFqQ39+d
6OP7h/0y2etTsXq+ucrUQrPK5DQM0f6ESBkf96kHTboFKKdehvLPPErtPM0P5XozTULapCz7jkfN
xvlLnsvW7ceA7Tadio76y4c/XxnEwb6wWRjpPXIjqMCHoUk8FAgAmUdTV+iY1EzPhZhrZF1yyEvw
3NrcmSFZAtEMV+aHclIabKyhWGndEH2L2WgjSD5b0GLy9KYsOitb/y5WRsZYD40z7dWJRUDHdO7E
g38zeZfNausdl2RHKIfTS54b1ygulk5Zyn7q1il0HPPa7mQ/ol0LAdxWhoPlmYTdMK2ALhzFXvnP
uAFgGb5pVOh48xhVOamaSQ+VL+Ffj6Jr7+8JV0soUjdtVfZg4c7sI1LsglMdiYoJ85CrLabBplF/
7drdEdaBVNyLkIKyfGimjTs/1eYDJnyYauO6MR0/4HfHaYLUzwZ5x2HQx0S/FgodpOO04vFvr8Vk
et4rtCqzIc8fKUOqPZ7ev2sA5r/xuRdxAjiT3AuY8zcoRUT+9zPD03SoMr7rFd+1dHKnvhapUxbB
UdAga2YXtj63jQZ6RMgSbccrhKuWzIE0HCcq85o2HBWcGgiLzwqrO4YfFLZ+FkQLQ0wFTqAWVpPO
vant5RXapxO0aC1tCfVxaxUaPio47n2+hXV7Z6sePzzsoDsaf7BRKir5zqtBH+PaRl3jwrSTQRtY
T7vIZ1JxXLF4J5tCyeudFChqZEYinvf2msqKNy2GXCkZ0CcNsKWxfSk3i6/DfDNR5ygoJCrS0Fhx
xgg/68nGGPEWzA/4lDA0cBJzIsgVQB+LYlWq7oGqM6JJr427VHD/lvcAv5RKsMnOGrEKrfbo2D5E
8xwcwt0a6sUjPXp1tIEtmcC0rhemMj6KJc1BfIdfnmZf9jjh7mgV8kOmjI1k/eZxsVEGMBfKEhya
H6wfHnpnGAXHxUk3LnFL5qsepMlsXLQwuipyJZKjdVGb97wbd2Uwqa3mJioCjDxMQz9FsL7atix8
qiUQR0s7EMcDLoLjs6gl4JKBGE6ki18jG0n82gfo8AysXEYAOJlGKW/ZbQWMU+7ej79la4u+OKa+
LHxpPUOTABdk0YXbVWmzAkkChFEwEW5B0DG3Z6yk0io+QnPVeDpADxwGTmq9Bg/Uq0skNcUxkCUX
9GeEyhs30nIPw2Jo9VA5GA56qL21qjOmW4WptakiOypikfGKqy2aLVbxb/0cTihwzwXsnRDRCWHn
4yhwETMGMn9WzwNaqUVAyFJOuKTTVi/lWU0HaYm3/urksTaCxkVOCWxrmqHYb38lqh63o+wkrv4r
AfwLEfdQCu/Sy7FIP4KfSywZn4d109VfOTVFXNdrTw2CKmU2O7nRnh/IiUU5WDVUTF5ogo96uKDi
3b20EIDj4ypLrWEQZzbbeZFIyVURmw2MjYdFR8PgejJPGkGhC4kTs3VHIWL8yFtuTIN9MLGKBSW0
H/j101mkQptyDcQr3xwTSUicSVxbLBQqiDnXVhCSeJ2uD5GkHgxdZiB4siCgWQLu6euwho7Hv6y6
Ai/MqnkYA8IM9s4BXcLj/eP1KAcwT3A9ulADW88x579LBMkN+w2vlLVFwhbd6/dsUy6oJJyXERwO
kIRau3M7tw3S6blig3qP8mnE/U2xd8S4bH+sxKGH0rVF1uBvj0IZLM08/opRmw8BUZrodIq3rBBz
tnvihDx3yQiHR0+TaTtYb7zHIH1TGIEmE4sJc+tcvsl+k6FSYzbd/djXfPotp1YZQ8iZTA48Kw1q
7Y1P5QK39Z7upUL2rocH9D1bNBihdNWQUF34ezIvYZFYWwjPo7G+P2wzQzKxFDBeKwlS/jipKLIP
3zXv3MwgYSoc1xaXrlCtnYMj1QgzLmE7UNs5+Rh9pG43RhlZXZy+Xs8uJy4K/ZZEBd1SadO/iUpx
GkeEsVr9H23Tae2uesi5DkYfM1w1FtGN5nHQkA2Zg5rmamZ2t5uocXh/USjOoBEKHoUJsmVcIvJW
mbW2QMT+ZzypEDts/0emXw5yEwi1Nj0Q4tom8cEB+4gnpPX0j0uLvKRHVZyx4lvmuvLGEv/p/Cbp
xiW7HqoqIc17hCaxfl/y9FYdJnUc3Ps+0mSrT11n7cUbozzQuuIkiEXD4whMqy/hJlOPKep54qWe
mFQgxm0XII2L21ZVxElhsxO3SDIK/8N8ShdoFi9nWeWqzhlythiCgClO/ad4Az3INQAi/3I/Qquu
7hrgdW7DlV7NmwEUEXC2ib3kA5F7ORPvcbxYBUkCXIG7ATyboGSLT6euIZM8urCGj6AQnRtP3RPt
/lIJk/WlxlAN/JEzLGtE7Ow+izpeUzICywdSN4M0PMl8UUmC5qIQUzUQboewYYhZ3x108JQowktK
162olOM9un6v98f9UT90w7VO/YOZUdlGsRMISSkeKJlLhLbot5xDg/O0o5CJYu1E7KYjSvtKoRoA
rCtnWvk1Vjin78+F2KB6t0nJdsonbflI6cm6wYjuL7zcvHtBm8yQMj8v5tcIF2kHLWA7RBsb0KAW
eQ3M/acInQlmGMVvCQpvsSs3XWxrazEXmePR902x0AgbDkZwTLAmla+a+inYy8TswHhv7wc40ITU
cao52WPRYIQQvEweQi3ryyFg5m9kzxVbJjzUY59q8Eq3Mxr1Qhnc67fvy9Ndpad/WPR+j1TlLcZw
sieN+LHEgAjw1pbUrxI6b9SOZvnYGol7c5w9gyXP+wILiCji69hFSdSLRxYXqaTBouGS6WAGnT0f
XDAZlPyR1OUqf3YX8e+/jz+J/8oABFq6CmDvGbJ0bmTRVHbe0FHLxGmEoTkmVLb59gAnS/CsuCEQ
sbZPQ+mJIIMRFToH47tXJukuPFNy0JiQJ7jnXishCJqRjL5bQzfTALQfNxJ+qyab9X7ZGKpKnty4
+vSiMHrWsrG5yGZIFPZfhZoA63Jt20R0cBHj1G/kUL9sbErgIz3NHEHehXWHIOvvWwsDd0TjEFIi
2gm86yMSO0tNdIgAeU1doyQ5Cy5b/gX8ckNT4/kENh/DCvj2IIo0QzpnQo2p4mgdWhaf716qmtNL
MPe9FlHM7+sSiXvAlzMj4ga7ZdNKe3sDPsdB2++Wk0L2YhnadVS59J+jIIF1O7CDj63Bh8AP7t16
wSbZ9PscFaYnBH5RskA2ybS5xLVPro0GZ9CVWO0PRusaF5wwSXtd+Ebp593oJ7cjDaKqEvGeu50Y
8ItmkqLUgx9BlR6D/iy+sYwh63wri07PfRPrP1V0mi5+d5ciXPVcKqex5kTZGXshKxUEe+0PGGpa
yfSAkQj00M1LBRHRulKFnbEjT1LL8KHgoHAbRw9XngP5fLOFi2lDKexE3X54JvARIBgY6X/3pXPV
tlLJPuv7P374I/WN6QgW0SPdPX1xj3LZCrnnuKtWz1rsoucYevoBfVXNM4RJXLtHGCYqaSLE8afI
ShhpB7y+KSP0QVGrHwGfIcVpZR6QwxjTYJB5Fo/8N2O/n/brbe1PnT3Y4db7XAtlaHfA5psjlcgh
F9aUJJxBDxEXC4Cmffe2eK0pqJMg4rY3bc0liu1gwxVCEN1l+mY9qKJSZvB3f53dJf/NfHAMg4xh
YFzTC0Z+eCn3xlggyiTolZxsZmOtEP+1pFL6pbf3xMf5Ht/I10Mg5yZiOOsxv+s77jtBIp5mBhyA
7OcCvrG2ysti5SAGOLhhHXZ/3FuNhXVfJjsG7dWzC1wi/tArik/j6vlWUn9cotuIteQvj3t3QN3j
MccKwhul6N5D8Dqp+0Inix3XcNL4VGGCbI6+FKir0pOh59dg8EDgQDF135CFWF5L5NktjZxdqNyx
amWXQJpKPJglX8KNA51o4KNOCI3dRucFOwDQ1BtqWxiBRcAnPrzQMKCLRpHbazjzZwbCQQN0wltB
FpYfarzXRof9iUFAT5HMHeSHXt9ueRc16tq0pU6hxmg0B2yWkXtEccjDoOp4XaQY1Mj1RWqqPyc1
nw/QioqQe1qWRQ56xMDzCK60kOWrh0gtX6YW237qOrdckTO36jwo9+jDX/yjkCXd2fTEq+k9r+TJ
UEZAbv5da9nPcP18Q8bkOOOdiAjXBrjnvu70W5Yv8nikiMGd6SqNTi6m/ptRLrDxMO651nl+ak7p
iem7V1ErAsRE9VOi7fItGhY5sEg+gQXZiV0nxq1PXVrX/DXJIfX5uFK17k8KjTDicCEiiaHbijtr
6mFhfaE7kZSwlia4vjo7TGafpjV+eDF1yP2ezIu+iF3iRy8FaWeLk5xqLx2C4GfYkkH4h2EL+BH9
Gwps2bHtwToHagf/TrbFa9e80268e6bLqsN7NA/FmVUadI5i1B7Ot6D6B9pz5jJ7jZK7FEy0xEyR
pKVwJ5ReN59tFswzUzewuTnSc6/+3Fg5jqcs8/QelBanbrXyY/9POvBIq+t5AZIWTzb3JUdEzUcV
3KpuH8y+0dM+U1pGnKqT7+qpT1aP3eP8QdH2i4c5UtE0t/+kzPphJX7RAvV22dCaUvcm0/Tm2k30
IlXdvjMDb+zbw4xAZCFDs7qNc9fco36QGHW69Wgqu1JBngH+EiD6HmdOKYXI2f1dL6OIDHZ600EV
Kw8orxjvLbQOayTePHMjt1qRWWS4dbzdH/6uSaYV0xtYltAsp3xP/BTInm0ePRj2PxNmHDa9JEia
Z7vgT8p0JKKi9xSjx3V3Z/gMqWV8bEYNtSV15B+mTrjexX0dZGQtECz1yQlgSnhHouBTzefAmmXO
B9w7cnj9s3dqnuPPeWLrTrmZyt3BeOA+FrQN5U81T5TWQBCsqJ3TIQnh8yS/vjGvE93SLxrNdhQb
eqalaI1XrRzyRPQE0BQ7bFEjNrHxmn6a5nwDfOM1eQJQe5O88XG0fCB+X1IY8T5oEZ99+BjO5frH
xVX48qv5tVfn1iYNr7hipPIjHzetLH3K9XmJ5J39+u88Qcj09+POw8bNXb+70/1Ty84ozfHr+Pc0
fUqGCEDWJw2JqHA2mvcse2uuoTBtuZZlwyN9WhOCyZGFrTBa6eYCDDwfj2mbYmLqlhLrtnQioOnr
11RYqznr05uRXGiD2fA8KF0XeT5mdbAO2OhQSB9RSxUI0SxBDZ2d/8Z/3hgRftB5l93VH+6lE8Vg
iTROIf/YLZQlHExIhG2V92gAausET7LHcNCvPG1ROHIeGB0PVTRB9WRVSO2DSNu04eIE57dtwaPs
T/B0tj9RK1uVSTPxgUTi4l88XaQfzKggAkqEh6oKgc9IIEvefygxTbiZxYMFajWN4vcQOo8nQn1J
Fk1/a+An7do50hCCh9bMkKxLaMspzBPoEteEWwKqWL2ouR6FcJKwVpz4C7rz0KFFq5TRXbzvYxM5
n29Y+iyaxNwvAquIb6xw1HvV277vr/5nF2aQFCS39QrH1qB3lDM1DsIBiWYACzteULbolR0ijRen
SywipqW2QOAs7fvyxeMYuVxoYqR1v0qzZPwuiwoHDyjtU4g3rC6C1f2nnYOqF/E89WiC4XTROi7F
jnVppHgAVWH9HDfLlQ9aKCbwo+STfy6qmXRjvS+LByauLCxPl6/MrqMcPBjHv5GqbpgX8Q7b3wbJ
HfidEHZHgURvDqWAH6mCG+GV/n/l+JnDuZIL2Lnjprm1+ltukhi4hJZFg2B488P4XDcEH28bp314
wdV9GUrKue87eIjIKcLIY7DSrD4wQnyZH81FQc4p117TTiqJTgrDMeBp/DgqPpWGvLvNe+awos24
QMgB1ujdGtrOoLtNPL3vESZ6uleXgrfeElRpW9hXj5KW5uPgByI18Mh1g74/8rTIJL7jjREzpSGN
g+UoLsAoBloWWFWLBl5FpKLRe+Fs2T3f5JRWPyN37aYdsJ1kyPew0lgvSNPYS9wnjv5RpaTexy2n
ZOpsYrfUOvZ8+AXDfrBD7zX33u2oZLljGn70NUmWSGHKBdoYvQgx/i9ApYWwaFLZEDoChz43cJqm
vAEirTbHVE2shueyPK/rat1BDM987vmL3mtIoJev1vLeXjZ6f+i1amdOaW/fPiYW9HBNMyGzzJ1l
mY5eDFW8knDleBLx7r++aGxSkYYTodEeWC7h0rzsz7fbh6ittq0eLDcp3vVtLzy/WbSaRl/eqsjW
w+v+5PFLT1TcesTzZWYkngEDpyVNqPEtMJatIsXwIrf8o4S3F6JxSfeUMYU+7QrgKUMN+6Ciskgq
h4tEfiNONmMU0csWKlYnQ497sqbJpro/ZSuPbO+SQ55qGeh/LxurhtPh3U92pvx8FASOJCdDNfCz
UDHyjFRhFM56+DLL0Qcy6ZpwtgkF+Hq46+bC9A/t9HjRaOiaRAi8qO3JGaU9di2+oQN19NtHsiAW
FW39dZZs0AfV8DevbHoLWMe/i1xf6jXm5eWAemJKilT4sy5Kc72ir9M6CTfnnEGltzOSIozxyoXw
1NVRcpjOcPARzpAaYL3aMs4q17K7+3rG4I/6sspGwOFHAm2XGpuNXFF9I/z9ku+OsuMqxenEeyRJ
O7kChtn9UOPLj7w5X4NFtxAtWJrXF5mMXbdknF7mi07EgFdUmN+375vFP3lf7wHOK1Arjshb8Qb/
dBypn17sovPHad2muTRWlC/gwElBvB0drhM5ucItlonch+u0gaO6jUvKL5X62CEGacMMsV8Iht/g
OILOS+QmH2Dls4fhMrpzQKYOWC7XUUDqSp/I2J1aeYq4s0VF5agbV2jq9b5h01m4NFacC86vLvNW
bIpfcafiFfWH/lRlnIPlj6GP80sJ3XTPyKrbVKwGWjRpNJc6XDpEN+jUGGrFeiT70xxfVzXgm5Ws
xpseZHgYSG5ANMv00qwEATCri9RstsW0Gof4qPHqzFnpyTHJsk4ljAY98Gma4oJOs5w4g/iLp6ca
nfFNtMv65eRwB/m7CoQ1nXo1BWHgPo2SriYzq6NjkECHROROdqv4dLi4GklfPVPDFKJSKFVrAKT1
mcWI6pwt4nioft6u3LY4f5xchlXAgkr9absxdQVKQHhdOvo8PJZjXzxj7Ry+hOTZJiBGNbuOptWX
FpCUGJVfw8sjkIw3y+CqgBv9MCvVmvM1DfCAJtLQ4kCILrZXxA2npmpISXrcTcKzO5sUKODZcOP+
C5UmlzQB9fVrgAevebR/15KV0IxDZbKbZtGjsIosjNOIHGyZmXUjVG7n6vowJGR0nW8zntMKgcBo
0ra4hGVd6orSyw7jK0EZiFeQBwZ6E5pIfSUQm/Z9h7ZgrC9idt97gY5cyt46ufRg8ibLvdUifFP1
W3klvvMneLtmgGYroE5Gsnll0oa3Ow4jWv47b39wn5hZYLO1W3JA3ELW4K4cd/Ss0FFUIY2jDbzK
T1EJHjQ2wW49VLo2viZDYQ7QM17yUlouXvay/L+XBIgTk+t0MaLP5VvEu/uUTGgXB88dsT+RPEW/
8J0Ds5NK1A8wl72mj8oxW4TzD6rvc5fn5md97ez4Gr+QKCYZXHE+7QinxUvYwjdYgoY5yeagRUCJ
hCjMhFyK999uo8AJZiHbsItwIy1XPBL5iirAb64riESVTuL+y3f9/SR62CuOtypAVg7ujeJgzhrI
5iNBenioqMCjsoDCeiGmVwh/st/T1G29uCqAdkIjL5Y/qTyEJe3jUsFae782xiUIGqG4UA/tC/UQ
fYAMAYlkNzD+jC1oXxVVuKimGXdtXNM+FOFJx9E4ioGm2N0qDrDDbYq8Q5H2htgTt3oOqxPHc8/S
LoLBr5k3hfQjlibJqKlPze1FJZ+/kvYtRa/nN+21JhxgGeN/M/FFbg4LP3MU3PXnoj2zqb8BiJSc
mahMysmBw/P+mZUNud7Jl6waijOyEphFv9YH4vrMW+7jALu5TTElOnHF4/p/3IGOE72W/q2gOnLy
gs8sql+vbuyG6nDS+oWIsedeGVfSFJfO35vABGeSl/9zx238u3kdsPi2rYfSFjyeAYaLynEYSYrO
K+PjU8Wi7n/+ZT50k2zbfmzBtL6uALdScuFZt4H62l0tMqkfGKqpe0mPi3nLn/4eR1JZ2rJPcFAx
POsDtZukzxSwmoJaHYSGP26xHgdH+oVxxkxxxdCP7UiC5p7C3WAkRZXKTAPU7ziWwZeodIjG6KvV
sPPaONI4x7QRepaq3cr+o14aK0/hUe6h8Bb++koBoUvBcmSXI3135jHrnXEonIgAVS9G5L3h1BSi
sOZmzBfL/DTQcZRA1fyvkD1n7f3H8pKSwcN6qlbJLLC1EQFL8gvTVDk5Q1u+iDTJ2KrBGGb57CrH
71okKmgTEmAc7Tni51KyVbTBSbGw5PvtX4tTfpjh1Hy4MkUyxUGsdYLIxEGHfaiwAWQMvTDBf7PA
2kfcXpDbzEMcINf0wlQZI5xCD4rOzxo6mp8SfdtwcgFP+KxseiIkFfegdJr5V500ExEY2vL9Qukj
UWrMH43veLLUFQnFmDHfpMwm4R6EQ2HjqWKysMSErIpUL3RI+WDzIDOHm9Mx9/rn15o/mPNVaawZ
ieoQsy2U06LklVoUyg0NhB0+c0gQVg8YKi8oIpM2fAC/qsKfmonL79jcxOXKkldUmkwM80mMpk8x
UcEY/DJheLcJJMu8fSI3VMOy4fNlCR1mtR+rnxcUifE3szcK9KvClKjII59130GBLbaiEk/2d5wU
Kkqx2ENfoB7ttbKw+Gjd+SVdBQ95w/WhgJrp8InK26Loyd73dAuQ14+sxtw+UzEA17VRTgSMFF5R
KVsGEO/3Fe0fnncLapr8ZyIzCctWcbmDJZOSPKdMgDmnDWjUhwlFBchGiSd5V/rkM7Q5QHMe7e6a
zMm7kSfLh7KaABHCzHpWJbfmltjDK3eDKoEjHf7GhgpOvEGosboUus5mNJ8nNApSUu58ddvFS0Bc
DGzpibBwYedfhsHSqpN2NVUCWuvhkqzKtdksIvWYIfVoKQeeZ6AJNgJw/AUOq6EtA2ygfRh7VtPB
jFezjLSNFgIZaR5rtZdUvkKa/vGsvX+9wJqCK1x0wQ7EZM938nh8U5fRvIIT3sTqzjwxzcUaW4rc
ZGgY8T6qsSucmlL09GY+KL12cvq4gDjlWsJXomS8VP7tXvQX2KW5ZiNnGsff/aj2FSB19LQfC5jv
x+yqKJ3cRZeUcb+ONtOWsKK6n2dRjl0RHMKBydMDkjwh7b4Ed07XjouefC1kCkAe/nXJDh0L4HTU
993NE+evJ936eIsKhXE0eEOWhSgQTbxsM226NwRipjeHqLy9HWbYQvVlIOtMsMpmexvwLK1JQl74
jqIvIB+Yn8SNQedyFi1m/8hcjLQLXBRw7MY55mQIAiPh+xhWZEbyoLSv1grQZid7OiD6C0J41vuG
hJllJzK/OAJ6QjdKR5Z3UnPIHUgjBB7CU0qJ6u6570TVai1BeU+y1YQifJ0r0xroaOSBV8/i2c/u
5QKWPNSQ/2iqIVkUm4aXsOHlyPLChl2SKx/2SUupIP5b+fU+gYSuM52ywx4OZYKOg8lus1hOoAyW
AOBdyDZt1H1eWgh1z9/oHBw+QBXCvAUUVSUaYVV5Gah6zinYYl0LSoer3CGiSGMgcd4Pn2UhK3NS
S3tD+Mvp25o+tGbDFPWIddODn5wQ+qBQlH+qsqFfsq+/MKkflVjGFBoqLpIM4sCdvK8iI1hr5dEf
cMAPAkpLtFK7tqjW/TarabPBIzrr4CTxsDWV+TcOA56YDT8TYc9oIadwaoRsOIuuYJjNIPImSM2D
6b/QANMFdohJeV6qrDDk7dGkXPLiCxkLOQDe2cf7ymlmm95GDnkC2t0005QZkgMqxv9hpjY/y6UD
CVUIPy23TKdcJ/VZT55fVQYWd8DN8fDluDajSiw6fvytBT9GO074QN81UdOxsED3YQ6hOgc8KKSO
6MbjRlr/UmvsmeyMawCpRfT889YiD81qM6qdex0smQ/5q1hcq4z9u1AQII9fCKvLLVbGakVu4Q91
RRu52ozr3/hq3OVffOZxQ9+Sz15AVp5Khn2wnR1iT2Uc0+tpHeDJGXpeNIRSq86Qp2brl8yxuezh
GNecTPm+QKzkNbcuWkrglXRiaItXd4MQJGzIsbdFOB+LT33qTiOFwJe/6TJWfDE2dfW2l9sfaDjC
JfRyHyY9BfY881OHN16xsCMD3LurLmV6rqtFRsnvHlbqQrKXg39kiVKxjVZmadwSytHeY5JT0qvr
koKAxw363i8hZG7NvT6eIJKIXRfAujiP6kn1MH9qql/w88tEOvq09xjaXc8COmdA5B7iTN70Zjag
qsolSmYbIuYJClzreksnm7dJBWK07lyAaVIvRw6uLYvVqRZSHfuv5e5JPGLaJ22CBw7hemBcglre
J1ESnNl4pKNgcN7KOq9VTNdRNaCIWBwO1Y2PwLE9OdfabbGHam2/8OKDFiRdeFXCtGIiKWA0dyFm
qu1umQODkULAmps6urNVwRAh5W+vnQcinaprPQ+1lUd6Rkgt1S0n9261jUCFEQtgPBT9JLb9RWvW
lnocg5tij0QutE6h2a0MB5A01LCN1li/5MHce4OVXH4yyZftjntL2cSfyA2Zkj+f6dRsIn35IQYp
e5nmkRrTpnrciNBWI/TefzgSVJ/IftPPdBBNtzUyWsgPJPgToAiSRKroft+G40mYPyIqElttcw9S
/i3E+JxK8vPUXmXVUq72NMX0idv8axK0xLBMXIJUWDsg3c2lYDzTu+5YE3ky5BvGpNm4HGbjyRta
axxIPiVdIZaWeUjX6AkKG7Rukpc52aQY9YvYtw5GW7XZEDbu7aFcuH6kEvKb1ZnQB1+3ISqM1sOQ
Je72g8eMA1GhDyn7RELWft3zau42X3m1C+uq0lF2MwLqmzOhJRoJNsga6zBMTKN96CC5hIUkUGTj
fOmIDkdDWPCRGnJODNq4quoxYWCeQCBp7RFuxuEhfqVBtWBTIz2MQtEBRwVLadko5rbGmvqyt1PM
B/Ut3zRlTFe/4oVRs9gwgKPB6As/yHddeQDAiW8WWmLeI/gyPQvgoSOvB9XxoZpNbVwLEj7KZcMB
DB3ChbZty04uKgM39EAvKxi9rM2y+tllEtjEF2cOc3gNZL0D66e9Kilmi6danJKUnlVisAJJveWI
XQGSiPA7BGHy8NaoCB80bdyXgzxsyLyeuA4fwKyK3Z5nGbcSJrj3chBV7EeQjk1H5RhckiUj98Gs
23bQffu4kyMTz8VSviHu4zpQtTEvGe1f1XtOgWKbhjf7Tu9LKX3BLoS7QoXAtKONBiaYWPxMeMil
V9Pwj8dssyaT1PRMjjOnkyzOzVsh26URjLxPDOL5P3PivHZrl7ftfztfqRel/jvL9yi+sgAUbKSF
Ydfw1AiBCOQZ6pdGg0pY9tLX+dONsjuNXJ2rs2IXC4X7KAXCRPLBGWIa2uAOqxSgi7fNPs2LSdjm
RC9LS9U6S8cNdiaemgin7nu7K0S7EYwZJ/a2QSvuxfw1SAD774x5eo+kZ9th3FZmoeluj50Glp9Y
XH49sMf8xbCf895NY+QJWZ3DBHF49zzXKuEp2HsfD+zV3bk2nyY53eJtgRPilBwkkka/OlfUjdLu
hkE3MLrL65ZH5y05auZSw0uEBxhJK4peH10BhPiDszr45uPJr/hOoKsvrtmDby6qi2W6ycVLo5ez
QaYw+DUKkvnlw9Jsg208LPZqdtLMMes3mYSy+WFVf2BBDEvig/MQeUM861srUEr0ptXthniXWIh8
73HG8cJYZ8HLXuAK+cQq8AggcpKT27uMUvcgzAD9uHImnS1UDdfIKnkmm+FCeiqNcTVjxCad+zEN
MPtIhMfJf/I1UT0MOwAIPogVjYvaEm2agZ3UU5oRzOZrwGc2Q41PToelWUwiMs2m9RyCRZX1YlGL
L2rcGLp3nhdwcbDrpXTVhYiPgTDn5PIrmuZ6cG88IF7b7/YDsQV0sZ0QKEnvm9pFsafN+JdBXPl3
31ufkq35dZlnLMET9qwIr4G9Zbvyue27DaJ0XZpfqV8stKw1nWoFri8Bt8rPnJTjLghW2fUcG4NF
DlpSRqT6EVv9+tWArjG6JG9gDJRPYIXWH7nM6AX3WDyMnM3FkNYFnORdtPM/MduAir2WjzR/ZDhL
cSxh+KUmPBCptpNBhI5qiYjQBNSvfprXRbOyspmP8pKFkYJ+a969juHhmRb0Ru9Xf9dBNNn3Ss4C
YqqAK/ih6w822jKUcK805R+QaRh5r20A6CoJ90Y7s1zQXEtpz+6RVkC1XFE8qwaZKMmhzAW1xazY
Wl+8cTbWJa4a6OhpDhc3LlTUS3qvhHhI66p+f0AX82hv2nVAPzyE1LuZ2z15P1MB2mUKdhZzIusl
ktJNj5uF9BimpsovFTIvd2X+gqfyOGbYAtPtOzvw7H1UonRtzj/1uHofxRmjo7ubPXD6MnLD2Q8f
h1yAMxBnCNsKmudNGdx/2h8gCA59QjzJlUXaxHmgPfT1UDSAxPaFV1Q6CuytMaQ5lCJ13yqDtRFW
37d8QQTAh7aZojv4O/M1Gy56vXUr9a5CqX35WMhN4nVbTbtvuj+7sCrKs1f+DiYwHbpw8E8z31YT
vqAmqRp4LIXv8i6Y0nNwdEr+CDyvA8nF7iuy8fD/WpBI942qdXBVrjNP+esr7x4byn0cNi/GOvvd
Wa28nJHcLeqJT2cRY7bAKCiBACK+3mUo/29aHgf+eV8Oybcp8pAtf9lYJPji6i1DlTXiirLyyBW2
Y6paUWI3Gn/lqLxAvJgneunnx44hohqEZzyPDafwQHeksUrp3qBSJB7jgHRubgiiGcM1eILwlyYg
2B30LTeOytlmpOw+LcAkr3Ud7bhkU+IxXjSQp/H0bHcBtD1g4kqnCNv6XMSjvdQYOKr2XxJIjH5w
tV+zSMk+k7lEVkYBFyocKnQRdpZYkdRmeBx5+jL1D/z6Rr8/T4bXeHUMAVFMewoRxoYq8ehXZSuC
DtG7knqqVKjuPbzlJI6setOP8HUdV5JLuaW2gvwUeHPbzvnl71MC5DlY/LdY3eUNBu4ZRNGXmtDQ
KfdVKAeRoGETkrR9MqQNPdtHnTEvXK0619omoMKN7oWdSU9gL4F6fO2FhFpzqPGqM0yBlitxdCBC
LiWyDJWCVK/IE/43jv0Qlpwqcq7i+3NHIh2kYw4uXCKzRvyKkjNycwiuMTFG+8feA1wg31e5DTTE
EREjsgqrXIz3FO4zf6ZwvfVDPXEM5v6gIjFq9mgC+V73nrV8ACalQRBjx+hrhSxJUpSpLQWR0H3R
5Zem4fAaAYO+ShV4Hj8IiT7Auo/5akMYVcEz5CEghXyAddoHthC2BRVSt84aXEkpNa6arddxUwWg
A4GfFmLPyVl1mG99UCt6mV6A1cEr2LgY0BrIBE9xTnPhR0nbXGVcfePtqzcoAP214ZY77O5OCbaq
6MlSNXs5PTQzKdoiupbsHyUSGqvoHZxx97mPgmcY4LMaQLACb0sBUbUJbyg4dMoB/iub0PDCYdVz
GMmemfk9IBrsSe7rx6D0f1WXnR3mcgTP3sWgAhJDwg+otym4ozy3JhN6sJOqTIdRcPDJisnTptBk
zQwe8o+FNXaG67JV+7ZTls8NGx1xsyJltDE4DAKnmP0LeilL5VjDIEIumPUAPDnUYeCoqWMrl5Id
gali0Jjb7GvdbH5yDOpeooh538h+xUtQD9IqBJsUnc6tK/MvkL/q49FhkchbwfJ4bd7HCTcNsrJB
pyERwEX13pPXEhbEFTmajGRo30rYuhIbSV+hTQjsngsY8iGtNaaB7jrwjDOdAlwAk4UGFM8rfkuw
EXyPXKOtTjKY7pMTxwDxQejwS9g1v5rxmEE46+HaQAkxIrySbJgNZfy6MNRQNTq2dOhGDOloc7kT
bjPx0bw+YE1o/4ZxusJOlOSmJAHM/H/UcITygAhQuhGM/Shl9S63JjcYGE2fnazjtCXS1pPcfZFk
OLYVokHI9suwzzkqx6CIs2+xRPv625uU1GTTQB54QPllxLPxso+AqQH7bJufgnUeF11mZsEYiKmV
/2WBmt1/gIZZfYAn6JrbjIyUoPDzhFwubwwgpwzhOAcz6bLJUW5xvd4pm26t2AnwpGemBvbKzDhl
gUNyIEWdOA05G5pG1TVzZJuZYgpidRxdbxL9WM52+BYMcKAo81ryXxggip9mq1tQAHImnt4bXSgD
nXBmgCvFepTVRdtKdppMTjDPIMpcP2/dv2cCCeNS/WbDRxs4gTmj4ElH1FK7ouP1mObz2ciQRGo+
/fI1DVh2gqORaVsDH+2RW7Pv5NQRpKTiT1i+eu0548V4WgegSNTUR1ufxZFCPJ1HqEOF01fk7gGt
7uX7ZJj553jznnutonMwlaViAmUro809D/uVEj52TBqf38+4Lev0LdDgCdKxjrri6FoN0XdeYLcQ
fh8VoYC9ZupusPyWF61bYHMuaQ1HnXCtgbkBI064lmWkmiZshO37Y2a49bQkx4goti6V2QVl8en4
BQyUC49nCalGTVoThL1QJHw74NS1UrbpDUkNwO2zG5KkV74FvwlEG23gs0M9wwdnzGSK5/clJReC
dFldFHyWnf2dYXOFY+A/VDwQ3OegvJzaoM4M0tUe4qBp5+YBxnsq4SJxxdsrmdNn7DOyupc6iR43
/Sg+DbV9GYBn22+Mk4EadwarIcHzLoHqQU7F7bdWCUioJTcGbdKuyPuF0EFyJv8LtFIP0hPOTCjX
T+GmLR9LJirWtjBPLtPFcURaibakI9ja7zEzPOnzyXvkHqIPk2W+vo1FpE8NIiMqPn0yWaa+45o7
bL0XMVmLB95d6y6uOuHe9sIKH5FGt4I/x1/uuG9TYQCvGfMLlK/Wi4+aTjuAYPLv2TuHKTDy4g0S
R6tq+uEgW+J8TJcUNKQ/cBxoW0AD3BaMsRI447ZUP1aeJzqMmFEI74URFG/+6/7eRtU4pkwSzDx7
C0J0DdRO/+RfLANh72pmFyGDhrjtbCdmslTd7zHpU6fjuCh8jbHd1786ugD40QkZS2nqacEFkodx
+K5C8+vfOMYLSacQI9hc8hVPIk/IhLYKIMnX3kPg9sGteoTFiKkWwM9XS7QEalYBYn6be2mSP2CZ
pUMDc2CkbKhq27LId0veLUvf2+oDWYnBchRO72CZ4SSXPrZzPZq+uWfCwyrEDGPbnOTbVIy4ZQCe
1lbTYW0GdsBi4gJrtcPf9SLleanbxxkSNx5aixwyUCEW1rT8KwG8rWGweRA7JUyASIRWzejUPhau
fLpkA3YPzuKTVvTeHfPC4erOiBYFwogMlYuWvphh9GDNdyvRdEfbWI2ErhdxZP9HozFAZ+obsCpk
tt7SDd2BV0NwzrA3DOHVw46LuB8QDEE119VYR0L+w33Oc1dVOg+tlNqLcOCxsX3oH/Su8FEyCEfO
tzNytOGIlsj8wXquugMNvfQ4TF11lX0PwFY6khJ387xE8BlFyRi5i3mqGioibH/AsxQMzcoq/ICA
USo6jO91rIHDK3fPtRXbB4Nk0HAQBSYOSGNooJ5rQMdA1H0No/RbHLQcCci4nMRtmsjmDbzIDhqC
f19XC0GGYRqG37s3snAXpFffQLZ+W/p5++Np/WokXYTDH8NH53P6JE8SzyAvry0+1MfQbR758pI2
2VfQx5FVYQrU+hUezpBREcLcSksjNh7kMNrnXdweT2Ek3U2isUyHQD13zEhM8ambaUmdRwWuzYbm
3L9RuLyLEiMQ90tU25FggRKwjA5nnLs1cQ84aGDJD9nGqTu9pdKu5rfh0y1hv5gXMcxsnxUyOdwu
r+DM9h9a3YYLOY7NBXrJ8PjA9e3qyNI114a/Ad8wfWS/aKdhr7YZN9vI+qs/R4WX2X5lHVM+UW1f
qvek19vjS7aeXjSfl4LQqldj07W5t4x++e4gDKD2TtjOqahvlrNh4j9UiOWZHV8EO84z07gN4eJU
MCopEgVeAIZKkkYf8r7Gh7LTMYBRhza9PR7bXl4dJGBpUOZ5KswQg0OzZkzqSONfz5hzk8Fsq52H
5qrLNCn623EJKfd65/CMEmH4srgdJeY+N5tdxxsWgNDVWXQxzaEXT7ASX3dgzPvrK0/0tYFi3p8Q
YmefFpuIQNcexRxoW/1yqSYgQ451nOmxe+aetnLPHUFrcEPCexLRg2rtv00Z6zpKOxwVdlN5B2RY
IlExX9reEs7N+acua/4kQK6BTwgC6U4HvQDVVFNqcDjb0bnaFMCik9gjfVTm7xdvAg/m7xxpIt04
g7UHksID6NMPUlGac/5KGeScbAdDL5d7p2l8nbFj460OTEd/dKqnQxlhiXS5SxfyTdwmpGTC3+Yh
wiB6gb5EPNqF1Iuqpjf3hvck7TzL8vVH8o//SE89/+FM3lGKLdCxJAWDwsl3ToZqUl9TavakyMed
jPsvzNWaQy9lEALOKf3wdLRf7FQsf4pzYdUd5VUTJjSy6NA4o5fV9sD+vhMzUEwhe4rUS9W31NAT
yUDrHhNr5us0/jec/lA65ojUF1SazePbCSv/rIwKf33Ifc/jexDlHzL8Aoo8UkJa0NMHcizG/XB4
QRYaToQr2iOOp44pfmgMQCns1tpl92H98vP0BSvUM58C006ILAj5hvpcQPGyvT/qWXNVYHwtkpwf
tUFZ+kexKm9EgwrYOc+au1rgtg7deXBVm/kIB2YdoiS2dRgUPgHVG/PC+I7Svz68Lim3qucGRhyT
OLo6r8rurhx9Aa7j9I2PEilU4irY5xBdkkz6a4jy0U5y9PwnR9x1PNOs12QM5gQtlWqIVD63rZZH
gA5zEN+kubVtMtUkje86WIQrUn1n9JT5S7OyLidVrbU1vUkihQrRSK9B8NJEc6xbxpDdrGgACAUQ
Ti7MQpFZcoH5BS5XiBX9CJcYlKPoNvPLCVbDE8AwjmWfrJUbGfg7lwoa4Dfh1BQN98Q+gjFaZF9K
GfpCRWaQdu5q4YYaFM/fNlbDZ4bevhw5XeKMeZLEP2mprdHAoUKv/UiM+vgO+WdTM6fMtrhJk48V
svfXJ0Pp86ivAUPn77c7ExYha0zOBCG5u4gj+dl/HEZbZTuvSADveqIcFY/supYls4ZonmS+iH3F
YR2qpVvpW0iz8Hzj3zMkOk63AIpB4mtF1ybUfHLskdHkuhfQfczHN3p63MTrUX7uPt+OdF6EiaBD
bNUojznDZQ/AXJ0TScENibQdnH9JkmpORYIF+gyZ04e2dIaQ4vj+dPEH2hTLxBSSEGFmPDzN58mS
gC0xkngGgDv2hKDOcSgBK9Gm5NbGye0uKBUHUohdUQ5UxtaL0b/5WfS6R2ub5bRS/ZeTSij/jszg
T42kq8tMTQm/X9o7LmLBmrD0nicU4wMQCA58rXrMN4FrvXEXfndHNQoI5pOsV2x0aAE7ylHE13QP
IGZx5AZnCq0HgDFfxwZUKL7zqupIt0YEwH+nEXguCcJXHGRirQtdkgMRB7yT2BeJEyFnObiMoMZ8
m7KmRkG0NpwIHSUcA3Lm3sjzKbvlq1EiJKrqdFJz/K9izr0T922KTrNeLonGIm7AAh6STWJ1q9QA
DCBXoHkKYvtBdJX4bsEmCGoWYyewv+RqPyDW+/BmdJLns/xM6D//xgjf63PozR00Wavg7d2ggWhA
k4fY1B81pGy2M1HdmZV9oNoEpvH9pxA1b0n40BOaNO47mskB6PKZn3cJqXTgEjCu4sbDzjkwCTqd
3YszfA5i3qDhgF7Ls3vwhRlWgmtUc5V7sxmTl0EcODPO6c/jAPqV7bT8BFtpjxLcHUEtu5IGxGFc
rjO/iX1fn5ZL3LCFb6QmdD+jx/Ij9jHZx/GU07kGzTqLelTyOU37410tZzqQH4S/mLFpc1PCLtw8
d9gr23ne5WVnXmYW8RUrKKaChcotU3MDVVktg4OTAEzyuHqb9+Cg0tIVPZs25lNFDn8jekBA6foQ
GmUH+e+ecdgB8Btu4R9tSxPS6e4E8q5fTmFe7zFoTYyoT/IVl+OrQb4WLuFlruhEqDvX7f0wao9H
bVhGfsnoeT48O4QudaAAoFOuxzUz1gldLyfdMVbAlUbO/uXdFDEQT/PKtiniij+dI7tzX+Z5LdNJ
DqAeb7lZPQuCaB8tu1nKO8mGU/j/KjUcwSCsaDy+fGYz3Mkb3c2KVVM2kg56frmt3VSkXZrN1t3F
mnPhO4NvC95WVWOm0RxDEJSl8pSCj+kPuc9KPaC2NGErQ74h1Br0+RUslc6UtoHzi4vkr18vG3UL
vMP+02A4hLBZdLVkPftldBbvOBPCQCSNz0qjm7c77PhIa7G9BDpWEaa3A6S9Al/pEF5l9rDZZsSn
rfAgjt5MjDCixqUwTAqSFRXK7Ot21eeyqFoy5NDNTslbw6vhZDanV4Z7+knixQ7V2KpSIhLVLpDj
sQsT1BxmC9VDH6hUMKB4hDGWfdkzj67mVuo+agLJVWkHFD2vqmNGQld9ZIgjucTcPoWLT8N/ari6
zM1x9AMW61CTjwTpp7adZUVP9cJJeTxE/cIkYCuP6PPcq/0JtaGzvi/XHasiY2eRwsHhTGzoZsHQ
gfMo3FvQL+ZaUrdM1INLSnmcv4phQE+Cq9XbO6ShE3bI3vKcnhWfrTn1u2d4owiCcJoobId6ib8O
USNS9fjHIACWCiNfw0esWJ4iCTfIZ3flGuLyFNJ0kZhsGX86qRIzS0baQnRnXH9RHmWczY70eCNz
z6Ie0jehgf51+/+pyRvY82lHYxNlFn++CyHniPJt5IDL1SFFdpZb7YhwM1MkkEb3vUFrqm8IGX4L
LI7bECB10BxsJpxCeJV+MEAGQ/q3aqmUgkP1GZqKoA1241kBJOLSzeejbFUgxIdaFVVatNZdK89c
2QGBeuMzDRM6C3MkxqAAhlVMcqzq9nkoeVPxWyO15OVie6dE79Bq6RLY1s9z/ErVYdWcrMxqXD0T
mhaUvOh7DsYyEvWBPJJSUA1jEA6wv17jkHpwOt1C1dZkkBQt8mIavCiSlQGgx0lmcGGwe3iG2XHt
vGDv3SnMxAt+6nEF+y7Lc1loJ7KJzuhJzzjWh9uEZ/+CFqtGSTBr2II2inEbXkd7/fVCUTPsvhHI
WGrdaGMfk2Z8UvGf02DEeICZVSSlo3mjtFwqGXy0f7pPLwTA5P8CdcDezoTQpzdglNdWEKVGxzQv
aQ0hXnri4Xe0Wz+iPNH5E5I+0jGZap8vrc3/99MoK2XAl20QPKOg3mVWvi85n/u7r8MeHfMAFj7r
1/0Ngs/rWhM437DSAU5wb+f4Tz9bmrwmS/TN3wnZh4T8a+eNFJ4x6V93rN8R5dX3acHc+Sp6Qdfb
cg4UaaywrVNnX0aDlQMhpqg490hm8TBoQFngbuv5ItdsITyf2QhxDFRb2xnMkiy93qOVYcAw/kWv
opwE73FXAx9OCgIuZMWPLWKkfQBQKDBYPUse5qqtXGRJ8cZhOanSQq4LY20aaI0heKKvQ/oNgttq
J2Tamp4GQWARexxOazr0odY8Fbjywo2ja4yXtu0w2ez+wKpX7iK2OcNS1ke3RrcLHC5q6TthYSRg
p73T5XkJeOl56V/Swp05cjaLXCW2aSRDG1fyTF9xzf5qXYyYF6+Q7ViX9bFPiAtui581l2CbGisE
M1GuDxRl6ryuwp+gqW0g6C4Pl+mtneq85mxzWui0lWn4VUN5irynNLBIEll8YX1IlXCMhQRS2ybp
cNhzI5b5c3aXpPK5ScVpUBPk9NfpOvKDZtHDzEkjZHHMXYJSma4nNXR5prLeeI9BrmYKkzeQJccj
f0WQI2bdJUYa1KZzxxCrAHKjsgBNZfIzKT9DOlsPzXE4RtZI313LZAOb1wcJ0w1j8E9eS48kI/yh
jk9SQgm+X5flSqyiZ/4leZiJcyAj/RLDsmeFXD5hcAg2lilrXxoSqh/e7vAbyxQl+uHiNsuVnGG+
h1dLQZ/8h6mGypdP3H0G12oqGLtz5284Nc0gFtUbcdqGYrWyozSuqsJjqaojzVnSacfxl4un+PGy
URkZDHv8PWQRYAiwlNY6r6jnDJ2pOZESOzZiEMkwEses+qvLS2Pmm0eokX0+Kx9VSta352cFVEwD
NnCuktbAcAbBiXQkR1QG9e+ZgHU38r9deSAe6KBKsAoXwh5lFbln1H4w7XMR014DrmDrI58XhuuG
OKBtZ4FeFUAvlzUK6+TCtd8QxMkr2hS1T8rrlucW7vkXmVUAuNmzCN1/WRa55QExylgk8gDeGF9/
SKx8xRFs8ds0ffaU69pRiftUbZYeluDNObIYaFkq83fW3mzJdCWZYn4xi3POoeHOrlpAdKjXyC2s
Fr2w6gBW4mWP0+IhQjR3if55T3V2+YYLm1b+S4SFob7D4dTkFEdBvs3P8NnzcIXTGjXhOBPmOsRN
6UKTMg9DoXV3w2G4FdD2TUZLCLMfoCzkjQo61oE5pZ8pxQ+PA23y3NpYFVjwBErcv1kJexeRdRIT
p3qfTHF/xGJxoUEupH7GJmz0hLaW8tmZ9zPqP/g2THOswDQCWthWtfhGtLFWcBubckNIQaKwNR0Z
di5kWF2mZTQIrCC+0Tnh/iJ1a6af92wA/Bme/MJWGgFkS5qw4KZnRcC5atxqU4ha6wmF75KhWbSe
2tle8N0umb64PgWUT/GYRKIiUYBdsxpb2/DMUXgmrhIEZT37aNLaKMJetfkX7OsC3lF+eapn4KFn
Qsp9/TWoI/TaOtwXRURrVs8ZikfXixYuby7dqzcNhCwYTaIDBxy4JJ+ChpctcchgvL2IqUa8N1Cq
nFccXLT1FBtHBkmYAQ53I4T4O5wtJRsMABKF5IFVihhpV/siy73819oXn5/BdID3d/o9EeZG2XAo
Y9udfqc++lVdd++fVGuXtwDTrM1gsFaK0ojShnt/VSYYmLMpoVEmMkFSVNKoOIRySjRAQ3lqyy+o
zc7DofjW1U3i+bTvqgopFYR7qF0bxRFWZE2MOAUh8wDH3/knoreRX56X+UNX/UpqRYhKRpqYs2l0
SosI0g3CohaS948ZqT9AFiXAj4VTOu1VBynvh2JorW52/Kjz52XIzdIxVp2p57CAIFHuM+wuP4tW
UOm8AqRt9PbL/TqnLXPv0dngiOqMlAX3Qe6ehmiuS9oLpbPRD5CRGTkRLY2E7zz2PGhqkK3ct5U6
164H6UoeLIxs/t53YX+YLjq6RtepMqpMdeG47UT2ciuSBWSrYJPrw2fZzM37TLtSjgUko0pWVasn
PCohO8mIPvUBErMm2H7LiLx86cME0M5ObBOoIXKn7JNmSQp86bQBCEQH5YUv+9P8b6pnlrqAupZ8
Q1nrPKodBg57U4yNDnc3aWf2UoHrYCskZpQGnex+3BiNWU//VXj69rZbwPYOfn4vJXUEAHW31x6Z
5UFUlhviMUbYz6gaxovKGCI1az2l/rqppbngFHcBJziN70MBz97J61L8mVnqLETrFxZ8fcGPgA27
wfF1nd49H3u8hajoJe/QzXDHXi3tUP9tXFC3ZWMAPstEq8vMfXiDm3v7sHeb0Y2fNFn3NM+9seTv
ep6hPGhHq1kvTib70UAqXJ+kxXvyjwW5cvglhPI/0BN/WEFChdSnEu+YDXXZluRvLFqFPjNmprLM
NkRg2m9QTcqUuMF0z59yHICitMvnwnUJnG181xzToRosVJf7YUp/rr3Z3fAgwLgg7RUTeOZP9cZQ
42uBfjDFtxr2jFgj5IrxnEhCzDYC1viJJjQhQbrV/5RkuKZdsRcGPAKXp8F6kpEQmnAx1N6kv8bU
RhpUzSavDOkIB6Xijqznb0HMVk+mkbhgm2aclGZNlawhazY/tdfI2CXeRBvvX9hEeQkx3Ktq0cdc
L3M3FQ+jI2bNQ9fQqJTTALBCZP0O12QOmBsT7H+ke4Dr9fx8LHenP7gBwlXbco3aAHIYuEnP/EeD
tWsb1zMwhIgW8Z5TALdu61FVRhT+TVoBA47gweaE2novvaNYNXd5U8Xv9Zyexn2agSvgRDQvmeto
fVNFBfiN2/yzvpLUIo8UfNyE+TxYun8ujfiWx1mUQelgVA+Dp5/zmzSN3BxTwezY6FTB0mKaZwKs
2mWzFcpcvIJRT0wk9uHZLB1vrM0d00oubACaw5vat5De94M/1mjG1wjedPeFqQW8+dyKZVHupCF6
4TlSfchaAZUukPwWKCushccUu0gorV5C3fjvFBsVy+zwRoink9qEbz/8YqOmMIYQV29ECe90MArD
JMaiUBwyl/QEjbOJcQBgVAJsBCxMP7AKmUkCgAf0NZemx8VNmW8hHaxMQ7xM0wipyuL01QQvsJUI
G9x0WBjpo0sA6g1b9KqPIeDukom/Iq2mhWosSDipaiDNBn9E5+LZC6xc7vkB+XjCsooaNba9QZNr
vCopCu3iFlIYsvA45JDazMsu9TEifKCUR5oFEzX/Vc1PVuAI+2YX2GQWZAatuXu4kiXTu/AOPNgB
otmhg6qmE86fzyT5Jd2DUVZbVmsGLEtBLeILslSpq5XLT1g9lpA5f4qIUTQ9VUC0jYW1DsxHWyja
fPuIjoonLZLqh9+7nKCGmE72fpegBHRCjrfZU25a7sO329WXQ4lr52FjSAuzSNBY4besx3I4YJ4M
XopcE1ANzcrEULTfLDu4Y8J1NTTDO9/XpvNTAkQ4LPirOjvejUmTzGgCIle/H6/vyBqLhPTLGalY
/BuLAFHfPxpBuqc3HQ7UhUdX3YDvLtnb16Qzk5lQgDsg2Dt3h5rmL64xEVybxuKMDVB9Cwk7WhEw
xqes6w71urHP9Eu0/jRxFxb1Is8tt5ijd/NmaFFlnZVnYuLHNzvots7MNYLuMYalXn4RdU81Ar4G
15z8wAK5/mt/ipZMB9YQlfaUrRbgqLuhydM6IYf0TlqQzmiruJU5O8/wiU7OpZqPh3no7KjDSLGM
83f9zGtRsC09RS0N2r1QQdwyqC/xHwdBANGF3JdgHOSiaJu67alpVkgwD1qLMONH5TuD6KXYVGbl
6rbNfnfLEHtyuEvMrzmBG5yvrV5ejMK9gK0NMiUix4qh1RnajkJhrE5V16CbS86RwMvlVadIki3Q
RmlNHtOCjbXOVzws9PBbbST+DVkLL0oCog63nMcyhkp2/2BqAWQ/yDsqtlpY4tw973yTvn/VGUJa
w+pTiYwYu79oUEqXX5AEP7MR8Foxx7qAGTHETTlnDxa0k0ZmndzNwl7p0eFPWb1r8NERkb41/WMS
U9WyhEF9mIAf0HKnGxu/59+gvOia0pGT5I6O4oqRIXQXwbemSPjvz/UORVksPLdNxVxDMnUVKklf
S4+Jajs/H1zJw+g71QIYGgW2p7v6QgeFYpYgTNKV/m0rnGQbE75oVSYulaIRmCGVpTNBw3aOvKRg
rxNdndv1ru8AUIVOpYw08qNVFVe5gsDAxXTBRd8MTJfyOLBXS78ymKnW084No81upGLgtTH3cs+r
HYMad0u/cAQqa/9IJjUiHfIyAO+RyZmGZgg3uWdc/dunDA8GY0URLoGo77ssM1CU2rxhTzs9+UnL
Ju47oJq0RNm0jbzLOaiNkMRczHNqjjxVbDA2TuJezYug2jRu1bmhTUbkzuaYhsWBXEqWWAfOhbvq
nWjR6/j2DvDALxxJvJZSYAf2IW1GEkThLx2uz1LPOxzHlAMqOP+f8HDBAes3Mh3n0Entos08p2kJ
PcH7mRmzxgR63GCzLPHXVYO5RMfyYUA7g67mhUcJCWuWQT12tjm5xixIU+QUXImhqCz2MigXaK6x
lKV9SUQxZ/3QZ2ZfgbdpbTDnoBJjiWVuOtHsTQSYeiKTkDeL/h+68GAmMoSN3SB2iU7aIU1HrdcJ
KJbmKxMnPaYgH0PZEXscZLvwxrKxpDS9wSh1vP86PEv17RUebQypD7oE/GNMT6lPU0bzjHmoC9Eq
eqLYOTCX7muMvzolB7LXnTmg9vYt4rsCk6zayBZ+yfIEn5AqWMZUEQVrQgrisGvAjtrQPvL/k85F
vO+0dOVBju/249hPXIJEQqfWjG9XJE81lybUmPUgxvXXdii43iXbBneFQrAxKU73dGaqJVdS8jTC
gdyLAuvLR0pHMt3JCJvPBdPatPy68X7nQBzKGchwtqlDbKiyulWhHup968AUwsjyPdtmPL4+BK9b
WcejWht7pP1xxIHWL+skq1/es2hh+BDJycvAlxUMyT4equcRhTd0uE6ceMbXeQGmhEloAW7xYAcl
NjYjlbkofVuD4vRzsGOOxIcJ/ZtjhttfdnSAZYWQlqcFWiB85VrDh13zx9CWV4fsKjGVDcVeIcJS
DaO8ghwcvoYUZFv9IdPB6DJicjmCdLtvd/d/z8ZZne9nS1sbywMc+kojIUv1b+pEW8en/hSyj9ti
LgDNdESJSHh2lu0aAZP8QLa+LRc21+Xmp77V9UhEbj6rPs+Pj6PX1yYuM8nWfom0ZaPgKKzFrwMT
tPGepeUVGhPuQXFWi7aPM3gMHWYQl4QaALIBZDoUaYiePSC99SUO36MIeJzl3nKDrrUCbnjSX+PM
BWz+xF3z8/m8t8nWZZqxCpdvr1ABK3wrrrJwqK5Lp1IEJUfDPv+ukm80p+pyQMy+zC+dbKP6QLLT
Qk4aTD3kT5p+iXrk6wXj55lubeKrVUnOXlZ81qdXAe4ZkmYWjmDbMt1wjPxzQQV7RYBz+Ws3n//S
VIfVoErUIApXJZrDsaYQ2TixtiymUygF+6xsnE5H+K0nJy2GigrWOzz9fSzx90L6twguaHWXU1n3
cBSniF5gUbCsngIMUik43Nj+eX52VNFVCdeFxdT780N0y+nM7Na5YvdVJn6F53D+0JlnA1l7imgp
6TlYqzI/wpWedHuJ+rTZXQd1RwGS4QwRNPiGx3RmMJTckRxatj7GXXWWD3j867VLMlBt1hTFM30y
Sr3Z1P95YdZjIleD1iUvELkMUsZ754wXtBUaGx8OwPHbwvUrUpkvZhhEcSkzf6izMBuE7Kq7uljI
Ma2DC4m4niRGSht/UUGQUP5Dvq4qEB7Kejsu2RfbfCEAi2yReqgGyDqQyIa8NUbWQEB+mLpx9DhC
vqj2EJ7Kn88sQjKXn13eEhZvW2zgvAVBu1ErNkiViD2nxFP75K/dCJl+wxopuMSOkNIwO+LsMfPg
GtvPEKSpzr5PuwXo9EN3T0DzPftvJBuvzm0ttRBmOfgIv6p14I4lmH8OhU4/RQQasiw2wAXdh84h
hOoSO6igBL+zvDPvFbSXI23XnRkir0wIWF5rC+EeBVjvWgiYiBZ5rTBcP8P58R1yGqF4SKbfCo3b
WRO8/fEna9V86pKDnAvYMctxtdqtdCdN5SoqY3JSKQNPPvb2sWJ/raWdywNYyZSR0ingTZqZA3hK
f2WVtnnyERqlESbYucD12UOog2ATSJaEMpVe7WGOCCLBhHmAuZL3LMnouX0Z09mL4hi9ExRNX7OP
852yUsS7hUE5i800MEvnryHs5hoaMAKIv+8X+HmKL5R3OgoLqeEUKwdyrRm71NrO1uJov3UHrjjF
jfpyghtRi/E1KqlMSF3Mg3L9tx3WryeiTMYv/Z9J+HSd6ctIvX4NV4XtrRZ8pDR2NT+tjtJXWJ5y
WlfudFJ9ZplOVal8gf2jUaax/7k0kapl8B8oPlcT1E5qbWqcPu/eeyhS4kWK/J42xxWSyHV89XF+
O2aysILfv1AbnccPfygAM97NpUxR2/F6VFE30QwjUU9R11syEf+ckAv6VpHZoTrRV0UuiqYQ3OlM
yEVg+FnAlF9fdcezYk5HbGrGvIuhg/BoxyoyeB8eCc0QCz14LBNurMlMCh60qx2NLaLwMEMqbuBP
fm8mMudxOu09qE7yUmJ7cPjN/V5D6zPvN2xvcNThmKLngNHqf3bYjDeZ8W7m2c+03EhG/3u+folH
Aig8EMcGr4Xbq3NU07KHVRnZMKVLGSSV3MzfQvBdSd9gIlfiGZUNhafvCyrNO/g6FAuv15Nhj2aU
g0qE4ppxWw4RIah/Xp1kiGxklVzF3Xp30r52KSe5glTXl4El8WW0+BY+jRsBZzU31ZECIRYRbnQd
NdjZ5By7YxcA+XO18uoQhPR94to6IDdquoxdgLryeeL/u3hODiJkIwnbntgEoW++f4pz0M+18g/U
OgBokT5Hs1yPFTyIkcqRprqrTno3RFXcG5NY+kKIU5l2zAz2n/EqnC93cOJ4vW1T+riAzFU1AZO7
bzEKoBPTOko3wuuqHzMSLBUQUgrZ+CZuKcLcqsr2MJQi5iKaTIo+3lHlsc8bDD70YAy+hnV56n/8
pd2WUVd/2EM3PLpjBDtvK1p4okSiB8RmQMsqFaQLr3rlUHpbDFF/cQqAbNuPyV9Ve+6HmfoUco2V
i1KVQYscOmywyc4qhyM5sMnGpWNb9qQblPL5Lxi5+Per7Txz4s3e3O1svAAM+KE4n48Wfx86iGH5
8B+t1RBQcWXD+RXLzv8yDQOOHqlLW65WXDwNcGpkR/qDRcYB4hZROdtg0hWmzMYRstw2i0v5uKum
VIXHuiQjgiDbO9+auZ7MvnHjJQpgpLZRurtJkks/G21MHlVepu7XwpZi7hIIiAZNp5biEA28E+lr
bnnlk4uQILTzFbhMx70CKDrgQliZIhoiSSB7dSWqtosL5V+uUuaA3vxJfkhvM7v69ka4BSMQSIJ6
Z4S9JTqDyybO0HzrA/FDHpEnhhD1rJdlVBxh9KHX7Vnyig5zMWHEEa7uztW/dUKWXfYvd6HZcagm
LQv24dh1M83Ywb60vkNQAhfkjUZwD7xPRznbDggtq4CoeDZbE89IM8fzjOE+0o1YtYQxT+oKdwzO
uAMpuJ23RiBocj4o04e4YaV8Gw3Z9jtHul5jOCvcOFmlhfJbqmadaeaIHXPRnZSepf6i4ZxXZ3sq
lOgBC7gPm24amyqNm3LKzCew9+0hBDE/Vlb/VtEgYmzAjxt+xi11fsVJXGmIJsk4ZixXavJ6r2Cb
rR9DG6CarXnjMBiPlBfbK4u+jZszFcXD0TlaMjeb5BLFd7tZ5WP8saJcmsSZ+s/TSzpsx72/0XQ+
SCFRap4Kf8ad3drD2sW/y65zpGpkeYFLQUublWKI7s2zUUINsjKr2ihp5CuE8oo2dpLDkfHPK6Ey
V1UGZClChCEJbdjoR6ZqTKppCSfcWrIK6IiDurkIch68RaFhqGED9IEXyWOxJanEQW+IES/2Mari
ht3NGuxDgFHzA4MYPx4sb/cqevf/kpkJwavM//TDx3bkLaR3vOEjrMmDM/aPQMg0b7o0m+bZZEI3
DPIXqtzLq3f84rc59O2R7/CvyCHIthK3gffX/4UqnCFh2kl9kNpc0i4IEH3UWdCQG9MdXF/u5/to
jZaz3eEtDPU/Idfuhiq0pfw7v9+2etWqbNwvQ+sv6yuAm6CYbvHWd24e0L7jjDpUIB4FVyKNFlVs
/Go7CGXZYosfyGOSPgOL8sva0zwb6PsQ/lWWSTGtw9+xnbYvM4F2hLYMCx0MU5fYLyOf7/9lJ7oO
DZOhQOJCwQjnnM6YM7EOkRw8mQKXVLBnX9E21YIfcrfmRScn0Aicts+wYMuyL142o3bVQpM6Orle
ku4xPs9LLdctsdCi7av1KV02lE/ysVoXDACN2LjyBjCM5EBj6XVDrDmGSDEruWLGhpahYeLnVj0+
jqHX0uD1pKb4uYWRkbi3VUvBqWhciwwDAO0tWelLhgaRx30lkUrk54wp3D7aGrv1YM2IZpwAWxsu
kHvg8Cl+i4chw1xkqz93hA2MtGhhaVu9ZfczQB06ihdIXmI+9M2CZeALhgeNusjgQvDFGSRyv48j
FAYiSHX2a+eCfpuy04hXVH7CgnCl0cIa34Sh4nyISAOc6E6rtLzcy9bVRLCN4kSBYrfgZukspGzK
YD5QjnD8Oc1XsN+vNvqRoXLf/XfDJazsyW0/HKeke1wFMCTU+OQoCzotfURYp0QZ4ksDbzkoYNaJ
A8uJZCKa418W7tKwZgINv+SvCECv8aRgArU/WM/v+pUlEKsvQeNa54YJWeMrYdfalwsDodA9szHn
XIIUeun7zcx9KwH73StOfG9JE4jiN7eMzyJCrwJX60BX23E41wE9Gyhond92eW3fIm1QHEU+7EC4
EhoKUe6y/1nN6RrbT+NGVPRaHUPcTErsbc7WNlAXxFpQZK6qkh2p7waUOrSjzTlSFtopJD1aysPi
5vV/cyIdUKEJnLWJjdbOlWjLapW4d+COa6UJB0aTMeTF01w4DkYLrOQEw5pWTfbuosnXVMwy9Kt7
JELTmxrl9f7Dd5rm8oG26mY/io7N+l3mpqP6ELzdrtULCkyuYz2+g2EIj6clBXa+EM2aD9vXiAiw
pp0SncQGRTbdzenfaZOa/NP8nGI5W7EHwlQLT0BuyCr8fWfY2tgSF9af2Ldyt/dc9ofbdYdkiSoN
WV+3/2LB2eOAgLHRG5HhjoHLAS3vG7rfXTLHwRhXwDxQpSnlXSCleSbVwFy7QsfI+ZJBGtqDxriR
SRQSle1rIvlGXVscPAJ7QEHltZgK/vVY7ra6MUeVKuD+Mr3zjTnem9Ll+9sxsccbNSF7lnqyviCx
1tdPJiBZ5yAzy0mCoaN18z8sPK3ESfFCoaO4sIQs0mvqOU4xEujL4uY40uTs4uCg4E0ngk/h+TIQ
HF/PXdHJi5OhOFWCGmDtZ1vVb+BhgFecN4zkSkoPuJBgNPdrbUhY60JXMPcQX3DfIAMA99H6a2V5
4LhM+Ywlt7FIV3ms2ctmpfUmmD7dxlujrrJPzWeVVEIuF4soTlW9zDZvInvFnCUuOEhCFnLhti6J
anGTKl/2UcpK1pXoS5HHGDBsllS6ODW0Xgtejsgp1Q/TO7IKhABfaVrCCCdSywUweNYaVbWaHpM3
Bphsv/g0g+RXwtbJA1r+XPxeI55B2YjwXaUV65ayUY+gO3yXh5tTtXLL8m1kiCHrK7p9bBG8IE71
6mBjBSDJSaDZzQzPC05K9wnj1JLFPrwGKq79FZjXkzwnveE7nCPwvULxFMLty2LyZXOb9479vRWg
qtnCZcxMOJncDp01a4B/8Iv8TuCaDKBc2foDoftMYeI8+bi+ICUGkI57J4vLccD21BxLFmQToGX1
I5q+RHhPSVv6fW9IECtXTboB9iOUgGTGs0KEH5kbB6NIRtHmmpQveP3J2W2nWg1N7XgjIID9wAj7
6VwRq26Truh1mRd55r8YezcQ1EGi86orz9sZKIZWIkEh3xyYzZa1C/mTg6NJPGTtVuq8Mq0DzHYM
RdZevt7XAdBCEZ8Md01TrBotv8XST57mAlnFwbFoDkf11QT42HSF9m1KZ3UAyMD7ucFAkrdwqtlU
jF6DQ46tktf0MVlWIG62fEqxukUPus+U1OlTssU1YAyzoD61kP8B/6KZs0nAktBjarE+Dv/q/Jdz
gve7Qu+VIhp4D+LTPjoJoEBXPuvbNscJk7nMu2TM8L5F8Y1tMa7GDPTxK86vC04WVMVo8uv1kSxb
+pxMJ/Z45Eiv8TOUIFcmkloIHq6W87zV8tIP3du3ra+PuHaBLj3E+2DmFYqzzFhsHAPnjWb5Yo0A
7MhF6gedT1XVkJOqyTS/f2vltgru6RxjnbsxUEUHsm/qOU8YqNqlP79wnWzUgbNhXgCcUwCJiebI
yHyB6QAzLsgVGVQLkGaH7C1BQg7y7Z0j+Ywdty92O3pNQFGXUuf7g8+PwpFBP7iP3OX/hLDfDWCV
jWVcbV9BI+NzuQZrid/1jmTIQeIymSRkbx34RW1BRJ4SoMJgbCWqci3MZXBMqgx5iih33uHl2zQb
gX8HxECaII/Hpd3+i6Tzf5nOhwi7aN/ViKNnDRWv202kL8jzoPRlZ8PJnHFwK3alpxCw+r07Jw1W
BQVWN7S/LUWR2/GQ6OLS0fgT2UhvOv/umemJitERqtXsVfVOiODAP8aZeJEbQMF9tbHbjsSWQNPZ
00rmuswzmqCx1b87XXZHoTL9rubBoYN7IlXbuWdcq1glx7Sk4v9XdtFNxR6ofze5D7YA0bk28kll
BxvEyq6cMD3hwNaL/w+y8Pb/6hAr3AXmfJeXhVqdnIbqQahL0/+CAw6VhGxldxzb/3S83MwhqGpW
do/3XG0fKSrugNqGujFfuhbJT+VUPhPjaKECo2Kmwn3bRlqN8Pfob5TSBDWx9rIjb7rjaVVjoxtC
9Hi1aIwqYECYVUZ1Q+T/Tah/hAqpDQkt3Yk3/gxTXC/xw9W5+2W+o8wfqaLbXN+sI55xsTCrqCmK
OgJOzcPR8eXwUDrsv2Y+tTF7fqBrmLe+xk9rMUrN+NmoSqwrCwpuSt76+pgD2xy6CN9GbMNAk26b
3I2KIoUqcuijcI4geOdy2X6MbkrtXvtzr39ZNdI6a51we5YRpSrvtBt9p7Yop7FANHuSzVp2w4Td
fmK5LUHocJV4/6S6SXLeBi5/V7lFDMyqIeXAEbVAsH7n2RkStIVKJsArWX2nGf5moZ30HifcSfSo
JhQzL18cFtNF92aulHQS6fiZtVBr5LVwNJdDXMF4AGTQqpaV1GTxXlSj/WPvDArhfVkHZAExX9xn
6ptPPIInwK9XJ+RYw0UcP1cJH26uvTgNUt/8HFtTiuuU3Fhn5vq4hAB51O3UpmuGUXmOH6Gl212t
lXQXrSn6uREgV48dUgz5KDBixDE60/vOhD5pMTL+475dQolFD/jrKQwBYq7XdcNTFTA7xmx1U4RB
BPfTDVo1OEv/3uXusClmzS25FcnyflB99+7spWOnfOOy/B3OLV5llO3kDRpkI12nBDxAEhY4Vn+H
HVxdAdQztYucrMCbWSsk3zfcsv6gh85gcnTlupuZ/O9Gyd/+EYEDFEft2xql6cGj3D8re1DUc6dU
jDAwJULV/L7oEWQe2Pv/eFl3HHFAlMsg2uTKbcBLmYtSm8nLZjTgN7iKOmCcIOFhLaU25S6fwtLb
5niG4uo0magrLIrEhk9FijhVqlR+wUAHZzbdmXtBxPvlrP2yIEfFFZ8H1eHHc5MgVmWF8qR7tpF8
JbIz39ECKPcLur1bWxywiqeUAWjfE8PGN+NYdEiE76Eqr7B5NKMeC6ViiA9yK1oImUFFdpU+9ZyM
tJ4L5/jXBv6+OtohlCq2fcynsKxqRP66TifhIns86MJCK4RQSUu0nqY0dxJTuA++0otgBo6djJ6L
3dcqpjWnf1o3/0IkE01H9BcC74bPpB+K9Dnw3UqplVPvIgQTskxTlVa3dizr+9+NxomvyCAvKoRB
iezb2VCned7m9/j9ILQsq835JefdaONLHmH9g4Uef7cADCzBIAbo5ffJP8V4K8bZYdds3c//I4ao
ZJNari0n+Kl+2NvK7v8yrML1CYGWM0LfqO63UspwfaZe/2UflESYYVvfa5BLR534c0jMX3RS0uP9
zKL0xUZExJSanNt5gNwZk4z+pbukAzMitRUfelYxn55fdo/EcPHIbgHdiMFrzXxIpXxJgcDsZJZy
UOChZBD9kkMWCNJli26kxcKMNlx/4mF7T8tVoo6EAuNgKtoAZHA3Ldis49tkr0asH69kXE/thWfH
I9pQ1NQejRdpyCGRDC7SSwNR/EDZe23GcgEi1aGEJ1NSt1wgBbMUED+EPavuLCkcKDnhpTOaLI5K
Ux1dRrHRr5li4TxUjtzZVFiYcSX4zygfCiQfAqEN/RrP1rOXEmxcr5s4jPDCxyNBFz4/YkYQSBrU
8O5KpJ0bMmDY4hymazr6jdJl3e3RDhef9M0wmd2lM0xYg3ciUJrvUZETo1Cxlw4oMZC0C1t/qL5B
eVB6LcCWCUO3ggZzklrRYvDMuvuMYM39p/J+EQ4C0R+S/BYDgBvnMU9ivqNgQFRcIw5fZ/PbdLLK
KuTvdjydNCXFE3iTe/ekJspy1aDRXKBhtpLQcgOOisPHIe2V8ZqsEjluSdcqt8isqoJ+XvMTshsr
zoKqFTZ1Szkw+1BMgvGbbcurgBAQ+cM/x5F/E2ZYigZb7xoTRw5X92hcwb1fBijqngyMG0ajY5r+
RSK70aMV3VdtxLkA27SZB3nsQMsDw0EeShK3F0/5BrmHOnHiPqWvo+IM4XvNKDXLdsaCwMvCOIvr
JsqhVhcC5mxLnNFHQDj5P5wShtTeH03aHd7YX3cklA9fZLkZf6v/m30hoTTDpgJrcFmhWNvhn1KB
pgFWrJbNiRiQNCQsDu2gTaT0Xz7KBn2a1e8PgCI1Ml7JhfFxmLR4D3vPtCMqhwhOnSnEhqWyyqEO
Xnifq0eyqibXA4jth1p2k6tUzrTrJBvcwSfDWAUS2Pq93l7O/HR2YNRMBY63s+zGQRShuxm3O1aZ
aQifdm6TmBIJh+i9158PDYN6QBJlis6uhNg2Lb7PFDOjFKgLFbNqwMWSvr8UaQnSMSpKSG6VBTLC
PZNOjDsbP7lGWMmgOEUBSpzTuOhRUhlZrmuUWRJO8gMvkuOHWW5QmCWTThMcXGKj1j5kBMRUNx/k
BPudPx3UoIP4DulvXtz1f92DfUqUCCvyn2vj4vcoHpu7lb+MqXfmdoPUozCHKDsN+VI1IPDLrMCC
I3fOc8WWkvBdD0dvQLTxuarTqUBQDy2oMXex2SebdHm3zdl1YnmGm0n5hsH+ByO/hC0N+nNSCmGf
G3WXU1zlDebUTdpgpVCQcZd52lxLis5ql2QCqWEdvlFWaf0WSnqp9pps5YztZ1bBDVJ+rl7QN6OW
ndRo8MwT5X0pNz/oba+VjesQ/5Erj+1WWz92SJvgG9clclF26OkfrQQ4lrfysMhGFwKIRCeiG3YX
4egMMhQZ9HD1aSin1HK5+Q2aZ2hbUci2d5/5xehRy9nQZfFui31FdITu8Y6zv0BLLAz2Nn3A/C/F
kGDY6rEkn8kVCicycNpWkOxLf7FgIWLfgoUxcD1GLUD0ekeb/OhBZgTnFsQf90OQvcbMoDyzXeT0
OSNJ/KB7zKGK0yDinYYf43sA4m7e+F6/GaYVg+i5jZRmm5ZbHR1nYQkxjoaSZVW0SC1ckrCUkmPB
h/VmwV6NVmfe6VX6q+FC+ujfXaZQ8T14W+siVPcwGpp6blRsROKRA3wHaR9Aa/+452MC5WyusZv/
ITdHmthir9PxZCirvgNqxDLL6+hUh7gYblzxaou2Pn9h2RHv42iReTRykzXS4UtB5iWRAniWbnr8
RWFoLZ44TOne5BMamWXIKuA4TmPEddqScPQJrjhmYWU30Cfhzz7837u8ASgN1762xkDmKHLT5oha
JCy1Kzv2aVQKXSib6C/CgSsiC0XZV1BC203uMjmLO2nSEu9q/P1CXcMZg9CnisFYjaH59MrKcjdT
5D74Cs0VEgnvGsJU+jTToK8vs2G1CQt60rPmnmc4jI40Tl/nfDHBQaNDUXh5+QnvqzQEzqHlT+7a
mwrOdOk2+qlKCyOx3hdqhfT/i7DvUOApXT51ZW8aiLHQhs92ZFucRBGMQXWcYecRLQv0kmtwx79u
KSKeufNcduVWCLK8MPSPnAQdfrwwHt5M+4X8mxc0uMdonW7fu7ybYcIWRKS5z6T+WEDFGZRFvpsl
sP7qoxOyWJynAgpRpSoe1BQJD5vQompSl1yeD6SWUQGF8r+12IK6z3yeLwaurMP2CxVUMsvjmxb0
Z+IF4R2FkAzw4fNgSUjC37dZi6W3qskSR381zLrYWbomg0Mm3VAtUvf868X9njRvVVnLTF9PckL3
/tE0EKFQnBv/tS3IyNdvqm/zslPl31gteSMFE7M/sx7wPkMUNRjDDN9E5ObVraOZdttS99trn8YE
mnt3OntfJLIlmg7CekAVvY4+bH1NS8+1P/hmF7j+NyhU+BaT7xRyvYUg1hsvv+i9/w88Qv8pL+cJ
Fwo67728Q43q5WTGnY/+9fKOTQZqTb4ECvg9jqepRE2FLDrArawEJEAw5VJVxXOF3xayb3W23vq1
EdQV9VaMMTZ56DqiRGzRVxjRwSnxzt4Z1xaSp2bve2ug+dH/nyItXy4FZldS0ORPS6QcMPTFn3Wi
6GcKZJEou0fk7WCZK97bE4mCPUma4uWWy1Gd76Pis/DCLwLCmYPFLx7RVNGvi66WjaovoYIojD1k
3nelLQlRBUeRNTR66cSdwN+pxXIEKhE15t1u/CKNvYDbsz3erLOAASYsrLCWUf+odh5/9Q9x+NAJ
EMbGYWb3WJ5uXsuWGctqW73MnTnW67yLJr5B8uJKrWdbB20E9285hKC16VKtau1O4B8aDBGLtwUy
oq5FJ8e8/cHeKE+7Oiym94VCxJ+lq+yBM3E/DjaQToGO2sznJ4fR9Qm1/c0IeAy0w9vBNDj6Cgrn
OezBz1HsP+YxHYAVGPwkNVXflEn/IIbhpPrUgz8xMPdiGBSC3wukhaYDMc9OzVTBFwMO5RmLV6yv
FJRrRFPZAki7nUwMb0N/zdBAIk7CVhr1LMZ9Sy6TjNEdDcjU6+OJPVj2WXoPtyMJbHdi9w51JKBM
B0Dep6gKf4uQkTiVAIOajnLmY8YmLmFveICxRw0Cpk/sVudw8StsEp+1q5N+TK+t1zYt0jPeaafN
xThlnHC58DJFE9tnNgd/e5PYv/ZdDMwlloH0paSROnn+PBkgr2T9W+7DI77rU3n8Xmf/VgKnyU7+
0k/ihF4jzgNcrRiESL05NEO5FahNZZiMDWGFHauTw2OBajno1muPUeLtTD9osIoovi9oUr2XVWDN
HlrcNqnBQ/sDISOzkeDRGBsohSRueGbZI0sTkc64fFgjciuh8uh2AnouJda9kOCYSU3Bc3TOG8zV
We4fsGOhR08P0r5z6uSfLAAgI2SpribH15zLzlrY9TRCgc3SFy1ct+5wKHHTrK8poAITpsD+vMG1
+2KLbClhV+1g+3dd1cvdVZP0pzGUZRDmtv+tap8udA1vwJO8GikLV2gFl61+/H7+5abaf1+5pXIk
4NN434iAyLs5zFS2bLX4PfaQ2tocHpeZm8boHYx/s6+kkfBpltHVIJQotcbiX1Vb9qvglV8mnIDO
3UlLvgN4rGRp7/L/61rnIfVRWYeYQrYICAySdEC6snN8VUxmcFTjRje5ogG7G5Vu/oSqlGStdjQ4
XLXuA01BO9fmlOfJyar4WQI1xFgHBk014j5H8Q4ctGW3I8R9PNFGGp0FmhZCxd4bGtcpUq1Gri4U
bpqWOds33RSVXJocEwzKm5E4SPO/iZPyclmbHUI6HkG3ceXCnzSQJi7Pql4AxftqZA/tmbktoemC
7snnMtA0ZUZxni5QUz2TgjWiok6ZB1ITflVOWPnV+ByaVOoqOBiwN+7SjjbUFan7uPJdHjPWtywG
A4shdcrFpgcwIf+eQCaKoyk/h51lCbFpC7jZB+mIV/xIY1wxof/GarTkrqQE3KFWFXkb2nn22buY
xJAL1z1m11Xok5ThHZ06OZSjTfjkqCsZnO5xB1XKbcMUZ8ypt4yUSOjJ+S+YKKV6nAqTv9Ruhw/U
VFUqxXpmn/0W1jdUBcf12hAR5YkhMN9zGtdXVyPIwwtGxJABZuLHh7Oc25zSMFjRjIk6x818YVxq
9ogaAFeV/474p7QpjaMtG1NbXS6Urrc2NR0v/gNDGArWXJeuwQg5nKnqoKiw2lASgJl+Ej+OxEVf
sUDMk5pTTXQNP4M5xHy/+UIJxyD23p97QHyvM1yRFcgqpVMFswlKE1NxLNa181ue4JIqTH+wZY08
DyNakLNV73uuaQTy9MlkUS7g04rKhSt2x6kyp+kkZ8rhPjzrUvuHdy2XKOIbiGgqNkx2qzHvq14A
xcx2geGttm3Qwu08xY75IvvoLbgPO9TH3tDnkJ+dVGdZrNktJx1bspgFndDPbu0kKZc4opStLRV5
vciR9tgkLWqW003k9YrT75otuKLkmx1qZ2LUm6oOGS3xonWuEf3yylJiGsEwfG5K+JBlsXAW0XeT
RQ3zfQKiLpSFndOWmhhVUOcxyhVOE8ABZ8tjEIMkjIoWfR7a3CzJdsulukBYiMobDtNuM9819u+X
Ee36jX6qtbcf5upDXe1uRHAHt0uBVyGOce1mstEdQg60+KpMSk2KhqqYOcgGViHNtp3mv0FW7sPX
iechWc/3Q57AE3yxVA+EmtgEhALcEm/9Cr9H5hLwb2chGRVGztsPtamHLgng3zHcUBbEoW3nq9LA
Ft4KB/Dc/TGTCK64UAiuUnRBa6sv8jBX/MRn255YpSka3dPbx80qsWDDW2DuICN2GK9+La9gNS0e
X45F4S1utzlI1puA6GwD4zphturCio6Uu10VlsoA6jWZGXsYlbVUSyocvpEq4IEQTIFmiQvcAES0
dpQJq0z0C9z3IVVwS/+WOrffJARaD9eL1pDgjIrxI5ve5LQCqMi8rLGsX6fGYbSivhcO+MlLIneX
hyGYhMZ3dhgDt2Xx5I+RPrPxQ+4Q+3+Mc8wQB9dbZedlpHAO/S6V3nM9UASxMhJLRcFxm6VflkAb
ez0mO78r+VYYAyuG4byQ/CdX6QvSAufr3h05ypkSt8TD9FM1G3E8CVmFcQ33Urg9KoySFnmfNzFE
tQppGwIl7t3uCJt1x+hrdXv0Qj7pvley1SIbipKEUB6htnxBGd2xlybN0Vr7QhQE3mDe5qvTCUG+
sjx4+YPsaWFGoNMHioKg6WY1UsuVxiyrqVpANIGPpDYFcOa+lKXWl8Sn7g/GpB1iGRYMXkgsb8eP
Yt/c1qPLydCQZsXnTWVFpq23sjB2pw6iELn2869tmwttt6VPJblASqLOA2xXU23fpMAQwzmCeTBc
De7MFud5Jok8+tJTA4Z5DfQPLQCV6jC07m33CWVZLEVBKgOtcZNqJv2PImR6GEFoFjc7C30/5U2Q
1tOT+G9sO7m3de6wcCBNUeD4N9zWEm42ttoiFqUiUJg4p7S1vA3N4VgJ8us2RDrWbnn3Lzdc3Ddm
EPoMavt8KhSS+W1fQc7B8rkb92cAC0KY+bYF1aD+kX8dn1OCt+9O6VMzQB+SW2aEwWCIx8NNVf5r
0H+fpUtVAbhaU5KLB0hwXyKe/9+rDKcBi2Vr4W3DwRANUmH/UIn8sBb5BVxZjX9N/8CXgi9erEXX
K7rQ57GCxMSjZKi//Jw/DiXsO4fOczgu2IyTVBEPeQOQ0jN9HRf0Nx1J2xxwLawbchTEe2IAyj57
nPsyD6qBYCUP2l5KEQLkfiY8oMqLv78rGLfjwu+356Esa1Gr6VYMDiCNEUgPKC01qrn34wDq/Qvo
7YcPCZ5FSeyP1jklckvjUUUKBMTY6rxIY+/wuGpH23J1dPVzFHN2Fpw27UTyC4tDYHHOxD9xy1G0
SU65Qr4mFwWAIwS65JOupeNEAQFu7+rtpsWsAu+VPaCoHV5mGXGC0tw9L5DBxaMYkNIsA+GutLMD
ezwz2c0U0d8mugYCTSJBzWRa7QBgjliRxdO3mdeFOLhveXtWwV06hAW+KGt4noBtkGCZgwLtsG7F
NlZlY/2aJEfnDmt7aYWwi7v4NJBoOcTY6YmOd/iu8j/vZ0lD8OnYCgfMik4jeqyMJZVwLZ2vS1jK
5k3YJtvyvN6TFwtx/IF2/DI4UEii6KqOz1v3ZGYEQAbjZGuBs+bELSeX6U9H/aJbLKmtfRZTo+Th
krKoWqAdb7iehvZnUv63M4UV4jd8CLGtT7bwe4aGIZtl/jogfT0fsE5SjBRmESnYgkA6AKITYlCA
YczR1uSkQU2sxg/qDYJG+9FIyQzVwgVXk8l0M6lgfzHBCU/UmRi4KX30k0UUlfjx08pNy1XamXRX
lAh2byiwf4wkGR8+AxYqCdYEYqD724KYNpj95SCP4xbnk7KIIY9iBaJxtwf6U1BBOOH+/6PGGbtM
a6vWSngEmgwNudb6h7ySMMGsKtwUP2wuZi5va9nTGni9viOUx3f5LS9l+MNF3ApvvQXCiGwmpRfR
JtiNGQqbhdp9Ra+m2744lNMvjV2Nrs5gJjZM+JuUgCsChFoGlLUvt29bFev6aCWw9yzNJqbiLAWr
3jXNA7/jVIb/xt4X8NXPGsHDyUhSpRzfqU1Ps+E+0AgYpleSHe3oQ572zBVGm683nCMq/3D4mVUG
VyGEN7O88Rp53AfM7OeKlmbJXoqE7QQtFkMdb6DTbOaxNJyEqHF24rUynw+n9IQQkdFtMbmu1fZ+
+rmbattPTE2kex9rsx/7ZTFJDcO7qeEGp8d9AQI70j9ZKNEwKzmZD6URWReQWbsld0tUVm8wlRD0
zTAlhgHL6Cfgah/LfQwKLooTPmcXdF0UkEwNWbu1XB9tePbtUZ2iFkPvEcZCh//cFVRF4g+Uhs/l
Jo3a4XQ+Osqq/fK8pRUioJnYwU9J4sc9dCsqyMqvbFX0q97yYcAShpD3D0+02ab10HR0FhB1tNs5
gMhW92/4sAJpCRhJvH9Ch+nyE/bPjqRM1nwmftaG/vH73Q0/k93GzvAzyfYQoyL1NAETfnL8d9GQ
Qd/tJjkJq9tsU4n8qiYhHF9Jm2SpcMXsqypgOI2jPHQWbC16Vp0VAplYe87j3fZddNqYi2mJSUvX
xmeuQQJGuzfcgTlHg+YJLTBa8k//tIr58333XQGGqz3x056MHWf9G+nZfPyCtFLENs15f0Fo4nu+
F2Tn3ULnUelk8/Xydg1EJUhJDn71aauFn9m1/1lt1h3GnntkvW6cjZ+fxo1PiKFxZIvxhHmIwQmZ
VD0hSXo5T2JWFsuTka/HQ94w6ncaVLgvAKpSavfYVS1qKwYzlf15qgCh47bAYvhmpX2XoVawuE+K
DikPm03+NTO+qU6akCkmCjNgQsiMtDO2ZIpkgU6KQfXQ26UupI51CeLKoL/GyHzR/vKyi99meJ3R
T4IuMapglb+IV1Exj3cTed70YiWG01/h1bYyyTmmcW+SSqd6uN375KAdKhoHMDQ6xN5qOiePrM14
c0RBcg/AKOtyGfBtGDYjO8O4nagFnqckosq6A5dyxrUQv2v1TJYobTbZQ7IVDRwXogsco0h6R4DL
B0TNtyG5wVgvpn17rhpqZv1GnJ1aKDAKVKpgUkn6q0oa7zwn+hWUhJyXf9UlxAKjdf+JFFlcKQB6
FavBj29BvD7pIhXqztcC/Ofy3NUBEjvMzLucdGeZs2oUF0MpMbm0jPV1uxjtTFpNW1bJ9D4dMPJU
aBTT1ckHEZUHLHPeMWxxB3+yXTjP2SrWu9uOX8YP329Hi8GhkzLo2NPlL9XpDY+3EwUSDL2Fjxe+
ehK6BsuW6SL7pAbzCUe7hlASJi3lr+itLnqF+eR9XP3h9qVXawyidYW0ELIBnd//VFzjfVbYPDjF
z+cNIjRtJ0df8t1iX+NxhsEIr4QRkI+OOVIJ79TBY8IHp6IC6sQGGVFDZZWe0cqqUaje0Y5MXdA+
wz+QVEe+67zVKCjVCn6IN3m07gqtzkaOYTM3rnRsUiVRFvQzPOhwqRbrHJF+IJCQ7UaEdMpa1+l1
h2Yl+ZRq0+313fIyqB3C05UlX8QzQvq3+pv9H4A4CfrwDcHLvB6ZKFrmvWPCusnTV2jZpHz+ugO/
8fo462TZ2WJIZ+ZHsHNoSpR6K4TgNWFlx9meYZhsv1V+JPVLvVdM5iUpV5wjAkTt94VXQdAU88f7
UOE4tsPyuX8Xa69ZCb/L4CRs8v1DEeAP0QG9RbWI69XtjHtwb0AMAvKHU0CncS91TkCAK5ahnwIh
J+wLwkVHq61hFnrS2XzgR/cdSghFF5bQUXsIC6sKy1VL7PMJtD5Qf3bxDXVwT2w83FeYl41qrLmn
AWisII8LFJIT622y0QSqtrMFQWVUP3h2D2qNgaArcUkjEkVOu7XJDGKM5aVT8wZQ9IHvtEn/VfmM
UW1upj3MITo1XSxW+Z61Gb4s90dbF1EaorBlwnESqN60vDhheeRkTf2P9ijcCuSypml6cBh7g86B
7T3GgyJojK1ILyWcWclcr68gsxW4Yuv4DJ6TJGWNxT4IeKxTmDfgJC0fZbwNJAvRpI4SUkuu9+T0
+LTV6WdSJ5fZvM40f+4jkfnkzN7KBALcx0ckSrx6Q/BK9U81b4adVP7zBp3gLtSHJ3rACwgx8JAu
A0NTMSsZKcPC9rfW8DB52vY9Ls90oI1EscawdNSbBu0r7tpRMIRYuIRTU4ZZc36ks/2GmBReXldx
LIy0sAey2KbdSnN8jv0RiHvI4enlHo/33j8C/Yq0B+zdqCy4G1qQ9ETtXlc0ca1ZK4797br+xp8i
gc+wD5HNj97BJhVWZBCHj7/M4wJLOHbrSo7gjEzmVM38lL1Ga3RS20pt2Z/YNctcOFqCdt2mXg5U
SgAlRSsL1hdAQR3YMJw6+yPiFFmKBYXAhBZb54K7xKrcs9XBeOhBBMaN3c+Kacv4IvBnTBZxhDXc
IEUHfX8Z4P7nijBuPA1EH2mDUfoOS9cgFAUTjuByH9ARgM8pgzmZoh5IMa4i1V3G+LD1LLSalCyN
rvLV0cwvp2QbdVTTNMFerE35k6Q5I+eOtE0fmwyr5cY61FDwajJWGkKYC4xLXGZVdz53gZayi2AR
D0nt2en0Xg8y53douw0pJ+yGUXef2LjG7njlIpcJUWeKZLbQVRuPcyGyzQzdPZjlXegf0N8DSuqn
CxVg8Ne1q8LY7l8XjV+S/XYTdUAmMKS36vln33UB3DB2aXnq86cjHuCQ6CGwf3TYpcU3X1FlxXhY
GKqSDO6QIcJSVnJfFuVhniDNwtkzkq+gDenLmhT3NkpPLPwGMffXHWY0GXzYp9b4ILYbfONif+zj
KW7GiF2pUEQ4skpw2i+MFIwSpiccknXBWbgXytHpCBuEBawerkuAJoKe+pM4STK4giDJt4Mo9DtU
CbfZTnPpVCcb8hbUKdeGzd8FbJEcg+YXMW4KdYm+yM32Vf6Lj8KjymTi+xUkKQDIVVsUl3UvmNyI
eskNQjNijXw0rda0qCRfZUBEvxOMhUradpTqMmWvTG87f4HKWXDHv4/TwoesqaYJsT0qx0zVPEWc
fINgGQZbZETRxxHwGXakrfSRrouesrSFyouF01jffzCwB0+yc33iWWTvOxsggA0ZLQJ/mDi+zXY9
GEsNMBsD4JXJBnHBza+7AF5SCWeeti66K9SwEbbHJO499KjOLHMQ1Zm/PA9KW9A3ufOu0G9hzHXZ
Nt/NcPt9MGjI8QRy07hgycyj+4vFfpMiowfowiR7rIP7HTNT+s2NGLKBPsXyldq/cWPG2HoxVVVb
FdmfhDG3FvL7QgBQdivGKqj8D8eG1ATPkSzQNL0lDH25fNwkLUZfZQKfrcaweAOeghfxmnZ6+Kxp
bnfQbcORTWPWIFONV+1WxMbWf/HHo/YfYT3gyN4awbVba/Vq73KXiFIhNkGGR9GIP/4D35LL2XRK
3ODKrF+1tF6EXSNvP5Dz+4F/OPeknb5XMNkkW2FNuoM3b4Pwc/iYlerQeX85IAWy/+Vq5RSKIQ58
XZ0Ez5m0Awkm6bDEKOOdRHXIayO7Ff83xvcd85999Wd7tWGxjN4fDE/KE2/LwSvuUM8ACwbBAUGX
WyHmtYNYLhGMEVVCdKyODeDT/5dpTe0XDGcD0Pxq4b2YAWQloyoQ/J8E60Gun4uzrbgLaU+sMSn6
PlcJWHlfb8ML1Jb1h217hqbGxb3+Fr4wP9ohF1PI2GRojk4p0e+kfuai4VPWBreMLg2fQ+9sG+/O
YEo9K3JGx5bzKz2OPrA/Ua086TCeMMWEg9k8koE5IhKgVgzQVgSr3NCyVVZIvZUc9rlNGqdBIpiQ
Kjv7GlHSnfj+uiiFow9A36BXZGe7DQllpKloWex2z0t2VBvDW06FXTuyN1H4AdgqyhwhYtsbdgJV
MDHf40jlfWgT/LMqN0XgHRUSAk0yPHKkKHA9K97evd9c3KTzBwya+GowKjy5MHZDAQlG+b3NFGmv
3O5aDmGG/VsmbD4yXpNiK/aW+4wqtGoVrZcBlSr2PpRJM1b+2TaAMWut5LwcoRZD/Rk3Z5S7ZrI+
oqaY6omiM2lbwVv4aDl0fZZ9bKyYS0OV9OK7N35XH6U+N04YhCocRvLu+BoIWTXvy7VajyMRzSs4
gWwVsiyK2UBMYNK63PP7errWBneHjk/bmkC0fDmxnQzHvE9QNxwdeYAAKtBaBg3qE5CyZU+C++R9
k9WO0TkBtGFbtQMeazbr2Scg+8s160HfZIw2wBnJ6JF/pNKOtP7kftvq1zoT438485J5Ue6ZqDCU
+tmJeE+pu2K1mvLQkGYMgqlh/04pxNphaha4HCOtmbr+/UcZSRAykNo/C/Nt0jC93wxtEa0Zwvll
arwS2twHRP5Me621XCrxjJ7yWo2Pig8NDI9JtTbrZTy+K570fGV5ib0abhwmfDXOEBOygENu5LvR
w0Rbk9a/4k6MZMx/I/w89cEnxqjG0Obh7h9lH80hT9FQazYb+FKSdLxLMZXmGZdsONC+GaNkJEa3
Cjb7/8VSytRFAnmFS8CSv6M0tNAxbO70N8kqtM59EIIZsyZXvQwu2EBMSpqe7Xxjr3D0WDaBEdWx
+9qWshfWoBS3jZKKsfAk3HdZCHktQzOhfmwuANsCed2Y14C0agdRO13Nr5MEfndVmbebikTDsqE1
65Lo1LBYPAUGzGF1ovPQCvdTlFBV7jDefQ601sUFhQQHvSGe8TboxpOhlrE6U5btqVOKZAGzdjqD
6YxVI3/iAHtU5QODwHVJ660fhXM4TXXW3RAXrlliudwe41rHby5WGqAYwj7mIrXXsbCAgza29vrk
VyZADSyodMaN7fPLOngT3SmOFRs+GPhBB//Y56b8xNk299ZlEKJZJjv8vzsYlMjHsCqbR/QXqAmi
yzJmchi4CDyO0PrFA63VQHI+6RCBT0j9VT/m5RNULIL6s46UnlU7pe08EaCIXtGSGDsTNw9HxIpk
1WPNDi6aOCGl9K2j1iv9ngB1DBZqT6xyXKDRQJoOrezziJOUbxPOpDh8iqLR/TL+rzgllLVyPVoM
HMVklF/xtOMnxMu3a7XNyRywp5oWz7RgMnwN2wGUubvSV7C2xFKuwmXNEmSSQh9ksY69cPU2RvJN
Ca/aSAgg2ztidm9Ou/Eg9Qg+/jaMUL4KS4Z/pjYHtexQ/vZ9p/UESz9j5bf386qQsQv21+KDkdD8
v5CSS67CpkkqQbUzGOQAbxnE6vJ87PzrWB/lVTYeRIaHwFS0ds8Z1WJYH0L8bAc91R8LTP91nKDV
QBmJ6kfpPj9By5vBVnZAuZ/1r874owGQhvfhWweXBAltGB8k39/SOenrXUvh0ET4apGOvEaDFDcM
U58OiHFw4zu0zi6f9CXwumXWCxg8fxY3EUiY6GYVs3DJHRIXPhd9H1ZKwfmd4hwX+ZoXjhNfQdCu
IH7aXsUe/rcrMW2CYo5Aa7xA78wj7xbIrsLjBNENw6ClFk9VEuQjKv9Zz6BmnW0+CRGYCp3RRLD1
2yFdnLBrsxZSQ9YilpNzVmEGaqlNmpSGYj/mv+WotAqTSta4SOX1aPnY6p8VVG1PvlVSbyyTSA69
aMSbhSiZsIgdclCjAxwT4YNhZOnUkFDIduOVwmQr5RMPZ9kQPaobwOYZt988j2nXjDmLnMp7jnPw
mJBnNHn+aR9JqaCBf0aY4qR6Rzv5kCDqS4wWLBCHQio9rF8HYt5Fx9Rs2qYpeQ+sq5UiBtlVD0ja
KuKWiCmnnoZBIMmKNBw2pQDNQJNXdEO535s7POC7AmO7O3nd6fYQzr3BVyAFtgoHcs3zEoXqhBRG
5e0lxEDOcdATQQmO9/Iy0yu0ESvbXusjAbMnjRYrZwBokq/vfbBhoJ1D06Tcsv9gswU2MSt+nWWV
A9/t7DmLCjUJf2MyhjiOjNtEY/ASl4O1cGKu0sAppxbfFXtpbYjn73ND9ibBVoe8y0miscQPBTNa
+/DXNSCht5rhqUA8GXUnoHu4ZM+gktX0VI8QLGSBBtk1kSBoy5FJmxwILpnggxC7sQsSf+7r3po0
bXeRxW6VsWMtmC+/CLHbrH88gdYopYMHn9kZ130bCDGtsdN52Za+wPw/8Qh/7iCKUsQtHR15aOXV
tSOaDIgUgRAsT68fbTBWjxYPzsSl7h/ks/kwHY71gbiAl53hDKlnfynojzKSwQUMiDtrQpLlMkxn
9UXv9SkozvLpUcD44Rcqzcm5VO/AzrcpKpcbS9Mxy4wSSmS5a7xd16HMgLaZs135yVc9YcjlVcbs
9RIdK3FDxQGFNzz25KxlurK8jiQnC+2z62mC5c6eWnDh25H/n3iSxK1o41+GDR9fkkyqwtr2kIhi
seDqv1HQG+lJpbn4tWb0kZQACh3Lw9ZQEy9gktn8/jEFYTsuZ9vgf06nr+ynlG5Irt7mGizCrv3S
6/dI/aUaN+KGTLZW3u91sOZL3u00J3LO4Jk/bLzKBgjctU+B67ONA4Myq6j9HoDNHYX+vntCxAZF
lj8ekcDzKw12uJVbzyerYNJ4Uj9hsvmSd7lprr+uWmRar7Md35cXAGG28MqRKPfleqAta3ToP6/N
dffbqUQucTOtlZMw0UEDD+WPTfiOg830MKiq5deEDNHyLfnpwbQxq/UfdzKAzwlzmcN5CzqkXbDT
VkVcXDXGdR6JFCqgHbwPX2tCivSJIuUK+Qb2EMM7KCkXP+T0cXzSY1tartc2svU3YYXskNGe2uuR
Ew8nJJFAqkli1tW6nmTlwNDAmOhbIQw4WVZrZ8ZbglE/WN8TvDgQ9rHiTIoGU9d/X8a3hd4xRMY9
ZtgkH9vv1nmWcZnKrI2l6AyRRnKgrDG51Ys89nbOHbBWsjtA9tIdWjGWa0N8C9XgpFcpuCPL806F
nFjXusZtLWx9isPLB314h7sD8Q9iMIJc25DNoJwjsCq+2yYzrl88mR6jTpiBtEV23XoEwqkYJTGL
yD7stv6wQBbXe+dpPidEigJ30QXlBdnKjvtOw8j8ttqNJaFI92onzWxbxWVjVpc7vgTHpPWmZJKM
A3/8JP62dwJZr+g5ByJiadYyLHDGabOHAt/LynF3fitE17ZGvWuULlJU2p1ehBnCl8snM2iSFjU5
aVdf9CFB6CAXMcS1TyOWW8/9CmaXdMOX2k1+WtkEBDUEQYyuayzHNLA1bUTxS0TihFLV4DrAFCU6
74r05lCH09L3fpNj8UZSca6oRtzR4PPY0dHjnC8qF+P/ekmlY3S1Vy/oDo/YCHBIy6mGuX3IyXnG
vr87c/w3avzK/4EpqX/JdDAoCxNTLIIaUI70D5zkJIk9EQzvDUuOySCQLOto6X0TUt7wRIVm+4dL
c5Cfd5iqiaA9PWWR9VeLbG0dLSK7ptoN7e7SE/GBD/mUWoy1pUCKhDBUwepEJ7NkHzyIBFo8yd51
nj8v8zcd4ix4fos8I8IlcdwVJoYNgcetK4V+Q6FR+yul9U882qbeMZ+A8FtaRQEtv4DrsrSjbYv4
lm8ZpIpRjwV9FZalcXYiQxvPHNlhWbbYp20TShXYdsdIN+0CA23Ye48C30s/YHChQ+yhPjYjV/J/
CIFFCTGfNSUNkMD5xLbWxqZsdN1v5TyIZWzX4zEozUZhHUS5tVevcXGJz6Gx9YscTGJREg6KTxt6
JgM46S8U3TIIRbw6a9baP4Q1XpC8iEir3qzpmC/I9WZHh3w29kS6g8wgYZYwyckIOF3MV5cwFeFp
igLr+JMdMiOXEMRcnjY4RJlOGjV7o1iNaxih2G/lHXn8/sbpBiZfZPxBUyyIWYwAZLbYQ/QqrNX1
aeEeQKzxJdPYCBSIXBG6cZSQ5G2chFNVNDW5m6iJ61RE80hDCK+Sd76/Q8YCLLqpS36ATtmaWqnp
YGsuMpTewUWc0LnAJqvAf45kESaED5CADFWhoFsn8fbxZtoOtT0gIaMWrOeB9NpnrUyZhMl5HgZy
qwI4LN11tuC8SYULnRYjzhlp5nP4OhyHmOrD725nVNJ8m12JwX3Q8yQLjLv4amk36p88nx9JTX4O
396VbVXtU6BEQ6LUjuC38K7zdF4U994GJ5xfGT4Lbj1StW4fts+rIPL4v8JarvLBj2n176+gyRIm
v0qKQGkp+Ws3cEfURaCYx8y31SdJoCQOsTQhIp382HOMGxbzLIFNEKttr7q/TRgQeOAIntyDPJeH
3gjMZ6XMSbPW3hM0EZTFHlkdReJadqizl4tOYXTqr83TrkI5++bEYskoKptz+A3nyuIZWmcZP3Mg
X3UrZ3SouO0G2ggomlAVRzldaCzH/AXWCBuG1ZrhM1iS4Ad9iMrb5KFOeYxQ9U/zyoFIEH0px4R+
MrISXLF6TgM0mvKYir36iBZ0vvWICYtcMgjXFoYNsYV7fgJt2hkZrNVqAK1aDtH4LD73mqcgwiCj
XXJJd7Bvq6w+T8OzUCpbJUBOkPBspKIXrdiZS2YZ/HdtLMCvJUL9pbdIoxz8m1bdc7BhhSp5TGk4
p5tV5T/C3NVHrbCguPRXTwtcO6WnhfVIhX/rBeUsphs0Grim/GzuuofTIMKlpFtYyij4rNFpZyox
YAQHhAfC8wemOGLO+uyhWH7fcbD5HpsGtzBAK0GrobfjJ11Q0scKSgbwBbr4y7EenTRcCv5qeoaV
GoyRJ0gJPeTLo6lZSphm9Hrdd7MA+gDdL4XvscJGfw74cE/pr3FzZoO10dxUWOJWs6BPLJRvVYLI
BAivQN5seZoMtRoTHquK/agDT/VsZmwHQzru88LY/hwaCWG6oN7gFyAv24tCwjpApah8zX70xpOQ
kTsP9SyFoipQNfzorNkp5B5k8w8Yhj55LSkYerUKcGxoGZJFuHm7pPzqI0DryFLvhZDtCLn+KCSz
ydu9arvAm4cd13p2dO3v0J5qdHYQWC7RFbabxg4ABU1jfISW+XR3CFsB5d5SJJbKeuOYmPt7+Uqq
tUli7LNz3la4FZ6l17wPVfkk+K+Sh1nQQzZKG62i6NI29Ph60LFP2gT2Xw7JwN8hUzAlN4MNyWdL
/aReJXUu4Kx2R1zcGMK6pT5yDKbw7YhgE9hPfh/1+G7egK8oVmorf4L6Sjy6yoBHqvW/SEfeXUn1
QYYhlLV0HYRskc2dwqts3z6sMYhNrcxN8nTG9dZPIkqme3eEtGGzqY86kPgEF4Z318Qloxy+UkCy
2zjfx74SX8Vad0lmvWiwmYyjwQyE4ep5tV+YR3ykjmsE14wyLtq7AsR54N8JiGsbv+8CQTxTqAkZ
nAAc4zPIdrlEUjftHqq1NzOrxQx0EZ1PwSzCJdv5kHQJ6NdcjLO6f4MFNQkb8EM4KSbgw6xgW6s+
UXAoHP78RsUNCBNIhM+JOmct7C0je0edhQTg6jZ3hngULD60ot0MtrNmGhiP2Jw99+MT0CfWTCHR
qYhrot+XUgMQfIM5Pzr6T4VE+EHdGViuzXLew9Vdriv8WKMnfXpDiOokNPZ7SRmU47gTc88/Qw/k
lYEPm3IaAt+dGj1nBkQy0pdGD1z0vfbZD3bbkqhXMvweGn8+YCXlnBb1Ou+Hd4HGJSaIkQ93REwZ
cV/nPK6b1wHZjqhQ7cbu+j1G4l677NzI8bpjQsqZeNSi3umrxRwBwb+JO7nqXPsAuVpxSa5XrcNh
4mV4J3iY3aoWsAxGvlVxQeYumb5qst8DeKKAIfeTMU3yGj0TdCZgPSM9hZVgzRxoDg9Y+dw70dFG
Onu2OnuComQVJLQb0Ii5Wd23jW95k/BgDKYID9K4Y//ExJx83xb09U8ugz5n7pCwac33buIlxlaF
2tLDYVkD48re0NP9Iz9Owg5wom+bYCyBHR0T8346IUzOZ98oy+Q7gjp71kAYJIb2AU9R0AYnfhDs
shw94oyeNdNbP1eDSeXIL7ytp6FWnQqIMhamhTxrVUzBPzyiwWoufAV+qFMANDlAKamrQVyJWlVv
MV7vvDnRuVhi30pTo+9OFsXIQG8iMCliMzrCoI6N4D3C/XlHjXP8bfGxDHM4AA4jqRtyEzc3dVnf
0IZlkVnedivpIGPZm88Y/AG4zPEFe0r2Ckt71I2r+UqHbdkR4ZTiildNWmnGjWI/zFq2pN4Wphz2
UD4+oxr8o0mSIdgNG8SbioTXLWMsiKyWop87I3Ol6I6mmunI62mECl4sie5ck1yMTMdD1wSZltxq
q7xRanwykl8UfUZvjpagDObJLz/imK+ELRpoFO0bz3hpa858Mp4e3F1XRyqi/CKcTyvOg9qlmo55
CSJFvliqqZu9igIOvtuvZkAUmhI8MkQiIiKPqvZ0Y60BRFhLdp6Pt7kHFuFdjKogzXQiI76arE5K
NS+V6LcEyEOKzNKL/c06GY6bSGGNZm+dxl1aLtvsSGBC0KlYppoltfLa3diE3J1qQM2DEC2//GvN
wuIoSo4egLucZ4ad7cWQLsQmQoKriIbWhLmv7PRoQmYe+6hSUxEqSmNtyM9aUPga24JDl1MSzFor
yIFcV7i2o/XfXngm8eZrFnrxxsvQ75Eh+Enpsfl8K3k0u8MQqr8Zj0vlcF5ufse2HPOa93IkLAkh
m/kyknFV1LQaIdK4/0jZU35GrK2Z8pPr8xJzSBLyVFzXzhnkb0Pr+7bS0tTmgl3y2yp0wXjqXB6M
xre9D8m/gn8V5Sbkz2MKiPi+q6BYfItIkRuTCktXyDPdXaQiF/j7pPoXtd49+pWgiL5Rm/6aWCQS
hW/mKhlWkVFfXYbKJEeWC7rH6GwixUT/Pkx/uxEKxsUjplWFtIWU+C2V0e9zY94WBP83D9GZqeMt
C+/hnQ5UqBM91oJvEvMO06GroeHZDLVNVjG3AuI50tFdyuAFxSfw9T+a0IZeNc08rTS3p6nt3RXl
6nf5mpgQjou3BXOKTDBH+X5K9aJRTL1gpUCyqqBQwQFJg4SpqiH2QpqzkYNHiyPtmGhNZ9ejHxdx
2yVDEqzbsVBhy9a177JiU17CLhnfCjRmFSXycbQdrpueR559NBdNo1RGNR0IQjimhhe0idkadC8V
ouhfSPMb3e9wgNLmMPP8rC9WgARbWVI3/uiqzWngRoCl61OzETScTOg/6HOcHwNBSN9+eHhfeUwE
bfkOXWg6YuGgPn5udHYyDTSUz/mWnmDs6PPtqsmEGBz+6SeMk/G4GFTZIqurslJ7gKYLiLnutBcK
DF/jJmOtt5FU6PmUZuJ0Czah54VGK8xHi01lYZzVPcGnLy9kwdlHBuH2sK4c3o6gUgVqkpehoTgp
s+rmKIS2s/Z4FlKlnGoL3zvwI9cChkxFbJgpRTveUnCroxp4wwAAOzgtR0ef4Acc70PkhVXHzLci
4VFRcIDNfJMdUigCXTNzEMs4pPwkaCb5sMD0isyf0QYfWBMPPPTYKVs7JO8eBFA966NUq64kjpkl
TCKoYIKLRS/y6Y9NEL8ELugqx+0DIHkwur7WQuN511697c+z2AZaSfo8qGoeB3VuJqkLmvpFEBa+
XTRvVsSM+muhEEZYE32olMbCAP4TesZpqBq7Du1Q63rWyXRpHpU7HoV3BJYEiP65kFXdT42qTf1q
2COHVN9tE2ts+6Jq1XPvrRy64NKgbeQdrClN0o1EWpajFJgfORsyWSjzTc79RRdhMHgqqiWCxJIi
xTLad+Q3GfkGEGGu7OhTOxKFDyqExsEXFSN6wp9/k1QhHUnHB7qBUNJVKgAVFaGCr5hJjUlCx/Z2
n6wkKvXONjaiauV5kDj1eh6jJCIhw2B+wwUAVeEVvHfABPacxrAOkz7OHEGdEZjPs2rf+hv4GhxW
kFcp9SvZTJJM+OhS+8CDjnDFsIgljF6dCnHEc6e1RyCZiZAs+XVQxCldd+wKiop+kP+M9Rgq3Bd5
LnV9ypreiYJSq+mv1u8dfIrtpVwPvI0krlHBIN7prJmkUn6QHBmg3jYH9euUYAo0w50WXFkOakeC
fNs7FOO3AaLARCeJTG5j4I+7ICNGEen6uSEi1RLUZnA6Iyq8OVDpXNResHVQcYUSAly5HPdiH3br
j1Kz3Vrhf5SF72EtP1XtUzoG0HHDF3stystzbMWDytVCrEQ2AsdX9ZaoRv7DEGKzPhO04TecTHnA
yRUggWn5Pu7U4W+rh1PLqb3T9kWKzC/XMzjWO87nT6ftcqvLUSXcF4eAdc/QiucNQ7HDKrbnzXe7
8NUZ95rkn1NfYqbQOHuHl68Uzuni0ZqeQxO2k2v167cPnd6ouk7kNw4wvijJsPYCD2mn5I6sG4N2
dHxUj/59KjzHJ3F2asfAa0qpqAvRqDu+nfkGrO+FqZnJl71Hpc+eLJ774w0W1m1QoaC3STsxY1dL
I6aDIHjbk/tSlVsIFpwvQmplJ20kAdB799bDpW0l43r9ZeIhCD+cdp2UyvuI3eVTLwMtN0sKI3ZK
OVdAZlqbdBdEFhQ6DhUJNI60AvObZhIiT7I+4x4E4oIxbNnbtmRpGL4fUOHVE8H/Th5GCscUcGxy
VAfaQgHlQhHV8+pnq80S7lUy2ZOiOgWhQ5yRWhcLp/5Jz+WiXIzdPWEUrWqxYflLKWM30HAkCG4N
R5hKQlFcefu9ejy/STp2QxKfx7xoAtVV4kqnLP4s4HTLkyGfkR0hqJfBqjWpxrwg3l6TmfdCRS/h
Cfc9gb1KoY3nhmjCLtpzNNYtPQ2wJmVqZ4PxYUlnw0p64x60Q9dkW1KC97zoIrpOOAMHOJ/yGeCP
DxlNQ5D2/GbuNl7HBjr/Uhi8hES2t6j95AGWPGHXoUxWSivYA7Ud16PC63xqCiorQLrVDmHSz2/d
fTKYtqcTD4FB8lyhqJ9XFz8m9YrKXKPm3JrKZG5sqOWU+zY4u0nuWWPsefEH/sxkvFPwLJi6K7rl
FPn/RlMBYvEpabAWhiXlfAqPic2ysgkEgMvteHx6OgDsRJ6UGUMptDms056Wu/63Vj1DpjZFTChz
Vf8STJVovgncA1WUA1PQeR06kvdB6SzwSOCYHeUvepyo/nvU/m29BIGAyaFLS3xyFlO6ITYkeqOk
nED90d875b07OiCCCq3txtHLv0AYVDcFh/a+j8KP8ASPpC/92jGiL8roiX2BuzSmE94GR/O6SvtT
4Dy2C9K1qso+t/J91qgMSmNu412xo93WYcEXSMg0mY3qcjfNzG+GzTe+gK9qc5KMuw70ML989zmA
vcYZoc/X3WRf838JSycmkZufls1Or2X0dfGifSli757bJI2FEG+w2PfI6xu0LxH6u9aedUg9fXgE
9lEgxzSQgBDoTmp63KjeNuwfTdmq270wDA63PAG5Eay8/Qupp3ahi8JyrGwE3XNGitrP2ycpIOXz
zPnrFk168rHeNltzQ1zge26vf38IuxTSjG6JvcOFmdf3K7EqGf3pi9cLfIpIEw/dQsen2b3d0rjl
08iy1/U3IempDIBmi+vomd4lzIblWAYopFfV57n6yYgF+t7qbAF3JqxMXDY+z6jC7A0cCFYRQM3j
QXLq8OH8VNf+qSKj1+KfmRwNxQDlUx1wZ1xKV+Xd3gtNfXy+f37OmXLPHX/sBbzib8A2zx9NzzYW
3DBaA7EueaDNDe47PcSsIeWKx3QNbf59Fxi1WDF1CKAgk9maZsPCoWGlAfJRr8M6EWkIJM6I3wrA
NDX/8gAkD3LYTfeSAN5REEKA8NF0OosRXmR5w80fwMGrtRlrGb+00E4R0W4xQ0rbZ+T2rxd5RQbR
SJufm9R+ZHdUnRIZDkEDSIa9OuP5OLBNxsAyW/ULG19MH4jRaUFxoe48PrpFow8vhTbg5QZt1Cmh
XxfHjEfiD2YG+SHKO5VEyECyESo2f/Tnn8F8VQUEfO0nUOHsz1BxA+ZiRaoyBIksv7ruNvpuD2W/
l4WU7d6lXyiO7yWj6P+dYUbJ7uSALzKF2XLPQeN5dF3gQdH7qzgd+QfxJxqzyKu3pfj7f0UO8dL0
4O0zbnoyA48/ajmv1YRmnLkuKnMh/ExUzjZ4aAgvbbkO9HhNbF7el+NUG/9cBT9xjk4VhNt+USxH
68CaMBnbIpm54XcG14or29ii9ZYWQ51ABFt++6qkPykClZWNNX+NW7cf7FxhibTvR87uDOUdMs0e
xY8sijjuym5HLP6pKtxz6lzYtzSKdoG1/8h87PSWym/haU2RoUXQSXxO64mA7plp6XRAjnYeNuXf
nIEZCXFtrEvqUYcbD7kt1VHZuxJlau4nZJL3eGcsqq8pvQwDo4SZaJWYDxORCXO3cWT2RDzpFcyz
M9SnAYb1srFrEOrQ2GuJC+bvki5Mr86x+2PPP+yjn2cJZtovVaG4t77wdosXJEdWeqmxAqMC3ELP
Bz+0nbtaDQ4gOnmO0Ui6O8Xgh+NG6MNL5tIh9oBvezyUq/SMUK7kOhx4L4vzEHD8C0w7w6+wzpGn
xJTLfYkH45lhJc2hufxXmU0O99/o5xBG0FzFekqRCXGTYXzt64XC+EezjT+uBvkkh5m3lqYRUZ9s
SqT8PioTocciPhxUEifyS/Q+LLLT/NHCogc3DuMbVrLOQC6FPxraN1qZOT1XkaahxIciw2ayDfGb
4WyqkyJeKtekDyNWUlRTmxtE13L0ua2NVz2w4ARip7uOSUmoBFiELsyfgy8WEdTaiN2QTu+J8g/+
sxoHnoSPVi69T++CvqnZbxqhE+EbvVu4hsgZyHSpDPOD06D+VneucZWdg84bEg60rUDbHCaCbEVR
BGHZvJTWK1pSjbzP7UHrOrG6lRTVn4Dfnbu3uxrn6vo3o1DJ0P8nRB5tdCivij5QyNK61QGkaf7h
9vI/NXiTkRgXzYV0jZUnDCmc9tvQyVMn9HDT6Bllvp2smU32su51hZsxY3E0/3IQoDU3fGdXvRCt
5y+cmDkWAKVu7JxcmBxjuUkJgsB6RmzYuiwtFCfTE8P12S1yKcUWo6AA2kwAsZrzYBetf0ghELwv
uVgbTPbW4TyN9bQzBqRz2jGzjxTlCgGb7FyGZ6UHuJK5ZbHAW9xPV+HNs8zAuIbQn69hp9ETuuxE
VfzP6WmkXKxZ6osnuuLL71gh07DJS+TpfAf9K//5zmFXdjaefHv7IfKM0xNwDGmGTU4oRSeFJ9qy
j3fiyTdy3FjAH0++Apg9s6xizgcGf+9Ts7DPAVX/MpwTxO8RLc+SCD65YnEc+vk7zdamplzCv7hj
Octl6gjSq918jjFuR/Ul84H++UMoFrbwjLXJurqJ8VlOar1zrvIpPboRFjF1MiSyHgILb/Nj9VHC
M8YoPv45U5Fs3cfMLDwOBB3UYh3WxfjqBO8JfVxWKkILSA53mkJN1RcXsy4h5yIWmQBlVO/a7dXJ
tw00VyC44bm3ZO2FThAroCfI8fq3P8BXBKZhjS6aBw00S3vLZEJTDHjV2wsoyVpcB79dXBz65hCz
exQoefyXee0TJO5ukKtqYdaeIu86H4ZWEyrFHto7cd1vOeXcAzijZ7ewTZmr4nfuAW1kwQ5DY4yz
4juZf9g+5SJVGp8ZbRqJvq6+J2+wW7cWNL+t2lKaUruGSrsTWIjlA3vrPdQ10azLV5J4ad+89+II
8kTM7qy4SvhEdXwx8aKQlUnl0PaRJ5fZLgOfaKwXxnvuwkclcNGjI/RSPoa8Bxy8wJZJTUjlRi4G
0kgdpxJ/jzYoBMgNsb8MjZpKwY9mCHDXq2IjoSQ5i4f0YhpeR30+sAZbIQYpdYbojzUY6Sfaig4c
42LXVNN5/l4ditXGRHrtIxIZ8BsLv81sUENC4ucWtRZmXfi7480vstbi7hifVyCfL+V4juSHnxuO
jhgPFHs/Oy1GbxaPjfFqNMU/wSuBuLxLrX0Ep+6tufTxAFWnLW6YHFWT1q7E3pnj0ivvtjXeT7aa
/2hecAd0wgAkwGtQg7p7IWFXmD/S1q/e3NG2LDTh7+uftfsiW43W1mTcspdaf4DnxT6c8elz2hmM
rcI0N7RGtJ9Prr/wYiAmfeV9eyaqkCLZpXC57vafTbXYt5PGilkULxsEmDqZPGPRMwfhy43MpBvI
1fXLrx17mC12KZosUaNraoZrdE7q0XlVFjfFwO/yQZukh4hEjk7gw1e/vH5NNblUcOD5I1p4zjZ7
X521US6cuG5C34senGRMWgXTfacPnkIGHZ1sbLsyHY3DPOYDv1+P/rI4YJjWF0KirBJpXd8z3TYZ
lJ/tFRWfHb07iICSz+pbz6742J0IJ4KbLIZap/SzjjnNjmPY35pbmWADgPeuEzcZBo6fP2wdG2+Z
NwnDhT1Gq2B7a4THVQmd5T0ptK6Hb9K62escz3zEMMqX1TjK2AaSGVJWo0wI5CyC17HfpTsBmGR6
SgzSrQr3F/riGvGAcfT5aFPE+osZW+I8tGBqT2ZF7uAusKPEFeAU6FHhOKcfprJojTnXUtJ7Do6/
vHv3rczFvvhOHLtnpsyKmufGrzWJgXIbbL+2wranPG+ezwYDHAATmaAdBdIfgUYJN+jhfwNUARlG
WZX31tUKxEhsLZWbKbmp8DchVTmwbRJRtcCf0TL48Iowq529QGyKIaq77PgzWagMGxNY/yMd0xUt
R+GAAbpC/a7j7kJWxII3n1hab+AHzI7druvxzaDJCJNWyTIJRxOB+aCYv4WPB9RnrzGHhdQo/xiJ
p/a9Dbi6qpk4wulGKPqIAaPmmttLALd3Uuo0hNvCiZRxYaKmQDFxV09kIF+PkIG/WNIsvMDVeRj/
JMPTeL1Tc0IuLle7KeWj7sVSveTG4Oo6DaOod9mTJRqGXTDZ98ew+++xC3VOneg7d6r+drv8sqcf
/eP9e3E41lPck/DYRuH15CIgFNnQ+x4jKkOG6UoUfHR/9NGpCPKvZ98FqEo0yL2phVnwVO4rWOuz
xHmwKzJnFFlfuhnTZKPuvXzUZs2UgBATuKpa3dhfDlPluqe2/nUzqhgwhwWQ5G4sfDDS9gpcnZ8f
6WObR+tOqFDEoOWyZ7wHQDq4XgWcu+wz8KQgyRF8CsSOA+XrAx9nNEDeCjQJj2lWMbC3I3gm6kCy
lQRieo1My6npRxkaRmHjCCy4Q6aMttausfSF8MsgZfyMe1qVV0AGbE35gwwGsHDe+1t4WpVgxtCp
l8aZrfXJEwZSOLG8Iu4XLmETGTfpkhJgTZ/uLZfJ9Jli0HsV8P8To+T2FrxanQo9uI1FE7QlLCui
nkwbQsl4Gh1M6m12oW2qcV1+Bhv47Ju8mltc7USdW/PGojK0gn5PDhli8FEO1ZXpz3knEfa7rRKc
64iHHbPa7dvXqJL4iU8rCTyCsnJolDsfnJSF1Xou8DmifHUTrbWLHzSwI7SsksFhkvoeOrG51bVR
oA6S/6DCe+3YEIqUyNBv3S45Ihuj12CAv66ClnrYky/8HNA9YF6TzSnwELrNlk7umH/JSMqBcyyg
XBT0gVICszPvM5K1688FewJocG6pf10QL+0wUoykJTK588mpXeMlKmG2Kk/dQjpu9sR7ODwErIdl
52IECPlrVmyYs3FplShkLlXWhe+EcBJrvgyqTOTkByTwX+g6j+3CkSPlW7UHkE2xyXDJn+/W0yfq
mokxbQeMzSdOVbo/9ZFTKof+ct+6plTj0sIWGPIUI0F+Dr5AJVfZUxKVme3ypIjFL+8xmdJP5L0A
OpqOxE3wHuyhjOx80RdIsxC+OsfFIu34aY7JNbTsKZof2DTuXP4Kjch2MmWX0VFDMziBM6n2I4gN
k8KucySnUwdg9Q77MV/NPYJhWDuQCXX8us3/o+zFxqLgmMwtTpMqgBI3cIksMtmu5reOE8LRi1ug
smmDssJn6bnhc3k8d8RSxllS46itb0mB0mL6GVckoy+DTXohexmFFlslENyNICdRhsSNPXUpv3bQ
ikjeFhaQdG54vIPE7KWPgXZA1FtorLqKB0wVxEfOEWTGbE4Yhfo+8wbeSMVV134GD/RGChaZsE7+
5DyRYAY91cz5CjiJ14k9AAtkVE+xUlJ4gvvkAptVbMQVcQ6w+FAx36tsTQlt7i5NloLFzAeT5i6a
eIi2Ia/eQUlK3Dx4+t3+mYXoiH+g4aITdxDxdPqKNXHcmkwyZamRm7QYcCTlqKBwmAd8GjcZXnG/
vx77flK/Fnt7eKvk8Fe7vjrKebrbxcmFs7BlRDr93YzHAGqHt3tYNGU4tI+7I1RFWK0T6VIMW5Ir
cHlt4o3ZzHWUsV5iExAZKDj6xxtVPoA2czohgMawbgItKjP6UoQBZKSwAPDznAm5XGWalNIiRd6r
W9cYAyOiSVV5PBlXDXcLem0pn6yf56tJu6z5rsVMZUEZgd19T27STvRfMzw+ATMVvfVmzguaJGnc
pWuVfMqdHluALXHOG9dYPGo6bFlCWcdQTN9Vtegb8k9E2lW5NOr6/fSGlYcIqJxiZe/wt6Mi1qUC
t05jovwlS++LjRIdmVnmyX+1JHol99Cru77TsPxHgSvFaW2cl83f895Do39NscO77F9Whxi91xJ6
uTuy3lf5hCmcevMwW4otzpT63H/DfPeOXa1/x+BF0zTjXtpkYLArS4b7RAggTYBVQO0NAXA57Coo
IwaXL8S7kF59ReORDpdreomYmXpryf1rNOkdRdhTkGs86LG42NT8P5RHhFsrJ0GJuNQMCjdCvBgP
FiU5JdlRT64ZqN8L0PmvVMey+KW/ySZhKxYmiu34poJKSujqd/Jad/L+zXrG/6kCiNZek8Z39Xpm
isquFgpcQO5gCornWUN1ZJaBEiKyXn/EdO0gkbvp9b0USwL8EXFryuMYxC7VX7Zwu7BKqj/qwT15
kVX8iSnITWy2h7sP+fQgHJDeIsERlrz8uQfrOAq3Xh57IRbrjHvoLP7w/szX7tH8G7CI/BfGwDvA
8UWzEkPdrUkHsUY63g3YAYOJo3Z3i5XquplSiOdsq3aFvJtJzTCRrWk0sgfr1RH8DbsYDicU67H8
UXkujPC2TXnru8rWFDsJrBpP9XQPJgZoygkqtzdkeFvGcTLnPqiKr+byRKTdfcHX0eXnpqmBQSvT
QjnX7PlVu2LHuFyA6jcXvs5VWXNAbe/5AeGJKSeib92Wgj/oNX1n/Yb66tzGHSBvepmeIiWwPac7
7TdjsEhgobIuvwnGsQlzQWF2X8BcUAQOZWY6zvQSxStzaMQOW4ZzpEs0O6CIAFRmzt5vmYwmvgl3
08RnemKoWg96HmeMYYd+thw578p959WHKisxjMRbQcOr33bk2hhzRLmRyr1vyTXydVDSzih1JGj+
z9Noa8g//TaU9XbhPC93FZhwszP54ZTPbkQDuUDY4paUN6DBB0eUoJtAiXgko9WtFE4mur5NhnRH
v8WHfBi2kctBhN2RfGWoTU79B7ptOUpu3alMK8CcUswq0x23zGmuS5TBw3MQ60A8CIoA8Tn78tKJ
IMufycYIBZVmBiaKNl7Yh8KyZG5KQpRngaEqVuQeYZyDXHmV6JByfby8aWLQEsVDl6Nw6B7eNey1
JATDFFVJIVXuZVSQ60RFueqquGdPzG+Dx8z5cWHlopQlYzZKJHJAmWXZ32XD2xUinqmiqjVOXUA5
zwCCzBZ9U+eCoSZsEYo25braDJi3WJRS37Gts6KCPkjwOYXXCHM2Nqg+U4Gq4GJ41DAcgRvdbeYx
tlTDLvkOd2uBW4yn4ft8bG/tL6A8sZM+8qjUJfJ0BINNJLA1bHgLP2KOsBZfFK1Eg9Qufzwp1twK
JQDqyWLmNBrsbTtOTvh20+6cki+XfUIv6jFNiv5Wa6CqwYXHdSONEZyD4G9UK9RHEzfgCLS69pL7
iHQOz5it5djP+u+zHJCDoQ/P6eVMv/O1oIgbO5/aS+clhUNK94bXO8KndF1zcy9DICcGq3RaA6Ak
6gxlvtN/n2lXZG5r2MHnzy30o4cMbwWf3qIWI4cHstk53OSDRPmixSoJLj3w5KyZBJbyejbHl4VC
5yfZ7OT4xgDXPzPQR9HB623JqBn9NK2vtqKuXNsdi1vK552H2y476Aj5S6UxUkzO+H1VHely7XvV
0IaV0IcNDm7TQJXNYdiMVOaoQiWbnMnhoymaP5NRM2Qtw6wE/DkH2AX8MQEkt9U5eK0h0nrYu+a+
WtdquoLpGA4aqIdrHqLzcqnNZwXJtG1ambj7VP60WLNcQcOf1aA1tNBsjsvw/PxhrSvKs3dHxyz3
UGcXQCBKjkopFRsAaqJlABQAKw5mfgyJQXD35ztEISD1A8JbSPFamHdJJeeDl36m7hK+BnR71hs5
gnQnbK6CtHuY8lZuYMdw0EFKjWwhzVAelqBaBpK9idFpLoOqov3qoy2mUYI12ZCmU0ju1dJ/2BRl
l4Q+UgiTxXnVf/+ba73MZPSypXyL1cPNKaMXNqbDVlWvct/0yWljAy1BISHnI90BVw3Ecv8l4Vo9
9+tK0ftYTC8YQpK2DSY3IzBP1xwhg0qQJ9CtzeOyzusAwWr2CvTOtEwLmWit3lX+ipUL+Fe1OiMF
4qYNZszV3kv+qMmnvMwnMeiR54oXujUWCz7zdo404DwU9CMUQBXRaU504GID8vZv8j6rSGMIGl6j
l9dEIqooFwDzlJqOg9rsXIP9/LTvmKdcb/aFKYrv2rurYk4yd0ePZ+F4FgxWuLt+1kYzr8W2UrU6
1lWwlMgqua61falLKWHVHjLDOe47GGG0RCmKi0Aa8E+Ikpe8Pvy1Zoi7FikbEEf58XUVR7q3dgvg
h7mP61J6uf3rjxWzsy4ug4zG2W1+IFe6CY8QaDmmpmrcQPQaG5BJrcWvZF5E8VIGwbkj8ZhkgFna
pGJX0yU+fzKrkqbLotnMhb0A0gEirC+GD+PIqwqCA3mzig9zQGXyhLHH7mT2s0cU1DhhWLqI+tKr
XeSQMaVjuv+9TdgA2c9baR9XkDPnCMRqfonC5QtUcT0vqQkErcPpgve00QdmpP/0QU+rYA6EJOaH
E9D98bv98V0sAB5us1GWq1LWE8mbyJcaFjKqA1H+2+gr0jwR4WvT48uRibwTNJKbxGpWGFU7BiwO
IKRgD0mWKc9ylpjn0L2TEuRGxbAMupZdxCxv+JVx5PMiw6XDoJrMETgafjbQYSZms6kUhxcyHx3z
O3r4s8FNTu67F2Xrclo9DxbWpP9WJPE4iv0iQbCQPEE65/2y6vCYggBEQ+50uAAgExX0Wl5nrYey
vl+kBmnd0JVSr+LDYIEvaYXQCOMmGtZa8q/jO2R+ZAo0cliNeJoGY4jGzmrPNAMesP/q3G1DHCqO
tMS4VgUAEyJhglzlBLV7Gbkcsp4x7hbdaJdlRPRh4nLPNmLnQ1YZrcnziPwFgsIER9ZNHtPRNIVt
IUn4ctYIKcFs6bxe0sB6PFi2ccPRXCCSDjhmMRPSMeRPkrcskGMxCHLC16LmaW0lMmF41u01tKFu
wX2wvNkJzDNvQn0VZDQ+YDep8nrfMthgotSQSKcjpX4OkvFrHQPEFFvklvVDHopRYX6iCDXXGtF3
X3FaY1WPaXm2A8YKntxetik/wl/3BJ+o9odkQJtJmIBBMz16Ee6b6AAuZ7EVZCiuf9K+U9WrZiTH
RUjo/WE/RRlL1HggPMgRkjZ5Vb6FaQEHYFfeAALHPnpU3H02JfG01hpYTmuw6qyTu9P11BKlMnXv
i0RWS69n810BzjfpDstMDOMwx/wNxs6dA5tpZ9JArDHrNup6CmGjZlGZCuzcia7e27fzg+JfxT20
eMF4JP+NvDKuqmI2C8D7VOhUPIUPHYqDab2e2Rrj9da6yNTqXABjMjGqdBxiNw9JHgIH/OfoHIOO
XxMvoeoznvS3ofFCGnFronoMEq0CiKa9wrpMzkaJX0winA4aY034EnG7pndEYxIm02Zo6PQqI1cW
F0enii+vJQCd8luMNpIr5QvW4mDFe0c41pEmLAxAUui8Kd14Cy+TWFWd37uD8QtRknC/Z0QEHRcK
X/CF9LIPl+qgyVFJ6f36ZofWvEDSNERQbBzrDFtuN/LjbGyxMZNKRkNdInO+87t4ymd17w3bqf7/
lNINYRBDj50vIASyQTLTQjioJytRgE2UlljpDOxF6gcMFf9PtX+nQH2l4DVrGW/2lkdt50S5aEvo
uHh0YIzdpwglDAXh7TARyNvjMq6IE0g2eZLprN8it2oWfJzhzgdE3msflxsybIJ5F1u1ATNTkNQf
STm/+vhH4FlMt56xRvlcHrQfPS/ixKifOiZdBc5985mVdpIN1EpHZGvpH67m3+e8YCTOpAbnrHa3
tXHakufkk9rZoRkSH4r3dNLOVt/VOm5399ILKLHtmWUJ6okYnfK8ohMnNDeZBDELfU2vQq1Vg++6
LL8qoOA/1051RuNUKi5Qt8ypdolhYxIOm4Z70avSI7iFq2TBiDYEgZK3MoC6KJgGP7Bp8E6CMEeA
fTmKzqHpu+UUxIICc+/sKpytanp1r4UyZmddS+3QzS+rmmWYztPFJQJuEUxVWCtihwez2aOtmILd
/4zjRXSCn8Loev3afVKFl35p0nq+7pzhxAEUJYi4LrB931sz9e73cFM0u6geq9cKQz3KceQQx3QT
jOO73WiQUMW3A+u3Ka6Z44WDX70HYy+dc7Lj/wbb+WwneUPUu4Sepzk6rfFBFwIaYXVLrvslH/pg
PABHpjmwrsgbRFR4X4lCnIxLOtkXW7IsGPBLvphqj6FOktjT8rDrpRSoRnntKtJXcgK6LPSHDcZE
Fq7cUJMjNaWZnNOyM0+aOogXG5Gv9taVVueOIVh1T3J9yZE89Ka78+9zeHJLKFcQ/llSFYuvzcgc
YYIyK66+U8Gmp0PG4W89oREx5OdTKbLdxu22NgotMVroPFGRPy8fkKUUwWRG9onofClttIBRqPHw
rnz/NqcmxcfA+QxuKHYGWZWV7YZFRMLhBC0rsoR40D9nsufxBu2gMSCfoegsHE5fxG73R0kBAkPC
uLbWHacWYXgdtfWgLHM11aId9kjegloxh46PvoYK6V/1rHmdWnwu2l2WkXr4jnvj2bw1GWPWAr/3
olHy8WyCwCR7TqNQ+Z3nG5xssH6WhiVQQAKTFF13UbgAyOpMMPAhL4wPwE+T5Qo+AAo0Ax6vFBFj
DC3ca4LVJ+m1O31AMWC/D4eyfP1AfYbDf6u+kwiF4L7/qyRQ8O4ju/Tm3DDOg/Jko8dzACLZPof+
ZXTQV/vhH5/5Cgmz9leO/Z4zd5BJFm/cIL0NoMGXl7Hby5hu73yOKqTswVQDSGbaJDm2F1Al70A+
ftpwgP8wV0zIN1Adn9DP37mdl1coKpisHTwxAUPFR76NxUsxt+JMZfqCs1tWwIkUGDR5s6cGG4nt
NJRAXOZJeJUKR3NvyNE4Yo0c5LjuYDhewcgUVObuTN+SZuAxbaxD99/dJ4hfT8z7ksd1Cvw3MU8r
Njsyce5cWs/hvxbUlJqXpscXMEvAT0py44fLxndVTItoMSwBWmzpCCKIj8cAl8czIaR+JQ9fmDDX
R+Xbja9vdzNmLqHQpawICJEegXYWXj+3tVSKhhnSgVBly8awS/9QhSGyMiF4SWLJnKu35JnJ1nGo
vHrpvztBIftobkKAuaXDrmGa1Coci1kyYS5ComfbOCWH2ieYMNUHjYGKHoDKu1BEFb6YEC0tmWhd
ZNEVPabQBSjKRU0gI1AwBx3Eh2EJ7wVscGqQfL3LCbdufB0r4gJ9dO152uoFYnv2LrydVI7oY45X
4JdXeo8/r6zH7UOTO139EXnI8JthMC/EINle+GC38BSMrKMfiJl1+6GUM5/uNyssO9Fp+sUlN2l0
GdIW6jjCsLPNMeg4Vb4lKg8ACDxEIW1iOuWlzvn9G/98JC1RKv4rG/rhHuAVNRyVS9G2RLpxV/Ws
R5bNzNt+PMhRoLmwbj+Cpbikg9qSZR9vlJFeZCduhjF2Fguj40Q6kMzQagv7tTb4ik4sfrkORlCw
PPUuV53NahDHWSJ4HW3wZ+j+znVy+Ujy1+zqiMevVtNqC71Hyl2qKm7OLEwJpDGwATt18yfyVxCR
TQQD6/kxoVa9NltrrEk7qPdI6jUgSETYWYF3WVh5bSd5L2mJF5g9stS/SgaZ2aI+X14CPetxLo5r
OTfjDn9pRBqKIvC3VEOc4z061Te3S6SxYS0Orp0AYfeSTV66my1U367BU59Y5/BP5VvmDqkPaKt3
a5xKquYsjIO4OOvKX2fWPHTrAWQVo7g4Ad5GvaE5wbuQ8SeP4UXKy3fCM0RPzKjAA6MIT5c8p1Cy
0920K1iiz23lAGQTSE7LFPdT/i0IEc/04l55e83OSLOjMw72e4HT7YUDUM/XFufWG4aHyW2F9fwN
1MLWjB30D44CmI02A/+/Do5zOcioBq7wWha3fhavn3mxuQL3zjIHV8qSaxVPL6Ne+tZIHCJ3W0RP
0qZkDtAceb3TWoneI68hQ/jFriR8cHpfVTbAxxoawe3zj5JtzoNiSQ66tCfFaUVS24fIX0v8ypdg
aAPJ6bLHa8fUvD0fX6hNgp6uZ6hmMN6suwQNsRFDdgzaPMwUIB4RKrtPhUWg1N2eOud5e7jirutw
/bJv2l7J/T+NhWfqtANbldZX4bsWM2P0SeEj6mG0GjUT874TA7m2yH1l8195ngB/NDE3YZ/2YFDy
hEcQZamzLsdcGPpXv3W87kYXEHn7gikSST2Ims4Vd3/BHZPiIyyRiWyzLL0aV7YxOtzMSWMwJ7HB
O5tL1znlj4+zXhMFUhv4ICSLahjsCP/5AaeOlL7tSGteWfPVLMCgL5vym9+3f3TY0Xu3T6/MB6sI
MWVVzPS5nUxqyjfIddmPbnucwTN8ZeiUMH9l69kY/zCf5jkiYgsVc+v/PYYDvFNW62atl+OwGJPN
SHO5ZQG+aFvb0ex3WcLDcyAQ2UjkkByqXG3YmKOWIsH0oYqOB/i5lKpWVFum00yUIrLsaxQl4Uf3
5hqasr1KMtWPkM8XvG3Yk+7d6/gRkp0jidU9VyKaBod2+dF5CYPZ7W3xmdT1qA7ES3WZpcsmozOp
lwlyu12sEwuP8gJgewbEzpgmsnh6jY2PxoNYRLZanDo4x74z2A25g+eXqvPUmPD2g2ttRNEntQuz
J/xf05GGH+fM0e98WXEpPkCkyp1aKSc0Uiw+qTN0oa/i5FWPM0JIdJry0By/1qV+S7NQx0P8Fbzm
8jXNzPUlVHX3ot2wEtpRy5DRK2+pMu4JLaYPVDFRtDknXG6jFjTFoQ3x2ZgkJr3osLDh/eUM1r3/
LJGZIJn8POAsq35UNXIXWxxaIsSEBiffCBiOgHMMwRa8wreBADQQlNuiLkoC/LjreNRCQFxpm3JY
bbGKpTlrAdiIMpiOpW8YlYJ2zpZMG9ty1j9EnRda4MF01DIeSFOzDhpRMEpUROwzXtAjnwxXPGcn
qYQ44zAqf4qSXPIaM5mQXXn0cVPdAKGJI6jcUnH6GkPJd0rf2WOeXwI7p1SbBFgVQca5i6uYTFYk
4LkAmYzm4di4IAvQeg8adoV+PxrtcySfs0rLfDZlXhQqqW1+c3XJMkmksHWHBKxr8hc1yz11zYD/
1m1q02+0Oh88W9nRdwDJNUYMnZO2lpeM+TGafqDEsdSiZsIjkha0b+74gASzH0YaBynqgL3xLqw/
ZCELp7qxOQCsZ1SAuJhqGMLyJiYjWDgopKBEuOiM2Yg1kJRY+c/jRItHsJftSPi+C6k1aDSUhVnC
qWNbeRafvc+PGmlVT67GgkAvTChccY+0+yJPDpm8A8vpBoQ752oEO8USy18pKtAx+wfZtFtlMU3Z
9Bq2EyD2Nzgva9lUVbYSs5qmOF1/cpqn2GDhopxF25fn5dsiVP4LGwkrenzRW5gaX0bz9bsWpzOf
O8K4bxBTsWiJSU2+GR7sPf5qOXnm2dmP9fT/U95iR1rhj5vN2Bpz9mvlCJRDvwRWzg4+0s5vUEU7
L+Mr4Co6sBxUtNh5wBJTQs/4raVCvakVtIECkEZUC0gzFQs1Xw8wzHeN/m3Z7gPL+Won3tuaKRc4
MpvfNKyDdAsuvafhgK8N3EhTPWbMC8xVFu4nTcOkZNlqibeIW7f6SkxW0Bv/rYw0fj4reiF9iL+e
8Yx+gzFCPA1uCXYPDtJV/HlLv6Mensqa4/dGxBvTfSZDOIYCuNZRjSPZPx1ocSt1FmFhK4vqQsgL
MuhPkC5RZ9FhdvWH6ardKCbN4yhddBOgRHDLfDS3SOF4XzNryF+NHrbvP9tQB067Tw4WQ5X7d7Ji
6xepnUux1tEZ77Tw3K6NAQeFqfFRtju7nS0uEFHRKMm1tYCPgouW5GfxzrM0B09EUBJaYaj49/Zu
rv8qfx0RS/da7eimZULGpwJ9i+76UOY/fIUX1vmHhNAHoEH7K2EtsVLG6Mm4GdHJBK7bZ1D/y8vr
IRgq3xS2RdO8WbOkx6BlBo4vTQp2PAarCoM1ePYHP3LEyi5EomrX9oghJ0JotfKEc9t2xK+WVCRR
uR9osQhIbcv5jfyGnxeqlk3P+hII+vMPVb0bptjlD9ZIuT0j99QaKFBffkrwL5i1rjHMt3XPhx+I
VFqpTKQZTbyrGVI7UGkDkVXH9x+TJ1gUAnRpdJqoBk1Ui8atBm6CC0pDqJ7A73LS1TDbdkS/pMmC
xKQa0Evze8CRGS7XQ41HUX8ig1wEhzWf3Tcxo75si3F9M0Z4a9+uACqXf2jLewyanC5nw2oQWBDD
LLlcorSMTifJhGHybIFuRgmH7vpUR8XyIyVF2aGnEs0Rgv33oyBt8CqyTn0W90BsMpKLoZvKon75
byqGiSWDioP90vw/f8E4DkA245aZK3TuNe6KoRlhGYssnY3YP5tjgCQ02dzbGhMrcu3IPVdWVVkX
tHPoMdQKI7A/+ZzIdSfrViC2oaev1WH4U1RiR/PXdd4gs2a289X2vlBH7owOyteOmVNOrw9Rd4Kj
llLFojlWmcS1Cg7bL2/7ehXqKUr+M1t2dtQOBIaI5yX5OR9qQO2QLtPspbsJEthSZmYXNY0PIOL3
zS/7fDBjV5ln9jJ1jLSE0ZylI2nXhHLKgCwponrn6UqS8q545n/a/6Q6Vti/pJqMhoMpMDnCr5gw
EK5+dHMRvtg71p59hsebjnWXPA0xd1YLDZrHKeXlRqD+KnC59amn6d/9Fyy+8ayDCwhQ45oUlPg6
QDlUiyyM/lVHlRSYVRSF4LWG6mSgMGEYeE2yIeEZuTzFgCfQNeA8ISSphdkz8B/tNrDu5VAU62wr
NgPnbunvBE9/XHVYI7b9/wiY1o54dJ9eUmNRA4yqERTVLp0LPoIgY0AZMYqoxt2WZtv0YJ6IuDdT
tzCuHH14eHKDFQOYYTKSogs3bZiQXjSozaGjWeej47aDlKVyG/o515lQ+VTJcVP0JPCt/6cyxyKQ
2aPgPS1uRostsbKkd7FeIDGoPHx+MrYXt8hvPbDEQvjKmKDwfl3CDReLASZTHj+mme41/ey8OGTD
OvcDpr9dlgFBwA+fBBYoYKBgyVFnGGGWM2LYxsluydiA3Q0pIAisJ60TiOKjtCEX/jP/ftqQLbgj
Gq+F3ZY/NrJRYImeXSjX8oma5z+Qrv15pLztfu4O89pfrRj/2IB24o1U+XS0XXv8puQif3wsrGl4
jhvdMkn4MYALOua/SIbWBsWnvEIIJEB7gYMrssvsLpLji99dIWAoY77xewFflIEToMM7J/09Hddg
pq6DVzMmy4TFjlYcLOOjIcmv9gmoBXjGtTR82NAZ4OX4zz2TOiFf8MC5B2Mwb8zK1Zu8YTEfwagN
wV+FizlvVVxePKv7kHZeanfncwd+6Y0AIcx/HYfpl2u7DdhSRjkyRCmZtlVFm97llnp3YKDN3GNw
DC0J02i/5aYukxKB/TBaqUiZn6JEwsBYvyBElZnRH+vsw6afTS1p+XI6xxFFhnWJIUGAJOO9jswO
lYFr5mxB6rN9847QGpdQCabGlL/0OvVsyfZawuf5GT9uPMjoDrIJ7KGYtXiTZDp+aIRKPlXjPA+X
BMMZjl/4VTi3/JUAc5llkLrKGFf2Tv5ZyFJsFpXrzexj0QnyxMWrfX8/DGcYsjbY43WpA1u4b7vk
OsQybNcO+t5lmfjebVZs5zxn4rwSwqZeWYP++YDPegYIy0uE+8Hpxu1sF9ZC6vjAqb5HKmmv0DJ3
yuMUqrHyeBQpq8+gNsHzB21fKfVAtCmW9412+JJpi2iWEXt1ienx16JHk5hbH6ERhvYx2nNuSYxo
PRGffzXym3Klx0Oix0dsgmhYf3TOxmttJhYzK9AMpwBhw6JC3/ApoOt+PisqDNk2sZtRp4ZtoHkU
XXLaJZMjw5tyep8lmlUNPJBL0GkVbNtUN+LoJtqEET8GeNNRVOJfwV9HDPrsoe3iENXw8b0XfBMz
1Wt3FlFJEH2tkZXBpCYwcvkThHtdbnnXy8Nk5x3bGi+iUaIaJVp6xTFAdJU5K6FLrmaOxva0nI9u
JuRsEZ1oDWepx7vQiJ+hMIOR0gouvPK3c3vPBXqipyT4sl/31H+BuxvegZtXYDmlzsTlLBaBLL9w
0rQNBaNU9GR7BWFvEgx0ME8Uc0F5AVXuBTY2ha1bDrHZ19c8RR9OulUAa15YGT7+R7RrAnoolLQ/
WubEDClmMtuQJCir9jxX52vhobbCFAvXycfn3eN2HwrC7Ag7vWlpNrMU47adeWYwxV9mWqfJ5we8
xGGMX1lwykv0sOLIQwCy5QMSNi+Xk2cJ2L1yC4ImSqpMCaQs43BQ5ywyJ5AKx7sXQy+W6Im3vP40
4p3gjBAVZ5EdY2KbX7uwR1drqeh1C3rEVa0PMMyOVEBpUo2Zq9pZ3AL1D/Acozy62sPMCDOTA+gS
XlYlN89GKRVgM6tcFO6ObLRPZTZASgZjQbswcP2hIlimd3LeHPUCiO40e/gCkx2L7D1f+hhJa7Bj
qGoC18PHwPnrvuTZYG+QAqQvlP9GHSc8pD7RXxPQZcYavDunDxk/bnxzH4WSxUbzO0xLq083Ua/Q
kSJ+iNYOgJmCQcPtSTrLn43lQLPxhzj4VjvhjVJlLE5VLzYFYux/EtwYg0Sw4ke0zpMpwq7cS58e
TQ3xMKKZ7z5GKB0MO5OWzBmkOugW8MfGwpPSyH0+YuSsmubcHSa9WwA/BruqxNwQyG0iUV3Ttcyz
LPHKZqe7MUr3CRv+nuI3rIDY13GVK/CDuxxmB6yxgSGkLZSDt07dsxMKma6CIZD1Nui693tErtRO
fpxfxcGQZ6ihWfCS4iy6vb2JSUPj1N24cYpLESj2xYsLCdMWeMum9VMqlQpi7Qo+r2Kg4TPzJ8MS
02p3BLTC9VGp4b0Nnzszjq2lL5VxG80ef2YulZCF2OerctUp+jpzpppZ3Ov+At0Mkf0LIPYKL3wl
Ch8GVzhsu8Afb25+GjjQbKokAjFvjyM61pjGu/tMHPyfs67WP1zEEUJIZMW20uk1dfg6ZJFaneJ1
0i+xraH+BrZASh7wME7X5KueMTIMB/5TtXKZplMwG4OCgQDTBEUvEwp6PaXaR3pz57DxoLVwePMW
x8xUb3GT2hJhJf6LMdUOuhiNd+kW8k5C+D7x+EcpHGeJXRo/NAfT9/Asl4WdU0f9/0udjTj9DUE2
8DuN9yxRVRAZjHbrFtzpB9HpI2M1e174tB591P2sTekLvD0v0N8NGWLlKvp9vm9wl+I5Rraibi+8
Wk/p28kILI1+26/WA0EhZ/cdtJKnRZB9+noFp2PhldUfUAxoK+YAWmlLkQb+v8REmtIvgSEfY/4k
Q8zYSvCk4oFMAva8XbL+pfzB4hHKF3G99U6cPtvEROKsLDyXpYTaOQ3+De5f5SaUSZxd/dM3csCJ
tH+rckpEvcp2tGaAv16cNerIHKZ5ICPYsqDWh/0O5X3x8fYLqApExd/IbmXRU7ypynQt6C/AjvBt
RjgZ4zmdXXpHP/xf90YSaPvGdws5cTaxubT9C7g/qXxTEgI5v1l1hsG0bPLiTGAy4SLIclctys/v
6N3ZHCg6f0LEuSeeBPZov5UFMRpln0ANM24LTUnsNfdicU41MguZv7kVPYFg3jXl3eol/FT+gKxb
EKf+AdtSEIBOQoH4RWxI1P2+kQdxq0X1R+otaw9IMkFls6CboX+ACPR4FU5P/IjsPqXB3rIeqxHj
ag5GAl8c1kKM0f9fTGTV0qsSg66iM/gTXvunO1rCgEXBJRrnVmpFQ5sZUM9OzClt0mSZkJ3x02ei
SWg+pyYOwOQzdc8b9vUeKA7VmIqh2nUtvXwlfRQx12sgPZbfMqm7nunoS0BPpbpXbtSoPxowtcei
gjhZh1PvJ0LOuOHSlLa7aDej7HIZkbQKpicntnF87hsvHvWdrEhcbJSNPEvf+DQXSS6fv4nUcTwT
WehuRp7McOfncAcEgfV5yoDgQU75mEWMOj9HbW6ufn97Rr2fTFr8jhetbRGgslNa1DYZD1RY5Kgh
R3sMhIhIwF02/GB2LKRdlWqXXTbxtXrZmVH5ODP0+Y/qd8CMaS8GTr0Vijcnt9N5gQ20v9O68+90
lEywfIXTrKzCmwgW0JCL7GXJa7vuNk/dyV9VYU5DXQpjGy1eZkPYCF8k6KBc6ZPZT+DfenMoXAbb
PlQvqKhHcyniJZSk5vx36I3sW6YeOO40hXxpHWIwnvgFfx8lqcsBHYfFeh7AkcjCb0XpkyDPnbN/
7vdk9AUJsLzqccyeZZ7JaFKZ1rIdIZ4Lvv1xqq+a1PlDxhn8nGENR+OAYlzM+M3LgevvuXuHZDg7
2KoQndqoSCr+Kc1PheNORr4WN9bCMhcR2Iynn0n2+I3MB5XXOlP0nE26dfb2DAwxwYItWOJtdD9U
hKj+qonfcKN7bNjPR0Sr1MqYit/zW8z2/9XdDIm/xlP1gmRH7Ysfagv7s00Q7pKAdKHiy/rlaCnK
B5qkVxS/ny7iyLt/HhCWRa+FQLSwWPpWpZVOu2RU/A3D6FWMUV2HYYiaxnaA7GryYZpZQIR7TCky
kVlCk3RQElVtaK0ZAOIIBPUqEurAro897wFHulCB1QgYONaFTc27zbxnUuEE+UGn1l7b4209AAcK
Xd7IV8mJurXHDLvBuw4c9RbdiCG1H7i+0UVS3hrWk5mysD8OnXcZHI9yz158Of2bDI3lc0W2VnnP
6mR7iVJlDPq64MoCyKqKeLeL1MS0Z0Jex3v12NDI53SxzBpWWJ/SJTOEJnqj2tVRfo7QiyGOJKz2
IDxC00eC4slCBWbh0n9ldh3gHQKssSXiQCi+Km/ebmyjSb+WoFzri/Z7JnF2VsAPf/xmO60lv9Um
1bch3uRKV3UQ+CSJJjcmiOUVevEFQ00Cg601F1HaiEpOyTZ0ZSceh+2tlnQS7WAETl2bxAdCifNR
ng9z/XJNpUP2IgdJ3DYQuljjw9yI8UGbPPEHOioztbE3j8RM2lU6Q+eId8My95xnRQJ0tXPu9eSa
SoQ9TWt/coCcQpIJkMVq9xiPqEQHLzFvbubT+99LSCVDeVTY6yMi4Zps3vbMKSLJgTzd5ISMB1yV
WbrXdVpnh9WSwB2C4GsXyHrQfdp8BS63UOJrlhCb+UiwyFH+cJ7BFdvyH+G6lB7GTFDOvRbudPN0
fH1zMzik6jJMLpsZYp7D/jQq/CBpeFHg2C1UusXHt0wABcbWO2f8Aanyja2UOY6SjQNGrGF5mY+X
fpp3i4bCjBmuuV1aKO0odLnrjKyS61WuK1EVYLEHXgj/Fs92xMmzv1rpnR43F69YTvOv5hf3dnsD
JCIlkppmjWxOtzsEcxFDV9Y6lies6nCT/kePZn7wMg9FkfD56y4/trj5ylIyPEltW1uCrp2zSHH1
o93oNFiaOWsqt549hafViQWaZ+U/q1ASr/0G6bSFVquUjE8iB4V0G24HSNoi7edJBYePBn4nsZTu
cj4rc82mU0b8EQZY/krZhJiu1qrUXbv9vTkjpCPDedSJZQI766vcG6cuQufhXou/2L1WLtaeNL6J
9bVrpB7MDrqyKeJjyuP8hsKuIEVYRdNajvjVN8P6ZsR0lh3HRCHMqySNKlecs7bgcvMoPzVDZQBr
fIu5KGXGX8UFBxMFjdIeOb8QOeCslihWGzXCIyxNVRcOGLATVdWpO3UpGvZMZ2dfFOuq+Psuoit+
rSh/gM2jSKC8nzQoCgtloFlhLYlZFWgtcIF+DX2tQox0OKBJyYsCk51WUnqgvfrpBYUL1HTqr62A
Bt2ExkZ0Y3GLsLNLTLfVy61hrj0sujexOXjvWYhwYJYbo3g3n8vKZHBiaqNgzJHtFMIKgyLboQKV
lNga7y09VyPJkPEWmETWrgoC1+naEjenE/p+QC6tm7qO96I3yuJYylcMtU1uU1pQd6d1nU5Ll8dC
Ptn/eLz+JUV5HBEUH1sQpHxxTkL0BBQH/72IbuLhjXp3y3rCCAHt2bNTUXtxQpK9kOK2xvYspJSZ
F9cKJFoEneHfHNEIZY/UHEOQ/ZNpWj1GOWdguPiEj/SKnG3ceOx5MHMKW1KA4w8qOZtfAmLMdvyG
VzMAnviLiMeh1uI2j94b1yPlKn0QJET8PFFMsEqCN+/xRhkheE2l9yAPvIrzCVMRAaMagMigoOKO
f6echi8XCHfPvnDd/LQTFwNWPrHxb0PlfapsykGAssnu06WyZ+RqnA0kPrhJP6AH+lFF1NP1TiWY
6i5vfeKoJQQgT1Y+zhNyehB2aosZRek8AQ0RAVpVd0pHEvd34q/GW5WlrXAPBp1PsjkOy8ueibmP
afzS1EXOu4eBfjoxJegCYKIqm8r/9oN2mxNhg9Yd81Yj3E/uqPX6DIm0Yd4MoEv0DeFs9MgiqQeK
0K2I0U7YhsOboAfCfaX9mK131QYcxGtql4siaq9n7MFPS3tSAngDrVdCNqpVlhvqCdPSgFE8ohrP
1GAXxvNNs0LrNsm1ssQbCDKpAkG20DIKYD8ll3wk/F4ora1WE6rhU35xvZM07m2Q3Fy/JL3YAZwJ
Q5pEqLtnN7pB3+Vxs5Fjvf+RfFk6MC/EBXd+1wng/ub2684QCeuXL1lSOm87D2zsJ/2CruxxxdoZ
Y707iTYDRRqnA9yjPSJSv0sNTBbH6VRdQlyuuZLmVKaO7IH0RpXCYtrZ+kJqHC5SeADc32d0DOXG
PCL6j9G0hp8v7vWkEHIgdCx0BYXs4H3cPnPLVCPDfEkCMN8dJ8WY9aXpvugVvPQLH3WVJKa0waPi
IvT9w6oQE4csa9L3yYGqqQI6nnb7P5MZOyMXifO+VoBqUHmT1+BunFR7eWA6bmolqEX0Slp0bxe3
KO1AKlVsBs3+RIQWBWJlpgipV+t9JCAaMgq/zvG0v7MqE7w8fDWKAF+EuGqcyaLC+IOR0wORxUuQ
l/ja4EqG2eqluCIqDvYiHH+rB6yJpB2XJWJwfR3memeIfxbjB7G3MtCXk/77/7UMzDO3+z6DcR3A
uB3OarPDOgn8K+HnP2Lh/gbhDttIl78N64QEcB0P75TxZw3Bnrz/z2fGe34urGiB7nTw1NDfqd8G
KVuwA7vQXzSWSAMlLE9lNhOdpDmp0rShw++iERG3LXmMkyVA4qC+3WrC7PlnAlkD9w/fMmVCc8e3
lPRl7MvGjBQ1ot1LILw3ycku8rKqSRyj7X4uFJ/8iBMEVHV/dYt7/8jGWgW0NWp3147QLOvh1L6C
u9CxZBdO0to/di1fjHCbfnrrNcOM9ExIKY8C9gIoZvu8hREpL1AIYLi6jQMvfMdTaej4x1plmnCI
Ln4cynGe79P1+mfi+j09HWoSwdkw2ggVHIRP+gsim1Rul9kSo65xtwS0cyOuAFz+jZEFyli2dn8G
bISdbYLJqlBZqO3iqMcvPK1KvEZjOXhnTSg6jCeo4bxmn+OtasAw0zl+lkw2QEAd92PP3RVsSHoY
3OEr+7q3SrkCqsVQKEMVwQ8PbtVPKZmER2NwJUozxyEe9Q45o38sNJ1MZVjgYGpMm1OnysgwlSoX
PLc6SQTPSQqfXHsOJzrcFJWX/a3Ifb9B2fFFP3gr54I/VlPvvzWZN4Y5BMdw/QKMxTpnG/PzHnmT
9/ZV0qNMY1NUly7XDBNG7mFbgGhNzeflwFGejHT0ROKu79AB5tps75fpDkTIfQKnW/NNd0CVmSld
ws09Bv8516lCORqIzPXniEl398MqWagSb8KL4wpeNaOGcWrFc78mJsxxNV2Qfyn6KbYsUUF5X9Q1
TQXjKlyDexgRvlDD8P10p2m4/IZKcplY6Im2oO7Do9Lrff5+LSeDaZ3lAEDNk74a60Z/BDcS50+p
KjmQlQW0IoN3UdOle68v8t7rsYiFqbLld3MwJYEwX42c/QcbncCyaqsQnouvIDlPXdzawuU6+F0D
d84S9P0HIoVWwra79QBSZObonkHvKQ283FUazVuuxHB4Pm3vpM2BnH9WvY+l+zcLvooakHTDNUdW
GNSmJkzRtctDoT2FYyO00MWwAn26fdTUQaGn5RfHCUngou5B1PPnr4idR0zgqJOnIERWXGa8Wgzz
+7vhdWtl/DszTsQqnv2rrokigXX+so6PA2KXcLMlVxXjZQiDRcIqxFYR0fRaQ8S6TbVVxCfG65Qa
7lWrGsFoZjOoEw+AZZ/RHoS2xM4gTzLMOnrWkssCxqlrgBmBfBNPMtYGlCXiF1GZu6Kwm74yYHf6
Nn9yrOwxykItHHY4N6t8Nl5YFpwzOCGqkawHyl7wqcnNsLnvF5UPGj2caMNehVBQy3PpJ1iTHkz7
yCrdXoIllgSWyJGfqVt41QF3LK/fW11H/mEXSL8U3LLa8FBDtkQVeRwm4kjZswY91MIpR9GWP0He
HYKZ4bMLgmNPsuthyK7fCQA6ekWxxv/YcQaBKfG2fUvKclpmNTGwZkTqfOQiLSTmCoLoVnXL4qTU
vb80bQl5xL4JG2qNhbW1nM6Zr15KKRbfTbqxqC/3wBaV6cCNUJNRbwb420GLlCJE6an42SsT4d70
qnoK7MaCUh+qcZgvAhjcyVHJ49ZPm00L6VV/LezqFXhQVYp3NgknvGzfGQQw3g1K6KeyH8AZKCwl
pTr/74+rsFSgbH888hVXK7db6RD9AQ0Q9BRnpzv3LHyo1UeRQ9DK3KPt9wBWP2kOjHy+fE+eMHul
P7BeZM8zM/cvHAGE+AVrmT2w690k0fPOZzs4XnuOCYzlZVxH3bOtL56EOxRuStf9/lcNK9N9/B7m
pfLYW6MaMZVJN7IdNIanXIDGLPZ/VgDrKj3+blmsA+y0iuo96UdGzzVAVGssgoI4jauYrr1HKMuj
0/IGOi+v6ZLilsZlYtQWeTgcO6/SZfVhkQRMNChj/Y3ovJBqPId7yRDUz7c7qVZRPINjdI5dWsVl
5FCUdnAFM+61L/ufEJF5c/u1ieyalkep7M27jg21gblbiBtUlmghhZ9OMK1NcGBANZXBH626gwIW
/Mye9LcUIyE26OIzde97HBlS4A5JuJ8wxnXHgDsIvzA/ZrwaQ1AvabgsXQ3j1H5Nf7O1h6mtBBfH
nalyDd+fqSAR9VQHFhwCMVmd2CqgYmj5ctB5z96S+yzgnT6i3onteKJD8adExnzce2WNgyox9ffu
bElXdOk/1gWjggC9du7x3CHcE2xtknXxoPpB08hqQ6paYg8gWqNrR0fWpcZVGVpXcytC4iRKsq0T
Wa93llvIIr6CL9uIG5smbYbgVMonmxAJALlboC2MwmNmyYWPJ0tHscY153eDu8H+1pl2lIKbD1AM
idjuohhmAZ8PEQGllzKuzmV1ytbVXMlXIraujvswhHypNW7TRuzIrAmJMK2uRohEo3Tqu7yKrU3L
z8SLHAgpW4P7Gihr+j48uuX9wtduvnYX6+/rjgW/gmzDfm7IOP2ILGi2ZZ97/pIUvAQav2WWMA27
uOSfvmZjyv9e8+TUlPIAv8VYlE3A6Bfljd/lJpZa7NqmMKBTVqyn2+EYOIrRAWH8XiF7xhVIHYjq
lVp0gOdvIsUFajvOVGYKH+OUX8Z5Mjad1lKZXgbSvUwE4X/B13PMcMFZr62wVsk0YZg58JfPswqb
CXTj25wuoY7EzWJq2ozWUOUxBZj3cZvNuUPkGE7igsdSJ31PabXywN0CsJa6+9NkOhzUT3Uu2oNT
2sLzYCdLUt8RljFIxSDTtmtaSGcbN5uFN8c5UEgk+exEl1puTWKzRqDmgAvajBn0CQ3zYDRYxeMX
2TABcBhnV/o/69nA5umIOWnCiRlqVhcisWcX813qQZkhhVWns0QbxK1y2DX1fW3e4a+tjEGvpx7l
ovB6rX13bL6FqDUrjDkVv1cnBt2owNKgt0Jdk/xa6zPaI2uditaLQTZ9S/NThZcrgkQaBXA3qmKO
0ik5jAXmhSKJkkyfRui7bJD2kjTmFuVQZXkAK6JSt87i22nWWvLnwSaG/qBH/WUolNwaVklwx99L
w+W2Bdqk3uOvyZHy0gzQR1eIsK3dXv2TGlUW4/bmz8elgeopDhUcZY1PG1x+Zrh8KOAHsj3S9vIv
U4hZp4P6Lc8+J8AsemeF1BsU6WyoWo9OMMEcKltnOQnns329NLW6exudmxQ1Uazyc6rWG1nN4TNx
jnXbj7F+QSTYLoHVBvVw1AUQyC8QZjzy6D6vwfIQJIEl32KFmF2WiMhdwK5pVZ1wq8vXAlDl0xbE
LsZe+oRlf9YRccgD6UQQBQxEyz7sXyvTYiEKPjyaSxi3eEaHzvu17AgVAMOcmvcu1tKOL9TjHXcM
uJxO/qmfIpfuedkQ57Bo8KF5cwjtL6h1tqdP7/00RYMXfZw4c9qRgoNmWXfYvPNP3YQWuPe8nVVh
7RDQJajqR3eav1zRCzvL1m23R+jb5SucdMUE6loTrJtxHHLpHETMLCdrIyuIUSwg8LmZyvvsrVIs
L9c+JgNS5VUEsItPlHzWQv3XXfr2TLn8RUavu+wFezfM2kSJ1b4tQRxvmJcdfmhoECqZ8+tr/dZR
mxKxmMGtHP7Uq6W1/vxFnh5dN3NTgPTfHwdS/TYfCTlGdaJvH5R2XCqdT0WHUWTVZhXJUCZbwNKv
7W07GdjbRxE0W/LDwaGAD+8ZZlkh+9+jN24O5dMhO8fP1aV5b8YgwdntJ5NcGKl8+UhaaSCto6Lh
7+Cpo2Xj9FGR0nLJ0x6KvglA8RdP7ded0gw+enXmdki5eDAl5hIAHq9Ktf/vkgjVD/HxdyRawvso
Qpd7WGUZ4c6Az02D2bP337FbfD1SByyFWnaxynfhdHhowOa/viHaf49FlvSBIZIzm+L3PQ/Uugbc
xlU3COGBZgEPx3uFfSJ7KznxT9tWKMmD8V4zFLI1RcwMjjtcuzKJlHas2LqbBkqukauOQifqgb6r
QsFHip3elDKXjMRD0HyecZQC9z6ZMMGnhMJgKEXmB/dnlB0q/7JR4TTEnzYRjeZOJWMKDIHnIt9d
SyhLwbhpMETs3txclJ8WqLuJdxXwiF4Qc/PB/XrgZNp16nAkLGEgr9EkYWsx33KwqCx3xNF2A+ND
3Vxbvv1MVjRP+bOK513njs9yfc6tM6Wk2bgkmrptnrrxnmQLeCmg9gt8o5A0BDiBgts1nGqPlq7H
B8Mp3KJ3QCGpvN0nkAwIwulVIdOFyOAK+ciqSpyHUEceTpEyfd4B/gADjZyggOz5QIudX2R5AZgA
xFz0FZP7eaWkW55i6W+5SRykMLhyoSgZA47V/NNtmkjhWnBmxSlkf+qsJOp16AdcPAPCoyMVNoTH
0znllMBQ4eVyYCGUy8d292NM2UUO3Rr4iABgvbXsv6xKrMyFd6s0JMJzQq5JT7N5lGSD0SS0ckcb
3xQEjv7ZHHo2idMhT4NnmP1A6yvpjMqYCbbDwupKBxugfYnY3e++i2BdmLCfCQzgd0UcTjYYxFP5
MVoGMg0ZaM0oZIfszZqpUJSnLQOfNJck7/L5womzrC0yiFbT6JXrFWdAXgjRMmHfbb6r1qkAE5u5
SX9B30W2/ONMEkWyf6cnC+zdpo3+NxnYzipUAwlwZ9Q5El3sksFhfe1KVjZ9zAUZQ7FinU3QRi+A
IvDanrb1Kznj3nTVigDoCWc0vipIFmvLjiyJ8gyenb18TD4hmGCu6Fz2FEmFAMAhADnPfy/+Sq9I
VNodFud4c2CHNNKYW+ffUspcW3Q+iZh6EwJIaQqw5RWVjEdnOJ7UnTlG33flFRb0VYuuWqbTkINh
roQdTHzfixVatv09UtEDsbCy3CCWEfwUB57ItzDDiD1MPuwNPa1ttvwwr7E33+FjhTSjrS6KTYhU
5Goli2FY84D4lkmiCBW3ReK0Qapq9N+c8mSFhq46Yy1ikep1xyl6QcqfqZ2MSqAlL7Q6oNNLTXVy
Ra5w7J2Ry6jRK8c35vafgmk1KxIe8jTZWEwQP4tYONlBFLtvBXJQgjlgRzoCyFmbKYWErBIiUuaU
NpyHlMwDGMb2jTIHCHEYei1ryN1ol6IU5uv+fPe1Z/0cwzVoZnca+QTFZ68NiwHI/v2swqlhPmSW
VnCIFaJRKSMNYcf0AapPZRd56BakZZjqlgrxIYCora6UTGC/evIGOhDVPu2jO/sj5Qkn26W0zpmO
R/VZdnr3B6i+/HlloA5uLbzWDfj0r6ZB/dba/Zkr6+L00OW8dXgzxmvLRe/6lpLnHbhS5NeRb7uv
lhZAUCPlUvz8gO1tY59dvAt92ZiXbEYth3IS2cZDn5wRwvEn88OZUFkcYlSSSMotitO9vN++MtQB
QtZdkSGFlPpRwIMM55GYZLVId9/eLudsPhk0hX6/SuxAjwgJAqOupidNXNXwybxIN+Tv79WkbhRn
rKfXNZDJ0jRiqqYOgBLO4SUaG99/yJwAyZiLP9dl0aV4IG2KkfAZRMKOG7NTI21/v3rTPaNBxKzx
yQ7JRWbpEbLR/hzsmQAuEI/OteaTGJz4RFTmxT5y/TEymOR1fiiws6lGg9/qGvlIPqW47x18OETh
9Kn0Hohpr6jnEYfyyY0LZF9KI84idpLEfNwA26Rsayi9nlx5u6n3SqK5udDX5FYXNC5rRgmL+IHi
Ab4OuhDtLLMIWlgzk4n5B9835t02+dn7Vm6Cmoj6OPaqZC4gwCELiIVYuvZ1k0qo+xx/VwGz5mSN
xt8Se844jxHPFwH8xvJztB9w0n67Kx62SkpFi6K1iCWsdfIXwzHZpBjSY0sQNMuORDIXeF8pvvQe
3rv+wizLCuG1FassYnlSF8AahkiAx4RdmyxGJAi2M+sO11j/QkIF6YbeGdICpKYigJQizZQL4VuX
GDzXTCCDFr6w5evm33uagBi2NnQdCUEg4s1s4+9bJs5pfVxUTHsqFZtgc/pd6moB/yu5xdmYgLYG
TmIp+3sOg6ZK2/xGyHVprqN27JHiedou4YARmWf6orKMZzv+jqwJMNp+Kg1Q91FUqk4y7OO2BEAv
veZBSYuTF1dirB4lXMWlXpd7Ed05fQS6J0sCXCLqCBqEob7ouiIVKkfDLxAnVrfOIe5+G9ewcicG
03aSAfvCuJUBUF7WGY0IDdLoqJO/B3WLzkXmZ0qxip9pPJuKgns/u+NXLIxb8swPov2kVmHnE3T+
UBlL2keQsJtvkCrsnWsyvdRCg5rCeI8p0HA6QuXGhT5mSSNj76J6zLKKG0Yz8zAspHllMtAFTEWy
tHjIMg1jaQ0OSN9DC1YCA8/p6NtAxMK8J8kAS8emjO29ho3rGeXRMlSPMK6N7qIiBZ9LpjuMdRVj
VocOTWlEH+iG7Zy6rhrtkMaEca6EhzWBupcI1YYy+KQZmsoMKl0rJVSX+klZZ6jqvO5VIs9FdmvN
NaGvosBVxgkyujNvMSKTOLKLqkytzT6upvDbheP2iKpKVg9U8759M0BuyuvFB86kDIrWhgkpnQ3w
1AF7VeWx14urTD6SmjObkGOMybPJd4qnsjV4I82wVG6oATWWKi4zTI0XzhX+y4e3jxWFHYwaD+fD
8BqORYXqiX3On7EE7YYylN6r2/rLdXrkU1ZXf9bNgll3QpguCRz/u+eRqJSXdLicUvg7JcftM9GG
D7DE3FLI+WdVO0pQgXuwsaFDjb+cyHgr5ez+Tv1dmH675ZyxiTTFDSaJbA7Jp8Yy1OJPPgbs4bSa
CUEgGJDH1k7W4PXgOkmI8/K8djBBZDqFcDsBXV0oLyrQx7eIVHi8iW4oIvlEgqK7YEmJfEdyQCVv
8wMcg2HY98RdWgltUn138SOjgpbJN9UHfBxgHk8qJ/vAtqUcUoX6E+vLG4+erwcCpMHdtGBqf2GW
TeNTspBjxot6YnR3HzhGCBLWghL7HINKj4Fo36bp5qYLChv/+gZEe/C4Jbs2cnlvjAmeknUYe9a7
wpo5yZ+g/A16RSsiLG0IiWzfAqXjdzed6G2pFD345R/CSoaXqGAC5PcAlIjVWaajHRec5KZDW+12
Rk+bVPCOZoK33GPCIDnhI3fDERc8m8Hh2y6CFwZ6rmqtLECAbFuq0tDyIt2OnRmquFHqklaV0zwb
n3WLw65cHhfp6aEZSE16tpFe784S5pRoLTti4XgWpMRwvAUgBLOeKOorapvVMgHnnJ4LhH6onrOY
mxeEmB+zPX5Xnv9H1J78sLbMyiNI8To7K3b/qKB+K+FcT/U+RrfNKdMoCyRAH4omJ3WvTJO22f5q
6HCssKsGU9YVtNQuQjVw/JUlftg2fggFqMcVie6rBBZz597f7gwkSheYLMKrPUYaZy6C8fldnH2a
zVXFxGfQIIvcCsxP6yGOCgtpCFzsdLYz7x0USnGg1UASuA9V7vRHYHa3ZUGp2Etio94gPbohLmNW
RkLduzaOjjglNtOe9FrZogocmSDFlBTQDwHLY2VdqEwCOdRohGCGss7C1S9dsGUZZGlgzB4u/hzU
CorV4BwGrHQz2lf1lmjY4fD1hkCycRWmXa715/J03QhcQ1Db5C2ad0TChpHmb9V02H2ze6whrA8i
jGD08BhHTnEXuzdDleT4mXV894HbzetIfhO0La1ZAUm6lr5UdBydIK2cQq1dSO05ZDk4BU7TgzCv
riH2EkdmKJs0ItzW9vKdiB8hgf695JB72gl3uv4fKCZJSgD6e2n/WzHEF8Lpztbwc/m7xoxrVR4R
eqVZYWteU9bfUUd9awQjdeL54hLgQCvGhHG3Q/pcE9MOni6W/hmkAMxgjHPUmYZ2cfY2T8VWlyiI
vRYwBnbTyELTeeigyye15FMD9UE5bKDBsJ9MeWepxGsGPBnPxs5LDsF1lgNoyeWBTP43/hwvtWiX
Ukt4RQ2JLQJ26kMtJZbQgj3CMaxgscRH1c65bcg+GiU20a6x8TkoRnW7QK3LjjpNsgi7+fo3L1cP
0xDpTRGXwo2TPrEAyNlHwGYJ51Pnlw9IRpkGf0ZorbDzCbFfS8hcLmpQQ2PMN8Su2drsTvlIC5vU
zdQIpMahXxmFduzWQzUl8DKhKW2iYhQzuZriJPbgjkOdeHA7cF5gqzTGrdsbsFRbCCm0qceC77mH
B8utxtxViXnPIcj5n78iT/reZ3wAGd/zxrmWfp62M6PFh6lVxaTatue1XOQrj2svwxlmnUhIQsHC
qudIYCENVIGbK5aWuRXHf14HU7yCST4KFF7JG8i4ianCBBC8vSRSQdEWGJ/ks8s20/Zz8TZyFBBY
nhd69lM4d7scq/xc1YKjP/5evC1vF55k0Xpa+5Cd0aBOXtXIL2QdeXzqoI+JGXFtrEc2rfQOOn6u
2EOxCYG9wa/EeA3s2G6ly92CSsF3oin0QHSlcnA8sNVZexCB7Cp022IydGi9PoWJTBWnmsqNnhUw
BUo978cEejYqF92+c4jiSDHTpfaw/2NxIAXJ7ehYaHLXQyZ1y9B6Mncy+Xx6pA1yZ2aNG1UxhzsC
IQt8NiDir1ljGPsgaI2haH8VkQPeWsO8EWLq/4zLp+sj5+eOoaiS5gxEUjvQJY0sJ03kBBOLpJvV
J3UMw+ge0q7ylfE+TP64ZcqfLvrU4sniTLjxpbUksHDlF1qllzQ7JSpkhouAzIBpiWbKPdY3k2O3
pyVQPmm6+IiDECge7bX44RNeKUkyYikAPpW9gSRNl9/iuUwJiyyHTey0KiWCr3UbDs5+yx4KyFKl
mvqqVg/VEk/UT/1mqp4/T4fSggPE/SG7/TOd7v3nd5omMppLdfDXPFpIJMJBa8GzefhZJPRlwLQo
mHLxigh7TVhufLGuCejNMhsaci8J2sJ+7Uzei2nRXIx8HWoStn1bPZU7ZXmLQgAFp5tvgbQhcKP5
RHGxXaYJF6Q7QLQbmNaAeEcheuGH5Gg1fgxGwWazh5YRZr5WYXE5vsY1jDa+s/KD5zc0cNvjDi2b
zE9ZYGr3NcmBbJ5G6ujECDEhgQJCnbB1uBAiL5FSwOgm63FMCI6LFNrEP3r2gJNFn0CfAXcSpy9m
a1cSDTWnqFlb8sWzuSqM1PAwjyMtOLB/B2Mua2lSOeAz80fMGD8bUuuMrNGcuhmw4C5Lqr/lrJ1x
+/A9EYe5L2P7JBMUVSmDGK/4vB3F2Aw1GQFdKtri1niVmfOCDDUphmg00AJ1VA369sHvgkNUj6tg
qp0JpcDefOV+ZR0MxqMzhOHoO76MM40snvq0a4qtHa8ZcEnVhuJxaCC5nv1TxkXtwW66bYpLZZj/
96NTpcRbIUN+4IwBEF/VmG2b4bDtwXJhNLW/S7rjQVhwwkcvHh9stwz3UYL0LyH4WBYlg3CQDthj
F+aON/mrCucLOLboIi3o/EuHz930VK7eXTQEgBkneKVV/j3fyXW3KXqp1uFdnVF+8KQjBoQbsCos
J4B37a+ZoHDo65hV8N5m0VUzk44kajH+mxiTu1/cS2R45R5J944G9D21RR7+kwN4QaGR0zdncZcl
O6K21oi650GZBRWvB44ip3Smvm3HKteYOP8XWSG1WMCT3GymG1tiIL3kE5Khwac/MX4hnlimks6Y
S64popzI9F3SS1kpMq8KNOtoCh4sYBmcVzKL4tIGiMb5HcqOap/txusmXFdoGbb216CPAuJSy5v6
fjheoj2ji+Cs/BPCUKhGvpNowGp0/Jq9GXyxx26QynnCaQen1L8wqbHIUU7O9W0ppiSQO9L2uG00
YkrHtJYexngN7cQISfmePKj0bjrbY4OH657KVU5sL132/lA++a7E2RBN/S4u8/RrXOvn7DvbYPDH
I0Pb8q6TxSFbKs+W0HGmKa2rl7bspp52dXzw1IJ1E6DPv+jKH5k9wndkV22jyXwyzlzGRHjTan4R
Ah/vQHknRXCs2l0gqduhJUzNFhTR7QTK78VWHWe4haG2Mo9LD3EaT5pONxjkvYnyTmCMxoOsAqgX
ht4zyopcgBTtTthJRiS821va6Yk8/Col2vQhBnR6H4sOlMxR3uUjzKbi9+1i5mf2AvcSDnjtHQz+
gHW26DpAswBtvE7zui6N58dR3RU7bW+8Bm+SvCwZe1xaAsdAVJ4voUJ7JToSrW9h+lKeUrZviu92
VIs8dv1GDYbYpzLf4+iG1dQIOM+1Xz1IZl/gCuN2HMTq6C+awelXY/R5MWer80IvEaJyeqjV6DFb
qx/83rBdeuZTRgTwuhfuYZEhj/1g/scV6A7VKDGwsyuOcxtWBeITHZ5YziP59Imew2taSOeaBjZj
nCFAW13YzwIUejOi/T1jxMmmy77532G5kW6FwBb53XhQwqF7FqULORzWpNmxo8D7t5wOBcPR7IWo
FNFlSOUm4+0DYH+sw56F8aZ7lEqNh9vp88ePjWaicABpgWh9pXpk4Ws8AyOKee0DqG2/gdFkC4RH
r+SnQXbcKeUXH0WeLndqLn7JPmAc+e5od4yrd6eQeunlCc6qOw6GjLHlEvoM1sM+rZ+K3rVwZhKW
o+6lyP65YAXqg909E+J0cc2yFQlRwW1hWONYM7wguzNb1aMBy2SSEAtzIVsuTkxja/I34CglM1l/
14006CdwMgHFRGlnDOgeg6jHWZAvvTH6rtt/nU6inS0RFyjzdb7gFjXxQPb17Rnmh4hEW5gHaiRz
PIFKCJocGBwEecOxhyzICRdfXXw0l/rPzCPSjHLWa71pgB1yuQ2KOcvX7TidoWxYrlQOo9meLV6D
98p5+3KMYHjmoqXgguNOB1PiflXqp4OJra1Kvd0bf2ADBqnLE25jkzJx+3wbzZDXc4Z0yziyGtdT
WgGK8FUXzMgT4HdBpl4/IBruJ6He+9KJ2Mm6iZZv9KZQJ6u9QU1x4iXBXjcyr9SfvffPLlYjxfvx
LLt/Qyf9RhXhGPX75V6hC0TqMDe/jUQRF96iBfBDZTZaHBt0khRh3KtGgDGp+KVredd5E7Lf3YQf
/6A8fn1+bcYh3tra68xYtum0QW+LAlrIZGqpIJYa6yGN8V+PeQam3TGjPNQW3GCKCPTw4h1NEONF
dFvINQgYNr1Nk1/Dq2ALl9aIY/vvtaomgNXg6+4rnrfLGvzzoS2R/q1/SqUJpr6QZ4zMZ4XEpkPh
uZT94cCpJOaquOEbrCvF3xDwmnTAVk1vrVOQ3YIfZpr0GMoOD3+tl65aFGc1Rj5CHGu/CN0YA5TB
u3SVDGdsObpUyHytFOI8nNl/K1dsofMlcOYt3OI//4E+xPjI4P3NSaXGpftT1zH7D5kkWhdJYO0Z
FAdmVzUbkywcsxh3mMDSKQGahjF8oykr+IeeRwy9Bfhxu98IGfvn31A2TtI3VuE5kuTSJqIiJifo
CEqkH7B/n1EAkwPyLsHqHFgL/1qm2VB5RE9cAp+XGmt2nsTqNi3ejvpoL5QF1xc65P8z8M3SD0JE
lm2GI54BUnX55PP/kxiiQcPgaNGJlGt3bGwkDQYpVSLcsBHlCmJ5JtRT8j1Uo0p2FRhgieDfKHDx
41Qo9adNJfetiXKdTfFKufV0oHt2GskoRVURiofghzfx+nCxBkSh9j+FwNhWY350+Zxyxd+VQvHJ
Vp8dITYdzweigpyNlyn8eVPiDnfsWK+fO0uNrf1gzivDv/8SK3aDC4uQXK/ZulskN0MoZG8xtYHR
nwJOEH4VNt0+XzP3bxCtvteNU7OyYb+yS2XeXcbJgW6hiaWQ6LL0DZHsVwgtRVuuzdNX/iF/x2cg
Mq+3TvsIcwBRlKx4XvlSCaEsKcKShoaPKqNyNbhACPlb5Zb3Op1RY3kLlGrFsmY7443ae4oyuoCO
Zl2L9Hr9vfQCbgX3MGjEKkGrXyfrHvkszCuIJ+aL66IzcgrJeq+2BYNT7TMQMCpPUe0SVvnw74Zn
32hNdgiFVUxQCBl7QrS/WgiPOXPnaaSJaHhAc/+qTLRzkTGr7NwWRoJ3F66GZM7XmkqRL5hYjieZ
UUXCv9E6LKe+etCZ82e3M1aopW85RYkI2QRdTJ5LJ9O1b5cXcXKSuzushexnNMTLeF5Te2YxDvl9
doVRJYkuEwgrN8z9IrU0+i+JDu8OmH0rRkpU8KgGBKYzgvpzc4pmskzMrLTV1hVsYpjzEZqjSC1c
FJs34pgr1aY4F0Yo7fM/91zXjhInj3lfHEvCDBU+ASPlSxY6YdvOM6qSNMkJfK/dZx1iENXsp+l+
lBX8GPpheKACGybTn9l1TyTrrv/b/gjA5KoJCSPMYXp2CKGatMVYrB7Rt6p3vmDoAzeL+pGhMZNH
L6UMG3KWuzGCy07Huaon6reM3P41Xx0vcErZ8ki1e6Bblh0fo48epNIVOfDLLF9Y7NGz7RqhLydd
IzrZw3AKNEPMv1pIB0J4y/y+gz9qsvB36lcyDcsSpxUNqMAnTe7kW1b34grXTAzAx39BhNlKdMPJ
zU3gZYAHoxrPbWlgCtfl6H4z1acxbX5lHZup7mBBaeTu7ijs/xhBpe27pcLOvkmnFT+J3H9B1vJg
gYACmmze68IEjOX703CVSUH1XfPMbVilqY6eTWZbs2EjJb9ydfiWEWBGAxzKkxLHhY2bNrERu43r
ppMfI0QHZrwvLVi1pn5aNtCJa7S8C2sPvlgKYhDVAnrQWXCD9m2brbtbAZ46dHLxH/cfE544NCVL
61MafmlZgrowqfzGCnNqcWd751I/dfHJKfHoMc7yQNyjCccInZJJkd//AtF9YTJvnLgxyh/MnqZX
5Bfp65wW3qAG84p1IF5KuzFGDZ/+txPRHazPoYXS+DfAvet3VrB7l8xph1gBDwjEHL9daiaLSQbr
mB7OGzoUUOGIzHD2IZe25LgiBp5prwW7OTD8cqIyJIOMfB0VIvCePh/GEBbido8ig/NEyN9u0sYb
I6b5aW8IhFokEF3c3v++UjNraGiaqS/BTugvM3Bba3F5mA1ysO80qEtgPwhZDZY3my4p9F8Aac8q
R0V/RebKVVpfouQRUQ7HDKOPhnf9/1Tj4dX7dVyVwZFvSR4GUzCaBMTrsqXalEBUzu2JDYuBpsrx
kp6t1qLOtRwi8X5vaXjFh0gxKOiFk+9EAM9KCITXL/N0EQ4pfEmV/4UWgpBKFAqPIFQ/dmN/9+XG
Yt5QpZcT8NPurGy/PdrHysrGsX24RNMhMZKdXZCXNaZcszYaanY79daxZJuJiEAQsyiLdUgt10oh
BuSFGjpsG5gnk5AS21s3Zz3rmWMuHraayqm5Zsuy0SACUApBRJetkWNrI8q81QORaXihGkRMX7JZ
dTTk7uQIfVtKMoJhXWwuhv1leEISrlxLs60Awd0g0TPMLxfXSHouMI/OCB6GR1PxYyXIW1BswEGe
5mcRrWtBVguSyGApLKWLXcM7+5Pu97sd1m4irQ/p3GYVN3zFzgHXdAAVoDvAOCY/7ACasmZpOjCu
3S7mBWpApZPEtnxDK5Y07k1nU43cUKcwpj4f4ePXrz5b2izvufUGWNPYLM4VoVhYYMAZr9dCFlrD
vL/1N36tlObHNeZ5yScXAaCHGXm6s2JoJIuCwmp3hSB3Yj+LG+G04WtFpax3yujYlfZ4r03emqoD
vJd2lXLh9r2sxFxTGQVWe/pPlFO0u8kK++YCJyUUIGfXvcDs7L12tnGfzgbb1vJzWDsY/KlduB4s
6W+cWwWiHvngQ5PTyJDoG74QYmPaMoVGNaQRc1Sfnaiy9J/7OwaDZRHlBUzKsvyibBir11QJroU4
GrgKmek2ns2tK8uR3K2EZwRZLLDjG4WnfcpNF8AC8oYOhNji1qJoUb3abmymCcbQnFPkaad1g+Hk
6/dg/IcZrs4wb/hq7dA9ZbXZEtXXTQcvc/g8Kqa9ANbnL0pWe4lK3muJklJf9PT/b6LIIQNjD+vM
d8u002g43YD9Jh3KP4eOeXM7HoL94DVBb2MMePqgvCi5Ggz3lpH1lhmkThRGrUCrtnRk78NSxOAD
/VQ3AjkMkE9+xQzjJ7Drrj/c7oUi9lFPlvB2RaAmXeKL4KwnGw2h6ogeNE6DDq7GUtxXmO+DDO9f
FAU3G+rMjb8XZ4jBkCuqeoY+JHNB+MvENqMNjkZA0b2XAA7HRnMOMm8F4ffPDTlXUd6Kgyo9Mqor
l2FeN7cZqwvSvTST6f7OtAvuq8V9pCWfLb9Q9pIxoTHd1qPeempGUEg76Codi2I98o3gs1vqf39i
DhD7eN9p8NfUXseSiTFliTJhGhsWR63/E4HqqrvOn9qBBmLQtk20u6lqw8tzqsyAe60SZlyc7lhU
s0qKkCxiLNeXHo10r5BH51k5GgpM3SBKYYzB3o8l0orcwNVTqiiFHdqzQqi++TeeKERx2piytF5m
uH60YwP3c3GqvAIUHkjgwgJC4qZWuCrJHj963m0fgFZfIap3icKRIygx2KF9qcmO5vuh+RuZdMso
k/fjfUfD7PpRVtt3TOBK5D/BqLb93/I2GmKTqoZ8DkSfrIc8hoTCQAWxXzSrpxcg6PbbURUw9/3I
UHd3aASJl0rl7C/5Gxj0RliQcJbB07bq8ErSTrWesdrP0P12nSJOo/voK1/ex5g/zmideKMMdfwZ
8ne0syxKouOpWYIyhFPk/pZu9SHbBD1FOG/WXvGNmlwT2FOBE6jP+YC+ZKWjzjeP7Sv4ruuV5Uo2
qG80jR8FRCZikmVDJPvUqAVdF5rdAxt55rdPYrQIDIkqN65kKiOK/LWL08PjfRiV+BOdRMNq2rRN
ZxUw+6KT/fQp0ZrOE0f9fM2VErem2b1/nmgcNGMv/Y8qrRAlPc4j7JNKpS8pAYT8vXdnHYlgCybA
k+up/Db2vgNuaeengh4qSncjBuxEsM2hmxkugUqMTL79Dpy4NDXsRHUOJuT6cfDngqd1B+LBl1oI
xv1sezcGajdAK7xLgS9HyNjphT1YnwcP//Z7oI1g51q+k3eDC7YzFvuz8IQ9+x/D3jGvNsJyWeOY
C1jH9+NShszQ7tjUanj8AcstIonjo90jZeTy07as72zzre0EGfLSy89FheMQzO3Yz8Hld9kReTtN
cj1jWqGnWhK1Lcb1Wn+FSRDiiMhdzZ8OZwb9pcwzVlmR1hEXCRVkI42lQBmY+IjU7HrTEKrEyQjN
rORUK9/V9XJzOkowDGCUSvrnW5b+y+UIbItDK0GseItEYMLNOcd/8Fg8gVoyaMTkVOoZNaBEtGfJ
w8BJ5mBUNO7F+uFgN58js04mkjyABlSNggWVGwWf0uoJYKbn3Rx0Tew/O1UAie6//psV0VS04uyh
ruZQIdRbZXJoORNUcaNV7THL3akpNJGWayFFDS8dKzu2AurffusevrB2vW4dRbTHSUpWPUcwUQ2U
EODeTyB0tRaoieno86fpvC1AIrOJR6YVIxUGzDgHNQmt+QCyMMMiVyK7/rSn/GoF9DfmqbGW23Yx
IRk1xhFq305HwLwn4A8PXY6AWR81U5N3uDBrZRqDFK4m6bXu3V7P5GJ+uk3qxIC6nmcr6CbVqq0a
7p2fULhPuIlVONzePYLb0FKDd2jOBfchHE9hJLsOp7GuNPkb4Fg8081oMzcbYx81+r/EgVSgPWqh
UnU5a0Wsw1o9twauZFR3PTZ3Kf0l+Az8Ok2PISsheO9pby63OPM3axukpoUsb02N8I1cW+SuIbiS
l95rCfLhX/gu4f9vx94aytlYYaYZKxSm10j7oxI3ChHBQ7KUxmGBwpt+0nLkftLG8+SHl0yMHmKh
NBPu4yL9lYcl9D7eB8bxz+Q8odXlCHFE3rKeJ4ZLp4VEyW5GD7GkkBEpYMLcetDGC835RosWKLiX
i3k//CYNF4nH4xSxiJp8Gg+jM3MMvyvs3NtbNrF7hJeFApTLNdgUr1L+8whgQdKao18rHmMHhjxT
vzMxF13oSgqVPNyhx1l6AR1ft8s4VtGoHrfYfWF2EhcQDXX1JVe35pb9CQsnhKy8imJGNJ2v2CQj
6dy0BSuo79m95/6jF8v3bjKsYA+CUd86ePRmoSO7WanKURwxoRuyM8/6Ike18wMrHLltNQM0BD1D
19/rYC2WXonnMwI87htQCRmtkSn8xIDAeZwl11Rop5nbGwHCNCjq8QgTSS/UlErzjhumHSE55YHj
3jIsBy9NDzg5UJl1KOroEMK45EtTkkWoWtX6wZ6EBbR4UJmMzBeDJTONY3BipQ6R99Hgb/fr6nB8
qVxRXZmeIgtIMPKIrB+I21KZuPNU9o1lnlASKY1Ou4TdGAI+K+yFu8MImBGxtS3saX9pmDj62tEx
2Dz5tY0ddCwFX3Exg6vSp2+TlvLfoNqzEKs61JVsPWmqJBmMHIPdCw9kpjK9+CBYrEkxs8hX500G
4yoF7KfNi1YpohTSLwcyMHu0nDCERy4+4P0h+0qcPve+WkhYMOpdjVyqzom/MiDaDqdrm1W1V58Y
Q7fbyWompZV5QjjDBUJEUfErhxKabX8J3VV8iMp+0VSxWPBmco7KG85rw2Lu+kY74NutbrP3L09I
WkwtBvWd69a5nKCN3uPYjVPOeUTetZM8IPbs9+mSD07OJcll3/ZLL0UyWQGbSRqMVxkgnSo5B5Sn
Y1ti9JqE2fsq8skEw7yH8a8JZfRB32Yv8unU3U8sGJuPj4oHSU8WNILFIIA2YrchqLn7UrUhofJ5
v/Ke3ck4F0L5bhdFTQpO7JOsZKvdpp6KvhzjCJ6kthVNi6XEJujDggxRrThDN3LHPnJVoRXFZXPW
xSEQ7cbHUgRy7HuZV4VygKMFiFceA3MgA/2Jcijt+ZuplJGopvzoojJKV2p3hgiVrQ7f+ryFnqt5
JY0NDIL3TyzS2scH6CCRsaH/Ad/MgIpoqa96BFZYaS1x7AEqNifU7Br4FVhHGsXPX4gZsppDYq7R
YDkr6syhtM+ecITzBpbh+EDZmsByqhwiMN8X47OsZ2gjr2jah4Ue3fzdVhbIrLr5J+c2eZgCTWlW
EwZy/FWTSYO3oFuuLsY6OJk+MLHu/zduB57CtMyN4L8lij7lYbLpZx6dmyMPxOveOG0imoZa1czo
LUxEYX86txJekVZCHE7RMCzgMfk42BzyQtb2gHz92u+a81lc5B/JLAEXs7eFQXBIdZTWu6ShFV6L
5lS/BLXA2A9sAPQ7uy/4Iimz8P4sGk4d6UWRHUcsBfA5lJgA/2o4u/lFQm2G2SjzTneEmdqlULGG
jO58JEmR1+tNk/Ok1+kOh83h/NbbidpfHluxQxq2k+0Lxqir8elqRbSAhANtwrBWEuSr9tF5zOEz
oGUZxDtVQVNuCCWGGxLhdxmU4u3arcump96GqttH5oE32KFCQLdKOtEWi1BpSCUOWqtBYdUSvLXM
advKiRzriCCul8DQqPPLwJBcW32Z5dwCj8d6oiMJBy1nDtrMSrOUB7VKQzifcOlMIVDTvvi3j+ke
pRcYhfU7qd8WgL+NwHAzh7gPbHFpHDWhsAQWPhltggO/Aih9UG+duC/73VXqME2LMjznR1nM9Oyh
u9XF0Qn8e6XYFVd2/WW9w7OrILRS6suHN5cjxbkifLnahyd3jZjeet2r2jT3k/3eCreVaLIJTT6W
As7BEkBFMh57/pvkOTPpoW5fy84vDJN0dG9VlmZw2cQ0EQiO5PmUjf5YkdekqZXnJdeFOWCsXB1O
T0BNUaux9dNsr5NpGXkVXWWK/zLgYWomzf4b9131THpYOd4piM7xlzvNxkT1TqkZVX6drIs/KZrd
4JIHeAjlmQk3I3wwVa+nAqdP3R3oddL+7WGsAzZyfsiUPOaL7Ge16nKtXCaZrLk1l08YEDv2McZ4
IrBK3ZxKHOjO9eenUFse8WQe4CbLBh4+iuEpT9//b9m/Bkohcc7i3IIjzIoF8tR7fkHs0RzHpgv3
0CefU2l+0YVlEfuj1AwkatKTSHRWIkC6oG5Q51inKFlf4LdgknFOjUGxlpEBBOSgtQ4CAmm66Td3
tv7TWj1eGuHGOgUiUOVd1fAKdoaG2rhP33/YwKppgZGgf/UEwTM4mrknBaD3yEjvvq7vWHu+/xnG
1pmGvtOT2upgGhJeVlTnwM7TpT7/9SY17p5IngTas5tAAJDiSc2U3jHuOQ1zkN7mU8NwEUTJWXIB
ZbgDY7zRDCQC/uu0p8Dkldpds6J9BLSdVOsj1OBCuZJ+wOeIF7D9aAAC40gK9FF35d0MYmrZBMvc
qhMZQQg/U88wqyhlswYUm6/elZ5Fe+TKIFJOKWiGOwwRs/+Erpcz5BT+C8nVffs0XuQ6Ks7DIjQ/
JKyJdCh2mYLb9pJHBJBWCVOhhn+OrL5khOH/Gfs92pQJywtngB5vlVq9go7RcG/o4rUlYa3RUb9S
J2VPh4VcplAe8Rt2wH9E4urGOjjvTZ3RYIiB0CMfs6D6m0GID4dR43TPD9WaKtnvZo+qGrwiLunt
lN2HgkGT/mlEppX+NvCl/LRWhRURX6ZVjrGwzzqlVqcALOCLwDd/nbyOyvWsV1tHFIfEohzGY5dB
/5h/An8TyradZHka3U0BDQNvV43KE/tyInm5ufAAulUEXa7tQl3uN5cUUbXIWMhkZtYiDH6EyyCC
RnVFuHxazSbldf3x8aFzX0UFWiKEa5pyXEfi9CRZ8bTMMt8/pGcosjXx13SXORDHZyj9kqYhqwab
Hp7QTeybtKItbBPjZmM7GiKyaOd5l8cqYU5MM553Li0YjHxwkNsyPm98OofIc/xzcvMfDx4MMPZ3
9s7zeIUwxpf3untO8/4Ezuw19fcuVhVDJW1neTXGH6rP8HABHDYJTvJ5GC0epwiThI0XsGa2XnIX
RZJQxphgvyOGRa5rB33Srs2tGy2mKASH1G6R4tst51L7VIuVPL4m12RFY4pwZqGiMuV5AfflUMtU
UcG04apAuIkyFvOVAxBG2mEJ+Li9qbPceCs5N68RSnBmnpVt8J/bEeoZ/VP+Y6npbXP4yIJRSPgU
/byxjH+n2NmOlRMB7EVlLnROR5u3vmCL+7k7qvlqBz3nqs+Qx3b/QHKx6UhPqVjUzukrcikKIYG6
QFp2gpGNi0JBFRKUuyUmMcA/UWwB4CPlfX5hjCxfA9ybFJib4RDzXpaxrssyT4VlO+ffYSunbKM8
SsM7/VERZHvpQuf2+KIhck5MqeTZrq1or3sjlrNbq1A7F09ewbDeMkq2RIAXZoXHdJyHcmJ+1+3W
eSMx7VAy/P/fsHMiEi/I+fShNwQnQldgKnV2gXrPuuoLafpXJfVgOtMSwYXy1bNcuvxRvFPrXhA3
3sAa5kLvsareiVfnU9vhvLTV4XEG4T4cPhejvtX3LM1Yec+N/a8OpxujnKnPglSYmLsUvAWS2Nbb
DsChJR3F3lCNa1Su/RpZL9CXxnQvs9zncuYqHalh1rwuUnUruQkPbtWDkczYHf8aqNsOn4lM1ocn
UpcynsastNdUb2ie72R86KbY+VIullTMCkcS7ateeuh7LKjtZHHVVP196gyEz+XXRBgqEjb5tmzW
6w8T1ngUtO8hpLdBcZ2LZ7a6RNeiFydnZYmnVVoaEpH73sBK285b0bwts3mNyz75CxpeeZN1dLGZ
oFKjeCIhwcDNB3OKnWnN9rSCvYo2bO9NZ0Y+6Y+69qV2j33FzyqaKQ6lNqX2ZzXM42diLH6Nmzol
E/AjaRNjHDis8kI09+S7b56dv1erN3hKxKH4mQtMyPjkxgXA1veBWWBc6Gldciz8gCr6xVKQMd0i
8udbyO6aCMEw/IIzvRREmxS32I5T5gTgTqYqnRVfd+A//6tQ+dIgPh5K7i37cBPloafTO6mhZ2RK
v/6jflGIfzt2Gmq6Pm85EKKqiqIX8CH2T1kmbIK0SJKDBKIJ/j+aAyGiLCOeDktGgCk3Zfwn0el+
oZrF4KAEFrmzWHQINgUR/fCNIaPWwrO9dEIyWv5rzNqTsB0Khf+uJq6VmxGhEPpWn3N0OQaAveWI
OwnlzmYZZM7MolYmp9A8ULVtDC1D7pCJorrx62/BXnqLnS/z92Bxv4D6r5nEwMthdZ/zWKq7lYgt
ae8JIy05ole9tlSRFL+J4/eC3ZDUPpOfi87SWX8XJNpWZaUSf0cYyCDSPF5xrbTG0/WtfUrWJsth
xz9pjfz8d3ma4+sfQzEW8zmIqRz9qAt0bVQLcmJV4vZ1UwlyBTVGuO40tKOS75R7n04PeC8PLh+e
gPybsoI+pq9b3f6qN1l3TyGAMbp9UoNR5uc1GfIjJPwjIt5p2UVS57Nn8ESz7aE/fqFveLofzUtX
iDLzJDTF7NJHfWryge2sr79ELNuzgag6WBUTTPtkIfyRgxU2Gzy5MZH4NHVm4VDXdh0r8pBH9qEM
ToDwu4Ss6of6nGbM2t13frDOkSDH2N5e1yOsa+xK0zHE7Yl04cNlArOc6OqqBYl3ZEKjXy55ISb4
1qq8yatlU2esKqVq6hMVYLXduYHjoXzrfo9a+93IosLeuZNUDS7V0O4GUxgjpnrxCyQaODc4bKZa
RR8KLwiLHJNdINWe9hsahWo+2+ZqnJ5QZ/2BA7097t2y76acuiFC1EKtLnS9ufavTFf/9sQd8dl6
+4Y00eXfN65zmtxzg7jAWeqVumPORgcmjcJAczl0Bef6HrunKF/u68NaWp1JuBJnAokR+LrcvUwx
RegCTna8zJU4bfsNo/9/IKWsM2pzDRr/exuBBFUCFG7FBL9Rd875hRL37Jif696WOe3gR9lKCT+k
IA6eiXIjlVEf57CdLZcOFl3t0G6x5biG7XdM0pxNGeaI1bKFVlklOizES8v80O+5W2ziHbC5Itpi
qPNj7qMpSRUOX91kY+6DKOOO5YX1hHCvwS+UkUvuQLutMxPPV5Ca5Z3iKZ6skaAlfV2rPptRQZzt
LknyuhPRrpTFkflSd5JMkj0x1gR+kCbuzf26voDzmH23NEbUl7EKCNJ8ZefCQ5qk/zH91rFAtMum
R8LR7i2yVnFSWGOLVIDDs03C2Hc33VevDqMz8U+oZ6s0COlpdGEgXMV0f7uNTTdozm+uiacxh9fW
lk3bE9okNd8WtWqjAQ3pno6fXzker8TWCKUm3P0t1/uInpWOieBtgKpWnydnGfOdZz6/jalLPOG3
Bt8dlioX8uAlZaXMJpUpzHqvdQVL94oF4U+a4JJ5IUlu4+cL5navRoqcqyMo/YCn6tpCwR69g2UH
7HWCd5aJ6hSs5i9AAnpkXug+tS9rl3k6LDXXTmTjj9DYEJbWWRgaQeXwGJm4anfJpqWWx4nJbw6Z
p39OdXd++42jqA8ZRQJK2HYoj2U1QJLFruGH9OAGnArvVXskxKoG3HJijn5UjO2oqcp6EYIdHWmk
0HB6Maqd47fJa9/u2MlNGiWD9AFC3BzvTLV8qzHMVaKh44F/u3YudxFZOC93W+M+M7UF5LpBdSBa
uwRzdM0e67yodOrUAyU4j+qLi1sqsTPNP6Gkgd38FG9nC53QINxyZ+KAG1btHlejrB1+t2lTuJ0L
Jez+emhP5sqlPcVRMZjqN/440BqHkmsdLsrvfuUEZ0VKpM+r7mARFppgeXG6hFja+G4ZYJvmPKLv
lCDFQoavoSCb+s8KlUvex4Jy7K6/tkiS0y8I7/eMrnjwX87MlBuGe1bnoKiHJ4eL3GmtOQsMtoof
jojviqddv1jG8wUMVV0z8Dsxc+vtjCNRRfaYL1dEVfJ9XisVmqhg+t5neZdOvZcltdMShKKyksJ9
4h7ZnKL7M0PEtk+06Ew1KmiI1b58w5adZqX9iRLZ8/zzWpwKJ0TfDG09BPQSahoKGce1YQY4XnQj
tbRTt95/XY1MQDoo4Lb3s79YVLBgHkvsm9vx4+3YzDDEKc7bdM/dxw/3g41bldXR2vy47Q26hUnc
VzTSBYdv/8BrZVxBV8bkcpNHeJujr+csATq7rQnTgKqh74el7aVH7sOUk0xxlcLcManO7bVB/hm3
bSnNXcQYfwJFac09H7lVLxuUIEOkBciQIvaI367InGCRW8Z4erkM01YrIzX43LmcjzmSXFnAKhoQ
h347DWLFelcWOkBJxuLguyLHL41Qyq7uHBZMpBhFvAcCuSQpVyGuzL3QAiN/8Pxs1Tnks9d0olOM
leKCzWr8hkKEyuDCFhapzh+S+ySKC2cjAycIH8EOgnewFjXfaGK9FTXZH1/BGaeSuocbvPiYOSI+
+/xgpoB42FPXh0GL53ePcTibnY4TAXmNRIAOPzmPdagPgIkK6Rcl6LhI0YGvncHIwTNA9IlIH9Z0
doQrtNBmQ1FbTKMGDwJcJ45jmFXJOt999xc/4gxXEFhYW5iMFA7bgIiJ+oj1hpBiG+Hqswsz2bWq
DTtkv+obl0ZxhD/HJcQ4x+QWlQOtQkYiZA/OqZ31sQYWyzSydazFJMkX5Yn38uE6agLDFdHSadQo
UCjVMHY9Z6GMOGGWj2YjYT4JK/7lttpi8+lVnyQCPS6INfDAyKVeNiJp+ktvFHH7/0yOTuZvIiKo
kaC8R979yeeByixB5RSWNb/0qQAVu4tww/MK3HOxhlc95/Fg7ckdeEcEvg8t+dyTudBj0m25APeF
N65UAIkv0DRbzLQc7wRXEtKvUsWjTTchRLUpdjW8HXt9cMw6pp0/lmAFD6aD5sIgvKC2cfy/36d7
CR3x4Tf1u5RGhdRazb7z6hb0NoTY1fFbq7b+D+kjuWfognu2jIRlTnTvdlV0RwL1GdvPu0YFgE9N
Kq4rkawnVUON89wtd0GkLs+nY0oS+ZXelH0uQANwr4Ogkw7maJ87OtpkLgaPcaioax7esD2Bt4sX
0PbBgyT0JVL9IUgbSwXiFfMjBjhQxbHrEytsGavCl1oUcx3Qb+BOqQTqXdX9ZOv+EuU6L3eUugvc
PrsBeSF6qkhjhYBtbAodFTL9VuwUTNWS0dJ0XdNxGcd8VkT75ETPuO7A4cXoySs4UlCd786H2Iso
YaN7cl8hbGYu1ew0huyWvAN4+HfdyGdEJnhPfbHf9NyPN0+3i+Bx/ymYxyJ7SQfbYE3T0seneuB4
2PRxWNDJyLIqaxf51NkEuvVvgofJ5GBvf1SeMCKBExPCTibhkdovLyAC+R7O8Wcs9pjaz8u9BKYJ
9+RZa7aMnbA1YUpHHKvCh3WxDSE5/CAZlUtybONQ1ALSeFWbC7wQ6Vu9n4ESvJ4+QSPzU23UirzB
MEBqMC4VBYPJXKLYzIPYd7VxyfTwwNeYt6TiXUMHg+fk4PkdYlQrN2qJlARi6OpaOFmsunUMIiOY
2iAB5hmCKK8Jde53IcIf2M/2gjooopLG6AGfpMiQbodwhkRqglinc7VlGTcdZnezDSHHA406Z9G+
4i4R6DvBhCpHTWIB+BnPL03SiS8fOkcjFwqGYMGdzOCOoaAU+0cwkIpk21H1Np6yfOFVZXNjTtnV
33ImYKBD3XNBkHy5Q7uASvd2pfg0iosTeVF7i0MZnIQJTg3dN1pXEVfvMLCvHc9qZbFu1MdeFv6x
d9XCZrvCL2chfvTO0SiIvNs2RlBnOWZnpXz8OA/IuVRf71rr/nHc8nq1bPGOXwofk3ruLXoHf1xk
E+64rrnZ1EO2GuHNABj1SVrEPZ2lGsmqEemjdxGh3zbm63nsmHo8Cx7C+BYE+iX9T/+ivVFNE08K
98sYb0ErXW4jUfX+jRVc8jw/iY6tbyYh5+5YSLS9LzcHvZ7ew4Eqfp0U0Eney4VHuhwQPJVovrkz
XVv6+kqcXUjAD80rEyEvEdUvkvpmJlaiRGYgRk4unhnei8wTt2c8arq29WgcbjmEM0PzkittY3VW
Ydf5GHBZkjWqyNKT5d8XkEWhwHjs4T1BfqJmVGHwCDrtqthYm7kyRjd9pWSuVD2UdZmHuNZ54TvZ
zIUrh5opBrlk3LzW6e/7G2PW/6KUQ1BVGymIVT/5IkFzkXkzT0oTScRjcCkcgIjyG1uiQDcWZbol
VMm+qPQv5LYRRcTjg4xI+LrOF+6GveJOO2LwHHIojviIaoEGRjf48TwuC7DQWYGsGWoJD6paUbgB
aKnF4VafA+A/fuydktksUca3G6Y9rmIxkEDlXFOU/fN7ImRgHA8bwmqIACwhvJgV5dvjk3d09veZ
J02V10nQ/H+xvgo6ABmkSEeN/btP9fxosFWe123BPwsQaA4nh9+X+ABj/5H1+l+NO8AOrdM46bTu
rtNEPXglaLnWBWLmAymri2ftjLZJvAlzB6+3/xV3cBfxLdgVKMkOe/oiOhTJxa3c6enFN5HW1gU9
g83sqRgrfeA3q0x+5XoYn6XyzAHt2tcLfX3f2s/BPZfIAAm06SE0qHu0IOU0aznNZZUmHWvC1J6d
GRA9vGS7lZF7jxk1rKBT4q1tL04ozUfqef2OdFofi59gv6hhb2+oC6XKatekpBG6WDcLpr4daCL7
H/ui9xBoJnbZ4ACE0/U7DyNjprxNzdJAa9Vew76pNyTMgDXRn3FHjZGL7R7paITEeoF8cTISCqs5
C+h0GjHO+AVS8M1ySRTb1eWc+hM8kmBilEZIV8CGBP9ow6r+NaYnI8j5s7xDByx1xRhbkycA3/RT
XR1MA8N+D2YmLZ4hkg5LmB4HIyTXyG1GP3jynM+F10RPhWXv6AXGDtmaarOns+nMX0nysWTKHz9G
25sFAZa5XqJkCqVvYt2X9xJ5MxTGgS/KqWS60M1twE7Le6EwRkdzAGkrOltm5gJBtlTLbJ9ykenz
I2h93iVnZFb9aSapSOgfYW8Osk0vzW29GN3Y0+kjdfzm3QjLijsfyBI5fiO4A8DBj0BhAgssjMDh
GhhRo4BmE/xb9HxcVgaXxK9GoG7iAIlC5VFgy0kOWUT6LFuSw/YwqfOhuywOuemoysxHnFOLaccR
To9qUs/LL5txMtR1i4G0gilpbVERnrHqmkIBnhQhI8O07pkxtE20goBxJsHB30d5Bx0OFASafH15
bKX2QZrAo2WVt7X3BBcFbrxvRBlH4TOQfU4a42ANLvHlEBEjDha8m2s32f9AAWTgN8GmYf3Vf60/
gYt0lyKErjNGJeBIht5HZXLaKgW1b8YpMe+bYI75e7Ydkrwntuu08bJpSKYCi/569B7C9PgvUw7O
77jPam03KKUQdvZ8cnCWNHgEZf8Qccp0x6CWNDxF/4y+a6gLGCAQYF/aDK2fJtcmc19HIhV6UBrm
SFyC1hsVWRfMQ8jIZVY6Y5w9A5WiPDeb2FD1crZZXwVKUUyW9yK+6Vhl2iKH0av+nGrHu390dZA1
dufUKdpESgLzTt+15bziNVOxGAdIt6iPpQlSTuUt4tfJVmC2TV01tUozoy/OVMJb7KsF3yKzSIc/
el61fI20y8dPzFJU+ynByWgakSraAQyGIFci9rON6DoTctxvo/NkrrJGoTi+BGg5MsjzQOsz12Nb
ugzQpGCPyEjW/H4sBxmjCiSsv28SnohN+eQoK0AKRN5q7SxK/MmqkaZCGUF7kZFRd26bumOag6p7
w4MJSNd4mSjKv2x71Qh3GqE3ijMHhGAaL1gD9O9CAP4kHbrfW+z1Ooz/dTsG8DEzrOSnFLhVVkKg
v8HQWZ+jb3kXgrnXj7bqp9o1tdHtAnindWH3RxqsUJGFTkxdPtpOaFpq87IBAgLSIRZxbinhlSUL
DrB4lJg1WR1XKxIQl/sNkb00Qn7A193tAr+uHjbl8g//jNV3At+JB16J0phozVIx/nLhiPvYfYge
0hqgNTs405ow3d1ejUpAOMbh9Yr/M91O+oH6ilVHAIwX4uFn/WHF+k0lLQDuQ0sfxIJFgjzrVecK
oqgI4VdrB9HTlYUvODDs4oeDtT0XegWavJnKl/oL0j/EHla/zMdxZzD9W6Lguk/3PDH3BOBhWtVo
JauGpx7Ovr4ATT3KRa/UkbpsUhexonr+yTkMogQKJHqGHTXNeT/cXLoTMP0SmI8z9cO9ekGHc3h0
RKuLgf4q8w5H5wI5v97rkyBWhKmo50Fhwdx72Ob0dGywLVtdZc78ZzPDdbOjIyN3V86a77zTdpXT
BSdU3gvzCCLGX2+PtDZcpQWB0DKVM1fwbk4hvsuPzqHzXRMAHwVWcTvltPrbMOYXdE+6kNaW1QQd
OL6X8QSXgj5YfB8UxGqxkSZbsdHKf9l9lEVOiZ40sr6uom1n+GeVDsXfCYomjQaLKJxQn3TbqL++
XUo2yhF+HO8Ot3I7uPcBVFImujyhLMjXlrVTDxckVTwaKD/yiX/0M+U7gl76zQ1/vwuZbiljEe2P
RbjjZ+vATs3DKuPUF/C/JH8XxMLftfAnpIDYvQSsfkuEZAf4gMlc+fNXkwxP5TTlaDjdbYdpBS3i
F2S3QL4ZObg0WacW9tQaO1mYVrcXcpE70LUd1NvTAR+nfPxzK4LkwYH3/dYeHnVOTE6ZRELyqdKz
0uMFSWwWuQmardlvGFShlXs3O8idHg5URw9CNdxg/ScFW5Ic91cGXlb44reZGvZ8pkAx512XuULb
qV0W6T9pped1x5txFVVInr/MFXZp0ROwO+L+G8VbISxLsid4poLOk4sHxuexP6NTCxTdU+beAuWP
onT0sc0uvC1sWA3QOZ2XuS4v/0opxK+MXnCGp3s4YcvZXW2Veqm3iTrh1o+mGR+UJ9dKBBxM7ejy
qPilQuBJdriddN0qkLaN7In6CNObN0fe+7uO2EoATPTICpNi57hObKXEYscsTzJkuQ61dRfA3K+V
JJOQXyQXW1LuSAE7cALnAY/kpv39APFPIzQqUhxTSSnDhVGKyfI+3/+4r0w16QIvFztFtqpNog0T
quDeSXown/UNz9VBtJCVzNp4ywZKxJpgLrymSQ1DkVlah9481x+fcqqtW+c2V93dN+5CavUFK+tQ
BSqjz1yOKMzFcAwTDVQ3WixOsC4bDG88t8UMQvTLkRNxj772tpMVeeV5clu0QbklVUFWZ5AAQu/n
R1CwTmH7+2hrHfwE3JZ2lTMiWAYexte2neJa7MrV033OaqwxdSMpjYXihltuQPrLOZvWWbWaPaTd
Cf29+a0grVWBREVw1FEQ5II3vQHRc6cqaLX+/4LoNa5kw3iCrJWFTjnmbA6ln/mpGxIFz+ziCFzO
rTfIhLya61ZWmiLW8+gozg9gzVDOhJKOjdEr8fMVfYLcxuNJxKc9sUbt4ZJfIzRxO68BbHBQdtWy
eqf77eioybLivqVWtRpN5M+arMz+YvzfFfor+3ZHXSqB0Lo7AI75eDwksmNr3QybnmTSeOmYa+21
ls1f2kt0J66OmeTP6SDsWSdFPGCSRY9PjniQ6MsDqSJJQmplZmRmFQ4ntd7B/wMh+/RwU7qA6DUF
twx0h+iqDAj/PZiprNr+EKDsXMe+DbtZUI+76sHrFaA/jMUNBA3LB1C4BBkVOqpOEYUuhhpfmfvB
2eDIeb5E3qoL4+xHmuAthmEzd/wITQKkSioWcYElcBC/cXTFm63bijrQakc80JOJtxn9lTyS0Kq8
Q74HbPkfJboW00T7Vg8ywefmtBmrwNijN20hCwKvR2UyFE3XAyUbHRJ1ZCPc+sTZKCcKpxat13vA
EotR9Apa8FaPwMNGSX4QtzGGob90bUCs2u10G1obMo7mKwUM38D0XJHz8/MUFLg1JLYizwfx7uu0
7IRKMbRfSuR7xbI6ADQWFEkIdyrYTKCFPUOdr8IxjuiwA7wMptmcBeBODKTZx72IgUvzwdbutKJN
ZqkNZLKwEbxBacgiDlCDqKJSetssyCSXBaqyElH7RuCsqQBvpyEnf9gnAgATZPkFlwVr4lOInoFw
U52CJ2b7tpFisKCQaXZkhz0sX09pwBPOAUfXB2q1PSrsd4W3fiRn2Ve/d+fAUv7D9eKaxjtXjuEQ
gkQYs1HAzkJlv7Fzbf7W/RoxjkwNv14EdtUzjJvTPTBwVgRqcA2CJekUYvF9/AfJXa9AdfXHcsI1
ozlFzlpMdjaOkmcFIsXiPjTRYDZ5IcgZ1lbao/dVJGDii5ALabiuea+tOsRpXXtOUIKz71KyDsxj
LKsf0P1pgrlbfhIud+lp1IFVntXiLo+QyEh7LPQRhJFLimHuJcRxyKOiJoatZel/V3iS1zRQuJeT
d3+Q48fgJQRE8yb+1y4zbuDjW7kCHBXIVVRMZgPbEju3q35X/xfm7V0r4arb8IDu+bkWwylG8OKH
ejbvQigLdlFAlweSdjujyOmA3UlnIxauq2gh5I3lNlQSNrkafjk6uTuVqggEKSigb5+UIL3TrnKg
0wbK/GbOQ4FTEoFt4bfHBQHld5ATLqG0zZiA4Q0nejzfItS1f+IDyw8/H9liKxCnAM6KufjApxu8
oFKFwo9iS0oMAs4JqQ4Jhox8R2cuEx572XtL/t8EzLTrqc89yjN7T/JBCeKlgUTrEpL485SjBM2o
QTuUVR0b0TxPPYiF3hozPw0M5pnN+5D2zV3QidKrQkQvhivEjfB613fK9mgMmEyboUryOnVH2mlx
xPtP9BKjbzugQC0z23d72B6baOxIcUQENoWFCcWbuXM9nvBY9oSblkd/nZABfsuQ6lalJ2GSVCHc
xtm2gWklbECd4h7MDL8eMtJueNFTa2FUKuZcrQGattEnm4zcWegZZfNgMIPWqysIu9PH91vNJtyu
doZuDD8nqDKi6zg8M5N/GYhElJklWXqlvDhyjAGg7EafE/SRPWmgfNQ2nsyL9nOc6+17yETd/2Aa
6LSwXm2uEh7GnBj1qzmgc8CGoTyy9ihatgSfwi1hiftuEtAfgAKENUdR7GiVuOmWmvj0MsrnRZf7
NAw7CK9R/rSq6TrGqWGXjxVBkTaN3TWG2rPM/rTXpDSfCBKgpolE+uKnfnlcCMllcNn2BrpdTtDM
t9QmVFgQhD20DugZLW3xjX3zw09xZPerZaFsdwP+genwRqQx6JBYHlA47UnuoeJv8nU0ATYhT4Pr
kf5BOw6EWji0uSIF86jruyKLO5rqyupiFJ0sA935zRbiwzdHnuJWvOtk0Ni9mygM8D/2P9YODc0K
1Vpqv0ikZYdhOqSVzZ7WOgXT44iSSrScJdqlAu/0TGdU9ZMtl37osG9mOJzO5tFeSJTMDiJ5FBgS
ZxoyUJYlN8l/1vHrx/FcuOvdDevTl1yrWq5X89Pv3ox4GF50w1mA7rGpnWCkh63QaJblaGVA5k0j
O3yQ/8qa7xtJqqA7+lH1c80n4OqwlCZPhh8PuWN1wykxnNNFV3Q68y68xfdiVcAFE7mpE2bRjLpa
K6pFNasGjhq15MHUY5PiXl7B3CroxowdjZ6owN1P27Mk024oxPXLH6EA6E4asUAIUXRETSlgDsZq
yU39FHzq8t42Dn0HMUr2eWmV7+w+nxgXxuWDQbL+30rE7GVkz4vGgUCBRDOd8JcDcq9R8xT2YOSj
PWznsMKTa69/2NdVQnHorIX1dM768LyYe5zI2RndSCk+CsJMkFr7VIDP0tCdwyLjew7F5xIpHp5F
gKHgprVhrAKxPe0n4e807F9wffj4bC0zkW9jPh7ZktZJHn2h4ujopnGtuabDcrc1c0BxXmlnWvz7
NsWBT/EGYZtuLm8pt1tQs9lEvFDnTE2Hrq0nv82SjN2jKLDLF4CrBRtQqgUKTr26va966HKhqE8L
gljjtZ19p5R+gjdcNtM5/yJbN6vu+DaHGlZBnveXTRp/tw2JYhJowFVrZpvnbVfBnVGpZNuBrFYX
xFYcgkj+LIn6/y0EmSeuiQltPWHCUhb+vrFK0FBDfBdjDpnUEdMl+tvaFliw63OfYRuvqStIdxCG
Dc/+30C0ugUggHFQingYUdcbwWRLAS8IOLBGXutE5GhdfQ4VLHBS31TURqqH43HvXD0VstNMhE2r
mYXJHfdxggoMuCut2TEBbJ1S+0T7RQq+BLAfRuITG3Zmp46tP/0/fgBfHUJSZMQOMvayx2FecewN
A2MN85ttYsVSI1ghzxa7YWsY5qbXwY46a6MFlz6dieAQZwUWwiOw9QaQd4QTFWbxoyRZjJBFMuZt
lVPpVPggQYfpW5P+0F2ktLy3SC8AkDpjsjSE/z7gdinZ9UWind04GsvjSBlt5gafald15XcsSG5r
sHJiCzVF1eqALVfIfVgK3PaTTeAYnJL54hWNrye0sn8h5phSrEWiZmeTSWK91DmoM7i3hPQxqFj5
WZakSP2WkFGfcY54U1REZ7BCRJfdFw9Ioc25z+HjhBhxrzgjfDBCLK53VHOIB0juiCD8m3xxFhHa
636K4AU8RVvqPNYMl9gpEwczC+LGkbjU6l4lykedJaR0VKih28mQIPL5w+lTt/42qRG9hVtiavWX
6Yi+7JpIw7HscN5OV6i7JIsQ5Z0hIcW/TXz+nzTCDehyfkpWAjxVhRbNOQZ7zTUjgWOb/IHfX3he
mpN32VeLrtDXRNOZ2hRZ5ZDvNN9u2oRlkpQig8R/SAJX8XQxL0M3gUn8+lYLyhp9lb1baEWez2O1
oUOjj7cp4o1W+atkgeVhSEuGSP3ZxdHag+HN8lnWBeuVRxEjc7zH96EIMco2NkYMFKf5aJpyawNn
9S2Gs8HDAWVCq5aRPjsJaiKhE8upRYF6TXS0cYgcXdHbL+N2IAuNT/lzd1hPVU9s0ohcVARuQOtc
ry0y7i5iIsNg3iZzPkGvRwR+4VYaW1pBaxyeP8FTZo3TSwYXrfbxJkMudQLgP1SWJJaVEUvbXFp+
JVf3xrpD14Ppmsl4thFoo/9N84+fPSAbdgSg9WdVn4An2Zt/S/vJx1/tepxyYgIs6OnP9lO92Dbu
L5tvea7LOOK71H1H5PlbnLAkEzoX5IZFUp8lKS2mBIMvaiJpj/n6IOTw7J37207GIzL2cn6ZpGeX
D0R+vCVjgK6f7YPjzpnR7Cn6aGFMjAPHsN2CY2QcwlirfssL9opOpDAHz6Wbh7EU46fE9hugR3b8
DEMTNaxKYYfU28mdTSsC9pCuYtI/VyE2NvNUfs1pmhxsDsdXo46JeQt4Z/Yd7LQ0baxgZIJCmbMX
L5eJyK4UsmRhaq1hhTd2BWif3VER36h4Xv49HkTeYjWcg47JtMtjmlLj//0SXC585TVJzE10sCni
HpkkWztkqdjISl3xvC2qhaRxcUb6EusaFIoggZRzPP/yh48gtqe3DZikhdwdrFkcR0B9xFjwCK9e
CNPbYJiUOCcHEFhoL72YRhCSzUmFSycyAuM3yMtcoROLoIbjpd/Ra8X8O8dhM+fAS1J/wwV9tOWI
bnVJAgM5oG/UI9o+jzRJTudp1rg1SEjl0MMJ9vEIOCyYjHyyzUaImHPXnkWdTc6DewmrvZWphdBE
h+7YvBdzdYE8fKBaxceooif/nOd8Zc5tE7sHhuL5UEqa7GK7DHf2ajf2mIyoHt4T61YMlbDIBfnt
12fA8jYxqa3npNcMj+tmGbf8ukpzKzUE7T8nWuS1i/CUN+M8I562BmgnzG53VMTbOjztDpQ+bjuI
aTOKoAwTowIJLo2fKI+jgEHJTrryLcuF352s5EEqBWeZERs9T5Q76cG/QphJEQjCVyNeCtO4uqP2
NYQO5mK8xPH2rB82OvTCvcx8CY19Aoq9kz5HNrFLLbSlmEugTnRmVaCYctM88ORQv0Jrs9+NKb0o
uUrP8Q7YrKWIn+LgkCC8H9LXs9vgybCDPHq5Vks2Y2edWmnzEA69XIB7ELAkmyQq2Kbpby/P0N+z
FB69XmxdyY/6PLDAY31eLFhGQTWlCKyRbD0s6+WjnF3iX6XE5phJg1WFGM7x/KJ1HtjTCs0Kjile
ghjln8ZBvroZ/iGGoODGx1Ic+b5Z1M8lLrJgwIfN58TcPD1yxXpYeI2JYsggz1n4THdNJ4Ea6zwM
FD0e0/AjyAEqybszTsIXyaPDGwmffUvaTjVhP7JcvHdUCSUeFfwPpk84SJkkE9l2eij1Y6hwL0NH
7L9X92grn7CqjlNJY2vNEVxmbp6ntmV2fhC5RdFWWSGh3U9NePyA+IOfCnjUH72M3IzFVHqWBET1
ygUr3a7D/AvSzYvRlA+VfTZwYg1WKZRLJyivZEVEKe0DnbPIA0D3YenEaM23kjZPeqvvLmv+wnSg
Ysk6zKyO3ACnTKIbsm79STZR1EjQr5F1yD3BhMbX7r10zx49THVHRHlMjirDPnSN9jT4rGWiGC4s
2VRDiaAxgNW60knwPD18RzE/nvN/9AvXmxB2LImcH6Gcdfh4NMr+1HxMzryYRshLjVEQ/K7iJypm
Y6nq62tNBtLzG9z4WrzSh4zynr5uaV3stKi7HeQoTi5M8wujAJjBEQ6fX5DP94w4Xs2bXhpq9Tle
JfMziMCHQtbre4yd3EF3S4eZUg1UPSV7kfn1t8UtybwzclnDpFwfM05EWLvn8R8xUoBkUoSaVRkA
FlyKmKUTkfdgqLmtgsFyEEdZLGXDZsZJPphscx0DcEVNBrq30h+lBI0g5MP4FjcqbFnUeh9T9l2s
SAe2sVL6LojCCbwVGEmEfkwZd0suOBvznuiNAi8muscGZQo3sS1XA/LCEdq2IZ5gPl9RB4BSHBqg
h5346dLOdZBFpgrsab1jnw0AZplwY+E5BLsnE0mxWiIXb70TmLYXYCHu+XgZb71cb/831GuWEu2j
l2W7/NgnZqW7zMjYv0tKSpwlpBsiyST7XgNbKbSIwDVrgXmAEEb8itQbyBpPHVnoN3sDU+qv0Aeo
bwOxvhp30fL5wFQCvYxVtc9bS0OeNpTiH0tKOwBn0IOf11MWGk/cCD5Zh/uG/K+nfs7uQeF0kFQ+
Y7do/M4HvgcAmYCXVLqHtag1qZXDd8q5VfiyShOCfWir1zGBtHJVZ1uUdrj/atKHwUUzBHQzTlcM
g/f+QP7u53kPLZQlxFJ1MSSx7P+K51gRf4cnvy007e8pdFvSjl8BAgfzJjo3F70QnBGoREU7KDpO
qpMMJIPAkb0ntjRE7LBLdNzfv1vTr4NXp04/+lD2pOaP/B+TY4mpj0YRWmSznMGkiVKm5zB2JQ2N
5UJaND86KYXHUPel9R1i23TvjwBEsdBVNPtEigxylNTDGXFQ+onRfRdDk7BgMlz97zcvqVXSvtYN
/9g8F7/mut+2cSQ8/HRSpoNDcBLxmV/zqLrdwIMA0FPdVIB00Uov8jhwvncP88XUhg4OLEwkf1ge
HPWX+nRGAm8RVq4XvcbvCU8Kr3Log/IRGmaFKmUAYwmHPQF9W0HDQ1wR8FskBXhil+TqivWmVrGK
/ZB3vtgOApgBM8nk0/eh45PD9rXAZMkqbugJ4x17BJOs0VkHPu8mrzZtuzC2qQyKz4AV17U49TfA
tHDux+rfVXsDVR47IKcOSXnb3dByLIKdCFWL+lroTpKZYjlXJbVZJ120bRAABgGPo721aZvOSLCr
yAFEspxEvxukaaJlYUPSp8PLSVwGkLTjbgblRb4kCzEecl5OPDz3UIb84e3Fzx4LruKwro4Lw7Bn
+GPcLj3xJixN6/gH1PQe+imJgY8CXLSRgTL+fQNsVQ7psXX9sFgUKhjmBPIz4vBSx/f0eaUew/vc
KHnS3c9WgCXB3MJyLSKtqlU0qoXuhgnUtpWD91VwKiPtxsJ/dCJbhCTyQDZoH85fBL67aWAtrCzH
/J2FDcYyEMAl/4o7II9kmokNcEFg6ZOq8lbJOcs0RtxzF0TDkekpmh5U3r7l1XUhJ7a68PtaBi5p
HzE2W82Hz4z7m/kIU8QF+bYz7mXJ3+z4KlTckUNpaCmUV1v2WjcO4bgScNWnRlDpksn0liApMzd5
YbaM2NtTRQ016rkU+7TmHHUcwYsasCJysnN9jm5EtkDedg1FbhUAZzLI/sBuL8N4C1hWDTC3bgFO
lCOI/YuZzaevE31FF/5GxE1TC2vEmWE6KJfbAAsRkC+3ilUMORXu44N+H70od4qBxL/pOwNHH2wh
8No2a8/J2CVa80VRoszTIgui3R7LAL03YPpBURocXFWGiIixKTytCKEuGzgG6zNgPXxW53IL6YD9
ql0qSY7RJS/rdym5K0F17EV7Jqs5BFkJfDgGCBpmcnkm+T/OsccNQwtKPq5V7Iobu0tZAT6uiASZ
s/LfTtkep2PYvVREXgisEM8Q9s3AWr86zrDmukxL2NyO73fzzO5Wd/fnuGkWoDRh/FeV3ePyrfaO
kwK2HkZIE2cG80z2ewQ8potevdt2kj+7I+irKDULZkH0ijXy9ggBNB/eBT8jxJrmpPrh2LcCbo67
nZkrRcFsDyHag+Wv5NLixOfacHvCu3JojNHNVTy44FmZvCEzFbTT3bihKGrjiJEddIWdXvJuTEH+
7Dy7zi04k18pxu4Wb1IRS0RIwiBrRVuoaOY627ROTXTCTDVw/O/hrFGXyyQYYKeSgTPcu2DQ/YRF
Jz/UAZzFVwCZUd4YfWElWfescl1MUznEzhRJOfQ7dRdE/urPoKnj5cteocMUVbBxdzxyjdhU7rQJ
np4vx4IGjogHbzxNMQTeuKw/fFKfG3T6ex5OQPTH0ktrZWGgzcNK+L524Cb2ob6xihE5vepRajJ+
ePNDoFG1+oxKlD2J2BeOphu7CcbBt2qQ8ZIG6GyhWRjNa/P1VBX7x5dLPH7PtyZ42OMp0e874nf+
RooSleuIyVucaf8CK3OcHSBk3bW4LbJbdl8zKEz2YoRoZSdA4lb5SivrWdfRBTlbp2IGraJVuNpl
gAaV7RT2eTGvR2YlqKlKL9EJTUX3051Pi2jUwoHALefPCwbG0Y+U2KlKuljjUa8zG8k1B/1oVCtn
fkYuFbGFd5XfWw/ArA5D+ChKb3FNbaO/+MgYVy7spumw8yZFKz44U7epblu9JAOSTklwUzrEh0J3
6I5jBicHa6+I5m3p6CSOdvyINEA2VFtqea8FWqfUE8WFdbllReOkS+II7iEW84QpuqQB1N25jskc
Otmrh1StxJ0/0ba9ienNBWTkZiKOjxZOw6Y8AdqwRrHdDR4lOKosFTtIbxmFNz1FMlq9vSXnEjgy
CJUXhJgIeKCAWZYBmRBfeu8eGLHj8Xp+eTvUenN2urPbOx5/EGRCgU0r8khBo1JxX4/9xhTXfXng
c7fXwZkQODlq4YGIULCsQJDkY2to9uNSmkzafihRKCrTDEjimXP9+L7FQCQFNEOnUEfmZvEB7dHz
8UNTlbfxnh2Wv5pFQjTdyXeCsrCpi9Rfc3ZyqgIUYWJqXHjJ/+F+JOysgwp00NICuVrHJHqb9Zma
nbV0wYLa2xCr0abwnnYDMwHrxKERayQzxry/xYgcHgEPykwsBWe1dTfqi9KayWHjsLFt+SeCKhIV
ism0UcnxtZN+ayJFKRRb2vlBBV9eoIYyn5uVenrc7SUoscy6WhUvzXNcwtyGJ3e7XaLrgmcJ5mkx
n9KwU6IrNztNgFe/Eb8ZlO4VF44u/27+r+evP9tULeXXu10VOOJFcIaodu5sI6gtjgxCnW9apEsK
SX6Lk0fmI3SErQuEAzbvTKb0L16sfygynmU2Yt5SCRg26tD5lQoEzVm0ZCjQk/1iPNwSzg6S7fkz
rO/xqsCdpF7IYEnGjoOOVdVIhLUw+85W+1Ikc0fprs5fTPHLAF7GOp3UHkPZZuJFv+7t+wAKana5
Pgc2TTTof70pmCq9FqjMMZo7AK80sKhuZrzfpB4rYD72gdLisvsrBmebv1ZwEApkuxKyFP5MDkBv
ypJ59O4+7gtLoAz4Jt6iqzi+9emwXEgmhIaCKCcSjsLZToU2791MN4KpvBPDzqfALSDX9v90J4jk
04Wo/FG8lS4Lp1pt3hIf3NUDz/Fp/NxhHCfAPanUgWJT+FBtf64zMY3sr193Y4ZaIkngQEHFEJfz
UakgIzLNjtLfRl/qvpbrqpIvBnlHYmp0XjwB73SDlPfEtsXaGutImqcQX4AtacRnSe7MqRmCqHBJ
Lq4rfN1BXansXMLCJnMBQYo1/iicNVoA8wTVGwcxG5FgJly2gxG8YukTK4HZbxInlznwc8Noit1e
7nrGa4aMEmhcZRCcq/L16jw37KaIMrKpyM7A53r9EXML84fM6YfBwunfmVwHByiKbzUwPLOZe53a
Tv9PwpS2HbvPRH4FfWaAjblD853jvYplkxOc/CWs6Vx70nto5ve8qXmEfFwSAGVvmiSOLQ3xpaR5
gSjNzMt9ovjjl8hQTxL1nDWjZ8Lk+jtxsCkSV41mKc/EEfjzjadfFaic1FqZxin8BcK86Pe4rs3A
GBrFAF18r5YeApPkj7ebZ0kENr58Jd7qu0ZsC2UiFA9FuE9qsiyr5hrj+kOqiyfDHmt6wmJPK0U5
RwYoGBW74ciiJXPE5SHT96NqNDT5+rJZ/kcjj6AyNg/0c2hMIIPSWPJWt3WkmCDBX8gpamIx3RcL
t1HE0dNHTQptfOPGAe+8z9DIaPrZ1at1sP2wkd9DbLIjr+5z9a5JVhqZELLCjpZBNCRhsIr5RnSv
uTPt6f55z8b+6XRBmsz+hZM/Lxbn76tNr3YtvmbzQQAdjs+8xi074tciF+htnrfLHvcnvhcGndbl
SakQ/Olva+FBx+NEaDG5mVoqPyfDmX5LXixWRodxV42+CMf5s2ECn9T8xiUH3n0J/ukbMqe7PcoJ
OjCnRWdxaVL/IUjBX5mStbjh4UhGF7E2QbOZ4cBqOnhwSpAeeAFr96Hr+ymYP8wDo6Hfxm6IJ79W
yF5IYJgpv4J78gIMyXSzcM1skMfSdUD4zhnLFDVAaYM18rdwPAQad4P3ryjV6FFdQ7Goy7+QqD+x
2U2hU8QY23T/HsgXwokwvrA0WD0461r9/Ias3NWEovgOHzNHoWMoRAV3TcRZoJ4FFGN7U4AZS6f+
2QlybYj4N0TpgD7CG2R5tH0lZ3LonGTPyPTY96ajxfr2Cq2zm5L3Z7BQm1Saq44EqkxnG8hUx/sd
F19nn4xz5NyXvn6XU8hGP/YuPUqtuTYAZ67HFv0aXqUB2wGHfI3SWgQplDaWylLTAY6swHwrVnnP
e9+Hbx4b72iUUAcNn0FyqJfNLBX7931dkS+vETVxemkiSv9Ln9OZ//0AZE6J/YCsORKXWBRfHqhJ
wR3bGHFsztlLd0RIWJwNlDoUGn2QKsS7OkHS4P5gwvlNZbbCgIBjnz1alGmGeRMcqhp+KZ/ZNa/8
E8P+bKiJbzcommkn1Z8RE4aXNsrAf+DeyviHRYwezEDtkLWzpr1S/GuvxIPUwtBMDe2bEMrEg7ip
4r0B1U4sKwsWMYnWD/Mx4Zu98UuGy3bs1MZr0glWz7sRRaKQtRzY+CDFd4Nb7C9MYPQfJ2gKfeiM
jKBoOdS7BbcZMWKV0KMR/r1lkeEjJ2mv7uaQ31D2ML04xEvhYdqEMgy20FIz1e6Z2yXw/H74mV2j
lq9dsqAZyNycssOMC3jmAqrVpjPcke+xeIPhfsPsH+pVQaT4jIra35WCIHD8OC7GtkdeSJP2buCx
sGUJeCu2U8WKEmllbk6kI9eGRr4h68z4K6BR4fQSqFcbhxtnTh8w+jJUmAJZL/J5vAT0wO8ZqohG
mm+wucppkJCORkXuWu9R5HXK2ZR+uOOcROHf47B7HVlumP3s3JiBLWbAI3htNfXkGDeR4lvyJSFP
kznRuI3nUZTSHOfe7lzlmBr1lmz9LoCMZDMRaO0iUO4EpskKdLdCZbClHcCJKHR1w1rmVryGyYxX
Mg9FZxSUNhfTXsZuR/TH/PbPgd9oHNbo1aanVVI2vtBRdW0Yfah1P01lsnT/3otrrY/fQLOTq8MF
ZKwla4yOU5kpq6k3+0AklGp9Y0BhHCb156VLb14SfWRg1RYXFWaiGAxOj6tvUtxdrg4a2hsnfc5H
mz7YMZwz4JKImZe91S8XkZqYM/ZB8TfdtX0CSXcOex5a3SJuHvnqXn78tUE4nVAjpjsPpVS/Fbvc
FO6T3YyKXywjcd1Suf3BawnRrANqMq4Wr93jMQUqbomq19CQ1Tvt4hJ2mzSvyzlT0KDh0k32/AC6
VXXi3ZOX0vx94CwyiAgga/QN4+b1YzN2y2c0eE60RxoFyi47TdprDwJ8rsCaHqAC5Slnzak3yxn3
rFJPfHNqM2SvD4lQWZX9lgfvW+9Dbm1T1Cu8s0qObj96cTUTu8a3TlvnnAw5Oo3BDLrqcTvj5l+I
JlnYDiGVz8IiYe3YyXFcn7OQkg1Lwkep3A1E56X2tX5siB9EOUJYSfrtHr5TSKNMT2FDoTFAOirK
VDbHChCWDV3HCcs+4gyMFvzjoPTg3EW9cOa6QkLrywlx97tABzGfH/Y4r8ipZ3m5v3COpAVNIFuC
m7oeQm8n9cI0qRd9I0zmuf8QBpfGh8wktCypGl70GX7UtwlggcBH6whKRwTq1tHqxURS7gDCKFUi
m8l0uDJ3tjCtVSdWfVoxO+ORJW2HcUuZy0SuxXgtKVqIMyOl44iKMOmASb+QvxPXE3MiXSlWY4ga
3zuleO/sKVcUGIz2TJS/GxFGihlD/kPHaQKo9xCyf1r/gnkUMRwoYbMDHKNTr4/tVBOsURaZuvHI
xPvPyQsNu/tmSZ1VSiHtVDX3qrBtA15UKXuzggr06JNxDn0rNu1bXuTkcLWSlIDJlvlIvHAoptnb
eoAihfUNnOeBPxoY/mRm4XhOcAZEH8CPYWSY3oRw/ZSYfwH9Q/W3NJ0XpaDFKws8qjmVFuDSst0y
0fK9brijBesnjUpCYJDbJldwEkfYs0aNPYQbIkWY7pryg+nMMjEVKDDBgFdF/SgmyAlg9PGX+GbQ
AdoldH3kezdsbA2TUpgL909phTDW1gwFlC4lwbHryn989QpWFlwEBf9TcGCg1DncJeWpcPDO0EyP
BS4DKC+vNBGcoO81oru8DJxFXlBhkfEdx89VT6Z5hs3ZWflvveJG8i5kM2UcDfzvBYJVO7mC7hqs
qqK4ba1DU7UDx3C1KDm6B+iX/8u3mC4AM+p/1FN1oZxsGQ86NyDbTuMUY8oSESc2LlSK80VtOXzE
1umbxWKhmGbvdnm0pdPwJBM10Cf1JrNPFNCUo5PbU6WanBC/JeppLYUFQXlC0IEDxTZV2+dOYIRS
s6R5RAuYDPQPjzV6V/NmtigDC7lwxAkDYaxAyP2YH11kr+u23JAN3AQmbC8Pl0cB9G7FLUapCRrY
kQ1xvYwYJJ6IcA/57TlBKmzDa5/2H7p3o93PHWx0CkO4exmv6Sqn4k8dHWVQtqh5Gea1HebeOcTG
2SsK45mGbzxE00tzHCS5+rFtpG/TEs+Al+0N5q7oRWjvr9o1DLTUcVDJ8WSksJtq6KwkG/ijzM+/
9IGfUEUBkebn4NEWnuq3DyDvmoPSehlLaOzdYk6XSWWdU8PjutT+mlrv+eUUpQhvAxHyXfcYjOHw
0n6xWLdINRVVBSBbWesJqxABfgHpxg5UiXi6pYai7n2VaU129ejmEEOO0C5JeU4c3+bD2I6B5Bge
0uKPCfZ3la3Y3TO6m9/bu2II5YK7FXYG1kI1mAHFLLJ7AXOV0tdzRxKulKoV/u54N22dHTNzZz3N
nS4rvyjH8LfcsMxSlkShGicRW2eRRyqid7tWWzllkcR7unF3UwrMkGTRzVhJmH3kdV61PFtk95u2
KPvk+nv8hWqkcOui6daAolhGAB6bnrX7vW7zPRN7uT/SagSU1ij7IE54D+C9VE7HdSVEgDuuyjG0
L9V2bzT5t7ArE6PLzp4iVZ6NUU1ZCkOErTIhlTmXTsWpy8nWqrBUzxrUkb+bd0CMQROk1Aw/p0jd
fJ192Ub8PLjVGlfd+A3qpEsr2Fmc4839xJ+JyqOzmmqGpeO886285ioMmheOK2tmGOSqdDYpVPbR
GrNjGZwk2duw9QJpbWgxFGh7eDTV4E6ByRxxVwATyjqxhGGEWm0lydFv1hf3DDVemCkRo0zIeXW1
gbW2cltqDPPOUFRYqFVXSlbQY8/yRpOelHPHpGDVnpLPfqNyhXXvGajXtM0/0p7xWusscfLLX+a9
0Vej7Po8ChaLUgdwr7B7km376t8Uc8k2cdi+SecHIYldez3/qatr3Kw3J4O41PxPrIyzRM2RFX2z
oyD6BRV6DrTD/4PjhUeATeIJlHOP+X8B0V0p+9az5xVLOyUY2Bq0Jz5lmbpPAsPhM9egxmsyVt18
3LRH14Nx9KaDdAR70scFgvS8ZN2VY0D9HCrf/YkAhGM4cJKQ2Be/RHzzYHlnWqYeSPLvJLHlfVKn
tqLoBX7eoO6cixdCCOkZKZcttX2d4fi4yyle546eYvTD0aVaj//0RQGjBCLy8gdY4DLbQ+ka7VKz
TiLydbxTht2h+6WMp1xv/XhnE/6vXNPngaEqB6q6bGes8C2RhMMlSYHN86rJJG6FAp9cFPLxaKx8
Dcz8BQ/4FHCJgSd3Ww0TN7zNk6hc4SiRpfcOwBnfn5y/w9QdDq+9Q/Z4DkvIfmJTnk9jAco+LMyr
NTb/7NIn6ptyx0SLdH9rB2ZLoAvLD8gQLL3G69HLbGYX9XuPEo7xi7xumbtd4FnB1raA1YRLw0JX
c6qE3Oujk5NbycFSZjNcdApXt5PvwIKfCibHmw91TiBHQeN4GElMySrcRC3uiST5/OMtCdDPF7RJ
VYjO5LH83MP/QumTMj7c04KBfl81KM4nxANTWXtwI0PKnh0Wn7LeFjX7C+s97sKfWwUcqnpEOm2d
r7JeUDhnxbqOl5vzJ6thOykjCJ6ravZc/er+ReCn32BNDAx4LuH77aOaGon+KUr/Y9RWMxYhSpEg
RWoTsMuTfLVfpukyOxjmL5zY/gTE73xECnCoLEntYgFbzpEzlzgtKr6V4aQnEf7jTB9tNZMYW0Uz
k39VuV3EE3h/8mjplcrM95Glq7CSXMxGjSf9TtHP18/Z/VvbDrV9KxG0XYA+CBpzi+xL8GfQEdLv
eIys7kdgcWp8PpU0xokwGAoeOHCtK+3Jo4EQZtE+JuaftlXaSBPnT+q9WAqr0DHKYJ+yerZDIwTg
CbLKDKbLElao3JqvbBgGVB5QmNrs2WQ1f3+e9iXHKPBsPOw0F6SGMtciX18RZJzRLjHfAm1HJh0b
AmrDd8bHm326MrOGtrOLpHKuDgx/0RMQh/5qVZO7OJ/CDoZkG128DJFA4b0EJRHYh26ziqf3wHID
KLG+1lUFJMuU63uNOe5fO0lfHQ8vGEZg+EnoXl6DLMD/Jy+Dy6Ob3aPHqvs4xERFsejx2L5eUZKs
Uw2NQHEt8kqmnBVn4KnxynQOB9Rf/sQzRzT0Zem8/eNPRnlwlSYh0bRc0J14Axn1xn7xQtn1eN7+
x9QY1kEYGbAVM1kHxrYcLs1Mc1l/a7KjlueNUqFl86ufQEZra8wmjMJ5vEViM+MMDWpUvGnIH1/T
mAl16NsQbTha9mMJA7szTdnrW5Y2Gea3V1hQOJ/FU3OYkqKApRLZJKqjcKxheL1yBddNwhB+Ny+P
s9Ize5uGVS1dGHlPGDCXkW3bfgk0vp4dwzV8MTlpdK0KFkph9h8mtaC+7b7qIy1faljPQgOY5lpJ
5/jmn4ALi+Xfrt/kldHL2wQ0x2GAtdvqUuOjUzDV4watOS3yKOtJlv+IBebhls2Xd7lpmVJF8jBV
mutD7Ke3pOHuYUcihBAEJheVXi1lGt2W9Sw5Vxpvos9g7zXpL/SowUsMhV84fzWBSStJvjUGkhXb
Kfj22PyIUbtkmQMiPU6Jjis2JE+ske9/rPubFS5uxINchSZ3o1Zu4H1zICajWAbVia5FGCKrMReF
O5zbcmT9eWqC3n/WKqvNwKmZgU3SFuym6xiYBO9Qzj5I8fkbNTlN0OI0g5iUm4EniFxaoi3wRKnL
SZk/6Q/g1Udri28XcQppGR39kMV+H6In7lv7rj1MNpEecuvsZAjVSpkDGqzlOkO1ihc3dIBYHKXK
lzIj/TlTfE0mXmBnyil8z49RGMTHt3hOunLCokogWh6mqPbMKPBmNRZqViedcO5srSNBpZEVnesl
lM+jH/egUFpT6i5kU19kJV7DfYz3vHs3ie6NrrAUsqPu/CUnGnZQrPlJkb7JssNc361Rwovy1MPF
GDTkrXuYJS3bq33IHtx/PTfm0WnV2g3VjRp3CmcbdW0+0CS7E25VDzn8horUfEIU8XiMLwuYCOi2
jcU910yCBYpOK/9rgUROcspH567BEqspfS7l76KMOlfsqpCZX6nnqxoMNkNGHpaw7FptdS8dLgnK
oihkRqlUorQQ7RdaZmWOxuDyYZGj5wQ13mIeegmYcQ+IGSEHLOHQzZnIGRILjDXByeXKHWYDozgy
wQKLuwGNC9h3XEGilKRAWBzg/vsypniFtU6+geideiaKGbZj5+qkO117ArTntuehoc2ce4/MQQgc
3v86HEgcnQOoppNh3PNxIsw4WaYHDOsrJVo88NtjiEorVmfy0hf0xhaGwEXrT1QIGB88dJVms8t5
BlvMEKqfmRSaehFVOsBTgowKrAeaJqYP+ky5n4qWXDMzv7SJh7Q8z+Cqx5yehdLoKlxkPhf2FMm/
j3XX27QwqUHivFbbdWzyVEJz4obRlDlC4htkQZzqS0YUQWGLn+jyYjcBf6pSxz0PUwkmOlAS5hKO
YwOZMfwyPp+uPlCm04O2099h4F5OuA4O3xJhCM/oWFv8W40wJA1LRDJCPegig2Qb55PQeEjqWrAr
LywCni0SLXUugn1aMz0FWa8UP4+tQIDQd8cuZxcVVofz95eMYHMlhJ6wAai6tg1nRmHrMkTmMPlz
ABQjwA88hWKkuQS7+K1m3IYM74lvHrViaoRkEYvurpvT0DCrXCJM+uScgL6j1sKb2FcTdSMdARLu
1z9RNMMpld/MCyG7dm7Yl+EjOH/jQz1vsnlpkbNfarnVejUPL7bawiwLYo5G6U4LQXn1wi0ab549
4AcHGy+UVFEZjJcHIDVz1Fwl+LUb5gwQLGt27J5Wa115mU1inQcKG0K0XKDBs5+Wdux95DkaeHBh
4DtAclbs8hCywiNhkHfW96MhPAbIcMV8W54B/XVxYwbWKeUk52Z76PvenfVpU4XoqmfphnT3O0pr
vTj+X79SQ+83qqe7IdFKxq5a61+uuSH/aQLP9gRKpPY8mRsn+CTlIssHOr51vYTHUAWINrlMeZa0
OJEIaj9U+ZfU5fTd6UfeFsdzn0/C54vAat+MafH/T3RJiCjoRQpehTkqcTkWPrRhPl75Bw5Sx0ZX
y1SrzCWJEDqhWmSNgwWVT4puk5eJSSqO5isya6+zDUPeM9oJnZ5Fwt3kuvmF3pODKiRhgqxdD5in
1myD7Dm0L1yRxvNr4XusrvlWDoRkbbS7A0W5W0Jz/sPC9tm8pvdquhY1r9a/y+RQp9bCXbCx4/cl
i+LB3M8ZdwYlyPqj9u2HPVtcP84qFS3BwMPc0BjzudESddNd94a4Gwm/azF6lCbbBjsonzjRj/pC
Pzmk5UFEkZCoRnra9VpzaYHTYeO0kCJDL0O40uV1L2xJVx7y2l1AoZfA1dD5QsifbXA7ohXO3vu2
bSpFnyMfa+3NBGy6OLANd+TIMIcZC7ACjZxMLClCCkd9Sl3n2uiJuPQgN3SnYrtkZmwg8VSpY57y
5PzKpLKpe5TF1x+nW//eXTVsBBTzO1NGm//iwgqCWi3r38GZJMkvu31wqcN5YjxX5rJV5ej2NL9t
pct/h0P3FqTFfr5CC5Qi3Wh7BNwTk5VttvKp+9+Q9GLtgDwbJggB4YpVuvkDVsIKPEp0E/uvRImk
rGZwGXSP2l13fASiNidxb2c0DSmsg1hkM7p+HYPCTIN+QCigP1fEimvOe8AmSsLVMsATydBUzdab
RdCuA8w6eKm6UpRTODzE9ksAi8Kjj6mE6J5ajMz/U0mqO+o/T1GDhf1P1yeL6v/zZb6H7sa92+/n
8iBUVMlnI68+edK/D9SaF+2ACy/0SAQxR3BW/wkLh/GyTJxIn7ko3tBj7PmgRwWlhqiMBgDaSS4t
4V2X2lAz3/f/e2ZFkwvdiI3LBAy1BcB/0Z4wTBFxUjizEi6rKtjw7asrY6igH5SA59mtfLu6k9tf
vchML0vZR0i2ArxbLYpQ3CvnPjkVnnploS0GXUvLY3Wa35Q9AcmzZvbxA/9aV6XBCW8fiPqPoXlS
SPrRNZYqXg4O6EsXdJCyTIZUYhC/MoO1dGB91Vw4YmygHAlXrZTCv7fz02r1D8w5X5ov5SUEwm5f
TshM1NS8j85LDRTmXwjMHViGJCBL6iG8F+dLi4Dgdv+x3goH4fiRd61EQPrDx8yQysXm1ik6MNYw
YVKB7HJkW8H5baO111UVSk87XJc9jFDsZG4Iu22ZO+gBVgSXabe7iOpVyVOS4f/fbIVrb2//JQ5U
SGDl3icDAuNbQISRavx0Hzf5dINx3sbHeSzGN2/0I/JDJOCd+36R6LKBWu6YFjTjS6A2WjUP8jbL
C7LPJYDST9mFZulbU5EuQQTUth5zOA6Y2LCxIRzxU2laTUaDOUqaF0mItUjwECXVsqH+bsjkGAA8
GE9mFkCryi95y/uWgn/pH6GNSFV/TKKlFyuLu7wHYXoKMzohqDOcW1i0P3a7Y7dn3TlhHlZj8Hdz
DTSYquvhOlMf/pQx4TFyXnoNBHCve4n8/zA0EUxLfrFxloMkiha39VsrUIwQ0c7Kv2NyhI4x9nl2
rqN/25yuvecpPbs4XC9b7lQM6H2e/PxHaOZBR5nT0PvNlFSlh2keC9Tcn9+mkNduPrDgvVgsYZlF
sCyrHeATVaP4GX7zoMKaELPTeoLH5yRvKSphztsXjnYE47FT03LtmEYcvUg+PrFDzisPusGi3rch
2nYyWsr2XbgXuUhWL//6W+Lmj880PclmUnykhRNAD4X4UNEk0ZZQFI/k4J1KXu8nTqipVIYYqBUU
lRkuL3+Wkv0ecvLHIz15FqfzeDlQac1qgdG/3YaBLePOErlsZq8wpOK+wzcucEtII6aZEmN6f+Td
e9OHxJGO6FFSZz41zojVFHlX5wa7OPOwGuTL9rQ07iNlRG2gwZi0YTSlvUaIUnQTBZedr57kGzIC
W6D1GE18gSxujq4gliYiJwh+3UeX7X8xo+qqc4NThoe1qpYLXcW+zhQLGHgsU86bENayGRQ27pzE
tOdgo4jiQV+vFIYa2TecwVq2b1bs09Z9z30gX8YWU/suy+tuNLH5bAb8M1b6DRJfRpJDBlHOxhuc
sEinALC81CRYy/NOtWeJGcJb7Y321hmwomgEQQ/xMZf1T2fMEAi5YflIFDgXZlLoKds4G8TTip2S
FgfYWcLBfrxEBHoT5/3b3JXbgjrz3GyOEsW80pfbH2f6Ne8dtKOKSey3tRM0Tb6BETTpjTTY0EpD
JKpPmdnhJCkoyFZlw0SV5VXqh1ayci6BZlraMlT62/34IdBXZjBIf6j8UlB8W9WKTMMmPnu9ScZH
x7SkqPEjb1SUmb9Z0iqkdMeZyNnF8eeOmLfUz7324MS1jIhxLKU0SW7mVp+Q2T+aDzICHlwZqrO2
uENmfBZuw4XOj8P8NjlI8wCmdae/UiYzAghDgkT85F0hfsrrH/ISYR07r3/PqCocFQvHkc4bKcIj
rfNw6tos5deqKGqMUWeVSQpHC+PN04eumlDxZJPpNA2dYBm1YEQ4xLpNnNofBXNz2BkTbeHfaBM8
qtZf3RIy2A9qXz9y/lL32kD5XcEBCaSsiIUrJ5jiKNGM7AVl++RVwC2TEiZ+glIEfIqvS8dvGXlI
uGCZQUdMDrgmoxAHCvNK9AKLp/A2BgYeKvq3o7xrz+vlpoHJd5uGSV++Exqy8V7fssqhm9YBYjnk
CRgFmzvA3VSBd+I64U7N0b2/OqEwLG7MJxehAUOut1gGIvsOltinD+EMnWp9c7559d+wkf/oO2og
2I5LIV7FprJQSMlklYXUJBrKPKk7RyJDDWOCQm1CQbDHLSMEIbwn0xtjiUJPlJx36guVRHbuz38/
4bxHXJ5GagUDagy7TVs1/zUGFZaVmogM+NXLV1RYH1L3OeOYH66R9CQ7YXW2ALMF27Vo19UctRu3
96vUI712O95aymONxholH2Ev17otDWhQValJgiVBrcM4wYncx6XX+cgZwAzLCsN7j96/QIX2TRwZ
aqne3ZnYIB/Ic0dQVD1qfSxlrIFRgObUgSo9d5ow40v+v1jIjmr/bRSzCUMH9KohrcZFunSICb1a
CKlUUZb3jcMuJlBQYHXlT3QGHzQHCYlnZlNFbQ9u3ZBjfeINLJg0oBh+bp+q7Pwk7Tmoatgn28y8
d6MDKkayYPiUmrk9nwA2Ivqyc+1JFAVsSXi97ItV6qjg+JNIKzCfUN6ChQOmmSBpb8UnqlEbXmd8
lWG+35LodlWM+xyxA8zWjdB3FmtwIGL5x8UdIO2bvlGv6RzeBrqEtRJvVvUnrIJfhtcwR4t05jMJ
npZbU0Adkqge9fpTT7LH7B7xxVCIogZQps9b/j/gcghUeh6TMHoyib8hX40ct7bddprTJoUop/sN
RzFVgMhHavHi+stxm3yhdzfB5+4mrZNpZaY+Co8igznrL3nOD8lbvtrzfXL+IlemYB4NZskxXJ59
yDVMDbKeCrui2dnXNJS9/khS+dkagBSIuRfC5UsYaqj7/pQub84TXtuIk5c1/T1z4Jn9qP944lHg
n9pWY5EqaYFxLtUlqVnW5RA6arEKyNxxoXJCefgLsSos3uj8PXIlGBV+9ICn+a8mwBKguKWAm3By
OD7rC2APd1DecrrD2LG0sOwWSijfcgW3Rpnii8BjeMKOrGXE9RwLfn1RVkw/6aSp0nxv07EYcF4O
rawd43Up62fHjeExrdz7/+Tyq7l4MTChjx+B9rMwD6GsihUbVj2eUgEKFopTcV75A6+vyRFhJUQH
unsfegdh74kVG40uUjWRaABRVLW8AuHFc3UAMCkLv0ATHSno0H7udqjykdxiecBNZePADQ1VgtpO
dUlQlpHiieNL9dlODBd/O5Drn5gtx66sfVgNdyOTVGzqchnEVVhjN4QgsvxeEzbnD1t1EdBkP3FI
ri2D6Xjt8/m99NCtQqM4x2Q8GHcjSjsKXKowOv8JDW31AiC8CVlDSdUa6PkQnGjdpaxicCxdAKAv
Tt1ZlmVIkTH3p2O82muzSt1qMFUM2AwxAjGKdHPs3FDZsSZ4/RDYboJG0/ZdkVl508RQRl47ey2P
nkzDVV2pvqdN+EB2ngDcFN1+GMkSRrc/565aTMCN/CcdDZOUpE3b17UUXGuKeIkzzUpS88rRAmAR
6yA6ClkojmIhHTSGSi0n5yQxo1LRx0VgZL+nFGAOZWm09mLlK/NwKYI3I50bwS9AIo5kbygQka0J
/Dt/A+HruXVDNBQQ4Mrfi/sDv9vY+CXjvpQf3CLdETr/Zz9jzmlwuRp/U2WTOXl2G5jOwniaLNvJ
BAe/DvPbahqNUWKLPLkKZiIDkvEqmG9my2+4Q0DfXfR6EKpsEoLsWEidOAc7Wnb1fYIl/Mpe/j0q
GoqMKAH71HbXeN4XcxqCUanx2YCtZqBoLzYkjEGcS+0NLhecr2cgG0Z8V9zTFedaC8nkjopqyc6G
76l8QSW1YOXFxRqm/7zmEemUByrSRnjuo7z+MNuiN63ekPa1WQYul6jL5VEFZDzhMB8FRb+B94g5
vl4kvEg3i425Lb+fL7Lf6QuM5QBJnADg/vPWItcGuKpB7qzJsRWIc1sB//piSkcBB+IaGfZjyZ6h
VA1ow25U5jTqsTEt0iqnT56qCCgU0Z+lYimI9U96ezpnh0FeGgPsLABHD/hrC1JQtuVHpb8jzIrJ
h+XCFg3Um9ljDzQ9bXLiSBkvDv+HPocXafqiQtXYxkdl5KG19ixx/miMD3ZXU4eZv4rx2kyPZUVU
OVltlHahURMnkMJkTQ2lIew3+lYuwIaf8bpDi0AI8B7Yae0GQRxfErRFYuUzTLPBkxDbRVY9/l32
6Db9nijYyX/G17yZn9C/MP8nRumDxSFmJOmLvVZsLNXQsq8gU7NuuqG6lXxREfjK0WK001J6w2CT
FHqfNFwa3qVrqDJNM8MPOM6iJRHW3WUELEJDeAWE/1RnDhm/w6O0Xl5r6fBVDEhmO4BDewYUMNHO
L1lDBys0VN5MjSgYTVre3LgK3gOUKwn0n96OZhL4mtNPLYbo7JMpthwHIWeU8WIdOCy4Hw4LJT27
0b7DQeBZaQNkEDbOe+F8bQfHHwrCBGKt5P2watqnAggWlM/M0+YrZ6x/w1YW+q2gxoxAmsBRxUew
+UvGVJYXbB1UVuhG+dnz4mC5IKyAQ6qcLAe1Soe/R7PdEPNWoD3nFRDI5ZV+30nJAhIbB/yHUffC
9eooBmjXfUbsaT4pcq0FkPiP2iM4MpgJ5XYquVUkIrS8Nprh8nNnXJJ2CuDoS7l89QZUpNtos5nV
tidUAmOFcJ202E4iQOKsDa/UwVVuYle45l0tqesViM582Te2ym55acn286x5Lz1RlVKar3io5ODJ
6KOxx373K5TZAK3Cb6gvlnRpvGKyfvDT/QMjwMXGruyQbT98axp4GmwQhyVzfvVt/LzGpITw8AAf
WvUwO4L+EqUALvHfgS3QCPvqv2uxoQXObr0M8hBTr6EzBpujybb8O+sE0NUxt2Udt70wNopCSYPB
pF9v3rRphrT5i4FOgsgJRj6dKMdyV1b81mfm0wsUfoHRhyMysputFyUvk3ELtsX9Pq4DEYpFuPHp
rG2KykrNzOYiAPnMD4mB3e0MvL3f5fURdgUIQpYhBfERcf3zkMQTb9IaSTyOp9agITwX9jEwf4HW
fDWYaSOuSLFryCSa6a3H9Hu1QZSeHNsAQESpQ8NEPiy4wHNN3HRTAQEyoRItsobEzIP3ZluG6XDZ
SNVnV6eRncOw/TZ+C3FekbHt15cCrDO94U4nqHDEoAZapgc62W2h4p5n52KPcY1de7bwQd1OFHJH
0BPZ2K1Er82dl00i9YsVKD1uot2RdRFvkO+fJ2pCxPxUdsUgdy+8dOPCB9MZjDZH+6KaHvdcv1Lj
QM/TEXsY+mMuGaA8op+fWuvwjFDKaJF1e91V/ujn4lGuIyGRKgrk1ZjWsNAsiN8gSoxs8e3kjs2h
zanDnZ1sVu7VHFed0jinHUpClbxawGHmFktphPbanHUd1TdpBlz54jcaqd3Dp6CUJQa1lVh++pVJ
hXqmJG+6wbGNwoelUTr0HPBUoqGrba8aPkntKnhrpW1OGUkQlvE2tELKJRgyWtt6LaVDzU/Ns3B3
olEBQsaLUNv5DuOZtDrOLQlwrzIzq/p1fUflhWPlb2LNSh9iR1yjJqB/y75aeyUUJ4qbKZjLBXxi
5X+TEBrq6Dipk89VwrD3yStsgcGSblSCBkLqQH2FlCl7CUelhBnXqQZc76m0bpZNLVO6JRn+155j
cJN3+D5VDbfILmiQBgag+R1ZBCvh5xqE0lY/Q4rMbN8zpHsSrZQHYY7PBramUUHXQnwL/t89tDeq
U8XPdMiyEPxgbQQXyzdlS4MoP/xKsEChONEKGNcCz0whxZow6TVtGEl/1USawByQUMaGwVseW4wZ
0Hsokj/wBgA+wFx1onK3pCrTlyNC+pRnjhyaYn+QoZXgDV7zuEiRaSM7tm99qAis9qiWk4OCZnAJ
3B4qKLINo1aWxMSKVuYRcUkzcpCTC5Ta5ejQCuHWuT8LAICA1f2P9mrahXO3MiI0+NZrh32nI6qy
8VL2wW/Lx+myKsJKw20euqlFFdadHSOjjnPIMTmj0VBwWRTIOB+uJBMJksN6UhX5Jo04GXhV3Kbc
WpUQblmmsrucicO7FzAIipmVO4dPLYQGOyU5Lrb2xP3F8ll/3JX+zn24PfiAcLFStAm581tHqsMN
h4aZ+oC5Kwsm7ChDqolA2s8wfxnE8ms4hJbOtGDGQjcejxMBKrR/Tl6T7RZcgQhquoU+uTIy15dn
OGHBB1ySXBSIZNTYakZojyOaNlOTxPnT3Xi4Z92p9tTs4/8ys4PvdH5Ez/l4RHxwKfybLC6fGMN6
B43zFrOQqgtmxikielXK4fNZn2C7hZ5jzSg51K4+yHhFTi4hfvUJ70hLpNY3QurnHxqGy8Vk7M5q
aZOzYyWKg0VvKGxpB8YHOldCsegz0DXGjKV5h5u8srRgk5ateLkyC20CeXQGJFQC96zo0/hl1KS8
Y/d1AfSaVSGT3IO9f04gZXetVWp/6Hs3lOzXIY45CgM35HeWLlA9nLlTYdT7bFYA8J2wdIY3R37C
e4EwQ1Ws7VwYSmpPl7WacwDCiv1CUb6RDHeN0v5uDOcUPbqrsDZAXOsctIuj2fFQkLEzd0u5/rRZ
HnE11EDcuymvTEdlTQidXifIZcAmZf0MMoy9YmqcDtMqeUQsXWxNLhb95VPthrRDJttT2H8q9CLc
y6T23g0L24POey1mQn1HELrWxHcxh1R3YkR4/+o3lqj4HX8DEzmgfQl8o8W9Q07gwPxnmE0ocCXM
SvUwDKG18ZaPgVseF/DEepwwopQ0YHbq80cOg1vk8EWhTwhSYYcxWDXj+c7eidSvBB2GY5qcXuiQ
OiiepE64GV5Kb3GllUDaHFTCcTNAKUPblTjCCF39bpNCTGOYu8ajkcI3Cq7GS25RBg2Ye8YuYAfp
PFefXzPs3qh+ke6AfGKWvMQOOMxnHe3lk9I/LxWPDyzFuErCSdiJkb9RmDUNuzBQ5cVC5JvznZhV
OVAyaJeYwCkRQ4fk0dA0njj9E3tfrMSLmT6ipVzL1cFFULgEP6Fv7ddgL4OrAr6ZP75M/+O//wOy
AK1OgAC2vdd5sc0xgptRzKh4gu3HOt0wdp7OJxEpiaKV33WbNKtZATO7eakASAeXUqQs6rjhw2Mu
36+UcqT20bAinaKPIuVadI0aHS9VUou72y+sxte7uWxiGnDH8P+tLy3gKCH2FTVihTgZEH5sGO+e
l0IeZUMT/udgY59S9xcLZSbf4pyirasbSbBdGTBMhaqW8IWtS5Vr1GjAnZ5g04oMDrbnpXr7conb
X/LEeKj//YYP4uSgnW0xrrTdjivSpv4U7+9nHCc+MmjxPAb2PEFHDP6IGjN84OSHOfnXvmEwfu7k
EBp10+E4DEV57DaDEeo8keNrWokh0gj0kZmBQ0ZMPdxWk6W/xZ460GfatO845mk/eGesnNVIbcsy
D4otJatDLPfipWAuyR3ofVjsX7W7wFAAENgIxhG82XtiPrr2WMg7UB/8xlGhNt5i9EcMKbagUrr5
73SyUFMYJPu9f3JFbUfUAjB9Dv6R+nk5kzTRt594+57zFlkUus3mc2u+sBbf/VkD7SqqtdclAkug
sALNWB3VeXuDgU1nPcLe22Dvan8KbaIjyUL0TkX4ES6cLO3FrALgJNclvhtyl0R7pkGd4XiAf/oV
Rv1zs6DEK4ugVAdhnRzVWD2nR4Q+xgtSgov60S/5Fo6LBzjKhUFK0yKUEyIOiWQvDADSRIfAwhvm
IQ3Y/TIrBYo/wLR0T3SqNZzd3rcJFN/Y+eFZl1ihXEWntC8xagGsZ7+1wGu5heMYg0u2C+VnTq9n
iW4gG+Udk/mQ+oDA4n6I5KfzTvjnoFMXeDEZ96AfLL+utZjV24znUsc+17mwpAHc/lAFlSDSsLsp
eFp/9j7QefSW3w3fSUIko2KjjGEbQKlOlLOLtPHTi3SqcGCHw7BIPhQlCTfG753bQ1iKPt7hZwhh
TJK8cSWV8VMcF/2R4pMS/biyYcyFyTphrKS16uHlUkTliwgBiDZKcB53mLne2pnwvyq5/7cTRpic
4QVTEiqL4pxpW8udSeMhDIp5QGfo5CR3eve4iOuTNePKNGYrQ2FTi2nHa/O3WlHne49VaOympca2
cbvAlAtKeJiq2Re0RaQAxWDQgDx//fEJuPrlQY3EhVX2Exck8J2+zSGEcAS9J77nl0ZnlTHyuV6W
CyoZ5/3JBdpJ2Hdpp+tXFwaf4x6qVj0v2dgHJ77hAt/OkCviRCu9ODouVs+ng01s5Qie2fM9jxh9
+cfCeVRK7La+F+1dxRIVswMKLN8BjhKOBTBEP7+54BzfLTGbUAHzIlUYsTYPAk4cahVTR8LO399M
BtHEDDuYLrBT73jubPkOpdf96ljBbfz7s0f/FqNB8MBcJOHExg2wHVTk+He1DmPNggfHBn7o8Gcg
0/26wNz3vUbBKenUGAV3wt7F7ogQZQH4ER1KlR9YYaRV+SxpVSoPNbSljQsIOzphLnHaSIB2CHmB
q+kyrD070NHuRRWaxac8MVqXWw43YCsysHuLqcfgxEshT85ThLMkXNlTz2nDuvcDG7Ar62rHaT58
E471vYIrW7paWc3zWFKarJczhoCnI8TPDPTZKMKsbMUUo4lIQWxQLsoQWilqFl2pBqsOXRy1gql5
qVJ1ZEEr4cLhF5luax47MWsAC8k1l/4WOfKKtUF4fARvNZRGIFOsG4hjRyJAkAD/lWnfZazZwIFB
9OMlhi2LG2Xf3+85CZNzD6/qbhKcxJhwSRUIikgiAkqhOJbbxbEU3JiyDREmDeaEY3YvtYxmejoz
gyAZuAj8gxwciFVg/NGjGTKC8SwpR91XbbjWFUjZD2pKwWNhK/1YXqwcmABtkjsOGKj17mhZncjw
vX5SKzMUgb1ZRyJJLXzFtTgTt5GpDAUvppxfD/8k5XE+8qIPxgBNdu1J73BbiFOijh19u8xIvkmB
IP2CoMVzT4KeN0NLSwV8alY4BZx63WcnEJ4sisnXCANvBQ1fzsPbkBni2KPQzCqSl+s1+nEGlUYr
48DGiQAAVBaSLpi4nBiWb2eDgW1vz+RMEPMbVNX8BAHhr/7j3s1TN60SniJaiCsPW+dP3XmsMmpF
8dTw3zakJ+LTy4NCUy5IRwSdG/JOgHoi/J78WsrWKaWqXKLbPtak823YWSsTMwabdN2dA28zyf41
2PVBsSX+VOjNay4gSnytUrh4P8nAjgrygPN0/oaryTIk1kAFRmBTOTbIp1V6yR0OT9yd9MgazToR
6AV+KiGc3fnB8fGTkY7bdttZE8pzg4GPSL9tK20wka76rGOwqRnsBp+X1pbBYSAo2740Fr8ySjvf
JUG2ul5CTsuEcPPwEeKqNdy1vsfebr7/V/Bb5CfK+IG7m3fWtNzhKKFAUgWxNzyUN4SPsuJ+t0rH
hijXeOqvrHViGN/kFfb5d7jGZcbR3cAXRoRA0Y7o852iXLB2lFOYhXGAWqHd+z0MRhIwoOj0mu2E
fx2l63e0HF0V5Dh37plsnqJhzaoRjXaUMvLohep5vkBpo3AgN0zGspN9eomM+GbmBRqZIlN7Ei2D
tMA5EDgp3Au+jy/4BCiJsULdTclWmHMZ5ZJPR/wyfyfEqqCJQNxpwr4GO+uOzr3W1ZRWd/mRIZhE
qD/93qI4iVSc7QvtdMAhT537tffK7VDQ8qLqtzGICpDGDbdmNjpCusPyxEDOKM7yJsL+lB1pnUF0
tfhh9EuOyqjuX3+LQygS7CTDw+3Je+MWKUQxs+qHnDUvkefu9DfR0nfMg10Lqm41zdVqoGpYkQzp
bw7pzu08WgkGbeDvp/NpyHaNjxA9cuvuUWKlrLzyUDkf56M9vodijIyXZGCe0CIrzVvLeX5wXWW6
TWGfdaK8HaymmUP2WdLNOvJXCSOGr/JIZg9Dp9q7YdQBApkR8d3supKxJEOXDiZLGUZLA6u1XGyh
IZQDTTQA1ykqkoJdF0ZktCS261gsGK0U6lhD2GDIfmCeNM1Dh0MLXH8Ipb3xxK+UC4NP2pebnyrr
7fWOUBy4h1qAmAbmTDInqnTYweNbhhewwr6dcw+bkNcOeIuiruRBXRTj1QoLrJ6Dvo6Sb3fA8ccF
3kYtJKSwEskg1KReGRYKiJd89lllvjhopIVZhClC3KcQFHKxVJhsCIRCNCy/y/uUay9Cg6mWfztG
Tag8SYMJYcAiK8hIPMNlGRUCYNEZA5TiCb27Z595wlvR+DE3lHFRvLAyNR9sDcaLV5hA6zn+VVAX
fkrPtPRJkVKhalXWnBEWmy3faoCocHoew6J8O2q9C6YmFt3XABnVd/A4mwHDzIk+aKtIMFZGrc+t
k7k+dVW0J++JKNj/FA5QvK6Q43l4ew0/pVl6sO2qQHv5DQz2DCpqeBpE1urNTZQyQPT1gYlE4ves
EIagnZvjCew5k7lASx8cjC4NPFuU2IxK4zO+afsthSi+lswaU4B4Ka80ChjSIRz7F/uMn3Fvmh2U
OqEKeHtHHdAJ+3YI6BDdn/dz5WIA0l3ydB9VQPb+dfk6m/G/6Rjkp8kbRd+TDfxUL2DtxI96i4Wh
J7TtCFzDUh63TC/qPmI3exVxbIMKQYAVVBNI7ECneZuxufOj0DsYpLQvG8LHOux9srPx501fu2SL
1jTtNOS99aPz+7qmROvMDp9HYaZkYY1llVJ3klxV63JaxR6KBfWi2kYg4EPk2TNKgsNpz12jf/MC
jrpmANU4KrH8t43W4L7rhP4jdLqzXkStT5VSWh3F0auX5QIIUAhteD+a8QIiX63hSNGwbiYMbiSH
fq74//smziorzrQf4SRJRHB7TyCvIR6NPXHxOBjI+fKeqoQddC79qtTsRKn8oNVhEpG5Oc+KMEUm
JJjDRwShfdj56NvHr71CCJVf8/DyJ78KfQlq/QslY9LExM7++DR6lctBAmXxjNKcjpteDK3D+sXp
BEsZ3mUQNUY8ATp8NezDJ/Zzo/2hlek9nYYlz8fudqHg0L/VR9kRzDay9iJ0e7xQgHLm05SPws+7
ICn4o3ctim+7t8YdxA6E4QiMT2O+nig2GbcT5LEXxLKJ6gKL1Szy3VL8IihCRkW36fGuZ2ejud9Y
1qhfGI+eN5+NAG5Todu0gRHCBjhUKX+NKTUKXfWYkpvXL4yC4LtvSHcLZk/31kHlGhR0SRYgwwWZ
d431RavpqzsDniwHEpBIvqs1zXwaGsaaTetEP7AAQEq7gjKH0IdobjCusMLezdQXktpKgUiu7OnY
dbzpDpjfzED+jH2KcKtZ510CwYJhMexok/yaTPwbnMPSwdB1TyiuwcPQfGRp9DZo5MKIdmbvRAST
LeQEI+p6TKmmXxVoISVgs5vchErz0lde22BpiIxdewkv0ZiMqhwEipaCZoEfGPXyNxx11LvsEDgu
mtyl8eRJ7aAVFcDxchztgOhGRdTKkg85ya3Wwkrs58rt1+c3pn3GvmAXisoyykLuE1sALHY7HXpH
P/j0FMegd4naE5JHOWVGxYm6Xq4xH2dbaaXR8nMMncXhBJt2Qm5MUuYfizUSToEp+7AI7UVeQhOE
mK1IpIWZbQ7DIEGe+KabtuAfIqt58Jl+/d3jcaWxk3ozXZI9b1R+mkt/kWOCmI/rS0o3zJSRx/Lg
4PvG2W5DC+2bLGloOZ2jWL3TR0GGmWBYp/9S0x4F/t3hbaMjjhOdOfcKdAdVycH6KgbRVkG5APDc
2Ht2jXDiyIE7EKYv1f3jPSkoJMxJS282oTpRwUrlzigkXkTwuHcXdRnzHTaZ2kn0v7I49eq7M1CI
6bbJAiwvV7reAKJB1ljmRspOYbPVd7u66ZJ7pVuieYYZP/NYPvabZm9TzOrzEudARReT3igLFn1w
v6BMOXXkjy+KjAivItJL6NCj6BdVR42ql1Z+jUgJWRwMWXIbTWddwpBIwCGnDf2QDoTbRinRTWqo
D9JhNDdzGlBJxySaY7GPVnN1xkL1MPzHBNoCpqwcjklkDviw5lShLMunEBJwr6997a4I503TwU6P
K7ISCwS+KC0FBxG7fdwxZKr9UDRQWvnJghYm9QpNdwmW60Da+1QYzNopOvbxYZ62rGNir3GxFTP3
F8ua8z5CTE0Oc7fDBvdE9ZMe7rgA4isl/kuaZiOJhb4N0jWSLL/OKUo0QdijSTu+DfETEPM8+KSC
Ud/xFHMFD0Xfy8OGiWqqDkz7/ykhQ0xMRloCpzDJ7XyOqx5XapNVGKfTgvBLC1Xwi3AdA+sQh4Sd
Z0SdJwCqbT7gt/p3ZDGVFZUVzpOdsnnS698+VhOAGyPFQGC5C1IRdHIkSmvBXTfTTbYmq8+ugcm8
J62k2P1K+Lc6x9p/6671rArm4QL62ae2rXsewb7BYbf1hOvNcJJzSB/VUGEEi6yIWA6Yemrt/szr
+VO5HK1zkjKrfGnWkUej57IQivJ0aS1Z7E+ZZBiS+fUxAzpyyG0jiCRd6TrD91eKlko2oYnBmzXs
6jaIGuAkJsJyfIn/YZaGD17/WK1LyFb1WvOJIcuy0uMZutCY7puvs/sBwqoRG/kb0IWcutYTV96w
jokTjNSBVaOtKBrzgsxD1yTHvhyOC1HrZpQ9x3+CAtrVMmbeqrZgV6fPpxIxLz3yP5dpXi28zWkf
aQYXs/CGXcTF00+qdp5IUQhHE3LmFmouQuJyiUv9abaUYcc/zEfiVPmGrr1G6ax1TCGn+slW3PI8
oNaiZCoxc+ZkrvYFwalyv0dafZrQDyaMdLChwpf6GD6DyGoFC6iDPF60/1uFw2MaMLDWH3qKhlyN
useu5Tnm+WVh2ntraBqPLtQrj2jrSTjQXN4Sv/bYdcr1uIWldn6Yst8okciUFdZW/1DIiKDgGsDY
ShK0YzNXA+jh8jP6MyAjsHrLCXU2TweAYoI4grZbz3ohgtW/zs5HqWYUUz4mLf0vO5Rt5r4CiIrk
cfMQ/Hb2IcuePnZaIk5lw3y/c9iovSJpim8iuWrh3EJV7yy80FFuG+A255cZtbZwzIMZsR2VOBfI
46mf4pKwsuhmeaaJD/qgEZ1CkQ+7E05gQE2emoNcsj6sYl9ocyalwJTAHwND7ac0WPcycaeuRZMB
onUR6KpbuMXi3Uka9xDTfWnN7sfOwX2xlE8UmTFk5VaYJMOVSGsf/WFVIrTwQgTinq4WQbtdqdXi
0XajsVcj4CqNz/TvWSXVXtry/noupBOa+b2YBXLjjaFgEI+7HeTvUrPZBLNniBOvA++h4JR8v2ia
VW4siLOaPw3WJ1jb935S1VUYFsfbD+WN5Efrhr3o8E+9OdgtuCrcZT1ufq6x/OGAP//c7VReLVG3
5k4jQW726CVPX9F+oAZ86bppey2IqiKoBrRK3OLy/MBuDR6NSnL0vjtPXNOIg2GfnWe07g3s1DTs
ttwgwXX0TCvqFULjXx7v40ZdPJ/54BJhjWYwVZ9GjNVhm+ynfH+h2PQHnBq+4Qg56/nwFJPTVyUf
6IICyJ3GvEJsRAhgB6Lp5iipD2/iSnKAgBbWvXe/tVC71TbsWvdi2AT3Utp6A2/xqog7CBXBWzh8
lOh/UezWqFKubc+Gy80UKxIyXwyIsTT00w0M35yIHQz9486RCTcy3Df7e5/nkm9eYjZpzN8hlfiZ
rPqAX5KCXOi0LWfZFhUvj/uHaFsdjxUh8rdbu+9ILsHDcvG8hFOeceM9n72XWofwv10RSUpWngJX
xK8guWjySKgRwFwS6F0BvA2y5fFV3m9Dc5UknBfmNo9r/W7OzUfD7htC1/qnmd/SlvLCF5Bqg+5r
ccmIupI9RoZt/bEm68hm140UybZZqNS3dKFGuMm3xpGo5PyP5qdoax5kLzb/6suiLss9/zoU1Ed2
w9vzkTLVtk7AqawMrtXtmvua6hXvXgeiv7hQLSSqYHFmHd30jXk+uKXwwsBobdduOHzVlgYcSCQG
sW5C7tTEUdfpfbHmw9I/jS1l1JlKMwVSwpTs618BLllT7E/NU3GLbz8sgDW6R8VGzkCjueFxfvYq
0Wy8v6s8FeXNiZGuXa0cR5UdWeyo0fsl4o2nRbvmJbX6Rgu1USuMoROvKJ22dF8l/K0YVGO8jveZ
BfS1/LZDbQN0XhNeA1wEEy101UQEVGMiu0AQzGSKXMYU37gxnv+XNVqTbMMJCYmQZW8eEjKlujt6
2fIdMcHJuraW4695z0XswncWyZ79u3Llj4dmEZpfqIT40e2EUtSjgQWQrQOJSyl/oFRW47sqAbtm
b+ZPa47qU4bxAipMSvYG9LAwwoo+siLtIP2XrFNesjh6wc/ThDwN7kLT+MaY85yqGLNiE/4HCs9N
qzGO6R9yYaYB1F7jzd25qItMK9kxqg1z9UrLWy80Vik4xKs4VFF+qCLpq3v/qEVKnR/CEUNXxa8J
4/5kX8HyK2NrqgI4P5CPQ4MYA7J1Zu+cOEB19h6oQafwQ1ZyVeQlO3/I2xQ1IkHnpU1FbbSmx5NJ
iJI3fJkMdFpXJCoXhGDjUtukFxDMJt1wMz0XrKJg3abCwvc4jDXJgPtmpPxF3HjVKKxwRIAiFBUg
BSTv/Bqg2xWZMjEiJcBuyVV9eFunkTYJ28h4e/YxJgBICJc6/24NN4moOpVLtuzLrDyKSIbq0DFW
hrfFDwoHnGTQJmfUrGBc/QTThUK5T3OHkNEtKqCFB5WsXLXTUsxye9zE7psXEaZxeNuFMDUFD/IU
QAl6nnI0wsXeffxPT9U6ZaGsIT4x5i50GU5DcF+bkTi2iQkKWov0RZ2KD+4rywD2ridjvqHtIiq4
3bfNTcbSVJZCvYjr/Boh4K925pQbADGONns4MJtvwiE4YYKh+1Wu9W6L/17UT86HWWsa2R8emMhD
toknOnOYhfFu6Ks+zU6vBOfa1RvKAx75MCU9IbZBY4I8xECTcDtryZa/+edk5mCMiEohOa9YJdjs
e8/uZ1PDqjsqyyOmenyVORdC009JNw4z66bAC/SwrUp6zKm31Q3Aypu3DUsgFLZJ6PGwYhaaf/jE
5B4ixrZa9wUQuPqpmagvpqirN34tdkQLUR5t4dCRWmgOunCDYAMOp5+LGULB+CGdqh8VbbpUt8k+
OEGrt9VGX5bk7JQ6zn5hhInfaHerwhzC3FBdifUFnkWI/vbeU21jFLuFVKfNZQlwsm8fBsLYhYnq
GqL2sw6aG/IKEmr4p27CY0tTTarEqzB4n42SlQroQpWcjCKGf84i2SWMMOHjEMrKCtOORL4bLgin
DOOW6UrxMZ31+BhuI8NZrmNa6iEfIQ5bNdv2riSmWI1YyQpn/ACivIpmOKb0XInIrT9zQAUFXQn2
h4zgnah6/ZQvSoGCTkio6UX3oT8V4wj16ix1VUXCWlgmVAh9pN3xf00FuxnEb4kE31hXml1pFW7O
3orGbjIDbfiUidLVu9BU/NY4NFgR5K13U47LRUdR5ZZ4gjXEZ5iuWYACHwFW2kfJQActtULZZ+Gy
TOMJb8kzTkBgczh6j0VxzVaBxwpXyfgarWVC8kgcwHryKKncjlawitPZPPeY7bHyrqT7n6WitwOi
Y0OI7bMsVQy39QOwb5HC9So/IemG464DGQD08jNMj4dfBL18+COVU/vqGiTFdRKtkxKMrFhk6ROA
X3MrntLotBsdq767iJvaroAcyrHl97wLco3p2nwzn3qyTVXV8/XWN+8w6ALF/5D5Np2xsNQGf0gB
NklLsK5g2x1nIsRgzl1zTY7GduQzKy63HkQpEiFQC7Fwr/gX4H0LlTcffQqGfitYHbyAwSpSH575
iWsvgDJunzvaa79Du1PcSMlXSmez1FTFkDxK5PUkjcTUiH7RMBciiO4AsxAZ5jNh1/4Nrhlt6J8w
NzC56PwwtP/Vh0RKVCUdPwGSilKWKsZPF+gZpgyu7xJVM/LPxp4OOOSeuOI2+kmFmUuKlntpQdyj
LFyKF5HYy6aISyi5xywK6D97t3igkjjBS8Vc4NSNHIv0wFBRt3/ERyKbPcrjzr9DIUgi53d3QsvY
sHjrUaZCK7WVfd2DDzXY8gXJImrCzcsaAMfY8AaODjWbS1uNq7ZUz0n/e5w44gcR4AJw1ne6jU1M
5eGGvJQ4C4CPPs83bZt/BpBMtc3jKuVZyzaxLI7BVF52sqQJZcqTsyoc2ag7cGr9M+sja1KBS8ct
7Atgzz/bgg8q7TkeRVlgyq8I0eCSCTTgkfUikY9vlXVeG0JKBBlQO7D9+BddmutjZIqwOTYjyDax
zWCtfThxkIqEYfYuEVjLuEPXMupB/4Hut9/jmkoBY9d+QnP7S14OY18/CPuVkbJPl0aZ986xTy6F
IHR11rX3LMsjSqa22kc3APKdgijH1Vg3orcRDdPBUnGxs3unIT4cXziQEGR/HIcZs2i/8lTQzdDw
XnigJAqshVU35LHidr7bc0nk/jeUVKjKXELWV48cKsCLeuTFiq6LwT8V/7j+DZOENInYvCL79+J8
UzW9VnGwwSPdT2Bi3DYTJgFgrFRvhNrsGtmKnR3nWUJz9Ysgq0zIfTYQALgJrk7PrR35sVkCk37w
9uNWBHKUPVX0XiRBgT0WpPcQjQ89nOe0RyawHPNXmorw3Hb2B/8IxOdl9pbZbIwW3Rn8exoY0fp6
PND2HNKPfmojiyP5i9MxDfiVU1KphNO56HB+QUSMY4LdfmChv8tI7qQQKMq3ImtTL0+4/bTpX++q
p0kgEAxSVDJQB2oe6ZoU5dqlOFkxFJ38G/4HRK1S2TnsF30JSwrFou2ro1qalo/pHj3iMqPMfnVj
LyOH2HTE1r98Dt8DsswpciW9vaezWp01uE1VTqoxdX6rzYmyfln5Pf0YRrE+W6sivb+0ZF3Ui2tQ
HmLJrVEZDvcOxGFtmdcQDnTE9hKN2ALHFXcFYn8mD7H37vyp+JE50i0o9G2M30sGVhirWvLExaMs
6gTpfHggiS5rztP9FvnTpGmp53Ob0+VaOC2tYXOJsihp4J2DFYKGGOJZm4Ii4kDDlWwvog9dgZL5
/ir7xrRQotskXrTp/b8iTf00UDk/Wdpfdvg0lk3koJCnt8iNLEDm+9eBUPMDD4vG0Fa03Gx5nihS
zAlxqWFTuA0UYadAdc6EAR9PqMKH1uuBvcHo1SLJ21FfyMcORSzTT31u4m4XM9QKld/PjQ+3BRbf
h+x3oFYPfGuR4NW42jn4+6IQA898jIX6p0eB+76ILvLwWunfacdnKOwu3eDci9FYJG8ymrceADgK
1FVjp1/qZlcB7SKgGAiRm901A5vW8p0eQut7572KL+QXCgJxnQioFkw1MzBX+izW1ztIBHcbwTHi
mjOYRLUSUGrg07CnmeR075dF62K3m8p5uPi++qYz7mrxaymc3+sVJW5yoN2d7IbUP2vFgeqgI0nb
irXnd+jFaPzPrDj9RqD3TX7hFCblixY4B/cjlpg296E/NVNULL0jXHl8B7InvH6Y55iQSDmBI4pC
iMCyJIqydtskyCaLSXUDUyBi3IImfjKWFVN3tSQge+vbB59V574kNTwlIlzeYQ++t9hFBm/d5d/7
UMyrBxVl2Zkuhr9SQkgSE5q/aw70BIrBYpoowc9VB7BL97f6iC/5MNF1BTgHRJstGokEYtq8G64m
ZT//oqmcg2/Osv8Ce8+3+m2CS9y6c8Uvg5rXrLyt7U3jaxuZjsvoQpAO1nPvWKJiLro6WQGSgGA2
Mlvt4OvisPqvKLzLyUgabrcfz/4AggPTKcr9qvq9B6s/kc4Cjd68PUN2F3SJWE8g7yjh55E8Mt3i
2EP2Zq0ANjiHwhT29xtMz6m8WuQE4qISK+Rf/yvFEQqCrzTj4kstxfoWAi+IOKyYGPA6KnIM56uj
NCcKYFRd5qd+Ap3cujGoAd9h59cds4TrWpeiE1kGeiFd0tZ4rT03bcAUmIOiX7pCTKrYNq432jmW
sjngXI4yyfTqxaqaJWC4inmVnsLz66YbCR6b85k7WjzOq5mp0W9NvKSMYD8h81UGFJS4YR2F76nD
+wZ8NhPdCpvzl0PQiQyORBKjFcw2mLd+I9dzmYiajNRzsGY/CD0NLxphrxTlfihG9hc+v61pnWE6
1Ni3YMx2eL70AOPzPKK6LRfmXaMI1skxiPGVuMuhA2ZgbtfRCMk2mE/e4hjjwEvWyp+NXfbwBtkK
wzYCwL2W7WTkpFIWzV+JLNZzUaosswKi5vInQSYxKxmkKlbtWEG3cozocKUdKE3nRBTnfSITDf8m
zZbFiLc4ZBRDRvoMSfxCqI/4QOCNWknvSe9c55zHoK4+89EBiMlAKqhgdV8FmsIshaIkE320lYaB
LhMK1s0y42QC7I57s4qmxK8IcmZVRs19bgCeQ+kKWUkRc9uuce6kMwoOHWEy5w5rmsbcKJy8jntM
xUlVZFfvRLwWx0LeTuTDgwsaxrSZ1I3te5N4rfVBjndWkmrBamG5V58qh3qU4zmQj/6jqq5vW4PX
T8ygTHb7vMNPYJx+N0nOOb84aV0uyGo8Pyg3SvEm3l5ETcdnr5EE1GW1Ag0JBwibh2f1SirVqMY+
TqbMiYapHs9GY3WxS78dmu3FsPgoiz5IM5JXjPx+Lad0A2QcBxKHszNufHn46qTVrj2r3Aau0z8/
pLctnFrHUiXg6F3whJNympvUqG8sUdLwAAIOlgnWGkMHdRvDP6kaQ6AaSzhzt+F5rXa74QQgtk4+
86JN8mKypJTOrRgwm8SgShzOTQ4AypgADX+74hcw6RsgaVASZL+scmGeh8yNgTOgmCLMZMaD7Jj+
sd2l3fHJbZIbsQlwqgS5mCnWm8qOdTbb83w7AJWCJr+2+ZtzR2C8quf++epay7fg3qi38n6UDgBZ
8nWcwhKmBHIz5uknV+rrY/5H1mKxjC6INXdYzJ6AxZCed3T+r0fH0w+teNpsvbuMs1Urba6eOZhh
p4lI2sLyvimAQbOUtpauJlJtYQd+N0A5tCuVGDf/5MI6kvjma7izzIjDyFV4G1EKO9VKXg8RlRfx
FGQF57bWDhzxwB0NFqJv5X6P5gbdgEfGmN0rAxx0lDLj2TYEw0VvnWpX3AseQwCJBOMulDGfNAhE
ByxQcO4cY1cRbuTxvttpZLnjkC3BNoa24++QpUOX2ZYqWc816OHP2rWhXuelOI4mO6nWBl+HWHDY
inr8EVYYfhUYwOUYcqwhIVEW/ZzmRg0Pe49Yz+8x+/lsbEZAAEeZrk4UasCBB7P/GMGQy+mbgNtI
4HkAw8gKPmDjO62f9J4JvpPO/YBjKxqOJNH9zc7Z2oEttwsMXSdwKa5dL90/UOrVd6ifLS56n4mp
xXf9GmMvixR+4WF3yk7zbk/0WsXKaIt/bNfs5NgZxT8C2LaCAWqDmxXM5h0zYwu7WbjFpB9bKyhd
KHc7OlACTn6wZsW+i120g0kzpWAaNrKIt/o4ywlgept8K/LCMWyizaj1Yzyu0MeBIiOfTx9y84dx
mB6q9DRmZt0GoEDY/hjIykkpX4HaYrMsyEdXEGNM8d7NzsVky63MBHts7lhD4eqJvHKf+T40nnNP
qRIfU0z7T3wqN9bsjFobd/Duqt5wZ9iBDSWMb0/XXP0A//rm1yvm89vu2TC+qqFPkePv3ezHbcjR
ziaawniOFBiEahEm+9x079TX78HGevXe8B53ns1isAh57dLwXCC31vtkkjplP8e1JjhXzpOt9C4V
E7+IcBbbFEm4E11tvXEIkidxA7oQgnuUTMAFNzA0+mzzdOdGfwsgAV0HDIc3EF59bOPNFiX5gd+j
kjJ9FA0rUnBI839X7S3WiYLPv4aaVfRPdNybC0N6erliDOkNpQ21gnYAIkVZuLRwEaCED28743mJ
ejw15dbDWyMfHzu80naWrjbdwRoVUO2GG4ZjjuK0UcjDKS9hmRxxNKriNwRgA9k2vYUJFU5bKoIv
AFVl6r8E+dpRhmde+2lyaogU4q9RwfVvEKoUxDkGzHal0xEJ1i6HuPvzFRIf+BVImBf8EwtPfJWa
UmAEA1PM7clNz86ih3jT6esumLjJ3gWNuVrfY7cB+YkuuXr7rGcoMmwyayCMPhpEB2fBb79jOgg6
dx/uuJSJDNTWW3JEGJ43W/eDSPhtCcXI7EylghNiwy9/Y2PLA2Js2ltdl+/W8NAB8ytqy8XQnIcS
LnY6CRrY/pw1cgIkoNhIgEDfue1mUOw/gmOUE2Fod026N4hYZ+m1ZsiuHbAXMe3ti7SPA7xFx0yu
g7EqzPamnN7ze+lmFi8Ottyq4CN1aIVRAf/4qivPgPwYYah9CxHd2cdh/GAB8EpjPIdSeJrz/5DO
8BkdQt/1dU7UxmO7pTV+t20dGsSqgoNgXUZBAiCLxCYUH74uSTQmISv9TwlHeJPjU+8WmmimmxRs
EfFaJZ2MqID/+Nfxyk1T5YBTlb5aIP3NzAWr7d/efFK5Av+pFM6JbkkQ0L2lN4GO14mevLSjcd4X
CxXyD6H8tvwEUB89qPEu/+9C9EKgqEr+8AI8pd0tPDyTQBP3Fh+2wrpZz4HcrnJ5gJRDCS/dgOWH
V9sbGuxyqI4JIMWGmpl3WfCUH7FSym+h/EstsM4O/Tif16mJNcAQfVsMsXe3WwlxtFPs8Z5hWqIp
3OHDUGB7deKyNKDTstBN/9Akv0z6j+lqULqE3LNGUwcaqo9FYy1Ng/2VF3Qje00kIbDopamaRm2o
5uYhAEvGX4bLA378TerCJdZtsEoQMCtHhXe796kyl9dMxumxbJDANd45TN8WkP2qCy9nKLnXVHK5
PHirakoBn0akrauZw4t0pNH+Kv8+j3qLZz0NfyJttFG+C/Azv3uzcrS6c0OURePK1+mAZ8E0lZ5V
/A8n/nkd2+8MkCH0chEjqp6HjA7gqXx34+gfKN2cH55CWyzrwbUTdBUZaurzNZAj9v5NNPOMrXoB
B4wiQBFeyHUyFHxhktwoiELyTdlgkh9SBCbLdiIk92LH1WyM83IxdXExwAZOWOc6CrsbhUX5JMA3
jAaYmss5JoQD4LIfXTwVIPujwh5vHeurJqcxBNTvBuJ61gVoG02BUZHLQTOUy80lAinJNQpwSv0e
PdPld/Vui/aM7V5i7ht6eurhT3bJE2oIvEiSw2eacWXEojkYtFQhPUPYEwySK1Lc75aktMvY1PmM
mkIXl5ajVJfhgAsU84EsywLyWaE+gJ9lYLNm1ZgAc3xLT2soAdT3SVnPh9Pb78qZvCnKmj676Uet
kBkE8TSi7Ri4p+TVkWfiYX2IuvxIga2rTXcsL4EoOyqUeMMBnmziKmQxLpUTDFMSkouZhrT3l06c
T44zlsvhCp/nusjHHfTfKxKJUpm8civii7UHHMrrTbaf+NFc29y1GkLbbBz2iBZ2XvwzTs8MJTkN
RvRm6numOly5Ww9EtV8JJ1JlF2nRa1szUhb3FIm/etAb3ZU6AgPM75inET1ZPjyUR9736o+BUj0a
8+VGQkqSN70sIP+M+lymcD+V/7KaQTKK/LqrZZsptVLJ7TsDUWQ2HHKKRCJgIL90KE0CKWA7g9MU
svL99iN6+/kQMHE+b/hPYONov8/MNJXcrYBuduWZTOAhBTKGvq5/9yoZGmCS4znCHi1/JI4b/v1b
ElPqmyGJQf9BtemCjn6+51jF2ZwRn8tixxBluq+aXM6DvfUTey2uiqAB3Keomsj+CjE55SCsxudE
5BObLbALP+n0dvav3/lWugm/7/qhUU12TJbdb0o748jeCNZQ5blIcuuF32lnmtvQwRDmfEvvEP6P
tCDfK7LTMw9DqAsn0a9PQpF9Jf9qIBW00lJRD4G9XocyE/YktBpCO7v+JZSo6fzWltI5JZ5VK84b
slTLBsieqEmRhk49lKBv2hR4ok0OJp2ugRY6UQftoMDFPidwB7lVKJCrozJxCZrmmiea9GklDEj5
ZlfceWVtK6R6lDnZ+mXcm7+ys/DJGVl3bIBuRkCj51GnoNGrBEjeMSZ7dz7nOS9beYll68mgt6/e
cZHKVCWjJ0xrsdJ/7Km8BiEgX9oaBtxdSlV+7pXQ+OiRH4Lm1TeNGX+nTLIAn3Pl+LfqI7rHutyg
tWyF+tkmSRfEhBAFAqoKr0k6Nn9X7ZY83SkIPTR1kNt4sRQ1YFW08NFjtoSBSmf1u6VB9mi5808R
ESRysuHcWY2Z0Xx65U5UE7fXRpMuehuEwkvIrbsUo7K1ZE+QiHu3eTTvld+CLqhcCRSf2zFmZ32B
DNTl2OmioHZgGHE+U/ECwqzN7vVKqJ67aSi7Z9FhJtBTTxiv3mAhWso16UafBwe96P4o6JOPSmAl
ILk53DGkb+W+XPEz8pw2mihavVv1yunrKqL4/IecVIQ4MCFGAujnPzZ53HlGdkLX5QHpQ/N/3JA8
N7NqLoSZkq6Wmkb2fOSlNSJsD6rB9+vYauekWFQGKKZmwWHKPR/MY1VORrY5oIbjvszvvrbuiCTK
fwEOSMRV2RCOnvgz8Wx7tuXlHKgdRHVmgyGBVTcGdEfsvq2DN5m7rRn4O0Osn6W8xNm1QYpf+z1u
QpZrQubvgLFMPEUMMR0AVBpMNmv666BvPpwdAUpQH8P9DoRQrgLVLpBhQpOZev9BWmycjU1qSYIj
hxiJTT8/3Ujikhq681BJaEj+3OhTHp9cVncx4yf+9m2T7cE0B2318UICW+FfKXHUG91MDFORT3dY
5bPkQslDwvOgVdGG6zvapdS8g0HotSnK1vQxUZ7SeAmATNuThjKA8HYFH5uUL4RnAT9uqpuFVt21
vxBobkkwLLrC0QYG97NH+tOH6rRsHR5FMc4+8PZ2XFL9jnNMN3vpxSTjoalE8b9w0ZbWTxn516OZ
cyPQHTRmRnY+5JnUpLTXyFmxSG20Nc0p0Ea/LY759DNLvLzzpl2lyjxQga8y44XnR9jWuOpVA08l
mx9fYZlXSESiDJSrm/MxoyyR4kGO8ecx4iVtJ4udQJVBRwG3ux3KSkrP4vamj/HJF3HwH2WNFvEj
u3dYGsgyzPFtYVbOJH/gUco6VaJOxdWJSmlfj5vmlNXKbt4XmaC6ULsQo4xVQ+WzBbBsH4c54DLH
4ifVMx6iEMxYKvageMhfjZfn/fVLVp8cV7KEg6ZCsDyYWmdVjJVWf1B1t4WymvRJfjiWqZOvFanh
pjq6kwPjcUgIYIl31wQ25XC7aO2hiPfqohNoXQBtMc0Ho7cXTfcz92vMmEbwxpI/rIhzt9/YwgBZ
Gumu3UfBEbnJvIIfejmyXaCAIIajAAUNSanh0dulitmomyTOLp9+Ce/LWiBegp6Z1eYTZmTP8pOg
vPNpEI2DmDeX1VAiV1JPsJJ1PACSpLxi6i6bO3PzI6HAaqZZgp8j/QYA8rYv8+pQ+r8jNDD8CEiy
Cxcbkn/1Hj0MZi2Ty1wbxs1YTdRaZ3Q9qUyng2+bq9NVf723xMJPrNztOuBW1V74tjFKuIAo6jgp
hu4bg/vq9ZtD7Qm5rtdrf1FvuYOqo+tzZ74tWlMQl3/ADaRRKNDOn9P2AfciGOiFu0uDoUL/I40n
/KrkKwrevj7XhB7MB0NAP0D7DoqZGMJJpzQjro+5RyjzMqTPtghcRxgfDIIlI8on/ZoS7cI40l25
lhgNJXcgNf6bCXOoBWPoG1cl6qh+yTDAC2ab1HORHxSZYEPxGV/B/fl/HXWqXd0Y7oNcgYfVU303
H2ukpVsUcdyFSNKmaK0E2x7lCCFkp8S172p4I8dUPQVn8fPAkHebZ+/HJU6ytffBy81PmhfrLFAr
UIIuwUg3269QkjmTyxztb91MufP7/s7TuOZ1u5Jm4k5s05Bb+U3+5p9cM9kW+O5oK2S1v7tTj5rA
PsvquLScsZ9v5Zq3+0YX7B1KsRJnBz5pWMt4AluDULafeJYsnR6Mnms8XuMDYwNnH4t7hGBpsiwR
TTmUGwTTgZt/ga6cmH0upF+EretIingdWqRH7s/JcJBWdTise1U5FCqlGTjhZIWtBoUdQ543/X2M
xC4vlvFClsg4eBM51DKWyHrwygye71LaoUaNBGsBhEQrHfT3Y7fqqUt52EcY5Y8qnuUrFPh1crAy
jbqn7/TA3vQHPsRk4rhGjwfh5AF4yLZRrEIITFIA5L/nN+8oOfv2q8H4CJsgIbAydNqhVfNLOvI9
GaH32PZOs1l3GdFcf+xzxVXpCI48lBSMCnsFwP92OlRagxku+/3eUwkqoIh5TI9KujxuRtU25GC5
s/NzuAAMcimtuUoB3ihs08HNOhoX7Xrb6XLlorsq/WroUr/LQU0mgIyOddwgywJz2Ks2gnXPKh9E
G6h+yitsQOgG7lrAQ+uuuM4q/rJ55YrUiijFk1k/UpwXMaJsrUmsAeEC60DDUnYaETUI+nmhhhBW
62JWisVxD4hVMCbF0JcfEYagi3xHWOUI3UadMy1FYowwrYcsekqw7x9Pdf1VYHFSglFQa9a3/TE7
DcW7vj+y3czL7fYU5Rl7Q3yGdwwDLMbF/TvFv4JRs4tZiZAj/r6qKjGbsAJDzGdNqbSoLSfURopK
JaIqHda6yN9Ha4jFg8e5iefOui6pCpnicc5SsF+uOeusByrHG3duiyT15ABElETyvvHEBVFmcRFD
2LDlNYV7L3UCoFhtu5cdszvHP1Ipmb+jTiCys4/JrOWmenlAI2TlQcOCi9TFRpVCMgzsUq/P/TqC
80nicj3HbPLg0wgtWV7256FVGKmw3dAyZCGT6VPm/rtbHeg8LHTehPNwKPo9atks2nvK3Duf1rrG
2jBPpb7ICnFLgL1bynGQNBusDIjFD5xRe855+VA1MvJkBAtkMhuqZmU5yCgYt5DAs+YIlVtdX5w+
2YvFSkxEv9TyhnYqH4/dAJGwpRrA+pyGmFq25BFOtJzOcvPMEvdqaVZi6yUDzKFLRoCHfYIhe+fS
gtVDOHpKqEAy43wNHxgx4kBkgdezC7+vWr7R2MW5NF9Byr9+aGHit3S56TVEMbSZI7fFRYlrDnzO
Wb0YGN42sI1CBFBb9Qn56CoAWd3qUlPusl6yGONFkTSBlH9CNFpWpQXrHf3lDau4GZquJvfoqcyk
TDsjsbFlJEgxgDkrmBVz0uWD8BxtHEv+Ia8g8PSB6FCx+Fy+xAig156zZhRmKlvKry1YjO5U/WRX
TGA0vd6ckhOcFKy1WexoARhkKIplhyq4JwBkfTlt2UJlqukxql8O6t1VhuzvYAdRFSbzmPR5c6ST
Rkbcr1CWx3irXnaQfQzZbceNx9tUjE2cvOSpnCxOYzpIZDPLxcaB3RrbFpwev09bdKFcNigW13F1
eZhsNoKw57V8zdO9o+l7M5avv3eYkG4P3sRFmP20ui3Gtm7JfzO3lr3wqbhy8y6i4GjHzfPfMerx
Cx4zMPCxUBrcfwAgnvMYre2sjr9K8ZrmdRsf/Ymw304I+o4SiYe6KrXzoWpmnu/r3ohFVeT0FPzl
SFbbvL3ySXGtmr0VWY8ygOOW86d84nSO/LP7F5yd/AiGzpaYx0NQ/zgNxHDKEjUDMNI1qPCxzDlU
92pSWv8aDKOBWCGk/DQ7GCn7qIIaUHMR6SIEp54g/FJLYEZFnl14q+GEgutPOH1klF5ZLxk5+KFF
Q3HxQpxTUNbZJS3NPAxh0brdQkp76/Ug0gMexN6cGZ72+9Z8obd8rVQxSSIlipzvKyQ8nBK1w1+I
SFIC7nbG7t4ZfQC7NCG+lgyVttAU1dkFV4wog36f1djemHpKWzDTUDEwCK+IfcuuEEHqA6Y0ENQt
DzoqfZcNgDIVGuZ+3NdJJm0Ykp80CrOJoriALuEDA8W2pkL9xTt1Rv4M0dqHZT9u3YaayDAOce81
6sDz0lNgMKS29hm6fXcUSfwrDh8aLv0Q0nbwpLajrOR/jnvLgaQe2ZdeQNYUb0cc4dowSkZd3bKT
kwnbkHtUdH2Gu//DxCQQBpFsa79FAgViaq0lsAuznBpvYvkpRF5daZLV5ZfyCPwYyf/Lc3BzbyOr
/qYHojX14jjdXrCAUR3jYx889wJjr5ZFbcNR5yx1agpA/z72Lst2r2dnGU7J0BxzsZDIk8vT4vIQ
rKfFur3DM9VeI7doIYqWlqcxocNA7iasU9aoJ0XsaSOhvQ0Ax2ZJA9H2D4VR8GZYP0KalTLe5VjE
ymaFGi3gG0SgayT/Xsr2jz0IN0+x57bUlk17wY040KRkNSaLpyRE2LmBZ26DWqKpt2JSvl/g20hw
KTgbH3ImCCY6dv5WNaFTN1cKMOBkzErf05XeL7VR0Rnmpfy2OCbBcB4oozwx1qN7aumuCfAjIpBG
qE6+7MIkkA1AJWfp8sKlCiRQqXwIVR6atrigagqaxDDFj7G+lIsF9DoFn44sdHSuB7NxqTkz4WtD
07aAN7EF5QNVcAbMZvhHZokqwwis1yLRHqxFi0Zx4rjgI0tKE2yoizpoPASGPfPaYL6xI6FQqI7H
yiD/sLqbzaxrD0zEFeYVAqmtL3BI4WyFsIJhKSIXcBab/Idv23ISGbWdzb+8/nDWGhntAb2lT5vj
jOMfxn36rIz8grUOmoCRc16S9n3T3fOHdSs9qoBPP8raR0NrKSMHVy3fuBACqQMz6YQ/jACHHoFr
qErHy8jStTEjJm/I6bSW3IjJY+m8Fbw3UU/Zg0m9283gNQGmFJ2z0CQ2b+t/MYgB2A5WmwlUA13F
YsMMhMmrJitbvLPLvPyci7Hg0sevkS9ICm3/5gq1/DGMohIc5B6C7Ut+qyMtwkNXhdRt/CI/398F
LilvGtAEe6ovi/STf5Vn/246TyZuSJZ5wbzXypYD4cvHuAEBevMUbA7eCHqZGx2q4I+UqOUjIKin
XvMcp6MU19ALfeDekee/p2kwzoN49DOOLr039Tz5yG9HN1/nG+M+mTnOyhZW7fQdQtzWBUnNF/yN
YttFEjArtEyEabicZaya7nNkfkAT5aAC5sxDWfTaDp/8zMCl3qKMIRnpslPRgVmjYJTbJA7a+f12
+eq/0T57MWZuTwPceQ0hpd9BEcaJFpr3ENOI8tee4TEBNRpWvddwhjaULZQSp2E3sTpWaN7HiJwr
UENzh5h0/bqisK3TCfpYf8mk/c6MoW9XG+Q7bWkf+CZaFbDCMcvRSXCpmquuSj/zW6didF11a5pu
pId7p0GcgDCABFMV0+qMUw3+QXd8egWYXYE0c+IaTCPBKppVBPpenutKPbG8n/RzZf8Ev4OkISSb
QyV8dl4zGtVKQwadwNckX90WkpG0botBuPuxlB9PQIfJfQ/20dL5e8IqabEeKLn4Y9LEAYP9S5iT
n9v/udQ6oCPjCaFGX+CCXL6ISA9vnT5gDwBkwc4o3B0/+fi8Ggn/rt6E3KnYGhRUrnYOv2Hy9txt
30q0U8tWWuBgA6KeE7FPe9VhMuRxi8F1lb+tlovAvbzYfezl6WProgWmeuo4fmFsj9V3WnIPsfQ+
WYWyJXUtP6VFMhFEtHkSY1K+D29BLD6N9SccCngT4jdTzqFdnXRrLSIwHnCVPRSTEe0fJEGQzT1U
VCtqSAeSBrGngJNMKm2lyWwpssZDjjkddMqftql+r3n/Dq74E6oAvdS3ttncMVnwHLafPfLp1p8F
K5aIIUc7zPr0TypSmzG48m3vCCoXsVaN1rzCNg2iUqrdAf81PTyU2mR2lBsAZ0nVEP3zCCkmh97d
XCp0RkgN1w4E/4W2RD+xmR8+6B8vltyheLxTvKwFny1kka8EMxKzvg6yHvyohuz/Z8tvQyC5pt3w
sn2BbOTkRCmA7C3ox5g+WsUJcqg/MQB8+kUbP219kyuFcvFN9McNA3+yQ/3+bLXXLuB4CNtmqwn9
LwRYmMOE+TzWxLzLJ6YwrLxWHDY8AgXMcC1giilFCwURy+P+xMmBZGaHNOUn0VOuJcBQTepuFdlM
o7gCxa8m1oEfi+CP6pcCXtKTQ2JpEw6aPfBAXQwerbC1Cxi7aoYgestElbMV4DIoCVx25yzrvr4c
H6ZOD1/dzRyUgoGHOJwIPuhZSI4gihzgPujdIWXGfd2iXIisSKi0hNDH+2OkeH7+6aW4LH5/pll/
8hhNdfusrElH25dDCRKIfyLc/3PLELVemfO8g0rGecx1ENjlFvoKMX4jC4kL0iF3CcEt8HP67bTN
2alpgqAtkadYFyUlb8oERRqnwXvFTBd98w1rlveD1fLXWZsRmkLbnpx9dMaXcPhuDoYo/nsoByjw
ZVM2rFREzYymPNdcxhj47YIjvK+8E6PBPKD9GVZ2JWVMpTZr9TfxaSkq6Dzyvnn8V69C5xVE6ssQ
NEzkEBtMTgV1IbK/Uu+6kDfxge2/2rzGHUYmnskTaildyubD058puVlsCC+MSzeap/4r+bZuc77N
5Tsw5RoUlP3t5JDbQWoWS+YwxEiP8XRIgK4ftBDZmisqt/NkdgDpIhrIwGFlNFEdyomWmgbj+YlW
9NhnbqHD/G+D4u+Y2LpVrUSAFOoH2r3vRO1NDrEwrz/VXlbqA5eBiRBVsgINmljTDPlnTCgt1VJD
tHA6/DyEhmlASdx6cjWkhZJyZb/btwmmQdlsw4fMimSJKF2j4oZJ3b3DgAIKK39r/7/Vx4RPHjJx
RLId3zql4nieVOsj494IWL63jS2tDhvOOi+xyIDCAs+O63YoN6z5ljSwV4bLf/t6CFpqf3VanLYJ
JPX2sslrfcONtBU6w2OtHvuyskJbTW9ep7y23frSk7Bb69aEIudFEc32M488EaEbmb9UKWpIvz4s
L14ZGPGFtnsyk9HeCM2A7E5K3asB9bd6SyAzljkWOSbQmPWztIUWQGBM+8CRlDAdN96K07fJqZHP
VwiVlURGSIURZGS7DfegDDgCFCHh6v3rX37fH10IiUYe09JZCgc/gVKoiYdUIg+pxuHFOoNM7608
qiwyTCKhZMHm8+JzPa0yxh2G5X5vSlp+MctR/GWbSUbsbkrvDnAfqg8Ph8+jGBlO2jHfCXB6GmBg
ymfrKM2yHGbsphCOXg78R9jYPiauWCvbQdBYs9u1K1rznozko1ZHQwsW8ALJOpzWLLCo9iJy6Kq9
TmhPggcB8w8fopYVgg5B5B5JmoWi4gSW9UldCJXHC5XvgspSPs9tRxv5sI+eKQXjEGtc7Kp9oIGv
PQTxy4D+N+OvyfcYPCszX3A8wt940bFeDpcenRoYMET+6HtvG8v5JfkKda68FtydeQrC+5CLmVFK
q64FG3GXfdNaL1JrUuqmcwLf1GzTGlXb15Fwv83TRDKE4Jol9Jap24mUtpDFzvVaeZCjdBOUf1Zm
dDcla8UCTTrGHSOfvtqBukO9gxHGfR2CSUJbpzmkwuLTZs+Bs0VGOSyEWWzsuqKVJsK9ozW/RNoT
EEQvwmIogmjZ6l/VnSNgXX7nochZ2FE2etK+ZzsQRNYZNgcsZVz/YBqiFDqRl5LhFrZfN7e0Wjaa
E9d+mdh11KxNh7k2fSU44HBWNojanpnRvGjbgh21O2IFj2EL0hnBOdv3ssp0/f+UWQFg0n51ZyjT
EN+rcuyi+87XhemQHEmlvtvdq2Sk5VXbytH+XPQBFnpeGhgirk9D5pAl4ua/Q1K+G8vV4JGOPgax
flar78lze4TrtSGaUj3DId7hbKtMwbsdlWFenwpYwbCWnqvS3cpVZ8vicyNsVEK31bPVrwFKuUNC
dEkbaWobbpCbBnEck2dQBLpWtS6WLY6rdub6qKfaBM16wBw6Sms5aBM2TU1NIpGYkAw3yAzEwIid
/GOnMkHccUm9aoRJb+xZhK6/A4x2Q+K0O8wLnhBoPHw3qrAC5FzuHLS6rPJkJ3U+5BgQ14JGHEUh
33IbbJvm5Fb7QI5whxI3s26AYBi+CwvVEleT1fFVfcOreY43ZDFQM1817S8CsuMdaugo/Ie4w86W
mNwVW09r6OF0U0v1Cvo6+bxjXJ9woVtidYWNMB2WN7J8NTm9+7l8tRuVuGkeKb3FotoATdw/d2uw
LZTM2B9tiwp7r3qSMErJP1kzXDi3Sf1jMn4uMjtjxdPJXpT+n6OFnU33ypqp1wyF4em5dCec7LQr
X35m4UpqWUeFQw0OnpPqULL67OOuL+IMq+6fE3thjt+bIpj/Wt8Vpqsiz4s1LelP8SrgPGT2pfa4
ZeTL3SESlh8knpWXgywfiK06PemMGEqb6UDE8dHocvXSxOuNjHgTBYSUoak6HBPUf82tpEo6kc93
/xwhIudkShXfHuF6wZyrrumcpolWb0UuRyMOAvuYFopRr8VX0zgM/Y+cr3cY63syvwzxmk3UPvcR
U9IZRR8RWq8RhMTuNfbWD+b04Qq9CYTFZjW+jQXKDIq5IVA4hEGeW6RAfNqJi7C7fPJBVhLQ08Ac
r7obQrsHOXCwxUVVw7PzA5Y5AV6tCKPUSh/HIpNXLxUr6QuspgYTN+hbhTe/rsxUgn+CmbdFDhzY
ubN3Xbcm/XBwF0AWTyIclWhMtwyweYLPlTV/U4oF4e3jqh8XSucHWGOve7USDvnTIHgsYRHnNdNH
hfZ8ymowxFjNn2K/cN6K7wykQF+/LWwfZg5gWRPxY5iZKoB40W0jI9Rr0dd0dPvYEm0zElyxEfGb
U2DGxZ6q3zMrgIQr+CHkcnB61AAtJesTxCWUVDTxapFU0nzftcRcvep5Bx/XBPDwr9QwCKA3Ygkj
RzVxYp294x+Cld3ch46uIsfos6ewBQ4EE9Xu07lyzwLS1GiKpTVa19C/L0lZj7nIxZJ8AzmzmcWH
D+FXDCGNdwtEjoJMoIuwlzSCURaMsCl2aSFG5MzuOD3y8uKLp+9N9OfpiwkYw4IC+2OVEcO1LvME
5YftkJdGYF7madRuyIMuWR2HDwVoRFirbSInBf29nO+pgKDLhFQv8oebjeiGm4lIHFIltXyeDFln
qfk7nqHMDAvObjYeq7LYuJSghO8LTHsEz34oMSMBleIh4l4XBtdfUd8otwDgNLxH1NgBpAdVol4i
yRa4u9OSyRVk88n5UTfITAWcnP2bidabLuMJ3kctuctxv3LRk3ZaEn1gx9FQzB0+Gy9nd1lSWHyj
3+tXa3aAgSDGD0J9md0284ce/CkzdyN7cHlLy7QtdCNPxKdtmoFA08aMFwuEZbm3XeCp13cqlTWx
QzUoP2B7RGEkFrDGvued/d8MVYtTZGEmdCgydx24t6vcbVBR608bYhqZROB2A8mG7t0Ala1LTHV3
dCVJ/4BxBAvG39N7sZseSwNptAyyCk/SClTrVgvyl8Hz5+MtJErfRygPrR+PA00f4O+FvMnw7o3h
jgLQDok6uS2Ea4l6sUA2UskMDhbVv/jqzaNrg2MIkj1XIC3dadOTe+7kjU6JZ9npazYbrr/R0B2n
q9+jCK8l/AixQYEPGz7rPLNhq3Z/+WRhLhFE2KGL+Rm+H3/SuloTqBJhviPas3iKwnBMAevIu8Dn
9UggcbpwN9w2VDwz7+AJxx5/MXIpzrjQBTKybqX+vWGR36kYkZov31o21BO711dTN7phqqOTVImH
L2y5oHXQFRh3nFJYDnfxSon2GGKooIUOr3cl/vx/Paj8G0FnDA2NrZ0lo5H0MD+tbA/0yNhATj4E
pQw1LFM6WgYiNmQhtWhr6k+LMt4jqETsgXcM0jhdnLWiY29p1G2sq7LBknGKVBxYnVO4Y12uAlJt
WRJucBYs/RDhaEtaKvbDYNWKOUjdjiotUOeSzDsMMg42s1vvJJJLgvoFtVDruTHB728A1iZ1ZwSG
X/zJdZnc6FA1+Jt/fH0XY3FpjfQOZIYgv85IySezUCbn/6XaDwGYYM+XNtMPbSwkQ3fsiDHFm5F1
c/1ao9Rw0vho6T1Wg52F68NyRQnO1i8AZSSRc4JrgC4yg3XsA9tXPh5CErVYQYsXlNoMJphCT90D
qHBWMVb6m5bLmsBecD8JaA+Nmlr0gf8uoBDlJtuJhduqBR2W/iviujw55iNxxVdxQtuZHuj/OnS7
khVhFTwGbbKrYPa5GtLXB2+kupFJT7GHtf7pzAR2EE7Lv+fikBbtCxcV66uf4VmQ19pS+7wTVBJz
xXOF5HKLbfH94c3ZeQ6faNsj7tLkRw20KPFX5ERiNjqklgjIa3x7KHP+aJoLUWjbi2aM+L1170YD
deHBOp9NrjVF5gUBKwb52sYmqahW4jR0eV9P/R1OL98eJaxc5OjG5Kmq/RUAm4xpjgCXbAgagKAd
4Hh6ePvoIbApunC1tAUloxvt+68E9g8SJlE16mUalmn6kS5Oc911cI8lBSlBmDZAhz8EmAc2LM+C
2eDSDC1CwnGT/Bb43AbGlmOCUldf27cRuBvrPL/pn0GmdyGdvbGcsdbkI4aszxnPRfcCGQRqfh8Z
meovTL0uEAmrXn78RJnwWG5X9UDjqUTP1KuKryly1myKR51qgGr6zXOTmv+8AanMZdCM/YnSE9t1
Sces++awBefhJo4emVB3vegYmXXtJDlP8MYmaZMZMe59Cx6uDmY8oFO0KYiy+kj6OqL6vLfQQ8Sp
gYwoAR406mnpm8BVe8Y+HwuNaoCnrK0BtkB9HsMoPdJR6WpbDT4yUm6mHlnZD/xcxfuXahBiyGRb
YhnfODeLWMLwLdqqZPQWRj6t/7s2BZT+YQbBmHpwruSUwdltFGMeNyDqmE2xiK5Ij5hoJ59oXzle
cRLxrO9pv4ycDnIjJrlL4QpmEUQo+hN5xP3PxVH1qbwFhFR8OGLelfzVsTAEDVOnIfYZHVFg4wlH
bjB79j0EXKaLIDtuwUnKkY4atmEjux4mwzdRutyYogicmduoO0vy6mIoWIx0l4Ukidd6gOWlU9dg
pDUW0cWmLUirr8uVkSUaSZjUA0zTqTBRSBwknMm/IqqRaRxHvBL7GK2MYHI09onFLolM/h/FPfaM
gjnfXePBog0+C3PWjkJ1Kv814oSsK3cOZS3er7keiH308wVyTllHfU5EkARSR3vaRbpIM3/vaw57
UEZsL6LBEsK1VObaH8EEpk4eM76NC9bE5jYiAni25F23mvjAmSmbjHEu+ngZhXcysbiNLCvOHDKh
D0QM8jiZq9eJSxDIpB3mE3SHnP6EcXCLwZlOsms9y4TX8Rs316KFvBtTz69Df2031q4r24elS5ql
0bHyITSuRTfXh1f3eXTvzRdJ9Mdy5lJWwUbwLC3/Y2hDTJiSzS01hsmc54jj2PJ80lP33fNeu5Zw
cSA3FyMtiKMxdRAFJNZ4lKgAjKLUPkYzjwmLd7pxNdwOGWSN8eXur0tmsEWHAYPit1kuB1bZY0/s
+z0gG2alhr/l58tSYBBSX1Wpkd9w81RSVycleNw+rhBgSZDxHGnBh5iOal6gdg1ed6EtoX9r12oF
VVPICZ6TyMqcuJJN83hB34jJefiHef/5vFQ7tNe32HOKZEYSSaJNhnpIgvLfr9NFtcW41gEd9b3o
mc4VOsuJMZhAoLMwlNK3X4EGlpOs0CCucKV0eNcUeN1CAeUH0/3rw/rk8aAFOzgdMT6y957RSefZ
sArKS1e5qN0WOG6MVoU3i4TEaBST26uHKMaSuFzagVupwhqeZhhoxSj6+WKW9o4Z4Pv8QN01FQ5e
v7HQQHIrAmgbyUDAgpHuGrijE9HXVEpWN1uoVyKxnX7I2oPU9CKW+nMi0gYACCHjRYSzzEYj96SN
NFWJIxOe9+HudrYH5DugNqTV4OQr4F7/MX4Az0K1cZoJGLzam2xz8imE5aNBuYsVl/QyFAK7uKTu
Vh09zZ5QzDVEVmlhMpcTa8NblZRA6CSYqV3hG0tq/1BSCG0wxnLqV/qRpAqyBFVZCymv5JicAaRL
VJfh9FxXfwlB7j5eqPipBDtpaXqp5sXmQwQEZi/kJl08d70vON5F005YOjzi8bEPqenxj9PGPbMf
gjrd1QANjcSi8s19JpMT9YX+b/FLcl99HhOWSrUaD1qdsCEHYOv2rMIUVQkbYOOTlt+ygFA+0vlu
+CppmUklVzwbiVWbkeDyE5MJJTZ4dixQWT8I5kUwT6mpuRiEVxTElvlLZO8ts9CSit9nhgXRN5Vm
DoBRUGAV1EEXfi7SRkH33etb6x9440bBp35RFKUCMjFQzvRm2faofPUXmVULunj9iNwj1ERUBqAL
vjNB2t5uQWoWKyNy0i31XLjVFyt7IakjKiEPs161F/DxOttcTBiFw3m9mn/oPy64hgglREC8GEBB
J7Ug/vvBdM4M8UOKHqa7YyRca3OadFFNiRD7VPeObaXjmRjL22rh7QKHIolfbn+zRea5Vf8M4TY/
UVf6IU6TSxnbgqb3VUp+/thlEnUQJ5MMTaiBaBkWrSDItgTxuDhN/Ry9K8jMDFuvOq5S5j8PyasF
fPw1/kN44qr3IZRMejChO7k8bguMe5fDzLdEuCCVwqemmwxnrcL4Hj4p5XdVJTR0weBM0AwzTw6I
ApLZdp1R/dWr/8Gtg2e7giniJJ91j+9MJ+jdv3FudCZu92sfYjp1UZKHIjJcyL/7Eq8+9MoTZtHB
QhxOoMC5LSchA9uv8b2jVpNl8b5IIqOKr7I3j8HVGzjAXaq3geUSsaK/9942clsgaOOx/7XoEAll
rmuyBYkZgKCsHk0uj1sH2UHQ0Ow6R3KlGngrYzJUxyACNiHPL1snxmQctsqY8JQN6CAIzFshsPWY
/Am7kRFSnTfzuOXUEUsazvHX79CsEiePLPtWYVYz+5f5Qdc5Sk7+4X3QXY/mCbjlCtmT3fJfCoWC
poe1N7jriNUEykU/PV3ALvxHBlYFhwPRd3ZHM2e3QUKixwg9dIMqGr0yoESQq97GecszWvOxky4U
GzNzz7dk/Et/BwCcV5x6jzWVnYMrH3Mosq0Fe1yUDbn175M0RT2om5/FY0FXE8WKkDNuZHa83Hm5
W0kDZDw1WugcCoZVhrnePrdf36C3IulUBe5rWDxcnjbdSirCQ2APjbBrS+iZvOVxz+kHpqe9CcMQ
DnszghpHlH11sfkEL11/xfnCK0x/cvjWO3nHWlWqXSqge+8fcEzZlVNBUyBEv+tJpEpzGa2MiOyO
4tgpbCALcLPKOSYw9+Lg1o3FrtVdPG1vdwWQhNGkSZYIrc6vDU/jf5tctOBp4CsDLGIc2IxnQOiS
K/Z5Vdvlg5CJcG4z4xo/CT8HL3Z5FtupIHOopVjnrdovbq+POImb+17yjCAsdgQov4EeB/JRgu+l
Cb9fEFaWg5sSeATA1MIrgr3QpwJJtcMi6mn0/TjQ8UXFHis6nflX0U39aNOd7sy9E6dIE0/9bsT2
tPUMubMgqyhk2/WWePtv6OAABxnWefnZGvlPtNVZxPdpxPvI5TkzFl0ZlqoMo6bvntNW2EdkvOcc
PqMDzDkQKql8IicX1ip4Y+UpA/6ToRKzEjA6IU2CadusBS74jWZjNbqlmW5UR9ZGGKzvcJi8yXA7
DfVrpUWA9U/p2mnl8V/g95WQRY40PiF1HXO+t7HXckVIlexxP6zpbfrcl+RxDQHeWw80eEKdpU0L
+DqFbabDuCMMkTVFkFey133mKdxB9XxPoP9gJlRxM3gHs8itfIzudCX3W5t8INf8GrSYjhJmu4BS
urTvLGIq1JaO5EO9sKHWlKkZdhUUUQ5qlBl0qMX8Z87GRmGcktSlTqcgPXF3r8lsYxtsFmeE+uRK
uQ58A2pzzvlcrn0X4eMAntcoWy6oSMjofqlPmC9c+X1156Rb8gWOcKBPn5rZQ95vXhXnwydOEA0Z
Ei2So9vmLy78HMwcTEgPQVtVkvKaqHdjGkIsbuM5OmNmJhXxtMXCvueGk++wF4SAsBnPUGp5FEVn
WHz1ko28HDAgWhy7PxNuX75qB5K9s15U6SEtAr1EHkEzUg+4EF3t8uRIswt1NdUJU6tVNsa5E2uH
2oVtyOKyN7X4iF4czTUjz9nItQaYLivRs5gpHh4NZ9yKMPXuXUoEEcp9/r0PqRdb7EQCeARhPggw
xWz4nMjhV9r606OnXxipqHjERtkjm1fdlk8ebctk94O0ljCiP5cLerGISgyssI1qLtLNV9yka9KM
lPxo5LHt0tTu+N+Zx9Crp2SVsaWfghnCI/ULNJMjjogEP44bbQHhOiuSycG0oKxxksmIuaTMU44K
ZmK1noi8l8kV7Jyn0qnk+pD8K1lVsShYSt1AMnlT1m8spTzspbpLDrXqrowp182/trVG3kOxMvGv
CP20MAAYYchSTVlxdwwekknHbzIk9Fvev0PXhN+OQOvIjsTb9PFegwhytbMDGhGbrp0SlSbxdu11
b+7v51E496MRiL7ZzZmvcnMqPxvIVQBt3mpIIX1FPHdSTAJVpMUtyJ4h3LP1I0BbotwkXZlUcQnB
9mVvD19b2YXxI+dSxvdl65H2NRSBv+MpGt1qXjgu2KXQGUpqDFTYjCZPtXwC+/nda+GN+JwdxXVH
xzox6YDt4Qe9DjHjyaRkfrCC9dVzY83KpImeCTQSz7pxZsHLDJlqkOndDns4Oeg2VM2papUlkKfw
akJtf99aUkan/pALKTw0NiPnu54yYdTJR68Lu2HOzSXiUXLpgLPii+/vumwwb9RAfcP8pVOokc6y
rMKrvuLJG7deYqCedMhAVkG6GtwtImzmuV8tDzbqTGvc//PA95jn/WGqJ1JPFodcxMRSC+sWMNPK
qZj8PGgygmEzBwPNDtk4+DaIakFJbHMjqo6NGR0CYkFyHY7LwB9RaEzh2jIMgt6+VBidM2mjDo3N
TFfut1U0tVAcPLT/hw8dcAth8+xMUfYOgnzWLWZGBa2LEkpDsWhA1lOSUmhCBhTvoHbGwnogaWvX
yGcwFRaWyPFTovylLA4n8+AUe3zeGF1rH1EA7w6kmmw8dO0EPe3zFA38RzfX6yt/yIrfHIY8hMxc
UksriwwdLihYl2KKPkfLOr93/xnTTHpy+BxuPDN8AQQvXzYbdDRilkrILsHTRD8qmsrqfixQVg5A
MKqOZ6o0GKIzgJlhnwDNw6TMpCck45rBOaKIWj+DEJdDJrLBe/Y95snp9gJMjGXnujWMFl1FhDVk
gUz2Rbu+e0G/6xdIiwNZeosTgjvHxuxzfE+Bzep76UHlKB36VkKsneyCX6hG1oqfUKChnam9o7Rm
RcHYv5B7kwiklU/sLEj6NFY40lsbjgHbNVcHvr07UJ6i1G/dt8ywkbFQkTYjnNGg1I7VVlbGuHiJ
pBYk3BIabHwY5Co423VzJUUas+Hr/X10qFNwom0djO8+fv76VOJNQ/El9e+bAnHKFSyB8k5WfF83
fyY9UuwK1Ga78KXV8UMG+NCMeZMyg9RnNETYf59vGa1QPBvs6ovM4o+eQ96b+ssgNFaiV5x26m4T
9jSFiBFd3vf2GxIsfeDDUUsEsrdLFJ1vGoo1+YOdzyQgqy4v7H0vaqa2svBc+vPnOVerSsXs5MvZ
BDgLgXmuZvvjb/ISQDCVLZb9WZHhWRuTl38GQ+lbqHWUIxyM0tFg0yeyKdWB2WelzPfDquAE0FVC
FFKcX15v2zCrA2X77MpPmQXmOrlROqKSgfZlioUkzQSzMISOSo1AMBNB8G1iEDGtu062+m8Rd71M
HPliJkqPR76BwKUih66VLB5BNPcsouhpm4TfyvhJHrhwglm0B4fzWUKms/+diAGq1GKouQ5wSUuW
zQqGohslsW+udCnX2x+ZrtPp0jpcxvMLeHBGS4f4d2DlIYO0qCaImCmqFHVk3KvdbMcJxvDhuuWL
lT+EMNhhTs51S5FC2fsYydmMYJZ/T+mjqmoa824czj2pi2BHJonYu/fyzylDXLH6C3VBmngxlraY
kCSAYYIoMFVUSdzvCNoIGqRmuG2KK7lgB3XSA8Gg4PkbIa9UOwO/pDk85bB/x9IvMvlsYiN5Zd4+
LKWKsNsfCYFiWzpRj72z+Rw2Z6A+aEl4Oh3/ZIqSNNDur/fhxmod5EnbSHknneImCLZR/sQ4HPv8
6NMqwYZ+dTFi7tqcpzQZnw2ms6Fv9VGIVwfOJhKza76aaFtZJV6yORWuPAQpvkdd+UJ4ENtPl0eH
55xVchhAp63e+5Ovb+AE0TdrV7x6sQPWgM/o0FJ8/3N0VVbu2IbLbeTNoyS1eQkiKc1x6atlKBpA
+1JX+jkWR/TkdABG1/NboOX4E56c9D6aCHNkt7Yno+YJmZpna4SUbYm1kWPLKpLclD5LOmhbJ0ve
phKYk2av/uwJ/9Rz/Jd9RDyuAsWfU8fswlC2HV7Iiy6JX/aqzJdRV6v1vcbQZbWHAEZvD8IWGPpO
Vk95/gk3Spw9lThlT/yQH+i2/j3PytviAVD1J645er438LKQCrOL1jGyZdY9zgNcbhNRpoZS1SyW
z0z5rwNJllBeKlLIxH0Qum8z2lnPmmxW0P38D17ApxP+73Ag5yek9kGtS9opommxxTe9ho1TzzNz
g3kUUhEhhXM2+c6j2KoTnqrXzucnGmwxpbQK8U4b9EeLKXPrtIvIFVspklDQ6aVQNO5w5XU0dq/v
id3Qfc/9A3iKvjO1ZR5CC2LurnKmLMzT0KAAM/7lASX+DePuRsP5pF/eKbxN/TH5BQwMj71RByWL
cVtF9LL36lXSqVXNMWq1CewgemumAZRerVo4035qCe5HINCXKmYcj4V1UkpUXR0CDReVFyt6jE3c
+ZaD4m6u5LBJARyB+ECptKJaI9IkIUkZ8FGknXbffL5KMBVN7exi99ezKLI8jXbbTLdYDfqbX3uL
XLzXVKyf9ryZylSFZvNt4UWjq9Whs5D4ndLzpY2k8ReCELeKOMrZwFC8by02cjYrlDT1J/qWt/8A
69ieeTviF2HQ7qY+ZnnlGqJFlsjMB0AmLX2YjOWNatjyHwhZzqpKCs+80/UHjlO5pJS5X4C3fw+Q
YCMhVo3R/CUXSgHzFCLhtcwwLaDujFZoAG474PHsCMK0sVhet62jc3mZs2vR649YtmZGhkQ/VvuB
OXIP1LghX/mvHbo+awP9p5gcbmikp5rX/riDvW3cIvtao11CjTLe582p2Zd5OG7bwLXvTHK4e+4u
DyY7rPqyvoZLwX2Br1dei6X/taLJYp17YEIjjbO7yTuA5q0PyAPxhkwvXT4vUrWOXNBMpikBa0rR
eFpykRk/t7SqPpT+f1jTFMsuRec6URyiq6pdmqeRWvc/W+qL6/Q0QyEPH+1zwHYBYVw9vtAZgDMj
riiBb+aWb8z1FZ2HPrVAHLQLQTw7Un/bmqYJWT76Nm2ykrF3G/aNmETEmg9HuFZPSrryVZmGbAOJ
nVjK3XUY8XHXID7X1UUp4lVvfP6nqiX+Yxn8J0wZRLhpw3reoDvh4VNegAwBcbYa67YnrJw742HO
gayke23xvVz/Oz0wU4C4cpSuqpflaNrGl57Kkl7B5lTxk3NeIbtga0sTNP42G5YoQgZI8B3boziv
go215FXU6osMguoKMM3vsVKy9a3CWR4jvViR8UlFM34ezyRjmCvc4Lvygdl9/li06nWV79A+HuA8
Sp5H6WBjsiMd47xMkLqMzYz142CDKFbhdyZEbKu+o+Uv7GDf8qnkRmihi+XV7oPO+HtuS2VhE2Bv
LjYzsTVe+w36vH6NZPnzKF431kBHSdH2/b7J3GV76CAu3in7SKhHz/t0foS/vSaCInxo3YXhGqWv
J2cXNc2H21SFTa9eV21fRbv8UAANFICnknRHwRxHQ+43PlRb+CAasTDQKGRSHQIbP3Sk6pojiz7Z
EjhH6HymNtr1DcW4YmcCua6wF61AAgHwEzmHRfJq82EBwzJFv8VCxseIZemQ1HyGqMBJvclelByR
Y3s/SmD5gURj6D/IsARReoMbpcq2qsm49ZgrR4JhN5EU5m9aPeqmu6YedUnUbaQp/cCWvOJ2AzlO
a87GiD51Roqjy2rtOD0ASTpsX3k/WA5G7jh/bQs0E0cgJymm000DTks9V2Y5GifqA//vjB2hCpf4
fJLaROh/7+AOoFLyqdyxdEImuxrCdnaTVlqsvzUhbJIE2deOl8vcX7q4rNDvs0JAncpSqvxjuwYm
wqfkAm1cGvEooD5Kfu21KJnY41RFH5NCWTtV57Te2i8m/6y7oxErnCvVQrw13VOFeTGnhBDDYbeA
2wi3v1sp8aqqP7s/8AgtD73quYIxwFMyJMxYRmQ93mf1WLCcJt0G/rlmUd8ko3WpUALxRBc6g3bO
5qSxvi8o+eCoXmYTBjq70knM/6pz+Gxz2W4YSuHIpX6BeiWDYUSPYz8blBu2LBdH0rSta3p16PD9
E95IS88sjUrywpE/YlI/0KNUmpkAQ1bYDhAt2B3JYscAqSXfqg8GFqkEWMsKqY6HDKhzgzWmF2Mr
8HFDUWit09FVvf5+U6HnCmwUHGPmEv0iTppDaA9Reup6GjsZ5/GXC2B3ezUoM/DPMsi14X5NAolY
Ae/YiLh3d0gMpURsLUFC0a8Hyp9ZT8ZYlfUGpNhXJxPqUdcWYgzNG3a83oSj0PR2WHBZ6qNEFjOn
jt6nFtaBT52tczbnPRrdT3JsWtGrrx29OP8KVKvCLTEbM7xbvJE4FaLqQSP/g7de+QVxRoEzx5VF
KI8v9bg5fo/S4flm6KZeFxIMm8FuE+LWtL6Zx/mcZ+pjreFxV+V1wekIynLST/qscDrrHUfd4QFq
zKVIJQAMTNUhj5INvx23TbMP/4/XzL1vErQyL+QtLqEoB1/2trwhJQiQQsJOahNK/x2yaI9AjCiH
KcsB/VzIuKjwPVeBOrnrVAmnzPNBdD+tsd7bhGRZ91IowQSSxYlP2rUhdRmCyGMs8eXmm/HIuVn6
F+nUan+8o7xGOXnbeBZyFaWkaQCy+VmOE5LAhOx6U717n0RFwMnwPEwZbJhz7P62Cx94ERlgw93y
OdJr9RkcrSWhXUpRAWkrxPQKxFIErzNeoBxshoJfwoSqVS9k/4KChXtXyLis+mo1XczFAV4UKYyd
EYlttx++a9+jDuLf8DvDXMKpGj0ADKO7BLdsmnZL6rZgWfm5eGNLuQw5VmsfbV5OwhbnGXy9BWB5
B/raH/obVk84woYUi1bzzgjn9UxgOLe+BwTc9qRnNeb/TCcD8R0fHLIxt4PxDbAzfo2NuBRDMM5Q
yr5rNjoohYGGXWUH9y2DfwaIFmn6mcmceC5WSQ/4p9om6hMN7wssISoHDOwtDdMAqzC3xWjEsD62
uundhgJLeCDGE4svuUin8v0hYCP/O4+sIoTJ01CaHyHTU06oApjrNMbyPZ55zObbWNyY1T73zGhE
TkxQVnPOblFSmaf1KBmsmE6UtZdqr+R+PPvMOs0zSoowBdmewQ28UO3WRclyubuuZdV6eu5Gpoa8
dSuF6103yvLsxWzH6PlonJnWJ/Wk4x52VP0W4tGxXsoIo16xrwPM+sXL3CmmE8mqOHDiA8H5EX/H
/BA4EoZW/rSj71Zr2dGqaxYspb/KnF/YBCrgE8/G1jGWYb6vQzCim4yaneGh5IvaPTc9nsnX8/c8
7jb81hgKIN9jTKVBCgFl1+jXBr4rHLkyJGHjpZFqfdY/xyBe7lQVM+JW2NG4dH7i5fDSnrvR3NH4
5lcrVRg5KZ4LTQPDmTOhxi4Ni24UUU2eS5/rV/TantlzX/TryEIjHQK9qyDMCfr9OL4tADnaNC+t
QBvVu6F9ibgVF6OMLVw37Km7nPusD7nW6kZblLK4ZuPsOTPqhPgCVy9V7634W3MN7HWjnGek679A
5NzbJ16JBkyXvcoRB6RnPcpedVGvqYVAxG+edbgkNoH+1DQIBeCxo5ufm0JcoEkzDCIWz1GlqO7b
3eMTBbLUmd5XH64V0DTE006CY0kUdfwT67tiaeGcz3gogbw8DPIpEnH7CNLTbtrYKfouMw7ocu/3
j4U4gWB9obyMzAil8D209VT5f01H9w4EcVcIR5z266iKAZPGx0k8K1QMiuedHaRaTbok6kEa5ySR
STJxfmCrtZT3wwpcfMZDd8RjQyNHL3SQy3WQ5muPRHn6LTZpafCji0cwBfeKwQbM1N4bWoOzO6Ln
UmNng85wnutrW8c1BANO3H+ry1SG4w417vlAr5pzvzQKdLxdqkkanBzp3IPmzjvKxzjuHFI4/PYo
Av5qYA8Nd1htGMBzQgtDsLCpqN1vKqeZb19TfCiJd6aHEq5LzWVKDnMGp3STLPg1CEXxUcyVqp/T
I6wcSlEIBKyOwDFmwH8/j515/pdRM6QOdbhbuF6zcbjJf+w/DdstJRkEVpZsxs6MFTIgL1lqWoAK
2HsBepMn4ONNy846ruAjCap0AeKhCG14srrKzrfIoYtBt/cqIDeb0izffLlv0jZmNjdBxZf3i59K
hGYkuoBrfx/fiPqgQV6VfM9B7y+PDi8wilF3cViKQrHr0zS94FNuIdp9RiVyJNnelOHsWG1X6oYL
SIK3I4sFGWve4PD2rbVKshscmG05cyfd1ElfeiIlU2S7SEi4T2fjhsuNVBH/5NIUdnrtoSlZDU0k
qm/3OziWSj3CCym6ZlUz6sME7OXXcBonkMxEaLbZ8zHunwlKiKyJ5qCOfa3lYay71PGcf8TjYw1Y
VHD/bv7s/GCvaEqNaLX7RKoE21XlX2d4b4WAQfly0mwsWXcdV8ILEsGM485F1M1RgUUX1/8+8iQD
FmK/fvKwsBQW9KWBoFxnMaQDI1caFapsyZXdDZTojtbXBv3TzWi77FZaH2bpgZaWPUAEUUsW63Mo
7bbnLZPMGuArFEuEO+DIyGcnDTV91Grz10Kq2DEVJu8zJyUG1uEm8kggo3R7ak6B8xRFVKUcbAez
4WyJ6/tplyeut5/lRUjIyS98xreEtaiGFaQfoAY7yiDRmsHD1eysi2F0NOCZzdhiPPgAKkdzo3ns
YjEetXbyfONG0taTecZRZ4ai1/4tXWFrrUwvbqBZOfyjLoC/sG7jJRxJz+Qn/PicHmAGnboUfug5
5GcnjQKZqnXhH4fOJeQag5jzttfH4mBMHqdUNYH3MalP7Edk/BPLDoZUvS36Fmb5lreVCR+IzoUg
3FFpkxTY4Ym4/2ecSbajKe5A18oOPnMvxO7nMZ1Sk7WFuATRJam+rBOeUGcLf7ZnM9hPg5SS8UPc
ZMGGH7juarKIvI+PEB9ltzR2+zd08ZspwN/3uWMBVTKC2owi4SDYsdWLRKmMWussIJMdR8nqxvnh
HfhM+gSbxWv+KIjmfgnTx64wiYnYuzrighdFKq81YgYPQuODPjzjSV2eOsS6hlsPIF9k2P4NPn60
a1HSU1VvHCZmdRPpKeXgwbn/YNeaUuUyF39Avcco71a+W+pi8KRoXlOCTgcWsiPILSbQynI30Oz1
6uv8d5VjyADRw08VaUtVfeTRQePAFT9gstpOfq9nl3w8IAwZ111Wh6epD/GPsEWvR8OgSWx+QEEK
4gQOIHxwJKBKE/TyMaSVKJFKUqhRzS2z3cb6CMUWeT731IWiGx6E1r19TxUwDN8bXpevwv1zzTLA
ek/HmMeClVbYx3R8ouqqJjwgzGryZgPZokeDZpsmjjzrGRXtebqXiVLxFWkuVVnHatBhSvHtYcKo
P7+/Tf4ixVbSQk4hBcroFvsz+8KzYWwj+NOsY6GuEZERolhOOiDQ0agv4ii3YPO4K/lzDfZgj5mx
rciahtHaySnVUuTTbAhMo3abf4pZHbL99xi24fs1JU5mvneowxdbuPHnayhEbs3mRMFE3xWBxV0H
oVVo8VS4Ert0TxlOV8oj7NdXwb5QmmUJX0hweQVP/54OqhVHPRwPI0Om7LTr+XZX83NB4E3Bxj34
Y2nhItLVhzuDdRC8PWxBnFqFT+qqtfjROiQczyhut6YBwFjia+4Y5Q9PHdvfA5x6ms/6fGFWoBBY
zlGFT/Px5+iBgX5/JbZjfq3ikaT0KUe2juiiqMxLKVDR1yCvp7vsKM/MN6o4SqUvpoCJyNdlnIt4
b+XguJCI7si+V0HYm7LWdCpaPyFry5BRijuIq+GyC2sAbFCBCa4ZN1n0OvpAguVT7zNtTWbCMcUl
mIMnII+TryyvTvgeFkd9IXE4ii0EdEJnFmqlWEae4fawRCPwCVoCKv2CFHelwX7biOa4YYpKY+qV
UbJodxY561nPMM5JMbgyyM1oZLbDdwNYvooJ9O6zljJF49VjeGYrOfwrt+LeNyE7tNl1JxTXLAlZ
AVoLkAUjIvWKkqETahvWkSKoay4ZWvuyY3lyF/+zzgrBvq6pWEYc10D2cwrItibqk9tEV75+oMaY
Scr+w6JCBSymTWDkK0G8YBQLII8G9lXP0frWpLlJSqsMWlG3Eviac5pd/ydavRVIOH9Q4LB+CZsq
DGNz/I2PjpPcRr2/MVE0yEshWYVL/RsDVoUFSwYUmDlUW9ODysojvEGEaOhfaKS+olBnBMmCMXdQ
b/gYvI7cdEaeNPIupG5Drr3WvOBinorThsa3QnaoG2y8UGQgjoiD3Ck1jbaccKEeEuF4eeTkrv0B
rt4h47sizr/zMGDZYuZGQ8Rjx7wkKAMXUdXMax4LK8O9bCKgB9oo9HtpXQgs9vCkr+A51NnaAeGp
dCVrnSdrZ0F57wDYpVW3rmbtuD0IJoPekTbUJWqoR4o6Yu52oP49oOo/3/h2FoL1ASXwNjSDVSf4
Sh/3xsIX7UCFK4qyEEsaZWlDctHSTbQuESMBPa0X+Jq3j6RePZrVTSWDdDKMknreYQC+qSHAwQuQ
nC7/EgNgVCK2bdeOKEBGeAKHWgcN/JbXVZ++yI25jTm7L49XNriNTcNFYgUWvaRuDAyRLmOzaQFZ
kmiLmadDlS9ulxdWuS6ObIqR5tISN6Zom5KHWWiMkM7mSm9rEa+02YxB7no+CkHUk3FR4ZohJuxQ
c4v06W2fYbh1No+vjAQ/G9zR7yuqtRmHGXkRFcn+IytX3vZc2FiEDF3bsPRyd2sLgyoWyzR/uxBI
5L7hIgJsUqtDxro/w5gewDuOTA21ckds3XVY/Qy3dkrD6y0UfTDWLOUtfYfCNFOhwgE8hUQRLfmi
OD4zjS/hA0/oEvcVtLjTh5r8uQNFv84EkAbU3lC2I4l3sr/CK2eCeFF5JgHeLfZTOWEguT0bZv2b
Di6oRpBx4fNTr1z/nw7QW7aed4O2SPeOkBKVj1eiW1MtmwiWsnQwcfpz1ZNPplywuGAqX5fF18pv
3gfF08IIu7Pcm1gzWy3BU2Xbogh2i1hUFN/BO0EQ6O+WhzYb/zIzpC3ebFHumLNDxRdHx441JqM6
9prHIcx6IWniqyug2Sbn9pMZ+odC1LVRK4DYjhFfUXLJclMldj6RJsG14/q7/ye4NOcOgAT9OoUm
UIH6t7wmXuBkqc9zG3zjdiM4fDm5Wb2wX/DFhnfqSmt0Ag2rqQIpJz5gan3TY6xHZM8MTYlxB3CM
Use6fvjCJCrl0bshdUdiOTe65pKEb5ohsTb7gqpjfIkIfsTUQtbO8lunX1zg7Dt1n9LJVBcGA7xC
Za68wQ7dg4rGHsoLL1aV4NPyq/kS6qYw/HuUOkAJjXu54pXU9If1dthy9KszasW4MyzqBz0tHw7P
p/PwnUkABidJrQa02FP9yYv510OQyYeHcpHsB/536qpf0desbcjLZyAT+XZQ9UYooo4DoQjkaxzn
cQaKppd45ST2YxArUzh5HPIZbOg39kL7oQbi8A6bJfkv1jACVnMZLpeKB1vEhqV/9hhm1iNSLgp9
VXcYLAgbSmDsv9RRg/DNtnx1lUtGwPVY5eC9ozqf8s/ZeSh86lwYsqHbd5qo1QOfQggY+y4U/10D
ZZdwlMoya4OUUq3NRiKjblAmHQB3dvZ2ZJs4mIbjTSMEQqsnG+ESGkztOlIPvlj1DdcOUshNCZ12
D1wuoHYhAu6xp10kSmcraU+1J1JWqAqaz4OoOK+EAIidFJWKEOGrQxmfHzKnYOIw6BCgkxXZBHfb
gfBSWk5IjB0VyEyFbSvPd31FM2ndX2igXgOb/gUcJquxAnYJVOKp5qsKZP2mQFUvascSDw8/52Kd
ojI2RP3yIDfgexQp/hVtFPdeS4vvZMVhaSuAlzb+sf34wzZEZ+3xIRcN8OC//GeliWGDSvbQ/lbI
kOxT2xKkEgISpXEHWtXKRze1G6qpq08RHztXa4yC2nIJWe/HH0GS1GsRirqTSjErQ940jJHE4tFH
4yZGfbK+fFMV4zlQQMrXqAF+IvpvrGwogM8Y4k6TiBoWVwkoOuCS5ZWo5NopqThfzhqNVKCjuTTA
xYG/lSRs0Ye9RN0SgiDRuQZNwHLOn47MKo8KMv7klwpwfJmtsQF6/zcJ1ZGDRnIqYzLy96H9xiWe
pZbaHYuvfbV43wXplamtY0Kxo+ikZkdKw11ACn4Df27pSyZ5mvFg3KGzWRwFuivzI9B3nKg0aYcb
CfaaVuQnb6CpEwDmqi+AzEaKYWSIY95LCVPTGvCsYCU8U78bqVm+8EptP3tXyEdckvzdwQGr3epH
lKwMTKMpN6CHO2SQdjP/r/zYFTq2okNCAXcFB6kLdGapKKLkSopYs4bXzR0KZTOqNOtX9Ucu7Ifg
RJ87ACl1P6VnMe39rh2XFq+R3aGbDi0R/RCHTABDMD+zxovvqrqIeRs4wJ+mEs8TuvA+pqHW7VIy
+vDL46xq9GNX1i1KQE0RW0MRqZ85Xll9wU4EbBSaRvi3jJ7EwXiousOxmToHDl/OghaClfndYgSO
OSAlSowWBXUxvTqzlNKS/vZ2J4wMLcgN5sNlQwY3+CHSXPO4in3oZCf1cF2OFoPHD3SSyX522fRX
hacOm7eW1Nt/XWxP+xqvkHJPVkrCQTeO/LxGFj1+9PlqfGXZqDIJnD0m0HhBg756V6EPIuFm26w+
S8Mi1terbXFGon/kqIQbKKtZ79qK9fQJdkw4s0e+I7kS/CKSJQysqjC70mhFDQs1iKpO72ax24Lg
5af/Si/umaJ6SzRkdRgAaJl9pBWDs0yL+z+OvAhzozhx5WdycUDAm0FWjHNp1V46lBnhhAFJZuJC
gnGzzv3B8iW6pVhgIQ+Gf+I007ykL7wyu/niKnJtOb8t8gu5hzj0TD3wDMxxOFthMrEiElOFPhPW
3n6+Ae19HmQ1+5o2Dd5VRU83J7Hq2CKjyS4qe8J0WydweJv7eNOjEfC0EKvQ8vmqiSsuCAGEhxQw
LM7M4lD8nqZz0nAGhnYtIDOY5EdOra388/OFOl7oI8x62YpG7V5V3GjSrk9wUozJnf5zIannnRqg
Wc+Cc63ilk1weoMVAdW8LZT7FuDF2wVgMgkURJrujrSeB8sdpW0euWX63Bqm5/rPl2A1mr1F2ATb
fjq0PLKkB74vXlpTnVVWXAVuax5MFd1eOwOBMiOclG//GuO8VN7YiVHkifZMx2x2Sx7Q2SDBMaJ6
gwIAM60PQwPsfIuc5KkixBl2/Jf49MrJpmI9u6tasV3TL3TkLhI1oKIQq3p8X58BfOVcqib9wVG1
D9UFJG/NzrL15dAlW/iqEJUXss/g+F6jpV5/2rmpBrLBVoVT7VTrzyQvqsrDE6tn6IAqQVtgkbg0
EVF1fRxe0Fb0hGYV4baMbFfzkpUllqsf4dgZOSixGCWDD1nU7WSCiKPQsSE4vNpX8VxR8bh/dI6v
Cuf0Ihvtl9dcrrGeTkNxOlXD79IC/y0iSzf8hEh+z6ligQ3+L5cYD0I0LbYlM+RRhzROlI6hlxBA
KdZgP5WC0iVnNOyIKPLno40mr6sNVwNerMYgP1Hm0H5d3LsIP21CyJvbVcQTwtmyeGkPAkuaPbPX
57n0Be+wO6woiWEjkknnpkujJXYgQaq0c44B+HhayVzWQJ7mdXyEtQLrNVrpUFWjsCDXkKVP2aRj
/l3y5/ErS9K/fWAuJ2qBzpbhPYdeQAW0dqspcmBOuiH5g8L0KlVv1Tg+/jiEAsJmzrbC1HTnd12A
jwLanDTafC9eD7EHuoUyy/95aomP8CLEdkmChIynCr2vMmWnEMeRweoIzvwH7bFK489FeCVdPAEs
BwzqaocUpChQNZhJIGID1bIasUyg0kS+BN3HoMv8WZ1QJ/E5rC4ispZH5bwN4m6VDtBoV7/p4Rds
MJNLiLW9MiVDmZaJPlic1aVNR5QZTfcCjKru9fgt/oJCzmVOwkyY3cSpZSWilFmexABaylMMHRAe
QhA8SqMYrKHBF1q3hfq0jNo3t48PPtL1De6OKemdcGRwUboxoFhT/MZS9jshQ5OIW1K4cpGyxkRJ
Soi6CqLFELGd4FSB0NSOwJhv8Xa8M9LphWdoUP6VRANyOwoGAh7o7EXL6S3haCVQwC6kjLALPdNl
yAaAzF1QmBRgIabmdpFSeluf/wXJdnVZYtfhpmtmg4KqFPzyKXAAhB5UryNROJS41h5dTdk668+2
BJaYB44hI9y5tpgyHEUvFE/gOpC4HzyMRMk1kPN6Efm45BzhmqGqbbi0J/L89LxKDUfjC6OvUa53
pOEZd6zC2UOgiu+GXV2Qe4Yhdmz5/qlX562ahOl0aflNnmPHSmBo6jBP1BAmC+leYRu0o7D9LqzS
r6hb0438R377dFycQVElFqOsJTSbc9lCKeZ2TO5KFS+q3hu6aL2P2htfw813cT/eVryWKzopow4u
m/p8uJj/aeU33T+X7XWb7M9V5GjhTVDnQlKrRdpZ0cD3LOIZ1Au6vO2kfCs4GpdFkjrul0N7rn+8
fgIhR98kp1rfHuFeImpBfSL2h0Bx+kEMdUXMWmWsc5brlyn+CnCpHV/aZAKUFbwHS++k4rJUx+gs
osk3cJcWnT1/5wHTz1o48avgav23XBMCr2u4h5E7RxKEtgQ1213+Na1VhXeUZoyTvuRHGlgOs6tY
NAXdmbr7yvIkbhfEzJ4qqsnHVg/Wux0pfsU5sYp+BqMLbbC0smf0jf8gKPobbtcadfXwJK9cYHEt
l3wtfOI5GFkKWgxZV6RP6jRp1bKXMOAdmiXvL6AWzv/uz1OLT143blhm42rswka+nRbxZGA/wMyW
afqWNnX0vtoBnsPIxTzgbgKKGnWO7Qv0VCpSjymzfMO+YLYlHHmrQdy+MlZjsOtxoLCq+vjJJA6K
wwvX+CiEt6RH71Gk8zyUrZHs9z7B8RrlGIIsxu+uaYMLUshB15LCaqkBBjAm6BZKaeSpLOruPnyy
gY4R86mypK7IljzseOI7oJom7IxsSOywpkHdKMYkCV9CcRI8pu7FhItnsFbHi0r1v7GtiHbU4b+U
hwcACQdKH/sccRD3kLZg+iSKVZ4oUzdFoKQYu2cJ2nnGeyP3ujGGvGYmJ9dnGxKDs+5aP47yr4gE
Yp/t8Wsrww1PI91cd6983Ws6Ej4+hGQsEU7JF8qIMIFj6DblHmHVrGlcpKkz0F6Qbjnbg1tGuxU3
zGHGxYqeJSTPyQuksu0GxsdgoRYFcFUZF2Dwm/9kcqAvzJFkOmXWr16FIImmB/4L+bLGoIwecpS1
gQyvDCLt0ldph0I9PF3WzOmhoYcTW6k+VbVgxRvPSci+omM/mFSJa840+u9sPMZJzzljoI/gtrd6
IIt9t76fbhXylmN06d2HFI7AJQrKSbYPLrYNDu+JrWB0ygDoWt1N2x26HlPBIyVVmKHSH442YroT
JGsTd0F3Wjux6lsyeYo0XU/esdpqa9VRCd6gA4hXMkZNNJ7168UzKSFsrsboDBei3KGvb9xTvr34
2pU1AASMrAwFIF+uF4VtZf0crKdu9gJCm0RZyena4P+D0zAUYi+aXzU9PJiwV+OCQfxK4G0oCnkA
wjqB+Hd0OCtnfygCwS0NlCSDW0lXqKlXHLnrM+9sbbPtpaK2xXbUWiWdcrMxK/+kTa1Gm5M2ZTHh
3Jd8u8u620mr9JqwirteoMiYu1Bt3i9CZtH+5/4MtFqYF/dCDLFEHjOlv6YFE4O7yqia/38EQfxg
Ig0XaaodUC72CCA/Ba7cK+iRwRz5IKdZQqS3tN6SECmEQUd6Q3Eh2xR+TbhRbT7RTkvjq8rQ3EpW
DgQBbtHB0WiD1j8d5eB32AfuPL2boztQP++ZaZwHmsuGspdsxWYnv6eGF2hShTRt3rZmyZdJ/ee9
i7/hd8kAst4z+ysdjpdVwvK1oSNpKY/NwYpeK/uyCeELzPPYZVNnt+l09hRcCadbl0kdwgosgAfy
3EcR8cQ3TiR3+arTvYHSZujmp+tYxuQGKLa9wtnJNSF2wp7guyZZaooCerVf8Guo95BJcSXf2QHo
81hdYA13NDuBqSh/zyhFT8dsh5Ek8k4SjuQK4kUYYhitQRhcwEuyTA7HnQZb3nZcF8OFObPDwP+4
7P0xXGDbnwWlSdUNZ4CSTTRn85az2yk6smmT1nb3ieh4qFimfMa1KG8swFDmQ4IeCzKdaVDdn8l8
/ILL7Uq31/B00vRt20RECWOiqQRSQvmdgQBw5dBiQdyNxBWH8vZ1C9jEQWSdqZwN09nn6IAIRuJg
WznKRlFWPZFUFNkb8GbKis5daDz+KTq1D7yQviH1G03T6o2xvyH4E+RWJFEztlXU+cYG5H/Lxsn8
Cc4GyAwtLJganlD/fdST0xUuZbdooH+1vXlBwB4REAsoBJ+8C4GGA6qppy4C4S2a8K3GAOnX61D3
hpHyDC2QGKCMEy4JzB3ukG0x0nVWjl9NpKVErYmN6GiCqQ+Qb/DJEEqaN6wWkcLgLMQBCRsJI6GW
Lo5liJeDIInEZyZcJ048iKGzFKepfxg6Gu3/bwH1cMNm/7mm6GRvt+QJuCPMNqrTxDBP0X2beXGE
+HmB0Bt8ChHsXJgv6Dxa22UsYunkftoLKzsP3etXlPkbNf074nwfLnQHpSG0Pws4hCEJWjGpfx+c
6ibiZ2PkkIvbhodkCqeQtJ+M8O0ALTiXvF4XxY67YZ2NTvVXKe9OTIGc6MabD4laSsOQhzdInfjc
mxYveQdXbFvLuWP4BgOuQFGeLBsZHdjkFOA0Zu6Ref1bHMIAF9ESwzYS7HR/ANVZ60ONXvayJJD7
3dHdIF5IYMDdbhEWmcXqoyJ39qyFC6BO2xLHBxGNTXRqfyvYtV4CKFi1QmRabfDAB4QzhVETGtL3
QJhV5kRMtut2J7ydPNNFAs9xot4IE7W5LCq0581+tWLt2V82ZSlqbkKv5C2JneX3zDkZC35udA2g
OksF/J3/xFdqG2Vqf3JsN27+3SPhZ526rUb054h1IK/wV/807o/t74GOYFJpoPjhbpIMHGaV6Qc1
ppSHBmaf0GkXMRL4H8p6F6Gb4rGtO+wc47JeGE2nz61Osn9HCYMFe768+Mf0muaU4FvNvT/wYw63
jxJLrMPetz6Ab3l0b0JNRSMhy5CSWidh/uWiVMI+Ufr1hnzdnlG1ktUqyQzy+U7P26o1w5kKayT8
O4PYq9HprGQVoeM/ewXw+dW8U3abHHgs+aMvnm/vcWIyjLsret/PWF92OeIH5hyGZDNJ7ZJQJwB9
0QVSar8+itndVpgomvZKKPCwnnEqUNeqMsAapL67tuhwr/lkv51YCPjAbNDYCQtqUOCuFSBZSzeW
jDvfnViZaUuc0cA2hyuSapaMZCnjvNFJVdhpaoBBjozRflyoKJK/J2kEJ9rrIcXwDgBlmd7+6wPb
nfXlFTBVMYnE925KeAceCEm4d6s7YRYK3HHYGMizM7XNoVNSKoP61rthZQtV8Hpa+U5mfCDGE2LP
cM6qvFW3nhuYh6FuDjKuZ84LhrAMpuQhdMyifILpN+xssERyZljcrQ0tiSxm/u7EV19lybjgceVR
fxGc3cnhq9ojChqMG75fCso7BDJX4MZEFjyIe9BP97eCMj9NZIKs5FgsFyALS5oT1CGrZh9teMPc
M2zE0Yu/YslaQ53fEA82RDWH9LWa36BdvmhlrOkxTn4uTdPDd1fvQg4Cxs+dlxBsQCmh7s3cN3BZ
mtCEM42P60HSCrhL4FeVT1YdpNkWFtxMw/+dQWG2gfhthW7/zIY+8OqhtB1sIMkMz+Ex/ItXppxt
mlvGOVO/HZFVYcXsu8urksrabzcSwmiCCObQ/SpW8wI1QeTdzTjZeoyXXGRSjZ/OLwqb6f4E5bqA
EXfVCjasJOY7my4Kgbv6sN4V10Y1XdOgMvhVdMpMdb7jioOjVuPnZiTdVsRxxs7xO5D3tU3Ju0CY
o1wFD34QpVlMkejDut90VMmrrGWRhH/l7up8SnqsAno4jpONdNYkS5KGzr1IBxo6DXKKkZsJp1FJ
q+VNfWX2/ASMdSkSwsFWhBQS7u7DWkgOKF9PcOG1JHCqB4PaTr0mRE9Gmc1qNBEFytqhRyAOgGcn
NmqQpU5ewyvUfpP9sE+zcXqLNlM74DfyOyWx5YZfHjgt6ECbUkSVSlA8KdGsbY27pFQki7IQyfI8
xeezbBjrnm13qRNxxFTDbm9fNFjYarDhSzBp6g57P/VcK/px7KbVTugcOVcsL4C9jyt/ahR1Gr9g
KEM1OyCS7z5P/Cl76JVRV+VA0/3B9dkR5gaOb/yE/k1Oi+mwJ+OhoYmrU+VgMv411kuUsCnm4vr9
7kaFAWpB8VKQgr/uK/E3TcK8IKIhj4GprrNegfvOZWIkM3gwGjmPJMsfpnMjH3ESivcq1ozStTTl
jxIgl4kY34eLjyqdtWoGw0fpvFuEbQLew7SuBneI3vdu3tLH2/2qF2E+fWJ/2Tp+WzQi0Ux6Pwsh
sdtIBFeRL2A+xuC6kyHdIZcquxt0s7Wmdus7ai5DnXbehheaT702yXo+OvgK7fxR2CSRlvifKjrR
+yuYtLPIu6wAyH3M1pWg//9DsBbWZqemdChY0IUCTkWa92iTvLi+mKxyFlVWSjzRJCBTVc9Y5yMv
6tPnJ9BwsEOB25Mdw63h3ziUW4taehPlLtvos2gOnO11zjcNMZYF17zavnyAUMlMKPYQCexBfI04
TL5QvkJdLwmN+3sTGtfG5q8E7oDQ1GYJyDyZ1+QBqpffi7OMJBUePYpdEYlz4Mz7cWTu0jd9YvVi
YULwJbtbPdwe0mRk8Iq6/UMoVLSLD2HmzdI9ZrUuo0taPmnGOcFb+GDxgxi0bLb8AR26o5fxfZGR
2dDsoGw9+6n7gFTnOHcorOVuzTfpUUNYw4JOqlzc/H/rDTfjP2yXm7dzgXx/bKoZZ8XS5GOdKQ2V
x301RRJRR35iswbPJroMJ3EsyQZbpjBTNpg06aWRiFxhva1ABd+Kq6prUr72sUnVXxyKF+8Mu0AW
UQQaCqrgl8kmJmHEaZkeX+r7FKeYpq4wcMaXZxTf95ocFs7xFidyVJs0JYajDAs8WlMhyjSJW7d6
wOtu2UQjnOctiqBbgcg2TUgi/VlH7bKEhO+IEA63CJWIpb6c7JT0YFBLeqInLzEipDxyRE+Cxq17
dHeUzngIimibWeyLRs6Sgy6qcHqODOTQ83CnlGKhxOA5rfSS1KobPKgtP6z2BWce9RLpGzkYlMos
l3Lq3RAo0MzRbHIg3C0h7kY3gw3olT+t25dHfy21m9lRhWL1EklyqvqNvEjXLHbj9TWqX2IFZ3a1
5SSMTI3hCXKvMCPioP/+4tC/mhoN/13DHiZefVhqcYNPWYPqkwj4ISEJ4N9XnRgskcd6RhfzNarr
bPesB9U4BXtgQELk4LbcMoOUSPsNz+LC2PNkVApu5n9Cj39XmqpxBX/lGu1FqPTKZx488iR2ckb3
26YqWg4ROc40AlCnmfYksnLJbFNBV05UNVpM1H53hSDccBihQIbvSeqk3T4+E/wavEdw1syrJVs9
VNWIedntz0/lwsJISsjX/VHjGdUtYg+sPQzu1y0LN4TnCkKdFKGK/08m3WKHiqiF5LOnQjoUyKLk
kSNiSt4EraCPqXoTbVapkLGSBjZdaDhfeQMZ1v6NnOVt6fQd1eB6VN5Brf3ZVonzGaAWVFuaxSDN
rVXLgLUzrC+prfUhiMArAMRxxMrVnxjaKIhzthpbYvDm4AlUYo/maOd/JkCRnQkC7JyjAOmJEW4N
sgg/eGqQhH2kjoXYkIeeyHSPCjwe8t3m63IGjh03OuTE+7ba9nV61SxBoxGOv5PLkOmaKZqt1oUM
i86vKJ84kscKqK85lzoVDCkn173IZksubcl83DyZp7D5MaGDkm7ANXl6+hZ7zCUCMom/8W25Y352
T6D/SzMx4Xx8YRJyFMB2lA1VkQejHWIxwywcDwawUX6Y3bvJAcj30YEdJOf4XBlRP+XW7wXlxB6O
PByDSf2kL/H9jYVSOhdhKY6XCvqFZTJsh9oBjTatVHLMTX8VO+mRx0D7razIb5BCkQ1ByFKnr8C1
AtSb1joPZElaz60l8V71wuRkvvA63gvL+0GbVTGEITSzSf7oiemgn6nD1a9R1oUgo3GipTehU0Om
VehuwvDBGSUfMRWtHmJmu33n53AQT23ICDwAA1DvSRS4rSH53weHVOPvcpoxkottwAyXNBXA/qoY
Bj6oNpu5qm19VH5DBJistORN9Rw4C29K2wq//1NHpqhoIglaH0VM5YVWPIh/IkpZGbQpa7vqGZ0e
dgrLmWaHHDy3lO+WsIvnH04DYwdB8/JDf5IzEXDqNJ6FK95BSwSW6PKYKMWm2XSjJktjDeqradVP
u81tIcidJZQnvD2bzzEm0PtLd6D8sEpvvuw5TO3t56Qg1SZwlACcwBjXc5r3w2ThC6TmTlKo2YGk
lq8n5qYIlHNwUtYmvzd9EONrvwJMqiWnPCZ2u+1kt4BwRsWs40cf9Zzdr81gPiyMLAJUcxDbtAco
nmfjLY1BjXeC1dpWVwGZaKeJAJuzIkYzJYe/Y8wdEOGXviq+IkAE3uWsQ9LqpE8BB5ymTIxdz1Lc
5LrzJDBlY3LuaVLzcrw6MyHw/OBQKRQ264UCaR3MfrsfaMfRzGGcT4sZiSGTSLeMD+xS2v/wCjEa
NYzKcZgNviyolIrQQu+8ogWNnYd9IK87SO5Bb5BA5y6EkO1Hxk61fkZ9wpyjMNmGr7GRHo8pJa2H
srz4hpDQRoOMfALjWzqC5MMXK0y2q4+fUOyRbkj8O1SSZxzPNhP929E9SKjGwSrKIVDQGG4m2ZO2
i+7CxpkJPpwTkhwFiq8hyR9tvepkDU16RhhQqnC+yUaHHpqanw8j2uhVhRc+qgrkeipehUHBzYDN
aJiI2eW8jZmkQ0VHcSptwewkE8+04Tq0FTGG36GBLLW2LaVKA78v+jIxXdHcOnrbgjPu/yLlfdTC
Ha2waPTor3b1NVBylVz1AjBn7S9etIPeh+LvVsICNZwH5HIrDT9049zODVR1+eLYEPcUWxkJoyoR
3S9vrBDWDwcVzx+k8aQC220EMqkM+3RKSBsmja/mDSafw46PKld0H3NDWfg5oDJn7NO4JY9zDJsL
1TU3n0AC0s2JO7Yr82gD0u5dZsbb3okEwBZI/9qu+zesdfI1YmBVrF1cN0r1fQRW1Z9Q0K75/pFl
NWxD4wHBgp35bwFW4+oF11iWUmDYyyA2KLVYio1vPWjoky02pAFv29sohh0N9+5b1CGyn4FkdgHI
FPnSDNo033JzuXP0E8wJfWR+1Fwtz2UcoOo1TPT+zjIZlsS5DswcnXL+DRhXlaaAjaCdyM7tmh9f
Ad41xZjVpsYTrpc6JHGMECi7TbTcRofMgna+1UtuZRZ3SXa6iHafHuOmWcWJoTwTkK6Ml3KiU/M/
Hf3B5OULvhNPMUyEB9MbR6ylsIpKLTdkzAIdc8PtWwuyin64QgDPofbN88Bf50VQgzK1sGMNMmvz
xBMxrH40dy+cv/Z9EUIfJEDo4vAtTl6LQDydPvJulsdaBai6Zzpgo1Rap2X4+EEBCn41lnZjPdK/
0GRbJhYRqu4RtfnSOjaX75j6YP6TO6OSouU8kzEt8g95WQRATkM5qqqtZXzh+LYzh6Xpj7m0jH19
6ImB5Q+lyLGtoMRYxDa36+CjWpsBygcKvozN4Zppc6g7Fqe+nTiLYVcUaLh2uYqvaNXHAAEvZFt+
CcpiRzdKIePBKfOTIaLYymDYX2P0NElq00ye6hrScDBibt/hSFwZmlFYhbeppcPp2d9E2FAgOrnj
cKwSsYS34ivWDrHQrMpWHPgO4U9kyDlTxjHdwraEd5RzK7TdZrCuPZNUBQ6t3WmK6LiLRd/O6XSd
fQD8OFDovuvzvbVb5bSq9lXl4ueABNE3Xgh9E64PjgpPH4SHau6JZ6yQydn3SRIxL/y0EEyw8noM
vwKF1+o4Q5HIylOS3nImo3WELKnvg7orvidBc3VvjGJF6XweBBokDdfV7Lqpm25qwQCjl9atGceT
GplPLKxtStFG8RO5pf8oDkjNf9zSuuRiKddYGDE2Q6qwtnybW1CI9RJ9ENsI/ppECe9vN01N2WHT
5x8R3mVVWWKJoZzTwm6NDjt7B3NF63Vh2cyoFSy6XMKapONeUPIA9yxxbn+cSwBxiG8TXrt/Eu3y
hPfLy4Hw833LZH9hpSEy2lHwVfNvsEmbMy/ea97vCmyVoveXu3creLwOK62FFSUYeYlLlpBGeRKk
vewAC9cx3ny25l70rKeu6N3nIfijGtsxqlDqfKTbM9sau1yMB1DVoOeZCyG5lZHeyanW60jdvgDC
UNxovFZ08y3hYvc9DPPDJBBP8/FP4MobjJTfB9sbqTMYMDTxHvkilngkqr8oPs4+Q6AeRgtS6lyS
RuyMz4UUbxDJp1ystaMSjyBXXR5vRWDLAPqa7p+5EIujnvwHApA8iiQGkpshFGBHnxOwF7TMqyf4
KVKOBQIUUXf/SQ0rNIrm7ritmKNoHTzqW1+0XyyWaHxOBpvVV+W6s6e9XtQmfBsY5w5+20m1FEXk
0kUah0SJaSyRKpNWzXNomDV/KmB09KJmBwBM/Q50pG8/h/w5uTyqBf6Re0+NKomuuQzpvAQG7Pj3
qFGpmYhUt2ZgofxPuobwTb0ByPZQs86BkW0bGxL9f4hYhrpZjhfE4qWfbs4dK0eif9I/l6Rq4r7K
KHHZzRjxxEIk/5VT6xwce7LjnVj4MHGvDj0zZ87p+X6QiWe9s514I2xsN+YmGcnS9wO47SCvAzuR
F4YeMALfM1xMJEGRrFjgmkgExSqqViMOOF2eLWJPkDN2OlqX6Rb9X534woTtakGRiDNmCzkd10KY
MeOTvCz0QB6TzTd2Wf5NgImzspGEMmCkpsc4Z8iBtE3mtGl6ykFFHgNkBcKZT0MkbvMfw2Mn1J4m
OZ+8Uox0EIaa/It63/ljrYwP0nvwcb+Ghr2aHB6IdZbDivnLHERPA+tRL1OiEyjAlzndoSmSu0em
OnYAdg3huGLd5Wi/nNsbS2ofgnkvDYyMjnpSbqKUOoR7Gu5+cIx23HuYZl/b40UoaopfAsBdliL9
PzUT6W9nbSRnmcqaZnyPLCNhXH2ssrv0VcKK67WERNER3pnLVkMIwuVDxTWwbzJR9+8g0L3VrZpI
Uc0lC4aTQWUM8hYY+hG0L0gfgkqDKAoHxQ+kNq/6cZP+HGd9v/pcKDVJZquNDSJ4s4mYWDWRIWHx
HeJxYRWu4msaQD2JtiDIJSdidben8yYynkFLlC/qqjFUeGFOvfEqEz0uw9Mmpb+scK0GOw5b6csg
UcfMKFsPcE/4I4cuDEnGCeUjrqI7+MeaR4P/RP3PZ8vmLzUhxwZz9JsL7tMsHylfkQ0/9F86W01K
1hAmtNowc8CAtuy4PEsQFqzE0mXQzuCxqy2jlWAU/iX4i6/DujDpVb3/aI0ADL2unKQViQh3X6ZL
28jSALz4RKvoEf/6OLwMNNS2LyPmJJpc2cYQfe4/2aBM5yIEUKAZRIMxrkTe2fh9emYx4ztCpcr4
mfrlgnufSqyikKq828IdvGESCDVzuUwChHZrAzaUHqhIWasvI13QIHpqVKaqQTRvbsUx85a5vR6d
LFNG5U1sXE8UJGatZghKLzDCz6keHnA1Tzu/sSalM9BMuWiJjwT25N6knVqIZ73YewE6zL7VIjL4
sxBbsUi+NdBtMZyqYFe0zT/KunUG3A6cxC4vIsdlfG1NWeleLPM226RnS5TgP3fYR6f4KoFL6KhF
VnEO6PsAUYLKeHlUKyHa6mqJ/yXgJ4lJfDgTLN5K4ATZ18Ke9w88ykDvQ43SsPvxWYzvuolWvRoN
Wi/J1ayAY2+KdGllm4z4z9iR8u4IeYCaZty9HWfMEgfQqB53pTXNBvN+viDNKhoGNQEnK0rVsEJb
gIttbVs7rB0gz6E3uCoa1jHvCXjGsgYg0if3lJbIcV1/v/XQGlEc0DojDnxF6pogaMkU4mo/9LTF
TMv5L8gm1nBbEBmG+cs/CSiYcfR8MBLP3a9yvUCJw7sme1KN8gDHZnmF7AlEK6ER88M5GNQw7FYR
gklAwJaMg0z5ioCILHpZKDIj8TV2foxgKTejvs7mKz0PWVcZ8q7iWEicKZcvkJ73dD+d/tfDVOpm
C+kFgmNYA889GJ3EUmG6c7+upPyaZ5BFhIc3Fh4F+qy2P4hfgspWU89OMo+6F/ibyuTCtOIP/Cmv
DA89/jWiii4xI0bO/F/z5Zm9BtO52I8/idNx+6kwFhqLeDlDSW/a+QLBAc4q+ALbbqL7spTnG/rL
HiUio9VG91bTUisQkwko55JJt4ScTOo3hyKNfZAVO5Cp8fFHTFfO3zrshf8lMYHyXKnnIUOGJcO0
6/VpALF6NWVirKDzvFHBHkQVr15tVE+HwM9/P0FzYiLJeiVbD8yozzFuhuHRk2LV80pAq+znUtFE
jiKuxrOXXQ9ZMEV6+Y6d6qqKGoHv/CYr3KyC6a2g3iZgDXOmL/o0qCL3BBEGeuLLFsdmH5H3Tnvu
C41L1Wng0BzqUakTfE56APddVruM9qosu6mIi//agdU9sAiJy4AjNSUQS1syD0cu91MIf9DoGSP0
UZbygBYHBRHIEdLnImKGVxxYO3EEIeju4DlP2tyan4KCloxpdh72mylFaw+ZrdXiKqAvhpzjFaSo
A+Ejmi5CAcxgZfqrrpl8EW7f+zCDP3RRmkTzdfHF4ggbsv5s1oQYn9OrscY2+V7c2XAI+wxW8sc+
0NQLXX6xNlzVvhoz0HmwF4RYXB5Bpk46t2o43eMfSM/ft1PUWocQKEquAk1prVAP7HbNtvfpSwP5
+OT5sRLA2A2/3r89gWjTaqg+ivzg2/Yd7hJrwBSdHWewSFCj+vlsSJZg1HyB4z2CRO+VZZUXkIR0
oNdqxxmyZqkpKltLI/tICLN9H/LIFRAonJhyuSygQwi66sbI7XIGOot/yphDB/Xi5wIp//KRBUP9
vOvui7+7BoSZOkiw3fwl7T6ZC2RN0iHpDbQ0r2kadGL2tksSA0VCFNZimLk6LC63xvSakZAg7W9M
y/y1DvE1yJjnnPpb6m2UivVX0QFGVCXiSw35f8s7IAqEawj9z3lYeFkVTM93zcNXl0BmlZjrPUHF
I2rRsAi3FkERhhiH9Jin7Wbb6Q1T05jP/mS6hMdbNrBYW2Z9Z8tzuJ8iWqJ7rg7iRfvY+G2Ok3Jc
wP/mtYIcUHvTSFPSpiz/fNovWPY5W96ThiF1+Webi+6WRZKfnlG8TA/TluoQK5mXtNQcJPtuJvmD
Y779q2AnQPpKMBN8G3hL+Zc5eiQpVCcx3ZNBH6t8E5SxZtTaQg+WfAbt6+dPdn2Fv3iUvZjvQMJt
6vrntymetLg+vK6Cl/zIFaMZiNnxcjC3mqfceOJMhutqVouaijwt6AvICPsIXxcYpZ/yqAY8u5C+
16//4ognK66O9CUN5XzWWRClYy0WR+xc9FcSnuh+93QZOlCu9EYD9fsQPmqKiNJ2WJyV9adof/Fn
hDJv4TmGnyL7JNZYVsUB7aMQwnuriI1hs1jJCBpVrkj3XQPy4KvwsRW0ZzeCfItuF3UhUeTrQcED
9XdWXDLDQHtwj33xjjn2QBM2ZtZllQGa2XTgFWcUW3CzSx5IZb+mIpEZOJ4JWtAz+0jl0P3FytZX
Q5SItiLLCvT2pfxkX0jTX+6L+8AURQLv/94XLZo2ZWa3GDtNnbPcxFHcbVM7rCjlswipNAFNcmiw
HvtOsKgiZoCzfr5BosiMGFgXOOAyC7EWLPVjCBJnL2S6Ehw7KNaZzhF1VXCzb/a9JXMmFthKZbpI
PTAqzSl8XujzehHnV7peRWrPhnmVEqjdC52jjU6yjZnE84+RBK7qJG9uWkjs7/rsbW8voqq/ECcF
ub4V+LMdNx62NaZx5bm6BIl9h9U2aobWD60JfNoLddincauNUi6gnNuI/2C9Spd9ofoQMIYswLJC
NYvx2fQFOcD3tvR+Q5YznCjYUDUha4p4Q25N+8JJj1xVWUB6aYHRZdkCSZheKlASQ4M0ciSqLw5A
QFL4vZda93Z/HDN4SmCI2klM6Vx2tnMWgi3M80f3jwwO3+/pvI3BvI5IjofxobYhdloVEtUu81FM
5HuFSEgVXUiwAvFuJ4KyZBtHXEr96tRPjqp3la4ZU4wWrcC5W6FC+fFYkcscKeAj6tNx+Smg5W9W
PDR5cDk7VSTAJ1Qz9v4IPEXcorcEZSyGYLa8UwlY4we7w6Ol1Sh3yiceWk9DZTn9dFsptLYaMlic
/kUAbLLhEQFHqnoeKHAicamLzJ29LfU9DJk1Vbut8aJRZY+LpJUKarTOz68HfPb4Nx1JMlP0VLTG
4eRNB0fFGFWkmVC2UvvKO+j7olKlbIKYG4XFzl9yQCh6rpldGJLc8asYtWEF7F45DygkxCuvl941
QQvcczu/Pg7Z4hKSzAzx8FcSC1R0dWrZnCeEmYuFKx4nFJoLyAstmKLzwZP64/sUQsR1uw9xT6Yo
c1DpXh11DLh9H8vY+woRrK0KKfZEc62yulePjLPh50MeMMM6KpzOdwRHwbcJWg7D6ZoQuT3q6FSQ
TalLWxP8QFxSZ3Xfv8uSV+XAe2JGPQQrnnNNEznvkXNTUKTQYMPNU92cof96TPywUDDxUdSNMkgi
Dxga579N0oneOcFIpwxwM5QgCyWGoBBaCAZH1ofLQ0RtG/VAL/yDZ2kUVEUIbNIiAoF997lGrf4x
knF0VgzvDqvg146TuzHV9tl0iuo/Ay0WaxZGYX2LDq4NELcsV78TrQU3+TjO3eg/l0Yxn6sJOQid
T/aUZrbDubuoOzQ0WrHYn1wj6zDh8NouBIswPu9k2qf9TkL+lmByTU8kMDY/SVH+1snjOMMJ5d71
uOf9knnPOtZdV8DVNAyKfHw+y2oBXVhz6qRZsZpOikPh7A2yqYilDhtunddKRbhMOqUES3Yczp74
tPzpOKiswEk5l/z7ANpLiVihNMP37n2pWy6njD99oqi65YrEOJRHENcU+Z3nRmAMQ/s1LpTlaC59
zCkLUJAfTvhHaOlJHOPAQC992TcmEHe8f4Ys2QyrW2WPKz1ZcHCanfpwIetQeo52x7KsJPCAzjdg
hrzqDTfUSLQx8mfV7+1Uu69LGQdcu3lR11wDqFaw+gQvqFsIDpmrnKK6EoT1MhkUZr+5/1V5mdRT
S747+vGfhguq7spjHFkWPeL6l07K3qGJz+c2+GyjiExJ/hrrXhuTt7ysCZ1DC0W4DspOEYNMQLSR
cGWO90OMZjQReLStrG+D+hCTmrQ85GlURXjErAPPf75BW7d6z/wu1IZdvz84mAhCcgKMsEnxP4OJ
hOn+5/eo3OlQhua3CXDu1X0cnrw1lN1vmFuu8+sLgLzUdjlY6eytW/3ZdxDfyeFJuN/Pcp5k6v0G
PSSbYpN6gF9lu2Hlaf+/3jJOulKVJRYBmZ1E6cbKdxCAUAQK9qTSrvLrRSkAY+3Ngk1dqkOvbl2f
i2d5KS9KLFSEIJ1tOj+OIYJUpNO8mnLkGw+bNPB5EEodEX/BJDdJ2o+aElfgu8daxvRvND8WqXmW
B7tRBTUeCNcyqlz3w20OSCvyDhcak9xx/9NoU0iB+a3f1tsIyWXrehPT4riDC3ycTsgbhszs2VlS
CyraJBQQq5zEuSIRTYQ9pUOvMv8bn2vzNjBQg+4u8WXBVKL/ZhjyL6sbpSJAgaZYKhFK/P4QMNLd
gQAikSu4hBrCumNImzn79Jt9Q+Fg0DX7tIYZbAujz3cY02swWUSIQYv7EWsm2yRg+ONNxhXNHzoi
ows3NFc+h+QKkPo/d1W0ahdqoEbUJuhPAzXu619BjHU/qBp4jeFf/Jm8T/XwoYZbaY0hslcs/MLV
A+t3aYinpkQcDOTcvWtM9yBjDgiDUp5Bg9s776TO07TL4fIVIsEb1AuwPbCDzPdZYAfKdv6ye2cp
kWyjqcrDl8uiRRSgbWrX6/jdwcewRnuZy3aAlh98dq0nKNSfMV53Aw09/YVdYamuga3iczvT9v2m
NIfU6VLAcboy8NMJiyi7K7HbljBtdcsaqKHXpYnScYxQSpRGvLhcPg5nO1RECtYnuwdSIbwddoEH
Qvk4aoxS+gDZMg0frP0Nqz2ME2/lfITCSywnmIK+Gs8k+92joyNNsMYl+9Hu02YD+fU9kEH7rCSR
8vu+YtE0IQDLu4D9+7/xIBA5fUpfalZxguw5S8xRUPq2U5KeMq9/ahd3fVURdTYOdypNH+nJwOQQ
MjTrLKJsYv8YFIZ+N/v89G6rkcgt78261ckNW9ieNZ6fxLv4QJ1J85k7lolr1VSkY9YTk3TOpnb7
jsHk/UGz8tKhQo7nRjM5S66Q884FROEIIzTfMyFRAqSsyceBUFUqe5b7tIErO3yfiyT8O25OI0qi
J75fVwgDo4kVlFJToknkk5/vzwIYz/9WVqCCdwY8oAQ37L7aXyFlJBAJk5R8e73iLB2P6JRECLeG
wyMFLTI/TMVtFU4/1zO3w22krtp6BQcDNpVbElhLSw1Vt9U5DXwwsFXqiGWefTpjjWrv1iEaNVkq
JCNf5kcdlVqyz3vikiVMdYAE0N4d3Z5L2DwW2lFcLl0mU7KdtZl7FFc2OmtSsrRdUTcfMJFWS1WH
d6fSeHUVqwK471mEjJOFHUAJ4HxXIfi7a4tuzYCzy/0lSw0wlp+wB9FMe5P4dsAYmeiAob5I0ijr
mxLZOIKD5rJbBKRMXej4nj3V/Kvl/m3pCkcjueaDC0CFqnbbRLDKCQSR83qHhupKQ7/MC0xA87Pi
kFRzSE/Djfm7sCDoxn9FEs+ibXzdPH07CKDrNhNibdE75DKnyrNZIhmXCBdd0l4ynVXn3UDfbd0J
GjpcQgr6se1E1bEB2QnqmoLw0HWTD0M3iazM3c/fWrV3aIF8w8UCx9WAHpJxg/WWlHpfxKTJDj7W
9qqIDBNuD5pARZBWWHWFdHXqtzIZkARsZEXShQTTOT9QI8Ji58JQk+M4szt2IlY/yYA628NfRP0X
xjjZzqdZMEJhjFWDKsbzfLRXH6DUCJGzMnixY9gqW7utFcBT6XzR5F2UX3q2zqUavHEKo+FVpYXX
SBfDxgxx0A82pZBAzSbeen+eRxm955pi0qb6qzkMrzPw3+e7ow/irT2lTBOsUITLLLBrfD4EaVFX
p/AMjIfnKBNLY5pJTMDtX7kAfkXmLGlMRJqOjzI9Yco47Y8ykTvAGt76QSjIPjUBsvx8FE1BOZUO
QU1vMDY1w3PwOMXmHR816y5bmj50d3UiKh2Kj/dT2MC/YoulVrSdmfmpToXz7e3gGZ/KQT6dtCot
7YL90W7WXDmuSGmgBBtjj6aWUnE/Eg524r+ft7N8xVHymatSxIrp8HyQgKa27rO0hPQFTHNSv2hB
VEaKr+xAxkrvYG/GHYQDe3U2HS+G4vBNaooSgSW1xHZGE1p9N3/ma5nBqZtCXX9EDc4702EZPOsd
lrCoMmW9oBqHOVNaPfqg00RqWCATqljzX5EKsq9LabZeSW+IvfahrxlWDGORgmRMK81UaDh5W5I4
MHuYwU0HJih/lhHh6Lp0hC7twoanJX3uYpe3lO7iZ9uHaAdFFiNF+Y7k+n7n70MtbgMnN3CmPjZI
xZ0gwEURD5n6Y5uiR7aHW1pI4sRsiAVCW2O4lVqbp2IkHxRhyYVFEi4IUpajgVkVC2quMIArz+CH
rBOru3/RaRkh87NO5heNVzlaNGt8J3/bJ6sO9Xlba1O3ofGYmxL3q0JFfz+PFXO30FQvCYIORDly
+EVeqoLZqoqBaHEwJ3O8ddfaYZEZUShljRtahslZsY54lUQrsAI7Nog79wbSEN6JYJM+Zv1n/hrh
x2IrLsKhEwGTE/kA3D3Vnvqojgl5a1wcVn6ilWwsKL+enWeNyxgWd4AdcrMakbScmmrBfu+aWpQZ
MiJF4WyOHEo0tI6BNei19RbhBbwbfcNYVSlJVh9nPNZI8AR9pFkOKhAvENCmf0o2W1PnuTo+Ddul
e6+TD4VujmBBx6HKItrQmAl5g6YA+vheRMgs+bVoRTcJJKL1MRWWcNaFsYzBTfe3g8dXP3aB3tw0
yp967GOSJ1VALaYGT84o5NPvYLGPKtScn68r9pWWyzvs7Hr9X61knddVmUDI0mVENDFr4VXmJZ/t
ppCAHZgxoQwDhr6OD6mrXSO1GsQ1Qnj5sWBZrlRSfQXHYuhnMvxs3MTCMk4CPScXMGZxuiR3EgLQ
Xu18k5LdX52yIiQMyFMghKM0jsm7dXjF5QNzOiM/00iVWRrD3NyXEb3MSvHGZsobejgh7ljE6Bqm
Cgxly8SVJLqr9fHn43BlMu3FQElgnIvw0SZCbukjTgWUEu58P3Th5Jr6pi4jqG+8owKUPLIQ/kGS
4y/dOjESCUdRCODUIcSKK7qYZHLcJrqjZcapEuh/CieLP2TiVoMVb70CSxR2/B5o4bE1D8nBVKd8
0LlZLNztsxLjpSG/WxS5972rmr6crrzt0Wpyn6bFCR5Ju3v8bOPMX4T92Lu8XDafDJqUXxgjdslb
2MZ/MK6ddvgVTD7z6Wp7M8E2fqus2MuB4BhirGYI1a9yilFUNktSWG/NdApLheYsz7rleVtPaH6g
r5hXdmIfgSECVUbF1qxQHdeyqrBqo3Q84Ts5n6iGdVAKzM38vti+LP8JvPxxtVO4hjdzg5jqKWGZ
NYvi/I7Pw+Hq8Rf3D9303BtSXOGvBwZ0+BhBwU7JgUumV8OTYphgvy8tiI+bXZe70dOYSXYHvpFt
oOr4WUvzsH8ik9OnlOBA/8o/ZNfRifOa1xGpxIZrnbp+yTw9fbmhs33ais7l6uD9QiTr7+KBoahQ
X3SiqyOqwQi/iOYoDjo8eoTjfjFT4vCSSfBjNc5bVLxjT9HZ4xz57hNugRQusaZRHjvmaLZvkiYn
ZxzP0BUcSiWZvOScW309Rw6ogvHCIpJOzGlCWdFKpkfkVBxATKcJ/jO8bFH5x1nSGeyxM9O7Vi3Y
feyMpdvN0eLsEOjs0AJisAZxWFfMTc2+vql6gMh4HFD4IRYF24iQGDi/0vdvH5Sw25PYeG+o9lOd
Nd1gPOhfOLccuhe/dhjWDxc11zwb+hSCvjZdHLmZ/cwu2QzeNXAwqJevqC/8QIM/pgX1W4JcI+h1
0BYk/wIzaaFSaBFUMcxrkVhXKDoHMrBBp3wB0TvYADlhjp/dqHjLC2srL+zvaaBPVrQ/N7q8msxC
YrTXKs9DZBZ283/RxMkJdPE8cKqJWbp6fcKyCmns092Q7B31bEcohhH0oTiLVv5gzOG+IlNm1ZXH
Wo4IUiQb6HsCF6MEvyaPm7Jsd84MvR3EB797hFvQ+zclWAAcdP4EsWhGI8n2wqhrntEkLoim09Gm
bFi8IQRYiT4mt9mt3mlRSOnkJOTjr4iqO+vi09tVElEAENFH72/VXTgFkpx6aLkSKxyhcDCrPwL2
ftLY1Vyejhp1Zyld9XwQVhTb1p33RoXBRmz6evg5kar/JVAVgWtwdxniVodZDHHo9jZxwIBIDJyo
KW0+hZT6HqyBN1PeQMhXtvChTrNJBxhvLwrRBJD+vyblsSfYhZ7HtVkyXBvwO8LCJ32qDjfoyv73
vRu2rQGWzC97/sFJbPqiICm/E1xhjPK/cKLbkmuUMau/alrIk2QW8DeJnePDJeRYGeqmYjuZkKAp
/JldMvm8yexyKBHjG4dwf8kXXknijce7bjkZ4NpdlrARjW9aXQjPFrPDHifXyv3gY0Aya5EYrn9Q
j0IYbz6MVtxXxDxEO0PMNY9vUI12r81mHF8++PjjPciXuBspNaJbAT444eHFOwDA45nidSG5V2LC
QD5MukPoP5wLyzxgNQA8PVdjM1bUrdeGriv8eBYOsKXYi4nYSmeFGaVumNYuGXAbkNeBONwYoD0Z
Klsg7h012OHzPFjZu08P3ZWvZwCo936woMtlNj4uPv5/rY438VYM4QtcbpHPAr+h3vDHANXCqMib
u/rTlpF3va+4x9EqxGIyR+pOpy9t/mM1+fASRSm1txXy8a4vHHVuGdIOdhukMmjnyFC1hyTZ0qME
M8y7okE0kgxEo0Mqik2QCkKaS7n4p6hqXs8cVYPD7EobsoYnHQ4C1Z5HRtBFCpJBDblgjSEm4kTL
AFwAyvu11eAmWNPsYgNWSYP+zPbOXmwbiZ9dJOu06EyMhg5EgfxQYUptYCc+0uU/zvnBShesTUz8
eYDBokjQiTmetHlA3Q9Z2NL3YZzrv7fNXKBaQmdVrZKvBQ12eLXT/YzRddHxPT/G8PLnV+HRhO2M
gwj6pFPVTF8NIBsPcFqxndWk7UqTzWXx9w/XfwqU/KFQFlhOnTdgKhzPSizNN+f2Gbn75OPGUXy4
pxpGouiLFNxO+REZhvbs/Ug555LYX7CJV7yjkezTy6mc+b10eLwlvpq8vAB8NSvj1uastDxfZWMM
3M8kSs0PJVSLbEsCwfIg9p+rdOqkiLhUp0+YCDUHaVUp2vSIZctsVY1KlBs4nLkfhOy4zOaXltFZ
j4sF40dyO1U+KAzIWcFhQJrGGcvyvj1U7CcBmfXM2ZuFLeO2QQ2hHxfGYtqcHRbWwBRsacWRKoE+
J8QTmvNuLTqlnHvetgzADckR9512758LpzRtBrqFGGhqsDcTZYefSuYUJM3uqTCK0DPJWL50DRyI
LuxAyutrY32NDuPPazg7h1d0UmTZ//BXjckG72XT4YntdFYYxF+Pn7IhAD1tJqdv6wbA8768eLFK
Zsq53ceFO6zhE8VSvJo/3TujO/M+AGa3n3CDnlAeEYFNpl2AH2ek2IySkWkAcE4GQodfmOWdGH5N
JfRJxT7YQ+tXxXuydzkpmcviGZK76ba/N0sn4CoYYdNu+hB+NEDJY03/pp4BRLtkIQ+78bxv+iI5
OxN/D3boPLpP/XmAgTsrcviNalr4oiacXnlymUWRAYlcxjXta8tFAEqOEqok5/G45QpOixly5F8t
9bBezis/EhbNRQF8sC3uDbX20RvM6/zsOwyUlRDlUDnMhZzfmp8OSc4wWT7+CTUFyocLLC2jj1e5
8m+49zV1vHxqngdgQiXyoZD5eU00QeZ94B2BITW1uNkDYfGilPZuxta4vE8dTQasnQv4Q1+LHGP1
fMi2G00adV1ydAPOcbkmDRNyNmaMj2XzNM20CrxopN6fOe349kWsvfJ1eQicXmS4XbR8WUuKzSEO
8Equ2XcIti/aPKYO/tvdyb7eAtJSJu+yqfIeRLfKNzzZanRLFxGuHDuFEnAAic8kybpmhk5Yb5nz
mHyvchNOwQtfb8Xe/SdjCEj97jWmu2sXndVj29uAfGtItGcmI+EazGSPw55+dBNzIAFrZOAwSPCt
wx2fR9bet6278cp7QCc/JPr5BS9TacjoPIAce5pcSP1uy1hdCp6VYzWtHVuNcM4Mc2gnWJ5cB2Yt
kjJjPEzlPtyWVIgmiobvvqWxpRV/eeyl9glHFf0y/FhobVZvmVLK6wXt1i+WfMO/5W8uZhmzvB1o
gdXwZzkuskNWV4mXx5rDNJhw1FoAqG+FVJUMBM0egk7risaEwEkX9TS3Bn5afM32/agb51UgvRhc
nmWm4sjGlYKBFhUBsuOhzQp+WVoWBw0YbupZ0enA6T77NXdyM4UakqAIp6INoTZvHeb7arME9Q1I
WY3BFcidxS1SfYBjjnMRSmq1dOSn0ar07H+C5WScxoxKZQbelb+z3fZ3UGk3srIBzsm+YCZAQh08
I5TzLsLSTuU3YocJxVxjKVK3uZDQB103BRMG1qi77/AceM1zaUBMhC7sWVdmwJoZnff6CrnGmrbd
k0moAkxStlZ18fWlJlw44fZJUPktxoQBZgIH/4wfhxEZDeDwu385e8qYzhDVekVSk1gfrVJXqxB5
Gr0youtA4i+9DqR4vrIwv/sbEXZD2bY3sYhoi0kmY5Vkq1YguIAOeQp0y6QATOPCGdrD+TS10tWC
aBvIhYO1lSiVb9dbzysXnMnSOuG86inv2s9Pkk5PVqDpXB/4WMykZVw6uYmxgtPxALZYapidUYb+
3EyiCYkisQtFwCA9OofldUzZfC/p1nd1jVjVTs24b2B0aLt3oMLry/OTmBJQmOcxHq7PaYyxl+uz
+pZ/07Oc16S6D/kt/fw9hao8mR5XdyaMczfKSZEr8uUS5RV8tBw08gaMnAjdznBAvEjbsdp/Gv6g
xi6vTNwD8lLWgubPZj2mpTHONx1Sm/BAJmoO9kreIvm/wU5f6khEQIh4Ieu5MOJ44qAsV6Cq+bCD
pDBJh/RoqH6ZckTSl7jg45KpvjDnRpuziEddkqOsLab1VZVm4Za6NOM44oryAjutpqwA8taQQG93
VtDnJjWIEN3Ulk/qTVhSlorFS6PqNNT+RClNREU6b2ZOMd7mM5gmNdd0pzvlRIJO/9D4b3QYIfvY
1w99ohyOC33KXtNTRf+CpUQWJb5zJ16SZnpBMWY8n0yJdUYM9geoG64pLMUBYWICZ9NES3U7rtai
VeBNfvskdCAszZA1jrHEu1luSmWrhaZWz9CBEThYrFQJLrq75njJV2QPAjLpz3ippbsFikIQEZ21
QeaFMz/eOhgkqBh9ZCZv5b1d50XGK+J47U7MRgrYWSrxKQZHQ7maDDOIh2yOBwLpmyonb2HAF1tz
zwsYC+vqulqrBR7SNBIOQyOKE4rn2Dzhsbc351UOTLc/p3fWIcyld22QpmIr8mrb9c1ES7/BYXAU
f4aE1azmDtUKqTzIBnNaGFwKBIiifcGOnhWZUqwdY13jZB35Awv57wZgv2/t1WgaMrX4m4kdx0py
G6vzF4JJWdMMFwGbGLFqo9O05wT/s3qJbIWo7MiqEKsKTKZhbIgyKlLFawY4I/8eikU7k4AvGr1n
hKxnRDjZdt8zxLV74szaH65dfHatx34cQKN4Vyi3hLeVMgWbsnodTynM2zu4i5e0uMY1aYaCHdmM
WKxXkZeAbSyV7Ea2aY4vZx8L6TLfpo/sSiG3y2/HuD+76Je8QphIfarab3lB/dpFCcgWdp5xd/bk
RdTTt+KDGrY2nzXFI2SscA/c+a0WYIEX/nA1Rdo+7tEJV2j3bG0HqZsqW1v/sR9bD06nvf4RNEVQ
zL/8DypgGsXvLf1n+Lz18AMvbNgJxJcxcZI8Zw4lFzqqG3HKd/8arJLAdD8Wfgk0dyZ/OGt/3ouO
RLdv9OTeS9aJsb3COLhDmRuFofLSVkis5GVTIM3J4maMtKr1UhNrW/D7N+YWF/TWMUeqApieYL/+
JX4v33GDBehTRWNg4P1gcjOCLyGowgvm6to+dYR/WG3BFUSwH9ekMyAqRKFQv+GOwtpzTrgRHvVg
SaYqUi91SUMAriFcxG7OViqgDZz0EHyN4bRJ8rurdxEmACelW0z+DDguBBhAWLU0YKR7Oex6cOWB
dUOFuKVCkeYFOX68KDyuHg2PI0A6PveXo9lG2jmZyZtGa6uThaOoPprrodv9dzk9/phzAE8DgHpt
73A7MdnMjYJBWm2lO2NqCST91kNDZkcnTHTogIMMvFmA2sT/rSo/qvHcIlZ+IsaTYlvvF2Ws01e2
eT1xxPoPdw/HxZQbW6SlNhc/qC6MJQZtt4sPi83LNqCosUoxCcbZvF7oILfs0KY2QgTmImpMMpy1
iT9+PPNixZi3ejT58bSYu3eJ45uoJM8w93rx2gJk6nofAorjfHqZPnl8tej1JarXKFY9tkC8tC7C
RihKCh9mbgK3Ana7uCMUC88i7WQvTyN0vfHUh+uocWSJanzE/z1l/t+r2Hz/C/fP1qMGG4SItRVd
M2Jb93tf0BCYFD5anfJav0XqEBgJRKW5/ypV1hqm8jzUjKiger5zBrRrQIvrH2osScNn20LFPxm2
gC+CyieFPkVUPjqSyrjdrYRnpGiRTFawJGYJwTD0lG72TgfUNbljiaMwydQb9elfE2SzMp8bow0G
vYKKtW6gjgGjK8aL+0Drtm9y5mS5nbiAQEXAJRDIRt6PtNrsKIJquzpOb+GEy3iK6kv+RnKsh0Fq
MEdfSSqiMtBxdctGj2eZMmXyg8ytFkKSDpwLm+abAuDr7rEDFK3isj6R8/aGbou+E4aOVtNiCz1L
tikd7/kmCjm08tk+XlulHMlJ/mUU/wHSKKwKwl+oH7BiAWBmtfZicrqnC5xynjxfvkGWPiJLItCE
kL9OpthdjzgngKJt0YWWKbmpRAEb9E2gE81Ghy/grjpGEUbdEb7fdFdIHXHiAI/gHxjm/0V1Kc7+
5f5JrQ033A25WkGweSpO08ZYlzmxTSqKfsa8vEMcYPicWbZ4r7ymp2e677bMF3XfxBmFELsRRNB3
xY7Mm3ndeqYUE5vi1TfeXBD4+o8M2t2MpXcAYPAVefjpszTlHUDuP9/JXX8rX3YrM0tVbmMXUHO9
Jw7X7/smkh7AJ3qNyj7MHO5IwjqKkJMWCgdptekQ4UtwQ30OnQn0cc+9+hqPcejFAMrAXT1EIN5g
Ujm4w8jldXL7X6Yj2Mn7bMgax34+6qhJWghhZkmsIH1YfGWiSHG9bZCkeB8lgDzYIAEtnq4lOgQk
q4dUxBQkV4HHKJKvurRlM0SOwKf4VwfnZHZcfYnU2pTpYMutZvsTCWwxEflSr4HjbS1KadoPYcqE
bGelzYDqGAy4HsBe3JHkSAkEc91OHjOny/kfCBRdeZDAIctDWK4a+7CPSSwvLfHLyo313PP6MLsc
oVsVnhiwUy8ldCO9i++TmXxzDZnPy1mh66RjucH3060lqPG1uv0keVSFm42jvNSa+LwjKmzLvhgK
oal5IpbHgR+dK1iuSjNAIlkd/o1eEqX/9AzYuVJVQ0FqkOKdETCrt3z+u9DVA5u6Neh1VbMeS8fR
bjWHMRaWF3R59/KL0EBkHnC7XYCXJqhn9Yfwq/iw58LQlDufG+7ln2+E+mZco3d3M7h6RIgs0K3R
5QOnh5+CI8O0yNPLQpoO8tScbFXx55KtGgiglVzOYqWBlNfr8FnAWhI26sUjMQ+SU4X/k9n6XS75
FKGBJole+0k4RNRxr0nVI1ztxNQOHmssQaLVATsutTQH7uLV7vcFtdHr0yLEu5nHkNIat0YSekLk
VUYNgcAJf9hasGuwWxPWIDPR4TPbyD6GAVW6nrisVJXB5oIbPpOee1xnJcUOP6SVJqQGJkUC9Hy1
iTvDsS5KTSGj4+1tmjW8CeEEke33u1Y7HVCg//yuAC0QRsT2Vb7NbLeEFVnbBTsSwcuW9jbJcQMf
H4sjaDE3GKylK9sOV5SWvo4ZTMaYZ9Zly7FuI0P4z6vHKGerN0hUYFHII9BjbiGcAOfjbDdqmmKo
jA2A8Py+xZVPxsyTzfIcUwOSAZrJmiHCgSTDVCHA5m7sW2cHIntCp5W664VpTQcgWCPqlKspa5Kh
6Ii5a+vg0crb0g8HDm65Y/VaOdnNHcBY7XRMljjF9McIDlzy9LfS6Dt8kQpNWYimIku6jPUVe44v
56bnY++lT22HpYg0ci9/VLPE4pj6tTHyim9hsOJbVmfavOXYGbEOcWM5Emz/zMR+iYir5DAOCHrt
AsQ+fV4xLLTaLeN7Vs0fVR79p9ifwQXdDOKodiPqpL2tBTGzNb6Gli24nBAftxvKLcz1WysTw13l
zOHQzWQs7WODTCJs2uVNS8eQuuR71zQrVwyjUSEAEW4maUClqE0bN3CEYqeXHHAdXJ3IRlMPiHO0
alwN0Alfxb8me2on391KpgSi08C/bXm0V6TMpLxroOp2f/pkzcnp14EALW9otvIRYL8HPJv7zdAi
nCIBVsoEV7RYWWybO5zfV7JlhqutzZpDcQR70sxpXmU4vUEd1827rS8lcHYpBvM+OyKL1Om4cAKc
vx1Av5HClQzIqXRd3Yfa0V00m7F1tsSjazxycX5IWyScHfbPRO2e5FntfYG29hO9mslksZSG4wr5
3BaIZ6ttOpwxCN7KMecJLIOgVyu2KALBUIPJOTjJXcwTvyr6uou6fJ9VGHpq/dJKQNt+QcDgmM7A
Dbyic0o9XYnFbg2/QPUABDOur1AADPjCs/ijXegqVPA4LmxxF3Xb1K2LaJgmBR2TXMIMyl7F7S2T
fTkOJghYLnHZGOVix7su0AKtvkSZEamNebVcbWUmNzntFbE5Idnarar/MQu3SzgNU8AFd5D5a5EL
Tu3azXGMW7rUZQfB7In4a9Ma8dRuX0bszr0/NlqMFbO871I8ML/rZ9stKW0Rs2W947yfG1CZcUnz
59sQD8iHGflt9vUwpvXoA9nQsnAkcTQR3+U7dZa8l0ax4w07bUrElzhlBrzGHjFniEyEkYR076wN
G2ZekpzWydSYico3vLcOVQE2esG2YUta1ztbak/jx05xELPho6uIKHV8M9eFF/M2vXRMV6aupzr3
blE8NKOs6OwD9K726dRBIqn//xSPE8UHyuYEwpPQxcfxNk9eJ9GLkvM4VMMKR+FR9xFTF5lx6y3b
CtqMYxqQFnF6wq+dh66IPPHATW2aTFL/CjGM/nfcNjIwyY4IYTQqr1am+5fE1RCJNjsS/cJ/OxIa
cH0xWYKlopmUmuLAhLKiXWTe9w7wnfUHvxWscheAsivtAqUen8fGQ6t2BOdHpCdUdzWfke9Ueib2
sRAgn8rNTkkDDJBIrIpM4Ism/rCcd4Sqka2bTCAd1sNKaVhB6KfqeUBxx2x56LagrIVSKg340bBx
4xJvRdz4maLGRqc6eSmA5vEnB6xrcVd4y8B+HjimhfHBjomWvDtuIgTBGYCa5c7q0dqmRBf9DV+O
kQ5Lso95Ky+vIC9kH2JIYAsQC5KxoD6f6ZtYa4IgLNT6eJSYWDULJZTAWTYBUoKtdzWzRpeFExK6
Jakf4J/eoZ2MjbkRQcQAuHF/w2oRCYwiMtLyT7l6Hgqo1Pm+CMdamBBu4VD+j0SDX0FlNaYB0cTj
N/daQh6dzlkdiPwMgwxOuduVKuAwBpjHmpe4hFdgDXeFvPNPC7uLcZWkr+3O2wJR++83/THKOP8+
Y6oCxVG0L1mla1ZzEv1SYy1vLhVVqn7LbLaPPVXjKBYiUjrgbIHDTVsHF59OnNMsEawB7y9hcpcc
QBzzPki8RDdtMuFbccXOCrT+qIxgGlnsxCAAnC3EKtgr1sKh4Ym0Zf2w53YjuKYA7rmBb7h9Aj+3
+aP8IwXxs+4YnP1555sogGdUEW7zs82avGRoYPXSiv3da8CbgYv6/Pn5l9vuIWyyxYss0YkBBF/M
AlWN/o147MK70/cTNRnp1HiUW6+tM6hnETq+NqoQCuaOsE8UssSdQGTR7b4wodNsV1E/HBBVkJv0
c2FgHUJG5wm4VQ1DWRVXJ52OwOYIEgd5NGfruWGKr2NIDFbU4T7UtYrjT4fjWv43Fj6BRv/Jym8x
xai/V8d3bH7gfQ9lB7SNr+vUm7BFLoXPyESivXOmJ6LZ5HwJPpxKiS/FzuZF8ie4+LlzGIozR622
I0FNv+Pnwu+VO0CMaBcHOg9yM2atEmr86a30cIdE3pijC1c5Mei4UN2CkcBkHn6qO7g6yXlXlUJ9
5zYdXRQkMcPg4Cq5ufVhg0jBdqYviVv8MrWwU+UU7Y4AyGS82b11SAD2FCkiCoPnEs+FmOHK7Hir
wH2hHAvj6pd12LoLNTtsQe0rNN1aBIPqhAK0KjOfFX4WLI62xtKmqQSSUAXeMBsqT25kvnWY1D5A
/xWv7o5YX1nAKq6QFhnuRDwSsNUlZzfZvIFeEyCeIhUT6rjx5O2JTu70p0KdHiGDLBlnvmwhGKp+
KOO9nwvbhS3lfFTyUv17/DqxAqQPb/x4ykLahduvQDJULQWXBGmHXdH76t0nM8eWOG5jXyZXzG72
yAv2w1JUY/EWQLE8C6adENu7Ar+uJxqf3VnmFH02sKHQ2GMKEiZt+AyXcrn2efaZsD0nJXdW6vyL
jdydj55dZn4W4xw6xKTqa3XA9IN6cSxslTXQUCqqVhmd92JJeyRM0psHZuZxPGAbpG6lKRE4a4j3
0TLS/YqwPliNO9w9bWxrrBMyn6L2lg56mx9FaJlZc+SgHcpR1EfB6iMMLveieWy+KivE7xznBlfL
9UIysV9a5Yn5KJ7xSoSq2VH4YeqmhMBiqI5i3ByWwoZngVXM/ymWspABa2YUVDfL3Qa4dEgJqg+K
21tdtv8E5BlVyvkEa4BKJnz9hnvjDoNI9XJZNGsst9JD8730uJ6oTeyxK1pTMAX9wp4iMS+PXVnL
r4YuteQx374o4ieawQQtN5E2qOe9hEqyOIGQxjZwX07fuiAsa9rjaJebx/I8Mt3SX149AhRUwJdm
QVDQEo7ZSrNG/d3xBKniTLhf+FMH61OelQXTo/FWdWg1sIB6xWXJj1tN1tWdsB8tRU5ra7rhT248
YxVsKX27yqo9K+ThOp5i0woTultupUvaKDXYp/bZc8YWkoBHXXjN+LCC+BEi2UkNHa8NBGuFCWjF
ixbCzPaOBGlyIYmeCDJFKRlvqZSPHOmC+aFtMflkUrXRszu3jgcUaBmuZg5oLIqdrNiUjX/chlmx
2eCj722I0P9FK2aynYR3Jk4zEoFakCl4LFxl8Vmwo7mGX1iT6SK7tjHQPdz01xNOdZDm4G5pKPCv
No+Gr60gdUYTLiI/DnUGJh+IAtwqRlflW5phFzWYp9UrRXv6jt4a1TaCQCqsX5uHU/WqxQvximTH
UajZ15IseTRjw7/NJELs6V/qRj2LPJ7ZqgIXPr80S2jkXLk2VLJlFFEtDDXDf7E9Qm7HEbSAEPtT
i/rpFpFhKcSC/A5j/ZH16d0zYNUe8KZ1dWrW0ikl1fBlA3IkBRajvK0fymZIhMEfJ1FtrcHxQf3n
auK32y8HYam5CyUuOds6d7+sT9yybZnqTrcCTEKpUiIozq25OdBzwSKgBxxsKu6rpV0UrFY+/wSe
3GAtpDQtLh4uq0LHO675Df+wF1Ry/9nZd84aL76jWd4Ex8hctYRQENIsxGD0p4tvtJ0mnMAhi7uG
z29Er53v1s9Lpe6Mne25HtvkBpvvBhEFhUnvrMXUZj0qYW2JtO0+L8xviyVTgq1um1liwlRu6S8a
Ya1y9UR/gwMKCacqOqag5/mQWwopbLGnzrmc8DhEtX2XpM5zzVKT+VfmyQQJ/dh6ghfmMW16wigg
w/oUZBNQlecqPbOpJmUN+6Nqo7LqvADkujWtALu80NAJorv1Cq47dA4M6FGu4hA++K6ZCZF6mqDM
qNIY5lcjs/WSeioJYixWfoHJOwA+41MEhFfeZvixPm9eBw9h55ikH1FpHNBUkND3d0+UhCBGlzsf
yJcJxI2JNMHkTOT/1I/JmP1nNXarPug8C4NfBr8PPfnCW6yYakl6+cTGsu3iK4J4pKnoAWMUxEyM
SVkzZy5i3EoXxCHEPk3BbzScjdlRpTzRmL0zvP0/UGESUg8Y2QvGN1qqZeUNnEt4x5nQYZ3gPQXj
PUq7p0/imh9vSmydklsHb/ttCltjPjuQ+AifuI/P+sfZwPyhRME47bsIl2Tnm97eKinqT4+jJ5En
R560ptXeXDExiTUHuQ9FbQVpp/wyjNSdY/01JxIg8n1VfxecX7q2xeYRIDrNhChQ51BlIh0QG1JD
6Yxavzt8l4hxnHMQrr/SsU4SC5Y/NEmKw3/wXTfVEf7EtscKpVEV6dSu4ZcrelQifiZhBzVbzEm7
D4iYdywr2mMT47apc9mdUTUN6nEMc2INELmHYAWGTV6FZ0NjMZw9mzzQme+YqkSAwaWk/Oxit4RH
38Ma05NcT6HRY6ieIVQAd1IG6qTaQhVHddUEdYWrZuDulHlFSU3vD/R6nBk1nMjfSVh/J2HncJod
EWYWKJQDx3lAazThWnhVGOJndMlbKZRfhr0ZLxYyxZDu868mNZObZTHP/LGLCRRX77VEYJpla8Nc
TbFaXFBVq8DZ0/9U274Vorr/iQq+I0SKfc1RY5JO7DnGHv7UY2LR+rXJ8EB4C/yqk5jCkIw5HFCv
FqYVgzdxfXr7C9RFJUNjKUQrPMRifEvEEdDwhJC4icdi0AXkHJX0IflHVKOdU9jFo0+yU2G2rNDn
hFOXYND/PG3E+gQ0BD1YsWYuacEsY5IMnRBhbf8oXqcnFMWeFgi65gke3e6dI/mXhMshumtgbqde
MCzzNXXvf7UAbSTfW0sd/U7YZobn5k3xPvIZ1bqt9bP8V9UdRtzJAvn58vdyWvf/X5aSQ6K8I0Zt
RLrULN4VqZWBM5dw+QQ55YBlPVONqg1rNJ2oTUXnKq8A8uIJ7ZSUJ9494LKABRAwSNTvv7MjAp4C
I3vERQFJqEI67avZPmEKbxHJR0jENdhGb304do2cpGlGjNDzAY4iiFlPmd/fShiaWAZhYpNMn2iL
RUOCDdvzbbIR3QXhpcBz0gfqOK2CqbWqcGDQBwVl22458pNTceZpKPgF6eYsELWlOY8o4GmaWEOz
KGnVEAQRCYalArrYiEtIbhFaJEvBoFhXWThkCC0t5aQ2vc6OgGXAFYJVDQ3VAzA17vGNIf2bZHIO
cK0r6P8MteeN5ydqe7YiaQFzv1CY4f+F1uHGqy1EeAH/nf/ROeECGNzC9OUqQab0qV4jd+sgFe93
8rSi7b/m+RNkovAxiYEq/oEAe14Qvn2kOvwMUWJqT44TjuhC4XhQ5hMK8zWT964Kj1X2Z5wzHnJW
DBkcoIERUsKv48MPXU7noqsyFQt/fMGN9rkViCxGYPuuG1FliAM7PUESA6zLj+t1Fo8AljD7/xjo
sQZAsUK7TS2sybaHG3Hx0YucjOTQQBxzZrnegv74LOdo68Xv+FfvHVlX2+9xw78NgluOpoLKPRkT
uXu8YUujPox5s1hDMnp6kVbUytD7ePAMJxVfhDFgpl7MnI27BUExW9fWybUO0JhbfEoTls4iYtnL
GpP1jP2wjMqh9SPcPLpsNO2P4QJwcF9VfH9VYRBiFgnllZxbyk0ugst119+9P7c+e6iagpI8TQDH
i57igvIlK3ZpcWJl1jgtF9G4wcj9z+8Qr1szKy4NiGmzubqYjkcCXO1D4wGhnAfoTpU0kv36jSVE
Fyow3ldmXDBl3H6Jew1v+qfpqDcZz7O4nvt4Tj0v7uxPvpXPpFvsqdEHzGWJy+mRUx0eMY8l+nP7
7YwNm4XfvY8Xe5QVvY7iXCRc11ycx38zDtUM8hPsH+Fhp+iueT99j9aDrGC/XPPXpOA//j8BR0in
Mu0XY1yjAlIdsu7Z6wlVPi1FZ8BTCBXflg4BzqHFG7Xqk79h+ZCTZdeuwlG0nf9Kpgy4THle02rb
TDKP/975JaXRhqQX513XYjKZgakvE/pf9XE/k8V9IUOF6A6C3ZOs30nW5CwHpciR5CrKf+u2qP78
xApw5VYAweAhmIO8hwT88IbPvppZ7uvnCCU2+Hq2NeOs+s6PVFjEZIXfdi4vopLwEyyBrX/RwKki
JhovdkuueH/dHM1hfQGNk5hUTo0QF8RzQ+KEuluKNWj85ZIq8CFMnMUMnQJYnp6q5Eeh1GBCLJrC
/oTJPnOME02fnyLNeF9pN+1UWD5GjxUCcmA79eIXKYz9IiwLIIeGe2rZe2K5X6EjeCcb9BGqd0Qi
IXPH24oImCZ/3IdFfxuQXRlm0jW+KneDLLuf7xIRaWHF5sbqc4lr1bbyFhgzVu79Oqw2CS46GFIn
w3ZuwI/zU9KfiIib/odwNF7RtQR7z2MjxFgJB5JJQYQ3uY69LmBEiKtOlYVNGuAdN947aRsB7JU3
XVjfUd//AzV1KIWahbnkZm7aLsPAPwjTqqUma3+S3JUBa8wr0IWyGJzmWhN8rlE3WCiUDrH+aPID
P5Z5mSL7cHDIXgaNr7kh9Qddlvm3RMx3IgWpk5AkYuUl3utEnJaQ4O9FK3CZ2N1AmsaImZen8zwS
ehmHwfRjO1+Ynkk7j9Qh9dCQ/H0O92wAB4w8nA2gr/8TdSwuAOdaNqjD0sBOe5KCUZDhjk7Z6kek
d2MpYpCsFGlJsxaGUwKKquVy//noqyUrZ2otj/4e4dMfS9ryLQF1hxK2A7cx3Bj5+oOA5EcbXcbl
zXO9hF0rJLrOTduOJjKA6cDM+a0wQ8zmLv5TAVYUD3ACpsuXJ/ynjpJDc8yKsAyWTelEedi9y8A4
k6TMHyAmpLrot9tRZ12G7HfGLziGD+ay9ja0C9HA4wixLRGsrOOX61H/ENEGR35eGBWQVM2nW15R
MN+TK/gU5RDxg7XM3NooY6YvM+wl/bUHm4fr4UGrEvt7De14wfyu0GfZwO9Ob7ziwWw04LagkWF6
JbGQoV/uCZuEKFMWjsymf8SRoCHe/2tvtzR8y8ApP7tdhwpewtKkohMWPGc51lF0oT/idNz5tzLk
e7W65okWnFbIkd5StkNZQ3ZWOuDePr3NEg2azKtILOYILTx2KSe2lDw2VXDQ66AucxUhECvWpGLV
602p8e3qHA8iX00b95JSJL1S7wrZjlKi1MmJwavdS12rL5tx6ne2C9rKZB/yvxYHXLp2rkEPMD1z
5f6HCG7U6Q3jWhZqKCOm6w/1Em0i/qzLGFCiyiXqA4nTbC9jlmUgVimLKfuKfr/I1DVINX0KJ9/k
Dx+fcgxtw/JSM+dg0Hv6tWvN1T/eBLJOsgh6ZC3XhMBs/vH6/vasKLw+MUIDAASN2h+bVMiu8Cqh
JxaVkpghOP8H/sOjeoVXhOWLVLixd+eZ9NHkqPxwXK8zeHn+WZmPCMl0vXBvM+GSc//Ocuhe21Lb
sZ74DvnRrKh/0dZv5Zp8tdvyRPiglW+Izz0TcVmn+Rbno7V3DrMxbWlErSLuF2mODRBUg01WW380
A9ZOgTvj9D/PGCDs4WzK7G41tlRB1cVzRm0V/HdyfnpiSVhTn6jcPsWLCNEgBVy7RJNrysAdu/bf
Y8UyuprxZCOMCeq0o6n6qa4nRfL0uY5IAOWlvBSif5VPAt0sB6P5XxG7A101YaqdgdWHAs5i62eQ
v+WydFzbJrUdVdPwk6JX29ni40rJ77u+Ra9A4J5joGWhjeBczaOi7og7GGKP3gbQmZQZNPZv9OAQ
GkTm2a4E86r61WeCT4eVkciF0/rC2KjHltQFQiE1JrLuAuBfn6bP0Z8Ly8l0cfVclIHV9EFAuNS2
e52IMIj/NTFx0qarlT7bjh+WHUo5oKaFX6GUHW6YqhcYYjJIRZKAjlc0MLBqeeFFDmgBEGIAPwNp
yWrKrMCh0uHJTZzMJd4SdXur2pepuW4i4/x6+9t5Eh2brzw3Z5oBzfzm1NDkMjkQWNiOiqxdPndZ
ISL/Y4TRg3Gum0nPqlsftjPq14LDsD/ckhZ7GmK9Mh7Gmnw2XxqK8ZJznjtn6kK+HjmEhimqOOmx
3uecmD5uSULHuoSuc7cazKpeboxyaZy768v0ZEqhTGsx/B51VAx8NZqu6hDNa0hBjqTltPLgP1ez
YfPLqwbChlIWL3qejgK93XicsSxndr7mbR7E7DtLTgk47J9+x11vy5c0XslMcvQy/toCCbMwmWD0
HQ+XR9h2ICNSIgfJ4N/1EHlkO2kOzoAQglfnej1BijC1/kLY7nFHDZwIg6KoZWJJn3uhYInKLNv1
pWQ1lijK+B2AGSQbNgBvWPw9YCKMCdaMmctqsTzKEN9wuGLu0UduSXHsU3zTGsITQCLxUVeUjWuo
b5/Prtt9JVOZFod9mq19rrm4uom9SrM2pdPan1DkdWqKWxevzvC6AGpzBoWiDpCp7mCRzR0J+Kj5
iZVDoePxYRwBVyZv0vU+2RVFIyZuP7sbYR9gacso8xbw5ZwCay+L0Y0k+/G8PdkjuHlgqea40JK9
aaBneB3ETbratGAX8TpvaFrR9Elgy79EoAezKmX6ftI36rc6uAApmGKRZwhLW/5KbhVplaP5DjVT
jOhKVL4NfC6Gu2egaCcgZgJNn0qweH8Vlc6R1ANrBZw3VzdohO0yfY8yGrcKhCOlR1ayP6RRx5YD
epTshDyCZZlZYPR4h4DFD15LToagjqrhvb6Mi4WSUx+fz44MUDMvNBpcPaBvLOulkCCc6VdxVS9V
u13G5C42X+Xonx2GhFQBK9fKVCDaxQYT9bfO+OhVEld/PpJC8ZFlsf1SsCedvBSByJvqIhR5Gcgr
x7G2vHxk88fOtzgMfkA7wZucuubxF6alFhzSqSQyvU51d8ChrUsqt/LpHv7M248UckZb6QHbxfD2
nnVmp8oja5QgWDWyza3R2kKmRm0mG9ZuKIU4TLUKEgy6BewmENQzsBsQE+Haad0LGHVaBBiHZVgm
6BGZBNXajDBK5Kp12bdb/1ELTinNWSeqy5kqy6Ru/r2VHozdGSWI+PKU5FgyKzLHTXcuDlUK641p
LLjwC1NKcUlOEGUKL8DLRfNj/esiHvBU2Lgb0DjXo0IBt3IZx9uXZzc26+2BW/NL8EwtniFHGEnt
1jO1UUNSN1aPOt2k8gBFJsSpRXeTft/dy5QQA245VSdPu2H6zUhDgpZS1pnb3vRJq2tqwYY+whhg
miHX0rsKDEI7dymcJvGzP6UJevzeDypdbnJj9wPO9pk+mBQqsrOiDe9o53vAUcz+RL/F2lLiBfQo
puyyjiDy/9vRY++XdVU2mITA7cAVFAa2ZJHCpS0GqCZCiIZhXUyj9yz1MiAXSLm/m70D6uxnai6k
CxE/qHJYZSvWEPTvdzOJPD4RSIu8CL3fyKSipGT+GRuC7P2RxWkmHOt9MBIt6Ce5LX9EvDEVy2Ko
PZOwUHC/3FYEvKXPBc5sbWRX3t5o3m7P+CVkPkjaBe+vXZhTbe06sJSV6vsOhJYwbsnvF/w8PzqA
hCCCLrYXE2pdp9TeIjzbSAILHTLaMZvotA7gmzjtK/nntoAydwHCDdFMvdSkaq2cPf9+sIJA88+w
auVJJKHG/J9/EGnfHl2kwjOya13BWHD8NgIsAsBRd2ySO73SFGqO9bSM94QIPWrg7EVYKNH4S+4O
N+0Ou4gJLqXTm0WwRFl+njYAKdxT+Q7mXh4hcwNxoroTAXSJwJMwE2c5J02aCLwQxsuEY3D5oZk1
3LC7Ojsth6NkbfQE06fPrqBH1rLjupFr1lqgBZBOfIIr32f2WXjv6VAyrYv8qS4BefqSQJWDu0WB
PKpky2Gj+5TcWVKsZRWqre8z8+CLICU14nASW8r2VvrmZCLnTdtl26cUrSSw+qg8rr+UceZfv5p5
gbRC1zQmJE0QCsR/wKGdRYq9uUs1xRjL1EnJIbr1E7kJd4f067qTKty1MwXVKDfOQIdqkOB+URzX
BuP1NbzumxB3/O3lpWLGoFl/RkcyMGv8Flqnp3pNvRd0xRFm71stEWaen6M8Eq/D4zO/DRRLcxA2
y6GNXUYqrPe3fFr3GlfpcCLFi3sNmS10Z4x18PwCb5GbaEVPiR0AiwtDHI6KOWGgbR4fvyaWaOCT
5jYI9kyMo/0T/wGZDJ0oTUFdRg8sTMTkfsf+kJL4dm1uo7uwnsXoopo9x+3iwdCMxbZMrWynZxVb
9VPDRN1qpQQ/ajzjItPVcJxHt4jRIibfFo2KbhvPFSHVk0dlaWp3LQHPaPEh3uTHaZItu3ReouRF
CHBxyp35y/IUSssA3T81dv8dqZId8hlDMuzmI3Ph/Zx7CVddLs7xjgJNp3WdxyMmLvQIidfOFttC
SMZaCxv7AdFNoX7GbU47QSMqkD73L2a2o8dnKijb692+Dfte3LxHKwvgkllGRcvRwkCIMjK5E20N
ZFC6hSKcI5Ftwf0poT5eIyDtihrgROtXKv/JgPX9+B6BfrYzJdv/jGfZRO0YFzAcpfvSTEUjEXYF
X/V2U9E/qt4uuhFwQrdy+kEx0LICS23eRQFnstQChcyOgzRynCI3qlbk02nPkUUCR/fINi+zodrp
VmY1W/6E8ImYsX/WFnUrR4VziM5QPdfHL9JF/ldbMHKcnNuZfDXKzPnQ8E1RiMpB3n6aS70Lc3Px
mde3r3kwGL2FFDKIxGoTL2p6SHEeYx8tEiXWZB21XQKElWwTYIUm9NCWeBkhXxLx3MaUOYmozXHN
judE0mcziwOHUWsXJr9oU0+4V1qFd6lhosKMK2/fKRbX6wYa0SYwV9X4RocK0w2R5CSO0z4NES5l
wCaT6aXzsYiBNjGme4dhZivNIcULL9lTydENMMyyv0uzGUGbzrJPbBXPzC6hIZ7h0PUDbGWT1kyO
Ov9GvbfTXcXURHSr3VRIkRNmPZxQfbmzDlkXCvzhNzHnjUf61h20iX9I6Ao6uGIN7tu5aclm5pax
q6L5FW7tmbqNok8loGySZf5jUWSVBEWrdWyVq8PqXc1lTIMefh8ZMMHfr5B2JzytiduV0Izi2Z0p
it0laKhNKyJ+U5HmLF4w6lZsZTkLhCE/98J7sABdNSRipdTfXEl47ABawk3UnS6FvCAxHyvv/jM0
oibidl8C2X5FcZEXfVr7Wkl4erYnuTISix55esvMgIlG86ycuMkV4qxjXB4DfGvpVPTO99GolIiU
dx35t1Fe3TnlKck+xRO4tT3o+S0CdK0N9FCCanDUIazQRx0I+tcjIaHqZPQWyLaNfkt1qXyBPacn
9omdEP307pVRyiz3ji/lsScuNkhtG+2gF3vBodMlZn7Pij9TsiwpIQvVk5xXtf0So/h0ie4jyoWX
CkhmqUMJlleWe49ro5ZAUH3TkmBdBifDWSQJLrRIFQZajh5vpJsL9Rrismix46gCVA9nkrmbdbfK
FtfzJbrad1favXnNfcHwb6bXS1ZOESmx4K3tyZAg4dlX956DvkzR3z7dvp0kK2oGJ9lmnm7DHkKg
TFM2hTEB9dpfXe3F4InZRYOSPidBYTnBRnIRCJ/O9dsuae1nTvYj4hLpTsfTheMII/FEHApNpa+r
56Pcx0lc0sPFYjIdyyWruorwOVoUrRIlRFtrMv02Kotl20RpDYgNsaB/FxBgKTmS94OI6LZvj/Eh
aH9LJbfemzjcLHvjK5RbysKOytvbQWKN2pVZVUiAqOZNZ1FjuwximHnN+tS+7Td1kch96TzmEPro
e58+i6I4VxjMZ5PEUma2WjhOlCYey6Gc0sVkGKRmXHDkN/BP69ujaWjxnSdf/T4OCHbue9p5vCPw
Ya3WSfWn5C3PTId9Da38QptIhMyCFGA3GdSbE+2TbW7NhOqYjj/U9hmfGYywJ+DoGswT/8xPLj8S
nmYbcAulPbz+vggRSUXzNtLwISTlI9DoBFbBYhfX5vee7KiQ2NJpk6fhbLDCb22/hMEt80Vg0Omb
eqew1IcVEfGnZs0Ba2DE3qb45mLRBrMX7mJpy3zGtM8CjT9xFw1IMJeh3fiuIn/UbY4Hbkeb2pCS
9NDd2REbLQUWB2nLicz4OoBQG1JdqW6oI0P9lzwxLAjSJg7vsNeoONHdioVV/lKeYoSo2SQZmw33
zYfpdQMhL9hcErTQPZXYmZ5eIMhLlJfkfptOtS6/7AGy6Hef1JVR/HFU/WnvyE1IIOWINcO6gheF
3zEBCJCzZmtMb/B3merl9sh1rj68YydMBsk5zpjxO8ZK6rc5mslyxKU+mQqFsDfMrio5ogZScO/a
toTzBtSVsdLbuUOmJb8fyUiHX7h3nFbfMkby4qd/OvlQWqJgm1m6MSv9mpKjsXJItpUTr/Gve4Vn
MGimXz1T0NSxs4LMqO1+iElPJs7X9agjcO3s5sRwKxqBuL34sguKzSe4IPTdvbJdGkVTqY/8EHJ2
yA3xV9U0+wDprmKksosXwrXmwMA0M2wcxlijGGPvYuwlQCCSit8RThreBgNMMRDadXlQU+qVqI4i
pJxwHYtOqiBqyjCX7ts46GuRwfZI7Y6Ut09WIynLirb5Mc15CYsA8xhWX6D0/4JsUUxkAukw1Q3o
IV3zdlYnqKCodegnfVv9HNMSXzvw31BRrTmNYXcO7Tw2MB/xbGzAFDf506fy64V6qUMS8WfWRDzs
QmeJGWe316VTqG2zsnXce0XMlPBoJNZw4Qk8SXCEJjvsNoB1FVnBLHqzcJy11aBTTHe0MHnWPNGm
BWaDgE80AMXCEHksHTJmTTQBt+ki/V6nkMHtNCdPCuIphjBLHk/L4fraXkot/v9OhurDXw3NSyap
N15Kdeejqw88/zids2ZdGmiCtTN/PF33Cdjga4NknzkAgp2yv6vf72WTgbdmFjMrOfg/bdikOXIS
DWlihNkvMNcqPQ0RJzzZP0+qA9WPZfN5nzTfE0c57+H8pif1hBuzFWEEse8+k2hXg4GBIUBSoeVE
l7h8ef9XhNpTU/hEPGfW3KztAHPUryKLa/nQ6KXy696qDCtv/xvx0Rw+6L9dqQRlUSBYtNfSA4yT
amrmX4zLtxOi0MeAYtJ066/EEKE7/nK0ZMlVsSSpkjcfoM3heHCwHe6uy4Ovf11rBfqxPVGt0Gf/
jhG4+C3EiCKVNztbkeYE57rD8pkR2JB3fgQ25vh8IbB2tsdyO0UViPkCNX6tZjoYhxV2Se1B7h+r
r2XLwSawjHUJarD1Lavqf1Ku9OAF8ySkIgyOCnN5lPESyLCe875tn3bOS77hHRlVxIFHI5XpwYP3
omNZ6W93GlcU1/V+SzZxlNnI3BXAXWSyvfITxAxGfhNKGb2dEUP19vmijLa7Zx8BkZiI8zJd/0Ob
WeTx7ItmgIAnxD4H460/W3CcgssGiVhcGma1rxQ9hWbyJLLIas4dVyzobX7LspNCarjSMvlv5dDq
iVOJKLbTTCAWqYMowyO8AvZgxze1i6wOwgBLzG2qXzlI90PTlLazJ099rIqICWesXzlGSRIaq/WX
cQl83MtM2ONI/PNuiW1xWpLbIst5xN5j26ygiNr50s7RQq0Y8EDOrSfa1VlywFHYdvG40U5uzDnx
u7rxUZpnPlZM/xkSDz+VRwigST0ycink45f/GvRl1+9ymfXhP0wJQJ3AJR+tGqNWBO//i9KSJP/e
TiO1UUUfNLUuO8NmzgjQdA9TNV2THS7I3jb9VI9MpgpSCzoIO+jNbz435kkgcxJ3zs6xenhGZSmi
032OvtbcEcx8SU8aCzisHWS1rXekY3HxAaYN0SeF6gYeg+lrPmmIuYHtM+bjdgrn5juEjh2SZdiq
ge0HVaiMYihvdYe4ws2gVfuH65+csRwLF0ADzlebRYXg3K7ke5RcIsB7i1y4PeaDcf6OvCd5DP/j
zNB+X3GwMhzwtmUM4Os84Xbi24FrSzZ223lDNbSzdHzJsn/B2jw2B9MCKk6eZUjSBm4tr/z/mPMy
M1f8Im4w81ZJCJBLXS51kwEVKRFuSZJn1yVs46Reuwo0mlAV3ld4JVoPpuh7gFa9h4mOzRAR94m6
5PZ5qY0sZe96ByMoe2cGTKg2xPcndUxXpUjdgNeoWVLl4mMbXfcWK3wX2P3IkDUmWhNU0PUZvmY/
ZEMfAbEM5JYmG93W3i1sbsuEKpEDecVVjPh83iUMB7NENe/qdrrg98SRQFOZcZOVOLWvbklpbAVB
jxBO9TuAcKo7tBM/EjFitjXvIT0ev4iRfhKkLss0C07nSM3OvjCzjmTUEmdvSSpGZdjJAj82EqGQ
q7wJ396CIDxCxCLv71Rwstw+xjabBwCdu/0AU7ObLQmtI4xcdI3HDmfS8GLgyqy3yHK0V30dodug
c9vvJoU7T5UeTVv/2HjaM+6GUHhrxAHPyMsvv78a8H8oE7NOQ88Ym6Ukl9vOhP+o5HK3i3fyLSp8
rwT4bagsD1U5iGL6yLXNegGp3uwdzpYUVJsmBpBzwFM6YNDmr6oJu2UWVDmW/z13VJ6upBfkWB9U
ANQebpHFGI6zRpbEA1z6EVHbCOEovLANEuQnf9hS07LebuuULCWdMYuOgKCXFn2cRnXl3quirezI
t+eIm00rjJEhDbldr6Yqhs9qCwJSml8OwYpRtTxqg62UGXkI9n/jYmgpvf411NiO2wJ9KMlfVcsa
O3Asct+5xLEPEei5uebk3JsN/tA5Sgk54I8Hu1nkHMEItdzKfFpa2DFmcMWlag32i6rNMdEC0CB5
K1CdtnE/dKz6Kl/FgSLZiJPFV+GQxClivjFzQ52pBO2dtjRsicitQ9n6j7cdk/JLoKpUWb290WBW
EGGOpslXkFITJCfJhg4Kzy4DtOV9g+6DHyFPqwYyj7ebvg3e4wWmzf3eWpUlMrkkU0rQiodk0UkZ
9G8nnkD+mf25V50wnzmreqIoY/pqextWGvJs1ILt+g2JFAUvFYYImuy7mSi+hpo7baiVtoAhtHlC
8TdAScZ47dTO2OozC4YHCseCtYZklIkJ//JU1NLoQnffctjlV1pv0W3iN03zYq6ONx8c/boC3FoN
MfKmYxB8CYYD2pBmC3FYiyiG7g3E3i+dnYfG3Dp8MosdlJ8nxDB7EK7TLvN+pclvtjGhX/57nCEZ
u0ld2Uqf+W93VDhBqbnv77bWwdcb2NSAGZabncM0VXkRhVC+c1k/IdFYvbt30JAOy4YI+1aJh0wb
R4EpCp1qaU0klxmp45mGeaEmnPZwaOWOKhh5YzPnu6YGe4PS3wOcWTutaRbWYdBEZzcPvYagnDge
utstqoNyJXm8bbxPSmNi3+vz55hjscGXPAPXXtSuhFClZb9dUQi5owD2+Sz8TsJrilZal9Ts7V2K
bT12Rksgtv1g3X46wQpjKEAS9FTehLFKeSr75/JTH8cbJJt8E/Zpl6cEviX1n74zUFFCnY3Rmjk8
yic2bmUxo4gXlGKgmIuPDOT19AxDMKPz6veKNyy/CvSKPWF7PfTrK/pHhZfSFMabkqd0xdGt0UED
+0kiJRRjE5UV14XgmdRn3u2w5zmZqNpTn0y4fkiEh98i9eMTHYSyqcNk0bi7VyHGlF9fJEnYahwh
7t5TSE4UNYxfj/38isyD48sWwH6w7dkfDzfyr4RdFUJx23PnFcf314r2nGqfVLo0ErPUg+yOfIhz
VW56xSmJKC9E0R5CwL6rOQGhUNJrrDoJD2I9eheOMlwaJqWvLgGo7SPCAYKgj2BPf2MVMdGUPcHY
wtHhSRPIlE6nXoV1D7T7osNKitu62AqC83wnRr+fp8Ugbgfe+q9l7QsmjkcXAVZJ0nRa2Zx8aURC
lFmD+K7pfe+HOeohQ8cf67DMKUKNeZjpTdh6AufZ1bj+OCy4ufg9n7pAJbYKO+t9O0/CKee5+n+O
lic5amBTyFaQoP6p6JIo7wa333NRRrp01xHTjPhSSaeRw8ye+tTaAZDiclI5drTlVgKR0QAhseAG
11GlnYmYsA1NvCGDZdt5srYkKEMwfFdsR5iNwiTvu2Nu9FEcjxoGt/KUDTtM38tj4HKwS4o2uR5h
1GdFNtd5uFiXa12Vz6Ya5yCbrFByCLZSfOiSnzZoWpQwKxMORNTb+RIOoJV3ok12j5+msR2MVD7r
smjvGIs6M0YCAozuccKQEy/oH79R729xLabaf8jXHlimYxy+Pa6BVW0+w0ppZ8UBUQY7jUKBQ5YN
PNp2U/YfvuWD0bLzXkeHnI4QelSclom6gXPYRSF3fB0qgpnsPTiNmvwdS6+ASr+mQl/x4fQk8oey
MahVkPaZjwIROvWPmMw8gZ61lp/uuyB+vVxBIj/pFaA/3k6BBxVsW+XIVCjld2urGa9FCmjh2Q0d
rVv6sHbRepaBUOrJPtbkLFZtYwsd67RvsMDoukHPaeIqo2L6uqIB4hLJImzaN2JW58+3Bsn1ahJz
tkx2Lx5wpCnFsuHKOCba7sDFc6s9LZVbKMX4GhO5u/37K8691LNvyPQqxfI9rqMtqnwUTUVA+opx
E2qhYYU4qYzEmiu2YCBKVL7UnAw61jJdpfKcNnP1qDOXoptjVylgWIV319AqB6jWgc8wiflBD4Eq
9QWjJQu9qeDw5BKEErXzV6Ztuy4q+ohNqsjUN21CZDKI3uj3qwmKzMZvB3Yr0SbmoiKQk7I/W5wv
7uMo9ftqXia2lNW+5Cdzb8t7OONEg7nsgUSBTRchON+hpCEAT2diY84sKJdfejQrJKEe42lfNR+3
nzIsKXOUIsqIVeso+eFkjOYEF3Hxc/Vfg6OHRwghHWWDxWaYdqKLMburkrPuUQunUNU2bGH41uag
wXJXyoJmfsmq1c8sfxdGcthXzLSyPod/Xp5iZNu6oi7kg9PB4tvjT8qghlZ06oST3iDK+aM9fo9n
K75C6JjSrbyL0sp6GbZjkxFkA7uPkad10L/aLg670tRJ+lDtiQYC8EEBoAA/zdkAgwbkBPe7Ag/S
x7ApZnIQEG6OVer7pwx5vbt8kZUOMq5Z6rjyYdNlCFXB+BhxrCr4qqQt5RlzGgp7KMp6GwBDmXqZ
V67QlLP0Rf6oSfx1PSTzR63xfRQL1GsYH+5vsOGdEXkmnakcevLWrRkGMwgOel3YGRr4UFw1XJ7T
J0nJl1kYOFk6lTyHvFEnLmeU+fEiFHturTAOXIfrdqTXzzUJ01SXofIj9eeMjexQWTJr00I7Qn7X
Uju5i5bn6H6wDrGpO+zrXddNAAJs5mwCldZa8RC6CHw/npURJXXdWvpms+FzRfSUXarAXrtDrbuh
9X4GhZPPiBAh8F9brElZ4mPV75N270SuotnA/iaWlemWm2jEKwMHKx1wGM0fnIEUpfpg53LIMwD+
qH12niV9+MYHMfyBNHIawB1HHgxaFEv8jSJJUxlwhNfaEvKGIn1oJpWj7BpaTvliWSFK2u2J3BWZ
OOguL6GgXjz9f/DKThlZZMyeVe5HSSRnSoZP8dm1FtSKucQqa3ErLtbh7AzJR23ZzRAb2LkArEmj
3Kj21E00DNtbCZjlP3DVLJy9PHifZUZyD+FnnKIMGfwvzNx7TpEz7GeX3rpnGtDa5O4wlOcgoamb
oFEeNMYW7MEXywcQUuo7QcK1mpsYoVWh9KRJeSH6KxSelIzKeMxOXoJmtHLaMMwWRFofZ8KGQU2r
3OSmu8uwbe8ep+1OPCMeayUK0JekFRH9tigw/L3TANX8sRLfDc2HCMmIx8XGY8URz4sy0R+TBKg9
VIRCuENscqlxb96J6oh2bPMKjUYes3cbOVi6oWxwsc0FtmlB2f55rqmVZhZMbPSckPbzQnqosx8f
9z3SgexspiUyUT8ikJ3iCSliPySW5f3WrpYbY8fJPxn09X6Aez9YunRgHaf0yDl22xgbOL2CQ5mr
HVUqLXPcd0uJ8ksBX3iI74il9FLLbUmoeHzIa6aMrvmcKCCNYSFDL9a171+lS3iaWa/5Lwt3d76T
dsVfc0Utx9n5/neSjTtR7+1wKYzP3BessCVmawxcooEUjBmyPkN3iQd8NqqwMgcVzpX/vCDoM13r
JTpHaTHQfZP/PbZ0jIZed8R5Td/tolQXjkdRfv609wWIxCEXliST2cq5Ai/N9Gq2fYRTLTNMbIod
yQuh2t70qhTE8dtUSUvDzW8A0ByRGFzvqcHBhp1okq3cXPNglOYdMpCbTSmSqiPSuAqAyKnfHTvi
JP9O/xNuadwE88JTiBaYMo8maytb8mW7b2P1WOM3jwhcte3c+258YCSMmjRFn2wiki8fKvbDSrm4
kSu41/SKt3ecB6ByrZB3YlxuNyvwkbJEukthfS+OfTrB6eSU6PS2VI1c1iO4T20aUi43HuA4P6KO
TlCiW+NqNEUuGXtXMeXqbc+fRKWxTA2MwIPkdRQJxLCqGseLwguS8hyuYAYIvOz+BLehNYoyKdt7
BlUjkOtEfnXm18MwRUPE7mvSdT23d/iIlTnp3CQATuiXrgDZdjlSbij8gtAiYsf26DQP7R5tqMqv
YYaH5OizIGUHtIC3gabPrL+jzy9UHupQU4khXlKZdAbsQWTRZIyzpumSRH44J57yVWjRzElW1Pay
i5SqzPLcDtq/guNt135ZLym3kEYSOOXTW6g9YJc+GuNdfD7bG6kAMk2caPDRRkdX0FskF9Yuukgb
3NWQ5qjz1rX3jCwSMj4Ck8mm5XOx3QYeJDeldO9pvXSRToiyK58buXVqk1KDbd/VOLBq2PJu+6kC
J/TL933rQfGN3Be2iqUEz3CD/QhOy1HpcoMsDJgI/0aXKGG3NhZWHfQRyg5DM5CeDt7PME+YILkS
63B7b94Kp0ElRNhlESkx0xugREfYOqMC45vKvDTZVTIDfs5+FLeF2pVJzw+3AmllPiz0VmvIFS7a
O+uM3CUZNPqiNpEOjiNFMT3ndphHAIRICmHX09xWVg/wZZGnFHCL/b/Qeg/zxUl5QM31Wf8CpQMS
UgcZHzHWPCM99zHjWpJ0qhI1/ew0GdvsNJW7e6bN7PePf2nKCioN9IwNu8jbs/QeQjLvMWZ1rRjt
isXuYByDAEnztWisdJlUw3seYyQyThLVOsqm4pezucs9htFDHCHWlC4q1S5de5rLML7wKtlWrOC8
ZTCVY6H38yhT0IVMH5ycwJK1KnoERsvGZqWYwWQEZUK3bMzsKK6e1M+9Xu0VqsrQonz/n4LPFLL+
+LP3piliQlZwSPnrNMfvPb/SVsNPiFTK+4REf8CxG4HH2p0pF+Md9IBXoi9OVFv2c08w1MVN4xuH
GAZYZSOzFcH7hftwPKKOHgOmxYJlWi0G3tH3s1o9Gfjpmi4tPBMFzVlDykLo6SmgI1u/AbBJwaWY
6m12FhEMeTTaYXZleSCDEpkcUITCEsDaVbYctThbEJU4o8exQ+2HFWHA/dlR/qWWb15sPJoWWUnR
iW6uEzoLkNf/1c5K2B/f+30SbcmVtneS7mTX7G+3kYcivBT9EU3f6eXolhwfFyyOPe2Z36Idlcbf
5IFZFLPKm/yq5E5z9QjVi5q7WKyS6TR3S0ACWob/v+ALBcuvJMDrLAbQE08F2y4FAVjF2vKWGv1+
MQ5hwRVbRa2x/Yif/jiONfmx8fC1EaqP1PS/A3ynusK/c/Psfvsc2ofEgC4eIh797AyNezIIYGxv
L6xD49EbN9jaO8bVSn+jwLMY3zEiLe1AT03fhCK9dSQDxA3A9y8lYIrPmLue+l4FhJZW8BUUll0U
AxKbPf069qhOgjO2zdxMM4DDZBKvyX/eXKeH8P5MLsnfk8Cr+ib2jgBfpaAzA+6MvNwfctkeHTQF
vC3DTk3riUZQT6b4R7OY0Mt5p2BiB3JBPcn8jsbJuq3e2JYafR4NashlaKX39w5bcMtaT+o0SUgm
3+rkJxSYIbWAWCSPFZ1fth41Nb0ff7xhEv0wf/x9l2Jqe/1r51XrWedwrfqWCw4uNDfz+IIzBPy/
pqHIj7WReGOisCWui+8PPv2Q6PQVLTiJiFpSZG7PCr0Px3C8V1FY2n9a7yPePO1btjzUZ+dy9IxR
xYpLyqoJ2M5ILfhRsEoYlb0lEjU3vDXxK/81I0gzqrixFyleJkRXnCKc9w0E9FQrKH/ds/3zP4jw
IoVS7jaFaMsF45jGxD4usAE4YCXpHoH8sGXPzSHyVThe7m2KybjtfZCdXp6PIf7ULPZASZLZd9jZ
nL/Xr0/vSGi9DaQ8Jlqq+P1r/Q5LJCzzbM3Z0cEzqFuOLQpItzh2fNY5or8b9Z0aT3vUBTBnTSCb
S5FDlzZORabb+7pp7+AVIpR9Jt2EYQE6/MRM8xzmqBUgU4UcgnpT5VzormsyOvLtrDQhZChnk5xU
lTnZwqzUz41KrqxyNZo24jj4F2dgp6w1B9TmMCWv3LpEjz4LuSbFOhuBqAsUdkJJ2DM96ZfWTCuA
5F6EWBjnwfCRixmvl4RECvB62J0VXj2HR5Y0lzinHxdkSGD9dPxGUbTG4LIlkll5KsR1LjiJzJFT
bd4R7w9IwTZM45b7Nrr9aEwgKkmtXhm+Rz41a3dxOH0jojIKmnmjK3zoe7qyaTBT1ukwyiH6Ug/H
i19uWvX3ujcpyBal3HMs/x3QtBmUqtZ+P56vz0GBrt8r8TFnCFi76OPQTtTIk3pyudZlfNhyjEqb
3ddK0cRQk63byPE+VXFFbXaOsGdnPc0yF/e9GCszamO61As3KTTbsV6Uph67jjyhD1xdbZ0mOG6l
RtiUhz2R3+r+ozrrr2dOrQo5yDNEPUqonyRBzFgbKTlQyenI9obX3OJhVXt9QlnCeTK4yYkUG240
FenaWiSiCggh1oDDozxByS00V0kFtlKBqDlAXIS7o8u6gwWoxlA9n7sSePHzOz67PVELJxVGz0z2
mBcAMk8NbGzGg5NtvvNmsMONujTM5vaVFcUujk+PVlL5nMynSK4s+WR+WKdwbP6OoyvcyQ6RVrTQ
9tF0xLuU7H5uGOlrx0PAEBB3w5wQU6WjG9+pfZOIZ8r9fBboOoUbCfr48zRwHpacMiEixdzAtNyX
MPwscciuhWwDj8pu2ySvduk1DOmy+8WXnimFch1f1t/q+5bP/BzSM5XiQ7rrr50+bx9zG4x1u2Wi
5C+LlW9Vjo1o+TNCVQmotLBvoTzq1UW/uEO6b09f7Okk036e0cv7HRpmTHyWliKZURAEuoinyidH
mIEuKt8qBy8IvEcEsHOH95D3Tc03MkeoZEtdDYofh4h+4SSrnoqvm9nPYInwexVlLnd8XMY0ssox
sXtyfimpG8rSnp6jFyGd7tYNecZONW04qTS3VZV7Ys4AiQGKFPzixDf1OSmfy5SOJ1cFz3pf5wQs
EQ9WasI7D5BqMrDsIW1VduXXTh2YZpdPu3iYIMrasZz46mkEkaTzKl6+7Vwo/nkAyYuTtc+GLBO0
xplj2dzMJ1ci/EKr0CG67277rxmVchxABwuN2lGVI+sR7o5oo2abTAvivTP8rOmNLG0bnQob+qAR
sqyFl3KRu2xPe0+9oAcxHXV3Vi0Z+3h5chL0DshTA4KI2Evfa0dINp2fJU1eY68Yi4t2XwC2FhWY
4DE7Op9otK/mjvIQd9JrUlMTJ7VjC4ZGf5w4DXF/AQoyd5FupdmPFmWNJ2tqfJn1vkA+N6QzXGaB
FzWY+5UyJ5L5TN5fADlizt5mQrgSa+F23WDNuR/7eYPFkOYeZkDHzkhPugS8fXLd+bbwlQFFKKIq
CNNnvtLTTJwXLLFv04dgAzR2R0y2gNlkLGrK0AUYJIE/A3f8i7ewq40U0kXb4DplkxMAj6Asfw/Y
nGMCCEcgj0HlTAJAz2P03e7+vjtBHN+zraCh53X3ElIam6pZ4WxCgMJnm9XvOFoHcgJVZYBD28MK
ocYeQ3A2xsQaHMuads1RxRliNDo4W8Dvv1hEImJgNx3SK/CSCF8vDhy29ZfZDy3VIXqn5Por6fae
mRy7wKlhTPQgCdSniDWNVNG7oZ5LHNBDwrQbR1upiW7BgMn6m+uYkt4hmNlxmYmn6PMYtV4+IQDC
tRWxYfK4Wvn60Hyo3O8aTF+md2pt3c0tvIBdt0djr1LuNRykuNsGFw2BovHpiBoufoXetvGKmKT9
uMdGo+HGCLOoQ3DvVigEvfHz3/PghMkrSGhmUMeHiiMeiP8KUDyF78Axf4jOS/M2gsXYQ/68O3Qs
EdQ0VfTT/c77aASRuzMndPFd2nFVvUH1Jw8MoDA/jyC1o3PmL0irk+/gFC+Ppp98eOHY86QrvOmG
HUnRMY2HglJo+R7krFDFLVNTQeDM5zJM6BHOnq2SYPbxsZyfW0w3VU37wpWqhfBS9oC8BlYPnvtg
Cia5eDQQrCeJ6ZpZiL6HlJdtSoocnIqzZLhV2KjGWPYOE8IHyN3+VrguYkjTayDYwcEc8Am4f9Od
O7lqr5Ixb2zrPmsBhRK0zLitg8u+oCI3vOVbHM+2zqn16AFdmeuPSQYOr2F9xXwHKZXzkmVA0q+k
yMST5eSAkkH38gc0DBhpgPzCfrIioDTbrvT3MK6Dd5s1FHc/tbD8uspXgbo6RrYoQiYtr0WwF3vR
yv3hGItzeuajwyOhd98xGFKRHI+JdbdKcMfAT0WDolZI/Y47hoefukYPdLK0ppPNSgbSZ2cnW3VC
WBw1ul0Pi+Nqu+iZ6r1rwa3Wy5WLiPQz6Td6IJRG5ZWBuHLav0/9q0pu0ITF6g7STkDUAOrqhxIL
pIW5C/USd8gwJUKPs3EH/PbvIhP6tJT58CdzvQpwwrV79keQORtxVlE9NCmyM0s8/lLD15vJbr/2
9IQwicCsWS5P/XhdGGJ2+nrEegf168fVPaEBBbnljdQKdK28h60TfDc/LWfdaPfbzrfTKJJ4YVvj
NdTKB3zSaBX89imguuBMFOBNC1MLNenJ/E0qm9Cx5bGsoonZ69e0pqkRpcx3cAe4oW5lQCyZ++Qg
U0suPyricl/r/82svCtiVMy+KZsEPvAZlGbrZUHhBjvLyllFMB4fv/yghXH33KvmmMPUE+Ycab3i
2sh5asCStuo8wKxqBhwaiyEwE/qbLpmB6o+Dn/SDUq+5t8d/DEZgfh1CifxRxkbP1TwZPs9yoM3h
6Zb3RQCp4fzH5WxJ3aLLrCOGwUXPZ+XQXAYbgcKHyhqVHygdv1SqpP8PC3TJg7B3T7FPjw8EVv+P
15H2DcTp/c5Uf7zbL0d0YOglftLhiO0gIiF83ZesgGXueE6McSq8oUaYpM5vuCyD6wGxYSE+poHh
iAPeRZT4fu8ir9vvSqavHjgiIUsQPXep3T27utwnWuzl/Telo6heYO1u29xyJ3fgus1vqKCqapRH
pkcob6qXQgpiiCwnufwIma9QLbAYC2d92c35hmbFSBek7iia9Cuq4s800vdeQ+UnHKte1hAXV4OS
e2pP1tsiYjhF/nd3VydHzJl7LeggDXIImX0eFSAXFVMNvqiVtKwRuDPXso3+0V+v+wFZflx27DHP
s0MkreYyZOJtdgqCKs1+q5rE58I+WR4VGKaY4lpZcgIOt3rCjn9wgt2eO63ejlWra0lWzVNIfng7
5QH+7ZUxP0bfsmQT2eSEQY0uL4jqmLLFj9BEMuBq0hJzvDn4XE+DPAv+8yAHUWysTQxEQ6vBpbVe
vWoXnqT01ABrc4G+2lC98v/IWWrKwLahbfHhG8Ax259ZxXf0iyLdxVBpXzAGfmtXyrfU1NHauxi5
lD315Kv2jJu0KipnDDqywHTV5GkfqcVc17CwC03aaQbt6y0HvXQBKe3K/eoDg437KH5AVYSLTfyN
82WbVXzLCOF5j7O9ag552r9V8dJILoSyIGMLDIpde+u0w9hqX0UMra2tcHi/EqW+4hol1vFXUsdZ
aDQW60UPDvgeGWQgFKLi85I18PwX6d4OR8oq9sxtZcTMBBx2JCmUNqaJMn3IlQnx7/c5uYTOw0wi
SjtYH+9hMksTQd1MHG2Gb9pfzfn5dUjlFTa2rQ1KcKj8R5Vivsrc7WW8w7FMdjBPMgDznPwJZn43
spLA7JY6TPR/Pyum+oKsxbAGTNJkgcJpIxQWrjNFoL6cZ9StLs6nw5FOSmCmlazAc1iJgMUKYF7+
un+MJPJBE8q7FVdet5Dt1JZAuiSN+BwynnVNClVNogrvYvPzpJQQxBjR8OyvPau7jpmPKDPhFYlH
/yhTXPs0E+U1MG81N6Xxk/zxsRMrFnT6LNvGNr0OJTWMDWYc5iN5PEJQkRNyfoYdSLhhpKP2ofwZ
eUG7gpefww9Wtb/BrzU85DC4/iL1hhYNpzs5uaVzyE0q5o8wPXNX6W1822Zc8Yp+t0WafJ7DOFg0
TsmYLXfNgPgt2U7W/RPIeNTvMFspW4ErKthHPQHXVFvRzAN0O6XK6/mpP6bRX7y8WA6F5uEuuY4d
cMGShao46qxjudj1dfZJSIa3fmthaYUJTU2mdef9Xn9AO95AOpdmJKI/jcwnudf3vArImGDaUrCG
50rFqOpZt7FJRVKKIVHEnJgVYQQxHeaoCWGGnMg0bHxPjBZhkbZDF4WC6sGm0dBzFd1bCFZyUZCQ
xfDfaS7xHdHsD+i1DCekHGi5QuynEDuE7w71dFuCG+C9qSakkSAudxFV9LSUmDMa2tpyR4d/ZigX
sipd99UvRWsoMBbWQvevw6r88xNjRYAHk2PZZm4Unn8toGI9TriV82X7j5jQr9Wrrv0mtMaBeKm0
iDGwnybf2/1VssCqHUQA+Ca2Pw3+b0pI3suyXcnHiaExK+Hh0lj/Hs2sfBVQmesFQ3oWzQs9HRUR
b9YvfI0sI13dyzY/ggCNRbcp0FRgf9qa6xpvM+7zJ13MaUryqVHALiG82OwqYgM7w8Z6FkXRiqRH
9flya+jRWJMALJV/+y1X/q7NXoIbcd4qVcwVLiZ4vP/BGOzohiJQJ5EoBqRm95w1T4ua/FC7r2eR
IFph3YyQHz6Ku4jf6ytEFbpTjbiZ2d6UpZNzsDjJx4hfXpY5IpVO2D2zFasQfTAm/z8b0QXrbWIf
LmU+4SHAEfIgXXlhEL0XrygBAvD1dn0ka7qthDJ9IhrTG2eqxqlrd3/jHrVJIyC8/ZSpCS5YCMWc
onpFjtpF/qTqGUR9CWqBaEcA1ugyb8REUd+9Xx4EYSvW2poucO+dOrwgDgp7VtszJU8GkHg6h2cG
mICw5TpBKWKaQ2UNeOPmLkMsG8aFZDgubH+1HoDgNyPxGhoWn4FYW51NHMagcGm9lrBxi5vBhMUX
eGA0Qwx3b+dxEQmUZBO1FNCtOTYsypimaE75sp4h0mwKeGPmH1w7x9O8b909/Ht6Mkiu3zeAEJgL
aC5s8bx83ikdHdzf1AD8lWPfcM04OiEGUhlcnNWuskEF/NvwRcrkbDl/ulRqoucuCGtdQxI4m8mm
5t4N2LXbrBNQ2CZMJVj4C9caPzi8nWExk6r7KErLY7xyH2adMdxAkx8eMuFnfxFVQmifXZwkDOXt
mbTt1uGHvFBjfHaf+LcRSfNE6k/W5CIqMIFdy9wy84QPOxFIdSchUpTDJXOQuZXtlIOJsfKtSBCU
NddUmySMjf2hzin8sushA6GcJaeaChEu0fAPkIwEZgZXJt+5eS8X1sFdqIYf3lrzWmexkKM/Ft9f
41rZ/YRdAnCJBkq+b7r47TjMuLF60isYeo+BbZ/myzyq4mIVPF5mQdJDgCKtVNOzgn6MPVAs0FSp
gMb9tIv4sN/bcma/A1lEwInUrR6Vb8+ppox9ugwO/PA37895plO7GTzxWVhwhIjPxDggOWUyD/0N
VCESwK/9dDvBXJz+/EQL8pB9ZBdH6qV+fVXx7QBz4uDFE7/sAF/2FWNwsBvFZr3umM82BYBQtLTO
LV2LTMHUPAxdR4BM1hbwg++zAzHMRIAkaIIEXhHJAME5W8y/5qhJWYgj3B6aufjAYHDMQ7eP04/d
VCYphP2EjL9qwvWea3ZgN3zvpgo2LFqUoFkS+NVflVO/tRi3HcrNVvzjRt9PGF29Rrqr1FGa/tSk
ru07h8TlPpTz40g+4z8mCu3/9OKsrdOHn0crvPRtXVcTEeK9oPFvViybWqZdD11Jk3jbIBVWfIZv
ff9el/v3dhrnkSONxAOGoafHRSbYNzoWN9j6RqSZjhbQXr1UEdA/yEn3VahZib9uXhLQVZzj8ZCZ
2Mf3Y1IjoN1q464ba91QQCAndpX3c/KQ9ZmxZ4uubRlNtnTqg7TN2DxjOeA6M11ArbyNT8r66OEq
wPBzdgFDEyny8ROZGlMjG2de48n24PHqHx6d6ZdRmZJ5mOzw31g5k20WTZK21mD7wJT1r+yX9paX
rc9/InKiCJEWxYM4priXbSTqG+cMHjD29KiNAIsohR0yuYDCqpa9zC4SL+t/Krc13nYnPrXubL5h
h/989BUvUCLlbg+j3rQiN4cBmYeZUF0Q/RQmXq+LRTEhPlYyUncu96QP4qUDtA22ml8lmG7qwgbc
1/0SaW/OSwrA3Fh1XQCBUorcWisfDtJkUhbfpul/4rRaVxjaIXXqN9fS57hOwESoulnLEVERi6OA
On7WgLV07AQplmNVuTm7XLMf+KqidxWZSptSFcExwH1n5oYvV2mAOzMP8DwV+WAWrEUkals0pjio
m7fKm/Pjl1NgYC1iCp7EHAQ3RItcZw8bwjLI3Wf/fYLcN4X7TxJ1T4zS+j0TIKb3cbO3xiJ//LWg
5ZLt3h7xeUHXKO2LkN4hjYPN24EK4WBQuiSrYfk74IdHXybVV+rC6I2EoeVnXNRy5TgWH213wPH2
ev0gDKIWFGTJaisQIPMnqSVmH7XmKFwn39UvILCmTi/lDFfcti0cYsG6Z9x6IreMMlEG8vxnNMPc
NpMU3yci6YPFLLDQYQfmUEaedJtQTIyfGCFkosLjUbvHBiXkYMMZz6rhzdi2x6gK1ah6Ixd3gfm6
yydlTswWfRPzjk3DhsdemWwOFhq4TeMxJPtKZ+LUg1FrifGNCIztp8ESr+IATBFo/D1ZSL40UjBr
rfQXPWckLaeg62VCqbR4MgTM50pI8ewW46gl0NhBomDp5f7mLjdJ0wewqbOI714O4xx17ciGqaPV
MjE45L4McbYpVWsYx84P04GDeVZwVoY2mABWQFRj9r1rqDRn4/UE8UqVCYHOAVcFMRrlM+EHJF4m
0sxJlXe0EMhqLoXte5QyX5W+kRCsVvyRfj/uNp6DaGKvW5Ysi4UnWOoHaQ6BeAxGD6xd+sJj+Sje
0Brw4LccVanYYugHJKI5mQhA2I9q6U3UBLz87OroBWvWwXb61U6SRa+ZDmtYsew4QljJ4aR5HlC4
dhuXmKPepimvXgadfNRMp8WnGwDGzqvUbCS69EXwxgNnyQhhZeJ3NQL7kHMQGhshKdwadgW1aG/4
5uHxbn3K9h+ZPZVMznmNUln9ikRmm1/SAJNPvO14cU40SbnhUlX7b+nDEU1VZramN61KLc26F4y9
6hzWqfAwhChwnF4okvKI/Xy6lS6FpFwbIKO4FcwNRCl/tfEs6TOOnaTm5rDaxH9pkssDRuZrubVV
GrpGfgqWE1VVgeycrmTJS6eOyutR/967Dp03m9iuToERn/1ZGcxSgLw5/GfsHYvCenytoExodANp
tKArOMx++ayOBUDhur//hi3RtLdIRGU8xIk7Cizx6mN2YNVdWmeg4j/ciq7ReOkIr4DF9sRqR9cQ
WF9FOMQ+Hk12m6MydgqWDb++FGTEskiF0G5ooWnG82y2fjvdvzUBrE8QlcuYJSr/Xia//7XMClqt
Dn4YZ/6TcXX/UWZ5ng5ZviwWiSBlewWM6qCTm9ILyKJs5W2ZVBwrcKGgI3eGPKXVo79a1oAhHL72
53urLB07FQlEOqr5uR8aLrwVFebtBZ5knC30VthNobkTfqlWPwnQpFyQw5nIWvql2RigPW4qLGOE
jOTXsKBECX8mUnx80pKHy1CmrHgN6TM3siGqMo1/P1k09N2wG+c9yVC/CBCjy3CYYHZfc7fRzrjr
eBDCkTSblJ5y5vofhBh5BlOgiCbdipO0YKjhzr3XJxlVlLIhoc4vvlqzXVBTHoWO/4729uknJPM1
8zmI9IQuPUJDPNE5hcoRzchzud2lPImU0OJ9Vf2z2IfA/ukaMuc1tQ7q0JdnH05kWcI7P4OC8vUQ
UkE+bHpbv9DoYtdhxZHYSc521Yj+ygNtvIzrhrfe78rHJttPMpeUnf6yqNfCI495a7gRen6UboKx
Yao+zbZKHcwVpyLDvcwvHfL/7hFiRgCH7WrBtgIljyLh5AIYSbbLvWn8KhifbUUgSqN1+5cmzSeH
MlTIlEu+1iWXSc/Ag9DTzU8brLKbwYHXDB4MhlOrDU66pV7PHX0OS8H8losx1Svp7f2ArqXbtShN
bPFTH2+0UTRpSn8FD+jExKBv8iOymI1XAW0u40qKwUYAsaWF/u4+t6WQp0LSzk/VVD7xxBRNrH88
T+R6Kbod17Pnk9MxNcTPxVKOUJwTUfBJNinRWkJCAilCo4XlMBrdqWx9UgQ9JhV41JBpIiHCYx03
vhlgjl0eCzZO38H907NZbKla887NyyuId2DbNAtOTAi705fw414PWqjLgIAU7unFLyvfCHudh6+F
pmVXm51jiGQmiYMiO2FAhjO32LWxwGWkzfigP4TyaoDr12yD6NNAgmQPCB4x4j17wGcK3Ahnx+xi
ScT+9fCQJSxoKOeL4Mx6xdpaiSbk8xlcSir+TChfkl2Jx78quHHkCarzYQPOHx2R+jnnYQgn45cv
EGO8+KoOfgWyvb/2H6ADdLGq8nwjVCBAWffmBdWqCnA0bwGmUPIUEmTrVmWd0TWGNHbfX4ntkVXU
Q0zm4Oie/oQB7Z+QcgQuoBL+9FFFkMALHa+AFOmvU+L61dKKvlXvnvINEkzu2b+WeXQ4LEKqLmPx
vwCoCeLIuwOm3y+F7jqCaJxs2YSX9sKgCPVJHABlMijyCsppS1cIhVvaQsnmd8jO3udI1w9sxlcA
T7m7qqrJ3qUKqsQWYqMk7GEdasOyE1Np0F071Qc6M+3is5zK6ayvKIIGJm/aAiojbZyg7pbeJYpT
WFUwNCTJMWYfIxf2/JIqH7cyjqSUYsPna7LjaGAIfAk364G4w05bfnEDG/x0CZLgZ+cMC1NN5B1G
HAjwGeyi/8+fdmEprJ3SIMoPMTpRCTaJhY9qvVjxg1NPN0xPpeXM8/5JogApo8hnvakkFRCypgSL
5tj4L0FiuOcbVn+LcL5OVs7x6WBfn054w+vO95Fv/paw9ul0BLiZlMOXv/afl8ug4/qv4tF2GUVN
cm1T7L5PZvatDUwqJ6Zr4Ihr9MZzeDC1DMEWUo8A2dIZeSGv8my6l+a/R9T5UZOV/3bscfYPohZf
4enqEVkZ4v5fgDDb09t8z5+yomzV81nt70ppBMGz5a6U2L9X3N1AurBRQRWV42HkAKRixWcRIqMv
mko5QD/jQpYFpdk953E+bTgrSs08XFRLOatKW9kI8fLLU/qxlb8nuANtOrotzQ9dLWW/HbLf1vZd
SirTgjPQbbqKL83i+eraPORWGpnRJK5aJ9CGwef+79imHJJUPy4VOl/npug8oAoA+xdezAQRxqCG
KVRmqZ7tOZ8xCyOkIZYKVUkx+CXfb7enrio8BJALvOoM6I7kJuuP5XSE1r5psK58XeyPZqswlJJX
cvlr/bcKSxmeJeYGg3kd9U9ilDYCSTQoH/RmodQUjkiCDcwjtlNAXBhuI/V+wpOzFMKAD31xp25n
b47Qfa2eeOfpV1knKU5d9F+w6XbGGympih/BbDVR+uSc4304UAXk1RJn9rUfGMG4hbnMmelvQ7bN
8PtuLWIaZ1hB52+odpetogiryfAfvFh4sTbkx62Lz9QZEyBqVpW2t4lvr+NoLZju5cwCU1DH1IHl
u1cOzDerbdkviMZeqAAdOSK4ICWbTZnHSNl3jBxuQ00/wrmtl1Xa2rgIIerNp/eOxISDn8QnMwHs
qg2YvYkn5zcu49HR8Y0yt7Q0TLpxAn40MFzxDuj+Hi6SwjtRwOWqY/mMzmrSSshXdQhjNhDPzUY6
rVfu1F/9O81ZPO62C9e9ph54bgGlB1DWlriFtmJ11CVhQ8q+zPhkGB9cAWhjWFVai0O5l0hJEEbf
Woxe/8+AJgCzeLo4hyrKhIXqmXBAtDjC4fiOQ1bL/GxDjRM0RAAp1z7Buh0OSH9BP1jZCrBX/KXS
jyrzJcDzFM4BoKlBzFl8EI/jVuUH63zi9DBH+kvrAR6gyKiRSx8ilZqium6uWEJCkNA77O35kk+/
FtZvWl8Ya8ICIgqkLESW1B4O1hGTFlopMcj6QCs/xhJh0RntMw8zChQ9HgmWDIfTvWSk0oieLJpt
D5ikJFKCc1pOMdH5ol+n+ocyL9zgNIeSPmx/jbvtmLrAv41T66d5vljyJpYk2IiI7nSKoxe/tL3f
q8EvlSJ1iaimKS8rEhFSjVV9H3XR/vJob7NtsqHNic7A0bxAtVBfHSqmKAcM87NUcNtTuq5C3uJ+
9NkK0MAlkP0eFTfg51rCxYp9TKsvMsM+lgA+DETGeoYKzzxutp3ABal7Okr3kUPRzDGwCCyo48Jw
GkZBbYnqhBLpO0fYs1s/IXGmHLC5BrBDk5iVepnyHzp5khGFCJPYTszbkzd2OtimOlOpcjUkn+n7
tgDj0XW50K8GEUIYg+Zw1ksBpG/Z43txzgjlydtkfhy64oLLe57gObiLQfiFkvUhFVPcJtANLuwD
tQDGG+XRN1k1XL5IMYb5X9h0GDiZfSJk6xtE20UAmdHXZ14CryYOcwIJJae+c6dHpivozemhiCr5
oMTGwFOcuWt/WWkUuaEJeIQtLPXtG1qwyHQbhVpoJDOGg0W+jOjlMaqs73Prup4AJ0s3fOwgCiBe
bTGvntDpi2mCmIC5TfEEbDJbDKFWljsmW1yMQS+zfoITc64XSts6ihVm49Cbho5RP2yTPmmNVNaL
nBdIBTaXpv2PGlks536lmo460whVEMyAjjsOpGKuNl5XbtUcW5XtR3JjfZ3MMNj7DNyK5FF2d80A
RV/oYpkTmBiwVGAxsL2wNQ6JinMhwdB42EKxVbGD7j2rEZgRyMl2XLQQpKNI9tlIY2eZwVPWL4ED
oHBRcD70WPTLJlU7AZiXSo40Y5Q5OgU2oaTuQ7V/IT1fm6Wfldmhhx2wf1q+5KKCGoD3IIAONDpI
awOD2E2VTgTt5/H8fGOyBg9LWGmcaRNVVPxJt7NqdcAozzhPlqVkMMLozdl2QJhvNZ6+mHEBPmdr
AReIlFG+tmlVzC7H+7SXprhPcMuRHcMkqJAHXUCIMY+E7zHh3myrEvwCwRb0bNpTJHzAOskwzofs
Hfz6XsYIrB299oBJ3AB2wkUXO79AfxKS6i2AWr28T6CXW2CG3Hkp6VjjNvdosRjxLbkKFQvAjoFT
OrmSP5AgUA/NCPShyyMPMZZ5Ds73FaPopBnJscDfFpFKpyTSX5KRvH6xOHX7XtgkegSdkjY2xDdH
9hd9+koOjOD4EC+Oe4rNSJjp3KI4tguRojK8g54kgvORrjU1FupIsIJD+A7Xebm9tRZkSL762+/u
xijt7pP6FKLB3ycpTWydb6shtHAhbzFOfxaC6LRRzLXWswciCzeAnhBtSXFDL0NtFXOtvpKHjm/N
fDsWQSO39GWQXvmlzfV6rcu7xWWvE8q7lySlwI62enctIqJouMehC4vl2JgRpi/8zbxEVjcuaW1c
uWWtRKjhZGc/V602amqSg5GjthkskAstQC9/tEjmiskNSaVPVRpXWO3UWgEP4dwCSorsF5G1jyPy
7+QbikY5ZQjok7BIVyGTjxBAS0UUa1y37dK0i9ib4PhYOY8NXn1yy3ZBdGsGQfpUeWAimYO7elaz
IDJPXqyXwjUnd6LlAGA2e/+owMmwNhVUlAnr5DRiJ/yZmyXnLYI3aU7umo6sjis4UDKBO+HWur1V
vALY5+ugE5smjQIiVK/K1UjBym/evKcv93UjkQGD/7HMHCf6jGTyi5YOVo2uKZUvmw2iw0K8Jse0
aEWvhRxm7pqpzUfFfZmPidjXxsXEkPlr1CvwgIZHCIdW2z6j1wngIhoZex6+RyRMyQDF61nab8dS
4yzKFwIwjDqn3oRJNAcMBL49bXvb7zShac/W2pD6dwako3OlndrVmFAAsftZ1qG6lCOpIHVjEmqJ
pcfHhTHz0HZ024IK3E+uexbBhcE+2/dZZj2yDlFT/y5g1AWfD3Gq3VJKVSYQg2EHCQBu3PTvLBo3
6RYU7XMlGafJFAkvGi97D2dD/B1QJaBubfS4hrmCn2zMuYogRaSNAwvOPcZ9z3/H2gfWGZa6g46B
18GdDmtU6LrRMcBTBlT8vzfsMkuHhScZmL8eSV5E0O3BvIR2+8Yz6LagHVTIWGPyDLHDFeifWZqu
6Safvy/qIiy7XhBr9c05lNl0dQfgIvulDCpgt6SiYo/NkixqR9IIgE5f5F+1bznGipnoBgBQMLow
I1k/b5xWFYRySTfyu1c2L+sJ8ZFBbT4pvFizgB/1Q0d22i2Z3KFPuWW1m2mqiN4f7i/KAX4dT5yp
bn5GDyQHq+xP5neICXt0GA555SpLL2Uj6rE+3RiObZDgDZsda3e4ds+oJpv+OIhHc2f+NBdGnD9L
VASqLLIHVVyvWr9j84OIHMUIRyOB6/GSo+NiySzdUvzWlPJi8g53KuCOn/9f9qmu4athdjxNHmI0
8uZvEPgoBd0zLAcFIGAvxJP+9hfPLVJ5Dm15ZkbmkBTR2W9fNtKAGIvaMYfkLo4fVgMtNJl+n235
U2Lruz2kBUWO9zYXzOsKoOi8TrsvDcAZY2ugkqC89u9OE6IArkdchRYjiW4FPyXd5oYs5tNQATcX
+NedElzgR0P0zF0bqeToJDMS9+eHJuqKqtm7vnxEOHo09oEnkhWEI8FdDBTW6SOsvm7G2SKzmcW0
jjBKnsb2HrjCZfpMuFYlAFGZ17pToNEnI2FA77PJi5eCV+If+EBXfXIWU8vj9BSEXvJGu5uaunF0
y2lsYU748kgEBHySZz+F0v/rOHZ4qpM3xA/Sco1fhglVJ8Zxeu3KEEQPxByAsguR9PH8rcicGsVt
1+wKDThVfhDkmf83T3PhMjaXZtKtz1F521XMEZAxbFaBTaxoA6VNL916XOUFfHohkgahkvycalpW
TTrB7FuudMCNf9r1XZynG5apac9reh7BV211OI4yDwdvPNJkO/qUhRg7TIaEYKNyBq0xRgPFGRzx
UbqJ02yLUEne/OmmE3QVxeA/nsnt7n8KEAlJb10JpNkzoxMa3KsgkmxJH34FYh3KGIpIHovmU4wg
jtseIWNeIxT8EOw6Xk/HkTkEvv/mkITO2CSQscly/LYjCxoZJ4F1ICgr3ZuKuhMxMT+ECvLtG1Db
yBRsGf07dUXSrUJdvm7Rb2IAMutnZg8leosqVwnTQ2pLiPgBKW6uoEL83mz6y+8/cGVJBv5VD58H
YcOQu2ArRJW9umCoo0rnIGIIFmjAwj23/jx58zz3A6XjQLboAOXBIvRmm0UGLyt9CNqjXjDJRsJr
eQArfrjjiBuXTrrxo7TQVrg0KHVXoIkcpj6YLH5MSqwpJxjNIhjG8lLf/IzIDS2JfhhgjoIMKdXU
mQi4ePW/NuX6ESQNUF9sZwD6Z0l6i7iwV13Rg4lawIdvl8W4zeL4Ap9wtmcV01FfkNbWx6M0QbJc
IYDrdR530KIMiMmGflVF6mTc+w7yk5qKz01xfxA9edsxkMZvofyeiWBwNuZ065nYuisEP9H+OT/D
9+q+meEZ3UL/ONltwJjhpMGPSzKYk3rm9IcX4NHhvPFrX/7IRrmf94/wmya+RsY5K4JyshASsP1z
lGsVKtMGhMqx/nyJJJw5OGJgBaZJ9ctmWrAacdJcVDClB7c/PYPX3unCYIcbqkhqKZWIcD3SFRSM
kFPWgWWOv9VSOn9pFvkYnsWTAi8nwRoi1zAN/UOuWeh4zwggdOywfFT2CnNl6wCR/kcWPUlGr0Hr
Vtveb/sJ73uqFSCTpALPWUWHYZBFU1owYAs2JHF/S5jzFUBWk6Vbn8B3YIdzz0pxosAzghCJOIlo
7/BJl5DtQ1qHpWgDDXHhZftDm4OD3ARb8kkqKGqksctge6sYdI5+prEqK76BKpdKVeq7ky8aPvUR
cJbPtoinPgQynoI0wCGPPV6wOi+d5FHOiXEqr309pD+5p+5UIopUCU9TNwVLBqDvEZ8WPzlDFL1q
vpRtRd6zCPzBhkEBZKzPLpdxXt36nkhoXtG2VrU0XdJtYeAt9fJY1TQWGhAwCNVFQ3q5KyCMw664
d9TuQNerW4Qz87oXHWOmd449uF8NdYcM9m/C/2huAoagexJdmfzTyzebL7N6PD+vwddcpwrfdXOV
fEKMLwhH72TgjcvJsRNzkTvzgnrpeXq+3ecpBmQEasiqP2inC+steUOd/AoOB/rVN7WolUJm0Iyt
/k8O0qW/UajnipJfpXiAL/0PO1n+SsyLW8+FpSFFj+AqjXtTRSy+m5mjEW+Py1gVLIovwZB9xtRc
AzMsf/uKaQbICcDr5av+OJVr7VrNdDPOGTXVeAjEOYlwH+WS8wi7hb1utUVplL9TNrU6N6A+8gaA
M1hMynYvkM4BsJyiVntgandWhaAOXZxjL+wGWMQVKBI+JkQiH0TnIKQiMgwTLUnwFZzQ8SPbMKd1
NmL4SKiW68sbqXXRxrBtHZB59cZ1EdVXTWKNiSpH7dGCX4sZsfObBrR60tbPDRRqRjZqvx1UlpiN
61Nc+9QMKrAeuBG7XxxlROAIg+dwkd2D6wtYB9dleuYDmT4GP9feUX0xIcHytcd+NcXHC3HSWizt
pLZLzbpCAH5vPLNw6EvUzGqZ1swrajQr32rrTLjM9a5FX7G2sKF/fOtFfjtinongpEI959sFoXe0
u5euSvcJnN2rN4G+45FK/cKwzECsy3vjOI1BBdG1PO3+xrG393lfYPXPAmdytZ9PxhaSkXZ40F/h
gqONIexcUHYY5Z2/GyqdPMxEBJRCIswbBntsVxVsZKLSl/z6bWczeWFEvFypFu41sbD7Dfc6KzPB
wS4IDqAjabZBL78XwUQu/5MoXNRTxX1ALohJPJ/9Jxjgo98SNXqWWXm7qPnQ7DLW1eMHnxksjJJg
/dyA/aqVlnChmXNjzToT+uVBXk3/V06U8yoOSspZx24YaDdfLOeWJfYNoUBMfSLK/OlX/c25t/GT
ycgOmIWEq1sqhOmR2Be7DMXUnl+6Q38Bekr79IJso21gRXfgM1Xk4Z30xj+dYJjf+Hvuk6+6spBY
622hbBrZq1Wg4cPvee2YD4D+YuVUBDIEECdHGxpdhUOM/NCwGoZMu/mE42h+/bZu8WdTpk9FJZkB
sg9Juilq/oZ4ucwrYnrLAPvgBa0MGcl6Cq8IUwJquEy63oc9VWT+bR/Nwsc2rtdLF1JdRN7ewPaT
zgoeqh/2tgsLdIffW7dkfRb+xv57w1vD+4JbwZO8z6V5999DynXUs4j8HETo2jromrGd/fUie4XK
PAjAN1TLbpXLCaWDTwzzCuZ7mNzfbDIje6MyXRd1Wps7+y/tvQpM/ckMSNkYdkMHwqChVQ6p/bbQ
u90X7tcC08vssi8u3N13jOunEknnyDTeRpkK0EED5PbevVwnFeu+g7bEFfOlUEBCmWwQoMOh4/sD
RwBG91iQu0bb+fubYscFEOaSNhG8kCkLhQMBp8N34OQYZc0n1NSsrvOGcNG8lU9r5gnHcwp2oF2E
4H5kxZ+CdK+/05TFLymXjwHPgEOAE5yveAtPYpy3sOSl1VobrE3MVohvn9h3h6eDWdSIYb7m74Gk
kviWWuiDaTJ709ghaTEdxET9Lv76CVcxttTjWs5TjC3bGeg5upn8u8ALkRU3pjlnHrnc3hkLmVdI
0VPaHFE3Dbq6dP/RkJlZh62dchbUKqtYSf+VLsuA99c1dp1yz/5A8YYr5GaDNb/uz2CEEdZ2k/lm
QgGWUL53N77vB4Fe8l8fbFV+Xpjxdh/opJbtK2G85vehnPLSNA5zMF2BihCCelPDkKaaeemmKY0X
4WA4FhCXsyc2KxR2utz8b9YQZtPcb9EF1R8RgunqglDMSBR8coX/GGxnpwccwY6fjsNMpt2P48Ln
/rp/UiWwOPIsx9uh2W4G01XEB7eB9j+XK/3sC8LOC/EHPZal77kKulefaJOofO/Uwjr3LAm2CFXO
RDf8thU3zhINdMG+pGycgcWIwLdNI8YGxcbwlT+DtpDzhmiec3XKkwnY65u1a9Ft7eI1sWIf6rNl
MZlEX8ijpQ1ZyXCQan2mUO5aXnGrRVEB1TEt2Ia1/ZLqBZQHjScmvMevDF1hIDY2sgcpd1+HfgFc
L7Rig3YD62Qq/Vmn0pXgVZDyBSN+QXWwBn3vns993cHU6Qas6nGY0nwJDuw1denB9f1F6vGIvolP
D82ARqUQMJFK22dzS5kFEvZb5AjRvghgQXVz3d1+wmnYFrFXBAXj2HrZwaGHvh4Eq4fMGgWUzBk3
WuEdaVxSK7XlzUD6QlMT2vYeW0Qm209SlehBR8l3Gquhb1GI0a9B70zMRTTUa4oXtbaiehVTPlzw
99MAhZfNUr4Jbfv4HCchMzA3T9qUyj4Z2nO4ga9AuWNfyQ0I57725+Dxd/ehvhVFsaWfahvW2nsl
9ln9DHSRAgyhUuWSNwQVAn4EdU7AFZ3cJWYpFnxh0YktMOm0wyxgX0+psZkLjf0sHkDLjCENOFFh
GjDSoOmz6OarETC4PyOVtUfD/h0FzlVHSMr5DHHYKz+RiQxpRFDZfhzT0rd4xz6SuwaXuzrhRBdz
dFIBuFt703+M3IqVf2ZMgIUZi2XbE6cMO0QFHLeiV5sRa8rmr4bawU8S4pMHx1hIRZYJcvBOPp4d
d+DZwjRHugdFd4InvlIZjwKWmhMIpVUnzg81mRTLoX8Pej0w5GhSSK+nFc3d/2w5dKklwU4Q9/Uz
fm4BF6r2ap4vnOMEYuijXLwPtdtrukJSgSOEhLehYPHsyc71CCE4pdxJEzh4dUJ2Kn238jaceuHG
t5RxRDzUdyDGKlHkZqlhWeBAy7D7MNQ00J8hZOc+CQEkjcEQoXYOUbI6nHz0wE3tNR5rn3wcrYZK
Cq4dstRNE1tl5PQsN5zJSsa6/WQdU8+uSp0Q/WfTk1xSueex2xxg2DgtZ7jXcd2Ec2Ig0duBdLb/
F45OjOwNfuS4wbNzVufH4ao0wRnsczbhFxvsaCQ/HWYHXQuPZyIZzgoPfXpNbNh2b1SSpWh+cCol
WUj5L+g2+wYKvWVZEB1Jui8WGlCbMnfdq/mZU9fjBcD5nSeX5iYdYh0zv2tj8DEEpuAd1WlY8bNR
/ufMyTCdOhgDs+8avGTQJYr2Sm8nJJYHD8TPot7xPWGGxpFzKsHf08M3YwCA6CkCx5Ceeb+eAjpa
xNPb07ChQA0SoPT2jMFGxNiWkUZZXagoYLGdZFDNUTBmYHaMp/HUOg0kLt7eAUN9tU84THLa/B8x
7nHVwGLdkrb42U99yP6l+AFwMktMkH20hozN0456YdQ8XOkZ7BgnOVW9pesyyIRCkBC/ltIpO65w
c5vHHxNJGxtyBcVCPKRyd6iYrLECaRSDQOtCJhhlmqLqCx5+T1XtcIrRitsy9xRYigPsIwOkkfNp
jqYosyri4QLWSFTuuPU6AFPD8sgoBuJ591Zg5UDpbTcj3775qlKBlCLL7XUcel/aWDUclnvcK8sN
5za/KDFddwFrofPRXmizTV1ZwZU9qQ7wETMmg0mZE1V4+V3uRskm8o+JanUzVZs/V6G6tgRDXJGf
4LGEMar3pHWnhSZE9a+uz7ek3os5chU8QdydQCkZId/AFMISKA+Fyk4C9TuC7ppGTWn9Dqoaq5n4
OpaaEfZCaEldnNeq6eN93hGivJpwtD905tGd2yJhHN5utVaNG0zbg67GV0VoDZfMuiQKm1QESLlx
Pz5bG6yCVb9AUqB2nKD2ZgF7/KZyT3USZ5vyWysHJMp7eazl2qzTRaVYraKkoSMnYO+ekb0N+uLQ
DsHodLZLWSu064oMAeKW1DgFJY22Vie87F4ABwHcBJ1+xdLWBP2UjGeE9x3974ACKYDV/LvApCYf
ZPiFxu+HUqbqSQ0pVto6sXppouiyS2iUtSyDm8cTZbgmVfL2y8tHzGZPPm+KqdYHh+wk+OpL/4KM
4VC6X0nd6fT5ACnsnGHD0ezabjS6Asu0Fjm4eJzxxdNMCrDvwymbzIHswW9v0tPReBkQQM4k4C0d
k5+IQyPXQdGol+S555yJuPghwEwX+rQ0VbYARLS/EAsbqFvlf6voAoRLC+p8OA384YP9angY0iDL
mA71FXnnfCHBDcXkAjF4m7sxtCKUUWzLH/632D3zPkMdOrk+yh9oyvQtoaZYnRx+aGb1SINbkHCi
e6qFge2F+LsjcXpHBQgWdjV3JlA21W6bNyEMtQoxFLdtjyxiRZzEQHLD8DpbCbYK/ux6N0GUeJGP
GkL768vQgb2Vwnmy/WsVI9IXf10/x4PQ4XRnSBcSfXzsmpUqHmfju80FB2VA3CLGhTYxfts7mVMs
GX20ACxEePUR+qjDpxRaWdd5CxSKBFrhTkBor/sK86FBh0Hb6L3AzrwbBegLxXdlq4o/jHgUor/E
wBJictf+7CdASu6LDBi727dL15/k/Q9k+O2mQxrkQqSXhBoF5coplOcb+AtLJQhSMIzEwR3lr4sy
bSjoNXAVdZ0NCAwiY3hzaDZ60Rt6MUCSBFUpsFwfE5omETb/v1q2LdgT+amsMSCdCNOFzPshIbXG
LHJPqzixequ0GASjGd8sp5XruvBvB5xzwFAx07RQ+Klzuy1yi5FsRJqXadudGjTpwXoY3dx+q/mD
bNtshDXLTIG/K1Jd8p6+zjW1gFbQL9FzGZVh1ytMeEYDMjvnr7dsxSIcXm7UwmFHHgOUBPMRdWSo
elPe9j0teVGyAycqLeJq9GKxVwHIHxuCRMUDo+jm95BOeDQtuJatC25NHhFgH5/k6Rj4DH4OPP5n
fEg1b+KLDB0Nqn90eREbdqc81XX7ey7z+qsAsxKoh8BKaAS/iTatPpXb4snMRwZoKSv527iYwlu7
2okqS1DKaWtK2c4rcFlF7P8syn5ePzGD1fy4zbqaKp6DRGprKqOxwb1iDpquC8bGaTvzshiUk+/B
ZxtDHWCnFULimq5GGo5Cm0Gw9tACuaAjebZF2Sf4+e9+QFvmBgBwB9hDUsI+qbutBkRlCu8yeNFg
vdzsSXBfJSv/Ng4nNBAzjKyWx/flvEQnhXRl71uAtOmBZZb9ONhHAoV0t0OsmGlFu27xYGFxm01L
C+Gh7zJWeitvz63gSyrlWj01P92/UzPAdYcx5plZZ9DXrQLuOUlktsKXCqK6U9YI4xZxJoTdp2UI
HXIw+kF7T1dKznlHNlHUjvEXMVixF7y4BegH28hIA4uuH/9p9LDdrKjHEI8R0KNfh0GTTlw8b8BH
Y4zGQWT3EgKCJnUbMFbqAWw5ikQw7trah6ztVTv/wRVL6BeJb36RwqAA2X0+jXewj38SsiuoVoiT
cxCr85i1rbo8XLJLlbP4SMF8mWYpXigUIWv6uAFBE+bIqlNVvrTPI6qt9A84fxcJYu+ttORdZNky
uYuX/KdG9S6RhKdpYo5QqDKKKi1DdpYyosOySVCmqB0DchAImlWlcZvhwuTJGaT1k9PiNBseaEom
/SFhU4t368QsZXAVnSKU0UUfq658+sQMQv/x0y4G3YVhIk+vuuBdZcgH4sBhxBNXbMSW2q6L2lha
KK2EVXd4vq8c0oWXiemOpFqhf0Rypd/A64mY7rRKdi6AO6COfBhWY3Dco6oJzqH14nJluoCh42Yv
IeEZ8+Cxc/E+q0i8p9njM9zd/4uNyEZui/BgxcfHqLTC0ghV89S+drbPWyHLpJU64wxIwgRUVSGV
zGQ3nyjUqL6E5Xx7LKXHE5Q95A1CbdEUYMweawSjL6T5bVGbDQx/kh600vFeuhKMXFlB9DeUKscZ
f2vQiwLwMOe3M5Bp4lOFhLEtV8dsCw5k2W/L9/KZEoqzRnsFGDM5M+61I2T00yKXs5ATgKdlS88K
8khtPpK1Sp67+AsKDGrtuUt5VElTjvsQoiwSf5Y9Y0REuwaClxxPLdBPRJF3XqoJc9jApgtWf4ij
lazPP2zl+Mz12xyFB6pCQqDCBX6cLN9JBxHniP9X9/LKB5GmBmgU4OiFOsGS3RvG5T5MOybGEBD4
J/A4s3bb6NEbWjeAliT4Rn4YOIjXQFHLbalfPB/SW17SIUe3USYobONFt+f0yLhv2TH6bi2t1Vml
yCZJInJhMLYlJnP2BrSpAHnneujNQBS552g0WV/ly3OZEFUDCyMZ4vXRfTcc5QuE8DlQ8yHlN9ID
W80JsM+3dxgs8VZ9pK2wRGtD/pJqSWT7XwwO+1hkBidapxnhPwNmDGgU8Msqm/Ol5AP69cyuWy4T
J3KTWRjfCWZRglzEgB2gl+5OiaWlKa39f/Vdf69HTPGOTfAE9W8zsxHW/21u25xg28uA5fSAW4aT
EAXKUw/65CtCuo0BNGW2WjMNuWxGr0BZrj6gD0ZPbsTIkGxh/eHNA5siqgGYcPQAzTcMqgebSwgl
5SY1oL0uSs1Jsv2mc5Uwjve2/OweUvoHQaiXGSmWxFNUgoCLivtabSeFPK+Ndzb40zsDEMQDsvmO
lRmQJhRR43qVyA+xMaNvXtn31UqgIA9gf6fWKonymgWjfnWNVx0CiG6PDq88m1cBHeBXIag2k/YV
NPpigj/Gk5GRFL56e1Q7BkbzaVjVHPrHSs6/K7txKyr6kfkSxpmLSS7MZwuQrNa3WW61yQfp5dIY
iDHuvV8T+Rav/j++HIHKOoyymmFaYNzxix0abbndnU0+orlLLJaqELjpV5lNSjnctoUiTq+vleSk
f+SOrq7vp5QYBQ+uqs3opE2z3vH547uEMi9qCH4c5YTX4WykDxAF8SKR+dhpRoatXb4gW0EpP8cL
LwZGEiL9hZPNjJOGc/XjIAtXAqmX7zxit5bSyiE8Kp6j++6MP3uwmppHYDMvGSlDD7QBlV6b4xkO
nS3rooJax0Tmchq6/DlJ5oOMS4lz/OX8MTTndiOtsJOmQfWqypJXqoNGbLckh8DneDpDZ4Z7ahOh
toNGjNfoFCQFgYsqZDum+fpnzkpySbaplbmAslq86FmGAU+0W5pIJNCAIgykuJZorBP/iW5d67l5
/38JkPpZ1wIR91ixTm3hTMn+he25K8cksiuimhHKM5B6fWUrTGIHz1mYwLGjeSTrmiSUczr30+I6
XuRTYAzZv0zpeYJTzLh9IMkxNmcMTpY7TFs22rwpH0Y7ivWBvi/xVRfuCEBt0EtWVZV2WZDa1YU8
wwIlYaecjabbK0JqUj/n+GKWP9nhnmfyFkJWbEeOr2Ta+1+9zS4T8BCTPGgSvJ5GyPfLqkvITluO
8/TcJIPPUhSLMvYmfWsczATuyqipxlwxizQbwDSgpecyGHBbRSWS9c4bunTRgFzw+txFfmbM2BL8
+uqJredJer+x0S3ixRCpg2fm6O+t15NBjSCnkFhnl6l/R68TXr0BC3jt6QSNhPQeEnD74mQX1Hb7
RV+F5M96lYNWmc6UJADCEq4WQL3ot+UjR7aOfhon/547v+BIjMdryMMcYat3vIqzvqKQ3Z4PXVQv
e9IgCfLEFMjAU855XaTBxCkkGf8OGoTkNEtRe7S7aAMJj2fQVRwHToFRsDytQUp6+z6p/7G4PsmA
njuWjcHC0PN2XT5KJNGgTdosoIkiZvtH/F4BCZQ8Cac6vCzQQCUVlKp8OKMqjMP5vmeeBKg74L4E
WLjQpozFnS/sLGRB2tqi05j2oI8k9xtqziYq6luj9f06NrHxicsWcujBCElTLjOd/U35y+eDhINl
a7GcpDoxe+lcsYnCmdd2c1oN2PF9pnEIb4BdCIHUiPG9o1Qz5NtQMuJzE2X7xtTr1tNzCRQ30z/V
WbFPAJ+wG8Uf/tY8v2hob5POQvRTzv1Q/yY0M1yp2cskUI9l9IG11XUCyyf8yXWSgp2CW529WJTp
X8Jn9wn3zbdE7rTItLwRQQ58M3zsZLt6SVxKJGv34wJvHiZ626E9L7GaC4oasbcWY0lfWPi3nK/7
3nLeC5Zh8NczTqoiau1ANk6ULsgDmSmP/0CMD1EswMwn0O0tW+j1czEyFegZ7xwKegwPZrlveWJT
ndeQjQ0dK2IalTr/0NlVtyThL0DWlpwRBNFdn8XGdt8Aosp8k1i5cRQFW76NgOLSvgfx3nZBNV/X
yTCFArRyE/jKMsKyqlnYRoUbPPntfRnNnqNDOV4JJIEVWuTnAKFWseL+lr/5U8t5+PhJJrekMbap
UAGC9C4fgxvja4lT831D/o1T71AqdorKvOT1qxRb/znRG6zT1VAfUfRTHV1zRibZz6QnmgXSRnTj
enZWFqAg7ZjYEgt2nK6wGsdnVpaYgO99fkgPUdybUibugirMOA0E89Yro/W7JgxGiNspOCfnEy39
nSPeD6vHD0hSsnyfRz5W/OlC1SKmeCvZdWT0ldeDxnZ2423xInN4PbWFyQkq/qJ4bLuoN4vThFYZ
Yb2ADijtDgK+S2nnL4Nw9Eob0FIwKHinXfOXCF6lgn67C6DAUsqv0m5H9NsfM6PIiwvbUO3a4bU6
VOuY8e2f6Wd4H4YgFQikCHq6tIJYL4VcYySxL3I2sYBOwSzCbhlO6zH57hFmqqTTv2BIpSAd81JB
cve+J5tUl0Ev6FmHJt7EBn5lhcXQxeBrC+9q88M4FpiTdja1JAEK7JzM66UBy3RjrbAW3Wvqeze6
rjlQjbhooufqjCsiQb4nDLD7mcAzqjHSKsjzKiAPPpdRwfSP/O6KEth3nu4668hkv0PoFo7DSk7w
n5DO5tE7WWIC1F9spPLZyKuEIUaE5/Ry6CMWg9lbUeNLPoA5cQoGtc57xpD75kSAYRjlwROeoKEy
3AypMr9Cno12GMisEc5rsHCYAp8to5D7kNP599Slu6a4nd2DlBoWPZjxlxnXEn1mldaiSKjqaiCn
EYMZQvhQZujI9mAy3sEmkLMFRIxcpNFJIR4ui8XslOvGqiJG82aLI8dtWywpU8qkksLQcWyRKqio
0czy198r2RJChriAgwuOXf0DmeXz6761nJNK8RBnArpBfzgxApOfdzkg/FAUJupqQ8JeQrAKasyf
MckGetK6P6+MFBsf5OezfM5i6qSibXhQB4r8OEmx7Cma0IBqoauxOwANtuw5q96ogmuCSPycq9mR
2wART/Fa6wmGTUGbSQk4jiobMO7xl3e8EJY7EqbA5UL7HcpODhHchsNVqI6y5Ra1YkGhW+5KX+7G
JPRebDSXVa7N2jwEtYrRTzqisW/SJ2nB/kppx8aMGOvMoOAutUduZmPSQWe8NtSscdVtSwMX90nD
HE7BbmaERewrwTznLRLSjbs1eIAdpxN2Yz76DbTPoUYtrZZTxG/d+1hTIlpUjw/K/nHd+0fp1TRQ
fN7Og5yVhyXAshvAwV8NP5odz0orPvAZmpmviRjaGLE9tGm4Q5+thsud5/UYF+H6eW39o/yCGGM0
AdUM5fJvsiYp4+6Uc63iXHJyQxTvVqjYy+SC6PNHGX2VFcfxn31LhuHAdgnpSg2VX0Vhhb81LbEz
RgLxoyS/RWliyEM02x8Cnfr0AxHlKyBeGG/dcbkkAjKrUCRFt+0u8KJNGBKDkMEPmcwsrXTLwfc5
an3cONyz8JgU0gwV0uTyc3jPk3fOFNBKhL/nHOeDuOAb2EwLlvG12SxWfBWv2eMVQoFBgyyJO4gc
4MfjbCAnSTigHD3/ZaxdgrQ07A/tFdaYLsvDO5yhcJxJSjRoFwbNttBLtDDgdS9BhsjBFWj/eGhc
TrEzIHEgRN/QDTVosPNcxclStTw4baKe4OwseNgLvKOLMiz5KqUazjUWtAGHDt5csyI4iQGKuswM
9tNtUCYGzrDoqtWcGcoAfb8QrOUaSrWNWTL69D2oYQthfUUuNvEH1KV6yF+wq4KHVH9NdroCK9wb
5hHIm5M+vo+phI8YGjQynBn334BfmCNIjAsX/9DmAN7Lp2btQLKC9cgKjF2SxkSFm9GrRQQB3imq
1pC+SZbpDyFZTHkI7629fjrdzWfSE2Qvm64Hz5ouPcsAdCF4hgJVSjPRd1JFS8529aIJyAdTg/nL
IuroOEZLFFMsGAjnXEgmIrvsWS6zeLyXhAi6VSb/WEs1Af/sIxjGfcunkbPS+dBrFusGLy+K83j/
KQZ5ep1X8CJcZ2IYA5qyxaXo3PSLhLgyAB34HeXk5a1xSpEblfssNkjnTYIM8ei78zakvaVWny1I
N/89ewO+LILa6IiIAWr+fCd6l6bHq8Rrvyburdapbn+XsFLy+5sXw5R3zsWdFdChq9yap/W/0QsC
QinTtSTDUTGX4vJ9I9Mz6hmopsmT36Y0fdg58ymDURy7twNiuyaWcz1Biar07/za0qQh57ay2Ekl
1e/IsgkSlLPvz0bGoMkmpVl9Uabu2aBom2kMuFCP6+Ehbz8XKymwzpxbeuY9yi4d8weH+mo3qfTa
ABhfrX8KYAI39/8MiD/fXOexOrovnF+qnGLWC7TYLAyn3NFHtoJThIjMVhT7389IH+IsyNrlebtk
po7uDXp7nX9fR8W3MMl001TTC0PnCNnpiBP+8oqkM+Qv3MfbLuy4IG4orJWxkoHr8tjhNk8EYEL9
Z5P88dGqUQa7KIgXxsTqMgnnyh+BDTPccUj09PEMN4ZMpkJKY3Jx94HKEEQQ+ulkppWsnS95qqPd
WLyqrIADLp0pMegQdqPxH6oA/tHxDZXsmlvlawM6+bB63H2nDCmPubmS/gC847JqAtzJSbU9adxg
8z2ZPnRPtuYtGHQQtmdv/gHfREb8e44tBAyJxHbTt+EqjyaYmXsXgk9gG4YVhEcnGC6U4hOl3sPk
mQF8mHs2Z2MVJgpOL+SNYuFeRy/JspeWhKTGkqrirAaf5IavplYBaiJ6WSQMuzUkOq8kfh1auwVN
LDYGHIERWl+8Zr/p0Jf0cehyPYWYymDRVoO6s3Q4Ic1QlXo93RDMePzz4nYpr7Y39YU3mRNqk3v2
GANSb2XKuGnXDrBPu63ngYO3SQGHCaxFYINJOnA3oJM4sIxLcPsOidedLfO21p5zyIKeuL99lQrT
xFSbSiPa0qqTJVoKcqXAaWkyS/mE8x7WB6c0lAaByWimD4ZaRrTIFcXnln2oXe9cFEX3R+UFV8x/
ES0h3D8Do4Vn1+bA8cht8puAyMSMemTsnzYKFU4nLJpj8mgzN1KolJzXDPw0S2BGEtxpMcQGPWzt
1g2e5UC+aRIZT8UrI5/vrLIIDVjBCU7hD5tKqjZWn8guM2Y+W8Z/f1PCEzdJA9FdrRbytMwp+qfG
lK94s4ROmDuCiKdupBD3N377a343UpzuuQNSR2mxFlsAii13gJT0OVoLSMgkXtaXzzuJ4hAd2UfS
KUkXplFptcooCpciLlJIFXoGnanrHkce3m1GPgs057yjEdFgOKoyapvVNGHklDN7Up7OxIK8svoh
iJIN2AtoD1iPSl3JvoKtUNiDRsFzZdE5Grfb8vBCF3lcZ2ohWlI9tLcoVPs6Gd0ijzgVbrZkOLhM
JbJWerz/uJJYHQCOlSK/th6AKaj5so+WwDlDysW0yrzSuyj3BwemMhuU1/kLR+lmNvOALJw00LZj
Fx6QYonZZt2sOynqwhACBqOgCbZEvYXHrLs2Y52fdWsFydOE+krq4ZXPouLECsigpPTayuFJD6pl
QEOBfCuhclubayWqUTIg1wq6kH+x/MISac6T4daiC26eo8CiH+IKU3tNuyfn3Ut721oKZeQAhsjX
lBBmIxw4UKsasm6VVpmiZU1BqjBTMx3KvGEjrrAvA6uysAz1Q0oZdG6RnQkBaqq9F9hv+5ky+XyB
CPC+VbfsIsSzZLiTrlGYUjKm6I9vPIDIzG+P9wXDlEI6JSQN76ltEKyCRLW8OwJp/moNwt0EEqtw
k7bued5nhDmgW3Iq7jDs0bIAnmXt44C38NfASSaSDDFTDt1S0xVlG+L0woKgCgfK/wB7m3KqlXFF
XAVxrVYdW/uDrhNUvn7/37nTL+VN+FjJOt5M0ZkzN0vrOOWBtHotGfAy3p9h88UA3bgRqMbSJL4i
VWpn4mWyYcYPxAsBhuwSEcr63Cn4AX5/E4H35G91nUB5VY3jpj4T2n5f8uYBp2RSr06qdoD/7aA7
gKPHZuH8WLwQgVH5R1eCw1OyzzkEwMTBzROYWF3WLWB+6zSg/d5MXvqUuJjnd+Kh21G3r2lr7dSK
E04Pt45up74wluE5UqnytcU7jpkSx2KZynJqDp+m3gWZfwGi0tM3PywdRWMkvy8WzG+SLuzbFjnr
Li9v8nkrKLjxncwKI5H4ppOolKvktGlkCy0nigoF0Wp4tjeqWfjsFA2BPiM3OGbjrKqcllUP5hhz
01TskJwP8WbV0hHSC1rSs6Hme37et4eL5BQkMcxX9igOZvN+CweZdk9wgGxISAFNb/2NQCGbFvp1
FLwVdsNDaRsz/6EbQe9UwUYeHkdIDNDVODu4eLlBLLdaBBbwMBjPgmxXV9mNhFsoJN15ye5Rx6lT
OGHwiG4dg9CIvxkhKiUOEE+j7HWv7xlFOe6Cmkas1bin0OujuOBqS1So6WarJrUveAgcTv+DlTDj
+alcrmzYLVR14LkftSRlhChU95AwxklxlwqCVTnsLQADwZr60hHREfKNFBXlQ3TtZNzaZsHD7bOW
u3kkhsC5SgE5PEPLjtGWKf1NS94nT3OiSlSQdXvTT9m73NsA3okneopKwey1RG/m133E6B1YaXbs
obnJvBsvfboD/LqNbN10PLwm8HMAt5sytFQsQkKj+c6sZBcAq7d9VTEbA/A8ih7E4MPaOLYFrVI/
WwnDnWG5XE4UBxnhwsaPRQ89L1Eb6mf2jrpZbQNIUBn4euvH4wu1fvjSj//GgP3IE+xfE0Gojn6h
c6y9io9K0MBVsnMbawjzcJJrfXNXiCaFZ1S6aamNLJMP+qIs9teaANHN5R/bhpWZ6nVlrFFtV/Mq
IFo3diXODiuGCyzV2gSODu3UNEKm3EcjdRaqKhn0i8zQ48iD8Af4o8P1GVWauOUSLZuRqm6F/Jrk
N0lHNjiLW+C7+4ZmkIRH0BsdTf8TpWL91qXxrIKR7EaKCRqH6nuM8xYM2urdeeY1iYoA01oejFZr
ePSGoy3R8y4pp/esLvd92RdBGPnyHX3J+GAqOHlGr/ia+TqKo/VlW76ZZmJEsixpp1EqCMBvyW69
4v8gbQb4jEYTx6x0hh+j3v+8fYiQuzvT39gXtPxZlq1ee9Ti4SZX/PzzDz3MD9DJja4QBqg2rPGh
cVDiCGUPYdxfsSXHv7Z9CW5WPRVPx0+uAv17ItgnLMlHLokTkruprEozxhRb6uhs07jZiL3AnYv+
dZIEUQaDOE04X4rbnWML0/wJrsGVOPy9y4PTGqigA7kB8WZWKfLvrVqLz3OWuu2n+Cl+ct1q5aru
natq93GaUu6MaRAAXl7eHowmmxwI3maVwt/iYrBbDg92cI8dzqrRpHCpM4xyO0ggfcMbGgzDctFP
pUVays3T2zMaxb3tQaLYLf+io9y2w3lBBxBHp/9xErHYp6TZo3CL3idypmxf8vhcrLLgDAy0ccIr
aD9ArphHFWmc4EeLpy0Q5J4sJ6ve17S8AoiG3lH06M+8CDJcCQvreh70iGktTa9jMg2DfRXIYhMu
xwrrNtZp6pRR7CYJb1F+ldQBP5yd3nD1cMk/z0txPxWBgHVsCV0XaR8iA5Q1PFRTtP72Vof3gNhM
D7Ls1C5RZ+DAxCBQFbw5BKcwIipazk4oOsYIGOheUvH772raLf4oJGMp5VmHZiecebZV3xhOOBNc
0NPr7q5ew93sUxV4B6q/Wd8ur4cE3cyWlUWFc77xlslQDe4OEud+SEtje5LmiWDZzEemUUyvukQH
HgpoFhKhKoEcY/TZ7M87OusjpNh0x/5sDBduEwiiIQm0+3m93c4NT5I/v3N4HjFwS3La9xlnpkIn
Rcj9GVVfSLXrrVl9fWoRyB+fuZiSE3QVpToCK5zlBghtETHsXbKjwc3Vfokz/b0vPnHEeN1wlPpg
RcnGJSWHHGz/NoCZh0NDzrb6VTiVEP7ngAoC9xjYPYYB8U0+QYfE5UCkTEkwY4TAC8gpyHD3aKht
k/8D/xIaBDEQP4KyWQhD3JYKSQQsrLHVYdK4y+ymAeB82/h/QU07yUzF9OATuiEvubYiaIGUyBJP
A+kgY/DcjGSOONfPPQtsA5LWVwX/n6WhMb0QUj+y6PZ3jr0iM7UPyWI2Ty231qEeDJI3qfNoDNNd
wcU6TTLMp8yTo+Gme3gpnVyTiVbLMo1M+VU7mYZQ8p5Tr5dX8K9SQBF08e+UxMIfAtc6s5U5YVXk
9ZzU0hSmFqjnCz1KHzp/tN9oh/J98i+bVH+bjJhAa5bUu2sn2P9a51Hta/MtS3/JwxDfrFGMCrsX
VKeDzA/Z2NIPpvfnz/uGgPIO2Pw6v9ZLHO6b2PEc2xqtnCsHSfJHZTsuRhocIA6S7OFm+ws/O9C1
FQE1gZGS04FTrbZCRabdoIPBXR10q0XX6R+daW1JkaOKtojRoRe6CRzTWlQqrFkDSJq/RB8EUYBG
Tnd2cvtjnZ5PXDNGqVSk3UwlX8gtiHsci7eMkXPGtkuKFMu/y2xLAua4oYw1XfFxZSZzTlLyRVet
e30UUjbm9RD2daR9CEYEWxk6XjL0l6SOWYPNJBl/2uq+G5BnnxfLg62uSPs4y6/b4kDu/YIoB1ro
Pd8Yg4Iv15MKm5GmX4oaMn/5S1L4tlD0zsxzFZu1Sc91Ji6ACgqE8wPRSQK+feBfLDEHIa8BUlwh
lqAhjemLKAllsZnDVH7uy5p7XHeCosDvC3I1ASv54MKOzHxlPSHUOjaEIsf95rKf9cF83UNpH9Q+
F6JhuXLIPUQ8FNtZLTvb0K2XyjGpQfGbn+22m40VcAXDnPsFOA/Zbh2uNNUsxcqSmEC/QxbS7Llm
3MU5AWyiTbI349MCk4WWz8cGGn0XVZ1svrmUd486GlmLm6JHa1wrL96KgjWe3yVJsIyw5Cgit0Ve
tsIwgvsHd5WqXtPTqHXpXStk9T3Qoz516B1E5u5ZhoSXmxGTFfH3fbdkP3I+bWLe+Ej6wFjF77PQ
qftMvTng1IVzb3z4ZISn86M/eWd6lNADGYhjkoVeHQSvC3iFmzHr18ovqK3ug1YQYiCpwSEqgZmw
XHvMqTKaig7E1wcOCQKTY6bBHeVjM/ro9OxtlVk2EIUu5+HcFXhtYBQ1EYkQf1yjOdM3+48YNZIe
eZ7NBI42odvWUDfVS3Eo1f8aF0l1eoFpvFG61m7AqzpaL5pmYEUjcX6lkg+ndKH9oL0PWK96tV0j
g8HmLeE0dGosuiMgetnN4w18iLslUEwVPVkBwnfxlbQH+v5Ji3OcJMilg9eRR2ivDlNzjIYkzLoW
BOSVGmnk0/IzpaKzbs14lkFMS1AwpNqpBJahRNrLeOuQ5cJpneHwcboBib+bGsGBNqbQP0TtwfGf
yGzIbcIQZUBJr05ybUEKVsR1ourNHJxNpcKk6PrjLWKysG1n3FZ6eYSDSKGJ3Jv8Y7oVBVQv52/X
cUx7SUJK961/fPHwT7jnMH4qBe5kZQefFI78/yhjZb6MYwS2r8jN12l/FueLvmNbffSH7U7m8HYo
7S4F/oYKb1B7bK/MMc/3c0YcqxaLomAtr7JkEZw8mfgYmhAWxSQM5abHb3CyiY+vee1HdOqVFZb4
nRjqetcJfZEjD0RHSoGoJ3F0zXAjLeM8qDR0FbCJkTByu4S0HJkleyJ2nPYfUh0S5DP0foSqhRXe
CG15rOByl5wbQpoN17qK6EwY59sRusqITnMZTTQZudqpWBzsAfIyeNUpPukXXWis48yYzeyB7xoF
j8KzMkVzN+YvnfSnW1C+9YK/Dju9+a9fyyJXSAlWOXsbwsQt3KmUPhSSLvS4jtpBwX6+A6Ah0tMD
wSK+HV6rbvodGC6KD/DeKqnh1NfjWawR6QXSW4qOWaKeg7g/WVo0f898g1i1ZlshwstDnFnZjaGS
opYCOu01O1si+6K3bWixc+p9gnejQvcsBQDjKscVHnaGUQx4m0vPkK9DKmsBafyzrihZr7unGXL+
Gbu/sfUFXqLn9pelN9I2FzMi8uV2d2SE/0JaB8jWMpL9N0UfxvkaX1QbdWBNcsBVvKDXKKvxOg5x
6+nlakd0+/RmuszuH7KizhFwqW2u6DcoB0NdYBOGMnzXBlrFeQPKJk9T1vohzgH1XG/ME6phkNP8
Q4B8I5diwarJFVz0RviWGmK3vGfFLlswvfDmwX8vNcRv9TCyniKG+5Dy0lJoNnruGF01Rc4uSPwP
7dRkTFVtZ7liwQFTHi2BF32ZaB8UsDvhbe/oUzfCO1MAdX3MsjW0DLEnhpFPLgR10HIaRad8w4Bj
AH4xfE2OIm/ZfBgrN+2aJ58utwNctKA22XkdLIQfDa6QOvEz0jeCdfbC758nWF7TKycejr1NkK7q
xX+VJQFlgHPjaPrcAx/ywMh/CQcf5GtwserywJg2tlIhS91+fha5Qh6z/mOK4+h1kbfhlkudIaum
HI5kD63hHpqZDdAVN/nVjRb1flW7IMZ8D+pBcRQRwXskKqCQODicb15k6256nkClwjdellstC8KC
DZOr9JHQyh2ccxDVB5Fx4ntUTn08RJjvkZWfTVS7hBIHdWtvzxqWN5W8YvyyIz7WGOm2k7p19o31
Njpk+2qRBU6bsXJqoveWUM6Ls0Q6vgcSNE6g1IItnMMhb6Pg/Gkj92MyfOxsh2HX0oLtHYypYsL8
00V8bHl55kRizmH8gKlBrLMI/RjxQAUwxE4HI8Pu3n6scX+vpCa8N+6fh+O2Hpl1pFrpMB1WGFxl
vLQ0etuSY2cBbxVUsdAiVqL8IXYvpamWA2qRbgc3hC8DwORLFDQvsKET6fOO9KBUKcsSGdcPPcyK
JUUeb7Nz5SKUtMAQJkdpxdjj3FIRlFkhj7CVkT8gB4zhaqU4/LQk8oS/6U3gakOYmjSXZZVKfFUZ
2/6B6Kjnf5WdrXvwQPv937U869tJbsRubQl6t+J0rfLOH4CUiOlmIyztrbsGS7W7bBfhsW6ftNdR
XLxYpz0cJccQqTd1qX2wQY2G7eXjrgM13yMVDL1Xj37JgDjCU2YgU2nkoP8yhfBk1apsP56lS6l+
JIdN475x29LsCvicmidvWGobETNacDH7Ykr797vmMt7G3vJLZyzaRHLJ5d8UhEP95gX0eMBHww/e
PLgPwkChbUbqD6fapsyS2oZnuR9Q8NkGu2oqJcJG8LVW2xYzPn3HCU6HvAodx/W0BR+AoFqL50pF
CB5CCNFQGGHvMlOlTE09KNKVTWnmMufRvbSl5G2t4zUGMoznX1b/mYD2Kzn+FELGPvVTdz4bUrCh
fQqUnEpbVnzbxsVs5zWiYTJv7yk1s8+0TgozwWl8EUGYAisQdict7oY9suJdIx8b3aU2kE+/6V1a
Fn9u1kPnmyks4IQ5dIyqXhXduET6Ck8kW89vPb1DLKn0WUz5Qd8gcJB98nZOdHLEA8NMuzArmhlU
yNwmj3smDihU8/6uSjh74dH7/5LlNSoF82iWv2qOqRNIvLCArhZNOAt3pA4LakC77oclsVvxP5Nj
bf0C4uq2OhMtLcVl10G0nA2N0sQc2PoSdT+wTUPqxSxUBWj0DoxXifrMCvxl8Mc7ZuNU+R11Yret
GzshUWLCL1rDM369KeCmCyBd5XB7rxx3nqOAHxHbkpfgheDB/3xY/UthC/Ho5UHDIGewdN6xnJs2
9MLc4h0wi5rTU30LKNORfXoJfQ9/53TWdZwIjEA7JJ8+vYfgc0ujuog5nCvw/DoMx12XCkXhLFrP
a69YcEfcZ34vQjYoFouuLjNR+4FiBPzncCOkHB7n/QXzG8ZVb1sttSoEr0nqspTwD68rdZqnQJKO
r6gkva5tYRrgHVAbBBtie5wO/fN8Qnnh4NejCr4Ecb+xQJ7rX93AjqWY4ym6WWhjNu3s+fRz8l0b
RiOfiLnjbDkh/lq2bwOeMJH9SRAiMDS34a0vwFc15FQZ4hsHIhVW2T5eSnIM19MyPn3qOGW8uvmk
Jfu6rVdsfp5d7BG59Zn1SA6fxFDMWfa1e+4FaUI7qabsoAE7QY5zPGHo4FO4/fJRPVJFVujjf/aj
nEKjbZm8Cs5t84IEgBdCbFjTNQ2LqDdT1f/leovEpsnrZZG5JBi2w+TXe/NCSPRM1TmKdvp6VftU
oyHTfJKf3Sephknk9MGSI5KfcHnOkSB0tW7wdN5RiHp9cN28WH4R3uSpe282iCi9vKZ2W2LNL5nL
ZiQpjy8QXWs86t6Xm7cl7pJPFm7l3q+O3rehuqHPj6EjVtOFzyP3B23Fe6F0iBH7KakLkbc6z+aM
ajomYQRzsf0QiO0Sj4/GgOm8QqBldfgRpUFZtVpnWQd6orBdHy6iAZjg1u2cojeeXK9Zzfl29ik6
RBtlFu0iQXxuAzgr90vJWgAYhcQEvJmaIW+1WhdHrxlILZ/MzMtbtgccpnJ7FfQPUiSTT65Lk49F
wgMDUcVy847Uk/IhM8JCOgCFw28PLEm+8PsaNm7jLSS0HU7jhQxZJjqHTqvEHeEoE8DfQjzVK9js
zpd+b9wx20f3Y2/RIF8a+5uBviqgSjzG26m1WQR3AXknvYnQGlHTVMkC01EV37wxrQJDpUqlnJGJ
e52/OgCKE18QFm6kLpvOZl+in+JXikFUw3pGOrV1Iuy7nAhMyOXwqZ7TJO4gxTMNyqrlEp8tcrIi
HOD+wMhFBU3eOdafBrEbkKbonQ1TD6Hq9Q05B0DLdFv3DOaReebHzKDyk4ct7gqvf4BJ5u9aGCvq
RRINtWxkry2x//eXhF7xYeeWnIVGjcrgco9JyvYUJUSQXYwXabykbsiw7N0eEAEeXI6utRPGMao6
6p+XyMcWeIL9ZvGCPvy08Bh1lww1rVRNwbaY3rEjsrgzaVd5lN4WfbID7/J3rl2gOM/1bI0lfZUy
OTse6N1tgWq78q1hJkcpkSYpTZ6VDaqDb24UWsL3LZwuUJ+ADesYirQDavZfpC248uLW6d8uX2QK
x1qeFKGLntAFDrlkoWpAWciwWfVcSL2gt772erFSnHcVVglVzLR386GOYXeYUEHufPxFf87XV5CB
C8mO/dgOqToAYjAcYrahQih8OQYzK0cCK4PnfE3nep517pg/FaWaWa4oEtG/oxdrVjI89VJ3dDQO
vjMP5IK7GdkXK4NjTKmSgLmvKr0klnUDajbqeTI1JzvokJJ99gAf3LAiSpgAqqgk5cnxVB1dDLCr
VVnm3Bz6FMzy/3eiF8PU078iq8Hao1szbilhzU1ZM58H1GlmeKbtOxZrFwJE3xpOEAYPzK0dX7x4
7SrnopOHew0vWuYQkKQiB3ppa+9EvvoQvumj/+mBeTMGEFSaJTP1SUrZER/B1Ky1AyBb8o8isJUG
9cUNWcgRH3f9rY+9aZUiwfNam+jag/0b/fFVNH7UQIbukOpPO8v9qonsw6/+FXg/zKvAt4vSqNmh
C5wdfU6/Nps/y9Qa6BXjKbhUgoClPvb7s0KoLoHUe33kjVsCgl3ZTWGg+i+XoJn2XCL52STXGT/l
GGKg7ePSD9bQJ03DuQQ4hAws/9MV9OFK7ay2UH3mdsFnHL4rE2IIA5LJ4kpxiP069wd3+0a9ovXq
WxHlQ/pENeoU6UUyiAIZSzyn1ynrjEhB2336dSSjQfA1exTTUS50DD24L+PemdJTUe0Yi1ZR9zyA
y2I94NHF8CJj80wAFak7miyBZiOFH4+t+OsQ6YO7j9VYoxu5bm3s3yAMcnSoiA1ja9N0UNvLE709
bBExD7Mn3l9jgSlDzISK9vvYMuhAus3PCP9P0Z0s/u8CwZ3dGEXAR+ptf3o98cHf1k+klkQ58Bhg
5IFsdjjZnhFftofEr2ZGojFG1JLB9t9nELYFqrgh9yMmMcccA4afsEyuH5hcdhkZh6fqRqD5kPQO
cWEQAnnKNk9wml2XvELLEx+3u1srMa8Dix5Yg6oa4lutZ4I1XG2EIQeq1PmnwV7XP9FHmt99Wi1R
S/adWx3H7n6GBPU+0dwPtXHjPKm1HVljke3UMDiBzemnkvOfVLac/EgDWihOXeQylNaRdOhffFor
qDdtanWUEEZK6gWpNDf+iQ0DJ8zggegfTSY62neUWPMJe9lLr4UT1RDjYYGcjI9Ep0s8zV1G5Oxw
88lpYiIzrBtpxKUMm9c1azFuDsDbhCQhK51b2kIvj+FyNsPwj6Va0DcnLcHBMq5LKtuWK2H2woG+
OqOGPQv1w3cgF4cKWk8sTqkW8k4gZC1dvyyQ7+1mdxFveQIy0WT9XAKvk2dTkxAEt9b1WZAaoM8R
J4aNGWe1/MBPAqeaR22iaHSb8rlqmYeTvmNbp8vlMF65zjZ5eIXhI87xLNgwvMnM3+kLt3VgBILN
RzBCgDUaL5/IucznbK0u0Jjl12FheKQ1KI8LxsEgy8+KqXSl3DfZCxfksYawMJjO5IIP3LJeVFnI
CEHUeaGpCqHZUKqyYARdOa1iIaRz0fLIess7/HZzE4Bet4rxjRQmDLvb65KJWFzh8ckgQwsuolVz
s+hF1rb+uDQu+v3COYCT4rngRFng23aI+8LhGrZSytwvbf9VUmhuu1YPnQiYc72mUIwEGmZRByMm
TIiGsgi+pNp+Z4X7jNNMvkUQ1jeqgYUu8Okq4maTMDq9qWlmLbBJY+vgv0cA5JcAU57nu4ujS5/Q
tn/Wl+lgQWBstnGcKywlUKmOZQ/sv3f11yEZCoJqWgO6R2pu1g9Rz/8HfVpQWzbhbyyxp9TnCotC
+0m7SraJlW0U0sR7mi1Ta+L/WGFNrOeU811Ytj9izM35UJolJBiGWM2f37y3ZLp+BRNBSlklIJoy
9xCI/QP8jn3adz7+hixwui+GHSPzCLOErbZAuj0mWxCkUo9NwHMOqZCxykMyr393zZR3RCaYzO1F
lZ5XtuRQCj5f7SbqYvAlOid8H1N0CecRVz94WshHJYmVbRv0MBFDQszlgQh4/+GN56I1oWiH7gih
93BTVfAeko+0a7CVTLoQIr88bc2zujt/IWLRgJ5xlQzCW21UkYbNokPNpL54DGbUND3cFEYyRD+q
EZlEqMMZpsOloEhCVep9tULme74z4zMVAe7z3S95vKweWytduQHgwrdWjwKC1M7As28okLbTWrpR
7SfoAj5LDogEfY3NGP+F5+QQ2o/qbXfLYXZ1lO0zFEOG+sDSTV/wwX02z7kJFR4T1KNO5nl+gJI2
D6hNqL7Z7PWmL4W8u6/w/3ZxZsLQn7IQxDw/t59+bZU1dkMQxijP9h2FYt9X03xb3Vpdaz7oTxKg
uSGfWqlCa7hrveBoJndHfWWAzHfY4Z3t2Y733qC+Mmyd87HWTZD3QKu3iVMRjkDYvkEGCaHWnnUw
c06xkpBEEJjuv+x/nee9tZ7fDELGsYTc+yInRhfzZoz+26ZskA7EeMOQs2yg7Goh2nALHqqiiFkh
Ox5InvLH5YhNdmNWQBODgMfxVUThQ44VRwLsMtbt6BLpkxewCU1CaQveKS7lDwlFv/rFAqGbV5Ax
EVpyJY7SwuF9ZAXm7tpkZD3L2QEO6XY8MeNErrirxoUd+74kTc/Jn+YP3dvWomOP/508kC3Eg5j+
WZRfA6hilcT6LAZCt4/V6j0pDu93m12wqNGF7VI4K8NAuIetoStf3amtd4xJZ/uF/kKKuKbA2Jxp
A+XpN21tbDWH0bRoKjIZmy3SpoYav6GtbGJChYzdLj/n2vXoz9Q3p6nOWHysfxDrTiKkQIQFGby2
CO+j0puRJrhRlFDyf7izwoShVVFN4gEoluo49J/YNLnQcnguRWcf613sGYIvgX2/AXeeKUvKwg21
x6LiCz5hi2WW/kYVWBj1Gaq+wDZaSYgIjLwTWaglLNHbQCEkccOnVTkJelUyKXzym4hNUOx+ux1D
KlC69dSsKF4vOmDxk0lo0zJaoHTPF+po2HuwKpXNU9TjK6EUlvVyYNLlmcyU3y/fuMc4iqvxY7zx
FC8Gzqmdlj8EnK1qnWj1lSU8R8f9igbNKk9eERDBJqnRCYqDCs3ftW8WF8zGpaDf3+7y1z56ZS0O
YZKABhbWM/jWnguGbEJObwTMbuHR8n/kdguCcPpEKAmdVj6Vbw9nSZhQYD4svp0ZG9cEbABnkctr
nN4C8Bpp/Y5cEb7xIK+teCc33vvmhrrX/cyTHzzsF8Wcn82LKFQXSV0uRDIdWqfcHOqR1/czP1dv
obZs54dm6tOeBaOxFrzv6BhvkfcotG33Me2n82fluW8bspPgsSRxB83gqfEICV0GfEDYboToa9P2
f5g8xsW1yAjW+lgzRXz3nymxUALotht/d/wAixWe0luszZXosqw81h0cnHTKJFtc4iDo9vBbNWwP
QLf23YrgR15aO1G14r0u2pSXECHmtf7oDSLuD/2OzzsCK31xn0JZruWMQ4W7RzbliA3ZFTLfTzGf
hfPB+Ea/7Loz1O5M2VB25WCcpzfe6c93HwOtu20shTAqby+VhhyzasuQlWm/sqsKVyRL9LQm7aay
xVgUWixSURa5ofOSXkrQTJpOPYDyGCtJqEhvEHMw0m3oYaNPYhYlB6SGMWPtDZBvPvuZtq7oetzX
MeZtwKMyE1ahxoOCvzeWZvzapFrtwFeWpwM8cxHb1dIBcjf9RuhYgmjhtjaGQ6hWfWoZLIgjPmg9
Kq+16kZkWcQVWtXlC1cfopXQ+EgVG5EhUSAII/R7dSkAL1MMrXj3KcJVmtR+BxCdc7A06WLmGANP
FJs/L4BbSsZCY1e01bg19OTlA9ApusyEe2pZlew5nYrQm+d1mMTZ0dpzTUub6MHEELghx7rqJx85
+6AUUREFj+sFUQTisw39wkbaTLK3LljTFtNyHKqvBRTSHgb+BFpXApxWPFxeLeijl7J6DyCgXYfO
xVN7zxOv09tIghT4mhQrvaLydMP1Eaj6yGPpu24z9G/0dsx7/zuAFeqSsvwbh2GmZpweCLEWUSSA
Wfvl0nUjpmr7XGjNNxaW+ET2+6HH2MA9uye/ucPWHNZrjqs/u3I1NdNGCTcjl1F/R8itW/S/9U9k
qXV2GYv7vvRmAi5UVunrvaRnIfZWiirVQGNdcHNZXbFLo385mJqGt4AwsPWNjQr68wbOkcRabXOR
FdlT+MNBycaV6Xfku0l09I87SDdmx5wJu2pFFpQkK8Y/Z0dfAjAUjN1XolzDgcTZ9U0ovNAbmHuB
FbaxyeuIjg7pDm9N5SxwmEnBBC57+7YGBj5d8L/o1Z6+YfHrkYjm7dsKwFFWMnmGM0Eb9aJk7N/3
gYRocRkwgOsJL/u2l4sk9hGnltlptzcm6+GzPbWi1n0oPQkScf/7PMQpMJUMGpsIpPsfJUu1n2F3
sqV9WtZa6uRl6wAQf1TGE3NNPX5azO3G85MYYlGKHb4FFBquHLlCsFpGXSQeeDpUtqmdgR49WGhD
iTv3LtxWZaY2G4VjRogwqN+8arkGqbGiawiU1hXn7IUJ9TLc7LKhFmgmNXPQJ4LhMdW7Hh6nRvxU
2211tL+BidebXqLJ6N4rbpXTYT6/0QaRvdnSOauD4pN2XRvn4NFRlgj5u88ZwsPqDaEgrbbZ5tZu
wWw3CrBPlb4gacegCcIm9R9Vm+xUph/X8r5GOgRW6vzWTWws81yRPMQzyyMj8S2SOL8iyj0UJClu
GOH4MJFj919MBSD8LbNLknXpAhIlFnwi07AgQz5AjHdgZztmhcIlWZYA6yVhFPU3QZxls7lFBgto
VrSWh4joKs7yVVGWoJ079aZ+/nq4OHjmsmyjdZrIXv4fYd/nHA14I9iJXsQ7w7yqETI1i2PQVF/M
98a+cO2bnIDZyRM7VejoudydU1uO5eENLss45kWRbcCF2hwDs8R52ajqFT45Q8s+xcrVVRji8SYo
tPnZBVVffECntTJEz5ZIXCtvuYBxfWsUpv/3XRZEYHKEPMZsebPHSEXk1pvqTlmDc+WOUPAtRwnc
oV3w0JlTQTJXV8TciBMhPgQo4aVV/25Ji38f7lBiXPP3PO7lF2qt6o1J4EGfpxJHUAQuWEbX3FO3
pXcGHdyWDTm4xozwdp9xQ0mlaCB+T0JaJZGlECz6xywbxtLT0VzoQwe7xxFc3s+HwHCnn5QKl9Hp
UwEN9GFSA69ES2wY+i4LjdAQqI7HSkdBIyToh7MZV3+/J3Z+3pgtel2ELsZvdPs63yDxiItllw+i
TQDYWj9baxO5RcBXs9jhbpgscnK2AjWAQx+2bGfTqQw6NL0+0jshWVoKFqycKkqybajycXR9eIq5
lLgbBNy/0GWc7kZ71tsRsjrYlfzShg77rs5Me5mfNVMwSXnhcud/jXMdiX+ahH/te9WJbG82ztPb
gnUbeC2bAEx6LzaYOdriD/A8NEnODcRbdycesOcesg5F1jv4/kXnojQOtembqSQRO17vlN6+WWCV
rKr7KKHWdoAKjK6Zb0UZQlkFY4VHI7x2NqeOtSDx0vCk/wYbfT1/myKsbQLk2+go+vAcBdkuDW2V
2F56/JZn9YI6ibMWsjwbpgN2eNIUODSm2FZ7zHKcfRxUaOm3/FeybWRTvEalTXokGNRx2MmpqKfb
AytF1jrEbnrDNsmAVHKyPV9RWO4JN/BKta69JSWSBaSPW4D149P/HNavbmat/vBUuuA4+gRVQNo5
zfstZIV3sV/xwMxms62JOoJCn6+H3Mjzt3F0+h93SbJ8DuiMXeyHS68KSGPkD45Zvm8ktMDDDLOl
+g+5eRvKZ0Y/u2E/RZx++nKfab6i9JqYvPUnaEoAF1XedUThI47xu5w+LxWuKKigk+6Ie5ILVubo
cLHvQHW6sD5i+GZX1wZY0CdYzCtjOSOEQPB9dSvf6VOdTJfHY+fBNVZxTuY5c4hEghotsqOmmGMu
xtBkC87LQL0XCNyYlnw9kT/6uIfet/x/3Ev3Fg9imHQSb+i2koPAY/2msA2O9iLqbLG/zyzGU4Qw
08/eCg2y4A5Jv2v0ycDA88ICxDr5GdoGf3kaQYBNzdrqOTEURAMsWtP7ME8EWbr6WiBzTMo2Bzg+
Ipx7qvfquzv8EqF9LzoRd1CYDfHtkiQ5dZ2qZa0+BPS+txSvsdUy1603eJ39Q2Y8fPjUibmtp3gZ
AFYxIc8PzGIgL9H5DKr7GsLTb0KSbeG5piPZ0hvhPHhy/X1ZFPQ+1FMcY4c0SWHgx3KPoy5rFJ4S
cLdAgEh2/SS6zVO4gpoFJaowqCdwFUiJsV1RjwtiybuinW+Za5mbsIGrJAzCAkFC7qEMN2n7Q/N3
gtC9ctRJYnteEu1YYJ/TXUGFxW8drz8SQLIDKkYhZTI9JgXvDZWSCAmPsAGpcZmYMvpj7lylCQd1
T3VZvYU7851Ks9iUJzxlhEVjWcr5t1VCECPmhu8PzlqAUsUFF3hNa2VQVK2ZnyGZViS5C0I4iZ/l
RPsy0RsnX9Mu1stnfdaW16eQpeFFLB8/kX/nvwi7sAZJEBSngqIAkPv6Ij12bSNPd2K87sEluayn
tzsqBdl/QyQ2qGh/rX7o4qqcXQoX3ZOFEmw31PtJPpyEB4EGy5tOfxUXO4Fv8HC5/mixG6LDXuy4
U/puIbFsh75HXW7awd6VanNLITYTXYJNS7U050qz7v74R7BuVgM0qNqIjo1hMTorhzzf+WnxioYh
wQUtV/Ym4G+p+ZuyDzjAIZg9bfLocF8d2zUHwYZ55vTcu4qNkeszJGJRGvfcEHc5ggwIgVCA7xeL
1ipXFY8YKqWvzfS5WfcS3FbYmHoBGDv9+GLX0Ho0a9wOvPHVEj6/kkrgJH6YYPn8pfOWvl4FTJwu
+gRpJPwdBl5i5PI196TBl9CCZVqg0F5qstrLWJLdAYYRqvegBX4wK+sBOdx+RG+kXIUBl8huaGC2
443TnROPDrUz2DDBpVFzH94hNl8U06gzsfdx315rGvqskmjBLs0Ti6RFSsjQOfSigDwyx8hPQaVX
wXddxXU7ciWFC2GiBh6Jlc0IP1C61/7BzqjYQgdv30cifeBUdI14qylbJDci4alDXQ/4ukg0+5OE
dM9FIf1xC9ViTe2sfh74lQElK4hwquheOPRm0UdEGwdyiVIPmDNanBLdvvYrlPuScYZV2A00FTpH
QiflS25J09ajRqYwI2CbxWIWj7bksiYq97ID9ObPaueOo6ZQLdqgZ4e3PZfCPFx1Z8nQI9G3smYj
CTdwRlt5tqhffDqNOGn4e5JJ5zJpVdmxPhwGNeKUrUQF548CtgfMmuZolq7nV3pTrX45l9m2Qbh0
qnYUEYmK7UPHc+omUreLddeQNo8AQq91hCkRM+NW0Dzleikqk6B8dUwAtC8UcsgeTPRxxsv1Gi7X
62f5+8idlZVDKKmSSzdOOyK3xO57fWu+iubngY822acrHNVXMd0OLabaosRDK+zusatFHJhD4SJr
39ycV5FVEkS8OnE+fTMOfO+90/vNW77VJ9x3K04bFXyYVX2bfUkeL5B6Kle7m0VuwZxk0mSmwjcR
JlKCWFKwX8xmApq6aGuX56WGIiUilUUFdMRz4pAXbGaRePkERaWgr4Q3hESCdwgJSuuRNSgIzBs6
Y3iZ+YrEI4chbNMMynvV7jN9fPGZzIAkuvMtrUS8n2c/ygo1M0psz3kNvzlVkiGKDr587sJxDbSi
HhMzr6bF2rzBZ9uIYrdMub5tMBqtTAX76Yb9EdFRUIXHoNOE/KXEZHtNj2C9NU5jan0dGEGgrLG+
kqvJ3DhCYL+aKKuxKHyAR15MwuMsOdr40kx8ILwc6WW6cs/uwSTxvQDSZMGY3PlpIMMhVUdw2mV4
1P9AfkC+kcVAAHAja+dF5FUJHT7UhCFBEnDSEeJf1Bd+y4SO7TGJjdCV3W9pURtxkDph4Kh+Oyhi
isvvNcA1hGY+gYl2ljDWMBkpG/oVCmm2AFh9fjCYZlx4NHCaaMlPNPhN+sZnBfEp5v4AQB0+FkEe
T4P+lJovxeWuxSaTpjYgpn1jAdg95QJAt/HECw9P5jTX1kFj8RfSAhvER4L4R1IbNZiZFdTCS9bW
DAbz2zz/MHkl9WdeYpMAzCuV+0rsRQTEGLx+jy6myjfZSI3GJi8/6J6xnzYNbKNwSkrGZQbjHgHy
9Mt7MgqD5RgToXQXgB/+8Re6UGwRe36suhOYWzHhJ9kil8JcNDFwenzqvexy8AK5G2QdvJUE0Tgp
FxnHANa96hKYgnSxDHjMpnxn14Xuu4HveoYClzvBrglknQBOePbr5SYxxhs9B8lQUGRqwenwvHk4
6e1pXT7sGTwjhrXz1/3uAFWf8QM/BYnylvf/Ni54RVnpymeCHrb5BFvf+0ST65DZDZ8O8Qz7SCJT
Rrpb9L7skLjgz16mfuiwCHEs+NQAzVi8vNgJPQ72K2Ie3SO9lDfoiqljYkXS1g1wF5gD2UDNVgCF
61ss3r+LYToVPXGhb8xXaPvZhzsefnB4+TBS/OtYjY2EbtweIGa+uhk0dPTGsqZK0a4YhxdJ5HNZ
5A0tAIjN85M1WgPt2Gv1JZ+jemW4fthnH4crSR/Jq/NGnHg0SIG8Y63Vv11h8snyTi2jN5rxMurH
6ixSGGpRCyufc0zWNDTyzYYIkjyhCWqPBHpKenyLl4MqvhOlaNuN9JYQI2z8wNT5kpRNTE16A4L+
AcRokXQq2BWS/KJ+Pyh0dXx0VoiwFSVBHEHmblzXuxntkleBopIZRYL88eme+urupRK+M3pc9/h1
u9Nv+/8J2Zl8oVhXXpBeIXNaeF+3looS+SZMaBLcjhdfw+5/h3bebryiTwY4eFIyFItlr/t/RKOZ
8hbX4ZcqqwSo4siZFH/zGfdwdvltxpS8N41fXIT9LZRYRmDwa+dGO+E+eN1iRpnKlomP/9R1j6tk
6NWXAPo3npHz/JI8TW3k59G6HJh6b3Hm8/MWoU9Yw/jl6nA7GZgUlnnGcQKmHbrqZtPoQE9rm95h
Uwdgbz5ljPbHHt1RCwmLLD5hp0hXM1AriY/dUgLZE5k9y8EukZ5TQznDRi96UreQNcP8NUIQmANx
ogLXnKcjkNyqrlWmqaEupcThYyoyp78jLskJBTMjMGWA4DNh2IbQsvmzOnEa6rNzS/44UCNZ5ia/
L44ERjn2nyZkhFi1SYfWFTrf7KOyBo7PmBqKV3EB8PU/xgnWCZI0386WY+7MoPFWh34hJXWJ3Fyt
ZRGp7DCTio8SDAMGRjszvRFhqTlp0ky5ezfTVXu/97b2xd9lPHrUItuVqujfwHBRpHoqPT1T6J2/
tJ3rnwCDiiP5gOVkPlQ+s+ABgCRtlMRNg8ykg3oYQKQRe1vTWqTBwlOCOjsocEr4QxNIk0XlMbHv
ykeaarSorvcFNKfb47585s4R3XXK2LWBTs8I7EcWO8WETrJK327T57In7ZwSUBu8gR/e1usbSnNo
VFmZ22mT5GebLp93aFl8cRUjD9SSsxYSwrbM/XxRWi7QWlkfrL0UGBzn3uX72QnToPqR+JK4xuDk
3w6EuU+qkfsC7UInEtSQooV9aoqCFJUaP7pfyLW36gTjSLaZ0doiCvxzPcSyk+qUyTRfz7bFKF/F
LpLE6lExjk3Mtac7QGkAUStwBH4tlHvHrLZgEk3leVCnS6IX2PNZS57bmf4sFB1e9mBhW9fHEEhd
EDnG8ab7szTj3D1TgXk3ZyNavYR7/BtxR5vUH/kbd7N11V1/F38r6JI7xNJmPID9qCUqQ0bMiHEV
R4TuRpso7mZgsbuX8gu96tbDQ8aUyVuJIQwB9ajwoPc0FjoTVi7QWBXXkzMxb1BQgfpRUkzfT4F4
vFgrpZDY2QpqoXa2i6V3ZYTw8JZPYDNM6axqVvNiGHtGxxB+wVACq4CncRRK/YhftrUVLgQyMVET
Xx8l7ulxxqLsp4bjCkFr1QBIH6JFD0hGYnO7HimI4sSgfTPW6hE1lpq8y2CJo0wGw+Gpi6p+9Ghk
np89F532VN0CRZ4epoxP+MjmoRmUIu1zcDaJExHwRc1I3pydSMuo/Idt+dcFIgixNLtpddkoPmeB
0yfSnIMOR8Z1jnzrfflNE/zujzVgCeCjU94kAOKylNzc8mAAuCVzgUQ8HnjhtufAv5USn7A4fF7n
8N8OuwJ/uk7s3Wb8FeawPKU44wmn/jB381ckMCvIXJCKIVZIRY/2bmUvhxn8UCWXywRA++Y5+ipF
Fr2UlaFrEjw9HIN5QPOHE+s5TfsluCnjIcVvszQRJt+U5x2eDlmX2lBatIm1N/odTaMkI0vf7yk5
zQqrlmRsHfG73xNn0gO1cHxIK4+C07oy+TRvzSCdZWwrj2R6iszRMmu0Wwa/XaKDLRF7N877aa9y
WgcEU0DhZs1InRrIGhBK8gpmVcV77V5Wkyjlu/+576ZvSPFWJyZIjV/BRsR1zrhzLcp0rKMHtwk0
QXO0XyZ9ullUnGHEZEv3FHLAjo65CZuTY7mBSgP/n4sl9oQNG7Vl/JiXIyDjFBwp6SXv4If+OqTU
s9HpLfcLlfJXDBBmT85ZDWdHIGG9FXgfEcR/v3ayjxMcmNZEXqWQlgy1jiykX3LMl2Xr/NeqnvVL
XqL0PjdDRTMSzrtxuV+3rDqjBZu1lYEdUNBIMxnf9IOcZIxdoc3q27771PBnHJ/sMRpXNc8GhKaO
syUIYMBP5LK3HsfS8CGZKmNQY/VYg53xpZmV664dSt43sXDIcuih88XpiGHMu+j5v0j2TeO4qucy
Mf8hpvZko0nrpLvZ3XGCXEAqA8T76iBosB1BMo2u/sMLUGCF6+6lm3icxc5weyBCjIhlv/MMRab9
cNQw/PyAUKFbZYklTxEPzy16T35grqW7ya61/mmHROmAFuxdIycce4m1OdKrrPiFy9VQeZJi4VcD
hVpBwewOhFOdWMZqK951DgTZfztV+7EKvwXqXaa083MIbRddcaIgRyx5U7QJ+tzsoBZj6jqZxTb5
YSG3v2a0VIah0YWK7JY1AWDq62K0IJJvk1AkTGF73U3U9xT2gBzj/iPZtpY92PMJf18qRa6fUXvr
K/scGzjlI8F99BB9QLfWfd5R4GyMhI7SLA84JS1kGNRadsyM8r41PPSvm1Ihrl5/n9yVtMQpMhmX
AyPQ9M01S2A9m1GCEHc7x02LaJtQmf8P8TYoGF+q+e/aTQmKmIKcY1UXrz9BGdVHFF9TmM/Ig+39
+zyW8ilEks+om0w4629XiIVSAcqHNLAuhZkdvPkswS0OJxCTjuKR843A1383NpFP5SDmFCXQzU3f
1Yaxeaj1AbIulKSJU2rc9Ajvs3eUrbyZlgIWNx20HlEPfKdwuvG1BelBEj5iPzcbjif/yM70CDHI
y+6AkQLYhJpdF6nV0za0CVFumY6GwxNHQh0f4R9oYiTsSqLTTjFZLXKBKal2kMyH140TgGbA50cS
Pr67ws/SM9MCNH1weP4BjHuMLoIkj8qCzEkcIiSLZCbLNEenIUW5wssKV9LkBTcxowYu9PtbYhCm
kHvtqflyu73dnDrf3wOHadf1RezAXP76OHavmOAJTt9BQpQispSpoaQT8bmwHtbEg/JS1GAxWUKs
xPFf0SJbyxrufnTpJ8j5tJNmLdxhMnVcCC2vZNXQQlRvFdPdnRWkIK2AUJ798Z+XM9W6xJ0C6ja1
8CUrgBGcoQ/7Y+wzOj3FlFMKn4ROZNx+ZTQONsB3eqVHvqKiNmTK1u9TTqUTvCe94eZwxQNaDGp5
t0pNF2sTF2APHmMwXPdleoitdAErdwYqdEsVG1jJmtPWk8uwhSuZMwstd2gUEkWy+2pzy/zrL8Rz
SD1JhtNwBzBBI+8o+bizHY5oicMcYKLpXzjJRmUv0hJiPHOS5bNHNE6KVaTyIVwwSqnK/RFJ66Vt
pbHXW2vht8lmrdhB9JjcCmcJ386iEt6gphluectBvJZswGDfM86KHcQ8nGBT8mRvSIJHpNccjOEA
a4Q/EqHb0UvrKDTxFVw+ehsFSE1SW/0/bvAycrc2KPUwwJkJIF8q7Ks8Vh76JrExbDIcXdZIzdol
Rca/hjslaOGz1M5rl6hxhtTUZ5boUvvnrHeZPkZrrzbXvrLV+aM3O+dTOWwO2XisZys5f+HaTPjG
Sav92QE9y2g7viBZnC32IY+dFENYAJNl7sZvZK5IUQWcgb4t//LZdO5tzGXL+W8wNON9OCdkrCls
ZC7Bre6rS0nvjTT3xJd7h3oAvc8QjxNjjMGSwB4ViUy8Ptxg10pInurDUT8U2YY05U62pMvbJrsH
xmN8/WJcSe20tx+CNa+suu1U6YlWIKhh0SewLoVWHWyCGLptsZnvQ893zK1UQzgNf1JEZN2U57cx
gHAksN57J69fi2JQ6UqnMvk6xZKCCMxOzr/911pa37LpXoO5pfw8kYUqT/Y8q631JiOWHqxybXil
n2VpCckTX5hnpchRkXqk2Kz5QJvnRIEzjn8iiozE8ttAykE1MGxcA3JRL//brPT39JLZYBJsQz7f
jROETYN6AI6XmZLNZht9JO0hMNjPRl4Ggmpx9Hy0ocAcQr+8IgJeZtFGxB0UGKdv1bjOrUXWDYve
VJ6LMuI7GwExP83+cGjmXacPzYsmw7EKXrnHXT6kqfGrqSzt2MYb0u4yGM11A3h7yl7W0qR0KiVz
wL9TigfjzF64CFMofHhJGc0jZVaC1QJXlbevKzBBJFCqiLtQOjbWlMf52Z+wsPARx9FqpcIl64rV
Qu4x1VPn8imlpvup5H0C8OQw/9hpSUzhUyezedaTxnN2AeQm317rOscFY/847DQs8GSdGgJYgmJk
7qDKvr2PKpK7cTm1NVrBO5WBp0OdxAuigxk9F3sLHVUTq94OdoeuhNG2kpLM+SFEtEpukSYuBCLS
pIFp9Ig9s8kougk6dJ/Big8MClE9w0/SLe6OVOglAjmbaq6VnsfhdnaYyVbwxREGX4bNqqHHFwz3
T5XPxR9wpYQAxKbf4ZhTNzn/sYzzoYViWYhYooXLBnf0BuqEAzN05wOE5I49eZ9FtbSJ6YU1p8ep
rQKXnKS1c8g6k6WJEjt69NAjoE30biRw8F7GXmemsEMjO/9G7erdj0E3oWoClsD1+cEuOYMRF5kK
b3aazP9K5oSD6zET+KEK8X4OBB4eu4YcjM0UqiYxvD9V23fZZ9DgMmzx6iXfgq1a1bvunmM5Vrko
RT1H/QfIrq3Z3E7we215dSGwSvsQIaC7kXz+oczDZZ9BE7aBqapc6IPVD3Gj9YjQiZgSowuWDewN
zSJ1ahHKIw6yezyjvn+DT4EKMOHGc5lrGdtoQ++80z/SRwfH/gmd9aWh63kF70EXkI/FC/GZe0nC
HBrqcSRpXVvKCLhOAauytG3pbJlMjo4wXDEmZEop6T0EsOsi3M5gvmu6mfxSxxo/vsguL5tGYXJH
1LzhdzAqqyuz/GEdTaTm4pmywtb7kXVuEXZ+HlK+gLsC2c/yrITW5Not9LDJIKjgvR1Ir8XQQjl3
qqC2XA1i0sZZdAHOFdYBZu5eGyF495yHAF25W6MkQYJDDLhgB7MQqoFNuhA7kI9PIszpi86r8y5L
ow5A9gf5hhioFgzRmIISUVLkd/4uXiVCZKEdogA6/SC/mz6ibV0+WpUwHIE4T1mG5KKTgr7kK7Y+
DTZgotyCOeh8rJ3E4PnO6EDU9QWvR7NOsOL90jQpm/nXsuL80/h1V4mNSzm4U4A5X7UtJ1WguArv
ZpZJQSYK1x9SBStidCPwb1mgWDaPVa8CWoauz5sPYlk4TdYumC8lEqTSUC1nkHsxzlqVgwQvr4pe
Fy5S7yjmiJwBTfNJx6W5LMfyacke+gxkn97nWtzwet/L8c2/AQO0hTJ4U8odgYGCfS9BanqZRYLG
BTwB/r+boArcVrQBqTKrPsaDefYTTVlnsO14OnZXt09icy9pXw54WYlC1yx83VPdxeF0wSnxPZsx
ERZbOFIQyQOdX3GaRGkZGTwZdnzZxFUWlrHfyX5PCzpx8UvBxOZTt14Or8dNxTsev64+GIRKEryh
0nbkb1ULnJYVcgiBKFw4hefzHTI//lAfQytRy5sa7SNvpCNoIVCDnb2Oh+DYNzyFH7NKFn1raVN8
uEfxKXC1z3m0v+7+icuMYRL1UFSNHPmgVjxpuMaR5Vdl2IdBXvCuW4/nncJ3IkLPiXodWR4R+iAZ
Ajb5iX2hc/BspZm2l6ly/iF24OWp76tOG1UxhNTwWKi6StVXSpHN2ozYbsIPtnkewSpkyW1RnOm8
OZhJdYl1KCSZExbSfbndKc6rH9moPmQppIAFr+4elTnCiMvKnUKtbLGcrCE0YsHfOwSpbT964yfk
cY3klikAGU9YpGbP6RE1H2UoaHVbFFLdU6n5ILikKerRLRzU7rKvsiNLHcqpdz92QMsH06WfH7IT
oe1XCKKZTWmhp4PQkqmmFiuZjvG64JeVSf9mQnqPs9yz8aGwRGJIO8uOs7YmJTyNExZuzvmZANDD
GzJYutzR/B1AitdN60XjkoYV5V1pdcr+wfQkLYrK9jSDFU3NSHcsufZlDy2HxPeTGfXbWxmgVibF
G62jklFlHroY5qhaI3URmm1QRdrLQsNdDT2qq5A3kYpLFgkJUmhYI3lCqQHWoheqpXGJe2Az+ALz
qN5vVhRPGZ36MxsmvIfShrjBZKE37D6SHzi1ky257sATcRZwa0rvyrmFUhNNFQ8Nz9fXpPvcPOVc
gJLQCfJfSUiuGdBJJeYzrBD21cchmkTtRfaG6H7fo1cNjF05olNX9rG5lbSn/paX40a/a/Wcc4N1
iowK0DC6d6Z2ZH4nrDD+ZbPemmDcH1XcJhN6Ft9JmVpxhlq3n5bwj1J3udosTE/Lj78M7EFOftFL
tPSRA4JPWueinvOWyASpFDDMWPB4+g2sPs/HDqoRVPv+s7eXIPhrkfOppbtuop5An/KS/sYwdjpY
3a26fMtEdRa+LK1RnajqGmwQL1kMnQcXHxmtT+8o7YkRJs7MVmjCcKZgkTJbpWG+WgnThtDt1nGq
Qn7aBdnVoBF+GKmyl3W61YHmf7eGyjKIEdYgmGUnk7bc/rG2clvIldHJZzmew/I0t1boSYGDSMBD
7yLWT0KtpU8Y0CE5Q7qIKm8HmrQP5ci6O9WY1Uu1N4hSpN1kfit9AO6lNz9i+dyE1r6A8sqSYz+g
t3IW+z5QMG4JzAd1ib2AmU5lhvUnUiLLAkz6o/Ocp8VwPNgL+we6YpthGsfilkTseZ/b9GDgm6p8
+ijcj1LtLgNAwhoMNsld/R3Krt6Lfn1nbvNd5wVbnrWXov2WGAW+wjcaOuBesNjfr05oybompNTU
K6oL9B2GaHoobcFFbEvHs2HsjyBF/gSpYDxYtI5rnUVrZ8N72HiBM8EwhKSybhXR+epgGZOedH8B
SLT/DGYXUYypZzDO3sEro7mhg0dzZSrSYAEZZDKnhaebwnKQ1hlLsBwk9U1a0pZs0sc/Gs1jTNW4
eGwgwwZwxxsJzvW04QeoNjF/5tRRzCJunv+OgVQ4Crf4FRsd7zj/KjGMVOlT1WmbANYe4HAg+c/F
MzdXTk+qJHPAqao5TYqbtsONrTt/sqIEIfjlWXvGC9eSyWKACqZ30k/xKk5Ci94rq3llN3Ja1WbD
Y7nX+sxL7oj9gR/f43B7bWiAE0CuIsf2NZ6uTpzWKPMb8SPog5iAQboibeCgC1MvxHIZxGN60JLw
chatxHxbnhN06FDgYYTAxvI+7MLvFaUl1z/39Otjhjq1JJB6lfSyWzK3aFCKRZY2VBct8DJ100Dq
DRaG/F7CBXYBmtHpg1BSyXexDDUsEdPXTatwuXs36agIgksrRNP5AJBH7GAIXrAy4SUjnlQwdVrx
HMZO+9gmDpyRhfTDJi8rGSq6E8/mnT3n1qAgFIYrG664YyhfyBb1oesqh9KtCem2cFJtDDi8xghq
FVl3AUvi6DjuZ0UrTmsmTzGUazx/JVs1ilLRp50ZMQuJqAcAio5XvYaR4UelwmS7Qre8xDHncTYJ
YthaQIvepLPXQzFl6Nvf0NyjXxLCSJM6JZLVkrw1tBlRj2nuT9hRKUc5zU+LVkLGEsGwdp45HqBz
wYL1zScPi+wKleJi8WnvFV7VWWfZdu36/NeYahHzjnHU9haIQFNtPKqDiBeWhI6zGm2csZBCtf6J
3uMrTau2y5z5aXn/dSax30J/7i6ISWK+dhkFRnmfL3JUtYA+c7PUtC2J2XweQilmnS/C0hFd7E2I
LAdWlp4lEz/GY3hK5aPqEB6wM2avzKS3hbXmI8ESX8C1JIfFWpOBjsQlbh4rhouemA0a+rm/qYpr
LmXjyRDYd4aaINLHBWsieCIoQ671W6HIXC7TBzpvaBF+BAy9/uEvgQSHt2BTa44Wo6keIO7risEE
PSF0nO97bwnv72aaR6ZT7TbjekdmzkTN6JaHYcQrOWmhWlSOWcfkFaDeg1eS/+wHcdZ6q814fZBU
0NdeChr7H3O+FcUVdxsB+6eQaarpvYSCDg5B6gl3sOyqNoWU9rnSBOIn6854YNOcCih0WvaCZ+s0
2A9fB9sIujsHW5wSSf19bmUd/00tntMgGwZIJHe7RA9QGLUwE1fNT9yS2QLyIw5rgT3RT68bzTxp
4DvUjxSz2V/rQnXThK0zkqPmBhwDFjnzotUG5E1zUUyjq3r+ltb7JU+280KR/9eBDL2PBWE22OUI
RzBWGAO2k6nL7+fQGc9F7WqsxT+LNdNnQ/xt7v8G966gbeUQfgiHDbCS7VaIkKE7a7QfNtBQxMIl
AQm8TBJHyV026Dn2StwHFWt/60Nl1p61a2dwPGeBQensoEceGT4mSMBASmQW70NcVUWGMjFSvbd1
GNy5TPvdgnhQLdE1Hl2bnFjT6AOI2LEDGKU84+i4bw9GjZ87ZninDSQdRlOjstBq3f+tFdCU1RjR
a82v67sQ/KMbN44kLvaIXCxuTKDGTu3kwdxNZq2FSuxhOvBOZ/EJy5JwW6yo40DQBbSzAFZ//ACc
ID8h+XHKZwOE8L5/OuKmqIIFyuYbpbUp5snPCqJIO4VdGx1VPaM+1KWpYYieTqxBdkioMM+1QVxX
1M3ch/S6UU54L7/rHCpwliwmkWulMw00s/1LbR7/02WDEbYHhZc/zQ09DGeTGBIZX4iQ24pMiQYk
zw3A/ky4+W6yD93sGHUe2YLVm0hpCzfDzduWWsy4CllJevnEzB4qJaDGNyQe/Q+i0JeXGGLsCdv+
nwcJVnI+fJUWXLQbwSeC8Kq6NUCUYal9BIx22fa5y0YpKm/IZ+CUlXuYpwwSr3xVH4kL/Yiz16Ky
YEJrK7+Z4K84PjGp3EySVhJC1XFSCEDEW3AyEVi9XuJhaQ7lTXTF64Eh2VBhbZAzXeTf2M5AgSYQ
FQfKMtcUOOS44UfaYrS53BsCsP2ek7eTcnyqNhRMTC4AQKWYCyN3ALyGT/d1EZqBAxglDOLCDKHV
sRrpfmGRobkVLJxPqRTyL927JdQ23v1ZAvjQZiyEkt6gI0YWM/X1Mp58EZpmO67imgupGlfHcZKp
DdrpU8+gfCXBlwQ2LMPHceYBb0g/nxyvBk6DSV4zSnPmvmCsLeOEyMU1x2wUQkdWW9JLDCCUJmha
X07O83HoqphU6v1Bj6+1a+D7jllYUMCD/D/bD/NtdIxpLT/2GYaSGdfr1glDb4lzqbbjqRiShSeX
MXV6V+KsDXVSPhgAerbNdQpSNmhjT1ulj8d5NTo65JPuq3wvpBiTeDYTyeuCeowurFNBcUWyrdiM
cvkY/GSiGKv2Ij+vwwKPFwRGOsyQvMOBfM77aBoNVwIhBAqsE8ahI9YXfcOaPDPqTZuoyf/lXQro
NVxJbsB8KHg82lLdhYWQZ2VWY8WRkaDGQA7h6STzmps7BhXDZaEBnsOqvLObSIAuMaScCNd+S9p6
G79dledrFuOMVd6oAI8VCZdQUpYhDWc1xIPu+a5WP9GdAEl2hR/hoY7aJ4H2q/O3peoA+k5VIpCC
hCFGUQhHsyVGEf9m4tdwvg1a2sn73p011yPy1T9QgTPQjQgn70dJSuXqv8unCcsnUOwlbBksAk40
J9aHCREcnhqTTIT/AA29u2SbUQ/+xHs8iP6miyvcN+8SHJ8PvPUyX4zgPZH/nvlOudA1zYMDSnqm
oFp8YGgPplZeY7ZWtXRiaKN4OpvXg/Ro1ToYo/00mG89O5cpao4u583FCsHViUqHgWJd8wgZbOb/
rfn609YjxSL1snX8nEoDfEWB8OyqVPoFm7kkuDsO20VV1f4/IHr8rP3ViB37NAgxgCvkh4o4Qd3v
qe7EKB05CnGLWhNxX3ujoAHlTLUpPA8VCXFXahAUn5mnE87Dcvc2H9npqhbOlzQ5MegQWgWIdh8u
UnRBgvxeNO1Ww+np5CLNLR0yL7Esv17Bilwmbkn1ABUuDwg9oFYCLKvZ8KAbC+A8X4cWNxWkLOs0
8Yc27cSRRS5iHYcyB2vAqog4yNqjN+CtE2gd/VXDuMpBdhToZ625325i+mqgxwOtGY7vm9gm57MO
mbqPzI3Y7C26M79RTPCxY2Z93gWSc4PTBoOsvPs70aCaplKkgsGN/KmaSEEI2Eq9SLNMgCTUW5wJ
0CBm6sFFAnDerhN943kTsmbRBfzBzYR7yeXvu3aizKaSFthk30BgQKcgapsL8IM0A4oHcYoGxgRN
4+v/hkKBHuChgvSFj2JrYrBIQguk3dNDJCg1v3XrbXkqElp+PX0d8fGEAx4OgweXjTF3jbkkgml2
5ryefXgmjYvvgL0dZWPm39aQ/bDe8gVnxGYi6WtYrStFhtS1YhU1QYmnBiN8Fi9pSNVqv7DBaIrs
3As61+yNZxFmaGvat2FcvlTvbNmA7r05FppWbgjY4JuNFG1zgY5RyAD+Ih4rsy/F6sfhlvAbb+y8
9h/BX9gso8CS3sne3VJfgCzq5WtLN9Bq+/fSUNzdzexV81POTmmnD/DclpALcbA0Gtsac/D9XQXw
ac787lrV0/jwnzrotiZW5mOOsNCuUoFpBehAV0W3cREUjiyhUgSjsV9ycEe7SzsM41ijIIoZG86z
ZVFx7dj4pBDToIokyvyQRLZYPKKkUsQFRG+42h6hF1MScZcC0x3PzY+21stEX80fp4t5UdzOJqhT
m0FMfSA0utrpB4Ef2dLU2O+RqLOozlxV25biUw16+utoqOLqtNMIemkv8cz3Ht6r/sLwv6OfT6YY
Pd1EODhv1hagINq0/FF5bHwI8EM91PA/Uaz6Gr3fNiSrlMQfLFgmnc/PkC2UBzqr6PJvQZiwdtcx
zFdLEScm0x4cEfRM0YapV/U+XjV7R46AMsDs1WA61AYhvPhdpRwLqQZCpRvgfXdwJ9f0aUpwJlHo
dAeSlbhS39uqwxlgWy2rpSiRqzw9Go0GNbuW6S2bZs+B/WYO6FyLAje+jFkb52LXwpXn5LzjO/w5
QAF/q0yJ7Okj+MwS4bv6aiunOI3h5jifVLUmKTVfDAFXkvyWgYudrrFL/cR0YMOb6iODgjExXY5S
fvn+gXXoxoj3tlY5jJdaJ+XMXIIMqRsaRBD0tzdJepDMfKWofAoZYs4jOTj+fCA64v14eYr+zJS5
nUs/ZcdsVgJp+lex6PByYBfSsJWgfsKj1FGjyXuF230Wm2NK8uIWlmN2jgDsBPPy+TuxkbAwbGsV
ZY4M5R6TXRIGHeDj5Vv0nfyNnPl1YB6ckYzl451bSE47F44icpmdc+gwIVvmGTgki8EBZ3Z9Jdgl
HOuJXbnKEPKy0PEYq6hsgbibhblmCCd2+NftefXYjcku9hH4Ado6WnhywDia9ikYDJTPxK8JHfpJ
deYOuA0srJU09UMiyGa0R4BobY9qa56w9/cZPaIPmcsVKXTOfQif9mX5vnhk5Hv9SWRea0b7xzDT
VuamPx5Tla6JDKbffCdV6UNE9n+2PeeYyCa6aeTGzXudPfMR9KgJupspL194GYK8vJCCQ6AZDpU3
FJ+F29WZ0RSPWaZZCundeZi2zatpqJL31z7N9msgeCYgd78pOrAGWtiLN2i2Zcop8JLoFbo0lrwy
wLABygBQlJR/2OkZvDrTGInXd2eDKSZHrsSYu9z54UjKOm4YwRGQ5sct/rvmPZ7fo6EYSjrvHAka
pctVkpcmcDvKyPZP1zC6kRxGnJEfAL15fB+a0flHfEFQaDZMe5sX+bfTiPIlM92NKtvNSF7SFU3M
a45m0q6LncR1rxNAqSIX5SRn/7r2bhCRAsU3ASVmjJXOpQoRyQGMVF4EZ/uXAumewB30ILZAhf6f
1o8lBBGOeUgMjGOYAGdHhQLs8gjtUhYeTJ7abu5pTw9LDdtE/hEgYVhPcAO8cGkLk4eD9O0CgYhV
FsxZb06WXU9zZEVyEzN1bRue0AT/llwUbe9dxPnaViqEau4Yf1Hpc1iDyMRwfUTXtZOfHxVeHt/6
ib03X9yDkcp23Laz+LucFZuXCNYofnB5fcUmKj8Q14EqBZUV2NHvNUMWJsFGHY1gqrvnnl0qGGX9
0oAq90P0Jrbm24NTP5f9hgPn4TtPD+bSx+VPVsz52rDx5/R98wQcGcoww+zKGJpNttklXvc5G0mu
DKZEQz7jucZzhSw259uWKQxF16fA+Vo9odppOvAAQ6aFTo+MZ7C/e9JaHd3jbDtDwfb6ElItbVf+
MD4jf7LWj7e7YdrqdyuGaLlHYzV6zPB1C+Bu/Gun3YrmyIFpTwmxOmjku7xDc7MuGEpWiVqiVmNg
/5Il+J/c4k7M/GLni19349vKVffMD9XDcTIEknBG24RmIxWsSb1dw4jqzctHNJXGSvR1qjiL+TbZ
6z5aTkUuMbtX5MQoTorzPN8PhMNDRXLsuvCj1Pzh4ZfVqdz4gSQdeLwYDZwt8gl6iZMYvdntGRMC
fHbaVj4yWxRraYXddhuLhRpXOnAP+AWTHVpw2OyvGtMybfeuJrp8Uxq0LQaBfCny+OWH9Znu7xo2
a266faLvL+e1XeKj0gxsS+eqzB+rWSVIPNBUYk0UVjBfhAxa+/VMkBsQEMEif2DrLOwiLSmo5SoA
LZI2g4plmuzUfLyD4jYxi7eqVKSwNthOhATtIga6x33Mnzb+VYOZp3CR3pABaviLQGbHkQhaVF/8
CFEkfV065gfnmqeFP9PKePAAByqoTRV2s5vSaON9UyLC/oKU4myDo2uwjiY1SmK4tgdYKDqZeGUj
zNvvr3sfCwZOc5w2b7aAGzsHm+IOzBxhoMgcD1aBFY2GrEVxCk65nJ3ebNtWoGvjCG9fjsxcaqDf
o9DC9jYu62pMfwl6poWmvcsy1n07A1k/Um/WxRhZvruDriYciHWr/9sPIHW4b6Ifi4Xfox4jbNfn
mhBEovkZUYmPgdSSqYVLOZe0q/n+p0Jxg6Tsai3dq1X7vK6n/kDr8lgyFKPKHJxT41Gubqwwy2v0
6z8Ys3PRnUwo+vIL2TGwfbn3+RdxO8awMVcbrCwbgxRh6aeJlTNmKwOUg8n/WM/b0pnrji4/jyLg
xRrQlNSfFvgpW7/m+3vOXCCMeNcOJZ+KMJMWXJqO7QE6Ytb9iKYtEeyR6UZgHBk98a2LB7WLLCB/
SifNFQ1JiV9GHrAhhsU9NLgJjBhepKGLXAtTgyrHyyZixMMbSGs+TLIFYcs1ttKZQugnha4E+mmG
a5UsfdLQ03cSMmd4iH8KTVkSgU4E9+TVUBkaFAHCYOXcPPLNwK03zO1d9OK6qulGTa6TWPU+3URO
4xN7b0rxGnLmWHNAHMlI4pLymyyf3nsy6AM4ERgFoAs1zAPZzbZYtpeQcJsPVJOYkBPctSP8C0Ow
91IhPz4vbKVhJzeSD5BPa75c5EWkPPW9qgp9Qs7kPTfqeM6N47jFISQ3hnTwnBW5ELiPqrLwjVLk
bHOLLrnx0H50xdNIDHHtOhcp0UEO1POhe1NW1/XTb86w5OG9b7dppK0WMdKWjVLc6Z4xmcMMpvgX
Wl0dHrnTCJ0WEkKBQ1f+h6hR/h284kAJauas0L9KuiBYLlIJY4lbvKPE7GJOSGSfUUxb7EZX+mca
AzvRvH6nBnCDG0w1GzbODNm0PPB9i0J1s8dvvYYmIsHLJAgbC0ThEmGRY6GzKGepKNbElqOjbeUG
C1dtvBpMdUwPd7R46lLrzDKRPm3hd5Pcv51bX2mC6XFddR0F5nPg/BHMUW6ayOFE0hM7YHdis4WN
qTHjW4Uk1LBT35W8hV3r4MgY/xE2ZzNnYy/rWzmnB77PtXeegUQ7DF8iZLbhg6FrRJ95qcgt9dRg
fjWuRcma670BYbglSXwHUetVdApCtFwJtCUOGMuNY0W12+zve9ATX4VcjGcJ8DvfrB1aN6kEdvmC
4Fis1H7HZ1a1TRbLfw610i+tv58s65dVgyM9D3G1ha37izEpVPFPG/XJ8RUF5YGwTazaavaO6GjD
ZjcwENX2vMXyzTuU14deAkhUJudPAeT9MIJkxNqNHdix1f0oklNWPe13Ov/ZZvZSaSuwTiu9ZiPo
7wiIBqPbQI2El9u/W9Z9RSbjiJrBl+Z+17866KCP4Rz5hNsjrFSFlCkj5FEi/dqFvh3Z17gUw99f
ZOyUa2Vc+r0BTIIJ2bZ/wY1r70uc2a0r+GTnSwyX40ZrLxT5+ouSF/ZyG++mhV610jc4RIN6FxjM
37WWxHMIOYdBxoPUmZNMLnWPOxL+k6iT4mQBwpTiZ3zolDd7N6Y/taSaKNVfZ/Oypp61iXJlzPOK
GasVb3QTs0deSV5N4BqAom/drj9Iard3EDxDTnRiDp0rxbkefVnsJ/mDk08CAzRED6dDOk50vl1+
/GoYhoxr/zmDjFlyW39Hmu+9cpGvDog4whwgMiOv7+Wse+7M9MNyM6LUduUX8BRldhjZfaBoz4ja
+F2ZAd81xidib+UB2SpDs54bZaLlK6k7fIsAJe4V8FA2rAtJPy12WZ5O6Im2NAEVBNXDv8Y4grTt
qpw7C5I9ohiT31PC8TvoJUzPijtM2LIKXdsdug/nEd9dI+cPSzPJ5CmBHd83AIThq5q2l4tvGP9o
tJxL/DrOIeJwIiDSYqBNj5hJFBpZDxfXGYKrF51TP2jNqOXtzZJX42/U8j6vD7SAeIpfAohb3Hhq
Jh8xUAsF/iWRKQM4QhexdeOJo8LlMcQCm786JrJ3cIi85OsWmRcm1dt+tRLnbnh4D7jMNxbnF5uB
vqbvGp0HPrgmhAeJKi7lpTl59Bw0ogMqEGFBaEndiOhqhp7DNBQxx1eDRHl0STON1p1SmZn3kayA
VkF/k+1mIOR+qOOUwIocuS5yh9eUw/nVL8qhUwt4J3tUwu7kyX1ZLSfUh3XOsjet+6OU3OMhXPKp
E8F1iZzYq6j+1T7laRyPaFaA+ZTV7G+JNO2PO4TUwxxVmhd78FqAr7s2sjpsTC8DfNkGBzo9j69Y
bTSIRvJBdfkAd+pEB3WFj57xJj3NKf8270T6lG7MIC/GkwV2L52qaOqoQiqScR4IQOHfYz2cQWk/
4+Rf4NxBSacwBVvs7VGXiCe0FQWnzGoqfdhNcv1aaKxHzk6CvU9Nch1On0ypKZ5hf5X1MK5rLb6+
NN7Dkby1kl4TS7WHP8NeboxtaXXIDEAY9wS8OcThhDWWChBpZRjXXMI1ap2gv0dfIJCVzfAufzDq
j4XcAhHC5q/yhBOVb1ZsLc++jrA04L2gJ+r6OuLPmZQlVr9bFaO+oHHQ3Ry8umsUtmE3ov0FiLNr
RUYktz+UOYB5oC8lRgNsRQkhuGzE2WFqB2Xu849BOyJpBcd8jFiIt8YwKQS9bhvy96ZzjHR7v5Xu
45akPHlopKiv329YFKDMnQsFnjLNT4ZFCDxytWd2hCunqJBIFZhSajRQY/98C4TZR2/ALOWw5GSD
m7ZPDxFKooDKxH+WakiaxDkNqfqA2eMz2SptGuGhsw7rlasnfv3E3Hkv2OIaytQWMIJiDIYlTtvR
F9/fykVBccfunPIkWIwiN7lfQeU0+/vBsQUaMX5Synfo6qwRHaSwn4Nc9D/GkPOw0EmMdd7NtKBP
sxEGelpaF5zOLxKNrqjHvEhNNSwc50zQcE9B5O/U+IXpoPMXTUjPcrK0X5D6SJWtOPS8xDjyA49t
e8+CoMmE8osi8GPTz0aCQ/cwQa7Mq3fLW3fXfwWsOUO2qxxdNVvUX4RfhqADlJ3FxCwDm4s5JHDB
I6GpNjSWWrWwf6IGZOpOFK9CNUKb1/tu/ARkZjWHF9Ega2AoGiYPPC4P99/b8paDp1T6boUqQ1FQ
5pWXEboJ4WcZ0jMUsdLVfqH7WXK/LEmrTzD8hSff4yeMw+FCXUo5np5iTbLJrL/Xg2X7sDHwOy7b
W33uvlVlxB0YLf8FouBwMn67clu0rGw70VvxlTrLHomUggeS5H6uiXMlkjgOzdJr9SQUKvaKEHSw
0JjhOyvG5ytbxAakX0bjtzsd53T1oqeWfc9PGHTpLzmBH3LdA5IqrVJhMqBZO2PkRQEaCJHGGJKy
5Gq8ACb6n6kyDviNxJxwCP8ejf54Cn+T2jHEdmAGVEiM92WNkhnz4sYEfJtm1bWa+zyMnXTOUB6h
3c7GH3BuTJvXndH7qh2S6DTjdCAZff4zjKg5hfyLM0CUEvNa4PdddYbcvOiZ5UkpdmSvIOQNc42j
UzXSlpt5by2ua9A8WSTew47Ngv2w8hDwvOKpRg6kxZ+nX7jOO3HYAOUh/vCobndkb1AKlp05L0ZQ
Am5yr5rTv1xw9uxF2cG71INkxb9HGpo7DM6cMktuIrsUt5Y5FaQ96Fn1LLexpjt7Vl2x5s10M/0D
0IwiRQj0bcpf3+dt1NGq+LDF8laZMMlyxV5/UnhcfnmD1OMULhs9pNaeDSi9F6lndijKeVnvhrjG
ax53b14hPwXMCrEXpQYegGPFzh+aFOw/6fZB8PIlBhoRdpdsQIyebCtjQ9imJPnIS0c6TsX+GRMF
f29OaLsPylXlVlURy/xmuKScOC8NW7jYSzkM+DuRpisTP68R7hdAHQkgG9dRywbSviiZ+rb+vYqS
01UaJ+ddgZQlE6tFRKDQRNkfAVrrZ4YMeiY3rdP1cn587hEH///n0y6QmeVgebaF2l5dyoGIgsO8
Hner8N67XEYHzdEAdWUfFUYVYrAGtZxSIreHjmelFCwLFqXc00VObAqXJ90K/8WpfhrjnDikLANr
h/rhbewvYZmZDp9Vid0e4LpV60dUo8zSwRaVh9C2knbaaR2GuSW5cx/NY0QnyepJjANYLTDTeuO3
GpKCm/vUxBbtfyF+CuLs27KdBoF/kq676WPR0kSi1tCeV92ZbG5IJibecnBK49q1UjPR7SmmqwQu
6bNx5o2fPLDrP+rwnYuT06PcmMbOJbjawt/lIPmZ1D0gfrit/Q+InCBvgdrpexMONL52Eb1WKoEI
PwVNFunj1hif5okrsyGs9vzKudFLjoX8xO1UkHH+PUoY/chqKhFRoT7Gdbp4YZXV2TY6T2nuUDoJ
+A8KJSq5zSUSfYeKhSWQMams2wwCXrIf6NvkEuq+QyDO1ME1lm0ub6ugpebwyjLklwSaSq3D+y10
p35TXmTX6xbKI9sqw6+ubhsVgWkNBdN+pO1b3Iket70h/OwSYZnj7rwNSb6Bchi/kYTmpysRDU0L
7w/uxzUFCXSyQ08paeZgZRArTA6ZckAeE/dstXl4IanApxkKMt28omJd3VLQjYtXzAIc2ESLhFiu
Tsvic6YFEDGL/IlOiQu97ya2SLkXFDsG18dkPZa4clYX/8Po89WvvhzqKvLc1tAs36cUJAL7zZdN
bn3Puku7UH5ljxy0YyBgyXNb8JecYg23GYTaTjqRmIAbdjdt1kioFNgVWBtkmIpeaufO54L3rh+H
8548K4qVoQkwXDNirZlVhsE9D4QD+bzgA5vn8xUIkx2BOJLmgeADcljvOR+fGzcxm6aI1639azRM
cZzHeDIsH0GQZof4gAIsPVe5SxellIBMmcWyGUEnoX6KivQeGqBlI7uxTNQS++fm2vuuhThDI5Jg
qf7KrrYbOF8FJDOuUZa11ttYU44cCi0bhQz3hJwTVRt4r38rDbx9x9DtHmxpRAzGCL14xGQWs95a
hCMg4o22Bi55gcQqV0nfrmsxRVRjlDMfCpSCh6CViCbrCbZcEQMZ4bFM6y3YHJ4wGJgPKHj/9TWt
9HyRWOSnwmPVDU23da2bpgJsdnLIHMvm87akhczSOYtMCdHF3RjKKKtN1MlUachrNPXgTSY/Rj3X
zsV0ios4ujMOUIe+oTm53gOxoe9ClmYH1uf6hAaWoyPjB9kQ+JPY40F/plU2rBWcd3sT8uE4kQIi
PSZxp+Gsrc/x46gFGlZLegpciF/aED4usC3qKTU6m0jqyLM8s+mOFxazbC2oZi0PPze7gnkSm4xC
TtbcK3JHoXnm/sHtKuGGrgFXXnqwWLns6IZ2cWVYW+NYfEqhW7fE4hE5dBGOVG1muJkJVabfyEbK
wsPP9sybqgTDdP9GtS+nulvN/+wyPwuAqCRiIMyg7to0lvY0g4zBxri9v21Ohc4Lt6yqeGWIXc8G
zg+An1FmtyLBYqUiFud0+FvTjbeBQvVi2pOp8ELovPGXeRImacDv4XLldF3NDojrmTQQCwnuFb6R
GXkOQFd1ude+kWc91rVI26pgNUIx68nEvpvc9Rsd9ofxeSemGLNtEuNpg7V4dGiRfIfjtM22qGIi
ifIp3OJ1mMaeZZaMDkRr7XTn++wAgl8l7WPmhz5UyqvuduKYTVzKDNmOSSLnPhJYtiyQNW5ZREEF
elsY7OCKci1jYfBLXrwcQE+Z+bIbkhdcULEemvnjCwVVUFcvtupk5sAszqYcP8GxZZGtYC4nyjPL
+RI3mPNzCDmIOoRyKJ/Qh0WTPLaf/Em3csNHXCPxiGOuV87COkx7AHWceCErSBazS5Fn62EFTzmr
DMSVq9ChRuE/OeSsthoyy9SsTLF9cAGZMxr3MCZ39HFlhanN1tUMF79G1YElASTPs4TwCH0LkKVJ
Qy81DTEmIloD/461BPfAUBrOdYcU1G1cm1/KEZwzTFhHgfXLz86EXmbizpIE4fF8JHq6UbELzPss
PL0mAWHuSi2GzJb/DVR/zMyAKV/2y+LlUeLt3nsINrVkZ1ZHHwNYHl6k7oKQRVTLPpMx8DEVwnXi
FdEO6LLAjJFOX/sleVbaJVovo6hNp67b7kdUTZyfwdXP21/r2CuKkWxH105DXejtmU99yBgO5Nag
oYp+tlS08ofERXxS4JJjZsfqbk3o26k/xpIoLR7Pu7UmnCFbvGUR+CIkbf56wbCiwTdEGneQygcb
Gr7R3fjKuvv4jZUnWbFhWwwg7/DpkMoq+IqDmuhCWKHBnCw/IQoAAN1WbEr/2Xwnzf/wvo2FaxQK
yqoyMI0lxNiEDEoZE6yxp3DnBvjCUT7B/tcLwrvLWj/DKR1ycp/KYHl4coE16mHatQCxMuL27j/3
iE6sWby9jds1X+R54Wbrw/6j4gvsSkKTDEFc3GJofLHPzSMr9sWhlbmAt1kcL2DnCAIxnHbFUVWg
9c3MhhEWfM8zfdrZ52Xl4erxZpAtXn7uOJ1jcETY4yOylXQTH8nUNziGmwmfzdoZQvJbOaUgtUBK
FgJZvTKf75tN1RqH2VEoXArOzsq3Y22u6T6NsVJSKlnJcS5PD5BL9MOtcTHoKEV2CxZgwj4OtLOv
QWG81c6+ZSjfkMExmwJK3mQQi1LE/7Hu+XR1ZLS4C7OuTNbnwXrfQfxSZWrzJpclAZhwvy5euCg4
tBmMGyjJYAyWfecIHc+C3s5CyaqZgn7zMqR7gEdLfXzBGTQO8YcqoTGTgCuK66AItCmLUrhHQmOB
ty82jnCR8nwCOdZM5/1zBT0YTIkss0cpilY4tQfv/x5kNE1bk+M5AJxnOlhXsiT8/4l9LkSp9c0f
hqkOqB0AkwafhAcMEn37IVCl/L5KJ1XgIDTVcTWEoWFLED1VArmHbFxIqY406so5vHEQPxx1sE+U
DK2FEIOAeP11lHrARxY1+yl8TSmJ9VE76Ke0GOJQ2md78QPpny07u3ppGM2+RPMaGaUSX7KTsubx
7sGBySKsRtjZQNAc/cdMZxGNoorH2agq9RYfiC1SKBOZAko+KdjcbudOroMzUuDgaf5FMJN5I67D
AyRF0kRBEJP4pSBWScDuplrTKUYaDsxgZK1OhyU1fgKKr75TzvbUt7qVPk1Sur69y10DsDs6X7yW
+dHqGzQljCMx3BFW7gCHogj8/d0fSzDAuOybR3SHA2gjXuBZWSHUbdDySWQ/OXCLh+jk4mWhuwuX
7PnOK+1/WMuy7kf4BGBLC6WdTrGQEeeUraeUfuNAeeIps/RXUWboYEDIa7DQtrFXCLlPxp/vey9J
1Jke0JD4Cnm9M1a78Vb1x90z02gWAQk5z5SQNo0nB0VGi6Vca2adPB416D8tU3lj8eo+pRV5ncaY
dL+2n8QztiOFDIf16gEYUul1yRDQ5XPqR4H716nl3XDcyd/DfAhDx7Dss+kDw0jQ2rnerL8gzfg3
EdTiw6msu4D9wVbVhMHhMxSUDkNU1koScTx36nhUbDqsZvxjiK3zAmeNOhMJ73lOJR703Pt+Sjji
ZowVogGtXCyDeU9lg+G6mNFAV8tmdPOIZIabuHfFcKPSi5ZZUXzulDOV5LfU1ySNBJtl5kZs6oVy
wLTDfA48t46uFGnhchnU/wFDmYhwFTNMZUeOr0C7rEyfznSdZQX5XJD/hiGYHCw+OkBP3M7Mocn/
5McjOgur/5xXXEVr3sF09KtEFq89IohnnqCCV5O1j69cpWX7EUiFBUx1rfiyOE+M3duHhmSbb2jB
bNrE3/Qs3Npf614OEaycwFUgpvrklK1U/OKr2QBNMEii+uUiXdzmua1U8cZijzwh2x1CVsmCSLTj
jpeJMAZw9t6uttMqVIwz4+C4HqI4DnISNDFwbEo7mvnBdG+QqPqfCDUpkq1tohFI1AIQTL6La1z2
aGJicB+yN5W/FnLEpLnjMiZrACyyI60V4hfJKtLDRiFSaRjigS0vxobMJP5HMb4v/6mb6IeBtzyf
LFwzYQi5+m0UUsBs8JvSf7/XIvsG27DYz0PnOmr3jg5VS00LPdAXOPZ7rAtgoC4cXJz4ReBfFpCB
gnxMPRarm+RyeSbFm43asITP6aHNBQrLLAyIk4KHYXT4K13fwHoIwIVQyTTvfx4pu65Xu+Vagp5x
N4/wZmgG6XWm78VYytenSiyhqKGLO58iM7PeAu8gWeaDcuE4/iBV/ax2G3hJVpM3EIfuRA86Lzfp
CHKrpnVrhwy+SOXaglVmBjQp0OhL+p/x8eJCa44bHFbLYIR82BT7lHNVu+vSPYCam5Qi2sK64R96
2b9ZV80wC6wIjpnlRmBL70G/JO9rF1f3H3FbOnAaNZCwQpftZsfs6pFJfA9eHasZZOC+mpC7KE7j
CYB/Q1TtFiwsinmrppPIUUNHGb0o8/WjByjrK+8Id6ULPUPK3+42mk/yQ2Fi9AlJ8n7nt0TN7uki
j6abVfkXX4RCdJGiHChAFhm+cpAQ1Q5GjEvVL5Q+knTAtLeWXGplZKQVJf2cthmKarckcx3FQZCO
oPgfNXagxapYBpnVeBjFHgUpmh9V0JnYBUZ1XXZl66uSeGcv76hXVq1+3cypzRWqCR97SUrwswJ2
VCJa7+Yor73G1Js8Kjr97PZEZhee1oSWevkEtPyro0bKpJDJ/G0sQLIUMAFAS0bHIQN2u0tXL9BU
jNyq7TEpkQ5GsYE38NHp4AogL/r/Dieym+byif/biNEZjkA1Ux7Jh5QwipFMsTzrM0uMxYiEmdaM
0+8sHNwqDVnHn+QtwA9MHEfGPkZTy/zyvgcaJENWeOArzsiMJVkDQRn4Owo3o3AvmwIhyP3A0Mh6
hqtDYT9Nc22Df/eO4UoxcNZPicXeaC4sqdt3AX+82ElxVAXdAnk/o6ka5qWqjRlgDDpDnYj9ncxm
vleR2SsZ1n1mkn6LBm2Pr0+XVjv8YJlctn767pkVPmvZ3dKbP7RJWYqL8J5yCy82HrM1HVUomu9m
haan6VVrfpQ+9U7r0Rq/Tj+4iI/AUrRA2Xf0EbQPPX3xsxF/nVx5LzmI+i15jvOVsOYThAvYzoZ6
8wRT5CzW1zHpWFRag1MstRgDq441dRhkxS6LQIv1cW/UsymJxMiDXNTLtLsuhAwiFsabK98enYXo
I0xs1tlDl+/dgfdlRBwR8eLgm6RHC5liKhOpq8p40clfNXMB8xHGG4JreQS30RXbgeaYMzCh4HMb
omYOiPPvNaQdJ096Q5f6nqOFQyoR/zC7HzrmPAsTMknYDWoXCFwq3xJ2gjvm3Kw9eDgIfGcz+rTP
ke5ZLvJQ9L80lL2IaGWTfBNSa+WjwyA9xpRQg3cUx2CkLXOXvHX8b671M/zQhpCGF64JRy2UZ7vx
JxY4BnzAVhAwYBw90jIkRcK9sZfve2LSKNg5pzoSpKmlOT8meSSRkA3ntz0HrHY1tprNIUvypVuD
aU7kPBeNSgZLHcN4PBDilI0WcHSjTE/1adL+aB4L1IyX6Av1FTSqJZIC2h3a8nNTwvTrto1ERdZo
/c1b0tq+6QrddS0gaETHf4WZx63DuN2L+41lFqk/ZN5bmDl0ZaK756cIc5Ndg8aBFpvYna9Do/54
n84rONgAmQr7mvFFMyiwBnfgvGKoiZu7El6YVZVC/vVNyt6L/Ziyzv8Ob43s6lVTeQbZWDs70Z5S
d+8EC9wANZwoBzl6ZiY8Gc9pEkHdEieULfXprKwu6aEi9521SE59ibwX9DoR1Lv2JlISlkkr8l2a
dzGqvj3l6iNJGCdiz+SyxIV3H9TnBSgZMMUSrOo26sPmIIV6yWKiKeXt5daM2to8KMFPauQsdI3n
VctDYoB/GUK74yYbNngAEHNZhTZSv4E55bWbW2CGymSjm0p8oVe2nmSt/+nhvdMPRFuGJuopC0fd
Wgl/3grsQ+eHmrb9tSuvKzwLNAAyD0dT2pHksoaJneFqLofgkWZ6RWTQ6h+QdwKX7ymZSLRo6vPU
a4l6kRcl7Lz7s2R9+6f+OSGlxynJld48In5lqmG1SAtQtpWULQKecR3MnkaKrMEhQUif9uGS0pt1
OP4rnK6FLUptAdy8ilzH9N54N4TO+ulNAkiZuNwuSgiykKeRTjIk4+GZux4/Te1GTmOE3KOmTnPz
J7fn/ZlvtMTZIOTZ5+3ysKeD/QhNOMCzQeA49T4Ntl+4O6ZjewFr4OYx4qDIUBY5V0m9QYtIFWM2
kLRKBd+ZNtC0LVWupF7Y85nqbiUsj5T00y1/aTuIvVn695q742dWztHm8qDSQh8GiTOmPPulFKna
1Vs1oiqwbgEqLXmwNR1NnCa54gpOaAt2Gj0KZEGSUQ3kooVaVNl5+kIYfGlKyncjGDv00tixe8MO
ARGLNvFVSK4iqYhaLWkpcYMD9651xvusEHWus9vb1Axy5Syu4Z0w4k/+DlOno4Duh2pTl0iOOiFn
0+w6XNun1ps7nkH2vSydFwCm1xo4qDS1JvbcVGea6gfUp1maXaOZOQde/Ffo6AQYEJoSG2ZQCIHE
3Z6RObeJ98n0ssDJRgBdDSA9ivGeh7/m9IqKudksMjlUmRbbXyPqLb11ZVuF7m9cGjMzqo6gQIFg
7AHKNGJXXYsNIfHD1P4PzycBxJnJ2+AuKIdN6ZB+ABrzhtjYGxdBakLsTMXlOwUyC6xit8ku8X5Y
AbxA6rf9syzobTqfpzPBLzA24VaMUBiyEwtzqap9w8JBd5Is77bzpz3Uu+3S7ERC2Si91C7iL6rn
Lp994738CEzopAl5BzTioZMNC7fZMAqcpjNkGJVd8R4POZqKwFCjB7Y9LtMq75yt94MPVgAernkZ
Jf1n626Hul05de+RkrVS8WD3JQDREN6gKvh10RMmPbEOekN3GuGK8tmT+5Ry94v0dau8nPxTMr49
AkneZdYry6OWPyfUPD/zTaJJe3f2bOs2eCx4WR7WXrI3WsIicvkXlB+fMVZTiCab5Z8/ThIgG2VD
G/IKWjX6ZVzBNrUW6q6IE+ccHl9JMTLWjWQAyW1y1lbBk3AmPgt37CVA6FMdk+zdGmdg026yvkp+
k7m9iKGoIXyXrVJkGVdGwaJ/wLBSa2enAUJwr7LTRVI+SsqULpIq5kJSx2SjBk/VVfFTXzEoqFCS
U6MG3Lzu6pCzysjZM8DRINsKCqDQxp4oFPYvbCdLyqjkv76Ljmti/gbsJQeZd9ZR17wHLiMGl+0c
hdyx5saZ38zKexWm/vuH29SSqsXbFGhF2LXj8CSMNaqUEnrNOUlh6zS1Fvt7U6Wm61kX/tQWz2Xe
yP8RMig1Y2aP6AvB/lJP0pHAFQTx1fNY7sgm1YrM1wdvlcxEz2O0JS3x8GBDbBOVjrwCiykvBhA/
Q9f7KIl+Xi6j+NW149Ah0iJYRnmLB2M1ih+MIBImc6KpoMxNPVQ9SRcld4q4VE1Zl37SEXt7zSSG
O3aztoFCkptwkjIuG9C6Y1sxy6M04JMB8XKFKHxigsPJqEbjgupw0eatcT9tfRmhuQzSbqkoLLYC
BDQIqer3eqUKVdL/3/9vpWslPnJSYU8WPabZZ7WTaB6aeqN3HAFZ0iTJm8u+q6mHS2L20suWLrEc
7j833J7+mAj6Tlp2VC6Rr/v3Gj3OjVqkOA4nJEfGD6zU+oKwXPAHy4QvAw9vnWAU54BtuMlTBTxU
s5GmswWc0VJIlx77RvsXx5hVtgQI1RHwtXWjFMOomzMyNMXFd+0RrauPAb2OXer/lqP5BYWk0FYl
fO9oubTjFO6dWIlfKH11Sfs9wZwyb7SIdXPEnUy1OUKiMaaGDYApNjLTV6+huIG1FWTfoGg5Hrxt
N1CzjHAOIzCKQqyuAVLImGf8Jv17NR7GtqRFPFXTaJ8YrLXQ7jfY78xrW8xAYCZMtLAdtqt6IJeX
tRBfiyqk7ORLR3uzkB0k+g3VScNRGxoRszj04Dy/wAMwD2wIR+pMw5kKm8tOlwyro/aCbzAK00W9
o8ZH0jfsXi9NjKrcKtxMYOzlhXgm8enjctGT+Mm19c8F+W3bw4UJyYF2szXMHzAdtoDPteDE3RDy
Lmp41VGB0MkD5A3e1s+hkoPp+oOzZky5GkUcDVg4A1HwHJdXKgKytmpN97R/CK5HyeaDZ30WIAZQ
cUNNOx49YK7BDP7pEUNsExguLPJf9YbUWlRtLs1TjH5MAaOwG+Dm9ohxGM8CEMC18KoarYia1GW9
NDntRizxgVr8pPGHmCuaiwNwJFXO2jagDWQvLLwyI7cxhApyKSkwUGd9SbRKBQJspjTfgiC8ZBXE
jU2xQOVjog535YGGVDIAI97JyWgF85/p2KdUwuEeGezjW0de9NjiqMRPxCDq5Mo9rcUB2HEOz6qj
OotyblImxWE49MrH6OuaVBL+h3i16rrgsRq8W0ZCqo7kjbJi705om7bBNWmhReKgm4B61qFALF4O
PSoAarVkNpy32ZdQ7VNpNyk2gb6jiWUBe1oxjtIsW4H+OikYA4NZY+vGlEH2rGwamknajbPpQkie
kh5uOhu9RV/w/iI1A0U7u+WyTIaAgYYqesKidRmnLaQAnB1BRBizOTnO49yNJpCryChIOTxq15pv
AxKkXbFPqc9AroIY8OkBbEbJ7wQhvxx6zC7SSeKkJmnzw0uyn8IVBlRhiPKg2MNp3jBT4/kv+TiC
2P53uUy/glSEUPY0Ynhx1OmcB0cFZjf5nAKG1hmCNZk6NnOPKQDEd8z0/ad4orXIfamFsSPP8HRu
ysTvq0bhEaxKowcVlbpSiiul5b4YLrHB9pZYzXzcz7loTGR3UCiz8lSj4pnZxwVC2dDu0DoPYfhV
LaX710hQ16yk4OIkCz8qZ2QRXXInaVE7TY14As19+lBtD66XqXF3ireDUXMM/pTm9m0+dW0JLACe
4snt6onlezglL0XEGzuzi6tJQT3T6lR/H4KREKox8xABDC88mOpJ4O/SUPjPWlJhnfgz8Ux1a7jx
iCp7efszMAzia59lsKsUe+3YhMUj+TYpemesACqoXTxwIAFwBFvLA7GaU21trHaFMbS8Abas+Dyx
hyRVntM8wrZWfWw/WvhHuN2f120gkE8/h9rXMbbFRAPaDSUYlPWwMCQM7nt7N/uFrqcxPuWgyLnU
7wzDiqHsqXCIoplzgerDYSBTodw6DAbCCsGt7eT7ZWQVOfCDUfLk6K9JuyNzp/WlQFTe6LtdcM2C
AXuS+Nb59qFTUORz4uGurTMHVCMa/JcbfptxtUL56ShfEj7AF72PyVpdbIz78KYkY2JQbvxstXAd
2rxMC6qAlMmC2ByPeNCQLeomNuaRy2N8L2VBO9XGS4ijsq5rSclsn+q1tZw/CHF6+Jv10CIktakX
Vv49d+cKLMWmUaJy8p0uMNkEv/WJ8JDDQ4JgbeTT3fWqn7eiHPtrwljhrvUZlhGC+Xo07o5qdmS9
ggEFWqMGBKnY0O2CUdkdmTgpVhIQ13iMNwjwD6jY1nCv7PQTMjPcYEzL57qreTETxRJL2++MnU6L
iSUVqvuCHyflQQ5bQGinCfv56h1sCeaM/H/fPhuhas1vpyXgyJY9LnP5gnLC9RDcScBP1iccqmDz
DGV+JH/yqHfl9xatmnICgNlFMjE6exAmNwKdCR7WbewEMy7eHl3+e1R4axNL0mFK6vPmaTcZL3kF
rjDptGxo84+XAGuK+NuYEjQYVCW3yK9NCrbuRvx7l0B38X5TjYheu5Y1v++oze7wqWiVk0bwWeso
ZSuwE2ifumtPYdkl9Ke0z6QYZmh0TfzR0LlUjQio1jBjiYSepp2lesgurPsPE61x0OIUJ+m+K3L3
humZAox+jlVaDFv9SUUoX9F4WCYCzh7FkxIfY2lIWEfk4liQpsyW2rQ+qNatRhRXzM9j0dAM+//A
VtR1szIgFwfe0/nYcQ3nD8T0aN86DHDlJOPIWr8S95GG1YDNoMbO2mBQjH0ftN2WGOImopkj4cI1
E9eld+DqGgJ03LAM2EGFSKFmX6ZduF1TXbHKarVZrvuuLvgDuOW8x6B9ICPdCi6lPXcY+gr4+z3m
Mht2i1SReNy0n7VNanIEQofMWayfOhM7HxoE9LJYaOZef1EMPJ6BSWNjg7x8XiOXSGXOGi+OEjRV
AjAnkNN2HDaOIMuWvOFKjfRJyLVIA4O5jqe8sHWXMycnd3RWAEFhFdzw/hp7SjST2SreAgl3dWWw
oPVQMuqZatNyOvRpQ3gArNf4ohsxkEpGQV5tYMW5alo6+aMhtVaHTVjfCLq2HI4+Q0N/spJ5UgdT
nhy/E8InvSlIMwe3F6SGY43CqSD9vy3H02b6B7nbiXM4QCsqjBvwQHV6MpnBB/Y1srYC9kUSIu+o
cNyM8+LJQ+e48i/H3lHCaonr250kuYnwyi3YDQQz9Vt+W0OveU9fZk4R/RZZlFC3pB518j1IjCRf
0gAZnrycpwgUmi+x4cA5dJqyEdxiFWzbHt5j+R2b4K4HzUxvxITzJRFFeyPXwyIIl0+Up4xkd87C
c3x+6Iei/uPSj/nWrBEIrMQlEdRkXJHwfO43Ibf8zx/vj4Q7sbjbjniVo1OkPJhnFcW0t62l3FLi
40gaF6YBF/dfSwCxKBWsrxFleCKWMXRIJUtDEuFZI5XqctfqQN0gNIA//cYbVWCH/SKOJaNd11Ty
O8wM12Wp1pt6VtrCUPmbRYTvpbuhVBPPSyL9xyFzM/+glu5Qjxm6PGFTK+OkDDAPr5gykq/jn9W1
z7xTN4av0mGF3Fi7ycZQunXT26mSqFi320AtvHe/7/DSquxoIfjlqn3MsECvW+9MMQzIce/izYY+
YQPw+8hpIlGJZb9GmQkRqkxUQ3WQN8qHeyDdNac7lCps7fPTn+a/QRsVXgyRfpdZ9fl3dv5PJkSa
beLw+au72xC1dBjQdS3U+fJPJiRd3qpLzqDeKIQbJB99RHzRjwwgMhGIGKWKaaVbq+jr3/BOsL6g
gFa3Ecxu9Xoj8vV5+E1BGFoZMwmNCwksCxozsSxgdZJ4HogUVx8LWD95KlWlULK499I84AiT5t0b
6XZL913wOlqjeW8ytU+J4EHrYTy5fJLB3gHA+BEB/5H9SZRITkkcafuR2sHh8DBwwaaMJrwDJhmG
f/3UG+qyAQm+EvJan6wKuACPEum82RSwjWmK+/2eKS9O8meAaVUZAd/2JiFpoe37DVNm9rLDm4Pe
O0ldhwjwn9IT3a7hEJXNOYU2u450UoVZ6kF81RyFB3uBG17aO8nkgjvs+6L6gmQLByhdPKnnJhDQ
mqWYhMvcbZ656pbzTs3+YakqcpYt5b71A27P4DwkHYP+lzyZzJ/Bq1bJbC8fqXi60eXPHsNkmUzz
wQjyCbMoJ7SdALi7WF5GtBuCx4fP3X8PAET2sixEKPmeMt149q3pWrgYmFFTv4yt/qOqvbDU0PEk
/0ohfH/UNmXlcQE9c/IoBbcm8AU3uyQhwtWPO90vyGIY6+c+9qenrndfCiQoISKvwj2eX9JxSnqj
HshrBh0ItbflSzNf+N8TlZs8zhIqpbVLnAkVWMW9+eWvwBdhDRtmZhYf8zaVvHF3CiuAmBizSoex
rr0URty3kIBvb/ps9CsSIa/CHsvXFYzL+3mK2shReIxdmG0rBu3dGz5rYjyKsGheWrmdEAxq2au0
tMcHMkxG282fU960RyamxGLunGvCVzhG3TsFQP7xGxkejaTsy7ZNuB3Z1xp3aqUNfTvxFkPmEFbF
oMIFK74r6RrKfFUTbjE1gWYO9palhDufWqK9esY7788woomXd3iGMUwgVOwXbqbZOxax+HWD11x/
6v0p5NCYm1oqHxiU9PC4y4fLzFO0l1I7QNkE9tXMNU0Ln14NVMTgZ5JzdhpIMmdobgNt7AitKqnz
AKMMGg09YMIajLQzmORqmIGLD9pRTKU5n/mowqaI09yFCTny2+XYGVvgn2W8qcRHjl3iuhU/a7Mn
b2wKMP4faXF2uuQU2kzIRoO58v4mwQSfKjDU4g3QzB1K6zrQcn3AEk87LEcS4P0Bepnm1pUKmkM4
WcZihOH97LTOtZhVyUm0x6HNH34FRVq+H0Bs55/y3U6zMW7J8i9InuXy4CqUtbYTLw6HSkPiIsZc
OeVLxay906vuwlbhF4AlynVaGV/oRfhuno/xVoy2GOVmfE4pGUx3aGBlYj2qeXyqaqa7e1rCuOIZ
myuhK/Rxr65jlRrXuUyWOSnRTkgcrp8GDPuJtTsCNFK5JgkB1ZQPgYiaw5k1DoM0YuvfokAh8Yhy
XWk/46zAgaL/YR5yIuWFlwOwDy2y4OFMWBoIRvd84hvfSb1hWRAH9KmJ/a0uhTpqkhMzQAQw4+pk
zyjP4Ozu6g8zT9Cq2lCVbNS8vyIUWZ2qB3fTqFZdLNZ/RUp4pCXDyP9spm3f6dC3t5KLtOHDuxr+
gtDvy1NGegi6LuEje8PScHW6NVshBlfVNUFIiGm2hlm1p78A1RFm55qsXsGiBgEeCby6fLv6WNRM
qmDoBHLwGOZlRPRv/bpqfMEJf3ZmqPQOhc2XRZ0SrpcDdlO7d5QE+lfQoipTCda0MU8Wdg0O+9Nv
toDXg54NwwSiBiLyXMqFm86n8hC3JsikvqBmZrhXV+IVWV81JqIyWUvOLVN9arDVHkhJtZwYBCEK
ycDcuJC20degRWhZFEiwQ+D/KxcMVKVMTq2HaDm9XdLtEDoZFhm9YnjOOZ3zZwrTaM/A3IgGksYc
Sm0JbViSlOizZGOZOksf8PHtzngC+8Fr+620La3ojK1xJbra431MVIcSlvRtnLoSsJ2nPRI2/iuk
knfyYr2sRs0ZliE7AaN2EZ1h5v+2KiIt0mnfyhVUnQ5U5JffxRbHUWEOeBINyGWSBS+A5EhSP6sP
ckUoWyPfWT7LVvCmOj8CJIFDU+gjMVh0PEz6dBYc1VzOZ0JTGTgt2MBPzZawUZz+M4qX6cirLOza
socSJ+G24pcJVWNuTor30kVDMfCQOqp6MuJusfRtVt5MN9BNyfXa85kMYbWpV2Xd7eNUSGwWG0vk
B4BIc5jUvbv1HAnaxbKNrGWedUL7+jsF+OojSZIZ6miGSwtWmKEp1TqauJnAo4litizCvdKNvdca
RYwM3MOnmrYXdzE5vkq9KGPHxom8jw+15FgEcvi3Hj3kb5cbPSBU2LssAUoFcFgj9fsgxkuoxdVr
8wnvBKUZiWocZM3WquEC6dFX/LXQvi9BIYbtKTX3w/vR+pQ8ISDn++XNqsv819pWY8s4UkMBKi6s
cZbLc9eVH+Xxh7fa3VMXZoX80u9+trLrJJtOY5WGua/um1YLIlBhbz1KYazOFALhKXfetwSOwrou
ZCW2jEaIYLzufcXSefOjg9CIvH1oqlQXtz22JvQq++UKasth42BE83zUI4hseePf0fjUxYHllVUO
J9HlTvVG/kw/r87JiEoQlAE8/xPX9O6XjGxPU2WymDGl/5MaJGIIWAyx/ovH+c9dcLHUQQzrHdlX
xnK7mo4XUu2GAjXqlCnRIER5KugAwLymxN/dTwTLyEqkCf060VmSLmikRb/EDI5IWjgvARjrEzB7
4sgdYnzqkYn+CNuBAwt7dSZPDoCivZ0VBmoN44NUyswZF9T15ZrVC8Djdgq4uXGyJK6FVhyBZYnH
o/LETVaKqFJ69DXxlvbZGxkcNBkb6tDF4xg28fOLKUpHSVA4yGeaaI6RGplwizqy/MAOuyfj8IDM
XDQ5kc72bTy679xQeatnvoPlu7VhE8f56nmYc8z7Hg4QM8YSNIg1e/5x5KzQsKHwTz6fUzA6RYkh
co+cBzq77AtF8FbQJ8xVoFXBaLYah5EoOcMjvSYVj/sSDfVk16skYJLG8cA97PCCZtHZ+KaCfbO/
CGV3ZxBGqsqZe/3nLMoCmO9P49rcTEPJGqTcGjEl933WZ3BNSk1D+PdOVgw9ZXwO6nE1MuvAk606
gWSr69Z7poE3T4NRx54nocCNZSiHKzaEK52Hu9MFB/iPWgbxlRkCvfpnsRYznJCiJ1P2sk45Ei95
mXHVWpD0/yXTw053Sc15YeOFsTegvEKq0CfKi7xvKf7E3p2TnDlP1pHvh8yL9BovgGd3K7aq+3pr
Md6qUSIzUUJZyUpc1/5bY8+dph//eV7Qp1+vB6S3N4xLC/xwImP14nmmkGlFPwKto15Ys+UjO7Gl
ruqcBnE+6uh3QHDia+DTITTFytdoIQ7pg4mqPHHJiS1v5AKEtmMSSnO8CrnAvhdB10P7zYO97HId
BpZQuqn3n2J9TzNp7UEg62cehIhB+emMn1VNSYcJK2Zbn/J+spUDEubPgPB5eahkKgxjl1hGxvzb
MUU34dFuSHN/Ft+q7GG7ZGMjGWrByelwALm98n66mvgO77Ib+diyG/utfzxfmBhepNSYNLXuwulG
okWxuK43KQQp0hl9IiLECFLp/kxCAnStYDgYxicslkC8UVtwDMOKELqMUTeRpJrwbMVrvCNsnFjL
rSKjahaeH50TzVMbsm0ReTq6dgxxTNJEJugIDsAJL2hTvMDdFk8oDCfddoZYiNZ7Pcy0uMRPDzoe
Urq9V+Y/aWBHd/GQJLAdpoITIXOti5WgG98eabhUNF7BHoYm2yIkkzxBK4uY1cTNFVbmx1PRyzIX
RafSyKmYelxZ0qI/uErNhCrunp940adQ2eikGm7en8BQtn7VjUxPlooxl9usOQUWw7FHnKJ6F0BT
ocvFtERmcLwAugDZx4FYA1W2wFsaqlHY0wE+Xcf81+f4U2DKDW6iWbDEMRfJGvFmwoF5ExMmMLQr
YhkAa+1i8Z5fITJ8/owxhzjHmBpBivRmU+cxHn6oRwNRFVboJnnOzGsn3gpm3HGTTh0rZqeMzqgP
CFGPRseAt3ckkCFHpcKnNLKyFDkvaeRDllYfoipuGfGR4pH2Ssvv4wg3IdxaciWMen1NaA5PC1y+
y8E96m4KzNXi2vrp2I95FyQOJxY0f/9/STvSzmVIvWwttvf+p2tUnGPZxw3g4GnQkjTMbV+se0Ss
oME7ve+XPRdD2DxnzM7VNDH63KD3Z9Ppl9PISAydEmb42ZNgkClqWhUmPytmLqpTBZm+HKdbTw4z
B/0glrmGNiJXUje0iB4o+zgQ0AWs22R0V6NA7L5a34krVt8VLnsoVEXSQ3Jcvy2ijwRjTcDhrPqs
sHdrUob+WSllL+QBbIXXGUVZtef5c0cs0g2G5zzg41ArpEcB8oVwT6kKiAN5A4i+9e5+2X6wyWti
W+yhPPICbWbI4mdXCIOa/k4tymtYFMhlcroH76JGTKSv29mphXcsyoG9/D/Vz0F9ZcqTtmAoKVyW
mxYceJOtx3tK7ycltAexapMYOnXWWqaOcrj61KXbw/6fgLBSPaZaDWq76OC3kpQtjLLLRXYEs6D9
z5f1pvHP5rA0m5MxU0rFlyi23aOYpaHKhBrqJ0b32GEONfVM3My+cZCHRT8ZS6m88G3QKxbfWdb5
fcQCKgyOmbMw9Aq3dmYjF3Vz0eC1KJt6nlAZpsRpfY/95IEpxqlVJASx9TH3kuar/tqsA+TmQnp8
fT0/Ko8wUMvwVEYSUTBs4IbMdzAh8epHtSJ7lRNFqtTS8X4liZ57D3njzTdrQIHFbNhcq5aZdxFk
gJ6vnvO6mLVYPoQYLXaKFyQ39lMFKxgdluC5J6ZUcTIckzJlq8BeXNhBUKfTH4m9dehiY54iHBJa
xJhEVwsNnpEupPnVvfTX6kH36cNQ++namDqoduVekmLfgu8/Dy/JImdv7FE3O7GZv5ZaP0sB1UEC
c/N8xPuJqDNEpui0x8XyaKWT+ebrZ1uPepiSdLErGF61dCoZwL5EniR4rc4WP1EfGEvpiyZZF8nD
L8cOPOcR2bP8qnmKvFYg+dBRgwLaLpwL+z2eI1CjPLKdP3wvNV4sP7lp85DIYIW1uGJvnPN5Lmuc
8B1TwjeGoq53A8bPFrtKvp7JcgFn9n+LTZQvdlabLEUwoWK5sXMls33DSzWxSb6fcK3qXA4PXDKO
mOhhqTd0XL+jMKiyWQZo/JAv8Fcw7G1YPEge9KjLfYwFKppaNQ+tuB7RgkrBvirSLNM8R4ZTH9S7
giJLpC+2l6+vZLqGFf1qK5nnCDvvnoflfjcIsJ++HZLdnzH2IgB4bLw+we3d/iwtmNP8zNBcNcZt
b+Dev72i5T+209hT43Ajefqw6UiVrWbiY/gFs9v1hEeN5Y9+V9mieHO74NZbfjl3uElggrAcHOdw
dzGOhA05QUHtPRFBz5IKpnq+msX+CfAfQquP13In4Lez97w+J2ELEUYtcGoc+vr0/8UwtAQhCF5i
6Xlh04D6cHN3o0pa76GsI9W5EIyaX2ccItM6P7YYZM7w+39VU9UumU3vrPzGIl4GVg3BXCakwl/W
YPqE5adwD/enJ+Q76h4hkJza8hVn2P8rs5uoQsV8C1F2Jn8XhCgl6WI8aYP9EneDJJo9X3le0Lq6
iQFt7yzVaDuG9RSJJ7QiR6HM+EAENZT1rggTjZTbBqzbvfJaq7CWEj3L9p1jEZjmPwkl2/NZIgh1
piZnX37/RprJW0d9rf9kjWBOqjPapL/KT31wXqnzLOeNb0526D2jX9KUJMFFwNWHIU5qc7BplIfS
iXzrx9oTnNIY/GU3vr68/dPepwnDEEc5c1LDWisGuIB9hXL5PiFjHH5nPRq/nfjYB4mYlPuIw9Jp
jwxAhs5yRZwpgGbOR0H9Rek9j3QbsrhCyuo6OlsWdBJbMnPom6RoMBhK+/Q/tnhr/c5ttqC1Lc5L
FnS3jqCFXIYZB/egbe81DtcGNPPXhkI1sSoJsGWwvXgWCEPrMemHmVYi9KADUME9UznPKXoB9PQP
nYmq8uJ/sGYr7Kf7I85/rJdwuJbVYRqUsTMYIqPIgmp5eSK8ifGn2zcDlj9a/Lfal3TQenPBRoa4
jQ+WSQr/1ryB5x9VfE+j8g68ZSYID6bjbyCOZmTP2YhDnGjbv8cNnh12Lk259GXN0eLEm1zJPJkT
meIdb7QnqG3XW1NNTfZE4dMlv9z+6UkMWxDwPnyuwYwSVVWi2OgUsMqYHQ4R171sW9+X9F314uk1
HTvLyi73GIvw44cPKxUFDY+dbrxLsqVeZ4lzDT98Yxlt/i8KKqYLqyp486ApA1Jbz9KN4VUNJLhD
CIXbEbptllE/iSDpR2cFT8AZVz4Nq411iyNR30B0axmvW0hvZNaul0/sd4tCIsFHob2tKIgi7z4t
4lCvT/SyCey0iHrY4WGNgWLf+X0tOLSpR9b5tBXRCsL7bKTqVHvTa6T40wdyXBteNeXjUaRqSDbW
D15n94I9nUpFASUIIdnoJyhDp2z1RGwrHdyN7hYZcsNo1aDPkqUXyMir68tY4zGQXdG6HepSv7Q4
cVglpwy89jNn6KWQxCA5r5cUj89yQlqVo5C6n0KvX1l9viAFg6zxLiVRulUF2Y1b4jIWlJLnyDK4
5IeEnquIJY2W0GJAFjDNbMskd5pCr6Y8b5G9Nh3hvqzrjNz6Ci3GB2Oti8yF3N/6Nl2YRufTKfvD
qrTh/jSv/47lpadnhFV3Gyc2+fVUV9i2HH3KI7qAoNjaiZ6lcjfdL4nQWQY5VziGIXXiZmKWupO2
Mvs0QW6jXaC/aTEEiwQDSm6h3TbUP7/UhDfP+TPXjrMIxxJAlDDcg3SU+Pg2tM+Ro4XrZqGIk7Rx
8tmwTijsA+sQ0tco63b8l+xseh/dQ7ttCTy/C64qLKOs6tu4A0UXEw+RMi6FzEYcw8LfCY1N1knl
Zb3Ge5/bOJrJgxKB0W4IU0eBunPftX1+qW1P5foQFX1409ddlibYsDjNq4Fdy9UJ8AxOoU458EeK
EwxZVSF3UD+GLofLCTxKQO1qKIf2gkaEJcVNzWgQGXcjMLWSDL7UQSCYFfUD6VP7NlljGBVKu9YO
lVhntGSdYjanuhvYz4LwAKnB45qqtuhHEiTvcOU6kv0TlhaPzvQwdIS9cM8qrCjW8qfRsRLYup3E
cia78buR5HQBlsnjMAk3we+Wvk1kIL4YniRmWhQR+F1ADe9W7bxLlbhUG9YQrsdwbZKowoyNkm55
tghth1Bj8c/naUnr2sgzxmXN/np5qnx6FVVJfxPvwyCdHp39CU/8+Rr6XpwGNIXRR7X5IjbulKAY
k6tMYKS8XFI7gM2f8HQr770XpCmTHSBVlj5mVcXDM+VXvEpIc/xGq/m9NDTKL5lZo4roWclArrLY
1M03GRwg8897t6Tz4yF4BZr3Vvk3TfsPhUTb3xvhE7/mfrjMsGI9o667CyuRvOR6SWQkXkF1OaEz
cKq4gThv6ATnxk0xCQ23Mdky6X8a+YjBddpLb0izB9wLWfZRuHA+5430wt43RHkhF6SZe7Ddmcir
nayHEhJKEGkWQJIhu4MvVXqDXdNDp+pL2TiPDSrj1DPgo6DFcYGPTHae6xNZk7zyRCe0CWOWdaLx
X4PfS+2yWA/y3UiP7hsQgLezUFdf4jdcgtlMpsQLnGVLDA/AgeF44XyJWvqDoBVnF2D544dLNwoD
OUNih5+4yGImQ5BWQgjIQ3yD/aP7/soDE63B4fOFsJogLmk7Q0uxBXCrz+E8YQlzv3Gbiad+817c
LPhaFq/acuDZv1GezJrHspYuOv8Kc1QgaIdXFizPfIEh2Ws4x2sruPKYks/8honNzdmtCcyztlBa
oE1MzYKufxKvAf/54oaV5kZRd/ZzvPF0CAh61v/PHF1pno2WnPvSaTvvtAeeC6Kl26CqeTTqr2Fc
Tx0I15DVJbTDXw/OyP2E5v+9SLx4TXAkWlP3+6kwQHoTV6bVArGIzKFAA+9gn9Ft71O2ad+ePV+N
mPA5n2ykrT1d91g15ThDyAw15yX8Ke1gSw4O/bzJ/WG71sZV16OgU9em2b1sZXLgNXZMnbHW06Iz
rqNxCIf1OdUkKwxiazk/et7n65qy0Ktn4PSHFUrtLncoM9d9qcxsIzbpvTU8aLQ0Q9/PrDmcJA2F
TcNFzumd7+gBLlBqo3z7JFVA61+gfJmqv7jgAOPJLPbwaK3rO94HB5IYvENJSGvWlIUkJyBcvFra
1f03SpY3QL5f+m5dDM8eHhqRlCmz4y7h7B01hnHvH+ogqQEbcU6R0/p31PHZjUjw4/6sD/6/88Cr
5/+LFob+Mc68RBHWdlXLh3wJobynEfH3373zKHWZTE83Zik8Cont1L4IXsFKxZUvWeY7Io7hbVOF
jFLge0xVuI8imMUKGZCgDCsNylz1L1i8wyuNCZ2JxRoGrlmW1wiko4ty7f8IPfgHSjchRV2CD1gH
wqByhcZ0B4NV1dzy985+ephOymz0HA+y3ML69sHdsajGSGzFtpq+Q0mY+aUoR6xsqXh1pcIpQjH9
0Ajga1SyYUcRPLtIrTt5jKr1eP+9S3KK3BBvTXIXHswiRy2gZICRa36Hr6B/uO5fHcW67V8GHWgE
A90ODjcJUiE45HnvnbNpMM69Yb+3j+1E+bkQQNLyK1Z02T4HbRcvZeIpyGD7DnaR10aTbTnKmFDo
SXdvxfPA5bkbMtiDxWgupQP0OnrHStzFFdsxnRxeFz+dSJWnDLZgr7yPoGI34n5oBxxst10LZrC1
RZhtnZIcUW0ufDUuWcMLSkxhp7o86sI8ia9JdxJVxCbKRVa6nDJNrXJWeg9AdAYyTKlXDxpTFqWL
l6MhUTjjACXouVB9np+aXxUHBTTUhzvOqK+3cZmy8bgF4TK86/k8KfKL1kOCE1BlYcw1gFBAhiKk
2xDtYRJ9YTWJCZO84log9+WoRVVakOsKT0YbwIkQzJ7K5HXL3c4RLxGoQoEQHExmiuI945yT8snu
1Pxh1SzY5xtxFkbut/oJCTrd0Gubj4d0rax28ljc9UKeBwsFLxXBYcLye0EAwq3jh60x5dazQ0p+
5q5nU+sXrOqSdaAWxH5/9vGa1rOs7yLnDnm+aD1/Dy148wrCPiPM6I9iSUD1NtE+3QEfxbMHgKuE
6w/ElQBSjoMPegnsM02bBRpPBfMljQlebmBDaApsbL5KxUupS9VZaRErNtPpZXjHoo5DGwxtuNP0
lhULodg5hWs8dR0T5Sf6GKIgXaqDpcYhrxoIEi2XjoNxnKo24XCkfWN4PLQ/xeutJaMxbsMMaCwZ
yKXyTzh/YmyY/DnX6auwnrjqDJMNF+X/ovt5sUjAwB9XjsMEUt3ej/2wD/Y9hFtx3ObKaDmfQS+E
q+k8AAkHKeSaTT1Ae8qxYWMm2ATkVrPO6yugFbeG/fJqsPUjq8VH1x8FLYHtn5/p8mRfw8Nx+zb8
AxTiEzLJSAY1r1yW57szu/O35oFWMgj3KbYXfoF0OiY8jF2StrjXyk8mpCbRNw+YDRLHpxMgJ3sq
tYPTZleuTT5uMrUEDmmHqRMGO0rXhZOwCpdfSjOSjVb1YEj1RS9fhaaPGnEqHoP/1S8sku6kwV4c
bnjA9kGuyKXmK/5g3IUQYtqf237bUDAlWXygJztXNdmmgWLXwVbkI1ukBspgzp9NgJZKNdPgvo0R
+zyxv4AEMZpMDnDacwgzPsAhm36Qx80R1zI1YXh7vVsum3RxMQvIezyhhaSHhK+UlZu/QIF45V0o
fg1TfAj2C9fcKXrBKRqbi5EHiR/JVolpErtsejRBLYVtdW6RquZYd+vO9qhPkAvFwg1WvGCsbStu
YumnmPyXYVgcLpbmmMIJWygWyNxeexG2R6DnN+hPl2CKRCms0cmGjAe6haxedm1PP/bDHMaUdqZC
hmP0NN6zCaXgB971Sz47X8H3PQMhWuS3NMYS0zkuYNZqLCzJe5r2PxD0kFThMPjHJoV84h8YHZSH
tSYHkMJnBGzH0yLluFwwkhI+lyFI5OvTFTwTHlBvj+9F6yL6oBaPClXEpy2pdUB6YBNi/yNB4Fpt
IB4Et5v7mke4CWxkLZw4Hvzx46K7eYMueg5LdRzniL6aj5JiovuTUvdiZcfXB+U5uKQxQ8eAk349
BCROZDhDOuTi8fNciOmd6uVCGFTeZAFdaxpVVdyKDYfgYp9tP4rlBW7iMRQA2ijckQcVEUCU/U2y
ZlQvlk4lGjOgMH2uZBZ9uEsvaV/7GdGICoJynrn80LOj8P7zjL4npynSfiKaIx3gtk24oGUHRPDs
gm0Pw/bZJc67N5VgfSkDsNTDrG9ou2EbOKY7G0PGM5IChZHMYPOXw6o8wfGSs46PDCdRzcJjIcdf
cBg0IQoiiWyk57jNHeYrshOq2VWBa4D3F+ytncVZxhioe4CJKFW6fzTYC54bZZXk/3R/o26MZyXU
4VItJMVNZ5XciSlS7zIdrIu2htzftuwfCGi3xZMUGjq89PcrGRK7Isb06gxxDA+Sf2JoJxpGbwvq
U8mJZ7jti5JkeO1YM/xM5m64vQ3uyQNyXHa/uSKUXxNcsxmj/Xn1uFLH2qxuU2uU7dmjKozsulmI
FtmlUsn5I5jLTPiR4KcaeEq/IvzmmajbS52tTzGEwA85UXMAu92eI82k6/Lbcp/DcfgGnoLAcdNf
xva0UOmOrCzXGl1xBzgBlLjNzAuT9g55XpHKckB0j8KWRgTDLxoNlB0OwjmSl+8erK0H+A3tci6a
sp/M7dYMtXe5qjl1Bic3t25TtlUpVtNMjENgOPPcb69/cld0RCFkBBmvZeQsdJPwp2Yph9OGvGZt
C3fHFpfTJGYMzfT2FvHut+MYFRE+zkEog1xHjRixlSf52ptAmd65XP1QBF2SNbceyFvZDLcw9Ld+
am442MRMqy7YJsWmPFPyddUz2DKWypM2rFjJ5PwoEh7OLh4giHuTQm1Cph++nVR+/OUa1gU3rX4d
XulMWeu0/LuGQs6u7h49zVvCvbDvulsh2Qj+gF6y4hBBRJn5ZAd5ZkynXx4uKlU9gByw4tsUjMeq
j1OXuSplwu0rrTV/p8hOEtrmsB9WkCYPXm28Qq4s+8YYg1dRReFrSphEem/nHefjAe3hi7EkvvKC
OYnhiweXrJ/FAYCRiSIf1HT/OCdci3dBfrlSgGJb/W8POv/duUU9tOMO+pigtHyNvqLn7PKp5Pry
3D0FGtSb5lCQ3RrfwmO5yQi6g3JjcxbP7++kKvuLxlf24DpcL9/p9OiArHUYrnY0l5zEXsjzFTnC
aT9e5SNj6WxkX9MA7sJ5vaXrXrJIwznAEyiTOT0zMr6/Iyqav1a/qd1fMmh8Ber7iddgGpoIjiVc
YbQSaQ5JSBrnP8scQF3/VmW+4aGv98yiFq5oPueXLP6LDhlODAYMeR78rfLNlfRqB0V+vDEfVRYs
QA1h7yW97+mDuaOxTE6DNDj0Yt3tUKmNMUMVAK1X2b87WRKhzzHTUUllFFt/6jyAphdzynrHEccL
MUxM0YU057QQNSLEUmSgXvdxMAFvGuU1Yi7KplfNQH8+GWEOzNvR0vuDecWB5YDBtW3nCFNFSqci
ZCE20yTWOgWjFg+0wIMChH/+oEi1LL0g+jDOa6zBhgFMlLvNu++Eo3iFfHDczLSD5YuGbdeTLH/P
GGi7cfmUm/jx0t6hO22mLsELsAlBizhELD039rO3XEl2IPL7obFIHXGg3BuQW/iNfgaK8xqb8sYd
88faYe4Sqy+G+kOj1IAqr4jtnqlm0naHt8KArUB0cSm0/g8ZlaNS18sbimA2Xe4bZgO2nPYG/lqF
do+3IW1p0M/jhPlMXDE2U77UTEnqZFGVpagdBqZGsF2joNOUZ1ZwrQMu1IeJUI+9/saxaClVSscA
fhNMEvjBuMFekjRiEkgvkRGSFveLbe8ByBvELq5MM0i2/ihnV8RkJl/TM7BXBDLZA/xWBuhx3Jt+
LG+R12asZGn7rpWwigmcVvl/aTqw0k1/XBaYdZ77Dmgjms6mUo/LxVKpOhAPLet4aEY8EQpfO8c1
9KsOafmFUD89xNahPloRt+B5u4+WQIR+8LR/cseRNqxyyHQMXZ0YDO/AuZ2RWfmktORAgyeU9BQp
/C1oIb3ZR0UVTtiur78b/mlmoJPnno6YlEdTPU7cuj0HG48ozJtjhfNZMWzxQGFnvr4Py97jL+7s
tXAbGJEmd3YdS9UZEstEaKNkkSOsg1FV3rb3pFv0MPob0TzzZSs97Tq+A/xCauBjwGAVYwed8nt+
W3if2hobzViJcQulk8yGBLzQvJX6bJBiHbbvXU4m8E9FcxO1uKoatBfr+TynLfn9W+I753hh78F3
CUzTgWoXsh9B38EZ4i5byyXRMckpAAjc2LJxbIAdNVJ7fwYHDNcFSl/tBn1SLQp1Tp8F4vibQfBr
3CpJ+DNbjAE1ANprVsRNzF08t4QSX4iLVdrF6daAtU/WqO95XIKQsLZknjltIPRv5GCB0Q2FIYsP
o2iQKxiaVY3TfeoxR39a2pLEXd9S3HSgIzjhsZlSQGvi4kGLPmUeEeZNnqo3UNe+HOdxoxoqPVwy
LQnEHi/4oONZVVJQrbSxBsKP70/lZWIEFa0sA+HLCBl5nCGtTn3UIN7t2AzUofA3IuqZgeN5yy4p
zMhT6Od2jP15RpTF/kvDfiVWuKqffYzZFu9ij0Me6bqBW/oC1X0KUTSgmtXcSYe8tLcLiTCZyHsG
QnpfWQIkaYuCYQRSpLfpcIA2u5SV5MkrA/HWvt5vuocfzHhcrHsmErd5a0T28T4wwrKwqT6AcKZR
pDP7WJEu5/yH12KnzJG1un37vFbZPfwDEhIbGrdd0Wpf8bAAX0+BR7kVGtrO/WROqMRKIAcQsPIr
eh2QQxcb9NC5uAU82bvmfzp1CKfznItahlo4cwzXB/2aYZM5Lq6wblDSupWmkeo1RWc3bZI6UJaV
tFdUyxGE27kPk9ZlvizOEbX01lJy0461DmB23eE7HNi9LaiMrlRcNXxPSgeaPXYVKWEOTicAAKBG
amUS6ouoOHgEoPs/EqkK1jfMFWZ6Jk7iJ/2hrGveN5hAdYKiGvSOSY028T5qk+I7PviOdN40dXuf
8ECP+hJYNGs9EmW0FX52/+OLgP/Ao0G0o+n7T/8X9reurlitGRWJppzISTkonhvpXTWGmXh63ptQ
h1k0fM8M4UIR/UHSdkRGxRBiuoMgVsBzVwzxyPngOPxaXKQERj+8AofKF96xWcKD9WMGmogTA7iB
l37HKA6cfmNnZK/JpIFhcp9VWSf8SF0y8uHJz/DHMzwpa6v+dBiSJxGefeiizq5N/gv7AbJTR+/2
UPsPjzuiqd31Hc9Ff3LiXO02wwvaKrkmzBant8b0sKORcIHeftiD3Fr9gbFmtpfrvHSYUOYq9kEj
jwiyXKb7+0bs/ucefIVWicK/wbUWZkK9pMcqMfM/UyXOHu1JPLkCbhC08iTLo93ZF/95eGJJ+S+P
WmOMvpDveSEhqgkF7QSZCH3MOGG39mKa8YL3aATeFHktBhn1Oi3DTJAIf5P/uCgVpXLKING30zdf
fJSfnlgrVQAgzMhA7UeMkyEBOdSSWcgGBSvvpoQy+Gr/sOqswYlh8ol43656IHd3WHAEpr1bw23Q
GxumGCzyaitgH9rf5qn+vExu4l4OA9/7by8Xa3uCXo5oQHkzceI//ugrqibSnifo3dVyKxc8nvmn
eUjmrDrRz3zLf6S1CT7AM50bgxL9uf9Ddy9kKDKlePocWHoYZ7kvwKTh11+aV+kVlrBMC9izuPj6
neSNJjkRulOanhkDbLxc3d34Tb8h6NLMDwOEAxCU/94xK7AjvtmEgv1qjV0mWYt/W8gkBaF/GGWU
YMSOcMXAvl1LqPy0+uxhZ8YuRt7cXV4K1cXQLumf7qsTpM1gjM433mIgqeQ+w3KjuDWfGZdkHKkA
AnVs8NmnkXXK5LZpMKPDN51gT+769ae0MHcvTpb0XoDKZQFYQVek/JJ8/BNsXvcAqFc0FrAJmc57
88C18f/8QwLRKTw21HuIHZw3RUm7vJjrd3S3nF/QJBFr1Nz6lT2PuxSKhywsxyATXUt8c+UKDIWf
wE1nxyV5i9mrd5mll8azCskZ5zs6O4gIb6EqWPwtX/2howUtuB1JkcZ6N1Pgd6TTTu6ViuZLF1n2
dSwqF+Sec5WFtcIRgR8L1exh2QPRDLYnX9NXR9b7q+RO9a7dNmu0VPjbJdSiCEqUJe8WnUqZjRgn
5z4WG4Z3n9x7Xjd4lWzyEvfWVudtTJAYPCc6XAwlfDj+AssdWStYpuEeXwmL0By8bYqOxuuQcidb
ST1Y4ck+NZjLL7yznpe1jGJ8h+LR5vUjJqToLH6ihCnSr8EV0+MyMtWdnWHARWZpAbudoFBPttc/
vaG6Kwr/qW+SW8ytgZHp+jkFPRSxNO0bPyzw8ePwVks1GTBnFTExtp5YaVBv7Kpg1vCqPUv7JgI/
GtCbpCqo22hsa4NlhtpxfOAt4Z9RUmvfOUcoaOvMioDwxOQAo80hNL50+vLTbeE8GOiuY6v7G4FD
bSwZoiwbyzBaNdIla5XRpqJHV5fTEGqYF7+kPKaXnnlABxSWelqhdWDUsPHFOLyihABipE7gXjCb
SpjZnPHzW/JhZ40ojoWxdUg+VinfQuy5aAaV9ZoFLKmv4AGBOJdu9HqKXyBA/TdJkm5vZMrwOldl
3P4tRmo00goZDpYB4uJXor4a5F3Xfz6jemoUsCLAQtISSNfFImMF2tm/iRdMRglwDVwnmbqmrfxN
9+USTQuuwQiEO6WV+x3H8t6946PFdeaPUfMAs+qFJEBoDXR4W0gruNBzgNUXAQ05I5bjb9blOxrD
BpiHz4/OMJnb3MNI//tF8zWUZlaSRKuNTtWXOURJqriTJ9ii+4jWbpuJlrooM5zPsO0o/dG/q349
qZlxvhanOWBqFn6DzYFHjPqgbAYGSsLNYXARk1f5kOhzZLrUBTB4QdvNWS891jmsVJslNlHeiaBA
ChHr3nN3Z9XmpGMf11qKgrqjblnz5WblQO+QE5GgRkqRJqKZCJTMMnBCPD6FOIX3+5ktPYquyPLe
/oQ8yrV3GKMQXF+6uY7MGWlSvxOaHMsWGMLnwZz16xDfoT14owyUGLHCRpObkBk1gjmcrmZ26yKR
jwbMI6Ip4TAPTpkj145E8lAXCxBFDHj7I4d5Rc8GPEWZY8VVWNocruFXHBoSKQjaTV6db6dgKLmt
JxLcN+dlq6nE9Jl5qw9EnMLUt5a/+gKUvV29qtCZJ1USOVFmxG0FBrJSEHPMfemmg+S06XAGWobL
v/CErf1Qnvhu/DO8NCvgF0w1fUv9PhQcMnqGHgFgjN6gnu739U1tOdK6/1LbOc48ONU6Vm6RmxHe
vrKXN5Yhj0dDO7gqzjKD4eZtsqPCLQjqABcV3cro/WkScdvisHM8qA2rLkRpQRAY0n4n27kw41Ls
NJuTIz0kPZ5TolYio4jIT4vvSR1dP/1IABreQnvNgXp16D0QuJ/CkTYsSkQM4e9hQat6LJStFbb1
rMYAUe5TCe0P6J9WD2xi/RlW6uvLS9lph02MoOC3A+7XfwFM4QiitnWGElV+abcMq9fQUvsrzOnr
9e+tR6XEflTO8ISlI0aIV5o4G6fjAP3+bZ20ro1MvRpV0GNl8GUv+Kr79w1JuYOo2ZcUQRmGReW0
0UnvmjrZ5YdTD0FeRwKWydIKcAKrrFtFUrVcHQ0eqPrM7bzv8UspUduMx284jSqRU152Cw4+w92c
LO2B6Uups+j7wbFIUujF/6ZNNgW/4VPPxMb7EfcrFwIvRLVb8v/Qaq38mMhERFAj9yffWcbt++kT
s0gXUXAFRbGZ4BA/qpXxCMQ/37XPseigz/s+XL0R1ipuqNTDBowA4mwdibo0bwRc90nzKscEETOX
TOwFbiN6hby6yMgzpz7WQB8A3J17Y8XBNDgEBYXipVk9WbE9sqlXMKOCK8gFjEMZP7LtBkVNcUj4
QLFFXRTmkJlrNai8an89G/VfRyXJJ3T2/BfFGh6uX+FKLSYzCrwwsbPWnsp27rVJZi0j8FfmnHZB
ini5hLo+XfssTf6oHQIin/3ujwrDx2Ayz4565cRiULJoZcHqRvcayvkcVOoWGLLWRde8pi9GKWRt
fMJiaFp4dLpEEzhg4dUqaAeew5F6jbMnuQn2PlAtSm2g3/S4zpBObRW8DbMcvvLRA2uwmV6rr3Bf
ILjox1AruZKv425TIjUlfyUzO7DzYPFvHvhe+rxk4fCY+9UKbRzsXJ0iNAe1yKg+D3qkLQQ0/gKW
DavJk81bmqZSmaALH4t62OTvrnRnrDanq3zYUnUW0s3UDtneCDn9iAwZimiWGuZ7RSVK59NPMTFV
fscJ7ReibEQG5eoxQZQEYSTh70/MGjNIgrsHqhGxqsrAdkai69yPc/XxgCfbTqoadRTz/zOiiY9s
0Y4SvI9IgRz4sNXJsux7K1C/phtQwdsTlQyyW4lmmnsoDbfu5AtHfLSVI3yMKyk2UXnLlilLGboz
Jbj7vGm/HmoXrLCvjAqNvrVzBWesFcuE2NV0DBT6rQTFplG607fPR3GYpoMnt8xQ/LJLj/BHVxFA
XFX9QRYgvzaNoJ5ZHzA0cPe8ZDZbjBoBbDyRhYWJQLi3yLnl62sw4J9uw0TPWqZmdN/ENeRW46PZ
xFoekhmw3dHLKLJKNCAfposjYFwzRskxX/ByKYUg1/PKCdl+1z0dsuOilbdba5VDkrfuvvduclve
UR/CmvdysX8Ig92wn80EH206I9MdRoz8fc478mnTC92NtgWYODQHcS4TFkoA80IKCvb7CD0hGQ+6
1yVj/6aAgislKZckFwMNUdtxshiqyHzvoJOUKrJ5bSwxVXNZKegiognjdeKmvq1AdwY8E/6yrrzQ
U8iDW7BdDQdHeCYQapCIU+FM5GRDRlvO/xjLQlJecA60/FK2Y0WJNzfm01JzxEgZpMeOCUZ+JKC4
edg7RsFeZQv+BnyvAKNsW2ZmhZ3bT515sPutNraFfxPOSXR4589j1DUhHV5XS2efTYRbVOW/yIUT
PYePZuZRmhpii+onrF9fYzB5lVtTOcj6WHZjQzsI6M3kgPvx+KSxRixf8yvadxUax+vC3wYTbhlR
pfjnHA60XKomqSX9EfPgsyLZFkhXlruNRAK9AeBBhLDEtHdmw2zhCKKdxnEITw4Uw8pYfMpKiAR3
7nzJNHX7ZQubBHdHkeJ6GyIsDkxSTRk8pVKPZR6/PenagNAoiFsqWNcKpZRNEgJa6qMUE+GByVS7
YDWd5Cn21aOJksPYO7ddVz/6tiZgrYWufhPLAe4fkdoHAt7NjBTAHj+Zm6IisC6N7zNYSzL+5iq6
4p/fu5K02q0wNzor+vACLIkuqpXgt58Ml6iI1HHDvNU7SE3481RLVoV4u+OeYE6oWwRGPcQlzTgm
49Or1+FOCnTHh3sOxxhL2scOm4l/J7tX2qlJKeDxiQ+zo2nCcpHwBVrWgK5DNry+wJPLF9JIAQMy
erZ7vE2yx5tXEL/qutf6yWZwXgHnbX1+OqW7t9pGFcPcUj6OhPrAJFoIschMx7eyWpEB8JBeztou
jkxzwyB10OY8xgdQXIXyFlZT88QypgdEVh4jewrsOpXdPWHi4ooGcGQSnyk9lvWq8Yd5Y4CJiRHC
ge+xrFekfQXZaIyhQTneuzyOgfCRkE5pPZFxBzYI4cg1JWxiTIxi+xSkGORE+wptu5iUJzkprj9v
N1g4iML2CXMgK3htZnvMyTMnl2JJfhYsf8u3+rvRC7v/ld8fZ7TOymDOIK6QGLNXXPwt0ViD0mD4
Xv/Y1WXcoyKdu/JJglsYwvtdtVYqig1veh9Y/W/qq/RA+1Sh54POAzjtn17fpKnnXWh0adCEELVu
IgJul6PKx6qOxPESCaQfGTNypL25Q35jwTAH3XYTxNXbum1V2MT28MfZSj74QMWzNNI3dvno/RBq
KbB8qidUmX7tlsVyfg3K+rabfIUQpVHFmzXu0COhDKxQlDTp+xTwqKGuHiqUnH+q6EuzfLIKqsgc
8Cb8KVI4yL6TR9xWO5dKYNmWdPOKRS9z7hMsBSAh0wBHL0NQxpFZj4ArYRUxXZGY+HZd0ApGX8z4
nEL69xR8OisBWmrbu4vcW5oYHyGsPot+YjkUOqRCVclWCnJnkBgSG8piAb3zC57cjKPwAdm1EIr0
Z7zv5uZ1UX7hMuhYGpcdyQIR5juj5oLXO48Md1rYIgW1cTZxtM1kHJFek0yNXyjo2huKqB85kPft
226gVwttaAw6kHLt2qgwI8m3hshGUssUt5yqwJCKG3yueEDl+rkZbfYAl0lM7goR1LrYnh2LXE+Q
B16APqB4dEAO1ja857JKhdFMOMnJROZWriRB2XTiC9Ltt0VBK/Ad3aSf6sK/otyQFskmFgq7t5V/
w3FjNuLihywRMk5ymQ35wJ96hpZIW7OWmdL8rc+/ltIsAAwm+V1pZPrY1N5STdhNXyK7cyEQ6Q95
NldxziR/3xldDgxwzlTh1SYQNBiQFxn7m3R6FjS3Ivwxa+ygu3y67f/S0KUxj2wOWCUIUbjJLGyt
j4dep11ezyqXoW3Ifio6RnH/GFD9EU8SXvC+LV99Ix3YVVq+UGahrSvfqrcAZpW0X10FzJE/8yiy
D/9VTaqVOldAxqWMjZgRmF0TgmfNkML+VdSPZjGQieLqjNeV1FQXC0s7Z68p95Y+QW3NPIZ+719w
ljV5ys0+uA703kGNnb277V+HPqbY8LqqFBki5bmQc9JgrbB7aoNyfBLsPXHX7jCOqFdqMuWHaXBh
cr/cB+oRvMrdCx7O3wV0FjUUf2EvgQD8kAlTbiBjej6N689MiNQ2lNK7qT3z1Y2EzWWRtaf1uDQ9
XhCgj3DIrSsSy5/qWJJaY43eJre87Raixzw0CGIVMIGupUjX2MWMhwOD8s7KH3QebsH063jZe7Jw
wnpCnNRRh0Ic0m2XI6EBygWDLY1IPskHV8yJgQW3rPZmUQuZTQ4l6vEHwmnHxpqYu/f0Mw7kf3Wy
sDc6NfM6VzOWAPat0WjJVSMdtGRimJOZkjxSw6sixSlH9EYXrkVZ8w+RvjT9mfOsDXObLYPUXD0b
kIv458ulS4AiKJ1iEbtJGXbNNgsghXAPFWKaeCj4y08ztTI22ZzmhLfvo4pEE56Fm62MymaEuDau
HSjkiSoT1escvo6JzmGh2ufH4/InveeH6Qx4gyqok6r0Q7vIPYeUwmZYXn6ZMGJ/L2zAfI/zMx6Q
7M0fDmh82Dxm9SrEHCtUu13g0+Oms+IVJheNIJJHIj0B2Fpu5zdSYcsKEF3VPgJhZ9ki2xatFnLF
c2hiOxfvLvqWOtGzcFEypgnWmSeJ4nZXkNjEV6Ed4IKe6123fUGImy6ql4l7RSA2MqCIYCBlDuv9
ucuTk2RQ0hoWysts8RIR19aVAjdJd1yqTgPa2mEYxJgUIRsGtOKQi8icVv/A1EWh/StYt7TOoyKK
yrIRRfN8lnt4kBgcAsjArhsxPW++tKVoKBeDDZgYjsx6+quAayCRYkIvByB9KCgpEvqOVxHDKXHU
xvs88/QISWyXCRpO9F5Ot692ADl5FfabAEMTPVNwZ+SkUnEl0p6U7xYgTU4B0HZrBjW26VdJXzrr
ZigVU3o15dsNi9dTGWAMMwSk440HQd56OVIGsAPqwHo0Ac4b1KK6Hvr8KO1rwoRoTlz+uWSTMFAw
zw1enIwb4LipjtWSNoxJ66ekbCRKgo4a+YQQZbAKqBWf/PlILs0biC58wmTCE0SmnOwHH6ntTCcY
u6VdInqkclr8iOY0p+tWcpw0SepHdtQ0Fu2x9FvTIT5yP+ssBlZXUWNL+hBNsOEIdhYL6gqgRhg/
gK0JbZFDvrZ0FoIhvhn6XfvxTg2YO4evujjSStsN8x25EFHqenEqS879mabGMdPWFSAim0QCkwAp
Dq+hwcMbBPwy9bQnEjK+UX4gKX4KaOdGgA0z6MhPmP1m0ibB2v85ZoZMuy61CsD0Jtg7Q+ROJHzt
Oa7TnKs8jkn9IhJQm8t+GvZOJ67rF5K1VqMxUA3My3P+nVfO2H/C4DaF+9KOazVKcUR7T3Zj6UTX
InwH5aSKCing3ELcp/SZdaSj+rpZGrDiKEd55ksOQtUM61mSZ9caOXJYHcakimoXdVEe0EHduj4T
w8ZNsNhKJgqfbpIHQxSdkzNLUNtfyvP/ukG9RDEtwKzHoDbjphZSczQ/FE3A5Ctf/N5b8zBCp+n3
80mWEcPMQZSVSZGmrY1Leju12pD21KkdiVuotPFmCl6+AnoX73RctHOWitH8Tc8ijBky4X5IsbEq
jMdpDvYjzxxsWjRw2qt7oavNk9Qf/lr34SwJZEFRTQtCBYQLmyOXWLpzxuBnhkiuqMkGnbT/oV28
1noHHviQMyydW9qyINXpISN1AlhQreq6teW9DhXvzJBS31YSg99HXdu/hoxJXtrzhighjAZKHpiR
zbYy9CeGHp4PqzDOWqtMLCYVgTNO83EiZOHj5i97qOGU+b2KOc2kO4v1M7Omjv9Q5Y7Lq6GVo+RG
s20fzcvWLNdQ5lRVPzQC1z/3nKMX5wV5G2qbZK7dPNWom+T2fT2c/CqQkh8QbvCUWrE9jf2j2qcc
h3bHk2t+Ms4cZxoIn4YcMLz/KAi5BplrTDXExs3zEEFe3iIY492QtMdL0vHLWMkeN3IQfweHpcH1
l1Gl0G8LYoPtwB08GjBcb22RL1V1kK+3I+kQOP9fPJ0IMm7tMEQX2eJlUupMwyCqaMca3FSmETs4
Yr4zNmi5CfrsYkR6s6LtwIC7E8TwomqJ0i8qbSnhL3vuSae/63zmHC5YjFvhlKlHBkAFOvJPx+4e
w146/BAAIOuVn5w5ZC/lsBv4cwSEQyFXc/hXSkohNTyxVAWGe0puLt3Zw2LK/n2eeGDeTFDvx4KI
NJUGPGJj2XoNMEiOdxiSFq5J/wFW0PFXyQyBBp6HXPkRarXwqKUCM3sdYdOsL5Tbb3sQZ/u7T3QU
RHSCbUen3wTObWPZ7nIcDD8B1028FJ+PAw6FGUPyQzi8lDVmsnYqFYTi6jKdhs8qWhcTadVdXKJW
iyPxkYiO1fg0WAnASQFB2nNA5FtB9a1ql3vKuA5AwevMQhgKMVDdyru2+dtofwZWy0HxhXpReJdr
9usgU+9MVYECyb1GhERGTYto58NKa0gDdNxV/Jqs8mC6tpBODSh1Du/Ig8EZS6QWnH8c/2uSyXnU
M4aSRkGsPtFigKyDmzSrPUymMwvL/t9aM/VIRgJD1o7ESGs4aO5IWIyeDSVSfQA/wm5MBugEsUUt
WbD7I8WOgfo/WCppjIu/CYs/Z5N769B0SBKKn1KFY3Zdp/yNIYmq8bWnsBXgWVcFMGqOXV8yzdIc
/zjbESz8Un2JYj5ETRkCVGXmanLZvi1rLyBwnXnHjtt8FjhlUz4GvNqkmJEUbt9UOjDhGO4uFRTJ
NxDIA+81LM6Suj4POGNfo/YB0TPJ+E6T3LdNcqdbp7acNm+z7rkjhWUxhP9j3z/FQgP3MnV+Pwpe
hFeiTIfMEX+UznHsl3mUQecToEXq0hMyi8J9aEul3Gf3Ru6pN+6vb6M9XfEKnos3m4NmgWEaB+bB
i/3E7fb7XIbkPASchzCu6kbgyEuzWu9/q7g6C3FaOVLNOhZ7uRvu2TgPhE0ja74qJMr+dtirmEDU
90PVyAYskt00Kp7o7/gfQkqFdYocl1eJixI7znrySrv98M/91x+vn169oyMo6A9Qq00HoBUo2RHI
e6Ae+eqkg2E+GTsW8+9QwGmYe42TfgLudfYrB9XduJS7xNglEXqUcu1U2AO8cXwbnItwUsZX28BW
FkEGf/V7clHg8GQsbuBv/iJ8UabXWxeNvwfsO3/Uu6xeymoa5SBvgjwy0zd84ocw37JEX5ZHCGCG
BAP953RZl3CIgkgRE/77UgWpjEIDpzt8/hsJmAhQlNZh/m61QjzeW97OQgAT8djvK6TAw0sr90R+
qOEBFLFn3ztArGz0ojOIMW5Oa/9mmz0bcvLlVatSzCvHKw2JjabLAE+u33HWNX19nVmQFFaSYAPj
tP3EsCuUO59Xvq2tAKZ4Zgjl5RpR6UsT6FL2CbXnKso1mHoIkspbYuzN2IoCZ3U1SRg95nxthw0U
CRj4H/MjEaXHpCkmPDWvq93zAEaq+IeTlRfgliGq7JAis35453ZwEf3rRU1/OeQo9vLLKv0MkY9E
HPbXkNq2ypCGKWnNpOEMmY+z4yIsoirrUEIPVeKcnd/EbrHMR8fZx8j51HvchZc56JeLoAtRioGu
LDXeKw/9Y1P3+3JvAiyEUGF8uwPEir8PYImq0aZfhRQ6RMR7ZHLEsXdBhjqANk8mTlfk0WFhSNm6
MVJ6tGzM1W2GJhfPt6HhCa9t8qmIQbZ1UOBYRP3+kyVM4iWK+gxVAs3uOn20CTFuLAFinaTQsyA+
UQhYKsetmb/IoB1KqHWZndV9d6vBGSz6dbEHkW6jWQp0CMlXANNUeZfGtAElfWDrP2XtdAQt/yeD
irvqWJiT+JrrWgR2twDhPipK/tVWCmdPsjhV0ieLreAkD/G49mCKq/7V6Pq30owisM+p1Ax1XviU
UJ8kKcZRd4nfN+vPeK36htAHZgGO8ceJv30k02uRXxDCxmZ2xPwyaZ81Tn2L3Pq2OLhEbJVC4X3O
X/Fe0Iiwhycxy63IhRf7HxogijaQw2vgOJhEnnAkJRhyLyTUBO/vnWBdB2IgnYQrCPkpf72U9OjR
69p9iyqugwgfB8OKPsBz1LqlCGxWbYxIvjevvIdvtQZZ6MqWc3o4BAwnNFl9SzP/dSPtWRUbhjwq
X16o1yHtjtqNDJ97rTRhDBDsnk7c9XQT+zN47P3rMpD9KFrxFOvnyH3kbhVmhig7ap7RyqXjeNY5
ucG94hU5t8uU1uTo2nbgWE3CKJdW0L4uyhAwdU0o3WR/WLwVkEYqQ8dVt7J7pRWPlfM5JukuptMI
vSyF5qvfIUbqoI0ApxWfP9sSnrkfsRNXGTjKz1Te7eIQqKUKwmSu9d3ZHH3T2WydECLpBJ70m28N
ipSwXQiW9ZDXw4suQDx0pkNBkzPz/9hf8ki4dzJTXIqRFloFXtrDOqq87YHKjR4WqnVGxXyyMiEz
x5/TJpeOX/q9JZAN7iGyOBPxxnTycEhQv6zy6XNK78IstORMOSgT/YvGeyHvBGh2FG34tsYiLCa6
3vzMVeeNq5lmAZne8Oa0rA7lv7VClRW9gxO3siEo5gOT8dehF8+/sFHGesIJGIBTBBoNX8ID+86R
yDU1QuA1Q1Y0iYhbx8rzVC4WQfnsBiOwHzHFD1Ksb5vQQfXCSGuQxwLUzjgf0bFSHhxc1FQZkuBF
3+ThMM52m40oOAc25luCPxLP+c5wzEMAGquoj5LfY9aAnU/skEirlScgsEwl5rvzjKkDZpNBl3l1
e3xcQ3SkbuIdHgDWh4sKMAioIJzpveCpTIr49ZJfiMo2HcHOeptPAuUOYlyrp77L74jleZlof486
rlzYad92TkbZ+9nYosBmVussNcXRWF2MlabVB846HwQJ9cHTF2YD4DBJ90mmdrkKdaNLOx8kzqlR
iktc61Ax6EfjOPay74UzR9J9WxkACXnoXVxJWx5iuU6yCmgPFRgeMr4Bv9t76WaKxxek2LmK3Bm/
5AUxOPWsc9GAZdqFqWS0gRQaKcthq6TWwHO9ZiIJ9q+kppv+llMLE8h1z+VGo1N6GqitdtqAq8sk
6pCif5PEgFad+o0TpJOIKkAAQTefE0Jy7pTRpwRFR72jP0+uzEaua5k8KCPffQ2Uzd7t373vs5he
0+dsdLO+vYf6MRFqdpcQmv+f6nXhecf2ZML9tf2S3A8ctWhh7FjlsHt9FTxQNUv6yjeODjZeg8k+
qoSpnnazgzguFqRb4WksSTHxeJn+WbLuvIMVnZFuVKfu3PIcJDAlbyTb4VvEGqATo9FT/cUJQEk9
y7CD5BaBLqjkiaqu58urWFwKVyL1c718fsRwCbUWPY0v9xYinCMXPlZYwLXVL4z5D418D9WyvaqL
xWJv75AfXn1H0v2tExo8NEsZ64nl5W1fq5+LCxFgWXs1m1ESID6k5Ru+K73RZrpEIOWcEmOlwx/l
lkPSr+8j4PwqSRMk1JigC0IN357J+hBRZO5NYm3yf+RF8+2o8M1HXX1TtWbjO7rFS86x0/8YMHHH
r9x93/+y7qAO71FspMhmJKIFe/DbblikQ5yjeJZvEjnfNUVCExzje4UNc9MTOMgtjN4UqpbjWRjs
JUtmt2VhVEoGG5Pl604Dx8ps/YXY4ClzJWLvItSogcbcjUSnI3LEXeNGBgqVK++Xk/5koH64Ghb+
eZZ1s0lg+ekWzSSDS4bnJx2JNXJ1figu5Sl4bxxHk2MxH7yi6DYlM1dW5hlRzS6v9i3LmNCGXx2/
ei0+CzofylW+ktCUP5SXz2NeqCpDZMtmyqM2h92yCGVhjidk5ajqbNH82hXY4gJkWkN/zWZ680xE
t/1IYA/woa/Aeu+WBVNYmA2tVXNESAJZ2VOtaBvFZ+dJz+VV7llmSRE3SXekgVxgaBAgi8a16iS/
x8zNMsvIYCgNDsXiUGMAPTomj/ijfs5Ml3NaOq+DcjBPhPYHj1Q5lAOrk6VoGUpe29akxMFsg5Pj
npo5bVQTeydpY89F46tOOIlEwfOSsdHjTt30UIig6W4Cs3V2uqp5xwwuMDi6Z393kcXoy6mf+jKB
PZouKuLD4uuEVlTM8C9/+lFRpFuegQZ5M8qbB/M+WDUVK50uJkPwj516wIT4s7K4VZyz6EQf1h7Y
boZw3EgrgaLoNYKjlqF2/YzPyExkRWjJDFKhGjavXh+3sS6I4+g/ZKIPwq7fFeEMV00ccJtu13da
oeGL5x9F12IPaDCqB8aNlBsqsGjaGogtfnMsVNOja5egajpCX1+GDDb808M6Di4JcRvmWK2dnmRO
NJqEhFvccseFhaSzOjpETpbE39kubYbfQa4dNA5hvs9Y335OBmD1YlmNmArxkpSnpMTcMZyjpMyk
jxmya0gdgFh9ZhEBCUFSY8YzXV+DJ3GT0WHIREYN1apEWaBULe0IJlq5/EgoXVpvgX6AYD1Jg4dA
sHrbP20dA2EJIZUpu4y0JH53oj4oF2ZbVOn32/HQiJdywKGeyVJc6uJOZN5NEsal1IfDIQ8+alqp
fsfXx6urX3/vgtjmdyDU/kLD3YCXDNwkxZucBLaMrl78DD2QW16yULV938NZ3fJ4qbChTjXYFNZP
00VS4P/f0qTLnYf5X4dAnn9V1ObOUqJvnSWxjJYbM7HdHquR8cdbLopsRaYZc+RQR7oPwkHv4aDt
wd9fokDtxnCuzmHTg/AZD5JSn6BIs9ADA4oubgdlLGYkn+otvkv0UIQtuHzQ6dtNEliXSfnAQx1R
wSx69wBZcpC3ETgG0r+MexN9EAQXvUxT1tRH/9MzrAd2Gb4RS8uwcDlG1uQLoj7g0n3kGVug20Ma
qLLKWEVP3p5BhpZX+bIilYWG6ijC+j3sH7YHYUN0q+fXLqEjUE1fx+MBzg2J7GjeOeo1ZjbslDYR
VqEmNKQ8ZyhFVWfe8fQ30PUJqfQVzqxCtoaMjscTIhSddBz9BFxDENuOUj5apbB5CS61lQZOeTNm
kL9T8sHH4e+xNkhN1+kRZZzkDwhhmbHid6NoWdnX7eBabznSlqSriLVTjyKK5oNb5OHjUZkj29uM
0vPp67uOHUWIWqIRBLIe9Vvs9vnhxvtLPS4XCUU3cC4SxpWGkidsJtv6b2j+ibPV2LrUQSiE9qZR
JcGb/BZ4Hb+QZ4n6x9/ZHrHPhKyhvJjnW+JAuv/+CqRoZT905jR3VoNb2L7X6cEBrVKLWI3z/Psh
5CygVbEQDRxZ1NSLYxS6RotU15RjA4EougoiEU1Q5Z1h80u20mfUkazKjraxXRdGX4KjhXBd9hhl
/sUIL5EJ5B/0B3cqX/EnbPiZ36/11/rvTwXTHTvH2ZPV7weq/CMOtGAOq9yYsUjI5rpdf+8yqkJB
QwB4AMzl9N5pSiHjF3wcS8QQnUtSBH+vADKnUfm7QiNuex4VB7wNzWS8C1BUPTn2XQSH+472RIjk
eN9IcYHoAdcz/kbCN0uE3QEvDvUID5atIKGewrkOevtxwaGiWTzGI4gEqhbx0kTJ2UmfOcTYcjYh
EmmWWpdlyleekU4QOfh0do1ViaTspYG6Pf83lZUP0QrHa0gqx/D2RoQCsoL3iG9Swyb2nm3nYHsM
uDvK6JQ3KOE7fTFaqLZSdI4l1+o+eZbFCaOv88jGns+e9fUjCxZx2tvRRJdcAr/LU075sW/NnSRq
ilQacTAa3wKYkdCIsuTsVF2KTGEA4oFX3YN56cdkRX8cArbb9kw+uX6KuCKvqqBvfctrNasYyJyG
ZbJY/SUdXDfQnVF+HnG/0m/ytS3Za2BDpK1NCEy6rosvFhoJ3sr3ebu0QFKGPm99lOgAs+NR1fLK
cjolUgOq2jiYX+fRFQRM/DJKw3RN8ULl6Y+XwbfpCiF42WMQxYgkprFf7xlcMZuZ1HTJ7f+leAVt
oPLGMWi4d90XdTG22xzoE4Zj105OIGMog+jD505rnyQI8peCI+EpyrzyQqVt8gDRVKShJmqfwGrF
IsFCUmB3sc5a69rfPjIAXFkwYB8RJTFsmaoHe2SSObqoT5JsJxfC5IVEQcRgYvCQOKA2nQLKJnHE
DvBpbnvoAYQwXr7QQtuTMwpZupzQAxgExq0xVIlboaFw54bN8i0w9zyud5EXKZPRp+o/sFTepwLC
5IHbBHrCcLMxvOjzrX1sHdto8/elnEycykLc2DjYnvAlX0T0PHvA4YYtSp9fhFYgeo/FEcWxUAOT
MG3CyngyzmT55o4ppf4fJyGNRItVg/R2KTKBu938eF2Ail/vKvJKtnjHiH37JIpD7mSEu//69Ynl
axjHNv/N3YJVbuytLo5SjnLUtmRS4kAIRf2q67ajyS/r4iFnZ6iyxyWYNvyOPrq0dctEG/WqnX9O
iKyWpKQMrwG2WQqTgVAdrNaxZpEDv9zeDZiaNHevy5bmPq9riPiBg9SuUXDsM1mcGAjQVXL6E4q7
OIKOWCDgU7NX540K9DktQh9nxqptrUCXhUsyL6PjUBBmUBfkUr74epDa6YGbZ7P152nf6Qo02wMk
fdjwbKdJR9ix8T194T1yT6YsCQOLCU7SaOpTdiuw3So5YygDWmInKiST9yRDiTziNd04+KTt7r4C
bXaE1cZDtTWU74K0c4M7ZIjudDgPJazsJS9UIgXbRGMek+6Ph0Eh5dfzkjUrbCPYRbARJ3BO2kRe
OLRh7N+mjNtufb4R/TaQYmPZjXB/HEwIbMxgkGvBGcB1BVfKxmv2oqj2C+EwsaSIXSl7veNURt7g
IYDXNcii7Vzdk8AFf6S0lQS7lgCc+uKwG/FTavV/NPgWWuybqxVSsSqyrW7Z2taIBXlhq9imjWVL
T6/jmA9psoTLmcR9MC5Eh2odmDLew7BY2WygQrf7nz8s3mlRXhxbqt7XLMUvI/WPQcPWTJV4pKwF
vzKgAIDIfIEN39hgcFUlegNuqDum+X5RCCcLLZQ08TAtw9rPJJXOYHQs97jON3fXod8cLiyK/FVt
XbJum7Vmzr+FPnw40cD6GVz/8AwshlND+pbaNVk3gQMJERYgR0bAeiCa5kHM1dLO5gAd57RQeqpx
Bk72/NTc4H3RX9Nq24cCjS9Aq3sNRR1cYjtCTiKHihspgPtZtQ9014l3Rnrv8POKS0Xi92jcH7qQ
UI1piaembMf7cpX7Kcnt6ZruBNo6qP8aC5htsV8tSjCJV4MaZDRXTTqNFPUTIByJ9syXMdh9ECz5
HTSl8Pw7zqJfZKIr9XZK7EuWtIizSeinPY/Rl9158Z9MTLG0/OOEBNv+uF0Bj3OexGeCgbGwiVba
eSNH1xYYDsQcC4O5ht7/2kvrdn966kZIQ+AMt7i+7JKJcdLpPx0YPlnss5cO01oh1a4d+GA1tVxo
dmonadU8Z94hLJr3WGcI6MsPNg3eYV+yQHlw6W7aMtoj5MrfKqVOBJUbdyL5KulXGgA3fGQyXZUx
EjV8byivPmWolb5g/2Y5UUUiIKu/G32e+NqQzcHMSvPjAMtMoNCBq9X0Je8Tn1MKUz0U6QXx3TBu
/0aiLdcsub5cm+mxgVHJHP0PWZFuYDM2Os1nVPMui2ElwGFCjxFp5B0ASMDFZJghQmUEXPSPGXrD
eZkR92/zE+y10WYk27qhD5eQlnVtlHeiDPTQE57AlYge0ITb1Hvogf7Kq8VSrawsi6OCcrtJSnpU
AjkzekA/R9vsCURBKuIREhPWeLN8KKsscWOBGJXmD/wy+WyqdatuEsxbLnzdQbd+9heH3sS72FJR
fk35cLvmPmb2rWiBAreIJlWft5Yqv1gNojSL2O4BCUNEFsBXiikQo707YRUJQkgh6A8/1FGMR2as
wbaYXgNPRkWVP6pnLeE05T/W7brQayNUVY2vgpHckiQmp8cXQjAoPQy5w4DWcctomK1iZH9qPRRr
9ZQ7qkJb4hi+E8j3v0Xl4zkpRMSI7eAK8E/Tspeey5vGk4nex2TUr1Eu7ERIMD2gXlH3UZW34GIc
h8E3SQgLX+xDOcqWLHCGlu1JKEw/JZvAP9LStbVhEl7xbgzw5cI8oGi/UVdRrDPWQ1lSDHdTWafY
4clDSeeA3/wbtNHGmKAONGzpTo+KNtESloPdUUA4nnsVLS87lRJxgBVEWJQ4cfHAnSO3Z9r/guuf
d6YhwmR9YNAcT3QaWLag7ujvKAgR2XXq/oCyYiqKQIQZv78aQbEZd/QboIck/1v54d1bwSPfiPeb
Hg5auKi2YNC0iNJeHW/FAeMt1w/BOjAyjKGFuu5wO49ZkrXB+mnzlrr0kQtajxx4Xw8PuZIc1ibM
mm6hLn9qUnp/+5epRu2b7MrB3YAnt9vP77zSAJAR1y7oGT8dzEGB0iM6donCkfgTPP9RcyNw9s1p
wpSSeMRR7HYsj/7Y8iGkQHYJh4+/oPs41lz0ZHzIF7UAKNoUgNPiB1HomTuB3hkaRqTVP8LgjmMb
VtVXs2tGxUc0SCalapg5ZjegVOYZ6Wuija5JBkBgLCWzntOUGZxJEJWC1EC3wo32rLFuufbcq3Z0
bVCYONm+zvseHVnNoSovD3PQVjmro9T7CyBGNzM61PDljk5WwZcTjt9yvxtHmjwFm271aJ09Dtb0
un0/us39SjiZSj0hNoxn5Yfm14qxr01hjKhx1lDHlVWUKV1bzuzJdKRJzqWTiGw673+i+30dIZ2W
wo+rOD7OZKFyW97YJxRGjxg23jv8E8MmyMcIyntr0rBuUCaIInt2Z7gJqcX5eCRr+Xj7JUK46aro
Cr5vrZyUeEShJ0jtU42/jg0SuUnvAdIjK2HaxVqfpjN9RKRq5NVxHJNO5A5yzRxvZUdhhIqSJITp
mInn6IkLJF1z+oLvKRsLhk8btsnyZKZ1p/GRlKsazcmc3xYz9D7OKNTNcsxwp3cwclV2Esb+wSMs
3wExSwcw3C33Ars4GIH1wzWdSFtdNkF63n8YSWrFvUmXWiAes3ZtOQAIZmnoQlRtniXHcfAv2k5i
hpCslfgCnmkmcr/lSFA5542DVTyeLI228lwyzn7kwRceIvTe7OXnEADFPAB3OIgrs9SSEXqbZIEn
UlJKNBs6rGzTswA7Hbjkdqsx8pLB0RC6jyo5/zzTO6dIhmH6KS2ILJ8Sr4CNX8Wm0GzWSw6nk8tS
1wVrFjeIpLdNIXTEw6AFUcuw0O6MvsEthwh/+dIyVEl8PYkrVITzRCrnlJXuzyRuDerVy4dZUEx3
YouXYbDkamMYiWWd5b/X2l9bdnYCPnsswhMW8TldbFOSz4h+hvMmaEQ1sihNItb65FcWD1texwNr
lDfWiov63oDKIm+KOpOr4nYvdHt1khpmfzwTDIrpWo0TkTi84RIE40VixEP388pBd3VYHlIP/Zxf
WB5xnchMZfET2jOJ7IfJDguQbiG3X5y3g7v1C857WhAB2UpIMWtZcQ/Vtlg3rTa4hvuCetesrDBj
m+TrOWKveY+FvTOrdwEQZNDmAt/zl0Mq8esZVImPFtG7NIvn0kyvvMAmpkfh40BsIYKiSyrAD7jB
FwC8MgLL++gG18C2+E3GC+2zhE1XJYoS0K0rYTqi++eku4O1dlyPhSID0/yWtRIKhTD9d8n9V+Wu
RW7ofKKfkEdRbyxP3s7CJep//vMIu3pk0KHUPKQN3V5BXsoM+cTm17bpzGO4iC0si2AhGiLiTlM/
XmNlitzZewolcC88vJ6BfofbFrWJSNw5+F4+SnRXUwOnHu/Xb/ktE6VhuTrt0XUyoSjjUssKHcTn
NVUhHlgOfph0iR5xNk/LGCiCNj+jt3aWkc0XrqQv4g633/hKbKKHgRFD/jW9+unHC+LxDlkBctgO
4E86TcYug4gblUTZY7o9oFrV15B59qp3pbF/shyQjFfto+gpwOF8+A7jtW3G5nESXTJvqrvbRmRk
gmcnleey4uhwwum/l4aHmbu3SEqWCE+kFWWifgJrcmahyqKcNe5+RZB1WsHeMI7XL9XeGMilPOwa
ddOVdMi1cRcWaF1x6wUSkNyQGfpA90tlAjqPWp+1PE6KJjAxl33zw1/ZXGJTzsusY2sZdadxUc5n
2Xs3SfWiPqtNuf4/s17orMFZabBLvahZ1xx3+AdBmzbKL82aky0n1L5Sz1TW3wHn4lW1PQKctAvr
2UwmBDta6cyJBnSjbR5eJW5ZuBP7Bd3kwsV82x+aVHyIxB38jjmOj65inlqbkTqfng9j2lNXtYXO
PN7EIrnf0J9YlFIi0Q5Oq9zIHRLRLBllp6yPdGJE0wEBy1IdeEP21f4m238ajNW4ndKNe4dSIn9g
jts+awg7z+vEZz1vsxzpQ+XQnmtSBjHaSvim5mL8gohXUYwvwhKh2N7P8VRlK3F0PQ/g03+zpYOL
RM1kBOHN6Q3onTJYJUzvpNIWxQg+RHJxO8Kc1h4Ca/U2WyedC/FPnar0aoRYfWh/UBGDiDujAYlA
COQAS4qExYxBwieEZ4U2JVVLHRTRpdpGYQWqoHZBDb0zeGKkgxzv8rnj0Iyu+jSQuUFyHcpyXo6S
zYFTK/LGity7UqZBWsdEReGFOsH02vFPV5e95VByGw7TmOMS5LGCQhxJrYJym57/eB7ezHSfs8WN
1AbTpkNkZ4eShorSNEGWHRCupObKFxjgozVW59JujlTx19718Rsg8BvnmciKTEHUzbJLj1Xxmic4
BkIViU0F0rUfLt+tVuXOdeFGomDmofBACVkGg+Q0mrV2r7zmal2vRY8TMuiK5r0vZ67VUexm1MVm
TNSa+MhtR+8VIS36kz0im6d7bloFNC2YZuu1zRWnI2yQu0RpPIQVts3nRLTHKMhv1GS4YH9pv22x
DI96JZqlGnePZ/J81dvdPQyeF316V4FmT1JlmuJM8QUOyok79Mrn/Ik9UpiwstW8gLzjrhjBvJgW
/iUsQBMuztTOhN9ekD3U32bL9so5AYOQgHMXrSkjeNb3AID5rvP85NufdMDHNoyYWco40+1uxKOg
v+5dRfkNWZeKYDsQQHit7urlI4a4CcCOUZI5fk5yKoSITJG+3UJwP2RX5cK4z5S9+lqBpJcLzG7Z
yM/xuUxQ6r1TPsHOtdQy8cuuqwxb1c3ZrNKloT0/mYW3/PgthER+iyNGl0uYL2UnrkyKLpEDR7yH
i01/SREydF5Fe4a5vtNHXEii14n1PUTN6wI07mfmDEqyP6l4i+/FbrbbxEKC+oJboIfBpQBYBxKj
iCL9I63zQrXmI25BRCtW/qKSq/NwBCG1HjRrpWwgE2XW9wD5qmVB5rkzoJclTgcaNvVRfYahM5kc
qt2ROgFKbJafM8Tp98cgTtZc9X8oa1tdrZkObZy8q8qn1Q3b4o3sbZct6C55Winf4xLIh9/ggiug
StvC10DCIXENVPQvMHv0745oIdcaKE7jLOnD3HipgW5BaCEZ1Quo02zYUhYnJ+L1XZUl4n6nnPUA
FXltErPRJ3CzojAMfReA0by4aWYVahzxArC3Q6wrqha0j1kjRPibKPqTchQ5orFUZ+ncrG/c+dSi
OSp6oRtDjE+h4o8Hicz54w/w2JrlB6I7yX4VhH2VWOIM9SP71CleTUqJZIPyLnjmWxqQVHepMdUi
KwiU2708IzRpAzFD26KJiM1T5wXKsB0fF3Uc1ibK/qp+dOaJ5jLa340/rDy3JM0AyUq/uI9XtMY1
xLeQt243VVZHHu7Q9cIa2sZ6udQDQn4aYjYAavZU0XvhNgBoyN0hRaUwykRmC5qvT714nc+NzFvJ
eD7kxxD9SnDxByH3SPhKbKHGUvfesYW9T//y1JNyHe4BFLLBzj3uzJLMcNSfvgSe3ZzqQA61+67E
WeomTQoWvaejapN17ypJ7jSeH5SP4RRVfdbdy8ca+UFILuh1bMi9aTEWRNarlRlkMUDwrT0a5e3T
A6ck1qqP1IRw04Ij2LajyrU19GOpigHJrHGlXS1e71bZ213CepO3uPRY8oa/JnbqcA7iH0SNaeaI
f6iAJxJyO1HRxQuce+w+62RwCLZoq/6fxre03LNgUX8be5wqEUFhMbU/sFmC3hUnWtwzASHqErP4
Oda4BtuKFzfvLpHpoSmUDuFTuRpLRnVKCfZvLP8RLuXUjJGoRLuB44nj7OOdRhEzRRPw964PYlob
tBr1qrk7yWkRLHR/CAd5qyAUVBg57Vf0QGY+LSiPkBiEBYiaGi4OWmpClaCAYnztEikd0zbvTb2U
JHU4YBJeyRkfHjimeSvXunlDmKuz68mlPeWqdlo2CqWyz6rMwkzcHt0/X1/98pvoHrM54ScDeALI
C8XnxRScT4CCAeSl9BlCZel6z/bhA7oEPkEa/TFX02PZdVPjrt3C4LKSQUJt7pEtExpmhzreCGOk
Ge/AGZyYtjGq+CNIbGYrAzWbTbpj4VZUyzGJ54iHM+y4Gk/KtL/80MxBY5SdTYKjTcOD7K70ORn/
iVBF/l3nOABKKdEXrw8RNVHLcPQFm/KGOa4XL+XrzgNopcbGB9Dwj0nj89n0cUGUyB9/JFh2LtOJ
8vqEmoPJuiBoA9Nw4eHKRzZBC0FfCR7YOKvDKJfCKZSW28TdX/SdcrP5miW8HO38G7NwThwk496A
jcFMTb0wylSxGa0bVnJhsEMYbBxZ35m6j+wYC4vgbdkNihT+94aH5ijWYVRqzuZpvy3aANwDH2Yj
XtfJ2K/j8+QOWlq23mtsUSPV5UEqP/a4E2Uz7b714Lh5l6XRQce+1umwlVNerqJzq2jAPY+xpsUO
1w7LUhgTQ8feQXDH5Ob5FkexiGDDZxR3iFOftXvG5Zvo6UityU7FLUHrSwVseHX5eDGGtRKUOUsk
0whu1s7XZUvtk5E+2YyOVZLdpQVC/setNu6yIW1o9JGffiJgVaNasXh46uE+Mh3EKMrEIZ5w4N9p
jEBPaJk7WxWd3CWB2VmJRrx5kmeo+s0MFY8P/Sy0iscM4FlNGKKTokVkQYPVEumAm/Etvzf/aaOL
zFriVI1zzIDD+e2BdGg8tZvvbwaTYx7d3OKjfqZqt0scv87rkQ0lgcyec+06gMALG8SfeT6xLUIg
ZGp8/kjO9Y9P+OvpZXzjG1MUC5yS089rVRLr2eXyWi2BmaMODa4leMoRazuYFprW31DSkFAYznFL
SRvMMYXMLLKt308/XNBsxd8aJv+0E5pcgmtu3yha1WJU8EV/dpHPYVc67g51c6QBCk5zOrMWkTnt
AuGoNtxvruG2j8tlckKovemqs/yWfLVR10c5AW0Xbf9Cflf6+U1COgu/PvAmEO0Lkul8zLFYKlkH
R8icZ3Ytm8LhEKuE3IS6JLmkVvmW3W1F+YC/vlxAN2VefGcIDt2LvaQgjiKGMCI91FsTp0joTi9P
UmJJg8oGcZV3zHaen6cGf0/C6WQKfQYLWGDbYfQiVl3nIxbre1cPuUOXaisaw/rYKxnAH5QEGj2g
coMpELk6mp1oVyv8LXVPuoeP8TPVY6FKuXq2tQgA8FWcpRo+taPwAxca41KGSMH5daMgY6CnVwli
F/WsdNQARNcx6z2PhCHoUVAg/+3Gj2jWOmfHWx2VVwiWWT/CZUMfmQSnD1bkoZnWrkiJECnaFZtz
DO4NNhSK4zZ4spVGSwNvp42sdHmBnim2O0PpzQUKMSqYYA4yU9soZW1vmLqJKV6PrbI7KErMJANA
kyabgteDNafwrlr9CwrufH6+zGmdTtk6KaHYRx2XXPkepSx7uPvgV/4XBZ8C/7ESs90QFu+RHzV8
y0eaui1fCMGZAdk3IeZTI1eqkjLeKffL0rwEo1ANJp/YUi08IPKIC0t6LCtwwyusnjLeHjF3Ly7M
xv7yyTJ0TNwGCeKG5LLa982j8vaP9xuPFD72njNiR+exSLTk77gb43KbL0lEMw2amvkn85oOggdT
Mpb2bPKSznkIloK01imp4HKtD9OvlfPoSELuFvPQySFpzIdrmd6TCOEPsdOXciWr2kyv7FTpMGd2
Nb3H0d9bBPhAmkQ1GFb1eMUbwtk3+ofAuOqnP676KsYHvmv6F65ffY/cTkKupSPsL0lp5HgM0SWY
3no9RhgjwvMV0e3jTxaBU6LSselJuqBmJVuHta07+u1ckoyYr+fvupcXoerOfcFLBJeB19uBWABV
yctW8AIBAsHevqBZXlc+553/9EKn6dYo8fELaTrVMKMor13ZJVSfiSHd9mTeMQKOK85uEsuKU81U
e9GBvHf+AV807qbEA6i+FPe38NG0MAqWftiMucQk9BF6qgkasKjxFOmY4vcVWyIsdfYRJfAj7Y6u
m1JieSlVB1/QU16sJem2O94PNt0Wu6jGKUIQoits5cfHGAgr/ojQSv6F1BxtaLJ0JQO4bMSMTcgN
UKmwAjauwtQp2VnOqjDGYEE2GRUd3zOJ81X1fBU9uq0bz4VBqE5PENLFBPFVkqJ+9QkOXIcdgy6m
0FgrkJ3H8rMrQJPBzLZEfVNBfJdalQ1w2Emf0i0ixmrUjfY3bufLYBjiguhdUfsUFpq/iWk3ea7Y
PLu5cN0lVC56FGdp8aYc2g9P/LtQdmm+8AN/leHKLwbVEz95vv/frFWlJa8LM8kLCV9S12eFPa1u
eXXT5OzDrbxO6nK2Kepher5DyZX4GPWv3Gj9qJtMd4qw0+EfgVVD3tlKfPyawmnez0Thby3qrxGb
CygIqiPRqpATDStn+umWSivR3nhNzD8T+EvDrP6gQ7hHiijx8SBQ4SstoZkC4Jxi5pq86ZVjuA8i
M7u2fV3BeF82O52IiY64HCQlBRCA8Hw6NdhC5muqyB5aSyty+V8YCNoAKVlO2oF7FEHSyw8jE/WV
Pyh/7sSye9S4KGMVcq0bI/f852m0RsdTlRMb9w0HQnOuXI6KqTCD62i125DwX+1dtJx3ALePvOem
gel9DadR8sb0dX8axurKaFQZFFbsYP8CPlzoyW3+WaAVMPp+Y30f9MJgF6bUJRG6MORhUOY6XiVy
Cdk2boLUtounLWIoGpjNM22YKWIcBN1EefFbBIQrXTGDQy6UgJYfBaDggOTzXvnkjHFmMPDuhMta
tnDo+vivVaP7hL82VUZaKMaVlWM6OcAPovYbMriklVL6vKvPqe70v0L753M9oDE/zy1F+QXOlWbe
E9TUF/Js4blVuWAdYDlLnxozBf1nMGuCDjIQ2m4o9qHSb5G8ndnrU6ndVNvwbFnNx+pJi1A3MDMN
kuQaO5tP3i/hDvl46RvHhltdHs6cjIL5IJSoxpifXQ61AuSGQDVJa8MLMHGWKxWiJ6korSHQkDgw
ZZknxs4Rwi+aJiyJToa3Hy5Cbwq3UP6kIbA5A33JjWlBdVSEaLNuQ4sZqam4XS/RheIRozfBASxi
Fe9zt7rTgRRFB0nfXlEPPzhC/28DkH+doPUXAmx+FNS1v/ifNRriDm0exdpmKf2C/1PjhDnJUZtX
VjswNa0SGJCvjo+terTxrbW0wgsKdUeyzrJuudKsyImQptCzh6EzsZM/QI7lgvN6eFdo8tZV0Vvk
wigwcBIFVr328knhQEBl3x2lKOtl+Ij3VZhrRrLB1QhJv12gEp2PozcGDK8R0UtlBu0aFzQg2LrQ
3Yl/otRChiK7ZsL6hFr+CiNWkTblXiwZmKpVqaBl1VCbarkf5QAG3dCMBUzU0giVfAogLM8a8Ph5
1bpyHCcKpKJ/6EMqc/UL+Ari0few9EYMA/8HHGqpQ7V6mG0wdYEATvx+kiChB8k1526v3NldFBhM
jeqBv1xX6dxuXWf8K18c0A7emZRbsRz89cXH2FDUtVu5tAeweGqZSlf7c5ViTQNviBdJ4Yf8Qa1w
DwP/c05zzOMZ8I7ENzgLQbg542UtaMailpvObM4suNxtFw0iHXGU4DQfVWckVDXLI+tc1j6HED+g
zdqL8eBIsJfABvGomELUh6p62FfJVKsZszVb00TweeIF3VBR28y+JmU85G/2ofXdHANd1hKUXHfr
IqMp3n+V9+qBmGsuIb0qolf3o881WOPnfEHWN7SblcppIKPmDjpiaF21h/2ajzAH/1C3S/cy9Qa7
dddKLN3Rnj7RUlVmnoRaT8TZa7mx1IsRrgG3IffIRWPOj4KJxUYYE822vdnB53rA8KEpCMlDgLS4
wS0GTVOFBCq040ARqMHZ5E9nHGy2qoQNhgOLmDrKx3//yG3cReJl5YgSCt8w+avWrHkXqtVGkvtB
+G6n6Nj5pTCbEj8HxCkF26WDGe+e4dbPbMky17aze+qHBUomIn20GCAWb9fS33NQgRvqUGIHnaQ+
wuS8HhdsBSn+4L4heOnbmVUN3O3hUE8RT53rRGJMDbNbTMtAvzypXveug+DIds+w10G9Ueskj6dU
cPCWElX0fjGgqzlAZ5b2l5DWWup9KY761A3vejyjeYxQBGuiPn8KXLfmLVjl4Dcus7qPxhEiq9or
tu09r4qHCIvbgU1k2MTOcC6BzptBO/HSsRPbCrdmu/UphcaAneXBh1NCQPvjBww0AuPr6vv0mvmq
wdIXveB51eqlZfeYRDg/Zes6/ZNNrSbL06yLCHhQTKgVrN9rU97wcw2t2zmOM5sfzi5112txxdTm
UQUsLWOq6LM290Yniid8NiowRaAuaM7X7wsTkBZHwps2WoOesH98v8na+DzXmeGAfhRq6/y/GZ41
kzBIdZUcFSHugEMSIUiC8DwvuLHtOHAT8LZ7qMJlElUSE9u1g58NM2PqR4raymZAPpfMqW55IQYF
AehG8SPNetFisrgAcSzuMpjbQTp+yo5Zz9rhpD7N42gtRRzEVBs1cmeHTwOEuMA5XXIkQlUsbCXw
ye35r2Kh7tGm5CCruqcbtP+DJ9mH+ZZqQHw9fWBlCwpEvV8NIwINsKIfYwP8L2rRRt/CXOrdCBtm
z7YEz0V4SBsw35jtd0nOkTEx/putubbH9d7jh04M+ueNroVrRO22xVH3HALd8F8bj3WDLJzwOZ6D
LKbcmaK5XMWuU9c+Je8869o4kkFBBg9T9hqBdxz3W69zmn/MGcUO3uoQisPZMxNjVop1ZXxrMc2d
sysDxrFEpjodIMEizK0EAIK+CuF1Ia7EGt/vWRs7EVNkFy44ZEpt28n8YiPJI+24IaSOoIYAuNMh
2EF3yBK2qIU6O4lAu59NvsMSktFVYD1tQqBg/Uf4Z6AyXSzN3N7LnPjfLBAgeUQXI8j8HVecDgsc
AJbyAB4ce3UyFrliXFFC9LKdVhzj7Y8TWKIRmEo1W8BcY1OUDli/HxF/lwDh412wwMh2dMBXQ2GQ
ZlHLQBaw/1tmfT4nVn7TwFnC+hBe2opfuOGQtYK16xu90aAtCV0NPr/nUN1jBJnQU485mCw9dCyh
t7gOYnDd5rx+g7MqIN2Lwnbx6U9RvbwRtXPpTRlxebqfDUzInyqQ4hbzUty0NLI+IHSXfQsSGtnU
fAM7Um2PTkUN1LuHCim8YocxzuqUclWGuY2lAUxD+Czw74E8JZ6qFclOrfE+Uo/6Awo0hiZf6v/j
A1iCI2RRlFpYbuxwj4DQsfPJ0oLwydIXM1FW9QJaRGFcPZpLuWCXVJaJfSLKrkdXfVRTj0jbqDlQ
gDlRtkq588IUjVSj85NOCVV6NkJgs9xKJIbsQzjwQeEQSQA4leideLntlP9mjn3iQxGeMzG/84bL
JCPvRQmL3UNRt1NYuI0IhxqPaXjEzb9jLDyGzOlonXl1cxaoP1vtRRO0B/T0oVJP6rBa5g3Ey7e+
AIrWEJiNBrJZAoWlgtOKZydZI04+R1whwEGTvdJrzu/yyca8pN0tqSwmQ8FSYEQmwoLXGdbvK13E
a3/7uwwH+iBRLKj/MWmwOllSc1JgSjF8f3oM4Tz9TmB2nip47pCtHj1IPD2gKiC4ORNoHVRkG8B6
zkze6oqELM4BSaxirDMTkC83/J5z/olsZ0NXD+vah9jl4mptQVgYGqRZsxTi9G9dwC7iOd0BceZF
0t/VbGN5Q8luM1J4Udv7Tu6pyO4ZYsHkuYUHBKeXibqe5Obz6s/YI3AYFfx3P1PvDwhh06n1gsxT
yAMz2l6MRfAvK8iyu3az21FeJen45Elb4BGK3Ffk124/H3x/9HPbRfy9owzwieeRKDI1SwydirpJ
vSd5n+WzzLfFg0uVxQYNxugWS3LQvszWtpy+q2g1heQOZrfJQMSxegCDlgyTNjFhNJlOKI1cCN+c
06e8u9K/UZ3/JrVPQ+jBBU0tug1Y2qdWtsgpacjUinWQ003Uzok4EW6hvWh7LZ6szwG7G7msEvk3
0mMxFM0JulzIy+9XWgQ4/+OlxpdFtFO/pa4pRcyY+B46SfVTGNMygZ2s/jZ8dggFNtvrjVxcQwxE
Axtz8Im3PxQPJhpy1muuQiLnbXa3rUG0unBTqDYBw4Mc6KDezq92VQIUYnvIsohWdFUQtT59eDKN
B2GU29LgpbUh1tFKXUWtyjd7FPTPPq6K7a71LF3Cg5mtUPk01aJqQONkfTcCRbWb6bW4uOipiOOI
HqmIP9sZlWT6aBdHwx8nCXmEBLPBI6/Bfm2j3PcsWXuEjsZiTPPnHeSSA5dLajWmqm8b++/RDQi2
Dt96r3zVc94KDWBV/YL8YpDtW004mtlAMSSetyVQC5GxubV1KjO/VyRUVKeY9D7cIhHCuuQob2/c
k7igWebPKbSyp7mDD2g6TOASe/gtclaNek1Go03SIcegMRDYPu0vE6cRclaGCVt8Lg0djci/X5fm
r6xYOw6Kg1yGwpIx1voAqJpBiOxRZAESoZHYv193kQmxo118MIHCUb4LOCP+NJZckTxKIUBuHupD
7h2wp+vFCV8/tbAEYTKVaZfEnZZBkuPIBSbcxWdy+BPKsJm/0HRsBgXKlTqoCQzr1XtCFqoKpH63
dLRP24lf4wEC4O5PC+nmf20Dl2fCJGsZb36gobU7jQRs6ws68mNHrsZMF8CBmaPecs1Nt+hV3Gnx
XZFQC2ZxFlwnc1i30Xxq6vdTt99IDieeWibKEqy8IFXbhoNZSMZN7yCUXq/LG1AOsZznbQr0vINd
TQzUs7wu6mbMhDWGS6B92wuUPzNYUJQbvQ6NxNqKK1lvGEBMfCjEYg+Qhz08C2haWXxgHLfFFQNB
Z/1buvxb5v52BZFgR77Zs4G1aNnrOjLtdSGSD1q6dIyegPFzHyDOecn8wQSr3EaeGWB396Je7Qxr
2E+0XHZDWmwz0uhCtoUngRyJD8o/csj4ZzooVxJ2qi64VsyYnq/YcsuZV6Sf7XPV4HfIdrVuIdg1
ns89mav53o7UpPxgj+7j9zpW+b+GjxaTZEmqEq8pwlRtNQxFVJvhkuphitgkCSpcLj/eujNKcV/4
0FaOLrrY3hc7k7A6JwTizbN2w0s6RcCqse4qwBgnTDbCniIDPvZ5hP6PTjsM5F7L1VJxibraP3oM
4kJArS40cBucARaTOX6nw/HV6CEquHSyj4WZlLQ4VKb4ckui8VA6q4pR9S5zLpvjOt45/yaWS4X4
KIMeMe9sqFlAhPical97WrhIFRV7AMkBjVrhkCnV+grxJOiGsOy0EAqzeVsdPkHL4d/G/Nagc2ra
3XHtWC/HS/uRLYlYBibyscG0G5NGInp0uLmKoUeC5dlTF3tlcjYgGoX9kaH74kPTvH/yZEzk83Y/
7iEXiJg6fqqr37Q+Akk6Pd6XbHGl99FuwX4US5xh1hQnMraxI6oZDOFaaBGtoAI2eP9gWeEGKkOJ
Bf31aDE+dzDAduTA93dgpC82AC2aKALrndbkGASPLCRnMaubDGmfX/MI4nJCAQYEvxLq+DQzwMxM
G89gzGLt26sll2qBTEPzK8EsOHVRPF7zGtvTG+aydQbsK48ItSOSNoOr5L6g1APPhRpV6ote9kR9
Z+lTxraZPJnzEht6WMjmaP4p2k7ixVh9ez+h6Er7xVHckNAmljucAI9Jkfp2lMO7dhSz7fkv+xLs
7exYrb2LUu0nInXAaXhx8SUwMw9U7Tj2IJlVJpuJHkARHs0dlEIYI16Ul8m7hc4Kv3RWGzD4T0yx
xy+Gw1WDOZKOnQhl0Zo7fEu+PwRORbnOXLq8PEGZRgQ+PiEFuL3OMqpZny6SEfvGB7UFzjA7elki
3O9nsZI4btVHlDyZdpFSW+oaDSIbSgyRAkb86Q2UWWYfWcxnMrbraIHt56RA6171tVUWwfgWuW5/
wKjLz2aumiqVMwsa+gW8LvVSO3jtpMepy2atMsDyQ70cVfqpH0WaJspR+Ko0D2m4OOPvj5AarKMk
mGo05JxnxSIEoFrSVW0708YPHfa/a36dH9g3i/lSTCGBrtM3k/Jm39oSKGdqlKXVttHokU7xV6rl
xG2mFIIOJjt0D7dQpEZcGZHUEwd553HDc1G0s5SDiD4NjNveMbAYCLwErbUrGyvc4yj3NYDZCnf8
axsEADtsVh6G9UoysJCMO3jnHEK8vH3tQI6m9CTUmf3NyQWa7YrsmA5X8GUqSI/4B63aRlHSzQKJ
24CzVer1XngEERNaT9k+bslknMj3/OaJKJzDydisbbDR6YosVH2TmIh9jlFoNdTZ98fiqVORyCd6
B1CH7FwdIbbfDRFxqpNw0566vJ/OPtH4d6jiFQh0FVhhxBdYcuhEiqjluCZ9NLMpJ46yKKq+5Qfq
EDcYLU2nMvW4zPjTUrJO1QVLkfoGFLMe/t886m1G4wm/MlUySALPW8CBTXftCa6FN/UTUSNi56SN
Tbfac+4oUgd76kybW9qWUKQfKp2pvXq4J7L+DTCPnkkHbCa+WDQ8B3BdFc8QF1X6hwFjEA55PdEq
K8ux7ZGU1vjfQSinA+8UeHTgr5YX2adUbSVNj/LpUltXQKC04pZ8lCqe0bbKL32Twd+MZENT3/LP
661VoqxoI+eteCMvzCqBtbczL+OzTKXVL6jBnfMgKcGXj1uTphZ/svZ1hU85I9wtVC/O8f2Fo9Xw
3K6seQvW89km+N/xWNx9ZQXS9nV0hSFFl8QP1rp1DBjV9qdHkMAPmgwjpOxlh2jF0vkYtbXYYLvX
rva1mECf9JJZ/g5dSJrLDJ0tGI80puiE1NBP+EVvDTfVnRPOMz5ZLfnPb4OFP2upIKO32eQsBsb0
nGleRp9cnGazvGrubt8BIWfxXjLmB8awrTJHIjUMrKxZbbmDh/JVaSFbtCrZ6imdmQOij78qT5nw
QEp9ap18I+Wi/zPA5tDOcrA5yiwpCZc2rOE+Q34SefRELof2ahuQbvgpmtXm7rRhGNwTOI5xFqhb
TCd7042uOPbUdZvTZ+srZgm0qdXWdPxM7hM99xlWEJveOQXRrOCL4LJvvWXpDNbsSMXdrO+ox78W
wFlCKzQdposiAeZpo9cKC0b0dfp91CPlxeCG/sACDYA4kTxkQ8G+4y5yEMgXIZHdnHx7FMqHN6BM
04YCac20c1+Tt1KxOVaCpzj1xNLks9uSLmmWYkOwvoTiTAgCnkzkWSfCa0dd4KZFZnlmtqoPtOPt
xSQOWLRcV2d9iivDQYKsPm7XeRrA38OZOq/XE8mFXKOKHRpjYhCYi2ugYfeNaA7oxrRSu+wNLxSZ
GbEC1Wf0SUo1Zy3xUY2A5M4cYosom8N/JpkPnwhcuUoNcj7AhnIBFnrTeGi85p+1HXcCLPgSxwah
dUmkEDcj9r7brLDf/7JA1y8Glrw3CpVn0lrr6btHkIp+1xLlx5mzW/fc76xTcRPJdkVvDaBGaXLz
fMBsZkIRk3UlxV38cneHzMjR7KSHx6Dy1AxG2wW4U/8AGbkrhS1t2Pps2YaPhNE1OUk8eldZHpsx
gWevyWQI5G1vFq+l2fa0P02Hp+5HwSFDPvfrQDZ/lUMrOzcZ1efZnW9YXFKSN/srogdcA3L9VXRY
JxP5f/wt+TvIxHvGH3rQ7fmJ59o6kDGk7KBDheWJXpadvohlH5nlAIlwr9sRNWMBYs2ZBYzdiQor
HxTbdwIWqK8eL4G4O1Hrgt86sNGhjd1eafWFtopxx/0lmz62S7eGTrJ8HWRdnqCRh1Q4PSuHxJmO
LKJ9MTE3hV/eDTrh2Ig3O+5+ctuewGT5p+TqqYouSm5RKD36BxSqDqY7cDB9Qy/NvTu2ovfwRizd
9ylAmi+7hjcWcIuqC+em6gdsPtWCuZLu3kdBXfcojMIYE4C5esP9o804p7TCfcZ7zmioUY9D8x5q
KyaZnkuQQJgf5mUArHj6W7PAwpCdwbE6BZUdewrMS+oEMaY96ZfOaXaUsvwtAWKkTjN1VuqWgnlD
nQj8ig8ouyi/DYktxVT2Huftx8X0TJI8wB2iaUaiAhOccfNRmFod8RY06HTpkDqk42nq9XJP09dj
54J5L5egfzxc4LZVnpKE6H+8nPirKxbrXNUF0t0i8zi2cBayyr0qT4d2PS8H3vC7KD4tqzJrdc7N
oVB4NWCnUaW2e/0jjglm15tSzW+OzehcmbYpy2A4jvKLSxOofkYistbOt6UnUq73c39ItdTzegVh
sta7VdIAonQAaFSzM5yAX7Lju6FihHYfr4FHmgo5pHJ9LDcI7n6viEtcsC80/5LaxRJ2I6ioC/hu
Jmi1rK9IXAD9z+ITfe4PPTag5milOjYRaA8PtVMr8a8dJN4/mW1FWMUlQiHAsX4pez3MuJLTkLRw
zz6VYQO8J6PnjkHzQMe0BYFRAbY2Ny3cI9KXDkoYgPwy9C72P0kdNp4mZ42DNNXaIjkz5xSkyYBR
8e7CA7DbHD63wsw+hDImWBiq3Ye0WhhOlDKnErDibIKGMJS5ynaCmR8nuINAqWUltW//zqPQKn7S
FjeNCk/wOe+c9masZCqtlOk0rXNf3Yd/xRvFAWEvRsGe5Kn6ZuznrDACQJf7LWj//nxMAd1kxuRs
UfA1R83eGIg/zxigSDeHdYTpMtRkGBf1zzF5uqrxis5GLDlUtPUYpYBIddMWSbXTL6w2Ssb6m0mO
2v2JzW0YrvkJfyw8YY7NUhnhbcdZQho7PznDPSj8Uv4zioRSMaEfU3w6IzaiaKO9VCdc3iwop/62
GFjGhqaD8jwGSbEygg5FIs1VDswGdE6STvCaSvT6ygeabW9a88OH1EJHtxxRA1BVTU8OHS5mYq/V
ygWCHW8zY9f7lImKQasMvYFK3SdvHHz+Z0XEzGjphNyvbmqNjVJmvyoz3dNbSR9zpgETdv76ONUy
Ll/DSwRU/4jW6D6Y9NwNXT6o1rD0YBtCAX/Pzv1qxhkkptHpo4IYyRdqOwpYKEXONNKolTERBWYh
JDaNeQr5UHepKVsDNIXE+vhnB5ToamAX3AN6/BTgVlZen3+7OG5sf8CI4O/KXnsQhcxnftXX1PPn
bTu8UM6sbqq9KfIKOjcOnW21QlkZAdXVRrtSryhr4Y8M97QN8tav6WowcAVg3G8lfOvtV67WluXc
079ibnNMYevVIMlvFpYCDhSKtTPOQNk98M7TmGyLVsCzXX5e6C5+FWdMB4X1z5vKfaYM3b3VE5R3
SzUpkzYa+wQTULo5EanCdvvHWe56LkImaDJdpSIr48I6u6ylBPMFqazLkC+DdnYWDIKh6eK+axip
Mrs3fYXdqyVGh6uyI7PQcNQNa16jVvSMzTFTTdlMMRNcl7IWYuHdIUTHvDpdej5uGV7h1WOHVKfn
xqIB/50C/BpQIF7NUIjHODgn1uACKHYBHf9X34C2ZpSRIvQNjxTNyfHm6JT/Fxu06BnJOiULAN7K
yXrl39FezGWZL48EKR37xfifH8vWZNAYhMoAoJDg0IRlW2na/LSUgggo/DyTvRQbZUZXr8wz7rGu
wyejbdF+V9Ne+qh3Tw15rRITeQdh5UAr/fGzIFstWG6Zf7FUoi2sdT6Zb3oSXg5hJjvJCK7NI/zG
W0fn3KR4R5ZCJx/bpyePL2CR2eHo7YkqZQQgOPCzgctW97MBeVi4s4F9mCh7wszvZ15qhr/5ePM7
Hmwy2BcTAUH2kZu8v/AkvwSyWSrjACXVJ1NxuIl9+jOol4WmxDuY5s6cYmY1xU2+NiqX7tf7EAVW
hZbvSeK8KCEFw5063xXQO2Zbcb2n2bxMLy5ZKpELX+epsf0M7z8pKRPzwEdUIDN6nfOQv7lVC/oz
EFgWE3GMF9Slv3mlEpH7pChExaDmd9Ufn+Ao2qRk9LNZxQteBcdrnGwlzOfXgK9kABGmYCRs7Wr3
3EYz+tfPxlH1hM9zDM1I0/DIz2UI1kzDZOxPNz/gxMCWm2PcFbMBUmkpZHHWlWD6QO5+UvWwfTvF
BhyWuZ2AIN1mHHdybqyG7daOL2BASY/7E4JsvDf4xk0OIrScv51EJ0+ICS8dUok3DHf4Dbtl7D7c
qTx3G4+2rPPe889O0ufL6ti9m+j3uvOz4VTFw/dSD7tTA3XExTxRXtO1A2OzdTS2YvTcLvij1GW/
NtrsKLVMHQwISPhVhD1d0MjC2YZfLhr6ckLP7AXpZXLMXis7nXVuEil2CCMDaNmnTXV0r/MdW7vT
j3ADK5oKlqWsYSqvOdMg7kWURMvDwv/2e89uDNVzws1Vw1WZ7Hhf1LPQ7NDfhaGzpxypPtz0zum3
lzs8IsthBf0YM9H5olfb3qZk4WY69Xr5aq4sda+NuRI0HvemP2RfjzzJGxhh4zjd1B8gs4Rd7KPF
86bj7z/Y6+fsA2o+3nFRaGduh3X6z9exgHUtD1Z3TBUzCfKcww1/EQ5ps0hp3m2W3ciYAjwYNiSQ
yxGRn3PAue9qXeDwuZwSS6MRI4wQg0gGAmXCvXHwCr+OG/TIQBjSbUOzFnyPRDBgcSSGV75w3G7l
lRbrkFVlffVL7OGvdNGkmEqYQpeRR/s/sAqcFi+eV9kt3OrMp0+sE0MkTgY0INn09i/RTlzU132m
yqgMI4f2IZ/wC8fYTaIyEkDafTwHETJbKU+KCeNsi7wmzRyxkV0JbbGx+v/deqvA0VeamEvIKiB0
BRhFKDqaMe10Y8j77kczMpTWcQ1oamTUjRNAuaBCf38YkJNfWrwbZ0itUFjPCnuAXSj6gTPGgKDj
5uZkVtik97Hr4zTKCRmhhcpIUtXBqQiF84ky940RBUlZGRJ0ytKN2mDrWe5+8bQyWSRRLD8QrCw/
Ccr8rnBUa/oRdCm22dVq7bMrT/IHc3m3GIxwffR/2vECmCXLQDf+cbkc40VIJojud0QBtfsoxyfp
uF4oV92xA7XAfZ0QWZisBbkE61KSCadNrWQdy1CFAGsHSFxa/o9GBIiD9Zk78K8NJrnwqIald5rN
pWdwp12kARWGEam+EAxuJisp2916AIx9lmhemEMprCCgFrzPI2b5rEPKr22rdenIAU6ggxinEI5y
kS0a3F5tpDk7NB9ZF6CBy7jgEj7uKz9YJqCNaKfU6mmfBssS6E1ZJhmFz2yfCdhVZoFYoccZEmbn
x+lNO+CXPOE6o4CMmPLvKNa3RJf+8vW0XvDz2cyULBbgsFfLeKlPvtzmkSeDEg7EvTC3FuvPGtq4
WrOoSMCA/Sx6i0K24HI7vlwdGIIcN35MPTNmMica9w3esrmNK6nYjS9mQtdY4yvhI1pNJ+ZYc3Ey
YhOMZODfdNX2Tf6NWWXoYs3aeRNyGkONvUuXCv2d1GZxIcL6C1IhDwxdaUCc1oRPicDbUbCsXBIt
58Pv4A8fJ90TRw2Rg0Z0orQf5qjFbSXEjsNA3XkaOew8DmpODCTlE7ZdXccTCZ0BFXTDY0lmHEei
UswCPQlbaZ6YHdKTUwnS6xGRCRISUFQHOi0yssf/BiF4mA3b9v9nf3+likHXeUlnzOdX8RL3dtLu
QaQ9MN3q4EFfzQ7GVFZ/6AD0oxomoQ1Vie2ui8QoXZpo5nlIT29Gkyx9tlLZai8vBgxHNIWejn9u
bPyba8fM7jPqVuom15DdjGc1GD+May7ouL7PUHEFSq7DZ9xHSZRNiJfnD654QpCQM90+Fl5H2Zh5
zGRm5upIKJj2Z2H92vBH5/ZWUwgmyHOmxi9uG3itfeezLFPNl0tc8EvNSQ33HCy0la+gA8eJ1WZf
FfbyX8mW61nqzi9ye6hAjN+3bmHcTOmxJukeDyGrCevjgMsko0U72udIXPlTBBWV9AmZJhHLllMN
2f+xkNRirrPgIVaNizQGDj1eyUUdkw/aTEeV5J90JmVIpXIiPmt6wFO17u4DJ1DxHvZ/GqAZJSrO
t7kLeJLiPrqOglMRfL3uuRz4wJsd6UOraPmsjDRmKCxfGwQ28rxeeWm67dHSeMo+m6NI9+ADMwL0
Ap+xCIpAswD/ymx+oI27fSMbH1TeI+ZgK7UFQVmY+I3dI0bEt/kXkvoLP6eYIgz6FDkhBGxm40bi
BHaUs0hS0Ol+acx62J2yXdhiHoxyK9ars4SE45yqM3tNvqbBfkj0VdC1vEuispwgrAchHR+NPSzn
+GXCVsdkyV8aQnYPpckjt3EV4hf7s6pHr2GwQ5GlY5LttSFWG2RmgKi/koJ3md3X3TjBGiNVMvIa
nrGxzOTFn1dbtcII0L092tl0203s5D49BjLex40P8i2oAev0N5anrUhhINDdwjxndtNz2rYlZ98i
ppHcKu0uTt3tSq8S9cgPBikRx4K2kkaSLL+nn3c8GvL7pn0QLfmXrsDBDC+L3aqND7WwJfwYXskA
ZdJ3LNdgK8pSKc7XFnpUqWd6UaToIImHz0ho4mK0NR5vXraWK7kBdDXZLGFIjOU/b561GUg267Od
qOO/zY2MYWtV2yzSBIn5MEET5qkRNQpd2PSGeSU0Ly6dVkMdLsws9lP5f1emCLDput1zjkaLS1pZ
y5rdPQKq1FwW1jENrbSnJBDvpXiwW6Wridk0mvrr9lhvhsAbPbo944IN8093+drymA+Z+yF3GzBY
r6b5DpX4r7+6JbPZhPCYytB+7UqCrv6ttZrE7syMZWrcyg0mFw6/zIwKNDAE0Zn9Ne8NUxVnIqdD
6z1OPFtv6dvGQ0tK0qJ70PolXc9nTH1tLzPkKv2rOe7tt7RkMn19DwDhlCb9grSusBLKo0XAXFsu
YyGJ0z6OLb7vxagArRcMvZrV5MdmxoWoQpXhif+EBlBZ5z4cqCDvM+QKMcG93zY3ZAPoc8kbCewB
NbAKiOjIe7uiU+gDiWawrzPW9C+AaciAafXGcGI5iQlltmnnCJgzHw9zG0nscmEeMKqgPWODO5QC
sarnJPBiU9z2ITTCUmGPV49pm7WxnwmEVovtwN1PvDtdm9asTDlv+ZzezwwbzkDPJVekbmHuAahw
/WmyrbCBnLFDlnifYBmDoRWA0W6D+oiUXNC3OC3m5Kdibaoe0ybg9/rTi/lCrrMuAmaXub83GoKD
RYHuWsSopu14Ps9v6z2TCUraLc5uwkKWtd3ozxXD+ZAkRPKmKKIMVgC8qotBSHnTU1khjuE1sDE+
NiFgpD04k+g/7p3KYngJt8jFfHUJaL+JCijVb9k6viPLJp9nT9txbNeZ7GZuhhnlqutiDI3wwvFI
CwGOlKfIDPYIvzcVF5KhGhNrCHX3cb+RLD1qH2K4IIjvxGHVzusk3eL54kX/oZ70/hVwlAwGazTj
RCubsLmvsACFBHcrkAPMywpT9RxJkCEdxbd6t0VomstiJD7XsIOrdi843qrxPjlXRfRtm6ERkbJ9
BNTjdBX6w0zySa/h7WonhVaU7E/WGO4hYQoh65LsP48zkdkDUE+f0r41tpom8JC4vrw025aLDIet
Zx7dKqSPQMnUxlAuMr5pc/ty4QY/PRXhc+egm80HlxUVCZJrHjlmSHWXpL02gHclYwMA2HLEuyhe
O8mmoHSJYMlYwkzB2A/hqs5FlqwXFCECYyT997jD8R+/UHlXoDjDla42+3UVepOKn0+wBt2bNfUO
rJY2V0LphJ9nSld7tXM0KaLyPDLmvbDuP7N1EXGjTCz1KrZA5uFEwt9O65MFpo9r9fbSuMqLKFse
6Wyu5ObRps/ZIRWdbc3W/ZEVIxdMOi+SksdmB5rr3vozlK5tIaDr9NcYAbWuKHeE98CtoOFH+yNM
JM+XmOccPkTPuiGObG2wDWbIswXWlBmhSpBddrIVvSUMypXEeDK/3JgqqeeYJowa81I4vLcHZWKn
VGZq2y8w7J0hCLCukiymV1MoQk5QmWALzaPmTTYUCU1FDBRiIuG0bre//uKUtyr0S28wFIbC/NZA
Qtmk6xVxCRhnj64PlEvWUXLjl5E8uhH/wb1rUa7S3vy9EixBwDz/6AGUKB82sorESPOQ6JlnFJDw
99QVjRLr7cJAVBcgGGTItGBeR+4UPB5A5Wto+Q3qpS2DAnpsocQYls/YoZb21JnTJuxDnorOvZqT
NsXbCPuYeG+gDG+Oc6BcCOQeTeJvqkLj1AUiJ2OpLx2yu6lKEu+gpEveCNI0AR5xkaES4jP8ck2i
r4XtD2aTQoF6JbnOKrWCCAolZjW5ywT6YBDqgZFrYwOO6WTWVxl7+ckTs/Y7azC+WhOMJFpFEjCf
MAMMpcmsjB19ginV24L+T44SswkVlmEleeQGaJjxPsLrj90+FVuQnkgcIfXOBapEbO+IMgtcMTPb
L01zrkFiZwWRiLhMFxOLZo7pgZBsSPxRg42258hAAk70enJGRQ35S6spHbMb+j3Kf93hAN2XzKZZ
IVta9ecYtYdCiVpPAT26wSHBOe+Eiey5ao7+DCK0Wn0RyaTkAJUDF+HKxGqDmhqtmYr4fqyfoyTa
wGUg3ku6r5NNzZi8OruV7rklzYQ0cdwS8KXMjZrTSCRVsNjLxJYPH0YbJ7rtqQaZeSk97U1swp+d
LvyiBQl3aiAHkfgwuKzW3kWeU3fhamBp4Ysec2U7y7eUgrGHp74WY/4hNSQbgxx6kNJOp+YZTT/1
TLi0LXe75pVxFVYS6hO+0rXsM0PwWki+L9rUn7/5eE8eloPk6jK/kDZpGSqU+OZVAqiKv6tZsdcQ
Y2wyu4n9xKku9QnJW7JI1cCmRb19t5Eeny7RNGhOkxIaRfPS93znQHO+gdP6grX0abZ3MaHpyrhQ
7YJFZikgSaJiCKwuckz42M5GKUkfvT9o+X4vdYQGendSWrWiOx4SiTA3WqR+zB8oZZIg4NnswQ18
rewZWjlJrfalFaZtOSEb3fwpmWqh8Yfyfwbh8wSsaC9h1/yBhk0yxJQVjJKhodv+MShhomb/bbE3
2SKhEk8offho/iV786ZSlna3HiONECgl7V4bTIQ0n5npGKH3fKauPCo4bP8AEKWunOFxhco37cMe
07mfzDa6wkCnrMb3ReWTLz4IaXXiQweBtSistGupTjcIz6UfnnB215cmNhne/1qE9hfowm4T1l7Y
9XcdEpCMZW4EVabVmKIsNfA1ZQcAQANMFiAjGFjmBMOy5d08mEI0UKMclhwYq3Xnw6bcNdooIF6c
Euk38+2oCDWvLHHvKDMBMcq53cVokMtZFiYEoUPeAKBBsWK6FROuQnQxHbIWi3OTzmK0m54oFenC
0Verk94JVynNImE2tZhrsTGPyHNWjeU/5zas48nz/y7akJaO7TxGN2x3A5fQiw9t2Z8S6fYlvc5N
rgiAWldk0iLskX/Z6a/l9hC63cRvXQW4sWS9d2hDTYjqxHoWX08Yx+yRXCi78ozT6UM7Z8ej+M0w
6lBjgkqdm+ISVtVy8x4lEUyWzYNbP4815EruLzV7obq11uaqFZx/xUbI5QaCFK0zJynJ0b9gQCtl
O8yJN8QPgT+tBjZSTrM9CXvEZrqDFjFEdqebBLvfzI2FLnsWhILxOVtMPjTjGtNVLhDOOxrZC8S5
iVAoBh01j5NAvHAn2zTUqhKEZY01YZKH2wLWUhGTFZZANbvb8xOMrL4ATUllnxg0Neu1b288CiwB
MHxW1C0fBO3t9N9eZTqQJIk4naiiHABmEfjW0DyrmEd2xyEy0asmLzV8wQl24HZLfqm98nfwm2i7
Eiin0gIEVPX/HLC5UTn5OPnQgBH/YU4Z0os7+9bYhq9snjjrbLt7dMb+ohhtAoKCbOqL8XYe0FS/
bsmyVZ+VXhWwjMYF1aeRvlCugcaK5bzicQ8xq525ty7Pi002GJoFEg/41iRlSrDF7Oz/ZcLRTGv7
/KuABylFm3gxysPWhp393qSNg4dyVNEOQnVuGpCDPiwqJYb1XMiE//cNeU/6dQHZM8clI88C1nMF
bEmqtWrGl0kxUCMdUhG7EnSIYYRyqxAZJFiQdisI6EsmGAb+oVyHVX75+jzNkieoL3945C8haLZ1
pJ26RZeV+o+JnkbEq+8kVv9EJ9JjwNPbG2asTsNomuRygRwi0uADCqwaCzoas+zJejpOxeud85ri
1Y8fo9161mhXeAMV68vcQPimb98u/M4AADZP/OBv8SY2GBhopodJdMXDunaPxKpb7ncLbGzFROq8
VFYCZx3JJvsnabhDoM40GR2CfKjJkWpVFWLs0O+U9nZ8LgeKEF6f7HuNW9FjT4db0UOapTqvSAlQ
3rOOZI2b1rJl3QW0ccDJFRBDYGjdCbiJHiOAdMkRhTNYD2DP7Fru2r67rTuW7JgLfr8lPEYezM9b
27xKKLN0wZVKQ/A2Nya6y+lA4HC2WEQV/jZgCl7qaTMugY0q2Baa4UICSvs0fG5ES40d7S6ZUQ++
RuiwZhsESrvpXTIdtEK+hkvVWJIuF7sXGuBrIBvK1c5czlbJcVos1MSESRORA8pOfIKtNidepN7R
fgsC1vbzAZeyTLZ8sTJMyOw23PNTlNasgD7S+xS/pKYMdQsplciE1/YVFzULRbhcSPLwCxz9v4wQ
x5aXm56g+2/zux9sJrhVg/OPY9PgCNU2B3zQH6082KEO2YctYtRnc/UBrwOX3Ax6q3XgZ8cwC+wF
gj+QN3FBvtTa7euXjAUxo4/AcAqqOd2680jFRYeFNdt76HtfHj3fJ/au7WDYj8Z8YY2bk1F1YyoV
f0pIxhNUwId88ppY5bATiQBWKkSdNyPfmsfYt5P8SgxoZyUQCJVPfmUYNVgiIFFQe2eVEybkZOak
KBmBeArlVJQQm8lncu8/7oyKrJiW+bnRwViLsJXzmYq6O0hSy8vDztky7TavB2yiO2rQdY51uUsl
G4PJbVYjRB8tiy8Ru8p5ftRUYRqkmMovOcijkh73dWJIxVHMJWeoK5hn4bcDJvOvkK7G/YSeFcHK
1p3uajZTl+8XsPhxiTKtKHdBWAaoM6+XeBDjUCXHKKTR99dXQRdMv8WC2Jrz2jMkMVWK8qzx3imy
Fk9EqrpNlKGTPR4awxKOP7F6ehtkKslvXl3HGG0jPI11e1Q9lLI8nJrG/Mv4dxixOzQLNalQQQ4n
XA8bm/ong9iowrKjHxXdk6SBcrmeAZTJzVP8TJQOjbEJ9xeduUp0+AEjTj+C2KhU8URzE57cab68
uNjNtem8PbUT5mvT+AsPEoMHQdK6Q4EwBKWGzzBgWSqX+YlHFrdWfOZohnYceJ/HK9jp3BIrD7WM
5v90o5iZcWcZeIDrQzDe+70I5GgxynbNSTRBqHYZRjD5WUqqDK8/4S6XjpQ2URHDPg6sFd6v8oiB
WfsnC9CCcRbHQ5zB+TeFJU7o0poP1ZzjrgxUiyhpiKh8tELdZCBiXYaqpeGUA5XXUhGXpfzQt4LJ
ISDrfa7L0ybP5eAKfPmqCblcnbUu5j3E0wG9d6gtJVTmDg8qEt+9Ica62gK75H/dxLbzYibM1T2O
pSHVqF43aMMZYKA9jr3kRkXyEAu8GPXyRWGI/PySfFd3ENU5D6q3y/uzPaBJUcNFcoOQcM2sj0MW
a3Y6eH265bXpTgtE7NxGfq1u2IXxwmpAqrMe8s04VZ4pMPcbsKq16B/8MPtj0/6CHjYesE5HoBjc
z6HHtb7dU1tt76g4OLcVJEogIo8F3P04dTG2nE34JBcKLETMdVhpWUFOY4ndqnda2XCTAJtN0rtt
oSwHweuKsmbfHfR4oRjo1DNYfabLs+ajXgPXPoYeHrRPKQi2o82IL5M6KIPFJ2AWZXLnuiR2TtMm
wUDMazzikAlM6sYQ1nTFolIlvmM0jQJa1O63q7BduyzBaltXXGLRhFb5x7B6mf9+pRWWp8R6xN+9
CMzzkCsU5Zw1rGOqeK5T7u9d5fYjCubXTltQNyGv+r/kB5VvLbLzRaG0wBeZKGXJ0u3pvEh7TRA/
+99kEKwmxYgnIw+WPOdfWQdGNNaX/Wb3y26SWbk/XBJEkRXuSSffzRkjSjcGYvJLbiNKTmBI4fDL
Rddkn4xBV5tJXfh+NPSiI8ksmEz+nNglipCRcpExDB08qgKzxWUWNYNspH5mwTmHixe+YoPOKFrG
4stGFl8NzkFKZbYWEF/13QBUTpvIDrrTFPVFofEI+rJfbfPb4bTCxPP2zygJth7jkSRgASsRJziJ
kvz097slaoBPebM+9wtc/b7AUg+RkRTTXy1G10+rpJLyELARMVqvahaLDozZB3abNzRQnKcxZQmZ
Sv3cVMwA8vMqyOGzZnaZEIjS7+Ci0/QKgtDyrPwmUr+1ZGRHO2/ypMZy2yVMKnC3jbVgGe3S32X2
HxTVc86afWhNeztWDUAiBpt/hi6xm4RrdmrPNURJkwJmBB8uyrM2s21I6R31UOKFegluM2Ba7gTn
hlzf2hBrVH/u7/IzzAd6KXnaSpcadEVBFFZxWy8cnbdQkYDlBRpE9pai0pn58oBlTBzD/KV5Km8U
Y7SSHPcromTOJGGU1ZU3qLOBCF6Ju+aT40Dr/AUiDjn0Pc720N2SvERrXbJdLXdX8E3bcnsIvB/j
bbz7eO8SfNkINSG91ohVU31kllhTNNXlP2c02OLGYy2cpqStJmgj9F35Iivy2oJiDLX++w2jIezW
agUAqYjGU1kYDxYH5FiA/8wgEZmEQOX3WrntLCq9sIgx4sl1Dys2T3UQDsQIpt1vQqQlozD24JAQ
m7qBA8vUH1Ix4cDd6ShGCMRlODWqXiQcIlbXpNUlHZGg4z77AzTC0rXGMwZ+Dn8RpDOpxDLhjtfj
vCXNNUv1/t/cxVcTW3ecgJF5mfROndBvsnQNIsfqQTAiRXcztxqfFxRxgjUIPDnsu897ltviUOAp
d+9trseVwHMbhA4WgarkD+fxT+1oxLfN2GShmkLk9PDWkIbexgXUrbzZ39oCquaHGxbsnqAr7D4r
MIyDeIecryFnEnpUnNNXv/5eUDbk0Ztd+/5MJTRgwyJbTfml6igtNKxSHOXRkjfwZeq6jWO96mbE
OhdXQz478vKV3kz+V1qo75ns22xoGrQWqYj8S6QuUUmKvUTTxb9wqD2Jn+QIDdgYJSwUtqovnUBb
C8M/4XnSOkHZu1VJtQA68AFUrSFsD8dLubQf0meZknR/fvc4FMLvp8CL8TgPf5rCWc5Otnp05veL
42ViLSRzuFTXyqFID/jB7oWpLCqboY4737D0w3X2cCUxu0BpnpNHe9XaCROyVqze5RFNbwpKrYA0
ki94Q1Ik41IxpS18NXdSQ+w8eH4QSAFTPo7gL3uMnsO3gcu56/b4IzD+GT3wUS9leF9jlDe5AzOy
Q4CQMQD/20z8Ma0NI2gfSksastm5IQJrNh/g89TzvJyDLk8K58lL2JJ5OZSduDEX+MONCUiCRaEd
rMbomO85EKA6Bx6+eqa8uivirYfvuQ1Ly/y4HRJE8XLdw5ZXDgsl8RaeY+uUTY2EKBsbqsri8Avh
SEAWmJNqZ7pBHnIeD4wTLv73X7dS7dA9DdbrWFgStim9DvRrSSh7SBl8pp4kfxt4/cMWes8+iszY
cnJvR2pEbuPWKHBvnWMLCs/R0R3eBSgqxIEeXB5vm9r0l5OJB29WwxKNBp4cBqHPqXUQn2S1ozbk
EcyXYvrtqULndSGtWmhrLQb+sSsaPSlWi22rFZYKAwi1tUqpPLJtD1NGpz8CuY4NBhWY7KLTOKvG
Fe6gwLadlMwPs6X3Yn2VbYipnLeV9AL0N+1eQe7puHxA2mJ9MeEZbhS6eUnmZE82oq+GSgzDuBpn
+4xGWCorCwa81k5c6ByG10UsWIKZNKVd7VtdL2hdpPrByXHIGWkC08+FD3HTMpiJDWrWo8ThcKO8
DctQ404ll461O6pYwz+LgcS2UbIOCXP6Lza1FZpZOs3EDuaWcS5BBrrXR/QIxKY6qp3U11kMZyyH
kwN78PrBKhrUmX52QBL9xEiFKxM57NgI0SzskWtTLgBPeYS1VOy+EipBIz7m8QKso2J0LLLugLOE
rP/PatNL8RIKvK1wJLk1MHX5eHPYLU+TO0Jp61fCd/WBLfImOly+Q4wyxrMczBgldz4adDE/hq5c
S2GMn0e0OuABhgImL9drwoZFDHf10sVJ44B5W6C1J0fzk08lVkgcNIspnSNwSIzIJ+FJwR40KB4f
+Oytle4T45f9TiP9s3pm4kdhlxPAoDj49FSAXy7K4XNxBx1KD8s+3KO5dxnmYPKHz40FXoY3fnJn
rQ7i31i8UN6IQVLUGWumpUUcAu+FBMlOA3FOWfhqQiDvbmlY7QlI9Q2ZHWw1XX43HYs1wQxACZnZ
lzkvFEOjyg14ZAFAh7FHf910h1AB/QPi/ADvDV9U9Ryfvis7XPEftWtE2SDLBGhsc1E7o8t+GhkL
2xa1aBjBKPpuEJV8IDhR288bm7k0rc+jAa+I+kvvDBqCoCZCZf0T8G1FA8yJAwezxnZZXglTjvcC
X8SVDCYdOdXnS0XYjJHT8/F5jOi2AaaSSPoWpL7k/IVUxzGcXMtuV9KBjXyFcgnoDOhslpTm7XoK
vrZrrzRQxGrGPngGoxS9HslWju6Ura0SIT5hvFiWwm0f110g9DMIEVxbRXKHKxr7ewDNClSqC4Ep
jSNAJJ0aGmdzg1AIxDuxxx+FY6RovNpxvD0S4FRzf3MHJDUHLlDS81Ffn3hW7X5h7Clz1tSN2Gue
/yrtVWQ6i30PexM5imhQ5SP+CY0Pcv23hEmMcqrlp+NWYX2r+VUK1VAOEm16zxjHkjdgkcb40Zbo
vahgu2o4T5x1RBLQIKr3oT1+Hm+28h1EsY3v6AfYtwLUFaAFXiqjb3IOj1bxFaUYPbJBDR2+6SXj
/JmcvClHubkwrzqIRiPG+S9RE2L5P1oo9uxDtyCLeVYslOpKXwH3GsSkNMsycRAu8MA2b9P31fl9
xwZgLVL9Lp4slG1wUmxl7eemFV/qlMV32i6Qrgvb7gHFUdfe1+hbpmPrF1IinzYEMeyferzSe+EG
3shNqPtHxXBX909AtUETV9e+qUtHcS8xTsFUucpqnSu4Senser+6O0p9e7B5/2pHp5qg6G/xma4n
LXU7G1Yhox4wvzJTBMhdA81qM57DMqNcbhOKBeobtHrDnmVW0AAiLZSCIkhy3Ol6mfcTYYGzbtaK
44ghtL5uWji0vog65wCbj4kyuCJISzHcKurDsErhbn/j7XHmiebMA9jaL0SWgvNIJ7wD/3IozRj5
KNrqdvojRMipULqzsJaYjJb0/z917OeXpbCoWCeSwmpB0E7cfuICbkZYICnmw1O2e9aO1gTRfr0c
HzD1qC/YkA5KXAIYfLQEpT/ysRVm13cuuH+4g0nhPaR8irsH84jlG8W0asv8jX4XS23VFO1oNsXp
7IMKxfGVI81npAcYUIOflS6OmTBvc3ZabY9XBFZomR9+xOVCcaBY1w9RIav70mAEydqTapnacXob
1A8roGNYEVE4h4sdorCEsZju5YfwOXXhKf6tJiWCude5FzTSZu7f85R4XZvyYm3wrB58OvrIMJQ0
hTwSU6Otck80j+vteVQIcuZOEfBCZGdlVng+U9Jv6aauCrE/1X8ELDPuLwF3cYUyVh9rVjMPXoXH
WT+zsxinZUqre3O27+GzVrSIivfUMXk2l9B8dv5a3LhN9hwe1A/LY+c+R7pf5DKSd0xaILROCIt7
gFt+8svaleyXHWra5MyYZ3rH9jgmMKoC3kByKJrH/+xigyuHH0RFb9tajHr06aNRIeq/rKsK/sfS
t5uf7eSljmVbaJw7pd7doQBk17/57Q+y1UGu7shi0spHiYWxJDjWlEqYV+2Zjd00fykIrKFizFdX
wQ0BdaNM1rkO0jcDQpUThWszB/pV4Z+XooQ9TLb3JvMSzUffIkNI8dw8W2NdFBc5AV2H+4LxqHPa
5cpSEL66a7NMPYkt6dRhxhIwx8NLqgOUFrC+wWqKU7iiTqV+tu8cLOlBLtoSWUOReHomEzQgQ733
8g8LAx2WD1yzxK26lnkZ0MswCVG+ZCypBv4vXHOP8A1YmU9KNd2Q88B7weI9qjvRTKXTXzVVh4yx
W5FsAfNuLBLOZHMBxE+pSeLWZ85k6M02KTTi7tBNleK6ew1AYhUYyicM2p44mkYB7gmdwGh7EwFJ
1zJD/2+g+Ul7T+Blk4QiDfvJojZ8to9ge5g6nqwS36KKSAiCBV6ETytd4kcBYVvgUTZ4Win/j+rP
ZXiu2KS7kYJTBjD9J3wX5j+coKZvI6B8cFRD9yRahRm0gMNFtNIlQTWjaQkKEfsC5Mu3G6+5tQTg
PZUHRXnKic09ODXnwzDZI2yLNxB8JnYOeOCW9l6uDYgl1kVjtWUGThMETj5tUde/TwhwB6iHgW1m
ifqC4EcgFprc7wWIaeozZFv6SvUZMxsUKZ+Y3qkhPy1bhdiyJF0zQnAIWkaf8YZKB4DkF6ihIqON
HeO2RHBxy2r+mOQkXF7inSS+tzNbSuFj0FgaK7DMCOq5JU/OknO9DZZ5vjcdXOUYnxMXpr5+JhsE
CsRRuLNnYHk2m1gSdhGNM5bAW0Iq8cY93Vb3+KUGanyxQXTJg75zZr/HwFJBvetQHVUMW3ykWr+H
kPn6q0hQQenRXpZ8oDiRadfM8U0Na6Gtve1oIk3HOKSUwI2j0mK347SBD7LAgn8YvAMQn0gs4Pk/
dqoYAZi3+Bop0wuUJYBpAoX0QJ1K0nEkYNq1MprkSdnsi8f0Z2EFYH7Bj3zLMIyI04tBHK6SMXFY
haSZpSprxhAPfiYQ3wL/BVJxUoXMteKDtnp/cEmnCgQ2tSbZubvR21gSsGzPB1DQ2ZTPDd2Wp1VX
VNMo6EIEw5FELQ3/Mdxn5d9uHQGQed4xAcvIX2vtXb2JedjYvn5goGNGaGpPnQ13vMWL2Rfs7Axv
P224zmhRF+9jGIcev12zjozJv4Wvce1NFeHJ5t8M9/cuW7sFhVe/E/jqF+NpJAHXU5dtUS1gSBkG
5yydKibw7kwt6INfCs2LPKqV6Wx1MHmRLdkMoMBar8yhsP8EkPHKiajO07uUyz5tpCAOW2YthQvm
tNnTzqhoUeFQfDx2I5Cjwfp8Z7xSjEfxfijQDaK8uOzj4592A4husVQ2UhR8hxC4o20q+NDlYyqI
T03x0TCT0gsE5ff8MryNZ+GijOEJG9vT4cxi4/UTOWAUN03tqG8cfnTjZ3c2ReS3ce7vALSxLYtn
Y2XltYW35+Eqo+QmBJbVL+qDLkRlVCvtv2HktOaNx+0VmkOO8YgUOV6a6YLI2sqoDV1TxqagAND7
WZIP4wED0Sb1yRzp2nrsaHBu9RJ/HqtU4y61UzMfKfrbQaT1ajQPzwX5qYXrq48BFNlP9Yms7qqs
eByFwC07OM0Dmrixa73JByFjXvPruu0Q2aykIDpmYIZYAFd7YLX8VcEi7kG0ESeUi/xaHpZU3NpL
RNRs6lGax1ic4m38cIJJMQhbasErwjJQYNpI/7UHOBAV3XgDk0fv5S9KViYEyYIX7nQebokiCYVO
nPCnwwBA8JKeFPJOiF+X5XIN6FEL4gzKjW+HZty7FZVvKqiPBNVyJq+SUZcTY5kJOwMey1fdG6lb
vAa7uoBdb/8Y0OEUFg/j3WTX5xZ3DWZvd8g3NUHS4b9i0uJ9C6FHrLtzfVR+ajpwKu2d6zltkOoS
lYUCSmAIZrbshbXffmcCPhlCR5N/TLXgOIkl78Y1W4RNLol1ptgtj5LeDfneHfmteHkeEC4BNgps
V5TkRoEvwAD9UF+nOS02LPDwDkvxQRhGT4aiE3V38av8SsRKggtZIFGeV03xUWIiK/Mtt7GNL65l
NXEVAt89dnldEmGkTT/G//7wCI5JCVEpIUqBvICph/dvd4MrEXCuCx2jgFxeSUV6A5QVCnEZrUXL
Uzat9e8n5H8Q4GcI2W5L8G68oqX3kzl9pjqbGKe5sZju2njWt0balPqMHKhYZBQ6LoOCwPTyC6hr
Keffkjawe2Yy/382JherRvWX+QW3qA4dp9R5HUD16vfKKLx66qd+p0WjyQUPCKHrd5xEZvq2XN4c
lDEEMM2Y3ziJ8lw0UmlXNN6d4zeKFL47VWCHsj3rMTlROSFry3J+A20c2/xdm96+WG9unbnrslFB
HZT6XTFXnrTy4muIReJeN3MBrGBwWxtXumPjmsDjHZ/fnT5mPkvtTftMXBS7gCo+B2hiGB/a7DrJ
irqZMdXx267y30rS35a3YsckGHjCen3Tpmu/zYKDsl/Sr1kmMh6YZEWecYlB0q4JQoSEvvjULd62
ZmBUdOnPlMykdhwGLQ9PcIP2qkDDD5YhwuQvVqurKPc+j5+eqhsnegIjUWTblmTDQt766jvZICUa
BDoPbYY6q4c+pk+6IOMC83yWHCTXkzJe3AUtu4O5rG7DJ8EnrvGWvYFKyvThNw4p7SnBn9YC23li
e5eNUECjri0N2UHge5Sd+9ZlxaSZUdPFyIBHqlv6WBqG5YsrFlyr8lGDtN/0henXQIEy4mgwUVfT
H3owLdi83KQycQLiJWfDK0kHNcAheHfsIpD7X/Gd4pa4AXw/iPGhfVX8d0i3oLguQuB1OulcifpG
Pajcknx8DqmdJ3owExtrkeT76y6bcogbV7o59D2fpDGLrEDsPc8KSUb4WhtFYsHsTWPpDP7c+A8s
3uTkRqmY0t22bxSONKfITUkVJSxzAJWoJWCF3u6E2MrAwKP4UcGLkWyC4KIJRGB4F5YGbxzDTWNX
jjDm5LBtVN1j7Jjuqc5OtisgihWwFlDxhZtZt6fxfjFHd/bodrbPrxIwXAepklmEdb7HXix/gk3p
jyyFtwMrFCuuca5ZqS388aN35i9rgFYmhHbPxV2uJXjxM1fICpY1OSoH6kAqxeCn6y8Rq20+r0AI
OqvjCndDYMxp8AZCllnJrtd2GFdtDz62oDPH7s2TtLfxLY/g768pwcLV//KPzoj3Q4kTvCbtnh7z
uXqaAauDIZ5RIcAzc0UocxJ23xRV6PrNytzT0x4RLH7JSv+hes+pTNp6+bI85fHBc49mKP4GUsS3
K2BqMEfHFtNIcupUA0+3/p6+zoRp9cl2PmVmsIJZ9ngjyjGfrqKRyyIlInZnKNbmQHSx6TWBxAXj
3UkGpIt6tj1C9BSiuAp+RiUvQonG3opQuIHgzemCyb+w1/yuzFTYJ1Sd9eS9Sr6EbWO2R2Hiv2vF
1uN7UEc3CVHshOWpeyjXqKiRB0Pwm2/wgAxkDmTszk1Adkwjrp2LUZac6cKCe/0BYA4Uvszhs6+c
B/Oj5xTtJ2Np7R3xMxHzBgIuIebLPGqvM0z6EElk8jOAjcG3cWT27XAPX4DdrBJeclezEAVOKIfb
cdcmvY7245z2YeXx8Iro7mfWEZ2kXq6mX10a2J+mDPMS1IxJou99MwwR/ppl6P+RqRO05RmCK9+Z
hITrZ6EeJn4H4k/hn5mPvwowVbcCxXzG8sS/zV/sQ9TdhGXotEWhXN8HFveFDonOci7ASeSlSiok
RqgJ/rBzj42F+gZOFSMwMiPfxH3Ep7GbZV9R/C3JhjOMNIZ7E6h3UxRAjRPmnr6t9fTEn2sLrc0B
JYxoQ3XN30HxFvzQCwy/IpHlXSVB8qyITP9S/nc0ojYlvr+KOdmwVAPla+EK6pdWT0LY1lw6x5TF
9bPlw8oQgLek+Zn5KmZwSeZR631FXEXAI8uyU36vWodTR/Ypmfb1aToNwtcxIbAVV3iBUojIh0Bc
yDKEqmX8Tbn3XH3xxgdYR28DSHskrzeDt5pWqQYDc9VkJhfWI9Jo79Y948kSxS7GsLYoFF9zjBIb
3dOUcEX+c8ey4OeRRVZQOHxskEx5l8bE+Mdl4hi6qocgO15h3ULeONq9JFY/UjpK1HHzJWtwdco8
+9u/aIhBWKNj38JIPBoh6oQ7d+zG/i4fS+vwG8Jb864vZe7+ShYgb9YX25PzqE13NPjgJqKbMvv3
Nje0U75hbO3dwBoYjjRyixlYGqbH8pXg798L9rOpicaayEOs43dVXXkDpo7KwkqCLmyBsW/Fg2je
gPU/RZZPDovyP/GYYb+1Fu1JW0BxBbVqbrvzRUPhPz/ih6o0wjN7GvmHpDieWjsQL3CmYdWdz2eL
uEQqyGyn601d7YZEemUC9T2MzcywpvHX7I9qykUx6E51fwtZXIIic4f5ApF0vpYrlrBtfxkvkmWv
yaZRyVcTEo7UcOM0+YJQePMews91oD7CwdKzEGlvOrH/Ub+uu5Ufl5nZvMBqLkPHef4/EkC7eef6
xV6Np0TzKfxqZ8Z2RX2ht5djx1ynMLqID1rj3XgvM7BJPOpqNz4Mn8L21BPeAr0zxi6ro+o63vSb
nmjoQeakCu8+HBiXkrGpHfH9NP4IE6w6KNt0CQS1mRctdU7zdyoZfF3IGR9K/9x5XDqxQqDhECZE
/Wyli7G7Vmkvq1XLBJyxbCvc87FbjTNZOGz+K3iybUpQBR5UnNdZqxH52E8jGL0CatnDl1pip1Lf
05Lu5reBxqAeCxKxLsUUfHgGBCWorRoDEhkWB79rORtWbc4uAnwQJXPNb1joXqmMGoch1py7ZQ6J
Wyl9WFAC+99CvhCPrw8T/8AGGKocH9XMbB349ODOD9Od8uEkKQo1lrIFy9AipjT8uLD6zIIyT5L7
RyiMZ/eE1ququzZzQ6p0sK4IMVj8ikiBN6IklmX0MTg2H62ZLqhAn7BEgFnEWtEpNniMEhHDDD6Y
I16Bl33QmGoK4sEJIRv2n+1nXlf6uDOaCubchmBeiAyNLTXF3yRJvbllmY19ihyf4JbiNP9OgJxS
3Ph98MvrJmWI3a3w3CJzT4TzBbDFMws2VAOqxSx9O7/8y1sw0JIo16vnmHRovjOEn2aVYL/T+vt7
lqWc9uhfgeo/Wsopf1bD9L2O/WTIx6EwhRe/r/+3Y9vu5aYb6JV4ry+li6vD0rObFoF2ALostwYB
g+p9sYgxBAm7MSVe5crG2rjn0RkzDQy6kp6YsjK9B0bCbByAqk/sMR9wz9U1mAzwsotVWIsjN/eX
9OU8KZYcuQqW3MhZ4XAPCqhaPijtyb0BXBdbZmhi3gCLUsHnHUR/dW5KCpqorAvn/tBb1vG7oSLA
wovf4knd0HbEWyyrT2UsldNzy31pVgqAU7tIS4Qkd1uQSSYhF0xvpccQuDzoDZcMxZjK4DySyOYB
mtlAJLmu2TH5Sz9nrxuuSRfpKXmcx/Gf3sXUE0ynI6ZxrTBVG2OXig/RPu+KDv4Iy9apel+e5ie5
6fMyDp95yZrWz3REU4ecmqMz2QtruSIy/JDrkVKRqzZyN8fKPmEjGdBQVo9/UGIP4FxsIKq7wmDF
cxaPxdibOdaWzrGt5z5SdZSr6hd24JldYlyrne2qv8EQF/EZEuFuYUa9KuZdR1WcJXPsJW75HHK7
+vwQ/NJ3151KJJ9IXb+VTpZ9arO4VygiDr+khKdJMM7wcUJqeciIruIPneUNCSZsdSuGQXqPLheH
6nM1gGuGYy2O7cFX6sI50xKRuKmtriS0z+Q9Ykom7c0x4YIysyKtnj55XChWVa/4U1ZHjFgahJvO
7rs3QTKvBVB+K2fSQP8LJpVfp5UsA13+iFs29Dh76esu6+gh/MuTDBL6PNji2ZXccZzD+xH25Tlu
649aopqzHES9AcRrDoqHLBqvOcGARlwwlv24FTW388qqZlP7hMi09tQlI6TQvO1SW2rOqGSvTx94
KWusymHPwZ+Iibn0J4UmYjJLPS0MXRi+1F6ZfrqpJgg4eXlmrGpmC7HKgErqbqVQ2vrbJEadVdy+
EsnwezIg0iaJSUL/JXENwvraHtTUegRqGEdahnpnfyk3mTknyt7IYK4gxxOAYC6fna0etTOEpyyq
G4eGrjSTMfProSCqXiy59iWeAOsSO4SiKH/iiaPSzXSd1D30OWEI4ADReTiWBCPuerHpq5SpFLDF
vKWcCW96zRhXeLB+b6Bskmyvba6fWKgDoUvwvxND7i4BiFp4oIrDCwxePBesXaFLAppTuJ8DlMe7
uQyuwtqJdjVYi3lswwl4OOoYyCA/RGUfC6bTeazDVlx1TD9pgykGr8Y3pmx2OyVJbvEReBa6+6zw
cSqi9i/X26hdVv451E4vBE5TGYFSEvF4NlHJJRsk6aQZ/EQwxqcxZhWTo1xa4/W41nD7gd6PXGKt
uvI0Uf0goO6gJXSmQ0i+ItexL5FzYn9gi/bj1WpAaJp2LWMl1g5fNS94eiiZciw4vI+8I/Bb+VY4
tgZyI+99XQyLu1gdpA+r2q148qetMlPPRhvbMMNhc66KYSAQ6bqrSXn04dYgaaW2jWdQyPXC+8dK
YqWvOBSg5YTSXoZ+AT3w8Dq1pq8fBzfFuqNLXYrUqbp64Z5V1oynCUZU01JK5l+GmtiAqIQKCCHh
3ql4bCQ5LefBsCUIhNTCWEIgCmKr26sko7kPaXOyl12Rh4FiFkdMSuQEiRVx/YZfaBuEDw3G2Aq5
bTCDWam2H2K2r6UJvvfppctP6CprWeILyWzcKAPytNp3JRSFoGJWmqIgKsekO5/UiKKFcayqSOSe
C+2xL9+ImbAhsjXwvj4B/zoEwMfOXxQH3PFg+WpsV1HoHFBM0JXZj80kQLvbJrpkTZY4hZJJDrJQ
rO1SkNxGy9pU/pDTh3vnLZUnnDUIXStK96IRyktvciwFWOpYvGdlWoBMRwsxzQh3n8jR1db+tSiD
clYJTGPPhZq8JscRxm/HWcuvJ4lLZkQmidpZ7WOJp5IulKLDIOiVgxL3mLPhalnH3ds3SREujmxR
gEfvl5MzftSeTUwW5ZmwK+k8PVmU5GEz54PyKYhtutJGSjWkka4BV3ix6bd7tykyakCpAG+wc5jY
DLHyy7pRjd1mqt3tYA7HzgL4EU5Iiiq/v2TuZYqvr/IjRgZ2HxIloQy/P5Bxa0FR8Yd6lZz9rUTW
wQFugWLrSXNG1HmIl2P0VOrtrJ3aHzgtZ2zkpDiSVDrR429f7mKdjjXgtAtfaZirwMublMR8Txs/
9KefuFutywed+805F7HnVvxbNB5UTB6mkGfx/fX9Z190zhKFPtz0wF3r8QyScaTbgSesN7aEEjs/
O/qxudk+BUCYo34affc70tA4SddHLDhaA1G9DaFfCF8grZJEq75CEFTR2wUO3jycCjrijms8RZY6
cALhH7BxA0YVSqp9OzUqkJLZh23IlnNuWT2PsYOMlfEySoluKm3zh6Oz+4duV3+eM+y1Gxw4599I
g3vjnHChM5tx0fqO1057HEX4FVheNd9V8HtD2KBKg9YztJ2+AU7fBpdytID+8I6bl1K0gvgLemlA
wdaTqw0RnJZOGUOAPFTSyZVRvu8khIovrSFUxEDCNSg2aep73Th/18wbxs6SCTFa2inmBohmq9QS
K4kDS8jTxE45JKyDTWtU+ezPP5fuf5r6hI0uoIaX0dssbRnHsbkuKMhSwscSwd+YGw1WlNkTi3Bq
ITpn9kyfm/wkzccbhnIDmEP1MepW+lUHzCsiRVDqR3uGJ1kmofxHlh/Pss+99W7x7+EUF+IUPgrL
Yrr1/oh7pOkMyKFiMmTiAHldRPn1tEnfpCstdrH4cJk1PkxxiB+sJOlnAtXz7gjOs6AMrFRAT0BJ
ER856WLHWEuCKage/8m5DgXH9xjfkIG1WeNNFuz/tp6mUx4w2lZ+rvRTKb4aUR3RGWFJRxXB2yzx
CKMtux7MnS1lN4loNSTGe09RFC6qMrgyLankS20RhUgyJRSi9XdKVRt43GFeE3RuRx/2/zUYMH9g
4CAFCKdEBi/8tICcEmGEJrQ8dZ9LNl6/zk/u3o5PR9/hzH8et8K9Nx4a0cL8RVc3I5IiDLzaDlu/
z6oP2b2UK+C6xSXdA1dFACMZr/BUQF+oSwPmSE4MH6sBhCvzJfTQvjPb8n8oDw34VRpqzsP9QbM8
bfJzrY++QqiSg3m7q+N8dTVVwPApsdbPKmsjbWdmT+hU1MRsFiFpVWqsEpzQIYK++++GUNqCgYOn
OGqj2/swqGtSOLemgwh0FlUzXhKSW/lzAvGV5mER4zcZs3OxfXPHc4H5gPBSAbEi3QEUNWGNOmlJ
oY/vpaL4340OOF061xHndW/pYv5jK6UN+XmPHsfMccvIiWISdTrr+PxKHRAe/Hkc/lr3cFIjNhTG
bblsPp4dcv3tBUDDwZhp9ZehB7t9xSrd4TbKr48XYkzPfMNlCpElEqcXw0P1CspW2xeZtPKcSB/p
UH/9gsd/4e5vhKQBUFHcVeNb+0u7fnXRnmcXwpcmD5yhzDM2P6OudsBmQQWV/9LRFaFqJbyD8YUA
Fwn7b//wnkq7VnYYCp2wb8zdbRVzX+dPYdZyASTGik1HAInCtkaVce/Pi9xuxkRp5kYDdBATialK
WnsNB5to3EiwyloeTX1CyZKTSAwYL8PNwnWbZ1uEciFg/q+0Frtzn0fhYM9r9HBqk8X9NufCBLbm
8ggTHRyqwJz63CPfzLFjQhNKk7gA+2KSR2hZ+1z/+FvxyS2EAiTQfpeSoB4jCMvp/ouCv9Dn1OU4
QOMFrZU1DoynJLYQMg9NqhBNdl7MB46UcgC/OmLKXUQvNYBdKgzAm6jARnbZXigQYJq3lpLwfpaY
c7ky6oIeY74VWAh25Wy05inRoH0VoP06JwkzFWtk/AzmsdYzS1MOb0EEMtEvhnexBdLww4Cvjk5+
wc3cTG3Fj6DO2/NICVXO4nOPtcFIq/87jDoHwnfog2UfxHCyLVSmg0gB5h2jPHUy2DZQv6SPdlJz
HgYkHM44Q91y9xcg02Fbd7cWJnEVJUqvobZUYXIFfBexORKRaaQ56EnqObmaW8cvL0scvjjqzn0l
mTPnqWCvqlzp32KgF18sPoDvLxOQP/pBMRPnYX32l6vBxgUfiBQeTx7jlQuPVsAANbYA7FBwG9L0
mgNCnQiMypEHt3KY3XL+hvNxPz8MzbIsOETF5JwJsO+WEWrnr/eAiz6lDNgVkX3phOMKuVzc4wfg
dCIVs26Zp5FZNPLTQjgs3NLZbg/txNirwfxMJb+6IHlB/EVHfARUWOY24//gO5S1LJhyqwxnrAMi
4cMoVGmUKqxPlMUBSRlS571xfm8uNOQn+HZ3E//5N7F3fDzRS8OBhDJ/weI/S+R7wdeodsqT1wOy
Bxzbzi6VpIZSTtHyndubsKJb1j8uDZXentLWT9P9PCoETj3xuZNZ/KRBva1hj05CrXKjG7ea7xu1
atCWVqOcHUXNwl8MMAmCWs8GQe9GHbAvfqdNmIv1Jeui77m1Bibtd30pr/CGORpqo6I588tm5AmU
yLi6DunxJQuH1Xankux6w75p9gfvfSXH2/1ues0/MozfzR1JdWPJEkKLWCYJy+TdsARCtuWwwp7J
SuEnv3y1gPmD8phhXbxm6XazljuvEO8aMgEZmdk9GTvcQdTc5TGpSEXPhptguRLbjkd4FzGpYtbE
X7kpIro0v9fSaEkxUZnwg0o4bjGxv234NZTtHtw5qhZeE1cbyZuB5JOwQOf5E38G67R/Eg5f3/VN
BPlbV+3SggVJRzJRffHu/5ZuMMDwELP5N3oVXPNQwwc5qG9rHJ/O/dAYD9n8IXGe74pgazU+X5rE
dqX6Jo3q8LaEpcU9jWE8Zae4cKaH6T/dXIS2kzNG8rNhhw0FxnhpIclNiHfoPrwr1WXk4Zf46+sj
SRpRzkl42oRM9XKMKaKkHmL6LsgQdZWPiWKWdYjFl6OT6UQIoG2zMa7v4cl3RCgAgiUYlB+x1znI
yVDSAkhAa1CxTfpD0t+2N0ryRn015Ig6JRY310y2kcXa9sLIvefXZJgHnFZYljEVfCXw/HFnobJT
VvXiHFW0kar/6FHn//h1vOpr34dudxzH+VLBXOO/sJ0H5SWb+4czF43TOKARpBN2pNW+Fm5JzSMa
S/5S/4t/y9sRBpZDjtS85KC6tqswtgyj1Y5VCMQfX/7TxLzmYJCBPmzz0T+ODbT1Ifz98h3uWmRv
MK8S1457dQx259Y0p1ZrgIQFsrmwVbVj9ZvjrKCbs1BXo0tbvR7SdVSZMKEKlw4yMhvLyRA8JwrR
t1pV+1KJPTKMHkahxPvKmPT4714cMW5/i6jZdbpkLqqxxKLwrVG7bLUXaVV1azwM57WmVd3t9uxw
pD1YdksY5Sd/sElqF8z4VuSCK4aOv7HGCUrayhTr7VcpBgHKQg0ORQxbpKan8nsqr50nj0bL6fHD
+1hUjC50TiOue/iZJ4sWPRy66IYE5JH79leSr6jMXyn7Ooss1YRVihQ5+2fmiYuEQ1C2xZvjg/+5
JeJegIc3N0dBMILrtNad7YyzwZkQ597/X3VamQyBSzzjuyftLjrUXPZc/o45s0Uja3IjWfBK+gN/
+N14M5VuUZj2YIGpZwA8+npgl3RX1rY3wAk06xT2kWt7s0JKXxODNnTX41jsa01aVdmnlP17mZh6
mIaqhOqCxjEbePEF2AV5m5FFsgnqj96XbbAI9ZFSbjLIqXeHj21kLFB16EOktCpYyf9Yq4Wa4+H7
2pClJ3O86hVQ/NIPRcp0vmwOI2++xg6q+V6L1strPArkvjUBZVo/aJJKc24y2eCIfU7AbPZ7Odtg
3hAfyyIond4eloAQy/lt7nuCV7ARqC1+NeLYuC9A4fiHGX4MiDFJI0RvIs9zmhTxNlXv04px6Uwc
wXCoXJbUqNG5EY7K8Yf61EuMWNQzipIlVKFZJermWJud0aCuSGjYAzSBD6TCjl70fBcKKY3Ytgoq
GKaRzGO+DJLYC2TJWaRaco64Rlhs29SSVJAiqKqz4X4U0+Nf8MCU/gwTzMj+qJuZW9ZNBH9K9lNW
/sMXemrN5Hb0Pa2IDWF3eKsmf57PtdNgTgc6QRzWDtmWd2TCtQNNlsg6whdHA5pXWZkhO17CCxQQ
7e8/BRN4dIDB6nsGOrrAW5IwtXYxQVJHNYb8JIirKU7JG+FBvl7W1OVxB/KIaE/v0FeHszUAJBSz
PnvNPgi1XJNY9qX/Vy1t5aj1cGl5Hj8DmADoaRELhy3uP8gHnN1spw2kzy4mqeQC6s72ZWo2d4dS
0jkOz6yvm8DKCrHjdj1j877KbQv09B+O1kftafXzj374Jh2XcEbUK/MSjYIYymd0FmoQ0VeTPfz2
LET3k6qHtZPn+BRX0r6JwtZhtjQeVHGXlEPmaF5L48LhvFp/QHIT5vwsnO1cg0SG6NjcuClrKcUZ
Q8SPj419bFFWpjvdEwKW+UJPk1NnJuYr8og8jgGYHHvhIgpEITpNM/gRGGUNGB8HnRg0b/mEG1SY
ya10zsIsIkQaxBoOPXIpd2RWyBYtvTvI7JxJD5aDLk91GGe5nLKfVRqrGLqIW23oYkR6GzIpxVKw
tEsmcL3qk+ZMqZn5rHsp7exxZOhpImU3eWyT7inl03IdU0UUiyIRjzTFIWK2qLreYXy9P4hw//ZX
5XlKuU6Dxe8rrquVl/+wFdJ71cjujfxepYHDloY5CCTSDHbYUwRKdzf+IqvAZRvQqj3mlESkmBOA
s2HGTWGr5tkwED7EmPOQ1cqc7bW+8+oS8xPYnQ9IrYPXyVrUSa2vJjO7Ck8gWA8cxwz16LlZzsu6
0/FGSRZOR1FP6iVFST0OTHu7zs00b2pVwm7bgh6f/9mTX7KZopi72Jg0BVvNjJ9OtgdbDTjPHubW
2hyhZs2COuupmeNLs4Ns4A5tu0bL16OFW44DhQld4IE4K4jtg7w+3pjh7Q9bK46h7V4qOeZt/0Jw
WUZcKtHJhGnctVxbTKm6uHwVb5/QNJtCppJZtfyts5TosuoUZI82+Az1hTm5mQbdhpIRynXyZwpy
NPKgXF/sgUJ3vWjgplk0o/KMkcnTovsPm4Mc9Q/filQHhYkJmjQstDUaFTTBYSSvdKNMVe6O5ePj
yGrBE/icrfPLa2BSprRjVDHQjYqstWsFQ+DTPL62tiYG94Ky+vs8hh+34cL3RNO1+qthNbWin+sR
fWBrKPqzR/aYBwuZLbQIfdDWzws3wruuVvsGp1wXN1eukdpjc3L2ULg941BIA2i6exYvSHqtniQ+
G9p7UQxBnFlmEKQpWGMh8gnUMqs6f228I12ME9sfwCoGri1f5IAYye+8JN38aW8DIqoXFh41eEUC
gi2htsYI2MwlwXzpl6NIk7+OemleVOHCIMkoVv1KtTeMpVxGsPobLKo4KIWUzX9SqzW0IAlj5lXD
wmCyQVPMXEfXrujTHN2Sizpj8qOaf5LZcRgjnWX9YyjmohKD487j9jcYvCXDE1fbzYDm2mvJYM+m
AIVnixOG9XSmezuGpVm3YnJA3o9XA6wpClZZlj0UhFLEIYhTLwn1I/lcttkiJRNFWwspOgS3o3FT
zQrjRotk6auk43l9GNs6vQuDCYQzUwNlmHY+OAflF+6HVIj5j2BGFkXaPI8oSH0m/dQFdRYSm9Ho
vVTbIkaZW+VjPmODOLY7A8Ci4Dzu6dWvWLRbmDNz8kVbQNu0eDHw6aQUnjLSzwBWE+dB/aE8kGc2
i0L8EFSQm/gNN0aPOlBoYKS1FOx41oZShSMdzedrwtjmXACgtfOCrApZVHASN658WV0hC5SEtQhB
m7xCnIbVuWJ0Aqp+DYw8eLC05AL9QzwR9FuAYGH5F+INe0NL+BnHITH5ZR+oVJV9A1cOsd9YxnSx
PdmznUpZ7tcAiIa89TYn+4DzA/VEuZa3UrOPaEp7UNcskND+GbI/XonhEHI1y8SNBz1CDPUBhthD
69gVZvWsdK6Up95F+lIswhmTpo1cpmV4v5djCWwO/AwusKVj8d7yH2X4RuS2j8FR6MXXDhnaDJxd
q0fBG246s5KVWsq/juPZXTne0CIZQWa43+Rsy6qqXeGK9lAqkqTrBIj8djQxmFWaZ2dqLMgbki37
/F2bAm8tJkjgqj5GzpuUGUouxT05qAmZkXm5jBlSpYtySe45Qkl8sPGl7gucYroFdNSqqQbu46n8
d3QtJme5rktLPtwx44+HQK8ascrPEACG/fk5x9Cl8JrjjGsKMKvn04ys3Sc2MwuxXCx0/SA4xpcF
sAyTKS/7evAUXXPoDS2/G91Uf1G97HIe3Fh60Fh0RhZc2JKrFhh7RjvKiTIosIpCHwfZ1R99qKcx
NpANraDeMZhogsIyjVZojK6vnVfAUk/oh709160o+1CWNqrjSuTllTmmwhHClw1Ty7DjuURzVuAb
N6kSy/5Al8mxVeEpETuScaODHgAezsmceCIK+oVmi3JGFLWQG3tX53bf8R1gzivr7LYF7muk8qLx
FQZE/PpqHcnuy2nXeAxzCcAaX1uzMcg/GP+d5G4DszBj8KSWfEtQ/taL6YPyMHPGHme7vJSFaxm0
F2awM+EuYEMjwE69k4jfV6v/a5yZpm//S1sPpYdXFIUYYF1anQvoPAfZhj4LPpPuhfAX5GciMHjz
tubPzvQkOn504woHW8GL192xPjLNYn1c+8RuhSFD9I/92esQI/FxJATX4XynexFUJmuL29pru0Vg
qs2hna2lfzVeYqTmxSMGQsv7rSCjVJOvhlMSC+2YgMlzsaLr970tVQAWPgFEjuW4g3BoQ0wQrezc
qr18IhuUosVAdw1tXAsN2dBWnGM/qfHBnybp0mL+K6eMd3AS6U7w4aWko2e2Ro+MI2Lx6JXAk1OD
ZIrOnxPJnruJPMC57hv253RDevzig+w0dsbhGO/wSyGjcoFQcd1yFwnCMDkixm4VwOVy7GtnFafv
Ma+qJSDFSnZNwDlU2hbTXWBc7PCN3hc5fLknd+yhCrvfSrRWiE8wWz5XjkToiCLo5FzG3/dNbwY9
DQSxulKXJyS+7A+llUM0RGjAw9qNNfPvmqukCyzzEfL3MqeaHPY/sKeFZ1oD2ZRWxsVQW5VdAfDC
COQ0l56oqiGdvL/WkjY2SGqHmBRTgz7nXKzeNeUMxKjoXZNSK3MFhpvho8xuv2U7U7N/ls0z+avM
vX8wgQkR8/PoHBeg5tT/v/WOHy4bq2GVofQX1kHonceTDQIbpZfN9WrW61loQfy3MXvgJzDua+id
oQYqUaKy/ssdB12IT5jshBl598aBe9gzyNHYmIHW7+nwsq3JxW6mW54giRcV4CLq0UMe5DkGsRXl
hOVcF1OrMPv6mba2TohevVsngpVrbnTDGvYWYhBx1TvVO7g/BlDSWq1ne6lFVYcTNyS1t9E3fPow
j58jtUZF5KI6wkSMZrg2DDILIuvAJ9fKXc7VQg4ascg1y3ABSRJlhSLesoVwn5sfucEfJSQKvhjH
k9WfSU0KkFZVE/epPhBMXXjEbLq+k5Y2OvdasKZmm525oznUp662TrHPqjcGhB0V/DKBHfa907IH
MB0I2U1W3qh6SyXWYdFE7em4lYaSCWuaENXbzrlM8H4Sw5ahRVQ90yGICZ5GHwU1Yfp8SDKb3urE
gMyt2GRz5YDrgLud7pkU2ebhzkPNx36W1BQuriPW4pl1SbXRstfNN+3dcVA2vC46n6gqB7rn9Xcr
CAgKECHK0kwFhleBEAQ0CiNJH3No+dqWrn20rk1Z/44oHEZ1kg2qL2uhc92h5zkxQKTlT7HLrp6x
Mta/stoPNBzr3QGzEMGjYzjns2otgQnjfFDb4m24ypgRgkgLJuVUuOe4VptVhsd1whT/JrBjkV4Y
1YgOLIkDex8W0uNIIg+weR3PdoI5vr1tJ022w89sNwrJuwENmrcjEbzoseFJVWk7AVplMs/fiT5D
wjpZJ3PZR9bKjHqjkNkxNbLCjndiaTjn6xvB2uKMfGTbDYY83qTg3B8Rwat5v905TnROJPuC4+fb
/Nzdl0+jFnyBZd7K4x/bR/taIgXIR9O+gbMWF/yHSALLvfU1lwhuLJZhApoF3/RZzwnPmvHqOU+Y
OqnJ8ivJqam7wPYDB3xrVKUTjQ+MPhU9hKdyFcIZ5ps2++DDDqmpUKNIEIq1gIhi34UqeUo15ygj
S4uw1kD/Qjogtg2/YU0N77vSLUCzImKeFcdeyj+O/acP/ZHrUK5dC8E0CUGdTOuYqz4mwHAz6rTr
G9x1KqT02qVVo6CAbbegMTgb+6kfoHWxTvVJfSQ20oajgGiFA+lGJ3klMuT05K3zTdR0dx0UwEMy
MUKVVu8VwolSH/2sEHKNs+/Ur4T+VM41LIvcGBTiNYquOlkBjSTLojF6N15/Byc4d+iehBihtmkp
ZWewXNJKkSFSmjymVF86z0ArkaJQ2KeIi2m4rvj11/D/uAyB3yb4q6m9ljm8KQcfRGYitU18Z3sy
mstSFNl9Rci3Tvu5tuY9uybIEVoPWvSUknEMMeInG13V1s3L0qJAHMyfaHUI3PrDuiW9Z5COZylM
xWMkf4rD3jURJ7whiVJSyBvJeO6KA7FIXbo/iJf+XBa3bHRgF4ECwVRHgsd2mil9sfsajv7+q70+
g4jBz20hXk0VeH70Jqz6+XThzdXO3a7E5Mt8/mgk+u+RzNTYe6CpiSXOYRmCGerFfo3g9wk5a3Tb
eR6t8GbGxj+NHzNlfEIWxkw99c9Z63fG/XBrj1tq8rh/WLOErcM9/NEf/5C2rTQS5Pneo4I4ZD5a
mm6EpoFd/wht0fBxZARC61IWELbnZOuEqqfl5w8FKV6RyeOtvv5utpiyXmjyHEsfEFKJoe4Lb130
u2mb8JYOIJuEZQhHRBDp9FEXNYBtkAnNo6KkP63uhFCyVtTwMTJtvIoRK1BJDkU5WmraVyZK6a1E
oacP7IY1dfs7VvN2dIu1hxuiplb8BYTrEYiUWA0YNVFHWuLewT9Qv/o2A/+IgSmoJzxZF7l4rZhl
ZdC9OjIWP1l1nFtgWmnyeqaW4k4EI9C0yVnrdEoaph2Go/gBtrDSmb8MrYl/E4yRFtfTZ8n8JNIH
vmT99Lt4ZthM9X49APOb6BCSZ1O+dkbpHVdBE0MrR/Eo+E2ogmilBEU7wF1KQZYbtPL5OKjD9Jyu
BNgwh8tctPhYJ1mm5baynPuDKI6inbXqjBNuLIVC9mXABFWo5jDRS0V741rkTmvy33No3cUfuPLy
yTFr3UHke055Ej5MrT5X0t0yf7wKF/R/Wh0Z2dQ/c2aJJItzWNvPBYjsLqob/rTW0IdJ9vFTxLkH
53WOO1elAB+VNEP4QzpXbTGS60UICZwgXJgUEPJs5IKl+7cIz6tl4dfFv4q2IAMTGmJZSXdZFehi
sfoYBIHNPpZRrdcTi3Hhz1ctkK7kSGyyk/TKrNzbHHMPPepCps7WozMWzZ4k1EyHW8ClVl4FbpGX
dS/dgaWq0qzj/vBskfVNZu4OudljJp5/ySL4vfxnMBtCUuAm02gWp17PwbVaMCFKwTK4nPsLXL3E
kBjbZtZaEuhLGtLhsPsb8rp1IduO3WQq4yyQQOYirwQsV5KYJOmEl5dSyJ3sTmKYMas1MuYLV6uM
G2IiNMoQ9NCM2V2FAU/4T2h0Debr9nJAQ4WObRPXzB7mp22KVWxKK0jFqIaano1GvyY5kQB3e3wg
XXmkJhi1JE6r8/g+u6XLHADCN5hovng3e64d9HpwC5S7Js1WtZa+ti1EtOjF5E5c0UcPGZTVrysF
m4iDbJDoIWwnL+Md1A6NqEol5q4BUeQY4tz2Mnp1rPEGJKHjiBimSAzKoEELG+nkTQLVwS0o4dcS
m5e2x0jF0Wk4DKICV1qhA6DKNlFQTAm3mUwsEPHNykBgkYtFipDYbedGjWMftQ2CfQ+u+nahfHZi
bvnjWNtQ1U04GaSR/aX9sLX4qaT8dvp6ZERyCQ8a6xiLAZRT6GnE7cdwBKNNuTpYaoGIjF5t2+kQ
4f/GzSHw4BiyqPiYTPZAFEiwQLZuma2BjmTmWysBNF8J6vKekwDuE43Y1PdcXtanrqrBLobWBHhn
sDP+Wt962tF24y5TsA0o7WIOiAaMcAC7N3+cEPV1ztmbjUiK+qowI0p+nDrnX3wC/6qymfgHLV4R
k16NOTpfVxqIYZj9UkWLBT9vhKUc8q9ZMGWDdnYAlSzUe6lN1lUKd6ZH2RuRCYb6LgaIxc1eZxJ5
iWRL8GRChy9UQbcKNBg2Z3vUUXFZnRNRGC+x0+kpjXGyAGqwAjvZ4/uY9yuRWdG5GPA6hbtAHuT1
q88yywjJ6QpIfDC5IHpBeYTbU7XBedS5qq80Or9wfCNMbtbli2jrPP8vIP5AVZcP2M0MsbN6Wbk2
BvZBcj9RIzF76IxiZ09BeXFURlK49HsNxnBZj+EdTOWNhFzKo6uieW9loRYAKCbzEFk6GjyD6u0g
ZR64gRTKxb8N36jeTAG55lKIWNv2FnyHtm91xU38sMI2bBaN1ty3wjpGhlq1jFmioqEakTJ5gz9K
zOK2na0+3OV8CoEcEjMRXoMLTxWHir88YYs65lXc2PaEdeP70q4WD2vCZjbSZw0J3CSV79BdJDeA
1CibJHa3UWzFXhLDQsNk8z2blqD/PooxzZlrMCTAHiiJAOkra6A71PhcmTNNfxfbI+6MqDWUsDPj
SBxbxrGsoKpxobWkl7KSrLi5m57Zx8Cm7xcSqgN78IjoLhXt7JsnQncmaGJnAr/ucaMobRAQfP3y
zuSh1KpUQXHvGwi2e3DIQmlsshlYjuYDJimNOpa7itpLRGn8VAEcnyBoHcy1cJGHZT+DNibvTARM
SGU7vDlqLcMm6bCyYktdm+RmIFmWv2nBixQv1FRPdk6XozddnjP6d1fqmBvA0Ff3690H7526HjAU
CNdSrRXb1yjsEZOVTUom30j3rL92JpUmuO64oU7xlMtGJfecdkuGcTFGs2H0Yj7TiN+DiU3WSbzS
FNV3Ty+Tf5ohq4P/gb71M/8f7MrMWnGYLSou52veLRoohlDOwbMK8H4j9I0P7YJbsinu9/dllHqn
rg6UrPSvQOEtlNIYOZ4DGuWUkIicCt5rEAHK+mT7bg+b2V77eiFFbyPro/hMblcyLKoUZuWm41YJ
IhYsxj8hUy4xKPQi18tE2jdQbM1Yi6J+HS03HnQxaw3ab9cAusblHbgVfEW8d85kCM3uQ5oV7A4J
4j1tHYjzVhAttcYU3w8PglZRrCWIRspxMTxH/wj2zCmFznIf5naELzR9gBcmBQK5sLvse/J9pjWv
M+rgxdxb+vr/F4iQIg8JCIWVX0bK8QSUfdDwcVhDPcRkfgRirt/cPsJ0C+r96q/1Vnnpdb3c0kyd
kwGTVfUoCfmz7H210V6kRr8jPVlJPTpU93LF2pQBWKCIHTIuS89np6pHhUsy3va0O4EJoJ4ULfeJ
jf7RVmZBaCQqFj3byKLWQkW2NfbP5OrvMXcQz+vVqJ/H5orUXLJWpu1pDJsw7dzTA8ma8TAifykV
uMr+/Z+916BGQ/NJs8PyPtCTAH9xcNCQeHIYZigdLnknCO/wlB8wIY/hfC08wrYR+/szHsjmqsHG
uyfdK29XWe1PMubC6zK8u9XNE1Ry6dhZsaKVDPCct2MVUifzb82sQBwEVZfwc0/QIsdiOM1DChbj
X0zedUqlzMuqNVASinnuhDjq4y6dOej2q8c03qyDubAwcCdROWKmtrZsZ9++5Lsv4efRqO4/4s7e
lOMrkis6ytdLqqMEbyLAv87fMj3jRetEm2i/r/Fsl6hzklXo0uZGHgxwJ1TrTDh3vXIYZwNKnv2n
1sKx9h37uQXjU9u7mXVDyJHN8CzMlCkTPSLnd9u+OdRWJBYKimxwEXRFltaEX6bl2cABm2uPw2ZG
X+u/KfM/Q7+8g35X6pbm7gnZmBZf3xWHKW7SlBPrldjjC/pVFMr0i7cwytyS9dAJe46bCe1Hlk1Z
fnc/tbUXaW2P0rxoMCYhklHjlEuE5l5Ydh0Cvy7ofcXVc5QD69d3kqIMCE0xeY2SDqczDJbMjCp5
MBlPairgS2qjtBqzFOayE1pGewAE/Dz1WxOGBoGsQLUeoIL9iwNy9xYp1MJa+KV8RnfFLQqBJaL7
tyXTUTZTyvWI8vT/yqVylNonErjQplTCnTCr2kU7XCDqJ7WhR7JWmdiCEj0GqyHULZadcm4BvZFb
TQeaD6l3AUAK1MBdp0bbVPgWcf72D3MIoZOaY5bD6BxntraCvpkf2daJsVzliTRXRH5IOvDGEEtt
zF8m22B0oMCtP3ka48wV4UAl42qACXTiUDDULEoTDWMudynorKVbVSSIHk8rh6vk3Ml+7pR9HuO1
I9r4D2ecUHeyW3FjQoX7BQJyM5crMcFeBuz5TYPosfTOivd9a+Prec+JE2N4uxKIhO3BH+sV9R73
YLSZ4cBfPKWQsbQsZqMjrZsOJEkpgYLWruaXQr7UWg1D7/8aZIUwE+cgeseCqOZqum7rkWcggWCi
rRJLzaN/n4vs3M/rCcve38hofDgSoxm7BL35d+VHglUlfBBESqoqK+vM1hoeG3NjYhoxenA3iz2S
6QfeEcXbx1SSPuAd2esZ7xGQLJX7y83FXPJ3hNt+DrI2QrMvC2SeNuwdl22F1zCz4VjOX05reT08
meBJg1lvdzjpe+ZIYVMAvUxVq+82B+DTmQn5WqDXNhFaJrEhZTdmnu9oiTHUcdZbNePzTrm7rBqk
0A+6ocfgqFoN2/pFS8O8wt5BpyKTd9GKDQys0jos4AbX1xw7zrVZTo/daVKGtvzmfITiSUdrwkI/
Xzn7H16J7/bMY3JwC4hR2iJ326FXfJJb4Q/Go9mHvsftdlBLCOKKSnJ+gzyxHqnmfKzBLjDVdxwT
I+ZJyNK4Vb3qX17wH6VtqarevfJaH0A8qoXJTocB4hfdEmC+ZB8AQClWUXR3johaLVFizqGaT/qM
A7589G1HgnSoswlYp+HKVD+Xib++yKi/VtY/4ZDDBzF/PgcyDpWYDhmkjlHrBdCCI4O9aAR0D+Fq
uEfxXy85ZdMDJBPuIDN0KE66k3cJejGYBvhfwMQYBanr/wntmSNaJu/armuZ+I29zn9MyRVYrOOw
r69dgK0IYOHOAJmcw/84b+JVKf5ErFjo7zB2iGskjCe/vaJ3TmQ8nEdhs0bi5Pz8IsZbqauv2cee
0IGJTLtYJwHiM2YOXXFJOrePi52fG4BpDhYO+9NSfycit9GJi+DmMusFNvmZH3/OeuirbfaPT6nk
vVpxyBLt3ahDaCPw19jsSOMcsyYGFBkuLn79m193dZkIIo8x8wppLTQY3LWEYEscMy+LgmVAZTAz
bLlxKsxzMCpram9nyFOZHY8O/3Zw1EFim9mHQSnbCvDtTUOZkqyABufXMf8CoG0vkOzHTGVLj8rn
IhnBWjaZktGodd/IOb/UX+CJjhqJV4ucWMUkNhx/FlNzUmnoD3CBG6WOe9wRm5Zqj6t2vbYRAkhs
+uBnJASLN/BT+vnpQ7XeNSBPu5PyxWTmLMNORU4mygHxIBkfuBrt80tN6COmW/IPUL81Kjb5qnnE
9xtiKdz20XkrCgULUW7uh+cK/rG3CxETmoz0TLXU3J2IrKn0XBDs10pszDOIJPoCXr7IRp5cCKl7
YULZJwBaIKBP7X0Zm14Qao5QaypZ4l1tfBbQ4zuY31C6ezt5A8P97qna5+45YPzLBEXA/zvfc6IR
kqF/nDOBCIJZbTUdTijsHJznZBkkCsLBeJq4zjj8kGPygVCxITXRhx84vb28tXDqNYpsNKmvDgSc
Kf/tIJtVcVv4kdsVg5Q4vrFB9RFRYuwxXkBskb52VMhiUVJo8LJToJSme3sQOlrH+gIB1L8sIZBN
BRwC7yWstfwHQKVtfqUgZgNyRZPFuJ5YBHtBR2GDjQudGqBaT/VTyjwsaUUVnQmxNwAWfcWIovf7
SE0Cf/S9E+A+v+E6tH8O1K3/fJUf58Mgfqo3D9lZePc0gFf+C/ZOCmoJ9zmgSxxFe69Ia6A3j0U1
I083vAaGGiaiAzEMwaZPychONkpt2xclT9k1mP053Dx8iEu/1UbRE5tp8GlHcZMo1VSKXHd/O4mu
xvsyUuQQPguhY8Uu2TQhBff8+Ies4MjPF7BxRxqboZ5R0HzXbS3KNSoFf0eikBjUTYatr5+w0Te8
CwvSSHgBa1iLjclAiOEDIHPxC4SbbFDR6LKHgN230QDctINKQwBn+fW3Az2Gn1FtxuVY6d3/YbiW
RzxLNIWC02N3S0vXQXKC8tpBO/0TZ7QcUBpgu+L50ZHRe4uv3bjbVp9XSAY/5UOqpuhIdWCZigdq
qe8r3bMSu1L/d4ProWEMq18pFZjBCM1uu3XPOsbIzSZeC5KkSBmzQBEyF456/rY1eV8Y7MyUaVHE
qWZOaXRjIJRj/+IDMueBh86Oa36Se8lfRexxXSN+2Ssd8qIA7s8/gILqe3UQWR2VYh1GRilZxRgG
eX1EjLScJ64PEquKKoECIi5KULXg94YEQ/89VR/CHZjxi0lG1fEwUt3MksyQtdJGyXTpaeWldVcB
mSNXH3OhwiCujn/zim0fmP685spzuGcnnhrDO7a1RQYoUWs6dENMusFvKtM2hwEwfA72clffxU4V
BsWHLL056Ip/ub2aAYgfdaevxicNNDu/cUwhzHIRZ/yE1Xj7/oBLGa+ABoN7KiyBH84kJdlKyyyp
C0MDMNQ605ctJ3zaXdsgA36tAL/ZmMOS2By209tFFc22yVxpteTdTuvBQ0kFu85J60v5Gc4VRHhG
7v2ttTvY8Ppl/MRQb0zR/NOuzJGktQQWzZRkORfKugPA937n6e08PMQLC+phMukKi6Kq+xyUbb4p
0PnuAShdgDdVANKXcn4qqpwZPkfZibCwypo/Nx+LtTBhSaXFrAyo6Zb+LEDUeuiFrOh5c19wdwD7
dsCLe2Rj8vLfYvSKaDMw4dpCGK/wnln0+hcbcEiI3oiMFiPle5PoQU2cRIC4OVhzi8vIWHeAU4XC
GCidWPjPLzSCICTKuA7Oc8fIQwy5x1DSzc2SAu0pVz81NGNyrBAfpPhc9Zx/zjsq9DLcYjGCJRSu
GrMl8Gf5GboDQXfwQQcVYfUbqbTsQ27Byq7xBmiW9beo4U3O4kOqvja9rOSavKefq0rs9tyZ/5N5
sBT/4VvzMCAY01LnXuITLJbsmhn6PtFaq4nyeng11tP0XQ/gZ4Wr4k1A1ymx3Zv1bvlP++47nQpx
St4NkxVcUfsQ1HiT1m05cKrdd3h8N5KFVwVxsErgWw+SKtG8cGrlg36/maz8lC0IK6+o/0gVfHSx
0IjPLlpBhN2goasyOxnkXfrk7LoE2NyozXPPN5+XRgKFFCfa3bCOZ6jc8d7Q2dzDjyTJwMQEaYiX
4TqHzp5wj8OgF/1AGzE34TWPQ4UWMFl/fr75B8FgAue3uWpqJ2HvHTLFEuBmFzAfebyRBmP2rDso
LkFVwbU9zxxvSdCNgGEgFzgAxRDYoTCbjWNiVj59A98kCNzn+FdXFjnVXWSch94NrG0Z6BaAzaO+
/ho2n6CgKJnwIo48vRjVjtDmq0eJzZEdWG4wqJCdYp9FL/KBvytIbTbzO+PfohZvMmZbrKIINi/s
uMaFz5ohlulDUWQams7+hhAYMFASND2b9n/dOZEMzOkCv4rT0GOLEHssgDPbmPcagHZqGEQgRImY
CEY0TrqpzO88qVWfK7+4c3uKrk5tKddNUErRIxXr6HABiRsuaAN5qZZI7KHPFIIsEqsQG77D5842
tqTNla/omdU3R4EMmZHoL/oxnRV0T3ysjm+f1KsSCodlegYLESAofG28vbNAFNVHNTYtxxVIaB8j
w/CJFzbS80JrcgQVZ/4glNORwNnwwroRa1jqwvp/84vLBcJlywOJMe630uP9G7dRewinY845O4MV
nRKUhTGQX0GiDBXj0pAZRAygkhYiRYpOvza1ZrWmhCwNGFvfXWzpwPBDbKrpZgzMhPbnDpF9RjHr
EjQcSK9UU1Al7BuwEx5APslaavL6MK9Wz2iETod+WqMM3baes4p9OsEl7OS+9UBc5+eKQYIhsXZo
teFDORfOqZNUiUHifaX6iXwQosWsP/SU/NsU8wQI0FDaMToucTWLvkjCGbKXcBYyUmX71lJQQUHI
DNbIeUo7iubqppJzP/jRKls7q5RGWQC+fCZcRyeK4ESHtHVRafLMLo+f+zs/kAnzof4hHSQF4CrZ
9ZWxBZAzmruOj6d1qzYYkMYcwVRvueK87lwr5bv7ytWz7TVIqtBxW6lrbe40wvZ4z8D+HgQIGm/9
HSq59Pe5trul7Bz3G4Mz0EdrarGxcv2jaBoAqYYOQ06QFKxx6iMNnM1SLjDpsdFssGdukXTxfp/W
vxFT4HT+kUrS+UjolwKNWuDwjIgyxFg9yjgedlC7xEtLfbnf12IuK8mdP6rzHI8uhyuxDuPBd/2c
lDbDkwttHwZNxgJ9webfD/0XDKPR+TGqrOTfkL8jEfj+86UWTx6Qd2DBTFHacec921KTNndGncc0
bSPL3aeEZE/Ks+KAboF6rSJTsw11h72RTXIh/+Vf5jk7v/oK3UPNMuB5pmG8/ywtYIShxG6EBJN9
GtME7wwAu5V0FSajpHSOUBlX8CDieDoU4vskQvFtwnwwoJyE5onrDeohKhkT1u/fUEIoXGVTv+Y1
592rUGv1frPxDzJENZCmeDwrqmqyJ8ME0xiBwA+2ANlGmbirWKaBfC4j5N43MFQwe7raG9wOTdTf
xxaYdRUcVzlTW83MM1wGxFEpMgQxVpzB8rq2t4Rh7xWyl0y7g5M9nKVofFZVPkGhOtZKO3/OCMIJ
rqaUCgFhsDp224F9D6/G/65Vg/7tXJqd9DX949busVBeAUQvFB96LcvfAENuaFdyPaEDXJS34XxZ
R2y4ce/kYUfjY3UQ/0WAFhiUQsrO/7ixvqAlI6Qh40OUSRE0EiNxm+RXrMnRtR0+yqJtaMkndvbD
1cJdfZaxoXW60eX4yuhV5xpgA0igO/eANBsIXWToKZCAZPdZNkNuavXODOniIL9DX44coTAvLcEy
2fH7WFOHEbkt/MNXa/bkzXDMfDST++CDqgPTAXXblVsUE1KhFeR98k9dkx1qIAfPz9z9YyrHxJfb
zs7TEbNExq3qGZXadG+tRoXATXCxSmLZP1ca1ovvirfm8Fwt30Ls+waBvvbXFF+O8G+uYGWsPEfN
oJvP+NSYO1wcRoadz9zbNcjbRP4muy1KeBlNX5co7J3PlhIBQD0C0BXASGbIj1nmWZ6eT9LDLGqL
XgA7o35DxQOiPD9NCe5xCysuM3+Q8rUtgLJjGzdGBgSnF5V3ft+jyUH2mQBCYInlgWImW/gf6UzR
DgNr2OpQYWbx0pwwOy+S90CfoObtiHiMne0bjLH0fXkcUjweYaSwgk2O/WsMoRdunGRymG53Fm5F
weGdBGCnrSk5pquNS6VJspm1e6KgPFf9q8jVndHNj2hna23Oz/53QjiPl9PuAZB6ro7uw2MGtmjJ
dCe3dWfeQLI/ly2fDAA4ArulvAgZGtfuLW/i0k3Oa1mnN6WJYHt7dWYPopXEJL7w1Vr2v1j3tj28
lL5zfyLq5KQTSgj/PXHfq6ihwjcLSmIE9ZkolPGTRI6NUMqfIkwPx99frYmgZ9wqtk2C/LyXg/XM
bMsyjOqedytds5yA7RsLgYiEXWWrTtPUTwHE+q45I4JX06V6IPjaKM+o+U/i4mbU+Y+ybsBjoAM0
mua5vvBA5brRJ/+l1arIfNnm0EkGteQUI1PHoBdZ1EWSna0ek66BZrUd1PFq78r+4S4RjH0Csh3v
6o5138LT3EkKJJQMTSRnGMC4FQvAAjkThsftmBQvu2KK0opBNmnoPeMG/o9uFq0LMl9TkuDbzh5y
X+fn7ta7Rj3GUmLCAoZ1Yj7nzQkXKst8fwWxTwjyTAh4730IjQkwm+XabejyRVoErqOcAXZhjjgu
TWiu8MPcVRR29RKtowU80AXz8yWspowsYRKO6Uwy5G3pP5WJ6tmiJ5KJHfodcqzhN/o3O80JxMeh
f7EcKBdx1iQw9+gf3HnySlg+on4sxg+r8Z6AxqmiNIZBkCuRpDI3rax1ixZIrkDJwktWUyUXtqul
GuAF2iFCqQeEr/7Ltd8D6WzTwebaHnBMB1FQe8L/efJxp4d6OcIHKdSIQYywtzmGeuVfgk9AqVRd
wcPN/uYouIFuQM4SgwajXE/7p2gjHxmPJ00kCMYAciJf39k44LQ1rDZ+yICO0S82rKMDbyoJdt+3
F8IJPsBBx9SSrUcbLQANU1jKZtQOBfBdv8riPEQ0dHGmtzdLZabea3nCusW1VAVLGUC9OnMJtz/z
zcsoy/DK653Ebww7kaTCZ0jLVaSZxDX2VxRBQjsCMA/tqED9I/zEnun2BNNINTHOTW4DpGt6WDs2
P+omzl9V5q1eW7RaGWv158owNqMAoCc2t++mMLLAm0leb+KWV7GMNufbtCZRVbgOdy1jpG8VD1Ac
lpzTAcRLn7FquhRinrDWlaa5ZFnx6+sct+KUYOXh2NMx7t+HjiyS2PL+sy8Fk+ylxWTfgRw4i4KJ
g9eL6AKD79na73aF62Tm/c31T4cx0mdF9Ckv20ZxlFw9bUbKvd2nRKnQGo9RMQLSjlLEl1sEvaaW
0+Q4veH0VHwjpZLJtQoic0mMCUsfTIojoJp/IE/zjHraAzKpVBzVK8niEzu78MTbXLXSh3HIv9I9
P44Q27gLBgKxaA2mRSWenkETgmCIVKidwqwT6V5GUaqS/O3CkpXnjxJadV1U3HSgV92sSPlvzRdn
BT28pXr2k/WwcFx0W9zlNqzBxWtJJcSvRsdXi7MSU8mTuNX7+EujQxPQwNUFtXoLjVD5+DMHGKxm
ktRuq3hiKAZIzc5eQWnHjSIeLWRwo29ntirNWbHMi3MIdhK+UllLIXTWkZtr1lZ/azpc2bMt75b9
RPFlGjF0Akc3g/Wd0hCYk+moQOFL4JIjORdfaa94jd4KGbeGa52VEKDjHlJIsRjYX8/lDIclPJSW
uLwXjEiX2xMu7FvaQhmFi9vlnhw4mXWgkQzOBE335n2FmsSSJ2TUB6j4YVu8vi2y7iF5I3uGXLCQ
NzUORZo3ZzeAPN5JdGaT0ynBbOrTWOcFwAx+PHqUhF47pwePaVZwhasM1tDyEjHWQSys6CnmwT+n
/USdP6BWwQhjwzr+dwxfo5kRGYkNgky3Wrr91EJdY23Q7NlnqIkY6jXhegpPCqqZ642LfLU9tLhX
YaRcECmXpwy+0+5e84FZbp3lcmCxNchIFSdz24Rsd2wcqDkfe2YAVquOWEynJIdLpTIPsmdt/SA7
sSqgOX+hjtnqlHV4MT+8Q69xeYQS/Kc8DYxdRSYEsbSVWsJX8xt5YHb74RHXHE3sHbaG+1ht+NQf
oBKIAx9Gt+8nSRPtFSrZA7diOOG1qvNV97rcRMskwCt/FVYx7/cmrLf+E7Nfs/PZ3UTQ+2IRquAZ
TtaOM3SoeG8TJw4GnA3twnOOzjqxWNwrmmzrwZFKW4fT26oVegI3LB+XbSLnDJp8gSiZ5mLYWu5Q
Llx6TdblVpmyvunVTg6JbJnss7JDhx+6qazbFoZFb2oHbcIRgQAF+QXMO9xqbR7ZIDT22vw6fFUF
SPrMbf0mkc/Hglt+vSCRGS1PRU7MMtbI8n8AZ4EmVUdFmwCLivMrnD+qXfdWeCte6W/0WWK1YJlG
C8aoz1m/FaAW6HpND3yJe9Qpzspn9pgcvm4dhYbClkPJ4SKUk/1tG40ZV3DSm4AesphaSn9ynmqo
KQIfyf6BRF4g9L/UHDUogEdqUW9Jy2fvPktOQMC5NOHWG0tOIfC7CUTXKhQZ/jt5q1OXztKkURft
zOPsB/UlxMLGI9ldXCmzOQoqfmfpBOo6LNrZ7j1DDYi9qjIULhPK9sPt563Jkraog3gzwVKQVwt7
TFzJ2P9OGE+37DGPafB414148rSsMQU92UqDJyeqv0dU+xE6TXkPKkMVTKCVFuMYIfsNH7SoOU6W
xW/J38Ul0RMsL5bulV6QCrVntU0cjedHIqhkIgZW6Bh/HDMyQvSDEWCZySsYyn2QTV0qcZ7yjEEA
rT3HdO1f6LYSnlyg0XYGqy+kjMI8/cyEWE/coTTRMODM386kI7gesiV3KybnCiQgYJ4nW4xshdZ8
lxRijOWW0NnuOVJOIyQvCLMpiuquoSBA4dHxJWzJQq0uBqV1QKHnN3Skhr5wnZUslXOOflUCcjny
1AOUztUdS/ts2fhWJCsbhSSPoTfNKSaRrlHaWVqWYYwFK6aKYi7UEBEMNe8hN5sG+p/1K7Pcvwve
hDVb+7F9m5jrT4yoJdyhBEe/kgRaz5uNOfFR26T0YuziU4hcPRlcc35GvVRb4RX5M+/4L2sSM1AM
1Krhg7oGRkaI8PpXfpgqTS2L03K5Jyt5bGVhceWoeqdIuL498+Of2WWR7CLsI0CMmrfjGH9CmSQT
gnYfr19wMhu7t5hfkM/dANZ0KcLngRw84VZ4GPrmjsCZeLmQfvypO59Rk9h3cgZ6BbAtvSimlgsI
V2nhYw1Qwrc3An9vYL/ErBm30y09DrrHAxh8r+RB/7C1Liywc8kD2jH1FzwVnDf3l2qwpQxYbxuf
PivAy5GZLpH4dxFveVCislESDCr3vDIg8CilZYSzaKvyGw+l2B0IHi3adW8a9LeWdFLGIVRrIgTD
DGlbK+krruIKpKztXdfnQCY5tLPw6Iazmtidme8VQhebnCe0qHktkaJx6jyXAALPoe0gCknDsfo2
fPvpe5X0an8nXjSgPLT5pxak2zsXNODd/av5nv0e7k5EwE51/7/Mpt86r6thtYaIXVuV9svYNRjL
ZuHlTWhVBxRltFBgU699ANIavkfGeDKhz+IufVf5vt5ZRAr9rHtDzqbvgYCCDGi557RfbM+dS1rJ
OH56uyoJtp2uSkFdcQGKXwaLNoCVhBHkmSe3kS0maZv9jmx3cKIoB19aAQnyFe4o7F84rxpdE7Vz
LVsM6uxKMvqkwe97m4vLkXxcyv9LpvWfYNeVrXjMNohmJUs+Kmf/BshpA7UGG9C9v6z879FhkwFJ
66rr3QMl81oAiIyhHyD5x9L5ipcK9XxE/604o1GGKwEZhoEVoTvJJCjwVyEa6R4jvMgx1mjxqfFp
rwLmywx/zKWsFnO9FMhufX5i6A+Tp+LE0KTOFra/JlZRGy877uTNRwJBwXg2kd2ZadAEx6Hyt5ug
ZcTt4KracDDi1bl+bq8AfrvsPvByO2sP14zjm2kxfRb67yymRciH9yrYUmL5bb2QYFC5ClLnjdoo
7RBBd7ZYroNgbPvU3ycfJWFA3EZ6IgcJk4h8RlyK4karsaywWRn9Db4bKmFTcd89uLp9IkFZSoFo
GViWZf4OKP95RmTuOSpP4/D3/poDME0sd6tvkvCzw+zfOS44PBexJcjZKxKrgnRt5W8XEP+n7Nwt
gPaOW/4IB7LSzerISfQyuEx3D+Q2wYWux4yKl18jCkzYO4wm8fucl8esfNupkyImNWFR0jw73Ls/
rfDjNpo4ZZOLIhOnMZ4wfMfl+uco6OYi2+5PiFTsxFHaIWrHAGJm7kz0WnXxnn6wPKYzGgIiVy3F
cZ63hCHWySP2caiRpwyB1NrEk8qWHhEFsn9Va8stY3qQFLP433Vke/6sfMF51OYSwVZWZURPRX+W
yPjotVa3oNYkxTNQHpVEpmYz6GDDsI5t5W1bBwY8TjaLwAy5U3C69Zgo5nUUpvaaVS6s3iPVOevE
NGCcNQdM1C6v0Q9kHEM+3+pI1B3YiCCmYzSuJoOUGKJKeKgAiBIwiRrTK/HvgPu5dbLN6Efo1Xs2
ryWcp7cpKYtlBZyU2J6ZtHs6UsGm+IPN35H3xxZp6Gv+DRWdJqkZfV/G9O5lWkhfZg17Ko3gmndf
eE4fcxF2ksOf+ouEHxKwYPPcBDiQeD0gstGdqOIVFAhoWKNcYaBYzunTzmRuKB9j4EShUOFe4PMQ
hmGO+IUBYMBRU1PHT10RYMY+cc04LoM2g4IHkMMshSWZRq3gJb6OSNUauJPJcHIJaf0cSzw3BARZ
5F955Byk1GV5pzNmobcLRhk7zCXWswnwv2i694hN7uQBy/TtNsrtxhICgjpbb56SfZw7PEr2XABi
UyyrrUhHZ3nJC8zOUrs6rK6h+hU5eWa1dirGi9OUfTbcEz08P4E1nQ/fxmNw3R+MyLB1n6NNz+BT
RnVEZjH+B+EiPklKnwcs45kHY4+mGuQc/0n7vtuBMcEpYUYDmPIwYayBZA4jPvZO5/cG6Rl5pVcW
gQuFWxwWgHRUpGB2AWXGLSDyTm1gWojMsmGmD6jCQQB1x+W9+g0w1vT8AjQ+zn853rOhUxkKSwZP
PjaUJt7u3JJWboMxjXNZ/Z62rTIQvi2tKAHbKfylsCbRNFFL2C1OUmFUkVldcuRngIxCc2q20unL
hbY1KoGSIqyJlRqm+OibmRE20HKl30I7aYmjlp1NKpbQPChImcPQ24wJJCpjvhmyjZk+zYqp070w
vU/YWGbZDSUEytVa6DZTA9lsdHYayw+ByzzPGcS+2lcgXebEs+UdN+QYr7FfR/Ovxi++PAF42ap1
ZWwQEVFGFIMAdTG5TOFkEh8F4W63kcvLvWNacpowj6fzrp85VKJHO14Z7+4xZ+kVJYf8vVo+6pL8
xMrTa6isOxIuvzpaoYt3omZ8Nsk05OhjJ5iNKtp67dLlMSsrnxKX+gHbV0Vevfasyzz9AwoQHhNP
lVbICVTzV7PCmVTH2zxLx3OfLBkxALc/SCSIMIOZQ2vAnoxNZPmkKZPiScSlnq1ATACghfUXtEfG
0LfdC9oLtjTNvAGKb1X1+uMNt/Xu3SoGtgnwmBhh1xW0e/vWNEDPbhJfPOHUqhEc5SexkaG/f4z0
Bw/bWfI1xIQI18z/vfZ9w8ByjdVZOxjLYw7mCgMq0OmsLFzp8vkeX88qbgkNuOadOvdsaN0MrF/f
aKi2cBM5MJnkgs6i7bla03MZeIsbv9+ZNJYSS5HCKG70vqY69ZqYK6SmdO3I4OdkhLva+mW1lphS
mi3RPwWPeEg/69hJSSL8xNazfilkqLtLDfNwYa9Ofl4jAqed1TZCM+yLcLjko1mwrM/OHffPgF4F
NqPS20iJAHqgJgOvLw49R6qOErC+0qEGYG52omThvLI8nzC7eikLoi7sM4OA0/dz7CCqVNysDWbM
iiqypdClj2Z8GTwQiqlAlOL4nC1YEZEScZ2aw3+AKLM3aVVZn47Q7s7JgEwX5jYDv8bRVtYEjZrR
tTkA332VKo/QG/c3/1v6T7Oq7iZMpzBpqHE0opQnbK7VDYGbNHnsa8nfnDesh+XZr94LlnijD4SH
wAy9TooTA1LpEfZHYeu57GdRDe3+R+h3e66huBH2Mx7qBdWxueo7M2KCwHo/vXj9BAjbK6KGZYLA
5B7HfoqBSZ6JUfXVwxBzZ7MRtGxJGv2BdW5X+fpe76NB9Lx2nur6Iur4Ou7be87gs40CM4UfR1YL
Z3w42NDXyma2Zfd60NK6LpAZIwCwUAhS6SJrKNCxgmLVRbBCI5fu/IeCPaCWGRytJj/0hqvG2/ha
j/+T+fg6i3NTWy1rWJ8kDsSQqXmRUC9acHcThvT5G2GxLMSXcFTtRDMg5nwc8JKkmtoiPC92tkzs
hnwyQvzKqv9qcMNUSTScllODWhPw4lErCbDVgQ9xG/yKJcynDjxbilH3RuLf9cFKxUgB2PeqjAps
o+ZjSmf3hsp9UuuG1GKYq25clkIwfZkZpTv1Ong0C7VLrr3foJvT3iLi+dDO+tgcBg1fpgFy8ow4
rWoVT9bjBggAG8DPCVIzOhT5DBeNOmfFzLH0+ZWQFsTy9l3725Wmsis11BQyBv8d5aPnTDVRWacC
CgbuoSTeg9VXuoEHXLaVofU9Ey1HOAqKjzNzHrhRI9wfdW1NMpx+dhdlLug6iV22Wl2i5FTaapyZ
JbwCpbYe7Y9sKaunipBbK92Jqxcy5bGoL+OVAt8I3RjSHLKSvpF+mjNdgesP9hkfK4VQL0AfvI9c
brfq/36ueRx8orxJ8iJRdR1Kf4ctkO2Si4HK67coHoblE+olK8geWeozlFCzX2u7DZdaW7s0fyL3
VtkRUPHtl/hB1ypolaoFGqn3Xslln5ahv1Iio/1LZKGTvUt/L7blpWeUw2KnfIRaJpoGhiIciQ5g
5XuxXJ2rLoE1iY7EtP1a6aUZR+ciWORbC0vYxLrF8vqla+80tL7sByXjt/AGt6R2XLBepambWkc1
bIpY7syoer/Rt3/lEneRJw1CGAapfSmEHEVvpEHGBy4X0FHnRbZjnDkiDLGTjhOndbjFzRjBpeI7
egkSZaBQ7CH//G5wX3mUGN6XjWYeeu5QDgOuTn0Q0kyvtxvEgGoLQcURXWRyWn9FN5W6YR49y8nZ
VMgxJIGhQdu5k9nPBgb5fCzsX9wcGG/PaukwkV5+E4t/AuN5zrr6SBvP1MgqZBfvJjk0IMeLwhqE
PqqlKMsS01XKjL5EWsYJ2sRtJ3Oe8TUpDNi3snWD+z2MxTtKpqNe93JEPk3+KUsSuyebxbvnsl7C
p6JRoN+e7OfQ/aaTanXDAwHUIZ717EQOuxyusRo1Pp7lJbOnW9z9nNGNHs2FqGP/URSnl8YQeRhD
2w44T8Yvv048hwvrj+f3VdpPC8dcHFTUD4fODoSc+4WERJfiLmvQg9XY1QguSriHTkeM7zA7ozr0
Q9UDNFlq8sC3vL84ogUaW3qHW1G9u6xGphA3x3W7JJKLGo19m6LWnoV0oN0YExmVBqkvcXKNYO58
K2OuAZ1aEoy+6oDGqOuSEBn3banHTtxIrZZlvNd++iLSHVdHYD88LxRcP8dAiCtrCvF4KoIRWq5W
Ex3zz1XlMTZRo48vch8y/RbiNXlOqzxeKMrUIfpdEZzmWMMuNGM2vxq5Ldfq9nfk2ROZyX+0xVwN
RNbJ5vEN5Z1s3l6OzNlfZB4iYIDF1QgbM3+8SDloRj99wv2iQzBUWLl7CKmDtwWrmZeE8iImInx+
kQzhWeohdc6pDn0kkmyh4pWuYH7jSvKOFQ47DOQHtKss26sIRdOmijJrsx0M7PfVbSYUbaLh2gc7
vxU3YHsmqBqV41LQp4BSrerEgQDXsk3SBzQB8w/9vwKCeE984G9SPXOxIECNoUD58jZ+y3VDXmKa
ysZhGx+Y/J4izVw/Q7KAVhyxNHUHaU6Ky5KQSeQEZ+TMjOq3lQd1CH9r5rrP9/isq2xrXnAO7NFv
8KrXv02mZIEpnjrFODdepMO+3KrYg8p4GKr+dXCusIDoUV8OhvGYGDCoFAldLu6QSGgrQYlSd8I6
+32DBc103Ws2TnBluQtpNMOANCUAwHvJmOnU2dMpB8zbwSBxdjmlCMuDP1jLVQDndhb0SJ8WwUVo
OAK2yFVe+QOPewtnpMWwLqxGN7w9IOkdy2DHPfeqN433UCPD07zRY6wDa3SvUTi7qKu50xLyrOGk
ScURLnpTonh7N6MdZnlQhcL0Rd5T4soYqe6ChPufsm7G0HAHhTKBP07pxa0xe2KqO/4CeaBXAvMu
TkKNG6WzXuurgVpK4fNETEvdnulX1nZVFLxPDFxmxoQsguzYSdYr3p5PWcWnJ108JczDLf2LfYJM
v9VnOyqUzzsEMri5xnm9zPgj9FxajGDuzajTag7x2eKHPamzW+hDAuQXwZA504ZcrR5kFTqXQli5
FTafUqvzvuIg6b7LMQT7OHx22rt55a/mH6N1PJPm4cNr7uo5ye5OJbdMx/+x6kS4iP05Rut27YmV
VhRT3XjpYHLODiFU9wJwLvlbw1ZqAAFKzMcWt+XKGlRPGvBZEtBZEOV78hqlPq0B/EK/rFGItlRe
5DR9cTU7v97YiLwTvrxS86Gdgyu8fdFbrQ4g3Wgw3wRljDccVnIDdM9fp6gx2mI7k1VGxMdglfoq
cFXfR87sRC28ffs/NJFRbus0g9orI9TRUZVgCbR/f94wHqNC+XVHaTr2/d1dFVR4YzIQ3/qO0vm7
/2G4r51qng6zcF3WFNNXmqF09MJTvj8sez+oQ0fgSWjgsd2lKVf252bH1p+b6HZY1dPUGaa9bF7Q
cu5fRWnh5QvI6LgxmHQXpTdJIgrmpxT1Yivm9XTZSAvDhWw9I2hOrmqJ2ziFi/P02i6byy9TKlPv
lcUAEfVyw7APKdZ6eroL2p4huNvDsH9GLoh9r0axSngIgEgukjn33tHgeD6tpF2KB2qu/WCAZM0i
NjA5wLOanSidEVSibKOq563FkO+7suY/+Dp2j0EMsq5l8LYoeRjbc469w/tZqxcVThUQY7Vtsj8u
0EvmeTY8cWEZXDe54WnsGeYlsc4cI5Z0XVAeV0o0kGX8x8riCsBt19NE3mtBqzznjvJ9NHJXoI+Q
Qs+Mlq3YkLTv9qYER3MOSFNpe77PWPKsLYCRl6NdoaoS+MHITeJqJav4o5YqmfQ7WZzGlOSvfDS6
9NaLlThkrtam206aWLBtuCc5LyAhBeWip3KDQwra7LL60mfI5RLovsS2qZDVwbyw49N+z7GUh1u2
/Zb2WvsjqJKjlI5bt6Lobs8WMv14YVWG+A2eIXzywLoOIG1Pe9LAxg5YA2r/ww4e403qaO/6ERL7
4DbDAXan6DHoZTDLmq6yRXo4HI1oNHDM+q1RSi0AlGaBbphX95bDMiX3DMrbIwfUop3Y6fjvlQn1
WRxIQb+BA+pEmy6UY9PhprBrYEpIJESdZircRIYfDQDWql7DvrDVVIus7BT4bpxDXc4v1+SsYBvv
hSHf1CzAoKWSBhfTYc/6E9dy0Akt3JA0BL9yVu2v6u9aZag5w9ruluh59oG3xbkplzGiNy4kqHBU
+z5CzeHt1MzlbZ2fZhlyWmTYIti/FYHixBwMEoUdeG8gS3tu47zhJX2mTtxcpT5xy5IBQ0HvzW/B
9gOa0GkpGI8BG8BkyHLOd3Kzc6zWso4MqGCqCrBU4kUctRevZm5/7DMH3FlbC0g9jBcxK2WLH3ou
FW9mGnigz4GWM5v4tDrWR17McLoBIv6/KyztSF4wBAmNH0u3Sk17VH4eybFqiJ8cQCiBo2e+LAOs
kJTsVRSbmhaIQQr7XMqxwpgoVlRs9VospYH41VEJuOllhH1CVW01WTIz3/IM7nJEGfxhUoI0Vg8l
t4Ro6Nur1utBZciZh6ENVSCmmSUBTO2dOlnY0o4KzVyLVD0vLlmzpQHmZE2vNMPInm2pU8m4YXdp
w9oCZoc+o9KKuJ5UIZrdbzB35bPrcYAY7fWS4p/s7m03NaAtaN7aDhxfBUHU0ysCEtt4ReDZkugx
hBHItqBETwvynVeY6QVsCNiUFWfayrrsgglLed5N3a5wHQ8jz9tkXVmLJLTdUDS6GmA2LsqWLkkm
towEkbu8ek4a5A3xzJhkyhKjM5mjtUsnPmIKTwEYM9+/UYagzGN0V+QPaJk0KzHY1zhgGgDQtgBQ
WcN+1TsaP3IlxUqcLeRPEnGUqw26MSH5HKfLK7rZBs306/EUOSiVV8gOKDceyxfhXvJTa7jomFgm
ADuH1x5yoFdTi/NunhM9z/N+glMO1WR9TLaycsNUmUNLU9Ee4FXke1XVRBHAjOPwzn1EKI3VPUjY
6lAP+jJf2kYV04Jc/nFNWCgICoOWBicWa700KCXTOJDuYRJl7OuaAFgtyE31Wa9zQuWUddrjG/yM
EILGX33mYEmNb6IkEZfCkWlJFZrdfzM5Yl0bDnfDDrEK2oaIU2q98gMgeZMbePOx7+rdilGS2E8R
Qr2m3anLSvVs8dnc4GOE9L0c7xYO7fbnSFwWOrWqc0O/8eL8Q7+uVAHIUyrQiONnOl8wb3LTl1hG
5vvN7hUDZHzJZxSi2K0K9Tez/zhc8U0Z9D2IKs+9fWl3Te5pGM+zO3hlGVGWVoH6/vk9852EzyMJ
huWpWVXVlQ1oRFXVzzDhJN1vUVuVCO0uK2MqbUkwVfDr8ut9qLv6eV9HjKe3qk01OWwA+IDXEAsK
h1VZJuQQWBFHXGcDkrgNpkWTFAFrI7G/Iv4q/1g+ZRAS9qpAZwIYVrGNHX9KQ4u4N9K6glARUc4h
UFyFLjQO+akCQooXNUDvd+U0skcQnPgn+WnrWRv3KBBig0dxbhk7RWK+ECEvXnm+J+mnN+IaEgoX
r4iXcnhHFZpNcILkEUd+fWu6ZRWMuM3hsLWKDMotkCdHXLlkqnledhkUVrIehzadgnFAszqa8eYL
Ns10z+313L6FQH6aEtvv4bN6T0mCZt0tIT4btY0Udy2SYPfFsmBr+6omyFIOArp5d1JnuaPtoRbP
UUF/1rRnhxFCWuh93XB14953pa/YR5sjCrggw1JlctzIOzSC2w0tjwwZPYYPQ/TCdnNETtabVo81
hRijfpuU/wInXp5beJzIdoRe36Me8JxwyHcRPfzyP+p+w0nyiTIROJCpdU7RXWhcViz/a0YqCKHy
K7MMsybaHT+Q8pL6fPAgPDljjWj58KCMlI+ax3mPEfWgjVV6IqArABU3nk7ByWfMd/0B2y5Nq82q
5iHK3V7XsvlHgvaE0caWYiILY96YlqIvlAc7ZEvlHVDOHcmGQbxQ7pbRCsgJqzcpWIWermOMqeJd
zIYWVD+dCgIiFbirgOh1BkcQSixGZhqZa+mhIAylEnOSSRH1YuAkokji8z6EybNj47D4N5o+itDW
X6UJYm5JNoCgRxqCNa6sv/AS5RrKBXPTHmNnTatYhpk6zv4iA3Fap3ObdrUlafVrzT70Jsey2lJo
FgOCLTuiFQsvHkc21UbcFvwZ49mzP3KNl6PfI3sDwDlrpCYQLXrSRT9JXed6aDuthsqWIvpGqbI9
gHZ36PKQVl83nvvpQDJg1k1QRJjDECZj4lgksgpt05WqzBLjpWkY+ZpUkQzZnT0BC2sPLNkgZMtH
XVjUnUxe2VOpJd3nagfMgG+YXElznHyBnpENgetd2fal+b85DEajK9otYGhEIJigcL5xm+Ms9IX5
v9WwU1T4dwtHea75X22BNg7uMptJlzStIN9+Swl8vJz/umFClJbIf3M4jKFBMe2Tk2etmQfVGG5S
GO1LYdX0cm3BkXwwzmfxc5m5x8iDxhqhYIfQKYtPJNvkXHI1HyQ7qzGTDgcaZ3GRCrV6MLV3ACTG
EXL7rTPtQ4GjK6u880kBbidW2v9X7LB/WLSbwpXhAzkEJaS1TrAa8seAMSYonyksTURXe/byqYp5
LBQMdDynlfUDrxBrfMWSNaFu6SkHP/I/1RhRsNqajyhL//Yk7wEwRjN/aF12apj/DHBFfEe9H+kE
o3XMadVk6SI+tzLMOrPVHgg2z7aR7Rc+3a+9dF6EKJau4Vam6b5tp9UQWfz8FgQHs3kF7A1oK8av
lCuOTw0lZwfKvbFxCdFjt8GDFY+t+ogwZz3ydwFl1cVjWJbLp2Y+zvqIBdYYlkEB53i8dZDpFy1v
yBGNYLGKFJw8l1VgDbsSD3NnNDcKFRvfauRvOovLwpHHIKM3QbJ+VtojYpqOS5dOv6kNZHtZ493m
7kp+oNAnbX/MeDrQZqMCkp60NywAjZEGgcuZxposDxVNE674lSTtGW3S3NC/okVY12YVb0IoS9Hi
7zu40lO8JsNZXPTlz4uvW1G4atLxtJcy4LWATpngUH1Pk2P09bGby7A8EDhHxlZSaNXiK8n4l28e
9eMNmQ9LIwiezZCtIGmu33A+PiAmISbUBf3CxeRMRLwjXbyYSofb5f9NHM1ggNuvT68o9AjPxCoh
3wpxX67S/DaKcGViNlJBfBINtm7gSnR9tJqXTkN6Tk+M/ZlqUzLtueY2RSW6OSjLMFIIc9DU0Ofc
iOxAxF3XDb0EJLEQ+VJHFAluSrQUkvwRKhB8H6m7jt9mqM2kQfIjLCZ13k1Ztfcj0H/Je/8EctJV
nWRoiBNKEF/SLURae0ReWu2Z0F+6VFAXmStDSznnDI+UwtC0uh/gofW1rTtkQ+b6OT0FUbPuRNuw
UgbqluFZD3kMU0e9k5Ecl/RTcbhiZaIlgZPOtdiC1fPo1yGGXs+sCrY2RCbe8SWR/6/y+qQ8RZCh
ZyxWVeDydTPK7eERSnou1G0133O6qdOGmVtVfrH8QfQKtqJ0Nqi5uWKTfogQBuUH/7rqIArU5Qb7
LQCbn3gzGpZXTJRTZqv8zbfGKEUUj30w8snxrbQXQPZBkJDywTRPocN1bubvVIlWtgMlEnLjSBs7
WeroRV58EANfKRiXKJWLijxbbaFqFBpS8LbdsU/0dxuriONw7mE5su44ZAInshWHkU9PjLktRSbQ
8L2TuTBcSuVQ4wsku3CVfVLQ/yHT+Pp7/InT1UiAw1g28mk/TiVC6zZAPG19g0+4nT3Sjpg2AfBy
9GljZVRSxSVnSreO9YwvCHYI1zUIu4/2nDTEfXEXExEFYRTI7vEy9k8d9Nlo2KOBl46OLdJndXll
5a1191gLcPVNMD+5K+a5piUuXGcW1LoCqVblVSbE/tKTm2ft0Sf0E8Wwco5KTaJvKcB62SrwhQMl
0wthRWOmX2rqRqxC45QBbMqRM4GxwqL2MkfZSxMMXIDj/vll/fDkMxLAmLlkYCoPD4+Je5reFXDx
kd8tYn+ugTaHNCdvF2fbHfBrHT1xztQHx+WpnSN7YRj/c4a6pYzOUBECtlIfalfIOIVWbJsbTeQD
Pu3MwyE8uPDFGU+htU1XrVrBr0rZsaKJ5SYbt4Mh3i0S1Y68NmN7G14+PayDZlSlNbPH5bBUQN2i
4dpPQStdEwAn2B9GuQNMN3oJEDSvJufD6A2sPLTicfqubFeBS+NVBIHBrE2qTqUEMvXQH0xixCQN
gbtdnpKt5eLb6rswge58YTNPztotbnmkCnyYFtPeVUWgWB3jGMRhBAzl1w7QgNNKX5ren53F8Kzo
WJBj40iZoA+411aSTztHQvM3toDgCTqczf6ir8ARu0uqE9D/3tjdpAOUSkl/xVXJPXPZJIK4oWeO
M2Bm+zyiRsttUbEdj47/o3VrHqsgOSzr9F6p/HEi7OkwDHYiZvcQSppJYzDQ3ePwL8q/PzEave/G
vNyW6YzMb0vii8qZ+3qBSyKbUGWfbt17lw3S2v3R43KUjubV8aLaXh1z+PDq+4R67LisoFOQt+wq
8zVSfp9jwWg0ybXX89+lksnRQU5n1J3/fPfcWTDRJt3Z0m+6VT4wUErdLLwxw5bOEZBKgMqbLYgI
1UUm2Sa7kKELyosDJqSDqzDNoNcbQvYK8iArgpVui4+PyWuClIR2HPBFSt2Bzjo9JILUub4Aa/Vl
hNuXlKd2jHANpplxOmQ844SUr9zAUmJtEbcmfQBv6+a/eXHiqrt58/bfur/8A7qIY7lPeDR7d54x
ii5XpUESOooSYf7im20ornaWx3aPcco8rjqhfziWC5ULaLzNbj3uLH6m233NQajEfQ31ZfWGGF5i
6eNldpViUtqm9phv6LBLz8NAhOTuli4V+mM6P1DTlId4jMJRq08vVEIN7WN3pj0nxaamXOJZx6nm
3Ur1nK4LTU3J5kz8e5WeWf/+ADHydsJfYJUlqPtGoWLCstVTGV4YfrDJuXarjDua8YpQ/IXXW87p
G27lYxuKbovh5AePz4jEpT0AUHVLdC5lp852+FvaNt+mo4TIyOX+yQLGEDvcLQOGJU+vT0kvT2Vz
RNmE2HqS+MUsvmLVK96sppbZrOjqWOWtIp7qpuRufiTXRNkl+8IQ9er2YITLarXBNB91kIYW4gTv
2gdxFDqS9aWCbXZH9hdZAK2M4dsTT5okGuIJLretp8OK+L5KVtBltpoLZ8UJfU00/4zQkcCf/l+l
qhhw0qxMiOLT3W2w32j1EXaUt5DLUfdz22xomU0MoZQIuRkDL0MedyyM3AiN0FCqBb/UEYbPqK/t
S/2w/ffn4jOA735ANyej7Ibh2R/o1axWm2BnYtTQjn7GxWhqRgRMchUDcBeDdNurW2Cvqx01a5d2
RYKqMmsCgYCZ022UUcu5RakwsSY9jBAx21/UUPhRNcIdf4DjSTEGqeZwE4z1GHfpiB6U3pfOhYPH
WuOngDa0MLKe3ksJ4iCUmevTrZ2f/XJhrNBWhqjXpOombeDZRjqJQDvaFW8GT+gGx7SiTzieoxUS
PLJs9LMH1TUKtNKAi8XR2gN4f0MdiusI2DBOMpVufcePaQ6CoIAWOuFHU2Z1IDmp9Md9G116HicS
tYfnUbUgc71qM6ySo25D1Me8OFTsHbEE+RJ6l0VXi/WaZGVdGcMp4bHpkqceehE03s3IoJOGnalR
bGSMIDW3rNB58PC9S4r/eLRrxrH/zRjFPo5bZWYuY4zVaFmN1NTcTnSAWNAsThgW3NBlAy5NphwM
DKdEA1acls7vCRDEwYQAl37JACyYBKxcvaMVAvvHVp7xrCGSnLmlng9UWdP3Shr5iGEwPp9PWAkj
z9sPeaJEGCcgOTOQood5qKpzNb72caWlbERaC3c30wgOnm0RCvYCKWy7apwT1Fi7MbBnsm1v7aJU
75pct7E9wHidikKmPnM/p8JVApoPbLNpxNJUwCyfzLtRnl/NYPfY6IDdUzy1xtu5bl12zX0wKXdY
pGhDkTvtJkHzvT8/EOeoK8K6YpQy+4edyNq6cXmbmGcvs8PrjvpBZA3h11ohP20RVZ8ZwnDPzDnO
DxnFS2ZNZfmEhqV3GwdGx9eEMkH0nucbwOsJf2924PMkpqdnmzWZfJ2wsTK6VnvaDV9zqez48oM7
Ye3d9x6qKNMvDFr6sjgWzE1lku3vJTFpNoaNex4SL+5Vcy+60WNKgXvo5NguABVnAjzmMoat0SXr
IYmBD0ftyR0HOBxNQROyCANa7sUpIeRPkRBRLMLwRFah+esrYB+WdDn3eXJzhckS8rK4fAS2qFHW
q9ULxgKLQfNraPSu8S7Wu8wwNwXf6AY97Thu55SowUnkO67VxOpXOTVBX/ism/I12M4LsRTAllev
tnpgtPY4D8vntW+ZticoV0HWuzRznQdG0p6OVgygZXB6UiXo2dbw8+tqe7k22K56Pj5tvEsMRYvn
MsULoBKqJHFmGgDM7AytOuD0oQxOytxtDrjIkYdq1sthJQy7bEQRfBowmVbDVydbf9YC4iAm0oaK
V7yr0qCgXXnVZx9IRjcui3JkBXS8fqVUWS4HuP6QpZTrKp5uA+PTsNOB8Rq9zc4VIMh7x9VJfFBp
MHylqtk8DDo79OfisEoVdZjsNe7EtF6Cf65YPNttPdghp+vf1vtMux5hfE6TvOWoPGCYKk/uuPSp
GtojxoIaBsVy+3NMuqtMe5594grsjdRha1/S97zQUIFeemCbC+TmaSg/f2ifEFCjex26/+d4Ih3U
Nmph2hmTZunhX5adqXw+4ekpz/VdHTV+V3uI82azShPoMDxMOC8zVVWgVvh6hzn2l5yy/oiTRGKA
W/BfnsJIm8cGYwZFabdb7USLpwGjiot/FhaLTMhEURvic9K+e4HlbH0D+RJ4vBcWDgHMcFTaBWLE
N2SaAPU642SZXnqKwMAaj2Gq/jb2f1GHDmuIeIEdBB7gB4uQRCyJUW4kKMhOQMCyA4L0ULjJFzZN
bt0xr5OkMBxHCvkKVpgU0/I97WEu+rlknqLo6c4EZo/+d92o3EwAp4Ux0v9ZL7dzOfrdOgCf6TNv
i/kNgcylk726nmzybbLNcJqUTL4gyIBadpl5Moxuq87JDte7sgxYl1khBoV8ALBoiAwxJ3CHYdOX
8in+QvdSx7qbS/B9NwaCr69PvKXYYMVhqBgx/xTcLXiiGdclb1MdntdMnSXypNSBfToKqezTzO0w
0jGPtYIJ3F5SNLxc4sOJuf1ngtkJwASwTV0bFbfYJd6boITK2fnMSTjcBpDlAT/RY5jTZfDho2sb
KkD016sFepERhBsU20XFMlW+gahyABKyUcSVjKugXnfOYd2/5dzlIZQYCjQWD12YjVFk8j2nEJm5
JDKfqOL8KWiQRDsviRP2MfhHHanLeXAaK1xswDaT9AjExbF3B+7Wn2TuVrmp3nkMpMufK1EZL7J6
mFHylTaCFT1UwqjQLSlnqQsmktZOsvolqKz6Br2+Z2zgmRedPfhr6GDi2A6rN5CoHZH2X/in+ypA
R43aXs5/5cJqwAu0S+i6F9O/+5QV6Qi84fcIkbI7QW+SIs8wYTd9lfsElhq1NwLsgdv2m/8tQYXS
T/aJB0ruuOcSoh27GtNbasULrcYqu3CZ0SLqUOCFaKAYwlOBxZQk9pDai2kXA62RMoIg0TdnFVZP
Vg71PKaiTcIXMlLiIKSM8cufOFYAQKUaXbU1gwndnAFq+/cK2baljWsx577wrMyrxjHx0edH0Mv0
bjIBOQMeY5Y2of3wESZAPDxiHJ41YAJ07yN32PrPb9nCOrJkn94iqPrmj2ZpMB7HjuS3Xu+mjpBb
kr9+OOrIEKFRcPeoqoNdTvCPCAedmOjby+20jqXkY7ieh1jJ0r9U8NegA2pfwYnG21CDz/KZWyhK
v03M4zDy8hSht+1In1+Fvqqyen1koYMshSf/IhXnzT9RJWdesd86wP9LvRp2dtE9nuD+sXFTNNa+
92jLc6eR4ucWnTEcL/qqX5llkHdn5y5x5N5rX1n6XHsr8LtBehtJ3JA8bBKm+lmv3NzuopHRJMDl
LKHlrIephBQVt7gZNqvtWRNmh+P1HLo7lOWCNADxVPNh4JbZ6LEQp2DBTGffpjDXdD2yPyKAA8gD
e5qLjMbwFY8RkcnNqeJmF1TkOaimGUP12BoY53l9QWCBcOCJJ8wdu6lhfkFKKNm1SHR1EQ0I3QI0
BKh+lHJdZxZOiAfQxby5rMjOzil7YEv4WBpux/HOi7gAJdRiX5SRMQEZXx0boVP7+MMsKOCokRLX
Uglf2zN6VybAWju5XRvVB1iQMcAX8l2eCcvOB5S8qAlrvtdr85A7foQoLRYytTcEUXTyJzFpOell
JIaFH68D98hGBXNjuhIu2N3/BrGF5Pkd+8/kvS1lCeYT/5JNvMWUYfISPISLhmYSrBJCNAx7sc2l
fbPr8Hl5EUZFCkDzLsnnV9q/JZYGlGM42T9kk/Mut60dhP93jJAuLO6v0jz9rtv5dZcAIBVRQaRN
vvEQjZArzvJWTYp1vAvQFBMhazGigpebVc1cA6UiHd6Dd/8O1qL1H9EF4rbjckPDRO2tmYhk/uQp
Kg5Q8B0IuDzyfdDrEvwrf7HaWD3bCu2HyU/if9XBEa686UFyZn+7OlGtq8UxyL6UI9ym7DiY/cO6
5v1VXbO0qKYYMn+CMhGVyIYbaZiJdYSsKrJ1PNSffc7XDhAhTqScyLQ341JUO5+rLzJkS9WXAc3k
5QpdWZmVnqAEFEjetxGSPH9uZou+uNJe0N4Pw34e/T7Kzu61Z1zp7B30g1lqmp6lxcyjgFBB0ewh
BLNn/JU7A6aW3JCbWakHOx7QHW3ufyXfZbBsmhy22NWHcTRly6JWrtjQ9jIoy2xBVUXYKR+C4p9D
JaHFMU1cEKr9S1a5Ist6yCC/KOhh5uzIX4j//VPbZBe4M2Sb/ixXykxS01yhlYnF7cr5XGW6sH7y
9YP0Umx/nzj+d3VnwTZMwv1lDsY5AIZgzja4jBY882aBahhgkuBsCL024OTcJ06HRvBdT0oKBAk9
rYUpRMQzg/8MnQTY8Jxqo3X7QVL2dnk0Rc/CNklU9UdKnMXjmlAYjlCxTNFYWd7SIY3GhKRb/1IC
4arVUlvgCUvIAenCi+cR8zyo4kui/Hj09GfpAkc4cQZjEQL4GEiUtop3eC7OWDAQYZZEr4FKMteD
uh6ONqGMkeXL391B9p4P4PaM7CHGGqNuxLlWYvT2xo2My2RYT3ler7aewCKpg0LYEMC8Ezsg7k9G
A2niblHanncq2BformCYkMDsk/QMgNUMJof90YuisXZ3tOb6EIVqva4Rxb8FrH7giQbgFWCDGllZ
jb+akMtn7AQTcRoFUgkezidqlhAGSWIassMSqzNggzw3sUSWIIdY/GLBbUkXp+zSBYlINgbvLd1j
G65w3nrNc628A2Vec9HdJ3CrjKqgpRRHkj8FVoTMPFbQpQF6nYdSwRotstiqvKwAmcdRMLRNf0eg
7acIxe6mqSx1pQIxzDUytCshKlnz/5U7ZCtNsPM53fzg3sk+eGHtudd9RQEac8m1e3FTjNUV5BID
EjMjvo3YOWvBVu0AH3IAfo83ZobwP6kyyusG2MEXrQs+mu6e5YdFoXwpo1nQrM8lisEim5WattDm
Z5TiBcPbmuJ7rjEfM/fznVtBMMeDxAlmW2VCfAhFgqrlW4GPhEDAFMkj19jqUhmVnVM/LnSy/GJQ
atH6l2BCPDPjShQV6HMRf39YEibbPhOK4fFw0HXmoM4Ze9jP06BU5ZIM7FknGDfOUZnCM/qe4BBP
nKsozNRlVEDAtS/77wYrkUscdGiJYS9erA04BScS8JbsPP7g4wp17hAhZ2L23P6wi/yRNZSy/y0e
TdAZB/d0iOMzZJnADTOT0kJxI09/Rx1zDr3J/p09OAj5D6OEvVWIvEBhcPEwdTUDLZzzBYr0LGpJ
s5x+ZFnNfPAWQ5yd9RnmdvQdefhmtnnnNr5QMJGr4vR7ClcPxpZtEVLG9pV9UetUDrNiVv8LxoU1
+C1QvhRdSIKr0Je/fZKHKrQ2fyVMuDCuJgKNfbz+NhUwYN9yRZNesSy5NaAgtq3r9Tss8eHO2IHc
nSgSiOBbDJzN0hR4Dqg0T6Eu8mfiOza3aUdCMYJkgp7SGCKtoifmnTCG/Hw/dDHNu26s/xbdF/2U
WG9HvYqp09nS34YjIgpE8jwAOGYkud1xApIVahpbU3GvnsEsqW7SmO5chJPzJ4VK/AE0dTn+uUbg
H5eihW8mX4LK0yNN3kkMDouYItVP332RLAKYi4gZaPr8ZJfJr2ZEB2iYz6TU+1EABZHLJR/aRqV2
V++H6c+G9aNu18de7K+W4/FZrwFJd7/AxaWv9xS3lmS1fuXkhKg/wQCHxqnw+AGINO0rYHjKV78r
bE33DWrTo17BdFCSIxSFaD5Bef3X1X8VkZzBJzVDu0lZVZFv2q642W/aKSsz8ewiqh0ev5gYRcEM
B/z6qCN9HudX8TNtqlZh+1/1aJA6l+OnYMxwQd076gZW0QLk7fjmoa4rYUJ2/x8fARLIWMDGi7hI
n/yFO9sf7/ARHHEE9/CeoCNGMwC3eAEHhcBUdR/ehpQEmRJD9tbLRoKVDjuCbI6u/urqzDQftO9j
wYxgzP2VwrEucZa9z069EUqF5atC9rCIEujAU/Kkg/353DGzpxW3PFbiXUHCPSxXnhf4u9Xb7pnR
fomkTEJjv53syeWL7hq8yOf54n1aZ7IT9yGt14iIPg+5QVtj3nZr0ZXOpbEaCPP6OvAdeoPGerWB
qb087ZhvUj97HsRE7AFe0j/TqgJL2LBx8ENBCLfXPx2e7F95tMmHSlrE0r+F1+VDBxQcfvI2hBIa
8x/Y26QpSbPA6zkhhx+NGrTfvhnuzUs8id36vACP9OapEvyt/mJu79ubcXYcZiDd6pgDHOjUKX3U
tC15WRE/b0xJPvtXZbzcYyJZRwHkkJiZx65kihvYNlKDWNw9KY4nTknhBprzEPGZnc+JMC9+g82g
Sv5i094qjq4AQJnPcpnKETxPJEeTokB088Nflauyi89LhOyLI3wXtOKQVpLXtX0t6krZJLlM6iFj
RAQZUuCYMtoumyhcXqFDU3Lw7315iIPuHpDa/EKTZdSfuX2ZewyFfZSATZJNh/FNm42hR2oH8uHi
0BFU+n5OqnVj338Q7/vyoSsNKrDPcCdFBgLgoL62h5L7krz9lt6IDrXV2FFJg09FIRN0VlCxbw4B
VFh1WRsNi80TXQW9fRCmhB5Ux/+i1aCgg98JKQuKe3Z6k1MsiMUHFRQZ68rW1yrK1q1ZNHQjD+Ho
7K2dQiXWbnwbuYtDb55YFqvyUSnw1kSu+jt92NDnA3t1+0Jt6JmaTLGfhjzG9tRMX/rUfEqTWBDM
BBQGVsPWYPtgzj6EDe9CqCXVEDW3w8Z6ux8LbaCKLH1ABpGDv3GU72AMRSv8Rl0MSv0eS1MMbKJf
tBvLrjkmHWJMUvn5Qlyux0vmIMs/S+OqPaG3dCvR9TLCOZkMTGJgpkZFFhNCKb2imlIOGiJdI+2W
OTzQifnvCvH5hyi2DKw5nGcq1R6voS0N8NbAbeEzOZDi3eYuE0NUTqt2mfpvKKUGgtpOQz1BLpU7
kLKSYhCV0gxCYvP+TSUVlIsy7zVrwx7GGNfKeWXW68IwTnSHqHIXl6tJSzjDxefpyOvnj6epNuXl
WIiz8OizFu6gwPvis1MMR/NuYya4VESDmh40lnELJxyYcUxbZjN63xKGdEFElfyJSIO+oxizn39U
s2o6Ht1KXzofCks9npuzHlIDYiP+9iwS7v7L06/IogQIovQD3PSR7SqsZKWTK2kPCLE2amInHjXR
Gq1Be8pHv92PsjYVL9Vy08uLv+AeKAbu4F23oGBc4wcybaMokVa7YT0Ez1bCfnODhZCdC9wif2C5
B47qg2Ly3ciQzwsMmPO2W/UkltDa84wTxdyUVJMsdGvDKf19x4jJoLHVNBd9oB8+gd0547rmOmsW
nALSBOOCC2k2agNa7Lq4XVwvRy6sgk7C0ax49c5GjPd8YnsqcE+vB69PJDvugQPH8WCIr+FuiFD1
SPzPPOpJ9TJTC0W/EzwoEk7w6WjKpxqoD08GeuANwB5b4rcPTEPZHJYAyx7D7FomD2bk/rAKFyZM
aNMdj0HybdejbGKbtQVtLd/OVx23XVS0x1yyaB+Zvzw6aYPShc6LrucDuIK/oAnNSdMWXqloehKG
DyWWZ8Y6TdRMBvE3A+qbKsZYxyq8IMuwJz5ZXkh7Fl2l9E5xcoGtG9dxgeXE/caWLsTGnlQwjFWm
7UJPGXDc1RnHTsfB5WP1eye7kEJHZmJ2bQSdt/sR4aBNMN30Eu6msLnu3E4vv7hm8veB7pARNdo9
5mn/+HtDdPntvVRWNvgpmwX+8dtUC1dT5YwFjvChWbtXDyJ7M+yyzX1zpAWTftxdcmWygP5b5iEb
mqOECyNoOeryOQ2RNj2UwrTx+BQMFKFo5FjIQeTkSdzRHhiDKGtqsi8tCY+xKOSKT1bVbH+Yj/jS
DjHpjrEhTyqGiU4VxTdPWCNHa2sAK8wzIqz1LWjgijCNRLmS/T9PO23sRraBqvQVdAGTXg8reeII
Ou6Qv79oqbD0enJpX18jV2hZwG3QbD+fyICrmxe6sTwRwqJydovikW8f0YcP3wy2S8yRfa38svmO
yGTDITg3p5cmsRRUg7LjAJSd+h3wvnuM5i0F3F57lK+oXBBCLlERUMUAlIJHUU3DExMH4664/M6e
QGxwspxO3Opj2FY06cyYzYeaY6IqIcT7OVeiScf0gpgma0Qyo4AsiP10VET7NdTtqsCAFWU3pYO7
OUqhsm9BDj3tfk1UG+YwzwtSqGlypAnlvwCCyMlL8czgVagMQZIAsAtCxTEmXFSzgjdLyU8Mygr5
L3WE7Wy/Tiq9KKhQQSBrecliRoj+mD2jEqdrS/pOMK/uzibjElfNpHkKzvGBrF9cCTIGXFDpa5QO
0bAyQzjpO+Ehc30J8H4nQoKaZFQRH9ra/wVCwZsIo4aqCdVs9lIeWCwVdYe9UBL0chMTqX/yL9hz
gM7YM4LBc8GUyfJLc6LHkwU2JoBuEZ15T8Pumbl14xamRoFTrKBN4IWS2WR/PuEWK8n5Y7Nnxy6e
bhS4jJYNEN2mfVMYxzExy3HqLwJs2XJRWZExDIF1RZ9nFNpV7S9ITsjKHcrhVqP/BkgRLX84mrFs
Bi6HWZumoUU5CghEzYdBzW3aPxYx9XbnUVo/GuDyey3vKne5yZSJE6ZeJ20cQ/PV+A15+88uqD2M
Bebu+9o8/QNW3LoLq5tsvGeddkNeGAOMAEqS14wtIOpMz1mNAQPt7tdLc+FNNYQPZ53GOWudaFXT
HB+Jily4HyMzkZKiJmKwE5ueNratark7FD9oiHuEWvH79YTqrUI/mjPbpZ/bGMLKsf9NKOC+qSnU
v58UmrKzMqQ6exRXQasXRlAI/YY9b4mGf5Sj2k1hMab5NHXYERauLq5Up3K52xY7oZQKAiE5AmCy
/QBemkOqDQyQeNc0JJdFad6v4XadJ5jlwyZgArxQ0D6v4acJ+djS1kIXgLmeU9GTIzP+3c/goiYu
JklfevlZZQrAuTWlDBP3hYx8JWPLp5TKdB6FpFWr8wKA6kSDxvijqlDHNqw9+1iD+NLmAfDywj2m
5Dm/Nl4tBM8BSecGEa77MN1p/oij9tZ2QJe/J3WzOzlX/0vFWs01vF2l+MM+wg+ZHAmEt4W2zHqq
fFL0qtzfglwG05aIGSm3iMLbAAbw5oHxn8nLKCMYsGbp9YG1457tlUIF8w6zHZMlHL15MqQLYf1o
niVnL31eBVU85Xxl+L//w/lr6A2sZi92EZxfnVHEpN+J283sY+IlnRmp3xtKNZzi0iCQGD+Vpmcq
LN/Ud74b37IGLyabTMzZeQbBDw2rVjzY0Wrm2Flf6n+8FGZSzea74nlDfq0yeUbWEgsJGiv6hzDJ
NTLosm2Ggud3A+BcX+igS4oNlCREzZTioLZSvxv0a2QjrfjkQw5lGZvzSSGNteK2gFysCZ9Z5sS3
XyRb0BLebXivCxNnlZcDRoALM1knKbC/tQN2K3sSWOBJ1CJG0DtynS9lnxeeRF4mrpMYnsVQPEmI
hyPz4LyDygnsJ696bXBYSvgBP+Mu3CbRYszPRmiVbnGcPeTIcAPPM6kp/+2BnvHNs179YRCBlizt
cOAzYEkCevUwCZl6j1vJDwsTOdPkSgzTrDSws4giMRpimI5rucz0eNBpeRUWfWNfRoWtRvSHBfdT
K1vLKztXlMkCRzZjw39mWKz6+ay6l+dFhPHakz+AtFHgov2OkZZmqsPNP+Zda3NxyvfxrAv7E4eA
9U4T7EGvaodHKIKD7moj7VmTMyZy63GLb1sPDvuHPUjgIh6iG6eiu2OizxiupYjJjdKoWgaZDKot
8p1Dkkk3mtgsli2ebscukyZQa4RgrotgbsGmtFDOJz5aF7TlC0cchiN6Kc4PI6v2RL3J7FR18I24
QgtZh65o5AftXsKWGwMYHe6RyKX8+QXb7vvt2WB6O9smTtsGjnOXSj1ynxZ5JR6CAbVvW4qkBgWB
4Yqza96nnQzO8x/Z6t/xDuECHCVKTrZ97GUsk9HlxjDrSfolZtLXFZLp5EnJ4D8u0auNHLXGaAB+
Tl2ZHDLGseK7eeMuK0vW+wuIlYF3M6rurlFbhI3CQw5MmA5gkv+py57tFNyXj4eexy3Zerla7iWt
A8eDb/b16dG+K4giew3tIegfroI60quNEkRyywxV3+NR6bXAdUj3QjHuXHW8XQAiL1aanIu6fdxo
W4I+faefTQgW3Cigi0zOivFoY3jPBhD6o0xl/jYbK+6BciX8nl9dh8Ug3evjZjG8h3spNi4IMFcB
072swMY11kgMl4ezUP1IBJjvdCC383CCRzsnJZY8GWZ++Fhkvg0DvCiJ8g2VtkIhGerGWTUPyUCb
1TqYQjHVMmV+1cGHJYz5v5P4QiZXavtP4ZexYJiAIwH02LPD6BJdLUbQkKsAo4fkeCywOAvNDNnD
VZJGl+Wzc9MsyX5HFut7pM7uc49W9w3MAS4qCGqCANsdYbI4X+U5ToNbkkNGB5s3mekNJDZvWQTn
1SghiCx86szYmhRiV0AxHgc0r3TQPF8txyPZLpYbKdBYBZD7K5oHv6NUmhwydlPSi2T/pNAfY5uv
4D0SYsw2J+3bv+lt4OvuQqG60W7LzGkbabHv/0MxX2uCKJU21bqQSpGNFMe5R1PRC0eJY2FKAT+C
qClJVFydI/2q4p/nYl2xjj4ve+wlkmSTqpCAROhWE+95GJ2UGDsLOAA+tomqgfVSkNboMjp7M/2P
Av8KRWcpNSvqAf0rDHLj+vCeKFsKtqxrchxucCFaoas8xjiQfCLcjFSsTt1wFFsZ8UCWSwjbkP0t
L8dJvG+YSIseDwPKG5lX4qSkJnvc5UDqMVuAOzqLOQdY/isBqpmcN5p6FZDaAHfAbttP4iwgGBnL
G3c93Q6LUIyZYAEcEglRcq9bOfnWNPqSLppGmfT4ukLnbiVvFKy6vKL99qf8NwWZ5jzYBO7mOQuP
FCiyrdGoHY5hD3qaTjHrOuNESc/0UCU1R1S9P9nBFZdk5M8JjFgsN78wMxU86vi2wLj6jUywS50O
gVVzxDDZGtdPuGdbk7EaO6U0fDPncUesQlyCR1wp47y9GRM7+U9onWGFx/n+umi3qbojd96PLwXi
qF1Q2SqjJUl05vmqNvxB4I4Fr+4ZODWbA50CS19F/s7GDFevqGtSnHksl69WCuck/DXGQcVtHEuC
PfDFJPBvpMlkhf9ajqYqk7F0CCHRyHJfw4v9QTQp0jDeZcj/ygUWFziIl4+RQlMWVk1zU7FV0V8C
CSONMGBi+7SD+3sFSXIsyWhFHXwNdmwmApPoIqGMgiwYch7GOfqKR8dyogEYtqmPmVwbAAUMGGJF
mvcYkT6lwJj+i648isyIxhuiEbuP2ZqJBLuFnsD9jwPMAAgnbaYzNGcpEl030Ehzv9oyFsabtJLe
W2ll/cHA7pdAd36P15AZawm7esuz4Hcmo1Hi4qfsi3bdiNt9ydH5myVGiJfyC4KCtDocmhzPB7cG
3HrW6Sd9xy1qUf3uuDlpuEmTtkBa7JLFQGzds4psuhVkn435yQp6hfN6WxSJQGjma53pxbPlM6hX
4E9G0evJoOGv5LshOaXZJ4B1kVA/w/+yUq3RZvwf3v4XkfQLjGBhj4QaR/SDK36OZ9d7Ngue+0bM
9sQ8SMVbLHjyyRlldkUaHNqg85Dd4RT3Ol6FNxmUVP9Uu7zHDIIptMiPRcgfX2ipuYuj+sDRni6I
xtTYjDl0VwQ7U5Cmoidu0rckSOe6BOf/b11+CsSo5U68aIeMxaQpyLBq5bz4vTlVN3MFE94zA1jE
pPu3PpORj1ZawTzXAdzhc035EYRqLjRVtfBKp2o9OtSilCCzgbXaKQCDLt7fESPgadRH1gfoIYU4
mZ0UG+zmZMGtQjdfoYo5Blx5tAm1a95ZPkdk5jhOEiyRR+iMOFAjLXrPDOdQ1197mbuuDz/H2Y2h
mXk9wpGs/qwyikVTKR89oCV/S9SLFnr6MXyR4P+N7ECqXdH1gcmKFfIGTeaOFybSyYv2mFFLaINx
DnuQ8S+IYpNm0KciDvBJ+OVfAyW64F885z1RhbtE5s2B28nWlIjI5U1xUAlpZ2P0WxRFJeozErOc
2Qunq6VPm6efbHsUcF8E12dnIXPZY5r/zMytoiDOFtS7b0ruDZdTacuqaeZpzQ3gv3BLDm8tx0et
DVqp1P/JoqMxX01uty4rYsN+gxn+Auc1J8fkbvCZwqiAkeaetL0fk9gDues6k89VUHa8savbQLV1
LGBpwzFJKqJgX56x0Uyat9W0cnVTZklefHyUHjJKDTaQexGc0mtxNYdbpLD/WbuBJWDoXPIvO69F
ImpJYUpeXNg1x1IgY041NBlnUHcUjmFJOMZ+wHVt4Z+aUM71J/E+QhoT9D2151mhLiiw+IG0iRD3
LAtsfb6Yipl1kNpZTxcjgzJJdGjwVyZ2N1qJrrzJgfTL/sCIa/p9uT+1u3gtJ7bcMNRC2J3gqMLR
8MF0s05z7GDQnmgQ1L+q8SeC8E7QVRmSVHcwzFsL4+iE6RR8Rg8qmnsWeySWiqgmvTKk9sBWh85j
I3pk/0ztAqBVunJFd8lEbrEmLZBp0Jk0QJxTMLvd9PN2JfXlG2jd82NHPywTnxMn2WcR4fiObeMV
Q7vSsZdVukV5bR9xgOF+CawHcx3OdifxvH5T3DBGoQPm2Pa2t0f7+rFj413cH85d2rghax/0sK3e
9bN373YdtTQO6oWNIsgMYTx7Ecrdcj4QB+7LtLR8qvvw3lbiAWERa5fGRZwCBcIH9EAfL+QDjEHa
4kIFoLzeHoPuK3H6QhuNvCCVdAVcZuGFJ6fxI0xTcTruq0JZt9CPwEp5Rommcj0+1LKorgA8PIoD
4vxn0t1EGUwemae2FISwy0Odib6DM0DNKFh7DozolkMWPLJTXrLwdI5inv5zZghvEExHuateZYSR
FANogIhSWWcMJ+SuS5I4J8eJSuKkNzFyka2c0CJr6Vp1RFWUr8Bw9zqyZ+xC9tJSayvBZqnpUFNA
7QxwgQFY3LQZw9tJf2L/3JI+h/9J7tec2whiNzgkn22oYvtuSu55wY8vCwFZmCnJ+SByHv8tBMaG
gbNr1z3jczmnkF6gmgsv/djXEpvdB8TWh4nKJeGv2V1+doADqAXi2FEyviQ90VGYz+nIhedZI6PM
VqAz2ZFgvgd0ip5pSPhvvqg5bOywkBXIAS/N6Fcti8Jx+omuNB3QyMPACOKI0gmwjdb4faXHE7lT
1Cmx+UZ6+wraM3PVg9fzwg9vlM4q07Vq+MZa/W5a6hj2AWH8OgYXUnehnDy4aJUE5bm6MD8anX+9
4HP8qtY9HsUxqMXjSU/6UgO8ZTfgXShklagbKFyjae1B/dgV2rA3NapyFJpaHUGLUJ4MZfZt1SgY
YLIouWvOdCXtZasRQ+X+/T3xzweDdacPTlQfNl6dB1RTAT32HeSgw/AcjUFyPd7axswdsWXSM3gR
GGC2SLKLd2xgIcr/NKeXi+tpQ1AJ5oeB9L4D2TuOup8UB+29SSeDtl8TKEUa2i+t3LcTHCHjDLE/
o5Eftrg/HKRD+OpdKunyy4D45Vsm8cmX1BrRk4UWeq8qULIe9sXd3oeKs94Ubbjt0Td8buuDs8OR
qHkrk2OnpV3sX5p26gYAcKu7RoLOMq5g8PnLjtp8h/6BMHudqzTIkKz7g4HUPuWi74q8gAHpG8uP
TwvfoOo90358HZdUKF6A3382eCpUP1Nb3JIcAuHegdtzGJRwNDHmz6XFs+i8kf0+VSPO7frrIEAg
xV2JIsyROt9hBSw3hfVKEHi+tLfM4lx7KyDRyI8edoCgDlyW31ixQCqaVESBNCnvBqtNToDGcN+F
hUdVLAkiPnjyh+KQ9AlRRv+RfzeHjBmrWxOafCMXygnmLdx3qh/cWCzuLVe7zi2KpDdAemdYcmWW
xMOTXFaLkd8pCoz3UMXXohHYeJEsigUI6fHc1xgghwR40l88NvexCvXaIz0f5JecAQogEkO+a5Z6
vJdgIrVklrZQVRJ2aUhqLqIw/vbPtGGB5EcknsVl23C8egJ54QJVIK4wjUrARWmN4j4W1u18l5nS
ce9VRTcIxbuuu8TJbBotXCQqxRlIzbjGsLll9R1X3FSiA2BypitDQwr1QuGYTVC2OcgLy993mPGt
6ZVGipR/MULoqjnTfXGEqvXj4EGcNro1BtmmTm5ScRWopWM0IgZAZKRW+I2zONaU/S7Ru7mhwN67
wSVqKw9MeN/DMD2urR2mveJ1kqAvF/rqLMS7cNE3XMpRSmKz53NsnXvFGeKgEgLslS5BW6X/9VRk
wPIlP/nXaduOZKNHXbZ8TXykGQlgrGhxK+CfWQ0Nk6O1DjQNf6eiaE0oIJUYCjH9+96cmoMog1un
4dd16/LbVwR0KUHk46mFOq1BjOpv7qYU1ihxiwzEZQvxhOPrdOQ+oHJtGxD5ArTQ3SDcHCEUUMPp
BZ6IRHcB9Dgsvkp6o0Op+xs6ousK8Mqsvlgc3BMifmBLd1kNxSeLob1fy3SasEdiBdZBaM/R6uOU
mbVVGspKwCKqkXgF47W3mtR6utXOUYNFV0idhlasQoGdm6q860nTWEQ7rqS5s0RJTK8EPbSsNOJj
pr6fpIADKdclM0/v9FY1YNVBtxo5q0X9ci+zzdJs8TwDqO7W/kEbbQog2qX9zESj95kWonQmTBdS
X7v7t/YVY9fMdq8PzZ/Dm511Vg7brfa4Odh4Wpb0L4KaJRuaAbnDjJR6McU//T/XNZtchSk1/2MG
8/gcgkW2mmonfJANqT8Cb0oG3R0To6T/HQyJxr9no82GVgOp5oBHDtbBU2ZfJtWOs0A/vxChTP1J
DfCKGy/EFoWFjqyt6s+3YwnSVLw6GJX8HVQ4NbJVgBYHJc0ps0gCV83eL5DrcpkaOlbRNDT+AeF+
ZW7vVWbywtJUyO+wvzuIPTVm7yZI2gL91ik8U5/bKUiahwxty4s+msIdhikwWyP62UYXeMxrE8qb
dja3G+w6EE1ss1+1HFFKXUlQTnQ4cYJ87HUFtO3bboDT9ZKbTafKqTwDVHQdFTCOljcjhFo+Ne9v
/d+z1qrl/9lphxzHrqIOyWA7cAPQ3cygxjaaPfoBiqfMxVh5YXd1/x0jZMGnNwqyp2ScZA8hL+5F
peorobZN7uASDGVwBkJG+whMqfy2R1Lg+GGQXNeUokClONaeQw6UvuZv+M7gVitM0+W81hLPtBt0
k99TD8Z/QL01kjfkF5s2ukTaeFBBrbWTonrXXNa+duGayW3E4D+3xV3Z+6Hy/qeeiJlJWn8eJOZ5
aUMFzdfqQz3Dx3ffhjmxsmQMhusMoVGuZQk36UpSzcSPymMH1IFCVIanUMT6oTKD+wnge97mcl5T
qgQzkNjCYSrT5ZLFYkXe6QA5/ORFCpqyhke6t2uiy6oesvHkv2+QaNBWLwiKmL5nkv7gV2aLwl9E
anuqrSGq+RrOGoSG2z3RCj0F4e+k1i3gUTa42/M3ybBHf+T1WZ1bhZWlaGVQopYAEH1wxZREasze
VJz3VVrBcIJMgEjlt7azOP81gLr9mLBFz50TeMf4RYCKzRTn2xBV+EBdEBAP0bOMQ2/+yzsDt3O4
9MjkVIlIiaWHHSbBI6qd8kQUWoacKUG5WLU7Gg3sDiRRZMDgA/7zQhQ36jxcKgwCjwPLDm/qnw1s
gsVAAdl0vB9ZbzOpm/ZehDyFZ7EVsjsehIvXUtJd+cC4VRvuLZ+fQavLFyYhDth42LgFJU/bXEnN
8JUfG6RrZEaNchCdd0itt/Cu2bZpGoYS0XaknkryJb10mCULo5B/mBoHTUJL/RSTMEblgpftVkjJ
ty5Ah/aEN2PWFCjMGkNyOrDY0YABBvU07XrGSZ5Wyj5yQjp3KTMCkLmTX2zVsQEhbDLM8qylVtd+
r0jXNKIL9Lp+dfZX1ayFXzH4jUj4YvuvMb2AqaJJKjRlx942s8uoAqlQMa32caMsQTbmRGA2yemy
xWlsZWBEOqMoM1v11juiMFim/NWzNzPavyK0YTSrmUWMxUqBfElW+Wjs/P8ziMjbMXapw+JMph/d
KejHd1tuGIg3w9pdDANYSR5q3LjsXAnpDHxbiKMREBdzEiwDAsnMJE1z+FgzA1lenn7i6kmiCXJ3
yU4gX2C/Mc7VnErbEU37QZmQ0Kh9D9PMl0rZUV5z2glBosgSlILKdLNrJiO/gmuBH4EN8lCa1gsD
THvdGdNT7jaIyDlrNyQKBPgkJ6qNsZpsVwYj1vLFbZsNcYQiXmj+sbQoqgMpghLM866iRGCTBm0I
vcxd58xf7ihVuOwca61M+JzOx1KbsmmISfef3uwy7d4SgTQl8dKWJoWt0f6YNnIopRK0CpVl0KWQ
4g+60U5E24JCgZOizNuRZb+LLerx8T8Olg0OE4cf71lN4lXBb2QwHwZUYB/IyggY7GT9kDR08gOs
ghjhowfk00b8YwRkqnKMT1dbxbgnHvd8qIZ9H1o343JiNu8hoiKumoTh7tZCAiXC4vqQddaT2Viw
Afa9LXL4MMh1XNtaOA/pXfCRQHEfT9Zna3hsbI6itIFya1d7K4CzYKqbR32nX7q/Lv3xdcxbla3K
a6zvqQ6uxJRmpqWNOANuquDyL+ZT9PCcIucp/2ztFBvNcEqqMiF19aL1lgKp3MUyQa2NcvURl1kz
0nNPyYQKpIMBJhDgeLnKizcODWveDNsjBrAI7OaswqU4ZyUN1hEmU5ANWpxDeiR+BIS6ldKMBj1s
vhmH/+qRImkYjq4OslmImD1y6nOZ7RUlII+DVOz5Vzo2h/W29RwFqViZY+WKERT5lCji5yDxK3Uo
97w+g/acRKLn6izeUH5PisoD6FO6N4ac0gzChDP31wCA9o5Vmg7Xf8c6o2BahfRuxFql+VWOMstP
VobgTHaIS8bAIvn2PNxkX3a98ePAyC+fKIGX9RyiyhroZYIqn6tviZNMt1x/LCU3AC1s9DF0gBFU
521Lrlu8DMeHB4wPUt2NE7Yw4/fV+yVmVUT3tZiiXEd10oN04iTq/P7KBfaAjdpJsfe49yeaR0MN
HEUFqrxfM18jdg87OWkRsBs0chBqOpYQCFb3PGw7mX7J1pue4DkkFkbwm5zQ1M+aclT1ufE8An2Q
NmIl7JlIhpfhUhVIpg0gdlWW4d6mOVcyjAmkxHgVUeAkVA7G7LBb2Q2qlEAEY0xbGJp5MyO1xi28
uOUAJyLYorEdPyxI2vjnE4GVmx9rUFeYVC48SAsElkc+QZdQRkZMbH9YeiyUdarJbtRiWGDph6HY
GL6QtEGOGocAhjrBR6qMtRCwU7ze2klIPp14w6kEZiT2bDLnBMSs79PpwcFzpHghlB1BCpz2FE87
NwNwtZfFNfhIMQTOZbW8lmLl73IWe9VHHq4hxm2OAxz6we97XqcqQ0Aow36KMXeumu+yRwZGidZe
H96mRnjRrj5ptt7TK0OQyDvneFvn1P/UkL2XCy28/KeqgmJmsXwdybStlkGpppHy2tocp27W3Y18
Gj+0RESkd5otB3h87VsvGxtNP+cNILk0E+cSjdu/jcm/UPXZZ6VeIpaSFTPMJWuNTezdQebH58nT
DuzCoI9Sg6saIilFxYWJOQNXLDFEVmOpGQvLGmdTKeUI8665w77PiapxRgX8GO1LN/uusfHtxiMy
X/cwHd/GXWmGuvQWAJFLG4cU9HnoDVnncRxuHiYj4ZrAG+fhznu0MSlWVhTKuMRc4D825MUiOCfT
HSEWFeGJKzURb0HjzChCFhgcZnovMZeEFIbFZrIo/l91Jb6QyrRK7JqIhlxXQARcLSKzKa1DPuuq
KnnawfeHvl3k+PntzXGrC+11clQ8woKfvhPm0PeZzzrUzb3xkIT/O/hde7l/auGIUiVoT8fuc74t
aOZaEqv5msnykmxgc26R7stj2d8yZhN5OxWrNUfwz8HcHSwv4b9eLCpmLi43o5X3X3p9bxXwA8Bo
NSSJCuIGtVxzdn7v8dwn9yWdh76+OccJElSQY8QPaMm3n8L0Ot+OxRVPNm6w7gG1z/f+u4BFtbW3
q2C979IBZfTPwqO+VnfW4f4KfH2Hj30+NuR/Uw5I6KjHtCFIFDxsdPnBGO7ERPxM1l+RmU0O4x1Y
gCLLQK/JhVJm4KeLKm3RuIixvv+6ohjOKQiqhMsDIVdrpjqX+nugGeFWEIF4NkjU5bBcVXpva/8G
TZ8cbrPaqnvTgEgBHay67tmOZtdaUqXD/jXqP4lzInsmLKR55H0N+XttITyVsCSQXtmzTj1jj31r
LDdL8NKDJiRmTo+uSha/yS4vJNhsrFFmncuEMGHIJCJVIL1pdTfcCHZtzLNLqcFbLIGzfF5PValz
b6XR22o8d9OBzTuLonfizbQ7mWaXkZU+iSFZ6DhHt6jEQn+EG+7+g4ghp7C9kjZog7tXPmQDX9vy
RkaIONg0rIIWXYH3tqTfW+0IlpmXu0V4u+u7MendNn3ZbtB4zu5eSQIEsu7tSVrBhPjIxL5m1iAj
kpX0pv09ltwbgXpki0f82haLCAPEdMh7ggIXkeMQx3WutZEhncqe5+G6XDuLcQYl7rKXsgFAaaSX
nq/jX0EG1kbQRljogb49QQqXE9m6S+REAwvK1L5BRasSWvHNJ+EhJarVT9tFQd5ml9OvVs/TIcWY
LDgn02fpaPLbPtEkswJ3WryrA+2pQAH3tg7nEhKT6K6HGLltB12VcBSo9tWgp+dITm/EF+/FnA+K
REaMpMN2C/CE5EFy0D7ZGko5LudIz18RU3BMmj0UM11Pm2ZXCKNtPujqEFgxax+8PgsIPHDJ+yNR
uknSlSzrl1ehPqDKwpR+VbNdjMjrfEtAgkTn0xETecvZePvje8SOj10gWtj3G1Kn9gALyldhMXZD
H+oP/AlipcyNL3wRH9OYpA3UG3brBEkNP7zhziZc9RUj/SqRbkgcfoGY9st16TQRgO2wpRobmcTs
dOD5L8m1O7MsYGkUrL4jRSYmPTIf/scpLpw4nS2KtPbcY2aPeiwGnbGQacVB1b74NtIt7zfT66nl
GkXj80H+1/SYlZZwD5C1w4AbbEW/kYNr7EKXyn1Hio9TsCcWVkd+NxCLq6E9gP/XBkbVNodrPBRJ
NMQ3zk0vqfkRGB7aEfTYV4pBeV4Vi/UTTPfpnK9XQPmeMc5nYr4VnYxkZF6b8e1cAuGdoUQeE/Nd
33CSfRLu9dxxndf5Ltl2ViDcekDpXiRnKF8iKOJTyINdUDU81Zxtir44+CgE9qrpP1CcuDRpEvwN
uMoHkRQZNUnA8sjU+G1jwfXRVXSnD6mkgczGYvvGD4+a+AUGc+Y2/hrx2+HlyvCM1hMo5N7firj7
LwjpVSCs29ExQUCZJKLd0ybLsLIiX6X8dlnF0tfWz1pbEJRKQS5oeuoFRrFW4J/sHcZjrcGW6yGw
AxVxbxgtmoSPbitGjejkLOnLHb+IPbOJejahaxKxHdljZXTSyFI6rS9L2dWmxRbbkep3uMZN7f4J
v3et2D9/KsEFr+HtD6FvWwtdINP3X6r+o8Q0M+SfA5yNxPsfr8Ew8JwqWkjmcKVwiP12S0fFymPl
4sOVScCaLu0tilWSeCdUI8WwuOK3xMlmMKCSUD3FTlXseIRq8vfgL5ry5gLxqyE8V4plPny//9lS
5mLPz3ESj/7bRwg9xE9Ljln1ZqowzFGumx4deHSykcFIF2nDcxSNqWejggy02KCrLmVL/n83X359
HQz5OB+yHZNnR4IhMAnHuUNYdpFxMkP9QGooP/Dxdx71o+xH6pr0GhP+sDUf4ret6nP2cahH4U6w
/TWPOCvJFsOrXyCIq6lEmKvQWLGwg9Rf9j3I78tgTCU3tl13I4dmMTKA+7AAdK9Si7vNcMin/OJo
+vJ9MYthkmYHgS9CBbjy2cb+Ouqwovqod6mZaCqVPUp5g3fs7Ia6klmwxm7YGmBT9tGtB6yvKxHk
tV4M9zx8xN1nuo0/5OP6xBwMCjuQenIx/pd9Qaw4IhCaczhzAX2RfqA6XgcPHTsQccJ9S0rj2OR5
pevZZRWi+ZVd4uDeSY+BUYIvJ4dNpw+uEjIyRmpu1q1bS8h/Pk4bVmxmV+RWwFnhSkqxxrKR/2AX
/U52gnCJdaUw3PdqOI07i7AWYLQFChHbcqsDhFS1MiXiV+HA6Qj+9u1807dU3G5CV9K0xiG6biF4
7uARsWYDIZlO3zq6K0Hp8pXoTLggdxIAJXGXzI1c9REcNAz7QnHjVe5DWfSeEdxQuaaYt36bk9uv
liZAEZv+pYlDSkJ23dmP3NSdgq8x5ZTpyXPNHPTQneGfDt1Qx7YrtsX00t9Ico072qAD45x8W3gT
h9u/jOliu1ziFXT8cq3RnVGKuC25BpjgbepPPWZP0ycNWYGuvHXzISn9o3H8hLrqmKQ7hFlV6idn
84THZ6GrLrKEl2beTAqmTTztl/gQU7wN2Pnfm8zEdAz1aHrVjVnuc+4XEAVapj7dXF6PJhM/knq5
yS+CAO6qW/gUvm9uEKEQ1FO+VqwBz38ZncFN3X1PmGNjwMOR+BgRlvSTxyZ1whkyokg/db3VevBq
D+JMxdSs9gBmVIWhnlWt6Tu3wlNdNRZcPlcv1MMXN85lFYe1/jXjlZf/MsUrX8bUdvWX2bemNBtq
7ONZFFxT8UoahlBmkI7NGRNDikbyQ59oup9TEx+NPBjr4VBHRAyw5torfvCa/8C+wfU+zyDiIcwm
sykaBPKlZ+KMtgQDZ6adgSvKIt+hlaGOqpkZYNuvdSKeEb1TRo1Z3GFme2nqkkwf4Wj3Iki/0x/X
T/f2VWolftjs6pqII7Nhffggzsf7XjfZB5Q47n/1NevNRNxPyafzW3ttome41xdgesDnyI4CEwLY
Mv1hswgA47TQvQZ2q4EFGDW9qI7HHLgtLxhHLCJIVTTf+Wq/ChEkCZ3/kuNYUhimGpBTKegAQ3du
EK803qKteLatrkHi3IHcWPvpgxEzTqRJCdogC6SXwax1YacDDjtACFibJL0lyTXWc5qwX2w+qs+E
X/ZUFSrUREc2N6tLhz1KYOrhEmHaefJ0Dv0UqxF9a9dtRaGDw3CTmlo9yupgzX/ZKE/oZpmTq2Tf
xNfI/8+YUWiqk1+vp0ZayrkpPbVkfOyow8fnwwRccpPDS2B60njlRX7jsAzS/lryuKxFweTdrqw5
wa+rQQ0Oe3o89xNPuz9NLxO6Tw+JuEcK7FC2EBD32S7ULpRTh1QRTkT1HfpI76eBNxSeftTlx+Hm
hvO55nhlw26lNeBQmbk45MlXLhcqKJyxTrrjeQMj2ZN1ZWHAg+9gJ/COaxvdH/3I+zu0nYtS0F5L
grd9OHLcrLqBsEApnqtR9wEp+cxr1XlaSV2zkwsUF8088KRHAaeYSlbKUtGNPce5o1FpPAbbex/e
8CWA0E+7k6BrrhJQmbhOmykd/Yi91SWDpVjfB/trBFAbA6fxXjNdknKwHPsSQYTI8UL4pEzzXcEs
jdaTuNVWRoFT3Etg0UZ99RTlGkN4Y69ci4CjVE/ixH9HojqadwvIvLx2bUgLLlm+3CdKjC38Cq2U
O5UasVA+ch4Gp/Ok6XvVACosa/A5zw0odOOt3jLCgE6xjAtcHrCznwyS1RYva9hbqZyM4qE0hHAb
pIpSp5xbdMwGc9NfFoaj2RNCmwXVgf1uI2JazDrt5AEIzVIktQamRWW9BP7ELRRCjewOqG96JbmG
Km5eFKw1Ibv4K07Lmmvsyl2xUjFC3VY84ir3A1f7qpgcVlV6VMCzm7+j44hHS9yki/N51SjSlMTK
tlHMGiL67MYPHYdqr9pTfcgNltR7iVr37M9e80sMXufUS4NOydLXLt+g10sOpV8774zC5FXkGSHY
1tOsCUfRKWKmYQNbzMhLdg6PdfAHwM8fVe1HbnAUFLQ/KFaTns2Z+Ra3AOXfSZr/HPf99pFiQoxn
qOFOnvBh8yk7gJwWQymQMMks2nXTd0h2gMqyz0era4RxbGPgnnIXJtrvNHPQmhCwvDBujh2LIYjn
j2nRolBqTHN9xCSRFTlaUc5kOHZHs8GWNP8tKwx1gIInMeclJZzcmf7vhAvnPSwfekAvfF8zYkrf
alvkSfRPzbco2VeCTg32F3PTQk4f3IjrUSzq69qbpZU4CAh9c6THrOQE/cH8GXPplXbdTEhwccCu
9WAl/+pW0sGCdJgcMUBgFoaP61OjEQU2TlbroU2N8i7ebSFpqlYh/7YADSBvuKhyywpgmfo/QheJ
14mzVHN8bsqtboyQn36Hc2whesVvlqOrU0IF9XmRbaYjzHT2xzgjeJHjzkiWuhgFbyJYYihXxQXl
QzFCgFgWB/0x6yJT+HBua8LVsEWyWyyufzhSjVPD2gTHQFvAuYL4za+uRmem0cWZpUEI6iJjdN87
HvfYhcHXroLacgy0z6LsqI+TBDjmErS+/+Qzgo/ro+PSSt4BCqBKEEAW89LNCXHrD17WHaeJzNnB
8xD/f7Iou9BqmAcUJkPAo0OU/qfqY3uEkY6UqJ4JOozw0Ez7Xj6yH69UJk6GTj1xAzbDBNBQAga+
ygarIEnLLJDO5JIG7BijaqiNZwmhZeLKGUnJaA1J5Pa4A7j1zaM1qGdWdEj63YKIpdbfF4E0WSfI
2QV7sOQYoavUMRBhnAwcIBTFZJohciUbJagXxCqyURWIVLS2shLXmzzamliKvmSYHQgWcntYcsUA
8AkOFGCZo5aC4q0ul6TX+RSzYh9zwKX2VGRqSV+kYMrrPRgUVJPwPg+qELjcsZL5DTlw/vNW8hus
rePlLnFzPM8NbVHhpfKPWHRtPAtrb9B/nsOtDoF1D8Qq+SJ4sVWNbl/6e56gshoYz4QDXHjpA4O4
4uajcXYXcITOVwwkGkYUSX5uQwkWvHux72geXwciu+HaJDQQV0RyJA8GpRMQdrHXOe8IeiyMGmdY
t63BQ008yZ2/xGZEy86NJOJJcLTzvs1jTkOEACr7kmUjFs18I55gNKfYL+dC7WBIlbWccP9cujsD
Oo6sWjjHSmOBI332B/12asU06oMzf8Seerp1AFMGnmf+CLD0dEW8gXxaAeA67WugXcR4CAgxPUp5
VaAcaCc9rJgXpMk4TVFZ9MbF+64STy+wQ/NOVT2A1dKwDlyk/ssA2Vsp+6OxI+QUuYr1jhPVKmBy
wbn0xuGLZ5nKlAos52PutPDbuL0C1VC5c8aIjR0U6/TIb+MXF/vyYG8FGwtlICxBu8DTGPToSTzA
P29NKDy53OeLv2UYCf9CrfeKP19WfsaLPHxP1I8DqRJ0aMvgl6Ct5HsEj7q0mVUWfGXghcMEb24T
fyYZAo8aaeJymDDsrjH3rlzlBy0guV1l1gJmqIAbdAVX3ZXRcESrY1Gfol+7wA/Hr7JUKPejBVDn
cb5iF9SwRKil+K3FduFuuBiI00PpzaGx2XSJsYEwvmouvXzUbcUJOgZ4A5nnBuhNHOBWwA36ety/
D/YvAy3Zv4r5bU3omgVz/XNFh3QbzNkimITHSzDLuquJfrpTMU3zhzCs18IiCQZnVH951c5GJuir
meLRzglfyxrXUVcgQZiSm6ikGDtpzWRaZAD4aREa+4BNcDd/aGXFqWygETIFGIOUnfm68yMcdgEY
+bdCRnpH3eG7087o3NnTSZYP6BOzAPOzUK3O4MyjNaGQxABftHf5FaYQCLJ15XjPwonC41r+HDkO
9FQLwl1aH6bNhB3xbllT+oTXTohNsMJsetWKYic9+XCasJz6FGETHobeBtPQYs3ES1a+OTTcnoSM
i21plpH8vcmXSShn0zGEbrP7xCaCladpK8h2ZimDlKI98f0lYQUw+2gnPWxKHKZqjYYEWF08uk7e
HmMpUsOAg8t2tRbSqTS/slQjB1EuQZUu7zdRDrCEMdepgSWYXQoUasE12HmXKRzfkQFDCTx2NRkQ
FVTqA9zo3icTDVmb8McTAVq4USBBZG5VjzYD8wvUquyFK8L4zJdIC47tX0wVGNm7fvQ0SR6so9ym
heRV7Rkwj4fOobq6Gf6nV1y2Nmxzg4UkdxNy0cU9CmBaPpmxUmfoKOC1vhu/MMVZA3UzYVx2deQj
GSeH+VRLO5w2/7jih1ILGCbv7n9Q9c6071AsZV3nVrFGDSXVHro9dms89L4uZqcViZ47JO9NeSE/
9inq4fOF6VtILvPg7kqfp9OeQ+2W+MsFJYGIxELs6nCXSO+invr555jPCEp90/CZKqh8jBPKsoyf
4H50hR7Jmo7psRDlF1tne3RpJZ8Ucf4euy3XM+Zc7kGB4JksWPCzK9to/zpKmycRJoPmbScqEx94
hXGtLadFZ057rvP3nk0V5m9FSTV+owAieBkWJqlx+gDjuaYlfKr27yifPrIo3MxCgZHeMslOiTce
D+DbdbHOMUR2KVw6PtuqJnNUgQW28h9S4Jtk8NE3A5fh/8LBH1LTYd1fklXft3B8xOx85yKq3vg8
lvVcEntp0hz34IsfOr1E2e20wrgygeFqXn7p7O2WQFQZjDmO9D/lxB4pQYiE1UQd7IJC9iFvRGe+
ZZHDk3XVNQ3WfKi3hu+myWuXrUrCIdgADq34XbBu3fWRpXZlM1eifeqJ/+DQKtvRBtMakyxlgpin
3YSpQwAi2Ebm8HBlbBTfGHzvv65WllMMfAPOADTesBDGfxMyNIamMVHvf4u+4hL4/1Iy6S/VImtm
Jq9Wrbr0zueegUQ+AtmBfwQoqDZ2E657gf9MhpY0Rk19+tuA6Ms0JcEc7c1+6CZ7hm0aQ5pcbD45
pyG1qqdobgrEyGVftj4LYGdvVGvCGNx6kxBtFOCooJM2+IbPvFMYKSA0VgDM/wDi1ZVJnx1wnuZb
BeobxgtK2h2XfARHkUqHIqX4LYHS9KPotUQe/efosXt1qErfdriJnuhi+/XEofxvuZbEqePgFe1t
S1yJm0lguf+xd20ElnKins8h6Nwd2AGO2gtnexDuHjj1D6/w08COIrLIaLgNC8i1y6XJt1lXL51E
WNGZw7aeMbM9unZh9/nkDgvCYUuhKorhbp/IrNDfgMNp45uFSMzo1oIk25xUv8VLMdkT77ChT5X2
VtYLP7qrjlduNr1IytsLpUW6DZOfjJvJCDSkVsYc6jhUaLXh8HG/7sQ8WrRxfY29MUheMeU3AQcD
+5hoaEw9VGmV78HSs96WyARt8AGZ3C+u+51ZIl5xFOGEsMqDiufmz9XNwBXteOeGsiZgllYVHwCA
/nlEEQqiT94qr64/AVo9NEwbl8Dcg5uYeLvyza3vMIqXliAztV/RBJ+3PaGYOCxprEKKVBdtJEHd
160054IUGSLodmrQb7i4WJ6bdS/U9CkuRHh44NoKJQfnz5QH+YqacIGxYfL2klsh+ARHZSmDDSLV
26oas7YHwl5DEImPHMNbJ6X79JBjU5R7iXvvDXBDyTze+rhxl9lXymTlqOqMo/CDkAdJmeZhvF4I
zFEFVplKdN86yZZoJlLmlmCNFvbyfZXnmI0PIvaA1QiOv+zLi3ZIZvcLk43+Z8sNlvdfCpsOfPlr
YMZHcwqYMThk+EP6zETlp8QbOU4ZIkXBPYcrB4cNHmdKcIvsmHI8CCbH3y/OD/00Px4I8ZNV6nXG
AsUaACtpgZQtie4Un119THYjTLyzt2MRk40tN3PBKd5mmQ25oK2O55Nc9jUy+MrMuuEURsi4Kde/
0+z9mpETlFQG9ODTvB8IrbdKixihpZYA9bBWTXx+u01ehzAE8qNHokIAyLMMAePt67W+pojntSA/
00P+VStpUWu6UEIDZdz1qXX3BHBFc4NoOCIh8Q53pELIHkxASg0t501vwiBcdcrFC8w++rJxDyfr
unoOhdIr6ckLd87EiDx5/WWWJmAJX5yW3pp2Oze2/WcoqFfNaXYfk+7spkCzeAv2bdE2U3G68EQa
TqFFXyBefsgVDx3VFPOmM62Ol8PxIqKbDvXwZrZ1Q+H6epRZ7S4lAfTVjb1myIK15uK/aBE0jQom
tzDTAJt7/UdUeA9ZNUkk536D/gq25OZm4tjegtjeZfhr492f7X7GIT6XohKMuAhgKk8/MxvWLPrG
0OQZr1EAA/uMUjtVqUxffHKfWEcUzwPn5ajSisixBqWP6t8gX1JEMJY344ti+9W8KKx8g59XadPZ
CYMOzlepu46TC2/3lpL9H2VuROrjuUTBa2ur3zwTB7fKF2dBY8wAvwTXSyI36jSaj0M8r0B+UUp5
lB/UNvqRw1Rb9Y079uOrKtKIukbNiO6fOCFCSrF9iYzQL0MJ92kmkLPJMencsFkXJz0hqa/XZMvH
Fuzr7Jtgf5YZ2TaPLZf7njlGUjgnb1/GzKmV+awKccGjz16P0DgNCc2XqkjUrdgbv63gKPrjuzGm
WPlMUOnI7ZdchH8mbN0Z4dfiY2oZLETgJv8cRfQN2E/Vg2ZnV8txOffLidS8Ej5BccU29O+YckwB
fcMtFdkcSjY+9HEqkswA6LM7l+3orGQW0p4q6wuyJSXHGRTcWp5nXtZZ6IcGMk7O+n2/iWMpyQTj
VHu70NEO5ADVmaivUuq/d7KgZrs13falH1MFUCGfSrls8f+VcL2eDPnSRHFcbLv08kQLwK26hIoB
iSZh0GPfyncmq0BYvLR9IOEpYJn3hc/pNXCe+bft5WjTC/H6xEx1AYVfUmntkwrgq5AIwXI7H1kA
hPVRhrzF++3nvPexj2qyoI94N9HiL8O6KF8cjgJBRTqJiaDzFi7/bJHgq4KSSDBmHUzZYGhjC3ky
H6pzzMOLEGUMjcU1IJsYtNJ9QOOLGofxeqx6Dd6DvwTaLTWTcfP8qDGbb3zeVCQzfcYQGdtoMKs2
MJy0jK/TrxBUQVBF+t1REKbRWLabkLwAC1BFwXbwPs8NJHQ21/NhMngZX1H2JJWHP9IGA1mmi0c9
NPKomj5f9YKpI1lwKSUydER+pbauc2T54NmMI9KxGJhu1UZPhIqMxEkZNy6/4tQvO8HSlCyO8ItH
HbmPAuJ5pqLZJpTXrdqwkRBRKUgwHUjfw7n/760oGycakrnmeRY21DvEcLTlCWZ8Zc/zbjCKd9sQ
NpbzIOgFgvqV+uCQiXAisjJCJQ+y6DcQ724TiK7/QsDQ7WC+g/bPo19UftJlRxPNriMnzM99DRB/
VrwUSxGQ4wuq9yuq27SMBWOmnOa7FMKjQ8etGhyWmtyvAQZaGthhoxv1qRQ8KcZD9GSjq99ya1QC
no9jWtFNIMdhnHC2tZh3OmeDPVFM9qDb5yonTz/o4NjppyYYdFHOJXooYIP5U5+GORAN0DodEthC
cXvKeFXNuykatIxHDDonY1vuVxZaUSXyclvkbdTBzaBDsEt8IRx6te7fEv161uLUNVqgL+RqTjzv
9UPjnYr+8ROoUha1JCJNRLbHakZmpIugJdAweexQ425dwCf88P/bKTCqd+mSHQWmOqtne3kCg39o
nRhLHvfC5TlhTpqv5N0m3POf+LE0ethS26Muer9TKV+o4y11F9RPTd5mYo6AOBTmeOeNPRadUesr
6dQ3axjBCgV+HtCXdAdmeHXBLWGUltv2Hn1/dM6b+zMNj0+0gg4AVYiAmscIh1q66MT627alDA8A
C+3Am6knbtk1TB9VhLPKKZV+/R1m017ZkL4Nw75MiI/cSjEguESDtNHSgLu8cyaU8QuNWHgRZrgH
xTzbDLGWFcTOBCM1paNtTxlobYWjAYiFukNSaGujypH/JDf+5ZawrGqbvYGjTetvQK1r3LxOPWUd
c5K9BpF3tLIs3Ajt0oNjc6lWNdcn5GaJKAOkLU9STvob5o3l8uXC2RCadc5kF67BYnKyrE1kumSx
nzBYUIWj3NLXX6mg9MSj+Q5HnugxfAyB39XvMWWHRXAL7ddAblF8QxULswfTPGpEAJBi9tN8b/R2
Gv6dGWivcOZr3nKfvakWqelxPbxyiVhu/ocnXpN/Jt9PbZmsrz81wffo7B5dpcOGu7xhE5UsXzLW
gYKepH2F08SEtaV79PefM0gN2EH4hngQ+VhlQrjzzKuMK7M2cra5gKT2aXEFDMryNPOwqnY/Y1dc
+MUuLxXC1rDibf4vYjQR/5MWN6WX7o5uS6cryx2JA1aYI6Gzvb3agECC9h325wp+Hp/5B/Eecr+n
TZnLxeFGyYhoCGKT3YrYllHaKOymD1tNb+lAxwUxNP95RugNGphXA7lDYF5aZoB2maX5eQbnifoa
EwPpzIDd3ZbVAD02KwmKO0f/eTMuDcaATCRgxOKPyNrwomGD45ryJ/Co8GzrYryBBz+YOkAIjjyj
nvaHbgqPFwRNqNnf0bXp3iaxAZCVqBOMkB+ESdtFYXk/xS4ctOUM59yzOw/35/Dp+W4zIrCbUCo7
3aGIcwxc7SYs/rMxuqKBLisEXzvgazrviPXthGux45F1UpIPOgY3Jjz84alg7EKOS/B08bhEVWDN
1t/0HFKp6i7sX+zqqQb7MUETciVLlcvCWBR4DG6w4bsWFF7RMKK1Xf88ku6vd/sYsyjtNpxtTv5k
G8sRds4BZWDMjTwayvThNl/mYodqJK2K/wQ+olRK3kFFW54V1CdrLoGfRoVhmnVXJddKiie0DC/a
wP/11IYWZAvTeH9ymOQINO/3twm4HcmgmknVfgnwUtSwuKUzmottZF+GuzRiwfb9PCkmDJmgHpmH
Btts+LYovd7wP1Q/T2uYky/zy7LPx9zvTVpXN8IrvBEDKG8uJcqNDiDGpsLzTplYZ99XLFHZ8hOC
u2x5rEJp0qO2qqvSWKYsgvG9jj3WRLvpwQ/vkCfg/KXHyRSkOyFQ3ZStp3DqYP4UDb64aHPtqpIr
lT6z6asccpZ45kcroYjeXTjp2tEAhtpObGsI77DwWuKnQgemLezlmXWwmsJiThJu+m4wYGtWUhF3
Mzlz1ipRPRWN/FGpOr4tKLDldcbKrR9By/R7tkmKTEkRxnt/fFJ4Y6crbFLCRzv59QxvqEf9N1zg
8Au+S1e1b/6RzLKOUAHSkqe333kVQBpR5Dp71/pbmdKxRmtBaEi21qqagcTzLGYfIZSH0KRpm1wy
wpOq18LRzxUB6fv6WkebUY0vLissnoGCjumvpuik5KgFq9LgUeRJlEkdNQMMQHHMYfNkjZNAEqrh
7vMVdVh8a7IxFDYmqKdCbARQEPlux6SP1kAC1MTXFnVrOCoWjyGR9I15/lNlrI/uP7hlT+iDi4OE
+kE1s42Z3dYqE1DHvIzBLiuKgv9xTpYyKaYIHEc0+dwA/qNRGVxpxnvFAN3LoBnUWcpBShF1ecZd
3wHAkoxGfkiX4AdXICGWiP0VYz+QsScJCPiJ5uuiKcUYn/FpZWF24HCu3UDvk6pP/DcwV+vaOxAw
qsL5FEN4u5+S6XKCeAjJ+H3qOaz5xvNZSW+ZUwuNNTovRKMFIq36hDTW5yENbrSmuTUkXhrRc96b
UK28pnetYRy8ParcpqxKYnIjCm4iU9i6820PG05PxUFQlnokBOziMlY0wQUFhN1wjF6rJO/liYze
2w7O1ZR9LcOjXVHPM8z62JdALswQVOkWHOL9Lv4r3V4SxJyjXgT5o3urH97gaPR0INBl+tOVYJUK
W25OoqA91IWM2eC+tQVqEGzFnDkAJvps3CITFB8W/0pY0414733ikwPHzN5gvkboGFfI7HTL/XA1
gfTPArQ7U8FaK0U9nkmq9F0PlOZ5cK948x0Lxb0Vp1uAe0R+DDvp/c3jAKaNiz5u2oQQ5a7V2Za0
e88f1uKp5KTXZ2srBnr0mB4U7nsUbS4a3WWKMOKOo4YFrF27EhyoHcip1ombvpfCfLkyRQ+SItoK
tfa6+Nty8ZnUv4xv2QoCvMhsR2gDsgDdk9xRVHeBwmIUSlS+B84iw39GcE5WeIwIt46Z29VDaPyq
8W+6pX0ZTW1BxNavQRY/68B42SI8BFS6orDFTCEkrZW4slJ+vDLtwAmEcn7R/2hwivUFAco0J7BG
IA/lfvJMtjRMHyMDl1jV9kheP/nc6hWZfNCQhnHJp/F50UbchtsXlK30oL/tUnwtjILRfXVFvihe
jc6fus8TK6fRkK7DMVH11PgKWTAgRrxbFKDrBbk1SwURzZoxrvRaAlrxM//qfrNMxEWey1Ymhgr/
QrOQddtaXe+w144zTsTJf24v0vB+LrDvv/EdoFSibfOtFH02861+Hh7U42QwJhmYUCWda17b0ZDf
DvQ3GXE4ktAu9U7CnKa0HujKh5Q15G4xiCUMBwtb1HYdyixUEp201yru9lXasJk6pI/8BK7AmsOs
lkaLT+Bt6Y96zhKWg79ohipYiNe7SpYE82lnhX5rGeq3bhFGa6JsolBOTX5zW1T0wd1zebuGveiP
Y9UlDkG3QNBOjVFB8f3B8YTFbtwBKVyN6Fkc1ET/YC4xPFysMGxwcPYfL5WZ8Cr9GQUjzs7ImgYF
Ecx9bP39S9tlww9OnGnBFg6C5Tk60lludTAZ1plvOAFSI/mB9tKuhDzIsdY0QzHRksi1UF95k7vB
iKw5Awc1qtk95mvUcDBmtN6PbFMsmX5bZ9dwUZUdHGTJt5b/pma+S3Zk4sU3DHiDB3yOb12OaiPn
8vwIPx7mQu+aMycrTtL+W+oaxRDCxYXDroDOkcjdTvh08IXUZgNticows2ZfYjc48rvR9SHviHQS
aABGft/D2cCrBzoJacS/eNXTDN8TYLPlnOv8HDQ9jfxbxdhMORvWfca2a+JP2vYXX2jD7tMmjyq8
oezy3RO+V/Mcpi8aElIGhMz7e31kZDsrycvN2Wrf0aZbA5/Cw3JUbAfZjXn83T8cuiTB5PEM0t37
DuINW0smM1Tj8l0jyNCYwSlcxc2nK9CtQyYCzyNOvyt3MBUO72gZ1/Minm3Dl3nF8j4nBMdKyhND
NfPzm2vYRj76vtvz23ys31S3kCoB/ttiGf1EUElk1iirZ6YFlyTbShmvNXSmPnYdikWLw+ATPlf9
PS7w95YkTcs3Dsg0hUBYsC+zmN1UJM6qeBCchYVZprd22yEidzVSxTzOEcrneQx5Wz6TNZpDDm2o
3d6y+Fhipg55JsAagzpRDhkq9SY+TMmREWJCmgORa3yqn1c9FwE2OpokeQaAz6rFiaBbQCgyy1ox
F0rlONyGCXz+pP611Vge/X4b4tCHA4mMtip55A1+HEKOcQaiDEu0K+Lr0v0jFPJF7b5iJkLF5ZXL
abENns9qXIolUfmb7JIVBE941KBwVholcNl2x8qWyYKyqTfONSPkqyvReDolnQ3MGhSipDoozmlu
0hDxwbJBnxjP4R9YUbWEvwGuLFBP7HqD0c6Wbguy5Qiqp09dtjZyi9BSH4bzhSgWmHZHTMY2esO5
qNR4vSOE1+9SuxywsTXZMu7v+GameRNy/PkvWIX+KmUtlb8htN5C77W+curFMugYc+2oZ+N4fkTi
bba41wipRdZtmACbQ54cmQXlRyb1V/09uJmf8/lnRKUtAWlx0Pj5lFBOOkOuVROelAU0Ssujr1Pl
Z8jYZGImIPJTAJ4E/jtoK6u8zi1fTERUG9ie2bU1wE8+NhZoujnE6t3h+yQU/EVeWyMv2uGjjwlD
l5w9bgv4iMr+Fzr8yS8ZSUf8cahgf9g16gPu8+dbTFzrFl/DF5JPGBD9MOCLyOurSJo/KvBPM0mx
7+S7Sl3kY0l9kvpt1uRrEEh19SG1ifcDqtOIwgZo5j5Zqg9+xrRVde95ov2vtNUHJ8Li2jTNIXC9
C3o34vl30qJaMO0Ck87mkTJPUFRMqzE30knC2GdyACfEO3qhMzAKWOaZS2NitBFwtXyhN+bULn1n
bMjQorwTa4QlG1PY/oJRayg3QORgGbdJ4NEv7NAzCkBWrpjIG/RZqwqKK2QNzHqoeL6BG+uJpU7+
pNSQhCYk8/ttQkMW6s6Of4IR1wIHLWCOVhbfWHngiSE0L2J1LzI2q4d6ca5b+6x3s3WyMLQHb6GB
fKSaU2t82hGarHdMP+MufJ5daOnj3tH1wfmu9bezig6Q3OcVzq2+1GHOrwsNv9G9M9sl2c5F5EBm
fw/lZ0JT72abceiBVpZr9ts5w2Q4jxZ6TP4UszDffFd3EMMX+iZhLv75eYfAjS/mzhFB2Daik6p1
yGW0kNQhVBIGoLd5fnXj0ZS9vDWn8nVEbvyWooo0HQo/R8oiFVh6Mh3oXAI7adkeNfeORRC8+WVT
m2peqkSJriY54FhHUBVah3zzwJM2zRGGnRgve3Hqfe0r8ECGgxO3EXJi8phRnc8CX7IldKbU5/f+
AzhgAIthrT4mO8hcsgVqbjqvkey3C+T8Dp5YixwmoArozNVZPH5G/0sBQh1B8Eknf8zCZzFh7ENm
Gf22Ysh8kqTBMhIMggiY7DtEliLVJFykSOaAx/Umulle++Yr0WWW0m5B950sxeLScnpKvk+NrdUu
IaHLctEXWTce/fRMcrG8oNcB4L79Icru4v4FElC/F/CJn6U24MbxD/F3gB4RtkgymvwAF72OfA5T
UHKshBegIIqGw+P8TmBxmwSUmBIC7vBLBXRJ2f9/lDw+6LU6+CrKUOqWhYfvlKbfYlJb5j2/B2ok
VshYM5u2zuk+/mx+PPeXpblvklKOlrCygfWoEcpb+eu8R17/PA2oWxnME1m3fM9vICvzbjW6gRnn
qxP4QJFUgI6dUVAI7UOh769Z9/TTMOJROSjghd2vq2D+v/yAS34KmnAQ8Uf/BcYVmSQcdaNq32Kl
g50W589B1/z39z28p6ESRxiR0kOdg+R6COTZ8DtHjvi0AdBSCCDUhql1eIYuSWpt0TKSvcbYtnix
VnqlPLfdFUpF2iXMDXdHxWG8JKi/4yez6NI0Yhz/7AO3f45aAjj7k1rhgp64uRafqJxEm9D7ealv
nSItUUJrEJRfEHwrdlTIK2I9f6zC9HIHMdAZbhllCyTdLVABIRmcXzUAWLiiCkC3KDYPlM2xizKK
sHGuHWfREiLTx6lyxxeBm3oQ9ExIROG9S4eqC3IQBjNJqk9WvisFWN5wxfdrl+K+psxTmGi3fpYk
b3CcrH4AsTCkCaT09WKwJKIu5wEV59e9b8uKfx9wG9zxCf6iUO6oW8KtzqZdNw7MXtpQ53v/C4yr
0pj6ODwbqadb3nWhG7gPn147GsAGFkzlUyQBiGz/C44xSkzb0LZVSIetqjZQ7nPXKRyYBqsLaBJ7
iqeVOtwletxhSbhLuxasI4+vu08y7EcSWGZipgEZdVHG8s4VnRVZ0WDw7yJ20yhPdx4uFSYm6uwb
sQJPOcaj/PY6vDJthxE2BW2VYlY2ugUBGjLnhibwXKFEV3dDlr1opP8Qf4wATFjLTS6hpOJsxOIU
Ii/THyrbupWePEa6k6UIKZ34rOKS4SPciNYlO+4qEixWudyF22cLrO3cZtkhEIgVRyN4g/pi5q/s
uyHorTXKc1T3xVjEutFNXazTqL/7Jdv1AoF05m0tAlMfwVwFb++Sl9Kg3gmuvtP5NVmtN8mFvVC3
URyklperPbMnr6wdz6mSyApm89zhCWpOh9Gw4pF5dJtFMcUsi8+NoZmf+uw152bxdbu+y9M0mH3b
pvX/oV8/x1wUcEivGih0F7Mk/p1GWnB/bm29CEGIy9045JlcgQZpaeQ0RjbRpjR2kBapbgfQP/+e
3noTMyRw0BmAPHQHJ3Ulhy/tV3/DjnNJ+jVY5R45l/h6YenejTWx5BHaMl2D2vcYIgC7FBaN67Pe
sSTATD/di1JQ+QNwH/1qepXQkAhh7PoynTmHI0cRqwO+aYH8xtD1Z45isntGa5Ed3bMmCsa9DGFZ
uCHYfWSA2JMB56GHS62CURIxb8Sk5e8bQ5+DPJNpFbzeXwTir3ZFsuogD7AcCCUPut7Fv+1t4c3V
l/MIdGVtJIAdywE1scFo1OWIsw+PqWGbfraH5/Pnjw4Y9x46BNbdZvVvk1UV6yhq9ixTlSF3w+yR
jUayjB3a+pr1taFSj+ig8LT1QUPG28qk9Xt+Q1cSmBJy9SNNXNrt8rkdf7iHbhqYtHPJ+qYXDHuA
1UhUVoq7yoxtv1R4kVxZJ5M89qvq0Juw3kI4TgV2W1iZaigTXLGGkNW1/gmjDoQuCIvByT5FC18F
FngMPxRjyNjrhTggi2DdCx97omkRWWeH9c0gI9hegMYDuBEkDLQ7HatiIO0dqcyNfQEgtN7DTLtb
jF9TMbRYbaaYQIEqw72yxq0RKj8Qpqj2HDMulRdOG3ZLNBzA1ss7aV0FhFocBm41U2L/fNRSGmLf
A4YmhMzq9dwm/BXqFR1hhEtkz1QfsT0cLA2RYgrfuXV87go7B2X2yZCvP19iKuRjHcD7cMGXPIBE
sMiJC6kGQIZAsIGOefWqc1ks30xz/CjyAqxyIw+LfvHXb4+E4eG0bPaMTwADxj27GEWWqZRU0FKR
nCt+2BYJxb4cPeqNOEHT2A6te4TD/5Le5R0WIs6uxO05uqBimis4VY8ShY9nnhIypqn52Ugj/dh3
X2Hnf8MMwualGxXyNuo4c9tR3a7bxMBUnChXvvI5BlNoQlmSIiEMyvCKrVNo9Bqx6L+w/EGh36pw
KVvKy8lLtqk+o7P3VIg3OmYhela1z1/w/zMHef+Dv0t1cJL3n3wToCaJJRXP7XPZj98SZw0s0n7U
3Rs81yLq6ADzLZyg5iLtM6aTOHwrl1nLcOEn/6LfsaJszr9O8mEjFthI8zT9w8TPrRkcnE3VOpYS
pB7PHC1+0gNX2AJ86CXL01NumuL2LVsg+Ot6qdeBYomVlouKP1vzKKOU/DD/n8p0tzMjQLOAB7e3
Qwy5Bh3qluXeZln25mgrV6inofx6v00WB1lK4S8C/QG6OA3QdSPYLA7IzqGP3mFh6Y6VjSuPdKkl
qMuqlHnkRFGybe/SPQv5P3pLRDqM4a+wZMTdnXPLtqx1HK3/1EKfZFhvAb0mDkxWpgiO88iuLhVL
11JhZnHEROlPxDRVi5icQX+3W4oZ2KzCXOG8EJr+Sh022YF5Ra8JxX2eKDXSlhlvBpsAFEAjzX5p
oUV1gx2TPmEcQb79y6CnKgCTFrEauk5pZj1P5E9GfMicRD2ukk2pnPwM5mgpuOZHfha53BspdSQN
O1UxVM1WY/6rvjMC67iTU92CeM/z8cyt0eAddw/VLHSSUiuao61CvmcMhZJFB1QcZiZzoQb4Do9L
24V4Yge31nvT/qD4D55EWOrqwHBvkBwb2pCIpo0POTyY4488Nb8Kcf/WVwueGyV5oC1J91yNCkHi
lgi/+jkZ/jr6Kj18RTMNr3yth4/4ng8GKEb1UQJSUMI6WCY0tAlMVTPdtY7jRyp1Dj8Vu8/9v9OW
GNzTuWLJvf4juqc+Jc63weRXyRh9S1Zepgk05h51sCdiMknwPPuVgC7kDvBYIvH69/264AgDyRSf
FFrGwl89UXBnfNB07eAisrVHttx4j8RTEe5+ERU67zT1XC+4Qd9dB/eMQkvWXWH8xc8MPmTvBeRy
vdpYywbwYH24ejPlqyQA1yh9odxyl4imRoQuFC+DWbeGf3TmOhxG+faADKIWFm3zUoq/yWnz9etq
LmaUXLfRAYv1WDKGamN7eVsslhdywDBspGIQuauTk3GW3tiaDf/3XoeI0ZqEdGVUo2rKBYz+nnvy
/xuXAf0x0Ehe01l2IBW7DgUHrb2B87w4hXiLzLPYjIP0v+vdQf0tw9EKePt9eINC6FPe9Z1dw31R
XngCEBe+n8yOKqbaiHDRsQ9B10Zcg+q/em1atnLDfuDFUZoNMzaX323xfVZ87pMbyGAV8i40iAO2
FkXHKJ3AOFfZHsJ9SAKwycRi+XDlTdSfsJaFNMz+Au++spBRzd7BFC/lNoJ8wXxEpLc487nIBxzg
Z6BS+v8XkRvUMa71v4o+EB4UshWG/JSEq3PlXKlrNkono7YIk8Tk+UfdJmFiiOKw6wZOLI2M/ebi
qE7y0BOgVzfmsGLt6No1C7wgLlym6TgrISy0161YCa91fRZy0XN1NRIQLpXJCrR78GBSHm2g5gNJ
8hwtVAgwjFNPMM0YwM8lv0JQOsWrGSU+IJLySmi898D4a37VRnUFCm77RnlMoX37nplF9v5qT2Ei
Yoib2c615begaAeFY9tLcizknQLfX85h75Ch2X5q4Wx22f7kMiN/qCvmKpP0tn8eva0XaIBEvwUt
RjmVyl22QbZXGNJDJPyGb69KirvhoqtaEVKrbf45eoburekc+KnY0tSRruKk1GKE1LQSe+0mOn+f
wT09dPH0EMX5f9BkB+syi2zY5J0TDs+pedwXx3osCI/8KirT2p83QE5J4NyEKeBNsmVfDgSKN4y7
X0WUbz0fV6Egq/GeDq2BbmO9ioMs+3f/UnUxCKRsNkIXlGUDIqQEpQy/GWyHmG8nso37/6ZZUM57
C6KYWZTrmtMO+cuS0NNDi0TV20cSbu2RhP80xNsLIRYqIV3uUFNEv5lRnGGWH7YhMzAm7X4Qo78D
YuFPxe/Bd/7VhBjrgMQtimPkldAkcb6e2EFAw6zatkMoZqWNdvinncwir7n0aqMVO9hIDaIHqywl
exoALIqRnNuNbNu2HQ7p7SxX1QU7qdKvST5eZodnkAD4g2pszewt79u3FBFa0ygObSLQVRX837rD
Slo+gdLqTlVdCKqoKwyrKmabR4z/nfRriopOu0hGgGCAOqoTP1rZPS66iG88c5QuKnPt2vvXTGfs
q/NLhDIAOHx86cokvgjrBG374WkWin/+AhF6kOWCMTwQLZtIgVd1nM48dPJnSyRfDyLEv+u5RHRU
NPLfheoqCrdvhFkVIgNRpVE96lSUQdNYnPE/UiwQd6wC5OXQ0xHC/fC5SYZK0H8OKF8+Pgg8PUKA
ecXF6pVJ+W8AW8/hUazcRxMYSBeSXU4w5YTKR4xcKBbRHXCIXwA/NsHIG0i4cHd7RlEKL8ZYvlCR
QSIaPf3lQv6nHDB41zNWp/B6jZmH0CF/1Ahaq7jp/C8z84/jr7AhTF7pEmw/9UlTvGo9ZuACAQr5
imt8LG3wABITG8BKq3hk0UD+9xuvURpxDztLgCPKda3MYn/d2SsGQRmSz/aMebTnU6owTdjyX7uK
oluulP8puic/TQjOXCsCsJ2WNZJTnxRDXTqW6CI+vW5s+2fhKuMjITn0rU9fWNQ5tRTCTHUH2ZGx
5HAMSKWlQQYJH2xz1Y7mZPFmg2S00pm8JZMoDqFOjACKrNT8Zi2/muQwUg0tCtO5KP4k67Bxi0ik
LrK1chfrxk0n7Bl9jKklt0hrjVC3xjHIGoW9y4FYt3vU36R30nRdqkVEMUh0luqMyWzq314nHPFQ
NNJ7+9QQMcZ0Zg1fzMV4344SsZnbg6b9SU57Lwt2ccaHGc0dCNRxU4SIKPQMRC4y7yPPZ+9/uxoi
4klH4S+xA629yiiUtFtBsONK0kJm0g/P0iDG4mQETx8/XBGmDySJsltkwOdYRqKwGrF4V8sdxr9I
1ulffyjHJ6EQqo6JZ8pF+PiiCUzwHiaG7knTpyT4me5tv24gzbdLnBP5+WLE7XQmEem+X9QoFjF+
oPrmf8PP6FwZYkWbVX6hcFpkS5BUP/dIQqhMKfX/mN/pUbmJowoLqY58NOgsaL/wFgDyhwcN5Lj4
WANfB/GXuEcrNxz2EBGmgoxaOr1LGX3YLKQiPF5GY9ZoV+uXHbblrUOJII2Oz74InIkOSNh6VDvq
IJJH7Q7a0yjVlD+ADjyA998iFP0YE0xcmu/txjYGJW1/cTfzUDMRzbfBhnuUwX/sv1nWpn66Ov1+
L3fWNUDu5QBZgKB+om+KCMGboifglVqXYQ+z9CpWcqRlvKqADs55qBhALyo+Htx8UMUDa029M+ok
RoJWMSDdjPCqn9b4/GscHWtCtZ89njb+ZWqeEvamMsTy3OjJs+v/R932z4be9RCLupWA9HpFbxT5
wds9wy7NOMNh5t/ODzl5pIGkumtoEvPNLO56S0WWBu37oiY+4K2RlokenEtY9i3OMI6bGWdarHFh
A/kr5YHnR78Am59JwGpvIglRUhbsW58CyZHRoZ5GGpZUO52fq2Wx3rf4CWegVxfeubyoLXDzS+o8
o68oszaifXBIrVkZZ+dD6ANPNB97JRpqdtTWNmR+By1uHs8v8SWT/+OGHnXmTKuO+11O4fg2Xg1t
foNCQcDR0PT5KdE1seNKmbQ51JzCCkHdS2CIHuwLjPuGOI3ZkY/Y5uG6QwEDb42QJzI3gKbofhe+
7CLqaodzKYMzmanBbHsS6mEGSM593R9D5CI0BlvuqNlMjflz1bUOpfsNHllsXkFPOxzR1d2Xkn6p
gsWChyrrPBTPu1HKn01El/ROMH2iAnSKuoIGvMNhHNJCB4TgRPi5X3whK0OLqddl5AW5/g3npo/B
+HCpgkgzb1kn8nnpCb+ZSgPNLKwGdWyTZH0ReMzUu0Jlslq6+ha4NNzgdDWercJI7Ss9WmNUS36k
XcF62S3Nhh2xT2k+t7G9yazrsk2zO/iNriP1YBr6Sfc0cTzCS7I7hVkrlmkC1vuVjbBYuEjIYnLe
XrDJEb6lLe6QLImuBbO0wfChxqX9nM0UBIjEwvKTXbkddE1VrYlLINHKw8paBfkJp2a7cPS5O2wO
VcpxFP+rBG2qM1sLY+OgSRF/2Vz9KbsB7vzJxYXybBf9kD3d2d0XPEURQ/n1BFEebfdptF80Go41
4/c10FUE/4iKO19hydxgSVAitFvQN4Wk//0ldTMjoIuswsYQhUX7gy+Brfat2NoaoX5lIsqbC8Rp
WUt2ulzlaY0gcMzJOJJxzM/m3zsQTQjrxPGPgqE+Fk3W8cxIwqw1PinxtKa51CaaudGOiimp0R5U
LSb32B/WqJ+l6Q72DFw4RheHfXNg7R5ObvNjAYY4xWkOt4aWOXCAAxcoOJLJHXDRDSVQE8snHP3z
A7xYuNcvnJbe0muEaLfXXv4x74ybpSbYGTeQMcY0GhGv4xJi6Aeo2NSWaGpifdZ/QiLdAiySvIee
GPfe0U1/UmEV3tQnheJpybraBtlMLThL6EwmLL+u3bMIDNqIwUKpCVkMBzGROETDWUS9/9phfaog
NcIfyzDyuZi9+rMEui+PeQ7yZNFFR3aUWkNws3mXw6SyIopOSHE0Q6zIwc1M5XPVHJK5mOTsAx40
YsAWhkPpXQMotAANpbO9Wz304EWoAH5f753cOiyqT3jEbImIPr8ytRYNNtnB/NDtHukZUZGy6umy
WGUEDVGhpPRcx6QuDPo3aONS50EwcJ47UJxntCcOIKN1bWMMxm9VQ+m1pTthLw3JRG6PmhZjC4ig
/uSbkDFaNqKjGMJq6DvY4ojEnAa5ttfQRQwfCRs6rcNTgZhZ1f21EMjnmDdQ0Hk8fqzCTBW3qQlL
YhZAnnnAHvnBN6c7XFUoIBokg/3WKyv6q7AOfmWoHp8Z/4Y5PjX2M2OLdWlOgHA0U1U587IzqgUZ
Z3jvf0nlCxCKewY3ltUwOgOVLEqhgBiS9psIVcayJsSViaIvLswcGzb7pZNaN+rd7+X3mb9UTEAF
dWaz5UlhuB9AICA0nAjoCG9eSkwU3Jjte0k8elCW+KD3obpXqCZS5grJItdg+hc8YqQNjpL2phhX
4SjzPvnC0UPYbPhasVy5m5pMVmC2SlwtXUWOLYqV7hW4pyJcDfbhUaBzvn8rRzK2+tNBHdsN4UKw
SzYqfTI/oa4u1obYVe19zeuqbVatRU/OmmToF812j05OeF0UGna02oPdLIbaoljOs9b30r0Vcpid
8n+KhCKKXS4tCuSKzW5TpcNjVfFPg5rJWwB7lHRH3xmOYQGDcOa4yhgG/n3yc5VspJScmsCUrUJY
LyfpGQ5l3/1uSQDLcOda3zvzwIM40nmO7yJKxnAKSIIvUHzO0Qy6oIxHpWEm1JFXBUK3PWmA9/Q5
Tr9QpmFQQBmVJ0NhXDkovr8+fF0MYbFX+3+qJgJYt7hIXVa28oUwqz+otcW22ev7qe58Cb2az2Qa
d128CdlEFu1Nrmt9yyPMxE60v3dasnYOaa7/uMw2Q3RQkhis85VGn/LZjF88sYkN+pXJ/UhFn54t
yDLtjoo7x3v1zZ3lWUeEFqYgQF0YJgPObUjH40UMkblG3t02tNNXuuEcBUy4bnOSQ0c5t/pkuk+H
L0Vn7dqVesxw8BbNbZFRyh+2wALZcOBQOJkbr/bI/1A4MjSJfKavEMHiwM0MQ+CTSUMuk3MjR7NL
qTA1Qplkv4DbOpkzGOWfYB2FfARLxjalGsi3SsSRBfMs+RBL0R6O7gRfzjvozQDqHgk6cvTOg9tr
wgY0Krrt9lmhfQhe3ToM6R6dveqPquDxLLCqCJiDwu6vMuJ1+BqWKiYBbDhceyFsx2/PfEcWa1wB
3RAk1FgzCaW+MgCy1Hwgdkqgrv3DQxlZXiYTt1ElJmXVPv1ZtQ60/iYWBGlAItFkk63DfLJlwnx5
MCG46Thx8m2q4lV5HYstgMtoYxaNgeaJBIJ6VXgURbhJQgwq6teUIV/4gFSLiWnwLU7ihMDxsI0K
oeFaE6xukMM3t4fjrr+R5TEUK8nVNQcfpIk9N0z97ycCDFXpSKpzzEe39SLOPzInRz2GgsBQPJG8
IAoqmt2J0fM4o24pYimDDstw9rcneN+oRApeLiXJqovHcVVLI3qorkBLpr792tpZvbZhvMD+mrep
iB/MfbkmoRdcXS5JGB3zkTlMO8caKzZlsDcJPcaYGQVEwcq27uo7pfFAmDUJdm8YKgHCWWx/hf6R
UQzGGryTDW8/2l3+7ZwnEQtC6p/rWbyd1izAuaZMolvzQ6YjocKSEs5vjBuZUfQBHBeKJ/wGaKg3
Hm2j5yBcI5WHDiRK8vtnTG3MBnxn3FbsbgmUFLGwLFJCFbrZXCNErI87x+iKIJgdcI9HL06FHVRc
PN6GC/GpnJSCeJW9jz/UDGfMCMgvkON4sinVlVubU1kQxOXxxDyXKujdAfP49kEz9fqIvWqzJsQU
Esv1eIn+dVByc3LhHQmqiKVDnC5+Z0u+Ygz4RkpU0bkSyQUw0jGDasL7k+tXgApTGrDV1ofKnIlb
tZveWmLc/4yebnKiUIJm8IGYJovAarPyQJkNrbuEk3LrkiXzB/F6ws0C7rb7OYNnEeXEXm1u43yV
lo4UH1LIcXojcNV9MLJGFRUCVSSN++/Vlt+MKYw8fzASUG0zr1ANbc5BIlvlVPlodKhibxYrTH4M
j2THC7HpsX/Qoy3tpGhPWFS3P81qF1qigZlW0hCUKuo5g9A7Jeb3Aj+2+Rw9VDDZYnwgAQxk1kKe
rxw0Tallu3Bq2iU2OSS9gbKdcGcEwcVRc846OEUyyZEW9hiRUPzVraA6LRXi4TKcihxzWKYtgAKq
WufLbeVpMujk/XQ95I+ZL8xWrQOsVqI6QFSDmM9nSI3esYHwbdfuxKwARYwT0aIQ4GkifpCzeBfN
Ij9ZMtF5MQJSI38M1bw66JFZQxOc9RjVycoBOpqWTrNYOuqTsZErHPi1P0/mVrhVW+ofUeUuhlgM
ayV90CfavGz1eKsajetDE7ZhEE4YtG/n/YBvpjVnLhzB4nu9RUWtyNw4n407LkqhCY0oOk6AV8yb
tBkji+IZgk2NKuKWof/mWhyVRK9k0PD/zWlnGV3biTjGjhMi/smf0/HeYG7xtocO4tazDjhtzDUm
r+65WN03r6mlsZIM0MbkWgoyEeOxeFWwIBgwP3Kr/CFujVNFxwLgwvJaYnXp4Dmt53Dtjy4CL45A
6I30TAy2I5jSSHasn+Sft1KpG2pEJt18EamLEUotRON5n+ZkBuv4HWdFaFtYzsncupnIRHegbDrI
65eCVpW7gnDs54V/i8xild8xMqwVx90X745Wg9Wi6t7QZNoTXb6DQDlrUiBHtDUcM+zxU6tfJXMM
YXJdqI2JopDNYv7LwydWd2T5abGnLKmR2q6Y8UxlY7NvvLaCUan5gF+JOe8DhXfuJmeVmQv/IicH
yIfZ2AJOf84ErbsDubLtdt7flzNEIpOeLIg7mGwXLkoYiGY9Yt8yB0PnK26SjzfLZjUQAzQfajAH
NfltC+DhJNvliW3KCHnk9Z49REOQyERC2Bxu/6zCziqCXI3DEECdaN4rJVmJmiurb4oezCOhNNGP
W6hKg0AyIN+reZHaAN3SEMORH7hrwDcvndUywNWvvYPxvFWwiOS0S91iHZ8xh56Oc9DKYoeRfisj
VxC5VmEIGXGnL5a4zhLhPQzL/echnoomwR5/fhOzOmnz58PwyEQ+cAiVCz1O4qAH1FgSVgNpBK9s
2ZqDmiQZJdaw7lKLEyfiSy6b7531CKK7StR/VsRrYu4RgZTnavQbPB51vLYJZIWOCqlaGGYseX1t
X+cm1u02Hht4+cqvHTe74N6F3S3jMgTvClgP7B5X+ws0CQgcJClwh8LvnxkedTwI/fqzDT9ISIS+
vejdL2FzcMgrN/Q5zwFZBmtEtvHxC7gkf4pjHG1GnSacuFn2sWeDpYyNKNdX1QMu4zXsJZZbu8fQ
p+zsUnRCdWg2wnYq6jpopUy26Caq+4yUtTFldLnF00kgE859E894KXoB9T6PmtOhoc+hmdLN82gJ
HlYi9jNaFo2ThWebi6RNE6U1OJhwQ5OL5e30b95nOe9p5HZdbmdjYBtK2UtjOKs0SYGXVudIT38X
SvSM/dzZg8se8c/Jxl7snyWpcGYwbDmlbevOzzYX/8btTf9FN3NkSHaj5pzy3K81tgwvkWyPT0Zk
tqyoCDErlOE+BCKD6LgYfnsMP1ykphcb+lviEhpEijJ9EP86mtKxVtEimWlpKYim0mB0Bf9Mfn0/
WRAvSYz5gDNEdwDPuIXjEgUWfk96/wULFH2+VeDxcp7IgDZgan/ukG8K9r/Hm8ZnSozMUmAtVRNv
w+FbXzEc+d9RS9Z/ZMhAn9OzCjByCWhfCJFQ9Gf5PiX70kduzbfau45qUDAMWiFfMD8SMFPPt3xA
+rHnZfSVWsIDzGtkQCf/rFtvem1pUhQVV6EnHOlnpasijZ26gCExYrlckY/wGdhnSeUH4NaKt/2L
B1TaFwXbwF4Ae4qwBnJt2WxkQgk9bpma76amdTVidMjA4IDAg0KaHyR/o3hLwGnphiPvXB81/Uta
NtIji2uECGRwrMYjWjDZvlxJUdiahcaf5E9qTyLHhiHV5xvVgq8Rs/lCtuneLu49lCLOh9CI1cNS
C9HAvan3vxMMtrYWSub0ZMiO7iGfBnBKY4FENbvq2xHA4QzgVDjGiF8mr+l51AhP5O+aMVo+yOnp
KGSY+W05j2JvnG5fP/ht2W9SYsKcDXS/V/hjgKdL60vGfA63E3aEC/nTKJOR1lmm8hz47ip/R8jg
07frBbmOEBP3qyJ1MR/a7tpPYI0XIx51LhCDXbkA+ilL9ohxPuMFCWXcv0JFqGWV2l274+XwnwzE
veWwB/AUxHNDoqVCoHZxxfvMgjsIQN+DqOOXNPwj+YSS3+7lY95nFym62JTtIlAzNvZp1fNp0jPQ
kLqM1qHCY9Qy0e3tYZ8MLKPMDb96OzWdaCztgfjIpVjbhUrPgCRcPU+ONW8wnEP5GYnHNmP4uW9d
QnOQo9bDJUfMUWTnA+OBivekxO0D1eABOROYub0zzcZXng89J3bB+F8c//v1GmOS9FC1WSCdEFkT
YP/Rb7WpobmJXCWY0bOXgnGmv5jCAvLreos3d/N9bYrOhGTIUtHWPhfkONOcwNHJwoR0us+uM397
z/BNbu4VYCf6dmGU0yAiKpEoJhMMSOb5x9dJ3oSTEWidSvyV5c8tU6nOI1xUCxGfaACaYolyoiTv
PK31QwOa5Wj5ht0ZYeG/6Y1ekH/1HVhq/q/PNsaxRgiDr/xFQ6n6VzsAtyamfcY/CVrxHvEfGXun
7M9Yb95+04l4qPyO8aSNFHjzhwNHqo2B066mWQ6PSIuonwBNrGyBixJEm5v0L81eCkXAfqC2A+j8
fm3sLEpdJM3uMKSQvrD71+/+pd9a6K1RzDW0CHhL89pvKay6Fuimagq6bLC4LBupym8JYI4DYpnC
Bhs85Cv+pgAE2ibVsuAmB6493k4x1MDg5oIRwfw/eB+FXxbVWEHulgEgOAyLCW1XdVrq379zfiN4
vzqNDee38P9DNoYcsLOfWRasR39aitzpxo+NHuG6tGR8qVgaq0vnE18FbOA/53W8tT84dh2JvAh8
7WNcs3ccnOkgFChgjM67/xFEeNFXqmwamBn4aHiC2IDjXMbG+J020BCPOROoZZGULtgoF78k8Gfz
7RpahHilcJhy0GZ/iU6fnl3CGK4qgwSogiWs8ra2AJ5+DZApf6NgRQMlAAHI2bSbhizZmhpVVG+3
oesxai68B0x4Xmd/9JE4iyTlFby8nfEOAcswaeH5/YDWo4u1UfQICZQ7BPFiFnTi19DNA2i4pLET
lQmc2yseUobIb1YPqA32R14jOFo0roham0ONtcit3QyqA+o+nz+1AmFg6mZR01vJ9wRx72jLtqUv
6mScCE9i47iYc0hJoeoCCyk4p3upDQC9jiZ5+EWwS561bIGAuHWYkBxgcjarINPAq987ptUFj5Ht
gwmw6zcw/3hDojXxwrgBakP1JRL19mqq6Fe9G47tBEJ+u5Ru4jRLmrt5m25uYQyp9ZDcrB49KLz1
x/gYm43gGk3VGTFTNIXhoJGOY8yTxhLnEtMoh9UMqcbvdrduaNlTCU8RPBp/M3YE2KSPBUwI3RIs
FpFoj0Z7d7UKtv1DNFLapnbW2XXbsRClwaaoOPRdpIWdh1YkLMOegsUp6euvaNUVlMjZt06db7PE
LgMgQK5wuFoBjOCicy1+F0uyXME77Ha9SWQm47fqkqxtpk6Ag7lMFH5OCU0fZuwmxK0NzB89of5p
KlvcK5KJ/78oOgjKAl8kbjToVHzZu4dmHQ9NWzHTpvPWRAbYOakx1I2k41gV9ncnVPr0O4nkBCkI
XabKzk9zePGjNPMSYly733VJ2I5NJGL1Yxnnrlg/+23MDXIJ2MYAyBDlOm1mXqtzwkBRCZr443UG
ow998DqlAoUYIILz9TlgIbbg5DpyKBqp2xPh1+S7vvYKaRwJHex8DnqotLF+jb40xe2Idmcm5Fa9
SlZpr+m82slok4rTi/QlqrRIx+9mt2jx31fejtoJ6g13OO3E3Xamcm5+4xBIk4S4+GRrWOlfXDa1
cQRd8cOsaUkyh99NunHQg5Sht/HEEq005Ba+G2VD9bUBEZPNWAloVyseOeaqGCiZgNP3NZV6xctJ
lve5pfdIdxdXo0xMocHqfKd15Vvq5hXCQq7ovdoUl9FDoVMaO574lrc0HHSlucwEsQs4byvOVNMs
n0HcUKzYSRExnRoKzvTTFuiZP7BckbKkmdPlayZ5JO4E3pBti4Nmu6fJOH6978Pg8/kqHaf00Acv
wOP+TfbpQnKSlgg4+UIrMeqrddKHV4gTRDuJuvnk9QNkwv5ODO8XIUAhl55hFxKsIgIoXiXZgDYU
HOJNzmVjZTeNkdZ8ekTFoKDrUl0IpVSpqYTJ+ngN1blceL2TBWncsW7Ya31+MpK9RPqiop8uOL7n
mGhOGhDa+GDWqPrHz1LWxexRPm97DW31kClRL9iG60AWlyRYQqTp2anC9jJMPD1vRs4Y3MkPJzn3
WIY9aHKXpmFilisKSYD7drzh2KyaRLPTmaLyqLiUaFNoBLFcr/dQXYwYw0tSuuSt4IdpAwNrg5iu
X4RS9kIsab5vrhqHhqd/Sy85tpq+7ToHF18f3eaC0Mza4hWRA6zNhPJL9V5syI0W7Q2ZnFSYWIWz
TvbR/7KInI3FtBUmuT3LWghCzudqv3abDWBXF52XJFC/UxPW9+9GlwIiS+I1TiQgVlJn54VIQ0De
O0UtZz7Y5LX3A33HdPMLCfx5itiXB7cIxeEH4MWE0q3Clr8L7+yFXarDltQabgZxYLtOTj1bwAth
JnxNxfXt+5el68YDcXcA7wXTX2+R9T8FAR5JL4Yp/X2gLqUe3Rw9anFhOeUeQsEdLSz3ul1O/+LT
CJpk1EVJHzZpPDQCltc6qwOnqbARHkNNOEUbKsAcDc1V1RDZoh3W/F/tjcD4Xr4jf2EJCOSpbrRY
6nI2Sed8pg+r+R85lOHw96Q8I6sUSsuVdH/6XzN869vhviu5YMuC1ooRqmR99R8QtJUbHxFyQ1uJ
utBUCZCkpkWa6Ivqf+9e546husWSYjMGxcbexXpB8k+CgVoq5BfLtm0WmvL8XNZvlhJ/DuW0xICt
4yFipka7DUB9pmEgG4iJKu4dRH3AMjHAwXYrIE7BZ3fP9UMv91bYgF4cGXa4P4qoW+B9sewTotJo
6/x9jXadvG0RoQXPZEkMHOdsan/vN3BAMUJb9+xymx1nkvpE8hvza8DEbFGmcJmb8eyWWUZB/NC8
NcLD18YVM1KBySvuK4qMZ9Bo9SpCMZxBvDOPmx4k3zv9Zjp4U4hW+3Ln4XKRvtM2YJWefkJg9Sd4
QzY9rS8eMOuK820POxj+JR9qsgkM95K+pMAn9VoXraswGGKGYyB0oKieCKxn0DvmT1zgS2J1YD1j
Oj2JucRjR9E3lKP0npJZTVh46S7krquRmkaxGOpdlhNyJ30PKQQnueLlewX9D8KeFMxckRpYIwjz
B8udHRIll6wQo70BM/lL9ENopOvLybF0i3vBKFn/MKwYlunHqhLczUicd6d1D/GAuzIfuF4lm0WE
s9u0IYASp7dB/55PDMbRNwqs0WuJOLLbpIlAkim0a9372T3FZx55z5ka5gsLIcl7f/2o+j0E7YA/
LFo6FCOGcTmh4ln17Tckuajct9OPNIKQOGxqmMoyfQDQISAHkf2e4/6OLfxD2GUxfuL1qenNHvt9
htNZOKxdhgJr5sQigtoVAejHb1L4EADWkJQAgCAb1yYFGv5yvUA6IiWVUCMK0tynXFg4bYFWamtk
GgQ22VDFOQ8mQqwqzUboDBBVnu2uvmaheT+5Oab1FTMcQf1QyW9QMVWIVvieqsYTUZ7Gd3skURLj
s8lqUIt1ncli0Cg3fkDVvI3bZohp9nvp0uTGIcU4PSuOwr3QqVpcIPZAiLlc0PSkA5HYgmpDdHd6
mRkMtU0FDYoHgDiZEE3fkVic6kIavJ8oOFoHuTqZ0Hfehj+mx4x8MlmxPUije7Goog/BQRLGkHTt
8pxHgzppXEROCwC/3+AL6pyYLVLIR9sjizTAqkoJhG/QWGNVXE80NOXTVWGjARtWYSzPECvIo6TS
f0MhE5mAJ/phyiz9VzKoZAd1fqEcLgFFF5CcEZ5LQB7ZKxmCWbywSqdtU7Kplwnc4BkN1VBR00g9
ooU72jqP9jRezsxPd4gGHJnjwb17J99pPo9H8NTF4Ad2IRmE/tg+JHQYx4JhWPrahKmuE46guk1P
oO2Tr/VtvKuvvOKDh+se0/dh1ce71WdUbNteuRi2qnN0bNN/ZWfDhm+9sdHomo8Vxv8QzRl+VxCk
4GSO3CAjiqcg7R3IjGvbbj9G6AqAj8swbAZWqGVrkDDrMstSdQz1MfG4WDBYL51O/8aKAVSNmrhc
OM1Wh+YXML6JDvZxTW2NRTy65JEdeSVb/y/4cf/1ORiqdHWyaN6WqwuIw3HUAJBU6xE2TAJ1AH9j
zOFNXMdRGqmzuxYWwquvPFeQ2oBm/7w/nm/YZ6XqAGsQlWbPPuSjQ6/7AFncmssOBCarO1pLogYL
xw0siMqxCiiN7hiYYyVBaJgmZWHqBnT3qjgbtkwHgfi24Y6ziNnOgzTu/rxNeWM2cs9cIAJCxZz/
iWVxjrBDbFguWUv4hUc4eUpInr2HymJF4Jo3AC20eNRUgxQC8Pk3NXzIjj62TqH5BodMbPiJQ7PA
7wG28MhFk1walNWVLKSSiGTSnpxgSk+exx1awZQPxK8YEEN3Q+0pjuo4hKh9hPiGoXJMFCZ8lVp9
TFUCn5j9rGQUurTKtfiGajqENEXHeSwOYja2fpT+AHtaip90VNbC2NY6dn1JhIEEqQhKiJRzlo1A
nN1NtGQPK6D8DaZfWWW0ChNVOXD1DQagqSbsPrfllNHrbFACEJeK1qbMAW6EJ6hEOJEHBGvk0f7h
pBV3QpG+VW1zruApIpYH3thlf+0gDa5T3vDAC3l0eJRODjOCZVUxoM+gKAkyVCHSaWcGj3JAItFj
sQMI3Oy89zXm2EkV9tPGkiweFXI4IM249yEvw94KxaMxUcAWqXrXvEbPt/olWW0vTMLxOMHvCrOO
b20Eksv/UStqV1+XcbLrPnKCZnVJzW+aMgwZLd9LeASDgAkfnsBEm9S4IyK65+tTvzKLlWodQos4
O1c8eYXiel1iFN0p/02nRx0F6dxiyelpv7HiDinw7RCIj3IG6RK18StnaZLguLIt7iV3qcAdA3iD
Z/u+pDgyqwjCWpitA+TZ+vZp3iIb0T1+XOtxaMESzo4NzxfvABxL06dFbpwEJH1AisE4yDZEVqml
06HxnxJTliABbP7KqZx+PnT1hKI/AdaADHDPGyp9N+b1V5bRBRMF2zfus2ihead6+bjXu/nQv/lF
TIVNz/LTLhmM8OR4lKXy05tEGCRcxT9FzjPmT1lvF0C6VOC+xgLNDp34irJq6nXlZkwXAsZhv9yH
aFEFCPnGDWk5h6mfKMntfXc4BBe9UP9HdLm4cIQpIsY81zVIkLKk6S2TrVfc4TZpwCvg/EVRRlV/
Mefu8QmyauYyrBUFgUHsTETO+NvJMxSiuCt76nosEzom873vRgYDBmwf1j2w5YoycbG1EXQAWpqU
6WTW7yLhrRi9YAni0i9CfBW8gK59vcVh/4wjGG8GLda/jT8oYj4/PBECHuNklea4p80covd6euPP
KC4hFHuvTdeb7ciRyudXTeAnwIhvMnAsBo69rSTzYLPJVj56Wz6JdO0egsUSs5AAiS8mOdPHosvi
OSdvg573+8EhNDJ+ikPiGO8edohiXad9eb9n608am0a3D3u4dUQhfesMebPefNXXPi/VFmKoO0Ej
KMj8+RYHZChhU+rq1/7RYsKrqOUwDVAl78d0y6yD1yCkebCiE2BWuaC+dV7+Wqv/S5LDhbnx2sX7
KGaOdWIgZAE/9ugCVOgAWKVVcRrFWYmEFFW6wtU0/h8tlK6aUbc8XaMydUwEVejfJ5cOpsNO0Q6d
n9ErpiBFJdThNsAabnLliTaKXcldquPrVz+sg/CrJcdOaXIzSmFU2GJ2jFwshvOTi40EKX9PLYmk
f/zVsBLUJvZp8dMrK35Ph8dc/0X773BhqPANGJ1pfAF6ZaUZgTPeOcwInGPbP8jHcSiOJtBxSW6Z
KdAUN69ndIi6vw7jQ6vViLn4Azedl5gQqYdY6HLlCxhYokERrxmBcddE4of/2Ld9LNjvM83l3FSH
p2Fl3ccOcNE6FSaMTMGUE+MIwjOlC7bcIRtQw/urB0E/8dznzS+tqEOnd5Grb84VrO+QJlK5mI/r
SuHENNoRBDJ2fsV8q4tsHF4lBA+R3FdfACSp319Gn2B2ng0GwfxKoA1yudQB1Qz0sWrCL7I4vh1/
OBlbWZmG08vS0C5PttRE+X8OqImwdWtI0UG/at2LM6/yK35Sri9k/H9NyP3SvzfnDDkXXQ2b3bU8
AV1hv90wJSHI53qAXA+n04t/0mVsVS4EfPH0dhN5r+X2BIozP1iCk+o7iyrVvfZV7KRExEGHDaO+
xsJANitnhITd8dF93lzzT9h6/oK9YN+q+q65vVgk3WsW8PaZZQBiZ+pQO5cgO0TVTGy0RFu4GLMa
r2od6Ya7FAKx6PYnvksAVx1QKIJ92pz3YJmZY9u/+sk78aYfb+niDF+Y8Jp/GzX/9SMFIBbsUb1N
VCSJN70MhTb8705zKGOBJ8z6Xk3JGnJF9RpzOrn2TDhPHNfXA8+yHgb5e7vm5KOnKue++5pER+S0
pbIDpfIGDpzrSRvyNW7v8EzbHvDALb74pDerYNCXFFhzLaqxpQGnaItJjciAF0XS6MOXZR+NlivE
I3JgTxskeW4/DWZbaDJZOyNhgDQwRgB4L/AhUF0SpdT1OnB/pWGp6XjzpqYIcwWEd6uMoFR3CKz7
Z4p+1XPSNux8/iqKsAIlG4F+FyDNfBm12ma0nnAMrzm6wM8yXjbRVFZpXH3uP8Zb410nYrtVIdr5
cvm9Y0VA2DIiiCwXEphxDfcwRF3rXzEypiOGRHTrldM99bcvKLeOUBtKsY+bXNg05RYLJiXRWJot
qoX3UFul8GFGzoWkGnCQwNzlAwJp2ILx7AjSRtUhXaTY7n3e/vcOrJRR6topeQTw1bdJXGm28rNE
KWXj59Y1+XCUoZDcVPwWhP6pyfp1mUbpSZHCJ0I1bDyQASVuiuDAK7IPQjxZ4Ffyr9SctuHiZ1tS
eycmgGHnq/j0udE17lMmILPXzfxA8eeeE777DZDvlp+jgQbnYPrwZM6gBamxB4U5BcZmBlSjL0Wu
nj4Hbs70UeWpGabWJJmJlnLfAXPtZFIAF7AdO+k2yONXZgDjzYFVRQFiYU3O8pK89IHjuPtZO980
beWJe7zNmZea3UjkRIRRiMtHu7DBcTPuM7qoMdQWUFdOqgmybsRcTqBj5cXEYrqzEa7ucqM9TYC6
ravt/5BrRhrM7lxrUJJKl6dv3Gg8jbNl8b270ohh9HkpOUUWxiZaOEJrQLiOMTlcqyBmyWguU9jy
xjhG8CszMyOJuWLjhBi7gcwzBIz/FqXHb/ZQTX0n3NL14jbygy6NYkasEsagKI3zOdLhSP+aJhaS
r56L5c8syghxm9lw9Log7k2RO6EbFOdRGWO+IeetDBbAEN/ALGbxGm2ganQGmu/Dm0j/WLv1TRun
8F1nYTsrtUihVKI3CzIPO7iSdr+AHORxEFBZz0TO+DWrl29U0wyCcP5SLAg1RQavZIxeHq79f5jm
onAS56lZCMAcZKIz/wQlZOhEobjeaAXbU3tRqrMexqxBEnjLp/aFJJhxUZnIBatuo4eUvGw7RjVT
elLBCsrLaQN4ic5isDPl/TmwA/pV1fjGIrEom0pG8QaP/NxWHMpvslQ6WFRlhlzo9UDFysS0WfjS
Edhq9/iaiWcRD6KyyW95svJxXEUeN9I307dY6qKQpQdSjSc5pEozxePm9Yrs1CRj8yh4bkyKWKTF
hKh02oKkLao1AHJtf0lfwoUNVGaoa882qgH8O1wYPjduwIqfnzeXIYT4tgveseNtMjvKASQtDeTg
THhwLMV+rZjyk88oJSh2RDqkfe3uzaHc/Qa/G6QN0+g+UC5Es6Y4Urq1MxSDC2crJbQzI/2D5JPm
U4v0drIOt3ngifC1zUTWokGz9Sg44OTw8j2MmydIjQ+jXJJbLIWD0liqUjOSzs+LjFbqbHIfkow3
cgybC6G3GV/QA9Ns4C9jz3WRA7v82fnd1MOEZGlLcGnzBqoDI6gkT/WZiZJ9vWX1iIICxW10rQt+
ovdo2AXy4V1XLXjeUDhirY985Gz1XoN3bfPgDRHEmBgZR6dBlW+IRgIOC9uYJQcii5BQxzlMIsLg
yak+TX+a51YgX5OOdDjDIN08oZGz3HQZE67HuIiMfoAUm1mczOVwbKKjKATqfQ9PCn/nzQtYqRXU
t8XWzoi5wB5OYLO6/ajuIDNvwcCJLc1DmRY78d0pKfIDfQ1Ak5F+pgGg8FX5F/2kbQ78wN+Jl6tY
YdjylR593lngafWbF6G4PdKkN33bcQgISDFt05t5o5aFkto2+F2w7lStWjk3zcbOA4Jkc1brrEcD
whfxmwQ8cRSn5bgGXtOPNDUmmf0bY4MdfAb0yQ3kcgNYBcN9Cjen54fFbNS43ZhMJoOGOoPiVvYQ
urelBe97ILj+8KcSD6QpSpGudqZwahYbdxgmeGIYd3iBJ3boNfU+OzUZz4hpipN4fl4dkneuiF00
Yp0aKckfiS3wGFW/KJPP4ltuMDQD6KSNDANjIv1D6izOtBxIMcdIpiyN0j/KSS6FahsNlSfi905M
9SG9VGvSQOL5ekDLFNrOgiHNmyFvJV2kETvi5TFMzxmzNyinh8bxFOEMfClwFrcLFl4nuxOTA5Cw
maZAGCBdK2gFBsXt6sgILTWZFG8BAMMbDgqngpagfMB3EQFAE7cyBJ8WbShE8lQLp7jcBPL+copT
Tig7E/g0AQIrdQVYUoaWk3wZLO2m6p0NEQOzcsNE0hqW/ScOrqqzk9QIKW5W94DZ7y3FY64C6yUl
s+TfKMXYBlEKH7kxhyR4zub60PkEHq552vz+vVsQMBKepBQPzK5mRiU/u8eNI6LYfvaSw1K8e3Jb
KhaLRfO8awUyu7iVVBm0NtOMb6K29v8BV9c1Ho37SsZwCcH2fjDIvI8cTpEfdDvCOY+VkDH5YOAV
/Q+bwmn37C/MI6BAX4k/YneKCLmBcnjM/k7c3Hfr2GhUKt4WeZZ/tvUYL+tUUZEWDZXfUOnPlezr
tjQYd6ERWVq67e7L66hUURZG1ZPRpA8UbPtqjSQIw2OGJ1ewvnlkw6VCWgqrRroD2+2wld2hPOl9
8J4F+wxXU6OITIXzSceZvggrvbBN8JYI8XU9vIZD5q4AyHzkFd47Xltysto15nsroRwyWzeqJ6Jp
+Gf5bAQh6/1ENPjoVVb8DFGvXjeGrlSdn6ZZLuwvB6AU6K08pQ1ZDecAVsVPJgJBb2U+jaNNsbtP
rhisZi+34vB0MKMdFywVHeIHrvSTx0QPq3Jr9JhqEtcxzApoEaKRajCmggiGtxNtXmsnCusvXUO0
Iws0ff79GeSSETzeXvD4OVEBj2WP/aSa4N6ttBrNs3szrX4iTgYOilMUWR1dqC/mgBTUyFKF6Q+g
WUxTQ5tSNQswpj5pu2DgphKV/Xz+Jmfi/ORB+bn/vEpO5K/2A9iMQEPYe3kNjNssOekUmt+PzZzU
CrtwzthpSM+Psaym214ZALwF6oE7B5WhuKAUCMc49hR1h7f/ndQWCwzvQDpLb5R8wE9sgW9gkul9
Y3950B5LAdjaqXhmtJCcAocFTRp1r9OB83QKU/fecLV0XeOXDLp2JVswwwA6GhwVZMozbLYGdz2R
6JyHDPkibWQF1Hskhvmy8PLyiPiebXNm6u0w6UqKkwy5OOAUGM9t0ORFrpwj60R6n1S0BESnLPrY
h+5JyXBG9YbNd0ieY4ESvHxRsyZelGTm0d/sdF81DdUwwhY82wvSuR1e5tGitxschqQd0YBkIjrI
k9stKtQ1wV96de6zBT5iHvijNV3R4k7zfwPiMt0hSEBVvqfgynBCjuPE2GgLM5rogkO94s+EUnKN
aqH2wpfpNZLc9OJ7nPfgjgjPGyMMwHWb8BPporTqW8mWpLtmMSSYTxV11k6ipe4mcBoS8fSsMJjv
d0wbfjaZ3slMt0CQ0WKQ7smEZeKOdmqD/QQPBHUKmkRR9bKEgD/im2HwPBxEAtz8LQnnTU05Fz7u
Z1ZehqyM6gF9Va5meEHwPqei321OC2pRxNxqh+QILEy4/ZB6kl4XrQJ19X/CCMEEa7MWYmfKVJE6
MPePaGQhmQlsqGPLkGco7YPNxJEqbXf4HJ6bqSC6fyBKVfACys1Q0CRCGIrka8SkoBm6H3VP+fXI
MMHxjphOHe/eLuVOBrtgr+WMuYw46KihxFcV541jxXjJugfJwNBoYDjTKg8qWiyZL8oUTt/Kh27q
SgofX4sP1KgBsKPjc1V0WXYO94Q/OBpfyOuzfqNdzEbx3GwqVf2pw5uuISq1/RQ1x5tzogsgGCWd
5/seP4QYnioYQe13AxaV5+RcyKHyz1cUer3fEY8/ISPM8mSZjWtiYtsbILTl7TakZsnYWwQ0DncS
HUsXnCBMxQEJHpPCI1LzbZtslaJ8cj+Ym4/g0HHVxrGBEMwuY2Yi7ZiJ+AvzZaIIS7JzEwEqeVHW
JfXXpEZGe9zihDEbJtXuL4HQc3GfjPwbNGQM07EpodL/AMfpdZbFCYURrJg6oVceriqR1EDSpla8
IbA7/b8Wwhvr2KCW/w/wnSvAUJrsHnTP7dj56kdCxv1lgqcnvYQGkij9wfdJ+NAmkuYdL3luG7iz
pJtdL754dpAE9dyG3GP2r/rkkrsStKAQTni3ebrO4jc59SDvgloNoGevZUSMO5tMkIE2Yi55dnd8
DvnuXLeEj2SFLAJBTm2tnIxOBIopQ6VpdT+lv5a6R8PQX4m5qEbwsMsX3a5Orq20a+iDi5Lki/I0
f0W6ZIyhLVEKPlCT6BL0tjjA8ssgoBMxzFDLqUFG0PF6Xrvj6dBzPRg5/5eNJqiL1My8LXg2T+9b
sELgcpeYIMFO2KRGqIyzOLWoUmYkuzYZTJlsSX/GEEozCTmm3ZkFdr/zxzeqMkCgji2oTcxPexqP
r08DX44Z5Repc2NiTAPashC/Cz9QmxDtAytXijLLOsJl6n3u7QjvrNeKB+pk/y3OfheUmaLBin0i
M7sSIv+MsrhwdpO7Sgydahmtai6/wiyvs3rEOIfvKn22TtAvC7KfZZndhg7DUhPVzUhgCczuuoST
VZZyGKzE+JhGehOqyoiW9m1DSst7pqN5ClTpjzqGXgXA7p5B6tWTGVaDiD7vgDfVHezWgVH+kzsc
TMo711SpjFgEGScpWXyFVJHaU0p+c3+8qIQMQEDkOvlOtWrszkWWRSgSEpJ5Sy8NSdF/eEBE9XmD
Ws6D1bAYf0ncggzOVgYOsXrlZ2Uc6zJP0kdNIDOnKuXxQdRabALI3wQ2THa9cXAs+RqcTnvcJlRg
j9mJ890AYTZRqOx2wUKzOfGAteOU13PprLgahx5GKB6M6xkbIwOPPKTz4MLE28lYaGyTaOF+Y1jG
qNIT12eG8ZBbX1pOTAvdeYpmSii3gG6+JmrSLi6I1QoshvSC58bLXzhdmgp+hswGNPsf6jAuv9r1
vNUVjvyrYFzhSZmweWiNZ02o2NuxvB2IgcL5oHIxmoD/WDVARei1PBQjJJEg/eMEBvf8qR7lDCll
mPmhpKdqh1KiCmi2alGTBbqnLhtG6G4XzxFwmKzB8oTLu1lISacPZ4/f2RqR+uwGoe1cA1ml+Rxa
9fwmRV4R0Y7udA/Uy5T/rdpq2doxuW+PVJIUTQXLEbEY7R0UnJ0+wuRpFuxTa7WtzHTcYZG+7kO7
H0pfOwWgxzOY9DMvrzYDcMcBw8AZaxJUbV7/xcCx9+eum2DQkaNDV9tMRbnFHWPzd4jKkTx2pFG8
MVy2BqsOS+6J00sgNRWcrhrIt/IHarub+pp7OCqDlPMGuoDL1kpYRwjpG2eWwYgkLCdgof0UfH0P
mxtwW0SocOPwC0ib9vsZi8XV5txvMo9sRdjiYRnT8OaSdwmy0gwoXuTGOy4rbhyahO/tG6zGS7e5
DXMJ6/0IuW2HNTiYe0/hH7N6t7OTFJuQA5zU2VSkFBJ02OhFc63F9rj50kdbf7h3Qeour1d8AQWU
mXWtB4wdBMBNBEut9PPUdCdLnF10vxXqXRvZODGlDmeNjRTLJz3dWyLm4h0sx/0GjFz8nSpGuR7S
gkybGJwDDqIBTZCwJubwijUd+F1a9OM8YbANqQHGm2hvSgIx+JiFDkjC6cnuo+UA54VQfSNKi2lV
z205FV1xSuqX2qIAWgTO02FxdWSwR5u6Sfc63yDyhdcy4cZHW5nhtpLTjKEx4OKfboGauaBMvl5Z
hSW/5hmg5asxiULGsZjyzt1oIZFArUBJpVlwf7BGH6VuxfJcS8ggqTHOaKM9YJJOpFNicyvbug6w
khPE+L9Tn3y6HOjD7ztGwJJUa8uFY4SjKSXa9v8wqQfoIwkMUeZxaA4JshiXzpUauYdEupi/FcPw
WEoT9zvlsMywuZz7szmlw1em1YH8xFoGbgbeSn6U4qS3W9pjoTbaoJAyUgY79m3ITPbFuT3jV9Mt
2iLfSPasyuGVAk2SD+7X9Xc2aUfdL+65aSFwHkxDsF0jxuvY7Pww/BTeuaj+tnO58mhfVgnHbTW5
dVUAidi+wxMLISfd3rX1T3LWx3knhWCF+D+C7h9RO9KQJxcd7OVAaSc8va5Ec1QmT8hJDRNSC9tI
BRnt6GVh6eNcZU0YTd6dJunaXt9SN27OrkkOa66xS5W+rqKZA7fAupXi+63L4wKKE4DZzFLqGWHs
/fcKcfE19jC7bdnfWLnUkbCEppxivwL7pG6p2p/9FTiCeJH61hDoc63GB76qS8URKnW22HGFhQmL
B04AJc3MsZn9fJC4U17IqUw6mvnFqcmnTzulxDrYLryE40QMUgRGN8k5a+xSC80LMpcRutxMh5Mp
lAexPELJ8eGt9HqotVFDocoMGOKYDUlQgiU9erhS3Gmc8eyx3BV3f693IHcPQ/SWyHTKFYjw0OHc
M+bEhSMwr/o/XrqZqZO0ihMKMFubg6jGTU1MobsSwG6FtnkQdDQPvwS4Z9hfV/Bowg23f5Tw7MNY
SsZA3lduOAfUMMtGNG0fHuYRUsbWaKRm/Ywd2hVZhiPWY72Nbq7el6cx4H8qPSeqiS2zR0SciGhY
6x9S2Li7J/tAwshuBTzoXRcsXvDTbeZECgiKiBrYA5tCwJ7IH1qDynptPkr/spVS6gfhZkdvSST0
ZW51izxNt2nBO/wKJdK9pF658JmJiyjJGvzufz+ieuGigrdNLq81csQ36GHtRNMsyhAXE3mgsWKv
q1Bhkp2YTJQjqtV0nhfolZEhT7NoOv9qwXSrQEfunWzRGWvw+6g3wuKNOUrzguKrg0+rqna8enbQ
g0YfjY5qCKQAm4AHXbC0CpHQ6jR/wZcsPJRIvN2ow2HqPpOY7H+x6Icf9O4gP9dhCmQuuc5Y9b6R
htIC62loUG9okCHUrY5P3r2JxFLwDe79r5KFOBQcJc7zFJy5VhpMLoRnORmSif2c+7boA7pJ5NDi
KB0iEMpt0Y1ZS8+XSkL3KzY4T7qFPMpnCox3s7VFOaHlSuOf7atUpnfwP1xdszaxBvyiGn+WPhXK
3SO3TKpF5zCUcIPHJIMS6UnjkHuFt6fz5ki5B1N7dOQ0PqrPTIFq7gGSzLiLEvHF2vatNlwtoPud
LZioCyurZm2ZppwjN2IwiobdO/ZnKYj/ndd/qmctX+Fw57Q5r6LwXIl3gsdcVkO8KBCTqyNTUZyD
TvzkMwOx4zU9MZlxw+9c0T9rYlisvLOpMHIxQQ58viQLTTLAXh4PY6k1gyJkgxuz6qjSl75S9XOg
fWW5lC86CJ8HJgM305jh5lL5ag5pZsOCq6kmPV2cvdQOydNIFZCdCpGrtAvNCeSsVEhbwmDi5I+J
TCqYEw3vuRU2k8fkoV5Td0Dopdsn2LEO9cuO7KKgPRIZBhHW6VomSSRRAPFGOS04+daGEGoMulYJ
tChKOUNXV8iNRZwW+mSaaI9gwPAcaR2TmRvBiRfacU04s5t5ZZqwPd7Y6o5z+AYFZLoEwrotgbSh
YA/FFyHjyB7ZlwHpJuZuy85fylKgNM7G8y4d+hT3pC9vokbym5yaJywsVlQPpxR1YwRi1cFOJg47
jrKusNFyOy2x406QfB/pONgztfvc7quniMFz5OiVPBz+o8Apukwrvm7DgWBnKenIAQysamJKEFqV
wu8FTWYhoEJYY582A2Niz/xedB8GwnH6dOf+4vKbi1e1+UaF16C+MRRTn6ISDnP5s1E4DdM2GvSy
WBatxJ9+rt0qHUGkPkgGd25ZDUruUIh8LEzyVPxudF0TSQpe960BGQQMk0E6TWOKQoSG9Ao/kNOy
3LFZpka+5zEMoYqiOqLNMM/nQGwEhJI/D5XZBB2jLuPVZHImL/NCGPksPf8arsBFLxkDZmBaiMmM
BLPYFEFYREmmVwjOIjJYxWZVFeTXgTGopSaqCtlvHvqsXcBNTehzDZpEJdPdrBZmX5PrkaEV+Q+j
dzxvx5aQhnS2EJCU/IhwGoWab5+288QDCRKT9npx4TWKxXcElOoqlXuVN4H5nkFWDHgK4sHD0sFs
0tU0zUcxBNAja671BdUhG7TOXNnW7rtILquCzX2mqwlofBNGb1dGHSrRw1XO35qXUDEuo3rZkGdV
1p7hHqEDxE+ssK+ZAoCdlzfdqhA8IjhHMrOmU3Zm1kUgY9XGDs5aFeF+Wb3WRGcyLONJx0AmYez3
vDH6tGeqZaGONcEaEC/oo2fqj0ymjGjQ/eDOOniB8mbNUzoIKJ5i1NkJkuoZXyDAAeaLe+MHz0Tk
/vAeb2IfMMC/ki30pFOLpisx0xZkvBJyPlj6ZQMHJXrIiQ0U0pghLKgXxJnDgITsKu29mG76OE4C
/VxSJoqd0s/g5EB4D/ZN+4Y29t78YQhEateYzG/yKReA6aJU1PooHnx3Gu5YQWx+TFjITxdabkfk
AU8N/KmzQlFp9C1IWNzFO8r85K3AkrkJOnXX1D1QtfmDTpylhH/ulCUHNValPeo4Xq70zrWICYz0
hhUurqHJR14rxweQNZV6v7C3CU56v4r7VNlaM/BfZJbKSIznTNIvaEOvx9wGu8CFRj+7JyWiLOeG
nsLKb7IpVKzQnoE5VRgNEZNb7I4anTPUddU0/CCAPg4sIXBmk1oKr0u18fBQt6G5MzXuIAgxHG+U
uXO0+1vafXYrdYRWKs7aD/AIyjXFiaoAC6we20NHkSlw4mNtKAk6mu00LcTLpY4NdzDG+ZPz0VBc
oppdhXSmvgYlyfa9sRy0e+zzQegDBRZm5BedzlwrtSdtee5fQqzC3RQmCQDGCsKOkNHtqRuC8z7C
GIdxEz5TGRT7PVhc86lYN0lUu5pUaVCCBDLq8wobjRWdPokjcU6Nfe7Q9Q0P94bXYAATZ1jSD+Ol
EDlMYAPcfFFm19zNFFglaBv57E4jyPbkHiOIs1YOIo8JzgKh1JNILYxR7jKKF9xcnrpbBNUtu7QW
63pLk6IbZyXBn+I6NbjSOcCqjofhrA25vJMvTMS4AWyt6jt2mfsxdeAZnTV6A7qiqfE+2jiqoZQO
3I9LB2PkMVvHs/pke3zwST92S9OaM9c/UJ1kBW2o5mf8I0t5M9i3UpibMBDOkgTVSSPBj0fDOQa6
IO/zBzrY3C6z4vxIzKkQSv+lWQJ0wCIO1k70/kykNPTzIrDXa9kzns5tif9V0MMz8sa4hmbaIkGf
ECV50TbL9KXlJYMHwISAZ9FcvGp5k38A3ebzDY3TzM4eY8SNf+dCL2w2cGJgc09JEEpykZIt+zOt
qw+SP3S5KPf3idefY209lJLo6skOvEzon5dm7ZZBT4KbBHLxFglFjwHs2naZR1SUfEJw7KuDYPd6
jcU/x4tYellS+oK9aujPvCd7jm+Jn/81RvOPJPXPWGb6GCvk9SU20Tdzkq9CONJ3yYpZoiOpiEaq
bzkOOtLRL6DvSTWDqCEGe0XBRUyxFdlkiIpLSqvnPUrGJzM7vUh9ikILVT6TKbfqQTX54aDDJvRW
M9B9CVfwnDCMpC0UnHGTkbKKrbwNqeiFxD9X7S7sLjVCZSx5ceWr3uZ/j2F1umKWbf8pe4SX3S4Y
U8AoPHW4wvFFuXm+zZjyOTccD1/CG9PHJPcGLsYV4b8ZQli9+vtGArwKFrE2acg95WEPfqQp4zmx
MahlQfRXMgOj1WSmr4vkXwFVomCzcUkjtFUZyH7UOOPc00N5rx8jWQXwd/WprWq4zTzu7OyzRCxO
WelMKyCMprfmrbHN8g3wrxV/yGHFYHcfj3ea+9B6jhnMDHYTqlU6noVfKKgl5kaUtvlc1DQ4/WMT
6MKxYFPHznHEzke5jWykDFmwHkcANXJbdmtSZSvtplVYIpTa42mMN39Yb5xV4TrHTMAu41zpNC7j
EJIlpn5Om1vEnjONxYXVRZUyd/3ouSWib3ARQOrinCWqDqFhp7Vf57axoh5ul9/G/3L67BUMkNqD
/ZWkwM9ZFLlJQB2PBMElHN6RHBa6ZPw/nCFok+MCCR9rzNvq4jhOuXXY10K5EnKLKN+G5Cctr6yN
O2eHnFn37xXmUfFfER4Xu+BxmkSRiFn1cpfV3d0u2NNxkZQZaGCQ1o7UUxmx0IEU5kAmP+MsaCJi
X1hzmJv+MJJleSGMf+BUDujwm2sOjquyf0hyuqKelt/xSl5N+hS4Um9Ou/oxuO6ClUaO0gVHskxF
TeW93jQb1oe6ApM7AGnu0hp23oo5Nc/23diyX6CbWfo3SHKDHvk43Wz/W2/U4/wrvIzI175KV2aD
W79ciuVhEPlEmIzVLYaAhOA4L2ypWSbJdvr7OyEYu6e48FmipiOVkhPid2a27WxERGbIhD3ZKD6V
1onBBaN3bWfEZx2WLqbKgb0UBA7yu4G5d9VGgaqRDz23iV56OCnUkLD5OkAg8uuFHrh5aZ1sNsOa
6gs1Iue/omlmTQ85SmsVhQe5mDej2kXd3Ibe0gsGIND1IdI+HPx1gqoL9jplK0/gcz17VDsfE0LX
13yKK/vrARbsZjwA+8k/YF5jHihTlEEkmOG5RrzJNY6MfddIoyoWz/ybov+ot2DiNWj0NsbpdMqZ
nsTvpKMkojZgeoRumAZr6DbesDBAl8D5T0kvpOHXgXVvWuYSJNoW7+Vf7eBvN7mD/SgF8rbsBhiS
jrQTOpiLjVlw8qJ6cX938mqQ012lmyRT6/sDY6xLuk7SQQ/1Th6sWe6SU2HCAK5rjELKsfEbnxRm
VATgSQ8yCNT0w4sJBJRfvljllyNrO5Ul7pz4gbUp1/YTyjBu3ceRRm2BGiJn66xHNfriOOS7UKyE
e+93zKjinREgFcbs84PLdS1CcVQqLsYR5ysskD/p7tTs6STU56SyP68sjUL+Vwz/YmtZNgm5Q6sQ
Dst2BPYLxL2U8uylgaFbvkR5DL5JmlPGHWlG6kk6sffCqqkSy700udCcDopqQqEbFzwTrLLbu7tv
yEQLi90dBmhzBNgiObzJx3IY57cy4wkzlLXGR7KPw/P9aQhsaSjqLCW6Z5L81mEG8SjL6U/eVig5
3s+vbFclhDO93Jx7t+udamQM0I/s+zWH/zqrQGvYxHQPI+5HvG8xitb+gxrfnuxcymKTddsBSzR4
ge5bkOHlBqRghSRaVhP/esARamdQRWkWwJtRs0BmWOMnBYRCf/lMRB4SIhGyB4KhSc4daCwa4Rnj
G0FuDnDplkUItLu7jkcFg9CY1v38stPWAh4tN3KOdtdiRsqLVfXiD+wRdZ5Sm5KfPi83I7SdhRkA
yiNHH0LG4kGt9BN5pgWP+lJD5rh8PdeEE9UqjHw94rg7XY/S2X5CdhhYq55kUBA1NsADGFDY/MhW
rajnYQFqa4FcmSpnj+Yu/60Zj9pQWYKpygKYGwe+86FqF22AANdhNdwyWR+cwXa6RYWic5fKSRyQ
50LSxo9/sFXpKaMmPbxZtbLZ14IUwCGkDJZ/j6/hvEaQtM0lap1FY9nRfKRwMcWko5p8ytDdl2qG
rJ5N/NUL0fMShCqup5RXLtd+RzceAQKxYlEIIOI6ixihrbfD5q11BoEYQI32lDZ9ofRVHNivzjoz
QylL/OdOas3pKzS/xnxTkwr8HKAvdbZ3ygLw6znq+PwoiOKzzKO4DWsliExGKY//mYtQ78oxZXO/
EzG/kJ8babE49xeJNwihr/BDKZ1p84YCZAnW9tYPEcxJUddnMFldoVKUnykTlpaSfIRneDwir5KN
2eVsRDga1b2ix9x+HxzbklJbmZ3rcQ7PJuvLfcAr4gX9Xy+wx9FQiOyAhVVPuEbsLimiOjn8SMmS
icxaq1ZyoqKjSwgc5wjxwyWC79c3n8u8EFZL7VF5BFp6hWbpIh4wA5Jkx7B5Yar4t4HWRYkQa1uF
w1n0oNoCN93bb5lFiYtISsViwCp6v8ifdw+VaEo5H82cKPuAwWWaHS1HEncFER2wx3bSxQsWIxsB
MMXrLVXdCeaW3pMPVyTvzmo11F+Cc1bMAkl9r0OAJTQ2Lq8HhUh9cYyJXNXk7xyAHGCMlPQAEyyU
Bt7WdC8D3vsjRXyMfGLyvpTzh8GW8pxlv7rEoTYkbI+V0XiHzZeALHYRY8Ts+PUzqOj1Yb6vYDMZ
/M4gCVJtU7VQY4iP0iZ5YMJnBoYanX7ehkTq94lgWq37vq3l7qMaU18G7sEaioijfFsQa2laaw5S
fOXrB0278o7Q1CS3qoVkD/PC75rGrzU9VxbaE4ConNjvBoh4Aj5Aw/pnnAEz/Svidua1Tsja7MF4
CFeuaON7cLGk1UNajZEol6ZiVFhJy5mRkkwbRcM9yUMmDF/9RGQBkvyd/yZltOdJIF1GXbPd9pyx
txSKbifAA9+XChvZ1Gb/6JiJAqgSw/3SRO42iClD7F1sk++FLsYBnwpvnc4DO/fU6ce9PgsCT5QI
k4mUf5p8B+TXrofN5bDGANO0uyg+YHss1umuFAmgJkNBJwJ6PuBnssulwulz936GBLZVpOMkWfgM
fvg240Ds2gBQWcO4+jqDoI3bjdRbtrBqRyc3320lx1ftGmtCW4BJs560iSGLI8U34jwcv7J75WUp
bBPg7GH4kIwX9NUSOtg8eGn+5JWsU2U3NqYJUthBt1N35LTRODy1hj/qjNDmqbQesX6X/Y04QSlC
fQWANUVxh2+JgONA8qVErbyn0N1esuRRhrz9gplDaLe1j6g0E0gsUuk/sN+1iRKORwOIPvyRphAV
KyeVix36DRMHkYcsjf3AcMzO+CRn83P7UKb8eubEA1aORCM/yTG3b2dRNgcP4idlpZsGAIlDxLuz
myHVQjAg2riQ+/R6gtJJSdEhXo8M2OBdVXbeWwCKZbsVdvfxIcHjuYCbJTtEGwnk1HELWXfEn3Ar
MRZWby/um8qYfuiloclg3MmgNRxkOZpR2gO00HK8YBniharxMMa/hl8zJD/gQee/KgLHIxvYpoVB
8fozDASz5nud0vPmfn6yJp6fa3KIWigtFv5N2z5B7G77M4iRHSAFLw0c2xqRsddHaXMBWMGvySNG
zWnFQ1qtGim6mlTIsvO5KmHYFlezNTnkf39uvWHUknKKDUZ6fXDVtyhnly7zmGZvlYMJ7dnDHPY7
0eS2v6v4zqCgB1IF0l43mUUKFZDddu0u5Mvh6oQeyXfmD2yXgf7JzuQqyycefv0uRWEyQvtQrLJy
R7nOPMil/WZw27DhdC+R1yKzAI1smU9wcZ1Io+OypJKUqVK3gUc0kHPMZUcxKrwR1e6mABZk63li
OAvGCAizkKzvT1Bv6u9HMvZS1EK2lDqyDtjQKF/GmaDF/E7GbGcm493c17uzGpsdTlqiihZLktta
ZThNrRO2IV9MZo0g+bemTZqJ/TfmN1KI2UH6tVO/BwVL1iCUWwU8SbiDXIeoi2SLMRgyQELH9epG
7pspcuz5+INBW5K7KFcbhSxloC49L8a6O/j/r8P3d6aEda0Gw0Sd5SHE4k+qmTZygjiVf1xx7c9B
3IX+9XmwAxEfSVSw9tfYVMHuyIWb0SeZlPHS5D8Xd3/8wtaXj6kLq9HK1DDmcsWo9ECmz/ShifSD
SDOusAWAcegHDNaIgfIQUXqC16Q9yi1/ipSXrPMZkR5To+mfGj9ctpntharj6pYg3DNM/WUhpys3
VP6GnQV4ldMlVgxWmnsJLKujV1G2JDEi5N9tI62hBNpDDDQPB7/Z4NHAP7VAr5Cl+jgNrNtXIHx1
k2q0OYAxbG8VFPJOImLBqdiBTV2kwTPxgSnc0FrIL2wTXPsz9/4PUVP6Kwk/u6rVs5u+GPhGKsL7
499jkVUBpmDCuLjT6muPLO9voqIq5crtz936N4xBtU6VAob/s5EaXeMcINIeb5fwmoid02XgGpZA
6LaxFq9taRKnZ6ivMkNT5OL7+cPW15I/ylHn3BKXRbiGbt1Mf2xDH71HuN/M6bCxlzSLWFFov6vf
tInz08Ig0Tr3O8nsH7MkxowGnS3BLuYU1AlWNNZfh2ZvDcjnu+05mJlVMMpDsenH1wzscU1buoyi
jTQ32By6IN4p2fRNGdnhr0RNddYPfvHg7wgOMSRrV7MiUmK6r1iiLU/PQZre2nvHbS0W7gQLAWpE
au8cb8dL9ru0KEYoaXg5IA7Djhd6eUxKlbMaKIjxL7QMOQ2vCziZLJoC6tBqz7D+OrgOP/2dNpsB
E1hWDk/2g3XeH1GKdfs0HwjldR/zc9vMAnBEpoQdSw9a1zzyfRRmrRAYusrpY4MXDxa379R90MHJ
qkgR4nCcKfEtV04YAt1oqehvPBVzIBvPuc4jg+ZbbI/oP1lNy3kn5IAOarHPrF1FosXhoYnK0DPI
yis2xsP3jQKLwKZybo7/zXd4jq2HcHWsilxfTnt1avQW4wiv6rxIcNKNTB1g22EEgNU0H1AC8Gj6
xq0phoI7wa9yj+aNdT9j+Iyk+BKm2bVW4ITK6oV6pVnMf4bwPHeeKbRzjaxY0fElocDJC1O+JDVZ
DHGUUHt7Dz2ICRNbkc4MIKsyWb0IUbE1peedyT+MHjT95dqHVFdeZJHG2WvdRKLcW37hh1fxpqHT
c+/QsLPzmIEGrM3P/lMoAoIUqj5k4zhnPGLQp0mRiumE8wNKmpfkHnCZpwZQrU2ohTt8gfxxvbeI
dSuBRhKor7BjetpzbiWPdRlSyxqnPKVjEf+x49u2TFzjnkjhP6jMertmz0ZJoZrL8XBIcUs7UhEs
4emzIh+FERZZUNNRAm09a3AEToG1Xkc+nAIeT3rKT/Q/ARPxAGclBLwIj6joBQAgbm01Fv9brnYs
ezzNiF9neGSBAfxDs5TSb22mxecju9GGbYGUPGJuSwfSdgZ5ma9GCdX7tzFI/jR3ouHEdTIQ1H9x
LUy0RrVenOfFgFmTpyqYkSs7mYaRZjOsyzZaiZL0oFYCo7KU09Grdz3TREzbWOj4rRtTpUlalCyX
g7eHlzSvA28t4+s5rxgzSGBj0enV3Et++0w5YUzp/3DFXbQSWR6lMhtjbUN2HA6EzJZg+Uq8bTkm
0lRaISk8hlcnjvqehnxESj/2ALHrbsghZA05L4M4UgqGE1uguyjtIrmQS4Nh+VdeeTmk6nMGCPJZ
plyn5R52zhTXTHnhO6SqFw8+Rl6j89OCzz0udYJaMDspqAqEnbrMvTWET7vu3KwaEj1KKWxQL5p1
0tv9uWmMljrJ7q7CpN4vn7OsOQ4hKyEzpo1SSkYvMT9u5exj8SaTrmUuIlfCZk1cERsZnKwrF3dj
JMii7ogBsmHU2cr3DvJvHwgBFhB1eNnVZhMao2EPDIb+tBI/6vqZXqp8uEIZbiHpB6LUCc/O90kO
LmuhMa0SPK2FHmMh6E6vJSDR31gPqcdh4u9apCxcfSkxgjXbr3vylJll6H1FyaDFMOQlB0EjfVWu
/JyFMdYf0JPyOik9IvLyHKvFAvOS1kIp/xUto1xyOEj+zqk5qgAF54WNF/dvRtj8EdO2bCrVtUhB
hu4Z1bUrGx2URsSARfBHTra6zXy4ttZIyYe9e2SGKoF9RUhkIiGkPOIiMz9dw6P5qHCzeTcZTj7F
nLsFZ48KmWMDkpKAtPB/+UY1rJNwsTQj+HyypJbT1Zpg4YuKQX5uMuNmQwHxpRrdZf43y5MbPeaZ
oRD1Qzh0JT6hdbR4KqBAOUB8hLtCu48UtbCTJYdx4giUdwvT8f5/Om/jVBuCFlMvboaj5r7UNRGz
uwdF1g/NcxQ09UxpWrDmOcXXNwZhfhja5gbm95LkeRxjhdQKmGNOO7vcgaP/GolOac6cWApgKm3w
+8rGvC3Vb7AbwLhiugIml6xF1LHPWz/hPGgkt6+VIcMVb0KrvNRK8aIEo0NaPX9nBNHjFPzJNsn/
L675Rydq7+0DTXohKgm8LJzD08dOE4u4I/MX01J6MEKynNBPQ77tkVzWEM7JLWGiPBNIz8IQz+rP
Q5HwvC2jHjirGH8E+tWd8GfXmsVv7OfQp5mjAVZse3/jC60KyAmM4hWkvYS4tx97xsZdjckwofat
32FsNTQ/jhAYc6ZegH6acqsbbasrmmpoLfLA+kW21o224WQsTP37vropVN6QUfByZMFZUYIYdMRQ
HsjpQ159+WhZmzv22S9jpPIR0XakWE60kqp+si6mpv/OCl9D/adCg7QyTRATtg8ESJHgp6FrV2c4
dr+EMHQqDFLh5GsEopqKC3QAOlKtKAbBoWe6Wmonsg8EiLJ9JhxMAiUfZDF/kffo8PDcRWOtqaFH
RytwgInQ+ShEjuSVWYdIkYEDUig2aPcYKz8/5uZO+aYWgHKTpkVWu+QdjPA/J6Z0KL3H3xg2cr7m
ROmyjmkSp5qqWS3+TOVfY+x9aU2fXLHDzDmYE9+E7OIg3uUeDv1kXL5oVtyelj2hrhoFhIcCHg3R
pIacnVA2DnO9HfOO7PyAvzZICdGASM/mEgAUC4LxEXxVMCnz80NqnrRPik0L7s6VpBeVxUW3rGtp
ybdcIaYZHGcCDpXuhx35pVlEHRS30C0mb3PGcU0F6bYON3fq/qO8mG1KijBzpELxgmYc4/61yX6j
VRw2yaVnzFs5i0/nTD+/ILfFCBaE4ERDteBMT8p/Gip4sCDnFQjG7vCp3Cs7RMuxEOTIkYZVMhHg
MQc8VY+O+pLFpaMX5xXoMKr9KgKcHArh4AkAtkzbKH1UIenMrngfuXb0UWl/xJZTffTLmErgGtqw
lOXol5k/kV4BsWNBncSo/grEgZWwDo+gcrnnsF1d1Tnz6yg0pVf2QaofPDrtsSWVfqyxjHib50nF
oLF3isOYCa0wuUrrtFzisaSKEF/WKK47XTsCTTYz+JfukiVy6Xjp3WQghYEj6a3guL6LK9L3vQvZ
yhCiuIerowrkOBiWyk7YKuize0BCUPs7p9aMq9fAqVcTjUTS3nmnSRhIRAZY6/UmEhbGlwM8ytQ2
jQ3S5j+wXQ0esWi7lE6bTDqlMfQ+jGpDuRQGbl98nDJMZaMzbl5LXRz33pi8pvMSORfAzijVdlna
BO5PzxIM61kdGd1Ayqf223FhyqPTDOlHcepeOs4thjvcPHfYnqALVVxGVQgClSlVndwXX5QStjmm
/J95LoscOoir9MxjvFoseKXPR4Alk8UyVMycrMGRF2eevlu+4cIq3M0x19GeER/gbNOREAeWuR2b
2s+xaIEly2HTDu/4z/PmeYEeVi0yOjhGJDlyR5KtH5/znwLs513uyhmTbuVVgJVE1k7EL3D6ex9T
/wltJIidj9AK1oJ6WCt+5UcfyDeOxV78S0ylsxHWXSJP2EWUN2ZLPFm1zmsvUJzD7QiA+XeSKbLB
UUrAQRE71oJqhfzinNyh+7tlmy7pQs6fv+iQFy89rUBApmoMOktezxY6R4QWQ4ICDFoTOJUGg/bJ
Ze81qsXxduels0ZKmbxAZMynIjVFuyMCUQWHhu84Wm/fDd5FSRU+kxZDg+I4XKIljCt81Fkm1FUS
HsmPBcIbU7TxDqyac+wCD3JeTaRupAufFi7pD+bwRrayEfSSsGf5awlfZs+2HRDfcoJ/fNwTEGeX
TmTwqjOm/eUXI8LsyxolyuXOX+d58r9FlY1rJ5VU3ttisIewiUXZJ0TjMwWOrsJCjJVqSN5jptIJ
BXrcopTXCOgAj/42psSYXSJM77W92/aimV9Klrlhkn0jZXQiCG/MI7EXAH+43BTlvgtMkaLA4SHr
v08CMLkbqtGrTddhHLnAuDmDGCqcudX4l8svceUM8wSAp2C/TVyzXtcILVkw+vPXXdM9zi+hVWeV
I+u0Njn9PGyCJg+FJ2Q5elibDQAkkqI1zClwCn1yU0d6041kaKbBoBJVj+G1Dnmm2LIlM2k6bmsr
mLJGbS5BlNg2V6hWQOwJExXqfmEb2GepUIsNr6kDkaiA5f/J+TzvhvH+N+jJFf3F1Tg2AHnL38f2
RsBYxVo3QwlnGwgNOc7jTyOLtDic4xdpo2ufQOH3MeIfN1Io0M6bI87rnAhqKRM/fxLuz4Ibh6pV
+aaBT/A+Ovr4OxAwDnKY++IQ+Bia2yxwcVHR4pE3oOx1ZBz9uRp6CAa+SzHG+nsbsnKN/C7c5FKO
cFR4E4WaQs9cBz3dIKFa21ezsptAKbIN7nZ7r55wm81P3Rzh5ynDnToK/pS3eEEKra513QiESVP0
GA2gr8JvOmrwI0TCSJfOS+NGng8MQx6azuL9B8fSMuGhELvjNo9LuKvtXisx/vvMroQDSrya0BoE
PApf8mlB7HdUds+cWU5OdcWDSe+ppOq7ldj6PV9t8s5n7UAOKvf0wBUYuMzgWugpcgVrZrQav486
nU/cTamFkfihEznEPDvudpyP1jqMknffzXsEltO1/467qWPlAqTsUhnLy1Wk8b1QUp89P5N6yfub
8dz4ovOkLN2pj+c5WXEkDiIo6cXLo+b6lpqcvMxWR/4BuKEdi5qYG2ZpdkWFLjSDLDjm81E8Bxna
hsdAdYdCCpcMNoo727ZA+pMLO4U/9hUwmymLmKOLqAbpWW41v76oh2vWm0upDyTPtP0rL2rsL9s1
Ux3LI8i/V7kwY8OmaALmHQWLCKLUUsMxVhUJAr4eoX+a5BvNPQRridWZ/l94xQdED5O+QiWh78TA
8ycNoajlfVuQfdajzlxG0LdpW4m2aN28sZyhoffUiQ47WAitqK1b/YeR3Nk9dLpX0f2H4nExi4UJ
4Asw/PcEW1Sv1+ergVbwy8GPsfVBSn93sRm+stiJE4GoF7EbiqJxjjC+QngVPrKB/qmajRM9MZo8
hobhAHXdPWxSVxVh/n94MdsHdrnwhr9k+9JreTqSMVqN2VJCoGyfjRaRy+4AVtVQjRvet+wqdbda
wI7BSj6A39q9yLXD8SGAPjBxfFUTdiyUaMkxNyFAbD6bys7Nj2V1byAtfnQ3vjTMcuQB7ee3LowE
WmqSDsv2trsblEjWuX+80f6wsL4ODL03e+GzugCPWM7TO0qErG71vMH2cMTwZDiLj3Id4X0gaAXZ
5rIK0H/bPOEOmWoVrDnEGhwdpNZXTuu+FpVxU90dv2QtVU0YSm1JC3N6emZWjX9xUlPFqSWgBvgT
vuQ9Q6igr97+7JXiUXkQkqu0UP5N+oKFornvv8clRlVE9u7pQ9MwDgC4rpc9EuYe5h4V6NRZNiGl
mWLYTrYqg9fYOg0Ac9yk7WkM8zuHhnQlsMSeS3eVNMrqKhbu21EL1yFACt4OaflB4fRStF/tA2Ck
lBoXunWApLLnzpTSVsFzS5DogsjNKxHs8NALKvy1oJx8PaaZC+mXOEGDVsBj0P8AySlEQcTSaBW3
3g2+VeFrGBy/TMQj95a5CnRzqdGogGCXDhwUpB9T9ZUu/1+WoC5K8wb54Ya2YvXpT2KUXAnLnW6T
Qlf60JcWrAOhrVZIX92Z0NGrManiWYJroNK6OY1cftg7pQ9jeM2xCM1R+BKG8K1I7rRmZePlNdcq
2fsiEqId9paSMibNz4c2TicFrxBg3C+dH54/Xp86X+IkTAbs4FndzvCqZgwiv11YEikf0eHBTtZf
2DJOFDcPYjwN00oOiSQ9EX/2kDm04siUEn8WOlldg8wm+e+XNpiTIx1uRdAgkhPSAD881SZVCoo/
KX3RMDxF/cFbIrT1E8R56Pkk8ZzSY8Vtrqdmdehz46uqsvekibqZwiI2VmteQxFmogY/HLROeypx
zqZrCNfvazx6k6zBUwVpEN5Eb4aK8yI3Fhk/3/QfYQtoXzLE4ijxsgk9E42dyI7hu/y3dmPIPmzS
C5t5PLQbdxYLCY8PB83eD7XDicv1qEPsn5+bzfzOMHYG/a3TcNjYO4c+6wQqEnO25aqv2q4h64p/
c+139DaW0o9fy0g00NQTe5Ru69Ex9wmrbS3sg8il9I18WiOOqMUfmKBW8zDcL9mAnvq0AB1kNpSb
k1yKCI0aSU0vKBkep/CVsam96GyKBurbxBNZmz9LuxQ586LUIjOJij9JAwpb6LqDQND2pggrDbtS
8NdFmfYAtD//R72zQ2fdTpk6hVRnp4FmHc4lb40lYkQkX0/1imlTCgOBgkr2cpVFro2dHc+OeaJH
do0LmB6JIdjfNfWwj/NKiXHbt0xUr7hTqOJakqugDGGoJIMJ+hMzmGR8HFPjC9CCvyY80eW6b3sk
NnNBlqWd3E4nEj3B2eh00fKbs8meaXHd5jJzfL2mbof9a8heO1AP6/p+pwy9N6LeHcWGniJqHHJ+
DoiygTtrGm3j9T2S4qn2VBTQ55E66bt6rFNpVk6KAPBFH7hN3uLoflBV1cuvXVCSQ6PpDoEIlFh7
Q2wXVV5IurC6yoTqiNOX6TwDAnO/ewK+hzTMqxTg52Iy7Wak0zyL2x+7m6Hdt/0xMsx+AATMHynd
EJ5TYvWle/ZdwH7r9ADqTFR+jc9mDw9lW05uw5RJkQot2B+DRPXxM5Tm1Af+kMoJ3rM1ms9kkyJl
a5M5HfgN+6v+lKxKGxCz+DZUoKTPSRYmc3QHXpW2/hFzPVRLSmTU3nQLHj6sDjMDstGL6KhSPrxB
DLW0LOnh/3WM00E0eIWmLmtJpgZnhtdYzjwr4sy2sY0VfC2ihl3nfQhzyrfh/Z8680xlBox1DABE
vKouJ1YGLvMwgjigik9HNQdJqPdPrYnzfPaBPprDjKmT5uOBm8mo8VxysB5G/1slFf9pObLvNf5E
gasP15ZVjgBHZH3JsyVHKX+9RM20ev7x9dKziGzznSaWmcJE6wKOLwd4BXiiqf2Nxl/vFvqBJpDx
Ma1EO5SSkFRtfIqh415scNBAi7KN60dBr8z4Q9b+LVncfCRVL88K8gdvnxMKLKRVhFL0aWvCxJvu
fgwTbn4FjtbmRvXiOwC/lKyVF4aDz+gm3fjxXdGyLJtSTOoNv15AvSJ4ULEEnk9spMPgU2k67nZW
pnOJOBG42Oeuhr0VF8MKLvUzP3ZNTNqp7oTepLf0sWm7MZkWJijWy9ESZCrdyEZJ3PUMUiSpYPDB
lQif9nhtIy4P1dZiVw4E1M7bPtZgOldMBBAn1hsjPg8hULRC1Pm7I848Zdk4tJoI8BYOzc3e5rEk
MRjNukM64VWN2xjv2d/vRLH8mZAdpEqzCDQpwHYUqmI43wEtSg+xkRKlyMftwXc2OizjH04llVA2
tltRPa99SdGHSQnR7m6N5mE7zpqJNalEJx565MXU4KlTb3CHj1f9uYOqUgw9IorhQ18Xgy7tpvE4
hBPkkl6Z9m65onn2Z+C9WMejKKXtYoJGysLTir7+QVIcjCxem6KfvFRKwCIJ2gl5qUftr0FXtKF7
ZuqYzkp/BMAXkB8VCee9yorBMDth3RVA9R1ohYab8ytDZpLavMNH2/Al8dlLDnq6haulWKFcfM9m
aXCLLXc4NfV88XHV/eisjG0sVz67RSqdXkL3A1gIMcg5ZWw8V8uj+HTQ5GRZm7ybJRUoetKMjCWd
CQY3tz5PFuF/lmc2m4VDZKhEB15G82XS35pEcDr1KxXc0RwCGbcg5JiaHifccwSnQf6V+PWRCSEz
veLD81/shcgMyswLDSmvGeE6BR/dmkaZnWRw5IQxboyf+iBlChmMA03Rp+Kjcrh4KTZoKMIRpfxp
fGmvq/c8j9G+2DRwZnxaJ6g8wjNS2VAVxMLyF/MQU9yMchqGIN9TzBNRGubGIQ+qFUaHZVkV57L8
1QLm4iLw2azSPj4Z9Ugg1O/ljuU9OeY+6e1aLStC1sP9ESx+/qgSy5sWDGLwLZ0H3St16uagc2D9
jH7LbuiePy1RAWqs6osWmp7KiVePYBLqGIG+Q9lQ16WwYYvUDk3GIFm8HwQ0uX21FxQu9Qh6jaw3
zewOMKwKRogdTJPJjkY2e2dXCgDMQVfoWS5LQAzd+5MbO4RzeS2Sr1pmmB3coeowR/QvhEpw8lpd
IkmT0zBMSTSc0NA3n3YGT1F4OgZhJqny6uXaiueEQg3NAHn4WNiXpbVhuWICygNer1HR7V8PVrNF
Q/qF3obf2o1AZFmR4nPPUzfpf5DHFaoQuATK6bO69f0wfEzYSoeUIEHQOpvDmA6D+0B3yJHDDhgL
5JlA/l/L/DuFw7bAtkSlozoDQuc+U45GwI9ubvu3Vq5Z5bmWS5g2bzFcoJj5hIrhmnWZPsjGbJq5
deOdn/vA+E6NyeRFSS9E3UW9Fb2+xubZd9D5VJ2GCF4coFMQYHO9mFYvrWHOCaGh/RC4xCtcUmtP
aoMVcsZa6+YtA0YIcN99IGJovE52r4NBTCihpa3Y0jfGjnGjKO+S9HSOGqCZwenqieBLkxeOFRvk
3F/xU5yWEfgckjK2hJ64WLt70Q+JZxACXPddlsVBvg11nyAYD2jDGfPJLCLCzF6AJiN+HHPPV98c
UuAQC6n+GTfchLl1Y89apULSCEuaKsV0nIwDegVENcMEsqj5WyVh6SDHCwBcHSiE9w25e24OviCI
Cs2A34AGCWCtCHOqKcMZkBIS+lsmYuRiLQZmXiJ7Jt/KkqksDX44biScyT32VqZrzz0gOuU7F57G
bHtilXFl5PvaY6AJck5Wns9kALWBLOhqo2Rp59WXToT4bCIDkTGgSs27JbDKp7wLy3gZIwK9lbEm
V0aoj7qZEJwnj3tQwEW5laTiINWGoti6CzUVgrRyITtDXVm9ZfnBV+CLKkTFTgpD/SwwF4qlRYxm
I7ntCnzzEonnIgD5tBUwNUaTb1LlRrxPSzjuPfXxL1HpN1iHIhqMV+j/x7xbF5APU3BFWu3pJX5H
ldQKj8aYdQnSVFc2+Yd/tRVk0WgCy5IMSscGj+nTBoepRhDQpqWvMCXGhkgO4guuUp+c9Ju9cngU
6cqnFT5/9/1vHafNFWEfaemd4MRAmkE+Gs5vosa+n9Ow8YF6oE03dch/pM2l6NWlHUMWP/MBPhB4
wtX51SsOnZkHIzHHIVtwgS+8seSri3bjZzPJyjBe0+0DlTfgTmelNVnLM1Jqu8ym5qF+cAq6Weiu
sCUc+rG/KGi8Y+WCZ+TOqnUEaf65IAdYbAvUqN+Nyq7TNn13U5UMwZptxQPC44OalPoat5uCtpgU
zMcqnJv7zEVFfcQsdllOV3cu9yyzh78XdisFrSpgQm1/C8XoXUinnzeSQicnyH4IN6x8KW1EFFik
rT5ngiaN5wA7RqC2JvUG0tKDxWg5EmSNShAHAhOmCxdsnph0ut5od88pqPtYIrg/rP9+VSTjAUT3
p4108yT9Ucnq8t476dC9/yewnCG8Ok/t3io0ODHMyfTtCjPygkGU5cMXsvpTLYChxIYMa24reYe/
E4hMAEByAV+iTV8U3nDvaF5xsMZ55ufgP1dUuOzEum33gl0K3Bxji7dzXHGsji3xCNfirJlhBUhp
yKFF2IDlX3cmQGov7aStMiiXOMI7qRWniukQwC/NkMNjVGp1E3gzBruOpv+vBqngkI0M5pmgCNOC
C4GctmcjorTEcXdI2jDicLEkLiuxsqa3VCNUJYvQSJNhVspwzqCHWjR8VQxsWjhxEOqxnjd+4ang
ZuKRqBQBMklEIqF4bA52gFCqIcTipXso4Z4aylouBtqoXiu3zaqLmHq4ku/xx3Pg4+30is7oj2PH
0ofQ5DbiG5zhb3aGQiOWaaHaajHSUYkQ7ONTxN7f+w3n3u88a99BJ7O4/dp6C7IWOcRRbt9aViJ0
AoJd72Q93q/aSiCNDwCGT9FF1b3ntKASEijOJNZ4zd/wxqBtB8sq4l9ZwZI3mOL7X9NRAopLJfcJ
nDW0oat2M/Jc8S6/HgqYwAotdtyzIiFbtLVO22w2UmZYuKB43A26FeHsF+kKEqDUqXQpvrAqgb2O
S1u09SSi3PFXsbkUDvkvWgcxL5CUwRYRi/kk89VxKYui3tDPekoeUPjPmgaRDwdZyeYdNWT2xFd2
txXhPgj0mH1L92HkQgVvhruWA1oW5xoCBaIMQnwd8buUhgu+mPeLTQHfu8fxrVBkhiSlgOJat7Ql
KiUX3iZY8mIE4vFqxkTvAo1BDaoZHKjj3o8bZNLsgB52qLaQNP3TQFunRImkfLlvj6B06lOCluDU
JNGxRvalK6/TEMMsbwQbp2PN1MxAVewhQlspdXGZFHhMY4BcNlCaeFg2BbnNcB+vJLA9nDKJwZcG
rs0WClKjr5at23Lhfr0ljGhhbfB0TxHqC76UndCtXs1bNCXkDfimErJ/jLE5OFA4oMYmoAIEHECR
6KncufucNjqEScsQxfj2iWzBu1fiHYJBV/ePmIBPyvjZqF5Z0dn1LMPH9xR+HLBNuE38fkyRi6Ig
d4Sd91pYMtzSb7gwrZFbBPWmU5ibySprT9+TGObvKeAdHvFuo+Ez6J8i32ULGaxkNjvWWcvlYDsC
i+EOpXMeg3bHoJJPGXKaoHV09/DPdhBpk1aG/oGb5wqlgsIgxx0c0S7A9tQSII5dwFgtCp+DQLe3
az5ffNuKDl+sSOaUOV7KFgaYdlYF0WDuqcV5FsogRIz3BbjR6xPDtn9pAwsuhEQqMvj8MCu3M9At
HM+LOaiUWtmnZz61Z+w5Lhi1lD4cEnWry5jXxS3DxGSOSRhS1VN/ZIdAoDCQ57534mdebC9je12k
W2kiNAvud7FRRtm5knxEV47okHLCU8S05DqdDlPuySg6TfSu69/Mz3QEmfoOQx+5fyoKf/j0E77o
BQFYQzB18fdhtJVAHQ8keJb0D21xOF70uAvVrV0iXav+Ldhu8+z3OxGeF1X7rXYyZW70WSNBKk9V
EA1OeVBvSO1tArDgZ9x+dXMaGOQ8ZQfENoKeLEc3kF/xJZ5mcPIWHsfzbU2tmg2hJL1M9y53c4oV
GSvOyI6+S2j3oaLlkW5LNwviUsEHl6Eyd8N9l5rFohhQ7EZ9xMVSoHPf0+FSpjedK4AZOR/bMFyJ
aPsKjuSURj7IyZhaCeh8ycnZRkUFlWs3gVYyXqA32P4WGKg48gQaiTN+Hfm4qMNVMNNrrjYQlZe7
uoMeYNe2r2uLBNG5+dhDu9KdNjLhSHI1k/fXh9ROoEquIW1S9KfzmTbla06Lz2XwEo6Ki40RDAvs
BekfkFXQZSmKIz+96la6uH52u4p5ooX7W/CgUyqwW9m7TsT4AXVNu3SnP72QcuuXyyq7y15s+/Al
JxxcxJJ2HrugfSCXD5Hm5U+PbNrX5K1yP+99tmrZe3J9/vqfJ/ahWcJa+QX3jwS7Ako1ZbNsYx4M
O3YXotJwzM0nzTrTeED/tyCHkJ9/QkffEVj+JRLyUqHf5uekJiSIwOPJZBvAUL3HDYDg9/uVAmM2
dlyshZyuprTLNH1rEP0u0ASuEtKSMl3HPmIV8rbb4XJx4j4EvEEQHQBeuxGASzvY51rMnx32578u
jLTr862tYUNXC5UrYi6mGsQ2GtCTFTf7w/7aoeEi5ZZTaNsds5Cvhkj4F7idhEe1Z1hzeVMSmK1o
3dtDROKM30R4svx3oqWAegWJnxi2yQuPh/i49+vdm8V8FAbZdnyODolMPfy22IEMAU0cxkqqevd0
IKuk7re+292AxjvGTJx6y8FhDH7TymiwHYDztv754YRxiP5Moj/QRUIc1SANg+FzsgTJuqQdHKNW
9d8BAr8+qQNiPm4WEIheNKXDA819GyBK2gtE69Iv+kiAkBMLKqikhLzVH2n8VqfrvojqPSml3fUa
mcUgWXUv8uO4NHn9D8HnapmkOl9t+KvjDaVuqL/PyFizLdvDP8c2J5hhIi3nKJ3R7LdzaBp9bwSi
V4ch8Uh9AA8zxId0uiOT0bfvZJK8XO2QwnT9Y3GUeVLxXtYYb8BHrGduy/MfTdfe8a1mfgfTM4gI
mnREnvx/JC60i+M1H6fPE0znLz+S+ufqV+o3Yp1mtMYkauvupDidgg75xm8nd2w1f4jTH1ebTRxR
RzVbmC6yCGNSx4A+L+RZF3/QfLwgrg5Fk1rahJp9eu2Jt7Cj1vDXiIvvTqWszcM2THNscPwbgDbv
nVXcqE2raYhheI9q35GozPqHa9P8ipa/eizcocO5sU0FO10+uIdT/wVZwAN6NJosgOLiafwl9Tq3
PZ4zesCQTXmKYZpGEVGqfXsEj8XizYYP7hxaqxydsGk6SuGItm3MQDyiPq9nWlT3WDwTCAVLxOV/
aou8wrN8tgzfklvGsfWTe39uqa8FjlV9ts9D5t07HBUE44ODPQbiq13hcO/RWH/+DHCZ+GNgIW5j
FTcoepWlh3D1Tz32yBh/x1w3SxIweKCD+sTctWIjY5dWUilL3mv681qWNllkwDeptQWMkioYH/UP
VOSG1vUJH7lznzoPu7v5NFz0KRDMN1+QKmAB6eMwYVjh+vFmDXyULSkXVxCOxXomctjx+J5DtMVn
6LMoVrnIILVgQSHHC3gCHWPGK1av3cmRf0HkIfTQ1luQni62AAIEWsNbfKMRiFkde7FjiGcVqXx7
LxeL8WzUnJ9jh+RHxJ1knbT20eGkKCpIvK+/t2Q0yVlV02vvhObbjOJ63nqpLErxW+/sRITnVWBo
XCWXQ8HXzOhXhlMGoPE4MQmKc3sx8iK9rN1FJ4DL6q/sGLU8AL6+jURwYXi+XsnvzU/5zPwbfp2r
xamteK5/b0KHly3C59CljYdWos5FNoYDvDVA69ZMOl01pfmtEUCF8DveH+qWs/f8sTUO4qxc2BbP
owGJmownnlJKnZp4mIWqnvIe0nrhplN+I0I1Ns27UvUDmg5Q/mLwZwhnF854pszBFBXHjZExuzZy
7FOc+bnc6XS9UG8BKmuyLkNiMw2NCw+HmrmNJQ5kuhGeHjf58z7ffOkfP1SGFi+AzyHlzvv3oACf
bqZtYGKmyJpLMxFbyqIbFQN6w4J1L+dPWj82x39YAVzEH0E5X7xj6JTUgqDvykvN7j6EjydFNm+k
Twtehx3LKnmyReMzt1GJty/gUlCAtpUdO/tidGp07/BM5gmN2q564UPkWARYDtiXhN5UgscLXinQ
iwkJcuA7D+2Sje8q0avCIX8f+3RbSLjhzERn5b+O+ln1dQ/tJdW4LrblNUWaON1exG4pAKdLtYi1
wcOvHSMXb581O60cGD2rLiotmZgHfe+w2SEdrsCC9ha5U7076EXH4Eko2eRqUysWizlw6vtPSrcm
IE0FTw3EnrT/FkYSftjFDNOMHxD7JkWWWuw6G9a7bADNsZY4eiR9kC7ciRuzmlQtb9ITAcUcvzf0
B4gMIqV0UYFoB7zQ1Y/oOms3ApaIm55wmshikKMXA8EegR/alWr667e+dw+UfDueFhkYpZwSbbTL
uZxdWbmpOWo7p/1Tr9hdouyowanRn9syLx6Y+X9FdTKbYMRHXFcFl54xXnBeEMrF3ScgJhIWZ37l
PWU5N4aki8lPTXDT5RbI46vHKIWQvhWD3qOovBfEMNlnLI+CulvQPxOevYml8wNI3eB1C16+ffz0
UVUJ80RcqAD63TXSBIG4N6YqgiZHLAqvz1h3vvU3ge+19vU9wavsa/NsLLF8l18ABweWpGDI7I9N
+fFmT5gRJs1m3SFODCi3a0T1T55uEUGZCrLyCLINeiRrJO/yVnppJ1o3g9nPoKR8Zp0asQG2MWsl
FpuNwOh3Uh3lSLYAa7+SNPXXGJxc+/U30snRLwz3nlXIgQBv0qo/I0Ptu7P080iEV6q4wApoxPyP
hWX6aJAckLt0z3WzdbOwU6H0frL0tj4fMqo0FZi8+BVagKE5pnDLHSS6xguX0PcqLWdY+IVoNuVA
l5kvd19dZC/NVdvsN9Yun4s8VBaC43C9OUIBKCB24BrU5e19/LULq5Vwea71udUk00EKh1D9pG4L
BRaxOrgBKS/LtcnvCl8CQvRWN/XHqvsvcoMCnkeqX8+spCL8Gnkp17ghybgfeY6BCyIPxSGAuh+h
W43GMN5NF/xS2up0RZSEgfEjKL02v6G7ibFBALHIqwCzcO8O3vCoaQXmULQtK3qoGxukPEvksWCJ
5664jwGvOCWETY4R7yJWSrAths9UeggIJDKs+SS3mMeJ/25SwIZALofbbU6GuyeD/p94UlKueRlr
AuWobXDsw1o79XPod58sAaWumTU9qJqth9YNcDbBsYnZPbNvx/sC4pVEYTYUHt/pNXz31wMLMhrC
LI4GaUfBdt2nUfIFS2KsdNI3FLDHBr7tY+uE6VSjLJvy4ZrNerhq/2wqZ9ZsSNU63ll+PlI/VN9r
/BTSX435FzDHiPydvNNH9hWPvez/+7bj/Sw+4Vs7+jqNtZe/jXnp5Yc5cGInofGG9SmTSDFoRf5l
lOwQDWSJvsTwRHOv2ClxyRYWuV475R7jrZFhSEtZUOLL8B7Paj9SWewbGrAVYB8eWTEvRjjArxSp
OQUzMe5Rz4ZCUmCN21mbCJO7+LRl9erlDwfwy7VbcdLBMG1Dcols6enHEc8gYbcI1sTJNZiXZr1L
rTt5wqjkSVyAd5Sae14auwxrqpB+J/jR9ngQjTKewluS1ywkwntU9bW/Kl3uko3eSH0edmTBFcQ/
I+eL7Jdck+2HjFe9xlRPj74ZZOySXVb8dnMluyqTiBLQKysuiVbMtxLOMfgsEDQibNxMPg8VdHLW
vfH3I/z45WdmbDZUa1uOE/A487j9pPwZB1aEanl4b9ND+O4fZd2hkK2vJRMIIZ+gxOMjDVDATrof
7BMPDWll/W8c9tirt5keF0hOMqVLuvJmT733hF167Ne20oUNhFPRcAvcthypyvXGcoX49R2oSYI1
e1GwA1JLxxyXgl7+muOiCEzg7A+QMxn+kp9NDkEqlCYzbSvqWtVmp0yA1r0Wu/qaCZm8U3I/yhaM
WxS4hy8AyjgbwZ1YeFefLNp532cwkkfQLGo5uCGz+2liQ1s2MhZjM0QWiJ3IpaqTGFZ3LoWqBJPq
WeUQ3yVc+Avw+Mq7TcPFKuTfKg4clKQ9XKeR1PpXDsrgSfVBDkkf4BeLUCImX8Ahq2xTU4cLpVIF
Xub5Qpy1WCQV0NAxKncGdsqpSjFbAPHlpHNQ/SFNovwTip3E1vI4eTzOIC7i7uj5vd3nk7VD4d0W
IaAMnG141AWtjLLXg7TxQqR/dp1w8Hy7nNI7IRd5K6v6S5xojrKiBvN31z0pJupdLYAZ0l3YaV69
Qj7sziDzwbGMXEM44gSDqsL59961AUdskJ2Os8OPLzpUnlRmOehl45YiFii6InmygPKRjiP7HLO8
g0vDn8Vvsl7JUfVRPXFRVKOFwjlT1nL0V0RKrWRSjnxyEMPBMcltACWTyx/7kc4KQ73apc8vdN4n
6PfTrNDo3gJN9eQg7PGR4hSflhzkXIr95EtUKgbqYsOmZoPACpH9xsShYge5MqNtgY68s20hrIt7
N229z1UUEGeiadvcWMTE+vSYUFe2P3h44upfFPIZsX4pFkX3P0gvT5gapxc3ZfrKXWXmEboKnS7W
sWtIqRxUmwrJyC2ii+886iWmQtWsNXuTT+sxT7ssHdkrIbVbY1rDj8W/RCCjrmqMW6xUQSeiFXx3
uzPZERNksNht0iVQJziuXV1PZ8hLzu+n7eba7GA6Fq6MnkYBAnHEKAbGn3ZaE6N4UTdxF2esqGHP
Hc7Vgh94wZLbn8A8kYplxIINjjrkEWnY77qH6CchBrb/VRfSvzu1WvFeh0DCZtcX6eeKUSKz5JeP
WBPL/4h1L8SpRLWV3kLVBvawQjiPhoXN7JbwONTyTA6Nzy9u+uFHS3mULBRbzJga14t7GOADW5Cz
89DRk124Sr6xFx+REWrlSnS4FttIK+eaIOPRrvxhazHXMX1xORPKdyeGKNkh0qath2i2JIYJPtM+
AuotZvrKqNQK4wMF2fXnBLVUZyYBWOWHn6gBiXV08DnfQ/CC2KpQn1/JqAyMzzZeKbXBEc9qqjlK
MDD/r5fFKgMREDolM0XNeub3AoOHBMVsdQ7FsCANJn2hLf5qjkCIFEoMXhWhpXtrbgt/q/0S9Bvh
uMdwwTXmDx/oKVHQ2eUbLFuklb/aoBZD6AazoBaelIKLXTd4xkmV/e/ZmLRqjG1b0ncwRRm+iyh6
bEu/Ouvx2qHaSu9KjWaoS3xQcs0yWYAQw4CxZSOIVG+3kKQHRyu8PYpD65TOQ+PSM9q8Eo6sPMuk
dZppfYfa1UJZdylNYBjCxorW0LikQ7rIsKJfw1auQHvFKgnrRkwem/H5wmsCLveD5Wl7LLy45mQg
A2G9xwyK7EXzq6CZa+cfOBD/XTnUk3XSrSIJkUnRexWOZXClIzUngrHAJb4YfQusbXoz4smY6j8g
Z8EquEp+OGC+dbTDGHUPTz47MxqTJBzuE64RkHdff2ZiYmWfaxL89pN/cel0Ew6d6Ts6jkoXkoCm
iDtp1qqKQNX9lQIh/xynW6H8509M89rnUiDKTQjGXranVxa4BNdpbR0ReJnSTvdsEbrR+ArK9+6U
qY816BTYHPL8qvJ9quU9S5SBnGe9+zWp9ORjEsRTtCRZisaZ67/vPAobKbns/HBoitAZ41wPGwGJ
WDSKFTh0lkR0Y9nJYwkawctuCcSCE+0zFGbEzW6BrysVtJpsbsUuugSsA9tYg6+JLSvWscRY2i3x
8j8LZLgVEeuELfxxvYPDyDv9bFxc4Assb+PEuZ7yVB9pKLNH0VKzqxiB42Cjnl9CykpujtUq4wqQ
sPJpCyQOnmyd61zb0k/7II0tR86aX/hpgKsGMnUcdA+7yXU2FCnv0vIjRUoYxKt5ZqGBE7PrsSJn
d3zAgqeeUVUwWxo2YZ68OwmiMC5TSxEAYu2kFpeAY7DY/18Bx7fo89rrs4D2KC0Yx4uSq0dhCrfL
C8J+sVi3eLR2q+xvLyTpYMUFv7nqqcFwicofgvshWk/JE9I782f3RzWTAOOym1HUU4Jcma2GvMpu
/4/R+Lk+6fcOk1d8zSgoL8LnyIrJ0XULqyFC77XCVnU2ZCbp6mwVdK6tZHyftfA2JiXxi+dOoo7Y
xgyFjBJNhXHfVvOPJKJZHDTINa8MlkEDw/qnM4WO3esfWYxktiCVfQOhhfMTodmYrW3ygdFF3HVW
ii1eaDS6ffl5VzSI2LL+WrykJ5RFdpR9o8KJE+ze2RA0Uw2wlN00i1iKOuTwA2ShGP/nWC2K2F2d
ZevTXmtvX+tdle0+h8SFe3JQLO3RcuuZiTNj46ttLTaH7gwrdxkfVBoMh1OD9mrrZ5KdjOoy39Nt
njBNfT0ZNagyPmlL3lFQnif8fGpTeO92wdeCxRgT2eKh+sx7t4TX4r6rdqxiZ8IfZDVgKk6pmTSx
FBspeQLm2alBwE4BqqipKqp4UHUmzT5dBYAHvPNb+OfjF/w8xKOjF1I8uDTqhaOJcpBPaKfVUs5d
D1jJ9lBmf0FQtNoTqT3Jvnvt13sZIK/qf2YfjK6HaJ46/ZVdB3LkrHzsBbtkgVwQ/hcJUuda/wLS
qqnc7ioB3IprseOMHstFSoX/iPWhk/35GCm38qzhfQPToPld96cmWsB/t2gxnPKUgOXlsoVJ4Vj7
UblOyWxZDPBdSgIILxCQEW5u5aSPVxLr5ugVj72cMAQZ0ApcVHLK5oeHbZSyMxuoErzHeHABcJDS
9Xtl5ApYYIeDY0k1XfhhfgoFkhFX8X6d8pQU2UkhS04t+BN5vjur6z3fWu3p0b7nGQ7R7owE++m5
/CoQWHAA7VCykM8yqGJRib2+cT1pXNxc8+e4GtqQW1bFF4jQsf2r3Irx6sTObOzBBvRmtl1fn8DH
+8977FJkwt0vqK/3BEtxrdgjUqU7d/U7mdAAjA/QJOHFd9F6W2ecQ1+4lfrlsjzniKJv1pR32lNJ
BeGq7WViSZobUD5QGU+iVKl2mQRKDxHuvICsba30oqpTLiIykZeaM6bkpW88A+r3jjPhTLEAdC7O
wLrzJvSabFcnjL0Q0jOHsU8xU+0yc0bd6+5/uMKehfBvMp6QgucVQBDj7YbqZibZbl2bfMBH+qxD
HOEZ6HOOuaOhJgpTezH3qBiaE0GO1QG1F2uZVxSE9INVa26o33hd/uzTxYwiKrPkgTPpieU3ZjSQ
+1UP2RFySgKPDNdMyb0dNpnLTr1P6W1yI+7aIAuGZKmNUnNQaoOZ74TZZZkO7CVwXs/DTE22sCnC
oByp6bbTPIjrlTgZiCfCPizPgKBamK75bFeT/5BlToHpYvSS93LiV7zZdOvpPjFM1P23vRgz++St
xbBdyIr6a3FFhNhV8m2+B3E+AYs32uYlDiwvSTQlp41IQLzvnhY34tM1BT20GbMIINAHFsM+hGwY
AG2XWYZ2V0vMj6QH65y8LKPjWnhYjFq8eKsv8KBHxXFHBi8xnbiZlLm+w8238UnipHQh6XsUTkUG
B8J+Pc2r6k3yQKY07ko41PxTArHR6LpR/+ZcLm/DkIT+fK2iF01m4xC3tOpEMb7MGyJvpQglvO3U
jXEf6PG5OVUhdDuWXq4jH18GoOyi6Ld+Pivc8hoZoWiCOkATypdtFRfZbGmLO/363lMknQm6beRK
BDxjfFyokp2It6Y99msIhC/BBY8YhNBGK97ESPFAcJgAUBYunxLtpTEeYyYmXpzZfkEvEjd1rW2n
jhe+sTV9BCSn6DvO6lkquUuHTbNAXTwEReWtiz2sK/OMRHVwYETa6j9rTGx9x0CUUngT5DsU4dGN
DVu4hHAqBFt1cfl37F1C13JJhsueOWRArQXUni7wZEVM4TvQSoJnmWRnJJkLJPRlS/boZnTCk5ZI
pE/JSkGA9FC+XSALFgob8SkiRW9Ut1zcNaQHSTqrbZ2O5mMdCj/g1zsJys6IFo9mIS6s0FyUO/Ix
memxXn86SEaJzRq0Yyxm5uMNKarxWqsFr2ApWghahtjTaaLTM9mbHhSeSJqDFZn3TEGuTfJKSa5H
iGvCA7EUlJZCBI5kvFw0WsxmNp6bIqHQdT5XE/oCPcOv/DaZVA1HzAfilLVhR6nXo1sO1Ix5QniM
daWkNIcqEMihFKzSTn0JgOvXxRF4/ij8kepoitLMR1AqbZa8y6W2GhKHtVfCvAwFJM/nGrIy/6Z7
nhs89egdvN/d8QSo03PSm4jOKIkHvKWwaU0ucTgJ0vhECkuXK+08r5vx3VEtFofhhsKKZgDA/GdV
lJAZ5uCMrO2ghHCDciiqpAkDWXEkhZN7YsOosrR8PGaaMwFvQ0tOSo5lx0XQAjqkyiEa9kUc+B6V
7DrMi2fUm3oBDBbosYGxgnvflh3cGhYq913RJkExLlDWzxM7mSFkzb72K2Qu7KbzXdtRph845Emm
CkC0Z1ADeZFPMcXp/Hz+r+VBNxnSuDy0mnBHYXbN36mkXKn+oSAq/OgutArJfLlrzCjfRcSjLsg0
fyS2ZKNTKbw/WaZfPGPm/V7ZxQtDYdvi15H5RrcLQOYkwKVVYwN5VmOZDEM35+vu/ngmlSMAMHIA
bSu01azclTVYa/PtUMY/SP/jdRNLJlySBW4tE8ehShtvzjCL5bBF7ZQU/e+AcnSsufgNNm1OJ22A
+P7iDtoU73lMzl6QqVEJVdi6nzU0T7mVugSOtaTTlUeR8s9IEKGjNRhAVDPeYvfUYNPkbBJ3j898
VOmHRTi1wjgWsakH8KBgvhgpfY/0azgb6fZK7cN7CTkCbHU+dPX/aksGEuv5hR9RmVRTHnFY055h
rmb9aVRdByrB5G7zlIpjFbFUmMyBkA0SDArfGcvW/otG0qmDsuZTVd4nPEB/lbBEclOaL7HC2NPu
mo6gCY921CIALn9kB+4uERBrTYoZ5K64s5CtyhYFP4SFEaUCQ6cK7EwJd6FsLWhwunt0YwyAbz1f
qCWo+J9bpUoIHoEK5voehJW+r8ATGkTeswucWsF4wmmjiTar8U/dJCI3msKfJGnZ2tpUOJYKSvam
+coFkDB7443IpXtvrapQ+g0anPgrZEe8AfqWiy5uARAQsTsWnrecYe2k7aBBM1ZyqPny9HXESpP0
Crd6fPtfN46u2oL7/VdEJIasQhtgCs3saBh19vLiZqLKeHFQju3PtFgd748hhSyXN5B7KYD1EZzw
oMvkZQsKJjLPn/5MxK+hKMrak68FgbhtVqXD7leV7bAtFVOuLodRaZtdQHJx2PLx8pkvhOOBB2mX
DBtFbPn9glgtS/YSx9LtGWYkAXQnx3NHpqMG1F7cIuI6ls3JsqD8RSyQm+vZ35pjINSGcqfkE16A
HeK/szjTcr7aBHkSYKDRS+3SB4Lw1/BHdEm7vg1ydWfsXrNlNoCtvWhH0zPSvxBUwlXG90v7EbMr
fESv5TYDM5pBGf3aKPsbnAgQzZwnQi7gdEbTNs8xcKZgw27NpmBVHTRUxsdyCHXFr4Q7E8RNKh+U
D0mLQ0CmU7hLV6LdmGvlfMKwJ0Jt6ePYxQQMivzdDtwrl11j8/TPSxxSEmcwRfcPG7JfXdDkY0HF
ixtQX6w24n8pqy7xiz+DHz8jTEeQCpFXSkORd6e8lnoJkQ6Ji8PuxESKlNQMX5qopURNihYp4XH3
qJsUOcXZcf3UKvt/n9pG08a1g78+PHkzF/WNtrGgDxMG2UeJTtNuohQZiYYqHy0IpZ8/75wvhTIV
9nSL2aLj2E+fjOMDJAhqzSD//eCjeDoMm6OeNJ0Syy7YB9F7IfLsCmZu/Xt1RGt/EW4USTbXGZu7
Pcp6XOTTA1GL+3oHVaew+iIrFT10U5SwJYS+bE0O+7l0RTomb1nIRg7ay0jsHpv3HD80KNi8jADF
WghUGxuEprxKH0vzkgcRdTlBY6rxaH9cI8iHpxa+jrciMl1V6ybV2DCafBZLIwH0/s4IkA8HaM7X
I6ldjxUispTG7sdF3SpQx0sJlNrf+z6GFcWLNO6171n+NeOvtlN53pJ0GRDIv9q0g7YZhWZWAfY4
7gARVuIihv9Rfzf9IiJb8J17Y8dTbjdes27mvgptRNqi0/PYZoYrA9wUEY8kVpCUPAJpaGPYI+Om
Tu1ciAWlflHfsHXjU4JyhxEtCbx44jaBlMDSbW03WD+6az/fr/GIlt/j20W7AzmzmisEJyhScrO3
i9MY6me9v/7NI7r3kJ3NnDGgGvBXUaqTjMi4aUWo1XkBoAGxTPxN4L0OzP8WToziAoZLjV2gs+nR
lhMv5X/tADulCnOyb20DFY7FlGfUqfZXIGgBQWVmwG92H8+nmuvMOvAmKU8ySdtWVp0GdaDTYOBb
c6/dMeW+M9GT641dXUS2VANTEHy1yW0wHAIwdMy0w39DK3cpnoQrYjtSQxTREc/Zgj4Bi7aACkL6
ePG52LRGyX7pCGXB6fiHDDd1RZ63QI4T2BzYjfCgDrqRDHTLDhlttj6f2bL44TYIEKLNz0YQ3rc3
LUO+2bkoAbOw13e97Odsdv6jPzqmPTTDzp6vOXHsVr5ojZGPvAKepGfUM+lyfUDqiZlTCkX7/26k
GgUCbhFRVgSaV8dlnvIwnQmK+Ad6/4+RDzQReVKrNkQS6bmj8AVic7zznrLK+AsZjFEo/ubDEfzO
1dpV9LAeAUjvjGjumc3vQimvz5pEZSLiNZ8Gz6VIK/8dVRj4gh4h7kh0QWjkmovQbACicb3m+RUJ
tPlh9v+wtNSI6ZQtyKKGEp7X58LbZ2XUOiAnWjVfKdQ/t08txPyepY1yMQJLyEu2POqJ7pkVkwkJ
ADtNmhqda8xzMHwmjld6eq5IdH+HH/bLsHnWCcLM5DX+aZGPFY24ztmJp8WuLMukCvssVXPXN43o
6RO+oDJ86rdIqrq4Q3Pwf962uDaRYkcxzN5Kucnrtm8QIun1F7fAvpRW+Knz4aGHsl+9sXrhNrHH
MysBKH1/nHxZkl/cN5A8TAyzKbZsVecsfokC4UW0GpsO3SU3QD9nWSObxtKSEYOyCDMtNSNa1y8m
TfXN8OSDcTjEZs2fJo8Tv3XnxLAIJ9QL0AGsEmi7S0wClv6dm61afolbznX6aV1dy1GEC8QFoX26
+G/PcoYr+YKDKAch7Wl/o2bzH7mw/nbUNaJcNivEwCjsJN+BQT3FxHUgRe83naohNJupS0EXiTXf
2mRDs74td+ysOGddKAvksJrMyNWdVZQmFOQ1eR634R5QhlbLLFcVfqGiLW3wZB49Fx0LVbmVXLQc
pwZhznipCTNv+f53gCcMKBMM6e0kJHIr5uD7UlEv2pNzpdV4iuhePoqiMXB9zJV7NEEm3GyNLEln
50gt06c1Zr1oPeGMd1QnNH64RC+6mKxbCWHJG6mJzSMYV5PbanrBhht3Nihf+8GquAjh90qwIyYA
uzxYteKKaL0+LiKCIdJZe6exDaLuShRbG+00DDfB1oB6UZJEx/+omdF1QSAOZ6hQJLOLFAnN9GQq
/SpAQZRe/hvms0nq+tuU9gcc6OY/JpFmCMWj1+g0FQ1+G4qN/qYDYhHlbvait9kSTVEIbBLNpYME
KNB58S4KNQ7Ssm7QiE5B1edZ+oKMdzd9zt5ZjmISsXht73ECRyz4ZK56g+V90ZbbfV2JUsrlhQxX
R52RI/jRasIvwADD5OcLXzNxR/JRFL45gjW+NA0n8IggmHAROZN1o25Y0mO/rpy0ShhEjqmaP4sn
fKZZdclbU7sOpU7RvCbGnhRn2R+T6ENcfNEHTaR5p8odR7+hsyggCbELMdbD7w6zvCJodObLtQy4
82uC2oNjn7bvNYYDOYVsTgPB6RdqJSE0Iqtmhr42EMLbOoppG+iLsgwUGQXtnqmxcDC57Fk7pDUI
RLEECEsg7oNQwvSrVaxElcolRaRUJVMR60UoaOS0yR7x6gb7sTvZjws8cZ7IAzQRxe38aSgV+/JB
d0KghQ3zrHQ2FNzbqQmBandGEh2GTVD8uvVyPR078zP28H7Gy8xK/ExMrrnjUh2jlUq2GIb//QMG
y/AqnaMfMvYvTGV1n6lAv5Rstb6ikGpBG/d1QFRX4mauTK+FCm0Oz9V/g5fjLq9qA85rYGvILCIh
KZfSS83g5BjqjuMDue8Y+FXINwFUWAG7M8yRGSJ8QFYvrGIUeiL2Xf0X18h+/MezP4eg9sMokU6K
esk/dfzkiW7rOXMx7YQX9Wcg5a4TfABBrQzaA6erVQ73E6kHRfi/ZRHTsImq4TjGfCDHgpglya1c
sKSBLqryCWHecPWmg187b3LaF7+BuNighOs0W4du4LnW2zM5wRuJYoXHO7bBJmlh+qUw+2aJMom3
4HOOCyKYMwy8B4HHxnZWtbwMN9Gwh0pbXInbuDQQtfqX59RGf0Y2wOk0dQXNdQKGE8npoXPwaecQ
sLUywYPA42IdVHZLBg+wbRtz+hjL/GeoiPRQWgksVwHWLVe1PGHkpuVMd150Uq1UepUun9YSo/Tr
eUfXM31PtpDwf+xvsENgE+ZhsYbJvopNkZ+6njI4PdoOQZSWCcE0yokdZsWzCgyCgQDeAelAMGYr
OtUqxRNABzRnQlNPAF5WEuMCIeDZ212ZB4v3KD82D6Tvt19YUDFHCo0z6Egan1PMYM4bsp3+5hbP
0GGimQ/RtV3tqxMlFldW55j1Km5tJZkUn2XsQyuJIt9NEpFFZXBFUgh6BF3RIYeNuTt7nyJx3Lcf
rfNqVEzZcPBciHwfVEHjGhpx2QZnDQeoxmCiB1xg9cKgDRoj+MHZwtA2IkOS9YxPOugK51jXNpeN
pZRPiedAC7hpNvHbdFssL25Ykfg7IuzMH8FBdx4zvzYtdMveffhbjXMShZBwB8nYqk1o/2yArhgD
DgnxIQFuTPLTitEH2T4+YdaStQoymOGcheZN3vZbA4PPKVB6xCvku7vfWBFwIWi2Pi4Q5voWH6OE
R1Azlz9nkmEBfoQzwny7bE+w1IL4JZi3TXOYGftva9F01jnhpe1EXRItacuRZqiGa8FV3mGx1Q7G
loe3TuER2LZl9QfVY17PL/dwhNDnhzIIyGfoN3H0zC0owKrWUDy8/wwKkKyBM5GAXhlAF+fq9x3R
JB9bKCcqixm1A6ckpagJtLLAxE4avOMJ3I2b6wfmXyUO4bDW368AjXYQ73G+Nie1/xEb/ArcrI1R
JTmmsRgkjtn1ZmeAqxO47+Yv8oIYz+VtzWLvqcmNMKEPGkissyV+C+x/xqgN7XVCTySKCJ5H40UC
ljmyRgAxtEjQJVrGGUMPLbeRNdtcuqBYTVTtEquQgdwqyHYIXgsEhP9XjFVaiKTLWx6ciqQmbftr
LfyYyb0JkhQ7NjlGFnoUGEMk3OMwzGIcUA0PRTqe0lyTORBvXhrhltuQIqDoQkpSfqJfNumqtPkB
99KYRcivN//bwBkRUUjAOHqGgkMjyUWVVmJirGiq7dua2tcs2a57brMygDA6Ltl5YPU+kiBaFFf7
BaM91cYFIEjXpKg6lhvHZ7IbXX97Mnckjn1kzfmR0R3O/M2aoTQ4JFP4zig7Vkph0+9xvo8r4/XW
xy75SHdozAWmNfyCqS81WWzKiY5zXhApG/PeTN5YTa8zvHJMF5xQect8Y0za1/5ZXY0RVcSDwpip
g80eGE1Fxm2n0uXjjBYX+gMOHAz732AYnRoQ/rSXKxr1gEKLe+SH9iJ7MMnj228QYDw9otymbw7L
LZOprZwMztt8aO3Sj9U9U3Z0Y2qhAOiAtT/a/+iTwgEGDGbC/9M27YgknBVpGlPg6AQfheI3Y9nC
gzYp8/HqsRoBzw0S2X6N2S9sd78RaH65bPqtXEfyyYuNDOLGjA1NzJZ4vCwN4+dZzavpreo01CI5
qOg1g6F8vIvgh9UJb84S43NFSdXUexBgXAjADmoPzyRLr3B3lt5tL2pvsS+Evw/zunwggKiSdpJ+
8GlrVK6rcgVkThC4cutWiVoi4JtxwJQttRdhMpIIxusQxGagF9kP1+8T7X1yWcDDBAt3clUjroyX
O/r6V5RoVEFeKManxsdXFVYjy9O1q//+p55KovMdrqACifcWly6JMp0aHHcN/sPy08d9yfnsBBI+
SUjRspNEGbkZobq5y8jGCXBg3/18XYuyE69YOdCjfMa1jxGhyJYwpBEo3+jc4Q5E6NUC4qTnWdOc
2VcDWHy1rWA2quMF9ypAexrdGAiBnnAAjxmDSH080jKGyh8PpWChApYVSLaCx1MPyNM8WpHRTcxx
J5XGlzlOTzNgIQsOBOgAyHlsPlIeMqX8YQz76QaWApRJxRpWBuawm43RnCmHWAbkm0C8H4tEPjDQ
38ko7wdzTgNMv7P44CsngF1ktthy2wq6SSoa+6UxXlgXGzExe3mc5Ai5gasqxRyM3apFHfRgwGRy
EYLX1FgGNZTfagBGoW88XWKX+WCBfDPhdMGXO3z4hdSahrIg65ajZHIIy47It1tWNLrr3ECoQv5O
C2CJnWFlSGv45EXsZau8aCI9ZeH7ewwyZj5Y9eUKZu/4p6lFwlrS53uVfJUh/FbH43zTCJXg271+
efzXY9TDOgDt7NXzPDhHbzkQ4/wRS3geB+VutFnBHDFfn+OG4WxDa3XZnvMNZTrNO0eGj6gxJ/+y
cbxgxE8Q6QuyL0+mtaQO5lPt5bl0qDbjKh/tcM4I7vTz4Ja/E0jA48Diu/UOobF3POW0fli4R7Xm
pVVJrjnYC2epikTeeHNiU7vCqjAyxYipHG0oxFL9jKFz9cUdyJ0IzXMIujSP5z3xbu6TY04LYe4R
diJPcVGbrzlnDgTCEwVkpaMrb33M5e8nTUgLnCj7FHJgLCHMNTN7I0h0haUshCQRPQGLaeNVzu/w
OOSeBpk5mJx8VG8ASySVdf4VRlXSqDwAAKzd7Wk1T7QSOcQYyEmZVOuxhjppxsCfVrEDIud0Ibai
WQSbLUdI0CO6PSS1pIdpB6NJ7dqNr8bzZAj0svxYXW+5Ao4Gzdcc2BAaMDDXiTpnZDRzUuysg/Ss
l7GAp9r3NxokncKZ6mhbElOukKYuLVQG4dfRIcnSBHg49YSQcubco/6LQyejDD3ncRFd13DEwkDh
U4SJtWEZxS9oxi8t8zimnzcFYfLEFuqYXs2tybrY0wjiw6DdWVrReW57LenIXrJtKp5DsEw/D8NA
YxYPlwuOgujVRwLljuPhVWRST9lheSstVvFQrf/BNRl40X+e3MCt1ev9bboe/9zOnKSqVWv9H7R4
78atwSZvkofs1wILihOCg3/k/OQFeeFQRDlUWPEM4iuvkEYSJgXfPCChUHwsESpereEZb1CCD+rY
d0tEjYW5N5YYHqd20nz57PRKc8nCwo3xzjyOAN8zL5n+HKnfa0H+pDljSxX7gellVTKIN3qPoXu5
vanzBXD+S01JYIC/mken1wVj8sbXUXlYpro4LVhu/zDYpJALOGMK/aWe3kNpQcDK5L7PqiICSogA
82xKt6i7kL/x3GKwJmrxAzZIqo0if9RCntuPqTNSl/lcxFuk1By2CHldghCeUH+eITPX4yfFZSv4
A5OtVcWXW35596itHR6tJsTAb6ho75AQ8CGqQNNml9touRvAVSlYDN6jFb6YA4DUY0aYPl/72b7x
DPSi+lA19gU9C7eK7LnlqrPhkPyCCBmVxu03WXVHhiA+zJNiKzeIrmaQ4MOy719K5FbiUe809fMZ
LVDwKmqdLfxUNkuFmLx3xF/qRuzINzrCz2NNauCICuhd9FI7ai8bjYtXO8AMQm87x16UXTBoUE3H
o1iCXUa0y695A+/tMKAOkIarnpVsVXn6zxa+qrg7bZj5icRCO9rnNa25sF9UTmqSZMqERJYnE0sP
H5Lw+4+VpSal287w6APdi3lkl8JvnAQmDr1SAdE6d2XFs1eLWD7oNmXkwHds7BewQPhfiWH0ELgr
zLccjp9zx/sYhtPxRWpllH7G3UDS+YXGiIX+pg8O4jFJuurDdBMqDT2QUfRKnO6NIif5ircM4VPS
lVQpCEWtwhKUqDOzrFkWip3gzYbWj2N3qfkbB8cxd3/RKjK2KJzJl0oJXXwN/40wi8yt0ebVhCpk
mXrHNLL16Krg+k8OkTpd+eJJhxFzb1quOgRkBqnO950LJNVa7ZWtYJ1Byn0h3NYwFguoTNaoEFh/
CyXaOGdJlNog3Zh2gMUYaGCW9mYvyXbrY1VwxPSiQnT7Ia0I4lI2pF4d223t4Ftrm4N9Q4iNIubB
6dUVS4tJMkv635NaQWVTOZfRI1210+eAgZ/O0HdAQuE3EuZFb/BoIFy21SANTcuRhinGiCCyrLlR
cRLeNeqX2yKRzrQ/wum9tpJRV3oWZcZeSQgrDxJ5eIaIWnx/fW3m14mFvMw+A5lm3h6t+Z4zDLfY
h6kuykBTALnI0xwcItIbxjnGvSuaa0KyLz17sNVUiXbhpCPrQR7bLBQUuYbvNpeuuILTrmdg+6L0
zY0rc+RZSE7R0Vk/KLZOR/8+mRxXF+a4QpbA6CimEkuutFFnVy1gbR+MqfO7ut0sD73BGFd5xRyV
HO11oGexQp1oKeIpsDVrNacgG7YtvxYLxV8NZZ0cj/Ro2HDhbvLFb7VftxTP4M7cHp75NCBjUgy1
3j1xaHjtiez3MGPmfM0Xu2Vm7wtXnCbezhDYihxPUtbfQsz73PJqS+mdtsYXEn0/rrgN6oOHFz7j
RPk1ABijMhLq+f3NRx28JrgB88MTrJRdhqIcITAjr/PV5ouzNFZcLaop3nljCMMq+8exEIKLWrBN
QGS0aZO8moEfTwU6TtJmMtw+UigQzaF6VtpuHNXZE1dbrGfk7DnvQoJ+gglVfeMsplO36pVcUNhm
tJH3e2ZStEQvPyM3ML1R+HVoaakTdamaRXUL8re/s1JCRUwFUUqaHwo7SZ6zgH66+6SASZvUPahX
QwPPg7ayxnmHY9t86l1xeaAQIzvZ7kMpqP55CV/GvWUP5nIFUS5n08jTMydP6m9m9vGZ7PMorri6
3YtI1kSKN3zNyk9qP+gYEnwusVN6QaJT5+WgV27W6+OCHAHPXRxFtfGNKAjfkHlHk3a6ZgvHoeoC
yJ+xq00R8aD8TJ6AsTtbDJP0Rfk3Baw6C1f+WI4XvZHOJs97DFKyd4drs9OzXjXajEHlhxEdGu1o
3Tqc2qQV4VcppuNZgJX3ydbGcDWNl0xndB78GjdU72KaMyMFlWOCJDpDZdsmHwVLUJYhVpAQ4G6g
6hJQjIQkb0VQah/CtJSQw4S+OPC4XD6qdWcBQmRtCCpyd0BksKtQ7f5i6ZzpI0TVCOsggyzCeHfY
farRtrdjBjlB/4U6o1WozmZS3t5zN3ao1PC9/yL1xnV+aShD32ArCY6OaiiOAY7YGS5A0rYngArS
MDommCmv5kJYjLX0wQeBATizFRM26bl6WXi+pVSc+NtV5jSwa9rEjnAbbc6coLvVyJkPMcit/UKm
2XPEoM5xcPM3j5VuakYAcHLpeQud5FuzF0vOEr1p1J2PQXG/rx6ke2ddBuwJ5mmEgqiNwKroRFfO
4Y/vhC5LyHYp1Pj0HA78j0F+22NE5qnUI9xVcNRpf9ToaWQaXlQLeHTfBO4IXYTfjAQ6+mMmVlo0
DxK6pfELSsfPMLK22HFJvIHhCpb6Fwn1p62IyaRJ344feEfURlD1aY+vljkfOUIiAWpJOfEfH9jq
KiR5pmlSC3zqWU7aQmipmiu1uyLp2Ix1+LX8bSYBDiLdXh7VHPcqZS3/Y1VNSfFCinbp52K9ctQB
r0ocIVAQfyKHqxasrrsngeXPlD7j4iHLzw3z14hhi1BTX3ewxl8ppUYFVT8E1dLjCXAeKTXj3Pbe
rCz9JtYKn6UOYLoryyNFxQTC3zj19DERQdTSv5A9KnLlPHLAuLqSiUJg7e3227t0urDuzHJuv/CL
WdlLpK420JBoNfAgEzRIgscq58iCn0fMBxegyngwG3bhP1pLSsYiArJZKLMB6dKLoZr8IYxTB/mZ
Ng/S117vrWJ44A6I5GgWdcqRWxenTF+dRZFylKrvthMdIIgohO1plRfM1sfsJ3lFCcbVBarPvN7J
PQFT395Y5SYLM7CIeGe1vAa26MKhnJ+3Pp880hdv9M5S1wKeY+s67nXbJvonXMkPpJdlTRmx4dED
nS/EU3eLKQJ338hm2FDcJpKscY88x7ItLY44/URG3n0zYdDran6rcKPvSBst3F6qGp48mjiHV3jA
xKb7KVtWb2y6V9E+hBY5Vh+N9EhiSME5srSvnoV+M4UWY8k9imej0m4MGA0Mhsj+eyGl7pOrnF8r
z+ReEfWrFkjEAxwCS1qURTvjMvMnYm3eCJjT43YcjCH1Y7nrG++b1s14QJEuhVNUsPlI6xXGxGGi
JY7jHZDNhsT6bjbaz+9b7c4P163TqfUT19WFa/o/gkCJRx7PBbj6tlgp2K4qYAr2+r1yFqQxhddq
8f7pkq2nZPJ2pG5bjLiCeqpVzhn+eKAxhm7J3d2jPF67q+MWnC8YxLfinqiI3gaP7rpain1FZPx0
Nj0IR3Mratb7SUYSxxK2Esn9Oqpc/Esx/dBTDFSTkryRJvuCfhaJQBo77HUbjfPYxLsJDrX6Qh3D
x9+gmFZoHzCT6+NQnTweMj2jE5ueu9NCCVHRRE9FzvYQBBmzv7O3KVxo/TzrBwxmw3eqVrEzdMj6
JSzmHL4pE2/ToCxtqG0tcTwYPXMCSG+xomnoXTCanTmFfB9SR5ruiIP4Qs4AAOxeDHS47J5/DEX8
mDSRgBnVfOUdXw4HXCmMhao4p08EWrwEzq2kZlWITCGkpyPutXINbJNRK9bD8y3v4r8LOZE+97cL
j4haweaR041mptFJTviqT0bc4e3nY5rz/WwUikISGSyQHlvc5Pnqvo4kCFjdT2Zmzt0rKdyEDRL0
T+39OHNIWGn+UzXgySgPjXOL5Qj89GqJyIG7EtpZhhwRe72zDgijdEljnnTQKhlZfsmNzdI9p3hH
bSIlexfDF+rGfLobBC6jEznf1mtFf3k/hMEhhwngQsvRI1P2/jEgWOJI+1Bs6FiFETkFtYdEk16o
7E/qkoWyGl8ZhgyPpNzghzDZNHwxfR7330vDfmUYFRxRTyKNX9FRbsLMVL3eidG90NJjyQ1xG8/i
t8wC6bWrjC9PULH/GiWXOBDGhzn1/5IKflqeqWE+Gnw+XCymvicp4FfL58OfMH01VcJyAk7Gd3F7
niyK75Z9MJL58vYu286PpRLBvJwQwk4p4YZhf3uYiNtPggr60fYZ6Eov1/41YGNDjpueiusLR+F7
aWwemuf38K5n8bFSVUt6tV1y+8cewIf8e1OWeB0FTCA7iW77DELJkkpGVVQJl2vHABwXTC58Gps6
JElinjcbQPAW8o/vqdBkYv5o+rjyM/WsgBeunj8rmdGFFZYHmPxTqmL0K/UKw/QaBReIup0mfpz6
9JYTubrkS1YUF/ZM7HxkJ6UXw/ZPypgwyVL2jCUE3JqboIxtybRsljtIV7Q/HWW3GCdJfZynfFeu
+T3bdbWumEb0Eo1eEXbOqisTfZ1auEDEnZEmGjewUKKTfD7wYdYDuFGpa+UkD/MZhXfJv/7ym6N1
V9UCen+J6d8GRnKacC7ogtRqz7HmLJeyRMxFxoxKK3u2Avk1vdV4pZvn0pg2ULXDG2lMgZuIsCPS
f5+cFT1u+kpBShyV/JywVhdbYaeeGHrs2SokIxqcHUjb8ApKuYw4P6G4GNETSYRdkumfvMT+1Q2v
eMNPwq9PqkbSzi5+uvgaX65Cka5kKRstzFfUP6Og8FzWAUjod2wwTY3zAxtT0I4iP40IUStfv8T/
15ksHoK7BkjfEFB1a1qVlyvW7aHmBZtICBIQp2H0fnoh9VWauDwSUsL0DonZP+sFHOK7RrrKbgT/
9/mSPIIOAfwImgGu8s4R/JC2UuiE+s/+r/sGvu51YYEVZAnJvVpmI6/RkQBwezq8apvDYiY3qXwy
BrhnNmXAraA1K0/2LFUQp5zRR4is7GvpNwxt1RppFXyIu6GxgWXnIMRmkqBmcNeYACkGGv7OI74f
h1RKFgM3y+jMRDPgs6wEhvbmWVYpkwWwAfTL+t3YelSTvZCTrE+Y0DWtZRxsbCRY/7PU5xGe66d0
X3JqhPEL1GCUtQf4RBFqY5sEoZZi58MlwD15p7bvhDWSVGC7bR9Z5zQ3H3fSIE9fgz88BjHKVQh0
A2xd4IR4a+PWS7gG+AQGrYHpB4I2fzJvVavrGRVsborkTeXbSy7PCyINcc8I34yrgcheNtwjLRvo
RrbztAhNu3Y0OefSuSRRduWLUjmpkb3GJ6uOD+RaZSz3eArV7AlpwK5A5WllPFhm/k3/uZ/qaptw
vs8HbEBYrcF8g4svbRxVxi9JpxDXMfnpUPbkSYLOc+kFLgFZxN4ULky3PJE7kA4l+Ld2WyYYYDQZ
qDrZpe/OVIi2Ls8yepAlXIQWY5Xf8vZi4QnkoR0vEWhdiPHioelwtzKmcPNRV3t17TUOyQ4AMKAC
aoMZTYqv5jI5JAkYQO2nh/MEmGWyVKvgN75tcsvhHaBjESXKNP+803+PxcoxX4A096OQDb048m51
J1H1xAi/qvMLa8jGZXKdbBUqNbmFxwZxylss8foyqqEt8s9J9B0jqQY2VoAdBM8hPNbYrh989qll
i3aZhZqWL72q7Nk0mfjdWZkIwMy6Ric5mUTasQ031/OKQs11GWFfVAti9kCDB7ZLprD1obFFn7Y8
HihCaGAo3fOLoh2tvf8JAC3lB9fq4h+FPA18TUpsaNxMrscJQqkEka8MOzOWcs5uGmjbKy7SWEgF
sP1Ib2FBOuD264lc7sMLRf6MRuoE5S2GiAyP+xUli/ViUGF3Fw9t90ud/5l+A1pg9/lqTgrrmQAe
lfzd72SdTmwV1f2nTeyZgmOTLZ+kU82+Rjmnb/tng8+OMsgnuTGhDi5b5kleaDAPOipg/7+W1qlq
ZJnv6H7OdgFU2nvvB7UA317HnzN957IrOrwnAHxOeJs8JLRID8eZFrOnpV4dFjozRrt52DPOPte1
dRN2P/jzVcLxobovm9Kr5iIjWepRhSYi5FXh3OoB4k0Or2Qy2YA9QINrpMnr/ThqtFrO+NEQS3qC
Y4wlOr1i4lsjndaarJM5/ulk94+iTw6jJWMtX3uGvHFkLzndQB+XUFpD3mD3gCtKLLCR4cpwjb8x
JF2IuNQkelDiOe1cnXGDJCnOZfkHbTG0k6bLHOT1PzAyex/pK43KHItyhHKguDVoL+zBpry1Zpff
TDprk2K2Hpnl4vVSs8wpT9hg3pvHmAhRPbIi3pZa8YbNTgBx99G8tmx59t1Ee2bPmdnU5KOrdRel
YKWUZ1zq+ikemC4Q092mi3Z/MYZgCxiwMC85TXZkrrWNwISdgjKfDvNkvWlZuhXR8SdKTVwvlHUN
zadUMFArdhYRoYI/Gq9mYiAPLRKyikFvSloaprh4TvilyfSt80yno/RPLlCUubWI3a5jKxHW9+Ga
/PSaTyXtvbs6Vaf1iFftT5zBdtWheNicEQkwOPcB7KJFkQZDiz08SZeNzGktjg+/LYSg+oJYhGXI
e1htbwaY6cC6srmxkEEJ6R3jkehtf90uR/5fDccAEJ4u1cHGq4YPuHlFZLfyJZ4gz3Gp0Dro7jcK
FomHcJGfZ/klgeM93YIJN/egb5Dgqeqow+lHLwn+SA7GZp9decITlVOuP+NWdaOL+RNgtq/Fv9YK
HngN6v99E/sszTsRELRyKdKQKWjp+rG/o8jyQ/c8cRTotEZuThka3nRjQg76kRT09KnMUY3gD50u
k+CiA92rUEHn8XppnN4bjsDshJw/VCmooQsusJoQP2NKv8XTHSctqDO7CkwijkkbJiu7b0abq2n3
wOzjly9riVyWdfmKmvxAAM0SpiPzyysw+hmro+kdObcb3h+4E2v3IPxl/FtaT54VlVx6GeUe7RUZ
XmAD1LLCeqS3l2hdkUQ8MOwdcp0QOZZNnETvM89BVQAOEIfaivgpSEeWnFcpiqWc72Pa8W/AQObw
3Xgt//lzTOWXkZPFhiyHlzeaZd870hcrPmAausyjjcwC0AMm3/5Y/7EFSvorv0DVpIfsKqoERq5b
0mLpAUB4ZGPSD7yhE8Pba3nvp65IYsLBiWMoRTL6BCN3RqcDh+H8fEd9ubn2VcyfrE5w+2aPe66j
Il4i/wvmeub6dgNiKSI+JmsKruEqgRKSTpZpjKmCpvgnc9JwXuZrokPAsUPSkiM5MuMydc6TLC7e
q4JWiEBQ/msel4QIpRSP8UyUAORfVCNjNmH8f89/ILiim9AHGasrxnGRaWiYkuGPA9IK4Sht33UQ
II7PfCSS41HchWCVtiyi7QA1iohKbDh9lFyWkwcvMMbtUKnm5dTdUMxbuaaecNUz/7Xm3aG8QIEI
z+OLotDqR2V2tUCsaPiBmxpU0DSV3JOjpnj1TZA+uNdXJwUdGpukas4w4d2Jt36tPIRlkZ/CAjbz
KKGgDZB1j0lS6w8J4qpEI01mG1NF9XJj8uj80VkBY7rYahR8CTfcJgJZphYvijZQfwmgxVRTzzXJ
Q3G+pkWjAkeybphw993zC6SUawUaR8y1177NhapbBG3uqLKkf5mQT0lhgmqC0QRdZ7RmNP5efN9O
GVicwFriOM0BS1wVdGeeHvAIbNDCYwTnDT1wItXEAfEvTLoVng9SXtTwxGfrFB3MxBpT0sZjKA/p
V7F4Ib4aKA9irwPng8aC4R8DDSkqOqc+kmJBX5/5wrNQU48jsxiX+OHERC6prirJA+o91MPP1GEA
bv8a9/Ysg1FsOiaUvWVNJXX5onKUjNvaBOlyqJFGy42uHmPvkwIoBjUMK5+pG60xa+8U9ix/bfSL
H2HHmvBmcCInokN3jUZjwZlSVnkuCb5NDZhoYWQJuUA4Bd8J0O3A1Y9BtXKZ7FruX0ehsBxXOs6f
NCB4HCwjIgVIu25ZXOCZim2kqrixo6YlrAHtOUbM6+zFo0aYSUQWh8Pi5/rIxRY5VkwDz6AnK/kr
YIoP+CrIzJy1KVMI8P5CtarKiyzAOWu36Z6ZZHKY+QUHio2IBk/1+btGh8fk3gpEUm294PZI1Ins
k1kUjq3IFdmLv4zYFr7uROI63WK3SgV8SI5akDjJ3je+EJ1JBPmiOjhbPdEndN48gWz1d1MnjHXn
dAL/OAeXuzPGD+nvYBeqQjhbgAE0vF1BxJ46Suu+wOdtp/HDOvf0wUm5BgeAOVlt+QxsFWEYYbbJ
rrqf4vzZMNEU2e20eWxZQisZ+z03EbY8f557kzkEHCUl/7ND8+TfENo0G37J02o+FsGbJjT5P6Ri
IHgDkqrbkq9X/UAwMH6cKpREnnh00Vxk+JamgmldUij9W1DFk19ztqJdoOc48oLhyeKaXLuIXEF+
bYLt+6/rcb8KHKvQ51+fiHZfcXyWIdzcEbcoxibPS5W1uMCNhZUgXanLyFB6lFdLyK1zItadM/nh
hIPKZk3ND3/bBCk++PdOt6Mpvj0lH5WigbAs8qePui3a6zqhhQsiToUP3qg4A4Y9A7FhhtPhHyEr
JfrnDSRzNlguz0mmJOekOHP4/ayIGMWwycy96SmUzUfn68NG/dlDheQmSbqejVRoR/WSi+BdWVCh
XxMchhulzhxmQ7kHzwXu+KEXIAbSS0038u32RA5NEjw4nv9SEExu9nZSelAnKWwAugRkISz9crwc
H9U1d2OfgHT3yut7DSn+7CduwoAFq6p1wVo0dknjdsT+Y+/MCUXVLdJF+jYyTHFx9jgUbmNxjTHg
RTeTzjDq/02zSyzz5Im9FkUsmrO1SktJ89ZwJlgOhAAwtbgoklPoqUte8hXvk5g4SCfWSHDNSd8H
AADILotv3uRsNsQ+eKO+Ob2BVwJQ8R1Z84knoojLBXA7HjxZ1r77z76J7Jo+PpQZtABPOCTK4CEn
zhwML9bdSADyTRAH3bbEZJSxBPaR/3rupCHNVSq+os9mjGvbk4HyIqf54kL7bqxihcaZXAM6Ma8e
UILfGLqW06S36ZyrXUhZu4g+rmnwU5gDxr+LQ9fK9yb72gUopBRSyLnF+CquY8w+/iQTyfTqPq58
2NxaHPJmMU1KVSjv0neIk1IyjD8/WaOeZ7WRsqe989B0QfsCznPG2beNPmKVj0PCexVS+WiW4Ar1
w4uL3wDl/Xb8HjVPOPJ810GFTC3O1U9jc+AaTLgdpHxAq5bJWIUgxbxfZrdAdibvIQOZYfxbzIMW
gqJvQ/43Q0qlYzOprtxG8Gb25veAsgS437pmycFCJcAiGUM/WgifYf5E9IcUsF2HKBGjaU/bfpd7
R7PkVYSc2gPtxu1ZUrLVzg53R0SQpOC7fldfAzvC92W4iIBz7Sv/Hdz9NDN9XMH57GbkAsUWQNRy
gngOIzeQnzED5BxZasyO2xTxfpnDuX79iu1cTALHp9ZmI8/witfyPpA0TPEI528bHku9UUiUiCWh
8AQg7muFTydwaVpBfmz6C0xNp7mao0BxUyNSje7eTsCRIf/US+FGczM9v4LLAYi3AZrCsALtsue1
0LQy7jaQtkKFJOjZZK7yVdnMMAVtfWVidC78mRu++k+qjbGpb1dYrRExflBaVePNVJTBIIeF6Ntv
NApfGhvjm4ny3DlglKRsnWNnmmAbuZ5/8L95sW1n/LAkJJymDPr4ZyGmNBXoF3sNPtV+fjWKeqOI
HU3WW+E1oauC4PUmewVDA8rpaFjYwhVspFU10OlLxQ6jOuiZMK+GldtGfjg0D2D9FN6tuiz5Ty3F
BfyPdI7xjf9yKi37NSOa53H5NUy20YPvFXQ+BmSNXdEhDxnYbjAvY3C/qFXEZNO08+tIQ6hL6p+k
5fyKIjsyrBxY4KDIEgrT/i7oQEFb8YiT4k+FP8qfjpShxEGQV3KqMoPRfTexlNMzQ+tAXWrZ0/4d
8JEL2gN93O2DMlkxcr216Ir6n32hKNd3KfBvA0x53Z5VR08XrU4ZcS8MuQKpZ5ND4rbyg2wUBdNZ
t92d93YWYgEJHXxeZtj6imZV/SmwDL6DhSGzOa+vbqf9lhuPwzHNCRtst9Sn2l2QSkHuhf9Gbw/d
7EJt5Ngz8UxIgfEOrBq46WPP7hKops7aJrzXs8ZJ3+/TlH13+wxKZiayXmMNufxMEN2wYqx2SAkD
VF5rmP1bUvMyFaHB8fFN47wZoNWY1rZ3TJ+HKcND8a3riLNdy9dTbJ0T/0m+6kvk0Q88EsZmblG0
7lw/J1SPxcm0gPL7Ptu8ykfjVYiShCh3Wqmop8oTXreIlop4+9vdCoQZ22xsUP71x53kBCXTtwrn
bQZu0gX5ANKHz8N36r+Pc6Z6JgHONFkSJ5EoJrcRO9sa8aQOjtGHu6O5crkfC3vui6noWov8TZGR
byk8jId7F8DV06ubziOOmNJ7F2Fd5L5m4f6KS0iG3zxtxIx2XDtjCfj5TUDN8CNFtNmuOPCvyada
/QRXsReMHM9LtLfebYuza92PhNW4aJcMAYZmVX3xMwkxymAR7TQQMPydFVZsI+Mkdf688ZarlGoe
jFie2O01x4OFs0c9hFAHsclFCM9zBOa7QH9J8/L3PYPuUrpiU/GuSSxqbTRPAVaEpoII4bzYPoIL
DXLubGyswa0zTQ2+I3ieXi6t0Lv2PFx5HVZJNQSCDWbsTPZ+qbfALCATENhNrojmta0+262VX4Mm
012oHYNxcyHktdjh5eCxtk2pq0/inOOfVA0JYDZJ9XGoNcxsxhUOU+im+3PDbfepfO6utkFDbdUl
jsFs44uaEnipBOYJeSRS4Fx4sZLBf8jeuRpc8CppeQgnCVnEU/CgRcHZedZCJ1omn67wORxzWvjP
CsVRax5anzgnBope5r+/VCL95+qiB87chz5SsMwTkqGyYr2bNC/t+mU0Ub64lW0AZ+qQc3NE/idh
72UU6rS/vtJfw6o4Vo9NPCNX0ou/gU6sNZVtnkh50N27WzTBLyT9QrJF2Lu1CbrqXQj9yXk/+g4C
GFcfSayjCZGUMpFFAfqhr2hIEeDlewC3K4lUak51jzbZpf91CSZW49+SS9Ojro3ima5kZ9ejuNTN
lf24nHcyfwpE8y3xMeBl6L1s7ngGnLHP2dyjC4+0XB9A3RVDwLlQsq2Gz0S39L0yHDkHAQle2cZR
8bduSu/xkcR/65rtRsBhc/68lKlEYhgSH8mXdSfJIfXS/PU6RmnyNr/I2sYhFDBKF4ma0TzGmz8t
2fOcLfawRNdmuhKNy/1kZlee87pBgQB7FOAuOSrnR6Nn71WTUzMaTUNg+U+rulYOyKOdaY18gryU
q6os6xCDtoj79XE+BnnL3l/EssLdgs3BWzrd3LSAWapzt0k55nJynAYnUaCgtSzKo98ZVz6wDPak
doXF/KskSfjzazqn81b3HepQqnNWmyoTb9daCi57maIpspjQFhbaSViyp0vlxbo3wDdhphDJ35PI
KFO7eJYkGdFW+/f/hTJ91+FGwxhHRhbgcvTht6brQNMUcbfrK0k5Yr/j4UAXTcFY6g4asTi26w8/
MKS7pC4IWKRekmTUgterJhP2UjfV/bre5SbEvPpqtXx8UYlF8P8w2/7YXK3f3ZQKL5AHfW093Qtc
QJnGJVJrAFCUjCFYpAgr4TXVnKp1wcFUeY3TsM7p9QxL7XG9mG5pPLPJW72Yriq7a2tdLZI34lwj
1cF0KAcudmNPjW4xC9o8Mu3REv6VPN8ne5h3vKLl22zy0MPABHE3VT/IYHN4laCcbZOLDGhJKi+e
pOyt9GudzEo0cTGqsQkGHSRPMJRtuxLtCNegYe5jeC7rky57Q/QW90i3CLrKndkTNYz+nJypXEct
TZbOYTgt6BOUeouG8vai3R3okkD/vcxM4l1IE2HBvYoz32y15+9NqT55Dqa1ffiJMaNkgNBQPJF9
IM1EPnlqksFRZG312+F1BxvnQ8e6Hhx8rAOBoTxzvsk2Pv685ZVDFCQl7UZRFz7l0hASiihIZXdU
t1+4zpoBfcc6e8ATgwegQxzjTZ0fWZrc4qMumziNbGkcrH9zQKU570TsRcGSM78dY+9DTf4uTnUw
XW/+byYj9j2sD9uRw8v6bHwcHCmD8v3fjgxYCc9IEMD3x6unAHJphuj96X12q5aSN4bX5QiWhpqs
rmM0yD9b0i0m2zkxkEVfGqBOug4PJSCAC9QOLw2Eic7gWESrgmAiYOnp1psNthSZ882qCjhO2BqN
ZYXy+kcw4+hVGS5NkyH7Dk2X6E3Wb+DfeozQUbvND5bPF7xhA7RiSBuqAcg/b4uV33LNf8oCtXQR
CkT6Q1mza1Qsegy1PIpEcowZIDLvATSc/sSbgPQWujrupesiGpgZHGiv6Ge7MVs9hMj3Uyf95OsI
njktdTIuPuNBUhHj6HWXsXQQJifT9nl5CtPlm5YTeJ6vw+RhxpLbmKRmjheizwk0R87JLMXWNIXS
eekO+Nk9f2KUGHBlm0fmj5CcjK8PyuqWfA56ZUpQcj9f0cize1+uvVRdShG9ai4abDEdPfnq8pkz
rx9VQ00qVh28xEU6Yq2jo5FQw/JyF0zZ1ZIhVFaoLagETvyypQua1z5gohNbbEWgVltrMjZKX1Zf
GyB71czSskQL2QOuK61RfInm2jgBHzEGpYMt9wj7297jq9j4VERJJk3kGKSI00924iZs9s1Foiss
/mmkKLK41XnGN2vq1Z/FCwLUPm4r3Z89OX/OuKn6ROGsa18GS1MDqjC8bq4diAaC0aOtyMd41T/F
HfeEqptO9g72Uc1RNlpwV8tCdVJ/uRaKrHpga0/75KUMy2DuluvMXBFLGTnMH7EL7pVIi8eFzy+n
KaYawaJfL+NN7JoPt1oYcpzwLt1AdB68lg1kJn5V9sJXIkE2kJSwGwqSyLXnBYR/orAPt17wzjpm
ZzNK7AeLmY8U6jbkXD+z2ULKOAqdIBGwgsVFF8LWuaZM8nX3R2Mh7/dqDmzvgp/nboTAH3FwYmO8
KiYMC/WBcd5GaT6FIErD9EoBWc9yGmerQYdh/ZKT0eZ3UG6BmOma9BF5pcjTRClZLV11Rdk5I8U5
fWlB1IhWT45eLnXy/wNXJCLscJCT5TQhTvEVslF3DQo7aWR5aZo6MPeke+hDPrg40aHmpT1eLhAu
FEQ6u+wkboA11pZ3PgNmvuHiK8rjvsuVQPodf8v6FU5MhgMB3VBLPB73XKpwmnQP4vvlMompfvAo
SnOTeZjzp9QvxNOYEaFNOHy9d3552MGBz/WE9GDDDFM67CioO71fhtQw2xPBs7TB+t708alN1fzP
ja25BjGGlhg6S0LcUz/+uiwvcX5j6FAgjOVqWy6ncLwE2EO+QRdU8wvyz+fxKFvP+lw8eivF678+
xgp4o+noVttk6mq/kbOHZb+JGRYa8mY6IfoGeNLm2jNU790aC90yUACHQqUmrYMTs051qHbj3UUL
uWrkQ8AjLroGRwGv1rSV76IrpWKW6ukMf/QbeZ7F0qLOUmucGjDhsqkSm0W0IXmkn0rabjHZ8Cwm
N2LOLYa7FlKODh1ImUM5L2qsVXGY/H0pLYGGRIe5AHwb9yMTYP0dmttUy1K7ftc2Z5ZWxL6V9H72
98ybeXeIzJ9KAc0fTMtHjiOE761UPMOCRJxdsT9mAsx2f7UhAYEyoY+N7kMeqWbdBqZqYQtvg3rW
sinzIB3kC2ssnip72nb02OgT0ORVAhR9/xk7RKel+XHdl1vSmnSnlMd1EN8Xq15msQFushgLOYg4
9jgz2R6x151hJ8ZxdexunNwZoRtdXVuV37dR9oiV03uWGwEGrovFU2OWiUSzSeVXWpJQvDHkFEQ1
VkX9UEjwz9f79U4b2ziDDJI6oVOhROj//6WG0361IfdWXWYo6yr1HPt3GBXkalA+ykNU5oNxVkXU
Vjc3uD8dXnJ40286CKDNo2oO5iXE/jq7ib7CLGzK2LGJlAJNecnYSwD/mc3Dit+11Gsjaw9nZz4N
lumyP6IDRXYd3v7+MW+DIzPMpEdw9IsFXBPZv6/qchUcANgFYo8tlRqBWkdQ/jaViOVgH2h4GIls
lc2pOcENwZk/DKoT6POKEM7rE4P2lHAsQA1OovzaXWhBsKYYo354OhsAgdjsgvpfMuTWf1n5nuhx
+7Xxp27XF6v5OvnE7tLyhE/y0OvChaU4usQEQZAWxCFctMuONuDu9Nd9fJXh1NuMCfkg0raVVPwF
0rM1ZxvlSJw3AVH2b08bbIzDx4EFspiF7hW50bMbeB/b+qMl9GNQF6eazvaP7ERGUQk4uy0moOiK
+3KtlshLUB/Pvl6HV8dkHP61zvzeA2glfxZHwnTeFLTr99sN3U7CXydhhvdQqu7YqubSlYKIYpBC
q8788gETjdiatsoaPkjaPdHqAAFbbJG34ClON8bN/ASF31WDv5YI9Pafwf0iRWOKujpkHTiJZiEH
e4jDV8uRZSDUrUARC7WSWGh6TN5YTT3zElrRitOMIjpG/GscsrprnakMDOykn7uCxKHAtnLrpX9j
6tzR/FRAlXpPAac2ZSe+17oCVTgtyUVTk1ANdD/a6Mylv9yqgNmYYq5hZhL4SBc4DGplXKuN8O3X
PzNUHxJmoJj9bnTQj5MX31qhKp11oSIoU9f5J7miROfb+5upAtSl0W6JuEdkPiSKx4IPidUxTteB
y1c9roeuOK+6SlWSbviHmX80HCjEnzWr/0Ex/BCl2ocEuFt6MaVNKfRBZWCXLna2iUqgRi9XzcoO
NUXVvwsOSBF/FZEMtfNCe36O3OUHpWjEs4pIMtdekNS4skE4ASMU6EioKo3hPh83r98duEh0J0KH
SQn1HnPUFHMoXshb554a8Yuayh9VBwetxmp7GRQfnZXdBHmqUH0Yi1xixqS0Bub27WBGYCb2yfkA
U+1H5U6E7j/QWsXxuNtRwJI6CpYPWlkmFOkaF5w9aXjENZ9KRsoXd3VXRhzhP1p9PfI4qIyYW7oe
0aDH6WTrcGHvE5PEEl+jjqjO+DnYH8EtriL7evo73hRa/ecDFdNrUmoXYJJUxhVK9H6U4KMAB3UW
wOTTYdkyzHYVfelHFWRo2trKnyekSS2J2yWGqZUrhtTi4sKlT5fxmwNapJ3jFUL5bSeyqrHrvltU
CmMDgK/iZLSXT6N5q/OjdQnyIX+IeGEx+732b0whieft+ZQKizh+4EZGbBg/PCbk6Gyx5n7pht8A
OU7tlfmeoInD/LWx3araW8Xw+pH9+6lJd7wPJHcnSNi/SN+VvTnR1LgxMrYA2ayCAZXAmaOE+4uk
WW4ckhtnM1HEV9EJo+2KNQsQX3p6GIijZYc83syDgAiH8aPWKhD0wLwKc+lTtrEPKFryRrfWamT7
rbkK1LNNCxv9Ec5J7hxnwWO2loh3ERLUXctST32cLrQWngPIm6cC/khmzEEx17F/etzCLrRa+8nU
ke60tpt82t6BRI3V8Kv8ETN6ZKSbR3gvUZenMtrXZtrBweomtdICjrvdLeoJFtfJJzFy83ZAnOWb
09UG671kQDwaKuPf53jt6vZpijOp4MJ18NV7cp9/AcqZTwbH8rfM2FktacRdCg/O1iQPoMzIPpLK
N0Rw5lkxasHwlgJlLipccO/k4C0FhZI686LJ0LP2RJYzHtEQ7PBcky4jnb5s7w5RGPp5K2HGyYoq
IAZpyfdlmUbV3A3Hi+NuiyKUiH30Q8WdhmFFCbInidRv0B0IeeTEHSNWiYENNKW9raY34FppZcYB
uLaCyp0Z4cz6e1H7S4ATJg+HkjJndKJI5kq4L1JZKc/0+EsgDaefwX2YPrzmmGk1E1rNwL3JNOXm
4Tr0mlC7k8OltvDoGa3gGf4qlSUAF3a7Rvozc96rvljC61iZgTt96fnDMWZvL2wxLnkbpEtXLIS9
i/SSnwIr4Tw4bfWAADMqG76LeIEhqf/GXSVJKsNVToO/RKS/ZwoFHu8GYz8vOwMl/Qrq3XV3asq5
3NmL1kiIJcOugD8KtxfcYLBRewoAweF6VNN4jVgsqg2AHKezyS1FT3SFTkSOfoFTv/8C7zw9ymDR
6k7rfFm+KpP4FaY9RLQHvOMcwm4BB2xDhKUoM2QUkM10zDl09q6MtXiSBK3IcXY547P8Ejv4kujX
LLr2KFPuVieINBTvWSpuJfhf+dXwz2rOuGblfPB2HWYi+Vq7d7vGs44QVDyeMOQ211rxz99IQqA9
mWY0Bdi5wrXnPqr1SedJeE/srfZdIlAbaG6k9WmQWoZsl2WW2qRDEsqHTACrQPSTi4bVevQ0YFf+
y1+8lgEhEBvPUtBuaGrPNpLrcwVkU54SxuoSf5c/kcF9GlaJ/WTw3SwUSOpnE2y6yro5RLm2klFp
/0Y++y7Dup3dDxEwF8x0JvUYLASoqqykpOaZPweISrL+t397DmxYVXj4vizkqph9p1TjmBWvC1Pv
ePART9JpaXJtGSDZSQZsp5xuZdhzWNeFVXWhcCCI436bkPwojdKzuSdPZy1+fxFiSEQNMYaSy5t5
ouzm91ZI72RohD0pCWvTbriEor0u69jVEiiTyBOLXCFGXi98oXH2uI+jcuFAeldd0RQSuiiKMab8
HKz3KjZ5YG5L5Df80w1Nc82hDk7Bn70fZwpq74n4VLYKQrHAQju0CejfFRaz3YD47geaEa2Zst8y
BqE0ah6hDpPA+j3Rena8rSwMGfGUOllRZx5B8G6dYWkycsGE4ZGE1duH8vTIvMU0hrCv0x9Hr49b
COPQmaOUjPM6tifevzuUkr3V+pfT9zK+z2KRT+3jwQuRPnqIZMQ2HnXdKMtw9WSOZbOsh5c3VhY0
ZJyi1KRPtTxoGgd/6RCjZRoDlA9hMGLfU8f0HWaZqiAB/02dy2kENcItOSCYKTG5pM3SikZSnn7x
ATkv8lr1PrEKmSQEsjvOceBE3MaI3OwJoADDXvnqpA4itxKIGXtENMQtU4LOSbD6/Kxj0KuGrwO6
aEXkk7jtOFEoOhFXbzbxnIBxU3rnF1Q1O/qN8PKLqOT61WijpFqeo+f/Bnfe7o54p4Rd1nC/Rjyt
o2C+gMgDZ761UqtsbZKNFGdWQlqBSeiQYyEXie8y40Ex0AjQHmjgGGdKo5hu21nZ5/+e/Zi26sjE
kqIxcQ0IOHN1cgJOnDBxp76niol1ee1NQ58oYZ8i7FJG8aUNXu7IBumXtaXUlYrkI2foPAADUl7z
XR2gxNZnP6q9ravTvb+AB6vvVCJDu1MPvfiHDGImC5TlMNIkxwtZFaTfFYJBQAqWL4L1OhyPQn2D
Rf2lVMyQSw+TjmkBbTp3Wh8+KAhQ/ttZozB/NbqfDvep/QpU9HVcXqOxUl15WTvSQA9wh7BKYlu/
l8wwowrNUEIORfHSfC0o43nWKludEJ0qTqciQn78awk5XONRrhvrCpucL8wB1uD2816JYQ/2vX2a
gQKje8WkUuIBwgYp66uziHmRyXq5cvPdofz1KZTx37attbPp7qaB/8tJiAiyQOH4qHm9w3d8kEHU
6ORuRJpCrgcbtXYfr+lJaTTTQtsmAoj+/GxJFnvzkQYx6o5q7mfBrThY18p+qhmQzq4VWlSzZH87
y2kJcqsuJLkIMaGa9XoXrl8jrgwZGQ/ZwkgJDP9f7+pcs3cc7hx9hOk5UvpV+Go1w2c4deOStKPF
VReXxfVELeUbguSrfxBUVf3z6P8tb9KUfE5w84vRJopQBEigfIc85MAK/Y/+9US85bxJ6KcnVOMQ
N7MVFue7WsT6Y06PBSCZMF65ZaK2vqHnvUM59te5YOnzd+09vIWuTK36PkoLq/5PBZwL1GzHqlfx
e7UEsHu65ySNNu9SWZSKaZVkLBFsSN5nYX72XYKDfN+zbRi7E7YTCVN5vzkWhr2U/NqFyhYFRRf0
tTTJXYdfoxfbgnVNUlmFvFvUfsn2eQX4TngcmXtA8KzfQyX6qEGgI4dTNahba8vLouSuT16CA6sZ
2pv0OOBwXzbys9e6VmMS2nQm5El43BXJpLYaqI2R54OI+yP8Y565fzoxZsQJj2ZlJvnaZmhzN8mB
a3CK2bOh0UU7vZzbBWbs5bg4gvpqwjGMLfdK4j8MTConqrFEQ3s08YtEHvXB5J0XZYNVSEycUKlf
k/9r7dJTCU4V03Nmdy8YxJ2On0JpAWnUdUXn2JkJ+lzi+c1ywjC0lf62dRuTt3yENnwNEZ4OKdIm
Bzij/AXbs5GymDNwW661RNClY1CbNCFN/b4xLtVedpsx/YOPtPBsUyRyS6UDkGPL6Jpq2o2Ech8x
ehef8dhXsqtFbzbAtrIygP6KdznNqOLtDlNLlIdkb+gR/qOcAXbgTWCaZAKbYLu6YwU/WSpXvIBP
KapquQvEjzBmcPdDqpJc5r/PZ07QXoWzPpt76Qs6nzpmy6JbWv/UMTMCEfI//Fh/6iXTHtTfI0aJ
t/yR0qP+3Sk5DXlPDjvDG64NRjo0wQeG8JztJ3E1vQ2hbj9wY87xfgNKOq0sWSOsjCn7evM0+yOy
uvos6OZuY9fT9Rbh8boi0SzIxC0JiLRqv1CUQ7TyNC/k3VO3oj9RgXtRgpJnXoNCal/NZ7odttl4
BXbODtTstAOKdtji8D3s93OSvJbyaNAG5E4HnqCEMDlpv3H7YLAzUxB2WxdgnNjcfESj3tTVsRrf
ITDL7g9a86/0yPCYhu2Kn4y3csRDJ9fQwo21WSVw5xOs8KL/aS9kqGAeRmwCLMgz09ULeBGLvsA9
O2Z8vmWSPlB/wG3it7PU35oE04mA+j3arAzX2AN7D40FJd7uTf0hztaorWWGE+ZjWskBLt++sb3D
zytYsT0Dryvd5rl7FJsethTp0Jw+YvHFupFLJ6iek0fuRnH8iOyCx/5kCkwHABmivHQ3BrCuxEdl
wEqyL5+XYZge1QfgC8ZAKm5cPcZm9qlpImoHubb+m8HwWdSayGQJ9R9qO4u5xMShxFhqv5NdGIwZ
A6lWILq/QOSnYVH1agYjfS/YWx99hOvrch7lJ9mPanMq8JCMWrt5anJWq/gs94XMY/1cbqlc52i3
AIQyMarai//C1gP/Ktxtmml7DGqqkFsgNcn2/X5mdnb5ai+mnfDOILNySnSLD0I/qfF4RwmbgRKc
RUzZT3TO46oVF7hgkLUyYLwZlA7S9zt6vgf7znqxxAi1ILvn+BSBKi+moeWIjFIL4oUevXNFxEFn
hHdapbmVQ5xQBuGGZ/7bbaML/J8t5GvZJUGW+sn1UXRZm1x8+6lwiqIoTIVUsoVGHs84c0AfG8L8
N4aex2TZVVpHy6JHP5oQ3u+9z8Q7dTrkihO4G+dsm4KRBuVQjmYliTWzdN+uMC9HiBHGn46kmA+K
o7xA6uXO7ql+vDyTdTskVoxt+SZXX0YLyV5n7cgW7qco12lYzHvX8XQDMvaX3OCGaSkNXDL33IcS
U8CWYiZaz4/pzAPCi/aJbfDlWukVqiVWlGloT64iMQYDkODVP1Y8/mKspDHd44U2ZtdirT3yid3A
O4YC6I5nd7yeejd8nVQKo6pnu8BrHG4cIcB33r6NAsSNb6Zat4gnFInTrtrBLwfKiAK0B0Qk7DOO
LZA0GFVFE5AErFnH+papFb8bKvpLwgrx887qefrwIUVrq+k7i/GwkR/HFXWMoex6JqObp5juvEU2
+ZlzoyZdGPb494Fz16kWDESNhFGWf20Ro62qZ8kzuGphUTXEX3pPQDriEOQ1xq9HuzPwc/5qTiwl
Bj/OFNp8h/GvGZDDtSQ3mnstM/1U7Mcsiz9z0aWSCCmcJzjYe+f3vq2RzXA7zK33TL5lXNh+4MOE
uudw1NSddWllHdG8OHAnwMEmJLtAeYYO2aAazcnMGnkw5YkCVTaikMn8L9k5qDbkHw9H8f3rWFxO
5pEmeF1OOdpdedrRl5bfcjIVP/iE6RHbJ4gVPdXX1vuIAWAd24K+GD5E7Jopgl6/1ZYwZQfIr4rb
d7cAKfZdcZ3S7f1DQujiUUftr5iqvFElp64+PkkDgYglMijRNt2+2JebDjcSDQ7TXu+AAKBwVgd1
BW4Osjd15KH85XTnGkafql2o/YLZwHJcE8Nzgkp9bqNSV4BGdmtu/WtCIGTLEHwembMbDHbNnwpq
69/7FSSMODsioOuMX6vliqKkcFBS9qIECNiBAbwcsZYRsnskmUGZt1lPRxDZH0D1koChlKF+TN6X
1s5p+i44UjyfHlqAlhsjDfC8EkL/kxGe7ZNmQjgzShvMih25VVbsonXUVXpTgmKmS16HopUcmaMD
7Papa3VbMMi2t/2ftvLUxkLYEAERAF8abWvQe0/H3eUHSroIkDfLYCkDNndNOkGuSwAomOJjiOWB
jTL1c0R0Vp27UjP54trzZg1SrGFuI/rEWur+fQSoXd8f83cDhbSBpqd0DqZt8UYDBXv8FlsiruH5
CFva386DzazDHSAENEDS4uLoGfdH2VMkN4/R1SerjhcQ3ut4N/GmybUba8kJqaYMsEQY7wSNcBgw
xw687nEecKv6Cx7JXDhFAACUHUePQHcUaS+whyrL3T4zgTQccXT/xjveoZocTttDZ8uWoe3A0NZe
sA7r8jF/unl5D/tSOg+L9iAfWvz9s+4U7m+ogD5/7aoC7rwebsCoezqgd9FrdRUExlzNozuwE8yi
ExDkBTtsg8w9MSwL6jo6xkegaFjTwHQocfbE8OUulQREEjSu9xLLLBqV8XwdSP6opicGhnQyr5eR
uoxsoltZVptEVji1i37uFVTtZBPBY3j0TSel2EclsfCql/nV0kUlIfipE1oVdFjkfFS35rK5MnlB
kn/CKaOw1ICmu0sxiX/8yzrd5gn+4p+Ij3BF13XVRVVzkaYatTfZYpkJc2EapefEL+pKbklobmte
Aq6k5a+5xY+303KJyNc0++WOcPRJzYHhThvpLkexUlJh0wCjbD+vCjXyzXthtwZwj4Dne23W8H1B
SRrS+SJJ2icDkEHVuC3hohX5rbtNlKc2IBZ5gzpx3OdBg5EzaBI48YglKsB2m+JPsE3ZqDpZ5tNL
e0n6dO4yGv+Va0q0P6BeGroqVEMK142w1U/6vCbmYpfxWW4YsC9phsMkwGcS8BJ7QOyFt4mV4guu
LBTzG9gUtiQHowNj/2Fdoen+MZHr6ysQM7dVHVt8gOUpvFuKJa+EJ5lzKxQofWXwi3fklQRqwIfS
QZNQQguYFCc8h6KUGMNW9l3erJzguZIiN8cwGSKB9frpav7bQ0Ksuewqv0K7FP35fOwsq4rwLX7r
++8mCkO2udDW+JbBUqE3AO9MbJPam+DH3IdeW/hQBgxqwg/zW4whEQIXk1jT3aDXFD9taimtbDcG
MoMV9CA7b6tMgLbh742c6+9+xtHb4Cg5VlxxeEQszvbscyt+fa60IN444cYNXcoAQ+z5lUmjqflw
L7Iqw2EczF+QP07ytIvMW9yUdBlZS88Q5ZO2bxrVi7U34VyboktkJAjDeRsyCfyLTF8Wpc3rYtLj
oIpB8kPiC5fzw2IsbcsvpXKSFobfCqbu6dGxQkVt3xkIlfH9cbAw05qFc7BHW5VY0y1FWMrDSDPc
NsmvMmvwrf7nrCd1wVK2BwQckxshUrTEebXXw3zxJJyfKwdj1iL7RM//AVhE5mpr75FEuOeFHyhl
pfnoxI0Ta29Wu9CA/JkjZXyabOYGxnZeQXPhGOyDEi326amJlPvBaEmhEimegNz7QKpPEws33kPK
NcE7RJzD7+8bVdOQb+H4J6AFx16GhV+ZjXzxGPJEktmbD5m5vBgekac6B/GKF2ZXXXFptI1Z8S+a
g0vSCUySeLoKDpOL4hhLLctOh4mF4Ng4wVxK23jNAH1uHEIy7sD81NTa/vL3V8pM0WUQjpBE5agt
ZTK2VRqSP07HVLeF5o0DLQ/L1ovX1qRyr8aG+FYBX2W/nx5wdDemKV7Cd5nY7Y9Zhv0KA6BHMp8b
sjjQBYG9eXnjFohYik1CBq1Sb305yDECf/dGcyKS+0W6p0vkwo4VD0Ivkm5CZx72TpGDh6opTuCk
lEV63e8WhUowUEOsIN4FkxKCw1B5QKlDgDGQXj7oho5knjdCrr0QfmVoJmitSXC8T0J20dR6+uaf
PODVg/cfNgsFimHvOFwf7GcLHxBAOxR69ZrWRPc9Jxyfn6CXeeErsx2gc6lCLZFgLPD6DEyA5E6n
WQVV4PJ3bBuk/XgtgPhxEEa7mZxs0Ba5vfckA/SP6fsecP4KB1nllwUn1VXlxn61Dx38/7F8bGEj
5AfX8FCwCDCuGV1WRJRvLM3nlOUgts/nsml0l4E9dEMJ5wG/qxgTNbXtBv+85OcwRBLuijTrfuRn
N5t5mnFwxu4us3qe2v4z4Omy0TSbfijILLCkQfKdjnhr6mOthSmR8zNmyhBXCC5ssT3lrR5pq9OI
XVqWaxAk4vNLi4A8giVjMfVPmwNjlwdq7K3peeR0sHQY6lUlUloPlquUQ16Nnzm/EvN3FcV5/MQT
/KKXv6qeXkk2vq9WEyoHO1rZHnXtKNkUSvheH0t7iWYwJCx9llQBCVLO/l7rTTs8fe5meqDUnwgc
kASHSqhUXW2KewZR6PwSiLRO5P/2zDOVXsneCrF4dKe3afI13d51B+4HMmEUotVT8PnGUQ4EKGxr
BvOYP0QrVfFGyPEZigiCvyMTyhjli8Tbp/Uo4tQmCBpUDJW9a1FhhjJmTM1EXjMDh4tK1MoGOLU0
gW4+K4mPhnx0ohVcsVpatN9Wet4gQ89agWWru6qQ2LKK9TcXrPAXKX2whEq7q10nMc1WhIGKweaH
T2pnfq+Jc3wFIYFu9vlWIVil0+VnuGtLvwjYZYFIDN/gLpxgSJbyH5MzRabOVg7oSPaiZXzF0xEf
6FnTNaOfLfYFiwJqReSlYWbGJlEzlYZPwAYIZTd2jvQm+KQkwE83NXdOP/C6JPNYZ92l+Qlsq84/
klyZY8Lz4mdaRtUnqtQ1UlvSkXda1OoFgUAXs2EOtuwy1l4A/KaNvfd4VXpKaj/Vne2nN1w+QONF
toVm/xQUHgf/rxFxin8sYbejUycyBAT7JqTK1D9uEHITQ2QakJDAC28CjiamfsB5JqdDt9v4vwHM
VNyWK4hkNhqBwkGEm9EBG95ds2qbho5BkEuLe5PhTIR4rtcMLRX+msTig+4T2nXFkJLWYoQnOexf
2sdHPKiQ6VLjJns+yMj/c93SBtSiCyKhCSDxTqKic4PZEGFbbm6Ptb+B/2Ez07SpUl9ibMTleR4c
2wWRBtJxbF9hoBtKcxkjK8b9B6TRRvPn9ZgudxzuX4O/UtM+SNCjhza822ODIIjkyS/6hdYg0qVC
wFm0nAR/liHNXDU0H0ZGuPMghvaMjvtLxtDr73aHYBonJ2v3fvJubYbWKITHjk+AoY6kaIrGWgcr
x6DGc0moUzuRItt7Wtwv7Xf1NNpNYuMggoQG6nuwzCyBKx71IW0ofKGr5jIWJFfw5efvWDDXrHxD
7nODDdW/NFHTQPwkoExj5rQEEgs1nQhCcOenjR3fsV8Mhy1z/fAHqJm4m5OznCUql5DjVq/Dqy/T
EHTj4rU8DZ2oJ5IFjr87bUYUWjTp3dfj8Z2gIXXNs1KG9TekIR2/Dvc/zhK2ANpjgIn2f9pvxLsy
Kd7pRzqEHw2xlsx0RJsHgV230dd1EbczyN3mdGWFk0HqAgzDDHlXIrWF2Kf4wGvYMEIj5u4Ej8Pd
Bms/6IKBTEbuLo57pXZnrgMKv0383vT/0KP6Ugi+fmRmQO8Mij2WnfIT33TRcevf7q8ybQ0xCdm5
FPptC3YphPtFo6c7uvLbJCiBqzhWpmixRcHZVN76nkQQRY1OS2BWGDxBgAEMe7nWxOvgaw88o9EI
AUhMWPRNORHIRqQ5747yZU0Tc5cP7rG0pKDhVZ4STqTqRIFaNuXOJ38qH2ICgwhoqPtHtsAGvPLQ
EiCM2RdSxA9DNmG1I8lqP3TGR7yaaOA423Sk3oqFFf3PBcZl/nTdOqIegFZ+sEYjlYmXLmBxMeie
+pFYg4CCuINAHL6R4aLVj2ksbra5xliDvACZtBe1l7aCWpz5MkIdfoMGn9KqQpvhaAhl46tqArGJ
Kf1iwTnOACvK7rqFw5desqgF8niCf2XaiJao0lYqf7DaxYoxQS+/Va6o3dvBvX36xy0iqCeSE5gj
VpojmpU3t1Wu/TArTjrhRd6/zEPOkhFfe+FI52WUMR+RQhE2/NCcmpOa6KctZkyye6iDp0diD6pI
fG6Jyc/Eg/45hLAvsLtglNgEzGaUnS4kkSQ7+ICdC54nKaUo1KCCLLhAkWZlR5eHkGXSmxPZd9/8
BdhfL1fsmtzZ86jl2hQBlGbaWrOj6OHz2H0LaDNeSBFcBc2lf/PTwVDbMWiopIPbiBxlYz1jlmC7
vH72OeDmvBQpX7H8l2bTHlOW+Pv+k+W6k/W2K3BwoGHNTg2P+IvBmKMLGDZTbKkiTnj4gMDa3xiw
OuGLf1tzz1iyZo7DAPWVPgBDlk6W8eQJwzyMFzBqWS4ku/E1GHJh9qa3+2hY4HrdvV8f3h/jvSiI
a2FKLPRl29LSMKGRImEmDruNZH3wgwtnOGVM9SnBg735qB2zd2xVpYnMUmNSL5vjWnk2F4lXQBhB
gpHoukyHy98q1S/KCQgNaH6UYxSNqjvu88JstHNJ0c6aT5JSjEJPo3dkRr0fYdMuXC/X6131OGQz
n0/+sWWyn0TCU4WiZ7MTEE/S/k6yg/+IPjv5MaJKC+mBwBZUtZBPa4QrQs/S60J8ETq1hMDqc7s9
Z8xxLCPTJwB29Nb95tPh8/tfpO+/giJjUKV+VL2GjcNHYoNUgeeDrvzka6bzceIihhDqNsA+i1ot
oOEEtKn7T3sOjMB40xYUT0jYORRjCngE5+c9yTOgxEg2+tJ8mh+CvHBEvH3AAvImUEv0VYV7YWuj
fyA2w8K+xGyuvzsOugy4wp+rkt8yIfYuOuzjOnP20zZkyFZSqlhaxaTVxVlFBHEy1Zn05Kfahwsj
gqspBPYcR87JSpB/nZq8M5FYA4qbnpZfzOkEUpSMo1nLVY7hjD2+dVPZcdrxbfVcrFNfOGosNMXR
csop0A0OgGKfE0jw4Nh2Iboy0Q2oXTA+v3H/hhQyfZyKeygpMTo0KKEo6bMr+3rvy9QaJkVi6Iii
uI7nl0plOi55MnLVQQyImOWBgizMOpmlIZhQVJTUUBV/d3KQQCQZ8u5aIYgRPh1cu7GQeooSGzqT
WUSIsUNx0sZk7nJaaCyFNV7rvTfPmCAsoXi7/oAGvSE5+DwM3V1VZadJhFg6nBOgaPHdR+XGmEuH
6eIom3xM/XugH5eLwfNSz93op9rOxam3CeaQF9Y4usdQa8qYC3byUaI9Lr1bJPOaBI4p7i2db+gq
kxUMrsOrtx8HmN6fBqxVpsDwFgU79ASohRYrOc6Qkm/JKtdLo2y0SX8cZJXZCvRKspwkAkZH0NJQ
bIsB+qa3I1cUWGowjmkjY/LbPEiznKFztVXUsJet+03WeCcP4OH7VozURObmwR9fWiZ/57290Em2
U5l2Swx9haMF0SKKK1cH8VXZX2HWAUkHLWoVND0hxtd7Bu/K32PXh2AeLwm1vES03Y3rKgScRiT4
2zs1A2jQcWpOfP86KPbu6baDGPvpPdlsenA77y1Zy+4ZoW1/TdXSQlx/mTa6ZrhVKjWmmr0dgNTO
0d46XoyrzWe0t6x25gCMvG/kPLTxOvhwCJZqThBW02bXER1N9JqS0Ad9ALvLjO6fQNCECavpRnAS
56uyo1oVP2dqW0tubTO8GBqEIhTzkwBIcm6Ayi6dcFIz7WZnVmy3k6/ACLmrDL8zD8qZiAYPbUP1
4eWRDRKhG5VJYaXKe4RIEkgOIhnez4hHSeOu/BEy4dQVvFMUkG5yilAhlYaVC5zBNZFdn+suq8u0
88MSJWczNrc2sJb47XGw7FyOdVnBrKAVinyb8gyVp3KeoJv4DznEKCYGVqYsmQbUZ0DR+5tt53fw
2O4jOZOjJ3FWoMZgKDAE0yECfZ7ldwKmnGWVCJ14xYe47uu4NMPcqHC4+fltY4N0Q7Tinc17lSGk
6t4CmQZgVt/GOHxr0hGy00ad4TIp//YExzkeuFFBa5nondPC8M4K12yxA6xFXw5MPILql/NtL+3z
FIqeHuzYAOvniCd59jZbFsrrOdM637AoP9FTKE/ABUfgzfTebxDYl9VXBb6C567thfJLK1VJzybz
ddwaO5Lb/Lr+QktlXJHvKEv8MXoiTLPONM9BwTBpNNC0MxfHNDT1D/7WCvU7PKX4DiFM9npvBeiK
pe4f8viMpIRNRIgwXMB7g6+e0NXkTr1tkAiUhgPkK+0b1VEn7hIOm45KNCR2RlRrpQcCoFik16eD
O9jECurJt3t4sQaJXCeVxA9ItqPrJyu6tibOZaqqUJEs/NCGhRBivsRrrZZlYaWON56wfmIJ7Dr8
eFN8HKZY0GiW3OB5KL/qK7iyqZhGTlQOK63LYV7e+FZvLbaR/K+PssYBp56q1go9Si2ZBrgXjzeI
BioQGlTJY2rl4XXefJQZwECptLdX4RXBLykzeB3qxG/48+JbQ59lYfRoL1vuO7Jz9uVV1tZGsZml
BOZ7Pea5sGjieHvA0FaHMcbAOD0t/ivfu4w/8maljASYcJiCdgQHLvq4QbE7QKfvn4wqP6Q6cvL7
9kqdFvFp25RG8l6KGXcHvOJhic0rBDJ1f0QdbFL1IEcEgD08mHc+xw529VHy2Ago3DvmqvmMLAir
6sdrOqyPxF7xmacH8WOdkXoeNs822+uia/nLMGge6wgYdnx5VDdjc2qG7kwjqcX/qccCssG3+rnb
cpr67PVo/KU0qW4BF3lSeyWbLaBDti4tFF3PDKRuc8OfSgznEEEWMb8CeVIEwvdu6VhCq/us3BB/
Y/++0RLbI8ej2wwuJwrI2Jf3qj/3fviZHCtioDesEFxqeVBsX24gb4EIrVqHyJ5tUaQ8fBOLF7o0
F/fTb5AraCSDO+j/qUrTnbjHL1j2fCxwS602v51TPLUxs1qA+sdSqiJso1Qu6XDd1CljLJYHOZgs
Y45At5OIT9bPYJfNoutw3cVDjj+dNa0cwt2yOdMhyDqufRbQLYGahLgTe5EvwaqEFzEZP8KNdHOx
1+XB6r9fGMsOBPeg2k/9mgMAZ1jDiNYWlIe/al2im875I1EazSg1Eh2fbWCxMr5HtQ6Jtha5EhjU
ITXKXzfeTLHvui3+/OENrRSSfUPgNnO2a9otJZs4GzYktWsiahZBMSjKlhU3xOfL1HgMHo426K5W
i3iEZAMs2x+PC59EVvfND3Y+kjRjOTbIdOSupfPgzeGAQfLusmkaYCmVPPgncA59c5GGYOS9N5gH
qGK2KHhW53SJMlkFrQUtc30rTl5bSLnLQSn7Fs+p/TrgpYICLYg+PXrLXH6iwFuN5+DFqwHhRbTl
qcRj16NPiTOZg6zfC/zj8jUm/h4/t5n3DvNy9EwQrWfGbnTSQNMYgpznwhatnG0yyQrbqYnuH790
jhR6IG9H9z5dYBuUZTyyKWz/7QIveFtNgrlctuQEhB3wpFor38dhon2/7YRj1S9jJ6YXmLEVONnz
/lAQFkgU3luZqQuDkArzjxNqNaUKJDJhegJvm6H54psof/3YhbX5YXfg5dPjmYsssg6BKaTK/m2s
G8Pt8pogS2qUW7i2sFi8nqfti6BZJ2zJ+LwzbcFKflYzoSIxTCyhLYaOHbQjkBpXHTnolwGlb0yn
vqwww5m3uLYlwHTWp7GA6Rz3FGQ1PvhvlHMhiTwR3Kzf0+mqUwUWwv+fM8PHHxm3lr3KHyLcaB1N
4iR+Zrnypw6v+Yh1+BopE8g0djn5eKNKD7LaBovrJEopjfYSwSLiEPowumYhg8sgpcc3IgbVOVPm
etjaszuEKglq0YHXQw+myl/nfbY645we/SxYq1fyCEn+OKgYe0/sdRrJ8j5Twli9hupnwLROjqwJ
Q6mBBvcGnTf8EYtI6ANdSDb7ICeH6OEj5WVLSul7NTuh3c63LDPgeubXQ6u+ggPH+BzhZfx+JyQX
5Y3JquzT1h8OiceN5+UyRF8fhoMvQ6SBJj+P1CW+R3+h9P9rKR/GcVuSbZe6FeDqaNJEnu8CJsWT
6LibH4cOkk98g66UqG/8BaMWwB/SXvQm+66Rb1UhxU4d1V5YvVRBXlw2AsEIWJzjo9v9NfzN04em
02ZxAcDvqi/fOczjhVAdxWlfGR/Dm7eTbvim5FF8oxtCMWZt+Z+NQFC9PCI2+RXHLJ2KEoCyLZwe
sCVma6DadGxBCROL5DdYX4WqJvq/fHpRQBGW2h4EbHknw8L/XRLKnlnP01087QNjN0zHKtRNqG6g
qL0ynDtHm3w3hE6ITFXhuY+t7hPA4NOkMQl64K+z9MHzWDPv6dTZ7jHZUhdCVjO1JBTyo8x7qZPi
/57OnjvinSCrBuE9RcYfvr9n9YnL39Za/42dfZTBOjrMDTX13aVfcc4Bz6jnu3HyC3TTC6TPFbnX
TRd3+csWMxnRVH+2Cgleh5Q7SXvevSvxdEa50QKIhMHgRp+5d12SZDeGWikKYcu81BKK6w8f7oM2
eTuPBmiMxM0drJaeWQr0Xc+22CVP8l9OT3lCzNWnihmrWaT9Er9u/jEgS3A4zAFOZrDhJvKdwnch
da0mXubjfRkwGvcukDwQDZ3y9Aw+b5YUwswN2qb1DH6gbRXEl3Kg4sbJ8M2A/CwMuiTIZsT/TiY3
d80JdARZbupC9+1be6+ZO/k8sIjH7hNoXNDBabIqePLl/UFJKhjLBpY9IwFWAIaGJrA4MLByF6/Z
FqdqUxeZDJkh/OqYhpKNAbofgSPm021xewnDsd3nlvCtSt3+OsJ5J3TnpgXjU5n3Ipp6jOSrzJM7
URG07wNlS6DA1Nkzaindm980oX1i00MLJ4b1XlXHk7WL0U33RqS3HKSzAE45h90ddVPPx2NbiKXI
IIEmEGbMuyDlDkJkNoAX4Sez4yogWmoJScCbg+tLwn7LMPENcm2tCUErgmq/haD2mKDxCczjx4Xq
gUxgJ7Qn+ISc4+2kz/bIPdkkFPzPaGcYP9W8MITZUZt6DCCVXDDQ9Ea3hFvhAiKVCT+bEQhKRkiN
ovOdfoUGkpX2tdZlCunFvGMDs4AW3U4rPrDlDa6ZTZwspHE0VnVz6DqYzxEEqklfSIpYQyxb0ftP
cUrr8AJ9xCXzsAx6d4jvq5HUDcW+iciMtOcQw7U0q66aP6Z5VpPNGhLKOWziOpJnaThB9yP9rkEL
8G3AB9JSq0WAbxEVH6YMQW9DZvfbYZiMhh5P+BmjJgTAawA2G8qRnqvcNLiTnHNToyOjkb4MCQzC
dtXZepnnK2yn7jFJ9CnshiBoGRzlYwehj61JFeSrEftjG5CHi/KHMySGUTvHesIJDbOcQhLk5G5z
JyEVDvVDd6JYSkuJ7GDD+t/r8X10H5IONfkSWvseIfrfMSLYNATdHOV+3v16ojRwe90Ac2tqaZII
tq2Qqn8SMCfIMOE0n95E0NwefuNTXA6lx9ioLX2ZSJRad34Zca2M6fPYf9dd05IJrA+uOkaNpVno
AgQ0RV4z1T4aTLPJLtf9ZmfqkbhTmVNGcx37hk9f0DmQ1c0ntiZgnVCFV2OYdX/fe+2qsBYfzLkn
ipPqYMhOAeCEpMR8AL2fNXunBmymnyzBbEWTwqenrTCA94spJzkXnxYyaDNj4n1DzFKdLfDaqGcz
YV24ffasnV/wzDQj5NhrJO1/iVhQn3j/QU68lCxYtttEdYrAce58XseTYTpgCGfFOu6wztZx8wM/
ffDOA8r17f3o4wfFUqv9tk1LVSTV0BQoq3PFN/bs2xtJ4bIAHw/5B8FaPmyvpR0tbm5TukJsDdf0
HMqNbDhUYtt5bBnVTyYrg292qEQWJ2AQaliVBH+vrrFr9xw3sc8SQZymr9ukjKG7f8NAChuu+ya7
IWNLer0ZCGq3f4NwJQBBl+xn6ICuHtlEjEwVa71jkxTQ4J5q9JO9IhvdWX6wpssaDP04s97moG4G
iEl5zWdWJS1e5pc8qyH0P4rpcck02NZfvvQjnNh+v6dDHXBm3ML2R9/Go8x8A13tJPIA0PbYq9q2
SUs4BycaEFC+3695gS5CuT30wM5RWG+Mu8OiI1kZo6QvIprwACWiFpdpGK8u+MhsVENcCsfWGtCm
84IQxBIo/EK21QkBQkW49Xmyi5eQDbzK+kKbPQUBxsfn5pU8VdGM/ZVVWErDEeX4YzaUiCELHQds
UbVEp+RxSA04nEq9FjJkAsJVXLtvoBKeCCo+m80lxbCoSQUgxwYZJvQ72CnrEVHDA+cdnvqAxfUb
sfXLTRQGcwmJrOgOLOWf+GR5Nsno+c63CeVl9fBr2AAUJYoIAociTMVJkc0j/yxn7EODtKVN7UIs
3tFxaLc4PMZfGY4OtP49+15dXUVgyarVbiP5uS7b/EF8tqbr6UHc4IEVSDhgsApiBizL3Tzzhfnp
RRdwSwuw0fgOly6EtEpLmCi2uXt4T/r+O5zpu3tcy4wcPH1zLVFr8eyB9YcNdkub87cYJJC6NAAq
esoHBqvB6l5uvwi5+nhTmUHPOFcE22pPLuRx/JVUwVC4U/BffFoM0b/kGUINlDJRABNwkcVLR2ji
6hrHYEtzQZB4c4hFRiG6gs381Z3sZKXWgeBZ/2mBSVpgXXtbXN+aerxnqnevhLJR1Hj98qn8AEHU
6lRaXNCy/sUMXa58bJ372z4segzfzHLhmYduRG4F+x4BV6NCKYYKKBAz2UqvQAohR+ajrtYrLEnS
HU3sZgAJGcp1Czy/Rr6bY/BTmhafI2QxUhdxvd3F2Wo3XMoSHhO6jpeteQL3v6ObeQDFZFL7Ry/4
2oFeODQqNnQ1KlhTJegJC0jv7nYdyQAV89LWOSyiq4uMS0mXGZmDGxAGK+pve0ELH3oPvHWc25Ac
N0hXPr4IvkJSWb762m+unl3SQ6TfD0kMQcdQXempcgUxgJdsMY4qOehsjGX/D13kvL8s2zoeLdkp
2BE7/KGpiWig+vPCedvCWQbnC5/k2RH8Tj9yF9S2E6npa9vKjpz9eNgO0o605kCKkXdjlEhkWNIs
HxnDYgQFvppPHq6svaUPlRsX3Hh4NUH0QW3hirUccacDWFFnr1/LwySvVCqgDmNuHi5H6xZVvHIq
1+jG7jPdb8q2fhMNEAX5MgPxLswSXvc6BB2CP8wa3JWyZaqI4LbOjDkWUckyhpKDaiNj9246Vbr7
xEYLQImRuGfRefvzdrja7fA9231RPYD+TZfzE01UYRevoVxZYNT+xAhO9CZG3dcQOoB+jO7h/fJN
VsMT+PzchnWaB+2a1PAOp6BPvtt+NQnyNVfi7dqFWsas+7Vy2+UrEna8vmOEW1CjKDToKTDeV5jo
t6ajX2kr/9yDjMYpNP3ndAAUhH7nLOCUa7tfgETK1+epGQaOImH8reogBy5jHBKKmRO8cK7jB9mr
boP/alUh7xpkbsY6/9RErbQUIkZbv5uvFbO/Tg7CMm936UlQaZ/ptqROxNFZx6A+nkCsUkc6leNC
8Z3GCF22EGGsTLnwMf45OoTRopFjwz5IB1q+WA6ERlSmPm57GpZ2081ElqqpRBiTf0bGHuAc0prU
wqJpsUv3vousnamXyMZj2dEgLaxhDQHEmrNDf1+JOAVaH0VRj1oVXAamGC2eUVFQLJWN0D0R1Wwj
5SGMNS6QsIZl1/pg6t0NcJLWy8g8Ld9cLFnXDbmoNY+4XpPvyejUFsuVYPHu607QA8lxZdE4XRKW
aGfKetj6ibgkWKoN4kCrAmD8OIz/WaZJM6+k8BcTfJ/8OUIFLntRDxFhQL5F4nFLZ1mrcYBBAO1d
/RIAhLzgXYej57HtElg0AMK+lHkS/coMlm/jFsWJhdn7Ujlidf56THoxkWU5f/q+cBhjUO7nXhOd
ENSiXDUI1GW6iqoBTlEffaMfKch5k4fJPakc7kAoZzMNpr2enzcHsOSJQcD/ZsaOJcQCkRPu9n5Y
IGre7TVJR7KBSxADYebQX/WF4n9gjyVVjVW2SA+X9HYHTvRsuR6dyGvRXM/xnlp0bV76P9ZfJYg2
XTpyoz15phR6FdNp0N+8RXrjlUmc/f4j5IXpVgJ3MuQO4cuoMpT6QiuahgeFrh60cdo3NZdDyEvU
3Y8gdspvbCQNoeb7LjRQhmukwlW1vm6KJZz/RO5p3U4aRYgGytRUDe7QRz2Un06eErJSF0SbY19l
lW5zZVWvt3/0dTvSthxELD5wGkqAPxbLwy3DAPT5VdefKvYChOhmxpSNlxtfrXJ4s3Ui8EiLbVeN
iNZd3iK0aWfJHOGRId/s8KrY3KW3W/Wq7VUWnee0nReS7grNqPJIwzcsBI3PpvQ/Tzme+xkV+SKs
AoTAmBweWRQxbAJ6rfvKMNReP83zj2IYCSjkq6r2zntutWnwZW9Griwk9cRS2uwipuWyQ0Hz/9gW
KQY9NeI3k1oxit99gHdvVxv5zNiKbsZNREI20KF2jerRr2bTDfrCsTfB8Ubud4aAR/B2N1KleGpZ
wpzHsUV+XivgG2BPbvRPX+9/+l5GZIEtAHPP3BrDfg2IqS+VdffUEj/WtL4Ol3788pBak+4dsc8x
Lv0qD+dQ9TkU8c1Hnz9HecEvfme6VvNeXHQ2XvRg8E+D4dVbtol1euSnoOXwvAp2rh4l7qSR7bqg
LDYfFr/3x3eWQmYEnslkyoCnGe2Z/47vcLVYq8MtndXfyc+cXeFRwS44pg1/ZIKu/VajazY84s8e
KANlUjcQG85+TMisL2TJHphGNtK1zuVwtreBYpSRpzxCrveRknIKRpZRgAhKSl+24EPHWZEztBlS
GJjizKdWgggA0/WD8S/SX5t4urBh4J3w4cR1n3UcwAfv6ti/l8XCxB+M5mSr2+fsnojn0Pn7u2oD
d0BbUZRZPu7ROAqnSUC0+r05VKxz9TmWaADpUWI/Mn5UZfrqOtVDFmZaCjYhMosX8rUfM203JNEP
aAw1MOvHGLJzBwM9Yj0VAazDsxcEn/2eDVo7pzSmTW3nn2GQxcXWdwuJQ/wCrR+RwPIAnJzmsFC5
HevjggDNmyAT+whbRDIq1qrYI48Y3u/zLpbeRjumIDWfHqNk2tnYw3GZwyLRjm/BL6/gIeZloomf
E0jsVeQGZ7XsGL847p9pWgfwo9YUwu7ccgfJ74fDTfRKrevv1fiVM8XKppBsAfOxFrVldk3rV/H3
YmDZQYbhmvoqkxPLGY5ZCeiG3AWbusigzfHCibmfPRT13pLtBoV9OGXbnH4NrvU+3yiEGtDumlos
5Hzi7CEC0WR3ewiwKcvDFuDQydN22ytJ86tyt75eDr/OPFBPumKuzxtIIQTWHmqmEI04GttmxOxV
8BWFspGA1SXX2T0BwgRYYe46pPLkg/x0PinyAfJO83XB580kULqOL/GErATXErs/HPOoyesfH8Du
H/mFmiFtCs087K3ghHxN/kZrC1lzeKLwNz5AwpubJReVNTo8k0h3PAU2YaK/XI0qCBiv+s5f6aG9
eX77VvDqhWcqKXRkeHYBHjtbiVHPEJpvtci9nPJWsqhIqVknwHxNdYXUfldBoFISocy66uxqsCiP
nSDsViAa/RzTzSTondYnVEJNZP/BX5otbEG91ol7WAVna+rTVqc28h0HothP9HNTahlj9t+RZ4dK
UGoFu8t3Jsyf0PxI2LHNn2kbY5Tqa2ZXrZ9Z+ZtF9bUYLuAPkqxvPhnaVFx4h6bobUyJpmBvjW0C
1e3oaS5exVupcGl4FkPj5RapMxthhyEN6nY/GTq63kUs81XTyupoTWFUPDkldaIUAuCDoRNAYVlO
NKBmyfNP6IiEr3OKTiJ9QgUCub0HLn8iVHzBaqyxrZAwCN+Bad12hF+v4i/b0VVCIx2OBmECpg2G
cgo0Yf02x7oQOuRgIaWyrYnBo8DsxZ8MQuaRfBfycWxdVOwJDNBOKz5Yj8rjswqt88D3UvMt31CP
r+hHLxgn/jJoYifUKCs/b+Z7bPtEvYx1W4SL9oDf1yyJp+czl4IdFwpEwIKzlx2CJpjheCHCB+ZT
ut2gTmwNV9cd6ZcbuoByF0Gla76hHHpgW2kek0KNzkd709mfhtxv0I4fP6Q8Vf0XsO96tpIdIHXR
Zqm0zQg0XKoT8aWQNmWWHYwOduWzIs9b4FjCMaqqkpHf6vYoxxKkVs4EAlBrJbkncAoUkBonLPn0
D/adVsfxxkR6vkOI+Vl9j8PWAIBHjJh/zVwzAISTLoaoqHdORsI6zY3a8wPxCJesYy8RKT61JYy7
P3CoZJhCSb8NG4mvqDkEkTMxw+mKikD7Qua9fRgXhkQVb6kUe08NV50jDzqaybByF8hncwOGdHDO
XxByJZAktbaZTXNM2dHQBGioZQo7DCLQiboCKIdTO+sTtBo36OzB1hKNdGvfahwg2x+60nP1qN3+
ElKkJMJfhiSnPJQiYj/407PR5R4uMTgPPoam523SLp2UrUbK0TAgpoZ9zy9qku0RavYLVYJXvRV6
979EMiM61swE9emPAGjf0EHFHmeknP27r2n1jE9S4L31Tx0QCgG4S00HVO/zKBe6xVaEmlfCuFcx
0inzCWNTOy+F/EHKp9gKfurnsXqBrbkADS0CDIccsqsiKy0FJ1/SozKaiExfCZI330EupQgQRYV2
2zwLH9kMLn0w2Q/XTZ8biyCMIjkhZGkTBsOR2bcYcjLzfS7iYGwMjODpWv8Q6k9EUSidFUgA37cs
+SL5Sl+iU5UeSdgUsSDmLXJgQySQRclPqW5UhCh4/CpSboYTHLg/KolgWnhJIhLf8HMRtLOZ8nDS
q5yVcYPG1QriBDdyJwgsMkkKXC/bzNpmaaPVt6m7q0MedIeAp2MuAancz4XX9qMPaff2EcQunNJs
c1Evuw83VIk/Z8Y0bgWlXh20OsYc09ztICn7zKrWDqF8rbEXbx8bJt20z3U5fY03diO0Z5b7CUBC
V51q0tMm3ehZFWlO8M+9ag+PHi0guzsPEz4Mlw7kJA8V81QsoU1FZ83h7QW/BRduAXMt55C2L9a8
bh4e5UYqec2xnnsAlvFG9xANUzlJpdfqVOFH5a+xqz4iOsMGU0TgvUit6YbMfbQdyMe6eSqovCwR
nDZvWMNZDfYBTzTcfQhBpQILL3/PettYCQMK7aylkPPapheGnwtRCcxRbvmluPnJFz1d9N+jDcFr
gUbUWesg6a/FMK0LQny64+gddEZmltoraBh5omD9qF+jZukdLhm0IK7WGaKY0zJMIa2+zvzuHoQH
coSatyHZ452o7lK3+EX+QSPy4Z3L4djUov9ZNP/7pNCNLbZjUjoqrAKFI13WdvTXxKAXDWTK1a34
ubbIFeQlUfIHExGa3jh+bALy3R6GRSFD+jL2zgsIxUNQz3jubEOH0ukquZFZPvW03SiVjfeldGdm
/deffe0+rTOgaGrY8XAh0LPmtv7raO8SP4cWPjNn39Xz+Ymo27LqhlIzXvCluC6NfnPvAFdFyJbO
hWphuwjDFrx2zthJ8ZaTd1bU6tFCt+im58nsive9fUmHBwOWG7tpJmex12i3MbfbZK3xElop8yKR
Qt35HPIGd68Hgjb+2B2hyBmsoK2mtSkGykA4+eAe11YCWYFjjgs3vmxU3MqDCbVp4fuVY4AHfPn4
XM8THjpYPvSaI6j80Bp4f82xj0iw+kStF3I71lgyHWKFczpw5mokepDRrDOS9O1WN1xgL/4TrhtV
e+hhP9ZM+EDFLFvOVs6sd1GHHz3dfA03o6u8WLhguuSTBdPgKYbaP//GC7hDW/AacY/WQnqYeHe6
xRHdVMHIhrvtQuQom9l8vsgAMvfTDyu79mHGJRXadPxS8ewmSSAtA7N3rzSnx7y34cntuiC3e2wn
qFCXzkNWUF14meZDDiYPYjoNqBN3lX3hcT4g6VxrQsSUEXTUtbTIV6i8kc2xTWX6LU84DE6P5aje
CQJTCgy+n7Ycdkp5cGSH8CDzXHav2Ou7bGNzHgpsqHd1xO9seEFkotuZhBywKW7zaE4SQVT8tV96
HsDsTxWbRlM5Kf76Z3dxsqIDVCJbkOga/pjBYjHwRdK24NnTW61qSzgpK3iXFD2YXsBn5oQ6oq1J
TOOF/13QaTOuUblSeLNi+PfPvWflc/H0RU3028PK2cPEfm1Bft2N9CIaGpO6SVgeNx/26lCcVIse
weY4Xtri+1EnHNUxzh4F2CBBUcUfs/3j24Bqi+oK8+cpnBR+LeLZZrCfdYv1UnH4eoKtfXXDdEvP
zlpfq/GqiyaxkTbifwW8db+EDYRQVKprXIGfrlk98s6RYjjnMNb2BKoQ29euGgrx136hnobZ2Ws4
fI9Wee6uLchgwdYRZw7OHwDCuaMgybuHc4ngUhGpcTdWN+9E0StUhiNDWI+iX/AHfbg5nCwNrJ6d
KUBVa5TS+5F4qJO0FaHNDb8LAB23/11xovc7RFw2Mt43yhnZFG0gIn/nK6EsUpS84JOecqv1ObwA
OK6o69S1yhQ97irk6vHPzMFtXE7no1kPhIiwH/i4Nf4TjIJdzwJWeXDzT0nejcTUii6lSPRmyhcS
oUajm8H98VBm2o3L7lw0LCCL+sLW+Hl9+1dJWYZHdu/oNiaFNqSwv50tpbcq1UiuU4tKVGMd4eXX
O5YLWBoq2Y++1ARSVyOZMhpV2qb5mJ5ToLpKuLnuIu2BbDPz7QfcJE7RL5XJDf/nt+/+O91U7PYh
6/jSJz00bxN4u305xw5RAgdl9GUFLvkuKRXFqKx4IhmkG1FtCShq7W2r+31dtpBNSYuGqVxzEcq1
9ZGuvnXDoFc0bO5W7vfNegZoA7xLxbdHqfHJaAvxc1MgJ0Iw+Vw/yDVoreKHhl9M2wtczSQxn/tz
cifTgbmDwKM3zQ9i5Leip/en+aci4rgQzAKy4s6POLNfCSi1aBMbU5rfcZTtaTnPg3uH7MKIRioL
yVtUkySsSML/MAM+O8LOK9iTxP6+I01wRFzQJsXumDaj1NajZh6SRErXQVC95TJF7910nMLRB0r0
xybGzLTmqlRSNzurN53DU4dw51/b9AbA5GS/bo+jJLT0ckN68b9DmI1GmSRumlVGmsITNSUlm30c
ER4RAfhRmPufWJ7RL3y9izkP5GyFnZf8QUabywlAHmdZo+7Km8NhlZzfwzUm1KY3sgIAH7rLbu/5
SULL5SZqgO5zc891YNEIfjWYUdXlIpiGShqsnCuAtVGvBe6iHuDEymEZG8xU8Y5rHtku4pAUCEms
33waP9FtbfxEyEXJ5HPmQ/0ooaI3j9bMAwAnJWD2Vg4VTfPls4OC+K3IaVvtTA0eeefEQAFcnQNZ
tI9E7XUtfgQmbWWbuosrg0N2ChaW0joX7YjQBM5FLdQP7VBiD5LHGQaVSmdoUQl/AGLhZEumMcVx
h7k9zwE7mBRiDwUBcX39GKLquVGo8GUKnkK0hMxKPURQFkr3+g5nwDXGbwhaXoelkvoJL3LI2Kjq
iGeGD9D3zrSAGdYZrcNB2yP1vYuWZoa8PD8SWMi+7w3Grd+klPTn3xalg0FhbAENGgb/bLyI6wTY
ho7B/2yyO8IE3FAK5y7hl7Qs7a34DZHyznmc9suhKjl3VSa0F4bDPdjM5loEJVLA8dWV7Dst85W3
2G9Ks4AQFE3pCe9KtR/71BeMkHfCD4S/3o588+e1r8bM2C5QvOjBnsUoOPgVKwiYI6CRChtywZRS
50Wu+Em/N2KPIzEh9K6UDEKazjDbPSPDGzoxWpQLzTgIFzo7xPGZbNMtIM2qTkwN6sXJHP/3iGrT
emKxFEO7uru7gulqD67mKfD5YMd1216HHb1U1Gp7UMhBFtknelL/dZuTQnLCSfTmFUlJe0YTEL5s
yQIfuJ8hnEcoReGZb9OiVzNpPuyTj07zi0Mc7e35C05E1y2+KTjIKt53h8RNy4Zcpvo3M9jZNcm6
pEZ/qpRWzWpnC9NLwDNidUh3vYHYIM6p+oWi5AESUoFrcJSv0EW/gsOf7yd7xLmQdLHnRdjTt9P+
sAi67oEyCNlzcbsLOT3nQ3cyVwJrHE2LyPTHdOM/mFJHShaueWJJABJNZfKIJMrzlOB9AgkOzINV
EP2y8DrLjW7TcoLtkTteCmcHCmdIBiUREZOJdr/NiTy5keu7Ei6/4KyOxD7S4ZJcyXJKlaP7qj6j
ExFjwVh4P06uY0Zzdu6o+GzZEXS6CpNlsZZW73+7uAaVB8WReMjmjkaATBUYStBtOOgotUz820KP
H1AfbfCcwBSlLyvFrSv0c2p0pzIrA5yBSvByfsZuSPVcUFvbv/UATRHGFHBeYEhDAlCSTIm7etLf
PeMIbTHNxS3lok4tPysixGaZE2suz43lCJmG/c8aZyFvQ0LLjZ0sIBvNZ0K40P8tQQ0IzyaZCZ4b
Ei3pKDVBou7PufathCdubpdB3RTLIzcnM11sq9gJxZz5mtiAxaxjIeO8YM4+ukqEjbg0vdAiaIpa
Yldfqus7SLuIpX1INkKvDai84262d6/aocLmjR7WA0Kptx3sBz2MEGJSca74Mtx3M+T7e+VTex6k
q8mrlzcWzY8x253flESbySaK7PASazUynj2GrCgCuqx9ez8lE5D22JMHpfmCp+jfIW4kV6mQ9E6/
/4YCpLo9MIScf13MY4Ce2tLINL+JWD2kTaeC6LdYCesrEazy9XKnxBmMC/INsjEvJzo3HoH1gvT1
0PUhnP595TiyWcSqqzqygg9qnOuoMPksWtGMvmhz2KC0NaLQLDHlzk9nJSctXXfo0rvHL6byP56l
nEzPfNOZkJ1dQOwY6kscfDnRnOv8KU3ie12zqHP7WFOt9FNu1QZ6EQDYjteCOhDu/PLUZNg3X6VL
5GY5PsgfMgosirfYXNnoIENJ9L2SjVyHcN7asR8tpPiwwH08De05u2g9zN+63LRV8c9BKoDamoq8
d0rvo4w81n0Ipy1Y0PrJm90nbxn0kZI9OABFIYqmd6zrJ/uUe8IWysg5narBMTLeE7a/Yaqz2H6e
WFQ98UOm3WI7SMsO/uM36wreaHaBLkNs0Y/wW+ep3jYdjFbkLs9NHAKq16+quhCGGM/xcJ1FekSu
ZMaRaYU3evBFnazO5/Kdj8KiCrpeS8YBFQ+5ILiW8CiKuEvWyv5bY6Axxyxp8lHdW7yjvlIe/U0s
6bht0gZwSafXxXc9HpYN7N+1XElZ6WpeAaze7RJqQbZxvMHcoAYcXQW5tgmvOezddYyv8GZ6Fp/L
m0hsPkrHo4QSZtOWOiG0JbsiNhTSlbwUFaDwFuWmE2p0LGbhFDT6lFTAtshpwTBx/mnXueqeE3YB
seaXHSVpiW8N3y8mzVVRM90CFzy4h0xo49kzhUWdky/DPkZp0r80xKDfYld3vWepH4Da6QOERm+z
hGMEcBU9BqCeugeOmiG5f8ZoqTQstLHod8O7a9DWVXL0a8uJiVyCzis6YkOY05It7BwLvCsomtbi
9WCAhZxKOcq8/fUi3+5JI693MLuUjvkIYvX+erwcamUBU2JagdgocOcjSqCQnEDOfQkO8MbuhJvu
ySn8qGOmcWuvyNsLLGJyz5nPeO45Z7bs7J5O4O3cX7MTE9mC5h/SsiYuSInekiHZqIsF4xeXwu4q
jYVv5Z4EW39hayEMoO0NYtKOKvV4HT1Qgl89Zod27QkezGgA6AST+8xvU765PkApOwmLM31CTTMw
6uX4UccEDNAkbCuYHh7VD6AKgBMUfQqlDce2CuRCZ5f4bUkZk5wYHgmUC5Cd4FCh6bwIoOe789IL
mnqX05b49is5CcAkRF9yn60+gDfIt6fmLdzqRSaoI+oli4sIoITaPdlOPyCxZrTG3/mugTHvxFMV
2MQ9pY6P7sxEaaD7QVMLkyF11ETKHZTbVt/Ltm8wq/DoErusAD45XaFhooK7mGUrWvXpfblyZovz
K8/OXIX8O0d80nEcsRWPYFlp+aucqQzemrCQ5TFexaAfqsnnEFfeGMPkcA1QokMwvQ0UyN3JPInB
+Mb3ht5IOPTg4FY8UsQAErwofOX0X8KWCYeKBUb509oFZNHjnCxCIuQCr3agF4REc7lfWm5d/TCv
PBXbp6Dhf76ku5/D71R0sNEHc8n8nKggeoDWIkW1NjwwNfOwE6RjcDAMNb0+4pQlO/8IexznovlT
eI633G9WlVY9qbVTQ56+KZf7Sc1DwmGAOFsRiSmW02y2QfhJYSP7WzyhdnAlUonAEXR0lWnNpa+f
zO+AvkPOkjeXLjN3xtuV2NFe8sMrLo16UfMojnXhMa8LQ/LJNPF7L+ktRD/RKO3VednKo2pzIrZh
cv8gU9eDijc2BT8hKZBxEMwFiBPh4m8rV0CK5tvaZuXUtc+RQR448gRP5WEtxDYtEPK2y9ucTm9o
Mz5iIEBOy06J0ItxF9e8aExQcEUX8Kuy78P8NUhebBrQJDv+d8VdGNup1xPJmIb13RorKrm7OWDv
L+WV9A0cVspdPyRXAbLtkxDwuuljPsJ2VJ/fa3PDU1uxX2Oj4Y47LcJKZsLtHDI0qxH/c0qRaoLI
AI8JimwOAQ/azkdfrOU6AGLBJU6qvxHOcczAoNjjbDJ6m6gc0nR7NxAFPr7LUWgHO1wrG6dvhYai
NUpxxm06jOtuNEDyNpndvRKGabZnhCYQk49bSorBNqmbChY9exHjOdAkfDDQOCZhJHKvt8q9hVR5
UXqHB8FX77wbnuEeKQYrV8Yfg25hJizJO9R0qtlnfVyE2ag0ytgWUeaU4p/ytG1coYSVykwtgdFL
N/ABKwkzrO2uKtBh2PRu5z4OfOZpCjCuVzaOA48dAQWJnUu/NxtPKDX0lulM4NxMIwvc3Gj1MvoG
zOckj2N7r91BKOn7RhF9rZmzrZ+uwiW9hE2DFq/2MfFcPqquGfkbeShZbRpYaZOEwceRtp+Yu7wg
VhQx/k5VvYPrnYfKtQitodrpr4++TEx40Ao9ALC9kwpaJUCgE57SsE9Gokn4j+rDBSR7pCr4zpNd
pyE/f9Lm2Addbga/nREzfjuW/TXwMa1OZa0sPZkNa8Isfmr3AM5o92S9j9yeuMvEfWbHxC+aKVe7
aPAvhiQ/FpYlwcZSCC8U4gkTl/9XfDegnO8/yFwR1NB+bXLY1eQJvERQNleTdq7mXrI4yFwECgEe
MAMJf3EGlH0ALgZ5cO571CfH6B8ZuWGn4uUXrWIBhtC4vrJXcHWIXwlnvXVE90m69Y9FwMQvg8Bs
DqvpAIyINNECsHM2u7LWK760BFp8D6L6zwomqe3fquQQOCUq8SUHxlQg2n6EXo6wTYsvPk3Zsif+
cICWVozLs4jz1RxLlzKpNpxkcRxiBSenrr7IXcGbOF8gcIbyF+8n0mK8XD73dBMfGykNJ4dR+eEQ
Dpp5E4bkB/EIv8XBlrBHIAExC2M6ke2jo1SqZGVn3nC2w8Sy04NTOX0TNTXJLCnngD8y5TdnUFM9
wI0Gw0GneJNEPQkeb5+hBKedKZ9IIOwBhzTAPhuTJdArOVW/DY74EHhP8uQgCx6JRFinVB99zpsb
+QDYwK5mDVHZIwVgLABmMnVZ57Q16YmaPXItV46ACE8d7avmkxdiLW0lw72KBbOyP5aYwQS1F97g
3/e8dc0woQEA1viKbS5bUMt3wt32L8qnGw6FlrE5C9jxwBkOspc+QlymdAzTCJgMZjFur5e8znPy
6aWQe9UvB1fS+9Aeg+X/4o7eeI1pDmIJFp8fRDFzokaYGR1ItMip6fi59OXNeh5GKcth+kOor9A3
CGRunTjb0F6vWY+GjfT5dqn0hALtyY0aY/0jWK9BqjugEsfVNaMIyWshvjgQdjtWSqSTjtXyJueq
q9ZIXMxXPtagAsHLLgHMM4V5sfYxWHg5FTe0L4FgwUWIzEMYq1o0xyqz8pUuI+Pg75O3WzWxSp2/
4ssZ5bKgaZRw1rVt/cTfsRueBzGm+XCKIb8SpulpTGaSSQpUdrjtpSq2IL7h5WHQ3uLNGgHyYLh9
XPF6/S/w/55gr4gomOxK0hOmJgZVT4wVe5gqqfqBmrQeYYnnitNOy8B4mhNeWTg+/L6HLB5sGW13
p4LmqOEgSfPKELDQD5ZcjDifwpAfbhwt4ZirMmyoDLjFLAa0DyHRJBabUzTWDKQy/GkERO4zAMrQ
O8p0p/3jbAGusgMzSkHLWbRAz2zcpfjs2zo38hK2EA2T4EI5t85fsGfj+2FqMohE23/fYdnN88Tj
iaSLBbkWd9kjFgxSiWIU8dg3fefZoe5hOC75dIbA5hwKFMo/X6FFyo6VkcGSP99mBVwLsbuqxV69
2WWk8qV4uJCvRrWyoqNd3MUGENP/G1Jh+g7BomM74ojkZbtLMvvjG/1C4JwQhlg1XV7ICstFVev/
dH3IVmLc1VLo/x9IpKk5nZwzv0tK607Kf/J9DsfumCf0g7fkRimW+GtdGWIF3+Dijycw0RpIJkwM
jC4wPUqaqA0jdmpoPNfLIntpRuVSqAolscPB2ZC1ITvDbo0jMmok1yuB0nUJ4x/4o0C4o5mXtWJb
R8BAATe+2HkSbQwjzCKikDEo5DISE2fW3yxLrGQpHVbybRfsKm/9k44IsC3FEaLuZ5dYLfHXmfXa
emAR5UUJ4clWZgNu+NqjIUhO7Wsro83+vB389Y4RfNZzhWp41zRhuh2KdaQUMLkPkSN0mfHc8lSd
kHzeuv7ZrNEjennJV5vYgirUrxgCohJKDMP2jK9nwNafQV1Fyfcd85R5anKgijEecy4Z/hbaP7bx
z6N/dIkdZ0wCv+8/ic72IPO+W2KXG8Spr0olSj3K7amysWOkcoZANSpFc7v3GkuoXpftYs/SSY2m
cpPOlWEfbYkKW3GtVuv+dp4Gt1L6djU37qctMGg48gug2CpwPFbMZ77YXcqXvuaazNfoB8q50D+S
cOfy+vMpozPW2T29oJdrIg13Wk1tA2GgXRcETvY5ievp3Q0r6XIrB3Y/3QUXJ0xROGIkstXRu/tg
I4FzTNde41MOeoN4EHpoGEdo9lLxpzj7nwzYg0jCq1Kz6nGL2/y4VUDMG4n1zjXljfNzr152f2FL
nF8TvBI5G96/iJeZQidjc+TP2hMGsa33NNdlx3i0AWiJURGSdmTPMKn7pMFQV4E60qED59vbW7D5
QL2u+1WRv5fgqMg9Z4DJSizhiE7PAg3tCcx4yObqweHXlktLjMZMrIflR+u8u9h90nmuf5E/7ebm
DtCBoj24qzymBKog9bPHBSsdQUvkNTPoN3EO5T4PzwmS7UNTbbR0Q9aXATQ+FOw3vZAPsZTBMjcx
VwrY9Ywxd5Gf8v7XFE8VH3AKq6onPHqfdjY09b5ZxPovl6grEzFf4oyQwHN8h9LoigJCfCxyv3Ck
kB+0MAUCRk8gc9wUL5e7Q0m5wQ3ktEQcdGYHjbtmGRtoAV15+yaRtsibO1Wd/hha2xhy4FkF3Jgp
+aEHNYGb0pH6KotgJQA+p370gudfzuLEY7IwbF4ghSOvFijPZQ+TYu8YgQyKWdvHt1ZtiMag2KLK
kAIX73aq4NTO+xk0YpsvNoDQjdPleV141iRsw352OPaK9TT4grKkdauYEwmrNXkJdgOZSoYCsTnj
Dq8tNnLgoAlfOFYimDa49GeAIxcsnB3VXU+SIE0W1jz2QYi9dfcMGp1UdRuBkbfg9kDQu778sbNd
MY0DtXBW7S82Y+OOEZukrbgeW+bJqplBCbLO974RENSNKDWvx1l9g64Q38BcJfpQKFvaoPdGE4Pk
5r9RVMWWhtVC3qEtEWIpCTgfU5AcFjV4E0rNGM6m/RD8RELk2hYHLCQ3KjWlkIb3vUjN4ewQjbDt
ixRHv/WzuArSJCCo3OO9SIWizGUYRjbb77BPyfcZr1l+YIyso5EoSpSWapwl9xjfkz+/YHjN4yQU
WZMhcglQktjb2oyaMNc9VZ19IGuzc4UwCH0Gb45kD9bmPmUr2B/OWAf5+JdXc4atJGUpS6zHsPmT
cwSSsbWNam0zLYW6hP4il+EZqhMqNC22RhMZXAAympy6SrxruC8NFJBLjj4/pSY4g7WCT4b8JoU5
0074ImrNDGkbc6m8FptqLTMh+q/Lin1XSgEyc3gGH3R8xwnw0WrWNQqvdH+/66O8ZFjdzZeyqGSO
qovzr/4pceIxfL70E69bk/yBvq3A+jeCkHoBt58WV4Gxp4YQkud08/L6bpn7B97swtuuVG7SAf97
opfxtGYDd/Co/JUwi3JHzsBq1garvk30E1PpcEa81xXkKn8CZS0WqnNb0QubNI9wAF/GQ1ie8R7j
7YWPOqqKh/nk/tuD9rVPCg0+ATKqoeLuKxW7l63Vb8a/Rhi7BUVUeFutoputxIk9GV194+kZ/Wpx
PSkvexRXGEOcn1hQXmFvoB5aTs+Zk/NoyhW7Kkfqy3OIlSA1ZLIpxaf0BZw/on+Whzw1oM723loD
xcx0lOMVs8bHMSRod7M1YPHxCqikQZyT3QVu4ajxZtFvxeP4J7GlJceIU2lOmY5DONx+H7h5EF51
ee40WLoEx9cnsQNXzeYkX8WboKtY9KP7YldOpKeBBNUJKT10upii6FkQnzw3brYRRNI1aKrUaz3m
S3pU6T3F1hqexDhR0gmYrI51S1bapxh77FhJzwZUicWyXiZPUw7PDIpH67BFKUsYsAoTJAeCw9sw
7xq8RUP5xuiBycZKgNAlbCtrU6dgj8t623J4ASWDVDokX6LeONsvuHRMH6vArmRdrj2S4zHyHvqt
XM1wCWr3teXdvUAbuZ2iXExbE/iZKGIS3kkJ14Yg3zrmPTLXomCZQtIPZv3JYaZCUkGLp1S3wCaG
dGeW3B19TqTkNT6BrLU0TwShKG5P/mqerYyQP/cSEDeYnxCNfhSNEe3k9Kn8RT1z4sdAYBlfBtqH
6mkAjmPdCCbfXNlqUJ6p2j1FKPuGpCHvI1fA4eCWdInuATTJ7kRUIwwL/aY6ubg+8P4CfXAVtTVx
ZnNV5YwDE57Jkh2DaOpxNzglFsaPIHU3wSCe7Lbgh2+A2Wc+54S7lf7MjS0CLQ1hMoRtgLbnx8Wu
omXd2NGoKY0mHyT9dt/nXM3ZM0ara9rlp1lJHDXpRDUETjag1ZPImUHYzskefvPYpElKjrcN/GG3
jnm5L4KuMAxxxXCvqaUd92q3xu31qXOr7BiprYaoyTObfnharnMxnOQFCMeLiHNUplbBTROh091E
ByVapv+w7/V20J4/jlHhctmYxa7LCPqWTDF3GpAji8IH76Zy1BkDAW1iPOazIqMLhUDxw4mFsFJE
dYgBiNIfK/hDZ4KiJmA64PC8U/jGolu0MZRO8pdsFsyVhqMzwj/GvnNtHrtJHf8mr6Uoz3jKb6Kn
lSsQvJ/gQUub2Bo+9k8GNP2Cx+a6S9n3i2UFdfO5A5fMVYJHmYiXX25hMl/ECDb9QvxnoL0snOX3
fce+KYou5BxsbN0YlM6Zr8KUxYg8XoDmJigc9sG8eoLII8S1FhdKn1tEJZd7kv011PwdBFRUP5sl
EPx+8VAcFwBnONEXNd1Dbg99pdsY2T5EvCPUsmc9wyDUxozAkC0y5qqzCCwXect+pDpF0N6Erf3V
8O9twVF9yzrm1DMLWqLEDo6tOb2uCXbc5zDjtU0yy0t50TWQ2IkAq9NA9r55OeWapkawJE1N/bsP
x0q4omX7wHdXaEqwRfjXiV/2pLphUWa5x7YKkMorUWJcnqAKpf8O94itnLVSPvAN45nytMMII0gn
KXxCI+ORowi4TtVrYINBaqx+7IToi/SRygpUAeptJKBpCT8SRnlhQyUibJCHaILrB89KtEYx5MJy
eVdjHYJMwTnPtW9GIDXsfC4nhQUes/znzz5VXX2QvaGgaSx01Qw+iHiSWxFbWHeCTTrweX7CrVsw
oP26oI4/vDaZShtEv5LhWPqx/spjLo0XNajyfCf5RHoM5vAl8c5czANAPzuZ7Gldz2LOUrjcM+jI
mzmCkAT5TTUYcqLN92IuUJDLo+DWk9JhKAKjCaBjVK6YJSpgq70D8tsQWSJ/GorI4H76k/UJaxb9
BDU/pqM7WjjzkLyW8DTFFASq7D8VQyr1Hv4CAgeaM5f6rUbw3iI4moIB0mKZNOtN+nOBbBplkjJo
9eRKSZQTeWBA3Ld7OnoExAKFiBVvnDZI3iVlXh3I161DSYjFC+NmAgwQsIMGGlafqBVA2PCHauu1
r94JE5b82YFhT06UBHmhELYfmrlN+mY5V2aek9z6nNPRypwGJD+QP7Vx1WnEZBb0iaClqIzCnRpW
Msx8tfgIgl8UYtLygbbYfoSk+xKEVJ7XSyzkqCNcvuC74+Wq4NPVunDSptA0+cStmfL+2kDepaRB
ALXOwByYHieODGpFOTDbzKCxl8Zk/IYP95txXF5JAwtHSOXfnU8r66l2Eo9MKD7X6x2nx/fvWEdK
oD6G2OZW6k6f3OadwgCKAiwmm6ryQK0HcYqaREtwi+24xcGTgV7W+kjpx2MP+uh0OP7o/+uV5dxR
kT5SSkddU400/Pk3spqt2BrqCgP9hE7GhBEXTQblrZ/vepcAbjMu4DLs9hNb6wfZhKLxJg8FZ0Do
ePdqxPnD1nWTgVvFJ/e4dO8DBuKN3Q6FdudDsRydJ5RDrt9mP9YJ32CXIZUhLorqC+rNL15vhPKZ
Q4xQRvdeyC1MIGC32I2FGE77mTAsWLNv4xy5kphjl/fl3xd5CZOTHJWASCLlv+Czg9xHQ9Gs5T77
BQpxgAYCuWMJKZbBUnTEqfDhrk3CwubA9KELAruoFzndjmmPHOjFs3Gau5GI56+nLhBhN5qAFBwE
Y/rQihyYxeS/MjjrIGhCs92Tm0F5BWo12kKYRe9TssZfs+Ni+gBIlXn2v23CuqhQls0wyVvZlKCv
OzZ51G5CLP3kk8hL0oFcvIHvHuKQVw0O1JglHLbK1qv+awyU7380iwm2c5vK1xzaWmEtd/phvLJd
1dAf7oMcKwPsjOvktusRdj8E8vudvcsyHA4NEDhc4YQCPO+NnH2V4d+3j2sEEe89weKeA/+LdH2l
iPQHuD4eTt0zGf9PH0I//w/Lt200y6mYtTY6jNQ6YhFLO4pIQ2yAMSF7BdCZAMxyQE7Bzw8OAES8
NnRZ5Lf0zRw1MrFuqM7/uiJTByMJiAVChUceS2vI4LJubmCKuGaDo/yF+of39oOByqDFzIieZvJ4
u/q3Jz5Z+MPujiwd+0U7xvVTyRlPhNUBifGyfLkFjTK6WX8nyVgRH2hVc4e2RZ19WpYg2fDfzuzi
RACw1y/DSaO6y0WvVyOfsMGBxvkkzmk8LeXLr5qqz/JkYLckuP2WJqwNuk6zBoIGJ9UcsCxDe3kw
YHd+ZiJWmiIDMhWhnD/eAgMFGkEceLOOddLWx6mgaOjwWbUbyXji20JpIsOMqdyVkInrPdCIoKJL
zVDI3wDRaYzgXkUILmPZBARvo3mkSxPzxYabjfhA6fVks3X0SIo5XGe+VcRRUEeqgZRcKtAG1X61
qaU8f5KMntrFdJwitHmsIA6pTxpGsQVyHnerG+04FIH2ocJMNWnYiWWX/PAmBb9EUiKDtkqR5JYC
Je2rckHHQxIrOBE8zonA5cNqIqFYy6olsQX+pxwliB2cEMCAlH3SwN7+gTsbtC6eZEEtrGYmhMfh
6O+IJrmGZyweEBBrLDlSaKzDTCJuaSauL8e9Afmg7eIWRSNJXq9ZqBm07UDghkkTYsOJ1MRkcfgP
9Eqr7KzDmSwE3NpWY2IHlNYkolmE9/tedFV4XYIJ4258n8Il0WDVms1vEzJgeEs74FsKJ2iL4HBx
R2gDYNI0TSFfwWrqwp5xQQDgjvaW2DQ1akKraiyNJoZVXVPwnlr/ioUbPjG8Md8JD51G0B2X8mBv
e6cVoiDt930D4dEvpP4Tqe9LF09Wmkx80pq3wuiNhvQfUq/CwWB5bff5QtPEWf7T46gXav7Ri8RM
x/OSKiEgHgwZ3NGEk+l9OzYwp8Y7RieqGJEiJEiOSlwR2mZEPPs9WOTMxATcrn83VrklqB9Umdkl
FbtsJiHgyMmOVR3CJg6XGNaudfMbwPryvG4UHfk/khLp+wjmH8PWt/swpQLHx1GFwEERc+7Ifhh2
QLy01yPcaE7PphaibFTa6gsaMpwCfbjPqFls4nYa01hkwwzsMYOFbOm9upqFZpzSTilmuTzOJBQ0
whpsFXPhZXqnfW6mBN/LlEYaoCkfcr/0uMSXsOzxPoOS1rQWns2oQmKghYf72DHAqk2iyQCb5QD8
nCK1iqV9Cd162RqyfVnMirSeBhuyEg3SYAahT60FNPciheHx195Qv46zXYnra7GpPTAp+7ggqJMz
gkEv4FFg8hnbk71Uak9maYChFx/nDBvtKT1zML0+nW35zojvgU3G9+FZP5jFHmcixtg0U1Evh798
pJkD4HBQp4cpg4ogsxll5pnVSitayW1PmKo76EUZ3Hdg0YZj0dtbTeY0y2jDfGXM9wi1QG2JrPWf
fCERxikEl1LHqnBSDU89VIX5NjYcG6gQne642YWNG/v3fLkqgAd4LFj8QLV8zv2O7BBKvmmEnRnJ
h2Ul/mjh4r4mp/2qeg5LqtkzLSQZ31wu7RZRRNl2PrVu/sp6QCBFcv+dkQzM/lJpTaeLDVjwixGu
xJEc2m568EV5JBq+t2NkybDWCtSTmmrbHqVP2Ski0IUbRYeGAw4gEIFcNCeI2+RdcYO8CS+CByiu
z0tW2+j2RvFy/fiyLQjSN4zZlr4axfJ892IZU0fHY8NK2sXQJIEznrz4GNd6NPPeiTR1fERJXMxn
5/aJnY+aHk5Zl9xS15vpfVHKE6HU00ip3krrdrX2lF7GHnrPVP4bcieeIfVTDvTjrlUVIj22PDqV
FBe/xEmVz8d1RmGR07k+DY0f5t0TfO1upkBADH2RiandKsSQ3dPPcRSQVSGY8ftpaVrliSzR3Wyn
cQ2YRsZ7uPxs2MIMcP/no2d2nw/QecQJFTizDsucWGgtZ1DAkEfhP3u0ZGUCsS3BYILrDUrN0pHU
si+v5YPDhaICkK0dyjSIfPrn8CgehAavaobfw+NHPwmzJuHvBzYp8snUJjpr+ca/06tn8fQMbodD
heaul1KZKW2KXYC/eoD6UIdckRI5LFXL5YdrLN3UYyd0nXevCBzMY4o/naTio/48ljiTnCMXxUey
0wvzMktprvJbTRCsr065AIByafh/S3RI690YAmliz6BvnXtqobo3Gs+oetXMcK8rPGI2S/APyKf4
2XTg2ng32Wx4kaMIjOMxL5KQQv/FQI80gqgtCSrskXjk7c28JlFjV36FDX2dkxJt0opfy9JrlAM5
H5pj7Tf3wF0QEhfqEm0qeuX+y/T1sLxiOov4vUxlyWKo2jCROvg2mOvwPGR/QpszOv3WoA6yVJfk
rfYNR4yXUMwFXuZWsiSTQA/QTqTdTKmhbGnhJBcOdZ7gjmBlPxGQEoCnj8LN2Zqg0tg6d8nNVj30
XUsqr4vUfbJTDytduFKE7qB3klqAgb8aJozQaRdYwv97BWMd+zhDGabOf9cXX40ju2UET7Mp6+rA
KgYpbh+ITZI/jTOvC4V8ID+YdjcCDIiqGiVd9+u10gAJtfecwCTc2t1ONqIoCawkw/yx/Hw0cFnJ
jPnaVtgn+vyiCOWImIck397PCYUTdQisgO4XY17W+RcavsQftrmrjQLWoYg8QU1FU7hu2m5jhNHT
C8Wgv93YiD+z2G+hR0ln0O8gl1RqiON6muFpo1ZD2la8noNCwPZUkRZt0c8BbYergup5xjKjSaYu
G8XSyDxhc4Zq/9yavfYZmTFiQnCmKvme5TxmkWEET/AkAa66IallSvW9s5QR67zguOcb3uZyXC66
CQFQ6t6u+mpEdWO1ehK3C5B8E3cOd1e6hggkqsTl/+70V9c+TBN4S3E9z5oxl+JwTNw/0B+gA4tm
YbzoCs+gly7Dll0ruCzjPNHRcCFZZBzbtjAtnLQINt3V498w9vVc5pfYQkqDZ8y+0earxaMubdq8
V1Vb4l1NjwsB3tj/vBLHPPeT0E+KHZ/YtZyVelQYXQaK9xdU4Fo4ieYzZo0XvbjtEIAqmZSBVXM4
Qp/nIx8M/FBUGDRmjrlmZLFS4q1eHG9WR93+8jVAiRDbmtl4wFAZX5UUgx3o+tiTXNspqngg8Ymf
YU7/WDW+J9Fggzahb8JoLNxAmRNFlvlam5dMbbZpO1dyP3upcJpq+Cun2SRZsWJ6Fsy91qkkB2r5
NOvBzmZ9qGIS3o4AYostBxSezIh3ky7DPJFYN06lCvteE2wXFPo/3CTsu8/VF+bZwVbepcAw2di8
pf2sIDj2tb6qbEir+tvGbt9WpVO9Uq0zGHLFXkXCLi/viq7SFI9sF2l3GHql3md/6DSS/L6uOmMS
dJE6wG8rTeswF9hEXnm8P3AODlGGgWNMcziixGf2UgYzP+Z5RzFdZ7yvvpDgygoy9eyT5/wwkmCc
qxTkz0JzqLDwA8Algw7NjgaOrfZFpVyCp7W0kn2YtxUpk65nQzzkO/ZBmMqhj3xTRf0DjzQ4Ojt8
e6aDe9Ux4wzXHZxXloihdPoCnKGhsMMikQ5a50UbT2ylrCjIh5IcB/XkdWdyfvaQoPteKb1kIZXd
Cd8EQo+B69iGcswl3tiEEfEV0OnAgn9mPqyHF8IZXcb8dm8T7InTcUip22Gx48WxTb11Ho4QnaRT
43XkB6BC8+LQM3SycRdrzWotLyudGjh4t/wpvoLKvwtWPnaY58KQU4EufGlycZzcXoiGsbELEf8u
31darfAphq2rAfmbnOb0kn/RKA2q2+6vkon1ntw04rrnCmIvrLbM7HGdwiSg/qaIiHYvgOoh9orO
6g3bv9n/e821Hz4jHAJbe6LMwNxzbKlkPvCAEG00BdldjY/TaG4DettrsL3ZfSbLhbfv1yoerU93
C93K27ZNiF1SJ/YXWiNCjTXR2Vvw2/DivTGCtO3yM28M7LqeE20yFNM/6Z7fC2pYIliTj7bfezPM
kK9p4+YqfFPc/1K9ML2IAzQN0PW5slbBUGPFoDl6E6vjk8Pabbp+IO2tG8NJ7GiGvJftLEjIFQhk
rP+z081SSfs/OBA3PBWJoP0SoDuLcmRvXZNTiPn9T/3K323g6JV6OA85SBgsHhekYr/HCsN2Ft+X
3dNx6FXAmI/pkniYrS2kEKa+A5f1FIog66G9lRiMLhlRsEe00y/N3sv8PhO7isYKDYgoxckHP6ek
FCrDV44uBUj4Zi1tDVxEy8nO5EFitO11s5GsAe3633nuV4bIiF0n1zHJSgzVY4TWsAh6DhnB954U
VBOxbEc+vQm3Fic8pnmUe6E2wCLP2bMiHCrCq3oFEAi7SeKFjDA6dU04BLezIenXvfQH7AaG4xWF
G/iyTHdW998Aq+DcYngE33sXJzI/ka655pc5wVB7DSIruNXzS0945ZhTDKZsfyl2e1WKRH+q9lcJ
pDohOaOuLJiyJLau+JIMIr4lCSpx6eJJ0jCtzKeh5QrA/gCjVKiAcE8OrAHyoOQTTI9WF55WOcRk
Tbc2rVD9SnfORDnhmzNe45z3+Gh613cZboZ27rHRrz+bR7LH72aNIKRbe0duP7qQWQP6w1+KsXoZ
4Ds8cM0Z38sIWNufJdNcb9Wvcxj/QTuYObTUTBZpBhNhb0WqoLPqxnqxhkj+jecx9jYg7nWyCwCN
FbbwwFCKEasgPPyRIeAR1hqJD4KCD62LSj1X5JGvImZREbpsdM6tFiCvTg3LKAV6VWJZbPUyeOti
3tn8sEckD8SzijIes187ap6JWtHHdiGR1+2wvx1uNVgPhwYwD/ZiBxZiECHBNL9RMXCpPRhpI+lH
rdeUQu93wV1iEpGJnSbSoVs9A7H5I3yy9G7k0fllWoucYhyt8pjDW9CsypDFyHVUcYhnS4JV17oj
6Ah9Mif1fjkduZoc9oU6ef+M/Y1Rm7rHjSMw/dvScdyIgMmZ7HJ4P0/jiGtDcDg6AXGz6XlOpN0Y
GI9Piah9+lLfBFs9/xoO3nRmN5sARb01+2+kUURdBPQ4dzHaVdVBZrLOawBU8O4NpwCEic8fvANa
RAzngIl+QXdQnTwc5uy/63BYJrfyT52cvQ9oFAG559D/ltg1/pjXspAhKZ3XqQgr/eVZycp9MWUQ
NhvIoQBIBbPCV3i1ftMcW6ApzbRPAAb9QTlLGzubXUqrqxtAlpIE+oscJQlQCwvvPzMVoydwAgxq
fAeZyCiXFPUUlNr2YxwiYEoLcbWylB8cnNJjmjI7tOVx9fWxQ3qXkIy/xaIekCRwQGIqJy9+rJSv
Cu6PXeCtJLh+0i0L78O+Uj3BJtEJ4pRiUtTlmXnaHw6/vD1lcdBywZtGcNciMIyQUnGxQ+cO7tmK
pZEmroxG11xc++SCNgavfG0PInUM0xs1d5lw+k9YFaAGtVPQhT4mBU9G9082DZqbqtwCP+0kY4AM
Yfe4jjCG6N4boHog6W1If/J/p7D/X2ViTAAj9TfiS7SMyEM0Rz/4bbwlSiV7ie0jrfVeN2zUYfxr
vJjdFEiaRmXqMbAl6ANw+yJRdBYIJrAnwR5h5GF8BJaAu1+RKVfRlnndItRU3OTQo2drB5yMpWaL
v4FTvkPAzUlQVM33Th2sN7pDHWdzlusdB0jfg+uUeUUMGB4mNgmLiJBOu91uKc9CmFJMzbVSKmZD
cCehtfUWr4QWZIXrl72u87l13/GkBaMLJYFYLubudzFv1cbletRZc68cWGDPM33+f/U48Ud9Bqz/
M74wRzX5G9i+EZOMNAVSl4PMnW06XBxxzCpIIrqjE1UvobJJnqTBUkOX8NnEXki07CHI2nha8GL9
Y+6uGhytFtYapYCjMhnlPM/W+Thh6CCjHwO+EjLXKjRNbaTHE+WztShqRtl6/mNfwNo1AiiCEBqp
bLLUKjbK6KAvIms2NbVanECaBLy9dzSOsfpCD2A3hgx1zR5FsWWPGY5/3R/ftyBQydVdur//riuZ
ep2HfiuGqocblaltLkjGSQLz9Fh6I+AG2q58JY3GhvwgIMIeUijVi2tRWadSQNHC7DNhM3ZvAfa6
5aJHB80AdFJCKHlSXX/OSdxtdvSlg3RPY5BO9M9axkbNXb8zRubVN0K3ndT8rgWp6sPxtVL3vgk2
40Zqe/JHGe7BV+47IkqH9NzDPqsfFEQZrU+VsmlvpGisG74ly6tdt8aXw8gEtlELKs7/J/OioElh
T0djSByFypH7Of751+xSykz0EuX4yIOHdr/rIQRi4W0EJ3hlGyXxjSpA6seMXI9QvGRm+JNjZCOq
+6xZoe9iLhUgYdKoy9sU4dP3tfreSMHY2QaCvng2y1zYef1ioEIBspU5tR7GMqWRk1NgQ1oBdSoN
+uGxV9S+ntI81l0EM2wzzL81+IdPlVMuJ3g1uK20j4MD0hDbpdYWK5cLke/JLBSDZ0Vgq+psiUtK
sx63wZmQW38s2gM2NAoD7ax//7eCyUz77Ygc/4TMUTuDO9+St2Qs1JEG9hBwsLqU5yJ3WkyTFKca
Dwq7/xCAlf5+jF9dQiiwemXRSmdsaxw2zbtFfLU7se5yDA1MA2pB3DLKmASXAtObU4cVe8fcQj9t
7GaVSf80BQ3fn2DViiW58Ks1YJqHt21GVllXY6bbJJf1mMs6wXpnKNMmlvAEP7892UbcVEGv+57G
z3trZGgCxaOswJvT0jHLkJWQ/jIfbSOzBWJZX7Ora77j4EbDvkHrvfjEfV6NWOy8N7kszwJ8+XaN
8Nt2YARKfH06Sf/uQdr/1+Q53mQ1wOQSxT1E2RangDCvm6RpA4fUPVjshVj5B/IgzdbLKPwsXXd8
pIf7UkE6cjvSHL+4ogVIV9I5Eoglx2e7BqgZ2xzL83IFUwgpNh6O+FWf7U79HiKD5DXcgjTMrGav
2ROdhXU2AfK9xbVI6jJPq97N6yXMTg7pwxj8QPf92sbcdheSyTPExH9Eq6AFSQnuWYkFxzW6Ad2s
aAfyYZjkP0MVi/TIjNW9NMGlnqyBuWj520zpds81St3Xhq4NJAXmtGX9DAphnHvU098yH6lfxTH1
YdgoSAQDnbqNl34YiJXLwGvygQb3GbohdzTWPhTO8Z0Fd7zz9aaHjz/tXOJFfOIdJn2nvRT7xBxK
6gqpmA2gJKlUZmhc5JCgjseQuxMKzTx6GCee+EhFnA45zB7agsgjF2s8cZYq4uuuobPgQwsajoVP
IUe32av3C9jFAvhTKHeg43XEJ+JeliZDCsp/Q9Wc9Oi+vNeJ5TNAo9VitHgVBZiBBm11WE9CawXd
36qa18DLueDBs3sb8tkjI4amnQRWDrlYeM2qq9pyNtdNl+Jf0XKBaU3sA7hm0P822g/nKyNZ82OK
FoKfiTWyuy3uSKupGnUonBMYfN3RB89jTt6FPAnq5htg/nr5Tw7ybU2lxPd1KoIJD3JGMgGut/Su
aTDV0fZEDMKIGlYNM8QAHYTLLZyUlTA863VBWB5bOryMFH3/MW/pCoSzjv2nzutHv6F5ZCMiMAov
8NghGIuOwHF/gPrWPk/JR8FRmddVLvyi3QLHA+rbA5RKnnOCBbzbmsTr+FPLV9KnA8qrSaaZCcvJ
pzYiyCNSm2RUsvrAKLs4HeLQ+Ypr9QBpST/llYjjjM3yx6aBTc2/anAEPSCq2zP/gztkgUlJuXWg
uuV6MA/GamMP5uZ4E9M5rkWp+eA1jdRzRkYzXcu9BJlrK4/fs3pzQg6NuSjo15arPZULq3MINT6G
hzv03oSTSrgBa/+yOGPfulp/SJHkFYEiPOix6djzD8PUkWtaMKmaHlmC2J1bvBxolA/kMzC6RfiJ
XRWdN3Rcuu+lupSTg/eou0Bk2GXO3mdqhourdFF/vhP/wnvaCmCNQqye7O55DVqj84gC2nbDCrNn
CwUsZgwR5Vc84ojO2uX3nH/PX7am/m7rDmrnpexf3Ku+/e4K3GIlngNiGTFMonp6t8NfMnl1T/Nb
gl2ilOLWCTjpZ/VXRVXxbgEwobrW6gcucjAAHzsHnAwmQ9zTjq7c6YtrHQTENq7jtuZkiIciAJqr
xJrAbqyjHJtwC/kMZvSZAYqel9JZX01w32dH1moCAmwDiFAYheVxkvhZQps5dINKBBo03BxQq7Xf
OMIxjGvQjYP7Il9q9mHE2u3xqhXWuQMRxeKI4K5XeccmTICp75jUaCFRLZR5Ke/n3QS3aK1Mznqq
BPSPWW+pQIWI47TOyJtW+ySjmxYHr8bqM89G1Cf4dnh/5oz9b/EUfxvI5fb0DzJq/LP5CJJ3iuN1
njknX8yLtQNEjaf8BwMdn47/rikoj14XAy27sr0kUyOpVs2AoNaPJ5uxz3NQkRVUS8rUWFNISUi+
1Lt+brDTBhgmhpbh+1gY6rm4iergyesM47ruNnN+f6YU8tLq0c2KoT348DN63Mdzg/d0Uqw5lyJf
kFkY/AqPjDJ+26zPYo6tif3uJU8XrjN2A1qWh5LI1qF0UJpnwW4cHtNGn7fOgO/z+zyWqURzOO78
7Aa+SyB3cGDGIzEgMOlqRei0tmgiaUYO/k4RA6UU668gnBjtU4MfqWHaxp35bW41D3Nthc7wBqtk
L8uqT/NHqfUBUQsrNti2xpa7GuZ7kG5efg5WOxl0tQBP+ChKWHXlB2hUZKw1KoWLiVrWn18vXUz9
gVkd+1j3688K7557zjhhr1srPSnyoOEkU5kiUZQQqegrO6HEYUwIEbksb1tuaFkTmggdByE2nhve
YBRIfBBKYHCSkv2jP7TkWllOf7x2CoHCA2xO/BKB3knKifHf48QRYAkQJQMBedn7VK1169k/Wu7X
fJhkGbbOWa/Mv8skKehAoKVUhxuKIcVCHEfoc14oLmxuY5SfAKkj9+E127c+6nY14YzhIOkRsxZb
iqPTyXeU7VKMP3VXJLiktcX0v+g5Khkk/oA3tjyQoZrbFzeTwGzMmGxrf2z9mS6dn1T0dvtqh9+d
/2/5J+YYjVALNQ6FZ7t5LouDM8y9ucUnCG4bhScwat/GBqxjNBNMzrIclZ+p10H6/Vp1yRCtirPy
KS725zQ+d0pMksrSUKhuLKI2W14p/jKf9zZUsJoRGsL5yLFfxSWLBLQZ0GLE9oaP4MiokwiTYU5+
s0reKgE0SdnBEK4dh26/hKGw9b92uYVMf+OYZXF547266UVuAZ+RmznpokuXv/ymZPACDDIXvNIM
LxjUHyeTI2vyyNN7p+otEczcBPPaVeLBtd7CGVXXrCEy+2NhF8VyZWWaCq3ucf8v0f7sICFiHH7F
DWCEBteERyjVR1fNzU6QOH3QK5SbrVp3oKSwnJ/bFuku6sQqlzG7uNFjyHM8/gIMrUsNatZwgkzi
aljI7DLgfO6LG470vb2Wz5sr4/wd26p+PWuBr/HI8czPHa/xCcfcD3IAFYu1XVo5jNlIhKLzFblh
DnxILPQgqNgPjIJGhzoJW+MLM2PmtmWF0YqM2NWWldiQICOMmGg5wwiIJBWOjnFtzA9+itNaUMLW
Pn0NZTK60G2xtwpprKszT+2WnwA4Jv+9FkefJF0c1L21zk9J/jLmfhOk/cp7SB9Fl+Gh9L2oVv7W
sHmFTHRxS8YneChw7TqAOogg6wclOcVo5+7D9RNxR60YWO9F0rOj6TtXdX4W1sMQywRl5gI2rv6k
NB4Izh/etb4Dr/5qtSzAAk3XtbQ8W49Qe5cncquUF+EQvhir1+80U1mb2nyth7q9vYpAYFV+A6lb
1PvvXqcfNJVK20paEtumGftgNZVXiX9Qjsy0a1oPtGUPk1dyM3uwccaJt+lV8Kxhhy+yfhDGYBgZ
4vYM2VyhoiKxywNPtFhOpCYwS6HbYtJIWKaVfbkQS88mpRvSZJ4+7O51jOXnYxLVUx+0mGREzDlh
n7vg/hQ3BNHIsUE2mLNLQAlxAA32MneiKwhb5sS2OKdV618gy90iNFFBzs4HdFR7noC5NEXUe+yP
Bv7xs53bihjLMsWjdFHevU9ljr+e1lEIldGGHORF69/vPf0Ke5EWgYNm/9IdeC0Ij4XPpHVC54mX
bGFoKv2cHsb+FLiwWWGM9cOQoPBRCn+WnbkiJ/eIspgODqtsBUO4ATJ5j6DFnSt62aZF2wrPYPml
TA7fgkUUkMmi1JtvSxYiz4NSnV0FhlIoqzhX0Ve26rzLmJfKa8qQG5jAh9CSLMPjevmsMwvwJDnd
3DKDlasYdbX1Eb9F1IMnS2/bE1EWTQiKFp2ZnkbVy2qi77NQs257OXjtG7jroMKUg4xjODilYdlX
rBJTCJQtEDuiD8gBojIQ17X5kMF3epr3SfY5YwnOXTDKWLpK2EZwNyFQS66akJ6mnlgPvst2N0+/
pa8f1mM+3bUE0zRD4zvqIJAiyEWxWUYw5hkgM06ZcvPeG3bwZFhue+VKtQgxT6XHB1PaqapZY2a3
QLi5O5jiG9n1sET2jY41xSoB0n3LuE8BZkJzqBNZ8nLscOmndp7vnUgC5kZsHPr3Xz2PENUhTnAr
VfslV7lBRTcaMhdoamjPMTH/4/lERmL7WFh4Kt8ZyeNA0Yyn/4T3MShSLDdxaXV9T3ux7nsHmJVx
RCMB19AoO4pRch/nZLmBOTBfL3KCLBBvdBgblvCt6AkDRz+6R11evP3HZqWKKT4ka6CFrGj63fIe
Ozfkt/yLLYPzperfHaUK5zLqMJMPo83ykzYort8X/Gs29Eq5CgyKzuofB7XZL8jIFX7KVwbpET6F
DqERg6e+PXsKaF00eCPvg2pnVHK3KWXH4bFtdtBYso87nTUKRztmR8qZ+vUOI6deHL4kzBeQR2TE
JwZmVY792D0kN/DyA+WjVz8/64AwP+bHcsSqt6dEwllGLC4QvvLxBGPs7LZOAKDYi/lu89pgnDL/
bKAtOXzc1oY052r8OnA0syU0D5/2DxWVf4tzGddgCrkgbEfrbXmsS9pnt6lndr0aSCuhAnwrFbtI
3YeoQ6GLdusdn4fJQ8JrPG9UcxNMNNAg76biwIrzSOQvJE3Vu+2uZsc7c2LEccJHSzHfzDO8VRHi
okqSqguQH8zgcByrrMLA0X/nO37pOhA3BXnLjaXChJhCEuJOAeV/MXnVpuRMizyfCkIdJ7zTWnTQ
70hBc5hPb/GGjp1Gnlo5H1iinp54i2zewjLpkpSzSqe2/I9B4XFqBg1jGB40r57fT+V1A7nQjIWk
ImGM2UA6Xprx+8e99UNIMDPcdwd7TJyFDWU6fBEXsqfFP5N7kSFed+NJcgMXypBxp7eBONTLVDTb
U5Igb6B4Tj1M+IYGzQEoy4Z8rPDFpYpWwyrSsouU/VhQZ0xIuVABqX3brLlKgdn7XXoKubGOKdtO
DNabnlJnGT4ZCxrXNXc6CUZQ8fH0FVlutz/Js8isVFsVNu+UiGoWNd9PFRWLJ3hNkbvKxz3lchrx
1X6jCicqAsgUff0f3oJFhSdhtTZTlFqrLr3fJpjj9ihu2RfiajLXnKS/mhnHdg9UwqLgRk0o9gbg
9ByGsFg3tM43KLRyQBevE9nPurw/b/R/LMpm+qBv5DfqHgp4N0T5LMo6pZnm1Av7XdpZ5XrPkdwX
HS3n6ph8w4SiJiU9VT2MtooQwX3nyLAsdCXPHyltxHjjZMmffBbbIoXMdt3GCRQUZ+HBodQefsPZ
dwbRTodRy/hkTQQ3k8jitGnTkF6H1qX9U5zmnMxTsvAmP/61mX+TJEqEKMjYovO8oZAs+4030Y49
aRTeYOeeslopfJLUZ/qppCv0aT42aNypdN7259NmNSWcGhGORr/pDm2l6YtWFkrEPd/luAWABfoo
52mGTv0ntPwTu6iGPnzUMYZ515Wy8hEsrcJwJnQo4JLxjf+/P/YLxbC3nM5MU9HxhQDBSjnUV8y4
BY3rCS3mxeWaNjXwldSyzTBk7sVPjWmK9CVGrms092AJ0j9kMK1jU4JMG7BUKoTNsFjwxvmsMZBQ
MVuAxz+7Pyoz1k413mTVjg9cq5phdVek8sB80mgb7Y6TK/5TzfDmIShufFNPTnWtoz6VIrS+N8Ls
eOvlXGl8o7Gpe9i4z4owebpPqzbSPzAHICYGaYf0nDZwlF6he6JQLiljV6L5X/irUIdCAze4qUj1
ypY7Lcya/gRVgXwKz2XTfjhkTiIpT4UpMTs+3jTFL+zXoYHOEM0Gdg2FsWEWQPuVzCtapC+l8vA/
f8lwCTdsIB3TO+iN7slI1ML2yP5VpaIEfSasf/VfxwllVGlqvPid9clLSUBIw6zuPvwTGCCCyU90
jplsq7K00K74Qxc8OKZWDMFsZ89cvblEry8w148tV1/sQpaoZKD4kfLDhzKmgKdNU+ywcSgcavnq
FRQOH9dewUu4hMCngdLloq/RRt3UaeAVVBYIwe3rwqUJYRRfagywnzEBhuSSj92nT2fsnSet3Qux
QhHIbsPhx4se4KucwZ2MuwsHU5QAJR+Z9kiWFBz5qJEbX5q7C6Zxq2CE1vxKF8H3VlRGCA3V9d8Q
vy9bH8HxltI7dYqFqDQOPKclJul8LEZsjhnp19ClwKNLWoUUjO8s4Uyl99vapq1QKCR4izDn9OG6
+rgShZAxWmuI/EqPI/oQ60DfmtSFf99q47nOnEa62zcz1qEFrV+gCRX1uWMGnIbEaylat10l65fX
D4t/+A1MWaWxXmRrpqh1vOJh3C//2PRwG1SuZQ+2vdUBdPnZamW/mC/7RiVwbbuuOKtRsBkOPDvf
ctnT3XNrWDvyvc66avUsLH/XGPni7gG/NY868Q66e7R9LvkDU+eYn00JPabEW/qIupoPdx2mH2Ca
i7vVgAtvcg2MQsfHWw17MP1UbT6lkbMgT01GX/E/s4VsFhFuQ2pj+mahZ3sj3jOrLyhCkaaWr/WG
qLj0ivtb5T02z/aiYMRCh6CKNLqjUHVOPqiVGsuOqicQU1ku6/kFCHTnSfGF96p2iHnj5E9fWE80
oc3VVQrjwpJu3R8MVuTAvXEqqVZu4yvdn0bEr5gO74jh6ZWgb4DDH9lmvMqUkL3Eaurh7OewGg0x
ySsvt2zUFEuTRoDhM65ZROrVD3xREciRsG9g59V2M1JXZflZGBiuYl34szTD3uFPghnOq3Uanq4l
HNBx70hP4R2ShhIki16P+3UTlpNUG4bCsBL71pWmRSfEpXUDQk+jxQzX9pjol/gFJT1NphjH3+i6
DeHido0eN7cf5Y85c38E/wOfbUfDqa5JxeU/MLd7afbaE/CZS9Vm5MzIAEdrlKiIRDb4m3R6XiIS
p/lrwJ4IP8LagGLGL7xwoBld8T6aFYKQKYCfa3qDzdpIwdu1tJNKM9KHQZwz4squ14Ey5q+kfHtu
KGBjmp1+zfHN8ulErKv1HIdFbZNS/Pj5VMx3MzEIgZ9gZCIMuHNZ9dukeMmlmoq6UtOhPFArF4XR
InSw2mHWU9c1y7Umc04InzD8P6AZjPOlY2iXpVVRm359ZMtvedSdaLfFm/X/l4e1osRfzU/7R8un
W1dk0nLlV+bKgTUdUfuqnKRMZdRJenXNcMo1KJX0Vr4nTrcRMDkHInwlfxzFaDhW4pMmjJw/C1su
LJ7wcgUPeugxJTYTZi8wcgHAn/jb9GJp+Og0IObFZfbtYpmJLXel7sfmYxzT9oXoRkFNrTj0ngxe
pXGjwNhtIi4YkQlU5gNSkPCkZOIyfgwi9i2prTrUN7jqMRlNwz92qYr0qKD37Ey3zRKEs0p5VINs
J4DcEEksv9C6yK3SmjtY9u5FJhNUQkWAJFMENU+2Y8nVRD70k5aliQdVHc0OmL8QBd1iv1OdlLdU
V8gNWX4bhxBR5JO6fWQet664d9pFCPQdlk4l2KeSoYt3OvmdNPfeuELb+eDsRbVGrqh3JMCbQeez
wy4fbQ6KgEFmknoC4V52WTzUpTDqK3r1ZoRUx73HY8ky28QlXHMJO8xc3o9luutQgyiJE2Yesm3J
aO4wGXJl9EuZ5J+fT6Sgbrx1jJAbO++idCh0aO9uJI0SJbyHjBiW+k83EmhPlv7lqTAjYrArN2Cm
S+i5BVhTWDkIV8CafaaZLvOwxqYRxxoGm6pJb/qN0o//TtekFflBmpw8BU9KboQ8mleFkDSRB2Ud
tY5n8ZAhb8g4dkI5bbnHdhKCahBZJkodUsxs5JqKpHgH1tIaX2WLGOtQ03j7DqR2IhItzOFo7qpO
RJDF0CtJWjh+zsOh47td43QUocFY49QC9mjpsLwaFX5AS1vBKHv7u4/2Pp+a3O0AqyQxy7V+0nep
wFNfihCc74ML+6M/Sp0o7JQj8Ug8LAUbzwU/+rmnKtmxmPedDiUEOk9Wupddn23PqNjykM4d5X3H
dEzKMliwqM77txSsbh3iWMcUhgy1nn2dQFPaChMxNKdK7ZIbiqhQ+TQHWFODKeDuy4OF3aVzzxfX
Tb+rYH3GAmn9av3XhFk39/6HiKF3xUtHcmtyrdEgV4bNVSIKlshfH8yQOTEPJkD3tJZNvLnopDsq
+Q0kCNIIMSIEF5N/gDk8IziM47Q/FUgokFtS1AzTM0AQ7AkWuj+h3hXJxkIsn1mrrplQMW+t8enP
bl54zbv+hspcdkyDRyzx1zTyNr38MvAg5rWrHqP/ZU6obhz06bNgWgU0tcNjmgeGUx7F+rN7qqce
ZG5+oIrViEFrqAIHhdftTEeYesyeOhFX3pQ/NvwRvFleKi8SZYaB12s7VGn3JMfCRq3SEsE0TXYJ
oQ/aQ97XqoCErneQ0fDaiy2jAufbVJvUCTFSpeEAhKFRxjvL16Gf3gfCl8KY4mCELDvOxvSgwwre
La5/PMr0w2TSAPl2riNleTlKq3MSbFyNpAJTMHDrvmsJHLhqniZtDRlzI/JsNC9NI0miYAk/e51M
52lI87jJk3Q2TuRkYe5YEjOTbSwCWmdQpg0tekbFgNczdeLUbZ223EqgEVmhUCcTyHIu1yyKRju4
PsosMWdW/ESS/EbMyJJFmXN5Yl8e8uZCinqWnAe0nzEMx6xCYrdYInGNoeTHINUa2xbQwZtiXa6L
SjHmcv0Dph5lPaAWCXjAE8mEbCgjdzGFjwPEUaz6gzjkzsdLLM12vKrOjK+z6re87eBteTuIP/J5
Q/pxcaxMgFNoDFgUX9i5uaQErGMTtrXOZjKbhPUBzUeGiR08i/Ga4HeMeKpbjMETRhtj3xIFhxOV
58xMyOnw4zn1Inw3zt9C5GU2cfBQrQj9WzsV0fKulEpvc0Iwv3SuInrpItYKph8IS3iRihoaAhkU
PUh2RyQFesTuIvyAMJFHk8jUhH7RbeNw32ZtolXaSgO6VhobZCWfeEgSivMhOeCMQ8c4Yrzw9768
Z2g1Cu+s9KL4U9frjip9pod9MWjJIrbCN7DOJIFbtvp46xUMN3R2N0fID1VNHaS6ZjRIed+tl4jz
+XEChQZd+dWirL82rlpTr/DdWz54gMxVqsRUM6TdmVAwi4kZnB0ydhhD3Tu+SrAVkwbnrLVHUZwn
buwLUJJfdQR32yb8UI0tIcOCAgRRMZ6H8uKtVuDkaLH3RG32bTyALNfudvdZiQW6knc740Ehs37+
EncLnc5drOPtcgpiOJYHEqioSvTertH1Ohv/oK+WvBqDsVX3qi82lOQk+fg+cKIo+TFAbRUbeyy/
0asG9ogpzB+dhu7uhFDAJdz7R2mmkIcrYrnbmqZz+JF78db6Y8Y5kIQKaCbjWM8zvKUNkodOpVlx
H+/iV4b7LrAYh84UiBn2fzBExKxuiB47dbOe3Pz3MxaYFIotG1eZCsRys51UiWZF/4xS1eGv1Ww8
w5Pc76oO7eIYl/WQbIRUcXT26Y224oVp+V6ijePLE3VHzoFZZhnMB1avbQMvvZFLcbGZhWNJKC66
tkTgr3sVZzjPEMQIywPISTpkhgdft2WjujKuKFs/YiO48gzF6li+D28432a4a60OuqlZlnVOLfYN
B6t3X1swDvQwugItzw2V7R2z3Ob+sQTx8V0J4nRhPCQgiLIP9sniFsuH7K/czRR+BHbBU8K9jWii
GkguBA2wHB4PCVs/Gxs2wmlXcwaYK28AE86IfL2I0qHZNJvEcO3OPQv1mEmWckYYuqd8PJMDxzhg
YY9Lh2sX5eUk0vk431XzYjthgze0FSl7qbMwBn8/ETRptVLku1q5BNieR+nJncxbO7GKEmmEMfOg
CJSx1/NQJkLCbwDIo1MIg8TetfJMobT0eOD1nU81fMR3bvqmfyyxLRJS/DqTAT8Elh1xyNKtBGE7
r+I4ruBu3vc3O1kpn0oGIOY6nOxoXVHnjkeEtM4Up25dmo2Srn19ePqfuxqx3VteHbJJ/RPKzUVl
MJadXenCQR+bRhFO7V1b9Kdksr7aQFjAaVCnq03GoDvhHSx/9TeJhP+wLIKGBdvmas1AwApHnFGy
VE883HYsPs6Ziq1WljzGJr41E6t8Dt/gFcTt8glfvYu/dbpcbo3pEt8yHCmHtvGl/Cli/EwtF/IY
iYNhMnyzSPDoKh5piXjqlcxK+1V4eDR8a+o23zPNs/b4fMGhXPjNKANheIS3ZEATT4QARYTDTyv1
bU2p4gm6Ej7hQPseLFKFY204Os/XaZqUJlM9h7OzR92nHRjeaSeJDUMtUblql5IlkPs4bwdk5sMx
g9+JMd5fZrGtmXXMPH81Es8G4Mda+gscRiJgTHspxviWwSJ907OS5rGfP9AxZp7bhNGNsF9pyU71
cfy+7VRf9ABuwRnvk0Bayto4TyQq3UKPaQVqz7Jn/ozF8qa+fIsF5ZcyP5lK5CaT35kIt0N63xpR
JHO3dlvQ4Cb4mpTZetNT2k2lv2mfVQQujW4YerVh67F7dhOSpRW7nXj7sh3ZMzwgtSWN68ZiqLV1
AdH7HbrZEVtc5RkpbWbvoTDrQ/5pYQNOS5JsVRD2LJ/H79U5gfHr3lIhdVJL29ADkGOMuHcGOEs9
u1X44H3FwyHpE1e9Lm2n69urjcSULQDoTa6WtjspysTHLXT7rsRRusWcztWF6k8vjllQfXjPvwM4
0Kv1wNQ4W8tkFKpQSxg1J1+NagTYF61ZhC7Qs5wKNmzGn2QlOXTMxQyCuxborZuoh7gPTeTqcQ/+
AE69l7CsbYZqQSOTS/QRPzef3ni7agwFoe3MSmkRkNn+plwFB/ZSa3O2qfyMgheH/7SfGpWz3Hlg
004vO03JK0WQnoZT1u8/zd8Qph8C4J/udImmWQ8jlegjWdMjNqFDbp208HmNo5VDpHSUkh6iClB8
yPGYYjixuywiBTFFFa7G+EtcN9WITL8gZ40aC8fxtvu7kF/2v5r9+HWJ9vv7UK4auxIi/I4pDBjM
+86CADTRcxouSbKUnsMiKtRTPH2ar3ETb7lVR1KoDqViaNpUREwFAPwAHUaorSfJRvEdrdbO8Jd5
tLbNmgzFonksb4eChakm5ojksQQXMDDr/2snNfDliNkwKuf/a0UN6KQ2GN5dRA2VqIqPkv3q0Kh1
BdoOpJNJkgHQqBb2zIvU+BpKXyN8nxXhiC2nOUCsk5nG6fjMNbTIX7dBjakAK5F03pFsh61v4Wyl
S+1YTTpYMYghmPX5qtRgi0rVShB3h2IXjz/XIz+Kkv51OziB9pMKEo+HomnP+0BmSdZwawpRKLGw
qMzHzRdrVg2SxozNIZNvrAIjpjcIQ2Ft8yNjRkqRNiUdQP1txiG/U6Vht0dBrlKL5ana26qab5Wj
8dBn0p6Z/pg49HwYIpgzTCRb2gdKoHzeyw2IqeaBY2V76vq1s9knZS3rrpEcrQ49IDEdlnY1Guuo
6aQM9RltbKdv31muqWqcSxdN1yxLe4n/DXQJguUk3BdL1Mg0TcboKoQBJ1oyZi+9OlrWrD+6i/LI
4hIc0Cc99o+Md/NHRCmi1bMFV/KjU0foDCyZ9EK4zBwhtSi+C11foii8v9+tkuK5BqKVQ8hf8/K0
L7wDLlpsVQlOGrmsuUPe1UMkV16W3fPuMA9S6HCbAfIh9jaTfKfNuc2C2L2eu+VmEJ4AaVBzZuJw
amdGwlxSECdyXps192qSX4ZJUT5qJzh4/X6u/cMRTBItLlApyyr8swhktnQC37yzbjEDTvZ3XmAs
c56MxWmLhNpFm+X1j0+OW5YMgDp4oMuPhXxvGTlk/UXkOZJRVujTKYhkhHA2IGPteKcWGom9VMOL
YN3gHQJOF3h10aKhhSvRPpOvx2eal01S/Wvb+l71U16KNS4xgM+mR4EmAsn/zkPQeJD5Xo4y6FHd
w7fHBQz6CNyMJMFGvmPBuYLbjVJtbRW0iJpNYqOSOdPuXDLqSAl1uiOXTLsVpKCPiZ0y1ne+J6/S
I9px6CYG79I9BB7pSk5dt/piOzq7cvX1k6Erflc1/m2p9Q7T1LIYPeS9dM+v53APVPGUdXKUfA2x
ReBf5e5u+Smdz+rwW4LhtMq4VUrQuaGCkOMsztxgs6MZjc0wua2k22Sol1NpyrVWzFu/D1hIwrzO
3HyF4uRzU4xT0hqPffeWVmpo5x3lJWK5qn4npB/hkl4qFHVtIKf9U/qtw0Txg3xYH8xPS0v5TwTM
cDQyy65YQWe7cskzwDyoS0E9jni9g1EEvrOv23Hkma9sb7CWD+o3eCiYFhiDPC9b1KMAADEE9j7E
auz6iT74A/kZ7qUBV+k1ig0tKxvwe4hoqY+bG3VXc5FicCulQ200v9CMDjvKv+LSqqBCmu8Dpa64
XAnL90/9xVz45DKUyAbzv/Tnrgj6nfBpxuz9eT/1uRZdql4ZYo9BHUtxSQyvT8Evhc/TzGmf4/mz
dljkpj4UcuDT/Mg+Dn2SvolPMTMStetO2Qglp4c24IYeKFZPbiJtYhmHcZvyPZdAB2hNkZ5IGkB4
jUqza898wKJRU3+XPqwyXvfDYchPveaOfN68PhykR3SnVRNuOiEq/0y3eacfnwUR8GAb7GERiNfD
xJIQGHBPC5fEJEKxpyRFwOUzy0/LKdCeIDADgaQdMpYygTEakxQesfH1mBf6+ulAVtIQ8jwyc6Lq
VfYTXsFZ59nPm1NGShTPkfwiDexf5ywA8BWyi5RSY8seNMu1pecTjFk5bd+9QU4U7eMExACVMsuT
1SBjijXO8lEoF+KOSwO1bcHwom2xMSgAYKooNeTqxH+TIOxT0JTiTpC46DYlHcHh1m+PbegnAvaZ
qgOR5X4obwqFyq/ERgNDmZ6k4QNbabKUm3iEoJBoBQC6VjXG/GPl7+DnmGpIytsjiZVdIORgw7wS
d/tqMD2A1m/EvZotr/kgr0UKCf+3tr785LVajiEbK4Of1ID/VoEj39Wjfj5p3MDISYBIFZTMLthK
05O/o+JFpV1bvjPQBPuZYfCBXwi50hAgx0295O1hxDFccVLl3MbsUCTO91t0itR4K3o5OdrWLt7j
GdWm/ZlHOF4sZ6nMJHtVx6NmF7wKngytyrIjNgs7IMO6mFvgSlcJg/sD/RKWAP06VgWN0vlZUuLg
7WzC/03/OV2DNEqSAX6cnofR308vqo67lpWMhinQ8i5V7nEVl63JYMzk3nCD4iQ4fxCKKrz78jeA
FU9d0v43DxSsW0aXo3Qk2JD/yYfO5g3uqQeKTBpCVzS/PQlbleW33BJMoSv+l6/O0w73zllkcTsK
vDdkkjA9kBSfE5aADBXDtsTn67NyW13j2CHBjdhemLHxYzKtoL+MLv6ws7xM6Ba2A/fh9gLZGCI1
TQEUqu7wom08bnpAkb3I+jS9Mmz7KGgEfEc+KB3HdHP6XGs99DzdQuAFhFMK3UvmjEzFduH4kePa
g0kZcUZNTb7thkMj330bASNAlYypCo7IIWx1yPy/UKnzKp+lczJlrKrNZN/LovNSQqkVl+tuZiGc
B0XywwTb0YIocao86jwL24rVafPgCLSzttbClYL1vHfQDBfOlaELcCtcDJmUp7LAF0FLgZROcFFk
8kFuUoFQeLqD9hwStyPVxailpR0i//G8D8A7RDsYoYBL4TtYtAx/0Jvu07SLhPc4TEuRJeIXrk3W
4AUAucu9JYDEd75dbjd1lyxskD5h7d2ErrWLNknpDJimf3YrgI/8zsHg12zhUD7b3wPpMsfeGbgO
Id59X8ZOvqfDkFwqET96MPzQgrQMJuvu/5wJoFp9xPeG4raP/lwNt6a5o6+oagjVcCtx6e7BKBRX
vrM228nutfO0HNzig4+SPbYLgBe0OgAH1k7k9KeAZScdhwNj7rtRv7PWC0mkWSH3C7cVhiHTpEWs
CjyuAbSOaPqUVewEg1FLer60X/Dqhx9jwQivHijcnBKVVL4XQiuQ05H0BOLW3L9T55vPfNUYEjuA
2D5O2M1mbntbWS1Vx62U2u7xKWpkBRDgv20RIMs7SdD1COJb58EMYZKXU6KaV8XRl7SP7UX5Sm2L
o6WvrpdW+a+mLmIDz5Tez0ndMGnXc/fvwALNXpwak6NHYEg5AdtStWoBRvX5GPzdYmpxqa92katG
RcvuYpGkSF2GkUjU14OmNAEzUkLzscaSsSR0jDzFltcchecQsnIzXaiHwaA3EJPNy5ftOENtE9g6
KB1LinVkQooJ5gMR+pQmH6rRYCyp1vWeobYelhMobGK3mFi30WkKsMvAUJO5smUaB0Qhu7KTZS3K
NjIkyyir3yPivLETGWNfXMAoTujtLbsGl/qKyR3fcsl4CRAP3Bk8smE3VU8ZNWjXpWoqcdhoGVGb
JI67LT6rH9edQmZmMURO9vPblrn3ciSp8icBiU8uwfjtj5iapa072nEnSCzkrJ0ZIbY9M8DYWnQc
NV2GOlrVlrJqlTtD6kUSvUTmOJnrUEK/FziAYCBq3m7s3oTzPjPTXZw51dZLJr0LFwiFgZEJWndo
AmTDVOfXL8kVMIuWdVYOvXMvrZ2E5nCmIkXeWla1GMUNtrYQUgjeMPVUmfj0IoYPS3Yl0X9qIt/k
uDHyJoQq0o17jZqxh3S4bE/zmFekPL91UNVtyfDFsAAKQrZoZL6H0D1G/nirumMFJhiNcXkNctzP
4gSGM1TBW/Y5K0N4sgGKqY//9LE9tNjJqzrSCi35bhUJB7U2wu6O5R1+6UWQWkaVnfAjCFF91rRo
clRWZ8/eHbDlzobvxPBg3LzsxmfKJYRzjr4i1CKnNI4zPUJ0azrWCkc1klpkDNwNASigmpGj/8zI
g+wN0OUa67mVmOPeMnPrvTL5mjSw3XjQ0KMXHzLMr1ovn5T3zkGB/wnVAjIUVzFDWWFVNV6fmVun
nu51ZJyIrL+XxNqDZ8qJXhy6jgWBrgKlsIpjcT8uz8VK2q9cmm0JFSLa4taN40sAzoTmHmkEtC8d
CFRBh/TIo3+rasfyPnfaalmCjZrKTFyCdD3h4r9DqiaL4uD/Y1/3R9iR6VRCiv77HeRDzDgWCONi
/fG9BMBz/kSM5LXr3KZkFja0ZGyQsQnTOODIwjKikOjW/hBIRVqgJAi8oQO+duekU9vhxaeCSr6W
Gqe3iB1hvTyYm1yFFMm5aWspUAAXqlj7hjagyMP32OKQEzYDvI1vmMWqJpjGU6s5C+1wVCY+4Luu
TpwBwviCb39irm3CUgEMLJ5KcoVOgqoWHgCH9JOHc1fnLWCZlNkCoMWOJ/ya2/9FLvP1Qeu7mP1N
QbToNH3PZJ8sa33AIJzetPFdHybiS9Xw7PJ40lHYKnxkVpu3tHBm64ZZFElUjwEELO4oI4actD4Y
PM+EWUfWbeZQldlvyEpequ74LXcHKehtGKNhoA5QC4VLRLcXwuVCWcTCVBoJfVYjE3sriUlIBZ1Z
tTaFGuAnX3yFkh7TRlugJJcUnW3xyuSW2Yfx4IMvKXH9zFz2OtFp8pJBaEgi1XLV1aK7+tE5enLD
vCgiypdyvfGH5k9aeUh7HDtETMhT13L2heVAttEhRARCj+UHtgtvYysJjr4zeq8YwW72knxwOk56
zLLhOZzshbv+akz6OElTRc4P45UeO05wv0iqEZYzZmS6cre3RWW8MoFi0NBefOMt4cI4hCdIuw6J
meCzCjWDy2cJuKlk67M6VidsTnDvaynCyHafRT6ag5yOD03gU8fBb0jcWgAOchEwwC9mlHZ6OI0u
6Q9kBBlAHq+P0vqE0s/d6S/EgB+cgyjCFm/VqUop5GOIsr/KEM30TQPdeqivnKHqVUeWTTdAwAXv
T8inAe3MnCRe5wbzCzlhvucGcrkVl0/WekEJ+/Swc+swJz5dC066Tf0Q8gdXNHkii78ZeEjfbwUr
rY8D4VcD1jD7JO6D7ZGi5EwjeeQl3svwZv2S6zDv9yrdlxvBpkc6GGhQiAROulbSg/vP8l6g2H72
w9pj/cwD1/NZK3lwEq2GH/Cf1QkcgmRZ+4VBrr/JwI9WicciNR/bdxH5fB7QGJK8wPYaZ0mZ78hm
C/WZ89ws4aavn932SuV93dI9aky268tWLZPp+M1rnkI2+r0nFG1rK4Mpd/iTCAAEQ+kBqqA/o10i
Z0k8R4wW3u3qqbHUc2WfJU63FF+9MpCCcaCQXcCz46PysQC9iDY9VGFx859yp902g39rbWBJRonH
ZTBDum+v1ThH3dsiSiMUCwF0tHZsZvN3eMfLtSbAH5AKARF6VKimv2KmTirgt8jFqC6ighORpVMB
03BSAdGHPATYrNX1EQuZSHgpPYvbfGv6HbStJhEHKaH5pPh34lccx1SpeVoX8VXJSwJpuLCEPWK0
tSZ5SAXgvRyt8r2tG5j8V+NbYGWnz3Qp1HObIoaMHTAaezdyUjYAGrVXXsmFbJfgOSJuuxH+lg7h
6YIGcHpIbZCspf+jGfMSfMnvOyGGMb3i3e/WirsAbM2hKK48LIcOwMKgQWEncgU7EOk3LM9B/fO2
A+CEf8vKsbHAKINpTFg6F7yZ1VUq/wa9KLqQO7u0BPTCuhnzEAEjbroDICNvFXSzCCKxNDes8/h8
SruhzyGw3ObCQzwJE0ELRFmWeO8PyJMRUE6AY81zHscVkZAkVyQE/vtaQxeGOANm7zOSShuH5JHA
2aBNuksl/ZuJ99TJj5SW84tpRwxRSNKtvTE/x6hiB5JSYSJwiFo7mFCZ3RPyLn/X3f4bLnIs/VQ0
n7a1Qc5ZMuLg4toRgssI4Y4Sb54RgxmgRrM7MGWrX1LJut1s3zDUqGgD9xMlG/fBZYMJkAxa8/Qs
K0u0s3ENzFdkEPIgJWuQU7Qnpux4qSHdX9BCUnu/XI/HiTcmD2caKEsqzU35QI11e95FrBaSSgUA
GkabAe0++nYL4eE8p+PDQ+4/YuN4vXkYgtZQvyqSoLPeXqtnRcpY0Te174U5zCtfnIB0sadoyh74
9oJBviqCrautY0zhjRXj0PSA5LrBlkvFOPpiyhv7PloTfS/5XFNjruUJyoJ0SYMwNViB2QiF76nj
IXP9NNvrQzPMwa0gvw7HfSx9/fgDckBQ79al+SlsVdzrzUsioXaY4rtNhBLGNIyg4aYcGTqR8Inm
RbIA/oMif5CNZ8fATNXqiWNgbJLbShs3FYh1jlqdwMUg0zEEPAgb5FDI054MyXTsWLLKyFH5IWp9
6HCVYIA4et5IjH0FYirVlN69gEzN+SSQ+jVnzdB6S5YPUeq8CHRhpuhpT90xNE4YnQshRMIVKSNL
O0OOk9e4LdBnP0SMIw12bMAfoRhj1gQtfMSK2i2Yc14Lrg1YRMcnLMIU6JHiPZssO6r47LzPuGHi
hbR7EtBUvKiqeCxiqMywCNb8KOw0+rzoDYsDKp6u7AGNg0VG4sDkNSAHL0zi4Dr+jiDx9eVsFtky
+MCUnw5o+b0pGAcFbSR4tMJ3keH9WI6BKMO3PxI1uTm2DgS+nUqmB269/WRNoFo64BsiJ/3SwRRy
aFUVuMdgoBiP5ItpJQIoMZ0xXO01Cflr1+jkoXHOWx66dmNTD8hl86LknRktpS/Cun2gxmTVJTbP
G0ZZz3l5WO0bxoTxrEqZOfUegYPF3dXEmC4mLOeBuDP904Ha46X+lFPbHCLNKMflUd5VZU8eXSBm
AwfXPe7jH/VTDCwKTOsTHVLNKbzomYorCiqZ1D7NLS8byEyD5ec5DItwurp6S19QSCGEmBwq3WrD
2IOX1Bkxx9578cLa1YH+O2D6CM8n9nWaYVuIV/6b6Tqo+i0rocuqkF1Vz5fSZK6VLKCFXe32xXih
dn5nzrmoHJlv+LlTL5HSHJhM5l5eIPWallyjzDahdoMMre767G3rj7IFxM9ICh3JIUDnCVreXLTP
hs613s/a/6klU8fDtt6ClgY8i5w1M/MKxgXftlvjgjLHyQkJW3sPL/XdE07v2O04zYny7Nk4HQNK
JPW4WJRDPObRkjXRWBEoFGakFkwe26tXBmS5NppKFUalnUu6QdHKqGeTbFl8ECl0+MneKpMboDVx
OuXp88qtTbDXmjR0qWXezIZuME5zpYs1VWarWOTa3gp7IksMgn3OJ6ArUilkG2MTAGy7Rcd1BPA6
eOwRukdWcpGS39+4L3aYaeHMTSGGaqlGmyzyUVqIZDPW7ZOisOv3hM4LtfP3KqA0WVxMu8QNfv3C
w9DoUi2aXMA2lk52HmC4y629+DvFk6AO7x7dUVGHFtVwks8uZB1j2P/byQ4MQHIj99Gp7vYr9LTN
cFsLAC8ZUISZ8SDcYc8EerhGKxqEZ74sE+8wPhTf7BBPJq1fQtdcV75j3YB2Xatk9tvaBkmvfwX9
MoTaEhsQEN+3lsMsqQCxEpCzuYX2JcqeGvdq5hFBMNqj434eetxniVudJ8G/U8fQVCU4D8/S6clD
B4TLzc7mnVvwSSriu4T7QCORoYMfHgJjeOlgCozsH2nihrMT7qNY/zXXOxYMvZC5utCg2HeQJgRW
h3gylg7O6VoIgCRGnBH/LwhpCrZZn+sbHOA9xK4m1VDq2sOnZxen09uoDgjZ1hN9C9ZTT4jOj6QX
cQ2ikMEItgj+EgBHuKWBlW2WkSuwui30fS7nVfqws22gto4dDg4TWunLeQRJCwTopFft963RN5I9
p2kMa98AYoerwb8NvQzY+/lQw25MYJjWco9hqQPgTUMoNw3Vbsrt3DoWeB+i5K6kNeibmbp/3T5E
7mu/H8fb6H0yruGJzoqxrcPu9Q3v2jbGx8M+73gHcer/jhevMr0s9E6Lxj0fas7FjSSvliUC3YgO
eHepUPdQt5ZVjvf49ZTP0YY8MYbQ3f1JZafbVwNAymqPaN+0eAQ0z2MSsEviAiJXQ/Ki1wgifz4D
sa89EgOjPnMqc4JoBuV9P3mnW58PQihPaDLQUJD47xnvMeinkAuu6kWZ+ZleVsb3Jm2a87y+Taco
sfOncpKdwiFDR/z7h7RzYUw/UZ2oyMf1xkYirOG8QEtkFffs8hG27HLtIkQiAhDGh/abxYONyEWa
Jnjjg8CXpdwSe6iQeXLVMnLdjWCHibfyHDmYtDYqAWGoBNkSGRnGHf81oCQNt5InMZhl0jog0eLG
vSRaGIJxxWBPByKgLm9+mnblYLqYi98FhaoZ7Z/OEPpI+Y8ctRGFKw1ByEkvr4gYh0slAwXjyA2x
brDZtbhODVcr/cSc77yLjGjyJ1TrjAr4yxf4sUTOG93p5MxlGS/IbBNC5VO1PClPBspnqwDkTUrp
aU5RosK5XSWvzwHqPUcHGXIIHfqvdvdbc1+s9OiMmPNGcEnxPxUWohZv29Rr9NIn3M9kWTO/0oZO
3zt7JU/whoDH+6fFRKRNfIDqYOkqCxaHI2OC5LQqNGpYV9u+d75Y7EZGqe/kX6BseWmdynzzDzxN
RG75ePduogCoB/dIDEMfxAXEJyAt6myfUdDZO2d/V3k28rEhaGrghoayxy3VDePylozIJysOALNk
g6TybGPvDxOeecAzs+jwlJQHlAiBGOXZ6ctsRPMkunUvUbSBWtp7i069SiHhOAFEPEXnl6uO6qUa
i03j3xOgw7zRuN3DZ+TLBh5fm36tyVZnte7tkirThimZUG13N21+Kh603N08wlo7d1kKg8duxqk9
R+do24UFvwjjayodfGTZf+r6kDBV0g8UrHxJm1E6OyRDcbnXzdcJACD2wpqPD3bMI6K2unReBY2D
Y4cImYb3eYy9SYpm1d4n0Ts2mjpwetWWc4PyyDlcfmCB+7k6ZAToAYGbhjbd3tZCfNS/xjdDBFPT
jlJF6jof3RDanwCQKnOPzrFXAjcZ4iuD7ISOC0Zkkn+5vC5hSZlVS1Gv/veBeXMpKPlDa2nwwQw6
D1hZaR3cduLQ0f3+yC1q23VSQ3/6cEzs780jwh7wYJrtfxW/t+QEK8U9rwl07aw5stMczBckR5/F
+HWZKDvRlm8IlTc3HtZ1dBcJMg2AG7aKV8i6O6OspckAFnm7vvbyhLb88PHPG2x20nlbbJiVc//b
iZV1NkllT7AoP63PtsDcIfmk/XGUk2vGkXuL9YwAENdNif9g1r1A0QDDFLmqaJ6BlKhYarwhvHtL
tnsnd/fSAkjNBdBWjVccX1I/9gXlWYWUJTYWmTwkfE9I5Eg8ZULvVMiTM6vV6SVqzATYeFrGyfIq
q3FwDI/AS6u9/Z8/PoC2nlfkg5D7hyX+7pjWpjecIm4f8i7W1kVLskzcB2gsymB1I76ojhwI58gk
EERRIJYfy8lIlDGDrIa+dvwIF73+iZsiuWvXkTtpoaSWCBcZNrwh/spAZ06rRIrh0FdIII5uSoWJ
WSKd63gFUzqSRJRWeofiw+mNsObIKBXMKfFW1148n8coPkpDYFqYqSnN+TtqHbr2fffrELW5B0wX
sf0endXhZKdB6Ii49d+uik2ivJv5ZRZIC9Lv/MStrp7147IH+LuDG+RqBABGZcHvvoxGziJeClLQ
D5U3v2N9aXUxdnkvGgdxi+sptVvK7Z0bxt/wg+bsZ0UD62dosnii8kJtfnjFshHUyh9e34slHvNa
Q64PTJJ6tVRyNCiksezNvp8WPhrrU3sC6hEjkS5hKIqGqat5o503w5j4XNCfP2EEthXP6JUhdLyf
mzhJVY8FxU1m9jvCuui5+yZRxvWofBE+lIi0WIU2Zl2rdl25xR0X0mITrrHn1d9gytO+aGfuxpE+
iL8UW/PpcxxN9Ynbl7AMwfNBNStXFKMYIBYFNPuzwbMZCHOZE39dAif3AEBEtt1URKmmSqGRA8z7
qolSRKDRv6vofiey185NdHncfBNMbM9QECgYE1sVOiWi6EeHs5AcWfdUhHgi4+zsxf+g/PvI8Z8h
TnJTin9sRZQbn6fvOfROHAf8BoemaYiwu3QFWL9S0TDhL+85Pwt8rD5WoT631SzVfHFUTF7kdXhd
sKxQekvrDa+kW10QAJTI0Qb+J8O8p3BP3Ia8UVP7Hh257z86o9aJHfqYXxWOOCaYZBc6JJSssv2f
GdbjK5uQTGkslFMeqi53qlrvrFO8jqIcp5oeLu97g0lm0M7ecxTZNwn0bm1rEoz42QeLNy90yuz2
bSUAi1hWe/pS70fmBFBf3UEAks7V48cBOnE10FFPXXEd0zWlg6YO2VXQG58Vp/4i3ggFb1hOVpX+
7nTJywqGytwRKvhjm/TtrEIwiSonhnwKrj6sVhjeobey8QZBMF43Mder/pjcC/lrdu06vHb8EIMA
bNq0ztzPHXMlapqIVSWagFLJy89qP/wsqUyjz6GR7HZX9iX8fcsbb0yN2NNCSRrvZ5Gka9klG9fc
14SqxyJoBoQJ50wou2NU7y+MzfR5/5qtTpavCydXnWzMd2qbGVzigP96MZcyjHt2qzRGKZcgtEn9
rknxArGmzBFPbE0OlmlCHvkCtTPIH157MAAHdRS3Ik5OGcqqS4CaiWFA/szTEWVsinCHD++hZc//
3QiiBKQP+w9oYHEsX7fzPS5h37xRwvJTKz06BWpLRjLbCfZeSwzIvqPND4WEOYLgP2brd+yVckBH
DWA+MwocgjSMMynK2Fa/XZ9pF2VYKeP9VSg0Sc4FU2mDOU3ROkt7SOGMyYKIuAj4dBL3u8irRs8X
DjqSKU+2UpXxg7wbzHdw6BlC0Wem5UP2+vOg3vuJ8s1RDTneqaH7b7CtYTrPwruMRjvBGepqzLcI
KzBsJbeapiYajiiCxXr5oUswHz7FpTO/F4rT5NVkS5KKdBpF4rzRLL6ebEjXC8jHYKtpsZQHYXza
SvwqDqliGoUQpf/URCkjB49TWLj+oLLsucP1POcmU6gDda/EvO+LR1HvbF7fuEDIWpJq7Ttglal1
o6l0yKrMvq8DY8EO/HFRDTRedT313VRoE0swR9iSVsOU7XhbYEGRCFaABpzXiG44d4JkLSoD1soa
AwuuseLwkMSXsBauGeK/PaVk1QAfRwtX9mr6s9Qw3PyNZrMpacq+D9qx4FwZ0d1sEIxXRFEUNcKi
mUY4p18jlBUx2KUjk2+WhkogoAyTC27tigfa+TlTnSK2mHsGMsiCvzqbTYjsoK9IzYY06mii2B8X
JxSGVk6iIJJ8TcqiIY/oSfpwTO9mlmfG1aO8szW6kdHrOwbhCinRyplcRr2RQxtWHDY0odIpvg3I
A6vhkmACokrOSqzWof9pMBKr+eOo0AZgq5HPTAVeihL0CAdypeCWE45HxUMQG54l+MzpjUMkyfqu
qTc6Rl4U5UqXiK3vRAXTpdF+IwfuyvYFoD215pDzIu3HtJBEyBW1kFj9pDZ11FpOHKZb8ob/3HcI
4tAvbUIB8s5awkjHjwEp+FdxW+ptov3R7pEQSIi/gkHYxEVkBUJ3enYsf1li3qASe1ss6UhYEYBo
UMa0STqpC7G+IMmoOSIhPWp3wapPPVlIiwF9XIpPDECybzThSZgRl0RhRTvn4ogLjewjcB+Z58zh
GGI1Net3cYaCXKx1VGG9C0BPBb6BbQev8ZfjrcKULX8c0SuYytuSD5l5VFCTZOFncBgQhhnLq8xR
pn9D1AEoQbMdcaeNXJtil5iUHOh9a291bxERl4QqWorjAutHNuFNNqXRMI+RZeYOizLxiJwCOzXB
FMJpH1zigYqcmZZ1DM9w4Kn1DMVQMIyW/hKLB2MKlTX4TY0nt5HzlLOEsREZRXfNUMX8LwtVyZgL
dzYr1Dv42N3Xx7r0k8uF5zWCtr7mmAihlEeLgRiZfl6hIgQZvAfMYe6A/aacM+GO+qnDVc/kumoi
Mj+9tXl5Z2p+AGL1qJgmDpT1mmu12WoXjUi9GZJQOSCeQAPphYaXRQtWvVzwPyyVQ7EprHQ9QsPg
vxzzitxSgFCiaE6m4Akht9I1nJTXEijD6wouBBtvAsnkLwYyOTVZS0FtfdtS/1jJ8YBjhw91kqRd
bAK6Tl7Bm97rHMWfrb4hLstZZhRTh7UBZRECm0HUmpiC3DYIl/QPNVoJUyJg5qC7cRzwwzN7sjCX
1So9QaiLdXBUTrhE243Yh5HNUe9FkWwhkgB7qpSHhSbz1MbkgbI2z+z2lPttAk0qXJ9D7ABiq5xN
YEH5XFSdJbnHF5tXeFbirxF8UiF3t5+tgiMyCD1YNCBGimTG+4L6FvA7FlhI4y8bvQtn4Lp6Es7+
Pi2o0UPhiHrbPE9/X/za5V65ZkTLiA0K/bpmx2LfryR6oJxCIu9g5lcz2saOZH3fL29F3SomrHIR
thB7mFjy7yZfuvTw4v9CePwApH9T11Nb+5xNdzDhdfDYkkofweyG7ZmSH2nLXIlLKyTSanu9jNlm
HKT0XULH2yOzFw94Q4jA7lmHcjCRoentQi/UuEFfB0Z24xWmc3m0ScctLbKm1rb4JMr7Huc+l24H
hzQzePKmIOqFuxgALKWhUx/dIFhwc8parLoSZoD8S6LMvB7o88H6bJ/9SyfapHS4fcLZv9WA31ur
MpSetZu49Y2pIMumBlYXYOSF+TL3RqKBiBcDuK8Oj4yjUuoRPR4kfE5xl+/5xVtRciu0ytj2eMwE
28HNi40vJH0JuUSWgnKJHmKOyzhgGXWxaO4d9ineXjobmLiTz2nT8v3UtC9OA59hC3s+1n0yFDpq
zGdPpT1irGoATXTj8tlKRtke3jQ4PfQY11NdEmTQOuZnCBk5dINnQdB9svBbytzEXzW7OYHVr+C+
wVc/WIDkdDqxx9OgGF/IG7FKaf37ke/OKDCv1kuw0N4YmDvxk2y/x2XMZCwffX2sgxaydUVuEtLw
TCesfcrmWECu9hqmcX53Aq+Xswrx89FLjNSzJ8l4wNXmUkjMkA7kZZ5a2311ti1NtiFGMs/Z2+Yh
zF4zQVoNRyq7ooWQ9jePkN6ZEbIdn9r0vAviRUIYE72I638hj2qzPoiYG+JAk2hc/xqDE8EPMUVH
IFCr2Ye6qn4wtf7hkDQ5L5/U6OWCkXuYidwOWbqg5WkvnQ+Cd3Bb9lhCrXbDCBRTwILUAtq2qnlH
heF69t1aLxjK7Xf6zFSWCmcYI4UktUEXE3Iz/Wn52V/PVYSmLYL1DNR6td8V3DesgG6+m23kc/ky
dHFchYrAR/TVHg9uJG8ZXw7lGzcrH6s3hM2ol7aZcl8YIl9pK0QlxWLGit9wj8F9ACwNSoZVDJtV
XGBIxgsJAAv+EsP04YIWQBhHVB1J+yjiSilonmZqPB+NZqVOqa2FHmBqN2rl8xzZlBup/ntRwg2j
IR2jAaa3Vx6NQKlUwHfxIV8AdOTXxLpuQiA+qOOdRcvzIKpb008USFTd/4BoDqseHXfM0XSbBhA+
z3qKstPq0LEKBSHLc0P9SKNGxW6sMtrUPkFJm57uyB5R3KHBafD1t6ltdtCE0aJE5sLxH/EdAVgy
NAaBQjeZdJ/OXhE3AKjGaxOHVK9FA64K9u07BoQYPG82h7A47u0hOtnekhgknAMm3z7y5AWJCb+i
+/cBekIOBADOSFn4UpM8KVzDGNUcxq+cr0Xql5d1mzvKVclPyvMZupHgWUGH5xEwoQP25F/3TdP3
foqpqyomiO2wJJLME8CCzgMiVXIfW0jdFAcblOGpsiHhVElA6CRupc1PZhOmRl8TYJPt6ko5Molm
WwljpdIZzuCOerU3YTyY5wqPgkXwxDtPWVVJkW9V1Xxel5kn9aQhpG2HgZS0rJQuD67AGw8JHo6h
4gIOTee4DaOTMoviJK532qZjAeFZ2jMHIYPGUKgVUd5oAcNSB5B1IY8rngEopXI1QHHMQMsl6WxR
w+34C9le035tBS752cD6T2H336EVcot9RK5e05u8r/4g4gR1LIiWVBworL+UC4oujlUMQfD3d15P
HFzaxGhVmsAQwq0iUlQlvIFo67VgjDeTUBuz+QVZ5T+ZFmHJmJFgJDcEdXbGxU6mHPQBd2feFpIA
4rryfhdd5cj4xCjj3JXcA6xGVJu2Hhd3c9a3yIb/wRjluxgjMKvXEFaNmeBEjHsGlgp4wI5xX5O2
bponyLotAUjEV7acRlAc3z3+6YF8LsCWkWNtkRE4BoFdoS2tp+jbO5c9BFYdFyzBLD/zRoaGsCWk
0f8Vwnd2O2bhnqWTdAJFTpgCARgY3MYUEhH2BY5V3XqbxeIa1KXGKI1/RtVOpm5BEGsZb5WitJ5F
9xsfkhrNXTDpa/6SkAH6QNGjweXEgsrhORm5EO1pinAuygWyXGJFolzAnPxNz/i3DlGfpN+BjzIu
10pej7YcjqMDUmIqbdKKadD0ITyh8dvtdyzU+D9UY+CAJt/17cG09hFB6dYjkFCDI7D+OImvLw9e
9FtkEgas1QdmUQuLhnHs6MV4r+KU1eOMQP47vmJCp/sOgJV42gIN9pGm4dWGB/kr67ITKupiDtcU
LUsQhRpvqqP8C/p+70H4YpTwSBS6e3qi049lAv8DJq/brxvkVZerWegGqxHhb6TwnWsaFZDp4DEK
eV1ZRr67Mc/mqCj/9vjd4YdmbauZ+SGtNWnD4RlJVDSFDBC+BYDebE3NtOXOjUiXFc7HaPig2r70
V39RQW5JLsWaFujO3D5mxnb2BvfhnmXHWgaeqfjKLT9wbertUsjs7unfX0e/mFcffBOl56GNEUnD
FjVYc5OJ+5pmBiJa+7oTHWYNlJ5cTkakuO9+rLG9iGBMhleWP2pZTBGuAHGAt1YnvHhrXYqyDLL/
nIHXniAjgP6f3adzGQnP12lbKQk8p/a8Ow3flnf9ASGYvpXHMMbTDJZgogKnbov+KJC697UQ4ud/
d1hplcCxgknB/v4TqzSplNXWAW5AqGPrCsfTRF44HGmfpS0KQEHKMy+D/3cNmAftwYDP2vWbeAfx
BjMQ/uhDZzY6Q2/a4ZibCmBm4E9U/0otrYr/6Br/ajw9R9BXxp4TqTXvSE0ZoBvQBfubiCg2WjCN
G5TWu2MrZRQhMVmMEtkz9khKwYZ32gQZHRcc01jDhsEwvHE49yWW2iB0v8QEGnEnbJbQ33UMfjXc
ftASNJ4tKGtDv3axvi3gEPIjNYWyq63GFk2vnkjYJE4dBQbBexyZNc8S4eklZv2uKfBKQpToVW5l
rJ8AyBNjPMNHXO+yi+SKYGmZOsWbOHDNUPyRNx7PCNwipJApjBD2kBTAA+0YS0bLbv9F63/93kld
Hb6SrUqvPz5Ywy9ZDVcGnEUvYagh/EPYRKs9meIuvOXrp8kAyVMxEEL4TkqDbG6sTs9CJlCh7Hnb
s98La437Q+obGWvP2/wW1RSIILTK2LYJ4oQOMSEzUCYCKLEtghtMd1+6CrdljCH89ryf3lbaycVT
UkWJkVyWldOPP+XctSWBQR28bs/bHGySbbnhdWT4iKbRdmZ7xpKtX2L4spZVH8HUy03ec7nPUh2D
DmlSITNBEjIa3uaYDyrIaiZejm/Aj1DprGwl+B1/DtsRxu2LYVhEH6RRhyMOgAjZvKBqgC/kmhik
Eva47Ck+kRnr2SqwaJNQiDC5m3FGmsmTbwiOU3qbheoTnXREbMMDKh7Go4Boe3md93up7RIdcX9q
aJmDDFvM0Hz1V9da4LOetrOqE1V1WA+wGwmdFkXy19fx7LG4WHCoJirbv1+QXmvHGNvw8u/3Aw1r
nbmjR67M8QTqirDU3Um//JnLxkVfO117ZdXkyEPUlXHfyB1q0c2sLwLaHu8HMGImBa1oAF7laYjq
p9aSBUfyozE+sDWbCtOo7kCquYtvUDBPRTMN5MmV2VaS0e7vxJ/kQUj5g7EkYbmf4kch406KP4fM
eEW+hC0TdGdjLtLPwaULyP5LQA1f4fvqSxNdfszpKr2DTr2jG+QycG6HrITPMOFDF1+u7OCyJGfR
mhmv/MvETH3U9sqHig0EDzDrcEuhPL0OGxq2CrgVe/5bCcIYyd2vnVlmBccpqYrIJsaBa3NZh9hy
TunSQraZircOOumnu5jkolZH6uyamtidzD7NU/8DeDwUHQQbzGoYKG7aopoaOeo4k87LnNz2sIJQ
kAHY2kengANfH6elsYyO4qQSuvaWbuNgoblu6pkEzEEdVPdUhnKbTppFlbDS0ZbCE0No731crQ53
IsCntapAXJxnXMA1nug9QGHuPYoB4oDE5L5Ov3rMgsxmB2zyYQHWQyIAnks3gJK4gXadXTUBIscq
ceqNTurZOKtyaP3IXB450BaoGc9JEgvMXf9sIlnaF7t36Q78yVQnwN6wMaq6eFUYnA/ibfki6tKE
hYcoDndI+0gN1yeBA3S4cVa9yXiO2UF2kPKhIiy2oWOqjcMxrW83puTMg7cz1YAEouNH+BsFrdtE
KXUmlwRcQzUxvz5D0d7dzr8v0AFAs3LEeX+ZDFjaFNTeD8fXdJQPA9pnf6uBQuY0C0EwvsaD0NI4
W6E3pDIhzojopxKj02bdNdOQ5AUkJs6FOWkvZHC1Sc62/g7Bk8hHomB6m/8M+ORy2MlCgY+ojWYA
K4TJulh+q0aUuIW2eLAybGScVLBopj25B+8TpnB1fY6cHu/9W38BkFyJFVbtPHbSraeIypOlxXWM
IBpetpAnl9jd+GVWuZkFXB5lvkkWAmbR05hXaG8v5sSNlj6bpUBsc2iHsfTrxyPvaP4jcZ/RNlfU
2ee2fr4MDg1p7QSvoXA7C3anyFa2k98B3jEh0HAmVMyl1LaOGPOGQjNCJwWofvcPYc56d5cOggm4
z+OQZ6D7g49p9k8Nk777xQG/u9WOMyeXrdM2mbBWEHwRRd/gqIeg3odcYnz5Qd9wnXObqQSJ3FPr
53tInNVjiFncwND1f/zkRZxvr5KeYL2OBxDoL5GQiyWBclfWY0U1SQDjNo5aguUtgv6CxG3ItoVN
RiWBc2gTysRG2UCiX2+72Rt+pScE6krthsS4eZBO5ZB/Rg5xnEiZMuR8QwoIVn/YTtSd4OeJFNVu
0/3g+lhaOnHw7+C87NKCjPs/c+hgMHCTNN54PuvdvVwLzDVGMSrQFWyM1uzCdHExoaPe9hr+S/3r
0QQxjTIM+7ZLBuFgQybahBcU2M5CwbrSh8bFONqjK4kIhI4MCmUp+nCQaGBVK9c3k3NzPIN8orrZ
DgwrHsyTXYLH/d0bpy4+k0ri9OnhTgOhzvh+jfE6imBA0N/eu+MOhMX25UpgL1etkf3SJyRiuriT
bTC0IMcYe8XE6WlZChTLcib0ajfClpEiepveosmR9VvzZTwLatoTfmg56yBNavEUXmRE1tTMTYT6
zi/KEBbTzKPhheEBcqCdVhX2ow/69DoKy+sfjkgHx/62sgUvw0aO4jWbjvFzaBq40VTFD3GhVM6C
EDtYetDVEf+H3KfW4XR1053fwNWpYa00mz+4CKlPexskRcNduPi2Vd3bJDzKjE1h5f96F/I+l34h
pqqal+3/I1HdvP3SsvsqSQqSPrJqtyX8DGLd00sykAJLEHd4lgVn9UZ+sq86h2B3JT2ZnRiap3fv
wOJg4/c+apGc7NnWW1cMTu+reC5+MlwNXqUCCtOqAZ3D+AcA94Tn4EYS8iiqywY7nCEHOKV0txU/
J2AkR0QrmZiYrQqeCdSJ74GpUHVfh8hL2gMVnEnLVl54UZX2hrhuD3oLaw5+VnrJ9eCP8WQdzKqV
zGOpDFhQ50LOGDG53/L43bI2rk/1/KauKpyoHDXUo2ppwC9EjUQ97iFzjSolwcD2Q6vo57WdmCw5
BBvT65IgXY6dtfKTFy+bCWOtZ2YV7F55ji7ihvKBm9EYeJpj9JnvA2fmym7UcgVohJ/Z64afPJ/J
X8ByuorzJ2EPfXy1yXB7FeQ/XJ1MXYd5lPbWnjUP5n3rZwIgbcCLLb693cwoJZWGq1IXRLkU0PeI
gJve+BDCsFEBYcPMbzK5ubYSDqJIR9P8tmNJQF/BI3gIugkb4HMXQNZYj05q5D3Yw2iyYHHesy5l
ofqaxqMtIT3oavhaaMEGOlTwUtSWwVZ/u+tkB8V4+IldbOPig6eM2WZvgSx4OK2mXwhzXcFmPjP9
xRK3XOdJOCP9VhOT0wbbRkLcrom2nR+iPiAX4F9Xr/hF5+xkqLlb98QzoXIkNEGIlN40OA2fQ7Xm
rSDfzJ1gL4WRajKh5LB4E3f2IiijyUxk52ptfwYUWO5v8KOZmDGd0no6n8EsZ1pyM9YHMM6MZQ/R
O+NdkVoikmzWg/p+pzJKRQj4UMymqFQFl7aRWF0qugkX0snTtwNe5Ksur+GLReJtfYah2NF10gWk
pKHVd09dsKq8348yzRmxLExODVnIe87wxWrGvw+QdUr2hgdnF2JjsjT9P3RyRgj1NDZZuBpRjdtf
i2t9HXsLEQAtzKPLgqws4uTj0TnzOEgF17p0jM5JxeZk8MUjKEarK/4GC4PorJk7HnsLYPLffpPJ
mZN45dXxaS/IZWdgCyYyY2G75zkzua3MMQGfPQ2amuqGO60xAO1U0LApOAADyhVqmN8sWriCGHcM
YClBujvMIfx6tlNo2ALzKpjtyFwzsw02Uzrdif0uSHU9YLso8ishAMafPgEdmoKcWXVXrtLOqxqI
kYbNtT059JojLd768dwFFpTf2yLlwDHKgeZOtej3rdhmPeezwYndKhPwSHQiiHutKJNkQa5gS0gk
YKUhs6GhWvnzNkZR3rJmpBb5PxYdApg81Wh2kT+mOmpLF+UrEdnTu6x2kKE+Ju6jIM07/xoXccix
yNbtKWsW/4DzUbUOULVQHRPbEMgpQ58XnLMFkUlgZDsUf0jZ2irWKf/uyrbk/3YyLPApVG+VYcGV
yD1YwEqSpCeYc9gYKjyds9wWjsm1k1rNSWdKCKI4y+20BCC7UK3VfAbdXHL/IJUWxnTXOwasG6dm
ykpCw7Xs3eVYmKrLJNeHCcDnSabaZ+PeQR9gqytxD5YSGs2cMQi+AHyjJAUb63Gsys0U8TOLprPC
4qG/FTKMFowaILVQ0UIi8olt1rIRj97jZ5ockPPpSov9yRFi1DCXizPSpO+fQAyYTSDoxVnrCKR6
KsA0nMI+n0Uf1gI9/7SlDKs/v0k6pxgA54v1ZmvRWG0ehS475Ttwr/X2QoQDkYhwIp7689lKrOCo
lYpqPm+QFldJPQTnFWOKq/GH+qJBqwCotYufBWPqN93G3NDrw5x/8ZzOu291NefhptwumpuzAQil
H/lEWqwQ9Rr18AFF0bkBTiodyoBypHZISM+4eIlOMeCP3T17tgEH2H9GnfQahBvgKLBNmgVdGwPB
nGGVtC6jYs+vYFua3U+5pC/L1df4eACkm1HqhngSjnvNGgPjKYOmCQNH4blwA+jOv+gkF0q7uiiu
Rns6sMbz/oJJVtmtM2UPxFwWbFXxM41/kB+sDk7/MGyrzBAarzxnST/vh59ZypMuuHTIgb39cokj
XcnqdN4RQuYCffaun+dUVzSbk1BDl7n+S8PP9ujewwSJCFikRkroDlRsIuiv3lwfVs4+lbN16z51
iKW5J4FwK93Kp2wbpfwbqSfnvH15CvCnInbwss9miu2d8iWAtjpW3wHtD7IBXWyHN4BARO7ZBXfM
mndBfjAl3zdhiD9Ll2d0+YScQPeac1I87EzREtpUKE786fLp9F1ZiOjzXU2uziWFhr4hCKI3vjzr
22nX8kfoym2TC0yTk27+swN+Kg51MwFWg2aA+UQUbdOC2qUzdT5ijYe8oMh3rd+DNEPpeFGGk83m
MmL0/Th+UAbktIGZMo4YEmNKkwUF0wmvOSEx7LZ10pG8/oeWXGNFrEOLqsRIuelP+uK+LBTII6Z0
6q+dtX4xDtGLDizMbFTjLZyL2IZZCbITnqpldGvKWT1gZ3yBWzg1zpgeSI/M9Um+H5x3cuf2iQEV
kNjA+eKPQe9J1VD4fYlU4GLtevYJrsisRN1b9XoO//kG3wrXVsaF9/UW6aQeSK+hdr/fyW3GN2/9
seq8rxWugCiv1Zyb9cx+jgnNgXl5TLgBkrg4YBeql+iTOI3bSd7BtnOGENN5/1v3dHU2rSwVHqlc
LfaV7exCTXCIaGyoI3j/fSEuljsvRWzGB4bADwln0MOMFdmAe5pGkIcBO19IpIoXoHUVi9gUH5jr
OszocQCNjnBNuNRm9xzhX/N1FtPaHSuK5k8MA3ifgk+AyU4vK2aZpDl4Xwf+DkpsASxOr6C491Eh
ZmkksX1nAuIhy3jYBdqxc0C5IySBLCaZc1YKck8WYofNMptW2FXmH2Lsb6S8tgu5zVjZKMWvAfhz
kmWrJfpeMc8COWDstsqEexGNzX711nDEEzIggqK6A8NELStqJD+q4WkxO8Ojv2eRlzRBsLd0tQ2g
mvElbLxrEIeZTKfdf3HzaQNgo3yUrVBUuJtq9Q1GCsHk6DDle72fRETPSNIfms1vApaEM+gI0MRZ
tcxJrI1EXMUumVYfJqz6UfEY4Sbse36BI1w7TiIK+sUievyUeud5dl00lukL3uIWKtB/OWvjI1JH
eHiXu1FyGSa0pA6rfV5QIpujAzmcISiTtmPmnLawsqo1PWP8mJ/UShyz/WDW7opPd6bSqViajaot
GED+KShcA67vGWbcxYoVMoe0vIsIfuJODfGgws8OdH1MbMOZ0GupsxnhHEFMgkrRE8K1bbD18lQM
T0TedKgxWj1NsVx5ST+njIMBVXhax5TgzCYZStpdQt3pBdV3koc/Hf49EwDVQuQ637rRL3R0txvi
QC1IiTDumGst0qJquoVM9Xk7lMeeA141bCCTGMcDIoTJktJ4AySE/DcUtfO18LcCz49ir1iQzYPs
n8Oy8boHfXz74L/2xSiyp/rL/3TT0buRfUzH+LJhdRmn5p0mDhYGjnvDjRH7ItlOrh0bzAIGBL7f
pUO/+1y1uFm8fKXIjDW5ZGC6qBocIgEH0QruGnp5ePUaa4QxCi5uRFZ0g1X46PqzhC1gAZx1k26U
dRiFqwJS4OIsJAzMF29efTWhNIrX6G55nFGdtZ6MxIP7Rh9GkurS3VuETAlfIEBwo9WWPM+RnSIn
rWsN2lqvKLLq/2CBv497oZ6mKtXoZy4/f/kAq6WGRNuk31lLNVh1bfCTH3ylZl8W4poq02vZk1LJ
nZ7wE5kYLbpQf8GMGb6rJ79cvPisBLDL6ytt9D1MTBnEFcHPDBe1TSDnsW8c/48UBEwpGOcnMFgI
zK7AcB3QBSgkoBkGDrW9HWVUTZ0nx49kKD683lZObltFg8ZsYjY8y+1Ziv9O/YOdqSF0lpKmBije
ND+/1f4y8hmj3fbgugZMHn+89/xmAMY/nfE8kATAE6eDRjg85+9obOeVspNT3FNJnw8rVwT7nqB2
sXlsaSiOoDkefZxwGoD16FcsdMIacox53oBnJeA5VWxs2qxAmXSS+v5pohtOvplpANhTcToqZ7N5
/msA8FXLHN7E13h8LNYtiF/31B7uRRz162Wnykq8I3vNcBB+PUvXYO8zDS5dRcAhydzXwsHHlx2X
vZhuvPO77gD6xpmhdb+xSJxnEVHMyt2v0nhtsJPyL7S7S1ARzv+nf4BaNW/y+8le/u8R4k4L0EwX
PyAQWsgUu6jaOXsFWGTodqryqNZ+ZbocGRacnYRWE5jo28Ye3KaNAYtcOkAlyjPTnb7r8qL2DVfH
I2F1lLbWdqwvypUlPl11ZUuAjoib3gy9xakYEsJF6RXS2nkrzFa0fQCITfSv05Zoyn5WaZTJgsUg
BNpJswb0Q57GLJQedDmwaY12xAAWEQHnSTqb7ahMBx/ediJj3YyLrmDDXpi1pjEHzK8vsSkGB9fg
H7oql/i7aqGb16YsyThNsGA4eiXPbGs+SSuwsxZCbC9k9oHntxe7nza5AdNk/GJn943Cxc591h5Z
vJji1XrgdDnjz6DFz4K/vui5ir25JAmNBhFX7V/cuwPvS0Ndl0E48HKZIX6ss0ZsJi1Eu1iRaJC+
u0tM5UFZzguuOkCjINLqma81Sn0jErmy2leOYMGN9jyEPzQ+55obW3jsyDIf6S/2eFAxP4R+39Hj
HnyH/CTeaLYFv8YphytmJ0UwkCZdKt7fobGGBdxRoBskToIdt8DwZPySEZOcNnRYvbjbRX1wvkCb
Pb4oOEIIq21J5DHCX9TfQPfPa4L3ct/dgMErGUovNZgF6A264od0xmzFqJonH7oV6g9gALNd5Vpy
mKn0iBeU/+AAM17kXNKd71hSMi9GvuIrM4zbZ8T9Ia6PMm6zhc7zwp5GMen1zdAvwtcNQiGUxO+l
vrOKfoTX4i3/Zs6F+ZUfQguFHQqSD9KmBnv10aWgUCqTRjq7edN88rXlviICaQC5b78P/gyuXUWC
Z+ANJQ+exrNwiUHE3VxrELWVQij6uTpMncvOB1dQ3bG6Ngc+BZs+woHV8H9D7sJ+spJ4NhMMxf9P
nk8Uxzd04FqZgoWg3eVvx+1szd1Kj98Gu6nAOK+TmKf4MOXVgMKqsslNRhnrYjgEJo09NeHeGu2q
Su4gyjxehj2ehL+kOP/T0HkyQPP+2vzm+S8x8SFYp481Z2GuBApJff/91rcaaU8fQ2vB9tCbwbVu
PkLyZXX8eiQBh1ckjfv0IS7aiFepFuxOYTWXHT8/WwXqrjfRHgFpIHcDYZ7OLW7dCr0vLVmiPgih
GKZnGf1EuKyFlGo7kw4K3ELZSaq2q8k1u+jo7iieLDmzS1ECB5blEXuxrCBzSvd91JXfP/LmLLdK
uFWrwKQINGWrjPQN4RMQuHbHxuAEnvMK3rlQlXXN1ekVNFcpasHkfVOLcI4sjKPw8IScDsri3CzA
YatVs2FLRzByFrT9MqqP/b86QsIPPBVKmsnliPD3UjkCQlwheUo4vS7hc9GfFnzzm+zi2CEVLSaw
uGec+qmDO7Nl65b8kAdqh3T/xawF/oH9IBgcaBuzKPjKmqmwhRfj6JbWopyNjRf0K6nnOiyX6jdX
Zm1jZ5Ig5hIu3iCrKH1uvO4t5Tafd9kkRvyZp9oUEQ6db80d2Y7i50HyYXG4G18cky6xBd2AIQl/
gOUxdhA8yzYz43+I3wBxjTtYcSlaby/X/QwcGMhlqHczD9BpAqmjCzX2Z0hTHlUEduhBsdaAfdg6
ToQVeIT/CsufN3VeNI21Ta2UM1r2zXToZIWRzPLvl/ukw9VO2f8EradCgj+cYoB6iRur9bEdg4P8
l3+di6IDBUuNavvJcdtIr+mpeh1K6xz+eYnECz6pDjIjElNTHRkapCH2mJdW1wqORc1SFmiJymXP
Gw/yJnXpodjwd1r7dsvuR5D7xkHPVX9YtNHgv95QzuqkK4WQk+QHd+1kovKeg1YBV3lpSbSY/pm0
mH3gEANOoUyfZHPqphhPo+GR65ZvZU3DZTTjBdG9W4z7Bv5lEJ046MVSfx9PysuEt5c9iUEJX0bV
l9BQn3AwWS6ZZNnOQLmNJvq7wGT/F/EFx8tpX6hrHoMVsGE3bwWW7TNFEhCfm+A7kGzy2SPZP7MG
LtJ54X6delQI7oEr469ZbO5J/WMx9C1Wi27eyFTFmZz9gJA2dYJ0Q4CmafLQAtJKWmD2n1NO+AQQ
FA7Tvy8xECXByFNxHUv/WrRhiePeIwTGchT74l1LNYYieRPzyFeLkYiPIl3v0FH7HbMHr861cdxV
7gmdxPcxvh9XiHyiv+weKb+soKphDVI2KUnQ5MIObAnMhFOcKaF2fXbzKhBi6zh78t1gnFEfUhTF
X2hKQXKg5BBP27XdhLihKq66u7u4WqOrijZU6oPc7QtOLvmxxVJ8aYwho/R4nGZadGgDyOEcgLUA
oYkxGlr5vBald3ESyVGOHo12HcUjXVqz9HtU0zPvPilRZ3PAnmz9PWLU6XCtEWYrt4QfNuyuLIUg
1ScYf1sxTpt6MiHcKn+X2/3OY8mg1sXVTPk5o1tleA+A4wbDzXzVEVOGajKYbDR/VRX23uq606V/
Ol39jIC07K1TCTtzjI9n2alIu+hnmjtAsm7aJh9zz4RgmLKRAmSKO4DEaesC1v5e4tHvYrv2lr0G
zU4fdgLBTV5PIaKa3iTsAI92VaH2HCqJCAwm/WsMWYqAJk9N/Gb8VwkUxbHrANQk0RK+Q3m1Qjc7
cVFeSmvlfxkIakW6bEFWvqj4j50/l/NPOaE+GGrhumN/N96Fo4Zacfasr/fpHj3poXfhlg7Z1hnf
Vvz4q3Tf9kkPqnsgJJrGChEghO5Qi9Ag8BCAnNVq025E64YYJ+PkIqOWstEbJ2lqDZJxgJTVwBkp
b+dRq1nZrZQ8Ny+Ddx0Uf/N7A98WFdFHD+Z78UMGhkkUTcBmCVCUpAO1D6H4CaNTxHpE6RA14V1q
YI8mjHSbFhYk2sbRNGcEw/rLOey5+VKoKHgtfrOdIFqqVC2YN6x5KuY1HMbkoTCd6Fb2RZWkO9sP
hMq1me9Auly+g2OOasNbfkKweDKRmffDpBAskcUOX9EAq5UimaJLJnyrJ7/gOE2S16fXpiahr0GU
OTRKkEzc7lDPRkqZGt5FZDclCVhZ8IlWaqfHAVe2kKiU+3c/fn5bOfjG7DJXHju5DbNhpTyl7E0H
Zpg6S3zy63DeDXRgZ5LxZUaabWjTB1Nn6ORjcU+/AWjOjrAtI+uGWNHMYe6V3U8JYbdaLLi8+vD0
kjKzQpLL+E6Ph+Ct8oS3sah1pxUP063xsQQoDgFmQC1WaAs8mrdrvnSxl3F/AaWAeFRsKdTLG/mv
RGrKTJbU6T3k/kv0cQmAMl0neQPnwjBsku33z7vBLzkKGMruW7rWC3a4dZeU3IUSEA+wL9+ci4de
+5Jl/iOB1KNC55+YN0vFSO+r3ZQfmVrqeTkDwJL6Yk7RjrWlzvbWXVWp+7egkjEC9vy7QXBs3Rad
uMdbGBssYN0M3etlFdcd1sF1dq7cIAPHt8eFMsJpSIuJePK5krObel26c9Avl0UdLh17N0tW23Bp
ABqnmxTMYnXLjiqG+2WYwxrMBO9NO4spNHzjiHVMfa+2Ot7UOU9hWfnYQRm0xWwbHAzdWRimkLZv
yb8VLVxeq9BClel3X9owgeSoWUBmAd7V0KqFBunrTKMKRMz5WwPz3pjLYluMd3Ah5vRgqCss/mxS
XooGh24eN0FxvIQT03skNQ+XEEY73SDiVPF7mqCUVsh0fnv0g2BlrqIMLliOBRWZSSv9ywQ8W71C
XP7RffnmuIWpEN9ui1Txgr1/P2UcZ9LsIBZK9iF+V7uXFNKLeI1VHMSKZldvhvikCiXMvIT8nOxB
4nxKmQfJhKsYIsH3wBje30yOtmLjFkhnK0BBV3kO3BtKy85BjCxvR+OUAdsebrPA09YNdQwvtqrL
tPpvMKkztTEGvZTohVcawz3SV9IRY3bwdf62y0/j+laxuI8dF8E3Xo4Voui5aXjCbXXo2HDZgmRm
xMfmAlwUepBAvr8IguPoQhR2Ipsg6u/e3cplIxdU8091inhdBHA+TswEdgGJq7+NwLppKuSluDxp
aGg13v/EiVIbwtujHqVBxIr99Ehfm17mZ7WtPmOGeXj3yHDTtpNRnWN9PkohMG2Y/JPzZJuZHqhP
zMqGo2XqKa32r890oGFYqrzNOMO3I7KAv9PWXXVNeRPJUCRtTvlx2w+Y3a4s49mEmLdjACCG6aVE
jfzonWN4ini8jOPz1/QV4Tw5h+gvclXOtUtFYClhDPYS8JeTTF8trYyKtiQUPISGF9Id6Ctx7Lqm
Tva9iGPiAYpBpT3l0Unjlo4ooceKrfJFndmLIBQKKzgh+usTB+3UTBexpgs9c6YHSUa8sQvS3wAp
BFMXOLeSbj1eIqmRjKcEeTuaUV+Vdq7kI5VyJPts8fE9xM/23Rr86f4cd/6lebZnzQYggLh6PKF1
RM9VhdmhvVS+3IZWBWWQhB08E7/6swi19RRmECJK4GYW9yQynnpyqZuGkpylQVIRfxcazd74XrzL
pfiXpQg1kB7s1fun4j+iCb5ay4TpVdiKwXaCLJ2eyEzqDCqT2ZB8wmqLqUeZcJVxEYUPsZCM6v4k
OvOuXtOsBf6sKzc2lF17leLAql3vSJV+xLeMUGAmpt2HftX6gAdNzgiX+urBqjZ38sPixu3k5HcE
5fxvXJVNwaZmSgULWaqQ1HviXcpr4SHcAKfCfCFKtoa8YRpqEzSvmxiIR+wgiB/Dyg5yLwq6oS0j
prnoyHm5T7XHvD38AZWRIvJAobO7vmMpH/QYRKQy6hznfr3ywKibGWUueOSD9qZTt+FzeN8rmV4+
xVf0ug/WTo+m6nTTA9AA6bogN7jKXmyYUdLhIF7YaD+Eg6HI1I03rRmFDCqJBIpb3cbPtGx2vk/0
WSs7VFp8U3qctVQLQk63E7oBMqOmn/8jSc0gkaxj9V7BGGwhAFu2HJgHnQ5L0d3Q7tnM4Xgj5Egg
xci16bb6JVnT+rMO7RTbWPvuR4BH9uEwweTH3o8xOxbrO1gdFyR43AB3bD/hPS6EDOMQ3zYlYe52
/nX0pkFywTzbJ0vHwco/1qf2PsDJkFIopXkJ36A+D10A0pg2aCj47o8lMh2nquMuRlh6mV3Aq3/J
iTpGQ3OE8wQjL//jGt1WQyaw9nK9JmJsxWbkxx/jn1EyWY+HbU9tPga0pLpx0EXmdtVQ7aHHGYY2
iFxJKluwj7BDZTBGcu4zkZa9hsKMG5elZtmdBxb9Ctfx9QN2LSzPlxwiBVNyU7ZSyGFQtTlOdr5y
87r575D14uXSEXaaKW8DiAykwA0m8Yyvm5DpgU5xp8L6lNUOtqYKD/phDMDsY4+zOM8CS7lfXk3w
RVN7kDfTYo9JkAojcqg3bnFhsuWRr4myMEoO5liO2uo+FMGW0aTFXiZScAg9dK4OQC/UEvZ2AO5m
uoSgoKJP/L4HNRQQKBfAboUojqGHe0nqwBTRyrTghcbLPkRkT577IQvQJj+E5MYxmMGtHaGrW/De
ByyS3x5reSjzkCTTwc1O8uuW9zGA7+/PR90j+LD4ATaHv2pOGJXdOBG7ItHxHAzKoWO5tSzHfpMd
horw/xiZS3WTKjbJrQ8SHXfXSewNuqbCpYRgkxUFSi5VebnsmOyppEyHgR7UTaUnw3luwAJ+X9YL
PGbpSI2Nm6i/6V4/AtmrTMxVolgy5WvUI1bmyjMAu+twAukAtKKVmkEnpqqCZhpodEWqKLDPKXhg
xlfFfUctVEVa1BQlHyiXXtTNyzeF1KhktMfZycB7mFsKfIrn9M+7atxubLDznZMHo6eNL3fFGzYG
Wf7mja1QnMYxPDL67Fw9fDfAcavi2xQdKY471m1ZooOlKDbbkkxhnE91vxKuIPrTRCk+R07T3Rc4
PPscASqb+7woFBD+G4BJnjv7r4QV1A+s6Exse8juxubdw3Mn8Ok4yaVPSxpG2AKdpxBv/keAG0LW
8qyKxnUkZ+VG3P/55z+sDaIyZ2E50XCicH/wWZAnc3epvgsHaQFgQLohb0Mnpj6/fHZseFCqcFUQ
gUppS2HdcbiMoPInC69ViuGnn2GCwP8XkOsjWc3uYky49OUfvuxEgnrwSjLo4LFsT/2NU87QUOXM
bVOjt5mmJ8zQ7wMoYGLuVnz9/dTCiN374tQPDXOUq00fu0CzAVEfxuaRu026peUddYifpgHn79AX
Kl9hSYpy1Ez4S4L/E9pmZM5UxU1F6JBexTrRBsz+9O0DzCZbYC0awoW5lCSIiIKZlKG5sumsPq4S
cklEbHx03spgmABaiDUjNdPy/3GWLjhYIDBXhuUiwRRh2iSss71sbL5F5ccX1cNJLDJMjh589Eh9
w2i2jTsnpn68nHr7qUF/WzuVetjAVhiNHzl4I14bl2K6+evhnhgfloI/40O04BwpSUHPpDvYdmua
fS0vE0N8TAMJ3nSVqIr9juY5CyWN5b2Cp+EKW8735Pt758vDi4xUDjhWTZOf8m6M6FCToSTFzy5P
hW+paVsaopDyyAS7rxrdNfVPgv2rbJeu/RM5avsqvNcxLQnx197xg4GNJk9hmt0PQu6WbNvNhT1O
XWcMdHSC2ao5+G/mm23AJ7pkLBNZf593SGdzyr1NrYDzf5cIgjxfFtyD2D9vk5hQwnmLB7cvpe9q
+4DJYeBpuj39OmXhlQu0Av67jlx5goZCVl28sCvL8EueXJC50dgzLg8bVSz3z98DJh934TqJZm78
kuYptM8qJGAVf+osc1TsGcBdNySXcUEFK6FFdoeaAxQ58w62ng8v5/rQyM5cECEM0ZfioYEF+dXp
u2NqvCly25F4nqNL6BXyEvhCgE3p1A3j7OHFuiCkEg473thb5F1TR8kq6BkwcnEUPjEbVaGrGowc
ZCqIVIsl0Rhaewctr47zlfd3/hBiumDe9jzlHoUOhHoOGqLmNew78hAe0ZKOtRKlFUeUNO64xuYv
gorEvkSYdGT1/bWitu/BmP1/CDAM5xBBPJMUmb/A/87LXNr3yrjA/bjPKK/zhsTzW/hpiGZEQyok
jmKmL9XmYhGOBPekEucK9RGeJyhVXU9w0TXubwLTPSWzRcuXOLge3fNB2l55bcYno4xq4TLKHXxQ
o0S4rYhGmvchxcWh/BAwLdh2KvJHQ4kYyxBunWTkVn9Idg9t83M/sehJcfwdYlkTejlKq91NFIbJ
2h06nttE4F3JgmiuQnsZFKD3MUEtFwQ6oXmR6onky+ne6aFnZt9ddRAGBnOiv09IBNSfM81dOGaS
D+Tc4U8EvFSLbZp0EU9dD7Hx3Rw5245NYH02DhJ088PPwIBNlGMn3MkqtDalYwerQJPCE1R1p+jc
u/2B5MXUv2IX3jhz5VGEnH1NXXFB07soJYsI6rqIYQr4umSo4t3cpyyQ49VW7ma/TpYwBNkS77bH
OV9tRB1YhenHeYk79eQ/8Ya9I108eEBOibzigED2eCUxRdwdoGsQReUqj6kM9krfJtKIxD5W2nT7
CDwI0kULxm4gAgXCB7FEVXxoNNiAQ2igRWh6jmZFd3O2cxm+07fFzZaua1JG4E0iUfXHQ5rqOKEP
5mAQPtf80mqLuatiGpfZbvNE6QFgYzrctaz5UPtxAUsswFr/i9iMw+zchaWwZvRgnMdmJZWZQsOb
SbKED65tEHrIARgotGp2dpCG/QHX+rIezkk4oMNgimwvenzPSAC2W0ceDAFGYAmFBJvHXqeyq+0x
wbO09an7SwceI5VMWecL3fn+tm2dkyrZFXWmRwHNOiPhrcSb6blpBkTn/jIkpX2XRvvy5cIlGFGP
VwNxpe8PGt2fna4UF1FGueqnIkVzjvL23OqAwwvDsVM/v2Y0vWkBHjrsRTTTba29Hi4ZaYlmlqHc
HvgBhCS4XOGE+c8ng11vHCvMVhuPEfvV/xFeQjZQFas//7HkFd76OMeeZRD1t4EzyXfeX1dmSqdc
AurXgPovq+07t8/aLaxjBn4XQaBL7sbbPGgZJFDLwpovOoFiEo7RMcnHsjUyT91Y1cQhG5z4uYHN
damQTAzgri1PLlQvRkGWphp1I9ZDFt9RjxfgjYVZvgGldopm8+NwEvz5k8RnlKTPjBy4vnRtujH8
+8o+iTEu1L5kQMKOYHdTASeA3WtPyLNKYC8GW5Uzf7/ADJOEJdMS79rpSOzrS78PkCKe+meD9r+u
pnaXB+ufgaFsOyLwIGg+kJgnhsq/KuWMlxM5TWpPFluImJguekK9SqCJ5mM/21Oh3wFJ1HMPTr0S
gPFqRXXxFQ9yE0bW7aDy5qyEN45BI+5ZTEz+0aZ5lQWxfTuAd4fJ2vU9l+NSEDpaW6FI9JW/hSuz
1Tr3ZVcXUernwe6grqWOKf2Pe4sfBjW8oI+Q0ZJ3hHM1BAyAY7C2iQPuHFO+Qv63yHh5ngadVsDR
+qmNmVZyXirpoW5UbuT68+tXMkzeSXh2l299XyHm9Z5cnDChSs9qj/P7U2YjMQGB8SUjS/YMPFkA
jezPbKPSzHAJ8untZvf5QTCtVSvESOwULVCzyzWScTSCo2JI9Xret2fuj79zVDQhLTL5IU92pYVS
ax7uBRGHGjPm2s0yQalO2L6V3vsz+kgQ475DOFWg7E4c5u7BDK6KJ3IRP9ymItYMGvW3kBqrAd8/
lpDH8wKqnEhxiczR3nQn8qbA2tgs/AoM9dgl1Dt+Oq33tSclk3jE4CN5ZpmwHl3scZF91GndxBiL
HJ5OqT1sRZvap7AV3HUNaoCtTT4EKry69J0HiwHQqVTd3RPohhmtD622CKwHyATsHr1YoFGj4eWB
ssfmIkGH+yLb1YQNMCD3bZdZWElxOpX3L34iAJIo0bPO0XL14hxVtmb3q6O8yXjXS0vCjKk9TwmW
NhevRTngwvjs/sVqbLZwNaJxSUsA/E1A7oHv025Xjn1nNzOZQS/kjjfL2reRcUJGUgePsyHUHUb0
84n1rPYAppZNUgMaQL5D+ymFITwKQtHjpvCUiSOhnPb3NZF/Mx8V58isJ9Tyrbkao4HxBJ8/1M4T
U0WyE3k2XmF6qAQwMEcaX8BH0KJwSCI7BZIR2bj9i+lvInnkHD6vN2vYLcQWpMV6c9HRQGURv/eP
IPYTLwBjfWu7oZhI/s6iwghzFxoWFcLwF71Fl04K2cA/1i7NGoSx3gqMDCQVJF6lFRFMoStuedP9
WroXOubEVicyLeDycEn9iv2NMtDsCCB22xgashx4Q7Mebx6RJTtIvUVbUOyKOh6n2XRcgZLprXSB
u5QoCVZFAiuGhZIAnMuuSHdankt2zJyfS1z6CFW5a47IdHtlJzUhfx29SLnl4opP7uYtyOyaZAnL
p2zjiMFiDToRkoUF35BGC9Zb/EjHk0N+X4nuPyHwdtP2a008MpSlK4CO9rqrpsj7ZmAfPUC1LQif
jAjv2yhMF4WcC5iSHLy3obIXBJm6WjOzGQ8trdxytzRrAqoJ6RSkqc+NV6Lyvze6oxwxB1be3jdT
kc/oHFTztzjDJqsdz1Jqf12obZtGPmEpqE7lCmrobA0I+5YBQTBWbtZz7wyb7gdfmvEUoGCdMB1+
NXkW58/MGyW5H8nzThFUpEq+pTKzhg2MAtBT7oSXinA0LGrpvfys5cwEPCykwsLMu1QYRZLrgeGf
rFtizankhMVvTm2dVbqskl+mXwWsHrdBlpwY92W2tKVPZFU1oygxanLFIe/tFR0qdnmdy0VETPli
uA/T7qNbepNgI5/PaHi80mQgk05F3CcEPn+cv6NEgJq3KbTS+ERhnpMcQ1nHQy9cEAaqO4bJMoA5
ZUxMi0Vvy7UEJpuoQlCcxrGZET95YgMdcdCe5pvJZ/dqYath7sl964jiuTCDCj3vrH3I7NgIVHSQ
7eKPaYmtPdcNlO4hFoRQPXNEezlaCWhv7k8vQMM3IayMN0W1oF7//7tL+MRgXZAto3ftCXFDywKx
lhwmDl5LWtPY+KBsYy1BGuBDUYNfPRsxu2Ciuvp1biE5xPR3uq9K3b2LL6nGd7EWQHiO3Sv81TLk
aQLc0Si+VoFw/bXn2vK+/TGYrjN8vRZ5YfsHxWM8cE/KdOib6CqXsbmDIQPnSCPbWmXlkLsZNFhh
hNFDKVNNQdXOMLMX3uGS8k4+qQARzRyKr5DCxw54JHd6s0lnLPZA5wYQSFykKYel2YDuEirMAdxU
fYH8doglD+DjFTebWtGYRo9jHlxONqRRCb7ghdbyczYNwj2+UPkWT55jeeozvI3LRPncJRZkxIwy
KWU9WAZETRc1LLekWI6GVAIw+Vc6dXFEDa+n0Tm6T+F18hdlY6y82Q8pjqBr2h+r1NxQDrBvKNj7
7IzTkbPDmS5GjTzGnT/fY+mzJ4yIMqtJXk2oxFv6cbcz3sdoKylFZFLn1CeJ2KtoYYAWUmCb2q5V
F3iwyXC2ppdNgmi6vXkdgPlPJlVJ8eGk4blvOo1YKpSOQXszXba1Te2wIcfs1H8lWca6B2LGul8c
t3sPrvjusfWYmCfGCPeMVXxB3w+1wcuNOZ+ioUHBXk77/chyUL3Xulg+C9qplnAWH9ThTrDPPjB1
ymLyDEj9AWp0xYBtuFGwb3EGpb6k9AVJgVZ0zjpHqn+8gW+qI64W5WLQQ7cTKbOV/C3U2ApZkq3o
S2fPNKUOmZrXGenOPuYJvoaqycQ6gq7MjsZhHP2K3T1SJiFKrFMJuCOv/s2OLZMIsWamcd51Qa7Z
9qo37/jvuhdVfBhONvkgx1GZ4pgjbktCGxSRfaBCvYoJYKnDLx0jcTeGXMKqgGo98pLz4EOxWIQN
VmO7IItOPAeWmMwRkfoGc48u3Jjo9FnI8z7OykYXlqSVbsbU1/NVzkjp2BLWgqQ/VwJGd0rW+ZEL
R91btGkKVAxsNDKSCO+nvLp1e6ZfH3UiEgtKtLpovGrCTG7KJvyE7DXizhs1ANvpm4/mprcJlFtF
fybiELD/CJZBlPQdLbwJ1rrP8B7P6VexKuTAwY7Lbe06IvIc+qy0KINSK5/DtXzqu1Zbuf6YLSWz
6NH6kEBCZHj8JuKxWYDmZO2WdJTeti07hx0DSILrpcIYY78M1sLNVsmfAFgnRLpZ14YK3v7A1W8u
zV0x50r+naC5ogGKcN0vdQIvzxxnm5m2L96eYnzbZn/NjFVMPgD998HtYFiiI+t21BwazIyJ9GdZ
o9SSY3FEKwroyJvF+XQZsWHpQgjnrG0ieXs3CVQHjmgdr/A9a2k3D9CwRWs3PcdRnwWGLXdW3uEB
nk1Znq8jtVmY00Byey50gSjqXms5eIc5PQZ2L6TdSUx9ysD5XC47vqvWXV9HIYyYZUVwWYGET0kf
qLpv4EH+2Gk95SIR5Fj69y0+XkVq6ObI0rr7oA3P43/96mgk4nTjCHFr1URKKJz1dYdXjmR4WY7Z
fhnjH7wN6MQa7dyVj8xm8BkxobOMRLELIshvD+tHf4LwZcw3N9P+ytywtsp0w26dnjwYqZtU7w5p
jCTM/ETWFvZ5bLSwd/QphZ7YzZ59OpDmlqho+qOQhJqElHuzcXQERT6TEi3IozIe1dDPhf3vwt6E
sm9DmFPTyAvT+p1hxBGuojSCHsOYjUofUPZonozU83LM6mrIF7CgM4b4bk2VR0WLKYf1hJuXzLdG
xnkxTy0xq+oMgtDg5NiTH6eKjVdmkn+2BpsKGNbkZ1vaPwTfs/v2wnm8eDo+glzkikQw2/P7GIMB
5awY4We8mbGJxybOP6TVW6fB3yB+pwBHaiPBZLZFX2vzR4taSHUNCehLOO4bdYH/oFwnjjYIOQWx
QQe1Q8OpvxqS6daHrwh68zF4AZEMJW5noCQ16I/jW1plxh0OtD8JxyiXAl5GJHt5v3ccVmlFii7k
TSdskuGFaBJabjwvAZBNRLE1uqs/UzlBluUvBCPeDGgeyHKCS7GnvEYvT49I3yH3EfFZF8jNnPvC
4gMranQkTO+Is4FjhSQlx7aHXNxHZiYpL2RaIk6+gUw1Zh9PbQ2Nn5SW4xb7xTYLluhW7cGKt6/Q
Ofu01zaqxU3J4mF79Z28CgKbkmxMuveHreNo9joJc1Y/ThQnQqVa6pwq65XPUakRxVoSNLryuxg/
4fvY8HCrTXwPggLnIZJcolqP6nCUvDBHJAm9W89Da6xqKm6KfNBkXXwdKjIOhmhdqpi/Bfeuekxp
9FGFDIC51FBmM8mIlgJ+0iI045Qaq4uYCM6ygV9dWrA99w9cA1UEw80Ju8ymj5zVFgmInlg8ijgr
Gb7XB94ggj/HUSe/npwoi+/fqwMcld0Jcp/TJBt3AgOVVLObI/ZXyBPSbt0GgnqCT4UxAXtIqUij
kE67g3CJl7myp/9fdadL6EbLew/W+ZSG1zlMpTi9nCM/PGC9fEvV7n+8+LaPlhDrA+Suj8lXekZF
6NCoLq934NhAlbCr6AWk3rtxLM96Kx6DrqfLmAVdguA2MQizqhNo2b9MIxVHv2O7GsqXftIxPA9C
jnjBEPsTLkXn8XAdEBcaArcGtixa97afJN3i8Rto3FauY7uOzvjWYfSfr3dbx7unZV5ZLY93XEnx
KvgKP0Txi/BmWk85JD4Bc12Fkmnai7JavsHJNwBhVsxH68e7AF/wdC+376J/82VqvU4rLx90ig+/
xjZGhidOVoews0TH/fG14TUDYmcl3zPKipdJL1WHQPV9tFEMSNarTtzCNUdnv42dNYqySmjBZDD/
Oyk2VfG7fH4/k2dOiK826gB88pcHG/tRI+r88OWsEKKqZ8kF/cA8+r6o0VwXdwi2lSML8iwqtdQa
TbYKczHqrtcBsoIpF8AMifIsPTPHiRXpbEN4O7KbEsN5UjTVrk2LjlJSuu4BWvA/CJAxvLm5w785
z5vZ/f80KIA250LENi1+igUWLHQLYpie6VYKD50R7RC4gzapeLFtC1NtrhrLA92zt19Ih0ZEqnqj
VW56T7HPhNlA95PFHtanWl224kGDopK50sSteOGQdsU8vdEDR7H1TovxYnJCb+fcYoj+/gpdDSsO
xuVCwz87FlM61d3fheCxUwnVwgRae7ISsfSMQOEDlrrcdPzJE5a05e2aDqXsiLoWgDDKbjYfVlXq
g0j6nbuaRbN6zsSc7mHXJBHv7NLVp6x3j36LgM5ei83vQ5uTyS++WBPh56tjE3ACoQJsU7tmavph
t3LIUmgCJ2RZ/kVM7R6Q5A42WjB7/O4jlFt5tz2pfIeefnE+2qhRUP7wi5hxo4AnZVXTod/qFQKU
4VHcCuM6EVk351T9vQPoGEoOUXER0n8MaeX03wlzQ4TN1/N/FX2ZnoGot0keAvHyiTizs8cHDxuc
8l7g0DT/DE1HQmRE0Qpu8/t3mW98/ZrUhVn/VjCNUe+wO4yc3v8KYrNVY+v9Otq9OwQvN9hswC7l
rtd3eZYxzLJD7NGi+n8FHnmblEv0opcXuka6Gu7ZAJ9pzwQXuSXFDa2j1OOfVUHqYkjCJR3nriuY
K5y4eDXd1b8CXgcxgQN6FYaWbAZw6unvxuzwijUfip12VciEagbPrZWdWam4nzEuZB+Gw4S6OQMS
lVIs9/4Fj56MA7isv+tu6yTc2RUDNmktvhB7caTyt714qhBORy0DH283xvVdY3XU0VYi0X04QvAq
ibJIfN0ahMJrrC1kxIMixyFMr7Lagq4QL4wEt1x5hQTUwMwKEOSNTSzaDgMveaSOgxU+Mn4E0uks
QpbrrWpv3kdfZGvI19EjxdtBf1NB9ETyjKxqWBvdVzLOsanW4YhVBzhcY0pGPMQwtMEBTY81CHxX
5KTBHspNkemwnyjbsFGQVBEvu04P98yMwgxHC9BAsEP8Fmq1twU0tsd5GgNOUen+KZzV7nEH7Q92
5DUefvvxvA+zWB/4Pds/7MstvW8bb/U4x9kSXCwos1gQF7Ov+m2e8H0hEaTlQUiJ67xFHlrX24NZ
HissRJ51Hm/g301zUiIqS8KCNTwxiMIzuY7ayY7Dvr09qntcyXgZunWwRxF5aK6JqjTeEaTlUHVQ
7t8+G3+1bX/6hotbYgthkZX+98/sBZVrIOU4efzpj2p5egrBvd/XE2mjQLtW1cZePSRAat2YPZXv
KiYDChQdCp6FZ103mJs4KyeKKA4SyLdiBk6cAyxnyfL6D9L39edTxydcfOBqtIA5tkHgcj/QNDV8
aleUG/FMUEhMIgNa8bIrjgcZVjg3vOEtfcJPI69uB7fVor2ZDEKPp6rDPAUZU7hivhIPcRSh3AY3
Ko11tN3DiKOctVWnY5qYlBAYXXrowUGZGvB41h/RDnhdlZjHWXoGCi9uAFDS5/sDaYOYiiKB3qBD
VDR7QkacfQxqHudlZpV6uILXrxHMm+yKuBspw5tl3odH1nsljd8OQipDDNHrHEaurDHhWLReiR5T
4PcJdU0ZXY5PIaRih5GaJScNgI6YNZVfoLr/iylE2nu03fSb9Rq0VP20vwofmktQlJxUQUyuUhwh
pt26S8R/mRttsoPyY1cCSROvVzFCB3ngGGuhUoT01UqZJ1nETQ+jYjF5pJcucs18QWILUOdcx3Tz
9xqlfUGj1ou/6zVw7iuA6IcwXliyzyOzb/oPVvFyjimH5kejWqiPLJViPaJYsXGk5ZFPdxv778i3
2HzfeYCkJHhaesIJ5uPvIxBkStD3MHLqjOgx2632f0dxsLK+SRFTffZYhwq8N766ZKJETdXFqiES
3+cSP/Rz7sNq+KTPPtQ/gDMokhiocBcpGLtlDEL/5YFCeV9fB7xVCxPatqj6txPHGH51FDURStE0
1KuxfRzQVKXJAF0/6NB2kUGSOZsbHLUVRfU1+eiWEJBvhLu0M7iythnM2MYGvCfJynxjrADuvM/f
YS9chK/nX6UkaDzsjB08NybnDy5NfyJLZ2CVs5R9wYEh96yaPAAJq8hit59AisgxpyTxCXc5RQtU
YvGYip607D3VXKTdzFc0+xTkHlrdp+r+Trt79SgaxWGMRn3Nnr2uM7OR5P1mfMIoj7DKX2fwNFKk
ypwXRW94g8oEAQWHwIxNmzwl+jVsvBsClhzQ0ECTWSYWF/fuiNGiiS+jbQRNzW5CWyqtcqWjy2a3
3VUjroWGbh2RGA71aAxeztoWpQv8f9caHzFOHRmbBEDZ5/MRytq6+VvxUBk6Dve+0Zl2J+gehBKl
Z7tNJc0FKA/391BPInPE+hOu1GgHtLef8uAXBu+ZTJAqdsiM6Mt/y5AmCcv+zpPkZBE6vUS/qAty
2g9I9dpJYIt/1fFK1aFkDqhf35ND8Z8+YInG8sEP3/y4heQDRcDhI+WgN+Oc4bAgugTjcyE7ssvc
tvozdbi7CCMjhzCgvUkyyYeJilEzvMj6++D1pJChTz+wauZemXBo8ibR8scz1qGu+9gkVoFGmJPy
DNgViYt582/s7cHdoSK2hJKHf13L+PkyGzsb1CwuvQWWw8QRs/gL6BT8JAvNvXxJ0RBPjK0EXmuY
Lo6ZgI1Np+diDuWEgH+HdMLvxn+mYlc1GGeN1glOvN2Iu0sUT2aYF8GsitrnJsHaIvvfMg6IveSL
2a38tbySS/NFF0Rk3Z3ptsaDLAto87/dAJGAfiRTu6o8GEwbqS9XKS0bPk/f8xf6YflC09jkyvuM
W37rXtW0bI0mRslRcAbJ4YX+ET3o5lNn18pxNQVU53sciIhotTxRdjWLWmZlOZVkvmZd/oLDONSe
UMohcZp21QncuO/1n7T98FXUXk906CtwcZjonBbZWJhc7rAn3TF+InCPMQBLWoE9L+bkEFlnIjWm
eqwbvjxPmfBurRGC+J/MEZjNcChxBNL4rymYpCh7SWY6OuhySGjGVZw+pFxWetxHJkCFhR40PQRs
0oP8hncvqzj2meYOSdhvDgToZP2LY0f/IxK9iHM6z1mnzcEXwA5bxP+BQaooqsnjjBv6QfVEJgKu
rZeV2mNygKdScmIo9wONvb5ixaoxSzram15ImoFCwxBwj1Q0DIEcsOyIfTeIc/RTgxt+RJeFjb4v
6mvl4emEe+lDtwLpNC0KJTkFGNgSiyzc+zIFGdoF5kfCF+duoKbCYXy2plvPh8JuLxhU3MV+3/Im
rbC/M4qAbeOhKL+ma5lcS2+B/aQ8CeSzwM/qhqV5AsJAbiTZyiwzBqbEAFdOMSjyZMNK9FJZvUG4
0Ou1vUyy+2g2WqctkAkSp3SVgvW0TGEwnM6MCvzfw7f2hvY5T+lAYf1C8V6aiwpLkHMn+T++MkOX
N7YSjkvGj8Nvf2WitPgm6b4OqcV8SFlu8Cn3iujAR7EfP7Oc9Kud8gtBKMksDeyCc1/21DQdrHCQ
enCGfU97qtWPqEtqDNLZa6icXbUsjtAhY9vRxYmCcs0DAKSQX7UnLpIFAcwtSLiR51+c+ziAfXC6
HXmjfIZBW1s9SauWMFDLjsin4PlI2ikvWG+UZaKoYrDGZFO+VKsMeJxfAU03eiMwJ4K3KFu40wyC
Df/NWmka5ta3W1FGW45LVRlVY1uL2cBaGeUbc5m72w7+bM7GA51uxgwDHCQ7HRKB9RpybbxmKt+3
ty47UfH/t4/2+a4OVX/NKcZfGnqz9cndGl7gx6dtbcYj7wVPZEvUAZLOuBRx251xoqMm6eI+L8Tb
/lsKLRtkrvM8sbioBiuBQWvYkg6Xj6cbRmdGHiWbBxiEZKFSCjKQa9hS2MpcKaRnYSObwaXb68/0
4y8cCQ90mrwmjU6ktDEhlVv+hcaOGAosWVnuaZWYMb53wC+gAHLdJmDh9+qjK4HmQZgQTMjgAjcR
JglvUgHKdEgajokqJhjOGecx+tFJ9VynUXMm8nVgdXD2XXU94QIBx4+NkyziQEFzRfitokzvtYme
gfEq7BwebC8/h92k+Ss5mBSGIMsrhIcUZDYn1KsMwmIPVuWZZbLM4WQIeTOROv1sFdQDMvNXUmGY
h9yFAvX3ontLJuIEqQpwT1fMTPBo2VD/S73veG3S2hRrm/UKjhu27Y24IOxfF7QUBvAL22ZD8tix
5AyCbJ5gczUIKnmm4ls7u+BzsvPP2JAkPHhaRb8EzJ3/A56H23FeeEicl/cTqptCr3SCUa9QA9QQ
0lNxuScnPKJJqQpZvM6th7wuC9vkCKPSh2B0iHt0B3302Rc5c7kREV4/9eKLccJd6jyaBUQD0Vjg
p/foM1qL+T36GiVxXVn6MSPLMDrnF9auOiLi2cQbhvItLwFcMIvnRx/ujuITcptqcE0g70jToAvG
wfjiC3Vs2MQbxuql0+/TbM7d7fUEb4veROqMDEZO517dythBl6Zz77ym6q5D5OEJFPQY2bk9Zhcb
+3apYVlf7d+IeL2B6GsCZC/fdWyHcolZHrv6aik3nzKgtQxBYb2ViBtZTlsqx1ymgMjHWUzZicsH
+rewO38lWDkYDXRRBsTUegYMzJOhFKiRz76oZY1ouO9Tk1edCMx7cDQ9LvY5HW5OYEpvelAfNxi8
n6LKCk4dubhRo/b4FGKlLJwP3nAyCm4vvpAECXETNBa4brNkl2+cpG/2d2ORiDed2jpkzzSPXpKT
F3ozGyCfb5SO5h9AmkXHoUh1I48XF0nnDI3d9wGkjjaEJLg7Es3J96Vfk/wiTW6GlyMDXtJ+d1uc
tMT6ivSEeEXzLC56EHkM0BnbBYLFgQVdHgO2vNJ3awCW4XqU7qgUPJgLrj83HS5zBMJLXyeJvamF
oJ6WW+P8LE8R1mmkDnAtWrrc6yNj6TgQ0ULZ5yzbxQt9fmXetC6/BPwsoeeGHUxbp3/priByeYjY
O3uljfYDanifUfLr7A3tHQQuv1p6kyr6oh/K7JMFPw7wt9ugc3BMs4egvQglM2X4y0CitEg8Cqtu
PpJZ0zjP/Y+HdrNJivYbVK5QQzh1m3YMe38dBVAzsf4Rr0nJAd3Z905Lckp7S7gPsgwmtIWYU9gX
8482JAkS6DO2aUdMDqm7Qv5O8DXrxc/1xr4hwJ3weq3WiyCEnO9RzF6IGn2LkwPhIRsPt9lQYxGX
rVZBH8oruBjTfZbe7vCz7hN3VowWh182W6lgpWJ1/ChI5PgUkkPoSG4gWoXrrsSpiHvH2RKZR49j
sRsCRonXd2WUzt7duM1VttXJHP9TKonvmYCjXXpF2IAx0H80d5FvITF0cq9EfUSeAtNCSJ2rUFVL
97ySybVKKm/RJVj+txgALVmKMEEqCK9OcRxWGGCNzUz9EkUDMJ1yt+WI8+VQT327nncuMaLRAqcn
6ZagAM5uG4njxNRydTV5x1pWyGZ6sw1hT/46ZeCw17lhio9mCuojTwFnyJhCM4MEs+CDYvA76fs7
wLXP6pnYFMS35IG9pR3RgaVGqxCFwop6/IJRXbfJk57vUqH0tiO0V0XspUfcG2Hvt4EZbfVS5R+z
C+VlQdM0Ls8X77W9G5hR3gTV8SbTzK4ee1mO2GIhQ8hhyYKvi7OfktcTO9YXW1fXTl85yPz6EJSt
FtYK9UIsaE2IJKz5n8BvBGmRAKwW0DKmcqOjfHhp0lmdH0pwmNYKsClyVQvd71JEsB2L6dVwj9cf
tT0rwRKvCyzfdT0evTEDLBOtDJonBUJUvOf59D9exTGRyhgzefrM5zzpkYP6tgkEGFrouHb/evPk
uN1k/UhbJ3AxhGUVMPo1mgZaI4VBGwQIhQ4I1NepRoHp76fKG5tm7k4fdbtz4LFX8fBINhArhAXy
q3joPcXl3vt69AyAR6g/CokyZPxompkPi7WTVoP3/c3wU0vsyzmPLd8RN8yIzzdX6xtuipNEdmDn
S0VuUr+o4zH+5XCrRWb5Of6vYY02UuMkPhKKK2L58EhfHmVIAAspjEf9BaSbQiPd/79qvjPHMB/w
GXNZhJyZQliE8v73rYn+ATHd5zAYvNYfTfgI6iH6rYHreLWsF0VyAzz4L7W2t3j9/fV1OSkqBMES
q8q7x8jys9dqfn6XMAadz8R8yrLYVksnA3PboRfxJONoNL7ShCubbXItAG10PmVLPidJEHZnY/8q
P1E0pJZYNEaga3v3LF57Nk01+ta5FJACVuPAbaBEm2yAOvvOvwwZ4aCkqWdfrN+gi8Cp1m10buNy
ArBJlM/dtwK4uy2edhhgrINXLxG5Xg9uP2bbsjkLN5f8SsXZeevbpJ1xRhbODyQp3git/CK0g4Bq
dRzqW44J3Ucw3YqjMW+ZreeE2tS+Ajl98PD6CwWWBUxhFxeACTmUewwsb55Y8HMPtoynyYPe5aKq
nGQjgxHqOwKuT3hcrOPGS/QCw4FwoZqi/vYNrN2t4ouKOh1oz/VD1w3cAJJpw6xXC3TUgicDitI0
Wriq3FTu4FtxZTpUZD5N7Rb23XRJuP6eUhDnH2SHfeNmN4MmW2cGcvRFCQcrH3Zix4XDyqTw6smb
eBBZl5icJfIk2AMkyjWCsnCOPRkxzvuNWwvNoNn710eV1nyc1DVyuRLv+lX4aYQfmvBwTzv7/qq3
iS41QoElq+msuZYpLs0YL8KGLE2S4kMrNx0XfRz9OtPOPt2V2RmsJ6Hk8fcWXtvuI8T01Qe9dneW
UumwVn8K4SHZelpZvES4PNCT36c17MuQauj86riK8TafymdFRjOSLPJp18bKIvfmFZudJGg0rA0C
IEH+OpEuuyGHTUKa7p3Hiea5ibooZg4VRi46qbFFjjVUc57kKoJYbdSH1phOyWFNmYTeQAsSfE/G
+kqt+cx/LzOx16KF3NlvVDCTVZIRQpGtPdKhj559f13znt9tWeo2yxqZtBkCXIVCR+3R17Bj/BFt
PA1wh4FddjJtG4uwJI6iATHCM39kSWSbxpIgu834hVN3ZtS+LyZFJCiEzhy0yomtm0l41dbOJu/A
/YFx64VVVuKD4jQh1FQj9t5rFJUVqCwMu9AU2DAt0UycEHwL+bpPVQA00wjFrYdKmXYO1ci7VfpH
0V961gCHIpzEDF6Q9NQu9Qvuos3KwFW0zw7P1mYbwlmo43kBJIRnydOJK+jwr+8aS8yq+HYzgFCc
HSsw4tbKSXER0S8TVAIs4khqlxZeFQerbCG7DFpmnWLtSZzKeMCeNnUkbRyADxRA536LUFw4B4LJ
mIDdPbItbPjQGsjCm3TuEQZwnFH392zGmIGg4j4DwMzYJZJylvLKSEIG+PlDPcQtQ1CJZgBw4svk
zL1Y1XL8sZfYpkxlRrX2+kTKHZVnSNRcsUhpmeuMWxZGcUzgACmHpGx2RkepMWTfhk84cchyyRmg
M6kx0dE9V41Hxy5gPa0vNEBjap2nk/B9WaIL0q9slfG7zVqyKLr4DNeMJhjc9AGhE8LgwQLKtEIu
TfsnQ8DyvcL2qjB8+gx8VqpcMLhzbgoWJJ6AMBIwzId6ZAG8mKW0Epiy4rMyb0XV8HC82GhyMOuK
feEt+sILisUF7+z6FkXeoZ5AekY7GXLeP4EbSK0ezjnZDlXT8ngl1Cgz113p1kD539hbLQaOi0an
jdKLCi4/UI/DCYXxCt77WKvek26gxPunYvB+AQUoiHm14KAZdrRTxldvgpC3G4+u4plnDM0IZZD+
iDSlxbHr2q7Qm2cuV8sZtsE9CJRvL7VPgwEVeCzejFXR44jy86fniW9KPCerRrKkQilXCxMyRVYT
6We5IG/kpm6crduCXgF2YbcaehlnjEyy9eNyj1YIzMkU2qjsT5ChGLiAUByo1F1rO82KwoPs46OM
T7n2WXyyVKr5KHROpWRFE91V2ZCJf1SWlCodAEjXTfSMWw3/k7uMA3oa+xsTAjojHnbhOu774VXF
B0QCtpD8m+LrTjhLEBC0ko3dEvpY4+LF0mZ1utvlS01Qp52oq8sUeDFcECFObysjy6MQrGfHNOsP
mBgq4znUtCNnpBZiLT7gAKlLo3qg9iskSccKEPkJGK3+vSWfCEziMHcsMv5oQ4bpN7/U2yExjhZj
SB1fq2QhIfZwRByuhPtKXNhy7IJAIrSBiJuaDsTeSr4E69F9a+/kFGx/DysHuNTWaA7NdfbW9eCy
p+HmTgM1AmBrFageiGLK3EeiLBXrLKw2MrO25IzkXORpcnmnPr5Au2fmYJo2I3k7Pulr9F5XlBQn
jgcOAgDPs9gbR4ob9vLwBdBFwBk/wL7flb7AcdhXGuDpwKhzke993UwNfDqI6KCaJsd9uADZ/qwm
ZQI0uvqDAK0Wk73UbRInWXecqMsE+ktawoX8UIn0c6F+HEjKWwwLCl5jAJN7RpUfD2Y8pv5P+BY2
E/2FWuYSF8Zxa6cBoLV7Ps5WIFx+DiVc4Qv3Mh1HQIRHIG9RtWMUK/XcKhf0MsQcNqbgxu8SFqkI
Br3ESqmntddKawMbpoCHIh+T5qVkEd82ZM4rTRsHgsqH5/fAOjbBSympgphMKKq8ArlY4Ij6nqjG
4qXa8k5jvVbcyKmwnlgka+V0CgyNs8Y58PboCwYYvTKSR4WpVfmtU6DzP/L5dp8mNkIdxvvym6SD
eZoTO3hIkVSjQpynQsED56m57l8vFF1xKHZL1w/YbxP0GrumShCVEd4BTGX6HYvmMSY1ITZEpJMP
eFCoQ/b5n9IodoorddGMEUxgYgQbenhW5F+2avICV0tsw1oAPqScQO0lQe8MamtVzg3oFMTmCbMe
OxW+EqzR94Ujso+EqQ/R6jle6n6fmZsf6XZctko5hTeTv93aBwFiWubRknekB/dDGh1bmZJL2+Cf
8LVLiDjZ7LELPIvg7hBUXCB+wxnR5KZ5AUN/IoKvZ2zhTk4BEZms/ME+rnRMvl03PsPhP5IU2iGY
cLGVjSOQ5MGqD10t1FZSHNIi1WuJZm9yVeSL/L6WJEMEid6Nixigo1gdfQFOeWgw2XPTKWvL7nOI
9bCEzdE/VPpPWsqI2rsvYLn7Ikkpujl3NcNHQBLZWDJIx1QIhE2jAI5xaZeEE54RwYmcsVsGZWtW
aRf7zSRfuYHFQJrN4LCjjTmgPJRoBhj7K6FTkJhVHmk72r1clYxZJ+j6XR/9iKET3pILzJdqLesf
rQaqVK0QxMRgNL/bBty97h+H2U6zc56gGu2rdvwAS+1I7Jwnd2HhYcKKqC1KWVGqux8HXsDxK8C7
jGVf+JWxgbwixzq5sDVB9Wi5F9saWj3j11bEWM7a9e8DvHYl14sVw+eG50h/jqu0y5BfZlqGSMPR
pbqgjN4OU+tOVS1AiOm6rFpZIp6mo1KHrdUqni869RTcJRkTt1QbLKLtEVcY33N5dsq8zWMut/wi
GAXROxRaPj1Atj0FO9fCnJHIobraMSsd/qne2vifyP0iRRGJoq89XbsRS6IZc9hdFZ5BcPLDB8WU
em6AGJvi94k9m9YmNA+feIPYjda/YcnA+Y7GG60ggO9b4mv6mMw/TM6QNgdqSK1245JknfCyN8aa
QVCi6e1alqOUXzBXu53LK9tqrD5VMhb6NyIv1L/lY2po39Mq1QYZAmTOQgRy1KKyeJGCtzRbjkq+
uFIj3JAYciCFXNpkgYRrr7Lyc9XDXyUzhizTbcQEN9CMZLUvNeq1zUui9LU8NTH2oW7jqO2eMCP3
waRPb7TNoAfHof/EpjjTEXKcha4nQFFMB/6Urq7z8Wc1a1+6m+zg+2K+YSz2EoPLvcn6Fz9tVEgf
QH1KGGIlT0M5Gw9Nm7KummZkj81BWhhSFRWXDT5k22fx+zrgVOxHPc85BBKAINW3MFnhRLDteFlM
mMUEQZW4CctahRl7mC9YvRuJPY62BK8begqmhLtyUvBok/SHtvKZ4fW6dzd7HWO/s2OvKG+RQ3P5
SrRjpOiXlEqpv2Cm1ynvBG0GpEeXSJFvpZG/i+cIFmoeMDHjmQZ4gz9Eyr+emenhZWQprQW0DHVt
1hNPyP5nPMdTmt+8e4W+45v0trZBjHvVpRAQ5BY+S6A7wH18tDctWfREnpa7YKJO5hv7k4F4fX3e
Vu00wJcZJ6bqgKgdTZjcY+TR3O17Er43IZwvrJSoTLqlTjMgkXHYBcsYMWXOxpIbpVb65Mo1VnGR
oKwzqabqLsZ/3HcVbSE0YXNVIRKq+DLv3L1JDmAfc1Xbve8UlumAoLCDcA2EyxIj6f+hN7rXDMsz
LZEhkiOXiITI8xszpwjwYVL2jENIvg2Un/mfKCHxV/kDf7RqkUt+TdIwEdk3M/oZUKvjRwS2/f1H
wimu37FchGonD5fI4x5PIB2lLjrIivJhL84ATEzEyQQQ4rgfr05C/kfVdUNKBktv85YO8na92Vpp
aZ1S7BxpkLMTQVhTEUc5BffJP1GBQJnanLQTCfEFOUZlDiLY2WsPPM3Waanln6x997+UyFghl7b5
X8f/TuX7B1TdXPeKh/aC3UFp2M9/fvN01+kocAnU0kd4vo38+JVIz0bawlVkM8ZwODL/s1Q8wrqI
W6WBxbKQ9bFENW6jWpHwoM7o+LcH0bDKT72dg4Fjn0Wvwg57Xl5UiAzVsZWOAbrZ3OrBnlVknsmA
20NZX1ornY1p5eUPmpFKI6J+vfGTrns7dyZ+mjEfEmf4AnIRYcBdKkjoMhxwAcUKI0NR6h1pQN0n
T1Rmvf/PhBEZdckCLd0BU2y00poYZra+IZ+ZVL2yN45lJzAKIUdbxrzaZEkFejmjoPvUX/hua+JJ
CcP8l8pjCtnGoURjjGAuL+6tS0tCFHdKa+EjOeRYyg1D82vTe+pImJX2GIzUzXRBxe1kIXS3Ejtj
CotVznmdxTYGAKQcKEp7IM04EO5v9VKlyEqlyeBD5UxEBLOloq/ubNYd6ZA1hPQ1JWZF/cUW5ZaU
9thQuM/DwGIVBGpu7ymTTZgTz7vKUpFs3zTqsnodg2/an2UZzJBN7rcaybpU1YKzUvs0yC4hDLSV
8E6l/QBpQyELelj1RMmaVU45XVQmShQc6/5e4OkMiw0byzwX90meotaLeQ0H6EixqKtaoYTdy0b8
LP7iC/T8QGXDNbdv4adaTyjA6XYRzctslOkpPSjt8UeIFmTwS0X444EYo6qfXd2Fj67w+0pCr3BC
GjxJ/l6I1mQrIYta1dEPGiDiB4yNZsUJ9ff0OnEBamqqbG40u3ksLCvkknHIepqjlg4ngM/1xUz5
pngcvQ+azJllPO6fQL8mtJctL1wKtYC4SQK5Z6RGV0l395Qv7oNvA0WTHqrRoEo+R3/LUbNJ33P4
4BlBWPdfZRsRa7mf2mdf8CJHQ701v4wyUYKnZiW9YH7TdfUdhPjjwhmkio+qhvwDa+X7NUyT/v/+
QLendDB91pfy2LHqZ9uNm9f9Yl2m1GD+d+iDQaiRuP9ROmLnseuw4J0J4H9BQDYgKXll1yu57cWv
W7nj2YHID35L9iuEhEULBLN0KeIenW8GN7L8xd7OU6ULEqL48zPFrIeHR1nplSLS72JOGO9CYPyu
/ikggT5CTOp22R1yp7869YVG2a1x3oMeoG/HMREJR0MtPlCtqAjd2cC7BrNzR1gmk6a7H2uh3rRl
Oii6olaeEtYRe4fBaTdUi9wBFARM4rV7thOS4FrgC7T1ndD+vLq5ef5BVFwtDftxqWpspFqLyCgI
EbXc6LL5NjlCP0j6jFDNCrxsb5uMUqp/75J7NxGxGQOhPukhXdsuB6Lr0eg5/zwWgSRi297rykmN
RhX2G1JvUPLNb9jwTPJ1fZFFF299YjVdtvny0j4G5zf5zRreU2GBl1mPthkMyqtuSgbiBYc5za23
DWOgVQnvDTWdpW1TUxdBp6RNHRr+XmqDX5vBL1E/pVfgEeYH72NWwYaRlVpRJff1WfMQuT4+StUH
/rGwyphoU1NBK+5y1xPtHRkHarGmaK3XawahWt4GN7Y3C6/XVMl4j67kXoTw+y7Ngq3ANK8jTMNg
STPbNbsbTPNvxlZJBi1hA2M0tNyzp6B8Lh9nxzsQgwSpDStW48ZPtIQxGA3j/GRGtzfjaXDT38hz
YUvWxmW2kdqTUXSOw6WImfefOml+0qyqFsG2tyhkhaQjfYMnqflifxLp8ksk4/utLS6z7LMyKQiJ
bWbzowzRBGhoXwe91NZAmLa3i4hGLm1WP96Ond7KinCRDTXfUdcaEloBXWGTM8m0ph9JRGqY+s2p
U2i7U8juL2973EPJrXmru+9H9t29p6Ja4dipkNiJqBapGJvYfi+W1VQrNyOA3lwqkUqbANxsKhC+
tXGLEgB7wlEmkxZYha+1yg/te09O/907kuOkqOlan2a/e3urGeoa40hnxflJIZZFPRxZRpBdcsU0
jSD9Ggg/a9+78frQpUmvxZ5NhLx0T1+jjF5iTVobM2sTX9Zo1TGow4nc3+uByYZi9pkfAgBotlOA
tPp9D5/W2NrCAlHODag+5cY7lW6NkR3vptqPcW/e2fUFFrlZZAPQvw8WTuSWnjF+af5ER9r6Et6D
o9klbUHWF3oBy2YSQ7Sw9Z+erlytA/VEtYmYymuc+EfhZG2DtQLJMaSh+gdzj8BpYdd0YhcrfJrB
9I7VB9HNqBhLssjvvHLIxv0Xy+V9aBdoO54/esiR2a76vROlNII9U2CDM4+qKpgq6Hkk4/z/aMNI
i23RURxlVYA0I9LBe8aZZlDbXivffdj/fZ6+o7MR5e5/uthgT3YcXDy6S3z4TNiW+D3PnQxVkJK3
+N/5YeEhoWtjwmw7H9/0OAY43bKIcPzbeWfPlVZgyE7wzu5PXZib+FHXkQNkMVGre1yMy/4QnY3n
eOJtXFm4/rvXP707VuT3iD213yarF/2hWvnXvTKYRu+2g+5yhQypEt4w0FvlGNuJptd3lyADCcST
LFZLLWgr9aDLcOzcVH46Iabpwe6l3EGmkZ4WVI6bGOvrDmG72xeZqpWqAvy8uzuTSyW9rPm84Jhu
TDIKt5PKXE4equcHXFCumOj2vZjuBVsB+tNbiYV3/VwZG0BDjmqM1u6e3hJgTjFWI3DMwP11c+AQ
bD7zzHdDPRIB9tL2AxepHaF8xEIbqwOEnK0+UVbpvd9s8jcpW206TKm7eJA1pidid/78EGoXAnCB
4599Q7C2AKcbn6WYkJznsLXVww66NC0utrbfvt0O0Z2IkhtgIzE5JjZT5JxidjEoqMagbXUcAvdy
K6QjGQNKKXGJbiZiGbMTeDM39pdw0eSfZDfnI1hZoDWB2soSn2PTX933PSu67lJZu0egpJQ07mJ6
fypPcaBJSoh1ld/fsU4rvbTCBLIza3r806LrMTuL1SIIa+q/yKuJ+R9e+z+yG4SV9ekE74kXnD3E
WPnyX8U7SssiDACa7idoKBykogjnc7Ca44jTJiJbps4KowTXxxyC3iDk5pGLpJ3P67Tvar61xUU1
ooit8SNm9SFi7zX5+6Xj5KP8NiyINbu5/OferiPf28yR6nAI+dPwg9n/MrY9CqGL+POTN02fFAVh
qtKivLbCDr8Rph2YmZARxUz4CMYNStRIEOwvnoT5Rr//QVwoReyEVwmDB4Uu1n9hoAMWvnQ33isv
2MORwRL4tbNVJbIXsIG0tnG282ahmDtBkeDExbZzaK+9OZzyz3BS3SkkwjnYS8N0WPqMHZlRn+WS
/X93/zqvD0yaOSU7RLZk9dSXoaam3h4c1R1IWEU5nCZSq573IUiwqwEB+cigB60lNsRHYOvxZ0Mz
33Tx54JVDOIVRKh/Zwh2rE0T7LH+P8ny17BOoAMLi0la0p5RNlws3ErENn9qM7M3l+O6SyajZLnZ
jELxyZs9SYM3IzX3A2qqVjWlNRRA0oz6iPWfIhQBKX0u+da3+bl9XEGTCiu75X3pyHlV9hjVx2sS
CqnQWFaZDc2eFCkyxJuTTpbEzsydp3QwuFBndCpEBPwFk5oMOskUbDIai4jBOPernD/DxHGQaj9o
FPtkF4/v2Q47QTazTrhM8VqiBiAQAgQVd7wbQ98RMS0KlnX18oSoyO6reEbO61fviPjCFHvMsCcK
Om/cY2i46Eo8bE783f8QILc7bGW3R3H8G2He782cmqHHA3HQXekEWPC8fY8P7g+4Fj/yTg6UiXCh
X7oqLtrh1fRw1ikLehDEmG7/KABEkS7iWB1v7GNfkkV3OEwY3KxlJRlPWddDs8vnDYbHMpc2Eyf5
R+kLcQjylSpyZofVjdCNP6pAEjlzXGDakrXwYAWsat34uzjwv6LluAL0z1bYwv3wJOq9wUIs7Fsh
ol3X7LBn82sWAZbQ1QYa6pf6cC/J1gNgJwFp8PIqnv6qjnUTK4lag/wZubg6bEiqi/Xu8JOaW2ZC
upqN5/KOoySwpcSHiotp3zfq6WqcRi+TeJ4/E42nBCzEizjyVDRR4LuZiG4RaCLvjWIae4MGkaWL
FWFxg+vMNvckOnlYPVRRwAca2uX7z515wjBgBCypFDLhdE8lisGejszPabZB/Ue4MIJkdV2ceyUU
Xo4PZMwf9JNYO6MMjBQZXRyeBtTAQ8O8ANa8JKzAAgJH6XUbH5Jh2pz+Badvfy+gUFV01utYh8t+
QcUhI+XT9MiCWysAMxIf6fKO9E/DRsbkq7lXK7/OYrpDRYrGQFxRcyWEuTSLXyaRW0pcQhRt5ij1
YIkLmzYaWE7JPFHofxl3yxYHdVGxqT9hiuGcXpNF+tQv7fvCIzawt+60pJ2nvVB4UejoZMaiHQ7m
uWncFzOnqdo2BIS7Z7VGRrjcz5nJ7UnLg5zeBEOUslPNPyWG81yORjiYbVmxhfvUywfImGhTqDVg
bQryj4sHGFzHdcGOZ0FE31qygZDwU41oVJ2v5Kh5NuyRP0rfzF+ZVbr2eS21H/X9F20f9e3kgDnN
avuJYqWnBwxJ2vbkiGsmOvd3N9KPLovBqFJwMJBWmcBBOgWyfYMjDpaSbmT7L1bmHnRkE/R63Z0t
00DzqPsUtL66VnpNfY+fzImOf9Y1i2k/45rNgehaBc6pB2Qs63eyiC/UZlDprAscJ6ViI1O/uhCX
4oaRy9X4qTz5THPEzEH6hLfKFPnFYOcakwbfGYW4lF5gCKW+tDOwBK8BhIMJPaGdWIQpyTSQFM1c
YscfNGvMnumsanZx79hxaEcHr0S0Y1Gol3EJQFMZEsaXoU8As5ioyhdPb9YGxDLC/CzpowO6rzNM
nVynqI0sMN0tGJbJhlA63gYnF/xXtWg+wSpftgteXdf1nbej8u4iGSH1yEyaN9o2Q8PeSoeN/hRT
5Zdf76ueCQYuoeEMMeX96CNYvyPilHjv6TZHmOJTyfKSN4p9xtwlzNPymqNOAHwN1GyneAa1rFdg
T3mQcDPXCmqfKrZcxlzJLTcb32ueBxhQIOVoEzwLkRdlottN8ieoApPONtYjPROdnxan9ChPzTry
G7F08oExeAihQVT/zRjvK9mYqhVT+fLT5s/0iUnDwOkbbtro2vUaAS2JU0f8Tis3gOJntYYs2JWO
o+ZCJXDqoKshYrSzCyBoeTn4CjbDzHF41ULTTi3h0QPfuJCdDJKLU4ov7v0caaleTCth1u96x4ik
YWpZc9dZ7ea+56zn+GPz+ZRpnU4bScsz8PRs34oKsi7NICapL0nZdUDZx7waxtL5tllu1lKX56gF
BwNws6cFK6GaUJxzM6GrU6DPqVxahZQ8LHvCJT2cY1nBz5NZAci+FWjYf91DPls5HCdoFkE5v8af
RQaxtpnRE7MKmH3KOqO/aGDkLzlwerLySxLZtJ4ZaTYrOzRug57c+gv4UsFXZ6MxBZUi/x9OZW4+
snBCi2c+cYdukP7XR1Oravsr1qE76kUU6jbX6BwEnY6iqoPEFBDeCwS7omoxEacVicYegTkeecUs
e8Xs0FyYGDIX09dT4+AoyefFbybgZEgKtF7m1KzNnrk/aT6x4OLBJD9HAzwKan6gFnVpa3JmMmFv
7Dixx4gOTRc7/kzfFafwSOH6cYBr+oy0PqlHZ5VZEPccbQpiRRKlCrXdoGdQ4fV4jwx0JbTuLv6e
iL4EpQqzbtliXAfR1lxH6XkY4XecYV5/GXGPUWYcGEushAFRUYDhAVVDnOv37Mc8kwG73Z72+stW
3yirp/K05KNyLZe9/avI+EtQVS3BFLFu+REhw/hxGjSPaNp4rWVpGC0VNR0LGGCRjOC2xR82CAjd
CeTxJ0SXy4xVHPYPQdRQRLdrpIBnl+1Txm2qYr5EhDuzdqv5OANWjRA57qhxTJ0CsSG9HeBWX6R2
V3EPN6mNfkrU1PWh29QHp4/aejv0xBQZRERK5hVCdnz3vKI2hEPTooi1r9HDeM8TYlDSuy+Ck9W1
6N/+Q8sIFfa3w3fCc18UidRjnzPT/E7BJ415gRyygEftkJ6Tbl54zL34avt52T28OEyb+QUdL4J8
AM+OcXmCs50p8QvQlw2QMzvWKQ/HUGsJMpVC9JSxXhYNMWNUGikXvMdpB4AUG1/SIdbhVU4MNJwU
cR4w1b8R56Jv72izvqoVaOXG5O6bH6S12Y2SvS/bM6ok7zBF3wB2VkOvL+tsrPTkmP5Vuj1qbDsZ
T/EFe7CmuAMYpvDyxlP1qR2skY4L1CUNbyikM9DQ1WJd16wxweISk8AcMCThjLKGexStvRQiPbzH
Sy3qni3GSLg0I3qArvxJ7AOzVclixsiEcz9YMTzq0Cr/nuF1hmPYA9MYNbT11NQNPNBT3pLvzM2N
XJDgSKDdKd2PQjNgzaBQGlL2GT8QEZE5k4cMiF7V/qBL/2Kq8ydYchc8TQkK2T4Qj4ef3U29K8RU
qvZ1IZLcRfkfG6cGPfVCXlTzjtp1EaVHZawNg5tAdHCEfKZ2XAUWvxb8P+fkcBXwattxoUA7lnv7
lpLoI6TyUsqT7U2ptck/eU9Isk1XRrx5LJ/ADXQfg+9zdRpQ9CuXvCXcbDKWMhQCC+BD/eM5zcxh
opKE3GjXC/XSQwaRd8oYmRClqeGWcqDJcT0+OhEafFILCDw4GRqiEdYDWonPPP7ACe34J89fJ8Xf
NGuuMEdEpQtz0Nkqrd30eeXpsB9V1vLlpgc+BPxOdkPzEBvORkOYNznbu5SF2G7yhWTdV/cI2XIc
aaAJ66gAGe9/yX12tD4iRgS3cXIxaSMwh9PFrx5JOp47lYmqIRxLKn7r3PQw7jcB4+9xl/HQQh5K
6akfyo2auYuBYTZWd4VDvLsHTBHL4GWocQehwo/CED9vREHNpHztFrOmPZtnQqQqR58mwUN2WkcV
9hBu2Ism1QtYpL6wCfUNo6dc801Lgin2o51TxUVc/y8Efej82z66yYfnoUA0kYm7bNoZFJ41TiVV
KKnboVn+OEb7UhHvsR1ik3c8aLNxVGWtr/Fga7TBM2ZZtTuRI15zB81qzgO4MBDWTXKemvqT6Rij
/TZgJc1RAEvhcmSC1aPckj3IteGEyfTJwYFiEgYuTiuwJtTuENJu1xbnBj9iIVjKGkhvyf9YpsAx
tagnOhoY9JoF+CP7mCfsFZCGlvaZcI1Zw/FRLabUVwgO15BcNjXpmEi+yZZggGHwCxhfnooBQJmx
u9SxsMSjnMPvkCwkAf/E9atcpLWep9Q7lMsXMyt9HiJJ+2lI/ZrLA7FZbf2VpVk2GM57qmumkMw+
pYvLgeBlzQEPnaYpDudPFbHkMJGwY86lL1cDP4+pPq+xp3WwkbjAVKgVpiXWaku2aU1yShJ3JpQX
5ACUZCawD72aRord+w5/kGb1GQHDyf/1eLh/SlZER79T/pA3SyBE50DGAEq6i5bqx+wUzTti21+i
mf/df853UL8gYdBx4dY4epc1AwkPs/mCG8XlxGxD19iV9fu8m8YZOFUZrjXTude+Vyndawn+2iq5
UkbD+we3ge6zmg7T+ZOUa3ChKDDaP4oK7ZObs9KOu8e9M67QdWkHgb7oQcracuLm1q29MMrx8Ap7
2S4h4op/MvAwBJgenJtrNNv3BH4iYSJ+Lk/x7XXvLlXEnmtEX2oIu9mpzz0HNoJeTR3VTR8m8eus
mLI/0SjIpJteZnsYwTK1Sc6sCRD8DJwqFRnXpf1hFhtyvu8K9AIAvWi8ohxIVxxHowE6dp25c/GT
obBnOrTGsjk61+OL8KT1cyJgfjiuHaDglO74MRkyTZw8KQWgA/vCE2/wZtKE62wo4HufqPt5dsAn
xliSy9ThggP0LVDZw2maR87O0+PBNrS8MKP0khdhaguyPTnI8vWXgyOwPHOrLcixk7BU1LXuBY69
Q+aFGwcFlKFaC9w6hdo0ymXu5PvbR1S9vjhkTxNFzNYcvtzqwwHZxljUYy1X1FSrhx+sAPQumtR/
3iOGdBeVnNRXFdxPlbChmX0y6flQH6yLrUJ4NvjiZro6GQVWpQQpfBXoxi4JGU/+4p0df6mzMKPi
LLTflvzv56rcWEk8+A4CBqv9lefJhvcwGUjpV7Xbnn2FWUSU3CyIRPtPqT6//2OuNRMJ3YzJ5kwn
kNUrfOfwZErI72HEaCqZRWgasTy4TAvpub8cEZd4PqxIgV+5f5ghKi9pGHuEa093tIxpDD90Nrp0
+kHNobuPg3TuRYEQfkRVT5dEZOcU3KpT9y4H2SULWUhxheg5kiMOcDmbYtF1dszwOPddzofYiz7G
o29FDitaDZckVSzBCP1HhNOuZEnQEsTSVSlsa//XKYg4wwGUo5FEZQNnpTiMF11/85/chETBg1mr
BKIybH+Wz/4ivXKD4JfbrRkN5Sogt3IjwOTEOePCHhcMvGO7rc+BFwfulS3VooVoIqPzHVEYB3L3
upVs4qNsv3z+OiMJ6kRaW8DTHB9XbpR4BjEaAH4AJ8+mzgacfnaXpI8su+XAnb6+DD9ZgenaS7Wo
YuI2y7mQ7MIDIvSeYT2uFRSImMXnv8jak14q3EmWzRSnmnu57xrG5FmLaPdlPR8VfGpCzmNaAlkl
P0hSfpSNwQwVkapQGD0EIOG9eUlUZuqXpTW4SG495b5EwYbW/qUUdpUk+21LLIb2ie9xCb871hWn
FE80LV0LWwpM5xPzdJfVYYlwCNiuBF51qGEFO657c9BxxuVot8t70zOhLau3E0khbbZchS9JsFJC
zodI668p0JmTbPaxUWpdAysWzIUPzO6Lo/YW/0e7dPOA1O4s0d/IfRgirpuyRxlY3R2p1u1Qj2g0
5Wj65CAc6Y9QpXnWydI7+bnZMx7UI4ACCdzayiaH4eImi9YZpsYB9um21PogOCNOkfnmpnZ6tcOB
j+mAbA74oH1zQWrldUzivI6xZv/J9fnc+9xgdPo8twctiJgEqoOTjpFT3SZMs00wacZ0Ato2g6X/
QG5TvyWtny1eB+Be2X39ro1KNVwAMwM27kfWgq2HYK5Pnj2PZlZyVL8ODGy2Qdk3msqQoPg1hOY1
DN7EvJgRXtK9f3gim7WTLdf1OSvDWANwolQor1za+ZZKjCVyxC1FQ4lX5hYTWsUyQPwhVshBjkKo
nPyXg0OSmYuwEEvanzI1AeTjKB26WAHkXzmsV+k4gs/Fd/n23c/3Nj69OvwPp4d4gJoCXhzRPFsi
FMVsseDRYJFmdLfuo9tPbNMyaQ9Op+AIwZEFTBVs22vyJ0qMyoXec47Xa4qqkZY3yRRo6lgPxh4g
2xpvOz6i/RLJw5cteGZ8LmQb+pnZ512xZcgoPH6UdUNb/XlbaR/g9/WhnivOC1FNTUNj1Wflioi4
PeDdJTMEgOxOCEP4X3YCT0R1WsLPPAQ2IeuG3Kpe5eukTKmCJVaKY3CTr502RgRNr9a3FCWMDrni
GOidu9ZJcd9TWhsBUclAPbFqHRVBoBW+48EUpllj7aOYwG+YSnGugpGZFdJVgRxWc9KnPIitL9Td
QjMwXuzcbpgdXPZAcDbtfPwQr5A64uSqzFT5lvTErVceVKTHu6mA872VqFZNJnzqKYuz301jQ+vd
KgzHSsrqKcys4SJdoRCXUrIJn8TmGNgdc3PS4Pv7JzKA7XZC9u/nm5ehLCziE/gweFqRi9M+CM30
yCq5vbfc6+h463Y8NpnJOsk34JEUHEN/YCgYcTcAtpxoQuQlYcleRVDKb++XaSMI3qi6MrxBVSgM
Q7Ivs99HwMHWfUHVt+Mp1U9HSuxTNdP0KNntjtK+9U/70WWicBIWJKUjmiF0NO0elSdz0cDXOJMH
AWN0l9yY6AAI31ZicggSlusls1Xr8DlNmMka1EhGhLrRV0BULFDLyx8E75tyRIkCP0z6Coen/6xS
VaLcwgitKdUZo3HlXKWitxtMjA80aGTiBSP2jtgqMcivNFKZq2fzJhlgxZIJHz6dM8iGMiPii32C
NBwylj1aWimcoIj1eLetwsQ8KjjK0iB+Dt3EYIFXoOJk3oxK/u0c4NjwVvXux/HGo7TYSTq9qj+H
mUh/lgEicflDPORQ68UdSFNOWAGDmXALDQerCn0Oa7UyrbrlACvP+dvvPKqL6sKnj2J+GraT/MJ3
El006ixtosOl8jftuD0RBwu+u4W9E65sNFwNH8663Nwyu395jrBuhQrmHgzqXTqP50yGPNgFs9+O
sTAB56AUkhnlxOqNfVmymCX0Ooh06tOzHDvD/I3aXcD0Jd1jJan8xnHAUrQZAzhFWjp2qsAhod5h
P1KEM8TwCkAfxpNnntcPh8p8POJxYCE6eAUK9+5xz4mFLWeUkVDdMUGt9PYCsOQMqabKi/ly39nb
rOuvkkXIwntG5v8sXvbYfuKsjIEDY102RUqEGw/tZxfzuPjYww7074Z7Cgnp92YsggjlduPS4olL
8euETgVY7lixMYvIHi4kSLn88kiQrpcDWrAFMrA4PUrUBOpI+1JHLOmsbO0srHG5bLovJHGOWR8z
68BytfVYnj0fLFh5KBK3oJ7SjvqVOfSOGpfzzUsmUxCGlV5tVJXxjn0RDZwNMSOiZo+G1sRw6XGv
x74NmJ21UUOdIQnsERud13pZiy8FXfwEifZtDYpjE+oVExvn59ygXdt3sw+MQ5veQvpA/9JenGA1
IoUrA4WD9swQRo5Qy9p8gZ3kUUWw7npRLeklD4Xxg6Jse1xki4kPM4aWrqChUcn7DS02R/SJ0jZn
VUK5QUGWWQBCbb+zDXC5t2bs8X/bWUSlxmkg7vzQwNcTUFl0VYpUq1eSX1IRqutDR5t0WKnBD2bM
y/hbzFD7IKrJIUl5RgxbIsar0z89ytP/FEzW07B12nXUBF35Zkts44QqNovmE4o3By9oDcS46lQ6
wiOryv7tSuplL4MRZ6rT/okgYmnyDnbkPl6zNQ2eOdmKHD+uSABoq/0GwgvQ60sFXJQZefW7rf7g
qcV8EErJSWlT6qroW4mQepOWJTJ3tRjpJSWb0uebEQSg+7vw5ZkmNU/2e0IYuuIjl7V6ZagCB7JQ
NPGufms1wMNNszfiIgMB0lHqYMZqAKbfcKRS8mbRNwulMF8vcMv4o2EEE18+HmpAWTKjSqk2Y8z6
GEfPK4Kn6jqgpiPaB6GFwD8XKCSXru8R82GcSrlCF/8VqtGWWCLv9x8Hv534SZreDpNyudNa05Yd
MiQhMn838JlTIe4p1NSEtM6qf4w8pGNLMF8Jix7qgDPVajxCgtAzc0yy0xMsCiSpGGqCy6tO2tDK
WOJN3oQVix5wluCKnKaxbHdG1pB7bAAJI7z3iFxPCTe7/qJ5JrbWSrKhBiDibutQynfF3CcQAt7g
fvTOA9TT14I+CMdqLrqXYzYEozKd15Uvhy17WjDeiN5pGjcTHIoYD/6YidXeHOWP+jhnS4UHhp+b
F4TsWBsamJIJf1FrTdu7nQdFRJLWm0E8ib8q0OXBshd1Yt29N7AQO8LzVtQl/bVqcWt0Gqb6jY2T
isl/b+JzQMuZ3WU8WNG6GNa4V8qhqTRUJU+zm/HK3dyOHyi5mY2KL5Ytignwtgo5FGkkcfYuLN/W
+kp0FQSQlkZb/icTj7PoBd5jLQeRINQMZfXUmQs6Eeh/HWLO8JFVfJaPHc89+JpHZpnC5eDGdVTx
CWgr3u8K/8H7wWuHI7QxMWk/aAXzbfrBBptgCwUDdbVkdKPL9GNbc7Lw8xXCjC6xmed4iFKCjfc9
ndCM6GQdBKq54j+jcEYy5GWCJo381mLNbStbgzzIyHJzdC7JIuQXsPVHC+e7gabZW2diC1M24Evv
pFOX5hFO82d90oOE4Q49SUV2UyQLJvNqFLGHOSGq3ko1LgQ0X1j0T2Bh5WbAc6uP7OI61ums0y1w
iGgVIeZj1Wb7eV4MrS4C+o7ggFsTsxk3QS4WnES54g23bGegN8N4vc5WuIKUZN+/udiTsQ1cI8qc
KWE3zYnp55/Ptx2URJq41423lCkRJBecF0xjPsLG5IxyWOD44VH1eEGTpAyn22snShN//Upy5ttF
Dxps19LOEFBXEYJVkJNXnwEtuBJjZOD5UYSHS/pg4JKpKyQ6eHWWOLmbBUlmCIhQaau5PeGuNMoz
T0RjfOWnxZoyHCqjzUv7LtgAegWBEISRu+w3nwVK6MGYDcKDMBX4zKZy3v7qPtUhIXCprF7iLsrl
8hSG7FGKgFtnzdxD3HWE+klvlQzxsA7cc9O0PQunY6ee3z17ROQU2z6jJK0PfgfOsWrNWMpAhMMu
RDO2CPg2TF0le9lxd0901UiDfTQZQN0FpPYAChddFQNyIvSSvaRQzn9pgHUO1dezlTgn1Bl0oF5s
Xy6f7hOuJRQEmOgk7R5KIq/YUv3RNQlfUyPJcY5lyLYrtvk4TDfu0ZOsHQ54rHyB1c5Uicjwd8en
2lxgHyLfQa7KBV26aY+oKhSg7xE0SZthNVc7NN7Nt5jl06zzmcd66zqxyfXVcLilDk5aYBK9f1ei
NL9kPNRZf5hH1EKgxKW+DNPCEN6hGXxCU+M4yt3aTQlr5El/Lz4glHtcZcIsAMxxqDVnYB1JpP1M
MYgFIrbiuBE1Kq9xivErxkZp/vBbCNu88VZhdOtsxqKTGW9DfSTVdnvbQAvoEKz6f4D0aeIeWMll
WNWCAnfIVagNNunQw/ER4BzR326oFmLJLHhGzGqXBWetxdFF1Bau+kuctka0SECw6whPE7SOgGiu
t5EX5tTLrIIFwugqdifKa2EbnXY5nB5TOy6naefv4lsrEZh7ffGShTyS2nExBQhaTlhvLMwvz/mu
jAJJmCabtZAMjeL4ongeqqD+Ag3U4jXI4xX4IAax1KQgjjyTun3kFVhEBbc6LDqTAsZRcB+QlV2r
Vv+Ok9+2U9uhRSN3F58IjwITAxblpa5SQOWRmjRDQkkk+LKqpspZZN1H0RkH6tGAOAqkzLrTdNif
ak4pJFgNz596fNkJCZPY/NNq8QALsabJwNRtkEpEANvmHhSsrXr59EQXDrLUzezsD7yGB44a/2cH
5pEP6tbWNRRYfILrHaVAL93bMApZvpZTJ/XqcV+ITGd0LHRJJgy8W+GhGTWQWvz0VWGkDqmGEG2b
oDkZ2gb2vC0E4JexIdWwhTZoTZvVhXtDzOj3KjQH8udAifH3ZfK1HdPw/1iaBt2HR2vKpZl7JGSk
eP+G+OoqfRKWrMHoUG6loECVzJQt0nT6oDIqPJlzkD9J7IVF3/0CpQ73PftTrzqdLBRuSGL5f1h9
wrAe0pX4uElyiPs/plC5xab2Wz7wbxJBvk20W8+yyqLevFhQjwt86WXueu8IRRj59WjU8MGLvIL4
b4A8gENLkZHzrnq/ZkYeupihu6ee9/2J0jn29pacysjl101BFNx7NmFyoGfCActKXDpok8hwG7Vw
VmjC+OxUk0xMzIM7Ppz2Bm+uTnDIjyhFxeFipk9gomeoRfRFMNPg0a3GQoLDIUCB2AkpEoUD9INk
N/tocN4wgmUOsMssZlis7bf3yhAsK+XTTS7xWr2uTYfDlWf0mjLNjUM2aejlmJwgn6lf+yfKfvAU
s3AimA723IFsgSqM9tIWnIkThnPZxZ3AhiyHh7vHdWuB8FEYyb90I8OcbjrQaaXQWf2panIjdFO6
q/8A4xS3MJgWT8/WPvwd1mMdld9VGYlxH+Gh8YAr3JHGqaa1Mj19n9SvBoRQkTFxNbtE2+3G22MZ
0tRxrLxK6YY2ZhRtcl8/RjCVOhnERIS5onGqrxo2bj1FGNbgRAGRR5/3rW7AJaOgqFEPDFlzaDIq
qzTj/LM8FJTGC2kLBqBp10yAsyUaCwWTE8eY4VLAj4V0ybrbPKtZOKsTi5Ap7rX8x58n4S0ZUAfo
JAbPQCuQeay8hs/3KZLw15F+FdWop36PmCb0+U5FOn+wfJubV2TZA5cnefyoyLw1lwZO5cwIvqEh
cgqqtsuDJzIcMBug77ElK//6Ge83QG46X/OxyOE/OONZwO2XXKZZZNlWQM+eVrbalpo8NfFx8QA8
U13uq2p3Hfp3Rjt+FvpxJYwI32IgjIy1ZifNHJD3KnwT+O5x9Kc5o+J3ZpAlyh7bA20/itan4ous
1N9s3txm0gZzgxGvXmr8OYT+bgr/rweSaolXkSqExQpkFabGM0bkd5R8ouLW9Pvc7wo616DIMXJi
IBDVAoXaIBxZXLDMRAd18wa1+jR4V7vSZk73aqLa8zs3lg56JdkBj4I3vwCJLwK/YYGVEMwzgEU7
j05SKJJF7cuQWZaDQruIN8r84sl+7Wxjjn4NtHYMe4EIch1Jv4oDZGdRc4L1sSmSzKVBpbf/WjJh
+HpZL51cw5FJOANZ11J74+ASa4RheHHKGXFyF6uVd6EqjEmtN62h3RY1C6k7+nRgfY+T77wjl55S
sT3E3nqbsevnNyBAcI7PtUDqo/PnjRTW/aFCNK/KNRE1eT8qre/QKliZXTIFcafOCn690C0QCxmW
ks21py+YzlhVz0qk5dgjslVElrdEHR5kKG0eBN09aeJ7EPVcFRIwn/LKgRcrlzkSkR/jmLhEGU1y
7Wham/R2Glm3SWVU/kXUiOo7vmn3UlXeTIpv6pRWYb2Ls97M4oCa4d5cCbcMmkHbjbkteN++a3Rf
YloEA39Mq4vviTyPVVps3+gatlgVnwSvLF8DHziUFOc0i9AbNPugJc5HR4dR+Rvo/J4NCMn+bciX
FneIq+pOKiMKnU0irkhLSvUEmC+9Sqg5BTm3q2u+NDSG7+0paI4FGCqmjTBW8mXmGAgJAHTR/1p9
3E9E9xIKJH1qFSWCj7X1BE3P5TIETXPNL1f9GH/bNDj4LWomiMn/djV/aW8csRHyGsE6s5IflzmZ
uhJJuvlWZpygwbInOM7FF13PlGqprVmNZYpeMxn+LufEyPlajB6SWZcSvQtS7AFst0+Ima3ud/XF
q4YHdcdYHklcET9f6X4z9zHYvgL06MgyjY4OhyRsm3mP7dLato8zO8lYO7VuZQMhi8DX+TBOFbna
uW4cuI0/bk5nD6bJ/9pMvHGRJ52IKV4baFrNkvKjk1bnKOTKypMaaOe+iDXuxW+Yk51/wBwearC1
qLasAmr77nnEk4FgjW13sWitqLUcT6v9gtRRdJ+y8Vh1jsyEF1A2IL4GFFEyoAezTc9IQBBCZp9x
hkhaOqGF0zxwgtXT19lkQohHIFV2UEQLncNUhnT4ExMdarzuYY3t9E19GhU6Qo7csUWE7C01QI7c
eriOtZiPFjRCVw4p5CxCW5vh5YlfXpe+MPIKJrhM2IzD2zlvEAkd8MYh4bXt+JxLWGRYFxkyOerL
xxN/P/T4n6bWVzF+0q5Z3bb7uI4W5PBa5a/CVw7gnWri/KCbClA+Lje4G+am6BHBLr/edEEqnqjp
NDm+9xCxBSZsuYVwj2vei00uG7Bipd8dYV+VACRkIxpoEY8+Z6jMLPYAmDKB2hJqkiRrVH6qHEFu
gWV4mH3QOycGiC4pQ627IVHhoSaaLRc+h+klfzckfKy2u9LfEgWlGYqMqWcADDziWlHeskQPPvF3
vpqDyThiLZx4t9LmgM9Bw+MsO0g0zTvRGgC8mTpMzAEi7FqCcOSWag9XrnaZsThAs4Ir3DV82ZQr
59JoQQ+2WTkTZnQNMQoOB9Ju7wnXaiet3NcNkxlCTNOB1g6S5KmoybWAq58DKB12HcLozlCJdL/6
9S59wLP8Z8/LdoIg35xFQk8G5tSEcZ1B64OS2XNnqgKeMlKMX1fcDp4rcN9zchVB6l2P07KOHuww
Tomb0Pt4v4afFEZdDS7bJwMwRW4Em1XX4OU8HtAsUTEAaesXVh8rDrepox55GsAUyG+VEp+8yhL5
Kem6x0Yln6rvQlY/MRcZ4NQrqmYk0HwvOJas/c+9aU8jKFg1Z50XfbgyrWp0w+fteXrnw671XHhN
RfiySy8zJFwVjCmti2X6b9e9Q3JoB1xLH2ZFI+Tc898r9ysQbhuyXF3Rd/XRDcgTOfdRRWq/vPe7
0JfwS3Qt8Y7m9oiy7tSuNHV24uc3BIsAWE0C/kKHb3a+WyVJ3+gseVcX/Lcxr85NhzQ6lMFK5KW7
BZFOp/KdMReM39fEZXlw01xY4tmd4LgVhqRb1GWPUeGhfoqysOWaTTtqRVMBj3VPbb8BViXzRrjN
e2XaXfJ0h8/+AaUFfPKw044E5xStqJiWjkRUkiGGEOixOinyeGSeoIChnEuXSNglwnoNPULnki6w
cj95PwZMXuofOLQNg2AmArASrAAilkzWNH7y0ZkZsNXpY7IuLMo8FpnQiFBm5E4kCdvdmlm+N1Ng
ucQSGqh1dHdFcED3/IyMmFt2BjTxh05kmO162CzvHF09ZwSZ2bwp4e2fh02P4N5M/yo5G9HpchG8
obKtZGKlJ0Bg1lSeXqXB62bzOYCbXXezQY4Vd64K6Y5DerBOJeHhr7xqvA1QFXhs++0DzhUoY4jB
Q4rk4hU/XK/VswvloD+qTLbzwpIfPS8Dqmj/blPYJN5v3TM78eMEJZMrn42zzEwixNFCWKp95EPc
FALrK7J8xHC+c+HsTTvzVL7lNw9bDRNiBsIWgWrM7CWdllFLPoMmcFeAJIETFqDGxZXUd57h4085
I+Zx60HQjJZHXXha8RAcZoUet7rXzbJMoLtnLaJbBHY0nbVlX/mHhcYk2DdOymtWi9Np5/+TLNSl
dUgqh3LkQ4r/kpSnxmeLTGfNL8B8Tx/Y4rODK+xRCIRurL3DmIu2YPCOJRRhbDIRUyMaNdMV1P4D
3YQHWyQJbe2mGlyuc4TFvIRe961W+4TGbfx2/yp2ysWrjnNf8BQg5bAfTf5UoZ7Wk+zn7B7EK3or
Jh6cY+GiXfskXaGIYGmRgcFqslY7j2PPcCtpAIceZDK30Ib4zC/UMw/yJT/LJHjXeoho6kCN3CU5
xHefCgsYN65X1FPA3Iej9FcyTtzbklxDpzt9jGK3/68tifeRCsWLixv40m0+OSCBxy6VBywaj0Tg
Q/zwpvenhRAD1R42aQL76N3ZOaCXUOxpiAguiu8KLe4jPxHrVO1d7J1Z8c0sit9/o4efQeFF3LN9
zAzDM32x7cyMAxSstpGVfpYvFLZx/llUJ/Qf4s+yqw1q/aeXmB7pzO0PNF4T8/DWEp/j5yHJWqiP
iV5rERnsSOEL2cWFDjMRy4ptwkSCPXAhrBn5VUsVu8jxdtXUZ0AAM7o21HjfvavzE2m+W2sivNw7
NtIVOM4I1YkdUSc10ySxL54458kocTwzerZuWlxC808EnzziIrMNrZBG1LvjAwNX4hA8rtXSonxp
3qdI53zbMs2lhoLQ4hMUIGabYoeQpiHcK+UE0+TGXaWLsO6cvBa+PK03Lk7CUN+fy/0qH4Zpa7iw
FjZ+vGklvwushck3GZZYEo4HsP78PdHTpdUE4Hkk9ZUGMcqy8PxbJ4k9olgCdEXu8zpMTBAV4S+u
q1ZRiM0VM3kjp6qxZveHq2wxHfNxmMCIx8QYu3MDaIF4C6WeryHiGgcQXudbe+8gxDfhkCOzvbfK
bOEyxQltxGPKFnt02obLhsVfu8JWBoQmFKdMA5Kunnp+0RO3CTe5bMwsNp8aZsZ6IpBFDd5CrMr9
q/BYI7pMQQhhH0F2G/fyvKtKxxYsX6+Z0JsqbtTphGQJR64k8XAKnFEK3I4/xK/yfhDxS+bbHGsE
A5GoeXD3op+Lem+jCrCwJMGhe8qmp+6f8N6RdIB7IhXRmBaMWwUv9cOk4sbkLaveXvJGAHH66Tep
JWbLDyIfc/fssMpqJutj+TKvKanLhEls9x7yIutvCkOkh0lfB4titMcghs+MjHzYNSZ/6KTqH2s0
7i+olc26ajGrlFMAI2gVzT4jBOvEPzweg4RYKXk/+erQ19sUmOrvtW8zvg1c4LZt5N9P0zMFQ7LN
vOMtDLGVqR3McdkSUMxjshnHDKhC1+Mj0l6BBxmdzimBUMmy6+v6sO0tODe5SrFyrqr78PX+yXtn
Iv/pr+/YVBpdZEUJm2IhSS7Np/a0SjSWV4Jt6X64vPG1YXZvL7uSVggoLrJ/V5e3MVUA8trEM18c
6A7LmSjam3FCqBZppiPpBMtWYt45R8Hxz+fQzaGayjbzYAfhgJdld7Recf9UymL3mYM8wmeArms0
EWF5ibdeHEjqmbnrtCIR3CQ1RJYZ8I1oybZIfzZ1B5gX33lIy5VeSsR7cfVxBPp0NeWEaslnmpsB
t0HzTedItmHchDkBERdDkGyI7hgnvstbqmkqZT9W9MX2Aly5b45S4Om47m57YkJMBW5KNc9DhqJ7
7lk8xinH19YX4U+IsjnWkNaVz0ZrLq7HojcsvVPtztdxGzrZKOZm5G6PZcX7jeknHPXYq9aI4dFi
6ce7W/LT/CWbIJNYB6Syj9ze10zC+BKCIn+90nJSU1p/SVBXDo/IuRjj2M07md/iZvd4+7vTDGgw
ryMKAV9TyXrCxaLy3pYsm8owNN3UMzkCB66wQMrMxZvXlS7PpN4iSfBzzOS6nbZn+YJi4usJKq33
0bkalZgUZvDl/lNiu/HRIGEpHj4uFCxOwWRZntWGpY84r4+XQ/p5QvUw5gemlw1HRfClF+C/abw5
Fau6GgrD+GbNvpN/6TRhNgouYtS6Ca39pLpD6wSoH4TVfvb0qEdebtYVhZs/A/q2d1K1ekX6p+LS
oEOSNQ2CnQJusMWy+q2KozBukKBh5lB8n3JIVYlWTH4fd/qkLWnAP3dIu+saueN4Yj4wYabi5YaC
619tfCAD5IVLt7EKi+VRWJufeEGJz45LxK3M6HNE3kDALoV8DBkGLoAnUojA9OheWOa9wooe4QMO
8y+J1B387ZKFCsBNQ3kK/efXDfIpTlBBDj0LlvS5mIHZSetECa1rETJgvN/yUsnWOBO8+OC84sAT
A4Ex0kI7QoDGenHn7yeKAwkCX6+nina7kyRu2zpUOc1Ow29DL7pKuYQj5oaT1hMMKKlb6qWYJbYy
NPwNBw6+ndY5xggKGLz7ko31FuFACiPq3Lo7PQ5M1px6G8XHqiB8nyo9R6TlMBXZvVSvLHooH08t
YwEt5XUzbEm1ZEp6oByGyp5gj+73R5YK6doRMXQDp+G83ZoseuhJQ93HC3Q0MzlgKllYk/YEjjMp
5/UmmCD7F2ODT79YtuSLKQ/3qs8DxRFXYP0sNILErO+u08AhaFKmoSCgWcrQy5bXkMC1xeljMdQF
o1HiwZ6cZWecQN+cfr9y3ONqutDi8l8qA9GK0ALm/hIpxTO8mOwKass2pQ5glwqarDV0GCvemluM
yTXdVz+NT0DzNzhT0LSYaoGHkNasGIfy14JQs/x43JodHZsN5nKuxNaS6wqEECmjan4IYGkpQq53
GY59lHlnlUb/55KtCk29ALUT2UGtOwRzfXhAAV0NbNisLnGBXBWyGfUD/AS4sdKA7vrBjxURv8es
y3kA9Jpo2vzHjL1C7Yq+c36A6IoMWMmeBVCoITZ4WUqkboO3Bd2UkJWGM20NoryqOwoKcpUfgdXe
/44nc4lIWPQelhbVeCVTX2sCEmpXVbqxc2MlKXesY+OdtgzGuCqz2iwySbd40Bb9DWPTvz95yPKa
PqvmUVTkqm3F2abNX0noPbZZ3iwXnosFfn66eaQAR82QwAQcKx+ZAAypf33Hqe3x5QyuQr6mkBj4
U9sv0D3jdXe4/Di2vKGkXrwJuDEvGLyyGQiJJWVazHMaMwL80vpusqYPCGcsZcjjAuuLsz0D5TGC
013rhaiJD1hwHwOIZTByFgdxcLIUiJx+9bYmp9776maOFf942K97Hv8GIQJOlvtGkO2UYkKWaERz
E4piGFa840CpzYaSk/V0DNm2FUTdpNeaoyqLSotFwAHuehdU6XF7E2rlgdvVIMiSWQsb5ZjlJuHY
2UsVryGUOtm+IdRjOtwZqfFywUwMtF7kego/u/XNU4R0MyY1nicwDmuNJ4yhS6+nFzc/AVuxbMDs
0BbMQjnk0unS5KgazXfoptnwlYnMKI/0qmqc6ecdE4mDzWFd9fHPRNcKQawSY5EcsjoinLD3Wr/R
DQUNu66sjPZqp1d95IrOmuR1SwXtTHAowG85S1N2hni/KBjhNnIEZWH3wHIHg9JjWdIA8i5xcfIf
SHExnpLQJfAqTeWseYy8LxTjwt+EuKpzhOKuHGJPEEsb0JR48AYtKhWgVmnqh9X4dW3r9+s/dPEB
Ci2soB9ir9K5rtGGGfQW2aqDqAyMNf7EHtZHz4FBcuMUeRqY85OIl4wQMlnU4XcLXvMZvwBK+9N8
+yTAY5DK942sIfAZq9ve4I8BsiutsQ+xRlPKqgjK8kIA2Nk5UxulP2m4EZ9E+G1pxR/5oYw/NMM5
UD2sVRgfzpvJoRgx1I9+h98lD6FPBkP6rYFhchOYyK7jcEQ06a0ghZEttDKQ5BNRzELWVWvKKn5B
XZxPU8Q6ky0dPX4qkaeul7QaNCRMu+F+XlLkyqxSUoPWVnT168SS7neLtOZ9YNcMh+XFwV+/2gf4
hsdsgiXZbQNugh6hf4/wipyTa6K3gNQLQ8vPQrNr5xd1bHSMCwCK7uPp/5OGtc3OrVj0XdgpRpGY
MJvcSrepiJJmbfHj5rSJzH+T4c1b0LgFhlRitWg5hhvUjawOoTRB7ZkEN5lAIUosAQx/scru1vhd
MgQaW03+JntArPwQ0vYzSW9+ZORvUx+rZQOb/qE14OqFzzsQvF7cnKrYNX920F3SliS23p1jakaU
G1vIHM/6p0czX+BpbGNEZ2QEs3nXhMBVlZ/aD7PQS6n1pu9QWemgnLDGorIKAV1b7W2BMpw0d4Ze
NrHOFkQ4b11ddRlwwlcT6DcoiYwIJO85CUQDJVS6/q42/8OkrVOVr3aSlcvE9xq3E39sIbfaPmDD
PoKz+mRFoGHSKz1conM0sN/CnO0xmBBQo4KGoJUsLCL1xA4/JPcG3iIpxLXqLfOzUrg4QmyJsENO
n/S+FBa47Wfn3McOmsuycT4Hp9Oab7ybEy43euAJ0Njh1VvTOukRtkkPHX8UStjEIObrtegaWAcO
smotjHa3ZBBsIaraCKUTgWyUZeQzZt2wYjk3ZiYugOxGmGBFRsxHLX2XfJY36W2L7SBv3dMLB5TZ
D2xzkuPTut5v441l3nKY7iU25OgJ4WuOyRMHSeFXHeGq2fJyiWwDw3m4puLsdmeNEjmzecjti12X
u0vL5WyAz/oeMH4MkDdEaXDgMljxLpyabdKWmKsRCvYLHnnGD+vmcrY0OIKFBhjAjYyu1anOtOF0
PHosqcwxMra91ZoE57WdE3LhIbBybjGxiEp12J05Yc4pppllbpTgY5MlOz0evUuAd4tk839PXfQN
SVWoWhCtluupBJQ0PTk6AaWhFSjBpWvoMN7FHQdiIN9wL9SVcIquYjfhTmI/ovIzssrC7yt4gbyw
X6WHvpO3iuIEcBm0tjdqZ3W2q6dRlHQZNehp1T5dQ4m4hakhK9vHE6YuE26BBz+e2EbI4igqKcJV
pjcOwLyf/nadIcJf045DAAxcRbCva7rsBFm6iPwa1fjrwES9NtibVYFSKl6++HCfccUjRVmD7YxQ
QnaBWWCGETbjgPX09G+BAOWMxTJ0e7SKh6s1j5/nArOb6CLn7b+TjKro5Pc5sjamxprj7YdfVpDS
Bvyax91sW7yfUAc64llMBnxAGsjyPchNlU/7Lm0f1kb8t08VxY9yC1Ofw+HgyS20BhlPA5ZhFf75
5HXIUf8tAwhheFt/RFx+ceq81emVDjHnFWPJLwJGvw5AsCoZIauIu/qnAZ7wwKMQwAVsXmJo5zAr
+4q0Jl3x/4t1Jehs6wwYsEBbo2O1IrA8g1GNSgmSF9ovb0kusIbGiEfMD7BA0gQq1vcHT98P8F56
HQYB+gOfoLy2xrzm+MoU94amVWAgE9p/JNL/GwwxtJ2T9Qzp4u/GFZZX+WnS9yC1GJF6X8LVXrSL
4PIXddn1+mqLwLu6zjDlIjW4PxG4ayGhVIBvD3iBMtA5rF+VjZyxoJrhmcGoyKtupKelKmmKGXyG
P+6wUMB2DZlIPR79zVwxi51FduRRqQ1siO5E4XMs6eD78J7uGIh1dHvxUsM6PmxMthwiis3akC8A
ppcEL6ciObQZbPVNWPO5MHCz8SjbA/P0ITYENIzy2r1lOvFJbxIsBvgN0vyB85oiBP5OXn0DwrKr
bLvDcrRM2eOuivbY0lfamjDm1jX3k5g1B6d1jnuXYOCPYNqqcBYwiBSR+Y6lul4+Yo3QrGyCnkxT
H9QHETxuL7g/NxfNnujS9xIJLucKxpXRANSpLWHfUn/VIR8i+EEecx8S/faL3CrN9D09891DQc4Y
XSLe2117G/pF7whi4jpskPlyKrD7XyxQ6dIyp3vhanUH1d1X7ECp4ZyrGSEw1Zl9eThqxLyiWqJE
OP1h7EeYKCRvznwMghN3V7Qhp9xmyxs9rxPMHsyn3ONKmQ5nrzPOj2IMXpbpdq5nTOYXMAUG70hj
U9TooZNRmGjlNuzKmmzhWZL7+XeVIWCsjh16qAYi3L5lbQezIQqmMHoi+3SvyN/q0n1leTDC0cDb
5BhZ15fRJ/Hm7djxThWu4LzsFirutjoxTRXZwCxkDtP7K9Bto2VEvvxUHAiJvPYgcgpunGOos6bf
gvLRgOCvCB9PB7AYPk6FTxj5Ekx1Df9fSd4z0eL3PM5t/8BWz57vD54a5XUuneHgcrD5IBw1GagF
EV2Bi9UNzsPVFBZyJDKm4VbjZmX+xxUevPwg5CCX5ImqGp7J63UTSKMl0m3ZTQQE7TBrSSWvg9rQ
JUz0tDHgmxFXSdnedzlDtI+LOHiGwh2sRVZMBG0htDC8LksXawK3jm7/xy2xsfRmrJhaMWEcMNO+
NCHt7rwmjZrikZcrAg6luYgB/VbkDoHSGkCoTmRVM8Y54sCJzmSeSJpbaV1ZqtocI0P9SiCgU6hw
kU8+FvblSSUQYLdfPSc+qCRNNwULX/RghZMwsS1cHHwHbfPVs0r5yqHwbOYWE9MYtGW42B+ZJkvJ
eB3rLvEb6uoQp+p/0Z3AOt+867LlUfXG5U4t15eyBrXUjUEmEEleiZYjdGyij2YhomqqOgD1KzCa
dunUYayg4aBfiL3pB/TQP8E3mbqGmueI/w/3XvBYkBbgMGPQLiYnZ+br27ZCO08M5hbWMsjlIDeh
b+qL1Qh97G9Vkw08ZcW4x2o+D8qVOPMSZSxqSwb86jRydfyiprXUoClwp45iXsrRDqf7JXp2/r07
BOkvbqudSHtg+kW5qv3loAxSq3YD9mPFCegeFdPIJaaYfVdYNtzyZ07awpKRnlL+c9vUFYqUfyNT
P+WXGnDVKq8QYTfNTGTy+bZeaYcgHUK+rcw0dnQ/Tgx2XaJEa0sxZRyMfUDK/P8jCD6oBXIVG5vT
h/vs6OtJVrzS/84ogom8kUnFlkOpTP0vgiThaPw+bHMMwjpplAffjTuUKDzYymefTOP3tB907QZK
KeKVl+OjkGzUuDAhwP5zxeFuV745czsY+qdFcY63WFMgiNUeeckzDe0BfqWu2KG0ft4UaBV55me6
J4Q8g+PPOQXsbzsuXDeLcPjlvX9bVRY/7M0me27dnoBa4dPyK752hIgTWG6Uu61+k6cqMxrUneDw
IVAZ0sY5hSBRq/mx4A/m3QXUa0W6NSE6EOqrrrE4ejmtrBp+ejQqF2K6lY+BIAvVtiwDBpO7d0vb
g6Binv1GQkBJHWBGueFuYHG/rz1HvpPlawfky23KA/VbPEXiCZeVGq7YVf63QRvXAdedo94dR9eF
fIJQqoobvwtJJkpmT6mr2qzzmBNmiu7oP879Mo76lL6/jOKdFgxYCfmW83DOk9f9SAs+V3ZM8jRo
Yz4Xi+fTFd9mIoge5TwAUnzCSCN+8vr3y38f448C2rBnB6zN1eDdov0T1fo/9U0vyGKxX5FGSq+C
8XPX3sdbkcuWJd/n7ZpHQXQJCEbLmXv97bRnztxhIqrbgizRf674Kb6bhhFLaJbkbFlg4L/8jnZf
6dzauqwZKzQ8Mcg0+kF0vn5dRSodJ9jySmlw2k7R7JVUBYiHj07WK9e0G0c3OoOcWyCZc1LgqbKy
NjuDuwwLPvXam89qkc4E6AsxvvGOqTAShDOlSIf4/eqA//xAPHdSTEUYiYLwv3HLO8iLEc/wLIUd
QR4Hpl721F8O7COtxwYdfP5h0gvOUmjDJ3dBC41M3UVVy4bfa7k8Ld6vsMlouYgYG+Rj5eISIifL
7o3aQdA67NuEQbsp7NTBSKZimnwjf5vMVZrB9xORrWY8MKylK1yr2OJT3xGeRA4lNUQjacFNhIsC
cFjWPKs4g9qDTMw4pbDh450wI8T84AY9wyMslkqJIKJ/wkqYB7IZ8oDaXL58cfxUNjl4xuJ2yht3
LuVxCdM7puXjm5HQ/NDGhUPLs+4IpbMk9bh+6hawRNpqTunl2UJe+23FXwv3UXJnYNym7BFSoiIr
/iW7MP9Gmrtm18sMmpTxw85Z4oWONEFa4/gEk7y25fFlR5bpg7kJAGxizm23R1CwezHqUraLc0uV
CvChqBwx2fqqYg3iXfxL3rQmPm6yb6G9VrIEiwSDGO4QflnUNqKip+kHfS9Nk8XICDTFzvXUYyaN
0pBmzS8r8NCjP9ZKvyBZDRfjkSuJ+c15603xypaWsrubqa+8tkPbSE5kb8QPWc4zghL+Oq13UGEK
9TAPCwJ7ZDRXKWo4wZN41H3z/0K2/jD1OSEwUFsvhF5el6xcI1KIA5fh/6RepN0i9Qr/fKwss1ey
5Y9RH72hy/ZkXBir+e9JY/31o06qE/VEoADrNTcF1+jAHlGlvXFhCaf+PcqeoKS75CkLewNpaLk0
cBFmv+nYrm/jjmN/Q4RZ2S9iPKvlQfepVqhllFKxdHP2lCQQlvqVrw3iLfC182kpzxxXxCrSyEDE
8CQh3TtMXSLXm4g20ip8eTV9SUKMzhzx1Kprvw0v6UQ+o6LjtBE8pdKoLvm19Ic+nKS6Yg1fMRgt
7hlUYGJL8i4S0csHgGOV7yEkc88Lw5rPQtXHRwUuPHAl47ozkDEEYfESDvnkVK0GJUQDr6ib6bzl
nM4Hpr6dle3Fq3qDDGl1DcNZsrjdYcM/e4zxcA/YIjdAg6UJLGYX+9jGtCwOE06zWekBHhGDmZAA
AJywGHzBLFEPmEesNkGdna3nyRQpiNJe3dcNrjvIMZH0/N7MbXmw39KIays/E2lK2jL7LxXDPL4Q
Oyy6jsh19SA//tKTVNa9DS1CfaX9nEjgG/tI5HM7/hffmlwNezC7jIDene+n20N9qrUNQ8zfjSMK
gJINouLndtTo/jYdF1m82P00X1jDOCcbKIC+5IpzrMpf2WTRl60y58WOmCYhQWxLIUx2dwC2iDCe
1R92wNx6K8bBh8Mzq0qlC+e/+ZbbhlML3d7pHU1bMTf/qM+gtAYd30jR9nfT02GkHOy7BG0rQY32
tiYxWkPnjkdxNLHzEbVsEV0CFxXMyfzh+b5vDhx3zJbB74DBKyXgFwD949Tx8wwpmagUvg+YIpFl
poT/ayZBSIFA83MxAglfwVNG0NMHxEnX0QBh3TNVF9GeuvbRPFgirVvjclUvg996utkasnGwMGjT
LjcsVc3qMTE4pnm/SFURu39o0hMqIierSh3XKYlgGJcLZkrCOZq5pGiYaGxEnL+goNWiI+cVcCfn
ddLtJE3aEyowHJq2yMbXyKGE2lpO8UrqOHeAE3Az8Rq6uDgClcW28ghrvFHPgQaNO/RlZ+qktCvs
k15y95wFdVlk1e9hIbRN3XeebGeRxtyfjbBxz35wmu7CpsFlB+3yxBYNJlFM/fxZmCNdNBAm9nha
H6xmRjNMO/f8YAr105/hHxDgx4QybX/Ln+l7/GSTXfYwZp9dIHDbszEV9822dsIZddgZJAfng8/v
pL7O8FwYvdM5mrBS9ZYPdEtPUrfwIRyvLS5HT0yWMdX9/9Vrzltz8IJJLCclmvtGmicZq4yDMOx1
h2WVl1cxngGCct/sJlFSz3zO9hUuPcLaHfDRV7Z9AKepBALqkIGDFaEgqUmvrij5RAD3f8Bf+FzF
0DKKlKYstz0WDzPppAEtzJwuzkTkqtrTmslC3g2IaAgrj27WTFCkVLhB5/ER+4XhMzS1JBefEvhX
+nYTQPo/BR2foC8ws2XUfmilZMlO+ak+1vnZ+sO2a4Ky5u8/G0ZmtNnjRcx+EE4aZY9sEHjVZjJv
1TRA2iMpzbutTgix2lbPGg/tJ/1k8OAm06P385bMuoHtIKCb3osH2uHVSGBBpRRacxktxR3ZE07j
ssuEDgWq2OTlshaLpNi31/KsVhIcLanVJ/gM6a+dXl3wTXQLh9kuoKvS6bgou026EhkZ+sq0BpQI
L7r2q5HijCxtOYn32UKdj/IO93GpFYNubA/WeMjm2okcQt0/xIefzlZtMSvIOV93mTU0qA5AGWcH
SFS5/2NGWj4rQC8CnIfraXVctnf5i3pLHMvdnFxFHfBXB7/21n2xhcDgclcdCNegl5rZQf2EfTp/
TRw6mbxEMAZS7OHHb7infegRDcycs/TrDs7BZJRuHiuFvu8MF/JyjLf41MM+3837+ww0ePAhRemE
qE2DRCDWn6aXnysGGgDKd77Ze3bii/pRAf+D2rqnwTFnbY8kTeMcZ3B8+dSVBddOPaQv0Sy1T0Ek
YkY8mrU/9KGulsbtak5EzghQwo9ak/RQZMxHEATk3izI6Lm4Apumhwb5AFBlHl1Irz9asLyOrcKr
yG+l184ER7z/yvNuHsbyglOoHsT8aUhFzGp+Uqo84N7c6g3GEews89PQPvSniVTK5yBMTw2dJ2qp
hMg3EbDfW1XHRw4gkyObmB1LKTn5AhxUVQNiURJDGxPwfelAMO5GJ14Qit0/F9PE5MABXLryJ8Om
sFZyJ10G/GOEiMGuQbQZefm+5yRcqB27V0Ox+dpVkhnrgQGlokhkvQir8VH0EwGj1TISJS/zNEtQ
G7oBP6z0IGY89CaO2ULNRRayj47s57lO/ZLVHPD4ZbCfKQSHCKyLXjR0bzvU4+wWr3DRj1s9adeg
eAcjoj5DeAkYPyqaGEds5TAlePTLFsttq06rxkvI2H0d8T0GrUsZAYbnAn0DVDtdxQDnIt51R83y
FdZlXIcCcJv7/hbUekQqssczv53SUtWxualZbeHRGNZ224N4nx+muY4+2CXbDqIQnY1Cw3mSb7cs
jPt6fVx6SIvDGCnxcsLErsh0Ayaofe9ZW0RofG+ACQ9PGjFCSI9us2WLzUpURFaIcKG6W5rEcVcY
SyZ0cdsJg+myUc0y7SPPJ2hmo7tkac9UoDveDGRHbczOcEFU7YFKSNvvSIy0qXEqj8I25ZcZpINR
/wI0ZnbQOROG5a0EGgFJiKvYzoM4pXyp2dZjuJuKFFWPHgh7e66gAEGj9fzuPryMyok/a8h1+9e3
023RhK59HtJs8xFo36mRpAnD6XWsz0qEGLLFCm4NiWqKoY5HUPDD+GqyuMqwZlhyalJefOJ6H01T
MZI2+MQqLRDlG9vku9+Ks5nBNv5uemIrZhbrTpoNqUVBHZcvSNA2SRNIAd+EwP6jloui90Cm80SL
Ixsikz4KlCE+2u/mxEAi3VejFSmE/iFErSHGqOnSxi2Pb+cwXLrmntiwDhCRRCeg2Lb8RahrCkU4
6INBdavNFs4cXNcEVN+F+bbsXLHwwBnL1XxhyMsHDG3GFj4X+nG4dRzp+HM/XKS20jxauys/yTxM
HpOL2wH7UTK3QTQmFENB+E4kjww8J2Zq9F6O5Xz1tVNEqVRv1g41HXoBSczgaptwnX+UPP4yyz0i
W4OFxy6yFb2vkVW+HendvzXRUdz/76e7cvkKP03iyw/WBlvRj57n0+FYEPt6DPCgFSIvb0Tyh5zq
Kx6Ayc6AO8huC1dHqR8t70QZT3AqMpKYWJ3vTujAhNUeUA4vB3x4MS910dIl60C/C9kA19Cy4s22
u1Mo17Tbs8qix+fr7npiPOFm2iMfU7UnVGtHSyb9p4E6WvFPKmXeqvvn814Ygo2XccLnux57bsT+
krfK5XDF+UAngdQmZ2wtZcZNrb/62YNvx/8loc2tsQRhq3/ToNOdkQ7MbWs+tOeTArF1U0728o7I
vBBLkIn/cyOZVooLC3IYwPp24uLQ5QwF28B5e0H9yeVWodwJ9gJQ68SbW8vF9dcPtbeeZ0IyrY/J
T8bSxY1/3cNXJqeQ1bEHx4DU5TWQYgJO7hEt92zDb3GhHlwaMZztDHultwbfBR2PWdRu1xu5L+0i
PufdlTsiA7JhG2Tv4i1obYhmMXp0dFz5ozjwv1hOTIrZwLUE1+YnnKT4GKN5ERbORb+diUl3lQqI
RGmhqEA+165ugqmyptM8HdySqmWUpT6NnTvXKA9X+DgufzuHlKRfAHF22v9ZfxURn30/mFK7rmiy
DexrJBv44pGNf3wXcXR8v0pPQJZ8bm+QFVnb4KaKijp27y2glFppRurbEoyhpsbUoH8J9K2mdMbt
CcSB3kcDL0OuDq4jEBRroo7oM/sWH9xMe4ocEdr04oqpnHb+Yhfb6fKjj5FPn9wKbrF8GegK5o0E
+KradjQXAS31wAa40YUEgjx4G+qLIalsnzDsxBUSld26TxM9x5nqebU+ieu8a4X/GdthPqZV7P/W
O+012PK2TaUEvPVtah9/Evxuk7Z3RC5IHsq2PWlum7AGcRvdobsWWy5+AtuKUjE81Y0o8BpTePMG
IF7XE6OXIM2Fbuv52TPT+2GwpO2Ooi1/pJPMSFq3Osr/TCgT5E4NnHOfYfmkOLBciqQ1UXFcxkJG
tkZt0NwZ3ROx30miV8wchjTInqJMMRcETHhjoAw7f5Ccs8eXEu0ETD+WWGFwLqObIzFCnjS2IwRH
Ol/vPYscxhRCByfHbDY9RwelnoKIznmupfBqFpenXDhIP7aEyU4VbVjgrsQCoplRa8EmTqlPERWl
RZ0taqJMxgySfFgkq3Dt5Vc7YbbzSJfoQO1OHecKuLyXmAwzxYJDPKnLCR/oLkfXaYmWM9c4mrno
KT2DuebRwEGHdYLtZlfsvJqY1jswlVWt99YLYq1Z/LO6v8T3uk50EKPnLEaLcqIT9+xawOEZTedI
/hKG1ueQbX4c+tQ6j7X1BgbVxNjF4eTmJqXWLec26sd5nYHDfApErMVd4i21ynN1Prt6InzH2qkq
0JKvh3YhGRKQE96hMjeLqZIMtg/EN+dGdpLY9p0bfe8W1pE/PzbH898ujQAOcWecEWiaV7AV7KX3
NfZX+40cIXukTQLq73iI4yewx+ZJ3+WHkae05BaGJfoB1MXi2FQ8ckbPuXuE9qUt0EPo+i94dyOm
QFdJmDjEGFdSS+o5sMWWelP0FEajlJtEM5vdlUGkCxYuT7tY2O9os2aR1n7B4XEYH2d48zzMUFB/
OIlh+unpkAT9oRQmVcw++XY5yEtHgxKbGgNbEIwbh3KS/+Elh8T9BrwXsDdUR/o2n/KQ/huoVHJX
pIujS+OegXHw2jB0qF+A44nJUmio0x4YYF0vw6c8iyZmbpX/wjBrQmqmdfoQ0xlxuHgbA2i9PB4t
Pyjw3wIUt82x96FsroxhsRgq2MNhKCE6kiWYXFOhs5UrvfUj5uDNr7kKCAAVigMkFaIECyT8omw8
YSIUHrPaWPV+sElRF59vFCi22S5ngLeXal2SS3VMm9IVmIjP0IoHAZjp5KtghdbEvPh++Mxh/5E9
WV9uvv9pEUl28uBahnxjogt1Xla/09d+24fRX+QD9xivsA/5eCvYIdU1vrbzi/DdJHHS2I2uXP4Q
KmtB1WI0v43YBZ2nHxsueqSGggshIyUBTdHfiN2Ueym8+odr0IO/x+SIN1IRPANlfQsG1O6hbmFG
yAHxTB/KYC27w0TLptx2KuNO8hyWkCL1dGKG65w0TLUvYzRb0TAaboJdUWkX6YhAQ2t1g7h4zPrL
NOhc16FGPzg7fY6egGuK70SMAREdbCDbZuW5PMq6axms318RoQWeXSbccWO1m+BH2uAs5pZqSzvI
ZZHmKqeJoUk6o1N66z6P56MBdMkUNCHSB3ulZj8r/QXvs3NqmEtl5NYE39G6hzTVttH/d3Aar3jf
ahEZY4TK5ejbtZze9XGpNtyFMqNKvl9sxZe/Bb5oi4gZccVsC1/nfqu9XO/ORzbS1u/7K8DNYXXa
IIF4VKUbzGbN/nHVTk3TCFBBQh/Cc1tfFq5z6fKIKXNg3f/O26v9zOXEWGv7l7qRTGWierwDki8w
UrYTQBX/gdI8QsgXPB8XUgHOlWyik4Yd9AIdww13uwmrm61n0DX7RCcWGAaihvCjrEqvNFdiU4FT
uvAatcv7Dgr7gFKjrY/YrGB8faWbvX73LW2eNg471pve+j3hGdAZ0PjKd/IcXZgMxwrLjnF66Zbn
q0jQ9RUGUU4AclOZNbkfDvTwbM0yKuuM7MGfLcBzSN+rX1ifMAxRSPV0bOzWMF/1YKTGpISK48Yb
AsArhmS8EEcb7fGWqP7NZO7DdvBwX04XgSIQM92eyJ5GzqH4c7vFv5SuYtFuZE+pjthRU/0iuB6S
OQVbGz9xN6KW0KCIUros2ncCTfSfCzAhUHaUxIE4su7RR5yMhJWcVzO5ZUVXffc1M26dyH/d9XLt
bh3Sh/FHHDHx6D2b7R7mhm8vU3NHDY0k7xnlIL2v2UOhP8ybWxXRTuxveWi4E6nlPflL63klVono
tDdPCgiqeBmOmxWffuy352KJqBMRtQFZ2Dt++9zWy4WAKieJ+c+vcQuV/SZB7EH4BpHjJH+ztsuw
W3ygbkqIFZIE0dORxTujfand+28VZsHlmxpHpdd/+2bndFc5zWLeOjXdfXu4CS4OlgMGKhF4dfs0
H6edPOBX5b+IHM3RMID09oIVdkFVCWaWAJdDTgrnE2POHua14f1QY9i5QM0ZtcSG82/SPpMBGt4+
4CEXzRmt4/vPAko2tgR+sQuFEyNKhvCTRsKFcY/fXIZrvPOXLo7t8NRy29Sv+yQ+Ief/LupZBSiN
yI9xLNw7HY6RCJWXsuripef/bTC/XV+dxoJV1QOU6i2dqXkCGtpPAkYuUzdT6MYvllAcIXpHdBCq
/vqycukneFmmIurB3tZzUrSjxDHetPKjoi00F0u5ebjef54mBTRBgdRFlKOD5WNAiGiF8PAMUPoh
wdqyyJhTPSZ8Q/9L+LLHgvdsa+bP4hzdV7QT3pNE1uizYSAPGAtJZ6dyAyk3j4qCXTdgyljCXpnV
ryQ/aHesIA1t9oHk4yPtOe2JYEdnuT+YWVv54Nz3rEZzQmdRuy5f3kJTJpbbg6/HHccODQ9VDGKz
6giT5GQDNJbjHNN9/0201v1sfCNdBGgfO2I5I6GdEvg+rKeNyR4CfQBggGkX6hic0p769aRycvIe
0fgp4zfO0mOQzcAV94C/t4hF4eLMF6ZA2RZwPc97n1PiYcwJzBmK6jNL72CuKSflyd4Oc6AWmZ0t
Bzc5GraRunQTUQih+xxWd/xGN7twHnCRJrpmxJAwFyqmFEzcjm9zlyAJuug6d0Hfx8EtnMyaML7H
7BHBIWSc1WPnzlpFd+JbF6Vpvk7HIVLn9ukKbVp3O3MLnFeZBGDtKxAhErjHKJ/wJ+EbpL5yJiwq
RV5zyKyWzWHcKycGhye6WPviKwXRsNWkw9671xYvOjdeGsZSxPrekaKA4DuMCsPJ8d7+IF7wIjEk
xCtOHop8hamZbtSkJtnsGw6NsAxmHurgExhFS472tjE0VJOsbk2H4BkBM4Zu0MtlS18I1X2b/4cL
uH9lQhL2aoSFRD9a9NavbxFxfcxVyzdyYZ8og/wfREiO5EEp0hOLKypbuy3ckIb2bv+A5SIMUyJR
KN5JpvjwA5gX/xrcxk1g2EqU9VD6SouY2m+syIzo6o416tQosAhmx/df5fjbH3Mi8QfU+lLcOZUp
gl01qN+n7krknq7PowT5axuJdR/NF94ddkZLPnxz3zPf7zRr+3U9nGQgoRtOoC37BGQ88P2efewx
5NAj4mbFvJBT2XHILVwVkB3gcIxmQ5+i20GWV+VfGAUjBqOitvXfGFsQVRxhCh/P9B/O+dv2J5uD
b69vhesPFfq4cRkQuJfpy9HsrPyrO2P9LLXmtp8phBzoxzExzUVM/P9r5pYpbiodnyCcE7XafWYd
GJYLjYhLtE1mY8CAK9JNn58pF+k1Hp0KQBMp6ceEkZnSgLtoghC8UGg1hIJRuPlV0Y4CLazh+7LU
+2P70w3tbuJ0xg6hfuu6Wv8HQQwcApxAWs8nXu6W4iNwsB7a0DfBCLyYWaHQ1/MVQ5SXN5Dx3CXE
S+eSDrS64zM1Lq7rK6VcmLh8d8kwqLlV85C5IHFEdnSV67OliOsmDpUquNHln4901JQWrXtMS5IA
TfLDyW4p3jn3bAl8y6T7r+GZVGZ1aUtW6cagsQ26jPktxxV6P5mWRB/r46hdfnlcUqsVi41kdNL7
PdmCZKU10rxn0K7PHyaXUGL/+2cfzpPx+QWl2SAciW3eAlVrqXTdiZUaSbTeuP2DVgSJhJlGptFi
ZmSxJhHwpiqH9B5Oi+7ahnrOFWvlFyudCX16yCSYgnqLyeYF5oOAA1edThZT6zcjVxZMgEBJcbUy
khbPwFWUcOzUkb31F58ToS0UHLrhlEBSfQRNyxZyS83xSbjN4nGeMMCrGWXhD3neYzAqAmRqxkuv
wwYI2whKVBJcFl15b39vsCpgFdyoZoCfepp44pTcoLt1NI+atwNoi+5ZY8BLiPBHhkqc24kRFNnD
P+578Eza6i5nON5OvIXYxhIwmgJXfhmxhQgDIJnu2QdgHrVKQ8Scvbrkj+4YaayCShxkoP2s2/LE
UHXRi4h1RWPvUIjUZXPiC3+KK9yYb6rHHx+uPA/U9Ue0/ME0v5PNm+ag+xHX7N/KoqzJGDvQEIuv
8yC6FWe16sti7wbNwMxRFR3OyHE7kI4bl5wDxOJYALQexpax8HlJc+hyDuW6My7z8sraIdO7B2pZ
3L13PZCKwwbFW9kkaeBAV+tKUTRRKT9ab1EwKfYNBOk2D/Bk+/N8TjfM6joi43X7OWtJy3JoRXA4
tDVfampdZYmuVkET1s7+ciMT4Cbs06QuY4nrvT32Gv/sMA5oS1Bo5OISD7DuUqWIl7WVTrPrWtwz
q4ykexWPkRwR12KzJjM4ga7l4IRiPZaKjfPUtFd/1Rd0xEazJyl8tryLQZWlXBXNmTj5rBjpF6aU
JVeANPMHZ7QYRr3eVsuOYsVxQ7KAJ4tV9svBh2ivpBqHwLWlCwyX9SEk/qPpNW37B+giZkDWkFGK
omhKqwoLHOu1qLXeMqseO1YpXjiYZs88qOTzAc05RCRz8ySoFi7vUTFjMSjIKG2DpatmZVKUVMbv
FKqdSMYVUkceriKO14hvi5LjmAfmtrPOAa14lvh1F/i7vjEzk/PtMiNIyd8QNRhRruatySs931Cv
+scbfjnJO1rdO2Zwnh8yzcqskGsGzsM7nENKt8LPzGJ/dwxOoDoodjOGVKxKjUeRUDYrcdZD9PDT
W9oeOr2axoCJszjaar1ieJ2jXWz4iR+rF6JRHji8H/JY8L3LeIA8IbVhG8RqqIPdZzfyC/5mf1NJ
3/TfudTJQq27qo9n7ZPmEZRdhYmXJ0CcXVXAj4GLSC1oulWWhLKIoIgm3nYbo4J3idaZ2WZ2c/tn
a4CIlHmDq24XViFzOdn8dW5kFoUcqnw99T9HUZ+x+6SRxC6xBRkhxZYjnL6MQu/ea+dYYKmTdvjS
g2XYxQJLCoEHAtl6pj3QPKuOsWhG2G07qMLVT2zZSJHlsoZ7ANxZbZ67ZGJDt1W1AY7FMLu6oAAY
xHwRujBzgTpFrbDVItn3joHdghumq3L+DdrYB0r7raXs059vGUnmVrdb5j1kQAVGx88q6PMXVwRo
tMPeYr/k9oBwoLvU3su/QiTjtoLDFxYte95NUuEFho8RbbE4JOphV8iBwOOSURLibON864c+EOhW
zyl48rBVnbp6QNn6C0BbfXVDGQJYknhM7N3fk00ASbKj4mH1cEZx6fomOMymhebZTZA0hPntac/P
25CWTEfbtK5sYUqIaRMtLG4qgaBpydHBvLNMpPGsyh3FYQz77AZtiWXx1KbIzvUrwD2aiCDVn5FF
H8qdfPBZsZY08n8eiUUJ7Ki9sh296/z3FEQu8EShx/CJG9mrnEGO+IuhuYoh0QFnQrYTtBmHtOKq
IxSWLb1I8ItsszxjZ+MyUP4hWLv79A/AWyCmohciMDikfr4fhXYUfH3fPbVJy27Cm9Z2pqsdl9ra
lij1RG7m7r5L1RGs/ZYhVijgBfX+l++Q2vyPtI5FM8jt7nuQ9BQxgpDZGrQGmsXT8xxO+HybCc6g
0HMuy4L0TBMTrx6tFpzkmqjVAWp7DlYXSm094dBVwHs1eck4yvT7hR0yRkYDa0L6q1Ysf8o5rUXJ
9PPpTal8goP0OW3yooZRTnuOM0X45rzYiKdDYiTUusNoFgmM0dcNhpbCets4X59eEauxQsKk2Y+3
YSkcANNrj8KImEUkSJopyr1QwOCNRR5Qay5MzV2vYzgaORzwVgIjEKakf9K6EdBmH6PG3JxffKCM
/SrV9stx9zo4xrXafrEXiOA57aNelDkqFxLXy99oswNeGIYw41PIERReXJD6Crt1qlf12lhs2B1w
kdEQQ/BnAIMR0aUhushFo7Nl8ME1yXoyuPr/guMR/BTMNTFUbTk9Agj/3dpmhusAHcM3StKv96HQ
JLlcK27YQ3xRRHV9yuYeU8eFDLvv+MM9Oe8h02wI9H1HFYJlILpnoI6c3yK+Y9MpONQDX0ff1Ksp
ZWwww3ExRwt7S2O0hKwadswFw8AygPWKQsGaGtwAlMucbRxNmpP5UugpKDnpznaVIPGlJaYcG1sE
RzCx+6fhIy/wN3Q2q1sgroa59WWBn+tpqL71dhNUCyncdXB4b6bWx+An1f9JUSEJUhv9x6/x6F0c
G3Ml+Mjf+RrZ3H5+rVnZFlHTfiOEUzlpkyuU2YAC61titV4KdkvwymDofgSA9rRGwTSyuX1jpsgO
nNjbm1KPgxFDJ+Bare/Ahj42inqhF2tZw3Glttm+K+vy0eTcXya14ct4RpubTQxCijg4fthyNYw0
dQbQmkQ3MiNA2WFsPzxwlxW7mNJYww4IqPijwJ0wHzexUxctoh5zjlOESPFq7/x94RKN+CaOcmea
n4uzJvthcyH6nAjiWe8tKN7xO5LrgfI4G0izz7LlJ3oVtlz6gNjEsGQ3KFdAhqOcc1Jw41P6O2hO
R7qGpmcks8E57WGdYRm9fJIuUyfGVSOqk6iX62FHg/SsOvNVjr10em6Haw881rF6w39De9PxOCPv
YfG2kBoAqxMcxpPsGN7pkBy0r+LvjmsSCi6Jg1F13QftUmZMCJhliXXUFF5R6eRc7yNgG8eGQDz/
x6R4uzxomNum/0t8T0epDNWAio1m97r0tdwF2noqJby52X7M3j99hjmpjRECf8+XuNdevG2pm6nb
STkPp9FuviGXdTxWkpvsBcYiBVUlIqZFiEBYGFOP81/ZnmvT7od+k6LM0HTk/U+cUcTdKKtWvMV/
zV4qmQOpQzrW0+YmNyThh94Jl63pLewY+YAKjZWCNmsBxkXg9ktUFgNSWmb75TWWRad7lQlXpaJl
aBQYsc0g4UWJiNHedf0YONMrdxgFAgqUXrsSUsdrVRIVNpn+prAc5WEZCiX2Y3cb9OYESVytq0Bb
PVm1FIY/FaPJdHIlg+Ya4YGp6JdxGsxvaE9ozb6GLczyY7GA6rkLyi6g1+m3vWqUEkfTPgGZtNty
m7AiaCG1ySC2ftvjn9Rgmb4ASQRgEIkfDUNnvcswmIkdktSVlnzvH84n0c28PnliqNNCbtwaPf9D
uvKMjaEqzt59p3ZJCSwQHnO6LIW6O/FMmWcDphcKt6Q311WzDD/0Cky7A7bPLY8Zw4nnhgDdyi8l
laO9QB6+RovqN15Y51Gtjf1b9EE8+GH3/OGMM3/jljQd1nO6ZHw3v/5JT7gh0P109iVpRMMUg7G7
SHOEDhoAQ+8ZSMu6ax1yJPte6jNvPB6ZPzfNNyY2D8xCLMLOpXlOo9f47fL8c46/RqYneE6Bsoud
pfLzxKnbnFr6Zzl8ABd+XySxEJXCGJKNRtdvhTUWju4zXfAjH6h86wImcKawaNxiCVDleOsabyGq
0RYbkQn2FkEDopO0KGUomtv5QmwRkr/WlBO49HfdShwI5gRBOUT87UAZNksx2jQT08fVeH56rrNT
VC/k4rlNLtNUZVguSE9E7ZoDT5HU3fAfuSbjIlZ5q3niEYW5UYL7ZAN2IyeB4gqbbendXQjCMnWy
kEqlbCiF4pmZXoZfhnd5gBZDwC5QJIpfZAQGKom1r1BY9bB4gU6boslKz8O+qykKsBKGL/fHjM5L
w4lrV4ewB5E5mDQxBnwHaBa3cf8sQdIai5l/0saDvcVjZGR74p1q2Ej5RAF6FR3QRNV8mGIJ9MGg
oibLrabre5pC3bOTOkNQstQAQcm9MTLH40DHWu9SK7WPKRNAqm7YPfo8k+Y+lQgLCM99qlG8oohc
xUy2DhtQq/CQsBd+hssdYcfIo/6u8XqyOOQ8VMqbmf+C5fzNsep6RD3kOR+KoBiLGVKA4idPRme7
cM2F8U/KYLRPrCIfzSEZP1mIhxO9FLbu9wf+dflPmAgU0pfUmrOsGvTIHcURffAEfKi8pJzYTvID
Tehd6a6/Ii6JizdVwwX/OIoypig4X6Zqmv5rpuSTl0ijJrEtRS6mTo7jpFrtG9yPe2V/j5YsTR8x
Fh87tVU/1npohvzvmQHLp17WGCNzjiemDuTicdkwSMnVJb0vPGGI0p7Q3Uoi0IgHvw+agAeY0Mmj
0t7Z3Q+QneCCIGMSlC5cNENo+NISbV7G85i9xNVmDx1sp7lkJSG70KB4esPQFPwon8nQECYKm/RX
yvezXiLVhOFh55WjUPs0Taaoc1vlSxtIkVAJZ19+rAJwISjMuW4IBmJceOQO5eK1MlBzmk1bOtxJ
ug46bfRttK3OCYRR3MCOMdAggQkF/3WJDRguxwIsIaeUVGcsX+Wubmt2RrYT0HRKt+ZSQH+OdpdD
zvzDZKKWex6stquPHMFr+5YZthrsw5XpjJ5WU3T2sv2OMQZWjA2lX++rXui6UG0nWIkadXDjb2pm
4GNsvbArcWbbGpisMAVJ6bBvhCUtexjO8xkpTj7ye3ItzagfCr1hrgwyryZmAqX8pmvdK/vROfAF
77w1BqqGTO5mwekHiWIF7DrQ4ZIvxsKURZCUpiABvsXyeqYVZAUK2reL6EHIygoEIhOvF4gsBEB/
ZIe+ItL+BK9IvB3bfN41fawgx5uyzskMxbZxfYut9e2ctslS9ByChNXEt291IqweOmDDpXQz/r2B
X1hClFF66yTtZXRYTTRsNEWw5BDufzvoRUyu87yg8ai3+vjpXwXTjcu9owltL88r2NmnJceuJSh2
njaU2qeKGJRP+hlyYbeMGOzVsYZgQaFY8/7lgWE6FVSc+Zv7dvFqQ2UZvwqXZhh318x2osjk2PdD
6syP+JrKBUU4XvncTDRXRge4L+xvxnd7tHE0kqV/DLzMA2ZrozaWEnVCy85NRlR7kEaf0kE0Vbvk
ZtP+4mwAfH8/DX3lEJToAKIjp7uTXH0T4YFoyQVWiM09qkeqq5ok/7lYQwjHAK3Fuzxl2jXSU+Fh
byTPRgwIV0rmoDXgjqfIV+skco48qQn1EtwxMOFTz82biyGFTnsL7SHrhwC5VQzRqEH3XNQ5sR/8
zfexsbIRsqsEl5nQUaA4Ut37s97ZdDZvjxVPV3uYBU3Goh3v7fk5Z569tEQui6DqnvHqfdqYMRzh
/V5UaSE4IIJ4PNl2B0OY1B407fHXc+PkB57SzAWuQXjIaWXiI5xYDxJ62ijL1uGWHNRNhl29gp1k
UdFBhI/hdVHrPvggkk5YL45klOPrwfNxYq/D42CRpYfP2MFXFb1RyXa/cw+WfJ90lpIQrxu8URyS
gmQa/KkZNn3p68bJSz9AqljYHZQ/pDoNAP7eFzEaXpoBs6dWIXw2wptaXXQrHLCnX1MhBMgebvF4
MsoRrnxERt/PvWP/1afjeyz+3tvVBwqxz5WnUH6gkoK9MvNo+R8P8g1BdmtAE2Kvywxerr61Jndz
ApBvh3NxsJP1hyqEvuVOn5z4ts4JiCYj770K4y9J6AdinYi/9+YTqjOOuZtXYJdBbJieXUMiwOfB
hW9jZhrvX9GfpSECjIYCMq7ArmfZMn2xqnYhixN/2f8v6lyA7t3BfTvi8tMLzpKlgrtDwW+Pe7oG
Wp1qtxvnab9NlNuHRXDNh3aUWafRarNdkavRfSM/cANvroYXAxBzSKlDj1O6/aw4/GaTc8zFVHH3
qiXKw3xLJfQ9MLEpNbI0VDNFzLQDffJE5Rrr2XVO0o4lr2ZMKx86kFpER8TtgfaB5Lx6M95t318Y
toFd/2VoHsX4E2fJ0A2Vd+Okg9gU0QKXDd2WLNB2jbUo27v9pAoaecXj9ex/b8xyLo7vg8dLtSqD
8Q/ctxM7BvKDyu05H/03wuk98tssUGV+BpiG3Gdi/9BXTMDmR1AMUBZ1YWLEtLJhOKdZGCOZq/Yj
Ttb5VjNBrTo5zHOUb1lqYIccBzsfLnlwgQbCTxXGAFdDYe5bxs5oQQOHeVUNpuSTJy7ja6Eq//ED
VVXsU64SzMHgaw7KvMNSBIp2cHnc7ffysTZ5ynEbkcb/NP9oL98UC0QqpJWRMzWtwWJeWVft86N2
j7DXZAnw+iI+3ibkRpS3rvlPP8BNgzkEZH84Cs4f9r7y0kLKYIkC6dceVQZ1n8cyrBOKlAU/1DrF
8BWBs7C7spkx2/CAwecKyDBLtOqRM1k0Xb6t4zoc7pm1okSPOC2oOgor6wVh2CJMuhNbfQ25NWDY
G3rHY2eiHa8uRYZukOueo3lpgww8nJ/8llonW+pHYvm+ZwVkZiOBBVW+AnphhYx6I4NWwuLk8Nam
YpPtTHpUFIT8jlullOeTjuU90H8gIO53cNkcoNJy+9d/WKJDqME43sc3HlavoMbqKtU7fDKbqTgc
ZPpKC01VS2hIMVht88y066uVXtCyMIzLVNljL+yocsuXaRENtWkHotxk9tMQ9V24SQriWSi6Hc7Q
Xj46INElSo8qwfUJIo50/PCunLX55hxYFjQKdb2iJl1xDFvecSYyhEW2l4NkWjNotAgldEnghIjH
2s5g5NwWSA8q9HwHNkFNxjf9tmLwfis2j/NwEUiD6Hx4XNVpR5IeLk5ThL2CEFKxpe6e/U6UE3r7
rmajBJc6oyf1zNzm+L9V0Pe+Va1/zVdGAvbJJDZcsqAn/mMe55I/E+7t5WXp0wFjQ0wdrvdRXcNQ
BgvWtdCJNnF4kou4spKlPNnkpOBQ3REP5czp/tjcWqTDsCOQVCT3UtGMAtIu/5XGT0LLeer7j9mG
uPmNBc1y53S9dfaCFa9Yrktq4Q7U+GMSanCfz4PT5ETDhPo1jzvwjZ9w2Gd3ef4kYBPKZdrY2FmY
rYWTmhocHOCaF8/lGED1/vjCKjYC7/cfQFTEdBa+24dRyNKIn68VTMUJVY+zg2z4dZZbR/O/6cbg
wYSE/pWTDK/qzVXxWNhgKtqVHRiwFHBFFaJaTfJD2APZD5uGhPZN3CXumBjZqsVtnpLLJYqHs4Cg
QSaoyqgBMJ84IhCbK9VrK233lzKdI9Cu+FpA7qPOM00nbIUO58emqGIDLx4R/DUdx3ssZQBx1nXq
wqGsY5bwr8AjBcYjvdYjrPphIize1ow9jk9zMlDMeclrjJk929B5p4TMjFXdyux8QAXG6l8nXHZ4
YLtb9jljm43npfScyTGU7EoqjaFTfiwTgLa6zI7kVk9ZGEvE2Dw7XbhtqFR/pHZILXFn0WRVQpgL
h079D1hZ9O9XApRQifvTzPNnv1eCCuCnuPnMgBStRyf6outp8tNmEkGwFvaAs9yOkad01yeGNq+l
ogmmwC1fWTlWCc1oKvFFVDwAjBgP5Jd9OpyTvJT+J/0AtZ3miMFFft2YTOUYLT1RJ78QMfqufweo
DFwuhwG6rYxj5bH+70XQyXmIKaAKenVgUeLloyyBLzdJ8GkV5RIXrnI9dgTy0Jnuql4wf77aUGP2
8bLZOQsgHZ0sekE89BQ3AOIbhBRnQpmaF0WzorHvvTDXG2NcdItIFRLko4I2odKpJ5RdZVwCz+kS
bWfNnI+HthpY6lgSmmz7zhq6R6mdjvERn0SyVuGfqRifzV465+J68UePtKPQTm5TZBwhacfpQs2V
UtXci64FurzDlkE2JAmq6QSxq/wBaVWdjF3jfn9Xxg2pqj5hXij5h8LmfbqqGy1yujVv78L3FwqB
RFBSaBEPOrCmfZ8fQaAFbEE0eFGMLQDK8U4VQX1/hxMjjTUwAlkksiDS4pnxnSJBqL1//hQC9/dZ
uojc7+0/bJ/lTGbJPQIu8eWmI65oyU7/U+YXy2/7juz/DvYY8+xa9QlbjPl5y6peXpqdAYP6uHvF
H+wR20F7CPJe8hmkaS89LQpLu+wGVHplsOSW5Z9QwZXud37jmni0qGbwTeYgV7eT2Ha5a5wznwkk
ycr0o3rKeitCs/4A587iwswaopsLtySVZELfo6uk/QWb/O8bcSQboF1glnq/ix9Ufl3pFkTxTl6d
i9KW37NAEvm0JAlM2/kBvNhi70t+KX2mmq8J+Mo2yX8QvEhqyiUVj59/MUaCn+4vosxxEg1Fhbj+
Lhpck53QFMOMeZEO9Qc3Tiiuv+dLya9HVE7lKauomxbeCSV99GhW7oyybtTKVeKl/IJEYZESAQ3U
AbFkj90vWM4kzdSPuXSFIMNth8V6sq6em4EBrioaBqxIl7nklUVaEYHg8I/t//aRgAe4Bwzn68tn
0ihUyNEKyzr+5BP1hBN/Gvkeg7p0LkLxTc60bKUMuVq3aPzd8ki4pMZR0oW+2ohzF79Qqzgl4GDQ
1NkVFILHc6iCrrQ2AhsvEDmo9mKb7Lrp6bHvToXwBiHF8ThDIGSNVgezaHS+S02X2AYp7pKYPrQ6
x+ycph5xBigUqalebvBWJgWH09qR864CjD5EFmuNcqmE0ctV86DaQHDHZNwTPmHFt6RhuGiOc1dT
cKNLhEmFEqKR7958/HrpebghXmsd6Us0tHYxYbUooz5kFbHmjEkA5Ns6FG9KgQt1tUgJuVhegdxv
0wrkPHEZ0LOKmtKi8KrCsngLhlcD2l0rD4zYis9MIE+rCWm7VDVRapdwDqAOLNA5g1RaveAbK60E
MhuW3uoOkLf4ygHV+wDTJOBQeBprfnjNRLqNBnTDB/LULxlyaxTw1BWsHHhhUXkZkc/5fc99jjoT
MIK88MKmi7pzQDeWct2SxZOks/AjxIubP0ndpkBpIyJWCrbikxanhTUg83HDspGzGtFdb93uuRip
ml9P6EoNviZjMimotMYuoqNw0x8/d8Xtafj3SnDnNJmYcV03hxmjLdD8HjYqJv/0OjlWQfwQKkp1
yetuFtVWDMklaQiDZn0kK0IptcCX8QKSJRy9YqfY/Pc0b7oLzswzGHX21DQ8It7szmNSeGPggk3G
yvGsc3NkWV5aiDnkPCYUZzqFmoPmOZuZDeZPIKwrgXQ7eAsy515WNGsLj4xmHIRMGKJzukOWOwfY
1zrIK2uHbeWGya+3DPZ/813w+G8Hh+Dv+vzXHTrzlOKi7ScHLA6qyfdBlWnLl9wyWiBvTpekaAyh
NWBKz0QR/Rut0aMwnwwoM9+b5Ncui2CCl6SaajrfHVXYQAl7aZsZUHpJ6hfhxoCm24zqVmKc/Hn9
wXjwKKiYa2e2QyIDLwTjD8SXs4DlOTRy3MuBIZvsx7nWTldNauOS0MsF+tk6ELteN9VhE0uqwjXB
qdAZQrIaieN8HGL8fz+Q6TUFlePRBj5nqUSuK31AZa2pSSuEoSvZ/yMDpP0WNdT0tPq5Tr8a80zW
mZJDeTYKWD6YTUcQCwy9FN4n2gd2nCvJPsFA2ZzBa6jef4FiBclj0ktXvN71x4nBet2D/cf8rbOM
l6aqxxcgytT+ZPqPoFa8GUZ7oP3rAPYmNFDjGemMKmNCH8eRNn3S5q03+h4IJi4Nmgv0XEYsyR1t
Dkg+8tQpUVJLjJ19OM57t2lEtGWGkTUplgtnO6XJqHrBwpyafCCiwH+tFUizVAsuStPhcR+vtAr6
0wsTY06LyhyhOQhKewQg4xk93wLZc1Emazc6oi3R3VAEeRrkdzwSAcqTS796E4a3FuShAbQKi8jm
a/+myPH+dndRgs1A9mzJx15yvacjqtUGItAGDqA+iRL6/Ks/OpnHZv0Nd89Wq2gz9PvDqe0DrjA4
c5F0wfIzNUB803JTvETEFUtmkRtglAQKWva+XAL/4rrzhD2kWWtAPiHcoY/SCWXkpSSt4KIV7TTa
ClDicP4OBl9TgOyE5m+qh4HfhZ2dnuEzpqs/pHR5GtnO7Xrs+BNWa+MoMco4H3946NBpsupaVBMT
UuFjwqkS4gwt73MqUC8dUNXwaDOMrz7iFD8dbSWHERu292kigN3EBM0EzaNqGFCuOuhyj0IiHJHj
uM5frb3K0T0vS/Ad4Nnr85HAlnn0d9GDdm1EGDA+ac0eIMiwzuntv2YxkzY67MzSOCL2cvnf2nyU
EZkOgvkjrvAPq6yYG5yb+tI7snFRYu50l/qqHklGfqZ4dSE8qHH3jyF6TS4hf0pWI5aW0pBtYpH7
rUStvbSwK1eG2bBQW4opd9ihQD0ZKYFlJKiGoa2nbxayCw12fUqtmnK/Pv72jM6z4hByJHIcJU67
D8/DWW2R2K2hZzq34KgVBMENAj41toMHNfNjdJW+CBc2nhngB4qSOOOcgxKop51SvRcKn+2J4QST
1uE3Tu3whbwYTbjjQ2xsT4HQhjPS6Nu27Npgrg/h0IeSctTLTR1w+SoFqfvGTEklX7B6W9NozDNm
dmQsT5wmfjh9zZkpYMICg2BOaUVu/Acp/PVl+P9Gq96L1WHRBLL/QWowvJR9g11V8aydojXnm3As
tOVwt/cRU6LUFX2krCeC0mobbggcaR7ZBQNYTPA+C1dFTq/skCPjK7k8mDXT5IlV1LXb93+5NuxW
Pwsq7CTdvWACumYg7E03n1wT4MyWxmMMqtielHBqB2Oikp+LrylzGDWVricbFA2UpzjWJj30IcCb
U/w5p/yhPwq5QUf84+6U+t/Ma36t7AUdLgoejVpV81jW3hHmj0R/jtWmYEOlNGM17fXIoqiUeY/H
j6AS6dUnzOS8YDnAD+KETA+X9IyjswWrsX0eLUZsg+txazhCC+l/ueA/9xEFb/UW175Pney24xxL
RZXE5Dm6EkOIVwlKdGR917x6KevLbAKot00Xcv3qKmSmXHwTuhjt+BEoyiRppA1iu7HUd9yKaiLw
J/fCUZAyLV88tlL/82VQlAw3CLc+ZzTZPEcpWFl8879f1RlfyvuCPPTQbYwTmh0HIxT8qNz1D+jj
BWq3zGhyTZb3qAP6a9chx7OxLk90KQlIL3mu5kKN7lSMe9YraV4heYFkN3dMuptbABXzuiaxV3xb
DmpXCFOfwmoqmmzZ8QIfH6Q1l95ci7bw0CCmGHeWvkPSGgdtypgl/pxyclYzswISV7oaq/SczHK8
ZbwQWKb7nydKwscjk6zykCGrzpbE0BgH65sL4AxZrOU+q+nMzVEUZ0KLWFpLY3UQzzMVDOfq/7sw
16SS1REJkSJXRQ655h0ZPe2fIrKZGmqIwBnHSzw+TVsPCh+N0gpD0NH7HorjLiiWjRV/sXYrEV1L
URzLAT+kcTEPJd7oKs97ryRGPiKxC5T2t1el0QgxRJlKIP/uHZJZRx0BwTNzkzH249vSP1MqaZdT
S11nDOtODih1QlOAba6wb8dt53GwZEw5BhqPh9sGgWCf23VOcPTOsmflCNehTDlNV9P9l0vauMQ1
R/F/m1j3DpQnD7NTNW1usdneHzPgcGj7BeUmKHj8R2uouqu48+pT6Uwo4l42BYG4LFQ1/WuTTUAL
6wdbkWdETJ+r69u63MBwozQ18wEeiuCCW2nBq5otESDS/6XotW4Yi6GdAYQ/8IcO1zyrxaacRWCB
aaEtf5yZ7ti+A8Twqv/s4mBYlDVa5CkyaYiZci+qUBHfpNH6E8f2BuZuAWiocmWqjD4ljYFevU6R
NgCkPIQRFpbQ1/2HWfgY//0y6bD0XanlodNSezVYeu4Pv99PuBpjVrA+EqiFOECzhgrCXPKKvM7E
5raW8D5zSR06wankQTmVt2nqd0euFfxU8IE36wL/5shubxw74LNG7Rft/tfGivjhG0gVEzJFhXOY
IIJIoystb1MvrWuKKM0MrRk79K39cS/mHaSihbGvv3vYPnCmn/1/nK8uEAbOel5yjIWjP/tsgSg9
74I7sAvM7ChJTlVxOrA7g+AP5QqaYEdObLmIsRyXMWswQBkRYyzXJ0XFRfIwPvp5BbuJ1JtDOTlb
qPY78sB25S0742b4BtSG6EIlL0MxiEGwPuti0KzIExC8hQoM10MSXJnmFG4agrcqS2Mwm5xD6FXU
FQtAZeKjmw2+WdtdLtzhkIFIWp6f/vCu51IbctgzUW6/xtkpIg6sonMPS5A2GFvcP9Ub9E/6zWQg
kFihSrUqp1b1zsUJ9W1a2CIvPcC1mnOoZuaGl6YDDEvGMaSYioEJBkVg22N1dVIjlR47Fbjo6MXX
bdDsnXvwGA9ipQjWwWIVcrEc/odo2SQKSZHK6bL72g1s2vcCFzb22PjITYxkEP5VUXyHyusjzWPH
A+wIKX2JhrjEXYnrrDnxikfxWxem+QzspgCOmoQG+eL8SGc+j3oTUomKFqFnGf4MIM/LY67LOyfZ
ExzxL5V3v1+Btv6BJcjaLNDVgz4hC81Zl5f2956lLjYzYvzj9LtOCPrjIMSSa0RfDZt6SqxdqCTu
uk1Tn+rgLW4aDQ/CzYHcaI0BzB44ZLYTAf4aQPhKfsmyyNgvhxr2D5IlC2vodNG0Fi0ZPYC6b1Yd
mj51WsieLWWKmUPWiUnFoSgn0pjBpB1zjNuPIFddLG2PutdH4T/5boqmknDFspjwN1ePKEKCO/Iv
nTFEBD5JqEowvQ3ClKRyX4ZErFY1bG0vXYnxktO5ccSkjan1ChfnZX2t+FmbOZozTRHSG9NPHYVC
FwmhjZWXqf1lrIVMM5mdf7y0E+tcb7sRcXOXwA6gqA9Nl5Xm8O0VSLeQv2WyN09hyxeSpQNDVJ1L
GsqIcYImMSC2EbiGATm8pEwPL/Ict4h35mtxt8AG2aQABmffaVLF4EUQzSI3TlN99OTiFWGWoBdl
PLdxOTJa/ei25v+I66L4cOW034At6jY9z0Lq/AnY9+LGYdvqNXdsVzD0F3YhfSz3lokXEX5wJhYz
BbVV4PXYdJ58xD3fsu2Gzow5CRIt59fcc05nPXeH/C3qWLbhEOdvORiWFpQRN/0D5ZrkrpmK4/NS
hOz1uJt9Vxvd9gLetxukVvOjVcQoYbSRX8Qzf25gqC/r1wo8qAhGr+TlliZGQtjMmxtdt4FaSogH
hRnUIYYKcBXD3ubS6s8Z/b/kkpCb0dHoeCdc5ZgGJVrU7SNJ9wg7005XctP/fLJ+5Vj76FNKgq2k
2Yg9GrebIu26JAbzFJ/BCQYv4vlIc9EtL4jDxlRcrag5qoVtD/OrjZMFY2sVwfKXg+v8SRMuNANV
r8Ujg0cnIawuP3X5FZz9HbdzHmz5QrEtpQsxE+oYA2mdNzeeIaEKMOJf1K70XNpl8FP+y44Gx11Y
Rv8UvZwqk7tmZd28+y9YFojgU6Fr65sCCrsal9dsSKt9beYgd4ubE8vgM/ianlFRLDWFOKe1D46S
VcOnATtV7yL7EVJ4SMwhA1JawhKUfCXETQV6klej8Ujd24hnKsIpyl4bhjnEMA6fHUGbUsHu3Gvy
rnVNxz+1hC2lcj9gUhfT5wno9Y0mdKYczG3oVbjKqNc9LuHS6dEDJvs/Kd4Ukn1J6H4/cL2VfDjA
JvgYckUfw59ZDnsAETWrMARoW3rziaBeHHJGX87cUYzwVn1Xkik2QUKkLgBngBhLZWL2Ss4ljgJ5
m3f3n1RcizI2Lds1Y2PcKVb2PKmkLY/Z3Z07iWD1anBQtgILUX8Npr0auFDeeUhAMhOf9I0c/Cj9
LvaQ5rxqrRzwMMkpYgCef6QGg+ikXpafuJAfo87HeGjiT6zmUDFUeggU1YDR9TzNHaGslZ60QZC7
jTheaqnTEVkMO+Q9vQPK9Mu+lidKn7fJsBIRnfRuuASDLI9XsDCNOhXEBMR41EjPuLW023uHRbHR
nxM4Foty2nWyf6bfhVegrgAZLfeaqSqCyiUFXQveuNiyCcxGhj7QX1+Hgdkncp8dQw3dBAoi9ycX
X0qMXNeMZjnFRK9SngU+Ba99tZtDNRU29Gl6jNvXNI0N0tUOpsYYFUNl8J1Ar7oRZM5K/4mi4/BS
HB6wnajAy6NWqZUklefLF8zNXDYpl0folDQ39RNQuFuiMBDt44WvWfbJLqW6GMyqajc7Ujky7Wvl
53DRbKe1VW1wFx5kMeyR4ktkgFgqhgLH4eCWRHq9fa71xQcLBNKcRfWKSKE5ARfLuG45tDjsGlRl
foGOb18gGMuEf2RFCFPGctT9gyt6czK/gx9YjeDVuQExTEG6tZ+5Dsu8xGgunzdOk+wkc94T99Jw
MYEAVcUOcQxRI3frEsQhEpRcTdJCeLoIu+rqVEaNQJUw1msuSeHT+0DAxTNRiP/D0OIf5TdYSjnY
Wsb8cgltY7tBR4x2moBlXD8sfo85Xww140drwpZXLhYiyuFplS8r2lDD7bDOyolOH4mnvzqil0II
lRA6CZZOG+hukD+v7Cai9cppmTsTWi2GtkBy3nFG6BN6SDhQ7PBqPopOInysghlTDVsDV/8JM1R5
PIK1SrDmO+rujBawfr2bdEiwEe/46b6pwC718rHjr+6hkxSsaowJXx8DTtGvzZVdeKBFIkE3VPzX
FlMvIkjBSLoHOWlD1TDpjTJ4vpMq5gUcL+pm8yDaxA16Ad906/2hntfnNdfitbbBC1thTthTGxmi
JOQxcf0pSoKuqc/MWVjw194NqutcD+YAry1T/IQOCMNaziCRNd17jGI3NfFEGYyIi67Mb8c2lq6v
T96nvr4cFA1ZFMfnkKS7fT6RLcwOGq957THtSYLczgo2GFqV09jlhkx2wWcUDEzrPaZb094I862T
/JQmZnnfaC5XBkENKoeGw6a2cpMYZuZHnrXKzqTxmK+MPAXMxrr7fasuL0jK+3TO4nNrbdmJKTHM
MagBrFRdDHrE2x6NQ/EGpbhPtaFS5cQB+QU+dNEwHq84Mqk/0NmNhFcOc2svIeC7WBNxyvRx8ct6
VOOvP8pQTCpAwunZdTenl4WSS1rcVjujLgbr96wrR+qj1U2lbhZX17Z2qG2oI/fAmyJSNw3dgKNt
Wal85faY+BZWDMsGQ+bDhyHSXoq/bm7LHwF1LZEoksk4Iuus4uoIS4oRl/0sY0OG3SDckmkSnZXT
soTDjsgyd33KJN1ghzgfRtgqM2u7hJwb52V0zHDkj8nNIS5rS8ujCbOUVn+/DVHVMQd7GMDeDNvI
e3013Bs+wlzJqcfARJ9OMnzxaKWPuDpf0Bit1tuijkFWlXG57D5xq1P7mH9CROi3SeUoE4h4+bH6
FQKcbv2WQIoPwxBZNBPb9vbSkd7mMBAx9rP9vtzEapZ182+NZlyAUTsNBlUSxcha4hozkTTldmLv
BGp6LeXTaLAxoT6fWVdqqx2tnfRzGTbtyzDg3aDaILoyQnxzHt6sndsU/6jSXUoYrog5WrLj5OL+
sgE1eWki993/oaKvKAeYo52amtKNSmA39OPrH78FzbKyoNqRQCTBtJtSnWbP+/RjdqGlbQL1pqhI
m/lh3tXJSbf8nVZBTktuqAmGC4MPBiYSku6KJa9IvLJ3OY71BS/21vJy87Z03uQ+8+V76tpbCHiF
gJsskrbsRZH8+7Ep5tQrifjA+FKaMkpBwzTCkU4X5DsLrQdQKKEKTS7VFvs/KlrCfL6qILT5T0ou
wSMgOYPOxmOIZFeg+NUmQ4O/zQJ3dEaMo2hl4W1of1yRV9m3C/Gxr7JiJC3PDv2I6cJgEoTMngcQ
8fefWV07/7ZDZBzWq0q0FFA+sH2SChGzlO0m5wvm2SKdE3/oEPoIgjJvYkR4apQkmr9jqacCGGo6
PEUtTUGIPRXKQtrSMwDyjV5NXgxz2h2XmjAdVmWoFVCSPmohsbv2M2K9dHSAdfvMYii0lqiGBZ98
6hhwYCkY/gpgjJ4HH+OczhftwxlIDBlqqOxOcGdEfGEvPHZoolBvZYRKRWYNnbqc06vpcrOc6g7b
AO8zB4HQvhpLQsdqmCqg7GjRKPfKNl+KBZbOGrV6eVTr9fLAcRRYtD5SvD2I4rhMVSTtGM9IZRSe
EuS9U2aS5qzTdBiaGup0MPMciEOgx/CH95bF/SMHIjJRfGhrmtAlkMjkwiSGykLiW7gj2qwla0jf
M9iCeKbDDKqsgtQQDnzrByYG8y3cLhfJ6LHvDcseN5UDT7ryqK7Tqa3MEalpBzseu5+nE5aoIMoQ
f4gB8X7Pzw3snT1790g1qcLIJzzQU6xtpRPfntpKCiCIGvjAC92wDGmM2WgHyVDw8C9eCaZqQR3G
9qHyGb09QuVtFKXTh+rCA1gPajeX0Wjs+lAUnZ3m4NeFodj8YZyCx3cbzFgfq7uhdeYZvuAtlnqz
pcrAAqyfkeXVf3ev01pyAYKp/POg8KPXf1Q4qT9qVDJAdMbVHYTBZ5d53DSPE0b5+w7C8TjWwCZX
BJLA4y0TPBiRG5T+puy0hoVR7KZSVQo24Kp5MOyZe0gVPB8lna0i9aDrG6cBtE2yBKDEp7IgOeMO
lfGHKg3AT6sS6SDyXVcOlXt/qiTSFk6e9hvTC44vunxxKc2KREhp3reE+su4EwAoamZLM1y/fmzj
al6wH++wert0Asgpd1lgG0F9xrO2lW3mxeVidSs5deJJp9sL2+iqp3nWMQ26fNTu5vNN5I40fZuo
j5K1unI+2vQGPZw94u2Uk6Bq8cZJ65mz6vk0+k1POmxC39UvIVB2BhEePOREB4ybvfEiWNydbPpz
0oowLL7H3n8UhKatJVC+vqpmU1ADVmaRAU/KtQTmz1KJehyhz1fD46ivS7IPDIxGVlJxAmknS9LC
Hfbmup5QDKrLmCNuUpmBzLFxQlLBwT+gE7TM+eaOQFacszNAMeRcK1UYirbTgGfZ3V4+qc1r/NrV
+eyrGMxqFiK8S8osRbG3SmzJPrtXA1LKtNHiufJjSEhpuMYS1Px8OGAQIzp0Oqu9EO9ZwR6dcaHh
TpOGg49KwusMk8bK12YFafyHduhO8wn48CwQwA1UpH1T6UumDJjzBgYs50FBsDJgXRRRCr4ukEmI
TXSTw8u5cG6ErthqfZCbJ6B3gggL2mUWYHpOfwy+iyzwZOtVVfbjydL9gV1MFiVAF+/24L0iCzqK
iWd0QVNPMfczVZGfvgUJTZwPr8KgG3u+Vnsm4rmRfZ/FJQYt432b6ghjeFKU1ATIBC9ugYm/HXQ9
P7f5ymHRie6ljuWVEhuGQrWYEAi4pcTqvudPPQkdFbLhOMCQRWEFM9W9Ncwf9IRHOq30Z9So264J
ZNrTsZ0nzcweFAzQ2CCGwheiRJVX33G6cffjZUiWdud7syO//dxxgsel4rsz5OVDyiQEq6KykIGg
9bVcvqOf4ahxC/zctAORSC6wtw8yFQBadyon6a1Vz0rxpqSPNXCnKDJsEa8S8zn48KnB+c1s0fgb
FH+HY6UFyNQUxYdWaDB8UDEXkU3JWJoFYwaT+5t0Ihuy26rdr5/1o2FKThafk7FmVrxUQ5eJE6E/
A5JGK3pLwDdUylNiIvn2JnKiv3dyh49sl07SkTd8KyMkraEUwOIsIe24QqPXStlmj/AuXbafhZll
emQU2NVCa8j1fnzvQK1zsqbpnsObQytsJMFphzmHcpLtz9bghTcLZVIy1mI1A01tGfIKLFH0lAhO
xe+++x50wrJDhMLPYHabBqakpkz5xWMBQlQXWq4RccYEUsCvhtirmXcRn5TpYVJGLXG+byn6zjQn
JhKAKxXS9cT8MWEScshraLMk+Cy90kAZ6Ak8feqrCPLEDY48ggQ6fwM9Ku4dFrSQfVRF2LXCem/h
nHxnjwaxfnsC6/ah006T158VvI2pm5lwgw0CblLP1PMXMePBTX0IegvXqEC4CSL9exl+nSJntsKr
E5i3Gz9mqYTfC+2GbutWb7SttPppycvl1zJc+k2JcfB46Nmen/oW8ld/WCzIwmvAqlhCw/x/JP01
eCCLatknqZnmozT4InVisgP9PdI/R/kFdtMg2mNRCqBirxkgLcWyuGHTacTe5+mGuZ5U4/TnLn4h
tPTsdYCwokd+iavTb9KajJJSTc8eO34DZUszX1b8oKgLTgUkb1FBsd6WoNvPyt5w9vKTKheAmG9N
dQq54LeEfqMOszgzJIXjtwRfUItE42gBGgbGXJPn0KQoRZdOZ1rScre0VDqI8l/jPktVawSzIcGP
Q/p+XcU7h0XzxnOWQstRUrYVhZjTQGjOuo5JdbB1fB8SJVJMDM7KhuWZB1SUIMI5l3GGk9Iao4E8
89JAL1ngWSCVRA0DBwXchmaRwk15OMAiiTtdjVLoxMW7dOROPACx8VgdFEjrPlaSnujTtzm46Suu
p4hAKqfD3SGOXFee0l+4jq+yspj88h9pPoZZv8Ko3agZNE1WXLOMWsDOe6SxWWVfU+EewNKAQXx5
uqf0yMxYkyN1Wp181J0kwMgIXr3QwK7QHlamI2lss8O5Z33kH/5e6hvTcmu8DOUUTwBhPlXutvPc
6XiKAuI9Wel376G8r1WeZUICOefzJN9DO0TJBZKHZ6dCNACX/NsGS96irrIIhnm89aLOY8JyEKYc
q7RxxBTc3hvxqc/pqSCUt7jWDAs+Mc1tmgROu3jwGGsM11z/G6GhipcElDHOlsHzIZmAoGip6Q2u
YpZXmxzruEyAYn+I7MwFXKTg4oQ9jZrOAnad2snAKZIJSt5bI30df02BeKZYx79oBMpdcY760EwX
vewSTx5boitoCxxlg683lLqR2GQzp1dLEDvr68BBVbh+uqYt3FX9oEdOE+qqMVz1x9xB5fQ7eUgG
Sm+RnLs47CLJE+rqOeTQqe7xMIwz84TaTuryNB8x5Uu8U+3mcb47wglAabFkP4cM4PjvsbCa7Fm1
HxThjC4YgEqfRFQdIqFYgRApIYpphkm22SLnwQIjVdGGJkudNTS+leplx+Nsj8r1TifFtAaid8Vt
Qx2n6QhqSWGdZe/6rvrqj3GArYiidxJZYBt3Aus5LhK0UgWQuqDcBu9iLjMCfp8rhwrZriywn3wS
5wfG+BO+b4YDsj/KffnWBv1PJtsQNvYtn32TF155HL1kRB2BnSJL2MXZckJd6ec6S3o5yj9jp90N
ltJkjn3QEHqGfN9C+NDnx1POLN2aMFz+9OcdoQ5GGksX11+ekMJauUpzl1LhF9FtvR6hVg8ANaEf
7wOXkSEjb2Ehknbk2aGwBFBCDTWmRUWEzN1+AfRt1bbhPMJTLc2g+d8VflyCGkVpqJwp3UxU++N5
rw74kcJjoCE7xEZVeJtwZo22OUP03EAu68lS6X3LI8dIJJwWWDDt754wEk+0GpTOiACKDabuUBYm
6xsaGEUMo/dDpfWVtAjDEy0h1Uf/SGnDe9E2C+kCAuUFaZ454Kd8o7OEzsdLH0r41IMZmkI2MC52
S4BCEaP0RxUn7HVXqpGclgrMYAMu3h2JcUpCTvqjoYUmli6MzeEP7HSzzyvMJBBOJsbjYdtain1a
IBHMtlkOnu+GAGxPXAUF/U9RxvFxZaC5NlVlsIEvqNq+MmqI16EhEKbIBoz0hZK4JR4HaYtklimL
w0H15xw9/g3arPADiA6V6xn1/p2T5/8b4QiUg/asPZfgonoSIgFT5HRn7kgjZMzLJklkA/kTr8WW
8eGVgsPw1DJO/Y2D5Pbgs5FVgbZu9FOw/FPxqpIi+WdmxotgotulKZPTYAgYXG98gA/xnbtaB+IJ
0oKghpKBS2sL/kH/aImK2S7rfeo8hIOMG4P7l4HxoKcJoLhq1vLXbip92lbSvQK2C5yma8gbre01
41Gd2QT5huPCptPwmKB8yLyFPW4ZTuN4DOV6f5lupU01iOGJaZW6Em290JyVmkV374Jact8JlgTh
xtlCNyafrvK/IZ6CDtloF1dHCeT2ERi9Xr2Fz5nxMS8p51ho6DfdEyF1SvNBOAhEJ6wPYsej8zQE
vy+zmefIgDjzCLxm8wew4LJxg+DJdVAJ6ZQPYVAxjtgZwoRQLRMk/bE1yuS67Mb1AIWua0ZMIguc
oq7P/yyOsgf2BnsPNLLe/OE55QGhEVU2nubXULmELcxsPRg/cJZRNP+hJDL/yGJxP6xFT4wOam6l
AT++w6aIdpq342CoTU3qNO9daJUALJOSvwsk8iFubjUbOHKbdMeC/nUUixkB18AcV+awp3jCS9Vt
92St9VIB7EQN7RC6qb95WoQ1IJUV3iI5sKIPepAwFG9yXKu4IG5d6a5BmqmreMyMcqO/Tw9NtxCa
RMQXeH7CODZt3J5auPKJkoL49DWknZtZ/K3iJGv/z8FUfkihk2HtTv32QaG2CQr63FZ76PfrpHSM
kxWL8aHFGBOzj4IRIwiihbWsIiDTrzqMj+K5c449mGcQB6fiVwqjEE7sCWL0Rm+Px+dvzKZD4BLK
zLpUk0NCxf63FDwK+Y4qKdBfrSzZVsg1GKcJ0vnZ2PAJJR+xyAkgjQkvuO1p6uKemSWRdgzRNn3m
N2QuMETL3NoWyzyL9Ys1AALTPIZp0IUzRkJtlkIp6i/xgZBxUyqnu3ZUnoqacP0Jm48ub5J342Rs
48drkTaAUWAwhY+rSWXwjbcfP3SO1mUeAzzWUvCIt0s1gbN6DvAOh55g0zVel4/Om3UOkUET9ma6
sm3iKQ/Pl7kbbTn0u7mvbDmgZPLQ5haJVR0ELuY35cztHlRBjcKyio4byKjUYFy/foOLWxdBB17J
yg02m09CK7tS3K1ujMcSdDWssqQ+AVY7iqJ7WU2HqQppH0lPLuo4RUPKbQbICa5ZwPneISS1MhQU
QCIGvvqmb0SXz4dxbfeJbNZRCTZ2taCHyU9piWWcnWrBlc1b6JIe5LzQNR2SIzsXRKxe9hT04EBI
3si6kvfVJCjIk+QaTXkvCizkEZBk0zMYggZ/oRbQn5KK2pHChQR2y9ng/yXOvITDQGNOh838U/K0
8RVHH46F94d6I2w7JOcuK6LpuoK+u0anru2QJlnWg2+UBHYnl0NqXYAXeUiUsrCgpawTWGT7KSbV
HJ4rj9TWzWrhWjSDV3MSdcQ1tEhz7llq1Ri5tdJxotvuwmPEVwHdkFNlnK0QryiApAxpSwxY9FL4
9sEg8Pz6pWu40zUUjC4k2bGYN9GrKXe7gGfkb/OoY6Twx9fM1ts4sBmO5xu5lbPSlDwPzr6fUJe+
tK8vgfKAYwdlcOSHghj6uzWD7F2KhyQrFK7Evv31FXl4PyxNKukIM1CqyRRykSUoPigLlDBc/MzP
pjzanI/8RiLtbGNex22klsFlwYFbWw6O84GRPDuCJitDG9S5xOj3cn+1Al/yeUGE0UArcghBsB7G
jQ/SOy90/vKOBgV9Sdgpv+wqtm4AKqdkolu74m4ENpa3ghWf7cJZcKCsSFXtYWOK9fMRIw3EUmSE
5h+KQxO0yufmSXmam8iYJwTeUr1fZXo7NIoyveoKBMkbYBFrbqf9p0LfKnFS3QFxktAceRPAUtkQ
V2cb5jYVVRkNUEud9SEk/BYyciBs7d1qKfYxcb+Wkz1Cy21w8hFVp1FAkBHZpbN6HznB1PdYDvNH
ZZIMc1/wD4uY+ZKB/eEPrH4SJUaDI+axG4lLIrmNgEbanC+LqCVaxkxC3oRhxLQ3oUm1MSzYW8dG
1XWX9fIFKLX283pwdQHRSLnHJUcsNLmDHh3ZN/btoHFrmYsOU21EB/MA9p9VDH+xmTG3ONGZRevM
kx+tBunK6WkeNcAX+QRdfsSlX2nehb6eteIAOh+a6fk5aSQYUmyoItOS5JjHjKqdScRDrRVOxsxm
iAjzYI4pYcGPt2jT+YvsBbFa/j0Y3PoH3IcFOO4iTbHAq40mM2HQgno+U7YUziYX+ijtrTf17Cvs
ZEckbsFhP1jzpo58bo6Dxe3m+pQV/3DlPxtFRplwkXOA9FQYJp+6EswrqQQyzT/SEl6YUlEQ3gq2
b/VmXHBsut44ziEf6SRpz0XIhQmS/51h1KfexiuvBCOHI8oulJ2Q2rCNxrWcjM5zuEq9Iy2rdVPo
HNDP/D3CUlvqDs0lXE2xwcHf6JF0oS4SUuLpfWKgHdWuRhR7T3jAzm1R+E/keB/FDlXgevuRTkod
a+GQRz6UIAqZcJlfuUqml92d/as4qUTvGJMfk9Llv6GysUuiZzVq99jpifHyv8fcpgG/mlvi++Y6
M68FGBNUkT63ofngjIROv8E5GYzUmiahX4qu/0iNzA9pOI+XlTHl3M2M9nDUvRq4inm969DcOW4U
31kxF+is47hv68V22J9L7/bEfogIJGnwB7r0i9H4kEXPX6/GuQim4jas7yCqL/sH23R6il/fK2j+
CNN6INfwa8E4Ft2YEFXxIBkcVe+Enp6usmp1YLLS+zwY+D3AY9UhwOGmB1J9G3Xt97PT8ZUM6FsM
iPtH1ZrWjKZeWv1Mvxap2gucrBkSGuvncY3kMG+OkMJG0wwBCWdwJIcwa3CIfFSxS3XDe2wOX6ph
Ir1afwMrnaHWb35dB3CPbW0v6dxVi60258avYPpnjA65uugaLQwj4pwj4jB7HBFOUCXkvrJ6+udo
ZH+5DmkDWChpGzrvHB4+PRWEmp+W3iUPub17Z8yFPHUyYNlg+5FHni+W//66r4SzNcSlnU0dz5a0
bGEA/VGNQBZ8xMqgHWXRrgoAPSrxSz3/NLPXFUZgphlTmI5rkcr9t27DEP6kfYN+9je2yGxjeEMw
coFlrCGxOB4ZL2PQSo6tLuiO+w+qrdMIf63f577NfwFgbhqtTHmjMw8iuc5MBiOW/rbT0QOTcnBH
6Zk6IC9brYT6ZX7NkTKQ9Yr2lZGQQfV2ZA9RNqd7pHOq+lpiRQ9n2wPoFTI53zSohaNZ07G40RqE
q3DEEDZ+Xzx2JZ4iJn5xX1FwIfpgRyEJu8V+nWCAL1l9IBlrgCKj0qaBHM0FH4ZhearZxsutXZXc
Phg5++9ThZr/F4kyKQuTjIiUwwszZov/VBtK9LN2CSLhJJRNF3dyHkyOnJuts/ZKiyA0DV85Eb2/
mJEQ7vzpXC6sR6sfF6POi7iazB8/YvKC5+JJ2S2Y836f2u9fuzg8CWpncYye8RbG4bd5aob/DNN7
9ZGsnVxEXb738tC0r47NU/h9a8OL2uVG8NuerYoUBBsAPFYDAi2xU4rpl3D+B/L51OjY/dFxfoWo
l6kveE3xUx0iEOEk3zy6W1M3Fy7KRNELxtnsJ0ycCnn7rDmV1EzzCSCCMRWXlec8S7BuCDWf4UoN
6Hrwwxt30ScMmZB1lilPGFfAaPuEafya4dIhePZz1wNHyLOL4GQRitj1W7seAorFQKl8JDc1UWGn
TZUbc9ZsYCw7I/whKJS510dtkxMnRm5z0eoaZv7b9Mqfm+HU/3aI1GRVw/WC19eQ0cKjwi3cfTbj
umKpaTJEb+c5h5FSe6ZnwctpzccwYxHnDAegus59DuCfpJXJWltwIA/vTNq6KXpwJ5EtNbY5GaOF
g54rhg+WPYAFI5OkfyXBANLwgwPPcdyrCy2lOpkcqtfLZ3Ez/wQaDywgjoIhSw0AX5oDyiIFCK+V
jkk8p/3p7NKXVGXE2cP1dOnwJdaVJva6Z5S71BMZK/MQvbKeXd1GBLtiHA/rYCvNY2sxjGBaPXgN
UywNf7SDKM1rLTAXcLuWwK0SLP0Mu9eiyvU0lAlF99M5/Z4yiSaQCJY1ylBd8AQadjUEDWp27Y6q
uVgGQbfGmZFd5Ho2ztsOpWk24/u0Zh56kKXUI7RKJAkISoY8P76XG6LTgFUu7Zwmi16nxtWpxCR3
XQqJeKhcaPGLsGhoeIrqkquTewdxTyxEG0/DPuRHwK6qQyU0mqZpSg+S+GXKAHJT05d668RCkgfV
O/vlP5wP1Sqtfxr0Qa+r+dNUZy5fpBXmauZTQklBDrp7S2e0qwZGYz9Gzk+MjQ6m+deEEFIMjRM5
Jx2l4/+l6dqajrHggw88sHTQXBVzja8pT+HVPvrrDORRy1Y+n+nHBT0HICNgdJkKWQQO/dbUvD//
o7rjugXioorOcuYph1u6rOS29WDWTfTSpmtBeQW1C/oic2S5QOTM8p27sBD40tFFzv8etD0bXJ2i
nefl1+K5jQjozKrBmzDz7Qjj7P8ZvTKKUdJHjSEbTk3WoQSGz+xjy+F0z3vbDQZ4kmQzYMBqlPTk
/6ylUvoqTmHDlRwJ7jGijU8RdkGxLZ3m8K0xmG9b5rZNBANuCCsgcycQujdqtbilC1SxRrmIzZuN
1k63ccuXBlLhgtz8RwMaowv8/70ltrfhJlQpa9clDmNzBe2HLs0I5ZOluM/zInO7NtEG0r2g6eRn
OwHJOYVYWgv/mTVXfTAep1U5V1euKD4UFrWLc9HOdsWE5Oxlcz257x3PAzAwuOneI3dNYL6xZ6US
TCOlbJaLmnsIIvnaph5Hv5qiD+9pGYCPAVa4DudzNClmILKdCQmLyXN8eyHkVJlv+m1G7AflBwHQ
veemQwgUqUL//xTQMljI01WBGTXI2QhW0SpZnsyaZjkvw+4F5/jwfQY5dIM9oWjmIpOgR+lUNgau
7qGDJxO/V+MTjJOULK5wkXcNEUFz2mfeqcdfjZUtbz69sYuC98af21ViQA6CVsp8wqqTp7tgoLYY
9oTN3zEG5fDoYIsdUpy5X1FUX29astHxTTUdg+LyrcvKMGP3a4XXxvD3lRrIt/TXE8oH0wwEpBGf
mvw57AA6BdzHUii0suAcpl9V/z5YtxcuwxdV7nODlzA/afaCrvxFKXjFCLXhDfWiGSv6PXKSwNyh
THVfDiYA6mJbM5EE6fO/NZLQG/gKVZ87VMEpMLyxcd0eRoNY5u1r/VUuXMzHbEDwLdTXsqylLcqR
sPrdUnK8ErnmNhqLmfFDAX0Ac/HhUVZhphTflR0IQpa2oNF4PXcsbNJPd5FAbiwANc/OpwExRpID
hmO6REApXkLtxXM7wGF1PRhclVpplNMob/vc/QdaZtSQtjMOcX36hSnVzf4APu9A3oXWhV/DpmxX
QcVhNpuPfaLNaPFIoMLhWxKSuxt6L/T2NiXPkT8spxQ0jF0gG44zyy7yhAhBaKrcEKMOnmkzuieW
0EhNBq06Uo+9h4ZGVr/0ZG/krZDeHqu4dUxUm+Wgj9zFzLkusRZBZ8ey8DjGsT3dfa83pzNjy4uO
zT2Tr5pTy60KcJ+JsmAYmLKZwXMEQCm+UdcM+D4kpD6D6KBtEikG9fosbXvLYb/xt13h0+GFFg77
+DHDjKXdYmJlrkWCt3h+Dav2/xKqk9MQoDfAUDMmbRMQYK2rfbfEZ2tyYh2+AeTdZW9nNCRsmUvN
lxshS7tHVTRDtMKp/c9SbAgCb1/KyUdXlUpqK3pd6ZK96Vb6hIbXIklTX2WP6ZnTZkLeTvwIIxxc
noRV8SDJxYQGgyGxJXmN6j/iNFONWSYvwQu2XlNKKvGWs8b9BZegByQU8lMm3pIpo7Gh10ohHxm/
fMo7Xv6AkCIZiYxynz4kH5H3DVk2x0UHXY9ZUFgOpp4so/BNvDfqjaBKTIs6AkUWhBlTx8eVwVJj
EoMr1UhXq2g2+dX7flzVZ5YubAk+hCNzOgW11Vc8AsbrRNNiN5ZVLjwhdwdKct4lEHkAozl+jTxT
Gn5TfOSIbD532Nfn96CLNuC3geeF2peVkIh1IwTenAysdncEMC3lg82RCszgQsyTz/t+Zbrlw/VO
rVAscIX/NYs7XIkBsthxbS+G0fGL8x0W9d0hHO11ONGTSUkxdJAs17RiaHilbQq1fi65mdGe+vls
3CTpBwhW44q6051iRjBsWMhXI2k8TCQMB6t1OmetUj0OtBFZ00VCnvSDz3o5aKHzKDBTD+iuUUn9
jpnuQ1eInrbh984u3POZDPG4UJb6N1uobyVBh5nr8VPKo7fBFn9JabuZXHm6X4FhqV2cDtTVXJqm
v026/rIjEU8BGg0DZtLXmVVjeICTASyqE58kSx2YMDe/LQc6DgGyfMCr+PcscXfXnhRcsnX9mlyt
sBR9fVFtz1fW2P1HHoaYmWfqoculilMEdADHI7Q57TcOQq7/TR9kbELapKV+/SkUkXRsHUJFBwAj
AucF1dyULQMuQQ3fZ16g5KTmoR2YimY/nLc/tepj2/i+bxS/LcHfbK1ksSMGNIEOZQqG02BSDsa9
7hcmP/skfgpz8XTvuEjYpCZ6EsrGANefyVs9XXTEz098PAckbRU6MxX3KCfiyfKYUbxOEoPcfmkL
0I0h7aT+GqDWaGu/6oP7u0A527mJMXOWfIa5B4OiojGoHDzaCvdMR/RQXgfEIa03L/o32Paxv6Ot
fuwvlaDSXapyGbRqlSGfbMI5ehMSvAE4tQRMpliaROCIZyciPCuOSsLc403GRNYUdRFFyBVB7UaK
kg7XfXTd409lmfm/JnWpog2K+87pUrLzJSy33wLlusT1GswCN67AFrvNjtOomflwwxSTUUVer4mn
8VxJuvlc64aKUBtYPc0iX+8n0//JqJi5PAGRw7jVYJIKchI9KjfY/OEYkyWMPZWUl8EyJcHELY7t
YEwHZdW+CsL2QxfVtKg0y2330wntdfCi6gCb32fbqu6FtKbYwKZ9tT2QogKkcIydSGc0ibBEYAO+
qrdy+lIQf0K0O4CvWyWiAdM33T6O89Aq8GV0Vu3kjQz9/zmzP79y3Tb1vudaHU6jAQ3DsFry6hrs
4WvuKXuKwSw8VmiFLZ3qivOOYDvL52olIaar1De7h3A8wPdqus8Zu0aOK9+Xt5bXG18GpVhjYewU
IqXXDj8yVcdYhdIMJrkG/ng9d4jz5lcx1xMAFaUjl72hJewba0J5OFKMlUAn6DO5Aidk/UQeWrXc
EiuRbSTljHcTPW2cwLLYhOTZ+Py1lCbFq9KFoP00ifyElVRnTMkryJPFYPsQtEF/eZFhvSiOzJrG
lvXz5sIM6pBAk8Vl2AxPYe8WGZRjAuI3jKCfIN4OLLgGEbu5xQpyQMprBIjqbbWpokSzPFoFyPTs
HIpMYsca10fehS71b/RLIh6l5BDj85ZKoxfteqAWzVt8wlxDkEa11zsqKkOEPOvvDAY5xVNPslvf
di8dDg/16U6NN69GqE7FaFISYw2dnOjToE8JdDHxou5HpCq7Urv5Wv85bFY/1auuJi/uzlO5NQPa
olnsJgoaaoTp8IfoXADBQ+1FQ0aO53Ce1290VO72pHeB5QNEsgp0MavDtcLEUcEWP4l3SxzHCuaq
4jN/Q90DPKuvNAdFZJeLWjzoxK64Y3ww8yrOKAA1oAT85ucGksJTeMlhZ6NPwpOMmGNbZsqu968b
qA8L0M6k5cIyNbUeawR5SIWFQtigZT9lz4kYv+psH81zzUFotRVIiiZOsiISOPEL/7vfduOunhnq
9NpsQfV9M1yG+rGzfTKi0rREmXIfVTtA9r89W0G5zwateVJTi0UeSFqGSo6Vr5jpzI4KPz5Ulm4Z
oLPd2aSyEgtIn2b2glfX2NPuxJ/cSWe+T7r2U2YKmEwT8sBOQ+cgY27tYbxpgHyVT497/H9UZ/r7
ExzrcbqphtECot9pKZ1mKb/YwYDm3/YZoUA1tCEHvqL4WZZaBJuwZ7N8FoU3LK4UYXMFXxEP5hFT
reclanmND71efid3lzatTlpdmRX30OhfaoS1i4FWlQQ/ZMSNPZQ0mDYLl0l8yZExJpktnlvzaMGp
E6o37//s0q03rB/AZKQ/z262bRiunPB5jYCHe0PifDSDLNCah/oH1HSN4lvqJFbanea08dflS6fx
J9F69wimGvAj0Q6n8JZLsFDN/+2qUIkjL5WAZFUgKljCMzAudfcPKBy79LXJK2Xo08sd6n/qPOSC
nAgDTpQod2G1vQoMcbzuxrtgLQl7TLTBiOlkEi7A6sM+jfMBAnTRqNdX9wmvHrn5fReOMrd61S1s
gGsk/Ppnd5LVs+u2r7gNmo/JSEmxi8+MWjNQfTuFcCSO1j0vbgUyiPJS+8sWed2CA70L18qqe3mo
tuz4TVyhlLgtVo9b5YH+/QsfyJFMAmrvdrmDfsXDou9B2QlZKkrXMncjZXU0ni4bRdzYnJQ51P3Z
blORXKDq42kYIJXY1RnUTisjm6kVLfHzfIZ1gHOEDLR9RyUv83glIvnpNPuhYDCnzMh4x+74Uyjt
0Jc0RHDyuhagTFSXKlBJyF6Dm5iPrjSag6OkpD86GM8CioiDYbaxpJyyWBfvLuZJVhLQpzI4ScAh
0MfVWGesdHbYf0cx3gzKQxrAOLSt6QRDN3nVR72TOp+nfHl9pKf41OebLCkb32jBE+evPMColIVE
+Fa3o5Sx6xjM7jlINtZC7e5pek70TnnfAtHGdbehi/vg1EID+rQSQwY8akZIsLoe5GgjHFx28+Nr
UyzngQUtKQz89wpS8DPj/dZU+GczvdSDWWaoMiK2pxGPcZ6nVCEVx3u7ZKPLV4Hhz7Js4xpihK/a
+wkvPzxyhoJsLmpXVpEo0/GiM8tLWUAJdfv/Hmsl14vt7GeAlaw+wvCUx9qK3plnhtnHHN4+QJiZ
5THgB0UHRUTMj6JcfiNEKrCmDlSepUvlyoFmpmbrbHnv3U8ZUAxUfVCFSkw0UoeKMcKReqe8vXDs
4u8NCfrxM2qiW13bkBdOvdgVRjIVeOXJrLzzl73gJ7iq+vXmLcLgW0T0dPP93bfWzjgCxZRoC9xS
e3I8EX4HRfBWtxLglVwlTS68uEr/Gi+He+aFPj6YEmXESjQsxgHJl9VMCqaA24AfJNuvaB4kK6jV
tH/eyWOgoy1fWypXxsRqb2SAMg6KyT4ANsLayaeAZL0eewjiU9O7RTof0hv7VX3peoJA+Xr5gVDL
Xds7l2dlgl2DVmf3iYes9r+JRLpXVsV8Lb6R47+GE+7peHt82UfvHj5ejnB47FCqXz+iAoEE+QeU
BIMGhtx8C9uXjEPhCQprf0yhWuwEV8HlnojONCCDDxRh8bk1/WIUty5QywHk3gv4zoRNm+VZgdCE
56s6/dmN7GXGEHtXj9eeErfkRKpqmrYRAaPB/ABuQfC+Z5EqjtQ6REuuti2eK3NhC0nkLeX2slX6
ET257+2ejA2a0fQuVdPpPH31shaFlUyczFuaalHbCIZWxliW6Z52qouDSzQLoK5ko/P7r/cpaNWH
81HzRpSqV6A+W2P+C0oWYklEFK30qTfNECBn5SgZRe5quNGXP+BmeNRKiRYqcNiblBOpaHcpVLS1
itVG1btkQkV8hiYthWbCcubnQb0D4SqTUpehVE7p19uU8JHBBEWNtlK3hC9hddGXd+/p8TwzC+mo
m8INxrjW4ztVlovsP3HCoxZkqDFh9/0bdSuVNN+0F93hNViShDZh9nlifZOeO+zGRoYMHxE1li9W
IHRhsu0CDI/rTIOu9FXBZpVt+PdmXosHoeh6rSZOGpLBJAhxtx3Q1t56NKyIhLlSDpM7NQWxl5cP
KR15xTuDEpid41MduJnhoxBlrPaLEK2lNrUFu8TT+wyK1E/Q4x1W7Ati2q2zLIN8PajtpO9Z0rs/
Q+vM1MDtjF7jOxZ9xYUqxZaHTqpMadPhJKc4+wZ497Vg91fkGCzp2ohRGuGakm6KI5dPqr2VQSdE
Zf+jU01FkkXVBK5YxUkG2q2oC6tgjDlwNhmlCQ+2aGdlK1WONFbbyXAwaSd3Gm4bPOEt8YydTq9v
kXkcfZmQ4INazS2QZUOAP9iqAYrW8s07UMoVy4tuI/MJlaNcc//+c/6jMwDPDnYwy3KjH+f7OfcJ
93qTWlmU8//+yV6E/PH+0+tvYRUOcN5B6qpjlLzPKCG1YeDDqpuOF20kWPvQYeONhN0k3xD1/Zab
Tn7+bUK6l4PiCxj48qHS5OYPx6+C/5US57V5cwuVG9RJB26VpTVdGpaixbHz/io3m2DDqPG9CWSb
+sm4nyWYJZkcTesqbZgQCrFWVx5A2coZKdlYQ5QWLQlhOCeDvSHXa0C3pUBT8Q94QTkm3R55+7vf
dwjnw8GaF0hW6PrMSa26g/4+jVRU+c5mFnRugw3k37JToY0qWvhELlrcoqFl6VAkvuZV0ERWI8Sm
PI9vIP1ZUd2lWW0c3heiaoxyME2tKG/gnRwIdWaRIrppiO6hd8op0w7exGJgN2j2kEFAHjJAN7rj
XYG99tcbqWXH9xGpJsO35JfpCw71Diag6j46dKO8ebbjv4DKFuOPzctypAThvYDU168zHvaOvWcq
CLFSFc+hijiPbU7pheFhi/KpIMBb2Z0AC2dbj91jNQ3KPvqlXEl+UzKUjanYRjmfgx6beikUoRAG
eawqdkmgv1H/9XT1NDSYvti5FNYkX2wTl0oLw736GRLNXIRTzInLjDEJKrep2O79BRRU/XN9eAAf
RXvBMFSyhzLnY27u7m228VXd1hVdx1OCK8kh/FarFnvoORQaXMk08VsS9ZzKMQs7V8mqtRqf4TNo
P6Hy82QFrBc3jD8waVgeiXpizpqoz8ryG3EePuRwscXQZ1twDVCFPpUllfc0kj6JQxqVh61Wkqbf
JgnrCVPXfvtVbMzfXUM2v9Xjmz4qVaOUAf0GOPMhgf8xAH5TPYVNcl6AKslcBm5yExEnAHiaqkxW
V4b7EUm5nVuZp5+CNPTrPpdC7KOUaIoO86o4E5UXZz/HkcLhJFeW9DOpHPjquwF2MtJVrbofomXT
UY7L/gLGeAWgp8cufsKO7uk3mgo5oe4exsrs6nWwGoobqoE+l1sFEl72Elb4RYPxnOtlUXzprDii
nrtOotHli6K2a+z6d9QpnDlayEXG8EDliKAc/rKQGaXVSBjZftwefM7ZkDmujwszypuol4I2I7lA
F6IUrTuTxuTcFxC9vaVrHbM4JpsfnMLLp+rQCAx8Ur+dic0eqM2R50SvVg+qBOJ0mU1TgHZ1Isnb
7KfDO6zoxYph4gFwYzSnDNUzgGMtkemgjqVacaqQqTluJ9YJV1dLThomLJUYNul5Jw9FtsFeLlSH
2lBSzTm/OOyobQvO8SniHFAcYB5UkXWBfLR4BD7C+sMeFni6jaV9pVRpBMzI/SIynhhbuTxHGj2T
viRVwU5l7RYXvtEFU5amGt4M0VKb+jv2olxFhzNSxdyJZucQlDBTgzjsKmsDT91a4A8KR2bk5ZQA
zYQU9XEhGHP3fUjJoDuATgZmScQK5oJHi8oDSr6fIJmXSv8seEFrg2F+3NQqtY1Rlwy7kYkaM1UL
4h+cL5hW5XAidqaP9zBvwCrI0HDLzJ+9YufH3YQxnO4uPejm6vDHOUorOPmA5B7KHqK8WQIvJfpc
XVvH+t9sCij76k+fo90kKrt8eGO60773D3Oqn/kgP5A6gFqsrVRPHMQ2k/CbdHKbSu2AK7Ft0eMN
xLmUITW1N5lz2qUazKakL/Y9D8fCB152tcAz3hZuyAFpqHOOv6ZDYGD30d22ytVyzFN18F6yOpYo
s/h/yb4I+7eV4159bBy07a2GLHr8IAoO/I+u0AAwi/mQBpIQTA3/PufNgQFXivPbG0ed9ABFlJjg
XtfNih3nAAZj81A2Z0dzXBPiu5icWWKxG8NpYJYH0Ix1QopbDpuTR825yHGXAK/VpuV2qfmu2rxB
CVA1B0Q74yKmxd3cdCds68t5Of5qFNXmQkr+bq+qBqmBWFDsqGvkd7X9rBh8c+cdpAr0MJAE8COW
5Bmz+ntqnOv/lBRNe70VJf/FDSJltlBNb2kwqOUoySrXMW8oIQNZNSkRDQM+4oil1V7S4bHEqvAz
Amu9BYCeKTdfSJtagTMt9Ylif0s/+ECGLCIA9aGdgQFSaf2zInQdJtid0rUYrNZCLMZXTa8Z49Sv
HaiHdOsIBAK/sshoucdbtDLlPXIU/tVMZc72Vnzs3NqDJocAxMPv7nxPm/R/uAQ5VdRD5EC8DfUq
1hz+QN+qLs6JA/2erAPbeHrAtiPZ7yBpGl5qM2fzMrIG3ZkewaX3tl3pg/UbdP09QxXA7Hmq5AR6
sO2kauyOVj9HWUlJHw8BdzcKhG78AV6J9edanZKKBvqzhWCoCR7SGkLF1lIdfxHq8J3NP7JsuYBI
ZIKBXxFjZ3kb6lVlvgfKQbFX8sf2WmVnYbHpkxRr4Jtzt+MuAxf7hKrCJOsteCUXs9F5SFLEdvot
aW7Vt+wK41ANAno9+y4tNbRyAzdad2D42QcctJ+L5oJEtqJ3BbBnI9gTUbb0W5ojm4qL0iNgXHXl
9PWMSM+enJeL4Lv6E7VIN0eScO4VMaSqhSrR5OyrHEcEbpkxOqxgNVlWPxoGd2B7/HvJ2Y/dpcp8
iprGgrI9CMNyRNzmbwuxyMiTkpXYt/TMDKCKvstKx053qf56lDY8GxEtN75Cvf0U1RhMfLBHSeoO
tZ99Dbl5t62zjPC22+teprB6j/QUXnZA/IcX2ahSG+eFKy/Q7EPIaeBf3wILiA0HYgOqGMEMtEkC
IxMkoz9PUY4jlCW07NRdHKmeZTiH0Jw9VeS5l5OQoO7cfdryosz3m4WayY/DdaaahiJO6tSVxI2x
gY8be/SEmUjM9DNm/0bNOtEgLUtwJsz2WxMFIPyOpzSBiKTO+8kt+qLhC8ztoQ6aqUKZ40zF/1Q8
ZvRBU5OUPP1X99feyo4enlNF5rB5hICRgxoY2PuTEIkG8uGx8YKNYZg7LTkGvDN0quexKD/ASxTx
N5fOFomomk7KVJHPAZl5NZH9wulcvnwCHMqJcrhaHZRgG48n3J0VAFh1BX/QqNEjHqEZCPnCBV9d
+jlurtQmKhQyy9d3GuEVNKQKcx32GGOq5gxMrFurqLBfrrBAoYyh/pKR11Qe6PnwLmWi5sMeMQ3K
/TIyNNOq4evzJ/42OI42zAij+jRw5AwIULyEyVHEUf9Bgrfo4HIsqslRHnVVAHQL4DpBY/2/PEG6
mhe4rNTTfGVly/h7kfnBZfZTePDbj5uLdzLHfcWMnOwc/DNzB8ZWia2i0QhwAG7DI7DRXRGfGbey
SM38ejQBcBtuCXoUybOQI75e85f95c54u298Bdee//bjTuoftF0GTkmUSnIxYRn/hop0P4c9XH7u
5VEPJ6qF2ThrTIdEOv657uvdXB7cuFAxTd8FEYZydhe8NHkA8mxHxMA0Z1VKldRhVp7Vtb0twIG4
ajH/KcPEXuxXWKIf6B0LoTQoHWKDco8gNZ/ndf2QfNk5A56WEJUJMyQOpDhdjBRPMPZPCKf6UNiW
ypYOsXN+NCvnoG3EJ68pm4xLUBLdrMBkSHfrMnI8WYYN2dZv0/ZXUAAgjf3QhBNVEHfgJOE/yXbg
BHaZk9SW6qs/91XS8fqy4QeOFSYbz4BWzSaBWuofLIPwG9W83YvgY1hfmeUyh0XGGm/XNYqZqLcU
TKiT9iLR1m4ffjrk4Du+5LIVamRgE3VIKdkR9c8SrBx1rQASE/kKVP5L48cviaIMOssZLMZDCwrj
TqfhjxwPmgD75GXccvuZUVOqKXFlhslXW7GDSqHw4VzcOftarOOxP46jJJgzZ85mfEn+BJnJl6he
rysrWfcBOG8AR/6xpHlAWsejXTuK9EayYPtxgsxUBHPL1/9LmcBgRNUNdtnn0xV+K5loV+NxWUew
tl9M6cI2mwFPmbgvnHQ+lljq5HVe7UJeY0UZ6XLeJF3zTM38DgimnM0nS9fUdQRdb78CNlLu4qB2
t1YyoPHMau5OeW067/T567u1FQPcYbtjeDcnRpQXFmHORHaOjsK6x3zBlQBlVDEN9vasadNiyUON
demgQ+lcxV02zSx0s/zGc4Y8UxfJNkNHmBK5rsaiHtH5ty9Vlwc2zbQ3nAvTXbrIN1VoUv8BwRJb
2+8ucerBKzCKyhPREXBOmW7iak1/1pOPuHxYzziQm/H8j6yOtWG5TiJHjqIPI1IoyVP34tWV2bY1
Ql3YixMjP0i40eqdlG4Ahw0PZ5xp+wsxltUAySNPVJ4GabtsnVjOg0M4QNryWoGnOrdLCCHUsw3n
uu8idbRZvtCsKlPIGxNOcwx4bSMU0/fvaeDCGPDE89qH3Cg15gWE0zAQ6Vcv98EF+1o4XIh512H4
MsOGHmIs1x7HjKUlTnlp5f1bp3RJVQ7kpAyX1kscXBVSaAGKJ1djFuB2vZtzvJa1pRpkZ5wTHaLf
2B7L7UQrn4QBOf1lPMh1KqiY2G2xfq6yyT1RLTjIRrVM1ushKVCgitnzYrXTMatjutmZJOfmlOon
hKLkqcXe0LeJlOTH6qUP4KWLYvN1HDkUMhDHAHmgLCbjRwihT33v4aO19ZKwvBuotfOqJxUa07h4
DNZ8Wom8UIMleYpGjEV4Z4E9tHiwRqOcEo3o2J1D/LuumfNd6sE3RhidcFKXO1YzF/MttH4leDQl
QciRm9BU5OfNUMVyyykdb+BBVDNezy1lHd58Jk4OqUbJIBHYiRJx/kFFtUQ1xHNcTOyW4410t5KE
QYRvspAJoaU75Sbp9ixY7tsAsRw33JGr2wJ+pY66Te9DTcnpJvQH+4O3YB3Cy6FUx1+krZGPhbVP
qFul58bU9a8PrLC5ozS9d3suywVP53pPm6peMVdxhlmIsTR3/ZDZeExVcx71BjtDR9a/Dnl4J3kF
LcQermXFgm6HmFU1lpJ6+9qRy6dyGJiMWc9Vddy1l7U3P/IHM+HjNA3UMGXQxiLzI6AkRB6ZbVEM
83y9yJrxmBfeKqZNf8mKXs+Ve1BApuESGr7ZsHC+hwfbuSLzW9ZFwzicJNpl/nxmEjDEMdolgusw
6TETn4jFiZO4lB8tCFCWVRosBOYdGdy6XxSBUNeMXpBxT0xNZh1n3yNtmjXfKGKhr7UgMiAGE9Zf
3RUfNEvb6QONK/gUA7Urk5RALlhhNZXXt9hQ+4JDpEHUXOKc9a/r8LX4Faw1CnCemOTAp6BRRLXX
XfW62DYE6GPDHAgR2lJdnHZmi8PB2bueoZsl4mV8p3zo+o3HY/CUHCgH/4jEPfuW8BN9mWa2dS/X
8HA7BH+ySQtALx9YpCnNPBii5kCFsjPk0lrmmpPzxF75qOZCwRdxGCuqSoY+r6udL8dcMPRByCrg
HNA0TOZwIEuPh6vU0sADOu3ZSn1oLJEOn9pxXrnd4uSCIqAoG4wOLigT+Rsdyfk4kME0/ZkLDiI3
rMzWwzMYPbB4F65NsnZB6r29uAi+yv5ieUGimxAyz1ZLC5IBO4E2w/NgjvSMWzRhpiA0H6oeZQX7
k4JYd5lhluZfURqhY3/qQStzrVBaskMbZitBzIIOdts27zJSovJ5w5sZDjIR+eLZRO2dbFczZtr9
AqKSVsfqtvs+E6x2lZYR0F2YTILiQHz2HWqUt/mJI/yNOLnZgKNwRq2AMjCt6o5n8JPETL7k8chR
SkfM9hxODLvqCJD+2DFSY5QqBoYeVxjPHyW4rQXz3i7BgE3Wl4RjoU7JvxNyCC5T6A97ZX0SkEtG
c9CliIbno0CcAlwHGLDZEthvFhD4mcTSUKjPF2+3LTptvg3ZmVbDkNlu3iF0HG/SVVYKeN65/KKC
MYc3riaUrsCuQnOCRurNQMkkZmBz7AQck9aK+sY89/MCyM8pxmaH0iVSjZNz5islLfVQCoez/PXI
YCmcuMLOCFx5ciI8Q8zs5R1K7C42cP/fFk7DCx48s9vHoL1BscSkPi51khwY4azW8lNswZqghS9V
gLomDUwOs49tsC3V0VddhCk2ExcJatjFQjsvJA2KCty55VW/la3dqddkPWqtCaYXaPekWzKsrxMe
BRqL2RabjWtsdhgtuJ8WZLOmtVBiTkOTqznZ42cPXvUz38T8zokmhW+J4NxrtRWaOHJwe6NRY3vO
bA0JSx1MGPR9+9nPU7PyHmZwWhhcc5OrtNiWYeSi1iAQHgg0qMMXkp94eTjNbKL2ZyPP1bpT4Gps
vuVQUwZD3nUA5PvjNWhCuo+jGpl4FFk0K5bl0wEouImBpla1t1eaxfCw8tpnh8nB5+iF00ku2TAO
5z1C4pBdOGLbpt1p3QP0ElFkNyHKuaIt756bQ5PsdQXYsqlYHJ1wQweMe1oKRri9lvBBSNduApDC
XbAcqWG65nWOV2zxAbt8ZriXlXIx1Dpzvbdq5ATuT6akUAMA9NPqMIKLrx9lwXTWxAVtbfuNi1BE
pqiUpxYueqvTM7miYyv2HsyOT6DDUklfRpZ4R6+kou6TnWDM8mltCoSZkcUOae2tb0c3QuX4jdIi
b5tziTcYI5Qit1wbs/4obzRMpdlgSQ5St8Mbqyfj2oJQ4fHO0cTxQPqOkq9uLAH10f5+YaZjL0v+
yogCtC2k4Lgzt5QA8dt52pHhOkDFgEHR/YiCwYasOAH55kitenOvynjsGSqZk+BpY7NAR6nsb1tV
7i4G/6zFi2qaf7pvbYBHcWtevEnxDIzXVSCP+etMunznZ5wJXN6W2P9yQNL4H8tLGs0Rb+5T5/L0
+4JzEGTD51Xz4yiygYxyMVq4482sLMbYUDHmX0RLGX1wObIuUQvYsD0DKNP54QZOWodxkyD+lwoS
1N6b3hSpTPm6HYzHt/WX5C6sT61DS0E0oro32DVTtuL4ymuNieUOZ44AWgqPwrZsDmxnfyL44mww
P/xM1XaDtV+8mmIIZgeUGZM4OLufRcdckdAUPyX0hKiwjnwlN0uXZQhRccoafFS7OVxZPusDuPsa
hbOgnV5UvIfGVuo9q5QPTpefRq07ZpKcaLKxzSdkAlLiSLiYUcr1klXIIO5l6+eq7TzJDNCCJChC
eVkXhSb7xcE1MaFUD4EAkODK8yS82JpI446leyaYRlBO+htYI20wz/O/e8lEU7nBHbjqO8/Iz5Mj
xTxIq66brMd6yqAk1UdOrPi7MyIpyUJ1rgdjSNdDElP69qlmMLgTkfu6jW0kAdT4KIxidnhxveY9
7ytiGvk3noQc3M1tW+bnDiN0FWa3e8LyPu9FVcSczuq0ib6Fv0v1i1+GVUT4+esWtd4JKNrvmOI+
DCuwOBnSOWFifgefzBMQbV3KSSrkmkBznU/WSpkpMJS/6WarUT2ZgD5SFOeGCETre1O8Sr/grPGO
EcAmJLWqOtWJj9pGQG4fAWIbtvnxpgSeVILOW1uR/0GIlhxkhJA6Xg43OiSXWmsjayENlgqt8J2Y
fhF+GiLLprQkuEkLNACIxQAg2ky8i/PHtjRUa6xqKFUkaY2Q0rhP4pIp+JOI3o4e+lWSK09Ut5iN
wdyYQvJbWV8mevej8ULt1NNCWDhYbKGimSFccNfqrLTR9CbiuweOywuinmL63jAqsYTq7hLaBQRr
eT5iJttfnkBwaBuON2CxB9AclifvnAYoOOx+WGrXHUpwYcrWqc30dnYpsMFO0aTh5pRNGv6Qt+K+
+LaJGGxt6ydAmCvMnpi2I3JL+P8l+Yqt97SwmkN+o7IZy6K7QMBePrG0SyRyL8F9vWgqaQ4GaYQ/
adX9p4kC591vAMmqIkid/6ByWMYsQv2nReZANrG3sTcj6yrAvgzY1Zw7tNvyE6aKz6yO7ux9n/9L
TxwmbZaQIxv63mDswbjmlLIErnYMc8xBuYrCwnHG4iui+GcanQ+Y7HwMbYMI4fUCEow7WBwSHWh2
+POWqmWxKpnNyxhayOkJCwob0yWd6BzLIQmeLMLx9emR31nN/VGpF1rO9YgxtPVv5fiR4i3orpiU
jGhAvZzY+XHepWiZ8d8gRjpfy5ux+imaB9YAyImFyqPFfi7rn0ZyeUBY1QnAK8vluDC+VARcScJO
X5GYikFs5ME+XuvX3R1b+08W9fwdWbrOU470hkOYyqXVNgEepr2Ef2USu0Nu/RSZcy0zcC5jKGRU
9aNuecTIQLbK604Q6772jvTltl2ZRBdbgxAsd8rwstiJYVPJadOMvtprYOxEPEJLmP1pT5JINZJR
dmFPv0NU134d012artXa6rkFYELUOe3YwQzZR20RcBsllrouBFRReCHgsESE1ui6Ys5jzkLs6eWT
WWVy4cRyZjiYfRL7plnSef/uWWTx5il6UocAJaEceTMg4zkHjgQ1JKCw0NFA6WxCtSDwQVmN/Ma4
/BZGKw9cMLCs5NYhhrQ6zM8w4bRO7d/4HqC37M7RQ1LGcydBfcJxK3OXjEwIM1l1a7D38B+K6UAB
+pDS1qSwytNvOFfkUFpqVjY2zlBSpoQ9/BZ74eO8TJGnQkGfy308yaR1T86oP5I4LBC4p8BoV49a
2Zj15XsWZzKYq0Yitc/CrQ/GEs7us0hwlQFD+gofGY5KtBR1U/4WrbQtEjiM0u0mwgtQKkRXEspb
d9/1MNI871APmm6kXVJkS8Lxvne/IyPXGI/YysUkmDEuuRJq1q5igOmj7d0qO7OcPlaNjj73f6G+
aPP9GIFox34xjpQiLAXQrtNnv3jfkGrhXtdmRK0pKktRHni2hDwPBNxK0L9+uOu+G+qh9XmAPV5p
UO026O2ExmPeC/QwoqwxwVFES/EN9YfczW1KCN1Fpn2HLrFsjjuLPj2Jg/uwq+jtSNcJjLnyfmMm
apMr6foSTfwyydH5k3ov1aMVRQFqE2U5OBwgHL8f6ZhS3kS9dks2dX611nFbM/13iZsRVTCATX4a
GMJdeKMaNGoWNm+iM6wqFEK3J+8TlXc37jJ1Vqvjk6JcwtL8aDrhha3EWD01u9+61nS6g7re8wQO
eda0MsDKA/+sCTKEPpR3rAuSVAYeXXY/2Kj1KguoJBnd9fbbBmvhe161KbxQFZn1oFk477sDAFK6
bEYYemqtmX+981XrwONHsBsBL3xh9gr5W/V2WvbZB/P+FjDuNbkdkoN1nlrZulZs3DzzkFKY6r1v
yJ7yPnfEaAmcAu9i2OoL33+xgBaeSitaW3AMzpTwZei5FHNm4hke/vsG4pi0O+TvMLz84f6wGC83
dQZT66VCPj4HXYuf7cFN2tNPSSpUS0MVumoQ9wKCXRKxLjewkIkrUPk0XVYEirslKVKZgN9qkdcV
6Zttqn8QK/rDDs7PrBHA82kgQqBHfHtPWVdYybwRln239WQoiFe2u66BXx4SToGpZl8k4BsGs4Pe
h7X2JRsvIWOnm+XeXVLdfd9Ayt5TNIJgH0C4PArAE3RaNi/ZQKfDcT/sulRa1y7sYMZScx0sX2uz
Rha3Ni6OWvZR8LzRs5cjIpwx5ivC4cDr38INGGBWs7TIV9vLrnUctnhWgPa755jrymILuwobYEes
OztShvwBLyP78sELDUbqVeR1r4hFJIOCV7CI/YoWEwGi8scgZVRJMIqp1tbMHnNX/mgSx8tfoadv
2mcIjUUs+E2pWVDO21aqBk9uuEK/8BSTrSXYnp0ls9eaD264FlDvxZ0FRoVnLjc1wYx8LXPpadbk
oFTP1153rTAWyBz8xTdD/sLiOzbFSWQny4hhY/BhJ7qi/Rs7P0GaRKlhrwQoInJ3KIkPoxezdihE
Yzng150xaD4dwHqCb+lP6TVihiXo4xE8ycQR9PAbQhVyYxmpGl3RcGqKbDyTkdXtZ/URq2riRjGT
6ZqmM0fNvcjZqNzfWosPLcFI8TGyhC7GFtxU4ubCXj5Bwo+AldcW/A6lH7LtvBHvy5VcwBYG8Hfq
Sy/9lfagDqMhxfUHMdQnmCAwMacfH9PeMGGMGQuCrMverbkpNAinYHxtkr1jtNhx3KMkI3H31NRI
gZ3q62APTgaAWWyrDAsGw22IVyHyBrp7kPm+kjqsyKou6qK+I2/UripVcO1zKQcYAnPYCNpF+GBZ
zKlMXBjFpqTcz7dAb1R9CnyqB1pnZHphIKbDaam1+oEoIoftQWSGZOjldgasOK6RpWN1rBMXGDw1
jrU3U7fau9Uro3SsuTJqY8/K6Y9JxaUSpfXTdaRsxMZI9fCHNcu6xo/3+TYMae5X9tAgu14YqVK8
X2PTpqtTlQuEJpbT35nLAmBh+x5KmLiRBqkLuOe9Ihf8e+urS4+7vJ/owi3pforQgTNCx0VW/CPH
sxGU386JSvOBF7JvqBXBMGjH+SohELtI3onVC3koMMhjeztzZdP8//4UGeuUWLTy8JQusNs/eh36
Cb97unmmHxPltt2Rml+zfzj1oJuMZ6N0MxjYKjoxcHwFRMyYHBmJHTcF99wlTBcZDXmKLUMFAMYo
+1VKs/GlJ7ZmD5s2ZMdfNlxZOhSOp89CO/dn+ZQOCzB30pm/tD7UXjFRPXd4hEPiJXb39lyQH5ZQ
VLwIenZcL9QBNtxX5m1769IjWovlf7oACWtoD9Tfyg/KEBj2QANwoy6e78IKTIFuzbgursjvpf7D
c6HIwMKMTAEOJa2luddeTExQZh9Uw1B4/6p5EJdQ5oU9F8Zm5+9cqbDZfO0wvMuRV+c5z0j21i00
K4Kygfv+Htaci15M9bTVZSdHk6VZVoVUFnWhR4ZJ1t5xSxX8BJ0iHBgogUZUbpqxfT5oLHsW+UU1
IrNwrNMJWTmDTnfrkNZiO10C+gHqrTiknY7l6/U4RkEZZ1b4eaVE5xnbXgNnuuyMwtO5zHfhGaT5
mkG5q4x7xydSegF+NEUv3YzJFe0GTNWD3XHrc1mE2axzq/SMLWvsw6RgJtNHZeaYbqNCNi0t3PYz
evBQ7UgSEcZejCWr9hxSF+Kw/KI3iTv5G3pxaw+X200neq0snMVn8C5nahNUGPP9St6gS1ItekcQ
BT1+BoqJzYYAAitFa9Mb9/27hYEpQOhk0DlB0HkgqxaUtRjNn4zh4yhnwF3wZOLKlp9a+JYFRqXI
4zplLoZBJIpcomsk+Q//Q7UK3+bQI26ZWQeNiVQ8ei9Ukvj8AQOPz9dnGUG4w/LhPyDKyPJDkwv7
Dvx3xgMj7PXKzwlw0gHxYcoGYz23EZZ19RTZ1ChWW22DNEkpmbEZN6Iba7Rz/10iIiBOJuudGkju
slA3P1aN2SFksT40km6tjWUrwfMRFdc6xsn+pPNnJe3oXvR4d9Oqj2Eut8nszOtZCWsNzTVjVO19
JHAcwKZjx7RglgKJyEEYmbEqU0GYPwfQ542wiPRs2zjsj6XWzoJnDE3OqTcUQLWJk8x7qntMGSgo
dLLINFhxBS1MPD0CxhKX6AhWum3V3hqRY3CVnx1qAL7OCZ3zdp7A56yHJlwUiIgVzKkOO8xrXK4B
vWhgADNx576zVEwKeBPqL5/rbxwor3y3aycLn3x2dIjWQWqkZomDj/ZYCGrNun99QuNXUVlDaLpN
JvIwC4udyDd+sBWj1eRp5L13M6mpgCyf2UXIRvYuTEeP3yx6/e5rbAEd3LGv7XaUloAv98cEn2uc
RHYLje8jwFVZBtnjAyXbR0QuRKcjNie3NEU8g7ogPNypMcUL8Bebrpc4+feUfPoSbBIiH4Bb7KBS
cnyGzaKlcoWkk9mi+Lbj7IO+4hhqWKEi3oCCLHc2jAg4wA7wzcliCQbU7myTLXsIc6DnpaxsMGru
m1pOsdSzETahbtETBdlf+AdMhk4EvwaInJ7OgsGevBen3cOIIqKeFAm9ZalocLSB9j/ukvainRJ4
vigEqFh83JdwbWCsXodHd8cHC/G/JtqVBuZ4IQIBgRif0cb1Cgzlm8wrOtibXq9q/MC8BxKuZDR6
C2nEVZ40m+V4lp7rOpRYDhq0NSZtaFGJkT6KhMMtaBxk9LP1PXRdOuQwWrpZ2emGImF4roro1wNi
HgEH066txKNCPVON/6j5RfXZg2ep7PmYFzfDQmkT0/u+3YQWiueJjrz6wDDXRHjRPgliY2J34J9/
zQCM7J9zsEyd2iSHluT7I4ub/f5jWcuKMp0MZ6c7pDEe+vBHREkXCAxJb7ldGq0zFp5L/qVz8a8+
4erHr8xw3XToqmaCDQ1IOJiDXou+tvxvnXDkPmBMKMC24tR1rFcX3N2iVK9JepI19EvX5X8rAF/k
1FoNiMXXK2iUmURn1yAoCfD3gTOwpTFAO4g0v73ztpyjxOShwiA8GDdjbOLQ2Ss0C/DH5mqYXSh6
/xrTpfCt3j/+hmAz7oW4MJ/RTA5WAdJ3tdIebURM4uiiB/zJYduKWknPg1sUIFtNKiCyGvd8YGLK
1FIg+1HfGTuac4dOXq0B0RPJ1CgYZ+L3/aepfPvChTZU/wKlmvXU6uGig679vaj2XwlRK/cVnhYz
H2ldRiHgG4QzjYlXVu1gddWi2hnWoCUSTsgasO7uFPtHd+hPaxfPIn4RkLle0YX9NLjuvtr7pusg
2sSIzSQhK+YLz58jjEVjuVk+j5p7uKDTr+ZSwcPqv9iKk5XS0H3BFxNqZo84RzRZKoh+z0k+PGSU
oeKMYGVBvniy8SNfEqAhMKutKquWT3fAYkhbb/wuMDV8GIlyjJhlEoHBukx2xgUzz7h5lEIIi8Gr
JPDpALd2wQQN9z7QYMcpIwpn7rfL7ARs+a21mfCae1zcSUSsFYdfywEicJmVo79UtRAC8KTQeQ0E
Aci08RSnxnk74kjApsTTg2XncxFICR2URIPeQVz2FuACLOJq04xil1kmsCOPXeKQ/QF4a8ljiWNH
8fn6ni1xXK9TdzFxlxVcNpCG0/bgFS+HKHI5zLGVkcVCjhMJ8fqIV91DNm/GKPPd+8EyjAIo2MhP
ZfLfEiiTZZSPH3c+97Z7iG8lMwdlBqxZYVDeVi0MMYRezgQp353SGpICrv5Ss+TwHhBSNzMRzkQQ
z2xchXyUyiferttKo632LMqM37YLSRs8Hl6HG9BpI7GHaCO8ix5Bo87RGIP5+c8yCj6uR3bzEr4r
NqamhnJXZUxqMzoEpyjqGK4rSqS4YH7daqK0KFAwhtKvP8HdVVBZM019EeCLa+WUNVlomb0zBb6t
fUN7IGn8XYJ1PU/6i6jpgmHFFwhIkgBJp4UlzS4Iqa6Bn2XSXtgMP22nZ/h+23K9nMeg2PBbg6Dg
9k2soT1t2QKnRBJbKt73Z4MzB8vzO/knqYsWSEewE2O/sdqw1jtODPNRHOCKUViRYWGejlR/9oZd
ngxTRTnrJN2ElwYgzw8Qyg622O+dB0pZt1vwc/HkLi2vxAvAvP13U33kgRXrjB8V5gFP7fxGaO3Z
EQ65IqpT9H8ZFn4mjzonUXZrGroIcOq/RCZdJm4oEkx4ytLrocYyycz/R6ASe3LCUcVUe8dSPpXD
xbRbYd/clIxsQPIkZJkdkcTbl37tKB4dKU/U0ssKMeumwvaqrV2MiSow8MMRLohAjPadeCK6tXu+
xnb7jPB89qB6bQ6dfW87HlcXuxwl+RXtyt8iWdWXhXgUQe4Y/8wKLeSmdLb5GY6aOTxe5fuWxdJ0
WxuKPLSRyJlpR7wxRMMmxWouxwJU6ofXCq5l7vh3xBe+Vft+o1MxTyK/aJPjK4O6kGs1JnDMGC2r
56L7XA5Vx5JdZtApG+Ql3JbWx2QnReWZNTVNawxQqMpeGcSPQlKu9GmI2N0BduSdARAXmexH+ghb
nhQ+DcBOXwdJ6GNinCT8a+/LpJNS9i4FmreJbSBIH9tcltMZb0142k2O8HVX2lwatSSz2GvpfcqP
veFMwiy58WTGEkCtbJf96ejd3rkxEVGep+qoz1Tr50I9H0m7jac0r1mkh2nxkuFMA0d4yLi4/nf5
nWK6si6Qo7xpRCKSrpz9pxLBbNT4kAw0XmD31Voglcfusee2pSsd+1kKcrYXeOsLFby/Rr+uWOb7
yphY7l5e+R4omFnlJSsvlhW7dTo5WT2w1R7wSqKH7mMtf/dGBezrkFWrhaTqGZnD76XGY+7SZSNS
QCLYqNpSAUr4Tm5bCtveR3fjUbBpC/N8xmS3ChAe7D8dJ3s57wnsrDK0dOzoEyKxens5SUR4ZLjy
8WsxBO2MUvLkCpFv0fYh6q+q/k7WjJN15PPrrocJmXch9qFK/90EojSRh2YeI/Lo08SyideBabZZ
/0Uvc1IuJw31LzG81ORs8vsBJJG2oeJLQlyBX4ySS5lRFxmzZ8VFrXk/ppL+Sp9LHkGuMKve3ReK
KVMXQ9pl/ADTVvIFoJRMx0kz+c1e+jqaDPiYQxAIy40JuT6vNTThrNbGlzk81S0ncXhBdCvlU4R7
HQUTDwtbABLwDKolA8gQrDzE/ZKsdp5nRZBlrnexQAuuPNGrBPYOXQXVxoCZc2u6K6P67vPlsau6
JUTMBUEhX78eXvi9qh6MsmpOmtlj0uoEpZti8Yqui22/j9WEp8pcSlNalsijzRObofjuOEBmJpT6
DkDJgHCrdl2WsWc8MONusAahKNtuEY82K3pRYs0BT0Phg+xi/4qDC4V+vQG5x6s1EacyveV00Qrg
guBSPLng8J7ybhVRa6aOCMlj76K5+4vBe++wM3P2r63micJtzcJY+fAp7X5n995GohLUC+UvYiTZ
+QyuFFUqTMygsGDeX7tS/ZR4T/Zr4QibXrta8oaSupRzV/mwTzNxq2VM+lPy3U7/lklGzqju1Bew
Z5cYMqST31EXgCMLI7sH+pi37Mys7AD1cwOKR0gTBJMEmv/2dM6pBtlWPFuGO2sVcg56W8+CjP16
WmtwIZMMmdNfJZnmkgfQBv40l0sNDYby1b3WrnE5RFQ72hXNPdawmGpYWBBcSz3RrhFjIm1E3F5e
tg1M1rAgq1bDLkqnNy7Tjm0K8IcbFJdXq3WoHMBL87F8yqvrxxpXOIi8R+L01vjHGJQS7AfEY+Vm
t+zp2vMRD8YsYWoaHAc+suKh7y7LakrqcYNeTTXKNMoFeiI5IL+Ebh6wq+veY1xu31Lo2oR5A5CY
2aulJfUZ2mz0fX/JyFwRV6nqe6iOF50PD6Q8mAC4UIC3IcbEyHRl3ddMkElspd2mLPLvrqcVjK60
G2iNZ5Xyd6RvsE0yI3qq7zT7ypVCegPy7MdZZOrywfABZbdra8637ZX2qdlN+CaINq0adHL3q4Kf
WKhUW7ckF77ZtbaxJ/13d7xCPoZTgVlUMRPjA8xc1VKw1kkZBqA7qE51eJQlhGTq7YHEGe0c+VrM
BOpOdwTAcTm+M9NMy2gldvEDTUMGxQrJiWD9ILUI+jnL31dnLQKM+EdGz3W0xUXXVA8wadg5fEkQ
nynA3McjFL2Xos8FYIXk7iXiOhxJ6vVEHbs9fB2hoY1TtRG1CgFw2rVhF/JEXu3vs8h6hWFhcN3w
dEMMcA/0+2Zp4CB2bAnZJMAvA6IuRHjbMa1kJt1kPcuemayc1uX3CXyR61W5GH7yAQ9TFVzdx2Jb
oLSFzBr64pc0kzpMmRnLKzvw4wwS9HTS6SmXmEj9Bd0ZxFd9pLaq5/9Bp7oI+kv7tkyU/t6BAxzI
/RLXuX1nV19PlrmLk2KyJq26cHzradlXgdDI4kHrUqFPffY2DMoc0NbYoI2sIRuqheSvYm9AC0Io
V8/TdBZ63zi7lF4IgaVC1nHNTf6mxkFDhPOPmBzJnxny5CgP4bqJyva8FFO9agLLOz7Rri7D/aMn
pFL8DWC0NrAo0GDg7nYc88iE7EpAQX6XIjIAO3zfb0bpNqkyWr+qEQ3X0l+MAPyoAgw/pfCEszTC
FRMFRK+TePDxKpsbfbSGPDvUyb01u3wlhhXygXWpYU7l5zKGwiIzsgAp5YhKVTT3DnSltE0b2SVK
uEVdHrqcga15HMjO0n3eVIfCeir7R9DKfE3uoczib3SZTvVbfmRwLo+ya71PoqH3a0yb+X+jEXKJ
tHfjkL1zoJ/52MTXsWwuiwcB2+FxwPZ5ADYS4qKJ6F3JD8qdn1GT7qiFSC/ZD+oBVHooQTc5fL0w
Rt6TI1rDO0GtacpDLeP+H8+YVMrZMdLNl4FEwzC0XvLDYCccg6TNyh8kP8LgVSWPK4zPIa69VtCP
/CYogv5Vx08YlYpAtAyhgrCOMl3/b6m3CP9QLZq1cxen9GEzbXCD0hF9Z0EDLHpc0h6xnO99jsIW
a4bcaJiWy1pjnPBVd1F1Y17eRWh9rcAN7hzJ+WgbCOl9ofFaKz1e6mTD2C0Kq45my86Baqe6MveL
IIm04filBNAu3q2tI/YSs9gj86ct4vNwkTXJPiEbrXLVWnrNyAuHgaHreHPgtZmBH3YeKTF+7KHa
4/XeeffQ8mSjYRo2L+X+L1PlmMoGC7SAq4ejC9jOBt3B53PHipRoX4iOQwNTpel+BBERURIEaU5P
w7mhYYGkutSyoBIvP/H0SSvw5VCmbP6zi6qh4cfwlAO9SbmkvuT/HJ1t9L2aoT9jIEhjhkiB2qRR
IixInUvwbD4yUgfuS0V886BHrjQSQr8z+hXAKvuLllRUmSUMt9JTl3PYDLsEPbU0injBViMI8DvW
nJgQzl2JNQmet9GUWLQQqmRV4vTJnv/ZJav8xFS+OPYfPZLZVdHFiUYXNyVFvgM4Dnkqlgk6vtoE
18SfQPN5kchbiEU4dDfkG4ZINCBvDYHpBLsc9bYiUxrZMq5K5XLtrOtc3D5o3lQMIp2aJbd6NQ3r
ZYCnTIdBcPZO4jh/Up0xQzEsnn52AQ7DSrOp4ccBoDjwn4oklr62jJ+JQ6qlZUnh0MwPsD048dt8
ngGFlC/U+7OYNfDrir4OEglARWV60uBDjC99H4KW7SIiMmvCc7CdGZMqAwjq82ZDpGcsrZRSerp4
iT/7XdowvahpiiGeIMjABGaqNh2Zcxq0VjUt2R0PvAAGCotVqukB0Su7uuJ3RDt/esz0o5C3Z+pj
xOuNEBBwEpOquwMjm2RqRtr6nTyBXh0ZqAcnEIKn41B18QueZj5E2f3zVNZc4ZwRXtWQPi5b3JyG
liyA/6M6oSZZBTmUoP1TJKN+NlSo9yeBrDghMqEdj8YHce78xmHHwWC3QqReuAPoeBudxmScQQjG
hxTQDt9AeDPMR9QJas66RGhZIS8SC6pYLk0ht1uYB8zQATI6ruWGW0wUzLmChWOw8Ag6DCr7Pzhn
sdqxMCxv9QOy0KBzIdHOoEnnCzd52Irm5iL9CHOSLw4HuOBwmlvhPexEHuDp2KFWK3Cob/MIRWJj
FGCAA+tXpQQxTFGaDECcA36AFqNdrmee1j7JCB8tWd3tm0b48lHHlDNI0NwOH4hM3Xp4JJNkDbi/
ewYU/dRppDk5ccFxpy4FDHdrM8PY/V1+U3Yx7VL65YlP597zwk2wftsLb5DP7jLM9+IPI/jTVQij
bh6F8qEpmQm4uW17HQ5PVKgHeiEtqTSzDuWE0nYUv6r4GJLecAQ53EJ+Oeklij9NHkwUGhbi4mKu
/EeW8laTcuSep0PKn6Kze8ErydimIJVN8NBi2xr0SR8+0hSEG1ezy7fCTfvCUW1e+2tojo+jeQxC
quPhgt7PbZxdomw/QV2+scLLq5paKKjQMJfa3G/Xs7zwJOweyyxvsJKJ1MjZaJhq4O72slGyvvzm
abFen6FOFEDwkoc3VUDzFfM7rAd9RlRG8mO9aVzVpsear+NVdek88G8/Sb9chic+A7tCP28QBKmC
V3a6uBFybm3DKwxmntgwu38El74CtwMm5wkeFLDzvC9v6hUSXBnczxMQVEF6X2qiBBA6bsO9go54
iTLlrpkAW/riQn0lSOrKT92X8oPYsIXOw3wLahlI8mnXqI2gADUzttcD6J7nvTGJb3LT8tQIc1/Z
9mZw070NFpUlpwyQklPV9xxFuJtbC7M27cjXNCdFmEtL+gXCRz4pdXlQoJa6pBhj1C4Xqfo/CxFR
Nk4osj0q6A9AC5HxhM+rw1K0+dfnNZdblOv6u8V6Rav/EVogdnke0f2EUp/mvkgyybWSlZL7He9S
FBiQ8FK5E8qL/NKO73FQ3JWQ7H7NKqJu1XdJlae/qPSWPKxVKhPEkwxZzPOxL/L+11IA/yW2i8RP
m8gegwfk0pwBBDs0vPPiQvSwYOOaAtprN72XYAV82qesAQvJK2RIuKmJxfz15gfdGLAQ57wBa1ZU
Tnpd99oe3mGhaF7vlkwE5NIA3aNkWnre8Se3SBiIESG859do9WGG2McWYGDXY3g8TMF0b1G8DaQv
35o/trL9mL7cREjWbdv55KayPHTT40iWOZRaF4HazzUlFC0EHct8ahNdtuSeK3pe7nlz2f4B1Mjt
/kuAojzonN/Bh+CK13U/+f+iVekt4IrN6jRu634Urrixfj1Np/iBLOw2wfsTDwrHbssyAmmqzY1h
LcuZNyNPUlZXuZnzl9+lSMMii7KMdXQxMFs/pbor7UIY0bVApbRrSsy+ELLBmVyf4TROxavv7kGt
uB+67xSiezBqe+17wJMicu6+Fv6+m8cSr1GxS4Gwz5S25Vms6aS/tVRQuHjcM+DsilXrhbu5XVMo
/Mh9ypa62Jy+ElZmHliZMobPLbf9sUPQvuIb7EtQWfXX4h4cOK8OYa9g2sPNvLlvEEvgdLgMs+DB
lgQgqG4HxEEp1r+T1H4gH2I5mcDTJJ/9LfB1IS57PjuAv2GwInhxbTg2jipuzyaSd/5GTLFPAsNN
kRe8hjohX77hRFqQRenKnSvonuqoc7EzK4AZyZL9cAyRMYUelbS7HdEX6FYiS33ERv3NcBYkdmS1
dangGp7xc1Wx+/TSESmL80UMLNgk3DPkFY48OdmFUTQKi6tVsdPZup2DhsEdeHQ4k2OjKxIOmqmo
Cq5R/diOBEFXgOWDqbfRx38oxvaGvmLaEQy8ssi1Boyx8o1g4TiY8BsCEgTtDnUqrV3v45iSO83t
NvMNOmEtc3npCJ3OFFAOUpOy2lBU/SVEfC/0zXdlSGlYwmP1iB9eV2JlLkaQqj0hA1CrngITT77J
RZiJVvCZ6FdqYAL3pPY8zLi05Ip4C3KrO88RrfCDx8KOqwzQYz/+sJ6SPjAi1ly+WwkybbCo7j3R
ByeAuQiVCrRj5CNykooA7LVNoqgBlIe2I6nLs5xyajU5cYHx4TtQOOvP24dZO8aXaOzHvMltH3SE
OnXHxUhcwy3X63fvNfoWey0rcQ4YNMkAiQqspg5xj3xk8/vflcRonBqh5hX0PsBy88X68ebh1QRP
bJ/Uv+oWgL1oK2/QDmgSqLCby/2Ij+kIfbPSptVO7/jT04S42r6RY8JZRuU/BNSKMegNTWwJsgBq
VzNSspEuCnhWYOLrbWotXSmcXmI0EmlhaQoT+3GhBinhV/LBw27K5ohrEif7GAJdJPNp2uj+3mrk
GLb60/xtsT6djelWC3k3qcTjqPEC6oCSs9VIHiSEhA+I2+l7ZE8kes+jQfMbH72MoBwasxoyWaYm
LTmRrRNuOKtVqkgGQ3S8zKEHi3i2x2+xNW6ALlpsWrfTYBZDhsk6FP0zgQVBQY5W97x2qGLfAynO
IE4/CEAKMxWqOXy6PR+YChOGGk3N3G/ij/4xG1y9JAxg2T67g/+ZE8Tr3nKJb8SeFv3NC6ls4Z7J
30aeqxyV9XzpVTJ/5RfkEd7Ofb7BFY7vcpL39hT5MBKF1unDieibEpswmeyctSh2JZ4Fgk+/P7aB
yDXviccgUlzrIRLX8RKlPcPVdAT23WZ/M+X6kiWjdfCK8nw0yktMMsHKb4wvDfr+C+oN07fuT5cn
hZi+EJF3URWMTGm9boS/0HEn9PfR4zTyYsOXuvRU3i6qVK0VYSe0bblV138Up5S8RnwU74mz6eex
0UOClGtHj0cRI1dLWInt9q+JWT4wJM3tqSq6OPXHiDtVy8xVUcVszXyzIjx7Eh0lNnPteBNtKDz1
jKnbiQld89W2gCCtGwQ8kZ23QIcZ7IGg0HpkjHH39zzRw0vlWgE5gtRygM/Dpj8oJvJgWQB8mQ4/
QaJrmUqTvIzLHN2pecWwI0CU4NQlSJaPhMT+biWyDyXkZysFiiYfasyCDBGceXAQJRb18c353GkG
1C/nlkSKQLGBQ2YA7g6KAii1LTmaUHdvrsTG606uL3sQQcY2PDMD7kI9VYJ4RQ63ebIe28Et1RGd
Dd37PtaNMEApn+sp8jWANyW2b9hCmQFU582kAhcLIfAqEZIKSGWirbAMRPsx00fcU+1Sjp14wWXY
m+dtc3vq5GUbob5fkX9a8WfYC9CfvMIzG5M+SRH/QG5X9PZgfIRr5RxPruxM1Xc2ABFPunuRzAIz
MYQIm5mBQbiyHqRoz6Xv5gdBLXCeD4jDKPflpOFKNXZiv9OyJKUjKj8L7OFMfOvqAlSJjijjOJ2l
eeXbwHADua4Ne7KcTgrC4MPPrFNfEZAHP2APzmM2/tby7c9rlfL0TVKM/dAiJpi4rYhuVhNLeHSn
wZCALUKFPsZF5q9cs6EzjrFHdCpRf+vO9X41WQC5uoxRMjqUEJvH9NNT92G63fgQ4WcileLl4pcV
1eLTVXVoOO3W1vmIaqpQK7KxZSzIbetaiiIOZOnD/qBFkVwoSdr5/IBySGmuH2OkDg6YrgbDVthc
KDbfBh0J0Rr8+NFX+/HH5DwJydIwrR7OOaO541YAdTbNGTlvTWhDE11PBvLWxrCoJXQJzvUJ2sEa
aXdCQhq+tLOdWZk0zrAmfd9qHH7Hk4pdhGVqNZaJ9ndNvIaEPnGm7MT4UP1FcYgVwJOfzVGpHCdJ
w1Aa6gvn8h2azXueKlBNgrSkH6XzDkBstzvqo9/wnLqI3Tgtg9rz2f99vRPbdvStB2eeCFV2/KHd
Ho9hCkTs74PjnRj5wvg8h7h1HfAGERbl9xBlE848QwQzdA6WmP40XRrJMx2yygggdQE3RMI/EwJ8
AmgFiDDyTv4GyQ+M5DX/wn13NvkJx+VVSb3/E2cjpIa5v+vDt+XsgOJPAgwMiLD+05Zd9jGtxKX8
bm06B7Y5ZCoFt28Pk86VhnDOHs1sJBULJ+m82wgEsHrBAvIrouociNHINaJF9z/rwoSlkzou88RS
kNUdXe3BnKDtMLinC/y85VYufUEXHn7QsM0LoROweHW2EXPqGvHVpM4Odfzti+oU7fQz3UNCXBLm
mW3Kcug3Y245ZrcxiTatBvIpTwW5ZJ2xD9s2F7W1o3/UX8tp23OUhTE8v6ossJyrQIkrSs/RzTUa
/owie7QmYiTM8gdqaILQffLQr7AA4qp0kFAFe7heBF61aqKHzPvNrsfRTVTpOqOulRgA2sBs2t4c
cXkLmCat7+uPtyu1Rdp5e0o9N9jRUSLSBKEo3naiNJ68r9SbCQa8f3gv+c8GFkfxpeC7GtGHPQK5
SOsm/sIEby2qilIgL0nMZMRK6bxKONnW29ZwBGCCDy9P/16LqcdUXNc9Qx8WwbfL6kyJj/rXXD2F
oyhgUyeRm5QzHOQr+hF9/hOByV5yFYyDAxU3AhdP0Xe+LaoRnqAPGS1m8L2UY8mSUSPYixMamTxe
9lmYwyyIg4kMoe8dlv4Ya8TDNdxGuSSTChnT7Jp0wtCHuqQ3kbZI+fjkCeeJ4EJWsndLr1hf8v3J
MddNkRLX3KITD5zVT0m0+i2sK9nyWHSrzmGBQNaY575E75GeORFIhP/y7laJVHP+OpD53cCvoYz0
+1JB8xOlspSNooWGaFy0beGajEEwhz9b9Iu+pcE2ml50kfYzwrQiGTfl38v/4wbJChSodH7a5urD
yvl/jwxCuobpYAbHQme0ce8VzFfFEXDOA+1GmEwFKCbipI/ofkdMhFt6OpK6DT9mdhBeXv+eQwRG
D1Hq4SuOoEO9GmF5fWKUdSyzoOSwao6umhT9aPyVx94/Zpa7MK3mijSt864haRoOreLiFJ/yWrXi
FN4bcGI8TxtHDInqx9oDbe32ylX3S5giqBfC+lld5VmoVpirgpX0RRPwKEk21lCvH40uUgGtUX3+
FhXwCunbRYrdZHxDNjKC9SEcoCYy9jeO5cg7Zx3Y4IPGyOC/cFoSCs6YRlTJvFQNePkWZRC/zpZp
WathwYNfpqSu0n1IGadlwl36g8ZFOWo9jyxBZldy7/Mz4wdesFIKSDd5uM3I7AEJuMkawkF+Z+4j
dpozP7dOISW8mg9ppTzIdMJv8oSVPakLN5lFlpU7sXjLamqQEyCOLN8h9Iea/eeG1AH2e9VSp90z
q4KP3leK8iJBn23yOP+WJqRrsEa8Hi5WKY80qj83ERutdiLn0PAXSS4VQIc3viHLah5FW0rxtpTm
zOk4SsCi57gJPk2OLrtwKB/433zETssns3V2lkGtjZcRXtKDgfiMbstPhAExzbcFXwDtRXllwSdq
7mOlf5E45tuSEcI6/0bKpjtNDuy+waSVcATjhOaSieXhzfK/nHyJs7lOdmWpxjMrAAwP8jKqUrIh
DlrUSiTp7vIJiqcqzZCAnFEhhaewCak4fRiu1v6T+OPgRTk2WIeZHRKui2ZwznDivkI8NUbNzvou
nMe6D8Y9B+uCspq7RW912W7Jnnpe24xRKNhkybqsXyUIDTzNi1CBgAZyxBdwBpEZXgocC+SsgmLD
X/gMo6ofTnXZdmjigpwXd+ihvNhj1k9uiZaQmY7rLwU2Cku1OizyqHx9ZLeNO7kka1v0Qvx+o0bc
Ud+lcRMPnVxBeG/S7EdAVyp5XUM74JjOsThng7nQlcAKl1ekPhmypKeiUrYN0tSae2ZVrlIzWair
B8p3DC+8dBH+GTMNYRQhutnxCN7sR3UuJvyugBNcihAxAPYcNBdMthY+DycEBoZtvAK+TTdgvh3H
JJu8Po9xRd03egC/Xn9XQeJ4T9gJj7IfFYr8HJSIjNFTr0jloAVBhql096vENDQyXuefidE/mrht
UfLtmd6SEGkh40nOQU4fLCir43SXCWlj0/CS8QUC7+kmLHr87hr8OGUSszXeUNCYLiNxRHmWJNuc
PznYK/U1HuoK66JVN3mxI5gG6CelcXIGhJH/Wxa9Ey0+xiZLM8raoFUv2g+ZxAPzS3oNN7FZx5+A
Fh/moa+vAxnND7tpVTXihkmCJtyOSeiSeNjZZCoAXIl22uqURKWrzntBvx3sYLFdDqcuOJOxjkXL
KGIKv/Yu/C/I9KbeDIrzLcE8SSVc8XkpOtdS2Pw6bFh0RwCe6iFtMPfpC85KhzhODhVrR8OQQm/R
cnoSBne29nZ+Wg1hJrAg0tA+FEp9ZGDPurKvpzMLIBu54OWazHQIP3vrssk/4vBv7CIxsfirX74S
51bRLq5jKsLwrcUVAPcqYFXI+gJ0I5Vfn4QbDxxO538k7/Gf63quSEpfCjIZ4fA+W4UmpgxRQEIp
Vc6IzJ1+BtGIhY7AK/EXC+XUPZ9Uz6oZ/Tp+99JkxTrGnTjc3m8jkxm6uKYzrzzat1O+wwNbw5Mp
Tmsd5MomUyaVt1+7beC1F4nerGUw+9Tb0Ohkenvg3o2vG30h9w8RdmH19lHq1QgRawoI4FJPHr3S
+jkG9JQdPQGfcLgM2Jjs1a1WfNrEIWn1XwJY0mu96eqWCjIe2+1PXBwIpOiRDWF/SKu2K4ZDb7Ur
owfgL/Hi9Kg6N1dJLfdI48ABknQDoDg8iz0I7btygRmrH8YUB6rbyHh1CbvHgB0xC6yEVnVxc0vU
Rv57hR8678lY+hPmQM0KMzoUyLJQWa41ND3guX0OVQfv8+7SwTS5c2buICEXE4sUjnp7tZxWRQff
B/4R8qiEuLEh/dgQCoG65KIOGd6Mbd+wtZ3EnAU393eqEehDh48zO1jKWjBYk7jRWFm5MfxqQbLb
oU9kZK05+46fodhXBDXKETk7hyFc1Z++/+DQUDLutIzSj2znLS8iL9cCU/0IzJZykhDAbQ01RguG
gg4LtyeO2Cgvj3LG94mJ+vAcAqDBqHqRjSQTdYlzmbjymCGHeUKxobcPh5PFQhctYbsRpY4/HWcc
hJ1TiHeJu+pCG/BqAjbQdepLaWKjS/GuQow0cdtxBM5HdP5SotZTMKCdj1Dcfj4+9wWh5Kd7xGsQ
pbb0XsfurSJ7vgwNodcVxtf0pBmMRb+lMpQSLHNmzjpe8CshSfoMQM4DZWwFyH1LkCduD0CZHlho
JSFtylukp7Ac03CQ1S5KYgQUF5BS7bBkqxN5X/DZxDileyTikqZfYvGDqRS3VZb0dsQEopjrU5x7
fQ2Q7YHPh38LxWRsR9mWvHOijVAhAszhmgUXEzhtqIQv/lUBJTfgbWtC35JDYESFNyKbOuKVnD68
Mqy5oUwOK5Jlohgg7BZD9wu/BdA6yvTf/GdM8zoB3jU3Y7Q3wnR9oLHYItBPBGn52BOz2QLFnBTp
F+KZSTXz0w2UKxliWKphUOPAUpWBFJ4tcgF+eujbrXHgnm1n37oujoWJJQbPOIqUHgYnOkPCABu2
DfIXho9foIzO4fFZk6VqxRKqFFf5WIxaz3ZP/9/c1Hi3APxzmWbc4m9f+63KNyeeWdpWkjG5R12X
NA0+QTH8Fk1+z1yTj/92KH03ubJ7ISEzFOLXN0iecLVkUoe0U0Mg6WxgxGbDN4iUREntFTnkveAp
r/bCKYtWz1yQmr+vlJqSAMtzO0wOz0saoMPs/GACT1vn6MMPvDvz04I3giMUebXRg6CTBycwPCUp
L8rXwkhFQNArojAsFbFYqJkovoA8ngVx5Sl0GKucH61O0bzsd1A7vZtPi039JnylMzll3lAfE/tp
CoFWm+xIwr2QOSJ4/5SiY7/av5VDD8evf3i0OSzIhq72djjXgkZnA7PlrSoVCHmzxCgq260Qxqay
6HkxWWkj+3frM6nfKWh8yyRTmYNzUnrCnU8xnEA/zHwyUvMkaQhIxNcmNaZgJrBe/4GJyY0cF3I2
DzKKT/95WkZwqIitB8W36+cwjk960wkyMnLdROMtaY6/xWaIH6C6SPbn1NDzvxcTa1PxVX8qrmup
vq/e31svuUF0v5Esk37m/DNw93giOf4k3PIyO5Nq5hOkMRQ/z52UVJAiz0ObhZCQfo2k4yuCy2me
+jM0qJht/CzdIDFoBNxK0eKpI/XoOAXBMWQ11rQ4weyEEauHRy/uWx42fctd4Fap2Exv9q+T1SLS
mWVPj/RjFNUWQ+eDXjuKQgJJgQklZ4T80L2pPnLawFk3AG8QorCuKWobMkGK6wd8qFARpvtacuSr
uOF/GMEjkeA/JLSRWxQ+QgPQMT88HkV1zqhm8zO3n4w/EZ8411BooQ0FvHnf5l26o4BosAvEe2Wh
/TwI/GD3+m0yzo9ocw7ofQqVg2nolj78lfOVcVg3iYMLPIp/1N8IjiqWZJ/WI0P6nHDAt2tS+Ew7
iXs5ulY/bsR3/WBlE4PhqBUN+4quXciZN3bIygCgOPtxeAFyY9Y/QxvYYtlFEgHBeLj4aLuplpp5
UDt2otiwpO4UVZHcoAmLvH1TJrSMBAzJpLKWzfLC5sg18dK6PKbEXkU9BhiXygKQrUG65s/sVqOd
xEaeyagRgL46hbd0UpPvlXN3NknXAkfeiKTrsNeUkZFBvYX+PfgrIz4XS7049qiihPb8JGR0O2if
yGo2vlk9sE96HwKrXCW6tYresAyljjMOwzQd87LhWJl0g1mo+KGbAYray+UvNzcmKZK+dSuQ77Eq
S+TPmpLTx2ko1oUIPGQNA+0ygbx/7EAbqD+p1BKJHdPfetj8wvwCmHy96uBV4mXuq903vrx9zkJf
oZQBxtNOf9HB3D8lsSXcItkqxX+np1K8y+rj0v21Pc4ohzFpgX3EJKUyAxmKZRv4156mhGWan164
iEvwjxSRkOf3aIYQ2lIwv8piHv6sR7bDSkNlK0HAtihMp+SK/oG5B/FwX8xELxxNJtb5xKgsmPlp
66xsOH6rShGuZ8gQIBQyvFG5hb9wWsBM8ve2KQgX2MkAZOWb/XbwNRq/zsnbkz5ySxDCfYpQYYB8
eXxMbppebUToKygLaEpTIqLwFn2zk4s2mRbttF275lQPfACcRVtM7rCmN7ozy88kEwLoRbryv5zl
aOlfy5PWciAbP3e4FPut9+kC7qqfuN6uFqKLUMTLKcmuZgIcLjm7Kfih+xS5248sA9tFWqW0eDL+
to8JdZNrUoAMfO4mlKPnRR8sDYqAdCTc2WfIsEVzCVzEmENwRz9EaU9IKEjCpC1nnuPdnRjaWIjc
jOnRZYIinQjefuFZsKxoJQM9BMgY6NGmvC1lei/5KIrW6P/9Ti+W/onRA55Ri6kjyFm6a1osg7YZ
29bmQm6utQzW5/6WyIj/BWXx3COACrZ/nu4giUailbcS/ncrKdVv6FK+ccapVzCS9Q+st0e/+5oz
Rv/QZ0CqK1N4J7hq2TBVhn2FtWnLPATKB2ZA2DdfJlePyGW9eS5EQUaeNffZE+nWDgCrH1dT+j4D
dMbZRwG63bkam87qZZLAj3MkqeaN0tsIFK2eHm9oZpJHiPqv67Mk4ieTKi/E8XJyyCuiEZfvGToq
E7AUPrCamGzL2feM3d9m8Zb32Of4vjzTZWVBasBsKgxkGDG0r3nuQKugqhnKFtfFl5hoY89GPjLg
CHgKq4nuinMDz09L2+YpBQwuxN+Kj6d9gApT+372J0ctvqtd4NgtZj0jy/XSMckBJLH4UqdZWwAp
ZgOuSsezoUAkTcDZxm9PG8OlpTdTkMac2u7Oqre+CbhuJfLn4UoNOkv+zLk+puTWIggMmeXrRKta
J30pomt61mZow3p/oFBEMdHvBMdMlJPWlbpnKUquTcPoyy/U5ztHAlx7gbnly56YOHhyFFCYKIo4
Cn5xRwi1vF8rDbuylMfsnfquMbMH2rCsIFPHNHVSN35lvLoWRytATqybYZ6eHOVybnGGf4kdJzrF
FTozttJDFTQK6+EQrIuC16iIh9kXWK6B4ChxUds9iwxDAyVjwVWXTX6SiBTEhvYaMceZbV9xvcCi
riB8GCjN95je9eoW5nCbXfZ+g/J4XN2DbLa11zVUOWDfm/xNVBOlnVuQG0mcODUN3uBtxNDclQCZ
lmAKptB0WeDJSX3CcLeyZL0QgWQdO972ci9NuC5Z0KYQzp/rYQBd0kN4GnaX2juxhEf+SQ2jZiEh
ZGdfPlWWuXYhq4EAxXgn3X7pmjDtIMFznfXmNf16ciOliKvMHZkXa1qH4PoZSDLQC9GPOz/TEF8r
v5I9/3kXX87JRm30oEPgW0Q99yMS/DD7JptMb+WJdiADj04IQ1i52OUFbL5Wd4TsxEdMt6yhZ0jH
7qlsp7TBngQo1xOw8oeU5mKbHT3Zvv0xRmnKK+NmhpdVle40x+7MdT9KGjHByLUdUD9GdL0S/2p6
UTEiyHRAgFnMD8xAVYnpZ8aOVJLZlBxpCwodiMTc9B2fOTAR2SdrKhY7hBk7Nsr06DbOnontbz4G
e7wK7rUw2R9/XLiG5EctEJSGlFB2p256ijMoSmcJqURe1nhkXyVB1/5HBd97jtZTnKLwaKbKUDi6
9cYUSija0LX5XjF6aamC2LD+iFrqXo1T/luJHP3+ZKFgW14+O3adozAnfWznqFDM36rOnbvWEpkP
V5V4mbGXz8q+VNGzEBCJwnHX9N9Rgi2yYIFiGNDQ8pRgobw1kgmRMHxmytOF89D5WaGSoFkMOObx
wsiHL/t4LkLy73ZRBeRq2xYVq0U6NkQ8WFtMkyBr84SGyXqIM+8Zyp2baPhZGLveaxO+bJXOKFI4
fRNifOV/v5K19TDViMmLgJXcKODCRtfHKNbAgGXSaGFX3ptmTqCYBE5RNNlJcYiDq9zNTH4mqe0h
9PrXKCVpBmwLDD9GhOPZw0nFImAgyAqjRgC8VlRPqa/hbJTsZUW2r7MiwPM5pPuPtkm1UrQ4Ew+a
E40k03RY6iIi6hTGSYkr5O2bONGBWmruALKoS27ostsEyFAauxiZsBu/YLz8ZEVrx+O9oEThh2cL
dqbP7MebOyltJ3xMrHJ+PsnQtTjehhRb2N28rjy198tYEONrNzxwFCQHrdM8LNo0qO8Q/trgtdnw
XhNGS9klfMyevnYKjwPP5znK5rIAy3siUYzFP5qBYWfvBEPkLNbtWih1yhxgRyRcdWfRpu2puA3+
GNlUb8MU+mfsFANCECrx831xkrFMAC/iWQ5O7TZx/c8SvKzE6vAyFYOLiDHLgHcRO0qNrcZLPFaW
5TUaHHH9d798DOfTlgXiZ9PL6pUSUVslZPjKzvporV3kIofCfF4r1k0rlSKVSOjAuI849zVH697y
x8/s3gxtn847gkXUdUyT1HJx19qH9F3/uZNl7c/kzpTuev0OhirxnJbbyhQoBAxBBThoXVW5h87K
kbtakQCFgSqpIXvhepjt4MvlcOD0IYzWS+jNp1BEIMk3iXSwCueoEf5I+A1pYPH1eSrOtybALqNs
gmMkvLPb6Wj7yCKqrRxF2UvJ6w1nUAhCJC3HeG/mNj23kihBNacknfezu02izDDF4NKrFf4iuq1C
fASd186pxhkKpswTfj9CWrvp7VhXRrGjpL0Fxu9frXJdNsqsSdHwkXMoUo4KqwCRKOB9fnbwqsd7
FQXyXM3Gai7Y8wdhrvfSksf0XzYlhxf9rUbTp4druC9ISqbNig8wlc6bew3FXpRkryLlbjnlolBA
NBvhNnt3uwq31qRMYDfqetC1cPDe2o6dOb3C8q1v5useHrq+GNWNdahv1XDhNvwROe3Rp06QxZN4
V3ZvtAwYaDJwc4rS8eg2RrHZQr34qwo1TPsCU5YWx5Zv9TYuG37BMSOOU9aBYD40bEeYprANpd2S
fXWmsY8Zxd3cSqai7mbKp0J1FZ15Um2dSWdh8FUzZlOAzFCyX5Q6alXaUzAzMLIAuX69lQSlBWH3
28JcT9Hbwxk4PGJkgZkjlHmq64KQ0gDNRM6B7tuKMcYzjxMJ/PAwHoQ6FwBWx5JwdqN8fLWHmmv8
TpuG5oGMUewfQ4Bp9zjM3kyXNPzfUlcVJh7+DcDxN6lYEwjy2HpFHvGgWUSwYrfWdQRiN+Mr3bHo
/rk4rHogkmFmso7l0nq4V7e/WAc/NkIPdNMvpUhMDg/JUIfIVfN8ls4vSzRe+VlizA0aRvQaUU84
0iGxQ+J4wTdQTwNz0v5JF3D6d5qghUtpFvOXVrsqhsfu0VccDAThw2WI8N6Jd28DL/XbFiRtPkOT
4NM4AMnO3hP/NB1zj59yVDUkER2jA6/LvOZDshP+bqIhoZQiphUD+/6x0AjcAzVXILic1UIUrRGh
NcjHPmfBmZj6UwR89RviAkI70aKzNw4dFYMK6Np6US1J99ka0sUz6R5cdKwXyhgOn883P7IpN2o6
QPvgxqZvv8htvEWtkZ/J4N0cuCUpkrMDvozpnsfjDVFcs3zH+KXJDPBjPmuOx6FoCobuxue2q4sb
yrnMRLltbxbH3ZtsCJfZcdaUYBwJMF4O0e/wMVLRPPBXSjDfalBNnrepdPfYRG2rzBw2DFkYtiX6
F6ZdSJejYqdZnqjA6vPD1DvA3M+4D9P+mdoloeJsHJRnH6HrgjvRmpt6CkTxNeS0zw+iZBcMPLri
QQrsn6Xvqc9PxhyB1uhH6DCKuLzWqwxtPYkAESDr49ZS6cfqjtI1NgbZP8vymnoglHO86eRpXIBL
KFZXVh8SR0HOYA70sE/BDuqTl3t1+rcsDoLpKSVKiPFWIcUofGgDw7st8GDaB+oA+ZUq+RiAEU7m
C9oxSIaqjvNurmxiNGg4yHWatYEovSVrV9WtY6LsXX/WcKH7oTXRBYmXvlkxntitKrHVJTTxlf3d
lu+KwOBgHFxEtqoOR3MR9lI/MFb7w466HvXx572k20QrDQzIFKV3UK17yNcEVf4uvkIiL6PzACcP
qy9QxOGztQYy8hZlqGM2lg4tQcDfQIlqmOWAJlgIGt4TdnRobZhWg7oMA4pVcZGtKZBoD9WJUBy4
Et2eHHZHOvIqoUyzvVwBtP9iBZuViwrVWi92fvfyeA5jZ/nbQ5/PuaymtC9WZ06z+kjN8vgKHLGc
w7+q7hKdA0ODrIQs5UaGHhkRzq4dJu8TglnKAPkAoMceQPh794QYuH0h0oYMu8P/qlhk7D6cdmrx
umkjjvge9eSlDnNAJnI5cWZ7Xp0ESfnZYNfb8RCTn/ev24YqpEpfsrTycgwT9LlH+1IXpzTLyiWX
TL0WZee768NC4wBpgWuKXv780FW4GUJE5dEzzQgsVk0blB3qQko1exYHJTarPQtiQPKRLyTVJUcZ
nukbzQshShhXj7y8lmDKBGyGNSlPCpu81mzeN/ZMs+6ZSR39SeZrjlNgTTwAd2R7JKyTphwnjcIC
VDtk+wld+hd0bIoKUkdt3Pt3jna78j2MZ9KWOYs2n9eyGIKsZGzAIhdn0Tel6CQunvdaaQTFAN+m
oU6kRfsiMeCpCxKOX3WsB9VODLSyhRMKQ1VFgCZwgrTqZYcWczQ9PPJ23ODQxZ8F7q1PwqnmFp+5
fUQaLb5Hxpdw2zq0mcIHfxx9Imlr7ygtHek692Wbddg2CoT+0cnyeibN+zeqSSLWYGW9klUrn46B
AgVXZwMPh71iJ99nvgvMuKxtfM9ZkedAHkS68lfA5Sm2sZVdm4eZ9nemanAmUhNZip1UDDsPIDL1
P4G/z3srfmjybL8pYqplms+OR5by5/Q8AfN7JrD3nRwbtDvd+fZtjXduy0PfXpD9rM7wUeF4wXnS
5kKqh6GTCFVsb/j5VoJLNBpE9Px0OajBUpRr7hxREzabuMprPWY8IHQIae3Wdr9yKWksj2EqXmK+
yiXp3t2IGSnoB16s3pYGbw/NCxspoJtkCen+4saGPnWU7cnpSf8twUMepGvD12q4qG+F1/rYAYm8
hUBmE+yEJjkQ+mS08geZP+SE1LdXMR/ULr7aO3wVKBImTk5rz7zeD30HAx0aQDVGDLilqelSS7S2
9PoObWiwO3Hr6i1qJyKHQ4WTcSqmAULTliY44uF+mBoFcs+Ho7eHKBALwz7sk6PXal48XRVN4PC0
Y2SaMRTTYeKeXBhkfYUNjRbG3m6POlKJu2q84JJHleiaCsINmZTIJYr2zWUHSx803TFlbjGEgZYd
2785GVsI+aFT9hxb47Iu1g5IFMOvKQgCF0RJuMV+u58WPexYMTtpFtPsjS6dnHiHVtYhljNq0VJb
0kIsFUSa62eJnyWG92BKkPRggci4ykIGY8cmU8pNgchwvng6MlrTzkGPAasmY7/e1iEM4V1LAbJK
IufoRNBlZjd4Tso0jnsnURXGvCAYTU2paTIsYqQorLIBX78SYdPa934Ik7yfGS1EHlGzkPB8ra7F
0Xm4jD8xDy4AFrBRaSeQXT0Ol0iyPgbJ/JrfSOV5/eIPM7qGfo4fe9HDegVcNKPXMkpaP5fDFo4f
9n1aWwVrURVTN2f0k3U+KBhalgjyBEqgpmGhd6JTqVCi/BXEhYZ4PQ+Jgr13jxKNC4HWV9la0CvD
rUlg8nwRJkbvivE4ZwjWZR61c/OyducA1BgWiEPgTBc53eXOJwIM9mTknvx+h1UJVoXCigTzpBIp
9d8G8w8bzzPobTechevKBgTqFnBFaLlV1mtGLn9Cx7y0vIjXTbteIU8miav09zO5ZWnj8Eghd/+9
5+CFtmXGGRbBG5fGS/d1+fsEqpbXjbR6QP4xZe/bWHBX+7SOq9ForqziXrX1emf2GBianLQZkJon
U4rZtuPrut+wNHp9Azj8Qa9n/VYM+MnNwV9omgToyDx+A8e0gNMTHCQsMjp1w7tcFik4/dITp6pS
4IvVroEhs9+Sn2bjgUzfVANtjZNJAI/kHKBA0LreHO5nyL8jaXClyszCLW4i9kkWiY3/Vl06UNGU
6Q1BCWyI3M5s3DdFlRSQbTpj8BiWcN3FNRkRmJZ7M+A1Gq+ToQihE0mzj661atK388c+BCMZhZaL
aHfAD3apf26mVEj+Kt3+uqhnU3z7zqkgqDLbrQb2PaAQjkS8jIuFohjDPHw46qvAE0DL40S0YrB7
ukBYz9H837yK3xTrmEhezsb2QhbxYsgaf0HaRez2SK4CwvKdatpX3no8Jtd4NAsDUCgB0wovmz0Z
YW0uGy9CohF+GxUPRrUc0ioFdhS8dw+7kMKR/g0IDiK6ov5zO3zgflKSiLJDAq+359RhS+Wv0Alx
Ey1gd7eFcsOa0CraHhYjAdVhVn3rp+rUmguMMRadKst9gerKxQbgCta5bsD87c6EEG49QH1gQjaF
8gcUrmS5+VhJsTIMyMaO+3bscHeBu3UQNnFXhN9zgFI4vMc88FUVwtyGCHmTL5edcx3y6xcA61yp
DxiyuLecaUEwEiyuaugTVPVgn632dT9OHqzUuAZeQtcKd5camgK4vLI5AcQk+Q+rnszSm0xW8rH+
IlZLCLaKB6SG/n7ZE26k6+3EfSsMHF2jUbtdkvVYBRVjGHc3TjYRNoOE2GsPytOUXKUZzsr3kFE+
s5fsvpXljFKeD0iotzZQ7mG0Si4YDjE7mFO22aku2T/3UY4RzplGlTEqNyD8MEPRS4UPmZBanPfd
SLXiFFA/jFa6NxZ6sxHctFYHiE3cTigEeL/2GwccZ2/mWHeB8EBU9n99QMqzE+KiCBNf5vqaX9T8
59CB7ak6piNXG390MrANbdkoZOXDrhahd7gJOqFWtAqEF6hg5Ijw5is/z6GQmfKu2+g37PLlrNYC
kn9ydY+0ORYqiffcQ1CL/9an1N1ReQe7+V+2l/LSg+RoaMElvWZQyiKOGwC7OOS12Dkmb//9mHzu
dvPIG4l6r1eH7BAU0Nzm8g8sC1ONWYcklomMrlI0ghncdTBw2Lowdqm4GH0vsgPTNMiRM5GX0Q8s
KDRhjir7wzqcquo2t79NQ8AWZk4UhcyvA4mpaDXsMyY1Jbb8/E+aIItDs3Fj4XX2UdrgDSVn33zn
Z45any6rxXjLQKUWTrS+U4wiS9+0hgb+wiBLVTTIC0E2yAfJG+E7z2AX/Z/DeDctNDKAvVqZlqA/
QrKMNSZyACImeMe6QSXafxn3sp7R5DrsSf4c0qm5Ses+YC29TtYSnq4clr60Db4gxTGoaQYF6x98
Sbno588K/JG3aR2aMKSZcGgGfUrIUhAaQbBe+IUrgOY0/1M79DQL8mdoALCOKypM8xR93Z2pYCIb
HQmEdN5IXoF2/cIo9633VTUd93XePVHBxA9pPRKovfoyrv7lAip2PqHCC+1eknN7ZOv2l6Tum5i/
2APJjcnxkD5qQ209Ly2ZR5/yqp2PVWzvzz4bZPi5dJnvx0Ks57l8wGKKz5V5OfKDE9EboWMGrCVf
3F8n9XVeYf5hfPcyAG1MpGCHWBR5Mu5syOtH4whwPQgn8Xz5caV89hG6I7cSCnK1oc+fh8hZKGj7
5Mft8icXS+Xc0guijql+jmUjqY4QiMrVYjetkmJaX4YUJ337ycCzntW7vrQoCsL+0LoBXQS7xqvO
A2G6uZ1zDq8mZcZW9ZB6vO9KOtHE6vwa3FkAY10NZ2sk/qp0mX46dckqpMfxNpvJIElgQdP10XUn
/HPa385vbCdQYQXXIc/xfri+S0WyyYo6fWtK/4pS2X4yKnbrm0lv7xCXsIo6LnENgTfqcpbZn4yM
C+mgTp1Gw9ExdIxL83IrMIqrM6mqOA8JyOFW0KWkOcRJoS3HS/M4SZHD+4GEqrahMsPDjdWkfNfK
15TXPZsXATb9uTISk51EVXth2SU6cP0we7EmrNgWVVe9Xw/EbDiY9Vn8bBOKq3qEpMEx/wSHwLcP
uWapwgjVEZR+pqDdPSYWk+DG3ApSJu8nKX2MN/YsKnnQc8JMJ6k7Qwrfc4bPq+L7xiTn37V5gjic
TxcPJFKnPycou3zVicfAjFji3z4Sq68BU2VhxMMBwHuXA0S4gfDPEy4r1Ma12Vmn55YbInJK5I96
ZWHpp1JHyNYK5xbxl4D56E3N53UUGW5SIy0xyqDPejdAL/wyuU6kTkeuxgZeYBvzmt/w8P+y1G0Q
qXnptBNa62+VUTgTW2lrL8VZ1+C5JSZFNZlv0uA74gjN7IxiheOMEnu1pOmdPTBBcvHPAVX3o+MR
SGles0ia3RIA2nDY6hppbY/50tpvkxAmc0IwYe5gHQ7YsTtIoRL9TNdne2pIjot8NBReeE7tbee/
UtfxRttaiqSeIdL98f0cOLHdsH6LjM9DGHilL7Zxj1qNA0Zyac4h0qGIVw6nBQqlm1sX/GNB4iV7
m9PBdXr/i/sNHvX17FYZpfTEv4oOTA9S2P9vGlRPpBOr9nMnfMdagYzozG6vowp/ID2cuZNB1dYt
O5qQRYFvc/plpTEOXmXWxg3J900vHfJYVGIMy+BOFZhZll+SyM7x4o/m1QFw1qdvSjbnm7lgD8cl
Ca3pF4k9PjySvzWBfQSxmgbrEfthgINxpcTDHRp2+t41S7IMm7fyr03t08qTlrlCcW8nDxsJtoWi
nQTx45de+FXvAUpnkxn5PczE8t4130wcF0dHUJgBrpXxBpP2w+h1znur/aetDXNbr1CYy+Nnuppc
AVYqtb/BD1TLKFKoFfhA09E52dV4OmGZhB4f1CIcWuxys5WTyx0a3o6iaY8XDJSM6+Lb5BV/QlBh
URM/xV3ipc+ca92l8Z+NxXfFsPzAxo/6QKQKhk3aGxSvz4GtclHxwP/Hrhe43xKmDzz8+VmLCq/l
xcPbouxHhaD3iNVyZaUfCgOtxUTB0pqvMISmt/HkMSY+OotApq2OGSE9FvPF071PYD56pr/ylOfn
Z4ZNiPGO3Owwkw1NXqDqRQFb3RkfaZSqmKP1KzhDyVcviQB66MInI6jxPrw5KUJlV3SSympn/DfW
SPUokWbCOeKfBdGFg9lmpzm3oIFZCuXk5U0TDhapxuzIBPUbTr6e/bjZENni/yxW0rUgPuc9OgSt
Fhe1jaeRvqf1jHF52aCDsALqmoiHCoS02Fvjj3hhrk0v8doISghqhV0WUtFujCiwlbG7OPtP/akR
aCSX2Ty78TkS35ECCBgDfyObOTAZbKC3dx7/gufmNw8PSnQb6uv6jlVOlFZyBDFTOainw++522tY
Xv47Q2u9zXCwSBRgoY7YU8n8VhmgDYkeOqGoZffraITO/InwFoG+Lj8UmbmNqOM5Q1bPu9jAbfsX
wuCsuLRQt4JI7jJhi5rZBmD5HBmx/9TWMcfEKOxMO0Hxdz28kzIhwb9NSowdVg249DM6ThnustFb
cV5K2ps9MwmJfycZD5MOVKK9AWCA8jXgDq6d5V05cCFEFqsIK2YrzBPVDYqIZBO9VPbWMhNgKhLS
qdsrjXmTHohn6UIV3iCSz0OIl6xhv3eLZQmqBQAMQYqy8XcSwnNpDLqG5enrMMdsrM5MPrDVS35N
THJwhQ3Qt8UL1YFIVsjhKw5GWqcPBNEIxxbF6F4FQuFwd9nLXmQuPO/JPgKCmVWx4yFF7GM/xviP
nRKMbXU+/ZrVdRGtnWQ7mPT2wg7cFsM9vtkI9/7CFIOxm9yIyRUydDjIj84YD4YcD1KBl6pLRMyd
LufONMyLT0cez1leewcQsISENA/tjUtuRq3Lncyw6joZivt2cgIleiGcK6WNBZnSzDXa6ocluOAm
X8wfKQdYoxwiO+mtYPBqybNxn9E1WzxUBeng7Mh9scttHIb0WMHkNcaGCuFWkySmpMrDDPOfddn/
3QvkgPGMEo+xLBNdB0xtQDcEpN26ag/mbKM79DbapWEQIb0EfOsna93Eu5kS/N4c1zrVyx08Y8hr
35YxrMcWN+rE/evJqj0kjF/oDNwelmRFtQDlcwjYr5YqQ5PF3fcZOSV5Yj/wr7+v5S8WVJVevsf1
bix5iXe3knZ88f380GhHv+N3Cybd2vMVlVB/T7koK9h8npgNBqth0UKB2kWq/Lh3pU9HF3qPqeQy
QY9jFrxAcJZLvh6jAjqN+m1ZHT97kePSBG1aobOmfQuv1/zEmE1eo7VXSoJmHpvcQ8xIBSgLMoUA
noKMzspSqdez2g7zUOlxT9o8ejNUBXbz2P1RI1ll3ckDnObT525BRq6bBHNIANw7AWIhkRwNxODF
O7Was6T5jkeDmbgPGvteRuTmw+zSTmkaxQpF/RUmShpXgDUd+zQjpeEknibuEjCftLa2kAR3eoGl
OULCxdsuejYemruAQJPc0aodaCMX/7NgA0ItOLFKOrY+JiRwXhwcK50IjL7bE2AmwJLuyTaI7NaK
O4OsPjnHJQoMWRbJx6COmyLhC1WbZuSCOdyGmDVMK5jGoLD4TvU4vZkyc4llkEUYhXS3sGF6mEbY
NzVEIRRDjcejEZb3qIInUQbNEYAZR1q6h5z9uttu0DSTTur6+fnqZQdon6Tl3q1s+ePMWYBhNjW8
g59CFFca3RACOD4Gzm76xHL9W1+xNZ2EgruZY++mBUXZvRU3Pw0ms4ala40d7t3YW/BFHRpmzvNN
TpxviWzCwKAMA7NQJgHyLaq7yVokIj2CS+jXdyG5evamqVxSeNZOXn0+Cp+HrLNIgYBkpzCBGoXU
4ZUnOmdweG8mDZZrtMmuc3XIlpv7cEtR4Y1r9stkiX+I3jcmBmnTMr7usgtAn0sbcuFaXpaGZBim
DnvT3x91zvWRSRWCbUmkPesfRBDKomoJPBewvfo7BAUfgBTDsdhlyltzYT84M3oUn69TueHd83Ph
aKGhwn0GOnrnYgTYRxTl3hF4+Cv+AcnFibNbbym7oV7fOqLnJZ+KVLVda2037fOal/Fb/dKHJBJP
/CCYLyUfOF8MhIIcg8JKpMRCQj6qI5zSdnZDdeuF7a8YtzGrb2T2bzKKT7Ptm3jAEILVIQwp40dF
NB/Sw0D7EvRzY7lgUi6x4DsHaF54tNGmb09FguviOq78sqX99AMXb0e+lBDR9k/r4I7kJe7w0CNa
AeosI6ywbIBxJddTM/BoQ+HcDrWdjXUhbhsQo0dKnN6Di60zbEa10baJvAj1pgfEIummUzc3PEIS
zjaXUHmcOIur/yVDKZ3HalNtCphhCCd3t4TGN8aBs46hW5khHoL8WGmUajw0vuzmxjvjeI7XAnuv
dTRCGdlVc86fD3ztmq6K4qRTVe8CRH1tttV1ulJ8/nYVN6lV095mJ31mHSl2sFgopjzEu5aTbQwG
a5ZFG62QDc+HK+P5awiaV7k/FiEa0g6vhXMOCO/bIeBOdBqwMG9FQwKkGkgep07Vc6Pj2JzAeuFK
etC8yz6udeuVohs9Ti0XoxEz5Ccjcarc+H3NaC3E00Ch8F+KHOXwtSRFiYCFeUuO1IGNR7P7LbXc
DU+tpz1vzCa4zzMK+Z5BFJN9kCo9Wun1XR1DqwEKIqbf1yJmJLtvBAnutlP6vuDyswxFTvBusN7N
SBsNOYDeuELr/278Nfz81o4LYam7Cgd2Obnh6JhNZAR1QAzAljwIBVA+1JXnHXq+xSv2tbMYx5Ay
MXR+rUDaHBjBEgmFy+3jxwsMj3r0/iSS1KKq7Hv34LFc4NtT0HYV9Lz/Tf3Hd5Q8EECimB6qp14T
oGVt7W6dytSZ4tohmDkxof2wzvoFNRLN0bBguEMeF7Nv70Jy2qnn11YSjpxyzAtlv6zHSu6edM0r
vt4gA8cZ90GFBbi6wwhbgFdiqFvvvzSV8NVBMaXMkbLfXOQwzrPHAIw7gyNuF/a2MonHEGpZR01+
DV16DxLxkt8zfROCEpZnyGgOEdEEOs79PHzXSwmVsvvZX3avZk+U8W+a/hHM3dX4cyjgPXpgsNTw
V0E8lremF2h1TKcOjEGtz/uu4p/jBFtZzX7byQaWtu4/GIlqzg0G+Mwk7FRd75FOQ3O2B0u7QKtp
xvdFf3eStLxmg3GdR1G3TF0ikxjIVBVWJyPPzB9xTmPjoinD2XVAeXGnil+4KkL9RtlalqK0FHFU
zJ6cDTFPBvv4KSBes4SgUhvKbpgycvYW1M9hV/qRDiDwx3ACU4FHxUxCcnPiq3/xStNOWzXnBOae
gG1YjBZsjelE8hGFnGl+CNqGJ35yNWYc8DzGqIB+ZHwsBIF2NckDYMQMY30R5cEFr5pmT3lefhXh
sTB7V2adFKafW4XWN/QiEqOqqGdI2k3kvczLIJeqyvm4mvvCwooK1sPqf+Xsgf3bPnxhNm8owZqU
RE81Pe1k13FE1p+9qKkbQ75hiCn0ATxCrxTheNFWMzwAGn11+hIey13FvbBqqEKPC5w/mqdxAjeM
uwI2PxHQxeRJWApGYpo0WDN5SshDE9QQMOzTep0p/yGT9rJYrs9piGM5pHvK7kubgWUEOGNOpDWo
DPY8/6cIruzoTF/I1vYyLn5L0OHSeIG60UbQhNf3oBxJk4V1ZqDk2ysHLJDEZgpn96Y4I+vq1NNz
VRO2nZa5gZsdkK7rxR6ZIfKgb9p1mK0ljkDcBlYhbXDKMAu6Xt7720MdO3bgfjTLszy4e7FimqLQ
zNoqRUJ1m8ueANYkVagKouY7QunvA3Ek3xNSCWIm8hLs9IyC/rhSqBIY7F1sh6vJkt1HRRPuMeFd
yT4zLLN38d/uA/QEBlBdty4iDOCVdMpbcbznnKI7TFx9rxqbpCRwtcbIYpNSHFRnk5L74uVYJ6Ye
5WkGPkCtSG8meP9fHDb2WnmC+3GUBOoeeiIwzwyBytxzAG51S4zlQH1N4lAqNAXamjwbQxzuMeqK
WBwb8zVJlXFm3BthmcPwEiYG3MCXGL1Y62AtzkqXkLtpeeHrS6WAZjfQ3YoJtPjDOBFK5hiFWyna
0oC6jbJO+DSJpy51BkQ4TAzNmnkMnOG5nwQS/cMkDRfEmUxomBoDmXpoMv186sgtURf2IGUxzuMu
39lcPwmYufIl61d+YMINGa0icODXCu2AhmEQFmAqBgjbnKwapeeJrTY/SDDBrqQ3Ih83Doh/WHTr
hMpy7AF/M5iA/1FLVOBCZuC0jYgr1EUqDgAA8eDiYp7Ir15zryWlBzN1g07l82PXJcXN3OPjuGTr
JU+M+e/ZdGh0KfPXXfWtkpkRZUIwTspuLJaEr4dRqrvpQEqXe4I1PKZtZ8UZ0ko2hNiOuJSb79F0
Ag8qSuY5OhBNR0HxKl8LWszJj5PBjO+grLnJvFW2IWAv8u0+VEscT+sKEDNG6pfsBXDCp03lI7JY
4JzAJEDsrGBddOtS+6A01NxlAsInxJHRRaQWfGoCWm7wxmPnJ2pl1ljcQ6DJXItulMxXqLEP82yh
3Dku6f4jMNA5dJMiLLkzPQgXsRtpI2bhMYGJ6kiPTCeWn1mHMw/iZiJRuilEtiYTEvHoti7NEQSn
FH8hW+g88N0mR4e0qklVzc0vcDx7r9ucr57QEBX6aIjCD1F9EJFOmIqbX3NN3hfJn7v8DvMoaRAK
0C3MBxyJ0cP6arPuQAwXzumVPy2/YU4W1t5c8COYS6fEKfeDeDqWAyDisyOemFN5EpfJH3dRS8oz
/aOMTOZ6qlziOySpCy4OT5x5HVRqkT7MqGhyjCxMZsaXeN+Jj/QOc44FpLLRXsWx8sPYEwWHazGT
MSygPFxbJvTev3ESAGEmPIIXfFgtf7gPtPm39qTGs8BpYf58Yxzuvz0krO1g2INqNGE98aoA9UOE
+meacJH3RSgyvl8YrXDIDI5qnPHhSfDd3/x1J1vOYwi4HM17cx2MuLdJMndSZWWcWKtyD10wVmVz
5EtiBkCyoOWD5/DZVbmZHD8M1J/AtlFkaxS8qk/ctHBgXg49OAwRdfW8Lpb1620XjMVDVyugqe3w
r1lR2gyY7dAQuWxwBnNOhA/LlNRMscQzPu9KUaQanjdiu3eX/HfhbJwdTPc7OeHx8Ag9SlDqIsYq
6JH0WnQ9MxUzRXXRvocG1xvU2eih9LIuDFZ/Ef+7glUvkQSwKvZJ9mmlalmkyINtr73c3YRD/YzT
JleFIpy4ClNC8k101Gs5DpfFp6WsTnMzzWADvK93jwHyIUxmOg+lWz13v8jngngxj1MIEIV1REh8
ePl943Wyf+E90c9Rma2Xv6FTC9MFCvd4rRV6YBJ6MSSba+s9gqZAkAR2aTsUJ9Wg4ceGTMmbnLhP
TBUVoMmt3scYNNa9XTvDufyV+CPvRGWlQFAO77sZ7JtHVsN6/tYsq9o/c2EDe7V4Y4Ue05TvBnlr
PrHZDpFlrs/C2+3kgizfsimTj3Qb9NV+/R9llWxFOE6NfvCafI+hoe+A0XvDvy+ZuS79VAFnkRq8
N7FmHE1cTQBwTVZN1MfFmyIThWHu8dn5w7nApVO5GYDmPm+URo/CsDw0K6uv4FT0qzUpO7gHeqyP
N5l80eFLCCnQlXeT+gqQobofvUpwNxmPOu6t6IRrt+GEeQ5ij7r8bHOppxoY9Vyhl91QzrUn6PIK
6GWYDV2RoTBfV3DmZyGXG/6/KjQhMezLNoZWjNBX+oj1tU+RoCnobTvxFdqmTlUIVr4JZdtnB+Sz
SlqZe0qCJbInmzGjbtsLxfrnoT5jMJ8+mGDzZkCXqjxACbX5D5lmFe3FhAHdUSYFL8CoMIu97E2W
Xs4G4zME46ZYFHh+GOM8Sngh7TyEwn4I0vC3jYYY2WObe+kc/6l5KwQQ/y48ysSJ75/3pCApzux+
d1dmo4HONj8ZpmqtWphow192wUeF3SPWeGUyoLFpSSKqQ81TYyr1vw81se0RamlMTMQesTH2uKvR
3fmtTGBZjsVR/dOBC2FdYeQikEF9NYV9LLRO7V+o2LyL1pPbAnXL3qOQ0Obn/qes6SUu6uOCLe2A
4HNFE7OmEXAVTIaOE5ljdq340Ug2CxPe4rrefUmen8m1oIm1rm7fyIFlLGeaLUBUwDDoXegV43M0
wUBx/WWsSra6fxavCca4IzR7h060Im61WHKTQwUF6gzdgKi2HL9KdzSuzrMR/k+puVi7IqXNIqOm
8otn/TIYOkmMamVMAd8MwSQmkRZk92MPZcPX+36x6nBAME6VDAWsD6SYRwoMD62H9tt8xJSuO7X5
iitPC6Zfj0cJF5xPp0hgT3ErHiRrEv6i6h2uiBbVXLkmvT1aRFM+9DgfM7mWo9BHNxSeyy03EGGz
E/9oxiUyVt8Xlk2HRdhx/x+FbbHPZ2chBVGAvidJhV3U8if7ubLnUpzlNVanG5ufG18bk0FKn5+C
mDvrzxCFSJps5CznCUKc2REO8zbbYYplEZW1MP4gx2IYGLraOkFba3CdGcl6GzmWjKMhO4OaQclv
QoJDjTF40NeRaoNRASor0S7lWSeioXOj+sASGvo4KubV469yvPNHLY11HNpdWnq3rFGvYBetsd8w
MTlw7ESgMVD9gbn/X1XOVRCXIbKX7C4AYxw7GhWDwR+CwhPjDdPZ0IeVTxmkosWJQHYI6ukyK5y2
27TuGmnlvCQZeGxyqlbPxEL2Yao3YKcULubk8ySCsHgapBmKPcEu6juOxUL0IVuWCkhXHLl7l9Y4
DYbYwtC53dquJtUYuo4IBbn3nKQdzhVRiXj+OXZECIO/p/+1RXUp2h+0MkA/GXNr6aye8ra/kAvb
q4+nUiQzC1Qxme0mofXcAhQNalXYdM60RlNuCJNFbiPHwbPGj4wYtp/nvw5oblIpxbFwzimeFkiZ
Xqcv/KVB4e0by3EBwwKiy2zDEWlv/JODKRjseB944DUz0mnydKt0Ob0e0KfGndgFoEZdTAwr8GvC
XEm3VBZFZ4UufA9edQ3m2af3cqZonFiiEjFdq+L6Cdz6cUXE8RR+cDg/0zDMpOCMgC2PmuGjU+1z
bI2gkT0BD1LxyoDRlijntUsckkPQ+WtvmgJWRpTw0lclHs7QYNcZxfhqyDhGDDODYaqLgrljAY8i
ZQFwgE24pxMMb5+8VjJBrp1K6Wh3cTEQiIFz61ga3yo9fRRVeHVXIeqk/xCaNGgKT29cRQjmMH+p
Halr9+lxOWdVdHT2LBJ5FPaRjqyP9Gm5LpSShN4HORUWR4ZQNtFh0ILvEVukK3hp3m4XXOlNHZw7
TWc+SjhqFxnn+6jZqnghg8ZE9euWVDFfPdTrMiFhft+bjOa7MoreXTH9yCWMZhfnR3IbcXIdE8Z9
sGM76kPc9ZO1GPYmZ0fG/key3PMElFWu16G7LcdlEw9YNl8O0CPjoF9RUkoDQkKhMAuzXMiTKUT0
IziebH/66vDSipiLN9pUqlfGNZP9YULuJIXQcFI+phPnn9iCwJnVdZ/5Um5PwoxmkxGGtaxImjxc
5XtOwVp3EjPSd5LaLLxJb5e4NJrVcbOu7KK1W22j79gyd0oRskc3A+OLm1hM8HTAE+wo1nwF5pNu
PIqjWLa5vMddU0Cu0Rp8JOtt7y3o2QdBjOTkOUKqvxgJQx4xUN3uCRq6B1LMIl8wBW1y+vkb8WiG
4FDbmjWZvC2/lIwklcBZb1Z8Mio7XvIywoQSnYvgsaypHRIYY2V8m0Bsddi5/pMziChdNnLHPpcP
Y1E9+28GtJIK8sJ8Ke1byccU3rLPBfHv45Yi2Obgw8S5a9eabznJ9cvbYN3UO+8goszgtH9TEMev
9altaOqXQttF+qJBpyTRWVlG3e+kL3psUyig5FYzHCtlcIiAGiVG27WOa5zavopzvbLYqIifXIjA
HbUS9/LAw3xxMDU9z/JNAl20IQ7jL2zsbf8WM5f4Vxj3h6lmNyrjOG3yve0FLyemA2rUaxoqRAzR
c1Ihw+T3mjhyy+lwNmWPWeU2afVVUfGU140CKXujUpPZ7xEO5vV3eKYb0z9pMWt1o+2UJDNMWaZ/
r+fbGzzq8X1GeqJE3F/ZjZEMA87QKOpqXgT79OtE0+H5cdc4MHjsrA++qHoQg29mRBzySx1eSDjB
gcskwYFMzzfsE9PrOdTfftzqm5TnsGTBiqP241E2L8kbr7cORhFHVSJmcbyH+dAS88wKNUTd72OU
BrxKeaUdFHHXu+R+J4qpX+Ypmaob2XcgmnYIL/NVPWQEEPPwTG0gGC4sYYsuJpPrDe/cEoA5PUWm
b4WYHSpdVlcC+Cf/n3B5BvMqKnuo4IIb1gbLYlHMQzHpMJ73EBeTlIunyRIbv4U/W5a9PUMcbUX4
nEcSkHaQYOETX2M/gSGayrCjsEOy8A6Btfjvxpdhu90DXoAMkCXTzt/iXTf78sBFR8ImcWEPX38U
3nlSCPTqiJJF1cGPJnICRNFn8gtgP04KBXeGRqGsOB6xL4LbzbRB4bvi56bLkXvHHKrDoKYXY11J
7Lr7C2DsKSwLJER046JKt27frJM9ic/1WdfOEzrnXaVCfFu0/NRjB4cVeO9axabXZnLMu7/dTPGL
w1oNR0ji0cTsvgqF1SQMraxYwlAf2H/pPsPCT4cQ6c8N0/YzdOJctxx0AOasxuuPmy440ifiaoeJ
7evGXa0Q17VeEasrZkrYku22ouCHzMQ3ffpf5ybDZm/+MTweOzPVUelktoPlP35f6Onfj59aX6ar
3fq1liBK13OGnM/cI4uWSdPq/s2wX63TE8FvZlyrikMLd5Bqy3Cer9WoXqHC4icjryNa5U6IEVMD
YYxwJwc6bNLOLX7MiVhtbQOike+HXW4uSRpbv22ovov8cw62mlsz77KywsN6CpQ/k1h4i7aK/IzW
bQbWe5+YkiwK14/Cg5Zxx06k0EKaW9CcPiLu9XqTHC2e+VLD/kQ5Wf9PJN3otNMR6li2KMZg9mT3
YZkBnNFulaMt7X0NTQNja37kG7+Tjyh+mDvye5k3vkCm9OvOPtexm9favcWa03bsXH/+kJW06eJ9
eeTlaTzWphiRaOi1yvDpqYeArKfiwh8zsuv/VB/RdBRIy/MkUemg1diN820U6AxzSPVI3WvS/Pkv
P2U4ggjKgzTB/ETnARnXxk95AeSNjUsoI1yJy4c3fecVKfWP3NcxqRKNuaZnoz7vjj5roCsuQk9p
QWbb9d1El+CQ1Q/fQfx6FtFtKU/xsNBgxCDJyY80zfthq8fdce7+qeRndpLzmk+vO1oQLSbML9Tj
UVdJPqv+mMq+EPxoTQHlpi2yVgVxu4+X8BhOelq2eukqt98fbb/2ABT+a3dOD1VBoJdYgseKAvPU
7vqXtL0UNtJcIZMcL66PfSG5FQt2pHF9n35zwuiIaAmHkGn8hOBNctYpHBQBDIekqkR1mTmdMJjc
isFP3wfYSOdFUM+r4Lzqk3btZrGZVeqATJexPLwT1tuC64wtxeFopvUyGETKNraRVofD5yf9jpAU
wJxjWSoLOCwom3GxqBz6xXX4HoRuIe3leT+hoagxpoi0ZHieX67Z/zXaj73IyEaRxAQ98GN6aTex
M09fhCMSfpeQ+3b7/PXqSgX0SA2siebHsNYNpokJ8rsHUNdVkoiP7JGwfQBTiD8J4cjgyXtw/CwM
S4Gh13oiKTNqO8cSxb+5OuR9oiZdL0ZjguYr9m8I6j9rSVhmdB23kWnu46OV8A0GxiBVf24lGJZN
RMNNNHtsGUMS4i3kFSCp8Q6UCBLn/qQqJKlvXqjdUXZWyYC4gN6LXpd5Cq8Y6YqRrCWKzNfFv7VJ
P2zX5t/MSXe9VOR3GoOVBdfAQdMBuZW6ObHOaGdGrdwdg3rauj4cgYEmkJk8w2CfxAQnmuJN2x4Q
BL8pRQhDqtUKDbREuAbtvVhubOXbZcGqVeaD3wvr8EgSN7b/AG3r/aNYMNbZKsLY0LWMEdMJt599
FfeLQUYBFl0DPH7rbYbsiAqahNDOIiHpiZo4a+P9p9FsLKP7/hEOEG5RkoUqTVV2rIjSY0UwNgg4
qkpGTToRJTPqD/hsPBRcn/cidhyVjc/za7cH9BtCq7Wmp+JNqfsKd7ZNp20jVzFJPOizpE68FFf8
O2aRcmGa7XhekbZ/P5KLywG39WQR5wWVBx/RPx7jPPSztpcoB7XG+Sy5QegbKGG5LgMJB0NG5EyH
+rRwpHhDaB4QjJJTywU1nBc+A6T7w11rQWGbIHPXmMRdL/JUYvO/HcGiNa7klcRXr4SEQdvwmrLk
qArTq8yl6gV5crEjbQvB1xB/J6nYZ2ilG3n4t6Sd3l5F0B0aKrPYaLb15kT3QIXefwIxaMkykU3k
CgT3XZYCn1qVouYFjrNmCcfjrHdTlTb7X/QCpGF3S96tzHLFHQZhOzVnM/qSYAWAcKq9pOIy44aC
9VOb6ECk9T934p6cNRdrYvNPieQ02y2N14DoPlv7LDtOeycUrdykmw7aNoLpGR9pQcEl2LCThu8U
Zlsx73tiP3PodaZ3WWPCFLF3zwdu4Be2bjmh/S8PaHyBLXBIe2FLFsqGrDyunODVpFcBkgppIjcy
BmxyoeRgJzSOjgm5ogNvXCrsmsavNMu/YKKv+qgmPY1cV4OW9WIlZNHzKnHvbYXaUeqtDzpQeNhG
5lPTOepuO5LuNVWTG37et/R1O27f+RCTrLwfEbQHV1oj5rLG2WZRYgTZpJLjduqBgRiviS3kBvRl
cLHsu+6QahxERuk5FjjhC2aFRcZupBVPEvUtweAm4gzTLH6kosKfwad4CRo5s2I0pw0ERk3Z0+kX
E2MX7KYwyMWl/3rA0kZOjn1b42nuRkTTb5TlQGNhVARnNJ9YnpfERGgzYasvutifn3RnhjUBqdBS
5lT6tFML5+cIjVFvVLqEWxk2XpA46sUmMf0bvIUvrSw01qEDpSbJny7p97hJ0vtrIuzq0EB/KPpa
oyHU11nLN+lpTCHw2DoeC/GYVZlSJm4E4vJ46vmxVjGT7BScOV9dVFQ08miVP4JvHaigB3asULj6
HG5CEACKNHuzrg+MCWZwHGPftfQ9JK4CQTlgA9riiXYcGr8HdEz2L3oodHfbjsJBgw7yJQ8R7Ouu
Rj7CnW6i75XeB3KVkiroPuywq7qUFUJG8uYlJwE3QuiuJ+5f/rhbr88ftU4bM1Wuxsdl1HuZ+dbU
2VWJ6v8yCdNXyOSuC/I5r51tf6Q8zxBUaDf3n4upEHuLTZjWCqgXZk69HOlAXkqG3MxqoVR9OEp0
mIQVsTDxTlKgHW+iPzsRNS/9wUmz+OdCdBwguy+PTYvoo92kTh6GmKRopbOQhw9spAkpZxwoN390
uCsN7C5uUv2FtteU4l8ltmIj4nAel7pBUfEvGcrmXQrspQIp+PIi0h7jNnfBKlvB1inWNEuqMQL5
X6MYBH9QedUymFtTutsRdL+rnrp5HjKHCcOAosgbbHI2Z0vr+UzKtVNbln5G+AXu9CYWZFfOE0xM
96fjaP1SLzWrTgX3MW/neP5fBui5yE8NRh9dHyZJvmIVTUWEGFg3FPIYalfyJvx6ThE8EUtXlPCK
ffxjjvOO0LEvSIBXqV0JTj0+h9OsPASX60PqAI3Pd/WpRVLSsOtPOooDNxF2Bh2wH1pEIQMhMhyG
RNqmWRG2M+v5q1tLgQnlij5UlT6kVtSAvkN9aLznPNnGlRCWNjMFXQOKkzJD+G2u13n3kH0HHNXZ
pcq4t7to+zUdUK/DWAMHgxu+thJQIAkaY/nsJNnOAifPQ4f59ExLpugHf+Ahoybm8mNSe9jn1eMN
zk4fO8owwG6imm44q0aQd3CTAxtDIdMtF9UmGdZkjKu+GhV1o99Op0xdPBeTUSNKaD7IYQCLUmk9
F1PN0e3c7dVf16xTj8qyNoJ+0uyuPvG1FQWoLaL5zPDa07emyxVCDA+UNpWvWgGcKCJZ4N643//U
3a7y0/BbEhvAc4ZFAkpHcKOReKjWCFARvoxHV37rkKd+80V8f89HvYBMHHhezjLuq1Vng7Y/n1PL
y+n8Rup+jwew0JnD7pM6X3f09/Aduo7unbmKMzLNEZaHsMCoEQtuh8DhpeUGbXnkS7Vku9I8+T5n
FqpB562jJBJLyCP+g5qDgyeWOfHiQmyXLlUKYO4BK4lFegZeAcsoz4c99gzwRfCVMzgKq2t4rrqZ
wyHLFayTINQ9pQMzrgp/PB9W1c4lmfyyDU5u1JvYYg7WJMJTvmF8FRQ2tocw+URjZWQPqxOyUCGb
PyTWaG/v8gRNF/FnBnG5145qMityOb06O8/Sio/wmRFBNsGlxG9HiURkOuZ79H229CxD5esEZzVd
QCdca9FwbWQe6Qh4Yf3rO5nXKF6T++HwXaET2HDv1mCGCfwx01QZw+FR4nsjCQAoANUeF2Zdcu8b
etck0w4UK1ZvFxCuKrVtczFsEUDtDy2vgeSKa/rEAUvwc2MDKq6dwkOvuLUC7HcbkNBA04/qbHbW
DjVoQrgPo8H1IwaznlCQsXA1COFSIwfAsnHwmNYZ57Xf8hmf51YAM9+qBo0KhxuOrgwt3PXlYMKy
l+F0Wkp+VhsVK3qhRknwbY5NTQ40F55ZRbnKLIFtOJW42+Q+je9pUL2RZ/yFCR2fbw/uqTAmoRIc
7hGeWSu40QBM3WRTTFbieKVQ7Z1xWT5h588Tv0gZQLwrIwjO6GWOXIyPLlVcpjFaQuYYkbiaSgZA
3cWBu0irlWZdXArq0joCEHlhoUI4768z+cryOkrCQLDOzJwfc0+3oynVhc9yvd7Y6XtfTXISZKMj
YCt9pCx3g9KP3n8AOc+/YUMQbcWluXrbwdYhUUCD7dA5q3zC5VmGjDUy/dPJjeplbN6ydMYWKRAh
YAEZKjTdLl2X5IRkz/ZVwSqjRRBZU+Bxoi4Wb83Xc5fB/3ANTWhQGkvExXOL/qZor0bqnSG/TBru
l3nGdRW4Umsl2XIb5PLhOpbfDfxsgK76ATFB3MzabRPOmmfHNoM4AtOLQx7dXmyIyzKvUVEmz/Xr
gJXSPYdRIPDUwurDYkCoCpvjSdK9ynbMiJ5udPXcBqUpPvptszfzXMC1y+MelYo+ktyQQhuMQtcd
Rrjzy2rc08lCoo2Tk6+JFMIv7SBSm24ezryuRCU5sAvZIvGQXnfQEU/1ydJqlL5BhWRGDIdEkdlZ
iwSM9dmKRFMoR1tu3iowjE1YHgo8OA/AeXfRiD4wVFd4QvJGZrpHucFhYt7s36MT6qg8kykvFHIB
O4EbFBBlxU/u2ZON/8KvmnvaSpENZWO5a6VUtRyRuOn+SrC+0DErIJ+C0KDsKTHnxQlJd5jcT/Kp
NtgZhrfzK1OQlQxSrcWjz8bbiecjAJb6ru+D4+OohfCbGbTuwoR9jlqsYuu+m/LpxNlaPZ3N1239
MTnU5lZC2vtX/NbxnEeFG9xYat67s6QVzVv2NxXsUsmB5utZXzL4a7vQiWaisQABfeTpMc/ziPso
6zJXqqt53vzQHK4hvh+jwSWIrZeKUcxC246hxFNRpbteZokap1zkZYk4j1gmDiL8EWUQvL2avz5Z
rtxwpJLpSzm+X5Ii4KsFIrhAPS4bVQWxRkGCB9HVBnE9TR9wXtnfDWSDq2XGyvxXi64XUH4db5Jo
NR0vKemMOvN2g3qO5NyVesRhcMHwrnHPFw3GbZo29ocIZBe7xgS5kQlXXqyeXSJOSQ0NS4gT8xaT
WncRU0T6YwU27PuuQ+A97k0zYdSOfXbzrWlr9JxY6wv4VAY0oRvyR0Vbq68QY8hrpNawLsrbj0Xo
NODLpBssBzKzkSIMoeF7z7QhD40Dlqk87ch0X04Ta85gz0vnpYAcVCYYJgz96uvJ+xa5/248CvJU
zkzh11FcNuJzo4WK8yuXjdWx0/PV7cBdouWjWHPRFoFUT0EfWGdXM+zyrSZsVpO8pANHXlw+Mptv
KVJY6pDoqtm6glvcV5fe/yvFHkGK3KAtMKqTjB5ZQueNJgng6uffvjMU+Y9+OqjnCu+u1hJL8r0E
1Vh7uh2owIVCHNLxfgigyfzixq3gKK4anaGsZ/8NTQAl3+9o9NHvQOz2fbX7dSNJbcTGz76gulyg
Iagdm1RUqOhs713lRH7EbiKuQbM7IJO6r5Au5zDXl8y91TdKIRHu8h8NG1CtmNx35yXScyD9DdOq
N9/T1bBS9nEFV+YX9qLVihWG8MF7Trpv/WRjF2eUSMyixFeIE3f9i+H6O8W5sottim5VHLoDSnDF
27KuzDQluXgdLD6LOmpDGXBB+ji+cjV62aPXHZHQ7gqVend2wc3AjYRoxIu6QX5cgT5J7IGDKFT7
t252jMk1IUCWmJHFJKkpWEceGePnXiS4qXhNExJvsCOLeF5tU5m7xYOZmoGcLk66aZNryyUXofLR
9iI7f525IlPSOSg2phts0EgJ/qm1XfQ+TDVzeFfZYDUqCRUwnsZp2DjUXRjs4HXT9WfNHCTiktNj
9HugOnh9kOySkcm11r5a77JC4XriCliPCjpkUCUJWbRQBUGqjG57g2vI5o2CwhuhohaF2yysW5xm
6ePXOixs0PEX0pe0xwyN0WHd094SpZXlTqfjIdKp/fNRA4A8KtQBVBm/RuDmJUFAcexzzlb4iMB7
g3iBinKH9x/QRCo7C9IpsMhNDrDwF2ZMbDpH9Bg4Eas3qy9FKpj+EK6qAW2maJC7kKF39pcYaaY/
jBl2EYYwkGyg4WX6wYgi7vpDo3wgQ3i9yqCjG8RDBlyZmXFJGqETzBGjK9q8/XqLwb67Bk7PTNns
WskPAtJxlE9ZWmSajDF3JVk7f5jxUtuBHHz9cW8meMIO50npaSHRgS0Hnl+ii+kI7KRirhJcb8qD
kbAC2DIqrl8GPrbrGZ6PviIxd4/lmKQPBq6qc+DWe9FRVot1CsfYc60ukwZ/XGEYVB2a28o/Im83
hQ93Oei3FUkiz2a/IHe7gzrgTvJnPPQZ8Cym5YhrFJ5u/jOQD4z/xRWERTEw8x98IdD/a+uSb5Lb
OFmX8gGZpcs/JADF65rG+4R/aCJEjyrhVrX7koC58cMWgzWhqbAp8UrfjCU9N/Ifd9SHUBUXs4y0
ly4ddmQomZ1hkbT7Rk0Z/IGR2NpN7sWMoH8dSv1/g2bNIP+D2n7wj13iW17sIGayymhRUtXgjn4I
TOYZF0QIu0588n1PDK0SdYG2M4eqZgDRmwa2I3U1mpVmerFPPSPKfHVYA7KWIOkTE0DW+GNI9/W3
SL/6kYS0uESo8ZWmJw4VAVHCirkvicT2m0WQFLm3v4hCo3a7QQXT+VCr0HCaT/5mwMyLS3RbXQPT
9OL7pHgxR9v8KSPcrB8vCzfrb/XMdAdB4G0IyyBHpmv8tS/0jX5Z58TaztHvR3Vk4pns9ZZ1Cax4
i09QkYajEq8fLKq3nyoZwz+zta8Qg5yasJWaqMu8p/VsA4ecgwX8r9fyH0FmLWgImzChxT2vDT80
nAY2e1v0bd7xe4KBqwaGcaYt1y60tudXBrvhR8XX4tHpREWVRTEykarnCv/6VmXWFYvlmX5b0heg
r1K+ieITB0eCAbHlXGWOQXMC61pv6ZRHZDj/JAs4J0X+sCUqSi+oFbw5GWgA2RsBAaSvV1vHy8Tn
wjUNOtA1uZlEhuX3EUPeSLLZ7nSV4o3rsyih/M8qAdicfO4Ss7SUPuKbzCg9TS9WeHx5ZAPkuQV1
fiSBQ+QqylC8vkCq8D7DQ/QmgEwRELV8FqQC5lJTwNCI+NDCWUBdcD7rkhSVTuiLCoWTfPAApoHe
JAJah0LYRc4Zo9mknhpXvjDrfxpUj7J3JrL1sX9paBu3bM19TOgnpq9l1/5wzdcTN+5CuP6Z44CV
qalZAWsN/OiHQjwCjpQdKJPRi06cMK3RoarKqoTRcJMA4v1Yz1gtRDTJYFwjJ4wYB4sMxtTek5DV
f57x1CyaswBL/vZKAO+U0PNBWDmUzRMCdKg3bwjP+3O4ALm/XyyIv4rRbej5aZLzwBV0dafA9+Ly
cNxS+b/ymJ3hrX21wd4u1cX4M2kw1UJmPOmvsOmyTWKb34SuOBtNye2ofCU6xOwnku2kwODoqTWz
indDbXAwQ8h39F+yulIp9vv07mwHgkHs2OoCS9JpJY+yup8IWc2qejxj0agh4y6BHaIIX4SE0hmG
uIcJ11wuGaUXqp4rOlGqZdHJSK3M9P64Tx3HRwUj7YBi6l7MRM8CSbRZTW20FcI6ugtYH7hAFNyg
4Ru4SXV8EZKnnp3ZauJHinmmogBKkLVMUAaC8lfaq3nDDFyqvlhPrZEQsZmkaBYJcOBILx83/nFa
JlqyO7jn5nmxoeMnY0OmZsp+t7BsBzeMTLOfGKsdm+OghDHq6bhgoI4FaZWyMendsSkP2JNfvsPG
J70/v/U4FE9MTjR+btW06EU7ugeD+/SNH42HkYRE7BWpMO9nFeYW5or67aXyUiXbWOKb6hhWm5pZ
BZ5gUB8RLmUVUZdtG23ZUwoddSTMvWdinNXXyFDaDjmIX5fhu42yAfCLIwxlpxyBzg8K3cVs28Rx
9iLsE4W1308i6chdYZCjzqbYdJlqc/PQ1za6uUhDoz3k1BCRmKZQlYLdQCS5/WWQFJT/ioEZ8Y3L
vlMNfDNtGuL/Fevt/EpUbobft604cRLZ1YT3N2pyezfq1GyCFW/RmLokaVhhy/MSccmXmNyXs7E5
WfEVV5yWs528GEfLxiEBW9GgTs2Sx1byZjkAdOhPMW0kycg8gPOyKQdrtsx8EyLVjZRw7mPxjNOz
JnI0/RW2i0scEtEAizM68Zn5z1mN0WhyxUAa3IZXpez+bt1gYULXrc22icpGz/enUbRYS+bDuiku
oHP9LLPcBcs9hLEF9h9Im3mkW3A5gP789Aw+cGUHHcqlEFw2xcCjk3mPcl3B100oxmlme056NPlM
mXEk3CZb23y7pC454AdQ9pxPJIG1DYlyNMrz/Dl10owWd6j9yh3JWQrkREVi4/mblLND3BU18kFd
430IpSrkzfEIZXqW5hdtzt6P8nntgqz2zjXfD4thcq2nFe8qY2kmYv+pG1MENSiLfSGaOzm3IWMT
an0SLB/ll8hFejFda8tGrKwvgG9wWwgLOsq4fyks6pY7mVdqoDGDbeNB6vPd+a2h9O0lVPc7kwt1
VwTjk8PixxpOlBRH8H2dEoHMhmk520SrDsTRScHHf62SCdbXv6XL3C/MzI9SbaSMdmiPQzlBn7XM
KwDABaMejdMB/Aflihr/pYLwcIimzTI1BqfnwD69rkXac1z5yQirn3gCI6WZg0v7Og3TeqFoROZV
Zyf+9xGe7NQkL79WJ0sWXOVR54mO5UwUa8rauQubwyenKipMSKDM2+MbCuLWTai6nVR1VSGNn9Ni
uK1ZjKej5yV0AeukVwwcr0GczEf+iLB0mXitpd+Ii6+jKW9a8kM/r6EI5eXM3QFS6iqai1/VDjXZ
bVF/ZsaZoq943obN61MYcQt3c+jdC8uBCOk7GFhD4g8L9YmnMQ+Us7obt1P4y6D9IQlxhx1ZVxbC
xN1jnMgKKECrGT+K3w7YZ6/NDKeoQJOEfOHXGV3t44JHK0pnN66yB+eWvpfwP0++mxIwDI8zt6k/
19qj8uNcxJid1NulVwO43wrvRqJeSZhHQx7xPTQ2EuvH2b0WlXX82sl70l2g6d57XMLpaDMuMRDy
+/UzcEFFLWWwfAdC4HdOUG2iw6qWy6RFOZJFW1nLkbIBPPbCb0LBfq7ANN129dWWq72/MFtNqiDa
EUWyjNKkWISyu4lohCgnzQHjx4zYLvmuwMGUGuEthPWmcXOj0ulpHxRDgnALTSpH9vYTbqye6Wtq
veY064wxQnY2kB3vaHXsiIpkzTOLNJCaFe6VHvJC5GEWE44uwYJc1P81vFwEQqNRqxopE8FdZQIB
LhcN7NkgqRfmrar3Q3OXVcx+Gni2JBceJlWlPA6XPNtKIzhhbx6IpEle+GPKoRZzvkPNU6/Rce4u
mjb0EJlwPytFuC0FZ+bUGJaibRqWLYm2VVtXGF+7VJrgogqPfyOswKMMPy03cbl3RZRc2zyvi267
pqQx+luXTtJF00wRXcQjenXyjO1zlBTwJxa+KAdH5tyrWY8amWE78J692vwvgWq6b71zckrUdV7u
n+Q4a5vlVxj+I9v0rA+PQpC43w1hIlDu0z0oacIl0bA09PZVGJn0r+9EsHBoFdbS5+BwarrLDI8w
KQqossHvI+3uyItzATjGaCMvIAdQNvZqk8cQlCuB69HKRkM+pfpSRhwNhAAWpqPzXn2Z7CpguBlQ
PDo8U2HVyYzU/RUb0fVt5eg7//4iAkFzAamJdeoTmOPHEp2lRhSD2CAtAs1PL0lKihfncqII/5hx
PLPeCVQwg8CTeZf4OV1MlPsTJE/CXFwRoI8lk97mvsXRLkWoklW50F2i25p8sZ3KI8QEwxAFVFM5
0vmVk1pp394deAFRE8R7+7UOqMWoGF4hI8uHH89aXOZ8AH4vXgPCbeyriNxl1zxkjYlEsrxKeysn
31ayhf+oWMRggrECdZESB3UYNWl24/83A1Pxs983uEpZNlOUvICThKUlug5glue0tsah13DDVVZ9
yfOVC573eMfvT/l8C1YgiD9iYGgljZRcNt24R+ff57n42hZpqLyfIgNS0F+N/p9LV8hA3H43Lk3z
0Hfe3OG1MMG+O2vX7L1xeD677gUiXoKn+hSc5642ARkxNBP5EvZJTU0iHBtTt4DYjOwae9YVOKGf
Lued9QG6xTroKkiDyLvGaBgUj4kdtnjyXnSGL7KPf6GtFoAeb2edQdy4HMYBly/WDhD3d4szbf0F
i2cuAClJPdS06Gc62hVK/d73yQqUE+knOhGTHhPGZJ8w4jU4EkLpyWGjNEvfyvnG2O1bcept5GO+
bJ6fyb3j3obT02KXqt/7OUffqx/7V3Ba9tvVguNvBb3F3j8gZTJGjHMYkUO2Adwx3Ha68mDT3hyJ
07f2qGWIwSQ66ntkoZFuHnK7FEqVxih8iTOYNBWMHVsRdXBNOYQp1IKUZRMPHIz9Z9dZNQvL/2EK
HneOajFwi2atSxOv3ZFqxiMI30SeQ2YqWCHqw6JVhdblvKMm8XXrJjSYV6w6ydKPCrODtfKPGnE4
x0cUOGqjgbvqWW6ZH1aw84OCNo2dOh02aSDLkP06vNJBBb8v3iFMi7CPgDBGz9neETVRwNmCXhP+
zXxfywk+GOgo1uyoBRNSl+K+JeYKrZm4fjDOkwYPEnE1ktCZEhgDkhDgTLmEIlACdqKYlssn4PYM
V5grHlk0mmgbsydIsAk7j6FE0wgId+PbLgm4c733AW/aoz2gIBuOOwChi/nw5Lw131LzSztKnEMs
tw8e7C/BodeXYrBZIFsSfZ28gcpOjlC26xAMQgafR3gFYEsUYKs6DofmK8fJk/YQhkosCILbtNow
sGLUKeffIvRVUMVl7enl4ieETg04LcUsczJ5B89+4WKt2iKIqKfeHf4yepEAZHVNTmVMS6+Ca+Ny
e048mjABl+tdL/syVuZGh19TeSLItONfvrfG5rKq/zLj5LoCGq/a9/ltlk0jaW5eJRWLDfw16eO+
obtUC4awxYNRegHJXMvPaBpjM7qFMzx69OTufL8AuiJVvXAqWL2f2mHF8D1ayf6d8OKjdjz05p05
3i7v3ibaNnxRt7cZ4LR2BMnKoDoC9I2BTYA90dnHe+JGMl1/EXLqOgTBsLb+qY3g4adt+21Dc0NJ
xUTWvziggKORvVEDxrS71u+RDaFE4Z0BUzsLT9yR7LlWzot9Tk6UKOf4zFye1QnO0dtuy6KMklfj
LTpVGy2GlcqGfmaxLYZ4a8d9qgRrK5wzmsZyS1+8JMibd5zZDKqJEAlqOG8pOOsBhn5IFxAC7cLx
zkyuCq9l02p+EX2ebEpFi1cRP9zUf6tBlEAXXyZAHW+rfqLxhMF6pGZsFwEfHRvhLB8GxehEtvB/
Uy+CLwNw3D6XqXQczY+q4vgOuYm8zJ+4HD+OJEscnkkZ5GuqMx566i8T38XYOK5IfJCEAaTmA5ax
dPhgrJ22jTXsKFwWDhtk+jE+TEhGT/jC8670MCoYpEMXo4BORFOyR0E3p5GtPifrrgTSoQEvza7C
bZ5DIERefrZkNvXlJE1TmQFWanuJgiS5V3sSylcbHgq8haTVqCxaLcLoYcvX6pNhDv8YSWaXqtKD
92cslzfRzhiSu5Smhbjh4/ZiFw+gLvU1UpwhpbGj9WZpB5tblyk27wDCmYgzWjbKzQTc5nT7avPt
SYJSP7M9QWkDfqsVKdV9R3sNZzJypkAaHu84r9N+TFbilRgO1+JaZzgjQZtWBi/A3ToLktTZ3Dr1
sLzkuNFvzIoJyWJ50qf4MU1g2DicUM4nQ/jSLW7o49an5S6sl1oqGGZahmkTM33teYPzhSNFEMma
1YY7Yh7JNDvoKetHXsqN4dzgFw/p12fTQtKg14GsVywSlrZZ1RDBNNA3DePtJ2MUnb/mp4bcOBxX
mVGzAIEJU9JkR62uatuIeGG5Xdjau5Fn3w3yGw9a0CMI2ymTfWMA+DvwzKoNbrA8VW9+grG70Vx7
njyiTb4vnkdiKujwLFHBUufPHQkGJyrUGFZCjQR+6fxqvKBESa7fnPI3KUpqF5wxrgYqNTbkf881
d37uBjdcuy0W2T1ULNPLxOU1aBivFJh0e4REQfB2xF183M5Jk34U2at/J1JD9Oc1Y0rApo3vSXqm
36yGKahvq2zb70fAcqwiZ0HPEXncL8xlqAt1cTcoMaz3b3OsBes4+9BVZY1MXy7j5p9y741m84oq
v8DR2g+r3/+vw7jtqLQNdY8LtH4k9n0pG0mzhV0aja4Dd/+4S9YvdtDUFwr0Q+TnxWAwDQzub3qI
KO6FPn0fc8Tzv9cL0zZKQPBf6r1vHYaM79uLxTnNEl5rn1KUu1SzpA1BcCVq2hpNYRNQ2Qa9zAGl
OJORSy/3Zni9fswI5AmB1RQ6RYmW+FDjVZr4VROIlOtzRJBvYjNzOWJtlZga/cvL90uKTr5Ybtqe
Vdff7KtUnG+1oEBcK17w22TIL+JDl9DQWDOOHK4nvlCcZG+44fkNT4pFUExR/libnO3exB+YWFZo
Dew6Vql1GuAMdsrnNORklxttyOfhqcmZxCl8m0hg+usBqYrczDRR9/kxieavzQYES5FoTzsKB0Ix
Cuzkgpr85kX3YvnRxObHNuPyMAntO43nuHFRAm8rFUclalYhD0PWqKZYav2wj7mKKXDVL1OwrIYt
IvoW6w5IG2fzO+RY9oRSJbROacszlrtawHpeYSMZYHAj62UHJDnEsJ9tkVqLs3B66YQwuIce6+S5
Ry+0G6EZUndBZ45vjxzKQ/Ew2qA49HEfgE8RNNZTTMTpsdJUzX2csNc8zAkEf5lnxw1b3gT5WfHD
m/dSOiPA75MDY/97a89BxrC/6w7H8q0vHH2QWbEHQDtC0D5zw6AfggjG6fAxzimWckmwdoZuV91f
B/f+N50uEbj4G5VLvA+sIO8UUuBZho2SHYRiY9YmxR3oMy2BAvBgrEBW1uPFeA0O+jTLMEDdfCJF
g8kuH3PtW4G06bOH2JYQoeslYXks4JQgAzaBPQtYiCotQlHBm9ztWquABm+rmH4+Xd1pZ8fhiweT
Xq9DPU+cGe/gL+7dXaCoq7Z3CgDLWeoJ5QxIwa4TWMvI5frFlyn1v/DkhowZkOKwCsQN7EnhNQ6Z
H1DBIss7kxtAMV9vCXre/y9xMZ5CRN5S5Hh269OVizMiU7yHemx/VPSFmf/A29WvZ/sLHMt3/Ptb
nmcY+WcCcObUy+t5AhiVPRKUvee13JWO1d/i9FwYqDhVNPyk64ceZY5uJm0zzkB0EIbX5oeokeR6
AHvU8snj+pXTm+mqPoCjNvGbaipnP4H7CqJbwb06WsbScBm/o/S7GuQerq21DBMM/CrgXGwfRd97
E7nQOZESiHcdBNtzoTNMwNS2+cdAgv9SihH4sZsJuFfaEEWSHdvajq6/V/XtXD+nwWxkZabarFL3
jH15yTX8gplvXxSEa+LKwnHDVZI+d64IToBoJzwCiNo82TCuMza+ltwW05nVDVXpeF2kS3dxec1w
Dng2owe1ebFjArHYXaAxXyw9WXOwLbsnNfVWKWuQUtQ+EpYThOHrB4BqewCkTZ+6EmIR/gJAEEm6
UvMx/52A9sG8M4VV9LcuLG4HeY1iDlutp1pmXC0ZRCMwKcMooxlMxqHEQ1KDQv8oD0xVi41LxQ6r
aqH+vHL9LHIGfAzMraxtIs6u3By/gc67YuksUnxCvIlf1Hg5qRQe5XoZjJTngepgPKj0+zzFC986
SuC4/wj9rEkWYk8BaSlc1ASXS+RXNBXkvhgcE3XoAQgXjis2ucxMCLfeozljDt5SKYIR5y/lei++
JjEaxa4Zsw6hdBVBuU0cerbCLEwu4W/8KnszGuCeqlh22qO2KmLAHaiEJxSRoLbptG2DZ1E6+9Rq
MzX6aSzDF7XT2EZfKmOApW2CWQLQI2/lTQY4pjXiZAZ9SQMcD/sHvn6pB6JXkeeqz9lhtnMQslxK
APqY7N8kZfhX+ttROqc8nyG5YdqspG8HpqN7jRPpVzsBqbQ08DCUgcTHcW2qPG736TvGRfqWKjuZ
FTKmtZ3euzUXKZAueWporvwl6dJexMm7t9d6dsLLs2MVTBtewnSJLP21NXtnpawoMHzkWSXYfHtP
95cBhZj14LCNqGZ13+OCRLDZPy6WWjOLjn3q81MrA8Furf9SYf7w5RA3GhQFjneRWWwCYVxQK32a
LnX6P7SMpCNxeNA9QQqSc9SfqFx+kTZ2Kqf+cI6rpuoQ/nWLs2psXXqhjfwghuY7gRlDqBuKaXcq
8Evr16lXH4C7VoY8zvVBw+aSqgyiLbgWtNff45WH1ZQRs4tI5txWS5ZmqRMX29RzqfhOghsUsWOs
6CCI1zpAzFoCv7VxkXdrpKizmlV23vKKmK4IquBuJbwJZiNaqyCZbMNQXTTDRlRmkPxzNeo5qdiP
Jmh8llaL4ZtKa1bycIvYseDKSC79rJL+n1qOoojBkEwHTJUO7hq7qX6F/kcokQRv9tApuXowd0kU
ZoFxC6eGKKIt8cQOy/2D1BKlJ7romoM7B7Bo4Zf1QywND5ulACy1GFb2yIrH0A1+4C8WY9MSqvzF
yP7ri9jpwVi2nroKrzPsvmeg/LtLRgH3ly2frETH3iwstNoJKvV5FqjxcoU/UjBFA9cXWYjRzUhc
HHwMNmUUAK8moL8uLLDW1KrMQwkUk9yvo4hKaVbnetFQZw5fSWD+iclbITHVCLVNKIRteBPHEH3x
xXkWpwJe5Qlfs4ER0+DHvWDlCLOP65VwilHqiT+vq8k3xMVwh/jnS/40xtcleHlgwA8DTCskprDE
8YPZ5LUai3ZppzHpSbM+rhluSABfeNtwBbER7QYg8InFrbli3SiUbGFKjvISVoKhQ8rS2QTQTKjO
/P2vmnUPyaZ9LsNzb6cvbLruRERd+k8j6BmO2IHxRobUvRo6C+2lNicci7fvbNTwqnG6Dj02zARV
hXp7qxTPkv2O6ekvopC88WSLUzoi4vhMEM04i2zS0ZTRvcEOXPossmppUkfrIPARtONztPjOLi6s
3W4cdYRk9hPQKwmJr+1wbN7g1HRLNRU6XpR74L+0frKHzrkRiWK6yMhKxJ7wBpJivpJC2c6n3R9O
VNLXdrP8GSK4H3KbpBb/Q2jNtdXupM8ZKebqpCCtsoFNaOFMz0llWtegc72PFtpaZsznfc/Hi8iR
S5VmGKo/0MEFnpsHQ8D5ixVTxzA2e/3a/wvmiJePD+Mwis2wO6fPUk+JyG3h1YJWcw5kplaNL0se
+M7RWCjPs2couUN2VKf//ut3uenQUR+p20MlfROUc9CVtthaAyJtefidtAyN2sspGlfiIu0utFE+
EJvNRuNKPnD1Aje36L0Ug7a95QYUnf2BrS7Syca0truG5u1j59gCDdlEveHV5olKVuRH7yYvz1kq
wKa4UqyOqVpIQFpLkRu6t1Q+PK3wIEvqtpUp/UsGH80ErR82aEvKP56n89LN35fvxXJ9GdRIVuND
WCgO02Rslhr/9kRBVuLqMO4RI4HYdLQDLdqeKRIuLoGGvSgRzGpPf+c6w4A0lqQROAAXRrbKHQjs
p82eNgtIJ7yM4cYgp9DH6FW6b/Qk1q4WYtvh+U7rlg6HjobFeyGLlq7BZwiJaELCxEk31o4tozl/
BckRiasAW3nK7+/3HVVJQVRpHgjwKDbKNcGReRonhySwxEPOvdz3+AqX9WjOgGTGRMEoX0kUpMio
9CZwD5ysn1jbQT7NHKYuwinHcpY0eRbbnaX0Kt9ASQG1vrzk2/2i6KiSNscqfX3wAnj5GvtRQ8GK
Ny5gZT7rJnK0wU9ey3SKFEY8zG8sY9E5jHuZN42EUNLig3Gs6f+/HGF4V5JZRGNvAkY5dPBqPdBZ
S/39qiiGs+Nf+O94JMzJkLNMqMq1ppPyZQW/AWw5ITmav+qQSLY4rdSIXDor/WIM4mNKkOtVPHbW
GTGa4Ekhpfpe2XZ8ntTtHRVo2hyJj78lODsEstt0OXu6yySa80V/GXi7y+9JiRQbBt9CqBsZ8ZeS
gzdHHXuo2OR9AupuLiSBgWDAOzweK02uCK+l3Rt/F7svNampzpjMxDaENr7WnV0PQ17D5Wh6r62A
JL7wHX3oJwUWBynAzDUXCXrRKdmWNl9zkpY57cwFYIqcF1F3SJ85+QB0fzXNBo3dBsWR3OKzqGaC
wQBZ0c+JsEFwQSoXwjZ0n0e9K0LiCexEo8jSTI3HRBxbR955XBeN4kkElEpzAGtFVdXg44FaZ3mC
s1WfRlQnwLyDqAw1iV4QhLkCkskn0T3/u7xt63PSB5HbNpN6ZB8LWxX3K4XiITMmeCGduB2XckKO
Yt0mS02yyIyZ0erYGLhllxEgfGzFYfUwDtlyBNUQAzFhC/nFxy7GDxyg6TQwpUvsWCfdxZFEDCZt
MEinpYkt88uoSLBUIYI0YunDdAZIicbpnUSJM3knJ9nNsM6/M57Bvy+Sw3RZD7QKYktpHCgxuqbr
tw1yhwEV0E6UOCaOvOEv9g7xb1cX8g6pZ8ttvrMjP5wXmmFpwGKZ4EuArJ/BEdS3i6uM1kbUub+1
aveG8fO6TQKvYrZ7RMdNQapI5vhhTi0oLCSHw7jNEa502UNWgE6cpxkl7BRdD8MUz553eRF0p3gq
tXLs0mI5f8Pz3v8EGzwK+BhkkN9BwEyoPuTD2GJ6zE4ZwgTmcC8g7tvk0Nj0aGEHzfzEtGKU43xL
wXTMuWyr9WMJ03483o97WoDXWDC9t93OsOON/+ldMTE6pl9o5PEss2kB/tUZUMiupD0hQ0jLC8Tk
Dp8TaIutoAeBmRXh69boDYhgsDP/YselDJMkzp844GhdeY8bdYylIFqZk6Lq/ebmUzYCSKfd3/fq
JdrTxb45c5l2CTLkNq5Jb9QxQZRbD5b160iBiVWN8cmmKj+1mxDVajMYb68fYYENmGIStLVNULOr
z7+SKfEXWVkB5zVKbm85cLlAbF/fbOQh/41ddFw6RALw+XHhH3nTYjesbr4OrZikFu0CDWj/ck5C
CPSL7OpnhYeye8iFIhaijaFaqZQ10fjxkbHkC4PXv6c095hrf1ZjTlw8RT+LbS3WXoVv+ABsMIVg
SCUu/sovqlOfhnKOEr3acI1+5xuJqBmsIJ0u4Bh/nX/b1IZT80BbJGv14NMNyKwsabXcjfkHv9nu
lmyTacf8H5IosE9oqYnT47j9m/eibKRTRSVIkj6DC8mMMvwlv0YJb0+vv5UPo4OINXcSi3/nEzGu
tEq4yjgF4O/Y/20lFPuCzxDDrqpGa9gpXSZ1w0OPBICjmoknB2NTqJm+RSmDlW/gx+i6i9Gl0Twu
ssju0Tm5Va5mC23aeLoVcULpLhf8KcMIe843WmaDpOHKhW3OWLnE/rnYeawDIiOzpSVe8DIDyELy
gut6wzTZm/4QgGfLBgUKdo6Y/WegP5BQR3GBV5NvB+b3RHm4zbMSU3JYIG7Yk93wpmZW5VhZclE1
3Xrp7mTsKScnsBx7tPiuGK+x1jhdKpHeKoGoJZzhoD13kYOBh0+hBnF9rlWxAx+ZRYYX+/BSKpvS
JbFKuehD8VJgfs0+JDB/Y5eCZGY5AoceHk3cZ+MdGLMaYsB5HjkjHyRZVEo0dlWImD5b3JE0ZolO
ufu2BnMjT1rXIcINnWQSt4ch6Hm+PA6C9wdonlBMAJSydveDC3EcoCdG0eZoL12SUcrTPhDvyO7n
ad6Nh0uB63mU2TsaDsF6CEPgDrx0dQ72q53GwzA92b7cvuJUfzyIn9fvVqdIMHjahTecA080ttmG
EcYZmYQNZsqh/yS1g5bdPnQkMcCpjYsKCX8ymSkAtsO+h3n1ZdAS5VAiU0On3CpDaiRZG2S07iYL
pw5n2E2i2g3tzf4sRseKIoMMowYvTYtikf004aS3nCstdXeQmU0VbwbBqU12pnKqLs4a6qTknii1
AeEw9PcNMVR0zd6lQeaOKnl9G1LEdU+db5nYYV4HFR+nFf5zibv9dZs3jHvOV8FHSxVV7J4uRo+1
Sj8s7LLCBnNaYSWuNSr2/Hs2QKxNASxTjRIPPrbtoenu72ISQCxuEff4BDMcqwFH3pqEicABGyOH
5i+cmKP+Vwh64e1Rj+P/bB9jqUCBjBd9VhTDgw5NsDQpg85QTUfaN/B8g+en2qmj+CbTuD2OvbQv
AzyzweOzPiAhU9Jq4uZRwXijFHCLxiF/17zI+YVi5vSJg9oSb5OFgwlE+eFHhKBC19D8+6AOYLZ5
dkWTs05cH8ecPDasPuC4SgEmOj2+tmJCIdTlvKedk5U5ugiNQcdsNktq/IP8WbSa2QHKZUgNphDZ
pPjU6+3E9C961OHEa0E1RDds0WSs2sFWschPUj4g/HyykcJLtetduR30LPVzm+1pfDSW22GovzGW
btPNWyf3aS3XBqbFLFHoFrFQ7I/4M384cDpE4r/dDD2QWvbPaUI1nJLlv97JXqRHQw1qkqEyl4Kn
jEH/Im7rWGX5UDnwc0D1iV6O9uWAKSQI7iuwUhSCFPTYewpe8rJt6SHIPYVH8Ew9pSuqSZVWVjOp
E6bsonGnnLtEJF0h/x6JbDz1TpPcLk3Z1QemDAa+5+JYW0tPYZ8CaM9YsNhY5SO3CDdoM4XruEpz
hFlOaSHrC31dV1dZTY3Mg2v3foFBG+7A/tBxzfPZTJakkPsZKBYEov7J/sblXzCa4g980mXmffNr
v12AcTYcZXn/G3fsGMBxKA3k5C95EddkZVh2HR0vaD4EF6LPTYSn4TNzV9WCzjqSYFO286sV2AtN
QigjLTVpv9GFzMjttwsP7r8/WiYNwv+dryPsyQqe3fgR785ZlajxzhqA0lxPOdvLANgCFsCQelRz
94wixnkzTYyv+jlWZbkdME5/F0tlIZzkzvvT47HAmjqg4lSSwQApDvhAMDv6TYJX9cu/6o9JKYup
0Sd6Ehch9a9LeVz50weLxOzuG/xX+oBSi5RiZ4TtsuJI9o8eULLQMkDNcpCX8RWBcRl5XfFyJrCJ
e8kLLkUTfDEf42gAGfOuqI5JVNr279jjvoKW9yV1mNskoOcx6JqzAFWVZXPhyacGDbewzkyBe7Gg
rJuz4GWir5e0I0RH/cDvVxsb/ql9IHdsUAKibj6/XQhToGaQfdwsCgpHu92gNEbLycX4oewqdBUi
Au4qmEhUPjpux1G/pxYi7P2AJQY9Maspxyj4nVDGYk+tQyW6xF6XwdCCJuaRz+qxBqdj+CupbqIf
19pzCkPKbmxUIKD0Tiue/Y/N/dAOLH3wT9WFS5pfAUDDP6Sj+jC+63TOYTbhC2lJKg13KStpCcNO
QTJxOJu6R+gNeLv2hB5jBy+YOWTsLaX3JTiMHMMlgJQ4wg1N7g6MmcUslgNf4bMPTtdGpv4NrZG8
hHyUUqnLXcf4UF2SdulvSOzOnaVqjGpVhbhfm5aQt20gtZVn5tCUsR0NI7blhkzwtfZnkInI0LoJ
24pua7CtYEMM7pLyZSy21RcFgKiIJTOLBHYWTeJqdKaAUPMHmworS18IvdsifZy/sz3tL6gLkd/l
N0ta7FQrxzi31wU3FTqBBQyLK/lNhBUPpAK3nfUpLwT/qgMpiUwYCi52o0BDpGUjaa/SKrOonkKL
+XHqER0PeXSwJycTUZ4SziM8+xJF4LOrwsc6u5tlkVMVlXK5uNn6hjgpnhxSJjYJODvLDev0q34y
+WBQb3k0qA3hLO0TnOc7kYHy+9s9y/wRpkmgYf/sSoCIKBsyfhdrf59kJtYX9skILrKoaNAfMBNn
rxkQe/9bI6PMRh0P37QlUd6uJhvokd68Uj2YsG1hSNRhMy6nLxg+4VFabELnDzadX67GA73G3IXi
eObzCpbhlHXcVwCXugz6HEJAHzr3FciHFekn/0sS45GUm1in2nH3iFMStCbIM0qTaAQnqMJHuzSU
llOZ9FwU+G7+3EMvIHnsAwlLWFYeqO6ZRMrRj4f5q819wXGWbcSFjVG9BB/w6JIDYfKwxlJpdy3o
KpEnS8GtBv+cZHj8H/op84PYpyeLebCty7CQBnyV5Wf4684j+XThci1CD2KZyHKiX4L+q6+2L1az
fpiIG7iu3eRCRqQ7oFNBuYiaeyWmdsuI0iFTy0nLvo+/E+VgF/2vP0uiDxU6lKB7BQf99l2Y00b0
6x/6KS0/F6OFCzA5bgMb1ZQVee7MvlzpCUij+CcSyKAkGWEPmzBz5T7ZHnu36Awn7d1Mg6t9ot1R
7tQfr07QavL/2HCrw4iu7lxLjuS2GuLglNes9D0RBGBhvI9R88CZprsYzZBW/Z+de1uCEtqWrten
pXUxsKuIKncAKmNEUp+63WuJQO0vO0Bl/hA4TXcBjGwkOc0rY2gMe/nG/emXt/3Mi/d9X4vUJ5m4
viRrB5XSoI0Ws77RpzdWIjd5FYLYPJm4n3Mz/2rPRgTsFVwJuNEeNCL0Bg9E5jAMq9Z37Oqyx+qA
xdMNn6jFcMnYPIV3SVXfrg2by/WhpwLtvnb5uMpMkGyHmzaiX0S86CBH3+OjcOBBOxhEwLuG5cV1
kRLMUGFf9uG0/X9tDVJsB47t5FW6ks/SVy4GLkB6HtbLHJbcY6e2lQvQV+PFkTFJHf8BRkI5zgfB
zFr7C/eGz9Vb6IW12pbmRCwhpbD88DfpCcZFA1mCm5Alpp2cPwELqKsgKkMiCvk3czY2i13CnITU
p2LSBx4KC0WBrMBU6XlATYwZu7pUysi/vEm90zuhLIRnmCy/3Am+95BbwUGhGyJRrr3nnCyvRhmM
xGgG2b4v6r3zU3+CgTIuhVCTQobD5JopUj9V+5G7lY5Kf6NZvRDcqYIqkEApt07N4dzlI9lv7Kgn
MeMbzzZm5LJ6xSZfOZPBsn0+iGI0ybIDAvX014Ndlia8f6byGErXOGZngxY/7mT5xLzrj6VwXZC1
7Er6KhQ3iILBkkUQgiou7yOQO6H/SftO0YTt7rw5ymC7sJzrqw+zTVtlzI7kRf1pP4P2KQZIM8it
n/rb+hMVwe0Hz11VCyjufJkIjWk/w+KSMhvQl6K0O9/J4xQCzeGo6lI9ISalrfkB8JvDvmL/v88Y
7CqeCjsVRFrfAFfUcYA4NGe84J+K7rZM4/MUQfhXeV0kYaMgwmfd8Mig6PVDDt3RygjRCSJaONHN
yYwlcbysm11HazAIN0QXG2L5oOHl2ne6VbSW4f2FUCw4gCYvOqKNjyn2HTgFDYKJRSJ6edfqXKvC
zmh6XB9DNNVjIie2ghAHSaNjtia3mExpzjWqA8tS7OdV+HENmAajd/+Hbqb1VRQh8SFX7CBHnSCk
CDl57eteGlr3a19BGubsg/1dq4ygKWmjtKm0sd8QJKtUjpvp0TDgQ6WBV2lsq3s/4dMh09JpYLJf
LmPNi3kYEH5S8PbSmBIRnZUAp7CqrXCAlWjJVPq+dxdtscT7umUfxaeIC8ymtw31ixlTfJMiiPdl
2Q/UKpk8mrFO+mwrajsCnxQn2DnHoI3GhgybDC0u+c1vwnwSIuog5Oc9Ta4nfJEyK57FB1pB4G2o
PbJ7cBlg142+oPJTGxuXDBmVMe9YaFYhgBp4e1OumBukyaTIsXf2+V+rCzUtago7GfUeAadgxcos
nD9wfs7SL54LnzQeLBApj6i+WARbM+Ra67P6gPwZCRTCuUBgQMCtTkoLRujSp+YwFbogDIw4Ci1I
KWxqKwzL1jYd1hrPnq3iMAvd3Oeen8MdbeXfFYJwFbLGS3LGx7RsJEiu4qvZbF5RCNk77aEz02LI
xxuZDgUCWm2bVvRenLrGMOqObRv9nK9oKkOAWycD0ZgY4YTIQ91FZinykvl80YtFiSFEM6F22nCj
fw1ksQEDqTOG3ryDV6jz4U3M7N121S98NkKdVBOPfflffoq9lpwZy9W/J+2zVDnZmitl3t44xVb0
9m3TUmvFQBBX/vIGjpEZZCjuVnHZ/Sixm7aENqRm5UYQ22y14rMiVRC9tEpBID60xktdfH5KzeLC
RbMvBUSnEWBG+XKrAQrKru6RJiqBRPZ7zGkcr1jjHVRLJozLObM5lnId2wY5ogFK/Pn7Ll1MC/yW
V1a6TGZ7YzmAXbCHDKlvjYReilhHhY3tU/hgUYBzJ3YxynA+A85LYfgin8dcHnPoYkE+UgyqAtTe
KV9Z/tzplbmz32eO9DpqGyUrxQR25egjAi8I74imv4+310w+0OxgVQgbn+LTOVRN2F1SsjmGhYTw
JEgslI/HpLZIl0w22Ysr5DcmhiU8L8tlPh/1jtTccioM9CHmnhtGCYgkBKDkFJj80G7sPq/Xt55Q
ZRZkmcV3fs3kTdg0OflTFDCgvkB+kYUxBaZa96Skn8FPHfoXpz3sMmbayPDIjNrv9eMvCIYnD5F+
H6DIxMxmUoYgnNALoizCnHdTSSuhBuo4xL2v4UtK+4hfJ+mzmGHWbGpUwgoB0FjQHCttMGUC1WzZ
ZE54TUbtrcglEeUHJOpEDFXW/90cROPJKeYgeklxPQDUibJDjqJeUN/J00Skzz11voIpqcnLF96Q
u5zeFth23e5Uxf4eDg6pNtKyV2zb5F8dFX1nWreQlPiYXDTGrN6nT1L/lJ8AlFd55sMn9gH9XQHs
dpsKDY7K0MuS2sxA/uhMEGL/i/4jwQQyxuqeV8iOYWwTiDJ0tCdEswIr/d2i6aEafbtuAS/OW9z1
QjJryl/hMMWzgXNPOIXs8qUi3a4PwbqpCCh9c8FDSqCNJglzlFgy9xaSZd88jmM0Fc4CaTBZ/1u+
bjzQIR8NhNZvaGBmqkVsObfjFIztj8vq1+wNmQ+Jhkxsf+vRuXVWUI51lm+m1MkpeQu+fdbii/ru
3MNqkeOwnN0djzz7wg6gHzhId/kdYapuVi8itMXTpQvkW8iuStGfVICrReWPuHl9hgP47hnMuJPF
kcICkV220OkRWbZszOi/C0RwqIFNZZ0FCAvv8jhhKv5S3p2wDkKf0aNdZL28Ql9ps9tdUYOLfCdG
r/om4tvsdjCvlgMEZxCGC0e1Gker6Mklzubhduxx7hmjSQ/QcU0m9W9ocKeQsAOrcinMpmhaCxuV
nD0upkaXwFAboc+wY1L45qeXA4pWEFtICl78sTp90/3Aq6ReNldhgoSxBULTxNY/3c1cl05qc3Q/
6djpHfrkE3ok0h+B2cRUku+tw3Ep1wcRD4jmggHfYqSAm0ClCx85rEWupXJKFkTunMYxb2rL3cvJ
SEGGWKLbrYL0/mUcr4vSqzIKNl515d1YZojGRIb9wPoAXDPkUWCoLkbNA2ZDEy/7C475UIptFbLf
KPhYqQe5e58m+Js0h1Ng05FWqSs2TXiHpBO8OGWLiY5Dxpo0B6w9VLCLAHVCwqKbU5o6fzPZW0Xu
hK5DPMDU0z9f1ANNqcYEsS1CqpQYQAd/3YaKvjlcSdUMu3Efi/mYlyEvAZe4kwygYIQ+Ao/0clA/
fdheTUVCCmZopQOsdCEZNmu1lV+1oPgtBDDlHDBUMaMc8BfOpHCZybaQbIxKi5pt+5OeeWizHFhE
kn+77iFPJAIcLhgB3OGwRgGBUzJeLuUrQznJAHaiajF9ak2h+RCzSwCPD0KriQBg5B6XBBqlxdTT
5w97BbRHXdZNEkQLw4sbcG1AgUAzGnVDpuIb1NnuV4ER/4tO32W50/iLLnb7Au051K83r6N1JwNb
jJS47YgNzafUS6NqlY/lGoQvow2qsF0Ap5cwbK8w7F3kLH2Njmuj0d3pSrxPgybEZaqejQP1TuM/
mLtMbbp1hrUPDhWkTMLvqZvsnPlt0aPIyLx24qlIrnMzQopofKDnEjz1m2ojmO6EQFTC8+kfkpRj
Eb0ygNOW8ETVLzvQ1vcwqaFg8skWfvvVQ+mKUb96q/542u/mP6NDTr8XVI4xPBxX5aYejVeqVqGk
sBECQocgK8BrdiIOGV1JoPXGIkOikY8CQ3tYDZCYPRC06sxBIbdB6EbwJHMl5HQD1Ebtv9ywcz7Q
u1oPos8F7Gd7bXvSQ+LdtHNIdom8Zs3phl8M3TwIQIB/WMWC+DVuKZRAjguQ6Dhufj4tjLGvOcNP
TZCHjFtxG6bh/5ObHYdw+rEOep6TyrRUAx4Nrgjz98Ewiis3eQ6iQ2yIDgQwBb0rGZYdYIE0Pn5k
70BS4WKyF3dv1DmN45l/wiAmuin5xfQrXZODOYIYfPqpJomS+LUtO5I8PJhTjP8bMyc54hTJpoeD
I4aXF5Dl7TVN664jFom+xXZveVN8WykoVpm4MKFDsDRSczd/jd5FfNPCj/eXYdd9BljfrEXvNzbW
bRlcbV+YqDvp9B4HUYhG8gcisXTH3YshhP5hthtrCCYO+vHKg72gtPoRBzRd6Yq2P4GmNukIJCfZ
5JB6X4wMxUok9A8jionM+Db4dvSg/eEZHkTMZle5zreyC6xfiA/J/rW7SZXk5yTTOaxntfu3Rd1a
D/huT3WOQUshq1pPB/ZfgOr1dX4A6nVfbyByWYwYaSkLhgjlqjz35TnSNAeGVajqtWqP6MUo1oq3
5UH17DT2rdMh9UG0JRZUlmUQ7X+Y+jJw5GY69RefqkFy4aJGsEhPuafRRYTRxXHsvQLb84uRp9hm
nhCrFs87RO/IDy4b7ng07q8SWvE2elPeGK3R1pJZTW6BTSCnCVY12J/oUXpGASXiEpfME5t3/0Qk
Vwfm3DKw4wb0hpBCQnR8iPqvJL8edY3uUMVT4yeURU6XXGPWVqlabF9Nu8Nucm94x4ZN2GyvPfeJ
x+8FwGcrKpImiDSOSPQwf7W1pZ9MITkkhg5Yga5OdUSpiRWSuggDAH3T/gKLdTkKwQ3UrVOW1GMq
2pt+CGOad4jPqkIDFv1yppKXkYwKf51wY7rLhBp+WBRtON/SIQhOshbmCvBBJ/INCljaBM2eKAp0
AjyhigsGZ0v/T/Atg8jIm3vp0yZgEiulJ7Viku0/69Rjh6BZUuhBiHRz0JBWy4iVzGdGsyhgxpvc
8cVJy25KOY+ksmkMuIsOsKvWXT5OSc+y02ukwTi/XKEcNLnH7W/U4SpQMRGY02xEURR3dt7eqSIK
4dh1kx8YRqVl8wsyV/WrQnEzMBb/5NRw2fky53esAT4A3UHL9bD8UdQGYuLIOA0f1ckXVNvQ9dje
kVUMb7lx87y6l4gPvxBQbURkNmBzLpbfwe8q7Ld2DZxjyxZT/7IBbAvx0tvRk8UNl/565A1zeNbF
SU6s4iFXCprecqAdFsReeJNlZTUWzFlD8U1KvCKbkqbg9dD/StjQxcC3YWFT5I6fq3U9NgMl6mqw
F8olVGMDQsxIWv6ex7mqfNTZ0byc2n56bkqaK2M6Fq9KGFZ545QNhgy6VdAFtXBuSB/vdnd2j9SN
NIwJ7eO6qvb/tpuUh/zsZ4oypWi+0won6ohoacEAU+XpFgn1EliMFCQSAnegUMuz8nP5Zp70TXAr
kui+XeJum/gGxlTc5gb3c/R3VYF54xJOOnV78ClGnmOkUWwC92CrCw3R2rlBgfcewcAv90Mk9CmA
oY4J4s8ZsW9wyj1m8Q5pBbFLbugyKgnXvPDct5n3Plum7QVS4MYg5fyiJMy2OHGTTLAS9Onnm/Bq
OboTi4jRVtFKmeqS+c5T9AwEKBO5ROb7aXWv4U29mU/mUApaWJLaXviBdtxNY6CLyyCilcIHtdii
jSVc251SoRPLYEtxjOrpYk4dA4WGD8kHJI144xEjAkZdCH7w/xWiTGOql2I6zxyPTkRTiQpzXo+I
dhNujWMeyEdOqxLfP6nHtcDdMmgm3cNH6d6oLV/zSAn2nlvyDqsS3S11g17NvzPnE+qd6ixyiZ1T
0cfLzgEaE38rwh0LW2PAlwwsvFduehS35YlgNQhYMlTdAxI8K6D1BgKxmUZJamacnqps+RtpeLkp
jeHPRxQdz+sbzxkMtpBne5w0kVLdZ8NEhyNMeDVvHnwXNHJUkcJ4H65R8SmDi4W4A4qLkxC4ZIYa
twy93cAGwMgcAv0GnvXYh9qi9x2d1u+Q6wuwCf2FoZbLBXD2sDffF2/sE54ibp+Ugr7+HelTzW0u
mydRak+4zDwIdWZI+qzV9JSpY0lNFAtxi6dXLqTs+1fX/kSqZGZg3nOXF3NPoY2Kv6ET9WPaHVSA
udZDWEnnwbyAQljGgyrVhWDVNNrmSvzHkJD7n0KEjEKMyXZUHhs1EI2GkcfSWrvo31aqqGujPjrn
7JhDEwDY+s8Pow493ZvjAjPLhEVOUbdTp88sMuvtTbETailF7A1WZfjL8kVqUH9aKAVs8gBVH2+O
bSWI5MpPGbYOfI+tyErtasdDsi3/VPKx7LeFR4C2fu+LU71QTzdKXT4FQDyO9GKnoU+MIHE/uD/o
+zQw21iKtIPiiehB2x5Qqtch5YrLHonLn09wtL9P7rbgVZy0HeZs7h3IrG8Xca+Ao5PV5q0naq1F
tld1lTx94T2gWCy5RnwYv6xPCBnrCl0AB6EWN0RZ1Gh5jfJxndm+Osjx1VOoqCYnEa0PUPbK48np
f5AzHiI5W2cch32ga2iB7qUvxAqtrv1EIHhEA4oFmZNk4YA6TvMJNfazUi1cX8YEgPOin2pjUCrp
QlW8Ty655v0zCIm1grcjfVr6Kr4b+M1PgX4rBAJOmnSokl9y3Qg3EQ6/hPcOmKghQxykPn6ogZel
CCm0lAvz5Toy1397fcwqNsmA/q2sKZOXy1K7Vl3R5Rw6MtTqmkMZVpOpYXQHCB2fvVOp77E3IlxQ
HVVneQCT/PqYZV47c3ZHF2XFJqhC5Kn3n5CZych33kvnnIo8L2ddk7esM7+ZYH/k3WREmDjiJ9wI
7c8opa27fx1/WxmhtEgYIRUGXIx1n1u7KSE4EqBbCIOEaDON1ejnA3KOr7yAfgQQsdp9sW66h9lV
hey5JjWrSqGF77WPtas9TCXJjoWp73vjP89001o43pqzXUjJNL8yLPr2yu8uKjH36dOknB4Yif+c
5xg790yyWsELVq9nysMS2UiFWebuT6qYnJke9ojCHf9SwEZr/wF3tsb3WvtClHD/O73trU+AddsC
sS4HivulynXBgSJoDy0cz0LqcCqiakl6YKSEHDHC+8y4M4l/m501i8rt2JMjxDS5dWXxR/3ha4AS
UZh4NhRdBBx854SFbs2T1wEsaq0tyBDFjrWOJbf3reVFHgpAqhKn4spowHJezjaUZqtt9x0KZWwE
7p9gjB04FpjOOtStszB0RmFINaVndp54RxkIFDb0q8LwBPwcrTQ0hLoxJbSaFzpoURxrniLDNTlf
QySSGAIL8Fb5tM1DhPa/Ki89t6e0nCjnR+isL1LacRa6qQEt1TcXpF8GuKB2jTeMvYY82b7WNyoZ
bp91BlifAGItnCZ5tnJgP6FP8zOnOBEXnTJBuY1KKV6SodsrYgj70GeiXlymQfmZmWP+tEza6AGa
/DubUASeYZtUY2CRKXbgVp82Tu93aVoHMY9fghUzsgy94fkZ6mAkpXnHcucdBjz1x4SBM5Ei74GA
+b7YujPSgL9Gs+k/1dAgrAD9byXyhE/hVY2hTDjZ4CgJqKPZyhQkSNqiRDJhFsCe4Ed8knMc8jhj
g5JVDzI+Nat4RnRCiowFUGQMGwQHRAdoXFXGIF/V8T9XEn5vPbUDhfgQXPozxJlguSj0vCMRtmge
pGUsFRVhQsG9N6qbGgH5Guee4+47IqVUuqTF1kHvLmxdb6RFS0LF3cZn42sHo5S1nl6epGT8Pu5u
dJDV9H7wYRbG7J4kjCb4YUxhvtr7KEpN+eGHzgQPB/Df+L6O0jPcpK0MEvoSjbjK0YXeuGbKr8Vt
yOMeyNEIOcaermcmlEDzhgF//5Abcf/QPQpC8LO/LiPULQ/PO+7w6Taw6xLygueS20nNg4EaQ9Zz
W970fBKmbu3CaZcYnAO4LTlzvHrw63iOeJhNKYpcKEj67jzy/R+uqMUDHrLoz9IP2U8bGmoJnjlV
tl13FtxhYmoZrxKNRog07yIdY54qethwB+G7EhWsSPPNkfoOM9ISlCLvlc2RilUodPlV3k74foKf
jNyb9+fklq1APvo6a1faWB7Mp8xgbnUvykNpYEKcJlEAFwktFsMG6OFNS4btpfBuR+KImfjhf+2L
6qzw8aQinp50iE8x9ZGmcltm92GhwehR+kBfi9RchI9GqK+syrTusdD9q3RvhaDy+1ycD2k9KV9o
EePTPl5iHfqE3rWNvFD/yeoBNxkLkE0aIgYt1SU7yaKKYshpuDiuk7/AuD7Xl/O4n5zVvXl1ZCVk
TjFnC3nfsfznz2wamV1LukABRkP4D5r6XF49tMqnPwEmoEGMNb9oA5OVPoFDm0Dnzr3vvTlzhAvH
a29uN1UK11kOkYKDVZtFfZi1T1vpJMCXM0TrdS5ZaEHJ0bpP4tlJUzRYeD0CsmbwCpDAVKw27gs5
NnSFsWanbe2JtOlnRbh46d+1IZcd0+2BYmPwL0I0rPjgIur69lVDFulv1/BNQpEk4SgtGuAM9CFp
1si05fLa4//Aa7XRod3Qa8cSKWT155SUht/Szn9jhe2MZm7hZKIzjj80cGMabzLTeXzihWHkmMCF
EvBhxgO0NJtJIimWRWjk4AHwV4SOQ2Mzi9jXAhaW6o9QF2tLLHB9m/pepb6rEBdgmUxtf2+6mJeX
zosoLQvlNCTiJMIHgTsOHT3v7X8gkp315lg3pwUnlw0QAZjKZ8ZUHwR/l6jrA5nAy/ju/O+RdTDc
E6NMrtc6O4+w8cYJYbRysyoxBLwnopQAbDfn1T+9r19TgQImukbyMAwLQZraO3Ew/rUyQ/AzcHpw
LjHEVk46Xycm/WNteLPgd9GIcj3DUWPCKCq+KnptWML3VN6o4WfVH82etZnCadfoBhm40RFof0Ak
1VtWl7LRHwf4DFTbwHClYpaIj5RxcgTpKQHaDRa9ED9T5+C8YTqdXrAzql5j61tlC108HKcoUkTX
2GOXSR5JsNMfz2R3D0ed59cPxyNmT1cgDweOU4zfwc1QnjuesqluIRveX1aYSd3O+Wdv1hcoWJh7
qaGlYcK4URT9YSScVJNP2sM7XFj4Q9yX16wKu58ZiUZHCkYTK0HGclUk5lOdDOam1c6RiES6MJt8
sAzlGPtPwPH1hmy44yPasJe/fJNWIlaEZ2EYaDCY5tsKzOvFiMwCdcxrMvkgvvBudPvuPVurbQFr
zujO4EgU0dosTefIRQ2Vf6j5MTNe/qyFC+hO+j2Jncrj6KWY39SOV9AvrBNqtZ1k3HoUzHcz9jCR
i920fwXGn4lWkMrbdZyt7bHGh16FOzXXceoiKICZwNRuelOSUp2ZpEn74yB9lGD2mlPdZG6QwTrX
Icg93OyN8ji2jc0Mn8P6FbePThcuedJr7AhS3zJcnDH4mMa7zo66dJUpbtdrCx8caLpffYCYSOCP
NU/OiqIeTCsuTnmoJm+caTCzcE4gHZ/y14JPB25cFCVf45/rqcwiaYFr/u5Y64nUoecmna4XLSn3
7q911OHgyJubXBmrj2b6iYvY1EBvDtZyPmXVJnz1KlkrSWfOFYTFnnFVdWk+vr2YsH/b3COE7RQF
kWCskN7BXYSJLoegfOPUsl2ls2acWjwccF08WMSkW5oQtYdUIjTTDA42yx/tEZ8U5Fb5KF+Eilvn
LHwNLVvZrt7Ojqjzys8re8x6WtbeaZMZ4NwSoX+FATmPkYr7/IAuxMjJD6ld3hVdyFqMeqPka76B
ICOkS114dIubj/xyn08RlgR5NQnmqUIY+LZt1D+Xqx7/Mirs7iIp4OMxbuzQa6LEaYgcklE14NIz
1VCU+3hXIetrUIv6a6O2iJMBrqm8iiANnXMUQdpwy/jiAdriiAnlf/dRyZ4U4rOAFaZq1KDuyL3j
OfFyewjRLGo8MXZuogE5468fVeMX8dirZS/GzqzsTPUBK9igL3uK9aRXxYs5Tfuc3DoKdsksERhV
7pR2QGWGSid2XyttTeu8ZlGWsk16h8+VgAxj8NGDRnNXrYdg23SfEit4A0hxqH8ddtUMvHTZ2u+d
qc/fejbuWhaHGSczXITmLvu/FmmiZTfspMt26uOC6MCYqkPttPRmz8CHZqE294Tvrh/ND2jaYjz/
f3BkOkj5mGpgTo2jfjlXs45s0BYN53xqy/8yKanwtkbhRUk4eLOZ63g7RIVMOPhzDFjA69aKS3Wh
hrtVmI3tzrB+YP8AzdPlAiRlGH8XpIHmYwOMXElaqQgJSXFooTvp7aTCELjuNHHJRKHWlUOt3SZT
YF6gvkEG1C8EGhYNPEZst2+5sc+OmHEGX5vq7IrNCSs5UCuMlkuSjeWUKuOrlgoJ5tG4mvz8vlyy
zGwobAy3bFuf38x7SYESk6cVtUsqglHgosEiDDdkLZW50FhNq/MNZyRgNeaDvK26JsUIxCD14CTO
tBzW2wuWgPmEoatWe4xnI6JnoiLbfEm9hh1aZYA5yf5tz7Sq/zfE3lz6d0ZnM1Q34zfsCu3/alxY
W2d8CoL4VVHPu9VSf7dTqxDReVzZIWCvoNQCeyAbOO1luK4034nLrUPcTI9CWNwKOEa5PYcvtZEa
z6FVlVYYExRnAkp0HOV2Ldp8S1bffKmLYojItyv6gJKqGPwOtY9WWGG3mrxFTtAY6cD5oYwGGgn9
UMEBsVxZlhDHfbHYCv6ZJmebG4E6uAsB1jQ5j7LAInLJWznw1xH8OOxPhTspqBWKLg5O96MH/4K4
lp4nRuvP4/YRb3ScAx5P1HVknlenpCyGanS/BFffnu4+0+6aXgpMJY6HykQfmib9M6X2nf1WUTzi
87/hMxpU3H0rWBu+gs6Dv4DqayPXgaSuCMLCIL/QLCo8VuYxZv2a6VGVLhFSDT02FnFj7Srut0k4
CZ6jwK/uuVNlAI6uRYofIWqyCoAQa1D2p0sLCRpJYM2oedEzep9bxHQNCWClueprlTKCiXj02lPO
QSHbj8JOP5zpIRtnpKgs/ZNNtfrrv9A+g2i8tNsTPwMOpqEI1UWyepd7zYVjRctmEbTiwWEfPzaR
kIGs0Nij/WRI1fmNeooBV23OiqiXwr5dLoCsyCO9zbM3fZR4EcgkyMLtWbnERmQI2YJCp19l+xJB
qK4/nUKY1OiYgR8mqyfSgHotb1KAKKXqNtjr8gEfhrFeyUeSx5be7ArbEvKO4Z8ieTOtAA1+fERw
XeiD1NiEyG6aD9XiPEjDS2PAPp2B60A96AaVgdTJIZhsCMZZw2sdLd9/YeizB03SuWv87xA6DbnI
ouSitL2r9YmfVyZZyuP6ngbmqEu/RaI0gpFM6WnrrnsM5CSzE+gbvGWkXGH+oPTD3Az+MBD18+fH
OOJWhi3TWLq3M7BbrVhxAmC7AD3QUVWKUC81YCAVL8Ejj45hENn3zIS7a4dc9bePRUQI3sbLiRcn
+pZZO9rlZuul1BixVpYkq2pK9r/rHIix33W5FONKzzyeiYWbbq2NiO5rlcPAxYHga2UtxSA252zN
75pbabvc25y4cEIlINa7dScJDd/Tc2F1W/l1ZpF8A79tmYfwtp5ZFRezTzWAszR59vljwaikxOwD
rfSiE1s40WzR5cgeCLGACo5Uma1YKlUKZncAxKNgZTsrU06hSRDwF/9IKgGRmqIurY7Lzy0e+0IU
RIqpBILfA2bQDJRlW1HXUbmSjiREqPKLeK+6N50DM7nacTzOqSpxeDZ5IBdRq5J/Pu6J9pcRP0Wd
MalfeSEKb39Qx+dl9q9drWoH8MF04Qwdf+GJSZE87v6fmZuc9C3i09SpyD9/cjVosFlKa6C8cAXd
iIX1y0pvGQbOs98Ys+2Vn16eA7ErxrLmzds5PhOnDvvO1O8CVcy6TWBGayqP7sHfGl4f2gVM1rVq
HaKVyyVr0gQHOJwEbQCc/mTx6ZQAtKcxWZ/I1LZS1FDh30J1LnjbDAYvmRHPSBSAbTUHFGVbprGL
sgQaw1dsyyf8D73f2SdxBRV0eGZgTES6iZTQgw7dyKS1GgAS8wr4Ny9NtgcUsuN+zh7IZAps2aAy
TKkU4EtEdsPsc90iMNE0FquBnlZwe29jckVKSqgSsIQ6FlexGW/dLy+eHVWfQpb44/j1lQlognxI
U/0BqCPJejOsIdfAHcDkOX9/BK9/v9pDUIeqvsDlJIfF3LCi4rXNECN9cjuNh63rCVaHgCtx3Huj
hUlPdxGtMkLcSJFtz9KIPXmt91IFww6XzvXwbx8FTjUhyW2u610rnI7sitVu0J88IYtMj5fpZ6yz
g4a6SF7/oi22eHibny/C0/IVzuea6Et+8rwz8eMyWUy/Gc6vZnyrYIg9/WwsTxnFkCzatDi73j1e
WN5Xky4fDRnwVvCvLALyCEjr07KlPbZ6r2eAGTIkN8iOWbOOMVxcJrCR2MYUC8cROdgffSqRzkB1
HcBMOtWCZA5GnQzDOxXiusknmYeLe3JsXx4sls5q7vUIVXFw09OaD3LypPvNbclHzhGxPSEkXJut
11Q4q0fO/MfOUwZVJQaq3bjonkNpmU29mhx2KYZtOl+QfLsUTEWg+52eztWsMTVpafaRE5J+uSGr
tS7BNDDxcEh8MalVOxCY2rUuJnfvcnaJwOCGBsF95zKyqVyQRmRC1l4fbssTSR0PGRaWT4x1PcZR
lG7Jqulrvz1wqIhJvUEBl7wyifky15AvD9VzC6vNiey3s5aPhkjDwKeehQH/jDLDn2ALsnkEAV6u
BS3gr9v+eUV9p8RFoygz5Yq2m78056IIK76DTuc3aTbU8AQvOesJqwIuL9zPpx+TYCyXntTVqL9r
18StULiz+QpfGLfX4oCFGx7bIBkVfVhQ3AeFN5e5zW/qZ7QaS6Lobv6aaUzNajWc/C0UiJNyqKQj
zPEcZ4AZ3H4zQ/Gu6FPvw1SEh3drDdo9rEyw96NzUTZUb/NXdoIkN63EBr2MinRIbi6waQBzt1xS
ArTnLK6FnZ0ZgGuj2W3NCu4YwbGsW5lcMzQwUc9AAENTuw8pBc9gdsSihbiXxmLiXipWXoXFtcfs
dpi2pC81ltxtAXcS8FGEOgEGvakicmYYipj7M3iEBvdMzGXyi6zkKP4WnSQQFPoo4JnKcZluoik6
camO0DyfB3+/Hid/JqpR3rm1q1j2V38xNmVAMt4yhGwUbp2cabBgpJuG0HAbrmK1kE+uJ/s2ERUK
jZ/YRpCVrB+BDhz+GQqXnacM83r3JSVA9WFCtuAgVKPBF37RUN5JJ1FLjn8mrXl3JCn4t3mQQI0k
ITWVUbuemgG8TC+LbVitSQFtifsb4Z68+2Gapks4zjOdP5Yna68skCxENkyisMcI3cocpCQsMSTI
nNa4umbdMneAPPOBteMAIsfpi0QTH/gIA7yMXq+w+cwMPTUe+3/ZtbN71t/xhB/8mrntqtNCPayz
HaNrUrDpzdsot0jO9sfNsoef+ND+7i+EjZojVFP0On8eM+m73zY9lBFs1AU7VfEvlFYtIhH3V+NI
Ci01uTbrw6v/L0SUfHIHWxY/9Zr8ygldq1aYiIysSMkniJ1ggVpwpvn/YmcvuG04tKiF+wm3ztjB
bolXWLsxGVoj3oKJQQMY+HIHviB0TzpPfzU8Ku+JhKsGXoKxEl7l+l+GmmoC8gkBRVklHCIPABb6
1oFCjFdBIhnLcKa5POE1Zp6fIhMsNoCC8W6teIChdlUEdknAScezwsdo+zaie4EjzsLh6vND32DT
6m26kT0PT3R4CWhZ0aPRWPXW5bDPEmij7XZVuyp/KEtXWRPm2OR6Ppu0LcX4nIx5zoSPTPtrQcEF
MELxw9YR7LuyEWkmYm2vPgeVoEztHV1Ff764nAKFPkKO86CU2FwQzqf+BjR1tzFelMdtZFjpzPv8
vEPar2E0Yg1/yjmf7Jdj3bPeMYBZG+NqP81MYfWAI2fimmTaWPKfS3YN/RSLs4JhfXO/X+jk7eHx
nPIbHN5MUarV/w3T1kmmBKBGnOxn4MQuvHOJx3Wal0+B4Gna40VL4gs6u0Tp8JHYppi1PdCx9Nsz
NihVgYun/CNKYqo+bh7SFVbEkKeQQ0BlcOeBgG16rNOKp3b75E14U5/5j66hv2u4ouT8c75MYKl1
W2LRY7EUXhhT7X0TBd1onsr9gIXwHKwxJsAVEtuEEJD3BusA1lrYyj1z8sZHKonArdOlPNiZgIVW
O7TGcntsn1w+AI7oCjamjrEAEpL/DlAmcfSH+paSpI+teWsT8LfGdS0Y8s4gk9tj3DS4uhINPnXw
wE2x/Bis79EeWmJmrVeeXn2XUqndntfApHefQ7ok8W3bU6Rvocc7Cf2Zhr8wcPIb6eYuD69k/Iyv
zTFiBH/DkrcNaGNbIikYxsVt0t2AiKoDySiDPVlkwe5lW7DNClehiuEuhyFkpn5liPpdpzSNDJnQ
P4D0qWOZYcluDlAIFLh7GWKRR3b26UYCwUhP5lVJJ12W8jds58bogUBT54ZN93meH/St/kbwlxLy
wUeQXQkJW5TGth85bAnVvmmk++Eeligf6z+M1kU5ACKMdgtLEpnf1h46KEokN5N2bZd7n0ue8jXC
41EXtjKEzq41TTqx3JCjEOso3ixc//9dhXJfd+zv52cqcS6UqQ78CE4wvIe/WKYfK8gMsF1VgOPg
/WGPFdbVw4+9NTOALFiaNofd7v6sEnf0VVQ4HHCF4s/GjPmNJZ0j6ienxXUoQ8cLcipuBL/3/zqU
gOm/iTB6rxAw6h5W7hpNpfKrv5xOTpyi49yDa5AN6/ttyKGmg7ph1UcBSipKnvl58yJk4cMDVUgI
lPeYm78UJDamGhvVs8pCA20dbig4Jtevgq61n9owfGUGrjPwtf3RSBp2eCbzv3eN2X0zjxN+SPCC
dwt6pKL8r96qpUXhTIaE3pMtO6SOX5UZT0MUGYy/aHqu0qufZ+U0ZNqBW2ydIX+VzFFL+RhKh35V
mXR1aqGO6xErL5Ha1lr8E3yqb0QAZ61w13pHRAaZE7GbkTuh8pzB1oR6en7VE9xm6ppV0rRu8aht
JcxakLhBP4T2oKnq69vj9WXqKxp0muEBKRkRug8bQoL1dcfmbLIKkQ6kErC9VuETMAMr+p8L6QS7
Sb+Lgbm9+plmhIJwMXtHz5fkJBU2K4WFUnJam8GIl3WlL6FsTRndtoWluHBjiaBnvUbVbL4IESri
FaHQuYSYhn0JGiKnbtzoF679UiZOlSaeKvo3NWSNJr/QVZ1CI/nG/YHcNcxyIImPf8Jd0XN+uwpm
Vl2ZS7oMUB0bEv6usIwLwFey/hMRDh5NIoLhJIKCnJE8b86dY4gsiURHMos/TZwPeQAKlkdnI+tc
6qFdPTD+wNLM2x0196KAz1Ebou5O+nxoaLkW44L83VRa1hGUOik5aStF05BWdRad5BGhBFGCxuA0
6IGig0GyevUtp0J2EpqSIw3pS4cOimLPC9v6NsF1W4exedjLzo1KET+QiWxMS3YxOuuSklEFQ8zO
FrdjGKc19nC6ZbU0e1ktNVVGOodlnsyGQEDav3GpC31hEiZaHtNK9XWWDGSAwFFBKidUU5mfwfDC
w9WFfncTLJKzXPGZ1dtRWUf8Y+JbMt/qjaZtksoZlUlrZORm71renfzWgiGjZHdxCW8aO/ewovxL
2gq7+N5i08TpAxSaty9sxDo9xwKTy+9nj8Tdrp35qDCq0/A2fWjIkK9Zu4mhzWfS054L+GXUVBvS
/9K4x+nqkdHaB2tfc4NwrVkYz+KBuMeK3SPwMGxQGo5rOkUoONB4CBnM7BugAELpZMeQX43CdzTY
TvsTMdMaedlMc1YWpLZRe/Cc3wcpHObBpUTdpt5OndW/hlpplTcTvDqrFfanoMhR/kDSYX8zPoUY
Jzx5wheUZWnNkX9E8RqCSRDMXTw1sPJMCaISh1BVeieUel9ocjK4w7R6orzDEgEwVvaPr/Pp5Ojx
q1Wus4ANhig9HMAYeTmWQle1MghNAKIBCtTHjiUyHQTg5T9VqSXPfSTZsZyPiJFbL5ohoXFnJy/s
LKz22/HG+V/gNnXdYv14JktvVaMwdjc0tWzcxg76NIzfwS96VMxX922PgfOXTL/QPdN8EfSnbf6o
hropZyvKKfQqpGHvTFW9ZA1ZUKifWytaifOcM5GuwByw9AnMmRzD5/+9zjiAYJIAMjtwy1f04sXe
Du3aYU5Pdu7jei+dUHdAi9V8X9srP6owAtkLGOuKlQqIR1DQN53aZpn0+7ejkRKuw52m7v3LGxMs
AKfZBoyZbliAIHh282uZQuwBZRyg22sDQ/lT+sji+mZgftPvOsibYN9vlIfsmL33ShT2YhzAiFZv
QkgmJSKfC9QI6KBz9jGjuNiZbyy8is49eSnsN8ikk/JWa5ge8N1YmUPKHLfRM+EpRdhOAA6OL5NU
BpnTFqHN5F0mS2zuAcrnFUkDk8+WA6Wy/Rrggv/pUIUmR4KlOuB2pIgNTpYq2VRwraXFmHk5PiNT
HnY4jPThJdDDyjIddgQ7tojUWsQUzQOkbFTHib76XyNd3D2ikthCnGmEGzqOv3BYgpdRJT6X+cHq
oB6AHPGbI/FHGOE65AZVf+J5nJLOInkVNEVBc16az9v2AKA51/7rzFDGk4iJof57j+o3iAbKYj0/
CKVlJIKZA8nFvjbeNwR/4HVmLCAhr/dMPd5DUj2OO1e7n0K0WXNfkOlAsyhS6Go3CEq7blaLKlZ3
KaLh/aUwvV7uVbL0LHI38JuPhrrecVURcailbWTOQq9YLufoJ47Y2q+T3ZXB3QU0/9FQX4E/SO+h
YL0MAbipiM8oNBQ1fgBokkoEXuRqsa0ICNg9lexXu/Ij+Za3ECpqyi2ED7fnXFIvC4h0Y+8yY4JZ
Ub4R+OS/aIHj/9/XzbhzSknoElzEv/EwQ/gl1ZKjxjuKwaI8/x+AvDI13wjTFZyOpaCqAhfrnOvB
fOJvs0xX0Gg3vetgMW/oHZgGprAiZPWpn9DH7RHLnsyOx4Knp6o8EpeW4G3jg2u5LcXO2KiddmeP
WLuiUZCdruQjp8MQvVF+naOYe8p6QRTOYXDIOidVOq0PP1hFB47HI4VWnXNP1u+FKdoZ2+8iPO9i
+uGtCpulRYr4+uHtXlofvkgyqXZSQ0H0Er/TAMBzFl7oJdcz8XbMv18eslsCBFpVluK6pSiEXDSH
BI4LoRhUe8Kk6n9WvHsU+vVRuUHJ27c030UpV9dH0W4NBFzEvaPmntGjHaUF7zu3lXpPEvCZ/yrZ
ihVAOq3fUHykj1uUWfI9D2jyFWfXxtbxZxlnrcx3zs9N59Ar0U9oN+QRHYYrcPYT8gmZajLx7PME
BURYrMWAwReXZ0dGZ98mZBrTLN6y1zes53DgZYoY90h7ylc/G3HqJXZrrM1JJDG0D57cV7ZrnRTw
xmvJCijrG0gG3Na6grPGbRidThWjLOTfCuY4s27Ta6rI6hH+peNZfqh7RurXfre3A/N9k6c9HG1O
XQBT0alE9wyq5oPxWBYs/0lohBSV54aSxW3VIDfzDgBqvCiUKURQiXmmtiUmGQy/bM9gTtFnI+DO
8FuCkMXJatsoeoctvA4Jx3p3XIDBhmNmL2DPyjd/ukI4iWsw8iJjpzr2jAfnRO24XrnvKdnqF+dP
s/Q8zCpOv7Vof+mp18vi9LTxW8MZLx/BVx4DiZq+454lGHobQQ21eTv3aBlzZCIpAZWCREvOGBPz
LOwD8HlPmWpeSI9ojdjAAy+87Fhw5rvj3mLMreANshBEht5I6eWVQ6H21nM9Is+0ztgGeRBiEjvg
JKzqtYCdEv4ifX7IFwtFHlGIONNeCmGb9VvdLyP8ponxGRIkjNy0OEJdIbAWGLGRFxPgB8D1zUxY
CM9aazhD+NWTtUSDQQ/evP+/SfodNWYAk+FPKXuJ/UEVwoxFoyLXI1EsBoP/zA65YwzIp9r26XFI
7eFban23GyUqfYnRu9gB9UjL9fXDJH45YFT0Oj+Q09JYZtFbbJRRJmmPvRLWGB0EgsfdlcMrTI+1
3myz3e7SdpEUkKlAEkCFV0GMJz/n9AEocNOiZ7o3R2FyjBpPX3PZt9kPqQd7lDnhf1gXv4fS3wX/
1HCidfIr7ZypjeggPkOq/ssGIgN+qe0lmRZrTu8HkVK8uhvFLLy9jJQa13jT4Rb47ggYeYWfyiEf
SJs6kt7cUTSS9H6SdVoCxE4pTLVXWvBk+wQc3NKoj6YRbL+NP5voppoUX2P1fR8tD92N51p8+rW3
NIJ+IEzE1+RZQpBvTKWICk1Cm7NlQJdVtcgZJKdVLIoOjY60wNVu/QoW2HY1wZFsbAMYiXrEeGOi
lsBN74X3ZyfEKT/AOYyCQ27aeHRjrhjeF3h1IHdAE34AEfXsV5EG+ADMmqYXRTRH9t2YC/sMW2Sk
oUig8lqlF7JIuYso3s0Lh3RQnw10kfbTJU3YPxuOHNW3xFDatuzs5O1xA9L2jopYvl+jfREikdfS
nSZJyDd9ivTQGXig9D/+V7+2mm6BLNd//hfOxNz3TX43kWZzuH8vftJI87KAa2qWw8TScIcTYfKh
Jk9mWq89QjmO+T/mwgvrUd9tbghk4uY6IAYkK574dStG1VY7HwP7MqMpTMrAKAM6s805DGESSTi/
1wSDXJn4wh+fzM5zYW6s9ZKY5F6899GiQ+9Y9d6uzJFuPs6oShI76wNM/nQQQFLOC/P2JUYLhfFQ
8aCcmavTMQCOdVx2NhjWo3mRqmir+gVPCaJ9jjsFuq7QWMeqMlhIY5DUDh+AxS0Nt4S75zmvZP7J
UkvHXitMVNQFABQMNVL31ISda+O9ior/gNcgvFLe5KOuIBm1VCeP+5gexMX1SaKEN26QXFwVCPFE
UB6RF70eLw3v8uJVB5KwVt25lG8coOje8ygALky1tCARChYUu8ffUAqdxig4D+TA05B+olR/OWvy
KxJSFZ76rVQsn0yjDeu1WW5ekt0C5AzjZxWgz9f/Po870oBdxveOLCGnBL8tjs+zsau7UXMmTooB
uE7Mpi0ROmUVzSDzFrI1DYKdZzc8AGq1zdO+AxdwrqqszKDmPqyMVcqxKS/K/oKUC01KloJ92iQd
qt1i8YhgKpZa/zO6x0uVSlDieuivIs/S97ZS/YDzoSRST4CZTx/0ZXFKZ9JnOxCOYpXUpVKsG+R5
umFnTWcT78+uUCLkSqHXpgrO3cG4fEwLJFHQVIm7IiqISKe/8yl9n6jlF8pUse5vQTXB6oL5T45s
rhUtGziJ+siA3mBRJU2AscUEYj+uM/XaEIY821GLjrPqZqP4Sxh6EcezCV3aSRQg+SkzUw9Hm5BW
RbWNoYO8GUNKrYJ2Xa53VqtWJMwnWineL4UKG+HanGu+AJEJQfXx1w3EsmgBPXcWtl6vdGHvbsuk
ZPBsJxnccfmLkFkDsN3C4S9a7kjMjrGZJN83t6u9+u8dWDR/RJpe4VpJnGSmeevYtB5HCEIPdNwB
RWPvcvrVODab10FrF9ymzNdUrc1inLetgvDouMp1IB+Dkzq5IPZ6UPz5U9mu1IEA4ynhpbQ/zITz
ZSK4MuxLg/IIOLAAIB9eDVaAVgNIw1mD+RAwqT+KeqPNzM+mPNtLCPxKqm5UCL/7WGrBEGeKoLUb
c0QyyC9+yjEg91Ocoe5WEJXuDPDDVe4aw2ERLj2GO4PdEoWPY5OK4v8KZwELg+hXc/l3Yh/oSmtm
SeC1LK9rTC1Oe4MhRsUHViYS9GFr1zVPcdKmDFZ8JqIPik5xLSYUN8rhsBwzGeJ1rw7DxxPqYUVN
LeNl2Kl/gfOqSKGtes2TjMMr/cXB03WRYdGMNdnrDIaw72OODAjiY0n8aJ8sTKX08KGwGISde9Ud
9MU6AeIoPXYaK0LbbuuiM3QQBO6zROZfr0UaK31CYVQItrgfHjVfyObVrvLV52zavZVEHd0U1R8+
q1RkJGYZZb5Kez69Kbt/taspz1XoJzXW0wqMrzslF3APTlSHweHxaiA1v4ToXr22gond2Fe4loN0
e5vTnMrsfOm85ZTUnTQqCfIHploJ6fm39uC8B3jeRsV43KRAPKBDgEuprehbTVXJVoEtFLyGJKTe
ihoyfbOpM2DO+T9WIXUIwMKSPiZVZk4nAA4GCtb7iXeNAIyhvsJ9zHM6vSvlo/pwZ9H+3cORcpVj
qrEFuy18fE/KQVnXZqp7Zjne0f5DHZOtpKbceZIo3Q/GF3n2K1gDA2TibHUgDPFWlPVm8ie7ddsW
ysSCE4u1xFIJ5xOSfgXlfUBsFi6bOeFC51EpRWB6gLpo4e7VdE3JegFxx80YoTr8D+h/HiUIwalf
0HXF8edH2heXNShF/mVE7F26glY5Sr8W6hNpKaO+pC8q2h3JtO0WqZRqEzBQR1feIS5EiY7KTtPW
9ETJ+O2rRgwphq7WLouw+bnJPSls3QyV6HdB3XjF/0r0qhGQovRilsnev0pJOhUsbzACXqO32gC/
eEIu0UQhINJNl6wik5wlh8iXGwo5Nzv2/6GlDx3PXp2gft9Nyzw/o6c65RuN/O0d9efPE4N1+Sx9
0TLycgdNLMBz7PejbZdjdFbfWUucuCunAJNpCyEAIdWBXGh0jZOd30XYUMvenEi19izVm1lWUY0l
s8zXJkETBHJOM8j6Q3TxZmiPfoTaOjq1eW3ujsC5jbTG+S+4kdHr8SK0wWl5BaqGECD3/80utqXI
wKcitf7B2EWgPSiXsZmb20Z2FafOmM86rZHw8S7YgCMiJJIM5wOKfLhHjulJiSivqQmWrbrc5pGW
TDgysPzMolyutIR2RpiDr/XmkZ/3ip3uf4g0frvV0TAvwIzDDq93NbKBMql3OFdhc38sSa8hnuAa
+9FSHvU/HG+jJaQntRWkyQNytEqH8bcYgXNknNgCAfRHYlibCzWliEqaFJ+XW+GD4Z+v24P0tR1f
KR1Gpvd3kHpw7QLJBf2ys8GT9SfjXM0uQ/K+KLlZaN3P2fg47X9FoCxZxSjQ06cLSlOEsVvZbBOd
A7YZJ82Qne+nfp3rxQfEEmoFCiuy1WK5Waco/GRW6/4Y0SwEhuJq7Bkh7jqRv1dlOoLM1ky0ae8X
wllXofklCX3SEPs0qxihreCRHA8R6Uc5kc7FTrpjgM93+63olaLjHeHKrW0XoP6vOAJtuwMnl2fd
U5cQ7MdCLVvJBbXy128zNVanyDN74pBzYHECaFjGW1wIBJ53LB0K+M0XJwZzg3pHQXuMZg/TPVLD
9YBftnYOKswv0DLyeU5xzO78Ry5bBSEPo0P6fwgqxwbUwHpBrqdLoKvb1TLaGKzGHUAIXVnjKUnS
FtIH0egIAMltAvyFUpkAXFFrQj9U3QzZtXMRfkBiYnj51FjbRGeT+ar8Q/5qriGOXWvE2ZjDeHkW
Z2rdkXp+dP3Yr1qhhaWm7Aad6YmdcI9uYy0Y05+YunDuXuEUj1JVKNoE7UL0t7hfTgLESYxZZJJw
X655NDdQclppsC0lnBibSpB8vtIVaMuTCs51P7NfaZ7tegEHOXZgbiJkWnOkr4kG+DI4+ce5TVky
X4HslFPFYobnm6wtoOFXWSce6quQ4R9/Nogn9Xd3zHOinRv6Apu10l9XVYMBuhxVfpAVOXL06Oie
g++1uNSrTtlb8/1pfQadhjB/Yue++4QJrUqmK7tkS/Dk1if2uTp1Bsy2zXG+QTpKCHjbNJ9tjtym
aTutWjmI6yIoLpnRg2CBRxouMezra13A6A/mvMT6G11r8q3A/Fqwdld4Kpa0nd51raFt1sefnW5N
wsbfi4ew/YwnJYFAM9bvWLAHQD9TTiM8/kpSv6lkSpjuNoz9yJ8s66mastY47SM4IOsOMBmy7FQX
nUK6ivCngERJQtTZuh8Ts/BKCPr9nwWOK8iVoLdE6pfEJg3QEmQMXfCuG/hQR98sEss5yObgV/tK
VM5ZVsTVOoHltA0JEWprhGnHEfzXUD1UYviyjPG+QZBnmrS19TgceB7gVbbrITV2bh//MDk2pIm5
h+0TiVd3i7fTWf5lMItmHp2fM7L45VNpGQFt6YIMVo2rw0qDoX53h0FqXaMlO26HcmE9s4rpmDcO
jVvZkQU7FhqHGNJ5rgebzwCpmGvNnOqJa9W+S+/5bjPxypkrrO2XbcSvZVuBCw0N+mUVSfZ5GwiI
K8KXs0kie00qtk5iBxiVfIRjX3H7hIY/dElnSJFMeJlQMNg1ZZTX7ACG9hew4vjMB3yrIJGiJ6mB
9VOh3qv1fcF2pDPi9v6UMBf0bRMUz7ubHT9V7/jpBLbpNcFW5JxbRnB2mMoWQBVjfc5m3Lbmg6qx
SzSgNm1fCl7Cg6xBQyWTc/CKLS4ZLq+P5rLtlOkkgDuw6S4ol2gd0Usa5QPb7wcYVULmgB3FG9A/
QYPqR9og5R2aCdsRnK9b/RRp9j07UgFYGgjqNLW0iKfhVbaGtDn4KAtv0vrNuprwv4xUKn9ZjST3
suy/QBgx6x4tvcSkmCarLu1D7t6mWNBzzaFjHmhWzL2nYrA8xvI/VSnJI88wZ/i80rThq0Pti2aL
s0ILBdu8xBMZ3ru0Y+8k4PAIL0lOXX07LrGNr6karzLvibgT8OAPjsOYjEHkXPR5k3Tal1+CbDx8
1Ew1cwSDwxgQF3ClXY5LphON81ar6vRO6sQosZYmG6FnG9QCWx/lRpF/AR846osV0Iq/u+UHt8TV
LzWXvs/2bCa9VlZ5rcaNtNIf8bHDXiKlNC42FmY4Iu7ZXaK1KQjUlGAqe8cQF87AwPh5VMrT5ZxO
XujyDURozYpb0eSDmJfc6e3jCh+JkRAlG8Mxijc7ium7k03hj5q75XHQefNm+L+s4CCd3ji5Wzkq
LUXK74F5nY7HM3ReM5qzjNqacZojdWtSlyM50lZlJG+IuBLaIJbrN37ujhWOR1FB0/lYIJBjCDOG
GRt3rSwysLRhQ+/k/sSQnUh1e7Ro+uznHf2VTphFsZwaqYR5Uzz4eKl9ZE1Dgc0l2Gf0MrlKlhDy
uscatdwPrj2lL6rQFA2r6DSxf1kd9HoX6sWCRVgEmUwsMF1vB9nVnhskVE6o79Z5D7K5uWNgcmEF
wju8NAgoc36ZfvBSJ4A0ZXKwkisavwQNhXEssPY/o32z9KLBZGjEbDxqgF+QqZ+Dbwd67SdKW2zb
mJ7gfob9IraSubVX3KOPadCGPkfkr4FHr4L2mVt5ocu6LgQLV/o/0llTuHPkzbhdLr6GZk+9QfEr
64H7meNJa18mkJZOFHNDeBZz4PnfqzMhfouuBr+nwrpv/xPcW/g/DT6UTpfqwb3VIjhG2CiUqFyV
+NLYI2vP5TMvqW6HzroblExKtGFCXlZvTqMmFmDwBkBxPRWKe6Dbw13N+hdcwWu96gj2M2J94UjR
53+t0q7j1fAeH8V0NiqBKcBG/+ylG1l+5/NC2lCKxlY4I68rwXHI7UHLjmy/OWIvhzeiR7K1iEzk
1zoI+oY5Vu9sWt36hZHzelM78FHWslVl5xrUcUaquD2evT6rySJWIVzfs0FLCabuKRy5lHAFgq/b
qyceLYYfzazfCjKXSvEtsufFwk6fjh9Zr+G3NZ0RXOjw9T4zyKmCc5CduPBjCQVD48QntNwGPt0R
41tXfvF2ShYT6/7TyWBOtEjhDKxtH31+kHP95jlYxy1L5Ofg63fgAEwTvmZRl64Kmaj6u+7+Ut5H
+kJD5ompQmzSD/AHMGsht1RqahRLA/ntsJzSYSi5ZE5ErIAzHljkku2nhU6O6ac5KhyodYIhwIhu
WUQaJfdBvYotSmtvecN9beItmkn+aTwOiow9g8/X8bQXlBkyKUt02g+naxg39gbgV9V/oXcXImea
VtKEkaHnPEyuP/kNMA5kPRe+d1fFNt737GIzyflbREBI2waaVNFOGeonQtAs7kKyJjWNt5FT3WMi
IR50xq+YIuiCbB4vLhxAGB/tXcP4kLBw11vVwTkV8xTr4A/yjgy1qiiJQ7xI5CnQmruI4XBgFpYE
uVwabFJaokpumzHwoyO9pBzxRzqfI9/YNeWWs+wqA2erQm4qRyNQkcBhgWtYu0ygUVJg1sn5/DKO
4CV6uTtV0/MbIYmuwg98fZb/mpmsJjkO/HW1RtqO8TIPRukxXSVRuaKq4njcoewmU9Kj9Tl0DGrr
zaNWMwJ4qwvLyaUmA8C9XaRwV/Jtq5RlNqUKoG+Tppbab5uX9lbIQPirD2ErGE7I1ymRZtN0aDbN
hpCfynT1iGN1peKMicooy6Z7W0VHCEYxoaqPaWeFeU53ixzxHh+y5ZC/nnB8QHSpZ8xwCffnQuSi
4ZMw96GEWsvgzjOBx/uRq4VqnNBNThIknAE4xRdZebdwTvlWYXuVPo969O55Yf8DCE8uAxa6ZoSO
v9t08WXcI2WY1S3ZIU3rAFPlE+DWDb0aooBSYJEYfhA1clrEq2/fUOF4L+03zDpQZ8OKIXuGqz30
k6Wb62FBSfQc8TqFzKOlNBfiS7FjRL9kWX/03IyBQdN3X+r/1kHa4cUOjliedVy8JomT1dpgEehm
mLOCVGoauPAF6cAZcKJtmir4024NoLJZSM0nS10/s/55+RxnwOogb8QPEfwJyceVa5f5Kn/mQYHR
t4pS8Fg2GyHW6wGIwHGN33XBBnPHR4LpShT5lcGQ/lSo+9jhy3Y+4qC9DNjCCc9d6u+cxpNejWt/
5F6YAjkmZPMFZ3LJDqsKQE3NqZ9ebuX0PGGAEzlUwFg6KNHhkEIyeRaC6JWmb5N95DQnJwjktgj2
UfKY/ir1kP9p0jakwmeFq8U2QtR+g2hTIYuvClhklcoDyQqewLWJ7OwusF3Cnx76tZoODqs8jBlj
VB7O+t83ms7EzTAwEEHaJCM775YIeoo0c5wZpauTEjV75qlNkuqmvSPP34x9FGG5jd6HfWY2jE/x
MPMIN/AtLeFTtqNcYBkhRyullem44wD7+0OpxL+9OdRolKWTtE4rjSK9s16V19SYmZMsAplclMDB
MV7mDdCFweoNypnuGPwj/vBiR+nC5Py6Bp2HdoWv5QD6yL7EVAwjfD2AzFYHwWjmtPOyejfSlpfQ
ecZr5vOBNIB/OjR7tqXN9PNkMrKjO9Zwb8uWu7zsW5eNDuDL2egxqaYUShaqOH2Ty0JCrEf2zyJK
JN4+FeHSHiTXuPb/4VeheNEwGKTaF7GUwxLXonoBZy/LDnCWccpdIBql6mAoCOQJ3ZOmZpDJTqwz
m9G2guIuk9OQjLZrpGLTkMNPKnS6ArHqhafics6BrCvBCu1k3Y3N4SzCUbo00E9Sok+4wDqlMO3I
ZSSzVbc45WQ8atllLPV4CHsbkXxmfjFK3A7vMhchX0UfYrk7p5ZE9hbWJ+bTuRLtmmrx/Nnce7Jk
15nJBmFwXsviuynjFe8Z+ap+Z3+X95GAEw0rioL889VPz0Mbx7OM5YBIyUz7OLQXQQRI1cGjpKQU
tYNPS+MFobP3Osi45PmW0Ia8wCaiIGj9RCRzqBY1k8MX4uDm1Rp9KCS/8a5eEKX1a8FxdWIuWNvY
R8R5Ga/pwUrnyozgI4WL2pYMh2wSE+eTEI0N1lRVJuq/ejYISMnfgLKF1riUB7+lkGvu8ZOlOn8/
zZhOepu9grNk7WqMkHH9OBtoa02Lt3qonb37mF08YQTCFDQJ7S9XrwUvTbo4FOFnLwQ6IGM5Q3g+
AeG9WwVmC0BRlxt17URK7ct7LaTwaJ1P+KX1Mtx7JjtB+eETmBeT21y62qaWRJJWKfsbBR4Kef1t
TsT36yDJAM3rYHgKdKMg3nd1jwOq0JL97Rv1nNB9YAdi497zyxlZbn+FnL1x//tKOUN/pug0o6MW
h7aGlHku645BUUEZKecXnLCXBd6xlF0GOG8quaGMDDVWpKZ+ZBhTBk8Gntk2VmlpzZVj24D0GeOT
QYzWOQaNKVOj2XsXpMMbYHz2QSQluXVVx7RDCnzGHa54EiDejuG7nuoDU8eCZ1URzs2JT3YedSYh
x9vyROteCuHzR5JusIlqWRXm+6zhnLyWngBJHREhYOiwrJl7292VoUZmQYuPDJXqJk/p6zzRF9rI
6Orm/yxt3iQ4n6zm5v7/AjNq+ZFXTxxH+w7GQlPoYWn7iWh4iJsVFk4axpnGv785aimUZJwApZbp
5FUzy0NeCf1LBYRHDj9AqnfNqnoa6IM+NNYeDFkItXT36meZZzWDqKWk3etgXf7QzUqjxrheaMyZ
vC1dfGDVqLCKlY5EzgsuTQKJCC7ghrpZEIDKgup6VxmuTQyqgsJvFCi8N4jmLVzHPrXfta9tqvTf
y/OKOwdzXzTMxV8qblCBQM3zZkNi0A0QaunrYp1JHDzqbpfANgHebP7VJ4fSLCl1n+U6xQDcKfQt
O2wX+AF47nYIMNdsHrQW4jvb8k5S2maKyS/ZW6zcu9afQSCVp1wE3AbA9z0rtM7dqjBG1DReaaMC
kHez++Q5BfDav0zBQd94PEVTYTXJFxXRe5yfp5qWqcSS/LjwaX5oDyBDFSAWw85BMeh/3si//MmU
jcqwBcXm2CagmrEBOPNQTwvohtbXku0WZ4ph4qgTtnSwGO099EbTc+qMIG0bdNBdew62dGWKv2wx
SjLkI+mynE25CK39B+TK/k7J6MPMFPPtnNt4Y46GQk6e7dnyNHguEANcoQAFmUySZ2tIOC4rI9lP
lnFdiE1wTdWdfH9ZZKk/TuFlaz/0ynQMCF3GIAnXvkfCRRqqrXsJfI0maRGpqUowbgkUw9IKGI2q
pcUbx+4WKM8rmu7QNXMNk296o3YUNVEUJ5oI8H9aS8POCafWdJobXYx1qKKYmCxsRSqwzmv8uUo4
3QniU7M+oGXWm5opwPbQN23QXUrkvACduyyRfQdXwJC5AzN1hX9pfpOvqSTMnrIWnWcGvt9myREN
2yHFXVNrgWii6QbT8q4fK2hOEJn88yGqkvzGrU77hlIffKlldP/nvUeF3+Qb0EQfFMPQCHUm7Eye
vvJx9Wt8Nm4MdT/vIm0tdFBjD71u0KkcIMGB6XYFHV2hqknkKxsvmOp5UdMnmuRVOWb0ZKoVlPp5
eJCU5D48SpFmh1AXm8VcZ9DTu/D42Ic2TYpJ4MfcO3A9sxrN9MhqO8KeDqPkdpK3YQaw08HcY+Wn
CPULVtRxBgTFyop5P/2mFIi0t8krhInGdCmiJFo1def0SuxNrKxCLqOiUIkrnSjshcdWZHvFJ83a
PUcH3FgEa1E55PnLdhTd8n0oWc7gE+nSqi+z/RubByESyF5oL9di0lF05ruBg0jONb+fgExvz8eC
JT/dLwakHk4IkSOWLNe7Bi7XqD1VTG+igAXySbLoYgdvtDtqHC9XmpOyKrIy9h+PlgD2eYyAPmhn
BmOvl7Q00xZ0RYLxVA1Bp1+2IILxqLD8KJutj0liTDhiWtAcjn2Vn3d/jg3x7IeFFQdpyGJg/DjM
/GiMUrupiVIt+bSTG4HR7gbyEz68+CLmw7CKitmHf5Eh7IOKOx3SxcYqykzUTbRtMlMP7OHR5HyK
jiWeluiUi9bU4NqrqGp7gUcoPPU4w9n3gqSVbc4xfwRfjlykRP9u3+w6XJU1gHMTSUZY+K22xKVl
1PkViLcz5rjejUvSS3dVRsAXBVld0AOuAu6ps45tI/GwWAhskekOINCo0kbV5bN8yj/0zD/QfAvP
4zuSuhTkRXU8qdj1NaW+KW+Yzc1g2PL9wuaA4TFXJj5aoVqvpAKSrbMeIxDhVv+wEmkucOtFCavV
U+azWILiau8tjFJT4S+HYNbhuJ4G8jHjNRoj0qTI/GBIMnguoX+kl+JxtUPfDlylpVmevQJbYhj2
axJuON9ieXmffyd6ctSGv/uI0Ear+RakDJYru/47YtmBDa6OmMEacE0kbxQ+ZGHz6hrGgFt1quHW
Kg6uZbsCGfiPB2dJsr7LTP7Wh7J5+RPK/kGHCI6l9ZlTKr0ZkVMklMr0ERlnwCbKgnvhZ0xwKmGo
N97ibd8sXAy613Lz5ylM3HqQjoTWj7SokAEskSq3XP3c6xIgOoNXwo/7YbYzkxzHTXRNBwXGtO3x
Fvm+rjSHf4LcFc2jaGYP0FgrRZxeOVE9YlToQet8btpUu+Acww0JpIARHT6U6oyLq7MxEXujYOpQ
KL1s3dlquDO44DQWpxJTDXsUUyKwGO+QpjnxVLFJohqMGu0M/fXbruPdUgfE4vxthdWxGUAAa2O1
yKTk8q81ltZMN2svuDCwFU3G2ktbYGezxaJH//TCCa92bTDhNm0R0xb0h1tqcUWvlJI7KQ5KvHIE
3aXcxO/Ie3eU6TehVGmApqJwSJhLSOVfVsO86PkYwFp2K80hV/GpnqsyDVJpLm8m2aOHTY7ElRNP
lB61rrCWuCAasajXVCnar6jgwNGP6ZtUri3MoeAGJpwmnO18fA8V2FhRx83I88BIsLG2pG055TIC
y3MyNEgMjk+Izne/NLp+IqYvfutidVgsgnx9Ml6x6ov02Df5ZZTw2QxmwpHzbc3JgW35K66p1BUY
FkVpsNy/Lz6j1xfx9zjHMNBbLdC7laAtkpW6V9/Q2R7oqZ7SX/8uKB7oHtqHLghUxcU8z60AABG5
NLZHwj5dWkqAsiv3ZgThaTk5VdS6xMCJqyWmTs+GkAE2tq8NrfydBevhhgkrpHR6AdbMG97pXirW
dC0zuGbWfPopEw9388GAqNfb5J6r+u0uIOXapY7oLFsh6hIgnT5DVZbTuHxg9JQ8GEgWGuOxX5sm
OHqi2r25X0AQVDTuaoMc3xV4/TlSTp4Ezao77CdE0rAxIvnBQFYfUj0PZ3GL6J+gOa3TwUhPTmSv
Km4g2VpYWYw1sSBZE9YBtpbNCq3u7A53O7SgG00fWOUlkBzMImHpUiSi0yKVMhmz+EhJ41ayjs1p
LY8d4O93HTdvKYllVl0wLu7CsBJklDdb0LbNOXFyh96kTx5sz6C3we/Rs0TT6at9kZixF9cE4hPL
HOBYFm0FfrchJrjjUND6HtvKKt09Sz/2Wt3Atb5ed3nfgUsXzUgqG+Fr2eLtvW1Ml5NX6HDP4Yev
eYWBddIipD88icB37K/hUURN9UGvPeBLs0hTgAu32J2TJ7ZxNgyL0ou8WxCsHkVuCGtSfYEO28o0
5D8GyYACYNGwsCWnmLYWLY++TrZXFy76LHIqBg+nTXbrSdZEts0GxrJh4n5BAtNKqPFWqDAj+l50
Zk+afsC/XU390AkBVkI9zfIpHyXGpEtZADhQZ6/TDjDPc6D2XbQ1fJ8x4CNR4IF5qcuLyWJKcc72
jchJ+jAAWYwk9ZbxQYGiG+dbhDHnk2negCtvyunE5nC3ZkUdMF5Zbn7vSBPnP8axW0wWj39ncoCB
IeJybjy5ZlbRXhHMkcF/m76B6Z1lRLFe2GBIDoguewVzURTiaJURYtysXuKXFCjmQDDkxmOCiBBf
jA6ra+Ywd/0Tjhj3tSd66btfyk46Ar/yTb1F28dKMA3wgWguEejTzCm3F4q+JaejUVr3Wzh7cgbb
SP/0XiKufH2kko39sbjYXXWlngywup5mbK9f5z/zRCbJCVVu0p9wgMen9kXdvrSVD+cxXzP5Qcp+
Xd9HDzDrVQoCZ4jw9TGZ1j1Gnod78PPW6vk/oGO+dpBgVztb4/HMBYRQUgu/MfYowim7Pq+5QgsI
mnortlDr0PaXdE3bVNgi+WQRDG8Ve3usme3LvYQVAdVLh9QpO/u/biBWFUtKlnYoUhM4gIbuez7D
VhKAIjy+s2ioLHIwJfLHIqVKEmt2tIQss0fWtCLK4kZc7fcv6y+uI9SLjBAp9sFv9gna0/EQPe7f
u0bdXnic3vzfTe40wAxR7rhGE6UE+nDv97/muc7yBIq4O4Li9iD+WNCzt/MYpWyWYG+o0npas+Mp
SzChX4KgzagNWLnT0vKiL1r8B/XfY+hOd3IdtKUYiH+S4LM3qLeyHErTrCD1ICsKvglZqy8TLQhS
NNeVb/OznRACe/6Nl/WQKTEbw0IY2wbmN5zZluB1Qwdze+fwMezmCesQFaFUWwUYKemnmb9NU1hE
oxyGR9FtSa4YzOqmYktAh0HCB6pKi+kYSf+AkVgbWZM9xx+AdSUve9l1MFZ/c3kVcCvxiDDFXfKl
R2P1W1+RPcV4gci0csy/G/5oLAtwwel2JQDMvADpchOUmX5rAl/XUX/R1hxJ11CJlfYXBdMRI5Q2
0WLpocunUzGx6Jc57az8tfPfywsusp8x336YhFXv/XG0SP2rdHKtcMsMg+dojFHau69rIORqDK3x
8ja5P1lPt44yyR8bk+2pHoMh0pAc5EvSlYFVseidM6DwN4nUdPxSV+Mv8vayiLP6OBX0OIv5DnDk
gykRcLkYt1fQltoEq9bbMKqiPZxbpi1eZ7Z2c85mQJAtv+85nFrSnM54OYuX+8IFuQ5qIRXVC8ud
Llw47ysUzoGmmk+oHY83Q/J1/xYWod81YSVugz2u4wBUzReeHyBPkxsSKlKWaJ6uCfM4sPto6o1M
Ec8Y+25kCS9KXiiEOda4PwWtektPqRlQu/act40VL/0FI4N4Me5PC8ZSKVv5y/EQtgRv1ZKKbza3
H1HbA/pinJDrtOtSGXREzbV6K18mCtNpMDum0/78jToo0uEH+MFFFncFi1ElNlkIB/DnaZNBf0Cg
tMFVA8sNY4slOoTYTq0mUbuleD5TABl8b+nNaexazJ5Eu4dioygqjxnE6YEXuo/aAgaq0bYStV90
PEGhTp8v5Eqly3gh2wHgJNNLQE26ZFsA8tYWuLwuV/w7F5Ox4M2+mBqb0Fvpsy+mCI4TKInknJUf
ZHCo8ZRlbwpAUllMEDHaZUQEJGuVaYwuSEdLe5l5KsP/G/D32g4EAzYT1PDjOFSu7tglGzLyJ5F0
SU4Wc+e4cN77PnVbkHQcDSG/7FlQTyBumdEfGnMcwX/x49s/1bNYzOa/fGyU4WApuWbWZd9Xb2Fk
9XOFCj1TYWSPCUBC+M2q7/p5Y3EFbjTuLtoAOG1AJPkd0/AfS6/Hms76A3atc2oXpSN3bEWaucX2
O0QXzVdztm7BmuP3FLjrml3PAjVucP3lvInQ+aeXDzl9MpHyVSl7rvyV5PEw2+I0r4nu97ryhIa+
BRLliMXAIIeFJ24g4c4zWgYkQGX2wJlFeEShCULq4g9z5M2+QK8K6fil+QSHobUTaettfCRNb2ip
E3exiwA4Fv+mXtaC9FoNRjac0G0awq/+0lF5tmoJDVlKOsJ0/gSeqWUllA6w6WXSYxl+YaK6Ij3x
Oyd1+kjV5FVFEQvWrshj6Hi9EZa5p/70dNilNJ5ve9LhA1JA/dXhU6nhjt1B4jGw9L9L8YFcpcnF
7qs8Sc+sUHUBQf8W3nMndQN7ceAYlmtJ5kBFfA2Y0OukCpGzzwVX+ILu01Hwc7EWokxbEWzRbtEt
wJGB3MehG63KKddlWiLA+jFr4lOBkTLkdlq7C+fWHAgovY7Imxw5lvK550J1kgZeYguPNGSFF4Fk
VHzdyLStil7c9GGfM1Wii/JWN2AXVsvW3FSbkyOF+K4NGERj0YVHyvqljg6yDuJ0kmwjihxoxxKo
xllUUhbMd6zaZMVbbBKRNEdU2osJVxo1zhwOicUf4eab4X3oBF6G0sPtx0lT0emA6Mc5s3y/WjCF
4ROVFFL3bO1hK053V6/4xLPlMmwnIhxAKaYnJIkFQPz4MHD7/FMCFSGHtEwbtHDx/JHhpubwq2tS
pNH4BsBENZKNIBNCY7bU2GU74lmF4/7r14GuOYuC1g+SLtHPfX9jvfsacviwu/8HxR443ZN2PQmF
7vwHrl1JU4QpE0GuOncxnDUw4PCtmap9wGE/QijD07QTFyhWtdujOJL1XQIL8KNYV2AWZITIEUYr
hatVaJNWicZMJjB9CN7+8EGNg1OoFtaU+1B1LxvuRpW1pVp2KJvFAvaiQU+sOiXyjCQHK505mM7A
qE0LSb2amzVK+/Vxy1P3fJx/1uhB9w12Ke8gWSR9DAvPM8ub06rGKm/6gFe2SsuZQClWqMY94B7W
f8yRXxLXfidT/O8nILo3Cksu+wD713TGWdAaqJ9+eIWWvkdRYqWQg/ybOOz9HVpcoL82Et+vkzbL
yzotRcNQK33hXEIgoUqIKOL+nJ7yDRP9xBmixvtNatK35TePsEEH53MmW/WqRJZMm3LMSxi8Iz/r
hBNxXVHanJxnUDghgFJYsHpvu3xg+rmY/WnsilwJz2V9QqWtgFqPEA4vKx+YJ5Ks8lzUHXbcMy2U
fPbm4eJHpaEGM77rTdAGZJCxAOVl9Qv7fIaXe6+tiQ0suXK8zKTM/K6lbgPGLbKu1tIMYI6wmiEJ
n2bVrtDNXbpqruE/p08FCg8/qR886W1tXHQmfCvD0coNEU0H9CuIlQlj6XR7FLCmin5FLF3dXryn
tjl/BTyhKMTxhJh0bBMWt3BjhAy94nfTeJVF2Y73faILxl0aY4J60sgWP+zk6S3SghXsRCEZCtu5
YxF01ICEDn5fj0ZLnAKDbTHjBTEirj9CYHl9DiWL1TMS/FMAZIcS3YP74RzNxbbYx1f8AvhN3sZn
+x5ICfE7OVbmji0V1EGXpcU1jcQL2pfFqSUHifmSwkoe+k70mXA1KDf9ZIvqv9qNMG5/hs1j3n4W
2jzyYxywUcyjAJa14q6Lx1RjWAz5uSWMas7TZE6VJO1M48f4wLBuoo1zbT8aqLQY2wGl4C6Ru07+
nnV3TCuEFGxgr/ql/MmX5xUiGZhn+0kQMi8umZmgbrRvBonWHkGsQqou4nHzz0W2Jt1sR+/ubCZx
yJ5afu4P2O5S5BhwvDiIv7JnnulWKVA8SSBWu1hY2VsbyXk/bLvbWr+t3jeElVyadW8K4iNQJNK/
M0GPAI9j3rD7XTVzReolcPOhpXTmSzufV2KDIxi5i/xs7mYdVGBtJr8XMQCX79Q8y4AXp4j0hW6w
yj16osa+/Mxq2Ktu2igOqxsL7jC7vz4jmSUq6NWstSPrk1EwLbVg0ZavJ9koaMVI0qkOMlhHoUrn
ycei8kOL30QT8CiN7+04j2TqVOyYNTbUDDfmCvi0ww1BiINzvQi9zB3Hmo/aFy76s7xxr9esmSlv
uTMbvEGZdB8pryR0NPES39sGel+XkghSLpuB8ux+JJTsFwnSp7P0tJe4CDhR4QSbVaA6jFhGHGem
ilYg5nZaLR/vE9eZLjzLscXfoxNNcI+BXxiSb17OcRj6M1ZBFSbFMi/1mO8sKzr50lzHrI9NP1VM
m6NstrEd4E+NPu9dogiuYDHTPMJf+/zgGHoNdTidiAmvjd8U0WXEWSPNve2k7V64059rrDcWw+gJ
OXB/WqPEO52Tr2HpX3v8rKvO4o60qa3wzRjZ1h8G+zSnLO6ZF/Gez1lx8MozmjUCO5ynatx+X1PE
N4YplfswerH3L78ok5QJ4iSnCs2DFEfH0JyGLbACb6Ad8qXTKmfs5AzJwXtYroO6hzDHta9mWHOm
Y17gMmeBBhiO94J9mx5OCF68V9HrbQbrgkzMp8IWQ62WgN4F6Jwuw0U2MNrIz72aQm/xnoxLObrv
pe9CfoJ7mXVJWMq9obtJ//AHh0MJe4RySyhs8h9URp2Ji5n28aJaI4vU8Slu0EgdvzKgWola9xy5
4ZMNwXCOWeFSemNl6MZqspNTwCWZRcN7Na8P01VVUtj3jbz7P7mhWV5g8esxfaZICQHybEGuU4Q8
GfVavO4R2ozvycuZpiWINKSjNauSlKCcYieNyKpoOVOA2o7UXB+dSHdLnw/L9oxNIIIfOymwpX3i
7gR7QO8uBk32BF3f5Rakfz/zxz++7avozdDzw2ugT7K+pipkgu7TIME3pDPhtmASL+up8Rgo828Z
2aynLIhesBJIlg76nsTCSO6dnF68OfVOVZju735RpAKgM/QRZAxW4L0oUoA9scfK8HmMnzNq8dCV
We1nCFhZ7QDMRjxq8MhljoGt6Km0LCIEZk+RM2wty6vwK4lmSj55AAEh5wTOH+KLviSoQ2vT9RsM
BSFIT9UMS6tztO80grp/qLrG2jMJ3e4k7ZfHX2cp/THZ095vFEQ+9aO+Pgj/rBy7KqEvT+KVW6Yw
zcq0jqIRlupk10nfAVSovX2UevwQWWE/wqhouTxt2OeFb6Z/7BiJmCfpZ2ox7sdHynhh5xRpPAaH
YtfiIMYfDGIIpMcoQhfXzU6FFb7CuHWiOiQGFwYX9wwQWAD+6PtihWVMFgbEulUnnPnJRMk/bStQ
6uYJmnL2aDfEWeqZw0dT8r/yf6ICmK5nxzspWnl/eqFmOV2l9cM58pZUTZkqK2HKecjeRah46cHA
dDtq3spGnKs/yeBJzcc4h5UIKIR0IIA42TpKzXn0pBRkpaj79KsOuw6E1HJZPQZ801FTO3kDnh5f
8EZDcGLziBZ/2pjGJ37wTNQufKrvw0Czc1F7/iK0BEIgoYjWK06x+IGMS2hnFahXldUEitVTqzip
2LJDJHXfV6SzXpN8w04lkfPX9LqcvZwEbIwGFIMv5DYCUvZyqCX5/W3zEcytsR12HPChvem9We5i
pfPDupnEUrJlBbkKv47HmDH1crY/A1BgLvqsj4QVWVUcB03p08yRZzM0jGCs1D3tTrg0uTbMb+mK
Q6gSTJDW2CwJ45X1ZTxbq2pxvv6MN5ERkMRtZADud84iuVPyHW8/0/G4qUctpWUaQsaLBXACDO0b
Dj+xcp/KtX4+e7HFqEhgKqTTseQ52D3pp4bvepQ8k7j/sU0hSKSn4UGb5nFT8DxTIPOH+RVmDlAi
yE2RBnn+99RREJ0QBQ/IVw8EVUkzuOjD6eDFf57eLiGMKKwIKu+zU5gARfuibNstdXX6Qt/CkSca
HrLN39hnbsWSwSUIWsmJvQ/RKrCkpj+6qesr1iXM9yMIjKcee3ll3ABTQb/QeYN2O9fmEQOECJos
VEazVgC7WcLyxC2EskGr4KkXzvwu85VqDt0xchY+WtxoNDt7Dg1P9dRr7vLS2tMjzbBQ75qg8srY
eHcp74XmDpnvtO/QnLOxIXvkQV3HVfqazveJtrNSrb23hsKWWY7SajZgbQa2IKYCMbF8/2jKLjo5
xIlx8HWtxr8alGDKAX69++/nnDt5GSwyjgAXoZByrRgSRMdp7UhulanlAlW7lYKDdZAfqeLra/Oh
ETexIBiMWuKAuvZF910vRIZeeqIu777d67w/K7SGEIo+guf7ckwZGAxV2DmSF0XAODC5ze0bbmWs
Dz7kZQKy4RyyMb9g6L7oc3WR5q5wHFCfwV6yG7MqPuc0tdzE98/XD1geLiCzz3pVKR6ZstSFGxfE
nu9lxTUTQx8gASUxu3MAS5VsF5sD/vB5R/0/olZR16G7CrmgvHOXUufqlBf3BPbAmQ92fVvEYKxr
LZ8x6955ilLknoXvBJaatJj8kDHAGHvdTJS3G7pkOI/xBZNyzwfNKVy+EadTWaRb8qAkJtyo/Ecp
SsrhDzIK6cHYSVZHY/3nKz2n+IIKWOTyy5+iTK9Zk5FGF2j4ygnNuFK/eWmmf5BzGQBp5BNz4OLz
Pxg4sSyW58W5+sg/lLswAo+w4zpaw14SgVn/sotOYIemx0Xs4Zb9/ydJcxM6RwCHcv8zceN8bl2c
5QPRwxNb3a46yM9Ud9LgYjL8BBtaKi5XXqNpYm6aXMTbUjsoOmQAq9PKaSpljh+InkE9txGAtwJ6
MSrFamfSLHxKnOdnr/W/WXNcoE3nB5XirYGKN1PDDmuWDOxIBMqgmU9c3dKAiHgJefw9vNwyveav
loN7tqiAMv02CgHWF3Ha+u4pAg4q6xulXDN5hXgm5WW2cEl5drVKeh85P/2ITpRmRCxvzHf8Ix26
MkdhXGGyNoAfePRG6yZ4p68xkrkR1R8Hp3s1o16bMu+mXswTSYUczkVGBy8LUD9FRb22fw1XvGkg
1eJVovKykEhb/Rs2ssdhtbRJy4JyHAorn2Rq93WwCOh2DQGMBLgdUeEsJUsHDyvYfe6MSuwpaO3P
NU+KtJkNxp7x7ifqmVeMrBSfLpzANI8p30ej9Egi9TYbGpifeZ3Em4Kfthh+5TMrlfL54MIqEmgj
J+jZ8AYsuwpTTFy1wG3lbJZSyXZfnskNriXwPo9QCckGTccBPXoks6Rblh4ItWTGODbBAaNTgwhF
+rN+R7cTR6nWJJmCJ6uXF2Tr/aVcw0lEN9zuLzoYzrvca+j1FrVlLaCTQcs82EJQnnq/SXZtLlFx
bh66Q9dIi5WUWHvQFN5OtbXP4b26DSBnPlEf1es+7gkJzbFkAl3/v9x27bLNORfP6V+sNs+GUSe/
sO41CoravrZMGLovfMloNemaJJe/gRG9n3331/09dEh4eVc395/kP1Ef3jNX/8oZc2ZKjzhSOg1O
hMRTdiG9X621+0CO2qaqNLzacY9vWsn48MHQl4TPgLelt/q1gvQjXaZU9zonXq9pqJizPlQDklAz
I3cNU+yvsTj5jhE7E4IY9g3h+N12gd8mvzOzSDi2lQTFFkSJCESt6+mSgFHax8X9um4GPGg/heos
HVAFnI1uQ3DFBKRh6JZ3N5F9xXyYGgfJiQy7XmeZ2GV0uEaB1H6Y88Lw4ASdi8RAD7DUOgTRr0fQ
Ou8O7GUauXD+kDBP3w8wxXnUtisDHVMexRDYWCu8aBWqo5ZdwDibcd5P6p/mFSDqYYddbGQhqOBo
oGX/E/Hegr5XGgQYBUMQgqA78qlsBC5V6SCqpfZEIj5H5kSl1N68ZkMeYSuYKO+VXRpAIY3PE4bU
f5xvX/Vszx3f4Em4Gi4RfSDNQQUZhi7KLaYfzsTCK6ijzTMU+ao+yIXfsuq9MbnvknyuWN3nji6L
XmjjKy5RCaMJWCYBTijbj4j97ABJx6hUxLzsDBAygy+NIvzIsmp+ZdWGin8uuZaB4MD+aGQSN0f9
LakAEF8ADcdEm0z2iuacDroyCxjlgr1UL1Cmz4AJ6zMoRMaD0kfA0/qk7zry+GG1ztGRU429y+kz
kfifX6vU7oN1Vk/zIfgcPM7tYViBCWxUgO+S7Hqm2M0oglqYed8gUzE5ioPvMxfqqXupKBNb3w0M
kIzZ3weLjxVKGxSdrUZISRarGKV35DnhWI9EfkYDQd6BK/gJrjzAVARGlRa+8WMVElaFZjZnQNQt
HcJ6o8DVQzYKl73wfgRlo4+MKwHUKHmcnhgFNjrdEapv5Mf1vFpx8iLgB97YqUA6OBjZya1awsNz
EV+PvyxCzRv3nnlwRccj9VgmrZjKFT+yXBfbAG/7j3CtFSbfwPBYZ67UYuYMG1O2abxfAao93812
lyIYWjR/2/8yl3NhGbji6qpizucpPQg1hwPiJyNqlwNu8z2Gnj766ZH+Q3kGNLC6bOhZHjK/WWCd
q8iTyt4gRQ66BTpXSADDq/MWGcCMD2ZzSVrQCPzJb9B3eKKCIquePZ8bCO6hRGOixGStMdEL9FlF
G4FmQ3trP+22hZbS0ym4+yzzfgBl840+xjmMQmFL+KTlAJ5s+E8VWhnyq1n24AV+nj30wvwg2HUG
rtgF6l7OQehUkmp2KqOSbnpi2BtFIVBpXO+8EwycUDEBhZiS0A38BEPjU7Dh26k6MI/WSGjzgGkI
1Jf/pC6Z0m5uajCBxEVM5hhYhe7fZDxyZk0L/u89w3ezAQOLvgXUZW6hhas09795WO5czmRb1Hwe
TVfmhW3Fh0Ysmq2V8jwDejSSnd0TiTT/hyE5hhiUxCqVa2c8ouTDv7XZzaCSip+vKNtFM5AsUaWs
ShHuufvw5QAW91VV/CVKYX9ZY3zOhFsP/oT0OH7hL6fkDpnpVlkBmfUIibR3hzOFI1IpDp8b3QXS
TFByIRTMPZLdRH3KOq7GpzD/7UlxuDGS9f+10AbvUJssEi5DRquFlcHH7wbKj76uwTK4FDqLhJQn
jGbsTWCG1tRssQwcBw2ceIhHZp8gJ/9gYzRPCgii1BNwqFsaVj0C/AMiYRr3XbtwApa2BUCSWOKZ
bKPXiXsL7ovlag3KLI9t2j/v1lQbKPNP5gt7FYsa0rdU/Bw3ECEUui770eLWKnxf+NIrgox2V3BK
iqs+1uZKSFOEWBh86mUzT/PcGibCSOoNxXJ3p32/YcmMiVhxF6QkbGCiTDFX9lNcGq14khuf99k6
HVBpHwcqcszzJ9hkzWqK6XiT5zA2oO7GJZ5GHbnwJf7v1AY9gw+pN5nmw4GlmLxwa+l3xBBgxnmx
T+7N17ZwGXJfRCacLrfO7GHEwySdlqH5uS29NgyMp8aW7rOoq3jydEM9x6izO0p+LOMGP6YhOkfx
katErTUpRqmwBq0ObFoH2ae7EYYrvq85prsNgDRQUgscvpoTj9jLMoh5WbEZrLPnHb+4irt31rDj
+j/oNPD3qEcrsJY/HjryNypIda+dtNdq49LlUmWXHEWShkv0NyxCN0siVexg8k86mRCgMICL56sH
TY/9+5BIp1R1fsq4kHAzKyr1X7Q0guA0ZijtkLpk/2X7H4OvCtDYGO9Ov5FNHtKXda8/CVVTXs7K
Sp5I6/MWPIakOFdOZnfOsvHdqpzOtwIpc7bp7o94JxdemV2D8L3eLRGdbt7t1utx5FfbJ1hNZBXI
x/yX3Vt9/9TL2unT+qH4jh8SF2SFCEnCeZpBkrzXOm12XSCycEV4/Zf/upUNQgGSqH6a2EzUxb7E
NgTtGBzIc6pEJx0ekndoey5Iek8s9c09POJGpwzcZk8YDIYl8yd6VfCCepGpGZqbjpdtNiTv4G3/
E7+YsK3oRP0jVAzgPAc5FaE9UhIVGVgKfgC1zTEsuxOtNijpoh2cgQt0Zh1//4c5twfbqnrX21it
+HZdHp5fSTLo1SxY1b/HC5bWZt9R3/8dGiUVJJUiK1EtH/UL4ZHGwX367Kzvf5el6lAAu9za4yb0
4OEYp/PaCHuRFwcPX4yk7yUFrl/pxfujHHOc6SDMWnf+8JhWI4SvQk8WttKThBzn7TyGWNfZ9mvw
NIcOF+fuHIT3MWGr1snjhuG0hdqXXd3USMt0BDwemuF161skEi6fyHMBI8WFkwZX9Q/LWBEltv6n
+ATxqMDAhPcGss6B3EySIEc5an+GQhhUIa3TLrlpz1aBnTi+lvKAZvC+TsHOKaBEF/Z7wdOnqGT6
OpxxQ7f2h3v+Weq6P4/CWL6CEO06s+/Wr/YRpnH9KZwQU4WEdEWCy7E5Y7JU22OmspsjUy2l/J74
5AyVUVSs9ei3TCzXy4g6UDjIBeHMcc9pKx2COsXJ/jRs7BMGJaZKyD2j3fcIZxGVQwB4rS0I6ytq
wOVO7O/WHw8FdJljlaY6jTEzSNzYkKHlpqdtbRct1WwF/Gx7Qc8MIgBslSMyuBnFnf3Qs1ohEtbo
F/aDZm9WFE/zs/urjCdo9kreWJEC6kxpL+KobzBLnBHjmfTP1DtxE9taGe4sbOAf2+UVJULjqWjR
3X/LtzbqWRxOyg5UcbhH1oO54v2llDDGBK3m0atR50oVxZyY3t1BijWEdWsRT1l/y+HkkklTXaRX
nFB1OIqvvi8RVRCfgm8/Xf1J4SV+IH9rMlOSOwua8C7nXeCvTtZu/tpbu6MYKsoihuI/4EgvPgAb
EBLhvA8HmmcpTpiBGvV6Nn6A0fPkZUen8y7V3kBLM3MXQ6EVai0kQHepMDD29zUV87PQ+HP9dbDh
eomg7GBQNswA+uPlm0m8MncObLbG436UfD1BbyAND0JXNRNoFRZB4wIvfsHuPMml/Bw1CHsqGIyU
I9cC3pBnVpojnLe+EJnO7qoAOvn2CrfMBoGWVWApICxR4e3RC2a5vTIja6ARIzAdo5FX43HNB81Z
TgpamBlaPQLZEXgkViulJGGK8KJrpMEQBgAvLOXKmxBRyQqrK6oQtmgH7OfoSKVLwKUYWPfE3Olf
ZX317ELqjVO8T5Wicc3tjaJHV8JwCVEdPLOokHD3CHe4oBhXIBPG2MY1wKZpyQtZ78O7z1pEGaWS
4dWKSUJRtMXyn45zArVMDDlRUYjin6y/wblZfXQuPavd2sefATerAIduRxtZCnzeCmVD9nxak9Lb
D0rnXU5/Ej9k1UFXDqainmlVz6u1CSYmxrZm1zeUda4v1lWV+Q8U0yh+oRP5lQKWXklJGLhMOhyy
myEFFwDVdLHwSjqzNw6vm7Gfl5xDRj39c5sEGipbQWoqty3t0u9qq+gwkIovB62AICvdPFMxCpkW
oqqLReAlOMjMCwVXZWdP0J1IfoQoSfOilaOKaUax5lAGEG0oLo0hOKkFOfetiv3ct8jLtnabW1fe
QxnM8v9MJPw3dGLhnxhnyxvzyOvMkPamBUh4b5COxhXs+rSxPy/fefrbZQsd6uEViRJl2LgfzuZb
WYr73I33A/BEdeoki3xfgBIUnq1HelWmvAcBbeapCmArvI6n6AhIVAgrRudXduQI2kjf7eGBRkb5
xHmbF+Nw5v+YMXa/T8bRN6sk0h2tiWE+Q2XQy+TAp+1ibUCWTK+WY62MuAXMKBwZqo7KvJpluUZ8
+IpVANtBDOI8Bf6/XLuhtIQrXxP5vA31H9YK8t6W71fNII3y81PmhkBsgHHuqCNg3ywfvviofjvS
5895lsSa/sk/c/hZkPF1yL34FadlJDBop2J7+AgedNfwf/9/S7TUH2Zvm+7cy9pFm8l2UgYAkrdB
Q7klV1YIV0Jn1AUC3HWO+uR7PcvXS0URKwYLMxRrbgg+cDAC1GXJPYS013D92l45ri50wMAqe/r8
H4FRUyfExC7/sfp6ZmIAD29wZikz0zlxo/6QdfozDkS6e8liNizzAi//r7ikIXYCDBI/UAgYpv2m
8YlqkABwwXpDS+xbbaoZWy6MRXbcWJosekPvyurA0WsTHJqCTHy8kXp/hn7R2KaUaDTg1V+6PAdb
BI7D52cmlD0cZCDs/DkDzcE3fT5AWWIL96UrvwuBrG1zrJURFagC+Z1zejbofZNY4YluAfh/5SfD
GhjZwMAWvH8dFwJut4BHEu1cs2XkAIz/s6E1kpxfJP6qAH+Z5HtHHbIC6vTwMxygQQs6GaL4Ajj0
eEwQAgXxLFfP1MVeR6jJqcnrr83SQR10OafsneQzxjbRvHPfKy/nc1BtwZ0O/eeB+EjF7N2gtcGT
/Z/bLsa7zJGk9JjtrwXihXP7getg5k+BWKRaDeNbN9Dvi6EV8IaZsbM9W6FY046iCFCsU6jrKJbo
cEb3RQta/VjlyG/zZOhADbUPf0f32Wa984GdhQeTNsYNAx/A8EoftoPTS40jJl2dKOLCCtpjxuVZ
QP1h26Wfvo4g4fkmIkwCPDYy1TMYebzRuK1tlJ8wn5QdD9zXJc08z1PC/hrYpRVzzo8DCznXhBEV
IZkHu0m6Qcfsya+2OOA/b/7MKuqyh1fKSfEU++5X9uFGlRyvLU3brroXzogUv/C6zujgxONyO9Va
YN1vOphYixyg14pvnvea0xM/uuPEdNKCoYD1h2bFVWP25IvKgKn2IHPWZoHKx7pRQobKwss6q5FT
ZKiI+Uevc5iytEhzd414Rj/Al0co3ibB+SUQI+2Nv1Al+jfcliKZeoc4nQL0EtAThE1q/U08Gvgt
133f9NKmgHiwogxqaW0i6ab2Un4voYu2jgahshEwHeVpnEjEDrOGYRrno2w/1/x6dnoz/UpayuRi
7Ody+RHNT+Jro7o8wEK9wZZLqeMkPLbtGsDPfPAiBovdXYVfS7PfQl0gjq9gxLCgA1DAd1AmctRr
N51f72Yskx/Bov6zL3oeOzQkREgKeL+0NZI390Hva2820CfeMntd2jd/nzrFpDt0F3NE5FoiOLhN
IfSZKMK7y7Vi2J8jXtRQaar9/PINqgB4rsNpG5yE6cCFeA/cKK6IKO0RwppmzyuqgWJrwcNAIJfj
H8SJbUGdhWcp6SsrXzz4PiBZTm6e7nS+G9wWZMFF+lK7BNlF2arFKoRAP6o1rwGHGaF1x/BaLlOy
nGSDDwaB8fEfDA00oBGXTvaqC7wpP1XT+h8+Qoa/eeVWOqYKVmbTrlkmBSLu5A3jyp0BIenP/po1
tWncHzc2c47MJcJC7Due8qFnKwJiqu48f/pk/aVzNlPEUvlobaliPsWqcK3Is3Jzs33OdMiff4/A
DpIkTN3USJwXEF1xcTISFUnGwhtRxS+MNQxpjXrFrV6HeByhdDl8CUFhL3wUa/5oMG9vtHBldP+N
J+kD9aFRAW+Sqx9AbGlTZnwUaegs7mkCtdqVQU/yFcy33YZTAu0n8RVU3MkDZcbWVTjy25UjjTEn
roMCLAyBmxmBY1l8OTncmFFm1pYvb4ZGCIFRLFrUJ31D/HvriZE3rmfUnhz0OZFF1+6+6iT4bw9x
C5fOcrRsD/VzHzv7/jFxyscDQGGfb12Q8TKptZXeGawG1nEcJ0Twt98JDXQvORVdY+LdL7OoOACL
MHFT0bQBGIWgDVUBfw0nEGj54VwhejLbSCu/jcUb8Bvmtb2g+Rm87QAQWKDj4f0byRUh339I5v5Y
+inx1tUzwDLBA3CVfD1jkoTN6wjcwsVMjpiZSueodkosyjGTajZwkTPwDnKIjqaAtZIrshMD9+R6
Wq5L4SBcBSMibdq1e+nUXkN9elRsRJl1UeOiAJIeyqTIgPh5QErFe9280mYXtC6SF/+wyAQlz3vX
eDIVAF/MQp/jFgGHI7MUyKaH1t5JhFWUO7JmAHfdusGaYXhF2ksCCmLhbxKgLZVxBdKB/QvOLXjN
VLn1pB6QZauDevinxXijice6x5m4wDjC6ThgFKFFuV6O7jV0T9jlNr5+CKZRoctaWLkKe1sK0+SS
lHTjv0c9BrU0KpVdkcNecCo6pTEGQn/f3pKVtnqGvRwSlEsr0jmABsWrbENrmqWO8oFYwf/ps+6p
RPpQaoJmmnSiVA6uejhac1yYMMV/ORoiEdSIDbfa55Kgo71uP/u715jcTd8orrwlBV+rghZ7W+ER
xNVLArgeLxot1Ldkt2F6r0bYLzT8vAHai/eg7A/SwyQptd+O9yBnkI1hPRtV33W3fddgfqr3BbwY
AXCRQrt1y6gQtGKg/QD+fu+rIhSmmox2OCFQp8fAdNYIjulGMiqS/iLnLa+u+Uu0+ynhz2AYx3BV
PEDwKmIHH0lQYOJytiCKQReEmkMnA0hJFGLG+DYmlbNplam5FqrgqFiUTxVCD9z8ZV1FlDDbs4NQ
uk46nN47AuKyqnaUPIp6lJIjO2qVEmwLmhwN8ogNZmtrddf3jYYW47h+bHMIgUHYaMzlQuOK6Wtu
CE7EOh10svQ9nDSS1y1gAPzP31RxtOt1wfqw4sC8xcGfJNUWK/+pqLh+Raq0KndFOATogYyiZjjI
DdAaNGt3N0yRGAvCPdJwbBc6sCk5hKEWjk72BeluUoIz7cNAB+57tJG57fmsP9PYJIuXhTiKpSON
DokR8ikMOgdlOItL/qv4KRULFleYegJqVypwD9w5mmi3ITcFY3tEEBdonnlA72AP7byiRczSvz+b
jIAN6jrfBY7WDZNDTp00V4hVunfueGLq1mxtFDHzJxg66/W8h6ygI1QGuqNUrB0LeZb/uYjE2OEC
yj6rx2//1PTusJPdSvgXGsNRwAuaMYm/3k88VWJQ5PigyLK8LjO2lTbrxYfjsesGr5QH8T7ZWALO
ICeDg+X72NwoJtZhg3H2/puIlgd+T8/eltU2ce35ASeJjyx7XARCZ9l/I8dHaYqthBJsTRMgKnKF
2kDnNSe2YsibpkqeX21zCzDl4O9YLyx8D01MsxSq2tHYgOF7xjAuRMcngSGJxFA0EaDIZ+We98fq
vbCMeNp2cttMyHfM+hJpoBDxTTEufdHpoVRFIlGZY039KbT7bbhQ7/b5LLZMIp7BLQoO2VDUu673
ZJQl28XMBabG69oMjKFqNmICWDSNe54+XY1hpdP4U+1hT3ITP6Muf9O042vVbhJsVSpY+Y4zR/Ou
Qp0eSUh60c4PsbjAk3BwugmiM2IJXqkrfgEiYZbVzvzZqL1in/f/xwxFam1wFflYfSHFn6PFwZh2
MYXgrJAhGW5j/GjTlH7pmUpiIPhKlV9qZUqjtHJ0TuUvAByA5GJi+QX4N0v2iKt0e0gnzfO0DjBQ
2Tyg2ideLp3RFyCBxPLmviuaLM1koCjNyfHHOPuKkrnGIvEyzdiCFR/+3hz8S/kxGDI57TexWsh+
y86a6YE/rV/I0AfIJOzdRqA1OZZTfgn/neZQABuL7w9PvUF8sGexURGGnwjWRT/TQ/nuHU8cL5f1
BBdI15jDd2VoCvBFyeNm57cXqgCDC8NsTpzg3By8lqFOl7CiscRi0v3grGrhmNhUGeP80YMLmhLH
y1v2qO/Fux0Ag4jBj8tETLy7SdiraADANJ5BXTP5ofutsZ0MoLgEZ/Vca+Hp+MTAHudAR0hGgBCW
hIvU7MLSgmFwcpG54r1w9eNGnBPmSoKxFW3gJnJeP3ykyfHoavfEQ9beCY7wktioqsAurlUKYCDv
6vL4mZYJogN0fSplFILeFa9BQK+CUCoO2OmLXwntBZb/s2/06B8nBfCd2IJLXhv4B1uw1qiwR24S
Heg1wu+5+hddKzFCihNZ09iuUuoTZgnMNPj1zIajHDHdguGEAPqNYzMI3+8hqkHaR81OEtzq/JNB
kfriGJUmuW6ycqKWzJVRG5tV0BT88r8hKXOYiyid/7lkLkaT0Xj0ySsEIJ7gisGTCrcKSXAC7CvK
jV7554LfW1czvwY2sZELrzLqe6lexXlDBN7VkP3BkXjI6CSDL4xcbbPQYRy/O4B/iHvCp3kaUSzy
X1T5SKAZr7X3O4VcOmFTH3KqSNFdcUGWbZNDrOtkBhoht+8OzfrgOIa9RNufcddaE9H1EwxWQYsw
FWwDO3MMvompFeqvuG/ak2dJN+hVT5yrRs8D2OlZYgyxSVTnuett+CFWRpt1XV/HfjqQwtMjhqlq
iGfTOdw0lOJ+Pe6KnWTasIL3gg8nBqYRI9YCiicK5CE3kzdVq51Uorsa5mNFFo540oX315zraOnH
rJpVI0wFtahCMmk4UseFSeVkqZ9nPIcBj7TkGnhkn4TVUsMJ/rFnueFvsfohDZByNHYe/7+jJldQ
CQL4uKKd4xu40qZK04Zi5uOdeOn5sPK1dPgUSuxqoM6Gyzj16qiUsl0D0+o+XDWSE8dAVOHT5vSY
C21WB6XvMsPfZttp4/29AbxmSf6J/a2rllMvvvOw8RXp5mr7v6dNLhv83Hwk0ryy3kjVSk1H2oCH
IoL7ZXLLTqIXosK2x6jzSdkvxdYSGHuz862mLP47aUENoCfN/iAAFeEQNW/HfA0LUDd0/nCWDbSL
+wb97V+YYoJXL2MR8xEYhPls4FF5d6sLRIo2hqz7ycz1HnvdF3Xhzjx/5Fv96swDAItFblaZdmBv
4tyZT8UDAVmWIY20oL3ZlsNQornkNAJNLLewMpzX/DJSOb6HREH88SG5TpPfMq82q8lv80GOdvPK
c2VdREJWXK/lKBEfK3pSnhK6f+5lFCXyKDW4CtEeMYyjnjQFrPbUHGkBeV6n125BFQUgNio4B1Qz
lizRGGspaIi2SGAEt03CZaJGsKf3Pqs+uDGLX64CakPKfXnoj6riNXwlYooLM+tdoXYsGnrXMy3R
ML2IQiB+toxvk7kd3A4an7Rr9QO5EWZhoxe+E3Ji7itBDf+ROMEJyxs1qoZxKsf5iP6mEjzFK92A
xU5W2c/595kKlKzulAPnbn/uGK3M/dcVNP7gsdcEjKgLBrsV/sO7r34Ot1Bb9E4QvqULPWq3NkiC
0HSG5mNMpTIkFuRinQZVzKGRx8hIuKhcvrUXamhBzmL4kseinWQZus9UAPM9CbOfSTN0UviMhpQd
+LtLa8Rs7w9Y3Q4sHqsqA26wJhYIpzuMOPKEQxqpfEtdN8hlQoIQiprZQNtOMbrjicbzvM6mVF5j
1Rkployvqyl0N0Dvd0GfW9lIVN8EMZL5S9ORrsx4nQsEmR4o5nH7nXnYz2ss3Ou/xii9zw6HuJPZ
1pacKa2/O9veYjuaXHpjWJENpflmdg1VQAAxOYlqpYWV5D1r6qn7KaA5+Adkl19v5Ptqp4iCDte2
3sbTR/gN8XxmbXpObEnPY8wJ5eP9mnSXOTxhEgbfIHvZx48ht14qQiO1FhVNsiDkztc1s89Jk4en
ZSbluslDXEqGKwxwhu0kZpxiN+kKGilixUgfBym2rvqCkVuq/QxTb8jLNyNgkR8enZfHt6X2lMr8
R1Qjcqhzs0NSQkK8/dvGe/pGdKuRs2zvfzoQG1mIxeXj0qg5QCz4Rr2DUWz7ufsfNpD+PI5JGH95
Wli8OCppalDV55y0ZIUS7t38FRrtxGizk1M3M4Nh5ZSgbICkZBTn6qHRH0A9eFEYAtCI16MUNmwp
6ZgxnTBblrgmu+CesE0q/F9HW3/uDTWC3EDUDyCI4v5GNxMX727bsIVxPJQpmxkxaD6HjjTcipPO
iszL7x5oPiRR4pro+3f2BBuH3Z1X/3ZhIIpO0JuzCELD+98m2dWZV0KQSaNkAUeQlCseqNgXPkJE
17yuAuBguuG89FTiyXKi3fjMfM6RavEe3rNshAbOZR4CfBWm+zbQc3EsVMGSYQMBli9ijpnPrxAG
+b8IDPeXMrl8rNM7yhW2FD2Ur209kltA/U+Um9C2UmBHBciVBBRW9lifoeY5fuQQIFeuFkcM0XrW
go3YHGSdLKa7PWG0gyryoOz3O9fIYkfaWsKyJjco6mRfqR6gQqGxhIxLcoIL91I345qIk92qYyI/
NnpJAwrZk+AamF3/Av4mSFfzZgLxnvdkICthEorsMWMWrOrcyXKw0ZPaUXfNXcCwBjJH5+OwMuTH
hF/iBvFpyYqbs1jLJyHkNx5U8AmjePrDvFxyf5yYMsYGlgmPwfJaQmtt4bj/8zxot1XQaDpeG6yO
N9YqHuvTL5FHiTSOFbUcsMevbJEYhz2sBnLLhYeTs9jGATQdSInfahGEpWlOs9ZxpY97FsOG5yJ1
5/qvg5lzKrPH1L3RS9DNkUHjeV+ACW1KLKI7iKEZK06kDt8oHMkfSuu+hdiVidjSd9nugnGaBhqV
XLwEsibS6BQx3v7v0ZPvvrpaF9NXOFp/9P6kUHUnZyFBPki4DLnCLBLiVHQpmoIwGtefzxVJ9jOd
qRwDnnCStgQoWg/r6uJKJjb02iccaqLsz2xGySCPMHpYYzgc2vHvF2XuRV1ZeQAdvussZHkKKmtK
Y1J01Sd8osGB6ESDMLVJyYJE4FVQz0ky6ueC9mF+fxkxwXqJN6MHtckIhAFUmqgO0mb6nA8yhmEe
GGNmdlSjs+3e9NZ+k14MBOw1hqQQP85RHKnLbGzT0EHvKtSeYkA27g7kx/JCtQL5boi1P7Y0HK+r
6uUKqt/TcUwZ9ZpybXp7yfmn8IDEuhyzP1jeBOxCWEKobywhXFl8Yp7RIeWjNsTLpRZvzAnIp/Ko
iYzBP5eMQvq2yaHHu3pBFwfLiQOCuhuDBDZQY8dmhz/rf0IwjafEixKt20GX1hHw5WW0Qj9rmU15
SqM7ef398LijFtcxTElGscQpHj5TsZTt8Qb/NEcjsooq/5+HjKHTaBHEX6/QD/mUIjP14TGJBgAO
ovTddfAhki/adsmVYrMCFzyA/ojeVNkXmzo9AfSpRWIVD9o/vZ/hNj8qXPLKpl5K6oAfZKCRFoNG
ydNhhYaf771Qii7VWh9i1kSBH26wsZmJ3okncKwxyS2f831mmpGap8QfFk5HP4rrcZqPPZnmzjeC
bCDbxSygvxDZ1FbBLqLJJQXNyB0ybdu20jtNL5vHD0n50NftnvsxK7wWh6jv1WubHpApK1wDELIM
UCcBLEf1WGrGa9ovXvGP+r96yAEXZGbYUqiANXYOvWzxAyQ6Xljp7ix+29yJVf9C2VgGZJaVgSVW
nyRbCxMMZyDR9XAuMS6DcOXiX0kyRXBMEdMT7vqNHrGN6NIItI2Q30hmUrAYSpxZO7oPQ5lLxsLQ
8nAW6uK5GOVWHgpxBKwyGCcHblw/OJAT2TDqwu4Vxbk3xPkqz4tiQSDcH/xpRfKV0523vfDfi9WF
HsQYpo21zH5pHjyYe8I+zuCd5nehcxTLfrnH522B5/fUJPI24cLPsWuRzjOaXsjNHyAdNFKm1Ezw
2wHrhMRaaCOPctjvWdYnnoyCTFmoVSnS+PUVXok2nmxyiu3PwDcTcuVFTffsTxlnDYRzXCSZYa5D
rhUzTZGhYJIBgWq+5yMMeTvFsg3+ONYCwveJiQjd/Qxocc3o5LHR6iMDM7cojWWjB7nVQ1yoRy1w
plA+LN6LCXdS636REbkntujjikJhHNWgy43QHafnJnszwizE3P539bQt3clqeI5TXYD2AAFWgWeM
Ma9OhBCQaE7KGUeoHjuZUmsop8Y4h37nUpw+P79hNI2xbqDYScWcu/XQIJ8khxvSdxUSqlxL2QYO
0oujGLDTuTomy2LhIoKHGPQAT7PV3wx7K5HlhJBKkf6lReGnjDU5RMPK3e1+bPwfdnL2N+7glQTi
0mMksuXndoYNGK7FBEAdr1xMgmAPg+K1XR8YWEMAWAc69crCcdnP+gU8pWegWRwlHJwSLiIljBzp
JNJvSvkhOTagxobnxCNJ2X/kEtwBqIHXDxBLQ1Cb0yROpnIxxt7c5JN6ih86MnQMqqNF173NrccP
seLQCC9mqlHeZm8HQT2sY2r/GlrXWlvn0j/TAdxZLHJxGQ351oCZ3OfDRfSS/25glotPxsGUfPuG
brlmMkJKbvMmeV/oIK1IEtAiVNiKIedVLhKw4GdA8IWeBLj2Dvz8rlp3apA+UbS4t2GYZAyNhMVe
02wEJKukW1OHNOREhTIrpblX5WRcFKKhrMbmnVRWZ2MI4+o7Bj+Zxx6v4X85GUFV3y/AVMQLB7yh
YxWoWKCFrutX+u01wC7/T6TLfwU+W134HPJS5vb/rncGVb5jO6SY7qDZcMQZPSxVWxPskFCQwFyJ
xfKn9kiB7ZHgAPiYifyxFkrUKkCjEZM9Y1J3AXiHB0CQVbknflcTTXtod/PNBPudA0Z2YZ9jFmqW
gosSPq5wJrZbmTEN7z688raSldJ0a0krA/bL111s4TjnkI7OQPCvWz7IdIV6BlMDc2F93orf9RZL
a46VRuDcODeBFvMH71YhaVm/Rq48YuUQR7ZJ1F37Z+9UvSk6mpNKcqY2wkGv2BAhZM10BAjkG2ix
4BOCHKbIrq/spFUYNJQN4bExrOa6AGPuLvPnlT4K7kx1k1YPwSPXMhe7bVFf3uCTMKM81ic6S2nV
t2wf4QBYfKg5uy9S+p5qGovEmjPddnm3ny8F4LCom6cKlUgW0CZK+C4OqA4HzhmPa8YoK75zjwoH
xIXg1UTjHLgyYoEBdE1fiQvVUVFG/poyeWYBkqXBiDncmpW+AeRf8C565CzOmTKBqw69F/ClnNzM
VVcyWDMWfNxoq3FTiI9Gt3O2v37vHVrUpuG6E+0lOtVN/EB0tNChBwAD1qiHc0lg8hSRJXwFbc3z
wNLnXAu1XfVk6DqJx6wuy2Pu+52W/Dy421W+4ZsvQs3DVMh0QcISDYSh/wHVDUwCJ10ZwUoTuWhl
t733pa0jq2f/ev88Vt3wgiifi4TS3vPVvfg9M1ZiRqopThW9U+pIX3u0U2r2UGdcnAyZqhyi2/hW
khiOpIHppu5i4RLDpHjbBc8VqKr0TvcsdwYBTmNFqPUcZ4ZsFtb1LaGiHaLr/UeCSaY7E1t340NE
7oJylVHLsvPp6P/PkA/iaEokaQLJgJpQiXTuE1YLBBox6U0CGcMLv8PI+WXSG0RZNfhrEjJOlj9s
OFUs7wSdQURyEYQeR+9KdwXYeMTsxM/hqM1x+N1ce7vXdqvXsfSuEeFVxed0uO4muGbCIvNHQhfC
zcKVCSgnBb8NMWO+bb1cbVgXnP6XYZoPBnFRahrJTKn+bTesr/7LlbEKnnMzCI71qXS9OBe8IaNd
CF345Huh3k0arHdOyrCi3qeMPsN7mOj7g/MlCNVVSMj+OzRJo/ofFeGivAaKFimd6aXQ8DWC97Bz
yN1G4NUB2/doVBXQeiLKzrLZHzWx1yWHNsOE8fEXEqNucM6mw6sxRvnTUUOGaUPGg6Hp+3o6a+oX
/Ppm9bAuBpMzF/ZuahE6U/JpdN4b3Bnx9R/O/uBn+oSTEzRLkHxKhA41ykUspFVipfhuGMjuk/QG
MQzjWmCkWEHH1ffXVNhnEzGLeIMRldLYrRrsRLAK31rCOwwYUePoU4YB3JJPpFDpwFgRwJRquQVR
GqMOFu7PH8L12tWW/XSJETQVGemfYNmlHy7gdYOuWPcQG6Il92uZ3R6IZDatosQiCEXpYykhttzU
0oGLoWsLp3XDbtq2PkwlLTTy2XkIf1OvfWKfRwI318ExHR1/QN9l7xs7BUjKmPhL0pAnhuqEAjxR
AV0R8LgNfeuDqHdtQMfG3dPJTtD32E3s3hgxGfWna/h6+TQKeH/PTdaXVc8+xBYhEqKGcE6Dxm85
r3GTjKIl/5vIKOqOzlXG7geRyFK0YYv4fiOBs+ELucRWq9R4SmfS7RIWDU5JUJjsGtaPLoZmRJBg
sjXg42dYMmIhdr2w29AHzA1e4tn5kbTj5vQexWaG08Wns7mzex4+yj2NXklO6G7lZt9RCyfsoVBS
2Dr2cB1YA/zrIPyPQVTYYrcWGLc2Dr+ziDVP5S0P/G3CwJ0WIZ4QP0Ps1BAHy6ReD9fr/HpPuWOT
TX+OrIk+6xZLn/BTSVV0Ku2yuiUx2EPpM0xhMjs21KTndmp9E9ilMrNP67FXpBjym3AqjZ50aFNR
ahenxSX/y9ovkYGSZI28bwogHcUQMWBo7Vu7eqIlgv3hTjPHU++8tVnqEXOu3xZ2NkAEQXwCMeGD
guz9+gcWwFcoo+jVy2miv2GM4WxSD/U64GmE7mAoUoZZs6iZrustK7MG8MZW6WnLKd9o5H3achnV
L89aJA9vB8+mRos63/w6Og55J2OSLVERJ3Nfd1O4bS0PQvsi/Ng6qFNFk5mzAWgQONkLzxHpjLG8
LQqJknyy0KWgsO/LFW2pH9LCR7Comzs49/ObngbH9CDoF3UFeLs+PxNd+cFGrLnDt0VM2Yij/AR9
HCtBKZwEi+66X2ZvqTM/EOP1IpVAdNlX3ubfvz+Tv9/4cAaZOU6Uh7kjrzNOFYZs7aV4JclYXq4n
zhZYWXwTYam7xzFi0T0ianv+KlsLtkGG9pW+ksDhAaHRuEdhXEN/MBmuw104FiQ19UaLu9KdX59e
k5WJIy6wOVkrPDoWR0efDDGmDMkgeevIgQi/MnZiwEJsqH8oX10y1YT9Ueb0w8d+A1jsW0H9Ha4a
E/XJ072lkkGlGWUc5YTDxYlHmovWKSFjw8FYigHmY59tu0ZCARdv6G/rG90JFtvOKFunp5fDuue+
uohPuyJpSuGBLCnBmG5banv51fVn5hBL/yyjVR7roba/8rBTV5nqjONhrF/Fo6gxGUQZe2IcdHVy
nt39Qq7iwWSTSy7I+cEqOXlal9S46EsQgnHUHY3AIICGfIHpbWSAddxAkNbDNTS1PfXlekxaERc8
AfthrWJAHFYicQ0AHjau4i/KfUXm4/pXy0PMbPI71AuPAopqOJQYs55Hero2tNFYz5KR6xfJ0IJ8
Fp+J7gnjIuYEOkPHDc0okfpA+aDGNmt8P90Kn6WaN4NSlVF4/I0lgKEKZk/mr+UfZIcU+84bj34O
fOkBIp2VTHAQkDeGeJlb398lxQ7bXhSgCmaTIvvM+Omf4KEGu6keyMqdOdLM80zSLEt1QgiQrwOT
IFwvvPzCFp3V1K3m8kPAO0lK8NdoSk05T094PQzbuoZKNoXy+h6DL2u5LMmpz1lzH/MCKxi/MrED
k6NeVdudSLHVDT/4I54V5crxm4eGpvsRsECw0WME7bhXNC7zkbS30Bq/cQVUN5pb5Qi0ufoxmMKM
SS9BnbNKOlK6oicFpK4BIDYdCqm8lz9aDV3gzOu9CHh30wO+BjzxqEKnZK5FugPcVPX/xXSjDL2I
4vn9MnaK1WaUEBz8hPOQA/7LSTkdvsR6JzU+zUZwua8tONxUmYIRHsyRxHTEnayQGka32f/LpNEL
EMdX1qNYacrQq1eIVfEXiTZTWxBJlkrmsdUJHbNBrqdaKWuKBPtFiGpc/sTjiyn5UaZJogPivi+L
eVMQC8ivdqUPqib2TqwCLFmVOoIYFAV1I2PjBW6HQf0KRe4HDDJsK8CHbH+hh5DlBugJKn/xZqwX
PevSCWslBKtoR9HMxpKwLOH+KukFQp+m86wm/5LX65BnkLeYE+95Ql+VuyH241YtLDhfuQ2Jn2fW
cQ5aGaR+H4nnD59SxfVwRiLzYFGjB0zZ5ZWuABWhykvMx87oSxANf4Hrbq4MT785I85OvtvNHwbI
kabirBPrPW/rg5R/AoRt8Lvpc+87ih4Pcs0vKLk9D5/ljfRJpLuUBtQzFzktDMc0s4KnhCgSjS40
FgWVdnR0eTGsxh/sqJfLefMORQV1s0z30f6TGSjAh4kgC2HTNqq7mIwadjVZI2zdDaXVjolfmrE4
IWNDi9oB9KGH9GZC3P0EVzCX1HNUhrGm3rF+9g3py+IIN5Jqdr6swRL/QV0lmBgUOkfYCfGkdUIs
8vbU0zRQ1ZUolIhp0iVajrbDoto1+9fxLUGGNmC7/wEP6FT8LSWf+yaoBTqktSPGDtaC/ZxZr4JY
PUMBKHJxfH410AAu84SgQvnNNpklh6kNu6TAgdN+FWTP3LbJcKAZ4GjkLRYdXPdvwjlmU+qxkL5Y
x1N0/r7lVj7ebpnsL/9iZ/y2sPgcIbtED4s5PUso5iUEym86Rrl32V/GuKVXrRMBu3ingHEXBnqx
z11xg4/ybDd1c/Qrcy98xu5DBwomJS19c38mctdeX1p6DK3biVsUshNioTRReyVxcGsiNFBpCBNe
Vc5NIfY3u29g/fCS1oMPTBirzeYsurcYzd3993hS78Xn9DibwaSe3/oLGpL2wLt7s3ye116krzXm
v5mMlrgXnLd1hsgfvZpXvLvETL5KXnWO9hItRV6jCcPnsSeeljSxgqG0CfxDBzyBYGFVxTB/oF0l
YceTcIZ/kvBdBhqzK23OccI34B9HhiZqMLXN8l6q/ZyjUQ9oaWCZtpiuq2qp3E4wAc4SeaCnWRMA
P4yz3zf1pah0lZcF5pHyU65xUmUG0LUWMv66S7V52YDX6aHuG6AgEF9qzflcWTpb1dhM/2EwdjxP
dOTwI0OiIdgLJek/p8DFi5blaeG1XwFcVtfeFLl2lQpaj22JdBJTxDgMICykhTLbKK8nZPWX6LxM
pkJWDIKQVNTUnocv59AYxuCoXPY6itUqopgnuVgJ9kxgUx+fvWxsIO5K2CAc1+5LQkoi3s4KwHG3
oAqNAAfEQutC7X9Jvz9JWKpukG0SCNFFrYJHGoPsAez9P+J26pyvKW98oLiQqEbZABWwtxOxn8ak
EjeoSesbzG88k5mTTVTL42xZNfvN0bip6XGCYOwzM0zkpJbmyh1U/EPzI+18j31Xj7xdmA2zb6Zz
cM5iVSwNoXenBdLtqQQuwpHo95y6MOoSwyhT3nuxuvLXF7Pk2WfuQmR6saXhfuZAAO5UA8HMTnra
BRlSgmXUfnwismhyvs6XR/5zUHw9VEWjVyBiYJdyuBfk58twMw/3HqfxHYJJjpQY1YRDk3xikGJ3
y2Q20VY9LInF+O0Ob6tEM6TKxoNG1WUgfVa3tXnFYgenmR+R8Dhkv1B0hPozVkTGSGGy76urbD7W
m5u6W1GrzjmDAOF53phr4XZWpwa98vP2HtyF4GiwN8gSdEb1M8aPVMRbovpDp1uySpDxDSw9Qi6B
Tufby/ggVtTDwH8OEMVMoQZjjYst8TqyncqZyyGkRFn6o4RjNyWWXxbsFhAUyNfV1x8y7xe5qtQN
ss5ZC0/gPAPzBZoir4mKB1xEHPcNK9nXpVQ+qEoqTJ1D9O2sIleGJSLVZcb9cLWq3/JoSqEmJv0y
3XzhS6nRb/S7BlnVmhrUpbPbetqQYLI2h/wk50vy/bBsGMRkOXMymQ+bF1d/yulpG997ekQ6kpOf
beLlQPfdz93WH82HrX1mWUBJOqW18jX4mUMZeoMd1Z6MBxzuLRCYSKAUw+sXgU/CiRL2Of0Klioz
p1O1Z2mTBT5U7uEexNjUjJe2hTcVHLNR4z4HAHbvz9hdqNP1pQ6VniuBhbXiYxbtOJkmee8jGXDs
PNPoOyIr8Yf3oyj4Y9HMTtBSNAwby8VZdbOzbf6RwVjyhNcQftZDjQnHlboFnInbQc6c6Hua32Ka
3pPQeX7PnzNGM1YmBW234zqWApKhVrn7DW3F8lQyKtmoD35e0Ov/aDW8n2KX10tBZnhHDNfSwtyr
Lw/uAeDYXJqL7XiyooOd7aZ57Vh+RFyAA8AFkygs0XhJnA7fi0Z/KquTW5gT02b38qyD9z/J87Ah
PzwH4a+jFyxPiOm+VNB2+uuhojnKuNL0CU9dshq7BFBBefsrJtkP3PnFfWcSxD7J1WgeyT8Dieex
zyOtGNCrU3orlPACr40I9cVP6pJtIWujq5RQSQ3PhC2OdJHiSCPS/tGimRWM0LOSS4XZjhfAuC53
d+nB3BHTviYojN+mvUOHOrbE3g8dnSXuXg6s6tkXXDQN2KhBcn+zQcM0z4Vc9wTTwBQUwesCUSAR
MIQz0fwh4f8lChaMOYNS91J2/ghIdk7R+l/vG1MvkMdqsKbbIRV31jubgOA9PwyvXOQ3qLgvrw+w
wkWPJpQmhXABTdomnxxvM1JtWZ8cfdnvIHuHZr5lry1UXM+6yygWaTT06H6CS04mS7K7oHIRg7I5
s+C4W2S8tHiAJt2+QxfVWVdQHwrtWVRbR53k2MRWEIbNY9crwqoKvQ3NmQTzJ2AltaOLDlUlJD6+
P+sP7UIfen2yxmiulYEoDP6suWK626e6NBPU4eWci7eFBidl13JCmq4/H7WUY2m/2PR/b9nELodg
RCuZHmqO0cTSOHPy0jS2rcf7jEJCfEbE86F0s5082gveDhCLVIH5mRizV1PlB39PH18kiTve/VB4
fnj5+awgxPmRB50/7WfBtbq3/0hcMdsgOKSvXvek+qAVXMR/RRmrRQpTecfj7eEn46yUK/X815my
KpXzOXSedI/UxAMt8PanZBtnSe++/ApLxZj9ViNrfbLKzxB64xhkGkexvmg9Jk0h9kjnCZm+Mqyo
D49xnp5wpLLamdf1AXXshlr6F4L0k8Q5oxJ4tbRtH0KnGHDKVWLdVNwhZydgINoZhl79Tdj4K2RN
vdXTgobDF/kxB1rl7pIUA1VODmboEg5v+hiVc/FrlgyOBHxC09RN8SevezAd2Id3G+ghg4QfeXd9
5uynsQpjwMRA5Q47wFdbvOytvdeU0cWQIcFGQMsvA6q/l64cn0TbS5We1bN9MwQ/4U4iBlZICNYd
XEh5CuAfFif0cKRppqMK1UUV7aDk/ltPscoSw4ThlDjYq1h82p+m9NKmsMRP/bkC8mEXRM9N2TGD
s9n+D6XUH7MoBJ2cpGtOj+zubOm3UegP0p33f8uPLkXYBO46sOChxLpg+9L4G5dedP5ZGuLJSD0H
RAIPwaWu581EG3asQWvUZIgkhhG6AKUNePkixoIwYMjeRylBOOvy4QENZyL4NyHXD+5ttQ9Fqn2i
Yv9nPlDzFv50oMC2j8dz+LEPrAUDr+6OOKtrnaUtrXZEMnSfI8/MTiHoll0b4UwHhdGwzUN9KxZF
9Z+GRwM5TBN5fse9ErMboH8hFfCqogmIJ5PanTeTKhW5WbLkrj5Twdrg4OTma494WW68vcCpUvHL
Bks33Vu4fL3d5prjutQ2JbREchmoygkdFxNO9jDJbymDRU30ClB6uXNsLp5dRwOUVP0+aLxraxZQ
yw7CNQboffZEAngS6qzcQg3DdESrnROS+0gEVRpClB4e0o9sjoq7uEf9pFdhgrAbbo1h/O8Y6KXk
C6pLKQxo0/SKOK4up5u/bOwWf7TN3f42rm99k/ca6K7F22SNlwDCiCQtQh2fPi03IUf2BLxQrEFt
jlFXkd6mk34kDDanautpIlB5YzvFByHQ75QDCjcBdsm2xT50Pg0XPXXlSQcrsfnLPe9cmJvNb0Pq
FZyNUNwix+3ezeEYP8GqJdmurW+NHEQNRBzOGt7nndGPdGQBweDH42wPaQ9I4vKBe4lkCwnrlnZh
p9YJQFvsnMggQ/Kjxq5LW0mCfn0ScgXM3fCSdIDjhtjWiQjqijmmZ1PMPrycQC2pnL/z2A8suCSM
MxTPU2WigacZZDn6upWtKUE0N9Db8jclZo44EkqnHc0pNzilbc9s5ZqUm60SVZpv97ksojanC53r
96NB6zZkbsD0VwdIKtaOPeYBCPJZe/9Vb1FQs9lelDtxZqDmJM5VqTsd0RgrX7EUcaElBKcqRbjY
VYqelidBqa0JSGS3GB62U/ttCj5AK2ttORBUJzUY9s24ytV4nueNxIpiRW+0EZbvnP8bF7pelGL3
gduRSE/Uk16EDpL4AtMpkLnuUFZN8NI9U0tQuYaoDxanrsDc1LraN8s3YI3RoZQFS5XKmzOTpsKU
PID0jOG6DV54o0FeulzBHrqhhdZVrt/EqwZw6/nhqz4G/TiQB+N3xn6qOjPfWY2M5DbSXErJhtf8
rkjEgRvdqdEZhzU7Lh5VGsVM8XVe0SYC8/oeyV+Uoeve2pjOCXBSo28NBV09gymG2I/eZ99FDQRD
+NLUVwPR+E65o3B4uLvguE7+l4Nlf7SsXJFdn+JiKW3DYKOFC/+is5Ao8qxjc06GCDF4/dBx2mBC
IvP2KPoxuYqnExciruFKxbcwf+EFX3+O9gAL6P1MvL8L/XT3tt+8fBQxNIl6Xm/XXkUznUWLitjb
9/OV+n+Auy/ZtR3eoMwXXCjk106hLRTIjh7Ja9xe7sjM6+qWB3yucw2irT27CEJiejlM/A5dnntw
fKW8oHcwmLMhdSYBqNHhNOdE7UBLETLvF5y9kQjKChsU9pyswh/koYTNkyse6iOwLWtzxF5A6p3A
/J/lRO2sjkB4vyyBs44kUCJid3i6fwPipjq54+lQm00hKtTdCAoK712jYj45pqT5qFmRvSdtXKjd
1e3S2uaODlu7vFy/pJ1bpUEW0ab2D/gV4YgpZHLGWvUvdog8A4aVhz0cTQHXRHcU8HCaSF75Votn
rdbAREkr4vyvzofz4FttkV1cCIahRrL8lCS2eRD2BeTWKP+LeydKGJ0oqU00YHRk2efJxYya8utS
Vbey+j49Hlvgk4ke8lvkwlepi9cuKXOr6YnRyQOQ4aFGtuKCmcIaqJmS9DI7BRCjx+6REuDHobAu
rlkIzESIlWgWXuQ0igj4wREApKJSOQKAAD7/q6RV+jxGikFWGNCVgqIyntiK3Cd+sWq83uvmKoN2
okdUqJXli4anmNqcexDWxoFavWBuaqUTicnjKN/9nqQsVxVnPS0yQNTKkio0YdtzGfHAQJJu877F
NjnlOLZhAXH09pDRxPgZzrWR1aIZ1s5HEAgJAQbzcxtOidsUbI+msh+CYJf2bBfp1ud/84EhNyi9
/GHtwPx9l89sbIWJIZwgEZcxvFx01vv6Tz/6mxAi5mBkVGHcZB9zQIjh+eSM3rIBNlSvWafpCE4/
9bzTUkoAaQjzVWvuUPb4+2TS/jhjyV+PVWKgOYKe/eSkCgeEiIFmJ0xQY5Xg9HYjuEefLAbAM8Xb
CJlsXY7u8BDioJeDnChQlUJCVd9Yoi6S82RtOeHHtETaeMqARUq9REcI3NAlys/LBfSwErXll8i6
dP1PscbgQDJ59/CnoxlO74AGrwuyfTlkdQT1QJBsqU46cdPysUEwffymKxlUuMQBmKkl1/0GHvTm
ZgTeVJTU1x3XNJpMJZAFtOfR+htOX/72iLBz5kQRyG9Mg5VmMWLAQsDIdXeaBWVbjTukcZLYW2PF
c4Z2EpViB1hzRfuayLqbOthiEQnK/HdFHpZNoVQZLCWw5XyJuIYTqxGjPs0JR9J2KwKzgS+XZGw+
Oa1giVcMHDO3I1Y+aa/3P58A4kdlYyDUGdLhC7V5aoQd8DC//rcMBs72rU08olzdSavqWzjcrSqG
hQgh9z/qj0Oligl1Kgr6lT5vAj3VlD/nNA328Iwt2IL5tPWmIyRJMCZQbH6Xolswl7XKkLb2DwAE
WcxKxpbM7lPsQtK+pxHRtca46nhAvk1EPKgTQXLsMijlgylKUQq+SEkwWD1pgN+Q5W1MiLuUfX7y
1x3YHoSDdFSJ9In5/ppvNSAMhAL8LnYKhdWYMg4FMpeWdlBxbOyL4GK9sFgt0H7jyf+HjlSK12Zi
iiSw5ueyjeYMthdxJqgurdjATbbMtnq6riU/Llef42wideu4U4rRAXTq2yd1rSYhNNAxW+iYHJTa
UApsoRtDu1pBgf+WMqhZTwLPVCyMz3DFYmV/vQowouf3uxZxi0CK4xXZ+ciMcM3a2/0p9NR8s9+5
7yYolS5mbiSpl6aSPuglgsHOIbutkGYSGulpPbQ+ECKWHNvhaqR0TTG9bz+7PsmiSrc5WkVXmFcz
Mv81+jD2Q8Pta9mNZf+WZm/gbUJt61+kCaiHtuUmGUX/TWSdihtKjn+iJathvq04S7jPwfKcMN7A
IM8RuybKs8s1agHzFjjevRb8EFFPqbTRezrXNWCL4e5RK+7rdZvhlqkgLsXCF7m0ehP5icZYmLkc
Z1BGMYxCr8lgXvM4i5YQ32qJAkcR4lIANxsZXk24oOd4vENHYRPM3QCobtYLaltD750g6xVxMyJq
y1ZVUPufX4TCFAMlR/TAbeefTdUtAshOTm2jblYnHpwZJ51zmeZ5ul4koSg5lyxM6Ekrvr1GYgKE
EvbvZg9EVmgQSk9mNbaw63VVJArGagQopCcxE7C5B8SZSL7nUVTNVlknj7drphSOQuhzJ1bxjQ70
whRdxV0f5RhcW+D2KBiOZf4GawMOEiJc+hIiq/Mfv40YXg2hYw2r/38Wz1Lk+tFkkV4fbxeeaBsc
b62r9G40oeC1UbUaiI/kljQc2NdL1BxjyzX/vls4U7JSkkpTD1bX+5bbSfY6qYiia6oR2iHQnu7B
eNf71Amw60/+Uci99ht/iuh1rGH/DgnAg+Veke6CNNT5H+SX4Xg1c2STPc6X9YWLXkVTlVxPxoOe
QGQWeB3JyhfUdK8U6+HLtEh6gRmUjWE36r4FbtDP6jPory7DN3zPPlkZlzjn4YJsut1NPUElMfdo
N+n6INu1Svch5LBQoPNSFFjyyKhfDvHBnXxxz7sYj7efe066XaVxSSeSkRM6MpNzjiGZMTQAi1UB
ZlFVFl05mTQ67PGH7uIgTbha0DLjGsIN+6OZbWhRG5rBOSjtbdh6YAeFQxmxwAO+WGbH4Iux+CCn
Oc/L9MhqpzIICchMiM1N7MtN7rG7sShDw8bbGm8C9ZV+XBMGCx/X6RjneFzZRaL5Ew7gt3QqRLgh
/jTXvIWV5JR8jelT3+22YT/PYwn9+Z+Okc8GJhbcaLwQCwj/S1H3ETyu8+IQ1T2jciPIRUgYZKuR
HWu7eoZ0DnqgKqkhM5Eco0URXGqiCLIVQXkiwFzIq/q7A+tllBjqnU3W5b7BLJXINSjm0rtIDLOE
vWpk49Yy3JiyI6d6wv3+U8XoYKQaJgbUJe56bQpNQ6tsuB6/A68k8vihsA/EP24hRtvH6EFM1Wn7
hRNIyk954SU80EIVnCIBC31COk1y3N8OEFjh4ejQ6yFQEMZcw21NatymLsFaBDqkr+w9M1Go9UUS
+S9RNl5vJ+Vcs5FnrrORUamCwTfVtFaubA5+QbmgP3rSrn8VmOne+Nvs1RQRpWPazAH2U2tCKViE
OILHPO2btoD9kigBpb9XbM1pqYuKGHbT177O2QABhqZbu804QSxp1nPEAFT8YGQl6BDzaYlBsJRR
+b2l5ONOcmkAz5cG7nfqAksHWD999C7sNnsAltoj2z+RnbBkwi0/Fja8T4+E2flaNMJntiNIvBoc
vXgPpyEAJ+luXNB44tTF5U7IrpF8EUqrXZQ+Hukr1VvhKqwiCOVqYJZMW+y+OvnnEPGW5aPmhfg3
WkR1eeVp704KldADrqWg1m5p0umUbBEp/m4EjqJ1xaYzBt0KckE9YjNW3Ih34ruMOD2qMt5vkz1X
ry2vdxf/OTt9sSLnlEcwB2m7WDCE8iEd7EFlpM5CysOdDdlKl3mQRBDtYCIicctFXrKRDM5CtfgS
DnfkQGXPRELCZd7QGFSnSK35hC1ckCzmpNfCgf7q105vNM/TKnZr2WhG+GBg7EOaionZxDBv8fxJ
Jsi6DD/SdiUBShyqReUZglALWUHKS/lzkMZ+KHr0uwYpFaPRKh0Qq6lhTPazxWkx9L8DLSazdSMK
qeZgrzoUoYPkqaRckGE1b01l61RB7aa94eOOIt/UYPt9/Q/Ka4G5W0vtzkGm+POJwXzA0syfPbHR
WDtkc6f1Gm/vs2pqGbBwAqVwpMh96mgyAR6Mj8n1rO7o9VcZNhq0eb8wJifsQFOcSRhBUq0omDMr
dz0PJiP/33+RO/uAHn0mMWnK5gx0FDzQfiu0ryd4U9+ddDo/hc2eUWqKNAXDCSEx9WOdmmUbG4Ue
FHTVq5UysyYcEp7W/eVXfuPklGAoOPal3RjCjpC06KrD+pus07Q030DdXNPaGqtqP2+2vbtrboKQ
Z/+P4HOXfx4wx/c6JnwNxUbvdIlKX8zGfs2yGMoUOUXEyO8QirdPy/Ghd6KFvKmrkQ5ifcKGZjZm
Xni36XNCZDK58KK355KX0ARi2O2pQ5/2SSl+XkKWOnYSPpSGcdNB71T55Y6bsTO+sAKo0puVPJYu
w6ySfahnZcmINTygno8qwxO5Y5VzYsxCQSeL1RhBZcMRQnQ2ccO2p1mnwhUYeiif6OBv6l91VMNK
9xduScymjIKeUo9qPA7USjunyqIW++d5QD5AOPA64ey3uTU8qEyfPhAD/I9NP/10pXhSL2CV2kiI
oVQTReP2BOFkordLhIcEaNFhDFGLEqeRoCNbpnufprAR+Vu811U1JOQr+D5T6Ct8FWm5V75h6Zeo
zdpqtCLTy81/4C+Gq66P1wUFVNuGSunmpDEQCZPZ1sdlsS6flJf6ahrcBfRrpDBumeTTTu/gvGLc
Tw8SqBo2gtstDTcZLG45E4G1mDFe/qsFaSNzMZFUFdNaL5mY0sqWAa1kf6RoU7XGm0n71tkzfVIT
ZKKxQapevUqsuBlbajNMowKbH8ytnSJPqHxcRKJASYyi1JIlAFReBFWisEL3jfUTxaKhF0ZITW6+
SQCs9BkYOs/aVX7gS1M8tdl8haD722XwgjeAz8kgrxrsqfGSbWUP9375i5w2OVq8gOuNh88orqbL
x+pDUVuT3bo+25OLEWLMh8BJ/zgq2htxwtVwEfM0i+jSXCbGE+K8+VOUCEBzp8xXKno6nvYCovQ0
0zu9cBENQJJCvCYOjc7dvDPo8Lt1E1wI4TLGan6LHqFtrZBs+jUqAmKvuTnMkJvedux2AuwnEiA7
It87vtEAME0OBLbLowYK7SkcjrwFzeSMgPtjna2ab8ycDsk8Y/lanURTRNRPq7/nlCCseRuprGxr
K04jZFD2oNY3kxkHADtLejsFm2L38YIiQVOB3j/9xexiIe7VbvlgZcJvcdXYkLL3/u36f8GZeErj
LA2g+5v5eM5oL2jrNmeO6BaaWK6Y9Tw5EDflaVoClsfG7rQNhS6a4MgqKtrax+7ujzeQn5tzUeiI
xZTbGO3MSDEGhPETUf0J1cFpwYBogay/as/Ec1RTjGUctQiYAOcZ0iZ6rPyMEc2qwCqkfbmRl3sj
Mpgi46rteVcLVXc/Hv81glSq09ZAPoLxRcBy/4BhalpIWuXvsUM36PA5127S/ToFMnVq3NvquPZj
ONddYsF2eHPsOr2ZFDvFvh1EX8UdWuyJOzU5cfwYOOWG5An57USi57msljWhHC+oJlHByMptejIZ
HV7OYqTj2tkWpKTsKnot9F8RHItboSO0ArocesSpbuJ757wKOAdDEtS//znTsw2WtCUA4l8xCrwY
0SLFB5dVSdPWtt3IqxJgnKS0xnvTorul5YFJrzQTzOcyqrTz/MyKrvExXc9ATitMIp3F+24dD+X/
eCMIRubDxMmmx1yzHYPCdoXzjwvDettUKbZMGodqLA2SC9MkE8Ri5f2kZvccbOJCWjYSUnPG0hYw
HPnpmqQCMmpiSN8w1n6JRMvCdWaN4gUCBvzZeatuwJJJXCAtP+leUkotEubpvu50Kbqp7xbbL0MJ
yx99Wjoa1eXq4fl83UgXe1HtDMhqFfFSLbtEZ5jLbcOTN1K2ag5xpCaY/GyOf53Q0Eni4lG6I+IB
3DccMuxgo/QoLfYKLheMkcpUNqTgwOLnCLy00qfymOCO/srzgMFOjLprDNW6W8OVBU4gfckC3ljg
rYV8UvYgn8IAaCdWxYI911lswEnpoiCwsfA4y61b7HaZgYmdHMM4aK4rR12iewRLFUW2EDLTQ5nY
RKys6C2v+d2rzhelLXz7t0jIsrOBT7bVzfqS4KKxnweZ/AgwELYDt4fBT4/cHG7rQd+IrcePgnCc
Sd+Iu23A2D/v0QSfePl/wo0MAdtMlDV2Iw06B3Chhnpt0tEP3cqCQo0ru1FxIbVBO0OfbfhP4MPz
CfW9JXqM8DutqYJXhdrR/3kWIpH24JFSv/NP2LSfTsNur6Rse0niMxu7PGsAmzu0gxvgLK9YckE7
nngj0NV21YBAvO/cEeYU9g5l5ZTxFoyubScjViGG1afQed9Mhzh6jAPr6q5kN6Mf7UeOEp5pH9sh
8M7btN36fs81+m6noLs/UNeWkZ2B3kqkafstM0CH21vasDyH+6OKQ3Ev69ZJ9XOmC9k//Ksfg1wr
PB9AYYro3LfPCAl5WSOHx4gFYMyIQM8RP9L4kQP7CUKDk/GkEBw0azCq9Aihnv6+izboMxhHYn3e
QBurRf/lMJswD8pBsZTaRrZvcL3hOpFj8NPlTFLjg2xTY552LKODCZKTvWaB9u2shtRQOc0UeSIE
oAiBQeBUpJPjL/68XY619AbrQm1E5RLAY56nDiAGrKdddQhDGrXYxTHnFhlMWNaSjD16w0+I1Sim
h6v5Gt1dCw3PKWBVne6xGpYxOYM5UmdPEMArg5T8VxSRTvGTzpIuWrbf9iw63WVK8MR7j2tr2rzP
5UOIP9FGcEVWx+8jj4k3pG06NsWW0vj0Rie+tEsGUDc0kmjOE9gQ13qWWD8R3vc2LqNoC6I99M2/
XFm/cHhOWuiaz0+jycLKDhqX7WsJMuWRIc+5SpXG2DNE+8t1S8izlAFFpmpIUlEfmbvPmq3+mXxt
pyyT1o/R97HonoS93ottWWTpCAIVh9UzU/MNtNopVWefGgUdnAANFRHnYOhoU7WeOeh//6jcxH2o
BrJrwUrLyrF8p6mzXMVE9IEDeva5XYeZc4Kolqohp1yK0+L16uAYSKZGYU2hNgPCQsRjA+YmJIFi
ROhf89ZmH3r1HUaAtMI3+mbZVMBn45Egx1rhYuyBYtT6kfRW/hn67mJnNSzxr0tJkk5vqF/UvuY1
2LkCCs8DYf/TI+mY21IADNm8ZCvWssUi0cO3yOR8Glh4hIUmHRlB1+nv7B+wJuFoqxWESYqdsRPT
NnGTDFXSNxsrYldXt72k8Im7CWxsvU58btuEdMNJ/KlvM7Ebgf/FsxOOBM/feYjhqGzBRUDh1mrs
dbelL9gdijYFYxC6tCneuR0P2WrKARgkVZvuf41IHp744NoFTxmDhWZElajxoz1x0hLIQrfO/AIp
x3vlw0pCzDMAMWf9P0RDMi7XH7ZxMcTypZGCupIetgOEZgm4fsjo/8B00TiLgmFc1mLSNlkb8TbB
irOfZZ/QQG3cdF3BiBBpuTIr/DZVV58Z2ziVE4s4FvuTbl8UQxJBbWUjCkIie7QNidwqPUdMxEFN
bicAgsOMEHmbslis7b7gfDHB9tdPQx2DMEXGv9vp/KCZebh61m4Hz7DbsLZhTYzcRzXB67FWaopT
P6+M7RnPr4hA7afoRHVufxk2tMO8V9CGhHiy5SxNwVCEWMW4Ufz8RNXfd4KT5/sgS9iWx7Ad5rQQ
x0oC0PLYCqwVvccryRuHBF7ewD5OMiv7AgE4JBT1KAL0HQNuWvttuICM2bR89puGMlhFFV3YGvd0
veMbwnv/6iuEJAHi5d/kXLkjDDxMzPBVN9fam5lM/LGwKVXF2P+Pu4uCWzRC0SjIwDC8Syx2zLH6
+KwuEr0F0FOCMDCtzxQHubbiR9o1Bk+F4mhsUFHA3vYD/+nMk5JtR5Nc17i6iIQJKz3zg15JGzv1
8pjisXqyVi4h6kQ/jaPXXLQ/EmDQKSpUFsB9MG1mDBeC74J1hPLoSY79JctaxmqyU6q43Ti6Fe8L
BFYHj+6xRkwHAtVep9kZ0HWTkWSQAN38vodrDwd8H2eBp2lg5OgiR6TBG4m0vET3uxRA5y9ddxFK
RCrU8Cqz79rsgqgxQO31bIQg06oA0tlqj2Kg3PhD2zfaYY+7pse/TOA0ARbCEFO3C9A6Zx+c6RYV
KkJ8YXoyd3Pk6T0V2DxfwoqyavNmC8feoeTtSIPLmtz2RmJV9FFI8eLKVLW1AAf+K+2wA25wHjV5
fg5kjrBTNqssL/f0mUIfsOFXwHND/VN0YuRiJX5hfpkwEwFe5fZppXZ3cDzevhQAIVK19mAWT4Gb
E46ez/Fulix0Dj79Qiq+us9Vxtn0VObwKq7S9LISNziIUykL+7C3XPSyr0PZfJbjyCBrxgp78ReZ
IPdWlJKbEgHjSsGrcGIIrTTwmhLsqtyBNMeD4ZvHNMa8zhMIO5Q3KbJSah6om4ndlLvhuFLNcsL0
dw9/WG3nrd9IRBgtp37AecKQmyPV6SK50x0gZLkC6JqTqSYUOdDkTJbUwp0isR5ymlIVPKC6bfeg
y/IvDgnizJMtWlWiSvI/CjumzYE5l/8fsfCVzw5LQfD5Mf6nSwyNpW5rYdEfjvTmDSuIUuM20fZX
xf2fAGHkM/JVcMZJi/QP7eBEdjLIi23Dhw1FwfNiVZ6vNuWVHolTubcdiHLoeDXNSM1OmZqj2nf2
1BZlNuhR/nXGz2JWBt56d0yB6q7OrGw5CQdpfDMKV7C+HppGVZPRgnWwgkHAV2UKLLRx91dRssmC
GWXuffYnYGrGAXfzcfIQfnd8aI2s53/mmNLh/7CIN4LzHpXkyGO/7t7xjLhcNy+dEwcEzQn405Ul
W8Hrng8nAvXP2pGJrsHiiJVHUTg9L0l87TWTqPEAsHzNpf8y24yFLQYA8/jqGOwFoaP4Bi/YB2yB
y9aiG+cSCHpTKbF+LlnSJDLOJ/B0qdh/FllHaI9kKwgIZpGDBfhe0ZgeRrL4U8DT9yELOm1lOq/z
gYpAVYC3AgZ0FnOQIuWs3SRco8bKLh3eODXKze2XuQwbVXERQamOIq3fIQ6Cl3w5WtfixVa6rBBi
P1kcE5615l3GW+I2BWrVcD6XZf1/HJCHmCd0alnOxAkBDRqKpKbaAyPg6ySWzlKCD7up9QEvjwg0
BQklq8w7+x23TClCvDAS12YQoG9oTSarJ2oW0n4yxj9pvGzEoajhJui1bpaNjlErQ5L9pvSM8xv1
Am3YK2gLMShWP/5JtBijtk6pzzvw7kPyPomkiVWj3h10VsYa+DQOjPCmcsQPXZ9UIHOfuAEvTVeg
kyDBesJ9tAwxqsKAQIz9upl4SVdYmFnbsqCsqGSaxeoBCnwFVEVcVeQZ7zmxeKWSFS1SySF0O9Cb
JQxnt2O5pJ9T2mK6A1FLqwdCQnWVRjjdkD67Yl92my/Dw8q/Y0fVoG35ZthmYojfNkLmNDhDfXoO
ceW+T1fPTXuj0N1gKAtXiDL9hEM18jWa9VYbc5VF18Wm+0ze/+1ASdcHBf0XsbKaLltpfGh9Czq9
EfVbDXOrca8olDnkQzUqPh4bcIUn+0J+mEVCb8Ca3S1v4+CjF0ACIg/lU8v4/Z034mD+jCVofMMs
j5QkU35qA9tm8J6wX0ijw4e3/+8fa+aRtPk4qn0QNujnH93rjywr2N2OYU+mLkBNUeeauXH/MfOd
xVrGvjLN0E3HaEmCcK1SqieKnlBwpVZWNUVXFbHor1m5HufoykN1tr6BfHGDMmZ3oodtZrjT73FX
fg1fJ5AMaadxp4xgNTIDZPUwTDz4k6y0n4DBllPgqAVb1w3bta1Zz4rfaVqlAQF21emosSwO76MN
AjwsB/HDCUDvijpxqMYceu3zM87UCfDzR3aZ/LawGL2Qz0a2hqDtE8d2iduiH9lgcCFMn1xExflM
wxELGxxgWF0YZBKI3z3d1HPdshW0sCBi5MxQFrjpEZOYfcO92Ojo6Bx9zr+O20z7OZd7RBIv3v2q
08aB4v3SYElEJAUt4kls30grxskxTcDHYCtdefYNTEjjRu6oOzu1OmZomJDnsdwc7p3NlXsImqyc
ghe1ut7aGKFM2xdnse94ibZTLyk1fPo62i8c6WNZhwvIEGCjQ/HT3eCecr344ZAZVHrdzRxZehya
obZ/xXimzC60nJVFWmcKVPSS/2v3chMxZVpknQIHdoFWhyvyfioGE4gTWg2iGIbhJ59k12jtOoep
1tX/BQ5iU+5xsTdnqSGIE/fyqaO8PPy8cR1HhYtcEFQjB1Z/uHbrhEZrf6woTTBA3rxmawdBxrFi
F5GEBlQYvwbYtOs7GyibBlHIMsJw+QyE5MTB63m704idvfyiX6jYAuo09zIxpPjDu/fagKxgoEpg
68ib8C43OgJmH9IBHafu7WwBS5hYtAsEjfUNIaNrAocAyS+Bto2SQKaIWtIE8Kt9H9odfPsI9fTV
AnaooQ1FSWez5v2uzaeA0M7sYSrvGy9f6/Zm61VqB51SimRHxLGMLXzuCI4+N8ldpKuWqUVFEsPc
NIbl2W6Zi75a8rkX9Q0DG8E59Dz2/hUkIKi2NvtIFHIT9qsmsE1x/BD5VM0LB6bK7HvHSyExS8ta
3FsGLvg2ubZG40ZfMYxKSLLKe0IeYy43mRaQrNya8zzJ6HGe3zhbgKUSNXOO5AT0dNzFzxxLV43P
qwguKGUgffh96zaR49xNxAkRJ2wCoH7mxrf9lYSrs7VU41LkqG9gYyUJdfsJsFdxZAhCPkpyggTn
erkmL2ZS5MXOjRyJHYeVBECrpVdfkSlmBbUkt2MtxesMh0VK6mGGSdywXgipVw6rf7GC0/6naI6L
8areG3Mb3dFz/EMRa5BamDkrv9s9zH/Ezr8EGi1/kRev1du8CkNAEEFCXwAE6cRCWk/5guU/9xov
bZWjjyXyEvGLZN9YIHwDoGU0pmEC15jxozf2kGhupsbsDM55xGdneU6OfxqF92TRGn//B9llTEK1
L2p+STV7Rx5EoptkOCRnyVfkKMZ5SB7HJbSQc7bjFlUCtCrrmKy4y/zxASFkNCsxJ82u9uDcZv3Z
0fOvjMQQEKPJIVkhy0rCUG6s6NGaa2WMjb2IAs6d92gTzKZCzEJX1vrR+PTLTYxknaAB2LYWUEO+
FWWE8HGbBui6b0jF8R7nWHN2xQBmhve43S1Vs2hRasPYEkTNwyyVeRp56mGJOvSZYLyRRXiHIpz5
uj8da0oLV649fozZZK1yQOty+dT4mQH3pSJSGIBqCN4hYKeAj66cJzi3zzb9dfAbuHrWu1WDnA2P
ZuPrsGxD+/w1zxAN60i1fJVMrmvoPgKosTMXuguAigUzG9txlcGsuVCtpWkX6OPdBn+nxqMS+D4y
zEgMqYuw1m5ADMEAgfW4KQHP+pjUaFM4Hw8bU75wARelSs/dWw725SWnDZBwH8N6/L1UUCYRDFY1
q/NpTjxwZSQNMk/0n6hTe2rqhLTu9y4EaY2n6+VTm0DMUuymuqokPeBKprtGAMaC6tilEEFc+Wa7
eZWq946w3XBJWXGzTAOOLA8Ntd72M2rHv9fO7GwxAvW1JO4jSQdDG4kbCu8vEiPExT4oONKG3rDS
CCqZaz+ubMCnG4tXkXWyKTxhozc3+6vt0F8LK8myZ8J2xcyqTBi/VoufT1NaKasf7N21Y0QOsKa1
dez/X5cTwzLuR5sLAbcS/Q2eyFUQ4jAxX0grwdr2TzT7xMrjVrl4ZdiSbNRw4lNhySTDezf2VPTU
0J9upQSd4y+4nL2G7b2vSSjMJY4FRaU/e+YCz52MYwDcUBHdIMB4jh3I8996cKqcqwhn2RRvyeZ+
8jYqOxQ6wqfmgVnnoRZtY8qCiZ8Y/Evc8vb0szJawArm2erxUbGLkn+46nZVLYrOCudwanBBefNP
rKUe8+fJe4FsjyDv9OqBQDCcHXCnsh/CZGMPxJ6rwc/d0VciV8YJJfjlTJX+YCOI/pgQiIDA/1la
daCvkRHOmJYfmLC3W8P0BavjHor67EKng5hSGCx970XBWb7sodg6hPIPqeMaYMJ618poE3gugQhJ
PRJGG5Ul9c88stee/fWUe0ALtuplqLt9PNhz1NC7ePJW7fQtISGQVx7Q0lkU6ZeqnnDB4aw7Cs3Y
1JekyOCLI58GNUA7NzSEimeLM+500hhorcO7kgJSpoP3KEULstkiqIpfI4Vr84gwDQRHCFgXu6f9
zy7B2Mz6KG7EvHSToVYEMAM+uwT/2b20DoO4uJl4W5++YlmhFaVr8b989oOrjSU2cMovINdTLR7P
kJ2PA32GzLAh6w1ENsVvupbCUQA6FDGshEeQpRRpIiuXOGoj47EEnII6osQRVUmCAxp3ChclLlFP
UgFzgHD/co+B0wsxELYlfIOg9qvzaTpZivXc5lex4YVQaaENuSa949jUI8khddeX2quE+JoDQF9M
r8gjM4X/ddglHyui5J12VoWR2dFrn60wTZinGxaiH2z7oRZYz6rCVR9jl/YWhba8MfBvimPlyjyI
absBJ8hHyQu/kCYLS1EL/J+ehqHE97A1uz1J4ik0JPFQhi2s9pCrhBkOiAAGEFNXPudWQoapyHvR
hPtZW8lV7s0dhFnL/buMGjlKelmhSQ0vJVZ80GBMUt5S62pLycACQNAvA/+vlIYfz0PsgtS48kaA
t0DCTp8F1T94x5AEmWYroBMjtUtmwdu1nK5wYjoXtzbrimVnTagzA0p6BqLDGVttY1fjgM+tEPUg
glAqOaBW+rACHIrtmBqF6ip2i6w0gKxw8fnubXvZXlcNxX5zK8y06LQl6cQcqSViNC5Z6QvMwx/E
iWclb+RymEY6PxFdpTXDzeUmvG2exbElE+PEnpt08/9MULxF1kOys3iyy6JbHfgyuY1dRPUDMCE8
5XzF1wtQeIjo+RLzthrf3FwuUmnwjuwC3cj3XrSYe98lBHV+DpxqkLvhSOd5YsFynMVqHuYv5xtS
5JYg0dCXpzGEldd6rnWdmsNRRrm6hJE7PzeCCgjqXHGnSixHuY1N666dSgRHoG7qL3/NE7PBvoaY
WVdjVC9TwFELluqU/7LfDGdILlRpjOC2WAu+Q+610p72qW5lkQkHT43oJuKonLeChwEgGeIvhxy8
naIsW+U9SBawyWuyFGqgX5fLNyX7F+8OQgpIbt/8z2Hush18bXDqUAwp2aB6L2ftHsUA+l3V1nyY
aVX5eXea4hleILspNj+nUGJ/LHpImJUZTJx8keMGH0TvW4HPoDk2nfx5VINJEyRvM7IbFORqv0ml
aYkOZG9tl8Q/Bsf4pWh0ZU9J38Jor8kYqTySOeShHhJamS7BqaowRiVe/2Mbta10UjFZWBDl+iKW
Ly3onyw7UhEddTAXPo7KJofKn1Ww+h5yVFpGIS4at4oBYM0PhVcKQNJJJTHJqWzBfGm+mWurpRTp
W/+MRFbqeGuE858aMDLym27jw2Z/MQwItLnuyBpQriLlftRX7egAzHIO04A8+y9aKX4/FYx9JtMO
1cTsbF1V6+kOn+YJV52pvGXT5vkk2G7SNOgN/jVBpwWLx4B0UUrL/ZOUH1HHs4x7+0xuxFdRsnLx
SQ95UjeSPsvjtNzNljh5+vawcMscbhUBAfTtISQqsGTj7iZEOEYtPodH8OMCxNjddJUUjrB8alOA
9bw81elqDVxgayM6G8kexnVH7JXDAzDcFVKNLXIjj9Mdk3l0gKVM0zzPz+/S6CYiyG3lWc55rdN8
WFcXitpD2JqnMFLvBPj9xeQMxwNWqENzdxdzxsUs9inl57WpnXx30RXHNvAcMMNOl+sGKsdIMQVF
LEW32w32z6yrmpH6+jVeDRRLRo1XjoCQlogfNpxWCz2RSAFrZRic3tGEHYaWhMU4l3c4NTCqj/TW
ZEioH5XeKkJvYtJrvQEpgTtbiJwgFkntftIGmrqvWvaW4qSh33OJHNarWIq4tdUZi7DW7E0+3mHU
nB6f//CePMRdcwtfdbT9GI24xxuM07mTQSQbbLjaoMbyUORPneuOvNhx/kFnX0LrI8cUPBP1j6WH
gxKTyl9VCTEDhq+CeZZ+yfD7DeKDjC6KIFIlgav93ELvHWsX8OwfkDbrn01M8W1u+rs9hZeH2KmD
LkqnSyAzSrmDwKqpkjWHbwcnD5rSJkPwmC+KfU42LiHGRCOa9mYYDd4PcWfvC1qRYXTKmgziCKio
oV3/7KS2fPZohaadN0NtYOYH9uLPS5DYz5BWgtqf3lbIGH6Id8oEwRpsKBBVgifmFI85RCrYo5U5
GGmUzYtYQYkod9Vki7pv0BrNoYqHQJadKraYs3JsWBOxBf3URPnVa0CtWS2RImY6w34d9/mfS5PG
9qHptvZNfJmbVuMnpnpMriH0crjaBun8pZ3ZyAsSJggn4Oprx0fMhfpC+1/AtAHjATUqq5L2o+E6
H1M5mLztPBfOpdOlfRJTQS8DNFnDwh2Ji014a96/zwzzw/Fu9+GZRLzjPfDn91GG388dwRWoZWuK
ZfLaArba/ETYruwdG0PH4xUuMsWT+aC6w4xZJnp9C7LCNe5kDH/b3gJCy7qxxydt1WMGvRHrlUs0
DIbyELn2WtxuYN8M6pPnqgXlxSMRGWvxE9c3EHRFB5qSa2QQU59xY6jmw1+gZbRbCYecHmWGMlco
vF9V/B/zqJM+yYNuK7Dw7kkMusCI9CjuRoJ2R4txHcGFea3ic1ZFhDyhwO3V6aRoOWSxNln7TO9l
zXsLv0jl9y531dN/nJPL2X160t5STE/kVRx6vtjTNDCyqwP3UAnyJAC35lvK/137DwkefBb2P3KZ
OEw2X0SoIj57q61/DyukLm5uKiPBamql9DgrmYdRD4XFHzwA6M8GBMOzxSNoa0775FLXM1/Ge4c/
1f5kvUNXPxNXf5sNXEaz5tsIqHkVvQQO3Zz8N0cvbGfY9G3N/MVxQ8qbmBEyOaWGKU75UvVwg8EV
j/WgLyCrRjyonSX9K6o6ErI007uoXXIe5lti/onRnV64tsKYJ5HsuFSa2tlU18/SGZLPo1nGqpMW
jgSUey6ee5ufl6mIQYoCQQlfFyI5ViULcn/zyNr8swCPd3oXvcrK41G0hnfweZOvcO91QywK9D+j
X5dPdJQ43dVr4JDsPp/O4JWTKxBLWKKvFwSdO+yMDXFvPQewehi5Ot8kszEHoU8II2paoBhis8u/
nKtlmx/ebL4pvMUSXFtmzeEogro4F9jAy46RIspwdvKFiBBM7lXD83EN6rAdWu/TcdMY4RACx2Gn
1cbe9scdXvoh6N/1xS/4Y2okX4A79FaEVrr33wn8V07j8m79B/b8VlYzq5t5Oefn2sI5Bwl7l51U
v4u0t0sNWbr0Khwo5eqbpdLSs1gIFAeC0ug3Q7QmgQZUGXHa3q7rbAR6cDSjtxZ0ODpJt2egOMPl
F7ZrCNWND12yhqw+9pVNJ1OZU/wr4xg6TqPQkZVxWuz3veyK4N5jL2sUsb66D4wzxsglp//x6Xoi
Ew9IvGH0xJXwMHULOUQdFwc028OyldlPY+DABG2enLoYxDaIUGhVK5CkQb3bIwhy9Itj0NTnzsrx
ri2NXZsXJvxTzAzZ5B4Z62EN1cUkrCaaQtt5sY5gm4kpP/g2ZUhjlqzryGB4tx+VETQEwpywXhc5
Vj+8NSXKTdC2TfDpAt1xWjDSPDJJB5f0lHhnQPN3qOwET4Yj78rXgxL7Uc8RMASzp6u9qu6qD/gH
/7CPdSZa2DeruRCFOVxqL2d2x3V1Ib7Um9+cZaVx/JeCCgurOjl7JVK2b0AEgZk9UCma/t+FMqgP
2SSbdEW5HFZ84ApQ0bhQYYimlP52bPpA6anENEwZThLn7afHCRJe2IyxfZWb/5fqp5NhuAbzkI4B
SSwsY1OsPmENzQjf2S8hnH20zypS1HEfnAEcyCuLQ3gM68AD+dTjEQmHrqKojiRUvdvVE1jvfIc9
H0t28zhpVAolXuUqAurQdLYy6kKHPAHW2bctmWwh6+Q8M54o2x7mTjNoXGdbnFud+0E4S6baJ1I0
r8CGin487+AON6LNOA5Eqspxl92gBHgIr0pF+TcKmx0w+Jos6xvOxE54nzHK+XROS9iNk8GQBfMp
3MY/gRnZiSvTXvkJdDMnlsI6U5dwkSPu7aENzgClEm9LEMhHv1SqZRPO5nshGt7gKmIaRzJBxXye
QBlCb8MaZhYDNrHWourTgi4zJ8C/JY0xUwta/TR1cx0winUl4WEzSnrIQBEtkFpSi6zSlRLKPZ0p
chTLZJ6uYHOM3Bcx4THUxr7LaVfEIZh3ZAFHH5rywQUn62invAdvrao7gMU0nyxR0SKOVrXjx69G
PtNXWQvuKedQORp/MzMJF4ZUALWmozrB1y9P+YtW8zagBShXGqsJSCIPi7atAa/P1MA8tMtx68fw
8E3au4KimHkgsob7iUYuw4NRqaSvpIf1vgkeb31StQyXd+PfOcj6iGg2hQRTkIrROj6HB8sKs+Q2
cA/jU67uWQSwnD4MRFj2UlCgc+Fm/daU7yiFInvdWMmw2XSwE6NlGdEKiOWponm1WgReiPWgwAsR
t5ixXQWIUm9b3YtwtwX8nkMwzT4+uXMw6kVreHW8ukzOEdEU2wKBJW3mfNe75pGkZrUKERzNI7zj
jGxrSce9eCY7nPfLC80kQDkxOgoJ8b39wPVxhcgAP+e9C5w2gFYucY1YDjE7H7jxLirgAAH+rX8z
2/rQyzVCfijpwkHmnCEped700etJf1ZLG9WXm5ogFPbj0NE9kKInukQbKNOa6KZy+H/xOgJYLzru
Nv3oktwv5zDLhmCgK6kzcEhOukw53F7IBVK9Ib04FZVK1irz39S4TfLuyaef1mhMq+bkBbmmVCfM
iezaPLCFJFswffD3/B6ew1NSmyXwtWD/xee1GTdLhD0G2UKMoJNLc91X8oAOuFTrfbGuqXf4+wCb
r2OEoEbLvIqoK3y2mgQEQXYNpK0Waf4SbQS4H9N7tDWsA9hh8HCbIgMXUKR0c0cCE/jBWGCEquJe
+uBjPDoKc34eOP1/VsGgK1o7aTfL0Pw3qgKJ5zqZe5gh5ahS1sFG5QF7/UCCurQfe58ovGrd6wIh
yflZwOiB4JLeS8bgKBKDmbf/KfwC0qmV5AKb4RE2it8goqJV6ErcgKd3xIObodOacWahh3La77El
2YCKGInvRbkW6dXRlBmzdK+UKizaa51fcge59Kai9Bw0yZ/CASoGgsup8/l5+R8NDCKidsb3MJcq
3TTDeMo0cm+zb9tGDISM4nfRREDBRAu9OJ9jIKKN3tS7S7AHn/dQN0+9foZmL/8K/rQeGya1ucPm
tTik67jD/06FP2hBs5YweoohzBuNvD9251qt+QFic5HegFOZuZ6fjBbZv2W+iEg+EOfFLrvqxiTw
FSWpAAX5kzAZoGTbsFWCX3atBjSeIoiT4GkXFH23BIXBuONgwsM/CxpPA93QmQ7iw7RUZkyxt5n1
kxsPSngQNRkEMPMAc0TCvTYgKTPbQZvGcX5dutX5B6SjCrlCc/2mIV+BPHlC7MkufdFuW2SDVKMu
ehJ3Oomdvjre3r9SvDq/+O5+Yp470mUHpmQ5eom6w/wUtulzG/ADl+JaBAqfDlmvOOY61J4uOU/P
Vzs6/ZjcRI5Ww3mkY/s3v1CRaIfuUZLi/sxrjJ83j0tTAHDOFfBw0RQIZ+zzlSNzNt7+BRXvFhuE
dVEVtLeqyVJbOaULvnEYTCQ+JJM0k+ztpkKTdQ/h2EhNbY5FFFnryihZcGig5wuWVQcs4y+nouk8
fx9/+g+T35ivxd9P1qZJ+Wq05u0dPWtYm+nczqcx0Gx/R9sDKFFPDUUGoXXbnLkVZvvzhjwfMcDh
G6hxRzGSE2l8nRmY/6KwH9yJ/LaUvqIkq7Q5/iwbmZPC3hWypIohynPvXKq6IMBXCAqs1TrQ4XvR
ALD/PlK2+YxomMAhDusQICRegioAWErS/tI6cy0soFm5AqhGTqoe3xP5PH7wgT9DvlilWhZZXoWU
dOP+lkhcQ0uOus314WX64eG95tCjccA3z1+lltt4nFWwHkcSHFAQGoGj4jGGq60na7OcaR9jigsh
4V7dgOYNg8ss39TBdnDNMt/2+41dZI1IfD2nD+7gqtVqlW3PpPCSEIChw3eAHlQMsGimqvDgYR+5
qVXs9XujZQEnV6F3WqVDGfCN/E+fnyHHr8VwuZnVnt5eAJ+2BJk7CVa7Pnq/MtacNMMHoiZQDgbT
eusjkrVrCczSxfcghSHj+cNk8fSe7lbgV2dbTFCAOlk1/i+GcRFhsC5GVMJl8kvU6sZNPniDdAGx
oGU0ouyJOAqNwIFf/uVRpidGdWeR3uP/cxPeSRIR0T/9c7r2QWYwHHkq8EVH5sxfwd3TZxzswXWy
4BWQyINvc27E37fRV+5pODJyIPGH2o3iGRMnksKYmhg0ZeHU9mZOayKxVD0CQyJm1ZUJIdCpKEUJ
mk/U8m2Dsu2YwkWED7jBE0Dz659lTgJfywnTnRfCArHtruQAWFGBLHbFTbvzIOf+1IuuWp4c9EEU
MKtfS2lTcoIApCPu4jF68QJtx7byQnt6sMY0eGM2TfdcA4mXZ6RGNw4M8ALS3zhr2VuVzLLy3kjE
UIO9NpkWQmJQR1Ea6AsqNgeqwNtB/aEkeNXzowEC3RLnmom7+go9PKQmiZlQcF5/+xFiDwTEnQPK
tU2gKWdJB0NntX2YULumfUneSdYT4TyathEhFTm+afZx10lfPIO9bF8fijvv+IqpOa/JLy8PbUdD
tzFXpiO2cctyKEhmHfPjQhoYjs3YrjeXu7Zfudr4siPcLtc/wu5WGUhwPnJ0AKME7qiiPI3kt0b2
gPLk0GBPZ/YCweeo72Xu4P2i/Kp1U6oEhmQV6oxyY/ftjyrZZgocW603OQRoXeLAu8Gtg2946CaQ
LAWT/X8TX9mcKj7rLADJa0K/eg3n5J8M2nZC+qpQzhSSdBXS0D+pd+psz9UnkResL7G8EQDiTJys
qMkeoy+YMk7QNFtnYGEOwKVXsax1D/QTnSTvnc4eAlT2B6ZbTFMWZ8ppDofrVgP3LCv9NDJlQMNO
ZRvm1cKKd44ewPz1Cqwfz8rar1w+5+0ql3uEsQM+ygZYLowXkL/Fa6uR+Nv4nOW6+I4o4JyMg8rM
/J/upuq+H/LrgrJyNYNxFQpnrKjl94+kT00pwu6tfgcU/6Dc/ldM347uizQKmlaklJNurMrcnNgM
dvxhRd3N/039vYkX89xwjT7LN0n9TAZnOKiPrlobXYo8uL0tLAowvE5YPBmWgI70VcSuXGfAuAux
3i10YWXjQbCEJP6FPIIZ7eWGaKnh9IaLbCB7uPxvPt5NZCkQl5l4G8t5tGAh3sjmAWUm07udy6YP
m3jJmZdYuPe+p2SyYE20+eZt32aYWUKSq8g35VhxjWujDWt0ZaJBmewvzsOHSXKLiPPp3ZGnPgJE
I8ij+3rhOnF2PF86IJofv+rBrL8jTjetNlSUJZpJHbWEAEQwOBiMeiBkUqV0M/z4uOTE9AOawcUn
7G2KnuVSNuGX6dLsKf97FqacOjQXK44MUmoZj/P8UEi8kRl06erGGXQACGtbBU/lgI92VaTP3AM/
SHEnGLtFj27VgX2ZPHMKYE4LDbZuZYlGeSF0Oerr31FFix4pGOQ4esUsuIDn0yD9sglJE/5rjx/d
WE4Cz4ivU1DR7vZKs04gkWB8ZYBzRc1wAFsBlCBIgsg8nsOScwymmMY5oZA3zJq9//1BxJ0RpsjA
2dFemckDORrVPjx8iT6vVwQ6zO9ZEfCjOaIoXmD735KCws1pspf5msNqZHawFLI4PIMV4lAeIDWM
frscPcKEvwx+6Kn5yE6v/eAb48xdBY7c+M2PAQE5mmfSMu8akT/vGChRPPzZStxIKz1GzP2ki8kL
L60WqrgoWmVldFyqRnp9G8kibxrqe/+VtAD1lMzVylhXUFXsu5Uca7D3otOm9m5pJD1pbH58SrU6
m2lVpfvqdAk85Hmn+rQ9qVSozG6mInmqPB2Nh2HDFjW7kUig/TyzYv51W+K8pgwMueQyYNcviP3f
RbH6w3igOZtJDShI2/cZSMTIF5kCmGDV0NMTErwLg8j94gk/GiASY0CTAWSIFWyIr/ismHiQGBal
IyZ7goLo+8U1gE6Xk7/C7OBjl+Jqae2NCABSG0ENBz747UfdJv6QQwhfj47o5WkC8NIiBQ+KKTp5
ZRHijB26zCE6w9WQ+mZbZ7y9tgprRVBuOoSHzNH01G/IwJZOcnW72QEvSNFWcJ7UdpoRdCE4Se+u
x2elN7p6PQ1n/dl+wCTwi2PBjUkPwyr4ztg2Xb32N5sHQFVk+8cO1XuqAAl/aiaEOz+Xn8UWw7KU
Vum+u8bDjAbcKcrtVRrYkTVvB2AJH3KpEY2RV+JZa7VQmetDKwVwnXhqg1AB/d62cCm2G+36Gjq+
uXdOQSInAit0OKvpnb8wm7vvvyLWR0dvgx1Hk8vTI7DmT7wXZrtdo5DGR+Ag3E88h/9veffFpN4C
Q8gBfdCsForz5h7LyXWXjhWeO/IEkMchzI9STSlVgvClR8s/0dqdmG9QYs2d04xSxu7nxq10QG3q
2wv2SaKD56JZ/8Jd9+7ukS4zP9nOu2hF97Tolk8jyKiUYU025VjG70dSb+ySW2cfg/JRpMLs0h3e
ISmBz/YSH+PEhG2HaOsqUeXotIdYHBu+a5aIUg5MxIXb3ia5FoHFGu5D116GsoHecT37/+2lySgD
GU460Ra66k9qnhClunEYbn1HDAOAxl+0yewq0TE/HuvXLDcV7U8xSsPAGtUo+4lWp99rEp7/SsIR
ewxm229qgNmOo2AEdajlMWBpNQJCf7jXiIfuxfWnAc+ecREpZhhMNGm7NqWyHAUPoH9+/8Fg8UdL
EZ8aFF5z4JfDkjOTdlLPpXLsGdVPOj5H4aI+Eyi0cTyFVMFSBIkz5ejlIigL116/yL59sYJg6Xl7
L0ZMxN2MDfQT9zOl26x4rmWsmXIowSbngjLNJqaWRTqDGHsPJhEmyYCBOGTJMr7IhUCElFVDJaSm
2mtWZbFZxsCBO6I50FlYP/8GXG4sN1tDzg5K51/7Zkc4Eac2KBV3/ON0gER/YMYRBfgfw+kVItt5
W3P71TFJj9t4sd93MCy/6lXJQRNJBRJPOnSMoZHoIPq4xPCxafAfx1vND/7E5b7Q5U1hkenKKL69
At0WCBnfVeCC1RTJcSspuOO8Zf7ZNLzhw5EvXQxn0HUCsGvNYc4I3mJxKo3+t804SH9dv4eQMnx3
c5/u5NcdKcgCI1AuFzAZ9VSP8P6HB8I4Mqk30zzFKAx7wnbnIeSPqzwTsy4dkNmr9uwm1mSZPinh
odTOIo1k9i70qCXqFZgiuaCbzZ/R/cb1NWUCnp6DU1Ke09zSHGvIwT3tCEOls8nX7q+laFyf313F
DtCNAYKvoe1a+UNV/f9Cgs5qlR8tzKpYLxD/XoC/slGUHj01Kpoxj2JYyyw+tPWag1+cCaobHw74
Ptg0SEjN3qFXMYf1gWhcYB0P5t/ORPMdtNL+OWCtO0qaP6qNjMwU5WoDR50qutj8HJEC3Pf7X74W
aStzgO1tdyyaBxuxVsRbX2NqNadAmwiB1oYnMDPiNVob3YFoptm50c0TsPfRY9SQEyk491bRX3YP
F0MCQtvCsTc3RAYyEOLJAcTpihhmMmCHD44ZB+z9ZswbhRwIAIqItlJK8ZOlBsCwuCndZF/0D1Ow
jiGYIP0iKJxmQ4SVmRt7+vbI6URHBZaqtMAzJjBrLojCb+lhXWwj4WaZsQxJ06+uidlI8AOEK90Z
KhJK9WUPTRFb/BYIYZpq2o6PdpQ3Ksm21NXhac4dsuWWNhz6Kj0heT/hLlIza9HShgGoptdNAQKE
xUM/I1eWPZnAP7/1ySgch5yCWXrAN1JYVF9akDBZwJIMnqW02jeuIxgIdEvXiuUgYBedGGUIqZhm
yQQnhxpSPZlfsZu7PW2Nvz2eSYhNr1OjE0XkzJG9uqWQXbzgzExlk8XWuN6CD8rmYSh00D+CDqV6
UV8XVbhQGPOwd60dIv7vPTwZYoQzfmsrpH1541mG9E7aiBix/EdaJrhuJwKYzjTqRCcgyjcVEfqB
NZ+uzze6eefyLNfRADHdL+o7eso9rVubqudTkt41tjDsr/XTGqkusS4cuFtW5YTpnV12zAG5VMwF
+7Z0lg3kbLeMjHQg7Es0p1bTMVg2v5aNW68EZsbTSP6LPE9VNPpqaYhkB2KpffiODNMvd2fRbJv0
SEgJo9UslzOF062mhxx3HednT023JXX75syYHAgu0uqK/iUTUB0vusyCnDr8XMnotqhGuhkhWb7L
bu3DEo8heF5H39VXzfibR2GeTZhx/uERILDDhY0XboouSDJ34g+JhfRL0IqMx9k9JPLtgGSr+hMC
9l153m1f6s4sd7Ea7ahhmxmLea9/jHIW8ppwZOTp8P4I9336ycw6aW9LQfDs5j+nXyp3W/wajBji
dFQYAPTT1VI7o5QXJamEAzpSg8dWcIFR3aVrSgLP2VDRdFULCu0yVcKwZUVx33MadHjCdXNYgUrQ
KnBzRmvDh/z/XaV0zZIk5EUm3QKRMDriIIj6u1mqWjMQ1iXZ9+pfBRZ0r2B3X9gMFAF51Or7kIbp
/eBhTS/jFKr3+J1Z1ohvL97aJySvodehpAo6NBe7DQai2CtGms6n5rJUciki2ITiXPwH0chtQDXv
FnbQBKZKIApzlgB3hUP5Va/TmjlDzgHXsmYFriIUZrypHSlNhoDJ0DqGcAVIWmQTZBeG3yKBYqZs
099cnFY7rDbvTnnK0EgqRGKIxonhvnfRWdtPelpQutoE0LXCpkhK43sCrVMkN7RC6CiR/dTqdtt7
SIi1pPVr9MS/IkKIly5Ir5Vy+z4DyWPksIWwr+/DhcL8K8veTOCdjEbl7AcCPSzXS04LN3NdoxWO
D4MiHNWyBvGxCS5aJ73Tkx1OyKAK2YEw18hP3Pb9k4Ea/b8jZXtdi1dqmXqIdc8oC2BH1XxV/938
hfTCucVtDNPsCviCqK5qSaSGo4yyPuj6ERcP0NbS37FU21M0jL82nh1NnvZpFaQ2/OLU++q+e+8F
UpDosBwxDYai7b2GtnQzUkrnxymhH54y7oU8khv90pwWfBVOKWssZVOYmKt9t+xcLK/r3agqQaro
tMDCoK9i/fjE0T8nz1Gpb5IydJmBaOTO9gR69FKp5ZQOUvL8WKGdx233lYbbZRMdWv2RNkmEldHD
hg37g80y/HDNhzjMjw+DANffJhgf8RQdX7aktyeob0GEjbeTvORI50MmpLoZsQdXgAHwO0x9oSMH
WYsfn2y3sQN7K64jX/hLRqN8a8A2S/0AKP8llWDnYW9mdH03/M9rnNnF8iohslkYb6k53+fYa/27
UHgM5lMuRK756dmu5Jeds+ze/PYI1HiHVKVYeoyeAqDZjPlU1v4joBm3P45F+YO/iEwayYv7VXER
O74ZLvJDfsiYC5JjDa3SxtR7S5IfXxKZFP8sM6Tuw7rFeASr6fTcXz0Dp2aRyl/4Hxom6mSQJBeM
kvVG9KyBh2LQg7ONk8wzkuvfZcfoEc6MZJ5Ll3IiYOWM72eopLZugQveFcK/Q89iTSGAPT1kyjhe
96dvygzZujYRs0WjD6GOlPkGqn8k3RziiP1nn8y4izP4fv/fiC7+ziLo1snEHN9dV5hO9RPP+A5i
lKLxSar3hgAdcceA0jbDzN36GwSNFiARF+r9/jBnHZmwaHx/MWq6O8C6u1L+a3wR5+0vr95j8ZFR
4XkSy9cYn209F0uVhXRyrnW2mZ/J7IY/x6q5poU/CngnWGsOedXklPjqDUW4YMDe7eYxFiiTARgE
by55DSvOAEEoMjmWdVK8mnKgOhfiJFTRDmlfW4t7NwoxSo8jTnkkjtWxaHkItWCqLkFc2MA/rmFz
BOihCuNbCb5reKyfO4Kzknn1ZfFMWN9BVpUiA7TO5kvPrPudshNLp/PK4KGvykhar/wBrqIAIpck
nSR0zxF4jE8neCvLfWqBXsQa8I5oVs1hU2yScpHYrAu9PMt4tSl8E/sTzo6hYlBw1JFX3sKmB2S/
jiGOrBwE79U8Azo0AABH/GMXDkGCjBUip7FfiHXhMXDs06Wa687BfVjp0nOaM0uYx1r0K9tF2VJF
iyH5xpLoVTWi0j+viCzb0pCKHqKyx0E7l/elr5tvR3hGd7SFBHenzkUyv+04l8IidFfIld6r1dE9
yVPLi6j1kWyig7OFcXLjD2lYwLhTSri6H3wq1cDGLBIrGjFlvZaBvaKQ6DuL1geG0CFQAHE3lRgF
n7IyfVxajh9Z4S2dZib3nMNodTMf9GZAYTMdgdDzKFmV66RuKNI0unCYM2zQ+RPUkv8+3tbYw/sd
GQiCxrgM2KvBIl7B3XITI+/DZFwfLEfOXzuxVyuB8awOkrxpCAG0kIqr/Px3gILsWINs8kSTWTjP
26iNd4XYX7xBFWDIMRR6hwb5NpTwyoE+sS6bp/OLAM+Ia1aVMONPcTkxfswDDPErI/iDNJ/CExsU
o2dEmPg6O6lRqv/VjTyGdKS6DU7Fc7TYmLbTW2sWRiBqe9YdTTuN6s7aABV/z4ULeQIRd8WbqS21
nMNEaCffSYX80gK7Zc1peFFoT9s7XAa1PuT8g9u8zLHekjdQRoOmJiPaPawWFUw2O/jOWJq5hyG8
2DXKRK/VMiZGsKr4KgjFJ6Yry9Te8NaQZnMBIlDFMokaCGivPAlZL8l0oj/0q2XERo41tjim9TEK
WMwPIW89UtC73Uvw+oVnukoiXqK3L4lgdECd0cMbf/1K17Cbk0hlvS0oQfcdpsJh5HjRw8EoBDAV
ozQ6wS3UO84kde0kdv5NEdYDQC6r6jF7h8VtOcs56EFM3iWtWa7MP9iq0Aq9geNZCOiPD90lc96T
Nl6XU7LxfDiGHwLsp5DXk5T9I3DxParO8HhBz9wpqtoroD4N9W98g1in2vT9XlH8D1EaNuVB5AVW
gv/sff4oN/cMdXmbx+D9uYvvWju/Xk3r5/tlsd8AYIBZEgeGpLAzSGawn3771dtccoZs/mqMtrU0
wLwCZDMEqUITmetuKoonJAiWkyBs0rs4ll1ZR13HU/9TPId+OoxdmVvKWj48dooNInl+M5YNwmaF
BV8CF8sCHVxXLnQE+xlf6pNBXuoa3i3mqP1NouC/VSTSIGhycf9w6ofYYTtI1gVOrOULQXkONH7n
nyphLl3Mc6A0cCNcmTn5ut89BP6Ug+tkkZAx3sMTWwj8KPuyxkgMvK5MZ7PCrB8IUQYM9O15CDnH
xDenm08oYujLR2G0mbhBkq3sLs74QFQyz1O6Ks0DHmIlYeBtFwyPJALfBaLg48uyTb4eqcX8tzm8
jtlrEpu6t1HB1n99PJXO5RVCQP2s2ezBr8KxMBQUSeEs0xHXdr/E9/KQLOIIfnLCOEKz+gnmjhG7
rhpaPZ7eoXCR83logihdjKefC7Tt8n18YXvOuanol+xd5ya2TVQHDR6kZ2uLLpgW5OtXSJgZHIkj
eVck03RIkTtklLhYblF9y0wbOXOF1zzvZk1l6p+uCa5F3M5HOOY6X9/4od4tVn8VbVh1aZH+R5oM
m+4CDiEXBd4s65D+PyEU8TLAVbg6x8ahstuS6uWFVupJ17LKAvgR6zir+rkoagWGnlmJhZcX7Tep
Rk6gXqgPqJL1KnxmYeW/t8X3SJT4zkzUY0eQAX7QNjwqlprSj3dSPkWhgdRvkg4fZjJ86ETA5S5N
FnTJKP6NWAt8dEEthcc4+wJJN00H3fFEuo8xKEPGZ1UGEvUJP5gwXE26fXu7ZP9c87gBj2qb12Df
9RE998ID6V14sD6uVvYpDBfOqim97tHySD1rAVqMaNBz5gStCsK/iKYxpDYkPAXqsxfA2JQGyXCZ
VdSZicB1AzbiwKAYimSNKYMfe28p9Q+F39wDkbntLR5SgoMAR7dgyYYzrCovHNDVVk12wZG+0+NW
9+dMQVm3vpvx5GFMRCbEzqoIECyapuATgCW3fxtOntRA86tsrfeXKEm8JCeBxJ6uriFQx2jc34zw
HAW0hgq+rmtH5OuoccIZNZ/EFWJDR6L/CRRGpOE7SUzXCwBovXcWCV5Hk8wJ5GWBLJaqEB3WC1Yb
fDg2EMs2WAU5B4T8eAqtGCevb0g72ZbeqyyOIHwGWNsQQUi78VCsuT4GX5J85bIiTefBwX7aOQG6
3+fFJxBkR+EjU5ioOQwAk16qqDpE1qkKqLzQjdy6Jf4uYu/lA9j/W8akOZf0u0X80tNPszl16vZR
o9amU2bpYYMCr3Yx6K91yHM270LWdqbJFYASGhwqgoQf4TBzhxzDxRq/R4kMJoJtCYHf/naxhmTm
53qYyNtWCDD8deQ4eECZHMZbeS0Hx3pV7QYuZ50lsFfoOvUCmuhaGd6GlF9/PfBPX5Wt6XP4Yv9w
bb1WhRpyO/tMFmzeq7OGVPs0kLBQXJqoI3K0R/xDIpJUlaVveZ+jwdlnHrYjnw6jsVWxNsT2vNNA
7Jhm6XrmJxJMBZdlikKuetEKIGpXMrONDRKgMPgPJACNDk4x8u7/5lADG1cZw/DUUs+UKiHooYM1
ptlJsroX6TL8JvcE62bOJAmo2dTpExZfuxtdR14ZO2RvY34+LC/83dB10FDsR4T1ZPgWT9WGz+NN
tY8ISZp+KqEZZDnQpE6B+agBYzGFqzCb/DyCcc24U3skpjwP/cBrI0ncfeZrAqw5PWCYGlWxZce0
UR9OgrZxxBqbRV8P57iwxdIH0G3r40Hvqt0T+HUaUY61uoI/K+tGF8LM/hTj57MWE0CaYycSSuhM
guNnTuPJJ2FsZpxeWqWttlJCGtgSCwD6MxhawgS85H8ZfOCp4C20DOLCnkNa7y2irdJo5drGe9k6
lfXK9rN/I2neFgm1/5osd4X2oeIoMSkV88uM+8+dPZbm8xCCPXFPkwwaSu4Off99Ty1a6vlcGOGn
czMQMUAht0rXYCQ5oT9rwPBJdT2x2Dop7Hvuxm0qCkQBTMqUevMHUR0e+YIe5Z5sONzBZAPlOeIB
cj0+EaeN64zGCesgcu0S8AuWknlU1h15YRi4oxHfhGVALH461d+8dBJ9Vz+w9O+XbUqRIQeracu2
IsL+KFoXop8rKIeob/WnenqOIVF3o5/MbVvwjcwNr9qSz9ZfkHGG6nOuPKF7S9YX9UMkI89KX3v7
jFHM6jUVJ1EnqXJ5vOi3wneFcXTgmWliwb4T2mZHAu9fx9Ny0Xxyj+Vle4rEv0MI2jPHMkBeWBj8
TlHxTP3NgpYn6P2YaYMRHC93eliDeY/SbzBDAh+KmaKklIzQdRW1LNDhIWwFwZ3p3iiuXJPAmptV
v+tDAqExLDH9WgG+dvD8sF1JsDX5vxP0AlC2oX/WkhCKY0tn2FgGZA20pCFMHj2zKy94ZV3OEwI3
iL454zpRk8Cu0kSQ6Xv9Qg/tJc8rJavVp/rknRMDX7E0yeTol2+6EzqDRDjv0X5OExHAaFZsK8cs
SzOxWSt7YZ1bGA13YN8Roa/moJwUgLBm8fZJWwVpq6/Lc7VFi709DXcnA/23DAuAxCagCr+FtNaD
mRBJ6KQByQ0zgr/o2XXn9Ag++lPFchWJZv3etbLsvs41FpstwjeqfvuFKfxFtRZtJXspJtum+WmV
9W7NQ7z9oAZiB0D8FwsXC56lOeOLW91+7EOnjQS6bY1YGFD58LPOsSzN222nN967cYB+l3YFL8A9
1iSFIz5RLfqobn3VLDN6P1eafJtc5Nceb7Lq8QmOwoTzrgbtdACBM9XfptbcdWKY+u5kC3neEGXw
pGQBrnOpoFzcIJE3rRUnbKXJEzMJEqcx8wpYzUYro5ZTbXD1jo1z4ypBaXz4P7WYB/RNY1BA7Tar
IJ9pAXS5jHgl6yBwMiollbkjkuZyMrd8DfXM3zgKMG2Tc2Vsb9JT4u0CHFX37Ohy6XrK8YCzeiIZ
7VQCRpmcdCg56PqqP8LrWQVh4vusTh/mtfMb9ArPme9DEhCJacKF7qPRixQoJIQMtRAFHHZ03iS+
pAsmZMysZtulvojZHlLoHfAunX2WTZ8cFL5us5jIySkVLJVx7C4aZ7uT3XXqvFwJfDxF8cTDYqAi
G7hrmaVJWVFOh5Ta3iYYptpn/+dwecu8zur3EI9HbBO83VrJ9Nz1+G1djWQq33GjiURlUFs981IT
wQa3rY85HBMbSrWl2FGcnCG8CWbIZEygXeFApJoFERyB/mnwc1Bp9m0sJ/yszxGLbKxDFfYHuHA1
BCAl+huaVoW0AGfpyK47BD6vTvtkfIXDWeBkGKzUI9QPrB+61Hw+egNwx/sOadlzxVIjALkJ2WRc
yFJfBY4k6WVTA+x9wQ5pHLghw6ranoQnYLHJs6W0pjnMkXsnPlERtqFlj12e1vvtVQ7pHCkAJYvo
smxlbjot7Ve19QHlm9WffBV+EaJtrXg66zBuvlu4IDL3y4PaeUy7ZxhbpOxKachUWUcbMB4scejf
tz6JPe4EgQifEH2NkyWaap0has5AmMTRNeWVRfaOWhfVgwuXJbkpX1QsNUDdJAFQQr4yfQl2d9hL
WEYNkbxvSNgnlXI7iN1cFX6TYUVCORsX6zz7mjJyeEtbdnRbOfDIsUX5hgJiG1f8QYXLlN8RuQL3
5oEY99gFeule1NSSZgGUoGPqH+Jz2sbL2+cAG+cRrRz4ZQwiWnOlt+aWCzb5AxCNplBIlyM1sf5/
RfmbFOEIo8s7QIprOeiaGpTbprtDxMqhf5HSvAKrweiOGy4RMTYJPe8BWD/fMqcoYgdsjsZZi1vC
ah5RkpZ4utcPw5pZhHw0kspLQRYjtRuaU8+bjqQKZxpw67RjtiHn0yOMZJM4oCbB1wRKukby7yHO
0QIaCwoydXg9NHibTfLP+cNuaYB/+8vr8bzC2EQvMJqroV+zZ750RlPQxFDd97Hjgsmww0l39Aqm
wlSRQLJM/ftpPhr2Q6EV5ttyUxsAZmScvi1wFuuPWPfr5xUEMEqGSnkk/HYjosUvbMeFckbsCodd
S3rNbkzVTrqMPtU2lj21faPIqjnKJ4RmnTUpPGLoUUBJds6TXo4Sr2Q13869zcSabEQnNrzBYefi
QA2GW95yl931WRHP62KpI0jn/+AMxoRtcQzk6U/LWbZmH6dK3xnQetZkr9i9qzqJVBUT2XEby6QJ
kJuMGB8mIIZmy5lL0/yPue6X2ncARWZ62gHSndquY0SriDCI8k0E/ZPhOoZ4WCloOoma3jT/vjwz
wXv1uLOKTRWEfc42bKFq+dDGZXBCpRMBRdqBlS8gdY07i3xS7EBw4o1Z+yt+1CpkE88YJkTbcuX3
2pH7yegijn13gndwAIiSa+nAM6sS4rjr94A8FSw4SAx6zYKBAYp01Sp185OiFgv1oJ9udLKkKzel
darKjMrLM3Dl7tQ2TUC1g2liJFNuEYirklMYjGe15Q5Y4Kt0jPgQHFMR9YwL740vQDwluUgBmVtn
V1HzuIp0xSyvhcfg+XCpFTRhGqRV6Dz0qaSd4O+KOMunSrysQa1xBLrS4Shup5oybfMwJvx8wkvs
inIPPCsIK6sPCYzaK+6sxizR0uRVAHyAOy5BRlSIurqqKSHQtJOasNPceIBErxLEts8BkhnYR246
GEe2WdHNNRtskIQuhIDnQBzX7eYa9hzTN+513Aw3X/oLat1rw0CIIzn0GUxBCDMDixpYy/UyN8w8
IBPJnf25QFgNhD9baTJqndMzOynN57pcWxGYU3tOIbMK4g07qmhuwmf/0dlhGLZ3YMFLOyQ/oocj
k2p4s0mIURTOb2BNQ6vHd+Z7P+LVNmqzyDm6F8xGvCG8KSuu4KJq3eRNYspMVVRBvkav29ZRgPex
KjTVLKcBrHw3v6HUOuSegj56pYs9B5xn0TT9pvmi597OnB5rf5BJmVGxNqG/c8Xq4PxFCroI/grv
ZfyU1Tcnilh5Cehd+2vLcsOn4sRlR6lvsGMXqU75IPlXU1W1XbejZALM05RRsLNYP0Wu3aso/epn
Go/yuTJyaSw7BWfoFQH2mEJwRvJ0gciv/sXdYx3JLzbhbGa633df4rCC7tr3CmhSLsOy1C6Mq7hN
pj1o+S3PcZArn47Lxeq8KAPOfOlLPMBqBkONCcMVaUYP7osf9ZkhRPZWbEU4IzwoilpOLrIK4lBZ
Wb3tSdnIACLXxGXzvzcuNxcPB09jK8XAO5JqhuwL5h2DwBuiEmojgEqyie0qNrGktw7iSlpjhssA
X87Y3UzsI4FJNM/vKtGCt7BYJVGPRH5PGLgrbUvVuftKK8ftxEvBga7nQUR/TqFgXxqq4M20xW9s
CY3mc2sQE55B1rgvapPyCdKlYRt9u7Oryo6feZ2HGFT2qurogwekIddxHvGdfUV3KJuq6jvP5QkZ
Yr2+Zl7NSuc1BLx7rStkYZN+fGCHGU+m1G/qoShWrhUgPjwLOky8xUb4d/xO3wUKzdAtWU3IoHWY
/5aCauOOKxVAdPZpxCMmfk4vahTo9c3mW/nkXBgQjEK45MkLm3oew+EcwZpoNoUj2GHf8EXQXTUV
hDcTRf/zwsvDKN72lixUaeER1qZHF3gsN7b1yUNlT2zeiTsvmkwd6vOI2vwOHgjT/Aoi16Kw95d7
hDCEj2tG8ydGGgOj479PjGQ+wSFx2JFpVwdcQJRw0b2lh+DTQafId61lPgtDJ2q7LYccvMG5Asha
FKrfKFHmftbox4WCOix13BAXhgcFd25JJVqCHuYYjOt7dfUpyOj5GDrU5Kxz8MFAYBNOtSTzC4M1
tfjbZJzq/AYId5sy2tC4gU0T4usK2f+L9EJb1bEfefx7/Q86+80NhloZeYsyJ15viy3UclgbSd3Z
/OUB4fTbqaP/AV/5j9bWYguXGmFu6yNFc/eriScMcVaJtoN32nalcfBaOpGSX9CYd5BYxC/FIlLb
ZVLWPnRWuaH21sMLuTITsQsunztwKYnK7eXkqFY3cJDSBaHqLtuzv4cEDwl8w3YYz7Hdw4lEB7Lf
NpHtqt0pvlY6DrtwhZfaKbjpgDeRvpF/wO5T1UIfQd+z/HYTiZf+Kx7IL18RiOehKWs3Q1M9ygCq
NT/XY5TDb36PkVTNYu4jX1Z0PLeyjJ2Qe8j/3NDbdzK7fJSSBVnVKm17/ENlq3PzNeAgndVG2sGD
Q60H51cMEaCb+5DUQEqVKLg3sWvmNbhkcOurJzt+dun5fSTMPBp8J3Wdy+iANA/VvVcwh7gn2tex
kmdcjWHHmvRQYkqJYFtodxXLZvP4yV1AVCG5559VkWtgZYDHRKZUb16/zCAcMrjujymup3iMMuKx
Dw1CXRJE+qYRpP5Uo9j3/VipNJPxnuci2R7SSxxfy2Ig2ahv25+YxQKJ9Wtg4k9laTikKcXLb2CG
jVxrBI4PwUktyW4WOZfDCz/++8Wej7pNxxDPG0bmgLafTkOdzrmsqp1ZFf5FL++j6UtoTujdXw3j
wcAnb6B5ck1djPTftUjAd9qZ5wxUHpYI9or2EFZa2QktXh8RqazEWokVHCGdqagFGTxWC8UffZm9
TuNhfBc48RcC2ZnXmwBSAJBjxcvSh6RyL0zgkdvDP14UQQZdcgefe/pvI4pCYbE8elEISbKhvkQs
ZY1Q0VR7azCMJa1zCpsS7wx6Z3kpV2UVrFGX2TuA0tHn/ShmPIKnnlMQLXZbjgUEbPQ3xEizXOMq
ijNW5YhJnEgQS6L8L/v9DnTALg0xu9xGw2ilsuVW33h1E5vPjoyEJdX8WTgDRuJ36OzNma0hiVOe
JiWG6keb1/BUEQIEAiOH5F/XY5Zts25XMXN16jv/YC+LkV/YhIZPw/rHGoMsZsHloZ82IKJlwLJA
81/caIvrWpIZUapKrS9raLxaqV/Z8dCQmVVg21thICnbWSQINRZ/6+Kf7MlKSSgrCoQ3wp9QCsSl
Tk3knKrX1LHUTlHOhxXmQQ7/FrlsWrgkb863ChjxOOWSU6r2VmJ+p3fVAuTQ7TzmsCN9ojpDNUB3
Yhp+I7+OVJMmnTh8RbV+/dAwob4sKq14U1cSkEQYgytifJKMaey2h5Ut8Sy/ZV95cglLKPl6Iwzw
G2pQcFeGOyRm08axcpQWbbAE1p0NyJk8DhQz4NF9EVstZuXQdd04BWohq5PLv+uoprqNxRaEsh96
AKxQxcs6Jw+uXQ14bbNrS8hLbmJhcqxqhFux7h/7sfFOC09EQbjonvbJwBYIyj9WfVtTkLsDubwo
yzaJ5vB8jJ7mwIpl7anko5o8IsmEODtvR/Kxo4DTUW1j8LvnVsfiq2mUbX7m5nwwZL9ai/CVt883
X8hutkjxirTS/eFzrow+h0oBnKOj9JXP9C6W1257Da9RWZy/RJI0DEK0R8ZW1+8o5AeEF8uYgclG
sab1jUM1x8Kqmmnf+TeF2yx7/dB874yzfb/Ox11/GmOOxFPdhx7xgGADP0pmfgpZthPuEzVnmUCg
WGVB0zXXkiK6jWx5RxwYcQn0VB9yYibVhaPx0LxW5JXN8C3GGWgRsJcM9T6B/Koj1gYlU7EJFl8d
jfPWS5AL90NUsZNjFB5LBUkLUA4BABTAm+Ybr09dq5I9SXyQ9TNYYPzscObCGeoOmsBTS0X5hTWr
PLADosdgyuoSorUSoE9YbulNr0LDQXU/Xjn5H+svACI2oNSQIWp+ZuzlhtEosUC9IBBeFcgCH1h/
GtqE31Jsbehlsa4IBDbILi01/bSciM+AqOURHNCTcFdK3ZJuT1R5Zl5nPwPYysmnMtKIKy8jdGQw
w7rvMxM0aSe75vrJMSDJojWsm8MwXSDzJtVJKHmAQ68QZB2AwE7FtQKfeB+Q1VfqxDVwDevGr6mD
lb5Pa/3xRzaN0qUxyHPKJTmCfLMyp4Mrg9zedXYLY8Y1qsst54kBPQozCUHtmXa6scrJy45IQUhZ
c0xki5M8qrsqAgsImZWg0OSPT/nnMg8VYoO24bGU62jyJJIv/mll+McEeJY6yPluTMeD89t2N6xg
8a/p1pTddCgvUJn8hIGoTEM0ajhgG/IkL1o9CnH6CUkfo6zVWyYfOMqz8o0ug2IWnel8V85CvJQ+
btuQHRc2AunXHRBiR3v4YFnOImLVFx/aIRQM/Rl3FcZ8u2Gyxpf2BwQX46Nw2bg9kTButNaXDBrJ
Pe6xo9NbcBZZhQpO6RHXWWSFb844Kxj48wydXXe0GNuGp6OrgCj0gaE0SBUPPGpZ37gKZqOotM8Y
y3repdodNOnGT6Hj9Ci01ISD585NL4CxH9jgpHe5XXe8a6OEEh76s0NJxitxVge5iAMaiqKIKdgi
dyE2LR6zjt10rG53AsrghpO6tUERXCcPWeylBB53OUhE2niYMjSlcy2eS8QseAL/1w907DRxZ4Sn
l7GcLEWDrMhLgKu+j6eOAS3SP+Y0c2jTJYHHQwpLsYQuar/F3yvVmu2zK670r58x1w3NXiImNA3C
Fv0UcgVi9KJ98N91f2cJ42vgDCoH0gd74sNKFwlkogkI5fIKReviVd8I11ILotVpw5FDShw+jklM
U9cwRVTEtC3XtiAUU25LyGHR4NQSCsZOTdyaF76R+qrWCqkb2o1rcLXG9x3yIgxWk8ZlaEt5IFaU
CxFlItkcaoexD5dt1jKWg1oO0Euail37bnhL5T61QlXIs3gzGuL6II4XS7O0jbOofrBAMP6TK8O2
rLpiRU2bR5slcVo4mGq1DIIl5vxTHl57mz5XwWGHD4PsPaIGPq5BceaTod6GIc3xGh5pvhajlSwg
ZrPILCUdQV5O2xqC7PluYmb4MxI9eMRMcYz48i+i79hTu/JtrMP8TX/ciZK2ioYJhn36FgmxNEqp
9hT6IcnIv3vG+T8Vava678K+F5cUFjapOsIuNY+o0GfiWGtHrbsnNZh3g6527j8xOOwYhBmGjFmd
uIEbKyFF2ZtSrYoON4UHuuQf/IrsIsX9/+1X2b6UbVpQZl7IlvIXSPzRf81VD0fF//zg2KS8eNR0
6thTD4EcwmosClKI4QnyRd7XsD5ddSSByrYP99Ork9kbbkjTyH21dqg2gDkl5M9j6JPMW3mLar+f
eFcmV6ccqT6Gd5Bi3GDDq+VHlXu3PrW2dODp66rxU+WZimyeY+EFT7b2pSwy86aQwBXNr77rbj6a
65AVBmw2M36k3NIFqPGF1Hk+wscNATYKa76r9tQkj6C0X4Y9G4rAwbF6T1zXhYfHzqiaLPeSku82
IjBxtNx/EsDC7R3yu/r5uMyixNFNZGhJo4bAjcHlqninB6WiwduzjXS8zquvfaQWZptolbK9BKij
nizQqwH4H+FKxgj5XccuMfj2MVkZM5vqjqguJh2eOvXxIRIOnN1BFKwa2x+y5o4WhIs/Q1Kd4ZFi
4HTLrQKjPgajKm1mWKPwcah9Rp+ANJ8byBXDhu9EfECjo01rXp05LUBkQHaxxiA0cblZgQ6ficGj
+68OpmP7mJkO24H3TcUKHkEO9zCeLZqr7RDDFrLnh7f4J9D5yJNplOMFHz8ru+NPzkoVDWiOYLOX
xRLLsx95IxkoLrWa1ZpZ3UNt5jKitrDcoJxSYy8w1NrcidO15j4gB6rC4oyqyHssBycYRQH7rsLv
m2V1IJNz2djzLGamIpqq+sn+j3uaF+iCe4oWQ+oAxhjOVKl8MS7QX2AstR8YoKMEbOclT6XxoBts
uxBcYoxCaeEmIr4t43pTi4iuiwXuWXv8STuncewYG//YGAaoecPwiRl0Gqmkt06WWzdaoe8qcNGg
zsJkFZ5Ha/v6atUp6bD/oMoErst2qRe+5RTJ27Rp5OFvzsffKuRmADn3b+aXYmaMo7K0ozWL6BpG
XlmB+QSff5Tr8nBTKyjn7A/P3nWErZgUqE1iLNE6+eLwi6JMrNgr+Mr4Zo6RD9efeKh+HsnLGnFT
LyCga47s5+OF+9NnL9XGrdXygTnpRGw1rOjGY+TfG8d1buYiUVy/VDHXGEhBlzX+2b5625T8D4+Z
pApva8Uf8nzDivZt+E5KnquSex+hEPRqaKM+8yf7SOF4jebZweWZ2fFyqTdFOHkJqJyU62aTxeG9
vMHhRyVvvJxWl9aOvZ5kN+m+g7/tqcy+QxEnnThr2jvkMG9hCS65dSIwkB11CXidf+CKaXkenwXE
1/kB3YGq2qpLf8f8X7ua/DxPCasizGX+XBjX16rBSWeqzKomvx+T6ldNpKeJKum6AQD9M4JGeU41
WsHqh5VLRKYmwkIfYmbhakOjrxMXbNwER6X4qU1sU0mQTb4Uv7Z2VQWXV/EJ9t9aOqZAfh36v8yE
ch6mOsxSRYWRbCcJcsrk9r8JvWe0OBqHo6zCjU5mqfOTLh8Bt8gGHaGauMOOBckdYkIQiEspok/d
9Mu+GZIoD2jr0Vg/wbifl2WG39+055ysyGEm4RZyaWZ7JHzIQw38VgY3J7VKv8jxKG/v8OULXJBR
Q5ocO/reUcePHErBpu62hrhkiQpoQzD0U5qqYE/7YhZHPwBqCoBeFeytQlGUPuiX2qLGj2+bq6Vw
3P7ywdovkrMBjNL+eGomA/TEJ5k5liJ5dZqwJPyi0JqEsnT/VReW9xTLngU16zNRAkvsxv+TTiYk
v1h4Oaf75rkTEqZ1AyhbcnLQEPp3C5ptLbGIRqUaTwZ+HObP2ODQyrO75mBlXn+5jCs08tuKX3JK
9t+LSAI0kg5GgfsU3sJA3r/VJMpfoER72Tee4OyGYesPWK4AkSezcZ5v2u2864WePFanjQUWTm/l
elHq2R6Gzh4i1z8XOCNIZSFUDbkaktg4rCDswQoZONBNlznp4DeG7kDLlDYKy55MvzwJce45K9E+
UtKUWyqp3Kcc51WF8jvW44irKfIzFwVkWx9SXc9f21igosanYlglPRbHWt/u1daDGvQz3igGt43+
DQuOlufiBkZne4b69A3PxFWIJQYpmh6LTxtl5XY5Kn4//x2/bX81n0PAae3Hf8nm59bWGm9lSv8S
VDvOkCjCbDKTABFIHs5wAtRvwSolW/fllnEcBxzM6qcfRpIv3R7JJPKQmZNKLsXyIs0K3zwyDLT2
Rilm7tLunze9Q3yDSpP13ufOnBzE7fScl/dLbN74O+uSa7qW8uodz842EjMqN6ewI2GFkL1RGEv+
masAussy0XSz7lc8GV9Aj21e2uS8c7V/M3bwmiFPEBkqF2cxysbG7aLYfJNjKXfju+cCXvs6BKXI
ZPApOAiKMTYwxtK7kvpARp+EIr6VJyaBC2smhtFIz0V5wO+H9vuqC1if+v01ktubxnyqdH3ivbtJ
Hvx3plGLrHsbeZB9ME7crckHXdbCm0NT2P9mH91K7P2HM2cp/rUtxPnwNIg8XHO+esLeGjeqnOEu
fwB16xFmHTXV7YvkTZMEjF86wNu24ryX/y1sP2FpJ20dRjaB/NAjFJqhUjLZqGopxw1GvUTznoYh
DGsUoebcfGzMjfuKFLOXBpAIBkCmOFCbgLmIpFKsAJmPbGATn2Ez3QtbNbWj0FzTDryUZ7+rk39n
w7+UdDl9jyozGx6lYKv4lwvQjhu0FyKOn9ujAmjKQ6XcUSMIC75huMzbWGcWN2ReU5gN6IaC48AG
jJqaUqKq0vBfVCy4qKiDfaJRDCKPIxerpysgXdzCVJERCyJR9x2e7za8DAaO4SM0ioH2f79pU7/E
apSpBpJXIDKM32apJ0F/2XJwNtMkD/fuxzFd2cxC6C9DvKvMQgYCfIFyfo6tLxFtaqT+vzNrw3Pv
on/dGnPSdHadQIJZkeiRy2bdAMIfyhdpwsmqdXhGsxp11ynsScVSp3iUgv818+m6nTLAD83r9fZT
TwU9x2AW3bB5y01oE5wJqbSvkgD/OHIdxsD+lDAuw1VkdYC98bAdpCuUwHJhy+7SLhI1vaySsH+A
5MSPFaAYXPGfJYycoWy/7oIxLFlec9qn6SxeRuZd+Edz/lbTTSq9vXvBq1pSL8UZyVrkCBpQicw6
TffwnDQ8vjjRh7SqcBwQ1n5RQiZC25EGahNmimxIkz4V5FGyYa6hErJBpGU0S8o5zQ7t7k89PfBd
XQUTHkAtKu/cpE5PBDtWZH2FI/Xx8DBHmKLLYFHTtGRePE7LKO3X/z737qoBSfjRGMPm3R2O9aP+
q0SsAW1xVoEgjVlV04dYMvlXXE/dtKBEVuBpWZUpChi4UW/gXSZaQ2ulFGF0VhvzPTdsoGkS11NK
5SUNN0/aRITUlL/ukThtUq4yjHnlzJyFi2uhoAGBsgGbgKohV4bVlJDl+T8ddVVwOMLmfac3P+KZ
H7dcqOjsHVLFqrUD2Vm0bwjf3Kci/lnekvjQ0SfQkc47+Vm8FJrO+K7MEK9bWw/VMPxtkkqj5SMO
lEvJzEPok7ugm9GiodVqYTdUQLtrRUAKPWeulcC+wCWoyKHtBSefhlcd81dvlXncqVv7HIwf+LD4
/KMV2xw4C0rLA4fhq851Ss7bva2oDjfMgasIn5RGz/8c1EiKhBgtkRU9f+YW3max/BGGU5PqOlMH
IejZp7vsd/QbGdrXnlYfdVevXfTP/185lbzYKix5EU/kr8CTlJSuSfP/AVggSpW0DxvHeCtsD/zl
1M8/BzckRWDJ7WyYBsD6qbkX9dtvXMMuTcUJyU0nOksnBFcAlMcqQkDAHqyPmD+hLhLZr8XlFYhL
daI03xjKZxVaIwT6GA0VdxUc4KmV2AwdiIF4w9xXogGtESWmyhv9KXZe+GiMyulAj8f74g84JBF9
Nj6Rd+2Uz8GJNaVWtPaedxruAR1fgJ0BAtg4UZHz/r6+qetC8npyVfnSfe6SWqQ11vsYJ7S1V8AM
upQjR63TMHTWAtHXqcXeHrJavGXZvEkjF3S6ecLnHUCHcDc6DS8aenCcyKSUNcCbIX3xvhjImNWS
KhB1C30wPMY/IfaY8W2Mtxv7wuQWatBknuzy/TcwL4HHd+l9YvWh0h1G7XcVI1/pJLwLROu8AgrM
4XmbEetjelDF3PaGDXLbh0fd6x53vEryt+Div6Or7xo2lfsA9of5RX1s2szFGNDBWF3Na0dEYp2C
oFIB2CjKb4SQSQ5aDvyM0iaIuzKX6Exq6zY+YubhZ4aGYIR5l+CUAAhAfntxOKeeJmFsK53xjz36
rp3QEQfhO7QDlgQxIVKG3Y1tMY3bPPJ3wcrRsHYNYO/wqslkxJS1KgqMhNGiqnDhbaVMn7fuAKEl
L+OzgPLKSOkfeUbYad4SqXIsw6h+ZnWC0eFjcGC94z2Em1/gyyck/PyaE2Wp4lMF/uhhmElZbzXU
A76IWq7vEjqqDfpxnmsAaYaF6pTveUig7cZZCuKcLyvDWFRsIm+PMlvreaqOrrPw6eRNA5OseKy9
9n1kdDE44cMAsYLhkvor2wSek6c6i6/FEiAGtOEBgt5DOUjAF7fpV8gVWvK/2S1ee7dDJhs0NKaM
YPlG17sRQdxitE8jruM4CPbSS3hcGHS1dhjcKjVlBoKu1yx0wXa3eP5SBSSNBzN2n2S4ywCiUEUx
rl+GzJxsZHLCVeAwvmm8pK2CssqxVeHEBBAX0GRfqJhF2vhEAigXXX+cijGCPCqfuLvGNqPgwwKt
UyFaSeGgpUBO9R7hTL8F2Uy1cSPvKX6WMRijDaV6brzUAigTunU1IyFbDu4A4cSLSBIiovoQb4NH
OxI/2J0V3lhvmK6iaMTZAl0xz5l1zbHYBiyRuD/wF3cPKsj9XMOgPlhle5rhW+CI6aXu4tbMJFz6
GI9kIPJ3ng/5IsXIU3EXdhkqwWemwVEvVNM3j/OlhtgC7UyYpVxY9EzQQ1mRFy2sLjEcESljWQEj
D0IAaJ0y6LCTC72S6sEZ6ig1wlok8Ha/dZX5SL241xXm3yg1TPh+jRA2QBosuqwR6l++K0GFNtke
MAerN8ZD36XICX9Vuh42ICliYQ52Atp8OMKyJsvjhyMrKJeEbWY5wjZTFFTYOxiZS3bdtPatSDjE
5GdOTOPJdnZ/php1gFbKi9ZtJtv5s6oIcygVsj3VwqrJ66qf909KvslOYwMxDsMHP8TXRdi2xhHn
ltvrw2LaZWOvb/OAmofv3W3ejcZxJGYwOWWnDvXWBCkvKOrvp2hlBb82Wmqjb50+7M0UdxbulJUY
vur4Gwo9SZ8/2oRzzUm8zo6A9JZXw/JlZ25/mBsIwQ7yrc8kU/ZP6A5mttwGDv0Ce202DVmsBcz4
+1prGV3orCYSUstpGu2EpqZuqLyrPympBJF9nyn81cr8iKzT9onU6HjEZZOHwSaYOx0fsnzeL0uJ
JhxcbxGZLi6MsLWW/eUs1xJ9WxvlBiA9rAVX/Rgxx+ZQnlyKJ9kZVccRTrULG/JUo/odH0FmClKo
dqBw/ixqGEWcXQvecYy0zfeNRANabt8SjVVJklMse2TC2LAYPQtWkqyNDr3Ht5Fcbd2dxZW2Dnnb
0KzegiF5U6WkaHYiOmnB+IxRE57JSS8Mzb2lCMWGG2nZ0x68FfhOLJaZ+PpB3Cghd2X8roHc0Ul/
K/indw/vxW7jNG5osuh3LaegHkoqR3ERyhqMYm5/tPILd4Axr+ALlRVeoaFzvvjlkyaS8klOx25s
cnm9PqsINTQDaEpUruT9U7WJSo8Wu0O4xQhDXs6usFFSnQ8Tmp6RwnXv24qtlkYc/ScpufII93mM
hUSRWeOG2Cv7WbqM30tAJHxKmmmVBmHBzBARs5sG7j7rNLZSHM9BfVEL0apEGMeKvGNIKQfclIBv
giumfmnlpi/E2XSW30KLGIB4BFCd6fI+1bZUP5RQhUzq8wPdZWowiyMoOxoI5Z+a3deKshgUn3pG
XKOp+lQC4hWr5dQqs9VKZQ+rrG8t85MXiio4XiU8I/mGwVT+oWPdelK0UfxZKF/fZbfVcANPV1DM
AD4ZX0BiPL0yrKJa7/d9x//SBV5ZO2YESGMh044jKKbUhatNkEeQZeOLsFUA3o+nb2fpeD+uUpqp
H+JCaF/DrOJUoB2/EysL0oqMJviR0fk0dW1OVau8uhjIbAvfsqVi6vYJaqDFyv3t2wfbnE4NoRfd
Y+Sp2kTW1P9nx6uKX39q5ZJ3MlmwYS47VFItoNf1uGbxauWeYsaQ8Kkk2a+ena5Oe4mZ9HWsHERI
j3yLlvBjv2qOflwpUyhLfszhfLxUY6f5ChiaBmfN3uwg521U7u9Z77sydBhIn8bTbodnLEHQEi66
kVQrTdD/d4NYxZHIOiyFOcyyqeiVPLoVZ0cPv8XhKy5NM6zg5vLyJuHuPxJELYjpAPwXE3cp1KXj
jCW31dQhdfjlOK9ZBttVGmLyYBT4d1PoI/aYQ0L+oVO2GuIyRBKNy+D4Mym8XSUxu0q1KOE1YeQt
mD38pykKB8WG+LuTWSp6Up5zHPuvBLujUoiGX0VLZe1JWLPqfCELucCThOI8Uk3E54tDWCJLBR8u
wb7DiJSWFdsjMf0JKVZ8wP4vyWMlLwcDM8f/WfxsFyQRcTxQdMFH2OyiEnc0pEBY8wbEhA4zQWKC
SalJKdxlV9xm8vcSQHULktPN1a+XRba0rsqXd/VHu4SSzgkL5bXJJo9sLkUupy6ryk1eVGSDD2PM
3T22LF/J2FaAXbFzo0ztI2WMVi+RnEcT8B1Iwt48ElC3vE4FLppUOXjZLAAS0wGv8cw7Qjj1JvZ9
lfs8gw0fqGGA3S3nPV6H/SMC5TkTKm+CnD6CXKHMXyYgDDfD+4Umb1bE1aOGrzbgUVdLhu+qSAX7
/pyRikmx6jOMslmJ1rn4X3KWVtwSvoufkGEVIVbt91gipASXMHZCivlezx0JKHhM7yluSZse/1Z2
qMTVozPjB8h4UglJcv5Zkv9Wxeczk4SrQ8MqThncCHib7V4tT0xMFs8HF2WnIgop81+vaUPcIYzQ
LNZF60+5g77B+Fcwqr9FpEteyKXfz4E++V27bApILRa5hneqVkZbmNdqMkT8rfio4Tum3NtXsZwH
UKoZb/kjFeH1FBR4Rhs6h+/qr3RTKHuhubJttrYgjazCEsbWoihgCEccN9CaT75v5QKTUSyWeW2v
f15iEe85wESEqlDi7TLt9mwEqGrzEJGGOPMFbW45WbYuz4m/G3CBVCwo+Y0MD0fFxKOOQELMNGz+
lfa2WoKv1W6rpIbzf7v+VwreASwKgjhA6dYxrr+/KW4+V2qlqdGZebTFJKeSAgUd3Yh5CPG1FjRg
raJsp3mk4jJ+xIlxux7w1YRSdXYcaA+Cr3C6PuWIrfc8L8eEMfPDs57TTmgBsjzyt2np/BLfRUe7
9wtI3hebIty1GEXHrx2IsbA2LLzXx807CoETr1IYqhBlh8s0BEcXGi7GiC+Qk0nBpbyMeHsoxbBf
xiMlgOlLum/LOfsVbm2RKBjtv3aJ9XZGx+JHz2BGa+mooFs8fywnvdTXJuUnufScFvvDtwFu4edY
6nHN50zXAuVJZpg3SEOSmegZjywOMCoRJM9tW5gS3eesvGJLR4duu3DCqZAOvpTLQltQEBCrWx3Q
Uq7LCQNsWcNsIEsJlGfMtRInNllXcVxW6F24dR4Bx+VJjZrYY15uFbcF/HVDV79yrAUgGfM8H9vl
WfP2GxVwUYURqNNnZsrQGzxiXWbQK4tELM6m6yGmQyJ8nL+z7KA8nOC/y/WbuF0D4KzFUcnZ9Y6o
ZFVhu5SEdWrtQ/Mg0kebX88POOBRZ9ZsXWcT8Hr52HirtYSHZby7sAccksgpPQCJOJhfsO2zhT1C
VfJjCbmsq6M3p9VO5nKMxbuq37x8A4+42IoI/ei90bX/wGPP/D7y0Ns31Y/7h+PyUdqz9onU0pv3
ROKQkcKswscbsQ3o901IOCQqJ9Bbcx/qFUPw+p2mHHbz3uARAtjNgJ6FF9go64srMbW9m1P0X04P
s/V7pEX9qxaCWxaKmFhqs1SMnJlSvt+G1bAtKuseW3kcgdGHipTwNolrwEuILMZxnTvOR+CKdAtJ
PjNZeUBdqVI1fS4P5v0FgGHqtso0/ajHfjiWjolfbfT2v19MDy2OxoaYTYkV+s/Ca4DRYg+y6KOH
QNzDfT/IZp5yhEF5jZKH0du1MLNQ2w0kSkB37YWi13cwtrmmKc/rl23pXOIxLLkxeOTaoLmjpEvp
5Xxp+APNBjDXRMjKWVEuu6Uh3s4EePz7PwrTSKIrDE2NjnlLh8GzUUaQubZzzP6+GnMfnyVv5bdI
nOcyG4doy40Z9RktZ362dNmqsZ86OsbJ2lE1Fr38PrQI22fOYmENsvOYDblKvZHNH5mRQaBCkyBC
wtqoPGYnhYhahlI6DBqtW6bicfc0srJQUlPKqYKgT+VLu89ywY0KV0KTKOkBvczjhh1PZH32104n
aL8CFUtyPRbLYXPbGZ9P3t3ZyFeuwmle22SyaGMgAstjfb7ecg6ueUlznBLd5YiDC4Ngy4nlnME+
OS0BBWcC3qrb/MVdsdlwVvk910HOswU3PLSZZ/3cXkGFwUXv62r7U3G8FNTizzNXXK+eM7b4Cfku
AEasbVLXCqg5JOFVyB7gv5VUMmuSvhC/laVW31V9ejMFO86d+TSJrVuxCBXVDo3dYtIioLiNYSK0
NRtZ5ABpWhDpxR1aQKjqj3MZys5ahHCuDCVRNCnicpOz+23AZ2UuT34EzVpUQOxWjoQPFNM4cI1s
YsHoMDZYQ2eY4RRisZ3j7zFwreu9WYEFQnC7LWFZcuO1S6cVyGSMPGaubExryEt7naJ2osFC5HPg
mCOJS7/CIj/tir1SKONtuuDIiPPPc/DJqxbwga9pd7yQzf3Yniiu890U9A4xwkr7rM2tWYFopX2q
ut5P6dsK4xmbJm0q99bOhsyT04a61HpVbqz40r0l3RfTWNTCaUI6ibfi3v00r37ZOZU+CXeHPrjZ
BccfvZelhdr4szmzVrwzB7Boo/GmLzIdJm2/SsiM5waLQhWn1tTrXiT2NHzdjt62+RGr+R0aW3Bi
HqNw/Ds+3v1Ofd6uul8t5DJsPmiE3EX123Y80NWY34v9dwVmhIIVyX7Stwk/VqUby6c5q3gioFnq
M36llqF0tYCe7iPbg+kz1u6evH0BiRnPSS5oUGkHFXKRe/69jNNO2KTQ6bZ4ZjpFxIoD/tdWXi5u
/fbEQ1Tqpd7vDYm1tFCnZ26pKxuS2wkIGYLDeCbWkPwjotO68V8M9cj/JBXRP/zftShrhDNQ14bO
DF0DHXGfZxggcgqzc9n9od3l1L3ymKPJel54mFXsbkSxLw889wt7mGH+5Rt/2c2BeYy6dea+bD9c
mi/7wlyBBgTNqWUEMId5mRO3vxYOlCR3omlPRWZDd5dr+luTZ4CDKjESn+7Ozf3j+0HUOTNH9gCA
TocgMo+q0ePqVZimz09nWp73g8CMQpWsMyTFKL01WJcWDn0HqiShfaBiY++uAj/+5md0OJ2QH6ck
FKXr4W7N5+IE2J+UbuqdaoydvTp1wQ6u8q+4M8jWsF3VlU4BspMPTVxzVuM6lWKPHU5tvaxd17vr
TlYSsxwkWI4+JHnKSm33H+DNkLC03qJkCqZ+Gq/U1VvLCGl556rCeAUP1Jn2FC4dVAs7zx1GNYVk
NhhPPiYffHGprhz1sl+uB7oXYnE7Guz+cM5yA4KkcaAkKCoT3sss6I2doX9VvoU/e6uIIetZz4I3
RLiQ916b3waaGlNa5xzD0CAllM7903L/0kbGr4P0EU/lPPklyw8HCfPUGq1cqrNOVE/WBNrwXGH7
g5i22D2EuSKwMG0XOAqoLqPg6QLsyLEUcG1lTEK00Xj8WbVJqhjzUztjcnQSg6opPAaFP52xta+h
SzpGds3ms1hIPaJRAbYGqBVlOGqWRr1l7QkV8MajGQ1WWRRiWcsxoJ//UkJDxuCUzh+hM6Obni+P
3AN843LbuA5tSeYErA3kRkzRjQKAZgrTUhxBjNenJFLmj2IZR4Ij73LyLS4lr++F6GcIOKU+yihU
s+UmLfVXD2/2gWBg4cGrvFVH0jxoxQwCY5iFdoD+N8zoQfpuDCW8HUoboMEvtJlyUyDhcK+deBOF
KIQpy2ifwS0jWwARdE5O3H7HriRC584DzpVZB9er02W6chnS1yn2hhtQP2H/ONopUvfz96Br5A/w
goEwPl5PYGSYG9ubjSI/df6nUT7RgpMzJ8RkgxWeHmYGOWUlCtoUJr5TYcEYn2znkxV3IxIZjb72
oehK/0IF3cDns5/jsatpwfYP8vW/7/uHzq3Pp4AwO833nY0u8cTuIiSMnzGij455afOM1B4JSVjO
o7OOlaOeg8PsLgY1FhmAjAWL18qkQ60eUCLcYw/zagHm/pIBcSsDhc7MZ8uDgg6Z6OHZt80m60pw
Aze6gaFcz2y32bYW/u1440PmATgJR3YmXEcgYt+652MIV9rusEEoTWNhIskdIETP6rr6yqjId2UT
wMJjPX37XCdvD/IVI0aOrMVPLNykOf1uBvvMPl/XNSPOWsqlJZCuesEqSCLs+CkiaE4ZYpZOMh9k
S8vC9t2tIKH9CAakiMiKCYGzYWWivWzbeSo7w/K8Z6vOlMSv+NK2gA5bm7qrBvD3n+3r7HNlq3gf
GjXD1L1/3dtmR1hc99D0pWlD5KxKorjgpnWCdE0YIzOmK5UZkv0Yt4OOccwmj06TgSkMH2Ubhak7
Ib3duPCy+7xd3vQeBC4vV904VjF5r0s8DYfZ5wrX3dLugzoJGmyGtRnyM45IiY4gdpmAMBvsHEgg
VIKVrarwIWhwv2wzp59BehfvHGOFSUJkUgVMW2zQ59kkpH3QEKUG7zVpByKRbOItIWDJeWsmRShy
kueFbzzEiom93afyciweW190S9kr+oehbDJlXBAwV9j8gy7/g4OqOQdlfJ7ZP1uMX6V4gqFp0N0g
dpQMEaRpbE8EfWN5oqtcYVElBSEsCN82475J31JxLWMDXaC7XSKh2WKQRYnfF8eo4emvH31nB+rB
0XUiWFQ4UxB5tFQrb0g/B4YLzxJchnLb55D1IokvcUd0BWcyDzPE1PgiVjCICrF7goJnNO7WqKZ7
fJUUNtBgF66Kxv+orgrA/YWYh7nNcwGpX0Ia5WIrFBucn8EflPLk9LbhH11HgrI46pEQqrqLFNfm
bCKz+9jnoJAzF0bfuGDk88iNOYYCrilfqRNCRFzF4tVjQkXf4qwhDn3xb6Ff1N7H7DuT71h0pZ2I
kGAAQWZxN6ILYX7mwijvf2wBgk+a6F7eC4GrNAOd4qW8vk2+51nWfoNzrQvofkXUBZ6pYHQIcJCh
dxR9fFosTuEG6HdHOFLgOrTzy1yX8cS3UMfZs/etWYfvmbHgZatrB1MSzwVXEydyi2uO9s3/VND6
Shb/gcTKi5dlY+qPUEbM4j1gnO+rexw1hH1XyFVMJoMVTAlTP1gPctgTUrH+JFOXtyX5+6pXMD+n
aAoy4hav2wk+pQuwLQMbnxiceN9h/0x82BMmiryjzMH3VsIEYm5sn7XE4jjZsJ1nrnD7jmKvLdB1
5jYCXGDlZddTa+VF+rJstCYhOIWzyiuHGw2Av7x0kQoyOQ+KJv8CqwTN8e8W3j/xGQtAVF9jXd/L
2tCJZjMDVPUdHRrY1DUgCtMyZLZGVeFqcbyhQN6M+e6B+q4qFQEtbljfNE3m4t2+7qWYVeTMV4RW
KdOQ9H9SCxHDdg9kvAcX/U5bP8YNIrXgO5LH1mvJzHcj1ZxFuypQqKJPhIU0imlahU8XbEo2pBy7
TjMghi9R3RqpNScOkrLPQqV4nIW0x0vK/CDoIZp4ixLyIPy8pL+x1mXnaPbOzndVDeHRt/Ohc3ji
na6/agBHZOgXkpimIj5gyR0g7E1dCUYJMLIuNCcAXzK6H1riZdQRmTfoZsCqfjqgjzyNh15+Z9a0
yoP3qY2l7fVcCktaSbps/G2IG604bv/81ptxTpsYh+9b0dr6UjKRtpCWm7tAKgO5vYe6CWauA6Ec
vqUaYjfhcKZCi2dXEZv+INx7b9vJUzx7X2Fvg2S28a6t7X8IFkHefoxXOrQIWZIjUk+jxHEdurcF
YeHG6xcBoFFwDXJ2lbJUaZmskd99nzXlOnsKaDK35wBotrNLg6hQn4RZiD14tbJ0np0V74BfYTDj
7hZT0B42nUmDM5nNdXZ4tKbSAtrR3WRA78dY0KXqU/juNZRsUtiHjpRvjPD3BhMNjjC9Njr2GgLZ
AZg+2KgVHf+sa/7KdtDjUKweXAYNQxEzgxUmNJJ8o6rLlEFYq7L1X43fiUeDOSBSDbPhghKQShgm
vvz0MVD1h6wMDEmTnYbk9XtY2rRXCHxIVJ+hsQdT2EMLZ53y1Ac7RtNtLGaNWc38BVwf9WbREvVW
b6tkhaWtt8WfW2U/dzhvo/k1WGNQgvamqOijy0nM6iZd09PfObe4joWj55/fITLu68qNzygwNJuE
M2KfCkrf7mZ98jpaq2skayuE41BjIlFNh74S17o475FurdCaw0cBGD+WF7pFLL+aY6OjoKt+CuNx
w1RuGm+FoMe7/jUJ1Yey/v2CGo7fH6LvZYxZYNgkxbKI5Dpm4fXn6IwguBxUf19C+rYTBhMr9uM4
9rwF+d9yZUPwXVIcbCIrkS4J396nc/LY395XJjR0TXpn8mJu5pJPAS42oreaLVXCtIzhVEGRAzf+
GyUe53PRqHBM7EkiRCv61PtaTUlq+EJ8pH+nIIeSaekuHUFc9i4cqRHrEdUUimIID2dieR95B6HA
NCtiwClvCuyqksZG3bEslGI6l2izz/QCcdK6T6QNYkBUXesYcT9MoIayU06DptThnAXPAVx4a9I3
j9HHTqFX47vK50F7tsRoWtPQmTqpYWm+j21x28Fp/+AERRRqCI6gKc7/u7jG8awFJ+BEuXAPRwgu
kDI0D0HNInMfqQ1p2RbuFqT9Ps9a/qvISN745MmRt1GKiQ/oxUWn0vIMvOSsArlzoY8Kj56fd7Yo
+TCWMZ22l4jcUdQUaN9/zG2/mBSvBttYve5fqTrtD1TyARuSmcuBAcXi46rA1uCbfGsPNUv+xEwr
rR381Cu3mItyLIfTfQZJVgjGhXW0MbKFzRF9hXJebk1ODwTawKAg/JdlxVPMq5BqyfwAmk9OJBzt
gkuHYl/oU2gBfUwgHwozzcbVwpv9A4zRoFrYBDaRD8MLPPXLvM/tlOBnEdeCPs+aqaxWFUTuWX6J
02KmVvQydt/A/GHLYw2ZPHbD61clhlXHehXJpBOxZN8XIqPz5ik4VX4gbRNBXzZPOLhG0JM56dpq
jlxotVqESsRnkMc4KmSiPq7KnuSQ8oz2DPn1AH4xXaJKxwY5mWfDpVJ7GRdPd3cntN87/mRAIlhU
svDwKb6WW1jk8erDkWiON/fJQZ/nW4eiiMunVPcerpoqUeJbtjvr3ZGdF1BOBZ+pHVQmCI/tZadI
sy9jxLgEC0URlPhEImk5l2d4pz08yQPxeBaGebTBagkgYoFBkPdaXj55YNVhnirbJZNADi5WmnuZ
C5Xf8GQSx7z0ddEUEpcwtcnDb9XmHGrIdpqDASYNcNv6fdi65P2eHJryN/ZUD88n579Jwab7xMhJ
oZAPO0nvUQKkEa7d0H8+4uWkzICAfBbagoG0tTqj5B+YdjJyxj9M3gJ/+vjpw6xaqWPld89l1vBa
yeaPesfiaZGP404Av23ZKGEg63zn7HuZonv1/muXuA7t/umQDw64/y0RXK1tN4+htvVn7Led2QIh
vg2syXK3Xut5768vfLbIc6BSLifQv0trIxDuu1xQG/PSOmXoyVjgX7XIw4i6pOlwp6rpUBbuUF6d
ohCIPzfuguYkaWlUMIBbmy6/QK4ArRURYToSlzeJhtqg+UAwZ315aTBmPw0FWoq7HMcOrgy5CYRe
9TOZVpN29/a9k1GC2kYnyGyUsQD4TyA6LqGSe4F25wxmXVGDaHRxKkXG55/PrlsUvsP3fICdW0OT
v85UtZ5ZUIFqSbEcdVg87Zkd2oV4fGE9/4G0V/n1URzAEl+2XwgI/mgJv68UZoU6Uw3WQUCw5mRo
vs20YCAuE/kwmzXHqj5LfvCze8mF6Qh7jxbj6ZbVvJgVJ706p9AQI6pwWGzn4fstgPH4GxYScP0C
VXDQ9XQq51ieEh6CxL2buzPJONNCMBZTrpbH/eItL/XVU702Nnl1uRe9ZSgKg9j4LRxcJCcUrk9Q
BI6PKNnV24J4y9dPcsbYx3SOXcwAahqbRXw/lZLVDQvoNHhs86TLqR4U45RcTo9AxnKHBUdzDY2x
mRC/qH1FRIeU++PwL/d9pECuS1wxMBG9Ld1KhlhI2J018giSKUMwily4SHUt6XFnsmc8Q8vFdKv/
BBKDW4d9IFyv6OkH5NYAfmoU3SR/73j5aHcsv8YhDgZ+OF00oQn4vtODb07K/Q8LL8H8Z1gvpMzm
i4CYqew8MRDIBCcw/UwxJWe6cdckRuYRKAGHj6x8WSO1eg/+rAxJKyHMVP7YZFPiKRCtUprdmwqG
NUWXvRKMf25yHbJynnnJMTo+m7lFkBjATbV2buNflpiUuzDv1/3QrG45dxjyTt7DQGSzltjEQODT
SCvXs34lrP2uoykCK/bYDQBfrLuG0YzcnGkWV/YFQwpVCglS0PJsvr3ncGuLa5Btikn+dTHs+XJX
+ihBrvtMTwCTgN/gN3mlgITLfIrzfaAqC2fU98KV1ptROddoNiUQpTyqDejYG4eoKRx+XBTPf+As
ikhkuKRwZfcSttQ8Mdsln90oIDNOVe6hDWKzCGFWCO4OWD5sWkTKR7Qs2K3gI2l+AgvkUNgiv67M
k50v5iXRl8rkV3eWcz52BuWuXXdW86vaht3VJnDeRhzpo0RZ1RLBztsJYq55XMCPomNt7S4E2wKY
fap3ZuAKJEoynQKbkzFTUOdmZNNAljZwRrz9eI8JZcaxSpEKf6D2kHBUDIsmUaFw0oLAgz+nthEW
I+v47cAGmBEqwRa2VQxPKA4Zrw9b9cxVhMIgeOgu1j3oa3WoYEN99cPhyXSzQsLeuw1dCMmg/pNq
ijc5f4JxNqGGtBn6IWFUT/IPKD6kb5QPFr8sIfD6F89bdGj9A3iHWabLH310b2Hm/+O+plJWfF7N
Ahlyi+xuKPOZu0obVPk/R8WVj5F7RSDMpdtYSclTBYanAw2IN0nc6AKimPh0O18wzHaOYLjWo2xj
HkLncH++qW5YQMFOUKcUQ4dwvOgcz+AGl1rl44VdfUKDAIyqLYeXDnRclqHSGMJr111BwTJH5dc4
q8XnTkkJG0JhSEgE0lQVx/PB55XUY5irLauQyhh10OqKNnzbONXZ/304wig+CgNtW2sz6H1Q1kw5
K9Jfnx9TeCWdUK0CdlFO1lz0IJGz2dol88IyfJeNpWpK5/iAh8f+CCy0Q/zXr0MPNKXTE71zGBat
7mIv97aDB2tf8p+XnKhWzYqUIg6GuBJLuf2FcQYjyuyxCXwX4AwOD1yBRTjX3hemL5kJ49C1+Q2l
S2wuXWzpq3I9asYiz6ugQpwxe5Tp+HOnivVigpp/C1DGTpJcZbJpn3BAXb/QG8n0HOp2Vi0912jK
f4NyLoOWQ5ZSh5m7bgOdciJWBZh4xeh+6Lm3MKby0r/QxKbqjOge6fVz5SQoGRViG4gZcQjluPfy
KslwamP8JedAXOZhOsVZWm2X/gl+oS100DxK+LUS5dz3G5DfsN3ZXQqqR6GwTsXaU9j+n324nXTO
uJCn2F8xfEiORS9uuEbmsvm2xco/VOlixtKiJjkJciqopSvwUrpzpzkrgW95BBNO9596jVdWWxtR
kVlUU/fEdK3JIHxkkDGXxQUftGIieK8rD7cZiV+k5iUcjdEaTiTtacZ/oYmW9lUOdSItyMdM2P37
9ZyRtw1mtuNaUETPgLmqKNMwPWtuQiwjnhq4NqBVAcg3XddluKQb1U/aoh/M9fhMdYC6RIt68A9M
SE/Kkl/vI9wxffHAYK4WbIKoSeS3okAOVQxsGEQwrGWexbA6LKzZGjzOt5a5usskHxmJdwYYjyJD
gK+tgCTevheGBOqPccWlO81hwJ3+tePhTGnUS3fhlxvhYocGKmc2ue8A/vcKNBFIOpV+XDXwGSU5
qCrba0mKIdBlry0iGbquAKg0rMIxjDBOKsFxYYcSTj0/aTwlzumyIoCwR85hN7sHzQEqRtcxKG2j
ET2ldU5kMBCtTRCKCH7N7eHRTwzLM7HazPMd3SWGdsSMou4OlIeRyg4VtQp0E9FMq7Eo7PhUsTSt
R7SkOLHGKVua/SaX9+6OrbgzZfz+PYsKxIxlxwCJNYU7wgN/iSjV+Auu8xxZ2CSN4pgau9e/2+hz
Q45mAmwh54rxmoEUqU7RGvEhKKuExwVae5C+HvHMYw0cPZ3B3F6gGhLcPPekCjmCPpKb7gRFZ8Wm
v9GtTvaX3RoccMWnx48nbPQSOyUknIdZDV20f4rvvI9mOPQV/FhXgI9NWMzRg7e/zvM1+Db83jc3
bMIsErll+KbsUPoqlbKhga3aF3UJbKYslNZxXFn7WLQ8hHyVOv12v1yS92rWQAsHbdFzwDYL/Yv4
kZVu78JxddJtIMKngMdKwXiMHu/kMi24p+1lIA0++tR6+FNFVXOOx7M7LAyzau6vjS6QBZrVMeAW
wPnVAvw6zds8bdJobDMWxQEWUwlYmR7x1CvXwZu9T/ox/8HWjHiPpfmJ4afhG65OEylWM8/rTfC/
gR2x1vD2El5C8QIL995ULXNnaczpdwXatTT2mzVua3p1I+XslO9veb5N4R7nBvZJYGzNG2aoai7L
QUYviFsckDAXobsS+CmVsOY73IrbxzJ9W/eG2KGMw0wtPAoQlXsNtJJWUU6yx4TK6Ka5BtMeVp8p
lp/f0SPbOkAe2arYx5UEs7k3LluPEboJcjffonQxBWuZ9dw3pQP4d1wZIrkMJbAEkHlVGS+3o2WF
Cu97WwtOXU57gE7TmBSfgMnoAF7GwBRqTUB/APtBOvPz/AuK0mPhN9S6cAA82ezb2ZKVumDHNmZy
V4WV8c7sgjEp0vBAilpfFwq04KcToZ8YJb8QLXg/Lei1tyEFAyA6iSOdpZ6+fThgELwYic5DGGJ9
XMmWhscx5OoHBrGMJ23UILiUWZkm2Q1GpZYKdDreorIGZ1SoEwvOlStddcC/apCU156ORhSFJrmO
9BCDRgU5LmiesXNn4zhTSn4Gi8XoNwm/vzcb+1TiBHBpuACiLFgw4H2x8R+L48EC//q/3Whehnt1
hHIokNRShNRnML+lNUgwhYPxNX09OA+JowHNHs5I7moFiBDNdDtvoocLMLKLjrGjURGFuYMs2H4k
avm6+jqUTdsbE6BJMcWX7BXjxczK35Xzxfh4gxbvmErKfvE5ZZ4xX68bVg0TUjG3uauSrW/JNEjO
aB8pfG66QYYkLSYPUwEG+xaNlbNx0x8OXXl2SXo3ufLh1bXn0uCSv6cIyWWm+8yq+lYG+5TW09xQ
fjsVtOyUC1/Zb4ioPrxyo10y48HhmUZ6QhilAjFiQ3Aollb+hF7ERvn0bW7jbtRCIUQ5ZIvlD+TV
i2UyOuref7XRu3mk4j7FfL8Z99cbQZGgpnCaYmwbZw4hJ9UdYLMP4PryFda4VMcL2HUW2J060ta0
pl8iijlMYVMi2+BWY5T6KRjg/3uJMUj+1Us4r5q1vaOKfzIsfZd3nUWZMCbpJdnYzWHHWrIeO86w
gjy8sbimNH+AL2KPQjZjowLnMuML3Nir8/ElfgJR2E9imjt55+JS18LjWDPsVUrvijubeOTsbS1c
mEkbUte3l4PJc6CB9fzhaMfHq+LMJfRvy/GikjkqopdLHB6gOrP/JSG1fDQtyUIa+mbN0KIBRpl6
JgU8h0yEitnKrujyZJy2K//yyW3gs7tWaN9BSGfxz7GoXsAX9Y9rX7F+ph0iI8Ts+zIRi1VwWJKn
rRPiqPlouLutdNpstrSe7rnObEAwpD1aVVzKx/aaxn4PdBzf/X3ZJ3VNElC2Ln6JZGcCWJ703GBR
qF5AIs2+tGQ2YYWJ/jHiABrvQG340S1QactePhWF0gFMRkkD7PjrQoR4CnB58/hXtkrBPS9wrmxw
JwycPUBy0J+jsYY9icCqHw06GfquF5Kn7AfXxFU+j19+AW/DDS66+dNDSArkzI6cP5PimdGmgTey
P/MojElbUxL0MUoVE8Gw970tawHhzCKz/ar5f22Om5iUHbnqIV4B25MsXMnyQSycBdricS2k7Egu
BjEFnnvkKwJYMnEgQ2ujYlSNyDFxpcXInp/PS0HPCf+D6WTS2nuPcLdp+gRlAY+c1AoUO8rc9vie
G0M9MXuABWIhx9pXbAwyN9ofYrmRtmZNyUMVOaPSmNJ4+19le9Kovy1YieMQDL1AL6x5rQ9cXbYX
5QwAQU0jWy00xyxpbwb53uWphwdCt1p3k86AEEP1fi42rD6J89s3t+wY72CQ++JXnbNv7O17B02/
5RLd6ZvXnN+FZiR9BLQ1lErzX6P5k+696P/3gfradLKcmg+dwhY/EG8cgC6gNpMBR/gi8Q25bM7z
98D8Mu3mDQFs3LC9IK6ebKCsHBT9/ezzO0tqH7NCJr2/wBQKl6aeHPpWD4/HmLAQNdUTiydKVZbb
BqPr3ndggENayPX0QASQUulv5w25avus72SzfCIZG44hL0B41UK+LRXZd0oDzdKERwYRgJJlfBYQ
VYrEa1FjUvjAUORzjl2XnziHTOmQyQJOfLsyWQ0YEgCtE8x9q8l8nDmhS1wz1Qdg+5Ul1Zdnyp42
y16elpLA36GLcQ520UzGqGbBV7XIHFtbEYpzdZRM6eECwzp40zlkMlug7iQxR9wAs+o/HYNkdy2J
FEaY+VcmxxuDD/m3WvXdHMvAEiTe4fHyPltGZzVlxofsaUF7yFVmuYJFz8QjE9zzpi5jzbwv8HLh
B+JdWHfjoeVeod8U4nRy2BAyFXaDL9D0vDdZGazzxF9L9Ve1CR3kFIN0TONwzccWWzikYeGGxK1H
ot1tVrtKrqA3HJ1VVOp/F8wAYLuyp5LNWBrEMYqhXbnk+5/ZXwNov/b/65VhgerqmtwV+EUe1hI3
K7syo+E/1jOtTykJ/DCF/3lMy6n+BiCUDWxrlpQSOqHkQeK427YvXDc/CE79PCplvOnY9dSpGPUd
BVskIp4l8R66Fh4YRK/TNMxfMf+INw8oTHlV6FDEA7CkNb7WO6vBhbcbZRxT24/LozcyI96tL+CY
PBmrqj8xQKHhmHSEsWoieva5XCpruzPsymcibUewk5HAfmz0eFwD5L88H2qoZgBuAn5QTGIgI7FW
ZzSxilm5qSH1Oi0c6fD67DTLq4e89OVTaJSsAIll6IX2MTdxky4qMSnlJmUHTYFRRWcW3wtL/4S5
QTkRjixWVw34lQl3j26uPOHYG8gVm0neA1PpwBv1PyT8nbxFyP9pFrIN/gRfXtH3XKdB1N54phuV
mtdJul/sZLiCfPcDZ0UIQ90ooFC5elTOJXEoem+86Nx8bjR0Vgq1xjvPbv6mD3wM2VmdUDImdrWW
BMHHOjigAtDMvdcb12UsozFblngvrtLawWu7/rxEOy9yNGTRDxQImoEMSyNvNyW1lIOyccp7Ey1O
IN8jYIXeJDCGac4Q2UWyOJKmyzJTprk+ksd5Kt94CwA7gClEKT0CG6drybMg36ewfUTLO9HYphqu
fSU5hGqhCdTvqvbmg889ir1Wu4gjkXzA0QAZjQvRvcrCN8oGnx8DNWa74cWpUcnWPZ0vF96TCf9w
fusAV1tjVDEAFSFmxlHo01VD7wstuT5AIjqVTRLz2y0co2JhFqSmxxWWpnJux+4IKJ8wNWwhXpUu
YQJybDuRrk3uVlqkWtOtQcOSt+f4uzeu4zsAu5q+m4jFRLx5BUvr5sqOmVh5uSDiF5OM6KtjBCvn
EmxKSBiLlyoZvDZn/It3GCtFw6eMMpH2v+3hm15pt3GwhxoAN2doqCMLLfs2FMQM4/whdUTaVdJP
ma5XOArqWEtxSbYdLpjCq1ibPKLwbUdo7Z9ZNbDESvsaBegpjOjwU1q+aj3HhrYW/47R8rShWOj+
XU/zK1f69BioaQnhkrbIOG1SiyjHiHx+HpWXSXSgXdWrEkEDmN2qLcb8We1Uh7xJE6oFHUf1hxqQ
6FpDVnW9y7LrQPzIffmMNL+KJBYBseUUPea18Fk8XfHArLoeWa0DDgINl9Ah2YGE/d1RpEps6tb9
hFAg0Ejl2o7gRXmm4C6PCClqP54eMvi4S2T4V2010+XHu8o+uodCjh3hMIyUwoyf/csRr7u8kHLY
Z23WzPAVADKge9ktaG84xyXr8U3d7v5zDW8mf+JnHU6i4eoDiJwfqVV1kAHr/FSR4VyLs+8DA6aj
dRlsrU7unQqGuZUw6KZDCJqxqGCEhk3MwjAb8ntcr56216u3LPYnh+mIajuPdRUtOL0EWYJtek1e
ZTKrg8dNcdyqq4DGFcse4YlbNe6qqfBb+/3dU1xpxMTVECRiI5zNfCzVMitneUGHYbWnVVFwK+cE
2A9cWcu8KHa2HyW6Ju1aTtRQ2loxK+jOkF2G49d7/wa+xcftjy08lGw5NoMAIqIaBJ2w5SVp5cJC
xiZIwVL5SR+js/hw2xDleEoo4wliy80bUlQq99EfMuil6hVRM2NsDtAJeCGtvvkkzL/4dEpmYBHQ
w3t4dv19iOIUmYtvRi5ki36X+Z5eIH374bNEeS6LAhSr5+JXc1gCZK1PYPz5P2cLo0ZPO5ByqJIq
SYv4f0dpbApKs6pLX2LNGablvE0YK2YiwkfPdKM2bTd5sWac5tA+Xw+2OG73rqsZGZFTpewZ48AW
gNKDcgGgDgu6SWRSjkz9op2HYzY+F6fg0HHm2omkTTKkiyBlLBsn9RElJXK4gBDVNeuNEsTOzXV7
mKi8fqCPj4WGRqzcDhsfYL9IBALxx3DtMchQLj7xHIJZlNP6X8HiG5PU2fSrsksOjP0kdXFt9eqe
W7u/H/MJ28+QGIYdf151ZRRbV33yNi+oU4Kef2c2M0Mixfq3RhfDkCc7PqI0PJ6i9fOo7MFisJJe
zTH43WRCWA778zxhRWFXzdd4NCh5KWzQhp7Ch5A1XY1on9CHDiLToU9pVd7phhdC3OD+62mSR2px
j1dHY6v35kHzE3/i4+WUJAxDZwqHonuWW58fgiqCpC2Y5a8+4sIDR9BktvLgYF1AVy6FdibFDlLw
sPstT5SkKBTZAyHqwIL/stDYuJB2qsQMfJgeyMm+8P6INxD4a5rvm3qHqEtOniNU/r9lrNc7edxX
3bBmBSdoRMdnKKUBBj10hI2zF544sqGHIEKkxFO8uAwAqs+5jMavU3nL0vtjo9ce6kTz8H80pxSs
X9L2Q+rALiwQ97lsN02Jjfw7FZ7LNQKnwxeCt5kTsWD/q7OMZ333nrIz9eGIVQxP84xMEEj6Vs/z
yNlUzWOs1jtCFukV0xNbjtglgJ7dxGSyUH1Ch7vrugTS/f/d7dAAkBKVJnz2NQicTl0zVpkZ9xrv
Vw/KwCpRjsY32fY6b7j7RTq4qNT8/5sR0BKJ5JUaO3FLhv2x//QWUvGUBkD6OhY7cLqTaegW5KIt
7O//qeSF4x/6WvNiHwnYMgjlsVD6afQ97DGzYpi9Jf6UDu7LVfNM60ooigsELCh7jUv4e8NtNpvl
OpP/wm8JXC5mNXJzygHEGA9572BGSGHWehILxi61GPjZLjZQX9JNw7yquuf6t1DtFdNK/hSD1dR3
1hNC0Anna2ThBB/fVASOeOR7V7eT9BnlFKew+OthAsb2pEI+jB5OaXMZJzLCV4Xfm+8AdrNDBguY
E4iLVZ5R+9f0AgsJK7Q6K5SMSc5DAhsALO3mnDF7+j7GV4OlTrILPWbnVK02hAT0CEwGio2qD43k
GOugoO8etPUdQ4a3LXuQnRGqrnDLj4EbWaPjCzPkAb+IScBDGEyLETP58WaykwANYWgOL1PoWxca
E/5d4rMuF/D3tE2tF6x16qFnFXaR2IYTmeB/j4vISQ8QAio/sRG2MKAcVDVBcfW+1hxEmoZXOoIe
WuDtIa80fn/kjs88aEtJE7BHMDp1otmdfINfRfgvxF1Iob/IOQLlSSDVP6DE3RC/OAJBJYfBhiyA
PJrBfE10ksCZLkKjUDFTBi8xO5vv9sxbM3gFKQLEPePGLd1jqgeKaWs/BKRlrM81syAnUgsTPnFc
3qooQs0ODiFFu9V57CKmDbyIni5HFRFCz/0G3p8zbAEyHe+0Yg4LforHqSl9jerxRg5JqxBGkS1g
ESqgn7IEzMAlMAKPFVJcLI4DM3MTO/8VVhUqtYaRLlSamhjTBX71oApoxJmKQ7sLi7AEopXcUyH2
D3/tnAk6HtfBjXQ4LPT2+2oh/7n9huYM/sqiXZrtaZghPfDXURsIhqDPurpDgJAAQJ+SJZn8gykD
Px0mJZOznDIyrQruvM09j6f6HR9VNJX9M7wO6It59wfS5xbajkDQxVpaTlkmh5YPstad7KW4eBk7
pWKIcJJnGd4rOAlRY6qZmEpyGvAE90SCEM6jNfNp8/D0sxav5AAaEqI71Nc/OqfVtepS51+XiGuJ
9SqIAKOTZdDKSvnYtKMV907DpeitjduDrdnp6eykbQ6NjoLMuyYY7fRCFyyKGUvBYr4EeXFylBPs
cIi1+sNDD7GmzGqLGDUIGamtLoNfKJENSI580Pp9rVPsy9h9Y9GmRHcKbY8jLi1gQFiBMkuqZrOD
PwUUyoGK4TgEo+0On+PO7D46F2DivqWQ7/iP0eilaTHM5JV61rNHXd8XqmlhA/WjNbz4MON7Pbq3
aOHCBYCT9x0DqowqL5Y588++yCg93LJ3M1kWsvxjz2mUXI5vd5cMUROVgNkq5H+Kbx6N9ku+2YFN
s2kF0jnpN3oibWg9htYgcrtg7I3qXcRWjCFUSr4NzjHgEashknDeFKNQgAsy4bKsk39arweHl1l2
YFLhCF3veNDJK728QyheSAStxaZxpYn2tcG/FLGiSvy4ZMx9I5Hm5Qc95Z7bZaqLBOtCwBMlmXFm
ksZdwDhzWqhCSGf05T2JNW+V7JOlC6nUZEuoS3JIDPk8lqcXdoXfT1rR4Ri5TvmCV6mcUC0CTvoI
/U5IXRTki+YL6PPRo2R4vzXJ1h3vIMYfgSYWxUCeMhfYZSGgKw5MLQW1ALr7H3f44BD9IM3hP703
F+bYFokdmHKdRo7MSVMYPa/OAkICGS4QwibYryCnL9QZDnHNL50mALmbUofFzYIiZxZ/gZ2xTl7I
SVA2IPS0EYUcBSaKvYxZjVoZ7Cqsp2ECcGSdUJoN0ZAUraGJeAbwflqFSxAR/dXNWSJWcxcwJ1nt
ZtjkI5jCBnr4vCH9v9NoVjBxXP/OpHAYy4LPIb9+G966GXTP94yvzUqjyy6iT0Fg00lE6VNx9+D2
s/F2Tmxz+zc9Tu6K5JS13ODQn+bmC+WP7n58eUXIcc0V0HHo22THRaH6AnjBsjmtJRX3b4an/T5t
lfY41kY6EBEjs/6yvXk8hVa6G4HCxYH4ypx4+0chgwtP0EIIA0t3T/yuScQ8xxfHacnR+CQUGW2x
ef3CHAgkQ/RnJcRpICMc4xXry5kJnngUj+6El8d+xtm7pNs3KC78g4m3HnqdGXBd9a7uq30i932C
wD2/swscp3BEBqlICV+XfHP7QAzG7mtyXWZ8ZFaxq/E0WXtSaJeC/swD1dq/14Ppk5uWZeug9dj3
SZ39IwG26wF64KNTQQwy2t3vhAetC9j2/LyQaYBvjBdQa5zaiBY041ySIo6s/CVxerIFlX3otJbv
Lw6N6mMqZViBnVmzefCgHQLNHg6fsv04YKMFYUOdzWW/NNuBTKezfCCoLILWybs29MpE4MjsAt+4
s8yckepCTky01zfscGWsCkCBaFgqv2N3/0k1KQg5dNm3CZY38bLkaD8Ii1OVOkw4Ar0pqjzoNrf4
ax5nKg5F2bMtMPLX36tjc8VeHkgxwaEBgD56Y5DsUPMML/qEueMa5xgNmf1AZtR2hyTzVtSVo9vn
WJN7xBoNTCJte8Dc6XyFPUs16zQvtanAysr//15dhd2wT5SmNQrmfJBqsl4MuoSboMRAKKd8SZ3n
/O5N20E9cdWwKK49NMeVZnoSGNBvNiGwoXoQmMyoJA7joKMPE3BeKm3S5yPWrbY4+mn2emhYrvwr
VIOgz2Zo/bB1FAdORm1iVIo2fr9fsKL2vAdzdH07j6A4OXq6KLgYIkZ6CB1pRWR7QchahHnILlP/
UGfTWg86NVInNSqWG+kisfRL6Cziu7q3RmXooR+DXqARCu3dMP+M3ujxn4ZlL64m6pPnOQupE+hZ
JyY3n5J0DypvrG7yIKCK0VQbvHgucbjxYJTXWPDWJla/zdm6rQ4LkdHPW3QA3fognFHUPB4VTjFj
bJZzF4fKGv1OYTWq10+dWecfQm3X2adKWyOHzGI7hx/XJdRhvE9M4MMHSYw+CPJFlRbg0u/yq8Sv
MICzUuApMc27ydvaQB8p2IhFLTA3aA97vpK7Vdtz4YZbs8KsqI90z6sOqFiP6I8RtGBcG57Jb1OQ
jMd+TQLDVxIbfRYycN17HQ9WClmERf5h4q774h/TeM4mqy+R1UFmAHm0uWJVTTq1IhHPsFohf75x
KDWRHl3lDSbt6X9OfE0+ZKteSdhtzKAy4lr3BROq81nJjy9EFA1fb7KB0HILDl+EpO1CviA1Y8EY
5upl8hv2n7G9ksDcjralRCX34AADlVadhJ8rmSh9uPIcuqA2EiK1sNlQuPQuEtIGJwIeo/AYM6Gv
xzHt30AIhWMb3rBWRXKS7UD3XR5DMVhfKF25xO2oUIIWTvZkMNltVGhUWdB6wZHjw4SPWcgqmmOT
L7jzorhqWS4ywgzhy0PIiY+tg1t4q8ZSCNpOW/Rx2oPLEGFAdiCckuKg9h6ZswF5BtStTk+Hl2nE
35MIzD0KoziRRTQs8SUl2ugSC/NSA2JucFzzGwF2eFi1tJV7w33enyCd2MMdGappL1ujOMapg7iy
sEKiKmGS1hzySz7Zjyus9K43gjrq/W9d9huJOFuHGt04X7jaJwAasCebye1Nkcl3tR9GDJiLjWKr
RtbTcoTY/9u+MEEV3d9Q89NnjHASgX5pmxuB2GAPybAoZJMPsqOw+oJ/548zhqZ1ju8nfJbbkeNM
iCLCL+Fy1X6dqBvT2tpY3am/Wa/vmr2J4Mpu+8v1SvhQkQobaepxA4GrKL285rEyE9zNWJKY+5mz
7WPA6asva/PTnK6mVhrzNkhXl7FbWhOrDC0Cb9L/Mx9Qj6FGFPPkJxa9i1MF6cNcFMBHtmNMbbiU
qG28bHKRhfeV2WGTIBSIbvKZ3Ygo2RzUV0BJiFxKXwtA8FfrmxBsKNk2j2K8X8RqK7uANUcrbyM0
UgzbSDbY7OI1LZWMagP2jgMNCEM+zVrZanZ5Z7hdyDl5PazmRAF1r+Uzm8F1gMvPn1X6Cl4Buvt1
M5m9YAZewUMFDGPOgeSaVObxdluo5yddhUpCH5Yz5qfIY19HEMyE0esKTCMNgHeh3ZtGwYeqMJpc
x3oEZnJ6gETFYZKYR6W0Z/IX8ZlmhoAkPxdW2wLz0byA87vELPSWEJu2hMyaNAUCk02qFEPSS3S+
LNeT9JR8UIB/X6qme8Af0XySiRIomL/l7Rdhmu399E8i9bowycRHVp95ExQ1gLIM1CsCmzqqwOMy
01lWVxCkDMqOp6uEc//00lNnauLqnLArm+5FN0MgModu0l0xAl60xgmD8UiedryY9drUYWMKT7/e
Scqn4RL1tqCozEXdJg8N3acfDJHXTKCv3dIxuyT8Ao9Nt8bMAJGWGzcxDALumCCXxB3l4jmFiHJ/
lfpOS5f0p5QW0p+voAzdswRHMKjXvC9/PEqaR9Ncei0CKECubQbOVsPbyY49vghdJBxOpjefvyU0
X4BuFbA7+pCK0H5P4bWxcMe1+I6KMBhfmfCfRfuuckqkeHtskNpeS9YOWQ9n30yvWMSUWS8YlCtS
5+1r2z9CHnsWNR1oV+R+Jshe24B5fIibS46Tf+oz2fLRaCreHuMEyb/5KyP2Zfl6/30vM2sxC2sj
j4flDzcip/NVNz8JrQQAsgjYJFziELXcjL3pWXe3h+6uks77tDedSPnZ6LzsRw5ZQJrmB18fBt+L
ys+qL4fjvyBBiLdIvG/Yo3O2pJofZlJI9Ky7jCBe/5MFjCbk5MHuVY5JALw1IkNhe87VnOTg+Xxw
a4cq6kvbbA3ob17wBhWxqEainEnIppBT+jdgEoFJkHD7WKuAL7TQTYV6czh5zuuHo3XWmDkogF6p
SbGBZPkR1Ja+i9LBRKN5k+kuIo9pA+g6YoQvBmGkALfuT0EoTctV2lZrIjqNLUM7CjRmzFdca6nU
86RZ9uHYeJsPu7SrgkNns0GRcuWZ0E6nZeYkq6ZkkfC4P++2ks4sUgfMnTldSCsGTqC3WRDQyBy1
wg+RNQxTgIuAtNyt5uEzChwoEAAOvVRLPm2fZU5W0MIhDg5jgU3sAOWsFq4vihJeC+rKl4JRWw6R
yq4XYlHT/pkeSP+5DT8Sa7N+3v6DiJnhWJytt2F44ni7KBiUBbVFyH+Ri99jynQ38Wl/2txCbNOU
tGykpXqkKsCutoagMSjiQd+zYYJEHbD36HzDQxfc6dRLmvySTVXYY5jfmPssp8w/Q/VdyliNkuI7
tpPQC8OmMV/4EpXiDcmJmUz+urrqeHdyKcOXa9UZQK4qU+Esq8Q1iHPnbuC/8o+GOeUt7Bv+Ig2Z
wjxEVEDDaSxkxD1OBaqsL1jLM3idnVvrlLJvaQ9WXD8jz9trRagBGemOQe7B2QcIWJJpLp7F3b9a
94pLldzM/nBYmwjXeRLZ85O9JWoty+ZnAiTYTNSkakvimDqhFSyJWZANBfhe4/tsnwaSvX46SGKJ
RQ5qu39Genc0XsyVY8H8g2fyg+YZ6rH/szloQPpWVAeXe6V5R7xQK2UfRODaTJPInV918YyoPnCo
NdK/h5yqS4yLbI8PQtLA7TWJ3/Vf0Gt+obdyoqMeurroNWlThj+PnYM9DDIrc1w5nWVekYMO0Wla
d7zZLTp86sVrjppy6VwsIqaLWDLVz8HWIVNv16cWVzb4Cx9IybWHswR7dO1So+D6aSS5LvK3sAkW
I44XQa94zCLXktY+bLHwFtQW86gkFjbEnSJrDFHa0ZtawojWHcLeqhbcu8waaG6jrScyY8COdKkM
tl8Rf4agyoODQAHJHqNlQkxubQc3qeGcShyu+lTZSfEbV1auueqKLHwT83bwdLOzhA5Bj+Ps91cq
zcqE/UBkHYZ13An/fQS0V7/bMLvTWyUHNV9k2SHL3EYKZRh0IsDk3cETMKu/MExdq8Ut4bxczS31
GbHZuKn5yCNacuClH6aZ5VEyEcIHWDLwR3fiidVdOoatTQoad3SPf4/c/ajcElw5AnlYUyhR5MgK
R60SvcTgKmc0THJMKsXs+EGjtYdBtxWkyh/yhBXIUtPbeTvplzc5XH/P53nmXl7eK3p00eZmiDgX
SQOWA+V6K7AIPR9dT0q2f3NNBBa260CCev7XNx1UjV6p6o4rSIXoRW4kTZPHaAf+rCdUZzgANgyH
xRYmJNBtSU8mVyNffEQtRRbcUMTnGk8qd1gJRy3+xlFaBrxLL+ZRJY0MY1WURPEpiOWMkJVZxuWj
LWlh6yGDeerxF36JDlWIEoAVjW7wfuFo6yPZV8NcW3aYvvwXJgzFJ93WyRDxufpoTfJnR2P51uDO
Z3m3EbWK22cF7xwKnJ1IIZJcIQsvhfb8E0QwDiNXZ4V7AD1xY0kL8gmDO2KPxXY/4j3r4ES6HTG3
vrFM2Er3VYXak1yz4hpjK+/J0/3hOoonL8Vj2/eq3vqIq4En3EjkNNyvIXdy0B8lxPd+GQIEVx38
TdcqekZbdAcFD+Nk1cBPSRO7yJj4nOHYdZag9T8YcLRrBlmlYc1IZTVEQwl9iHJhWzfflw7pxnal
upZ6C9eU+l6/1ay34HRmm5Ruih4mwnJJ295j5JE3m839/e/tY//zTIP7EWD75T8wdfF0GUXvP8wP
fDZrimpur/dz3nFkwgOCoSRE0E56UrHnrAsHE1wEfGdX31NdL54IAZZTnmPqLsb+x58InOa+RpnU
EImRj1ysjSSqQYOsgOCX963xo4je+NefJKFc7aRQUXb0HDDk1PgMQq2hlofrhPTPfI+wsrAR2jY9
54H1MOlVW4kIcaJCCHMOXLYl1UosBnDVTt39mgXEqnnUU3/yGzwPBGYTQRccqa80ncWc+vBZ4jtV
GZxC6ZPvuZ2QkkO862mUDNUOPosqqb//4QJLDw9iOBEYd7zWYMiNyhuaT7Z4tjkx3nrIcWkFqbBF
0JCDzJlTQHoM9E2JByFQ7SKOZOZSHP7cbiEQKokuWu4oUD4d1eLjpz1pHG13ABq2Z+zHeCuX/VVk
9dkV/VmquLUYOROqdG0RrCyUG1pqiQzPu7mnurGY1ApSMnUtZ0jTYkYTeG95x/QGE+OV0rmeFMQl
GBm+ib7KOGpsEoUV7m1Hvd9IqNEnZsav40GS/o+Eu8uCOhaqzJzQjcbXJBb3svPA4v0JcdAb28cR
ksYN62dtRToYK3//x6RNmV4BRxJYTuJ/G4RGiVdBLRXowXK2hK/fFGp1VDNeGL0SRxU0x1YuQ7Oz
s9kf63SVjv3T5G4Gvkfcm7bfeZYHSQp/Cbw6wiyWTR+TbZGBoPEaf6ZI36CYc4aSFUmiU08Oe/V2
8W3Xqn6G9VCUuiUM1iGKHo91HJhsjFqNVBfE08x4e51sLThzSVtMZkQGoZzPozdxNmnEjo+YfTWu
JHbZFqR1GabZ6wVm8JHBGABJBsTA4y1IuPKEuJOMuhon6TmyNDcVgNtiLzwimrYQL21nG7nZQHgo
Ey9mKTNZPSmut9po3ngcOYg0iVWgDLZIl04EjFg9jFtfsoMz9bxEz+obDwWZLcHNtpM3FwnWhTqi
BzoZ4RqB1ic6QnmAotMlL9M5IfWIJH/LZ/ct6UIuZ5nZm+vhAoPITyzf8Yanrtkux1n9G5lysgIP
AZbm7XgvppjH5++xw4o5ozvHfuZ+51k3KhYmpWTXmCY2M8LTE80gtlmQl5vPIBwWpqHHks1qdSB7
yyV9VcIrTERnbeo6v40bFFv39Oie6/5spMJcdbDToNudUhQto+5WADCblv3u/nWsN5JegKpwOkPe
YxOK6fX4ADAlpgjXBZq3QihQKTVMBtNIiqHug7bJc4bRPvCkLnlsktvNRRlhw3aM+RdcKGajq4jY
hXfpfT6eiCXdurp3eakIwqbMMxysrRMVVrssBK+CNBsuryyXie/e2i4Hq1kg+XThod2zbp5wtnfx
J/hvccXPcAw2mXPFxZwLwxEgenxCxGD2+RFn6RULG6ZRVn41g/ezWXe2oDukqWHz8UFIkJzNnIKH
DZFpVlCgBEW6tdbBP3pHKMkafLJ3Lh48NP1MzzEk8stGy/Ou3G8yFJaki9lwQjxCbOEeIH2xTNzy
5ICK4aXlVaOTWCisIG/RThezMoVcIf2t1ktF9IGu0NHANSf0kzRHYHAcfaD2bBuqDX0gBfKYysF3
qn6Wf3aOh84K2Ft9gT+u5bgOl74x5WxEtiZfErtIAqrynikMc/165xDg4X01j6m8UrbQb+yVl+zU
73iGMsf+oEev8he6/UotjUjlesqwIWd1TntpyN52xdUDCMiFtNLOIoLCm2aORpWIz4Huzaiy1wzL
vaD73cEvqWXHjZN+ztjbsharhy42BW02Js5x4dYFPg3ptoXW16+itw2k5VKqbFZ/oSi20Tsnouhs
c40c3i28xPiuWsTPkk0AtNMilPHcYkpIGHZK4t8/frwAULltJ0/W56z1WAWx5RIbtf0zNWlYGMvI
oH3cpOdInWrBdo9Pt2joYLGagZMzTsOYlBRuxxdq7CeW1TaHfXJAZpo5FC1p361wGaEhDkts/UZN
JzWhCTRJnE19jT53ofPo6jVFDLLRTj8i/ukcbz35W9AdB905Xb56qG7Si1TmSodTGFIGooOt5pey
jFqDQjCyYQsQFIAGd65SxREOW30GHmG30l1J/LDGuASLhRLPB2iwBXdJVA/diEKL2m2ecnMlr8vk
vEF9ZlJDUKt3PNWy30j7W7gh3C01TiP0UrIVnqWXkR0VzSF7GYhh0MjLp82ZJ6Sgt7lV0Ajj9XkO
dkgi2IurBSCuVpc3s9mZb8CrleLPWsHcwR/3PRTub9fDzomyZECDlFJJf9nkW56RK6n+hUZC0VGS
HUZqqFLanHl4CHCAJWTxoXBHMERXNBdT6xfbAVxcIbdVQ1VI1zat/Uad9qLPi5mho2vMEOrgJt4J
pEJW8WbIawZsMeiNMUCMzeOKxn9TlhkGHAxMQ9L1tARGjnuHic+T0yKbZZFRF7EFw/FhvIrIEWWj
qAkFSGBz2k6YVli1dBcbWiJgih3zFdbyhxE2uHp7oCOyTIAAcJSmf1hHWZW4b+awf2Q7CDB4A4wF
GshW+h+ysL2QYpKmFNsy8E8skelI4Npb/BwQmsYsEQkpz9WwkNHm52KvTmBjMyp2SDRy+/cP5a/J
XWn6bxisaWHx/0wFaWYY3T0uSHu1Jgr7UCjdvw1eGbZ/gaDZ3JEeNzrWpXUkaIWNixMpF9mEvo3f
DtPVzgBEgaY07ba3SYTJCgHcTNAUCGeeCpODgdcnv2mziaX8e63v/tOFWY6QQXg0MTYotqeT06Ds
Dg7VLUhoR5MVdBtBxuzZ427nvU78SpoBlWfDvs5qE35A4eH9ja5C+It5V5OldW4sFhu+fvTlCG+F
ceffYzvtqg4WLgChVWZaGBSnwEImAKQlUYJMjhD8Mbbj5wnTMgSVcExmZ9Z21Qu+lLtU5UTgSRlU
M0gATl+JwWs06uhMpvjCT/qN/BXa4NkRkeZfnMS3JqdVxYuejWTZcWDKv/2lechkR/JQOetyTJ0I
fX0IbD1knCpZrtxH8M1SkBSleXJNCSkfLa3EaKi1HrRN2FAkKdqGTwaWUe3VnFSwwGEn5pvbhrz7
W5ZDJLdcJhWAA2fF91TX1rj9tPsCJNFcJECQHhhWpZqceAdws2YZVHToI7G7W+cyc3FwHKP/OY8R
EXTZc6BUG5so+/oZf9+/msk6HO+wtZGcx9RcHieoQ5QkfZy6nnbV64uloEc6RSLHD8JgvHgTcgsN
yhVoA+WGVTqtjCkR8xvFeW6GKztnPycUgu0WpDUxyTE62u/CQS3PPWjHmNc8JWmYA3jjcsSlEl9V
1OMkej5f8XFx4EE6XinooYum8VVo5z9LFxaL950HDQLrB2vPH9r8Iq61En9BFx2v0IBePeNHSwQe
Oyb6WoVSjX1op0/B2GbV5EPVVAPieW/QqkSG2TLXmBvXBAAGRJC8CB+qiqopXPqdPuGaIJbps1R/
13h0FHxeDAtBdXAVqftZjjPZ5XwGz8E/RU2C1DAncU6n3JgHm4HarQwDkuPoSNDx0tbP0WRimGd/
Ay+XNjrReKPpssKIy98Q8chnQ7RAdfzfowJ0WDwiWdHGKcyuQgv/zkIIq6/l8Fv6hk1DRZ3CHYxG
MH5kkAc8ZtUGIObY96OgpHiuXSFLjyQVR6IW1QLswddRhTznFiR+MTSFfbfdEnBojNBnjn8Wi42l
XE6qjRhpLFD6rS3/NCJcWazercPmK7EXrVea0Zw1RQmxWu/9YZdo4Y0mq2467JjibfjXQeX7MUUO
IYbAHAJYn0xoD8YYub4zGW+BU3jprjOKSsgeqTfmJvDdOj6h4dYr3Y+/H/cUptUBBWloH9ei7Zny
nO55tPhX5GbW+XKrXb5PhyQ0PyDfnfYcW2s0+K62dU1vJxmO6VOXJKzCA73nfZ/ceT538ZdKMais
nR9Jymp5VoLeXgAz4WQMFiVhU9+OMvN++pQpOUuL1U5AXTBXfNRRVO8NNpCjwuYHdAqELmWPoNa7
a3Qiyl9ntpczMntUSC9CMXUXMlO4T7oEV8U2buw+taibbO+10yPspnc+aUyJCwy3x/FPrzzhY6G/
3b6/AyXBL9aGdf+zW4IxqXzxz6fdxtBeblWPpeNx1AD+yJqxQaIzNaXu48MuJLcq9g2HEIKfaeix
yOfE+dVBMBsBrmdMlr3NSN9mq8HeRhO7zu6Bsu6ttIaCiN7P/uOSCKDTHKNTl7u9ardjyPluVMtk
VgdzDGWj+xMVpMgBtjK11aEolMekFSq7JUo0zSiOp/P0ASF6urlP6jMdjh2vc6aitKk2ytrxP64j
jX5ikjx8E0m65Eh6RSzdSozl0kV/oMEwKqDkWXbENs2gpMvqwajY68qo6Cc7T+NC+hdk3wNEP3vr
Fj+EQs9IyYh4UtF6KupkXBrDuiAp1aoBudibFY2i7zUL1/DISp4fPMVCS6E/oKgu5wZD/N9Boh7z
WZbI8nfyrnAOniGjxKLsYq+GbjJMEdED0iDqvGOvshgrifn/UkO6qiJ0KRVErtc0aLyT3wVinyWo
eRRHsmLd2fYBDdwq/aYhANSQutwBNIexhTyX4e7ArG8Aa4aTNWXdnbsLI6mWT3z1bv9SDTtD5GAG
utVNgbHnYol2V8LzaUAwLrquaRijFQb7XXr6huJcBTthCh/ZlTB/2GmlQzwEWI/FTN97NEAfT7sf
8F7H0EB975orXxOS2XK5xCXIkT7bV8RDJMtfGDTZUskmcFZmWtqZsURRCNEO1Mepu3/QFA2XHJ6p
ndYUNDCXgHhBENgDpwpud7HplTuamym+cQZGcDGji5PRRdMWJaEMTqzbeAhMbgtNdvOofHhqlX7/
zPvKiej7tknLpUwYbCDrv9jOV7cS1g7jEbYVXNnUzFClHAQ3QU9Xg8NQePw786C6TqZC0EOXYDj3
6Nq3LKn2kVGmQwHX28/diOuyKVg7W/tqjxblPEc5yt88uGPMnJ9AjUH2Bfm4jN3wlDei1KRhFiTG
til1HOHKJnKEE73+3Ytl2G4bqPHixXSIBDWuF76KAXwND8pTbvDh+AOT9iw2faaSTxO3FzIGf5eN
fXaFCedqc14gskNldkSG6seen8CQ+4RPIkARBxrd5SpjNAs6JSsM5LRj7Zzs/wkDrfcpe17ads8n
jAt8khpk60Ayp0RRqFsUax1QLoAMJn1x95yZ4nb2idqr2wanTj+Vjrrova5gxZptA0mca/iSi0gl
hp3FmxlcI7oBZeAqi0UqCz0ToI2Qa9PhoNNlBiNrWbuAO5kC5EmO4SUPTUVs16qHZmF7D3okoMnw
B5l9z4upVr6rrt9nnw/kLKPNfB/dfeMkvZUImljQraV96CfPTQC36RiLx3yEF0+9RdwY4th5eFXb
NRo63gNNZkUVj1C8OmsC/fqyZNObYKiLZUQM112lRhWCnaW44Y5zUFXIxAcbQ6V3s2pEY3Cz/lxH
DsHztz9R7BtAOeNKnwSU8rgOMacts64FnR7qMDlunvgcGVa5KgYjF9Bei2nCl0nt/VmPqsrOyOhH
PqdphaDzSnbZQGW0osCOFL7gwTohxTSgTi/YrPn12th88taVHv9GpuiEKiWtSpq8513bKu0P2DJU
1poTxRj8TAWz2Cn/snk7rTg2ZO8F4AqTxpP1QtdqvD+F8+8KVCgOTNjl0K3Nt6kd4QgfzJE28MpO
z/br79JvDyKMgEqU974G9hrFGvY5D2kBLTLmkHophY1Hx9T/KgSBghw0S5ALRfCSBUdFnY830w7Z
Z+CJ9CaX4RG7Xmd9u289UPMs1XOjSQ6eesVoQQ4xNq8ewdDdC8SFmiuf2tMTqeDTWFwHCkrKGnii
qYB8blVhl15atHmBGf6y99RdVZufUXWuAnfqWAvenrLWw7axIPfqpBkXA84v8FS2ng3l4ucIReVN
qmOziuSaZ1eOVpRs6LjNYNnUJlI5+EapRA2aJ8OgPJWyVfKGbjT8/N6+uAAc/EQBR7QEh7nmEN/S
mz45hRzK1X6kcQTPK67TOJxKaBBGRMK20B947z7OaDy/oeBFDFF10B3rEgiQxtJha7k314HRSzUF
HB/hV4uIhvwXCGzeGIGY+jJwQVqqK8tS695rsECpLRyXwMuwOwNdB+iF10aK6ICPkE1kfXhzv4MC
gOZ3sIChakv3GIyrA10doIgusyi8bdmzQNwxWrMWwQR3awuzubastCQzMnPcV/3o/dkcZdptwQ4s
maYRHvExSMSyfdMqTNpLq8TEZhmwKs3gsh3O6M1Y6DmqFHukW1fPCk1vLHzUceh85Bk5Uj/8QpLQ
nScq/vH4SkqIPcQQ9ZAf6DgUnm747d5T6O5zGEYjIKPZesk1bSzIgN1ragXg7OmcCYmmhqTBVc/E
mGNABV3Ta15jc+VOiv9jc6m0s5RGCkY3YEdrMlCR9+vmxlTIeRm7xA0SJVotaDyoq50OdGnLOMph
9RVoxZpm2Tgmz6LHZQL0wbnJMx1RiWwSr11FxHPAvVTMe+Xhou0xIhqlBR/uIoHxWBD+0g6ZjXUU
TgqdnwlhsQ8rT9JzmUgRfSpEyT+8AxI38YNK0GQE5992bBKeMjN1hCmJzy7JKCCFceaUDK0f5Myz
uexsql+uSBTW4ntKvCV/xPQJt3XAaA+2x2Wy59/xaom+jhezN3Js3oJnSNJSeCAYJvncMULHR6sb
HZhV9ZC0FSu3vLzpUvqaCSZzNQrDC31Au+vlBAXYR3h8cZD/ej6e8kzZu5+5qgaANY5QkB+ohoE+
aBsPf5luSTt0TFB9yMQ+qTdXxtVs4EwqR6C6D3RIRe5rT4sBDFVA+RPNGFRvwZag3ZRzDebqrxbU
c4iWRmR/4dNmSXda61r6StzajOec+TKfbw6R7uEX9mc4l074lNtUEZSsi1VGMH3Eb38b8kvDMk6L
3k4cC8KYNo6r8qmAsxdd/Q2vkJX1WAjTk6sPVxizJUkLdioZ8uFUH+Grh9MhYNxK4zUq+JDryJFm
iBBeOA/PnsRpritgLHGu+9f1k9tGbmLTfulf1/rOwz7l+SK/TQciqeL29I/RwVK7Rh603Or6tL1n
Y74wkSWT8qajjRhR/HCZ9Ivp6FU1I6nStUCE2ddPZ5Mk0+n42DFpE/Kn/7D/q2QctAZOH0fjkf28
gm9KKFAAoXRfdehi+csgoRpfC57sjVpY2bM42Dk0p5Mmu1Z/ToE7TX+QsJa6dERBNGlTQztxrdPr
ArW8JQg1pr4pOHGgkjTCGGz6+VFWD5pTGWnS2zftkYcjNm8AWoAMZS8J2MO8hHhwrcVCQP+zWh2H
P98zOGEkOJ3sZmNKY2fkEDEU2OIr375r+/459/aCTFk1gPEdvp6NqxODxg70L9BQF8v2tZwnvO3G
yDVGpXVmFnsU3Hd90ZWZcsYJM5SBQwpL5U7Cf8ZtzsV6Fqo9Onl4/hwKR5+K1t7+/zWuSzhLc/y2
+h/5va9UjuQRC781I36Q5PDA2++IaZKPlGaz8NnyJ9eUqvVt1TUBUL6A8JfNyxTSJ/bfEF8/4SBR
gLsmR7cNwBd4YMUTP+30QcqGssu+N2K94LtZeJ8trJmRvf57P+3HyPa8rXhTRjm+Gt0v6pwuMPCE
ojJTHbWgyj1f3n/j6hYZ1LzaFij0rVaU+gGDE/XKOTyQBxULWhwHJh7XLEVGkQhMiAPqyd48YY9+
W7rJW7D6f6MmhKCZKaYZKQiO1vWCKTlkWbWKADltc/W15sJgIQQsCy3p6LH989agH3HeeBmucYuw
ZsIb3IsLHPqzbhkbo81hbQeNwLN9+oP/6e9LqWR5wsH3JZBf6v3bhXOMx2L0dF0mRDD3SgaAMYK/
VgUURtiOeKSHcZkHM5v4DFRBOSVFiSTXcf45AK1chSiC++2R0FAhu83VLWa9hoGeTvwA3x2ISolH
YinwOBDQTSXLmXxtTsZHE/WR2A4IkVqSQF4OUUca+A1qjnxLJGFmpNzE/5Kwh2iMATLxVEmTg+7L
CwZ6aCRq5t9ilsqIKm/Flu8EQsV5/FVj/LuvOkR62HkpCRTWAPvtK9TuR7ZdfzXP30lNU8DQ88nz
2isKcMbSp5UIxOAEh0QCK8UGzNWKUh1Qyg3cSyvd/kLc9It4e3RpWxD5SzEJFkbnDUkkkOt2zCUY
xTVo7hpiCXxsSgglzilBQzfNaifGT+8mJv9Ser6S3N1HPuyPzr1BCztw8TdFh6il5S4OJbboLgTG
i1eIyyJQJndBBlSX9VorwVI/+w0MqSLITrDg3A2GF2VjMPyrJREVCWC+zKleKxuJvs4gJPChYk+h
+xINut23WPTKIDtDnXByBvt8HDtE5LiXZ9g3zuN+vZm4ccmBXE8u1mL4hg2MpjhWbw7X3dSmQ3Ma
sH4Oi93rBNpBvHX/CAz1oTycmZhZZnObFO4PPFc15EQrHRZu0SIrOHuHduKwYaY24a9Fp+SviHfF
d7vtc+gsKuJ8SNrEMWrTPZfbHcN4uIQJRuaL64xDx70locPzCgy3iFAHGdFAlaieBSU0cJ6RIAql
ES/0eWrAW8++Nycrnlv5FTGp++AAnI0S8PxYrD4VaQ/PXqJ7paz30UD+FIhYRv7MiwNDNuqiv/ia
EhiLKkfxE8SYOuMmtH/DVoyfrmSz7zBtJ5inHzuI6maPFznAWqIGYTA2FVrapMQnILQvP2+HCECv
A1cRVmxT19QaN43aOOsoPXNHdlD02AlF5VGOdVZeevhkt4agEfiLZcd0GVZZ1R9xuvPEjyB/HdqV
LAOQhYzJZkoO3TeNCsOcG3YxUr4bm6tIgqd9Pt3EY+Sd62q4BnThKLt2FWfMXZdjwNc7UIZDh1sN
WMPx9UgLKpqG1IRQ9XCGd2o10MTCnQfYHOoN18obEIx6hcvj1OnsGEjPlNbFa/13m9dxGA5dqu2g
OrdRz/7TcdZq2YNXtVURBuPBRWV57QgtQ4EyAoCdn9qWflDn1J3662znw1xWG+iFbXW/Pcg3aB5J
5cQK0WfMcIrhrFS754nkeWFdlNduMg4DsGbmn6toxd6SIyWmD7YeFZnSRv566NGWk7/kyWtTGZhy
WDOa0nj1qf25bPxrlmvktd8FAsbTs5oLYkxHimrOk061H/nPnk4kG3qZIp030BJM60wEf3nITfza
XKSZRcKdnmsibfKgKo+CBQojMQvfpErQniR3Jwn605Ez29PlFJG+aeUaBXKxurs+7F/gZWBj37zf
5/rNQi7iKnxNkTHsNZBzGHlTNz0W4KPQg5daq3Wyniae18Ygy/lCUfv18oAYHtpy1S5vCjNgVBgm
+PPpz0K0IMgDnUXgarzHmIL0nhbs1io99y+LV0gPOcnjnTBzrr3m1FJW9sAN0JEvhLcbWjs8Dax/
YsKgfalnW6F3vLK0akLr6p9WbH9t044zVr9XfFigLrhxMF9+hQUlg9xh/iIVAflIqP4AYw/2uurz
2JywfHfoQC8S8AShdCQ8lKH/RdnpNr5IXsU/l/yeVzrE0UgXRrjd+IvtHzQiEK/RpHsZ8iQnrrn0
nUYqUz6XUItsi8eCGd9KJIl6BmzDXJMm9CNYDNJlA7annidHT9/q+Fwrcxv3gjrzjD3ZqJqPmX3R
YwahCvmtJ6DeTlQkbskhpRJGY0xPEDFm1jn9cDdUOVUMlR6mzerGzPPV7okzCgMhvRb5Fp6Uu8cF
qItl9hXWYmH7bi6/ud2nzyHiOSI3cB3p1IhoQuj5Z9zlb46VJxMnvqk6SMmrArfZemg81irlwsF9
7qyEgaweqZll9sSnwWrgb87H39/WiD0pl6wK2DrZbBQu5UuIauURkkTvxUlGWjcruGmQN7xAdGgW
nzaj7XWSLiEQ4eHiUO2C2yidNiDPH4k5nghBOKiF0+RScglyL67qz2JFzrPzB/nxR53dqGGEjSKC
n5WNYUE0FxJfrJFmzk2XFymKruZ2GHSDYIX7+8dkA+ftEMLdLwsKtMjJcF6IUBsV7VgaYFnoDZka
DjCQsFQ5Ied8oB3xPqdpwPShY/aHOZGQVure/ddr6jBmkY3WtDI69WYrBNQzVZtsfZdFq2H5MDjk
viD6e+hw1+aNeG3ZaaaoBWhdh98j7tyTJ8DbscGy2HIUvzAdC8XnNAXjK1RxbJ05J3E2PzODJpW+
VAy9Mym16lsWnII5tzoqjfw4zIR3zdf1hVoTg5vO5js6+NbImO2WNf0meN3+s4hv+8Ir23OJaHHo
S2efoMxI2eSTNVSe3d8Wi/FfxgCQoXnlFVCL7c9eEb5Y02bEr0K0q9RuI0RweRoDIH30e36OFiSA
MMw5lC9LqPjvRyPq8zTwTsxmjHkvi34BebUf6RxHJ7PfW9WG/P5JT/RRPhY/t3rEuRh8OpoXsMb5
3XrkQ2ODVn2YfNsv10D45ey0nOJPiM7pDoAb15N6n5teIKCkEk+Y2UlemRR1PQtIXnkvJ012Cn/y
+cr/AWZ4HA2AZ+ML74quu+aYkr15s+2Nn0drc4M/ZGOo8KEuRB0E7ucaw1TtdxTboKCX1AVGlPq8
ARzQ4g5644jDgLls1JhXfA8+/mojdbOkp9P5bNkd5tHo7T8b9cvvDZshXsPl/4LpVSiM6GACa3GC
zx6EIPXHj4ys0TiOMyLFqSYvf4mIstDNhYScu1xBokvZpT5WjU3jHiIgjUDR2wpKGiieh09vbTjD
jOKHN7fanyEJuQ+fwSv1lPlVkzz3V3BSIDIAwLyvEfEM1qzUvP90p+9AOPkaEQEf6DYNs2mSTJLd
TByWvvAfsPr2vk6hpb2sodRvjb3eoTp1Nqn5KbcjYBxmsk1Mukpqbq1rAnAtDlYbYv1BxjV3qrB3
IwVNMibt6f2Lq6N+R1FAFFNgtWSBHjN8mY16b1wc3QDjFKXbeybutJfQoRc1kA+vwm9pVHt8e26J
iGq3KkBz3zpP/d0huSEI0bfkHB3MynxqovA2DOzoB8AwyLvQSd2655UiOOQs8CXpNZFnd8O5hyOe
JPTgZOR0pyuuaikroQEf/Mx7rFhjtly9Cgy3H3w+NSIpVvDAkSNx9EtNvDEFPxLMQT9G1/6ybPxA
6BsFxSbj5rzu3dJKzTUEaSxQQUPBrD6ei46ZRPv05yyIHtXA35C6jtDKTeyB6VnQ4LyDsu+h94sM
PwNvZtDZd8NiY+D+J8ZLfNOfNlqWcK4G6qVtISPBXZYJBiJ8K8H7V6d4+5wtWP1JltV+a8jDNZwu
FLRkQDipmWrCGpKrNQLvOYThjmyfyS82NLjUAHuxB3D6lNhzRz7JCA89ffR9p4kf9p6nieYSEx2E
b4/kmEQ2xgpyFlYbwcE8Z7rCzomuBpvSPSAxjkzB/pOmZf8b7g3X6wFa0uD4w8tD6Q2h1zKokGfP
jzpiPQkMwYUOUwdzPVOE8ZinFtjoWvFU3OmTVUuTB4nrR0+mSFWmzpl9F3naqN/oG4nfWggdn5on
acQsMiJGTXmmoMW8mZ4FSTlGq5uopef8d3G0BzpcueZjrEptlTbMCHbdge9TE/0ULNos5eYeKTrH
7yGTfdWTXmO13c5d/m47lkwThSxn3bJozYNmKnwEBZaEmqiIVxSUBZkrJJF+mSdyLIskRsFez4bt
+oKlSU50mJshqCwSRZA4AH72NS6NLJCpNkoiEG49Dyr/PwlxVfGcl9/fzBrSDRszuslKKXNTiVEE
KRrfBqSHn18NV4BpMJ4l/dpFhIxtxs64Np6wkvhtyexjN4E1U1xNZC5HP4Uj7DoVWbS0vpm7t2Gv
DP5RsxQIOMFFmiA55nAfFe/NIhzdQkyM7Fhylyn7R6X+QzU0JwhDBsEL/AzHT6NBNb7hfimA1lbL
blrVazHsW//jQzOlp9kQGdRNYXpvxGRi9q0F1kSQDSvdRXp9a23En7AloUDAkpxA8SX3n0tKfa7A
rVFfsVw9/fitl4MCK7F6/NvHtkR3PNllZmwNXyWQdFtzSGDtQweKK4JTgbiuCOADANhd93p0Qpmo
3Syix+UwyrUPUpILM7JRkd2oA6ZIgf44jvwANPiu8NQG2dl+PxwMQeLYzoRXGMkaGPkVEBgZgCiH
8J7858aPXoCuzOpk1uxVSNeyAalWNeVY1sDFiE3PcSm2p+hVE0uPOl8lIl7vKVYjoui9rR5OY4Ub
zoCdxcA6L5cNKo+wDWp0nNwYPMevtB9y15yf5zVIaPiI8EnwXD3ZrDO6zTeQEqRe/VnVF1CLJ/kz
CrsCloQbKOomMbJPR4VvteLdwdraHrTRDFll65kcCL2/mSu6u43qpfbFiBNFXEKlAjuMA4lIBkur
h8+zHVG7YPK0SoyPoxTHQXi1D6MLYVptE8PTqB60cmA+Mwpym1t91sRA+q9WpqR7R9EAzIB5mH1q
BcbGJMVWrUWhdXpKSVIRCt+dVMegFsiBF3i99xat2RxMFMrgbc/KoDCtqbOylU41Beclw3ICXSft
MN8Of4RXFbPSAs3SWKQU0WqAa7r05StEc1Ws4wxZDCHDuKWYYlM2PeW6LduwnYqfkt/BBvJDqbfr
6Dflp2RoLqm07lHsYc6fLhJVqfhNjU1BY78QTbXUNgrwQVp0gcG0MJ6dlxgL91vm5ngc3R1SxHaB
y3vthmW5xRh6dnlI0I+PoOTs62AfkfjrWPcajnsdJWaOyEGpJVKC1iBD1PGip864xiLXruysXThg
u8jPWwQpmAZhmiN/KC8UWg/BKTp8MVz5OslCbZBKoVTRN58+K9Q/JtFQOccQ470Fl8RRCMp4O3Ul
Zph8g8n5Ua652oTH4ftUH+uKsM5Q+sZ8AMLSPgYEaG7/nvgJrSfjKdwypdaVcG34y2c1sZd5TQEV
N6tozvLIuXuuIVtNW1JziaSpRUsF3n66a8NouyUTkL95kpPLjprG4OlYmM+uB92kF8AQiOAnYdRb
wR/SJQcHOhL73xcg5xOigxbEo07gMYMNE4gCpRfu1dJflsxosBNTndha8qvrJ2kcWiaarzqxtR2q
YSH0fpuYJlYDfzHEdZ4ATT1rrEgAz7ikX/noxx7bOiH1r/s/AqEvali0EXlIZtxRtjQFek5gkpfY
h1eQhJu5os0xuhefsaVbqpurITDnmGLg2wMv/my5yo3Wpl/OJcJqK9WYLkcehFBUpEwyuhN9ibQw
ciULUr3WhRQxjGnmuSKIzcj2OrNnFxlldb51C+ANLgeh26J9KV1LbrQqbcEqjyWOukATwstvzVkD
xUBYw9u7mgHfHLoS0gMX0G4zjLO5kOu4pnOrbSKxIjVJ6CF8FAh6fDSUJ97j3M+lB4xdl4H+GYGs
yE7RwO/UGoNPOHtLIOMJ6XJNOVTQ83asc6iUcDCx2R8Y++dP+hPI+kFW8+lNoi3JoJ5fBx5Jm5E3
pbQIqaevgry5rPDRr12BSdX1bj4ySMFANQfrs7sfsYvcKmj/99xKompL82nll01XfNPphyr5rkbW
wcThEfdNDDnCBp8ieZLvmgrNabrV8Ckct3XgVsWeBjnSHdWE2r0KPud8owUSxyy2EQS513k48UJH
kthN5rThsBc9YYFMrKMIUHoFif68w4fQAQ9Scr5TP4b/jUsCMYUjyWxa7FOrBq7ozzBT47fqWz4G
mKzfWtca9JRD7L4HRf1JfWlCEvVGO9tAwoUSGvuCyOvHXl+wmsfvgLv+YhYuLcDYoHnlvaErsAOI
xnQLDZXXm2TyvGPpNyI+kXbrCwUkTpyX895LuGsVeCYPYVYCxG1ueC16wINyxhHWSHNJV5wlO9YN
fljrMojkmGevE9DMk3fLxNJVxewoiPsYyd6+94OUaBXG6d6605Dv6suKtjuNKft2WhmJXeAEUVVA
8P0UQF8oxprsgNghbAO8aHNAIlf78ug/Vc5ELg6OcXZ/fYWvcpuDnEkelTyV0bXIh7FRi0qZLAqe
cvu/xQcZP4KfFOZi1f/r1YwD4EIPK66safEY6IYY3SUWZju2hhO5I8mRBojCBlYBQqOOHcDmZk0A
TsUfrXu5UmOsTRT7tNxIO3Jd0VWun9AdFJENoxJNrlcRDrQAl6Y09t4QwfxP4Ljy5xxka2MV3zYC
b2I2Aw716+DPnRYWcBRiwMt15rwShXFl6/BTOWxUR5kiSHBfgJSTwViGxPf18+NhYxEwwu3F6WsD
9+0V6buRRIBT0/zgC5t7sdkRBP0MGnt7WL+55hFb7Sv7a+ZhAZFetJU+yHyKs3YPm59k2DEve28p
RLB83/3RoSTz8QWf7Ji/qKCNoT+kS3Ocz9V1/lnInMgGFyyjzPm9IQLSij19p9Syf/HOxW52SzDQ
2bVmaO3IarG4OqNcPhAldl+4USec1AIOllka4+CzhzKUsugPstNH/R8YT8XBh37VeIXV7w+1kIEL
+ANaHImBP4jbXfws3bocMEuAjy3T+XPDN9jnPQJlD7gCoo2NKy6woL07saJ9kZCBJ0BC1gVNlLlo
brl508WuXPBqcC3auts0jRyzq+ucvnR8ziiUcp7JBb/x50XesWDEXkLVtSUa75Z9BOgo0sTst9Oj
T942J1G+D4G86jicl7yPFPpRvC0zalMv650zOaeZUXQrCMdZGSc6o1xmon7DPZVk9eWxCuymLIU8
bjwfWCcQP62fYEkY+kisIbcKs3+GBXNWgIk6V4KXloMdkdGOkArV+FEU8J90sWozfNAHOoZafIEE
DG0YijJdFilIRcPaNJ1LpnatUJleQto63K+lGWeuj/qBY0/iexgeUCC/kagWTUfpMJNLQycS3vJD
quUuJY3FZoyvx/OeIczOTrFleUvX1A1JhIYbxeZFPPVNNVeGDRuctjhzIrkGQTHxUOuu0kpq3c25
WCB79AWIkLbRYwAYxsIdi4Ett9WHvyZn1qnyMLtN1dOKbuVz/M00t9aBbuXRz3NafGzrs3omqY8s
OT4QenU+Ng8id+2ajX+MCS2HFNC7/8gh1TDduPSWKYTGZ899R6PyM+GwTgNsj8sL3FU51k/B+urJ
KNO4XAVj8/3KGNC72Z9VPiUIbGolD75SZluGQz1Dq0yakwLJm/G/tA/TjOKXpmu4mvY0N2dohbtH
LPaTJPfL3UXkXNn0oi5DDWpdpbrwDjy8/LUY0tYvtlCTc9eshVTlq2ajQ8TwOSAkk8Wou4i1GR6z
xonsE+3cb6DDc/em9KQVtPQTKb/1f+bV/nRcpcSl4vsXeu5gtMGBh2+LQ4b14dbodKBNuw5lC5Pq
ZZ9jbMuQiW2aGhBtOESrkUedh5DqxdnB5CUMP8/692xz5/NjEZ0AAHwgRkpRHTjfuVzgyH/P9WOn
K7GoSEudm64KncYXO4fkGLK6AkXS4g7R/TuN89RNeS+IItfQv1ZQ0PhKO9XKvGllB1T2pNi/gkD8
l4ZnMsDpow6Ga9mMoWn0vNjSJ3XzGF6Qp/faGwEBICJMJyZo22/zS/vhN/c2tqNdupZXgOAqkKFx
GDyCBArQj+evxTvohYxDPdyFJaMVyJZEdd3UFxFns5KxpynSUpEqneJSkPtRJ3d83+Bt9CvfYJ34
rU2WboJeDFneRGk8skKQgBaXzFyp4TkeEDkQJRYWlDCs06Fxg03ihzppChvcbNuhbepcZR42FAd0
vDpVQaWHQvzoc/2N7rl1bRCrYrmPpxMydSis6aAHTqUMGRPhRrgB9W4Il3NHBYOkbvwRncgq7/eN
QbJfE+Lg92+HP+8aUFI9ta36BPzQbCKVEA8rk+L25vBkHO30PvozIJ9UowqFQigSWnYdT7/esGRY
EgnBzF2dRqABWdz5Xpt5LwnSTixLsqK8mEjt+aS74gOq6o5Rnd9rlQhtqq3KY5tcp2nffWyTDDW9
fYTs655/mh5XrTOO1Bhtf5luxgSt0IVcgbqRTn+WJHfTEoUbbP3227H/uJv40+ZopTHuQcwHq9Qf
6u2EQswDBHy1V0d14AYa89fuaX9RHLn2KktWJYQJEsz9IyTpjgD4s4hcaMim/FQYSAA1jLqZ7922
CYUk5cS8z5q4MoE6RgsiWPrMoOj/Agk4zneBEXo2FvoFEpxRhiKYTrsOOZWP98sB/GhzD4DwBrxt
779hC3YhdLstvPsHUxrtjm6pjN1inRYHmiMxiV/T5na5okk93zIGS+vd1Wvq+xk0uDu3ye0AG2XI
JgI5CyIFYgWDBA2xOdnP7lp2EMnGTV4kFdXu3kHS0xmUxg4wIzwCmkYO4s8g3ZVXHsUFuLYWEs8M
e9U88nlr6LjA2AxqlyD85uasNXTf4sAOsLm9/gyrdTFX/dY5VGeG1H4hZA1J/B4NDCKd9rU0zSLo
KPsWG4WMk9RzFynI427kshrxyt6z4tMIn01yo9n07X9I88gTSrbkNdq86XPmEAvymlntlgN1FTC2
GZJ80gtX41xVL2LtyHWcpIC8jJzIoJ40kwLf7W5aXrtcn3MGR0ZQoh1Eg3fZSZqCnV8udo6ivqOj
uJ4v9aRpODQjwP3tASEQ3FRum+a+e4HFA1DkSkh2aBEHqFWx7mqE8sx5BzZtJGKzuhxwk1V6+T6G
IJlZ8Am6JvcH5hF4jNMRHfmrZGnv05QlxSrjK4h8jl+2PBX+zZxohbFGysTJrSRvBNq2XnDPNkyr
8PZvWyW5rjUg3Rgpb/jse3MyV4zB5JbrcXKOUxmRiAG9LPp46nosF0IOTmFC15Khbw99H0QDAUDT
eUU6KzlnUlYIM+agVMpRDrtlceO9ZKz8wVyIxD6KkHeJ3gaDkoww2BEWGsg1WL+Xd9xTSaetqgM9
vJmMITo7zVEMiKMtMbf9p5gvqE0hRTU8elwcuFBx0niDEUhlq3sJIHQcTK2DTqZE0sPjQR0BBbC2
H3ZOlx458xwp0fh8lDX+9Z7P6Hz5GzXD3/So4Qeddc0fO+sgobh416pBQyPr/IbAOBEloPAAmgFv
7ng5z8IOtpOFFl9jer0L5IozNfHZNxfCwe5m0kzhkEvbxF7mYBw5aBQTKcmNh7fHt3NRDH+zdsjg
4iHWpc4zQbeX8dvsahyVf4lELP99BtRGBBWyPkCU35tsgx+uASeuo+d40gdF4BKZb9+Aaj3wzVop
Tn2KFAhmgv3wr16b83I+jjspuw3wKT6XtDxGHI9Boul4iunZ+yVeVQrQPKAAKOxtJPN7OG6eGZR1
DsTTtPImo2HcdU7x8liGZBSEfCD2r2b/RQV36MdiL1kvOTkm22a3O0qzfyOpUVNaZ8tPZ4B8nb5O
CHFaJSTlYVPguJdgqjUcWAxuzbU5LUT0iCU828ng+rVWOGZQPor5B/bUOnRqoYaXNaDEVYYP7m7F
3DkIU/0eCjT48UxVwsogmvxNOvz+oP5JFuILSlYO4fIrCYnWbtvgxHpNvpcZ6NVJp+t0+Y9z9ooD
Xa06+GM9qBOwZnnWR7iKWNxKvPtXxwNlWuwdRMQN5kpybbKFiXmm0c6/7uFrZU2ZY07858VmIhB2
EcD9+yK2o/aZstd+Ms4dCIimuYG0QmkbBiWoZP8hGYMDQy2yB+LjQihKDmFCnmvzZQv94v7/XXXV
wXG/te1ndcG3eliCWq3qrg49Lyh6dJxHk5sVcgmEkopRSNpWy3ZVxif8MzYMLA8VrNWOxXgDfSXC
Xppl3NPx7DbX3AghgiFkibkvm/ovSGBC7X8ySumZm0fxu+SY986O1l+H4+SQ2945BY+F6kfBOnzH
hvZbNgL0iE60X1f0e9GXyQDa3AmWTnGerxj+1Y9k5ANPtWs/OOonYmcPqTRGY0rwe0sAYmHyOUOC
79b30MlOXusiX7+z539X0wscJeet5Hk2WsV0iJBjAup2RiQQP89ZN0wUzlGZxEOT+9ZsfK/2AHQK
OhcsCaFOT9TRciSGyQUHUoTgHt/GOaxwawcYhyJPLl6OPZQzTj2xBvBIEqy37Q2TTePB6QGqhWPW
xuk8hYChcdcNe+6Q8zUUGjIhRntU1ZHm7aQGmx9xgYfh6PZiBSnbOE01mKIqKxb6UdVsWDNQdiBW
tE4dr1IGwCv0knhv2gXgpm5sj4nSariha0ynMpabuuwejyLfY5RawAS2ZZD2S8qYIGnh4nxG+23R
BmaM85LL6eoQRG5tR5sK99Z3cKJMZOfM9EifFlE6lbnIzQVMScSgwOCo+2Uk8oSZWYCSFNVhSLuR
Y/sNVv7lHnZ1qHXQbdM4ZCNThR62QUkOPVOJ7sJl6AHkvq1YKZOtCYN5Wm6QFuxPjoy7lEk9TZ6/
rclW4VBBiumMfNSOTBeoJbYbkh+k79hbRztzlh8SJ+0EQsraEI2s9J8I/cRJlVjkWG1nlt79ory8
qnYzUr/HZB2bQWgBW9oqgX9RAz3H/IQj0hXop1yDmcekQ+KG2ggGNZCAB3kzbCs6R/io0cb1cH1V
AifUUZEl7jfRMkIaYEgnzxxZ+fZTJ79pn3H5FNd1ArkGLBhk0UcOdnKTPOa3y5X23TFkSNAZDdj9
BqEv2tuS0hVgapMtr+fZwt64WhvGwesWIwy/4cN7UtcNZjWdn6H3k/ZGEnDLo9zRvZDR4wRxnanp
vX44CDs5lmp62Bm6g83OaiYSxAbJNXn162GXoSAYZHooA7KSEPEwS+E5He2nIfAGmb871i8g6Xzw
5+C6p7sJs7+T9rMYSK/GAwN9ArE3hx9MvbLykQf/MiToRTQc/6dcHCD1T6lqLmlbvr5fYX+mBhIq
y0Ou1cPD+uX5TU/975m+zUMvMAkBd7DMS+qeTat/UkMk2vVeXV4M8a+i4iMAeJUBAoR8ipEAailK
ffjcZ9eTtoELNjnwRL7hkeQZuUzKAtgDm4qB8MI38J6qVVqAZ/OOhj6Kn2ZHyMWQEgHi23RdEJHt
1EBSDdDRaextZmhdKwuNBmBYSTask9vRpFvg2LgyB4Q7M02T/HqV4vJNhZ3mZuK61WXnSl5P3xMM
7NWPAdSbscO/OQxRYOxRz1TA5ggeTfnzjkM3AFR131qXoyoWdxyrmZ7777f65YESOuxFx5DvTDum
CHmtq3JGzHxEu22qO6wGMXMAPerJwUUqbs3lglQl3xB3ZWJaF04iNj2yzB6IFco+3WuO4tkug/jk
KejPb0CN50BebT2u98wNYVa5TnkAnYYJbHKGV6lOZ1ujqk8bhngtrobiPmw7kFSJd/XzooPDgkUt
7aXyKFCmbiFiQpcIbH32z9qqlypNTvbPVLFbEvGoFYzhCyjKgZzumeP4B+rGDPLi/ZxsShEXWiSC
fVOLLtyWj9Pwx0NqSQgKZOwcipfYKMeCuihhqEkgN6cyei/B+DzQYkA/1I+FuUuKOB3kJrpah1dn
OkS/64Anw5t52xyw/blr9bS13PABGk5wjqJv3VDGTeyaDMsmLu531bwAy+zkYjkTfHnepfrXg3N5
2DrqEwevEMuoQaWO+SgztCcEeiLdz4BZoPWX4dax4NE6PfC35Kq+AvMbbUO2y3JOV3/ZBdg3IEKw
1gkTWv+Bfsz5+OIpYEdTXip46RY4EZvhoBR64qNUN1RJNAxgIUqN6YGecj7kVe3QapPam2i0rmVU
q5Q7K+gmbxcrSc/usu//vEj+BUElFHWZeZ11YcgGLRDyU/0FteNNJRAQyjfeznP2/8mrusy9Fyab
pDx1YvHjNMkHYkzyUQAAZCgg5P3wkCDySphk76FuOR6+s9hw32ysw1gENgO4iaQdXPwDn4R9I5hn
wYSc8Y23D2MaqKbCcvffv1732q2ywBGclgCwkobBUJHITQCjPIDAk+zoRvGgz965ZUZsqQC44JzM
Kebtx5FqFHo35xiTIWPouJX6Y2QkFU4GLYq/dZgrO5WS3juETnvlTQbllG+NQwfvYpAPBIaeqf3y
c9rCm0kP59H13z9vUz9IMHwqHg1qHuveS+LFniOZ0/xERAc4/3sVbk8bv+P/lh8oxzNFSsPSh0kZ
qZ7zsuHwkXV2+i6e52CT7EtCojBA/N8VGpSTc7S+ULmfuOwjVk7+gtxHYXq+O9Bo/lmVYz/D35ww
Xgh0E4Il5lN4TkTDvD2JUF2il9qzTcRLVUw6FGTQyiFs5gKn2VQG4Somib7HQGlbmlwWPBBq3J3d
u8x0IioAE8HgniGdasf93EIhmGJuhU1CQIQiRuDX1JRt0QFl95SHMRXU1F1UQn4SZURHgKqdzQT7
089pZ7aAPT0BPUkB1ED6JCZoTfU/IAUZa9T1l2b96xe/XaJq1IjA6rX8ymQjDUl2zNaqJo7teTRs
CRNNoH37xjEqfzDJ9627H6cC9jSKnUV3yD2DtWzR4Pzs/dY1ELAb4ZChC//KAyuLFbi3ayW8jkzY
chlLKPWgMLix0NaIO7YaBv0TtRB3tHXH5IVv8LEk/v07G15ky6nQfOJZ7eJd/utWt/6HzVDRiqWR
cJJfWFLNQkh5pI9K4RVaGMTEfn/k4PPfDA1cGnpMh3cvGaWNdBcZrtf3EsIJHocKmjzOo+fLcoxR
i3zbZ27Qi28LiTuyMpl6Le+XiUwa/CcAsfSsOqiGdg/FFyuFmMxyqbRdt0rEbuCP5614IJEUeyTx
nRbfzJjp4cSKdpK10I5fZo4eLFzTPRkj+1cfePqJHPfiMRgAww+SltuWK4rj+Q3prIO4jZqpnREi
Vyel76/DYKem5JOdyIDMtQpi72E/gluNT9818B3zzEISu9RC5swbQ3KJXDNOzNi3NMCuAtSVVPaY
rZmpBeqK+f76yfPoE2C0SM96H38G98Nwuq02o43BIB6bTZNuK1dg2Kjqxn/XifZfPBuXHsDJ/xlY
RRitNv23eW5+JtOl2ualI1tT2qrGjH85AwN01aAntQSA2zQG7I8MpoFOEgbmZQ6O5zHiiR2sSXwG
zqPQMnUQeEtIk5pA6SfvXDWFCTXxI6IbjiH0Ttv09SZHFvUj+jHwxBS1ImLRigkllXuiV4AZ3Gaq
bmmai69ukvXsO85DLjwDrGq2b6tXqLVQ7MGZWvGeankWY9mdqh05zyubWnyQ4aTSw2uIlfYvdnWV
2cihsUZQ0JOLTqJjbyJ/qeao+fU3hVxQExX4by0ysUcDOMhjKzMfuirEpCTzQseyBGBVFw2kmA8V
7hd5oAMYJ9kkHngiAL/QkkrCdiUklK0GFYGWGFIMPjUwlg+gjETM9x/RmHCq0rNoUlTg+o72SHHg
/Svgp2v22upPeF53+AET/zihbuvg2vnB6T7wv3cfwyriXEEfexdM4r1lsx0oP8MBJu5sg8yK1TnH
+VtvXLDtnAlaZzYUBDfBu8mL16jLcMA+o8/GbgxfaZf6oK+j8YjN54jv0R8HkKzMgwK4EOf8lYTY
YTfKklQWy6yUmU9WuPKa0RGJzV3Ze2R6sz3yD43ZL0dc6eS7b9BYsGKRJOBVkvtVCivskVOmeZ3/
/8kcIYG4TySDIeSaX1+YRDX2DfJ1/PiSa9MxReJBrGpN2g3cZXNDAJfSQw4JmuZJazgCmtZO+02g
kTf7P/KbCF3QjRO6Yqb87GRysunagP2jy5J65lRVKvoyXajzsVL3W7K6OiBkeDV3kH4w6smGDFuX
x1o9ibp7YoBWVPNpPW25W9NvBy/xGVDeQv/ZjtLJzDPUjIfhGLZmvCBKECVUxVEAKOkf2CEPKHeM
dSwvA6qN/PsU7c3DgI0M3IzwLvRcY2o5F0SUke3EluktSpBn7aSgNBJs+/AJctKFQdte8+yaRlKs
/1CW69Ayrcns8ERoOl+EPgd1hqvIM8DTEnzjvFGouICvgN1xCCEENFKjRpvBGL/0fEwk+EOHxVJa
k04+amr1yK6wK+bql+T9ASSm4pwK0UOvetSZabFIJ9M9XbHGMsmnuJ50my/JMcOiY548sb8Xn8yg
8yY/mO1c8mRZ4+9kVwo+hJPie6r6TooaGmzSkjrOtvOK2U37Y+HqsWtMUnihXgUlvy8wm6b1BP/P
MLcnD8G6wU4yklqXm/abQo0QDKzZYoWU/mPx509eIEQP0aD2px4m6J8aymbZdJZM7I0cLlkuxR1u
iBdbEhXuPdp/4bIqNsD4BHJ8qoAqdCBCrJRHzqG1SyjFtvYRZNQqHC96VGyGDfnPCYSJvgK4P3Ic
i19htCWgQBDqPmDfFkTfuhvgg22rjN56GOnDW5lQb9a8iPsWO9hq9FVWpwXuOwAI4gi+L9C3QJyu
pmtOku7YSeqTrfLsI8S193x5eqylZx9+l/D2pgI28HkDZ2U06caIQ4OGbRuZECWEmdXud65ZQ0SN
nF2yQPqG7oxbgV/7fOMrKlwi4t6tHRE9qPZBtA/djPm4vh6/LxiG+a/e5nsSA+hB82T0dKANZBCs
bLOOoaWtTHSI72mmvPpyizu15EGUn0pPvhR3RkIjXsueGrEuJLq1zf0G4hAcRbXq+QGOWHQO0+k7
FXfTLi1rPFUmbi7etyCyypr/CM/tRKtPUoxTPfNQErmMN8k5Ag4+cKz0m2MceKYosVIFa81yNIjq
C0GCOx/Fp2yCcoUkeHwByxbZ2IPpIiUecY92WLlsRw5bXJg9fPAdd8ViAapjqA1Uf8jtCwfARfYT
MJoAayCixtfDQ7IQSyQpQCbNo23oJzGtSNV4yX6H/UolLXNCXxi5lfu958SEUBT5JAg+2bAfcEvx
YhRCjd9H9HvjtK0H5av7CVmVVLV442xOSlOdVR2gTg59NsahnfECAK0uS5/p8H26ZPCbqfPrWGaT
15Uyyck1fBvAJ1JWXuv9RZba3q94Esmku9s+azZHlH3E6XvoRNLE63XXx4/cvyaVQpLizka8FphK
g2d0eEG8B6fNSYuI7MBbLACHtvADLh2jr9whCLydUj8LMp6wN+L6N418OR2/7eXBkxLdIILSETzN
xA35Ya/7pS4NdyjlVkO7lDKe1J917KyZE5qpaRAWXE75n2fH41BgMIOqXpPBg217PxjBeEvVZ0IF
kHk5JGmXO8hL0oD9R0oH6aTFU834dY3VjenGiVWVq/1MPTMnNuJUDJpzo1orPWzFS3HIui7pMMcA
+8WTHJqhQyvUdvaQNKLeHels0Nx8SK/j22VX/hllBkke67hj3zihbFHbgU2IEjJ2hL5yMxgq33ko
RfyDzSsz0Sh1uXxxfdXbPxn4mCyaegVI8yhIDAWaF2lSPQmKJQ7ZvQljfj7Q324h+oniiH4nWUUH
eNFRtc1cVq5cegOr85Z8a0TtYXAnYvJAVbLx6p7/qpKHtV2+gG23Cxn1Ndzuu/QL+YZOEYsb5dVi
5zGoqWESXBnalaEHfuBLo+Bhe7paRf9pxiCzkjIVq6iV192U0tWRuTG0Z5Pjt3SPFZ73VfrP2mw6
9DDhdIS3l8zqo0r5SP/FCbZvZxUXkOIrz/NKUcXhvWISeTXnCE2Mh2KZeqHe5OMaZ1a8kiuidERC
jVynQ1SMEVbw+6q5IkuVyvpPrklLoFqETlsMxXqM7UDVqYjbhYY0QSFbK2KAhiBcXjObxjWRxfjC
3e9uOzfT4XToJFmm+007XOLrJfBHH6rycIt1oPdtKaA4sBWgGBkNNi7weDleGwE2FUxrng9xyLpE
ey2s8UupGlcHyNUgR+BN6GowpqLzehWYp4FH39+NJMSsZXARb0aMnvpbXatMs7eym55iIOl0B/Y5
/6XN5fGIG54J4i06ndzqexhQWHAYhqK3tvz5AKAyLo4Z9jO8CWuat5hOiBR00bE6TH+5Q8xLG7QD
dKVVxNaIPP5HcrchZEgyYtByFDUWpvUxgtQt8W/yYIME3WgYXlMaWCGucl9A/HlygTz7PP3YLKGJ
vbNL3Nng84ZzMDiwVBEDVMPGdBBx6eWwCzYoeWzORfqYOKpVSmTOeYuxqhmlwc3czqnqYLISaEcw
OcBO5P91+IOKOpKBFtSfET4vexMzjrR72goPN8rzas6kMLzFeRNSB5kHMhDaBN57ujhMNnAi4AgF
kgG6ebr8nUuVYO/3mpAXGu4DXcInryKx6YyJng1Xip8kkQh8JVA0cv5P4DC52yLIWPTFlTGxK9ql
tK39JKcv0r8tww+uaaYmoLlmE92Fx6Xl8thN7WsFqRsoO3Rrqw6uPKvEZb4X0a1ScUrY2txzoVad
czmWRoer+xReGyzkGDC6i8wf+AKV95UMg+AoZlcPs8slFSK+BEKvw1x6ZeQIspOJ9FfZNm/FWh60
7zoDM4uALZev4aQqbIM8P1Cg5PCgDhrZo/JzrMEKPhsb9pdzu6FwaOLro9W/pu3c0ELRke8G53wD
MNV2ybHZgxfB7gULYK49jnOf+ZyRt9tety6czqzME0dNzhysWYRXO2I45+wnA27Xs9aCKomu9sNv
iEo35pqD0cKWd6vJo20o70WcO/Ffq7FWmuTJaUxOM47esatFQXJl4Nm8wudA8oHsb8aMKtwt1IeM
JLKvQaz4pt/bnUkY2hhaeUQvV9Nmqcb69pcG38MKDnoms7BHu8KmCCd8lUh9o8Qx1LefrEde87vp
2TpaiK0+Br+WMZuKi9yiXoEXylY+8W8I0Z1ZaMhirjz1ySGwXwVNiOa6KcCn0KPjHdxKbsWTbQ/Y
oVzzCF2Rh2JGaFLrXl/VuTI+z0F5M8jR7XnJKJsMl5HFTEZA8XedLtFUCF1bWQ9VuJKGvkznh9o/
6w4QGP7bZFvbCH2UjQdsfxQz50P0e2dKB1BZvWCMmKzVZ86L6sc4kAzSbi0qTdwRfNVMjXAeystI
AWYzWIdRP0i4aTLS/kEDRINkuolVCUzhX9w7rCFDXvebcu+C3satSQdz7pAI/Rlepy0ehdOjQfX9
Ny7rk34FwkQV57bFLDmjk3h9+9QLR+Kivmmd1/dzdH8JLlYHh90mRgFvOT0r/+FO2JMK+VP62kyf
/slJSBu1yuuRAPFTx6QstS7y0R5mnYcKTL+7grKtBRORDhDhYyWUvSTbHfEH34lrFsKEWsxtqDtg
kW4d4Zw7CVLtS56iTb9XAGU+6dW4P8uPjGR8in8H56B9ol05LPD7d2YI+2ZmRRFTvKSGXlS0b+ef
WNhKqljR4k2XSFRRz+gr7WCYBwwwo0ZyJRIPZsb5EU4ZFwGArfl8iYGi8p2YldVeBa8wqcFjDd6w
w3wLRep0bUM4HHLzxspcRl8gaxgeDQS1T3ZHzgKT3WoBT7wGdzlGLFhk3rWGUukZs0Z91DpVsj7w
XZoDZgckrSbKZ8rUoYcrzqzuvY8peYTSzlA1sFPfDit0MpeAmA0eLKvt8FEhdstOBEHqf8bcosqF
iI9BJ4FQNMpBb+SdOm/SM46/Tkbk4S2E2Dzg4QcPdbmd9D24tWM9Z5ENPUTOOa/p7GlwTV0dACTM
Vx8CjnAo5BRSqSj1l2rAfL4BOIDGWvDF2OKS7YKEe5Ut1HTvds3Ss0J8x0YoRhbtHzUi8HZCvSza
Ot+kmNg7Ix2/kzGcTETtfIVDhQkSOMquiRzwefe8iM7AAuojHIH3VRKy0lalf/JDR940+D6R9PV+
O0uVf2WKSPRTmJ14wxBZ0umn+tb39lMyQKhKo2Iok61qwXkwDRCBryjsKtxLNVj4BwY6Pwe0oIv5
jZy3xvYQAa+cHBXlvtn3+4nLGvJKhEdQXQoHkGTb1MmIea+b1gz3ikBEiZF0cHDwI+e+2exUMiFv
RkehshUoYWE4Dl+h31AzvJGFn5MCuYlHmDURgNAhJlIPlzg0KqJSX90SP3KDBFIKM5zIEPTzCGZw
qNIrVbbGjSQakLTBIPq0stZJx2d60zs58YeoizKvB36YFGTU148dgvMnF7t2NVb/Khf6OYKX4ol4
lFP0jda9hF6CE2FybbxrTdTI6QBK6MufyOKPz+TEhL64DSYtpO+NryVeuakkKyvu2+AymJx4sZYX
jZfb3DCNixuhfts6ZMuDsszGzxsXFjMaTC39YN6j67ozYdS3T7z8mWArOxM7qnolYOvnCXZ9IG94
03Km8IaSeDHwtBp6xKOFJcqpQqrCNVEHJ0OT4TIQsRQVAKUyZn9p1GqD/9VkynwlaqwCuOUNE3RO
Y+ZSZ5c2jVdlekFyUfA5UoRkOD/kpn1GFPJ+xgOTyZbHd0eX0sTJdrfbTlpMMsUkczuGqJaN81by
B3jN8X6T8OE9S+AavWrPnHa5aoGjgk58+rrmk5JJo0ByVYaG8mvSDj1XR61c9BJRlUvR8qcQVgyZ
Hn0nRPXbx9h03A5woFOTuBkcvXzmIv+MbLEjbM/LbZ3M/JPHtTG/aVL1EG0UwXqC3chYCOtfMdP+
hAKlVqkQBpStRAGgF8WEKqowuE6hPfsw8FPKrkMQ34gxlyI+sAnvCFsU4ewNBzOmjocNp0mPNAQ+
X/tYMktTerS7pHYfdRK+eGR2LHsO4/cFGv8JnYDctsTT0JdNcgjOPdkiJqaFfVZ7j7WsqapgN3e9
gcz1crRlVtT65ExzMg43NCKeD3M+X3k9t3KPlIinymTP0RDNnKiCAZALAqnkgGqmm4B/idsPi+bR
7imi699epWoWAkuTUE4kaH444M1n1sKPYh3tSult+ubXxCamqmCV0310V5h+f0vTqu++Arhc2C5I
3CRgOsILga/Zu8N8guzODYN/t/zoAznxqQkdpp8ZC5/DgKsMX5CdnY1dZ6vk8JZBhyS3R+D4T5nn
hh0QmqGfh6J8Lwc9MHyUALXlAcnIm/LVbDJ3bvzzLvKWCdhihGoVn5a/9r6UnyRgQrOu1Zez6AOk
vgS6fDZhu8ZmigTG8ZMf2k1Z5Dy5xae+eqpnpqZEZzidXO6XkssI/liEZSqzo1Iv8I5cy6cdZtbM
tNqAD1ps/nUyRVAI54LYVvT4wgVZjROIvCEQppCgLA3y+j5bvMtNE6q03busr6XoODLVql5tTjjT
zGP210U/J/I0M/CekSe1Dk+RSXJhd83Jf409cmPuxKFeEKKY3Q4vXJHhq3wZAQrWD3iVFoGNZOO5
mKs8qkJFilZcy5aNXb3r+AGj0sSrJZqIM6Wwyp3ZUAqh9QVT5Ep2gaFkHNOnrqdiFNSqyQto6axe
nGFqUEqPmQbnMwf67DihUoaq7oNaZywRpsD2M0uoTYG3a7Kq9OxlLOhNq0KppLt7SvG8iuOpLb5s
AFuteLMYKvua0IyuvoR2VsmsqG/G+CEHcSe4Am6hyOLgQdBo7B1mU3LFw4LHqWYEG54jQgfuGO5V
JxqtghE2Ouh/KDv43hRqkjDee1h21KJPWI7SFMlVHunofQ7HilJ6WRDKh7ZB3Ftk6wnD3wjKRCUh
GOO44MmYrQoX8RX7udg42HzootE/vjE/XnXryKpwwngOKTz+0L8cg9rV13GWH/jOxxRa1suMtIZ+
3WS/2BBW/MvmAS7EYgrFhOjDlr+GeCohKXVkHKRIZdN9RDPsb1thVwmbH6DWV62NZlVAN6lwmGLz
l6ViE9gLUBrSmHzObvHnVVKhsd1NKIIA53maToGVfJ+9CR5uZ4ScGCqRBWN2WPgkQ5nlpEVlwqvk
SPp9luC7pSi7KfopQv0+ZbhvoA/B0ZfbNuWH8VZOslvnW7YRd4ZTXc3z6F2Gi3c8MNVLJADOuEzT
QXvH5dEz89OODDN7HDyxgZjmvE/UxuJa0/DMUNezu4k+wjvib5Es6D67oQwjhPXuDBl8+hwBes+M
3XyIBF63EaHEM6gw05buuoLAYevkjUu8oRhzanrL0F+DtnLAN2/v/MReAE3/QaaWYcy0jI5yQ8b0
Kpdq/ifbjX0B7iATDqCON//miFjdMaqpkNGy8beStYrE9tb2AubQvrfV5wyVzHI9UQqeyrTY+kUi
3Lo7y75QoqZhlG14KkaNbAjRGn1K3ShjDPc3mW2kebcsPkOMZZx6dq7hHcss+nRK9y6cCXs3PU5G
/veMJ0Gwe8A3R4KM2XIngzQrnWkD7vjSepmz5/7vZuR5f4CAeAXFcYtw0V6q7HFevTHFVhn8crAJ
EcZg+gUZxn+BnLtg1Jvq7JKEjcy8Y1b2XFwRjpZIROya1s5HdXqJHULSm3PATjxuSENoYSAw5Zkf
8XrXglVvf5NRPNqWXToqKoGXfhvt2xo71v483VBUlRKZr5ZN2oM9ofSpFxzlhp/iOYEqikQb/48U
vOSdCh7zRvGE24axgiW98Upufg/vpJH4idm/oBlXiVwMhmsK5QH8weTakqcqZDBc8RwQ7z3W6LS6
b94p69yu9hmNRNvwBXLsyLKhsNAZWVDdXdvGRPn09s9sA4BuEfBPRcm+SoONgL+svfWLias6CPSO
76LD+ebGLkR2RE/e9pfXw7rSpEOsaDA0SEHmQytqYyLmhfxvL87VjvVqyz0RKvBHFpWEQaRr5PhA
XQYVBvAb/nPlTOYyf4N308MetaE1jqcNEeuZidakm+f8vEVKoplvleoDx605/EZvaWMCKtvOCrhv
959hbfaGv1eVS7gbqLXgFEZFDcsQ2nwLRM33WmHRAKe7sAl+rQXgrZclO9jKseOSv3u7GkVLVhe+
FAby+cBfXwJMaQ27WmXdhMVRyp2iuo+sa1HdwcM5tUPjATvrNu7wk7kTwKLJ5XkxYLXqbnCswLr+
edWHZb8VXQN+olRqT8S37Tab+Shcoxn+4vonq1HEGfKw5QDNvJMLXT0fpoFXhrk1uJrjoJ49LJo9
mVB2bN6rGGraFDf+t3aC+62mgDGOXPGThsZzbHn99MjxJFkfDcMsb1xhgYCcnJbeQSqRlccHw+Kb
nNOGt874Fh2rufyaWezH50C8iFw4SwqEeKs5dVGd7XBrXzM6bl+48QN8mGgdmNXGAhmk2pCBWREM
Vykvf0oYb/Z/6yLDapdgXG7+eI42p50BxGhi1hxIHPNg1kwuQY2H2PNp32wG83tygl4hDohusMDb
b5OilbF/HmjkQec9biCch8ilGxmtERO5Oy1vOQvxirFsC3S+sfZjGlvTkik9yPg8mCF2Z+4EXRSD
s5JCfrB2w44c9Xb5DNnXvEE4N+sJXEl7MH/rG0NRKUU6FhwZ/oyJZR5QU+tbzx86iXv+fsG5MRLI
gz1u1+cm6hJpx2LyA/6ZxPbwFQFj0WD32R/lrviBrFwT0cAIypp0LzGPnCf+2M6VVLDMzV7q5hNi
/NIHLN4Xaaw32zH6JcNs9n/FIQ+fZGK0Mi2q+GHyRNBzQRyY34FZ0yaTiBSJ/q3GMig2WkkAje2S
Bq9aDBrjP0LmhfmqDhV2Q98Oefh0XJGxS9A+jvIHvg733wXALfinoQ7uspBPd0il7CmdubggJ5yQ
MQyAJVQwbZdjbEv0EJV2Mksw4c4DkoxhP30yggxL6P3l78HTyfdEwIiQxDG0ewNIHGR2OBOO5Pdm
morT6DHbwTufXegif+i2awgDqDV0EVV3dDQNDsEh9y26vQQMtIXkz57uavErAMN48D4vubAvYNoP
ybQmfC3dBRSqqcDWjHqH2+GH++cqmBMOkUKPsHDut/6K6cG4EJpTwLb1AtstgiD7g3ehuBJ25xtB
Y1taofqcsmLxRmshc8+hNcIc6OWPaUJ8LTKOxE3WNURCXj40cbROMhXOq6Qy7P1cHBJ2+kLrtX2j
H7nlsHlzA+VUH4yyh7RDi7yGrdUcf9AHICzANll0D1W6qtozsr4T5jQmkXm/ptfv4/wOk9MJ+nkS
am4Uc3AoOU3hN+5oHwmQjHmvxDFQAywr9jw2tUuRXtvBtmS0HOi50C1P3Ouj55Ku8a+hmYgO3lN+
nYosEIzuIbhdP2HOMQIbC5Ek6OTDJpz+66DZ+lvYDTIX0bAbblwsR5/ihnecsI8N2f69Pio/VD8u
2tnTpUFTV00tHnEX7/kaKpCEhJoLhaA7soHw8jJAg4kKyn/NjX5CpJxvd5LIJL39VY16IrfDibMS
yywBo+eyGdkR/C/PI++I3qm59LDT1gsPR3ZKWQ3CJh72tCSZLXxHWjQ17or6EmsBH2MLktirRJXT
42fZVyblbGihSsn4uj5hv2Hu0Yl7VSiJ0EJcjnwUEbntmr/Bkwz4vad55SUMFEvluDT1MJbe1ZVs
O5keAsjaFSgUcDkgBS7t5PgU2Jy4cqLTkNXcSRV21dDPqdJJe+itvOUGB+qaUgCn78U1NjI3IKZD
vWYvqqTUefjYQJqy8Qb/ve+QJInD5NDJBPExCwTugyGqdstrxu6G/XTLRqy2lMjIdYUEZpqiO0b4
G1Wu0hSo/fEJGvvtvw1QrvxCSRbbsYYw+V0V3uDTofjhcgF5MaRHfF0b/YwftGMarGMQh3Q867ZK
Qr8AaBOGSrFztqANca97UoPuKtMqbNnuy4BeHPmMZIJHxbWU/l+kI/V5yDjS6voDiUjhryXFfWB0
r0q3u/nINxbllEbncof9O+T30qmQhQpa/n+XvxvB9yBh+ccRQ4ZyP6viO4NlK+MlcqOuGMYaWcxh
U9OYzhyCRwyEH7Ed2gjZPoiUKdYviPY1o/WajXoAMdo/hnFGZvqevzjEdlQkNXQTv4x8T7NwQ2o1
zY8U9WKqIH2OP3XYgxh2/ykMgUYVZ/xfgLcnFYutZ2VFZfx37B2xDw0BMpwdsoKyd+W7nbC/FenY
sz5fT07wp9EZg1LVxmx1i/29TvrWiTkA0Npbks9Ht3Nkzl4kTL/g32vf99AzOOrovRU1HwfriY6Z
KfzF5seMA6OpLgbsWfA1trYkcG0YVcDckApgZ8iHcFGIUTD3i4CqfRqZPZ3ahkXMbK7Mj4GGJ5nz
iwRerm2QZ8fFkMW7/3k4gBvW/vOio8QXvpWch/SN0JNq+sNi8qXGvlM6XOT/rpb9Ale66ijrMGvz
kvaXCEyS9leeYxe2ugNTK72lKr5B0DU1V606MMymzlhjkW9oRsD1LgD1EE5O81mGqnxYL7dRWrvN
RGKvg7f8mWAT1RWsWIc0mmKrXzetoMcUPUDJgXPf3U2geFv8Qv+1yyCnXQkymPAqPkRKbcVUP4Dw
8Jnw1S1elI552cMBsyDqh9ZDlOrvV/z+GiNFBFNbczHUMwoihheNHxVEh7NnBvq2vu0Wb4vZGfqX
oIHqgFKrHdxYBUVfy2HEhjHuW1w424+5+AvLqd8Y/4Ae1UcaVbnU589dnFm0v9ymsIap3+eQ7DXq
ZqlUhnSCP/RTDtWc6ACjISyetBFrAusZ3V9JBqdVbxNXY+ed4qN3L+SA+F/SiM769cDXl07HjvHQ
Acv8om6CPY1TEgTwpoKfKNsvf2uTVDdIYSpTifTnpCkrQ1M+IgVvvQjPfUkJPiUMuTn7fDT0IgVM
MvIxFNQ7VgQkIhwcNdDuiPPMvfjE63M40TN0UwXb4JMVsNgUeWrTTiWzXVkT3R4JEE9i818mJsiq
wF/mpg+3d5tIsZiQG3y8d3wAMTrTACHtzl+8XPQRaOyaN8eaNlO48ullxnJgNeXpkdy6dUmNn0H7
hpLxdLg21ysgWrM/8DoJlReIFprf80qvn61yYP/CRt52nMx3+ROK/+xjgMJOenbkvpYew6DGLa7Y
hWlBC/Vac5jvtZZifSji3j08HPQb3sM1ZuXcPmRec4mV89ujSv0FU6C/zHL9zAAPMwzls0c5MMGT
PWNSFpmlL+NAj12fkSSBrGqx8noGbQVsNRygpwl3quzBDt0robK1eg+8DfBn2/GyoFv2Y3vheA8C
0z9AL2XPgldkp9q8/z4M5W1JaSORMAwYnNQD/L8ORyyK5Kp/W8o8TlpjM33//d2gjVOvtYKh1i5T
Ve/q0FjWnsp99yBGpsINxdK3XcoB1bO56iJKSdoiKwekhnkHaz64qIMPQJe0281GznAJqkPqPiAF
sEu0s6Px3NOS21R9zITCjE8aL2PDK1yd1T/zeCCVX5Uv8yoFj3db/0hufcXp4N26NA1tYky/Ikb7
vmlnQZ0/ldDXrw/007WkWkHQlUP8mxa0u2T3Z5kvXwMvHyc0B6r6rWooawe/VK3c2X/8zOXwx5ND
WZQBU5tpSVrM3aRigSvamPsa+VmZyT3LYiyMKBTOjDSAsGDH19sUJavU+NDndoMHwIyOJnkQxppo
VCB1cvJe3vUGzFfTWv8lJfMH3g9/w94gkXh9ztsm9bKWmLYKt57gtWdbvsdnqgx/YbcW/iKaD6M9
5q0pVG8fR4Tw2fMtE1Lw6MZk2xYhUkQGvZTuGdtNPNxtjTPh1dAjhF/Z9dMeeEWtFjPxKNZsv+Ow
79AI4ssV+FbQvBZP5dliHbDgmhYTBIZZcbn5NHFxeWCIktmevdPvY1JL35KPlDRD4vQn/mPsVOGB
CIAN8fBhVVEJgkCBMCu8mefycWPanxyosdY6jya86JY3QohzqRHMIYBqQUZNdAxqgerKfKe0EX/b
fOEHKaIXfzY1UtRUUQY4NocmM7tYrYmjUA0S1M0B6fQSggRZc/SubB3CYi5lAFDR+SG1xD/UCZ5B
O134nmWZWefJcuyzAl1rU9uqBIQVAHeyd3TMI8gqbUd5iMiLDBjin333l3AfQN3pCAtNmE0svKjf
mEIyxwmCQyB8cMclel3hzBOUad0X8rdisw5Cb1n2rr+M7rrg+1AYWGDOHlMPSK3Yp5Zzs6tVDqWl
h4QKFvE1CfJInuq/fcAgIMFIpL2BuNNvV4+hHu1DbgEWDeiaTS1z3JiHGjYhCYF4L2tCvtcUxiox
/5tL9sYMmreZMI9TFvLMVZowd19V3UzpbdKolj4Z3/qI9rsCx37U1qSD0KV9CY9nAWzx8ycThxHr
/sluR4RmyThz6eWN3+5bx4ZhVmLxj7qYJ2z8SREFXq8bVi0OMiDtPejxD7Lj8yYsCrUSXl1dntjE
7poHh1ZiVm+o/L/Lr/Z/n/et6zQPjwZs2u1GKCM6pYXBuGPEDTIhJ0i3yGWg4cECcex/E+q3UvnP
CoWoRIExtSHavushdRJXhvtxNY8yZr6iWlQV1STQdsVJrJb/YKVNEIOYtV7sR/zFoUe258dBInuY
TIW6Lq0+JMlcgYzNit0MHPVYaCkhsDBnt7QcDgQxcc380harCPvy8T0FerOqCbFTK7Da0ubWN4BP
GVWAH+7FIbtdXwjgngD+kBpGVF1ZsD3Ns9bADwDPbnAZjNx+cs8hnEfBy+AYf5iRyl8ukIqB8PDm
zGlOpoGUpHjwphhpDRaxkyX3GL/u4P60oAEnR2a/TFve0Jv5t35+zHvDJGNON55ysd/wlTB7bmMk
gI2UKVAvcsYhfDtDY1t06zrGFuTWCRVocxTOhk7oyD7pC1EKs+Xf/39C8ESvhXXw1TfHLpBLgVea
D/mZ7nL+hiS7HfbvJUVkeROZzb+6YPnFtxZAlhMGt2ZTBXt60qYmu5fb4mAzDjFmlYQB5O3g1krb
nv71Z3OoTVGFlIXXp8/+NXOcUSDeG4opkNV7S0BIKl1tcf47drrAEtoJ/6B5V+jRGBepAyzDz4kp
LejL57zOUXS15K8QQk1GSwQgYxpDLEQdt/4glgUHw5pTiachHYnYR6tpPLrOqzQNRh/lY/UpNu1a
+2a8BiiMPUFofP71PIuLqWK+pIMCuZu9ehvoG7MMfaynPBx5/ZuXStZJkSD/7qctTTDrXHIxJ4AZ
R4HDphDCzhabwyNMV4G7jS+epcWjFJiwCqAn9bZ8/UysPlvsOdAmpIeFpmpCmLjl4cAydkcKbfj/
NJ/NJHEv/7pBJWghaUzfZtTuma/ai30IWJ58xx5bhAFKVgbT4CnCCKts95WDtyePubnOb1xgfG9h
Uat5PxF8EDhIWtqEVUue5s2CE+N2PxPs3vrkD886dbE0uunFxPSM0tBZyMPWhyeN30rMrzZPA174
3TsNlAeSmNichz8rAMbKTspCYn1hBJRHTU2HKv4hPiZYjEU3kKapD5qDoWJpqTFIPckB8+ZCzFdm
Hl/I00a1DGM3wpF87giPtjNsqamNlo4GeAt9PEm+f9dkW56J/dGfwhdA07bvgHOjraBRpqvfP083
sYQqrY3Nvx7ejjF3o5ML2U2seLN3Jqqh6PVCuQRHvDO6H3zFYc6/oWceaE4s5gaLS6416l28X0Re
aRs5dHZLDbNNZgoGS0CPbjVP7pXUXO+RIPmdvJlmjBO+Dy3HcYh4phLnzMr7L4/WHJaLJXtWY5jQ
gCwct5Q5cCnDFaCTAoau/yeLIva4l8ywQMsok419VcPyjwv2xusIb8HnEPjLTloxCgPwca6ERgYK
VXPuDFnCHbTnZdu2yvoECxLKolyi+T45QDwn2u5DiBLNj3O3IfTCB7chQSL9bYPUt83U83nIl3HR
pTQ7kMcIy1FIErTCHReeRGnaRHACanThbcmK2fmCz3FiLkhvdRzG5SJ9X3+SD77Pi3Y925TBqhKs
8KuSESIBMiZ6waMHykkVjUd6DilwMWtmLJhhZnt0qxDaQ2kx2V8nSB0oFAdNDi5xs3orxVPpvDa3
E/db1/Fesa1OJZMbIAneso5UTWj85F603sVK/NgyHdRYnNnOJoIVTNV6y1IRO6Ufaoqw6sz3L8kC
FHBEFxZTiAdyIs3mhQtPlIZEcgguPHS8foW9byLC+SVVUFbXuUnYHpZBBbi5B2ODXHNVxTb96cD2
WbCDakJ2CIMHYgq809LjQmg5eFajsUAHuTABF6sCzhFtok4d7BY2uJUP5Rj7COLRO3ajK94yBIcO
q5ejgJ13wVP1kchiTSomg96eUlCPAt+EHOQlCKx0sTPjJlpThrf50zWTsGd8CRdDxXaEEpOeadhZ
AtInVbeVk+7Hha4XsDEev4SkR2FE7cyXSjv4TW6A9j9mkD7HDF8yoQ4Z7wd/4MUQtELkzQb0hImN
Uvz0SGuyDmki01+WX3fYj3ZKlC3xJ3jvU2ogGuWbSKFxWStukF2Uen5yQq8Ffv4RqjNfeoAYcBzl
Gl0rACOc2iWPVdXb00Wttrzyd6Iz7LGpy0PUnjTLM0E9rhn18/CmcW4uOdUlb4PGLMNqB/3fMXQk
7k2+CbqaNZ6A04eh+g5WqtFgcIGq8WiqZiGU21alBo1pafdJr/gnur8l2M1g13ChNL0PUpHxDJA0
PBoxqHa/u9bOBtdLtV9F44zEr6LGlbRM2R4YNvnHWX3ijm2T4Tcy7yZvZHM7NUk10Iqg3r0bvxCv
Opuj2UX1zNMF7aq4GYyT8URjFoegR+ZcNjZqL5cPHA1EjzUbx+b4CFJaR/L+3HzMqage/3V+UZnM
1Hiy3I7Y+tX4BUl9UL+AJj3xQcasg13QtzabwXTQs5FPkSUBqRea0KafDqTKqdKcIqx9lEu1iILS
cj3vtk9UEzSwb7y1P9EPDYTEhq8y3zByLfjvxWu9fy8G7ziuvhJnUhcPu4Qai7ljyDzA1EF/BCwh
liHvcq7P9FI7cIujIIH7HsTuxpnC8LGGFxOJAOdW5ra7UdFQFLVVOAcxL6XqQhYszi4V9dYul3mq
mEuL0orMspzVDkLFT+OL5CBS03LPM6ZE6uRqPl1rMzYFn1yF90O0HVwcwbj1M8GOewTW4KL3r2O1
xB7ku1A0UpcIP1XFzklZeJTqjS+RiB8lstobesKsq2xxV9wE7RvS0+AQoHlBM8nvx64MTTt9ULnS
NhmjOXzTH0T3cvO9m/CxA4o0fDdDedxhirV+1T+pubiIgh0j9L80DxZ2Nz4h8b8ww0WppXP1bteY
BI/Wrhb0amgEcgwEAz3bO25C/X5PkCqPHnXyW4ibBXoRnf0YJ+ufoeufIQFo6fugSlNQZ1oAOzE1
MLsQ06d6zvvaSnRX9+gO6iWzJ5Q7SjKh6hgAgxPF7QZDC/9blKjDjWlR3SvHhSBYhOSUD8ttCrnZ
BqkvjCCzKZHO1RksdSJB/1eLRAzAMQfqMqHIoYAEfFCfQWk2Xrx1Yk8Wl0VpiILoVF5AG0+yBnxx
ClQSGzN/kK/ofQmPru3oOPX39/XjuzEi8BCR/v0C04cz1kKPHq0LXQaIXqTU1Ze81iEj3DrbXm/w
+jHk3YzUDzWRg4PIOIq+VeBJv9rJyTm8amjhW7eqQVTd3NIJpf0nbZpjcLV7paIFZnd8Xy3z/zhJ
mev5sEijFyATVWOH3VSN1ldI5mG+KEHQkU60u93TX6r46ksxbL4z5w1eKO90PWi2lcgOD30Kq9XD
MGxZPlW7ngTEt2h44aWH+DLiFqXFddIklV/pAilzc4VsqwDQkZWTtqhc91APSLzU638yBEDb1W6D
9VEExLvkftnAo6NWYMixPyPmYQcNNmjP8plgSQ+HScDPMLHw/is59RLzNirmhzKHKLKT7kb9BttN
Qde8bR4ZYenkKZAdRlwZQpUCP+F+D2kogQXTTcaJN7LMLOyLtMOvj25f3k131ycf9QTy4oucDq+a
F9wo2xQl12lhtDQV4Q2wEhPmUN1ljPflbMGUFi5MVJnYQ0siZ6g5QcgihuQGN4rhbMQEu23JCBgP
OkBgJ2bvpSHZofUB0o7QhPehqnqIklBinJ+z6Q+3mVu8B/kRylQhcaup3xAsdAMPR8LPUeEwUaDJ
ChyC3drundvI8BBmI2AbE3Avri44BU8lm0dFvq2+YumcaQyclW8ibP3ak1H3VV84ExEckvDZ8Fn+
LEwqKAMrGZpS0LkyAJHGRK3bkBGlzzHBDYt2kaJGRDcSKNqqNKcOLXhRd+Wl09tiWybXfm8mwt5l
2BpMCO69/nzKAi+FBWLgy2gIKHKzlVZMMnmAEDLZB6uuwgb2aZDQt1zVe+dlYVOelpyOuTBYN/lN
QBG2VQtaZImoRikDcvOguybAaqMgraEQyX1tiwUziJDfiuQ3OZq2WFAEkYcuPMAuTN9ifnEKaIOQ
5G6k4tSPrEIKNqZ0RAbOlsD8EgLXSj8Sf30dwgA+jd7R675qjlWZe8W8GHy6WU5xXMrqv3LT4Cer
+k6K6GkPo674IF4lfTrDk1EZ5px9bp6ylAEVNYNWmo4iuFpyPGjaKFnabegaf4DoOmXWt+6l++Cn
L/dVKnf/A2tJxpv9oQzQlmoyHj6AyYAuLp69ZThTDTNce/hqqVPbR/KA8GyeZQGbSxaMKHDOA8Ln
TH5iialBuKYkPm7oEd8B+h6ajhkobjXfL5Sy6jZSe1Ea+7hvP9WQACtZBg3xU9FiKr9AmnIZNfX1
yn7oyzsHnKHlbPiGQJWDzMj0wPJHd+vvdlrtNTEmZwXwZ1TGxffO3rMq9or5jk/zQUke739D+jFy
nY7ZF2+HAV1XxAIxgbq7eRym0uWRdjyUlq4tiMxEitUmDBxnwdaXNCc4N8ZEqiZcDxwF8X9j/Ju8
jFz7cJaO4nEYmgOsGlzFLv1Z57Nhy88RVe7mDuXWsaKn3/Ez2Z6KZHE1wkf8WMSzooWmEjKzvj6k
qbXQ6tx4PGFjAirHEj7yi3/9fdqHzQc/eAkJuFrsJ3IsZk2C60j6Ygr98Bfj3Sg6OxlvoipyW4WR
vapYYokgkIkW2hbR6WBiTZxjULxrJnwpqPmKhnN2jIv6ecUISfr0W49QUU1PAfNwwhATNPpoR+tu
BIwok5fG+FJM/b8u7fn4WzQ8r5eC7PqS57zcAyGbWC4Fb9/3KU0FL7srmMIs/mDInrieTj41hHOL
TRxRAKiBXS7IxDQXY8R+2XQtMrJ8nHXhRrIBPFady+/LrIaVDTQSpXdCauaJdrUim975r2wNLJiu
Tt+He2rKM0Kf9BX80lAcsmQ33hRSQDzrB6eyeTONQhlbYuthB4vBVCkST5TUinie/uxB5N4eurrG
pFfhdbLqIWLb/t4Qoshc+0Yb8iUG3SfXfUteMO0Dfa1qL5sw13DVQ9ADhOujIRc2ujPqNr4hrUUo
Z4W233v2TH9CalNr8zVBeHEqgpyAk3r0KMLu6Tdr7Y57ejuVgeV8h4TVd/zREnyXSK08BIE8zOf5
80bxVTIgzlAmU0pFSNw2niLcHYJNnnbwYVnkowYvWkgL4U2+8kCyuWpymjqUWV9/Nv12xsKtaqhN
l4HwiB8CaMOBZHqq65kfIObjOC+YjYs/q0MDoK+/Rq4z15daoAFGeWMvj1kivP4WPeCMQucki+vI
ZlhowCXt9EDWLxkLhpZtPdLzHjSeXr/tNK3bqTfTVTjpSGE6dxOOliaW8jhB0RsgLG9s/f+yxu8g
BjP00a4WQjWENJQLuUAZKyi/1ntCDAUmYau9HYUNKbXtPdXUYTCc5fviBJ6xP99YvDTFXKjR+hCV
7b3wRxX5oYI+Yt5aVPH10Z6t/Lhbsxpwtv2Nb309oYtd7u8RY5clNrPd57ZJs4Na+AV+UyP1aARn
HYsfqSMaraamgFykeBY3E0/yFHtn7R4d+FoCZ2h6V1j3orPCd5dzqZznErHvUCcTsUGGYvS0F5LQ
/kuQvOiQv4DTDmtrW6d/3uGvw/Wrg88kgZMkS2FpXPiZ9D7Q2VyyCoHDke7J1FSgsWAuhuqFHEqH
RpMyH/EU0IChtWbcDO9pj83iZMwDxXthB+yksp2y55ACbQNGlUiTRyWDzSVA5EbLyuf6ty7TUqKg
CIG0rq92m6shn9/7jzBRdHthDlT3f2xKJzlM7fCyW5ZaNC4+n+vxolSKgHa6dd7yPmBlV5uHloxd
51irL6uz9rEduAPHkkJ3mfffmP2Fa2iX/N8P4+CTHgaV9gDrbtSNB6SNWZRYaJ8Sj96r9HAECK+5
faeLaSnhgQJPJcoznmLScSKdqG5fx6LWJ2xtJF6q93PeLJv2bOCFCv3lvGdp9YVZzrh9nV95e92x
I/Xm90G1ViTsGCOrhGerwjy5PoD72+iJnoCRj/NivTU+JRIVe56W6BfLUWzoh7iOc4NlbZ05ZKvj
+/Vltm+IwOfKT5ufAXRQLVsS7hvS1cLEfoP/AcgnmO+89eT/x86HKLQYlwCfhV32cNiMNWR5tFnM
DSoV2iIl9/lJnTLfq3jJJoEREsbTYYMCwpaohEqT1BdExxewZsjD8mRehXD47xp1L21IBQuuPM67
5VCZTjGU/0uDByw6zzNwbJOEGlDv5S3hBWSIFqAXf+0NH2ieoljW6KThh49zA3t7WmAjECB20MFR
KibH1BDaWCmq9oOSbNyAqcHD3c634BusH8z3FasUTHnXoWv72SwPlFEujrL+rbcPcn0Mlrf+hE5R
M8LZ8o3HNWUYBKTb/ZIqlf60Sv009iFni013+VqlHoam+ENY0YyVQhoMBmC1LGNPujBjObjOAzkY
Ca7hUXQbtoZ4StLjV2AkpKV7oVKdlp8zypYi2EBm5oQ0+o1qvYkEDu0hSgSD6DF8D2NVmKeGyG6A
alIfxVqZkBwOsAcbqzViF+aTR8czySWJ88R7Z/f2810QlDJI9cMW+O6g5qBoKi5/CHIQnd6Ef8I0
MN8rW1D3tF3GdLDH80OT+e+frXLIsZQmKVYy0wGmDQsKtaaPQ3bwHqRM6GutZ1IQ11MMohAeviAJ
3JNDUc+8X3h4fs6PNKvRRGc0SwHPI5SRhQLuAviI+5M8IpfedqV/c14qQAqVeimcDerFY0/egTWE
kvBC73ykc5nKicPm4LgYvi2vzyPnduz07lxL75OFP1CwWhEKOU+KNr3mvN6CvkOSJjv2A+Nsojzl
8h+i4wJAc7VaumoPZWQ8UztzMhjdWinexi+56A99QjJ6IVNcVmmEqQet4nLhQUaZJaRQIWxAwW+z
XsUi8NYKL4vhSmxUM39oNPrnhW61yVLIEbLNi/rmU88SKiLwIB8SC+VYmq+iYn4M+RXlRZ8rh44s
ysNPH7WbHkVTwYlHiOCYDo1FufAihnVn1V2vUlPtENJgY0WQrGXe69fLgbr3TCLYMrvzSbiXWjuH
JmTLu0PM2HRssUpS2NnF4kF8x3xsS35ZrWRdNjKDwAupsbHnNzvLTD2Hjq4Ue/zE6i7zBaam2lcc
SCElCXTqVbMjc8C62epBFR2K5gmYyznafolE8FhRunQLkppKxPEzfejwOMymUXVjVDYCj0MJiJgV
Ch06/mP5Tpb5cSdThkWYf3q9LhyKOfExSRbiRMrrsLizZNvZDKBhRuCjnlv71us0dXfw0vjwOniX
rEk9xVLFcw/DdnpiQrvGDcUn9l5S/SQ7+Dn6pkUmac0WNQDspBbwRE0DZqOMwK+qQ556qkiaTt4n
UHzqwBaF9hiXtq+egqBfa8TRXMa1tY1rKJxBKGcj1jNqFLR9lY75//d1F09se43uyL/dp64CYC0v
2IXAMwy1m9WntJQHIV/WCo6DpYaZ9PIfaMNv3ugcuzrvyQZWE3VTjZwDlgeIaJ3LiMagX2Zp+sNu
EyV0/8/p8bOUe+nxbLpvqHxR+u9saPJ/AoC8VnovfLSU4hZKkXMe/nCfgl7aIeNA8kF7jH4AOj2W
uiAK6VQHaImuWp52s/WmQwvh93xbT0uWJ4XRvZaPn2ltV93ivB92VE1+3P5Fj9JJ7USjPOgliWN3
cipx1RFWh7hYpmNpqdLqpfVSEea9VOBFyTZrvr9AZ6OXMNzutSleAIfuGdELsaXha/axymPIfFhS
1kISZqVo+Vs/j2X2b+jnpnz3ua4Fi1exUdl7pYmQHSozd+gR9rpnJUPNo/Xf1qfP9uqbgDfa9mjg
jTTag9Y2A1NvlcVq7Fwok+DY5zH5igs4MJVEzycM07A9gdQykgg5yKgbDCSVOvvmkjj3iIiegMuD
ZQkg2tHxBkJN9kHtoku5ea761EmD1LLIU0a2aWuZ0Dl7w/Ycp894cV/BsatqRXbusYIzJaS2mASd
IoFo9U5NWWY33FRZcIP/op0iP7sYbzjGhvkpqaYFC+Dg8rgLNI+UZbnBWoO6x/DDrnmT8rhtJr5P
jnTTED1DYQS2SdkPXQDqdC6jzeGIzFiznNn//DOanY5Rg5hH3KgiJpp9UUbHhP69edGPdO52uzJe
zCzJv7ZwoXyCmt27d5DTGGkd3BYGLSyT2NtswJvPdZfR5O8rVQjD2DrDYuneyxJqVubQbtxbRbJJ
HKCdoAeKbQOLtzN7sIc5bN/wZDpjC+hbx+7Zy+fInapl3jGTE+wHcXQsglGQpmd67EgOjAlL3ZK0
H8G8uxoENeAG6Lm5Vcn48d62s5lR2CgennkCK/FeFJLpvxHgd+OIL9GEo2PelrJi2akj9VJPFfKd
YMWNWVO0FAqyjDS7dZjm5623SE7+lJ/E6/iwSZ1smCN1lOsJ4Qs4rke7Yv51UA39/YIm4djSCUh8
qnFAftppRUoJc5/0SatIk7zkeLZVBk1dWDZgilDSbsyj6i0LyxVlKvFdqIJBa6c2fsEaeD47rEbg
26GBm2324OTo63dV/uvRs2FUfEpx++MFrZ0iSQssmEIHghyOmFuSldHwy6MEms/VgR/cLPjn5XX6
zuw7kDpVJ7QQL4QCokYRFRogwqHHtOeAOMKZg0vi00VzOS/fA7IMCNJH0PPFFfmuhirv1XEop+/q
/w8g7jO00aLmpYOOlhSVKtdiXkqMU+HPAXluhYm5dY3r1nK0WB9ais+clvJlRe4OGCaz90ALX+0P
YKXJICde5T9CiNaNyk1SmAMAjqjIDTyr9FbGMoMBxtK0iOe2AwwGl0esseaiXHQR9ZxGKNmhNKZl
9mfNqJNtaa9WtRKW3wlhobanuib1X1b+A4bO5CtI9nPwL9URzGmwb9iy5862UCi1aO1JKxush6PY
/Mg7jjBKMN48MgZ08JXhlr/yyVkL/d++jzFisS5c1zWZKRTqNwvppxPt+A67ogpGd1wFTs19Zl5J
btAfIw6e5iG/fa0SBeT3uzJRv2RYlzkldG0omSfmpN6oqU+FHdPfk8liThZcYoGkCzVToi6un25b
61UwVxm+7GWfrv6fsgY3TnYg1gY9IMXO2NGSpcz8HmQ1pY5KQEQzcRiye499s1BAUmMz3WsPJJ0O
5S9rw9qXtj1VZoJ8kXsijpzjUQib7aEqy5xqqo9j9+CMXt5uAx3Qsf8T9oePFszksYCu389B6z5b
iLLXIlmR7LmBJPyUlIINkQIlwObedcHNz4BwYluyfVhxUVn9aB5IR4MMHCIMw+UWykp+spd1Nxf4
X2nrTIpLIZzNy2Hq31kN19IBZbftS7uMyB3Wq7NhQcq934bGZiyOdN6of5CthNceJKaRfomDbtuO
cGtZPGWkaTpO83artCLp99/KaR0bTrpx6LXl6Ynmd9j64tCllV8VDFxNcHYZctFlQKwmoniNc0xt
C6vPF93TnQj7cgK1LqRqaol6kxQvGdx8Gjsy4A1NLh40MRuXmsA7DnY5XkobxQOQ1ipFZThFtfgG
tP5SlfJnz0OFzxFURSJMG4g1nBboU7TcRIwW7jtVloSg0vQ4W84cuk28P2+Psn/6H8kLmEw/OA+E
EFK8l+0daHb4n5poI2WzbI9/Hx0/kcwO+67uwdFYtfaDU9WLog/++UJVq0l6oqdMrrg5ElpO2fue
5GehtKdnoKRmgKMJ1EPr1mgDI3zm6xQ7JG4NWPCFDB3zNO62hWQIc1sIJbbT6xi7RTNwLWvmJURB
HsGTip0rnYk5PZUq/BK9oN3m3lF7kDidbeaZORtKnuIsZe76JBYYHj159rpvnktxMrKsgxTzya9M
yHhje/yFPeEjcNkqsvz1MSxXtQmoBlKqtT94gUiChv06gPMQBzKJz29s/gC4j0YZovEIlB8fMhaJ
XaJMsfdGk//gPtmEi+u/V2HtHYAqh1LO2HYqs9CGRPiL5PMjtSajcrrlx096M6LqARzEXFg7hW99
pQSIZSa+yo0R+biLzsMrJypFU++BvkKnprmQApEJUSJyidtq3RZCpWzt2MG5LisLylVVIobc4his
8x186m2SUiIWI8FS6v8EDFrbNlTNNVt0CxcxBghQ8xdB18c0CzPOh4rUHKy0oAU4I4dQzZH0J1vc
eJYHgr7dBlLPEs7NUNKM2Nt1TWw0UGrcuMb0DPMhOrbTWpelfKJW9cjz7laBqPnPnaf6bKpcNF3L
kOf5sVXuOfcETndNQkTE+0b9qaGe6L+ZTnyc/EBVlnOWnOsU+kSbpPILkpWNf6lAaz7id0/SlyMB
CZJOsZ4UV2csEckHZrOWudmM7NgtbQSKuyg0SbUelqQvZu98Gl3VqwJfJjT6W5cNcEGKishV/nNQ
GDFDsmLGagIESsOG8MFndVgcQ8nCNU39YwtwqXcb2pW75DRjHgixbXAUtDj+/NuKXT7YMkcXgvC+
wvQOTlfZAA+7lHGBD5iXWTY8sOPhHzRRW2CnNByjh53CDtXhGzAPpFTEKp94+FuQROAtA77leSi3
frrHrKRPI9IQJR1tnkRkQfZ/No1k5IfRahFVSmky/qy9i/nLvuR3OEBEgircUnnil89TkBjqrcoy
vGKfJkyM4whw//0wA4fa7JlVtHKRBNmGT1vfIB8bGs2FUJ+/tZt84/M2FbrIz1uO/x6h2BNptDdj
mF+E53qH7CVYRMCk9W42O4NgoouLYvduvKoFcMU4ukPWKBX+PiPQ8KIXZ3rCGVvdMRnZR5Ge9RNp
+J4kAPIWAe9BZ2R7lUzh5rYDr9wTpP1bSvIIguonmu++A0DDi2R8ASPX3ujGF67JK9LAAEh4o5gZ
Mbh/a1EVEOMy672NUohVxwCcPuPkDtiF23aHuwZHdhxCHXj9o84d277NmrUSzqPadfGiBSOTNsvs
Ylwr05fmRSWSS404Ch69vtrEtc6EjREIDBehjYiLcYBUxwyd32yugfKnjaQCkVBDH5vbV39MUo5/
hedJw0Ki2qa01JUVB0BJxzIajldNont7hocblODK503ZMPEhgam2cMNnEm9np78tR5TenBd/etMC
/H1ja9Rzeq8HQvUp4cxltc3pjmTiRJiYSZFmng5vuN0GkkkKVbh4Mg5cLDt0buJBed1ZOMhdNVAY
8SwVcTc/brljko8jMbOrsHAdrcLdz0XlG3yiMBFeEusO0IGPANFVHP2/XBMtPU3g+HdYN54vo2GA
ymzRIRsjlZi5hqQemLiVC4pHohLxbEw6VkRWpAU1eSp4V/h7UmDgmLynY60+IaVPF9l3NA/VIoLG
6cLjzS/EtqcU+9dRNjJIOOKh6stL5Aih/2+cdNpnSPCkcljqxY5oG2wm7+nnqym0gIzKAL9I4Qn+
G7lnYvvUOf9tQ9BeF1ru6o3NhuwA4TjNi1aoK0wt3TQ+TQKrojc8tQ3oqVpJ+a1gIa5YjosOMFl3
rZHH3p6pfWkQgyxIX2Vok6vQ6Un1JZZs5KJHOrolRCN/izs3BSLxxmLzMSfIai9Ibz8vDG7+Zjbw
g/NEMDOUlSxV45+k14aqZ8hZHe4TXLjI4GTT+22eVP5npqf9vAG83U1fBsJGyekKqVsks4dsRUsq
+pffwk9vUBbDgDguNFPupD7a5L2jzJjthgYZ/VqFWBz9fpM9qH3IlyX6Hj7cmyzZ6ba3vdLss6Hi
wgYhcx9C/ysaypt+4/1OdUmemK8ElykEzZkK062+g3x9dCYU8e3kR3V/aFxJtUQthaLyG+AfB47u
UfSST4uxpTI7aH1ejk7X9D0qukz2riV5KVEh+s5hkOusf4Jm6ZUMR5MoacDJMZ2sRzzKMLq4jaUF
TzAZfXuTakkdOvwNex5qFDCfLdinY11DyJnm8EWJ4TUgnCjHMy8B19bbpA0biuPQC81Jgezg8CRm
1hoa0DkGWR8e5ZJHEymXgZQFGNfh2wEF13/nWV8wbJuA7+qte9nbFFtdPfPhew5a1m89nhybmx8S
uzGsP7kmRnps23o1a/pYf5zlAR7frFIw2kpUS1IbFZEHGCB42NGI4YbCKPprwsx0y6GekG3Lbkwv
VA2FgIFaj5WS7ZH2wzCGp61+ai8ackJi5Yivyh42znLm0xaS65YBbiGPKnQJU2cGchN+nRSuEPtw
VOEilUuu/G8r/HcU/hTvjU5bicSQTy7wD/1q53/3EnX433GKmBUCg3jx2h6rMSJo2zCXC96Qnyhb
qWcVtZpkV9ziJJR1MyYAl+WKzaEfXMOKI3H2Ca645eOjrz1sBtKUBAibc6H/IxLg8DnT2NXAe/5k
VzDtiq20Kz/WucXnG9pKPzDir4h95H/RyQNqC1ioL56MqM7VEcKQ65KuoFmeoB97ExDniibcicVA
2p9XHOrBlyy9NBc18dURj3/PE+E+f+9A5eYrkunMFsVAmE+1NdaOpgl8a7nYagROUeINkpr3/jmg
BK/1HqHwUol3jVDlib8Toea5sT18joRpkqW4+d9a/DoXOSWsMbgtzrM8AnoQinCQfQkpUAjGtRt0
BTjNjXVWCvuXahrlNCDZppHkdC+zm913nIsjnbHfXc8EuJ53GWmgcaYYnqsGnfBA+1r4X5A2HzoG
vUdCcvZ2TuMLwdpnKzSBtGK9jkv8u0iQvElBWw4tvdAx/+utituqfyay93sxFwOguis2aoA86LfH
WWueb/ZQcoZFnbhkWXSlDRfAFEr4v71vCjh2VFsux2QV8/jMbG0LbQHGk2NJgiFK1gdUMDeZCvUw
OdBRMke2I2dO5kap0ubGY2UlTi8BBTS1UYcOTiaOCBRU92ck5JtTZ2H8bkXdO9PMBMPI3pWUP65Y
Ceuu/sss5fikL+pfcepiokvptX5BD0a1zaeh5pXJIdF/w7TZAsY4YQk9ZYspTyqvwopg2Xt9CyAd
/UcAsQ24znlH/DBB4BPOVqkp0U3HQdesATGNKyVr9AmCk0bfUX9r62OILy1Awj0DaaH7HBb5RZiA
e/GsEWm6RjBBybrHsluDLlslVHaxxyw+vMxV2VIKxY10n8tzaKe/kzCDfvBl3Pz43oNnVsXe1i4y
/g7Y3ugE226oJoGP2LPPWcF+Pgz8WMd5Op8m0jRarnesAmMWu4c9bIh9gKPvnr48XcC84Hdlm0NS
HBZOHA8I7N+xI1sd10iFbXq9wNbk9pEsuJfp7CYOQc+SxiNHfbocAClPDCeaNCgIeenH1aZvylab
4y+h91xnT9U2GehATJxlhVIQEtu7xHbVdpfjB0Agt6cmSLA8LZEjg7OE1dismGmnSnGY6Q/iiwII
RaZfaWDILZMIetbvocefaQmGTPEV1gDILAyKI8BjF5Azh/u7IHQ65+7X2pfYty3LGFPP6neqttDm
ExtMGvimIF2NOPfuz+4X2yOWVGRozztz7d1bLylq2VLjvWqczWBnPM8VfERaTGJ9Zlv7gXssslI4
JIj7NLhRo0H1KQQX8b9K38aaK6iVNwg8iN+qzLNYWYs+1f93UCwu4q2LyZSOUPcgnoZy1DZRT1W5
hbkc5M6HXZDXc3bqFOcCHyng+hJsKe4QKiHXNjf3seGpOpRZofDIu0gxmv4sIHrHrXiWhI6MUwNw
tcXoSpmU4qBpDXsHusbJu1N0swHzN8des+GGPyK5XG9NbA6teX9bnA2k0+ulNGEq3QZageDgRi92
KejWoEzLGMNcDYi21oSyOM8DYihOCB020ptEBJcJzzILClw9d5x3M/xaq+O7zFC3x0CCTcjkJzRY
d77LT3bE6uDD7dt7dsMuACZqxy5ZolI1nzLH4Fkr2u9WLm27XPOB9Hmkr2Cgpf8zntyhyAkRzvXu
tIQnuAVF0538FXAQIJUBm8U3/1Sq9k20SFB0MWCOx86LHCsKUyMzU7ekMSYAUxyB+mFwjv6wj8eo
OjmHyQdZ5Zapjk8MOSq4XWXnZCmn9K7Faif4ilo4SulUL+AX3cMUNcx5C2ba6FC9rUkZwGIRy/i8
N7ESBdunySsY4n1pX/8yU6375hkNFIpVfjLcX9gz8cLyzV1ryHuEaI/F4RPXEbHz8RQefea1ly2f
2alOVon8lEMil5lFsPpFVVJeI3/Ufj91Ze4L22gBEHb3YTUV5ktNMfeHKFPRbgIQRvkPPBue6uac
W9aeEuC91Mb5+h6eLPdcoXIP/6UilgzyyjrNDijBwamDdUtsG6AOWaNpikpEfdu2CwPCnLHEmBoI
jzQvCo+30rMb1+wPSzyZQuUkQciIKJSaaqrqr/TARHSYq3Ah9O6TsrzCH11+cYjDiYp6dM9pey6h
eINhjvReYp/DNsHqIKr+ZaYY9ABFfqeDMmGWad2Ul/QMCC+HIEsaSEx224QzraIoJ+ujVO41cDtd
RYQgHaB0kVmpSidCPSXlsKpiEVSxD0M483Ocwak3OK3tYdGRnSUHtUjU8/x+kd2XKPyNyNtCchLU
d0vtZCkILgP08vr/xTwbEjCJwG1VKKbtYr+SC6il68ee7udz5srjXlr32r7F/KD28jtwvn/s1Q3Y
jIc055oul99SiaK1w2lbvawDngTmpT9l0uisGJfcQtXHz8YdAVwbx3xaIXIoK5GITlIKQQoyxYxz
89I7MCGjEUmO+HJug/M9cjoztlXWTaW1WHl/eUn4VDZbxrh3LfHVtcgh/6Hp1Heey/JcNFxz/C9H
SMQXarPu+UJlzSMuHjCyAvWkMz/OFO/fDfiO5ov2zCZGvqgoomlGEZyFx8earC0i6t2OGuZMmKX8
G2VNBa2n32kfKYT+37s2SXPRJdgxRXqSI+frJ6p+xfMiwd/EmuefFBKyWHuQXt8Uip0o6M7Xa8bf
UkScYiv1A7dNbaeanCnBjwaKPIXbR6c/rQ6iWTrB0ZhIwG+LsV156y0eiiVVW2PJgjzJs4bcm13P
JJSsOVjC79TRT5TDiLz4UBqykbgyZsoJRKYdxt8pHOCaI4aFsNTlhon+yv974rVCXanOBTY9juHa
lL+mXY4NyomeD88wA+ki2/tEEofUa0YHaDMDayg7t5e+UXBpxViLfKfRdN81/ygccgtnmKyyEACs
eycMcpjgJb2v1AqWEGMJtNjxYlgX4A5pI9b2a+OudRkKauuMR5Fx5qNeaDIelGlKLaSCUx9F5jjn
G7JPyar8nJzEdg0ykz4RVB8rG1li6Hoha5SQDjKV3YnsrrvTMEl6JLXBQ/82qAwCiEvtewM4n0gc
LvG1osxhnXH5YSwXE3MfYi4LHrGEz30xmxha2K/+OASdfN4YjGs0jsT3k39Uzw7XrLxgFSona+CI
3cRVGnY/JqhUVrL1a9EEmpDC1QsCLl2e81KYTV1lnJKS1ga+ewQVu16NirY3igI+kET4ZannTwwQ
FzNkY2BxWGBoRzcsXEaIN00qwltgwQVmwri+OWtJj5KOI8Woh7dSXYEC2JZjhHSzgv/5pgWsvn59
JT6vEx5Mad+uHXw7APitpD+6Y4csb3MDwyttpCkshVlYz8A+wFxmw/Pp8bC+5ndp6klINuIs9df9
fAlEslpglsLeBSDbJqQ6Q38R07wNRm/0RVGdqxsnAI5GneB0qK+cNIelxL3A0p2Hljvke2ttevwj
s2Rkhw4mOXjGDOm5n+t4KKFWZh58Ipt0gy0wQ5qflZHnWVLOghak8T+FGpSXYWmGV04mV7mKBAYC
X45sC/0MAG2pUx+b43Ya7Wh3sp5JtIAQ8q8lfpIFhFVqKkB8XcBegMJe6aEfi/+4dsMxYOrR9HZh
sSyynt0nFv5zoidTVi3DG0xPcQrdP1ZAhvo+dbMtoJYkvSZS6JI6IPYgHvfMsJPCwJDtpJ9Qa3nn
vJm7cqZH2Yd6lo+WjEypT2xRN6/+lia80Safn849j7EWwvONRbdvIaffPfuP3hqM5FKQIUGtfvvY
0pWM78jseKZ9Lny+i7d6D6JhEJvFhUbSuwbB8RtPhESCCc/JRdZcapjWRsklVmEQprJMvd/Tt6NF
7btP/v7QgnX5CROCwnwDAC61Q4UAOYKE67B8qsZneTIGjaccWeIyo2cZ5eyszsUyxqqtQqvqg3CY
L2cRYF1vqIGA+27oAzloEzaBkiR2W29/Ho4aIAO+ml17Gj2sfLoZKHFLr1EEvTQ0gCussxg2DFyy
2EFRRS3uJbyUZACmZgMkP270rk6UdwN6j5kGZH4y89GL3u4P20EJ5PozOgfFIiVjZHXX6VNHAL9d
XqsYa1NH1qpYsRCZBTDySVTTGCuIFD0PV/S5JJVNlOh7yjzEAN7tMWuRWHFC01xnVIpWWSWhc8gc
QZas04PoM1v6SJrC0MqGfU/1Dbq0auFOgWFdIoeKIEL6f+g4JdL0ragzczv8XngtCr0foNDAh+Zz
VSHdTOSdTer/q2SNSCySE3kkXGKi8o1R1JlC6iii5bMyJiyftCkj4AAEIkFwCRkeEoOeLvAxmKuf
Bv/lj6CyVcHIs6gUp/kVqruqBcPZP6j0A7UMORj7ZINR9v6YWh/4G3x1lfN2cWbMx4p+vv5Ez9Bd
eCEOea/Qj121YgBr2zc5SjY/UX0DPBLOXCnTQFRwCCRVR/CbkBijJUuLih1tV229LdohEoecQc1A
ornMHu9g1Vdu/pCteG36bzNaWW2YWC7q2cRfWi5o+ktk9au8MbxvC5J+WMncgH5xFTIDFp349Jjl
6btald9764pQmqT8N9j+XccQK9XtNsiyZdy5+XLZZClz2Dym7DRillBpeASnCsmAaTS/WmYQqi4M
VQkDBF/YEQcwsCjfhk4Rg07Wrpbc0lPpZLfqlOF7Hm5wUrCtQMAYDROnAwNXfqf8R0qXK5fRJ4kY
Lz2pMehaybf5Tg5krZz8k98uxqInBliYpzkRzgpzqC9yLKeVkBabi9AXRim50rRgHZMaksURERKa
tobc7m0XngXYvm4PTat9HorLG1t/8OBbrUn7alpCUSsrG+s18I3S99zvz5w/TpVKLn/P5VOdaETx
vZsBGJ7l2YkmaMxtkwLtlcowgm7bB4bOVDLuGThuF7pt+i7TYsXOc1/yyGQ5UaBIghbsvmkEHu3S
fzWCoQVlftPkaNgafUL98riAZu1wyQwCp5zrQMlwa/3J17ZmkbAQGmt1maz7mePos6khUV+Ylyln
zmcTDGcrlsYw081n8UdPKvN/pGBhKMdY7+rOByd6CLucF83LarUyQUDvUb/taNluGd+S2en0v1eE
md91nzH1HDG5Dz3cGk2Wa2nB4FiQvRs1LfLVIipdkVmseFHokH5mwvKSLFP/ZrCdiJCb9PpkjKpO
9LAOcFSBG1kYsMb6zw6j7DMBGDXV4CI22JPdbSrdTzgDNJGJ6u/05oIF/nAdLmWpjL0AcbTdbXi1
4eumjb3ySS4Abvx8NLLnOcZcFW1ZJ+QvMRC/UB2gRJVm+mvlX65puTevxq7b5a3Mgh46Rrcnib8I
6Qa4yhUbq8sOzIUQdNEy1qhWlkKCm7wzpD7aRNRXxVj8fqGfMXmnWcHiLxyIzzDkgJfYC5AOykLi
bIFBFNg5+E/3xBqUvM+zXLKxZetBsrVwqtqCkuGKt/5EifHrs37j+aLwa4CPvMYfJC1qPzTTUk0w
PmmsNx3mn9gxguD3UT0fXEm3ecC6Sf8DxZKsqVcDBheVpmTVCuUcKHZRMp9P70ZNu9cwfBrdxd3J
aWcSPONdBjLF4Jn7W/VvzFQecrx+ye23J6X5/KrQuGtRKd7XBVHHtDj3ePulTqKYqp93+Iz/BalO
5HzMLEocDEidNcBeQAY1j5SvTYN2MVoxQdImhk86V3K+eXBHN7xq5t0W68o8xSBMMloHXP0Duwp2
y5CWykUs5/LKtw4lvjaRWn1oAzpYt8BIlSKY0rGEgdtN3LRnVid8dEj5+Ck0OTpjQli3Q8Q2i5U1
kOkUjpWbGMlOFN0FklwWcZ7JvUB54fMrIWPVPVnIjiul0gvUiA6Oye9sysBwTxd6s4GfcBmknqyV
enHuNBnNxtVR547JlCbbC/q/hLOyy0OaO3cWDudLql9W+Uu5jHChVX1kmZBGhXgY1+NWXVJluxFC
EuJJamK3s05ifCLWfawW9Fo3fJ/TIUzJsku3FSVD1U1C5axZ0w7d2rUXsQwAHb+6fhHrHBveWNMG
LgJeUUer7Upe2Yy0U+eWUM2/LVabHxKPV1i938SRZ4Yfgu+PZH1CSugyjvnEfQe39x7k1qWTvdrp
vE2druMd/uFwanP1+nWx8OLbD96vG51Z0629tiTsu5NfIT5AYsRhRgGQW7jtOnfyUyyPAey0OyBD
Om7HA46q6bd38bMaqWkvWtVZeRh/SI24/YOuQT0+16ozU7IlSXT69bOLtjh3NhNJ93jIH1WoMXcj
YPjo40/MC6EvfuiOJaTsv8z6L1ot1gGYv5mo0Q9PajFpVua0E5oE+LEwMVi8FN0WA4eLXpCKQfHT
f6t5x1ry5Zr1jzEi/on9Uu/ET/BGPTFpcaRjiEccs0lXIPrG6M9H9SxLSp449luJ3iUi87j+T9Ze
/v+qrvU5CBeuixjrxzJ/C3gM0p2Tal6l1TcZVcVonXrQYRmzgDs1Uqo2U1tzOyZ3qxPqYHesnT1T
81mtp2X/77TIIYKz70dzKHq9yQUbgmwJcoEGiLmhJeMF4tHOJPDhbyDLxm4kcfzpfZgZlIzJ2RLI
DxRPnc3dgNN99SZ2csP0/NWRk9w47ZTm3hvojKnh2i2vPaW/f/lu1gBB8WFDM6YK9sgcCT0t8o1n
YcMd8xQ7yszarNxhbP5L3spfCFMOh5p4tJs+c312CiHUHQAV7DZeAxGES0Uh7lzJv/QKEqUbvnfE
hyqXtztASB1cRVYBpz9ApQs0NZGFeKZbYzgwF4n5KspBSevDP1/Msl20N1Tt/DUqeIq8WEtkPaXU
JxM/EkqfZI7GQgYO5Cug56ZFGSYBzyauZBKe0nhN3r6QfsLCBnQcbW9gl6E7uuIsxNWgAzdxgBTY
F7ra3THVUGLRpWZs1rtgxTdOVYfrdO836agnRw9jt/6uvaPv9W+PHTB8REOS3Z8ZAKtS+/q4A8Q6
LtBFu33QPNyYc4xmotj6ja8VzNCGB4ovtgzQj/IF+4oyCPo6haqn7ohs7t0AIqIK4Ks+JLGte3sB
M1W89v8CQpquyjMrGNy7euNPszUXQl2hU55QUx1X6q8BsVAHYo6DfZm76Rph+jBDk39Wk1pknl0i
ypM+XQBmxWRuhbzuNu8S4AH5IqUwj2dmZ/4oi90JxuKODC3uswoaC+LzClIsAppR551GulDQ1v/Z
gyR4XViYUdKWp8oJoVeVkoMt0uAIXhxrsLz+5MzzNcAxvYL8BIjcJWbebyIAgPJ1CyNNk0KBzJA0
bcs4zGfJ6tnXHM1u23lk6VS9dh8HaP4Uiv/uk/r1nNPCiGBN8wKQ0yv9w/QgEsjDzP8BPxy4O1z/
lpolJQo/OA7CuQdOuw/eJOvqg4M58l2X5vz8KpKQ2TAm1vc4Uks1rMcKQ/eRNuHdUU3t+DQwcHsl
MSDfkZDZikCDZ4LkYJFEyWCuADkgrUHuKez5Ff0gRS9K8AraezAuJ0o30l+61gDyS+5WURXiKYOB
VRfaLPnA3easFrKRIDdnWiy3i/+xPgigO8QO2ADkvGkddZk3goJlPCx0zKiw1W1VuHCGoPNymbQ5
jvlJPjJErUTFgYg+iRQPaCowAY9mMH2ru+r68tAjH1116oQEDF1CWHZn0nn1v7DsHBqZ8Mw6G73V
iyu3lJlGCTtXHL3uwsOkd4HaXJMxf8r0Ttr1Ze9BvAjfTBG4Rm50bSW5NmeJHFcrRLE4Sbt236km
Ywe/Mb+hKtCQlnA90adIaJ7Spmj58NXsvG7FA9hmbbnQO7gKwb7aBUKeQLZLCfY5rVQe9kZMFitQ
TFmkCKqMxll2a7LGvMTwUnm9Iq9myjfL58qXo78HwiF+3fxtmq5mYOSjzhahBmWrRJHNScvBl63I
qxzpQ3rJxV3Rs4O079U9Ay247RQ5e8f3HtUUcnIhWGCiSPbvx6Ta7eC/idrOoJUxO5+nbcbkiUm4
yVV+nJDh2UwwlsY6v/UcoFP5j7hQhzlgzSvCbQLHXx1YqZ8B1tXE8onhRMQoaexv8O5XkjSKtJ5Q
LPnuT/e9fKGJ01qVJArpMjyR0+NhhgFDXvN82rxnSvrzV9+dVY280S2mBzG2SUmoaYC78ZIZsgBu
MxxalSzqluEN7eNYlSPM1vXWGF2BmztwQ8NrGEftUNB0goZzf3zN6yzjqEHqwKAZJOmrhSKfLZ5P
C3k3FuwiK9hV3ItNopnIDxDKOtm+kc+mRHQQuROvbx5WgJIzuO9nYC77LNF/9MCA2JO9b9NwGQnX
MvKwuV0oO+/hsz29RZYwdiRMtIvb3bh3MX6fS/rA7lPKo+2ON9L393d+/qKdNkqvzDQlR2ydSpBW
QxHn0u4I4K6DMqVRDbg/azVJAUeBMIEla7NnBfEysRvGgX3RjIf6oda9w2eN1cNsTONwNzCWU6IR
nNsjNAvfDOfvI4wD0GSDVXvBAElWkz3wx21abE2fBSenMSGkDXRnx0qf+r01TfuHQ/f3qJoiJUOt
ZftgDDetAWAE2mSzyheQtTBqVDDdM7GIDN06BZf64aGA9QiWV78EN39Vc9OYoqVQTN/7T10T1jLC
SUaCYYzzHHjdFSXh8/vKMN6XnFNocRXW6lV5zybrheI1FCcmA4XeTFaMUqAdX9MrSNOh62jhwPGc
BH9W3S3ff2pOfgzb+KY0xOt/Rcnybu7WQM/ouqcZPiIQZwlspZTmkWoI/ihm58BkwpMgouOkEAbO
qkQ9RJ2jPq20+65kJKrn7TiFSSHZJfVa0TLFWSHakUp+JZlOV/6gf8yMvn77O3GOfjHwvID0e5DB
1tdZRdza8ZhWQIslnURO7JPvfSXWFIhnHGn/biQvYwqCO3GA5/UhXkculZuMo7gup+k2Arp06vEG
oigmUozsucq0NJj08LwKVlGEKjAod3GW4HB0wqVPHvazPNctslzzLbLvhnZMB81rgyzVfOB/9KL0
nNsN2jA1yHnluRsiSSz2wbBbhHKCl7NoPDgrciUbSyMw+hLxBWIRNuFYPj94eOs+zsdl+K7dD9zo
CvMsIp/P2jL7HkO0Y+Hdob5J5uRbpX1Kwp48Rjkv3GbI9EtBGa/kc5kkyFTYPO6gNu6zpAI5R7E6
F+PTQspykjo/llCPupr0X3dz0IrNpGd45eLHx3KDMKxgiiyTTfYoabo5VWmEmCSHhXcBPhtrEu8n
siH2YgPOnXpNG7IC7jnkgY4axOQKjUvXjiKf8GQdrPtlujzZBgvO6sM76kHpdbxV3IXGIYe8366c
qZ7E9QMTXfMYeMXFHhqEvtNfvwLoL08MSBuZxbDFm7sayePDqT/YbRoTES/e72Z9UeqGgmNRfYKN
Vl+MohQ+EtlkSO8BKpainwnO9sU/9rY3fGjGa2vUsxJm5YusOHE9CZ60kH4sVVN83HmcB3+JAiBX
hzAXaJ7JJbAloT870iM2o9ORAT5kdwvLyXyHGlww2uQHEygkK1ZhI9QAm+/CxSS+gfK5uhG8NNM1
knlOZhYT2F5td0im+MWztwglxlIPP+K5orxyIRPy8UcIt+rcbGZg3J7ThIY6DCK3wdO+A/ynPn0s
Fd3vK9Sm/WnGlPDoyD7woUgHBPGsemyGnh46QomcN6FrIu7YW+xuqsT6cELQQG6lz7oYEi/VN0qo
D88oViDaQkZOjQTHGO+FL/BtsbWunwlCa5+s+YV0sYWTvmm4n0A0B0RY1sgCqInbH2q+k0SoGzQQ
b4l0VF7LGJaz654bAUO3Gk+SlQD57VMVX+PBSb4vISLBTvkC8L24SgIleoWipZ9RkAK/9f0l0XnA
xaS1WwZi2umfRY/wewh/Ey6uLJN29i9GXzvg6F3xD7Wb0VO/vFKHDMU4CgS6fG1T40J0zOkdhW0r
/GqR0STPS+sO3j2nf3jm5CIbrLMRkGlKJ41VTnOcaZVWIiTCWUK4fGE4vaE4BgQsOOEru25WF3qH
3iYsI8miZ/Fo5RhL3nE9AzpTl9jIfprbGt6cywuSJkNQskW6LE2rYZ4O7rEduoEnnJMd0lOhaieD
MyDpLIrfFKvMhq0cAppn2JFQtfvgv2ehwoKlOHZXvHy9tSLA/rdDZsvo38uAZ7lb0Ds7A71GrURP
IPqF3LOTTssHHWn7Wv19VnnZhN3rjksrRQbKkybdhDgAunUNJKQyN5ul9pc1iISVpIQyWxW/ceq9
Qgn06V3zt37fJ7UXtCOeqx5GSvF8BMdvkUBvI2X/XrZqkM10CgF5gCH3q34BUh26665lqQd4m6yt
eWUObnf57x/WD6yd+bQQ/3+tir9smiEE7OPib7oyz1UG+FA9f7qJudg/vdeGxGbOqb/hK8I6tHt8
aRKECQdSOuo8B1CmatDAFQGe8rjlPcCPjq5/Mtpg6HK5Ovb37n7sBvAdWjWgvN2gp4QiF4n7C/yx
1UNrQa+BGhQM/JzJMc0ZghjWqy0tMc1qS1mcS18x/Yj+Zl1dzdPoIfWqdNFFF3Okp3M5BfZSWrSd
QqczRHnLsZcVn9OfdCyTKf2Idc+DkAqddruy5PaQDD/Ggh/TZGjoXyo6tJ95k8S6j1bm/ytnhcyA
rpawf4Kmyo6vl6S78s/zxvVRZp8QdN5MpV1RmtwBLgIjrclfgHISOHCAaeA+BcuwOmJBaX3cNzcM
2YHUYzHE9MhgqxX44XZBYw8ftBkzIKaf0mz0ZEFFIjJ9rezgFxiTeMjWPS17JrIRlf49SLD+o4DF
+FYVjZRl1cWwSPSNyZ3bdEngRXHP3sMVPnxNm0iQYaN7g2J6PxYJ+3nayIrmTiDHHo3ZlHUn085N
jhuyIaocWOEm/z4PrbMT04pc+rV4lwP/XUkQDlpelW0TLJmDY2a+53XW6QQtd+7nR0/P80U27ZTn
8Uw0uO+VYiCfS4rD2c88vcQrkEClNWdYh/l0xLaXZ3FTTVgC7JlPEmHOrD8jki7C53jHiOP4EFEg
+2aFYJLdcLbc7srdm002q9vKD4cAI7luPxe/+Z1dpwQ2kqngrUaNlVbK0HeYHO8gyM1gYt0Ug+on
mU7Ciu4Rh+gdiCNmDPYAZXqdK2VTzAoz1wAoMRa6RjuS1KfaLwBkhbyEI7JtHjVHN0w5uM28RkyQ
GT/dwlW0cUPQ2mtIpEwIqb8T7fChWU89nOAmLyBZZxvQCYCHoHpOjFmculJLnKdOGCPnXW1A2UcK
QSAvJckG5KUmjH47LCdeLG5DS1JgPlD7zx3Alqbdw7SHnoIKMwV1lumHo63AIDMb1y724AiV0ao0
b1DpCvMm52IGvzbLiOiQeh/9XqO3I/A01PbKjC7iF8KjnJxVL8g+spIhSbMeF9vEmm1iZpNuRSYY
QVUX0Bv4qkrobfFlGZkpyn9rv4GywgKeMeSeHQfpDnL5cJ68EKCtpLLzeSp8vorUnZ1QduUY4NiI
4GKJb+yRU58bSZzk1JxZTwpHNhrZoQDnPDbnQBkpaPQXhf4QU7xP0Ng96WIPquXRLMe0SZwhDcoz
OpyzvMphJuiTavuTZm65AZC5JO9zjzpFQbn1crlVaUNQQ1V4zkUi2zVSUtH/UZY95IjKH59QwiLl
GU8e61Q7AauwaegRksjExCJVlWn+CZWCvER6gIInE8uIv0YwzmpWxIX1agrR5q/y/P7+41WZlzp3
9IVTrtYfEJDHSHaJgNxzb2vfFmXdLWAUkiuawcwrU9/Wr9mgeZ2H0Kc/FYaplExZynkfh5SI3/Yo
zkT+O/j7fe6m5pDclCOWu0/AXLCo1KZTNhDGKGLa8Lnh8hyX9ux9Jgf0yN30XT62YAUKkJ2iiK4c
Bg4YdNNrGR7pGOXBX/zsisUqFPCeICiqnJF+BXKVkV2+siYQY2+I+EX0uXX/0MVRIsJMfkTR1d9d
W2kUHYrBOpt34sMw37qnGrXmfK5UtYQ8I76OHNsPGBUUInK4BMRd8MpOl47stGWFukvDootn2Piu
QRn5dgfGpgs6yAwjZOLJNDvFmpQg/zvguB6gOmYfqb8MRCu3LGgR/9+v3OVi0yMsTHDBpLg4RN3h
fc6d9pMrcyq1AfwWluuUqyxpmionQ7dPJCGHYOkA2mEKPafUGjglxXmGvT8f+XnIVaTy56ygyfMm
QFibxhF63OQOGS+j2poBErDPYx9pQI0k3MzIqTx/yx8bT5n6Lgpo0LyMrphfBsITuQDqnJ2QZJgL
HVHVtLzb9IvOahp/XgSXJr9Y1IuU0ppD323UcwOW9JAwgPzON1JvwnpJqwjiEqXJHFFM0FHFljY/
xdhxnK2cm81mYj6brMTrt0cnIyCt63HqgNGSxrdUwgENo9GCD7oazZ83clNzHRUEleIskslB/hiC
NYEOOc/SzTaLxf1v+ERitB07iReR+5BvxsshZUh/+lfyArdSunZKDOFxKJWMLlF/LcCneyGqSYOi
YQ0GC6Xc8wbOZFLXC42+ZsDWpis/seRNvKgatO12vzxS2nCJuPtQqjU+JuY9/OLy1RsoU/zsoP78
+Kc5Qs7cQITg12xtl0SKEtqvAuY3737+85gdZ88oB5mNdKvq2vU45ohakaOmqRW3D0VPNXXLBO6e
GH2AVj9+NdG/U+OR5SC+ipalxWov/DyssDuyCOPnlxUtNy5Ac0AryMK0eNcc8rzJ2NCQWuuKslDv
ue/SuUP/i1gO2AipViKpi6evFjj+wABKXxCfwDVNT4WsONWERxeM3iGii1iw9VCeIiHcjUN6z5iu
JPDRre3Y2FPrwlCUbTP1ks7W11UUzT+/1U2t56PuF/kR/hhQdwxXgJLXdePleUS/+mO9qODb6dH/
ZYmei9erwM4IoLw9Z8zekI26vD1vvKfCy6rYv3xZnUv5ZeodsgmnzbdXySdStxXGGI/A2N3LaRqY
2Z4+TyUXFBG/+diFY+SWJm7tGg6AGv9sKN4a27bZ7aw0RdJ0xCmmdM2C2WBfgXJ9IuiOawaPXLoP
ESFjDRukEDhO0fBxLR42Ka+VxLKcrvsbMc8enjtfLof6JLKlfNxy4hykXw1faY6mvCfAr/qTFXJ4
MBt3oaKe5+kh0d6RZ6ZHAaUcpHB+Pd1bKTbcvFhkOErpd3fkHu6+Ja0YomhiJ0e0b6KfJvf1mHwR
zxs8ghg4CljI9U1mWIuiPVHsOdQgSkUkpSJl9dxFUxprvS7maqFJ020OQ3paavcuRawGwFq0UNpV
zkqFf0i/TUHQ0QredZNDSYnQbizkfYUWp+/xuBrioFLD4yBXH6ohb1UmojWMFrS7vYafutaEOwSJ
29Txo5WqsAYOKS+doDVXKBZQmNUhwNkRzeDNhRjPAVGslsnv/K+eKWt0hkfjPYE/tJ9dbglJZUwb
6ur1q3/oYLgvssjXOuJE+QcCK0Sdz2D/3FoLEq/JX1Fhpeq2KnArNPnrqwG+elKDe/NYiewuTtyk
9s6yxn2BT1aS+uleWfSh4UkD484jwfNxYuVsoqFny5aXlulZAuW6TuWhL/q/TTsgROYZC5uwLhZ0
Re7GpaRZNDlApM5nh5drlQO9+NdcnMmlt6BYZRlfyieBnCRUEBhVM8Po5M6yYGrSneAN4iyoiem6
c8KAD8Wgamibu4xewobVpnNeO1fuimNaOz/voUoULdTYyJlHV5uX9kx7kpOsWoNM48oaP6v8XcVq
wX7w1yAizAKnZwAR/R22I1y+50A1+A3ktIH0C9jqy8mbOnMm9yDHQ0R112gjK7IqdK3I7zR5zanh
VGwqiT6E/FBn1wHLiQecmznfkb5StKYwzt4vsmLxIkGnRFICk/Hmd/lPYXWyREQgYDQJMtyCo11a
l/7WgcGDXWCksWII9wr14HmpcM6z6ddg6QYsiItLmYpF8aQfRCwJEgX1IZxXVueAoBs969RFmt5s
PCYQOy3coUAFLVadxG+7VOJg91B3glV1u0YW/JLNue4hWi2TIgI4uP/4vzFrim3xesjYfmjmMC7A
HJl4EwLHym2r5FHyJbwez6qUY8IETpWV/VYGLZrgBzb7YNZkQ5lrfIqkh+H3nwNk83NtEuzUyiwc
NCdyy2oD+rQW8LGcUprJN1ErZhsVUpSAIspo8c7nvd+ThF91Hg663IAiC/t6975FFjkA0COfxSOO
H4NYjDL/veUegz65zkX7vj9Jc+0+NLAqQIBanUiZc2ncnlN2se0avLrnI14ee1vmRwZQjpw6u5Ih
/69XLTNBBUo8gXm4G6ALmfajjIR2H2SKBmKxsgSHxtKlnu+2gXnkByplRgSvpdTDiCGKZ9StFnbX
DaCb6HPPfeRgUw76BpHyC2gEfV/groeEAcEYnGbC7AlFc8I+b26vblFlk2LBR9c4v66ok/ivYsy0
/Tq9l2pZ4tmRSPegrb3iLzgFraka6NyuxgoFivTijNubZ9O6E9Q1I0B9VSryp/pUVb5l5fWIsLwk
ExAVzTkuO3vbcxwKRXBXG3u3H2QFdXeQp60UTtDpLYsJJ+Ftjv0//saLPOwy/dZ0rY/Jd4P29tLg
3rD7YXvGcWEp0JVq6C0LYsd7N3FvlFhP6aim3Legv2xxZLPohIxjb/Ec6irdaJ2Zb/QiPz6bGTAd
znr2vpldPxubsT6FcZ4bw1EHvUf8JhMs8EikszWD/4/8xDUKX5GtehmT0SVphwLD1uLuRp75LkiU
jAScx5fh3i7PJu76IGQO5q2cAC0h9iKkXW3GgUkpEamWvTAh+NTcvpGTHA8VEjW2LIEnkDu/WDKS
Kr6EG2OL53VAxsMY392TvIuvSWKWJLCsV3E97LSOKp3R0YS8mdaX0WKatU237QXR5DQ8NuAjQPoV
uATQXswbA7rbkt20JdL4H1mAdhTKFUBO7wkbEHZMlPb77c0Mr0ZWplR7Ovg6mf64Ms2a4zXTMV0W
QfYUuB4/pC5hysV571LnhUC9VJv4N+VUI8IXWFVjFwLbRgIq1TWiPLZIi3feXqyvNw3pAW5O06Q5
QaKn2t6FqPCQY8aSGuQsQJudglC1i4duB3Jfo65qNcUspqLXzAw2lH7eHz7e4FWU1qR0qG4KJO8+
bWdAmcHWCwpQBP2g8f1e+icrpasDbTHi8H+5woNMM0t90atNpBVZI/fSZKj1y1J1e12EbC0uf2uc
hqZ48LA5bPRfOh3vHaz8DJIzNQ2KHYj8D78TjlBpyXJ7rzsxZzfYhfg7iim07QhLPwgNO4D0nKBf
5I1Rh/7TjQFLqsIN23Tdw3CBFvSeecXMiavUv1FOEHt0J8pbbWwLDb6D1xCvGvTnd3Jb/UFR0qXl
KNJhEFUgt4gPnPOfKSTA8YC2/vH+9tDhVXgc61M4oXULiCUW5jz9XDHcd+ruzG0pIqYFE+4hgowJ
X21Ju2aB7Yhto4TcnnE3xW0vBr+e9aUg2Y2//0W3nCzcuPFmvqexDe6GakfFx2V39P0wY2uIWR3E
SGiDmAIb157mD5C+RYvmnBW5lPBqc6O8lQg38fQQf0VXYVOAqHtJ1ERLRR1wcNhD8npp5rlg7K5v
+yjWHi6DL5VHS3HGHCiQK/J2amkjz6UJs+aY4I3TKd/WIMiD6F9b8/JKT/uX2L06ojES8oiBGRR+
9raVyjMueNijdfwxNDBiP1ch63FigEjpaP5ajAG3aBL2nmHyJ7BViZWIgksk5Qu7UduNWtpOcKFw
YO3gGhwy09c11Fb9E/466nD/Vpeqbxjt8DMo5e8d07wuZqD/Y8pmOJ2mC2bYdZpxFTMPFrFkW41F
5Lds8UyGMFrJ4R6wHa20wD2Ni7nIixAKSlt2FI3DMhIb6VUqbHK2d9o+rdV6PhfmtKTdOXh6Il9w
grndAHanSjZRF+4lTp511Zl77q5cDI28LoxTBOBsrFWRS88I0DQ/Mv6TtCfxVTGKYWcdYIWiGpef
oAm2N1d+F8KieOmm2AhTAtd4+ymPD4n4R6hLJ5UcgneP0MHMP8x7zXSvtuaIpOoCUBRe7Zypokyr
jzz7kEWkkbIT5XQSw9JNKGMdtLY115lzq2BMh7LPeiVn1Vg9ncYKEME0BN0PLYFW5VXHudP/UaUI
4tWjSgB9sV9M/pLpR9yoL/PvoTB+UVFN3Pd50KGxVNr2T5vepd7R5rn8pJ8XmJxywe9sfPiK1Ftc
mhuImOwqygp13Ifju7P7Kfs98qhB1NdWkxbksqedhGN5pkOlT0QvaQGFKBP41GtshNsZzM0gvcLt
8LxTZ8pH/1PyBnsESQsLWKvPBHofWpwuRbN7J40QCUvmITcqlJATg7qnzvduWFqNbp7DtILMzCdv
f0E9RS6TmZhNjxq76Z/QcXHGKhL910JeyUEQF8o9Je8ridqyij7YdoTD5xO8EpP1CRKWXCMrS4BW
JZv5UPZMnFTkKds8vQzYueRnoMjKxlwoDtGgMcB3dA4RLYZsGKTZzsYedmVYWvizMJ84zDvyYepX
Njeu8TySp4deNPZ0qcm3NAjNw8awQk4cG7n2mcRZA8pTR/WwG+TKhTdJCxtofKqo5s81nlKVDeoQ
/M2+UV4MoHppVVJBy0+YHAH5G4WS3IGSjoSQfcixVhEJsI3AdZNxvSJAXrq+ieIIA2uScEPr1pbx
yO7zbDBq22JV3HMKR/dxY7SyE4radibpJYhCkUQwWlF4ljGEKIiDPyIN94LK0Y5EInD7H+G3I60Z
a0I+QRL82GFroj1I/ajEOlWpeJmmIzt2ou7gloWpCTuKQmny+Lc8FSTBF687tN7f3aoYpCpYUW//
XI2/6zi0frPiox8GIili0obuNNiMvo8oK1HsJxpnbBWvCDg9mRNthh4kGKD3cj1fWAwFqPBEaE9I
u+AeY+LEmtPK0vV5DwzlB8SbigdynhViGsASbsabSM2+B8FrJjX5yLMc/ihBOWVp77lwSjV4q3n+
s7Fon0Q5FKEQdvMXqticGsF5EAf2ETFMip2LovmbODtyhCbNWraNAb2EO58sfDrHWTHw7iB59pd7
41r+9lBRNW704TqU3BGoC9qOAk9SgbAlB5LPAhA4S2hUpUybRnwVPJcf3ICUzitgAjDYo4rZw/z7
G6m5iahUV0eP53+JqvGvNTpES6uVnl62xkgct6q66/pXp7KhoWxaT/0Yqg9eNHwgi38HlBCJlX7m
wMCxQS4sXEUCyibd/xnWr1y93iEFdtL+NlUuFOrlySex0qmCjgkJNgu5RSpfsO/ZokR1Feyn74S3
PCRWroHGjXdj46Yx3bpFc+gzQYl1Jei4Bsd8VN8Bg6Wrhhe53RDiYyg3to4Dw34MoyEEPy4GJ1dC
R82g86puRKcJeiXUxr4drPFvK1zVgSYjumKmSHUw9k2tIVlCC87XLVS/Xn5aWFZPqlOy0OFdHaGm
Qu4002ucvlVrD1bKOepwLk2gRXnrzfJXSGWc6t8Bek0VYbnrpT4pfsqProHntTCEoQLylAIVB2fM
Xu8cGF77VyBLBNh/rq+M8hTzeLkQuO5his+6d5SMQl7E8wxOrF8fmOznTlPcmEg/xHiNG8atoK4a
a5YtG3n8VWq5nUbc+wwqp5MjSWxW05MaGYW/0mghttbcffHLYVHsnmdWn8cSNMCmahe0tWVmBlHI
kT/8vCPE7u6rB/5FPpJ+n2aVtWaEojE7mD7oPkixfNUV3xsx8Ctt82V+HiCUjCIIllyGMkpHgKyq
jqLn52NgAj+rA5xwJnV8pwsT/LLBAOa/Agd9MLdLi4uNPXLPSTLzkxiGGXzPwSWFVI3TEDXjUBZa
PrOLTQ4jqLwgSvi7PcU1FiE1pogrhzwqnak90OUGm2Afkvub9fy8qdkRRbv3O4bHCJ4daxmahT3d
R60e5dMS2Y3CD6NwSH7A5pciLEGA7jNNDbDQB48SBsRHph2WC3mC2hxhsyABdyWia8bXg4nIv22z
8VQ2mv5JNLxn28H4Kb2IR57fIwQoxA4cUUn8PIylt0aXNXu8y0aurCiu3InUyGdTiO2/qPC1gqWy
LgZFnvVCMLzweru9nEJIXt0Lsq1qsp2n5plLA7GABGQnHFrAHTJ3eoyO/1rUshIHUh+1mKtjNmy+
kqVpcZu0909VBz72B2D8lIsiDt2JkUFzbn3/NwoLxXUxULXCR5Wl889oBWzGOAkMUsfPBgQiPA/j
kZ4cEfF5NtGvzP4K9lrnFN/9d6XzXd3gDsim22gb1SilgBrEiD781N8pgVQhBZGJE/YqAoc0xHzu
GHb+QOCJxHEwjmq1PNgr313vhbjIyfm+m0eYCiaZVKfApf8UiS2LzelRnYiH/gacAI27/d7gg436
22WHz6D4r6uEloAK0LsGxhrUK2IgBxNmEoxxiM+5ICNth4rCDxKWb8Gw0rDht5sBxEvq8FXGVZIu
w4v1kWjZhKYIirDyHGB3cOK0ZURVd9uoLnjb+Wv4c3Wicj52/D4aGhe/uCkENBPImV5fqNav1IdH
Bxd55je9hlPKD/EOqSLr4YykLW+jtNWlnQA/qdD1p7s/d6H1lAoFPVQJu6RB/Yz/2GmCEgrF4lrn
eXmuaPZuEAnuj0/BrfchpllfpVcAeWB/vqKmeeOQI3tSVcxqG7j7vSZzer7WDNwyHarCo6kZXOOC
RmYcthSUTwQ04W3agfyplZvv2JG6izyOpCJWVT5/ENkFsrI4c3b3MEIiN/SHEtprDKVEdD8RIT9F
Lns8OVPgxRipcnUOwotWg1UpeRSFsO1pZDBpeVZ6CNxVupmL5Oi0vJDSi7cDow+snHvdeinYljGv
h2KD4W5oKNPC7MINhK9N4X8m3YUz19CGS8ucNv+xRZzP36Z2kfjyzv6Aq9Hh2DHpqpbHUuzJFqYj
YU5VCIoBLPd176ycvTKPG54TmOvqrnPUq0fOVfl+v2zbnzTBY9+MIt1xbQ2accNtkKrd8D0glApz
/kMki6EEm7lin2MedqARczDCKz5ALvD1iJqZg6qNlnJdQUVxXU1jGagzhVTnr3pWtCGgDWlSM8Gk
QMXiaj4BsIr66zIvXqeskueBLdgbDJH918giuEzVneWejX/paKteLPClMTByt4nxorrQMTKwMtRK
Q0tPKo9PYqd9hqsnTxjOt66rkjKgEKkHmartFK2rOQyIm+j3lMa6gfa7FkQgxIlHQQuVUgducU05
F227VPQzyZLjPwn2jx7Rc8xy6HjSczJX0UoAHwmZYPK48MTyvWMWi970MaU1h/E+hLJFahXbIFl5
aE+7Lk3ZpvjniWdl00Zt/721dc9lmkAHQRrVNtMrTm6xf+AawQxL8UWGtVL3NzwWSjXVIJa8f9Bo
gzKzz+VY3PB4TNBTmgL2ilcgsJlJERNIiW2LLOS4FDQ09JYXJjOVlCOI8MW7v8Es8OekPF3LMnFK
MFj6DgPLtY7Ys72yghNn/OphrnVymJOQbqitCEM+DcLQXFHsJ23sUyJVN7s0Dc8nmdmiUEgoq87E
Ev45h95KWF75C/unHZv+KHlX98oFaPYlhzKfZpSf/gzPbWtRPbJNVcrJ5hojczFSqNSIZYqorh0b
Qv1magNGIY+HwguTp+rh9JOqU06Q5oZ1vDJrhDhcTGx5Z8TRl/oK2QjV+eu+eHFpFS2pjuVQ4cyc
WTssSaxyk/zBF6+JZAeQtfV1mRTRG2bnfSoyl1xZgiVn6dktTADgR2iAwcKXUw4sKWMM0dEHtR/L
ckD8LqXM2zwzy1jneF3byPVnyy8t67HwH02mvWHt+LsTsJeiEJ9JDrkqhzKSCtQU9b8UR3xUdDot
SeX29JKYHK3lGJgy8/6G5vFH4TjYTrNjH2OP4//ENldvbkqTEEqjX7wE88y9vdcnMfDLU+GJmvPU
zhXonrGquSK/NFlaKieeMAxhQCRrw5B1Xu8f8fv59Tp8ePl68QCzkWQ6gBcp9dGsYSlzhTYUgLU1
JBrI4Z4IgMBAuvE3UugDo7ICz0oJwLi0hP0jctBJs6Vnjjkiw37nd4mhG1V8DcXXcZr5T7/a69tH
p6idDt71JECeDBVlDQACsOAO3+HfhtU4wsUI5fCBCTLf26RSKXvG78rr2PJCN986mKj/mI52qCT6
OwxnO6hstUJbDiUGXghu6/Es2poxPXjh1wUSHZid4JPYemCq1LmVGi2xkCSOE2/w6JRz58DwyaWn
JlbSgh/qxYharOpyz5d2wBd1hciG6hQIjTs/7qMgSAvZ4JJlP5pKEryMZseOFOTg5nFtDT+G0vna
SRfgOZRLba91DgZpfQysogZKB6FiUrU1BxSwd8+JJ7H6FoGf05ZjnuOkuThjm1UCW3PtoqE1z0mE
3VbCa/aENw95o1ktol3Y8NEGiSCliyL6sDJro/Sn3cL5TrLER0z/QYLQnqujAgwPVK7oAcWOxlZP
ntydPAeQ+AFlS/E1yznh8PqZcAuHg/+IWASG3edDekWYRbouca8P3ppwAt/dCDdu8lYlYYA30Tp/
UnB/ooIH7i0XFRnNC0THMqrahR3CRzgRM4q+9dkX6VlHUZfZknCNqEzrZhETBrkfWZRazPumKdXO
8+Xl/g9QjfS0XND+ZdgWSzrT4DzYTRdd16FCJI04t3QRHc+FaJR1FOM2BoFuvg/xRM0lAXWrEyGL
Tm7C8+tRPn+W4bJmyuAGk4Qh3dZcA3rEa1rIdVetfiezRSKrA33s/nqNv9vB+PBZppEM82fAwfhw
MsuCJxwKHFVDjIL0uuu1/zPY9wbfDzsoigrEuxScBbXkHcv4Tj2B0gurvk2nkATWL6JfH7tS8LV1
RSnLrKYpOE2VgC8sJh2jMwkY30bkFjXKRJYtSZRz9nWTGvtIFMVjfRV2APi9WeuXVs15oFD+9rRj
jNUeab33I3Gc7Yg9b85Qm6za9Jz8koVTzbuWe9kxXgI0jhrUkGhv5cW+PY2aja85G+8VMNZevQr8
kN1LszMBlmhmm630RV1bDvte3mpBpJc03YC1lL/ofH45pS10JeT96qyAEm20az8LEBMJQghR+4rH
kNribIyPRDaTS/FmapfWU7SLh9Y5a7p05mtd7EYsE93MWISWBLJpx4kL2sB8cNdPd/BK82swuU2y
Ag1tl6xTOMWkoN0PzjiQNgMO1lk6571rxc4L+VgqA9U7XaARGUywC2Q0w6Yb/KHB+e8zMYHuk//H
xgfkW2G1o3V3rIJKabPxA3WoFHRvUphHpY1bZdXumhvM8eQd/IYXke5uR02Q+qFpIWXTimWY921m
erelq8OgSvOoB3Tae3kjiX3QGxry/uhO3rpSeSKbeXnAqnZoYvhTYG6+/bzRMse5gkE4YgrtFWmH
X0ub75M8PM53/frFFsBewZ3C3yU94tOWNw2I/S8IEhrjZrMMqx96xniKtet9ylrb6/5V1/FEwYEp
AkZH6cePFFJT9VEDntCkIchA8VN+egsbKj7nvW1GzgObYyjmQxFCrE0ksQrDk1wH6mLLGBwybvkS
yLa+Zb4kdBhE4y1cRxUoP/9fd/63bj6k7FGoJNf4FjPJ6qxZOK3ERPeqQL+2bZkpzmZ/5EKkatDB
7nGisDf07hDY7hU7FlKoJoXJ9+nwKsuPyICJnj128xxJsulkavWT+67MBRnu4BZA2JZbJRFyK3el
pziOtoKykOfhoPVQdaNTOnS4KVcXNZiIktMND697Z7ZdiLt2gtXxY1LWpBirbJHV/bCFshGx4ZNJ
Q523hiltcZQIcblIekq+I7VnKTapm/sLeMzEu5cnIT7ctj4Pe3g1dhwA+42DWySJYPrh+6HJVsKC
pJ1ZhGAFSW1flEjCru8To7SCmc0Keh0vylQQXbM4oUI0evKCK9dILxt2s/AZlCGaCdpsF9UsWM+A
OcQZ4xuK3czqIiQdPn8YSIsszXPptDvdguc28J1Nw5YfpGfPrAYaa1aEY8B8SeSQFp+myiyEdkyH
0plUFR2lzJdiUth6AjeZ90c1U04k3LlFCYEzVcloda1qgiKwrasVM8BruiZn/PJD4suKIigc2/d9
yV0RhyIlO1VV0UVgynwTlqC2CECQN//fkiQS/IhuzhxR4m1umEoMNaY0QHCeENRqQOz/EI3IIe/i
rc4QiVdtq7csAbPVXHTsTFLAK+TZyYJioguEFtwaK696roSzqqSBDMgX3E9sbAiT3vaG8pPcBWKN
VayqDhwQD7OWR5qZeHaKaZYoDI8EJp+3i2XWkxMAYnN891QOhJ7kmjMlA795xG3/JFTDAvw2M5tW
yv5u37ieAo1bXjq9qJ8JW69qfzIRQrJlKlktKp+vsaz1m4/zYmuUbABYE3NzvBmL2ZYg3U+ckd0b
6I+4SXvRVS6gA1WvA6+BID3xvSRKILz8edRQ+yMwwxgOJEx8kxcJwNjWDzz5UQA8tbtCqnzY2kmL
vA+Yw0gugkCHWo6Fw+J7uTqhFTUsO6rq9tG6s+Tqqll/xvAMpNyK0RPzRHHjZ4asPq96PyPSNYdr
i8dNto+HlU8RI79RYZxXvGSvADZoW3PsDPeGXbeXcunMEtP+tHCFdbgJSZjHLWvt3SyInN+ttaY/
ktuvUeIrvBes5Kwqp4eraqZ7SnRw/67en1yONQsjehGVC2qv23cqeWXWa+LWK6lRd1vfpJWKuf71
PV89e13qFjKZIUfu/v9NC45//LCJBSaiNCVGU8v7mCgMhi+fYhjIqKdjDZm8fvzNcmt3vSi3SINz
RZd00o9rpRWhmFrjkSoOPXLjfSVjFsYQ19BsJX2+JH/nnXyPueE3tgG4XqUaGXekPIeuKabNqX4+
Ybp4ISaoxBv4wi7YPsZwjaGlKSnDHN52mWT1NhuR2igCqyjneC6vIdWQUqySpQYV2KSIK0sHl8Hs
fiUDL7jqqFvWAOvOw9NIA4rqLpv5uW8PQcrEXSxOpO5pDDr/685jJ6uO2/TPgLueGyUrPy0WK+/E
sWVQYMzU4DG/LjokjTYcl1a5AjpIvL0tZf6bC1aE6Sl7LgPtWsz+59TPxDFryZYbWknNyh2kxWqj
0dczcz9mLlJdfcw637ApjzYLhBji1l+DjLkTNTeVwgUSJ+Y1BLfRsEvtDCuYusKCCwXG0pyMvHib
miG9GZZHB9FzXPsmms9/XZRb8zKTxa2ztHodsLFhBd4YagCum5oWCaF2+yJt5SRTF6cF2IJ5Tmgg
fkAjZ1+g/yls464oHb71eVyFsb/IB5QfdLA5CAW4ebZ/jizw3ZdSiQhp0BDOKoV5W4wnsBQPb7k6
KnBZuVUN9k/+F097NKYMnOgvj9S3d97myBJyIShA/Ih+it4h07oKDMjJu1vQo0IICl91HN/5J+zM
a6N6DYl84LI82PvejAqz3qy8PJqBNa1l1Otd9gxNkKJiDceWR61eUqDxOmDy5Tha2p9T+JNGA0/7
XViE72Cd/KaRjTVQzRzO7BwKWp2AAcp4qGlrU8uyxvJGgXUbSj6UqZu5LGeDdUZpif0P+jDtmsr4
YUmM2QSRN3DVRtABV3gJDH8Cs7LOkFwigD9IeIxnSEMCfdLX6ba8WeoKctDM74ekz/DrNJOYWUxk
8HtnFYNO9j61gXO28zqn1sA0E411Fryi5CmUM3pxv7iC9C5WOl2ocN/UMWAYAhFaRpEVj+Ho+Bn4
jyRqAb6jCQ/XIbJn8qjKx5sIbmy3epQxMu4y5b97LftSpuS2l3j+O5l/gh59N+HA0C9wJ2oG4k4t
9kMKJJE/4r2IWPzP1WDu+fct0j0sLGfDRGmpzIVcWEvc4acQmZe0eGUGxwn1bz0dLPhwIUoPpwe6
ZaaMADwjHKWIJnnq0cTZ8byaOmGtJPMeaDqe+9RUhQ1iyfhIvS+ecXkGtLSuqm8TAQVS8kczMgh0
8CL9h8U+Y+Lfv2TUvfjjahbjZlfR0zLo+ouzwUhAEUriBmb19TP5JFRZBoxHdTDjDg3MkzXLCYld
N0csF9It59PonP6wdwWV8SH6eDJ7gjTl4csUgPe2qvD4nPEiTasw/9OlVU0o4zqx5VaHYiv5VNKt
lfWSZWZz0lKSaCGEG9GahUSISg9VQ42aO3SAtsCbTKXIKX6ailiie1dr9NAD3iIf9P0Coa0Zgy0v
NSB6kXANlyowiLA+m5UqIIlFxypjsToBM2K+Y6I7JkKnH7t6Ca53974K6Lv3AxIFjk/KusM8yc/H
gTeeamXC/AQmHSlTUdVxr7GOCFfOieUcp8TPXNWfcv9hifSASVPRBsLUvePLsVU+H68fAAXTa/vd
uim7IUTPBcVhTB7k6dMfDj/7eEI57ifIiFZOn20jO+Vwb25LqW0uxOqyGsekTQ1tHcKxcP0+mwW8
AtA6WFSyoh2QjREWsTVg3Cg2all+oYoZQKqZ6NghZ4QJR0x0+lG3KupK93AJ1iZJaFXTbEDHVMi0
mGFGdLbpF7UdG5aSN5Rc7BDFCsW4l8LT3VgFSRtrCIIxdoAbldcii9MhGKAxD7MfVoZ1mFLx8/x2
d4FmI5ryC7YnUc4MfAMjVFl4mw2M29LQTN/1a1G8289r31hNtPM6N9LHsSw/GlacprCpY/kEtz3n
E8Di4CRscMj1IFjEJRC53pOBpQaFpU6nJJF/fd8fJ/W4igGmYuN8BRiwLHzT0Bxc5avlccIghcN4
/RKF2TceXRvq1KZxFJebAD0HmOUVxEcjCQzt5VXv0K/oHDFoDDYr9qGSOoohp3XjvY9RUp8MQjvF
n/ssz+xACqMFYQnMtVuZ7sMjg5MP+cMFipA119WBIdxGKEYdQFZ+xaiy9KI4DAGXRh1QXhsBeJsv
Jyvs7kqWLNFT4W0WZlrgckzzbSJqW8WHFxJziWX2VmbpoMNWcNwF0Z+o8i/w8M756q6qO6U92sGF
l1LLjKUMQe0lLzedwrnwRy+sTovIkY1SN/z6+HuzY0g9n1vG1aGrThrMS6tgvq3pugjtg+AUjxMX
FsF64X+aOm8eF0YHrmaZCswKZzAZxv3pUAIKjyTWIZoGfQNZXGXBPWS3KnAchBT6a766FEwb5VAm
dXmNgQ8SE7ipYT8drI6j9/4QXrljh2jmVWtCfnz9o8qe8ehzqXf9EjmIX82syKzRqUL+AyA+atBa
fKrEDoVD8iodpFGPfGo/xL82BeDq63S1gTDwF6T1abn9zInR+6wQPkAKnJICY7nCaQTIKAUVNpvM
ZrEJDxVM7zvqVRXNOGb6aRpnjTR1fBd2D8MjRVBSFkXGTPCMe7fhqKFZxRIFs8dYJoVaN54xpr9+
Rvq25SSZWPgcvFunN27VqggBSm4poIR3JQXN4caQ9ZKfB715i+xZsZlb08tn755HtrIq0tT8kBwU
0VDciIk14EpUIPq25y38AsobiSVnTOaWGnznhGOWDrPcBXBCzDvgChF8x0DPnFomt2vVsRO/umWm
knGcmzCwYbFUvbsyyF6ozU6zeoCNFaKjxiWIf+bNzL87g6JYiQb2B5jqz86jwxrwUjNu5lOZh0cG
Hfwc7/r+HG1JI31rG2tbMikQO2TMWDIRO66I76EZU3ibHef0+Xh9aLqOjxOTjHZPs8q8cCFAY4c/
MpWNK0R3NJ7CBDWlS5ONbXMWPfkUb7P3wIGUfY20lrpuBs0abmikmr4oFMdjs1YLPfzh2JobAdnJ
S5z2Y1IxPpThdGK8v2wq6gCshpAVHdlN2vjF+3to/ncK28NVQIpTUxxL+RZp2q51er7qWNE+QUrF
SjqqYVxLTPdGiJsSUOxp1G1YIp3rETGY1Y/W3lTUAriugb0os0HgUfDOh+y2x6FNUq0o6AenUnYZ
hH829Dot1eWARGVVT6lhfEpRwHWt1szgz6BGnADaL2ZJRW1/MByaLhDWSkT04OvOp0TTCR/abM1N
eEZLkJ6JtoPiZbsKzcdsAK91fskQv1kR7k+npzB69mSEBYAl8NrFbBVYTQCv5RI/tTlcPIgfEtdr
vOKalTuZx1uxtRF/lxe6Buxgbade54OIrduRE9k15sOIqNc/KAUKUGLJXy9v08P17oC4c/RP+TpR
FVKMf7cgGSAK/nIKbf0pJKVJZ4ISYlVteX0kXtok41TrmxPJPIgMcfbJ/p3/VRFjlvMWX7Enp1o3
q36g6x0HF6eQwO6CvjWoHJ2JseQ6E5ppK7LCAjNqpAE5Lxo47kmUV1aM49+IbwkVeBLjBMMVhUV1
OS22IceRty4t3zpyqqWBch/YIEn9EmFy3H7yom9/NUJqUDS4Ab0+8SnYgWMGgCpiNnC3bR6FdRS4
KoaWBnXWYg5ECt7OBCA+2/duK0PZMI2JslzVeKP5YgE7u0HvhabFmtX6dMdTyVxCCqRwa6PeKhT/
TrFAPfhwdnr8tBPhNIbq73mhc3jL4LpHC95Q+Ywjflz2M3/WugMCSUj59t3pcI2D7dy58+HTqVUe
6l5DYAh6+//jfvhkKAwd2R909cc8dPG9ksd4gxHIDVpSSR5wyBEin/H2JMzwmIIXE1PntqHSOz6V
/pv6eAx6OGeuvS1Wk3SnBCV6et4gqD0SGYWKltFqqVBdFy9Jikgr1seFAFTDrCZfMxU+AbVVcsdu
BKVCOYNIJ3SiedSjqB50N2Gr410vfl0DUEPr89NFPXaGZWTdXKQzdSNsuYEIQHxYB0Fo7Mfvid2J
Hja5qlXjbGSEd3E5GkxH5Ye7e+s9FGFUzul3qD8Y6N7M4qT2hmpBtQ0ZcIzHDHvnv0mx0huufo99
ElpIiiZOvxHH9k6gZSQEASzDzB/DXSs9Z+JvX4G5ddr1kXo8mT+FHZeEgYS0bguNEJRYsbTVx7JT
Tzkz4F2zON7tGacFAY8ZCM5FzYp9ZiMmqDWgZi3Y+48S/N9YLTfNhlZl6WLHsfRwfeDJK5vsj9GB
8bP+m8bBtJ2ft+MvlzX9Otjc0KFO80w1ZmT2ftOzeatIy7QsgE/t1GkaSrbRFFXydnAqsFCeS5Ns
w8YCB+F6vPj3+oU+7sgJ18QQJD11CBmbDzJQ6BL0L07q7PfLmBYME82BjlnPSsL4M7lfowX063cU
+QLXYEZQlh0GUAocFNOCB1yTwiX+xRvjVnJ1OwlLJDgJ5eiKSPhbYT9vk550HU55Pvc9l43vovnf
mRg96Aecvjd/FHAnUhHDoDZUmYs5lQYFtFrXcY6/np/AxvaWbwWGC9d6C+RCd0rFBZIfPDPSe1/E
DwwfCHJgDvTr2qdmeQ2WaFAgSFpCLvkMTwqUMQCyR5nbIXcBYDrHhYKJiObZdxgUum1U8M6hj5ra
zGg0hfVyevQYO7Nl2luCKL4bkgry5fgO0AtnAdsP5xHOQDJZeRZ0kvgVKuFqnkGvk5kFpBi+edwc
AZR9OisIUB89NDcdJiYfqvBSGtC0PN5gmoeN4OI2w77/YW7YKzS8RzsviJEMdEsNTqCmKQswxjIk
/guzZ8qyhQclQQxQiJIqKUsbOOgxEsKMPR8mpq7bt2phhUK/A9Jj0zGcmPwez0q1+htVs7K4b2hp
Ae0RKHG/ZDt4VFNYh6OzunkquVprqZVmfd8IWgt28EFe9+1pEp/fwsKc0r0xNpv45RoKxQSgBolz
Q6UHinl1dXDIeEfIucAwy8Bp32gcVB//4NXzuvAY97nOqYzbzqOpDSWD32QALKDMktWeL+zkInt9
IXx96Ky27EnlIWOeXAEXai/Xsat3VDea79+EyvGTkIkmzucJ7GiHWZB2D0hDxz1HOBBT59phX/g1
FhZH/XFisqw9Ug7oaQiJjGKOXJPLuAS+kwrwmjHDrDjuojoXEkNX2zbMs0AJVlDy5oQ0tsPHcsox
pXJIFNrRMbSKUz3fFkTvpv9UCVhKz5/tCTODLOJgdm+JCiL8QthHsBeHE19pG7/kxKre7w/1IrGM
aE/tVCfUGZUprMIIgnfqT/W+hiVCfKNy1IaWF0XF62QdtIpsI8NREHAvSl/9ah0OAODcJLbYZ771
+khT0sq/ysx+8xDUZ1cMFyubvGIvmEaDUwW28ocy6/e6D6BXQbbu9fnkWv1kAcQwAqzC83XjpaZw
/R17jUz+1IbJzmzv5/hbaRNN6wuVJo1l1G8j2Gl4R89CZ1URVHzbtSp+h64RuTIwrK+ChUUfPJ7V
rNg5FlQmaVGEPAwSW6UkumCyvJu7KOFVxPQtyXrsVt5hNmYWZIvEgDVKPpa8oRbp2O0VAd3jffsX
AI3wLqZ9W+wE/BGPotTx9lYEIGBJqoUuytKGk1fAowdI7Rg75sAr7FZc54MDGX/pHujTDzSqnjgP
v3l+jwF3GPy2VK8A1uKmEKiz3Ii8FgQzrNjX8I0YordVZi/ao38vHGcNKSLWk5/WLAJj/TOflrJ6
zEd/EyoNkohySs3uo53GhH6h7hRhrCtlTfUbuyXW4tYREJEG4fZt13VKoVguXCRKFu85xgDYBYOr
JvgyMaLttWlXuzZfZrz7a8Y8DuQtT27KFWlZuer9aXVSjXhH7ANSWaIF9q+eu/nqBXN2sB1CSeln
SE9r9BcRP/3MkGcutKoBPJjdYUiUPwHlu+SKwdoZD/5tuYN58LuKUvUeHIX9Q1dcLeGrsHhIyjbl
k1fNMLhA5N/bM4CVoA+arCpbOjYoXsr19eCRup6BVDCgVot1WlxUpqCVb43Qdv5oC3BxxLgUkb4I
rPR7VM3DiQfwyX2ytCrWZ5ki9sdBn7alKk/Mqtodb93MpHW6MrH9v9ncEV7OaPJaOb4slkv1Efsh
GTOk4ABRztQ9xY3Xpzfm/3HZ/0kxD9AHzqgX/Y9BWvytGjVx4vBo3n7sFypSgbD4aAwf0iZ3CcaR
hI37IpKoufPjpL4gOB2pDSkqXwuM4fx/8SbERDYPvHkXeHOtyc5Luu1FhyWm32JEQ/xhwhDcC5SJ
DudHcLcnbxmOVMMQAxC0jw58wScnfaDgyCqrWw9Eu6Ys3qjwzhSbE3wUlfjyDC+3gM6o1TExp7OJ
iDhMb0oau0omVfKG9IrmUSeZzaKbwqfI01Uad3jq5QAXAiJ7147DCNpxsa24jvr7UIpAr5jynjo1
XurfmI3gPx04huoafmzOFteSnNJQ+Ctuty8EBM0t7Kjkk/akRHhWzuD6ZEZGAdANmziRt46IwViQ
HsisOgr00r5wmW11yV4bTvqZmVndowRMtS/kVGPDYalhC1oZhdQjZltzz07jtFSkiLeYnFF729Iw
393OM2o+xnajz3O7U9G/H/HSeQrEjx5LmNjk3l826CgB0O/4Q9cXXkY6BJmECW8uG4hQ8kjSmK1r
t0KgnwW4MNHq8xwUD5bkp4iRTej3qejhKvzRPC4fM0D20BmvRFY/RP//SA4Uqhzmwb5JDPslNcMx
+sogvOAfej8RJ4tzbbm+ypAqkKneP1a4KqgshDBLP0M9sqvze3j3QVdxoUSVlvuzf3786hobJIWD
Ar0oHfVrcbb19JEPUlMeC8amCCyPM2gnkjoCY8wV62phlj4hA95mRO80bv4XESfBBBFITQkTMdA6
8TYfjgkyC5nw8UnIzzTCmdu9jId086gjZj40HhTixXmxruLyfHFq4JewP4WZxwaUiiniN2Hc1FcJ
WQZLEJ66fyGuPm7kok/Ob2aHDkUJGp6NNRu1ey+NpKaHwiygre6EsCE/ZRUuC90Z7yeFVQfhrmJ8
zDokYvSRmKbyGQlIC1P6RXnLYYfmOLcurOati0M3nIeTT3V4dFVH6FXN/ekbyLuP5udJFKzzRYgC
6zx9+ME9czqoIlt4xmjxtOzMWh6dzjl14suYt4KSruNmbBrzxvL9iwzyWe5dILIVYnoWr/YO/8pb
KTkgrjs5WByN7RikW/PYSdF+hr4/2VB/vZuZ9eCFQv2hjZqD/U5tMO9YNTmG4AQvy+XkfJrZ1PBf
TFbIaHEqQBaggwl6J6qJYLsl/vJ2qwXEyt7cv1nqbQeX7IVbDEFmAPsG3tATvS5DQIW28ZCe122e
TxcJOpewUUopICWzVl+oW97bAGnp0BN0zBlZu1aQ3Npj3WaN+iyt3ME0rYRnlr+vXVqM8lfjRVJQ
y1EkbVcGUjkmgtMFzKFmddAP26j+HAX89qk0CweZvfCj8UfWQC1Fr6ZumlOAXLKrnn9EpoDYk+c3
F/ie0jk3viiL7KWoN5OebtS6XoGEa/mvUtlU0AyHhKEPy08LU3M3jXbt+Q8anWxFwomQNRLhimc/
ii6eO0EkrEcRjYmWrBQoaQMkYqmdU8dF4a6NEiQ3LKo3+6AUEwFsua768UEKQBZk62aQOJ/TaUe3
U+24tiGjfuh/94jzo/fINXQcVYaAlH1ETVd1xXHZ0MGH2Q21C2YFWqV9JsvsP3kTx9wLcmuvYCeX
QgcORKrEJAs+vAvtJAdPkSnGKizETmHibyg8SwKi6s/O2FZEIXzskScHuza6Sy6LGIRsdXQqCI2s
4BV7BtYc1GUBkJdG2aGWK7my9gaqpY6axBG/EhxMarSveSUSlkNP6CMQunaaDnDUC5a++prBBToz
twF9LXBQQ2x3F3+OnXwP8U8rtiTM61EslCMpnaRpH8/tS6rC/wA/wvuXII0wFive+2kSKbfkoCY2
VxsbGp4VM1b7iYYySvacNe0BzQPLbfFVeHuXSTB8Yo5fBsXf1clNAMwXttnYA7lMpZJchk95aKf/
UbwmYECWd21RSjFT0gbM+6Mg+NrgwU8cUS3T5UroAxMyfV5yIWpyyknmIDcjPmv/QkCq82R8Ksca
MN0A/QanxO50HwxIxhr6cJ/TiKLKk4ybB6QmRLr19dS+uwUypLkZcSr9nIn/L1L68Wn9dUG5JrlO
PmTLojVtTJfOEuytsRXZzRaBoWzFeONgavTo5lBZcxfG6dBY7SZGWw8u5BjsiCQmFRzpcEWlccUY
D6VT9/+x8WSjcnmGWBnEgSV6pvsW4Ae/tW3fta/xVXTY6C+pRHJRx8hxIdKXH9yTqjiCDzavfYCB
KhlHGKx7WUQfXzfp8vo8U1FjSjnB70rqjN+u7vT9jeFax9WYW1cxoheZ9l47KEOgU6s4ToMUBcIK
/LKn64EKASoV/MC4Mzl+urQ2QqRce5zWU0zpumnxUtBNKiI77HqVt6Y+s28rUN2mhnqRfW18X/wd
+O9+YvItl5GZ3Y6tZHORqFef+ZfB52iYS+G0e5CeKpJO116lBzEfEdFK7NFGh1cK0RPatpovE2cn
u1Q3wSkTY5uUn+oKz4jIzP/LnGdaySjNjSVH2yOUTX7lSZMfQM5RVlC5xafQD2r4t2iR24WyHPUy
0byyi+/Utk7JchOwl60h3ZPRiBs44eMxP/M+q8cje9bWnqhMNQpYGjLN2RjoAdgcnQhkbGR+gr0J
Jf4xYFMBT38NGNPMFeUHthHQSsBWdOCoX4yIMYDK0njHDfZ4G2L+rdQjE6+REqPRSqtLgPxYe4uF
vX2pjU4qZkJntmDORzsccIu51jyFu9HqUTKisQdigEc0mXmuOmR7NwneuhptxQFz9czISVN54Tpo
mXawaHC1xriARbVdLDD9XoPbKWsMZOraktKF/7iIUPqjAl9boz8ub4oyt3jBN6up0FlW6tP3A+NW
nhsg/U3jTA/hCprkiAYGslRPr1QXsDXFNF2d5NW4kBwONF7LhdeLmsvxo5Ug6VMCwVTJXJmVqYmg
8D6TRj9zWgkyOxgI2r2drm3PHoopuzD/n93lr/XPfYU9HXNe3xtC/gWvg7xbC+PPDf59C3Gsl/Gb
y5AP8gCJtPLBn44euvVRLMx9PdahLASGo7EvFumhX1kjuPtqsoQHywl4U0Sp7k9f2cHAWokg1tL+
wwT+X5yyQtVybmvfoFnDJvP92rAtx1seAjG97e7HFyKzqpUR8zY1VLxC3YmIdxjlSSb64a/1rFvO
whGJH6ufLc9QskWaKXJde2hcSwBlEH+HJ/ZjoLRGqsAIev4n35hjN2eN6OxrOdEFHLeSWNSs9EyB
fEq0gy3BlrmF9+uu/x5nfkykc7IVaSkBXClTeJ65dupXJRlNvUHvuzQMFgy0Sd6amGPNkFPIO8A+
UOf+11PmxJdH75D0vcqhxr+itjt3iCWlkV3FIadVVzQ3rezIi0DgK8tgRmlPzF68PXt6E/ra67mw
j2luQhmx6CstG5X+SIVjFgfIyW6ExzepA/B+iu5/M0UXthFqkIu7iB2qlljc5Sxd1/SL1WAE2a79
D4smw3u9djnjh3l1kVwK8CqJSOXXaphYp0Kmz23ubLlqyoRIsKQpU7Cuaf5VIPB/lL71R/H5y5uV
kMOR1v3+dYRb+yi8pZSOvw3UVAhOcqKhjco12YiXO66npAZhHuSBqZpD893r03xNhoCGnh3cB3sF
mN0bIr/HPtJ+02d2hmPpbvtpij44boha87Di8ANnaJSQbKWG5OozdVSjXvPrQylpibe2DwODQiiE
LXTP8l762po38t45RQByJ1D31AG4+bui+ve5+Z9Th+ZgPTDjSnxELxN/ELcCB5bZyRT+0Q6WALtA
aeM5SP2FV7t3lh8u+sJMirFKyfFZ8qglo3cQ8sG/0q5rRcdNQlewo9JDH2Kmh/yLFt2B/zPksMYu
hwtnnxbRdFhlroDUDJJuxrFpeTWH+ZyqCYfQ8ZTkS89yON5SHKC4bVm8Y2R6bp4M78ZWGI5Aox1D
wFTt/TdiwqyYGl/f6NB9mWwo+tOqbAFt+/eyjYBFqzCxPdbts2g+Lf0mT6fH9/oD0PbhVtUS4hbP
MkhVyxhVKsP7KfpvJ8h12vTTwp2ENP2JpAo9elHC4GYkPvbmYH2ecIBjz06/OMsCJVsJSRwMxa02
gqqc2lR0+cx0dWmADV/bmar3sMyzL90XSI5tOQeYVf694vKcFpSFBX/VNkmXcMtBvlMqwdyXDQ42
SRbVwfl7n3FX4nDKXkXIJBohM7t3QnSPE00RYr0FXKyJlsUVCRqGBPbPv26yi1mgcE/3dNlbguU9
spHFbmNQ3mvGPPN0KjPwtWAFaj5Oasg0F2p93bIRfJCtUX9FJEJNjjpY6vZCOMVGaYPFFyZT7fH0
wamwDy29yPMWLeYhFt30JvBNxrcloqQjkfH1ciHYP/F/f/h6DNXSUTId7jiGUT+0VZe5mFetEQYJ
ZxpJiINs2fm8H1L4fJoftOJiNO3rFCoEedkHoXiX+tCu51KnzyEHQ+cpmodUFhjVUcZDuKW9Jo3o
93JuDof/hm4i8uglAeVupz/asH0KUPsuJUFZYirlqu1bfwgY+UbYqA5oA5/weWat0jey42aOU6zB
voOuOXtUZn8Jm+9Hpzn55tKbn8X+3v2uAAk5b8pOvjqJmw0WJlQzLeFkKqGDjr/R6rkQKxTFp2pI
7nOk6hZjLbxHsANSvZqXusqcKPbjEZTc9BtsPtdU3O4VxVUrti0ZyYc90VxifiUzu/EEq+hAPZkc
Avq14iNeUOxxKyGRkqAEAA75sP1I+VhgPgV2FnXT3oeMifQhT55YbOxnR45Y7RkeMzmnIVS8S4I+
orXaZNXa68q3yZA8NrYgicZzFJ/folved059KzzHi66eMClL/zdFF+Dn2MOD6Yp26jeR1lJVYxyL
VZuvBVAB5ttoWBSUU44i6qQ8Q7Tfz4xHruWhQJyglnCMl9szXk1N6QeNA0byZRRU8tF40/msI4mn
9rFQ/hwuZp/NkRHW9EYT3VyDh6+44QhB0QhBaZw6IP0CU79sfUvec1wDfCpLuh+Z16oj1+nVHlGP
v9AY+y1oIY1BwRp8BIc5DSCBXwSWeXwUUywnon+Bks9qWlRdZiZwSInPkL7nmge7B3vWOtDVxRxW
nwLcmpyHw5zaBU9b53UHOoVH6ph8iiA97l9B9nyvcq/bTzJmYRDrGt4Dch57CUivKtyWZleuZVPs
8meW0h8cG1uZv3N8rrJEUxrE64gYHJFvDpTMJmXisd6VQ86Whxdyw1izUJIRd3PkhievpDzcizqO
g7MSZaJajfgNHG+PTgJgmJjdsT/xu+7hgS9MDXctrfvDtolCCXVQBijf8LNy+wUYW/Cfx4p7HrGR
cmQXrCkKL77qZgW6jfOY6a9Suyrzr5TtRzdWJ/Fr/WTgCoA0UBVaffhFFWjCDWKcGpWtPqtkJ94O
Dy+U55dklxQFcN9sJvM/x+I7WtePthorvwWD68GW9xI3esuBzCwUM/4NmiXndE8ilg0LxmoVayQQ
atzgq2YSAKm7+wRolEqafwpWLQZwMF3X4dPz+6QvC9D7UA4ogps2lBIjpOq/DNXNQLFF4yQRgNoj
FavIDM4IdUMZF4axmdt8trDjQI5g/VLG54FtS4IkJbWa1IDS3rIJl63Mcd/tGL7UhOhIu4tVW3Rd
wzCDlGVVrhQ3bKnKQEbM4vfgxUeKLglh7kh9cxLPDi75CKqla0u1TO73qikIvMNRSMqGl4bYMLPz
s++L8CRs0go31+Z9zM639uvh/f6eiwFuWX7ZrqRCBgUYKhZdZmBdoss4tBs5JqlULDHVYVFm/lou
pr1qHTrEpJ+jZ1Ml3NwbC/vJUN9Oj8CLNqeP6ixAki4zbNOK+tRQm3mAkhQyrEfTaUkIqEPF4hu7
PaiAuXMPH0U00NXCPpVq9w0C/F45B7JRXJGb2d4dNQaZGJHMT8SN2KfgS2dlg189JWtwW/uYOAHj
apQagelTF+dDS6h/FhXdyEPdNdzabHWKiF1w8FRJl1UdztQOpiPExYjq3RTxT+g18fEATZPw9qFX
sA7uzjMvrhpUfshhuLAs3lVPHpNoTlBkTMja7UeNdTMB7zKK2cn2gN99PUlk/0Q1oTjf2mulRjM+
sxm3Rn2XDH6iI5LQXxDTLp/99/wrXiDiIQ6py5XJOV3SstBBXKmX66oOubKlB2eMTjzuaAFxAdgr
XZcQjEzh27lFbRZSSFRDD9v36G8SFmwHWryk+yDnH8eQf6NoFjgmNltCbkNsG/SPtFc7HgtuJteq
k4doeHC9Q062IVHMAl7XaqN9ISCwzTt65xFvvytjwJBtszXb0/niQCK+XoRe8rpk4q21YNgcO6Ty
N2OyQlr7nkx5iajdzq14W5NRc9nxOZPNyBgV9DIrIXm14yRHKLAi33NeE8MZP2WhkSrjvrBFqbk3
NkoVlLmxndN5GIWqv/JQHZYdQRcx337D6rH8/zDVeWiWGSqkUL2ioD407IHHNN026sMSIGZ9/47F
qHslkwW3LPx8O0XoGmnzkrb1QWoG3tFgOUfwKz1zlut4aM+QSREiYcDnIhYz8PZgi77RYTcv1qtd
XwRxF/tZiHs+8H51zATAjM5EYJYndi2k5Pg0LiA8mJk0ewHIwj+rUFKXVesKsSNl1i/fFcQUrZqH
Eru44tDgEX2Y/2yEsO/kYJLyPBCvywD24D5HjX3OkZ0KO4uZW5cegupI6Td1D57z4lqtTqMIhXRS
2tJiGHIx1tNTPs8/RLN8zD2swzzOku+wi1J6jx/PPnLirJm1gf4tjApaNv0UlPp+/4R1TI0/3C/3
ooCG1yzQKCBoTbC58c9ifxuOWeX72aPI78MZHwiySKCC9RMMfAy77Jw13xeDEUWDnq/TY01ikCHB
cNnBFR+Vxe1pVYvUnxqCd/XrArPEmygwF5rJKF/eEOnJ7ak18LI2afMTa+bt/ySa3a35YCKnTjtR
EGCfVuLJhPLEilRfKJAUuNmXTFVWXSEL9xtckkbPdUfQi8wEwol83ad4ZNSNXsmiQATfy5c6cSto
qPnKA6otbzX954DZTYFnzaWsVAd3FHujOWQYnKadPqtb/2KnIu/JLz2quMl25Yt/fCQ4y1GqQJwA
BmVjIzMvOQrRrYoxdVIb0THGk5gRnXk8qi0phkwYoNGsmUMe2m9VfYb/Ky3EBh/iW5z38Y3eR2Is
vLH2G91c2GtuB6iJE/rMGT/nVkt97Bqhyer6FD4wVd9nPRplWlL164JxvsWlixGIq74h7Omxj5nq
YTSykXpRZiZtm9FtZpoUWGylixMRxqYl7Yg28aRsP5Np52N1G1oRJ366ECS03kBtx7QAnnrabzOi
XqXgcV0HiAec4bJXP556cj6h8CdMD8kTD8jm21LzXRxb+MdQjWQwZvQAvWgzUm+bGhRx/g7DyDQ2
etXNDm7pOdA4g9EV64pDwMF5K05WYMSzEBUrE5qBIDOUINgOq7+oC285bRcOAkszqWu3Z6ZsQBba
tCUguTRoJeGkZCapuh0b9M98DPtZFUd1xnLf8Tk4lRLtl0cdSrG+lbIURrwdXexgFw6TegZbAksi
8IMVYzQmhpJVbIspIyWHNHELhvW+hGHQe8K/GVfzj9pfmqF5MvruAd2hXCcbDceNIjiTh1LhyD+H
l1bJzZY2cmYN0hPqBwGOREN7mX0mdOm4jHjQWpbjlzoDmJti5cCAaNTkWLa8F7GvP1IJCU7gs+xq
gtbbfQRWoTLYuqhw6e5VTt4arxRHAkcht3cvM/cxrGVXqYdunNn6LivUlH/JZUETjV+uPNWVSLsV
0WLkHDriMbU+8IZxaCzUIsAFKG3MROr28yfiW6Zl3/TP8FG6RnGtZ04x/36AOokUedbbi22X7tio
SL7iDvIp/XygHBJAV1BfUlLp35BynoSQEVeG150+aYPmXKoqKSY2lSx3PstG+ooGmwfbKGnYvEHH
OU0WZ5gAkmuFIV878n2o9WbSLYGzHh0GyNzTWjUvEaraNrwzGM3oCnwYG/CPKhThbeh6BG2iTkhX
YO1fx3ax6JnYhJ0Sx1J6jEHoc8X7cEqq6KFllk3arucm44DM57ROKZlYwEx2P6HQK51Hosuu7aK7
Mc8dVxikU6dRHx74xnHs+vPzRNRTz4U5UytSOTzWOL3l4tfrIT7/iTGzKRzt/fIIM0X4SoTXa0Wp
fpf+tTUcqXlabhKNVlnmzab3u+oNqqq8SRjCq6JyqzdDTjZMmR6zcxqC89U+98odRRpnn96h1Cvm
1vwPdqrkJrMhf3xiKBSqAfTKuBLMbW/sjTNFFPgpbBVrXRIVGNuyApDn/ajzA3p8xSCzcdbbCHqD
BgkhZDV95kb9K/URjYsUTxsi25TkEwzb5E2UBloWkQVtlj+y8xZEFhp9RcYMFeL+NXFTzLZ5GT5j
hh4L9mwMUwJEu5daXx9mI2qsT9JJlx36ZMjWUQyf7BnQMMS2MUIePNw01HI4mHRUsugNH/brYxlS
wr+EH/lAKcTrnSbA5ZSAlfHLh7UbtJBzKAGj0kglyc21tcDVPrUb1p9W+DoKwtcABge5K2k0Z6p2
qn41ZnoIkYghvPI26aNEssKg061hqFSWgJSPLW9U3ucuy35jpzFQlb0TJJyCmN5HrIGWdKbYgl3a
t0E+15/qn+rqQ7AnuZxdissaBMcyVP2bKj84wUvEHJEnFT1j1k7G2h7ZpGwz727MroziLVvHtzXe
/4RlwkjwVNK4hvQBy/OvMn42wQcwBW7wI4I/HfNT09yrWSpb5251Rd20Bsazj9jOzcy2ZEhIBOv7
5cFqmrTL37mj5BLyV3ZMm4kTR8Vwrj0qU9HF13g8shn78IyE7JIap4K6XO5xlDJVEzhYHjCQ9Pjv
elLL4UEOuAW4ikW8G2ZKUrWC0FfHG6fSHuvyvHe2YKRnjAC9uMzV621SYcb6lwBzDhUrcA0tU99p
/YdFtHsIFgHmiytTXQtzbH/cLIQJ56khe8Eao/WIxWmyWCcHEB/OkAhquxHOhF5L8CvWoKXUcsj6
PMAzgnTpmqkIf/DsUnB6pUhcnMc5bebNyp4ckOGrucEDxNqcP7s4ZwyJJZTbfS1Vy3f2LT0gOXhL
FeiDwpUNSTRlIQQSe1xJDvIVC0hElNwm/wyZ0gO4zUEMc6h3FKX4C++rfvFrdoc+c1uxpSJS9h1Z
DU7LriUhWfF8IvUvbMQkCtQZMN15rUKue6zuGEW+DX9LmXu2wKZJxzZIsJ8DggQtgvA0HJq+3mwm
1kkBAFViUh5cgUTcsxkvsbcZlh3PoET/rOdOkIyfhlFgYIu3ItOaXa6+J+0BN/WDdNkNgejZYpje
c66lafgV+jJvrRM1GhPOyR7WtRAFOFIZijDObg04kdhIwvnpOHawxGHThxTnY2WHHnJdqTw57dwT
LCTTvl8qHa+EBsGMIQIDevIp6gtcdpQG9fjkiWCZ3Dha/LDTZxOUIxunMdtRyYWPqm1p8fzNQyos
NYvBLY4NTb5x3Rca6C/BiA6OKwClNvo1EhK+FRsdmG+kqUAvq912ZzLPe7BSvugKq+fruFBIdD1y
M4nOl4XynNrJhtfJcadw3JRzPhRJCtzStdgfjOvY4KyegyHRYEuDc3OH66cFcwG7mVhuIcfPzmon
eMkUor65fQ7dqGwSKQCHHzPWqW5pRYC5ZVSy+4zkaOijlJnW5/KIH2gdVnQIM5GvCGmKNWrnPR/K
1grGzCP7Ii3dFfVCxVIZ6Gi7POTDiA1AoOJBFYShU+8jeE1vw1zuLXfV9oxNsMNlSV6gimKwIZt3
KRhgrdiVTCqfqDEo0hSEvPM5SJHWMFvZshspeJ19SGal0cE+hPRD66SyL1FD4VLHpsqU1xe0lLnu
EsPG6mpOyDvbuLmDNuIWp2rnqtzXxJ5pY+Q7I+qXOXcF11zX7Q+FbWTn6tgJkCLjFKQbJlVKKrfe
FcSH65rmhDGo1bjah+yI4SN+rBYufQF1xhGLmohPspmpO6jY0VILdyU33htHFHObPrdPes0aVWO6
covpeAvnHZ4rbv+42wf5v28MvUNaj8yvfu8oBk455zkIQBvbXaNjZfuEWCrBVrLJ8uH9GMHKuF20
sYkUqkP92jThTkU6BDqZSRv4okiuOjyw7p2Sgm6GGnNnvv4FWUzwUH6yQT3v4f3lhtCGZk8Yw9jT
971G0HBC9W731wk0lFB6lzDAuzQ6rQ7wOAp/x4eEPwZQj1+i/bx8hJsLK/igemZoVKVrNvP3WEln
i8vMHUXHggWV7ekUCNGbkX30hkeyLtMFKT9jpv+bQU2zZqoN2Vgtwqry9KxsVctRxq+38IHCxkHA
YjzxEtfSmPhunUaEpZcz5XnHWotDimDBDQ1Nrpx+yIzAP5/ebDVABfzsA0j2u9+tvssP9z9LdmIz
5D5MulmQDE+rdU3xa3TuTYSNOWWJdbG2tQpAD6i4SgHPHwvU8gB/VKfGv8cC6BOIkSSDMh4OfIJM
tZOGqVoNFm40+Ul/UTgmYGSHDog/FJKw56j9d/i/gyUI6GzWl0o7jpDMaxnGB0rOca/UkYdOYmpj
Prw+I4/DEs/OAbkhPotA1CRDOkZ/RAeUp7xMJJwlwYYFYVEu7I2t3h1f5qzqDWgjbcL6tBSpZ9De
1ShbvUMDToUJ2WgK0hcGhYh9f1vnAIHAfKlSWgciYsjzZ0vz+wnQikoHPdCOEvw/Aarq53L4bt8I
l+QGsJlgVtNskzUJPmjfYjVS7V4YyiSwGLOzibAMxrhBc3QNNDly3a3B4+CzQgWuDMd9ebWBHkhB
7n3eou+6RrW8kqbNz0/YIGkwMqAJDsBHYfszRJtUW9Zgov/sVeNQ80E4x7gVF0mp9rOo8yaW34Gv
8qGpbka5QE9iKkNEZBznJhKqSZXo9RkRHuUtJBrwu0N+FQDWJ4vDXHGU/1yMWmsmjMl7ABkvAxOO
zq6gs7NYJ5kwlHXThZuBIM4KjAcxgBgo8M5OK29xLkaz92jYusiEYcaOkwi4sdr4jzP2zRrnEBYA
2LhmLaxVk3SLSKnGXjVhSzACJF+MXCfFefhyhDbSSjv6F7LUrAwBJ6Sy0jfAK58XoRVR/wTErNI1
TBNpjFOOS6qi9ocq+rkmJlYNP68g9Y6jAmigyNK0vf3Z8yD98XydvrADj1m6er2UPVBTL9UrwHjL
TNQdW6e4djKfVn204EaxXoZKm/IGJt6fDiPNVPdr7h8TDz0kyshSkL0YMGSYBUftTlP29DTmnOIP
2RaAWSdOkY8h8qAu1oNQATRmi83qyRRiNNoUDscYOoFUZyaH1OBBeMVBj869VQxbNg7IHyX9bn8b
6Ko4RUezq5Pe0kodXP+SvlTI7C8b9UJRAn2Ez2KNqgZLs9rYhXrGn1iLxo2h9GS2mjjt/Pfvofxd
2dyZqOpB7LNjQhr5myFzk5hJ69FbCmUNEolEgdhom0mHYr1NhLUfcWJiwi1Vmb6OChWbh54HHR5a
RYT4KhQqsLL2NABSTn8ZNbcCixcqQcR6iLwXE6CkpMKoCcIEZDLZNNo6/OtChKyYLpvpD7m3GKpK
+AHmG0VkFE5SLq3xsx2k/2aJcNQ3vJYWZZzsYs72IrV75z+ULxRpolMHc831TPhVxjOK6Ig3sABA
avh9mnjLaQIbQ3zP/hPYpp3HMNRA3jZ6tgdc6RHg2taq2IhevZShwEQfy5aVBz4a4titK7Iy9le+
NMvGk7cIV6Pxf7kr/wavt8Lce993U0jczcF7wkCnS5k+iYdWmGshokZO9fxUrG3rZ1tCqnzm7JDD
h4H4V4er/RQnQx6kbfaf1ki7+wjBrtFXmiQf7y2fQdoRYoI9Q3094FNYbrKtpCBoNOoGaILByvqr
Hp3yIjEhuD4JH4MQ3lzLiNAzqRCkw684LAsgt7784hWn/CDqMuxfQ9tYUbf3c5tCfew/W7f0NPH3
zXEnGV6odwLvHyhpA+Tf9+GBZE9LT/cSr3qMk4VjqnSQnxeYQIk1ZSg6nzODM6rWYBZES/izNXQz
QvlXzR4wKUMZ4BaFM6lcfY++dVctBG35dqyUvzK2CpwukWfkzGqiyVmsoWpC8ozAe+wD9EQzOocJ
3wVeJdfXCR1fcED/beTLftGljET5gmSYFoaDXbZmryh96KwR8WN29aX7r+5hR60Zs5kz4z5vI8tU
UsSg9qHHxAeVMOtmOXIMoZ/kEKknLipI0P4fjdgGrh0KDzqJPZleSEkqgr8tCRQUyE96AnOiapHv
iSdbUuuxOMTsNMBjGgbjQP3WLAKqKjzBKX3sJjiKWRcOxTdact+9pVRwymSM2oCsopoHk6XJgsul
Sw7r3TRkENcvay8VpQPT5Mpa15xU/ZxdQJFPf72iB+ZjPdWfWsHv6DI5cOAAfX2YWyivxcr0Ryv1
y7edEggchlGOEIONpvfisMzfgmVS/z145SLwS/E8G9yk7xGbXnhDT1clW2DjF9byqX+Tr5o4koqR
hxRjuimhlm3neQncC5JbknHu0lufsFNnQwufrHVIkJBG5+AJ0UutM/D9KsG0HUGoCml6b/Ko9Pxg
+aMPty3fUzcO5pFjzNQbmzKIJ48AojcJsBdMiXy7ZS2AqeqhPn0WO6IrXyRFugMYh51Esy0+nFMQ
HDdbGFmuEG7RBsrKrL/dvIffmsuBDQikFFOGf7sgRyYB4zTlZ3Ruv7QfaysgCw08ey8zq72gIi32
H/kchzNp+J1zEX3zA6S6m0elngREX1ufMOx7MfF2Lu3SOYehPhMjL8NUuAQO4VTzKElRQI6/CT/9
04Fwy8GsgRLZeY1daaUa5Baad+lKf6+7IOL5qNNXO28dZI+rtg1vhqQYo9j+8gFJjfd/7LKoerdq
v2/UrKqHGoPVWV3Q1enOjtNuXP1emoNnbpPqR0592/SbegTJksF7BkE1zAoE8hnR8VPy49nRsBP8
32otOcJXq8tIo7C9TxNNvIy8L2dDvKFerOCm5v4Zcb6SH3bYcKh3DMWeHKtmReWX4fjjrwdV0hyr
AE3xxQrbN42IoJAWMwOpLutA8ZzsJk3Zbwc73rsOXbO1u58HM4PA4CpIhv2fZeANTv5GQ57djAl4
UPMrcOoppmeiB4g96Ekwc4wCb6RCaMjuud5vZ0dkIV740lgV2JHPaBJgAX7y+Kl8zSVmzGYowqZw
pIJoHsqvfSyylAdk5nqaVAjfnrUggNadERFuT9K25/ffxIoImB/2DDXfIBzumkazGa1PF8nUdsx4
OHG1UR03/8mMWqMVwbOK5TgGg8DPGIa94lsp9Mu+ccC+v61iLHsfxTjQ9wfk0azT5oLzfXE95b9g
0qHGE4a4wapJXdckCzIoh+ctwz4zWursv49YAr8vLpkd7qjgjR7dtNHJrc1Cmxi7xCHnGH7vTsbj
DTa+cZMP57yCoEfT7l/II4Uo9g861alZoq+oNTyraBguV33iAZSNtNoUqq2ntRj1dMTfq+26MOR0
3IWG6Wf9zKEp6Y2dSZx+/dMOfs5c3Rj7sQt54raYHscs/zj9hHpFdooChN+PdtWTFFh7rfGkUQ0W
/ETWlARTTLq+wv3Xt8IUC6vW+geKWsCBU1eeLJu5PAi8msh9e47nOuGwdqeEg+W+OymSFyJU9EFm
+1TgB2fWlglo87WuCxuLfeOK8Vu1kUYF/U5+1eq5heeM/D5XiS92LEbkBcc0MPHp5XlUzKNWlmIy
+6zkmswvYzG4xtWqBAqaGXv+LPOfGQAjZRtGpUH51YDAXPaKSnDUY1+oAHiFShMaA44lSLrbE4qE
bIwRkUEi42VcBUs1zTXywwRR/ssw5cGyxALtmk/ZKiWbs6WPHBufWkwD/6A2UwvzlG6/lS1gDj3e
vuNfdfVDML+RPA4Srvi+1iRySJHwTKzsGHnjHkn79IR8aUEyg/Yxjoz5rzVXCXkq28sUU+WZQFxh
WmaESoZUKNF2APMmi9A25nywXQL/l75ZQmgmh7jE9jJFE72svHQ+e0niXkQW3MCiMEkC3XVgR4Fj
AS2jR3Rao/VaSRFVB9qjL1kNpBWpfMhlzrqVtK/apU760QX0G7lPQ40gm0FLxtHbx7g/EtgoOtQM
E1ep096+n2Gz/kPbt/R4U0UhFv6PTVq2V046sn8i06tgMs8CugszG1F4eEzpW5QMTDeKG71vmJIi
PMMYUN+dBxA+o58u+jeC94/6zsUebLW+3Za6EU2irYPWtWGmrBTVJ/kde5mvRk2zYoHRAVty1fkU
+9JE4UcJ+Jt7Piuu6ZWGEu+hzfBjDEf2Dr+arRBIaVhAXblYjgU+ZuEmQAa3HO/nGyXiV1PHx3TQ
JK1gx1Bivopxte4Jjc0QDtRUF6UipXPEzJBt0xZ5h9pb+/f41MBOSG7CSJlNDXd1MRMcOeYUw4xt
c+8ccLQgMhhJ12ROSMT7ejMIFtkcI8SFN794ji2bNLasU6m2T0jQgcxOnAoDi5FCJchYGMK9sxvh
hhXWjpCGrb2/AhLmwM3H6len0Z3s9MYECMIc/An6OLwKemGKzrxPO+zA4vWxvirIAxdlYDTnakBH
GFTA6wPUFdACNlzpHyN1zawybdIWFaLoyg0ARuWhcAuWs/+a9ir7KaEDozv6IyLyLcfI7ZbGXd59
jvrsVa+23UfSmr9WjYYbiQb7feXFhDZInM9ihSx4gyAvtqTinZlyZAQyWIkSUMkumm+6B+0sjeol
OtSKyGLay2ULhk5TcYrnKw18AzGrE03kgN9BQ3VfKlCe8QG8zGEgJmvDFH1qYciszuFTYPnz+6CS
wzQoWI0VMdHAlHhiRELkvz+FLaQcotuJ40JjUdNV8ZIcdRt55swvABd0AGF4XfJW/cOXmW0GYY7s
+O4FdXy78WnD1ShronjYOiTM+cVxvkEkPuT0b8imqzR6Pz2Sicl7xU8aSuZw7khLHmVwOL73Oxia
dtJQazXh+KvtBJIXbODSB0rn2xMY5ZaoKuyRz5kmSi71sngoOYEc5eed6WW8hP0QlWVrNTY5Tu26
h1qssksN+fMi6VBTKuRzYJFawadCQMIiRL2bU0bpxZAHOuIRlnN+PPQUJKZAEBM9dOkl3AmELQ3N
6otWhLMeBo+VxfTV2CZrcoJsLjCxP9l7QqC0aUEh1c3p3/4oddIvdkJ/tnRGStpxnZ/EfXmlwrj3
+BwO4/tVWdF3eBwJ922hA7WjfDG4+NZQtOA6X7PCUsesvKaOz7G7sDmAtfkmizBYme+Uua8VOJCV
5MhZezfNRCrAf7wh3TUhgPvwQMu1cEMrqlIWMnkCMN9iIHZ0jdHVfyvvRe12Y1TSBr3vXaQZOAce
HlcoTfH2LBZ6kfQRiR9NaXNRbJIgbjc3NTw1PRhJ8Eg7mV5uW/eX6TQhKcsf9Ypq57Q1wCo7SCJN
UW7dHvYtUcmFEYSR2a70Tcw44YyLsUG3bWw8WCNmUwEFy3ipzq76Jwz0ITsr1v1fYaNqRJlxNH98
VtEQsRArFuZcrpXE7A07U9iLWkoU5Xly0rKoRwW7v0k6wM4DTha4C5d7JyRLRvxq7RZfEAya+ecJ
XlFPLvpKtpZJsBAD642Rdam2nRSSrn6xn83HVg0XrpFsvGURI2e+gvKiPFihLZ5AtycsDuWPGfsg
KFH3rya5SZhA5ooemHTgKy5Jpq1X3J2l28kwZ0IC9Prh5y7QwGdDuw8lsA7mFYx1bOcQvncvJj3L
tpZRuzRVSMhpLfUOjU5NF56A4hw8Td9hW32lUzhM5h76mBx17CQvjsJ5ye0e6SErTxHZWjRsybxa
m7dtmj/trcqiEhbvJgQoU3pP9nhVgxzRZivTTzqj1Pk5V1hYxt7puBQHxjsRmvvPoz01GVc0eI04
FfasMVDeaWmpDTHLy4zO21cqvan2Y4FZSOocVePW9PMx4DRZpforxBW6bEouN6+dxsIaC50vHoJk
Jb8f4yyk3+wAYcKxnoIyOSZWrIcpPAz63pN7Npk1ZJBTL4T+Q0yALhSc4aIMLE+COb/sTb5f2x9R
+Qfxqid1113b3rpRIIINEU5IRm2a/JmRstaAmCmYdsd7YR8B9WFeq05Ig7YEp+JAbPO3KVWbE0hC
bGxP1UG0og4Nyg8HkEfaKDJ4gfNkCzwDY3IMlVqXRK/36qejZNzlc4bgMTHtZfL2/I3jDyEPzul4
wWLmrf/DE2by/R03IeI4Mbkt6D/+uWBq7JGtSSEFSZNo/eQsOloMIpPy8Vv1jra/2HnOy5mxd/ZA
1HD4dj5Kgg1FR9lPJ1xuOKXank3WTQ9JNB2Z1An8LFLeJ0UDXaV8clNseZ1SzDt5hEQ5jsgeTpCI
7NQzLlFL+02cLzxyVD4SgLkMLd0RJTj9and09nhjt+VQyrD8xIuOLrIXPGlQiooTPusqlxEso7P5
4PWK+sO081PPd+WFyxZmxVxEJbRZ/YxBQkeVmW3Y8Z3jWvqDhJH+MDcrea4OsqEItO5eb4IPzfrA
UWiBaPio/mJ5qXyteNB19sbBWthyOX+s85LZSyfEGpeezK41M08YZ1ysjhk1+I588uTT8+FspRkd
D8ZJX0gV8KzLEowNcKB5ZefS3ZVJH1Otx+rkb84NGwN5VM6hPc3EOYh2utsI8w6AAmPFPqBpPdJu
Pkr5W3xlwcWhKtEjnCGRIKRFmFb1S4EZ/n+uIMqYHayUghukUAgJUw6KyRSFz6yHZrFTSL6ZDxao
yvvh3fAWMZSDVkeEXkWXzKKC9slp+yzqNnvMoRkgNmZFs/wtiJZh4vhP70cUhBJk9aihVnvqMkbe
hl0rWzvvl+vvGJu0hIxwYSCOM5M2kJRy+6BqlAisy++zNtuYKKuksTL3UvNms7Ll9DoIiCseDoSR
VBNTfqtyXGbz0Ch9hxZsTTFqDRJCNq/s46DTUbDzVTXC3P+UWmBR5cNQZkKsa+HJ262u3ooBvNC+
b3ETlLy84BNm2zksyMA6IrX6SwVfgF5OWS8yDyJC/DHJgRb3j4sP+1wQJdBiFJygNFh3r1d1ykQM
eiELnKn04WraadZ6ZdqnEvTGFHVvGowJcUQK+Ne1dq7CgOL78MQW4p+4a6u6w6cFSRnKcKLCHSzt
+UuldD88Y7M10C8YUGxxjb/hzhB05Vxnyqo/O3HNX8C9eYjUICk/ECq31Ur/ZdqsOhdEwUgCwI7Q
CaCBlpMJODPyq38bh8cUsS5p8eL6aAFMWn0zT7GLzaabwwB7w03JftJAGu7eaCNzMeJhI4c8kBUJ
Gb7YvAJhL/9QF0ycL7urmVeyPUyh8zUfJiMRQYDhMyp3//sDRlMyBtbeY4aaVD1XsbH4zQUvzqEh
8naa3jfpHw3mSs84zySRQSIQ751W3HQmVP8IIRT8aEx15Z0YXPFGXpd8JyHRsLEIrOHgqoaJx4g3
cE6ZioGMOBhVDp9m3L1s7WxZJKj5bw53s4qrmNDAy4Ye485iXHG2yX0q2Z7zzXaNOeouxGosWA4Y
i3GQYaMKI3ugf4I3NOCMDDC1xDTHbx3sW/4A/cmw5Xmzc4XqVJdAkUlsJx5ZlqlD/WKLORBVhTrB
Nx5vO5eBNKeYsV/FKZZJdX/tvXzuM51mMWUGD1KZc34QU2U7BXWkey11z4M2sX0EQ2y2B8Zx+8Su
k/tUGXz2L1VZXCUkUHuqX/1/xvcccEBvGMUbofHxLYeU1VUXZEDG9UZ8l5IfFK5nlvdgNIpn1ozT
iKEFbIV/MN7y76riOpr5U9EJbQzeUNORAGkx3FLCzr4pn0ssF4X2NsNof8RjbighfpM6sW5BRetw
yAiQRO3a9psaLP4kXmPpyKiksvaLoGRPElVoFQnMofhcU19ux4WKgR9yvWxnYd7ijy8xBZjMubxJ
qz/8ZPSsW1+5XI7Wk8vAX3RBaey87fyZvfK+FMUBItBZLTdplqS9wrm/xsbS86RO9Tr4y8vEfmEP
HAvr5sLLThDaxfNZVMDCSZDhhPxHLg6CXtNv86DiIFIvw5cQhImUJbs3Rm2AUT8LcKSzXnFR/N1Q
lzznUDs6WQpU1guaS50ahK44JP+6w3MCw8n0S4IHljyS4BbU02MQoNo+KRYdCTwK7gMD4f8NdwlT
yUA/icesJB1T4ME+9APfHNCIv5x7pSR2SfG2yV3CC3EfOUU0YI+7+Uk8wmdkVscYqznP3j6bbCrb
pjaqRtlUylrdXoqlBnizlYb5hvhizvJ6LlOwkmszLPqDtijIZ1lmFFZGjzHb5YuJokDZUzPBOaDR
67f1stqFRxAvAu9MJybSzAkgZN1RCmQkcCh3zJ8OsVMJxwTsa1rD3FrKHfNsAX9eRwRwLFIDtJUw
CAAcuIiYZb5Uxf3MJDukZLW0EHk+CWnOy3UJJ0UEFaZf1BBAbAMeKWgcL0Rnrledy2X26cEFKZmC
KKGlWlP+ruPz+Eq4/6oCC3EuNYALqr/QnIvyR7JLi01mCqMwFjkTH9uxIVa8qXCLTOKOEc5XF+DI
t9afks+EL4CLSEis9qh/XjJvW3cm21D4rizFkGxr/trirnTpRZGksU+ao4cZ+s5n8Ni6bqilzG1T
RcxumPeMuwfwhlizCjzHT61vxcX2NsqMvQQFwrbSnCNDSR/SdVPNdz00C6ZANvlfbudHrZsi1gjP
Z3JBw6FXj+5017PnfFcrVDOqANyZ5nzlnG2cLrGk56rRv8WHIfHMMRu85mL1zLjxlWR3wWlaUsEc
tiG4X+XhUQfQJzB2tboeAZ8rY30in+mOhD1dLt7gsiEauxyUuIgm/nsKiC6Duz4mtT1qBHDKrTZY
nCmjkmC7Oz4oUlkAqZOPtbSjtUeAYvIdAo9j5SQ1NTRe30GaEaeX2919W2gzBVJ3qe0ie5KBxmF0
kOQR3gxj6onDcjWgNhABkXopeGhgzak2uLmH4aX8uWeb7y3+nQ+Ec3IhyiyTFgDqIb1OZjsNocP4
8mguj7knKWIli06n+DGsKtgLMwLLBzo0QjJjGfdfX3gCk98bxnCLHRgizn8WHRGtVofkksMrQ1v6
ppi/i22UF10/2J3w4HL3lWCmJxvNex9vCX9BPgk8tPdAoVQPRJmQeR80wZTOkv+i8nUU1C+cw8wC
uwMJDcEWcuiqSc7CNhbhm65w7xYOwcsds/wKXsK2+QG093iIvitinew/dbtXIO3fkjCMWbhJTyQl
BuYJvMJaaUMzBOAy/Jxyq28hUwSn2FWIKxejZr6Q7xINl3vA2cV4/dXEKeg8FXGCUhq+gilYtLaC
AZ62Uh4potTN7cWCk/RKR4sCwU/ej0AeoN3JKTazvQBwThk+xsFThEdjZ6fsY85in8hZiEeJXMB5
0L6pwe2p5t9Etk+gQHvsmWTDN2oLvYqDbQU56UA8+p/i0buTqA9bGcbJ4m8Vc6Y7XptIM/llgPZ/
fw6GWqP6jTlQb0RUge6QG6S0LSECHmjkI4WS5Au4UCXCkTMHhX90rsnq/A79cG0go2Oqq7q6fkX5
o1LzQIWJR2i1vcp5u4gwmg0nQVfLCx7O3jEMUqwDcys9kvZYGtJhg1NenrmdNnK0mnzVYk3M3HUY
+fQegSmbWkXWwyZEWZgOutXv5q4oPe69cNcdhIqKhjPTTlhzxw8R8WsiklNe2rXwObpNNGs2wL6Z
BLQSuCJTsDGdKw9WfKW/e316poAt5cwIkTjHefOkMjSQu6kA7ontgIPw2x1BY9hEbTZTaQGQAyZd
iKFZ/Sn0ancarqoDd/rF7SbceYYp/XrrlbaJD/hTEc797IHaaH2d6695y6847auwHZ+HGJTVCRTB
W753oHf9x+Tovm+pAAoGhtiPGkLJ41oS8TBeR/lI42TzflUQwsioFDLTdl+g3hnG7hi9oKTdMyAU
sUZxuawfBvZFy4uBVFhBYvbIBQ76GTPkO75T0hLp8R4B2krhEYr9olcQh9FOjl0Sy7Cn1kznUqhS
m9kWii86E61wIObdemPa1aTm31e2CnCBbmSGaHW/bOPeFFm/xZONVkqF6rBZinfIb3tolMXJV5KX
IhYgqHohgTmVgn9PZ90MeWVqtIu9Cq/w9CMeLKCYio8qe2C8bi1m3fa2hbnaUJfBj2uLLDXZH1np
8OP+r8EaCBWnF4decUAc81G5dJOr5k8M7Ivw1XSNBx53yS1N1cd7Sbgg+ltaGPA7zKMdRjHjlj+h
5ikTLBleOhhOGCcv4yTjYUJQDd84tK2eNL369Maw5etDThNJPnSZSRJbdyCIJQT8zztEZ3MJ5Caf
uzaekCJHb7VVIxYT0ubjMcUXeQ1LQjyGP7chczpcV1qd7HeyNXjDx3NFlvxawICC4fQODJxofhB0
V1NEAlYJSNZqzBqIAjr66u/ao6YhaaGNLSNdYia/4wP6mARibm7hCcqvMwzBC20bZf9o4PiCBE1/
Qu7jbTBXtIGy9jy3Dfx/bikg10W7sPu+NqamEqkYf52wWTo1ejVMdPgZlnrD12E8egOaPhybOq6v
tKHqCEQEVKIByX/TBFA5jEHumq3pZa0Aw0j5nmCapfztKHMt2OWjcpoBQEM86bpedZ+S6wJg2/9w
w8b9e/oWg/lMD73kGU8gjk71E+aYIA8cuFlt4K20TX+lt9GEhL82Fs6iIlb46gsLNZ7kuus31txi
DRbOssA1W05ODQOq+fid6vl0ozgYqSVG/yT7kJjpIPsHFUOoz+py34Jtuu7eiMjKFMzYthiWJh/g
edEAZrEHkpZn/NF4ZnO16nFXAkcx2UotxHPlBMsce3TYhfqmKP8OSFSpa09dbzBnwIpcG6XLvBNl
vY9lFahgFfpJJJIsW6vXRmQptkNQnKGBa1aSnW5eNMALsDbKUo9B8Qejy204WxjwCkxQ9JDbOJnH
clrHAI9SYcyy88qZ4FvG+/dIiNDsj2sMb2X//lRqPpJALKuhQtMssx+heJymK7jwhkJrVYLzH4ct
dj5WDOFvsrfRB+AtCgHW91YSiWyQH31iXYa3pPYs85oxP1t6WjCT8PNNikWu5faWOWNhSZntyWEk
F1dT4BEyf0ZO/dhCiKLONp+plZE6kmTHP0ipt19EKaa3tLkgFf/o+K76szSq6x9xekw/DM5+xM2R
ZH7Eq4epBgQ3RzcF/auFIws01LyLEP8htYrEmDMwcYE8jWVTqVgrXUUQGc6rOclv+8RbRXN9X2zY
g1bL/rbACN4Zdt0rcGF17tzUKCvC+mRp75LiYBL01KLC05QwRuXalkkrysYKf0TDHIGriOH+23TG
6Enilf/rdV5tAawH130wfPZXiLh13/pGfk/zFCks7WT6akHEIfnre9/OJWuFD8EeVF8Fq4YfAhef
Z7KdK6kQfvo04E+uIHMh0l/NY/Eev2AWo/uxuZTbJJMFpIHfU9oyZYDLyKnLtPy2BO/aBA5RNRBx
VjzVLLgv2B1uFe6vZOtqE8wlN52Vcs2meGhBrIrWydhPE7eD2ZUWXbMr0ogpvL9jzSfR3KD2KqhZ
MOjkJCuB6P+d6wIeahebrw/cdMM0axTe9tBEt88TZil+bprha2CGAzXCph+73Bw085OEBtsyH0OY
VOQijeY3jApXN6g2HGTObkAuJSAvIN77yfTgpfBM7nNPfDHRsKpfNI+hGeVYnDoVFKDeHuEFG4Tl
hK0d3sHwiBKcrzselduR+4iCyOux2cIzLP7et2AkhR5RqMXvXscJKinDhUND4GDiAU7UpzFFURJZ
eJ7t3CzO+RWvg2JDraommeWHLUhaGcaWDjgC0c8tIJ6ZL3wye5cFfCx68DgPZMqbyAG999GlImXP
/FX2mBeoOtkW/5YRLQ/FF5+uFWzlKmkMFnC8rooi5NjBAZc1F/HOau2eowC8xj8kFkN/qFV0HldP
L7WuSSNAXhZ7pznwx2v198G/7F+334cICQ5F0jAujTn3YJurQwt2Y/8dJi2vM/F+iXWQUJIFocZC
gTaxb1vL98ntk2FviOHTG3r1FoO2G3DGT28G1h+nkLg4WoXl2KPea9f6v7/RbH53wEi1d5vbUOue
X3+MwWxkA0HeO35ic2iQ6kSGh8bPdiJ1z/D1y9PS4IomnqFpn6xBrZ03o9PSpzeE9iRDXVTfLo4i
sWwXbDwjt3OaPZy9+Q48wDalb6q7a4GYnGXeX7dWDYk/xiiplCEy5lo/54MK+ZyokGNGTFTSCJuA
amIN7Qm4LTJU7h3rlLE71FbK8osMGEYJj9DqSuk79G53zhUBKh3Nr16f6PHEif9lGRtRHbgQ5Xzm
ajGSGpjwfzP2Zyz4owSOfJknpj/ElEr6FyFpk4e+JM85BWMar7e2SUVyKPjLfzGFQvEav6xZr63N
pdADm9xPIozrJdviOza4/+r63xAMZ5oRrCVLT28/l0kC2UEJmi8bnOjtzwufLZyJgQmGFvKnESTq
LwPOutJjOanHI2cg+ez18JDC3xLEIzKSCVpc+KmreSecHu9BhHqMtmN37KKRcC8uX6LHVPiB1uUM
0u78Vp1wb6LXcBmy+57cTIDi8PhU4QdJPgpLjJGlU8AtdAL1l6ag/OmPr0mmWLEwWRge1B1eoXuO
5VMaTQpK5hzDRj3JoNkFsmHOyWwM7DmDrtK/B16U+YJzhMTcq+4SxxejI2QH0V4mnOQB/wsLRkSx
bFA3wdf8n9LcumRBGSKY44rn5YyPWBoWqtJ1cyiBhE2gRzS3BycRDOwm5/QhADMrsmSx9AxOeoWI
lSrN1MNEzIcZefD/6l94Cmryh76sgbsIk2FAm9ZQgZcxMdOPw6tAD0UXGu9H59AFg7AfWw+HEhSs
DbRwtBVnANTIMweTemk502AUB8HJsKCdlUP66mE9ksOwsXiFfZIMeGp4FGZKnr6j+CShDoGzcVHa
bOHRHkFbiA+swYS0qPb3BqmPpPWrWmLMwOnufrlBf0XwGtgazfq46KaeGRyOkEav1tXBGS8zSXOf
qHFX4oNfjAdWTx1p695dE4V2Lj5cga0Sp24GFF3aVAOriINt+iZnw0lNK8FHe3gE9ZBF8MehYsC/
wJuOk4qVXu35LR2jpwSnquGXXzndQ/5xzxUww0hf4h5k3QY0TsgmSgIKj2OimO49Jl5/X2SVrxDK
4ehhf/Z+esYwfdTHFcXgeL4zHUdGk29F7n4K9Ccq+Vs1oRX/Gbi6v9PBPkKQWcMarePhzyzHv9jj
4IjXTPTtOxioV75LTSZkfWaX/Fo/q2xoS8WXDW0r3xGacBHt5I/A9/vpfSJWdaGQ0vTJuXXqCnQT
tgdK+SRUdLkSnYFExWapkfKigJ1EOf4pMoiuBGQuzyNuBjpByYVIU98AeD34TIsYJ+KDbdf6UE0u
UmnPXrT2r5YuSYJmsO4Ppib+B3iiGVrv6TG4iutC+uJzLZlpNPKLk1q6uz95pBK94CAmrNqwCGrS
SNb7VLH9qsyhTrMwofwbt2Ca5yrOYULYv+GWi5qMtvYI8N/no8V0Gh80zpAMz5QJ+Eocx2NccLMH
A9yUcvEzRtdBHFCWp+EUyddkMEtgB+2vV1Cx+n4j6JOgtStgwrCnnwxA3+7RJtBViy3r2YUHGvXF
gKrXKI/MtDIOgVG2yHTu+5rUrhvGCY81lej5ARbc9Vd1clFfmexAkDhlKi+NmkQRrB9CUxYESl5W
DZMSqbClk8mnVQghw9nX9xSBFUGv9eOeiHDpsJmTN3YUBkJ1fqRl9POka76+vSNN3L/rASyUKj89
uZoN4SUGt2mcnk0eEiETTzxDh9vhlmWtRH4HFcvQzuhokyIzvMbKS4u3F+qKfr3qgGWynFQ30T7r
rrqhd0XcguxPmROwgJWtFg7mmeRmOaXuDbvM0oCLtCmmRh3rMsPL4HYVTv8kECY2wBf4FP7zPmr6
ISoVaOClTjkRIk20tq8l0gfzdP8xZInapWHeLQeh4SLBqdTTX7U5sqVc5gwPpgmabQCnaZKBvkRl
mvaqdmRwbTSfxJZ3XkstPYRdixE6TUJNRXcBtINazWrcUoyB7H1fS+l6fsdgNi1AvETYZ2218Jfv
94GyUtiyHPlUF5nGgExNyI5DGiGxLsa7cUdePWYvIqxoXm/LBvsx3t1WW5+VOycwwbzXN3pR2syD
vMbjzMLKta9yWmRnZbvMXVQWhK/liwcbhXwB/0HclKK/mVPg4VcYNxCr0zArXJ+rMN+FwHYKO2PC
JV6yr/kWhy4KeDCQWbzUPr34w9Ql2PsP3FhVMfuj7mTO1OKG5t8Lc81C1///uKylwsS81gd5sMC8
8X+K47SVfZN5fBOWqWTCZbxvnCeiX5b8PuBDnzQdPey4pV9ioaELuRuASxR8ETGSnYMS0I762Dt2
ktVTiTgYG6FzZPxTRuvuPJzTLNN2Ezb+g1KUjKJhbdj1s5DgElGeJqHt/T/2gx+spV6pSPOGnVW+
6/G1B3RP+0WZhKI0HrpEj8CDOTzDusRsar9SRoH+oaZRL2HtP2xYLw2NHiOZ6zdBQUbCo4oo+1BY
SoxZPSgS41/bAHvuOjvWm5t+Daky0SeYYvOnXW//PYUVNz9zrkO6iIZxsk9jkK2ohuQOofrm4hXv
9d37jiJZ9EIfgyTUBsthq34gOHm/KXEiC5NnfqSbtAtW/VFWGtDR6w5p/zSZcTkA6kYIunjWUT4u
IO/g8obqqa6O0NllQSLfC30sGD4hpIAJR6wYfFQiv/keP9LXACIeFE22QDiB+pg5ssBMGwRKRiC8
DsbuLXtcP9qIveSVL/IpfIH+JCvLqGLTwSVeGLPwnXWSqmltvXRvU1Y7uwcbEbTB52m5Aji48z1I
DqaZRuh3XJNuJfpLZEGsWD8FwssqHJHjG8pGsQ8wbpoUterKr0IttNyqckk+T3muS2fVKxHM1rpz
LSWdPz0rYXqA7jdNpP6zhCieUdUY/DTZ00vT3wy60lMYSZglzQ6d3dtiGwtmioZn6dMNXXUVbcbu
HCbzn12UvfVct3BjPFjMfhZ3FxEDgWQbJIeOWNGG52IBNJ86R693DXNYDBuTLVhEQtQCF7lSEgoS
9vEtHgjEDfog/hWKvQScRrwuZpl7/CmD2ngxWUDXfDiMsBd9mf94eoA0+yHAHfig2FMj8iaCYg2t
VyOTWk0sx+v4nydD8vygAerDyirWVxzuGd2Byavuhk+6XqDpL57stM/vyeSsRtZPuuPZQlkwnueD
84bPhc513tjlYX+98VDVDZZkR1WyJm0Aze4uvhY3gY7b2UKORsm3vzL5SG54vo8sNfesBaQB3BVf
Xls4t/owG24xD9s6ss/UOcYPNjlKEGBpZihMtwR1O+xCLItLr1KHZbC12RlUpFnJv9kK9t7oHTfr
SmxT6UnZoAt0N/YQeueDolmlu6H1NBMCoar8os/UKl6Nq8fuHcB/76Az7k+i5OXEwgdzJSlA7vsh
ellhq97lB0ulLFqrs4NqIZhJB5Fc8FsLseheY/hRyrs4nnIY4zB3OMqFEQ9yZOA5ykSa1RkVZlUk
WucmDFe2e85G15J5FGl0dxT1w8mKzWcuUkyKaoi1/096IUw6OCndGTqbti0h8t6+k7AFXz+dPx6S
fWRz6MQsi4MOhWR6wi5EBLFGBBv1qN5sKhG93f+OYXWZ1SAmrKrbgzN5o+TqOiY1/JvjZ4HK4MXl
/YJubVgNPd62waapUpWpikn5qDOmGR3s/ya87NCDRgFhbZCiwAYc6IxzO2p9f/B355BZX6FFXkfK
ZyNKqfrYTksqwyWeiHhy38eNuDVfwOgxytpTTXXqL3FPl+paU9SIl4wfQ+trNM64zlwSsw7nOjkt
SL4P77b+oiTnzFLjxA57BxOCwXreUdhdabSlGXTVQa9upX8xC46fZicYSbxs3ArU29TD25huSa7B
Gfh4Wqq8MbLyMFKLQAaKVgjx/b9z6trQ4Ezy5+pyzZDPojEbYJH6wuYtCO3WWfpTvZeZru2fBLno
nvT4JgeW85MwvxrY97msRyaTJ/NLdJTuNtn0/rahuckF2l+t70K/9HGBEYopOQbs3g/ST+JowIS8
49HP4SPmcEj0dwD95KPgNpF5rUS5CNxXFFIEmWVgIsrfyaEL97I0ORk+me35fDaGWDGhm8fGOAeA
HY/HZI0/BusacD4laLzobplKgV7AC9LXGwJ8Ctql/1lSwK8BUG5aApb5riupqbgo0CYpo/JeyAfq
HOiT3vKk9Z5NV80i43eTuMqd47nMKiohG5eUFNienKsTSC083ETKp9vhNXXH/pP51lKqH12dDNcs
c+5SdMN44HnwOIKna5XqFZGgBSEzuCyaSm4R4zeclngQhaAxoO7umLZ2S/QYYyK00of4bGQ4dob/
ahF9xyXQmYGASaSG0L98DVNC7GUc8x5XK1hPg9uwP2S0bAGom8eAMJ6wAewnk+rQ1Tdq7MisZTp8
jGqk93smEN49hIa4bpLdJwJJKyReFf81kOAufMqPWU5zjrR2Jga++sT6zjKuhUlico8mXO0n4uE/
RQFIpXHP5i/TsXeI5E4ez2freBJCZ0DxhdEEgf+qAC9b8xZBMrklRs1wQBxyOlEAOrcpuvPCyxVO
rSpLXYpVoVT9KftIG1at8xnBzGzgOHRIZmXWDKPPV3a5GX7sgzH0TTSzaU/jdbfa0HSWJXDlkqdv
Xj/ZHUXEhyS9oamPxzrWiD0jHVlR41fmSzxS1yN5Wp7hjPqjblHOq9rhftsCvPUozyGmTEvHA+lu
G7kNHA0dkiCJblSveY4sf95oEwd4PDOonvhg4RPyRhInOEp1RqWDUAIKa+Kgp9WUYoXToH6Hvm6a
jZGp9aiHgZOWzAYxKLpWbH4rbOV5MWbUaEEIsxxcsoofkAeRCcVRrSo7W+0y/rjn27Y2NAVUPAXk
HxJeRFMPJxSAoxkpfm9MujFsdPt4UQRJf+4xg0YCKXW7ho32wVMQ7p6mUYsXSK1+ypmLvGOgHs6K
Q4LlScZlAuoV+XG8nnOF2UgTmSGSRLDaMj6mdr0zjQwf7dOPXGTJsm0AUjOZR2pEBuneetVvSvNH
cWBBlQkAtyGPgL2gDakRpQWK9r41J8nGdyG3Kgp1t8tWnShvFZZ8IzprKdp0PIphjHThv3M8aKON
LtK8aiypzlviy3MAfQoFa6WRNMI/VpliPnjwF98poHAlZyAT+z/RdHrFzrH+alvaZEQ0DpTAlegY
I/x1QP/5JUKRZ2My0nWGlyvkKrVOv8p51u1AkZlkut0i+ORMPEtM7ohDL5HYZU5VGq5bGB4NNXht
UUxX/aJqKmTtWfTVDi2+5v0iJMCAuG9OtdLfwZTCSz7BGg2BMts9v+6ORpyzLG8Y6h6RJJhtTo5B
yKnFn3gGC0H0zpqtNwiboMRJw4hHYJEKUoT9U/OIkBxxWDtCMstCJOWwojry0hYF8qzgdqeHKMcu
HONXJVSslSoYqyUsgfzhfwpllXCfzWfYA08EYr+tojo9ug5EQ7X3IBxEuUWPlQQCDeGvb8YsDBN9
1PerGL6jEX0+70whyh2ow5lSPw0z01syNOjkC/DEm+JbflxftHC3rU4pOuKTAObdBla+93qDUV5H
i+pwrPr4jbr4Mh56cWH2rTkP6ahsTOkOzfmvANaNEz0fCz+dGH8p5ltaYLLmj7ED4C6Nzd9Qb0k+
XIkwZjj8bX1uE6fdSjNHErY06nARqGXCap9JaAITrSjMNI9jRJ8kadfmgwyWSZfSEyB3fzOXLnBA
07glRgntUTUCRcl0Ce5zV2Qmv6CaxyNH6c/4O7vsQSIAGQrG4nQ5qUE7dwl1QslYhdKUJnPPjc3m
HoJ0mh/y3o/O/NbJYd0KU8eDtDWLH8MzuytNs+K+UJiNgvF0b7lCZ6ZeJJnLlBAfaeixu/SeuPd8
TSoscUOgUIX9Y6Uod3HwsQmlOWKghHCVuioJBdFvjvdb54QEPaPeebFJ+9+Xa4s7hsmOKwZJYvjV
FDgA3tzXzVrEwN5IJdyvGGhxJLJ/u6FgN35BKypjzqiWYU1jTrkBYsK7+MOp8e1gjXOBWHMVX2wg
Pvu0tXelMgR5kdza19cCD57jOD6gB8/05EYMJNA+oiYqUFRzRX8iWZz7JngSEdMulBflrtZsb1iL
Ru+bV5xR7eoUAyb8rL1lsZWjQIOWiPLuSPSVFVAvdowJ/rR+8QW7dxfRsStm2UIni2yFqCPHMF95
tVb/kNlXQ4fEbpISZLqp0wQFZrBxfwcr8oggH36WsF8731xXUCJWRYXibuitP2w0h51Hm3Jo1g60
n3NVOV+vxaBvCROaOAtD1hEAIn1/lYkoGK+QznntiJqFUqzCENproVYQnYgwcjCGSNw1H4VOD4Dk
tJ6ztb6C20MZrCE/CEotpt5BkjJdiSDy4XtObCQoRAaUoIm/Sd2YJmyGYGOQK8JF18bWYFS96ZqZ
2euRCBO0Iu57RZlc4/0W4CAUnSVKxpkasd8MBT8Gku+iU3bPwguOMl+r3KltfiqVrqKu8AC8j4sn
wgMd9K5hB8E4mxx+ap9eJOeCO7JG5+ISOhYS7C5gyd9F/TnmEj/NXBIkbKJdpimnu0CAOIlNRb8D
S/sxcTIxLhK2JbdECYV+r6CAwv5yJxZeNZnwCKxe1g6op22rqgSjNP7niQg6bb9neWlecmC85fc8
kxzcDypaXjRhxW/1BAezD2T397Ms7nZiJnmVycYs63n2ii7wpDnnGJ/isEtB5cBa7vjyoIQKr+xc
ZYvVaGCCULF41oERG4i57g0Q7vA5KfhjWNaIAO4XiAJW6VhHjuY3GubRJArZ8F9WjytVfI5TBSgn
uI7Vp/y6CjngXWwdyVHYdnh+lZxLF0FoZXXJR6rIVmnLhbEIN6vQVHQvUkEm49cC1m4zNzyZ0FSa
xTcWzQufmRNPIYCMlCLKRxinv9JUUSEIW8o2h7AmanoPPEAT2xNYlf2mxcca0xmgkiRoB6TEwGgN
liakUuojFjSq/puZFHWOyiXs3DuoiWzjzSY3WC+M6AGPKQr1ujmz6of0CojEjTexjcq5Of0PqzBs
N6rSnfMlHxW0Znsa3PWWGWezlZFN9kQF865+UKavl2uCetn8btmqoC8/mB+UIkt++OsGtE+QrF9Y
PRRl1HfKz7/kZPGTOpz7uQpJNI99M6VEt7yjrSY/mjlA6oB+tOoglA9aop+/mCrGpIRp4Vrf8gtX
m7n2jVSCmY/eJFd8dzNXTCx9bpD8f0hOdc6S9OFKVzHscJBfNXtYLRVA+sZ3j57GWoWOHWBsyL49
qhSzc0cqbUeXVMCcuOzGhWY/ofQlZWq1SJ9fUIXVmS7iZY4rvvIC6o0PkEoLR2NvB7wGBQa3J88Z
9akcYRFue0NUIp6F8hgUM3pDMbIT6FkOP5d56kbJGjAjHaDfeRj6zuMs5Vy/FjB8fUs/jqGOidcY
Spt4UMZr+7uhf8y2b6Vvgno6OdLAxSGmvwmLNmuwfZENUEaEpn5MdsROFHEHvfuM//kl6fF5hZSD
JiRYr8CbEy06p+XEvxwhCp48HbCDJlRh5IuJmrMKYzwUtTVSGpjgBaYPrfRWK/HXUs7xfCkwPji/
nk64xejgcurRfL2qp1mchvBgYN5A/qtRl3prQxxrLoM6rHa1kQqVDsAFbLCID1fU+43JagGl7oM0
e11a7vrXytOIKHo/yPot74HzisbLbvQ1sUcFsG9IWcFuOWTkdBxZ+4MPBfayOl9nW4fz4MJiMaKM
FdukWwS6jHP8MfquB12PxcceG1tO15qDEsUvwOYlc4BXdIL1d/9c2Pf4p4yBnRUJxcryo1PtpKIK
5GZE8FUk5DvrC5fi2Y3pv4m8YS1tNpsl6l/aHfPiHC8T1R5D0BMPXwyQAnpsG4FQl5TrrCTml32U
9aAKsGU9dUsxZVB40YaEHoYnfFmK1ThFRfx1JSVX8b6iC7F1VAwTKPIRI/DutE2CwE83IAvoCBVs
5d+PhaQwcHXSbdgyZhhbOcFmRNrX6iMb7lkRfvZVXaGQQNjZhuZ/9MSHttyAHQvkJM6GPVhwUjlK
/45Gz16Tlu6aFMONLmgYwL4ZVW6L3Q+fymf3wM+KO4YuQfYSqVqyPtBAdafuExai/Y+9kO0BOiNQ
tHmvSrJ/mr2/9jObRlxcnY/4E0WmPvtG7Lcw+mzElJ6uVmEWVA1qyhmJ7wvnPtOLJVGnrizYtXOs
DcU48kQ3w/juwvAHRP8oN5pZVhPPB1NC0Loi9UAHndYwACdAHapkXTR0SBVh94B1kIGU3uvmj0gu
SNFxrG/06zwpALdtvJ0MtDcEGtS41s0OmV4PCLCvdaFB+mmVHtjmM7JTafVUtEmJ4Vg7dqPGOCK8
00vLoS4lxl7Q6Vg1d79jiweg+kH0erF3dTfBj5eyE+Hm4EkFaVmcsb9uf59ovgQxEiPlRv+QBB+r
n7tJEfh3f/gx1VWj4lumCwTnVU9iJCSnbhnxG3tRZwqinTGpxTALBRlg/Si2nwru9WlQ/4lj5t6Z
6zqjjNxg9vniypcjMW7Qa2Ru2t+cok7R6wMih2dBmgAgxTZm8+KAqXhp+fvoebnXvANT+mlgV3Xr
qoZ7EejXuGwPRx2FpXXBi94WlB/8gGWnyRA3T492LJw3/pkZejx28LqK6M6jZDhx5t8+8Ask39BH
0WOayzQROu3upYjWbXM9WhojKYSMFD5W0Im5X9Z9uyBxKBewKfoVacdi5uKZk5zuKwGVq8uVru3a
7Qpp3DStECi3DGFpowe68o4i7phJk1cdiuTzw3BgzKRO/ur9v1kgIWu+PTf3ZZyZoT9uMm11jffC
w1m5Zvia85CJzQ7LE9GpYhwKpEKfiXldpkdzuK8I5FPZvdNLzw9ynKKTTRCfVQi+j+1UI93yl2nh
1F7rpp9cpFU/ICnltObwWSPYvxB4JD1eyouTcSYTZTRzvQi5QjHFSWrD8YaVpGvm9r7/kR84cQYB
OMBbcySWyffIeFIqv80o0YLlGzjTG0/kJQzbTLPNSLHa9Ka1nJF5YOgbaQuDd7LfGrRamIxrLBUb
ani+7rbSeWWi0jwe8RyKKLP/Zwe+xif+hqRqtye1629ltCjGv9AdP0Z747CPgZtIhdqHAUJsFRcb
sNbilkcYA6EeKEVpqWRTlsJpOaqRwTu9LDm9NCOQON+iu3a907bcCWicwWxuOEAl0sez8LyOp010
LPu3RrpbtunXdYT6tsrA9LoEIVnyj69INbTWlIe/HS29a8pRBDF/ZyBy37kTj8jaPxWdxwzYr03E
141mVvMbFqTLSSS3lLoBHboJvxTtPJ/AIH44Mm7s2cNJfh8d8oATyZ74IL1Uft++HFKI3zv4lvXH
pMo8v3uFRAO3vxZ9wLqYtTG9Qol/64Yjvz+chtfuvkStizj9F4YZdOfizsmtYSGvU0hW+UykfNA5
o2t9BZVbxR2KcvTOH2qyKZschK0Hf0d+nkkiI3QatbgOn3vVEgRtIcEKcZ6cGY16XLtN8jRAZCEb
qA7jRK2dnRCgXmpMWUM2+fLtXfbOzhzYTP8yRpDcQcaPS3qEkBSDLHCfcxH0FFjfPZHkn5kYPdmJ
XaXi/3iNQL64VD6HX7XgpjfKinClHS8DeoS6L+2NVyTHS1BoHC+MYFbd8qzLAk/9yJ/mjQ3CGLQ5
RFHMCafOlsf0FeP1QvdEwfZ0CSufPNTVDRCVL+iZv2qnH2qRTQwfLo8WUx4GXCB/L4NPnieJaFUc
vWQRXtreaESyC0sZa8UhPNJozvQk0FVrfUoWbO9cU0SlKvi8JN7M3+h3eNxW6MIucuZU7J8ap5rc
DJYLrTSwofBU3pQ1JRzLn+eumQsPDPmJxqmD9oi4qwU/ec8fkx+HzG3Ml190uXCmmX1STuMiUo3h
74DyG5gReiS91xgP4T4MQepsc3WvatUWl49dRZrVKmurdf45yiHHd+oytK4hftT4biNoA8aHyH9y
sPLV0U5ExpkxKoWtMcXst0lYb99cN65W15IMp9IBggT3tsHOk0zcyN6ljl4eBOAYIuHB427gzEJY
56fL/fXh17+X4UmjbSH4cLCKf5xH7t5TISN5vi8gvJ2k9ymuD/WpLUz/+dah7OXst47z2bJw+JrS
2uKyGem9CWWkR8yt3AfWmYD0org8pMzfsya4/fDrQ7zdqvF2ZgoYiVj7EoNsiRWtZp5Z+Utb726v
y+a/Oj47dpOBuxfptlYuShI3Ac7DMrFmZRtYgxVCVECjacoF1wZA8AKs+YPiKEMzPMIhYrS7UaxP
1ew8hBOva6/SkBpgzoJufJEirY/zlhmIqqPJqVYU8OkSF0OJ+dZq61FaiDIXvMKELO89F/ePpaVC
zesee2xyTUArfFOeUM/rvYA3tRR2y4ETC0VWPt8suNh7aEWLzhkHyF4kgywvjInvVTy9/4Mn2f/E
XN3X1ST9WE/DhmaD+2P0T3lN6a/toT0dW+ZchTsQ5Ie75wmhdge9pHXa/HFY0Jnvq54MiMkZKpJL
/A86y91AJSVfMfTq7zFfxpvQ5u1kohRDoRj75oQ2exdxv33OT3TDaYyMJYj5bogkcGxvcwtcZl3D
ZuuQVBqnOtE18pSOQfmBH47JHB+GMsxRQufQdqGRMC/kjQZf/dAaj7qkz6yPEONOwP9mqB0rpAbQ
KIwVdDuXEk04wAjYU5cPkTRQYf2lFHF0P8G5NHKR3wC5pGSzy9LQWkPHF37hrUpePlaw91QtIvlg
ng15AEeaQiPaF0rAS2tS3zi6S4tfBJM4f2BDPp00mC81Px3GrNnQgT7qDZTWV0tIp4CtyjqMz7wt
1HR7SzwBXO68iZlxnpfHNlJSD8nlt6QCHj+fiTAP6MKlE6OXLKPbovB8DgbBV8wLzJG4IP/YyGdf
Dr1ChdBzCfByCzansg7lmOMVc8dMCMVO74OJN4AOZD0vEwW2++4LY+fuQBhzVulAN/BtmT0JoCvk
dx4v/xdxOH/WMLykAGKFRA5jcqVMC1o+FwMEBRt1Dxx5jdEZgcJXT3VmXcmaHaVBdvNp2FHA9yvr
BE1PKyr4oLrKpP403Z/Hzgb5TZ6RyrPufKAUnwcuJ70b3MYA6uZsz7A2rSFmE5CihnFr2FgjEwjW
RreiO5FQ1D1mbGG0r5AtgLJlGO0b06vTyEPwzQruYpBYNbrm3Gp3R5p9RGZgaUO7bvoLUa3PcCkg
VGGc9wQ11tb3DlIbRgMY7l2GSKsf3S1VhCsD73xmGKufinxVt6tbHg+PL/O2AyPBYTexhMvEkX4N
oeqBNKX22nnTL1dla9ib76lbhexgb/auU1hl6bCOQu8r0yUCHZf49hHGNm1oaOyJS6cY42Gen1Sg
ukOxWRAZ9Djf3TzhwhN6zczXMScXZ0NywAJb7sV9/L9u5x2It5JdogqJE1/uN0NlAzlFa91ueIwG
KKtVOOUqEgysYnoofIpw5oPtTR0DA/M+uOCPiG9dPVBSvCjVjzV4rIpAY5awv8uzwTPy4cWimTmh
0sEuBxQEKiP2Fw9Md2q9DEUtAwC3WR7dmd3/8QUY5nwP/G3oSG6+2KcnQ/PfYLHEB1WrtNzHM9aD
zycBIYw2cJEXp9srDi5Ro1c6gOpp1rC/ONgttgoZPDqAZJJFoV8oD1KYPMQYx2CxNa8pgXRYm3h3
wifHq3uTo6Ki8Yt/EcxdkAzwxGEY9FILDF0ZMNWV2lizgVPcGt2NCGssbz3fcdFSxbmjHw6iO4SR
J0hIHoKSrlKSKA8CblAo0AXHclli+RM5h4o7VU2fGI326jMnEghhDpZptI0c3kBp5Rp9ej8EhQg4
HMbDNDuXzMsIXhN4SJgiakBOxNIwDdB8kqu8Ea352IDfR/GohV2Xs/yDkiX5oCDgLLwgbHJAtTj9
ObCA4spmL3z5vRoxQ2PheKGVHXcojbJQIfQBIdNb7R3cSOzidNhD6s6c4KKlyCOXdrX3Z1fxkxPY
+swcvvjslerzfzSZLCG4coM3jDR0lnJZA11VEcvV1qW3HU2WxM79zulH3KUpBHOHfmnmja/UwZ6o
QCjyFkGfz7kCjxSW3z2Z2JuYdN6gf5rY+oDhUhQEcSm8iT3roykcW7vzFizgI+cVSGfYLleS1aqi
7U9b/fEbW7UeEY5q6gkKPFHuEmKRWjOKtph9X2LggF4GoovcZhk1+6G6DfX/obORIKl1u/ssemJZ
OSfEgu1oryW7qHMfdP3PnKaL5czoZ6QuiAgYnf7eSc4A9diXDYS9h27rBNK1vkuaqjZXg2EuSrls
mO7RoF4wvxr0FqAkYC/0ICeeRYSXihnRPZxnvTRn8WikpwlXoNR7aHIUVHQ0yy1/Gnhz+CnVtJXH
IHB/bbbDT6uWsWP0rPG3W4xtO9Viro3WPpVxC/hoTuoYYlE3MTvu+7ciP+OEAWS7jKjDz4K9B/Re
Z8XzYl3PfP57sIfi2ZhF7SLgGyWQ8qvmgJgYyxrQt2M8qmWYZMHNH9O/4CYT/FlGlWwkMHLFVhfq
JOuslzBidSzW9dw5GxemXuO3OZ4ugwzDyKsG8U5k+qJncA9S1A1z3zhUukkMMtlFWCLeUSiWwpYx
E83EnyYiMSuZG7Zv1F/FX+vfn0B8dYT0/1nAmNcmPczNroTS4D+WQFD4HwDRs8sE8oGGQmiBnHn4
F2hsMjEFP52Y8YhCYkUhYQtS8yXUkL3WQTNWNmh6jVWD/IRaxmTfZKLPGyD+UaaTqJhm0g+jtd52
uwuZenv0b8o19jOYcVRK38d67jZmQka1tKvUVy4VsUuiPzW3KpgqLZoB7hsjsvCcvFcn3upa9rIq
gQGa+GqIvjuuVu61v/cYMEx/945rD4OoHR9kRgBElFdSYZnzYelw3QW5SisAoCZ8nE3XS8DaaJKD
usgnqbMu5xQfmm4SMvFdL7sTE1/WpDUiSo6a/QVxjlVTQ3kwmqRtyTxCEXQjDlazEuERL2hhPqIs
hDOgdVdfWYppMYMt8ufRtyuBZXvcXf6rnvLKNbzUqVTxb+OGbwyKDFgkcHiTvwCxEk1PHMVn/pvy
RfzdEpmXhmknYYyzJRDu7/5/K8VwkS61t7opcx3cLblu+2o8nAPctlsO9MvL+gxdi8718sb8w3Uf
BVZoF1/g4TRs77tlJLuoRioIUwq8x0wn5jOgNyNdsuXLo0YNikYAf4mFe5IxA32WDM4gTjzYI5k0
8iW0f3T5AP9L0ukcAKixTCYBA/eb5Veh5bhGOIK23jh9A7igzAYqGlOVE6ijskFNO2VSEKxoOQPK
FcXuZbkXUbQLPsuMk7ENcwLHUSz2/0p4mAVGcBeQTt7iD/FmMuHjV9sd9T9WbBRcZIwTcRaraV0l
/oODm6Yt3a/5HxmJqOcrah8+BM6gOE5dZ+0ZQOR088HeFOSBZfH2B1DpuXw7IuXkEq8+IFtcSHaB
kqwZnhC+hkDuudpmTlqZUWX+LSgVMnENZecyujtVcn15hH6grIp7t4fnrXm3miy3Bq4n3qbkZY3v
u/z/5X8CPhEJ/718frSnDFEKDx9eVU2nuecaUWDA1paI1bOfzDsjlBiP1Je2XWatcoXSwTLy8tyl
F1N2PRQQdhnBdfDNVywPfAMCIWHOGhRrupxVgds67hOREQews1Nfbc6RxjfGT7cbk46Jxme08t3d
CDzkt9ZrAhHS2zV7jVCOlz0aHl7QpwWJ5GM4g6bxeUIjgAAgwiaWFBuFYck902XZ2MNioL+aZL3s
r796RNuhe6B65L5JtKyxZHjhMCsuy32grzAmriqgMThWQrjY4m6EOCpX3dFakYaGyu/lXEw7bA91
eW3Z/y+TVU67kwWIfe6sp/Z4laiQNKawaaWmgb/TSCEV0hkVhhEpdoXGCJB/b7BXiqVrjGGkljq6
kI473uqMXp67sJfz2R7wgH94tMFRUWHhWP07NhkrhhqxE6ZbiLdDm3Ds5nXXNYcHfAVPv0N+fKfp
5Q+0ScmOYvUTD0blu5GXxiWxMuPqdEGMJiZROx4Qe1ng9EUszQ5EKz5B65EBq6gLEdj7kR3iYJX6
80FR/GKhMNaL8N8zfcjxQkTRz4aXtlnpnGvGwIvP/B5eru3XUNaZ5Tx2XbWprWM4jAQGZglVnx3T
HppJ1sw/PUp5z0YCDB1ePTxK2tkDCZA4+lSLbZ9J+wRW4jvs25pdWWy5BKVCEkc4Adj8xl1B0ixo
we9quRHZDGS0QEGpBBeey5jwuPtcfJuPMYbJUPOESZlpbJyukZFwojy5OONK8Or0Y+HY2eP/yVZL
hZewNTDd7cn3T6+s+SZAnDOlQOKx3U941vRlIaYyFAN3+3F/K1Jn3FqVviv6W5xATWUI3rG7Le9C
0FZllXQoXtaG3FCcu7TPqHE7IoBjiaTQNrvQfLcdCtkoqgIz2XtGn2cVJaDyQXvg3/RWlwK7HQ0A
JRySjR8nTL0HXEh25qDQk6ZuqNHpx4wduStwXr3P2whV/wSKLnLvlg1/zIWcaVrv5aoY/hY62AmP
NIfpN03E6PHkcx6MJi0GJwDtlvCIkt0fAqw5vhv3yRPiwR2Bd6E2ITi5IJS5zaoQ6bNyASeLYOQd
5mXed9OFvIg25d05OgIopdTThvrH2+/gScHA61EU/29oVFYc8Ph2rXHz6Ih9OL6IOQzyLKZrc68D
BcIs6o0mj1xniG9kkWo0YLPRXttaRsPHojevf9TzoiMbtiAK4zROqrU4WUjtvCe4k3uZkI+japop
VMq+0wrdZU6HO8WSESyQmR/JkCCB/OJFekXhT9lj1Mx+7YNTDZ25XRp8OvYulS+OLWSjn1E+cpNp
4fvVJyrgVwbU3mHcGmFHs7//kBBz0vBoZ26R0LrBn1tFgB/lK43EC9pnHEuFCNdEp47692io2Dk6
hRaS3Nv90kW2FTJ8sQKRwKXnsuGNky+fnZCSYGmsA+mM6Bu+Fiq2JJNjN+MSwxRMFBZY1Rre04PD
TtPcHkd2EP/BNWQkIyvceDzeplFDxqhdt5M3eWy4nd3j+NqbYkW4+AVr9k63PFSJw3aQgObdue9Q
S55f5axzfWKRbPHhFerHMzzTUrlB8hq3AjGOLckHinspBFn01N1ufD9AzuHWGzdMUuAFYG9epYhi
HMu83rVeLbpWBVlGJw48LmcdFKFdcSCg4PAzDHZKnuU7lzjTthD4n7H8g+06YNaHo2XXG+a5Ryw3
tL87PKdFyn3RdcRPUhZ0rqx7sDiiBCJnuob65hmYdCLm273EtivZKy9B64z6ZXm8qg2rvkGCG8TX
tal6FJ3gatRXrrvOrMFIBe2vgSGVJQtvPuA6UAD3kj0yyVATxv3WcLaTPV99UMrOfPpqgq28g8i4
vitb9t/uMiGmuUaeX20sIf5ZDKFSaRtQy+gGOsAvkxIfpQYiVLuJOxmlY/MfoI1bm7JulmSvzQgg
RqM8T2iaggeoYLDb7J0y2iLVvS9XvF0Hy1NzwUD65cHn4aV/SpDVuH6yLvj4uT1cMVtv+Hfk1luj
PHMAt4Wda9QYeqqga9oI8g8W5S4NzT1JdP7OgjPPvNVM+FdbeUR0DoHIpIhFzVEkTv2FHXuk7BiN
LFAuR7W6VD32ceGZ5YqgeTJps2v19A2F86i59NXYuJ7sq2VFftJ9sOAtmSVpLOaGEuexsDUxnuwb
xNUGSxskL7BZWIuIxDKAxNVTqxuc78e3HoRT04vNEGX6TCenyJEGJCAfmBK38d6wt63UGu/kPY4K
E69wS5rb77uzJPHHWmJS5knif3f/6aqU5P9Aon/gUKxodla5p7Vhk2zDbga+pUpMrTqxqbkOJkCu
wvnBEytgYMD5IxNgcwAG8eemNaTTG7fujSQrf2QHSaur7wHwl3cZYsGUpVGelXnfNCZyd5jawp1y
yAvv3sy5NcAKEjUtZ4h2IcwBVNYKb7XAxrUtj+7ekuZP6Xz0ONWaql7L6LIlpPDF5VTvSJhb2BWz
rg4IbHk7kLKroWvtbGOGj0tcaEK9WcxkWwU+oa+6Jb0biTPgx+zA/KOHCqZz3PGoxZx5ItdrYTMh
ebGGNQltriFSQCld//kcRrWXJ3h6lv/V1sr/najDNvY2+a3TO2oW64B2/u1GaGPEv+Gtb75+Rdpf
aLqUT0ZKI8KtXlko7rX/jn/qQH880I+RKGwsXV1CwfNI7vYF0o6sZ8LkC93gdq4eBcr1k3fspr5K
OjfhG2XzdpYDHDsL68EypLOJIRluV1gx4ZFWSwGPOInXZ1JOy1Zod7iVdckGE3odNImHupZ+nfqG
7qpGknbrOX8AKvOyeorrkWgJXODMrH5ceAXBtYdvdgOIbSw8o9aFaGwfXdw7h2PSigh2Hcp8jyCC
+SnqR4PTyqrXra26b5QmS2IHbGgic67gesVUcERKlCWXEJpaozcBP4TBN18ZpqO6YO2/MGNcMLGP
SeN7GhbK4LK3oy2W9+gVj58muoyJB6ETTiDlWMcFtJbD/IESSXm7jKgioPB2gaISpzvqb6f06+DP
rGIeIb6abLirygymj0Xmkw0WOAIlk0Raz921aF2cYi9K/Hm4ivOSHV1EhsnsdZfzJPNbFAVtxOq7
hYj0CErhGFDhTJxVMaAlFNNybNsm7ba1kwlHm2sWIoE+8NtbxY4xwLcVcLNy24h04FgliV0+wx0N
e9Y5dBGYk9qAyjzEM0CZEZADD8xMZDtTmYOgOvdf4QXQ0i1MWnGTfaDC6y67yKHe2/OxGdChQUZM
nGRHGVPsgn0GsgML9UH6N9ZzD7RgZbxnOztWprx4Xv4sL0ByYp4anFRLnWKC15WtSx+S5gfs2wJn
5C44QYOWo7L5Jju9pT16e/ar6ifFKWi4bmXJxYL1mjO1/QSOWFS8nGql5Lt7qLqg7lmWHIOxbRrR
tnpZJHG8jIIWRBCDvcCak1cRfCCLfhUsK/etr79LEfEQsC1Epaif2jsvb+8KGuFKz6Cw9TG1UvN8
7og6XzGaT1/O11jfWUAUa+rBUDo3ze1NC/m3dEnWqGu6ls3mg17tFKRsCM08MBBptwuONVYOVbS1
LJq6/xjn5QsBotbfgOHtuBOlnH7rrhdH76l2DdbWUndJkpbkLfAXAG373mwamG9MeIC6aiUFPmip
jlACTdFlVZGOwHrV8QApouqjfXX06g2rNwQuu1tJ+ADVg3DaG0M5KH9f1yWnIRUHpnelFn974o1r
br0PLbF4l/ffIP6EzkgYjAJTQc7XQxiKVkRicUJj1lrQaAcDPfdfkintF2C/1JZcxlbOfFTzklGR
1WvnfmPN8XCginSdTdKjmD3p7G2kQd90OjLmRYH19zcmC9pMb4RLzrxL79jfqFnMI/rMzADj4vYo
S4TfY3LHHGQZekb2mgAJHwu1eybEPbAqCTAWmGNUwX6oYjyau/TxZ47PZ+FlT+xAa2ISmYFSKhre
1RvX8JDF2r5nZ//RPnKfaeD5zax1dvVw78xLRCZT6Ib2ANA5FO7uhIvF+0hxuAeBSoTO/9m0pvwF
k9wFqGlISfu2nrgYgDUyj1HBPHK+dtz7rW/iBub8OeHaiCTP09yCbMusNWkmVhi6fkok97CgrC0Q
HG8Wo0Ro8x58f3MRCoM0EM0Y/AaEWlLaUKlcByIGY41XFXlh5W2O644xjxobbTbYmuI2aGIJdYI0
1bE8jyu1ho7Inx2jLtEVb+Q2POe3cDMztZxrxB1Xskd+5VcTKkkMxKG5QhpWXiIV/Cgo6nF0YuoN
Iv3LYrSFU6q94SsGCE39OnFEwh2fAQunv/OIldB5wCmhbtS2u7UuHD7UvMao5U7uI0sXZotRC6Ql
Ipty591chgGP5WtwgVkiYxvR7a604R3K1pSW48QAR1lemHsHZ40cH0Hp7dkLOTv7gqeo8brsviHd
0wPGE+6v5gB7iQWUSU6lJq32JFKiiMqViOt45IuMb+qCNarfwM4cQ9B1UMC5K2HFMye1ZSrRxEqJ
Fi76AOX7oQPZE0Pt3AMYyhc4aEgPcdCmTArKCYKQmLmpfVSCJmqWg5kvNOtBDnMN/0oHFvwnWQq2
/WwYWtiCZBi6XtmV5EHtsUzRMFxNsMYZMvt7j7MuUnFxqja01L9emd24Baj+S1J/fvu6BriZ0hhw
lV4XLh+Vetfobh+RAOa+2ec+I6WVfR4w8q51DPnGXFa9PPYpu2hdXt51CPxgonxrG/Jr9nqverZ3
WzhopQHjYW/ghKtlkVMb4HQPIyMgOWEZfw7BpQHHt/IYiZuh1jUYptQiHIaAJpjfiGwYWBto94b+
I9nehAQ8se7LUZXLQYzv3SXcIGKGSfYGK9RQ9jNESrYMkcNIfytYtkQveIMRAqGTD8NG/hNo7pPa
UoC++sP+l9boDtR/q0UkgUPeZYU6RI1HiRqc6PRMT8z+ViIX0zIXy/T2mKyJjm1e5VR6t9kVfY7p
7E5DAmqnGQX/I/LOWXGVUH+TyZg6i2A2s1xBnsGPHLOg2LP6JFQRlneUUjnntug8AcBWcoz7Sb65
3rnvhFQIhhxP5xq2xtGT2rj7QrkvqworeFzwJB8YRvoDpDAr5ue5+fB32r28wMCad1mlVc3KJcD5
Q74WLPbpj8I2W0XrlGy2WTA/YiJG1PIfQkxNaa4KFRVIS6cmC85nnWyOJQ2mcA8sZ7xqkTgOZUL7
GAnJ4cmU5t2LDY/6RnpuXZbs52Lx1s+3NO6sBNkumMEs52AgYav6MHwgaVPFevjeO29o8htQC0sA
KoPRbF3sJCKdpo1PVWZgGck7nq0z0BmpVPmO+NaQotSyHPul2gLhuoiqm3F+to0ZesTz/6ur4ln6
EQ0p3xL5WwxaeGLnnInOc1xz5SXpc12P7UUcQ/rSiMdg0u8BFCxa6EA901EgHZdMHpNYQMkXuxGC
l26RbDuhtoyBkVjMLI4/Wz3o7zNz9Z7ScAExQCvVqn25eXIau9jLgiSVC15mYuNufm0BRKzO88MV
l6b9SG/CoupwmYztW0BaX1qcvSAanleM0UIo1gNBfuSR5JoOCsAGRnFyCfbzpR/XeLaKBUzQCoOp
rJZfXDGSDT6BiiOJaECFEVnWapS/UtnASovoS2NB5L1DlOzGn9urUn5X2KaCrJHu+ihSG7z57a+Q
AXIZs62Q8bmwTl3elR6v/P/KZ2Nw+5mJVF0RWLRYsh0KV3QORI2L0029A+pcYHcfil7wGXdQ1BL6
BG3mIXasvfdMSEBZHUXxdxak+qaAkJQuwi7eTKySXHY51epHVlAmifV4I2O3Q8pvExPqCZHkgB/f
2Ys26hObyO1ZE2jkaLyCry2LVOc10q5QPpSX7j1EzE9v6DAl3vI1Rb8dwVLERWYjDHU/jLnplRko
fI2pPaHSKjuFd8mRsDAgg/UJUKZoo+rkS1dF1X9mPgPsWxH7TFYkdy/ywwlkv+BmJ0aYNKUODjdQ
aTJeyi8E9ermEy+MLaj0aUoyWfD23/wBoi3NeCZMHfNRoiiyvA+LbGIDPMz35kzWyeMaeg1XEUfO
lCkoto1AWbuLjv3s6e5X6cWPrXBX3LkEiTlc423mI8+LU/9XPumWejqZbfFzUd04yjK16qSwvaNl
jNatJ/a+O5uuI+W77m+amLvs38UGhmvfyoTfl8+tHZfKCgxgLYUwMdDuKPHDaImmHo42R+FqtRIh
Dra0GL0H9jXk/fkURDWcMptPQFvnQAAUHgY0ai79MUBe+u397Pc8mPv93mqk857oQUvX67kYGq6l
1DqhO5KMRcGab5x+oQWr/In7ZbYpFTcXiyEKVn0r5J5vtjBxMJguZdWvGJYMjYkNdukA818brCw+
PYZad4Xz2G8QtI+TIVUNtN5JPusZUdp1f40579yJjiwz9TrgrD5JsH9047TbW16yxKNk8UB3Jf86
mW1Q/BBJiIeazILOmR/qBBY9g0LpgFcqJUoVgXRWYN9Tr6mtRLreYXx8Kg1xoThj80wZ7MQ7rTD9
0PEtdIQ1G+NMvuLH1RhjCBbUjqkR/fjiLeGVTcCYYZo0lNRTYVDlrAGQs6pzQbq4VdLda6JhjBPN
drfzJ5wHq48GYWU+HlYLKOO1Mx9PB5QEPEqzQSvbbWjOtT4Jq81fZ3A+jSFKlwcddJXk2WDDRJTr
+zCvHLq73iCKGqI8Ia975CH30/FOdWWQlUfD7JzrW2kXNhWJcFG5fC9gpFfQdDa/WzcKyCyc5yFL
y9xeG6vbiNpOH91ofy+6W05ekdj9KdUTdHIk+JzjG+WSS3BerMnRz/wiAAZaVFDItfX2KXWT1k76
k6YSGCurSZ5643SjzCEq1LRSYJg8sfKFgBK1HnG3la8gSRgkC77/oSRMU/NX6+zEikgssMv+SDE6
jnBHBmwqP4rCIbhDegbihdAI4DTQnmuHP1scECJXrN+bRP+AkTgfMIXtQrgKfln78uBZ7dLWwp6H
jsvzJOcDivrEmNKnD0puxpthUJiIlG6zJnW+scRQrlosxMRpKt0VIcNfrO2ohZTYgGQvES4c8gHi
6K2kRnh5F7/Oit06CbG4Lvy9zhh5ssu304ijoZ7PZ6thr5tqnJMZWSB7gSQOXEP6/3r+BHGyAQv5
iTr/A4bSatwS2g3Yl//tNF2mCPjbWJi9V70/mt0lzSgeY0GX/caqwbXWMaYym3uk8uNm8fJRnVf0
2lHTD9NC11E/WG3bUJLaFgr4GGlickhLwjWQFI6EaIWqeTLr6G0MI6SRH05X/DFnAIFluUmDERuE
pdOB3Vk3JA9R7iIjeSkg+mya6gAIUmVSJAniV2tEJEnZ0D/9jm0ZHGA86aBogvi2ddz4mrYWOPiX
B1VsJdArmQK8x20IdDkPfnAPuwyLMzAc57Qol8vRH6uPWfAgFEIWxs6IfeVBLbob/5VrymeA4SZ2
qT24E2caYuimv4tfHPgE/kD04HVpKReEX4ikUHa2d0HVNESgEDkUq4E3MJW4vekynz+dwjWj+SWc
69ZSWgIK+KpBD4TFdcppJOu1891ejumuNfB7Ij0o1I8zdd+yOLKY1dI4dUYPQc9AhXakaI1yKzW4
ACNiv/vasdMcwHKegndwSyNDO63wPDapq9VKWZPXI1sI8STnR3lEgh2fGekYq7TxSW0gcYto9Axk
FUdYdC1zFrkkQw5DTe3/SjjsIYzImOScxdw29HQ9BjGveiSjqtE++V27FCx9MzfEEtgyn6xJiPKw
XEwdvj+X4XOwJW0OfDGcS7CsdiFqQ1HdNHlQ41Ima9v7pCI980YI7+7P4UydJ9VaGBFAaz6OLsSI
8Hr1XViK4gnk4oW7IuEMZ4J6YrcfKZCQ0BPLv00RjjQ6H/u5HohTPW+P9X9GARmtFi3mmsFrgjs/
gaLJ4ziYgsWEAgID7WyKc9hkNg/ow3IICrVv1904ikZbW4t5+QfYooeoBtFGy6VtSKY5QRe/Mv4Q
4JVtrB1RYKY9GTkjxXK3IUp8HpFOLY7FP7UdRv16XouVVpbbXr6WSQCLJ+JpGm5KtLjXugL1cAS8
7fyEgtbwIFT8fTBwEOeFs0JPdUOl0ym16zedZcHiIILt4eZYIeOevJZ9zkD/SzOMt813zlx+JlM6
WGEGKmOL/BMM1U82wvHtk8bN4QZcO3w+H9Nd4I4MiNVPu15xLqlnccqPF+nVciC1b6FCkWoBFGCT
raOjRv72vttYErs3GzmYI8f28ssdnS1PV/V6JIA3isWLDEkogCuMgnHuE/e1gGVUmCvgTCzz60Ce
0sB3hKDSBCcr0Pp/hVfqF2NzNSaZqpO11Yx6AYKDw5liLH0fkbV3725/WgdcFL5CVgjKwzmkj27G
jDmgrYTfQ0dnaW2utErM0OeiT7RbNcGEllq7kduqmbLa3RM4jA/sGz3/D5bmdXzfRIUmtd6uZrFS
sMtceuhA24utCoinXyoKyXmjO57MRXCu5B5t7AHwNgsvm0BtnqlcT5jS7tJthQh6xzNtyRdqJUJj
yGxpzSkm9Wn0pa/BQqbI/wruVg6dmumZx9d517c/XdKM3uMdGbHNwtHkKeXgMdryPQ9O2k+45hjN
u2vWqOTtgesqqPxyiPkEyK6vofJhL1EWBVPrGDKC++cyA76m+f/cr8D3Lp2Fnl4lqw3zE1JmtL/3
ZjZScUbZtN9JDYybqIFRgSP/D6LOJ1UXQ6HXZ3PIC0x7PTJX4xtodiUxYxrfROvXWOXs+jciXE5a
udzxf3rb9XgCLi2loy1OywGkV0xSzZxPI3gU54ABOJYiX6mZeAQK3Ecn9b6F1/JdU+OjMBB5CESh
5t0JBfciw3OGPT/LiihhBlCTFKZAjJqunT9iWWtqMjk+5ZSasnAmrI72IAKG+0AO5Uc5SijAGhU9
UCEZueqx1Ok6q47F5cyRMfbKNP/JoA+ZDYGcra2p4D5QeZpzyp4g4zpk4w7+jpsvNCpZ4K3PbdNv
UYV7S6+MbMu0T8oQtPmFuqQLDOBDhCQJpv8n5r6pH+17r1Ub0rUjxm3eULxZ4AJlKZANuOSw6OiW
x7hP7pZG6mKdx3UN/fNgnp3aTfCYPwFAOFH7ycozZ3sip3MLBQR1fH6KzI52FyUO9ASKp+PLROHl
R69PWc/5tHTxbE/BDhWEbdCH0eeKMpAdFOq5gMiX7qGJTnEYLhrxovgurCX2OTfhLs4cNoFBIvXv
YF1paUXpOd7zRr6+nEjaup6iPEeSHC6rjL3X5pTrZtUMbzTcrlvLXshnHqcdQwgr1toOgdBLakrW
pAFynB0TX33WpQA0gFoPCwdhPtD7LP/OXVJDnq0/qYMC5ur7clSJAJ9k+7aC52SKguoo3oMm8taj
WkqbtoIAb2kOCv+plUGyOJP/3MO9rrOulhEi4S20FW5lrlwbsep/AxVpC65+pvqgcqKmq/rJYla0
y0p2ItMPAf/vmbv3t8kEvkrb6e9m3+4lVEMyN4Muz0oPkGEzyLRpR5iVGZ9jGYPLJkbEWzNFP7bE
hmSIRw4As6IIk+I6vWzLs8vJ0yow/iwUkZbvD9oSYrpYTEaaI1JzN3TOEC3Za+riVzI5Axj1xjYT
O8eCTZuYWQdxsP+Tf50qRFZdKmuXJcNf3tUXQt0zyChIcJP344MN6CkQb0pDuNBP3+Cf0KyB23lO
4pV2iKlPr1KmXJ2tfoom3mGOjFNk+65h8kM9qUGBCg7ZbswC+UBsOnblahXN/UKFHxqJIoCqDq3T
tEBsL80oWt9TZrKn29fOVtuGphKt9TQOnZAjhdU/igdiHeWZ2mPN61GwO9WyATOfNKWPeqd0VqLO
OIhzxuUD7mNi7W8sUKLV2wZYwgzLdJaBJEv84IknGRTkk9TJFypGZYGkEc/jKj4m3syyqhYAfcK9
vJU3I4k3GX8XNWjD7xdKdJOH3/lPdKIMKfofeVq+5a2+MhhmW2eslP3A8Jyp8Vs1YSz1I+9FyJqQ
clszcuY/4bQciNp+ZE6sKQi0/NSAll6porudZq9Egto7WoCnIHL7ELA+FtlZ8Gx74LiKe893WC5J
Jg7bh4J4lYamqAobMT13ZcEu2tSBOyMkBPdwm8L5w3VWs8wx6DxA+JsOOn0aB5xqSqsyVIOiD1aH
tJYN3DDGpHgMj5xVCQPEl7KnZWmGL9WrXOHYBNYWdm21+IO0DDsGEduHjoCqmM2tcpL7DFMvpJJU
rPaVF2EiEy7sG/isZZk2pzrd3mF2JB3pNAM2sRlfSdrIaLWtpj9zVTNSJ4Ije1p1iciLrIUUqBRV
yNg3B5nmgSUAfVRu/cGEEr6zAssSer0WDx25yCD/RowZRVrSrURD6WkjZl5t4wBcLXk7oF39x5pc
eVaM6jx1jWci65gyKyxidtvKacKyuCqhTb49cnO3iQ8tacoMAEIVlepL2oOm3npjoE2RNVvUPVSW
bdyLcKKXlmTaOBB/Yx60w7yPyEr54ZZwGIVafYoYxdZAIMIDmXs/2NJ1fBCARrYWJ3tdF6S2A8Ld
JZG9zIlDEBjIUTjUClFjUfMGJNl7+bSvyIk5X10W1fz1aJSVMRJEqxjaoRETxXu+gyw5HsmruXEP
/LFftVWzB+QiWiNVlul5A7UeeULtY6hXPYx2iz1gWGnSpdc/6Iv80Ui5HQZL8A6xs5a0hYgHSEMY
4RA05DD6yWeVvJqkpJLgo354P04fsdtpzqUGHw8ItgfKilILGIMf93yxf3ZRvxpPLyZ+gGXhEZVu
AWQJEjZZch2V5m2kFOqY+NdD+KnyP0nD+kL6XZTlgd0AiB9RbVlLvvxAOQ/03EY2y/YFgO0qHW+T
PkGYCOMFvYDNPXoaz18iuBAeglytDcDZ5Lza0R4xnma0h3nGRgWyUTITtC/XFewi0x21DdLGhL3O
GVa6fQGTEaHfXQe6ndIDcKeQvrBvDCN5STi743z1D889re5DZ5Q+ybeZLwzVfcwzg+jXzV2d6+dj
gI73membHWRYcxdmpX0MfiPI/ItkYwfkBy7nQzkWbSzoFl2s5AngjXj/2vkdPRaXYGfiqUoaQot8
e51YB2DxEJAefPXnS/WIe+g87S9+272dVG07ZSLwq/fuiLNv9lkUf50RUjRKEpKBf3A5klJPSOub
ouwwMKYdiESBufuJDZXRdv+f5lG0QkjVt0qCVTF479KyqqQ/mxuI2Kf3D71Itu8dgJWGrsZ8pZSD
kP1WnUeC6JLYnGryjAzDYsdDavIHgEGvD66LqeyItDqPU+38GOxUGBYpacKczR0zKqJGLtJGYDBf
53NYg5mDEiCbh3kTHTmXmOmxhnTIOhukHuR0f8aifjxUhqYyJPw2na9NrMPP4eWfby83YSBZNPSN
JN0TH/27DAsi5vjA1mQ2MgWEuahIWStuT/13OZrkc43W/sg+BzapXEJA6QpfjwUpNx6CLQL0mxs+
hXVw4F/D29BSePMn/Ij7uGEzll214K/V60KvA8QSFWyzmYqOtQYCTQCDhgMEw67sDPV4Z90yTmvP
AeA8pgT+qB4x3iDkvH5kt9AVU3DcNFmZTu3OFD0xeJgeZ/cpdSr2y3F9AHhyDbqeVObnti1nVgdU
3BLuQsy1P/3wBYSwk4i0J9lIOHoLdBH2krQaMzdoIsRtEKj1ufFvacsDyLdaLRr1F16/xfhV29vO
eSKoLzitIDVTHxDq1SKw5g5B3NS1wUfvTXzp6cQO827lk6b/tD8MobcX18yR7pcxfH8MyzP2YHAi
UzQCAU+XQ0MusfSIt9ZA4nnHi9TQ8ZIZg8dDcbMCY/GZu9dFq3NIl7SZTcdryWWH9OD+ORJ0hVYm
8G1qNeF4czLFnep5qMm1yCPRx2k+THcYw5ZfqnerFc/VgLy7pnWUwxdNTGHYf/Fj9juYfavU93qM
vCgWyTaKARCmWKAhtDI2PFP4CGyE5zypliTxHT6T1nKdXF2MI9hjb692XJPNn7ajEvjABbK3OSb5
l0Tri8j+iBvmi+fO60n7nI4nxJJu7+mQyzK1JgVfkHpQBr9DqwIQ+3U/f6IhV4/0sniRzgjbYiuZ
xDpce+bcFme7L2ZbpTrTMkwwaiXxFCYVSSuR39GUuc+mt66m+iwMAL51nyaq6f25h9YNVBTr9d3s
4D8tnDMWSL7TpOnmm9sMtYFptgxgtn1pRDr92b6/mjQJSZjDCQzedgsIG+aqgzCUWpkJTOF3DXGz
zw7txgS9HDrM41YtN0TUrzst7XDEj5pthqGRf+AbXylzSP/zfZGO0J4v2Dhs2G4mckcYmD+Bdbbg
ysi4w9zLiTGxyJY64nHqLW/Y+wicnsz1Olhfhxc7DQ4e2S1VapN1iFNsGMJCtORDJ+lsNUI+btAl
HmTyJOlirRBnZLQS+2/5RJAHxB2cEswnWNwjdVaSHhXpy/xrm3TXCU1dObFz4VFEg58OSHmUhP0V
1b1sfuvVxT2SPEjnepj6rrf9qxQT0wGA/oqlv6BmCmQ77uID0GvCIKt7FlpCp23mp7sVc8vg5fil
SalrsxbJD8wjaabfj1zwRMaeu3PxZ0RXvomHF7PshmM5y0q1wQ+OfDnpRJ/HpXD8kHyudi9mTvLq
WqkPA6WiAy/59YXzgvGARw92Duf4qK+lgTho5Ldk8G6lWjBPcx2gBPMfIm5UTmzn6pCRePiNDCNl
rDLGwNEmJjC8IU4NcEOtkfHD0vnUcjmdNk45FLxu46vnG3Qf1yXN21CWASfBSe6jGJjRsdGmcqXv
iesW2zQtV9h66QBlIFfWdgwApPUXYV81+DBHwAcGNzkUITmTrP5svo726dMJg1gQNAaCYbfYU5jL
rD/mb1LtVDnPkI8YSsSLJrwadL/oPlsGAhWphQ/05dTtF7iWXtYRBXXbIbJsYpxuzziBxcb9LLp7
a3VOVMvuLJ/Sx0GZW3U20RX/4CESb7nprFCQhysjSFBLIVWwfKUkgbMwOadRoBEpQx3usJnQ+tKc
stQAeXxIQtKUOM0LFcjN9KnUR+RjCwFDFdwvpsZlaFV+74pTWsVf5dn1krqtgTQmGEf2clmBnxju
0FpGIA350sbI5JxHJ9GmIpSoRo7Pz7Vq7Mnr/OGel0Gm2A7C1TYeJPaniki1qsBWIPukV1BQEHk0
HopxpE2aPPZAnY/Oq3Y3UYXTxskmArz27vkDy3I8ttIYu0WY3sH8YTalA5yhdlrQxVTAlDsZWehz
kLNUGOqrU55QORxxN3wsEgAkuXvl02TpJ2t00NV+CAkyEHtlbCpcecoiMK1Ho+PRFiBrxPSQ3ySc
P4QFq97dDaFho0Li+n5gMwWTBi7BwxDdCw0HChiV/91hGpBwvkLLVq2SV8DZz5F70C9ZWfPgu1D/
W5effq3uTF9s6w0MItwVBR5hrOHq4Bxk3UTfBfdaVZI9KaWuxvsCBbQ2qQ+LLHor3B7ygoWfk+DO
9xDN8rZNYyzMrF6vtGR33E5x2ElSlwyp146HC0R3IPRs2UCElmrr2RXNH97qQ88tAfJZs1Bb8AZq
5bEtyYek6ZxskSPuLlRC6QK1OcAM6D+5yCCAnoi7A5H4o/4U4LkbOH5pE4vWOYvQr49AGEwj4cVA
x5MRjICmoYLbtGDnjHkpM+xVp+c5K0ctZEIt03suQwc84q3wSXTCOgnd7ZqMw+N2Ny4hQU1EiGb+
DO+3U8kWz3i0Q+zN9Im/Q30/wQ32FywqgyM4WdfYyL42AcqQ74JYcHksvptl8m28nncW2M1ElQBJ
0g44tnuKV5gIlFOWPdsv1pjTlqP12z8dJdKQ35I/1OdtuekVLpcf70g7tICwQXhLyTPLzBMvB5u1
pbKyGgPq++TvQg8zqBYUBmDokbFxn8itN23Pp14BnmpxxS7vnZj+EGGTpY6jcS5hb17po9luv9qW
/13Z4Q3wkIUfkNeHv0p/rSmJmRGa5phdBnhJYlyoYaxiGjs8PRBvlWaR6VmuYq+VvYZ2p34IX+Pg
BGKov4W2QQ4MpiGDdvKXyBmZwhweASNmt66Atx8flN5ZDnhyaLVK4xc995soX/ATnQ10uPTpXBhI
58SFFLu690ccZjld5PPgN//5D1RKdDg3rdfH/dl9eXbPKzKWv0VK9LldF3VNINq8DqskD44Np8In
ZliUVHzm4TelC3G5Zq8t5/giIhHJnJUbOLx9C9KyFXkb7tbccu6doMlN1HrGClA79gGhVGEpWAIb
Yrzq1yW/55QMsAUJctbN6ys+f2y/p9Mv+ezKd48icWt8EoknS6BNxWuku4Te4XNJhLEwcPeiYJy2
EO1CmWQG+LHNavtYlKwzKLC9h/hP1GVJsoPFMyEfw6fBMVIQNF4v4jA98vdzthjPBuLFHUwa1tus
fq6Fy8qRxQMf8+qIYPulzyZRfXQDMg4ru997rpViYWxv6W9dIvZi+EvzFYBB6A+7PqumflGTx4HX
UeasT+zXjn9h8MfqebU7K2x+LmoM83+fkegwUVZtCzGTUGrIZ7ZECuK3ddrh4G3+vGX2SgLme0wP
262F690wOL5mU3Opth9ocvwT4kZdfDOewkCWbO/YAo3yKrWKd6bDKtAtrh49Qeybwr/0+BNUK3mn
2KbgSmhZumvuFogNTB2wFILgWiLza+vZrZk3fNAoEjhmMVBITi2obKc/VnQkvL+KbSeET3R2tb29
Gw6kSGWRPm/crhTZ0V/MXGvc+bmGnrOp8+eDFXjZTfqGOerfa/DQW3wNZlFsWBxfhW+kkL287P+K
5JTofIW64zaAEQxNHnV360vkxB34mf+vIK2E4Hvw3zNCzy7UUgfwvD/X25GZFGNhjbgjac2jMlRi
2tzTaohJOIUfbMO98EkS8qpBh6S+GULOkPJA5qhnTp4IOikrr2RKNBCheeBjUoppBpMnhunE6NUu
Krexg6tI0VjX82YLdQsZ720zvWWyoBkytz+YXBGAZj2Mx5oQXxoIE5bSr4YyvLMbkQfRm2TxWUKc
/mjn9ccwlL+ZvfOC19D87xIltTFJbQrK0RFJ8LK0uyrcwP4mdG9Z9dTv3xH8/NmfumTJt4gq34OK
MpPpd98S82GNT7994RpQ1D5jCCiUqtmRZdRiZRRtpFsdt/A3ArjefJXUuX8K/cKDfCWN/7gkK+Ap
oB12WUmFIO/tXJ6hjKoG0i8uxLiob9SD8L6XXZ6W8Upw2ca5Vk06O0YHw3fxhOR1tR0pNDNGpuwf
4eYcRmGcKn/ynnDAIHVG2dsVYbhUAAgF8SOjPHHC5o0d/5yWhSvJzpmlbWFuL7mm325tE2rmLROK
6aUZ8z6T76rrRSgUW538AXoTL+0Iz7iN/EjJ4lfxH7FL88+1q12FArMztymje3MyWkA5TF97YGVi
+dteKD3hq6QbAXV0LH5ros4MDt1ShYf6UjB2wpdrVRO7Pb9jSBNO7MLFLne56YNKdMGG2PMvErX9
McEokGY6OLmHIeW141LO6SqgRjhzjEhHmS9Jodd/YIVFzZQxWbk8jH/7GPcr8YJlPjymedvBLQEF
FtGzR6ZEeWDU/rSw7VzJg8Lrl62kjmVoJZ4fhu0Fzt132UbM+EEWYZFWmaysiBW5tGOsoulO7sHQ
BI3/GVopZetF/6bV+88lhblsF6ifxQEiBfK2NNLrWbKXchDMdbX36434ymJBxgSVSjZeki8rOBa7
Ny0Ne3X6Sf1Jafd77faiOzzSS8FcqOhCgbQ6f6I9Xeg7qMxwwQbasugCD2xGkoz0OvAgVeXkvbiT
JmV0pc5VMZMiG7vzF84EgfNy2xX4Mgn6PAPanqN93bJ+XVfzORM7F5HNmDkIINVifi3iL/4oY1iu
huxcajbgG4g/1Ly5F10mVhjBih5DK0eiAUZrBOQAuufLo1W/1yO0c1H0jiWJUK3HP4saWVesQtLA
wVr7/v8D7fDE0KAnfkjKJ2mvTsADOrNoNvI5cP2+G7nY3RzNngLYT1M58n7oG2Cq93RTcQfewjq+
XXd4Chet3kzWROilis0DVHlT1XXXhSVuMagAF0/r4FeLEDWCYHsAFJOcN5BRpIHrVoddkuEaL4y/
ZKMDVL2gsGTj5/ucNA3BKQBEgNXbuTzycZrhf6CD+e7TiTerHa0quRRtk4EYAXkcYvRH72KaA8Ix
I3iYbSjuFCYg+cd1X+Jt+A2uDsLtSRr/UygM5pxrkoTeQZR15bTsF/7/pVcGlLm0+xFeVIAFQbvc
p8HifMtgozuFKV/e0dIfA/qaSx/MjO5dyAtWDWRK9nRM/SrhjGkTcH4etWh4xsEuL35sJP/Os97k
POivsWg5K1fECQoSsGc9rRr43elTfVzvO1JOIf+u1K/KqLJOkTsFJTUfAeGmMh4ZtRXTWGfj7oyF
hN182HIEaQW27IisASiAeJ4tYysEEDkcQt+ZaudnciYmRYOmQ99N7bxxTgJSL//pOHtfEQV2sk6s
4rJlmPXJX43VqW4tihzHUlt9GZOjVYuLEP97eq1NMvURMAwgm9y51boy7igBiItjtUMyMqJePNhs
u3P7V1Y1rmaNOznQajk74jkVVkgkFC19Z5ZaOtDEgTFE/NVQxCcRafw0hNiTlSm7YEMV8EuBzSIJ
pyoXzRuYUtLaQ0OCyskXz+tf5XyxDWsw0K+Q2Fhzy/HMHWw0qvHRA/bR7ZyzgXotnAZoE4JC6sbq
9gYN75qlRZLkEoz86WHaFBp38ixaX2SXh31ZywKlwOcsBW4G1ORZvidm2NkCzmi9soUIF75jECRU
u4hUaqoHaDHSq+Q2N8yTj0kSTwxgOacPArfUe/TU+dPbp67dsqWyXCLcp4XOtruBVOfI4yOSGtEm
IyHXEoCYExwql2U163B+EZLdvVKAJ+zp9/uK/TkcWQWOuYRoHc/d9lwp7eUhEsalNKVu8bI0Z4Na
OpBtXbIvIXBPWtIQeJALu8kUs1jTznuYhokv0B2MfQrgfJTF3ASrC5qDi+SqQSQAME6x9Rkgg19y
3wj1IptPKEj+5tBN42ijizI79L5ld7HIfDGyMBvoWbwCYnKgPv+esdfNhZRprRrfc8DaNKnQiodz
8BqMXLP+0HVjbaRq443/kDbDk/kWgY7rwdth8u7mc8Wa7f3UAnzyTqPmabyJxP9ZoE82IzOc4BGC
HHhipAZQ8u+mUEJaVS9ysc9yGpCih8NO0qnMYD2zzlfc32+iqcUKvxxU/Urm02RZvXyWPM7xBpxL
CvM9Ju16xPlQWJZ2CzK1svg1+wQrrrWTcpIVoKQ+shOKueQXn+2MoGCWoP2qd5zuvk/t8YvyWsfl
JC9+9a2Ii0GoFBj4hxc6TNDfxq0+8yW/wANFVYTpXqQRl5DeCjyWTU2UHQfKYtwjaGY4R3dQksFz
+EYUsM5Lt5V/nqFiIWgAL93fC1N0gqzdFhWQ58KUeyuA0cD6MiAlJzD18xQc3Rdreety60BXOJvk
NJy8ebNhdGv424FoowYYKeb6cpKgfHwBQYZfsEk2yRVLbvFDki0uAH2lRaZ6PKg7mLi3tj5WTDC7
1f+KirdRxNrO80V2vPWX+/aBLHz97F3ckg3slNB5xVgwwSH/UV+r/oQl2tj7MiJD+E5PSUAxDmVw
pG9nlK0ozAyUVx3i3llkINRdu4PgjVJeWyOzFtALiI+Pfc6Nb6GoP7zyPxgnHF0YvT+DScuO95R2
HUlBmqEjJXM2JOlk0QLWQ/eWLXSh2cdzxFuBJpkpcL8nqiKQLO74nJn/oEu+kTheslSFkAbZrOAT
S+ejD8lYaY2QJK63TrspxG85zxgYZRgUv7YvZ4QcUEB2fWBbhHjrXq43kRzN5GIgY01UL/Px1MHB
F6EZyZU81qKnQ3q2KPrm85oT9WW0fNrrJgtP2DHM7tbhNDWQxWdu0BQbrdNjJKx3AfWzYp1Er4Ae
IqRSl/Cgf9XfZU0FzFehcV6bsuzm431Cd4to6ducL+c58z03ernFXSJlsE51OkUQITUdDMdJ6JDe
n3jiAv7ZClpUUTxHoUdjW3ZelilxvTH1l4fJWy1bo7NWlU2HQy2msaqcDuLwnDM8hFU3w/sBmJZ2
8Fi3Jz9Y0kXuDHNk8CfNKBHbxPo4dtZlGhwjGOoYOyu5FeEFaWPoA8WMdomncaa/JAaghdqKOzsM
Tm8ZUx6NtmnRhGlRUh9sWTYY5soxVpmjxagOcQU6hkKCXs0fkEtNGIrzSMV7CD8fVMBkucntfIDo
hQpldkBL5Yzho6F6ldBB58GFOpHMJsUkENtLKLY0ADmuXrtVHi5qKncmFN858vPoS6wTPeLC/DnG
M84FSsQrJNfU/6iAy3Sunos0cR6K/pa+i9TevSFeZEAASLo13FiX+ShwmLNbFgBKc6ldNePglPzy
2U/fygn2HEhpnS1Yj9SCNGHJvb2K7Nd6mZoJBGiX4nlgtBWDk11b7nc5OM+PHnQEdOIXmZSiaA+k
HEpKOoqmNmYS4RA/npbrwQvQFOEcYaGarttdIDvq9AbHbw0omWRgQJ2ZAtQIEATbFJ4fBZ4QK0eo
jlhVOeC6s17pdBr040tYahMHk8LfCuGj1R/97SRahhdMNowuLz6deefcQnLnckxZQe2r0iR/gHsu
stkKd7ZrkO+blsIugT4Gmx7dY6G9M1qTPWwIZcNEVVCwqUOkG/qM0SkyBh1QyBAruY02FlMn+tuw
othnTYvdFDQVS3afCJR6EEyM5Oec+HYaSUO4cOHP0+dOk6Qk3hmhxIkngdfLF7sEQFN3RZ9+9FIl
egvHKlvVOpkfUOHJX5nbHlNTC0ZdlnV+M7Ub2BGaJLnhh8lJ+gv1lCIMbcgqM32mYkulQ/RoXeBZ
6epnM15OBDBmbBlFIEyFfkyZMkZZhqsW2jkr27abOj0brBtKqDyc2yZrlBwVE9RL5C51IZ7Doi7K
QtYGfMH9zNCvUEMJZrdDvQyjKub3mGAPDmjA702kBKEKrcz9WVZIl6KOAlBKwl3AjMB3Kzx4mC1s
v9apLYlRgmG/PnMyLngPglz9YzVlcGebYCka+QKS/+0ZAa/qcyunX/Jwr3azEnJW7LmKbYMUwoYP
Gnd1Xzd3p8MvAqu4DSM/1n2Vdd7Z9JZIbkd9FaG/RK9edW2J6mtfccOB/IbPBJWTr22FDxkd+0To
Ron9bcb7By0LfGypUgBbVy3/DtlA4smviVyxlVophzqbdJzOa9Z1Vnu4aiYDUmR3uEFvLEVJvI6K
l0pvl4uTHItBVBkplOzRaFhbKlXKu06FnKwvtSIqoLXjCVKpZtpHD+mbYPxNXKoixeJvCeUhd6xc
yNMxbYstK3FjeEmx658uvOV4B+pU5/oMaPU2sLu0pCfjmjZa3RJTMJ8bi43in9wdOiz2zud7rZZc
UZwkv0Eey/VM+47N3FaA9jogtZniis3AJHJ9EkWhrxJSH3PnYxaqmhOwy7DWOtr3NQNlbIaeFg+b
xaJ60O1ff3qZPHLMjVGGbY0/5qkS4Y9X98CQwjuRbinqEv3uDI2VPX5mr4+OdFyFag2dVpFDeRgs
tjU9X/HHO8ZYtGLa4vPqOi3Av0ZdxNrwM62cZlgBUqFUeg2QM9urYB3HJmSOVSJmBjEo1DS14xD0
0A1aEv87KJAtC4MwQ1xjd/IKfFhYVcrGpJXAFZ0xJTxEmmY3P0Z662AnB0tnpl99vqqcVIR23Wok
56jZZeu7JHEhqbtqYwzWdVWRg5X8VXUS/AYO9B2TZF+iTZHw3Pqf4lPyvhA4sQceGUnDa/X95Syh
XYcC72Fsn5v03pwbiOTG4eNJZhryCK19wDJmua6M7iFZv6Gx606eNqzJBQKxKTIVP+r5vJ8cJXQF
iR8LpmMS9KacbjWPEHok3J76xUthnqqbLji8E1kEKjHq4YiKfqTPwzPY2CY1BNxviPrzc87yFY0F
tjYyyvDOOlQ86WFsgiw6xnEEDnIF9L4Tn+vgm2BwNnHfIPllyLOU9MM+YQdHThePgBtcKO6iHogk
OO3I+Rv1lQyD8MSZYwjHTNxP/ucTbyyy+SYARlyxLg/O8XNNBHjlBdpZe+KJ45qLNEQDW4RB4N8P
2QT5sWRGtjA09XatWfIWdbmmOZyy/FujBPd4ZIb6zT4hmJuC/rwObmZCieLqo+1e5y4Eq4WaS5t6
WMUqZW/ADyUDlTBBq6w9+6t3/SaiKtstKTOZgfoew0032zAl0T2IkdAfY0vS9lUWfZNA1hKAwYK8
olrh9DA0XJneMaaNeOHiEUAPzrOOydXI+RpRqDh8En6OynHWHvtcYrpsFrnucYyFmow5unRf2KWi
AyRapKP654w8s7O9rNgJdRYDe/lVcAv6LmPO9jXClbkEw/VplVpXEi3DJSholNj5flnBauKc5/nB
AqRlB2xa6FbWhGDalMh0oUA/HJSi0zo54zQ+cOr3WaOvxEjV1VV60GWR8oq4mYPWczahN+OjxP5l
H4lZmaNa+jPnN6wLrFjOHgRf3FSbDGmgiKBLrwH9wGWxBIbCF7vVE4wNJqNDsm7RD+JQ8ZZGT0G7
2c3v1FKbjZGFhsM6vSKoFGK2m2+bEUP9QgFoJ0LQXJoMt+3FZCdFQY1ENW67EApepzobPSMXYrsF
CGogXfXCB+eq02wHq+XikopGfSGJLSLqg115JQNkyKL8QAuZRlS7YDXMin5FRRfYh9TQhy3v5XYD
UrIe/vXuweAIVrjgdpnfZAsq2RqkCvhr0BiyAQMeXiBdbObbKa1s35QL4x4PVodBuGF8dqtfpU/f
AoNDamGXqRgd4O0tdSjRtKb0/8TfkPl46azXo0F9jjVaExCEcom/BccYwSopt6MqSaaPh+hDpD9Z
mjEQN2EGRHK7nea+SO7k8zFZ60C1GRanB/TkGC5WP5YbGh3YFtrSSPCEafBT9Iy9NMd5suw7Y3zT
UrmfW+j9XQocFreMDib4pt3oHgJjKU2ved1H2BziNB3Izw5HUWIOr7kwHphpXh15fwJUpS5mxvrz
FoWYqjMCEzR8NjtC7LXF29E+Tb5AyY+fsrEc2DMrarBoNzz0dBKgQPKCdc5MNx9czp9rMbua3GJU
1SEoUWfUNF7DuzKFkeVwavmxYlldEV4esY+PYCdgenUvHvMy6futidXtn/swK/B6sjOOUyQSShJz
WWUiNQeBqpMRpwfavukAfAngb8zAiMNMdiJxWumHlYpKxGw2W/fARKK0Q4irpbZyYAt5fsTrKAYG
6mmtUcdUaPKthGZg7t5PtUnTNBMpRnqE3W7ssmrWuOZy73MtIv553RazZ01Lrvzi8tn880VUerIP
agmDPK/5REd3DV8dGpkm0k4DCTF26OdcxFZTxn5eYakrsEXHOfzqJvnbbv0KAXF7xu4oabq23c5P
NK4waoFjnJMzSAZT9CdZu6mLySG1xP9onOf7my1Ogxx9xQzjmqUOBYgULp6oMTmnfq9nOk9ojiX3
/a6ko3HXPiaWnpMddIgYqkET/Weh9+D/oLyx1y5dTYmaq2jCriKOWaj18C8smOTL2DGabmo6vAVm
dwChO6YPXeLyuZpWN7qWpghkYg9ifMKXGccFXqyxgDsRb0t3Qs4HdurJwhf0Xt6PjoKg/fMi4vw1
S+tP92OscTCU7+xpCP1L/OjApkfn6oeO3bWlXH1AIlUGsfcurC7K8mtw4iZ22E7m1m2lgOslnCMc
iLC0IvuS2NvnN+UBI8WtZyZzA7lCd4D5vhWFYDh77zmBl1uzVUPYFzxrgE/IqLddZA+ke3oN36+A
ACjaQC59K+RPRKopgb8QKHIQRLXCwFhGJaHSYAYt6cieFj4AOayBppM2D5uFeXyBcFVaG+Yk4Z4O
8LLJFXZU8SaeGe7z6no8sNoMAcRw67erhgHaLjepoyZgwZqtD1gHutnAH451RinHZg3bBJ8/7cCb
cOsy8VnDzr9im0jcEVIk+Ma/FbKTvipi1zWr9afzrnmTRdBPlYVbO3KWPTOwG3kJSBZRwEszQ+Xz
dWZw2hk810SpEzpXl+Lajvt7+LC5UaGi13hQBNej8gkQKzuFxB/QmTbhKo8Gopzjzi+91XD6p16Z
VPEMA1J0X/R/wdHQvYRRbDDmKKpbYjVxvN9CcH6ThECBLc4NwpQjLQGZ4Ac1RgOfrmbiA1XhMJTf
J5uliFAmC9bm1EeIMte+wxQgWZBksAqndA4dpSkeXx6irJVJsOAN87IOhWiez0WUl1ThkDX2fKa/
CXMmkhj5EiID0q/qRlcbxT+X6cPR/D9y5lF6Uco4rEVxog3uOT9yFAFuFCombsQwKYbNw8eKDHNJ
AMSaf1XdV0mCr8vvdaQaoX8hOfREQbEYhSTMsSNgFI7DuIeqX39Q/GXwGNyBbkELin27DeoyQPZf
rdND0qKZrLE9hYsPc7l0HHMjoXSLe4xTDr5kS3XTt/dseycZ74xK3uHWf1JpOEESVz8rF/KxPYHI
vivB070f5er2GgM5x642Kckgrvklfwgy/Qmm7E39LmWPfDrAinX23yDjfgsb9G3Pw1izQIhiglpI
07lAPv+vFCG3DbjSoaeKut8Riea0Dyziqj325eUb8Y89YI4pVjPPveThWGdTeKe2DD9+AsF+fj9r
YJcxIFNYCqZbDHT1e9HiSIiXKqJXR9i7slzip1R/IGCfSpDbYknig7xQgonFFcC7iFmVueWLVG+W
CCuZmveof3lLzob0hr3Slw8ZKuPD4W/JaetqhYC/h/dHCk6YTq3zcqyGWy6gctd/cLo9OC4Tb9Jr
vgXuMA8pxWFODjnKgatnZN0izqZewxGd3sJg+j/tBir5bMIklzsKy70sKIEes1fKxkkPGaNP9Snm
Iq/dU0n+o2PvT1S2G2+E/EkfSQvUlPEVU0uHpHO0xBneGNUoUrCscfedl3xQ9tZCaHphdnk76twP
6aN4uxLowrCaESj7sq79MRi+G3vrrwiU/yv6rMvt/h5j1JoaQrkqWf0xIgCZ2OrUFnDULYnTvz4d
ah+sBuo/BnBY2skUi4WVm++R2N0xINeGJj5CnkaXqNFTd7MHr/ANAouEhpzyS82PtTzoBWqryuGL
9XAcgkI+MukzII2w6an4RDIStGaPSNO6Z+Qfx5jiL3FkQ5UajE8wNAWsn4Vu3T1yHDbiOrjDdLU3
ZgtvaY5T1twtIAXZpC4qVR06eoSdGumWNHpZqKvBL7jJzRNbeH4akpY/J5eVfvIP7A6HjxoQ7ppk
KRuwUiKOJTxnyGJ1B65n99BNumL4H/vLXRwCD1ppRElElKtfnQNZtfeEs6G7Rt89I2QNuigEg51h
Lm4hG2pNdC82uK0SN8JATBPM6Hs8rGrQckNZvD89Wl3L83FNhvk0oPtxOrk6qn/6EPMVIcRHzncR
4q2RPzYIfTdXeRwQU1AeXUUuPmGaJUtyvsS51ifVJvAQ6KbdyVbut7yI6XHfVSi9tIaqSX1Z8dmt
p9KHqrj+7Q05Mksg66d0fTGpuTgG4uFAvI1NMS7ng6LyyrB/eFuRsjZLOBtn7TXOkvj5zyk1qF5J
zaXrkPvPUNJRmc1K2ZuLU3ZFyOCkyOmrTqvIrbLZMI15Qa2oGTYLBnU3yq9T4nY9iLy60eHeIobs
TQkFRgfxMT3X2ySPmENPCKFsspkkOj4/RwQdmjyYL8zP0faM8XOR7Int+6M1cJ0cstHVuoIMp1jI
NPw/LyXNxcmjOTTkzJRoD9x6hwo21eEuYnjKvgDXREeTN2PhZt3gef+cYDizK6AjICUd1YObznq6
aOtW00aoxAMS+mQQC9cN105tUtHvSwyPJ+YAjjZTre4xDYJrOrKinTCeg33InryFFd3zvkwU44M2
h8NwZ5do1jMqeR81O4/FQEWCy/Sk9S/AmX4RTwhCw0LXMrBVwKO+l8GaEbDoa7bAXpFEsLZD69g3
5YZz1ZbJJpeZLj1GU9xbCbbT2+4yImdrfhEbgbohKrihihV0/6tjvU5q+3wTkPcRHnuj/g146q5x
+zQL05fgQHBNGPYsNY/Y0U8xVWIZicm5OvF0Ne7oHi0E2f8MmxL6nNN3FmUOoPibi2PS8igvCZCD
j2N3OCmyT7s8784wwxVZTP02cpe03e27boUa04dPAwK9v5vuWVyQgYowoS2eJpmzzc0kXXrZNf6l
0MfKT8TP2ch1PIyBQM8C0oEzxza1JA82wMOMtUZBxFXw/CM80OQgfOYwgW/KqwcFctUpOgSmkD3W
UUMHKjrgsFfC7ChhDOTYzf+WVmsjxXffOEZrs6h0++rDifIPVNHpTZZPIJGlRBmBTiTaJWdXj9TV
qn+BSRirEYKXzYt4tGAPycW2IgZ6YusSGs+ePB82zt3+IRhQU52z1W05uRMVzDvP3lWDAIUtC1Fy
6NaoaeRxnn8G5fkJRm0ZV1JO6MlhCzmKh5LCeKIYoPaLD9c+WO1f0V1RLOpXwn/qoF50wdlsd1Dk
cxPQFgwGkJvMxfiD3HvJ79dLwE8qYVp9FsesP0tkTbNyB+tXsSet3w7A4iHt6LZGRCER6uveujXB
NUP/YV8ogEVXUk41m4N8DdE1JkKFuVLsQYDwiIj68OzfA+Kuz3j/u9T+eX1tcRFTsLziWmwh1Xoc
55e+bw4Z19nNOIoK+1Zo4AaMCnE1mUM18wVbGk0p5CAGqSRGm6qziYlhN80yoqLsaA+8Wdbv8ybB
NPmv3xl0MeV2y9kl3qxH92nKOxcxhayeUi6HZydEypA79yIi3+WLSmp3GcUzcU10fX2vbEhh0uu+
O1DZguaRRblmnO7FxSqUJ+ImDqB8Syp/JGJvXSWvMa7c1A+tg/Uf5bi88PxAftTW0GqqfzWJMZqS
LTd/Zfbmkc5UmEfegVvtNjRAb703PoQJDoq7RDc7hSC0QyS6RWDKqg7h3dVxD0yVkGlBnsOp+kCq
MgKFnhfdUdCvEcMCIDYozH60bZ9XCvOY8NROK1LmRw636VmYO/oPJSIvQSCmL+/6wfiKI1h5nAh7
8rhNYafip7iDtdL+WsmPm4EX7hrgcxKQCL9sEtZ7TB5z13ul2CXkMJYavypLRRuoFLBkDj3WRa2n
tbDBvuJnq79FRYpKUXG6fOsmAcJXL0SLYQi73+pC51fuZbGKhjtV49xOBaMGiwXBNGNWMHOvRgUo
x795qE19ZJqc1S77rn0rQ8S/QMtvXHLM739Ay/P1nE4yCn6X0ae5Ph0mBQTFd2K5rejmvSSMJhIK
9KkN6+Zbh6Cha5Z25JgRxqS/EaXBdIBZsXCqoQ/bYxbhLY1F0VFV++tN08m3bUErsnj4UUgHaKay
inaFRb8Mts+6KUezk1fD0ppdbkYA/KzFlKp4QR9p7KEtzsd4gR7apOLB0m43wYX4K4fYYU2DRz+2
1AuGkLR84ThJU1nOFLmLOfHo9afKPlGoewDvtCTC9UayUYez0T4shJ1i9nDXbQNDPLZLLpXSYDE/
hLC/tU0b4lssSr+DSEMSDIzMxR9cotTtB/2gGpI3ws6dOKtuAqPUtNbec4TjBSa1cvw4szEU83yY
TVsKFB9drlsE5NDZ9eULySY1prA4KxiDEzTYW0kJorp/MaifEmSHyyJPVlqbulNryUiTyLSrQ0jw
5/LgJvx8M0AP/nJnfAgnRsA4YJkcgg23K0w9O0JQNTuQqAHyZ9FPA/vMtRq9EaMQDJvXWhecR4cg
z6Rrq/hmmI4DI5by1cfvauuWskLERyFd3/coYqipHOHD5R3YDzMzm7bizUI6l6zojJpSIdgHy8FZ
2L2+y/OxRvzdvzbd+u3bQrIX9Qf6Q6GLygOeN8GlZAW2h+fqnNUOyGXUZcQag27Kh6zy6vWkHx9r
7XM1q2AVXqxXhvtVYKxFQXVhNR70dd238M0y6ARYFNIo2+RPmjprkKMasYTTDrfwdGA92oz9pLLt
jUm4GrJ3it9GNhJ9p0eWz+O7Df4LsHdJXMn90NAb7L7y+E6DvVuq/yPEMvTYV3qzdMMvgYcTkxmf
zJQsBSmvyDfkysmAPF93P21DJ5hrwQyO4N4KY23s961YqeFRd4Y6aNW7xHUX04049Hmcg8rdLjop
97OI327qtqIdKyh2VSqXVaOn3Bk4EvAaQCfWQPApjKdQs96ZylLCBBuRXCBAu+Bn+PPC7joltHWZ
QfioxRrIujxlbNekiDsZEHxzzoiRKwAS90O30sL7dcKihtFcQwQrEtvkle/3HVPoWvoW1L/lFxHr
mHlt16F+7hriIdlF+nqZfNygNItIcQJrlEugobdMDHb4nL4IDbuIp+qS79kqYGNL7y2juMiMAuNE
6hnfCmpzj06awAmTW9wnkn0J4j0XfNxJ+8AMwOJTXYZC6XSmZzXs+bI12Ow4LIdkCNO2AYvUHqXX
6YDOY9hHDJDiC1NB7/UiznU04Oup1We5ZPmg3kinu4Arb4vjBYzzg4IAXjUQoTcaSCoGZgtVvzvr
eF5r3G7Y9R2rJjAkgYLHkGlPL/OtBo8StdJSA/InACyI+HnToFYbZg8+GgNpRblS8lqqj8PZY2Ld
HWKnXekhUbGG+XCrwwM6Axg/0J8Zsei4v93pJF/LF78GmpQqD8xV0msw3DKJw+WXPd4ohulS3sAQ
i1WgMkBQNrf6MdBxiUjmMGNkY28gsOxc7S7njAL+K8b+WSANtRh84srMlzZi3IcBuaRvF/2113Ao
2kVfnWTDcchS+hm5rp2qYL8EqXJ1dJ/LbylwyW8lUbOL2Vhw03KD9RhGDsNLGiLXXhza4rqZTMJX
UzGi1XWJtiZaARdiSsVqpyjSkqkr+OSz5GphMhUcaUrLOJzJEmDriS9VfgGCS+Le9cfaoadyqE+R
KyFcPcloDIVho0De7SzRILGRN+U5OJEamymjcnJ3rmRGiE2NNV0Pkb4t1ud8CsausQ+yma6TW3s0
VylFZUqQcFnkUvpzW5FSEwG8JoS6m/CaWwx6JIKjS6Y5cG5ty0IN3P4/f8Q9ktmN7ZLrut3HCf6s
oh3dIGRg2yasalbp5+5N+h7Eie8fs0QKYV6JLymt7XNaH0yFTwsN+DIOjyS7eAiAlJqAcYs+NZJm
Wpa5A5wtoe6WY2P7Rqaqg/VbM7fZOPIs7aP2kvBa8f5sKDSXveQbq74qwaXiBygKKUcW/XpbuYQk
/vGBl+dkniAODx6KfMGe1ir5Rs5svk79YMxH749z8rz5RtU3HjhGd8p/1NKxSFcRQpws+h56voF0
QsDTjI6BJAc9j9u3rWnD2AlgxSjdmpSsNBPNb0JHfnqo3Kok7+nMIt6BsIGD9r3Ew8MAkC2XGnJy
VMnSuaDyUch9aNbt5sREmebSuZH4SPX/cy12BIOr9OfveaXn1bue9U3RKJbhgpjGIg+LaO8oj+eU
N2WEhrhnZeHmK7xdpnNILzJsS3nC4xcLcNIj7SbWByZQwHNQpY3+XFi4h+eSRPTwEsNf39BewUen
hBLSgGz+OnoJXCZ/UQdqhxcDIl3Y0rYv0p187o4lTho7+T/yC/DRF3Z72snwkXNgALYNLL+xaB+9
zNQCyC7ZnW5TAh7OmM9Hew9OFHZ87Jm0d8oFE2+OjZFmyAUkCKkwdo8FTjktSnBV2tqF8+j2TW9T
L8mrhJyaUf5Hm38TROxs9zwCASBRlTlHiG5dDrOL4ydeJmsvzB/isMAAf0+ae4dE9RRctyCBJtlR
Gn8p5fX8GiJ2ut1w8dutb/KGIHvBqfM+B2vrMXRR0vpFBIGSiol1+olVkV5PJTarv8DhCRkk9F8T
7l/iHksNfxtvxTMOj8pF8t9tIMjY49ZWNucCWEpxAX3lq9LVMbkHVXpYc8aGb+p8OGGUyxhTGLpg
9I8WT57bIFBxaLV2FnVR2HT8xKcllTMyGO5mShHjixs5b1BtLT54qXhRok891/EJnvoSDdW5GZw6
ZHXT4nrh46INWfGwK03kqqmqM1ArDBS3OZ83Pt2evx/j6svmnchLGg+9vMjg+dmomSUVh/4/54KN
evAey9e5nkX6KBktnDXc5o4WKAhVG7eku+C5FvyVr9HyIkEHz00KbgTrSFkJSSjW9mG8h7aumWnu
BGQ/WXeAXQMIbfLDRjSQT0MMQNM5H23p8SPG8hRj3gC3uNx/cgTIu5MnkE1Wq9k+OrOzAowe4jlS
x0Y6477+MrDx9Eh2drM/c3hHSotgdlRx8luWw8397xIvZQT2kwZu4v3KyBl9qEqZPsmZ0Z6soZNh
m36LfEWvUbOL+3JdtEtbGgFUi//wZ/wyQHF/5BlR89iFAauajEHS3nIgRRp2ATuhlpS30TKcZ1iI
0D00mQOiIcXccjEpOyh9XbBMnXe7M0Kt+JUxX3De9q7xHWsH3S63qR9VOIeBiJOEleSQgkVW0Shh
PgpBk1ExQLhkVl5eW7pALk18rDLanDkZv1KhGfIz+MRsXt4j2+UAXPdB3g6ok5iSO2gdjif0uVn8
WfteaYy0Y9sWwredlQDlhITAhLGmqX3KNXSMWlcXx16MFcjoDwxAAgNMfsr2lgmffdLzQC+O7R3A
hLnRQchgtzrSyYVO8Dki2wbfq1UX8a+ljsEk1FmoG2fInOQj9IG0Bp7DkLDTXRasROp+zfzIpOSO
BSlPS/X/1bHVyiL3/qaoZa+LcuKoBwZWPzsGZ4QWulrA4KnZxWgSiy17BZTXpL8IiWLjfRoN8jt2
flkSZHUl2YBnG+4ZQ2M1NvsiGARR+O1fuqE1eXC6JIsqp5cTedTlonrxAwEgblZ4t5yJAqUd68zu
zZJqUxe2WNJRmazTFsy6hZeJv9fGPTFcQdN0S7KrKGTM4oOn4kqGRlB1ELqab1rmwWP25qa+n2w9
3nisGrftsABw595+4RHvvvaE5GGvQUa7A2HG/dgrukP3Q2Rxm6TXicFQC3PsqE199oip9VPfkkhR
tnAG15kOxexzfjTyBuFAytyi1VtWuTPhWkSEzNx3MmFKO5N95t4g1m/3csIHVGGr9+JwzGCa+Z37
Yk6qSkDtRIA3EwSIA+xxB8ikP2jL1FHdWova7sTt44FAeBp0H6f9ZBsWvigsLROLX3olEczHcMnJ
NlGmy/HPlWKQxYG039QYXJq7XuIHisrAMwLl2BQcV4WXxNufcDc6f5pLr8irK0KPAshIUKGLwpPB
PYEIoFvpNJI0Iwut675lwfdFd7zH8br+uOA4+/AuyZa/Dw7NDFlLKEYiBYj397h1vACLt03ND13A
S2d5lmVbmrPnKV2hOHg8GHTe5MZVv0Q6Kl/z8eVlFohLiAH+hjxdJ4loFkbGKkpUS6WjZdlfHL9O
sX3WyEKFIx384xD7458fhfYpDMDe0Yd5WFTpM4YS9xr95oCP3TibyQ7xQNBmKs5jTYXrnlJQ17hk
YxbcH2NpdwvkH4R7t5ypsESdAwmmkoyfC/CPPRrNwhxPwyjLZNu9pRSXoGPqieWnNKN4rA6j2U8d
EX6tqVkQ26iKEODPd8Zxp8h+d8uT4MKHaa5ImDfh//H76DzQc8pgRiSrcinoHCkqBA3xcuGMA+Rz
W+sL6QkLAi10hKO7RvOHZ/3y8nVs9hrUadXTuaCLumDRKNw5W0VB5FrGOhcO9+MSQnUQQeOQwqha
10fWarn8vQ4iLw/6BB27EIasyuNpmFJjKXa7s6VxlrGlJQ2tWKMIArjW6f9Xh8s6wNwjCt8DJPkM
sKumD6OYJt3wpv+hss9SsISgg1p9vwUpWPXqFZZpWqznX/8+gnJ75SbKDWyEjX3Y0o5NY754BS2S
UPXl9ZIV+dJQmI7DtBR07lB6noCqC9Zk3sO2jo+YsMf8bRL6YcE5jNzZhpDR9hkK+pQSduJM2xkg
xCd/fKBxwGmRZmZL4IYD4EPfiMTP8LZDj2o+gKghPddv1p+nX54s7FPqts/d0YSuIUuljuxdwEPo
dVMey2yKxR7nQPsXxVoD3eZ5j5eImeeqnzsvdHA1bCyqGYnUB8F/ppOkW3yjUyr1P26XMGCyDepv
8tVIGOw6gIAf9sTdUsyYhj6dWk2gVWFllj4QuRf02UZusxyHpdPMioHMJHhJCeTgV2sWpLQvl6hZ
JrM6KZfWsJHDwuj5fKVSJFzUNdgh9miZ9KBU9tgjLbaG8gSGwaD6tNFskz+6dXaWXzffqC8Ttrli
BvryMEjCFeQZiHBrmjtgGTcWJbOHYAkEVWQg2esM79UZcvO4HSPdj5A8yYJMRD2pnVYhf4+0va1y
WPkHPKmutgX44rySyNiyOhvXn5KbCXfyfSTgoB1PxiOe0lFxIYZlyWttl4HX4OdXG58DxAKinsVu
kF3QVPzz9JfyRHzTbIbOmBx5rIczarz3ZhHZr3R7eaFHmO+ijUVpPEsam8FHN514wvXmaJyRVXjt
4edWuEBtaNmCarvm5TM08MZ2nHkIlV8MKViFBNlaorBRuKTJQh3qiomQ5IEro/91NoVzPbrxFq0y
qFjQ5ACKujBEgz7rZok+OY/J8kr/nOg7sE6a5zqnoWFuVKMZvB3khkwE8zik9mbGTOS5R6AOMeC4
u9H9NFZTcnz6cn9LoAd2qUVn5qYbMQS3u58bl8zk+dHv7M68KdMj478ziHFCGCaYAQUR2B4v0+6N
Ru4NMVImbWluRBmgZph/be1mkblJNII/AC8QluCQA/x4xO7ZLOtAAaKa81ZkYw3fyRfm9wq3C7Ew
m92OX1AVcY1gDdtJH+kIlqqRDTTPpK+xqK2fFpYuwY4EJEozXzULyPA9a6oE+Gh9l3qwkeni6pxA
4zXR/bsIAr/K3M7HLH8S3x3kIS1Z4ZAdNZshcM6MIdDP+edxzuea1CiKkGSMl85im5khCDk+7J3f
esYQB+GoB+hYDYBajzNvHUQyZqAdIG+A5FL0B9I10HAC+C93jscmBBqDfIkJ+ULhmLFiAc+eT+rN
lDs7Tm9S6V/VQwX0vL9oOXiyPgDTVkxbSJsr+xKJwfc1k6Y9XHtXe+FUpUQfBzoZ7rTd/gerVvfp
oF59xm4Sg2KOd2HpxAYGZ1YL453qSpdRIOTjKETfV3uIhmA9y3ITYTll03iQiuzEUWeEeMzvWehm
HSWnqHcQUhQ7t1Q+5fg/g0VBzzZXtDu5UqBvjtL3s9cHC4GpzuIsdRBbXQX7olpXP19Xn1iSVp7A
fWyIUyoMJKCBTzpJDPkr5g9sm3/TxxvS8zM7BkaKU4Dp6fF8KsTwnYGUjgbr05UTXHzECV5iPJEC
dfcWnhLv3URABfamNrlMxU6915Qtv/as/s2MczbgMR5bveBezbSvh1d6zqxfHvYluiviMAetdkkn
Y32U6rVADlq9AVCiNUBIsaYT3YBJ0q8vqd15wo20MWCrqFKc6U0xLWUd87Pl2akaxGZIS9B7y0uM
BmYw3Kmv7TEgnVnVy19Ir2vdHH+6smBeIaMp+ai0OqSoryad1kvJrD3+314nHHB5kP73XHDBIv7g
jsJQ5lYbTvQfSqeuBmPV1AE4j64zrV9/1BdlnkWYquPFH5jCHagl2iz29vIm3zi5fOofAYLrViJ8
s0Y/72FmE7BoE3WqhN/EWMYuO9EbZqQih6o2Ll3qgR3/hnDqIgM8yXKKauJ7bmDAcOx43W8lnXa1
hhP/YhfC3aEXIdliPtZ/7oCy2EgPJE/kD4EYFlqnsHEQ2Rsby3c49z88eUqsRtYtuIRID/aOcLo8
VJ9AeUB8q/3ct1fTb52UcYiEZ8BC4jQJCaF+fyoXskMeMazjbdWhJRgnhoTnpAB+O8cCOVZBLIeI
NwjjatGKEsEsgTQug2aqCRe/HetHYpY/0GyBPeht4WnK96CsOFWO6OpWMuow3eTESxGAuO6g+/u9
s0Heq0Om/ZE57P+L+Xaytk5OUoUKF/CJnJG6NbhuxMIwCyi9sBQ2AcCFyolx0fG2CRC8qSAU5r/D
SZ45hT+MG2QrLoRWVq1qRAjmBejQF8+Vh6BBN8OqfEy6ue24ncdjSteoE03ks4d18RxQdMTE5WvZ
1iXysFBHfnrosGRmORlN1+k0vytHULHFELgAofyVUG/MYnBPJH7Ttv4xBKR1Cz6ZvVU5AMCbkmqa
Gr7HOAAO61UfcGmvDGBsVgnxAS7HMI+iTlWv3Yfc80xtZ049jGcRTmkYibydZvGyMRavAd6MEJ5Q
qVbNfmKu/ZFlbO25tDeztGBHbT+gEQ46ISY3KhqbTHzwcz2HuEyd++qxV2R4ZhKQDI3/J0+by4ND
Opc6FRdC1Ay6v6KVuGEi/18UzKm808Lu3Dsyj4JeUcUnessg/M4JU7HRchiiz6fjW8bYdiv4uwI/
chEFt5wrRh3MH3kqmzCOneYpYVPNHokNhxbMZIcEoLSlWU8YR+udOMZS3/0kJE7Xq2yEqyhLXJIk
kVyL/vDOkmXZSR1FeiMSSyGTdjnu3f6fa5rG01WafWQvT7P1awR+ZHPmquI68evRnMuHyYXgthuc
h8k/ir1HPFKlRw8iTsRQu5L5XWaX94jltfyS7tx3NJ6cwacbBotCFJKmm5/I83o9GXiRsOb++6wG
mGLPdSePg3c3GrP7M5bRNjC1Gsf1uDiZ7L2ERFC+iJL6siG+rJGLbgxjUXywOnZQjfZ3Qj6vx4dI
EoJEe2JUWy15XwS3bRHGCPlCW5z8YkZo/h846zPLj5iq2ufSL09g02uMgtyn5fCeOy5SKKjIhkRw
DAz9ZqI4WclxctKMqWs1C+hhfLC0kmnABz/5PR9+DN2CLunQzlQOAoNQVpmyzU7RCd9JTVmOdayG
tNg1fP9KEYM6QhGfD1Fvl3MO981E/3rKKBRHKVqGb62S+iRmyg6XsKu1vEcv2y+4vaKF6j0KrDyc
6WzEQwUyZye8n3h5PrU07ACcJuY/hLVrC7NLuUGvJqLgcUjdd3ZDkVGtyogR7+W/GO4v6NvyG5hB
93muCVl/DrPwElaiZ3U+h8ze2kFJJK+Jxw6ebOswmYM0dZKksZObhrwe/gXU53MWJvQlUWLoJAjr
wJJI0QPAxEwXJ2YRPKiZ+0dJcHxknbJFEfNxCwV4nHUPe9Ob6unFk0H6zaAlqITrt/XQyee9YWS1
xv465Ba/Uk/yHu6vCXqNyxwG91Li36Re3dPpAfJEwKUBYiTaNXBWapppEiy//PjsuiXevKdecBjX
vdn2eHEsz6IELWL0ImIiyswmrrKCMU2UoWqGRBQJepwirRsP55apUMJGzgLOTNWMQyr00F2mPJA6
j+V+MdnizBJegGYp/at0Jjsihr7WqkYcw/SOnVx8Qqnn9JvylJU4SINee9hj6x2bBleAryFET1aH
LkEu/LzXPOZILn/u37KAcwgiqo0afZJUC/noIwW4DxPWCjtosO/rRh3iNBYFELrbQV5ajhjv/Kcb
pGD1S5o5rsDv4TgB564HdQVQH+vPpObaOETgxYU4my2MOeP1YIe900VRLIDuQEIMaY5QVFc1XKI4
pCNLSioFjAkqeJORYxiBm30SboPP1r8y4wwjt5aUJEoYd11vKEVd2vy/8Y15FltcvsJODipoLNNm
318SxfwQwhTSYdcRonwfSpTRNmol3kjufMIv1IZ0yC46NCtX3GyhRAZTDNRBlnCqWDtbSt6Z5ypu
i8T2JSwFPz6+57q2reg00fh8RgiUPFXqcuh7hMbeI12KOx+D1JqDg7007TFH9N8dywn2ffm5b58V
e3Se9GwN96rCcbjKkidvJfvEp4BmbJNWBjIjQ6qOmNDt0Vt+IGKTQFYeuG89+2toMQNkbew+jBmc
u3+eHpBZ8P/iUHM4o7h4gDQnIBGDt8Z8brLq3v/VAwLKv+7RLU+fZuDbeZVKtinwx1l27XlFIzhY
wcRUbcomyWPQRIG2cN31xy0DSDVl45cfjVYCGcvuFX3EkNYBYfCNKFjFhUTvlV5edQYqnEGovKKU
nSZsp77fhA9iOSjYPLJPZt7P6t6R1xm5LKX0sggHtJjiFKAOZZf+GccR5WS4RVUCMfskkBmDa8lR
bWdFs79DRurB6wxAbsafc5G8sRU/2az8tUO0380kq0+nTQdH65pyA2kPqa64bAaFZPkq/fIvK8jx
QucU2epR1cTaDCIlA2qnIQLMjGL4Z8yjj60/9E9//i3CnKVURAklM1W+tFIdjeF/VZPnogNbrifP
SWH+Z4QA7UwSf1lE5UuXkT8xCG0ME9eBLme9RLZbakPaBGdvxR/FBakHZN/f29unzNqyzivXLoaZ
T5LlOPDxcxtLSSz0KGNXTOSaR8p7iI9j5zPvjWhTcebVYzud/15qJEtBgJgtU/KQe2IxzoK0hSYZ
LPdGvfU9jvjPhfptiWa6F8jKuPcxZ4wZU/yLSYTXl8BYlTZ0EFxuStAtFOOVSO6xazF9WA8S8ie+
8xocBtwJCkRGknROhA2V6cYLXPzfCb7DiO7ycoKSiTVd+gIfzvaAWP9RF+4Km4XY6xwFxTNF1KoR
xC3PjJZFtxxfKSiLdcDjTRzWNbqjpen03+KBJMbhPY2OH2yfZAN8ImKbbI4dk8RscHoLwi/ONU3A
kl2oPErl4dGG+dHBJXSU0Tyn3rLfCGYxZ4MOyB55mhzYQlU/S1apUSx6g9pIeXNE+GUFIMAq0OHt
JucNDg5OiovrzuQAraDRPwJPP4axPITz4kKIUtAdo3grXe0l2PXeGie7GSp5+FP8ewhVeOtHybHx
6DHfZYlHIOCoBzQ2eg45Akvqd1Zfub8pHebe8rxS89sUOpBbz077CBePB18nKsGPVkeAR08bBaCE
oFbCD/9RWvhOgykHrBA1u/Ja4NiTjK58PyM7sz1ZQpV4JcHW1vS66emYpLeSSJHs4fJiWGRhC8nc
VQVH4Q6wWWUwAgN5xylc1/dsLyfel37289XwENrvd7KwoFJ9Bl7HSUICRwE4A9mvbQyxkVPFwt55
CuGIRN9eAboNt0GHopkaYnlp+RIxDziQzydCpEgYnwDBU7eMWc4TgQRCcJ4a9FLhc8QosVF94M2r
Q6SPu1LplASphXsDIxb7DIFOoABDBup8SOAYLtN3O0XTVrUX9v5/jxXie0uKJ9lFUEUX6xeBPyq6
Q9QeaZ76vvv9kAdzJh0VxnVu3j9U3v2osk7yiCB4NkEmNsG2xHvjz2APGPUiMc5EB+nWtZrUYxzI
mDk28+3OZ0VJotceSklIodcgQGRAcoU9ZaFVM6jbrVtmtatYBd6/80wBT+BUl0CDeCE7DujoUyXl
B35d1zubFwbqPP7FISJ92mYTGMj0x3uf6iXJQBDbviRBezFXZSUCF6kszUjMf4byGNQiEeMLaZne
WOHNUUMxo26UayojgKfmVj3YNx+d1Yqjm3JWVfHTg0im1shTufvkrkLzSFePNVOKQ9J3ptet5GKq
cjOdBkB2IhUpC9XPiUA+ONiabMF5OM4OVYPc/2NUA10UiGwTe0mCWGIDd0+6zWE4WHpstoIxC1PF
dR9LHqHo5X0rwOtb4CweC3JnUfWlnrwQoIEH2/4AMnMTbY8vkx68TMvfsraxcaNX/0HZIMr+vze7
ChJ13pH+v7uW89X13tD6W43h4ZwkccHhddSU+a+wbRDtSIujI3n0sCf0fqeYnnoDqIT0D7rPGkKi
uPiRxJKTgEp98Vn8wniY+E7xbdplTTAQzGmEETg6N9BFpaUyoakwqRyj/nA5PKit+H1svyy70L5Q
tmX4wTU/qT+i5yPGFcQBpeWETSERBhySXlpDUi6iRjaWKgSTzc8YFKhLH7l+jPabHWzDHZ9u8zE1
Qs+oONYjzTf4BLq/U+jDkv7HBy4Sw43IuEqeIUKPk22zrQBjRFH9MCEXEbvMXBua0GSqk3p5pZlD
XRiuJzgjvu+55xiMeuN6A8oof9UeVd1TApP+mG719ym27XK0FudOoBc+3Q25gMKHhcKQxLAZXG+d
aydVTtzsSq6O81Fa3bz+C8+vXWWA7uEVq9oefivhoLHHu6mAW/0pPIEDPz4gpOhpEJfVtL6bONbY
3JCrdcuY/L1WY4bmGthn9t6QPoRnUS0xamtvnHZxcrEoe1VUBRhiP3VvilWkj+QzTRCTkaaKf5OQ
F3zjkB4P6b9UxF7B9fRX3a1dUmTN2Wazo0Vc1OKK8lTY6+V0HJIF/FdvEuiBT+VLc8N3SIKFj0c5
4I2h/FydCv5agODJA0s7f9+43jv0FVKVRFuebtF/NISPMvGvkJvxVNryoGzAB/bj25WEX7uofayx
SjqRoGlClEZ1slAy8gZDbS5pAWzhGmgU3/W1R2LKcyD5nwPFWewa8CP8c0hplLHiWd+D1o/mJTCT
zLhdaZQS0bbNdOOgHbawsPY4HgVlacgAUdFw8JtPlIFuWXBWTQNB+w/jNdEZ+2ljrutYrX1vRUKO
ZJakSOfCOpQ/5X/Pumq1COaGeVXCnKxG1feixeWSBGtHB6nekxYb+40pHRfkSQc+oT3oB1PJx7rj
04zZUH/6mfL11/75CW6f8kL2FwrFxZc0DO+w2JOUW0n2QiP/P7WuWG1F/wHzMO4YRsP+UEwmZZEQ
bMPYtFwMjCC+9omzVYe3nGe3FULT7LTxsew/Zmjbmzk9Nq2gku0wEz1H57wHwPBpZH8TjbVf9mX/
ZUgp95u2FJraAqsLjwH9jx+xB3JTFU/JUa06eXH9vK5g9xLeHDbnVJbQzKrO+cJ5hGkR9zxdYhcy
WXQygtb6G3w3eODTKBVg8D5IXkPhp2aq0+mgXczxS1dAg39PWi2vF+w26J2Vvrqan/D+6vokcGWi
doFRKsJk2L0rkWlZqV9Aea3We5OmVdRobQzt57Gm9c2JNKqv9Yr6ftTiL1VK8247QQUYkfaH4F3s
MRF1aOuUPrDvyE1ssuCXxB0aVNokWgUCKxpbZzOSpD3UyjS8geD/AaVF1ZaLGOZeqwAgWtIDyeMQ
frNZNppMfZdCURjDFPl7vf0BQaWq0C8Lurt26Q/d0T9NBk43av+zqZNdjPjV6xfTdjkPvrbqyXzG
yQM19DN6HAKipTo2WdAyeI3MVx+Z266rekz8Ck7ps57r4tdfke6WsywxoTvC+/+RpSPj+nTwLpuH
aBAvcbasNp/r3CQM/Vr7B1Lp7PkwkWOg2MhS9rZz9AkgM5e88HVkoZuh9zQ92N4ei3c7RuGaUeUy
LygdsEj7XuWO9B4ZHGupvToARkSDSJh+CrFV4+GJgJBXaJnN5EojHwadwq+kmnrCMeNGVv9PwPKQ
UH3aijOU8PuIaNY5dPC8nRR5WIs2sjY5QPr1+dJHToteESPTIVVaveWJpyJo1x121QSFFR1ranXe
vjH0dxW0w+j4U4DpL3zRt3+IDcG8ocK9apWPMiRHFRakIz4YQb5vzqN00oU+5Yob6vzIuDZtqUoE
A4PFAgM4yMwk0ZeDxe6esDDYPz9R+/wOmKiWu/XfD3nXQlCNG0/94prmDXtp0IE/q4QhSRXW75im
9w6FOREosy6zCjmDO4qRJxb9tg4sjz73KZH6rr71+WupoihuxSbSsAaNCuGnnwrCqnfqmTYkjRNM
qKIybAk7cU6W1gEii1idN7Fugsln4cCABvHXDPsyqpxLzr3rUbRZxd9UZceMoU1/7xP7rRaqTW0Z
phV3Xxku9UEEVnyr4wAtGON2lvR/YPqq5w/+DEFW1KLPmabI0gdo4jhgrfm4D/N6IF3s89LWUnL0
DGKpuOz1QYBHyVSHR4A5hTYnh2pajfWyfd6/MEPcPRnHoR2sMtvi3r569VTG4j4ZV3rxqeJNepDB
5kxKVN1AkBdjqXgvbfawQKdmfSndrXH59bPfnKGgxBvP2K/h1Z4hAJLxKlwU1/1eucRovJHniaF6
mCjIyW9koia1U9QhgtT1w4om2b6viVo3Uud+LBhi/EGhjene/aQwqckGqCzrRwlrWaCTR4B0Fh5f
RupG6GqT2l/6lRPlnG1pPnyl6/eCmXM1jIIp+kRgeKBg1+NYb7q+rvAAd92zzRK7By3n6RnOjoV2
jhljxD83s9OdgKi1CXzYbpEkRLZG60dEF1YxkOHeC3q4FmG/0DMp1d2NiQ5qZ9jNjUtjbtC+bSir
jIMLkjVxPWFRwgLxDcUzZx8vqeaDmjU2aDcQpoBujDYBQTOIDVjlk/yy1zGfUe6W1JRq1yCxN2hl
/77zKuGT8/pmkxC6j5KdY3GGemztspKwVXGny8WjmpbrqvU+kvMWRs5MpIV6mrr/cPsWnuv/MB27
BqVCptOyZ5p9Gv7aon0oWZEu/5DOZLA//zGRpRhzM17NtNT/z9zvFQPUr5kAf7g75mjJ5A3nhan5
mUhU5V6G2gDIpj0HYVNIdzAfx9mvTtsuUWocyTac1fZwABXk3pafAecib6Wdj7Op44kaR97Tdcs5
NRkNHwkdD7Grk+YSp5QVpdF3AwaDk6n8oDnQUTWeJDrDQKOQNPeHjTxr5ei4SJhqEu1IHmgwRwOI
quoVOtNAHsVXfCjsb/fes0T+kvmyxDY5ob0vtaayzv10pIyLNdEScVw5gV+EjmlOLHbiJ0NP6P3+
BdeNgPm69J2m16nvZrIQ4sRFjNTPR4VYJ+sinOF+Vta9U7ZBjwhKBX0HGGGXufgz1rEufOHRb8ML
fy+t6PS1bAztb095UgDkK4OZnzT9VELCT21aN8y/xBIKJSHUkRimti4/iaLJlfpHEphkDqp1x6ps
xRKD/llMtzdbTohRJaRc1wwNisadeD5VpAlNdkGb7nBMIvmaoFIgkf1ShqV9axsRvMc85oqgi8SG
5oNPgASOJz+x3IHRbeYo5yRngnsCdzfKbguwQLsr27HmitCUnAL7J2OVs0ErGxd+RccygPe6pUpt
o3mVH0zyV2dDAqyDlLTaON0gZT7kNT0K4/qvzgqIxJPOrig5/jRwgUTfBhdnDUNFRaBtySBSUAa5
MZcZcZHnYB4IbRxvW3UkTkQoVWlVEAiTE9KuuSadFcJfT2dIsmXnDrDfPBggNDuUXxo1+ukXu+u4
8No7IZNNxL6TTNRGmXrVL+8S702smfg+06aZu8vsWDD4inu+cDBQeuJ9Bd2u6V3RWVSI1so4aYKV
vKmBsaCgUuvMx6nVqkBE9aKOPxZmMCceZrbcCPLvgGe2asfhajzP3ArVG30uNX0VGTp53ByTvJm7
v8DU0N2GvDz2HqRMX+w6eyvXGujFW8i3HhQIqJDKeGES/kzgP8lvMGsDqxvHuxwqyxxmW5V3WXC6
RRpC9cbOuzOvEP5vgcQscBQW/Qq6eco4JCkNCI4qPV2S3gNPDNmQKZbH1EeVhFu7jnsYRiqDmmdv
ohQ8sJx3gUR22lnXvMR97EA7tf2yKshrZMfKHMA6AJR3WsbJud+vvi1qZOx75Pwpehdjs6PbWato
SdjYMpNcN02qJoaa5x0HgEru8HTGUep04bbaqLQja+ba8W7GJSQqel0czpEQqLpW/ukH00M5H22I
9itDijpRwTHaiZJ5A+/L9yLVal2sid9Y7uYJ06mc7DWDjhSq+hzrpRR7Cpy++zp8JS3ju4+UXlfK
UayoCKPDcXsBlDZudjoJGIGIhNE3rqGfiXQaUFzWJJwT0Jph6NABshDzO2ZTTcb0GYFUCfrD7MDU
+gVJqDkEZE+BUzawniInBDZSngj9z/gghlBp2/S+cIAuOQ4v0nkFDmc+OrGcLqi8LvmL1Ojta6/L
PAhTInsh8ceOEx7gSPrbOXvKqArWzI0EoJDsbkWBFwaBCCROu2NKNgsD9tKPE/xDhosFRaGXI7SG
gCDsAiavbBzDIvOrJvYPGvqqgGjP7NVw3zgZ/3gNjgMGix0rS88vH6ZwA2Q841oZ9uN3bI4sd3Fj
bcnkTep+iGmYQ6RrJw+Sz0otHNhA6CItRUTEDunfrvkTrAFToMx23vrzOX+3hZXjVwAp0ZQH41UQ
qrsV8vsMrhm/f6AJ8ScYjBhXnXaqFg9VIujWgLBJY6ewLEAlEaEnb7BtjOFjk6/RvNGmDkU1iRgo
KDuM4AbEtDfBqohTks9/ppuDIRyA9mxueCvAS4zBXYI7dGsPodmMPxx5TkIdK5an4yhOCQxxu4vn
SybdXFvS7jIk4Bz45lURhDy34FPbQKl8Pt/5cdT/7/udLl9Eu6ti2ALNklfChteH/h4PYJ0g+5S+
ueiKNtkCEC+hTCqIThSpLfWkxB2PUJp6hWjJKHO2Cc2EEPFAKRHlaJMQ5n38Ep+U3sOT7+MUvqrK
/iO+saxQacFnxq2+QOEE2eydT7CGao7BJB+RxPNQqmR4GouFoliMAXymXwa7OFQOiljbY5qXtpKe
bBvvV3JLSzOq6gMaGvBslcabYyzloiYrT7bJ0mms0JAiGmBROSQTswgTmlD/n+2Udbb998gHDy06
bbXECONOkIyqY1nY/v6HTZRCSmmvIIb5vRn+lpx/PgKb30uO3jAy+fAaCx3G4Bc8ctv/xaf48BWY
EL3V/Crqy/lGIKC1kZw+UWGGww83AsO/C1/EP2y+2Xaws0P3Vx80++ojnfbiwdW4U9avGK/yi3LH
NrEyR5tSi6aI4lzvfGmwtHwKGxgNuDrqKZVh+DwQxwCp6zDoQnI7qAbIFEELahD6GCN85YsVyxFh
IUojvxRkPMYzfviVWG8ykBrjESj1f7Pi8HGLJrzAppGeF/xB58SxgRTxfZB2OkxJpUBaFVg8wzvf
R05dMQa8KAPgW5Mz9j6TyZlCcscEDyEgpYG/i5WS8pc5gyD9TD3ZMerRaFA4aguKFPQc+lUgLeCJ
iTyV7cQ/vLsersvdwhjbYuI9P15ARLlh9BdkyHiF7aPdaLjcweXuzngBW5OoqnCuoH/1Q/gSAkAB
9bIi6UAbe28N8T47phhEpzcR9gr83kB45DttTaQBRJKtTj7TDR6r1dPLu9M4+N0mEaLnxrKW/N0J
KyGtGKhLjj5CM5gEKzgn7yzH/Hpy5f++tdTSUeouFul9CGzVk+T6srQxx03cbdcJuVAXb/PJaw4s
aORio0hH7/NlG/UINrpegoKexE2pBlVjpT+798xJl3aEEzZlhgr/zqR3iebgapOAjdEGFtSTMm9R
Xpu/Di2iZDqS1E8zGb4bvqzXaxz8AN438hEQSvsGMhKILHn5FqQDkdf0SIi3nnACEcXxlIcup4+H
fChda/BKOlMDFCBPqiiIlH8IpVcUEUB3zhMkQ/zby0v1LcO8PRBUXpmSzj3m3O6P5CwYV8Utc2XW
dRvaTRNJif2SGi8cnPltn576FIejtOj8heZuGh7kEEjVW63nzIHQYjb7e0XvaIpatu2GAX5YdeZf
jyfiqaZ53rW9yfiUgurOkeYXF3mHzPoZx5nP3CD6vG43pYGtmkUT6gcCy9pmiuBsUZl2/p3tutgi
L5qJCs8/hqNI1f6UO48AEE7aluMLfSvDuB8r39Uf0ruic06P9JMhEP8Hu+wzPnyISg74SwyTc/BT
mnUmjh9ILhqZwkgbGrwfttq1/me7MFBXrrIuKDWAyvAnJJqTz01aiTczH8so+FitpRr2WFDjDAuP
us5pW7eDCED43UzKAg8jbUDGkK9DNLyokSPwt4zD2toGbIHPJXV8tUrcj+oVaNxEKmv/LQG7UaLv
jRB9lFv3GGcaoapXNphJHG+38L9aygSTGIbEfXYQRNY7LtdSulJ4IOWLXj+eNsKIg+5KI64w5LLP
1gGfxaTVKjk+yuAXVX1hJxpLxJQ+tJGu/WrHbFF9FVNXVq23XEutUPSct9he99uNeH9wUHmAb/ma
7dNDmh/IYN9mtDSohy1Aq50Kgc9v0GDVVmV+PVY91Nt8Tq640Fkky60sqayJzhdkiP4Pek1HO1TF
yPDTe/P7dHwsmcVgCb3U+gIldOTH05PCVDaFz2l0blg1FIASktT7RqAfdKfY26sjaKcCU9oA2IKD
gCa4VamesLZo9oZ72lcdmfkyd0Hfp+trOxtrbz6X8uS8yribydarGckVdKtG4bBzZBz8J9Ji8sne
7jIxmlcczgMvm/dpGsirRdDbK8lQz9lDY+LGpRd5S8nig5yN02/xuUPpjW9J/TCkneeWTrZ26mKs
369yIiUIvMQia+zmo9/L6Dhtgjwr2yBy7cghdQ1zShPE8GoSZY+VQCt3/lqM3ybNmEMovl/TXCq6
ouAxdKyKKjvAkaSBhrih1kvkSftB4nSdc4k5exF3mezvn5uA3Ax3FP6y9u50KfbDpl4QfqRXgr+b
UwA/m/smbPztHGZRW0kDqoArlS7YwX5RMAr2mQHHXSgAFa9sP0ROMpKyRk9WDEAo7U9Ft2ce/dcX
6m/UuTKR3aGSSOeejFVFjq0QDsUpXHKTTnwMKChpKfqNdLP8aPSLNI6zHi7HYcMWmfDAH6aoaBzh
UCBHfvH7S6wiQL9yN+TD8H9vcT5enCKLuGGQEbpN3J6Ckh4T3SfwfRUdfXpIf7Orh6iG6vtKZxBB
6R8todySs3+9owM2vEplTFSe58vJ+IA244Inf0OiPwQl+Tsr5vWRtFY3mC3S0DuPjWEjVp1mOLWN
h3DC177dOjCtoc51t6hcqLtwDzbIz9mNyQ+b0aw6TH6e/ondvT4q4V3KYMvs1/UyXFJLfzJMbHF1
MDQe6vkOojpTBfs5d1871+yYK6IScF748B83A9XZIeDQOYbosCja6leUDWJjZP/X+8DQTANoE4ha
l87yOwleWRc9Iwt+JDLGjh6OTSP0BcHHLiZGNiw6EYYu+vLTFEJJ6OFCp+NOCHsnLE9zLSIfk53S
BwRLe71y94lkcMBtJiveXy+4Lk9cqUzHpOaG8S5GLKqjKlOaYZkCdSTHz554fTPtjPoDrhQ+NWav
Y0et2X/ubX4lU45AxMoqXhaJGgD2G29T7ljq9Z4ClU0G7huGMw8aTo6dAbTFOT2VRPl9VDducutE
GajAgTB+quT46bvhJ0SsWOAjebEkGQSTuGCPcoBO4W73Hzl/L9tDmD/e1iKHU3kN++9ssHFAEtou
/85ToVYmQNobAAl8HBKpro9Wqq2SaGqTYxoEiyVMJivjlJ8FbRrRh/T3dML9dnZHyIBfB/UajYGf
dJAwywu5pteM6N22doqhPBgY/4d9UHKMxYpRiulBp1LCL4iX+ea6LjvWKSboGkpKZu5kHFpdDNob
zHUVqadtdfEmFjx2VqvxEGohioBtSYLOrxdUQJMw+ej21VEu2vhuMUfSrQ9+WJD1/G/oKFLu5Sxn
zj9rKUrSUBwKMqg1lXF8hURnyowUJWx7XvusJfWkTkW1nEhxu/aO1gZIDhG31pi/um8wBa2JK+BH
8sNyQdd65I5nFHf/A8BWWOuhZpSnY6imE9Ju4tqYL0pqimptIjfnaoR753zrk2E+N4b8bVyx31wF
/0/PujQ6rj6rhOD9h58/MxDTX+Fhz6Y9iwDgIXI4p60AJb5O+7ffedo+LLszbr5bnxTQD/ttW3M+
+HG+2KXZ0AgXn9qCo0s39t8TdD3oAxMCs2Xfjhut9RnC4cguw8ErQJE5ikoCrwzGqIi6vKjwB80a
+Ta6+MXBLDC3kMA1NFnzP1Km8GCaBsV9YVPnQsPjegCXd1qz2mQHAd49IsOyMP7jaH5k4znfO4ZY
thVLF4yNzwRGkBxlcLJpfJmUVnD/x+RF/pgynHli5BgataipSbMhSL5PRnM8ndC4PRg6KmzmGDpk
y2xIwCe/yfc5e5nFaPOfSWFnUNZ6LBp2LXSXNtFKXKL6P9Mv5yjTwpBHYGG9TrTpxJvvcO2jem98
PZrox4ETXr/UaZ+k1SrnkgxxQY99SgLl9RIvsnTwVbebonw9b4Rx4XpqffzxPTqSZWyGD8YXKsKn
pxfnGZKhkYuX+M7rMumXnQPEyCHlgfQh9h+QMQSgYcIjBasIW6blx9dji7aP2DUM2HEfQCHFWFd1
0YgdfbvmrrsoBV1vBtJG9qKSbxovyVymaUT5wmRi+prUulPM4acL6d8czuzYscmst9w+qRk7NsS7
Kx5u+w3vo0zv7q7QzBOtcylR64/bIcXy8xrAPjx9eNuI52hnC8XCdOz+aiyGVFSertackrB4GGDF
nlWJashX73tB4SwtU84xJpw0X8UrvsTABZPaqcMprkOmL2nBBgFVuZKvtiZME1QBRXWIoLxHXmSx
6Dcj98B5eyHC9LyfiEaXNejHAWPWkt9JT5ZyidH8UyO8TIMXjeh+O5fBta/iRedjR4OkTsKWaT6Z
+nD4zaJJrd4lEiKyg7/Nvh0YqP7+6mOhi9U4qfYeRjRD/rRees5WYUUtIsYoJwolgJxm0nLUIp8l
OVa4q7i1jlcuFb2/qBrhEZQuv/QsiyrL13amtlnrXakOFVQDY6+TzcBiMZIeVBKw5UeznZSyduDU
lqs36dRgjbsT5Ow1YQuxkV5YtRiF3rwo9pPEMcyNbwGrFkfYw02ltxPUrS2/W8SwfmwEqGi3k3jb
yTuMsKejigpM3xL7e0csfxdtq8CPO4kjEmVQ10LS5yYxql5WVXMqwuI2OlJlf8XRGcs7KML+Lz33
Knjf/f24wYVN2K2BKnDZqfUEVJAQogpJUtkatTTxBcyH27ZssthSxTlawTt5GUDfpYvn6Y2Q1mtE
m2iacxAF6Z8ggs5ZfgZsQ7m3l95gNn440QgolBTacro/gF+6Gmj8yjWNmeDQ10L0dA9akOZ6ymie
Qzba1hlhye4ij6okvb2yIXYZGlap1RhzMvF5xWfSxqcPcADaGlzDr++TiVSqVO3SwYxruXZ4qYiZ
qU4y4CJAsc2BuIM8qj2SIDKRDkTSL+5Gfux+C/YaBU/rxWoOSVThou9Hfc5zQYa8OhMJ697TXZ9d
iJCOJOQ1hq3kAQw+XjwUmKNqX/JEmy/t9fVPn+tUjUF0T+Ekopw4Osl3FVTbPxw2FGUYwl/PV6dn
SoGlrF/L84Ryslv5jEN3JH9lnQEJZJMRMsUpBmykBMd/PgHEd7ozyVgALpF7qXMZsa/IRd6gprR4
t+pCE7aFnVug9R+e52KMc358sXiJQs4RumqXyUO+9zrzRANjRuWOkuN84LCKoqW5h7MhLJjvZXq1
wMR7SPlCvwTv74PhnAoq2bq7zRYiG3f6MjBz8U5PBDyVXYN4qd1gYmc+WgyOOBfJRsWAztN92FJJ
My6h1EhpVPIJdN45AGCmwgZMQwuYZG8bzP+E6uh++jdM3dBIlla6/CV9e9cV28CRwFETeAYiie4q
dvTVmJGyByAAyn39V0Gsaj279p6rmOobZ//GMq338lWVKutpEe8QNopVO/xgN3GWKhoiCmia1fK9
8jhAWxpUtdt9l7Z2nnC9XMHcND549zkdmMF5PLand7lHngGTB6hPZFaC94B51NM0R6ns60wgAXkS
Jqc0qvk756il3cLcq//ZM1WpHTOOkgVtogS7LyOS3uIbd+l4rH76bc6/t+1Nce10fiZrDA1tD/m2
xTm5mJETROMBXAPX4YCeTNc6m2cfR7q4ZUywITjAozJKLDiawGHjijI9amGRyo7ZFvr5TRGospEX
XrtQYPrTXUwK4F07lvrR12v3kXfkNIDBnTlWUo807JGPsRFqJZakLp1ejLAPGED/aQZsXY0hdNIN
PD6UaZHxpaLXVyXFeBZAhPRM64NXI0aGFhpvHFhb8TE/7p6U9bOxGVGxdtTEWxiZu/CzG8iqr5nl
JG76wtEyZljzEx4JaLDvET3ONH3xBn38LRaTCtky3U9eagcF2oPD2R1yWQKuz5mOX1AcLjEynXn6
Zjm+/QesvH9iBlIp+gnAxinaBzMMJmrArkRgrgIdETgtG3Kx8HEicDxjY7eXQp4wWzk7yilEeZ/G
VN8IKhwK6n7OQ31lLGZ68a9lIAnRACtFg+ECqVfEvtkhIPc084CGdxqrJVR0rw/qymD57oyx7KRB
HoNGWfM4jfKr1XSmD4C/y12JUmed7PTsYbWjXu8qw2/99125nLYJ+bCbVc80ge+DztSxTPJ1DnPs
YGwkgoDo8KM+adamkyWJC6OJINR0tkEy7IgDJfyVRB5989dH+g20sHHws3C4wyyE01iDjuC9J5wW
T59HZDSe8QCgRvpUHmEgAyWPtr0xFxbpUvEjHb+yjJl1MmOOpV5kBbLUh7ehSrbpaGw89MXBD8ri
qNu0oFK3VeyvFzKdaGBtUhLtqaId/eO4JF0LVupKELAY4YEQpVMRXhoYJIgs9hp6DfGUWTzwGuU0
F4U10FKqFUiQ9FoUC1TTQ2gsBG9ifV5EHOxOXD6VOPzyKLTIN1wUm2ME825mpXTPNXxxQGl8gQvZ
gqnfDTJpBHeMmLOFckzSl9uyPjD2ULoBIpI6sU9cA48QFhDqS6DSQSzT0zMG4HBGQZ/ottMCivj2
BP8ybH16yM5EGqih0MzMnWjZfbmzTQdUmBaJJXMf0uvQcMQoCqtmuGrVRzkbkKaYQbYdVJiGix1r
WyPupNlKbnWy3xBuUHOkO9gOFSvQVt0ijZAl/UHHWEkhtAo4GqtmK9lVlKyaW9jcG6OYjyPh73+x
BsizeuW44kY1s6YmjV+CoGKQ+s5Zl5fJunEyV4l50qnM3DtalvtaErJxiVr6gUSFSupdeqExancX
dSTUB3A3GYu0FVKBm3MzX8h6H5w1dZ+sEsEOuK4lXMtpUpU3c4r7C0ByIYfboyKaab/DlBnyPMEF
YLs7QzwFVRUOZng9WOUamyNPdFlB80pU/bpfsOaskIfrCt3Boltr5sMNzS1ehhGgw+4On7E/GDJv
AvTrXlYnuwkBPaSNpWHh5DEG/e5GHkygRgpip8e9C9cbK+fjwFQfUkDf8AjAqUrRX+dmf1urkkze
YlIn2mPJ4l5V/BAdp11VqWfpYK2WC/A9/MsOlNT/LQP4ggkQqOi5SvWl1bc3a+fHzIw+CL8frGTO
GzUeM8TSTelb+EyStj9aiYBT4/VMJmimQ/AnGPeLNhRN61tV1Gop8/OlXStzOs8aYt+TYnRnRoD6
iSk2fHKlNjnEuRLlcZuHyKiGSDmaNQ6u5/IlM0/yALPnqP9MGg3jnNixM4rI2ttav1PayQLiJ9N4
+KTnZB8q9FMTeAk/YU+0CNu7T/FjdXPHAKkflQic2hA2mwPv1pIOa24uPMr6ojhCHSruSe+KKlPc
ylF6dcKKknzBqAqwcIAnpjFaRgxKlk+VOvo46cuwqJO00MrzEX8xHd40vgxViClbV2M+IHuEEdsA
0DiILYLuPjZ7Vo57xWcA+MZ3N5e2wrHrhDGQ4ciPxJl4cMif7njmxUF11k60QqJMuvnK6TYcQk4Q
0jve/v9Ghs0WhAlFMJAfBmXn85SvADVZsNJQ00MvA5Dz1ELTNMg5BDqAAqpoTAmy6pzHXvCNBjVn
hJi9PoAPC9mpZt45nsDYmOGn3a7E5NBbN5yqABGa5uXgiLpZDPep7P3KYzEuqczqe/9KIIVlGZso
D5XuzuHfhHgDdEdSslQjmCS3T1cmhqrDVNhbq+NTJJEtws2i2AXNHHd1YLOCRgGJADcyaml37k43
ldCGWEzjrynfKR9PdZZYiu2XsiILzvUDihoSqQfQn6TdL0v+Z2hu4GpksdhqxWv3XqDBvFlACqyz
vHi7rLdzFm/PWw1n/6z0dy2sPckH5GMPfsynxhQGNQsMMUsfRLSNmnSxAPOFn4z/CkQh4Fk+yVz2
lNTL+ObMvjcGtCKggGVXF5HPDq07GDFcF1SdTr4E2GLoRDElwf1x2fmtt43N/zDv0wNR/BCLbrdB
hkboniAvbWAWMWXx9xZUz3L2DxiN2c5Ob2d1neJptYtOIAKBFHEtSOjD/HnXUQ8qv35eMLbRP9hl
K9SFiOHB8ODMHnuZtvSLFDPAXYX0ch40UA+DmtFt8SXxrPZ6VKfzk8vEbyrz54XjneAynvxbsRqR
EiziPDIpdVjpOW5PyBFj52jyBS0zJv6X1IunAzPTtSEBuIgvCuccG/d5z7I0qk9LjFvsJFU7lmoA
w3ETEjz+vY4aPgfhBvLsY3OCzbuL0UjNXyFPC/Alhlf6cSwVkwa4uYOOmvaq8cGXfCs/aJ8dBKQB
i8SYXGilSbnRRev7Kcsy2pd84BOzdZfxanojUxB8pK5m3a6oeadrhzTcsz/8DYqt7wrMJoeqplTO
fiepduS7VQMpT4wxL5xQj6igqC2Xn/BMV9n+nWf2UocYJ09nLXvLD/SB/eDcyE8w3rvLf6FpSt5H
c0a+orXh3ufc3/5Q67y9z4QRVs9yWlMna9c7CD3m0l27gju98xozMtRJkkYTH+dnNEOlXC1SfMUl
5IjtprDwnCnahy2mXKMTYqnro93ioxlGjOii4B2/o5voaQU6FIDKXo6YzX1vljT5GkXRqJ+oA2ea
NbbZNcZKK6IynFkssvHVh+/zUxrDATgaXyzcfQROsUiQoKykX1yrGLI6KKxnzusNbeYhlbzjhWQH
t8T+/9PRBWlu8KpJvKgOSFnFf5bGe8eVz8y/fyPzSIYZm6yYtZog/15XthtBCv2EI8ersQmHKzCN
wtCSBjK5rCjGOnsD/1dXkQx1w4KbFKCED12F6nJo3WdpF/k0dIbLX5mmPEPn6DRfO/EIaGA1sxhw
LwnOgjCQKQYZPYgQlkN5BvoCVL+QeqnaedXB4qpeL1gJ+TpUxOCazOm0LOPk6cpBJ+zD3RaN2x+8
KbWQ2RJpE2RFxmLKsr+5ujfiP1anLYAEEB5ynYjROu20AY9ekpUDy+ES2GbpmKXlQl3E3Es/ecvj
B8rIydIjKR1UuMw15+RogZKTNuJ7B9JvA7PFGQFMM1B1+FVxjjWheuR7ULj7SYzv0yZlD+gyIB1X
mmLqNhGi9/vQAfE55WDM7Vio32xMU6hO2MAWT4bz4WiCmZZ8DAI0vn6slRNvRCLrlNN+86pFo2UO
lHxt9S79qRTj5PNH6W16YkiG//XFGQEWPumdHOZMuTzQ8BBFYMMhSdhbr5fs3OVJOAji6jrxhJvl
remjLHtN6rBT3CClfHk8u4rcJIuEnvSP9wymLChECDdVtxoDK1Zs7ZKdJaoonSy1oK4ipcOSzJ2U
Y0EVv0I5BWM5XYCxgEAHr2w/OVD0HKwQIuBSX0R8CLpNmtGY3vrJOi2CkbdDFbE7ozxiwt9V/VXW
6RJmcQjO//Vo7Ow42OiLcq7H0okG3M/rXyD5jE+QlJEDje12sgDNuHnkhf9NmBEIQ+bn9IwyNYTH
4IaLq+DGFTgUnzYAlzGgmGubK2ZHkXQqrDqnPVgf1zFrMVJh2ox5nsmSlhGz9Vv3VNqKZspctS3v
k/lvG1pgy0Z/wlNKaHKIhkLx00Bkoy7Z6UqATFmrIAz4BzHejdXgKOvKdR0dnyiB7V5fP0ly16Gr
ZVMCXXMpL387OiwWWyiCnSnz0Qv8faWGpv7UsOpmYK33O7FAeJE1IOSjvpS54d1CRbTRMCwnVdcs
gCdXC/kWD/Ax9EybiuK57GU30AzUXfulVKOBEcgI6slbO7Fp5K0YoI+6a8q7w/g9vZllPsGf4ycb
2yBkqe54B7ntOQ8Fmd/L+06hyY9gv70oKlnxurbpy28hRQyqvxyeg06rwbfZWZNv5hG9QYXiwZsy
nyk4S08JRiMiTwREbwhUuLO5TRJwjMnPxJIyUpS6a7picBGSMxYY9o4yZxXOLp3bvqz93VrMZp0g
PBWt61cU0VDoyHhDY8/w7zWEvMr9+HeiUjlZ5eatZyLRGJ4MPlt0/SzKzYPeMQZI5yQV8bBCVtr3
iq14w4pfdBc6RG6R2NWBKwpYvfMcl5QWXssc2GWf1Mfpz0Pql92HfiC1dOxffSUUNZiMr+t0JQUy
jY4bbrN5Z80I3DOVbq/P6xNbw6fNh2N3JfNvy8/KskIyFnr7xy76saqkm1XPN/nCKxi620qrnZVN
t6LmG/2Nr2rP7sqx5AOIwR948ae4JXeBEMZZmJr0amt0858T8HIguzNxDUZOTWW7mg0xVBqGCc3H
aQx6Sj6kLA79SFgc4CtNiYJayg2j8EASwSXXE3bZ9b1tJb1cXCEeoiOrFz2esz/ZItfMfQ9PcSlS
kjSpTvDiuHuAxf6kq0JAiebFXnCGgj2aXe+y9MPHwye/FtMzo263turJy7npDU3OZOkPoJIkSU5A
RPGPMvBwzRwplifKiJjHBaQR8pVq+4rYOu6N2wX+DLVV7F8p+yRM7J0btpVwfmcxRaI8B0E1yIaL
cKmznSnXGr90NSGXDpOO0jk3o8QLbuMw8Vj5OUzKtzcTE7tOg/MS+dC+cn2NH5w1q70gGSjAgcWZ
KeA7dpPZPHJ1B2gplU91f3deq9LCwfeZ7bGjgveFxXdf1Q0DV6Yk9OZ4twS59ITQpVzQ00c6hAI6
pyfGR2vWWaVWvTKiB9uB+8WfB3BCmKTKmfGHLfUVpCqBk+KyB0Cn7+JdzXRAC0JQgWMrXCU9MU2k
cJLZx4H4qV6jcJXKNonh+F3/bR52kWH4zcdJPPVHsCmBBpiKN7K60GG55m3bZE24OdA3uDOFGvy7
rXPswMVo5prJJ9bvQeaSOfDI5dNpyr96wKJtuQoDiwR+krfyMiOky19tWaHyifCbIt9Sy2C+6jrV
SeUpe6inNEn0YPJnLrSW5l1zQjxyi6Ehfc6WdBUYGlWtwcSrvN0a3OJur1DtJ6VVGScan4HeyD7O
fNMK8HNEXi3DKxflp10bKCUuI8iC1FB23xSymaUGc+r9+rjaonnwhdsONBe/gpAFxBoACHtPrCJx
fcEIk44sIKPAkPWLp5TLzvaRHoIRdBA3nvSlfga++Xu9+8OPafzg8sHijMwVo//apy/FWqawB6P/
fPrK8FQo24mItVVsQ5UXw5eGR8o+8Myi1nXl2PjgykPs+m6FWGXpHERMJp+XoK0+lSXRumHuiT4Z
n+No/RVcH0ow4mTwwDbOHOS2sw3UtKLxSyPJyRpDyHKMMJAwgT6I7Amte2s7QFQocF+xfDFtqy1V
zvEDAjdyVvmCXbiy/erxIMuzBoMKyykYazb8fJaqEKfHP4QYGbqog5D2feozxYRMXqziZamjUEUv
OXM2URQLLc+M0scjg5xAiKw4cpLIWodGkyJQw7FDfAyUDyd1Pie77k+8UeuHusLI37eldPhhE+ej
mjQDm0KCkAJAIFDLN0sWBVx7mDfo+ztbpV6Cb8MzWCbe2DcSnL5TNzqyhk21o8JSZ6EPUEeWMJn3
9/iCU0q4fvOW3wAEFuWgWOHQ5YerWQF7WnpRcttK+3Q39o/YDQBlpwSR+tV7mpaZ/+965BIsnfTa
uBOHxbQDE2qHOrQyH/veVJTN/6pEPRqD8B+NAp9VJ8fiCxXRem3iOMmXLodvzPGEIsIqU0rIANz1
xQxMcHXUTKFfOBb0EbB0LIwidK4qqhtmbGiE1VqBLAzvJRBLuOk501Q/Cj+TsLb5AUQMmOupnWk0
H4Vzvmek8/jWzhu21+rdunDXu3JaVKh6b4QP+PD7aUPjBKjN3XQI4oA/BNuLI/rfTC4TdkYhl+bv
iNuMDKLcy3ffuK8626MVWKfBJCIB4PW1J+XeQTcQF9EC5kEd4AL2FvdtnnMMOf0tJuTEvcKSHDNZ
Crc2Ir0MR55Gbrzwacs8xYVlyeiy0EDSITI6r24P7FzzZn6oAreTz5o6q8WKCBFPUW9sys0QIIJ+
JBeYeAAATnVNQUA5JivZHZy99GqEC05PHT4UMSs4Ku8+mUn5tzDhzhHAQ6mJBo90C3QCp3UiWE0E
lBZYvVnv5yeEGzBYqh32d2cZ0YAmMBoTRJ2ZL//JiC69mrpzMYFullHGekvmeTbb8IVxjgQJs7Qq
9YKBLesq7T2TmrkjhvC8NglclSttClb3xXvnAa/yS+ik+NIbwft+TogKsq8jvW+FTOSlGVIRnzGx
UzXHXD9nELxELKKyStHtLdP5DLUrHZpxQRFwFfsVke67ZTFL5caiMpaInmgxwct4gvNnmQRv7KtM
4TbTp/aMReXu0vAxcqg/wvuwm7SrlQRRi/YIrBCfx4H+V4xdyciHXoeO3GkVpDUa7c6qTsnqgKMO
Bg1TYuQ6VcpLPD1uBCNFyeT/BxRBofClZicD/CHAajO/QmxEs9q4V34Z12bQNF6PfB9ovLEnZ600
t2ZWUaMl0As89OZpHph/fM3vFpzcyq+C4RkaP6llMo8o0qpqcLt5mjOASm2qK2UizVXF8IVdW55/
WJoXvieI+hrJaqmG2beA8GVnNmWT5evT17dTy0lep2hwJPouMzNYFmKdEI9DywG2sgzAqMUgW+bi
ezrDRXo20x9IlT4mfGyDNsnQ6tYeXIJrkTJ4084VbIYPSTnl8bef6go798ibBLhDho/WFhsnv3s6
keyJgZV/rMI6dsuaxoBX/PNA1CzIhPsxhjJBuO1BeMCluGmmw/np/4iU7fr9fjyiOzNaZS5MIomW
p9GuqVcDyNTx/FYknMZaHO+3Qj50c3PmvICVHEk3X1n6wBwapaEw/RPsB4dCNETQpzTHA01zpeiT
xNAv+3WSt7vUaCrD5Ou+vDyEMLKAue/OOXjSOWrqpKAtHXqY+z0t9OzU72xBohBLS4l11yKevJj/
qG/HN86GDljjDOCgSJCHR7YOFv3XI7OBDrW6Ve2IzEfETvlboz0IigxgtnOcO81CsPFPig8hln5W
NYuT95WyOxMtm3Mn5LPWkOpWPfjdUN5ru1mE6U8Ctk7vy3+ZeYS3XWtPGfdAtRl5ck0RAxNvG5lg
hotmTVuJLcEMDy1GetPmlhSyRzb6UNm+pVHFcrDJ4y0BVOZAwb4OKyeiWJYWlQ7VOS7h1cWylmS/
yGNkp7RsayOH7439IQrAo+bzXxf5RNVCg2stVFcpSz4T95r+7656Mofex3KTunw20i94TCfo6GLF
51T8sDtXZbz8iPbIbvT6Q2x96t7kgxl7rgl+jt0esUfbwuMLF6bZQuW/lBGZPdFMrg/Q+tbOzseX
sMK3ky3hhMHDJlBFty9/amAW5samt4A6YI0OVpcf3TzguyLTMkJR/qshgfbeetR116qkMJOhtzei
OQTbQn8nT9Oj2ayOTai7lnuh9j1E+JgPChgCqmd5AjNKE5lL5cE6L0E78HYoqaJYtdhjunWAVIas
d3gg5QV0p54Ih/asrkfGdOn29sq8qyJlMvBL/Ks2zWXv24zd/PMrOmKlrIM8rL6axUPZOrUelRD6
XmE1HVXea812ItAym9NLaxt+AMAAByH7ESGKhEd/86fLsoy/bKnzBzb5MmlNSvkkqxpX0iDvx2Gg
/6zpeI5iCf2GVhk5+f8/VOD52MBYHp2gt0gYjOJBAF55+AeO07QoraIakKxy5+hLN4Uq/2TOS+75
y0KoDVyCi/36S2mAo5qiinzXOodfl+CbRIoJvpBehXIUAA+e7Yau7tkoXE4YzbBBJ8/uX83ske/Y
DXCVG4zMqsRLmYhzba0Ina6wJNXtrnhkVjkCni2pVV/2fHqfSLYL23APjmMmLi0KCYAxlo9VVdSA
Sv5EHbS8GBpK2P6BWPd8xFOuIx3Snfhkez+9xp+qE5zlGaKkH/wbBvO3M5360+0CbFYe/sMlTxVp
WApiIBw2BAvjpgSlsm6BytGcyOpnfLqxaxfqNzoWVkg6GJf8HOvjpDsLmrAxnzTtzT1NN9TKHNRg
fLfRTH8WIgEgGAmXUcDkbJWYzVj9qukgTKq48iBhcmWY9q787tkxocbHXgY8v8itW7ZukqSmICfB
PmFz2VdoCyzjsxDo3hSiXBikNrkNiY3vyFvPQifs5dHgClehGXTyXpxDgP550anB2Uovhv6/GXSR
9eUm22PZKwfQwIzqaAB9ONAMof/J4ipiXM338mfzzud4b1rR3Ib4TBaqCnv1NG1fzcTqMiYBPG/n
ESxR+E5iKce4Jw1QGEcxAoPOVtq8PAr7dJYNL4dORa7eYI1/gw6VQ2xWTLORPpejtTt3do7XLCsw
s6EytAW0CacF3gRpREarMfD/OTV0R6hvzykLVhDoFnXB/6i21epA8mXUb+/ewHF5T93ZQIierff6
cf/M1A9Fk+i8GkRPUfcvXfwQbCXfVZ7lG9LrTBFslXtO2CINJhrF4kLLvJJ1kj2hvAzbOd4OaDYF
s94KP+igvyrBUIc+lWxVCsDKsbmnzBy5y8qChsAJB/JVHi4XBR2j89mpDekefAEvyJ38D5iPKOFZ
GE1rkg/gDDeDsWCKtKgyD0SiZqaVEkVfgcUFFIII6jv2rJH127/gqLw3WpVnmBnyq7bVv5Vd8EH9
jFcN+KIeaBmbm2drXxRT12xtU5y6Z1TQ2VVpmfmydx4Z0VI8A1qyCVeDhTj4WsBrDIZ/5PSUHxyX
XEhnd7A91gAC/MrOSlqD0PLpKyu+JJtQQ2O3bvQbBC+xnt39LFdZnPRhrNN+cOLjDKTv70PPGQRW
LsdlZ4ZxLe3SihHzwj9FHzP69NcuTxlxHcEzGtB1+JFMQow8AdUePqNPxn576UpdRe53E173hl+K
bsT4wuMla/JwMAhOdAdBCpFC/e7Gz//U2la3JC1iNafzHimdA5og92nqe1+EzUFVZzOHlhex5MZY
4QoHSglmkxCDZG8gyipYJjKcvYlzFfpAvlOxiAMR4s0+SzWIl1Yutt+OsDKaks74cFdUchQbNUU2
87lWHB5zpXsVFldk5yLFMZwniumE0o/Y8iYM3o99NTfyQ9p4mTvTVO8xo/sFRKVJKyi6YIOcJRkq
HJKF0+++bLdk4mG1PmzoG+eVN+2OYGRUtefSXkqkS5C3icn6ZiMzzSpIaCpPyLMUDD7xB55GCUnK
PWT9PkCVuTpBf8j9EeUqUP813OnEiAvCefkvWwRrsGBr030lZ/FQze/JUfY2fiF2JPed7UNJVtVG
59Nb9jOR9ef/tGvy+eIw9MR6QDATQ27Bjpkau9YubyR1iegjLDmTwuKogF+f09PPlUlrTLVSvQhP
oCHoWcU39dIQw7GFEdqbQuly7aK745Uq/2vc5961hHGpnxgItbK/hHyC1w/RyfZrebsogI8NIiN4
hIeQysiWlAw4sIVHK04EUtrX6t+eL9n101FAjgUWzFX5PEf0a2cjj1pRczIZK4VKAN6q//v6fB0z
CoWG4t838iWUm3Vla/6IIar5hZCmri2w4lNFTe4EKVJ3xY9nU933KQElL1/qYX+Ic/acAZyFgI7Y
bPAHCx8uTaB5rfGUXEt59InWNlCkcRZfHcKcac+jnZtXNVKM1n3SX/MxkDrfI4hCix2mFmEDBbpy
YH9a9l+ZDe4r23fSul24syEC+Adq7b8EhduEQ0SjK1vVdubgShWmW7wmE8Tk2VMzuT2tiq1tNx+A
1jjY6Yv0ZzwcbOPoX9PwQIaZYJJYEOcY+qWPy3eQukpTh3SRTXJK34FzgPCcKCtUUiwWUTWIqagx
70hrlp8BZE6YWg2n+0g9o/1fUKCQ03bF5wlqAxNpfMO8B1VzBMXNLzTm/IOwGRZs2lmf8jSXNQiL
dNyvN1+fha+vPulTGbB6QaAY/ggtYjWm/+/N9AY7Izk2ay0ZzHqyciEsJGDpA5Z+PiTHLqMSGi+X
+8zl2r9gcQWARGLhCBphQSM2v0smCkxSKr6yR19vCkr6t6I/1xPkHoxv8XPxc+omK5weEf/4kPxP
o06KewrwJlnTE4Ax02wE/G7ySHioJUZJzvRN+tJDEl07ohayNK1JwyZOwshOcy4MpWVTi9jicZrX
k72SZjvPAtXkBYwjYvqo8v3psVuC5rHUgZ/2Lo9PC1mnOPOCtYz+k9lKjBWKiqwC6t1OdNElXZ7A
2bTeJQslzdCJ95jP3W4cVc430Hdb1uKe164z7eSU6bmX+i/4H8SrK3La3E2YEm+a/2lLJWzISVzj
ja+n9I618He0dOW0SX8+8zopTkAXIRZPR/u4K47WzNuaEhRfOGPI1xBGWpovZRHlRvUht3fXYwei
2JSwBwqX3255MhmkXSyva/N5QScwD40DjPNT4UUQQV34oJEn+qqIahauZbVGNqWxdiXn6JcCEuz0
5Vjqyw4H4tUoLFxOVMWrKRJe/qeM53CdDS6RL+1IcpW7q+kySV7vSFkhoit2Js0p7N41mWN+vDBN
EooE2l2hVcHOLZYGSYiRI1/6FmlUBRLbkhYOkasLXWIh1aHUyuIB9EAUUcjb8QW9wDGUY3Ip/Ff4
vzxTg74VkAnpupbj4sMG39V4rX6wHNLkRm/fczQjUBbqcBK7H6L/CAEOREziGFypkqJCbaeMHT2X
8hhB7ylIx8d4J3uu0UBUO+uDwGnDcNOckrMTi4N+Xfa7KcRrBP4fZHBXhCJVWeE/K6v1OgHtUMdB
0Rd99CBlRuKFys2RNg/rkgrqbvPlEcudF/AzynBAF8kQRnGtDdF9LPWVC1/sBX5hcDOww27UG3vW
rzsWg0L8fMfgGiAvA/ozBsv3jso4mGAt1T6+5UuKdIX6kqFi1mLmJMvY+R7P5xburT7EBVNs2rRr
/nNQ/L8lMQNIWVeFhu+0wJ5NqRcH1LKwhUtQu0G2FbXjQmA1+jY+ozSwzR9Wd9Ig4cK6bPtmgwHx
OMBxe6qzHX38Qf6Klme72CBOiDzFdQ64Lwx8S8GW9fcSlKgbfuvZmhMUbLN2+0+yrQ6NEeqpSRuG
7v124Yj62HccbWxn8mYvYrMK+tCwQSk2HPuyl+DaD3TdxQ6TUcaEfi2NhUo8Pook+Q65qJpuRvpN
A0w2hqVE3wZNU/HgSZts5/kH5oQ1f4CzLnsWMzZ38z5EYkVn+yPfGPtOOr45zGEYh350vjA5VwCl
mV0Jao8lwkMpSZEzTI0oL/1wNld5U6reHbC3oL60wcmmHiY7MD2+yC15/MXTjrIJ7+ho1r4dB25t
9rsBi7HmGvqI+Xyeikbv80wYchQMydX1lqjYMnFVd7v0kiSI67wQo61aTzfmGKglkxwI2Iqwjz6S
doxmYAy+0sNP1TswPWSsiOx3SxK24heDztj5+58GjY/Iy2jMi/PtveUAXU7Z3wB6PXyiISQLMXHK
Y3QNv75wN4QSo/G4OhWP2TutWynHoIneYWLQtxtNnbRP1IJpOzHkVlZTr2UgULaAl+9e+xhSCqqU
GjHfq5LyGBu4ac/qWa7ooIxyB3+QH1FzX3lg4Zm/hFQiS/aH0s0bEkYovoS/ew61EtxmPZCcmcBx
Tn94EWWujqrBX20Uvv9PmoVp6zPVHrLBfOsnSKIkAbWabGstoHHXBBcjSDoLFjOR3MyODrHGvQxY
lWivzzuwcQNhNGOEaIITylwOGe1LW9clLG1C524ACBWgaXPMyZuUsDb9BG3pmVhoVSSJFEJwxuYr
3RAgWYKmomqDCjd+JGELl4WTy8SNfGmNo3X8ZPAQZIQT8b4VS5Vd1gmNb/U+Ei9+6t0piMzL/bP5
JIuHeaSEWlBv4NEswiFaMLbG/GqYV661k7tDBlwReeVZF68CmsQdLQdz5KGH7hVtR0a8yj8H3JU2
LVfrln785HC4c6xfq9n3v2CdbueMZ/7VRl6Q9HcpAzqRwWRcktdQP1HyMbGsq6jS0VVZ90d8okG5
GJPjjatna1YmUO2m6JJkC2duXdIM8LydaZi8AofgObJFG6DWvUBWKzzT70TtmK7FKWjXKuk4ttdh
MAfCtDQpWHiEnOkDTlbGBHloqk9pOqCbULl+OnlI71lZnW4qiKOxtXH78xlXKHqaCfa5Iotnt6nd
ccfdCxcoo1kJcPjxT6csCdrN/vD6YSZomki4nJLgHi8iJ2Cq+Vxu4YvdkIIK+J3ddV9Vq5btrF3D
iMUNiBHQoZVWUtggeu0xPUm3GELRK7W6d6Os7V1Kockl0CIqIEUS/f2M2eR/bcfTb+Nh8+ru/2rY
OHBkL9AkKxDWHzMVkwG+hHxNUs0sMaQ9Zf6dJzkZS9YcmBuVdSlwxrtmudicddZGubCOX+ztn4Hu
oo/lUYlVwujF00VGtPhd+N5dxWNyDJA4V5BA2WfHQHYWqqTXpwVesBIKpllsS+AiVUtNJtsRvp18
6rVV3/jDDfD4llNn4fQgGh1NfimtxiJFNNA3X+ykwQvN8UxG7rxNtOZzPIqvfSL4Gox/fyq4yota
vgLLoxqqPNMLCG6uAPawt/hFtmWL+uYaw1SNRpfmcUnoR5SlqKo9UMAJ/T8n5Hbm2hIi5qSPgJCb
GTRkRa1TJUkN4wTw7aP7qjHdVlW9MMNTqU4WBpTwfPS2m/w3XLSOGM6Xkmej0pUHj9Oqg+McbX44
IXhsK7P5AMgghtfNdta9Rew4dWRs1rEPWfVyz87zZHVLsD4jU37nC6dMtqtNEUJvlYodAn/wdS2A
ti8gvD9XvDZiPfGFdog6wLUoJVGkTTNKAGmVf4Pkn1SqJj7x4V7o7koLIrvfO3fltWYkNq64Dpii
foAOJLcD8lp64ZkxRmZIN2k+5wV3A3ou59FLKvxfwpOJr8zWbdqbRj0nH22uzhT2tDJ+r8+ieztL
E7KuOASF3ig3hTIer0coMvSHsiIj3UjXxJ06n94U39HlhnJmO8g5Tq8eYiq/OeB89jik7r1HAkiO
TIcbNWzUmv3E0G7cEhpUCOhL/VOpb0NSnOfaQvWeezNiSgJDedpZhBfcPCEl6G8NcQMs14n9J2zT
PZsFy4QVn/13iBS4/GXcd47Q2xvp3bKhnUnA6b1WHCrmzJ3AKtKBzvcrhVs8X2rz+lr+hw7+8xeC
MUMpl20kjZhtv2zvIjOOiE+1GYuqzJoCM/XvMcgKEeOLGohasubBOAG3zd/OMyc9KhkqPttZycCr
8IkO9x8pV5n7YVcH8sX2n5UHyriliks4bKEQJ7T4kv5Z7mi3VAjUNs5TZLl1Dy9OKdlLxe44ivcT
G3gYsnJFZdifV5AD5LI4/A1ZOHTiM6VY4pZ+bG6WM4wIZvKArXTs+JRIWH9FRZtMxkeHpoKjeLFv
zbjuQhPEPwpXnnDYlXX1OQrha5rNenifO7i8jRpHVTwMFmyASh48RmuYBI5zDz2NY1o0SkzSeLrt
noZajp392wuKCn6BjVtWYhHMMunk8WpucpQijQEE0vdpWAF7brjQhbxalitT4jKN3LTIbnvNinrA
BzFIJcnqfFZQR3W/61rc5O8Gw/JLAeL+BIXv+p+ENoB9u9VrSQ3Vl1uAr7lFjTke2fN/mukSOkWS
BnbdRnbUKCm5kkkizlGrw/uD+/rpeIpkqHL72SMZpdHsiNGE8ZKTZynsRbmQGgaQxVA7RrqNqFzU
a/COlyi7HnieF1Oq9/KADV91wFecl3HKzl7CimdwHsSqJLXolbz6kJACMQYQPN9IizCELC0UCAIX
Q+JWJwCqzn1fhWF1nVB2Vgl2+z0poS4fkN6i02sgANnf990wTdkJqo1F7l6Dyuk8SNeEymfSWxOC
QRo5dWHR0NCLbO4FzrXvAkt0vvPmDwUqP50IR7odMRXVx1cktsAjCxmbGRTXqcYmPRaOeXK24ad0
MVf4FuMANq4HpcxqNUbf5QxonRhPOBY4El3dQtokenZAel7CQ0j480v195xbSMwYq9Z01BmnslZp
AFYHmj3L21McOT79iDPajK/rrCu+af0gs2HYht8hC8oIbSxtFpCjLKbnwzd9Vt1xQRZsFCyztpIb
BaZvz73qQQx8f+oLaUYxVrafE4lxuphTPn/rR+kmW2FjEyYyqfdvOkQVcHQ1Og5ggwynhP/IeDAP
wEFjIJJWG7GAaBZLG5NOUfIj2DW5fKRYjSFQ7neX08o1z8aWGITOip40x39GriJ0g5kiugQ5YxiW
qnrWozf65LkKa3J+0FeOaNDCvf4LfFQPC7eP2OFYRlz9qIdOfU8pB5E0EGJRztGXySIpFsXItXFD
i6NA5PpqxOQI0eaECvB6hOhfg7yg0LsnXjnhzIJVY6djJukaMCqgGWKzpoOqAjywvysItcNfyrA1
1f3vST6dXlM4glqQ4gfLGLFd6zlut9qgm2PD3p1Cdt8+wp7oWgoxtHSOtxAcLdo4yHe7avgXNiZX
+kvwgGtYbk3JqwdKN7fgXuOaTabY5i8QQtjYoynpYMO5yKns4THr23tmP5v0Kc+S6DrPexmCv0pK
O2Pam6khscaXdHIkKiWuZ7xQU8PTlzzfStQYNZjxPdjwe2zeLwAygmC7+HLue35iKqH1OQq1im91
+ZBBsnkmoMEe8FGzFDsGw36VfMJxQDvDdU9RNHq0b1O9exhi4zKEPWyf5I8LOYNO83FZMEi3uI5j
9MyK99qpJnOt2XQkCv4nJGgIMx6QGc28tKkRGoGczLL2oDq1hWBww47/Wo7OPsdRLva2E5t4BCd1
vmuPx1cBNTnFlVGAPzpQXbTfvZFfSjHXFS61HsC9jaVpectRjrSu915pZE+Qu3d11UvyPswthucA
foP8Ty4t6FpbCHJ6jQiYpiTsngfNn+JoQDJnYCLKyvsKTrEfKPLyT29c0a2ihsJtDAHeusZIY398
RT56DxVNEdVZ4I/H2/yjW8iwKNqOcsvKnCfSrvNWIWFOHtW5fp4mm2xOE1J164TCS8A14Qc/nfAZ
XSujb1L9hR6rG2msCxGfjzk09N0Lkopn04M3m1UO6vF8t0e4vgmqYgshfCWXpp2s4p0rq5En/OsD
hEIcmIUKlEHyllRiDA1wCs/iv224rrxIaLBXUKaiAzASVYlL+ckJCqVjF8nXQilPLSCjS62q10bA
T67sNCkBh5Y7IRQzr/ObrRj260DpCaUfrMEI6IhEII4IDg1t/nG2YzI5gdMz0RYheVu6XlKNha+W
U4BiC+1xrwkRC/e0sDR/rXZqQSs+cLcJPvcm372t8aOyi+++clWycQ6oY6ItU56xZXEPq3mHiEbn
FnMx+NhqZsJbKH8/UelDnqios24SQ7OsnL8+lEhaukALkDMA5JkVKV/PE3Fy/gEcwuztW9LIHXuw
XLOEXtEBBr6zzDL+MK6SVypl+w69gqWzIM5IyM3G5ETN7lsW2pz+9Kdaz0TqJheyKv2QQ/Irc+Ce
K0D+HrjwseyeA8eoMpJcDujeZl7REZHkB3I2koIIYLH9LRuwk+ZQJaWHBHUbgpabFd8VW28kGdvG
eKorl3b59zQwokgxxBunwsZ9oN9lWFXGAP463W2rgDoTyLKbmQdNZI8WRjGJeROH5fTlnThCwPB4
/+29uatmQ89rixM7TNCRKGil1gj8hZACoTiTRYrGHya11H8bJtdei/yjss30CWMtfK30LdhfrvR4
YsBoNVb3IvoR25CTk62n9iDstyOO/8LzISH7xXgW/QIDdzhpiUSBEGgDI5yZ02dHJrNFFoDtmQbL
slQQl+N2KAoEAt2mFANXxdaktBpqlvQf4JrTT6axWCclb6/hDXTTFews08kKPYnWTC9o58vtP4UY
G+LnjUu8LMlFU6FAbDrhuJFlBhU3ln2N69WaaxLRgVuP0hzeQOwt2MqJSCB0QXoopaalfxet0HBt
7lOIukkDejaKkvVUyMfMGR+HUNKZk/esPgv8hNmIxsFOd1/mZ0o+5aJb9ECihSJQQ2E33F8mKTlZ
ju9D23YW8Y0jL5INUKch9DZWJTGQpURLmFtWy3PNzaKYpwuPLVvewCaBl1jya231ErNH60leHkz0
u2mWrEFI4dl56MDAUN0jCgYNDi2SxABUvE0qQSgS8Rop7TWnZm/tOCaY3eRh4B/LCGZtpjZ8Pc6t
5fqnsi3LZJFEVNqza2e2cZRnNf4tlkAUramDRxjJq9DLERVwecHDH1qCh4hdSUee2M8LbQlzFZh8
Y1h7i9AtfkFE0363etLupDIYmlnoGnhnsSBEMsrQIAH3c0VWJ1Jsnbbu5wJOvqeEzGibubtqTC2Z
VbJnNlcKXyHMXK45hHU01RHZ6n2LE/cnQ4jxRurcmJA37yK9V96eVn6Vuvfv2QUWUy88qMyzsgHD
Zn9PacB1eVog6oWjyFt9lbXNcXjUap0B1uvtCeH64EX7Tq+xkGu3TqRtYTRqRzgr6rdIcF82RfNa
L3ANU62kpckAMxCMeG2ZCW71ZCyjsPmnCXt+fySd9bAOCbpKBZPQDZL03N2HjDuAxbbqfEN+2Wzo
UJbRR777v0znr/Angn+cLqVPS9QsZhg6o061shqn+/S4Yngmh6Yp0uw1ZYnz3sASvotijzIDlgjT
rkX4lCtf9FdErmVBtYdFZy9JZGEUKKIqJVpqtMHLl3Q827ErtXS6j+Sdc4STZaJCpoJd2qGxphEM
0WRNP9i3s2wL/pXuqc2YCA4evD9dUGFPTfHyF2HoG4lq3+QEuz3265LkVTRVciHZuhniFDlH7iCb
y3LkXacRQY7eIluJ4ZvJPfA8CpvQvXxsus1vFW+Fhq4xCYIfX7AVr8fz/rerTWixfGtulKhbpBOD
5ldim53bY0grdyu+I97zetf31JJ23DKKwZhNgwTbbzPOv7xx0exT4gSxP2dEt2XZon+ornJdIIW9
oeZNSWCJP4QosfhitkmWGyzA88f1+Qp5g8mO+24VE5t06spPDxf6Npz6uUlWUwxfds7OCaSjXZIU
cf6ALkrCtE2PV43tNAIu3AF2OjZxN04bek51z6/MjCx57xxdCo8NLVVvUyt1sKIm20Kr/vPPKinu
ELZLXvYQ8HGllH2sSSSFA9tabiM0opLSn1xceXCsQXi3uko/tG0BJ2bjqqt5wqflLszvZWI5hTzA
exXlvcc+5frRlkV+15MqO4RsrFM6WE/lIieea6qBTTcxvdCphTGADlsddLNS7xosoDa3yNGcdz7Z
5Pivfd8RKylHgmMRLSA4xzAxkk6a7sdmsJ7S7NCfN9ftCFekEx5zGXaRWzOaQrgbi0tawcdpJePy
7vU1rSex7tNz5QHnCwteRJQkHdpQz/u2DRohEKLJHqZ5mJGqLqdTLmd6htUWLGieQSSdBu7ySkQU
wVLgLRCvEY+LoaS9R59ml4GXQ1PmlQuhwRmPvu4rRG/LfBe+s6q/K7uJQF1a7bFCATySBi8jefQ+
z7AdmSg3iTZLcHwGmvjydD/H3P6/cBLEBHyfXa+gVpe7I7NQToWrmvlk6EQDIvJ5ii8trbAHLbvV
l3cpzXKNAL/r8NBRXfY98hV+vCkiDtqNyo8nYkw+TBcpJmmdNvd2ZLI5SH345brY+SzwRB8YYcW+
QuSg/D7T5KNe6kPGhrnH/A5RUEg959RczvnFQSyTXCi2S6Rxjin48d1Z31JArmpT8gOXDUzSS/Fr
yrnAwNg+5n+YOD4lytRVhgBJAMk0hhZ4VMlpINscvWVNUJvlpEg+CXGRtbT7SyNK3pSqcLWBa5E+
5ZRaEoia+k8B+YRN/sgNfckumvi9rT0tCfPpn+wy7qvynOtqsMb0JRIW8tBviibZsap+c7+OntSI
DobqqJj0tSX7YaB7u2B+R63kvWQ14HDrxTl3Oz7PsVM+AhvLN2gPB+k+vrGtrcuoEV+pq/hPhsp9
Hf27eTKgoP1QpK/Rxpjpcld3Sp59BVM6pl9dRqWklCqDuEDxqYFPPz4xieD/GuLnuqkdJrQJ7TTZ
TwgtmfsAt7SUhBQrJmGP8OGtJY2LEjlyoWB4F5tPuTZnS85bmd1WKSnXqrT6Q5SsAFQ9QrOLseis
uwR9Tu82WJOv9OHIJxQTSyS3JfZ2XBpb9RY1CqiZVcwHKkF6hqS9KA4jn0qwVyUOcnYKBMjj0qb3
df4ff7m0GU0vd9uGSBas03zP0DzujwDPBVrMEizzSaPejtoBoB+gea0LcaUiGEU8fEmBDF3GrslO
QWKzI2KRVt2TSUUpSk0JsEKjNeFxl02eIQJNrP0LfZqzaPlsrZhu2g9WsONkJkYh6oJMRsJSwkqO
KvDDL3OENVKuJqoxpY2PQY6X6y1eBJCXajOGPWGmOsTl11ka0rpmFCHtShBCCvHVLHyQxOFCtzes
Kx0guXG9PFlkd/gc/fXeaWKJVw//q+7NPjScZjHo3tbQe1eHGtCKbP534sFldxgBkjgUJLWrax50
2uH3/vqYUoL4YSFFCJ7+8I6tyPfhyL2YG85lPO2VLXyAlVdz75c2ZIOJMJ78gr/MarlCbXItQ5l7
1nk62dESuR2KQWS8JRv9ckhKwXbqk4sTDxvW/UgAJx28IVmTkLx/sVEO+FLW+mz1Qd/iWukABhA5
91HyUA2wnNp6lqxwNriYk+3dc/ds9ZxnMMJ1c2mpP8c3Iovr+qTqOmlvBFfZC5EIqVb95xElsLOP
Ney2KZeIeug2ir7Mpc4mGST231UUFDMsYmAbNNoH9BuBWHtQSQGLYbhgYAApcHXMSbZH4lz2jeul
ZxoVmbAd1eVY1JTCzICPP5OJbUDpBwYIUT2sevC2T+pFdbcIfS80bIztXhwK6RJlJucl/miDc6Yj
o5ElOI/WhOEGNGZtCSxa21ghBrBkjEg/PDogT5m61Kd67tlm9LUdWQ7Hf751Aecg+4W/9XeJMrco
jYCadQPMK/cPhiP1deTME086m7eTXKx7GOyp5TcIVoPxFUH7QDCMMyRbyv1EF4BqlxiNuIAImq0i
GVDLLdAC4p1mmFuYfLGdMIDD//vV5O3lViHf5Y8xW5CC6JUZTo7ygpoZqCceYPzoThga9ZLXU462
cRpvXx7MYYQOqlrq9vTG9+mty6yt88IJPxDNLpfbVu34QALd0hy8LIUvTEr19XLzrYsjIKBWL+Fz
kx/6Mf+UsHUG3cOnV1f3TqtuL8MXGsiwsX+uVNb8/8fymNYI09fbQJab0qughUDrtYvWCsVM5Qzn
vvKWJ4kTuTv+13DAdl5jCRRTXrfl/TMydjCb3f5c+eUXceA51QORcu/BxpqpOw/1fOEYys/F+vdm
Uq7PAtHseLntSG8DlA/RZ/CJrMJlkoA1ccLd5KoluWG/n0TfGT0NZqhkbw/89vrGnwIssm49ZjtR
pJ6/oJmGbJWflbjhmJ1ZjBaHFay6QYRjjFIHHr1kEk2P6Mpp6YQUYPcUZ8zXBSkOGKEQ2ZV0nm+E
TiWogiwzU1zhbkp3/shVSe66DAhDxtUps1LH/LEtr/4383P5HyTBzQo2AS+/imwa757iy45mfux0
baGei3xEfcG+eqiqfU3rdIdDMLwsXUb+5QRzWJpYaQ93YPxI77AhOiI7EXvIokDi1zx12C/ymLyu
q4D7XshSWOT+c5MsC0b7fzisjoM1Evj3UTJowryNpXNctUjw7z3PC9wlb1FcluIrvqt5rcfQ3urz
5eC6Y3LCQUDuiKpkH/OPTPg75aFhx8CG1UErylrB4zRYtNX+W2s2guWS/eug89lQuEZdhSyQGaz7
+tcHKG7iw1gvWfFnJ8y9yGxRC2386FmaEXaCKu7sWt8JsGA+G63ethUviWojhaIMImyfaj5A2m1q
/yoFBayxhxo2ecAQ4QEEWrobYpJI2nFXaJB95OYU/Mmrbfq6RhhdibeU1wv+83FdFadMoUMbIVuj
lVeeoascY1BbhiHURNXGF/4Tw7saRRd9OsYFkjOhfB7hbb1IgZV+h4I4O/IzPKnhx3R9jKQKIru+
g6ZHi74apMRdPk6e/LSucJjhzewMTko3lIQ5XjTs/E5HMkniF7rxL849zkIzIC6kyeUjh4sR5Xc4
DmzHjkDJ41QO3P5KGOA8SFMHwk2ZPS/SBDO60x4Sd2Kv3pUqXia2RHn6Hy+AXlfazk+pWQAVj2p8
fTFCjblV/lfd4qVi+wMgLj+sN1XwKVy/ruwhZmnByZeTGrjTwGgcd62qOOm7xUYXD1DjPrIRF6bJ
L93CztZNMvi09W6it8y5IidSR+wQYVNxs8/sx31F/YnbQJXRKuzd13vFp2soPRTM8eOsrqfqufzx
Xbs6uaR2voyJYtrMOIHDfbX1omI49LJYCaUAKqw2AI8J0+tr7xSNPYtQiJNtGxNB3wxeL0cAsJFz
4Q2tGW+dy+DqT3uCmxpXpJOqqUPNkqa81cFntstUC1IwZh77aTfI/2KiDjM25mIMAJDAa2++bQrl
5WD3LkvoOd9sgnr6WaS3NOVXeZv07BQOlb19qtekaYo0BbZUesF7y55PzpdJefREYKRERxz4fBot
cjxVju1xntIMjKUknEtmFtsJx50OVygVD7UBl+mU4XPo5vTHWYG2lKshKp+XLJcCAThddeLR5eH8
7irGxc5xYbAdmJpVuyp2tnUjJpHxRU+yVp4KCk36H7sqiqO394FULWjaSyaJdWUDZiE884KEGYld
kbfupcpbdnoDarRHMUgNQkeR9/IhZjDCW7kNUry7gvT82aoCh5TJPxetq4Ct+3umU9CvCQ+mPt0t
2o8Jm8nBbsPbBd7Vjb6omcawYdIGFyRG+8GqY87vQN52roewoxUbTP9cjKpnfYG6VpIfvJPFNMkj
iNEozMO1Tf49VHJbvpY604IDY2kjD35HVfwroR/yNFsGCCIXMN2UJwIl/tgN1VExi8d9/NlgrJvs
Y1afsqcZ7HMUuLZ1n8rHhgG8AvwjWDFtqsPcwTTNpntdz0ACL7NVkEJQbtWgds7T3AStMusKdCIs
nNWe8KLGZMj3BwNWZ7n3ZzZHacOraAQs/cpSEBpY/KCXR0v3XB3EZFZ150FgRfilT4bBC+xUleuP
nIyWZxpjM1zAwyD4+YLYBWwc4RpiT0vS0mFY1gr1sb5hxfvskfv9IyENMRpdia0sHGi5fQKohvGB
1RcdSNuuWrXDS6yhJ6aILCVRCGUBXgmXFmnxFO9vD5CM9lina0swUfj3NMXPXqv367AP1tf35tbA
VgLZM2kbSn9IXapPcuVIyFt5WzdK62OKOGVizFdhe90qmOTIsUNw3DJYGmRupQrm5dvS0JE4H7do
0cBGdxMfEzFWGZlXtzOyOn3IB0N3Bq+2P8/IQ0SXZvja+JBSoPgNKZHhfTNVGZtmIi/N3wDW+7bg
y9aCUiW7wR1TX6g0L5yBdUQPLuRqS6ikoh0WeIA6TMvZ3eMFBqRB2Ii/bWjErwdkSTQzFMaXLbJ7
uiTidACAMqhkN93VoLjCsGuhA+XBVVo6FByyjDWlZEAAC3FrHA+JS/HTY/i0Tv7H5PJJOkhwYD33
QOeKdun6Vr0M82fbc+mInAWJAiKG7GD4JduTpAY/VGTg3aSyI1p+65CDQ2b+gXLfb8vokBYMrXll
o60ifPAZ0bUm+ZjCB6vRIDTHLKpzAfNlyYSrzgjE72zxGDV9NaOnwyqUZ3SKTRcY0x4hhe2iMeBb
B1wqDEbQQx9ap1Pqo0az8xAxPmSx2pLdBoG1qGGuWJ6UC0+z+W1nsHTJ9piNfG5SiELUdKON2LXw
zSNz7oyXIT3BRV2sl5jrns/kum0rjdRiTsYXM0qjasV9UICvq3g557ZWrf2z6xZ6Ydra455GT8Tc
3H3GmZswOyZtHvouXp9/HcH86YuR+U0fWE3860OwPoBc88qi4lQEJYfH5WpILjjlNBkp87bn2YBo
DJYgbR3KGopgiuQ4GyaNLtcQCwVkdvjjND+LLN6gueCqFfWKSP9z0hf+Vff8/cmrKc2BUE5ejKgG
aRM8V7zJDGCcX+psuWd85GZV+ZA1EwYqciPJp5sCLUGmW4E9GwQWX27naD0nQ6P16TFFxUll6inF
BZOA76v0L5PyMzQOqfCzt1Add4fy7TYxrcZg/gD5gDfMP63/Pn1Lgw75FRR3FufhNe1yZbANvmuR
QM5+DsJK92r56vOz0sjHgKFufQgZrjDsdAlpoiVjWImeYaWI55eoWH7XpK2dpsEZm+9NhKL4OA9n
WNEevedNHMt2GKK6W0GkhXmspNno9EivMMX5clivHsf4C7b2fep8XmX08K5QIXHcTzlybe3gH+98
Snuk0oNTUwyGz6zbcT8C2azNlIH393wWH8hxQYrfDDH4fKgjuOJ87Us5eSmr6vfUdL6FskUYskzG
1262mtWUQFTijGN78YnU4JASnJUO++8tcTOyN5N39wwWRK6irRulkgsNRVp/PeDCZB810vxLHz/f
ZoqAyZogVNZhI8VGDPqaCrt+VkoLATxR+8Z1DUl4Mu3J7nVA1v3N0hnilV23yFURtSc0srT309yU
2aMRG3LiGuDtxx+dKSQGezVJjA3Fx26l45Y59xeyozXkK61vbpyQvjymWUQ0kE0ZeShv+ynZwXhX
iQaESlj3OLbAJblhHw6capytCiM6Z02+W3siD+Z4cjomb9UtVztz0+4lalTmN1rcAgW7gyx5FArJ
1apAwd+LHlRlgmyYE68HwadhD/HI6VtidXGgijbSVgnShdZKKQOwf/Tby4PeaLtxJ2f7loKFFjA7
0OfQgx7oJ4ov2O+CrNjf9osN5XxDRO+UuVhrp/PutwdHNxeFr8kIZ4FeFB/Rmo14UPobcRGjZZ8C
znW4Ylq4Kc/WR5pPEP61AIbPp3DlagwKi+yOyyPb4BFcrSmki8o2ZHw7qGqqFdxWHIwUAIyk6CWT
WusGIeLG582JhR57iUBF19dpSrO/wptRpXjFh0HZvNt/E7RJJxF0G5WMaIHXUo+NXVKsRjLlQIDa
mWyX8fTvJ3sNJZjsTrtCnjjF7JqgxXVssefWUwGYJCEZgIoNIpNLzrNGVjaPezpSbdctHcEVL+bE
GOXGfb8GLgcqvPhxq9fekF+GdQ/C2EemmchTwQo/N8mlTx0FCi8Cy0sDDT2eUfZMHWGOVjNoMlIe
bdhycg5mfnbD6bf46wKQzwSBSO0CekwkHv+ntPBPOw+etPaoH312dv13JKgGMOm32VFqsNH1qlAc
Yw4GwsupKum1J5uB1+l4CUoF+8QnLDhGswXj1ihGZl4wWB9iR48BqhBxrr/KGfO98nxgunpuajBb
eQIkT3f+lauL5kg1lkeQhHU0RVkNHJ/Wbv/KYS3pL23apsWnb7i3kAlJzahT+iGa6RFjJiHbFW5p
XOPv9mt9laYkOw+HY5D2qdGePZsQXHgkyTBx3cxrw/8Zsx9ks5r96h8PdtSCM1jW9XHApsPkMgIn
EMBQgAIFpTKL4WVyC1W79Q7F+Beh2SmwdqjEGtwFi1JYMxQCCxUM/YUzEGJw9B3XDxSu5EgJt4Jz
NYvRpNtoXXoO1cRFZ+AiWJnKA2xh25dFwwnAQMviwkp+CQxyUEgxkCBQyu7bt97fN/jKjMM/as+S
awkCjsZvt99lZxyD48fXysXxIZaeQmHSP+h1pfFi1OWsL+tZunADnI88gyMhHqkcQ85vHuoCYP68
HDGnNqmEf50CEGuwPytw50xUx3NZKQFNRNmlfPY34KphWaHQb9lNEgPVlOF9iWqry6JXTqcKMvoj
gPLI5+KP2YRkHs9iz0eSciw6SjvjUasPUiHWn2FWPDISXAp1CW+5GdOb4c2WZn39jPJuwwEOmN4c
BnatNNH2mBPrxM4IlZWoC1o00RhoSSuWmQZ1cwU3eU9r+jKXRsNrTivrPp3IbpzgTQrzzeHVnZx0
3j7hm/Ksfc12YQciO6bO7dUHK9KyegOgAg9D033iWBX6yeOyi5Ky1wyJNMmczU7w71GXGD8pVs8D
mG9yq5v6hTenGvWMFMcqlCsMMdbbG8ZuZIvZekiS78420EH5KyJnBShVqsiTYI/iy02iFk/uhWlg
tIvb9xiWcc2Z10i8Y07lic46HR3qd4wIVR2BhcdguLwP9RE+ZQyr9A7SeQ7hJQFwVn9WMRXffk4c
i4jrGr5Bb+aG+VH5ySdjC7rYIQzzSq9n2wlLbNn4InRH42F1/oLnhcdaHtJsAD3haIy7EmGD1G8W
ySfmZnEIUQE9VIMY7+rsdXlzRmjAtj5scR2aV6+yNukJbCQfP4p08eBSV6aSDhcfHKoHvzlJm2xh
YW42E6YpPLrxWZsCqpR5VyucavRITUGqBoxY6fjO8zoMD2cWgmiKBOoRWZgjKks6Z0UY8pcCLeTt
SuMpSE3ZfCXa4d9M9ibUpWjJa7f6Rr+opoNT0UojS2jijL6DeYFJyFaUoVwl7DSes8DjkDeG3HoJ
qPs910uzqZcVqfBuFxLRA8u0xnwX3imGQXkNMMCA6tMXzjncYhfPNeOMlDFCInSBDDHlIzFBMvLX
p0h1NAFdG3dcGuWXpwgoy0ROlecsrebAOA423BY2OUmJcy7+W5sBAi/Kbcl+Fedb6BfEddTvhFwe
IFWSJJk1bc7ksrVWM60gxTKffW1cjIn9UwtZb30u7abcWorODKF6Fkx9KTDaNrgdVkR/QvyfJJ+i
R8T0TWEgmuYrAg20qANAOqV1NSrJFOCgdBHbYR2mxCFSqgj2ofB5EFfpGtFhTfhD05lGSfjRIl4T
G8q3+H72WFxX6GkzwBgWEt2SRfjAuQ6dHRdZPoWH904bbwUSTWrAYAo3EbCQhv4OlrPG1z/5rRZl
eJ7+AzZZuwA9h485uGKZoWWcyH2vh3rLwPMy3lmW1oAC1LxZ+PaLft2zxJz3LUuH4vGpFEXuNcgX
t4y3lGUvU8sc+FuDJQZffEQJzu6oSZf73IDRmWVIz2PHGKu33+dv2NNBJBnjB4I2NQzL9H49EYAz
beotiLLgNDyb83T4ac6fkswRHK6tpYa566TE9WPFwz6uLkkuH9ZWInNENSwY7ndh70eAMq5zdJSP
sMdWgiiG1SY27scOBEnJaZ/cK87FkRY8x6PmBHpKN6gjCntFOxEgAkqnMOQp7OMLv7nobjjSCik0
qEac/Ghrm3R1afmygty5XWHYFDY76X6H9vQOutvP2kqYUW9nBCCPnaNDBLcT5DdAS15S2fWKgRK7
nE8hl9dDoHCQrKMEwaV3NzOYKZpW+x4a30O3vrwKRTnJfIkn76ENkShYfFt8V92m90mwplX2wbxo
6HKLtPoaloplQq87/HMLCZ+jrUV7uwr6HaWtvnAoU2PybkIIaD48RLq5Wb7BBplRd8iiZdnHj8SL
pNnFfkjU0AUv44IMPP0AXvQQXSa2li2WS3zCNsAFUMQLHfBmx1b4yiPKMZykMa9xjDKOslOHOWhw
w6iB2FI49Vn1SfbHK7vgjX50VH6bQ2JfmqRT/Wg/squlbY/5M32nhuoNR23yO0ynH394hsc+jiu4
RhBKKoY/M/5SoHnaBzZgq6JIVPuqBcTqepi+5+qneXx8X5yXqfriArZmyNyERqDdzWgEyZFhvRuR
/swhvKmudgad1iJTZ0fpYeP88uvy8bAM1TJhsTWVe++lYc6t1vjtJRZ7X/IzWcxs2Q6ErdVpGVFh
hoiSiSP/t8aymLEs7mf0cyWgTpDcWk6GmFKjHcLlJZyz1qAmzqAx8Px8IHBPbmdy40qIl2rDEj+E
Svpe0mQ2OKaiCBe2LbYDG65U4p3vu7Z1pWelAIy+2iuxBMrSBqoXOIyby4KzAdPEPBdAfmzUUc0u
QPt4vj9l6G9hxR5ADKO6/IMxcbiYWBs/Xecj4G5e4xfWb5vGMD37wuP11i+dr1/bMdmkpzXwsJci
/An040HevTeqDg+wdAs8/RILIrl/EyNXxXIpC7l1tSdLVDuFkfEiw95zjtEQVGUTIC6OYO0wozX5
ZX6FEH1+KhTArgbNMp6NujJ410yR0sf+OrX75uVKGp/S1PaJRWeSwbQ3ckBWvvdl3bJ5osrxcZDg
O/54Frv9W10ore55dKCEbaF4qeqjcI29PHKBpS/8QnvvoZ+5gndgTtf9d5dnr0CLdAdyVcmcAKlZ
rQ59dJZQY+5XXbmLo0ph/kVBq58HiXUXtByx/PRDhZCoQdAJ72V0igEsVV53Kl+/VvN09C7sbOZ9
re3TB1ssBENamZXHtjW7EQmoFF59OOepUjTX9sYG7HT59GRzhcc1PquxNchzD1He1J/AGpgL9tyw
7fdsT7SjKao5odxb05kc7ta5DRAuLF3P3HLstFAoWD42by7prbY+wg9GkatqoTe9NfoiE3O0fskJ
T7FeWSLfnaD2VnkD+na4z2U52yWskfjgYb8FiuHw1IOKVzmIfiuwTlVnegXX/3YR5jwE/Q/lF+4z
tUwdZloVxcvX2FMF5rKyeT0OEo8lgV0YHI1xuxepeIyL1psCkhRoWSlCz8nA9ypoWwnPNnn0+xiQ
i7AQwlCgpb7jTqhFgEbekOul2F0XhHLbvGiWhVXeTvXMkc+sH2SX9DABpxe1kCcj2tB+tSgskkBB
vvL7AiwAABZCIAPu8WDcLeW1DzEWt58WTczHl56kVzgaUXO5PmQSJUrdBx2OuHdnHnMsqsOvm/yI
1zkEO9gVp+WbocTb2yLkWTOJ093YSMgqifD50USL9hHw4w4+vlrLSDNrSUavnECsJUEwGr8RQIcZ
Xh317zK+zEu1PfiJcn5p3Q04kj5k0rPQFuTYNr3uUJ2zCyVo5vZTVUf9wFwKN4kqIqQGjv+N+/aP
LIF1PsD84TiLRYh+R5w1AeVwHV4I180RA0sTWUfK4GR4h61vqbS4EK95WC0Vh/GzptI32aW31tb3
tI++LhJlzPy9HufHskoyYUaDP+AjkcDLu4ujMuwKrqWtKLBMkzYntccWuEp4TyVKIQGkOdjilkun
6an/QmxxGGvv7V/VY0FhMujWERohvgr5AjGCN9QwuGo6jlhawIej7AtmO+s3gbELhqmCDFfECbqG
EqbPrPxklLQjWmvmc2JYBQCK7MDJHlsSKEU0ftxIk0BD3Y/Mn8XKu+T+qedSfddVbfl7T0Q1L/yo
RUCdfuY/AJz6Zqb7gtJM9H7Snw2c9Plzee4ARuGrBSwQiAzQHA/XI2N9BIhOVu3ER8Ra7HSvXPig
5/vN2KTM86FmuTeY//fNETX9W3gAflh4rK4mBYxFwyI5nH71BElwmaFOza2Pl+DUJUVLig++3lVl
4Fo6Ugya/qzIzHg22m30gTYXAKhGfPg1VIPMPfAIgR6NZ47S1Hc5UVicX7214eo1UTPW4Y3Wmwhd
tsvvChK2KV7hLeFmsQg7Kt7Y5OGYK+XhbGtKpiUXF38a38Xb5MP7d6XqU6ivWCEj2DxTY9lK2W6K
sd5JJlG1EbbvRhO5zd5hl6aQurIQJQnLnxlD8OozDvYzbltnpN6/B3G3uUPhWOw6lGJPHaElTG/H
cE4wqztnxgA5eyi1AOX0urTnqTkwL/LgWtGuCfL+RQ7WvneZzNOs5xUfJCPHTDnKnSuTvOPFB/qk
uDEyxlRIvyMY5G1GjBoxaCfVRsovhCN6c7ZuJGUiVWRos8vnAdqG2zlbLAjcIbt1tkBkP965eKIk
Js5p9aRThh1so63jG9a/LsiDec0xT7bpvksXMaDltZgGErfGDnSpQR9Xg0o2wvvBm1653wZtd+2e
ZvE+sGTLVxrk0bWbQqiw5RRUTZQw7A5op9G2J2Hk++drFdWWpHhlgsHCzazUMr2IvRa8iIXhHfjd
eeCBOrywSJ6XsR2bXDccH/l0KbsmKArCrM43fTYbjfuwdFgCmdtVffkI/aKgP3ASFwZtEqsThTnL
9T4JC2Asf+EqZuee5r1UNCHS6EshAW0Vda+Gx3A1E0AVjA+fX8rERYBvBgHdYxKySIWlchwloHmA
vncE4teKCKfj5TT8bo7Cv0unzTCnLGXY/0HQjxrWzQVg6KC6m/L8IJH1h8zxU/daju8KVa7lwRpT
Qvg3EwuMs7qs/5u4bv55ZHAMI6ofDd7POUVgtV1F403qC7ohE+MH1serCDieHdGXPc5Xex2IiLUd
F0XU2ucNX7ebRilz98IzVDeiAD+bn1UWRZy48DepbmF61vcoT/+F7bKnxMQa2iaLoJT2Q6xv3+qq
n3QliZgvE4oGBgiR4Vu+6nYVizScEQWVFfmY6PH47ort7r9GE41yYgatJFi/Z4WWa1EGUknABUlZ
RK0EsmghDmX1uufEuvsqbCqBs25mkJF+zHV6J7YXjBP8tjQ82hlmvm6j+BPcfm1B47eu/AyIIL6S
TYpoCRr/A+a+eIGrrRnGcejON36Z5usTtYoVMx5y65yPOXeYnG4rW0wP6JIvPO7LuyEc9+CplW5y
Dhe5VcZYQwZTg+R7XzTGtQt4zHPEbgVURbWCaf+1vvWRisEg8YpgvBUEBUxxmvdG0FjxOwOVMym+
ZengMfSgKZ3SHr9sqgSvClIBuR/J94e6tx84tD6+RjISzBynqTf36oko+pGz0r/9563rUoQqg2Hj
aFSbtILnp98Jy10JaA6kryqX5kI3BB/KNz8IhVe2/qbde4mNlq4ueoAX2UPr8D8UFu9rfpDF/oVp
QMi8DGj+M1bYIS4Hv4fRfUD8RwGEbs1LIpcKVeXRjg3fI6joYzr3UAefGwUzipmk6VAVvUCPKD+j
Cj2UP6gxeGxSEQToq+KYlpJAShdga9jpmZlBg5aw0mPI+FdyFNdfplgiiBNGRPWLMnjOrgmqeWqo
21WN3kwp/3CtdadCIKXH2pPhM1Ji0Qvazc0ce0qZqu6wYfKIEB7tU/EZGd3kaY0n2FFV01Uihfvo
QBj/fVtqnLPsa9MkHQjL2U3FVUZCuqw2//InBPPpEk7GvHqNrssnzdMdAcdAtUBPWcQWnYfjCqgd
Rm0q5sebkvBiYegmG+knLtTbQUCH1TmO8G2M5alDLzp4B34QANmpSNXh7vIc3rktG96Y9efbVomj
rmiO+n8Ee33kNqmYmMP6zdeBS64A+HcEj4zCSC57T31HTNCdENnjGvq5TJyrfGEctq1CYYZpoUVC
Q5D0KT01jKFxROj8qmaSKGq2z15i3FHAAoP5T5/vDpfZNORFBiEy+SGUSuzNbhZqtmgQ7LDZ6ph6
hQp22432tfwBI94XcmEHEIlCiZ+Hifpo8JiSucB3CvzpdnyJT0elHhfHSj6G0P6WmGOqDQNKxdFz
OVPPtOn/D5GVLIKgBh7lUhKrzqn63ZGOaCY+nwgh8TdrVw+jR5ERGoJNKhEb/8obNJ8+zxEgLUMX
zDhOegh4vK0DndWgfx0OLFhcuUnpOto6Geng+X3RA+qNxmh4dWgKh6IVc4LFEFj9bp4w1wPqyhC8
bP+VxTM4UKtXRItFqiN3S1zZAsAbN4Bbgh8G4q2iZ5E5Ca1OEIAdRy3DbNoMFarGqzDXGL1HcIHC
BMiAk0mPtMNa1MvS7Bo5B3VdM/+7AiJsp9A9/KW2RNcibXMee4VKdQU8aopqvX9E4XGSM4lrRF6x
gQTrHqWinf12RPjcYWAcXDweHvtpTTGEnGpbhdHDYYBmHDFwOI+QhMeF4j/de6QtLdl1hRWy+9Cg
RuH8HY7dB2WquM9YVkhQOE2WnTT8Sfv6x2rmA7yygL7DVNKknh5GLyUchXvCCKxmbLR4mp6J0Ho1
B4Z109tFKuyimDuHFSKss7o0hXL4EDnMItAuyansT6KIoBqLpCcsB7ECxUm1QtiZ0dheaq0YrBBK
ok8T59QCiX8YLq+0NW1aHqrNZpqUQnUhtIp7MeCPboqnrkO8KTmW5sYEkVPAskb98rn5JVt03oPd
PNXpHPQtUEkQnIOztZ1GWGZeDBioXYhh4DDFZhnLfhjPioLmonYMC9oCGMN6E4DDhMKLSgI9i7Fy
RaZie0FmIGAVa6VTUQYrQ+YNIKIr+LWhvMhnaIS+O7vNqxEIIZe1rSVGgzPGFmMENugOmD0ITKME
k0qXGRz1wbvIc1RTDSic6BBqEyJImsryeDe46gnRalVMt0G/Y/HNAY6FZ0RkmA8mYJMtYUJKfFxV
1EX2oN2ZKJrQ3gqNwfCKiHFdJZGMKbpylQjdyVNL5D+mmjPHU1lAbBkKW8jN5anOKzCkuEIvfFom
Z0uBEhBYe5pwqBZYCTP0iKKco5FhCwRcbt1H31z7qnwbYwiaH17FI5aNbuelvS0AZBbDwNkUv4Wh
jVPJCSz/eKLAiO2gmV3xfIVcDkXfYqPBFUeo7MZmPDJFAzISw9T3owI9GpwIhUSQpkKVbDJq0xvg
AxndMiuSeVjdkR79Qy8q7onWTHnQO8uFH+q+jtvU4UPKBUp0uX5k3N6zCK85tuao/Uv/G4qIb8tq
UluBQrslRG9avWLzSi4AO9vRfixFtHmEdyVFsgNIP1pz5Dy+1H5slzVThWdwzK2sDP/NsZzuBiiL
cSW5h/odgKtKJtNgJt/9Sc/NMb4mAR7CFbBTgZkNoAGMwqmmDTEIrDikZu20AY2jAUEPCW8T8Z9W
3uJsMznrNI35LTY1o34i1pq/W3+4BR17y1oZYEnMyQsk7o+2RSoJq3ZHH1NAkApW2lR9j+DWQgAp
orC+2Q3mlIsBEompYpljZnRX+T/i+yPi3+t4fcvOjYpjfiHjJjqjZe6O6gIgXJsJlf1Gi8vaZL/2
SUh19Ybg4VqsrlfL+El5X3j8vdHDfBA1UqIvsf5OVyqb5unsoZQdK34gZmXt2BjkiGZRmFzWQPKe
biGjgZ037R8dDLhFStCaWvqCMYmBAzjysrjqQCg79ixsB2f1Wt9PRILBOELS7Y46CM2KZgOSY3PB
iNG4yQrhZCSOPXPe7LFXDGXx0m6Wvox3xKWJZPYQYa+TDKseNzroHPNT+sqD8EjYGkk1BdHLP3iI
feSonW5OEs8UTqNNfTOOvpy5aAzSRv4IYWjEivlgyydzeget0XtdTIo3BhvCBd7FrlaQrK8aO2iY
92SHmiSCpO5MFydHvJLLtV0kQo0JrVw4CDKCN/m2XguNgGWv9EbWJhIs9d7gmVzsLy75YO0Z7Oku
NdY/osiWE4Vv8LICSpEQyDGFH2HqHxAcRBepx4XWXXcuFYA1oUkkfZ0FU09Mla+o11smCH7It+d5
N7ZI7CGgLWCCd5+3KTMzUPAGFxHc01uhOWxi9Xcb+M8X5xDzPyG74MEnyrZ5VBgS5f30FbRq5IKc
/9ps5V9ulHqEgS8iCTLxOJlqtrkHjx+XG5aY7NLeIxoWFfs00PfFFMzapi8veTBvU0vDzZkN4a8b
3LBTnQNNdf29YtlV6tqcX33GGSPP3Jm7/Ci7Rwpf50tj1HphCRRaWK5zKE8LPBccl/uOKZnWN0Go
RLLZIy5wP+oUtEHWl5mb6ywnlUulHQ1K+87oe/VKDgJla8JfNHh+9pKB8aUFwxXWVg6lvI9yHjcG
wybNomCFr37xa1AmGgeeBSsmnKe7Hbz+QXZ22S73RwdyGpqi4b70ldMKponWDknkjUBwz+2SVSq2
I07ii2m1kdDlOpltATR8kSQD7qDVxH9WHzU6cRUKEOrVHlptJjQiJBQzn+HuLbQIGPEdX2LfaH5A
GhALe7ES+MpsVd3dKRa3N2eToCvHU2T3NGSh0d96koLASeNFizViv8y2/AD53PSwxZnzLF3xzBwv
T7Z9auZFhieiIHZUx6OddK9MyptMgWvQNLqp3mIZrAWaMyMZSIlX87sdUiYR5afKwBX6tqBDRpvJ
HyffaerbRw6mZ6rbHwVzziSXrjCffl+Oa0KEaSP6Czt0WrdjH/LZR+2gkrg4hEKWuz5xFl/PD1Gf
40OqUtQ4lKjbINrLpqXWT/spd2UFtwcPy7jksL3ccgIUu3UngDffv1MrbpS4k4VlPIEeQgUa1Rey
kPuL/15viwkGv72V2fEfxjG5CNGsbM4Y2uqE8UmsMrQRM2xfoKQoGBzHD/FafQ667qqCjMpnHxfJ
3xPVQX4UlJYosD7BtssQV2BYn6ZeYcIRQ8U/OB1VKWomCm8zimAwMKhMDTGcAI5dVoujS6sK/2s8
R8CBCyadTQLKj24XYT/WrBGt7xAhfUAITGC5+CnN2iCeHxlITWRJ8qKZMKGIFzzbNu1lWTrLWcWf
zHm8cP8teGbo9lDxX9n7s0uq8YP+kB5VpdCUnedhcWBrIzeQ0w1A6injf2BmqSJC4ggNZvuxLXA5
fCJz5GZuICioaHGrhmpR62A7vTGAhDQkdpqQiTdRwAGN2OiTFxhrylsLTjSkV5NSA32D91zuoVoQ
ksrb0DKjQTWRmDKGGIb6zXIzPiPh4XlHEtCRQT4YUbuSPdmfPATfDgBNleKiE6osdtY3NSwhcgNS
JZEiI2NxiqDwbKA1h/aj5WzD2A3lL46hp1zcUIZx6txRwkeoCFZ6eVjNWP4E3x3tD3/XlmW+CeUQ
Cn58TZwSqG3ghLd3G6BQ5Ble4oIivS7m87qk41I0ZLMOlorYMs8UK7lvpEcuFGijBeEUuutMFRgf
EXo/8y5LRV67aRgXadadaAHhD6GtmFiOqdfbPje2uS+Re0wqb0wUaUI+kK8mCowzSPedvGPLN8zJ
S3VBR2lRDHKLkeO859S6IjlQ6wEy27CLa/SQNqYCXy5tuDmSVBBNE9udd5WuPvXI5ECd7bmelkud
5gTSScQgiFKV3bb3HePsg6pEr9iyryVQBZjmHHa2PFq77pShAaGcEu4RTxHpI5lHZB/w2mvLLwxJ
af1/wKkmZshT6S79adyQPk2F+H5f/HLVnQ61lxU1MEPvfT4zjv2VDYMb8GqTTzAzzzw1NdVxetMZ
k0Rgh0FZGq0BmPpOKNsh6rB8rrPcVI2bq1TU69pOX44N/MUSBqljo6/Hq3rltCCxBXGDrOCc79z4
VqyPNjRrWW/Pz+4oZnAqOeZLm+uNRK1r7r8hoKXv/Au7hJsq3AsiLYuzhtshOoQYSidBpDLfndQV
3OrlnaUEaw5tuc0P1avvYxKb1185zL6EZPix/Krzs6PTETuxfcootNFQ4VKckUeJHtMI5ChzFpQF
W8eWOxf0Dl+xF8vwO07iVCUB9bNfNTqijS6silG1Z1omIfegbjJOOOBzjqnFoWWl9sRgDqIg83XV
0ZysdOYrZtBgwweSj0ylnZ1Xw4wfINXv7MrllXMQTxnYf3AXUtGxXEOuD40REOupknYrhwDV/zMS
ulQa+c9HN4n3WFO1j8etHVP4zwZLS71iBbpCsHf+QthxB5izx1jHg2+eQimEkbf8QpFaXa6QHHSQ
y+zevLuLrn1Pg+0yjSdFgwxZFW7eLAv/DMeV9JDiBPsnpkmkW6DUAwEdOgqZtvxy6UKguFjuPTsf
WOgPfCKS5QWZTh4VsxBJstTW/wN39pZ71d12lRJV9NmBL8zJbQ1rG9z7LvuvmxpvQ/mbsFlE6hyE
bR50nIFjLtAYxsb5u1YGKGkcQwKlW+oX7c7jDzbCCCa1vvqZvtdSHN1Jm14YRziKb/Dz7fWVOD44
K5XliLTWUt5nB8OZCbuy+UxD716D/4803azukWrNETUVviTumWi3BdDzby1z8pM7zzQiLT8k+OOE
x9rI+dpUC6PHHqyoBTrCkqCEYKncWp8DUEnyfZU2FlWXSw6kaxhGEFAo2QP36JsHDSoaskyyUQNG
a9h1r4nMr5mewsuU0Jhh4ZWSl/SMoKusZKpK4AUR5pZlbB7aCgQ5lTLMgh+IqLsE4ERMR1bWIzT+
aPmCRVt607O5I1XfBzpt1ouXMyFlKq9znw7IOMMlbb9OD7+Pavf7BGfY64+6Xp2oFZdLm2fkV9V/
XBNCsVrnsrLvLnRW7W3YwLdny0EuaxpzjU7+j9SGpl8cPczXHVz57IzBNKVSa6dDIx0CGtcqsu2i
LIc1cire7aROZiBe5xHSCODUrYmXJ2DV3LMepfNL2NSyMhhkQRjKZCXruqffCMQ2W/MmBxnc02vo
xZny3UTcl5u5C/PYHC/H3C4bTe1cLKAFngdPu+aiGMqyNTLQzBRfOxfz9FkSnraf6D8i2QA+wXhA
DIuVJuEszjFs1Pw7tAlJCnw/KUReK/EVm+TntsHFzycyiH2KY7+ViFhEEytJoBh8MOI6ywMDdaH/
AHUUeN+LD6ZvtbYHMd4lZMnQTlVVUAaHrNJ8NILvQd35Qc5fA2t/M1ATQnn6DbgbUT/sH8k02PwE
M/L5T3ck1BMakNoA0hck9+FI2Uc6EbSPoeE7a4N2zM1C8lQRqeINRO9XMFmMGf1098xReViJKGBW
AOFIWCUbvqR7whfsAhP8uYEYq3b77HhGmFRAhzNOP2fuXNFpOk4HgKrYWXTerKJTcsO1UCutxVip
vgq0ec+heuHEht1w6gmWl4QM6IPIc5Fvg1cOAka9+G5pIYl7UAR0nZOJdxotDMh2NyNQXeMViCCC
Xv6hklI+bjlNPL0HjkEzZ3ZUVzqUJqQ64+dHC3doiNqz9bbSqvsy2SYlsMBJh++XS09+a6UZDYsD
VCi/12cfo0KALdHokhp9Uo1Cgstw364WqlosvhNkaFd/IS5TJnUyK/PekiKEpSlvQnEmEDmNoPfj
zMSC6mc/Vxi27V2aVxxvWagynRo9pmL1o0WdAkn+ljQG67F61jSCX2t9j/ZtE5WI9U5b0xgy0yTJ
h2H3eHF4m4TSvJeQz+MzaDrDnV0pHGVWlNxk0zlPul4dnNQOQngdklvkM/nr4wZ9pWT9boOATKrJ
8TgDro3Z5X0MDVRqhK6zvV9qarkpDE2xstt9qN/Z54igcjMvIqkHiFwtcW3YIxomuS5LmMAW3M6c
Hm1NlFceYvGDf8Pq31wlG6FT0mBxI0qbmedaYAiwRnjq7ViD66UqWCaf0DESa7FH7kp7hONf2wuV
pyEkoQCgcYmH+P+xTw8wHrMNDR0uCiXZaI4vItxpafCKVXuwimVm3sjzd3WSYhD6T/M420tHqFyd
kyE18iUekeEPZxDe6ziv13mmkBbAhWtP2ykRhcpzlZ33hupqZSWgIFI2xj25ZlflOSNSwYEbywU6
1CBIlvwGdMuivoH6MJjx/AydtIH4lSfTnw+XPwrPqcgJS6c+DrEKw7Xct9JNqNjMa374Kfnxcgte
xmyGv8WL6bhnR+PA9XsTWKjF1S/Xj7CTZ14S0WWyaQ4mFy1wjDZLX5BliYPUcT794+i7mixAQCqd
DlnKyUEBs5IYHNRtU+nj2XjIZdI2ATH8dFlHv1LUw+7xf/WMfVDe7I5+JizRQAAs74F7uPrxBzeL
RgEOJQHj7DOb1vN4JAthXTZJzV+Os3zQCgfUZdDcN1XXUwjXJpSofnfOWmVuufVHIQ6YNeE2+EhS
+99fl39c7nHl1xzNsc2xxwHCEOORgIti12ips0l2nqpLWd4DIve1SStLvSoaylgrKYL31fg9vgk+
SYBnv0ZIcbcO5hC0v4ldg+63fc74xriBJCehvwneaZrrREqfgWtTMTQw4ujwP9ThL1/0r7A4HBQj
WMD/VF/EGewFhrsfWFPDx3kF5rMbgp3pAiT9UuOipKfPIdZMqr371aXc6aK7xuCjk1Xw3SlSLoWT
5WBbQ0y0NU36ANK3Lh9Z+6/JHiv93JveR4E7clNtkHBkQm2gADES98RFuXWEI3D8VJKAJsSyBDDd
g3jtecWXtLljuiO6aJFAL/wtkbOOndYPWJJgmEuQ2d3ENNATpfcpZowFc6g+Y1HALpqf2RF5cC6g
IxKoJvVXNxoR1zQyhYNnwaviC+PVEURXqXtzCYrmTjLUtW/HzHWgWd+jeiecYginLVv5Cdy3LT8D
dWmJTCuleU4NLPGCXNzHHAHLNIGxbGR8IuUaE5RY8CIrLfApFjowjW/pht5BN5r8hi7x8wJet1fR
PHlh2wTr9ux9NQhwQx5mtFfdYPRW3AYUcyqyol/fmP6dIjiBAx/08sDdBCYc47+jC+dtJ0D+Hz2B
RcOPbI7LnNUJ/y38B8raD79KvxySAbYsJHaseekkGY5ddh97NIun6GMJ5TAmYQAOI+Y7pNbUUYfU
RYr/1QOe00Aru/kmcik4VVPhsW5e+heHJn7gIMMc2wWQalC4ZaYLre22tROjemUiAXdwAhGZP1dK
K3TlBNekeCaFkwUaF3IKM9Pwjeyvzrq/Dt3Jz1ggrNT7KtolTo8AYDr/O9UlVuX6VG2yrrlLj/dj
ucnRnGN78udpGc+ACIvbCzFDcbfrK6OvP9feTmde69IFAYPWhoMRdNwzRriTcOCwK+WKNpp1eF4j
7xcdrVpapTJitwe/TePqmaEAFTRqcPmHBQPRH2mTz+2pQ7Vs3gijrdhq2/eAOEsyDHP8lMGNjn50
L7U2AZfvFRoMJa/zOMMF+nuHZfRAncu26k/uo8n7cKDra2joRiG/mpruRJ51Nn1mgL1Uw1F8cBRr
iLCvgg15jRcG11hG6L6YVnTN4cBt1fFkcNWZsfR1U9xKFoXHnP/ZkgtBuyLJ8JRjlcOMYG4fAV8T
/68VgytIpZcMmIH5i39ZbfiRNiPzoKKG2/blFYh/f8oyRs42/5930Vi4NcFofuk1gIhytgowY4JM
JccFb75SwGBRMjQ5+2Hlja6j6sY5kuIY8pJ/6Y7cQbL9LsKznSg0A5qMiYv5yNXqLTzFn3wQ6rz0
IlqSA5CzL7S7v3H1OkAL9V3CtDAIvIHtXyW0FEniQpB+4xzWEIrkVHLkrTgG66qOltCr0IB6GoMR
wwLmDs7XWEu5RhUhZAMAk2XPGcMFU1vdp2kdaRmPCu3Q0/v6tZVXPYIMNMzOpAV4QnD2jRZoOBmI
JJB39r5KADif0/Dz1nP0EglKrCIIC464fwZYC96liCa66IUVO5GsqxUDsdlzeS/EhDZbibqxHXDp
2lnhxYgi7LSK1T6XAf1IvvXDlm7czMAnD3pqnF+zTNh2TOOIPL2irJ5KceH7KY7F5XIJ4kyZDzY/
4WIf0oei93TE4CaQ11vDtFGaVsQTRGoyCAKXr9PKRUw0k+2jmV9q4EEa+puIrEjVGAkVYUa2dN/c
qbu8U7vJXKS+eBW00jzfChY2NcIRPMHfkZRsSoMge3dUjAkW59pzdjlpnSzYyfwSeyJBMZQtez6V
0W0vLE6trZUY2LdAVZIPt1OBDMYYgwdXRV5qm3TL2dDIP5kNk8/ZrQTfN7kzT78/E2M92kyC+547
xN+oa3ug9mE/TK6OKL0CUj0WunizF5kJv187b3MCdowAlGuGbJG3vRaQvcM68tCsKyN+GHJgDVAg
+zZA6XmM9umu4jrnTfz11gq+HbSuEvCGk57HSrKMWzrrUqYF0Mp2Ryg3mvIflK0ltd7I0a9rZWBq
Vd5Tk8oHhTKeZJWirBklmkAiRKxi6FvuYxvOP7w48Zoh+MBbPGmf6J9Wj1uXurvjSXpCyr1g7H/S
gXb5uppTArPUmD8nRUcEHgtoMrChim0e4vpsbveb0etFloTE5XP+AABLTb/uI7ReGb1mfAyAenXO
C8sQB1Bc5MPSgxdPfWoRzoFLJNvS6uv3TWGgcanoTWo7bLEojpCzO+fsoFjvgX4HKx6t68lIg4w6
vCR0/Mn4cQVGekRedQcWrLKjOkTi3rwtv2vsH2LQnFRGtXmLj0sqJafca86T1O6qIq6qaM9tarr+
f0ZnE8FSmlspjXsnE8tqzcVBwBChlddquzEwMtDg4M+98keiYpjYcvTlzvFdFpjiUyaprhN8DxmN
MzTFaXY6Kil2hWqJZ0M9icvmKzf2MTE0Z5ggXnNOETrodjpae81qlZLijFZ1aufwD2M0PE9NwxUy
XMCHnfIXajQu6WS7G8ymLyO5TYuKHiy3rGOQ/w0Gey4JSiQIL2D7Ue9LoiNq/s9w1Iv/nGzjrh8M
k9ralObXZI7CJhCElhL6WAvQm92UVW0ACcVeGbB7qW+w+I5X6v7hL37G7bNHYtD5Az/7GR21h+KG
Wu+7fpGGIE42xrtQ6vU3rlT7tUs24qNdEh77TqHss5/vKoiyZku9qe+6PgrAvXbR7Vo9zeiBdtFY
1J9WGiAxBUB+u7k9lZsKCrM/G3R0tIpDlmn1lyYDT/y+hNrXpsWe1/aBxAqPPkNpf6+EZWzre9uD
S9serHaSaXgPVwm+A6ksj4e8jg8oruhi4IoMvnRptjtn4QWhcYr1TOt/F5cFOwCWHbywHh0DIZqR
Yf3vkhVpfclXJ0chACWX9n7G3KJ8G2z8dAHa7RPglfdDSX8t2PgrkjP2Z6DFOhpLWVEhsJi/Txn5
ZqDKGbeeP13kyctnfUqnNzDIj0pvBHlfh0XoQkV4ZbDMI4eOrOV0LC/cnjMsjkboJYAE3R9mTBmG
YyVIiff7klSTxOcJyk+LRgCtlS9Kv9sTwW0DGfklmsOw7tgB63FzYnN67MFYIwWxOPgDnJIEinlq
IUCYZkWEgSuEUCGUHBMLpDtsibwxyY+IWxYSjBV3D2M9LXyWC0ljVcT3/MYw1x88DP6oNyXbsnXJ
RwaDLTRDwxBVa2rtVEp/zvEk3hFemGVKeq/R9LUG/gajz11qdm+jDF0ciUjYpJABxiNvOYwUId3K
ISVeP/eEy+bSLe3MQih4Zid7HT5PNd2ijQS6UBrvucTEmKwC2KkTl3JZ7EAFL7gHD7tU0wVFwKAg
bJNIsXlQ4uFt270No1y0Yu/N9lZUNHjGDIwX5gtnz7GYrKevMSlTAG/paHu1UNRZLE2I4JPqYQy0
EuwwFzcBfcgXgt15FVK3dIEcv4xvC0Vp/BN1uuxiuOCxQMQTTm6qLyBebXy6BNao73Q2mn3JlpVD
3SxTEzb70GwPbYRM9BTxw/f3hm6eYInabX7hK1VykOKW9gQvJ1R8BYGGRByQoy5UftWITQifuuPi
WZ6lzjEfIf3TUuwhj/UvHo7sAhaI4qFT6gsADl9jDg9IL1FXO8tuE5azCkqUaQs97BfamNd0Tnvb
bnWIcjb5BrOGrdTwl56zhoq06CE+Gw2ft1KeyLwyYlOQCMN4Y55vKm0EGEddb8JvKUWL34k7q8WO
53aGQz2a78MwyPZgvo4xT2Bzt6x7GzSNtulk3xuuk3iNjS8nNYKjYiLHrLVEotSrlE4XQKo3kRBP
CPEkzEwsZLzkoCYT1pRwazCYhsI1hHep0H832mllmKVkl+nJxl7K9zGcdhM0keqGwehLXDkEGb6g
nCUDNmWf9eNMACOegGTiQ0w1MtFL1iowTDWHdf7fTH4B4sR9HMtaGsHrdvUuLbZHFTpAijRrYeKr
T4uwYYDnI/we5KrzNHC6cRaVBd1i6U4qLIUK5ku6czmlkezMxEq1yvHKnP2IeXNlyWq/2fplAwy7
pRzKcRftlg5n+j6twnkvz48LW3psvbbf6PcenXzTlhdzysI9prCipdkoqx9DkuTcvkrJav5fdr2r
b+jx+eGF4weIYXJlOnP/0okeRaithsXhwqjLGcf5W8dukGEEXv2Moea0VwGTUnu+4KLlygkRADQh
TUXhNI/UiT8VlkFxR8wQsTvVySzImQ6ySmebuvdR4C3FnPqqtpm8U6x5DNCn8z0TXNiBQA8Oy7BP
20cYQ5ncPVVvQu5XiNFVBHvsAeC+ptu99/a/uqgZVmVKXtlwx7zUu4DoE/Y9MlgyoHCYvS4CBS6e
/Vmz6wEMWhdf26024nnB0I40oqaUUiPQaQj+792LWsDLmiYMxdXwyWUgJO0ssTpXUzIIxDSKbe4b
PkiaMDjc7Jf5x7lK6j/IoYqvWEO8PpSLJW6JOVXyYXTM7nh5B7Uh0H1EGlAnzmHni++sNBBhjkZ9
DlF0UmJNo3vwJZgiDSk1Jn81xEyQ5X67my315PjF7ZvouuiNMHVeowF4BNEXk4Y9Jn2CgMquGByb
4anGj6rCUMdj9iQ8mU5nZgPlQ+YAuBoMtEjUK3jKo8ekYYqhN2dW5Sh2B/GDMxsP2jAttVUg3D7h
tnctznU83pD9jp8/WGs5g8dymlxDOJqaVvqkYqxZM4lO1QMcZfzBFKiIy/ATF5k7YPsVqHdSKtpV
V5XAw4lKreQ5p4yoSDZdPmGhYMGC1U66Hrc+nMzwHE/HvFc2LXt3Ar5MwYypd7IYteHftswmacZm
cfdDDGqi5b4KtWBFuhOUhqh4oEoTizMIci5NxXBHyreGrrQdzYMCxiYJ9zQZ5qRhUUhsymE4uIXb
fmry9frHNIBbnkufQry3TcHeo+mpvxeou2cAzl4HwSinP4CavUUw8cnPElGu/JiFPBD/QWWLyglu
bdb57XX2S2uLz9Y+1oN/jzo566AjsIO5LeLr2SxUZuJJKaqsYxcE1EHcy4o9Wpdkqb4VWmZaRPkI
XTGt9cDxPrKC8xe2CCaXcwgvAw9BItKq6X2McvOqF1wDpdAKe784ZJOCnTjVVAhYsE8diIPwcoem
1YjOR4CdzTwLvZ3bOAziSHPt6w2bDQxToWNOKpED1a6IaNavny51NAIxd++WZyxCztm1cm7aU4zp
/bh2f+PAeiOoM5YkIk03p8+wieA46H/6wp9tUNQUa0/SLcG+Q7pIP7wZqj5q3hsUJYXjhj0NxATX
X+r4BJTEK0gYIUVDDtev2RMR0aAaRLc4l/wewp50adf9LfRuj24vZ4UXXx8LTENQARMhr0X+D+FK
KODAC62vXNqhHmJe8cTpsKTDJQbzSOS2lFzeP1V0EWhoICKCCHdXuWNQ+8YBNhrOkyGjyTuwdF7b
0LNOThhO/GIHZ/cc4uekDdc+INBEgCvlMkoZiObKQzErKHSUjD/5rPkQhq8WHbgeIdcp0pDlyN1V
23h+L99atFh6HUY/bJQJGFPbHRIoM1pP/AaYRxYow5IPogK0baU7ql1hDFPbOjk7+y3kJbgYWN2Z
Jgy2thz5s+EpP9w5uvOgUZ+b3HZKFJRfpEtk5ft42QWh8EEUlttmkJbFraQ7O5wceCTQa3HyiOsB
NwK8qNN41tvqbkd98efjkKpE5SYuamOHRCSuMzgdtBVLM5ZiOo/i6Xx9w0THoSPUlw47z89aCfqv
gM2iM4/epIwUy+94IOWfzXcxbVV/mfYL95ZEAX6dWjmr7822ADBQKchqIANBYjU51Bum4+5nIX2q
AkMC0cfMjCDfD1gN7rhPYcSk+IIZOHOsj/pLzAdMVtyJTeOaeox0U4/iQkcVfvUk1rYU787bBtoC
hqzlQvps59dv8Mld8py2UtAb0D/B0130eGSWxPxoPgXH7nQGzR4I6W46TlhbJPWTRknQNKNB8nz2
ZC0mT6agGmVbu7mHCuo+8nWRUrKMCfnnKky47Yyv1aCkL3RW+/b1p8gKubcVdZp6eJY/BqIPhkoI
46csOTTENG3DcilWyyWbdHxojzsPPdJgO/zJ/qEbrG6nSwV07uVLc79EOMzJUMPc6qtEh6bnYH9a
nxKH+Ul5t1vKtYwzSelp0F3eJOwy893ojioVmc3R4uxFOjqWUSPR+aA8138WVgMh1INTLgl97k9W
cxAp2YWhhvdYuFBSzC1/u5shNpCNEaAboC0xUiPEQJIE/1sN2g3+DIFhhCurPhqlRHrd4mbbLVp/
cCL4VNh6OqJbtZ9fpG5ZweddPoMoqnJ8Gtlp/kcMCYzd4uSG95F05wspGxgJB8N9iEnZdy50Hyhr
gaaVvF1tw8O5u0PVwpAJd03qd/zfy76L8qDyNUAQMMcfziZKxDDJVSdipPQvjn0Pvlas678GCswW
B1kDembfO9VCFlfIVJ6rmRKiOmqn4RVwjZ7438DfqfbAgs8JwyUV2nZAapVQ/vngD3wiFrHwThtR
y0dAnDR2RILsrLCLsGAb0xSWz+ezviU/Ucgtwpa5TYLNzKpurDFZTyj3OdkOGSiWdt7hEWTzXoNU
eSsPDKVwSEv+buPPK3yduAbWPb8U3K1eZsSKCkBSr3TwbtFQNB8kfqe1vZp1FLBDmQFQJWisUEw2
ZJKRMBWkVaeywNPJ0zQhuaIP6SZKth3PrdBSOGh5LgsQQtncQVhD8900Ns/6s5sSTABt6CVV5Kbg
RLOcvdOZyZvAO0V0j+8vxFxONw6K9ip0j7QvYsnyka0/DjYIwEDSvHescSW+2hNbX2oNbw3BMTEV
A2JtAfNEZVYEaqbXhH7YZfZkb2R2y9kC2P/v8+Eyq7vwHmr7PaeutbKey1l1K66sU/ArLyY23dWr
nQhRTtKZWJPBPB5VqY3VYcVdb70t1/dic+XfrRMX6QRB73Zdjrn8YqeFkN36ZJ38f95UZ+OXhSoY
zi1zfb0ZKY4wQxFM/GzIgyLvyy1b14TulcVRzIxfCI/jlsAg0ZhDGQLb1r6bgZ7n2XpUM4ZG7RjI
3fNk8sCaAFoa21mny11YtufccmcehvsTZgeXLiwaAIEVlFvzfQrePnJW7sBSxuFUezMEhL8YVXU0
5bXdxfbBnBIKrY1pNa3OKtTSR6RBR7/pNVqPVAtuIRzeW2yCNyH7aHTp4z1Spbx6bhShx7opX15X
h6667Kcs3VR+SrFL8SoeWHpXXza0IMCiu0/FnKNU50V4onL9epc5zYcJufJMlf2FDsIo+4c4cCXX
j/SPN6bbRqlMNT3uQdDYn9xPMmARAQnQzyXwe7ZXzgm7jHZ7GiT8s6nLt7Cer51b5HtYSpzU7Lpw
AbAwZxTeh3sY0qgHDhvgdhbp77j8AwWqWVhPMnH1VTYkC6gumnuxuO/IFX/a/hU2nCMXHEJs/8U0
SQGkz2J5XbJrVRsmhDiknGa4Xisa6KEqwmMu0EdRTKdaUbz94MlJVvnAokqqmtIX0vr6BqGzX58t
jAMEEwjCX2Ztk6pq0M834HCuyg68Ip0oOm5KHK4fxoO904Ogw7KA6WNfHFbC1y2LzTCfZ3V8eyR5
XS+bO2iUYgEvfCXzeWVphUycUcwqZP8ZRs3dNkImtJPiz9D01ti5t32P6WKVgVhvJqQKukQchzkK
ssF4D4sCQRSVhID9icoLtqLrtcPSgSy4dtz+3lcgtphkYdr6goqPJFqgV1TedbZsxHzkhUANyHOE
BL7A9egZQEaxdoOEFR2rtI0zVx63E5WctyfknNDV13Rp3oMu6ZC9OE6Zi5jUfuXPPmBBZ6ZJphYn
YjfihkLst4UZhK0TFRIoGcTm+zjuJbppBz1Ta0VD91xrtroWsGElpo6LKEgNlJorHEQTPP+0hG+Z
0hoMV9oS2UfIa9KjdXjlaG+FDLGkeMN0jWN8x0NeInvVSr1w3In0LLW9EeZbrJyl5ykCU2QTFLVj
ykDn0x3vip/NGX3ZvtcN3UjunLbm0Aax+7El6XiDEzQpYFs/Jlye3BHSJDYqWmUWGr7iF3pZjEBu
35ww2rAf2D7VFOSF9FVad9Zd9qrFg34mRooBbYxWhjMM/1ApqCbzYHzqsPOHH8Lazx25GTNbhK0Y
aKRfbP1I3ICKkhH1somZ3ydve2kafpgVg8F4OyaicOsLxPW8RiFTmZGIyRsIJI6ZdG9aA5WmUi9U
yJsj7vT4WNu9wUZiJXXTCoLYsjFt4Ez85Lg2uRk3ZRHY11oi47nv1YUo28gYxN18I+G9grucv6eS
LcM0KlUTqqOc+2rKQ0jZ8S64oiRizPF/Z9IqhDHFi9k+fAgaq5Sg514eWeDxr67ApuP03CVzAnOP
iWjgCEreZMQw04cfnN33Z+W5nU+ZHxaluNRYJQrWDWDK/QNxKYf1bWZBZ7n41Qr4g0sCQsEWRGcJ
PbGVg4FxNS0EgqrOS0LNlTVkDptl1LUJSKtTv9RwqFqJDnyuoVJ2oJ/U0bCoy6gunKr1ffpF1t9u
xs9xkmHtifo2E0ZXgRdTCc4AJP70WfieY6wj++PJkTpIyBpk19jHrsI8jaGUFPsOjD8PLbpgMEiT
ORItptpvsyvg5PSG0/MgxC+mrLdGWz7YDt1GsRjPZ9H4wYQKMbm/OKtw2bgaWjAGl5I6aQXdzjMT
OnK9Ac2eHTDrJu2H/TKJw043yQX1FbgNAyUshVS00ipNpSsiZpTd63BQk+4Q3DwNTJpDpgT2V8kZ
JT/vV1i67+hgOJFAZqmoMIoPiuyZCpnLo7VmgkZ3DdgYO/JCIKhRRF/CYxzHfqn2AeGgi2xbgpF9
pX0kZRDaoJDDxo+m3F/azRRCs0+YVu4u6Qus3ba3btxj7UnfxIbK1tiMTuCmKRJViXJQW2pKVuqX
MF0Mt2G5kNmnZZKpfkKF0sroYPG85GCqokrH+EsyfgqXd1GuLYd+FUkB+dNuH1SliKhFcXbgNBhe
ku3dRWsuK0l+mj4nFPIRyHTAiMOncSWhebfMrOOs0UKdttAe6NL2eyimZ9zIiFhLkO9BWi3MrkGS
EmaXyzNiHcrOR2D7rr8mvTkheEg1BKgYPLkWM+hBHpWqGdtQO9TSMDYAkEVYJ/U5xlbU4jX31cBu
I/ilQ4olyMdMn+zkx/yIGV+/ReDt7zetL/raif/7p3RblxjBVQRqD2Z7t4HK3U1twR+b8lapsqz1
StgqCqkqRyvrF296e8z3nWt3CpA5cCrFoB9pLQ8Nun6GuOxeWugzmOq4ApnMQknls6Yg80+nREqA
gyuRt75vpfsR9S6VV7zv+rb1Qe9U+kPJUpg+2Cn9tmxcX0kVUSGkj1ZaKmYcqhfPRNWiQewg2foi
AHtna2CsVAI/5/c0j5hVmI5AN9EKuecBN0EhuQ5ZVphzOfi2jx2nydxEMMwsbxZ5fRloQwaXmM/X
9/Fzl6eeZVDMvaznUjIafcmhkbj4Iq97JeTd/E/MYBqMuumnlXCmrEXBPdmOw7CrZOy9FOMUW4CX
OPgG5BZM5S3okzkizVKNgg3rZz4Bs5VcQOoBtz1GVDgu8IC3smdxXzlDwnFMuDFjU4MMnkhdLrtL
PuW080tEQSh7oggTFTZefGVOwGKiyXcQD3imRJSDnLCKDRf0z4NPZh9535KJnoj/CA9sl+9JN0Lq
16Xz8Tv/VmsyZ35IjmCV4jwc4QWyT9SYTsSyskfv0OeD/RTAcXvNcUGC2x0VBVNzuOmGMUQXYbCH
Fae0kOwAoBBpUtz/Hv5NpxXsmpdxfcvs3uWvYbLv2WIK1rd7j3loxfpAdry+zNrpCJ88bP5CUBk7
5ScQ4RjM6/T4awguXqR8rujoiWYLeraLCMa2f4UqGg5aPBnfmYz0p2Dc5WzuaqAWdyxOjrGuPfG8
N0KiuhU6vBEj+toiery7WEJUm3OfP5EnkX1tOoBk8bLBSjMatZpEckOoTx235PEaPjDz8IvgbdbK
78Vx5w5dsdmsLn/ln/LpLLYluXys2AyMFxcVbXMRluBbJxkwVgWaZ2Wm0M+F23uXmpdt/sF5YDaq
kIikfQyVmIJoTzXueaE8OgiMeaOyNzdZels1Fh1rlGgVJFqCpKn4Yg9LG9RFblmc4w1d9TVfLDxq
G0Qd5XKA8bz5nZwPskxmiryQuhXVurHidP5eQGWoqSHKHVoq43fLIouDLtvYnncqbxY0ZB9V31SH
hl2uDv4P2uH35m2iSfXsBwrUYdIMoOTfsr9626OVrRikP4zCf3u/m6j2NAL/RU9I6mdOLlOGYfEs
4Sl51d3to5ggAgqjXzsLMrET+v4S8dyYRcmBaRiZX2FtroGIXQ33+Xh62GbC7etHeG1nMUn6xI+t
/e03EA6ODldwGyxRYY3D6MQKFONMBfI/yQBxrjwCKiWfH4XEj4a1dIUamS8zNyhQKGi5gsX81Krg
UkqY6sHzjvOHNQHYjd+soBD0CUd9fSLKKB8r61HowAsXVSTvTHo3De6qsq0i1xP2DtYMLzUVFEtf
qDVkY4Z9s1NkIsJHHakvC9kyXc0rWrEDAogvijf7MW24YkTe1ddovlww6y3d/7dufLnennt0jXZ0
hVa9W3MGIr90m57RDe39GUEuwE1B3GJXEjD8oK/aXLj3VziS1uubVwDeLV0xgUE28nn6tpZeQBIJ
cNXTQjYZRYDxeozrOQ5ysf2rVpRQhcGsAlNN/UpyOrTjd71KZLywUFJ7m3fsHJ69zXBhwuzj5xl1
bNLJ23qaMN5ld0ZARHIcEy7DB56omBGK0GidllTyUf7BIbgHT0YfPavo64gewLpM4whs/wxda8Pl
o5YNjBX4IozoyGO+jnJFCwIvWEyhOOvdrgTbRaumHYAHLTn5KR8rxHteElQ7ClE6IdWYTwq3+nug
ZdWcuz39jkemBBymqvCZdRAMO274VuYZM4Ww0P4FjKq9apEk9GJSO04lKMSYXQZ82iFX5w0co1eG
CiyLXEH0a8LySjj9YMg610auV8IvDmUpmLdz58uBPrBFrbHOBL/sbyvMmebGcjSh9I7KbiBqF6S4
AAymVHyHjclblsg+EJ8H/pKyAZgQfDIkUNmxgjfWiCvg9aUuZQSf7JZxG3vI/c2uKOgJuXIJ70qr
nO03jYq+qf+f/diJcgkTla1/K7bgaB/Epon8Li91dnxTVjTWP4X/T/eqKKgSyxdn6I0mbWJcH0dm
or1wA4YP1BVNfTRQq/I5IfUhU7DjwuSVoPHkArO1Wg/JJ5Uv4LnhXwJdNbF0H0+FsazeuxCIqZ7F
rupgnYX4wAP2rGEJ/Syjlbke51lCZaLA5EIDpmyC5PXDqAnkax72CACZi7fe2h9z3uBY2l58fyZn
ttPSkBuMnfNs677N0/324H0NFmuixpVZvc3eps/P0YMD6OyRaWmAgG5uI9SQ75uygt2V1VachtdS
EcbNRWdQDyXhSW4AtPcIafwxwhi99waCD5Kq8kLR0aSM5FtcegC0I2/NC+tr9yyxaD4BvnLYT+2V
CknrsVA4LR59C/Ox+YMgyp1GO90S1zSnvVHUfKz5x0hhFqUBtrf+WewcXFlB7aUdI5/X0fjD2DKH
jX7fwI5AgJkcs1Swjfuxd6anjcPWFTNJc5QDz+VJtDgbcAU6ogvq+2isLjY/7fGea5MTnqDdoyXW
jLdpUSHpDS744x57rcO/odedOiBqAtc8UcUIfhJn+4FzGwbXI4THyxYh9c3GWDUATXUq1tc91pFM
8bG/8h0E1ORrOJ8djzbARqiUDAb+QTau32mb54+IZMJaj1ajs6IyNY/PTULuFFS8mwWnIzlnpMdZ
a9n8yNMsh91V+q2sds/GDMNpLh5yc/+6r9bBLiLardqMzYEIPCinVKmIB7Gb75bqtRNjWfAZzsDT
ATiB/jGlDUNguDS6/hS4dzoE1DlCRYubBVpq+3u4qMRoh/dwjgA9f6mPliv9mpi9Z+pnGaMfpc0W
2yaEFZQWhKJ8srkgf7RjPkVsl+yLFS2FCXm7+N+kIZboQeVY8JygBoBwGQ3KCmx3X6RIg1KXXEan
EW4Gw/S7oebx36u1w0kJ/NBOVconrmR6d9WivIYpPCdl/Ubb47t/5JaZlRHCtMFFj5OLATDb9OdP
sdVOdPahye49oWH0gzkD43K5ToRDvT5uIv91oS3oP/azaAx1PzHb8DYtyU+uAWwcQ0iHGuizhZDw
99UCiR3B9WNAiniDivgrAqap03GNEjZHwp8667YhfWBUpsSCsqw2+j/HMiLoqPc5mLFp5s1S97SX
wwuzauk9sv2qE8KgZD3G1DIkMG+KoOgaOgSzmH9K1fMLpUeGn0/TcLqSh33vMTJlwiduxgJ9AOtr
y65bksPz5FQxmwOiyRk+Kq5CsTvaGkwi44MAGMF3dheolsWEHnNH+GzUSLYqkweNIpcPFu1egNma
vArGqXVTyR+/yzHqpwU3NCd9Vum/DZHIMeGgID0Yh5y5FiWguR6OnKwrTHddMMR0Iq9uNJwq8Dm6
vQqD2+HFLS9/N6vaxCS4THAwXNfBgfIRT6EbjVy+BQB2j5khO4WWd67vTXyKoODahHlr5KjCzfVl
8ByRtznUY6nYoM1ZOy+/EcgytnDXPu+zTqLf4jPVnFdV2xwqyaxlYTX1Nt1hjcGMLLQZr9Sprlqu
YjOJ/US2UjHU8ucXhLNCo+TevpNLQIXJ0B2vqr4dZ1Ywj02wXVrNFYmE0L/TtrgXiiUghuhlSOWX
MfQM/vLyUWr8iZ7oxd3v77aL9sbN6IDGqy442OILs+mG/cOCO6T+E9q7h+dFmRlMMRDdh81RBZna
tz6pVCoBHbC6nsua7RG7ZhhPYdBES7+DNuyI1yw5Hvj8k0ha0SOUdKvo6lZVMphau9oPCtOtcEnh
x9EYNStwvP/AUh4JoRlhtP0atQxlPVtmF8XBb1UVRypLYGEwAECdkCOM+DCGHdV7w1EVQhJIyaS1
uth3oSCe7MXtU4Su/3c4mezAFHiGqm9uXPxDEoKc+MMsmaoHdRF2iUYXKhKk2OBp+x7DM3bp2nqf
GOe1Cniu+6xNcs5d3NeHlzNPqbY17NBsRy0mj6/symixUDQtKMtyVOFphAaGUOgyaFnw6/Z6YhDC
jguMPlEscNRBSnbCSq1ExmLgBiiXQbHrpY3bXPEvj0itH/7cf8wjXEt1AjvvERUKC04yPdh6JZJT
6R/OSpcPOAgwmVdqngYk0M+VE8b5afcbZy27TGNFuM8oOQ4euNPDLwNqRVrIcsnXi3IxxXfgbrrR
LbUVqX4PY8qMAL099fg8VPA8KE1xNRC3zRWqgimC/SZzT1vLjdljO6ejXRPvzrjIkaiJ+uoDlR0Q
zDvYfO4xHm4Z7AxIhmU3w9gP6RNCz2xD1tLSqSnNlrHBDtfB58ZKskVfoe5SjD+VbHyldDFJpawA
gsNoYk0ut4hXEPd8CwIfxNpEyrzlSJT/ua1jYghI11Jhe8Li0gjGj2Rur/lzaX32Qn24MM+juO+F
CE0DNicaqzYEAJNpIdvf/hYep38SqIhw6yJ4T83DVUHN1SIR5f/zNIDn+5DHKX8d9IddPfHXOD5V
B94zaqfz50g+s7v1wQqi8OA9vgMfJSxNc4siUWQTNe+k7bgHcp07U77AtxhB1f+EMcu5CP0b2qru
gI9zxf4b/ra6iKQ0rmGgxOj7O5gVbj2thjcEkED4ytGnAjB0+lROMUnq9ZIRLzRCPz6EZ74O7lGU
NKktoLt7DfUC0DU5zu9uvENhCy9xMdSqF0f1kUh1/JJxA8tIJgdiitB0lsvvZ+WBCubGYoM5qJxR
X35TNYh8UyHkivvrZfeHPa/0Wzf/y3Vk4cwqgLY/lsGOOg0Vg1M+DjfEpFwZAtjgjo8X+N4oDLsS
sY3XSjMVGgboBGnW6yWSSVGC6Qiwf3DeS2v0sc1xVt5Y9bo5tlInBYJWsvL+LLTkS286XwakMsI3
nNgVMOyeF9mD/zx4iIuPyiOK1kdURHt8YKSIT1SgZbAFbGuEZNLXIPK6v3TrJAHeGwripCwXNEHY
j/TdJEG3PV4U6j2gl8ZOm3w8Ith+x5cuiEiJBVe6DKd1RXEwej/DjtXVDrbXi3AAAY+dlHpLaaiD
Rm9kULrn1BxjIESAvgCmWF4fGEsQ9l17Ym1eHmx4WtLEgn3RZ/nthuGNJn1MIINQ6zP4nNOqz9U0
Sb7ZDGxLA7BxodT3UxlWVMU4ef6EeXYATc+ZZP7LaaYU/I5u2Gs6tnyXh6/2tPHgKiYZOKN5xe7R
JgL82TTM4J08zCamncOtVdTLmkzBKkOpk8YpKfJ3OZGGSSHyMOyTtGQqQGiDuZFD2qs7Cj0AQW6x
mih9DlmXPbbvT3sfYx2sd61avuy2Nb3lge+g2KqSW3DaqL1FajZWzdBOCA25QvWF7q/pHEN2gTHw
1xI8r2fEtX2mj7PkETNl4JpI7zfFJiah3bHpt2Q2s8tXERk6dL3bj4UnL0NaK02hbGl+SRoQC2fW
DO/COp64Jrd+KcqjEuUuFbrWO2/yxswC25CBxDhGAeoqx685GrXK+x/azpF90hiiPuhgwHSxAsjw
+GAXWMOiaIxMcPmXb3iIaWqsnUETOtcqVo0QKG42YN6vgonPZVL/ARw7bzU9h0zQ3AzU8YoASxsd
kul4zBIy++6gAE46qhehcnRn/r45O9SSbxA1J5JkwW3wSpghvTw/StHHUIE8lntP4noc+U5OrIFS
glVr+VZq9GnOKFQp2uRldqsfo9iWWfGG1v1ttel8tT79dYfNd4xSBE0aNEVJ30FKXrxvocwmwY2P
9pyFDK88VUl6jpVnVShx7LgzWTuAwwRq27bDRxUuvIs+AAtjllRBkE0OJ7T/jLtrF94wG9LEJ46e
xgbKZgoPLybsq5TBy4Tu4TVlIc11Uk1NgxMQ7W2nRSPWtq1wCmngdTnt1Dy09qsnDs5uzIiEdgUp
ZtwxvGPvpi6xWITe8HEhh2SbTV7QqPTWTYkj1BlcRMnEQ9S0DChtwFnS9/DAYWjPq49oH8SPTgHl
Q6AbqfpP7sioGr85FQZ4wrx04TR52N0NoIAVoYAXYs6jJtbeRauJ8i9PELXUer3IrWLP+7arA8u/
yMTsIN5IuIOEenCTEPo6bpmHfeoEjalKnKERxTZuL0OZPoPsIxyDlipap3bg/Lq4bj8yYLNvZr/J
ef/g1jLLmqhpUMP1rHSzVT7wnEX4MYnv2RF+HinPrCEWySUD91faCy1ZEPYhPE91oGJMoJv0DUym
HwuaMTMGzLz3+meX1CD3Ta8XTrf2Qi8gfKjoWpsFdSKhhSsESbhbNa2pIBQyqUbtV0XwSCPwytdH
hye7BaY2vtg7GN8msFijB3EO5P9d5Zingk9r3GD7JxArM19JWTociu6dqA3srwPOoiK7rYwnCrrg
P2bS9TsKb+q27y4U6xcDpg+vbWtq+ynXbw88CPQJ3fRMMj6qjxKq67gwA7EpYr94/MaMt0CWkxRG
fzZXZgNKC+nbbkq2GDmXVDrZ2Gkic9uEv97NP8woFu+v0jFEAHEJTMwHkGu+Zt9x8IFOPIS7L+O6
VIBrIAFSkmrtw1aR62M2GhqrMhs0ODsC4EBy0GL9/E9knD+Fx5AeJJuhP3FoEqVUSFu5Za6m2Wuf
ki0bbHw5upHFB5ng4M9MG85ZF/68OVWYkm6LsLlt3RT0xJv0IBIEpalPFR8MzU2ybYK3RxJt7s/x
qA6gyc47i6Cf49GVoO+R4VTtyGEqRn5gi/+1cEeEM8VZpN8C+/9WrAbHCIxUV5ZeusuCOLIC6396
mTux6SYmNqtU2b56oMh7BouVCI22Z22XmJ0HVt/czES0uB5TiaKCGevi5h8A1vZP4SOoEIuPYyPb
vrzyRHggqIZUOov7QKvcw8ussHbTbwCZIsFbqGtgoK+qH5RH7I5ty38upkrGqgkZqhsPrDaf3ERQ
vHiNX9e2gPkR0lz//syTJQdQ+Wz4v+jNsV9AZcMikGa+u1/M/3dJjkUOb8/wyQI6nPKdvuPJQlv4
ciacH5NkbbafukKlsjldPyGmcZEVkPuzF7jZtlSeRiHgqpNRtZHW3uKlu72k/JCw/mfo8m+LlANg
hnipe7pI3hklP+n+6MxOxidAEyM83o7WHVg7q7Jj9u9eUvUQUMcRIYBMcj58hvpFmF+a0x0lggab
DkUnnTaHCE+imhk/y7IKvJwkE99YeIfN7VwSWJpc3O06+kw06fPE36Mc0fw5dsBcd2A5g1wBERWw
m6dBj26KfvOxDX2nTw868GEK4gES1utF/9UFXTBXcEJr8VQ5NPDUyohHxbrzVJGvxorrSpNl7tXd
zuwFqMTVhD0wEDq+TkqCicguWVR4gnDAjmfWMs/HGzYOfDydJJOzKg3DFkBNIvRKVYgzWrucyCL+
zW04xNTiEnl/sVieKQcBPjWw8U+F4JCs5Y3wFZyLnr5lzLDELqri/FWX6xJeP68AcxdYRIBJlrWk
TZOUHmNOoxfplLhClRDjpZV0ti3P7fBlHiZV6HhxfO9Xvw7eWBQwiekJs4eDygRAhKmdRT5f2+x1
eIniIGuOJR7H3hO0wtQBgEPN/DFe24tG4IYqlIOQhJl8YVLK9J3fKHV+VsPJTY0zldX3Ztk9VWxP
emVOJgU/yKVJRBlQ6UNadxkoDS+Pas7H8d3jOJ1cB/f0l9iAEGERBmWdvH+wcXz4fCvWojV2kwm6
hk1GTPNqqC57kplie7pHKQxav0pjpsAok4pLCxlV1RZgN+esyXt6A9DHBQnt4NO/A1ZcgUlbPdW2
aFuiDprLatIkiOUr2Q5bSvPPmucH8Nn2aryvtVkahDA7ivOFkVB7tSaawDLOYZswcluj6mRq3pPT
IK0bfs8Is+AnvrAjECLE0Xilf//A9jkE1FLjPQ+mBdB7u+3N54VGVDPHr+j77S0Nxy7glwI34XCU
LftJ9xH2Z3rlSeg2ef8oLmjQpL8YR2d1r5UNEuXQITU3im+VYjCNln3XCHF/4TB/CiDeA9qYT1/O
Gift0A9Mer5XLPrhqwS6beHNV4fM2EAIewRIdXxhJ4p4GXc/HUxdbLCBKarg+8jb6ocoh8T8tKon
67nmwcPDN+B42XM9MVWQPsRL63e5mSR3WaCdu5FIgPgRkbvF7fNBPoqXhNkzwGOTkV0BhCrt6WfE
fQxNAJVfm+hq5pYMI6PmcC2k9pdu4AHRSM6cLS4haF6mVA9eVapfEHEXKr9vliLdxJMeqCAVB3Vf
oXVPGgw8yO+9/aJl5aPBudK9gdGfZPhba9bZrf7OilXGDn2oTlm+U3JnlV4nfK2kKrh6J5NaBV+L
XhTJAvnQrKpy85WrtNTC8WLcn9z62LE5XwI1c3Td9UoDIQvbA7Ep2YC8mxTKkpG1jS3J66TS9fGf
T7nGW/F0E9Ph0F4+BMVrtrYqTcO+byDpZCnZeXupIl06rs8Y6G6NYYGw9gzE4YfLsmvTVU4zDu/u
n5RL7RH6B7CL8YhwANjdEYPnN+Moc0Wtmgs/g5XDq5vmGAF5J3WWBOuq4bg9Tc6Z0ufTO2vSGhLp
HF6VibnrL9Stqw3UR+6Tvlnpzlv1U8hTnnXc+cRbQOkfXIxMbaXQ9l9Bkulh49RKzo6vjUGIBquC
Qme+lWdyvB8HWJO4w5Rvb/hXYX75VmvNOTPMoum99HBdImGoiXfDPFAnpPpKOSEa1ome6KdT13Jz
NUyU77zSJw1dig3IYOioSa48zaPtkF+Ih4K121KeuyE+poyG6gFXqbEaNDPey51H3dBQ9DT91eio
cqYAouhuvk1I2dUhXH6SO/bR2qMOnvdITPu5RLI6xrFJj1uEhFe0g9CuoMvcwygv7WPRXWTvuDMS
XHQLTe+7fgKX7X7wcVZjEbvICkBYBdXnLbmjJXa7mYZ3+DxCTHC8JuXT2NvI/YPwOm1rO8bLMcLa
oAHpXZDHwzUw0zwifiYvqNVTvyUZ0ItF8SNgsFfOOKF1DyG3sQNZ0vDfBjQ24n5GjVTwv5U3mjjt
90Kf8OGdXAZEGKq4n0HMkWXwpRygJV0Ob/XhVhFPBTv1RkolA3xchpVCBd9dwZfVipb0U9KWWEaM
vwUPA6htNFjrVsVlzXfotMPlgt5qo041XM8LdpHCBsYtgrcbgoQKw1DAF/SzZaxY8GyXxxD+KrvW
teEB4DatS1Fpw0SmH/VRRb5e70RmLMId15yOE0LXyWDlFelJjfz1Gv5PbX4CW1CcyU1hRoOr24j6
tlhfF0/Lk94f7ESAKPmtav9+cZC8Eyvg245RDQDgShb9dys2+8HHq0Uf1nZlB8gqabXFM+9BX2I/
0WjRyx2kOOZv0hq1omEjGmKc3EZK/UytJW9vafE9b/j1Tkq5Wb3P2Io3HmZ/5k78jb1ZSxIwaPnH
Ci/9wrqH+i0c0Ju6PAtHX6tUV3c5qT2P/W+ZloUmRYO8cIi1RQ061a5PmmqGxovwTVTXlajMY5T0
zVuhVswfCQLDgq6KbrYvDSU9XWgYkEkw46ElwMXjl6SEjpPckGwG+B885LqS0vPD3PJiXbAUkY2W
N0CxFH5O0G/xkpq2d5/3h/eZV8TtMoJFBLozxxYBfAG4EkFAdJijdO1u3jClN+OOYOHaYV4JhlTM
T9YjldROmH2SPfnwcOqIEJ4E2XYZBF8daHjNrPp/L3GqfsUvMNLAyl/zq/Y52CTsLfvgmIE2NDm2
mpkx9ZdPxPtQ5+/SXx+zT535iLVD7e+U9lq8cKCRUYy3KlZvlT+ptIXdyMYONc5Vegb6bLh+Zd+1
n2jI3PcmM6Mg3L0NVa3+SJ8Y51lv/v/9RhZIjN+sxtSQIS0N7FDX01YzUFvWarrvugUC7URXAamV
855eU/lJSF4/GAMc3BsxahX+0/DsK2TfePWj+SkqXR75m6kO5hhEMnbgF1onOe0Dfow880r6xdra
cz7rqudKLq4jYgAF4VHbzs604C6M/6cVYEs2Bw//SQSTKV35mgNFE3Nu+Sog7QyDKKPKUXjETmOC
AewxNANX9QIqGvgv53H8cY6FfABUZ52f4IM8d0kq6GxtYc0XB+OzacNj6tIFUkvfjr16/4JiRBD4
bMSTFt8B/9AqahACj3wBVvx2qLIycF0vf0cK93ly/f9jrsJId1insoshZxc/Ij1S0rN9vcImltZ9
cUCv7IwxhWhbpOXUsViyRXprCXJ6njhVfIejk5usPMeEet6ite8dr6OlZX6nXt+SGQaEt2UwNG0c
USkTmtAzdNriKO9zRR/4rzyuEXBNnfP0bdGhDKpq0OyOGCZsoXtSJSBR+8X+/YS6w9+1AhxazJdp
agMYTfBZ/vMcp15q0SeMsKzusD+TUXSq3qTLxXHS9spbT/f2BeS6HKv2TN9bvRiN98u7mh0tElmr
8tHVtBCyDCFvKjfpS38VYBUllFu7xcLRwUPyoIY2Rus9Uh3XIwkSyjFBkH7l3UEKuxZQhRfzQcOu
8ZWFhNJS/t2LXpj4T+3+S4356lp0p3axgwQRlUF9Sajm+3kYqaNoUhNCxiPjiKnkGcmv1V8KIb1J
jdSSDvIhimgArKbMUT5IZRPHniFdF7qU40T6WBhrk8GVZ4J8i5FyPrCV61aa+U0ZtsdNaP5GFLxc
17lDCySEYUAxQHxv8tRknp3W2V1sGct49B/WnVDVay01YXPBU+EBj4L1XKEl1dMitfjWpnAKV954
5GyIb33heHcmX7XAY84IfgHgbWZ8Ut3ID0zWpk+tQPD2FiSoGo8mzuJwzCrM/xbUAER0j6M6+t2n
yAygPZPBV5mpDWXO+jr4oAjO4FXDePQ7m4msUxxzp1FWc9dzPpJrd0cLfZbgskS/LTcsKyaHSCKt
3AzOpAKbbmmustzsXEFQQvV1xKbK/kfgLTCHEUs2YARCadgr922DR4WTcdJ9jRmSqUFBtRymJPP5
ujOU6qn5Ga2bmK8luher3AT7DVrQQlqBw3MFyGD0t+BClSu+AJhHp0qYiP/nUDPpxhMIohwDSGMQ
ZBV70tknkZshvB9txY/pqSDauOrzHnM3W/R9ydskBfG4ucZBgfc2TLCprkvI3fE41xShfBD/U50Z
dVQZN/QfK+dG1PWo3cbFWtTon5lIPd0WcFmboPdyimEI5jJILUBxyzG9JeHphoFVBj4SawsOFept
qMR6fRzP++iebTo4fzKh7sBI+PAfBtuSnxa0G7V9l/C644ZQtXUZxr9C2D9NjBZDl/3aHdvhhcyS
jKTIDE9BvbMR+HfTDHh5iC8q5mndhul7Q84OvmuY5o5TdQVFCyK5eS7z6S9bmJt4OZ9V4GsNFvYY
EwQHBwVqDuBxGn7W48/nii6WXhmTDO+nDXcqj8lW1Mrnv9s0vuxQiO5+s+PF4nR0Al/aq80Uu543
NDkfStRwsRgsVRCHXSuBQQtPPcDfo7jwGw4f5gaZSXNIEIP+4AHqqjvngPEPWZMCpFYznqm4gbfD
+5oXCVEFOK1n8JTsHVonJW/VMnrlVw1Y7UTrlyayO/GJjqkLGzzvTHKq1eYBtBxBVb8PySTyT0NF
nJK/MaWBBTb6piRXShPm7pbqpr+wfm4vuCRUIzesdCqgoKIbO6dNIqmnq+8mjk23aS4sSYq0Uw/R
bsr7xFEMa65MdvvhjL5fQvclPmox++CZ+qn70e00T8iQkvv+spuLmGn3BRFzhIWYSyroVBrZ7smk
A1xWorHxwjh4n92Ob1bfGa4las6hdDd/pRrwek3/wtRooOzXNbKRICHIdGXgkpDq2mP/Q9yxWkq+
Qz7LbeTLl3jBu7+mQBI7Qk0l2vDJxbVEyWxkq77AQ83hkZpnlf2EtbnSV1pK80Ht56VHONIrp3rc
oXnuCXq60ekLe170GKM5zyQtIW1FEZ6yJZ3pLkz72tNAXxU2kJt+jKAws0INtJt78OlgfeRd5mhf
5p1dSVXTbCmkit6XGy5yFr2Ff92f6YZkQSpSRM01DtC7lYj/uXiALFHYG8zuhAO8yWeKT+r6HLmG
ucLVIPPIXkUAFF9rgAN3EeeGzSr3LL4SWzaf7RzWoy7A6cdpzSxz+HB/t1HXX3arOP/BATrMeGAy
oO/ATC7up9RFg7E6McUXQwMO3Raq6H2got8yIn0MU5q0rfr3r2HUZmZ6XUYNz2b+LjrtdxIp6u90
+cnDfzgj1zJIzfj4p8xcX+qk4ImiiUiRFXkRztpdkAXhDtc4mphtviNyEmEEHRjyg1uiHmKlhNUF
uJocR8MYPDhEMW6cJVK57v9L/DvI/cehvRvbR2B9ex7V8O5sJxUGK6w3vQ5iKMLK7X+03MGc2kRf
en9cJMbIF1quah6r/KNZ4v1TRjbDvTNLYP0Hnyvvt0exFoVK5DUy+ZJq2GgR2PtxIkVLZvEBF9o3
mfI1wWzo0GHYKfiTpIJmS5DkA2qKJIjWM2jX8wdUEwPCYiZ1LG14sGO3ahRDQ19DoHtXELl1tq9T
CUYyePcsiMTAi/aGsMCTryU2yQbp3ja86wJrR9L5RAR1UCykBiVWI6c24GMMEK+nnQ6Pk/ma8AC2
U5DrafauYIiwc0DyXZNIiYGOgw2w6W7JyFaVeDepAVDnu5agiQ69aoEV5cpt/nTkWbsxTnTqNefk
QzlRdeE7LuLv3B3xAVyJ9vA/ImQVNraozrTcQ4haMuo1JSqWrBT9Rzc+X+zRa8ONZhVr8WSUNENe
VuNrR7soKYY4VkTtk3XUg6ZsNOaTHhNCw8t9MiZisD5ardq89JFs/ox+FULzOEfSKaXd/ScR15s+
Vhlof4xy/4AmjGNeF1BM7EtJfK8jstGCCnjskaNaWChWQxLu9AmOCndIsaan+pFaKGIudqEkZl8J
B1qGAPqzm7FnzaVxkZ+kVabhkBjGk4eXauExiHYbzPoWaqWrnfCbYXI4fQBrrcgPsqzG+rwc1tvo
VxUkfEbybBp0YoVDtoAVmN4IYNiDRWc3wKn7r3sGAraepAKok8FD+8mt6DRD+lokqgq8dOMkwLCF
s00KjWxNpBVNnry9+R69dmKZDGPpbTZCapYXL1+pupc9Dhc+IvsWMhvUG4XkSdYyN43FIlDyrGWx
jP1H5/cwQagt0n6OwR04mgsyOridBm0CjUnOxtS/8S0+fbV1ScLF8OaAVzkqszJ2qTO7skXK8dGA
8oOF50Vldt7AjAfBhfI10c6VXPrGV8PKiKh+ibBq5xc6tpYiFvAHS14YfLq6B921Rl7r4dRqR/UK
uvD1C9q4TBg8TPYczchjrSlx4s1Sy/13WhKhhOdPkMYp/l8yCLRJMstup0IUR+5G0GYDYbkpcXMX
1m8clLiaD4sWn8YJHQ/ztNxIWl/P1WztsQgVn4wGod2bBl9ER821bUMe0zQmUG/z+gjYK4XBERJv
OaJnUjWlddwTMzbGx5ffg2TESVX+2uVRgeS9anyW1aSmREfODi6xeeBCMoKg1OnTRjV7SGUT5Zvs
g/ByR3hjf1oIGjtS4N69S2MWA+PL3EJAY3U0VITpgYL8gbQMFePJDta/6Nc0z9B0DNr1kmVlwm08
bMO736sBbnmiHgCxCqP2uvaMAhgtSmCVAWbe8m225J1vwGUmzQKcExJzs6eUqto0v2S7EoUm6Qwj
1gOMKqF12OgG+/wASuBubEGFWxzXHB6gzdtjTJxLy9+n579Sl6i8vGrXxgoflD/bM5uTOMGu8Z2o
eIDpgqOYZ8DPeN58xY7IAT9KOPluMKjqudv8q7zjWHlpOR9+ICVS3Rdw5lKWqQNLJcXEv33twWVd
Gw+FdJmY8HBoTTD+eLsAl3+zqPRegrEwfQHQEy2jpZdmm2rmOKJ/WAdCsEa65i5zD0z0+gnKdKQh
NR4k4o+mk/OsGHKapGBTvKb2LHmrIP8xAWjMSx44gR/uINHlVJfXzVakYn3VSdoTiBq9wtzazR3r
YjqnXkXqsqBDD05BFPmTsi8KC0JqOVGDQbypO9Iehd3p9nd7hRhP9JoiImytwI7wtLL/xwb+YbMi
K8gpeGwNqcF8d/hO2Uf8a792wlFXDPnkWEZYzJlpmgaVbk+jWmtqBPZtbfabvb6mhNFXOrwvlQ1o
Dobgd6uzJdj3bjBWDcO1pxQ2P+jplbnNUgRI57RXt/NEH4uIgbo7TpB/pBt9nk7vz8kRU70ZZI6Y
tC4GONqFSHXqLoBEBKkGMdl30os+53t5eR4H4HYRHzTmYALtLMhH+yWP0RGwwIEniZxLa0K5Bx14
Bmp485JmNOLDmEDkS4OQDZVYKtvSeA9a9ccUrMIK9SkrJdv+TvygKJ0ooNyaRO0mM3smB+xWg/u0
tXJ46jHOrIkzcbi7FSueIaqBbFRVRVN+AN6QhhvAQSnXiwYXak/H7//yKf5dyJ5N11GE21ekWcQ5
M+I24NpMtbwyXQCbGjDgjCNvFnysUhnytorWlUxNVO+ZfFNzpoS4DeO/fVqx/ee2p2KzP55SH6Js
NAts01zD1V6mHX4sExjbIx+cIrjcSmBtTKBd5UXZPmFA0lkEt52Aiqsd784iYfTapaxIA23mRMNo
udJhy949KTyUNeHJFPQ3/FYAphHSqlhAO2OrjkD8md01qfnA3vVGxgNXdsUufr5BQC9a6qeWYoL6
2M65CVG+tsu9kHsoPGYMCcp4ad1JRzQSZbquPPqcWki8Qcmh800Hgi6+HNXVH2sp4cFGIOB3j6/e
dL6emGYMU6QwIAaTVsaFxXY2lSySoyt1MgL2pAeIr9Sudr97S1aUF1+UkCKcrMTCSD7QYuEIpxl6
TbibVMvLCtgZ/iWQOD1K/K6NV1Fsz9lvGHbwS8zZlCC3eacN6TVG+JSjwMab0NqE4cOibfxe/xW/
NmXp90vIZ8JQiajpLAx2XpB73Gm2ZZzXbsHja53uxIqgtG0KQnWTW4xEEPlYirbtT0DOliZkL3tb
VLqyv9uzqe7UT1pUChXpbSjmA1VLNy8nYR/j0654UvtpYYRG6QaUo41PMrfGaw3xpn15/ZlCXOa0
O6UBUb6ek5R897GKnF0M4PIy8c+l5sS1vE9d3mxkFHA27wvB6Sw7hIgXIxAyJwywjmLNddreeDT6
fqkbgHCmsH3RQpJlE/gvDeCmxswB78ULIu8THIbTJvNq3EbD9A2d1jHmCJIHwyfqf5vdTvJCH2Xc
g0NGwWY7ANb75kV+GV/rTmR3k7VSyTmvDjmtOQVT2ACdciNCjQwp7c9NkUA1r2RJDhzmHD0EsPry
svTSmeeowMld9iwcLUgAFMoB2JHlCyD1qZIk7Y9jYlSGMGmU2iRqwX3Nl/OFsYW9GFpzfm86Uokk
F3VnVF7DnM/F5lVgjUM4nbJWgzjBXYMck07B1UFJQ0Pq3PolCc9pCsuxQXEXxxyWT4gKJ0tDOPi0
8rjC8jOOoDTMGYu7wI5oGc3+mb/IPMtknjByHm3WyBbphQv76s4Opy607VLhQKrkHySozPwEm/ey
RGDvCFutocCsj00IS5vww2qpm1C6NtmbfcIPZlAUfbXchp+BDAzFF1QufqVVvulA25l5rFqcsX/K
XCAWvvXl4r+dmYfQaD/nohpgQCKQF4vek2S7BHDg2TiTmUAo3sW8tCpK3Uy324X6/rS8lia0EM3l
AiWN1dGj+A35Z5z7qAdZeSLOXa4Qlq/ULY45w6mflwEERLNtefrYLqB9hhlviKLoXkrpDzLEX5Wv
gpmRirK5BFVjNeOIhAN6JTIizV3jNaQzJDBieUiZdrKDwY7ZKJnUcH5CdNbdOQxGbXbp3YTfD0O3
QZveH6c9du3riVeXX3ZhWDToS985//WF0Gs3ZjwgPtC7ZsV4iTEK7vv+R3evzVMtTgz45Ou1tVIf
BFZBs7YFRYqTPiWrBCU+gI0LPoF4O8DthMSIi45Kq/Y9acKr94zEsYFeXo7J2/hArIZmUKKqugKL
i8yasrElPyOd2QDozrdKd4+Gf8CgNDCYwK/bpXJchNr1LO3WOeoynQ+8mANUTLTsC9AaofVhYO51
4zwjFB7mvxFeVPGUuEy3f0BJO6dU6If5hH3CxqRct+Vrxej8ofHkzkhsEldh+37pOFO90/tk7IYs
tdIolnUslda0zJ5cViQtqkjG+BQ0cQy1JyfUPFZRpTb1Sd7lSRaxzW9fNapKXBQtaQaX7hMx8j3g
3cYYu6maAzxMTLA4FNLX1TwLWc9qy4thW7sWnWQ7FlFjPA8anFHAonxFyQZ2v0GHRQmKcQCeC4UN
49A3YMG8WM+oy3E2rOxmHVoj+eBs7oOnOL28MJ+th8abszFvTHi4J0XUIt+FCWzaNMlLRZlPbcGA
B0SGxbJzRGoyZQ21sOJG+OSisBaIETeRReo+x5csKzOIqqvwUGTxw7paDYJL+wYL/71/Do0RA9sH
1W4ugyz6uBKvH0wMC8kKBcI+PipDX6LnrHH1sA9w9LkPDnXywp/wKD/maMxxQLKuJKoar5C2WJfP
9ktDMJ6ICWYLl4AehfqDIkWYZQv/6NWxxnquf9i+TmpaYMcXr5gYxyh9UmSl8PuPccI82a7pkQU+
iuCqvNvfmVGIwa+CRHFw0OrxzzGxDtvcrQtRwLBuWA4r9h+7Bp4qZhtygR9De44MAyU5Fcoo0u23
wnDjRrlYQUXEW0TmiiNVOO4H5g8ZSl0Pl1xZCfyc0wmCFte2TrDGOIER96KXeY+rvXQ9ezpeIp6E
315GhKSNSw3b3YJ6wnm5kgxWPfu0tmnCYpoYtIhxYlIcUnBvuOh8Y4fFMKs099ikqIEHg7yn2nTD
XHb3FMqgRZPKiorl0cl06ZIPM0RW4WhZkxRXrzmg3oOqy9hyAf94EgUMU7YOLMXFKfnL9P29fWl8
1hlfPsQkFK+SJV6D3Ch+2GYS72AZtdrq+vyJ9vOY9Df+AXvkTFv1uftRefuAz1i2AX7eynVP35kg
kzK3RAnaOHF/A0n6+CUBPYV0cg0Qxmnk9x58eF33wx0LPXSrjmagB+2WoA4N2EKmmJMtg/6Dy3yX
B9dFmV/4Ll71fKopj8KBAangP9FxFVMaPr5XLYeTbRzy3OjFjvYwJoXrzQqf+X+g7u5WIu+fjPbo
fv/Kcgo4k56CCKVza95zDPEjvyGpgIhYw8k3dP2q8nr4mMGR9FyqUmsE0M6uVfG/CJNbOOL7wyEx
h3RD2foTtbp1AqGf9jctFz1tOyuLkSrwxe9KGNRo+YuQ6Z+rrU2TXoklUQHNuVBITgm13Jl9L3GR
qjVi9BfcxeLpdthfeRzI2jF2wLjZfLTyyjWFukdNJgE+G0sivcLZA6Bk5ezyxJ6Q37UWc+1CCbQ4
YLHRte9YtY/+gtTA8LtDxkdqL59E3cHgpuUGLApDUQApuVtpJY9Q/hVvRD2aHLmcCpaDnRpqhAov
RnA8aAvRlRx14x7z9EHff3Hhqn4qrMeIb/UeAOMpqoExiGVggwqw6Yn+TURB1M9tkD4ySLO0SGEW
ruxLW61P8p2ZqjaKeva+vQR/UDlS6k5ODUGu1SkELPuHfiy53UNMJIyTjYDw0t1+WqTc9Q3HxTLI
3o1LwqR3Kc+86FiXX8FaAUkQx9XxLmSw+nCq1bNzG7lIvH2a20HY4QYBpMxgAykL2QH1KIrbQsDo
OxFDtNPB8GU6Dg655ozZ1fLGSYrnZYf7/6L+8NC7s1Qr9maLq7/Th547Ajm8DCJY+vsdjmTGV6AN
ZP5dGa93VFirF4q9LqwVojkbikDV0gSubrQ4PAbDISwkMh8Dcxq6sblqxzA65WV4PZOQ9MZ+DIxr
cOmkb/7u28lg0UZNGPbAUJQ2mUop7vXmJyh0zgqKKPaCyLi+nTl37cmzPWIZAsJN/dxs/2/+1m+z
meSUq4JBEo27KzUDHT97IBFYm9irRuark34iHIEAEvSoNfPP9kbGW/SVOmdJ3pvhiTAW7q8sa7rE
pl4V/yL8ohU6B88dhFa4C+2+nFp3vsBlE2em6QxP36OfaYnL2s6HQD1xlz/pN+FerUbtI+0hVfFA
Zdv4x16zfCP9myuPl83C5yCN9+Py2W+w0UeTU7Kr340PQ7u9SMz3OmCB0MJuLGqC0aCfc15ndymj
OrNkBUB8T9fBGlJ9BlPplOD9ChVnukQZ+eQ8Y+oarv8QfL1+gprb8N3Dan5QijWRaDBFbwwT6j//
0Nw6gJTjQRzlV4QlUnVEF4Jtzx+KqI+873G0HHifx8lccsPLqr22MIrIS/oHORrB0HC28E0gAc7D
IAgJW5SA/OFfcGTPmUXFmsGhPsuqpB8MFdEdgsNYrXJej8KsAKygF/1i2e7nYEUKTksN0ieQr+ap
BFYgDZfITJSFYKU3LQWEhKGqHPryQPyODaHIim2Ry02cMl4DRAo+MY2TnPh+1oDI6DTjgVUcVW/1
5ABWCS09BCoOMJq2E6/BiuTp8gARWTOVZKXXMhNRljlojgf7iqZNQRD8xMNwr0wE6zpCsomKEG6k
ii16fVRGDtm2k4X3hzy64jxmhDXfWcYlpsrk8xs2KczFQp1N9G9A+ZpC4A7z3sbjNBsZYu9pmKV6
1hNkTym9UemHvmcldj4lYcPWIU4l906PvsqMaxWmJFXZgju0Q8/pHcJpIkPIbdKe5LoTFurLaI2M
h4gi5Qx8V0pI1obxb2H6ecF4GDq3Ctskzwvdk3367bk78thxccU3AFLCSsqBJ7i50EBQFq5jxt6K
hRUQet3zu2PRiKvmKyh+lPWIPDxpeLiJgGa1ijXqbNC03EPrNUCkkqP2ymOTjvoP0DIILyrgisYh
wyv8/dHu3tzeQbKe4aihlQ8zbNZb+kyZsh4vyq0L6Fz7ykLBFkdoDzJJCrE4g2kabe4DJ7wzrtw4
EZtLh958jZgfkcKFbN7WlbQObSunQ9VhsWczBQYvBxClXkGNp4PxcHG9xgdKZOUXRv/th7Ud21+Y
u0k6Mt7Xf/mhmDvSqnanboIvDaixTQNvGKnCYkUvZc8QWDmoqR37fDd4kzeuXOQs1MfJ24VTTIsI
5HfSJ1klKQvkjkTWqFXVnHhZZJNelVYPoWGNaRoBsd/j2btwuauGWt98BGULBV4y8eAJB/LoWMKd
F+bQfF6UHmIN8jK8Nbj/1Rydzl+JqUOC+36VpqtdUEGEcy/GYtBkjm/5ePoSdEaCkBcIW1kVMiac
xoQsaqvfxopca6wgV8O8PzMDm6V4Psa2swgDqgok1VAW7Pk2ef1Wo4+/O6ocWUgm1I9hZP7/v54n
I8//dzf7DeqNFOvn3ndMrCFCRWIo4tpCrHjcBxge+SKaWZJ+zKzxsY++6M+I5KTjCfRWJb7tcUTM
kLH2xmzmobWvlGaxWLxhZi9rFkNhKfJQ5i3sMBZSjJ0O5upV5ZHWrwp5NhYFFqxq64qZv/L2MrkU
HyHtTXc3zibhVE2UUXuQRglwxrDY23VqUQd5vAPHLRCTpiQE20sdvt4K7oEWkPgpURBwWGbips4J
Qx9hqwripCSmFT6/XAXw++vEofA4cjPL0sR3GWnNmbeNbfpUD+LUJB4q6UM6BEioQbh6PElaVJlL
SmjJBN+RzpZtc55KdbecVgZl5AmMHduuvpJG9NJfdqJA5kxWyiz4AH3B7iamQG/2mEolDSJKFxui
RsH8q6wTNmb3O5XpGRutmdJxg16HYwWlVM5bROVQDtmzgXVpfL+/uH/RnY6fBi4eE6rQneoFQFOl
V/bibEEs2s8LJwxR8TmxDorjnmBaOTW1iFgcyq4h2ZtlCWbWkFibi/ul+AO/8qun9sq0+C6mhco8
n+OOGBDmr+k3G0PrQGknquBABgvgf4TEMTOtayq2+8bWxx6AmUqFNHmiiIkAUF0kcNjDjxdpMBzN
zW5bUWgPBnu4JualUu0SzopAdKdDuV8pZHlbrMReyd2Uw6UX3OI1j4Tq2eFvPjtEAwa5Lob4ioHO
eahluoLY5pphGrTqDDN+21ODGNpeNGTsf40W/v/X/1urn2PMo6B77jCVeNgFbtWyMyTX3j399mtJ
FTO+9OHYnR/c7KqeTw63SERH539aOnyLz+M4K8R5roGN3jttpjLZBdRG7FiO1lu1qvb+SgFEV+Li
YrGfwQe9TfYM1LAKQ0yq1iOJA1RKiQ2pnB8ZliTUPnVfsctEOVtMgH4mv6xgXL8pqH28S0jJ7Iyp
mUVOtbMv7xcMxTPq1NvST8rob6YRZpX4DPlv7uFtZmdWr1hp7bfrxB+ar+7OT5HmId0+K5NAeo8b
RIET85kkHpokE4l+LMj61+Lt3fN0CAbAt9SZD+fqpJ7mHBtqQ5aqN2hb//BgEh96pa1VvFN/pbm7
8ZJxxHS8CfhlziRWYI3qTDIQ6AAZBKjbA9sJA6VPAPk1NEcMydBbbchoOo2LFWi5Gkey/x42K20C
g4b5HZli/nJVbu5eyYx/wouXaRRvB/vva7c+NEyFtJ5tp/Odw/jh/1rqshciLvcDwMmg+gBmdPhW
IYT41UClPCzg9rndYBbA5uQO7HL9xw1eHCpFpCN4fNOInbRVaUIC+t3KxLXJ0v1tO4EN/oj056gQ
x+C5EDQG1eI/vtcsHdWqeI7ZXSuyZDWNXJ4OktFWvDHzB/+LQR6xUDJEBYM2dXsHyVW5uqeIOlPF
z/3M6zhrRXMJU+3B7jHZkoH9vjOxOtvtTSLQxd5DlfrT3Vn01NbXg/H/rcqmHRTMXWeZfonMhnBk
bcyDwEcIiDIsfpFVUxCEajvWfFMtJmHYnmhAWqGyVi9cbFsjAALLcf8RDrgY5Tqct+GmqAeX37V5
eJrQy68I1fVPkNEaPVHxR6r4RpGJIhyHmOegdZnzj7sNHdhpQn4GOuyJAcKJ23koaCcHIf+AAEt1
1H9WpAWKiuyDAr8ogYRdHrowHiOGnE9YTiE3MWY4RES+yO3q2cUiN4ee9qtW8nkx2XLp2V8cy3rc
njRqy8xKjFQYyelIzqlYrveS757qRtIOPJpSBznsBGF5IC7/McKU1ES1RmWLeq1MpWdn72rlHUm1
zgLP5zEg57Cbf4sM85x7Epp1sXjbttJTt8cbwE80XzkCbjeuhjqTtSFjFG6aF73301jk9bNTOhMY
nxDo2G4KMdYVz3ccXr9cgCsWKXydVyK4Pf6/+7uBswJiMLP64jHgqGhmTf6tl/KZcYmgHm6olDbS
pBk1GRRspY3NMDHXa8dWoNvBW/IDZvLn3sqYGF4av5ZAHYHph5y0hJeugofLZSOffO9z2ujfOd7V
+preQ5ZT2CW5Ai2zwslsrPa6YeyJ7LjrO+bI5Y12Bt1z+Df+/P3mRqdIhT05+Ysd6iilbXXJzEuf
Z43PqCz7GEX3MejZwwv8DQtHo4FxVYksqSU/0/+Maea235mf8rWbm935ThuEpRtLmaZcG1iEY7Yg
+GKXmuO9IMs8l8pPtBhwOWt365FGGHcbeyQW5qGVTRMcu5GrSjEgjRQrx1XnfyQR7JMBfjPcBFSi
+kthRlmVfd06dd/aAnPp6vEfhJuwwFMhKWjUGFhJrle1tWvJTEvQsKrdgFivW8GlUEKrwA+Hvu2V
ikSF0Rs8k+wFHv7RCweO4hVGa9q47V/gi9BPugIY/sCen0QDacVIN2v8+ct2abtjm5aooUV7g7U5
8HSKTOQpxdZTG8OhTuM+2k4JB9Hnutp5e+MYv19Q+zSHK3Ui5RCGWg6twaoYtMVNO+NMRyC/9VU7
/ejQXjvKPXStIP4v8bq7/LzVfGNBgU0JQulkRp0vMTWF+y0HSpmHJXZIwKbduKN82JJJ6IOlZqN6
VTzod4E6fctTfU/YxuetmQkvAyCGU3YzHNhV2RYV69z6lo5vr2vyfYSKm7PDyYSZzei6iAgnsu80
eBAmvYih2wMHSDwKLhqsu3o09ecL6hr7K2yWLONHVAQMCkK96QCz0wWzDb0YZYPanCoVD/tNYGju
0Ra9f1E8W5poD1R3GRSijeJAMmQyxvRF96Le+mwFnBa2cTlSr8HdXvarcZfhW4WZXvxuAzt7gceL
iTdM3mUfxymJMnuKazYiYHftMUc0VjSKYXUtP5SeUcTYCK0GOy2ChgVLn1srdCb+obb59QG8iB8n
74yYXgzSpoY52JzMIip+DfvAQPujdu/Vf0FJPB+FpOMhu2ptwJ0yef91I+UV9/UshDpp31bPxsfN
ev3M2f+ScNkPKTVhufHRu3bCiSznwcOFFw/mrhslAARZsCwOck07EpthBiDnH3aGS1JNABYFFZJY
vUZSEwWtRit1kEnYsRcxso/DfTcrkKEijI4gU0jk7aTiO7lVQ1JBwxUDnkmfgXVn4Qad5rfgDXc0
WxFq+kUTny4ei0Tm81rsv9otePUnjuQg/Sw6+d3ZI1jyFov/qPIYZ88u9QjKLWTxzPmREsV39owB
oHoKRNJRt2nwBQ4nlXj6shVPhKK4NzrFJ+42JjO+cHZwhd3JIjrX3lPlMTXmgBFqLJ7zyqwCSic6
p9VGsEg/zCfGAVxrhmKHWjTggEGW/bQBxHPJ987lmL4a5E454zUsjgRXeH1IuoWe1D8rTUolyg2a
2/Lw/GEVvSgscSP0UQLpGLTvECNCmHMYpmK5y9Ni1zwCmVY+nPGlJg35qxPPI5bK1OQPCtMgHlPp
kGQsEJJ2vU9ZZd/F5hkZwd68dy82M2RQLiAx4yrsaeMr00GHDHIHlPICBjsmFoufTVED+InziQzQ
UTFoRPDAkD2n1aYIQQSJ4WCzhD6RxkceXe39Pyahb4AGf9XjUbBSLFM6cL9SOnjMMS6Iu5NdPqgj
bvM9Xd3KtCLu43LLu9MGUqWsITsp2aNFqiqW//1+1aKnDmTftIjA6CH0YEMlUe711BC3TPoj9TVm
ic080r1CgmaLtWF7pnK9cWwXnYZvRAUeeCg+LiVwwdIXMGCU74zoYiRtHZZ14R3YERgXjk88+Ajk
7EUntNh1lsg/vXUpQGrMjKapgjnpnQrx6j3MkjOow5emfzEqgNCbnuAQGzFmcwgIjybno8TdaKAc
Jq+iGPTOOLV2S1x/sXHhLcJkVWzoYT+8UJlaJ4QOXMfuez8VcjPMKSF+tNNYhHSh/6Ui58k/G4AF
J+mGab4Ifq7De7snd/eOXb2KqeRlAVvbpLCl4nYMlbo6w7lO62pbChfUxlahcfli1bu/qCUjbpqs
GNoG1IW7MGnPTm4mTBxexmjlj15Nqo28nXbryFzExlyuC12zS1TQYpfa5wrDRLmiAsviBFW5Na7z
CBDq/ZtJaqExzeabAq7/016cZTo2ADqXjSESwjde+28YyGfrBR5/kw1yRD4VHGBnWjyQg213s081
o6ifGPUD6lDCR4ukvdsBmzl9eJHmp4v0K21c6qV7Yl6Qgw1eFpJfO4LSXGgo3up8FOvKuVhiZE0q
/AQtEowzy6xmvniwsWOEkGVfN5Tu2SLo3dIBZapeGLaKbQGsTowgc9DFaxuKSK0NrE0ylCqy6y52
dcUHo7RMrjXDsJ0nWmCuZrC3VBtuH4usNOru5G+hC4zjYE0wnMclvO4zEnF4jZCOceoAdUIb+QPw
YCSsmMnHdasIda0NI5tbpazxXHwp3v0eiWrVYczCaWRSl0q8geHCrOqPPMqibBL2pRTkwHUvvaVF
4QrLYXdSwN3z1etqRF3z19SIb3pBWME0pUwxhkxXP7gs6urc+r71IFq10AlmbhmG34tGWWF7hHHI
JR7uw5brs6+ru25O39w3oSN1UdiSPpapRWH9IQSgC7oh5xIgoOBLGTJ9FXs2xa6n+Zhpz1s4lV+y
lfGyPOU3mPKpS3p3HKoQ/clIqowyMJnbjw8etZFlyXcJn2r7pSSosZEwe0DMe0BOn2eI2Q14j3pj
obCU1LB9XtKEMqtMHvGgjWYvAOW6//hXQ1oxHCT2B05yPFzkXP+L75wunK6k9khQhsdXIGYgZbUJ
wa9jR6+muOMaHuRaTGLfWgExsBG+tpzbGKSF8/9j96eHz1caqVb+f+9SiSCbpNJO9kxOCRG00cQA
xP2h0FKaRTEVXjXv2M6k7ysN1ofLh74NzbOrW5PVjF4EwQ8jeqrUm3MenxMp3NVvm7FSoBAetnsa
ZM+cXNTuHQVMAntNDFkp23xspeQQnGoJE8eM97eaaH6ZMRL4S2vtfjPU3BagFHwBssdtcImxMXwl
WpF1ojE01iJzNzUCxFN0/WD5Q9vDcj9e2inyY3yEe7LNiaxe0HFmds1jLd1RXVU5Pu6IQsld4S2B
3cfTq0VrWob8MUspr+9qoXtfBN8yNczaulIzI4qrvbwPxR+ISDHVOYSQb4xZS7MJDBnVgPcm+C3J
u73iE974vNJZnhkS8uPnAYqHyx6LoWk62ZyGM5dZ0Hscu0cYr0jjNheHrr4zE/JSq+ecowuxNxLk
r/mdy9BSJ1VOGFud6vWnR0j+fSEGgvZLLiA71zpUp7sTLoWhiFp7kwnDrUNYhFt26AdDp5gymnul
vlCNYyTKHCVkdn9JGNcYWCyH9m98Yr8LYRgupSVRWkpPYnq2beV5c/uoxR/hyttETJdvFhs3Z+h8
XGzd1kgEPupLIMgLv0fxF7Md9za/n9QU1qZC4VPTeSq3ZdVwFTX07vSZV8UpMYPYfn+ZFS96rOEV
V2cT3sLTXBZB3vAdWBH0+qXRTNmMuF91TBFYxrEzqshOZYq/VFgpsRvyokYEAxySZCWSOVz1/lpC
1s2ppWaacTUJh1+ogzO/v4CeM05rdAOGyZkaB58600ab+aWM4Qs5Tl6au0uS6IDCPT65UUHaJuXI
rdkvRMvP9/gaQvBeIaoPcDNrF8HuyoFW3TGseytBSNGskUIPJjIWm0AeNj7BB5P+CmI53DCxV46Z
oiZQUF4F7f9ePQMIxjtBnwFIyHwWFRgvrnUF0vLOmTJ4F7WMZrw8SRpmYAb0S/6JBVrKNQa/qX3p
T2VknFT7wpNlVU2/e26xg8DwSz3wKMeBBrrrzRcV7RkFGzuacDezpcZtN90AtpN6wvItw+dYRfLI
9CDa3BM187Z8nrugDuAW2mW5+ob1UA7DyB6wdYzGtBMoSPFqi8zaPofZ8a3eabholc339hfWd7TC
YRoKxASdXZUXlx3gF7b7AP/Tj0G4MrtSZCl8haZ9MEmtvHx4/B4xZTUIHD2ZDExnfqE/XdH1vh9z
qGVN8i55Zezg9MxF96MXK0zzYsZtX1SmnmE4D+t9ybaxjJ0GSfUL/+OFmzYj1KLBu05IeEWVVHam
zHdgE0yF/iqpk9k32SplNc5pIhXyfltxXvcrM8Crl6QsvSt3SsI184og7xhmkCaRcQMudEfroxL/
HYOi2XaxtZSSDAEHhRdLkkdZA62725X6OmOilTCh7dfBUdgI3p/TZUvXhdTVvGQ1nAvoBt7R3ilh
Fu4WytgCATUjCFBmIjY2g4nrS3Gf1Dee8r4RpgNq6y3bW2+O2hwh9KK9dgZ66H2bj86ZRhG7tGqz
aEKNCzyMWSbV4Z+XP4/LEQqDa9ji54ryXhkE7euNFkuOZ3i43PCxGU/4vopGc5BCGF98AOXlZCuf
n330ArkM7KCd3PFaTnCD1LyrSnbwtUWElnw44Dj7XPL6/1Uv00QNGCzXPFn5I1uzQt1xci2Gnq/2
R5Eid35hZWStYkyG7C2n+EwlsHwrq9jJW95kDxbI5SqripzkwNQtuFlj9zz/fsORhL5cE4fa7GI5
+w9R8U20qHMynV8UquucBPb+VeXCM7YaORJBXX4aWkcQqXVGPWHuHa3iOeI5sngUbtV08EX90zAG
MFqDWQktPMgf9nEKT6tchioeglSdS9jjG8RwWTOnrBvVRLlJJifMsjNPBA4p8NcvuUzOs9x5uFbc
q1KTgWIYxb0hxWV8FfYMNlrO7/sAV/CQI3U4TXZHe6/pdbq5aFbWDUejHZ3MWRsWGLeh8MT2rEIw
UtRa9xTlyI7VYwq15nkkmOVxiwmrnqNxBrBgvpuzp/Hbb0zKkHaeEbBolj4eNLVOuenTptUWzAQy
wGXOyev52KARavBKvIlTFmsPSmHdEA+T63bfLFrPEMWwc/MUa/Vmo1rl3l/1fieJgXKUHj8HHiFv
Obb2jGvv6zt598bwOG6ruOJx1z8ZcLzEBsFL1DjiXQsVbF6iAR7/pE6+j1Ao3NIOhlZNWH6WVkw0
qvZJjbGJOhzbzjRHY4ySgONBz1CT8KK2u1McMB+M33o+el6qOXtT6VgYQ/RRG5D0/R7DyTBCD8kR
qGCyo62MlOQIdSm546C+Qfkxr1ogUlgXe4SjsOxOHteyZvQ+veZsdMN4wIcOzFYinnW+ZZOvrSwl
4LoHy3VqptnhodKD6Q0HYmGzco+MkUYDBqYNwDqLDPM0nIAMLBnglw9oe/2b1Zci6nSIu5sFgnQa
u0nJS38hiZGU+Za5DKYsdoDcVcLaW0WKSQkKkuuIOBgvR9MrPt9MmrHO9iDecnELtydGsJPHUUVk
L8tp6CaaK0/3D7Dej8TpxlaXV/HcC1f5kBIOBOGY05bIOC3RDUKRZ9uutA8mvQtgo0t+dkPkpNyl
Zf9rbIO3qSGdtRL/MPu1NzbZ0eboDC0BwX3l+c4iLADYlGEakDvsO44DC7EAg8HEd/jFJaD9eF/w
x2BBO6H33rWr+Uh86R2RslxXtwmiCd45dbKRze7Fc/zHSq5wWhyb9JlRRe289Wl00hAWxxQtX/Ft
JCCrbHsXVrCzCDGmA4g3iivswQB89EC7JRUK+pw6z4tjKlnGCUUrFqAw0kys4TBbItmmK1kNfd2e
wH5SeMpCsS3id8E6+82a0BLewlivaRGADO8LnHRCnxsXDAY08SEqtQFdXcWQmZkimwhG+5RMmw3Y
WEvksFTB9ZI6oNkT9hDZRBD/xHhL5clZ6i9phwD2+z+CL/E9GFbXYTc8L0Jjl8kXCHCxEzCr+Qnc
pJVgs0mQUHcs37+bxJaSjaEFYOToEfzaG1TDuRvhdzFda/bVeAN3yK2iaTgpDBn/gF6rj1sCzbIK
IMD9pNIf9Upn2fUHO8uvzFQVsMjWqkHseoMvFF+NMHztRf5BbQ0p++yev6XSYxbGVtnec5CgnAEO
h1oA6i0o4JKtMacv939HanRuKbOviQkdKfZRKvEn6sxLo8oI0gMDaRL8CeVc0MToztY+dtXV6taS
Vj4nZA7o5saYWk21Qyu+tnAl5g4eNdPLDnW+ieIFe85KaVCV07UaO/D50PJ7Gop1UB7d94DpBQZR
fRLZQwTvzE3XKn/KdjKbQ8gcLBZ6G+JH3LTIfV7PLtigCJ27cmHaJFTP5bOiDmUgMVoRoHN+BTg/
ZP2nUVcD2WS35b3LzNFjPtNhGbW1GrsI5E9KDfvFg0yOPkZXPGu9e/5BeGLaf7lcprxFQdFsxxe2
vkNFiMCEWeUOW9Biljz5gQYXJ3D5JyNKOFHKuPcZ/L8pF+fvzHiUx2TegBb1KOnlglptSjZFVl2+
RK363LoUn/qOIPydc4F3OQoblqmTfKy0de6yuwAPSMJOfMsm/iNnc6IgLPY2XEtOtG2ES9lMVRHX
UPfGmlRPYg6RaVyK7JjeO7LaAATtOPo8Hvugd6Kh8oT5H0gHgap8OrW/kZz9P8Qb/PtNY2QA0NwE
c4YECNsE207CYU628YO8qUOKiAdKAlSBwG9nMjztTBPGwMYvEDZ+204ZYJArf6DxxwQGOvNiNmHq
HObc0nLGIc73VQySaNMZBLdHM7V5AwYXajLhlOGTxvt+IerhFwGw6rd6KO1bzJBxyv3HH9m7HXmI
1u7nLfIZmkHK7LIl2/FlSA5PbpUjgfJSkwD+O7TYC3kRdqcLlcwBk1qF7wBrJ2Dq8k0aou1VN1M+
+1p9Nmn3z3O+SBMeNZYSq8fvVJC689oRu6/3mDNeehPMiNrmVSyI9sdZ12tWF9sYHypD9Nte85Io
FjCE0/vdSCWNPNAwosfnR1dVaP0RuDOVzx1raWsdkyrNqEykcwM5RymdCaIisyzpBZs/QVbGOFph
VL76uecvouYy3oSUnB1nKW/RC8cT8ew8BWffC6grL+qSSQ/Iz5VxifjN5ne6/tZBw8CxcHYWpEsa
LZ9QnV7Fh6julUuyriddXwTSjrftJwl2Gt+OKCQ+Pa9s1AIpi9CbZZfOc+xVgblAQ9ze3T9Wexka
kZRDr7E+NjJOE7bGRPTQqdp977xwh1+w/tNyZ8U4dFLsiBfjILWpGwbiRnUMea7EzpB9h4LpYRNV
GrxoR6BMJXo/zlhh7nIF70XlaPpVDqx7IRYESCKycICcdj9npWu/pUElt2Ms059WTVIRlD7fyZ3p
XB1NBLEg0LjpfTG6HeCPIsW/4XfNuMy6NpzUnsB+py2duG9YDtpysgT0w8sjoM4BwoyBwz1pcYZl
qT8gQmmGwEvhXnoHyrZuPdZVGLl8tFszzJpObsHQVY3q7gUIov7NVEeBqo6daADeNpMTZM4TUdoo
KcXH/SITQKwlVSF1x1hoqSz6JR/CvMpuFLkktp/lEJBgfUjPvZhoQjJS8Ag3gmrU11fATGQA2nnu
3iRNhbPtni/e8LgF11khktxIsf92SlrO4kUC0vzzSV26CNfInQ3k7WHWvQwW89COdquhyePKmjBJ
2Nu7W+Gh+XTGWPdMgXNXuQdOT34Te+2uT0YT7HIAOPZasuvC8FBiBafVnL2AcPLLw/nK1xrcWOPF
AsvYZK8fxWfIwUM4WAiPd+o0eiwuAWsOyaU2ZDwBwdQc7BXYVTSBIO781GQmpBi0L3OW/CI05vhX
9CIO1PEoipyDurRVDshAw3VCW+GtIRxJvFFbgAUpNOvCy/LYw0Th6bvPSSm4cI0KFa9bjwpJ/oXG
XMnXv9t5jJ/MCqyqmmvnItPdKlF2DmKs5OSKiJtHWN+cW8iK30S+ZxBN5GEmI5RGiMbC+aHau5GE
8iUyxALsbF+yV4MQhvtO80q7vsHztmfr8Tf3pyWZSdYKo5ac18RId4FwUYGq46025JC7Mn1fkxJJ
+YfhDoYdNVoZo63cqsMnbbRSv3aUEvnYprBpVF8vPKijjzLhiHt//q+1pALuTFimeC2ewX+opBTj
7u6ksoWbmaiz7HQSf4X/JAwvM1b/6iq9SPclupUcR8LeEvqCyOKF/Bw1YFpS1C6v3kRdLGmML3Eo
DLjzCZM6/NAZw4u9VooAF8Oq6gNHR0paVkH2INIO9X6qROavV8gwmJxLLVHx+yo1MHi2KzjOPWy7
gyckP4t3QRtCdS4+ghxD50Ybuo9sxcsthHrKfCD3zOkOtqltfSyrVeH4yyl+DigNM/w/7fYmc0ji
PzpiUKmZ+6+2laxp6t1UvSiqVdQLlRGjMsU5qo5UF42rov4qn40D5tN15u9c5JvdJQNfAkWhjCqx
TQwfKIxOh/SuScnLJUqCR6eO8WXlCABpuirKd3U7OLLvDXtM9Q4cZw8+tvQmbNqOmXFpRKS4EnPh
PjmqXbdNX1ZSe7eYWU2w1oKywQbbFF/Jap/qmlsstISvkSbrftA6l3cUhe+Z+KgCAiJ6rUCrDACL
r/Sk11f9MWT5kIDyFISSJW0rw7SCttYH1+hxzKW67exUSEppNf5v/kncVjjkQ8Re7XXPoOOKEfXI
vUBePB5af01Vg5c/AyWHmgrNoTskWWd1WNg6YvQ4zx3yFo0i4eYVxHaFw+d9eKjBGPcGbtU9X3t2
wl4M+Z2kODsww4ODDNmjn6AHfdqL6gWpVvSq9cCf0oAWs9w4WScKPr67S1fxWPfrMpa2hjmR06DE
KM3UG9ADOr6GXzD+K1/tgcCt/4pgn+j3jhVtgDqPJzEtmcsOu/8PLqHAaGWbE6neP1Isylvzc8lT
tbXxmal1MHiRsggqx8U7t5P/GhaEuDawNrUHkGEuTdYtigHEcQkWq/C7vPbwlKn8RYhipfVj1iK8
++UXLgtUFTYneGFVtllOXgPMi1htkZwj2i9f6BC7rHhmputRPgs/OgqiQ5nDivaCOpIX8z4DJq5Q
UajOZFuKGpKiK60dbTKpQ0UYKzL602WI0aDL+uX4iDe6T3DqB00BDyBaFtJKMUYrjHx5xxY5yF2R
YZrb31mlExNnYrdjv4AQPbMlmzdk+XS92XVzxm9JPQQwvytYy7vh9NIPyvs4HawJuGq5yMs7ZDKA
kYt1aQzwW4iMJqwgXc4t957N4uwHwrtjBjkODmmZ5F5SgGkp/HQENvfGIdM1FxswN9q55TQVYIqv
SgTY5mfzMdtwqI7SBRaEY9vrqG2Xrj0icxtU9DmLO9s/wLM4JyTeDd9KmvYsS+6Evj795jGZ4fo8
OF+85QPhVyTZxnc0J1DHOG+754qQlVKEWMsSNfEIEWhrtR4nLeDEcFZxDGC//CD1l77DKDt82y0u
xZebOBf8An2xuF8xgdDyHM2OsiIPfQ/XSGDW6qS5PJKzKdacYEAXp7WW+TpbDpzzofR5YeCnTMke
u0ci/RB3AxY19AFPK7DcFpgTNfLH0IuhcyyDqRE9LMm2nH0WkgBD41O8kpWollhBTnRJm95uVwc5
z4mINtEts1d/Mie7v4uGA7b4/9J/17jOBGx52Ep5WdAqAILPCh2TVWSY87V3LzHXAKDyadvqjs8Y
LoX9uYhb8pnj6VSgz9KKcbQs7rvXWT8a1Gvc20cqQID/hrvaNHW0CquPLC4z9nNDAYb8Z1Z//gX4
l8Uy/lmoAB/89cQqHQFGvtL5V7vVqhVoSnRi3bpVWdr2P7Fi6aE5grNv3XKiNNpVCMwNO8zIJFEI
QZbcy8hxugR7wOD/YC8mf/cUxmQVy+oMd0iWoE8ro4whwYwUDfZtim4fnJHsR45golKcxa528u4j
FIklBVJS+1rrnPdWmBFNdGjNMyN5a+ebgMR6jq1bRv6HZZHpscCvFQUmTXpwbAnKXCiPJUOqSTtc
sRm3bn8HR3aCISqzAL+ewcRmZ95y//UHJJCobTOQsrUeI5hjMK0X2VNOk6/dyb/jjXLYA/p8LHwo
4/qe4+7/pQ1NjHCdiS9nCZI208l+R/xN8yzbHxX+g5zCA7jxBh84yRedcJe95/iQGm8NK1smGJI0
JVF+y3JsS7Rlvz7DCk36NE/HbzrpBIkuWA4Ka5g1hB38JdHui4yM3Wep1gYguyHNdkXrtlzjt17N
4r+xYoA1sFsJfC61IHq4NoQ9jXS4V+6iTrf5ySK8kKcV/Gb2tq0r0QzdPdA4I/yXAtdmalleoxnu
4nctbGKlCMHP4GOZBZNCC3rgEVHLJsHcUrVrT4UlFMR8iWtNqT7OQmKYg5AfMeb5PbwsDH/kr8Tm
lCxxd/M3iE1jH/BI5jrhVAnr81IOeTCqWU0oXz6CfajUJ0zDhyvXvxe1P7l0TVHAtghrdZrDvAjV
8n61iUBc80TrrcxmhoVBV9/QWh4jqs6ND+u0fnlF7x2QKpxWKxVUoZuE962mM1kMDa3SBEH2vLmq
/uN7NuUyiGpLVIAMbUffSjEyaOXgLfHbrbQVJCTluhukxgSfGdKWhUw5povq0E/LgOstbw+E858o
CixBgJd+jC7GH+kNFH13RRnuTKUR2A39SdWp+9A4AYWTRMstkwZ5xC+035+wogxHRq/2MopJqDGX
iIduEmqa/klIKs6CbEefaG0MyVQ9aomfJlm8Oy3/zn7elkzKpxix6b22tdKPCwgQvBGeMAEZGqfk
yx3fqj9ZoIwEeio6bYa7a9eynyanN+GF2PtwcJalqVcFg4osIiy7d0ZcxftV1A/1jvgSrW01yGmn
fNHhONgonm8kGYMIqxWEKskT0UM/C2Qp8pBfgsWWalLVhCSpafoH0iUkF/xIPZdgiGJlFpoancXR
M4uzPcwb2wuHDL45aidgnJc6UvHaKsPvFd87tGUTMD45VBHr0vzOwyu7UHcfyafKISHHIneYp3zp
6xsBWVSY7sTo6MxQmZB7pDvY4RIlrfvXdMPASFv4ePKLoGt5042Oz4ovoIiiKqC+YQBnf66eSXgo
SOgGQ0p8+UM9HntjEw+FnNB6RJsNeZzhhVbnMJ1a9/pefEqa5VG2n2q4GNzSOk0mtGRQL0QXSE5r
Y8CqGDeBv81ibk7umrMgQc2KWoUqHAl9rgRWrmQhE14+//9OW7P9TVDaQo8vjqiJg3xmz25ynm3R
ELBbsBU5fjZLGj7mbpOfsnJZTxhlcO5ZBpxsLVQcAOawBZhGGB1WflCy/GnozROpsUDBjLi4lrYO
HosavDtmBfQCYXmXNsSkhKs2LsKjIK+aYupgWGVY/mRJ77VLdOfQFrbnnNKzuegbptHeP+T/Wukh
mlVbh9RWSc8qVrqi6aVXmNeDliuPZsAuMF6FdqGvJEqhxyP18PGHrUeM8aV7DqmMYSusEjxRr26i
AbdEdEqSq8YHyr9+VQdlIKGHLATL5UUTTqR4o2G7R/DzgLktUs2Nj355nqaUgNaxozLYZ67EqA0G
3WKkrxIwiuURg3iRazdasN6WZVy5YGHCMkkl2E2GClnee9GAIBrKO2KOzdArS0hCf9Sdo99Np3hr
7Nia6+sJpqO9CTscWqEkH7qXouiaGmLc2yNgOXhucglZNGSFyot7qI96W1HYvmTPlhPBJbvJXM2L
pGRKKiW6b9GpmRH0Q1EZ5i50fOrzZAzRR+hZRkyd/Ue5et9GDX0TbRXOdgIwMF5pccwVMKuyZvPD
/aJBFXE4oU1rec01BXy0Dzfm2sQywpMhgvHDc5f3Np/A1rx0QDB0xYnIO/Sop1CGyH+n0RJ9R5ff
htNmZV7+v4NY/gSWNMnzJnrHX+X0G/KmtqaN6LbFvdbTxrJ7aMggaLwBDZ3RIHyMk3ZCGLviJfD2
n2RARQcyucIomCj+I8hteZh19VopS0cF1lsArv0anDfVbkWp3ANxrb1U8BuiXYRA1NxUCXoFAq2t
6O8mG35pcsIKyGvH2D2riWcCR7KGOF5rY9l05TqGy0uneEWwbjoCa3zjM0C/PoKIsBdrYsR2lG+/
I+o+VIN0kmDvrpCuVrUPzI0LEoTYyteLwMSf219sDvufToiROEGwcfvbuTUamTcKb1KtHZuPpocs
UbcsXs2s9ky8zhZRHhbWV9yij/0EI+AnTH8MnsCx1cwR/7Dx7qDhUf4TA7GCSPJaSKvr6oQDJ1l8
ve9iqtLcELHHnKRwTdSMEljOOWX9OoXHEN5MeBLVEnTEGfMWXmPGmrPOnpjWY2RKsIOI+wNKOBIu
/WyyPIqqDrgDWADOZw8HezBnG0OBF60pFK+RsWERCnJ4FH9FYyHPQSDluuFTFvWqSn824VyfP6Fy
Xov7SYTxgq7L1ihrAmUU3/pZUbmhWo94ntpFXjLsZ00Jlp+pN0oqwDl+eSo1c1e8qH9XOarm7i1w
Mu8nkoO3Dog9uRy0A7GbyQvNOMh0GUf9Aw5+uvSsJSLII1+zEwpUIeQCjpZD72vksI6f6NUZyEfk
Qmk9BkP6iuADdR2A3UKDOISfToKpwepEJ7TzvVDg4h2j7oJR4NAKCtes016MK1RFDtfClYMurQfL
Z/eEPRCAdkbSHQWsvzrNFADXKnySj4zwuOpG5iBDFoNt4HYTJhrWj5JKM9fiFgNUraqWnGzSAtc7
+fQd1CQc95Zl4Vr+X9GaKPy6nOEiIV4MTTHBSQT81SBsHaAVEdSpzN/PFjDODsw32J+ZSuZoAuAx
rGn7HY6ZJfVRA9GxFDpjFj00zrdtmtIT2gwAGkoRxVfYCLF3dCnPk7QCisxIWasXPJ4YVxakMIet
WbhX2nri6/VONvbs2cGxWnpFB8aE31KvEGnxoAg7xbXZRieLJnCaVhqoRZV+5Ap3rkKXZgkrMgm2
VjybTdVglETshxP0+C+mOlOYwpIaaFywhxgCI5G+p/tL4tnn7ebr3GNklvTho0WJz+8AmABaeb0p
3YdNGLxFR4H0J6SAR2WNhBOAkVYbe398p21o8zqFKejColixALRLKibcXRkzVqccVL8HmK8DY44x
XJNnjB9eGmfcjWkUh44pAduGdA1rS78LmOp67tfbUUTgFYqFPD5KNb7eskv3Fk8ubc67+9jQZedo
nefQgfLDBiIz9lAXzjpWSdxmc7XSDeh8XPp0+XmxeGjSIz0qeY86cVWjnVO4YaP6bGi7ObmmESij
E1nNYNGAa6EdG5HI+d66BMWHqaM+db9JYUH+G5ZyXJnpVnqwjf56RCIpzMNHc3MQB0oCoaDMSHKe
Zy2C02nQvDHWfcij7755xephrNYJ82wrsOXzCNXMhhkcG7yYwkGLOzsg4cDZBdtNuaeGH5cNAAie
p9hM7NxzE0d2G0jKLTPARSr96JQ8BAUjsyFEV/ylRUCvwnBQPliwHlgz+gBbgBqLMR4v+YjHl3ED
D1IrrR75yAWGTjbHKyRZlsVwDVA7whXb0y4NDw8JyjqSwj/nfK3Z5FIdnPEcyISBawCyIG4sYgJF
mhP5BB98Q8JOybYvOdrvDRk08y/CM/G8ImlzYmRRAY3eNb5lAmUEP8Oh4j7p79Hewm39KN6nw7Z3
HSCIoqCEW8dVJXkbJrbR4sEUCgsrkLgESd4jZNNsb4e4kBXG0lj3RotytU+HZnuvOeQMc5TH4n05
4DtgNBv8SA+8g616htTSbNetYyKaV3DiRYb0WtPFDHNT7KL+4O9q8sj5rYtt8QRaZqdcKpjP8oT7
mZhgOj5olR+J0eMValM+Yp06HEXUp/9Am8PjE19OF5iqVNfAeVoZscOHkbBajlGEk+qhf0ZrE4/u
iMaj1L0ebETXiFoaRM51d2Ey7hsgo2jOrieu6I+o5DRCCNzcFDqwRfSn1afEiQYZPQ3GHXcaW96d
qHyEIL2VBWARRwrbu/YZ2OsQ4aYMZW63FqHgWahJLs0nuNHrRSC7F3U6wB99Uo5pTSpM+eGq6iMT
Tocj7L9bvekoMKBRwjke7L9b0K58qSrhS9KJwl71lwl1fLwVoS1ue0HChU/fr/KaA0amDHHj8i1r
KcY9nOu5ZdG6/uGTBCKa7gdYku3qa1Ccpx6NdyukytrkeQJ1pC2TfAmZiGKOAacN1j1tD0C2WMzj
0mF8HFGpqgJAmacIOliPv79Y6KTJf2GmeaOvGFpO9ynNcU+rHdv4MEKedCAakkwrYXiKOgxwJziy
cJ0q0QRPauAY6qBwHZuZUlmkgOxCFGGSl201S3D290/Zdtethr3lZs3cCfsL5hxCh8FF70MRCh3J
Yu8L9q0xBbMV3IpDMSKSml0p97GkteixqZtNkWHl1R01r0NND3W5FbKs91jqWkx0i5xBDcKCvjlr
F54aFLD3e/1X2DWxzbi/sawiDL8dJlHZ96eD1WySPV/ulWP6RjRckPlsyDMiD+3uY1sOxxoBPVs7
bTH8oasEucf1YrbsmOkMfOGLQ4d+5NSLdIqsXqbCFWg2jxh+6tVyqpaGWcD772whcqWrgDRDmnDU
edgIWfTGf0gLO5D6pHlxbkShyKSiIOPinvmF+88quGGNH0TIoaIN34SbbskCTgAXFhnw2C7rjczJ
d9mrnBDFKYw+syNFkTIPpexkAe7MzOYtx5xy9RvR1kRpPCGETTvyDvXOHB4GyEbiCunwn4gjdpqf
IEbwomhMSH6fo1Nrh9e/Mgl2wMnae++2mKRnoRdrq8b2o/Ew20Men10pGw4B8ilAO+OzsoXsZW+i
zmxZRGn07jmnwBzt25DkvMfYxUTNKjtincSrDFfeMKa70ANEJfbB6xHRBfzkHWVwS/ebXc0mQMVV
oEsKC7TQUdhhm/bWelVbeXp3FnMeFKo52AkY22jlAN1j5LAir90Cnf9buptythlvWu+623xMCbrP
4UzKe9CFYk7ib9Lr9c8NIzLR5neEy9+BsoNTcLPjoii4L3ORdcnaoz+RdMxnu5LXL0LV+7vr6KoY
DJaFVjWTThMbgsDg1s3nmk63tIf7sRW3xbFHtuhlOzGVdRgUEU35wt2ttyEz9QPRt5yIiCHUWPXj
EOfbnPsr3bDkZpLgNO67AIvvHot1g78lZqAbWRZ1IdpGs05ImQF5PcTrH1o226jaqWR3yWy6CnAV
vgL+tSHs4WRzejfFwMKxaFiTmrrFqZ7fnosNi5c7z7Dd+gVDK6rpTrZhhuJ95vFaA2tLa9Ou3bte
a0837q/WL8fbJGCKmr1lMT5crgWAgUWWDnxCjWri0pklGO7z6fU7VMdCyrTBVnYOVc1xDoqj7lFw
y0W3gYH+zOgu3Xx2ZgzP3Kl5cY10w18uKqrgV87NnGD/R09NYrGPz5EEHwolkwRG7eHuaXAcc50D
G/K7ZONbvZMpY3yqjLMAQ2G0J6wDmZflbsDXh3a7gbkMcgUjP/xsnnY7zadPMc5/977RN7dHFfL4
/KISrI05ctUvBMMZmpWt+ntMxWFyKdksw9SUc4jHvfwPaullU1gl4/jfqQifl/b4BQjAN4Tsvi0B
tniHZL54H50VPXgxHbwVGIFfulkd1E/G6tC1mNJLMVab/AGP3UWSz7pY2l3pNwnVX3fCASUohvkj
8PvVmIZqJ5RvaixKrNXtYVpn5J9PnC5y/ZUx9W8lmS9uQzFMOb7warYTcbeHBlnXEjOpJ6JgVYBz
2w+7oXGmoAEZQA/MzDZHZ797p+KC5CfJ6oDNdwlankYeSOlDi5lf5dvvxO6phaie6T7sYAInK7Lz
BtUUai0tTpO1QSTnD8IwzCVlnqXK20rrjm3cR41kT3KZvLAHzdUARa6Vq7SZYc99OP8+SuutXmqJ
3nNk8n2Riz4cIMOur4DUqgEYt25NCgUrYqXIamT7B7pPNDlwzC4Y7FZssdFdx3Mp8Zdpqism91oI
aKBiL3WEic/wX3G/gF9brT4GHSE3QbWruPL1ygaeJYhy1Vmx9/rbM/C6XrT+F/5hpKb808IKHP5R
CF2ls/L4olyLhx6oVeLqCxk3wPEQS1p2uW3RltTNrKE24TgdknciQSeTBn/v7rmQtSni54KTT3fL
WSI0pdYn7Pcm0p/s9jlh3q+iTOlmck5zmfGvhRo7l7upWzIx1BW60Gis5pGYtoCCSGergO8rcmft
8BYJqiWEhTFMy+0vkodBajiVVnS+oZdbUX5vCrO0KVwt108zdAa2IW/BE2ZrZ0FTOyjfKzc2her+
O2sIOja6jZfVDhHnl4be15jo5Ukis/fCSlXbeZoQPoAuUb7R7ozgOl8YkgBjxzmlAWYHfT4e6iwp
1gA3pBe7aARzsCfl8z0Kye+QIEdomWrFBacUMBfIhG+KRpd6C1oN+QueHvkxKM2Ops4qkVKY6AqD
v1c/qr5oXtj9+h4s6LODU7loBZmqqgwsCNiUlMF0SezC9mmeof798UDk7sK8AjR5zRggDVpn0jxl
6hj6VSqgvYbik7JhPiZRlWhopcIhB5eTD8x43AjJO9TrlQYd77zS1ludz8wiebms/oHSI1zvAe5o
/QT/b7+h8N+rT48nv9VNC10uYc+crtEHl7rMCJL0td8R+smAz/qEplBe5TUSX5NcF70FJoX8Pimp
+TUO9dx7nrzPvHO5lh5GJCjx04nw0cFuijh7dahCSBZhDvTsg8ebhRc3KL1lr5V/8nJ54M7kVEak
2kJSvYVTZTa8sc77xgWveGMi6VqR4Q3JxnO90feBUg4CZ4JBiczUaDcjRh54F4+aiUvj0h3+MOn+
dmaH4jQMescuXBZTjU5XgBc335j+9HTtibX9RmiAR2zZUxKvlZDYxMXrQCvPkm908v31jcwOQcoj
7gZPzuhelTyGaKcHoLDJipkWtvenJ0jnmdVClFoA77MUu6qd49Rl6NoOwrN+HA673tbMw/pB4jnd
hvFZVjQIPx2Nd8qD7/XvmAS3Iwy0SxRXXLT9Zuvbqui+FVMrt1qRekH1FYsSpZE7xwRAz5Rd02+n
5SAGvLAytyjqshGwEdB4eURc1T4Mp/ZaPILN3q1PrKEVNP7jj/o9vlxAVI6+mqCYIgLC+95D5WNI
DKOoJywofFuFOW/CvC2ixq/adzv1KRrWCoWZ7p1KlcAFmtbi6fELdvEfijIB9S4cCQ/UT5/2R1/J
kVzxze94HDOJdMa97ph8O3hClXv0+PZNw1srSUy5OJI92WPvK/zrFqfrz655kW0frKNo7r6CEJd2
5P8SMAQtsLHrw2Yl+o1FfRDUC441cPUsXoBQhMqJHabKZlsdEyhELA/YYg2GBE8aiR7/19nOkyFY
d0qf8vNJ6uGrkJS+NoYRRy6iusWZm95z+Ke3tGLK3zir2urPSNjCKYXPFJsiek4XKQWj47cYYV0P
gofehRfviUbsyR+Udi9oWo0QExCwmFa1EV8nn+6P2+x38ZMfA7pj7IlvyuMBksoW6HA49u0w2XzY
ThHWSOQDSc6l8bWInqlsp5YqpZho+Yu/Q4flkXg9P/5b7FlfF9UXXeZaEug4GKFqi13t+DqW15ZG
T64noyqNIhaRN2XpxppW2ZxJvo4puZuQhT8OgSggaMs5wMU0ofPiqTvyJTevKZ1Xf/9NluwLkS2K
4jaL2zJGY14Q4+b+SNxbp4uMYqiIpANcX4wwOI7WxFICqm+EFEuNiPm2kl0IMrvYSdwDAqz7gohg
qrjxlBq2Pz0uuysAVRUk4b8TTnteWTSQpWqFFT6gYa3Q5RSV0ssksxvlaaVd8RbEkNTO1/fqen32
1GrMNSSSqahyvqzuiDOgh9l+Aub/4dCiXPmlO+NkmwyOhmyUusFiKl932CSf7dcX7u9Ijhrr6a7h
5mboGbq0lcfMEDmIzy9xVixwEbX8Mssz7q/7O52DHhQ2Ne3NnC4xVQUTkr/7RSSoIjyBJ4+HCTyP
ysU/TgD3ifMaBMmtiX9kGq9kliIC36L+3Zxi3LeCDA0RG/G9/87ZP8CG7f7oi8UXQ2VabwJfDn9D
XR1szqN829DOASdR+YHzb/nz6Kgq82Axsqf4iLkbNLrDPvWDcE8x0sjNbafraQj9Xj4D2iLCD3u5
2WGPG53udZk4lJ6jQxlOmgOLtO9MRrvW64c+2oHiFi+42CDtnMHutYVJ9fCRrrlLPeKW29vzg854
CafiiimnCZyN8I4HXOG8+nFhXzUlMCISMboa+itBG7PENMMSuXSLOsCnC8kmFbdBA33VAigmOt0R
UV4W7pYyWvAikHSOf3DC9ftNmQEY7CmlfTWb0tGy7sl931qZT7st0HZXNnV5yKwm+VTeIMTr40He
aBTEGc20gcMcyh9bc0SwVnZeFifbwfMOF/UuC1BinR73qNDDk3BgIVka46LQo1L1oSyuTYyfdFyi
qpXpwKjqqdFRHqZmeUQh5JxV79Zib2hYMEuyB/G/QWG9JvetXZsfD9xOBkY5wIUtpTvopwcRD1jY
KZkRko4OEp9jiQNl5BdohAort8jkv2gigNQcNCazmc0VxAifSiRuLpCepaekdHDn7q+oTh+hUzRS
n4AhNY48ocxeUlsN9ThQiPWREsC5I0A/8AAFHekjjsfmAsL7sACf8Y6WmMntEPWQF/60pCkCnAjB
9W2k8fy27Elo/cKb3PyRnKIc2bUbCOZZX6KYPTIxGTLxdNfSeL7yUy4i64ELndNwh1NzF/C6/g4S
ZBYG0zlEEuApfeOLB/1HLV5HCcaDL2FJhjEBDb2DHg3ZiBClTCCrDFD1B5x7k+AaHKFymx1wJ9ix
4O3nTIky2U8vGbUkmrzfB2zbDybamPQQnsF/0SeeKP4wmUPjfo0U4BOkOP2/d1iKdpN5jMzbqb/q
HH2TIuxMi0KrD3Hcfmr5ODH5frJK705FE6a95nft2XCZNtiIoorerMHvGauoKQEZUj+TgC3VLdkg
i7JbUKyrHHtKw3o0Srs+xySJzZJlVHvZ+aRKN4wsEw5pg4TZ8wcUkawJ13jE0WfHINrBUjAJ+ImB
iQl6aKG10Em6QqpimPP51b75YW+B/b7Zye89Rm1deW+WrcoJmbaZ1N6uuSJ2JOg3VUIaEqd/az24
xwEDvABMqIqHtSq9u/lKbeXLjvfD+v+0OPPkNA5uFQEyC+8pjQt1vw4OVLunxBaPm/2opEOvp/9r
LSy2elt03FrMNj6eWv+ysS6xHUEEZBUFaxaUc3nsijhSlRAPZ/BKhxIBjVKZ55POu9dl0r+tRMdg
Gh3dc1qpOxlg2lWaP6BN+owMqdrs/RFkk3vebluRQj+/9dprsiP/d3a8p4esbK+YG5kxwoQtJorS
3umwag2f6WHp108XrEtZ7fffopKY+vFfl5JvEHPGEqAtxJl7g3sKOx7SlhtBehiGhJIP9mzy0oWH
2Yklm+JJEhdhiYHvYT1smXxmilA+PYoWLzh/aBHMoR6fL8dW/+Dqlq9bjTTcdbluleqCqIgyUWqN
N6L5WdgVjxxh9Ie/VhIvyjfiSbPnhyukT8CoKKRVEimJ7c/H0cTrc+gTtWl9bmMYI0Cp/KPRLX1B
wthQacJS7bV2xqyI+3lU1fiUo41j+X/GfolTDHN9rL0tBKqNyIsN/35CViTWESExXg40SKdN+YHl
GIqR//KCdOTi4KSBfGTm8t2PyXyuohhuSelvns2qJiA/63MgirO0Yo2/6fhmiGrsLTUovFAt+fKD
zan6ATnxxn5eiN1bdvu1Kuy3Q4dIs0wJonmxh6miycgGUHmjXv+wPpz22ALZUREfGQpzguTMg0Al
P/ZldG5vdzRSvLbLDw6CwYIIyZTQYz2Hua9kV3QPDJK+FfEMeSElby+bvV0NqVckFyS08cAo+Q2L
4xw6JAKRnJSorLcMrv8431VNDwzC743ElmYcm52ckDcb3tr2w2cIKgNKhgRwwiXa14OzPSBevg/M
74+C2r87UZs/YOYkHmG6bg4wLqOuAws4CG93xDBbswB6JomHYi+FZDn6Gdrm30E6qSe3iizCr7BO
irVFj10zi2zpVRdageYBfRwxi38koy61DFsWJ+ECO+esR64Nmx3W2p+VaZqxDWiF5MqFsTxeDjbV
zgFUDpIZZMgmDXYNkEBVnqFAelkdpUyNpDYwzozN1CPtDOZbytX/PBLTnFR2J2rbGvB1OKGseZb7
lVMyr0kqZQBaOL4l8nyyrmQmSTCGirUA/MiFPsnnorWmti5HZIn1kXSdoN55NnnbB1vMdrzfC/g7
MnJ0y19qbkkdxdyje8Ny6eaWBtr8LRQ/SYo3VvLkwTAHdO8OOrVVe1gFkas8gp7V0IjMn32ESqn1
YENYsGmJPK6ewPav7nVNQ7e5ASBeWmfcQ/LEulhZT/bN4rCZMW8DjumTyHHih/EbHfCp2D/7aRde
0DOjkbTYIQePlm5y0ZoZlFTOK+Vb1BNN2vWM3B+sD3l9/XZFvYXKgfi8zg8O3FGMoB/JyhuyPeNp
Q1FdnLBkFkRBRVw/0cX3Eh+tnCOtUzmfhCy3jYwGY2RV0nVzh9lovJGejuonnnhhLnfsHl/PkhkU
u+XQ0o/npM4k4U4kRsN5oHi1ulJlaN2cBmJmTu7OML0Fj4+OE6R1tdXjqO/0X9iz1a+xNDO0gFK8
ypOYuEKXesqv19eFwqDI/toEBT1j1Sw0ZLHNtAkYSqxPzhRG/eB9EIrG8KOeLF3P3ttjSf5TjnnK
KfVOSBXZcPMPe0OeW33yT6Hcv5vYUpofemvD4xc24CrNz1lmzYjgkYOkmI7O2lPyaJ7N89xy5zvY
gDMdyWErR91DvL0IDaIxdtB5XuC/5WLxa9pJDTm+6XD1C34cnBuyyKJR5OAu2n/Ij0uESPpjNIfv
5aN5VX6hAhfrVdyIZ7bDIPeb0hI9nQ31wzujyi2YI9aO6tR0OI34CGRPyrEwsztmWv8M+D6YC011
KKH/HAijI/6U5TwHke2FDmi83GFEEoDZgyyiCnHkj58tRaxsbNiqfXlh4+fIQlQplB+7n0h1dXUu
5KHK6RKMP52P5aTEInZCbRMhDAhF9nI91WFlObmzGHQ4Xa+3gyDcQQlCwmR2XqznncRR85Imhk7A
h7ZURWckVga8BuD9j7RP85qH49pQUMiB4OxdclP9CtZa+w/b3/YpD2EEF5IEVHdYUryAqHIIO/y3
FsD98DHKOQc6/RRPw8fItYAgrXKi5Ze8YAuEL3RZ5G4CC/vxmROMVCpl2XeXccLq5GGA/tw1KDSl
Ri6mn0RENM9weIfcIFilp+Rtttuy2YWBFo9qqzXf2otuexSi7kKL1tWJjIKn+8yBh1/RkhMjRTM2
lfUiSeubW3hOziO85PHJiK45kAjQl3S3dCZFNb/DNt6TMdP0Vr2eBKt+Uhw3YaChfJ75lMNoCUvn
cNeiYbcLEU7i3P4ZE4eyEKEAGFhupl0bPw54xXcFH0i4j1ATqI6nfwDIok7f2adu2y+QXOApQg79
NUoGBXzK/ZUyMhk45f5K6u9pqzhu3q7tUCnEYixJxfOiwQKtrq+xyrql7yWfiIySbaJXHN1rX99L
NM57SUv4XUGgjUQKfjABjB75L1MDsfMgHKhs0m9QXtPSKb9fSncOr1coczYETI1fZqmYJkxNPMF7
B8JFF4Izag/lHaDnFlvdtQ39jxNWdQ1dEdFLwMuxxRLgYzl7xy7O2uiDKSdSwsvPN8jmtRZ7FTNl
BYLpe0EZkyrAhEioE6yIlqS4fBvMMK7Y4RaHe6bjesLCVAVBx240pZQrD0ACtCL3B1j+bZnj7Irw
8z7i5qQa+bKqBXeWWIE+wp2slAUMSH8nflaZicz+VIOfZKEDlRze+NQaLCaWthA+Ms25d2e2174W
hWBokuCkvMklmxgDo4bNL9T1pYcSAzPvv4MVSlUS7mrHXO2CkajuRsCQpozudRAmOCO78WqN/9Ad
dHOwCIQPh7OQLZJTy0q+QMfV9IriVMUlIlGQdinA7x4XhuZazzy1IMeRCshd/pPigVG5biMclJrC
WLL7/iLCYmNjbz4DfndYHSMdlFBHcaR5bs39Rr71iwuWqIgR5ODFfHIm/8kP1vt41qGvMHXoYaPi
PIETAoDbrU07GpO0LRRhIvqvc5Yns5/7ZPNVmQ0uPkkw6/E7NYoQwZ8sn0mfYT4n37wRCQVPKDyn
Ug1G5qKnr9t+Y/KkZKUBcEVkbr7bwBdR4ZORhaQBj+uawgYRY353JVUfKQgs+puXT9h3rQs+Bnyv
DKRavFtgqg+MEz9wsE0R46RdIP0m/Bc4/T0LFyQBIRntU25Yl9xO/qseyhsNAUokrrVifEuKTord
vlMjt63rmpEw0s+gesM76xIEU517edYNbSchZyTFVebBdF7EdjNG5g3X46qRvfuF7uXv6+aAfmrk
GqEfgFw2r/vL10wNj3eWa+GxoXz2z5DDVwlIptM67eCpVb+EmAXI3NqCclcJtSEnejAnjN4l7riL
4zovGYqmfFsAXFdYrUO3Mj+o+AvU4kIIwa55Xg3O8JqtZr7+qXapPOR3tVPD/7wDbYSQ2u45fLfl
dzsgyVdnfknuAnIIr9RVBvUwvyXDDv8tt1OuT0/Xu5yaqyEmSv3+O42L1SglfGYYZSTAjRl9W8FZ
nN+3iK14BflKJ2pC7tg+p4fHdA+oBhu6+/K+hgjyshnZTeRR6kiDlJHcbgIAhT3ZuPMxOSePW08n
45Nui5r3L5axl37LkZLw5glIKSfqaSFmYM5IKe342sDEsp1UANqhWnkIw4SWydUJAhTUjXIhud+k
LA3uyLQSvJhQ+8IXxUDNAnjbqiT9saRIdWJiBK/Cwklr7YFhBtOxCrWqC11yka6lu5lUl2RJ6ZmU
sfBSEn33z0RWyFNWIHasLdRkoVhFZrj7wGgfiy7Bo8wKRdUtZKGM1kfhpSHp+djyakRGTHIw71H5
6wVoq8jMrweWoCKk9R6znVC+eIeGmzOyZS0IwcfLg+046sFZyK2USEHqNdamY28L9hvWl5YVuwkI
2EKtLaPm5ct/3LajXB8movhRD2FWiRI5qYUlqK2KKaJKhxa/qobZKN7U9IMROvGRIXMTozS4XLKl
+NIG79s+LzD9VSAC3hS0U+8bsIyWynIqOzcmD69DBKO5+YqD1BDdb/okt3DwrddCe7AY4or29FYj
mDyly8y5hX/MsIGYe0ERICMQUvYOJiCoaSOwwxlSdkWGX4+SQxrS/GD4LjXks6U86mc4sKv/dIiv
uD3tzSC81zUE2IZPatlwNoYpIqOws6dpXv1rrESM4p1wKok0aBmO5fMQD3EeKn0OL1vHRo/6pjH3
ydPeT8vjBAXwQfvkn3MC1y6i3zJlWdzsDZqW7RzwTzVkYUWD7jH2tekR+eH4hfZNU4h0kd7+P+rh
jXxKiDLBHtKn+bVpL2r7lBF5eqAshRNpqcJ+0EllzRssuhHIYWMmRcOrbtgnofhEUxE26RhQ0zsT
dYumNLVg0kIEzF2dgTJV0BAu8Rm78fzXYPwwPh45YeC/0fJBDvZLEPwZVAZuX5sN13tQ5xNAauUa
C/rAo5REunKoDRfCPRXs27MzCG84aykdWkjIDqjSz8QBQ456Ftu76zEXiwy9Z4GqOWNCOCLBdvig
6eJo6SWOrUqP7eGaNIZFo8shHspsHWmsG+0LhOlONajvAdZgmVOfJfOZdbTQIL9+O9iqUDFwDHni
K7DGeu54Jqi4sDjzfhVFoer6CrHfuzKixo75xALKk1sim988+1+JReJ7sRArPFDkuFlK00UeBGXt
g27PGuzvCyKG2153e0rak5N4Yo5gDj7VXJrvH3dlmZZao+ee+BEdwe1x7TOSpZ/aDg6ZUrD2vr2y
X3AaUZ8ex0SPbBkTxqRvqjXSePJ4m8ftIfVzBiRrNj9pJj3auZblatJTvH5sH7E7cOhnQa/oF3/q
ZGjYqJiJwhtRfSq7ZTWVcGfWHiVKqFT+bIkdCDdlB4dEWWsh1Y7S6IyT2ibiF0JxrMI4gGpFwWtm
Z0QG+6jgJvjJqB5Dl+/sWifC8ioM0YEZVc8FGGFhdOpMwOqcGpYfaZ/jHxB+ZQGQPhuXblEMC0V4
3y6qOz4QlFOBL/jWc7kUudpOy8/4XpXZ6PqRYC9j6KaYh+QlnjIqMoeCBAZKGo2gM5hDa1J9UFma
n3QS0Gc2R+pds1EqwbnoILFdqlXBIRitOZvHbZg6wOvuRlnhuLAqDeKlyvdWYYSt1zT5k+8UP5Eq
UAfyS2LUY2f/NSHfT/MlYngt+yslC8N5Ej6Aax3YIuDW3myO7CVlPnd54vJgedy9aAWTE87Fc0v0
VaZlXY6vC5PlrL+fRwQ3s/XdBb1WrahuVXLdSrE2GDsri608523xdaZizN4qc3BtGmuALKLHGgTt
tDzHWIi/Vo+t5qLhRbCZOW5h8mtwpD2Dq1FeRepX7HWeYcDsXpXoMY4gmWyXpylu2PvkYvSZ93Ms
7Gz3ycQJLN+ajgI+OE75ZSMnURbIiSJwegbfsslZ5Ia2pYN4iBOeh78JIRG1CIsapdP2ovQbpS6V
YVo4Uff3Dus7rcG320HQ8S4+wyDflOQWJbGRIhsyCTj6VlSE1cDPZdNtF76EQzaLgZ0SB0J1ACEu
OyxDNPyrqKk8vhQGL35pkgked1xLVeSo+etVOrsBt5P2AGmfAbwp7KA6b+x2Aznh333SUNEYLOvW
O1X1XnTSvbDvWoJA//C3UkGtNzJMKB98qQ72mkLQf6+5W2HsziQfs219WxaCKI7uzCqjIgZRZE56
rMaulbZ44QT81gaDh9CuOyFvvYKp0gw8QQa9YFVRphzMSvf+3oZyQPDn5p+TvfH+6Qtcqixj+z1h
rjoq/zob7ngZiVAqz+vlX8gHJsvrG7IMPiyWJi2qzKAUOo2yBkjhlbypqazi9i2tf1XOvw15nNE1
LP6bJgiTJNRU/ob78fyBB+RBSNSKIhttagyLKHZ76UJnuy9VPh9ZUl4h0x4xpSgB/tdtHQ7im2fV
WEPKpXsOI95Gi18Lav1PjZx4juk2Ws9Tdb+QMfS4TLuyHOh9b1kgprPneA9K7Jpj1VKVCTzKEkMO
gBU/vsn12+fR9woBgpkAd20L5gxQxVqnwpzzbC3I7NFNrQZ+kBqcGongkEygGApTgmucUvMFitIv
b7+OAuxUrcVaD//nYSR7uYtPVMHpo5y/cXX5HifHpyEUN0QGZRchDHUt6ETHHN2HsVYfhG6w2uqK
iHlHj5Xv/Qasv9gALYFK/msE8m6J16Hy9pArUyBBjx4meQwNqWuCCsMhvvZg40/yv79v9Wyp56/u
+3XycVPVCIL7XFdbYrf/G21dPl97IdMtfBwLdnHTfOKgn6oS1evmHBrxYCTeuWrTe/YpRZRc99NP
NZXsUHgzb+OAYQyWvE1a4pHkO1Fj++WR9bdYbc+Ys+VllGM5QOyYpt834IL+Jpnz8MZ7d+6fDFmJ
ii2AXIPLHxJbW3SQc+6rOZEzBAXzghRe5rK8BpJiXaw9BGHjEQLNPMPukpHw59VEp+8lS1yXR8Nx
14rZR+VIwa358gWxV1b+9MjLVw4LEB/CXn2VaMOgshpZ+hK7WHFE2nmekUzwXoGD3JFxCEpgernH
GdaSRjuhq6NOsVZUFaIwOu4ginvXjgi4NgM+1xwp1rR17EymJsXMsiLIQ5bmpF9RDXfj3SvYmiV0
EXLVO9s0gGX/CWc7YomgJGsBLFCMkMui1bRZMs8UHex+q730uORVdxhq0G9xViarfQ3Qxda2Cqbg
0JECI+hGCdiG01D+yVJmUllVtzXtL/KWJapQN0Z/p3e9Jn7NOFS2rk6xfxb7UJ7NJSBLUv1SWTwS
aBYxbQsqIzgpMpPNMA8Sk/p3LLNMt2XQ9gtFwE46NgH02Yq+7MgRDDlcPHybO979EZ30zTYkDPHv
x0nrCQxDzOOAwQvh04edB7TGRH4i/Rmq9F2n/iapgccH3/rUaw9TDP1Npt+aZze8/f1JB/N/J/q5
3WgtRTU9aPRKUPGbZlEHApJBLUAYMVazlA9QGOi5g5YNmSM/03gW4e+APig9dxqlt8etSsRWXaGe
0kaUPMS3QKMxOzmTK5U3vgI2A7i3Lr1Tb/ajNGC7+PUd3UtoyTSaO+Z8mAfbagSsm1RQ6rHj05T3
5VgbU20RD9qHtTstahFFHNqIvIDgVg2wkyJswcJuznVQu09OsMOZgYHMlRwgOsmzJ6oirOLoxhI5
mRZYNu4nA4kd7Iolj4l5Au4A8oJ3JrHL6/lbVXbe43b45nmAQWlaieeDq6vjG1D/k9PPlOaCGk1C
gITWF7/lb/9C9EqqR0oe9Et8avDBWaH90MtN6gwCxzfnVM3l/cu2K7zgycrtcUgbOCVURSlzUVtq
VznHiGCgiLF6rF790DP9wIlttb1EhEWEJKTm78eGiY05a6Yu+ZmnvCsUQw0v4F3kx+H96OIHVXVz
VkWOqEo+4PWTXEjUiUXBpUZ28sVnGa8ddoP0jS5MFxUg5nArM3YmIZCw8Q/id6tzkl6utAIrRxll
ywYDCVN8qcpgymUeXqG9X+0x7cE1i5jqmBNtW3kT8adsB++niNmJK3MQql1yYzV4S91IskD3g4PV
3BVK2Gokd28er51jmPj2P53e0cblSFWfVE0/nwhbY3LHZXiN/sK3MRTVxNuunqc2TtvlhtDIyxdX
zoOCDshdzvaPawDLz9GVQDSeKY6GJDTkM/xNXrtIA2ha1cun+6UO/uFsroGdXHmWEYBDCMCpgUcr
N73BbindCD2wg5EITgQnR5XYTnDKtBxoRmoMnkVT7KOxZi5dezswR0+399ho8BdzA/K0B84opoqO
FToXybKkAqE6mO9MpZt5FIsZ292vTLAmu6UDrw7/NXf4mun7PGJsR68cV510ZDr8sNdQu/0lSL1B
f7P6yRJTNlH+JwH9DzGvAsLLbX1IWmmV7CIED/0OkDTt7TjQf04F81BoI1BKQm9GuvJ31XxERcca
iOSOdAEonRlhhZcI4w9J0kdcVRedm70A1x4sZSrOOsJM6rOyoneqrdFfuby+hi5wOP1ZNEnmBgey
RPIrb2JnBXpwX2HW3cT5Q9QE26A9FzRDPOdLFG10PWHhJXrIlEa++2cGNc5irCrSxD6c/wl8/jgX
gKEH7zUCWyXg2WZp3aScFynWxLLpM4mPuJsm2rYzj3FbJ6GV2YZHaesanqOYUIos2Cr46Ar5zax6
c7OYT2QqjxrNcuM8VpUkitpYgq5uMWz9EZAF+PXt2COWydYXxm31o9GNzEDLG46cTw80B6WJCGfy
SMEVTZSYShgQidxejbrZiV+QZJNVXMjEckNt/o3+mCNulyUOzWlIUPcpCstJ0iIsibkGtRVJEUdc
cr3p92DBcvEeQCFbR8PQPTEz7A1F3bPuEq9MvArX0JagU0GhmKwnw583AE0T+riUAsuPrk1VaRTO
pEY8ALtt3VN9zuN1JYstXKDLCIxK3QLcyP+YX86muGR8EaIUm3S3s4k/p0k24DI8VqRfJfnIrH+T
UMonmyIqisvtm+4l+IXTNebC34llkbkJ8BRaCNup/szIrWg1xNqjByHveuYLwNnH7eS3lbZzPS0a
gw0Nqw4QL+HhJGASY/UeRVg1txQ7EPI2D5Grrni1vxTxjNWgnvJGrnVm09rv5MgivXsqxui1eIb/
5Ffqv2bu8iIV6J/4JcgzbJnrBDYNKmbOPNMbUVVbFDZqiz4HOYWTFRoT5QoBm3mN3a5rJzsZsXHD
TufAyTh0UhmgyIswMYnVYmigSvNC2GZupYl9LNCJPKCJzDz1SHNpaTTp1RDTDAvV6PmFrp/fSq4R
OFkJyRAMzh3NklUlWdZ2LvrdtKYNzaEHzteBXHvDDrtxr2TR3ev2h/JVBcubIwxS4pB/O0FDPSvd
WCDTZaKrVhG88uBeojVL8eaoZSGCn65EBM9Dj85HW5vFkdpi/VUOgz2NytMNZzrKoUzExPgi7W4E
0Gbsrj+WPHECNB+s7xUKCa39LOut43x1fGXOmy/OxJ3TxZ1LW+QXkzhvPqei4jCLurAq492UjicY
8xPWK639Atk6F73L9UOufgw9V2Cl2Ky6+kIY5kY3/TFcB8gzPg6GdnG12XowvARDZhHpD5XIvT9+
++VJYwQTvlxpiUmOdjpZu8DHlFJYafRu1I+PjneQlwvSOIXuCSOuOkuMiyqpN7knXmotEQudC+CY
I+6B5RA2M0ZPDOsVFYuhykC4NxT4EAt1A7Amw0+2p4b12c5lmunmLPmY5BFRwv6AXM3t9cK0VdTD
sHWHacUgb0kggIqTQoXmGhAbkuVo5wtUEUyokJp1HeTaeC/kqI57lHvPF3IOsjtVdjfH+zYZirqa
/kjcBWeqdsX6X3EICUmKrhKjm2FvdhjxD+QV+spem0W6T807WPsPi7qZT0CFh5zNls3uOt8nT+iG
uLSlOmokkBzyuNAqGN7tYac9A2TVfghuAcpnh1XN2WURciH2w5WOSkfSoYyeDstgGq3Gjz48lXZ+
YfgayZGMnSiD6OfGL5wFgLO7q8mplDqURt49ENLJJ7vT0HpUrFd/IBftsjx70rrHktsO0PSjHf0F
1TyNjdhGRraBPAlww4e17fCdV/yKJa0IOa4nyEEGQglLj9tjCRVrd3S9Y3lOQe/+WE+dYEHqhzpM
OdiF0dGlAUkb3jwEpHCSSi/6b0yeUQo/Unf39nhmJx9RLWTqcpSeRlsnEi7zDfYWi55VV5mOGWdM
hQisfer0QITBClRWKU45bDOsLFRFP4JtD3MY8ADp2nRt1bDt+TP695OPW0AKwIRRRAscCYmcFzl3
HtaVEeWE8PyPed15K6YohpiDxBl8UB+Ee6LO9vPUpxlEsk0h2OsuW4rAkpXQT+t996961Bl5youG
WBembemEeCHxds297L3WuGNMUmmZPYFAUmyjIeV5FW7vMp9Y968jzzBlYtd7MENVlD2fVl0M4Kfo
1xU0rhV3oGn3eKhHrRnG2nH/7D8/eEEY4D+FZ5US0cyf0Ggu289yzevGVSxRe1tnvvyAW/Tu2fpy
MkAvwaAnH3K7QXPx7aDGsJLEGIfbowbsC4c6Uwbd9KsNm2By2Ai5t/mEGdsU4lQEVUX5p5auj0Mt
dfl3CnS3+pc/0wTjByMzSQwwC8xKtIXwNQtTbBlgpzIgp2YcqkeJ2kTOpyL0/M7LCCCb64SelpLF
tViI0LmqnRvSm5G3fSgFo/5AigvAiKERCe1urz2NFbwf+rm+V6eNdGpux6KFxTV5ss+V9jqi2LYf
YSd+irw6Ys6wAL8lIr/XgyfAI1EDH4lJlOPLE2omtNws/7OF5e+ro60SN2tyrF16RNbVL4SuVrrP
JGOmacAMSu1kkzPSh/vIgZNS2jPHj33nsYZkBv1ES8okx88zEZV9Jht4qikAcIERBYwMIGDxzuXh
E4jygEefKFuNECvEmMH0g7gQBMhWu+d4TuVoUdYxtVFXP+fq79gRRIyLEIMx1hrsBkO3FpbuZw2x
uAKfa4w3VMYDgLgfHiET7BIR6tpH1z/AkR//D22Jif0O3UDTlrSosBEo/PiCRZnSGrlAmzR8ET+a
AJyKndTzmMV7HR7EhZaRaK1IQXM9olj0H19fCye/GHuLxi2FXYsXXSMFa5thNJ2o3mCuwlRWD6p5
MgFWKN6tIT2xK69jKUM61Ea5zcKxDBdlkEqqu7/4oiwv/zONGK2MQVr1+RO/Ld3KjaOQEUmfqwAb
LYHl/Cn0l3pPt+kHfcKbVlShvGNIcxGggShr7dj6VODb7xI5ipY95+mkqYQku6nPS+FIq61tc/9t
3tCipuMaMP0Se2RkKpi9BSAx4xYeRkyAsP0vxKDBMLoAyg5AWJ9OWfqUh8AIdScKtaKmvKuzYN1Q
5ObO+UVif3gXHveVqw6lv+MN/OA7xrvL3TeAJFodee/LDPmSFJOdBu8S9+HwlyYIcX+QErfbHhDw
djRELC7M5JPssx14TUJSMzm6cmqF8Ep5g7Tmdx7+Eo0VK0ZOlMRVS2AM67hAEqwANwfYwTrUfdmu
sCDTLaX9WLIV7ZwzkuaUxDOcIqLQyZZV/N6m/COjPjfqulzi3HnpdFAjVn7KEqghENUcECVtjDXZ
yJzp+0mPjZ1zH3yyD238DBZ0XyPmScZE6T/SN9IE6QkQ0AfLY4zO/JQsOa/ZVrCrLukSUWJ+BCo9
L1ARt8b2PKwe4MUaJwdeDMBQXDreHrBVjSWRGvRRXRUGVgZJmtaOQOAV+rMiMA7uxltB7SwqZMDR
EAPqmNhL+QVVYN6ajc9sTMRV1URoJhk2uGy+/TeNTXUlt5w1YHvclPSFXph3heHOcY1FIjVPDQKh
rwVIKdqNNw52xDFx8Td2XOB+h2x8KA7X2qAagdMYEJTNlmFWpvZuO+b572ujUZblJSb2vA38GmrX
Vi82ToccF+hozWbueJR7ndK6RDNZ2o1QZ+GCwQGiXQ/or18jexUp9O/yiOy+o/36bVdCv4u6Na77
KOoR9/cU7zmf7dwsg3flu2HHk2SkU3mjkJcJA899Em1YjvoJSG/Q4zy33sGVt+IyrWo5KWWzaGaT
22xSfpLz6m9bAaP3Cl7Cxh9ZwrO+zMx5Bg6IQpU258/y/9mMSHJq3i+srXWizdECbwyilL6fVrx9
5SpUQy4x7CBILQsr2DGQekXKMr+OBCs7AB6KaNt8GaqQp844M3v4+BfxdMtivVk0o0N940pnzUSe
vRHJxOQ7Sn/9Qga+XLtcBAF0kxVQT09XClFliTr9rNUTZ/d/HSrEqeKa7x6xPxsFQzqDMi1qheqK
aFPGT0t+2mylYpemjpvnLLRzP33dPK1ZCtRPyysjlhoeZAgf8+xpjAqXX4qdujbR4dugIW5wRkKX
LdIV1mvR9V9ecvY7aFTvH/gAQ8QgmsUESFOSrIuA8xS3kOwXfzADpvK0rggXzhGJxdHLESPppxSN
NX+9+kudoN3h/pGKWZmYxDkIFvFRLaiojVIvf/a09H9X/0dbOr7dJRFjLJ37e0tKXDSGBP04JQlB
OFISTBI+6RcFuu8K0rCI66EoNAMhdGw1D2EIr0zj5+tjDKYYmU2zW2vI366y85dw/zNSTfoZXWVQ
wHqSMFc0cRqqhl0F0ZltapTUl3ST5gAfQFeA4vZ7uiGmg/r4Li8oiE6SU56QqJ02hxap45Gr0BR8
SZFSbITZ1owNHCtJjLxnpLuOk+ex8ZwyotLspgS83PKDr6A3sJZPFv0SJB7zZat0XpWng3PWDAum
+ag6DQQkfheEDR/uIIVyzG3x0rAwO5V9euzVqL/zrwjugDiNxjFY0qGuhaOCd1AuThozrVzD8/+f
UcSioxIUFlgvZOzs5r4cL+inkzAil/DicsxaAhinvjzFN4MupJ4EsXdGidCFIeTRhE2SJvDmCW0r
9G7YIbvz4NJBtcEi0AbqTdulVOjetf+e9FkZrI+lkERLc62GBoKA0Mmkzl2kwLp+WskAfHzjGZoe
0e74UmyvZc/bxo8aSlIZgYNW0ZVHtw1mu1hRP3nFCD8L57E/Obz61JJLcaYVEF2I97SI/z0HteGV
cJH8EPhMU0pDVBsbRhM9I0OIXZUtzWud7PBk/2gkhcQCvQPvRq95VqCwXJMUGjJSYiZAppUzCRqN
FtQ0QXBH9rZde8qdR06wlGXk2D8GbFfsjQ3Ky/4Ew8ag9UY2jbEkbGP315SUZ1ctpHTLSg/hWuDI
Z7TrKA26CHHHofvjhteZr07wtDqwzdmvJ7lc1/oP2+Wrk2At+SlS0nQe9ZKYUsrDrWM2DpPrYICQ
+9BePD1vERZSYUT0nR9zZhb8V/AJHi3XBqrsd8C/KOxkrtJ6Ia7qlge1NS4caaoh8VDOfVcCJPcp
maT+JbOAcZbewxBKkVhq/htoCudPkiE9rbrsWJ7o3pI2QkJSgfUP/4z73Pr6sQVNlPc2E8/4WYKM
dXXBMX27Z/NbSnwhrgjicoIuBdofnGGVX1Y8fa2FluT3Bgm2T7rWZUCfbu7yhwudPaB/jyLLLcDf
LP1kkj4KkN+lazgVLYfD1bS9i9cKm5+chTJe5qrSb/NKuFHOhukNp8RVhJYTcAYZGdtCVJh5xQ1Y
R3v8b039DE7Dh5vIAHJRcJ+X3kTzFCgm49nPwXepOuER6OWJFt8yBaDlf93M+9m8oZyUfG4+5Ysb
hPsKoHfe/88+5kNwqMtBVTj688q9m7x1PyGTc9wE1mJQVxxs+cu4GAGPfEOrAvKOF935d50Yc5QV
bDWhjYFgR6qWllYPu8VRO/9M/4i7kOrqtPCP8DKcfwbKn86qvvhpllQVBvuUuAtnm2I90Cpa0ZtD
aolxm3MVGXmBNTd1u/cSGLLW/mpcglh/KoRwHVgJV2I5zMOahvzQ3MEjTItsH5OGX1AWc9uFtZ+a
pCdKKWboOIWsoM224BV6kCVwrGPVkRgtZLej9Du4UoAiVzJQGLFXVxX3YQYVr/YOz+ny8PNL38gx
W9jAB+CT8o9rd+IYA20Ex3X50fJeRYttynPIUuz7qSj9qjCHz5ADjD/oQjiDvxxveTuRWJh+Og76
dujQ72ed3NYEr3jTCuy6sXMuxRCzj8nbVk+yCfm+rdQC9KidgV4/0EjLIuO64kXunNlfSfJe7NjW
ASifq+EfPjf4mLGRX/M0wJJNUVaJWiG4FMbRd7BxYM6wPu+XIXaorF7f1w1PDmnUTLMvH9EYZaVy
+CKQFJ3BveSPwCpNY/CKmpW3lFe6VV1vHsbAYyT0SrY6qzdV3kZbllBQsljxWnCEsMNfvZebDlZv
H1IgeCGlu8uSw3eeIjvC/JF5ERqKiVlafpGGMnw8oWbSY/U2WZNbx7njIXxGRoDagYDUAYvXdTm1
/kvsu8U/xVDH/BaiKGkMn+tJgIx+EQPBPyqZQlxjZ9hauY49tTm6/3Pmndo1zpM9ysJJ05AsrNNB
sgKJsHP7RphaTxMzVzJQbjflUzx0YJCK+b0fdzBM4XbNubG2MVLKiVjaUy1FoVVZQqyYTT9cXGzM
Xdxv6gsB3aloGfPi13xeR26UZekTnUim2AjIVAzQCtzZC+bPB3kVrXMZwsc7/JupXuxX54lM/ATH
x+F6CCsBS2bh1As1UzO7Mdbma3+lECsHFNxQOEw2G8CZMnxzKtQS8cKO/3EoMLlefiPz9W/dJiOl
XQitHpWIPkfZm0OF3oeMdsJchl4tk/UFqmw7FyqE7ds9nPp3ITfDfojp8sBpwKWJZaEJvnGAQ1LD
R7Jj3RHBWe2lUFiZbeBpe6b3MNUZYecgdGxyxHKdb1KM+dLjfCX2hN8uzunm7k7/Pt3LI53w0rWF
0pReik+lZiSZbQcr0HhG1C7xcqGvrwF7CObTOIIjJhB/RvbfWHX00p1b+q8YesnB5vj3KD03VUpn
U/jv/WL92wq0NZfJ19U3MbgZF8F27PmOQ/pRs6zSzZW4wVAxuxdtUMzQgYPC/dlNqTMDy1fewPsD
9ApMFcDFA2UtmJdEtzOGZRyVZJYCnvS8xV038/OF9idtvrSfCddx5Z3uYokhGf+5/XbXaJYXmfYY
fvDIbiEThV2f8JfePvkm8RWyKesH1GrFyQRBQkOH2pNUDyH71lt+4rtTLUEoZUChhNM6XCvUWTO6
lbmZIHnKeZrXAN0hPb8H70H88PVXCAb5FjwLerNSZ9woR85iRDMd48+wfV+EfmEkFHculLvFF+5p
tmFyMz+3GD9f1gojx9x3xbk3CC+tZjGNGOgM0yOea/AXB3AW//SSJbQSYmrOqRuju0BDMP3X5g8m
czIlZuNsyhCiaXAyUMVGXqtztsfRGTc7/KnrpbtUt2oYAc0S05olKKoVlZxBzmlHU8Km4BvV0nlt
AIDNjAOxCCkfnQzbyogblRvKfSidLTqvCTP+UTi6hI93WyXnwMmE2yjNzQEJA/AA8ZQ9aBdpmvwv
+TmIzGA3xgknQVgQsYayAtqsRr/37nMgGiJbwsBsuezG90k87gEZOA7SeZGobFlHXVvFvjlFDRNn
4SQ2lxcRTag89qMPpFm6BQ8gY2p9K92vvj0+5/YTTfL7y7vTqdtPhvb5ELZzp0ZNx/fsIBkdaSyv
bylHzU1eCfGW0b7wujf01UtVB87Q7Xb/zcCzKpMyzocz35yamob7p0DzqjUhluq9XR77GJegcm98
13KZql/oxP//TbAgwfF+C3vNF+AkwZnrThSBdWVWCXOjai3Rx99Qv3XOmxR13G/1qT/5vu+M+/ed
ZiiFbOHe8NtR9WmD6x8btiNmT8XIpHYissbsDutRfp83IkmJhePfITM8AcWUandDHww/maEGt7PV
QJVjEKzy6gyxRB2ApjwQ+/us60ddHx4NLwJ+dQAZZfE6wkfs7Odd49QGwdNJK27t46kHmQPjq4Q5
fcmGOIJd7ffkaYyyv3loegWjz6TxS7pQWJAoM3vu9bwZPXAF1RfQ9JteKHHinCPX5ausJWLJdYu0
oiR00b1AzHZB4T2K4C3oxlc+wHX9BujYYtyz/gxN4PIbb/fKBgikqBMYTp2gEFpvSp8+TzFF5hfu
LF03YHVhKzdwhwH74d8OMMeNu0cX/Y4QXAMKUqSkVZzqyS8QGMd99mbjI9F0wzNtyqLI4ivkobZb
3QMTr6iCJPR3NPVai3ngqrtDQyUqF6dpCmzwbAlsQHiWVEJO5mUMG5U2Hwjc6Is2jFtuqufMEITt
SNY1UqHDiZfuaKwSCIGGNfdTdxFBcwEg2tiz1u9TOTGEGicGT2CLSsTPnuTo1ITOTW8E2L5fwHCS
Orx5LOEmTDKdSi2BIQlXNzcWA6zc/W7A8UY/Sk34M4qamEzRJXhCOD3Htu1DR7ckhglFIqkkq4GO
kNt+2MnjiDq/ajaLi6Np47TFdzvzoOT0ITxYNbTujujwQwK8GHGZ5TTGWobOx2yA/CnXkk3SKz0C
j4qrzHatyl9a9xyUdwoE20HVQRv3oE0x1Tbe4LrM1TNx0zV4Ft14PgUX8xQq+qzXd7c796VPfwvZ
zfl1wUF33O0w9fFlC1lfmLRry4zs2YXQH6c+EIuLnUOfdfYZoPoCE018xzA5T5olsKGJZAItDFS/
nrPgBKvyJ3s2HuNdP+chLiFbD6ky5Jad4Kw5xoUgASkiG+cEaeQIEIqV8y7lOYkCSQ2Z6TAghVFn
BL09c1nVUxpPJyMSYPgvJR/YWoJAIkSzkhHqm/gyQcKmWjTSbhYWC2ifmbIFOcxYpxNKFiwspD72
0cO1ZZ0sOSFGAmzRpPG+AV3zs2kE1rTcJgPX+/gO7R6zqomE6dkDvtmyVe7I1V6jhL6kpgm3rMyK
t/1fli9q4NQSnAXUd+7nCHIBgEXTc8bsqoP9dw8ErkqDOL0Eq6LDUui4ChA2YNZ+sVIDQOhbfMpy
EkdMa/j2ZhBMHDj5n9uq2KcpDmYkHUCffdltt0bw3WaC7kbHhbNMkwlsGhoZIpead/DZ8q7WMcQr
6Hy/DQPYKHXIwotS2PG3IDfHqd1MzF4g69D/sDamRlvdLm+SPVkyEc4Zie/KXAWG9EWDbs/VHDLO
E0sDrdB510DAOJiIWYULnoQZuevD5PWFUYvJksaR7rFOoWCB8jLObOYBa1lwWQfUsiIckvF8rFiE
iZXDQpJZBIxvf2iQ0RgAfp7yyacqCJwMYMU/n6grBK7DVGd9D/CfyhYBhYgeUdYB9FD6eS8zguUt
ZltxbOvDdfqNZJI41Vk0SOLXdq2P+iD5FPRap8Ffzul0wCoks3b17d52/BkbWxtfILl7Hb4lDqR6
/45Z1q8PrFdz6urhdMPTqk9gHHKSoLmr4Yc9vCaQouIlOngBkVcRswySrXoHc4o1yoWteNtJWm9B
AWYeKIw1UlBncn/sI6mBUrsGNgQAYN0Lb/PwOyenG0lZ0z193lRbMl7BsGhahQ0X2AQakaiv1JKD
UCCHsQajCX6FtjnusaHP58TNnE8GhWXCDTtZ0iYX9x6+T2vSL+mqJ5N+QYhgbSAMbwfCcZrAENem
IxQ/XK5S9dynMk9AQNUttbJkeF8jKaUD7gS/MOL98qt/Xh0HqXSFZVPqZldj5uhMrMLaJOaODizF
fUQ3WMK795G93GiK5xTRGPDXcN6/nmTdOGmApksHwh1krMYrmt/CLa5aVLuNUJjGOdi8SPREjFLP
aBdxeA31vJqnSQIC9fm61EXJro43cjvBpWL+ORzci1cRmz2xKJgUju98UiqcJw7m5BkUz7R1v+sS
faH1KC93Kzso8FUMKPStwMxk/ufrK4elaehtEgpBVeG3+oRaJGOiRct00gxZJ2Ur/kS/Q7nGvPBq
p8rbdyvGHsASqW4/xKahgBToilwjoHekZWtdhdM1AnguO33WBlDTfc6eAGfjQIzZvisSa9AR1Q44
xsElvrLqRdai3MVrmSnyQOvFnLkgvYKnQSiqXEXqyXfa1vNuInNSovaMZ2s1FueX71WZ96VSHH3M
Po0WglT667IZ2JDUbsa1AVDV3Jlsh91lMGxFDhb/OhRVldMQAhTQ3R717ENdCAE6D3VWsuESAYcL
SSTipdUV+cWHQwLDxXV/o9XR7mXpK+k27kZi/OlpWfLgv64QoGHtJeniBDEx0jRSve3AKhhM9aQf
IIMqroPAMQt9FObP3ZgAAmhHT/tElYz1VgBVEqlJtGwRXY+L0r02/sWA/sQdxxv1BQldGnQpitTU
fdhIV2hcuo5mNtLw3AO53Ae+YubwhAeg9kjKUYA7b/cZNINshljgpaJCRnZj8YbwjKor2phnuCOc
AZRJkt9KLankwpxne1uv2E/U0w+yAltcIFpK5pEaTKXRKRdgkbc/3Bx0BxMtFHe7aNL8JhjaWJqo
qoupItMYqh2Mxenq9UZk9wZ90/a5h2gbhk4SbXt3VRHjbP+Y5PEi7AVnTfbKWcLkFCyErNEXSHw9
hckEJTPP+McVCGgVnG4B+xdeDGZ1Q48QL0fsW6xDkQBQR5IVAw7v/2QZKEIGamnFOtFv5iWeRzZN
oYFLYjkytHX9YH5Jw48uK04b9BhLANwcQdzcu8m08GI0/+7jFOnbo/EUe2HiNxBDmHnyBBR/5J0T
9b0XWqJzjDiYF8gkf7yFGDl7XgvSarh7aMsjdLN6+sx9x3oe33Jd72qbSR7WjRyLrul1b/TwOdps
Gm9ykfT/jZqbpyilwhBDA7YkwpvhNfMUVv7nOnt4mRAFdDzGUKr+I8+eqEKB4cYhgq2EmRsKCBcQ
Je0OtVm2wlTkwHu7k5irValaI/ki1kdfEmh+aHy7pQhTczAJ+Qbgzb7psTYGtYyGkvEv2uwjyXuw
RYxmSanNL+3nMeJfrTVcI8wXOyYeah92PUEvtJf5dB4RBqlXjfd2wHdWrsxP84Y9d1J5wcYSYVKv
+jxY8eaOfngM+MmAUJ9ogTFFFgK0PGENAHFYmJtHlKhGgslw6KcuONQzFpXF1Z8sM3R7ZYa9/CaK
eD3jocsmnU8zNTummuK/NzsprRNp9us8OQcrJ5fUckhwLFMuqD/O0A4+USNLBGT9cgh9D6GmMTQs
s9AaWdXqldezs/udPNM9Imrrb0GmWh+qFknEiDfZHrKijZqtCDf3nnOA6dL6/PP5Z2eNYdWxlbgG
ErSx8Q/YxDzKqFH1j1YqheR0LXo93CVKagOMDsKakjE8iW8yN19NhOI6b4DPnX4xbzUsu/nozwtG
fEsYtsTtTAJFbyWq7iO4Q7Swuu/Lxousww5JmqtM46VI4IL1XaQBoAoIGDw4ClRWPmv5Q7Bf50lO
6Yfhg2XCzpZ4ZkOGGv3mqbmkIca/AJJydkaAs3uh86k4BG7tzJWFFtkF5QL0vZ94DFKM8Ql6SN59
Rhc5kWJnjh+J5OaPUCbJwS2eIhLpuSgNf4CLDB51yIUcScax3tZvBI0eZHJovwLztisy3m7QzFae
2OtfptihhPUT+y9niviEpguo6T0gQU8J3WBjh7vvPZv+kqeYUEnf5LOVM8Wol9Ts3bmxaiiJTHDs
UI5zG/WII5JVfqWTlhIbbph6HpB3vLZ9i4E0VdAqQYpuRPeIDNWrjCE4OXBt/FLvNXJllq7y4Lx7
7WwrQN+XzJz+Wq/5alUkIvWlEvAs9NyPlOLHpVgQ+PPIv9yeDxsQafApw4OTXkHlT+HWWFbReDIF
Po7sAUakgMkWdDNDQX0U677P16mLu9BbzzRxzkL57GMjjUTGcIA4FV/P1wdgSStFhPxXNK72K4Ww
DzqmjltgGvFtMaHv5E36/yokjjg5Nef+NNdM9z77fMvDa3HA8SCLRbn4h2Yo76M7DLy6T35EFBmV
sTWCsdhLGMHkN2AhwJxcs6vaL5VNmhGkBLhM3Hu5D4MtfV/Hncg3c8y2p5fSSWAO/kdCwLdJZDNF
qyj8ZWmKiIln8wAyoaMremHelV+sJuGXk0TDKK/ObYVl0kx0V1WJEdkYuTg1E0nmEubdIDXeUc8r
mcy57CCbiOpdxP+gCxOK6nqq/LR4mzws/RUb3zGXs9Cfjjr+WGmIkZJdsXDC6hueFAonfNV3bXob
RBkeESiQj0o+XQ14sz5kp1S/jMRSmh6KT7WzK8OzJnzVsZDZHsnI9cSkGU1VBp2/5LEzMW/3Ytxs
TPTW3JHsSLIiqCTkrTcxV6k/wtJcwFMT9Tl6s20EeATFV6FEOOmfAnFyVOds++A2cofh4qFN2gQJ
98k8EmmfNzIiinJzUe6xFER3luQx0GoSLSIqIsF6hLx1Cs2qu40ftufZcGshPc5hV5H+Jmj6Ffrj
EkgNxELKeBSv7L8X5X14j/ekH+tojT+hUaqrxCh/jCXmGjPbbzhngDMVqeeWGmNZYE7s2Ug7/dYk
96Mj0hFI7euU1Qps8CThdgC8DQOEbVfei+icmgzDWHEntAKy+IPypc/Rb/9EiopnVCxE8IMCr87d
C4sHM1h9YzLd846AnULqSc99z+ZLWe/HdvZKkOsr09RlfL3l0h3x1td6yBIpyWauGiYUtOzR+rKP
BNUvTRY5xcI+T7R+Woa3TQNzBa/SNAM2A16B5N702N1ect1UhAG2VPSuBhs3w03dG4fnqy8ren8B
9wGRCpZaQ4EvHp+gThSgdoX7iaa9jJr3PNeLkBIOlZ1o4gLwCMhdcvg+CP9hFHBoPcL6QK8pPlhA
5y88JKxJ3EXk+B00gLVz8/DSLVzTkRa4B4DtWevvNAjfZuhYebdoYZnW6KSTBnj9OMAxVMd3C0wu
u6LAI/0s6tuZyOFm8Dqw5wxy7TQfDWci3pdcNNKiNyIy3vkkfr/wyAO5vKHLBLUhE2yQ3//0YvkS
EeluHug/GQC2lPajxEagQYAIl9vsTrjHNg6ByVqhYHTEOEsVMWl1Bd7pN+MNVg4ACzcDfZZ23ehi
canSR+Vm+6L/2AwQu/IQgp+54/S6casSXzo6AT+8jkr0j/hF0CVslFRn2v5+Japd1/Ht01fhpyHL
fzUYxA418O3HhGqMOVDd3ex4OSXGoDq5rumplEKrzaUoep8hMa5bfQaviL0K5ZhbxX9v0sAkHRmv
JuyI73PrxkHH9c/TQriJ27slPfa4SYHYINdoH23NMLEoXXLUOnNgg5WWnFbCgBgLpixJ+Kio0fK3
rpSs2DeEmIjunfwb+mwb0iME4uuhiLOXBVlWnfg58T+5hkzOczk7zAUJirxW+yrPqvyGD2N6YSMx
PhSz1pZ2uIITAaC7lbGwJSsf+flwwnS+lFBfD8Ca9jrJI81yfpG5kflQfuw6t2DTrpytLNqlvK4M
Y2zHPvR8fpzwamdCK+PBSu+WBJ5noWtTyn9UKJMGUpH6axEqU51gKges7HPoKBds13lltl7/5kjj
7zTyPLC/37Eo4MqwvE8ZCv9OB+X5oRslcFya2NbUAUb4T4B/4YtK2tcmKxJRpZGRxItlfQoysvFf
iHYkZW3o+CxyNnU/Wxg6ZbWsJTT+SepFqZ+i+drNLRZK3jWTvL1bpyt3fmP2WuB86t00YFTy5pLz
eLAUtqfNrFeCvqXbrDFlGW4XkTdVfRs3ToI/cUU5SnZAu1rPqAgbmRZ5GQMJZIMT4Onzs6RZxIbV
O7E/PxKyffe1gyykGAHZjkf+E49Ws/2mz8n2G2zcXy+Lko4gU7BbhtxnC0GXpffzgTyHbZVcqdz3
8v5z7VVXNo30CC4XP4JkMXEDaUmmN0b4fv7p8c2Vxql+3faWhMCBICGPNdWWVb8KdLhJCQC6M5pc
LlHnpF0rDor1lZvK5NsUu1iMGpbv7gTWcycWSQzew5uVPRNX8RVXmBrmmFzbLPycpGNccQD0eUID
8wopiHnsHNkqoYC2P3eTYjfAGomYW/OUcVtWllk40QSmyAz6bOL7D+Vxf+KZ5rozVHWoKlDu2m9Z
9QRzMVVILXJjZSmeOWCPMcCnoSaLzbsdjuEKTDL9ymypCl0nDS+htkscpUa/AS6e3nq0Ntasw+IU
hazk3RQ8twMU14GtoC834cjmgxZZ4Tr4Mnx0kLOFVOhEaRXxIvrmXeVc/MTdqitqgMXJv2O9R3Vq
OqRK1Ql2McFBDeEwkSak6oyYaLe9KEtJ+MAZ0aFMbq2uynsrRu0L5LDBrayM/fSTkHnZ3BkhULA4
fuxryvxVhXERxNno95zA4U9ZnXt2OKUYC8DZw2Oyr3Se1kn69CRgqVHbYGiAXCmcnXsZqp/g0yYV
cxRtauXPlhoCbSWTFAE4fqG5AwSJTVVcE9/gSgbZhXiwXIIhsWxZlwQfXSByL0Qg4KMNtXddyoNV
Oyx3jjEBStygXLXe1STq8nuunGPPuGpF8sQoze2pncbiHmPzV+MGt2D6524PbaAXlusE4IxmobIx
pjaEYck0wG/HsiYR//WGNFu4rY5gfYwjstMPuDEc9yU9S1NUD9VSeNADDMA0Jb/gOSBSzxxSJ+ao
H5auDwNTlOlBlxtSjoQ46k1q1QNLkLj2hL8cM0gWd/ERlEYN/CIbjdS9LyRZGFwpsFbdyhc9U2gd
sUmc3iskCpzGqE+ZaFNkir72XQBoK7D+VIfYvacQxdY51Hgwmtuz38mLt2kw8TiforKkpK9fQoBc
LmPPISugGwso+D/spnOYpgV8WKR1iZoTU3mGJaCKgUEK9ML3Uy6Xt+C28AAcHpDQdvZDZb3tT/Pn
G3Bxxy88bVYuzLtJAeDM3qGqh5B5sF+TK6vn/czdCVyPMtWXU4I3wdQcudkwRdYT3I//3GaK8ZIi
B9ufyiyaMg2izrlajDXSFp9bHgdw5LGYpH5bDD0J5sHuISo76E8K0OympjOM4JOnVaj8WbPzZqea
Nj+53CKNnh8p3ON4HCluIu3Xb4LUoOPsOZzUvTij9Zf2UNriGXIq9A74kxstZYkfiILwXUsWoN0O
UtA+2D64N1OftalD/fXCi/IU4689n2V4qkubW9tk1fthNxsj1uV9eLeaQ0mhlr1vJlteyOCkSfbO
6AWWbmeAQ5asBqojwfrAp1FcReM9GzEgWH+kp4tP8XuRisKw0B1E10RtiYOPJca5nNcFr3JG2v/f
EE3+A/22V1oWO5u83ryspKRXchFIMX4qi5to+6r/Ax8dCUF8zyoHd75s1Oru629+Sm0gWII9pFyO
SiQa/VScDi9c4ZagMP6dUupzhOuKM0Gizqzb9j1a2F9PDc7u9v7Ann1OciSDc+FQpwg45P76PTGJ
8z+Hf/eXRlnHkXV29tCIC8UsmNxVrtLm/IN2gKqg4vCvTQ9FWSO5Hq9zLQnYXYh/Wa9XLZsfAMhe
2uRSHqgqUJ0WMmm6zZDYbR7Foq+1Ts6BH29Nbhtqz3Kkwvs9ypdha61SzMemWitWcnjejyjovn7H
xgChswhC/jJnlyBsPKgUXHTb6xChFGvdaGjm5QjZTobA/DPmHqzwMlefvzRSaFHmEdZbK1TrEmD1
pxVQBXG7vREyBYNLxIYU6u/jYNJV4XRvyEKoYAvxbo041uMUNAosgQmOpYRMIG4NejIitRvQhwM/
+KREtVkBzFrODsggk5Kql2ls90ZEd7pMpY4Xv9yuqZr2GwgS+ZB8WDhTEThUg5QIVJzLDoxWm+Fd
Fkr1ty3gpjrByrlkDuvgH8SW6XsS+0JBzEG18fZwKZs+VdltX/x2Z+ldbF3NLYgRvVRKbJWf4YiI
M0YvirR5BquFxtBIJ/WVX3AirlPmrhTWF2C+FRWhfQpJJuSoDTc7NZ2/+mm64eIYbOURW0pfK4zR
Pd6ntTB6VcXWTXH0sJx1nXmrLjlwYjSgJWgiIz7KH37/pE+vHC0sogpOrbVOuWrakHb/2iMei8hb
mR8rfQNETyb6AcHZqC4vd2dfZtPSPceM8eGXvxb9ygEIB8C2wEywBHKfxwZB6lu3H3efyrGotSoo
tLuKd+b3l4x8bkeptBqYIALxnLW05ph36AfKdkFdtL6TKv2JMFZQAOdzRrfNQHjOlSAuTyN8JfqC
Iiq6yu+pE3fhsVySZdi4Ug2ePy2Wz0ewj6g5JrhXGY7Pb8aIP4oDc6uB6ZARc4SM/P6uI7WT1E5x
SPL/q7hLfPrxcSYqLBlA+tB50aJeQGgIlCGHoV5uvdG0qZxZXwS5ITlWlneFTXSlITt3KRyLIOcK
81fVdjQGnpgjC4wtgAjLwwxzd8CSTQQFTjINk2XR/0grpq5pOFFbmRDCZ8O3LucZRtB1yIaJ3385
RzrilsthuRQEUl2a9sQCKXn24Qsyn6ek6TC8pliq0smsYGEi3BZMTIrzrCBm4X32qP2eTwjVPMoJ
rO83FA32Kywu4Hext+Vz0+9VT1MFUMjVNiq1abriNQK+fZsL3usjaJ9ibyqSd1Y8fk3OvGSdWCZ8
j3NUHE5GgLLQAZ53/rhu7JNAehmUkVV4cPyYRY7ln+PSZJ73b9unLoKVfhYmB8uqZVUUzjPYAqfv
EaATBmhJwiZpWbaysmHznQ1dzQpdHmjXqSHros/vF3sO1/tH5F96olhAnQQyUmxlkSn5NOYQLk2Z
UV2zD/fpAnc5n6JqMgcQBPog7cU/NM8K8mCLgHPc79DSO/fR7/6b+0zifQ83x2/uG1uIHVqnPtmx
+0Tz5HqMoG1zUd26KgoEF/r+Cddf8bbfmu4rXXXu3hZaJmFaD6AXj3dqXYKhLZcCgEnAPSCNFrYp
H6tgHTNh+G2hoQy7ZO3qqte91SwO2AY/TvpbiLong9a6qsBjrx71RFBV4KfVyxxySP4dZ0WqzcYg
+Ot6ObcxC8vv49YM2lCx0x+dkrUvaun1bw4HRiybCbhtcywfcjzEe3nSLMjipejcyo1mIiI1OWx4
cQVk5YxbiCuFrUOeirzXSCgEnvAvU8dePG+lyBV4CsVXV3qGdIsb3fLpwn0F9zweL7+z2fNL2bcg
zIv2nupZrXCYACfnx08i+f58w6Mb/LqIlc6RATZGK78GyGcGqZPMWCAU9VHBGrQDrklVbZO+FdmC
oEzeo8ZahrF1Apk3LmH60q5/zlPT6YNze1OlYJVTgfaT4R1wVe2BGiD24LKmmieml16S/aOAhQ6V
Z9PAiWsatEFHGoFHtC6/OSSMiR0x1Gg7P4K6hpj5l0DnyqOy97Q+w5ikGo8e88Q0aFZhMX4cSD/S
zxEoTPLtFsx+6FEOYE4iJj1HkeiFyyt/m8MWcM8JgMrqjfBLnQ7OxPCtm4I8AYYJbsl3W5BQkgk6
4wxTNo6bjFyEpjpNlcsseUH57RwqFZcMNP4DjiSvJnp37QMsdk3bKnxA1q2QiepAey7bTvBdcomw
v3O4+vLKon6OaSdqLib0iRpOHCnPfKBTKftvtj+OhSIZSJE/xMV30CHvDUbOtpfLDJShkod0KVJI
cl0kWYqmnYLf4YbiFADQJ463eVK8HxR8u8AXSNWAx9xFe0WFjlpM3zTy/1nQuaUYaefhAuSSCHPY
fz0gPtl3OUw5Ko4+0qqeKuQQkRr1moOlRFVPAC3b0eu3KGAlYnuAE8E7qLf7WZE9wgkU52WpwKKv
2RzbdDud+ZjgpOjFwov2ScPjuCeMcN64VIFoux5qdGWkQ+rcSvsR86zGvPoF3zVmtldgBYceKsy0
3ysSLcHiHuISNCfmrIkkjAMhxaFSQ0OmoCr6u2iTpuJ5fn6pvUNk46RahZAK8gMEaFhV5wfDBfjN
qSf9BkXGydkLr9DVo0J/UaSsbwzqlpwHxWJvV4JQA1sSa+dJi6LYoPlu9TGezwEkkPoT7L6YgvVz
7r0d36Glwa/hZeJGruK0pdpGSlBVFSaXQQqDBnhtZ/bI8kXqYnKh+gsfXE4L422/dEPsdNI2SnBO
GRyUuL14ciDuW4zT689RA1q0gt8YABZkhQSEIfY49vIzSZFUMyFxR4pDrZsd8ZnRiln4HB/qQqRN
daenjrdEIl2Qh0BipD84X60OsowPeK/SetftcPn+z9sfgKVppDPEOSVpnX0ZEMZ3EcuRfNbXs1TO
+eV16ULgFlyTr9XZpjvl4zF5WrgPJUuddUq/ZBbzMq+lkWzUpam2QKPhVdWDlyzhgtDjsOSBluw1
tqNhOXNurrUvx0YFieMGtGsjyHljz0vKS9CY/+4o83iV7XMkvzqHIyQ0mwo0H0a/S6nLMTCTT3Ni
Whcnn/Y8ZOmzwBY6S46JiMJLOcRiE79CpUpNtawx9HbSbWoYTgxd3oxeGrzO0yy3RfzloTaehSkN
W0nIOawu4fLbMQp1kdzIVztjXf/eoajvm8OAbuslwDy4xiiyZUlEV+9v/5UjOBmHmleegp5dQWVi
fUUkf6g06gxMlEz4lyEsseIY2En5XmfIlD6/ZGVUjqUeX6kh3CdQUhwDZB82U2ixaDQ065bx8+RX
CyHQgsizp3DJdJQchsrLlJXlQb37+GKoOjcmj2tDM1Z872iqfOgVoU6L2BMbdRLUJ22Xkw5HyXpU
yhXH1qf+ydmv0M1x3jjw51CnHXhoiNo6YZKma7tjWBrJvnsIaRCubwMB2mUu0WXoZZMQhfFzGQGK
eexZBWfR/Jnif5G1fwBbSqZDsHEyo9JNPaeqigU2YQkam8OFJeT+4b3zZdRIEhuP9Kdbuc/mRFuj
LXJUxulqkTYrx6ff4UIC3yqhBPYSUg8vtMMFehRmrO1LFqY/6Mcy1xUlPDQZIllaarzEMDwG0NXK
c5/4obvlwlyVyWzPSJcWo3q6QPzKTmrtKHLKwhZ6mt1+Kx7vfuqIqQMk3/dBLBSKW/HULhpu3P2K
rvrKDp2f5xRf5UXkqYzf1GTSqbYjxZ7y+ouRmnlN+TBR4kgkLyePx3ZXXePcSe1iiQF+TG382F9X
qmu2F7XrvLxNRP2Lek69nSMNK0h9L82wxSnPSUyLxOmPtgfESjXIKv5eEEvTY3UpcYf8gJA/3a7v
6GUbFCRRb6lnHawhdtANiYmpRfgui6XVYtNqLBqgPyZPVCmkYWEHObqM4oyUZxRC28aSBVZFEE3h
VbsNu/EbMg8NMPujKiKGJlEspkOtDwHdmeSTj6xrnl3FKfXpBd+xXvpbN42yi+VjRXc7e/ENSRUB
Sv0WMS5djj3tbUM15w0UmloRhN0BRrkWUN8BDMWltxvkaVj+rdjOcGpokGzaaw2FT4etsNOYnzGa
fUr0qDRp19XzVfcr57zBd6lPZmvgkQg7NrOd1Y8+LmDN8/Jl6f7twTCstfZaFu36Qwf4rfuJiUt6
nHFyEulmNQcIYvTVtxZQH0cA/RiLalmXvz3/22DfC6QCgBEDPdVfnNu7cQYbl3ROJ8rDxG6h2uNl
zx8WdOn7jIwYe8Eb3Ui315o6My+NedpXfJbuI2vo5SloSBPGfe+CGaQaXqAYSzuH0DVQKYdLVFNy
Ax96dYCxpLMtSShd7hgvcg7EKpP3lb+17asK2ymxujplEZ+oT0Yvk6uiHAnzRSEjU8SnTOu/6A9L
hJdWUG4CVyuf4sd5iOYylQKP8RMoJQr3tgxZWc4Wmw1vdywf5GdI9jq2LMK8JtPX3WXNGtjS8L/4
kv9tJD/7Hq7VV/CY54+VfPLWcUprW1j5e3rhY89rcnsSKKlZFxailn9Q8SK86M+ZHwZNXQEgeO70
bu/Z+UOpQCpGI3e8mXdaBAa1X/qxmS2rPJYpqASoFpmxCjQI0H2LDrXqnB12AHCvt+Nb4VuUcdk8
tavNDEq1LLdsAhv66cHPBAfLfFmizL3Etbwji44l/eHA+Px0khii36g2f4XKUqlPIS99Yteh2N8X
Xq/3b8wPn+ekNxs87EEtSENStn4P3g19VT7kx6zRQ3qgxLg3KJ2CYICXXkPY7djiVCrx6pF+yjZ0
aMxopYJI+2LgD4dT/p6brT7PwrilGLrwybbCt42nbQyfpIQHL3C+Wb/zkL07VAuvae4YM9UG3DKR
+OzrkyQy//OMJCVEJrzmJXZ0nt1AToYG/f53YMUZdVYIM7LhHyO0BzFLPJ6Qxh1X2imOqLzBSDbE
kqZfUAC3p3CnK+OakVDY2noUxDPtB4NWW3eAFphIQAo7dRCTs6zSTKxDuOoyPTmfjObsDM73MWlh
XM1DfFLaRRVsz4gnPPVKg8V+45ptXk9kXr2QJjaEuAMVKiPH3vyxExjYG/8yLLcGV8p6NkdP6PZs
g/zrcXGQtfhHc1OjcbvaTOxi5suGgo6yt1z1WMUh2ZXJfesLifgAb2Ta+kCdmn5/pkSmg620AOxz
OGboUAfOVyOy8sR08gXNzHtnQ9Motu5OMdIVa88E/fxY62xRFw4Ngu8+FENWUgkrfBp2UYp3665s
VzaPgGkgXBsMX+8jDEkPEecnXE0oFGbDnTLXfcboAX+mHj+sjPFdpLFM2hK3HV7y4U6N1WdVhOZE
3wHAKIn4mwosSyQMNKWLs/NOEwHXFll2y88HQeRUO5skZ0/P6QzP0mBDeMFkLoSzPDENrDp98lHz
nQowQYV2J76PeAl7ybgqKjXgCHkA4XqGZqmxmuGpJ5c7a2RiV7FfYBHFVZJZTQlEQAQEnrz36xRA
tX68Lh2buvpq0lpyuO+ewge1K3zHJPNcduIe4BCLxS3p8HaUMRNpUaUD7ETl9Uq3MLRPRP20V2PQ
I0xkfkXfXXhil37/ubXMExN+8opNrfWXzGWg29kcvMgwrubtzJhKYcl+QN8xjMczLPWZAn8RhPki
Bc55vMyOVWLlBR163QWD1NSHHkOtb8aHYBXAUL+3plLcQfzLEWTDE6WOncCGokGjZkdmVoZdF3Gs
4WFekxrOONU9XHSH6+EpSATYWOqKyBsh5T4fRZeXnCqo/z161fwiUuw3ep/UVxWjsW+W0I/tOWfn
DLtxCOXru5/faaJMmzFLoBSojfJtRtV0XueQwwgxhPhIxeNhIItjvn0Oqm10HOKHq6xOKK+q3l2z
mvBAw5OiEQz6Bwm9Na1QDQgPC3YTzWVKBVp6DNp/05hxcJqxy3nUzD1XCiGjWNvgGBo42Lj3QJfZ
rCrHj5ttwpaQOxJW9lzqJZgsm2acoFl/3sZiFeRCA0P9eV53/KITCS0tsRCEogfJULPLQcoLzxLa
TshlpesN7I1QP5KoiHIt06MLxbseOx/1X+r9UsFFuqHSVDlyudoHg0jeYXGp9kQ78Ab0V/9Ovz6p
RXqEVmYROZDB+FLHB00ZAfX9L3F4rtvfPORBAXCAxd2WyPSSK4vWqAFkXlI/EYvs+KMO8YeJh5wX
mDH3gqhKUkqZLtDxmvaMZJkKQ6Vp0NuolEmXlIlJgTNNmujvVAJXwlIqCvX5x7OotUxu70Vw/Uk7
l7NTaftIKcSnR8UIQZC1YgStce9ivgPv0NKd5QvxsQkDtbp1+YMXaxIWiVCPphtJ8XQVgg9wj2Rz
BcCeYPIQ1i6mxqxAjQibRt3fr2lJTOmw2afQ1K1rHRk09dINkghY37k4CpyUteJQ8lTCnOAqo4os
1tVYgIFUs1TzdgeMlJH+XggQljkKqHqHLyotGUHS8KxFmkEy/6WLs8DRi1g4OO9Pk9N4CMBj/8qZ
cufKc5qRk2Au+5hV5dutCxKY4/o8V3EqcgkjyMwpBwJj2puZIUNzUIVc4gijZTzqnOxDLY29cYFS
FHdcjh5IP7Lk07m2yFjS9xDpokHEra2GTkN6siYRX0BNsecrfac9yTf7ORwvppdPj7UzeKGpHSEw
WPjN1TEGNSK7Tflq6Gl35DM5a+NX67I39bDjgvoUgY4km2+NtHwh/FeLlz+q6zGluzpQQE1wLuYK
KVsGmTxsUjOEPkEdZ6LW+KEaLdddLNCsD8xjN9VCVwXadbIAhFxql/aJaujhIMQ5sLt2rYvXVKXt
ccah4DFGrQOG4iP48hOs/SjsXf8udOnjLrv1jeh+lDVnQZumDIePb1ipmX2QtoqUWVGsKEpdK0TA
kLyirgoKLTqXXTfDaO9NZH0e84f7SYbQ/Qh8RsSpJy0bu8uxPiWN5vv2TxaMESETAmOb9cPSJEcb
eXcwbupFFKavO+7HhfEuKP2VeYq42RVD2stflaBHDLV7ub4QNLv0AqlXAWw8nraM4Fmt8FrM2BMA
zWfpRzZuIxg3EiqOXUspGSwy7GMsWNAzkNTq0ZLHLZ5VxZGf1N8dQg0kL/abQu3btSmQnVwEn+lf
0gAbIE6Sr00xiHoTZK5Wt80/dU3RcuJpZjOqA12jRJ0vJAwARD90NjKODKoOOaYscTiz1EEJVqjI
E/nHZPjrhT/Run2PXCEBe7bBVpDKvuEnUb+jEPdkDgK3t3+4tnju7WuDUGzjrlnbH1EE2HEA6QGN
Tk324VV2OxoBQvwvhaMSAyQqEc3I5uqLQUU7OJsJErvNkmhrXw79/JjmTaAzGt3H2bLqWsnWx3Ds
enDa/IMFWLfRmiVr59g20hrRKKh72fxiFqPe27mMGaIHdYzkFXo0XaLVM+mNc4ZzwO8v4FklRdyk
R13FcQM29p6PetfbI19kVkkFCeMIm5fWdfS4wnUD6ve30YwwA4NuXcGO0OxkB33GKvRcyhF9AwV5
SurEdCMoBbyZyzFsqBF5rcgynEx3fBUP5xE4qQwhiwpJO2qQKu21JO15983Vri6WfhQMCCyodHTm
r9wXXYW4dQBdJT7Uc2PPhJGj3qCoDr5rw7xZH6KKcGiwV6rkVUu8/q+QifidjpuhVP4U1dQUQuGj
VE15iqeHSl/LJvEwhmRpf+IWYpZjOgPun2P8veyXiEwoC4qdzXdkuxxHSmM0RO8SNvG5mYazCaIh
idiACOoEPopP1cUGEOgEBHFeHQtKZfkQf1s0BcVePW62GLKO7QHyCr389BbMQ6Y2i6JjRv/DKYrI
2FgSZU+s9lKJjPWFHsheC9BoeO2Ug4kYr0Z4Fyq0aZHoIKbAhuj9KDjdv50WZUI8xq7jJw7YmDpd
3Ku0+LatkKWiO0cm4jiApyeUOSm1/t0dpWH8Qs3ZRstsMo8UXNobcMGbXrUwv4Dn/DImpX6ZL37v
UbBNAUWrHQ2wg9guL3reHIw30MsVXp6pPifbQVJHLZsCZiHPYYq4kdXnlnyEbHW4U6osMlR+oQXM
YSv2ylX3LS9P3z1Gro2/ik/HySdrC8UfVKcaP9oqB+vm299zLMHcwCcPNWa/lszSOyPPPZLpFgY6
rVv5nrDPzabvDbQd9duWK9AdqrEerb1PuVnefPzwWHVosIEuHPGpSHQ3D3m6XCf/wvZ7lgBA0EV9
porWuQW/MShVyQTTvnFbNT6cl33QBwFAhLU8a7/7XX9hZyloqQyenRCdPzX1UJh1u61Wy8xUDIol
bJ12Zpme20Yw2MccqlLssoccsknEw+kEoZ25/KA1wjuZdMHH3VttA53/gGY5tGIGd3mnwmbQTQk+
25l3Kp/uJDVVJ5zsF/fTpZ0TMB67wd0TIxhIV+42OaSgVuC5upRCe5gOVfNWghW9NBAA5npjWEdw
w89UOASnnUSJNTfiUQVmErbu0oSSkVkJ0HFAYw+0McuPHj3DbcfKexYrBFCbDRmaIyooCjkIWb57
gDhqCsDZB4xv1U/uW+fulcpmEzow7mO7ZSPC/xgXg3UrcCpPUH+VHMBNynFp4wAtLjzituNzdfAG
zs9LwbRoysyMSljDTzqwQTFYgGQ2SWBtulTR3TDQ8YykqGWIxm3R296ApwSNlJfzspvfmNogk+Al
w6ph7/8J8CS47fJESM9Owy+rAiEuAhmTyMWPQ0/uKqEMsYnr2Q+v5mlKqO2tQ5ILEFR5nt1Yq4wg
ZIx1DHJt5bfhknfQu31SemJF/Kq9G4EmGcHv09sjg18Yk63hzDV17XzZb54qHcV95Jquj6iAAyHq
lRW/Ik2VS/ZG26VXvTEfVxEQ1Np/e9HNlJgtZAV6HRxgD8zi+YfrvzP4+7g7aQU+x7Tko1UdUcSh
AgQ5nUQfiTyWNdI7FJ6sVI+lgefe94fW54xQvU7kWOEuEWUGhZ6D1o38unEjq1HF1UqF2JKelPqj
e/5lbmI/RW9LTuuHl3Px7/X8ie6jEcN+Uy3HpS9kBiWOlTkDGBWS3rYoCTEXK1wfL63HDEa8tsdc
2cpS2Bxk47a0YnAYCaJocR5YTmLFowHuujedCRwGJgsgOBVbU5TfGs6BBDJgyCX6MJNxQcPv7xeD
+cZ2Q3iSfzte+trFG2tIxcosDKeSy+bQ+NyZ/CRv4/5EXgT9wZGr3/jgAVo9n7XrubujqtUt6DBV
FsgOokCMKRezILn+xzxaiqIzME/jJlfDtpANgZ+aXR2K2H+EZkiEGzk66IFmUPahMdgF7cMQt/Bj
p1DNYfAqpD7LaL3mYHbbAFAGRxlD7nl/fBPLA/FyznURybr8QQjiBNWWvDlRkD/34lcFzZIuxlow
GY9MCWz/hXj1pwJtIoAfwV+k+uuYwpUakgGvpitj+Ojz+MrnetOAsjJ96E3DirjceIgRin0iDfO5
m1d8fEGB0mi5opr9pE3BXLcUAyZN/RCDxEU9p6J8GqWGbe402C1ZWAnx6Ag3Y7Kicq6lp54A3zVm
afaS3jZ287pTohJGgLXJ8le+0DL+Oi4v0gRgCJ5kpnW81+jIjqN73e4Jfe9herzADt+TApnJPYqr
JJmRzinWjTTd67Eb14w7N8tHwVgmguTHuo488XaMbsylIpOJnkWoYIVUyboLEw32VHk075wWPKxC
XfKWbfiqJzx90XUBp1i//PEZdkVvoCWAg/WoGzvmaT1k9cS4F7MCpbdgJlWc/7hGPkH2PRfI/Vow
CCYtD2zFyfc9sk84JweDF5KPXYBKlUcz0OGc9CXt2q2TLxoYTv206/2zy05Z44wyaDWNugbR6f3U
4ZHd2QUG1QWwqWOBsjNC4NIFMqIdzkL7C/jsYpRjP/Za0ojYyl03p53v8Gi6qIEuW5u9070evx+Y
wN801mg0oSs7iVXUTPnE+9Pjc5hsWE7uRJF5iyQwjEkXZhCcWfCYHz8vPrPXnGu+hy6+KSEpi/nZ
qrEU/0BnArwvw+t5LlI8fM3oV9u3XZjBs/KTC0Ja8id9ePlhG3FHTGMZTO+xIlmnOLwATdb1V6wQ
c6eu4YzkysEIliwgoLfj0HIFS6s8nW68D5QQOdsaGfXvqnK/cvfz7egWlziueVe7mFrln5YXbJyA
ow8swM4iXv44sNwqAP4Se33h/Rq+qyDPEBTDXOvl1li1/HaeHLDezDAdKTxz9IcnlHqFJLH76Z2P
0CGFSWJkP4vbmObLSTyLh1Lzru1/oXrzTefVVuR8ifNhP2g5xQVBUGFw32RqhX1AWcLtaBsFa/qr
UGxaq9Uv9XOgmXsNw5l9ni+k67aKPgwwg1ieD9yAWu0qLTnSIWn8sr3cVo5TvjbMMooyuUl1NRVH
+02IaTTDXDl+zyvBOX4KpeQjPWrYFTk+CHolN0TGwZ+h0ODFyovMfyEW9jpVooVAN/fod0KJGHdd
4O8D5IfpqEK/ao2EOi1PamhdiSTifouiRWZaS5E9mamGRQLPDP5LP38BWPhCVUP7hYanTT937oRF
hXFg7gY2IGL6aFDeD+j20qy3YyZxbP8vsbLwpzJSVN1Rrnx2FGCIh8iaJ0Xs7TKAEmI9RMjbi+5g
hwBBKGoDa5E+i5uMcA2OU5ZMF3pF2mAFGzZu1vz/6uv0eryRd1qOZFMZ1obepny8ttq2UpngpoH9
t8XcmzTQfDhw+DVbBXN7E34bcKOKmeSvxtBccCjgHLw4GBWtAIhJzDcOcUvppqBdvSdOEoQh8xnC
0dwL6kn+9AcEC9jWkyY7HBU3eaoZle4d5P9xtpiKzdqkqWVl7luaCc14o1snEdz9Gd0ud3dpZ/Ss
VW8nCJRJun+KX11WhUunWqDAe0jL/z9Ld8TEXFYmnAxBLuxMwQUokgVT+wUJgPXoOkkz9iJltTd+
Qlt79XCurAzgMJyiYFfIrgrKoZQ4pWt2i114F9nzRoBvXmIXK+NuShnYLJIqV7dxDEa3/EU6Wp10
QnkCDbtRopp2YpAbI+Fmy/4uP1vesgdIa61kmooasP+jNheMqABdbBuV2LJn6ZNeEtAJgBpN/DYm
i4YBQz61L690SxB5PR99kMMccXc5xgNnYrU6v0rhSKY+kRtQGe5w5/2Cu9da0H52yEHxSHgogGqH
NEZdayV4MVlNfCf7cTKELXQ5bnS3bD3SubFMRREJ8MamAJeQaEtWn0w5nti9VXsXOI+2MlrMO/4g
glHIR8Vwfb7zMnz1ybE09dTEETKYRtT8pCIpyz9w6yyZMt+vZ1pLNVB4VlY6sovRXN3T+jlnn7Ug
Uud8p9wFZI20FEG+1FfaUKqyq16ps1rHtL/hXAbqw3nzBALLhsi6OOMdXI6r0vjcWXseXaJDRh3I
eiKfkuGcbhylM7lASSQ/L8HYzepN+Ja4f7AIFaUCBbRc5iqjd80o3YqrrTJ8nVxgIUvUM6rvZSqN
wPVI7GCXl5kpEoUVw7LFIsMeCCcUlTfwa7kfZoycuSt8P/CcKSKZ6h6B9AUmqmEIsAGpZv2QGLY0
N4jPehTUQr4qiElO3xr+F2i2FnsDQ60lVW9IJHLA2y3BNaME9/LY9bCM+Sz46XBUqa0k9QH/3R5G
QS1yB6yQWqDIK7wiWM3ihezmetDhRwKUKSUhicMeuKUgnaaEHgtvtU/w8NJa841BWvwXUFGteDC+
2aWKQjKRbgJ/dgJUQskxYuk4l2vQ0E9CbmzOhsy5QgHqh18hNbVHxi6F4/NPbDH63aOgmJJevB5L
keZXUgZctdSYERhppNS2UIMWKktExyF34IfYUcuh2kouhaNGpNnUK1zd2vpOu8s7f1jJsXf+VjKA
yyYtoZ7w/ODXOr9mq9Oi12zXgPhbi+RQGgC3LHIcgh2GG47vcNh9f64w4tLveLyWNhhNufG6On8X
eWia8BqcO46ze4GcmfSvg19ED+bViYg3r9HXJ9f/8zivuNC0idrH9Z98vtD/YNMuAETT+7SS4Sdq
q2KiqgSkT3n/QLXYF6B3qYmFCD4xCNCrXiZ77iJ/PZs9ZjpRPszivA3stECRSQ4JtWWu1v6CMxdb
eWK7+J24Hs/KwlQ7IJbQJPBqhRzMgH/IvszW3eYwfBvlOVYZKRkE4Dbi84+HxJ3GruednUgh8Dbb
vnvTMrZCRDwjtx5Xmu/73YwrbkmYGEcEftRs1hf1IZgPbh2srgIAEHVWkD/HRpxg41SoENmzxOLY
AzJ7LlkSrJubLKxDwbfMbJ8Y1GzNDq/KiM/zCfqGCVCwqOLWcUwhxoN7Up9OuOJavIo8tqAnCB6M
m/4XaL/xrENi5x4WRlWau8/oXfFdqArvWhhe2siCRdAWXl5LuNISY7KvDv5G95qDH7+dX9zfGDjH
Qe7dF8mcYCavtMLKuR2jmnscU5a32mh/cykXY5QIpEfXATg7klCOCEXo553lGUOAZn99BxgUui4l
RqUenyHuOX+W01kcZusyhy/5QX0GT8XqoweYESc7RdBZGYKstEazddYA99BnOQraxDdTJ2jLDyYO
ZGa/bjC0J1zmA1FrPV8CHpbQFk/Sx/ohm7Q48YKuWjCdp+SJW+j7A+oGOhYWkPDKCEc6MYswsEFB
MFhVoEmaSpXuyCeJFbw6ssuMgYJx8Y80UV8GnxWIzszPH/Nz98OAHBcWzRuav324wXB39Ayauaev
1GrNqQ9LH7RHi+9EGJdyXXNtv1RnD9y7GxTEqaBXE5o9QFLD8qcFpUDgB4Qpv4fVRIKst39dc58T
VFamLBk1VJZuKPM+QNQqhKx9JpxHqJW1nsoesUmpIv9MUehmQtHTs3E28RrQJ9tzOrcjl6s5ggOr
x++9CfA1aq0fuppECAlQ38CMXFEIt8wLLk30z8irY6NMsdqKUX1x0RhUMFFJUE3FEGw0zzpJ7nsW
erVsOZa+cCf3FmJivaQWZb9teNFiW50ILzkmTvqBeamn5m/N2FkiZgxGQNrKsgvqPmXOL433j8aV
njKJ/JXa4Z+1rManqWVxV7DbzTNMuHC7TEgvgqlq3oULQ0hPB7Xv+ASMuoufjJC9lsVzqxB9jwuw
czySQHwWrgpvFfpL1BOqLpuW/6qKeQ3ByRU8wwX0lT8jBn2sbEg1QzjqWZ/fR/bmHhHq42+362td
fDLUp6DeI/ToBC+U9dcG2nEPW1RaqE7Qqm7LAwJ7BMeZ8RbaCSydOBfj6zcKfot2NxMIBVHZNr84
rRV314VWiEIJvXOkX330D72g+CmuOLq6Zqs9vFcHmSSDnXMCvK1ibfKMliJngRjwYNyAilxSWRRk
EQrk9uEXM9nl8H6xNvkmgHb6+h1z4UcGFflbzLa3KK7i7h9He0PF5pSwU6ip3af48nPOPlZp0CMz
aloUQw5nef6qo4BSJ279hF1yhTUjIB4NWfRxNr4+J6Pa1brdAnYydW8c8RHGlBN+EXto7+M13c9t
evcBO3IdJoWllTWi5f7+irOSDYViXsP7OwJ7Axwno1IXsJ2y8cIuwJkVXud3jgASE43aMteeFFKQ
Y27KYT1HNJX4ghjbs3VYzJ7ipr5hkyU/7yQWSKZj7HYdBzlBA6DcxGWb9PGoS5bNr0JTSpsXJ3NU
RD9gr1zthWUh2/AyZPusaKgRKmaLQ132IgZzQq94gcmxrLmT1nKzQUi6ruIZ3wJAleaNHgC7Upof
E8U5ueOeQYZM9iuAUlFS/qp7L13cFXmJqlZru5I5toR3SJVeCJEQYB8+q0gPB9KIpLVBysgeYr20
uTGO0c8SloV0drCyiROFqeHfowRCf0Ud2oIWCbif9DldmOE5mpK3gvGOmoBGFEV8ZQdsRF1T00p8
MISatHAzz7wiXYkBdG0KXXmAFPg/ko+5J57EKvnybJRcY77PLOzMjct0apsXWxPrllgmJTHeNmRL
FrPbyWLDNSDTA5L0T5l0warkWh9zKfZ8f11smHxxPjEiL/zRuL3qF7S9/2F0NHRF+qHo1W7clGHr
LSsnMyiItINpcL29DcZHdXi5n9IH/gAAiC/y1pC5eC4bpaqSETrs1hzKVz3dRKu16N6UGtUznbQP
iEaNLGaVpULEuwYT9i8T/D/QlxnnNalaU6Jc4LXqbHVKD0zw4jFfMbkAxePbiL1x1gJ2HOCVyjgQ
6KEN5qv7pOq48hJvfyDJigzaLVMZQ2YYG4VR7ZXCOPeueaUVTuxzjnTbEeNe8/f0AtbiVpdwjJqS
NP2/zWgvneD69Du65ZQck6Ta4zYf6L1a0nKhyixTVv2HqQaV5AnUpLIOFpSam86DLiHXeZGTFhJ6
UoO4SA9brl6wsKAzgznudx2kVe9361RPjtI6vtk8C3K3ONX8ZSr5E/aWEXB3M8RJdkd86nklAl+w
gJLFV2t76vv5BRxC18clgTivuv6hMrdr3YDzEUAHAHAs+dmsr03zppP9T+v9S0CLBSMzfnbCWAL1
HRYVNP62SWzFQflbWr+pZsBLfvE6j+NyiGl1FJVjdPHH/StYx4fkvkZB2bWNffnfCOfmVpq+fLEM
immv4+5y6/YM+mLuHGxmD9QoBvTTlfNtqxeZA/Zc/SIhuyHTPZBjmU84jW9YchI8kpXCJVs7XWGt
7GOSv+Z5XeaEVvLwN1bRkZ0CnLZSxYs8+XGKqEl9gK+YTXWZNf8Z8/Ps7EOGsrDAv/LJGW+89Ulu
ROqzV7fYb6tGXrN/fqEL/96YAWDh89Fmj9NOnkJUsD8FsvjEc4l1atDu7VL/RaQQz8R5rIztXVZw
v9LEXcB2FQRL+D2Yey/3+b2a73DjCPoo2/L+6Z7XizTd5zyLJDt4ddPXYXuClw7I7gydLA5dfPFF
BvxiZwHzwHQxOlkewJNAgyxYwSwUNshvxHbxWb5bw+J1wKYFX51QTVHHWivQ3Q0mEcB43NbQ2Ets
yxhQnRlqPtWDVJBDohak4WF8wFUVWmCPcR9aQrUUy0onx4+4W/thhAgBVleVaSVQDwLl3GrNPe0y
fZb+fRJiewaiVn1DUgaQAF+2NZSGe+7YmhCO1UYW1ZpobaIA+7Yl01tEfFqL8dyemUp5rA2GA9+X
/8PP4KMau/vRE4/L8AsGfO5vwGfpj+oNclvPAkIOJTxfl8eRwXIIcxdp4Pk/xcYxeTWAbyD7mJUl
h5FMMRwMbNwqJcQ3VY3rX47ME0dm36ocBJwIRiqTNDYoUDwkxGnSZcOPZ9MtSjITe67m9ZW2wmZp
3ZnVe+z7ho8xKDz1MVKNT2Lc5H8fJS2JRzxbKk5Y5IdVDoOTf9CaQlX0kjSzvwtXH9TvL95+LBlA
CpFkOOLHmtKB+K0IVFzmorv2wqK8LHd9y/4556IdILdM7jNjcOYOeYnvP0vDD5TllBNQtAUL6P/k
ucE6CxFSGMcA1DJhG9PV2iNMKJZ1oR5gzDZ1/N9XTjZOZBs744tuIC7nR+8TymG2T4jMwvjkgFfp
qrez+uSCpqh1jucpU4LLZf+59pDdPQxejQuaY3FEXfHjXWqWLA4LI1l//fOjj3OgtJrrV0/mADfZ
VmxiY7k1akau0Auspfk/euZlvL6azuKUFpBF5368dBVeK69Xx8eBVricTQsvPl4+ehZvvBMBgAfh
aNy4b85PUM++qD9Yw9ZOmqXEP9QasoTlD9FZhrDjo3ADBy4O76xg9R0JBbS8YmWkYpOGZxVnQKST
HfxeNuFiD+z/H05RyzQlQxA3rHOmJDk8nD3Yvo6BSVjTRvZA2VR2dV10TnChonqASI7lDq3osdp6
U7NTdeF43VAKinP+21rTTKnX16ACC3a8jGAK4JdPAsWu666DNlQ6D1RoTiXX3eTaecqe68PoxvKs
kSnM4pNxQdv1kTT08M18txI3QiXa+C23vJXHpp8iDciCd18szzi54c9Jsq96an0g7Wg/C4kqsv1/
PL3XBuZ3h6E971zwq5NSfVPy9+2IOzvketHMoJNcgYNk61GOCy4xMD1pAW/+QRWvsZSo0+06T/16
W/Tsn9fImMwOxk6K2N8hgfpxrIP/Ge3UdM7RP7Pn/dfB2p5QeAzQmAmi2wz9znbTVeCD/gv5/4KJ
z7BBMW3zYRnm5r2IPZ00xYcAD7vtvF/+xH/3jROzZOi5UkO7PjtUNeOyszdeqNtmI2ZYKglK+jVe
tkrzciM4PIjnNUDH6sjNmU+U0sC2hw7CRdf85Orm9alxlHWjRJiaoc7DedwlNFs9w10Jb/fH51jm
/Rzxw5jEyz1xV9uZwBq3euaJ2H3GQ8ndm578KmAa30A/KRWXGRKGYeEbYsWrMQ3FueWQVleT3TIC
I4SN9GCScavb1+ft6P7r1sI9ln/tn1ypse+gofkvMlFKhZJqw/aCWe1gzH7x3ROPXUZPfthmi2li
c0Wf67U/T0HKLCdPDMG98JkfQStUeufo6cErpQ66t3ZaaWphd2QPQEItPib+qmNCVlDjvr45MKJ+
2gdZOWGUkKDrXHjvMyPV7DgbDoCfiQ2hqJ9GRMWbDOn4wOYlwmQTyFHDBLZ4S1nW82yEl0MBL/6j
SCzfFb1uWY4G2GOSh7wB/gSmqLlX4TikWc9g1B4RVv0uKEo+2Vf/rCsRhLt1A9Sh8WAnMaowapns
/mxGTcWy1CvLWqpHxN06NfAaKMk7GBQ1JMnmemYDwwKmbiwk6iYtFhjp/65P2hFSXO/MAY+I9dPA
6GuGQe2euLLb4uCUO8Yxow5J4VcHH3IaWRKP6VR1i7PWnIqeZY//eosh1l6XLQFkPioJwzYtCQBz
sLFichSupc4iZn+xc+vWSiz97HfBV+h3U10UmslimZm5wJBOpIGnR8Kl8QAPjmEjK0mZCYs3frUf
7M2XmD4nATcXyn2XXHhXdzt+lw+oYIa0touHaFifamSno+6MF39f1WDzK40rN1bNOQHdKNQVTga2
NGNx3dY2wvtUhRSKJFFNywC1/WhA98eZFY4csl/o6PDSXZG5HQEpEneeNlCy2jcoNicSBUokYd8k
pDMw/dOFx7cTPSUWcKoP6wHiKtrUp13aiIOPyqtWGwOv8EKQkmqUxaNSaqfKiZ2SbGy3g/7PGyKz
LnxzO4CSy1FPTBsBHGXO5lpjLNPVrG8Qul9pP/h4iLlGxK7Sa//poNp2ULEz5ZFoUQMfFuUnR1Af
fiPHqFcsPZFIEqaF+IeZebfOOjTcvODLdHyzJXRn12vuFOUICIvEHkm3cA8aJwWt3YhAnRQIBtwA
QOornh8R7GvquMjZ8+GRFGdCrr/+rYl86xSqLG4aiuZIl/NcaOM6VuwhLvQHkUVkKpub3brZGWtu
Hk8BcQKos8ypCdLk29wb4iDZj2lENRvdc4Wyij3sqZ/KkBo7zqsyTkcbP/e6jSFcBpz/ZrMZnlhU
rA6+5A1caCIBtLMZKdLxPOqMqyIM26B0QbK0WodezXjgH41u+DKLfMl2CcVUTdBNFMfeFc0t81Lz
4XiawEODgJ4j0+MAaN3MydoLAYLVYwAHZXKd5n2JPLvnkKtw38/OYwmRx2BbjI4y3VR1WAEwwaE1
KhVsrQOUkAQnSbNbB5ZQByyNHAn4PY/frCN0ic+bImH5xi+7UadcsRVv41/T+VfZ/KvOMBLMZ9Wf
nqclMmsDIKNsKaenaa43GcXHtJCgs5M+FnwAznH4i4V2vYC8QHRCnw1pC3zf5RVo31rjOzkQulrB
yyIWqm3rmoKXTZ7wd+lMRFCbJO4N0/PYnPCMMVeLvVprS3Q3afSbxeXQEjSI7Tnjxb0m0Kub4B7E
qluXVqzRmbG2zmXMZQ9FXJL3rrEG20GWUaMBgzMh1yq3IphhQr+PwPpuXUGTIhX+pitIXHpNr5fm
szCPbl459jM4lhbH++bTnu8UgqJ4CSW77EFtObNVfzysnGRliaLx1lpfh2qxRTBCDzlVnLHBX2fd
km3L1ob6qkprfjFmh6YHQ2WuBmDO9HxWQ3BnhW+xF2bnMdGgaMEXWdY5TRs8/1kueFS4P4bcjJLj
oIbnqiWr8Wr5/1lkV8dBBDi2bZNusUTfZc3av8aCtHxk8rATWraz/22YZ3b/pIbY6e+Yw4FZE8jB
MTKQkGbRadbdN+duVtbfCGGMJupfFK+xdhGSh/419gMe87C5g/oEp9NIeNQEq4uP6WuRUK1WuinD
zQ3g12YoxR3wOCnu50DK+lVZmhrAxgnuvDhfkxhN+D7Se+zc1RdKzHnxQIc0pzLQ8YXFG8uj6pQ0
5aZQ/OuFrAy1LVqDtBX6bDqk/FiufdawuZu1WRhWD7K+N2kEx11gOuJPy/7pSaZZPkF8mWr0GJO+
IU66AiJEKykAJV8F6dPPKoUcQOlMvZHtGznDc77fbA1xYJbJ8Ms1nNjl/RE2BiA1Do7k8w/uKfgn
dfrDUfuODyfMHmi+EH78gyELfzkrjvQ3bk3GOV/9CxoQko8i6nRioDkIJ/29zVsJ4TYxGmgVIkFW
/hu/lb1vHWZ8Ffwz/at2rzR14kaxKu8BzE2t8PpQTuiKSyiZvGR+tUfQSuTSRZ4/B/R95AQp2hPp
mLHXBAUJif9tCBSoBLfyR6sA8yp88B5HBurmVjVu4AMKKbxKOtzjd9bwI5u+0qnsMspOU195VDGf
laC/ezasH/VRINnf1fHUYYwvDeER5uEeDqeiD0tCboVoXW51J1rchbMuw0dik8GBB+cv7vU/Pt/u
sqYh2HpJ2BzrggI+E5VDrptcjKFaRVdZ8jIsM4QvT1Wb3ER7Ssv/Jcnj9UJZ9EBpkj8q940ZZTy6
T7gY/jrNU9iK+W6tOyFlA+B9c2lUoR7CZkDrDBlBhBSubsNQKCtV1dRk2J2LM6d0efOB91vIwy1H
jVdvxA9yAPosIhGd1UbEMn6l7wKMrlPNDDx74SIy8NkIy+gNGyYDosG8uj87hAy6v9NEr/EPvxuh
tI/hV6gI8NBsaqajf78ccfSxOFDz+QNcY3/SpyRMzEWyOW9N7IPriJUglBdv8xj5fY+p0ePVIFv9
l+bmZWUz+Gg+ZbmnoRbBMK8WL+lpiG81CNsvAN0XnnScmYcGZ9JxG88QEUtvGrjaGTv1fA4cQPC1
mL2thBLo3hEdF7RxAjklUCBA5wIIN+zAcFl2Ej6xVuCgYvQHvMpREY14TP8+yBDwTrfIiFV7xD+y
G9eio+gjqT5gWnC4IVFuL2G+i+F9yKdOjTDMDH4WqWbTWfNNefeJuk2AAfFfaROcCrfa6/KCCk7k
cxgyL2tchqeZHpQ2MSXvbjsAigdLdVy60L/v5FJZvzEW7kpPXBqHFCubQU/V1OChyVQL0HZEk/X6
WvVhOsC/Lq+yKsrXu2CZuh/DXQUxYmrgxaOy7nbAOsGth8WUYoxaeBoDDnZTMvW23rKOEk0IfzQQ
RZBE6xu9sCWhLl6eC/IChh3QyfcqYrUqzsjozMKCTupB8bPrclWSoHNZQjLXJpRmgcl54joPjOKQ
fN/EqWP7P87iZYY3iTrNRsrSEl6dKC/T7rDYcvM8eMHzVYN1bm2EsmzUN4E+eelzoJ6A0cVKyjqJ
unMVCoo8ho+u58unj2YAP9QrOPwR8sWK30fUSGZUMAJeIBeTPjio+pTeUckNvKYgODBTtOPAz/CY
cuvo7kFIJx2DFc8wr8BOFE5Z2Kyqub4WH0LMUWJ3Ki1f29MGh/DFz0I0P/8b8elaHDCLL4SmMOLP
XeUMyBss9LGGCN8Lf1wByfwxBfry558cNZIJB/PZy0MqLrZcllY3WcaokvZdMMCo8xHqvpu74zDV
aqyrqw+oUquJVUdkp/TLgL59E/uLDq7mr3ShGtdmTmK+1ET8L0gB9SrH919a0ESKz9olZFKXGr4h
6mg4XvH0pK7P/PSw3BRJ6OJLb3mXUXJ7bdKvfIQPJfzd3o8f7LRFlWBw1WABF1+zFTIBIvVOZeNQ
eUT4VxPG7fk/ZNVCwoJVXsIIw1znBlvFguEP/8IR6mloSsASZa84r05hbBmKv799Xqzb5zzDyM/c
vBIFP91m1yuWsb1JTyvjGVkehlUFS8fM02+Qgh/P7uKLbzSgqVyLPcK4MU+BsAbu6AFn6TyU0bUu
o3fKtemkTfe2iF04OjVMdBMgmhd4nVVasq1EimpkNl7eEQwhAh91YCEfYBKz8bhPin7KzvhKmaxl
j5f2Sc+B9LMOGcLdxhva4ZyAlM10mMjpBJLwy1AVk1U6/08JUZpBivmhkNjcd3f0Xsw+DiF3N8mM
gIBFuRTp8fRy3rAHhCqOyaZ+OHsySzHTYL8dTkqSXbIr4zbfDARPRiRZXOPMF5xW2YmLxow2sAp/
aY4D16Ot4fT8aa6FellQTWLx6jlD6dyO4vGSUFb7WWKJAZ/nX9KxpEbRHyaAhBn4I+xnqjmodzJ6
Q8cflhSaPAq2NfuNl1GCDaS7S9P3Eyk1GLhwcFH2YOcimiZ1LfeSYbMHTSxmc0JeGrPFFcDIQBNQ
cAXarD3WOoE7Be9/P4nFiTvKmh/UtPfO/H/0hofIJRvuzTTLniJBwThGy6PP+sI0NMA/K56nlhsX
XKyP6OEEMac8VadpFD2TuCsGTcAE0p+VNm/tOv0wT38S3GkPFZSyr0eudnXko6WS21O9jFUd1J5q
NjKMNil0u7+Y5VFONgL9XDm8WKcrrOcAE4+/z5So7bCNiDOpu7fvFtaNFGIfHBJf4oW4j56wA0yu
6LA5iuJOS8yV+REXNjvy09XHy2O9hvyOVhWN+eQIJ1bywdfl1HhyuE1tnXnAQvxDVKdrfFZM5tXf
gsdjb567iOXPTTOZl1D4ECeUbxp5N1QMB6SB0ky9AZScD6huTG6xdb7mcLOK5dkei8Ekx8NJVx1Z
7ylkC6pzIGJRi+wwQM1/AEi5zBZgXdJl9k3R0kOmZYe43tHZt7MJB4vvda2CliFSQwTO1GeYwXvF
rlzE/FZL0ypA9vpP6PEWMfude2wSWo7aqwMioi3pzYz5GmFYWIDYicSJM180GrxRcvNd7TjLnFO7
b/Vqmz1/Ml+7i9g8ZZQZkUWpwkVtD4VsNYK95fruguXHxNV87sY408EJY+VMt5+IdlnqR5FScjMs
WXiuyKI/hoCwZYZkNXFBJj+AjOEREBfSAXkHDgppEoL0lmXKix6Yz+bWEln6Gyq9i14oVoWtJ2Lp
hasFzXu44IntVxUysHy/pmj1opPVsd4k1ilIySa4o+/nRdZTOCsUB6EE+8FctaPmCrGdzBl3R+ih
oizAME9kokBCmWVyjnYjSHW0Lbzct9aTokHeivL241IsVDVzQCt2xP1RJpRtzkgCyVSKqeogLdBg
TubNLG6CnCBh7FRldVsF6hpJP+P1rZG/KpK5x9nNxbb4swSN9sD11r+PVJ99Jrv5MdE+6O/71dBx
7wHFJ9dDLSxB3/RocdfP/owu4fgDghXrl4ZCivpkTg51pUEQl4EbdXaRlPE19X26Pv1A514LvOOE
8luv2pNSfMw8bxMZjZj76bByo2oUpd+LQRqlNbDoVWhcSJbrVlY2HkQ2mAM9BoC4d7jBolK7PUiz
akK95DSwHZzYQfPaLhJFxRTT9LNGIQgjlE8hWzBggxToaGSES7lellR7zzNycgYqIm49m9y318aC
eZnwO1IKns+vuTetMI3GKY/1hlbRa9eXELqUXPABqWRWYF1VvSIeKefU7KNYOibTZjqD8ytA1DS8
DHJT2iTePMsqD18wujumxf3KJP+q3jm47fm2WLyCcqLLccHh+cOfBoBIt5i/+oe7bZjjajv4jZHm
UZc+5ZvfHUqjJaeBF5cRI+96SOhOmFg0X3svcCTTsV8YUs6nlR3v5Ls+BB5E+1xGKPvpl1hx9Sow
IialARebwN9z5A+69c6dko5h+QPqg1HiiZ5dEPH8W3CdkCeruOC7+PSB3BaDF/jHOzcUScAywCh9
9u4zVpkAFmwpPkOfPpLMw/TXSIX06Ac89d/ECIXzBBSN+2ocWXnQ5zGxS8M0FvkfE7MoQheNcY4r
KMRN2WWxeY2hfYrKM46FZlhhO0cs8Ejy3yKOUMo7Iwa6zG2drE+yqphyISHvXQlZB8UMDciy+5Dz
9OKB5NdLxFOu6Od8KqtVyyoi1cT/ZawX65rT6YFq3BwGqFRkr+nSz+RJwo5byayKVc8J21Y4wLNL
fRFbv7YcS267vx1KZ1XBacQO+B8x8nJ1JrCvMTppSpV488xki9VhTnvkkXx+5Lnlg7Bi+wRPLirz
G7dLBeT3VdD4qr8AQM3Gc9yo8FyXLhIg6qJOBCuidVXg7jhVrCFrJwWB7cBjEMXaZuVvNv01JrO9
yoERkIlb6bgONG9D+0MiW78mWM9ELidOBO1tkUTgH5orwrGMFIsI07nBH0/r6Lq2g8FA5cgCE1uy
XoMaKzvfY1oHVLH198CbS1NupEB6NwKgOo0aLtUqvo14gso0wS1P8Bfn6ysubiK+F7lynQg1uo0d
oKQbbTD1QTw1zNuyfT8MvD3b84un/qA9pQQYz4v8LkiY7e+biTDGia/wjzzdZV3EFzrSNHleqarj
VEmdgLOfi5pygBJW/yapA2GHBeZ+JccVgKO966DutcntFmp7Ylwt5FPGwewPT6CRQeCv51Sl+ana
2FQF5KMF1i/Hl6ya3AkC8T908IWpnvtuAGJ4lbabpU57Ti2317TnvPyHuxX3k3OrhshKXRm5kobi
foUDKhiY2m9ZUcoiQRRb6LPOCiFMrR+VGqd6eW03eY6i0j2d6iLylV+SNMB1kzUspZ5pShrufAIu
2sHmVnYvVi6x17ksR4b2iA8/CtP69sIqOj+UtIF74FY5jdHP5pfFkCzDpYD5QF0xSu7PUrjuoIbL
X5r+TJAaw8p/gN+Fmy+TAYJLGaOH5l1kS9rpdwNta9B5Vgq/ocHnSnGIO/NZJp4w+IQi8dArOXfd
Bi6GAnur2HZ7YeupJhA9P4ZZEXn3gSKaOQznE+rvoZPynpp7IzVxbzS8OdJgzAuiCaPbEt8QCoGR
5a/iC66vF+rxEHASXipvLGQl/B5APG4+57rM6cOkqA2FJQ6XSGGIRp+vZsIlb72VVvcu16TMy9zq
oV6kdIWDX99jC3x05FFVBqN1hB8v1HH5/VCTXV2vbWkyTiwXFuXTAKnv1hvfwifxLq0Wjnh9jisg
MHidAG3OwD9k87w2VKT/cpMUqSva0GRmOIUISvtPGCufWWQzjiOP1cbIEvwf3S8AAqxO0Hv8sP/v
QbiPm5WkNlatzewbG+odb68dVZ3wYAsecwoYIxSOK15BSgSSlnHZeNmaZkqI1bpg1fMfKeSKJCTt
OKqMEbiIazQc+4mSjaLmHpjT8fyJWpBguxAma9dKOrVASNpa8YBk6bsw7Bk03ld/4nGLSibovXcu
3Kk8eKYwZ8waquTI5oiHwivH2XfcuILTFQoz1JCCajcA16hoJ2B0gZ/Ixp7YDgt8/VZlkJkorIOA
+F4fm/y3MJ/LY/IzHRzpNbPLfX/1qZYqYhPkJcBa5VsmH7poAgetf0cm4ilrhayxesGZbkZsLV29
ZEhAJ3T2WUlQu3jRDYNLAbusqFx8gM9rjEsKGoNzC/ZWKOSQMmcO1m6jNjsGUQdBGTTOEDINyHv3
W9DtcDVbPlu4GxfAmbem5VxuT+Z0mpZAA0qRF9CvRHuHBAJiwP9lKcwMZYKjI5kch9YlkDuYy3AT
ddknAPb+xNM9OD2aWGBSCE9B6RnT3OB7IH+gN7EbRJpwQPCicoAv8h2nMPWuDPbrq4XnLjdmtNWR
LtIvms9QfYJvQ6DIsu9huwfz4raRFyR34/kyWyLMilmQ1cVI5mdSQtyLj2hGhbv+p3rdnzxg0jGd
VIAeszz57O/3dltWEDr6uACZ1NYWtAADbXLv4CnYPwXcxkNeVyHNwWRMwXng3jYqDZog8qDRBZjz
r5xL3NEKRE3eHT4NsxCKexKcHxdiF8MGx8dhveV1Y9A3sE05aqH2RIgEorLGc+BXNge5n6Q3rcd5
oXN8Gk20PEr0J9uG9rSCbI0qErjMsvSXEcnk0jcE9+8JJaMG81CzhH5aSEKF15iTDNz8LXvxgupk
t21ycNT2uGzxK5l0oDQ7KJP66HHM0Ril/tOW4Gz5LYgHcCbC68mOWw+y0KCggSdBCPAUsy9J6Nuv
59w4b4vj22T/J0EA00OPezXMFd4Yl1sKblBVGYs+77zdBiDcTr/nGbhKxpbNTqC/u/zpqMqHLcL1
87MDGpoXSNFP9lgcMunKAotc2y7nitZsOVs5XrkUNeLtrYZwg71OwQc8p2EKkQ/c8I/DSukRp64j
zGODRhc6WabfD9Z08P3+DUK1NTAilQ0MSgZsktPpqIzD+CqwZZ2ftWa8DgmVRBLXsPZYblW0iDrx
ANLeBUfW2iycHKzjDfM8u9wgQJ1BY/qazHzkOUY+imQyoe6UMi09zb1fL08hu9YQqGspGxBZCd85
pdrnMSiWXRM04HrrHntRqcr6S9CdtuF9cPKJquYuEXj1nsWa+qflDC2jokN9dqOHDZdAhI0zWqA8
dueJcAm+uFaXP3oFal19LbaMQuOn1alPS+qNFjdGaV0+RTHIdpOPgCgHeg8N1j2caXtD8J6bIm8X
G+LJf4p0MLknmJXGoX8Tam3Yaq/TNwfbigliJbQ+njL3xBSQl3A+HXIoW1CfCtzeuw0ZynYrVbsy
qSPvCjMDCLG5CxavqV6iONbQtXp3EYiNHQ4hv3JohlIEjEDIRrl4ggyigFa1piuNcx8e8UEUPE0f
xVxAwDOf1zj3+sPTFd4I+GNcs5FHGwztK05tZv4+Q6/jfx2dwZGCaNbwacQF0PtzlP8ZWKYYb6zY
Gk/CR1e3csVGrtGNk2cW0Fw49sykqAzygCcnANspHzomyo0D/YdeIHLBMq1L7SHhergfQH0uZ3l9
o8qihLbt4nTU7Z0tXeHg7QE//nX49zZhd3aMucugStJWEv3BBzeC/KW7yldjXcj3yP26NhHyO3CH
B5865aXs3W6i+Riohb4HCbpT1zg90OER9sBsymJs+Zadw8Jt+N8DWPcyNlLogA9nTLzqAZqIR2SC
ASNCtWHHaONN4Krvi+KDntPb/w1wK4wwhE39BHEcezYn7bJSB8eE0TDg6YLd2J5vxLmHa+IMJcRY
pR2IsrTTOyuV7hFxKEY1Jt2994D0fqD/YQYRY2hBWxk2HRtJWx6Y061BOn9nCIxfgxgj/+GHUngk
UsA8XIh9tAMrhwC6889dr0nizD4PGZD0akExyyMDJbLSYUtZa2pIKoDOe7PsqGwXbnGYCLNRWz4G
L33x0Fvr2m5D96fHQ9QNi9GJlU9saSF++7FWpCTpv133tnwsa5AVMmIKtjkgW+obrfLtCkrxPcsq
mWAR8MsjF7DGX4BPRzT+v+MdiafiXAYNQKPCB+BGelmhGEwGFYrA9qrodc8uN0Rqy8+Rp6IkQ/IC
Pk/ZwOk0FHAw5MDB7YozvP/NEeFlH0SSLFqvBWtMOKQ+bZsxcPRSwd6J1vbuRsCBF7/IczaQOZWE
kvjM6iKTOr9c3xCVnE9LptIZqSGFpykonpEudeD49HX1QhtI9N1XugzqqWSEM0p7MX2yi1etCSVK
Zd6KJerLiypzxHJ+YIMUlhKuVbjrWDjTivOt4EPBUpWDVvNL26AwmJkYAcagRTkz0l9KQUhXKXa8
x8hwC2N+kYXqpyP+FERnLs8OYl6dZykTmxuadKx9yaf61zDvgg6U4abryDFKdbzm2RUJGDC3VWRB
titYYqc1blF6ZY3q2Jdb/pXFnQOumCnb4kfxS3WDzG8KV3VF7llSmMJszOvN5OuUsI2z6MjyOaD3
tLhl47b98Rtl9fC+BUtjRlM9bck0Q9nwLWb1AgSYTPgEmxST2LoyW59mhkoYcbMotYeN01sXVE1H
XwLw4iJRwU3CJDofogaM8JJv7WY5KQYRcLcP/pOoop/GRfYTUpqFNQ+G+elA6asDEMdbLYaVMfHo
A0K3L1DZM5zs7C/qqnMM2Nn9QtR21R3Yhy2C/gzGKGeYM5zF+nkhvS1z9npyBqMNy5CbwsBiuFIh
FKTEB3a/zr6T6u9mZ+3Z/Qsycb7K0VNOANhSsOkDDe7+ol6H02YEtY95At/QLjURVaDXgcL6YFgc
MBXv6q+ggt8Y82kIXsbtTSFLPilanCTTVoHaTzEC3B1+OBrBxlhgloU9bK2V4m7XunBpF0SEAG1o
f5jE/9+rgMy3bXSX9YLDoOvUCnt8/5Gwm1KhhPMN5PuOlZ3ESts4IQti22AwDMsgzmJnIBEf2mmh
96E6TZPOmR2Bh5LsaE83sb97bln7hLptzK5tT8ECJ/wYeRVM2GrHdvfKZEcfCscSuL4RLT4TbdKg
8MNYXFpDydAVx29q7Y5fz/jqRVoN3JzRdAS4JTobSy/9Nwn1/efqbbzQAI6/9Ux45u0ICnCXr9i7
fz6M6obKnGBvRziiPt/AKYlTRqpqMQuSXUus9cN5SIs6qMOO1rpWfyFvxzFrFULSb5ZOG1EuZyFU
9so3jpAFGLNZ5wbWCkyeYfyPiT3B0fpCS6HlRVgDHlVaHHkguJ/tP9fwla1EppZ9X/vCyvgCNqoV
YwVqGdGWSCo2kVOLObl2twSaOqTtCURpUEJ7UT6N/CIA4HA4gEedv2SwJwFnwpv73DOdHj5KMNfM
N+fnUTruqJGIZDP+EDX9rqU0z58mG0ozSuGpMxqCLMlfozXf6mTRpIVGdjMSMePaI/0ocdP8gaPs
7mi2hOUkKYZB3zvlYOxhmkg7ZFkdJk3M2tMFMEv5ZI8HfJC35VP5CyZTZvciDD22BF25eCEstj7D
WnA0uBKYdngUFGnwsQjgZKRZ4eGno91ui7KlQJbiAS6HZzdqbzWDB2VioWl8pteDdZNOEIjDgj36
irW4RSlrTncKCZoig1k3IO9MJ+TS7ILB3PrH1igIzNaNGMVjKX04lYL9w86RXnehVcOslt/bIMRc
snel/JxxVsfxFZLUtrZ91htro4Ww2pAHdwxFds5Y2DcCLSG08M5hgxJyzC1dZuN/cCP5aJokwioL
kfmrhwk9Sei433FmiV8JxBLKJs0qnX2sLld/IqPB/w0R413eNwW4R3qymmL/wZC3+SJubH1n6yoM
G1YxHdqqa2js7MfklTkj5eRMl6yygjSkCTZdBd0bxLxov7G2aNYc4e+5tlwxHw+AJOH8N0xNK+mO
zJXrvUD6EaDytupo+M0H5zbgvhW9YZirMbyADXrbU8YDjmlVhm2KAkPVELaNpc3G7itHEi5Cikku
nVSuftuPpQOVAp7Z7M8rNXg7nBJkLMRKqyBWVxtsEsTLC+jw/0fZES6So+otw3VPXKMDAXVFkDC8
sr8Y9/A5sHLUd9vAN0YqBK2ddUQ2xOAj3MUcbZfLbCdtk0eujgtMnRKVbdWQJkVQd/hNSH83QYpc
XJ7RQJF7LyqyD5o4rpDJ4N+5Qo8qYZRPN5TyicaZNiG/6CrRG2ExIbXA1uynTsAGN5530dumFni3
9Kne+Qjo9JV1sFekQA7y45S59Fuy13mo0fDfyK9HGLgdPZYzBeqzC1qsEgZ+EcoygGVr6e6ddBMF
k0wfLOtVJRXgkY54PMcZT9nfiiAGyJeiStiXGHbdFPHpwz0gI2nDh1pW0WtkTCAWVCpXqtJAzuKL
cZ5TGYoxGPnZXGe2jkhp9Kky1kUppWvYTIwziVskuB52lp+1T5T6wl/eZwPiotz0ybSP+HelmTBP
lUMaWaj4mIbIKmCXd/HbmYk23byL3f5gDCA5gNoacUGwekGiu4hQxyd9rU7+rDRXbhkbKWEKS1ch
oYgyhJxYcEJmEM7SOEjTpFlJb/GvTZanEeZE9oxyA8R0CrukPSdZVSitSBSFeppt+2c5+LBtbft9
xD8THVnB6hKJAW1veE+7fBQimw+F6fgFiKreOl1T+JlhRUlAmGG2eWQZCtxP3qcSJ+ksDVjrPsPR
WGcwOxOxMiW39tjJRtaoTwgsIfxbfLShPdK1IIjTFBu80/00cXNLeu+Oo1JM6JqfxL2NmEHwjUTm
XY0QdClqP+aSOoGl3WIUTUYn/t3sRYi/EsOD6Mn50hID4Z/TXZ50buOL7JRJcKc9PLX8RquM9szp
27bnMcBU/tLqL7H8IS3uKAcgKi2zZQ2DIrytXJkcAJm5rBmU88vB7k5hlZRwTL+ATL2aLWWHR1OT
U8BxGtvOtHd9NreU8f6e33/4hxQ4GLjHbf6N7CWWOZFxFphQlvJA+rqHj0NFxti6L7eUZAr//Wc8
5RBAuPZCf2PO3bPHEO9sj/ufyvSKJc9tmcaAu2HWDYWpJJmJpjSPwg9sjwhIhdP4hTaWuSK6W34x
KjYNkHmjWUvUPeCOH8FVs7GFOiCC+UaCUXx/LELsEvsCoaujlAH6Y7iHdJQR4T3z40CYKLodqFc4
SUkZQuoo9lJzaLs6d2cb4rZl4/NaeymQv5YpXQN2O6Z4SA45n+TzU3i55h1pQbSDy7EugtY2t851
1mGccrpnmMQ5ZiH27COmM2QVcDp8RRHJEj+H0FrcCdmDPoUGR59dtcuF7Qam3IWDDC/YAX2E9BZP
zZEbjzw8LFDCYou8YsIsfHgQQUfBnqntL2DwfB64wMyoKtOHrL5pi9Oa5lWehGH3CHgKy2LCISQK
2P3DVtiJD6Zf5+jZuQmEeWTZV8j1XY/R52DYxzf8tSqUbUE7Wp9zpJQiFzLPdgbUkrWEGY/7BKGI
Z6pSNnDlNqd2YxRbE+9Kq1B+jbfzS2TMrDZjAfx18txBCNX5vNd/zpaAA7roCKXbHSEcHo4MefgP
eYxboz5S0GkWl8IHJEx8gEb7Ex7ew+uCJ7bNaMdOv4C6V67mzjOfVob69MqORqw485aem2LdwqnW
e1Dv6o+sfDP8lDkGywG28/BvfT05bqyWj0RrjTOno9WQX5eOHiwW5wtKNFfQC0MGQL4PVsobUoKw
3MMKBoUf9Wd+qyqoKJDkrcQmbe/Erb5gaj2zBrKKyW0lBVxmJjrE8IVC3JemG7BcOkDhzQEbMqg+
GLpnWDhScAopQ/Gye7lhZXhWMWvNjd9UCHwDXcWhi2O+qinEY+prLB6AuyrxktXsa6dwAon1gShQ
bwTqvlwlePbmi55tPc/ZBe6WKkNN1L9u0dwbKHcGrMeTBRRkwU3J8+ZmG5k0bmYHydE0tp3aCRcX
YLc/FAJveeEYJaVSrUVFZAF7yaRPzceI0cUkaEWQLAGQMJCpyh08ah9xgdu0FIf4aRwmuNTX18ky
ZNp5f6JpyHh/nq/VSNHLgQoqzbp0Q3oLYgpQKfR/vd0ZuzXGACbRBLtPQiKRBvHmYdqkmDA3Jx62
oxeWgRxa2Eh8f8KI+R9TSWZ1g/TSHvzK/PmsfU2fboQqwUL5DiadnNnz/E1oD5iHaM1+2ERbSA6g
6BsV3fjCkDRsvhfBZVKXWF9Zg2VfyUSb+kg0Y+4mfkoX8g9SNEq3EGk3AfL28v2fl0Pu1UNKTr76
PhS9MjM3NCS1ePerY+Nml3n/J+34Ci3NhpcHddw57EFOJ+b+3523Kv+n0U2+SFtTqippscJP9Ary
XdY7dyBwMhaLblEqOh+/XjaRBk3Fwo6ZYY0bmNWfhC34o7l//Yfggp+t5apmK+wTIpgivol/ihtp
1th7xckI0JzWB18TmXTGGw2fyL2X3pDqFKpXqn6FS3pKUqaLfqxBO8jB2lUs/6qImBUFxQBaML+X
TuG1T0BUJH8+OzlJy3icKgb5hakyDYlgY+aF2Yrioj7XxTx5OAk9fM1cXakANMhHdrNlLOSDJnTw
d/lMQrUNaLeLDCrzUM9dGgCJABbP0Nz9wNPY+pkJaqbJ5/xaCD3LZhQIKvW8a+Wmu+GlQQMmVsuF
3fzlYhWtPZ5Iupz/xUEEPfzzANjzh3JFCJFi8Hkdx8OWRmDt9nsEK8id2skZ96O/86cg3Yw5Kcq1
fbrGOrPGFwluvCD7iT5nSNubV6WiEM7cXDolp6o5OIxe0JLXiLnhZLlq66fDFfZvlUR9J/GHJykU
vzrNbBjkThOBzz+zmgQ2Z/gdxrmpuiRFY8sToK5t2lAMCmrh7V139fl2nw7WfGMPsNGd5teFOEIi
ko3p6C0aLqYmFUKBkLgqaOAOAxNCtHBcMFLbIiGBEFZLiRrRn9UOEzAIztLnNnVdudfgeDLtl+VR
ufEOoGCbTYqPcn6RGa3wOULrdpZHjKAibp0OKFTdGWjI5Kh5rp9RAQ/jRmBcfMR/7U88BVJ3TMbt
PCtg37LxkodAosBSoBNflt5Jtz0kMd/+Npy7XR4ngzvf8U/yQBxxDApl6H+CFiuX5q/zXMgClNg7
hXKEd82eixNW3dzrdI2g/IDSrTNHq11cAMHBTURYsXw1yy8Kp5OsyuqVMuEyXIPir22YYs1KOCQd
BmlTzXCp9OriOEcU7N8pjAnEcsyv+iJAg81tqNiy1Li6FdqzY+0/iqMAfN0TcirAOYJOSD6LOR+0
fJ2cTq+tbX7tHKx7FqBQ0FE/N/5ISHre08XbQsb6+vqYgTBdquYKLSf0J5xZ5Ickg7vd1g8YHGVs
w6FG/8Ddsw/dW1S16twrGLuU676zi3UtmWS1CpqScjJOQmneKRm/9sdgccRGEBC99Q6N8QHClQnh
M0XbayeDABfQnGQRVytiFEh2/gQ8k+PmsjKdU5T+Y5df4ifjVUHmTdAxATX6N/YI7o4Cujcx5izC
kUG6hGynyGvczNVwJ0akW1mJf4GIuGSVuxwtCC+E5vHWUcHpoJ8NVELjZgP2xJEG7OVuSwHqXl+d
bg+sMqYS1ts+S2WpUxRMVBYb0Yq82r1/aOrsp65VFr7tk3vT7+Mab6hiMHRnao+j2qnm8H3mWL7X
Dw/gX5gub5dTThzzdNfyxIFN+LUKVc3WWsrzNxPSZt3GAvxAq0iDhn1dDfulwb8DG/K0nZDn+4V5
OnrEAWS6d+1pvSgw8Xb3mPF5rsHqU0Qn0eu+WtQ2O1BGfgrQm6CjvyfT0t+778faYFySmL0+3Euc
pX5Z3zl5NcwhT6H3wHx36z9J/T1NGOGtHJO/g0q65mTFuCI49+996KngDDIb3q2izf3zsTIxKeJX
rAmIc1LqzI+UPFhbozINiJ0g/1fK5s7dGOlvcKpmnpO1rsYlM8T0pnkiszy2L3sATYHMzhwN9F2F
wmcVaMiiAE272eUq3Y30Jb9okxeMC1wzRN++4pcdiY5op86ah2cw0KBN9CBAG25ZcN3XY2IhgSi1
/amoJaSZEGepzT0Cn3VJnK/xI1iXZfQJ3APigqRws8sDRZAqDpXKsTXkL8vuXObqd/X0bo1l4sVV
kk6HMBvqL5YxjF2Ydsfmg+Qlzj7rWb76bPjyHJFjZ21VM1sPo4vjPsCxLFjWc45U/E/cF+A11XEu
sR3/x3NZ6UcFQJ1+HUQc729Y3leYHR1PSoPngd0qO4fl3Yp51PLu2geXjmLCX27qod/jpX6evGrO
D96TEqwyztWFKQrbPuQ8xzM+49M7tf9dAHCdZaVbG4Np3VUfSu5q0nmVC4kGDlfBmiA2pltSv3JV
qvvId5LHo9muh70lIhOKePPiSYkxLiToY5R1pohBgOMnr6711ZTf55CtmSkdzEtq/TvV+qES9OyV
gwkh7cg8UuPBJHBAUobS6H7+QQBGWe0+xsQ8qfp0Bs7Pee9Tifqr/G/qgBCpafxZ7pJ7GOSDEl4L
8xFduPDFrw0GALnkYB1115/Fg5bxD1DZfIYz/OgncPfwBCJMOIr0lXz94TeMTGEgQUJu3BKVCdFV
UjCRKyfBgUdlTcwu6s/6kE8a9ZTOyny5P6drhN/5n6LA+61stZEAlgNNZzZIW1KL6dXFGsXrlkxx
WE+4xz8t2LDpwRDz+Aq2Ie6KCGBuoDp00yB72RXz8BmYgi+ftckfikeqwjoqNWBuW9CUPA81ANkN
BXdQhjWdTxGx8Nz7bUvDnaNPnCXjNPgEADeGPMurQg+hcoVBz3kSddJJMpJZcbQs1Hcjl1mm0CO2
N0/vpK87vLRUCj+N/iWkmDmJsYvxFwsuE8i0+DxBftya81vjBPiygDnmcKdQQnTLaGckxTc+3sgS
VhqLmbeJPI0HiCTpfUX5NPlovJM70j6fEr2R6bCPOJ/MuE7Z9b7e8lF/6g0kAjKHGYlrtxfcOmWi
2si6mBsYn7kgNLXWEwLIQTAIKjrKPI/Kq/l0Oqh1dwaqZrhYInxzUO1iipxPPw9AEiU3IWkjH+Fo
31KhbqcP6F552p1G1d2Seu5TqxnH/cE0627b9diNvKwuLbmqoP9G5ZYoa3zuaUibD26cX9vXECKo
D2kRAYt/vKKTgpphWgMgCc5j9nd9lOnXYgUmL5mkwuxE1zTurf0BFErB4qp3gmDo/kZW6vD71Anx
gPlJE4f8Ds3vWUnUzEBsWDRNcsHCdFPrStAlVjKbQBT7dGPqZkOndzMMvyu8cZ/6TRC51uNSYugF
LpwzmarLwc6zxWbLPKuZPCwtoOqr2LAWt12n6Nt21Iledtw1xcg4hZB8Vme/xaI9xDVJrgDicKZI
f6nkL3QU6gtoPNth941E1D7nBXMZqDCcPZePFLbzzjeF8+b7prJQ8gNu6tire0FKb6na+ufotssE
iulr8tgIL5huX6sJEGF3T9GUaOMFpcX4Tl4nF9jpzsgXsTvZCdjDo5t4e/U4wyV6qbNCSPr0UAvZ
z3bRCco6I0IgZ6p2YYfmRSxyg5eXt802HXK+TqsAPKckclQmcCJXWCjnE6qmXsYEtlxgSqeXZMOJ
MG5rAjviUhCB7oZIUuNlFZE9cQv1mwrj1I4oa3YI3IRpOLmZ0kBDQroLiTtotFwmX3Ps9ctdbW7a
YZIhKoB0gK8XbGat8MQZPGnAh/N44BM0gGLo5y3M/T5nUT/uphGm14HuIG5OVJvQ+tdjgStpR+Jn
KzTG9tJgW5dFuuP3JBZ3knQWP5IoyAoCSf65S/VZZPGUT7rbRKUWiFoD2cJyyYasR0sbfSzJ9RpS
5w+DHWftqvzx/1h92uLu9h79ZmxWakaYza5hkG2TkYKC/F48f3bpGWIJRtn5ABliRQswX8tN02gO
ZcXBecP5AI+NhgrTAgBJPTRLgwSt9SocIOncVe9R8+Sm1gu397B1kpnremG1gucfvqXtZyOVhsGV
XS7M0MTpMhvl+tRMaWVGcM9TCt24jOqVQSNh1NUrV/oxovThpha0p73X6xeTghxVbmmkqDxgO85p
+Zx8L4tJ52yl3CB50PbuhRHpTTzktpshvds4giBLhu7a4OstZELDuV96Zw6PAt7wTMccp9Mq/z9W
+CqII9Vc5DgpPrkQr1dZYDIESAWq/sB3bwDjoRsnCzuLzn0fGSbN5T+K4SIlue5rFkW1r5MUK1cA
qIK9SPOkZuHVvRKyDnaaaSLtxX5lhAe7PopvFET1uYisyxKJ1sBo12Qc7y6iZRU7CnfYdkZysDpY
ZU0H7n27Npu4lVXHte42q2gqYEWjq1uw5VCIFAVsSk73wHmRVLTeuR+TUDzpFZVeQ8wa0bC6MG1w
CZADxUc+9LoJZoAivDscxcr7xFMEWIwMZX9ovRbSORa9tiTy4/ghYYD8b5QwRV+xy08ltwHA5AI0
ijA8c0LBlCvGEKpvFlQ53AxRotLDGhlZp67LkPxgjLVRxGZzFuXcnBSIfe6MY/MtoRtJEVq2u6ls
7K0v9+OZCpFlMPPYVf8pOJFokMDFR7rISbgQILFx93vaavLuKp1nQcXKgNz/Z+/DzC4qOUQ6zpAW
p+uoKkwPqr2+O3f1dh4eRwNWCiGAipx9Spq1u/uCRbuOZTSUq+IFsUu3NfAd521bF9uDyItJkSu8
GsWSRJvsrxogYS9XkmhaSB1P5Zbqbs+mAjkRqCfFEqNQK5ehkvh1TZ3yCAifm8i559b2s8MmWHia
GkCD4HNYG1EBjQlQClmUO9uLXCBJCH2xH17VAuVg0GULO1Ly5sRNEk+ymh+Gz9cffCLRz95tuZYj
AY02LoR1V8q92JFcwqxwGk2L2bc9FOLW8bbRDkddiIhSmB6SzSSg8xiD8fHZcn6wwVSMhTuHE/cE
bUlRrxu09cjYSh289XN01lDST3J+fY6umJvXEysWvnCopb88W7YT/5PhPvNlE6SIe5kFcx5CHap/
Vw1tTNcUdXYOMWm2ZI4gn7TIhB7Uxj9TSx8VzS25IwbAtJaZR8Wg6YcOn8ZR+dQGX27zmY3DwAUB
8cVyTF11RHFlo1ItHA/46ndXMGbeL8UQeTevRTbkM1FPC4pOptwu1aq+JyxQeEhjkOa3oInttp60
WTLnLCo57IsnpyVEFgZ9mgCo7Aci9TVc+FG3zrdQFkeVxXEGXsTVRnuc75LeJhDFxgVQYJIMzqIP
HygovO7dNbYPNRIeyy4/uQnaLGytgCHMlaQpW2eWN1ZUL8cYbfXd2BBsCIH1yAnvN8Yuydz9RBuI
u4/NYD0ScUqFZJLgEO9HQjVZ6XumJ5h9raHSdZM6PZ6p0WmHSF71z6hHXonZdxsmPiTOq5EshXn0
GgwYpsYKWxc/WnOo+JSM8AdSIGnzw7XNtnLltKPU3BZBBBP5IHT3JLq/0XK9zxwUv00ivAbZZZWd
BtoZKfI8340lOeCYCkWatkWDB5nEtWMvwb1AzqgvwUjPxP27DNQs3cjjC2Nk4KLwuiIDqeCkB3tE
OwXbHZdMJ72phZ9ws4e43bfaWcwgdxrrg0Ypmf3HWIFDKZ7tr7fpCR99wK3CK2HG8c5q4c/7JM1V
Sc0Cz6aqPO4+BbARNYPyhQHKuDWLX2hFiiT3X6dC8lZDIIuwaEgSYb8gvu9m+cVqkwR/Yh5k1XYo
ilNrrrd794K6cc4Q7ZxDqYddFuA5juhsxFeGehtjFLtzgXx8lVRnWkU8ExFGIvUH9scr5hZyES7s
r+Ca52rMInHSRBd0WjvdNX3uIuamJA4uIuPsMnKnpcmlazuLaLrHqtj8wmUWdwV3A10nF2ibRIC5
LxXbvjQqI8OXHLRnHzELxWN8NY8H0zPnq/iR6YDqkTvYTK/VmvdCVT0l6ip+UunPqmlpE78Azojy
04OvRiR4pbfdNE7piDYkO+aLyp7v0+I7SGqOA1LTM1ihDGlCNVkE4tn7qlyh9SBa3ua1bTtEsB6g
P510FzcTqU5tuXvuCXblr5hCSyWzqiUL7FOmKLdNQPQqXZxVjPS5LGreMVmlaYikgmKGJ8fAFB2j
rm2YlYSgjunIA+WIrqlkzZCaEjypa0G1otXcxHFMfOt/0h/tvJl3vj86VWIdVvG+iw779aKj5G+2
ljbBTIZy4CvCxZ2owY6fHdfZGT1Ow3gLF+JC8TGAXwvZScSCBAMwH1t7vFTvyVddgswCr5OBGNNj
SARVkQm3eM6zmcVojst+ptyMdPEi3N/eDs8uD7Cj586uU4xuDaUo240dxML3kpo8aXGQVhLi19Zu
h1+w78KDwYEAigXsZX9LS5ir583HFUDnxfu6Tq+r/UxRQWJcrAVwZHs9AThtRTek8XX08mDygWYw
m9FAk4i/zHRpCrSsJLbGlgvP4ogOIzIj+D7crkbOQIO0bu8LLPXCmtB7NzIv9Hd+YjQjoxKaA5h7
y5NaipaNNkNi61CL4qtWJBKKGnqM47vV6rUmgSvJ+JhzBZ3ZCRfnQZ6GXkyTOzQUSM2TYqOdtGhq
EhxZwuCzsFjECyhcw4kgn43P4njmMMjBOrSiFlvyjzkXgWpAmi9tFMXRUQjssA5+zy8F16ObEwST
OlcxYeKS4IEis673g1gz5RQ/DjentGqnDa/ngNcsUa7gDMIR2baoHY87/RUhpuhFISJsomStWdN+
VZe2RLQDMa8xTA3pV+EXSkpsqu2ZSZjFsBXjpucMWE3+QQ3au7xifLNM1g3Mq11GNznV/L92RRxp
iw2jjVipy1ZHOEWHsJP94QCvhESlI92KkCkfLn6abAtAqjAnFBdyDWdFNuz+5tvQA5ju1BsFNoDV
hM0MRiT1ZhzFMrf+GIEZwzYBc98D4dTPceSPChH2uys/Gr30HDKH+F2OLs3sxCqdU0CSJExarsFi
7FHUOzpG+lGZqCzyXuwvVxroRkDNOY1Zha/9K/oD6HZlOHfdxtmOIfQurG+HRA8lJwaDi2gwCK2o
B67Konh4t1acRuxpwvEOpJVpt3slaJ/5YULpf7+N1T/pAzAJTQt+qK7CTc22HreMyjd5QsBjqhyo
4W19TqDodeWpMI1/T10PvcMCUSRhdVmCmeDwAeKaGmJkQ4AbbSlWnHhtbUhSLJaabHUIWIeCrt/C
GEGeXZalbYwVDJnf8em9/f6mDZAmEkZKBGhMgGWYS521dFgB5SvvpbQXi1Hh4k2fUGvpaYjPJRZ2
95aPTHSWq70th7gyYjb1d2tI46fTSZsfR729mjBS9F0Q44Trtxu6gN2C3JQhpszKxOvrXksyqCa4
fKvegvxyle/ltn/pqKBDqVEls+ERAyHrP0C2RmbFMlNyABloj5/SOnv39BCsWxSUkeoZW2UXGvK0
eZM1wNFRFo15N+uK0rpkkWZBMx8pzwDD0trEhEX9+4hqeRTodR/CPuxZWcc9gweNoqXSJM7nR4dB
kZPT31kUQQXn8Mrm3XjWZy0VRDyZsQaAu8oizXiF7rG3VgqprQT/YQV/HVEnx6tUlrUsBhHilaIk
iAI2YhnC+p65iDO+aTCZC03l9gmsvr4sL68z0G9GBW7kvt0SLCqQImvwrj/U4dVpdeoMmcwv6IRE
d0mtASAWxxJNkKCmZfS3uwKO+44/akd9fTZ8kLn9rctZXeNcu8PYTQiedmKBg8Tbow4SM0rqJYzy
sB/lOMoDNOwFCCn4tMB7dmB3ELWKe1Iw5BHh2PKvKH84iFo+80ReFlRg6sAHhPxAKnp/JIQ+m9+F
OFUYYcIe4G11n9O8DgdzWRcLWh8Ww2f/pjqhdn7+nETAOqk2d9Xqxo1lKt8xHQVuPMD9Ik0lIa52
tw9SbXf2RCLTwmYTHM8GwRYqseX5GFD+iwXEqHIVWby8zo8i+avcnI0wqEBuxCO5gUglWrhLmwSy
SS/xvmzGDmpOkS6k/ktSqXp0EmyqDEB78PLi7tPDGBhs3eF/Ks+7/Wt7zM7i8qlHPZGqdthC+DXC
648Uqn8QcJjsJ1jw1vH/tj0UWdhsPGnxsWH3D9RXPk86l+Q2RTVBnFqVVtxVw8W4cZuXTXUOBY0v
pOWlfEoWnrZgS3QyV9S+EeBkVQ4yiPvsIlTqohRGgV5HR+mU+kj1AwW5Y7Qjphp0HxccapaRV3FP
C7zgH69A/qxMFUZV2hAi36x+R9jiP4D02mGj3RD38pg9wuFGZBagMuPrKsGnvn22+dT8dB1VPSIA
hzCE3otBwLWRTCiXQ4PJ1Ky4yrcVFq4bw+XiSj6rTs9MGtsu4xJHlUPWZ0f1JVV/a0ZZcWCHQYsL
PZiEprogqTL2WXb9k4eL110U5I+MymDneqpU5hb22eJkVOk5lqU2N7JssFHoQoBhEn1VbZSX5B66
TUquzKqHXvdup9nr1k5ilF8dqmeI+66zgOZGBlL1UpvV1h47DTTp32qKuWy1VoGPs2f1dJ1vyhZW
5ACmxlvmV5usLZH9uDjaR0hbNZkGmfHPOpdlGoo+MrSOjuMPOoBTiNqz+0YQtKYJ2JpVjGc+Y1x9
yrdMuSxXIDPqSV4yS0Ma2VOzm7spe5VVYsutDHMpc/suRLcerNMC8Gp3956Pih1Fi5e9kZJjAciI
l58JnY2yOCO7a6WJzrUTg7gHpRwTCv89PSJxUq/xqPMh1eFEV3aHUa/8dB2uiy5frgZwdBKmaWSQ
1m7Bj3W9M3YVwVYs4t3xyxX39B0plU+snFF71RdQ+mFLGnmlv/bpt7Vsq98Z9Y4AeC2HUtQeBZR4
w+x2FWcq2q7h2083AMZ8nair6tEUtfmj/yPH1hM+vCSLx+lnOkhCx8hocc3Xkb4GyT+7UpY9foRB
XBxO518iNjta3IN2lTx7xIvogVXUvdV+4LOG7f+U6WHAJ6PZz32y4JIxm9tdXVfEmNyboJLPM/o9
7MW0WkbME+F5T1aXnqInEZ/ki0K3Jd4vVEXqW/HQAj4xnQZCN5D4Spj0CHXSPQMQNtPT4zwWUqFL
0l+eKvGN1uaELkpo2uibSpZ6/EvIk+7FdngNHqHpRCU48CDSG82jxsHJCcyA8pyNomNycSR2fXsY
kMOg7p4+1N5fJW+JAdbEbFzk/3uxCco/AtJn6QMjYnEgNxzQfVvotWZ5I2VXr3cfanTcg56/lQsW
7qZlnFnKezqr6m0U0oNVk8VeLaWI/2sxHttq5dka3ruGByGbgr9lMJIGww3nVaLIK262PLbNildi
IB5X9ISdkCbKIvrAEElQ9Mm2SWF4uAX3pD1c1Y43H9CN0VAXoIYvYAhtb0ucFQueRwwqC23uNzqx
5g5KxOlRfNrT1RyBuOlLW1PYHzoYMrXCSwj0pQTE7yCzaPllNsR82TI7laaZBDMJRajmddZXvL3e
SdYXkzgI9x4ubR6CKo5Oi+O9oFBqBkVsvYv9RJbxw1WK+He7X6JgU4wLsIM1OrO0p+istyoKwOyc
GKEBzTcjiGP9nC4rQV9k8NgABjjsTOrRNNqinBzCFItqMCOJUWAmSeMSl+QKRJ/gOWLAdPkuJrSa
dTuLLSfwiL4SRbUEH8ex85fNPn0oQ8U6P2TK/uCq193KDs8WlmKuH+15jAgmvH+sfm2PV8IMzkh7
nvz70s3/06IxsApskNIy0IwgnbqIoM4k22PLQ/n7cf5Pc0tKSexWStLhclxHeVNNJMZ95xV19cBO
XCLY26H29ZTVJEsWC0tS1n0J2cDww9TlV8SinmuNWWveL3u/7DZJiKt+x5OhoXLaJSo0RluUIqrF
0quUbamwTxRd7zVfBkWnqwjHF94w9qxZNUMWooisMEHb1QHKaavjKuP2IEu69QX419N9vyIwU0EP
3mvYQiIGHXpTBiHK8Wxuvh4kuUt+LJjxaRX76cK3tl51kxVh4J42lPePWNosoVslKosVw9Gks2Rw
kjokQ27gwxLXEGhf6Clq6niQWGObAqJ/wkmHQS/BEaAX8GtpPfYA2ksLuBkl3cKcLztiwilMWTfQ
LIF64msE6ESj+ZBjBQU4jo9mRxQMsqMrbbmVCrRr8BkhHHVh7SniXS5vcmPPk2g+0kWMd1D4mdj0
yQkaZDiU/m4gmuR1m6Q5IceCMQgQ6ib83c1LsTQn+PDCRNDDl8mJp+MCcGNPB4IqsrGLcFRQYWQ+
aCyfCCS10q23F8gBwCfEPqQ5VPCy1bwk6aSBgD16mi8iDmDhHACWg5S/DFJ3ZXY+Gw1frZ+QV4bW
JCIrJl0sUQF8XQrXITMtPRio7yKMETLdfsiTUqoVqa0D4lmkLJoHZ9LP4y01fIdERcNylRr1snXI
vTac7pkxMpyFnkjfV4zc+wGE240ug4vk6zZSUSMFDEOGzbqi8q1J8+d33A0o5HrTMxU3JCNPAVI7
k69uRaW4vqVa1s3XYElPNCrWsdisqUIQZPIg2ttW4E8KXBP/UqgFVlAZQ3afHZE9m350EHbSFAUG
cdtQklLva+BYbNem12b5yi/kRTUhGwTIeibDAv+ycdazk35llXcXIbab8wcWh+6GWH5DQdRVhOYX
ueKFihy8V+TP0t773qnth2xesh8j4/94+TTNFQ4vZ0UVunpWo7ZXwsrhJxkSjfdQVzAcEZ+3vEus
oCUUmpKwnGQMd250XSFr6hNlzlSYuyBXGEK73wnipH5Wy1e980v2lBZGNPmAQsQEd6je2o0Wijr6
YOhSELPl+Ax4PZ2HkReXoUQ3a+S9D5QLorVRgrfP+uK+QwHuUeLKpPv4g+WsEYY0llm5nSkRnZbV
6ete6Qalphsy8RSwJcV4iX+5b0YenMHTDdfKTYIUvfjavweXAj1rnD/zNPCUHontQ4lxvHuduPD1
xmqBfKN9iKyuUhKegfIp1Pc3jbY1Nkl/OtnFpEoVynLa9qo457rIZJN/JJpHLY2Nq0lYIX9bBfrK
gfWGlNJlQX4TuCy1ZcAsjA0rXecCOU2B7teQSXzNKr7T7vUVi71N1jDUokqOQ3MeUPOBZZIzFEk7
6rHWdNwqz1LqygJPdyLwcNA2qxxApoJe/Bmq/8uU76UbHs1tpUhaQ98g5MQiX0H11nmEMLtKwU/U
NbylxJvZurrL9buz59vcFq61CYyMYhaW5UKyCnr39iwrJmr5i6k0P/cf5p4n3zAYfpXmOhE7/1Nn
u3LTtZ8u1icL90fZLmldNE0Tqj796hnQ7TPU2TtCK/LUT+u/Y7tI62EvEM2R3ju5KbjNrbM/Bn85
mHZ8N/ZXVbEnj4/jKmu9WcntzJa37iYE/91URwqO1PNSfDKRJa/tLwDFgJmSrYWo2T+XC727veqO
4AfgV2I1VHAWPTbnYnLxzyQRoeR7AjRTTHY2w68RB8uo6CXvzFF9Q9avTdR2HriYY7xUI2hIYFrp
oH727pTG4eNOb+lnnzyDaRLQg0F1IBCPVv4iw0ZvnU091sAz1TG/h1oQvm7W1KLC9wdOZCIJ4vjj
C/9s9JZC/hCqYS4f712c5miUi4P2nyK/BPAfyrKFNIVhgiQz7h6LnutydLXDGBRtd6HzaPEPwS5x
UVZxeORMVjRa7tI03Q/jKJnD03bvCy5f87ROjsiT
`protect end_protected
