--  Module : ldpc_encoder_pkg.vhd
--
--  Description :
--    This package defines constants and types used by the low-density parity
--  check (LDPC) encoder.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ldpc_encoder_pkg_1k_45 is

  -- constants
  constant C_ASM_LENGTH : natural := 64;     -- attached sync marker length
  constant C_LC_k       : natural := 1024;    -- k = information block size
  constant C_UC_K       : natural := 8;       -- rate = K/(K+2)

                                              -- n = code block size
  constant C_LC_n       : natural := (C_LC_k * (C_UC_K + 2)) / C_UC_K;
                                              -- M = submatrix size
  constant C_UC_M       : natural := C_LC_k / C_UC_K;
                                              -- m = circulant size
  constant C_LC_m       : natural := C_UC_M / 4;

  constant C_SHIFT_REGS : natural := 2 * C_UC_M / C_LC_m;
  constant C_CIRC_ROWS  : natural := C_LC_k / C_LC_m;

  --subtype asm_t is std_logic_vector(0 to C_ASM_LENGTH - 1);

  -- hard-coded attached sync marker for length = 256
  --constant C_ASM : asm_t :=
  --(
  --  x"FCB88938D8D76A4F_FCB88938D8D76A4F_034776C7272895B0_FCB88938D8D76A4F"
  --);

  subtype circulant_row_t is std_logic_vector(0 to C_SHIFT_REGS * C_LC_m - 1);
  type circulant_matrix_t is array (0 to C_CIRC_ROWS - 1) of circulant_row_t;

  -- hard-coded generator matrix for (n, k) = (1280, 1024) code
  constant C_G : circulant_matrix_t :=
  (
  "0110011110001110110010110101000111111110100000100001110101011100111110100101111101000010010010111111010101011001001001111010101000111110100000100110100100010011001100101110000001001011000011000100111110001000100001100010101110000000001101000011001011101111",
  "0100001010110010011101100010010110011111100011011010000111100001111110000100011100101101000110111101100101000011110100111001010000101001001001100001010101110101101110100100001101001100011010000001100011101111001101001001101000100111110010100001110011000100",
  "1110110010010000000000111001011101100100101001001010000001100011100110111100111011000100101001101101000001011011101001110000111111100111000101010101101111100001011111111111000010011100110000010110111000101110001000000101100101111111000101010110011111100101",
  "0101011000010110000100000001110011101010000001100000111000101011101101100111001100000110100010111001001000111011110111111000101110111001101110010011010000111101000001001001110001100011101010000011001100111110100111001111111010000000100110110011011000101101",
  "1001110101000001011000110100110001000000010011100001011111011010001110110100000101100001111100100101001000110101100110010010111011101010010010110100101110001011010001101001000010111100111000011111100111011010001101101010000100010110010000111001101110110001",
  "0101110101110010010101001011010100010101101101001001011110001011000000001101000001010010001001000001000001111011110110010000010011001000010111010111111001011000000001000101000111110001101001011110111010011101000110001001011110010001001111011010011011111001",
  "0100001010000001100111110110000100110100001101110111001111001010000100011010011001001001001010100100100000110010111101000011111110000100100111000001000111101101111100001111111010000110010011111100110000100111000001000000000010010111001001101101011001101110",
  "1000100111101110001010100100010001101000010111000001111101100111000111011111011011100100000101100101000001111011111100101110111110000111010110011100001011111011010100100001011000101010101111110010101101100001110100111111101110011000100001110000100011000100",
  "0100101010001111111010100000100101010011010001010010001101010100101000110011111000101110011100110010011100011110100000100001000100010110110111110110001011100101000000111101111110000001111101001000100001001000101111010000111111111001010111011111001101010111",
  "1001101111100000101001111011001101100001011100100101011011101011100110100100110100001011101101001111111000111010001110100001100111111010101001100011110110011110011001010011001010001001000110001101011010011001101110100011010101001100110111100110111111100000",
  "1000010010001011000111111110010100001010101101011000101001101111001101000001011100000111111100011110111100110110010001110100101111110110001000111010011110100101101000110101111011001001101110100010010010010000100110110110111001100100101001111010100010011000",
  "1011110111011111001110111010111001110010000000101111101000100110100001101111100100001100010101111010000000111001100111110010000010010111001010111001101000110001100001111011001001000101101011101110000011000101101000110011100001001001010110011010101011011001",
  "1100111101110010011011000010011101111011001110000100001010011010101110100011011111000010010001001110111001110111000101111101101111100100010111001001100111001010011111100011111000000001001110110111101110000000000011001010010001100101001001111111001011100111",
  "0111010111000110001101111000001000011100110001000000000100110111010100011110011010011111000101100100000101001011000101010101111111011111000110010110010011011110111100010011110001110001111101110110111010011110100000000100010001101100010111001110110010000110",
  "0110111100101010011011011111100010011111111100101011111110000010110100110110001001010011010101010010010001000110011010011000000111010101111100010100101011000001111000011100001001001010111010101010100010000101000011011000001101111010001111000101000100100000",
  "1011101010101011101011011100001100011110110011110000011001101101011101100101001110000011010010001111110001011101010011010101010001000011101011010100011011001111001100110100001000000001001011000110001111101011111000101101110011011000001100101110111110001110",
  "1110011011101100100000101111000101001010101011111110011110000010000101001101100010011110001110000010001111001000001101000000001010001011010010001101011010111111110010000010001110111000100110100110100010100011010101100010011011101000100111111110000100100001",
  "0100101110111010101000110011000100100000111011000001011011001001011010101101101010111110000001101101100000000011110110100110110111111100110010001001110101000001111001010111101100010000111010001100110000111111111100000001010001001101101101110100001000000110",
  "0101000000111111110101011000011001010010111101101000101110010001100101111101011010011101111100110001001010011100011101100100111010001011001000010100001111110111101000110110111011110011101110100111110000100111100010010110110001010110000011110110011110110101",
  "1101011100000011100100001110011010011000101100110011011111101010100010010101011010000011011000110010101000010110100000011101111101001011010011101001001010001100010000011110110000111101100111001101111111011001001011101011001010100101110101011100100001011100",
  "0010101001010000100010001011110101110110110010110110100000010000110010110110100100111101001000011100000011101001111011111101010111111001100100100101000001101110001010011001110011100000100000101001000000010001010101011010011000001011100100111010101000010110",
  "0001100011111110111111101100111010110000000001100011010100110110100101010100100001110000100010010100101110110011000110111011100101100110111100111111110110010111111000110010101101011000101000000010101000111001010000100111101001011100110110001101111010011111",
  "0001101010001111100001100001011011000101111101111101001010110010010110101101001010111100010011101011111100011110100001101101101110101100111101111011111111111010111100110101100010010101100101111010011101110111011001010100110000010010110111010001001101100100",
  "1111111111000000001110100101100111011100010001010000010100100111001100111011010011001000011100011011101010100010111010100011001110010011101001110101000110100110111110011101011100101110010011010110100110110101000011000111111111110111010000010101000111111001",
  "0111101111101000010100011001110110101111011011111111101011111010001001101000110110111010011100111010001101010110000100101000110000000100000110001011111000101100000110100100001101000110010110100110000011000110110111110110010100001110001001000011100010100000",
  "1110110000100101110111000000010101100110101011101110010010101000101001110010101000000011000010101011000100011111101101100001000011011101011101001101101011110111011000101111011011010101011001010101010101001110101011101011011100010101111101111010111001101100",
  "0101000101000111111110010000101011111111000011101110110000000001000100101010100110010110011011001000011100010111000001011011000111101001001101011111111100110000010001101110001100101001010101110101010001101101011010011111110010111000101000011011110100000110",
  "0110101010000000111010100110111101110001101000101001010100000110111011110111100010101010110011111000110101010010101101011110110110011111000010100100100101100110011000011011001110110110100011100100101100010111101011111001011001011011001010000010110000101110",
  "0111010101011000001000100111001000010110111001010100001010011001011111010000011100001011100111001010101100010011000000010101011101110110110001100001100111010010010101010000000011100010110101010001111110011000000001000101100101011101100111000111111110000011",
  "0110101000001101110110100001110111110110111010001011011000010000001001011101000011100000101000010010010000100111010010011110000011111110110110100100101000000110000001110010110101101001110101100000001111000111110110100111100101010001101010100011001101010101",
  "0110111010011111111011111111000000000111100101111100101111110001111010010011011011001000001001001100100111000001111010101111010111010100011000000111111001000110100010001110110101111011000011101001001011100001011000001010110101110011000100010100000010101101",
  "0011001011111110111111001010111101110000100001100011101101110101001110000100011011110001000100001100010011100010001111011111111101111001110100111111011101010011000001100100011001001000111110101000001100000100010100101111010110111001111011011000010001000101"
    );
  
  -- functions


end ldpc_encoder_pkg_1k_45;
