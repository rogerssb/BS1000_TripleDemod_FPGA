/*
    History
    12-??-19    Changed DECIMATION from 4 to 2 to allow 20Mb data rates
    12-18-19    Added reset signal to interpolators to avoid random resets putting system in unstable state.

       First pilot data pair in 50-50 mode is -0.373817, 0.128822, -0.361626, 0.0697403
    First trellis pairs in 50-50 mode are -0.360298, 0.167099   -0.361679, 0.102417
*/
`include "stcDefines.vh"
`timescale 1ns/100ps

module trellisProcess (
    input                   oldNew,
                            clk,
                            clkEnable,
                            reset,
                            frameStart,
                            inputValid,
                            TwoClksPerTrellis,
                            estimatesDone,
    input   signed  [17:0]  dinReal,
                            dinImag,
                            h0EstRealIn,
                            h0EstImagIn,
                            h1EstRealIn,
                            h1EstImagIn,
                            ch0MuIn,
                            ch1MuIn,
    input   signed  [3:0]   m_ndx0,
                            m_ndx1,
    input   signed  [5:0]   deltaTauEstIn,
    output  reg             outputEn,
    output  reg     [3:0]   outputBits
);


    //******************************* UUT *************************************

    //----------------------- Detection Filter --------------------------------
    wire            [47:0]  df_tdata;
    wire    signed  [17:0]  dfRealOutput = df_tdata[17+24:24],
                            dfImagOutput = df_tdata[17:0];
    DetectionFilter df (
        .aresetn(!reset),
        .aclk(clk),
        .aclken(clkEnable),
        .s_axis_data_tvalid(inputValid),                                        // input wire s_axis_data_tvalid
        .s_axis_data_tready(),                                                  // output wire s_axis_data_tready
        .s_axis_data_tdata({6'b0, dinReal, 6'b0, dinImag}),     // input wire [47 : 0] s_axis_data_tdata
        .m_axis_data_tvalid(dfValid),                                           // output wire m_axis_data_tvalid
        .m_axis_data_tdata(df_tdata)                                            // output wire [47 : 0] m_axis_data_tdata
    );

    //-------------------------- Estimators -----------------------------------

    reg     signed  [17:0]  h0EstReal,h0EstImag;
    reg     signed  [17:0]  h1EstReal,h1EstImag;
    reg     signed  [5:0]   deltaTauEst;
    reg             [17:0]  ch0Mu,ch1Mu;
    reg             [11:0]  sampleOut;

    //------------------------- Start Pulse Alignment -------------------------
    /*
    The start pulse coming from the pilot detector falls between 512 sample
    bursts. It indicates that the first sample of the next burst is a specific
    sample relative to the start of the pilot samples. The alignment module does three things:

    1) It creates an interpolate signal that is aligned with the first sample
        of the block of 4 samples that define a bit period. This signal is used
        by the interpolate blocks.
    2) It buffers the frame data while estimating and places idle time between the samples
        to keep from over-running the trellis detector. Note, estimating takes 5300 clocks
    3) It creates a valid signal timed to be true starting with the last bit of
        the pilot and staying true for the duration of the frame.

        Estimate time = 5300  clocks
        Incoming data = 13312 clocks
        Trellis time  = 800*4*4 = 12800 clocks

        Since the trellis plus estimating time is greater than 1 frame, the end of the
        trellis process may aoverlap the estimating time

        Time per frame at:
        10e6    332,736
        17e6
        19.7e6
    */
    wire    signed  [17:0]  faReal0,faImag0,faReal1,faImag1;
    wire    signed  [17:0]  faReal0New,faImag0New,faReal1New,faImag1New;
    wire    signed  [17:0]  faReal0Old,faImag0Old,faReal1Old,faImag1Old;
    reg                     estimatesDoneDly;

    always @(posedge clk) begin
        estimatesDoneDly <= estimatesDone;
        if (estimatesDoneDly) begin
            h0EstReal   <= h0EstRealIn;
            h0EstImag   <= h0EstImagIn;
            h1EstReal   <= h1EstRealIn;
            h1EstImag   <= h1EstImagIn;
            deltaTauEst <= deltaTauEstIn;
            ch0Mu       <= ch0MuIn;
            ch1Mu       <= ch1MuIn;
        end
    end

    integer SPARE_CODE_WORDS = 1; // first output is bogus
    assign  lastSampleReset = (sampleOut == `CODEWORDS_PER_FRAME + SPARE_CODE_WORDS);

    frameAlignment
    fa(
        .clk(clk),
        .clkEn(clkEnable),
        .reset(reset),
        .startOfFrame(frameStart),
        .estimatesDone(estimatesDoneDly),
        .valid(dfValid),
        .dinReal(dfRealOutput),
        .dinImag(dfImagOutput),
        .TwoClksPerTrellis(TwoClksPerTrellis),
        .m_ndx0(m_ndx0),
        .m_ndx1(m_ndx1),
        .clkEnOut(faClkEnOld),
        .myStartOfTrellis(myStartOfTrellisOld),
        .interpolate(interpolateOld),
        .doutReal0(faReal0Old),
        .doutImag0(faImag0Old),
        .doutReal1(faReal1Old),
        .doutImag1(faImag1Old)
    );

    frameAlignmentFifo
    faFifo(
        .clk(clk),
        .clkEn(clkEnable),
        .reset(reset),
        .startOfFrame(frameStart),
        .estimatesDone(estimatesDoneDly),
        .valid(dfValid),
        .dinReal(dfRealOutput),
        .dinImag(dfImagOutput),
        .TwoClksPerTrellis(TwoClksPerTrellis),
        .m_ndx0(m_ndx0),
        .m_ndx1(m_ndx1),
        .clkEnOut(faClkEnNew),
        .myStartOfTrellis(myStartOfTrellisNew),
        .interpolate(interpolateNew),
        .doutReal0(faReal0New),
        .doutImag0(faImag0New),
        .doutReal1(faReal1New),
        .doutImag1(faImag1New)
    );

    wire faClkEn            = (oldNew) ? faClkEnOld          : faClkEnNew;
    wire myStartOfTrellis   = (oldNew) ? myStartOfTrellisOld : myStartOfTrellisNew;
    wire interpolate        = (oldNew) ? interpolateOld      : interpolateNew;
    assign faReal0          = (oldNew) ? faReal0Old          : faReal0New;
    assign faImag0          = (oldNew) ? faImag0Old          : faImag0New;
    assign faReal1          = (oldNew) ? faReal1Old          : faReal1New;
    assign faImag1          = (oldNew) ? faImag1Old          : faImag1New;

//------------------------- Interpolators ---------------------------------

    wire    signed      [17:0]  sample0r, sample0i, sample1r, sample1i;
    interpolator ch0r(
        .clk(clk),
        .clkEn(1'b1),
        .reset(reset || myStartOfTrellis),
        .interpolate(faClkEn & interpolate),
        .mu(ch0Mu),
        .inputEn(faClkEn),
        .din(faReal0),
        .outputEn(interpOutEn),
        .dout(sample0r)
    );

    interpolator ch0i(
        .clk(clk),
        .clkEn(1'b1),
        .reset(reset || myStartOfTrellis),
        .interpolate(faClkEn & interpolate),
        .mu(ch0Mu),
        .inputEn(faClkEn),
        .din(faImag0),
        .outputEn(),
        .dout(sample0i)
    );

    interpolator ch1r(
        .clk(clk),
        .clkEn(1'b1),
        .reset(reset || myStartOfTrellis),
        .interpolate(faClkEn & interpolate),
        .mu(ch1Mu),
        .inputEn(faClkEn),
        .din(faReal1),
        .outputEn(),
        .dout(sample1r)
    );

    interpolator ch1i(
        .clk(clk),
        .clkEn(1'b1),
        .reset(reset || myStartOfTrellis),
        .interpolate(faClkEn & interpolate),
        .mu(ch1Mu),
        .inputEn(faClkEn),
        .din(faImag1),
        .outputEn(),
        .dout(sample1i)
    );

    //------------------------- Trellis Detector ------------------------------
    wire [3:0]   tdOutputBits;

    trellisDetector td(
        .clk(clk),
        .clkEn(1'b1),
        .reset(reset || lastSampleReset),
        .sampleEn(interpOutEn),
        .clksPerEq2(TwoClksPerTrellis),
        .startFrame(myStartOfTrellis),
        .in0Real(sample0r), .in0Imag(sample0i),
        .in1Real(sample1r), .in1Imag(sample1i),
        .deltaTauEst(deltaTauEst),
        .h0EstReal(h0EstReal), .h0EstImag(h0EstImag),
        .h1EstReal(h1EstReal), .h1EstImag(h1EstImag),
        .finalMetricOutputEn(),
        .finalMetric(),
        .outputEn(tdOutputEn),
        .outputBits(tdOutputBits)
    );

    always @(posedge clk) begin
        if (reset || myStartOfTrellis || lastSampleReset) begin
            sampleOut <= 0;
        end
        else if (tdOutputEn) begin
            sampleOut <= sampleOut+ 1;
        end

        if ((sampleOut >= SPARE_CODE_WORDS) && (sampleOut < `CODEWORDS_PER_FRAME + SPARE_CODE_WORDS)) begin        // skip first trellis output
            outputEn <= tdOutputEn;
        end
        else begin
            outputEn <= 0;
        end

        if (reset) begin
            outputBits <= 0;
        end
        else if (tdOutputEn) begin
            outputBits <= tdOutputBits;
        end
    end

    reg [17:0]  inCount, dfCount, faCount, tdCount, outCount, inLatch, dfLatch, faLatch, tdLatch, outLatch = 0;
    always @(posedge clk) begin
        if (frameStart) begin
            inCount     <= inputValid;
            dfCount     <= dfValid;
            faCount     <= faClkEn & interpolate;
            tdCount     <= interpOutEn;
            outCount    <= tdOutputEn;
            inLatch     <= inCount;
            dfLatch     <= dfCount;
            faLatch     <= faCount;
            tdLatch     <= tdCount;
            outLatch    <= outCount;
        end
        else begin
            if (inputValid) begin
                inCount <= inCount + 1;
            end
            if (dfValid) begin
                dfCount <= dfCount + 1;
            end
            if (faClkEn & interpolate) begin
                faCount <= faCount + 1;
            end
            if (interpOutEn) begin
                tdCount <= tdCount + 1;
        end
            if (tdOutputEn) begin
                outCount <= outCount + 1;
    end
        end
    end

Vio2x18 CountVios (
  .clk(clk),
  .probe_in0(inLatch),
  .probe_in1(dfLatch),
  .probe_in2(faLatch),
  .probe_in3(tdLatch),
  .probe_in4(outLatch),
  .probe_in5(18'b0),
  .probe_out0(),
  .probe_out1(),
  .probe_out2(),
  .probe_out3(),
  .probe_out4(),
  .probe_out5()
);

endmodule

