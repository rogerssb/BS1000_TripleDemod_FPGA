

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U71FUQf0qAsGxfI811Hw7L7fy3nJYTd83JjuLrHeStKqJTUSdPESLymcfn/cVpzfBW2bF3BmYXSP
e5wyjUbgzQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pWFieWO8oo9hfHkPbS1OEKBGvkAlQMLueuSIE7bWZbT6M/kqq/dye0/px/MdG8aHt5pikgi/t4lz
LuwJbIiNPyrhEa+tgcCOd+vb3cYReHlWv6qj2tNDsdeIKt71eaX1vjVYrragxGzIIBpV0lV9r6kP
KVvXjylDR6lRRoIz//M=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NL/pTlSg2Og5yC3YWVrNMxiSfHO/GibZQp2PQUi2R2a4HnjEylonymvH2vL9j8JouAuk0EFB8tc0
FPakv3CX4TojFCd8gaptzO4C8j2m1/36bqI9Uf+rv6QJs4sPJKomGGlgn1W0EQ98otaSuLPzoswO
7QVhIzc0r7KyYZieWEU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
iV99aGfQcwtekMk3L28+vYpw9Op8htG6fuBIg0zCTnTsG9RIAlgGEYAJA1TMbtP7znscQ9vJtEfT
T2W9slLueLoFJZrjCE/mxALz1CAlD25Ec+I45Zew3XrwE7ALGx0DdVLFvX6rrGYjjDSv4DlIm2VC
6VPRrT0nE7FzO45hOJpJqvRO6QHlNl9OA4qb1iEgAVoqUDz7Q3O1w5yurrFPSx5RObMnWO4Qir4o
LgFRirYZygtHGrCnsFsYiJLWkp+GPNATT9pDv2lpM9NKbSvhFFiGIbQHHydyE66fjDOgmN7gsXCA
UeWavj8i30EH4Fxe6GGfWT0D/Qx7pcscNmPo2Q==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GLCbDl+3CBTQ9mXi3N7iILMMdha19N1H4Xq77fJaHrjhhEYWFsrbEcAlCnAn2Kh520BkwISUGiHX
qhiC60l5dQBrHwPyukWPv6JPp600q2D4tTB4YMXGX59JzIzkFA/QrfOga9Qw0wCvItdYTofCqKo7
eKX3lnG98TeQJ8s8Na7clQL5NcFlbPxzsDOkoCF27W2dAEoIvbTv31NrWkRzh6kEnyUtVfJH1NWV
FG/ORKXULCX73nJx5iFYlTmU7C0VjbqKgPj1iuNvkn0R5JLIQMAtS6mdCRMQoKwPKsaF2wBBoBYk
2rIlVV4P3Xm15ZXC0wxW6lucSgd9Cn7JMSmKHA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wqk2o9IWswI8gqaghcvLi5Mb1OEEF1yuuxRzIAnMyN65arFFPQqZge265OnuRXAV+/iPV0UMsEv6
4dwyuTpRDf8wwbS873M0Q40Lco2/Dam5vuo5sBSb7YIBHHVlW8FOxDEzR9E70T4b82HLX09gCGbS
VHCF3MaIuKHgKOwPoM7xio+IRTmw/QcyxV+ZWxI4gbBzAdJw/7w30WQHXTjlOna/N9/0AC/gf+Ze
AGeCmAx2NVq7WHrX30TUb5uYeV0v1qhZcimC/tGQVg88BfXc/+4efXGKlwNimhMDrAakp9u1bwsa
V8i2/qUMV18HAwJfOTbqZhmb1ioPKYJivmvsDQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 103440)
`protect data_block
sUhxUjcPQ4hEyyDk6WJNmVur1tmjOXBLHHWAmvhRq6Lm8U8kWh6ym3dl8lP8aVWyDS1WFUe6kab+
C0+4a4p8xE0BYjgkpCNEoM4zxbJX8fYAjsq2z5zR1+hjOYQnvqO8dtHlAz3PYmP1s0lK98eK8inD
Uch7aLJ/5QxMccpO1mnswR0Ieppv1Fg6iWx5C2kN8a5Ho1onijYaOFnmvabJuIfuR6z5IMGVtLtP
Yjc233FBEwekSxBtLUZqrd63WpEjE8lAnWsSCk1D9/HVvhGNE5yKJB7cGJcjCc/0Bf/q44Oaxl3w
MY6eoMKm4ZhNk52Rvr2JcDKDjEH9TDWx5eUVuWOB3ndG7UJfmy+/mJoV6rYrdjFV0YU86C809Vmr
4+dgqIlaNXp+GAkUD+2Aq/DmGXVkBPNhabcCkqayJqFsLsZ1uldtCo5GOb3WynAzJSzUBWjUi+P2
TpTQarCNFoUPzfnk2i+oxpaKZOQdGTN0/z8sLvTendOORpYgBGXDOO+gYCmAeqMunuLf6zEFhPKv
ViY2lovZq+9A1SC/Br9AgQq3pFk08W4FNh55vIRI+FcoNJEuuSRM1E5HVmPNMb1Db746RDfAenV4
UewaXYdx7CdnonD8xDwkclIvyM4bk9y5EiCgj6UI1vNcCs+AomPfyQn4TjwSgc3QgnaGoKyRgG44
tHr5HTEeYEGdkBnJYITQxXhw5p6mPMYR+41Px2l0w8O8eR0KyDlf0Mb7DexdyDn8uVUwHOF4Moyl
nsqRXr3WbM/W/SPxCaMw29ceDM7ReDBigNgh/5LLL9L+p06+rCgI9Hs3rSKZohNQVD9g3iiS/GGm
FHgJkVqI9sk4Buvc+4/3pICq+ERVWHs49nfC4H7AWw/7zkrXiiJwMa4cij3LVT2ryotW6WgKjCVA
sODbv4rjVrDhEjpwNoPewHKqsscUeoXO4/wRFyacKWvII52qbeFpCNFtoCJFmSbXC5Hj/DtmX0IY
07fIttK4ujinO+zx7Rvu8JuAPQURoVDkEr3wDRHKngj8o67G4m3ExUjlXiAULzpLHwmyNIyRvx6E
26jG6HNzFljXqvu4+FtBhkU4p9qjknp6C11NzdMP4MWWXb+1slh3PjcnDXPdr9TrMaAAtAuwo6+f
h6joRmPvpS26uXSbnq5HpQJVMNNz1qpbC9CvfFLYor63wQ6wE0ewZSyVnkY637qrXuA3MCoCHDO6
8l0cW4BTp0B0XbmYFspPoRPl0WXu80aBSOHSWyrIcwRnQIZtgs+QKGRxjlWY41jAKX7md4hRELUJ
LWWoEsK0Ev2ms51mHDxs3o3Enz7U4S5inQtgp4hqxfAkDEF8ilC47jo3ePTraCSUiKEx1zoHuSaH
8GT3D6BymvnkeyyawNnEJj9WElVBZrszA6uidTGjOnAzcK+mjVi61iY5GCM7RVCtCpniikhe19iP
TVWYyZ3nj1hcDcH1R1Tyq7OcpYFGGRMuUbOzO9FKMxhz9TF1nvhh2WpeoIra+c3HGTHvbLYr2Bej
sIraYXOL/XPXbXKAMSDJczk79GVKctE17g7ojgpadbBMwyfHVfv4QFysXYWzWQPZ49uxzJnh6Vbt
53RX9s61qzt1PU6PjLwQttwOj9BZ/LBbWKiToJ43hrDlH3NGeD3FfHrQok08g8EPGEe36e+DLAdg
/kAB7vkhwD86iyt6aBVnGX2vwd+BzejnlTUnbUw/zTAieMIU72rQR2h3TWyZ3qKeQZ0ed5q+Kavl
u9/dUdSc1gQhXyENiS64t7fYxjQe5Fzm9UPBXbuiFlNq9zudzQMp0dSXnSpRbbP9AmobcR974anP
XV55ruAzCp7z99yIe4z5ZnAMhQRHgTSW10sRfmFeBeR/aVVZ3xTA0scZSO4d3knV5TfTBYtBOxcO
b7El7l9P/Umpz5f4qseYi1I26Q4Ug1rbDBKTySqeCdEPbHyxACo91jcJ/i3Vl0qSXb13gczW37Ql
4jE3TABhvE33q7Ik2ZM1C82mXP8q3aXFQ+F9weDG2euu5VbEl4ggtW/UWGEsd5aW9D64h38q+o2N
U/7zz/1/VTbfNjO4cAAE1Aa8KKZXGS7tHPGMWUzb7EKUNXulSeinCMvRtKDJ+HrlWNOrRwyMnjQf
8NmqSYRQK6xD18yvDPDbe1xPHwcnCCfbogD8aAUvThcI3LPJQrz67brZKcA7QOcPY7hfEGyS5dQL
yoCeHT3jaF+NK7zS8bSRBzZjb3Uz9UnNM82s+L/MV/x7X59JityB/gVKj+tpNjX8thqsOZgezaVE
L28JEdtq8cC6/g6ZtwQPpsuZDHH1cWbompA+7ILsUOf+8YEdKn0vtnMlM2ncMcnp+htmWrcggZHQ
3LGaxPSw678pOTBayjp8ZO3eahR25BvpZjmyEjGILk313eF3yH3RuOIGfMkSKf4KXpCCAyZaCYbM
r3cZGhXUxY0D0fAigza4r7K8JO2aoTHWdOfXRT8oGxZwFzIlw3q0pWjsz0yIaiS4U29AEJg40Uuu
SSm/TF5okSbs+v7RLrIfsxx3JRCKG79JxKVOXjGrTRf7pTlXW89Cnw285GOBMgS+KAKryygMHFpt
uOxOoDwlURwyvmBc1XUiJXt79wSRxD8w7whWplbiudNhLb3Pooidv0ZVLMAI21Q5ZeVoYJZOQ6Y+
ga5btNqOgIpkl/ZViS74P8m1iZ81hbViqBmoSdSh7by3rdBkh+LZiCsxw58BLsATtlvJxaGgFNSl
FkLP8HeGfHeCc4P8EHC7FqhQrTS8JfvRNkMrrF6tROaOrYk/C4Q31IEp219jvEkdrnHYbYv2Hy71
JtWyjXpgSdu8tzUJC5vMD61cEsLkv+VtK65iv2BMgcQGlSePZcULd5Svo3ciCMW3/qJeOOZmI1Zb
AuYNKGGCoz5D8AKlnIV/TRaBIVack7iiLWTVD5w2rikgm5MabfZQ0y0t/4aASedmPlXqlVZsre9E
+ojm2+3i9bJ6lzdRPTaSMQLIuzaVqaq8L9RZT37GlAfytsu8Y6qBaSKu4Fgo367iUrs9Th4USZul
StaRi6LUd98E+lg2TYjP8RmU9JFYY3sp8beY+rWjfS+cgGHtV/dxOVv4so4aVW2d+pgeGXvJR9ES
OD/eoKTlXKB8LbijWELw8CjooQ6Me2YCQTklch+8mOYGgsXtI0dIAH4tQ0cfki/kTBl1cCWkTObY
6CdiDENRCKDSKonqqxZAiiyCgMkCBvOReQLsAMgdZcALrbD+gPZo/gFauiLWa/Ut85YvgXVEq/R0
3rQ1QCHE5HUN2hykuNoZXyeOLKZ0OCgBD+JuYDow42PlF5n7TSII8vDr9TQOhqZfWNjgViARb+jo
Gyu+oB+Gq6LRJrWFChj7e8WQZzIljq0aZae+UjvIS1HXDAdeklrIAXQTVpMh/MBj3SsmpCz4mjGf
460k6vshFDxqQaZFv0bHOP3FfTrr5UDXk24qfE0xHv0KP80raEyp9RY8rXl9WDpfVunahfH3b7GF
5QCxjSxQ0UOCHkSQ2IC8xTQKCKU1hDZyAFy73CpveWAInB2CM86GF7KnRD7xGbCQNrEKA2xuP7ZN
72RARlD13Sh/8aRMN55oRt2DqYtnp4O0LJdmbgcrx8RS/coLeKKZLZD8FPRHDahGykemRcIkPiCa
GfmU3HrovO17mF+WrjuZXtmvkqsIW4Bu48JqOvaMqo/5L7BYAz8/phbnqlFUGBo7lIq2AmfmShXR
6tDCGxFNK8yxR1lUs0BqqaLrUE1HmxuUO4uMyRNEQSKFxmvEV/rwBdFmEG7Mdf2z2vTmUmwFZmIh
PHOIyIGV2Xh9iXaESEJNQ6isrph//dBLNep6agurYuX3LoO++FkpGXrcZYOMPq1Zain4t4CKigc/
iwRTWS/j1RUCL011BP1gi9KeTw6U8eOgz3lHcBgT8JU62WjnmSmOTWLduOfy16fRp1X/UvIjr521
0gTzaZj4HO2u0A3IsQ8LMdogt6qYbxoE5JEO36bsdV6O13w8quwHqrvr/lJyqezM/X6qM+h2kd1l
KAPyGfrW1clCyYUC7l7THEJqOrGIvqS3tuOp/jtf3o/niSlzy8nP9X0a55vCgJDpcF9Ww63Upqp+
hU3m2DEw6+I691kQ0TJek1QLQXwNdt99fXewt+nK7MTK9XcIbtby4yV3cd1I6Q3iAoUmMj/GgZv0
F3peNuamqNlSQO4QYQow4Tz+Q5g4Q1hCl21Rh2jdkhqNmL1LnOMaFlbUbYECRXgCbGSZFTRMAnk3
ZbVZcHxgScQf0e6f5ZeeToZfxkef1t0Pvzi3PipGKNYbbe/Zy/sEUvNFJfJiq28G1tzqxWuIyD2Z
P2RUEs4ckDVA/WhcXbb0/w6WC+MYlwC9t7vYMgzvu8KZLjwRVU+aHr5kmpWjJHgfC17z+MwXOJ9S
0EBz4lAl/2DO/ZHFIV65s52IUCgdqmfPoP5L//4fnhuhhVvgDOTo7OQDtUrFASBWgUQT47MQknU1
tbimOMvrdJ9/MSsGba+uDRvBEBmcL40MxFEU3BYIfCvAvfojoZvHSf1rXULMnpBmZex8j0GAwCK5
5d/JYMj6sMjH/zupVMCDRhj2nmy07D4oDySNnHD5K+4WDU6W0AqZzUNaf+OfctPUhUSYh7Pc+Rqi
Q5U7HMMuiiS1HPwwo8Au2He5d26HUFn+EvfODBmeJDPBo5KrFJ/v+hIGEgGDzdtYwBn8mpRhpo7d
rKxDZUtd83x+FE02OArePl8KaLTrt7LQeRLyj+LfqJTuL4sNl8fcXI7vJYAl3URq5KfJdXT7ZSVQ
ed59ye9W3nlJm9gW6SsXY3yer4AtH+VfRG2w8wETHKwx79Lu3C1SfRGCwdadwdSe6O+a+mS8kPuw
19fRD8cXLXKhjT3WsFQreT+N+fofAOK2Yg5e39BRCWWqmvbPe9V4tGQaBI1OWgNcWswqciHqFqQY
oDXBqKFWIaVZ9j/Y+nRwzySiiRXGckhwZqUQ1jhi8+kjJzw7+xUL6H7hY9el7sgkbdeKOutP7GBq
ZSYz/R79TZN3KhPt7GOvyXhMgLL6gzKJCsz0jBQQc+q51fo4CuYRZij7EgDersO2MHKujA8/vVmh
ELJVEW7pFH4Iut01KxHquw2uDW54JEQHz9jF93f8sIkyXLGkNEhXwHQmo26h76v1UUoaFZN1s0hm
izbBEj12ocx+4w7AaaDIIUA8Q4abWrI8ns+2cYm2Bh8f+PKJVFdQCsF3dl0oibbE8uYkK58B7ThS
cys9s0VyTN7qjL7FI3DUwYotyGEZ1V+ZzPbht8ACIv0ahipwFKwoi9NonNEfxiYcfRB3sf6zRSix
95UJSH6akBHTjj2LKO0R/oBsv9AcXqLXYTLpyoC5T5uWwfMqVKQ/twO5mUcnueqJZ9EJssfjiRrM
ejHIEsW+5Gc5M4B13FwPECv1Sjd4RIJxX0ww0sqnKTBVTtsQhhd0TqbM0/CSTzXJAxB0lKDhunGw
SWIiZHrs3vOnrh0vZNkXuUyVSnRCiFeaL7y3U7Q1PwkTgOzGp8P+0uBAMbkdh3z9p6OMWy6X5kIh
ibwNTuKBEXtaFZ9dyf2m9YL2Soo8hpIj6QwlZg9I6wZqDlRmE5rzfaAHfsxOi7fHVf7p7EZ17CHY
TDRHSe2gA78OOQ9Jax6t7t2/rpeA5tgvVLkya/kGDYb8vJQjKNSY5Y7GABmiUrgnkVKO1veqYbAR
VVzbxtrar2KUzEzNHK/3QKWO8LCLVS/GwzQZjuVVsdxijOE4vsk1zoS+D506mGNFAM16hkSk1E+8
0aMRCoTlSNcorl2f+edJ4+RmMcQt1LK812DMZE6yVfaORfhvNyXXsaV446KlLHDmVYJEBcNYwGhw
2ZoSSFf+ibrAFhgPCZbKGtuxpZJnksykS1Ht4MGsaqB41mAvLyIil6UQbv0LYAxO9cMF9TwM37mH
DPkDZPOXgKjaIAXLG6GsZ6cBxhlWTnc/iP57CYM6kKVPR/0udWMcrMx7dmvgtty5vIaNmR9A1XyA
pqpUm2DMXx7oO5utRDCfX9Sxd+jp3sMpS0zHPDM7+YWk70rSbgwxgHFV4i3braalis/hbF+xuLcS
9TOKmMppTvb81JM469fw/VLwTO/b5LnUyLd2tMtP7uv7yfakUbxgxQhZmUMjKAx4yq4ZpQQyrP1W
jum4RCSGEIsGpzwNqfugPehXFVye192XryE74dILkZQHvGSGmdiskAjDR+vX6/GKRkIXYmV416pK
sjdoGar4KwvOqlwDvjb2IkyqhqOpYHHcVl9ppPinXXuvlvPJesNqJ0PVthYx5IFDYdmlMJ+LW92/
y6lcWol1KO74UsBdFApO0y5op0XZMdSwcE9HKk1rg6sXPnOhK8DKEoMGqdujp+D0TfXm9CGClry6
oZK1r0YDcXmQlH1jg/L+mPKU/n7rTNoQtqKBhg+gm5KL706D8CeLOOVqr7/z3OpaCCHuONnw+sYU
k+VqQTSzQO1scBvIfk1YOiRTpm77PJQlxT3/frub6DfgsQQyIjhbNhQWMcbYhRMSdIIaTETHIq35
69DCjaKBcvMB4gqzGlK0SSegELybS+1D/EmFmfJXWb9tNwogYAXuhSfeUhRlLFMVTFpHE/RwNdA3
HPnTna2TBTmbxYkIOme25GglvGc/Sa1wh7Xr0gFU0oVUCX4NwiF4roevTdSH3TXx47SfhYkd4VOe
jgYbNKY1iV0kEx2f8G4ThqbGNV6Ysojn13TnoA8uEu2RVKuQ0xsqMgo645hPjr9XmAgahsevOwVq
aCuuP0OtZblcWi2oaF9m4CvkaHlv1PYTaPaI/J9yWJhr/90ztS6Ro4oZbI+oadOnv++zE3UpeJU6
jBkSK1u2G8riFQw3Vsex/7FPAth05/dGeSgk99J+mJaVeYVzOvTJcufCkyDxP5FMuA1tFMZSFy6F
vhsrV208WDrU8Rd3bmedWFv+MFiyUe/E/Z2ose35H0P1wW916mH3vzZmy6yyhZTUd7uXjSgn+LUf
Pmi9GM6dYfgAHL2vzc5nGE5ZrF9wKwpgfDiLokSFA9G6elOhOeBV81oVwBTAJ/eHhwOaYoTXCyhR
bBfzN28aQcse4xHH8DdGHEtFuMIdT6bP3dvdeegP4a8y+yDpq5hB1takHnKYSl1/iuFR2rKi9cZy
RUoB2Ga78PyUas4NS9XKCBZQY0nwx4dx1U56bLzpEKJV4M7Wh/EC9b4Jt8M49KlKDTOhCD7pEixM
U6PqcNwAOjIfUqQV06lQB/Qtws8OcFOJbRaYRqVER4wJUdZtvzs9/Z4ZJcnWK3Z900BsxGd6nnRv
biR7p+SAldzCvYK2E0Qkse3tidHU+Y1Dkn67W6R3WHVEt0L7nDE7TyB7g8GrPbFRmkgnQ0BwDYIW
SdKMQC9KWsJ9A+l8XXOxkueV7sgWtths31BKNNNgWrI6ARVku6enZRTEGWhAKMFOEbqomQ0jPOkd
ME0XI5hLeXpQ+hk4NcZmXeQuDwsgZ2S7WmxyA50zLNjGc5f+hOgUct6GaTZPH9NuI3mR0SSTdgDP
/swV0Ygr9JWRbqEQuhwxBVL3ndWuvPtBXJMGyBESyr1qRbo4jtIrM3icGct7KTgFr29n96yscC8F
aazIWUEyHncTTkgMyt9/kRbVw6xlv/JJRmIXmgl7iCpx20KxnMQEF+f8VlGN8vMsfrt98kbOfPqL
0CMd3kO29mjjDBBWBD2lPKfgD/pXFm4CV5DJ62uZPsxNMHJTeP1Y7o6Gsyuqq5pStLMBfWTOqKl9
TuImodKEO3PhUfqY8O6EU9QgxPGKs6AHt1EZuEp9VXjiD3zmlKgLMioSJEhRRE/whw85h82s7Z79
NyeJckuSduvU8T4UGVfGDZk3QKIHnwdPf8IJrfV8jIrR9IZTZOGYJr8ZFQ++vwqNP2/u6IsS9wLa
Ahbw2DEMN7b/KHBJX0DWV2xv7BQdcsPwLn8RMVRGDqiYGmswo6FhQq3UpCoZkQR2bmy8CzXqamna
91+ZA2V8k9E1OSK0GVOw/mEYqPNLA7n1ulB5fSbzlnAC0/vo+iGalhbtFUsBe/8NHQkMN7/eqHt0
IUhikzYTgvnXDqnaLCFGLYGBz3DeohjGoMUh5YkW5O2AwDbWyVuQkilU5ZbWz+FGqe6wlEk0EdTX
JIpi8fzfLBTpICH+QqCYNmk42uYbR8o+51K2ClWM962wKG5LzDUy0xTsbLjTa5QBZZvALi9uKfQ0
Sa+uDXmKvCvCpVB4FB/RsfFBZGdB7iY8GT53ciVpEZnA4F6yC0BceWm3IiWroPlbFtoyvxUb8ck0
qz6PCAuT2P6A8FT/DUqS+uaS+zo2Z2EdMgcsUsLHDltXuU7hVGEcJGf+joFvgR7a1Q//7tI4w6BZ
4kMXBqouNSKijQxPfp5KvDkzf2Nc68E6oQl1Iop1N2Drp/2j9m7a19hqVYjH9a6Po51v37wPyGFH
AYyWF/sDf1r9a3oiUXuz9lXHc3lnY5rAMdN8opPpLJJTfp2uP+dTsbbjuiF85exqeY1n70nLzNqc
Ks4GUKvYouc8od7JAX0fueeYbSjTpZgUZ7gwHuhu8XK00YCJC02wiAq0DwrnpQGp2SPD9Rx976jh
HewWG02SM+1Ck2s0td3XA/BtSUZbo7H/+nFOYEJ0kp5p6PVb5ZxeR67uj+fW0TDEV9oUSadKktT7
kWEmVSo2mdDYMlGRTGXdAPQEjwqSYKEAa3vgCdvZ8LSQGTCxp3B4mgUr7tlBVWHGwUaydgCT4/iV
AdtXHkTjqHZUGqwkfzJ1sgmKn8MKdE/vtzbNFSBuRmvwHHN9nbe5On7vibeG5TYZeayfihnfbZA4
m0QO4D15ZXvHZwD+/+fQNnVhVypJ1Zwq8JBs7rL3itDClf8O2+mnf+ubrYTievroBJlhL3T4vFQL
7e8dWtUlpoeoyiTw/JOUQENOtdmsZdu5Viwb7FndN03EdwXAVqdGHLIbrlmHHkRURXPUg/8jVi1z
h8ii4EDTThKjDuhsVPCGkunhnddTSOAGKcEibQpeqcOxjpFNj/he/QbnpSi0TiMjv+VjfEzfDd4K
E8sDrgpY1cbLBswyZrH/vdGay/d391N0rFh3IlUXaglX37yUkdhzo8DdAPpX/Mb5XBV6PwIiGAti
6/9jC9hEyJduwAMUtDGxyBzMTDY/1wxdSVu2Q7dvxrZyQy4JYE65SDxeAPA/UCgJepFrg/Zu7bq/
PXfRZOSNQVPq31R+X9JLetV1LA2d7JGm1RC25Z726v4mKuN8aGShCqGdeoSdWxEpp0vYZBEWiRwG
mstTY3/zAWOyfP11W+bQ7ooIxXbdJ1IGUvET8Ms9DXIuhXT0wZ0WaYCp8QvB6hd2VgSUlOB2euA4
ZJ0XiuJpnM1MatFKWtc8BHpktB/Q0O0bFi0/sJmCkkkd9xkfGn4znJbf1jnCS7SjpzbaRWCU0VT+
Vu/WaWO0hI2bJsidD/yThybYUR9mCVKeh4bxbhCA2CqmN8zGaOfO6W7Qc/rk5xJNA4cSuLIlPIEO
LwZnm7ZO1n/oEtZaKLC6Pbmsum/B8nN/bSkgFWRMLmU+gHaxSZZKDl6S3CbnZ0/I8TUASA0jYuUY
QDZ4f/2KmYgn4Zlua+qbu2HHt+XhIu2ABnhLB7dHNQ2urGN7aVxwPbCXtP4gHQo1Kex51S5aWCwl
lKCFL4ay8jR7N2urcbKIXsL1XHA+6HYtK16WEV+/gaYXmtXL+GLetKOauJkhUTLjSHJnQliduCco
A7Rj7aqBrWIf3WI6gi9i7do5KgM8BY/en9vD/u/0mYbAYsv3E+OgHP3Qas9ctvS4bXpOdMluT4k9
bry1qDRKsfh+yeyO2nmDRm4vjXZu2Vbfl1yd77RM030UnW1S6DbJeQdyvt7PP3AYsZbT6hhymicO
nlEhEju8U99eRRVLh1P4R3ch6H/LxLY/ZrR4t3kgMS3gE1HsmZdNvKCWanrYoteT1H5qNU/OfxyH
f8ExHtNVHSgWGwdxpyZn5t0f+WfAT00Ug86tvQY7Ks+DKw/q5Tr9cInu+gs4vBBZdW2xyEGvdxs9
8h/ECK4SAf4gM/wblZWQCrvDY+5gAD9JYKZkdmKsoCTzoS9z43ZCR4FLq+L6VP9MxBtmFFHigteV
lNp+muVmrvMude2i7hLsxalUftfnZFdsI9Mt14b7rw1BKeb/nF2O4r7/bUNxqw4arDBfeuhDF9aO
llmrx94yBLy90l7CWLcpFLFNqCsYLavxt8j7WTXVQviFY0jF4AvU40I25jpvFp5jHTs3fzvuA380
k17N7VwYlEAIjBH6XVzBFU7LxPNY30yzcQsqxaYLDhrLJ4kOgu7wnBcfTUmgUDT9dzezWzR3SQwX
WKUjrNmiGYCFOgFbnscOsij91KLs/JNqA/fse6inIgv0h5HyRUmyHM76XO59KSta7GLfj0/Ae7Oh
DFDtXaujjMZPT/iimr9a4l4eory/F8rGcI5DgJmdQZE2N6nDhWpq6AdUI07n2JuinjPWPVCdbLIp
uneaIxbQ78+r6pzTGtzedb4Zs0eaG79K0LeISKR+C+8XpoeLVxE9ruJNKqldwWauKq/rzrfpwkdB
gvicqBfJYLE1ZyPoYx+l5VV1m4njO0qztn0RWQCYPutvVaTqCzle4NQfgQ49/YOt3ohPWvFBHvmt
JBsawz6NZuPnmtry8E2s9mrVwZ62rBVEA6tPfm4fvqI1KrYGvAX8XoNENKm9gmxPwd5Re9xILtXG
FSu0lYHxfmoHcNDKJa2cy0ovchwc53lnbTwSXpwBxAH1mRldnFK6pyPoQsEGW7L5/BprKbMAvOqN
aojheUOxkgy3R/6eG6RwWAmQ0x1F5D3fwbMnuuA31zxTy6XwVZkf0X7eIaOBDoIvVm7v7Mvu+vi/
mBskPxjYIsvwdV/NsB3WhYazf0RcMH1Rlkcrf6NxjZMxrtlpG0usBuwaflhbWkEr0LwhPcuRKPjW
XZNpTqgieH5oJ8ethdYHVFsYIdvlitliJ4wXHoy+KTAx12zI8aHJtpvTKHwwIWgpJuhCOq2YS3p0
+2GanLE39kVLNA7hrul2n9HDR7iX8Kb65hBwvnHU1L5dsyA9KmwT81Z0RHSe2x+rY5YuQ+FJuZaJ
ETO9j1BahViPJkK7Dp62yG1VH1VyhH0WsN1m4OR9Cyxs/vue9QmLab2TVZDELafnIIO27l9Umkzi
19R9hDhPcrOUGYLn8YfIriF/avAJdczlR++cVAFswRA/vxwBkj85EP/1wvpKzhv6ftay5D5vo+rK
AWLk4NL2DPHfX785XJZKq0NxynCL/i48XybaAdtDllPKjrfnHAJDMBy2vXqTInERwh+6MxtIioEZ
F7kBDhz13TEV52jiQXJbZAs3XdX9f7ZVjkWL7WZw9+DzThUyDCH5NQnm8G4am43MVtmIu2iSAjtj
j34jjd2lMC0gzCNRJoee13dK9u7UwF86CW4tU/9IxP5zJwtF3z90I+3Ae5Jp43/hriVNXruoQXWP
1FscyVCLGtotaRvkfK62h3K6F5bIURZhX1MAGkt4Kd+zMbntMcgh3QYSyIRY0J7MsiCSAw2Ichnv
/3CJ944Fy0rVpuyLgFIdQ7aFxnRkIUTB4vPqvDlHhfVe0RXa2rp4Gbvwk1c4GVlwWSmNOslX0MEY
+roP3KfxQMWXOFMcT4xiLYPgRcjKV76F+V9jfI/Q4QAraWQlesIl7OLSoqj3CvgkDJts2BKVBWz4
SVNovgK8ptIMgj+zEt+qpBMjjWI4D17mQVySmRcNv10F+mWbaR6WdyhOoK8XLhIoKcstn7Clnvxm
fagfPWldEsyDuU070JZ/jXcrKVSbdDvtSHnoJDqSNu6PXKIPd/kXV6xWq3AhKWwuR957UvP9qmNr
I9AXj7lfgyO4KIb6DyLOh/W2snn+3SYoHpYFN/5m8GzWooxJKv4X9cfM5EIODdmG2OoZlNOr7987
/1qh/fCFOULtz5D6CsAERi2mkZcgh/hNs3dfWm6e4au8SXRhEKIhFy+fnQCcPDAxS65cNiRYeoPL
BnV92DW/MW05FfHRr/t/QuDR0C809iW3WSGx523/MX6V5cNkkw5ecI+4j6pKKmhqcbizqzfQzYzH
SdeTslDpWxZPU86k2HMPvWUFv2fH7V13ESDjzRAUHjIWKxwNgSn+fhwaHHzxyCzgrnmidTtGMuVh
cxq5izUdIOcS2KlwzuUIXt9hMHxNm888bGx0xQEWgUhhi43ihA/2ORujTyzJ9kfxVZdpwatVpuAF
KEj96jBcRXijHHt5aeJ0rIUw86HMKAlydBCo+xVnNBU6+4lAYTy8x37xwN6BFOzhkV6MpgcagGag
r4JAanHbA8lgOnATVeupiZ3F6nx/S3CNr3COtwMeXR4XOWHYM6GN3I5do+1bSUD3wjwIYhQPw4Ex
09VldicplpM5eH8VEZI2ee533JEdz+08XJhy2n1KmDI7eRcY3J7XiAWS4F4H+emNS3wYAoNt8LMM
Pw3NurxhQGLsbjAYklox0Ov7FWI+/wfmrmKMpbU23yJ3l04veo7pCgABjFNmXA+9y0bLVN+/m4bz
hcB/DIVMdCQe09ZhsOYhSnM0mh5mT+zayrT70XapOkaCbNOWnrBM5WWVkhyPveNKAa3M7mjuelh2
hKMmQYiK5bT0T61n1hJrsBHA6EfKKIU8sBKXCYwtgqEI1ZdUhBz/SEpb0tBlwDjUKaoZW/H3283i
J37VSGCMNxkenrvK7CUJCveCC7661A8PuUKwXo0G2ta3CF4mThjhvbsdAh48WgM6UbYsJwQ1EkgS
3PPVZNFyDR2KdqPpeiYBlcGj/nB2DJjl1UOT9F/KFywgiD8/LH2X5XNZp69yY/akW2IqoWjjyoC+
hB30kFppCLXjOH4z41V97HAo1t9B1XG5zLNiWDkzSVgRwMooncFFNOcP06lizbNmRjO+O/USbzXe
lz9jZ+zDtZehcCNUWAk6Z66prEKdJqr5lIroTPC7JS61wptsI2qOdOXsD3zL2O7tCy8PNqlPfhNb
3GGmcbYt7I4h5aQz34rHIkWKqljMgvwIUmvyDbzv9gRpJkcwEQLNslMoKoUvGMRIGHll1fjKl4Gm
Z8N/bBnjKkcsp8vEVjRUdJ8x4Pl7LHfuLQOQcINuTw44dd07aNljNfYE9njTYcNf8ev0zbaasj0y
s/821UsfbnUKeeFh5vwmKFhRS+J0MwwatzDHEvQqoOaposuTzTIWwfZWNK/V2xAf683xToAwkBYF
Ootugox/9fusZruIX3csVicTHGyTqtIP89sVrV5bdt6QAl1B2om/hVHL6IOeQh7PZVpBXu/B+OM2
8r0ORTZr8ANtvg76HJSuk3n+FCBQblOfBjxBnnZf2Jg76QjsCFM7YWaa26BtNleLnSvCWsNrad05
nfevl9A4+blKJkRe60wEBFi7gmoa/gM2N8W0TV5XvwtCK9bpqrAw1FPghroRKB/dnCjwjHTnmfoT
v+cdJJnyO+4YmVRADA4Aw/u2HTGQvpmFladCWmTJnLOVBj21VdKDgboLq7EnPeduu2d0tSAZEoHX
g3FWsJb9NEwrjC2cKjzCTrz6S7r0qkstzkhIG9HHUQ363S0c81lcUj0mg0BIW9H+eFK9V8weXUCP
qxxel2Z/QLDgkND2jQm/3o3kDFVyVC+W0YNXSrVb+nOWNtoUSWTbSAx57vweXtzDSS4tPEt9SuPL
ZRbNB+U1QLVF2cNGJ3ugfmUiUVhqWWPM+1Mrm3Aeifsp0zxJYALpPZl7ceQDAcw0uKAaLggCrQKg
OcP/yss6eMiuz6Ad6LFm6Wo9vjQajVjMR8XfzOGHT0/1EnGVi7nRfT8tWnccTYLBqP2BNcUEMXXb
JXv7788Ja0IErkDlKVMIl+14XvLrWDWFZNUCj0mSN1ZX17lsN671J8CervhNK/2dxNKYj9AcZGFS
QlsDK0amOFfvJ5q+TkXl0N+ERINT899Lgubm7eUokmmdR3E+xRNr0dOlaDNJfl7bzIZq7yMTmySu
20me67zq7GV3BbWrAWcvb6ZjHs8S9AO1ENyGZD77JY6Vtqo/vD7pJnRCIlVcVJ9rM1ycToeKAs0y
AfRpbfji8diVZQmTHTq9cYu6kC83p3hPtFOgB+AVrVhE8VhraqJ+h+37XVHOAMFG0jBvN/nvTUxt
yRWxaB1felhEGSAqXyLJM6EaFk07SjzU1WIs/QgEWDFX5OV8uuMnF7LHKeg4hClE9toGpMsVLNnl
oFM9OkRu9IjYwoFEfxfYEY4SOGMK1VvFiCD9u4t/qxSbMB3D6DyAqMOx48nsbCAm5A/qLUUXlGU3
baCR+91ZAwbww43ksur7l8eljGpMolYhWjGG/A1B5A6SzqW7YYpJgYvZlCe42Pv4Pe47o1fb0YyS
xg/fsmYQ3FMrhsMq4WZj2BA0g/3cr6xKkZ2DpvWedAFjFw0mnDxC6AxQqHxqKS5TIGHH67bXs+OQ
KqdYXwzMS/pFyLBTBfXr+ZGr26M1d/Ix4/UHh52DGpcWjFhccgJTOukZ46e3Vqb4mdp05IHEHf+c
ERdzujsKMZ6UjDQF6H2AbHhcl76ccMstbiHWM1ybiqROc7XyMQc+RgO/7MutdJgYsE3n0hmxnwUj
GvKwc1kYG8rAYO2AFPgLeCJFO43KW60nPqs0ben9k3iFUoBocqygk/5c9DD5yRbhgbCoUMErtKqT
jCSPSNoAXhe2uBy1rtLexzKxyxK+h5xaoLB3y37jQjIS4Vcu0IAMPV8fyKtLLBo1tyavwCcETnIe
EmvnNe74MOJV/ZWf2ekXUcK8tFzmxyCsoaXNSPAhspkp3tIL+q1x3YTp86bPrvFK0UOKKCJwZnXd
4yVNQ8ZVXUS0bJXnJYMM2Oq5NIbGH26HYMMsk1nDcRFyehHabhd82DDjQrvMTNou6iw9jCD9wj3Q
afqXSRwE+n3R016xEGSul3qqzDFjMJJ2jM7A/geteyL6inHOe0msmWDX7MNAhZWHpZKsAzZG0vAS
6TPbESKBdQa8o/1lA8U42OyrFpW+q/BNYVj/w7cHfH6Revn9uTfV9ZSdsqPk2j1QGEv6zSWJFEXk
q5SKzw385in954OfdPBuuLxoshJ++1sXnMZRypakh50GNzLUyCDO8EaBj7OXY8DDdDtRLCPQMdxi
Q8LWeKkWGi4Wjawe3Faq8G/Cb7JfiIQmXWqICqZ3BvMEWCq++ERYFrdCrypbPnWhJxdMJImewHhL
LVfSMgXeuclfcac4ZR9z9dPZlTMNQwTxqVBVMdQsUF+43mPq5MKCjIZe7jjUjYuNomsOBcLtv9Dg
0YFSGER59Bqk2Hah/JqX29zpHENpJSCrepXfeD+Ej6jcgrlETGTDw/LLzekiMwQSQvqJn0CCiVEI
qvwQXcUhNzgpvGjR8pLMeQHGeBgTvph2NiTRx786Vf8+9L/+iRan95T7QSt4fFvyi0L4WZxPRQtl
bxkMkLZ5nLNcCF87ThfgWBSTYc3q/R8QRMIkhK2rwNQL2Mmz0JzqBdTLjstH/GwdVHDpaQrR9RHq
GFom4YcwBM+mNspogeF9/mbhUuTGODRR1Nx07HCPXfl8svxWGoiScax2qGde9DLBeg49dpmC4nAd
ZZ4LKqxSvP0PbRP1S9LeIcQOts7vTVU4Wn295tlZSG8A0GR53k9PsLPOWNDkdQorLIAyHIivo6hm
rEjd4QldA0anXu7YlmdQtcgrO/x7UbRQL+Gg2q5f3RFqVGuqhMIEFya2q5g0Zc0DjQU8HPylb3L9
y9HfLIaZU2OLd51HwVgdROkNIs+xjXpFHf7Q0wtLm0iLHccWVw+xNgMAnE0Css2xRZc/i0JdAFwZ
UyheKaxXfsGAEQJGIJlQJSNtfjMpytTPjSJ6PQBRvY0NmYqb5l6kZdGac9ZT0qGKJPvi3xF5ljHk
Dra6ENu2CFosLdx5kdUzD+Zh35ZqaSB43n9hnCETqN8I3neq0QQyZKwJquatOfd9abr2+hH0HCfl
bUA3NHUh+8AgYbBQL0mjDVBKNuOHxTPYf8YTlRhl2Qwwo1IADp5GVHG387f0Oq6h6pjKKdWm8ukb
RZsuQ0PYbzlLbHC7LysJmr+xWraRBAU97156nLAOHAjbjl5PTsBrxn9tZ8Oz4/pU67y9yfpp/G3f
xpg1tymGFRoMX/JbU7NsmvSuujXFgE8B6m6Xoj4P0JqNpPGm/pajoMdZGaYxozVD4a//xp0PNKUV
iGK261B9savNWwV5PMN+IKKO9CbzsKFvHtLA1s89HpZrtz4Xf93fgY9fmfUct+QC1Aff4YE+a7Sb
uHnevyc88vbcWoJrIza7DZ405pU5OfALyQi/hc8mf0djXVLIZ4EUiKkcvweB7yhFVfN+XCGTwSmx
Gar+eXAP2JqBpCHsEDbsQAKjR4ZSjMxbKm8LTYpH5TNq/GuhujBpDuCc0TsbhO1Waav5ADZLGx/k
rqHFFrKE58kUnfjFg6+/wzZ7ziunERzh+E8jz4p5jJHQRP3Q8VKs3+qbzC5VuSzPGEI9WtfMd67Q
a5Q9pjdFbwcxcWtysDgqq+BuDwjxRurZHqv3s96Q1xx6tDjBqVV91Gl2DEyBz+f0gpQFp3qVzB3y
HOu6B6M7piqgvvif5O59TebGg3JnFf3OfCKIp9qbX7tRkgNrOrQyZ+ZbRKK2OVoFOp8mdY6dTHP3
C2yvMJBet2hNVrThuTdSwhOPRLd45jr8MxcY3B0501l1xRY24igyZvEGviDJxxbl1EiSbMkSFJdo
EQjEsD8ycLMkmGyphbnYCoaycSxsUFfEepbnpMj1OvPouLdvBnDPrioOb74Pspkuo+lqYlwcxhHm
6vwRbLNY8EsnZkW3lUnpse22Bk8BUtMa1Vl1QMv9e53HCbULgt0sX4UALE+/hqaa/c5b8dWsKq4L
6Qtju3Qn1V7ZlprbZxOzDTcy/0QRh0S8X7zufaVFrrfDJ/wsJpJrLbVcz0qTcj7S4uDOEZ/JN1H3
sgXscZML05UZLeBTaCs1Qq+ynTHL38RPYg+Yts4Zz7JzV0lH/4mxMfJLSHL0/5SYaIQ0OlV9sq5p
y5tGAK/AfR7RDf6ZLsSBgFkS7CTtB4MIMOP/hDilvSZLAQDjgFrH2UuzcON8AIsJSQuDMx7lnZ6k
PZvojyalO5SBX103X6RVtkzOwqGSP6N4Eap8BPWhP0gfEds1C8CCM3L7r4xRK0U2D1wcHbPyPK33
u/3PFjYlNnsbdpALNsykbMQOvFFUWUVi7H/L5gPxw6jwEuyON9dXTgS/jvEJSG86+UGnUN0Qzk+X
UlhmXjjOCrfIPsPxZPX1DMiezzKjKDFLjeFCl7n5tLfmVItN4dbnD3d8vby1OF7ByZrp0bg41TE/
+5jCSOAqHymxkNq+skSkwyzOFO/SI5dijVNfDB+m72nlXZWtpnN/7SsB7HWdZjzh1P2gdLWlEFxj
dkCjrOjdLp0XLJPxAgEK8ncKKbBXvZN3frcmTZEvImoocek5YYaB076r/V7+MZSEhB8NQYcsM4QP
QyA4Ri+sWuG2FI7DbX/F6e1rAkPz1l5AEe0d7JCBsSFhEfTkzeSTCRqjHmz5b9Ej+FmWz9QExejr
YErUddV21fw/sqEGL4GkaV/y9Sd8iZa9MevbMHHZBG0SZ783LcFb0irXrc/UKsyY7vLyByUH6WQc
+jk8+p1ufLTUZfsz4HE6jYsY8kKThCURaL/UOk+yIZ9yQ+R2vUFS+NFvob8gMRDWfTBagCzoxohE
ewR0hMVlCZ7lkNSuxLPnQGPbzufiZU1FgD6ZtYswjPCmES00MqBb+JHP13L4Zo2mnPM75eiVJF7x
Nb7P9lxLade3QEmDk7AFizeivyukg1tFhs3v2WwDivaw1OwdZY+iCj/P1Iz+b5SwYLCTVLl99Ucg
An5DnN6zkVjLHmC+87CJaFtBArMVqQJGL60lo8gBxTh9+OFLqTX0d3VsUqWamtf/HnWu31Kd8d8v
SMCYUe662wh+eyJMH2EjthW7G5Saaagp2ELv4NUHryWk6uUoUgvv+7FW0bQgzHfReL7vtkNQW6V/
HgLeGqDQHhwtkmO0B2njLBVo4jBCYRji7g/7dXcrujBDT4gpuo4RYjyFwGD4ch1hSdx6fLEShGB6
/M3B8lBbLX1n2zVKSGPsb0CM+sYJv+GsLtoJDWO7txdcxc8mhBVk/2C4m0dGlkRVs1FHGb3I0N2y
9rU0l/50Dlx3anm9zbUESEdPbuLBNfSHeavaAWGDirEd38LnHclm6kcy4d3Z6Agl4G380YYf6z7o
3eA1OMthqCDK6lhzvTR3HMseRUVNahcN2GJvYXrwr0H7CJIkBRYJojvVLMAHevnBUHbeS6Jl5DTB
teFshVOdgVLbwePJ/DbxysZKBmKrle/IpGm1Hb2h5O5SO6FZjeu6xBskwng6iMvhNo2gm59UU8Ww
JyWLWwBppGm6g+vK2hesvEW2URKhgpXTRx1Mng9CeyhC+xKoiOqrtRnPjNowrzD2XgT61qtGYPdL
xJs1LLiuLuWRPJfZ7n4nO8+olThBclbm/i1FUrgjrLzmAKaIeaceMPmCUnxu9z+ROwa+mX3VgkTH
W9vdDJw+pNTe2tAEV6XTqeTYdBPeMC6MJBa+9dqvm3VrmlzWlTbRZmaJROlC5WxAZZ/KdQEwp8lY
24GY/6rZqzczpoTf9NqNoHEzNHvhgST0wczmIVD1ZG5krWfOveeWW8YuEIDcxcWKMxOmqZnC/1W/
A44P4a6JDzZJOMWP8C875rB3olCHOI/eCjT2+4whA7GWYqT4wMbZmI01Ckx6PeBgaB1y25gMoBL3
EnyRfvfOPzbPM33Fdjnb1QYdy4YEjui40LBQeBcGlcKAzr4FXd3pSBg0fSbkMakbeT0sCQhFNb1c
DQmVVOLbKgzi5RUmz89gif/bo90Tt0yWO04JFqtoKxR+h29JPjHRKpBkxdrVcJ7l2cW9s8DN43VJ
PLWi3wnVj9JOIAzHmH/0GUVSXPbJICqqiEqRdF4FIyDxrW2EOOOy0gD1ePz0Z5cSv9KHFQP95b0z
1L+bjoUaj151Pfi0jsQKG8tQ6S/mcwIHqWBlDFZoHyCW63njxCDuczPwak/GBUR3heZceoHi82Jp
AwXxRJwNazc9EhYmTEUvY8anhRU7u/81sy3YOjtmrOlWEeeJNm3P9GVSvbuZHtsrOrFAq2I2Ry1x
UkXmHaWS5Oo3pl1e/FcRXXwchLG5BHgcSxBCru810oVF3tn9QkkLUZl4kgBTcbHnB3Iz14VjoqXJ
9QnWLrZxwpLH9i7PTR4WCvvp5UnnySt3LfRVgSEHJfqtWC6mjAjU9t3tHFqYAuuMvraP7mmqDCuR
9ChaN8C1n6XeILZbsGgSbzMQ/ss1DbIkiavMAPwMVxrmG/jEOZW77WSFjb6RR996xPVfKl7b1n/C
ZeSRsIxGoKxrh3wgrALdTRc5t5kj6nodc6KLqmUyhq6Oh+CK9m4nlQS2q4xEcUE+OJ49rs9HCDwA
BP+hkf8GGOb5df3hfZUNFQAAcJDCx23tC/QvuTQqzQEegGqyQO6/fYJ9dB+J+EHu9UsD6krZeCt0
R3ZJez76zC5ADXaObEsut8WIRzS6lMO4OQ5cjBBNKAUKZ8d7MwiN4BUYlRroT2Sn9ykZhj260RZE
7eOGmy2jD4eTMJUAI2lIg4yFQt2Bep9OIVyZqZ7kX5fobJwmyTLopWkMefQZzXTBroOBqbFtrNMq
N0n1DxQZh8o6QCHT+O2gNOnkeJPZSkTe9b8Jans+XR0Kf2zeR58dPItjhD+78zRDiIqOI0MrqQGG
vH2SvrVbX0QT9Mpu/6UjhUyWOkhgnSEGLG3H4ipkDFP2MMG9WnTRYJmgFvvjWtXfBKkgQfFtHlKw
70eaFb+33tPVCoV54vlFHi/RH1/dd6V1GSg1kWuYnx/L1dPx9AwI2gknLyhB14dBIWF/ZIC2NerA
gnjzj/zHVw42mMS96YDuQrRTZ/DETmIhNPwuWa6daF2qilbX3qYA+ss6HT6RcxMOKHAnLbu6HHpM
cC7tNlnp4YZ8MyE5jXmmWUHkTXpuM3/Ld1QCARcDyW9aW44UNzlQdzdPLcQQDoJJujP/SZXMRwiZ
MBDgnjm9wKBAMcUY8EdIWMrBfddr/wz1jhOLLed4hDM7Hp9QI1VtUzQCmqj3KebmNttCwPG3srgC
tIyPdvZ5nYDgSSvc9RNGr55VVzWKe9QZ7WBOY1T2xUt2LkvW5lopYnlBDvCCpg8lt2q17aru7dgF
FxMer8ln1FUQsUAHOnhC/Bm/DJ/+SJaUmDeFxedapqL4d+x6KuPdWmDq+TUrCghNmwCyP5A98GJR
y423RiI2zl2RB1UrXc3ubvE5+ioHFqQt7ENkQll+f8N0RXh0DM39qVB6S5hFRXA67Gxok5vBZiu1
obqfHolZfhriS2Lr0+202oJmgUmfnbBhYzLKluAgJAleBN845zGR2c4pOcmoYcfr2AiwAcMWVwnA
8kvn7+e0m5kTWQCKTBXZxgzW5pKMerVPc9mFz8mqlardFchM87sm6hB8XsaoLGnRrTfX84d82kT3
5GYX0bBQGpXOotZ1j4H2HY/mproDO1Z2o2dLAMDS5+qotzWauvIiPK8RT2+V7pH4VRAReNWhv8rr
MnA3UQERSqDsbfRunuythGvPtGz3k+CjhK2VYKxHcXF7tfxHyHRRbCK4KGXN5A2NevCiosOWR4Bw
z2ppU7LVn8zfvADszpb7H98MyrwCB3fe9B7QViTbgy7HVwFfDk5ShKv7v3dSzEAQ5Mb26TLopPpG
dU1RjGZD4Aj4xJDLmUrI1An4G1abeVD9br45ysNjxWb1k7JQ/OxqgUbv6Np+Gl27yO84BQKKpWzb
fYNkMnDuE7QVp/jT0ILNHzwnxg27TNG60bjTBfCEL6ZzvzxfBjXQU6maMKviirA9fURdT4sRu5PR
7MnzRncIrup4mGskU7vFOJSBpb5h4M7kD9HsXmsFvD8RxisGNWjjVyZRtlmurJwPNS3E4C2HF0Wa
KjPGiz1u0YJATG21VIGHO6z0Drlx8Hf8hYH/NET8HShahCDQzmswQ6mmH8V21RtdWAPI5aJ1bVnY
yXjZUFAJrF1fqZ84sxabqVFFz0HXkTXDn5XeW5B8En/weFMhk13eXOB79ur6ZlnOF0qc9ehMkt6C
igEROzREWbGqKb89uC8UlHcUbBHjOoeoukHxI2OupIT3SJvBKoky29tAxUJVWYtsQNzqSqcfKmhr
Q1PuyFlU2VAvBQEXIY7caCK/TmipdEV8Ba4iWqsc/ATOEuaQFyX3wUVi0XuQ+qGBBgqBWAPTJ4j2
wZxq59AJhBhYq2DcYQDAR2As1XxV/b52GfFH173n84yo1NoUeukgPg3eQaUrb52W7+ZRz6rnGZR0
m7QmAgDtWFs/lfoL/uJaELG2Kqja52L0j7WKFsb9jUxEaYReuvR6uANAoS6l6JIkRFP1APPTpRXd
23P4w151CH5gHzakeN0P1XIMjJqjR9fYcxks5IZy3Z9QNVdzfHKg2F/h1k9eyrtrCWpAkaiS93xI
n2aQJqigGUyBb6uHkNZdGmQd1wfA+sfc7Wnb1pOAG5byvITHHvdw7C4Cu86gOa01htDR7SOIHepp
TTsgaxKN4s/jgwJ4MkkcRRoVquTgiTGg63yFzQn397JSVx7Ec1qoGjqyaoCXn/qZeRMD/G3hFNWk
4COMvOfna38PfjuBZHSHyhditzm4EtUYW4qItqtlid0OKGImISKnt3d00/6y4kTOA/v0BWrK8SSi
5fJ+7XmIYKC4JnNXAnUXiWwwWWjEe3B9Gwi7MAv8foII7SLLChl6ybOl6o/XjBzIpkPkcqxdHzSB
3znZr4rr/sRWIsaejdI9+VZBZs6pP1YM1mMa4RJopmU9daaRgUN9bShZyMQ2xpLHwVNlHpldDtah
ejJa/DmPjNn+iYdockRMlOoTm0KORdHsg/WCjt6yqNFhLPdZ25rD6Eo6iWf+35OnOVE+QRZ020y5
akZnN4Jvo3aibM3GqAGKNrOHrQ6gkaFz8QNzPXcUkaUhdrMk5FFHYdlVCNZrvxfaXRlBVu8Yne8Z
eEszeaKn4nYF+2vuxSZpAMDtn9s5sSZUCQpq5eJwv4nwtk5h5ba1PK+y3z5hWEQRdut7Rx4hSOop
6a5tUpnUfK/KMvhbOgLkaPKkNnZKCwxclm+8A/ttbAWG/v+UFfkSrgmTwrcnITxvGTtft0UhMYro
PdDvnE/KTxmRlwRJPWhaVNRQcdkXGuxNknnDYli57PMw5VFziFD5vTE+EeWw2dqHyTcxcND0ZYIz
nV7Q4vp5G9zPwY/r80M5tNVoQFfVtmI2oy9D1I65HJMBYco3KGd0/+XcxQvbVi1KHOU6es0mkqag
JdC3aJsHKvkI6ObSCcXei+lkp0l1Zb8rddlVN7llyov9ao3tkDOlOFFvWXcHKD8yDibQLlolrgi9
v3THIc0zs/YX1TORKGRQ8PoyaC8b5pZPZQ99zKuJQiYLYKr9vyKa2awKM0cMRFME815lt3mTDZy/
KfvHsIvA/OmXzqYeTFIgklg4bfL47ZFT1VSdoAuQoeZ0hYPACm4bkA4+plOxiJ+3y/v7DoRiqh0Y
Jy19JNLYVC1TL62KJOIUCNgiL6PlkZTU5b8AzH0KarlxQopO33mnlHyqBy8Q+nju07/Im/OdTXVc
iw5sISRM5naykd9zV5uJBo50EzjPQKgOZq6FWrqIhWSc8tux46Q3+y4KeRzhqySUELdj7+gJQjfQ
nMx6LWLk210m/tmr8DXfjKTzT2g5EbGKZCI4yVunmQfHxVdT0OKCTveDeC0zmAIpeqQrmZd3Zoce
zMAiVufCTDpcWT6lmo4iAf+E5W8a3aUpqnaZQUYVRD9GxcKxFk62hAxpAUfM/Uar/oy36DbCZibw
UP/L4mYgsDL00/88BqLvUFVz65qsRrDv3V3UHGyjhDzQeAnVk79upDwtVGalXzGODF0MgAtJgvSg
JF50xOhsb4pKUDHuCPTb4Znzuf32dYpdOD+gy3o+0r8AbNDpy1XIDu5/rvhWVV9UQ+gguppFY2ZV
3tHJOs56VQkgtL8cZCpEP3EqGH6llvNkbqExftOthPqw53J1jUrOwhj05CsMkOvhWk4AlbPznVYt
pvOGDlWVPeEmeVJeRltY6UDddgFGj1Jo+jKlwnA1pZ6FhUB5BZcGNX1PDu06gLXrW4MHcNeETDwp
E2pk1kT/RWivTIK2EwHsGsiqxhJ6UMx+xSu2kQHPv81T6mxlhf64DcOHzOxeMwGSvZFxbrYM29Sm
iDiy8n80wXqjls9LV8CGlDrU1mPEu5M9YLe4QQtXn/HiFEBac9/u3OkyEkbiFrymMGig9GYyGO4t
9vUo7jOKSy16ybEmlPk9Y09Eb6kOZAUvmNvEU2Yi4vhJiJhypHJY1+rzJ0Cgft0C6mYt7JL7LTKc
CF5hYclInYZfBlWOYv7R8VlJBqdZ8+i7b8oPhhlgS5DFDLPLiSWA5q+qK1MoJ7HE4Y3ScCKOK27T
ydGNlpq9oSx2mOa2ZzAUQgDUDiI3/VJS97Vm3ISxvtiu1fa0SrYQc69gPzbuiCjBjR59ZDrJONgd
f4qvmMs9/Ow9nMfBFH2wh5FUbVau4dtK4hnboS8pBulR2T/ml1H42mzkYNd7NrCkDYIqjJ6/3GVm
xj6lhsfRC/XwWfhrrbXJ/IqZ6jzQx4FAjH2YEfBChhAUhHoHctvVzY+y4v3BzI2QW6SXBaSqPvdK
ZsBEzuIAJN2gXHZktma6CjW6G8wLVnR42UUQg0rTTAQs/8nBUy8EdvhCrSuu3MJ7kk01un8FqNHA
dvdksi+tve4HdArzaqN3MCItczWxhmfPKO+U7Vyd7OTQE+qaGR8Ys9IZeyQw7JVh6tpExfOOAFmG
trS3hxrfYCXuLvRr+8uMM696LA8P3YspWZP5ekDmE9sE6Ntm4zDnOFfOFVTkaaXphtNroVksxV3/
mkaEJaFTWEIJKGKh9iUCcg5YvfXdWlNtwue7clN5hId0Uf9hjVgKP00TcPKKE5aUNYxkg9TZMyOs
clqjzsYYeYF/ookqMyK/UgQ4b2htQs5xVWuCromSie/RJeRCgHiM8b5HIe+DsE9Cl7si++sRNSDk
AKSalGrQPBV+eU7Xe6X0O3pTW4Y33yubm9z3fTcgIKJjog1cKNSvk1HT2PupFf6FEkf8DJiedYFb
r6ky5NpwBM5H8rAYW85cW2FnODhg/h1+mXbmbmjQPUJx0FkkqjaSTJG1AZjq4mPAXN0XOmY4QL6F
1hMiYhDmbxSjYl2rTTXPHauXH8F6S9mqD95IbDf0ou0gB6cBcQ5VZK62Kc03XB26PHAjMmv2HksD
ueFaCN3fWK6NLOquYVyXBGIdyb2bOpNpfljsftYbeEgtHiEz7P/2vF+sATS9wv4wdV1SPgk9CGGd
2UhZZibKmvJNkB6HfApEnD4C00jK+qFktfEwMI6LBfPQWY+97gBM64p+f4BE1e0yvmLpPnW8fZr5
GHZDVTri8swnb4NUv9OBCwBWTo+G8t9CNu52INe0OR0CCLkeuyV4T3+PhgPe7KG2lR9Rn8wVvMeo
mgSzb83CQBmvHZ3kL9Qdt8qEL/HlZaiBS9Dfvjli8Mh8Avn5s6dVdhIxEAkbpVr67cg9S9tiBDrC
5hjq9tD5pmjoTezTaO6YvyNZDwYT0xpduFgEgn6TXtqTn0/3eVN+bAxoZGgYgKf3NVTk8daO7elB
rJq2V6boj5GfxXbDloFaQX4bo0z0ldvw3tSONZ0rUruuTKYxTWzntMlcx7mqQ/klts4jgC3CO5TS
HbcvTp1MsY+88278axPcKp6Jn/88BIKxINe87B4HdE+TpejWICe2l9kTn4n6lRxcKfm2kQBqQvEZ
d2zE4u5ZbHXw3mRrBnBabTPYgWFA37p7tProwUeFFdGcv3Gu972yHln4aHqSzH3FMzhe6yJp18gs
69MxcPm/hhbM7lEqdpc1qu8N4UHdC/Mn3s6GdmBQCQnvmLD+vbMQ5VBY+2NdgXdJrcx4vJrydbXz
JTGDmuwoodjbJdTd2qVW5VmtnbFi75+AcZPk7AcuFtoOh4CKeRMU1mB7cpv9xKJaP1e2c8+sWATo
w3h3E8qjmom3vDl2LBho3e/qqFGYSg4vaYZllimoMeQGbIY4rsct0JqrWkqC+nfSV/g6Mu0PyOKU
VKOPMj4A5pONTLIiTojmKBw3gxut51F8F4ptkFCAbNdcyYbNkemAd5E2gapgX/TATeql3G3dstRK
w09ht9QH7VRokUPtuEtUesmg46L50RuFY6ANFso7KbcGTYhmZRG4UIn0biaxtTTgEJGxcCkJHBPk
VJ5E0HIBiUNmXnjClsU0eZBa8cr8nVXgm/Ya0UX/wgKhVI0exgnOvyGGcFSTVbi8zTrsqHl8XR27
lTek5ahM6iTpeICT6htRDcuu89PqcFSwNKvoPGBdPtCZ9NjyadfS+NqbFT15rMgcjQ4Lnsdpwfcg
35Cta9RCJbF3hCaVGhBeYISMiffdjYMr/TkYUG4TfAJDmr3fsFGLdAPgIsHrK2gfbT15MgZKtQrG
If8LmxVq/N7Lynsa32SAgP3whtrpckiHdmS5ql9s2SMFLAeH6J00U6ewQZlrlXeV1HwkWQDMUhdT
BDPHy2jKe5FHsVsuLpbyeuslPNDI1BX/oLTI4qp5SbII2pVuA4r0p7HUpcJnxcq4rEFnxN5k91GQ
BRBH4I34Tz3F8FwNOh2zjXGlzMLO5iqUjm0eaOEmhtyXtzwuMMoyi2EeOhCOzz7vl3flrQHXYS1Q
+ccELYkuO3TRt22/o/50HC/60yt2vwIXhh+pWMdgDZPyhCdKqHO5XYlmhDptIj1Eu4YTyGmRO0MC
TSAX2ZcVEwyKQT5iIdvLv2sRAabDNr6xNwqSMxWjo3RnWUbPoiqYSGiXv0slf6WRRGyvzhfnwnky
su+F7gvSfdhoqhX42YzYnwfqx1kfeCsUf7vtMQTApK91t8nB4pqnrofpS7MiGkcVi79LQJINDcPJ
Y9d93cc/uY5laTk+/bT7VaEtXTAFzHj9Yo9FrTSdJBpn0GNFmNr/YGO4yrLzw9VgLDgp4rcgz9YV
e5lQUi2VEJU/PUyOv5pko4QsP+lcvqsQD/C7clNDE1NiuZllZnllnQ9HmbfFND25RiPJifyDhlcF
fS/pMOdUEZw80HQZuGbAC4GNfJ2XyFk8vT8kBm4aHAjfad9ILVj32bnkv9uGPL6hA6v+Qqy4Mmkk
z9GaLpTunnUwODp1uMxkuuQKS39Unsc+bi3W88BYotNLDuoq8EK0M2TfE+crq9xkfUDQxSJWJ6CG
VWL1x+tGdDPSJFMMo77scAvWGv7WzgzYufuPkNySo56ASRXepdV1QJcX0oWgMEDa1J5oR/ZrZPjy
kl5IbD8E8swH4Umo0loaVEcu4XXLvBThg1uPZRq3IcHyFnbq+MpZNXQR+beqQOH6s4tQMLxieZFC
AxhT7T+0mzh55kigtqMNHecR9c3/I92DdBBQ/jS6pDJFa5tYP5FGVpZb0pJ6hPEADBRc9BaU+Efz
3gJMXJYz4ldihTglsIukjViEQBAM9shAfkyvU3jkNnAWbEIN4qF4hNp6LlpEpugcU8XG8YZa4gOE
CTVdw5Gc0bgPKZhj9dg5flP9XWm78v4aDuQemA8dyNBjIUHfkMKwlzk+tVytQjM33PHwhj2ARg61
FC7wENyjp23J6+QE+RIfPBjuvWeIowzcnNIijtSEAiRBw7RMt+7dkPqlsmjn8o3CMdBok1xZTYhn
fE8c0Co2s5lD6R9ekNBzE0wCFBIzuGaVV5m2BKKoZS+s+WWrKbrn15Ij26LCSf/jkMjenB9Uiz9q
fToBZpymvu3weJcLTpUlrdaOSEYoiyZ5w3c0USraBs+lLe9Y6X3SBQGZh3i1g3JNGv+Wi/GSGXiZ
Re+HBZ0+FvyPPmMA9iLGnZH8UTbyzIp1NBru1azexDcRNAgYJuNMJ15xQBWB7S7K+zEJP0HmnGI4
UxePP2DUPNWZJoEayqzwmKXJdEPMThLgl4jiP2B477znmhTxBhOgl7XLdr6U3Mx4I6NApusp6QzW
RG+g1MubUDZHdVXIWx15L2QiJqRrzT9DQI17O3nc72698iEQO0gzr0lDdb8jA6kArefgreh8ZiVL
sJfHFCeJkPPdBC7CF7H36W8z17cms6sEey+roxFZpfJk3JPhDJSHhpyCPGdnlxWXB70cTTUpScLO
bBswAfNo4YdPxI6gd4hj8KzU0O/gx7ZMwP3yMXVVvxgkzsVLkKf4z19aGg0WZxc1p3ebLTrQFuZz
0hekH0IBWjhz5PzFbdZZhGeR0JjFei4SXqh0mBPQ4lyVXNat9IqNeQqA8i1zqSJ5ZvAjw+2T9woJ
kN+HafXhs9WiJ84TYECRSex0e3oM7xrcBFVXgyw9mzpCFFkBoJQCmJ/jeHKuG0fLwmqJ2ms1CSn3
Ch65aq5MWonorQLu7OCPhlLEkcZ0ZGfmsp5BnTWrlZlC0ZWsPl9adb9jBXPqgtrAcUyjlKuBisre
ROD8gi7zKGz36ncSL6bBQj2/sp/H/ZtFAtiMALbr53R3HMNSne4dK1lHxy0pLAYrBGjezYER6qwM
/n7ZukdoeJYRAXV+kyQAGayC55xEYZd5UGDNbHNgZW6YvtpKNMsUnNJGjjDCqEhagjrzOnlWhxot
F14ujh3XY6BRy2oCNGgKK9mO4Jg2OQfRHAwU4gk8vDdgI7FIV0PhhXXPCg3qVwXuGdYAh6Dz5vje
U9Q5JtFy4Fcde7SU+ssAcyJ4A+vcsaXUcazQJYr99YmYYPMFqpQRbTRpLv3wd87ooU8Rxr2qrjz8
L1F2iLt/pbnK5LD8hTPxa2V9DLTyDPNTSsxinyv0eptiVCJ6cDjaD8S4TQ9T6pctyvgxgOkOSh/7
1eaetkAfc1KHKBEZuHjm7uDvL5ZCWRd1tKy0Dws0fwut6jbjAvUW6BpBWMoj9G7p1AHOKdx+Ehyn
F6dCWesaUR6Zm8jHHrILR5bvplEhCe9KEH35CboQk9YA9WdBdlHKTqjuPJAFHUfDCE86iv/P7Ktl
Zr/u86qeUFVVWM2B2ytDOCtcWOuxDgQVtlOTOORpWtuCyonXgMzjqa4bFjwUDjIeHk/1CCyUzcNH
xOgiOHvG0Qxbu/ItqdI2g/9mVYYCShGHPecN7watGo8hjz2yrhwFSfjxtiB2k4pRDsVI0ncM+wXL
5DHHPrnC0VoZThXso7y7RXLmXeKf5qHSaRlq7x8uZPSYjEjv2KqM4vuXhPLmDxzM1bNOygAYnYM/
spYkdWbtb2vs08YKfeRhMp4kpOZ6gzJNXJBqGCcqaGgnI8HLdgl2y8vSQZPzeBndlmVIHssgZIUR
GAHIWxu5HYvm9kYJWqEl/PyAjHQVFaktjCgBpacZoSLX9g4kb1wUyNsB5PQnue6LlSw+5uYbmPwx
pZQrv3gn7153Kpzzo7ekww1emeuvkvmTnB39lx5rCLzR6f7mCZUV3udqkly3g7czrkjizUyZMXWc
4NXogYNVTiGiwL1fewjSOEp3Rq8V28zGzr+l+Is3y9mR+PBtTuFjMJ2LSjDsA91lvY5ELM0sEXCm
bL/uNpaJYU7dWQHYFPdt+WMoGzLuk9wvVVvLWH2DaHUNntUDx6+11CFhoDZ4E1jbh+opio5punW5
2MksixVIejgjwlU8xv/TVzldt80EI+NMmbmRdZ1z76nLA9wpJPkqt2Lfn+tKU6/iRBZPraIFO8PO
ZhtOG/YRjJ8McRUa8NctIt7qtmVCH8wXz4h5VDgmxVaIoapRv5Ol5vBMUKXUIhy8rDby/DgxGX/j
ehi3e0S4fMwHNY5uRrSy/PP6jY8eyHTkKXO4npmvNrpU+Yh4c4Gx/hOk4Xv97wiFIWoayIv4R9TA
vORa5cuWm1zfFQI9oICOoi/fcp28+zLTm+Jm8+QzTVhhxUiI1i6VUtsuvsfPz/EOBN0Pehp+q28P
ZsRzRRq9M83vkuRgT1vyl0aVwSkuiFNWAXLLAAW78Wj+3EdsyPvEE+kz5e7lUQgnchujt3uwO+u9
aDHQKqk0Bip4ZcS3Io6gQ73qPhDX8tPui3xe15hUVN1yh9nUK+c9EqQzxmI5bxSSBBd8y98zIs2T
/xVXWb69TvZw6eC47p5OLEOsY5NNaz0nBurbXUkO84PfMwjxPYQuri/yMSRQFwT4YU78wed+DNQ6
Ko1eDcS//odhJfEgwZNc9CX/pxIhHw/KT8fqrfEkit/r0hpM3Oakiv5T2jqUX6ULGMf0CJ0BbYY+
+XTxjdbDYyMertIVaQShQZj2eZPhY2Jur/oq//r+UriuRnBE+zUfSCO6tceZzHNa5IaVnKyQFkZb
7R4ZdB8I26+j8xFVGzMACRgMiCWV6lMjqwv8xjSMaCbmTi+RxoxOhtbwWYy48xakrg2tpCS8TfiN
vAHWk4UPUAQGG4PprTsrXgTRgEWtfr9/UbgQKdnvtFDCOvt9PfbVHp0lSen0G95MGlotCXr1ZLrQ
HbZRpO/3AxiHzfCOSw2rJWE7w4ogbr6RuiMoXHQRG8aazKmrxTxuH67XoYGFJ1O/v1PB2+SCtO4N
Eu9yEcs0WAGnADD47skFneo8eFUTNzGggC0O+bpKL5luS8NNIJfhVtL0oAsW7o7wLukz1+Ge4zDD
FBydO7osfSmcPzazHH++M4RhsvIYocyKx806ihgwnm/Ve30X09g7c0MKtd5kRwiPPGJVUra8LOH7
5R9Au7lcHq3513w5/XZd0vTg425skNkx5S3BCIse6uJJRucWfQfW70X611frNKy83nwfTLco0heA
JYj3ja21TmTm+M0bA/y2vx48/wGa8r6CqgctpWKUoLHb04JVJGB9qxa8mSZrmB7/G2A6GfqMH/WL
UbnLPag4E6PcGG8UyNeH1MEK68q9inioTLCfGsfdE0fkT3h8q4LAQMPtZbLvZMXsdGEls3sQq9sl
kC5s0eifCFzpPmEiVdUm0Anyb8mgKC8aYqzOWF4QJaq4cl49aB7ZquLfx9louMUKPzXWD/EW0EVr
hLuhO3ClM3Qvg5b0Jr5FqpwXUUoxeqHEvM+Pn6r8vXharezX8PPlxXyUimtv0oERyvVbELk5XITZ
GJG8DNRnr+ye0GtjZpB1b1+YKjfhLjvRTxjJLRFL4ZNha3Y4MuAs9W1Zy2q7xkTSfu4vhUwXt8QZ
YtamT1rFd/XGHlb3qZW3lRicm5M9TJFB3rfgeU5Gr2NXNeVqyzbZCkMBXRGJLM1t+7mZ9PwcBQyg
x5c0n0vLCS3s19wt0yE5IM4HFC5r2rBdhHVa9SRUMNdVOSVc74DZ++rMOeUyCOak9939g//jG+4v
2vV8MUl+5IyD59z8sWIstaxJ9SD26kiCcKTGr+Cmgw7urbJ7Dj+PKQKCUYPb3ujfijZfx5I5kMCt
lTgaJZwbm3eWDZy0kZ2TQrEkFlktJ9ErEh7tZZcm9POv3JnFus30fcPBY0mxq03LZAlF8riAoIZR
59cvVzituoJ6Ovyiz2sISPZnl/+mP0FeWFNudCgRfwHbL1xGj9bvD1sg9jhH0ZewyOh34lYfNyOM
aqY9IRxdYR53byjhYB+1bbPPlU/oIfwbWJaSfJWUuGmHC5dPBz9jsdViVtgyLNeH0/6pNY2hmJa9
6am8mqvqDwaQBcoI3wU9Hz0P+v87R1R1/u2HehGzbQP005ykbHpDVZEqIBkYr1vWxWi1NoPjDks3
TsCWFgCFhXTiCI3xw+lupAsR/BD1VOwPC01GAzW7+a+F22SwlvOdGuhjlXcTe/7haWVqC5bSt/YN
f9GG2ibeA/VRWlGjUqoupKu9eyKvAh5gM7jMn3Zz32+MDWJTO1oqhUOGX5CaWPxRbI9A7QTsvYOg
keSLk8LGextcoBw2vCW4iNoZWjcjbeHzVlMqx6CkKd1y2x9oMxWiuf4QHtX6D3+td9ygTysA6fXK
voMMOF1J+KDzeBthm7nJgFhoSp+90hC/lIb7keF7Z8RQRMLhIwLBy+JOOkzn3ZyPOHvdiaRDBB2+
odi/TQnYGyuMK7Svkk6abN5U/b5NL7/GvOXVuDb0lW70H8HLKIXUeWE6Y6swBLw0D0tz/ONUJl0e
CM+TNJybJ2mCPWqZnIc91auvJA3tmOIr7quRt09L03IXXfHRUtiPuNDDCZuo2+2cZejmJHkje2jb
dQdliNoBRmKWzbIWTXedsjnipSgQu2/xRT+zMJiNbcZqtVf0ju/Ked50NwGXIcrEB09B6B1UzoLP
pg1x6Og93apD9C7YuNyJHJsMQuOYyj+wzNEX30Q0voS9hhnWfLGyMs60XSWexeCjk2x4i4VK7nMS
VSPOSje3ZaakyfEjbTo5XwQ42s+h1tmhET6WN+VFjRJM4UYLZ6w9UGejw5Rt+iBO7DWTnhdGZIKZ
1rBHB/TN1fKd4Qaq5alGzs7DGzfcoYRsjw1WBzdh5ydccp/X71jMKX64ar1bqNNj9CS47bfthIpj
FQNNcj2M+RmE/aYXeWFHycFkTRs2VYi9R1o/rcJiPNSI23/9RyyRLWHOtyELNn8dWn4U+6SAA7YV
/SAalpyrExTJIgHS4EUDrxXi6iel+FFRlkM3vWulEFVB2ockIklUyWmyKl0JuUP7zB8RNCuLKuVH
VZO5kcQdqTY5gxH7hHiDuaGlFz79pxhDpoggKJ+kxgHjL58/mXICSymB/nKikq2DEQxNcXKW+0n/
nfaw4cMreo3TdBYaLMAgifLLldhhy+k5s99a7P/S0fXsghvGoiEbELwwUd+ODm5hkpM+yNQ8ia68
BYfbFzdrpDS3NlU3RJOwEksG2QPVirz3BKOf/X4hWTo96QfPxL5kBPzCcEvdRt7XgRlGZyYzqc/W
GVB+4iINtNhaIg+fG5Xfdf9qTX/tnmsfDx2NBJuB1adC6ahtXaW3LCaiIQvyt0p7ahOohGzwdPZL
lquTB+1hmbmXHvMtDJmAg+4bOo6h8nxWe5hH1splCnZkfwLr1CDj5HMn7G9NeoFlhiC3d0yA4XTn
i3oFhBb40UrjJ7UVQaNuZRR1u/V49y0Cop4tj7qnyLLkl+wKowaiF/z8HFo8ZDvms6PmduazXnzj
ZoyVNFyNdQrwyvfaadqBXwhQPzMf5nYNmLEGz+eU9ECXmuZbwPXGQJ5ZwXTmc6gyjjixCeuuOanw
xpTh6byCBtw/ByvMQkiWZg+wFDhT8Ol0K8+JKFCApc1vtwLe13fYatthOpVT+HzPgZd8Ue1xwDO2
YDpELwjX2C0oUn8NRgge4g1Rj/0yZ2tkxAbN5sPqTyfTCU9t+jOxv7A54ZJ23EfSinTzOpXVvQYF
eqJN2gSphy/t1mGKxFVvSZqlDWYc3D6Yn67d++q4ffwXlyZRw69XxcqO0Tbt6Wg0Z2pK7gqT7S0L
J+pvzVrg1ofzJzjjWbekgrBQywo/yGKS5/rbsaNqfFv0cb0DDmxp0ILlI+YnT9btDMmnaZVWqWZV
OG4wS+8rCuw1SvHZNiWn8Lg5B7bQi+2/s/Y6BbQae9/y91Oc3O61/rFbd5yJDo1DeLYieDjfDbxM
/z99uU12nMgfr9h8u+30ZscarLe6MbeM0znvIkR07H7K2eEtA9DXeBCjako7O934JClivqAwmzp3
VFz/CbmSlFpspjOeGnDEiIEc3sm9O57oubCOHTsj4N4o1W41q6cdnpybOYtdpMqrz7Tj+/saF/HR
g3PDw3LVDebbVugtvWMsUI7ZdKiSSmxrqqf3roeSYIApoaouTGIf9AjIaShrMto954cCUonNYzfo
bWRzngw6C/+D5Up3b8yQd37wT1vPbAlq20eaFEh+Gns4u/2nswDIXL/tTuf778BS8YgNeDp5XbE6
y5D7uKvTQpT+VB7q51vKooWwhvGYrUXHXlEoIrlZ58MYmiKiwxKcOPKwuTOSgs1z0+o3E08jH0JO
7wrzqAJjwZT8vTbM5SwS166DmbEcffJpUxi9VGqYzyKW4CNNnVi0IsmjN0tfQtBDj28xOLRUwSRT
EE64254WlUAuHj46fIvW8p/bEdSlIv8kv4pVFganxS6ih3TCxM0qml2Q60GO18NwKEjOZWps6xNg
tA0E5lvmKQK5vRKxlEaw6zBI/TlqClcKHp3Y3A1JEose5zv5YlEbkCpK7nJXFCmuoxEFLbHXtimP
Pa3wbAAu75kr/untB9ovIjuC9DSU4jN9rwt16o947HpValP1Whtk62RZKUGNUnf+dgT+JbDix0un
bw4sTzChpgi/RRyvnRl/hulBUDYLUd8uCUZr8sA+DrrEJWzdJuwEPvS5YUmoMPKPKpvrfvMaVYaV
BXkdBfxvQXPEJXgO/5F663KK0i+u1E2XY0np0iTzi0Ud1RG4jwrkcI9lqSCvrZB+fyLZKd9Z0ZGG
RU4vDXk5YMFJYhcOEqd4TeZqiOiYHrpE4V8hWuOkBwI0KmwqUnWy8NwEve9xEvV3ERp9Vt6iB29m
66UWReGzDZY6Nc3IYbLb0cWzWIPXZirg2OX0NRA4yVL2cWPStWaLPKJGLIP9PDkGppeHXVe6fo7W
5GXSiDpAMPAdGfnI9UBfLOC8ON8Fb/8lFRLdMRIDmCVYbCvU6F0TR+q7BfHC4y4dMZpePOpHt0lb
+GU1DgewDPV8QV9A17rYW9EOrfsABVLT0eaNwUtdvLMtOExt0/7C92Uq1631BE7wLf9xjV6txjzD
mW6POWRFTqpn432BdhCl+WPi9SUxFXLn8ZHr+aanSqhZF8RuUQoAl1yS9WYpkLrVfAJNDp1nqTTz
RqqhxaGU9bv25r1jYv6Q0fWHP/vbMcWo+nmkcVe2aKUu9LY7aVI2i1+Lfa0JUqPBeU4K+fpK5ryD
MvnQf+jZHW6E96hisbSp84HNylL3W2bkW1S7Jcpa0ZpJ0pUPQ8bdJXfcFpWK/sVVar+Xq9At/F2L
nHXI7LHv7zJ7N+cND5syr23+5ykgZfOM1tqy9ZDWPH/tomfIfA3ZG4yZBenhVvxrh98gGNFEyOHa
Szi7+z5w3scN7dc/vR3D6Yw3pN19X9pkkiohJGAg8x9gYvJGcSwm4m7/UoJHwUUbes3t3LSKt/26
AIxO28ctCQeWSqU/cOdH6Vs5ltTKXjuiyE8kJwRjYrP/UppCuv2sZGur+Gr78DP5jcl1Ax0V3A0Z
XFxVjr6CPRmBRxgVOZNxy6bhPFK2N6xpsPisDBg9ZVsd9FUV4FDzjjyUAuwDqVUfnaczZu05Ji3E
Ww9OFcnGISqQGyL30m+S62AydCO9KQ7qV87E31bGG6yL7AtwJdKpcDGZZkgBdAXKT5ZsJyVGn0Gx
g5K3it6FT+Bz8Miy5PjGd7T0Zkfo+5IDV3dtdGrpqAenxekRsLglsOYnuFr5wAm6fB1+SBRvl+69
fFRMPEpcAHiIvVwRAIpwNkaMk3QztGy1WxGM0q01p1TQYwhn5PZT29o4pRS4GMU+MqcrWtutPk9p
A+azZXlycgv2uNeskACcrjX7k77XYpeHPkxFdpgGBsPIzpmT6spS4IxI4GeT6zO90linu4+UfzWi
U6zOrC1HHEJiVrCfPaN7OqjeQMdr92hbGxJ/vH4FU8A41nV0kE1SAOkumIQHpkmqkCpNlJUafYRM
z2Tbwkva3eu1CDDUbOvNmArKxWYa8PNeD5D83gKdRgAdW04CB+sXUS5gVqs605j5/34XBP6h+8B/
v0RjFSNpU2kWtlixWfPH0PzK5NyfUMa81GPlYea9z3ezoZ6HGmekapCYXHAtqrm8CMOvddi7PCzC
tWHtZnORkEF/ULxZ/69ARaeVLNf2WBvlyezYCacreM0sM4Btl/jWq1prwKktYOo506tmmRcfBX8I
OySF30Y8aFsHQWPMD36tmxSoHH1COG3+dyd3uARW3aDQIr5uMLcABi37atF1A5sZNF712bgPnCiY
Y+lzt2UIFX/cc/pklDDJC+LtM6yTBa7DAsuFb4oxYB8tcwfI5ffC0SWyJ09XqFAKCVdSPH1yDjTy
9Jk0Pfkbyilk6q+Ga4GrxrpriTO0R3VriASJBz1k1myPr9bXRdMjWk/djox2m8rdmom5+bOvdyoO
Z/yaCWpDapRYFamkhEBeVSP1e9/HSAGN40MlcMsJmsbSb7slzA57p2uuQiDx+1lS/gPCMnc99DM1
1CWt1COMhkMxeZGCGBn3Yy7taXZEGO82Fv4t1OPUqwM6lt1Jvgg4lq8K4loCpAwedh0WCy6R8uC+
h4bFin9u+rYTlzd99LRh9/zuVAws+CDykKvQ4vCv/fzCeKMoJyWy16s33+WIyHwx1EeXlU7q3vYV
16CE0+b795sUiVkO+YSsqJ9hd/VeuD+E5vzgEng9EKsiExi9daJGalSHxvM4ZaJzsfU/CwssgbDZ
BR52AfUiHGxyDaKZ1Fm7N1bR7DsD07B/rjv0SD2B+Tfpc0M2Qb+JgTpI6xKKzCcd23L8huhLiEVn
GY/e9Hs22oKiUdygdonOOTlf9aS+l/JVUttxrSruPUax+x5PeWIEqXJ5/A8AYATcyjhEg8IQAIIU
SXXaQ+H5rES8FJ48vJWO1y1WTbAyTUA2wL4yy97bzUkHnvAZ+P1ff1ETWNjh57kaz/ZI3YXbGzO/
rQDrzcmiD7xirveG9oEM1QiwiOiffg9lD1aeorluftrAHEpKWReCm+YCdI8eWGcD4j2X8ZVSQxMr
LHB4HX5h072FVoBjaLyjQb81c5YMIV/lilDldaD9ZXrOipCDDesQl/wlzUo1Nrd+tbCIc+931GY/
myuM8ns//fUaHgsQ8uX/0sy3caiS7HqGTgz936cCBUFv/1/H8DkqczhZy0i4Gd/6+/sCw2Wn/sx5
cVPEHLRdTgTKuTcaDROgJ66H5gSUAUKof9DmsSdVaVIaqIrWuGynFZZGMUhHyDokrhKyHeDGC4/R
VkBMJyfVspzv5K2aoWMDiHYnyHJJYpHc3lsYpIVjqq6RLwoMu5DigF+xEajawo8VhWLNEGM10urM
KlPMJ+s/g52cxJPunzJJolB7l2Pe0w9utXD2wbubtILQ8IWNoKlV/Xxe9zefPMEI9WU6HvBMrfrJ
Y5dGxXuIl3aVywZG1/EX9GHdA1lrlwAuyJx+xyBGKrEhDEF3fWuvhsNsv7Ki2vEkO39sJfLctElN
znh70ctBvOCS4vBM2GLCUzjSDORNzvbvCKn0dlvz9bOZvNrBVnk51dxYoCDE5dxdrI25N2Tb2dbt
XDwjs7BwyEC9eit6fse+vL8i17hy+2wkk23B7IXpp3jAr8J9Tlmab+GAu7I3wOX5FPQZRrFI5RsU
OWLMHigujH9Sp+UnpotGCXCfAqm1yR1/ghAJoYEF8RMvBKsU6NTaAbwt9hVRt5YAm+e12q1gKhSi
BFA/17j5J/PvUZUZrWZIlg7v92KYgzIOkR9cZP6yf7vqrgjjqPW1al/tyuwwIvefQJAvdjONBBaN
tSY1uqgxuKdickTgtdUTNGzPEtGYtJnOvyuxIMJ+YZ6qyp/Yxy4a0kJQzKY3V1Y9aC7oruIaw+Md
+cdms8q7wDJXyt1B++W3Cq14Af4vbATj+K6UvdG4r+LQnx0nOpFwf5KcFBVft0vClKGOJWI6KjLP
hbkzRg80tiArble1437bbnE0ixIEe7qwDhYwjZPYOc3QNIK7qB3HRUY/idcL3nzyt2BIDDbgdtQ9
MhfC1JPsslBHs4Vs7f9AiLAz1NEiqZVgxaTQ2RbaAQ1g1Q/gGry6tndr+J5HxVZmVGomKsoazEBB
wWTFcDWXByyKf1ghKqFS/SytfJyP3QsYhmI2zeXe5bCbacjbsB3uQ12EKc76dJWxWmeyoX1MfW3j
torJyX5IzTwXZD57gpfMIRcS4LrdFj1C4Q53adk5QFEJqJEKqMrxLkSlfA+JGfHE+BezayzbgmYd
BB4Y5csUAtQYB636rKPCsN4k7phbalYRqDfDGhLPBqM9gd6X2kIaT7xhhUdfiWsTBeiahd/dSvNK
KyvhOc8dz4Dv3/+l1b7NcZea+eIcKbWxoWW53Pfl+XLx86qBFrP3G7zrWiJiEGVRBCt/5MifBCNh
Cj4CCoqpPOuGW0vbok9NqVe/zp02uTtmBT7FJ9O62ciJhXZSjWL3zpd+P9bVV7arvn6+HalWP/+T
M0DZvrnqKkvRKdeh2Uc//0t+MAHkpLiV3/zeEip1XLS/ts/PIn0OakQOOkZ1UI1n5IG6IjxgiFuQ
IKSrojZLQcRQItE0mAKkqUS26zjTCqx0SKdykzhpvYb1kwvw4ncDKJoWRvRjPV8Rh9sdYixZEMhg
mONylaU53V6xSa1AabEqFSVaP0gqzgWbDOTgKkKjGaPoKhWO4WIokkcXnJuIe4rGpYya0flzUTlr
cUkzj5Z0BwHkhjmaQGuXWjPWZOUSv851wB3KIR429Z9IR4z7z33rIyx8CswbJS3TFJ+0NytHC4dI
Q4IyLTrMTQdqxZNfdurPQe6OZf1AkwkbleUd6OvG/jNpbdH003F4HhyuenjpqHpmrnrTdoMyrBFx
8OnpGInNivEUKVZi+BIYeWuntEdTgRgiDF3J/j6rXqOKXCl+4KilOSGQmsaUSR1hkCNU/flRU/Dr
kgbXen1QLlKhSEb9v6GUyLncVV4yaeLN8kJoTwSjH7zkhpR3TSkpqYITQY7SFtiVZggPzEpjCfxN
ebs9L3T1ZGIe7fqN2VBPbAfzxF4NO2RPy67kuCAyTALWmhaZmU2e2IzYr4811L0dO6r/ZoqzNwF5
IvcY/e+DLwrv3VW3hSCAxPI9sO4Q4e9cWN0jjzrCb8bRvJIHiBqGEb1NJHmPvs/grygjHso06B8O
uiF1/hw171gtn/pwnJr3waqv3+gJ1WXJnUcNo6K/coQaIL+mnpBcRosaGzQvY2bxbvNmG1HkJF1w
vpIaGMzyFIPQCowRQnWbYuBmMcXWUb2EsCgAoNOUIx56L2NEtdY7ObdcHkqdZ1kZXktKSCOkjMLR
KpLLoXrPHM1ydIjw1gv7BXITB6gurOWCp8lI6cCucP4I7xKDBdFqbsmf4sQ+t0kQ2J50PlbTm2gZ
D+wrvx+VJYIsil6/x8Rv7ljgQpeDtEA4TQTPy6fQCgIw4zPxM/xue3nRDX+ef0X76ONB362uky2P
2KA5BD+MzpUX5oYUWYfPo81Q79ZzHHs25s9OY4q4Z1dgzyxfjoTiLHnX8ZfgoAtu/MAHzMRtM0tn
S5C/e2YtUGZwECrhuYqalc9qOgTWCn7uRkEsDADFY8b/wunSq+rFTfcWLezFP9CaDPKLE0Gwgm3Y
/CpgMxSi5nITKiP/A7ttxFOP941xRUgpCH83wQENifIFchGFnEESMunYQ0a8r+bKcydpw2bN1gNJ
EYnjY1BtzauU4PTH8sD8xZ0DWdj/K+Qnd+mspkrBnMjMxGc3oEIEnkz4LRLOIJGPtwAB8OGUqgnx
4NcJtnu002DPZRqsRnMpJHgiw8SSNkHscvcg+likS43+66f5idS8xmkhjbRkow720tteO5/dEx67
mv2bdyGTgH3UytrrXmDOlpj6Zqui0EiRgU+hcvKdCd800EWpHbmt4AWeT6pNkY+5UykpaR2nrq5R
vF0er7WAiTjlfjWptx1+zOyQF+ysuOKQxLmRr4HpF5xsu30ILDo5aTekL3rFpGrPQismSgWZYyOq
7UDEqKScdMgE3qpvkBjYx/wRqJpxvsX6u/386iVi218l3okqENF5zrlXk2gHaY05O2akSf9RA5rz
L5HrKMFmSXdXyubd0i4/FCgU1NMzgv8Yja8FVJfhT+S3fdstm6+LSKKnTs114q2aLtD6l8qmQGGO
03layvjq8OhTo9o4IT7oXhY7kEtidHuxmo3L7eiZL40Kekunrl1yJ15qoxLecxYSyw88QfW96FBs
/fnQomc62WZ8D1b+iYwGnA5d1QfADqUyJcQ/L4sKGtq0PD2ChZy1Kn/cLIwj3GBD1x7cmJzTiRPU
AVxYCNr4U7xg32kw43WWRPPzZpKsilJtXms8wZ4/5V8erEzatZMWcTCRElNwrtL3MlS40TxBFWp5
4vNZUTxdV96qrMHca0gXSmMveEHs/HTeOd3cTYsaO/4UCW/gUoPBUq8CPUsTb+uT79/+axsCMuwC
WlQYUGbIKzX3V99AyblLHWImhHjuO9ItSNbqXThVR3VI52ALTQjtlqEhWLVdu7XmDnm6aJJY8Ke4
AjB1B+7sf/ElBStuz1tWS27BZ2fOgfeDB2rQbPBU/kDpv8FSdCZNsaVFJCqocfc0ENXtaWBlmksu
eCLggB9s8Y/pri6zm9jUCSHvxeho+h/dwSZKWTIfarBaAgmmeQ7MtmvY77mE6qFpkUlk9N55EAYH
RTAdWgueNteLBeUDnkZkwLXtDGs7FECIdbRt5ZzPMxRMZkF1ajbbqhdBZ2CKfRSrR4BAcLF4BRGA
K6UcDPAjSM6Cb2eRjWUccf5VmVa/QTAd7R1facny4yGgOTpYpRPCqm4IK50lnUtkJReawd+2ozWG
1cH2jb79TRhiRCRTdyeYj4Eo0EXwPp/pgpgrd3y5ULilwEes9PBQpq9omlzPdbd4qq2NQOWselCg
osjQjuhTPes44s/enCtySUj3xlJYNk5zRDeQyJ387SneWF8LrXfIXkYSy3WiK4Tc6yrqrelKxcvu
PQ7YigAKOrjBKUxSzSliazVf8cOOiEf5i8yR94EEZ7fa+vbTE/MjANL3A8aMM1smJSeuiyFIAO+U
Mvh0NkPkSvEQZQ/KVkzXPb8WqxKdONlH9Hqu18ZFY8shaFfh2He6zzLNpnb0SLAgjJtxWnVYCZ7z
Dfs/4FTJnG/HOt6e1VNkwASDoEqcn42pZmIXjXRhaZt9wwT0kJXd8ul50rpoWOfUNF9Vf3J5IBUV
R3AxlMd1a7LFVqHIZs7L0qudq8SS33EKmh4N4r1ryDY/XPNjMWOUzw6gAm14bEktpEYLrHGCjfhC
ukY0UE2k5YmB56hSkB/N8ygcBSEnn2QqFnA0uDKT3xPqCbQCEdimKx/wu4TNtp5yMhSlMBz3irJv
2CF+uTeqwcdo0rNDxL+x0L0WSm/e6FRwTP83L8w5WmztsxLbYryFVcQNGF6iIqTmXG4Q6fNkuqlS
Ouk/c/pxaW0Z54iyH8qpmcJKs48ukQ1r25Qq43qdyj31ndvmR7IJOfYNOL8TZnekOeVHJvLZ97mu
nc535XP0LSjDAsYH7ql25LxvGeT+VtJ8/8qedRiRDbkJC4DKxbdE4jjasAMtUzUxGJ3G8BtJgE+k
ctPbTuEVFqrvz+Y0I+qsatgrZSGXLIdZ0WAFJetwhLF+ELSDpIrAhNuI57FECq3f0pzWDRaiRJrE
zbMeLRf72Jr81pE7Pi7rG8ngugjWzzSFftKjK5wEZFJf78x0zMMzEKUfV+8XXXfyPBu3bW3FGoul
Cs9WDRJPaIgA/CP0tFhrTAMqp191/xLpN18pPHAVuy58NT8WMlYxFKwNWt0vP3/IIx0+Oth4aKWO
/ID2SnPl9vDpqer5odxr/pjfEFM9Lg367feBxPD6XHOr4RpRjTBfsH+dZKISICRcGxYUQL/QVeNL
OdENd5FZuvMlhDLQ7gJt+GwOoUYuxl6sELVNHSCixQ2NGjtXgjg8/S3apIcwnutkZnAuvY5TFXsd
44slZZkhBvpPTGpJCkoiOnVL5mM/Ga4zy5ikHEh75+64YyCsx/BB5PzmYyaFZaWR8DWtUFYTCOUw
sZUpDhcyRSXyqCvuuDN4lMHM+pYNYTVs5MTwyyHoVbAzje8L7P2ZZ7eCdlB4DywEDyrGbvhYjVkO
Qyr48mQ7X6H7ZGvZuWkzu09i7Y16qLXDoVyYFSyUocMJYnaYtAx7GVbraBmdHQwAbXTz96JhPuNK
80cK2K7wcICLbn44R8JfB+K6chEugmE0aEA3PM8Q2Wu6l1vhVytk6k+NZYJTcecdsDayfqUD9puC
9AXPwvunVDsZvEEojOn++MkfRIC/90GRoHHVFOefUWCv7pZIlghCoLZgvDyHNUT6KNQ3UXfTd/OM
ZGE9cDxYpfGKWy+v6vQEyHzROx5aQt5EBlD5swYIHZuPpww8n3IF3dBQ/0MoLBToIvOJs3bo3wLm
XwcY3rzlZfUGM5fKHWA46e5aiRkWYYNNaWkrbmPj7aC0jITkfFanODImPVqf9o2xz2n3mrhpV4v2
hYNT6s4yNMkMQKMIYbWU5HaJKdu9wVhQZHzPCC97RCEIrKoJiAAcRBfykotFzZsR8ZOXNoVanLhs
r7VQyzCuoobgGzdFobAUqa0pkC2bb87IFoVSsZHO7sIT3B0eqhsPr5vYzxf8LQyAJYy37w0lZhI+
+g2gxg5jT7/TOy6qapCEUYM9oUv2IHEpnTeSIk+6Vr2eBwNrGUQmW/2KUfyuLTGoExIO3ekH1qpt
zq0Khk9DplkYgvY+g1o7V5zfXwX9rrmG93/7d+xXi4FO9591AAMmOlGTGVZDJy466+ExwOiU77cb
vGKfNqZXeIO1dUW6ZGCK2kGChSLpHkwlCQ1mWJ3OOwUQGaycV2gABFYkfhLc5P9W9HpHh2kHoe0M
SD46g9chqn8FgTmRd0P4isgb23KCZVPtf5juiUL0oMd9eUAwVnPTqOavG6tG9jq6DZr8MzGgorOS
rawZLe4WbUagyouGKR2BZGmF4yt6y4W+vVBQcHrSbqMfHdNNgPqBkArbW8C4qvXbNAuvAoAlx8cU
/DjBvz47+3DE+iF452vvC9lbw1ENdkTovzaDVHQZjjBSy/rrpDs9wRxYUU8xgu1HUEqUMh7zLcAK
kDCFarrMoCCjqUcDWbW+PeQ3WUXlOBtKbb12SZaaSQQfb/VHBGptxSCMqBaRSc1xS0Fy2yYL4mls
fLChD69bnUJIj7tY41AW4Ko8eqU/w4sx2YzR+UWrYpRVbPc2mvIpeQDvoU2IWA9UraRoX7MmVIXk
Am7Mv07JcPCInC2A+XObX4TXLul/idmOTW7bHEaqpmTrpeSLGuR15DPZ04wD47NA7akiAO/37kVj
vAyci2tsrd9RI7PZ3KKvk9SlGzAFhsD+CCkmiHYhBmwI9gWQT6adcYQQ/v9CV18MFj5F2i2hVBEH
CQMPLlEvh2rCWpJDPrWVbcrWvDNhJwEE+tGTmEkL3GUcsv3qM1k6lz/ADTHFv1qEPfDqx3RkUBYD
c0f7qszwd0U1X1J7+Faa3wAtAYAO9rXiTs91B4b1SvrW/TpsOLkmBd8MP5R2Od7W+zP9/GR6fEQH
4jxVjn3DnZ3zz1Obi8ztUEvhycL5ZVlyIZw74L6u7OUtR8MhYHtKyM0zSDKtxv70RqLnuE0qX5Y2
OshH0Zi2G9px+oZ2Fkdatn6LBQ5O3jZ1aL2cbvv21ebyxgQj3aoM7m2YwEQEA5eL8dS+UqcmG+5a
7EsCGVDE/F3JbhPraBARLQPHtEFZuCDVZLZBi8eZ/JN+NPiSk8ETU3kao9I1V2C24/kr9uQKgbj9
dAtzVIIJ29MFzDpEY9B5gE/dbD5npYDIZrTzBhAtmyQX3FcUUG3le+Q02uyJrsGhWV6kj9D0HBcc
4RHA3WTJYvGi0Np9G1X8tDKSPuGLwz8F7tHdASF7RJUgiuViyK33zBj0cbcw8tRKeJ06AByd+7EM
4wNrDKb1dpWEaC17Ee2+UENND4+8ZlhLBd1x9//Y9fOq3tU5BMrMEKuVyjiMTxBxUsXgszAgHANx
AOHrPoI+QPr9P9586JbBG1RbGewbQA96inabGjhBvUFfEVlSc2nYghpvVZ2ycZJGjQhAvEvamldh
FWT2I/TEjDsT3je9q4vhD3lpxjUskKNqJQ9RPZQLyOGMIgyKdcCgOcwwoeggTNerWWZKfwoc7a6O
GoZ8JGmsLCJTvYJB+PG47whM9XCigdNKmNBBzE4NxH/UxZNAdDZsKW/94J5YEI6bFY4ZMARi8tE2
rFEUEimDUXstctJc9EekgfrhoV7YBd93gmZJOY7lYtYADR+jz933N4Ux/dGZ+n/ulJM0tNPX5Gq8
Qhwd9KxueX5BQOxY+an0ScoCkx4ADUQ80lekw4xGND4/srf5UDcbdVQZ+NwQbfB9/hA0HMrOiV5K
m5JLAHpV4djRmJMBjfqNzJxBoo92xA62f517xNdgwmM6oYXzv/+MVJmnoYQV2zbgpLvyuWAbEuDK
XUWMgJLtFqDpF+easbKk6tvudcjDzx7qlzkFFTLb8D8RHnPc3eu2jp6MUABzMolwtHOilF+Bnnxq
iKIQoEfymlTkYHt4qqKaQerp08+BYy64ZsAj8Qyj3xM7rRpa6QHywt0U8oxyBf5iFjdEvWkfNsDt
E7MU4UEopswbnEWuZYwSSu63oQkpzp/DbsYpf1ZnM+Pyou76yMYZzxcanQZdmcMrSsqV7RTWNgqt
y47DNQSpqCrftToEzucV70yaKe9Ao1rIcM8LjJVkcJHwRpii/727TGpMAOVeIa+37eE4NczDSSc9
NAR4TUuvfk/UFr4KZE0Zsy+2rpRfIeAuGR9Q8BDrRU5vUt54BVsy+r+lXI5WySpAsaUAgLb/G+Qb
3lBd8HL+aOPoqV9ZyT/hSNndba/vhu9WGc0guYds/Jq/JbIyoKm05J2DJq9RJPvKfBGDcdrvqCiH
36VPTwqgvSKjYAKHfsuUHLS096T3LsMGLd8aPol0FxEQCLa3C9AE8DtVLoSljSFGYkZQkb0GHjeP
fRoWVpXczJ+virrVRjo+B5QdlzqzoEOL1uSBUwLrgoxs144lWDzrFalMOsKqLiKqCt9S7Y6GAHS9
V260LFVm2CEmMNRW9LDrDC6hFNfQoDyhVPVSmUNQrDigcXhZPrRljUwy/6PgXOaRE3kuFSMb3JPn
eeM3k0l0PvP/inOCddJ419ECnElNyJwJGA5QuSPi38h0owGNFW7eii3yBwoda1X4elcWdDKv5wH+
nXedh/aBPQ5AowICd0rjHVN32/UFmtlkRdDA/q+ZFOil9SL5WWm20Qts7XPEJzzRUD9qKZAN3NKM
Xme2hwx7H1NTvNd1qXnHM/Lq6qxO0nVQktqX68Nhlo2XNWduM4Jma4eJMRlCAbCqL6qOMyAq+bsN
CIDXjSr9GQ3ISlrvVFm8uUEips4uiAWXGhqiJh3OFO6PEozWLeRZOXxKM2HIl3mBuGSLTxEOb0ph
LXRa3G8JF57QiQHaoeawcDrxuyK2tDAfN6V3Idw3Rde2RyKqj8QXd0O/P8Wo3580qxjlBhknUCQ8
eDI9WvNPujSliFrN5GaNPA5D7zQx1HMimyl75ZYj/qT6MrDW+LwEp/T0DLg+FKJCJ5aDPu1XOPKi
BbbJHF6YV3TohUUioTnX2BKxUhfzJivIqBTl/iw2kviojMIt+c18xGWyuVtWq+l9YRNiuFvXebP7
naO1SOddyriMDhDBSA5+Ukn2rH+0tdmoLJy3ipeDWUi2N4wWCN4W9LeOpN+w16LmoG/gXT2m5G2w
s+1H5Rfj4M0Obi2FvoyNeFMD8tFNr17ljJpN6F5St5j9kkhBGHMNhot9LCCYBtGRXgzbMDof5CQM
cKsTa83lOwxf3KAQZbt+3jAkc14qqIko4xlJXgNOyTQJcpsvdo7Qkn/mKx0oryfoH89oTYPU27Dd
sG508MmS/08mrPeXT93NbyjDCWOmHcfGzWx3RJYhxTkopVPYXHXBFahp90J+Z44QoTV9bN+1IFIR
NNy+9lc4VAozvA010/Qgs0nG0AQKGJGk+H4hEEITGors1fpDw/wHYCpwKhIngplxW3fteuWZP9EY
Z8df7OawYLboXVE7oKm+x4LEX4TyvFlkY2w59linz+8O58NWzLgwNziLqHJ4mXSa+SwWbp0NyVxG
3XNVSXp5WKFNy0yt3ChC53CIuZksuWt4PiRdjdPz1ZwCWoeb8RiXwdFDGmEVGwaQ8SwbT/Tu4OZz
7SXvjCR7eP91DvnTi+K1AqvFJeOiEZHgGR5silMwl5u4vb7AOtgjyKPniQm0LIj5oNoS6j0246Fi
dfsNWQiTgvRKtwS5SkiPMrz4rxqwPhnzQXQa7d3JKQzVmvqZahAVeHyxWRtJkMlbPdKO2S9eENAT
OObR72ySN9gEWZiKmKnng916DEnjW93u6R1q7ureF1wi7i7jrueb6T3MJ+GinVmmzIouTPLKtc9v
st7fC2kUFkM+A17Ku3DNt8qDlVnTaxDvAy1GMXnBCGOJJaLmNr7h7/8jZmNbjWT4HIaZ9K1KsBzY
o7DYYMSFEOpdspqjkE696MwtnZdrS331mjvZojcXBGmTJh8ZUhdsYFP+OQ+TSFDhY19gUmyZtwtM
3wTSpTVm1PAt06Cts7b82T3+IEPyQTbVWkrNt8KpYe2zCn08DCB625ApMc0U2RLJzuuC+Q6ca30Q
4iVGN3TZ0h2/BG69YCObk14unPVlAoYPHM17ccyEB41pQc9r3exGICjgwsYcKkW9ps7ZqBp3+Uww
4446L5/Wbzj3ee+Tfq/Blojxe2lPdHcjgezg6AdbObNLcBGYkqa1Q2zg+UWbrGFAgOVfaa01HW5z
YSJcjgPEosHIVTs2CBGg7POKs9Nt8GzrH9P1kMKUiYvwGe8z/3J9nZKCepQXxK7yrJ6zztIrjlAN
FeUcNdFsMPIRqr/ATWtuzHnKSfA5Pi6GhUOqVTXSxva+u+MCqu0/QlHEXhWSVFmPO5/OooqyXRNL
bLRSAWxEbJe6kk2veP+eCvQfrk31jUUH/9OD+1CWWPBezsE2/W4BD2BGhHdnoLGalE0DQYJoSf/T
50bpiQ2Yv5+ax/+IRjtqdHpVLnIeY0sV6uY7Nz0GPRwRyc5icdvBPKgXX8QSws+YxwfWa90Sb45n
aRBnHULHl5MTEvmj2qVaka8IW5yazz61ByAsQPC0H6Kesgv5ZDVS8TODsXEIrlrSasXeFgjq+W4H
SMWNPUhP5zFvCjLspEMdc5usXVHY1rOWtrPfGsSptXaf9fSeuNO0/T3SRQwf4DdXDUag9zi8jvEt
bCThACFzQGjh7mRtrwEiZnVOzUFR78dl0PVQU+3kA1noeOBEn3/4cEuB0I4lHDe56p3wL2HQ8rzz
3CfONdSokod3DiDW+xeuAH3C0s5UhEheI4kf2Y9VCRvxe7svbOqAMQqJmMBPTc4d553JaN+hvokY
aAD0e9MWlQhyclUSlGqoiu/tOnkuILo3U7d13vinRv/M+szGUl3YINFTqPo6G8uIECq7s/7ONXw8
HPgifEtW0SsI0b+/jnVEF4dcBccBYWGnoZPk+G0Gw/xAmWmSkMPujXLy8XteGvk9Ds7M19ZFt1c5
0LoeS5HGK67NaljNqOaYZhdvYnrOtSOh6+XhcTtrfQnm83qq1Mn0uj3zjcLCGKVuJCX0Jh1mo241
VwGJ6TuXDrQSODKclNgjveJZwAZbhVW1RhPldVEYD7MXgMsJQWd3IKwXe8UKmflK1tUnoDB1SIQD
Dnwt8AJT6965WkJqsWfgMPKytGu1m9OtpscTXM1YKa3XdjbEz+kgSSiuLkwu6kdsY9ZU9colPEM4
lASDaVBs39lnHdpTlsrSX2XfCduQBN60rLetgjwgqA2ofkc5BjYXOL8H//Ri6PVLCjKNkBaJ/K/u
GTFwXr87kpFfD999LzlHgnUsKlL9uQFxblT7ck9ST5K7w09ol27/VMndLyHHtfqLAguyXqJ+ja8d
4RIm++dP7PX73BiL2VsHwVJZNo/fFpxWcr9EMXw0tRahsS/O5oWJx7rzYd3XkspO3LYZjxpbE9F1
n0rmSUNv1k/XQOIQ9mVaUzw/Q7a0Be9J1/8kgStItuzjKQjRVYv47wLfJem3ABzCaTKJrMg4Qnvs
9Ig3uL1ZrZwLx4ahrt9yJ+0qPxKVOuXivTiL8HM0WqHpys7gbuc9U9g9LmX2uzyeQonXMUO//62N
bzkzrsvjdj+qr3YdL5q5+xXdTCNwWaQfsiFTQN1kB+R1d+py6KcyWXsQEA0gaEeG1D14FXcK4BOM
dbduqbSgDgwZiVme8JFN8uFb6Z3vEW+iwDAeLXkoaK2YOvL2DRtFLl/7zldxM+Jmy7C2kzQhSnDV
XtfbIC1yHhfMDqe6PzHb+xe1CrlCyTrjvPou8Ql6zLQJP9hbc+UDtBSPBZmwxYyiLY4NPoe8CKSe
b6MntMpuzjDvre9YrvjfY4xww5gNg4XwM6OIr6tkvGYbJpc9eWA/fHFjX3LJEhkMg26qlkXEiEEb
7hpfoUHe7o3hu26SY/K5Ij6/2IqeUO1PSdvE39xQKV0Tp1lC5Lgtn93mu/oSonBLuT+ffYnlrE/L
paAcJy7COYtFU3kSz9NynuVXidruOnhGOX8uEw0/nH+kF0AZBoj/Q5BWHco0BtIbmaBJ6KsvFwAh
/UJii8i5yxwPY0JQ53vmdhY379ORuv5VESNnzdfxs0dO9Z+8Tc4lS+fEJ6c8Wi0BTlnmxYndt+yF
pEEmW2WlOsYJTrwd+MeIwRccwj07oHQHDxWnQYNme7SElRJw+8N2UWaj5kWcQDDE0BI36PI/t/2z
iyJKMds+SJiXuwsQcmDotwfX8o8iUK0SLSeJ1TYu8UZFuH06fWI/RgeJv99SAVOnj3Fk39aKS7CB
IKDrVhRW0RGKLjju+hOm0JoKAZgicJXWYg3MXXAis31YVJchjwP1Wm5pxdAt6kcrHOkOvQtUeonh
is1udhz7sBf4uOT7BPEKcn31iAw7Kmj920t4x4KLwVrHvk4z+NeBUXmULUFSC6iySO2c/H1I5zwn
vM+UI99080pb+BzwixLLcpH6Io70w2AhIEI7I5tQfFRHazJUzS7KlLMAX+vC1wMNaMhxvMNmrorv
j7q4QXrBH1RX4MZlkDGcgfsL2gNVmX3l2PP1L5WArgVg9PR/SMJ6ek7ARTNLBOtkWUcExmMN26uu
t/ISZfihN2hfxLOjnhiYhiXJIGdjuSydX7fUL4R8nFs+ciY0VMB1z0eCOqDgsBkpfdAHWgaIQoHQ
wvOxywbT35bKt39oeN9dCj29Z0XtRLI8LHe2TKys7xnpXf6NVbNV+lnffZsZdveBLgjlAdj13gnl
d1irwmWYZxBfOFzAo79sy+tYz+5pGXiMKnGO2ApUKaHP9YqjGELH1gu6NjwPkMVATmst32cr6vqM
Yl2UAvgDefei9yVD5p8vMrjL/zByhG01lCtE/zICuHMm3JZelC/pjntzbUKwt7Ov+E8Wyhi6I8mp
ejJOZaJbjarMqU3LAW9HqLArEWC49sp0LnqdpJK9/Hgpqnne4QxJBSDFqtlmV5b96GF3rBCIxM0v
NOzx1B0T2LpZEth/RePKXn0O1za9aRi6t07knm6fko2RdcvrKP3C2VNkohNmxf7byVfGPX1FPFpB
RZG2veAo40oFH5q/dmRRI2/6A9XCfgC1jE/BAUVdU7Q+cMmcECO+SrDyHTUyg8m1a577xmSo/Pbc
nNg4HVNxzWA4OE4i1OEBQ0quue9UOP7AWHISnNYTfF6SE4OCMLoJOkERJ6lJ0vtbgkj9McZyN3Tt
FuLT9N8YeXE3FWAuWaNEUhLr/EHlNsqK1OvvBTnxe427qbUtUBtyqqFgcyOf8mQcaCBcvS4XR4dP
BhMP9UA1a44tSJdpS61cL8Mfc6zk7Pd8C1j6/y1Sy5JGDeBmKd95L4ZDRLWVRv+E65DpPzWfARU6
w1HdpILVC5cgzBaMtNfonifgajkssop4y6hba9fSUg7hsLmFAfVIO0LXJOEPI4kXyQiH+Q7Kg3I+
ZZkfgGI2b59kuEcsG0dHxNhSvfmtUvJZsUFJ7uTIdtS8YyRkc01axblOupzCNHum3oM6GOXilaXk
it4r8JNstbXonYWX/QDFPkaTdZlldf24C0L/YnYxCagG4QesC4CYdsF0p3WniHXxUnLaNSUOQFND
04g8HM+TExcmPcFt+CNmHQi94mhP76tY9xfZJ3eZaMZjoZCqFtr43gsyCzvRJ/fYM14gP/VtF7Bl
aIAPYrTZRonfKt9tdB2jZD2c6LUj//WcvL88samhF66WYFipXkkoygIycucw5h1JwziNZS+F7iaj
UYH4XRR6hhcJ5/qqC8AiwvMRbWlUl0BD9+jIeqoOw9Lk0oYHGcvKvTKtzl4BLVEFwjkWlBxP5MoT
/K1JbviEN/rtEreGomfWA5d4VR+bqdd8KqFxCVz7LUgCQRg06Zb5SaxiLkl1Xnm6dQCRVCbf0WL7
52WLh4tnLY3toETtJu1tDfRDTHRAqt4bJnXQV88WtfXE2T7TsDa7vSfl5MvxHr7/7yhsmn2m+NrF
Oi91tPdd/ZNeMxfaow4474WPM3g8udz6A/BhfNEVqoBb+OK78D0DyVtt/gln79spmxIBMOR2+eJD
k76ijhEeoyE6bpPCRicXtIYlDyusQ/SaOZyq3MXN2X+6qZ37PlfQO/NtmjAXMGEdRxC0o6BWOHeb
/EctbNfFc9yqDVneMIKqJpzhNAhfQhtCyy8D5lH6kb0uf2REPz0W8Qmi6AooaexIwQSTxTKUJRge
IvZhR+xnoWnGNM8nGkdjxoH9KeIZfopdaVCrokH1g+Ou7EEh+AF6dFhRjOWw8eBcQqdoN9XHprHp
V0jHudgavUo4beY97Oj5t92t4squweqUKwj9YBgEJuAk9azMcnBrkAsGYrRouHmiEr3bfteI/Rg3
Yhn3jQ7gczyPhdp5pb76mq/7j7eagShlDLHE7nSZQKClp+h7x9JWrcalqYayFaDpMMaRjBZECLpE
4IHa0D+Y/lC8iVDfmBr4/27W4VecpbHGFBkZVaYCvxe7gpgGCruwr7LjUM+oczxRmv9f3jSVWJfq
1tHA6ugZCyNOFLdvcyFI9cdC0fm2OTiseBH9jnsXKW7ZgrdaSP3ShME1ICfIb9looQWt+0OsReFx
vO0KmueNhshKHgdtslp7uBUe9mac4s7xuEY9ctL3NsEmKqBbSNbQoucWUxUyCl6ZlZz0c+TOL/B9
VQY6iV4tiOqRhuepVozmG4AP/EmDzryyaOXl+oAVTC4NgfI99rzKlpDkUj2ppAMUXknPrThRwem1
A+ce5Ytuz2lPhrKjtsEi/mesIJ4BZ1MGrxeDNRSVjbeDoTjwEo6kDrDE7jFdSGox1OQogdqz+YW0
f5GSxI6QAnhTY9oLG6AYhDibiKSE1LJqfpPOH6WzUeVIBD8B2cQASRGwm8EVPpw50Ml5Qzp7Lf+M
DmGSOTZPbFzNoeRFSSS11rQ7TtL8nCcCDsL1BJGv0JitTV/riokmNSx82NCaJXVEs0Dw8ODiCHt+
5/6iOj7QvSleUwEN8J75JqZ2bwnTRVRz07Ps9fgLfa8RXRHyTia5FwBQstm7x939qTp3OkTBPjB4
L5jQ+rTjYlrnLbBGL3hnjZmyUBDf3keTd1g0JJoA1rikO8X0FuIGbeMryd4NCFVVdOxpgIiEexlH
lRSS5iLb7p4sqXnb2zZTLKifCbp9oXV29LGKbpAlPg5+EGMEE/fm3hMWDhEtGcvDJ3v50xaX/KPr
Pyf67uazW0Sel5tXMl4Ahe7ZTaqdn2ThYR/YaK6sr6c65e09BCCVSbcaEqIrtNoDybn5ASFf8qSw
JbSsRXhw/hdgY5mpaFn4xbMlST0x/vo/yNzSHouNcJ+MwCzWHy1oZ7/hOQ454gCIifEhu7U+iOdV
4OgossZ0E9HLtsb/tFBElbq6l0EKxuzSYgMLBWGJ4z8Cdn4sM5OpvuHTlgZxq2WDZgTchZ+NJhyJ
fEjdwAAMxt/goHA18KRLyKraBqengzL3t5b6vamMrGaRyQziyC+Fc5KhV4bJieKcJH4+lEY1ne+A
KeXBxU9bY2c/hla6hifHdcYwuf9YHp9c5wIN/5DiYWmJXIwwyiXEJuZETXQ6hDLfDX/yVBFh8cLo
zClqw3OeTJBs7f7WLnmE15qSONSaYmAc52toer8wqovl9+yz+V4iqIJXsrNprnWpy6WXIAjpGess
dqRC3jkeoQb5vW8RjWn3wIVjuFnaoT+t54ZJ/K93oDmRSfmmazuLXMPALQC+wCcleF2LCr7sc+sr
jxYr0c6JRG8uACykOVaJ0CcenC313NtT5VGGE2HC2C7CJUZQ+6dk/A4N9IbXDSP7Z6nRVcx5cAI8
3X4DiFwRRQlL+jQBL9T4HojwlyWZmgZkLrslwm0gqNgeYBAXAeHpKlLGQmT4RPEmUGJ5tMEyUiHO
0fRhBz2mPbtWwub2wEU7UcM0ktb7CIG7jY0PZClxO13P29mb93NzDe1tb5sBbrjjjg926kS3VlSE
Lnfy374nfh2/vR6MWOv+KZOC/OQ7Mq7HB3/kuUFqTbU4x+l+rRjWnCJSlOo3d0YrRKMJAWUnM7X5
O4SP+7GmGT95Pv2Y9aZ5AFNqEHf24syxgVIdyJPgMO+eUDy/o3rDlPascfWxx9YOfYtnDX0fTbhi
fjA1zW8dNSMZNCqK+N2ICECsuTHRR28rkkKqYE956SBBSfQY8kc0rEk6RxF6nF/+dm5+XH8rcEJg
Sa8h7oIOWC+KGdk4uhm8xhaoqsmY3wuWtSonP9a5ON6tfuMWq6JkH6ny6YX0ojwRSeYljiUqwkQi
p56hz6wUg9y86rySR0iziqjcU/9Irpd22v0WS0oE/1kX5h6tCOdbTXT5e1hrsHybO0+cGIDTdnKC
Nuk7sy6B9rVxXHigWykmuqrGt2/11y0w0bxFEkC5mhLdUKjG46Z+plb4d5kQIFon4T5bud7d3hzu
mZuSYyLwERJnhgNkEwnUSLqcWOuSEeGyOQDIf9HuTOkwiD6t4HvahSRZwuCoq39iPtYw9LKdEtmF
XhAc84zaSTGY3omFBBq6OhkrkUSClEGMHiNqP9uEx2BjjKtH4nOth7MwGF1PGweDspeBPtecq4VD
PCSUEXvwslSGUCiZLG1CzvQkFc2pRdP3V4+L4X8V1G48Ze2uY7AlEnGftuOXy6le7v/bqIh8hXqD
ybrFoBYGQM+WRcA8FouguywldcT5WzCBFlPBNN7IGYsLM6jNqRNVRqeVnTwSI+rnfmrZxNNdkntd
IjZ4VvOC3uyxxtLkTf8Pwx23Z8HV2I9Ysg5PusTarK1GO8jlL8mvzL0fDb53c5ufTyA9YchiCe72
q41HxnM48KDhJwv0jUrWiUFeAxgCXDC3akRqDE+xO/SZPUU3jjsgaz92uQk+KaiIMkURy6bsPucs
VQ8PgXfP2h0+rmZpO4bUdW5xGUl5yr6GjxeEBpWl2H1HGzRo59ZmCxQ742bOdo2O/UWEsdwzsbxC
hQFnE+ovjCXbCA4GBlvHZhp1xi+oBoqeYRBxW4hFdbjrPCwZ0vYicKzKsZ/OBtYFEgmglSAHWX47
oBT3pgnwW72lqGtWgphiUOzTwrot2ecOXIfk7CRqyXGrOYYgym36gnvyHNpVPzK3ZpPlay2QEYED
hUMfQiJb9AiUrriuQVSsLYqmTuCgZPLllvN5FsBj6vSWzsCOprYSVf30R8gK7cvExD0xfWx/IJ7E
bcXYbvEkgdOImfUKBzfg1nJw/2o2KrCh/71sdqSuaQ6IaFm3+cTk4EgswwR7HXYN2vbAmHPPjVei
WN+/f9k3bkG57vLkg6BXNnzW2WPWptpi7lpC2/O4j1bs3G1fXs20wSelZwvHIF62qPpifKl4uTlR
Gzcpc1ZAb58Na/YPFrz6z/fSTENSUoNMHnGMkQhDc91MVCj3sV/jDJNbsC6vjvTjCwE8s0owYWa5
xcTt+2lMiDVb1sFQA3YsmBORfJk4r0RXpqY8fMaPlwRHP7hUh2j0IAr9jdGu/5jtNlJt2n4G6i7x
0fMMa1WCKiIZtxBW7PfZXTrxQHCTLpsFonmgkt1FH/VpJFXMWFnwT9PWElAhKpUGnXzAfLi9Ue01
sF329qsumu4I4HwKXh3UG15sK/wvWEu081pcrHhJ26PesrnPMpGPmWJflpIfLM1XqIBi6BnNvdZB
IhiWsw4bVp4MRdSJs8FIlEt5wPIsodXy0aErJW5FA1eweZE43/RcwldEm3c50rkF0ABj3ZDo4KjO
+if5H68Dn0/VywZQ28R4PLTNZx/NEu+2Scht0xlKnS7NlV/0ec601CiMkgUwX2/8xXweyq01DHpj
6L4msVxx6/LUCLnbtajwR8bV7GmFk/oce0e9cDhllV7yvO6HziYUaxovG9/VyTkRLhm2v1oio8nc
JNfR1kC3BkvtVmhXdAdvxIxpKSF+3vwFskfkM7F/2OvcjrR0lvwbLs025s29TqsnYcBzY7McHW7c
FNktbIME1fZNl1R2GQbwVkDllatCm6mhASRP+o4nww6LVkv87RyUTfN6TdEaaZYui+3h/lYhWr91
Oi6DEZ6TvVuNaVopXvKCdb/xZiMVGJ9fgNIFOP6EdUqw5WlWQovuLP7j75YJtOzRgJKATh+mUBvQ
tstDB7Se//TxYLyzXjPfKXjlJXGlJy7SHTEGWxo0Xy1GRMexnoL+e2DbHQAKoelHqcVRvmn9UOWu
5w6nroSqWvIMC2zBwJaBu4ehuKmJi0Z1TLx80KZQRuul8nhu0+jJtmjzhBnHzAtlujacTUtgj7er
D4QJND3s5KXf4S7dnk+9YMjVGElqQEh2zFtJOB0RC0W6mExLMvStFeIvlva5kINXafhf8YYJKVG/
lW6Kgzm/LpESamLmgXHw89wwaZ8MastjU8Osqy8QrEPPhJGOKkkbTI0UNwLCKZ1+s+QDPvPyCEDu
KMC4QA791w9lwH/8uQS6nNpW0sv3gOmZvhoFbnzF3Ymm3RcPS7n5p4/jpT57VB7unueXhcIm4Cg2
K4gl/YoBPDK458hfEI3CHfFPgLmJHtGzOX0ujPrqFWAKOKMCtuFX1iLMvbpg9B6HjnIj2D5p+yPp
o9uVXoanYtHySsoUnslW1Sm2qQFnG/ULPhs4L+vCZIfgAXSkT9nIG6dWRv+ynccIqXTgsmMD6SLu
eW4h8yfI6w+KiQxSEiiz1AsZ1fbeR+Ofdx19lQITFloae3Tva5PWQ4LmpMbfeD4JBzOgannUu4Xm
6qfdnEv0L+D3PItY1TpyG1G1whyiDB5V+BgqhpIk20yL8QaydEAL85gvCplP0veyw+dJbxWjzJy+
SdEOV65DJQasiQT4EHfhrjSPLj3TgSVtrRHup78/AB6JVF8Pj2hUi/JloFso8hZnVvLDml1pbqf5
0PsRzuKihleU5Dk01kr7cIvvJ/DkbsjfSfOioV9uuHMQE9c6iFJENLT0JdXnvQqz0kT00SfVGR2g
QeVVTyUw3Ffghc+IJMyjOsLgJSczBV8GrY96ApFmaLN20mYM1TuZ0+uv6+EjFSAxFPyHWFLveXku
8mzl7rMdyzLd9l0C93rk6GwGoGjemudPmbx0aS4QM+9N7P6yzxmtQc8WQsbdnhL1W0uCPU8Dkfk/
/dddYkkuYsrhvRD7zXHT/+neZeXCSE6itF7m3g7q9Vxsc8v0doJQJrTmc+E1h0rSFxfMJsxYigUd
UNYeRF8fsPnx4c+dv2R4cmG5VvyRConxz/psammvumHC+eun/BKH4Rj/8QskYFxk1ZPNtzPTjTEQ
rg/xRIHd9dN42rQqmVn+exjqpD1EvxXRcEfWHd/32QWkcK2MgRoVh44jy4ycVNua0V0z1DZO+NMc
DFSL02bHlsHRwhGeRG0GH2uv5Eobm+EhLgyDecVQoA8+3Dwre3dshjbUqCe9Wp5vqWEc9V71WjGf
i1PLZOzxlEn62ACedbEPikuK3eTC4ti7SW+QY7rlUYu1g86IpxcaTkSrLDH1fVIxHigqUYZyu0bC
y3tU7d1MDjDY0TPHD7GY4I8NL2E8syJsCORfIBtP9/jrOw92llc47fJ1o3YXz/tq2S8mPfCIBIay
Qg9Q+izYzjvtlEMq83JQCG4LtsXh0W1zsI/jqSH6vVzzXNmgzjIQkkR0y1vdbcVxHFxsIt4b4zYN
9yUq20i9wtX0WzTdjmOwhR8r5mGLlq//7gdGMHhnOE/uPqYuWbW6NcM3zKKHPXFT34bhHGAU1z3f
Gj5QzKIbS4EVOtVk9AIQoSMhdyYHadNJkeVAp0XOuQBfpRcxNy9mXsNe2rwgyLiwLq8jst6sJXHz
7XtdjzNUcCDUIBCr4Q0+ujUMfvkxC+MiTCRurD4mQaO9t7d5FvtZ410+cwF2RUVhh71nV5Nykx7/
fVK89JZG2QpV2bPmMB/nSj8/PL9ZmDqdlWACUnV3PMQ0AagmJ09HdywHej+7fsPd7T7pWfNeg2Vi
Cku53B21wsLQ6qY8GuX5IeDdRkAV/YGVQ2T/3GleOiOAi697+CZiLU49vZQG3iCT6VCAZGCSkkGD
wGrxq6aph213chPW6QBXBFzjVzSfcFy6KUk2CKy1QBYwcWHkmF1HwjKHoPU02aJPreTI1R1z0UwL
55uxb1pf6QX4alIm4Wwawfk2hUllJIvc2Rc2a2TK/iRw7POOys7zpds9ruu881gsI1dmMCw8vUdY
3UZ20qIJoNdc10ms8Gq3CDuUUkjYfI+LtVBiLvE3EgaS+iUmj6uTgAfB9iJfwBR7IVbxOHVI2DqD
8ffxdieUXwMKu4QwnyIgYsiMSacFY2nLHOA18V+SgobzxG7Q2ZSio7/Nda1MLWpfZzYaSYjWqdtK
nK1CNFkBPIzekouUV0EaJbseDc/Uu1PoZvNiDu+pANv54l40YUd74AGJSB+rBNHGNHEkkdIkN4kz
OYZ69bTHnr31aOhqLrdmNXUtEDrptzBxUMoECWTVgYv9+Sf0ALVQV8Qj/iZ/xKeIE51w4CuenOgQ
G97LYm9zxsZ06UfL33zoULl7t/wENQihJknXrDQXBgyh/tOoWkhzbioEsNYz1m4UF556EUeIyChq
bKAnpBiDhAe8pvCW1jKv0AVi8Cgm8UWmvQ2V6hFIPlZa6aRWkOEtpWIxs8rVlT2s9o8D2O49o0X0
aaDHBx31KVBLj6NBxa17QuvIV6ONXhbvWv31szevTA9PdcbNZj5eWbTchcpDY2HrAExy4PcpIkpM
3aEOFn4D5ILPlRFXG1X0jr6Fe1u6rESYXTO53+4GfxadEpQHden5Uk7Ic2W/tl4H0WE5KViBjHpX
H6lCqOpmu7bywLVfNLydKuCosmPsnxvtbV3fCfZ63zOVsR5NF24J/kmLXIoPLpp6iwyFmGbr/Om8
qzauhY8Hfxsdz5Y5SYe/ub960/85zHOeqdHi37um8/2XzPqW/SS6vO/dg9qhd5PqpD3kllvLJPM1
Cc/uyzC88l0C2vr5EEC7X8uL1KZ4SPY7sKjq6mkGlbz4PcxPw+d/2FW5YgtnqICAAF4OHBkf1CtE
0H6Wt6z4N/WTWaVMLhJNds9f2HbEBapQfJ8eAOP1kLo+tKhfvRo2BIq5xKlUXS4AbD00jpRh6XEn
pL4KteYRk2b6jdRl1wtDyYo0cn5jBquFnKWPhdlbT+XVjJLkVoNgGvaRtk4P0IAPaOjx8F0Gz7b7
d1setH5CQMjcbKRreAwOZx2m1iVbBfmRfNifteESUxAquKmdQM42wdNwtrrkmXIn2AQr5Hj/Ifjp
kTJDFLynu/63kAEk9wLCCpCkovrLbKCDPBQVgy8DGMkvXIIkIW7xOdLe49x+TThQt5+oF+Bb7Pjk
OxKkhk0BvleBegEkAmnIMG10KHq8QMKE601FCyjVRvGMKCU8i2B2C0CCvG+eNZ+Ei1apxYKTKw28
fnD6epm5vcx7Z5ZkFcvdB/qL7iZyevVzfyLQd1MSGwS/VkAgysd15/LtBQJ7Rz6S7A74A8YZ5B/k
iBbrOMAfSfGNpMpT/qjiqI2RnPzgy5YgDaZJrNf4Z62qRtvX349+mHwtFB3AdvgVK8suBtv4nUHr
KYxuA1Gftb2IYrhrnQHw2A9NWnwxjLSekT6uyAcCuZ/LnTigWE3gAuyFwDQlUv44kS7ykw2+o7kw
r+klqj46l7p/5DqcXKWtnMCxgH+5UbaAKBXPVdDLWfybR9B1Y4qh8gXp0nY7QAoSowNTHWlL4Da7
nEPEybd2s2+EUCbUSiUf8Nc1fm6LcqOfmcEYkOxzG/nssMezTv3nBlvBA8sdy7eKmOznLQlWIZSn
bSQcGhzMjQYQONh5can5ykW7riAvJFhNe3E9au7jxFq75blcFcUmOICoZo5t3yq23DzV2Ppa1IKP
pNbb3xHzUtacc6KRNc5uslAkPyDYXlQL34n3ndjMQ8rob5tuTHISRQrAVvf0ZmQyWr+ASdLkt6KR
BmmQ28sVKd6RAsR67dlb9XhiAOa50nlgxHEA5/1uEiuP11O/Ez+HNWha4j7/BnnU+YffUyKPRfsn
eOmxr8nkab8EeW37ooLFbHajNxYMYqtx6IzJl6mk85XRJulHOM/QOThzjvWZUuzCkFN8QqloDXvO
Xwikqxx2nhzDxWjfVvmy6GEjw/CQn9QQV9Xbt5YAiW/wNrB10VXT7odJzT5uzY2aN2SqNJY7jNCc
Lh19iU48Qq06SFNt54XpNlK3wWQQQwS4gGkHtVqhJesU6vxEExfTqn7fvhxtdKHed/oRLms9NMar
kv4VNA2+gfnpkCW7l68hDxJcE8OkpygV16uDxo4zcuBXQMuKBbM5eJvYwcH6ZawAp29SwTh6tSUJ
4I4yuoRVz46f9FhGqjNyXcRBk5eJ7ZYe3LiNVQa++DxW4KDN4m10M+Q6j6CLvlR01ImBd5RL0urs
+hXSKuKXPE+2y3qISlgqCJ+sdNGjtpjTNpUIzep7RFkBtJyhKfBwxwfGSGOuAzJHPzHqyiBFNdH+
ksi2CgaKf5V3XJxhbNddHMdT8ZwO9YPji0AStmkOmLOaRfN6sHo33hLshc9ZsWGSn8FgTladT5vX
S1ubi+nAdtmeyVJmewjO14bXyiUAYTM1elBySufYNh6hn72iRqYVkbzDnmgcuEOSXJim/rEBNsUW
cVO92Beu75bS5s9UBBBhJxAkAGDU9Di/cpYMuXYae+daff8tpxvCTnrOMzXhexL9oLvRucrb7Qx5
mpXkplGmL7+giDaZgCask4RVpDOqXvjhImJ2RZFjVbdfRhN020BYGUV8McB8SOobPy+umSrg6JJ6
S5EAjn5CQGvIkw9lD3dbLNwqiY5M4hYwD/PZtqvMD1jVzctG/3xfyXjd5fL+ddvmICudwI4HxBTV
OBVEqPGuK+s8sd3pDY9bWl6ghZOEIXC4ynMjqjw/V0icVuep38GJl/SbLfUvIA+RmAdCgLxEK6ui
rRGyc8uaWD1EhJ2ncKqnsWMAXvSlWIeDdWEwsdZBYtotUFZMxTt9gmTIXhMbqamo/gGbKUzKfKYa
UKRcYDAlHBhstdLSTeNSHDW3ug2njwtf2vDhA2JJ7V0q9uzD65+PQSZTFMM2yPn+3pqI9JFH/aqi
vICGRqESyFzOACVWXrAh7YIreVBexacfgz8l4E/3htj8B6R7S9JYiEng5O7+9sZwf6ntUG3G6xP5
IIbZVWgXZaJu6tuZMy2wj32qqsJtMKEIcTU4EiJjICaFjZedigxLg3g64lgFlS3dWnRxG9bjnDJ0
949ykqrucLqHP6xxVRgUnVmfouzlkraXaALpU2cL5Cv95nfO5zB/YFG0EQUmsJlXQwtSE/3TnFVz
8f51wNmfB4go6fXTMY7MZ7Z74rdxg3WtLJLVgsrtfKiEjVjEJZ59ukY5xT6o01KdgRg8XwMQL/WI
V38/O9aQLMfLFT4HfvUII5UqejgKMkBuwn6Hde1TPvbAD3BoDpYyX4MLA6m+2evTsB2L+wIB/qmZ
9sA3kV8VvjBltFH4VEIBnAPGuNZrE1Fh6EMZnn1/vTEmlWvzLa96sfdoQAkAAY1dtlqsZnYIltPn
hUvw6M/Dmafq51q8mXOyT0P8ufur2e7tHL/9t68UyaEqsl4AHvYCbE0csn1xnmzxubgneR3y44Cj
6FqOsVsOl0/2yivD50cOtr5+pzwCs5oWz/K8nznppKBR/94fcCQKbRq0Y4VdE3FoxnHBuVWqFLdv
X+hLUOKaL+MNDwi8w15gKb0H9GcsVTJHAfM8ZjViMe352RHamf9h5il+w7k5gNHJ91L83NUlTIW1
yvh2eaD2raQJSjNlxxnKSPoOp3yx8swfx40lIxGkd4+Mn5sy6xKDyGSNLfm/VnwqAmEwmYUDD9gA
LXJuZnOiwbvbzyt1fBu3Sbr8dPlr5SLISJxY7xuZtlsDJHEZX1dRPaOrbq9gkWE/27zVurrUkmF7
eJ82ncL6vpoW9Vl+w4AYgUJyu79s/H+1TofKzw3/KtJ6MQZLfNseDh12L1Hzdd4NAQx6IQ83NtAd
g8n7z+1JFHjsjw5coYcRQpDT6JCq86Q1YZry7SqOyDbWBJOGbiXnWZMa+SnpBp7dew4hAF6EsmW8
mZy/xqY7uOXQ/hSjZejZz3R4zjB5qIzLpGY2Zl9DjyYuUXT96np70g2PEtQ/Gm5ROFpJDsKwUUu3
7z67KVxGyxpwXoBt5i+XkdrNs36H/IYmlG7saVL7t7ZeA5Zm+6TJFoyZvi/vEez5jRQQFT28wQZo
xMTbG4lrfZjfargFn8sPeZe20rLqlL4d4NNNDzEFckpPCPdSkckM3ujYwEQFKT7Ien+WspWydzrl
GIm/lW30H09C+SDZrn1a1BJ+2DOfAhRXOYE9BVRGu2Q0o2Bmo9LK8tRRP6xCUXRPfMn+F8TR9HrM
uhj/HOlqgXeCcea8lAl+4GeI6bv2sw+5eFBy9BJPy55GRQ8t4kg8M5ExIghBO+EzQOMw1q4E/nX4
YTThAaBz2QkD2RcncDvovYivDGWbUzEvOU5Zpm9fPgcdqxLHOS0HNwP2nFtxB3cWETIGPgKikAEc
RiDBoWkHqNZbMKi4csGP43etnUsSvCWWlNKhRU2IrDSoVhE2sIija+s92/vRUBAZ6f6G9ajV4jAa
DvtMGAfV4Cs449987wAwlAwHC7kslN1b9lvDFE8zMY28n3xW8YjY318eloK0Ty4+C8iXHa1+b1fr
ZHvP3eYmYC1sMPu+BFjO/CG2yBSSjW+NgH48+lHaJ9XWZkq6vb/Ktj2vJV/AO9XzShLr8V0T2vwd
1IdpjmUpLgIZYRlK6FVghCnR+XcCR/PmZOTrO4wi1cAzeKXUhU+BsUZjTURRj1etU8TmAguzd5en
2pLYQVJWc9B7/wuzEyDTXF2G4Rl/zUprYiUBoUuULhKOe2FUsLa65ZXuxVKem74mfSi63W/Of28/
chK6jJIUf7rMT2si0CYUNMUCpB+Szq8vWZEQQ6Jronti1fxDvQY6YzXWasVS8eq3psixb7lfHcmP
oYDe4lKfhMxS/Jgds13H2lQFYWlWlx3Dc2ftS59VnEf7mOl/s9PoqrcQUcdHzxY4GWMySfz/Vv0Y
Gp5S/dwHnDf6iGMgC+hQImLtmRUP0DsMB9Ou2QhBEwpIWdzgrg4z5gekF/kynhow8aKJQa+GPpNm
qKDyrfOi2+DII4MiWvs/t/RWjRfAgMAlRocpGHFBlDUF722ZIzBmYGFOzO57odKnWh9nLofni9Y+
nZax0IdOrjRTCAvA6ZSmXgFegAX/TrLbYBKC/LoNcXKPIvM0drO0yu0QEXP16sPXZMQunKIxzR8R
m/V2wivEofdt9h3aZTfwJ5nR/kaLkpxnoJiAG63Jx/d1GhJcVTepf2J3urNkFmA6sJx2Te52q2Yv
oTriGqawbT7f09hdcBmT0uU3dyLzG6IgDDKI3kzyKaiYis6dLZnbCGRMgGMy00QDF+EA6OmKPcYY
drS1SperrMxGiW18H7Y1w70byqKmdwmCUux+hPzux5Kia0i2gwDB7wkVuRMPTit2Bw0FRCRm8ATa
SGTBdXuH9Gmd9Wtv3C4OvGC1AtCV4DzX2cTfiO8z3xqo49F1ZU6RKco4PkNH5zaPesdWwwB1P29m
O3+fyrTGAZq96CZ1crAHwsnTl5WtCRBdN1BIQfjLc4P0VNa5aKm2lIsPqYTAvNBLUsj7zRtyeWUl
E4ldY9ivCi/a+0mwk6nCmakjcB8DZe54mH8vDHO5LBivDE1QO41h0qzR8JwkEDSF4kRVQ/ANtv7A
p+hp/w7xKUEs4iQZ/Xm11MRgs4+oZkCKvR0wnW9f1Gdbnk7zoJii32YZ5zUUISqWdQO2u47b7vnV
9rDXrMfDPFfnQFlT00JSh/7EXRtfFdyGwjKoyeouJ+a0/fTaAmL4NhzPRhkjI5t//RY3Qd/LJOfC
00MSqyYiDy1zpVyFu+I1mwboalT+vIompypMmKm20GhL4/F1ik4jjZbRGZLUw5VaruBpWFocx+wD
TCUOmyI5ncy7X+YnKRpBv3WYJTH1GfkgRQ5N+tF9LJSsM4M+J8XeZwSmHOKNZX4K9G23vC0yGA2D
BH3AMu9wVsqHvM4oCg9nzxssa8OBboarP1fjDebj2tA9Fq0UKwmlLZuz8nxmqStKBh8GdGXhl/hh
jlRhEbw2sr9XORs8PPuAFiUDUAABoJSvMRmuHmic7ewO/XRdriCxnq3PGkECEaowffncWBHaJ6ld
GzfF8TjOWeJXfXfDjZCVal5/8V6SQifr8s4/VvPNyA5U2yciFwyaEOohH1j+i6bVXytVCphERDnq
TVj5HmVNU0mk67LnCLszjObs062pe1CAqEh7KfWFSFBT6gVdh/OhU+/hJbJ1FB808Oa3PjT+ld7O
jTp3EZeptJ2Bp8y3BMkNM06IhcBTHiiPphsZJyj17YH58JV3DxfK4wv554y7R9ID2u6rvZRiQlv1
Xqro8AIBD7LS1vMBYlpnCwtw8++XjE7Db6u5FeeeZsVt/ZvuwLf6wntH6RH2F9d7AVA6O8KnLgq6
3dsRdQ9J33JHS1zUL9JfoK7JVVNYpajtoKYvIAVeRnd399pdA3MNxJfZGICkqcZ9f4ZVHprhmG75
qztU6zVHHMeL9yt3Rv/73VlduNqQx0AX/4bd9d4HIpAfFAXMlAaBzu0O/ZoxkU/ZWGIQano93po2
1MBauwVuk5VyglxieV2TExJW2ohscNT9mlkiBtmebBSI6V/4ZN7nEr1Z2CMUIxkQBwkMvKV8HoMh
m9JFczShPhOf8JAixIzWh8Ur02bUHN3AuCRAz8tPTWoKt92fKmQqt1wQITndASsg+/3Na5OZhYJc
MRblqq7cwonUoGsBHsVMVQAHh/Hl1/ABoZ/a/t4JMDAOlsjr+ReJVWgerkZkrXgJzjkXk0qZnNg0
A9j6mO57F9YF5hdQdocdtCJyzPiErlSfTI81lbdt8MRvE8v4pfj/Bvx0t/XnCz4u5DSYxRLCrwrx
RGqMHgRkgphUMubUJ559JmdeKSy2saN01eDqpbJyXKSr7SH8tBiFC24v7mbdTNdRrGPfx3xlDbPE
1ky1Oe4iowv6N684I5fvUH8AQgXW5Ddx5wDa25LilkNSp1rjhyeZZb+a8tWsZkIPpAmG3QLT/xnM
QyMs6S2oiuY7F+mwsOLEXmh3k9VPsBK5QaP13W1pACD8l+vauWmKdZnTMjm4+ci5b/5lDzTXMywI
gI98W0lrxB2JyR0g4VUM4SglhyP80X3xPtcJr9QUB+hOv5wjzSEyn8mrBH9UbAndHwx0MU2KiUvY
rYOfikuDzUi0Xdy9e2dv/h/95SSiljF/QtOBCpGPdGGKpmcnu0x6+tavUQ/tFKdRhRtJCWeNoqE9
/gRTLLHNzi0rU6e0YtVSAR5e7s8AOVkMFz/8S5Ll3YXA3CghQ5/esDUS0kQ3hLQubxldRpH12OQv
JDrgXBvv1oa14V1fS0yO4smlC1M7efDw5iShEcq+6np7Q1riXFZEVgLz28K658Sz6vKUdGNL5qK/
kC0VHO1f8edKttIhEWi6I2uv46xVjn9EGt7HyTFFg9DX7KuE+AJbHcvKXOsSirGaTVg7u3s0sEMN
M4Zr+h5JRa4KQKr+qn/54sLQIXmS41uoMXBaDClu9kxDFFzMK2047fLbUVbjNayTkQo2PqrpDe5v
6Oy6dusb9bNLm49kizeXyFxPewgXMESFdYbqSO+qwMM+JnkF7A7sy8YRq60rXBowNyhkMvTVddUs
XpbQkKeorLTHmhfOGxXOeQ8leVlMrF9VIPGK6dEuUM8eGmB8mMQ1Ul3bv7KISiNYMgH1QkBFpVhB
0c6odLysIAYIDS/26H8blADeUeCntTJP1Qepm+nhHkCNf+NxeZ9GJHveHvwht/HkiM+D296voOV9
3zlM1AGIQzzJbydm9tnsOSFrHCTVJO8/36J9TeZXG7phJT0xSFKepEL5iHvCc+tePdWqp/fLD4Ve
/sJF7tsj5+sFInykHyBc/uGw4GDINjXdKaEwD1X2aJhlOVSIbIVOydKaXnrFoK/Je01xxhSGEmPI
kepnwNhxXev+KRAmZ8G5dVx/W82/71SL0jPC9i8IKdffgadvGkNUWRii5OsUARpUeHWKlMRqs6hy
nXraD4c/QamO9ckmQdrlk4osaflyI1sM6WEJd9Wfd1mFtUZpvb7ZtbHdXYzkWXxQ3v6LrwlkcCyS
Z4U3WIb5KD9Ve/AXdTYTxH6XZUXB163pY0xXWE2lap412Q8DT+DmOAuodYrtgzZ5jGAAY6XtcGlx
qiTuOmCuz7uqUxwC3DXBRUeuHGtYPRF0HxGIp7Wk4KpwyHFN2IiMh+KFoE0FaiETWk0VZAvkfq4F
oqLVj+W1RmrrmrN8pLV8pqXmKobL3TPXORn3I4a3dCbGLT0gNzZD6JTo0NYZJe8rd6j9LLUKAoCh
b7p4+tNkYK8/3Pkj+vx6WvKRhm8X+944xiZ/YjV4mo3ePCk7veFI4xnfeC+Z1Bjkzu0u2yzjkbki
nYtO8BS4uZem5lotNF9xLbbv5N1t9BluicY9+N6tu4S1EI5sQY16OBe/CuiwoEZV+BfDbK2SOcj8
/RnR01saOnrrCmPudlhxCa7fBAZmDynMWWvQj9Z/XNAlQxfl9pp7/nC1cL/QzA3KzaFr+v9iI7WX
2aB33dnaQDp9/HsbFTTzj8WwWwPdlLLDH4VP0hO15zgQPSiwaFKJvf7AOcj6g13Yo4Z350LgaVKn
FcslejWKRKjToZnaeNed6DBREe7Cqc1WAx3dXohA/qk5VXgJJ2KA0R+k34DU+f1mNq2porsLXy/7
95SrLuvPm/yRvYJ6df173NBL+askv1L+RWsiNvXziteSX64Pn/U70XBM2ZnMktj/0mXA1X0+un2g
G8ETeILdaLZF71bNiKlybPRdnPMBejUwIamXU9xLHXS+f9Y1XCaCLQ/wZa3WUEtsef6LvY6Wo/jC
3BRwdr4I1tKIPpTjQjwZ+gIairZq5NMRNjcpRhJRDrS4Eo3hyohLXoUM21v5Uq8X0/ytsFroa5Q6
PHQASTRll5rxIyi8XK1L/bCFZzWiqhY8ENneHQ3Y4tEeB5LqEijsQilzeBOGEca2s1wFbA9UG8Mr
DcqlyBWZ4pSteR3tqCwZAFE+w/csN5ALJY2e1Nfw+NsxI4le6zzy03Wve5huhikKdnvvgiuMkm1y
NW7AqYoQwhKBNoS7dit+SOMn/YG6uckqXno/WPaTGV7prfh+5uvqPxzpVBsP0FzqW9jl37sf04Po
tLSPn3weU6oIGr6gMFzXvPGTnVmn7pnem3t1dSOU0aM6U0XriU+UQrvZ6sYG1FQkotZo6r2xyX+s
XRMIfpFFqiCLGuwUsQP9k3lUhosu7De1UXiveVxc+OIkQ39bSMnbMQm8NW02JHEOu5v2/yH+fKKa
6yFETJalMjYvBttyGvkLs3zFQGS9dO3K+FKDEN3Fr2urq9IA6azB3Z3Px3ol+WMR8CAV9AsVNj6Z
0avPIX/1HnKfRdLLgXTz/Tqmeb+bW9B1t+jBYAXwAhXApdd0yY8Gc2NTnLmjbCE4SaXZmbgkOv0g
jDbpd6M/i8y6vS6GCrnw5UJp5ZkgfRIia7qj79dGVg3f/fWpYNmgqbXW3VI5qFt/s2iuqUArr1+L
trYWIbsyXDFJESe1SwMehBfeo4x7A/C1gJKgHfA3ccJxnlcy0RLTl14+hD23oS7zbVWA1cEQbjxJ
4Qfrm40Pp6DW0BhWtIkNIdsLK+btRwTfKJDyDSCiBHtCexLIfm/TrqWj6E2R+SBusXG4gfp/kT3f
Z2prhM7kzkdi429e1u8ZGeTgdMfAmgRp68HHMaSdeSqu4aP/419JzX1m5xZ60ON6YH8phJDtePmv
t2kXSBQUJ6i6cj9T4Lmc/NUwz1lbwV3+FC4jicwsQUFMFAwndqPSfOfph7RFUMYtB1AIldvZ1Z8o
Z0XNvEodF5Rk1Bhq4rp5StektB1/F6SCH8pN/qenWViCNzZMfpKLD6fvtzU6uGUv2/yXs1RztSYB
UA8hU5V92BfqnT7Kbe1PRPVWmRIUbuRdseJGW7iC+P/GgtdcpNnCThulG2C919nU5rEmVR4i6zzh
ZD0KfvijxlO0iRn9aISSBWi50bDuVfYxyzHcAOKViTOC+M8jWFmbGqalbQEtMf7soQcGl7POLpvw
xgLMnMOaVlKcRLOnc5p1qP+p5wkC+f+Ytsy8LzA2XctZihQ5APoDSsOfnL3ibNsH7bF9uPK1mb99
qP3LDrrLCMEvf1eRFzFRnR6Mk2p2jaxbiFp9zl2iiGLFZ8s4p4lYLBJXgVVIQP/lEBSZI2/rjoBx
0Zx/1WEY2MNFx215+iO8DlMCUrjiMMOfoweVW0QnrPKB2tbAD/TlMjf/65MZEmwzSbhsD58qWObl
OrqvMTGTUZNxaQGbq6IHioEZNJndUfdQCDlnTPK6iBwoRPrnlRlJgMz5U/bpd6qPNIWQ3c7O/fC7
wdCHNZSTqjy09PyBIm+J5/0yfiHzeoyKmKP0U0DzreYbwRBMAAmU5GWeL31RKh2sK4BSeJXy2JkT
LqGtoJ0LJj5RW3HOo5ngGXswH+R3si7RzN+gK0S3y3RSSYj4ImoeLzNeVkl1cgAnQcfb7/9SFpoq
mBvYIXgscrG3u5oxUPdGwE0dfqrlFiawYRZgCNwdUcdSTvMPVc5c4qRRQ47hqAWTHMSFv1ErrfBr
kc921+dvTs9kOcHbycUFzqXAMQDN9a8xP7HQkkvYNo2/n2h/YgWuYT44EHnQM0oZKhvfnrEslNYh
ta/NuoMThttJS14u1sV5KM6cGyNuuXMuIUoqzZfE8wGdfv90GQ+KN77WEnsqMjDZXGd+XJGxLQvg
GHVZ5jtYvn9deihVt8pDDQ4iQO/UPYN+r3X6Iqu9i0cmtAXSYti/lbXQnD8UWtDbCbZL80wG/jhH
+K5ZweZ9he6sdTjtzgU1mUgoFFIebQwMKJbdZ8mXhHeVppNbbt2h9qBdi9VSlmuC9I/NLT+CVgik
5bjvqnZLvtkkTrL33RIiCl7hIZrXF3FZ4mGGAw6/fa9r9SH1lYxTzrPAhBOFrT/ZA6g0IuvRG501
SHPB3lEQ5OqJZsv3Hp8ORCL67NpIklaZ/dCJJPou2NSGOEPcdiN9QWnxekfa37k1fpdN8IWV0+e+
tEUmjkt9SPLU9QzDNsoSJUtJl+QblKIgfYG30jTQ/VYUTQDC+oiHcdZckaqb1BUJKEJKRAxIRbkm
RgY0WRmsnqe0XLotLhduRBruZ3OhQ54oGTSVfNCi9+nxBrE2ywg3YajCMl/C6uy7CMYShjgKwo3p
xCVJVsEX/eEs2EBS7DGlyqYPJoH/iSOG89CVJagNxu5h2StPTgPQc+N+eGDs6b4xJISGrkJpdPuE
BEx6oXUK2nUEs6MaYGgX2VAr9V9QVUHxeeX7e3YhNeSZoKlw3I1lUsL8RIJ5el4M0yIy10kMHt+8
taJqjqrMZEBtxJA6kpV7JPdfzV94F61X5jkI8caQ7gbGjRlgbI9qXhkNjCsdhglfWf9qOkgdM8tt
lbTRLQFxGDAtCAJFe744FT38CMFppsVmApCDEzEG5t03ZT+kvf+KBIarzbr7xa1QgE9uWZxoavHv
RSfTxZGLWrmbMSCM9e/3oCvZMWwYJFaC/WFVUdoLc4358K5gv7WTk0SMHYIj6FSq7QYbGTrFStiu
Gf0EU45zPpsr9OGT7Ui1uIEIAxED1sXEDs0QI0rTHsnP/JI2jhlswO+hCTr4ht53DB6zi4MXgtjv
SJgY+urS3oVzLAJ++aIBwlRe5CoLJ7AKCM1IXtUH+wrcLUATuL3Q1zhaQld4HukeG6VOkHbqH33E
ekExg7iKNkc8XeMqxLz6K5r1DAJDpFDGx3hc2IT5VsmIj06+2pIf/Y136UjkCZEjWqRbjqNx9yMF
bInVOJfs80lGgGRouXmv/PJA9FCngU6h1ukpdkmyleMFfUXADyXmgJP0bPC9OmIHUY4o2G4pwNuO
r5wWo1Ggz4d77VJkZCEOlRIYhsS/BdCLERJM+Xuz4UgEirJflDRgqaRHvtw4/SvAf6+BvkUbGCx7
QQXI8ckgdXpRur54KG9MrvSNi16vZP30PT+uZ+HDrfprlQF1PSu4k/rsPeSo5MXloWi6f/0OKd7t
V19hcd6J8ca8ofe6uEdYM82VfUshNr8zUHvupjjBFBpYocZFz4U4DjDMduQxPgo2V//B9xAce/6w
1PDjrG3pIWZpSM9n+RWNptYfqUaQpOz1MZFfJw94u8GG7JXTO/3NkVWydR1PbYCxwKMgj0P8xUCw
O2l5abzKsHEV/0jcb6rECd+CVLaHkGv/jgSbuhY158tuiwKboJfJ0h/9uw4uIyaMDuWc0G9Y0H+/
8ZkgZqXzd3RUmQgPw/hBMe81jZKgSQ3L/yeeZ5sA0XhCKkYQsHTHtaXs71c2j2CId462rnms1xQ9
8QLfHKSMQ2X3Zj7t3lJK+mrlOfn47AvtX9uPY+W064A7cVjrTE4NtLcQqEQhF2NWOEHybkg+pBHd
V9ccPQw5Z4LlkXvzGywBQpDmLnxNLJorttWrGl1HTd+R2KvxvMw17K/5OAGPaH2EJsPJf7Rk/Car
inNjmlzk6To8hcZ7StrNmm2becnzAISDBkZDiKFGzTe0FOVtwHWs6pk4G3qLiZKq3eIkao4PrpEh
QNLDdIDfB7exEVZQmt4C0Ll9UKquRkX5avRx6XQXYlw5t0/6GqJFIvTYJLtR102pFuM84zUcAhk1
097Z+LNgkHw5JYw6Pt5CkCKFOiU2/ak7ssjNqgAar3NUYvXDVhF2SqB1K3FfBzB7VdQuSlCmMCmq
ERVLqMfMBO5SuiY8YsDlAgvSCDJJW3IjUFuAfoZ/x1qCY7EwpHbofs2uP+GsCa9ME4sKt9Lo4FLP
IHVhWMqQz+vU5Po7ebIjPanSsrXZH4yyKn+4PVOJv+2CNsZj3FXlJVRfrfU9eg5EL4reaGWV5NBA
5aUdRr2jZDea3+P1ge/HctFs060gbajIkmB9eVck8qBXG6q6vryOR93XRo/Mv8o0zDqDbSZ6T9C3
9jyHAZQyXSLRnAKQqGWEKW45IWGjnJjaAxRTFOG0yKza/m60QNeBJAKCrKz3HAM2sTnXldZWvuDf
tHDPFjI+fQ3ufvQol+V0HU37b+Sj09Q8JeQ8Lr8fxL+oRdU4Uu2Btu84i9Jhm9OpdovxvdlgyPO0
EmWuHdgNIq21vLNa2LiT/slhDSTpZ/2iRtw+x/oHP3c1FgIQAZjhefv9+OGg07zEyGcxJCHUrOtL
6JPivfZ8XyUe1p2eFL9YOnigSpP2cdqGXoH9yMJsgoA1x2LhvmOBHo3OYa45e68/RgfSFyJ0KQ+j
y5J0uCQ3LEdmozxLC534y5O53x5mEoxQW7essBM6Ws3/vHsh8HDRIG9t81sXxwvCaN0TmoUQaqDp
ExAZyWNhlGGczYJuFq8x9C5oyq7Me2rgF7iSHyOc+m0IQ1GWejR2pDg56MJ2oSFanTA6pKHfSpXM
lb6+cKf5MU8HoWsrZrPNdmuiPxdpWpEXhvGy0sQs5m4LAOuVZp9a4iCoo0XqXTuhsiJPW5Xmbkr1
ACOnK3SbVXGLDxdkPT8L70/SO17tERewAPwKzvlXFf9gfFxIAGHso0A13cEQJvz8HH5EVtWtkE8W
sYnXRIcM0cZCiPWSaXOY0exRSBiKvnALFIzFhP+P4GTxaI8Q9egUhw+aaE41jN/W8C5fojlKzdqi
XSQwknw32Q96yrmGUkL+ERDq5o2XvoBPQCPJ1f9YQFmGi9/GMGH5nXIBBlubiD8RsrRe0rh6qvpi
g0GYjs2cioF0aq05RHVTUSkv6jT65GdFVaGLJtoA5RZC1LAbBYd/gom9qQevBkzj+bM2PXaP5/W9
AD4FcRFrtUg3LFqBs+yM7N+X+NXKOOwZ9VMlmg62ByTxYWDvNTgkz1NTIUKCe8kEAwjvknxKBX8J
ZYNX8Hyo/nlW9AowoxNHcGxhFwSrnUA0D+M6LRkQGmTLxFShFd/GEeBUbAGWx1J/XzOIdd2IToAu
fGZC/FYTRc8g1wfTi4OjB7AUHNFVKZ7OuC/j6to+PQ+5NZtwOrOExZYgZe08ULxh2IYLduyNKfJy
ZkD9V/nymjog/vvyIxqHnGXnOt2NJHEeWZkVW5NakFlqpjRt+fPKgCfVQFe7BnlKQ0PIdf7LC1/3
PBkR1XMvzFqsxrvMEZWJsnB+v8U6VAcA3NsAjjdpTo/aFtWfGw3cpuUcLmsB7HXI9hDa/ON1Ucfg
58xwU9w9feri5Fvauec2lpmbz7oR3l4qIU3AOHZzghJVaWLgDuF55iXndx/kkqsJBH/DrzJviHf8
7FXlrCWW9dGpdusexETzauMSZo+0TRaN8blp+dPycuIb+0zGSJvXsZ01JyIQ5y8rA7gZyN/G2bqc
y7aGRd3YH6H+orZNCd0nyaN2Glv2Ko0EhcxXG3+eISUwHXHQx6orP4j4SaIf+Gif8qyq1jaTEZ8A
1bAa5QY8o7m4IEYbmvI17RQH90OBVN48V9LFYC+YQj1QPB/W5FSyf+jXA3tXobQaJsmDyTqbKCqW
4ZHgiHqaVxvniDcR4QUv3czsJtVKlVc1yKr5eb3F3Hn8Qd7iVFPLvxH6iaU6yxrqFBYglJ8tUK1m
4l8jfwZFtZAb4eEdIpizTQh9imlEH/SIs8D3aTuBkWRsD5Fq4tzC2nPMkDHmqlVDt7/kDwUwS6sa
M55K72jXzC1d+Yu6tNWmL78HA4LM54cn2lltZ4nz1DajbLzAchaNrmfAR0i85nj59tCfxsnxppMK
xNrG1r9zILivOmkn1XsJPhivKY+aGhne2fFuSDjBIx0qa1kMX/OLvwlSCsc5GLMIh5hVBsFRXrgC
I15G0pXdds/JKHBIm6qlZtE/JuFtczsuyzMqRdDdl5hZcMQGUISZE1eFaOkti0a8muCmjLvyA9BC
UyMBNmrb0Pd7W99HTUqB7vYWLUFiCrbBd2zraWBYRYeuZ9dAHSep9Pt1CxhomWpVwakrtBj6oJKK
Y8yu2WVIWSmhrBiFa5mAJR88QQzKdRcXHZbFb5o1o/L3w/Lb36S/ypuBH8LBPNx2rapQM/ba61Oa
dlRXC/aKexutaqyLIJZFkeuKtSVTrz9AfqDzKz6gyxEW9l34YAelp0IqxtV/kQmVVbAflctVmYqm
SZ2od9t9q6HBh1uuEBcCR0hibLQCNqQF9OVs6+LtI0zuE/k/pMShot7m9M6u5L85SCEcq8iiHmuT
nIlPILgmjq+pEA8d2fWe2VX/Ci+9KUOtZcENUscvfNzBfaBR0a9NNyDgqEnwBe0D9ZoDjMtjO76Y
sVuM8zdjM5WW57NMt/6aQAy0MdLuTIDAs+XxhMK8sYoHOw4S8ewiqWOjA3Og/dLVcV1HCXukpF2j
Dc6ztMrJNUHA2jBGL5uXm4Mg62nUC2SHMfvQXZNoHDGDv5fPh1i3iII2ZAoWxmUUICEZSqrx8wGq
4mewhULU/jNvXDBkBekFJx46xzRawQ+4CK90MlbSWpGj98xuxWHKTdM9ov+d8aD7rPm96SAMaT6k
OlgIhGJHH2sRt2GQKuryOF0ZY82C5qZy6YvehzkDlCHuMKA4bGLsGFTDmsNJgBlcSkpE3tNZRLl8
gtoUVGoB8y8fojOXFwAC8X6ZmsRtB9s4lBBxydaDWro7254jsVS/MgDWFxnCd9bwdQsqToQIvN4C
cU2OXeF6w+mcWBRVls0fLn4ajiiOJHCsGbhFCPBiXGOrYLYUGxte6vaweVC7JEzIfPCnvPmcVb+n
QJmxiymEtwf7TPR7Y2fiyokqjSOjCMEe8hJhNcgCus8C83acgBIUt6PIo3UNcg0LcnCY3XIPgouB
iHV43x66zR0hrHTKTtRCnhcpr11N+CAqjvE9sYQaqhrzPwtRD2UcqPpg98XGR3yKBH2zmiN/8lDd
KiSGlhcL3aewy+uc3A3jPXt+l0UuNuVu3VzfE8AR6o8iBtpPtRV6kXhy2F3c/B5FkgC51/6kMdXX
1n3xT2OsBKprDeHTlPRJRUlZiAqyv4Sg/qjjpEk4vAoOy5fc5KBp8NZyLVLkU5aTyRv/nZNntxsy
lWBmKf1cfqvc4CPntHqkXTwS3LOqYHZ7H9uuM49BqIZ2XyWvsmlabpUqtQToNMmOIsHEWrro/FGu
VC84KRG/taCffRMhsCI10PL0od0Jjm9fSqgxjsz4PSga584qRYMs8dPDInwybjqw6GMEPTCW+lnA
QwFW0lkT5RSAPN6OpsNxbB9WJEEYeS7aMqfGHouW37JhNm7LZulAZ4uifAeI9dRbylpG0G5P08AP
Jvq2jzWWehXcq+7pxm9hrMbG2ujx6kZHJhXKOWb+cBQYjifmoZN1GCb3BtZQGWKi11dt5Jj2jHhp
7/onLqiAXVRDbrc5vkqWelQcn9HvhY48Sk3LnMN21eZH0fL4o/4zdC4J5v603oumc5DAbz54WIq1
UG7LLRLsNN4t5pIu9wGf3ayVjjxBvLfoMdvIA19SJqSSO3pbO6IJi/5VsR9jHNhGmfZsIsd9AXza
LFN0jvChgiVbBjwBmMnkaxgelkPnEHnz8+VkW222AmZ3S4gq8+7SfOEazdTfatyGuWs/QuVTD9A3
CjXgTYSghFHw+3ALqNNoiR30ovU4zdmUytE8O+fo1kF2aD/IXhfbtrLQK2cXfgyzfxHfAFNhMguv
BDRon1l2+1UtZFsmlf0BCnAKQJ3eU+g0EmALUIV9Cmtfn9DwW1nuVsnro4CJPbxbSTMR5sF10ClH
xPsJI+4s0FYNpG9VNkQ+dflksBci6gFB/aNlq0/gOzRq33E5wF2IrqbjKEq5hZ9OivMSAxe1mnFa
Spkef2UEyY5bLKaPl99Ns+4EwfccJHlmtjGIcrrr0clmgGDK+wHChh4S+Juhok2DcXe9ZJ4cjAgC
adOr82jP30CqAsxH8gkNcetem58wXWy7wRx5D8slt47n19JeplfsAhd6k6+ONWhr3KlxF7ki7eSl
2+/tY8trVWXFjMJ45MuYJmG4MJgTZ+UyUIx14SDFoXdaVHbTvKR8/rRvEg9JPMLUc+c3b/xTreTS
ZDIlYQ3eLfRKCVVGIKjePM4Gz81wtUYn4emYfe916L2FCq3/h1pzEj8AbHQxqp3LvSfh3ZSnDFdm
nfDJ6EzZQ2Qt3v5fXBo4wLx0fQEL9VfV0aGmPkMKorFRzeftHErlWda4diGqFKJHofE2oyYDUDUy
xhdCbvyVkp4T/1ODEGCx35Zv30eR5OukAHo8YcqsBREgx7rw2xhV1qp1xA3EmZ9Zjz5B2RzNpO2s
j0ZZ/7gRZ6X73pk9km7srcfMNnDAcVDKoeiMENbezS77aujT640zTyhi+gQi1ouaAY8suJFjYqm6
ysvFuBJ+6NCb2wBVp/e+oQIg1KYbUBC+XT958DDsTncmXF6306/Qf/jwSeZ8Et5njapnGR/W7lrG
ZPblx5fgend/mhq8hjN5YbI3kaz30ZXQJAeiXkRTdO4J0gfmnHkVc+AV5elwQJL9plTi/NzOiwEP
5vCP7tdM0pzCRfWrWDHDv6rYsRvedwLRsm5MecXCzyJwO5FRxJhWAwrTW0Ez/zkMkW+uR86JKHr6
P+HyfZHgCFi6kDJgeH8u856Bq2Rjnzpk4Vd5YrxkQsyevepEGN3Vuf7MOwqfkOnVUOu40kNdH7un
UhEPt5X6LMlmgFr+VAGdZ0kui5+7IiuBBktc3BwreSTVa1dnhW9BNgaM7+IG4cEOKOBvfPoVLy0A
XEZtBFU+f9K4uK76F56i6rqqZ8MkA1aAOyeMOy0wu2uYgEtMbFmcSnhfnQV4Oivvplc0+58CP0+k
ouyoc8aR73SI9MrvoyBJx1Gg52wazjekM1FQy9HCc9DFw674/73K03gaVPMPm1Y+0fgtfEkc8eMe
bnXlxB43qHOSF2JB3smUQyAP9MDKHL0jG/5sw6LS/idM3u184oNZlUOmcchFDNB3ZGIHXgt0ePPZ
WbNfo0nn85GsYMsW5fMytk2aZMtBU8Vi3CkVbWSHd17dmfzWwxkbVUzHxBwrlHhXfNlaAQ+YvDEn
xk19UGVefXwRu7D0HJREl0o3w5tEyrot/wVtEEfLF4QELVolGp60Ua8ECnq8041kStG6/Y5WdERf
Nq4odwVN/MirJzsYRualneW69I5OUICM6GrxqWxqXl8HdbR8Wph6D/SjxVW/MpRDkxyGXshTWJBE
wtHqFwKLRysRH12Yx3LQuYbdt0MlWz2iBejv5sBI4hWyLaRp9NwTvetlbK+//cBgdnyKCmAaBmuU
nIQw90Rhf/1dhKR0T05N5pvLHJrLQrTYMMDPAMzonisfwZ/Bp7FXBjZ5wjvYTjyQGgFm2vYYZY77
5A6T/NpqVz5rAUE0uRt9evHbpQkTOa5K8cHmk9dalx3vt41fmuMXQJJqPTSaB4Nt3ow48WL4ioB/
a6RD/YX5s0LEkLl8MmHlH7YeG0OCl+bui9RoWi9SqM64iGErh/EorH53VsuVG5l21DtIfDt5hKGT
f6epMtMA90yShYyRT8gy9paDfqqlKcsI2fo7CD2WnHlfFNhe8tl/uXNPRzI6vdKkWtfo0CJFYKAX
OGcruigtrjESKnWVHv2wElseeadRfP4MJkZ2DMlxD4yNJc1UgXXWdOSXZ1nvIELjaH8ggNuWiA2H
alBRueFepKsRI0xbmpSvtRDC1tZJpL++IgaYy4IAi/ry34OrcAJvMYNykQ7pqnwtHICFb76rFD/W
exrNsFv4tZpvp15C1HTtnEYXLVp8xF1BYRHni3CrH1/a4W+eV7QY8ja+JImFQMvdrHy29JxpJpQ/
AtptPWVRYyfQ7Bvuu6hxlCT/Q0hFFXAX9hcL+TeSU8RfHFvxY3WqhRQqICNN9tzYNoif9neJqC0c
N4qT7/JOPsfI1GrfgM/eijDE/SbFJRtzH+CfK8R08paelZhqY3IlVfBsuRfrhbZJXsAzHS4buDdi
pyvR/uqXyjIo8g2BwovXV9mYB5wFs6CfnL/KBH+ZKbihvlCg14x9f8KuIToOrLvDmn+0XHn3em7p
8kdorlFA9jVFDdT+TS7eMy2MZnZYvj+6KCoc/1/+uk+67l5JEZ09XpRVMw541jXqdUweOdHLgreh
+DJbbkH+a3i+U6AczZmKiV3v1tnMo8dVe1Psieirryj0p6vuFB462PtFgyrlJU3k0vfICs3E6sZB
vZaA2oJDUwmKUicC/H1BtguqFtzE8FqxiQAUYge5agMQHcKVBWlASP55MYpo3wChc5Oz/cDO7RG7
iQuLLlto5DQVwSAhcqOzTMNJW3Ozh6gWdF+n97XZ2LX+p3hqPaZ/CD/3IWjJvx11Z8UrxYB5lhh/
oEXOX3OnDH6x364IOpfLgCHIo4HyKO8Ej/wNHErCpJQ/yFu+nj4g5f2sealP+ZG+aMugW9xkovyN
HghAMGLn/9s0U6jJPguzyfe5U1+I+bP55ffNnowHccKZ+6KXMHbGXG/V0p/ucqbKRI3Xnl0K6w45
1g+B3iD6mnpBzQznjYW74AjhbJ96P+sfAPQFu6a/SBeYdNQ9U1BjkcFBfj+OxWfV3rQZl99aZvgu
uC3oyiIb/DKnv4pCLp+HYD7eI9/g+njZg/wnOq/0eouAEIujo54gExnEkSyNHUR9L3aCKxT8qIMu
JB/KP9jKI+azx+23J5zhFeuppLtO7rqdAPmrY0+53YcMdDvD6B7Sw3Q6LGu+SFvWUT3izkuSWoF2
z8BPn8wjJ11GrJqsKseWoOncxyBg2+DtbjwvZcovnIpN0zXu5dk2x2e0Gyt2oLRO/mOpYemQ5Qkd
kYTVNAbR0orm83LRqzRJTUhzoXS3XbYQGhEA3vvhHNg8sValsOHjluzlhUW/LQoI8nr71B7qHCYk
rlzUUc1v5xVQxYCCEKehEIl4rQhvZeSYdkcPqWGV4+KVI31uZNIJJukFGB3AbbWotJvdy6pt+Xe9
fuV7l6pHji96dDKGeS+yd0pFLxugc0QNI2ABjrngKpyMf0ys4DRvQQWst25vG4IqKqy4ydLhOWsA
xGL5lDjLx8xP8ak4oBuzFI5leEtDeEahP5OSNgiz8k1mVWgJQ7a3T0Mt8XBuD5ofEXqZv755EaXI
bcFQAcqSrZtQk0EObGm/c1B1kfY49W8KfXgI//LxqlhUGpu4Rv+iLiyQwRlYnMdhuI+ycJcYTqwU
fZsXIDUyq+KlrHtxEvzcIvJZig9l7CU5Hq94d1+PSSXhVBAvyS1+B3G5E6ByBOUzhXm7E7+qVViW
gDPTGwd1xPvA/PRqwWwzYe/Jo7oX9PDOilCcncvD8KqzGnRvbhgJmSqJj++axo6SveJF9Kr8h/X9
/lD/Jn6YOrsTyPjS8Trig/GsVGXbHrEpEUSjnfUGiQwZu9vXv+WxwlsHAM3ydW/VCXUu2Z7FDh+0
RbWtUvMlwXmczsMwUNgtXEP2jVUmhrJaQW+tnwHVoPewVdzi4mXzhCb9Gs/V44GgELmMqjo6OGrt
WKgRxAS8NARXvr9iWqh/hNWp+7WgWGzp2QsEod9DZ0iiLPd9gFSw/YxCan1VdFjXuV4F1FDnqhFm
b87lIZRS4JBHwuONOh3yawGNK+T2FzQm6EbnDFrISpjYe4LfwalP3nOXsyodsKMiOdMT25sBbC7N
KnG0X57FpagNKigQFxhgoktD7a/OpJASZeYWTHkEbf86xZtLMQO+Q278J2UAJTd2UflO6qbF8UlT
1+oujKETwkht32Snv8IZWKEx4mMXCEp1X9fsmFVGciwmyy3sU17lLsFm4TuQkGFwT/qf2Ck98fY1
+Nc+Pgp5wzhEYt8jRdcmIcefUe3/e9srakq9WDj2U794iFEcJAhnj4dJkDHoKcsVahrJR/Um7kX0
fz1Y+cBQy76G5OzmZS1FbfGvhDQpnGb6LlJvvcsp4o1+ZQ50eCfB4DjUsNxmtcLIbZ6PXQlG/5gH
/iFpRRf8bkB6pZ2RvxxDDXqZArlYRuCW+hiMqMuC+xWanY3tRkUg1tDtq8Ofoege8cgAEmV1TsWa
+Q2r43h+wwhETTKrRodUx1/zGPz5zthssgO1HSPaaPbMV2C2A0Fi8r1bttvnq/o9E8AULKidmXh2
ogt7Zsl5hviUCH1xQUqqqOcz1QhAT2o9d7avcstxEWApCPI+PJUHiS6//Ht+WXwJhq/Ft6PhPO3x
rmsI59gJlCrgdkyyB33oIUiO6ZPOJM6t9jnveEVL33b8d3UWwyV49fFvo+YTw6BpbEujQw7zrxjX
k7QdlFc02pckvrQo07J9j+o4X9ieXBg1h203lIKsjRfMMVdoDpnw/qJu6DFf3M12co54VyXsg6Ev
aVAhdDqn+j8VixMNEUm/TBvvLu6Fi7HDZKeeHxMHDN4tZzhj2ym86YPgIPdhQj/PrJOIx6/v4EZm
UJE27nl+mIFHUg4PXrzzHj+Bm2AbQUMZnLDz4b5RTwaYbvGgBheitvGVcm4zebiuT/dKkJfFNCsi
6c3xp70xYtUt4I9L5qoELJcN/zhNObigaB33TaHa4sZvqihRxSttWC9v3nt/i/g3V08NSzKMhsEc
p03DgIwTiKckquN7iyI5Im6nu/PRZqfLvpGH2E305pXNsrxia9YYbaDI8sqQM1mcIPzRgua10IEf
2nHByPmQWGtYOW7bzl7LW9nahzsoYjd+cLMuDTS2pE6Qh+PziuJho3V3FqHoPCHY9W4aoGZz4c3K
YCDPCfLY6eK5aYEcXSc5YKFHLChBLU2HGPCL4zZAoifV3wTNBMuCmNEcwG7OU4654HnOrfdUBu7k
x9o0ATstDHAa82mOc1zqfaVfuPxbvBGIu1yw00OIJomT/KscCTT+BjFTvik2MKO+hiOid+R4TuEc
wEeIkZCvEi9wwuC0ZX37PeV5gX0kbirEhyFW9GMwOIbz0ZZKwYJNC/qAmwEHkuglP+JvYRnnTPAC
aw6mcJfdiCBzk7Hmw0MXF6HUGRHLOwUm0ghaUXKMvpzRUeng1AHUzHNtMGSa6hkKanCbba0KZyVa
GuSndOpLJEQlMLzilJldWaNpj6kjZmGOBzepAL0GhBIwLyIOmZbTiKE11ZmrwofPW+drKmQXAg5B
sTvMbOapLGZbjQRiWhSdhtQ7lvsczCCEbJH4xAFwIR5y7pnIZfn/uSipezMXS3qdiAFpJy73W3W5
9WOCmF2ZwIP4qo8fbjY3IPAhSCfMxO9TsZxOwgOMXSUOFIk/DkTGt/fnVe3TNW3IZ9i6zLPfL4vI
1+lC6eYY89hMz9o7XJ8iHfV5z2g+faDlSZxT+SsIS9iadUbVfyBfKfUFMtk/7NFTqQ9HyDpTMnGd
nWEl3iRSjMEAhYHF+YfEUspAGI/do6vMGKe3ZY0E9PizdMCPnelLFadA6nsglliMkZQnPAbHDEU2
lYTdlYZzcSHQAWH1s+lzZcig9meXdgV+K081jwxB2Ekkz/Gbg9mvufRkW6JcVOauYkl1GQtEul+g
dUY7w/YpwMJ20y7cwjidZulMf4sQmK1W6EorA3zbyja+ywqhiQul+6VN2CSrIazCz0HWJPpte240
7Hwoe8qNytxXwulCkqt2O0lr8Po8MZEl2KtX5rxUdYOQGAxE0IIxvFktGEla5QSjZp71kvGfiJmo
XyHJ1J9QAaiB5CnRgIV80AQ/7POHf9Uy7tKGyN5HfagiXIUl8skvWhWuhs9v95GLmcUTm1uPmsIH
4fxgSkX2/U5vApgDLlHsqyH6xacK3L1tEprj9WSIJbfbkETQB8WnhrggnNqnt6SXn4tqCMlNmRMI
1nBAWm1n4BrY2vd5C7jfp9hOn/PLIk3N8S8rhbanM3OW4BgbPwgcbB5s7G530UhxmqOuIX9XaXLe
SNBwLmso6J7f7qADB2g17QyZoD8cAUWcBIfsG5x6T4clr2KA1Mn6K6afkvaKb/WW1nbGho6DBC3m
SKm97dXyQjMwR8PdEgFLuVN07R0/+RDANWwIPa9WflhSU1apfZsrJEe94INvAJGkKlCpqOCBeef7
BP0dWB8IxgwDA8UvYj1hDfUDWHPGrKbOW/SZ5JDNlsnqNgfOaqu0UJgcsUt4WkLtLlB8arFNKCzU
9DgYxIMHEYb1Ze4YAURvkM5USTkPzd4+q+chcY1fFrXAkiX1AkUezJBCWyfC02Nq/NQTcxzrnrYz
JSd0ViiJzISHT5MDtnM2Zw8BVZNFrm27jPyUdb7g9lixSqjvctBaJXvOBpRgmgybelEXw3j6MfiV
XngBytB/nTvBMYHyLZQDMsrhA2mkUrI1BQyPmTDEP1f9rnsJWcgVO9WvhY/Kwd3fRGdhE66UML5/
RnqaZvEFius9ZVB4pKhEit3I85NKud9F57JVZ7qlmIc9uAJ80FVwl6xScnDumyMRZLgzzr4fHdDr
jEzRD8Z4u/qNzsIiFyKSf2J+q/yj8xA7L7XnGN2Qbg2W8qtHJ3Bh6dh0E/5ipSCW8nsWiTcebQTO
cb9D0V1VWFN9cEcjWR/KrGOiAJSKPFOUdCJXQYB3rNKDtd6H3XemsRuY1170rRLNU6f/K+Z8Sbkl
b+J2aXzZf5MEcdZBWc+vtEHxFbZ46EfmDXUVrjb9wP/hBHfwA8sqib+EL1VBugCqdMhUBRR9L7SP
rPNFo2bm3VjdfAFnw7xiHjEmE37uNMWDizNg0+vSKO7pK4z2HjeZvIFPl2Lv0iKyf7m5aWalyBvd
U4oPmqNpcgfggyZ1+fEioXCKwtiOtK1Tyv642Upuq5z3V2g1Q+FsWLnzPvzGMyT8jjO8fF/QT7u/
ScTWzL8amKOB1B69flz8GVc3QJnfOvxCXaEdrpklaEEB+nJF9z22FuTlwGtH8NjPwy10hVLj+7IF
kNAwlVmsrHRkJvsP0exbQka6HSIKft6ycHgeD3eVDl49/fLEmBVEF6D/kUgcCodyU9Y60FCnl0rh
NQ9p4eCiqnGCJlUcB6MYqdxXSRjcMWVJZLpym2eF0z2/dkObwE5NYYtGmKWRO+v1ZQjrmAnD+pkx
DwH0airdrJuaL+GDo3R2QCCDUbRf7FvDYzM+/62JXcmfBl7ltHBH0pRGi8EBatC4FhaXAXDYUYPH
hJyDh3vDGac7p1e6XPywEfTCtFl1gnjkMPnAPOPkvYwMuR4L82ekpSCmvFL8MphyRAEVxwXAgiTp
xOa6Htmel5NT7GqtelZRfUzJleHtiU+kjTDcgWjR+ebqe9imFSmrjlcbvHk3rigfxwlsW+3ATQBo
Z83We00ZcuT+Hm8dDnUFHk3RnQDIo0Zvifm5hRMktrJfylIRIxGds7vJNBfQVDCb6mzxY+INBWUl
lOc4O2V15phDpb7a607VCNIFrSf1SBBjJKd2fy1AwixNVCub81nqRCsb9NGQuaTY6b93i8/+Ffb1
QXEnN8sULvfslTjUdkqUEqUPQ4xz71ZMzQPBQIhkzWs9B1niKRiS14DF0VqYx/pWMxEFCjoGdcUp
nqdHQ3SU14KZ+WlsV9Nc7YYouIbYnWK9zhHMWUjDBpSLT6hDGzFiHvIwAGZuoZx5OXoZt46EU6Eg
4Sg6I9ObEIjNpRKSMV0GMrJ9mMX3r0CHPWrGjWi1crcYDgQu8B0eJzODCH6o+7y1/1ciT/Zk9Ezk
olNi5dmDU496gnuePYvGAnF1n4nqcepLLBSugdZsdpbOUigsSjpYyJN5Reoab2wxcx2DdkZdCyTv
dADqGK4QhA0yigXzgdKdIwONCE4Kyefabyzc4omKzV9e3NztCePWrkRXpZK3vhfx8iMoCgjVWYi9
HrYUl814Ksuu/QrDpqwYZGQRZ3RYr3lGrJTzJaIASQIiXuCGSfl3Mri+4u5O+zVkW4NUkb7XeBkQ
1vPM0H6WEuc0bS/1T3dEzqjnvSzx+b1LZjcdYDRC8BMYCH+2mxW3XWcKHj4gmDrCyYQEaI3vCDJo
/pUHox4YLX4gBstzgqgGdynpzwbASRyX0NVp7GXUXTni5Sg92u4uNrWWjrs6qz3nAf6B09D0wVGY
S+f7el9dYt/BWuZc9et8rOujPkiaU6Ty6WhifsvTmqgqErDquhYUFQpyVKqGr9nsimDNaTLuAQ6r
pS5WZBOsS1c1BjAUbfFWbx7Ev4EDcKgsUSufNLBz5HFqzYQtNPyvM+gNHP6e/4XrsK9crldQgZDL
NAN7bBvZ7YZ+k2IcjknV7lfW2DYToJOfl8SsZpe8HT3nP+WzuxFsqMn8sYXT1jFfDJQtVLQkVf3s
Unw0XAPiBKYAVyQCE8ppfAReMh83SbJkykIm3WJIOZMZChHDUhpD6AvUGikUZ1L/xTXqaw4s5M+Q
HnbTJ8JJg2s1a6Ll7GhUK/f4zC/NnPe2hVpLdOGbtQX+8ZJiz3PNtEOe15RWab3ZE0ojAaQEyu93
PT0KQuiLMPyYpkqOcoGDgdM9TVpfURcSXOoBxNgPhX/eJtdgWxOGW4+9eJEUcO7uehwjUfGYha7b
UjHGvMtisNMZTXUU1v9WutzjrpA13fwnURj1e/ZU/VJ+bsKKpqJ83W3sYPAplGjMkELqSppjldzV
MdCJqn443fofhtDedowuyADBwhzelWgHRXAnE57B1Tqzc8P1jIO2deWKLQGUdb2uAswl/awtmzAK
EfBQGn2EbTmxW6xdm9/f3ZnRvvUOIzBAITDFzYjhNY56ekg6rzX7WuxKaNS0CwhWjwX6HQNi0BUm
AQJ/M1HPcy4KQ9OXO7fE2VeAJC0dBWMcxCA4tXgkpQfDdQolFBMErjfFPGInWZky/xQD0QREhasL
aNeiNfAMFm7onzEtXiGX/LglbxPDIIRvHc3a7hxi1O3NcxvNCix29Qfp5G5kIRAUPOJ/HlZiIfX/
pdxm0SS4P/lOvl1YMt/SHI8zTWIKB6q5CusFySTTZHkcN/bqy2Da+91+NMIfKQg/yIrwdyWoAfIM
TEiuIe224UNC3AgSUfovMLvx0hkSS8dcs1Dbf8T9GMmJ+qBlDuowlY0Dsd/AoGROI5iQ7tL7hFyY
DobzyNQm9RZmJBXs0KbXF0aUwk2rI/9G+mgIFJhP3HEJIRS1qlFwpa3mtZ/V5dHKNj1Sh2MmEQoE
Z4Eh/00i/6w4hIBgPbLKbaJDyXbgCu6MhVi5pEHiH8mRDhKyMqT8IFfDGaLV4hB/Y5HoS3ZX1GM9
AexDsnPkEBGoIiPblQxjgOG/aICwq24tVVG9gEqxE2XqerJMc+LRgamjPMPstg3RV3TnKwFJ74Eb
8/1q4MJ3IyvJGtE9ZOcYcgTpIMVF6Zrvpjad7JcQuh8JrbwTHis/u7jp/6+dB1Ehq4wTUbGCuMMD
WNoWoSmOxEO3PaOIloQ1kAqVCyUMOtvWmZIo4f/j05vuCD2I5VT39THNqeZ6x77Q68w9upBxJamh
y8QZRWPdEf9w3+ocEkju1TKkUTKB9lma2sCG00m7zR+fq11wH58YVgBhmZBHFD18Dww56I51q7kz
DgFdFtYMrG5OHAPQmUZ0xZ+GXJxqcENfdkmGZVNiOOPzzDL2sGK3A9b8IGofSEmRR3qRNCSxz9qh
Gt8fPTDlC70PC/Ka4fBMTkTjgyd8v4uHt03CdzW+mMHkj2I9Mj2tPivhr/W52ihLYaqHEVIgo3eW
/VklzcmBFdwfaZK0IQEqOfHWXqs0SV+ubJfHcXl32xwoZz+LCLzLKqM6Y2vfa9scioWcFNKELROH
J5c6Qq/nN0+xiheRagbJaV6c18tXVq0p5/H5W+KrVo8Rl9QmMqXKyt7LYEB/pYWTIfOnkDjydpzj
Qmr1sc5CzKzuYyiQ5XxdOUJmuNm3F0FoCtxch8sEUtNKvJ0bKGe1XiHDL1IUA5jxRE9S4MqUeS0Z
EPJqW9+JclyIum9Op0wLzN3tTWS3vnt5KJw8QlARVFPE9A6OvJcjfl05CowU8wOJ5gM8IKqOFW/3
FEuG6TunKCLE7bJuS5JR7Cbc22xghd1k53jikEk0+D08L0Lut9WTY2nR4kBEpoVFOefGwtEgl63X
Uq7RhSWo5XyJa8B2K1PF9qWMBbhz8vStgy3YWy4PAj8T+wak50ldI/cbBNzdPgL5tbXqMrG6QCyp
v3S5ilOcCZ5wMjLrsa9ffjfoYraaYuHZE2cx3MSvjMQdkBaRDlkjJWPx8rdXqjXTNrQleZE5wbCl
LM0znZvz+SW5SFF2bf/FcfFXE+jqGdzPKe149PXaPmP7gutuZS6WYFy0qIBBnS6osrq7BPuzRYms
UGVMG7m3KsD4yp65uuZCs1KcYl4kd7N9lmYRN5jOVpiH7Z9Rg7747/HlnyRdT8kskhKrUZ0OT1lE
WGw8XQLsKW2CZmFPIyBUpfF+TTnwawlSMdIFbH+Tty8gLukaqqBiZqzQLPPNCuLO9IrOi6UQFkyX
rSioZVQU9pvoNtwWxZ38UyIg6dDAh5z63CsDnWWm5dzLZbO3PR7VYUcPZ451zOA8Ffwi68AWFUEb
1xK09dfyyYP668QmvMPxQE9Al7WnAppjGYu/48RFwiWzLNFpxOVJePHMKVo6wTQab7y08QKf/s1g
po9iXtwuRtWv2OV2tulU189Uhnq59aaKGb4qIChz3QANOA1mtc/AsVjqTzhX2EIkN2a01lXnXlCn
9uscfRNPx9ryPIA2dNLS4sfyhxJe8ZULBbTrf+rjsKDz3uvgrSLe63s+QWTerpYUb8AvOjzXMg3q
S9BbqOSXvgo+bdhl5ZEcSauqIQgTLPNErzYgFYftsmktXk4N5WhPpnEOZJiz+kC2Xw6Fj4xa9m90
zCJChwG05G3n6xlcG02WgqZC32RXHFT5RK7pQhz8568n9kaDoO8YtaBk7wkAxg+/tBDakJDDn6Mw
NRmVGow1JiTkgiR4QkxGMofVtfls0NUUjIBlpaFZ7wOJgf9lhdTbLVPDqS+muSUECjLDjnssnjnz
ldedtyBzljfMy2/Xc+R+s1p56NRTZ1cBPJSHpymWUKaWI0lB0od7gCsrrMEHDEsnNvxbK/+F47Xl
L0SJlFMeeU5YMg1e6HahvAQPpEOX2Fozlowrbu61eoweAo5dflzU+ALf7NVE6DzeFKqZ7v7vvaza
DacbomvRnRCW38CK/9qE2HejxuxGVITxmCDeUNTDaRt/6uX1vTXqIferzd/sQ2j0KSVLjx3H/OUW
qn6vB2o9fp/PvRz9VCQu5i41QGNufXIlCSIQtp4d0wLYvB6MTdqtGpeAfcu5cVsA3BUFh7tXs0lI
t4GBIw3v9vWCxonYyQg9adZ+x9Lf6oI8zRlkf9Jv7zCfD4eAtFKWeY/KSITHXrAxnwivOaxnzwL6
P43HHvnQ2QVnufErn0TBmAnPVxiQo3tvuq3T0jNAGq2BOdOoR2F5AEkzysq+xlKu2OCDQG/iMnU2
dQTymtPGaM8jEXaKrPAdO1oY+q6UlqpeWgOII64LuCR52R5rfgvs8arJsMGD12rNutQTG/Z7j10M
SeZyz0BEjxDNe5rNqcmerXK9onuihs0cz2aA66sBqB/8t7G5/HmJjCHaoMW0ebvXS+htXLbLE96k
LzrmZ2J5xaj1Cy2QPOej9TukTAUGSY2RlHuASHpnxHqnWBO4lyltpiwrXlOzWs6D7pfUivSHy/HO
VIifVEPeMKG3W2NLuVZkDCZEr078UGdIaBus7YB2mLp0Bvc/vm7VQLw5b3dGeamvN2uYs2Rea+lH
ha8ysaLZCErn6cp7QzjDkj9GWX6hXlkfpoRE2YdKvGHr+WKZ3bT0t8TswKDdfvsyjaylTarINBVs
wW+KMN726IroKfFUPTOzYFXiwT5fppfZ01r7iJ17QdvPcXDt99NVG9jjUPVf21iA34vAgvhRWwNb
5vAsXbXs6Krnr1LlYwboDZJ9zmKRDaI4wlUi/MYnvGBCAHBt+QnPnyfFEdbHj4dDR+56HdcDwG6r
0RAkyEfK6xFwY5W+ufbaykSGgzYntRvDQsNubsWgP77dTuHMYWzBt5sQ+NWCACnu+sfVHw8Uf87g
1vo1m2fWJRaiSWqTy4nr4cUMjOW5ZVfYNrE9AlaSEaBLprCjjZY1PDVkgb0vVVSi5XwON0h4WHEe
W+9ZWNVOKwNAwqYn/LiQJh6JMzLbCCUhEOA2JoJ/QYWGJdeDuBREpZfZInOpknA2+OWUs1TxEODE
qkNCPTTtXnMZavx/7/NGHrAxH2Fym2Ciy42ffR0XaflotB+KFsIDzQ55PwP1lmyyBc6u2VnaGxsP
uqBwIVnjUdaCT/Jw8pN4k7tbWvQ1YNVD9eu3ZJwPFcyd9SDKVw1Vf42TeFPqs7n5+ELUy4JA0cFd
M3VRhCLwMm1Vnt/aJgSHgu8TDg6wd+Ag6FSs0p7XNcH3xt9uo2z78OaWdqjRhs1itFhBEZSTCSs7
eriu/EBh5yDzxozfn5mjRuFgPgJ4bAJeOn0M30UKgC/Uuvg/tDVKhfFrtgYjDIjzLi/hRcV87ssc
xL/xUh+iF9TrsDc7x5y1bvdS42pRBY8b73H/1H0JEkyfkwf8kGyuDTLkCwy6M0eYrc8ZbWAU4Elu
6NtONE2n4pjTo6YoDKb9ifcTxx7HK+vfD057fnpL/2D4cMwQ3iuEkooGtMTX2zh5ramDITdgzMu0
ikPeEudJ8qDEkF0qDJ17uhMEZQW4T6wTmiNB1mLVJjxTTiXSUIJq0qTyYZoSY4NC741qzhAcuOxY
rWkwn21kWxj7NuLrakScFs/naUnGgTRrEPLOS7dkp0yjeD3EZqybW1211HNWANGT0EmR8JmIANUO
RX85jHlWxU/Niptj0G9gqkjle2YozpGcE2VoJg9X5UthskKF5T2Kl0NxepjpGTDRPPlXZU6SPTad
+T+0QGzniVOnaO3InV8YjV82XTbdU3EUSYRIEBInhFy5+pCVEhtyjO/rjIax1nTiw9YVuhTp5hqP
rxA4BNQrlANGOies7fUQd5cbwgDYOVfLUlAo6CRVS+5hhj+J6oKlUbsGI6uPLNeggy2UWdWiKP4e
yjaF0VxgbUvtOJwj7A84318XbLKciULdtML/g1jn59BncuVjepRvhwKOR1G5q2Gp/i0K4bcbrKYf
QbnHZQNh1Ltqe3Z04vDcprFVr8o0tNRDbBFO1TFZNnf7+hCt9Pzuf/Pd1+V7yjDYBEGW9HecvmfL
DWVR6uLgc6HtPZlyRxg8+eo72PGbsYQb+d+NURauReJzICkwytyDg+hJxrceUmDQ49E+ZxPSPS8Q
vasoqU65eemxMDGj5MYgwuA6F+3USF3JT1TF+fgr8I6Q/2pgzdOgLk2jXNUv6Ws2vc9sBvMqDfIZ
0rL+sEZuoaSR+YqTU5i2yaTUFIHlYMJ95nQ2ylS8SUhkjNwIpyUmSiggpA2SzOB7RFBbPwFdf5jo
M16d0atv0fk/mKjXUdHWxUv+hKQRrNGmaOjbuvlubAeyJ/JZ1jEhnfuKFO0lICtjrNBrRUPXSBVC
7sSftG3z0GMR5K4Cs6uuC31fcmyYjGvWJsPSsAmRsCOq8qYO//KkDK8adU+RoPlN3ANLu7aPZ9/o
7+ul/EhOz+2+7juoSHgZcaYx/6Gmr3F0x2+6Hz+CjJqb4p59PzryCJLtwrYp343K8J4vklxUqVaN
X0OhsYZ2cx0USdCi68X2a6yyp6ft723HnrT1VIlZs9AvW/wlk29RBGr7HgWFA2uWz1VJTDKxmqzw
5FoX9kBCdiOJJYttF1R+15vfVL9A7kpsNH/qVVNvAf3C5o9ZphvKnWt9bYnZtX7LyxzkfLg3kBh/
cFVEcjgcDg3yhXhkEV9XktStck7DbHBL5Au6Fo3WysirYYhUtJrvUWn5DS7x+wwGsJeqtDWOa+4F
kaFkUfYVNoceGJu54/Uti7amriBmfcdsr04+qoOFGX5eT3Qsvpzs1hNk0TdgBg+7dPG6L+RyMiu9
cABQiCBK5tbD9rW2MNB890tI4HElylHkGIf8RZMJk0xe1Sr6P7/YhjXXimwKIUeSI53CwhAJVtE2
25Z5mVMcKcOSAokgdkIg5E+t98cbchRgfh7ttjxH9b8AN5li3493zdR/EWtllRUJC38XuWq1Wm47
9LhmpaH12MHjM1uoWCVzZnDRIpSzCU7dOy0xHKsSgQqkUXl401ArvhIb5i7FZIADpUBps5YYwVVD
yY97tXMf97dq/0oB1rCvWPDaWS8vRMko14YKM6wIE2AsZn+h46lY7ZTht0gpK1qcv0kv1XDLltCS
rzBe7u4HuH6hqeuLs1XRNT3wignWYgYoTlfHAIfEojXTZOFYMHuYfy/5o/mA7X+bIKkTg4a3V5qn
8iX6H+7R2ERQP18Bv/Ds8h8cJ11RQ1Rqn+k3iRu+iyiYhuqrvjQSgFRd8d/Ht6wnrxvX0e5NKjhs
efI1jFyDnPezdyKNc2GxoIDaJHSr8WzOUzySG3JB2vDUB+Ay6b6P4HXSjGTITRGglD55YRa63rRJ
Cukju8MzxXSvMmqFnJA5qYbefolojo3zqcrcrSq2huD9Ai09tLGA8S/Ts60o/PxLNcGiwZbOtrWc
FlIanNX8miB5IbxC17CIzHY/Nl1mlgIguWuP1eo4ZHUAzScMXqwdy33T0/aXnjsID1X1EJu8Qeos
gCilk9fUYYFuQOHZE8LkLxsK4oFEj+NPprkKvDd6Pn/svqLY2UWI5d23TYXzDDY1QiPIAvQSdwSP
hn1ZaAycoDFEyA+q/cWbffWelGMWk9/6r3G50uLQDdGBren3ahYpQUXqeVmHln5rR6aQac2l6v17
4Vseq2BQemiJMM30Ec3/fklKsSlQPWKibAP8ug4g5SOkgCUOM5RkE4EtnL80rcAz8XMSoWFaosCK
/aS20eOvMFYE53bBC3I+R8m/IdMcBQvcSbFiKxiyB6qn40VJVpdg2fmQLgjsjTxvt041q/ShisSe
GpAMsB6RAoA5/aJR7FX3z7XtYvIn13zYoJUfASp6zjtKO1alnrqHZWnjD8l4nrZ7LXKtMpYdxtc8
m2/bSGbw4u05IBCUBFuPCrOO7jeo+pfyMS/plJImhpXUdV04O0mejOsKa7z6jT70lOLxj4vuwP6x
JqT4qDb3jwANVye3j3FDXLPEd/q0D9YYBWw3MgLo/lfs9sTYbigJ5n1WCAqw4relny59Ycuiwb61
4pMuy1eqMUXDbo4XYooK1rWznJL8nCh+wJqfoi257zRi/UAjSQTDQJTwbsVXTajMgZL5BzSjbMCQ
SkWNciSVRcTKoLibL5LcbYhU+T44zELLeZ/CDxl+aA1Qu+FVJ6ixfGe/KD0c8D8omxr18jIvPSCW
FZpz8SAFGxeT11l+Edilgs0mzXFBpVjHtpxeZIvG4hTEc78blPHB6mfYllXpLF+Ab4IMZJTKQedB
omb/0M2HYa5/Pf8CVeHZdwWTNrCZWIlHgspcuIg4IYi7JttyMc2L/bdvEH1lTtWc34yHNjsOfnOK
g8KRCq9OVPufgtNQmVPODxY3/kJLu1h6tqhBIATOd343rDDAuKZ7rm37UJIrl37cnp2uUVg2yp2O
VcQxBeoZ32k9FXlRFlwD+AaIEp657xnghGMyTwWCP39qBeK1llS15jobQao3YKGm/NNvBkU2GC7G
5e8WFMZ0gR7/yFFzTwRrPUkv5PnJ6IGIKgBbCbeXVPiTpMnMTOBLmhxhvSj1XXLK9eT2wVpIbc/W
Ho4IpcfMW3WYLh+8AZEIXXIOpfFhF9rgPOVFs4AxVBhPHPgbOiQ9n84gcTz+LAQBRQf96wSBAGM6
pYi/1Bl5wrRa5ot4x0SvVXmcljwHU9fonRBPCClT2Qva1RKQsZ7FsqDjvPxlws0Ws6xR683pdDA/
sVSbvOoi4xoZGJnD7jDigcVNQoyZbbESUD8N7OK5HFzoLoSb89e62K5bNmBQzactlYbe9b9e/Cjm
Ikg8CFsZDepe8xhdsze+PMBmcvYJe3Bx/3f4eimpEWnElfgCysZJQ0xJDQka8yU/BsHi5UFz1mSv
MAesuDoSYTMEbquczb3xvMmdDPN4O4EdbPoi/zELOHaPYDRbiMkAeq4n5RTcmeJ4+Clbyb03P6PE
Pych5ABOylTfALy4cV5G5k5cR9Hxn4y9dc15d/vBaWP0dJheamU1fHPzcI1/xQ6fKH6eISRbSwq0
esutYzKGy9s8R+cRXxkl9NyTU1ZjkahetIOzjokdefFWRODRLnX+WyxE1890qcRWyN52bpC+/DHl
Py1ZnXj/F2iKZCXDd9V2eO9XiIAyuoM32DA74ytjENdG9c5zCwhr0ucZ0TLXFFFMdl5r2spJbR5Z
ewBjqwcPjtuUMKJSA28b1jtgNEJUry3tMiW2n2J/pxBGOL6osyDFZWu2++Wsdtn3aETV5W7NF2wD
uRO14zfrnmKR4h95QoCmgXZOw7Rk8Jgz1q+Km8fEm8O2/hmLj6psVD1YPrkMsBXp66YoeYUwTo/Q
LO+yJe1B7uZu1nApLFFY71T3HxKBrk8OW6clrqBmtLWAGbf+jQWe1IutEUz+lm21LiNNV5qoZKmR
pyONNKK1WfjMmU1I1SGf9Zi3/Jw/fIyeU8mib1mPuAPPH8iGcGvPUk8JUoPGjqBafhbI6L25YyAE
BnZKzKIgq5aTQac7yUSNy5E2oss17t7qGT4xxajsZR0V1zTm9m6IPRwPrAj8hv7gqpxmaDU1ZykB
8MBvR8drRoJofAvQ84eaR69pgPdkt2XvyVz6+02F02oGnWnPTZyVY4kvXJSqLGOWGIJWlWR1tIFi
oQMXgaCkZBUtPy7vk1GcLlYoTxLw9QclEbi9oEr55bhp67SK6+VfwYHJ8gyy5uZKrNOuh+eR2i5o
Yzzns7RZjusZtgOPTXjmZq84habldJtLszcQ4WXj4qtWGZ6gbI5lvkZ28QfJB6MjXVsxu34bp20j
ZRyzy+FRJU0W/ehWzyyDMNnmeKa1Q7izRSfgvmXODIcaGOogq/5oLa56wy0jb4+FfuoRAqLx+Jmj
QZJ4YTCzJA58NqjuFYkvRpBiLBMusz4Wc0ZUyXcxE9Q9su+BNHXpQ8hAf3P6QVkgdh8+ryq/IDIt
1Inlil0+u88a6no9qcsQuENdJ8m0MnkG/raybnjJxERfZt7DTJ4ZjgFy9dJW6UVxVpw+vU8OQII0
IIg7c2gVEkCTvp1zQ9q9DJgcTpgAHcywJY/20pMrL/aLtWvC5WyJqQN0TgNsySSEUkr0Re6m0Duv
XE8k7SL1nP4jgkWn1Hmtm0dB0A9E0k4TLBroKJBTxTHn4YUUSPbe8EvMiZd2Lg1S9tRCBmRvfR2a
4BHZYAvnO+67bQyU+4PVoC+Rkej/5qIGw7tpMvS5KNSgLrY6X+WSzEhG9xGPhLYfAyWplJwbAnGr
xG9etSyVhXsQHDIcbJT4dwnA7bdAzS6hnBTjihDmAed7ju43C0QIqpPX0PaxXfovGNwZBe1bCg1y
01+l8Cm48SUeE/1ZbZAX7fPluj+0Pt9GQ2Pu3noWiAGowpaAmHD6wfrPiKqK3afMX8AFMOuJGd1a
p6wI2QnBOhMtXU2GUmnX9FrEPiKHyDnyHICjQSBHMx9gBlJnRq5JGROJllRQnZdKqvh6QlNZwXRz
mgijGest0BHgxqKVljiIvFX60l6k2pLTxvm/k3WK0Z4Sx6yViZ9FgTBochiJ5nSB6I5qKQjMLMBT
+ct+nYySlrT4qoeeiK9/vq1aDYWbN676gKNHt3mLDtCIU0vYGRCWRBCjlwha+3y54zX5/hAikILq
aPUgIM1vHnuoNWdyo8V4xqBM9GZ6LoJEVZwFN+xyYVpN/5r+HthiGerYeNV0T2iI2ncN1ErKyEW/
aRnNa6lehX/kaNYLgAomR5EqCqUQaGfKjHdvR1A90yqSggKvax2vkE2OQDwzf9vFrMLTy/8LmCWo
mEWuRW55CZ44v0ab6CtCmAzxVj3aRd9r0J9YHFYopjwrIArWYPPRiC4kqlViAxLNRFoFHr5429ei
5t3lEi+CFD9XadROUcPJJoYNCiAoVuEhOl0+FnrjiD2T2BkB1IkXpQ4TF7xQtqwVaiNZHAkcthKT
OQ+Rno0J97H4M8Hf+oYS7ZC3yKrQnTMqR7FEz72SKCyrHcOHaGQgIi+A/uyHqmKrTcIg6w82vQD/
bqRTlXvvFmWnpCDKZUxaATNcUCxTJCnqWZ8yUru4dJJnNY2mIQmQE/mxPHKHoSfQ+iJOFLUXUKe8
6Aa9529McfvX0P+LaoFw3q2nBaaXHecl8D7WqUT2RA6XxFE8Z0B2H6k8iNmjLSIq1/4uX19Qxjf/
c+I8RgkEl0zGQdaFFYoJ/TP+KICpsDtN44jwf7wWvXUYrCmfIvNa2IX6AkZVWmiVvDbaEwY5wCHI
WhBuZYt6Eoq8yU982tJuNC3TDGfyknVYeTduk2bo0IJQZnUFVOp+TKUBwjgSDGTdt+/6JZZ0ptAp
NpUQbVx4xsBD0KZmRvQPRSTXfObErqAUOSUmTkjwsyDN6f389r/vUindl70CX4giAVPNIlWYntAS
YfhOWtPjfENY6iS+nJzFRuG9tgl1kZWzbhYVlf4/iRl3Xd9+FFj9WHbrLNubwW4Id6bXJtmdZo0t
3RiWGVpYmGJ0RjMvh+ygpqJ+725A5GotwSQIxmTe2IcWLihqqlpody7OqnUddhx/wgWJ9XwlOc6f
lwCzPbHvVoZtfVJE5Az3bKP73x+3Zycci7HtMctRKKjC3zwK00pEWmLnA4OPXIsnIQIjA8SrW0Zl
YqtSSkg8kZAEaBWu5rahE8C8juEh11uBDP320hVbzFy7tkG9hWZ1K+/fITxx5ipucRw1gmcpGNTx
KEcTAwla18SXUW0pB5jT7wzS2OBZLk3FJhdwDPtjUm2h5GSa2q4vshSvllRPQlRVw5i+3WfAaPmZ
xiFOVaITN6bzd2yt9M3s8CP3IP3oCPt2kIA4M/oLm2VI0LbQoB3MaG4B5RMxfw3VbG1n7FtwXqcz
sdz4P/C1qKbYcQHgmakP6ZNJiAC05TbforZaLvfnI2c7Ik9pqGZRFVYIZBe8P3wbIDppJeHadGoY
9yLhzwx7KoEeWvWxQws/h5q/fRoqiTDiIKabfo/zPs2Ru7NOywwyMkJRh5qS0ucPqe5oV/SBatr2
8/Ij0QorZ9bPrkJ+gRx6TKzLoWxiCXHXZOMdTQwmMfim7AjDwW8mGQHDhf7feNz0IMpjLD7V4xpB
UFwTvHg/tbqInOxFD459m+pKoTh/ofagchoQhL6hfubiWwlRa+fyzov9/hAn+11cUKyAoavjJ3A/
40AIXvmIqFWnLwYOMhOv4eEIiK1uSWmYQrcPT+kmp3HlNEe98l6dyGyOgZTlU3Hmn8CeLw9ZPa4U
UJbLO2iLvKT8G6nbIl/OPhA8IqWF+dKgyS+P5YRj64DcphNGDZB0yXYBTpHtxDqgedqaOS8GgaRY
CawZF7GhZOqj2MAai1jyk0RShXG8tWLiBL0oJqpZRNvzd+FhaG6fNgXlGguqGPhvq9S9J9UloCht
yc9H27Sz6rl936x68Cloyh2nS02ksKNy5OZCVuwHBt8PXZPB61oStVS69wF+UA1/Sd3saSXzSmql
iT4nOvPlwf7Ybnh3GhBqebyuhMU1qOvntDjc6Odd/h1psGzmI18My41LBPwmC1vH11b0V4p4v7OJ
jDh5Jjw02nKHA64/2Qa/EdCLUIy0qWwpbZ4phoHY6K/9wXgiwysQ4EY9ghJAr3vnupsB0lZlr5o8
uah/u+RDWIxvmu7lc5pyB6BQlo16U/TAcWL/iCHdVhbuQ3n5dKkqRzDfZhcHqnubCWRQ7ZiotbNv
KyHKxiTyhC9RfaDsjNDllZ2aWsgy1p+5Zonk/1mhu7Z9Agx3OegSwmQXvj9r1XoiU7RTSIuwDt0i
t/iZ3stjLuzV+zn9xiJkUMYpYRNB6kZcSN+lK0k3LGSl9aK+Y5bPVaN0q31Cr0d4DOQ0ASHxmUe7
8aPPCHmlbN8IFg3iju0EMVlEenQltS7Ww4J/WDm+9mDjb1LKPleknI6PLG6xmJ7Fq1Ywew7Rd7kf
uyXwrUWx/dC0HadhB3BwQpRBB4COwsyC1G7LtMrZ2KwPzCY8H3q0NlB8kN+kd0w3+IQ8QgtbT810
eqqmVRGijGiWcy6VKZyKyJdxMenhWlzEz/iMCrzwJrysFLFeuncCWuZ9bbl+eLk19KfKo0riHzbw
fGPdKYpOchSm7Jjd5rLCGY199durq0WTyZLT3FbBxA9XjPqs//6/w9BndCYW1usPFCvEkTpSidHb
bdsCL6OuGD8l3lCh5cBeiY4DYLR0Oq/7IYrO3HrmV3mnDyab1pWbzYPiE/pRNDO7WOPbc6Uy0t7A
jGnDElxjKHHSDfzucvOJWWXLMDuS1RDxgUIKWvvxz+IQaBnUQHYyo6oSWkVWDISZxaGMZIyDE6Dd
v30j4pK5wS+x8jL9VZIpE6NsLcYcfzUsAH9Q3MqhgjBlNWSjvp9mc53vnLXoNoMpw81gYNBI1jjf
eGN990YxJkQRpxVsfL8E/CHVXT0Kv9NCSLkD9dKxLhWnyFzozl9etiX+KDsfzfDqCJ0zIOGb/qdG
VsYtWqIN/qEsNyAyWW5NE4rMaTsyayrf52anP/kSWVTsl/3i0ur/PCWOSWSP/5gxsjJXfOMrqQ3M
PoF6kJxURuGkqrDMY1gIBRZ4U4OFaq/10O13tchd7/+sSQ4wlSmB//3vUU2QWJQnB6f7ndKlkguV
hfdq6UCYBvDz86GPqHlUDtNnnq0puC/dZ4SBhBf8yZJaHgYzg0NG32LwQwgnk4Opv8kgz0uqjSUL
lRb1pr1Lmv3r6kO4BTJsoRi+/ph5kuYrb90maqFu9IiXTxdEYZcsMLjBParCjpn7n+enKPUQsS93
38mJiTOO7Cclu/xoUATtKOb7taDQJjaWjODpAXyVicR2WOSMJ74juZWahI+ViOGDvxWRbJ9YfLzR
c5l9YLd4fYbUxFE/2hrmevxAZxHscNJ1OANALUPKm5f16sqdYMIiAhaNgN9W4R4Tku4a8IJq+B2N
WgPt5pkJbP5EEeyMVMhvgm6ZmUDx/4Xj8sVQBH3ME+ebKeh25ZMJ9t8Fw4md+bR+cCTam73WYNAQ
JQ2wB4erLqeJk+WEIwotAc9oN0BvpSd8vQlR+Q9Z8zR8/2m8J3wXQt8bStYTB2EEuAx/iNKFVoZW
oEtJhM3tEm6/pcUmc2QTsjW2NH/fBGO5gjB0qecikUhuTYiTb/GSV/4L2fCi1Oze9s6boCCprI7+
LTIDfjzwtWw8HxrIARpO0jG4zzZH0DTGL0e1euj/ynBTiGxT5+WZaN5jK/wYbl70VH8aGoSToLfw
duty/gMeTJRCbJw+4Y+UXiA0al4YC3TkOT52a7Ur3rllrl2Ux/xYiCrT3Kp7yQN7P4zZMD4rKcqZ
SEIlPkDEXwzG2Z0keDKeWb/8nx8oVnSHGfvHgTW0Qw3sq6/2vCxexu836Ni7341wHESHkk7RQPb1
A7W0ypaaWbUi18NE2t2kXRI1Zi67ItRP9FBBId2YOVnLko1M11+97hT2xXQJPkAS1aVk+Bgic8XQ
rfw6e+iPQN0JhLjZ4TUB/SVsqLw+TZvBn6lGq64/Ghw0Xph7AMAD6iZIxQtexEo2laVUtpqjc2Ag
S6j2BwbNWaH9Pc2EmjdKfZKgDw/MXa/i5CCnf9HDmCaAnW36W9c+fspZXo+eiLJhRlzA75GFUFXM
NALN6/zzWlZezvCN0RQJDcmrD80UceLUjcSquEDyAGsGgkUywuGW7yR0AK1W2v//P5+1yfQqldes
arfBdvoXU/Ju4HnV34lsVHBF+exst+U6z7PQ1yUjdiSHhdxOelcZRP5K48GbaU0NQNHAiiqkQ5jC
r2wLjaGY6jGRRDAqy730f6VT/GHk6205svtoCBuPQC0CYezZZP3zbi8C4YH4wcTaLfrl1ZM1M+E/
quBOD/wIY2FiCNXCkU3eJBPRxYkXAvHiDEfKzfDudj6j21dQPtxIhnew2wkySQzUEbpvWC4oMG2t
rvcotlODqCxVae36FItIaxHD18u79tDZ2WDDiydmgGFvaC1ph6sa6dWsBS8aDMDK8+HQN37vDBw6
s1H6ryvUB4XPyl82W1RNB11zGIFqboIRaHPQxgbzRCqEjSj3/1AIo/TaugLgr4adFpuLzM0T9LuZ
Md3B0w26QLNg/DHAKWxHzboHKP/2ytDRHkYfqmxZGVT/VXZF6hkHsS+evWBNDtCJzqBCX+0TlffK
PvZ1h8X2+lo0cWvuXjW/zOfC37mBFHCW20G/C/m5FG/8BuhSf6aJoNKhBvuGkLsaxzBGtcwSFBIp
kCH5rYehro8GvlCzuhAUfTFsLj7gEz9ix8F27C3v/lFRqgkEW8nMXUJy59pD8nVfbXjrhyS4D87+
XxEvDto7dhsCpmkGVI8rQhp28vvvpZoCjquWjqxw6PnpMidRFSxdwXjXRYroh+ssMgwSWrKgI2fk
rox8DkFaZpHT4UeaTQGLuMQp0QEPPj9tbpg5Qt/r5KAFPmkPp7MuxC0qrOnC69cuyGs1DanQEg6S
B45ub9uLsdhuUR6q7z6lGS7FBpXOIMN0v0bAIrkwmd7lLU4Aik7WTK1CApw3a0azib1VE8upoM0w
430M4nkLAQlpd8Fkrt5IDQIxY9+oYFwn/ySfilhmYMMq0F0uo04Sq34B1quEGfXdjebvZhImPwTL
jvbJ83nse19ZlpjjdfglhL2q+jFSxxj3778ZbSqTMd3kZikpovD5FrJoADStBuh5vlHRg1MJNDlF
oBbM9H+lkRe0AXFuhhnIHYOScxAy0+LjUJwGad6vjQLvQEpSUms69YvRJ4s8NIgCkTL+ose+I3SH
B8tBT99pP0dlNpFsW8wSEAZiUVkJRw9OS3E5kcU8y4GwhyDlDCqAWQWT58257920p90aarEbeUc9
ZJezM9D1BpH0J20V3ESSBilcbXzIEE4Tra2qo75wpTGG/rUEfn8EHfRDE9Hz1YisBCeGrP9M3pkY
VhVqxA0Bxek0LrY0t16Y15GGoIzLhyrRqrWUFJ8EVejF7fezIUOQZBGW96gT02NTwkQ76rIScd8m
5xVrFGUBAVd+pDUB7hVuEv4pk2WsYzZt5jcj4GmH3D6s0DHd5Pmi+kfbuSJxqkxULyFTaAl/rpID
0vcNRJLE6JN6TES5sX0opN9N96aNU5xO3KJj45hu3+o5mDW/Ck9hQmR13HyZp71fDy0yzYUYCs2i
RXtKIzl8ES5+pDcKYfwmCFT8OgIWNawUA7ka1CPcJLlCmNxJN6Kt+hS++O2MpdBLQlAAKvt1wy4q
a3dkknbeUfUsu9cX8wzFaLHBrrN6BwSSes5Zp//2Ean6z2XqVPnfnxpk+t+dKc014BA1DZmrBYcs
K4CYj0S7jigshyTYuSecS2+5eRcHA2krXJ7nJEViLiizqp3ehvjkCL4pTR4oiTekVvoXmYKs8snJ
orRET+KospJ5uUfwcfQxlI4DnHMG1WMi27ymk9yA/+NdB4XfAMKLchOLmopEcwHDVgV8099dTET0
inFJ3Rw2oMqx4C3J2yKzqcl6Df0Vh4OFu7rEB8AeJcPWOTgCgm0Duejrmube9ErTaXHzy3Q2bU1S
udB7prv2q+J6qsjDUYHOiKDk8tsbmNM8TRIgh24QGVn5UFJEf91ndANEUyO5vaRbxJ8j294xZa3w
huAVZG7dK9mBlSkNRHsFHhyESZyJGD2JQO0HKVqm3oujiBbun+OnmJ2lqCkBJeP7eka38T8/Eolj
JhbM4Y5CsrgbvmDxa9bUcbRAwQxXL3gxtxf281AlV3+2SMx2ZOMtJF6LFy4e/gpBeIBla84bQgpS
5pRipR+jLX9WOKy2VxZEvD91Fwrls37weW5Q9DFI1wjxq0w5CnzyjPpzr0Oph0YbJH4P5qq4IbXQ
txdLdg6zp0ZzlzPvS8Qfl7nV4CwuRY1wsUVCUeemtQIVUr5qzQ+XVxkXeMYfgY6C6FjUhNPNavKN
Emu9i1TYYPURGkQF52caJsQbeB4GNdlWeYG+izVgpJMdwfQtYmKalZPxYtdqVEwLq8a/NDNGKBUP
v9akyi6SE/MewyDliCxDPwJKYya32bHDZ3mZpoOShcXoi3WQQcYcAhYxI3w+T/i8hguJ/SVZ8red
6Sctz1wm3tdYNSwIUYzjX+bgJuzokHHRPd+1kMpwTLuCIP1F6rjgxMzkLI2T5xUWOJ3crvoaxjnW
vcaTzFCGeMxkOGzqtu/iHKAIGLbDcTctUalj2K+3dGzIbI9pEQ/6VjeEdIubJfNRb4hO3tDoJiUR
yCkxQvDfSA9xjr5miX3YqVQuBQv6M01GuQC/xG1i27drK8GXcO3yyr/tQb3wYqUfTEGGeGQBgLde
muVzMiW0gwFRvgPz4F81yjY2MYI+3BNcY9Nj35Rb6a/FflBYf1YeUv+J5Z54yqPMZYPBQ6u1RJPZ
U2j5o8tqwjW/26Yb7PZuxMW0k6Qd7bthQD33klXPHGG/jO4QnKzTZeI0fzK5M/0bsiP3K7Q8j/GJ
CiyEGQkrZ/hULlt84lX0O3ca4029nsQK3A0PzJf3qS5ge9Aa/1ztx/J4ypKGuOTk4BRuFWW5FUFD
o9vkVjN6pzvw2VzTAVljWpFHH2+uDVmpWMkWtUgO6PM/1qNe+adkUAyP9cYkAYcMI1Dqj8H9YmZa
aCJWUX8uN1ImTxpROlwKCJ/y2tjpdrgGZh3Nxa0ieDL0nSDaO/LqDH0UwrsT38GtCDA4S/uyi+tn
Tr0cvfCgecs4fbQ2ay392AroTSmbU8PRULWsXCwClAqyTfNinYHA531JTVr2HGKQObTtW68XmZ3/
fUWa9REZQByfwvNPKfpwsWK+HfZxdbqJVkLyjiNUFuABocl01/eYtJoKS7ROJ5ObzdIn8EDnzL8T
W58/wTJgWXYOVDGLKERrcs2FpQuPZ9/2VVIyAB44ISbxDKE70kNdwE+ux6fxW/7MMAZOB+uh6bBE
nqd1rwOjBWZG8a+UrXLQcg0ObFeNM27CHX88cSi+LnBTdlL7Tz09Ptqi6HFylmhO5x/JO/DnKAu/
NZAZ0cpBcFfMbm5cgd4U1maZ2uNdj1nqgeKSk9ImG13Fhmf362M1hdTZQfOgqHUFMllicrVu9Yyu
/7e8NtaxH7QBHfTvlMVr0s6eOwUmh5VkK6pDbEYQB30s+wceZU7xDg6+M3KkhetSC+GQdp4xWddZ
mN8s7yga5b7HCl+spA2Bupp219iiDsJtNTstAcdWxHihf07tPUwRwLQJw7OjUb1D+E7N55JiIBZ/
kEqCn9KihWlXGgDm746b0oJfBh+OOFNSI6EO2WiPKCG8ixSie6V7gZbiLcwC7N7J7WWKpBsXajjq
sJ1vequGG10Punx+hjTuV4H59nnMKoia8INoL5udziOhiQi8YX+HFQzTqFD2CEYMdc0LIXQ+kM33
cMp1cMO+6Mi2gpVKstUk5/nm+R9yRoJWU3bZjFxvk9zHzcgUJsFxCBB4YoQuvP6U5b0tcVN3SLV0
ntyQ2HhQ7xeDZrEd+VubG22nT//pe4aeA+yKQEGaQIX1vCiIBoOpwV4t30DC6jzG7r3WWkM8OPPQ
BweB+4Easisxp0O/NDdLwoZzTmPTciPC+y2Ew1F3OewzFq+GxGXfszHw9hliKetCSaUodB5Mp/1R
gNK2p9sAKzyAYqsM9/VS/2TIUAmlPxn65bUtxn930pauV3Iir0ibpTbMHr17hXM8ibkqk3lexnNi
zX1RGHAwkZtNtoqYT3vs4Ns3raE0lIvT0uGOB9MdRt3lfWrYYnEBJ92xoyIC1f5l3mcZ9pXuWHID
tSz7LAXBa2jE/nnrI2uVgtBuauCbGyvrl4WC/8oU83A/J16w40663HzFnLZwLKbVjzRLhcUzIArf
RFYTezuj5yPqs6hCOerOIUntFFqFpnWUQj2ahf6QpSQUD5GkkpL4pRqbEXHiH/j5HJJiJZurHjs8
euzTX7sri1BIKRm2biSpl4sAQzEnbM2vBFs3HDufXf9IzY5cOFgxXFXDYndDYU5cYBI8+UA42mR6
kx7lZ5PADU6Xwp7tOvOO7btmNanxa+sWsssmiYZ/nMhTgbDymmtZxGk3BhpPnYunWUAq4A35sE4a
4cdPynzzKVmi85tA9spVK43DOjuKP5cGxxN2ZM7VpZRgt2PvC/LpqznL076R+RLFbJpkZnhj+MYQ
0IFfz4hvsnac3XYE8icnQDPKDfpLnGlDx/etNDthvU7cJzDiKNMzr3tNHHqCCRdGbv+gYTE6tVlO
GnJciVCKgWss8hTIjbbQ4I+JHs2B4o15g9AUXQ7m3HAIdWW3ZG8Vxuqs6HLQXAszQqx3WLztJ1b9
uyYFG8pIHQHkIb0tgCXcI4HZggjh60mSEz45C9JBWyjvTXAutFw+m1c+3dJMOqidZVXVY2iQ0NGn
ZFUWCMy7oundIePvSCpfc3wueP8DsoS/xm5VlaF/EzMmziemxiFEpq8+wDjX5D0Iny7PZA3/H8dR
XUlnVeY2yjeEo7RN35fk4wLWx1HQzg6OJVIRkKxASwHFlCNlGJdwwY9m1GTYuCG/JWUSEq43T9ft
upNap9iJUADBLF57jS6M0F6T+8lE6OqVwWzUPZ6hj+5LTAIOjyG/v4Np6exXcKIhGP3chkUzYOp4
DZBm+BLbFWt83zVfeEVzM7orZO3zgiW2v1aHpUcn2XRWoJnK/1LtCZ/kuHDWov7CPJAtMWqoWi46
F9dRAEQ+XYehCjpx1RTk3fYcj46XnwamBcQtFhEPz69CUgifVVP14e6P3pwpJCr99qrw0s9w6+Gy
F1dd/hzBbOEi4x1+MndTuSFwKA81rD9oR8kW+rMCDRx5n8AC8UFUBazdBebfEOrQ6zbB7ug97y8G
qyPrgJkk55X4fjySwOeqb9V+5kAw8GqTRRD49HBBt3VVuCDXlz9DWuZGIEUGBpv3FF3w8/4tz2U/
M9UsPuSX9j1jqjDxc/UFAXsY9Ww3u7se/YTr+3ino+xuptG+9/00zjjZCIpE5TTgXPIA62Yx7JVU
s64RXX5YukOd7MOshxdP9o1S7MLLygR+ICiHbX9sx+zUsPnud2Dh+xBhb+PAk2C9mjxZER9CGoNS
z6+chEoj0A949IorLYVRkl7aYBFydBIEY64AVx0gVW0zNtOwpwfbmGLsCSXs5uARBUdMNJg3UBrJ
zIx1zPiz1CBYIX7Ythm2zLpPfQHZFNorJDR6gwbNehNHU4cicseiS47nZe5/4bGH82UhuqotMqms
KCdSR4DD01QvNRpj9y6FCD2k4a+rLt/5gCI4HoZC7/wsQL9WT422wE2I3ylYexbSLvS0pGHxCH/j
Ybua2PwEAbRMFmxx2X+E9Qdt4sZbGCYPqm8qpOHNJa0eE7/AIFBYTFJQel1FRGJXljG7vWwdZKkh
E3E5EPPHZL/DXDmFZ6DlduWkizTSirRsL2Dde2pbqBOlWmbSki/VJA7GpmN1KdIRwrilPjMSa70D
3KJcVwxuddO+TULwjlq4DQiusVC8uSHCv/sLZ2I5R8IJqdtjjjleIISSbld03f79mZErrNqVFNdK
E2uVCfq8g184sTDyiPiQ+QXPG2X3fZCMFhhQ7bWLeCkw87k3SIN90OxWVnhC2zLChqmNmsAg+nUW
CiyE/Dup5WnvDCijBmcXjxIVS1OgKbxrXlcbQvZ0gsd7QcWP7dK/vzYYxRCDHkLuWUr85MNjIqXt
x/z5grBjKZNeETNXmpd3ksx9vbcgE6qEqNFJI9nO+a3VRa/bYgaVhNyTjQ7dO8Nc2Ajk9sfeRFhF
yLedMbp1tJRsxo8zUOTMid6af0h1W2ndjHXZXH6dJyRtf1QArqzGKp9KmERsuriZDKmYy24QJ+XN
oJkzmPE3xRX2ugxTvpcfT4a7JYfthSQkJLEWj9+NCoO7C7R98cyCHX0dEFO8cBwVbxYD+Jl9vuHi
vDWL46WN/eMJaKKikvHCDrXio2OHzgiDAapgfseCb9Jg+gknuMHsgZeq/TplMkoyKqKO2mLI1c5+
SbUK/RBZw8nMjEkQExtQOQkbiPvOLLQHonpmbZfs6ofOyjDQJ4p/E27oI3kzKGBCUqW4Z7wE2gqs
+PLtExA/KiuQsnYjaMAJcGVfpQFq6spgBaq/HavGDedIL1JDnCKZmPU/of3OFG7+RXP0+HcbV+7j
dw7a2W4UONW57Z2sr5zvZtP3ttVy93y8jdeKIYryCOP9FVVKZ0o0M/lNkOe6ZRB83toMt50XmjQh
UdE14r/yGjFp8MuPSZfFg7Txdr9j3+/60PuGnTgZA1hc+9KuvyNSnHrtCFDc6HO5L+WKLf4QBU7L
2dH3F+P8DEpjlOqgWeqeJU3VqqwajZiwc2ATR0rc0WntiiGSZE2qNyKNtwK+OcyhTmD2riAYCP64
Wt4K9Kot1cLcqE46rfz1UjKpZv4kwm2jln/oHfo/VvCzJ0IggOcY1yh8FQae5RJ7QZlXjGAw6W55
WUORQfddOHJ7irLPUpUQv4hRv0+zZPbJlFp1ePg9C2kviYSGwFD6jKdFOvKZNIUmSPA64mjERGLp
Ha3j306gUWYSU8VbBVpQcuaQnuQtrbtV3s0veVys2McfMH33ysimLVQXtiNucLVM7CIpUVcZiNYI
czqeaGFEdgBE9XO9QoeMqZ4IoN17e52IFz2u53zFqVksfd+d1CG4bJuViwd42YxkabtUQNg/BI/j
5tVgWu8BDj88Q07BuIQycsI3qkpyuEMuV89xLqgSNNETv/ikO9Khxc65EY5PrOVltUXE0ogFtLJM
XDY5rkbWCiAV6nuk/nEkIzfJzc9ua7aF7HN2Cj+oa8RLoB7d5Z6G31LWUYhK4PAd4yfhndWPVHWA
RvSh4ysQP2Vj4H+wDggTf8fUDHyINFNCS+IIUGKhqZGcibVS/0nrv0Ntk/G+OnXy7wH1CWBMukoD
SJ6JdZ4P6zt/3XxVzVA5ZTBEPFQcL9S6hTP8E+RWju5YLwLEKGQkiDNrTR/CdYhnTk3dyQNU3fFs
YZd3DlsW+vUcT0oWJfw+ECm37eB5CRxcsq7xLKzTN98ZlysSCSNo1V936EuSoJUXdeydbEDkBveR
HYa/oHr8w+okjmuwX+kLj7lLDWt1WHMx+0sEfjR9YLECV6BcO5bpdmsFrBnLQ/krAYfif9mp4YCW
Qh1ElAjkPeRvhzwjoCO5hMoy9KDCO8XlmNgyeRS3TJ9KsFLnWF5cmNEAHy23lagDctjGDsfR+8Zt
36DwPEjEpPEF2scCGfo0ecpFyv4jYRa4eLE++9lGvj9tIaAnXY1dRihh64U2FbnzOJWIG/Emnz63
akhaA5e/Aw2DhMuW5wpHP58wlS4me4oiipmOxs85scoF2tkBRxuF9349L71taC085cD3m2L4HW85
UrH/fuIRAq8dA6HyY4DjzURpN/EtGOK1hMU6aYKQ198FGUL8mJ+PNYfVz6dD0NwJFWwkvjYxFAIY
zj4M896mXy5lPFOpCPUgGJQJkrAW7XfU5bmVGUJ6LZIbBgu8GmckIz6DOJo2CHHmqPGz5HgOY0Jq
aW08OIh/xEqzTIIck7j/l+HsujWEpAm/bpv6K+aoXDVVsVN4Wd/XSHnbH1U2CWcKtdEVK+Sjdba/
q1Q9/eh57VFfWYynqwyiQxUm1IbEMsAelx3RBEKS1J+YmX3xTPkhbBR1z4DS0DBlnZmgNIJUaMiW
OMKH+ARgTaRffbkEznM1Bd5dhCP8aXPucsDy8w+omAyZ8pzl7dFaRDHzyp40oTyCqwGamns0gJEV
qyiPzvJVkICpOVhw3rSFdd39Goqgtg9+JgSXr+k/TmHfkL/Xd3v0JP+LFBS6mnD5UoXM5re6HpVL
ygRyiiv15guDuFzuhSM/DV+gmflpdHxDk1B1sYosY5HFfbN6Dt4P+8OwIWB+dXtEibhBKwm2f0Bp
xwNzSCUPkg8j9X+au6nev53ZTLol3IjI8zPCmhnYr57GjsiDTLvn7GMSIeZkTxgrPg5lLm0/Y3WO
mlXrc0jFg4u8NluSUqzZkmW8vYwXJZaUl8CvqKe+46WGouMUAESaODrNqpVfU/RNWaRVwu2L+MOb
KvkiayIk8nr08/jwRm/YTC72Swz2n94rpAp7rG5BAioQE12Bpc3MQh7f3n5ZO/6dxaF5wJfQx/Db
n4o4VHJSNOIbG1HVUW2iEmZUz7llrI4Fc7+jsC2GNMINPHJsFbvP3H/C9vFlKKY4rcnTRVob4+UR
/MqMHqO2pJ44+HB6LC4dySO4c2IYF9ezFfriTQlQXdtpV2e/cVjgZkn/z6NPuNqXuQYhXYYnKgVA
BmEZnsStu0Z+hq9Wj+wOWP+pfzOzzoVGIePyTRz+KuYF/JL/5vzLWFHONR0gvoyEAqTQm0pUk2jW
cwa9gyXh4P0XEoVhMMaBVliHQ34Y85LffxWKqDutE9RmYyzXrK1xtYWuXGIZhjMJ6pMzYqtfs8Xc
ZSJh4xjnOX5DgLj6nDv3Iynu0GheHwuopnIHYuEKicOGZXYvn6QO/2aD2HSduveqbOzvttIgqvoi
Yox1xapGdtb3RCdlCFC+JB3VA4BYIp6UvJztK47XkBzvdjcgEi12Y7NS6Z5y62srH+hcXDDjeqhj
izB/KzvSb8XabqAZOWdtrzu5LAJRqKMTrKEG+ji/EobziP8E+NIsGbjslc5Z0qiKdaJpmxEHOG0E
wEcK/TTB9XwdzuapAJfqiDluwyxFMjMf3KOT5VTkzbhkVax3Zibxslp/1E7Nhxq2fnLCGC3xtrAl
/LEr0mlWil2rGFvPqDW9/WIDxaKcSqUPPKf2U5jt1Yf889jbcypmsQQnKWpMYOi9GPquC4hYI4uC
iTGCaBFLREnSfZR9zQOI8AfBReVpx8nCXlox5a3HyrhpWwgL5DzUxGnoa26E/gjwuswq5mdRbJNw
QHOVMN5Vy5rPv1t72bUxbJPK4o6KgKsQNfyFb3gAFd9mrVUzLQqOvtT/mpX/S1Q70mxnw8uDA6uA
NWtJX+uEox82+wakLEqQR+a8mg0VhfzDY0pzuYDcPf6Jv8lON1RFbIb+IqkB3T00YwZBoccyI7jF
ZIyh0Z2o82+jLxXDRLKW1VoQ1jyXQb0DN5FGNi0py7SeTRl5HGhPWxOvxEFgYRhun7MX6F1AFzcI
RMJVy6xD8s6bUfS5XHKnt/sTk/EQH6AeS+awMLiTL1lS8UCKmGyShgFVYVjIVAVN4Y3ezZHcHEd6
b2saKoV0bPgH/OzaGhDIWlFdMIff7h2PradCfPrCMZm+qbaPi0kKWletrTYdj0Bp9U2hqIe3gYT9
3BkhPYKhQJ5NeqaWmXwSfqoW7rR8hd6a4dTDhgfP7LTY9Y/cV0Pd/9aOHqJuZv10Ql+8MK4YduUh
P17MTNfgA671ZF2ohnXl2LpBnOmd9VXqCxA5PH+GxS6W7Q2RXtyuQg8TA3grW238roTeSjEEgZNv
Y3TtYDMqt72O3XkXRoTY0mkpNx9jFUKDLNTb9HeeRxIPfi4AVOA1ot/qYnUce9G2TyW0MWa4Dnaf
KfQlkHVVTQZsHCHdBsn29BpLMT/fIOdMO43XZTi9lfvWKEljImQs4Ffa/XDeLtSl0r3NcZlE4HRf
k7P4MmIGg1UbCG9kZcmrWUOYPvpZIKnNVmVCQoS89Q2SzYBZmZ5zeeoUtjVsvhKHb08yqK1gJvTr
YM+7hru8ML0RZXYVOawQnfOLBbwzFB1GN6Z6yluKALZw1lRS5HLCpJUeCVpDgEWVnLVbIoM25hZm
v5w59wmSIMWYqLERUTQYhK1sAffS1dllmCh35TLf+l395pogzzpZpAWWnaL61clquqal+DqIx5LN
ILH58pp96sM5aRkrtQjt4tQXAYJaKNxIzCgR+NAuxx6IJ4LuzJVrCLNn3C+2Tz8SgaJu7L3j3cee
zC6DdVcIS4ox1xg4gwrQaMlm1d1dysk6O6S8CHDebKRbKtC8eUbgj39Eg6LHrs4xyEgtOd0YdhVD
8A7zGHEcxokEnERH9AGvkfEzi+iOEBEZcUffXDZv9Xf4n9bzWrXSQXKsEd0JUHYyM2QkambGkjOQ
PDH6IXLnUjNkO4Ks61OxRAI8UY2I5duBppu7RkV04B74O++JJZuE5HYrBNUWjyEe8Q9Anx/pTRkT
jIMxLWH41582TGrTb7I7iVWQrVvts9YB7LHra1VojcO+myYHW81jffQWXthBZYSU8RG2Xp5g7QwY
NM0we8zSh0qkxd92REKx4taVJbhlDGO1lnAGoovSnYmH3r9hyMq6b14GjW8UMBMYczHlcttkrFuG
C4Zs4RoO7lf2YEACKQyWMu/KB1rX6rchkJ/jWgyr9QbQjlptzCIa5I/869YGdflleigN36xVBshL
kV5x4LTJSyC7TPHQwGdlmwCFLuCn6tFGPuInACG4Sv3+z5fGCJUv39625coNj7jDxaC9hawx9nfm
ur3OuRkfpfr59ii/ZtNvIQPF05BZIIsS83QZfIJLPHbLutIi6XkJ8Tge9w0TAOs5tx+Cl95o9O83
cdEeeZkJrARdl+3x8sAaSDP2JOitBgg8oxZYklH69zDGlpDbzFMpsTy0PJ7G6W1pva9d/vaYEddp
mCjIvQ11WyXDoTUsMk9qE++IwfD0X4tCfnMuzkFcBiRmx34dSnd480b+nQSZkmErYuDwdV6oGG/N
UNrZo5tWGvpWCq8ApuHibilb/x/YJlqjDYvGMCG5XayYe9+zFJD9d/LfL4wbsuwLQuykoMPBprBq
dk3kTGUijLFieY9VjHFhs6gwamJZdMPt39Hholc1YxsZMxb9QNqYu0f3oPcOgeQYjIyhfT46/mnn
k6t5+RrpOq49raUDolv2ygGiR98wUz8QF43vANjuBqy0yOpsuQgYyBpviVW1/4f4lux1V5ZFP+ZB
WThV20pm5lLbgRXgfvpkApxKxD2YcxQfa3dr0VMEjI6X9Ne0rhEIa00qPjTISUSDIYDLXLT2qeBq
9kp0U1AgCWZUVemniI4VTLBJG0kyQ3ziIeYT+fTuUddpT50LYQgAtZZ8DGc6TDoXdIESQ/RD4wk1
pq+VQOl1dUl44qmIC/fLajk7A5jBOPET/3M3L3slJ5jiQtBE102isfKgXYYM6AqbITKlha+g6ryy
EgLVw8jeCxyibLfHZo5m+lhQMyIehFkkZ32c3k9JgSQjdUc/blM0jkhIIxEEcFJ7Gj66DKBuZHsZ
/ycT7fZvTb8inmD5VNtYQSnDDxwgj16GwsbVYFlSZuP+WlK/VKbOijAb4kow2bKTtpXUcsOtLMFp
DTOWlWgpAuxJYIUFSb41W88YKZPl0j7gFzBD78P/2p5hiXpZ1tm00E/bQGsEp3Im/9/P/67Vb5ya
Sp8kvhyKVOkR8vvH5KpJUdQ5G2+V5OIuSiHSoL4sfGjIBx/ePS3zHLh4MV2mkzmj25glXEoAaXOG
mlzvUlN4ERcLqkhrah/jAoHNXJBjXPPuitPwtzHRch6m86NM+UK5Htt7Bi30Q7O7W6FNodZd/RBd
wTbWSUzcQ1OfKq465OJhw7wFgfH18O3bneXW22Iwr/MuQy6ynfaH+tOr8BenkxsXTlydQEF4uLUV
PoCL4IEFPimD2MByfE7dZZnd6UZ045VMYS2VNHmOwb1lNp9QcPWjX7YeSTXL0O7dV/fo8zNebpt/
oSbcgOZE9mRVt18tI3A5ONPj82PDoKgKPHsu7CjN8M88C0pTTxP0jT+fyLyFv1Sjf20yslBrtv9V
9DNT7qzrGcHUbwxphq3Bk6xCLa9Acw+TV+FVbfWRQX44dim8kWoQpCffjFoBQcK6Vcn5LYwA3go2
k5XMu9Ts8YzV30b3FPT0nynO4kyKq4gLdjnfw6nrudAoZUaOND1PHV/VKuklAAH731ucWIIyVNO3
aNvuN+JBcvhpYAupAFvPpmFL3GUjEcpOmWU++5xWemPY9EPHC4uPKx4D2NG/iVxpWF5zKIDhLivF
RTmeScNwCBOQqVKceYuJdymYJMEuLBnP+IgNStNpH7aWU85h6D4HB7WRAg/dNCO2yreHxXu+ms3T
nFvOziGcquuI2hPc8BexJZidoTXT5fuidY0V9PVwMYUL2S6cVlX5cSGcdIvzD8GjjBvkcjVu3zVN
TB6Z8oTGkT3cJNGygS/JpDMCaNVcfQs+p83I6c3Z4zachPgwWWtOuKFKUqVUn97ZpukHVqHvtTPN
eSajAVIVlhWrjV79rnGy7zN1BiVIoV3XgdFOJISL80MmxpY48sfN6IUz9okStN/dK4YlesK10xaq
mWJWcVBrzw37gBcsFPmDgHYXKhfXkcrcD21hiNsppIaDwQYVP7uK+G1rclYQFbwHVbH9Twx0Zq2L
4MwKVg0lPw0lPuW/GU554ExnDI+ZVMBl+qGtlkmdidpVBelKunxjitVrDRi+oXOTIvW8v/OboKQ3
HK3hx3xNS8Io9KYDFxlIHYaUlPwOqmVZCSQarbT+G1yoche8Y31ZJmKZ4xJ2UhY4lNb/rRlpqv3o
7JJjkKAX7yc3+dhPV3Jb3m2R/fBgZf7nzXQEF8ubVNv05h+j1vFfXf13ODsbxC0TYkH7C2fEyCAe
u7uULFeRxk9DvF2x/D2G9FJlR6Xwrq+c89NoLDHD7d9MMM9LimVW6EJ0LwUi8ucWK8fEfoE5M8NU
cTfn0YFwrqE3ryyD47HeUNs0tO5PdVAQ6vdoE15wlAciOEBfj/UdVIMgHQskVPXFEmDQdbKmXjrp
30lzD0bsEnT0s7Os/ttGdO5dxP1BaaxD9937ZQrG98PtQrNiPFKbS2geBoK+WCbiM7DUo53BZwR4
dK+qF44tYzapX021BA/6j3A3kpguwv3n+0cHTwtGco48jj7u8oOAUJAzM5I9xhDXNBkzQF5u9CPm
601eb35kh/75Ke5LYIcB9wqASHNSzF0I+KK+aB8dCm+f4h8y16owxSI9EQD8MGbFCl3w7u3htm9f
GRcdsIrNMWhxiUZz0j2nZ/W2OYpt3uJcV9I/yVtTV9paDEbNWBMffk9dK7Ux8jB3GEruWF8f+0U/
uk+Oc9hALaCdLv1oFYxpbYDxW0dDpwtWiyj7q/kfce/vG7NENHE1h8SuLuPMzJLwfHKqqszKqoJy
G9X2pLyr+yi3xX56/BBfA3oHHczfSd2GmdF4CPh6QzupI4qimfgaTshBHlsMTC+8/FbEQrWop+ay
ydSVW53Is1FBWDlVS2JGOZOd0DD636fFm6Dfviq82HaH1No76/ULu79MeG3PpXgPs+hPd9urx4l/
pFu12w/8GxRD2r+MUo/KzDs8AJ9eSfDfLH/hgb9eAeMicLNQynNm06tC/9hKM67gIDy9ECCDyYM6
4eSIC+GGMwE9/Rx59ChWcgHmMOAMrlmrA0HGQvu31Hv2BpIw4/MaU63XdJ3P0USqBlgXifhCc6zY
/wi466poW4gDI8OvuaZp1dCkRSJ2LFW96nouG7SOratcSRTvRxOwRBnAUvNDEPffSwrr4Nf6m54J
qtpb3c+jwRlJWNluc3UYuNYNnFF0LgvqiOtsjvWclSqixLoCGue3xpWR43qlrjmJgVhanSwspHyw
I078JyGlo7NQnc6Ht7TD3yp9WNz6kv16L5OfGsUlCy7s1oxucUkalFpTbNkjTefAR/eXN6MOrg91
6EBeK68JOY8o0/E3Rd7s6IUsNTgY6X/ARJKl5jiNCbrLeR3/in0b94Qbyn4G/WCh7h3crBGJLwHX
9PM5WT5WoZaKOknuZDe2nFZ6GN7Baa++B0hYrUCYzBVTxDKpF3tp4MwtAmBk5ILAwKV4ULu3j97v
xZ/KLhTybGBhg8nSzXtG2UHL96SBzI9pD5n5hMu6i6GBIz6QSE3vyCgSCHyMGXRpTEKuybBSQL1Y
P2vVAI0cL86LSTIC86o9GtRQAEDYYOtMPFsq44VYSgdtqtGmslBLzGN8XbcfKtIkHgFhzkfVBi1J
8Rf8u7dTUZm+ueXMU1Z1AaHSVQeaFgeIAH30IdC5DXQ1Z/7lIiHYPqOJ36WsV//r2/sukD+EyEQX
G4Envs9ua0G+WRfIMS/n0klv9CDjsy2mmjVbpv7cEY+BKT31d2b3UQVxEcEx9z5mL1z5JgkJ5UeW
OSirB3U2C0KM4NxZAy8UlKQ9vJOXrDvXxr2YVuztW3I1A9AWLN7p0GrproU/hhIC4ywJM2mxD7sO
3O6kd+uffTFR/Ih7PXuHCMc8LrZlCQdYLKlr7WTt4D5TWiX2eVfPYCSiDt83y3NoDq1RsinZtHWb
EimfZC8CjZj0C9NLDhwYB2MQAvo2RFuCMd47j0BKlwRillXe9ATUBEOgKom1bqjfLD2uFTzOTAGJ
Rdpm01pR8vouDdlJRmSBanfakQKPXk9Z3sWEi/dHyKf9E4eonIt5pe377FFOhi+PsWa0JYPvBZ+L
+/FapnUeocLowFo+qMxhLleFoUiFwSrs5V8hnA9qMpERco0ppf+PRu0cptkcT8DIdqPhn+HDJ59D
EpYYTnRUSR4j+TjLoyma/6mBd+a7lmzoM2OZj/Y7vV5oA16Txi6OjXaNV2pCWP0s3uP3CQ2JJMzs
pcfcRxeIybiHQZDfN20tp+ju4rWM5s4BY4HF3ERG5xhRspW2Iw+PEwpuBzl/qjKBGCKB/i9P31la
6Shq43neP2IxNs6s5gZDlFLwYaMLmNRbR5QM+iBKkQT0payoqe3fcBk9naYl1sGdJzrGRPR2oAPW
81Cws0sFDgoTmUBHI6JIh8GaTn+MAmriX06GTvExcmPJxz7vXi38ulEmKqLtNWnip2HY3T4NPTEr
3+pnXwl8gYb1nOh7GGuaeA0F2aX81jE03EggYzjVxKnZHbgd9zXw4jZenBIHj0HLNgbUZFlJiKMg
1RBTCLLtQ5ta3DLmFpE9l0j76xJ9UHsObhRfVLvUerEI8Utu4j6L0KX4ZCLkeX5dvIL183919y+m
6CoWKbV3erjqsFHoGOjYdvQrkefUZ7nGeueYt5iT/4/E1sOHH2DOAFiAiYBwsrLbI5HnkY2+jYIY
Yjrm/Ns2VCQk9QBWql0xKcN58oIVmgw8/Y5Yv1FSi3diQqOYGK06wCHRBao9bEM2kfkttvqAChR/
5/O0SyyRrUhiJFZp4LvnSn8DVxE5Fno1kDrhucMSagOp6keZ074qLc5juIKWc1s4FZKxmtLBOJjH
32ZpYh54y2FTDCklNsgwLKAMIcf4Tvc31UGOBtf/GZSU96M5reqzlElu3MtyGUXAvULJ+afU7yBg
DcwPJzPiqft/eJez5EXYEdoj9vHUlNanD1/eJCUHG7f4LNIg9b57PXB9FV45KcRNZq7f3OI2STMl
7/614doZCMohLelBq71lEB2Y4B3fknKxyTom7xyKCy4iSOkbWYun3x0WRLTYHSrC52sHk4FRwHKD
l85DbAvkbNRfU2Jf3RUWZDrlybIreJNtdHzVPcny+VwoTTWQunmen0vz8PuefwvNu1ak6PZCwmw7
5Sz5XRbpVA/m0SmdYQm203iM7j5Z9ReIZ1+usgr+indEhUlup2NPWxMGpe1mmgfQinw/i7qpVqh/
6YZcytHEUITKkNF3MuiHlbTr2ndBNRnnAY9JfSGGrNKJZq0f55e6ojPiy++KA81M4sX67ZVbzX8L
Gz8oQUT3vTH1EuT4DCl9MoGYjngiOIH0Jk7NDY9NZVSjLRHm+qQV4F3IRsNvNjuU9BgfIXYrMTEM
YusWj1Xi37WsME2Ru583n8DEVLdGJzCZARB9SHTlk3yBSnBLUZqsiryPTPz7e71R4mimxzCEJ6W5
zzd3KZk4uWsmQRgcXwSpXFRgvZoOT0fdBUnSHFMcerr7ORqCc0/7oeQnpCC1PlxYdfYXFCxfSdT/
ybrC28MLsLdUR8ssJT2METcBkrLvXEfKMhV3DLoaasao5KZvdA8lP7PtRgxq7Byf7TjdNdvEXMp8
zZFOV5X3Auny4LSvoymu0TxqX5BBk9izIf2VJDyVnkzZK0iM1Jidqsthwr7m5lsCNlgGvrbRVRX+
RShDijHTTtafnl/XrLpIzotZAIQAJm2eybOPWB50D0ipPiTH1UpkJq86ZpFozSCgBgyuKO4Nv/xs
SxyfAni1P0DMO3f8FdeT9Jde5Qjmo2WWlwPB9OlA7dF49L6xye7PczmAvmC6oaH33vs/BSQe2yuY
RkiQGAFXdiexDm3wtZS8E1mUbJczetKEU00Xv7ZxZRRiJjdMiFnz87bLZzo7zrOnV1RxhOTsPR74
geq8XzRfXatSos0p6Qtlg43e/65i4c1hUEoTJpD3qVE0UpLhlrr0X/C7kldnj7+IOPttFEVOmrQj
fwDIG6AFI8vlXPuDmIUiFGLnNnrC3bzhQX3840wqyic1FDxT3jsdtWfguu2iBncUWQePB8n0PSa7
7njZjuzpxLB3P8GsgoIPhznbNCmpfQI2wcvbeV8nq11EL1p2uG6/RombgNmj1lWVQXavHbJ0BvXR
/Ts5RXp8D/ZkGxRZTYpALyajaHtlERzU1swGEGuDPyURFkOUAPJjognCoTt79KA3FICpfRzqZb7I
SxoNY2krVikhMZs8i13m4FQce1JQvx1ihMD4I8UcGjH0dZlMJPQROW4CGm2/l/jPV6tEeYmGpxlE
Egyj5K/Hhz8aeFwFntYz3s2I3cTwFE7ylUiPeO17xxZEXaYqacsb+0KvH/dftH95AN8sa19t6RvE
U4sLEdon0eIH5auPSfZO93nSgw+TbE/2C+Y/IBMSFzfHGHQroNp+xC/zEIqbn0kbaZKT2jxtgZIQ
I8MupBJN0HNa0/Gp+3/vKMqBKNcXKi8kxEZl5pLezsGHdHra2HkKvXF3znVZFLMx/gqamDzvOzjX
CRCYHBOh6smWNlZAEFn/7GHaIhckgHGxvyBPnS8S189UNoRKm+TXxItUlPSvrbrStCYH6def/++1
TLATpc4LxfN7NeyHTwv+9WYyjsNLWyvt0/zVp1M1EJ2POpVvMj0QBHrb1z8NA1Sae7LrTD+uKoIO
X3q1Wct3Fa4/nyPwLz1kRdq2378LJYZn/hvGa8GE6iOQwr1kEILVKS1l0WvQL7XjsdfEV1prEazc
US/GV36qF3wG8oI7dW37m1Y4l7TbHw3rdeD2BrInjUvQLB05C9/Phpec0/v7sxZrAUZRgQhzJoGO
CWO82391CQGaNfTJscZB6drpnHUMsmc4F+9Rxw/8xgMz7sATbhx4FtKXaYyGurM1uj6ijWKV/y5+
VBW8XfDvdL+Zipi5WWZxe/zMpOXZAtlL39cgUJ7Z6ThAX9mbupnn3HtjuvlPrboT8gA9aHTgejZ2
Wpq9+W2mY5nIsYGt4WmB5QPphYk4dJL+8OS3EK05JsiksCDIRXRvOv5OJK+jwCtTh2BUv+7vAo/T
tp00CwZneYguT/vHiRAu/W/T+NsA5P9mFVtRh3mvpTnmb0xFCOBcFOqv+t1kt8W/8AfgK/Xm3mXY
URWkQBzrNrZEzBgoP9K4pqcjGdP79gSPZtoQ4vxUcl+nZsmdscV/rrfBzAK7JLdWTmImKRsjNqcW
waCWzAgwaIc/b7qiZjhrHiDDUh8RfM5PxZu+n352zAQ79D7AxKJwuADc+M4ES5k0uRdxLfpMNMUm
eNaaW+fsgfBuIzEGH6N6TAbPcqAMo9K/LOiPUdHIrXkMmajGLdbG7zCVb9DeU9tAHkhNQ5lhaJji
biPYrENhbeUmz6F7N718ztkDiFOqxQz6Cx2/vwGBo84KnHphddzPir6F4Q4RxQnsBtLjcVp/5HSD
Zz2A7lqFFbW4hJfVHX3I9QTGnJA6mkSS8Kog5hh2wcQkiVujtkRXx/PLtuVM3kZmEbEDboILdh2l
It8wCeFqOIyXtq8Y6IThDf06RrJHW6lzkKrcjNIvuFJLrglnbOyFIaVVF5TQAQlmLkfa3jhojVXh
5DaJIKz2YR71Gyxkr4M1pfnaWT0HVeWw1+50b6D/fJW+NzZEro/C0qIpCY/tAVH663Ie7+8oObvV
8tLUDKC0ZAaI7RZHcXmLByVrTN44dAPtxB8UPNkbQKCYisezCs5UdCcQ8NPms4Aw/VNmcnuPkn9v
W5jblKD5nQ0wIL4YnGGx98t0CXByh1BLO/7qZpVs9CdmvziZWsvAcWCtih459FEeue8dvAABm1fq
V7cQ4gmH280tRGdOrIbz4x0ZE4c6XoAUINfubUJNKnClI+bcqF8YFmJTK6GwN8x6wKdkqjtrSOfI
Jmk2wF78ha1pbhWb4BdWCYK7pyEf3z8c++Ga1gryOgW8xRzICPayuNOaVLzxs63dAS+wmb6XTHPc
l6btM2gGg8undwBHwR0rggMPvOyrgg3l4aeGssgVoT2hRYmQGYvyx8AzoD5eRIwqu7U3rCuzw/Ba
YfeEDEwYAuSRxStJ15kZxnpzw1P7BQSYX1ot1EfKunQ7SLjvItH/UZUx1vI45CdDKN4+REzZ1C+b
d6a1f2CJ/IRf+6IL9RJxpsjg1pEq7R3RI5YsPuNI90iQg/vKg1d25CY1vnLTis44G5sN4IQy8nml
tiIMhOOnmNni/NZsBD/M+/isSVdLK2veXOqqx4NLHX0yusKxkjhkth4r9nnHpKtX6Cu17FIVm7/z
b0Lo+m7MNsNgf9iD6gr8VeoulKk3iLeZ/W8K6bKB8POlO97IRnikD6BCxfLDXlqrgg4iGmjDQW3o
B+EC2inNm1Q1BjVPZDc/z8CtkHB3ukimQ4KGVYs8hla79/XbmsQ0/HZY/FwA5HQoXnV10eECeQKr
P9t+2+9Uy1f3w/V4cX+qOoacimfvjcj1iXgiHdVJKGcPbqQHg90Xo9swl7oQ8WbmCMqR+gd+yZsd
TGppu3QU+9wigE1eVhSy+eegPb2nLL/FzMZ4EZTJVpNpPjqg2CnpuUYbd7fVdWwLmz7oRviZc6qf
5tqXs9/IqP04t5TIHyAy2ByEbIEUm/kKSjTTUxucZ0UbKfE6j41NZzgtIkgJyqM8f7m6s80j3MvR
P5jEDmrAuIQZVfuzsMU8Sscb6Bbl8I5d1JpMtEQMaNEGzK2ppcX/IoeVYL7RvcQqLGr0UNPKm+YR
5eOhCxpg6RdyXSlnErvjnBgQG7sWVbcEGiqEZkKADmidbGMN1xZKP097RgfgIDAuKrS1LVKl3Ewn
kGZSgK8uIF8/eYAmexFrrOC8sg4GWhtVKmtVeEycIdJu0LaubeRcZrw1NROW+eNlK/Bb2zcmbP8T
BDucsdDgc5Goqlwiw+wRfG41lVCnXVC0UMedwX0dzaTs/k2i6qoD8GTFZs27jQGmVg2xHUY1kjQe
jADgwfj6gHC84GGAyqNmBBFccqIBo5B7ViRmrkDHjzPt1zv5a6kD3d/VnIOtmiQTrKF0wICBgP8s
TFs3ip4VK5jFy0jm2o2RBp1fef3RNFQn9gxyZA0eM8lG8ECRYacy7RH/5KeoTCjmv9Yf2fmgfhYZ
S1niMqC9pm7j2RYPNyC2+7ChgvV0KhDEFXKV0acanTlH7tmkyvTIjvXAhynqAKQejdzXWGHkcQSb
Mr9ewo5m5LZ4t3nNhUAdomt8jaaHqK3WxXPdoKRbcCP1m3IW4iwf31rUWoEaVwlSBDGzQptVkH/R
MGikMmm4+Oruguic/QjDuta6mT5sjXcnehi+lwrFXB7zH+/8aoWWrvQERTFp1fgvJ3SHvfrv4pu3
vlH2rEpYqj838V2I0nyKywc3XPfj4457c6/68PFXGk+R8iJSdr0dnnYu3xqp0e/GriUYMHTvKNDw
7yyzW+uDqjxlEPhY1vY1rbyK4O7wHlOF2qGXXVg1L8ctsBJhG65iw1shJo5d5BXEpRV99Naasm4u
FecZQkBndb2vfLk5bbMEMFdkEb/EcNjt/19pzaMHkl66Jz3PiN167Ydm7CiQTcYfQMduBPlI7/tz
Cv2ia2j2Y5DEuEiNztmXbYYI/9fcHK2qhya/FLZ87hsE7zYzkzwruUsw+l18MgGytPNurg6wi5lo
wK0rDboSb1ayVAH+V2SAaH5BXPSJWa1pxsqzEQ6AiXtlX+i8PvqHFfDiPspOoUaJYapy1BiFMQhQ
BfVDVEcnK+Xh7BWAs5Gpfoyv1Dnfr/ej/wR+H5ovV+OA2TLDS2qbjS3I51bFV4bColh08oTys9Qc
HlDMqR+e+/QfyippEYBidhOUHjgcgmY4gyPWnphh8ehBx3A3sbj4HLuTGGmoSn+lZJ82HIN8TyUO
j5GeURgg5GoCW1DMpooU742gS/Focr3kJsZvje7mzwFzojJ2ga4L4nQGm90n90CNkv/0HB/DCGLg
bam/sJEoR9sFt56iVPTCJ9pkQnKExFACk1eoRoNNOItkK35TCrNJPbL3lHuAyN5dc6bBzH3z3ba8
KvZL8ZcQlaDf9LjAeP3FUM+ylfJOlU89fiNSIFeNHPnyO91knMPmM0SEs+EXGXbyhpQyvcPfA8lb
2fHl98WhYAykDl5LivLN1bMAhrEaZl823Bg3Voqcb1ymcSZpwhkNZvDyNSWr0MC/ystFqnBYtESp
7bC42F6SaY7cB6wPsm8/ScN9VzdtVALm4hBeAxwv+Gmen+1wa3cjkjnGTPDzsm0SpkI7/GBMTPYF
G14v/2X3lp8LXAxDVOxM8LM11jXd7VBlPQf0XFPTsRlV+MixmnGSzwouZQ+N0LQypNpyuxztK4xx
NhNQHas8PdSMR+frtZyur9AaInM0dS4sZUJoj8htXnuCv0+NhMZ89Pi1WoVuuC7LRJe2mcBjvMds
d1pxABNmIoI0vYHt4oPdhX9/Fe85p3e7vjyW3NuoABFqP8rfSWzH/nzKb5PL6tjwYL8stSBjSrJu
jAOHwAwomZvlH+CYxnZND8Mv/WxcwC5f265QPHTPxLu0frXTAewy/tekeitpgbN9EzwtReOQzrvj
7m/42oQaOa729We6DqDGP7imU7u3bJVkL4qOpr09nfTkQGtJ7pBNojKazQjlMNgdMGeVgeJKKGVJ
/DxwaNfSOpFutrUFHbd7HpR+Ho1JJQWVSL39c0UHau8bDBmiDgBhuz52eLH1StAsAlBj8jMuphkZ
EMyUiyo+DsvzBLPp0s9F0Z6PjskY9o+swWqi0eXfChfvK8sFqliP93986hcIBxJFJNUOr8iZAgbj
S/NZbBzluhkotddFaJK2dy/rDsnXPyJwIAqj6o/LmbYA54Jt8NuynoRPBbGTWrLCjgvAnAam3rb/
x0Uuo7vFhJMIsG/UGfsmQROuGCx9fLxhuuueUI9bbn33LTQRwqcovqzJOiUBu0MoHhbwtjXyp0Cv
pP2bvYLcYwXkvE/EREzjd6Vk1YTK+jHe9udspmNBJ5zxTCLTISrz3bPX77x98VDdn3oasCM6DgPa
IWZKVmshB94x1QwoS5pUyzeFTlqO3IxLGAkf483LSDKpWOZlPn050PoyCYB34Vi4V91mZxrFjfGH
UYVsT/pNZPronzvcGBA2QvWeI0dLpyhfK7ibwB+p5Hkyrag2G4SKzqbqtA30+laC5bw9/H59Ssiy
sMp75+Cy+SovFB1b/t0bCIWfEUae4ng6tw77xV72sITWuBtifHH2X5Fxj0o4Oj1oDSjDR+DIDFUi
NKNqaIQ5sw3z5aK6CPe7hlDbLhqB/8uPjYowzaHgGqTU1u2WllPHpYgZQudG/VGMhXYsJPxeLhuZ
tVlk0sdbKBECbSwkjHPb7oTRTggcT+16yhKsqAqVI7IYtXdvU2aYujEvjEThBzNQ/zC+4TpSB2kC
DyMBwh1d9TxusjoSYYJH1g50URV7q3DG8SXMtN5Y2OKG1jhuSopK3jO3lqkyRbsfo/vyymcKO+eL
zVmBZxRr/Uo60qGytzJxwYwv4NmoAZK+28UwiCxi88QOm+Vfdq54Y/OT8xhrckj6OZkyBavhCI1D
UApPlrA+fhvqemjg4UCseuqUl/79IZU3DockbG4C7ZZzMphtOGhUtDKItR+wFvMbinLzymCmVS6I
uW+A8W1UUPV3pl9vOPAseEmjGDwXv0jx/t6c9TiUflV8LzPVRW6bkQmJeiYpspBFdN1TFUmrsuum
Zj//+AjsOCYRPwHqtyzWZ66AUR0854c6vP9Q+GEgC8RNaG4qcRtBBTTOwK17CL4dAj+yamLHlgQK
WDDZu+Jo/VzJo3RezmfewMkkX+1Zw7zTzptRqdPbqaO9pX9oVlhUG+1iT2T/Jvbd0aibkfAPl++Q
D4klqT+34n/vhL5+Pk8hhoX5mSbEY0kwUmJwt+ntviHa6GyVTZ6VCKxH/E+8gF6hBsLuDnLozxZI
QeNMnCEjH5lkFsyRdhQAt3/pDhJ6nRpCcroebN5oaWTKoLbpCce2BhWJZq/RqFf9HB27SZptBzfi
VldHiTn5GrOU5GA76ZidXwHGPuK/V054TpMBiM3fGc8pbjHiTBTGZIpN/HU/FUZmnZ1KOpjQFZRE
ukrYInXYpAUZC45Mst5k1cJT1IwbO3v7Hr4gSUGQcIvnKjZZ/9I9R6Mj0LBzeM1xqRPRLH6iDYff
IvMD23yE98o41uu1C5YTgdpdubizdJZe61ENOyqJK5HuAPf2ubI4gC/e2ab45z4J8z5+0Z5yiqm8
lcfq3CffXhWDSstPy2YlKUk1mbi7pYsu6YCLw4d6BxugC7g38+VumSuYZAlwhILrN+MHKUz6YP4u
86M33k33CZqAgele2OOAAv94+ik9SgDeoLe5XVZeylThKAJxE7Tl/euaB6D4vkbFTZy0ggN8Pk7w
4N9Uk1sxKSy+OjxfvJhcSNPl8rMsKycfIONa4Sc+DMO/8ikkn+JhI95xMQ94iOlDb4dg7xI2z6Hi
vNjL4lUSYqjZYA8ryhaSY4KJicx4LP3D+whzMtlY5dEv2qzaH95Fjm8pC8VLPQQnI7wdlH7/ov58
r6/4euY3kCthUifqrSlCDfU1XIGA7G4c8p+c0mQs/3zh59QF3NZDQEVTrPjawwaP858bvdEvEzZL
qS6JAyOWf5dqF+qy+oZ8F2Z6szzh72Ram+qwvK7rNMV/jXLvp+7GM6ICxY9GFAmpmWSULDu/9Cno
JVsJKg/iQ7MM9v5q4eyo8Vc/ZGa95FceELaN/dSzRFyVnUhvEm5VEWtthxzgM9nYPCC9CVNMrtH6
71dk3XkG2LyS1cE8DeQFOG8ky6kP57gF7imp4oLCUqc6wAYlHz59+247KYLICLUiqAWrcrkMbRrt
bFypwvF96qCZ5wYtjLSpwNZNpeI3NmBiHw5Tde5Ejb/uCScw4Zmkh1fj868AshhTSY1G71SESI1/
QjuItFkaKRLi2pLzPLhyCnhGeENQmYjf1hCZq5aiDHyrevzEH2hothCbSopy0H9Px03duwt9tp0y
+wPy00/likZ2ixlOQYi/13P3PHUJpFVt99rAuOM/tugdb4xu+zecg0tjyeGxfaJXj12vRRmcbeqo
I4sppP4UlsuV/AOlUhF+IypaoOAnWicVy2cRR0j8VP7ACaH9ciFa1vGjNqfx6axECY/np3S7sTcx
n7Lv92WHijS6vGGho5FlwwIUgBacM0whKjKP/2nQKIt3PNDDN5y+vav1bz5DXj2LHfUV71SjHIpK
5PRqG4et//zEwgwo8tbFs9PY8mFIfiMQFY9jVJMtly3Moy7hDOSumoutDxcKNS3CQbByk+fCDnkU
i7+kxlSWuFXwBZqP2Vl27A19F5CH+GY1kzUV8+PJDIPxUOLP3vjgYVklqB2B/7YSeieLWJWV83+2
7dWhAflHaVfWYwDQhavyKMvF555xwBs0wecRmRNxhug8rcKtR+NKSL5A5Kx1RYcKWHwUKSPDnKZZ
51io8MyOtJTjOSlaLGN05nT49SfYN+tyWcAmqXUS8XmdeyV/5qGOqUeyGK0c1E2ZAAeNrFi7qa79
nHhKqcK5PpfMPmOj/e+fY8bBoZgqepXq44B5TnaqaKE63jw9gayBG3B+uMtBq9577aVbDfG3E0GV
89q/KxoRVhX6+naMFdNKd7cS5TBqzsfQQQIyZrfrsJOF8RKY+sKVq/rLs9tSgNtswr50jVJowh7Y
Tf37dRZSxjTTCuu3N6qt82jz1lOjz2BadGvMHsGdmhripPrFLtcqWSizg4fEzkz/dWBwzugzWXZB
sEXQB0c6x4uO60hlevxCgRc3inbnaN1CFEgKy0CKxX0cJyfoa4OMT2my2ummthxDJtHAYDsaSjaq
QL8X1FV4CJnlE6xvJdtU1PhHZJrskwoS50lZcXnb2Uqlc+qj3DxbYr7HKGVoZ/MEb+ilShhdLpoo
7ucp+O2UiuC+ToL/uqoODSsAfLl5jeQ8Q2aQ9qkVE3hJ1oWej4BQs6TaEq41jjd1UvD9N5Eu8r71
8UC/z5BCEWEuZN2y55lQon0QGNI4+ggZkOcQI/SazxnPf6uEiRtKD7jWnYYXKmX0h/3sSvbq39pG
SbEP0LDstCL2M0DvuRULqiHpm32JL2irq1zJ+8g4y9NIeDbBbJwMFDN8Zom0Zc/G/C85Qgc24NNu
9mYxo+zWzC7W/VcI7R+klNHJgUHUQS6ffk45upXchVKU5JRUxxpfxJqPdVhB6XmT2FLLok2BJIVl
0h261p1c5/YoM9nHj1XNXGeRdT5zoDSFRy21e6LJEq9dBCs8BlOJD56D7VgwZsIzIyqoFQ4vltXi
936CsZvVwZ9CLcnCtEUv2Qcq+Ny98wysuzRWnsRHaUhyO/VZsmv+3c4RVrM2bvWm39WgahEvD5Po
lceXGxcAjczHrJ1Pnk/SA4VtSnLD8C6ImKfvNEEcsu3w88o3PU6PGw7L6khFNC7t78xMFYjjioK2
u8zq3fj8boEgNyvgCSf65ZKuP3gUFKzncFPxeVH4DRZ9+trOmLIDxeRVWaZ3LmYHx3pBKcdaQTjs
LXZv1N0WotPYFGmHmgMd8oZEmdQvN8BkGA+NETMeJDm+a57k1P+gnrxcuSvRZRwNP+Fs235I9F2s
wb3DIo7h1gAsUgQnzJo3NVkXZHaV3R+uvkXXTuuADAZ6jPBCORKTrNZz2UMjEcHiK12EaluhzCdC
mY16N3yLWLMZhy+oZ1AA5h2GKtx+bP4U7G8QPZqhUybJXcM856vLIKy/syzI904OijUfFPyIusLh
08dPEAdhPX7UOcsTVr+hdTH62+jUGZdk7j9VGtFE3AwWVPHCZbNiR8o4YazbV/DZjHemgwFnGX9E
CDFMaLePD6ge+3uF6bqumKiXO481mBgRUF5JAA6p/q7uWyBgfJrIKCo/rETyLTKWEcP74gMc5Ho/
n3y2czJQHIaPYfwJz7nwPypN9o5mmjkAl/VbIU3UFVjLb/Ek2lU7TE+nDfOAhkaPl7b6Ua9i34tP
zFD8Jo6BOZHJELECJYxAJEgFcndqljrmft6CsJaD+YM6YtnRd6FOebP7yOLK/nZisPur654ToZ/v
R9VE9FO9scS27HKqcoorbvK2avOHuThYMjRJDYo7+ETJ43CjiO+iWcuZqZDKy+S/tycmfZw7um6v
W/bZJ22jKRlnHdJSTqWfESEQcpGeVSrR+Dgu3gbFpgZwlsPh7+PI3/ofj+msGk1aLxSJDtoboYfi
bCeCaFmFXkWx5gWcU3/P9cRyNUayoJwOEdJUlw+thtOMnfB0XZMNmJ/nuWNbVK8m+18+i9mttwkc
BgcADtKwsxQae3GDjCX9peCE9OzbW7UQ1gJsNmBBylSnEmTioAzBafK95OBs+1zb30nvRT+6y7T/
vKyObiEz9dMyXT2wUhit9t66T3KBAt8TrTXF94WVC0pQtvjLJ6xYiVHLL01rRdsJvVk1Quu2SR7t
AWEmprpxL++PorhOrvU3mXIic6qAUYHYDJby6g5WQFxQljOMH/c4SvznEcnF3qGqKi/BnQwVwuMI
/GFzz1arNJBpYQdgx10PUsfRn5Azj+3H1pCvC0mVeKBWZCxQPXtHv5dJhW7mslRXlMHNdebt+xLy
OHhZ1Gh0GzdHurxIlvTioWAhsHkvaw+E4Q4CFl2y/5Ovwl2IvweXvejEBi2FPN8X8Asf2I4Md4rk
azjwy951/j4LIKvEGzyGTLuWyoCpskFG19MCvNXU1oUgl85SEQZc7N6uYOoeJOumtnQmdAzp3trf
pJe1qyq1RCE4279hGWJMMs9lK4fCw6sxuw5yXWPla+2W6Km3gC9n2uWQOoDayPhRFBWy/aDDcIYk
TVrngfHoyLoSICj9OXSSW3gCRgYlvx7C+mb9ygitvTEaCM/Qgtq354clWtKHbQrIN6AHH/UbRAkQ
l+hbhYg5vAxIhXe3F2DNWCTyJWDMtBBDst9IZu/DhbT3FEILqwJKUcQiUwqZcECs3hIsTofvMgYW
4KShwTf3B5ZzudSTONUMIBldVsrAubAirYQHoIzAv915jDfBZhuQ4yCECrTwfpqr0HJTBVd/rTiL
ODtIbsMnYqadROEvir9Z6XXvGnYBhaWZ1IGYjXN8btWpR4oBsSthqEY3r+O4YGCZlzDzKmKgCybB
F7N97fhNG+5Q/vSVgRWCXRX9HNAYe8a8pikYwTqIEuyRxWJuPR1g+OK0U9ijFwv66LxIJWCym6EA
gb+bb9sDch0FAluOCEOMr78YE6Q3n3jZsP/VKPuiTggxz6/PSMGd/LIPzZIFVXL9zZ5Bd+gCPyPw
uWWrRUWxYDz4o7UcXKKDQYvmgwP90Rgq7MKfRrhQxRxC+O0urnqryyGlMP3JI34R96u3gX6OUtzs
6LqyW0qbos4idYrXtn6lZYCnZK4chSS1yMBacv9hz6E5KktRrQM+Cu/nMalDOpJNR5lQDuFislCC
SPN7m048+kuth3MTuYyauCZ27eMXDe7OGJS8zDvKaqM8cFSzAKOGl4dVOC9BZjCCvWeSgtMsIuly
9lU6ylkWq/TrBD6RVes/96sYdPYRLo/80x5rwBQgTbuujpV+6hnremPHp5OvX7NresOJdXd/PtZU
XGjo35qTSqa2mg54gdiQUtywPLeFaP8D+f/JVFwcAUYsbKIDoL7g9yUBCcETW8lINY7emVUhFRko
K0fpYXYlOBjE+y/0s/dfVlDZU7s84j65HA2BrLELXJ1sHr0k7U9Z/8HlA40YkYaoqsPtpBVT3U/y
u0SPTMFhcITbGZc/qJWp9zX72Ledv/r0p5VxhIDCzZKKT8vd/62BIHpWCnRpyUuqp4L4SIUTARes
RiZtmVs47Q5stdNEoaO3nsBc0RcfO6IxWNxVgiOiGHJ0S/gmRaCcGhXnLlQ1lNZRt19tEQX2Bvrt
3fW1v3j4aFkDUdOI9Ia6Z4eZDBo/ujvLDrTAc6991sH7v4KjHr+uUEpVkQY5+pH5GT1HQ4+jWQDs
ZlRSgWq76W7gvI/U2/5gKtLXEDQ5mRKsmlZqEV156vkGixxIqMwRpAf/aoE8eFrtR5pJjS5AwxyZ
27D9Uo4lTzVs39n0WGII2YMtL6jVqjmA6L/Ks62jSHoRcJ9Q9b8oeNAoUWWojMPJPLviRx7nzqBj
/3QtKhAJcPx3qHs+epJ0RwQJpERbHmne4V4Fr37KT/EISyBkPZp2b+Ilwmt2eySUoeUO6PMAY6NL
M7hACdUqOTZGEAhZK66DyQlRz7iAD+qRF+XTx7jbWphCgsJKQvknO0+n3ACAAj9vukswOb4RIpik
jp6tPBYuYC5UleREIsImd1zNHexlf+ncXiJoRliE+ElY4lsklFnmyOCOCFxxyySztxjvRwfiCesD
i1iwrENci1xePsjGiZhQvROiy5UerfbzaxsjC5gKUR9wbvQr5F3NItDLt1/nnsJMZF3QnNewhMvR
ry17VTE68hOWw7mBdKvsupAXM9Nq+/D04gz3GzEra8ljLWPd4peQ2DAIPgkaTEecWgOHoctoJe11
nfC/ZWR0J77vQp9USYv0u7nLkI0M3swpk69I4gePrEJtdNuzsweVAz8TiC+EiI/DQp7rZ2ZkAWXI
gly5LkqxOIjSe0HADnmY9SmWI56g3emyFU7fs+IZgH1aZpZ9G5ZMGC+5DJ+7D7LVI8dnI57ajJWJ
H7b08G21+0Brz5tlvWbt2KFahnC7ADrYV3GLt8QmFCikvQT7rE4NK/L4NMXFYhUppxmvX0uqplVQ
+ZMbackSVfrWuz9UCKutPfXmjVDwYColRhhTU1onGD6Iy9RnQLvW6fGd+MJYtWrHfCJug0CvvcPa
piLx5g96AgRUX1CZRyyJAXqGjXpAgQZf22vYivjZKRbZIaRvrzym0Bk6b2sPbIT6Gjv5G1odqMU9
L8n5p74dYOikbIEP5D8RNvsU6CuDjgjU0j4yGH81kAbBi3il763huvNmM0RiH8r87Y2J4ahK6oBY
jWXBtZUj96mv4cVyrwZ+fJdqbG35LCS+VmjFFXavFYiPODToTC0JL2VdzYBQtCBbAZ2EavMS4lO3
ku7mWp6JKvNCfPyCWHQhaqYIzLXkdgbFJWNunYw+iOFS8iLQM7xaoCn1qVE8o+lYQeMInfvv/QRG
Ll8zSja5ZqcezcoLmMHHgqJ00ZowyYEk+v3uSm98i2dkNpXHjTFmUEchNmj4yUtQHMKdalyOWz3J
AuDnZzZEMTVYY82navDaVSj26br73Vjd2xmZpNWImu418VQJ5+6Lu9IG4lEX4gDDaQREhdy8NUXk
/gvZzDyiD5qtwrvnhI07sf1IuR2UcJ7o+ROdopv5PnxI0iJPDFgFgcgEi3w4HIshXd9IuZjaNwvC
3xyINY6WrmDdRivKY2Mf4DrZLtl0332a5ZiSTNd/KtBU6sakYGE+gOV+Ud5vmCz9gIuIv6Zm86Pm
1qz9TuRUnh2FS2qTbBhIFnBkWKO3tSh2Edb3sjcdzVLVLO/XeIslJg0IVeCSkyWiw84llekUNlE8
5LbLasWhw7IzbajbXV6Ow9L4sa+K0uuYuNrlqmW6alUpyrRsnwI83XJjfao4xckNRmXoiL1rebCJ
j2MELIDxgNiVKpbvK7y8aoj1GP+VsLq3BjT4lJrY0N398GHLldzimhVBnKLHNurRbHbAaokqSYv9
MDSLoMNs1wmp36zc6Qu9FXLj0rtc7FY76ucP2KRIjnBg5kpN+25/nh/JQ8Cv5I+7ob4ltW/VxFXf
6Jc8iWWdyXTtQLHsYl8dU9HyJjFFv5dY6UDo7USbw4ISjizjLJCT3voKg9k6qERyqg8n7g5XtANx
S21u/+WEi3Hp+Z7KO/uEGp5v+2TwAyqzoNyFZ0MMu/YedEKBACjp3hLyR2SRG2pv7/nL2tEsgUzQ
68+3S3jR9YlybHeH1GaUtQYtyxOHTzmThjNrEA546VOweTidbDTBCZ0glODUxcNer4QHhBwVMC+H
92U6Hma3V5asCUkt6k0yyRAIKSNeKudUJwfOD7aewvKZLQIf/YenfyMQ7o3OqaPG9NT6QKua+IxR
XrsgVfqsMVsbWOoaUWwv5F4/Jpilkge+Zdlvqz3yL4cnwxuSuWSoBT3XauF9gs4xLFJoc/vO8hoB
iWZkiCq8PUPochFJsofraL08efaSzgCuqhzMQVHoIIuWhvhvqvCwjbqBnofPkSuU6rCPwmyuf20n
Xw20nyuTWA5xyrEtwvluQ9FFNnSVehQfJqN4giCHU1RVF5QqcOXxZKQ+H/iM2n0dbBbN1QsPluSS
GREPqP4pCTUxdVyVzfSQ1lIIvLQ2bqHljMiZPyF4Ubl+1O4zNtakqyvXitdchiJ4/6F7ulG5xffj
JiUuNFGBLU6pab/V8UHmLOH3kp3h6oMd2WWN7e0Qnol9yN83i4Hj6Q6sVY5I2IF6RJHXGixiIVQ2
hXWyOZ+043QY+BhRTraibdB/xqVuQCnEH9Cb4KGQTmNyDs/JBILmXyYvW+QosrMDMGf5OYeE7b9m
JXj7ZIN7jz9lO7NB+y3PPKHFvBFNusp0RfJnQhqoPiejF8/6uxLCqX9pwdGoE7dCcnsjOW06TyJz
6wvtg4zbbHWD8JAVj7dWDNaDHvvCGM8czFkx/l3IK0Z4d60mbKFQ0htVQjmxwRoykLmilX7KxXAq
UeuIYM2YP/TIkIi+clq7/7n91I6tuj3UmkJAnv4TEvbMzx77HjtVCnNqG2aFK6Oa0p61iGgv5ACx
MpQEAYNNEMo5OIajkI5D9VDWUiUP4hl+zYgJ1577VPAzu4OFPorDb6mnr2PRcwrQlzMsnrcqmr4C
akimZVPlraG9wmiLZFKNuytx9siCCrtWYX0we120stiAQdmZrJ0sCQjjAUrX1eJRDri/m30gjlOZ
HjppU7A7QLOeeG97HaEVLbACHPKLw1NIBDPivb1yQ56zkcoChAOuL0GM2xZE1cl3QG2OzNC9oeiv
ajf+nxLLISDZY+UepY6XF+a92ecil8k/pg9CcYkC74t3gJnaJrAHZhz4lyvX0prk8lPJ+FHvfY4n
pXhFvIy+Iwq772MyD9EEX8XeQquamGkq5DdueNiQtPqfUn/V/KTr6v7ynYI5ICXkZzv0RFKKJJyi
Au2ayJcEGTcXUniLAz+B7hKkMV9+BJf6kfua7Ieap/ZOM+b4Eum46fB8zyGTFDeX4kl/zj6vVtft
IeJiFkEGhK6ipogTuP8vTmjHeOP8pCp4nKSOTUXBm+w+S2fCluzUqi1zRtdvM4vioLrszM5EOQMw
PLq+zIWBNWxVP93b7n07oGMegnaPRZy6wIedhhXTbfQxwFLtuRtNfBYLCYHCP6kpZml4cGNntAGe
4epJl7MLhaaXXj5fyu5eFMNhfNkp0Jse1eg3HKyIpMJBLBJUCBRUMRPvOcKAFBbIUPcAjUEr3Jxd
jpkMNzOaBLHMD9lZ7aTgGWweExI8IAB4MISJ0rE7mlenv8MXVXuP756wk/sD2L/wt0HpkZQJm9Iw
P9b356e9saJ0ERS1D9v5ODIQhAzZv08XryIoxYN2dz6S1YG3HEUELYNNv3DIiNNzOEn0DRlptMXI
30YTkKLfM/WCRv+p2h1oIAnVi7z6nEnWh6+t5ygl9rpn11Mp3e6Wfm4J9NoiwyUbaj2RXLwi9Ra3
94coOmj/6tGwO2HLtFLZNmf6V/q0njmHHw55YtvEPn3dGNOXsE2RZWsVe+Db+bs+rUjUgvYBgjaz
XZYznJCQL/FiwehzbyiYblxM82IHHUFKXwHpKLVJtRi3IrpETvg8Ekys4l1Y2+w6/Tb5wR9qa8uY
Pi8xfpEvC38Qo84nC1csa9swQEMhyXWurvtPr4LFGnCDHcumdBklOhzTxWCxZ6QFXPgHhH8EKyIk
YDrZs3UYoiWrnLYHoBXNhcPPzBQqv3oURvBug9RE/ETspGFH8Chvv577Zo15YaJgaZmAB3XEqmAY
ENupaZUcyl3PJYnwYVZSu6YmaAd41cie5OQ/MuRwgYPxxKpDuLTefNCK3LNlbwdW14RJ07NPvBMc
TjF5n149ypjU0StAHirlY6dXBqgwDHGtSeT8M66aHUX1hERoXZnuwCOIcX3DyvIgWhLJltGEpND4
wmtIpydFAR5gvX6L8AJFqnWAh3Emtg0dW89TQgHRet+rR4OCmHtxOQ6okWuVf6DQWrk71NqocBwC
4Dbb41dEL4BliPG4Ahg9ipatn5I3p56AnyJT/JOfohlOSRs/LRvqMGwJIohdgCPVzjY7rkOkJlXh
WgOy5uhhVLWyeyugFZWAV59fhbUIaC7SfnNX8hHnmHiIwPuMshWguF2UTBFqayWTIUgEKjqQKI2b
vURGMB8mXIfVxKaoCyBDRoid+RSSS6zHGspydHJGy58zDabCfXOhnfRJcqbsGXO9VNHRjuBGZTix
9QZDPNbICUGQqRGsuWXXyX7EuurYsWhDHw6S4kraAJ+QHKk+/jCbQMD3+fYCzK67omMVWXseCLxE
Xo2dtaL4lV+63l+nsSmJNXAkFaxXwLH/Q06yCUWWoR+gQkFVBOumCsfmN1Kwn+N0YbBBSTkRxEJt
2YkNiAOTyFz+TMIzHEIy8NQ99h2CvcR4fxB0k1dq5qU+Ma83yzkLVpMpYw4DTB4hDq62slACTC05
iOSOS5S+qzBQCLx1sLsOLqTDoWjkACo9vdxPInTi91tpLO5eq0V2unjhhQ5buQyRM81yoZPRbxAg
OO+7S/ePmX9vPP9vUfictQ/bius4E9z7hCaLo40Y8T7imG/PDf0deq6hAag/yI4wM1ytSuL4rquv
5ukHC/zmHE6GLN4id5xPVSYKsjsni/j5XN5E8vFUnQOqaAjHI2zJWXfth0hNxkQPIfHAo7mBifAp
gJ3bOZkt2d26JUfKBtglwVccQvM8tKNEjIwajFJUgE03qPv3wJtC2kPQJSFmGUPYzFdW1FafvTdE
9+kxiUtPR5ofZWH78UjIiGDsGVtB35mSzfIzIBbBiw9XdHS+QipnB7ty87E4PxJHLwkj3Mg7yeaN
h9zUceRuROYv6/782K+RB8q3nw0+fMCvv2oi8LohBZiET1QZmhtgbT7pknWfAxhCLE3mtt6Bkpz4
BexbNeMReS4t8dnA2a9D3NsFWSIcY7hdzz2v2hsM8BJtatsjzgIuHaSrcmobhum3xp53hdaz0pZw
sPpVi3S1Uh0mcs1RWWBmBEF077eWqZnyXUn9velQkbIVIFdd2b3F66T54MV9DBQAEHK6E0OOYH/F
lJ9Sr8t606g7DgzsnyhuGHVN+58e89SbtKXsZAkKXHHU+dWFMbie3kCgz2vMWn4OPWUfSCyzcPr5
TrB0+ay9ZQmxpwEVYYqs/+UjDXCOVztmHOLkr/CzBnB92doe0uW1axkoCnWlZAVjEpJkDnmeCU0/
MANQAcaQl3ieQJDSbtZTL61yR20q0JyLi9PdohOTviseZzUfrmGrNAbxG2DPcdZ3j6ojDisBaWCv
kSF55N5lc2EHAVSOrfX2fTnTNfjuNgnZR3NIAPXBrIVvIliKPTlWZIPw1ujvxQr9Ez9DuGkaAcIb
Nv3QzzudfJi27SKU7fXuVoPgjPlvHZDIo7CBpZ6ko6AuCZmYupAnjxQ5f/atcYyuxdNM6GHBRjBw
yAuFI/lDHQXj2ME4kzMZFni4OWxrScVSBVsTmVND26ADgMS2WXJ34q/vEtriKv6YL4cvkHGG5F4x
qn5FdrNfxXWSBqaVar8jv/Pjxd3zezCFnIeS9mGSka5hpUyQhmtms+NEn3MANmBSM3yorPb9GFMq
ynDeF3VtMs8KKTYKJCekpElmspirOlL7lhMx7TxS/lDC62bVohfyhlfOV49L0l3Op4gBNWQT3mul
twrusnoa4IZA5VYZO2NnLMkneRn+maAv6DObQGU1ub85NzXEcTcpTFDJZD6oZE9Xcp8zAfsWskRK
Y1qu8mKvU86fKiH9+OAC66Ca7tgMsAS6XhdIHHuKjNnH7/gHwxM2+apXgxZqJ+/M4FLp+QtpZSNj
JKthK29zXE+aJ5K2jPxjrnAFX2SMPGpCK7/s8RII7T7jXQK8ltDbVnOBb1qXOWzmq7xskGB3AVz/
N/ec3fSkZFAEjZxONB2LrMPiGKKJXGbpEi/BsqlJ4htJLUz9vkpd8bFMjjRrGy/TpaWeaJ8rbEjr
PrVzSZSNlMz8k72H3lXTWbcj0k6feZOkgXuZnKM5eyeut298rStyRTkTCdY1rRjEKWSWJIV16/D1
g5YXkiRfunLQdVXvlqy5NfN392h4tIHRZ4pFmq8rs6YVCDqkuTr/THbYIMrz17CDMuyP3JsVsmVP
3XlnUdqS3VoyYWRBeOl/XqWruJfteo2NGLCkqXRysBaD5mxF0W3uVrM9HDP4281zQh8nUdHQIOU+
IlariqMXupXTcFsK3RTCdjgJKac34tR0SoN7cmEXKINCF9cbvsSzky8tmO1OF0y2A/fkBU64EsAG
kSfOdmw/tj9al9y4Ofv3Y7S0Z4LMRVOZ2jhc5o58dNpNlKF0DN0Q/MIHY/Guwh2ON7ycecniieeH
QzwD61Yx+8ErXtSIxZxglptRiiiPL8+AMgfKvR3CK27pxVPSbwD1avXeYYxciuVUIAMRppINddSi
cVQS9zg2a7lfSANxgR3DBCB5l9HRLII0DrTNnUSqZyeuTs4uU/oU+5+ihwGolYOWWSmI7iOPzR1O
Qvvc0o7gu6Cowm+1kh3E0R4Ep7zjAumExkRZ33Zr40+QwBMsbqLEqmGRkteevjz+JBpGblbYaaZh
DvFXMXxQG5I5AhSU+6a+7nj4ENZvxoc+IYs/Qnk1ToWytJ8m34xg8bc7Zd4yzL21Xaw8vt+q0bpY
1uwkddS5ijpPx5m42mAJhEHalvnThZOYBfmW2xzVSX2xlApQcYXXL6WejoZI9+AQhMbrr52W5+ul
LgPpYbEc8/41eftEHF/QiF21JDGX+EO9yQHy3l7KzDj2DPwYSDswzqL0U9rsiTdbuGXWOABOqkIM
5X+X3AA+LwOQ6rjYExoclYP2peGsqwh6WoyZSxyURdv9sdRzb3h8OoEBM0h1En58rUvrl7VnEdFK
+G7bZD2MElj627Xmv6TXmsJvnJy1sKXi1PTOEEY/k0fNp376i/vbez7A5nhDYByEgXYfzjA5NUIm
J0KIEgl9DHiWu0NlyXE+mCkk0Dg1VmQmqEU9lfGd0Z5pBCOSQ64q3TmgpCklSU+03FbnAv894RWG
3dP2IOnUo0iQcKRFJu0NcaPVaYDlYfQPwy2dRq+FGNeREF5CecZCspqkeUT3+KPVzdaFhMIC0h4y
cqnW/f5UPJ0lPns6ByjKQpkWcgkBr/1YifHfPm6Gagr+5GYWlN0RqWiXI2C1FlU+FE5RDeuQrrCK
Y67x4jfejZu7atX8z4NLg64ingqXq5KGt5XGWM29I0pu6faYwthWMjLQ7ivvLsRpnI5tMjLOQ+7u
Gt1cYO+QRCp6TAaSW0UvsZEyggVri8mj54i3l39I4bvkctBPCrjvP78+j2y+KCnftg2wmWiAxCdV
9n8ORB2zAW//1ICNcnVajWr45NSsXZykrd7Mn4DICq5TXzaKVvxyZKWvRsGp5n/xehClOTKpePRn
ALWlQo7FXzV4VIJKHbemDX/St9HT2IQeqotkq/IPECVhp00pPLcicUkRSc4GBvMulyqjj5mT0KpN
u+MLFd43ZWHevJmn0JkcomrK7yy6BxFk/mqpU8K4J2kOQ2N/hG+3ZfBGDrtO0Vz6HUXGUty9tD0Q
ig9H/2r3YOlZE05a097bybWwHKHoytoa2aTO3CnrGwNbT1+A8KPbPip704nCodV3eVO0ZPy8yVIi
gslRwGM+Zrxi329dyk3pwpot/aMjwbYFk4+dmJvAX/40+hZ3j242jKqkPGAiaTIXDpeQch2II8EH
lNk2zpq0PHZaMGC8QfX+Q6w7oWi5F/dvGxwDJ9JxAFxldlXaJrT/OnOgV0cD9EDZwd1Zq2SGd5XK
VZnB8v7AHDovhc9VtbcEyGgjjq1a+FBzDb519uc3XT4/Q5ifdLh8gDVfpwZVuObt6yWh0EC/hwva
9omfSHCWYlxoRWsRKKfeOr9qOMRW8/wGdJx0RmMne6MUh3S9uBg2P/gpFiv29Z605vy4JjM9WRbo
AzMafLwyZqBQ7N+7VwRoIWyqk73umpL837gQTxWj2Nl5q4D/2kAckn1YVUI5HiogXS3vHSKDZy/o
gBvwBBgkXQHyfgVFWen4vdA3ylADUtsTk77tXeCailuu0zp+vxLICKLpZIligMpZg5p2Xvi9WIhc
oMmAIBsEV5Lr3FQ8UIomGGIShzTh2nuw0r/TKFfUstTjw1orzZs1FRkVKY6lcNKGq0SWWqmjL0cf
rq9RBN7o46dt+CPS2h6oLJcAb6jo53OX1lFPk128BklMrnto6bXTHE9RNCAQ1C61XWv9SsiorIre
dljQav/6FaYeT1A2ACvZmsDWmOQj5oZYGuHVkxvggC5aGvpKGT5Wlow/+yt/V2TQT8IY5uSX8c69
85y7of0dIISLGLOsJlEOcPdHyEZqoPLZwBbBdqt7hZk61hc2emHQuOS+kgS9nOHzjLUb18wSNGYH
wYKqM2zWv15ZQuZ1+nKtY1e/AiYJiGr1uvaqiLLe/opJB1s9K+VI7/L3x2hC7D4DxvLHLn4plM1r
tns7J/Z3f3ZTxZhQ9n26EcqjdzFVOToWTbwVfm05mzLwsxYIlgDSH+10ta6UR1dz/1Mkqm7h9MmJ
fXHKqSa0SM9BmRUpOy6g1ZNHs/1o2cCkRcrwDJzY3y0FBQ69KEQov0BxIlJykLFodlmvO51kUBYe
OCCtxQ/49GNzuzJOStUbMbQ7RCqbnO3qrxOXm+q+18ZCnmUKuxcFM6JkNKRnuvWZhlQ7tIwXZkb+
WEOOa8zty3RFgmPJBOPRxWKUR0fcvVv85yvP2sJDotJ0R5ow7EpxfsgG507cjQFUAFLX6bUQrYTG
5dgaqmAUZMpIODcTx7HQPMl0eOSS+uTHURRmD2/3dxo5OSJw1kBqOn/dKOr55GSgbCAULHryZKDe
J+hBWSwdEoFeKhIFck/0kxmlqLcC9K4HME51HhusZ51dOQ6o95AU/MTQT4r7qHsuDRXXzyU9i0ox
4BP6VXOBgzlsLAZMpwwhx+8fvfKvWhUMEIbH6/m1mjgaTcjH75jPIZ5ir7wgVb71/EFD0krF6ZMH
YOebOCGrsl4WmLPKPX78IyVoQd3vrfqRRKhre52ToaR4fliL1YTW3bMGGybzGURg5sx2djYTWh3o
PwKwbnBS68ytculRN27zDY27MC6wpbG5dJSb4UQMpwhPIjiMw58O4fP14rsqOSm/6wvcxSuw3sGD
8lUu8fc4GdT5OQTiXBqmc+EqxVnOhFn6Lal8yU0ovrr7QWK+2J5J1sXrdD2bylHgEQZ6kjZBm1sM
ipNlvEYdtdTnfHOTn6SgqnycmfsXVg5maDgTjZQ2tmAJyzUlQeYfR07iCh520twP0ozNEtpe8CNV
Wg1MhU17NCRHEckauo690C0QbAHREs3N8Mvuj+22GysJmvb27tpH/7iqn3Z/CloagHmxbzKLnwmP
Yor+ss/umcyKqucf//dLjJXVflYkLxLvaK5K7frIPjcZW69gKRXYmHPckoI4ZFM02dGPSNmTQRmm
+HbY4EVXB2ndAIvgRCfvQrXxWSie48tuVU1RlVRwFMf/cm78+at/SFg7m+a+ZO0KYHTZSYe6K0kk
UNSXzfVLOjDOXBeDpoR425AYG5ggyt13v7n/Mtyl9wpTT6Kaaq86cnYEda8dKs1IzM1XATmbHaC2
YZ2wzdAtH1G95P51yFQmgM1na0ExvZ5Ktvhj7pkd2LJxKuv7FzzZK+ILaslGq1c0uWcf25/oBx5S
ZDOhF9lPbCB5RZ4EJgHJD8KynvoXWWCXQ3LjkjWWwCWxqKxn32JTUITZRrR1VNkaGcMRl8lkzVT2
pCuzfbxGex61nrfQo3EkDkL1FOlpcI+P/nOvxDUsZppY5D49NDwJbi+3VwINwR/iUicLyOHkxUtk
9a5GZJufnJfszgi6xKFAhBGLvpHpt0wbu9g81t2s6UxHClW4OxzEIA6yXT4/zTDOb9Ue6p4ZQApM
SDIPEvhyxQOeBY+GcxizXJX1PE1cFyLEOLD7D2HF32Fu3/z8t2hHx0MzuYmO9axgADWJuQw8mxlY
sVfhUY3SQY4cQb7YNedRSqj6eFR95YeBfpDKz63lgrX3nFv5c3H+NHgAjkcULPPQlo9U/Z6iSn1i
gwUyFbCC9uVLC9w4v+ghZMKSXppQ7VUyT528cRwr9hnjveqL6vJPetIPHPAVkW/XJjOSGFhUf6Ub
+mwCp3labfpJlJPq5G1xfzkKBA4BeYDcVxC+6iKBjbzMoPFWc6El4V7k/64/0ctZ0BVMKRE+nTNg
+3426b1JvaP23SM3PSsB22iL77yLMPplHnxAlJInJMk/VqiobD0SugY6sXQgLftGHDN2Meg7GDEu
5aHYqw8Nizgtp7pcc0sT5+oznt7g5sgSnu8DnehBnZDpTKrangEXVtH5zUWoXATUUIfJXEUa6F43
ZperJ3P5zmVi7Q5XT29YnwEjWWetJS9XLMzsAop1uNosU7kXzOTLS2UZntRBNkQhHvOvBqEcIm+E
PxGC00najFsqB2Y1XV1p5HHt8xT96fJu8h1+sYtAL0rvjrE4i2dGgA4sYTpW05mXYHZo62B/dVSJ
TmTkebu82sJyocMgdcnt7mz/sgS/6CDJBYIoXhvmPvh9TTTjb8ML14mfOXxj2zXPX4Z3/DCApeDP
zelkA+F6TPJM50BpeQtO614inMpFyX+lsNZ4PeLRJZ5dgwxxcbbeSXkuib7oZDPFtCHRCpts5XKu
8wTPFgNvoxnRWPjFTJqs5OLurjXQKw4gTlKfkt4+CXY9V97qHuumr8D5Ui8uU0NFz4QNIq53e3ze
OS/C1RMa4lNRv5MDYWVdKDd55FpGeMSWgaBV7TgXW2XnDaaPSXmEnhaK62qA0w3DC4IL/irg9OVn
3aAXu7ZK3b4z+qsQQBnW+hUiayCPcn9NNwzAIwEYiHfHz649U3Ou5I2aWLG5spyQZ/VSSpKQFV3n
ChjUIeLKiFfkdyWRoEerLQT9ZY8aJh5sAD1mtyWzvjD4SGD5sHO7PDj0R1iaSOhgTNOZptSDwRZD
SWIkrx8aAikB0K8vW/dJ9nEzvqLeauFB9n0yQtpqn0OS+lp3rVgTQYE/ffMgmEZe98PLddXVoVWJ
eC4+ezrrc4rZW8KUEJdQBnufu3j12ZOYQBF2WK5a77LCnYEZZCvmZ8LdCkPHTPC837uXcQUugV1D
Pd9UBu/kTUH7walwex5vgFZJh0UY/68lgeR2XTsTF0g9ubKstFPXRKRX/+QfJyPSA+aLlDFS8uqR
D8//xRfx9e7UYIFZkyM6BC6zwt7n8l1J5zSU4UfK9CrHpZ7pNNfUYgQxgWvJ1FnY0u+9EcIgdhda
Vq0m0QbqR4XXoSnrKxG8xEjUWoCJL/SurQrf25OXAbNtE2vFZEf32bwroiEi9aF5oJlV8agP+TeS
LWdwdOXAnKfzcZY8ksFdcUD8kmy48DDmeMH/x6cfsQu79kEtzj3gQ9jTo4fUoHF/sncb6gxT0rew
1lFNpTlNUbgXfAS5p8Gx5MGUUV4iarK//kxQpv+VkeI50hsAwbwrUv2C5PHpj8WTvYvskQmWisRE
iYZK+Lx6N1AWXNTW9okX6HrXO/oBlLtyufyBuwFnWiR8T4TjzOuIVqkZwcNaaLORdxFK/JY/1IwH
YmhvHn6o1NwywjaMzsmVa0h2a+czehdD1SPg8zriW9/rf7ZkZx/uU4Nvpu67FpwL+b05E76czN3p
cOJr4jFFoZQ3xV8CVIA7DSR5Q1MzRrLONKb4s5oJVLLujJHyLs+CnR/0mm8MWAAvZhmM5bHqoB82
LkdkyoNmbJUJkLK2RZWsUbxr/wUZxfvsVFLE1in2u0iPmn3a6cDvmD9BeBRnPtBrtqsL7lVGNMcR
7qqLXh5NamRRBhiOzZSHPc6Ib+WrQcG+hx9lgPrKL/7D3VfdJJhfk/C5Ir+wcNDJ2Tsk5yVbWDPU
jImRvFWrTBFvi7ytlOb/okZjDPTY6sjZ+yINfvqQHYJwZoO1QkHrrx+Ase+v6s+7mR6BuWOxhqLM
3M7DV9cXwJ450H5AIfyTJJsec+WOcEgK5tljajFvZyHpdt2OnKnpv2rTwJoKaOEVQqnurCdr1Cfr
a4ClnLIER1J9yLuLHuORKYuAl8ucoxDi/UIImJKWtiSAvGkK7UqjhdGQG8nbwSLsluRIJxOni7Fl
gzoeH56unlRDolhTPA2ny8tTM5QFe0JGuULgmvKrN0ZkMyTUbv77IhkcuWkhTcc1NsR3DqnIUXoV
/9dvRmmr6GhLkBtrWL4n2n0yvqPHiMgn6hSWznXZx8Tt31U0ZfIxWrJ1tI+snfLWWtFnJoGgxYlz
5/qw52h7lmaP8YgC8oHykMpQPhzqR7Dq3PTs0DB20cPF6YD49bp/EkZDBLR33pfs8e8mZ2BKg19x
umHIzHiqm7pq0+rZ49/asUqsOKmD63z7za1kEWuSZZsFFapYQHSvP0maT8jUAacslqmr93bpIWd6
uw8Dh2sXq/ktfTljv18J2jDWMiXbHiSdNw/yWW7CqTh1d6goCMvdVdCbnusKizJ+afXzephMrBB6
cwgElQDEkxbXbK8h/QJjK4UNOXX1VkcVASGNzcAy+5l5YVWcvW3Nq5VEw0bGCDMNFgMF6lCOeHNh
wWLkHsGlTMdniNaltv2sRBxgAPkHXIndYCatBkBMGdcm6EYU+EnSwNkniUEDv4/8NjDHg3i7uCSU
PFPtRrmhyuxpzuEM6qQ2lyAK7zNg24MEiovQF1gbnJ/p/Alr7RajnxSv729KSmhwI6WYyZPyXDKp
GdBljP72nMyXxiXn18dupA8w+PBcHaFeUjGH7bhOS5JRYEN6tSJKltVOhoxeFKPhEtflceNAg9PE
WeBb2+8oroMGRftzc1Dhc4ks2ZNV1fBjo7pfisYHLGUgHt5+OhmTI5ZaBrfGodNLGapefF86oRiz
BX9m0lOJHJFaDUOvVR5I90xXfx4s9hjZT8cLFTRLcE0AFPJXnxmi0kUtf0pprhNlrSkyVw73M202
/SJqrVQlHnsT7KzYYYj7z7Anwca0uWJ69CF+R5rX7TSnaGZoSNTcRDCx0QuqNZAVqeTBswUXPkmO
pfCbqcx0RL7/3051/Za/HrkblEQlnheC8TcEY5mKT+BtrjidwwXTxsK7/Gbv0Q0qzsrWA5xzIMkR
7MjMRw7nOqAPCDznbXFRqE8ES1rLJuRclWB91q6XiL9oiFsXYyuoyeAwLAwlCnEIA6Skoy9r9fdG
eIsKqSkxmltXGmTdtgBuDTIC3Nhl9P4L/BKQvAQfeXCsv+Pv+6GI9CdcHv8+4xuHCQ6xzHOJbsVP
hrUfbr2U2TKqmlzYYoTV5/02exSjqygZ2ekMRtub0Y8PK9yH3wiQIQr/KT9KhS3OR4gboRgTXMga
iWt2RtpXXm5YLU7XvvVQ+vCA0mtY6E3amvbjanBxABTiajui2VnqVWKXxyjA77eff4XixxIYGA0U
thmWDjh1mG/NHnvdwNP26BGzyOEw6DXyPYFuZAqkh/3nDt9Wu/F0ZULUarkXl42/sSRBIvQDy4g1
MYQOSCbQnszGM5qxLBHRVwaCicBzJslJDZIZ3talMZOcM3IPGPYBVGl0JK4tyxrM51SbU/QEs8Dj
GM27Ox120jtoSjFeVgJA5cstMr1LaFTh3LtVYA/le3pjY/m2Ga/5ySAyycR8aWuOvoFTMSZJIur9
OTHALTWT+lOdEPWA/P/AaVOX0XcesNqU3NYysNS2AqPFJHOzyLYfAl7yhkuBUbFx9g77D6cLyPOp
Imox4ZFi/4Hm4laRYLuOAqd46jE1xIHbQEP8iKdDz4UkHRWHe8lbErYXVxzqOuqZ1XhmUAQL178i
/hUge79k0wpbF3tqQoIwUozWr3O7602bMVIFaiQQj+0HhkG2IzTm2Yrl49Szrcp8h2LbvwL13RlC
azLfmyclNfZDM4SMmPo6tGOHrXPPKeEgdn3RcWxVk1AxK0DjCDh/y3kurAam3Au5Qe675oymrtTO
bPFM9z0xp5NFKoZCVu9o8+UNiZQ63yjpWwkPuBR70LNtIxh/GuY2gYTwOrxB5UtVGPVAFRI3+C71
4C9FuB/WM7H0IH+IEBZLmYvw/8TndVW36IpnXFssnt63sLfRFQ2A2ZrMNQvWMFV3i0FYAaqGdN0r
fFsyCDqYQvXF1gnSoSOFcB6pyD4l6NXqiRSz+XN2kIjUeLHh27Onf17SXaevld9AgSy4WOh//MBi
6vxCnFNh4cA9E4h2HcBy//RMk3X7MTJrf3zH3Z7KOCRHmNGnTvS1KgkkyVE/tJITmENIi3Ff39ub
IWiUY1iC68ELsSpUA2/MP0FLqMdDKlvadRUSeXo1mb1ffDjHIS2xmdfiSCy45b8bFzgMdufvHf7y
DnzEt9U2hDpctUkuSn3opU3iGTjaSFUYiEXoa/YUBeTV8qgyzGha5+WQIC3M1KyZeTPKdjWu70PM
DQSelL5wvKDXJMf+V9ZY9XxUYa0dvJd/bxPDWUhIh1OpPo1f156SYKBpRgIkXwo5Kk5rcuBcQ2+I
NhfSmhKrUbJ/mFCveyMt9SkNwhEy16wMYlYGL6iv6B9ntDEWg/MLD2i8+zynYHu0QB/XQ+qzkx8L
eer1Z8R/xaFWyydFuY5PVfFKkEG48yx6FrNsC5mPGYj96u8fIp+vr8SPoUAQb6Ci/qdtsHK2Fil3
GGOcL7S98+pzZYOEYmdhU1OifMFOk5x3E9+d8oEtoDsLmGYNas3v2zhAqRQd+fwmTmdc4feJZ5E3
mYk62qPaK1/8SACCDptxu9/RyY9T8VYEryk54g+4KQKnmh85+s3P9uBT5gjw+9LV3jZ00srGSX1X
TIbYYRbgfdRX9X+Ss1ajGd5r0LdmNm1D54zCSumh4zhp2aw9cDfKvCax/uNRTmsRp7f4KLCUZuN5
/rllHOXDLiU4FBqZX/p8wn8jtCGc/AU7UpwI6feaa1SsMZhwTCbgeOBQ8ohs2ywxEfZXGEzqeXBP
92U96WaxuHnP7SbCfc+lN2N3IhGDM3EcC85WN4eMgqYG7O6QO8I7sn2aQJk1+cis4wJsc8RokP0X
jKSFX2CFKlVnMa42ZS8hXAl++AqPOe9bIeodZ5CwzMMolgJ63tD9SEZSgr/B2Hx0A5oK3oE/c21h
Hx+vp8sss7WvlBLAM68R+jgHkVju0fvB0ZNSsrV+Xed/oteJeW0Hmf1AJ98UvaZlsNvNUX64+oqm
zSf5m1EuwWGHE8KNUs2rWo+jXkLDWp9WVEckyyJxzfZ45ZcdQ8TXzyICltz1Uk2TXwN3Lt0jf5v4
Mc9O3W7TxJfIm3T9D6IWf6/Y7piFdkUoi8or2PhmzeKZmKxSmHM+dum0nSEUFSOQUwq79OZqapoa
ej0j3kKoIuinnf1yPDL/jyBx3Ewzf4I/XllS1FKTVWKuHtLUgjJNsapfxusLLkT6UgdtBQy9UGE8
NrMuFBsB9SgZmTRvPbrvBEmiWBwCmDkk1RlpNhPKoJIiWA8YQosMUyDDSWwWU7FTRnoEihDGRgWt
X4SHm22jUA2UdybSxSxR5t5eGQc9iQ0RMqO2YUQlmWHMrhBvkQiRuYFRmXO2/gCNyWbLOgfpo6JO
KEvBDxIB6iE77/49omO4N65koZfJh6HiTJm5huv/zwXXMY2CUGJif35qVA9pBNyFMouivOxAsndQ
Q1N5x4AjZmbaEQ4tPHtofu8CMOO547b3tLsMd3dtDSQ66QWp9e17dUXY2wGKk1Y3odh+/YS/2DSh
brYe0JF2t+0Y6ysf/4kb7EaaX+CQmdn9iX/sy6mkz/A6uGCI6vr4RoYHL38zMIDrXNGsqfk+NNav
nboOpxdvNTN6nqqhQtkHGaQF7nFDXqf4QbqVWtjjwko4uhyze0VXB2Nia23Awmi/oCaR2ZzxupF7
ZnKLQFHBW/iy+be9rFx923iuCdS4tZVVBK87SgQBZ6vK6KwUdLIi6jdR8cgseR7ucFJdxJVi+ZwP
I1mBadWdJ34jxsYMMBSxUU+ZDciu7UuhEXUOuGPsmM8Y8joNMmPuCD0IQyiXyTZr0UzT+Io5uYOI
/m+M12rUxzRV+bjTXnYVrXdaqsAdZc+8WxzBK84tRUC83YYqSi1UDPC0QKa8FMDy6HutkE3/Hy8R
PRZ98SXmatDhrJPxKp4ysjOEU+yU+EPIv522FXkm77XiKJf1YnDxQTvu/v6B5M0JaG3N2RnCZoG7
+FQTBGqw4bXU8sdgAS+Z3JcEjPS7Qym1n/82EJLUPnpEFAGgbpDO+z9WxOfbMYdudh9t24k1LkTu
oIwgN2Z1Qczt4Xsq7WTQ2X92FVOgWa6Xy2ubqM3vkDCCjHF9y21ug2/SXUyKzgLTd7eycdtskryV
M5qvtDUIfNq1pkOIP8/UkVmT2fJZgLgj/vIhHnYwnUDs3ygn+BL3DTt08LB9ksLgRKuJE8mdACqu
V5eYPRDl0OP0whlKRA8qMBjA0DBaqiK0d1M7BavEAzz1DWQQ+z6wZNDMsZW6iy6YNVG46BhkmUFN
pb4HS2HK/6HHwDublNhyHszujmDRSfaBDgd2MScuWJAQn7kAOHb89SQh
`protect end_protected

