`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
NE/TPAheNKTGVLK1Jq6PBGm4y8cn9mtr9qqwU1XHtun+EIN9yGGadhR+kEqDeylJ5T4A1qG/m+Xp
O38T6E+1UQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jU9GgCGuMNz5Iie7XSQBxs7Fk7Cd4/rpHTrQftmu/g4iB0UlTrSrSHtw+iLaImkVpOoyXmpIj9T8
HveqgokD+3rF2YmlbHV2hs1FQo1yzWjdqSQnoDvM8ErD1IdqJowl90n051cMrsoJdTOnoe6PPklq
NfwVGWc3OoPmqcy0nQU=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cCa3JfqWCxYcpHQVbu0W2qsdW95BHKf64tjPZiqPO93O2Jc/B1qlFW5Pq1wr1Uq1mxeohm+hMqw4
+ozsDRpyZyztECBL3Y1XPtn9UccnPzrkmXk8mwX9+1Ac7OvdGi+IjK1NRZJPSSsJbVWif/vqVPeC
Y1FG2sKi0DdbTZiU9aA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zE/7Xn0KELPzIlv3aivoJkAEuix03l2xYHaqi1eYyNKKIcqO0RHZY4ejZ0koXxWLy9HpUNml5XDE
RfxMEV83rQ5wLdQHnbVdPPxr9L5b8286Mh0CnlHN9p9PSENnXKqtvQcZ/s3jIIslbn9srgpw5kxX
S8bTSq1G1IfxZb8y67clI7ILuHt0YkuJo5Q/NdMHf4DjdjrtwMcjTknchBIQBGy9VtqQrrKmPpih
m16MNcohom8rB1cyX+FGoetJiinmyYeE/n6CWyg8JLYwZgEB/oPOf8dCwGUNJPdKvJK0j5aYBm0z
Tz+3siK7kBDS2O+qhdn1zwO6Qdkw83cEmfwpPg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZPP1UdRI2C6Dub6sp/yncyOSUiN/zMD5kdUY+DABM+pKmsyDzboDF31rZVo7GEf7XC0OyUHtkYyZ
zEBfeukg0/SCpbws6ThUqCmCiTfWVmIIFTgiGING8jk27N0xpW6VjIbDBOy4lbvF/WUfY/Slb81+
yMR/kKlBSpdGbFs44oxkiZvOOrpUboSfWc3tTt6DvDK0MBjm41McQZHTcKNXgFyWnrU6dwiLbLZL
ZfPsqRdWHolJ59BGPXkFgWw6W9zGsFjgurkhvjMMkNY1wE9nWJXwALk/2+p3Q0vJWi2s0jj1uiif
p6KNbR+ljyk5bJE6LG3oaRgk8cRMgbqK2uNazg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZWzveu/poFKFlxbXughILx+N+c4wCTsvuA+dCRg2hnejRzmcmHb+4Jh5DlvKvcQ7p4GxFFdwrXug
ufiXwThjraWy85vr+Ne4l6+5ABpLSCv7YSU11hcxEZHjV/zAxB/CgLuOttR1r37yoB0PWWjZtSSa
NJNvrgtFrxfV5GVQdeiDllO4kdNcIULvdsEEhjKinIDlNiF3l5LsJbmplk/2ShayXlgEnqe8WbX5
iwAoDytOAY+1oZMeG6Hn1i7k0UspTuGaqcJfCy0PEimkYDV7ONj38MiXKINKD5wM0RI2lL777Snx
VrG/GqnwtfiUJge+2j1y0aF7x06bsEMa83mlGg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1558368)
`protect data_block
jkXLEaHWLnYQj0cPn/maEgcdU89tQMKps1cEGLKdtkCie8zbgmFMxfULQsT/YmMr5f0rhqsOlrfA
vwmYLOMhhmGhaWOp8PnhB98C8dcAhhvIxmkjootfcgk0WHY7GOwFDiXrX5oXFr+l4Y8g/mzYGA5B
YcSIAJmoIwVmm3YMDLFKLJxwomdLIh7h5Pve2Qd38jmfYHH/mSRVSRZePw0fcN0EPWFOkkwc1uur
suZ7XxMhXbfRdRjZ5jev3ZyCWH/qNron/KMWWNi/AXfz7Z5Y7rLSBX56nTtV7IWxR2mHQ6FxeytZ
IXLnlpDt6d+R7GNUrDGls4sBYX2DWQ8n4op0opPAqoZq23z7+iK2n83QjbwDh+zCvij9LISiQ1cF
kB94qdtC8fgroPC5RTCMu2d7ZA757R1J8JEi3Le3/2VYGi/cNI4khSEWPs1TCgmdpLLzXwlOp0wm
8FP1xMFMhyf4MTjIOorHiwqMwAIs0cuhZaM4SkHE/dPjOL6hp3X534UM+OxD8C8Ukz1j6BcHTjsk
YAT+IIfmKlywp2AFhHosYb3lQ558Um/Kt77D/72IpQAAPN+FtV12M9MSplPThWrLqMUv4KVX1iMi
j3R4kjEddShvLdcIU1uF+2LjR0M20fpzD6hmd5OpRjoyOddT81rNKuWfAXQLx8Xd9s7i1zNJV8KJ
sFSYk2hIYuaNIqWV69UAIQJEaJi0RCCVIDkZQ9igeZh5KnIxpAYctOjKm/nItJDMjoNjeEJsM3er
4qUSpT5b/D8llnzL152WfthwSTqm1y+k0bn1f035TwXKtACeP924Exo6zdNImRKPjM09MAyGX1Fo
gEPUHgrXweWLpedGKU22LpbksFUE78JvXzUjuBM/T/mtWJ3hNsimjYA6KE8YRDhcd6u6LEqI2eL8
OpKC+HOZQW03J2YCH6FEP7OQ46xSZ4LKPG6g9HDCDrz2xoyGkpW5eSCsymWlWv6hm5RNwPwgbeLE
z74IbaLG3kdtHMAK7ImmPwOXVkM4/x8lShcWHJY3QLwqA/QC8iwaRc60r047qGi4Q8lInf8lZGde
tGZIrz/ZA83WtF8lsUk3XtFFDyaMe1tW9CDDZxibZN6m9CgQwUle+Z2L4at4mvD7nI483rK18xvO
pKan6zkj/AsK95mhtbIDhPfpelyW6xExKtI7BtXbWS2gknCBHOwuxeCroMKknHBNGC617GJw/aM5
Qj5FI22BDMsRCfBUyJfqY2fYV46At3sauwriXJ7nLj+UaO5gxSow1RCzGCHtvjWVmCEymeQmijSg
d68cFeHym/6VaVU1InsybmlAVoX94JRC5fUKeKUVGdNr+Cf2QI+fSyzTu/B2pYkn8V0VmUFTrPUO
4uK6fgunFjR296zEp+Z9MUN6ZjSvCQHJdjv1SBbpvTqC7ydm5Vio6JYhIWOKqOOJ9oNiKOx7+56W
p1PxFURyBnHol7P37/m3Cy8+UlLrEC/mZva6ngprcmF/jh/3bca9rTNpwEfr9ON3ev7upcuocy55
zV60v4MOMq96v+WWTkr4/nO6b4P0FaUv79kk+cQ5TcU+TX25Y7hIcOFfhAkhyYQRmSmPv2Wf6xUN
bvCUqWtzD/T9gWawSp8HpdJGNdxrPViZ+CG6T5JsyeTMeMo/BU/brB7ZO1HBqzV1QZVJs7K0ysU0
qjhRqToyi/wy96A/n8+cYDBYDK7xV3eLTBpVOOXdqF1Tx5AkjZNdWCwR+cJnGN4Y9jrJXhJAWckb
Njtaehd7T3KUSZ4DioMYuCEQSqDokVeo1stbij7740nsw+P+TVfLHYwtO2nH0kQiI1/9esQufH/R
5NCUJmIgGIpcup1hRBUL57brLtyJEHrRM+SouUvHgwQD6G6eLg30NBTluwwe0cIY1qYo0TWWpAbx
6QHDFG0ThB9WnPvSegIiaZEE6Wv3ICt6RnqEzt4/uOi8sbVur8ZTvsyn9tbyI7LUzPadqb2TL6uC
Gmw72B4nTzFRh0Abm3ZwRRgVGc+HpU+xSzU5H5vOjjLrAonq6jyxP5MwvDTjP9iIBANr8DH1BCXT
9s1dLP1opEB/06QQv98WwYV1UIiN0Y7Is+T4r1igabw/w0gErfLf/Li4w51eyMHugg5XTZsVz3QU
U6Zn6+uXQmE8dcYREeVSM5PYDmN9qQFPCSGp5S2Snga5Vaj+6FmVdQuGWoT1X1KlfT9Ohyxfgen5
CzgwG6nJiMEwgpI9ipXt5X/MVvY4hsExYWv0F7lpanrKyGeUcM4/kPbSUlt9Wf4dAsqg5MlpXuBd
w7NTUcQvIFr14ZGzhUVmTw5MWAVZ6XwdhNWgmIrHHnOogxNodqV+Rsq8Yqh7aQ8H8UhYNZQdFips
RvQ0L/CCgj3OcsoUTXHCNs95bNfx0nEE/bzf+z1GiT87gOW3Ic6BN22Sakl3fPQg9X8rie1Y35pW
5wL9A5XkonNaGTNU26wkOc3pjTqMTEJl8Bp7qyIGAe57bLH2oAJ7xsNhBJ9sOcLNYH5fT6ghqT3P
7+ekri4fTY01RlT2rCfbu83JeCF3+Vkk6qb1rHwaoB1qnuRps5jZ3OEhlONAV7MeJqWi01nCYY87
pxjD81tX+Brx2kLhjWUe8e+hTlakJ5eraDOi8DaR8pe5YrLzupmmY/hkUpsDvDXkMFPjUfy5uzvb
1PswMcLGFeTV0McpiZ59sO2fWwZjdcU/RaL4Jen01ZnKzSzTVA7De4ZnRFntujuPvYp/zHs+Eqsd
wxmCaSSGlRclIBwmG4JtPtVx7YQrOjuYw+fe26B7Akgkpe48RDItxzchsY1HnmJmr+WRHXnkGsyq
3Ldjt2UrM9+m/WlCAsXqxA7ZkttQookRC7RyArEkopDYWk6anhdctBEEvZBXOAGVB+psuQ2hnv4o
aF3rgTaiFvSt1BJnF9SZana65gZjTxYLQMG9mEdJXbimPj1bCTtIhTcoBsBqi30b4+VP7TDi0/UO
Py4el75MooUi43WykY3TsXe2oupCdNoj0GXEdQy+pybkXgclOHrHy91uUT/G/cwW2Xv5AGIRLK7Q
eW3gj8h0Q1PzcxzXhSR6QZ62DJVeYZaUQZamNxMvzkDPTmZwKr7N7RRe/gF62FQSImZvlDSzwStF
/FUVTb+JZA/MwhwWZOYRZum0HPkFIc8dKZcq8GUC1gO5beaQaN9stOVT4BCKJGqKrAgkqqHIVJgg
5MKFizFL+FiQuAQFQ2oQ/2J+LTn7D4H05iXEbuOf0lUODSawxjInz4F9Fk8f/MgkWhDkaNBpeUPx
1Gm3rUoNDpncbvPaRW/i469J8or3GtUkCwZKQy7+oRyb+azijV0cYClmI5B4xTP6bbfhh1jkHryr
aED89MjJJ0lbGVGDDTC+9ykEa4gyrOe7O/UhmH/HYgsglKghvM3S6Mnf9sGcZiRKrBr8d+cBA0Xz
8F6zHRddCGHq9To3zk4owqG/QPpwPCdGKGDuwslEdLJoUD9b5J5Yl9FPlYy9kyR1vn5nP3zCZpw8
MU1a3Rcdrc4St8fwpR7uNWBiRC0lwwbc4k5fqrcn8kKRGx1w2aI3iX2i+zaVN0bDmeMnCtRYMXi2
KShxSNQX2Te5R8r/As8Dcp1a5ry732invyFIkyBn5s+imHZ83HxgG84OU3MVSr78TyiN6jGXI5qn
AWwS4qjEfP6AFnAMrdDz53YIyfZgQTiiYO+m7k4QwR94Pc7OzY4lWDifAsadHGT3XBrFpShGT3Y1
golpoDSh1WAyBPWBASv9rqlNsTnyFjLtgeJKWnDCQH3E6yzTifAOasY+Ig+N6OW0f/jkKkcZuJJd
hRNmWaGZW3YtLEY1wCdnhdjQfi8jKom4XNS4+srd2ar+u1rDbCyW5h2NdDwausLbb7y7S0ar6gVK
wQ2g+vpqqsH515jtECsnXrTMfo8drZeCHkBVmLxqYqzDzBV0BnfnTdWLa8aM/nHs6g2PRANp8w/2
HTYnwoXZv6WpymQwuwpJxJcONCzAVVJTzDKN8E33eTCieBh7wi2NgBwwxytICoe6HxXA0U7l5TUB
BhXEPKkxsbVtjJXOVKiSD2FrmbWA2k9hO71sLJcv0GZFwJ+JBBkjE9NfuETIsSsWlZqgoXEfHWwE
7yCwsA6tSbm+TT2N551B0ClCZzGdoqjlYGF2N+kZ9ip6VVv5FEv59oDaPn1t2KlUYbuaKW5pEFSh
b7YlhEJF3wvc6uhyRRH8RqTLZB5EjAmEouYjsz5VWMoWuODrGMQAoQGgkBRaaIo5xLehqTs9CVwc
/6NWjIwHiwCbYyx33Tpn+RlA9zxl5rvrzQd3jz1L+0K7XaoG/npOoUWgcp57BZYexu9P7iCF5SxF
moeUv1TAYDTZvfg0sH32Gb5sPmFKyJw2hPwj/799Wq4R+mZewmvaET/aSE7A0GpV7ICwLeM+qVrl
QOAfdMi4MP/EYjysWiJNfzKANQqQaamLZsg2wySlbrKnPH5fx5ZDlPSixx6vDYUbN9kDoH2sM3Rs
WfuLkoaH8+g7EbLDDaRr8g6J++45O6g1CD46HgEcfGe9C2jEqoLKub2DNEnZU3UtN0Di1dUKjKlv
D2cDG455SPhndm5/efd/EY+W4lDLebcLVAZuFmH1HUDBwPDLhabXgfb3lmUJnx0LOBkxe1cBly9w
qA87K/HLeZ1LcPd4kDpb2q5LN0gmDYfJqD5dzvrGi1zs5quUytwRgunabufy401hIMzfpjZmcKDp
QRM7zRLRByi4jt1XADK083SCMpnBsWPFnCuBZlQ0p0z7Vln+5ZjdhqPa+vWmqYpOvdfiGXKXUT19
sahfpcSXhh8aqSd+plukg9XlV0c/3IF+u/bYVU6SupJoJqBakeSuSZ6OtBTFsDXLJB0cjBY2L44v
M62/Xi6ENRXFZLTN02RhInIbHZHPEd19YSdQksj7vdnvndLKZyODJxFB4KY+hUHGBbxHX0ryx5ZU
NRN2+bT23srRscl9868pPHfF7SoGMWhbLgfEpPtQIwkmDqQRsrfTOLTmJtuzxZ8UrN+cwp8C7ZKs
gAlcs2+TmtI6i7TwB9qmErNyWWdDUpfWl+Gne5lV+CSDqiNMW0oRqswUPOTx4GPDaHLfXnh0qJBW
2SGJ8aQwduUMv7pnIkFrEBlDuT3Wwg6vyuQVrYRJ1rtM+hbuYwQKGSAZrbRlR5ewCpOFs/nxXvfm
LJ+nvcqC+ZLPp8WtpwBt/dgkKjT/n1/JecBEOyDaaHo83d/QEt9OLt4EqMtJsHIzLnJugMblimro
9NyDqp8/NXGz/lGQWngr7MeY2ZVGgqscVhW8S5F18H0XEUUk+gH418fWZ0RqAXiTa96D6usyqLYB
lfiMLvdVEybz7Zh7EegPktG3MdHIKFNv+HoLlSyp13EJooNXaRyakcsrAUYla4burZQkS3EjKfJc
m5TmIsTk9l4sYe/S/Dm4zbTpIG6IWXOMVZNTpGdnGhbCN2eCYIx4KPviRbqBlyTUnRzwMEoace5r
lwUAJOJdgTz2S3CFHzusquTwibIBJ89PN12ZvF5+pYTv5QxDVnW/h1qme6+cjnhKoDcfsqoB5mdK
J5C20zq1R33R+cpfj3igy+55qdTmIlV/6VhCytCzOWFW2JC329saP7qLqjHzJq7Dhwc1BMFXHUJ1
bhCMs7vBVXLITVzRnVCrTdDK55GTuqj312i2X8PHd0jTmgzt3NpZu8o0hHbm1slBdHpRv9OAeJZV
zkz/otvt1t9qUmTnO8K7Ld2ePp+aEc7TguiKYAFJfbFsSbGUIkQF2QHFtlA2+PLI9mcx0j0fwtMa
r4B/omr0pITrB1SWTab2GkYaT77aJlL+t5FzzbI8wLT5ClpUi2AeoJgKJggc+weH9OeFipC1ONYf
pZ/S6S0EqF2Ptdcxomo8d7YjltO85Iijg02IyFmtnZdeEJs3qJ1WjgBCGG2LEEyN0bHHGg2m5mVF
rpHvQ/siZVuvwaqpB/+HBrUWdsLURdF/7+6IQQD8yxatt8uKbTuVbUd7hHAd2bZYrKIMim4t2GGJ
8nBLjqXhfMwETapAkgNEv2Qx0uCjU+gNbAAV6nIq7GxWfuAqAmvOrHHs/3RXjfLWmtXF7c/DErsH
UG+vJaDc7Ni7hqxrUK6oE1tSShAO+r1JuElUgz2XfbIzm+S1gQMbB2rxSzPfNBFtJFZK4toNChDx
cf/1Vc5DmwwxjqZvAoDGYO8bO+GRcncBEhBjlCvDMXRf3a8NVcaE3GXGtcr9G3qqH7qwfpk9h7fJ
t2zzIVE1l+1MqQpgPJoX7mXxHvUy0Y0kJHQ72o9foI8FJquXetIbT3jDelz0PPw1Hl36IjhK0f5Y
qJnzADcPTh7BJfxRZ1ONmxRe+yFWhM9ZmO+dmP/EAy6sWcvdNLy2b3jwHRRIcIgONey7zJQhfUOx
TLxALCkPfgbhXge4lgEmz+w7OgbkFRZwFl3K3wnIe/IZUyu7AUJG8ac4R9jyFZhCpIDyzDmmBPnr
Oy9Ya+vXDVZYPKIz9Zsx1jgY5uvTcsGsrJ913Djd3DxrnsjtbJKmX9+9x0fXstdKUzm8H9t4okfB
dAp/gsX31japSr5EdeqH9fiKoXqRZQFETq3Kyty9DKTYFuCrQOsjhA/SB/8HIWCp3Jf7H3/odIfX
znSvLV9xfuo6nQ75C7rOoE+HcETWMIOLpWzLxz6rsZVWEi7ylP0/we7BuvmuIpot/q2dt+AYwQCh
7yZNet0FIOzKaweYgdXRfMuMvLtymZDb0ThIoosBu4mEsGS6Hz+fScKdlqtavELpyR+0zpXDC9bC
HpuR6+/HctBKcTzliBtk7dfm/UFTekO9AnSWaJ2IqkFxEr0Icg8FGPFY2OTH5ntpphMV9yS0ktKd
2/VICmI9IreSfsOnXvbrBte3PJWjIsgoVcorvqEqNG4loU2COHKzLOcTCUcye2Cl7QKsE+6pdaBt
XxhxQZJqJy6YNBSqda9Yf9ae5I+IDO5gKqUNtna6WLVG8Avg3A/ZNkWfwBYYsWS95AbHj+jdqBZm
Kk4mjH6ATPwVowCPzrIhnEEDQUzJ1kPnE5bWBtIWKyBnKWbRFEzfGyHFDssRYzBwbHZZ3L1oRRzC
QRYE4j/V/aPFcaNYIDkKBfcDQyU8rqaaG65xf+Fhvkkx/1NUypseMWL2W4/PUjKhaxOHvhEhy6vl
VuZVC+fPjvw+hcekcTydGlWJuzwtybdMqjM/F0hmhQoX5qayBfvy1VaA5RNBTgC8wo0wN75ibv//
BLx7gnImm5h8kTEy4OrYfWv4ROsm7SD8esUzLeGoKmfBXVGZStjBuI72do1SqWi3zLRt1FsHyP7D
wZJ9m6YZGmmwSBoETe40SqBbDZBW01BNZKJEHZYrtQr7ImQgMdAaTojeNcmtTb/U2lIHgJti+MzQ
ihsHG1oTWn2vr7FpmIhTnaWiMw8K1EX/hVAc3LUpP6zfvmBHTrZzbo1bjyxCi1Gw+vc4D2nGcKKt
rEEEaSM7iGIwNSpo5WOT8MciKR4f1BVjA5+7JznCzucYREbh7RtQHQP4mX1SQanCeC6YEtTEBI68
rinLV3Cqrz4K594HaERB11ev+urBLZGIimPMAC4F8n1Cs8nJRoJFlFBT8GB2RUhDCn4FuXMt2l3+
0BTad0ZLZRrZj6Wauu9NcYb2MjFgfnrxvRAizHdb4Z/f41c7Tuzwwdg2Us1zId9yzlohvhCmAETN
WWwlhOpa/ZCgfbV502WqA/2hOmExn9ppYTbqPenHzVclw4pqBZsqfKSfd989eADmU26jV4Z/I71Q
W9FcjVUy0MvuPe3QbYqJHxIuPWL4Ev1dCbwlZyEaiyMf5vr7Y+8A7Hz1HFluGwQBCi7T1EZHrgSh
YNFa5u8YgE2FvXbum+kAjBuU1gHqDjd68bemNYpb9ggGU7kuYEZXs4FfF8fdWdUZ+36SUHjVvIzl
Cp2fpPuxOJlPNCWf2bpxwDtGwEndN0VZrIxNoVr9FIql4Ur+OVcKILX63/YAkt9hhfUJUa4ppo5i
LjbFGhoKowSJnfJHuk/yrRpo9vmg9aBruatrprX9msOa26seOy21C2oOXZoAHAPZiQxOJ1Jh/sAy
BvhhT1ZMtWEd1PgNKdLooKLPHVbmr4lhZmACxZmPV7mXtUMa43DHwZy/fHqH8g1vUCZHOGmQGESz
7uLIn42TW+XB/aQUgFgWieSZDJHXOrTapbZ/ZBRk5RotOoKsbx+nEPNKQr0vSeXcvapUWNkVn3kQ
sANJP1oiEkZddMzb0RwM94JrDx9is8XbzBvrivxHEL+BuGUlcjHfTqmdxi8a04OBZ7DwwZ5wCto8
NB6sloO/cihnVg7QGP3sNElpPag48796WaVgOu/Xa8j46vRWGgpFAJl3dVDdGyrbt3XiZiiX5MqK
Gf/sckxH780n4GdHmwFJIcnhbI1FixRv68DjC7pWBLxP+g/GCDD5KNF2A6x3hoQ8VARJhWgeFfjw
ybtijcC6pos0qlxCeLqek4AJpDzWxHevQt41mNaoc+DemX+O0g/TZNTS2zDANTn5rJqJePlR2Rvl
ZLu1KuvjZgoF/GpuX+kLtrWSQjNjEnetnRtWByd7PZWtvi3nF11Hg1jHT/LHxxbl90I8lcIwQGFp
UHXaQw48lNMR9orGD2khyxJzzme0cwKVK5ADzbNEdxYQ5bBrb3+Y1W6W6V21RKrvyRZHrugqfdz9
e2P9tI8uFG7o63Ha6xq+DiEDlH7iAkzMmaQQs4XF3IoLOi7ubDxDbSqG+9Q6aALnpzU1cnRIYgNI
Vqi+QV13dxhoVmrgUNTNbvgCMjDq4Ey4eP6OoYrhISJVDaQy4jiB9T7Lpjuh43lkHwVbT/UHcjXw
XhFyh6X01ipDocCQkPrkd3pshvxuBVgtV/U4D35hiGElD1jsYzYhU/kAIpzvL3xU3S3ID0qSY3NW
kZ+PeDNlTi+JzaI/85EnZBjB6hbSk9DnCl1w6ckVI2QPDLbC/a2Lh/m3LBC0pUDPIZ77N347dEoy
x1jFfJ8pry4vlSchKLgEVX6ESUhGzUXkQhk75xCfx8MaYNXQNGdIOTaxQH9osLMkOt7KljmMcVTJ
wecl8ttBBs15V9HcrAULEuiPkVV8ShgQ7FmT+oTSmPYR81irK6LhGHnaT4XMmHDIB66fi6Cm9msG
o75lJ718GWC/qieW+wreNztyD/5HZFzbTONd6DaAnQ6WWB9w/YVj4AIoNMuLmagI6CxYCJrWDh9J
oUkHrC4ZhvolAoB5iKqzoJY2KVz9khZD3DoL17bUEiYTw0HHj4KwOLt2tx9kkGseI9/S5i3AArHt
lYlBRiUl2dVylp92K2sWrwWvsT/e5+p4XHs3k3Pr/Arvw4b4tvXDxdVK6dwZcYo4kYsUrwcfLmcT
vAYrSLvFX4pFZXyxbj+9KXoGg7qX8C5id2ueDygWVvjn96IKAtVx8+OF0TKN720rxBla46cEZ7oP
JsFXwAGoczbXnb3fHQjevTO37m/ZSm1qbkpGv61LZXDW8xclsCoXuSyjFEACSj1kDh2fzgfrVsQK
7TbI8uOZG54ekq/AHFtHZ7sFeOwydtktsrdI/F+SyDmmFeDQL0M73UZ3p37UxBtx/m9p9YpDOZ/j
B21AUWnTe8TWjSv7A1AnhfvZTPAuTeEi9ow0yuH1/2UmwOiCQnuA62dCDyPtkOg9rFIZNacvnaVv
5GrB7X1cTHvbswjcd+7PrMrkiONf5AdP+B4yZa59OF4kQDDygPsmG+1RRoAABGjWcUtsxn0pTi+E
YvFig4BZrzUcq7gisaNjY+/3FYy02m3p5Lggk/LB/nOjCqzy3QyZ3lszJbYujAWYfXB8qaDH6jUH
tBZ0gGgMHjoe9+pR8ZL+ffdXI1VqmcIJgeHeoFqnFYcD7wJSVnr4JMnbBtjBzw4pxtC4UXJHjbxC
SaW9ozWmn6jdbHB4A0Sktf+pSI0I66wAbvss1a6X+O6OiHIuW/MQnq3IlCG3uwqkpx9uc0o1pUxI
AdF92ZBWhkn6r+WA44cBQrA5LGyU1pQZXg8N3VXrCEy5TkzfW//xN3ecopfqc60YRwlm2734GdVc
dwxHqrbEXTjhc439tJvrNoYElQKXIp7yAo9c11jvlI3+wvs91TjXAytkrw7oaMeClbjXvX3ZjmBg
F48IvJ6n0L22KX4WzOl9Ui+R4lZ+L6jSVCS0gvuCNmqvEDddBZ44dDilVqVvItRDFwKkhQeq8DvX
k5wBHyQYoWMCoIlYjJfEOrSIg6yOJRbRrsmo8B3kyKBjxrp0jgf8/Dx9JJ7Tg/byFhKXSPsWKIAd
KxuReHbgluMAewghdg70nrYM8ClTJytoH4JWUz8Z/rz752Jbo1rAcVkH8QcZ+BAFGIufhNK3W3lG
PgjDhG18K+LdZc+lhVsAq8iTUSA86AocstoLiIhxloD3lN7cEr5/tSy3Pguh5xID4LZAADv/dAY+
Q4QppT6jLh7sUNfQ51Kcx0YRbIweHehiLs8L03e54sWk82WPOAosTG02MLQIyVhf1cE+T/M7MK5I
TKzJJ2T9/VVt+72G2hjMDdIk3DUek9zLgNsxDk967h76K6gq/n8nbeZOZMSngLwUcmCuVgmPKpcI
N1a0DzGUvIOd85D60oMKttnn6NtZUhnKHSI5Urkzy1aBZ0XYAF2TWW95es7YfZSq8kQN7v8RBod6
wp9HVUN42TqHCJFIwtkWPj7HpJ93rCIJyV3s4sdhx/YmWd2mRl01l/LDtvAOusUV9NWNQFciJM2P
JFu8rCZCHHdbMu4nDmCU3E4hQvtaTgQuQ2erR7sUW+5QcECI59uHSIOlnDJ9K7ixrH1cmNPrhjIr
oyB3uEtt4mWmAdbu+VIORGMFMRdotxPodpTx7YwxMKnJbMsGfJjS+ltEHM7/S7wetnSiBHptmAjU
160t4SP9zsLy4Ec9MOEk9GaBsYB1zY/jbk8sJfuaXFPe4NgSqifKslEoorCFvJwC5pAjKENX8U1Q
/bYoK6t6RYhJ+v9r7UqrM3+g+Js/XrJIUP8CXWEcvTwZxY9DZI6H+i7Q54z0JxVkZ0vyrqETwe4e
N0UI92BxWJOMdC9wIZ8do2aSSUhqH4G82l5blNuQAZdHyIYrlUboTAX49COr9/vtubBx0GEyHBvT
rZ3uwpxIScqHzoMWOOq3REHBZQxkC/O9HuU/Iq8+oFRXSud4DrXGysl9tQrtowd5iv1dL8ofambZ
C/jDxQH3qxXj+MbICjbrFudwKGuhEgRosxOrER2BMwqrYtNSELfETW4vo3j/lw9Zgf2rz9YJ9Mr3
vopS2urIyr/kS2QFOUdKhBVB3xjmmU6LFzp6GcXb7uGnOhi918tLpOzEX4ShmdywYEAs2yYyG7xZ
5PqP0sV5Zq+O0LPgh1HcGtTd/vImpq9uLXjkId2XROYWFeOQHdoqF3dDikyZtndjpQUqgn88bq0R
g04w86wdIxopUwsLr+rYrS/SzRlsWrTE0uuaW+7+S4NzO62lDAcWd2giTqLawJsKxKgG62xaqt3i
MRRv+gM9mKll0NtY9bAo9eA3ZCAF46hH+hElRLtO+7mw1OyzWK6Tb7L+kOcnhwMTgT+cIUDRLQ2f
1kRDyotB9DwZdICjC5+DXBAWQSk1x1ToZ/ZK4DIFefC8cLHPCTLy9DmFYmC3QjcvFSbPF46Zc8WH
gBkqvP5WTsC0okpfRaGqipJ5FrEhIYACO3E7vsT2JZ2umb0dMqOnrQJKzR5OID/OOX3to4t+JkgR
Aw/gGlMpmSj+KD9VOgrN5/VNynQIA8MTdpRZ8cWhEzy8hCjqzz0x330YtGDatcsVN5mUkRmu4O9V
6XK4/kuCOYvSi3auGCq6b+xu0BlDap64236uPCBppyQE33epDEzpiEnGhr6JVCJpUutaFx2lbJLN
jxLoUPbYHP4ljauFE/Y9JbCW8nZ4JYPYiAlpkfZm1Lk+R4ipV3mo//vqn1Y/T2VaJoeMEWqB2DCH
xxEoMMbFIgSDoX0CnT9yWby7gFIxMfr38bjMP2/aL7Ur8XInY3kYgx0SBFpfzjI+tSAnG9ok83G4
JOQ1Wcdc+MMxG7cOuWK+Xc+Gd0RbhnADV1NNVw6TIT5NGsffmsk0bDXJEi8YPoE+M9MuHVhbxgu8
lx9YQMB48/ZyrRxtTzApmrsCygLaufZq63MG0oXS7G9MwlNtmpf/ArxILe+pE6/1QznjVFBNdqFq
95X7SnKiQ+JQdgbRlgUiQHysDjpEbhYYjsKSXWltCyEAbWSyWRaJ3xVXteQKRofl8Yh4uegTIVKt
z2oTOEZsz+GdcGTHxTWZanNPkMKmvsF63105wp4WreAkgUfiC5iwtarqRcXXm8quJfJhrNpcrcye
ppiVZ9UVzSyvDOn6CKwZIgGXWdQi0ytZAf24bpT1ctQFt2WEBPMudAiKQKxukcowuKzbrVBlLiVE
5S7XcdGWhao49YyrxHZHUKCu1OKUYTEKOZy4SexdR/QUvxCCD7wZUnn5cWwmzjR5QFm05TLPtmV5
84spJHkrF+1/4cljeA09W/92cIZZMkfePjAsRyloWjk4PSZK3KF7XMLlgOBsPtD1uO19tpOsf45w
rN4z9xZjj3VjCZEiYXKf4+xvBGhn67spq3+m+aE65cGaEzL1gMDLFgPihoSN2rnYU0FnOs3DIEMd
fJrLr7/EpMQbI0wacRpEQhJej4t6Y3s8U9KmYOYAOeBEWQ6aTSd7V3p3ms1LRAqmQrlyTIroq1/j
ePUHdJUapCR4svOyo2b1r7E1bUyzJtiGpiefzfNDfcuE2EO/UgJdyyulwQbzO50TpuTTuHQB50aG
qFI2GG5OOq6PmCJGvaDZhDUAUQL8pVGlBLwFfXlV4iXIBlEKV33lpRv7G/tzYGs4wiUW+qZOJLae
7rlmnsWrV+OZ0hjh2LApPlypPOaTBmBfYZ5p95OD/bSMnUTM2B53U/j+2EvQaKXstC27b9/17kjW
xDiLmk/6f6moB5oXGz9uQBCSYSg/0wzgZgUcJ611c7fL3K28vCrd8RkJ4cyra4CP1+w0JGEiA5sr
q0Vj7ITgIPpXtWw01ZR1AxVXhTsSdFKwshRBLQnnasWLw/wJDmeIQj2LE5NDes78TlP2MFwUpolH
hQRcogr5w7OctM4aL2PwI44ndkFnFAZJrrEFZ8qKQZ55O2X9WD90hJXU6AVH//Tpb/rUeoyc4ECT
tzrlL+LU4x49k81MQCAGeKfjj3VVNkKROrxZy3Y3suJ5yrwka9UttVKMkE9viCKjdvagFgjYKz6T
awKXVmZ6D4r8LSqC1N3HJN4CWiZMQZ7llJKW+uhQ+PT2kZURixqbs9g+DWpejGYBUt8Ul+l0gIAe
pHxR9OslO0UHtKOEp1mRVgX+4ovULCFX22iTVmv5r//YISUUORLKNNnnTWJWe13M4QbauaHlYIwh
KhUpSRZLFt9vwliCoG8W0f5zd5QRlWs4meYGwaOyweSYYYNv2R/sPSrsUu0DjC/Ji9B8XDADmjQm
XnjNakyY/h3U09Zwfa9BY8bX6ZiYCZzRuFw5FuUPut8hwTuDkCHfLdZy9vZblr46hTN0tCjHTZNO
wy75RjbTuzx2RZYVU22QLyJKoCGIRkExlAaqWOAEcGFYu0GUq3RgQ/TQ85TIpEXlKzRzlEDRMJnU
rad/u2bxuDermKn0MY5VqX9+2k2c5lyM7I5v+Ix5WmebMpoQbBs7vh2j0kXmOOElB+F+F+1m+SnN
06rmR/2Wo2QLQMTx2wycs2+D6uSiX3JHq/LR0iCGqTQtce/0mkwLWbN6DXjUeOH6knDTdVR2UYVT
isbXPXp3ZiK5IoNExlRY5pALVTeFaxdrA4S/yU5JgzYnCrTmb0ikw4Q8s/qaVpYY879fcCpT2Ptu
Q///0AVH7zcLN0Ami48Aq40ysui199hWumAI0YJdwPacRY30IgudzlbxspTJPZP5n2piYg1kChX5
x/ryQtPaCdHXDJ4xkzH6GF3I4G/Hxz/2pVoB+1ijOiCysrBc1PZDwbG1t6Y0FdG97W20a6ZaXnUQ
Zc6YC06h68Uj7PID9Hca9zV6gQgh/UoGz2zF2NBwckk/zXqo4FpmvX3hPuhv8LDJPBrj5LgdhN8C
6ymfiiHw1ki8bPNEq+hg6Fx1XkOw7cwtjP33j3JZjRHITyeP2oYB9kG3a1naVBRAfkw1VibVqHob
3vP6hrjxDHDeuu+VOPJ8K3HDR6uwGnxfFGTVzXcYZ9CU34Kqv2YrvzEie4bh0NotxjmqQ2wVgJoQ
RzqKgB7utzciV/fO1JLyoME0L2wf0sSFHqCycc3Hm0RXp5gsR6JqvQWsP7ATghcMDOm5ZN0U0AtG
l+ntsRodPmPI+4l1ZnxznwQHFn5rBrX+U1waVxDrdKQytc1PjXcbktA94ymYzEfixj3NjbYWAAM1
H5ggAmHa75hqpj0olAORTzl3lB+jEIQ5OePYFTOVPnuTEz3sX73rRIALRwluoJ8QRwNXGCsP7JUm
sI7t2RPYPsrjFTMBwAgkyzY/PoHDpcp2tvPC+AJebqIK29/b5bl4yBDiXLIZyu2nBtJpGswZTTtC
BY2GUURy5jVpt5+ugNP0FFnNxCqoGqgx79HvqdZVFfEOHgzvL8DiP/Q4O4O2BhCHa9XgKG/IrbRk
enLiNxPXR3bTz4Xw5TAzKLV7HAfwlwUNC6JDtdfSO8MyXMacyx6f/0IXmluddy2ghyH4CBp0mFoq
ANcNddm2y766sZD/blY81BWXKTisNcu17Q2pwTQp8HxYxYpyFssGqUPi1ZPu6w+O1uC/6uLbgdK5
oxL+LEVSUz+drn3jR99J29zuO9T3uGStgTWR98tUYUfN0aItu+PgiiErXvInS9krUBWiNa9F2VR9
fgSbp+hrcXk18Wk2VYD2eQxS62o59RdeuBdv/3a7UBHrgTTBjkVEQ0MBvd7VK6TOqk2IgVh2VZtp
BOg1wV9KLc/FP4pmmBBXpmJooeyzygHwAAcAkcEPJGZRZfVntQnqsasDtUSG1SLdF+S7421Qexnp
9SPcKMCR9WeJ1AtHAzh4k6T7TPwwuTzrTWrFhS+8nKGloO3onA8dMj/e/xgkRBv47mVWyC3aATXz
aJTTJTrirnteS8YU8FAtV6J7EUmmQmB0W59URLYdejFNhzxkzfYgcG2YKSORxH1LhBO1pp1n7aWL
XtwDTifik0xYUFQogmyvh9vSZdpT2Ur6N8ueCRCdDg0FLyEfVW0kBfSVtDPNluXKJvcscuaZKrLE
UU+ddAXTM4ACidjVQPecH4t5JspEx4z+meeCi/dmGps7h7XElBZTSHX10whOHwW+zcotA57CXyt+
GIt8iy9G5qFBEIOI7pDoG0ICgcrYQmyZp5hmoSyKByqgyT7lW4BxhIAhwBKIjJltUvRBi0XkP37J
paO7BdIzdY6W3nXMXPJRsbsItpnl+HyBenvNrwIfA06N8v6/UmDSB1K/ycHewVNUF6X2P0iSg4u4
tNj5DXBgIqkJdQkhN9rzgtbYXIKpyYb0z52Gu18Lga5snUS1gaPqy5MNfaGzzh+LkKpgTQ3ZWZ3N
afbN3to8MSlP1MEzAoqg6JV3TByPBREz5HVIcwp+4RTAuUgsEff8uP6/MKv+eRXcIPR3camgtQa7
UGbnERcuzgIi7OebLIXV7gmZ3CEizuNIY66RyZPUmdzYOPhz54j/k57g74B1a4kdQZtHxrGVaFvH
8epNwo+jSPvz53+7yJok6kM8cE7NCIdiJGmK9yAKAvb/IwbPynuHgSpK+uoke2L5WFzQqhrcKbqX
gJ2ECuxQ9LMjSzuGRdf1nbDMazgcJySRGIWyD0KL+zdGkNr4cQrZwj4MCrckK34veCEfprt84nmC
xJ6M40N0csdNOzS6RHRvUA8mGdwmKF7GphiwcCg6rd3DrMrOXNJ2NzcPgeZ02QyxB6a2KjL9RATa
cuVAZISs6yanCbmNlBd1QAH3aSwMWb8WkZ62M7O8CwgSln1LiGgn67lRi1vwHUkNzkvHD1jw0AQR
y9Tuvxg8lM96qG2OV8kHUHG5CmZraDNG7NJSctAiAkL52/GlD8uff/dudQCXbpXRh5GapnwYLoR3
eqhRdGsgjPTiNDAUSdeNSuzC1oP6TPY1dkas8IT2ybIok9FYAT7sEeDXc81cBj9xpR+x4/7Hz86Q
AUBTQu0nGH8LyY+7qpdjoSJhMMuUEYAHho+V75gp1Af6oVVQUda6KU+gKa7BCJgu1ERLfl/TGGrj
f6K4K+fbDgqgEnuH8R2Oqx06zZaR71KYMgx25QPyw5IjkNHRk2rxQI3b1S5WeaUs9BHa7Et3kHvj
xs84iZcZeqG0KxzqoIfl+y9G8+53Ly09ORsH79RuVwnZbhJNHoTgTnOt7dd7M19gB7VlHZGWRQWc
yxZWY14f8YDp9K4VFa4QcGEYZN6+S+Uk5n5Kflt0TJaCw2ZfUwur4bvO/mMknAsnNzKaFcWDDiWJ
m0dTPc+0+AcCLpBgDyGZFy+crolmOhjPKJ44d9fGFxlJWSdeWKmrzZ/s32zjtC/GVk/5CeOrr/Mc
814KnME6FGcljxaezE3BktwO73DMj8dI2iaz02Mrk2GefASLyKkUMqOckIpEZJKGkxNj5ssrCmL2
RgeMSnfj5tj5LZLvAkad9EkBGD9/dsGUKdSXbrBel5UmTBZ6zF9VJceJFBo0dSp3A5B4OZ8BK28R
dYsWfMmO89yyUBRE1mMFpRhW6R3C2mZ4jZnsEi+okS1VMmPhJ8+264VZyPZdk/CPsKJV5o344x7I
LsB3wa4wbYUEMGF4k2dAqB1L8tm94B+qtP6B0gNudZGKbmRBHm0JDZFx86m0L9L9lWeWjt8U940a
DXdQAQkUfPZYxe/aPXdtNxOZgzf5DRMZhDVvrvwQX+QqjkKahHDDgUUZ6ch3Jo1Tvs42TBThoodF
Fmbn4X/WMykFh/+4R8uWOa1x1zXo7ncN1KRnLHfIDsEywoBUqvXWQPRJcU1sT5bOPWkJwHEiGs4S
LqDJcYgXMEc0iDcVz/ZhY4PO8XtT77c7IiMt5TXso+grsub8zIkemndCfGzNFghgvbAHmU9SDq9r
pumibmRAyF/hOIB+RTIchgx5fbZLE5mfZrxyJjMzwW6ArOYCprP8R1J5B+c8Svcw42IuhEKCIEKh
bqG+lQUPP9nSkcCYtytJZHU59QhiQPoQGcxu+utrK+7TD3hvBr5F5FxvMiyqJ3Nq22E/tCq6ydx1
0nnLtdHXQm8IZ3Eia+8tx4CiB7gq8447CM3dL1GO4Ej63J5z/MIf0K0i+rbruuvJjIViw8s0WIcx
R88ur5plQVKA8OsYVh3S/xnEwvDR8uioaDDSWBbywCm23y/bHge5MFpRPqnXGQ03S1kcHM9xydGZ
lED/QnXiVuc13hjQT0KkUwJQb+b0gZhdGpSykMHeKZ5IuVl/iD7P1m96xP5tZIdBv0fhI1ki3dBm
+qGwfqOfMRiKVrBJAGYJnl6kblG9g1JqIXXBhcv1uowdfOtNobTSBfzjT2k3HxpkJZXgaE1JjP6h
4Gu9R54DAVs6QpDDYoKy2Ot9w7eA+3EghRAeA7LZCGwqhwBWlJCjFZdnoPv/s+prwrj8OUbLDaUx
fD6Ka6huBpTgyoyBySqxsmQUvJmjuwGZ4tXMxBvYpF9oL4f1wGt59dQF31IJBu9HfyW6caHPCdmt
iQ4U7fVWoHiPVkmctJojMM7EkdQV2XN4kvJ1nGNzcQPRXR37BDEYoCL2a7nM7cfOLNV4/1sAP6VX
JnGkLbBo9IHOiMhyOqrfbjwuBKtVhKP3C9N3AmRMXPO9ZW/ZvQDSLfOgZXPAClskQRsAXAtj+zJK
cEr48RJx/JIqRjokDszfkYsfoLh32Y39D76/vwMydqlkKEEUk7CQMOra0aOfreICRhmAt2qnFZXf
7xCRsy8tHlYKLRrfgSD4tEtatcvRdcL4s9QYtSP+TaeRGoQFuZq55P16rwwC9p/o5h+/Up7kYXak
yd1EPpZwIXqwFfI/kgiWc0F6THmlEWbVkJNN5TdkQ7s2R9pa0Z6inYCfxetwRo8Xve+pc44YtANU
NHVMXokXgqmJYFo6pVn1UJUqI+0uV5tHDNdr/GFgWUqLyvEYZ7hwyLxmKhVfdTXBXwJSh1kubrLA
lWB0E7atD4cO3P9M/EoyfGjgH24hkUkPd6dpEzHy7o5hAlUvLTidKCJPChSD2efE1IBuT3LXvTv1
/WIf31XU96Qabv6JjF5mzFNOHm+CBnUqM8tJTTHK7V8FtCGE1QQ6XPg3FcSC+3teosEnzww8vN18
5Ao+f3Ixohh/71tjO5k1c1dsiVwTqfeoO7FiKpExVvKhiyXEaYvRBt4PnAvDLZ4bIzmcKZYlL2fx
nKcQ7hH5FD03G1e8PO2sZOmmPhuUg/D36qZBPlBJ9YwQc/u02dGrjwScx2L1y/65x7xnkX28LJ1f
sSs0zKYk7ZsQnIjp1Cepf+mA7253nh7PCtn/9qS4D1ffR3aXL17aXn+AbP8rmNk+vOQ1UaK6bLTm
zN3Z+Kveukf86TMtZK04zrn45phsxOpCYC1jKJp9n3Kbe14v6oScrrP6Meb4OsH1gxF4zs2Zxtb1
3IlvItGNYgEdKKZUdA7ATuLHq5zLgiDDtImkhjbnT5spvfcS2sQ2BB3qDAXmdQztA/saDrJ7q4to
uLLemHSYPuHGDqAlNKxygZFjI4g8iLe5RRBZxtM9U4Tv76/P/JgbwJd/JzjJoR5OSSX2RTm/r8py
29tiQZnxn6ZkRsiLQVc4/Bho8VdNcNaLdxi33HbrAOuWB6aJtWkEgnr08kDMWH/RIT42sl4XITMu
R0Sd4lPrTW7g1vEkZLJRUFjaVsxU0J+KEmnkoo2k8hiUZB+ThvyDYMuabq/Bcgeaku7mi/jS5SyD
d7pCoUOImFH+yNz67TfJtQfxYJTLaCH1XCt2QN7pnEVAHvZ73PBh39ylnyh4IAMe3vDAcF6jFyOc
nOHPIKmxLESaEqgvia0nBtNkw6DEjJimE4RtenNcQoX30sJXh/WodGC9a/JLaGCR0WYhGYPaIIJd
5f5P8oHNOVmsZ9sFbRl1eUBiEFZcVA3vvlWPpGhZQ9W0JbmHcTTZUb3nL+fZsuM0bOnJiKwU5KeQ
hOhi3lE+4dVYRGSNDMVHcGWrDszoyAkmMRRvKvuoPNQnnuR4N1HAiLmZB+tiCFKhaqDd2IUwNga6
Sv1MXQyg+KXbT3m+Gx+ZGF/mcWUfEWSK/WjlZadmwCOHb/vVBxtm38E2MU9xOQeq4KuXfr7cIveN
0jOMFg5nI3tWGC/mX4RrWXkny/fW97+xgeGAOaK63oUFLPXt7ndMyDjKjrh3kiFiWTQCGDNmv/C+
s7BWOUVufbveJnRs6PWw6hYaKJELZKZWBYPzUEBwOJJnJhB/0nZuwxgot237NqcsCAqATHEXUcmh
3ePQYNdu7kE7Okw9fzCF6y0ojHjF2JRw1HvQxkMDZN4QgkqJ3aOabMHRblgxlwjxKELq80kdWwC3
nOBvjYhtvWJx8Ap3HDHr1clUcL8FTGqa8ELh4ufs2CiwF4K3b1Q9pcBNfIT6SvA5m07mziRbmX95
Ksh9IagzDcRuqFdDqpJC7CWu/m6JXwRk11W+3DeavSNKHuOSHGBN3nxOzZllr0hWOjOlnKcOYZKK
oMzghckn9w69fpoqYuhVNOQcVTvaJQTJ9qIpJG+ZetjHEf0YxU8dPrn8PVdA3K3hfD5F9KEbX7Nv
oIXjsIQTbyr1yeZP5beA2i3b14Cm8ubJGX6gkM6ijlvGLXVDCx4KEsPJHLjHW8Zd/YwLxCk1d7yK
NtpLbr0QDvQ3na7gJd1SovejoPCU+32AacZaxV1AaJ5UX1u1vxEEtdILxLryQjEgdEAmr/tLpAu0
H+M4pzcyJZex244bt2GFD9yXjROERVvwJ0roSxTu1Vjb9j7cK0iT+xsB86YkrXw4CEc5qJc27PL/
wytvvXIZ8Gkjby33lYOXTn7aU4huLa/wSd2NEtu2gaGZ/AfLUGpwu6weYRirlPTnnquq2I8z5JI/
c6dwy3HvLX4AuBpb81TZO2qPkNSVh8S5S/4ig96KXF3/ZQnhGQ9xjXmkQczH1VS2mqomCFC6Jjck
/EDuQFFMcNAW459q4OZW9/N2djex0tdrLdvCsuiwE5HKqHGJnWemzD2AvRU3bIWBUld5cDV5OQE8
vK8+C3xd+I/oeYqOF3x0kjZP7cg2ILF6fSdwR8Rsx1x/ZSwei8ssqAbG+8N3X8+C4+DQYNhZ1HJv
T+xeAesSTWiVOqCNsztMz/4uTzwPkUouG018+hhSUDj65xc6Rf42aNXhQ7xZGgx5MbGxHIje8u3h
ZOOSHJwWUj7h2bDtJUOg3srFF4GuFdxtBzC7QRGFrcYV1CBdOTz54ogv8VBfEqHEQPcUTrt4zMZu
AexCUWjE5lY/Dm1zWK3OEW1TKTCHg15EZO9GIxqLqDzpa4O7WtVE/cpv6uOuQ6HrRF4W1fal/01O
3m7MXQJTsZ5VQ49s2cHciPQ6bh8VrqFxK2avmVQBWFTd4BtUw6Quc9IkieMz4kNsq9EmEhYlCUnl
8u/BEI8K16eg3D11X2HSVVhAO9KjVdQRWHsuinfVy7oX/HUI3+Nz+53VK+MQZyyPfklI+bgIkgPk
gNOCN5fYdWXCkF/t3FJrybitw2BlmOG3bwdRfWyyXHNrdC3m2mOwBCLMpcvXmF227fLZQ1tqPTEU
Am7f+t7Z4ZJvQVSWvSz2iKLih+OgVEYg1HIGtr2iFSP0USW/Adxeoq897fU95+lnjxaZttK0NTXr
SZyYBHDSr59MGy9AKKSjaTESM9ctosjIi4IMZiYyfl7iWCn1g/27mw7sithV3iVcddVvG6NMUM9I
bDN18Ql03mwL7fYwFrNLD/hVKfT1pIJTsDtBCSRlOol0XlvqR1Za9Ep240gQzQCcxkE531WAT+G0
ndZwNz262I3B9wzLOrY64kEMog95vH9nG3fcY8zIhTHAsACBoRLl0EhxMF+rEvyxEtcEedKOkszW
a5/Z2IoMhj17yWA+qYecs+bDd8X4oHJj090ig6BDXusT7TEhMsYW5ctCT+etO2dPGuz7+zhuGCxB
L7LKqWr0KKY/WKAkjRmsLmu+W64kgdDJ4I79EagujKixPDk8NJr8SzKnlC0cmx2eQyKs0pDGxDTO
eoFmNiJqHD1rexJg/KtH4syiMEsjmj1QC3qHUlsFGaGdJoSSNnjjH0K2QdTcZ7FeNsDDoy8aeVvE
N6kHICm57IBQipXD3q8QmkfqnUQfySDwPood33UP7zYOQZzVhkT6cNLajhtFaW7DpxAN1tFUqaeG
wIsM6OqK4pkuOlmG+QVcwKhQQK0AkShq39M53hpQaFK5DAde8sxTAoflw9SzDNxej7MdgC48s88+
/ymMKSzUK2sq9VmpCCfj6ILxbm3vC6XKdxjrd7/IfE+VY4EjvIhLYwF+/rtOzDuiJl/GpihxusyA
Eq+/rW7g79QArZAFBcVFRSSSxRtlgOKHBaqbeYxapyeRldF8dzxqQaQV2f/fAGRuYShveD1aGxQU
9Zej+/M8o7ivtqozZhbshZbFJQCwrC3+cZrA9QDTFrmFOPa3LSdr9dNg/b41Lflu1+Unhux1kWv2
6Yqz7JuXRtKUkcI9+KJqwGnnKtGdbnCUKRgPZ3tKP0KwQl5bv+qcYsj95EQttmFc2v6nWiCpajRg
anKYSdN+f840dv2D8ZCR0g+xGn2TuCBEB36f3AkxsXuLbksfFynx46OYWfjHELUb43zY7PbaOTmj
UIlLMU9+gQ9t9mXChDtMtzOcQKkULuPTaWpq8/CzmqB80KxT5Hk2S4b30fzQCzIAXOzyd9cIUktE
JhiElhE5P37834AHFjUaXpN/0OFY0JVxVTBAf1AsqqXmVsfReCi1ZCF++zaF4gplwL1tRyTmrw5+
owGZSGqxggnhfqJcLWj1pbclRXUDkTTqsmgQjZboo8WJEnk63kK8mnmRKxodbLuocaQo0fJzhShm
VcQyi5Z7t3UWcsi8EhzVd0a90Mjzq76KhZF6U8yZLn3u/+8G5sd7oOamLFpYgHyj4JKWOSIQFawY
S4KjHLVdKBg7HXiREyC/v1yUcymN1hc4k/CRbRMqisLz+mPdPm9GyHsLLZC/4XhSzewzybX8Fssi
RWVekDE23et9K2aZNWgpfRI5/kl2APlNbf2lmtVtD/1Zc9RqtZJVP4JDrn3pYVrjQN8UxjNA48Wv
ODpMfFBJpn2jvVh4OoiuZKi8xEdHYcuCi/kCK0v0TDN1agQyCbfjzrbvADcsleYer++S+c6niPlr
EqqDRugFOQ8827GgR3kJhVHVzIMswOGwyr4xCfwMPRFb/uLAylMSUF3hRzcTfo8WH5uSQIFJJCfq
DfGTPMTmsi6n7P/anQtTBKrLIy+Vynv4sXKOK00D1lquo6AzvsUt7RsJYJvwW6yjJ960ViveC+kA
q4axyX24H3d0iikJbVTeBSwFeRNYVfy3aRjIn1j8upf1UwQuwoBSRbKPBsovMl1JIwXQNP1RValv
WlGem1mZ1ZRsyGQpztxssp4ruVSlO65XNQoIz4rxZc3iaTyKSf6+142GUfXVNOVwdcYcSCuh+WpR
2TtkzHhrMBBHuotLcok4AMx0ymmQDhVhMosGjMlz9vqMNau4fYi7UhR+g9Yt40kGW6u8YONKotF1
W5BEAppjqVUM4gvPjN+ow9B2Ykc3cQSo9qJsslBq63cAz7SdnMq4Ht5DzcT5C67+Sh7YsGaGIsNb
gR4vEW1yLINeJMMkg5bWy8ddBXbmjMZo3cfNUJAcUzOLVFhnYebVbxPRnzH+VB/cidwx3n0k0sGT
lUIYocpMTVUZ7rDr1RstGwhGAmcAjaTxN/CDad5Ld+UlUT2GVzAqNxQyKiz8FH8pORDvI29hTr8p
hGRKXiJ0LXtLCnTF7zrMH1VCk3HRAvnEyz3O/GkH9yXnII1zv9ETh+pH1BeLWT94GGeY/xoMt322
hqGPCcyHwnxyOGWQb6boAYgohomjUcW/h6AVpSoxK2abQK3aQpZfMhu8TNJv0kUEXI1OFsFts2d3
XalOuQVe0I7T5tKfXxy7qx4L9i3bFwJFFig4KXR+THLitnD2VQxpJW+cTR8uP9R4Ozb82iIYg5zJ
VOk+6t8htUy72j/jit5t16ho/vgSQ2xDwscFFXRnEWxw4Xi9bffZAAw/AEdtU5spvQunCjNfc8c/
aChJtrq9dm3q0vgzRCCaNTbB3fLjYuYSYYnCQc2eQEeBWOOW30n5tCDUh+YtN9Pn20XXnuQUQyJP
MglhsINUg+33m6Q6Wn4i5QRFnUO1m1HKNsTKh0teiNmF5qE7qp3lphh7PwYl8J8kpqH0p3C3pw5J
sBGMYvMGie82KGDOQeVa2lFqD3v0KVi59b2HU/caWt49pIzLY2XvQXEb1LJicgFq76BbgQdXek9P
DWyAy05YrHqnbyU9nmHKWj0N4GWqfpg9DS0KSrN25C0rdjsVhede9KgqI/EJH4hPsqvT/vQwwn1f
BVgCF/CvxrNG1Awm6CiWwEVXS+myq20bLi5uht0rTBpylP5GcbqlDqmlQbV3gK+ByL6bE4DTqqTk
P0Xt/1V1KPNBDSJ17hkDAZ33Tft0g2p0Ot+9LJ+nkph3nsBcWMwK4ZqnOXsCr2FWQOVOL2Ic1i79
BbH98eJgAzJg8cwZWJZDKgb3G0lj+Fac5auwq4zgviRgxDe3S8VQnJKy2CD10SUFLNf/4csxjkt/
KrVer4IpQWIglai8nmaqd9khaf9bDqrlrZLyiHr8UWkmgCgEZH/fJtYUfp6ti3Xnh3shvK6rdS2M
cUcgkYcbB7Ox6fZK1ViyvEwvvsPIoOh44arxVejMiv3YXeYPww7OsxnSHvOk+hUy37l1v3xbydsw
RD/21sybHBIImjxIr8UM3k2uB+Wn31UgpVDL8LXNkf262ICUrQQrEqGABxWC/2dEy+Jr2/oGqoNx
me/15BrS4Yd9qdgWJUAyfpdprkRfHcY0+e6OAPu0BP19NT2ZMrKLCLkQPttmNcX0PEWdF9oHy3Hq
R6Z0p07fbyq0X/G/oaelh6PGMjrl2xlrO3qi3+cjNrEUywFNwhmTNevWsm8oAhhBIH257R4CMZM5
eF2bZ/VqEgrQ/6jxKf+MuKVRl0NOZW/V2SOCGIryRFTcIJlSMp2lpmW32ovec4wqwSfhpiLf9FQg
vxBfvrNWwZO9R0Kzz35n18OjuEyE1Nz5U9d61gzKimKMWgE/nIrX+IhcIYbTxzMlE7BhSg7axl/d
xWxj6qE1JZ1G5tG82sHnyt7Y88XOyne9zZxjAeJt180R6xxmIJc4jPmPp678oA4mg9zzEDGwLlyQ
hkeNhDbhd2bsGFqrphU1SITs98AhWGaL9tviMXkv45nL25deKxwtCoN/n2k/Vy+cvp/fQ5+bYEkI
XAISphdIIs3X+7pn538RjoqnMi5av0tKnZ1CsqMSypI5GtTgvCDqbZ4Su5hxAC+jZ2MXAu8Bfl/h
ddGCPP/LVE/rlE6vIRCvLY5QfalOdfLxjiYRqSlOrgqbL/89sDTt9/XwUcCVqrJFRAWXE/z0ADPr
wJ0aRsh1Bb1jlH8fD048ZpjJO6UWD2NVbxxFx8LqQTMPeux/hAKj+DoqJJ3nmTokqbsRnVxeiazw
luAEKqrSVuH3KWd9vgusn02qOI8L1sSgcwUq76MRk/9Iwk22CYMxhwH2rAE+onsoruiJgClbd8K9
H78RmR/JxpB1MuH5LeY779VEW7jUoOSaT2o4VSgWz86PptdWvtGgYxKbZhDd4tAz0EaZeOXEZ/+7
SLcghCX/ASQ3IgOu4F/BgPbX7GCpzgRqtZoPf1E2LJGFObQcD2PiJjdOpM0Bsgst4C39xgie+Ufe
G7kxtsSNfllYg0GOoY+em58qkw/3m7YiN/khCMlafVxe/Qgh6SesUc6x7ZV4QPclGGheHy0EjiZO
QhKy27yVRCRLFcL1p1prOEEeMQoxx4K2sqzGpqtJDEhZhP6B+nSryqSwFeq/ThAcDySnRleN6krM
ZT9pMVSEPkDOR4lIWkH5IjEcRxQgvDehWEAapEepxA9H1J61jd2DONZ1EYDBpNDXYwPWTjTig2rh
i6hFKoQJ+egr5E9WiNP9hzVdPxI1WoSyOJ8m5lJywA7i78MDbrOUYCWo55wemiMfAXbiJvl/y0tT
t5ha71d5uNszRUHdyhxzmO5SAYb5f6Hy64Kvj0lyvAqr43YsGJXNQifsTnliBj21K9RZ1g5zkN1T
VKgrwVWeVfMWa1jFd9zSPFHzKtY4bBF03+IXTbHKYvM2hUR/jZqFkZltVvhOTfK4Dz13davU+Toi
3aKQA7WLETkzvPlSlnteVG5oQbho9ek72kdoDbw84pyieBns9bcj7oaWaA/RoTj9BM5AiCJ8/WI3
9zOQ9mpSo6yBz/slsyijEn1p6lU/qY6mohLY/xh/7ZvSyBsZoPA57zrLLDDrYGZ7qScdkaZH2ycD
TlnHuZyLTDsD3Iffur3mRY7dBPhfS0ITKkFhqsvGNhEDP/Gf5rJ1sOK1EElmJC1mwd/+B19fK/u6
qYiPsqcyjyATVca9uOOY0wLqs0WxcJQ6OYf2AUT3XlIpN9+SauNjlGPqCXpdHcF0LzxNViNz9Nsl
ZrFIDefwY+kkiMjs97CTzElPZhkQDSYo9kJWviGyaQCpJI0GnOQBFqgWAas984GpOt6+Oo+FLGpd
DkQjpD927RmCjZYbzndcXPmwFIUa9TOCgWC6uADlS3LdKqjDOJNGvsGic2DykeIYGeZ0Avmp8paD
IZMBXds6rb2INIo/nto8QrOSCb1kNbkixoH1J65ABPO5+jJyeXZzlQaSyzaWJlPDBpxIO8o3RyzR
Kyn5vrJTOfjUXa9VBa8F2VtWFEOd5d2rDzbd+VBTk/TBHo4HjuJEhNItnwV2+gG8AH9tjsGAN9AZ
O6gqhOcjli1nZkSF4pM0AydApwgfRPkEl6Gh7vO/RDgaEGd8zvDhpV47c39yCdtKMH6P97OHg8rU
RECRgrx43mseuWXbjPYyvbHtbGYN2K1NQWS1WmWWLNwO8ixvjb9PKyRHBtZ0/s15+QwjJOg5dPuG
JDds2jF3kDa8n41DgdB1tr1bNiqznoataTaN0kop9PJlMHYy7nIvh/ja1jAtNJb7fg/hbCiFPEN+
l2WRrf/UY7RWYnaAwQVyMzzGKyQKmjkFcH96SqeVJiJFAimjBNuhBzlI0zTmZMRE3Bh7V9/t9k9P
53kmwRxrMQ85FZtly+mvnDhiKAq0pIaqfSBt37iAfIvsPvgF8+5nRcfAgow/hi7gk8g/+od+xqa/
Sob2dtfFZk11QPJaYqaF7tCxpAliHkTup/wf/37XwUdHwWfoKmAfgeHS2f3NHH+tFoNKYps3CqJG
HfleRn+725Kq6SVxdOaE07472hsKkbf4/PveDzQqsa9ko8FT6xNRq7mJWV/Tk5V1vCXQRJyWGNbi
jx2kDOQMRIC4dRCdWX1faygbGkFPsEWXLUw8mmr1SgbXuwoAYUj8y/ppNl0TUYjKCf0wZpSZf/sD
q11CLRACR56Rrv1rvOJspdDHPz1llYTmN1oQkRYuUoHybss7ufQw0BUQxfy8JfXbh4/OUEdWxDSQ
8Y+T/XBiEBA8hNTLqEB2aZynUVLFruchyHwkzJF2xc5at1AYWTiL1VlLCbXOeh0yBXCGb6OwSyFA
oeh6n1Wp/MAnuV831wdldPpCjWYTf8znlIHnH547gU8n5GZALbkSVVGOkv5gGQwuozmRZy0frMBO
kz9CGVR0elj/hGHnV6g/V0DZ+nKaNW2Ldcr4C9eLMkU3ennwIVMaK4M2b1yV35UgPyHI2p9nCLIW
XwAXKe3T2f0UXACu/F73TPq4MeLAhtoP7ZdLiKv71dn8HwErc/NYFavIgB0loHmtXe1UgUk9mkS4
oC+zjgRLIxr2q6dALyag2+3cbj2vum0ANgMC1PdFYKLDJX23YPIc8z96fGqzMaFTbuSu3zaBwvLp
lh0VT/2GaWcy48DQhLAReL4bfPZBHwPmTQ9t4l8dmGo6K6+zqWFRtkcNPaDSUZln5xvhlz4u9mZb
Peeml/50TX3QbJws5/FiN5cNNMgAewuHCVq+3K7KRVxkxwRCZMfkyL9sIPlDyi+OfH+VP82LUWf1
KmjBxCNYpAQklUqJ+HlIkWN5FdyJ6qfCSIn1cFuagwGA8hoUW5GQNJUa6XWE2Yk90XEktLHWLJTZ
jXpUBqvIxO6bCNV5uLoWkzSqfcFZSOo9roQo9IHXuSbkglwfz2BHOeJkmRuXBSvRkOeXEtBh4FAh
2QmzUweunT+sNl3sJ9L4eQac8OwC/zQL/VTGDcr998bWt3pD3hF9T2rouOId1ShJ2HqRElkPZTHQ
kC01r3ykWAq11o0hBmT+GO0u/9RP8db4L9B6V4DKu0WEJUFqS7oeVYbRleFuNwS9hhu2b8OYYVZp
wZshlI9P2ywNchcygYuw4VZLvWxrNGqUBCcs/t9EjwE6VQZDN/NkcyIo2cxHgoeKxwRfRXgBUY8h
DhOvvjnvr7cOv/VRY4h8ncFzV7frSugR5n1FRMp7j+wiFMu2xqPox90VWobsjaEQ1QRFk2MfBfIl
qOK2Veoi3C/0tV1a8H1oMARUB7whqA420nPt0k4WKWCV8ICsJv+kpHtgI29wmZV0EZ82CeIXke9f
37JZJKU25QBHV/HtJDnO/OXxsacPOV2he9l8RBvOhFFYXQKRhxJW6rR2AGDFjHsSpJZLfLEdKP50
ps3GfzFvSBC3oXMORw7JI69/vjPTRvTPp6BcfPwLjPW8WqOHNJnOPykMrioEWqbmLFw8m9cLb0jY
cUT811LWhf5qcHxbPMnvXK5TyYhzJ3VYFOxh8YH8/M1epUBVkzhP//aMnj4daFhejHfT6CTPQE9r
0SgvSdNuZRfeBtxll0L6dLDhdRykw2pysDkg1xwHDgpsi89+vsJlpofvOCyga9PH7NT3qJ3ZG2La
U0sXxqKq973FgDhvayb0/vvnNUvOOO9xrr9oIvLGS4Q6vDX45L5nGW9pY07nKlqiqlnEkBnURG/7
kOHarH6c6RhRrxQN/05YrlI9g+G0wLJFLu3XtiW3uLPVfhGM2h5FQ+umwsTWLoqeAeCIH5reFjkS
lEUYz4p8MWldlq0rrjsEM06Kk9hl+n3WUICvv/9//KT0+vHGeXdxpALuXuAITZK5jMfPBGEbhQ/K
bzq7rymEZQFfmI40vmTTJpJ2+tDSbLmIrSGMKjl5DRLbfSIRo0Je/Sp1G+ONzfIO3hbpT+N/Nu9A
9bAZP5fPcSre0m3TlZDoB2PxbQgyGj18j9gQiksjDA1ymiY0uGRUW8xT8Oj+Uh2GXuBKe55eDkur
SIvAUdlCvVPJ9nIVUkJUo6u8QRpw+SmFkjUwVyYdgeSU0+1UHf6H0gexe71vl3r50LnSUrGoQ0tK
MIiwr0HUuRBudBnm40n3XI15+bqfmj1DVfU5rjXxYAP6VuJk9sTkFXpQdiW2AptBdW5l5jn9kHrd
c/b2KyAQJl9DXFw6U7iUUdvWTwO6fh9IG5npSQ1MyXgW+ljarxHULfrkaO7x7D/ClbO3rh3urFnx
YbZFn7F0wdf4KCmTEMXjX5YzDn0y0JEo3LgUmw/kbdIM+Ctv5BG6XWuWJMnWtUA5OQFcT4JSbJZ2
SVWQg27uiE3Khg/XY8flBHN+IHPQDkMdMMZBhpKLAgsYsRHkp5YOWE64sIpEU9/Vb+8h5PRSOYu2
TM0NDxjN3HyY5m7mPgn91VnCkpLmEwKGRkp7PaJeU1A5eVamNR2Yl0zKQtnURVAopFhVcBVdzlTD
Qnjr3P/opuPOZH3XSBJSkmFLKYaVRqBz+xTE4OXzPmE30k52DIm1+vPjnMU+nLHyZC/exxD5s/3C
qzx0QIBBH+PvB19xKHrnkBLNF0ixVZ75fvvhcNr4V7iQKsFY76X4qoj2m+KNj6/2RKOMsNng7M4i
r5SRPRSude1+cSOL+hOEUZ/5mCAOPlmbJuiERRWTkzLtOg2Gti5gBHAmLK2uK1AKMok/LdhTsCgi
1sS8Vl7l715YBeIyoysZu89YOxQ9/dcx+0zqYK5J0Xd7TPr0ShtLf2f5DELlx0ONQjho0cIu2XhT
jp7+faAEDIDNmf6gdA/EN8CLQDeGdmPJPam8yXkk30a96rsQVR41Op6c54YWPxWF3AxCKgiZ0Rth
Y2Pir6iuaketoJMNBLKOelzmCdX0p77rmW8DWbcIQwBJunKqivKi/JiqqSYh87COLOBnXmQv5geX
UGhpX6vI9GpdbGaNqLrnxV+U+F+ML1QZX5QbdzChcmg+QFPMfo5tk70O7lzwdqtfly2wRgshzDrO
K9zoqv8CbDIaxWRUKcGW5YRkKAXLrGTy0oNQYI2VwzRx7rdZ/UHXOAaXZfWKRrAZ2NOFVNEcXQ3g
yPl2kiDAPbF0JPonSiyKj5yBLhWJgd01go4ek/prYA1XSok7nzjB8EOaaR30jbtS8LShGtuF+4PG
BrccJKP53OlHXO+/3DyqjYRM393PeCc0Eva7e79zs9iy9OuoGqyExpfAGmVOPHX3P8sdH2deAD8M
x/uIZpv3CsvwvANfahM1bmuaH4xwnTkHv7ZzO2f5M4eCFZBS5cDHw6pMgHQa1Okh0qdaRIyRfyoM
dP8NBk5Nv9W/R8pvCWodeXOyYbIw/6OFhqPWJ70B+ldtw9NA3XB1f/T7+zM+f5SBCY1LbBuQpjZo
dkNnPCujBHkXzfLPd9q1c4fvi5cLEKTx9ed37XHyh1BSS3fyor3xSt10TNdsp85X/CoM7A06V77Z
ZdumVhtaOd4C68z/2seZV79p7+TAMsgGi3OsugDanJZ8kCOZvdVQ+Anf7plwQvagWmdxg8yuqfDM
btgXYIoYZ0UPcz4FrpQXMkjdi0iP0FpdlI+MRLzdw/UTEAf3KjBOr6ArctTGIFywm6e1DYZLbjU8
NLLAqODQna2/DCWcsXQwtDlS05NRDvvLVV9MD6sBhEYO1coFq4hfFvvUGFo+37KXpABHkCRDGY6o
4s8EWVw0eiOdxC/1Gw6uf+oNA6b17o1BMu55lJsnBVN4aCtnatw/GL0R5HGvnbuhwFfo6tgboLCl
5kyTNosTa4i9/98OuiWBnLRgTQ0FkD0a+oz0IoQcpfIs21YviHSczN0rw3V3pcZZ7qeO2Q2R7EGl
e0H0BTr3L7cHJT9YM9G4OQBs6rGa4NpvscvK0jdpCedxtgi4w7p2cypqqb0P35M8yhMZdIfG1hMg
9l+oI3qyB6ElBhvhU41EhlbV8G7onJICC0W5K8NSf93Kh6SB5Hama8sG2qpBuQrpjOVhtJqVSEVd
wrQJHz8BaDD1sT6ug/l2X9g9ywNUw6jDgUqmx4nxrTrEBmqMVxrYLKw2ZsEtm4Z3576L+W/d94Zz
J39ul+NzMpdDXifhZIn/Rz1Q3h3vfHUpK8grVjAihgzngTC25bGPay/Pcb1wu96OlRaAPU48w/0R
jOsNMvJ2HxqyECPMas1CpXludlgBzDx7C1sOBq+G3FMZpTmiXmn6It+rRZDFeA2uslsYm6J3/dzN
I8kY7Up0JZd2QPxtRY0hmACtW9tz8N+cBEWg0s9WPL6wvpGV5w45fEr8Ufmm/KfeB4lS0I7wBsto
bKIpxXgywBkHuh7oeFtq2ZMORjrqL67rxiRPqx0mxBqm58qXky6wqglNEuQ0iUpnamCE85nPMpxz
MJbQ/2cjIpN9WxOKtm6FJwSqN6LP8255MYVdKj+OsztnariCea1pr3PzgQK4nVzZrVD/2+2ah8M6
kemJgEUiZ9+Lj8/y4giKgk4HHgDZcc0nmlwI3Uo3G4O5D76VMMZTHrYcSMUadCVlMqhwJ9NKZKlJ
v4d4EVbTFAuJLPosCqyq9bXUQ5Tx9bqSzVQfSaifZRT5fwcPrk3DVauP9sbqP30yFJK5zf3jRuLY
RcvIfdmlZxYb/nh3m8KKUw6ZVoKEQOyg4AfzDRiNhGq4w4/8wsCNLBzGmRA2AdlH0JOJ4qYDjTmH
tncrAkQS4CmdWVdPVJTXGwnlWwS5w3bXhoYXCPYj73vEdoaZ4rwZSdXt3xxInEhZh2g0C/2AKvpI
YcRWfQ9IxZfrdxVPwfSg4sOSuzdm2xV85nPRYQXWeJDvvwQDMDVHFvzdnulg7q5xotx+YRxUbUFa
Y6afz/cBPQhssmQGuVZdpJp2/4Uhqidg+FPQBhq3zSbagMXozqXJ1/Sk4yQyG2YAbI7M5sLTGAHk
weKo+MStFhav7hOR1w3qeVfYyig2ryix1jECMhMUEPyy4N0Dwv3xAmf+G+xsIjMFNizRgV5NcTyX
bS2sjbmf7l6elNHTwJNw2boJJ2+tYtKSzxjXikGyJOQqEiT2DVa83Hd2U6hPkIj3aCGEpyt3dLJB
Fkd8/aYb+6X+Ci5cMbMKcbkQQdR7Myc3MZn/gu0rtM8FTP5yjtAlXyQnDuVXCiL/66zaX0s9Ggcy
TIe+WTsVwOLfso7zy3MkHVnXvnL5WxQwN496YwsnjCQ1Pnf8eYg8vKGd/0dLP3B4Vrks4ueQXUyP
jDieI01Zws0FOEf3WwEt6rz65IYDQ5ISSmCh9xyJ8F0tfhTgzCJOmf6yhrjyhEwxWcCT5iwS1gWc
xG0FwcAvcUH52F241xx1/Z2InX0rvXcyGFKnVEEu5fZnxkJDJTXKwz/v1ySlEamV3wRm6n4N3PUi
UQ3Wo6LhI6gQJF88+YCoF69roA1RoimtCR+C9D/JvFRQsT43ROBxuGtaDVWnAVubKByEFzAmijBD
g5cPSnfImKBgyZjwE6SE/YpvrHNjY5ezUSWACinqUwqiaYuyruNw3Ebwirce7Gcc5Hj1dvB7ZyWn
Gu8yVTyz1K4BTyjVchWbcxCbimRNNxiH14Ey0lo4DmDOFQqhbOjNyfRIYCYnd5iZsPVaTEBaLIbg
FImkNmo6qidLRlM40C8agkA7walfF/bIlN/FzDOiXKi18Mqd9dE+AL0yIo0+dlCVFkMtbefo6KC3
XFuWmMZA7Ao0nI3tARMR+6j7k59pOzyoNn5qaJ8Abnmn8yAG4Pvre8acwsOBP3msrNaJWepYxADO
jkMUoibmQspc6Q95I+nLKfbMtq97qmnxOt8bWGH3GaF1jR2XTPM1/HX5oqm4UV+MnKI32qD7zA1L
vCoQrwQH6fl1z75pWcQhAPwLDodfjlEnFCaPGSU6ojZCpcflXc9KKknU6lwDYJ5B2AHPErpe8/Lx
yt9tqHo7HjRb7Mdq5FmmVaBI6nYvD9fk7Qf2fsMuxZRw59UK7HVqxYvHvb5gFomHD/iGCuvxlia1
90zUK517OOT7mC9zsVEjHxZ+aN3jYgSXnfOWhVLJZdQIOooipnICL89ge9CI//r5j6ZfWzXkAusc
D7x/lLjgPE7cAXQ8Ph5SMz9ESzVcaaxVhGFa9xoSaMKNcqa8up4TDNmKVI6tolnURLzv/QNUDV6Z
SbeLpX8o9HLLHw3S7sS1xVz8NXRO+ghKr54OH0kQuprjTKszsNhF2aChP50j+GcFnprmEERQPvuY
1u/sx3lN22Bm0ldLIb3FzW4M/zilyPxsKm8yzR5VlirvjUmZpT8dlENFNWB+FoxHBaBAP9gB/8X2
3xvodxlF/nvGKPkGMTv8d950WIiMH508pOSLkIBDtIOwrR3EZSnSh4US/GuybAiCs2Hpdf7wTqjR
TnfiyU/A2mgwDEbpPwVEvJ2zHoN7uvnWklRZhE1/6fbezTz8nceKpz8tlf3mcDgiIgZ7dey0Ze5C
RWhDgpaqSUQDV1hZTvwRcKOHtGnqD6eBvI6fqnqv7n5tilpMrnytEC7JeYnpeyzEpevRH7WLQDUT
YlJ7Gy1qB5cAslrkezC2Kbao9cYN/kUD/tl+kY0RJUagiaFDEbFElGiiNzWp3iE1PgyeFOnmVs0r
LOXAhxT03SFf/UcAvkIleNlQMk4BLNeVz+P1RM3LHOL1o2IckqvhDcCAsMudtllx5LRip4ziBFME
tnWiP83EtWVAAXvHMIvMObs7cpw/pEUKcXV1Vk8o5sMX8OWArnFp1YUs/KJ6ZKJPd4MnpzLlpyxS
PI+Z9anNVtbof9EFx5NyLJOFyFj6VoJVZare+VxRX8pZHAHDO263IPTeXB+DlcynLNc5YFpCzwGM
hSxTXetJbLOV+x4DiczKVKy484VfJOol1e7tL6CKYxpJ+/xylzyzUPpCxmLIgDApgA8HACWGi/bD
hXRlvCwsoxhDCYPuOa9MFGuy3DyMYE/5/fVT4vlelTipQHVIj8BxtQDYdyz2NM9Fm4W6AZ2nNuQp
02s7vDS6abEuk2/egRVdLVmete1pgzTnwlEueGbERi9fnZ5KlzeOFFJppfNuoy4ZRLn+6cN+cUvj
x3IznvARO7vePMyQJInDhYjTKPLBerc4579+yJeMwqv8PnzlyOwN+Im2xDgF4BmrMlMZGWaM4Yyd
Oa+k28J4Dv8C5JgDusZI+hZU81BTdX3njZ8k9OSjU8oUp4DA3T62Dx0lLdXGSlbazlZAWW07nk6c
MBt6Wpz8M6awoLoHUFjfa7lScKB2xoYK2OZH3TLLa6PkndQYvCCIi1TXzq/Fxs3ulTtwkWfMwA3b
c2Fd+UKapMS35YVprVmDZ6YxEHkuBz69CuEhGnPihyeII71QzSNMivwbS1bALyTbJ0STjc9wH4y1
+LloDcXXiQk8BI56TGg3JIcZoBTN8j19etNoK6A34PuPmrOhWMee9YdkmiSXq2BNwpA6YZ0LQSFu
o3b9dOreFBM3s21gTojIVZPHw9nW8qdLETOd7jcCvd9VkwawHC5OcXuRKsKu0hh6VCgu8kG3kiEb
XVFOBctECqQZa7QelGe10Gba2WFhNapOGApzzngr6jAZTb4KAgdHnZlM6Eq0q50iZIyeNC0GwHfD
HQRiQGev6bxQSjh8ksz1oaC12qAM+9KssqHEUsnnEPKYtKOfB5yHer6CYEf1as9sSREQcib/bP2F
CVJyRnCOvcSJJt8Zdu8FSzz8WfZprO8FGzFMOIIuVKgXjI8R1FNO8e1So7AUVdq4BttdNcdFv0n2
NCu/nSOR8pOrpu0eA9LfkUmPdQOQGl/N+epwPE1YNy20is5L096j+12Nn9TkZqqPbn8wNktsBDHC
dkKv/5UXVRs2WpCsfHadCEu7/XFy5n6/Mwis8g8OHLuxT97hB6gDK+AIrnsCluhPX38RhErCFuD6
LWQU6Y/OWtOFrVM3sUH9LC9tyQlrSUdiFN9/WUf8nDqJ+R6CCC1Yd3X1H4LrE+crln/iXyYZRCvj
5AH42g1J1zJCeARuA0a0TmLI0gVVEdRgzNkmn4XaHXvXe7vzPUneaa4T58OSZ0Be+3OQ5NXAU9+D
CGTKOoNWbB26L2+0ASB4xlNN5K1/ZtPVVm2WkxTGIKSFYsIM6BVEPDcQBnpp28GcwJiH49YXmKOV
AqwglbNThLlrtCtl+/m2BCsafT/z5wmoNeL8l+d3XfRLEv8euBCVKkARRSffaUe776MGiz45nvrX
KGEAH8wuePoaCozP8LRTkB6UrpEi+kDZOURZzo8N4ZC+zLpFVc+7llRUoHKgEwnHRjUMdEsbkc9n
8/B5oYSsrRj3Ur5lm+hkrMyoIKtdRV3magINSxKlehJrASdcQ/Rd1ImDjopUkXO7MnRerdvb8m1r
6mY8Q18YTBDaSvPYIOye1h1/RGxzQJo4SXyMx7f7U8q3sbf3/W9czCdy81xZJsg0JGCyyJIsDI2P
Pm6uGtDkOkvJE1vGccDOtO/ndx4FQpKXl+rNtg8ZEZ+zHi/HkGQ3+5H66OkI6CbJO/zIqd+zXnX9
JnlgQKyyhnoDyu1fc3G/s3BfL5/cZtellgquhyIJDeDebxE88HXXyBBscBkTBuTAXE7fVbGYmVjQ
Jn7+oUtGc39eYTw3zfQxYU29YlK6X0k9gKjUvVOBnml9arYaT5XY+VczvGoLAH0Ohabb29XdGy5n
y5znM/SyynNrsf80K+z4LkyCeVJYuEdeNx1PoIBa8F7F8ulphx8mwRAHYBi3bprfl3cCLELXUtbw
lesln5lK8TvNIRKjAVjpFZTlWNqIT4ViiIMrKeptns+buGCfeCaemnGmwFCc0kNrtcgdVL5W+42v
MG/U1B0Xc9WkFsEQk+d/nY640huHvMoPpKEj7Gyn5tmdBF52WpHNvWWaWtqMg6k+GZyTm0qkz/0N
X3b319KUAr0I/1EMKYuFA5yzigeTkpazyjn2tWy0lHsDNJby51ke29QYXWbmpCYe5IYn3KxRhjQ9
JNSg1lM3SiInI+cdbPt+GT3eJDLKSI9cojsqLAGIItKWOiMfVbnT7eYkqdiyV8fAmR7t9V9+9Gue
PqD2gb+7KTqJe6kDCuusL6vm9EpcjESMnS9Yb4qiG/u6Op35zvegW4GSTMLNQxXmfWFGzCcEYM1v
GBL+HMVCdejACgM+/Hm4iJ3575NmDWOLPQWsaFwpA9hhvihnsWJse9/hjxb8TreTCPgctOJHieuM
qWlLQ1qso8eo2Ts9f3tuv88NuI0WJKKADdHd6Wb/l17LIqdIDRqDq9jDMxi3pEp7GMeFZM7mQkZE
/eekLDjfcC8d9pmlSf+9lCv1MnVh45CbC/3S4rvW1tLQHM1kWJnHYZ5zRITwiILCNpdn/cpJCSOZ
yk58xRAr4feQYQ8NZfUD+wCgxxpgkPD3Rb/H+kqSKPZBFR2Csw0Zi0kgz34rqctk9dp3fE6d0Tx+
+R+jLwAg/3ZrVLImvwK1yzouvlUfi6EJUoW/qx/UCzWUviOSMuQgyEjqPIFWYMOOm6V0sBSzX7dj
o5wq8F8dKukSf6Bz9Do+7mS7e7ZBoVJ4zpwCmBLfgcPbtqude+BMuwv6EIcS0nsVIqXfPvjJcFQW
oej8Tuncj+DLxrwiGOEsklE9bdyz6UQydozwgNoXvPOr4inqMBC3Gz/LDpAfY0p2TApyYxorGP1d
DQxeVxocTu5RD72Gdb9o7FCBdpfrEtaCpTHf33FgAJlpUA/IoLMNeVpg717QZ5i/3ukoZ2skQ/jk
WG22CtTL/rz6KuVNvxv1/AudmpB3HVDN8RAXNRsQxRowUFHl2j5Hs06OmFcdthXJuyfatvw3akwB
mP4lsf5gGZ7guJPCGBVB7/z7fn5TsioD8U9M2aUHWO+z9c8MczxEv+JvXoAqI8EoG4jPag+5iSDR
jmRl4jiru5bfgQ5hyxrOlR9bt3UxxrzBYaiX1N4KgDT1LNpGNibsz+liAWQztCZmFDm+kILSum2W
ugcsO0O9ilwG9efTGGrJ0CK/Yo1BeN6mYP18D9AUdOhrZFYtxswEwKl3JFl5xhYo/E8KsvxKeGU5
SJH0zSIeYll3eUMaKHu5uokh3Bpx6BkkFYlHk0BmZednhTofLmX7Exq1IcjMYkGXQjUwyCeGMglB
z5sKGgMFGrNcI1mLrIHZ38d5mKRSsrI8GT1rIJaqENUBEspF3psQSpJNLtU+JGa9Litnr8W1YZJ2
mLmdTNTpEGIqZCDmTT7S7aV9HrVmmnJ0NXTAgvlpt6QfWeiGLcGmSbjC5Ikw5hS4lMsLIjdJUra1
piol5NbYYjSpoinPiA9ResZdS9lSiCJtSwy4LJHCk3XdZC47brKcnzerYLxB4ssmUqMvlMTa2/zW
HoYan6fUSfIC1jM74MrJaVcblq4c6ZAUnKFKMTLdgDlL8nF23UfwWXZbqi9+dYB//2+EaHGZli/H
OBipU4GtLenxxbb5kkIYVxC/WzbmGJywQuCgUfGh6olGkxbFjQ15QzZ8Y8A22SfiQzx4+/U9LUo0
iUGONTgF7k4FxK8bxBOwKI/df41OBVFvTfAWinEKbtVaNf29DIf9U187742FwkC672HMDsvq7V7h
DtrqTMhnRTfHTbhP3yN1UvTcJmiMIHVMZq6kgWrNaA4q48zsnE/lMXJqCrumGObKMqwrDVtQKWps
etU07VFCtrVm29klH1TECE4lIqYJgwKgMreHEMGs84IkMrNNMtcPQkQRf2wJYcpsrnRvXOzXyrLF
xsP0nAnoppHIb6bcO7lD9CBwyg1gA5AOpKs79ZYJiemjmT3+Ecoho43xarVFDfTc6occj9FAz/CC
kfM+Tqylelqf15pdEyW5W2l1di6YYfz2xZhc0BA5O07tSa8bHv6khSnjxD4XYTzEr8XBaQ3/I+Q7
eWarBZO5AIljRtZFF6KWSb6UXqCmm3Z5QqUSzv9SFLHtQEUx6PHPbJU375c0DDP6q5jNtcqD1chm
w4K5pBwXFclkakeHUHeJhzUpb2Rf3NIKKvoEECl/a2KNstzBKOTZwG+C1H7FTNO4x1Lu4Y+qeudn
D3OTNtQQ/iD4V4Qqvzv59lfNWktRQFUCCMpz1uhz2unSDWJwhbh3BwcjqApUQk2JCG8EOtDiuZJM
VuQOm9wm2jxQZLaS+FVMuaiX5HJizB94RfRug6ri6Gqg50GmLUfd+2xHTUYfEWG5/k2evzQxc3R7
ZFwb+RYEwnjMQ7fePmj1UnJS2opKyvnHk87hyyjmsIqGFCoYlCw3o3KkHMf0ALy7U2fWiJ3JFXOj
UZhtIDlP6nveC+zWMOoOAxTYNfUqI8qS/ls9FKmot310dfasXTkU58vatY1jj0rCj39LANBMxSQE
tO4pqIYITNg0hVxEfnu7rA8O6ZYE2gKu+QZ5M+XEqGcG2p/phEnmYki8cIkKrRBZzFi/b5AsP4hv
/zWw6W6FvCwKMkfGruO1gyrzODas0eoEJshdyqVv1y/p9vzg0WayNatQCvNhy6PreGY+NnE0Ulg8
Vkxql+oQB0k6EPjnKaTcK82gCbQvqLSyPkOWsuWW6PCGeAM9g0sgK3u0KJcKIuMgVp5LMdDlmBQm
j8OQa0D8gOgxbRH/XcDOOj6iCeEuhQsDyqBgEcSu9TfEt3Aof5zFGCpnKyV1py29H1zdXv+v1eAE
vxpcJVNoV4a9yfFuxpy4mygqWdeTb6AnNgqQ5Z5i9qXmGgu1WdAcutnYMohPryBVMsKnPgag8BHh
sfnDUVOGQE1aGMehSAlAIQuyM+w70eXG+2RKJXKnrlHyS7txa8Z8mhr17Ds0iEgqH9hnhGBTNoG/
7Q5FnxguSAdatE58jz2p0y7nTqOb0qN8QXCV5WPJjciqL+Lpc6jGt1XhkI9kCO+jCQBhlDWOIrM6
JpBKg+vHu42/hznb1vHnbaQXD0brigvMRwG1NxfOVnk9EbYmaZVWlVn8u/WmRk7dPgxvnAUJI13P
Lc8pbF7lb2oUBhZ4BrX9YtUNh1ANWCxHl6V/UDhVM4rOwmHqYnjYakLqHx4pPN1vIx4Zj0Wa83Dh
tq8qixtdDiRQJWWU/HAXW1UUHTdHHshpe8q03E+SYBUOC1UnM+1+oeRuYQ5dukj0cMNtXTVXrxM/
BNz9kjM0iaOpgm32JHi6S3t3QfXYP+wPldOgEBeI7IUQQwsXLUciaOxfnGFq2qoflboEi1VLe3My
EHuBYqVURORkYjKl+rAjW2Ekm5fORYGP7SlVgLO0nmg7nK1Tc38qGW1RkcgzYiVqkH3uuKgnOuFM
+rErLY6m3Vx44GkVzpqDzIdveRdpl9IIuG9Ki55z99XRrqOIRytgZLT1TPrXhvZYwysVPtTRHinG
7FbkCdXMxiCwwezbDaMoXjd1+0qLakKlq8gsNjFtpruGThaV7XzElaxwATGV6TPJADidRnZEWlwG
cX5FvyDcRJofgy8qn53i3W/4mmyelTTX3yQalvXDpGMNCsDxgT2rc2b407TeqfkZYCxUtrXuYhmw
cNXKz/wa08huWb1qkoi9klvY3YlKOTCZH0o0Idyg3RbHHiOiqBsuNf99D2V5F06dA967QCHFs2nN
Eb+6zTK+d5sWvv01CAwoT/ZWPbGMTxOsFM7CfMXC3R+P9iO9sLd9XdEsIgB3s/vPTQ76Hqq5KVpP
E8gsPoRd6jNcl+PSviqOPtxD/+8FBF2yxfCoiWKOLpd6RC3M3kcB5zzz4etDS8O4Z4yq7jBlp4vc
RBHVXUmOMncHYTDPzSzO/dXJtO5ZICmrF+uYhOKRovcCuVAsjY64xe0r0z6Z5Xjg8lDkFm34Bwmg
yxishazgJAihJaTumsr7RwAROw89P/8h4AwJbkuiNHr5umf+h+pbATaccI22wPDbWrwO1JfatnFB
3F39AMKpAsriTpMaTl4f1M+MGMsV5u47IBDQ2cBQxunnOCFBi3hfgnxufG2Y7aZwhZDAxD+f3m1O
CoXUce0DjKKdu8HCuPgFG4I1AfGUQkc8xbvE2Zc1GsE93az99zG43/eN/iO4R91tVA7aNmiG3Hcg
HdSeQFDXpk3Luna6m3RiuISl4zF+A9WWG84ZWRzLkku+MA6ncbaBMJ8w+4bbJgLAsqSVLwKFXVPI
S6rYnX1Hzb1f9ArQMXNMar4fNTY0lbmSlKLd0F5YmMVfXpBPyLyd8+OTW7taIO868fgA3OuV8Uuj
pSXGHgXCh9SmR7IG/phYrbseP/d3cwLBeH6lNTQCcq71R/dYi+oaDPvHhI6cJw6OH3k6t7eaKiDb
vDLqy6iS9KqFXMjSs/99eqvboHxnuAEO8kkB75yaqjgC/msw+6+8uctMoyaty8n5q+h5EyHXbJfN
yH+jt5V7Y8T9m6j4H8ctDiz0D4LJL+Ub4kPlzxLN7LwehKD2uta4hOml55GxTfjpwL0OwMyM2UbT
s9GWh3ijWoPPr1C8+Z7OV8ybWri47+iAIYtyOXTTkfanhbBmB5l6ZVn4qxFwEKtp/p4QKFVjH2dw
M1TeZMI1FG7iRAG5ReRBYFH4ORR9qCUJ7RuPqf5wukAvN2kfNYrlcpmILpwGNZvnr6sQIxQRG06q
YZCc/XfDsWl4wKK4bN4m85nePOTllgfuvIw6jqyhhA7km9y4a06Q9R4b5HaXwHy0f0gioJICFCzG
2aQMkKfAmRHpcnok4MpXXcMLF4DymsqRGwBX34ee92YifT6lPI35+prIGLm7CRD2JqAn9B9FWqq3
Ez/4JVMOh7KA440TBU0gNeUOTG3klAYwXNZQsNmVyWU5DTcjEaETEd1MRudbOMMVwjHWmWznXG50
s1FsYeLthJbTgK9kkNsXY8VQTyNb9KG6Xa2rMmsdd4iuDQZuRHUF2GqUKe1GTWNInWWOhqJYDKFE
VTrRv4RJ0dd5rjl9woMJhQeOU0G7BHlXnou6BtN+Pta6axJJTMVsSqXscyyWF2CmeUMDSu4j0jOP
U562qnGa0YD5q+QvPJpgm988SgGjucUiHFDBUOdS+B4WXLmLeCax1V8oKiilcfd6s0bHQp0htr6U
eEWN6hlq6YGvPtfjxC22O4ukCqFlJbwGTVr1kV4GfZVhKrN0VLSenyNFuB05unWe67GCzgRPRFPg
pAw7wWGlr8UKziXqdI1GBZhV8MFSfLdQ1MuD4Xkbci0Ln75zTpxjTUOPAV+ZM0FcErSKEUGRSo6G
oMsMZK6zgRsWVYrlNeExiUsPtVKBMrsqNE/NI9vXinndRlIsyqOAtuO3TelaG9uy2xbGY0zN2U+2
tAUw2sLhp5+IId5xQonZiWXLohNm+Yt9dlQ/SN2uPWl0nV6xMiLXFT47ZmUSLahCpDCeeRh4DoV3
ZWIFzcAQQOLWY1tK4G6bf7orlzRtkFMQSDpvuwgQdBiXco3PHVbJ9448F0zBkEj6S40hfek7NFyC
xXF2Jqr9fpW+WXF3kFokcFAsEaDC2UBTNkjYc2rKXbBo6bEVdN7FCrFvq3wSNRaUC3HuKehsovMU
GYim0bN0K2DVRSq+usDfglHVH9Zoat/RTOl55tmtyyey2dCbYNRB1U0d9BxFofxD9ewu/eZbZhKh
jIwNGZG+lm2Jc3rQZ/lUJaEditZN4ea4+QqgfO2UeWcCX0WJoHg9FeSzaSq87zejad4KLNOSH5J5
1zyhODeLejgp55b8kPbGna8s/ooQgGtGwAiErNyY+jy1rxbkx4fjkK/TlTX57XI5zgZhOzNlDOv+
hIjO5u9RKV5TPNS2BJDqZOtZhgPnv1xhdL4dgMiMQPJtKamF46O/ILZKU1AS1ckWInCNOhNpFlUv
MJTu5LEZIY7QFo8QgLNeOaHa8RdqJw7GLdrVIvsZZkZfQOcNAtN8Sf/lXlLHQxsN/8kfz2ud7aav
cE3uYVB/TMINqzIuZP4H8+5/gKcVRmAKjK9ECuplkrrmkNjzISaqvD5gJCE3ZlEu0h4mM4XnGiBu
eH7KsmR3dhJP0dLFYTJ/ULbYUftwJnJvX24n5Y/y54x4vXS1AoVUe0JMLvD8k6cr25Vfqa0J+osx
WMjQPXt+aCfyMZblMZbTsvlwjOKJrwFimqA8WaPiD4TTiTQJoqck3vPocls/JnTVq7meOrTZNPBN
VrpyRlbJ6gm6LWlO9M8jzhNT7OXf8uyQjOUOGic2yfTOfsKuGCsTPj2p+9OqR+yLA66mTSHYFMNy
6nBu0yxkJl4bnLfCC4bH4v8LUU3bdIxLWQR9pDug+n+oXJr08V2JCbwdafcA4ccbSuI3GP97yT+t
3pSXwPCmhmbJ17e+ow3h8Z8oizueqQ51y45dBWNU8S+CItR8NZHcVjtDGxwY80n1Hac+Iky43y7N
IOKCQR/etq6FiXyTpyHprTcGfXSg8x+LOMHcIGFgk6o4gpMQgTFSYda2bU+FTxSiPo4DlSekm53h
lGKZSVAUSbX1u/r41W40u/3WsakSlwTvNGHIIGp4lgKwO5v7vD2idBxsFbCcbTfLWvcGsogLVdxn
+bwujsj69jcSgf+27WlyeR9RPBArcAsffxl+1yAF2GifQGFhFok+qUYOiqHOacVxj/3ivrFGZHEN
YupNE7PoNq4zsSY1HqK5mFMg0JnGdjVTjE7iSrQyQoScRGNTqVvR4r0RS+A4Nx2/RT6fLupeRHAG
Uo1YQLxWAcqm7SMtKK7iP+QRf1Jt4JrjlGkieAyPjjhdr5DypPPxIU/s7ih9fH0hdLd7HwC88xXG
LF3kczZVsPTZ1+qtf0eypndOnYCU1jvYpGH0zQfDCQsxAP7NK8BYc11shwKvcks+ufN/5jXrWMqx
4xgyQN0D+JzaI9ceBYV9O+J7+66PJU4j07HgkXCiq/khoEi5+eYali2LwInarUpQwFmuFr4mn3mt
t2k9wCdHTedVPqoYVjfigGDTdouaX3gDUdVSLYX12L1PYANEwoskVfLVuCqDHWyT7jov7Fho9yot
4nlFRBMJP3FOP0xRTWvN/qSxuuoaf9XFwYkMfu6yjVlL88IXSwGqStaaaW0njpI+tovGu6prqCXQ
XrAg76Pu7K0PTI+DhektgDmLXL2H2g+y2YGFFbqZWgV6Tnb3pOv7yRZqYF5TdYVj2A68+Qp5lGnB
eJ1PrL3Yolx0SVV5IO4KowWxSJGuelba5oVEuZEi23LQlNI2Fmzafb3Jbe/XhxRN81XoHQVFlPI6
Kl9lm5b7CnRmHSGrXnBqrj/YxoNma6wGV0KAceyOScd4vzuPNO3QJKehbNpF4Vp2CNVZi7bqL1cj
85BNlVoEhwPRaYy3djmsqWsPNwVvLO1f3Ci1L0KoXcn8aCHlBIHPFEckT0ut93wmcYK4x7rTHOpW
MrU+ANHdIKM2is5F8FlQeGv8GFARdB9v/sjyZlXVFB9LZdkWOE0cWZw4R4udIhaEl5vevPEZdoBX
mneLanEIQOzVk9sKvSH/2bfEkwf2EqQGU4HE4RcOstoPIsCxRLcXZLk3J/Zx4q0I+ZZaZ13dzKRc
qfnuAqxjEMK6LU4USDjbMUfI/gmFJpSFeRPa5VKKBaCE6iAG7hNMNnP146NzSESPbkW47SOr9/Wr
+Z3mrmOayUqpKbQ63XMqsCPPmqQjGpg3eEN5rFekMyma72SJ6U6IBYM1uBb8/sTg/52IJYo/6shh
61nlxGBkEdziiN4Mwzquu+ONZPlaeHUZMrrINCaKWev+FyJ92CasMPYnXJYkaqHo0iMc4L5XMkRs
oUpqR38PmgGlSow4jsoj+18QlTHI3CPvIfxTxd6H7Phr3Eon3/zcgl9Pj8Jnn8MDkAj1TKfzflF6
PCxI9icxI+GDqzCZD8qKdBu4Hel6/MI+Nj2FZP/RhP+YehNYfm1mLgVQsdGMPWvmCis77HL1F5br
yihx6wV3EFIRgQgaPvbOfunI7aoo5LZgB9enX4L2eM4zT/LThZGyesyqn2uTaNa2Hh83C1Q7ec+/
5VF6zPODVHjgTKWCksxI2KZHsMmUwtoJSKt+sVlTJgCiLiP1pRkMEHpNWOVaytS48pRTcEAm28Ne
pgImyh4wuBTP89vFjL9dmNLnncQRl9qOJTZLvhKY7Up0SxAwyrWjAZ/svHYICsvRxdvR2m4viMxR
oYvXCw8jaINaLDZtdyA4TKhO38h8XOBAzqRpoW+RAcCs4dlkP0gse7jJFcoUzZq3SW8+8gHgFZht
Ir5aNsTrMgV99VpFrDcxVJp42sUXnP04Gm5trJiqTM4UsCTUIAQNMp81WfDs7Ufb/A68ounadUvW
7Yq30IYOFhryRvzi2BQEPl8GnLfm+S3mh4/K3V0ju4UCgtb4QSJORY6hCJoh5SXvB3V2027Na/BT
i2OiBBI5/xplRRxWSx7ZqbFf7lF36m/PM6fk6vPf5dCIwjrOCqcvXlELMBYYQdqHI0rofg0jfLfV
Lm1skcKRP4VYufphdJY4WLvCv+xSas5wBrH3AmH2ofVem8Jj0o3kNbL7FjwF4qsB/Qi0XhZ3qrsu
5CeZB3FWK7E3jgbwLxLmvVlCuokYJ/v65LfdDoOSlLbZ2SUjeLvuYr0bQ019pGCMxeAh3kp6aAAm
J8qm7ndkrKIO4DuCiHCq7TGjFCVPcbG8fDJ44J7DtFYR0eg6u/iS+VEU9R7vbvzrHMYOWq0d4Gyk
9H4ppZjplo0w+m3Sm3A7Oat8KJ/xAXxaEnK6rp86Ys9RdVaGXhxrDA7PiURHB/4tG4Gw3UYpCR/E
dW6EBWGl01Bl/nMRuXSlRBk6FA0bBg3SeU9xGVgRdbvgeJdZv1p+YtzYsQ77aQf5eoI/60l9ehTW
RqFyveMtYIYuxAAb3XYn4Wj2Hy3hZsXKdHFm/9KEE/Ki8BNTis6lu6bP2kQ9iUsNKJ7lptihQpmz
+6JktHTnOYPJZ4U/ImqzdcMke+NpFEnUrMqulFjSQtpzIDRpkg1KgRpR1xzJABn6DDSjQYWVmsZs
7eT6tg9uvB8TXgNJKckZ3AKaIwciu6tFBVDSzUbptsgSD7xF0hh07trqebgPnF3C5ltz1Zcn7csW
fmZ0k7g5tJsDX9ReQZaSS33eHjspOr3P4X7DZe8bKPMOPIvUIIkKVAGADAqgUpIe42MdHGyE4KTv
1Ju33SpZhAaAccxdC5/4hv/sKPx3erIwCQsx8MjSZ8CVNcD7fZoTyf2yiL5lyAd+WA9Ypi+zRTjk
XSjYxvxLLaADcmoBaeClpl1a1L/sRSuywxYVANgYOpWT9Z6vmV4hImz9yQNn5/IQEeSTIczzX+rZ
TIa3GdlyD40xFbzhGVZbms83gDc5j5e5DThJqacZawNmrofT7Yzd44zOw6giNJ8d417JEl6uSxDd
/korCQpVuD4wovR9ZNKscRPzW5Blxkc7fG8A5Cqpkb2tRBq/QiNypdv2tAQz2qln9kwuE5tZLUvZ
1ofikrzwDcx8QMN9XdoSVZ+wJ3U/xcnBgV7Wwh0p7oVfbg7moyiroVmIrH1pzturvjPHAN47WzCm
pS66aje0SZ2n8g1lVT3ZOUsoVmzi4LAMHfwtb9Ihfbv6Nr6KJ9NX5oyHlWJsSzeZ4Co6xRQW4apZ
eFO3yA3kdPOSh568ytCJa4j8PQX1p7RUlygpJU8EcZinyOLFIlp1lZUVBMPcALc3kYbaK+4++nCG
GQXRAZBXGgM1N5nYumENTMcAW165ZWTEsEUPbJI7ZrRj1HsfIwL6XQsIMyZn2pmM0J5obHt/+VPM
G5Ygb+ZTnCFb27WzeZWxl2gYkF4b1c54JvcrGTzXAEHH1taRFaduwGEwFjCpsYgfVmBTt9UoZuvL
cx6s1nWRDZGAJcLkeURc9kTsG8oZy9pCfgeTrPwIz4dA8XOgJHVptX7/8lxkd2s7FSQK6R3f95rV
442cR+M4rU2DpHstXQSQCgjKQZav2au+DIq7cMggE+UJR0h6qsqp4qWdmUegQiYHI1LWkv7jPDJp
Pv5jjDpxsqGtZEkb0BYX/S2ihrXKh77bLmplWfiLgwku0O7Zc2fQ07aNIo9No367CAJx2b7U7+iY
mIexg3DkrTQT1bF4HnHbeN/NFvObAuk0Fwi8coiGRd+T29m5W99ebDkJn15jm5DghGtjAgFnn9si
azZux88sgNKccw5vzOf1DdhLJzOeOsjcZ/VHggXaSCCECW8ZVuKxZKgb7Ghll2sAjd1r5sTRfx8U
HvHTI4gOYF8mVAyvc4CeazMB1qk68eqoppSWH9YsFXj6wwTgGYQF6vs4TYAIci46/gVkHIIOkLd/
RKm1iB3+FZJW4n0MIJRpFqLo15sDjRFI17mb93oiKlvFGkLeEaCVz8F3YWKBAnfEGgtCFLAeMQzT
eW1YgD+Ws6XImteZab0j9F/wf6FVeN5x/HzZZXQqVGMxjbv4UC8hexqeL3MO/SuUpzUUc5PtnqCB
RYy/3autFqNwwKCy/7o1UwE57E5LN356j8QscYzUPoUSXkFoo243IJqQWREdjpFGiX8Gi/v8ldmB
jx0eWh5VrcauDJilgWscnYAB8KaS6/mCW0OWkQCBY75ZB8Ri6/9nHk87CNhyV3sgNnhOBbbcpSp4
yam1PFrbQcwU9bi+FcN/VrJhbB5RAOiixlEwgYgQ9Y1Z8TDKdkdeXansh1iOJd8SHKyPCTmCPpSI
1yLRvRSXgUbGToGQtN8/zWYvhdoP16hL4vCzpohLkkN6VzOgl4XwZ6FhUucuEtaeR6ukCNRO9lot
Lxi+1jHiO6mrN6Tw+2yWV1Ic7aBzRvGgZwP0qkjjg4P59C/Q48OeuMDjxw4Q/g3+3bKi7AQJbh3K
lgr4+fb2SC8iT9+R+GdLGXNzNEqrysEzhJrJ9TWTOV4gsXhuMPyxg2kNRfX+tqHZgLOTiyLM7HYg
eHARsnNZLnZcL+F2mPqLoMRu1FjXlr0INdimBl1u8dQTcKXec/6gcIkGGjhauUENxpC+Sxr2WGBh
SkFm8SIAriH+B3kQG/ivRuaQseiaMNZ27v8LxUr3rQ8owbT2A3Oq4SJ6OVSc8apNYbYRTQSKSE3w
b8UQrA3Sc8eZcFgeaIBRMK3jHgY2lSxZBc8V6iXSrIulVGU37rP/tye/I0esdzNMkCkb3rqMFiO2
c7Jz0ksOAGR6s16vds9p9j90tag34xZ28b7sZuJKrQcVAb6mdYwYf7hJOdwBp5LdD4gk5abG8rfS
OPkSi9UCOoSR0nkIutwvGBgdS7AqQhqzEZjTJZEFQHK8Vydpt5XjqHZm8jL3G2A1gHndJMlvlsOq
ADJaza4eaaFetAqlvl8gVl+O/Yn8PaQ6esIfO7ojtyslWRXvuArMr0YjVXHVh4gh0QriDQqyr3gD
V1iLFW6+ucOV+Z2Dut563VqG4A+9ZS9tRiWHO8yg9wSB4nirjJotGIkU3velrBqUEp2RbhcwlERY
BaeA6GnSvzjlW9aoP3A6solNnc36FnF3MEZHB6aKE2OUDbfYw611qRLKW6oWwRn9PNvG6LXJc0LX
qM26yUOB0xkHNYHrX/cxh48NOOWWamiEsr7/IjY2fRlfHv7zyjRQdBNKiB5sR9MQ3G0XTU6+2RDA
6AQA2j8XqjBvHXNK/pQ+8OhPdc37DaHTaE3+ilj3gtFWnbupUeZQkWaTMFTfQqa3+/U/2G2NoMF5
Cc1E9tS6kgne4Wd6xJXepXu+AsG3KXC17DrQzyJMzoJQOS2xE3xADhmk8PwcJVFtK38ZKSCbZk+6
N3smOPCaHGT5L92mVEB7GPqvJ+8odSNdmLN3226Cf4TT8ZAy9EkmdFcYYxa5u1VNttDKdzII1+Ff
jEQbLQSGEjZCiN/jE2n493ntV8mtPllZGvmrqDEqfj7JZdZVAhDWwonxqnBsfxr0KBcmSZNzj/vB
GuCjCaUU/krKUqpxPLer00TABor4IDnE66D/P9WIe1Cv3mE9Fw8TCHtvKAWcZRU/VAaJEUu3idbw
BHW0138nb7xhY6mPBspRlfqcCih9j/Z2GZ0mIrO1Nl2NMOLDiXYsbfO4o1M+wVWILAAgPREojrgX
dCIAQI2Xb2i/jxVTIan52Mp97weYDG8OH7I/zi7RUediLgItfgl+EA2A0apTb7TInlwj/2x3kgH2
eCYIXZS346dJHKmWAKe8mO9cL9/zHKAiijPWcxRKw+EAOc1F+xUxs+fTTixxPFUA1P4BR9rT/Dul
nBtaQdrbLiwmzj5LwJUGEyHTLOhTusPjrVhdeCvujkzNBqya4YfLRKikSV/Nbxe6AYqYkD5aSrC8
Y7dVh62FC35ti/QIHCtKfPC7n8spzAz5PpanoxkaavheTS+PinxJp0mVoivrOJKRw/YXAvtyKUkw
1JPnJvHPt7ma2ExuaLqPVRbQYdXASUazbMIVOaELa3p1zud0ehWTXhZehcYeMNR5YO4JM49AxE6R
76xUr8UQoakCzZaadtUeeRyVFCQkuQ5dSyGtt8GVpyOGNnCIBwZF58RsQb8d0UW04+IJR3igsNoY
e8USsbZABawDIZqSs833B+vfkNJaG0wy/N+m9IK0xGQ0nrwirb4V6nQpdfIHb9UTA6WUNaZXd1q3
+0GcIAytx69l7w08ZPb85ec9eKqf/xyiBQBbSNEyicsxnXpVyy4iMw7uXbufdncBrWTrqWRwWrVB
iCGkkDHxn8E+JW1dOd3HfaGxiYnCAv0j+mhWU4/fZQEMCVnL81tBD7lf/lmGsDhnkqnl6cPuUUHt
Zehk3HqI/uzNfPW5b50yEyIo4guKMpCaRGW835bdDg4rl/9VO8WqpAb29NwP44A3ItNmhkapgv4R
7cOz5SnCklhXhVN0LxsEcw7/D53FaIc6haLwhRmkT7WHu9zd60MJDWGryw6gVyuw7kTG+lvZq+I3
ckT5XDdA86l4rX4GkfMG9r26iGklpB7+LHf88gADsMkzOvwvFvCmjDvPJE3VUU9U1BH+v3Jkp6e3
NeJ0CL+Bhihi9ucN9Pb5L0uABh/13MWAguUPaBGz9Ro9XlhDW25ncsx4Hy5WxDr89355kMqKDu7F
pPy59/HBYMGGzvOX+wm8aeicWmOVvkmXUQnXm6oDTVRKOfw/VAl/9/33ZcqyS0r8cVQR4fYtr19M
NPdPJ7bk/6q6Bye6TjkstWIDmmv1iEk6sNUkM/P38F8IFQz2UafR+zn6nKG50XeaX1XN5FM8mooC
75pld9Z4yiyZYyZerP7ULGymq8zvZkTJh964Tr4PJY7eOouimp17RGGd8V8GbVCbtHhpL8VnkcYl
grve/s1+u0sQ1Qr25FCp/kN9G1vVysMSZdt0f4zGX9QalBatLGp6QeoKWkXIcLfevtk9lB2U6lna
nbNnfuiwyuYPwQpUCpwV6SXUdiYrGuR2U2OeFVLkDbXW7jM/vUKM2nFCyxwp6uUi01vmeXlrMi2e
CLH2UN23I6xkWC0bnzHYEySFp4i5W+NpaCKjM6aW0XOptrbayAK1HbsqTlLOc1fZ6lhQStqrvsz8
NdSTXUSrmkpcZQuQYM7c7+qGqemrhwzScKEm7Tp9yuq6oYJ1paD6JbZlSVbScBmQ7BFeEba7BDQl
OqrrLHW5FVXt9HwsyYQKeu6onfp4CTGIZDY+gm6RjdlgpMAckydEop2620umDfrCBuz4BXvh/hg0
lnMnn5xqkZREdgAx2nJdPkOsRSmX0Zb+H1iae6RWmUdEMTcyvNsCjgOkF3v0P6zgHDUaeBvsdaRG
mYqSSED/d1Cq1MViT61t1Z9dyXzJ1R7b5sgn1dxrz7bgVpmyAiubHna2JBxk0lc1rqOts4h8Ei8/
zdI4S1/HWqW1+wIEyR2OSOHgTtIz1Q8H57dIb7kPVSUwFSN3PZZ7TZUT2AY0ks2WCRnh0KEbFltL
PbT+hYH2lIbHQ5ufRBENGabWaK5r14dzfMjU9ZRW0GMYU6Az8tkVNc18YAD8A3GaRvhtud2oKNDq
3veeeJMLqCugwu5+wIFox16z9lMnn5pwd01otaFCPR85oM+3zUrKZxX/fiJuBsDD2JfGUeLhXnNw
hhL2KnqNE/snsTM3dgCdkhPZDtE0my1Dl3l5HnjnrgHuJc6danfJ5q/k7LFOSJeS1DIJZ+qCMuzm
dlL2JRAHvrSn9HPUxFMXED7o4qFTcIKXEO9f387am506+gqZkG5wOLH+H3rOPQyNMwLtCnmpgsXb
EvnvK2PBjjvLoLd/bKPxZ4lf4ciHWyHx349pBBE9K7ltBpkg6bSSl7Kjk+mqu383JaZ105udQZfw
K6CqM69cFXl+agqCV4wWWGLXJbaHoy6Fesno7ablIZ+7bGtxM2rjYn1jhBkBKvLp3R8qIlA6IZwb
G/UdycbZC5yg/MT0oAWHbUVV5ptS5rMlgqNOO/VfZ6yY1ynuUp/+lrCP+GlDyG7OxWeBiUBicvif
nE3yviOGJ4ZBpanswjVDl+WYD+Tt+s2m8sR/Z3Q4GMc7WxuX/kIx6VpsbhH4YiLYHNJEQwexpzK7
69baRst4i3UsQUOP+xhRt1dlYtrQBQ9nIdWaLYp0LJyEnmq+kdC6ItQaNYOw/xwNm9AjslYAVoL7
S8z/yf63EXAtcPS4YHI3sIUDArW0qShjwp6acC4C7KerdB9JXZYmuLZjC2Sys59JwQY8cYwVdSK6
qPTR1us6beXQavIjpl+MgzbrpZgTyosdl/ROTtk+qNQMZ3dIkwVgQC9vbYT+0hjJnai2rK6k+KOr
Okjq8lhVLtHWGBiXx3NRj3/5lx8QeQdD1bVogYVpenK0NeID4wdnIGT0QeM3XFDmXZXH+5ZEGxm3
iKUWsJkMKAs3ANAJpKUTAQCqvIShe46fSqvQXGsmk4imwJ+dhxKu2b/F/MHOhMbWoCEgMfM0OXc2
Q0zUSDgWHdVGIhVnzrcKUeJQkxPY1h2TTRGlI102mk3FQQXIGzn/XNYtlYaymhF9USC7hljGlxpb
kBjvz2Fo0wLNZGt+Zuhryrzh1FkxwpMggmLtFgalV++gpR/zfPKvPou2zMpVavfwwt+KZnj+gHlL
/+eIKe7usG2oJkCCsRo8BBSlnDU2FoVNfe8p4qIyaf14Y4jz0V/ShD2ubFHpPTRJtCSycwk2mPDG
xnhc8wM5DIrRGOR7gbJmLCcJVekoAVTxG4Mwn8Qlw+LF93KhbKSpqmuyUx1waJwKxfqwMDtm2RzP
vlgS8zQ/mV+aFgr4sz8KyRxe1Cy3ns9DVqPqjSmZQwRFv5zYi7T9DS/fqJK7ASYpqq5EAbZ8U4V2
IRvM9lRAXzXfcll9oDb8J2cgC+P7T2gNZIAT45weYWXOMhWl0oUzVIfjX85JfT/P+hLD6f3OD6HZ
0zLIP8+DQOTm6u3H78WYzj1drG2OGatMRTyGzBSMrY5P/eCtyitEeXrC/Vt/bmXqZXfl8kty+lNE
nzzTmCA/ZJYjvLWEn+o9dU7JCVfUnohwUjwEwg5yozSMLliYhQJZwXbkzo8g7XcZ6deSR8EGE7iS
OdVJctGn6esXVFqz+3zS9i7Z7KzNLKT9+YxxeegXqEeHszCh+EmzDRB/2mOu3uHAAXUlLJVlFRQ7
y7CraQ+l+ifnqGaqku01sZ/F7P1/IN2s6YhnA0p/B4hjiOmXCtWooG5Qlea4vA7NCG4iOKQg/3Os
5oXq1N5PEU2/ek1/PgdkYG+Bii6tXb6fErUfHjyNpUquQTsddO2tAE5GiOkLPvduu2lJ+ZyQmrP/
DMytcNolaPpqGvJUXoZOPVpfCD/lmfMcGbJG+hD96F8q4JRQtN4kLyY/TuOdRxd1TEgTFcgxrq6i
joZQGh5Fwv/bBWMJkrLUZV8Z9+GFDRUE54lhw4/lPURDfdm+w53oLdDYS+CslV4NPGwm6AEO2sXb
JgjiAiNyj+r3FksGqx4DRbJk815Hobn3gQ4IRSYSsKWxfhJyiT3LY4feJj4S0pzSCB+VJutcL+mn
uxIRauNtcwhlsWJgXZ/5/sco/W7v+ED4YDTe7JQ8mHv2adqPtcQ7Vde9ji1y14DSCc6+okjnJ5bv
9zHa5x5o1L9IIvKgSB0YBWfD/SS+2mAh0FCdgcKmYWJY/mUVugOF0xWPa6+psQwn5tIpCAd2S1ch
C5NfSAHtGsrSzcHweX0NZyThjtVk/NIbvznbq/fCJA1jMIHVB2Do5n0Qh4lOFOUDFJJjHEvHCsCk
bMsfsIE3+3IegGes6pclxRMIfFpA8aUgHc/MuiXobXePKUF4d8xBlS0iS2OdrGku7O9Yh07zL/5Z
MtE1DJns9kI8riWmOqGO7/rWiTnPLdfZZAhOiO5eSdlCv6Cb3Wh3ihnP1DSJKohDXTen6JZY0kjg
73w856RMP/AgETl/aY/27qc5dSLdbhmMh19ZYg43TQoA0PCd6dC6Q3VyAE3k8xmvZDCw40a4PKEC
OTyURKprk7QwWPjfMCAJt/hbxdELyEZpA+hWY/zzqxrf1GQLwIpjq82eaZXX0rcG5EyAnYP0b20C
2kpVyIsbZMocMe9p3nHBJiHicZ9YrepY7bQb4pxKOUsZTDQndPyUA4evXKo2sQlrWi7XdsFj0CdP
uweLbnSPi0IlyX7+wgP3/sYfk8rbEPwD9Ij21JIWkS6Ytdlq5nY0fJQOT4qOBo+rKj+klJ2HC0Ek
hL0lq7ozt5lhBRWT06FjSLqb+/2QEes+RBBgZr8575xJINYCjbBW9Uvk7lLJkRhR/6pT61wcXeSy
1zE7Nq8q1XIbyRpuhxnNjPwVnoAptVMtPjwpjfrGLObF5jTN3rNpu3OPnrcVvEz8vC8lFtx3ItJa
iocjatapN/Q7ViUSLTCXycW6M0e0tmdsMcOtfU9SzuWo8f3xG1HUrbDJtrwUU1jopZp4kMICZupS
eEKZ1kdlCYjDL+lHBY+p5CnsCyg1f6xwl0rKelWBx603xh2U1WvG5UjCwOkdKqNQBN0ExvgJ1wTc
7yyu4GrzpPJ0iQ44XmYiteI7VCbDU4D58NEfUWPLuxQyF6GjsCU9WS4RemaibNE1UD7dT0TSTyd6
FxdmwBONOFsMOwQ4ysDawe09M9H3t+Q8qr2+At73VuY0IgvtgXGYp9zDr7Yeth8qFlRMewXP5PFx
z6yuV5WZN5XtcCqkCG4xctdQTAgoavfr3rHRuJnAKSqkVZX1b2pmJC6z7zvZ0h+h8c0txW2F0Bta
3lJjh4JpCJv5vYFWa/UIeT31z6xwI5lI1FtQBfJf5KTXx0ejM7Tk3hOGqy8Z58LEOhRLk1xsXGMD
AD5XQZy+8C2agBCJOSjuAHBVauuaouivHZa6F3zSHhfB9SvfnoPmJM0gBwOxglUQnCKcD2pMXgx6
vrgC4n1rsm0Z15ZoRpwa4MtwhsAVbe7Rxai3kYvJhqEfywl+zBBKMFqxPtcrMztWfMGsBlRwPJ4U
apwlEYXvLMNMcRyTG7I4xFwRMn9PxrjQ8vFk6EfiBHW4yqxTe2h5CWYnT6R55c2wsgSrdyg5l8oB
+t4oyBGbU0O8ZtSu2fY67tbuYJ8/1A3wmRNwYeXKZZgHce3brQRJZoxtuPZZz8vZScr4dq88rV0F
S55al5v3rXFyFWhb20W1otvQX5Ae0AvX8SzpyJJs6Ye1UUoro0GrGjn9ouNjCfCi7yaYn4txiKgQ
QOG0Fh9Z+cEwvBqEP7xs/9SluGASUIJBggf1QMF39tQic0UCVWUne7y4hQVmyFTzuk6IpSDvsSkx
Ty+4x/SMAwDDePFMi7LHrF2QZvPpqGRGlyLXwPWu2pPSMxXVMjPEFNuhIZNfno7lVf5dcDuupIva
Ospg+Ewqzmq2IT1fXPkfTUyA0noPqQdSL7R8N4UnO1Gx9+zh1sYfRjSiPULRRuZL+KVJe5NJqS3b
+gKar68ovTIJJQjFgTGkH3ZIeh3BthR7+isrPh1u2ZJJjIEQmB1pmWlGsDW9MWtijzhctAUQZgpD
m0bjFsJhX211WT1Ej0/iBg2eixIy1Ay6SB3izx7QIFwoKY2k6fI58r+G1VBXmdEt7QcaVe62kTA0
bpZ7ImmpRNrcEn3JQbb5lXr8uWfa5gqWE9QT79usgohEYpuViNNvJ3X6NLAnTVr4LPCroC6S1wR3
3Uz+fUvJsVMDzgM5FhVI3IliEe6GHmLqHNv2f5KHicd4DJ0bfC40mgAzbICzfeMjPuve1dWbyGgM
e7nJmUDoZiOJYcr1bce6MQ0a32uYQh+seqFd55BkEzp1YG6fN4jsJQGtzn7YTDPBBmJfXJ6bcnBz
svl7V+XdCTZ99j/YLB0ec+gdcT/185ZAXurZ1A8h9eyLvO/hfPyqMVP5DZUlM7WGHwtE/Kh4W9/m
RwX+dnovG5RbSIQQ34VxTGin9UpHlzx6krJhNLtmBSEARhFmq7EwIGl/7pJRcd425wERKPiZFXVt
JUHMZJeH4q2hDsR2v+eFKjt4RhRLKEnU05gRRSGoI9UIPzSvtRSCuimnYAxq6SG7aMjiHldCoSHK
93Z3VNtuHl4G2fUnJ/kwSktPKOiEk0QQ0QQdN+RFjb0hrg63EaBQtL7IL67Vzh+Zdj5LGkZ/5hi+
fS94gPrzQqBjK4kq74KeItsvlXQURlKv/6FDq71n5+lz1LkKKz5JXaM6pNO/BK1E1jymuCXPi9w9
iTZVDOOBStaiHu9HEo9OpyIgm4li6OM0ajwKBmUCHaHXOK3nv0GhAzv5pJ6w4IuGwjVg5YoFaZ3I
ehGWWsawR4ZPer+761s0tsMgPMyHnPGl1rRIkvrwC7TfqK7sPXyEzU+vzR3FTybeQPzl08IfOJWD
gwRxuC3TV+LEclJzStGZfZEqY83yyb20/JCOnPKhQOGJK6jJ2i9fE78mnsbS1kmbYb+AwCd1TyRX
DMwnenRfu7OesCUDcDacHcCO55TOO0A0AYVJ0fwDjWeKEllzaOC/rY6Sup1hNNSu/Bao1Jog2VSz
tepFTMWdn6kfJYagW25Qv7fcU545wl9vmbM/dfMjQZGs1EKbnLOgjma+eLkBlrriRyPT69lC7l4M
Vl0x1H3nbNRJ3LUQnCtCcqo1l7oEfnae/uCnYuN4eRO8viV988OKyr6vNWDSUO7VQ0RhTf/+ToDD
52aQwAKwHiqLyz1vcXMXOYEUEe6oB1HsD2H9vj/LuTns3v+qKHXCmK4GXgfsZetW2B+/lNjprqLT
ih1yiNOOcvdZOfXmHQVcJ2PNpKLbRS93XGzU6gVy4eu3en96n4WF1ZSFsuHk2+zWQdHrD1qyOQn0
JwKMPY4MSTnb94zG6H8sBGrBFlQptVEznu926PLWnosfCCHKUfPNDaphlgNnntiDgowwAjIFACH4
CGfkiqAA3Tf0rD1nJXTYDNj1EvU1xaFbba3GQgtVAH2CuCPyNZG31W99Jd2pCcxWBUuZFQgh2rAt
slnxQyEGoeJBbvuXjudQ4Aen7jF7g6itHYbGLyRmD2qKG4ei+QGVuz8w7I+OaHOZdxFCv240Sa0g
Zk7j9JO+0Tfs/Az5KqC9KLe3drYVKffs8PCAQfW1GB+BBEpxHCxH2F9iycsZCr3JbdgTVsqQBtfG
lw1U9V5tlAEG9KkkUTjeuPFRvwWOszx8JXr8uFZuotQozaFqao1D5U0xK0Am2iGZcr5bguTdRRNj
+DGtwyB/76Z6+jXxwvunZ+84AtFhsofz3muoi/XQJ6UiELJXqXh8iZvB54W0+bXtiC2dghjy5ACj
TWRHqtwCipivaPsPn2C8aBWBb8f1dxMwrqktf3H9nMlT6I6e6hKksNP87kkCSdpSMng6cwFAHNeu
gy8jXrJiQ0txDSjj85Mphd0QYSM2oaijSrqR68UooZhCnjrQooMCE19Kist+jVbQhT8Ly5+yXYhq
FAhLmHEpJdllTtdrl2TxruyG3llS3S25+lvgyzaul8b6RUt2eJqJTvH/5nDRRDf1HoRFXeW23P2m
otl6PF7X777ZharOIdp03ohYs5zQPBmKHoFUmWPq+KkOPK48cZfgMeBU3dLhDMyCg1QXrdDYq0aW
ZUgYFjuhUIP5OdniH9ATrLWt6DIlvL0xtkioXWd/RhFdQcb9ceiyEHrJrnWBX4OTH/G0ytFTGohz
Ks9EwlY13F64MAkK1rDtXYyd/GPCPUtrKoYLoALKVLMJzzwEgF6r5rxbn5mvB1lQ/jkrc0Tjs0/k
TEk6xodw6oHww6U1ZlwrHNThVH6e55jlMTkITHBMryQXI0g/ORGcCoFAwZp6dENKvzjewKF3dnmp
9WC3Zmpk2W86Uctpby9IQSBIVTmDZdfdJs+9NvsXqXqOOkJn+EXHiep8R1GXO5yNLPvgxtb9lIZ4
Oj9+Dh64PETLN1W7iZ2NrfZJ7bpjrKOBdxsJT7ncD3isPjY3W3QxIkqBbd34PBx1JUDe/rwY5s5S
n1QOcy7T7maT0ktEmdh50UzNU4M5i5ppzgDTZVaElJws86D1Wo/taX/zF39sqngr3AcElsLnsDTp
BRlfdo3LnGE8g4idzjWn16jFzfS/osPUmmTslbxiuL6obB1X74veYMYe3vvhDoHyDSc4zFkyohqV
s+pUjIpyxA8CygLbo8kJAt2XeJox8iGk7N9bjet46HJ86guhemtI1qJZ5agZiplh01vFcjeZDm6G
n1/gQ6JysEXTGu/Jp0X7JttLFBvOQY7mjiTQVITJRoAW+Hl2CJEtvVkXnv8xUbzGhxKZV8oDc/bx
twprs0DJM85sTFzIax0tAFNP8SKF4u2XjJ5TGzHGUgdaqNczhKgCDINGp7IFb8isgEkc2hCwsAlZ
If6AlpD72KpjX2Q4kCmkUAyOROSdUnyqbfRRWoYZrbcCanPVaokj5rLLR4oePk/fDr1/RMclrg4U
NOkCc7ieBJrn0cdzybUZBrGZnXGO5FsaXVPshGl+fddO1gAiMilVZa9Trd9EQjB9gnPk4ERTkWMY
wiHhc4jGkJEzFHXDwQ35ynn+RRwCVmQAldKenDD6t6vAxwDgAz3nD2RAbcIK4W2p03vleprIwy7N
3hlTLqLMxI5zPa7f1+6QlBRhXpfu1MJtfxwFOkhy01vfC+vr0vX8BKG+vRJJDXGNRUtIw+7Vi7cL
/OLofrXniK71U9xMxWHB95/TB8liv2lDHRN3BK7+bPk6LewmjcxRNc5pwrLn1z0Hf5erI2QIObMO
/yMaVwdOjqjByQG1xU8hwuxlNfjeil+302cSwtOXCn/tFJYAYWlAjIaYEhsbQW9K0VvwAwDRqQJ1
NoYuZv0r4C9jsn23mIYd41dNarBIMM73paXqanwKMlAMqmQNKu0gYc0lRUr75q9VH/QYPmrzW9Dp
5pM6l9AEja37lqF+o5MmgErD78OywmTNg8blkV4ASqBLrd7eWJXO1lbyZ8STBn4EIzNcJQOSbwAe
Z2J6ZEUVjNZZYSUDY5C3IEDMSUqWzStEkH6dQkg/NfO3EXOCJVTia/fgdp2Tsham5FqEdyZoCfVJ
yoei6jjYwzWrtbWflFSdWeqN4AlhMHPL5gggidqv2BRORZDtpsXGm+wRv+hZ7wxOdHueQtjGAuFp
B0fNH8FE1F3jnL7chyQeHQNwkuGwfdprF0YFXpqWyhTss6GwQzhIiHHFlp6X3+rHZXm5F6PfMNgy
A3gtQQtY4i6zAazDE4j0rsdy5iFYyuFodcyBlRSlvnJNFDCqO9uCpyM7BAnlLZC1NbgOCB/iDfLY
1hCn3FndUBM/drxKPSDvdboVHuPp/exbD1KO1SAqB/UJd4IYP07hwUc42NKH9B+ipxebXi8vYbYY
O3xasApVzlzcl0d3poAyz5iHo2BZ4WknqfRnqGpC7SuMU2eYM+jtAq5mEUd1NHb4bwPr7l3rMU6s
aos14SItZcSFhEouPQaHYk9wUaSDT+KWZRFiqyU8BLPQx3pzQbkcikWKgQ7vm/djREpFMeoqxz22
KhL79K1v80PQsLHy01R9AQzBUznRiW9yqPnvP1oaFh9teENRq170NMjd6L4aVj1eTYUprt9HcxDx
4pxNtkKUX2oQ7wNDs7BE8jz7N6TG/t3olDUu5ZtTh0OztxnMcwV92x8HnJSxmqsd1Z/XxPTc4fUr
CYpE3YgPVS+Ca8hbL6xAm3KUiXvGZa3uUnmT5WgZnaPMy43adPWbu9KVPe20nCfVHqKtFEJJdAgw
2D+yLl5LEVSomZLt6zoDWEYtaKtPuw49iOFeV7hhOElRszhl1r1xFx+pFuaDbPtHCt6BVJyXY3CK
NjY+mNweqav4+BW1qYLVxfUsm7Vi8corLEqfS1b5viGINnXUapKJoHEqBAkL2WmP/7mW2JBg1SQF
cjrV8aDpawWUK+Ic5wJQfOJBOkR8EFJPhM9W/mOwd35287ytENd5Jjj1aODF0YQA5vf6huFpHgj0
7Dk/JAih+wygvhYBGJNuFMWlsSZZHkeH7nVqRXSHnuO1lkkjB1Wk+/bNrDFVS4Lm2AS1uap5umPX
9PbdVtKAa5tMK5+3yCMH6Q94fuf1jYto2BmTaPmtGjYFvEYy6mEueRmPWxhzDgd4C1DeyZuWubVU
9FS0ZtGdggaI7R1VXhro3yNDbP0WmTXBvPV+O/boA4+PrSs4+lsUv/CFm+DPrOWcGMTGnE1DRPdO
LHOHEvHi+16C5+YDqroNJ4KS4TjFOJZPMJJl0b1saxKLOK9zUGEydJrmruhK2Lj0xjssxlqtvwKO
d886HoYSW2dJ7A/6ZHyB6YTqzI5MAEkPE1dsJuoG6GpD+dhSNrbNRaS5PTwSxNH02c8Xq+re9vnk
MldUD3nXJzJZYiaWca6a6m944eQtbdWCKlIqOClQjdbjzeqqdEzwmHygNtFrrTvsgW0+WxxLtz+C
lEjBI0xKWhE2rlFcx7hqJwXN04EdgS2hAyNv5aP/+ezOgaaLHUmNhyrgxrp6zuPoQSDTlcqYIz+K
n8JHE01oryNDilZcC6FeLduaq1uu7Moavyi7TVuSs5fxm57M1ZNsTom4rdyjq4180VwHR6fGxZiy
4E/H4EEAR3a2O+ncNj7gC83OAyIeC85nWOBUdhH3cIpjq3BxEcw6miP9ahPeIKXt44Eb6+zMVRsn
NYGFDFJMtyFuEXpzp4AIuvJ9rL3iu3iaQnYt6j6cERG04DUu06b6B4wPa8GJ2G0WiklL3Xt89TwS
jb8Ks8XAjuheNINnEk2Th0TUd5X/D786csFf5aSdMqNm/EZQwO343ZREtBRFB9ZOVkyohH2HyGM7
T6mYtx+ssIEWrUBHhzCfm5XeCxMkpXgd/QsktF4loOchnmpq+cLZ5AUuYXHqknQHEGEMmpGNEhoM
in/bOsEu6XokCxU6Avz5qK+n9A31AV0YUu+ZRYlQ4XoxTsg+yGdrQ8R2zpYslBpSkhVLRCNv+nvK
FCCptl5oW49vGdIudPHtED4AJmqj2nLA593jhjVSYYCJQkA5kuo447jUUJGXjsEnDIt9pcGHC5+l
AbeDXAjp/NmmXD8wgQYne1ZIOWqV7IPWDLU/QHjNzNfxiqE5et/s0EIkuLeeLzCmtZsVO3XXdaig
O4VqwRMXbtMcZEgLxnvL7F2u0khU7vqx0aGsCpOCvo4THuTtHszrzf2KCaQzJo6wX5bzQLctSZMe
WFwANzgzE8rpXBinck9qqfyV3JWz8GndF4nx5haQojvI3l3ip/aOyAo4MH2T/DUMpem5pD8b5it0
3oSkvfzgbHLtfGRQuN78SBX9Zu+1FExeS3lfJKu5xjV5TlYuXGFmihfS8S+0biAlt1Z7ZtVtE49V
FjFX69BP9jHFpYxbL6cXGYplimV9q+gE0BwN+0zNBjHf2uyArf4jArSzaYjY3x+kT3GFYSDas+0h
Yd95neRG7FGFbdpNntm6tRz06fSLTbzbSv7GYfwxB5kcbAezot/JKZlAkzW0/i3VZfaXrghdUvq1
gR6JfRvJIy/RLkWyh6ppMxfH3ksFALW/+rfrdy4tpcqToRU66yQcT7Co6EHKe/+rexp7m7EmaF69
fjZfdiF0vG0AcpL+QUpR+AAEOS5qHx0VZANaMCp/0dyPqXFizvRviRMR+x4qqraG9wD0mDYCAiHc
h4RGgUZ0rIsHlB7OLIgeV6BPGZC1zxYn4/b3InkC/NkSY+s6AxrF1leqeHw0T66vwG6g9rhlPUXl
sPDLtgvrIp/okM47GLCz/juiaYdLsu2sKkT/IGAhSMtfu8BsBvyEDvEUi/QEf5MXZzmjpJ+7j/DJ
Bgn0M7RhUcsGivSQRlSAfVRzxLXg15x/vR1LUnguZ5vaowYeA9vwrVwVvq197jqomoEYRADFIx7e
VysBsUPBq0MLt/XJTnNaZYWsZbhxsc5R1clmqrAn3tVNJc8Pj5bcTu/OSno3lztEoB3c68lmsjQJ
GRb3/9jqxDBSLKBaGf4y5Y16blZNFoFXw9GqjcbwRHnlryUg2s1daizutsqHkEI9R2weDHPVMpJ0
V8lp1/bqn1r1D2uXfL3kEr+MRtOmHUienhenlCoRdMgkRFGfWhGp6i8QbER/MCmjiVKEc+2EovV2
5MfUJSzLNWeEhMqSLIXtJW9QqVvG/tBs2j376B98q2QEq/adyzudKL8ZyGo3ya2WJzs4dRB0hs4O
XJAl+4x0/v95qrFhXyTXh5PQ2onr7UV+xE+LhFOT//ojgXznDx3WvXt5QkGp+hIdr79DLrTfHMTg
//MjnqRXx6w9h2WsiSxJxtH/+C49V4QE1aj0vcNXcAQMzhAE9OWLuFH4qZn7BijBSiZwk6717Nsf
ixlGg9Ne8R5pFZVQhebFvsYjkJ5T9eaEyHLBAD9YOwxnDznFtiwIW6fff5RWXGVbs026JeJWlEdT
tXpiqps1yIaQrfs8fRJ86wujWnE+1WE+T30ODoJQNHKSlV3rY0ZQI8Y5nBLyVxK5cAzRGPsOnTz6
uTkTinVB6Zdc0Ks9rl371/xRLdj8T4xkg9gVbqAcOf9QRyA8MsCH8oLdKJMGNaokkoB/ek3liUOR
6aoXK6peB8RFCUUUEIxkennrGO+qilo0veiJ6ZMsLeDkf4njjKODJ84C+g2Z1BVDEWK7PlxPWuYj
BaSqpcPA+AqlhbU5+13hQfsWXyP7jM1SVXNvnJfRfPJOEa0nAepVgSpZpDmaL3NSHh8ghhT/3w7T
wzb7H9x3mP+N9hwlPZ9qbt0s0WPwgbCsIJAE7WsxSZ7SA+ESF4JlWEUyWOXL6nQavkAplHljZcUK
Qu7uJQ/9t1QnHabUuvdtFWmFrXGObzn/da9aWAZjkB/1b6FiO9P9ZEJWsxFAZ/FggaBG4ifXchXW
QllbEKZfg59VB3nGW4OPfRewIOCiX7KupD8DgZkSt25lRVgPoXT3GOV7mLRFF44In42hywOumAsz
8JkTfwHUjTxwvnUE09S3Q9Mtu0OxmQdNpK6bjihnYgfc+cGwG/CuLA5KSXI6n8sqQMSd3sX6U+PW
K9PhGBBgD9N9Fdf9RUNIBI4w//9c8IsHE2tDPyNAE2lrXkJK6zw6Ez8WOefYl61FevWMkZFiqzsa
EoWMfWYYgBQz+i53nAPrMFh6il43WhQoRRx6ckmo+nFZk7yhKw36MtbOQyNj7tOwhQG37wiCF1uj
zlMuGpA8TPvd9vNkYq9WPmANSyrqHj1GCOmUjwQd/ymWuxdHy4iQUow4pPXXz1plJI1/8HzQzYek
lFAQT9tXKGIU0MMfVLxwsbG/5dYL+XkcA/3p4X74c9IcaYFy+/KA49u1rO2V8mqsijpeDOY2yv1I
Wq/evBgeR4DxavYiesKQshGEvVIP5ZE9ItSjLniWuLLUE6iRdOQvvCwVhcKh2oZ97PhSYVaR9WsS
2eDhEMUnh1Ca/UApUSzr3kpSMhmdVY4733j37bbjFM0LWwrNHPqj2tlX6Ydtk1VswxsvoNdc5/BQ
1KMB5WGCiAnpedajb6aGgX/fks7WW3rgj92OsFZlbYvLzQNsCB/q+RfeW3iU6PzsOuRo+pzmyyar
jpl0EAI3CklCZ+eZfJ/PvlU+GmetqYNLCUsUYSaaRTvSTY1677Q7zfgjaFHbKXmUjtiIqBlCQgx1
Evl7urY4z4O9azM8eMReK0rLqYOixUhALTrsXQNtQz9xIWraFHiJIzZVzkQ85o0XLvRYr+vZuT18
2n6e1yQhjYB68VPh2piKD71wuvaZMGyeXPBPbiOSogmHoBuP7RWmmrom807H+ERf0YO9LQyw9Fbp
0cj1YSBoykr9aFh2IykpRhwh5qtOodt7oTN9VR+a0X4Y2hlheYA2bU1DaqJHswFtbCt6oEu3F8CP
2lHZJw6kURrlqHqDMm2zKEjtkB87uTJdnyiPilofk2yc75e/W1tiILFjxi/OTqN4l8SudG0gcr8i
5bsEqSQPXTpR3gkyefgH6rPu9NwSfNOzNrg8rK/jrKayHLSfJ/oC1ew9WuKU6sXgEcR1w+ry/juP
GxQeIZZQzKf2HxUmIUKZbZcCkJkY5+YOBR5QEVadbA8/UylKoMxD1+EaOIGjiudhj+22kje/bWZv
PDP3dUv9xUGbaKXy9mHMSkm45xCQKFN3eYeFiGZ7/SSVKI0A9J/LJJVYvPSaIdHSIaCRCz9TUCN1
nASn6zlme09Gqj2YuJbwG72r5Xt0OBlpeAft89/lWFvXTKZMdVMsqYnixLhD061QvuKz3kGndAdC
o7WGHpSvX9A7MNryDUc5mmWanK8s4j480Kozbba18E0pNFqphkI3fKofqaKk5ApCYYTDY3FFoqX8
fdlJFsdaav9FS/jKQDamDxB/yaLj6e9TFY8Ba2LQgrckcfMKXFSajq8ubPabPArfd9JZZkQEnC/y
MhbAd62lzMGmafbP0DKcPr90r6msmmElRv/alKpVZqwzC3giVZMtg0auKchAukD5HnR2JvgzTjQx
haq9TvzyS/+81ZjJgNZ0p5OMRKQ8azZQlSAXJRqpY6OltYTtPlCqi8X4Gx0haCnq9tzlr54nh16G
YCIu8GUvYivD8ss3PKmi+9gcwsdeYd1H0ejjuX8jGj14+wc43yhAK4J7GLwU+h2d9qFIQhuQeAIz
44jj/l9aEbhoqgu0W5ajx1i1ysgOy5jz+hWh1TZeQxPBTjx00hJG47FSV5AVQ2jbnNMUzqycietJ
u/HQHZ/GKie6/15XE8rRpOBvmRI+cPXRaW/YhhmtPJrS6KtVA7ijZtbK1d6RMTKFZ31RaX9luGvY
RiIp6nZsD3Y6YlfEGIdGn604aNrp0ZUTgy4Q3j2mjbSZSv8yoiJZ0REQeeayVcc9fyxml1eS5QYc
Gp3m8ppTi+xnId0saK+WiYM0RzL4LghyU3zeCsllg0qutISf8yMZU52XLKEaNso0oJLS6cwIZ1VG
EV6wGI1I2YJ0qZx1qsFUtaqEW89XA0uSNaEGGsNf7hvKAMDHieK62Ez0v5kUCicQeSE73D6BvGeZ
TJrIkXPh869x4R/rS1gkHLeJ9wYPofWx5XT7aOu1WFeS2+qM5YQM1PHEYD/ccT2GHcJSc+jkftuE
kaQXT30jHZvA76TsVOu/0X5qMIpZQ+lZ3oJfDwe/VUyvgG5+g7fpUzQ3mBeNAHthwezLMAA5hQYv
IMNuijk0tHP5c0edswNRoLnVIF5b35tfzLpl/pmmISEzRN0o96CQ1TP+Z5ZkmZNROzcIDMHbVsgo
mF3g9V8CuJFs0Kc5vCeAKtSpKteqmsiHXsGUy77eZmYQoPGSbCMd19O2pl7wzR82lhNtVqNPyMEo
dWpz+jP8QR/s4mraYSp9KBwUYaT8VRfCzc8twUzHaMm/6F8J3GQkf2NdxgLcxDNZgcdiSMeGdaKI
7hzq/2kr6Hrv6I7UZPXP6wXZqer4GWYW5aA2odX37ODq0XTe9J81PwcPSqMR0STBAiOWZ8zJrXEE
kk5oZvv7bFRxYfIQszxBICx1koq9oXwr8/2g5fCYXZMmU2DAtcICJiE5dGwUavQHUgOK4JJJfmC4
a+xIGwmr+EMmUlQMnv9S8yoMuKKloaptB6HykZHk098nkIKjCbiJgVAAa4qeDfHusYY7I8yjOzb2
jdbrk+9ZD2Bd6n+0Rxgbt6z6jzq4gSnp4x3EO4kauRaXLV9jDXwda+8Iqduk/pJtOF79vg8yWm+F
DXy8SkPPI3fhA07s6zu1gzp/zzkzxtUPzEZtFfUWRAIKAWtrn+cRaCTIoHygHAQaFBITybi1LJ8E
BRAt/4rSu3tn9aiuPbBSBLJJuvrHZ1ZnQDwtSY69wopYF1cz2e0EuVGp5ca9PtlxoP5T6VbHDFn4
YBjZ6o3AUCyRo6ZHn7bWJ8nhOHoaanXCBjbFmNGDTiIp2CiTCtRIiX438jRiAIWuCCIXHhjnUxnJ
sEKZkESUKLJImbQc3OCPjWa/KmT8lXpGgwETXCTFjku2Kw3WmhGhr4qKD8x3EFLwvJ4hNbQZdxCc
uYCozUUJRPaSJH82FiJnviCkbJU9aCLmrQMlMbCQ0yzBP5jiMvUYLR7x8rjNtWKgHvH7lJ9Ufkfv
bwC/0A6mF4wBxVl+/lK0zaUzyS9oSfp4Xp4gmyo1ylzxgC44XWPFK3lisP6LFB0bYR75YefZ6eSa
rfuepd3WXopIn6bauIy/r3rt5Ss65AYIQ+3PZJ5idgpqzAR4PaxCnK6xWR7ZHJyUAXMvpOeR9tpA
ggYH9UniqBLlziGPZGuFkeU1KVtd6SZ36aM0sH+YsHlYfWjtrQsILig3DUMiW1IhFcB1BDCwyXkY
5kpdeLRl3vBR/s/JfW3J1rE6NevUY8bv7SVKws9DVHobQRUJd1arIX3F9XrZuCSts3CY0HcDe/zS
vM/FXGO097pr1ZVp6q0oia5cKp/4SQrZuc1xlLEWFoe/VV8nkWVcSqGSxa7Y+5UUtikAAs/+8CB4
MRqVeQvXj+nQ2BHXDizrT4/1b/NEkoOWtLpYiVC5EO/PV3PmWORr62a6j3vdkX8utckab3l1m9n8
VzNHe6+nQv/zqUlYvaKvcTMDb8VB3LXDpmJcW3mceMyg37BQFIFIaTJSRQYmaoi1NEqGAH8Uns8m
yRE6R1Qd99uEJT+LtjilG893suvnCU0DgLW9sOR1r3eWTcOZGQY3/iCIsYIoGyA+KXuFmlaw9c14
12YZlC7f8Puxcd2/o52sftDi3FXW/cOZzYSIMP+TgDXAXIMLzTMXsqdIMkCtmtEmy+TAxBY2WV7p
MHoMIarlFCA2IxEfc7hXwjbeZO6BsLRPlS4RGa2uPrqTW3repHvYR3+R7S3IoIbKKIYmM+1v3klg
4TfvWMicdbT0fdrsZ1YxaZX/NQuBvV4qyQ1yZBrHCIJ08i4vcNa3Zj2BDWEZrfPl8wsnz5rnk3qi
15FpkUsuiyySbLrraNu3GlbwiuwSMXhHsxbwl2lncN+8TW9tCspw9JeL7iR1CkJoE1P9HRIMtcPW
EbfIfZUitl2KN8K/c0T4j7ikKAYww6l/+Smq5lneSVGnsfA8fPAtGP6KANaZegH+4iNRGMp3FqYV
wATLXIVojv7+LD0B7QigBGFyQnj+hSBFivxWejK5uOmQ08JX3rSM63884YcKovZug8MS6M4vSDco
aOjK4yzpMKff6lgyRg6YR7TrB9E6hkOV6P+Fzbb0Ul4BErET26+darLYMkpZwGC31exjo0T7D7US
5jE9xCdeeCZPYp70xsUR30x+EAkUbv0u3n70WH6ci2LgyvEDi2seHyJ9I+qZKtZQdstZO1Jqdj2J
Lx61HXpw6i5sC5GyDn7SrbvC3P5/iDoCfe7+fheXS/wfrcqsNmIU5zAcvK9jdhTUJd/p1a88+tqh
++Yid5xESQP01ohlhpZjjmStKwN3ungWwPzJcSzLLvBlhdwxM9Enu2dPBzzteasLdaTQd/tEwNqU
gaUsPLENviaxYH3yMHGLhqtxbXgH0Dlg7q8GKROBYmY2xui+D+ROeA6lQaiP/kDlt1OtGdAvzdbi
s4EAaHvZsOS3/+ZJJyP2rkCrwjewGtTI0+V6ZWq/6Lug452B3KmS4l3ChSUKclgFEhGnVsTqhigr
iVOHx64BR2QOk4X1100HHY+n0mJkCs4yA8X4e2LspXN2uAf9VD0XExwE6JUrLoJVqmkmips9FRD2
rSI5h2TMNhYTAk7KBoESshYS/CJaZ1IwrbVDKvhlfX437FstKR+MNYqDWzadyxyR8+3vq1IOLefr
0ZMrO9avNLJZJxT5G08HTq+krgtN27x4fOEudPwFH/1SyvmBqgkt/1zM4GRQ9FcGM1PO6ELW+flb
gKa4qHchJzojjOs15j0iaImZZRCSLWLwH19QhpeNsYx/qQCbsRz3nYqTiTwci2TpqVbTJIDOLOsM
9sLUnwXP/6Qm+Ywxr9e4gKqv+DX79MzniJ0ZdAUd8kGqiZ1UTm6oqQ2uLCB6mAJemrzpZkCFYm1z
esy+nZYhdDj4cnz8AATSGNMX/t+hRceCzlPEbwLmUh6ecV5vzPFiivK2oUthHCzJMcCc9XGQcYOm
A7qL3cfb6feDluetn4zYrwPPYe/KUVar/IZp0W8oXQHjRlw/d8cHhkKyqH09GCDOxys7dqWXWtIh
3c50LjZRzQOcavEJhyUeaPvKPS7ajCR95vAU/Ecy+cQroEmo8dLXFuz34Jj5gLqOWyw2ya6xbp8h
F/HmT02pxC3at8E7OsQbxlQbM5kpQYYtZTtNv25WgrBm0RHb7iW61C/0W84PJWjG+C7K0t4beBzs
2fUTnqWtZRmoITJ9jR6GKxnGXmf7u5dHjyO9qmIDoa8vsGJYzWSBXmZLQ8iPWdT7XHlejXhG7/ot
dnHltlrA9WK933uNsstefYiYUqUVPQPeLx58RPz+ixr6F7APGLr0X2TkdpHZ3+MM4yYwXP1V9Dpy
A0j5dCLtTRU1iDDI/BS5k0MC2iUT+Ue5cSLqMKwttH0jcSW5UNwUODx5xSLzMV7EG7CLNVPuxDb/
j8d3RKxtw4vyHPXEsG588Y8HgPPzWl8i8giwEzhvDqgTfHzmmiwyNn9a69pJkzhR3afwblNmstfp
9JVcqJtirc3HtiHK4SsdeJyA7F9DCS0tbf2HfMD/eJYZbCZuk8GjNDcRO/vFYzIMg7R9uy0Et2zK
F3jNqTIRpAepzGUoNuePuCDW+EuI1tg1i/vQMccJytVOYIBa8eOk5HBy5/8I7t+l6sNLxLFun/5a
KDOmRLZAjSJ0QbvRhZa2st01sfXoX363jJbcc96FdwkyaVg1Kfwa38+tWZEz9xRVAj99w9UL0nDm
w65zedcbNJNuTKF6It5Kthf1CoKzZ1s3pssRB25xixQBv/reOxvvXkF+Wm8lZSiy2J64C+1h0+4X
GtzOsMc3RoaTqV0cMHNcL2I+nLiMzAgNBjmMO4cwsAC4RlgMDu1ulA5GOSsMqkuu/XEoTN0OqKzh
pYT9QB1K9sKlkdPEY+DSo7Kis34QT4fNHWIrydkoC0yzynrzKPIewQ/jT2SYME5mM0RhnniiktSm
87hV1aKHoOvQ4+P3GM9Nb11DEXJiANppTG8oW90PV3G4a68oiUnuAjw+q70vuj9KMY30WYwcw6Dw
KFlOX1tIkypEzt1KCti18mGM6z5dQEdW4LeOYa/Kig+p9RnfyCG3rEThpDEDcx1DBmSzy7qpbCwV
uZ/mp8zQh3WmDiLAgI4zMt1CPAw00/UlKRTexO/+CLjMADizwh73Gezw8k1DZi3iRCKbhQ72p8yB
XTUkKuZJ3pj282MNMTT+0WxPw0jY5W/8DilnIeCg3TCHjFDjvfGd3dAezTVMoaY9C0z5y0ikd5Tz
KISleGjmexOYcJkYcMFyWrUM3Crik84d2R2yDr3nRo40OWhyyg0u+4tSiJXoAX8mKBvIfNgCtGnh
fJe6J04v2q9kfa04irsjFKSTZfNKypNe+Mxj/5o1kbuJDj6paMcIxFpsvO966YalTJNhmQA1z/8M
7EPr6Ln2sA5Z0zJX4P3m2zLeEu9j+2v5GbZuCMgoowg6Kc7k7zYyHKkiGfdH7wICUlChQEO51wml
6oaGKFbyKq1DrZVQVfT4rerMbQ1lkv7OaEI1SQcc6/yxYaTi276ta/Mciwrz4/i6dDHS81XaISJS
MoFoyq7Oawyax01bUZGV5XLK7tDiKlOtJ99rMGwbBH6zR6ykERrofs4uHKSafmp2pkmocIIfgBPe
jmnMW0uYTmzphwQA69uOSRIajumsI4GzZkFRA9eWP3tyam/gIRxnW629OJFjnPYmtxIZQmGk4TSr
nMoQmAvf1RhCBuZNCglZFL/ENZvTmM/Gd5mYgTebRnoBbVMSdGRyL9QYk7beMOIPcqIhTsUf00pE
y3uGCVNI4CjpIs6Gm0bDCaN8b+3jSV7lnqBW5RFaqelClWQ2S7rDiSCJNS8OifArCU0/JDULA5tv
XG1P6iyJh5Xv80pv4MvRKgXBJBtbQDXkg9inOh5jnWwOvtd3lAQGCX791p8pNONqKy3VXbkkVj19
+QisEgirpKfMMUvAJKm6af3FfCC/AclymiNR4L+RvfXm0bLl1yuad0/64QYj6eiwfnJ/lTUm/BYC
uHybH29yAAOpVzj1RoBX3i4aNu1Mlc5nd7QWJuC52DZ3ptrIh/gHzrYJGuzxLGnvzuE5daQ9MQMa
77txu0WWRMffzpsGVCg9amPWfODADTjYpwEaunjshzPLitJW6aLVYfg4/UOzHPZedNjwkkCNdD0J
jIFAUcdLFdMlFiZ3gWA16rZ1WFVNL1J4ZErRrmTNgGFbCtQV5aNnxkOlcYydXMW7Z0Ez6aQpksLj
jhEEBgbOjeF8UR4EGDbdDH6gpZvZIkimRDgQjeVFHU5ys9zLabZrv3LDP8/FrYiMi7wmeloAFKAL
QGyaBdkTK2CD3J3L2QAVm0Qsht/M4gS1zBRiQLphpQDSJpmzdoa5wDNCWP30aMt3+A0nYFULOFv2
qFeQhtc0Lc6w6a83pSnHXBTq1BlJceVx9qSmzplUxq+50dGhHlOk2S8MUF9wUmLQerjPLA3/65U6
I39wh7Q1mYKLz69JMkxuT8tM7wpPRk8ZVd+b6+1f859bJd7MxD9xSXTynsyT2/73kjV3aeAUP9QU
wRTcR8D9/DiCyq/ITIsgcycCmSXaeXVhlqILtUH/alXW807VamG7A85zd3di0BkFhUrB9MjH+MkL
/LDVzsXV0SpbOnz2SlntKBJs/56kJuZvr6fAcqOqZ+2+brpYdzP8NLxIRyFQcbj2TGi2NX9pH3aT
L1F4vtahf0LQGuLmRcT1OBJZBG5YIJrGFDZD0YY2ZjY78hrEx7h4TglC9ZQoKVlb0/uYeKbtstMo
Nr/9N9cIj9SNCjPeWJ8/jaq2+Sm2Dj4TfuALtQqzPPplht+KGmga7sDeeoUPEhPtR0qWkhqKv3yZ
Nlfx6EMZZFIDoicXhWuDkAHFyGfF9vKIpS3Q9DDihEFhwj7XvCGFsGD1/C1nEZp/W4l/GiBHfpx7
CIV6hLeR5r7IB/P/gfJpA4B3KzeC8vfdUBuJGIF2nX+LDK3AGOb8y7RUrhopPeijtsPpdHSyS2Q8
NqA3igTb3VLkSx6SbOBccSCBRPTU/NJ4xdRx3QXz99pbHADp0/9HYhI6ZZea3MmksbVsq9BjGmSr
TaN9kjDtjNPL6L8F4MjYnEyM2nnCPpmrWUGl3REBSkPZZxxLjAC4AiPAd0cxzOW5btbUJdYnI6wt
iETld4e51mVJFkaLAQ2nP8WdJ2q1FWdub6LCgVFa33BPg5iMGFnCC7ob1LsvpgR5fLkBQFbiN9yh
bBY8UaPY1WSGWpg+hktpJY3+o4JMLEXiqRmFZABCF/6XmZDf16AHBUgxapUl3QGEIbZ7aOt+zGgN
UOb1tjH5XoxPrfU18usrJjoi0EiGC96355MZiDjCtu+KY3LfuZjxYR52H28nTaOlD4Lu1ax+NxO6
6YIRN0GTaCFo8Kq5iaiRBwSmIx6fqrFRwiQv5fcZZ9c9NoROoKvmKFaxiDQ/Jg9ulDIt48lUHyLI
+ZdtFtYRJLyB299cxrLbPBNaVHHoO+mOTv/vs/UkgD6UrZSTvuzJnj87LH2AafIgLV3rrbljQCl5
FoPtfGqHVBqPiBxeIXeLMsf+whBhqRBbkujK69yRHUDzQ/0BWcpaG7sA4LL26KwBgf9L+pqWLLF2
JNgtH5XOxyNeO3/MRzANlAmYnTiNYfTVoKTf5OZ5X9IXqcWZljOpTZ41hNUXmE2qsHf0DF1Lzdrj
Np7PYLJV/j1WKpqnJuipQZagQ8Y2ctN0ke6rWK6CBqdB9ULtQc7gjzvkZjRAmhLUtYCmhDQEC/oj
nyqy/19jl//oKGT/x2clO3sfoSzopbii3HZrcXVL87Si1FxgU43/p+RjFuy6Lta0asPhffLOKzto
gmQ6MK1xp/seRlA7UZPt76mjpBdrRcKFMfeBJHbLpkQ8WgDQvEIIuwpyXBENnmRjFXEwhTbngS96
M+2nQnCfJXai+JYcNegoV3/E4JZcWVU+pSgdskevKU1x0Lew213GMkFy8aERyMr0OvHfMxr+Kmg2
pglXaoUpBlDnRGuvAwHM9ERP1wgWna/Ev6mEB5B5N9qNA0VP59CK5y7iNHpx7zJwwussT+G9qLHT
MnX0SGUIBljtyYmKaYgmAuCNie9BpsxgVOgcUOQsS++Wy7ZKHB1wSst7h9YluSiR0JmoRBQ+UNam
ZdWejzyYEYN6wQan+GEAETbFXpg6Q069llb+NVHLOuS6CFoE/9y7OZh86GOKPNQmUSLfK7rDySU0
OMdkBh5AQjWFTk1IWBMNYGxbmi0Dkg+NihEnB5XGnlxh8VNzvwz7PwnUS9nhx1omqGnIotxXKtaR
Cl4O5mQPrFPbfWJPEd8xXUWSufdJOUv4M484jXrs8IE6CNMrtS5h7o6BSwJljNEwWGIOmVd7Ojoi
ycxmjWSrvZ+205HUwNi8pXyLp+z02s90PzuTGurpg564Va3AxawiRtc7eij7fwPqsw0b3bC/Xd0F
xN8EHg+2Ti487+LZ5F0S6YoGOZ9DkI7XEMllN/GVBG9KeXXC8TtU638yS+aNHGYzIlnCM4EuL5y7
vQvZ+1ijFXa8KJEizaooZf9m2Z8sGZj4gLgUFD7p+pDkHafrZiOHI2SxFcilZ4vlqJHSr0cYPWDo
8lIN1JP0T/8XPPj1gLdn58D1u1wFduhiC3piCKMDABRZRMQhBZhJflr5NEwtQTo73lbDXsX8E7hC
JPjrrVxFrl3u6vu5/a1/PVJmweE1itL0ebbobcZ6k1JjIVDISMeKDR0C+g5EqcRczhz35Qs19Yuo
0ETj0qTdRnuK8ABbCChcf83pAQP7ttjPkokNFtoKVRUPBNEmWsOzcu4cp9xF9Aea+noYuiDQj+7E
OBIBnd+crjebXGmGJs3wA79WdNpQieQ380h923lolBCqEi4OFKai3mv3EGh52ZKchKVq6Eca31gQ
hQB1tQy/syDFb35m/1Uj9mu7PwrkZ52eQ2EtG/8KcC0E7R93SguOiW8jXrnxPS4XHumouuMHYDZz
Gg/htYy4/x/Jme6mrDvJJ4dKD/PDkJ5jryPTteoo+w1G9P4cV4hJfDEmT/9s+aUjzCs96zTIp7pk
shaBey4tSgK6VNkc4XKVfyFgePaysH9CzJV1hyIhXakD1+MN1vzgu2khdA60BQqrqAggFwINIaxQ
FeNTg1ad/hTHP+2n/8Sm6NFFwVVFLYuGvwJoMulCvpKEJF9P2sr2Lfdiqe3JB8Z5JyU7/aReq5VZ
vIh/OHlPWG3EMptAcYvEvRQIJG/sfve+F9uve0rRYnbDkc52pL6l6c25fiJFIBMTLu5aHl5moV6+
ov77kWrGIjVlxZN256gpLYJ+8pqLJ/gvm/okQ50Xd4+sATlGG1VToUxDMXuukNSYmbDzpeTLE/Qb
MBnY8H2JCK6We6S0WfXGwTCoMdmkRq4hruIK+ihFu8T6aWjTmS6pXRhajtvm1h156oDzRNC4aJ4w
bdDUSefZTmGD7SxdSHwFju2QWadHtrV1Tj95lIfZ0xQ/oJsvmURObmpcDNb9XaEOSfEpi9nJK6S4
U6N/2lc62SvcKrzBcCjCvF2w8R8h1fYNPa9ceO7md/xSespA5CwmUgb6oRbIIJaH6dc79YOjHX63
XiIUkuJ68oszrR1YYsnP6jsoXJ48wAw6S022JGpJyBINkr9uPmIDt+U7CI15DvvZpvf/eJ/bdXqL
HKQ/PcdhpJ5y5A/I3iRK10KeIoCtCA/XZWH4VKFlDjwe/wv6QKF4FhEMd6rupK3FhHevlgwMM+sa
p1/nH12jYCsm83aLzmTl3cOdU0/QDle1kCjiXezOtR6LN7qUpEpEvBnbBv4O5v84jpZXvFzBKLgm
cvJE+uzKNrMZWn7VjdOLNojhXi3p36+5NXHhz6SskeWryH4VQYVL0hUfltzYTOZWeLwlbOc4VMQG
hQ+Zpz0O5UWIFxMSqFQDuFC+B4Je8WKjVKTcIyrUs7DM6IdyOVtnbV0tLg7yVczz8dsXj77xXctO
up2gTeoJqgbFD0mHmGMJEXFOL50i8BDbWQLvFI3vfkJ+iPnNBsL8eJPYjw7H4tzRdm3ki0G66hUx
X4IhcQ0wJSaHhiqc6kkGrRnAbOVB5V1myxGXZ9lWaDEJ8hNcct939HGnmp4y3YkK5K5tl0Hs+WZr
Pd/fpZ+jJOIs2LMK7UvxEhTynYIm6CirEfHxRTTyqYaaX1EEYWnL69kLQL35WcW9jafUNivbrDPe
86Q4K+lHsn22eBG5MF+hCmwxVoU9kcLmj5RKf6Bqa5A4eakHIaEV5cLndReUanwSDMk72nA+DppC
G+9cQt3uVgHcMmJ/4CHWo5mc6bGI/lwc5HTLnOx744TADv06cetf4ADrrSNyH+wQEpvbilVdewz9
xlmrAeD7SmlUZQ/QZER61aFN5MdLWSSF75Rc4k0/w7UwgusHcRvqe4b8kxTPMA3+HiFI4dJwaWPX
nvvv2oZidcGmkvbDZzoISjTCEf1WRss6mTmwWKtNUPTFQ5amvvj7vWoDkBiUN0mLVPx9HfIwFAO/
2iGUcL9vN/ZZM2nLHsamMI1OY2EKc4l2epr8Ut/rJMf4sDDa7rlkEdcUFJFxT7S8dO0iMd6qhvXr
TIOuiwpavF9wRXkPVd/lZPZkUIvvVmk9o+C+caQEwVZ+TvgPYajy7AMEsAmKp9PJm2OTDkvZkRLt
7N+XeBlgU8iCNnLM5A2sk+bYCcu6c8KATPhQfFHU+ai1dXddkS+Tx5OW/iYYcS11x5EBN528gtUO
sx6A4EKA5LUktSOlMeuXgHsKcr19rZnUwiCNco6HRksWH1O1KJ1b70OvnDVrmFVdYBuo8zhI25gl
KzY4ObkKbqo0Eb7JSwj80gJbp9dUL7heIsBD2xa/5Wn/MnKQqXfGiE3neBmfL0e+2DDQ86OnpVQw
ltu9aqbb6Ud7P0BSh36swWEY0MKnK9lo8ekTYRZ7H0w7FPESFwWD5gAKTI2G+AKnj9t9+uRYwWNe
87UJ0WhOXwAaZK0rl0N4M7V6hFq49EeaWF7gnHf8q/nlCkNV5zKWMkqL48pLdSWNKJ2Tn1SJvweF
GMnq3FF84xOyYbwMRYayNwf2y19qVWEhT//foo7y7RVoIXo7/ivevICEtbYIVmYPtLZSDpfpc2wr
pERd4kY7En5fhhbRb3hVPXD7sU6S5FUy8Eoi4Iy+Os6b43gDUNC8QMNNtcbskx17x0bjTmsDBxni
xqoO8mN4d9ljKqIWo+lq2hV8SH5F2BBDw8t8EAXoTPyfNVhi/xlAg1LLfcOxKyJctPBHdeMxJxOo
tQ1ng0CtaZQ+WxOX4xeK0NjOKWcR+KeyWJrFnGrtVlaSwJnaCrTpmctfX3FyCHMUlS2tJk10fKDS
mAbwlU+MFy9VRPaI3e0PRp0iN0xnGOMmsy2KbKGu6tl5QUodRcbunBPzIo0X29ygzEZMds1OhZ4s
YYLBekfk4JhQorqJ3BS1Vc6Rt/ONF4XC4ZS09Op+xCbHl130b0Yxpo31oEJMvH0MqHwEUOL6lh/l
LpVIT8Ybmtp7y+eQkoVpprHxMeYutZiDQPCK8Ob3yGqn5pu9xlLWllBvGE1DosSIcZZfvyN5NjPK
MgqI0AMLPFC4ws9an/P/y9iMp2IQkR7E/GsFBYbW56U+ulhJvxHdNf1/xuCeOmploFV6it2bcOjX
D1vcbYrWDj15Iz6a6edaQxjLRN2CGRV9IWqSmv/W2+qTCpuCwL29upgbqFQwZySq54OhTTg7FqQG
sqdvp5hRIpikTi2hXAGRs8hhzbVlI+wffFH3S6NeKsHjurxcQQSWivWpwkMgXWDJX7axzX0yBeeX
ysqsm8kZsU5tUUhgyUhv2arvxIW8E6+HsFMyQThjOFVMJSw8kq/ueWnSDpuZUBVAJ0uE7YJqHYon
UQYgIacmNIXOpvSfAzcVTq/sKDmWRXGUGdb0wgDnDZNlA59Y6JNFZX+VybK2aby+huwffh1k1csw
Q4xN9UHqBKhTFrEZORPepK6mdPgPNAhOYKNh5N+UI4LcddcExkdHiIpvBtCHa4McUVPpltVE049j
E45RcHtPM0H2FBCXUx0TnTM2+pXuZ1wridqh8tZAtpRp7SUSkHz4CPc88qlHrNrXleuZzWqWXAbl
dQG6dhcBQGrZSY5RyFeVOsfKlsX/RllLDEiin2EP4pILYcvoICkHXDrIt7jf7S/44TODEkge2dlo
dRaI1PmR0X2jCaay3U/dg7ZLdbVCrUwCLkC5EHih2O/Bo/9bdU+JMAz3I5AahM85ArgF56HCfwAw
Y1R5/mhRG3MfaZUyP0Dp4uNfC653f5oTxVqBd36DXfaee9vOedV0u494ZeoPOqNZxx52BQkzDtpL
grF2xonop3hdneOxlakazA0WcqTSoZuzfYBYeYGtTj+ptQLoVVeMcbLjAFG2cDrI7APuediLJ8QO
LtI6qX8ZoavaEhIDb1honfRKXXyl1qS+STzqeK1VS+hORZpeI8XOD8xaEiv0f4PTqO1pni4gluUA
P2A/0Nx3NcgcAvk0ExO7T68Mpj/gdJ1cd0DlbOeWdbxuvZvLDvqzSvxde5sR6tGCFAeIYNDmh7te
ecBR8xe6zgrdWJmxCuzZno8O0z2UxXVJC6HxYP0Ne4dXNZhOKpXCOpxcGhp4r+1FbsNeCG+Z07Uq
t5ysnSrcF3LHZZ9CLFoOkHG1dlIiP24XVhwr1d0A34fqQyPC2KEzQnH5CZkMUHtFD3cc5dzWunUz
jdMaxdOot93XPmCAsduzNHv5jlGywLqOKjeaZ3Jp2L+m2dXqFswmJcLQ+kgqiL9iEIaYlKnKukWf
yScuuZmKSx+KyRSvwbInskax1HAvQQk3Stmj2dSAwbc89+Q7gC3eF1Igaa6Sepg4wbEqtHLCJ7qe
GMJkZse+iWAeE9h0YIyB50oY/As2XI5uhXZfBzgdXQPjlINONPAzpXN9aPoUS+pzbU3wn7I3sYiW
mnP21Trds0BKJCm8xVVKwPk20f8YXHhj/zCmZyhCj4QwVJ+N6+hZtDVy2exYsufDi9uC9ODbS3DE
ws9zemY6keV+Tg2BxtxWkMY6i4EEra8IJxYpk+N3ACq6NLDgo9h3xpoYyQSSb/aqbUPEU+XrSv/j
aiZVXYBoV2o3K67jjJpCcLN4/Cg24aeFLhoXDCU9V146CItvQqCO3XGHI05SCWptX+cxio9Y/Go+
E7JsqLVnxm+tPc4dlL5j0hf/RKrXm9x5zZovEjoIBZa2vSP+IBkCV/jDuSddJ+rHjR6X7nrBxRcC
aDUNBEzochWvQE1BYNaDni5pJdklT8DME+l3GYm6XFDxSsPd7FMVBYUeOasJjdQqyJ/yWdSDdPGX
EXgmp7HrxPH2yUIImaWJ4Cy2zWCi9AaTrSm5ML4O8UaVoqESRsjx1WvqDmEstVXBJ+SRj7OYySao
HIVDXArYiGenpOC8p4Fb+ioQsNwdH/WzL6edEzb0QT9Ok3oAjKUVwPkl1oSeZcPgpi5r7vJn5Jxt
BFSgnrX4u7OZyUv7JMIIcMjYWmB5fK7SsEwJ2WAZ3plQphqdEpXgQhJyKwOXv7BAjvEzP/I3yrGw
GuVNZEo5Dp0mgsMXHDL86wMvzEFLZeUR5J2gCrAqQ4PVizX2kq1mvEFNVRntRY0Tzm6h4sxRNNnz
kxCtqdH0S7bqPQSAamZyAQHUbaohb2fCi8i5smTpU1sj7pcyydVfnU7koF/ajft9BoDiSsbNpFPS
TP9wge9ife9d0kw6K0krOQvqp3SNSyDL7YhEqJJ6QryGxH2EzfzFR0flyHKPxw0b2Hz0cSrliui3
AwBYNMm1+hABAVGM3fTRyhftlLMoSKgSeTt0nMdHFyIJPhhKQiYBmexmeDp8iAY3Ku4ww+HwUZgx
BEYZwHdz6oershIPuYgXOWS54mNKxVGPaCRF8H93z8h5YBNlvUd37a7uM15UzUTjyPHb3rSn6RkF
oOufKKnQb6Ukt/qm9JwJ4PBwPJpmhgOBV9htpEC/Bor8g03MvTqNnR9Alt263OlM3xdIxe4lzZRQ
9g40Jo229x3gmrwlYwmJXuHDXjMds7SzcNxVqYhpQ2AaKeP1hq4b3fqCgxleWLEqNFH+QDbAEnBZ
dfyXsBedMJU+GbWLdlZbDNGGBdyVnIrWwsQtIG+G+d413XIN5l8y1IWcAbxXupvTonKGDVWnJCk6
41Lvonq6N7ZZIoxZU8+YkkYTIqeOppcXhFVHWT4EiQwzjJGAGk4hXZCpJsWSTa8LqTp2YzoE3ha+
EHn4/KZOQ/tCTdWzBq7RdtNgTHEx+Gw/fDuiPN73+yeIp1556tgUPyHzXyEyAVvFHP9l4U4NnFbf
H17Vtmqdv8IXstik8TdFS8UDXhh5PWRT2yeUIMFyYqlkl3cGYr5GJfQsn1GCZ7MAUDMTQ7RzeEeC
sleuHi7Dm3EmFFIkDvz1CB2k7zw44zoQEg88O0dlXjsKrabGnfL0EgdJzrGOp3Yy5pHqQ2zNvO8e
e690RenRDXEv1GjWA87mum1OIHJ9/1mxFmlZuiWFSy3yYlFE2p4SsSq1LnCYjMLtMp95DVQUjT89
OZE51RyN4VmSRSANgPIn6rbxDUCyRFdr3dcbC+8M14Dw0xHAfUn6YEZz+/qqUaAVolzOJz1L6nnl
OuH0PbRSkhQWROu292kjXxwrTcAIr8ylPigA4kkObBOuOp/T6CDNlFIrikIc+PkmKmMqTYC9wOsm
1OlPmZNCy92mJlMuML7B8s1lVtphmXSwzOtYXKyuCdo1vSG1bvL950OZ/E8on/bwpELRVymaF7+T
z85sVqIUZh8wcoNCFZ3wO9MPWbAPcJVXqy18Ogk0B8XMM8YLG8y/fGrr+Swj9K75hTHfFe8usQHv
iFEO7yfcIDo9cyeiT3vX3R1cJ27+u77DKlNqPIQjWJj/BLz0G40xVwcCMiuzJh7/apbNJOmCdlXu
q6H+NuN4UyEO2TlGdNxBCKU2OaQoIe/lcfge/l0AsGdxkq/SgPPhiX5dxh/pu4FmnFqjc/yVpiiV
ekNTMJEG9/BPbhLy4r5ZGAwPD58l65WZA/BI0CdII+cqp07V18gyvIDo6/2NkXBH5JoEZYBUmNLv
WQW9wxzfgOULX8IK3qjnNwoa3AWeudYLc1troo75T2Se/FJxvN7Z0awOF91kVU6qfoePJ8F+nWvA
DxVGeqBWZLb3Qclm/jnu353s91ZI7MuEbmC0FYijMJS+MLrytp4u+rmLoWrUxIbUTPpf6mukbZAm
9k+p0Zy7LlPzNq+TLDxRrgCqrejCPoyYU/XS7rvHXYWrLIqvgMotAO+52XiVnwl89P6n1NReoe7l
NcXz4JGcmto+8mMLfXKw09sa6iSajnFmbvUuC2tWewWnv/J2Q4oJIDqd6tsDFdXBEFboJTM5T4Qa
C5dzNeoph/6pxQzsoi4q9JSPs+qKH5ixew5ysG/VP58O2W0ChBhQy5VdMHZg3JxDV2ogLwIExomd
hFrF8tg/CYZMhuEBa3onKIy54FoC1c13pdkYnpHfCLVw0ZD3M9jTdoIoTo5vNNjwPKHrD2boTpD+
iDUzQcOBVooVXrRPHJz+mHQF5IlFpAKZVf22r2mzfoV+ZSxhUyl46/wvRv05gq1m+onKJLYNj0UC
qej4EgR3SjYbaZj+0eITq+jDH32wpUfBnQc1r7wHXBkoIVkFNcOy4TNU1qqqd6nnnDmUtDXPZ8qp
6HmK2qeulH6Dbgconl+PxD/22u7FiHwTt+Q7/HN3j4NSC+VagOzhe0DWBxNtTXtoAAOhDxphkhNn
rSmujNRBeahOCfQBORCNSWQ2IAjGOWmEOUPXXrJxAuvMZRSQDXzmSM3UOq+Xpw1AT7qAKtQNSL4+
D0ioLzCGLcqOF3jjgsqVLQU1Jt9icjEDIbbTiyC+pwjx7ouUE0QRBN72Jxh62QoMmqtNbLLXgt+f
XlR8qx8tUa8HNSNzSf+Rj1DmxxYaVSFhSiEARvbt43u0y9NtIqSj1UiEi/qFL81njHlkC8kyyVfQ
nt+lQk5rpPvvupKd4xM7hCLrrHMQQJnLisjWRREsQ28WgfnMrCr6N50586HHjU67UKkhbLiDVzxk
z8pOG5yQyp86muKxmTwwrHiu9yzHWwp94ITM0ORkJDvzhPhpvgxyG4h2qbCLRa00R5NY9QNhBsO5
jNt7jALXZBWjiWIkV7WhpIIVz096KEgT8icAiJFkcz4VD0fTYTOgvpV4qO2i/WbFfoqAocsWeiDe
ckmB6pctXz0jjHbDUc3cBZBX/x0/VhkbUN5SNwGGdmSFTkdiEMW7yur4dxQwgapBqV2NR62ZaAYm
YiCU75+Ma/5P3rROlOvONew5YUYrSG1OwZtKcLZmefb+/wFNMB5SupM0frW7Ai8EeW10asi/DgFD
ChdeWc+Ilg3TNyWrNCJMvjT1W1HjdU+lDzRbY192tK1dhBCNTT5XDFT6z0lk8F+p8qfaPgNgiKEi
5M+DwjHL0C7Ud8IgL0lHHezlPM9HJDdsAzix8BEAVMzvEoYN6jrxhIVk92EoU7rAmAxaW6WRIPA9
t0ns+fD/Udo1ojIZveBerqQ2QIE4hM4EJ3niqniKKg+0iN8J3LxwH0sbGBrU1Jn2Qs1KfTu/jAly
7JVOJqMB1LGlmCEFujDh5tum27lA6r5iQQEE+xeT4P8g7Wl6eh8u8n7JEIUg/CeqVk9AsMk7pBum
jwq5puGgfe7ofCvLhaSOJP8Qq73Ah34dnxpLpR8w7XhiiYpxlEkL06WnxseKVWdDnC9RoCcAWpEx
pfRO7vjtvkl7gf7Xa2TdSh6xd59VVzQGduIlMNSlWilTYN/JEiO3zrHdI63gGPKX1fdU2t2leBnH
t1LQUIjc0WZuhd5NQd0/epNzXO8Cm1P1XuHYDylyoM2vvD35fJnt2X7lfv1D9KD4K1XTr3X5m3Ny
SD5XwutbXTxMvzqTVjsLm3nFhA1+GJkSpud1wTdFn1iwHPEqUgYIEpHpA2TrzAvafqZuij7YA2FC
foBhslEQep1b57nsaGPu+LwFaLVOQlJaXp4FB3QI7eEQjoeY1exlduLlKfQcS04cQBiC2Nd1j/sJ
0HmZZYe1l8bJt5r/nP2GvKrMoMgl2J4Eg7A6bId0nHey59DRZpfwH0R0JV7XVielRwksirYCVC8/
BFS6TsuICFdazGLQ3W4QdIFxBAGjDCdxEly5m0NNW4zBDYGgAEVyoSuMhzYXFiazz3xW2SGqAM3/
fVTpDRkptf3PHnhhmO+tTrSbEWD8rcd8GiLUTys8MGCrFVOgLZrlt+U9yZnmBaIaAPPvpCQKj0VM
bq1ifjXghv/m+RNOlTE+vGLeT/lS9KiVVVBW4Gn1lrpxjGsdU2Lk69rhG9TZqlsGG4D6y63SDenz
1cANLAz45XqP8Vwie0rMzOQ0ZAm9gEgUQ1ecHrQi60fPumrVQ+8Xcutbu46B5uDCdfmi1XAiK26H
03qaTrq1G3DYBHgutn3AXKEbWipW5ir7/9aFVoPHdHs0lWWVaxrDyjhUb9GAleN7o9nM0nn8D9Ca
HhDxIWqhaPqKquzXSqj7tGitZA99GVS9tHrPK8DU0nsO2cMWPDyuHx2336jh3wX3JZ5E07c7WVBl
LD3yvaEJfVKziWWaD2KTSj9KntmxG7zGmugTB95uUVTSglY+wYcn9YO6Db5euMa2KWxyva/J+PSW
YmrtYqLZHj+TtcLGs/Yiftjh4ks1jCfrLqe9vIhbMTP8wJmezSnRUXbJzsQBVSSy0H/rgVltZe5E
b4s27ltQMXEJWQsBU1AqrZQXW9tJRdOG/pf+iNDS78TDBzRx6tCgPiauVyMf4f/qmoCSPBeNG7H1
fRRtvYJIHqd7ePHb0ou+p80EdPQKacPLvXN40LAvJnT0SLXFiqEL/0AYWv7bkqw3JEJhPkiejvnR
lxtt0NGTfG6NVS+YYKMQpmGCjaDjnBEBuA9bPzRTZkOQl/qmWpJibBHEbyIFEem58i2KXh6rLZy4
idAKcuyJELCNPLmh6RzJSd+xkvlZ5HeXM5NJvuXM0vh14alMXb6sJzJG+1rCsbjGrE+hw6mFPE3A
dAu30Mvv6h6ds11ivi+1UjtUw/nJTvL1vrfxdw7Veh+jLX+184VDZQ/PDu+78fv4RTRlY5b/0jjx
9CS2SB7WZ5aAyK4zfhJ8/7OAl7TIBELGL9ST46Kea4n9TpSjqxz1o4ok/0bomWWpuY/3f10nM2yR
oFJakyaXiq3VaTcqS6Sr/WVLdmLA2Y4RnOOuYPnHDxb+JA9476u9etuCOCZLo+nUYn5KWJCTM/mU
JUzoeHfodFysT/lEUItP3rC0nNFw6SVikve2B7Npj9L+B4ctSEzrNeMP13ubAsMxSP1PmDhWNul7
Uro7iqJ9CTbtDo13wAEmJsyXFLApS60bSSrxhzvXGkPpg5EX0GOEwuHnZDM8gmT9ZtcR5dDMmgMm
67b47DHnYKIdVdrR4y+/3IVuVJDwaYGqk/zk7/yKIIymfx+McOD2LQ/ztx9VD9r2tdP9ucg9Vc6E
B9eZzg8U0O2doWi78c8wgJmbvVUe9EHATmbCJJbAoSuyW0P6l8Sc+KNYPIGcNOKbuWvwn3+eoeXw
YWeu9pZWaqmj+sHohMvJCrTUiyH9SXfCGBDIqSm4KvgV3kgWxvbFRmf3qcnU9s/Ba4X/1eP88MY5
Z7o5um8hn2Bfgs7vyKDFWfolaHs+3/+ToZBMCy9pi8jh58uOH2MiUy1Rupx7ly7WNNPOyaRQGltN
OeuUtDK+/EEgspsxe3Q+VjcKISHkxvXW2RG5bQso1GwpcfPqV22hKy/y7LE9AxdXVl3sV56NbgvY
32GRL7kJbCbBlC58Z3FpPUa45FLVfww/t+ouTclMMSndUaulMWQ6hnO+nu85D6+RiSKYTkPs7T4M
16p+XnFGThfFfdOkMtS32k+53QjNv2VSXkiX4CfGD7S8zgomh0oLpIAankQi0RIITfOFO+MUtrLM
vn2Q2jiRQpiAij/W/djg3x8T8v9kalDJe4umZHM30fZLmFdX1xpnUVy1tXpaXOAEXEswVmr0TRX3
3h1dpFBiMSaZAv3hsGAhmVMD9b3NZWxYmGE5ZOL5r0fVdGaK32UjPWBlHmfSlgXeTXi45ZfYqd26
9H6+1vtE8A3KxrIkle5wIbJvSSZWL0ygSp45mgRn5YcJ1ew/eTBOUORZKsFubxRuRWHmr5/k+8Xu
7u4Tujjg+Zut69FFyPLTX1LiVs/o9PLWr3We/+mMRHQjE2PK3U1VH592j2JBRCSYQ5ux7aZG9RI1
VKRv+nX+QN/WJeISE+dppjC51TNVMRaff9+3q+fZ+30XCmYRULeoKPKl2uK88YLgUySrkf3qqWgY
ffu7hMRpcbeDR7BwKJfw9Aa8ZhFpNHrcBm6R+qvi8W0t5jj5LSVSfDhj9ie24vDjFMJ6EYEb4cRM
eeBOMPHunEtI9RyNlkQXcOzsMfxYZiPWp5WjhBZFeiNz3KFqjcFSKZVxRRHBNQyWEm3oJOXIdOu/
YU6Kol6KAfJFf+2NxAHY19aFL11Qcq3amVvukq6Mld15V0ZtWGNrHGW3y1gkeGskXeZ3uNj6DQxj
jWNEgAt1uyzvF6VzmjWiDcxYLRoIve9vHd6zkzUb2vQMFLacv//UTdGqAW64ZXPBxCSmSDRlSDFM
fqDaEVLhjPf6PSUaKvOvdG6HLIFO/C5kF3rQgldMSss0DGIEouWFdTYBjoYL3nePPbbrGAOnGMV+
u0S8UsExe/IoOI2y9baRIRg8WIeZ/GuiEoL01REK0REw8gOHWNYMU04cNJc3Uk70C0T9OadYxIy4
f7k8l54Ave3ArypzehPFR71vOU5q9VfC7ASbhbM1KH01g/LJ7VTUWFpi6dsFwIURxiiLEhsmgsAv
kf4/X4uNHZ9LIzlKRnaMJ5cLPgnAasglvZU3DivFuHo4zbH1Nyx9zZl8p7L/KT1zOV/uYaTrd0rh
EzC0s0pOt3yp3nugB6/U7UxJrybttvF4VYbaHoRjiWsvm3MogIOvRMUP5VsvC9+4E1WGnE7qCFsf
VvgCGVRjYhaic6UU81B9LiswHxIO4qpZYeEwS0AFGn2LGdXGojOrcfO1UZ3b5F3aBnDwy6/UKT13
k1objBVZaEWrzz5Z4JGKVbkU6cEW8cZRHnPQezZWM33Svhg74kb1rYHFMP8MjuE9odSNJXij9bfX
sr9tV1WAj2Q+iKs3hJWFVe+AvpCNmWVfzOKkD5UUGAZZcWq/i3Fq5N+q5iZQz0U9Ci8XigbMNgtn
m634EQ+k4OsWH79bIFbLEHtHVkX5CS2pL3+6NZF3kCOmXcNtrZPMzyzTivJJ2rDVeeXiW7k8wvO2
83hWbEqgQZlWFtQv0ESOb/hfYzfIYLlI3j+1fJ+HDUaZ1/oxHfCX1B0b6kfPmQ711A7nSz2mLmyc
IOPvcOzN5y/gLQlx0SZ/JpEJseuqZ+Qq8i6iqegTa4uXdiQn1HEri9g8NpBNRYjo9PyV8jB0dRTs
/I9RY3CbQt/tfVIlHXjR+bY6LyWXSfCHZXud6AGRK8QvuVI9ZRh/xxRQnf9AA7eSJkucDjhSBpY1
e+ZjAqtJJ7W2NS5Nnj++L8kDsP2XRGp6CqsF1oMKOcoza6YtRr/n9vH2HGUPdCMgjGwhYRdzdR6m
TMRcf/cDiYJ4m6uCbEFLVzHw6V1Re2kNJ4snuZbar196xthV6uLYyPjRh14OAAIg5yb7/tWgr+Kj
nEBvEviqdbRDt+Y/74L8lWIT7kO11tzv0Hfid5ffIBVm7xCW/0cW1YR8d/44GZjk4c4OMKuA+sAV
eVn6NBy1wSv8+ftDf26IsugFsvCXxj1I2udfNOBZORd9zaXl/CM8G+DyqavRIkyuuugji7MWWv2J
DANsVRaJ62crrh2MVWUT9udFY/9dcvLLe0rYjuPgiQMsrQxjWYk25Qx4+BStWDCuvMD/4BpBaTuw
vY4TVwAswM9pOPZNRM6quRj+vnfSU4Y46MSwguqI4uzsAQZMjXc4FKRbGLVuJ/6MXnK8fpUdKB+a
B3q3CIunkb9l1h7t3wsVGpM6jRMkHylOqfglIXruY0zDEZXmIOnl4mgFoVu3kMkKcp2FcJRt2qPt
blBrjQMahfJDxBAg8LO004A0Bwurp8CI2bEU/xsQ2ynWsM9wkmwF42IX3j5vDpX5WGjgVOA01SH+
u8LQrkG98zqXGqN/+0D6AUIiqZDfPAi5DS5RnwgiZd369otNPM806XRshWKiZtq2iW6Cau5mcKZg
IeTvyQJnn3+ZTOC7vkslHUbsvZUZnDZZnge2mV25s0pSFbK3rmCNmreVaNGJHZ+WNQnIjIF1Y5Gg
pMNPObNIGEatKk2V6Gm2iRRBE10Z/RgeeeCklQ9bJxQJHJuWAcT6V5nJNQQFZwCdTaG7gRs7oFaj
vxq2EcqhXS1XoYTmyg+faejdM7alFvcw6Vz3NYEXfwQ3zgUutzGU/iHgHuGveMDmZL0oZJPFqtEU
fhmUWNFlOgW5j867hYU83NTkZppuWhOZjXhWftAqemrfTt9nAUl7dnymu6Msn8imlUR6QqMiDhK6
214b5h+MalrepmDjMcHl98CtotyvCJrmGYPX5owcC/LGqH966DfrG15TD5ixgnSXHT9o47X8chT8
Rx/x5XlQoUK4qpIqOY0ykNNVAP9vkzJCgGuqkTAhMJWmd5cInFSKzH6FvSX9TYSDRPWvWsZlFqcz
mgTs9KjVotvnLBJsgldLatuM+6X8Xx9Z9hCcj8rPOuTKA6Zb9wTiCYtCQi3tPwBmgq17MFXvYiLG
Log8wve3T5TNIDG+7mASl/0fm/TPwo1Ne8tqOu1Vsg7EZVk+I1ycr8bm0wvN2xI7Wt5SDiupewe3
JAE4+iPosLhz9WFZ8TnwTE+CzTwbL3cK1YuFC7kFtPNb3+f+4vZA2REYbZYGEzgFXh0LCH/04dFb
ED9ADQhXBU35unIB5QielevVEzH3mDb3pQtTRDDshTh0mSe+fjYmA4O9G5QUgNGu2QQfONRtrf3m
95QTdgsnZWAap56bRGYZQjgkcFnM8x1K+1PwmHmQ7prtHNR6zBykDwnuTNq5Zk6eakbOjq1iJVuA
/0ek9CG4GZUEBLNmzx9jV1IuXwlIfL21FUJUic50AKCgVHHWK1PGfvuM1ef2r6ZHWK13krruF3m7
8X4LNXJO9wE7jhGSp27ssWtirhKZrCe98AZLtA5cjVBMS45sazOnkl/7bz3w/jKlVnx7YM6HIxV8
ecAhcrY/jgSHFfzJD4Vzl9f0jXumG0vex5i6tn5AUucx2mWU4ND5sts4ZiWVXa5T1Z2Efee7OTqx
65TfaU8DC1VdWmmYKNvYWJG3PTnJ+aHKz2977w2Vu32srUT63t4f3qxxjbM6FISs/6mI7bCAujHU
aXUu78S9vnRYxJ0qh6LU+O5YULqTjoAB5VRCU6+puxPe4m30Y7eFl2TSKKgsRzbuXzxsFgysAyir
zySQwMNfdQ+9AS+FpJf6u3Rro6GmMGwsytd+WZs2vOA+Sy1O/zD6DGH9XOPlNK6CYOKWAGKYSa1Q
lkAjj+Eu1GcckvzpflIwWpeFyNyap/vykrK+V9G9CRrBm6Mu1zw4TwvyrCq8fzgdaQlUV11cfR+p
McMiRYU2WARudU8HBqrKLqTFgNxgEoxzoclk6IYh/nlftd9+U5ALoyvtPrV2yzo5HWMMErYcmtK0
/V7Tx/QR5+gJLpLJ9fwKawpNXUyrZ3F9N94N9TCra6dYP6mKawyrUSEERSWT7fwplHzXxLtUpuOG
NLNy/NEM4jbkpXQVjsN/dQxAt/20AOnRma/uRtcPr8ssFeISSM2CIAkNvW8hAgXQWj2Sxw35Xm/Y
gWeDKu4MCQYSYYHmv1J1q0dMjpQOjdpPaZZLMxJYce8lbrAvU7aWv88w+zAYTB4OaMhgglXo/GaB
JLvRTfvmHtyARJZYlbrfmv89NVB7125G3D9Kyg+blcH6nXyPv2nbKxqDus0MOh7PnXKSgbWJPfeC
fA3ok7FxbsmI0bkQgAGkwQzU2uedKbEfybY5CUHQadn7XltaE95qcYbl6GdatsotCaYGOdqrFaQo
uwUplLmcqhpOBQ1wy7EKZjxYzWrJKd4s9Ojjszmu5lWNSIi8envFVLo/aTb4fAnYi+rBtt1v7dj4
uco/AzpSFtXiiAPAcjHUxDzlH83R05vAg0vPVEJloDkQQSVLSQYQr+QvKFSKCf9p4m4AXVzMW3hX
Ag2N457s8oEgANjQrjkkFXZYoNOkF+5PWJgedqLyYdIPEb1Ch0nJISiO25TpOmi7dyJm1t7eZi5O
xRc2aByQFygLqwMM5jAQt0ezmTKrlvwhS0EVCrKBxJR90GfualX+MxUgXm/oAARTZDs0dYs9ATJi
sNJDJ63cQBzrcwqVE4Ie/1CygnbPOQDgl35ztNGuRK1B/hlxxGWr4waImMCOWBLYq+B1Yjod9X2i
dSTI0pUDeigq/xQZzT1TEbNDgQfiOw6hqvooiFmsQZ8VptEXRmQAXExtAlGMneL+bKnMent6JOtv
LuennuY1Um6AwFiE/wH+xsH4isQKhusmGCc8lVqDToYv1HimNUWXgR0tt5R4OO7ACz2eJH2tYDcr
bsWjETQJn8MTdgMQhFJcxn8exwfY7wPa1JBhiKRH3jbIPheREX8A6h0at4+zOg9k9DOBkwQM+lj+
Lkr5S3vIjxSbKAYb+tyqs4dxTcUkW2KUMW20Z170WM0F494e4wx+DS5Y94/E/mqEzpM4wnv9v5ZH
a6374466SkiMAo7c7rkADQmyBsWaXUo703ChxqQHV/jLBPFjWwzGnalaFLP9RGU5WkP9J0S0tGtd
+mx8LRby32OmgyS5IIyybxwSEwFF2EtUqKKXRmLrwKOwhARqnBzbYWACaonQ7BN/2/MEHDtDSCVO
r3X507osgdu2+utYLcRrhl+WUQd+tUWjT7Pcj6GAwstGHsP1o5P87YZF+FI8oqvlLtTXE5pmi48b
QSrAjLYhWuRSt/IX5+TVLbfd7/gX0GJL6cLP6NjATXjenrb6AI/HDwu4zMOH9pDIGvNyzUW2uz3O
v3mLVCMUshTEB1GbjXuoJbkO7N5M8ppac2DQRfaWGe1lCJaWV3VzBeeTLhri/oU+i7qD16I2cLBZ
NtLzHWQ2RlJb4Cr0uAb6zSiDMu4DreimzDfgS06jlA3sL0Vxzcg3fqOabnBmHCwD6ImUjGkl8ipE
403ngmgc1gjXQ28AbtR2rz0fmpF2KLCc1tNTgc5EcNbmXqGOcr6xFUqdsue/CZcGRhJbT9Y83y4s
W9z8Gzb7wg12dxdulGGJXxAQPJTRUsLRLT3MIrwgZF4jV05zmljIzSLPSwP99RI0vP2B1FbWYUbh
kZLfLmSHLhaTTJhPD46E8k/DXFo7R4GpTfxrT1vBZuJbo1B5qmrxjM914z8nZZBf+1Qkm/L0Ug+V
Rl2gPxsnK0O9iQU1LtKmPqW3CO9ZLBvqabDKzQr7Cw+2Jft/sE91XB+7ZzyzyUMpvVR7G18wmV+n
MUaHAoIGwgrVmydmaQJXNPw88fB3RSVNmivsPnOi/rEnD/tK4ixg0FzTSIfvqMalY5rnQfUReVaV
HZibXgcglkcG84Hb8xtb1bC5B1ZWhIDYbf/IiP+u6ySveJtbiExcVFucZn0yGWLWiXJt6aBSE/1g
dieuoi0l74vdqwCfznfH0jNr9NC4PBXUNux/B9iwn32xZKYcyrEgTHf/BOMfUfzErL+hTt++fDvx
R0Dm5sQ8Nf+vYnh4Unm2I74b9m/ALzmOfDHzkssheHgrCTAxeL2u9TrQDky6f+zCDnF2aJ/RX5fU
ZZbu3LKb0mBsD1ZmWuCb4EAegqa9Qb1Ydbtfeh+9YP5QhsG0VXgzk8oRptGbQ1F67WDHjQfPzst7
HhIFx8k/oaFVInyW/WOI7Uw+zxuxlO2tTAM+rvA/W16NQnLP87cvRhb9gVVymtLclXP+bHk1YgHR
RmCRWKfiuvWLUg15y1e+axCcNrXUY1M6b4zHdYLgNwyM3GUWEpwxpFyTP6gDjKwUYO+Q8zBZP/Lr
1XWkjJOaAv2A+C2k2wue319KTn7kbxzKQ49Jz1BI0+OTqo/r87TZyGAwmMut2qGaNXomKT3vIfUM
lD6zM+uSIuDIEedieerS4SkgB2A8Fhcgr2bgxFuE5bcIJZWvKlGGJt6CB8vGxnJAwPgqr/TL1pbz
WJg60znHujOVaLm/6ut51Tfb2eHMry8lfFA2RwI5cQse2d377BIYLLlgrio0ewVsrPDgHC81G4/3
gyeCYAy2ynRlI/ma3t113LyNhXr5olpUg6umkYlrLQIAGr3gFNlAsl1u0L9YzmkTtvnFE680K7mH
aQ7mOK+AwS6vJO8j9rHfmDpYbJnKnflrFK6QXXoSDvMWZgQVmyovI4yll4lN/WyNcHtD+OIdereZ
IHpEu+TDQATEYmXko21xxMMDVO5E6Ym3uBCmak1V8PwOXqX6N59jwSAisTRwUQBTX34B4lAI6DZ0
xeM6hRqbjGoxASb44C/pl0X9BzHbk1ysMD+LhXV+O+Iw7nRcKCndbDZu7EIS/fkAReFWn84gFshO
46k4xdPLCgvxrjmpZQ875YhDTjHB3lsUbNjfXiZuJ1yRtN0e7voBKAvsfV2q65141Bbay9N7Y9+l
HP8dCeY104LIpzL/8mpWctQPG1GdGzrj8QCJTAQr494IV1uFRPF8i+TFNF+EhrR6iDeYP1lF2erY
C3RbUAFbLHuQ2sdtgeCGDCpoM4EM61zmP4EgBhRzZjRTEe3Y/o88RIjmxGLOztQA25ZSUVMlvA8n
VZ+M3OsO60k6m1m/sQIOB1zZ+nvjloC1ujVKXSNXpodTYVdb+OmF9SIN2F/IabOgP+TZxffdi6xG
37fWnD43j8qy+I75cinO27Ym2seJSlbkr8jhqA6xBbS8Q8XotZkYu3evLot6Qws0wLByDhFLUMKn
on4Pq8FS9E6u2KEln8tbhYQ9MPvx92XA1jftZwBlhT2wkmUsHt2F3NYRZylVTVfA6ZViaBenrFOH
izyR2tcLGNGo6moluvCqbB/BOyOKIzGNEh8uog6FJCJ7Z0DBex7EeqeuoydIgZGVb2AgCZML08xK
ZXmRp7+mJmM8CIMNPkE2iKk2T6rhnXE9Uf6e5yx6GlH8LirIBoInNiQFafFWs9iEfDgOwJuoGnR9
43fYslArdE7jeOq/pRIp1z0ZG8yB6kzgUhI0eoO4IL9EBsOuBq+9+HD/LNYXVXLejOOW1LllJqyF
sfHzoSxyjADzvpDAGF1C6NhHaSPNMRGAu0DffbV2w8rTPkJKkpajByKgrSzwXTg19S1jHYuMbpun
UtYX3UlI+gFydoAHW7N7oxPazXNzmnlaM0hsq+n/FN0ozexfXj7w+l0227YoD/Ti2wkRDQjywKMW
GOA971KLoAByqN4CqLAW8MZa+jN0nohMuL0zTGg423sk2unC9ewwIbgVTVwSpunMqkdu/IVt7/KD
nSzRYbaVPWb+5ODJeDde0osVE2JYoS4QWmCG75px9xz0r2BOCGl/MK3IunwNt5M5iykQqWox1k86
rWSXPUJyU6GXcuIuN0OPwDiWnSp5LL1TaQgFDo6c7bAHnZIDlzRsNLEq5Q7dCSLLAwSYv3zimZte
ihlJRzUyusAG+rfzZ8SQKRJDw/m6XdrsB9gm4TOpxZD1zCbGgmxQnxo/aKI8zjFbJsf5covMuYbx
rJJjEknlIbSsHLovAxoMKwpuh7HKKL/mi4gaXkRNPynYTg3JteY9QAYcEkH4Ap9eIsZXsMKlbATN
1skHZlXbQzZ8QyteHtzEaWpJJq6+G0I2lH1Xv7udUHbDdMTnApJoejT8jALJhA1JNpLQytq7nSzT
Vn2NRD1JQ09i7KPwRyqGfwxGARERCmWDOX2e0jzpgflVqVNkEo0N1QYoJyzKvW1PWoPCVEWWPRsE
rAKjjLQ11JEmqQ2QGx3BQR+UHFJSNPSzEHDxCrJ2n7djo2N0t6bQ4DVCAuux7gyL7vAwfqU7PoTd
njcM5budoKpe2OciyoZLZOd6YdTl1mtzMOFp+3H/GEHDUkm305TdFlT6EgTF7O/sYzzfwNG5iZNp
1D6gAXJEeDWwfTp+ABKhbw4Mhcj9Vo+pdw+ccWEfCJx0q22FoXZu6NHTa3T0It6xmmkRHyCKjleO
ShPVPcfQs4rCJMJqyZ1CfIUi5bQQtXmk+qTBvlvt7D4wEN/RKkfEb50omoGqDUMEuNg38jCTPu/L
Q9bSu/5LfXcfScEDlr7GggBEQMUKOyIAJoodwhAZzD8LWv74optcehhUJj1GOT2OwO4p81NcqYAz
NsDd2oO6Y5/foxyQr/qVgxq7VZHWToJjOTLcXEuv2tR7BOg9n0awsMq65bI8Wbi6JGLLggNIRonU
2LWu7KbPnIrsvb53GsiQo7oiJbN1tauN2xDWk5MICph8kn2zRlPJtgZQFLlshrV1DC1Pn868ZuT1
oDlO8z4lxiHR1sPzP9/dzxof7KFog7oG6arV+poHftaLTsvmrN6LqHgQNM4hsJWd8PZe9puwvM3c
Qhq4T5PJ+kcClHJcvg56a1S1Mifeke++mPZUeJG1KjtmXCCwc0cFM+U0RS5ITRVFde+xmWzBhdot
ijdiuyKe6hr7mD5enX+vincAxCaFpVGZmtr0Bb8DlFBK5Aq3Zi3GliDBrAMYADmbZ2P3ZK+ICzC7
yL6kQzcrKVInfJlAz0Pe6HKqtTHptY0JbG4fLXj4qjMl73nLdNlegRazhDVm6RqOwwbOIu/oe5DC
M5DokXvjqXJyAPey11k8+zDdGGJHKO4u6Z0WXOwRI9D0ai4b3RLZR09fWxCBw/LaI2LTeUsuyTu0
ySkdfclkRtXK05x4Fybn5S/1t86WsiTA/ZaGdGdg0hlzAe3CLBVVsRZ2bf5IOTssjkUvArkQ/Dl5
XcMLfjfNaBuAoTC/68xPEOpuWcxIcWttLBz2otWugAxV52bxP3d5+YJ1/AvWxDPPvjgkdopYt3ev
G6iUJCfDdnbbt33phMHxbytv5lT1e7wYYLmrmB0JdGhbMtmHkpQXaETygJOrRc1BVtOK0daHHwTB
yHMqnXEENBd2ZIb10ir704s/ed5Ag8AvCFS7yuLWLnKP2HwPVCzdznR5hfpOvWZoISp9a7Gg6VRl
qZxNruCOalIfSz2N9JG1W6a6aRXLycCVzM37eYUZyJdNvocGRiJN7LBH2/xsAiIjzvtM6WsLNLIh
HcTmJE2jZ7wNXzQJfmo7cravqm0CrOyFURakVMPCMGi8yt26bVblxr5dVj6PUYU/nwEogFpyrbe7
3ulJfYWTKPr7e5PB3gQJMeduyPAox+0nrWLj5rXe5n29zUQG0G8KiONMnN1fgM+WGFCMPZ56ZOKo
oYlsMFqG1SZTyP1Mbmc7s/BCDhnQAqN02vS9Gxb+TrEr5/m9Td3LhJPKVlo5lQoVwpXU+OQbCzZS
xoazqMT/QzW4726ZMIb7+xP8s7knWTbmDW4VovpR7+z4yOvFKLJF9e56VCXnfija0upASktUUZEi
0bvMXAxMpgXL1lzabY+xxnWS45s6b9MP6/wupWmeU1xOCrat67frg6UlWXAPxqj1q8CatRj21RfX
l5isozELBsVSFx3vzoHS5476QphEVhMz7C+aklTiiTeu0vre5j4Pg80mRtvKjxzIVl2MIMNgdqsa
70QP7cjswyWID3//FdS7jhTe1zsel3xl+U/0M2rd9IR4t7Gx7KCPVlXnZ5uh07Khx9mnvOuQj68C
RswXNffAt25K1Yje07zDzJbSghToN8B40w/XJC5IEgBvw4y+WbYbn+cTqlD3DwXRLzPaFusUzkSw
LLknorIsR1vjPjflFANI89oqZtffA9+4gvx55mqJocelJqbapR73W8ZXlTODnvx2LvEOxJZN/CXf
gZ6jgM9k//6EHS5ilAR0ulXy5oWKf0ItwIno8iOmxB3KaE3k0pEuBUm5ge9Fqq8YS/Nb4mawBEIv
gVCep0VLLTxn3OwrfP8rrzqWAftR763TxprXgiyd9lyThDtSCpkV04A2PR1skCR7oH+m6kfv/SPl
PZ/eUaZidr8cH/VaUzIRFDKP9aa49/rbA4eMSIgx03H3fkI6qVN21YpOAHpcCcYCLbRybBagZR3P
wdCyRsCSr0sFvE1C1T1y6eRqgt9AjBhB+8QOKX7sjrci+hObCGAI5IHdlFpw/4Pl/T2nVtiEXl8Z
+JWBcSp2T4gicfk45Abpi2qo7djwP2m0Ke2kndnZHR55LSGt1LtLEi98mqtwa1oj/rqAf0xoF3Lk
r322TwjhPSF2aIqb1cl/vfCDvgGelbCzP/1i1jzRL26fPru4hFQWGbuLIpKMGXBwgSCf1TcNKSQy
hiPnqqCrjBgalEUdfN/ftXYsACzrErJraEpK827xtS6aqItVEzJqXf5c4RBG0Fi9w/1eU9TcSNLR
pShsWU4p3GcuONxKU4wWjT9BWyUJRPReuvMcD1oFczyyqM68sdIgDJ6ZCExja5AH27LLdrTIRdqS
rYxctodtundwTy0xpX3fFFOSL86IAmdwQs701VqKiFWiM7NFnAr4ET3a/eXXwYEEEYG8VWiUwuX6
o8PxvPL0JZ1n7ZRq2ZyIHm17zWFgta4n5cFVpHgFg/bNvNI8Gb5Lgf7KqosoDvl2xHcO+Jo8Gh1F
LwnmMvZUeQFf8769mOY2m32qr1QSFR1abtX21tRoJ1n52LJJO0PEyZt0bKgrXcIOYEHYmEMSAJeo
MQymlkvADHZVjV6okkJabpwC5Ga2vz4ElIs4GQQa79mqIGJt1C3aEPKPRWipHtzTsf4LZ9cbaUCo
CpH0c4mZ+Vqc4EiiNTFYBqw8SuM90X0ewdJb+0uFoorRyNvQcPT3XdG3VoYpB6OuXKtbCCaLWrgm
gr5O+UL7Q2oNb+8uJKz9uaPnOKaIqzlWg/MKUP/h0nqJjL0YLPryxMdColxx3eExjw34bmuemN1l
R9oNXTTWrM+RXiiMOuZvRAoMa+OttenDjrlrbzICB+sjJ2oW0uG2wrxIRWLkd4Ed+itGUTLVg84j
2tUWU/sVYPC42atq9X7370lEpTmswR+cBc1iAUD97piLGLXHBsrvpNV+UIA3yewftyjTCp4bVsqp
6LV3YJFFL1sVpU9jFoThQgxcyEemPxS0qEltjF2g3dOT6AJ5LNq8hIs6aFOJQ6EQD9rIXKd2ynDq
S75xHTC3eG19Mcxqef64iFt6OuyffVMXkluKzxKCLixqbwpGoWtfJY5MjxP74aO61BS+SU4qnr/j
BN9QdlkojnbjfIhIDvSgi+sC5Dq4YT196X+IFc5pQsOQKfOv/sS/tdm/aqz+db/9CZqCq4oxyFpM
6AyQAkAKmLpM2oM2MgGhcW75iVFwuYiFADJdtXH0sF3FB9wAQjAh1B9CdyCLjbeiFrDPpIspxIju
vhikYGu2LgNQLh0RMv1mfT0vtSEvCDodLe7j27gNNpjNfE6yumiiWgWUDwK5ky2YOWX/se15x7ap
CPVRwmK9L9vCakMyeUR9QuDHeu8eJENXS3QFtQ8yXCHAY085iT3QwSIlovIN8BfApU9/tkeLEiHJ
gcUgfQ0RgkkeLump7FOtyCM7KzYtmZpuStitzv8sBTdYu80bpDg/3ZgBAlog3nrIMPJ5Xwbqrc4v
ZsTkyrouU3Ykgyg6e9xttpfAt2E5jzVDeuaiH9P47BvOdBdE3pugRKIGMDBoeqPlBC1pF+QcGfS0
mAPbs+o0mliaLz0tMphJYqSq43zUvPxuxfY8gIicibmzZgoyeTe0XWDAt+pdL4oi477NTueXJTs0
HOQEdpGypeNTkQ6Asu9kfp6vuy7EYFandZzmhQpuLnFQAI3lMX+dOmGQJ2MkUr88yFdDeYUUC1+Z
/GmtGT2vD4+0L+AwfmqOtHse3EjNdGFaLEX4ViC5BCUQAmZGr65pcEaZUDFKEQTEDkXkcWX13u/y
VEOVfw/V9tsKKDbcv6ITNK1IK+wtMIjmJ+9+93mTT2oNkL9LU6wMiJIm+XtEkBHbJoUoPVHB3S37
EaP2iR1LXKVCX60Mmo10TVmBjQcHP1OVkTeOt7KXRhIXA0HJhQZgbw10hlan8RGFqB4uVVBG1aaE
P+exNfgAxksRRS9OwANUnFQs2HwVNEbFmZswZ+hWSME6sxCK25spK0Rhft0yHzLm2wrMAha1lvm8
lu/if8vR/XjFY+aNjaluMSPIKMKab0B/e4HDTvZCAqBgcymokcApZKzk3hIiDuAjMoEsNny7USRk
hr1x/l4XSWav7/3re9HcicF0b5n5vOEJEUwT3HPAm89wDn/I/mj0i7ZN48OoeYqOq/+xiVa52nKT
qnGmr+tv2pAdy/XRuGzDoXj8CD/tvWN4PNDlo02ByS2F7qjY5wFc1QTjzN3cvA7xrC+Oide1tzv3
YmF2MiLaHvn7JJD8Bka46TOspxj2beAwVicheA9x4pUKNTbP+4iglTsxo7m4ayazgxO0XtqyJURY
K6gBBa+KWjQTw47Xlz1dSgdGvbtjMCyPB5SUTcfuiGNmq/MLY2rpuqnbM5NorwEgsLMZHgkZjvh8
GN02KyKU1P13b/aHkj+9fWTW0mESjS1g6yzu91sL7k4MSOzQmM6yMiycrIlwepLBnJVuh9h8Pd7m
pnMBsE2VCuX0WNtC775+9irJ82sc18nZvot+i2vLEPgbwgKzxwvVFGYex/hRuAMbiHNOaPyESmA0
BTbnk26UnEuif2W2pL4UFEFp1JgSQTo4oWceszsdhNfrcI5kVknPhOjz/EPEmA6EKkSu/xBOdRbG
Yw3NgDzynrLGWL2i1Oi0PY0xWTRW+3eHqe+0zaFWQRXk5l0XQfYMssxM79daYMsrZwZOAa0/XTul
FIfj9Y1BfZ1Ly1gsoqBVjz2TaODEZ73yKVTG0wPvg2E8ZR7VPYYAyCxabVTyiQLWUskxUb57g40D
lHNM8VXW9HcfIzoF8NoV54sQ83pDmWSFwa/orYn4WW/ZoZ3duF0WH4YS1S6XcQv7D9HCPRyIoUeb
U/KvG57F8Jf9i2JyvkmgmQpcqRpfZxZ33eBlt2Q8IwMjMeJTQaz1ZEy8jqq5nEaPmhoZHC0l3KYC
L2iSU2PDxujmHTWRXz3pyfa3i0kF2NPrlKQs2CoxON24NvOzAdjsfn5nOderhE8kb2zhUcpsGvXE
l7b84x/8OTVCxnj3HcdN8HK+61CsaVZ/opjue+hntkRTGj4ENy1gvSC0Dgfnkwj8QA9ZhDw8WlF6
b8cuD2KGOGTxYvAQRsJ4n+tfqn5/mnyy6B1Cl+hXTv7otwKN/qlcGRESrNpTwpYKKktk6SHALb+Q
0wKWo+9+sCgknhlMyeBg2Oro0Qiy2RBSpYfCHlNZ6KV9+G0XDSAORQumYw/y6SUZID7rc2CBIN9P
a1+QGFHecYEAks3cXNnH2OVM7CwGNXm9uaADn4EDitCFTf1CUmT4qU3lB+/gYmfVoQnR3xhxMF57
myZR8GTgRruEH2IN4Rau2ZOroaBgGRiXhwD9eHGTQ5FQTtdikSv5VhfyOE09LPOt8+SxiGkOvvQy
QBCHhyr7gwpjUfsfQPPymVAuLUUY8SKoFYesq/RXFvzEdY7EgFF1TszUswxfBUXdF9fNtogIKttW
qGMM/CrNKoZxVRFSE6zpv/3QpFi8NzPtFxI0P0IsX4B8OpNHzzTiwWRDOR7zEYYd8NDJVNjQiJ5q
59C3AjMt88A+LCqbSVMnHr7H3itQUk6hSc6z+dfmihonwlptaeVq2+pH9pr+rMylqrJv2YSlT9WS
nybwEtHZgNVdQ8KEbH8nwlwNijJjLDs/KXI3XNWWptO6jhcApJD24ngA5TRGM2vSyEThtHXVobF6
2VSMVUyVS9eh9MQHcW+bMGPgx1tdYre+rY88+QTcPIfcDxSybLq7YUAZlSn6K0SNfhaYXKPF+Eqd
jiek2gcRWugqTYeG9JLJkX4OVvdg9Axk5azbThemXd7gaDwLxeVv6YlxSzY9A8nMJEe8COuEpLRc
WH2bvEw7oA7yfzwzWPAr84ZRifiHYhsfBW5VhuKQvbD71rsPgr2fj+CE2svJkt4RAJIf4s4O7l9N
mmw5pP1+SdmHl4DLtKwfaS8VoT101JO6Jgo2praS+VanLMjzRFXaQGNrjYn3EqdipBcqugxlgCEJ
2TiFH6gePOYoadhiQ5p62WIT/UbpZtBkamCOkuz8CFa0WSq95WbjMQ7aDVtU4CiCPxJv6aqMLgtE
VhzxZKaSTsboNcvPFNIyhWRdtj40aPMcn7asxQDB9aGXZnXZ4wDyO+PWXU6In9F3fS4EVxVb6BAp
hkBrgEZTQcqWGBdVsjIf4Md6f0C8gZE+FbffsEa/9nDW5n0KQe6qy2nNhS75rfYyz+XVIw1XU0Be
kAytNRhJiv7HvdddIc4TWUzOcl0sfJFOu5Rty5lsgymRdi3lRQ6pxWzDedo0wPc6gNCZoWN/fhpv
gYK6HQbtzveT1qcdt734pu7kLdbrq21jWzV+cVa9eqyR2wLVVagEYNsuHpFQY0rtftF5HCuLCg/g
u8jTUvQ6BCL9P3shOPFCThaczZR81Fp/lJ4RPwi/FsClq2S44ghhSpE7J9qUFPvLl6ZRz/aamKNv
OD4m8ryOZD1MvQ5f3l5rGYcpSIoZHPPT2sFW/Fk/VU3TKlZLstuIEiNnwOdBrcMEXpHkDCM0QMjw
J2Z2ogETaawhx775qsoZiO5sJxoPYjOUFCmHqJvIpF5LOzrnhlEX4Qo6tN32H2If/FXEf0D5T0aZ
8d5cSOwDP8cJDJCn6NR18+/1Ghjvvc3ksx9FAPe7QFTn5tIWuvYWIsB/QEUN1kI2E5Kt7QKHbG5g
sF50D2A84/klAU/mOQ6nXcn/Oml/vHoL6cjHI8oohi3q3R/hRXqkp2x/ROHo7V/rYa6Ep+sY2Ucd
F10Jx0cCUjGvDnaoSwB4Zzucuqy0bdkgHQYRymYAqfX9DACFTlDLAmU4lMlOMuUaxMTNfYzDv96Z
dPMnLz6jv3DS4kp8wcVO0K19lAds93oQWIgJFGiZduy0hYYgxWS/Wo5+/Krao2U2Ec4/hSwJ+VrM
lk7rmU5yg+Q9XBXEpysXKIvkIDZ2MrMmPebp4t+oKKOutqRZ0OsBtJ/SpgJI/yrV/qdsL1xkaBF+
/fVxw3328hOEjCYMMVVEW2J/4FvUyEASWcOa1JmYS1nFT6hdpVVWVvZnOPW/9a476eT6+plvFcwM
kx09XmzRNHQ0Qqy7uSoA4X3qfWLisW89gdNKemBjfFDJgThUz5Pt9AP0YSsSiMvSkVqT5x0I0DU/
tz5mn8hIj7AdJlxXfUJHXMbS4sGYYNkBvBgXE9Rw4cCGOZmIe7boFaST60OFUuh1MEwtC1npC7Rq
mkexMFcgk5FXdnTDlpYTNNbM5TjWiAb25FK2vdRxTFEPoxgAATbIVFkH2lr+UiyTMgrFv1dVcSGA
y9bP8Oai+z0SrNki4xYDCO4GRgmeIVBXINh/0CD9B8ApW5oOsMZ1FAQmGbi5iYEnlPimH9BZDGgB
NAJH4fwmVMtmJCq5oCaDm3cdg4FzvMhpX4iYuZIsDRwj3vs/wjmgKw+/DqtkIctc6GkyPIwRS6pz
/gC6V4q1aTNkKZ9CSV+7jFRkzmDh8G4iJk1UhsUf3WX2NmEEtu5q6pHUN9teMH27jFazXAMaRvAT
UeEpuPE+yS1sqq/3ohYl4peym3KPdOBNQuXrImY7HSoi4m88SKFfB9ymgDHgPxwBybx1Khh1HTFs
3aBPRUVaLBcLg11CB0mW5NUMgZBGdb0FhvaRxtuVqFJL8CRbRtbMgpLj2kOes5ull3Pn3h5E2ODQ
I3g+IF9jOHIYcSfEi9xc5HN90jt3YnNv+UNN8+ZuMz5mPdDx5mJEz43AuF0GddnHpQwO1HdA4vcM
rksz1G6+55hN3lqUUUWtqbOhlmjgaZCdu03Gjb7vt5uDGWZQHXGzB4M0ikt1Yjf8/d8LVdti6a1e
VltOpOP0LYS+bXgiXq5PdYf3Zk2mm9COJTKdoHYeec1l/EngRvFUifAvhr4PClu4CuNQbOxNnpJH
KTgFKgpUKMKXCfpt0lc3dJdM+uB8lY6KhlfeSv3TZGvmJdaLRbgUxBsbZ8t1vbO2W7QrPPluEuPn
m9oTa2LSDvYDqvFbDxZTYrXazc77oGqdtnjHz5tspGTVp7m47pT9AqqFBmKzHVh86iQOdYKm/yX7
J4mUHV75bcVb7gAFMIhjtV89kTnWK6Aq64oE1+9hyb3nWA8Iyn2sVnf5LSZC+peFy3gWBfjzz7ML
VbGsYMGgQUWC30+J1nozU4alQiIGHfLNGOnwpuNp0Evxta43qLgUD0FgofW8O7lf7QHj/kAahm22
HvAEEnABQfytHNPYHj7xAOM5wbpz/5sJyTkEnewmkkbpGcj/6G/8lnCmVtmxovC8GA9kugMr7Qvj
8CLd1voDEL9YPK1De1cQ2sWopLYiN7zfnb4JurbRgyaOBT42CgraTtJ/aB4osHwVo++O53TRMnnY
CMO470H0Z/bMBJKGz9nJSo8Ihpr0pg+Luf8DkTArxtNOUW32/IzPIMrZLLqj4Vt+6GGKyFH/idNp
qC2t1f34HO9KpkS/Y2HYwRjUOvwwEIUOU4FFJeK4R9H/rqMzJu34v9djrmm88AgHUg95g5HKBXjp
sthEhywLTCQgw2Jk11u3I+zREEvyedOBPKL0qXaM6AV55NdxSe1Ytn7fNgvi7x/tRKHGgY04oquD
omnNxdjWlxFxjEDfvINr0EHPUykHNtiasZm896JLKGXspMSPDbqpaflmxFAvpAsyoUSNEcF1nyPB
lr5GZjY4/L7O4wk2ntHRk19aiZRrE8OzDSX3wHJUic67vIho22extONTmC4MJJHeUISMr+6W6/ug
uppU9iNBuhJlHNyx0x6wyisUYRinW9azjl3zQT3HJLA0Cr+npOk3QhHWY49PtrG+47SJyZcstxa+
MPmp8m8bz4hGDUfsS/r4BFhNQ9xB1JocfCyuf2NV5cE3sh+HOyk2yB/ymv4277ZSR+hustUZDfJ0
G5ZTCJ9bgDUwf+KNnxCZVVpEtdXcaoXRPjS3gj1kfzKhNmKpJWAYSPtXYNofGMdFKcQs32AI6iBH
MgO8l1IxfxDxW9MicWNTNjmOl2gu2ebMyIAjut31pkGu4FnfIHOaDMNbjL17OBCV5dlAYOFOlVQt
iQkeUX7ctB798+j6fKeSWpP8amL7S6To5NqM115F5rFJmiveZn8oydK2/wy0HqT35T31kb2Xo0fm
4rciXNNeeMvhFTmBzvHYi8kcDMkKYaWJj5XVhpRtY1lJPyON5lNgQXyyl3GBAL2TAyeGR56auOoq
g90oVtynhgxQsHrRkR7xdGl19P3QiffaZx0/A5+z/WIrZ04prLJDtus893cokxNjmm503L2aOVWO
jafDXrIxpmQkAUS39/j6bmGK4GH6IGlmQqmoyXqolAT1HWxNLtWyFbEWBhNSuO5uAmVmx4FWRz5s
+vptuQcwzdSUYx0mejDjzF79Er84zhVanpAMnBE0SdS0wk30FekGC/SRCCXX7N8O5Jqc7SFYoTl/
apa/tY70VVtBpupmkV++UEwGhYp7XgpMzABOdQLY+zPsoygBCmbw58wIq9X8LJS7l10WwUbNm0b8
vCzQk0UEsAycbPgynuh7Boe74f4GkusyoNdIc0TaHZqfw19srqyGXX3C1Wc0O9B9ufOB8NzZKxzA
PZmAJfsUegXUvxNf/I8TOOCFd3W/o2xRwoIXGllk/GK/JqkJp9Ha7L9GxpZEn7OaBfzvLe90kuhc
n31l+ALEEWxbTyMXpDtxjVs9TbWJYQG9nRuHjHaouvpHbtNmU1dsEQfhfYxV9txn7BxvYm6jJ+VE
OERm029RtdbhQLLBOFxKXRNO7eCHSQYsT/ruUjQff14650SOo7GvXEaWh4vld0pkE3NAuJU1Gdge
KfgHFmE2KvlSzFiisO8ov9bEOxCVItq8eT0aeNXEDOqQn7wLwakQ1Q75c15SalQv8vLI5SItw8fL
R+tOJOhvW/w0ek1lsF7csDRDWFzDXAl3eACB5uf8yTJ0nViTcK+Ob5cl8nHKDZdLuNgJbiMNVbaX
tVI2aAQBoXa4QBA0EQkQPVtv0fTK6RegOlR1vU07jlQRKYdtLcka8XJRRS4R+EBVO23xYt1Uag7t
sDk4iRI1yzi9zjfav4wuy3rW713fDxcpWrz5JpAfvPcSNVFGsG3a1V0O3XgD4ZKBON9pHmyQiMC4
LFtNSX+8HtvFcWVWZHPLX040C1Q+5wkfVkOaeaejdaBYZ0QxPG1BAatkqsUTVUUuacEh0npEM/Xr
czs/KrEekKe7BfIJc3va0OiAGe4PNjXoLUx1PJ339Bzj5Q2oF0HxGf66YPTIuvQoZkwNi8yg3d/O
y/PoG4A77o4C7n3glNMPr4BqUX7vt6zG6VXVMpTiGhZwqYra34DHIN8fVEDRdtmjyKP5SpTyRxmd
kFgOhYQ7B52AQJ+ZggEvoYPpD02TH15jNRLv2Amp805jrdePVU+JCwsXoJxOEfBBvxMkhGwRwp0R
8+ljdhMqJ4lH2SJqm6IjNKA7PkhXiBQAMRiJM4WZhXev3X+m0iLa3LJ7lPgHPItUly8NkPu7AdUg
kjSU119+X0iXoroG1PIiyKdhA+zAoa+BafZgcoVT7ahH7mzxMl1u/ZkwDEthVu28Kaq1v0Db/FI7
V4htzyos7etofjsiyFATzHk6dyhuoC1d2mUBYHcUaTWse7YZJwPN2zP6JYThfQsJlL3x7Ln34I4k
n2ARmVs3WrzrA1mDNjHCDpln7YiLxFvu+xzTmJdta7cGfCQ/GcxXKP/V001EGXSjkaHuWxFo5csM
q7v90dcbJmhY0NNhSJiqOZkpTVjXk0PkU+uiqr25wyMd5Ac7+2cgAkx1xtRhBIwG9m+Tfn39YGa6
XaTbKMeDaz0Hyy6haSp3xp9XYwvn26XUiGN45NGcq9a3EmsiNy8TTX3+g/zUcBJ/auUvLYBB48Z2
ZE47APKCcqaXeKBowj+tI44MCT6WJJECTCxpuo0rwSO6TYUWGbh2C2Svn6KSJrynvmKnL68I2wtq
pb5ebO/vFU3dG45KMtbvj5LGigRQ2PFofUtWqbFR32d8XQW145CSxhN8xKBdl80+uY6dnlfFOxja
HO0b+RTH0anustP8MlifNa12FBcxW6UgRL37B4r9NXuiBfPGg7ViK/0XFBzwU4ESlCjXS2DZfhiY
GR1IoS8dCbzldbkfZPKk6qMalqCs22rWO9q36A4WV5owcXrGiIIO5PWZyndTL8Ua1Wb3m691hwFA
htYPfBcB+c4ulrHF0VJYzQ+rpNMyMeEe1MKaqLod+8wJfZlxd6SbROEhAhp1fnqkt+m55WEqUvqg
dyrNoJHWVa26cvJ15qtDe0J8yS514xc/+HdF8koIvfECoodAKxQxd2fEOadkqd3fXYIlkPD2YLHW
hxXWaiwu3hcKv4TXY4GzBmO4Ihzt3mF8XAzjeACsdVuUxItc6OKzH+bVF3Wycnuv2Qc+d5XWUn6a
cQBUYderAWEmvRoQD/f1laX3/IejuOmEBhL66NZm8rciokB0f0IIY7Xhs7Wb3mKRJ6XXt8jI1V7C
MAygl8zXDQbReaX/Qe4iHWgz5OCg/Y8YOcIAWWCgfex7gNYqcwHTs0uoN29dVqot3Ujgw26/4HLb
tUYa9vsa9KF/y0ZapJDjOq/wX4NulDzeX15rSPzRbyNZFrYOmr9AzviJX+uOaMn4F5R4+wEDEXhK
ApMXHnNTY8werO1SJ6PkvqILUWI3Qp7pn4P5HExx3gNUupb8ycUzBu8BYWaD/T+dUCJqjwyuDK1y
FmaeUDjcam6CxB1M1GPh4JdK12U2+FUmPuJjni7pn1HM+b6sCxMsyP+13oeT4z7Zy6UZ3lcD4WmW
GHo00PbDv1Q2tvYjRAAdJvsmjHjoeZycd3khYeGl8qLVzkUrDzXwB/vvKE2/L+Nq/OgnByi1m8g0
1bfo5BxY7X2tojroms1iT2boqFBnc31+FLemd1DV2/jiywdDQYQAn97veMB/ACsNge/OqiqTF02/
HAyccLYOXR+C1lNhG6LCMP9el7DtZ3ld46QAk5MOjaTIxT+LCKOhg6EA1wVMuDaQCbIYkpIbmCCo
lOTo61QeJFkvhZWgU9yVtRdWdX8ErZIulmuLCdSQCQbu/TsPnwjRMgeaDehRASbNrqI04RzCTs5w
DfxP/XS6Uz8KZpLy+9+ydrNPvPYv7JrT5T1r8ws1R0KIuyBGqq9BVCHPd9FfB7pPGJJMJt7d6VQ0
x0Lh71x9Mk+qky/pdx5U9zeDBLQ+nqBKquYE2Rv0kYrEg7fHdUD92BEhNcEosYruUwUyc31/bx5j
jI2Q8Ei593nB2Q3gzVv6FOCKhqLhkq4R3HQaST1qd0AD7fsiqTpssfv6pVT4Z4fMJBmUPF3HYQ9d
mjUkyn6ZwNZDdn3qPNZkQAUJWICB7mmoOcblnqwRnV8qN7maYVX1dvafYQ0BpBMrUR/PAcMm6CCW
TprkQaEHfbft68qpMq2d1NJx8LrlvEXW/VSGrHbsZXUMnilTW/BFTuMVptA+qfYwfs9nvWIiS/+n
WPvpWJclPNhmKMiiMsLCpkWlokxFCEkJqRc2ElweBSPaYxZFuqAGnQAQvdnVNhOW4Ag4to0+d0sM
2g6+tXz6zJsYbh1/cqa4Y5IGjv5+8I+66dZwFmls/iz2TlhnT2PjAbhzBBLyTxwHzOxv2GiPKwdq
usvp9NwFAatjJzSFj2vl26DkTwUXFjrM1bii9i8UBZ8aai7hVEaS+jg/s4XDIjtA08FbC3gn80Is
5WG+YfE25+XJkTgGVazvip1DXWwZw0PLuUaADvck8H4uLMp8lItOMXAqH9nnKDzyMQXuIsdwsn5v
4hGaGYb0drEegxlC/iQdMuL8jLwOoPmA++aLIfIDYcCSw2JHAOub5eXwxKimq4tL7M/0zFiWR4Fd
7dTbYI5oEeZQIceG+lU8RkVcPtaF3ko1s06Fj4wkxK9W/rxwtXnK4RjppOjxS+9J4DNbYuHZWa0u
XLnKdQmkYXJZRDliz//5merFishbxhWtKrH816H4scQjjS6rhqSkuSKpwx/p2RXDWIQjceEfDWvT
iVo0N04wwdO0gZCHodmMTNqG1NCJE2QO/il3X/+P/r7HQK+MqaEtFAvDsG7+irZxImG1XVNUX0Aj
cmY56seSg3+91Oq6dQ1/0wIgFy5tiZSCk7p3QnhtTNlLaZeTCmgrvNCj+vVNL2YfKaEM7ENnvr2J
UqQ/IsiZzh5gat+FTRJrC+WGgBAJ7wpGskdf5ip/zUeCKvyvWzGGT/Abh+B0why3oFe0D3bFy6/5
NeISEt+gw2FetG2naN5eUNM95Jj+KA7eGqLVvuVmQM6EhUhcc2SyWNJqXLiX9wnk9/cXO4s/V01a
WxDudLSelrHwItoB7By1fFIaFtvrw7pF0TCpLd1xRMdM1HYlIoAR1k05V2IqE8AtpmaraQ5aUFh/
PvwRWfKDrHmkMTQyhgKAWl29LD01NzcW3IflR93NmKfHFLzzQe4PsFcNQjNYlncn5Rs4+lixWcP2
UZj7oFObA8Skw1mYjPFI6pqAH4Yfu2bK2SzJ7wIkxYPeCh3dzK9p7vkSbuVkfBnmN2bikI4qYVYy
NZNchuJQT0yDeW+DQphCjZWlBcex5NqMOfaP8whehlJ94MZLq+J9NYgWcHArhy2KeK/Qb7nH/5Lf
GJ5XL3yq5iZkdFNT4+FVEcxIXAK/dhgHyZVdj2Rot/QA2OAxKMZQhgiHsDACKmsTgtOU2CHg1u7g
WFC9OuV5KCwLP/yOqT+DvSGO2SVlCw9/Uf1q35mZCJrMfYuRmBkdFEzkIiKU6hEV1dTK5+6W+y5q
+7jykcpO77ePF2K90oeFb2dO472v1OhQilUhe00TIPIpgLRW4TSwwz4viBjAA3LDVkX6uUEzCvpm
9lhHsAW37hnpis1L6XqeY1kez68p3Ckt7JcDtX/tjBSpfkiv9ZA2J74gtnQSSDZE6P0gC/j8ykMB
415rc9WGvtBVLLkQDAGiVGBWYnt+q03U1VRvrYpTriVJkrUiHBBIYtAKJzIk9MmPwoYxes6iZJQQ
XbWFuccKOSSFdqBXr/f0e9LbdgoxfR/4r2OewXvPyUQbN5PS1lLJsSGCWcRo5iccu71E8YGtKv4x
sIG6Kvel7nAzSJAlSsMMM4vi74eaIhcj3s402wzoP9pRQdO3waxtBRarf7iTDV1XxKXY5bVn4rSl
HqSqI8rBSDz9Uorwdky16rG+/FPm4j1UWPhNdt1vNMjC7DVuz04emypwub/X8yuHC9eLOrta1f/m
Irg0qqJfA6V1KDRTeWjBAIpEVh0o6PqGUNbqarxxUPX49EduEsDPNoPay9Nn1sEdDq3eGRtNzgv7
bbtT+eUtScT1v9gI5PPz80RkV7MHaoAVSosSwXfDmE7uiBfRSEd2X7vDRY76he4v4mzhU7VJmkqE
0b7s+08Ymfk5ZQ5sf1zmOmgAXVRuA0NmIEKVLbsD2ynawL+xngjyCefQY8Uzlp/Oe5W0NG8f8Yce
E/xSg1RHBMd2KY490ul413rQ1MXOUta8XkcY1t+nFhIWVqBtp4G0UTdBO3GEVjrYV6Pjwvx4IiJI
MStBvKRSFQHX5GCpCuqb+3yAl/goGUoOBudb9I7Nw0AHZJqihL8MvMMAnE4FqH0Vmifee07eW/wa
/vqh400aqRYOk3/JzDVXmIcSL1sPvRVHWpPisXrYFXM33ei4NPVZa2TJC/Jkqh+NkjIgPfy03co4
p8Hl3OD9wSWQW4gYQIFIHvJkTetw8YQ01eQolnIrC/c3s7Fd3AbPkL7JsGTWxSLzhk4w8fRVl5EI
MHRl5BHbBplGa7FCaKKltHhIgDsSdtw4eL4HPPP1suq1HT39e/vMMMPiCdsV+eQzMeydp4xYwElY
QL75t33vnb9151wjdyOaKgXfUmRvNHcuuqdji/mcgrL992ry/aH69/JlqiIrpRvygyjAlBFsuVnK
sna3ilWOlaemqZpXxoJtMWv9oi47Xe3Q50c2jyXcPp3Zry95pavNeZvUKilVx1tMAxzQt8cRV0dt
/vLzzsJQgHSX2PhJ1g40uLXZvMMlBMJb677ptaa9hh1TcOg9F6lTRy+kL10h8jCbqLWQk7ZPZ1mS
AX3pxEBXRzlnEzkVL/HflnyUuv+4DFxtxqZKG3jktXs/+HBxYEwP7dWUSfA39eysFJG2pNo2pYdb
74idjwwIut0LFcD7+RN2GwQQfPVF2xMNoUIm5t4+4aVEU4hmXtbWp20VA9zKVPY26Y+H9E+hvmo5
PBmjdzkV75MxpnPyktDCrs/Ywr1HOA5CeHMrbXzUpCXahMJphFhcA7wxzLGtqM+6z1JrKMW0A5BS
hWxuZAGE4MtLWobPWk5ObdPLyDazpJOM42A6TbVkSy6mv2dDYemyhifPMvLtLQltXfcZ5xJENWig
YGm1dEiV/QHwujoWPEPrZj4LZ5pHcI7w0J1eCsJBpJQsy2JbZIgGD/dFje5EMHUIUc83mpDPtQtg
8VIkJx9FZVbJOXUS7cBWaCra7R27j+Cs4kmqUJWdhrjMJC+03lyE0f7WyMGSa2b6r040tD2+YM5c
AS1e0UqmUwfpAvr/v+Zq2b2RMYkroSK0Xioc88AZZPd7pFsAjm/YGI7JMjqHXYc+pB0Qxy+Ayrds
YjzlAQ0M3fu6lQT8ocK8m0x8DP1gVqAG7rtbaO1/7lmvvSwSVOc7VLqT/UYJZGcMHNU1lIw9bYcX
D9JVRkJiPup+gEtZpB/yuz+jIEbqX0XSuPinvGGVhvvtndSOQjfxyGkT+zqFq3A00BHrSfWAjmZq
BsomUElEegNy71tHWwc70Jqx9w3IpvIwDHE7/LQzYSaH1iUB2ejrFuLMg1meLtg9J0hruMJY2N9T
kRGCc/oPcmbj5GwJCD6YKjBMc/oZgu9DjZfqpNicgJhfFZrhOPFeB8vCRgB0Wdo7+9JwmuUPMojc
dUBom/PzpyUNld5Kx94V884XPYf7ST5JOS8FiU75WWBt5sCqGn9Pr8fxZ6Mp1DWv6aJbsuRRpwQH
DFlv6hetmbMgy8aRhEYEN3ZR3pxtzdaLsjpPXyGzKSv6pvfht9vD7kqk5FZZKoIl/D0J9tkl//eW
HSZN5OR0kIVjqpe8x3uwCJik2nsjoJhMrYd9sr52jct+0TxrIHhlT/6iQqYSLTKWHrs2t11VmdTD
SbHfhSIYZkMixqHJSdSDSHos2KiAT8fBV5fgoeZkzUIbEY2S8OBcTRdPkEHteHX2eq8ud7/o0EFt
m1cpz5xTkzHqagua0T8m4r8lOU2PNnV4S6q/YEsZGOnG4hrFV4+DTIL0GHLHH9OEvaQvduh6oKn9
I6v/uz0tDpws8mViS7Pzq2KCOofGxZTA8OErjf3u141eiON2jyWZlxCirCsGWTreIwjk9KBwZQKc
RkYtUCFuviMedvoSjxKdjnfDbCKHbeCilfJeOPy/HHCPQEOikrRYpHUzjNoYtNLBbUcLysjzwXwh
BfwrGwasEx8MITLJs6av1eB42H1kiQM5RnuMw0wf1y68OzmtEbwqu78puN5xwFtyGcrBglmiwG5/
dDLC+5Gh09++CrQGjVZiB1mlxe4NwVd946x3vH0VGA9SCt4+yHOg107lViCYFo+EY0rQnifLMdwt
EqTyX+33S5Um3KRasve8RAoQaBM7rlvRbuC1YQf1cYdHJ145jbrGjlmyi8YXONpasiRTutt6iBJl
OTxqEcNjtY6cnGB+CwKgh5jUuSeQs8H2g2SX98JJr6WhrrVHEeLpmNGUdnPA6Z2NMSV+rT/bE9Dc
cfMPbGyhmlubfvlf2XjuIle9UUuE6a8fT81wWIluXlu/wSWqEB0t87AqexRyBWceGkKECaB+4Pms
DIem8oMdkQGai7j2OlVzh8m7Mn7rHAYd229y0IWZDQPL3R6TNK8dgyHnqT56x6pH0E2xa9rheUgL
hA2y85jTyZLgiZoC5xv7qho4nAVKm/FkK8yLuywxe0JU3cOeRTnGiacKBMSyrtXqdNboF/MAtGM6
HOonTFy1Lsll+6E/61u4w3pAbN+9dq1zi56DiMgqJKuqsnR6iaOpe8UWO1CmqSgrJz7+MJh3fNZp
9mudt+16D3X2Oha8Xluut7G139jNt8wCouogv+U3uTAm8nMwOQxrZEL7RCyVg2IyFuGCEMnUCRxA
2rtNO+YdsJefB3DB7/SpnxwGl8QFLJgCjpVc4KiUAfvLiWdSIo/9YR5hkSy7KIoCtBEjKuQshpt+
HLOxckAOdf9W/RtiSx+MGJT94iuLUYviVQ1tWNaEVUTpXUa6uFswWAhu+AnMQ0+sPGQ2kkrOYPY5
IQAR+WXFXI2TaBawA34IVMWQFKaxcpgABlkmmEdILzIcpi5BfqprEqiwlhxgj3PpoObZjMMis4bc
PG0azfdolfkAdGPiAzwarMIK6BaiQI060+/S+FoRMiDFmaYt+mVhej3P2bsHVZOTd/IroeEKFWem
Jg93A3wzivk/QSAXPtWHfbfBe5qZ0r3FNq0mMbarstw3gmW/5vFzQTa79IlK6UMSDtiHRoDb+m+t
/WQfW1iyHh1nM3x6EPjwc9szAHwBItkEoYieQQVYEqbCMcsKJwxEEa8k8siUcBE9AHriDhxb3ucK
Yu5WAcZh8tiumi/QzxJoEB8BKnC0eQ4ppGp8lrCswnnkUcZotX5zOPLaG5PQwvSOacNlvSiMdVag
0QFzKmAKK8puiamx5svkRYHyOVLB6sveLGQjW+TpzNJSahUzfcQtxvmZoxuDy0ARGlspZSeXEaP1
+BNw42vMQiLF2mfzjdUXcYHqpMKCohUoerv008+zE9BWaXqjlkl3P27BwCa7qjGXTTkI8CZVf3cY
iVCR15d7islzdIPAHfowOfZFHPRNnRRdEsdjoNqpihokXuos0rVRoy7yzyctiB8oPcL8Na8JQ2xv
x6lraWK7NBqNs2s3LhwLtEdMr93Ksh8Yw4MOZCbSt8jnMOfIUVNF9UxRDO+LpFU92+FeJ3ULpFY1
jvtfPpaJzl0NefQff/E/PTz0D3X549kXliTwbsRIFmqcO9/3KhGDchJwpBQ60ci51V6YAN26B3i4
Pa4+FLB7YuVNpOH8IyIYhLTRbN7TjF2Y4PJdyuDAt/Zbn/5l6l8vjMUHPGpB0q//q0eXrUY57cA8
mc2xwA6yftgenBkDKtvaY+CRlUiu/iOoAEdnzlFxbgiBP8eXxSNyj0dnFy/E/WgPHcsplmCSMKfl
RlQBX4N8q/GCK4DLJMLz69eaJvhecoL/x+24jpEE0DjmM2JanAYVTWSxesitamA5WB2DwIL3RA6l
+TXK8V9+TMxTZ8BE9hkqp1lQAD96YqJswq7332bC0N129FSCgq7vK6+Hpclco8XDX49sTBUH141S
IVdPBY5Lh+UNoFgMNXR+bh0xyx2cg1bszHmPFfXJFoecFBCztZrhrr9TGHSVAXYS4buAwrEH1wk9
jMNnMJmLPFSNstOZEZsO2KdNZYe7w3aumh0/2RB0A5Oyg1Ief+TJyKIvy95NVJ5CIky0BDWvMeHg
w6m+NckJEkP/rr3+XUR3WQfHngVovHLJeeKRzUxWeFHCbh2/lCiPfNKMHupHrfe/KHEU4GQVhuLr
kEHjo5dVXd6OseZ5s/i8fss7y2B7nGmujNKwMgXnFc0+JJ8IWfjSgN2D40thct242G9ag5hqYyVU
UQx6FDlTk2QRuul3vqlaJjFjtDxROz4JWAdd+RRGWq5tjVdJMPQuHWa39sMtjaXUzfYn2oWWdc8p
ZDPiDAat8NgVNVtCU7mPx9ZLG1B5nDjiSIp/9eIH0+G5GWK19q/dfAtV9QhZWX7NbVWq3bxP0Stt
T9B7dBOxQfzM9gkzPaI07mj7AWm8e/fBBzC/CTd7KGT1hzsmqOAKZ7P8IoAAgkkWNbcGIZT8uiZK
bCjZ0t2PyUQsoyvjlv5AJNrUQq58AMM73JFkn/N/5YK1xelmi4ix955VouF3C/4UaNSOONPIZCcY
PmWXj00BmWld2Vm57K0FuTxn+X4tgpWpAlylp+D1DqoO/zLi9cRr3y1g4eNqztijrPRcw/UgeNlb
t/KvS9Gu56PjAu7b0uJI2+HrHbhYjBd9vR5m8wHQgGHOcxbCFs4EAYNnHQdgz96rayiJGZKPQYRr
lgAakjpHJIrP+VgH7OGp4dKHqfQIJwAr/sMzeIsDP4YwKcfgt2vYigj4mD4f4HHBdVlJixzDfT+J
3qrYM47d2VZ5Gvi5V3l8BWJdoV1huFZ9cUwZJmbnI+ekFSY+h8XWP2ilbnITOkYD9BVcM0MdiuAd
ZZMMD19ODhRe3j4G/xA6gR83mO7x8VpGA/0UeYa5pReqQL5FAVC0/6uL6QNXOuhqTOrABf1wdLWd
snVeCAnrh+XKkiorq8ZLkII4FFs0rkZbbGCgoFAqWhUN1xVxcIgn+d73EV7xru88CaN+zUMm7w8/
lwRSae6u6fE3cAP05hZnCHmaMW+sCTbtwl3W93yJCSwPykn4n8m/F1tTb+UsyY/ye+nnX97e1bcH
kPBXQGgcZ5P4UCl+bU7Dl4gZOx9uBNS+bydT1s/BVlxbV4QxCCXNKyC0ekKk2owBIWYFCapzMoZ8
3TJwcod0tSX/0h+CkHK7ALiEO804pLPHqvhkieleZtFHQognEqi/R//xX15pKyQrDPA7LmPcV89B
0QRZwwGOHPE1GKtvVaDeVbLhWvRH9T7YpCu/zRXtNggaL5h5JQ2O0HROmFnIcUGP4r3SDRvhzn28
DdfkrJ4etRUOVv4YkQRe6E2FBTJ67WsXC6G2adjYOULlaH3VVQ0DdqMcMTBUfGiSvHN9AbkH3Qnj
lKOa1sEYzIdU4s4rGHVg/9pxGgi3AZFF+7EgSX1TWGIYYdGEqbkkXqacqK+V4GBillDtneWJX5+f
LYPKGqLznroEkLj5Eg3tkXXFGByci+Pg0tOkzEdQ4BP5wppU77Oc3VvsvyXY3qZ4KWWpUlX3FdqJ
cN2aXxSivZ8Cn7rRwNWtTgZaKqETfJEXAXlwDzZA7q9E42VRSMwIa7jOzqC/L3xfN0olPzhnq0Xi
fde56hQIeuzHDuzabFG9epc0wak8nsUcoQ9mBVsX9gjEJh+oY1YP6Q9mCAqe6gSUkrrf48ej4Yv6
qhTKcT724eajfXdbjVd7o61vDfxUWM0PcPcf3vdYJNqVZXj7AbdV0MMtrz7YlJoQeljK1rAuBXwN
ORrHyTQqo5cOzRVzSUBWv8lRgUmMaCFRqgaaRpQJDVRS3RDX8PWLVsAmbcerLjw1pvpiAwMndPoC
sCyahyspeaA8HEnt2Vmcgr7dCb3wy8zgFY4lDA7Dh4SFo8dFg+Rpr7VKyH7Mo+ezmrWUijtDOCmJ
UQo8AOQupbjiOGLTJ/i5DwQt4qgDvlh+vDcllUs0WnSPepl5qZG5QO0Nzj/lkOS2bSc6vunIAnmM
moHH3kfgLqiNzz5u2OkOSS1+Wxjz1i7stuwl/R+cc6+H1TbnbJxqdP4wkTXgytTaavwx6/VcAuje
ZpqjYtJI3J36+Ywa3PJ5/fI956dCFbnBPZ5PgfwhyO9pakpEbNwWfcSePYsoTYz7d/EYTmTCQL4v
N5t/wGcgMa/Zj6EH8VCM7hDS5c0XaoFEqYZPGGGlLBbK+EDKnHegyXYUY8kSRCSQSj5KLa9CxUXf
ng5aK800aZd9eTULxY1VQvt6nVJEgxZ0Lt3V9LE/usPzggacPZcdr0r7yTAQQ9DbB4LLN2wQPtjK
9OVS/ShE/bVV0zwFiMd3D0rmsBh4oUb3RGi3M5+1DLAHxd43GwL9Y5JHAo3jVGTbL2dA2wTRNaqK
RpNK1MgpREwfqGZI2X5f9HtzVJr73JJjLbwcASnvjJk4adumfiYhDtKFEu0puYBtrcFtN8C50FCW
x+ONTVPGybkMmxW8RP42xBbneF+4VPgw0y0+ZzXqOq2dWZZBdhSvnrCVfCrjFZHPe7MwHMifjbrX
ZPyLxjwePiloUHbMRjBNpZ0vr39NtMbwVE++DfgSc1YadKs4H3J2UdUzfwJxA4JI+8UlLVn5aBJh
qmOgtzY+xu/pwOvYTP14d5egqXOXrwlP2Pf9z9IrZXKnjca+r7DSvApULDGhpgvnTZnTimyIGQA/
PVOfdhZnxlmmrTKOoYax3pZ6FDFd8LUDqZ2sVjn9WpK2fmLaJS3q1TruYO3nDZ3Ob5hhqmo/iax9
OXolpNaUMfJqml++f1bApv9NYq7ifXyYOXCEyihIN3PS91eAnIKe3MUn1UZuakge9QY98to0gnxU
vS5LmTFyhGT34+Cf4+AhvVoMCEDzM+vVMH7ZsCNW9DWvdq5OT4WQNwAFgVg1noJWb0YlJ5YNodwX
DkPxtUYGnBRA/oTI08Cto9/UAjjM+bkYB/lH9MD8KaUlmvKhtkoXfFpU6abC9agpv2r1Kykec8bI
We7wUbf4WYEAkFtG6YvsfmIgEIS8EvB1L3qG0EFfZag1xpaFA+EXnhSHVD113LJtzf2Yc8AlYDIm
j1danGBpVTMor/WKPb4SBfo5tm6bq+zJygYZ2fnj2VVnnhU2x2c/wckmwMSTujZCBX60UB8atQr/
BJMsTDfbtlFbAPqCn3NNXwuCdds9ZfpqYqgP3E7EmzH+axv3VVOFTOD8JnpIUWUQQQISoe5+5bht
F9KAVEhK5vslibgixGMULNhG1UII+wWy4KRE9H23GMdMudqE7KjFoPMGPhmVxoV/3fAEGD7KrjeY
QOCka2tI2gst//ykTpTubxgoGukClDLs9Rdydioym710raAuC2g858Q8CaZDwhRGDqOPwOEcRGT0
lEKfwRDKYuhri4c0ABe7S34taDqEDQvLC4uE04fwLsYNhTNNVZFydpjLWUgyEtyvxd6ndBlshuWW
THsSPUgwcLTIDw+LKonXZiL2VzA4At7WNgXnSKKNqvHj6iE6bxQ3noeFpOVzPupUWtBykEyfOAi0
he4DoMs0mfqXaElneT1qxLPh8+BgXopJ7HMnTX/IPYfbZwrz2V/ZX7fJuXeFyX2pNaEc9n1/PWg3
IIMyTjXxeRoyRXXLxMRGc+kYrhQr1ZoqYfWMBmIBIYum3DBTvrghKOxQt53mdStcYBFUoi/OXlwC
ttt0WU10R071u6W1YxZtQyGd7tFbldFK0tyrJ6Z4GaqLsOclEo2xYUbcahxQdCuaqUXcWdtq7N/3
446EkFEVNnX3Jvl4okhgXwrBWqVsY1/nsMOZ0MetnagHIKEIxdujEOkuhrNF+zwhHS2UfSCAZ7wI
ZUC3QdlVLRezp18oRZIJVIhWLl0sOUV3O8U2Dmrsk5NBCDWHSVdxcnReRtwa6y5ACdY9/V9cNRfR
yI2Ix+BO8JTTo5Du41rAtXxMlkWKJAcemT4lAH+C3NpXcRed8DXTC/90rUjNw8ZEbDTkT6+/DLQT
e0IrU/ewDJZGbt/PoJjVFWF41+IYlsPor9OVX//pRqdpfgieEsTZttP/YOUklEtddefoDn9DCNUD
Lu8hFjKIcuvSum7PAepbn65A873eLQxvx+6+gMuT0bE/Xy7NXwaC4o2g8P/3f2YHkFOuhBpzvakj
1/58srMB3l/KeIjwS/WaccgxYgLUo0stdSzPwMmKU6MX213n0fkXbHwjLWPuCgiSSZU6XQvKLewK
D1PkScMhqqcXAWzNGFTvOFItiHf5IaImyq5srXm39zlrAzgepmhJ/eArGy4m/wa+Yn4gZ+IyPLHm
m4dLd3LcjsLEmpIRveU/8ej4rZJUBkYskgmDcmr0N6thnXbeVUrSxc+lafbUb20qjkeLPfd3izmX
oyvv0zGl7udIplRqi9/xrPGRZkMBELp1ghWqPmKC3QQT5msgtkkkmGGxUdzRwIHLJmBxwyAjeqbD
04lcb7sk9AQIA/KQRMYqWNxktBLxMTNFthJzAy/dAPpRUBMeDS19/sDJm/Yc8fpo9GiLijuvtJyh
aqznvgCbe913klaWkKZa5aI9b5zE5cugr76FYEZNfHQ0S6zI/SsAdYu8+0HtYmRmgsdEG9TS/Oq+
HZfaW+7VF2Q6K5daT3VhmdMpBc2Gk2wif9KWdb2EfS2Yu6P2iYr9JdpC0IxGMMy6SLv0kbvzxXw1
wTuD7Tbfq/rbi9gKhYzSuKAYUhMniiqQAdluKWfPSXBxTmP6BNMhfdc/FupkML4Bf1hQqIKHHrA0
3wLI5BdXG1coJ2pK0KZDUFo4JJQ+T2t9KabIOI2thKhY/J7cE9z2QpYPmxw6KLLrWT5OdZY2LJh5
M0IIUIyUyN/GsHcICRnM+NhGRKF/G0zX/1M5Te8gxhDbAVSFsOMp9AJnC0VjNMF/Joh2u8+JmBeu
1/0td4ODng9jLdcj0fZ3I21DhwlTkmaOybSmcvwFtC3T/HboeC9867//hut+S0IsNaBlE/XtUtvj
+J0NDF87j71BgRf2o3EOv/THsNFiA/8iK5PHBq8ABW/NqHhIHFnVOq7rkJCNJi69mh0Zq3KERas9
A6QcmCAg9or1m1aqhq1bbqWsRsd9w2FEcAVFd/tAb0BCAn/JIhtFtf6aXEP312OkGuse1bPUIJQJ
3VrWVGD1lUrWDvQcvVQ48GEUcVW1OeIdvCU4xYvTOL3rogTgVRk2lcmcqKOB8vsUz9T+Boo1PMhW
jyDM60GU0biibxwjRy9hTNkq5vR2vNZb1smv+oMZfHll+irlZvGIS3eooa2zSoDHH5Z6V2qMuna1
qCoFxjhknjwHGZD/NZybhK+dUISYbxOR0HzviOx7bnMsZkvm0stlS79mhQmJzQ2MJmaI0AMqDIAA
xSKGQUXaiCU5/+Ay2rdQQMueKei6iv3FKqZ1JiRmmHZhle0n2f+WZ3LjY44JM/+kbg/Y23MxNOUK
l87eArZfkwtMAkYL/Y0KmU+dtdsidZIE8JxJK3jzICmlWOkzBG/1pAt9C30+1CTHKl7Of5WKqMet
CobQy6tAvyqsFJbePdTEhoEazaLXVni0fDBYFNpvnnVeOjWagvL19aL8+yQgyeZMNFZ2/oO3L+MQ
yPGLRUovfx0a7l56UCxPLVY7mX1yo6PeFnZ1NUAvvQVn7QmJUHIKnA+gbB1w+pBfi3qq/TzH8zP2
UQRp5b52uwKWyS5LxnaRLPyRGZiu4FG/thJzoa/vDxPBfSP1IDMROZVfG3U6eUQF4cOFKKz/igOh
BL3BZqqI4fiXTXpcPb0C/RbBXFiQJQsMypvDL7GFezttddZzK4yh1uxsscNQXxICZP77/5LBsjlI
2zbY5Whz8yA1FaI+DiEAz+b/Td8RbvlB8f/yoVkZ0KQn9GKoUjb/TexjVaGowhUIVuCAwPtKiGUL
FamQ8nqEGw6038Y/Bq17EyNo0FpvrZwqNbn2gJ2fDJUqOX8kpQpSLoU4ubaSpRd5ol947FBzS3j6
3j8D7DI566Li5xWZ4fnyHFrVoOOboLKv4DVqzGB43L3VkpS+l34K3qCyxgfR4KlWKu4/Xw6pigiH
f7Cy5CYTkZ4u+kGA4EOc+8x5x5eXnXdRFNkNd0cGu8Xv/uI1skmi5IIiYWgp2KyCRsGgn/LI5kY/
uGzw121pNYpqSmqbu13tihnhAxTOqFWMn3LgOzp/MUzm/P3VHqxwHtZaLyiDF1mc3LrwP8jFuHDm
3huXWW730jADoG512n2IB7Rzzhys5R5mKLIMyZTwJABMqUO91LQNyEUGMJiagiF/6NhI5OAaB/VM
3lZvjr8WKI0Ew36ahodVdwmxnDFCCQxFfgehq2mrXACzs/XdHSs1kbg1Qi4jf7iN66H9oOCaEBZY
UHyc/6AK0+DhgLI8rURhTTwUd6eHZ2TV3OYKdFwdVglQP2wzvKl7jCWQggiBVxZnjv9t4JIm5A36
Ir+tQCwwLiWF/FcJIqVKVcOzczRhUQTL0jyvlEYMgswN9TaQcF2BKA147dmoZUuaQb2HGECE+H/h
k7r+bytlfHrEH+IuATrb9XFzDQiiC8LPWSFy4Li16SeOE2JeHRZfUxLiZSrnUTx/Q0xgy5jzZFbv
oNS2zk5/NfzpK4e3Wl6fFyd/PVxQlpXJA7BT3l3iKDcFE7DmLMc6F2k3S4+rkMYm6hbGvRpx3PYI
i2ZDA+AjnsE9aO1F3sgQ1WxQV5c1OZJ2pZjinfuiyropeylvmgb9CZiFIGIzt+podJbainLV9kiL
FazyTrFNT6NyDx2MFiaUWA5lulrIQTqJmDlyzSmoLpOEGgn24NjMASwJAIWZp617WaxfkHDpt+BO
9dZ1hKzqgAktcgMqh3L+cLKCO2Xjvf6I7cUhYB0bEHfT36mpdnFo7XUj25bQh2VMyFMyJ9jPLGFO
BAtuh3TH3zJPbDpzDRHlTmS3Dbee72oY0VP7Z/iUqoPIYoJNc5q6kSR+7Vvhs0zF2uyuxft+cIuI
i8ApPPNbYZ9ysZdzQsA8d10xO5wFbQdWqHd4qbJAOwi9JIukYIxc6dbc9+/96/mzkNbw5oGuGRTk
81MWW8xyI9trjCxJP9ojeBaf7fALuOcX0l+qILTT83tDFbhKab7HKx98pUN20osunMxQ+DRPuCvV
RqqYXPsCQU0txCKOV0tojzchX6U02JjZITI0wiHi4zVWQNNYLikN7KTZwPPZRQrqHFVCvLLBEoX3
E0Cw0B7bMH2hQzGjXOhL7pg7OwOc15HJso1+p2+WOMSsscQagJWhlgPK9gL2tXZcM70AQX2moDte
OW+lTJRcdkWdcaMDdHKwpYZVWCo378paNSTnB+kiRhJC/S1zloJnWSmFqklSWSXQ/+URhGH5fIxT
2riDCiUhkczwdXhSmX/Y3MMcnYqE6ZM/x8qOTfLPwcZjC93OrIiSKimWE4UMj9+UzD1/0Uar76gH
1Nmprlu8PA18IJd4Np1kDK7YVxctLgzULhCYSqJ0IyujGKKLH1vZXhJsucTtG0az129O+9TOCWSc
n5rpQ28Ld3+A5GK75bRi6RLokBbyi2PbqCsErvtdYKznoJsP09Mp+sHF03kVK4LNpRh5RUGc94Ds
3cO0DOnBBAljMFRSpCqNSJPMhIHmDU82Dque+bX9Fqhlw9ANh68qFLMK9oXrSm3apYvHLjAKQJGi
xDa76utVf7hXYE+Yw5Bylrlx7Unqnpx3Gol0sBaEEdYJo3OJ4XzqfuNcc6ZeAnHjF99BBw+JWKGT
KJweTT+iGueKDwrfGOwHbD9aruQiwba1ev1PH5IYIJwnfCqDsFwZ3wL6QKHZcAFvbmSkK2vCh5Oc
kormk+lNXeQgZD/ClR6IVtnSmqv8y5SZTTi6SQIjAy4jDb31uuXhaRTG7vx44hq0A2m+1uZKiaRH
uJOSFh0rQ9zPCySIWrXzWtMwv1717KTEhO+WzEvfnnQm0t/8w9usTu9rK2Krjq9sBxmucxACxMmJ
TMXYE5AWaUyL0JG1a43GtdtD0ZoF6ES8wIN6qQVSlGuqRhyqdEiFp+E9uv6ow6sWDcdNALdP/sH6
oywsmb2Gof6jTKIAZIDy4Ya7N0lundfy+8otgIXrozz3IoTccErivnE6IoIYURdDTWY9psqx9oHH
tiUskv9SBEQJK7jy9SSyepBdvX0TtO0Bg3vKYKZ1oOtPfPJYoRZsWxrAobln14L0GaXyyOozkn+P
Vn+0XTopi5nQYQvYRg1Lbk4DNxtPuxMC/XmMDgU9ARcp+q49y3RC+cVGTP4jwUyLIO+5VOZ0isPC
ecIitCoqre+4Kx3rddycxBctSZapZJopo18FOrlQjUnczKbwlw5bGcq9e9b9okqOxGUHi412r3/v
43/LdgC4XnZMWkvA79UinBtGn9Qns74yhd9a1gMUufB0E4PooyZQCkAAXdBl0AeLfOcL0iZ9wYnk
S8CH2IUeVAuk1ePxGwjJ4CJxAvtOuPmN1UL3hhaESUuz8ROv2Aekc64q7E7l22VXyrzwF6JDvOvj
cy1kWZ+cdKbguAmNnYjxRddeCvJqDBCPlHoTTwOluEOIB/NzH25u6jE0qp8wp2n/4apYEdgrCZnm
7+txU6fYWWH3DdYNxzXRCA1G5yzqN/xHO+GQELAJwTiFyaQaAwpvuVEY2OGwW3B374gxGoMQ/Tx2
RkfbJ20Z9K8ofs1EgfxfF0DVg74oUT/o3vyQixY3/+p66ApgBwswkDTC21D4o8WDbfl4fVSaFOg2
s9VIEiSDTOxtFwFiNnkPrJBD/uy2Vlt55NgOxgnzOBLzs+RicWoLyIZpCbFAIktPYmfO1KfHcDtl
HG6AWHEFjohoZUNiQoJnrMZ7/XCzMWI2epQ2bIPEJGADiL3Sabid+2j0YF0WsLQLtt3aS4AM5Seu
0HAExBwI3k1/KwtLAFKWttf0LH7SPiw/AeR2OHCuVTfJi4Bng1bDsvb/q3xf0JzBKbq2ZBJ46IMZ
/jDRmQIEKBLEV2do9CumooDXKseduVtCwDidvEhqXLwb95L3hm9SwWmqFszHOCAhuvcOrH/dlxjW
2z3DYsbsD8yWnwQICrhbGz5AvgZAJqskylCzs9aOnoCKFtUifP/5+gWM05K6uUiFYJF+5qIEg+ed
nyP4kqw1hOs2EUTSbKK4/BcVtbiMgng5J/lSIwNKOyGhZ5zo5cXYqAbfM/sL+WZhXik46L5y2JcQ
UjxGeesaCu+o6iRZBR2jq4PCHcZYXDNjVv4qVx+sE9OmkC09QEM3eiHHetrHNY7S+XX+pyFXwqvi
4wZNen15wSKVAMvHL/9K8QIiB8twJsaAfOkEuln5TslVBboh2OWEQYuFnSDzCbTHhOglk92wdVYk
JTeE5XwjbrOHn7Vm5SZRvjG14YWKYSwVJECVUjCYfE+0NinMSBrebDp43UhstXGYllCCg2Epl19H
stehiIkqJCszYJXiALl+VzOje9X14FkiNteVxRiyUFfG/6/4XZnFCfP1dsleFleCuM55mr0cKdb/
7wuWW0Jhm4EzWFT//rFYyItC1DxOai0cRoFYIPfImp4Qdch5x8Bg7x4OqnrZNDYFQa9Q3uxEEDfU
NScLJcutAQiDqU6TbMPTFJZNBO1+QClPXaMhRp2m/lg3NqVNIwydvJdldMPZHrUt1ga5iouhG/1w
b58beCRQKjUDeLISLuK90nZW4Cuj8HZO1r4Tpel+gPpETISvjFo2PxUsKUP6kZDmMTLValE7UpTl
FpBbpM1AZsfG+D/ckuoKgFxK7ClhXShE7I7ZNaO5c9geZT3k/hLuiOqyWAoJHEY00ANRQUgh+uEP
nMVK7LTZjLeBinsrQtMSABRi+x+tXDFw+cly+YD6GFTGF3aUFCf4oQhmGyWHz9ldNmAJnjzachk/
4/fDehTdDBTXdQDMtzDKjM3l5bggZ6q2QQDPO1SbByWVlU96y5a4x8bZbpaMFNKuMJyTQ1viAx6X
PhBhBwByhsF+hG7uAYmHiD+KhjLfDbkGWeSKBZ/5TXQkVtoIZ/wQbfwEzdvh6JtZ9TYD5ENx65Fm
lZ2sZn0k7DDLHIShDq354mgojVmM5tysFHbUIm2lx8OUNNWZxSkMQhOnFCSV84tVJzDIcr6CxBOo
YYJhnBcTeDYGLPkQrSiYvUYmIGZ+5TznU+BSZgDg3ydXByC3nYoSIrAP4CFTSHy0HJhGbjhFAovU
FS50/bWPL1XA5fzTKQ44bCuYFbaPOdIJcR0c9CB1roAg3lU0Bfjpx4cHIRecaDjWSXi1ezMtLJ2u
mSqPe/6ht0MXaa9KGBlYbx+wjK2CAxg+Mv4ZR9h+/Vbq32YWa+YEiAxea59Hf1FqkCFVfb8W30zf
IdUx9p+0L1aR+DRW1qVbzjWnvzcftejIr3Lfc7frAD9ydYv/ZP98NoMg+ZOOdPyuEdtMpNX3LOsg
Uo6FCTeHLWdEyJCoDMlIwQhvJd/eUOGaLMHn+J/NGVbKlE2V+4PoijNwbmJ/GB0yjrsT2VmFQjFg
a73YVuIUx+DSTdhukGGfdoeYTX+LUfVEAVOR5N92cI+LUICtYUDEIYZylcSF5RHXPVGPhyfgZ39G
xDXp1QN8gqNVFkNMUmuleyblnw1zItccRxWGW+kc3F5DZNiOaX8sRMP2AwsbUgC5wAMXXjBbvP4f
MxCAAPY1LhPN0w+4mK9EpC7AUdIoB6WqAkMAkEIrLLjvcOuEuo52maPIvUbnYxARjqaC5DvcfBS5
7rwwx9p6w0kcut98du06EsxfFKCg09FVYaN3gPAb8hWjIhErwK+G8qw/DdLFfCPrbFXGbIw77WM3
tlP4L2OjjpomMFm7ToImlPVV3XoXVk6kZauf8+TPlcX91Y4I3Le0R7XHrhr94bGtov3dH5HTgho+
MmNqm4x+qcwN2rtpnoudCRGp9pBv8ofTQ7E5/vAS1d7ea98XFioIx3ULPmS1/tLw8zTNGXQ3fue4
EJy3ujFNlQbp+xZc4OoR9pbKLzTQaLGJzahm+K3tU0owDJIaqeK7Z6Ga7EW8lFf+5Z+r5+Lvc1B8
Sfz5m63O3Kyt+BXcaXdEGVSCbHO7xcQEhaI2BouOvyrgI22APPXr7GId/Mv5BZXJfPIzX1IALLYD
8WNIzUXu3Q51MDCOpJIyGoitPbKUprpvHWsSkveNIwbP+hrIJ0IuFGc5xEBPGvgWPKaYZkHFUP5d
QHzrurKneiSJsj2ZXtv32oZOSndlt5LpYik96lAU2AjHQNqXkT3H/Jsoskaoe7ZEmwipx7yvRKdz
vGqsu9Bpbpd5d16SAS1FiEH1Jv12ryv4IdKpPHHoSkx+LUT4xg3q00yhN2NNtMKsF4ObHvhe251U
9eGW71PeVRBcvXj54eWcYavbcwUhZBXrs5FCwXfa4v56SZ8pK33RFiFbDnIBJnm1E9q/ijS8cth3
MSzTW6WOBCf3LlM0fmnllJB+CKLi4lxArSIBvys5dDsu/ovavFnfNltJ8hqxoR7uSotvhurmo+Nv
qC4rnlox44hIvx4PWb3bdIFRUFkVKflxcTuYrDI59DBLZer6BdevRUQeB1mIJxU2I87JRpwZq/7z
799/gtrKzXR0C+v16nPnoBqgPZyBBHs5jliDUWmFGJM8AGSgstTsK1wDkUrqf1ns/oozwDXP7Qxg
IOtrbrWr2wduVgHN7/brpMp+wssvDxXITt2GA7ymHWM/fBkki70QzzOeiHO8G8SxKu5ngxFqO/m+
R92seQPHWjRfpAM3VkHU5M2QBcG6CXm0sGw4ClrQkd/pY/xaI5GHeQNn5uMO8eX9zkJH4WnL5bJO
gMQrpF1snBP7DEnbuGBciSuYw3THQLbaGxeSFptHNXfZaHKSPGeLDUz5K6Bk9y3Aqv0YzRHv1MQw
0Hs/dkj+EGsAauT0wpVW91h1sCMemieA80vwhV95X/6CS7gDJadpqyq7d2gBmwJiyBmp4Xs5EOy6
9wmfOe+/A1F+Nw7vB847A1i5EgD5yxXPROGCvthdgojA8xHiPcNTYtAUH0kp4u2RDZGhErQdUPhO
On/zhsdbj6lEkr3+OJhxjOydBiwGOvtcZ0Evir4WhW9W+uY+05LRXF0qR/Diu8pkeUrTpkXJBvSN
aR0PhkYwMYchht0N1gmcWjmw34aWx/fiue24G+3hEEdKty2noK2tnryIGbQq98v2Mm7i+9HFEl5y
GKl/U3wcJTdGXv/fKG4zE9RS/vO+DQkJUvPaRdu/M2yhPVaJ2uwdkqB1C/quKyRJEvOqgC98zdBV
6K7dn+fHzsC5uQz62NvsHU6c0PKqJKB6/gqUd9d3SN42/bQQkQ4amgCriIMt9nV5P5yVwbENhNx6
G7C92CdMrR2PKDx5wltBvjzmKSWejTXDokG/+k9iQCkYR/zpxFBKgdNFNnbN2rvf+k9HDSUBpQKj
x8JOBO2cT18iaOuKgvQg3JDaMZ6ryFO198Bsp0Fqt/ya5UXF3siE1e6lqFMNOv/l26VcM03/W7iF
i8Hwe1sRgfqpt7LmSJ+i5UDkbM1Hafxp+3Tcyr7HyLVimy3T/M77AMJxJBtYjx37YLOrjXMhf6iw
CFF3suNZu3b0fNI3pAkZh7RI93YPr47aNe1L3zFzHtCGCdaOd+CinLzOvgqRTw8c6ewBzYHRWMns
tQ0OV2DWXYtdWYEtvN3uHAErR0wTkc3vfRNlf+bMdO69kdQmC4r2OUHZpEf1HuBis6pZaf+hp9hM
/vpnHJU6uGVtY4IDM4yZrAP1Q69fRXNB3QWXl5/42xw4AsGIXi1A0efxvSLfNHtw1aKtItrXe1q1
meCiVtR/LkRIPxpqVo/IvxToOooDcdz6gMV2YsEz3w0PmA9LWQiM5jVWdFxfDK8rekQzL5mnfD9y
gtOvJYInRIdXbEJQ0LUZ6uNSzn1WA5Cx8sPVj4aFG/Bq4nHaHO2G4AvZJWqkyJfrPB+tcjvWezHk
zPjVILmZeY5lAH74e6GLunNKg5nUeSmNKHPgsOksiio4hG0OeLt8iscXmh7SwKxEmyZI+d9CmJsG
UsJQprJgsOTMcycTw1c7LWnMHyE9H0LKPeHjXFAyJai2tjTj8xyomUbPAtKY3eyzcIJDTkHwVmOy
R3fP3L0/tu0HRYknIBfPLOEYlOqlaidkp4uSXx+uNv0zl1A4HekLUccdu1Sqxp6DV0UkX9bKfE+v
b7tIp2bEcy7Y3gyZxggDDZlcxXIYmelKv7Ko69tt2gHSH89LfQwzzgXHVin0WMbcwWdHUHR672Tj
MZDqraFEUqlDijmj6fJKurorAQD5M3sn1hGM9rpuomE35Vi61AvMBjb4dbQIPsTHlxtIfrd2ss2+
j67odr+GVe5+PKwyCeAbbshOFIpKN+Q3Mpjxdxg9s2InTIKfBjG5KilQNyCaYFxvx6Z7jvBimICy
vUmMd9zZgkxntetZ4CcN43xLXCVnay7kRw7IoF/ac0R/iepDLXVpdm7M6XsZmlC+Q6PIFsutORp6
2xcDBd5mi242mt5BWU+f9obf8kxS9aUdSbG0Elec6NfX9MZxllZyhMJ58WgTRS4SCeshjIL/zN3R
JPyQ5MBtbo7RVim2U+WaA9lrIDhBz9CYO2wKYKos46dZGrEIDXXZJ6Tt0Evx3/N/+vDb/kn5Luwh
HExRopXyYjgrPApyB/RTfyT2dnE74JPaMSVDqULeUQsugTkJ/Pnco04LREDq2o6cWndLrSDl4ms2
8wL0KbyiaAyM9cQ0tBoaaPFmA7I9e0nLB9ZgVn3EE6bFp2SCye9xUl56XHlkhvGM2oKkK56tBhj1
ikMIDB0FYX0bC/VjzJOe03MmP3UM40RPh238UETYKHPVvqEx4Z9yf/E8ZKYy+KxzgHoSCnZy1SO7
oT1RejExFUJEK++zPkC7cR41VP/4IhczEAYhgFdEcexscN0GUzIuxzWglZ/dYn0W+CQrUMbflHDA
rMTSnvv3932y12ap/RibFiZOw/n12OWw/0kbYO72LSGXv7BvfDbE8qvctb+ZogCfEQG7kq+vYzWf
ODzSWWrwFVnJaoE8LPqgb7iW5FvMSAGAb6tQkHu/GAjZuvzFk3VK5WDz5beiZe8mslnx1hJP6UWS
sh/c4OoWJGQn0SvgIxe3eIP8JhUgrzP1jOutJN1GbQCZ7LMjWiZn84NL26r7KkdZDTTgZ2K9X/s9
ZGdWZUgMN2POVPAeBZSaQVewOpk11n/snIA8OVZqX/iVMOiHYroU7A5L+n4AHnLKYPqIdQ1bprlf
rVz6HRto1Pbq4IfOQ9t/LkTDaxw3YKvsB3BoKVNIirgaGBeUgCULDXkEivFinOwyHWSvaVM7kY5G
E+Cwqtejs4QxRYCqryt0gBod9A5LrIuT8Yt5cUDyRjyjhjNpmMop35iKkaM/Pz9jIij20tvdznXs
Wdu4cI3yXp84eLypFSeUbvTLSSfhnul5JuFl8KH5vDdQJQoIZLkwFPqoeXM6A2HOarZf7urgnsCK
I1wjkG/Vt34E/HF/P+TzHs/89Lg3t3ktFcR27eurC6OZfODxKz8RlDpmZK0tvwavEgiPxidDPmle
rMXnJSkSIMf2Fm7obVLBAwifHQcNw2oYsvHtYjslw0SzlTMaQMuFVx3r0OYNNrw/xHqIlN1ai9s5
Kg+zz6Z43IuL++WwbHz5DWavswYgmVZK7ZgRMzW7wOTNNoGnjlY1u4FGKhZbpaqUyw/mlcqUYbtM
LSzioUyC/RHM6ZJCzWRUNMc+loXysyN0BJawTkf3rDH87Yu+gYFzi5fELgauVp50grnyLzeo/RjN
/WoOHCI19lHAt6JPMi/YOJL2UY1ZqMTpbLJQs8NIguChw2Vy1Ih6Uazdr9VMaN8xYI8++9zBAfjt
55coB8OLX7hlxGvd1QVdK8Y/G9VoQ7FMl/1n4iyswY0k6j7ttm2ihD7/ZMwDg/z28JaCN8ffdr5P
2i/7YKSOmDdgLrsAHdwgZFqVDOt+hH+01APL2qlpMfncIyjw/IQc/vs42ddzt3zFK0O3KJyXfEgF
XIVxH2xVr/Pn/gmg5y1WCH2klJrdMy3sexOhkXlrpMhpPw0h+Lk/GYArKJSzap12UqmnOKW48bcd
DrfmceDr8NlX3uIcyAG5gN+/fOcXdFZVYDXy4m+IaIRCM8/YMke0qT/t8ThX+ORr7HJbwOReQlPy
rAzcfGpw4gGYdWKdqMAaKi4SX+EKC34AOBXFv/xTTA2MMldDPX8R0ereCixd71O/VwaJ0HZutCoR
DrDwUx6xPRlm23jfRUKApQx4AsupxT5RVnBv290GV0FpSXQ3n/BnUAyXQnNnBarC+T6su4RwrDci
9DTlZr+fl/Gt/9GAE5buf1A8PSIrRWavFJVOvTRwv6deJj7oT3JD+jX+4mxMoGSK33Rg3dX32Kg4
V5v4fE2ljR19w3JSdgbU2L45qcH1CB6n/6K6rHnnsyE0yvYdLeUrYRURl9kgq3f1vSyPcFTsovBM
uMT2YGQNXVkEpHCyimOzYkX09n26oHF2keB/AcJmynbw5GNXKxOCOUuYD79FA+EVI3iXJ1u7ZUUL
zYbxeygYJZPgzASa5VptRZQhpm+9DLFs0IBp8jyWCaXe+b5biCmjYDX3pNnDuSjwWNuluokbGKaN
baANeQTjRnabpQ7XuFbzf2tBqMX4JIc9ENVEpRhNS683n0CWGt6Fv/ZprE7gqze5XiT7sVHqEwX7
roqT6Nxd/ev3rREY1bURDIhFNJO3lm3VQ/QRcDW34WQxEIP2dQca9NscbJW/tQw8+avU9qiu5dcG
AzURtPqn0X3VeYpvxbKukxnnho7BlsHoOirGvynU3n02Ptl5tuI0RwmiXnyYhLJ8pmPMP8ea1SHQ
saz9NszVbL41gU4uroEFn1TVo1AGWn0bn2cF6F+dsZJ6O8yItoNMnlISqCVbrAThHnApMgdg5jKr
GSrYfeklub39v6TQ6FKaVSorGz24LFm3/EkY3lXWD52OeYrCDiye+Z5RW3+hpB7cV27RQQrTHrZd
ClJ8UFeNHmDbp0NvgtQoiy1Na54InxXYzbOnQBPn/JKIDGTXfaIuNP6MS+GJNB2tsQUcN8/3GcAO
glr6ZHgPPvktRqZ5iQGfH+IDjFOKe886Q0K9hTUtkl0A33laX7rE6YeSnqbnDDm1CX7oq1IiphRI
JBRLayvJXWcKhtAbio9tqz5Mno0XzdHm+dFzhwnqX9bKhreEWmy5VKM4feBAl2UvZ27GNYmDLFWq
61HmO04RRSBn8Jxows1BX3Jbyqfd931LaYN6TdeCigw4FtssxHmon0CMRIdgKpQD8dhciOvHwsMX
g58eVIXZYQyYqNRsRv9kj+f5EiqoXeI0chY49/ZDmUkKYTR4IplrvyOEScoqB+PYrCrG/oNasMWZ
dFGR7Zmv3jhMfsOY4JMw+KmJ73oxhMQyK717xrFQNcJ4VkiaFkWFrBCwrLl3ZO4uuVyUGMdlw8eS
7y+ZlVySt05Tc74G8T1nAk2aIgazuMSFD78AVDE52n/FVsx+xgqpExnuLY5Lic/nsQPaWm5jP21D
iI18XwcCsl2XsUDfsG+iaTEfHuS33KWNVyeZlk31u8RMXSfUiJUW0D7pVUzSWPbnrIlOir6YtF71
FmYzJD8ccvZ/MwNAMCBcX05ep4b6WkKPnK0wDlbPe/n01oHegV1rjrJfo1ogC+DV3FOspu8VXrLB
VQceKmPPxdS4Q+ikQam+ZAbfZ9cUk77r/UFMFaKvGTvW8o4DrCBmCo/9GuaiZXhIseCERulP+3lf
QxDyU7fE0k4IzH762CdGwdj9UOOaazqrrI9Tk1LLqe2LK/2pE4OdbZaMzHF1u3H1ELKyfKPyGVRY
uIgOI3JONQQNYspgu9/NI/7yRF0DTE67DUPUgNVwxTF8I/K92pPu0XWFmpHU9hbyQfeyFpgik+c7
WU4/ygwWU4NopTIP88Fo1TQLK4k7W/yDbGtIps38gDxX3+deIzE8nBtEYnf910B0Bejz8YWa/u/O
0J5MrY/cutK0lsL/WO1gcO+lNxrV7dt+uYapP6iEgGK3YEfdnn0DA/6SOyIOInMnh8cSN4/86qTk
+DDJyepPdHUJefFvnuX22fky3jZABY7HHfD8oDTOS5Ig7BlUAt1KBG7paAQJs1ntMGfNnTD4bqC4
lsgMHMq3lEoQ31VbiVWpnvNB5vlvInjcRCDv3bQ+x4tSIiGLqJqpUBsIF0ni0LsjZ+yj4ArOtrkR
eKUibsB6zSfa3F1XIuxeg0qH0l4C7f/6PCe35468QJYNVqHt1YaWdT7QijIw2sp1o9rrrjbXL6pz
iOZIpV8BNtgdKm7PTI6Rnw9wtpGushVgCuo8JoFEEXNqr2Vkey2+K+CUb7dY3jlB6GE3jtZlspD3
kYu6BUISNQ9Yge0AZ3biuItKG3RP4ZVvH1BcI1NUEtTl7ocKsrD7UtQ/RifZ0ImGx+XxOulqvvM9
zV/JuUxV0IXNGu4S1Pjv0pM+XeWQ+yp+kYkTptPQWlwT22i7lGmXNfew4PzrhAudN1f3mSFlMr5e
2I2MqsUsBoIeCQ3x/G0nZU9qLVHs22uBmdWNtl1YWEoTvbKLlQDcamBtm1mbvKKJQ7YRZ+bz1pE0
fLVR1WbKrGC1RI49+7DagIB4alLB2qGycNX9+RKF86iY5o2NwW/pYni4EvW+EDqUbTB7x/U89K+i
tJ4ShdceRGNNm4aTWw4GraBtGmk+7Qj6H9UV8fiC9p8NUfHFjY4lFOezrU0Sj+a9/777pjldNFF3
Woa5Du7YHRyZJZjZnMgmxmFDty2T1WNrdOQyppzaftR9r44kfIDu4HIefNXGulPtD0RdZpx1TDbQ
+R/NDW/gTqWjn+WFslG0ogXwUvWre4mhYcS1sv4rXHH0EHTCT8v5EPOSexzeRHXDAbeBTuRAjpRx
jwFux+ydibGHkVZgw1ur42E8RuWsBotOHMk97pKQZNeL974IiOPI8APhBljzm8A+gjjsCrBbMOh3
Q5SmXCyDwQDQUSSrtMkgBhtI/mUBChEV4nK/qW9uE5QRZiAROm7xLbeX0h/oMNe3XoS/Y5l0+0PK
Nmi8R+GvGD66Kn2dzkseXOZDApn6t9lmUooj/HnIlN9te/CfaYySzYrN6cpSL3DawhjbPLu66TeL
6ILyZwPequFonZebvuenXNpAJuaOW8ZTrRHjdzN2J6LFmVWbsmjOHPsP2m5v3/w9KABUdHKnZHLy
uOQjwEZxH2j0Hj7oFXPacHfMsaK/eQ/PhwEiWFNoSIeXEAapKtoyY21bkQDQvkQlm41qBlnYWpxU
jTzLMhLHYUIsbLlMHowIGWPiXpjh4ek810ZwaBdeweGVT76a2zqcLguezfroZiqWe1uYZftIjCSg
8314tWzOa9Sscs71mZvZX6RVhgcoMw8x9m0XGwEVQu8hJaeFYFl4E7cCgdXkVF6jeJ36J8gdGhwc
gJTZZv5THQJGtPHcY9o0KpVtXWgHER4pxIL7b4V0+BlIvt3e9Bdy+gEL800ZvP16TUJMTWUS9qs8
T4GzjmflB0+NDzfK6qCbZPPZ91QkIDLRMJrgP9HHhRpUO8aUvKrSezsGsQ8s2ywYO4vK5iVPS/wz
X8aYjTShzkgjq1AbNCTm273uFRVClygH2QC/E5ZOwQcxPBLb4Bd3/2qw1iRV4jQncwqXuJWQwLre
WsJOZ1fsLzqP6IRuqVxa/u6kicM1xvJmWOz3aI5WUziQ/udEcXK1JlHW3C2B7s8/z8QiU3aG1skV
vnRC/vaOj2/6VwK1B7zAPj5TeQ7zK8dm+ZHOSHSft3WCpxKRiSJn5uSq8pClTl+AZzZECt2z9c4H
ifpYlzm0fhNkK7jC+uR7D+Kh+6naeZpvIMMM8LgREFCOdrHJUnmK73s3CdY+1B4Y2Vd7D7NRSsoL
7XmUdhQwf8bjvxkecmGBFkuTX2MgpxNspQFq66VuJ7FyCiqH3FTPlN+/UUVwEnyPHkgj6aWIuyLf
LP7e/hMOqhrj/ntD83sfpwWXzRtWJj04U1qPQXG69a3uWGl3XB0p1cH+KP+01brFxsnVdf/YX9fV
6FeKlslJ0H2yQplXFLrTep86y/Aez6cEQrvb0eTVJOXa82XBKcasrdBN7rdRuvYSufb5nFJGTM7t
Od7m+OTsc1kSOZi54I6I6hlBeHkw9uQuRZrrux1h0f5ow+lmPpXRaBN1V4ThZ7gDm/R/yw9jEmeY
2owyrrTRws/e/vqXJ+lb4w4gS+IDXkrXlGd1UD3v+2Mo+EB3Vw2tLLeFzjjAhwvFKZmmw74WaZCb
FfxyG7DhAqvyoB5wSV0pwPPMOguNcAxIHbjGNvxbJl/Ek+J6/KGQFV2YzQArheFwwNcnLmWN0RWj
3wgAh66Q9hezFsG4xvLJlq7ARgoICTWJSMMyz9BqCgzCe+S0OvHk4XTQB2+3iwcLtrBTPyBabZTU
8ZJiB0VoRUa6OdVmP+PHg9vNbLMaAtC8wuUXujR+AshxztwxsIan+UOseK0K6JUUXQDpapUIITok
0+D5itXoLxc0aOsil4/1YIYOfPwXmg8GlMYJO2eMSm03LTTjYnxocbAqQsLRZPgSnc6xS7Uv82EA
mREY84vfC2nDB/60pSDnlxxT+wQhF5uoWqeJlAqQ9TB8nCndFzeMU03uI4bb885aEK3t2KxGTUe+
cShNXRYkQcI4y5FxHrXkiXxZsBYDKevTS+T/QQLLJX7pBjuQnvQ5dYBlzcZ6oeaQpKhO38FN5SV2
jG9N0AaXKFxDMZ1alPv/zYyNGuToogEGkzvwYpnl6SV7+JK6bn+0UjZMN539+NQre5i7Pl8XzbEc
1q57h/Dl77Moe2vNVIHuEIbtG16PSAyVF+G37aZTvfxUKVN+zoZWM5UXvJEPBpY1Qa4EzA/Z1WpF
BDE6jggNJJV/SYmKIBfFafwzQbXp9l+sjckAjUA5UUaBvnbzrLIUxNreD333BhPhp4n10iKz7TKI
d+e5maQ6kkdagkX3bsc8ium3CcC6YQs/3Im+rriBmEeiZ6jdXdBNteAZ/6DS/e3tSMImCSmTrLTj
YhAwFv2sB+QhVw54dPMhY6FYTnzatBf6nLalUUeeCUuHQ4RsUrhOS8sleYd6EPC5CcPCBxuU45Vu
KoiWvUjMkFZF2hbo78hrc8317yHiaenclRNtKNggCvj5HxTXTt15uhh/DhfVsxgPigFkrPIK7tSa
KBsbn2lax+Hj1MP0j2RhJFxk3X+AIuZSxgDpD7QCISqBKrJQCe6JHedC9Y7dKYcmJL1HcjSXpmIa
DJn7jt6VCNg4v2qKZuIY8cFQPopBKdvy0SBJbZlj47XFIe0cskSCB8WflbrcoIORQirUtvWIqoKu
Qu1YIz2v2N/neYukT+LJrTAhdTi/kSVeFmgETfDYiX5pT5e4bUfhQ+9LIzgGN/dkk6pgqpjNIu//
FPPSkrRQ2OqLgRPYUkPeFpzB6EEom5A0Y0cJ+e87yA8ivNP7FknwDEGzrLBuQvK584Aesz4wZ9q1
69fFfDxlen9lD2HJfybxYjrfxKDflgpvJvMRjvvT9Scve0T4rEQqUaNUla0B5OMpXiX7HPlo852X
u66j/YMwaDPfqV5+yj+cd9sS6WUIxUKyTEPwxUYwX6n9a27DxT6s2Uxd/ZqvB4fb2m+ZoUIY+04l
ESM5sD6BFIrhApx9jQvNs9Kq5M08SeGwuMt0lDoL5HS9U4ybmvBQJw/cTogGwDoq7m1qOT3caIRN
olYTYpHxdshAjJkXSgpFBdP2ImUj+y2jKtuDhC80aRXoYT2WS1vpTHkfx6xXC/J4HTawHv0AfR04
dt22+JWulIXBUg+PZ7PJYmAvwXg8SgCsLvl2GeCRs6l19/2TmYx1PIe9uYW6IGY1LKSyQBbXr819
rBxoAaTT3Qzw7iFx2Ti0lEhlELR3/Yg0UqlmhRb1wAX/yzjsBEVu5YcFbLeFAxDZflro0XXJBe28
D4AXRy/WulI8AbAzfySshzD9SzLc/zPB7tMicQAUL/mQvKdBZ7vPTbDiVgx4aBrWawByEy1Lf6lx
fH32OrkUCPDSu17zA44ZI1qeM6VXPrLRbFMHOA3nikzwXn0fdQIQOtI2Ux2z4OAvdz3wpUt1ljpE
M0hwMxjpj+WH8zbjq3KDl5Kha1O3MApjPy2SH1njM3/h3XrDnQARMX6H2jZMfZyoZfCjJIg+bmHT
1H+IN39R5CXR/9u2ohpkgvcR6hibnuTpM9/B0ty4XwKD3xF0Mkc9BqwZJNaybbbGaT3rLjZs7rPD
gdSLhU53Ht0r/7nk8RRT+mFgSgsOVPCivT+ZENEYO9Al4L2TOH4UrhMyjC6DjeuWXI/4Ll+xis3s
YyLad580U+7iEFIfoVCyGgZkp5ft5jEylT3gObGKqlTUYXq6txheGUYyRzc4qAVi7KdiZvvO3dUL
XN8bZjBOxPcqMTtIWhCW3obFcLKx/7LIwF9wFO6WlWj3h/jHV89ExhENOnpCEYEoEk+P+kQ/iX8B
jyY39wHFbgh9veT3CiH/hng9ArmixdopKLh8X9nzfl79oQPVc9wskNyY7o+qLRd8Rupv2tLJsFjE
mroQiBrrDdVdC8SAEoym6A5He9nbgP8HtIVcXUvOUnBdFJjcf8zV5RGd0UlsaqIICFV63cyeG1Bn
zBFukzq0KXy1xy4nZdWDsT6EXshM5u/GX8o6AsZDhMQXHVcKrviVHUWsdwH5l71tRbrlP7zlBme8
+Z+Aca9FjdTBE8JP4TfHLmz62LkCibvElA4aTHlC5I+vRnB58n5gjPszLHEj4ruE6iqPf1UiIjpJ
FZNnN4Uw/x+toAncVuwKG2FeKQE84CuBASS+P1f4ovnwb8dvmJfPQkOANWp+KjxnE35JqvwjCh6g
OnBmzWW/L6L/28EapjbptjmH8AjmR9SK3+zvxq8qbOMqUgqBtJ4xmyHm4g+9DLyB2Bsi/x6LtoxJ
Vr0ddAlRbSfblqSgnSaIB42OjjGxIfFQZoJsuuIl9GGC46obSMlYcrJ55J/dLw2XOBw2TTraXOcd
op0h1404zXwUIILparPV68bNchzDXw2ehCI5yz3Q57Eou+3eGStErVeURAV5wOTUENOY3WqWm0Iu
Yn6CIinAarVksIWx2+G4XnqYrqkitNzGUCxyThbOCrzyGuoWUuQpgHGXIdvUlmSwf9lc0+LJq0lJ
E9pg1xSd4hf2GEFWQCrN0wZ1WIhowLJk2exDO2ejNXJ3SChD8WtVvWxKvYdx6w5umb83xu193YTY
LX2AYluTvGF/A3Y/u5bvaqFussuf5lujn5qSBh9pXQn3TGoyBwB/JJdzop7/C/iJcauPjyj0AXBK
UjS75Pg6PhPcwJoqSWMQwgtQ//0huoG/U4PYjmIN3YmxyH7cGfqCZJ8NuQ4ngtr/AkXEr6p0fNGn
OFj1mGbph40HFXQuGxpWhLaphoxYT2Yw2mqGg7nQgYO/Wn/hjnQ6kovlNQ3e2csgPu7rZ2t9TB1G
QfsP3WnQtC9ImJqZP3o3Mv2HZo900lNRIQY+LtjY1Izm4kdOIP7d1/6k86q5a4jOoLzjuf1OT8oY
EdppmiKHWXXgAOjQELCF6wxsZ6M7Gxrl196z72iyE3lFqLMUYOS+oUEhq9UFFCxVxvKRGqOCnCsD
oG1FQIc6dSskqDFBDdfWdZjATogTeN2CdzyyYZ48Jq9f0IfxfCGNGbfCz10tosDJcrErkdSNjrVc
EpckRbXVLwZvKO+uk53Fc4+PII1Ixk38tyWwhVSL8p3TobTZDwOZ8UIK5cqFamaZ04is0tL/wFbD
rKJGlcYU5jW2I/zUW2qNMP0yskOo3shqIYhHRCaBYpViAbCubooOJd0cCbljKFRkFScKKbAG4TeI
Vb7B5RxYbP90yuTHhfiADk5aYJUqWbZberRnPmYci1bvvF3fOJQhz5u0AiCjKsaa53MQ++d/hTo6
AiACEEdvpxdypQE0Z/BTO+mK4oOFFO1V9YD956p69ifSxTQWkMXwkuW5i0fAEdD3miZ89rjO07MY
OejD/L6UEPdFc0ungPuAh20kBcZ7sJtqujP/IzRsXaRtr0aiDhhFXr4rso98pTk72eIuikf4UmD+
kQAyg7YQa9hjpEQKyGrnXUTFvA2xHumBsKA94YcK+IyxpiwBPIDVyj/+CovX8fQJOjLDn5VjEJbL
6P1jfTRwtdjK/JfJbmA/6CMxiOPxyUG0FST3/Q6VtPijgfaGkadk6cvU2nTAc9HWa7ut4nrKDnIG
0HXkCJOd1gIgGawOAGWc7mhB0xyW+/dzwG/0lJc7+iXWJCwERL4x+m6LSOkzvQ/Oza6eeopmKn1A
tVD3Jz2aHy2eqqWSoTeqJBit2cs5OgkxEOaaM5zuQIloNno2ZuybleLtztFHdGT7y2xoGDJUJPhe
9ThivZxxv7c8UbtnXmxuxaQWg2eKoek2n1Zr5R7jMSwN2FFKs+Su7IdepDXnemyh0KH2+KHmF4Fm
q5w9L70ZdDzApc5Pc6xuimdRw+QNca4nGwlL2lVYx0a+6I9gzQTdBtuYQ8OZ9lofKKJMRDxr2SJK
D4RDBsG1xcgJXRJTyKTq6NyB17BXdR5jOLkgWvgpN/cDyu1JtE5mvtLl0Nked+HzFabeeTuWRVE3
PV4cdY0DVWoEFyfNMFdyQv8m2EnWjNrXRZVmDRdxSzHy6M44dAHWfWTrTuQYvmjSOCwjkZNr4qY7
1ULJfnZcBRUXIXUTPQ5xt/yGkEInjX5Zlm3n1Wg1SozVcGSRCyJBlQNbcYJPa6ozQEtEKL1KEUYy
7yV3bC1pb2MiMoxrEjzIFeq8bRPKiK5CJORGVvBW+oox5HRtQV9WER3kKU1LUNzrjy2qQWpyhSbC
eegMn5GiEztDh9cxqfcW5HjYLM3OnR+fix/WECAdTi7Ob0t1Ylrj/Upt7E1jJftIWljDSGpvXaEQ
lG17gFvad6mAMk57AjDSiP5Jzvu/X/IEW2GYrp7OI24VXXRPYlr1hAMmPyFg2DM5oiYFVSKV1ika
k8vsj32FvGZjiuCgIMudAOogg8yoE9elqjFfoJyrUFfONjetYhQs1bgo+oh1J6L0ui5F4wTHNZ1T
92fKY/WOn9cOuWJYt0ARg0DJKCB11NMXC7RGxrqStS++/1btJtvawid/fiLzegjjQv7jkA9O84Sk
IaDWgyWbsQGNzL7PXjxpVB9Iu905NaL8WIp1LptcuiK3Xup9WVkc4+kO5+3vEWmgZSEM//W8B74H
0WuxBDCqe9qNxG3fKwnvBYGWbV7TbMKsqjpY3XAPMlCxlnBE134I/cYCMaRvTfsc3BxC30q6GUZs
AajD1gl3ZTVhTrGdMZwFbbsWpvNQfvqfidn9+I50wVigcG/QlzVGL8LTW25NXfq3fyBwaa3D7aOM
RqR+oZdCmFGwoSKN3svrDMm4lEtcqfv87+7egNpx7f7lAIJ8/sxJMsaZ6DNxlgvvH4UUxUFCLql1
HWDxTpstA0q5QjnkQ3XSi4PpUoXAQYbOWLpI0T8CQEpkgbvJBw4bOnvZMmt4DROvjW3jP31SCTEd
XKROriA0KJL9ZPOk2RJbcESTIKYwg1vCu5+gZ1azfP0aT2jmLEhJfXVJu4QDllwN+R0bYEggmiyn
iXvrHrQ6f0NuwFkoAwVfoNIzZERchl1iDDpdx+98MtzUBR6xwoA9aVPrfWY3Q3qscY83C/Ngn5td
jFf71QYLzmBjT10EaztHZ9rrODV6IHvY9EmLGGjA0Eutx8pCwhkd0aMwt+VxNThwZ/34064NeAzO
3p1jn5sp6jX0rTd73iJOhGUgxfbfMLmaQQar3LVGQWSsSGgyTlkYoIrI1hnTGDTv6psLIDyjXTtz
dlPnI87f28jYycG1hBrHI12n/63OkCWrfNynG801dz68xfzfaFrAFtLUzy698W3xnOF/agrLrQi4
9h7rhGfc0LCLFJk4s3l9m/XAIK3xLytFg4t6Me3NPY8NuYcaHJNcPNRHR9IJFG8qP6smwBR7Dbff
lrOdYA+ET8ULBEfSoNP5dLdtYQNtqN9d2vdBR9D8Z3BjejKgxGgsJZJe+bAuFpkraBc2HEtBV4v8
zvjr3RZFfqHwf7wr2FGk3N1RDUCq2Xh+q378wsCTzpnfzSNGBG3lmezSPO8Nfxf5NDrrO0PXdmJc
DzuCu+E6elWjDBa2wuO1vC3H2fuz++nqM1qAQKOSW9B+n5D7kBMCPgP+Uw5tdM9ohUeksuZO+c8F
1QiQXaAinkmAIgGnEXo6qr/+csLCYwCoTBwpv0GcBgAWvrLHQRbsSC1jcraYWk7h5frV7Dou12DX
ID8QX6QTKEAcnG6r4FMrMKn1K6ZolojRKoq/jHVvsXPM91IXkpHSFE+Eukk6d6F7RC/cSyUb0Gch
DeL/bINFj1JtXceMe0Y/HHwKlFlKPyB3nwtxZSLH7M3mkACAW9M8qRBNPwPJu4BWrG1c6KdiM2pC
g9IrKA8+0Dy3xOTQDqYiI+Fpgf3nWQDlj6P40L95gc1jqQdIXhzQuyTV7aQL7YI4hq9h26woBP3G
WLpN7ESKfr7Jo1qI0lOTQlk7pQBsCzivqC2axVA+crYdItv+4Wh+38o7baEiPNJqT0kNmp64Shx0
rbr5slcaaR0bg+/OEyse/3uvfOsz6ZkPVwBW6SoEijIdmQ3V9LBb5sIjF6BHb+XaUHUB3no5l6pJ
RmVpcXP7M2jAd3V8xZ4CzMy3zkVIVg7GWudnWsSCva42FmElno1hGOtoNXgRSGV1HBwx8nt9ukp0
f7BxtPqTd8dTDwqLfczVqtODSh7jGlxTnVhn5u+cCwr0kI1/TCUArADIJ0ZPcY5t59uDv+oww/k8
7WCZKlhLIKoRzf3ycASrtFcyiEATDyEsC71ZzleXNdbofch4sEWyZxW+MOOcoAcTI0xO7191e9mL
xHURr7TvUgYgnCk+RPFdTDAS98joZ3SvUiXI9EmvIl7T7HMw8TZJSnoEt+0b02lXtYDRQySrPchR
CIxNk/j6BwAMqNs/PkguoHm1OFByRdT92DP1m84ZDJUNbG+mu7DnzCl881o+eDnY1tF2Fmp0zmwG
2MKbcyddZxxSpzT32P5iUlKMTgUIYaTrKvqrzZkR8qSerhlKOJiUdFeKBM/3QPiUK+fgfNrQcCCc
o0l5TxLdhreLgaViSHoirPdbUvBsRM9aBBap8+4M6OdtpDIsmN44gPd8NFk+4ugrg4ybJWLwcDdP
VB4/qy6c5olgvbbEykj/hk+EB1Rr7rZrv7G/uNyJt9VseGQ8/3Gp/acmogK9hE36W93n7dqvF3Ut
xc1XdQZ4ODUbaOhlioDezMTClx1FfzafMem10tJCKZY/K4LAVad6ursd18VnZdwE3Oo0od3F8Jbc
2q9n6K9f7pU9FCxx35MRHq7chKfwTPBGx7WVBz65TfwTDCnFcHd+JikjtRrgHCwvxxJRSj5CMJDS
Zd0shs0aTBD8bsDystGEGg3aXTrwDJFyVG2ULO0JuQz1yN1e7+J7E3QHtrfySVyz39nLJI3TZ+2b
3B0EjvlpV7OsBZjoc7pkwt8mwGSFvFZ9ZDhg7nGyeNsp4IYHGkd/zHcVDPebVZ1FFNKwvr4HvLX2
K1porm9wU4Tkf8EMdH4fWe1KZawBWMRCfQYdiPnUmGear8AJbKDT4cCqaGgmoTFtk82ECFvOMi08
ICc0QiZ3t08TUUN5pcHrueOy6AGZcpVivYATQcZ48GTbSCS4LXX7L6Of+Ow+U9e7Lt1kbBHUqoWh
6eIBeWOS6Eo3F7RIoXeb6TwZ6UwVEJgAqQGi6ZWb0PDHZdoHL3U1IUYbFAYULhtQkggtqCbPS7++
P7+BF98FbauKRUKQU2VpEx+ZYgwRkA3SAZiqpGZcWhPJpKQCqoc4ViYs+TMokwQxBIZyvFEZTMjZ
Xo00Q5Ofk2ckL1sIyQ6G6Qf5yaAbazdbbPbe5ixcQm++2LM/rtj0nW0OT0N+HzUXk3e/msi8dueo
Us23uxgmKQPznYKMFhUi2RDepjYOPb8D4Mt3H2K4BvhJ1/xfVi3TtVlRC5xHuELhdcNqkf/K493W
Zjrq+yr55LTABE1SwkwFYlt8zHhvEEwVB5ZeOakZus8nUGg+du5LN3CeHdHD0hjhkkM4KKUPbu4G
9u25sZhwJpR6fughfoNp2zpH8FvkAJhkv6bAuOO7R+U+/IOx4okyRS2slH4E3Pjj0huFVOLQ820N
ZqO6k246Q/rKPCG6vn2qcAgxJA/GhorFye96GP4OlDSTq3iRQurUa850X4oYk6s+5s+M0Z6gbb9c
DfvIVJdY7lyhZlG/45Uh9OmQGnA3I8W8Kf2E3at78W6+F37NMxPLWDWPjU660O7NQBlQl7iG7F17
WOo51n0tjGB6GtNQtzwTZzi9ssVunBDPRoO2Ac7LEwN66L/xY9sdNnavr2e8LlE6jJNbhMBA4lSK
UWIbsYPidUCTjA70dyf/YiyNc6AnBMOlLpO7BvT6mZAy4ove/RxzcreWBSdPkm8x6p0jfVXqiEk2
t6Vl07cip00MMuoPHP7rZYQlFE+ct9yOMqCFjPLjrWTXQyxFDOK2d5FTX6+7KkCDSD9D7F48Db9W
18DPYCtDGPdFsDUrUkSxBTl/aD2L06f/8bPjvDBSSdiB1hsYbPiIPleQqaJA4/C6zYiIkl5BL/0o
7UiUDnfAUxhvIeUAT00dkMsI9GDDb4JLZydk2xzogzPkUHKtUHj+VLtiUoFP1cOQ3luOdWd3JfXx
Exn1mk5rj5bjwGYfBX9QSP+kWJu8NZlwWVswD0SlxiSuzWqjkwlYwl7XsaAxoEaBeCk8bayVY/Ef
tV8/rEslGm0iHVS/GVq5uG8/ZQm8XVdY+KFfZsl9txHHyLSdt6TUtKUVo39jyPs4HP0eTl3IH6OH
RcIGUcgCyvSCnF5DCSuqlJHDIU27t8UPmAyS+nU88XXmBAPo9U4w21WKb/AGZtDAUcMZ2JlxUqZt
N1f25pfkVy8gmiJN3/dRGr0Fs3vgdT20RII1kreCpXegaKaAaVDmh9/Zcd3avst48k/zpfEj2lcY
cIdTDRWgFNOVnaS/m0H+l935nfRlplUWS8t8qrZhtQwBlzhXMKotilQHDpfZsJE2VVmelKMqUgie
a6CXZA4Wjo/BCnS4HrklxH4iEzwg1lwJUyr6VZexqYitJcRrBzq/B52A9MYb78ivX0DC+prOII4B
JA+xVqXru3XBottEu4Oo4rbfN4bpGs5m79ABV9cgnjxQTg757kjgtf/k8Hmr+aCh9q1gQnbNDtpl
ascqtRSlhC9reimVoCtPUJRe5DEY6TI3zj7GL0IM4IeMB2nIG8PRpz6XOdx0SARKRstNAKS5OCxR
VEQ6zfDnhnm45m/iuK4LOpZOwvuQQ46MASLRxAHxjxwDoDyF31O/+Bs6MJqz6ni4LEphfiex7YHn
SLlgXcj7OwUB/CCGkUeGtCnvAW+TdIabc2v5XqUzXjeOeb1RsTuVKumOz2DMJkqGno+6Cv5/eCVi
SW1+YR0NWJd4Cz0fmQWW22Igc9puZzv0ugODRNU7PRdMb0beDC9yG2XNTW4IUNvsQr2W5cJwaBRj
sLZ9ddQmHYYJEbA04mFV4GLkdD+4iPAywbloSKgpuwddYLpMfwSb72b+UqcwViT+0N/OniuoqG5/
V9ll5QtsVMGRg3ctFw/i12wpniqAKPRBFgxiaKrKlqWTAGP54knnd9UfrNOU/ZF6w5UFMEV4DNtW
SIwJSKMEQ6avvoS8zimSs8E2VuDqdI8D0i5Y8XJkUHiA7iXTmvVZGYlp8N16lXbc/YM5LlsEupTH
QYUwuqg6/odvzbq5B4Dct6fi+neglrzVp9m3uJWDiGfY0zjPDo5ts+QSy3p2xWjESKGqt465Uafv
GMpPL6N+aJxF9IiynHIcvHfD0I/FmDMrCT+vR7C25x4SeefbeUJ4HUB7weig1O/3ufLfWO+piBNp
OS7zwRbwqGBXS6vgB0pHFirTWNFtMNSeNNoYhAOeivflShMGtbsAI3oi5HpuKF8BSeZQTmOOJttF
eQiMBcoBb/pGMF7sA/lQENCEWdRzybJNpvcTrWXsS5YtuzvVTOkjqiv9EzU/YiEGNjZ4RunpEu9C
TT2G8YiNtAqsj/ThXahXr/pnxQqMRAYiug4DfRN/PGEKY62zBYd71nrXYFAH5VKerkge1aomejZl
klw5o222YUMb/WZgbqzVf4udbOgaO03cRpsQDlfOfFV+KJ5h0dh70J9HSm053G9jBzCmC93wP53S
nVOm2uRTiEhRkUHU9frFUdzK4yNAGVq/VdRk051ONN6A46pNww/2WyaZszRm9WC5fjLB3CvG7mGe
yMcoe2shflK4tzRPXJ44Rv12RwCNQB64ufSucPOhYwqRylrpCdlkJsClbZMfj4c20I5HYxQ+Trfp
B9LLuNDFwKLUx6ENz5BaRkBIB49suUsz3qH/8SGHvUTbLcR/i8hTXAnLSqjjyXzEHE9ipG4DUh4O
oHIHJ5BCfQVbEgOs4jt9MN4VrKCHKnX9g08eDl7/QR+dc8e78fSFPcff2OEQT2kcb08a2/di/nSX
EZ9DwJnDvPzlbaNMG5jjfIvaLuGW0Lr2e+p714QqIDScEEN8XLsfMfCM/sSUG7RFLiHa1Z10ylWH
JdTFz+N9JGuwoR5VYERX+MKtIlqxEl9J+Ou2ZMRBBV3A21mV5FxmhzxC8lDKpECcy0MiWmhStwd2
ngaX8LD+Q6sRE5F7QCb2wPsO6HCzYRiDnYYsn/iieMme0dkMAGUXSrqEGqQKseFnF81L7QvgCNFk
lGYg/xvEoflcMbqap15aGurev74/CXo6Hjwjc0u1q28vy3k9zaxZRjzk9PgVm4cfH7EOIVyYZ4j7
xmOHAumnHIn1j/i/girlzmoFK0BmXmAFAlSzIo3W+Jjl6WBJYz/GkFDazKWxM/ceOUlKqQinF4zt
MLZUZkoHhIAoP78lg22F9n96edMW3/YW9mpkQJ/f3rXpERwrFPMh9zbcVUFd2dnSmpMzpridIT/y
3ONyRNoBA/RBwZAbSoQYe1KS95DokROq7KxuywvtfxUcYtNO91BRpSLwWOB26s3tZnydg0C4nfnO
CNwtAVjpJBJ5/JIWkJ5AEgNBUvIKwVdY0s3NR+cUKRpnwOF4ULg+/91hcHHnjS7HKiBqrSsIa+WG
Tn/r+htHIw3vslfdDo0bZNUboG2BwvrP8oljq0xuKS/EreXvEVoCSMgQYq6MJ+wZj1LJzL8Q2kSI
i3Eq2TnEI7PHMaxdOElT6yewyybd1WPdPHj7CD6L5cLKW5isZqh8caXucwlAZvk6XErS8idG6GBj
SuyKqu/XkgcqT8UiHQoKnEdEp9zKXjdU5iolyHt9a+8OB5pehzuSzz/Qo01+M5RFzJj0GLNLYpHT
aQdhFvPTe1MtyGIjU8raN3M58oFY6wiEJ1Suh0UuEzoFWQTZws80gijz6uEI8vNiG3EkX+jYBG8E
WHU2OLZkgpmdAQHWvv0Zm72qfnQoJfsI6ohhynpzTTuiS9P68wDHVoBZZNfpUYfZSB/v+bAa0EYi
JgEzGCojgbmca6kN7iGdJRawOZ/OyqjVgip5zTZkpAw8xLGIim/nttFVWanwyC3PkVflUrdbL5Zu
eITYIuJvYCp2+HLBi9+OBOGK7ftFU4nwQetVE3N2+Pyfjr9RaE15aFIMOC6hwYUKrMN6RPiL2aHq
f7k0YgVXXlkm+qddVL44zwRMqsK0eSljnxShIpmjIcAPrvYbS72TMxdphc/mZTHyJIyOyAQcVJi6
X/ftpYLFN28gAaiA7HMwvXtbohBDN46+vFp97S0W1RK6l3p/bmUv6Qd/egVwqcPN9ibzFJhe8TJC
qSTZdccpZfuq+A4U8YwGizOJU4MgJSpHnWF/xBhH+rjZcaxteQitOGkeUf9SbdoEYJgibOxZ6hC8
pHboKtDMm5MKTmMj++VX+120Cpnj5027E5/fX6uJJdsVd5ig0thFmvPKeIEeg6Tdedo9Ifrr5sXp
c72DW96SGZwI2YllSMsq7k9HLfalyNqN9zhp8glvSkLe/ETrFz5/ISDoQdde5tP++74GdzmcBbeM
DwTlhA1EZ/E/jlwT7Wti8iy6qEZ0EHHiKQLFiSr8J5LfSwLi8A56xHoJEHPOz404Tn261AEgI7y6
2HQRqIyUBoT6EteEtMlbZJkktYcFvCyyrDUNkTaD5S3rIpk3w2aZ/sirJ/TkMc/CJv5ZKzp2648M
wGDWkdL1+9L3R1f7lSbwtsI4WLRxoYdPUI2601E8s6Et87phA1h2rTlFMbLoqDKiUb6FyKXcFSYX
pICg5dG+s652dIXa6gdwfBVA2w7QBwhacdFWSJPAqg7SdwIH9KMDDnk34NwWTzbJ46GH0xMPPKs2
daqMc+4Lwn8RZCqTs6687a6iYVgfRWHlfZl4l0AjFZxfmcrUF5JMvgOL1nLYDkwOZHDSdme4LRJf
8Ps66HIck8cck/gBMCtvYsQjXjsGqKrOYCdbcvPHEb6bp/3R4ZJUy+LA5QP2Cu7Tu2pfWlTj9VaR
qtLcADOUTgbjC4SKHFVQj/DdeIJNEyPlHLWdR3D7zMqAWj7SMpbahj/p1vdolAV4wicVmrEh+XRP
n4t4FYeDAivGNYz/+o1QlmMzA1WAnhEULw/6wYb1apVd4b4Q4JP/qSeQ7jeJp4T0uvhPRDy9VRkl
RijBCRYTkKZBM+zbPjsnf6RSNDFz2r26x9N2FnI0B4NQ+Z/WX19VYgU+kavHglhrTkpJuF255Onn
GAA3HgWVJT1SULwQnp2dXFGQ6lnH4ScAjT8ofAgu6afR9y49mcToL/VlFLpJiSvyaC8TJE/YhAwE
QhKEyd9lw+ApXwMVBpRVnN0ZOA/03dNI++2ZPahcKpW6dsP1i3fHsvINhBa7Yv1XdT0Q8x5HaT0G
55hsrgVO65LyD6liXEG67Y8Txv9c1bXSjtRKz3B2NLdB8vdOVG1ic2dAjO8dnCmin23/mj8GhBFE
aRcTyVgxKY5oJJHHk4RF76lxk5CclcOS9lAcyvaMwfzBF56rpasKfatqONtVPq5eNxiWaGfzFZa6
6u10Jy1YbWV8QoNy26GosqsIWLN1pGsljnfh94mRCZAE4mfD9pAcJNoO5YKdl1/TBevYynKhqwGB
aM0+1aIxEnlUDS1XA6GhXm/R7bmTWobI4NQduPYUmvxdrYzU2mG94GAEMMxVlUn0T9jSgcPf2Uri
LXMIzG5Okvpol09EmLqylrywwZvQFvux5PXud21BwlICVlfqXOj8On0mh2U6FortC8rWbXmMFwEK
c+Sitbc5gSCr4U7J9zFM31A+e/Keb4jeqmnKEfvzn42w/x4U2i5brE8ipNPb+ID1MDkdbJXC+mqx
OZV5VUXRThTraDJ3S9m3zG4/amIAhlJVG//GzFGrl25XO+doVjuYwetEIjjPfTZsgytwPKJPY+Mm
n6+HQbMf6DJb1X+Z+joaJRK6K4sUtBJ3EhwDVVFLSPf61jqLQ8ztZtnARRrNnQvcOLHh6nSZh5lE
uaVrimTaCeyIYoexvHc41G9iBacXdbwFcTZz6psWe+qTYKQJTBJmpxOs7QJ2dEhk1pL/uBtyeHMW
BC9SPX1zZ62iKhcpnQvv30VE/jbKSFmL3R9DxbzoqwfQ5rkoorXP0h9BH+tyERR/Tl+EPCkJGaiy
duabtwwjv/OVPHqhaasAa7A+YhDUTjflk2mRHTIiva1T7Aabgf1TXS81I0k3FYKzF56T1a1vjvNE
FZXk94eBycb5SsnOHzTCMzHwN5qnBcv9fAqYRGEWQv2VvBr9R78rL5zTG1AHpt2UIFop+xwWHNoX
Os80DxQEHRTMgB0s4RtT/7QCsap0i7daW/duncwbNELL+vpsRj0D2Beyw8snBzWXWBw1qe8n1Vz4
edeE8pa68pAb+ktKhiS649VxIRtMRp2u0glAlMpYr9Vn8Cwf/HnvT6EgO+XW7Xdtfbwx7feSLiWP
wMyvrxeepe0SXUbT3o3E34OLF7GYPbcpDUnIYFfsfvuZXv0Psg6yUcdvXmyWFZh3WimHEbxSgda8
Vzhpk/QqQMjPdWls4VO/h7cDjJOS4V2KGhiY5h2LIAXTik/YNixD7KkPMCYniCfMhWlKRX55kpYT
Hm9BCYdfD6634xxRjZqveNPWeTunl2lFV57z+TvGJrbfmOPfyvxo4ZwyOZNhOrhV+2Y/Crowq0kI
keg7FL8Ss72RM0TGEG7LZzfrrZs0n2vzFsFYbscqJDfpR+hbq4dkzPInVsgiE4XzI++r/VHMkiQU
lh2xgZI7OdtPwMmJgB69Rve6cBYxCzqAeaH0Pn+FmXeApk0goX/LOy2f8ycm9jSTzeM4qHg/YZFx
3lwpZkXxrTryC2GhtGkOLfCZQ3Be6VLG6h+AdXBVWAQ2B9NWs/UD+xrRzjaKwTzjnTRiEt3Fj1pe
tfH22LKKgriXfhdFyh8mpd6ePNBBjDVs8UVt4lC89mjix3Yys+RPeLmncWZ2j9FEkKXKuaC/PBKy
a2kuVBQEy+G8HMQSU53N4LtSWFMSDfRb3fpIcIN+Ah/v16QpL46cA+XlWTMd7OPJEAn9Rwxk/sIq
GHS3VYVILqPRh48/ffCOV95HuzNHncIsFr+Dfu4XQIngCzz9Sw66bHWz2z+tSvX3k471p+LAyzFZ
++YTEvEBOLcXLrfRzc3w4FgtqtiRx7DSwYfUP1fJOaE0+0HkGljP7qsokQMvykTaRy0mLq6UmjL2
dmHmf1dvD0GTmKHqJ9QTpdjyCfJUx6H4iitwLg7vSxjIzAmuj1QCygZpNN6zO2VRlOYNTb1dY5f5
BfLkvN5o+k6eO/oRPMABa+ZJWHtjg0F01YjCyQhYzM5L2eQrdXBDtyyD70jlLgyl7czeN+MReNbE
Xfm/uaZ7CJrucmp3p3pfQHhSAt2BE2Ok4wLbZ0XeY6X+utSMLGE6IgiPTNB+4LZRNE7riSg5TuPo
PqZEAcOkaSkVEPK7qW6cqjYdiNujPqS7FrHS9uTRqARsm6ojnOrHmfYSu+4wKYyIHBQPBDBeHATk
bCX8jmwT/FWulUaTX40NqmY49e9+WX0/0ieuM3dvToKJG5HYdVeQ1MJ5lGSuqRPRTFT7TyBWyrKD
b85gtGWxUnLI/LFYKu3R/Ng60jmuXYFrRbRQ47KLFIb17mR/vBTcU5N5rCuSvYPK2AFizxjVZb7f
a7/7TN7lVBJR9Ka2yRXYvXsCP8PmTubpCENHW0x7ebRSsypajoxDKJO7eb8lFYQfuSb0977r9Aly
ga6MbtqX+OJp6LYqDp2sgPd1VVIFPkHIkK7dZEob+WKIElyNcN6bVMDXsrwD4gs0qTnTNz31W7Bv
OCXNMKLdbKfaIpU92b4LzqN0sI5ROSD+IdcIRy9eqD/ME+URxF6gtcTP4pjTWXytLhoqGULwMkkS
wmmvwn9hjH0csPgwQktXdpvK5/8i2jokacHw+qVwydh4g+cI+s4I3vPjGmmROuI7smlSod26h/6V
RWKoDTtuYyMHmEEIBU6H1kR+0lccukpbx+DSWs4/uW/ml8JZWQPHg1YkLwalfvdog6T3PbaxyZh4
fPDWQrVrso82thUvnKy/FnLXCQKu4IIz+Lyn7ZVqbIXpURfVd7AjzQsABizQlz8OWTBCdlCFRGA/
c8AXbufsMBl9dJiQFyYRfVB0+eW2vJBshBYhoMXRXfcMOjNT0yxaYaQMGeQbFRBEocpcCKXA+QVm
dKxv3eb83ICdPzZT+IM6b6fTH5U+CdzkkHjnpDnhSnq5Ka9YU+9IeUCnYlbVsxESjs9fYO5FRZIb
OjFMQDT1Lo8+lw+GiyBm5y/7KWl+XE9i+eiTkKMmMSNXFqpVb9Q20s2iQ6T9MPbH/FSQMP2opRWG
llwEX17sMKoumhubLg1JExMpp5QOvTyfbfmh7OZwoAup1NLgVr1VfjFmpOuID5mbGlaAyMElo0py
Qjv9ZvK0ic/x3DwuhUHpD1nqVm+cWmnTM4VDbZ5fhuTAEfPeE1EN1FP1IaAzr5vTeVJxuAOBSMhx
4G5gplvluJ1q2vWp9+VNCkR3/rPimW2PJKuZIFzfOdQ5+3G/4ivdAZcQ1QMdMqV9CWdXJkXz4vMJ
B6j+r557Pps85VQNknNcKi/SnuPIVSO9MXSPA69k1ToCQjXMta+eWpFraDmCUaAnloJKfzKwylAf
jG7ltDAaX0zilvKgdl65E+7SumGa0E6i1Eu7IPggC3PLX7ARHhSCg8b48DYV0cmvo613Ep2IivKR
1yU0i+mfkrC/QJXmwvaCwXA/aJL7YIJzFSjbaAMqoNJt7RUO3Z5gPnB5cjad81yqo/3MLtk+Owsx
4ow4JuqUykVTXejIU3sVYDllPE1yY5Ht8+z4j5Al3M3IAEMWEsw5MRc6D6vv4KNuTCu6O7qpbqb3
bM+ftM3xJX9Atz3SfPUYhAT1+pfxmM0IH8tUOmZ3AbmWL3avxdPfXYEJdoXQYBSlM8QygLEPcQnu
CZ/qk6ZcQL5SHHU4vn+eOih5Cb5vq5si21URXGf+lhYwMOYU6QWOKyYNKwTPK6MOyUdR6OaOybaN
QGAFDbqzbnvjSW4g9374wzyPiCpbZXu0Y3tHYSY4uYXQnmSCl2TzDaNwGTEhAlBdiiOBxZklNvi2
x+i+4QL43e4W1ySb9gZhTU4B2YHG+UwSKcihI7LdKOxPbYOgO++CdWAvVhVna3X2KsRwEufFg9NK
LYGaiBhp1paSeEP91ZXKPYncYtcwuqOi4uc1Sbm0vROU/WjVBYy0MGPjckYLjXeBN29qtlIosJPz
7exN/2GlSVehyf+qlEeQWRbQQNjuUBLFbnO69PLstFOQD0v9dS95+uPChIgOWYKQGnoQMWrdtRR6
wjIKs8Bgkuevyu2mizDUrXx8qRL+/hdo5HtdQFgV3GBIzfboSSa+7sk4NS9b3NLLmiRetrprGAaq
OcB59hW+qsZaYIPH2vAb0JZvMCXA2dsjj7H5QiMSVMYOGUFzplsUX0UlZOgL2XM2uDEEfEnZwsrn
m50CYiyWB+mwFc0Zq1PNLdBPCsrA9PzIwllFRur4Dl3XfMvog0M6xDjxiCwxzI3UUc3EsntcBU3L
v5hQvf/YXRt/i1l7b3t9Gj+ovklvxRSOwlxUj17keITHqwGopQf1urTivsjrNeogzItPn4SXZNxa
l8gCZRjRg/Y0v7vLBgmBYavf85g7+YjUn2OMISLvq0OHPrTxfiHqm8qgc05Ntcn9oeUmEdYxOFH3
6CIgI8JRz5psc0JJrONtd8Efoz0IlFPzzSnZXJdT4nNb3jf5kIfOEHZFopU1WTbcSgaa+z3HDXrL
ZZMaFnByGzYUuTZGoEKpUxBLTocqgBOz9Dlc/RrcrZ0L/t1alFYCBe4QstnahmkL3bs15i14/sLj
yeOpAMqWs387O7LloIuCCXPUJGpeY7PfRqJdRM/jYBWkpgAxneq7nwfmyUhaVkvns6mwGh1/8pNH
Z1JXuTsmXfdiqx9IieTsbuXOh4aCSgv0oiSX96ueyQxBU5wicyS+A0rmdX2NYM6B0H3l4F1HOgUv
1Ybp5Z7ZFb2BwNWB1yYHrjlMlgLFBUg1qw/8+QJEb1OlOFSALks1UG9QnKFG42k0VUSvPvSogYBe
HuFH7+1QkdXfFEln1cNvJdVti56IJyuGr1uGN/M+pQqNd3vd8KoKAA4JKXil0ayHRk0HQwuyl0eI
afiVVNsnwIyzcCtRZ7quEAsn1seqV1t/l6temtvd+ycg5hXwn29eOtpEAdUJ8AOyV+9tBzx7dL3T
7yEQsofGIYMwO4zgti3j14FqhB9ua7Ey3Kqqfa43w6IBat3xco3+sy0wTocPJKcMDnEekZOl4FPV
IbJw4yQVi7M9uUrdFkqS251kJUHcghY83cYwbMhlAsLWgAz/ewgbsBwjniKR2+VT/Kftjy97j9+b
8Ng4TvcU9liFFnM+Nt/wDI2bcRIQ02S2mcWmqB0afK8ShX4ZonHdFa1oXn/FV2Z3lxQzF3jMTJ7P
K94MglWEP2UOG5OlAiFL7WBxN5SrHdeyrUx2KhrKD8y/lHs75cQdojkOoAbzlOsbq4lfpMz7p2dB
Ht8ZF88w26PUaJ9WEjDEOijQqM34uIWs5iKvmaJLLO3m/HDgg0W8ityM08SVGXFrHKt5SpCaZl6D
xc6VXI/ksbP5fBqE6YXuYeXX++VPtihnBfpET6jJH2T2QqPm7iqvCD0LCGWcvALDA/25FZM/itpb
qSXH9B3rUPHPtsOVXLDD2qjIrirR/hOZOkOnjyjBny6IpPQfevhIkZaywzI4Z7Q+71cM1GXRGGU+
IhVnke3rOmnvunWCzXSOOIOH7Ik5PI4XsqDWusXibED5r0msrLOYi2YTrQm9PjzfQ9UDqSShRiVn
uJm8M7lt2e9zMLUxMOd3kLp1s3ANNbh7j50dZy+NVDekKxmcCTRql6z+JcoWW3L0CAHPwOdSnIOC
DD6IPokcCRgzwJBBeywtd6EvVUTDTr+ryB2LX9mz1NW832ed6HcJoIFv/cXXGBeOH/Uc/NQDwF3u
V7mykAE/6bKi8JmPA9nCtYj66GYA+qfIQXd7L6QCIvzdtvogICZSz06XBZhQk5/jiq1yniAIO8u+
hmuTj2TzrbrmpebDfgshBkyiQmR5P8gZl4gMBWWJ/KVfu09KHaRn+1zP6JLnpZnuZwgP/7Mo2UfN
BGCUtr/oIqWlhu4TT/RYvpFc/TdIq/Cgp8HykfMg6qofGBi+kwWrJFnADQ61STjS4V1nryIqDINl
IOsDbKvhlNOfRxkkTkvKOnMmN/Z/2gQlDE0oNOkDIvBAwOXnDiYbWagnkbBPAClLDRJo81+JRyvl
Wr5l/yCfRxBmtlH27+ycHAmTxd9RaNWQRFAxfBHo7cRY6Q+pfLrNRUSGToCtaRtIK/7c7eumZYJ+
kTK4eKAJe3Ej7r1ItEHuhRfkzR7SzrDqiqQzmHTGvINw4b0V1XeIqS9ERnrCyG/STYy5ROB3Kwbl
4k3bqejKM/gwvJCM1q0C6plBWaAka8xfVt4sM0ILBpqozWOvQqsgjTPxeSvwUwco7tjNCumtMiqP
J+q00uVRFhLihz2Zcpna8BE0oPYITvsYJd9sQ8JYaC6HvaMqamylv6+7q+Iau36x9CyW0zkl2cB4
1Jag4OQDh66xKEpLE44/y7ErRO3Ppgypst3Y5KTISb1Y1AsY8zs0sYMSOAeHLggSTzyydJLkQukM
TGhBl6J5V5FLklp4PxiRxVv1cmByWo7iAWpxYvwe5mTvWbY37yPVn3hydxw3J7cDldGSmYGcB7ck
vgwMdUQdJT8JvDJtingvGHg6AcKs9XSu1V3ELGJVK6iQ0NJqxXwC/0boblGNi0RKAhBPEyXA5iBT
n0INNU6oz6zV/HwbELGbLSgeJSEJrumr7vRlDUVAv7IJQWGaM3EiqVdzmBe7dpsFrXdok+TkZmhI
9fmCUNODmDGKQEgyhcj8ggTJIbVuYKGg1uyh/XCcan4QwYmF0izUuNa0gKBvyg4YWBL4tfeGub6y
VmNo643IgUi+jBqr8GiPPk1Oa9itiLazxxqlyDfdoPzc7AXk0jhD+5y7H1YdXRI9w2eJs3rGY2UA
/dMrIVRUsADTpKJMYezs1Ho02sigWlry7lsPbT8Xxb4CbN8rLXwluZTKT1tSRcv7+1Vah5091A9K
733tnVS/8HohHKpkTWTz/VCWxzANU7tda3Cgnh0QA91Ei1kIKPgHFSKJalhY9qf03GywhSiFuT/K
PVp2yNA/UlRYPEeB7c/yDE5QmFH8o1WMOOY6yb8GdPdTRZh9qVQeMwTSyWiOul1SVUxwr7ZYnMdt
6lX3BiF9jQFQj1CkVIbg/bvMBevLYGAhVGb36yJ0m9yZc6nZg6lR0XL8HkfUXIXClxnvMmLpo+QE
Vn4nILayCWi//WyY8BJUtP8cwUbGUQW02IL3Br//CCGEsl81m3HywFNXvmxg24J2zuaGhVgAlck5
GBARU7CAf3+YkmMkI3SiH6rRZM1cqj5Kf0qItZLpqqH10SO/+oZySmeJguHLNReEc5hax/oRw25P
l4xEi/xbTdl8Z+4cLnzA/h6fSHrr9oihTomoeS3YwOLWHhPvHl/Kfpag9E9Kar8mBvdLJxqLLZYr
+92/7O1Qg3sxJDgWoLzolnYyFFdppT9J0gXOo8S5StSOtxI+mLKUecVG7orvvd7n2673R2rITJD+
rTUS8ykdv9EC/JF1tkqEXUxIvWzeUwN4m6Wmr8lAyqgisKEKyPqFS0/YGPeJhOmA6iPAPm/3o/2I
nOINUbNzS25hCwI024qovN9Es+WNOHe+DOQMX1csRtawgE0fe+soEGp2+anoRbvGH5Tg3fpF05V+
gtBxhSw81R0ZKsUYEDTfGH6503gV4yopMGlTzgT09QFR2Em2pUI76oOntfxbdy/ILn6Xya/fViZb
LeO2ySpso2/K0+J4xFJ4Y1UDgVu84aN4/xbEzHl+QqmDMJybD5sJsRgvKQ8FR4VFb3eizLE/y3p2
tNqOhKtsE1drJStaXH0+gKb8n+HR/Pms6V/dNROOF00BC14WU2W/XKlNLpwDltSTtqD2YjQkBm00
WQfHocs2+OijnyHvVfdjVTGs6Pjd4aLIQYkDh/biXTA3ujf4bMWvWA+5Wr9UGUBjunyD7e5Nwh6O
6mhpUnTbKgaeGPBPcr7qcKH/+W+YiGi9nrHso6Y/XjbyoL45pF58xqkZKzdhNt0WOSd6/ZYuiinA
pvjmM7lTste2geRxBu+fjQ4W6MMf+RtdKi93ulya0ZcEOB9YiSC1423oR6myw3/Gev9AtqD+u36W
darout2+dH8O9Ku71O469fLlXcEKgWgZwgSPgvpKiunKJi/kvQbWwF71D6Ta9j1X4yzwAgT8Kq9/
8dMAIcA/DCfoLmkL9ScBBDVzcG55ofnDGcElpD0IHrj3FZxgA3ccf4bDgO4KY1T/pfHxR3wYkJq2
EU0wECBka4Yp3Kol59pglUVPwftmYDRti69FnWD4dXiS1H0dZvNZfrhRJKSewN8FwKL+h2+rX0MQ
qYi7XcUb1eJGod8QjSLzIhwFfakIORE3QpqOIDMg1k+ewrn52P0887/fEVFx9V+U6OSwiOzwksHJ
xdHJJ18HgSBCjTQn4NUwxhM+cdovCnLjPbQMfx3YyhZeW5zWQAQUTXs8RZmWSWEZ6jo+nv90eGw7
aMYJDBY0rts1616V+5vAXz+GZs1cDc0+Y1H/hBoOY2dtxGWhc0Ttj7IJ939tnD51ygHL9mtfBYS9
S1KiehkjMaiH4qT9NtbSjjDM/Q/qG8VwlVT59X2/GBYwOGP8L3nMn2mJ3AxC74bWKEB9/yqySTYW
AD7ep40w6oQYPqaBGPyaf/RjOwuqcvqPfLtNhi8qeXWDiFoUUNR2+UNSzx90jA/X6PzzMZga5zAC
i7Lnrl7QoSYJpouLSYrpE5tSK2OLbV7td8aQVZi9pyhGpZbii7+OJrC3H5AkZb6t7wYIV41ni8eH
S/L39j9K2+YOzrdueHi/JxTTRQSYXFU9dN/dssoEAPzdBetz60Q2vY1sLW7dzJg2a68Y8ab0N5cW
fKZBnuts7A45IfMGf88AHmqo3zqczEEkHNdvFs0pxSFUCZwzzNXV9aHTyUjIr/SdRqC/wSZ/Hx91
USS0+hKfpdeZrQZHP1wZF8Gvr+ZkHpN0gb2jc1JJGDev8Ft4EDFvghKaX2fyteOd/WfPu2mP427V
8DU2ZXVJjbJWjI0mFKHguMQR9tyP7v51p7NjlL6Y+0TsTlGYmCdNS8gB8R4fZsslTF2ZGKXRDgtb
2ONsx4rrVvSHAxSBNQ1L/fgBImbtehjmDszx6TXnsTcb/MwNqNygarRdqEkh3Ubmixspp6cqMiMj
SnwrhK0h1zzzGRZ8gk348CgLBvsrgay8vs6epdJR/yIZuyogUw4eXCo+ZKBuTrRx9SadHMsDkSgm
iTRFWl1HmLG/U53gUEiZTH0ICGuaOBwr127istfVTVFG2ETey62nGfqDpBVJt0eiF1uLIvow1URR
6TRNjB/OT8TIuhEFgorhPqBPYqjmKVkk1HiuDc2S479KHpoTYI8bC9+G5z8xcKpvtmTlmKPqcvvx
4SsOjCmjnBFIkXutGnz1QRLEkViQsZD7qYqs2GgVba1xRQDpOMN7QhvlnhrNWtvV2MiTPS7kdVoA
2Go4aOKuHzpEqBdVG2gmaUtmqX3CG18mtrJzKi//d5Di/bWduNOPWIFjSl0vsGjv1o9A8VVskd75
Q41XzdS7b/sFezTtc/atYn7D3Zh77cWvSyRk3bk40/pj12YRcJ1KjxDdHg65TpipwyOM6Gr0LcRl
o1V8KDZMbKooZh8vGDSgKYbhuap5qDDN90h8e4Et/f/yKUYTGW/HpWohmlrA71D9ssnN012znFyI
bDtrv7UQ/wgVTVeBA0pv1O9P0/VsAxSIqZ7GOzbB61AXnr9IpXOndF3c3JihAZM+FBuqvBMt5Kc7
Y+KQh3OY94q6iHL3nH2ffFw0MYLviEp9Xd0Bhvl2ouXO9XWa9DVBs4VgwSk7WSmazPYv0vA+Ba4O
iF1beL6s+8eT7Ny5rYeC9iSQBOlAEh+nA1/Kd1U94bnwYz77CzrwQ0iYjgt1H93nyyA3pgaPfTPS
JkDuM2uxQVoLK8ymdZazo00C3POT1WWdR6fmq1E/G3Gm9BRezt3Sbmyov9se24IQc5YXSdP6QIoX
qH2dXXkkjchvflfX1zBpIr7auh8LE463D4oC7Zcpd1gDoIXk0HAxM+/0fSRBfnexhWqqPbde42K7
0MP4tPdjDagTfTOTYbsX29Fsh3jFNEUy1x8vWmLsbTtT4WA+oIfVVc4OX6RoX6ClTzHOK1VX8Qd2
wOGAKPxNMV9fGawZkkvPq8JmMG3FuKgBsEpeptBezKWIl6SDxdLAk5aeVBTUCPMe6NzWzOAhot1h
QxQm6agGxSCpBvarom/iOT1IT8b8Ix/QS36siFlKwC0KUt1xILr77REfu2t20WNwrzg7TCUgp8vI
MNXUItKiJo8GNbghODVfXj8e/D69Q+jC7H88K0EZxWyN8091sbKJgjO2IJ93DRMnjteTZ6XyZe6t
oWyNlLtS9PzPQ7aJ4jD4rZM5Qkt6YR4HtcJ4xTdSWXnCLN8pEIbLbRH6ddxrvrPWdqU1PZ14eLCq
TTMC7tE0s/4q9ClHjfTWNYEVs4Bh/hVGhhU6DA+UgudMF//IUGQ2u6Zv1haUVxN9oQzHa5pIYdXP
1reqBlyvfDHmnO0MoMnK0MJui+tjHFzv0qCYR1GjsAR4Nw+2aBag78W+FRPLnC4zJpXTrfeOPw4A
EDn2nZlaQj3CeWIMCp5djBB5mhK0zbh+3EOQz7Q2omLatD4I6AMcOuObirSRqJTf0NZWMbcU27pf
kVQ8xwsGUJElMPV/LHUciYOYJlmdcJgaDDJSclvD7KQ6lYigE+tFUALQnybRIUwu38QKW0AwEb0R
X6UCNoDhuF5Lace+o8wotsus6I0ZX2mnxzIZb7wPUxvMB7AK9qbpfe5z4JjNESnC9Vq8LNPIYgXE
KSlXNFsuXUgPXq4g4T+5O6zPfDiJ0v813mxD0UR+Al731+y736nPBNsjlsImTyoKayELUKJAI1vv
EYZVf+dqzR4kmRGoEPqXC6zMJqyQunzlHswKUY0wa4qtiOo9Zvk6/JNCttQ1IpgHW6HR9IiK6ziS
D7f+yaXKhYCT2B1mI9yS74dIJ84PENEBcMKsykOASwR6Tqd2k5ldd+y2yM9I2u/wlCUe1yMzpYAM
8LBdw649RTf7DST8ncbrjxZ2e/ZxTRCt6+ELYS8zhkFD7ly2Y+3+WqH6YPvQ85YiX4zvzRUcSspp
3wrbVjUWwFc6x8Z+HfGsY/ql62ajg4c7KiwAO8njbdzD28Q3QQtJ3KbjezZjWSUguCtGuFzKn6CE
5+YKxk5DgpcGAEjTzI09Yalv9LbcSdO3H7dwxUDgHaDS0kSsSFpH7WxV76drlpkqglx/J3MEhtbX
Xoq0gRgoIRmywkl+9ilLBSYYvsOzr8tBkGGafVgegpvz5Q4edOPFmadWNoM8+F9oAv9mI+R3K4JS
P2jy3Sz8K+Y416I+jiCK6xYIxhSbLaIDuYviguru+31xHKhZF/orYukoDO0VJROu2YvrqjFrAUF+
f75TQVkxTs62hcBx1m0LICePzoJfX+cWYSvMPeWCxPUlG1MrwnMNUeuKz87wTie6iCObaJNE+zhk
9Z2Yz7M/vrTNKIYPYaH5bB9ealSJWhoKhY6XIXHXMqY4TlhO8JIpXztIiwCQ1OTyvlr7bqm7XX9T
xYvgb2W2Ia3DB7t2SWJPORdZBbCGIZK+xzqah9sbBj2ZWfPIpUKOYeIPyf8Y6ZNXodcLGuUAzOC5
nmR4yTWILem1nIiaCS3JdAT7ODqz5KbQOTeR6sVDJvtWszLyhaJPMJ0AXU5+dTEix3XWHZyPy9l9
HVKv7wDNZdykXt0j7qlHpOzy6K4M5MubOaHx5dKvIM+MkUTbxzuwheiRIdjMaGzqToJinaEDgweq
eiJj4orhiy2ued1+u6mkhl9zUuCrZ6Mcrn+WjYnTS+q495cs1zw7FC6uFU3AvpDhewMr8tom6X7K
wKf9qDP/DyKWV50avSIA/jvw5e65okrrX6YcwdJTCXFo9rAQEl28grIqyWPZsMyh1iF5Y1phxexH
271RZCtYneNeNoCv6ZA6ehh2RTGG+xA7MiwWS14QuPd4gAPcKrcZB5bvtiZuxVHzKmE41cCvSBu1
VBq5SLro9U8WJmjC4yV/HyZNV1EucP5DTtlSCscWzkE/udIKVX2TtqgCflbC1SaeQZ5TEE/OZ3oV
P5TbqtvTyrs4PrYJdPfk/xb1QnzTgx9JpFZA3oYo2ZciR30US5/OkUZKMeGoW5uqFazDRT54bE0f
n2fBzV66pE/91g8bfRl0HJxqqSxkQ7TRnRW/OyVOI6XwlqTNkYPx5+Fe/x/KD0Qr+t0ikfw2reYL
l7Z++iU0KsN5tuii0Htja1JDLyzyqs5WE/+IZorFsWP4mx17ZVwzOwqjZ0skz47MTJuW3elS0gNi
YsLqJTuMl4Z+zHLSSBvB4tlvjoUyRgCP814E9d1OI6G1iy9qrIsWGm+Wh5AalJl3zrRwZyUSClhs
01coOd13HOcX095mURnFI8o8b+8E2C6r/JqzTfbLHRBR8Dl2SGZCUahsaIHBeBxHEAz/Pm2cOnk8
6x7TjAu1shjBNpwor6rGx6RGsh3LR3hpL8XZEp7r6JjZcjHy6xoi5D7vq/mF/stSr0s/FJRZqoNP
yHuucEszAJPxXyKx1icUG56h0J+ZJkD80tc9BeKmLHBSyim380EmIpyHPYg6E71ROgHlji6sdWWs
xYJrXR1lmvPyGWbvtO61S+GkGTv+YVLMuk3k6PzBQQW4kmduvkXLN9PQRc8UhQX7kjWhsHyfWq4f
HPDnF/WNmg1shHFGvIRdbNgVT5zdZmemwvPlHp8UkCS8kZICn9FMeptOlixl1FxWZEgifU+bxfYR
8oRDj3ERoshPkutVLSWtNcOoyqISKgfADHKFt4XOhDxtS8dyjk9XXBTMkbuy5MSjda7bBnkrAtHg
UFl0Yo+f8kXEFVPLV9RNIHS37meaDuoprqrjQWjroKa1ooH0vzLAgzVFCda1JkZJo4exX2CcFT1n
BWKDUWy4oGCF1LUfMnREH6A570hmgvXGTOgVY8e9rMHQltuttx0sB11TweFoVYcsYOpiPibmYX2F
r3hQLbJt6SzlemmqB/OiRIwCiyrN82FDjKfnPkxKDVDxrKONU2SQzGwhKbkXTuRDqQyEX3rWeIgs
fvlfAv8n5KjrSPrRzGFyOvxTjDYpb8Tn13+lcK82Xx3HmFAzOHrGmxw142SnAQ6KUIDEqt2kY68O
lN+WBm+TrawTYUDF12pmQmnygDGOSp5cTKtvK+3c23v+M4yBlvX9xbkGrLJgaypQ/iAg8tjjOZtZ
YgLGVhjhW1Q5GbcWuVRJlaxbxcpMbwQHmZDyWF024jvNJOoO1lzfL7Bw44lrseSgn5bxVqcBpVGC
3c2d10nhl6d6mc3xIQN3uQdd4yuhZtuZLA1Ew+13H2+syboSSE8pV0LUm323xUc57LzGtVBIhN6f
diOIOpFTPmkTbZ98siV26aqqidAkmDPWCgYvF0MsOa2FATQu/vH53MqO4pBXxPFSn3JxROhB6ho4
EcN3yOiA9jKAGM/6e4KAH4Dqixj3C9Bqo0bQRWU2N5VwxolCS/r6dSEOCTJN/XyO0zZnvdhcdy8e
ZAbYJoR5ujSnMfwdA5A2hOwXraNElP23lrPCUJYV5r8ROjqa8p/1h4+WGDlw4B2DcL/loGuC8k7v
m3z9u2YyT9uNDoGFUSde8kh11sy5JENp3ISHlFoRmeaN8io7hAUw4S35NGv8+02xvurYC6moQKbf
ZOpBqC3VPlblezrZuTaX75jQpOtzvHT+x7AcSCuS2sA2OAMtI2p1Dmr57wYbDpiT162mx/VTRkxn
/qaH1bahbvHalPdoLWwTYNEOCpMxJbFt02Y7/YFp6a8bedPj9vdQnepUMzunqkukLQavTpg+BYFf
a8QXt106o0d8llB3fVsxmP9EH6T8IK6bIUq+ZRl4PshfTZVTGVy37n6155PHxiG784RDg6O4/6gO
XeoPJCXSWLxRe/ghH/ctGiEex2hH1yVV5QAVF2Zz9g0GT2An55AGzMYQYfUMVjKTItMBWdu9dwwQ
OCapQ9a3o6STtX2b1wwUoW3978bkdJo2shNIkBb6wrSRbXuxEQsZXFS7cqPN7OSnecLYNaL1SNzx
m5AfYwWH3jNGAj3p+c1aWWhW7D/JfgMS40NkSBF3kisV4pUK53oq70nzbOUAbHyAF2LTBraYZfyR
jHhva1aiUB8qNTVgctEbX7rlRWMAvYlYcqUKy1rdw8OU052C2xAMz5VL3XrNklPTsw6UNAMenTcd
l/vJMzI9a4txc1YueQjqIoMOnch30m/a/B9EpTF/yAnk69IEtW01YoxBlnfAZk5hWtSqtO4m7E3U
dpzQDIUKCGZ+R1OAuJq8f9pY4WiKjJwbyvhLgYTlK5zNhYhWDQVP1nu3cAwJhdD01dmeAuHJ7Lfd
81y1xm8E4+urpViDMnAGwpit2eXkJdWLaIlWvJYpzWFGQOsIMlO1ahRariz/NnSqJY/la1GfnwZE
k4HfCTM2Co21mdKu7tSE9+0HaLHSZTTpWJAryFR0CEuL+PLFGBuLKdzuphb5RCqAkC4bvBE0g6Cg
PdURU+4wNC5MBduMph3TIc+D3b4c6yH45+lce+5dX32lVfXnYbjTHsXtOZWINnwxouCtaMVCgx08
vy4Gv/ezlJdjBjfUlgxLt+0fxVtqBj7V2+n6mTJgRsT+3G1IfYaah2dmYSB4660Kk/2hDuwQckYa
hlUzmTlLUEXgF3evqhq9jrt2Q6YSphs0OpCI4yhfne7sS8M0+qGS3Gi11XzM8a90z5/LATLa+uw6
na/kWsxqZMCLGvw5P2LTlyG7i1bW99fvM1AOgvsu/D8k5mZuXvacpxoNDLTPkPxUSWMwmpPCgzkW
tymiwGm7HXeLqxfQxIriiqX/B9SbD02quveatNvNzcrTidbI7XmTTmY/mscShcs7RFWco7VZxWxN
Iv+AI2cghlVKt3ALEL0IbtSEI3Mpzk3wW5e8NGKaVOOASwoDrDDVYxsuKYoJUEQo7zgbKQXNk1xt
4MmPD6nTDTVHYSHkVOJlj6LfAhEobokcFNXzGPM0H0ruNJ0D8uUjJrDFpKBFtGhiYKrr482X9M9V
suQfVTnddil66G33PoOFKEhqn2CJg6HfZvBLv6+e1RYuzJT2fngAFga5lP/z+87O5NReLlBQAoK8
YUehVhuRl0OBh7SNoDz5yBMQx/3Q2oSagwdHiqySwWdxOHlmI+74CkPDEgU2/OCvqoTxGAk9KUKZ
d7H1ZIcQ9w0tQScnguuKVmUlghE0oLQR9u/RG1W5Wt6YC//R+IZKgz/7UiFJvIOdganxik4hpkzw
GjlRsCD1UW8KEq7DYwoGBKHn+/d6woi+VPW6H40DtWlrfl1uiHq2bYsHAxWewqr14KKclhq5BDjS
Wugzk4Sh4McjYzqcvmUqTi3Yt0kglYsPlceL+YrwJV4HzqG7dh1PNbGwfaquRj+y2lYkgdeT+ZS6
e4nY1DsOywq0lu7tMtKun7DSl54yRC9oiukqbvH2xFaOwLUhlWPHYN4jBLU4OGj2pEpGSrHYe9sD
Bwp/SGYwmC6Tj74cYG5SqMqxYjM4t9dySOyHfQvkZpvDjl/1FDMTAnyrFt328rEGmG+bo6LY+Drw
clp8SBA/TjlYgyd1ly/H+HZEKkKaOy+zCSby3+p16vg+mcKgl1CyZd9uIZaH3lPp2r5Zkl6Wqd7i
DD4x8nyaif2T0FxwpU1V6iKlVsyEUEHwHM+mrTDQvyIlQchP8YOAgj2uR0Md68WwJPdmEGDAdK20
NpcWVtB4X9Xq8rJ5rkrnzzT7GHm7Q9CoH5YVRJQTrFFo6D1dhDsDIRaata1ih9rRm3iczfAeZVIw
Uj1ozukXGI3ogOCEh35ehAqsFnIEsF+8XsPLKbrlSiUxBzkxEYqebVge5Ddcc2zpuaviJpbMgnMh
9hJRPKlN5Nfw8lsCGk29UFoDieH1+d0T46sqJVFM2WWMu0SFR7yUv45IiuSEWPXUEIwAA2ub1yQu
HXQBvbPxUPcstK0USnVYgyDDl/hJYMcff9zaxT39M0fu+DcFMWXmMA86twHfapuhbPsHns4xUE1W
nB/AkVpsoSXC/MLb5I4HND431hHf4Qqg4nBR4iNXLtQt8l5I41DLSJhFdoWVsaTV2xeKILlrzXNB
3I4K4JZpXy0Mx72d+ls3QzvlnulEYR84uYc0spoX0gqo2ChSTwzM9PbMPNtIOZ4NIyjvyGnXqMj4
Ku+WhP5EyAj/33NhKfSUgAnnG7qdCl301tmPfkdZvh4tRtBInzPUFlDR+oh1PXsNhjWynAVRVN/r
pvtJD53joSZwaWnAuT+2pbAeITI4l1Oue9JIAXw7u7MH3ZGaY0TMrYvXXzwNcft6yT+V5djASfxl
oax525RgyYAfxjNSPe3ws/V/eagIueUKza94AUNjyBknj8yORtX41ObvMGE5Urb53UxnXxYtCO/s
KwH3xwj6HTSrDzvwpVKFw5/QeuIKdqR1xgqCcKPi1Sg9vDASk53lgMulszsEFcwSp58MPPLVVLTx
lYWhE7gM2QuvDmdiXYD4mYysh6cZKRLxxRNGdthTli0M1bG/cNGgRmSjsHzVy4oVX2t/BpxlE8hy
1DfJhL1YB7+9rHWiLC09dNghaQLvZR/ZvvJ/R8wbnJrRyWtWO70pkrS9hmQMzyTq/s1L5dWavFnI
coi4fEZL/pWIVjzisE0xfpMroNCyB7ob4B+HRwV8e9XoDtxA9TWGK3DiAu/1gef9FZ45Ulq2yoiH
CqOB1xyL47LSVZIrT6IHhvWg2eQyIH581RCNODNiY7a75sNkeQeVb8/G4A0BVeQ4LYSavRdHDtZH
QzrNbM0DlmVcECJGrI2TFoRG4L92BUnJxHT1Lhr0AqE0OZndfDhetcbC3ZfQSE5QecYI2Ux/H7B9
9FEmWrU+IShHnyyaLjkEVWEDgKYA5KMtMjlWXUAA+J1QLdxucRyOudp3lCkXcGd3ZucngW7RP/Sh
OccSNgoIW8WkZebh21pNe2/k8J1eCB4tiaG8U9QonY1D1pi5/0cB+0RUjftd6r1/mfq7mr8eFfwH
zG5WHdazjU4KSEwvdqE2LwCEMiCLDG3vDfjGqOmGIc0cYTVpSzWIHprsVwhtCikThP/Pag8nWh+E
99qe/zlnhnBC07BSRCDurPmPO23PjcVAnL+2KwtHNQUB+o0lBkMeiwDIBFhgMukq+hPMAbTwN1f/
zdVz7o3qKqtlY+4BvkVnKosnLztm/TK7rF9vxTqaoYaObYJ+mtp5ADdi0czudxaCSjIm+IpgDf3z
sp3yAX3zfDs1zBSz/PJrqrKf5my6m4crqQ6bV2Vfk8YRQz/8G67bz2QUu8hSlUZPk32XjwDBbLx5
wd6rSiKARFAApc//fBu48MP+ecV4bNNLoYVtFYZB+3ugStBlXU+jkXVYfotLIWbQxWmxx9MnhxiS
wkCk/gjgGAkX9h/lmFMwysH1V61KLxb5naXpRRTb55tUaz2fyq/xfbCvRfv2u+qiUHsdn7k39i1/
BbHGCxIb+l73UAx16T3Y9vcKQcZwYFGRs3/BWqrNFPHyt1bcVxFaGOq+IeiSqjkSPUq5A9GE+oyq
1gjYTBeSszJgftH+Nh14m9VMVJ0MupfR0PHpjVIR94dSaAODFCaPRDvPnj8Gbuqu+FiRuewIxJf2
DhmCWAKOyXdDKqhMC122WHVC+xLf/ud/83lnpg7IgOIKql0uCAYhHH+MJxaTLiaJC/7C4cwHBKeA
QNsmSP9fj46qqLfsaym7BSYgq4mQMsj9xLYhhjSm+//nJg8Yzjzs9XRwDIfToJuf6M2l1vg2++bE
vXGZzIMoFscBtbSAwY0DTtKr75sKzqaTIdpruQpIAN8PzSZ2JGW8GlzOjyK5lada2YZhfHNM7Bsv
6QZRks/ZeJv24bWoX1DM1tDB2tGuGPcdBMy6EYR83CZ65H6EEnKWCOMPp0xKL59lKdelU4GHEZSp
ZbsegjseX1n9SKN9hGIH25umdgLTUbujvc+o+Wk7X0pkGnxdq8/rRU7AC21wJK1Ktmow32cRWqMy
g46k2PIvpP7SNYFMnpmOLgMf4IvZFsnlSbW1sQjMHC5D2oDoGG0ZVUzMz3ULAoA+RlfDRzWqn3Ia
qW9/BhU8pg8bQ6PQi9WYRfu/RNpZAb14eWU/8iR2XVsNV7JEX0LrMjeg9nO9eOVBzYFwY0OSAzf6
exuK6Fvd5/2lb4QsVJCYe6NBRDBLCIT7CQmkhEow3Taj7QdrDDjqhhKYoRuEa/xtuE6rlbok3hR9
hbMq5ttiX22D1s2A2lpDgsEQoLvrcGkApuymoqQCeOET6mlrg+FwkNBrp4yGBUJKnCfzxfRIFSw1
6C+L8bo2BNMz0YnZquxEuAcpVWCwtnuAWWhq4S6ywlJrT1E6mpmxJvCHvLe4Y37eWcx9Njkg4nYg
QQCzqImAHaKKONSzGH9Vct4VYUJCP0wvpW9/jXdxg5i1UfgiVNCmsxvlZAqTkS3Mk8TiRTNjdnSN
vfUQ/rtfGFUFCchwXgcRGD3Uj2NXBErV+aNRkxyU8t3XLJRY+4OAD4+StwEALElumkIPtCYzvVMd
iq3vbaWb40wp8y4lCYA/QTRy1F94D7SBXpf0FP4AqO8pgeNfqUU8kNawJdwofk6JwLk4lrJFLpUz
8ujIVILelWezc5nwCxcl30MYAQIM9Vp5eai+3d+Rr7fcTeZTkD/y+ycghxMPFjPn1Nkihz/1H1NF
r6dM6A4f+UoFCV219CZAnZ1YKMDOT9kXR4LfsWLbBSbihrvcfbvdjVHpcSsAMOmIOkjkCFYjXp71
SqLWg5OS0YsTXHcHvGjTybmXv2ht/+EX1k06/DS0YMlUo/MVmSbgVh+Emf3UI8Q3m59+qPiAuqj2
UFjOWCLcauoE10g4u6w+HrMFKzUSlhKjm9/Ax6kXnV9wp4r0Tkv83+JVU8azlLkBYFr8B80bxblP
iFrn9pBqMu+ay/sxjVqFKIXf3GPx1B1p7iZ0jYm9RuEpjbOBhPEiJiCx7eA1V1l5hY0sgdtRv31S
bSyPQsCpW7YyGlYg+xgp0kKa1bWBeBUoo0K8mp6nwyAxWnCTOnTzQxemqLHQXkr8TZhfwZT9tn7V
tfJBpIDwhMEZHLrZ+klxsjMZApkrleW0Fi3dQia14AvMSPQV56Q2o1MMrpW1hK+3xMVsBeDAyXmo
Oui/9tISMI0MxKt3xhWivEmIhMW0jHwml9l2AnsTjTK3rZJVFsZ7DVtrImMEj4HQjui6/VAJSlUs
1BE2mhmJMxgfv1RiDXXOsoqSoBkD1pElcYwh8fQezHPJ5++5xfYLrgK49SPPNgD0w2ywU4DX5pes
FdsDg+/3U+Dcza5VzyqDRK8HFL3X812VveqAo18DrgQpQc5f3PrF0g6au0MYetBDXIvdjc9zgD4i
59sdDm0+RWbclyGRR28h3p1tMw/MA0MY6UDv5BLrn4H6K8g6tUScFkM3rWOSpvcVam1VA4i45yz+
mX42pZjDFWzz7sMHCAmjlmGJmpIzfV7FkhrOzSPW4pxSBduioqkyHr7OynP+Gt9N+sv0y3GOnl6x
O+T1ifEWT0iCVV/NH5qWZcIBG1SFjHavwrflpvIYn3n9dantdNfKqKnkwicYxTACeR8qR7kwqcKd
NrYVYyVv9xsRkVZUpNhNkzcG+0DGUr/F38vZ4vuQV+k+1I62mp8WExOBmihkqHSVR8doCu1y1q3O
foZUl+rdb1vGfwGEuEWqb1b1YtCES9PXC5EXrbsq5XDLEx8wB6PTzxp4HiTp1yN7pnwltPqLGYlv
eQ/TbLBuW0WBAGtKi8JpouIgTdlVp57CpcFiP++VAbGgvzCaoSgL9NzEWYKqBrwaX7GiYEM6B9pA
tNQkrhkw1ltlFKSJUggaCdmQkgQw3jkPIN0qBQHmHxn+u8i+Yjro7Pd+OO8xCWnb8M5JQu3w6uKT
TvwQZYrU7Esf3Ir6BmTHLn0VenHa6sL4iRftVJiru2LgdXAN5awDF84/TQ/1q8HqBqE2qKjExELX
QI/Ne8XtZgkyjengiIty8MfFnwPuhdXBoOwIpnbs6836uYDN6W7XS7MADEyKUGuQTLE+zVeEVDsG
NunEiuY4CZFcdyZCQrXVXpCM9My5rf8GgOkm2zvBU8eWHCpP2t2KdTOmHVvG0f64C4Kc9NJZaAcN
WCXiZ4vAOLsUzhsNhzVydMCPRdcn534sjSDurIrockZA2WVyRTNTmXOixUd4D93MLFHv9T839w1S
oWgvVfELwo2tuuqUQRn+VGd9EXUqQpOQeBuZz7bN4Q/SH7UidmIW+I4Q170+HO3zdGoFYzQr+rSY
78gfte9fgjR1jtF2ieil9hxT+H8CEyNCIeqr1Fb0RWtgP6NNZYIBAmtqNOWLHWuvovsfNriRhK+4
uEjxBrK168x214YmSSRs5jDBRL7uXAMyjaI4VfxOcr/az7LbN337HsEH8xO1AQOMTr01B89sST9/
mJJjvVtIZ1Vjozswb6JiESilCBcxWqrsAW9e2v0c+K+RPxSXLRCVJk/b559bm2XosX0ytjmiAplk
02AH7Vj1OEHVL3JSWr32345J40zx2htkxNYX+BwafJK3qfUI+R1fkhDlb4h47b79wOUBeofL8Rir
DaLO/sUFwG0qkmRM+GqB6x9hL2lkeE3Tp2jOFA9kIwsXWKCgTfRapZhERcEd9q1D/qqrsCkidB0O
g/jTZeiZtoTlB66Vnp8vZ/cklIoHfCq+J+xQgLBj0VK2kQWNhRWSPQU6ZnIdIm+KIVnP8UCuelUw
YLngrZBOsrE43THsktZwn3yxkIf8q6F551gH+S+/O8kfk5iwrfO86OQCtlRDuBuextzQ1jRGvQwj
w/O4ViJ0+xsUrgOSJOVP/mKOU6IR6tJPslj2nJaBFTAdHk+Uno5vaOWkiwT4nlZwlfbCB9S1VXxx
O6yXCqRu4hPiQdH8ulu3PIvwIaJFHAnPdVgmaVQMrp70xeF65mBfsBOxVvfIkcsuFc8IJSS9aBt7
7I2bp86RX2Vp/Ike9aDYsqrDU8MZz3uDjd0dJ5iQx9FGex22G0Pow1Ky3GPEf15ZhFPpzy9QLYbG
oLu+UA4lIHzqRxUoElp3b6QRYyKyYyvOrEExh6lw+kQZqbw6jdB3P2wFHEMGvAKhpYA1NPKAOrT6
8H0fanWJ2EwuOPoocVDzDIxmaGQEqrUUBrEUvxSvdXZeg1da+i4TryoKO4tEuUxW8p+V9vcSRJzy
j9P0beglSfCtk8BUP/qWbHFtE6MQMC/KFceol1btA/q2RfY86ZsMXt8ZxPB+25lx7b1VGHQbunF8
m009y7tCV1WuMsgN869Xwtu1Hb7xO1Uf9A92vuXEK0QcobfSBZfq9n09M5RT5PB1+GUpcVQZN0Fw
BLdBIHu+dhpH+AUgyhg9pHMS6x29P2SypRDKPTbuDrtYBLvkDI7clUhBwhZLJ9uACuiubeHgJJl6
3DA8DrQRdMtaI7h7bvE1jr4GzcrnDEluGlaGru5TmFbOjNXMpeURxUbDF9KSIp1NQpqSWDZ7ibwD
8enx7H4v0UzZI9Sj2XC7t1g4VQ8na2gzESSL0GCjEVBLE6jagoPDTA/X+n6iU33kSn9as7msHq6X
8ZPCwWDFkBWtiLv3z8yLvdnhZYyAJvJPJ0Owqqoiv/ht6+sDPFbvywhlq8tqZN49deO74k0SZRZb
5jTiutEeeSpAq/lxuvZiAYXA4DRRtJbHl3nJQdXAFI7VEyNk0N2stPAjQHH/8bHm1NQQGmPeaOW/
pzRDN/WBYGI0BY6kpoUVW+K6nto3qosyviRNpeg8j6dRhxKFb+RMFiUdzBCdBCJm9yd3K1bRAOfS
UyA5CgXZuvbOG7We3Q/GmEn9GclQB4LdkcgCTUt7Bu/UFG66THS8P2lix0M0BHy4ij+dhfbq6FvR
36feviUzLRAimN4fbc4bebHnOCztGt+pRr4RDTjP1qvFn7aRnZckJdKXfMzZOH512XJS9dKdzySg
93HJ5PzDSJi8USOkkY8b8nOfdyioFN1/AxSlPCVJO4aReyLGIj7L78+FGs/4/P1wQN+WwtzdvLH+
fGsRKxBPgsDwh61W2g1zEYWQFVr8FD6vaLEwHXAzVsb/ayPuOHDFVCTfqfm3v4cX1DYp2ydIozQM
+m0IjyWHAlMImRxWZvaMl2cVxdqBB/wZaBIoY+RE1IpVbnd0mEiNmjxAK+wuI2GhahLVAXD71QK9
ZWSrGzenKHX73IuOwH8wkSxmnIIrA55pHD3ZPoPBGoiL1iLj6xUzee+My87VINYMoCx//KgX3GgU
Q/aNWLJSMnwLQ+E+zmumFCzfeP+3h8XGSjWqpbR3TfYPaCwNFX5XPuw1FQwouhOpxuiGpooQHbj7
EzePiasN9PipelLFCwLaUfKwiE3Y14glqSdz+j07NvBNgR7tKDL+goz+nWJzKbExzeXZcosHYdpQ
9GjudXnjF08cUn1vf2kkW05xjgl5nDL7xeORDKtVqd2PnEeBJ1R1drN1zTynFkNbjB6ltjWeMaEU
pwJbSZc89WL81lbjdAF6pXN8MErrK1MiFEySI0K/kwnnmjQC+MMxESdocKZVIt5IXTzynxnSDOFt
Ijs5yIfNHlArRitIAsNRsirJpcpu7QWqwx2vUCAwOOTUXBY6e1cqKYS1wiLxAXHumkis7g/DlgQ6
kkzMcBjhKe8RwViV3bWiinzIYNN+Fo7bfjFkXXicwIip8EQ5zS1IrUtBFHvwaagkq3pEpCxYUvtH
WyMyAagQpSJ2K16Bvj9yPySH5dRU8njN+3McvmB4XNkZ+UEDXWXHAADQ7LPNZyHbzRhBQlc7sQuj
jmd/7568SuY9ddyxORTfIskgBNr3mUfHz37xMbpUQhFouUtFxpUGtq57SC1fay7H3XV0E3WFNPZ1
h8A1RlOh8h5YyFFzrqbIGH9L1GlsTqzc9onrr99Pkea9+5bMKDZEyP8VBP0QGHmZcGC26Cve5Gj/
6VRabHqH1gXeF+7FJzmJRMuBoNtoEzSMb4C1fxcz9mCXHmTuRdtf8o+Be+5DM0uLCNS3V54eeO/m
mkV5F5gS2bm6IYjC8iYzgnf/KZxjypmhPxnG5/F9BlptwJAwU54MLF8qtydEkgbhr/uo0vCi4N9Y
i9Dil70+dnt7aQvPWcNqBe0clm3UIiHXCdKBeBzJo0B2c00kJOPVtYpijQaxhLwnwegMvfPU2H10
oheIvXtfB8qfwbE+4dFSodYeHUbSD/Aeo+YdoyUXoTWfkvXw16Ma+dY5T/MLN15zk/emTM8/laju
651KaxrvGyzVD3lsl08XcFCLYEj+v6k/2b6qRakl6R7FJ4fFTVV/oPBak4GEpnvagHSyBml3/YFu
vO3TaevhdsfyuhXcn0OUsIbQu0CfcHO5a/J0irxw9MiydbAJD5sHf+e8GNOUHSXeNjvlx2mf958j
ov1QyL7Unw4UJYNc5JbBYA21XhlBstmfMXP9kjX6jJjEMyz3jWgtfcgFAzFNm3hBPtePpjuWU+7w
+zUBVhRhjTvaezqC1STFxjDi8TNI3BvQaA6Tj6K0ejwGQQ8mFa+1TbWp0ezgiRCSIwM3a6r7ghB+
ehq5YF9kivWwq/pUoJl+1QKiBsRwGfB/RR1pDC/c6FTJhbpB+rlwhJPt6Fo/xKhfGTlhWp+1jwau
Huu3jST5++LO4VY2lD3v4unJ1DlrZ7TGHy37BmX5RAFTsnqlKUHbOPXN6ibN6jceGbAEAMRWBmd4
ptGeADtzNxYeG5zoCSl0/K0ItfBrTN2eC8vDXDV0aaunoqhgualxFKvAEtgaG0SftmtHXz9BNROf
vX4FQnBoaWgrweD7fjZyMqyO7PUjKsweeNJoA+vZK0FR/MlRZ5ofv40YFMb6RIbJJXrv0lKlPDp1
9WcNjzuuSdyAZZgUEYvHURyH2eRP3TMwfOGCqAG3H33C11CzX1ZNLH6M+wqwF+9CJGDW2pTwMfiq
ppxvxNmRwClngdOyKZATAiJhuEYbJjoynkrs2opIv9jwoKzd/FkPOkzjpa0yuAUudRk1m+3OrgJI
nNESg2McdB48Ok1rB6hVEIzHwP6uAWytXJLsQ4msk9K1+RM2I7x2wBVLEbqjxS6M0HkiFPMmLeMP
h2BqWjZ8anCzapcVHVvJDs4YNexExbbjZrnfYe+jZcbsqjR4/6/z1EG69z/HwUhLj4hlg7DTz2C3
J5mvGGT9TW3sHwgV2lw+Sp8sLAx3oacteVnaors9iUyCOJzlKUaJX1/crL1O6TNsMuinPeQ6CpFD
THoIJEsBi2h46Gd2OYJgW9cs93gJXm9E2v7xpFXMzrfviHRKpKLxl2T+eeojtI74jJPFNL8KnaqJ
oQ6btmOz9hOz001JgqFI5xlTYtFZFLhXGzFAwNbNBYv7cfILr+3pM+7LXnaRVFcXT0SSulD5pPsr
wUI7gGP6XiAgNMRlHrzMWSW72lbbO5tdP3BXHKbSOVBeC/BxLj/rot62jNFiGMntiFCk9rufNgPi
EZEcs9yJWhKSHlapmlIOS4nHr/FxJH5smKLUAZb7F2oXymjYFyTNwd+VcWyxlWNeNhHMH0CiJBP1
8RFkJu5mnNObrPKmZFbDIDygyBYFshdb9NBnbIbeEybGvUPXuouGqHisHS3I844LNYbkNu24SveH
igl2IHmIcHcKzosKSlESPGmoPMRd/1MbAflAhfz02HfanWFwQVktMaXV5FkdzyMubcGalsDz2vlb
hF7i9qKky7SrlS20sZHBmUnrYNY90N3fQhlrsuKOY+K4uj8pgDRJWj4QYBNKlO/EhETHBOHMvD2a
wFvCYL1MwmccrO4oCv+GKqbAQXCWLNmOFHs1evND1yP86piU4HBw8QcSdT81HQvtr/21MdCrTv9Y
n4v5AJ+bouPafRTm1f1eGXXTK447NZlqd8d6ZQqpLlk0e9x4x/r+3TEOwjX8OY83EiQu9kegvKxw
TkFgRZORvwHtF8qsreIyaggpv4UIp672Mk7+f+VjboQ6MsfXvExk3gnb4J+Vc5EPrQmu9MONscU6
S5+9YbquHT62jBwKDzlf3JZFcaJpGO23uTbBB8Ptn31eMhtxwWiRnJNt+ym7x0w42Ituh7+kx/SA
vNUHJg247tXCO4+top8dmPuUXo2PexQaJp7b19loSphWYiB4spacLF7ne2fa+dHxTYXtslv4P6pZ
j7nXdp60ou1zFnSqMEIt2EsF/CsYFi6SiNQTvwrbC5Osioj1bwU4b0VZ+EIX5Qm/ZYqbUv8sPWIy
siFf/3NXyro2pWDkObwrrsHa/4eRssELbPmFIRPCmp62Nkxw4aulCfnE5SAtVq83fgI5X0iM6q/m
HBAReZjaQLY4HtGP/Fz46SnUJqrRW9dI6MVErmrT1ezXqPorbejdrht2VHyqyVK+Yz1NFcxWoeJR
EkVmfNtqIblibFTrD1+Vj5xpISoMakFrNeWg9iAGMIBRLl9/n2VqaQs5zGqlRlI/zfUujbhXuIPr
X6AjE7UWaTdpV2vjaf5MfCCNJ2NwmVjtiwGbSIWb8N2qLdZtDNf++vHlInj0xn+V5T2iyJvUr+11
FTAE6ZmsAqxKxtdQwKa9cHZcQ+Zjr9v8MVMrIvBaPvhiaWGFQOeC8sAQKN4ZAb3pv6X1ghIQy5qo
HWegxuIQkevjpZhBd3/vsdMNkUtOUCAtfuc3PtV6LO0/aE1duZxRXhwGuYGhyts3WfkEUJaXrXkB
z5o5RIayr8iuwiDlQbgnCz6eOlsTVMQ4a/WGzlRVIWwJCv+DMrD8kWE4g5GWsHSaVlr4FH9k2u2u
hOCE40eiNoqEls7uPErXt6NxfmCb5SwBVQX3lfhBGGj05UiRz/R5ik6OeO0zkS/33P3xusC4mU7J
NgKufvnWgBmvIo0+Z9hB49+Rn2OTEhiKX0okAa1PnrgTH1zwjmq+hd4UcrSZdzu0TRhqcOyONxeX
nc87KUCIvSIPULyKedASOtWegMgbijlD0im4NRMtREHeHfjotAhMzYGRdZRg1UUnyIZGpdYrKPFj
U1wcpmD/MkTS90HjwEL6c74CiL0fdQ6YmzCmdNz03s2EUpBUFTOp/4kqDqhyxR0wzZ5WgMCOELZ7
AsoVmJgQhs38rx4mDRAgBkLMpDr0irlHwFgMZbXtMkFrE7pMeK60r6+VBSCLo6KUjgabju7pjOhO
TY5TFuGyIpQYRyozfpAvoFZbG5urd7f7yEpB+2Ygq1EXxYcjAk9izj6OAdu7Sw4o0PrD2L5i8iQe
608pY3tEHQEh01SEdHQ6NIVPSLRbltFnOu6rGzQWmVgH9Rgg2+3yaeTRBgiI8Hgz0IBjCgV8rsGY
FUe01+bf7JKKd2zcZ+iS43wMr+oWDjHDBo+U6VViYZzeztToO30ZD3Lp2b+BxJhcahpkLLHJC4f9
jRMn4w3AqcLFxULD9n5x5calz+a7gVeGjNYHspdDI0b+Z+PTuxkIvWY6NMcUdkPQJy0PtTKMHbZP
dV/kzAilnmDeodRdBUjCXCkDY7uf6uwtz91YNsUWbSvS6+CWOM4ECBeJC9DFRrve5u/gx9oeN2D2
VSPdD/1zZydqEV0Si/V1PbS1Y4L+A9rw1bhf8Yupsy2vvKyLiU55ZI+2ZBVYDhzyxYFZh7gF7bdX
3J0RzqMctI/bVOYlZ5AMYGgGbDPlH+qVqN8v/LdCbwoGLI+9usPfX5jXwtZ+PFrPI+uTTZWYJKGl
ncg/V8PufOMhr3kHlZUf5BpbV9FZSR5bWJq8aCsyWF0OGS/WevfUZxnv2Im9otVX0TmAKl7iCDAd
KXVWwdxqvDFCs+66FLaDzKvh4r98StoLUqOBOULQ01RaVUJfmjN3Dya98A0xu0V+txZjuzP0XRG5
JgJ5hPdXXpKZ0VszuR5279gUbRB0hS2JWuw7loVqzWV7JVcgpWnEPsmmhycp2HDcXAWyp3mScLMP
FTAvPZFNX4+Az6/SJgTdDguiyLEcoXJwlCizujt3n65qbB+uwr6zBpXy7/+Qs8XKXGhPW59WSeBw
U0CoXvXB870liPDjf20lVg1IOpJzIdJ891LdloTqDWWszW8w5tCYstxUb+16L0K8u/J8A4KiuPih
lB4SWZj1hBol0O1MR7mSTLu/Cd50ZZ/5zEyFKfm2gHBqlfaUjpVwQNQJGROebvKIwYFmODMb1iXe
p5ChddI3Q6PdGMipYrZzsxPrkfsu7R8v1JrsIquYQzf211vGk5dl3G5dAv5JZGUowqNZpYGzl+OO
VCo75Iwf0Z0t6G75nHt8sbtcAAeHq1h04890x7fReG2bJicTv2gdAGA1vl+IZfwbNEHUGtegi20H
nl/C0imjAOeS0ZwV37VnfTYTjbT+GzhjMEBgMXQZuKcURIc6ay0Cvlok4mbeCYyP6ALd4euNovYw
UD9WJ2GQ5L+9l8tZnTC7dsK4G78K4YT1ZS+n8KVCtn2IRJe0RTAMI6ojk7tK1Y4lMiNg22Nvdd9C
RFO8lDN0Q4klr1bVbgO2etZl08sO2SRJ8Vr3D24JUsHaz7WTcm7VJ+RxtRa2WlDTOeoFox4kPyyh
S1he1S6+vlfKPzsyO6YxBZvPOKnvdSPZHK8vFsni6Z7ZFqpH+p/w/mZZa+yxXm9x5Zs/4griTIjD
wYzUw3Qr1NVPV5/BVLPnm6q4X1qsZVHLm6XkQJyyljC2MyMtTUDBVeqNCyLLnxkE5HsvTTcPq5f3
2OptSc7xgLPgKui3abNN7fdWj/t1dkpS4GMuuYN5q/L2FvvQuZ8a+/kQLQCYc8T3k5g7dlZo4kR9
A/w3qZiSVfcYtx0k+shg6AQX4SiwLLaf4l1ddFyoW+eDcChToqM2JYXojAS2eFkgcCGGOq9rqB6N
gH+6U/u0M4+pd26B1IRXPn4f4YbIhMlVnbgUZjO/kJilozEHzG1Ql1D6gbsDUmJwW94DHuzgKeyp
zaYEVl/RSGuxkohLQqL0B80UcSJYngwxPvoZkTHIf1uYd1dibFxyslThRHVvGX3f3B1gCr2EJ2ma
tHZ+kHTt7eEZUVuRm2FwqqjuGrRkZ3HN27sFlA4o3pGTKBL3g/+F627xqQF9OOOfV5fdVuDxxOmx
bxwmLb5z4W4h14TAlVQbXEr6eU9w4aZmFtvSpFiX9DxvO/k4d1CA1+KNFA8EWuYzzGQ51ceqfQc/
HxbacKE3RI8MeFhivC7fZE+sreCdkN3FMX7wKIMHUJg4hcdc0RJjrA1XCsszvEy/5A4oU9D2AmRz
nDRdu2S8ROM2nyhHRwlso4ljGl/5J7VCq4zZgJ9iEHqidkkTfca7OUCPH98+VWxu2VG6VCbIs9Dh
xqXQDsSE6GGkHZJQ00qju5j7HaweEde7ShZ9V/kY0GKWC7KlMDeCTCUxYDAmrhKnOv16VR5I+U8s
Sd6U2EKoGB1s3BGZ7PsTTc1JjKvovN0H7kK2APp6rLRmxv0Ta+975cs1Ll3Q/GKui3C8y05gDof1
o1/cTJVn2iUr6uwH1qkxLHSSTJ0azCM8RXJqk7jf84NU6ghcbeZJor3u+SHW/jZEjSHxsrh0+Gwp
p5cK3yIavbEoJV83b1YSHiSV21eGqGmizh1ytaBj5XFmjGQB1i5+L2XsKnvDlA7MYbmC/UYZAkLZ
5iXzLRZVYeuA3NOvr8PcRA0DZ+EnanehzcanDYj1wai7HPZJMYo7jgBi8JTzNrLiVf3To3ELFL+l
ml2j3lOZTCBwrMnuOY7J6QuboogAhWIfGQ+uhPznxbCzvtNOaUDC2mtHuqv9boRBQ9uyMprRdiUw
q1S8kiKmdp0fIxUr5cm2nI1oUXsoZR4gSm4fRobP2rwgvKT/8R3p2z+dLKoUiWwnwnRoQ/VIwLX3
4WrglLvObuZJh032AZ96BzWTv6S+s9t3pVKdLkRfFBY6eeIn3CGbZNUr++k8s16lRoN1gxIerfYD
bGhGxpbgGwa7uFoptATI3y5e7BWyjEr/VJmKR0MOCcKFF2fupvTj+BCDb8NCR7hVjRN32zziKnVn
5lyOxU3mfmBQM0SKnVh4yEo/i7Anm+w7EdkvLLqfs0y4LkenALIXV2POWy+CxftimVzVtH2+ueDP
C4woIXZ2f2FcBJBAeXIhuK4ID5NLmKSW3gRnoPQBoPN2oXnriupgglgY+7X56wb1vbWplmLcIXp+
zQm9+HB2BYf6Mz/oR3uR7epOn07aIn1z7fZXqzIUUeuuquRPJynH8ze744f7V+P7H3PYCqTLUuoP
zimiI4yNWA1hxcPb37lqKdPkEpARh1LNwWL36yy2p3QVZCjz212Wg2K4fypkaeTd1nID69tEFnSU
/zjNEHLaVZ5AfWD6BnSpmvXDNdefY9dJSYd7xpBB57/3BnM+G30uUsz+zT/IPcLy3DrTSlYrL1+D
Dmdvc3Jlbb5urk3cxGP6Kf2hBBFqotWz8d6NPSgiDYG+HmZps5oCDGfIbfCZjdX00pbzBd7vSzYB
OR9ecD7e31kypiLNrY8cxeObo8o5f0IhbuFWeLN4iMEcKRq1izX3+aTdGxR8+/y5Xva8MrbPvj5q
YaNItvHXvXEre6KDCzyfyl68ZUO0AfEvSzm49f5KDXfZxG12UvD0H3l7ztEuczyJ4ujT8HGvrUNH
x0mqD7FdmUDoYSGbUMryseCBfSj+6hmoHPnao+VvHath0AKurNviYvbq89X7y5rejYsivz97U5KW
TzRSehy87M5m9Df42b7zKAWLQ9/uokVGyC9xIPXrtQR1JsD8Fo3bbLC1VSun7QDt0uX5qkpFn7kK
OGVB8Mcj+UnkYZYwd9FzNMYiROUcBekz3fHuYinuXJCnnBZTioGM6TuOsBrARVE/4hV3BRq0BWgD
36sqAFvwSYL9oHmUUKquilEGDEXNHl+WaE8/ByA6g3RX0to2iORB5uxVNt0U1JAPIALnToUfrZXs
jhYEaBDEEb+7ISDjgYT0m2iB5WfIc6qK2cppNAnkmZCNp+mPGh4FpNJGPdktnr2oG5LjypeTyKbw
As23PhYsS9cVXhaS2U6DbCfmnDnGhEf0ZzSuq/1wvgzSL4nzs68VnfkCWWZg50oGShhZZKRxBs7i
yFnsuRm+VtU0xqUuPkDaCG0SH1qNPZcBt0/ahWZDDNJXYFfoEodNQ3Kta2HCPzqEkLjQOSFPiOYp
xlSMM3yz28vm1UAPVCDaFv3VaX8pPFhej+jnxPHMC8hVIQ6qefj9BfDo8PkTMmxMD2NuXpJizjqY
rzEH5OFfH3eUCmRHjvf4BI3V0YnUOXouUVhOICYxWIjm5ZAZa2DA3QpjWeB7V6m1iKSxBxs3gTmR
Xcu9PAanyhyyaIaEyykgXnC9Yvp1odyP8CQZBbRv9uoGJ8wQtcGhAHOVShvIVZmMzCaMd1ruz9Lk
iB5jQfp1ykBmn7bY/5cnTmgFc2hWrPvWDxC/cPIQXtnYDf5gUm7cmN3Jk4rfqELY+RNAvntOek9T
1llS6T0DUmDH6w/yb8o8K0qLS6Uds/I7Ms6Sv6cDFWsjb7l9hEOVp+aLqDULrOcEdLcK/yUVMxT2
6Xbki5q9aVKZXBakgqnh0rhO+E7jXMyUiSKTMBzUNHDk38jAXeYNUohNZxOcepWxXgvda+MciQLS
d2YpudBez2mWSIfMRq/xdEtRuR9Nu8Wv8AoCAoYjm48hAovJlTP9aBIp6mBhvLhEtx/d9+r/ifF5
glhIg/QITl8C5QvA3Wu1QzFY6Y2AUaHJbMT+/baA0Hn2ksxBEKDEFhr3BT3dvLlvCKInLyRu6jiE
DPjMEoNVITEVhTidY+2YA2f+Uia4bnMSYBQc7uoLBRG6EK5euia6Ar0Oceh2b62S9K8TGd6QVHHS
bsXfYvhUERBp1HEp2GGUTndfd3pomq5jVJir0O44CZUjAcB9XYlmJLT8u03T8RZUV5wo47kMmrvo
53kzlfdTJ7t4XEhrXIBv0eRHeyerMkaDdWOBxS+HgwcOR5E4swrLRdUfUcnZpt6d7xVbZIq38N1f
AedJphCK7Acs/rjO5etSEQRoQ5RE8J9pUspkNvcj8G/j5CvDNqBhSfulyUINc+IGo/bjDu9fKcwR
+u6l3vtinPzp8w6uiID1ZKFIlafLFDbGmpNY8O7nUJXdkBzw+WPWZK0ZFbIB+xcWW8gjlNQJkO30
96DZNSeqZNwEDvop1n3N8RQ3yK9oTAtnFMBBl45nWmJHSnFHWrm5TlhX+DTFfRe7LaGuA6cp099U
omgqOp4ZQolmW+RR7PVteVQpJqGVhaU5IwQX9lcBhFaFEsiuvPY4jJdFdLekjObczpXuhHRd10gB
MMsJt5dGy5l7x4N27oTuTy6K0JzhdZ9Rse6oMHka0f4ZnP1zWXKkDJjhAjYuk1AUSxOheVnba1z8
vkP30HtYMqu9DRdwDDSZKiwAgOGh6tT1lpNDXXRiFNlVdrQiADTVb0dUu44B3JlvwO46gp1N4FV+
AXSQkPGZ6LFToydy+XewbLZeAXBwwXDHvYqAlCwr5l6v6ZVXpisyCOfoGGWYu+7z5e4b6klTJ+GE
dBv4puigyzhbEWsvFooeWXxHZuup6lLxQ21dAFvLHnpet7LOmm6dXKvl4ebcIX7llbnhKGDTSQhu
23LH8itMIAl5+jylkxfuNllfSiroE4MKOqg7ap+yw3qFmzKFD19JP5dMJnsUkJksGkoftmXV0lse
w6U1o/cf/lPBBbBcxYZmEF9vpLZnPcX6E/AelxmpGHKdpZ93bRgc1BHKctDfhPfOnXckqltQMOjW
2+QrHLDbsEcDYKl8Y18N5zJ3JyJAo50rznxwMVS+5Z0zezx1tyCSYww1uhI1Qn8A7aiDE1OohDza
SC+kp18JI2DlFgMC8W37/RVpO6DCHuk9T6LCvzMtUCB8YNZPRwButcUMnOSS3Bujn6LpujIk4gfe
HKUGZZTwWWIZqg1fD0lSV+1y+A0/Aj7QqREQfa2j8jDHZS5ShL9+ipHAnr/m8XssjDso45Su7YfL
VcgHxX4YW+0860ySxi4tleMlOly/iJwtWovQiAZAvwfQEQHbxSRDD9Np3VogXYcmKiIdofoFF7Hj
4OevZivspP+agv69Uw8LcYZpAzxKhmy5wy5mL1ixxElE50ZO8r4TJkKm6sRT13wf5QBP6DJGb8GY
Pa3oGvQEDMDoMW703+nhpQmD2zeUW9BwHpfLAzM6NiXhz25bKHDoybbpxQ9I0kyliKOciUf5cMOL
fuxJUBVWl/Duezh2g1m1m1L6+jtq/hEzbg/UnMhYqoN5oLLJdwFyuEQdYmFjEwUrDBcJyKngR7x4
8+01mnwroHKa+AeUgNh3kH9yp7UXY23c9y1at7NewnWJC4AfCMiY1QttLqRCOoqXcLq79S7jgsQA
SY3ZWqYAsSI1wWXZ1YuaoVZ0uLfkKA5moUBS7tE+6MXfK6hrHhcYAtvBuFu19Xf4kaZrD9nScqTF
e69PEWIKtrZzQjvULTylXw3xNRZuDF3Y1gsoC/uoBbddywoLHgqiUFDSL6Iyb54w+XrLRqVOS+Nt
OkVxZ1FXzyL1pR2qytKuEJeGTeXitQPPHkgkc5Dcw3mjJhHepraqIq7Ne08ufBqUWS+sNQG1rfGf
2/VD3hsge9qe0p83EFFkhEBzh6FC+O/LdtgWG4sOYkLH+dF0XZCO6N4Jo9WW2AkxcD2BR5jOzA73
W3WgfZG1TQ3QObyamNxQJPUjGqJz7jvqdbzRZzc9MGP6CbjccixDNqt5LRkvxzxBvE4phxcs5qp8
oByMPfKerYJH9DbVQs7IyVv56Yed1HjyB/v3JojgYmCfgvOOtvQKKVY+5swQMh88KZ5kKqOt/ttv
dTa6PpirKgb+r65L8oad+nvQsQsbXJpgGScMk3Vj7KF9xICcsaDzlJCUU/Xf+eXr5JBS2BgJvRyi
pUK/3QCIyD8B3y75cVcO6G6odmKCAD2XETKLRtZyzzVEacb6Z6qfMjYwZG5TPwlb/ZF7WTnXD2Wd
IBCkR8i18b4HpI8/UC0sh4JmYvPbl1d6exMIiGSKQY40Yqp8A5KXnM9nlIK7f0X8X20NbXJ1KMYH
9Djx6MZ9p34xPG7AtgLjYaatdMqIFki20dYmJSs92MWRvL2Xp2oKUcJ5ZYtg64rzRWS3L5lGI7wP
8cJC5MnXnq/VIxgap2CTWPic/ri2Vwl1JhBQWINdPVhF7ZCt/sNKJWq+quTwpnoq05xPA7btBHyN
Y84SIdq5BR8E8TSjY/mr0UvXQbzeqtjdUaroSXu43NBPwDh1X7UCpKp3yGoAwHPDP9FAUc6HejPz
ajjTyM2TMJPlCCH26Kku1iIyc0ViUJKg7GVcL/cb35oSGHUoEkscZ4WUJGzziSQqwPvG8ylz1FBm
hSfwpYhpINCwdz+qzFOBk4LEwFtZxqDCYkfucP7D0+1W43MnYXdawv1pZG27pk+3LlZa5zBrRKOj
550eG4H4hkzDj1StuUagPdkUEsOnSQUrRO+AEwTdyNbSyeoI7+7A1y4MKa2lVSgSFt7VFekmhqsl
iiU1i+pWPu66AP0b834fYHrLr1zQ0/PAta/wzZXN/7Kqwk3iP/gkF9QH2qxHavWAVgfPwqih2Fj1
uHDcwVIK7VytExK9zDRhnMX4zt2qk3lYbw1FBuaHUQdnE9UOvTl8CNXbIG4JwhEOoBILxq0supp5
IePdDPcsCwJ0YCP9ATo878+pIQXAeHCce+wAVLuAVsKMY0ZWP96Sb6jnHzvWSy5/sDWwO8rkHgx/
szBiWh94dBQaFkOG14DRPF7lPyAtAg+P+Q0/EOHE1DQCWaHu7luAc2OPh0sV5Du8ucsfiUDx4Wb7
JbWMalkschbfWLXs4UJ1g247r5CvHzF8Gt2M7aUDn+571KxSecGOXHADqKLjMuY0vw9sqAMuheaj
6OtslmZqIgCBEOzYfTgc2rrL0HWmqdh4zddNj3lPb3aoQBo9mI1+Qrtg1FUvlL1WGGdu4pT0FGHL
3wQ/D4WbVxS6XqLqkTp2KH3SmT262e9tIulGtWKFw/JvyCob0CDivClt0quG5vKZ7w1yOF6wDwr0
eNIBxucCmt8OKzBSfTsSHff8c2x5l1eW7TL+Z8fhO5yybhlzMF9n4qnpBLOeWq3nWPAsPkwiIKTT
fgZTf6/wmfEn1fp5I31WTsuSx3g4BLRVTMP4O9mmDuf6RKITxUJfBbHRi2lawEFjq4zdxagtDA5I
v1nHf51zdi3z8RvgddKm3I0vg/vzI0arevKGzw02ckiv1i09IDJryrwYo3jgQnc2DxykG+2K3eVm
qg94Cw4BMHgBlcjeDyHwqYAQUzGEGIwDk2vpenZwFM2IP0S3LCIaIjVPigkeos8kG3VFrckapFJN
MnRykgWqlpbnxNq06ACm0qrck8DH+X7gLfooqucSrWeFxGDh3+7xnaHow9RAOGpgkj9wRF2H59NL
F2NPq0MR1Wq6Z9Rd9O5OqHiguM5CTOrZJmJjZf4iLpEqUCXNlthkwb6WaFjbGxDBgmKQSVs+hctr
zL6Mhhjx61m1HwKg/hge4CEaBiLPjZ4+e4ck/o+RFKpp78GX5c+CMkqABRt5zlLKXhL0cj/turhs
fX8gdJTW5paOfMKowWprlfUy3McGrFE3BJo3bt8SlwC9KDysSU7PVMr6X2mG8pW+3ahKUn2FqwQB
2A5JaXrlA/4PkjtskVA0PehDkS4b1hCW9rYqnpG6q9c8gHCNRjLUchUpn9u/XnFeExvG8+2UIGon
NLhkuxAAROYCzj4jVnP2wIl09zQ+k5YSERQ/7NV7NnmxmrRuJpD2ttc+UgP3KTtL/aVJzjFwYUEz
HWhSk480ojpaxSmgSwWO19/LCnWVNKk19uZDifb10eJfrxTHAQcbUH/JlxMmik7KX6H+cWtkKqAw
A+jSu4Rjd/xr/Gobd1WJuoSDKYEZ4Sezk7gnmkXZbQA3FdCy4moLXO1JfOBflT2UOk12ybI/DHGL
1JB/JA5I0xZk/q5JjWZrjFCe2vzggS0sua+ngz5gjfb4i/mdTne7FNJGOYvOHdejwzjKCy8MoUxO
TqgQUSo/ASldnH12Wup0iGPBI7jgtgDFLMPItN9X+6P5bHLAwdT7LaaPKgfiXj8TYfD1nSbJbSl6
zBDxxJjmnOOYdl+RbR+mArzwpSXI6RBtYx2N90IGuB8n9fb+ePkLJ5k3t4RQ05sAtFLuZOZlm6t+
lsxukJtPLAcTSrfzs6gBwYuA7+eDPz7tslKT1rJxSVGdUNA8meItxPsCNEPdEf0rkvvjS8+n4Fvl
OPxRwyaeDvcoSpHsss1p2w/DA7IgcmDUyVTGAvFVsILq4Hcg0t+4Jk+Qw57LkaW8nglmya359haS
jcckjINtsFkpmKN17A5SpeEgJVlBbUHuhgCaajh8Ow6FOUE474pxvWl5oy5aGxz3EeM/QbYBsQ0/
LXG4tvT4RIQKpyZafIgqG91/Zf3hlnPzDMaVkRxoJVdHkZIvDzX4OIC6U2ybl0AjfOX/WOPYsJ5q
WAwFVATosTUSuVOfGnW5EJY6yP+lMIQBnNawSO5TSGk0wyP3BwUChxznhX3jYnnGJCF+MS48dQjq
ICKImCJgoitQlT0ReXXSNZ8L8+VPp4EC0aBsYW/pVcf/251iMTW6YZOqJo4az+QY3t0A/5zXtA3m
O5gPkMXueU2zVwFgZBPZ4qVT55kbDOBxTr8zSMuqJgD3b87rMcAFNn0rfWZKrIdySl4t1ZcOO14O
cbpfV+6IQUd9FhkbjghuhyqVXFMZ6pamSiV/1nVOqLHneTvhbCDQ808hNfmmigx9iWh8NSdh3I4g
cW4/PChNp3+ZEJz68Wjl/XbU6wtoBRdA7MLXZIzLRBmNtDCQJOtEf4Lfs8iHwasrKad54djGSjy/
/HDj7rs/s05Rjpi/HxdSaVl24k/TrCVD3z+N7IzhxnIcEwmm3JLurPAvC8pHQ88lzEoTDdLnm0aM
DIQ4XWxFz2d1digYMPZkuTtEYfIg0kAE9lMlkfQRLGkE6WqhSEo32Eq+mN1n0JjMTmRlyjuOJ8PI
PoB6XLXbKOv6DqCCzHM9l7zjpl+FtCAXKVcpNy7RxVnmGez4ZRNvHoO/oUMzVrX4TA6Sz1n3A3J7
O53dkMzi1vw2NYfHqGtop9J+TNb2u+Wl977Khp7GC3cGZ02NZczH7LCwIrKbE0S5YagNwZsjqEur
Gmz4wVH+CLtsaqiiBgCQ2tUoef48DZh4unKnKXmpOjGWGfsVI7G6ae7csb1hhHKKj5HbkDnRHicT
eethKXtm87AIJd/sNgk2D3ilwfD+I/QOQ8hZjnSYOJ8rFY3Gz/KuRW81McGeanatG2mo+gkSVGvJ
x/mi/XPKQn2VIGp7W1QmjlJpU/BHZMIdLrlfZ2eJ6sV0HIcN23/5/TaCMx/2eqqaku3lVHmREoHa
T5ep+nokGEUmQvTS/1r7OXIvDh7r9oR/d64QypK289wTLknX9Gw19m4iIWUBFUqY3o2v/v83tVox
EOchCGM2kMjrpTPp6leMdR1cUPlCLnHC+qoQs18apWrhFbM7weO3h9c6aVRcX5KPYYV3Fr1VSeZ4
MoYNN1o5Ub69l8/mQh61ZQ0AVW0hQDumtkdbme+iAdyfItUlHQdFYPng7G7o1IT82X7nEXxssxB6
SH9qOp0ldjKlriNzKjuEt1zpCyVcB8p0awBP9cuumqjvxGAXHuEO8/y8wG22IoOfKc/2qruWbO3Y
5FOMENt8yi0xM+J0Z/8V+j53GOR8a243y7oRfgA5OWVvKhwCcG1Wuz2/EVAACfCln5vZvjEjVIXI
WlRdwf1cFX9etkPdDcCSDMZ7MvUc1Uw2i59iJvZ/NqSh0gK7L/Sjx7J7ZL2Mn4T/kYOq7F9ks989
MemEj7pqfOM5Okc9TT827wV0ywAB6BtS9hzKqusW/Kac3x3diQqRDoB4BYkjv8J17xasdRVekrju
jgnjlOGmv7Ok+MFwnZ5fu9Cjodb4KqZ8ltFCo6rMat6CzhLgHvxY4MpYOuN955F+42120d8ucGd6
OugNxNky08q2JBBHTGQoXL2Af9pu7WCxuZxpOV0XF78h1q9gqDylxLoYWAleOltczErvL3SQLbFw
Cu6if9Y9Vspoj9ld60XZ93KwtbHtuCmLKQZjFltLA+MVI5PQZC6rDxkSjBxVek6rRFxzO2yEihVA
rxSIbMM3/Y+kSCE8PVf77ueKBsxL26BUaJ+GW8m7kUMGftRoys7QLHAZEC+GgQZQeB3JTuBLjbHH
Hw8DqYqj3pcmfl9BzssPZs8TWypn21OAhpBM13SQEREO77T9AZfOlFEkTjgvngHUMVArk5hOpPYG
tSaes4J7Z8yaBmBCqrxVN/Wo7CkzHGETK3l9R7eyiGrqPEkSuvHErofoRCDqENVQtAN4JGEs/SjU
9vt7JS/1xNREwwRzy48uxlysFoFK9a6bpGibBrSmJRm/BNTktyHyqaotwZE248w+10mSHje5ONC6
IPQPSjzH6jIvRorm6St71NKTaaYcur7heYJOT/GzoBLLIHJO2XyGHO3OnZ8+glqQbhZNEMHdCGMh
xLC2mpixpkNPhIjkVc0+Rda7IgtOj0KQQvi/Hyx9GHs+K98Cg1Gc4vyxNXjbpLVXuTakD+TuLh53
n8Bmo60rWR02akIRbxM5q1/sFvEtP7Dl0zTKd9yXf8xznQ07Ej1w0F6Ttxsk8W3pKeL4eeSmt/T4
N1yMpLy8serMw60pskPknAs8h+RydxoDOf/5K+YMmzFwRMaMDlZEaDjXnMWB5B2/ujC2995YMurm
LtWfJFJuKsW+EGZIAGEVn9RjjACMHr+tkCuOiU+r6CpOa5J9rLqP5Do7j+pE2p0gMWLf2Twu3iFo
LEYf1mxwHUvAc/iykR1QV4X6UafbJXUnMK0y/0W8HBA5TuPoY8b0o2k+fvGEQXP/dgGB0UsYjW9P
EAnkJlLUblHFfPxx7uZ7bk4M70FAWN11K+i2mz5hV5lBK0xcTRqeYiRo8NirKZm4zvryQgqnoU2F
8j/xIs7NRn3OpoaPJrozWY8Dc47uhF8cSCRlwbyWwNJ6W2+gNdEofIr3WUDLPHkQ4u/0lTI0eKAZ
N6tWdy8fEnm/YX8FvjZ5b5ac6D/0SaS1RZzg5MHL3adLCmKnPJWm4AAdywEMHefLWMOJLdeouXCm
mnwUIcPLK/mWzSKImPrGnDrPMUG0jyeLAj+IOdS5mAMhzn8tZdDKIBB01WnMxilp/IUbefwu2QB/
eac+3/uphLSEWCmrRUwr+n4CEc6FmoREYYy3Hp5nnZSUW8fO9h0k5VOu4lLAIa3ByrKxPoCUREdT
Sw/yA0LOF6E1QvX1oTffvEcYycfCPHuKue1sFybQjgSN28wTCKqlD82aaFOL809cEPdEoX0AOCnP
i6K/zFuyjBtXUpgfhY6kHtx9VrxSg/pbA18/l6/Z78eHjJbHauFQSSuFfSXt5Fs/vmh9L20uYUGM
LHU52N3s5qe38MONzlKvj9KH3kt/x8tpmlzq5VhMVk0TaZwmHfrusLRbCqneA1HT1oIqSdNQ2E/c
N7sL0pxR1XcbLvH+YMcR4i8I3/sQQxHYgIswDD+BbvT53e50IZLpgGnaPOpxBoiXYQASbPVAnlr1
QqCQOAyllRzLUuPXUM63LTWk8yFU8P7LsTNCd9wnsnnm080H1c4N275GnzPEusaOq83RUprZHG2I
2T0gz9gljsfQreQwkjwDGpQQEEv6cP9Yr6818HaVzLOM4uhakUqJ9+ucliSwxMNMWVgZzvVJMUx3
mx5AILYp7hWqvei0GP7vvogSlJUoEiJdlvxVO/dNo/hfUrXcqhfCxsCguVlgBjl4YVSEVzluhutm
EQJr6OUdJg8ey2Pa4k2Wlp2NE0Y8BHazNLE4dO5EI8IP34eb/rlH4AJzIduXhDRNlndMmtjwDTnP
BdGxVr1VSBNwOF5yQcjbMTNf9V2hKtj5qMh4w2Gl/uGlpIaDLIfJB4lfKevYW5ioTyI4IQwVZfDd
HsD3BIKxUb+PR3niM4oXN/Lb1+qx/n2LZ7p82DU79KK3vH4vShV3rnmIMlgM4maWt7Er+LWmAmmd
O3sqMN6u6+csv7ah8jiRFpNBeItImPBva8sOce3jQ1a0UCpWyXhPZYt+4kfHCQL4pX63NC/UO0AH
zuuXKzmR/UZk7VYX04YzgJb9/Uqav9pysuAnckwq5fqWceC8lipmb/W2KbD7+z0G7AVPX9FdMcwd
7WGGCBIlUlwR94my6azOJPxqCcE5SCkXPqy4A54U8b06C29kl8dECX4y15xos0K5mRmbb4ubGgnF
SHqIeLHVPg5qEEu+0pGWMzZhhvGdGQjgr+eUF9vcTMiB5vsXygq4V7qQIA5jwPY0Ra9G9QskvcN5
rowaqnFEHUc/Q/4MBtoWFlfW+S91r8OXQJWJ4XIyE8Ie1pBxeYE+KekJOKMkHJM9NnZncaY2jEIO
0fqbqr+3B8DdxDsejK7jHienydeIigsQgDp+BG+DXTMyGL20w4jzpUsfh2392h11XRaeNfTTcHY+
t9Ig0MYvhJGAMKeZoaSm6xDGghZLT9/phYWyOfBU2YWUdxqTw2xYizrP+BDo5TVaNXVpa4qXZwqj
axbQ20kQhz2i4l/rxOFx/boYJJxDsRSl+5/MWWCvBXhgEjJd9ck3lKw1cG9bcYu1X5AMm+O9zlgA
mrjvYmTMWwfgXepZxqOhIkMARZ5rb6FLYexQbU8xXtEbW1uooPpmzPRxFzbGLR01cbfvFFulcNE7
eo4QnMOeU/ATD6eKfJ8W4TblBUUOkUgXlW1TRpgy0hFSra63YFs6NN2o0nF8PSa/Q4Lz0EhdGl9j
bCT6lyITUrzX8I0EX5qrq+8v/5XXx2gOsK7nYv5ZszgfdmyUv/IZSMj0+pRTnf3je4jPZzryuMYB
0zxgFAhvh/hhuT6zH/Fhv+PkAyjAo9ZSs7YVxeLfFYwChTWc55/9s8uho1E+1Slds/mGQAwJApKe
stM5BDC7e28Dpqvuy8m7TKoh3tEOva5WSRBHNx2BqZzftMgKO3N3YCRh3xDXCRVtq4fBfLX1Ryer
Adv20Zr+qUBWNIMRN0aNa8irR0UTJW/Sc2iJY3bpnjiITRhhHFIP9O8ZiKrxzYg8sHr6Te9RQg9q
hRjc9lwzD/PC4Tl8RpuC/xewUcJNeIu1NPCleVsr3173K+48a8gTe0xPaOQNMG/Z5zP5mTKG1/Yc
Bqb5APscm/tOSEsaguO1A4pZiSR0AUrqlC12LB0N5BC+G73NQ3rH0dT5EWXOKRiGqlechosruhKh
d4a+3b/6oRTAUZYqmsSM3w/TxTOYvJM42JbrNv2zBvrHnkBFeZePDfnTZQ/A9AhjXv78MXhVZZx4
kPrB0XBgZH41M0yy6tkgFfrxt8GKbSdTCAVGQSA7hoc3aOmtXUBjPt33xTof048RU+spYzpLElIX
A6GsQfk3wWq77EIuowexXK95OZyl7+2dEsFItn36NDRGTWIK7Vk7l9QsAViGxMDftZ7Yc6b3mf8U
0kFBmo1imcQ4l0I9/vp4M1EiSYTZ3ZF5YOTZxxGfABPl5af7gMHY4+rvjws3ipiaU2oZDd/Pq91+
igKaQuXik7swHdMBU2PsJpMg+RV/vIhuD4xIX/cjQ6f1iVlzrjThM+81V0+CcWiYNR8Y88N/pnoK
679KuPpzwJRY+kxqnpnYrzu0KNLb8i5sQMz0qM2uB1qswhcYs8rzYHPWzZKIZb4nQdfAwLbnbniq
yAZkYf6Tz259RvVOcLT5qCRQ5c1ETOIy2K8tUeKxgsL7nS55P3WDV0O0MwmmJzgmCVQmT2mRIJoD
A0jsDxJqiz6K5HKIfMrTH/omKZTVyx/KXyCG2fklqLsKnk96MIh5Iw2ykxXMDx+qPKNK9pLC2NV9
ze82Mmoh1F6zievmMsH/DldFcM+Fq7PcER/tySsfHlN3vrbqKv+yUvPHKaczbleaQSqnWk+VmLt4
V39khwAln38s82y7hQVCYfT7b4NaMzJ9zv5oiaXAgSwjqgbKWwuVBsUyanUv9Y3RBtc5C2UbYSwR
I/OmwY1uPVDLZ2upOr1StJM5tj6jzihPdF8p5uUXyGTplqu94D8glbkG1HPTG+S1mMs5fZjRfrrL
cZmvLniuU7/sVMlYmnvmzvDroXa4i6oi2D700RBYpEVoatpGFElzCehaFyWmcR4a23rfN9I8YSva
vu9LynQTJ7PhGh8o3PQ/7EssBT6tMlP+EKzNfFYAAZA0aJjv8r1IxZaaNcrqw9k4CGpeCh59/NsT
8t9q/GHvNCsqYirNEWVM2r4+VyjjnVZWAMelJJxaM+p/M+A8A2016LSlyYK6N/WtXrtZAFSeFrRZ
gMvycf0uMIJ8BR79Pt51tO4tNbXRTHDzXTcVC8uKacSmAJOGCMO6XIZMWTvIGOMA7NWLcNCOWY6n
QVo2d2CPMz78ILXLwhu4PWELajffTThpIs7mEM+iMsPUj63DBvDJHSxtfQH2eqS47xaQHW6MO4ED
OERWu+pNyK/fuEm3rrQXVwZgs0QvPdfgsm1HqNvzybjic3eG7id+7zgXP/RasCE4r6mBLrC1Miuo
s/RnWB2upsBKC8GKHnhPv8w4va4+VRmLPTHG2ARJmlBHMCdOW2gPfh0PPQ0MVQXbOTSkui6ocXiK
R9dB0gtQgtt6Q8o4CaO4oiC8/Fr1ob2XoJ4X6L5rTkMcIy7111l6+2FQdGQkXWfmJCFOVkUG/ftK
g8LWo4UyG+hpRx9F6IJqimE3payEeQoiI9Krzbn6LDlvR2s3Q/r2jFyYCU3k2Zy4wGoxDBIe/U6X
1Div4MkCtJKuFZ5OKB4c8N/DOq5UGwunQg3clG8dJU3l6j9vsDppYWy2rT+S6yJS3I6d4b8tKWXy
msBM6wDlYUxXNTzqnykBB+HedTrDU58wTCFqEW5qv/Esn/YSf6JeuSxvQO9PZJ0cwXok/CQA33Il
dtnAjp84wu+K/FsOqgzynKgz7d62WVQLL+c7WHp/aJVqX4DlVYoeGlKWxcr6KXPLqy/j7zywcRRV
b0nj1C+LrI5e76JEKUVw336jkVKRGhaA9N4kdATRIJKyNbSxXZkgu5txzVnuhoyzq5viPcf/f5+1
Y0lHMNeRcFNIjgMITKU0pCWd0Fg54M0aAHQrJkTfxcB6Rnz5AImLiET17irCT3ewg6SMBypedb6N
N9vXH3HOJov9tbuKPHhYwZPESJ4Re8OyqMj3lhF2FgML9hjSTX2/Jz19mjePYLmOrfiNy//s5pFr
NfqPrwouA5X8Ln8aTBh7Zt2aP5LfCfY4fYoeWJ4HiMju2iTcGy/B98pQLCDrXoHn5MinZ2gceMZj
B1l41LDAOSp5I5aJNKpvsL8qDmzcTlrocTyqqDNfWLtDe6tteGvs5PiYiB5uegdmwwqDcHW1o2cL
DzYwI+gqhTFH64IbSw13SbF5ghYiQqQUREJ9rqqoLVXzqk3/zXIXGjyfyVkPtHBilpNupPVlEu7k
zfvf9oTknBmf0Jb7GR1/AmOJWjXIC7DqTP3U4hWyevuutUr4LErvkjvt9wm5l6mx/ueQgjmjkeNH
Jh8mg08jfZ5q0TE9NvSLc90VVbMEtYVg4zXNfhw4kCF82ndF/0rp1GqXNemIpfG1Dp5crMo4EOTR
ngyjJz3WSz2rvvaIpDowzwkqzgQWPSRjpnWz7p8XiCM7zHqQXF/FPcpAf2JgorTOuxESLv36HCWv
wIdJGPGnYM+VkUXgyR1PVuWbGhFwcKTLAGUpQOysoWPj0+c/L2jG6dXESdlIdO5bvhi3rB5hjRoQ
DGbCYZtK4oW42dvPJllX9Hu5LUduVONu8o12Rlr1RT6eBNpspLhMI7tVVPtZYPAmV0se3CYHxyZQ
GGsxuN9erzbAA50EcJZO4FRUvICWjLhKLV+pwCrTG3fzkf8f/st2o7iuEsa+QSJijzj60S1+6QI4
eRzUPAYE4SzoLy+Whlw31H8Ck1eBhZLn63d6JSEMzPgl+YNSgCg5ejCk9hMMVK9o5gQCsnFv1rE8
DoXjSslWt4OX+KKzmovtrPExV99BFWsgEabhsbTWYMS7yTKoLB9lUMOnPQokq11eaI9F4hRayuGZ
MLorMMezzTkUA45QCiw7de3FcPntqfV9i5GKLiAP6o9/fI6NFtYk6qZnO0IXpfrj3ygdaHlCRcYI
cj9Lc3JXAcpTFch/6xziG5R/+2f8u4a9kQvZUxfZJpeFd4qSO5QfQ9cuj4XRPbjlYzVW8kW2Bw93
lNMjXXWtWAuEPDx2TnJ/gsxnFci3zaGa+EzpiBAO5q6tijdzPOwUgtoZ1BV6lgZxHzMk9z+zQRGS
jJ8vYndTVLibn3eEED97qewm8iQ6cWzcA06Z5Lj3hW+1lO8Z3eGAsLIuE7tMf/57VhKayI9A1Q7h
fuu7E3auQtvd/c1Rg97hjjJ4tEb422dQHwlMA9aFC9z6+XCSoDohWCcfXUSHdtaYQk4FGYiOvXKX
w6Ty3lJTYLju7frkExq9ip52YAPslPJ4dzwE6OdioaahA6PWbFpey95wTZSTlSa7mJnwQOF8JzH8
zdu89MyjaTB2asl1hH23Pfpwg259sPVc4SSDO5LiX2Y7SSZn47laM25+iDi/WuWD+z1WxD+bW4yx
c+Lo38ZePFrhDReF8G3579JgAcfGf7oBFuMWEnqu3zJxXy+Y//QmaYS9gWDaB16vcFyZETWMHgQU
PLUJbvCMzTJjfRuNOe61EIiIlxReBUbjrNZ7gq2K9tmniRUL9kZud1NZIgRWLyKWnQ3Y3E2olsLS
IHOCzVneb95M8VEqd0vyBtM+Otss7ZWptf+U6uc9WTMmN0V3qj5Clcr4UENEeTObrn2P535tfqrn
+uj3exeCf8mSTv8e/y88dli+ZMw+s2XR63HYaVV0WtaYXGRVl566SBRqFeQIuPaz5W0gLL2jdP3I
HYhfnRs0bCYERF3rGLZ0EUx8qAq/zPe9pJlgpjFXi7WvBAqVE6NJiorXWRsz5Y15YEsJokVQ01vS
HJGi/GKc+lh5mAUcVNDZaX/s4tEr27ER9OaG4qQ1yLwGsBcYBP/Vw9VMfSJ8TSWIl/YRhCaHDihZ
JW43U4fV0Dc5mVYedxmykgkNw/JQ7ro24VgxF51y/Miy6qv4Sd3O8iG8KDsGXr/sPII+Kk6CroQn
eQf+Uh3rTGSR4cSL9W1blV7uTuoRaUhEVpt3OpBD0LH6U/F6b2dtAPgx3Sa4rn27nrxjc78cnuFr
wCKLhyb0O16LNrEulV9d0jYKZ+Dohp5MX7m2VmHzv/5aSvXOwssiassVqiVVQMYNHm8gc5z0Y6BI
p2TZlaDMDmUuiDbLLLKkadrZ/md77SD46jqK/gsIVwTJeFvd0TdY2UYhT4AxCnIWl/JXB1ou0U2m
WjN7tS5AubC7TlfTQ0G6aO7CT2TrMXgCB2brYQXHkuoIO5UdiljKtaLEJRDWm+I28WQCFIWib/zM
cWI9HWNZtRtes2pRkJcmXaiO/ZcsZw08oq7pM9qiWAH+vOeYzZyRMWpuxlibJNss4RLdV/NdbsU1
t1BrB+VLkXc2pr1kc9SdLvVNwpZtNVhEE6VNdjXm0srjcpG40g8DzfZaaW2vgFg6z3Vow1Ys2dv3
a5nFQtD0ElrzdzeOYmNrf5QzwoXjTkpC/DAge70Tys/B4ScYq5IuQrdXoGxEO3H6TW4lsLXm4hWK
sozwoAHO6jAkaqd+6x3BxC+qUUYdH5rLGUwvk1qHwGvXiljZFho3SZs5Fbx1gMpbeqgEC8V7Mier
LdxbDcurnfWlgsfegiOP42+hyLo2cHZcJ1l7TJzHE0Sg0MoGFbZNv9FRRLmn7mf0AHzKF3hmkRlf
898ESOZ4SxBHFySugtpU9dFjX+k5/6YwAThN0P5fgoGpbzx2ZCjUa699PpFEzO0d2P98gtLu90Zw
EnxozaYx2qlPd4jrK7dkQu4rp5lmeLiXvdpR3RrYmxA+oZVS5/aZ9TJVcbvfB98k4wITjsQ4/CrF
EGyrgcyNhHF/HqFX04xcdJdJwUHAPq4QUj0knrts7vN5HO91BGM4QyJk3S42Asq4z54dYqCqb0ia
cNG1SiYHwYCFXXf7JiOlX0lOW/GHZ86KNwIQfG585KOouqaLgE0YO7mP+Rw+LjDPiuAhHUx+1Ns+
IBxYSuP7tEebpk1p6dU4CO+q5o7ImvsX8fU2hbkBEnw19/wPqsVCZJ6WOsSYQmGvMmOqgrM3TYlt
VYtrDGtkZR7folRejXl2TBjtE/YLwEtUDNvU4dZFSfvzJV+/MP8Jg+Kc8HOlfVfcWIlo5H18XS8q
h4OOYd6gEYixDrzG6dZ5WJ+LatrcNIm83UXCEdLXDjUK2Y/6eiOliKEkiktfHWt4jaDbMW11XTHk
N5GfNrMPG6GwpLWyCAqLNHr7ChbklvfcD3fZbTJnpDZnqUDL79lOfSmPvPpvvFAIB6+JBfNPe674
DmH2euxX1D/qhSk3OF/Z5TnaG8o42zWvTdPtO8qtES0YIuA3o+tcJxi7dlWdwSKhZGjiPUib+Wpa
HUMdEcZseQhjcjcaacjfUf0+4zFoD+QC1R4PhWiOMIcflOhFW010D1oN+XsNjOn8ysafBA5pLZLe
YPytrircYUGeQYmixRNMlFoC7kfZ7/17fqJLsiwzr69dI2SVukpzmhdP3bXtwdTTXnLAtyRr3RKZ
CtULfunL7R0+hPdVbMe4++3jGD2JkCuxMHaAZJC8l+6f5i844SIH56uX5Dse8CW5uAp2FpDI0Ge7
Fzzu4fqVQCLKmuFhBxl2QtMbp59AAVo53GOyaPA1/TlFO5/5p3ZA5YYEGwMzH/T0GT1/d90j5nbl
wLIloDTy79jV7fjCcCcTjJDyrYSeqsePTXwPgO7dHwiBaXE2LVkDVjRnxa7tD+NjLb/39pPXWBkc
7sf+9J5QDnHZUObsefT84BqO3Qm8m997ALqqp1kGT0JHaI3m5794Wj9Z0mAmKpvOb3xuG6ePpxOQ
/QuLJnHSziY5WLOJMfpvQxv28LvEgiP3cOupfzJuAq0G/NDP5xzs8xvxmUsmj0GDQrkpV8NW9wPq
gUBwiWwQRUmWgC9ws+/95afSLG2gvcV8UuC2KNI6Xwxrrtwi2fdVayUXE/YCIKsyAtp+OZn79UpI
Az8NUFg6G3pw09MJEH9g7r8+mUxIBJDXr1a1tlFWN6xILdFdWAEFFyysDnbHuR4rd8qSpyTvNlZa
Lw+WFszHztYKI/iI/mUCH+K66blsAf8p5OJaATlB/UJ/y8zfYQrvxFkQue5yG/btjG8PtEbEtqsc
kNPt+xfJODwUcHCdF+J1+IdZaAnBgkVFj9xS/9WjEcRU2jLCEZjCnV5qfmDNtgYt3Ky79iQSIcNC
5UtBylz3aBCjvq5S0XGfqoQOkJItPsIYkYSrhwZkwledxCiVPaD/NnaCcwYKD8TNkXVIueyvsj0f
tncu2QqoD+301w+HYt7ZqGJlcIm1WjhiuI39nx1Qh0hadprX1EdOe9U1heTezZA7tuw//tlnLSq/
U8i1U/FE43J/xsi9HCHrkIiEj6TP6gcsO/bten0OsO5CamzKHFKmp3Uq5dK4c8Y1AOmkfCDS099x
Bj4W4hQLO3WaVenC+N7S39GpHdhtSUr9XBIsMPzzJsFeGLKb2LEQ35Ebc8ahbxniiDJG3jgjNImH
vzV2MPTRy7tO03Cv4yq/qD7EeHhabZt3nVqhWpmly7nAl9S/klX5MNpSFoHYt4391TQ/RSNRUOBc
zCOGZ2C2FMedDEJ08lJHepPGL53W5ShW3SRzD+6/zRLpPF6Y1GpgX5o4+H4nodz8CEC48NePlZn+
6R2trmL4d7jmL9kkvhGwe0JQCmuNWaFGyNeGGfWDSDPvwC8MU6rk2AGrelgROkiGVXjEiHQ3/VW6
Un92I3b6XAjDz8XzO98Ga4OwCPYzxdRQmIrKvdXqnSf0c07H0yE1vBlaRRUo6fE0VUuW0VqBCLu8
4DVlX8DJt+VUFWsf07fwWjb34uHEGXOLmgOxSDzVdp7NSsLWGyqr9kBqT+ACznKHqHbinQhfcjrc
8LMEGOhbzBg6W4oJq1tKMOClpTR//tu8H7DtNGpZxQp6dbPS4c6IRONGR+QReM2o3RF2WhcDn+cu
0m80Zo9ywzxgwMCCxNSbn6HVVxNuD3HRAd2XasVcebeaWi7LG/0A6B8Jl7dOK24J/9UefRt1wUXV
pEkVuFpInuOvkUTX0kEBKTaVqqRaD5fveMxy8wEbk9eDbkOsijlAziGrczrIZHGuH+/RyANwbkup
UOmlHs2oQS5YU47+T2VH/T1aYXhHLLaJVFSd7SxMkfc7X1E0mfXfjzk+kMsDJr1vgXKfR527a/Nw
9XetRUV/4J/2fbLEvSLCf8GN8/EkU23fwT+UvpDY5hgji3lfJXt8bDBdiwtIEljsjz2SIcNiPqL2
V628cOKqZHHFMMqiHK7blnyW4adICESgBxO8eCRlp6lF2VHDMP3DD1NjktEsjkfeyp8Y3MLVfg25
PvqlCARmsLZ4YiYORwodgt+kUdYqEDR17jXQT9ITSTvy4LNCENRIKUze9zckTqEAKX/n1jECBm/8
GrraEH/EBXYbCdGchhaiff/xZpwdog9v9MVgnSyphWNCAiNgapviQVth/z0XEZEh9YpxzFaiodL0
vxJ9pwr/S++n7AzG+nFodiZ8i5zRW00aiXTpsB71G3vE9NO3F7hpyGdlaWjf8aTufjSCnpexxIBc
60A5fjT3dSoUDS7zQ3CzsHGetaMxd9zdJqstffrGB943snvcGkNR9dNPrRtKZ0tveyKYNpn6PSzC
8ikp9qXOCS1RmtrugAQgu86PMNmkm72iK+JFI2XyxqQxQG3GrIbsnG1689fV5xcjQnbdMOhBJPC/
HKLY8Xxk6Jc5iRg7TnW2EKCd9De4Aq4gqJruD+sGvh3mAMFSwGqOlBJ0JUHN0Kp0d4deeWPz6ZVX
PIY4oyrNTfbGgLdbuz7QtkrxzUW79WbPTrNaoQpHY3ZVWTOHSOn73VNJNZmelUEHZhPe6PiGCpbS
P+y67xQx1x8CkHp1cO1+VECARgjR/Yjl/tyyc5YjK21YMfRZRgNgJy3PKdA8fEh9JVT9Aluf4+NB
7Yp0AOiLlQTFDRW12Jort3asIAnA64YP8OYgdSkNDnhA2/aTx7m0PpiaDEu+xJRI3uW9BY5P0ujP
KDEZ3jSFjtFs60yVQtj9x4OFhXtpOcI0GVlq1O5bYfh4bb6aXK+27jj0DAQMuSUs+rK+jGsVrBaR
7x9qyjtNEzbcQ6jnTJKzHdaQvWk4jCSy7Qgldy4nBmgJrws0HjxDL+RM5fQpPaLQmmjz5YXvzL5+
I1yyoxj30Gi9EhDa49G7xHrJ8IK0V27fmWoy+0pIorOgb/TDVNruW3MmnKrud2u9A5drimSXg4qJ
oyf8QElQr6HEpg0nGPapN8u6IDV+BwY6W9KhZiW1bTFt5xOwF6K7017IlQNSy53bjpDgguVjp56t
ZB18UTdubAzI6FkLMMNtkJBSnq9mmIOYAJ7qKHgR8WoH58qzKUuNom6Thxr/upTIhQP0ybGQD+0z
r8i0umZ5wDmNIR7L9q4WmF4EPePEO13yg97GGYo8oOomo5NHXU09eUEMJYrrMLQxProVrFPzbLZw
tjk+bkE88Do8q7aTKlqntjH7qZVJlPXW1qtiXYFyfgemOnfEqTOrBQQZnt9m95ZnhoNuzxvhIHns
9PESekieDkxY6GrxIl2/bZSp6TjcMCDm6sQilEA/ivH/cOAx+WqxaMPD/ja0dSr9NqBgOdGUlyI/
BGHQnng/VTkL3Konb/a2I8TepexsqTC+7NE5SRPKMmv93DpkQPFNT27NFT6uRo2+4/BFBZWnO0yF
gAGoe6z3TjAK6rVYjNj+tqxOAkJlUSq0MxF16O8PBWuzVCup48MqP2Ub06UX8D65IOw18Islxqj3
PPnjAFIBemQ1TvEpATRfmohflxTUTVMz64vL0814kdGtQttsxqPmnM2slyRZVKtuTFju06DoZTex
O163Y00oLj6R64iGEM1ZCyq7g6bKMk/KQ/7RBJrmH8vDy5HoImFZYBe8f0V7f9ziroIUfgiyPzOu
ex519mVdXwZl7i8lkCXsfcUE0vlQOY962serrXUqknHpBujnr56VwuoPCOyukWq+8MKVDdx04bHu
aMIsM7gRWv7vN5ihpi6/NISkJvnl4MZfsOrPyJTxlFbUu12rZU99LRWt6SCRBsXOUjegPeR5ESKZ
8tzxxPauLAlYB2MMj/jtzmtzcGvf14IzPGlRl9H6wu8gHnFRLffvZQPtBPtDQ/DS0FRYYasNcbTY
ch+MZ0A8Mn0A76rGQrUvk9N/6+Z5co7A5ikfjZBjrGCR7QQoT6gMkTpBX3oKWU+GUOn/W6xSRXhI
tAkpEG/WTXiCgs/sIFsPfC8tvjd8ARvAAE/A7umnSY1/VO6Anwn5c0WeCuL1Wo1pGssproZ8mlvC
pKBMhjKtkCQUNqnM18EgIggqfFOpbtq7uKQkRW865BblUSf2xNiZKIbxR/iP+4cDaAcCUqOeq7fO
5JtmcO2AZ6cQhj8Sv04Vqe7Vs3A5uEE5PIETLso+bajLjp07rOyHk3DwIT+Qn2M0xzyXxZNbHS/K
YnUol1Qn4ATEkjPi0VT6Kx/I1xZPAyS6Yq5baiOwAMmMKNk0ME7Seo+i3XtbUIvkVHtjmw7+8jHn
9gdGk+krCdxVf36WM9EROuW1lqLeVmJz5tiW+2on9HtJa83ZknzbuUEjYkVWZtPZUUpco0F6khgj
w0mQg39lTgnccOwbRfFwrWjmzQyZ6DNKizkLX+Gw5ZPx59FJEvCtPtw/n5O0wHlraNoNtbxIFDg6
r+TAZODAo83+2cp0berz6hj7zlKuvSYdvORqwWC1Rr7r/6HM+DuIncEc/M1TsZNlc/VeB0qi77hU
9wFiKk2LndC4sX3y6x9b3G8OQPK/pHI+F+PQLRlOy3FWEZGXfnAaTxUsEvhBVIE66w03MnTOx7Y1
WynFqC9j4XiTm5hviXmXNLX2nk6iWNOnQpjcyDlX5GvQQotAQ9Uo7Ops1vtIoK55D2jIJyEW79Cb
mK1IkPQAch15G7DsjuagtQBJULV0xNzBQajMC9oiG0+vUgwDsuY6/Gj/lmcX39DK568n0WCWVx5t
Yw1mECYAVw78UqGfDbZWe6g6NUzowyJIrVLIPN4+x3L3gI4/IVFnC1mQSCEx3mbFpxdKZTdYMYE5
tHcOeyMCh0DpUfc+iSsEHXpfxKlRg/38pWmgiyDgum+usEgf+MdildAjLgURtvGpIqGY7JYVGVCr
8mwCIfqVy5M2gfhqhYuUiAZQqGhekyiXs4TTavKV6z2anGl6dimtoHVo0PjODrUBuxCJ6Rl/UKmD
KM+huYQxLkJflxCDZZ5JRMWxBVw1FMMrQqYMNUbKuTOkVhn0JCaXQ5ZN6nRjkpFZ27aegSxQN0YD
hn/CPLGERKDpKZ0iFc0jjtvmHf98EUnirgbCULgp/AKgh0cYA6vb2ezqfI6Peb2mEo4/tso0M5z0
Ts3hBtGqQ95eQycdr+PWgYQDPBoJNEznVWmQMIc8t3CCL9YMTEWbaQV5nFfrL44vbN/nZSGMDWVJ
5Phfho/DeViJXjDg5GWxDltzUwQ4ta/K0Bv/NRSYws7IbGLbV6QXwdv4q3FcZ2mCot24F7168ms/
HNS20J+hfVM1tkqCrKuDCgKB4xpIT4UT7fMWeRsT9NJSkM7kJvxU18OZXdr0vdLr6tjNbjO+SQ71
ckspNBWKh4TZVwW+nrkZWTT3opkffo3glK9iu50LJhteHGe73qJDISS6O5UtdyOHdpVcL+3z7bAs
qMUjCFmDq0SyZuCR6Deyrjutpacv2zkOpZVLKlueEz/eg1uSukTiffTcPrNjfLRxk1OP89es8Ala
JT2XlFqUz7I8hp1kDHkoFx0x5XPn6cCVuzJUTM2Gc+xMLABPrXGGls1+7N1Dtur7s7Evy3c4rMEw
KkdjGNtbpaVWuu1GlOLJd47sBRnUuo93og01VgRWzaxRUUGHi9qDmu38kzylcA/oklBBSMYmsRpi
cZaZ5zxn0lt8bnwCnIurjT0UHmdT/UUTSyMpawmO/eG/VmrI7dUOWNNp4Yu2PY3nLeCvDdCKe6As
JWhTOFzgbQWNtaDb8PG/yy6ysRoP2TkiShxxyjnjrl0mp/WO7pEp62igkUkSTOIKHKqGt8eiEULS
kMghoJds3Tw9775eRLKPTS95ngmW16wc1oTqZBiiuJC3bGk1Q21czSIYSJCJKqE6ANIWgbUiDCOZ
FkN+PcY89UVlhu5pf9e8Gw9jeeXDK/4mRREGhgUHEzeIl/6IDpZAn97iGMBA+AlFxZvGWYnfXAy/
3KpQ9inqerlQtIzJZbyMrm3qPOy6vNxsCjN8hZQYwgqGxk2Mllns76q45oh3r+zSGLsifMcLPytD
4FR+/a5A5e7XqcUI4sWD8rk0PZCu3J9tgADo/ZrA5vSAK9/xPFSLELBrQrcSK88Y7kBRslpvnjW1
ai6/Mys722cCLdxKKKSy3p+2bknSWCjslEve00Oa3uEcJWJXbZREzZf4aE7LpT2cFQPoCWn5UXKC
sB7KAjgy2ezOf+HZIrGfPCNiGo+6kjfnw2pDIlS0CwshazPZaPkKn1nNdyN/B4DKZkRXb4P0BTOV
2aEv/gWoTkNBlTaIDu+pH8vlZG5eJ8A2B+DMqshiFMIkWPgU3JKeIFxDVcRrsYI+Y5mMjCL8A5mO
tRjupHi2Cu0HQU6lCBzRMdHGsAjMrvNdLPmZwb7Wlfobs1QxXINWd7T9TkRMxRUdR80Flb6JisnA
9NRVXbJNgeDwCfVA51GHqCc49x8h9Bp8okNvR2Ysbu0ARk5MBFC+Uz8YtXPo3V6Kz8RIiqYR4Rxj
neRivHpkLp05pVaaAEyPUcCQ5USVuqSkrqq6c2wgARwdCeHuEre+6dJ/RuFkbHI55FhDlM3hOTv+
aqBKUdFUHuutKK/1fnCtGyb1UZvC+4Jvs6O0GMQ2uaOVy7ETKPBkaFl+MVdoVGNYzasvH/q9eUmf
unj6H0uL8k8wcHjMVxaUejYPtZZPjaddYdoo01+6/r8kcadILZ3CfHpYBuPALOUCXaye7KE1SoWN
qaqghBjY7TeM/GZUbVAKbj+LQNy7javRADgy63eVk8OMoCl5CBjMZdllS6nx8jJLZ80kMhhheFc5
3wny52D/7Rzvz3+NgRlAkp7eDjDD6muQ2tFxEx7ZPxogBalVpC9YRCUAfmTOXkBdci1ZRa8q+VQF
qRIjSaCcoivamZ2b310gZNLUysU585jLkB6W56m8APoIXBAO5ONZ7YXpWpJlrzjapCfSELiIBN3u
tBKOt6WJcvryBcOVwW0wJLoCaUa84sT0zyxDdkhQYgpmzKlQniTZoSud3EX6XhzhP9QafQV2Thtn
88QzQ6ynTJ4+UhGIBnkfb0/QpXNPmeqmHPKyTSzFEDY6XE9ZqXL2IyWndIE2NNvqVSZvCm4/Ugq8
OYCXJirEzCTooNhbO5fgjH0opkvRlei5CKjuVXYZJBzKejmj7RCR5MSgFdzeYpyxegmweZuZ7yBE
/sLcmiUOFPBRt3E3+skXPZuZhLcERdNoVwEyXMbClTbheQwC0+6YXGtWfNH7eUoRPx6HXp2Ys0oW
FF5p9oTqVI/W2WMcLajo/AF+rsXMdUExl5HNax/4Jckfe3KaM3FTAq0BAVfC2MCgaJkKTx3eZSFA
DZbD5g2rFHkPLhWIa8HSodiuzKDkrrrlR0hJCMASgIcfNIZ2REdc3e2eADtnmH19s/DxdWNE4Mxt
i60gzxdA/mnVPzYpqOHCRhWQbyeChyuWDCPmUD8sIZHS7nxXA17i2CCgQxzYxLPyOAyLm60Ufyex
Lcv8AiWCvruPWcLw5Flv0HNPcNpcfi/kR2mAx9AIxCgJs2rpLF4IdrVOZEtrppW7rKIExbIFz7tX
BmyPLcJ8wZF1QGpBjEdipqMeEABNWDuKLqhEzYeduxnaQel/6TpwLX8kbh2fEnRmzM+9OPQIVQzY
kY+FMQqlV5Y9jIYgjMLrXvb4IdINfO3u0K7c8w0+JpQbotS/iPd7Bad5pA9oR7XYBzS6sSfvoQKl
VRAxNbEbmiSeDbuuvcmFocD2VplLXim7wXU8rlvbD/7UVERpvVKKOUIuYPcYKFradbwoOpZeQzzp
mQrrB+N67fGJKDRCFBpDVIdK++IR8DyIbRNNjfLtidfhlvLFhWZMj3kFo6TGDulCpMIAvcIX+HwN
DFMRclFmHw/z+PXbzT9RIglFrkAOGvS/lp95kPehYM3gAL1Lvs7MlnYsRyO0BGCfB1mnJEJx1JzY
LpCwlC03jMjoZrQBeRdDAAQ4hHq/bw6f6ebv92sMUuOMQnnNkVfTIKAD6aFJzRRCYRep4zLjhMGV
IXQJlkw/SoxjkhIOJvSZSoVWpVAiS3rdHUx3xmAieY+p+w4Ofn2Kt7NDbiG5PJYN/GeKZBlacEZg
GfHlJLLm2gGRU/qUri/S3DpjkuSZOZLrft7wY/v9mHQTjv1fn37ZL2aUg8Uc4wL2ht19wAknnhJ9
3D2F4wcCxtX0eKLEgydAYMkXiw52zMyGlVLCbcGoFxJGD2UXujG5ydPjr47HcSHKQAP89Cabb9Wr
VkmhYkX2WZcZ5HPSmcfPnUPk/cjedM0NbaqcqqLsyrXy2DJCnKJIMCrPrm8u7/Lp+1Eptev5yWdl
s9QbonYhDml36NPhJz5xwVFSXp7lYs2WPkgofp8rieCqEao23QCv9KNWgINN8N0FJhFVuj2c3ja/
Zzjtamv9bvijD4ng1m+Qc4ek+huaJn+Nyd6VbfbEqfO/jV/wQAO71KBWCE8a79OQNefR/L6a93tV
j7K/kEpReK8BHg5ZW9Ph7PSpdfgUwUZlYYdHp45D4Zagn0X1CQ45wlpx9yF22Q7zO0kRXcgcJsGW
ScW1CY2RSIgGtOoj5VuCH3ht6nFg5Mx6ZOnb/578WR8MONDH8BMvXSPGnVn017txc27XdqY4VNvB
gTv3JlILCSw1RwURuy58zRXxdvG1+k5QbUTd6h2wvCONFpCye69hWsyYAxOyoLOKXRvds/OMSCku
xLALYvGgJ50Lolz/dwzfJxVJS7H4z+vtnaLKzuxyiZNtKRkzOMCv44uutRk4k87cVaYRb/lBZHSp
L5uakilsKJjhS2MxKMXCfJrLehGaDPHtFohXOBqmH+cMjaCuPa2W2fZsdKXDnWnmRU4A90+fCMqM
zbfH7EJmkr5mekpwyiL820SWIO4z9BUOthik6Xa95bdoWXDxVB2n93fqkXtZ24x4EUEzS0ORWINn
uF9feVlYxymsCr1/iv0oF01TUItdLtFFKoYJzi/nW61+SejtgQevT1UqBsCV+T5UvQuJ5Cr/ZfLa
I36IaFF5wLcvSr5xvJDJt8vVB1TcZFTBHAjTvWP3ibRqOFncfsC9zz0sk/2KsaQ6THyckx2bb+bm
8NGnYzVCSrL1EN6S0cmgeC94BgMteypDzT+WK5fnCdn4WiAR7CGaYtVpxFo7+RVetfCzeRfsvlOQ
vGTHAnk5oylYekRsN8wHFAbsvuVRmtseF49w/xqyBXiEqG2eLesTog2z2f0JS++n+0giaIaavn6L
bNGky4HclcwbtHPhCY8fBajQ+LTK7qIh5qSdlCJZueHrCCsrf3pYGvqQoCVD29lA9IEK4dxvLnd4
a0dlkTT2Xz1eoRVk3MiVDpeHnEkL9fKNf7iOj83ymsvQHIteZ7LMsRtHY3ockVBwHmhl+XpnKj2L
NUoshFM7hJzHhbfSThv8FzyAG3NimcrhEhBr/bIPvyl5ikMDyD0U/yuBfOIohZiBjRfDa5oHYVtE
0QM9GajqeHCORSLjeuAeczlhgFFymUD/qlxkfG1H+Imy1RFwC6J+wqFVOXd0XsdhdsAJ+21lMudC
43OWvhK3Y4LdpnStHjGCnWxFwgy9vni7ukadyTkbUdynvVZKzTX2VxKpJAjztaRXOq4ttAhv0Cn3
PwVd3+dgQprMyobAXcuni9/3andq4UJMPSPEPvaDs84aMv/1SNGkkjmJ4i8LTrOgOevr3oJf9UoZ
4Fgbujcrm6UYAGuCfJD6aGBPZAKl+fbp77y+W/GSYiIsNh5qxPApKv2NTyBt8afcWVT7rbjKshbY
242yEBbIxPea9warax8TAYvorQ0nxYCxv8UB9SMxIdnpKY4lKio7LAKe65BTfLDvcbAwA+ouGx7M
NUuR+hNYc5Uq95ynICQQLnDmzwZDuLE2O4QgWRj8bV3kZwQ2kwK8FKsqkd9M8GdSCrkgu6z99U9c
TUV0msdVuOz4tzQN7EYA+QQZUvvw5enLxb2WFREvkrryBeufuHF8CV3a3Ry+Kzo7fu1qh6fqJNZg
H4hB2DtXHqdhBqIsM2jvcSvzBr7ONEPx62ia4YEjNsovFLIrn9lHHhbEnYUcyugcoG6RCywixlzP
+WotonrSaJ4eEyFxL+o5tYyf3paDD1KM7u6x3Yyh/rBr66CPy401bxqcgs8pLWS8KKFN+5oJUW3c
grQ905INrQC+bA9yjMsXAzRKClizg+NsNQvR5twt1CoO2jv7mChzIY9XLdiQf0+YuIvuG3jOTWS8
yrf/FKzhMQ/Z8dslSjMNksWLvfs5/Fm5y8BHKd7mMlU3ORD4Lyx+LU6cfK1r0Yn94xa8e30L07zL
m28M/2yOXUU6GdWBwfysdwhywBSk9NTnIYxxEPf1YOuqK06SfqRg+L8ozaJ2FtaNET8Czu9zgdaJ
lwxgy1LS4a/wKahUkiy01R7tQs6p1Adn+K9ZDidjx7bHbo6qEGHEncWnj4We23yDECiGa/nvXytn
iZ0Wht26hPesS6b7RLgmg28Wp+6tIu2bOc7eDkk6wUwJ89lTwwAUL4kstKXXqbcDj23EwqhrkPuH
Q5pcpOK3UbjlV/BP9x3I8NXin+CZLW3nQvVQrk/yDyw0HXwspakLuB0g/pN+qg0l8MDZ6hx4iljU
jM6RJgllJCTtoOGKhZvjf9pqDAECvLGHPWXWVhnv834I/ilE+cI1nhI/HFp2tvtRM5ar74unuVW8
CkfgbLD8p62sTsstttadIQhqRzZh51I05IWOZzvRv26m4nOsa85VBMVikZe1oB6CGyLnh+HN6p2F
DQV63KsNMv7yIB+OT4gzssJ3BZrpUKMDKA01x+fH3yYiZBYMY7xPAoCZp7QMqXZ70CBSILny8toc
tD8pa1zybxMi3bbZ3/ZPv6+zjbHSgkt1yVPWprxCtacfdzoIyDqzP00kA9aoCqav/U/dE4TtYp4s
0wKZdpZfbA5SYYv5p96Bko10PDa9wGafMVQt7YBToO57zcfkDa2Jk+csNDXvk0ZJalZJmDXqtEtD
NiE/I3SE2BizH5Tf5Igbdl+jWGXO1o7uyZNEkmy1i25GgtU96Pmd9VlcR7h+57PFKtt19O0Y2rMt
tWq5UV3/PRBFZD+tJqUuim9u43c37dR+RW+M1Cd8kGiDiuPnK66Zn8LB7hrpzFW+EXp+Hpj2y2j+
gRiOphXH9wVTkpR/4YWQGu3E6JMwdsE3qpegvIDgMsV65WGkLGVCa4qGNxmTMQx3y4XrJcR/rR2N
Q6D8PvygNxFsMKxxjR/lFqd9bpGIENJJff2i0BT4Fws2Ema0Bl2ct0IsN4CgcZkfzalwCbtejcQM
6plaEcdStDQMYBYbxWTPFueQpB/rsjtg78tGq7Jqy9oILDnes1Z0AFGf4tCA+qtXnohY4gMWg506
GghM2z5B5T0Y2xRSMWNtCSwEjIxEAAma5tNxsx3NSlP4KkGVGdIyC+YaHAO3m+vMf6XrKkRk/eOv
79iLVVUbPHMhi9DDlx0vaWBh83YQyVzHO9WwfzwlJbELq4xli+1kar5mfX7fUWG8bCl6LHW2cuOU
7GkO0SwAlTOUR29hf2X042xT+DTQcIhBp3Cx7KQMyDLIRiN/SC5Dpf0UxgCdQGWguzZL2w5ihugZ
g/+b9IGWVvrzLFtz0mc1zCs+U4CIi7KzpAiJxki701gOfQ+O9yj7rquCSEdQEcBXECyaht3NtqMk
wCLG9osdDU/6AgJs3wl8jPq0cCRrGaSzpZwQXd3uiqNzoss2bV2Y6VAVV581Z2S/rOPjGdi8/mTb
1fODr/aHDfDmEDZMPKrErtQI5NF4wOXh2aoIUXJ9e67WNxYe4N5TDvfkuNiV2qurgPNiC9RIWpYG
4QKLOvgvrQoTP2gA6Do3HNqnW0chtw7V5+/Zv9PvYcWIzh2yA4Nldn846/QGQhKzEM2yrMbhvu4j
oCo0IqU0GDwz69aiDd7LhOuxLGIW/v6N3Ntx1La/JBL2hRzcUww/E/m18vX2y/dinh7ptjQCyPe6
2JRa7+TzW+LzkUuRU2C+eIPZ8Dh54mTD6H0k5i3BhmNJMi6G7Qo0mNk1RXJhpNFWtgfkyBfXQ9oK
dfvDZdfhH/U0IKdbKqlUwLwnP9gEvZpcoQhn7pbphNqzxN1RHEyiiR/dYFRcbt6CxMtgzjg17Xaj
EY+rkrvcSzqLz6SLm+J8APDHOTHzxamTW09ETfXXHiaf77riCSIfTqR2IiXHywADI1cFmZMyKfwB
3igHTSjSavMa7WOCZftA4JKykj/yX/YFjLP5T3XPxeZsHwO67Qp5K5IeCekvq9dZhY6LnxP4AFjV
YdP9Rku+Oc1oCeXW5RI3l3RL2/L15t9QbzSS62EMRmni1lxbv/rAC46hqtV8U6h8bVb4ePDymyOJ
xCyilJcN64FUn5cntDy3oM06SPymRiMH2Gk8GZ3dggMCJKTSgiTba7fU6HPJu9X2sJq++/bpok2s
JJUKo3I4bX3Rkf1/6zCDK6E0SjMv56+ALsLumVOwP7c5WEEz0BRwTMNwAErDg+bN/n3NjewcONU5
pDatfYJVOTZHJK1J1PUzUesEt7JlHPSbzYOPO1reJdArtRIlOIz1PQqURXiJ2Z6JBYRmYfFt8DI6
TU3FcvHOC8+/lFiFZRp/eIwcpitLA8xBl9hKtJ9JpLEAsh1k6FcW3ulTsquYriFxyDvAnSo5SPDn
Gxn39prFfSd+NJ2myfk5284B25ioGbt3FxFFMte5q8CH5klk8ljmfLmGI82l2FrvsUtx+sGIX4Ga
DqAks5U25ZhK8dbaln/ChgWK6BfehXtO4ZmeRAIFcrL0vFEZitswl2EZRIvlEWx43f85iIA/JB48
CFKHJ011keS5MExjbpECyzzfOdQg5jlfQd9hsRxmI4G/2XcfdAuSDoqmmSDTyEZ+II2606KHkUf4
j6rCihbcDvZ6ioeQmnlEEKEuY/U/+7LizIb/AMmZRHBYFBXSrmbofz6jEXJL6NxLCnv1IEpQ6opN
24ztbUe0IWytplO8/NcabwD3mWLJqyg7GqP4VGnz5OQXtVaOVc+JZrDcCwF9gBXlgbo3ISKYohEd
Y6qAQ7SJq3ED64j+TXaPdGM9g0XnrYcEo0eF/gYy2BxVuU04BLeTD4WCLeGYewsfvmvJQ056Axzj
QCrB9zhY3Vq2Yi/yvWCthmPU3JjwBLlJh453y1aaqtupdqHvwSKnFjkhQcN+c3OTbFQ30YFrnD/n
f8b0R6PG+n8Xeh8ugVH9rRrduyEW/oBXrvcJPBPqlklo0EhziifW7upjI0+tQPFVunWodHsYyfmg
7tgTjdRUXnhfYKKFVLpBGRqZIIOkZvONOC4a9TEzCqe7kl6xG8Wp8OeaS/pXEOXiRyQeOIhoZ5Ni
rCaqxnUmTbqpMKWB94Ew2eSfOw2qqp4q8r/mssR3IenkMp6yZRNevObNVRU/OAaNKbjW5OLBSS7M
L+3DyZXg9vRwrbasdcB07red7fd/cP2/BCJAm7BkbeYzeEQcz0reZ3Bqokw86MC5awOHHCIU4uAH
lTDlQaeJ9kL4v3zT+zojFj0CUjOiGLr3tHOC7mgCgQIYkx+Xb10awMqvHZ3hLtd4CYjAQxNbHXp0
oeOG7z8mPmf1y8UEzCe2qU4xceGnOCdQXT688T8lDaqPy20RwLKOg/yunSx3hFty0ddvSA8x6uw1
Pp82GyG6nHkfTK8Gl9gwPd5MeQJxYhHd0JR/yeuczdM0AFNK0bu3CdPtQEjcMMRLgLaW3YQ+5pcy
56vAGjZW/zBHPOmSmoykGzQCgvcxP1WP85jG5Xk4f7MWOR7V5PoSoWlFjrPsYwzjvtX28kARGVVC
Stb51rF9xGIVDDqc4XmI/cidlfXr7QR5/mOzVDblSxisY0M5iOMU+m4d+J5UbixEX5yF0BVcSLGs
IEhaANVcAkZCNm7BiHwL6bM6taXUEDCdYmTcPQU8VLv1+k79nZX8x1QCw/rfv3ojvM5l/xx52bmy
igK0M6VrjtQfJAEUY+jpnkzWDRGZCADxDJVXPRcpgT9euApMSx1P7ADisZevJFkhY4iT3ywtW+m6
msJYkq4QoV/2l5Iykf7uzkzHyHztRswHmoNwFmYjmDNedHI28NxJhEcbuncWl1rbl6ldwgr9Dm6w
iqZgvoFbkhy8s9j0E092ehSvaKMwNzMJqihphsMAsUBdotHcVRdUHvAC/uOEEyVksF+HtFjjzCtf
yt/Jhieg/AKNmkV1NEJNlAmbOobeXsG5P0CxeCcb6We33ZL8w14z8eoN6uoeeUNww0/t/wtMfEYU
JiZI/qYAf3pXDYE6q493XhA6c8nvQy/nJEACq6GqTTI32R800E0YK68F48hcFVaDyytrqPUqKvl1
w2pnRNKGfTCae5PG2OrMfQzWS/3AfNXJQDSbbheBPFyqaoGm0R4EqiMMGnUrAAyeLYT9uVFTJNtZ
i8fV25593O4TL/mf6Zk9wiBSxLVh4Atb4eh0uGD6sBsNy51Umhc2a5z1OuxSIeocJHXsJx0wOdSX
CWX/lGPAX7wYrwYVx9t4UcuhSeNlNX1PnkjUqOiiAyJW4DmYX9dd+juWP8v7q2QbSNHrudsRm0jo
zjskvFKzZr0TnmEBqJSSDJr1Mi575N+nFj/UzRhWUGb4hgAOBTWyXsmAsy+lm8BmM0ADdD45eODK
6hayKvUg7dIU4RybyO/wYr2Nbu/QhCDrJHc90tbOjFmL3udMlm810mmG2vs+NQi6Tdz/nWhYz3ai
hkCnpc35wRv4TGUJTxEpD/zuYuJAKrsfCoaOKFhUiEDSuxtx8tNlOg1OUBocCsUsYRIkXZ457d4E
qd6cgbTqgE09+t1waO2BKUbyk18SUyD8aN5IxOkI3C4Lajphp8hdLA4AnYlgxJglq8N2UcNVxPmG
4ITsU+ugixQj9mGozSWktkf0B4UZHo7TvwB3VLZvRUjIVyZwul6bMawU1UVLtg2aMs7ZjBLWySHx
ZXvljwr4bmJGJB8Mk0W2dYaAVYc0EpqwpGsRHgIrdKcWIys7H5JyoZLWu8RJ6thX09ezwtzve1Ht
IdpLByyaoAHkPwMax1OMDa5XisIVvwnphdSNLO8hqao1p5eApz+khpsIbWZ8V3TeuWcOBy67SIvR
4jp6SH4XOEZTPGhTRtTbP0s3hAJvhmPexojwJBRWlNgr8WBFvrL6tmq7QMFIvJqcTVoVMe6/9uZn
KAvizwtyEZqLtXm8Cf0WbpvVL8NqwP0nL71VFPFEuzOo4+Dv/R4FszFh6iy89eqCW05MPORdwLyB
WBhIWC+HXnQshtQwxofQqGGTE70sZ+fzs6hWvTZjHuseTXf0FQaMvvtHt684cbyWw9ZT9VSp80Xz
jl8tAmT6pwWLKRepgFsIPRaSI7/ZRz8yvQr++Gu48jK+nBsbo2Zjwc99ymXsTyIfvSnHEdbfdrOJ
g+iJJXnv4kwgems2e94t5X/7UXK2RM3JCtHUYXougldWspXEkUf+g50LaFU8HshDUI32NKLbCnmW
AltqOMQYtns4YsUZtndg6xD5NzW5AJhw+V51vok3g8aNGZe4IUNmYpA640th2MWWSevYuUoZbij+
qXd8za1yOYIKhSkW4ILa1/qiZ+2yai/zINvQQYoU9UBIrKXoNwszERz/ww78rk56nhQXphsfqZOK
ecFrDz9XAlG2hy1Txq8xMFMNrgkcHdwb9uxxFullCOyWm3idAp76dXaoFKcrbcghu3CrnafejRv1
uAxA0s9nQnmvmt9Xk4Sq8gFpnfQUHJePv9gBQv2u9NFwl3Xv0YEnHTpOwzCcQR2pdHr+bFrUhXof
pTLyVUhDO7dkQ9eiU/QwDH6PdNIT65s0oK/q61V2esQnKD8SZqSuuF+/tLqENWI6Wst+RC4R49G9
GLFxiDSYxFAc8F+FnAuNyZBGbjFYPCuSOeDrdeOt7zR382jzkDssz44zj1rRjiiWp+7SX117Cs98
DEv3yqpudkvERkctuAlPrNkCEWuTsjzl8WwbXVuhn9m3H+3hMfdQ/GoUyTpnZOj05hwqDK9XQbiK
wNcgsoPWXuTu3G7Dj+w1p6UfT5GcwEWGu2hfPDlkcA9q51NB7cyPUkuywRbJREjijhd6c0ZalxDX
do95zDFEmnfJ3woLG/8vRRwFXKXoBe5gAryuTXThYn6e5wIJhzRqGZ/POvivKzV989e60X9pxbdv
AP43BvEvjRKaQL+DpX0jJohjxe7VrS4es3xXMWvt18qDLXniLdaq/UB2wzmacauZOuLn4rvmZUi6
AAvnfd332AgXAXzSjk4cxz44bbNhdhBH/s7hRapqr0TaRfZ2RSUZNcMCy/YUD+AY+a/U18+ZSu1/
2DZeNkYnby94X3bK/W844xUD8ktn6tPC9Qe0JFJPZIKUI4N/fc3r+BZhh8uRut+e4FHw3duGKuOU
fgL8lTrKQD/Yngqm9ciMx5R2QdW/lvzL0GdTeuDm0a88dOXEo3cB8OcJZycT0W+Fua5Zn67Ickoy
egA2Acq39mdGUupscyRvrPNJG52YKZVnfgByg/rmh2fPhyvRNFaIJac/yTbJsQJEg57Ffwdht0gZ
OWDcH63QtX+JKqLa33lgEITlPeJsCWziiUCX9+aNQf/bpYXipyb8RQ2z/nq/6IxEMU3/AXmAN5V5
0hzfsz6eRnGpyuqkxCZ4xLj5ms7HqFXEd1K1zOBTRFdboHlpE2n/SNKkfflTIwd5A2G9nqsazc7P
r2K1TqXxiJuAYPAdDorx5/o7YUJFA6Tfud3HxSlf9qOHAS81ZJlehiFRpWrV1tTAPaTn3VVFESon
N8s8DLf2qgrg+I++SeWQpB8kFzwrnSsWIOI0g9fDW3zpz/W/26jDzDA7yJxAEtf6pd9RpSLzO4TV
EUHVGkfJsRcq99BSp0YYEFH2Ag/WoUWWsL9uVm4EYPrE4orObazKjwhZUh4YIMh59t4ulGmXIHlZ
NjzA3Il0/uxycsliJOQaHhfD/eA+Qm5pHTvp26Gkny2x6yMo0+eM2xn7U84e/4hHlq5ZtMrCSMl8
xnx0bdx7UFeb1SWlMhfn51kZ8YiuLNuR3W2cz7neq4qsun+Z/wIXGABXFjQQTopLvl7laKpy9M+i
mTSpNFSFIL9pxaj9TvkLgSghVTogqqnO5a2jxme7sJ+XH4ruP1Ic39pcwQNs/cpKAy48ZJQIKdxS
W8UP2x4MJB58kSy9kCdAz0l0/1FTRdr4XPWqMMyLqVuSVaQZjE4GBA/DwRlaUjKxMzcHFopxXXOS
i4cKn/Isf/mYoTp3bymKTTATFYLf0qJKzqMgXr8chDhOzXI4owV3oiOgAs8G2mauJupbwwzf7JBc
M/brQjjnSl2gUZRZuRkRgl7mWg1FoBcCe9zsVuZCS2HOLu9J12NjgD7nm+KbedrXQDj8Is8XkT/M
9j8e9ERUBfVgo1YNLf0k/6LS2S1qIYTV1iOnrbYWzyXVpOw1K90VO0Ghpf/1ScWD6peGQWoXR3HZ
PoZtW++39tTymRfKLOqiyJuGQSxXlImlHYrIUILqkNI+7wfzGinYVOmgqrOwb6Zw6eRQRsKob42B
rqrwhrWUc04HiqvTMk+rVnzXpNWP7orPdR7Q5ZaC2YvFQFL+TuTIpTOLcuxtkrPOLzVplVoYr+ok
xSJ131CL0WVNl3aMjaSfageDk1AeJgfCCEZaOHSvFZZ43UnjEyi22r2O4UEl46hjJ3/s0mQY5f7D
r4NXfO8mUfiiyoZCAw42DRFFBm3xVSql8n1CLOcul8Co8YMkXWeoLm1gNoiSXVzX6v3Iukho+Bpw
FZretZUWAyojZhz3418WskXe08VzQ8aIywGTmijmJM9tP+GEu9wlRhISigPvfW11Rgy2pM4hoZXp
2MxbCirUJw+NfuEHIc/FKkQahtb4DjibAoJ2xNgCs4Trw9h3bD3MCvxcqOSsW9l5uiA2cT79SOZU
i7yd/zwCXrC8YdS55gncEdvY1WLeJzxpPzTHtIDA//yrlnCAxEqqu/oO7A8grJMzcXmdjziYjnLV
Fkoi0jf5yIsdZ+IYN8Bw18u/Fx7DseNRzUrvPOd6RQphkYnlthGOdHMNRkHMa0MAk/G87dQ7U1j0
HfsgKBbaG2QrRYVtCMa9oXa1S7giiAqaVlH6NVPqriBS17PmgsjGn2dNEDCOjzuZV7lgovqQHNoj
ytuybS7I/b9ssVlda7054DAhz3knqJ8loDf8HuyNQ8FLD0HWI+tAFnSFp8HNj/rcR08AQc2YrkLp
gpbacbbLNP50m8lLvfS4dAmKhfSf+vgzzooJr+G+jvTk5Rv0k7hmRY9/qSMhkrHiwCAbaRFYswxb
xtY7C6r7MdLAVC23xgvXM7a8KjKDz9YDXS1vZaiHZds7/0ahnvqc6t9EKkipElgGdoMYU+hwj+4d
AsJ0PzEe5rzAYHmwX6hdBuj/37Y0QWSCzZsGAZPuVmSiftDX9RGQWKclE7A216ocgUF4OQuEUIRT
7QqajCzj2wnfiR4ueEA/kEKhUWPDjWp6CVGNi0PXwLLTVPjJ5aismd/imuBStLgT/MYpERWRsnXH
4PvmDOcGo58S9270FFGbaPJbxCGtOFG9s89G2+xCZ3HThGlgZZ25NVfwuuuRoaW3kj2bRzMxm/Te
YgwmEYDUtyqRlYPq64ZYb4v4eEScAHtTGd8e9MZxSmxLfxXtzH3JBzjtgH2N+eBfcvqVJOG+qnEN
dLmR4DMeubsnm1qf4LK5DiotUAC7XitYrPOVLrcuBJF1SUW2XKsK6g+gsN/dRLzKm6ShuARB3wl9
S/r1ZdodtNrgiubViCWpHUxezM+dC6eBUUwhEBmnem6hUa8apLuIv2CII+KSjXBXvwBf4c70I1kO
BwppFC3QuOQpK3Kgkq0RA7srGk4aO5EyqpIdw/L5cLdSzZtr1lC0cPb7yxaiTM17NA0DtAa6YInu
BUoooOfADNp33Kxt8vEJ9+uLkI2ewVX8i7JW03Op3p2yLTK090ObUPjiZo3H/eyYm+/5LVwov7BZ
mPp9SsXRorzZkwDBN3CO8DhPLj5l1vKcrjy/HUO2MoPRkg79nGrtGTb1XdAZkbQIfuG1T20Tgsel
RKHno94QpVXz+YWwhopOyqof3pREShnt3sh4G7TaIFaU5nM4U3znXYUFVxCUZyLJvCtfjyNG0lpu
obCXG7O+4ELsNmKefvGu07win98iK9ad3zJgOo+hB6/ZW2mmVAFAygznfVSWnsKhbphsL0diFcdP
PJWzhzn+nv4190EFv9Mfu/du2bXtvrLXSWS0V6QrI8Ln937ksWLtS3Wn90lWh+0i6kY/NTZoxKTx
x0MucPr/XbIlGzmuoAY7CksPkTBYbjqsbVRe2WTLR5AJlxO8g3ouRpJRW48oC4ZQsxd97sbyaFxg
v0JNNgT73jdelEUlfnppBYKpchJsD2t0E1uXf9E9iy+/tV7x/9ojNq8OlXqBbIJBIM1FsMxVKqLc
RpwfGdlIVhPKBH0LJPmnFU+00X0BBcTr5/lLZph9d1FLWTBKYldZ76cQdD3tyk/+gmd4FjF5Z3/o
Yg/fGdgOF0pUYtI8vUL7km05RBJgZpZ9vsb5gDwu7CHLf221iac+d90xmyroVBF0nBJoYszVCnPa
Htpzt/ACEcc5g3QkODHdQlif732oA16WpojFgp2i/20VAVlYLqkZmTfsMmj0pgaBRpH24aOq7dFa
h77amVxk0qiRBfAthGEEjmzkRHBGNf8vU0jNnOtYkbpbbMBeom+asHcGRUTaCLC45BeFbM19oEW5
GcOWf+gS7ECnGoccE5XgidPuKn7t5JJloz4sRIJCOwg3fOlI4Q2Qbl6eEvsjy/EC3PtmmY+YxjFo
Dl2fwKsy+4r8hcHnkoqA5ehtG4fBpTlAU0d/eB4SoFYwJS/N1Ey7EAFF+MIRXemjwEINb7WGMSdr
rWSB5YB2tlOITqrZthIlztjXA1Yfrz/rJmtUt66FkNMNMVd7hkOrWEdKPOfyJWmBH26nEq8/6/VD
o4E1fYhdkrL+h9+r2c8LCWdT2dn4FkO5vsYWN1CAY/v85w27+VQB5eByy1BDoZnsX/wSQbkERr8V
dlukMDaTCZ5kavVA/G/+34eJUIJj5OL8lEAqd55tkdij1dkDtjIQPVzKxzE4kGybeFj/z7+8gHYm
Z3y5haY+lTNKBbyBzY2dDBpvq6TJvmqrnzGMDOJei3TIki3vnMjyrm6KQHvqlIzP/331KWHtiLPR
6t9OyHfgBs+ktONPV9Utv1OXzRLt/W4DAI7VR/wKx7HXpW2Mn8IYoZWdpCwMqM7+fqcHlhluw49u
bSQeWvtHpn0+rlcDW17xgi5tiH9YehrzKKVLnBu+OsRWmU06YSA0kXCwqlqq6+knasR6dbl5X4NR
/+MLGq/2M0s6/LSwBmeCtFEplhyzhDNyKGIIEkPSLdVKwfaej4NvpOO6tmr+S4qKdRfuJdXC5uM/
rpVOZDmDjokZDAD0g/JARLzKhgShT+SH3R8haWqrfIJqfsgvWV2HbWn5Ng6EjcMTCV1kQ3W9CEHK
IOxQZsz4HeJagWM21tqskfiLQ3DVnj8IamD6C4i3LGuFXSiOUo3jEXRkhmBb8dB8fwdbaYK8f/x6
letWC02g9iM3OvIGvcG/Kabkj6fvKFfwYfcMwfwi0lI12W5P//kKPd3MqzeS6wSG6pwEcm+LdBH1
uzeA2Ewn6Pglhu8AyV8NLrbxLig7/Ir8CkFSm7NhEpmmUeq1amnnz4u2fQwZXQIoXZsgHfp/8Rf/
tK8odL6ukad8vKZKrES8dGa17rcQXXwE5OmyjwMCJWGdzOkZZOq2OqNas43SYHC91AACgmSEK8MI
mmzMr87dpwqVXL0UF6HrnPV5RiaBH7ybLRlFjASVUV/LddGK3A7oQjZicDVbzrwwuj7QdYfvwfDC
31Yo2bqWOA6IWz2npQLPnXtZpitk8TgYB6LtB6CvJd7Fnkb2Ot3/HkT0KJ9JpA966ObG/7w2m19l
YuNobsuVybkcOmfY00t6VnPNp4/XcCWY1SsBXrPzId/OnZsH/yYRhQp4nYvQJnbfxqcLj74LHi/O
iMfhEpcySSup/SRmC25b+PU6JvPS2zjcGNECMInJq8ayZSaiSosJ10d3TZ2pSUHiQhGW9rYaqT+U
Ngar4V05EwdHDyYLwhAvZNfQ/fz30YSYZD7+viD+Rvin1vI7HPSI37cGfSg3UCezo3yYQaF7j2GX
nc6E9Gewn2UON8BKSjJkWj9lKETLNRjYCVDdLqfVoQ82D1dVKmsgeCMse9/P6ti/kRTFDaUihAdv
tB35QZ+Avbp6YckPs9lc9ByDOqa4ZKkD+VdskzGK4kQZrgL/jDgGLlI/bRojj3ySzJXu03U5GXo3
rgBliuNWsz/yHemmRJBrxjA910u/QLc+x11V2sIA4B2BGkuLyszRZHE+FHof7C084kHvZMAun/c/
IrfWkb35FK97v2a5DFofAWBCjVyc+T2sVcPC3M720MvQnWEpyO09gj1s4N9i6yFLYQtEdSnh4Fwz
vSL6sQKlG/Sfi/eIbd0mc7OTHAhGc4CaamglWtFRgvQwmQkXD9RY0eNaS+zbk/QvGjNP/j+RdoUA
eyR2QecOKyNBvuj5mEuVm5GCJnH/l+U9ngpPjmg+91EVXv1k8w5CU0pRsmGDlBen+2nsUwToBMSg
w+ISE657aysibts9rRbbHZ+9V7r0pPKFOZr51mcTB1fDCgfxSz3AWcWGZ+I2vT7wA90NyDmHxYVS
yCg4SastNrEb/f8523APUVE82Cx/SAFhqrWPcUKSCZ6FSY9heayEoFOVOohiTLDvEhOmdO6VGnyD
N2JhIwdG6TXy47CUcsIThXVJTW2fIs6F7PRQjXN7MTPQwO387UQwc3qYoc5sLfeDFFXNH9u/q1DX
+4EQSAy5G3zAEG7ybv7F1HGsgiv1ut9QHcQXcQHxQc9nNuDhBpRgq+PdBaNfpRyB55ZCIReao8fj
KW6boJuMxcx/k22d0T4S/TpK/cecAHSYDzuq6aOJlhTU2P0Tpd2QcASxHDsGX8Sf8rYPvvXBabt2
yryVheVmGJgpfIf31gdKBvzSn06EzikdB630TRXkbnpVoxu34J6oPSwQ2Wku8Dr/2AOqRuw/Ht4p
wGN+fs+r5dQTqMJqXYWQqkvDwAGI9hV+xCE7JqvS7duxxUSXI2ITTpL5YKXk73BMp29/DCWUrbo/
gyEFoF5DcBFq6rn9Nn5fVgVXGGCzZ8GkPREyeYGA8A0ln8AZCTv0Lk/RVv/VWAWp1+93sh1AGWIt
/F5di5dYwU4J/YCyf+gbzXux3FWmnDZaQ61K6nUII4dBSDXyL+GBTJ0FvB29rkMr+kj5D0RVSWAV
uAMevT6u+I08lu8dmJ8jrlplOdjaS4p2a3iou2IEXEbtyjDoUGiAjYiLsckTDW99GTPdhp/gl7BR
i0T2O9ixP2gLz6aZPzX8YklTjQ3zDMeY4QqYrL3jNZe6/QIUurrtlXMBkiOAl7324usDOdb6t5u0
BC5yEdYnactEiTYB2kyMwwzkPfaH5Q67nt/nOyV1KoFnwdhLjwkqVjQtmIDpXfzxIqf/jcwHkGJR
OxAXervpkRbcV2p/oVtN4kRbGmkXh5ipWUJaWQI46pAsrfvTtnIlknXS6k5CJurOV0T4NKuuslQB
j2pWIAHcwW96PsMj2wpiguAEnk8i4gIBXZ+krvGlRIDuRfPHMotRcrE431PzQ8C6vkXWdr2T2e+x
S9gl5tupqjYZnILF6j/Ly37vFzoZcyg1ltBUkbOEFF2GHUWatzjx80tfrY0yGX1lafRG+ZMn8tPO
ASkUptluUKSStt2vQZ2gCG4J8/kqzd0wnB5CJ/D46Wjjmz+5ejF63oMhPle171VIsbi0tRgpA0N5
tJVqBk0iC1kaporBpRHgdNKYK9g1xykTSFG1NxgsiHYrWf2OiApTwEQX92FFkZ0u0d+cU+xBjR4h
Y2qoI+8JH5FRTwBfzlJCwgARPnfX+6jZq42q9fiDfEySrNaBkmN35223j9dTvCofLyBT+upUTBoo
7d5Bc6CEpyq7Pw7I02iGtyeHxAwkr4h0Dx387tlEDB3vbTepS8yS8theygZK/14cRf5h4HIV+YYU
e0cuad53aZ4fc9Wqb7eDTF4dUZIOuykPFVetJ8g19wYsTzABE0ckM5tTHhyk0qWCzWlL6gg1zqf8
XsbnnuNBdN1WnjcefHFB8YsIb2B9WxI6KH3ejiAFHynhFvfODK8M2+yeyhefMPcreDzZmez+mWHI
WZUbh2zztXqOTVnxcIk0vF+Sasxep+WRQHiTajpJSbaWI+frA9pRAe2U449yszBMpGuEuKU1/lFo
e2mim5lOsjGfAc+lUnv4AfdEsYSD+l3FW5kGvw/KOlLNFGPEFlXmq7sHbMuD1xa2mUX8fHyWK8i+
m8GEeOyfd7m0ZOQdhOKAvOmBlCEo1LPrxXiVh3JWgtStKZd1iPBc6dumVJguQDR6zAcuyRe4jVAa
SBJl+s598wwz6Ai4EZUDJkS6J5P/3B+uGC5STQdsFXf2lEVoFcG2a7/l7CSVTLwfTrxq0SMtOua7
agQujuu2+IeJWzNInGBJkclnpgLIDm4CpAs81CBsRmD/kGdPrTAAzzvxbBRba5/MFH4o3amyiRwb
oMj/3kS9enDoRoApZQLHlHq6K9LbJ7HNU3eDDYsTmYPfrtU7VhL0vcKoKeATQXAHBcqUGQaRAWa4
aA5zVJEiRGxiMB/kFXy7At10+CC6Momy2GkydYlt6xMN3qm6RFLWC4KFRCmDo/WWehSdJ02urlDR
IUm8l5lxw0L3PpJX0TkBgDC0gRrXyiCntu3I2ujAdQ2XWXprtxpV2kwEw8qmZrdJW4wAWusbV1fd
uQ4m1Zf4bLOABPtNfpKo6q+t6ikKKSOXNC9aYKItHrW4kaiuLQIdFX4J6JTCGrK4NZGp1kUs7hDp
VZgDb5sQMR/u/8Be+v8VqocPpiTZj59ucmouhVm7FoTHweBQAxbrMq0FMamFUl/lVfyy7RF4FhSL
kfczWNrE9ufw0Sy/hCCQVdiIbmkvriDjAHp5MhCGlC1vYMFR7I1pgILKZ8q4kWuW9kRGvQdToLB4
jSL3ErHnVMnwHsBw4g7iUClr3AmXKlURFQONtgEjxOEObXpqmLp/d5HKsbFQcUNm9PNNcVtQn3WZ
09w9FoOs1Lc5X641LYnyYCnOdfmqRTbxuQ8HeLXo8PrPdxXB6nyjOLtqV72OoLyMRewSq4Nf3/ze
O86QJK4zeJiAoArS376jPrqFlj/8KP3gVO7DE3As6U/v1BdwmtdSBw7x5kIFCZ2MGmg1DjwbbD9j
kurhtdd5yspK5rlSWXkpL/dz6qQ8w0PhMpLANLGbvLBD71V8+Ufbj2BK/i+dg8UrQakKdvMqsxy5
l66Me1Y1uXnFdMdV+t2EuQKA15hRxSU1UEOQDnRgaeQojAlYP6Hb6c0pqKaa3DMfv0ksclZdacJb
23IIbDmK5OqyIjuly/Lu8lNQY1LrAV8rirstVOybTAnMHKfyqLslm3HqHuuD6RYuwtErCOGSPZ+c
tiq7cgt5uxH3WJj7YXWy56eI5nNzRgLxFxj2BWFtj+PXQgNswudOm2FxAqEINAyV4O07EglKY69x
5mAeb31EyRVaOctYQ2y3bTQAWqqInvmrlYa1gBzvTulqwCjwxQoPeLx4sCAPrHHGx/I3stSoLcO1
gqKT38wgUjtTI1UckibyVr2UeLz3cohhqTyFu1Japb+U7jQ4L6FeY7eoua5QKowQ9SBCpnKZYNKV
W4SbqSnoe6PuEL9fp7fA1/0Fj+5EoxauEJlcbqr/dFavtSN5xmYTkBtryvBa29PdZlQ7ngBGiT/v
rJIOp3Rz8VgXUB4IdKiRfAm4jXPj0N23eej4VlJ6W6MLisFCjxcoLIaGy9xjDbMosJrmpb8Cw6yD
hPLco2WBA8j4PaaNzzGH9UMEGO45aEf2YCZ6JPBAMA7u6dGR3Ipa84fvqxL2TFfwIMR8hGg0TQ63
vArIvc0mwRLwnvc2cJ3eZkEyDnNcSBtcPh7n+yLKBjKqthCc23BKC6zdTVN29LpKMGywtnDs7kpG
BqydhpyeIXLmjgR7FuDJS0m+3Q8TDheMrw51LiaBH0pP/MqU4jySid3mEtUPMehTApnD6dZzc9ie
/Etu/Icr7KrViJntlAWA6DgU+UmQ95rmbfiNxbz08RCOoXSPUhvkbZfPblZ2o6JisvHlF4+LCinP
/LMEuk3fKqIAVKzxLSgNwhffa+F1ndsCDAm1FWqYTVLWcKyMUYBdrNg4yPFYYlZTg7w56pkJDwoe
oCOdtY/6w9q+2KdHW5WqeGibJ5AfWY5az2x86A/mOJfMXpR7S67pgQXLkoOU+MCSKaz3JJuhJrgf
eCNeE0hq6g5CpyPY+lFj4FPr4gvL2/4DED4PKsQ646gN8yz4d9UargtSyvxJ8RHASbkHJoyQbrIy
Y3+0Wbs2Owruk9LZsp+nV97UXojatE8zOJxmphYN6CSrZUh7uNy/NKpgVvP+xxKlRYjQdao4r7jD
w8VXVrsVRln28wCC3mEDvXZEwnLqQ/3uJk2w6tj4qwCupbYjzluseWnY7NlOgCM4A3tVSo7G34Vg
xC8pgez7L5wWF2lekjVwX6Hz/wGN0tj1HI47nqFAH0VXa7mjemlrZSRL793tX3grqIDNZmFCMS0X
6wSzP23bBpxU3FF8LHD0+1h0C0FxaMCgqJUmctqLNqFQiH1ZPncuLoUJ/Dyrfg/vVTEwPx2sMmfG
iGvZH1ZH/TYj8unNeYC4jZhDCdnpfiJSyNZ/4bFFqCba77Zorn0XL/G2ZSXT19mMjxOF5OGTZHiF
23qVPRWUVqgvtcarpsUoQQmybyFYON7aj6wf7cHWz2GWNIpODXlTYG3maW3K09IbLHZ8A/7vVeu6
VKy5q0U/hhZmJrUQg1t2vKU9IvZg/e/L9aZ6kZPu5zDot8aAwlvHeoLhXtlaobYoyku75Fje5m3t
VLqUYZv4bYYQ0PkWpDb7efNu6OlFz59LFGeT/4TxujNnIZQ3sKQbKkiWdEExrM1YNGn4V5gU1INO
jaGtxp4y6uCJMW6TgtMDLW5qBcy1cHnH1zgLmKbGX2Ui/LGJcrcEohdQrK5uRLGlrdFgmkErVC8X
+0azV5tD3MAzbtxHWBBmcvwRVEHZL1pIB6VvGucu4w0jTXLSW1UMwrjWfYS4vjJUwnU5RpfJ2HeG
didepNVBCYEG7ZzAiagh/h3Kt12WqGMG8rTH9f2DD/xErnwWfAwwe3bWin4FMaWVJogNTkaZ7JaM
MgPBfRAT55FnNX4tKHuXJZ4WHPi6dHk83uM3jJwCv6Xznnzu+SXnt4b3B7yOt3HVsR+wll4BpEWr
H0fXSHNBaTm9WDRPWlvI0CHqfx0qvLnmy4oUnwZv+jbmesd9Ahs2LGRDjK+45GH5OJjKHUYP8dD9
CrqicsSwTe/aEp17aRfr6hRpjjzVGEilThRnaDUsgzbpJ+zafwTnwQwz03ZZd6wUV+D980+7TRwa
ugcYCDBaPS75iMQC41KauqbxdZnt8qmhEe7A6rgZX0zGpVU3cNePMfGNjQwDHbK4u+UzPj1qGi6G
zRObUoAQmriADdLns+V4R9XsoGv1HzH5+kcB6yrTlddYfhahT+sH5Z5NMSCSog2vpUWWTaKaBVv7
uli5fpGMqEnRp72i1xTlEkMEAhLu+CIG8h/Z51MfftZ9F1H0GgGKcUP0VA+2lzew3OUbp30VQ/9E
idXO+DDdr7nyPwy/KNuxzRR7kcDyNRCOt/8+gXmSB54AAwj32NmOGmIStaFq72CqCipocnaJPET5
4mb3/hMHFGXF27zOp9oQzXhX46/iXOKMPlu62mMZ4in8a5ornCZb7djTA8+DysiJzL5a7V1HNV5z
8fv7sEor/pRo6Y0R/79+4P47J59mn+DgDTam9whf8t6Xney3nDMOOyQ9ibU4LbjWFH1kPhjVa+rW
ddDHR7tuuLaX6f6YbDzEbKdp/GjM38KUXoCfUcRscEvBAuSuPxrYoFcw0vNa7A1651IHQjpRSHvQ
ojGW12UgkvyscHn7AEz+BM/yNFAaq/+Ki0u8zkTCujYl5nMQhNK0WCLfR+KOaajUE/nBpFf3Ey8Z
cVKdBxgcD1oCdueaUPCTnNFYymCfZRJBUeohMOBS8dSqQp6p4/ubo99NgA2SjZbQ1Wq7YK9lqIw8
45DFQ6NjkAy3eAU2TDtxnJni2gpt0LzLPxaFBZb9T0o6ZUy2eOowY135ajt/6lXDC9VWtc9tTF7X
qyZ2DKWQAL/hGitRzNx8yBiPYz+DJyX/WUL4HblX1C0yT1Vy0yyOSDVlFYa8D/Pkr6hkbHp0fZv0
fpIA2OzOKUnwyb6IfmBxGO9kARJjY3RxT+ycUSUtZOLQBeQLHsyx35lXyqpxc+MTS1x+3B0gOozF
MyJDiOXJTRq8NfJ9cSMGboC+4XOwxalfoWe1SNNSzQNe0N0YIwV5rr4MDhwePBE0x2Ao64MW8uTN
4P1/jHc7CH31eF2kr2m/RX+X6LEQiU4TEMax6f4g2e1Osf3JkPB+w/TEfj+Yl2gjvaime/HSC360
n5GfJh2xK4JSYxLGhFX1WVNBFmNNzIWaIicvZhtep8eIDmFjwH2/oXEqYIjKYBd1lhHsYK3z61Te
f3KiW6Mv1lN4HG26Nx/5SMcNHwY7TzIVqHShoKu/AtN9Rn2iPW+ho+QlJ6bME5r8DaGxe2xun8TU
+Lz/kdF2lVk5ar3MO8NnQ1v6BwFqQLiOjl4JkyrL/wLN3pjZQ+kPmJGcydly3FxzPJRjZi9Ax6iV
A91F/G0RTap0tUYwN/0vGP6QpswqH4Fmia4UrB+UBnmpHDzMEdc7ObmEAwdhlmK+Z/koLjRXB239
lHdRVEeuG/spPM/oVOu9X3czAndj+djhXrF66u7MZ0dsiScb41NS7nx4nV4GBZVcsnAe19h6L66v
h7A4D/eDRRd5egMJ9sht9bU62VUS+pETp8d44duuwqTyi2qoCQIV0eY6Yv0bvU9qNFt9hWSYADfR
ooT6iYEy/uZZcW35FkGw5ihyjAXlo0j9UivlRJkqAC3YFXV6KX792A9c43ExOP3o83RPVz95MbSK
zWFKjjl9mexxXVtSrsshTvToxIy1bd9r7AFkI936OtCFK1op1rCORfUGleL9Ix7YD0Na3ZLuzpZ+
0L1fSUI/X+8UaF5R8cpZUkJPkrUDIyAm+hMD5mI07yhBuzySFI4onlQLAFCkHPbFUx3pWojIJ2/u
POfeTopf+CnvI2WWnTS/cVDLASRIqVKI6YVytH9hSnBiSSXoedb09VxO/pghOPDirGGNQJXqA3ia
3SI5EsJMuoxw7RaagMeIvWDrwzcr5AGdi2MC7CUOrKkt298BuERdpZAqhIOYgUMaVb9tK1j6fAlx
dLBC5N1JPp9rmqrZ2eKT0XN0Vi39UZ1YCgJFNikOpu/l4J4VhTli5DARM6MndGAXh6WASClbXUBI
MsCPzYgzSsmS+UrAaMV9tNh+Hs5OVO61cBekSZNK/0WaV6yqe9URzxpPKMyrQIKWgbtrm7ascNFb
XdX9xd6PZLW+kYAmvhTNYti2cB+UzMSHIl8rRr0iwceMYpk8E1r2kvF1BZ4PAPS3fffkbrpuXx4+
+utk+M3G0OrNsnTnjowJNjS4Z9yp7FdSmMWiYmOdFjpg1672E5pspAGAQNQa2m0g3WGqOWNb1Rut
44BcsZyCNo3VraordT+MNXum9COlTJxjbBVbAaGy63B6okzHruwO6B2rOvZSWsST0aJNayvZbWQR
nEXZ2T4jlO3i+KwR+MsBse+ikrGBI3fxSVgt6aBEHvxnGxZ2dVPTrz6o6VAwANJMH/GYOkauonsn
9/2HTxp8lkGKxGwKjv5dEO/rNa7C6N4/xXXa6WYi6K7PJOqgDp5vsQatmHaUjOEJmeYSf7GG7fTG
zDc06jn9zxY4Ctczyvd9iafYM9j4Zq9EH1DHarZMdNxWwiNIq9WjE41pnZB2rIjbUFkEVQJp++m8
XoaVYH4tPc2eKD7wO/QzhOSW3jo2Fgl6eFgp5yNoEJSxwguYJ3zZRRtBzWZjvaN51A5rYmnEJlry
q5Kc7UiyiUYu6tRokBrRUoir+fMgRmi0HBBqWJwYAMk5fbTJvpRyoSb/GsrqaHuT7/6i5fZPZ4DK
mUfgCETZXjzCn0aJV7AUO9PwNN97midS19mSLMk+ytPYC4fbGmj3D0+Q72TpMSZmq5U2kHllHYAs
V665VeIVp52NPD+Soss433Pkjt+QvmjCbOWtkdJr16m/pqNTYKCEnMldpxUH2IDy6N8v9+Rl/HiL
SLcglkKUSTy3Y/l7BdOtml+PWaolwI31noZhZRxzw9sT7jDLDF7X35FO6vISFnZB1JCM/ErtR9B7
GV3qLHS30TBtJ8NiEo8E2V3YQbSerjWZjqKajr6jSUSE8A0+dPmlbeyFCtHpx3DLIjMNkviI6+0Y
axbJ+hSkbJ6FHv4FvaVpmcIh4E116fdRRpINwS4bJRNGJ5YxzuXnNteP/TfCkTXDtdRKqCe2Ix9Y
31vGbddT2DE0Stkcudv4/1E2xRbddoSBZrr+80HBVmisj7abTWm3ONxRarxxjSFd0mQHGWPrBpnI
dkQad7F4VCe2yWBrJGt/jtERlWKloloN+SQIkLl35ZTVXbcvV6L0r5hUuKyP7sSeynKNRi/Y5SBu
a1v2ufsB0zivUyoC34W9tZYQYFinNheIaKn3i1yHybMdI5hhkh5O/hxxaXzHC179Lpm7aTtvfYe2
1OZ+U1Nn2b87D7dK61dIQrOouykGIEq3HqvQkNn4+la08rwtEfj7nIdKxxIljelpn6dSzEUnzNcD
0RWk/a71FCPekQLoW6x4VRizgCwkT7aWTLVE7aeU4pqQmSPSQYTapxBbbzkPN+NDXTSgpcCo22YR
9x+2GxVJ0n5WH6o5YpsOnyfSNpTl6j81g3Z3NmRLBpUJoWbz//ymVASupXDQsHznx41yHKe68oIK
n3S58ZfYygjGXf6F3CEbzSHBBvS4Vxoo9BI0N1nFkb+chkiA+I4OdtvIcSraymlHeq6l/DN9sE1w
FGng0ZPq0xuVraNT9T0wIR01jRujKdfWVYi+jtIdPQU8ejtggjuUha5NNWYfiJbPiV9EICy0gT3g
48S+L2RLRhUPCrZdenIQxArcw8BRlZy363rqo158kpz9dlJqaph9sXXG53+B1C0H2C2q4pQumJ1D
eqmiJKVDjK810nlgs5zns6XNT7AIQFchSfI/DxnSpf7AnO3UZ++DE8DU3dodxhI0ur9i87mVaByG
1WRegXWLyAy2BfaX/XCncGSYhituLjuWHHJjJNNVfgyrbpEAkaL1mcm+zqwmAzKeW7k1iXDmy93m
HiOEAFNE8N0POe6/wHirDQ8YlKC/HRrZ5YVt4FRYTpf+b86KQ0gsEbyd9yI0d+OM6oBOdYva7hAN
Jivzh34q4PKgkRYbDJD5uvKRheQqeErzkyYLPu3u6N6oBp5/UYMTX8ThUGUsLVyjamPSC/7Wxs2Q
UfvVgsEOyJ6URuTZ7PHCVBk1llaGV/KzucnzKfbCGMgKV/Xdhp0YGW3ulF82FG84aHCKRV7XuK44
w2HM6mF3z/IE56QsdPEay6o07lkuqLhdtJt16op0uDPQ2Au0ZY80i8r3m/oiAbVPxjDHKDBwvP9k
v8zpK58+GULY0XO2WVh+bkaRHitWUDe4gSN3TLizSc1UkWUx7U8EmcRYD3qknN4+ohMLZ0slPoGP
Rjw7eIi1JteI8P9QZMdHRzZQLYKHkJfgTiR+CzR4zopqYNYAYGnqU1HUvv0PUWtOv2xexA2zoVs5
9S6kXwf7/bn4s/JIOQuLIgmMLYThSwvHeooERKoNtIb1ID1mrrxUT60/M4Dg+E7dYUlyrHG2g7yR
gsyTWVp0Hwdorxp7R+v9IEIqEgYasne1nxmj+BM6FcElg7PkXrCy7a2SwICX1aKky6gNsb9tLF62
dFt/BAEUwbSC1XxLoCFiUNeLk3inGBrvydsuGH4GUpZnQ0DxmNsVcWZXdO+HiF+fCdy+2J8TprMq
5361QvQQtdQSWXBVSDWRnHQbo16nffPVWlZjgR5SOLvWc01XWwa4BkKHdONlVlYcBtx1vY86OZ7G
pmSzNxyfWmcXaG9Xj3UYvMn8PYof/CbGNEmEYHie09HyRW2UBYZXTNcop2lQCLlz9OF9yUTAGgCI
/iigiC1uP9RMv4PnKy61J0ov9TxYZKKw2YafOd8snDabrh3+DAaejdEw9O++xsXw1YQFvOPLmZ1X
z2BdUgA4/i+3R7G5GAxBSCi6AB/Qtc/t4avs5AVKTla5FdTNfJjHx+mezS3+47MCKzXXEW0ZOyIO
WeTXTemSIPamNnAKoremYzaruE8sMxMK29HE2rPy4Ju+nkJEgw+I8DtqqZDu3a7ioktUNhrVueqd
+hxWKFWakCcBDGfgg8kM2iVMgkubq/Ds4zZ1mYHqMKOyKB4uVXUH+FyCK9rnzkjX4wvMdUCBE4Re
55cy2cyeoe6Oo344loLkAw3T4bUlv3tV1wCgrU7lQd+kycfN2ss+TlP7Hv3xi68+KTqv7Wu1u0OK
g+bRwdxyFeBU0VbVFukrZZEtCjxwpAhpG0H3+iZGOdKDxQgzF/wpyN+F01Cjn4hZ6rSzXNurC82d
Bcd5UyjH2HKomstf+SOlBUeIgXwPvxynnt9q7jBxHughtf91L0gijU3l6EVgWGFP2kgXWkRw8jm+
QZ0kSCfb7n+DfKAqnfcsp565MdxSfJV88l4M/ONXI3tOAbw0oYK+GREK70vMBJ9OHCRxMp8drixS
uj440xkXWBfAM59x02eE65bln1pM26uVs8xXJ+sOxFWmvgVfeFNApGS0BGE/LB2ipDyEqX9EFBKk
/RKNv9EcPvxjsWMZemm5/HbIPgjV0mnBJKEH9/HQs6sFiSTRlWxW5f30rk6FLAIzoc9qopLPNzOq
NcjTaSZ03STlyWqXvY6sN3Gaa/jillhoWR5EVN1EW7uO4MV0V+hbItA5gcNq0tQsv50eJHKyyJmj
By7gFPkK1zjUKugCF5d6CX3QzGOMz6uyt6BYQXJOotGBersAlqhzzRPV92umFqGdrdXb2jc28fXO
ejyKw8Kt7viXgd1iePT2cPbUfnQb/gXjPS6/yIfB07ZNtBJsMwPtJv3kd24mEvyNsyOcc945YDQz
aQjjyJ5aUHk+g13t0IF7tvro4Qc45waHBcaUTrnfv8w+sBe26PCa9xCyDHyVj0eCZiZ/u6Hj/02n
t+FaavUJ5Q5Zyqb75tnvlHraZ6J+yK0wMprUncFAEFIjmUlCZ7r+BqUsHA9vEmbXFSRKaRuVgWBK
PPdm1ynA5t8njR821UGcuTJUcZoydE128FPYtr9PnVhs8hBjk2HeOzV4xxZRAELa2gKUKzXShTbi
r+6+LETgwjBGrp0jYHGnrMs+RnmHhhJ9Wp1swUOcA3Z+8PXx9wEJI4QaZtkFBWgJhZbMTw4/RvBP
XJ/YbTDoguagYF3iOfh46vih4ftAt3kkojGYi1eOXjo7atFvLgxQp47boXiBozaSR24pxtvve3/0
DNFX4GkNQTOditFwzoLT4CoUnd3Myy8BHbZRcQ6ZZvI0E6DFJZwQoqipI8cgCHl8rPvoiv7VgeHN
uUi1FiOWAQNh5+crrGD8e2VtBKA5Tt+AIpvUftz+Ai8Y1xxKmWH7Uw7iTq4bI/uJcd0COxwviNyj
NDLtk2eFkfzvINGGS5c5wkxXS9yWtKHQ8KT93DtqEFwjLoQNzPQN5QkeHdixt29F9eNJsIsVDeMO
1SVu8+k38rFjbg+8YJzmHw3Y3wYSiUyvyG4I56i+kiJdVQH92fCL+/wGMDSS1OMS73xAFekN8Z1o
KFu3gxwXEi5qU5yVSLnk1cSsQlnoMqjKgGbHmAKwUP+mTR1k9BJOdeU2fz7wxi83g3geXJKB/HXb
IQY0+NwSss5UJkMNAv4JKKwAPZot0IJOFoocEkoCVr2fb7VmPxfWg5Sk45K0FhdDLpJpwQgNJPhM
El46iteDvgVCb1pIuUn7gfEuYzCkeL2WXnhotXnQBO9tXnAg1WZVf8PcSk8H958wdpqFsB/by7iG
2vD+BfcT1xbZukFsHvtJLlP+vVXYpcUXTBCgKYUgHWKdtBKGpjEm3KYvCb9C+tgCZIid5I2wtokB
gYOk37C7ZkuYeGzcqVKssNOwiBPasHcWiwoZvGtfpWjUBxxNiXGPO1JBCF1OAsqS/UPBUIyg48Qd
uamk2Ci5/S6p+FKwmEsnLWl7RVs5fCz6cPlP6fgrWeFdY99a0JeMikJWg33uoN1JWVRT8RypU8Sm
RcO+D+6KfUDTeOUcT90MnYruG5ADq0Z7oKfPJ4Bvq/mnpOoAPI1JehoLg+uBuR7xDZXegNowpMYN
9REcNOz2nFbPZIYS7vPsKzN7q2Ou6wyorhsAJT+6TnERaUK/eVHsIwno2DC+tsA3U9+8ntwZMUBW
cdhlbHF2PYeQUDK32U3bfXl3579uSjUcPoVo+GaswTBG98AliUvwTkMwlPurYB17ymMCad4+x2KD
sP9aUvG/JaQ94XlJfaQj20u0VlVs3YUkrQeIT9cJfFIkKMqBO6d8b/gIBMOfC3dnaziVQ6OMpuQ4
whfwnjcXdKpDlOkGH8/I36pAin5MsIOzAukiGZbvmoc9jyIs9JKiGExgdHNd8ItydWEh9axxa34j
xt5MWymimb2nITkD9pQX+ueI/MR5mwFAD1evlM801tLQFketMyrwMB4o9xUvIGWqEV1sR438LoVE
qE/R6V8lQbMUSPWauFXEBN3T4paCO7cbzs3m4t6kA3z/s4To41dcfI3aAYNdtwjreo3hIzCOSHI9
KaqLmQNekxNvmVy6kStBBqkc1NvIV0hA8nlOzW+lg6MKY2vXLz0nvtoXFIyyC1BF5yKTbYxkRfqM
wdnsBGSkOqOZv8G8bR5F48tMk0vTqAbAipu8SIct5tu/b956Csl99wYd2V+i8+vY//lVbL5dcIgL
gW25SifT/sA8tXp9V5CBucbYxUYpbf2yf1UnjG5rCxtU1Me2WpkoQ2J+UL7FBZRaTuuQU8jIO1d4
0fv/RZnSwwQ9avYLa7i5YGg3nU7Ogv2tOoYJzO7SMQ2p1kPmvdKAdou9/06C17Q7oy5ucQQvE5MJ
3FUa08Q+8veYgh3UuI7NRZCHnLG1FQ0OAdN2ILO4kV2mj8EJ85W6srKQAMxVhW/LGNOBnDMtqgvV
JomCDVmI8JjOciA9xAfStbVjY1tgpyrN16hbZI2F9KAHM/O4wl6KdbH1YJDD9IFd1++YqfS3mdEe
KZPSriQW7jVFdvzJ/mTEtNDXRK2RunQQcuDHYBlCZDOldZ+qNE5GcBcDf7cqqyXq0w5lYEp9+vY1
BsoEE+8lGpx9wAq5hk757ByiGDfNZzKDo9lgV1qEmTQJLQYOJDgdKfdOeAbpU6DBaB61C+b+sC3s
bxcUcSRyaGj8464/AXv+R/I1Al+Ohz5ATyGjM4E+t8qnc7DiqQ3HIAS/Xk/z6Q60IQyQpJCz10+U
q5QPFTSUlh8dUnPYafb0xI7jKulO/Ps7JBoNhgPMDhsOIYC0M8a/NCt65NZLTGmROYIjsOnn74Do
or2ynC8sgVnSS2A7FRI1eSLUIkVvHhv8PToLEro60SqdK88M9d0w/zMgKVjh+dBwaG8u/4Z8hvLv
5bbKb9ym2ELHsXgICLnunVc0ulp80t+w77OK0b2+f/8ITsDDrAQKHTIwMXpCMRgmDZx3njZ/suDl
8an7UDoW8D85u+Luz1A75u+KxCrWVmzP3c8f4phIn42kFj+bdkJ+1IiFd86FLcH2P7m3Ze90LVHf
jK6u62j7kQw3e3LhoqgpXXWDq99F8YYQ6tVHB31zFbLZ03xA6z2PUrwXyHYMxL2bmx9U0zBoLnzH
gejF5K/ha5o/DBS1mhN6+X/EbwFeOv4OXMJTgK5AdGVJrr3B9MuK2+BAebd8sI9UogkJ5g7HlhmD
Wk+q1plQr39tP5zQczoD+ToIbaX4Ilczyikuazzqam4lOAwKlZoi2OUj4GWkhqYY2ypjBQT6muvP
edXVXipuvPNQ7FDfQ7zn677L/TVmvVjRd68DLVhWzV9LpUfsdEP+EYxwD+P04zaZ5G2esESap7Np
T6o1UwDMwfp2vTHLs4yHdjR63Kh+4ZplLWv/65uxcftkDCXO9XhWpjaGj6WhAzeujEbblkkdPfLt
RGEefw8L+ZMh5b8eqjGuoCVGnlGfXGYKLiSUHUIKUEN4x39T+6iU9EGdyi6UOd2A8gbtV07R4cXX
01BTC+aDQ1QRRCGnWR4pNihqLNyQ9yJ9B3mxLQ6o3ymffqBG4jRFEzkKtmHRWvYFSz7SQD6G263B
KGYydE0MQnXaatvKzBmqyRIm+9L8qyz8kK00mKXtPt2yBj/+60vvt5xQsmuVoQWx9PkLfXhjjY8p
S3kaTwFcv4JssdGr/bxDkzCUra82jEukYemcv2DCuBdHUBdTEDgqXlu0dDpGvsyq3nkTtnG5zngl
4B/Q/e9Z0hDmiBgnT91jahxPkz1bL2nvZf2n76Luuv/n/JPZXEDKc/Q8cas9NufS5uPyvf2W1TFH
NrcCAxciQqIWr0Vft+NKNfrnQZYKnXWv1MliPtD2SfEowC8XnW/LU6aS1ulPsXNI9oO9/cs8J2ZG
OpGkY7G1WpOdmNVRVWiUF+6BT2Yk8TKMHFqWzlCOX6fiiyd5QL+lnMbDBVnDdVeVLMKXrnDJt8Je
EjyzY9iinMVZpomq+Z2CEPW6S94kqZmrcRFYK0mwO9IclNjndSCESy7QGETAhnrdOsRQqsXlAnZg
nbYBdwllT2MWGHjouDQUZPW3JFLzIgbJiPk5Bwp+opLEiYj5LoYtBNinosIatDhZjbjuWk/gqDuT
cLdjQV8gz/mcg7VyoiE0+goBSFqXoHxZkDWGnxV+T9IG4fxg3+EEzQXyYA4Hx+e8CjKG4gaZhtcq
EkTD5vhu9hncnGPVPRK+OXtAJ3mKoRWpC9T5Iz/dsP6M1PbcZ87P75Jau7Nn89R4ikiA2MtA7kCB
SLsd6ounG2BMs+TG0Z4512q/0ctfQT9L3k4oAlRY4osesO8iX7m6NX0fMuZurLWjPP8qdNccoo05
91eAcqWpa2rS3/J0QYP5EBYmA8/DnUp1slC55IVZ1R5YcA8kp+ZErGMXa7FyrmUu4VLJdGYnCIT8
xvgxT/fD3x0756luBrE5PHQ+fbHm0N97ornWcVLcbETgoJCjIjNp3w2JenLNhUZNznX/d1AWo4Wt
+b3nWw2/g83Kv021ypErWgT8q1zvSulLgjePkHuE3EF+mT8TeQ1HB5FL+kU1B0/z/rKllm3ocuHp
rUmaaQV6mjp9T+k7yxxvBAvGELKQ5+GfvZldU9xjtq7NKqNZVoQFFotuIXfNn/sZNBm7DP22aBDB
2zQFriyWZ4FSjMibfMN8hWWKuvZW66cZPC5eEYDP2hJ1NbnuNULGxwPPRQ/IMAYM2ZKUIB6ld4Qk
6gv1Mqg5NUYT1gGLijAp4RL+WruBnQojitpgL4WBDO/QQ1OMxbQc988tAH8GVxD56RrSO2MVdRuU
Thtk/8QbM5qr+OJapPEwZvJG+HtKYWDrPk8+ipymZ0Heyz5W7Ucs6dowpfGEy8GNZlV0S3IUXNR1
h+FiHCgZg87MRnh3mM7bCsTYhCnBci8U5OQ7/4fZlHc9zfRPxW2dwsbrAU9DULf7EU4535GEmQKB
O1AVm7WJciaRFNDlpv1RVus2+ALgUIYyfk8oz5y9yXC1hRMat6bVsxgp7hclMe7UiOpqzqM/pa6R
D2r0r3XIfiSL1BJoNoYL08O9THPxDysi8q4D0re0MqSThnQyCtc4P7bIrqaYNh4zBhHcZ7wJEK1G
bl44kjlaJK7J5MaZrb2YhNO4GGuK0rzqRA8CI56Ux+m8Mei0yOi1r6s9M75rUQgTiuqLQ9ArpopB
519B0RoRYrKEuuz8KLg7zsZ7lnK+wX6X/eOFADc45cTf8GB0fyGjcTHtpH+9HuBR5dCHWdt4Pl5/
v48dn6k/TUPzLxlaUSZ/SZW9NWmmUBPCUomK91blT4e0Q14AXK2Yw23L5VCnQtqbqA0SQwd7Abvk
X8A6tEScQmW2egBa/RJHbhX7QQ2+4+H6PRXKAH4kQIg6bD6io6YMPdLB9PPujkoePGYe2rHqEOFM
72QKZiApQVD/iRSuLCkb9dShXAtbXZv4WwHsmXn/TsbTD9SgWUQGDoa0vrRR+mav9XTEccFlV5tu
qbTIL+wpOGgexlaHwWjsEYQf7dhRmYsnQow1JZaKUNjOrkFVgvBVURNbdqQJqeiuw8uGEBo+mP7S
x218d5BWl09kANqiqB4J9HKFDDaqqMFj72IR1Vzq5NcoMUftZk/ckM/h8Fcf0TJakI64je3Yjfro
rnIQsK8COEmnd7os/AhSj4NlI5Y21t7NixtQoON9MF0H9GfD3feIIRlZgECF7dF5E0efI5Ro71ep
f6UeYaVkAjUGJhqX0rwhWttaxmws+OiEdVMOBosnWPwiTUNOdk6YYMhfhAuaAjwStDMF1mTCjVBN
GJv0o88iA+VE4w1dHeXp3fEQDBoN2SHxZr7x2e9ccZI3KgcDeZIOhWUE504u0p7u5Cdcqq4Ne9rK
LtYf2vsQ6XyyYJqr+W+rgRttMM4R8WdDbNP53j9fIrI58bL2sP7lXER8nv+VCERIpFZKMZciOn1+
/x6XrQ6DW7fbZ7lvRD1J/YuDok9Yy/XNCGlRwUXbQRH/z+DI6KigaR5E0aEwTnJDnGjo5T+2tY7V
Ex2jZQ73zvRdosIMS4K4HQzuyjwDosvlXp1Iux/xW2jqaJiWeVRyIvIi02CNdSNMhHmG1+7SMZs3
w1CYEbAT66qlyEvbxOPYVrQZhnjzQm8B/rH1x1TMhAkv4qlbvNMVb84LP10t/15+Pn7+k7zs1EMk
UaiQ7KJSy+VHvAMjksZe3/HWdi8Y2mfhIbO8BNqxG4GZEpu1P2gdIasMRE65nnEy2V+rTo3wfaUR
2Md7Jgfb22kixIN2EjJxCHSQ67F4VV2ZsxYZDxEzUCeaawM5qrIWvoXR5Q/4+WiwZq2siiehurkf
RPj1HuK2q/WzO+S8D/eRY++r4U87vPY8+AlOYf8J0Mlh3mkACUefRRfWHfzvSH3AACJNuPJPsPOW
IVaiizq7+IbyWMld0Xndip9uXOqs69KYR+iGk4vkeJmOgCsCeGutXBDlh68h4GFHmllQOu2/PO6Y
47bfLRtXk+c4/7+9GJeMx7CTY4rs9iLXeQnZolOLeWgp2IddUkWf+LWAYvbjDGfz2y6H67dtt8as
l0KWv3YX0stytdBXFtsE1Ak0TH0QeN+lLV+vvTRbnLKDrGBkYKZMH9bTZlOtPog92Q77aZ3/kVjc
14gInoHP1iMQAwFcgZ+3cYg1BPCaFS0B+GpLFYIITe0jtSzYfrHCbK+nk+BygllI3klHdASj4Enw
Di5E3eRO7BaZ6kfZF4GrOoqAXLdZGXuLJb5+Xorwu/kLTXovBcTSHcw1m+f/FTkYRjyEgtLv8IRr
nZNTv/k20pcpskgZHA+T+IOAqrmd/3pv8q5IWrainbjBwhbudgHdgoORb0Q+MWCIl4/XhA3xkydj
o6HWIckp8aTX8MCEucG+U/J1NnGlHTRBb0gUs7xcW46hPDTNRszY316mU6I65/dhQW8Jp3pR5xot
+gYxuOPAPJXPp3AIcmKsjnrV3FxNbCtzlxOq9SHxSJxNCNjwJiqfvYZocTslmqs3xnEO6xtbLPE3
gLuLKA6GboWZax6jCYGMW6paVszT+zmP62fbuIo63etEokAI+myfcagOcDdfuksBSSLl7ciYs8N2
vpHYMan7LfzfAYy03bNhX8pH/K7l0SFdAlL0nXlKo+NyBkHNctz7hOFdi96hHcjSvVeKEwNIh8Bo
Z1d1/TEKdZd2ddhsIUCuNX9/bIK+88iHtYP/UFiMDdu/aoeWUhvGoBQjEbT9ggLE4sMldTtw+1fK
jLGf1cO2NMWjEfSdCc764/efHiTzgNLmXcsZX9ky3mdcRbeDFdypTx6rUDqA2vDpRO5gcUnRqwNm
MdtctTbE4muZ6UIMxD7mRXuCCBDTEvIqVW3QVSj9TpbR3LrGrOySjanJFdR6XXOl1POzrjSNG4rq
9RvWNtvHA5hOHq8J0GIMB8/o2U+AFPsMYCyzf6ctrFYhN3taIt3Zk69T73HnnV3m5A9HG2AzG3g0
FJupQoK0Q65kxqGToZhABdC8qhch3f/J/uPcm88MbAGi7nkrM/9p10QvFIgf44R2YGOB+jsb3mdm
NqEcrC1WcW5cZA63lFrbvgswjUMxZhaVNw2t4IYarV+TN0p3dioP5B5gEE+gt7WhLs5NSu2+WzfJ
YPX8cKagNh5m28vAvg2BIL64fMcnGftAa2fif79+muv7Yw2csj9uDHNDSl+5nBiQGAf1b4yTKF4n
Bp6/QU6hU+p2420sgUPSoHSwBEA8WTZs177FI1LELuTuN9/0zVJbgQ9MD+Rt5bi3bu36+ESBPLWh
ee9KrDM+vPaXv2QFh6OewBg2ThHIKt8aC25RLr8mcnVAmLWRizQnUKsvVY0mbl3y8hVCh72ojT7I
/j95EaIko/6KCaw8nkiqXL4j7RNIzXeLnPtEyWIH+UkqFKr+ovq6wH1WN2bxiRxPmL7xvFpeqx97
RlDSiNFf/W9TedXKi3RlYWsT2njkXUd4xsrA80CugxkxLJHSbVkY5odxXjeI0OCH4UnpqGAFPr9o
TEiX1qmMKFpr6GQajHa+aROvzI9yTLJpm5WS7vtqfWYj+61COil7ETXyshDc1wJTN3L3bYr+iqvV
6OhBwQX7xflMfab1c3geneYAIda9HdtVL5PTZI9LkQYxvdqSWL4gl7HJUbLyVE01vtvIBvMDsz+k
r4u6gXcvk1eJpdIFstWPvJ3Ee7hhvw3Ol3Qn/Kbz2bNgH+28KEgMHg2QFGX98KPuc8TaYghwfNnQ
mupImPsCDZQ3F/XMa+VTJXVj1U5iD7nIPK6NlpidDNMofIUPYo3EybBD1XV/1hoOIALP68R7alXU
J6HBw6TWyGSRJc45bCFzbJd5kftvDQkbJaOAieRtKTjOjSN1ofvElUSTxWCO8Uex9g5A6jY8HVsf
Bbc8bgCutuX7Q0ouWiuv6/XrpVZG6JXaPTpbvxVG+EVK3KoWhQJEjik+GA13PkyMHl/QwoCbV47Q
mRssqettGgU94afqY9wKMX3H8BC+rlQlIcsya3PEzwFEDU5HCdT3Q7uVeDTjKAXiw0IUEqI3xwsJ
Sx+SjVOib/zZ53nC9sFa8HSQ+P181nekGJwYXf4Q2RunBJd9qspekQMJzMdUF0EGN4WlD49525gB
j1r1AuyhILCoDD8EwAJ+AeibQfBKqYfFKTeXZK/vqxI3vb/oHtthauuozVE31kQd9X7ZFY1ULsH5
6Yzk6M6nFXOgUMuHALD74srtSScK9Ij03OPHi6X4oYPllLmvm74/QNAB/0hY7p5I71IthLL1bD/S
Q6Z1+NvF238PwH8ATdhOXtkvLVd47A5iPtdJzrEOc5/g5Gw+S/AIFuiWCPYlE/hncoL+C0hDhuip
LqTF4dFF5ZFokjJ+4KwdHBoiYFDrnX/dolfGgAJ4r5sP+rX7M4bKkflvWz2SFMtpLvgJ40zQEA5Q
2Ntfc0AX73I70lSN1YRf9hMP4IQCR+ut2zVfc4IQV6EdxfjG6lrUfyVGNm15p0a1Q8o7Of5qrwcg
11qEJ79gdbMHJ1sza8MzcwUpSCBAEZZ0AGr/6AVwvV8SI9Pq9usENNuHAFs4IZXpM33niP05vIOy
O1ZezYbuJ7T3sTts+LuLlTnlncfL0X1qocVnhGOmfNBVqsyouRZYJM7OLv8Dv+Ie8jzQACUzwSU4
uPf0y7xXuKcwEEFIYOJbp6D4WCRi1niYFK/F5luTh+PtMEUE26bVYw0BnBhHKSI7xhUeiYUHRK3X
9a3PDinU4QAPlPvni5O74npEwtTa+rsSqSmkDIeXS1ggBOarVbjn0sN2qm0fhqq65BOwF1GbpKpG
ve8inVx2X2iy0AUn5dn5KLT0dSR61w5dGGbGfI8z9B6RBtTOocE1u8xaUMv6xeslrKaNBAHATwGn
k3SIC18B0RAdE8xi4KDXzUb4+cOm8Q1CxYUUdBsXnZw2zi8NDFlDEgsyxDk3exOZHTUHse63FhaQ
U0z+dqdNrWyz3Tthp0o+rpOQsEElsRtbLICuy2+/P86UEvXfDc4N3zOq5jLQZwJX2n0cAtZdqGtM
+a9Oafp3fVXizvFE4leE7j9WV8lYoSfNmGuSDowQEJWJhApcSnt85uumlNLD8/og4Tr/4vylhIm4
7pkP9TZXGTV82AMrUlFYJ0upA/lEN2wl4urdskY7JdnMBlicBAiQWM7O5cyySrR1ylgFgJfLz9zg
KfF3+M/uYoLxo8288fl78nWLrbtsHLxVBF3nyAdyRCyT/V0uePyIP08e7G0KDBRYDBuOjO1k295J
OB6kCiMXo30rnpCzfm/uihgmoAnpae9LMooGHWOeO88xYCWdJuPTsOEQcazXSJDNZjv4zLYZrdIy
ZrkEZLXaIjI2MJk8JlH73/7na9pC9Bw0uXRZfiKw0yvzhByQm0JXtrzPFqMywl0jMspwfhh1akWx
6Jiw0n3ciN2elmEMMcZNDlzNESaaehP0nrLIYUlT52WZNz0nmnTU0xMzHdvqJQ+q1dvw33WTy7kS
+xWhfVmLJgLe8ruVZtfR2G67hDveocfVHiZwI/A4Mduki2lvXbYxhSYCtD/CRVP2BrghIOXdwuuA
ijFohRc082C1ghNWeL3aSUHayQ8NvMF6Inx6GL2a1aoDeAdnR+kKSeC3xdCmRGxy0VP7eUjH3eTf
M9dAKLlMdxlhxsU3DrNAImirVOf8jN+6QHULp4pGjXCuVcQ/BygqUEuXy9v8jdB/WHxJYJAVvOji
/ehsDAf91ASDYr5jhtYtcKemVtugWeOrHHMr/kc2ZLIhzw25K1dQUnMXepEdMmp6I3X49PIMatVR
GAllQzGJkK19sXeTLxPGAiXku/4nLUHw7I9aNLJZsdJyqVGlio7XxAjLoQZkI9Lok5Ll5Fq/P7O5
ur7Y+A78kAeT1VnaE20O6znUx/6U7Gw+59cTzeAUwUtrKMCoInzHu3GP3zXlboONbp/bkQ22t+oM
vGBuvZt7aIva2QElD/BPgGUgZ6XhxBNCO6vVeulXTwQzB7J5+H9z9fC9UX7I/aTa0Qnf2LxQK4CB
1qLl+eaej1MGlWTfaJGpud1n/uecjZJ0VRyU+XfTQ3+PKGy0bmO1fRHnhgYUANUzlgf+dtsbRdlA
ZoVPnhI9c0WLqFv33pZ2TDv3XdQuUmAad2KMlrxx32y5LJ1T0yWndtBePeeZSGjK4CWPtOLmI1Of
WiCSiup0jdL1g0xJv9QJzx3FGdP0YmYutX4UJOV81IvP9P/ORFAZnTOFmWOhsZjTFw6ePccHwKLT
uvRQyG8cvCBnVubIIAbg+Ws5FixnmkXs/kyDW5ZdDE7CeEsJOm8KA9SMk4E90zjLuG/qVsXGTwfm
2ns2Dm1y70QbimuOwxbJ0b6MA4d8tec+k9qgwZkmVeuYEut+FvAO4yqXGg8iT8VOx4ruhqJq/dyG
zwGgxGkAskfx8sQXhFyS/QaGGKlBPnQ3+yI7jQE9B/klR9YqESEDpu1lnESLY8DSSd6uvbcp3YQa
CeHS2ZMwQfwMIP8SClmyI5OBfkPZkZvEEE9YGAAvKAHUyyrpyGKXglku5yMYdnT0R1iXQa9tmvpd
V5gFyMcLalEAeG3dFe3q3oWM13Fu/sGM7dAmz6fZX2ae9mVGsLr1NO9+wd1h4SuD6J+XwhtEzVc/
3f336zHtLfqfzSOQe/Jbc4QyXzItbEF1bnalW0EClu8MzLMa40BjrxUJDbSSKRC5kws427AnF6j2
e3QB6MsXIt1fBg4kyihjfaYo5YtdY7ra0OhlhnFyg+vBpyoNntvE8Cw+CL7Ndm1TMGXhyllUYvzb
j72pyTpiCGzrlEAkcJPdiYSLimsBA73B0Ay3e/92wn9Mk3moJszqgXwULmvkejhog5Vkm0uJ2Rea
jEy4SpvWxNaSl5yhfuoNa+56WmRlx+smNSEn9eyEOsAiMYC6VugxqlkU14HZVKk+mP1uRaFrtWty
l4VG2xwSslxQ1hkP/SIlWHEREE6gDhC47ifDohoz7uy4lDKTbVsRVJvOYEWpAAI3vC3MPxbi/Q+g
IKX8UGXfHljV3g01Zx4X48nF7cDPXizhzJmfqtQ8XTZjBd2iYTIU3Axc7Xv8QcyfkE1Koj2ChPEf
nP082Le3NkM85/HU64CYU0MJtUgbOeq5F7BOP+1Q880Oeyfyk9/iK9AMjJo0/I6Gw5kWdIYl38lN
wOn1suoaKqZ6xftP+QrlRRAMPMfkSJBnYWAVbQuOWNuDLMm5YRrJOxDL+QNnyiEvrXO3fIY+kY9r
yjjYGtTxBSwkPO2JllFuL/uEvSmUNs2D/9NTlt8WCOKhf7CXe/03NkVOQgSICOmFdVX/vDCL3x0/
kJl6Tn1iBZm0MxiPNxXcQnXVAcqhRivtYf4BUIKc7HvuypeBF2XIvTa9ua3dXUQTZhDx2yz5i9Cc
wnTpqUnhGG8yq0Rg8XTVnTIWbYDJx1YLTB5MMN4fXwZa8glXHh5EryivTb8OIuWjp7MBXBk8NnGu
46F4eJPMBjsYIoTy9lZIivFA/oUf1HC5FCe7SVrHUzwLn9lgKpAeJtrZe8nNtr0jdmN1rUoWCM46
aublVJ9HHZC18ia3F26Q61VGxxyDMoi3hNIA/WoBRCOU1Yr+n+3nPpFu7M2hOk3Gp47QdF/4AbI5
H+E7Uxf8IFHOvl+kFuXO23TNTTz63LACDny2RAYflwThLA19eCIBTWXr07h2gyNwPWo57WqGgxSK
VjQpqn9TRytzyZ9NMq8JwkX2p3lMybUpG+LV/6nDJn4bRp0z3sGL5mpiMHtuux1dGmPGFKUl5iao
i6Q8dlvdA16ZWZsVX6yOauxxowPZI3HvyfDR5dxE+82xE0gkhQBWzt8DEP+zQMBwSWLCkDK62YRK
/L1Vk89MIRMQRR3Mp8v2ww80mSST3rGqnXCfltXSXfvll5ZgXliN78aSOm6Q4imXwgDofL8AMd3q
DmMu/nKuxQU+sr/bTL+aqoL541r+dc6m987ANNTv6YH8QqpqklZVbUEIr96e6Qgnzq1GKNQWlcnw
pBwVCAM3E9PZsjwYMKq4pnaX/ha7wRI9GCNk6z84Vhp1R3ECuiGiAibK9QM/6TnCJHCFHCr1NCi2
enSDTIkSBq6dkvRLQdMHU0S/79IsDwaWfj/md3OsXlaGEQeauqFDz+kXKJYMpdv0Tn49RrFMLXiT
HHcFqy47Tocgp1B3Qv2fLfcD45LxFGbrmQiCHGz8Zrx0pjpOQfjDOVnDATQ2air0lrTN0Bh744qk
ix5nEXDW2fc0cBSRqT+09k57neIpXAgD+OGnA8Jgy7W1FHKmCWJ67aKolQoulkex0i+eYUgUXE8X
k6FnSWMUdMgWIbJiGrBJOiIvy7P8fUWdt038FRuBncP4nyzUWv3DShqGs8ZLyhsTblygjClMNtKz
AHFtovfc+kbwFw5M7udQKaccz2DXvGx6CldbfPghD4DUbd7BLDBpBuIsFXLXLVNfNlNEdOGCSdHm
VkEJtJO4nAzfN/FaIgqDEOYLv5FNSmEN8GAuj2Lls9Ifei/HvKMvJZcmoccbXG5MJX/1hUAb2ykq
0T6IkIljouVSooA3OJUwMFKT9zUMlr8V/FAIxW6Oc+xk9pOOkTlUvIS2JkM4qhEflL2wadgQ7yS7
L2i1ZmGm6xe6elnbp3fLxJcZpina06Mb2H0LZzxffA73myQDJb7ZF8hAugvnviIJx1/8V0DYEvtr
RQmT+aQ57TCCyc1zANMqoujACcKYEYu8RNlzusO/LpRc0DRTg3HktZKR8+d/XGRSlnRU4bAnzunj
8SXyfGIvFWA5q3WYY9v95Pzgnn0afI/87kEHLvxg65AMK5qC6/raWdMk3CTkpMB94s8+C+PhR4gJ
gf2N0/meY44Sz1bLE6wZPo2AsGsO4edQCOAEmY6yi8xXF2nXG+xeQQ1aSt4zWjDPV1NdelDq8DPh
kNs9tL5DVVAksVc2OKen9scx193QIecAiUDVfcejuAuTBPUPY1vqbktXzucuHJ5JzqZ3VBzmdStR
sUJJ0vjBVXPZ2XX5rxTjts4dadMX7UZqsKfD/FebY6l2M/g4ru+/kjfxH/HJWDVPJfeMnKtZfRaF
TVfjexs/Uf3ODwcH1bZFr5xBkV37dIi8Q4RClfEojycd5R6Zld+GCVHrnLp9wIGC2GymdpIAxcom
PnzEPXUlo4jX56Z3W+Sqo7FfPlXB0bdirNrgZchp3IJhJaS7kZ+K2HXNZ5J/wkz2JYp0VKAoOZ84
AAk0i+feKvwUHcmZIoJVLgWc495Ka528LEvt0dnj6vsGJVYwAx3hdzqif4ANvW9lU3L+KtFiKfgl
xN+a96efdUVsCRAwAsdNEo1p5qTkRV8YSWzzyhc5hJlSstl9CzYFMOIdUZX0FPM/CLwtndcDuw+w
lLSZtdQutUPwRiPt4OVQiu5pBcYU3vYPuG9gO9u2Ohe3wACsfNE2FhxUK0b23kL26ectYPzwi4bN
nIJmV8g4ZnuLmYNFoiehHxvzQVVRDsvpeToqd+h2OguhFC5BuwTvvi8CuwGFOQHHvulMQl1yvM/J
gRttHWUCFEYDt81QuM/jZBc5yxKsB7cVVKqQ+kpNkZlHeDfy84QjqzPe3VA6BA/U/F1hSSB3HObc
aSu36j/n9xbaL4lc1Sg9qPwlk3Rf5JsefVHwY04r09ADla5SCmGkE6AcywdUM2QarUc9gPyZ2rXM
qE7ft2lAAEvF/YGR4ByBGySEB8sdBZ3hpj1Pi+/9/4EHsDWm3wWBkITQAsFWhEX7c31v/qDeocYX
+g1yB2Z5+z8KgsJxZZP0fRnsJS6OOrO/Nc8Tijv5CVS5ZlZBWjjiagmn4nllttrb79xd5LyrtU9i
M0cC+3dGSxrZNbitKDSGzEHet1WMWYUPmvnlzECqFbE525q4soBZoeTlX+HO4I9aGnL+MnhFoULa
xmp9XqHMlJo0TJ7PTJA7J/3HKQSkzkNSTrs0SRhhjt9YAKEhK99Ymu2iGZVuUMLH4F5B3huTjxDV
pWTzL2JegX5wB6UgXUEKV1qp7++Vk5ocH8yoX4h++oD1eF5s4W4xFyRnOKPgHryNW0JSeTcMzFGx
euzmd4+cFKVKazqRs2CN7kxmQ0q6jLLoA98Y9N8SCtFHW0Nt7lOArIBvDOhc6RSKD175DvDVZu59
iNCSWp9v8CuVqRAjmm6OunB1XYRDb3pVaKmAdItu8ssNjORzFaIMnPq/Y1CC8am/JN/Pv4/jBpLu
EVwltGEkBsKlAFYoYyLhEn9oGIhpYrSlse85yUReTyUskxsqo0gcqM1r2efxISjm5GCJimiMmnB8
yA8H6VlcjtMZZuPUGvOXz+hbHAKMy2KhbZxAY4iDD4pfSgCabdvSpsd2NZr8d1lkDZHY5H6rB/p7
1YaaxtBTf+0vW8qwjgX8nM4E0EWhCbblxn79dx9r8mzrfklNtnyJRMq1xJ73F2mbIE5JUEbArz6I
kZuj6BxwOzlwRZ6SVtyORvr+hWv4EoFjyQo1cZ8wbncS063H6APGi6G+ijEijmNVHNPjEdg/OyCm
VOee4s/dVL3Vgao0zw99lVifk/m/4X/VBEE3sMuSV1FU4XP89liaGqiiAsh9v2Phd/fQGzvvTbp3
/myznAHOP6pOWv/eF1AvTK5/gx+PP1Jbs22M+ktABXGlkCxBtHr2JUXaVow5fQKspULX2gCJJwxb
Vc7vmTi90GvVqUFOG72sWto5xjC75BjdBjBCxR0Ui3yCNt9qwQDIpzfyMVD7fiXlpJU5SDS7UpRD
hnq8HiIK5U1Qg/NLf/nV/CXc2iHCCCJehxKYOOGB4CW7mDuoNPRVshH9OyjO1SPYvo3nbVep0wp+
MMFgteWcKNv6u/wEHtXkyXaTH8lTsmfxyyg4UFeRJpQ6e/weLqiDGH+0Bi4UuuOvH0FZs90yF6nt
RMVHo+thj2Kl/p2g/Mm/MttvonkP9IzoKLdtwuQMZ4lbFW3+cvY6NygNx1LHVWqoA9tT/BmHLo7X
LIFgsEjVb2pNymDrTrZc1fz6uLamy/k7dDnCWl9ktJPUNkifj0vU1//eGdeH3EHDft8nuqO7PqWH
G63Fpo+KAGo4eqQgmbAMdSVaQKjhnnjlW7T/HbkmCZYf9XlR3sBZ5AVLoLxo2E5jDHBtq4qoraT8
qL13ppiv4UT+shGEjBFZyxSWvkcziq5LM0qBR3pumF5Yr1msrpcE3LwmeIZY1u5AvytnHwa9pSwx
Tx+bHlQDHW/NeVwhV4BVwA+0bhnscgaEGW9+yt6qaWpSBBjxyXbFY/5dLy/00hvbKfCxEuE0Bi5P
90EFOJZvcBS0g95TV4HZhLAYQxuiJHkis78GSzXCD8/2GTvOtgf8xTJDHjvfgD+W0t/uqGhhusaE
h2VkB2OijHuT6XE2/rHCABtpLY9uRR8JUDrTOOGnaryKckBu8nWqKpqmgHCw2ePNVnhmf8eUAJT6
ootNdPJlK1MFsj/dP/1xwzF8yu9mP8OOhb9IDzGDk2M9FBmEy1lQFeuPZzxn5TMmvVt5pBxbCDmF
5JJ0VhI9FwHaBGBi4yWbT+/iPbSuujXg0A9Z7wMNRJQxJIMVkfswr3rFbbpaI3oTSsMC/5FKteM/
zbE7WyBM5DqV1XCE9ab6adw7S1ofM4Kw1RQhdYx79kISAls1nH+GCuZe/Y+GaCShiHxnHQHM+bNo
1ZnK9jG6dFBsc3sAf5fVM7+cN4aR9+neKs2HWCr8FS/1R3Wh5AZkxuZFab5DVEEemcrOOQZIU/+Q
5Z45agRnNcFj1GPLnk/6qajFZPYOG2bhb+VOT0vmPGbsdri6vAtFxCVZytCJwFkxqz+pZxigmn+N
1gSpY7lFe6mawVf9SW0lOjl8fEWCsQn7SbnTxQIC1Bw1ZR3ZNourOZz65Fuk07LKd/LuU3sKOaYV
riuT8pyemi+N2GdKv6bJ2hACpBNVv4tBRusBzQwMnP3IYEuuzqm4zkJ1t1AO8O5XdCfxS5oE2THU
rpyLBjvDYxL11lGPc3+8MV5UDq3ElIoSsSzQENwCmiqMsy7sGQhO4ImdyFs+GNJvtdGac1Hoxfzq
1ne+aCnbGimbRI2kfS25zshPYZmS616UQM3dDcg8gP6cX+uuRdWG+GuR2i36TAgFJ2N2QVLVnB/7
yd8kmdAcEUub73uWufa/hAphHT2Awg7Hs3ga2PDJKv9dYlB9XgHSJO2L4wpAV649RfD9PoWrbiX6
jpAnmjAv+mZhWdjSyzVsrYdms3E8aWeq/Vj9YpNURMFmQyp7WHynuVhEhClLjxfC0m5H75ioOJcY
+/3f5sUH+Ox/M/dPaoJZ2MmblEfU6PppCLu1vIvT9FMPGGi2tv9LHswXIMLM4rm9is9UwlX6jb38
VDbnqPv7RVUSiHxycPkz9V64MpWV9SYNNJoMVELEV0j7VnUF1Njjr/w9GjCQyjiHOVZfUNom2XQg
7U2te/iNhRe6a0nzOw1HhHZE4VUR73LNqxceS1rKjKLwaLPNv5dz1zEz62DRv1gxAfSfgnelLxBL
s1iJN1sEh7vDOPqnXn4M/wG/wVYqKjDjtgKcPUSSYNEUYOUvO/v+yaYxB8JYMVvHcAhSVNlZzO+A
qxOMufN1ChKWy2o+Uk1DrdCvpPq/71DHv1Dn1KxhUn8gltJIpmVcivagsGdNFboX4hUpKnNXElDI
HRTHEYpJbPLNwuWXmzQmzZdUHHmkGkyFINBlG+FXes8r++9nKxFhlPRquhCCfIavfnT1FYPZ38Iw
9edheFQI739AbiaZtN8CdijrJ2hXw+HsNn9rOM+N2BU8emQwhj+e6gpyh25FHu78LmpgCd7WKzJS
fjG4uK9q6rjS22kbHkBsKC8ZLIot0FeSMB2DKQDx5kJOCKmQuQJkKLHy71ZxSenLtot93H74FUn8
TtLM6mipDKpJQoVNnpybc5HHDNcS8jzxW7uuo9J6+msgCmbwCP86MgLAGLGGvSGW+WZ5AJay5tEk
lU1YaIfuu4mefo1tMR22Pkbtj869+VADB1csxckkd0M3avPKg/Vtib63Fj6opwMhWVPJyP779je0
TyBhH5i4t8NYGAMrba+J0tsyW1W/JmbEpjyE0m7LLJ9gzHOR8WoAtMMjjSu4Rr454rCkiiVFelsA
FKCK8nvc6L+rmxE+RssSoNjr877NbEV2FitoRBmBYk6ga7J/cVPtGsqYscyBiDTG6/0osgVKHA4o
fbeAId3R1rOhwyrsaw76a6zkZBdf879qnnfnWon4KWK85WpItCf0xM1A/Z1JQpFTTkOmSGDi/wGD
QYCoSXkmQFmX8JRNn7zFM+MZu6YaezKC7eTgOeu/KsAzPj+iW3ezBhoBd+Ew7b3WcqL1U5H1MVkr
tfcpwmU2DE6GkN0vdkoP0xqmZucMzO/7yNBZQEg8y2CsTKuy/sTygIHBZMh+V9trTqCxWhslZOhZ
BA6Anznx3Hv4Iwlh+X5GIZp85gMJUqaTcRSn6qJWfuF3cK3sPOwbZ+OIR1OV/dmJg1V2pWZDUHy9
ktqXQi6tVPzgGvgd1aEwGtSepEHiJKqsvwZ1/jfMFKr4zK+N4coGSyqTQADeF9+DUyaw3TRRNGTi
JnRmalugllrF4X8DzY8w0EiQdclKj+6Pppkp8LuCcfVI4IX6PkAkfo77/JU6f+MiCrs9eVcv5D5/
SxgikUoJRVasqQmEmou/n4LIlr6JkRlOwJ/Om8zzpOy0cszLpEIecse9ud/HtW41k6pyKbUPFhDB
vKovlslquThAinSb6lJXz05ZpSDcXaEOF/satjiQDKxH3jg3A1QCLlJpysWzReThQ4QAkQtvIdM/
qOd+PUdDKwE8tY0nDsIKL9MV12+05y/3eOCoxH00d7PggZWMf82Zyuryy6d0yfwB4veNnuaa6ySl
Xt8n/wyIbo5vFyCZI0yf3sUbFIJYZNGaRIH66wy0njF3HEYtWc+KvgdSouQ6tQbmVQrAjYrGaQNF
UGgWlGbnoh8wufEBjlznE14+cNP0PFIuc7bAsjEUMsEu022bAiNJiC7pwLYER/9AAKkOo4t86EzP
6S0cDvk0MIJUuBDVGQyXCyfVeIsFQrtOcyZ+qvwV7gRPSbRq4/s/u+EHVAIpYYPVMFEiyHwbtXuW
+O9Dh58BGSyzGJ1NXIboZMLmg7Oop6N0WbUFBtj2UUIKEQ+pCk60Ygjc729Z1ToYq+jR3Ne1yBux
GOeaupc2qubdQXEHU7Xq8TFLd4KKKBLdSL83WNYSu58IGEtlCCqJ6Jc9KkW28ixY3cpWh6aloiI8
CiRhc4VOfdLWxsRdVopq74Q8bejEwMhvpyCXDznhMmvaz93qYhWVER4cZsHCn9INY1C1FxxcZTpC
8WRZHaKBMw7BlDBSimOYPhRiListvDAOX31XFRV16ctEOfCNXsMPh9vXfTka7OeZ4HB9P0drg5t/
KkNvU+c7YiZEdRvgUHDRXhWstmNHYaUKoUqGAY+XeEkP98UMH8AVa3eJ4SZK+v+J3xr/rCj7Dzbe
tw811ohuBk6EdfARnDvj241MHYvRUzHQqC17arUIWWacUqUj6dcd/vYrAlZA/ZvtNerktRJMHQZb
XM9Cd3KkaOyGAdzXQkLfK1MSYkiB7j8uwMUpEAm9iOiFlE0Zyke+WoEFi/qOq1oefONzWPtY4cTf
0A6ESt+YjFzMLmT5bwGSn9kO+QBuDizAcQTQNevveN0LIseJp5Lqev5WC8JoSGzLjSlgUk+o2c10
nMZmMlgIt5QYytOMmkeCCeNbwBCDjyQu5I2l68eoTKHzSrcXFMhX8LclYvbwX5GCnBIAHPyCQ+EK
HKK4KflSOemo7aRiDmjTzMVuVV7gvbwvgcw9ROGs+IoHI6KFK+3EZ4BQ5JF92D7n27oMVcFXrWB5
sVDIFt1LciPNC0kttIckyc199We/XI7aG80mSCOwUurVNhJkVSbHlcc5kphPyKjHd4PBjfaCfpz+
1xynWsp9++SDnrSJfJWHisOGsL5NtigoZb+swLA5mpofSfgCofkHkOPRzSIU+27PHqcLyioAm3HX
ur7wTbqPFpW5sgyZ0jNut1xBOSBOxDoya31724jmTtYr5yPlgayCtlnAmHZbH531Ore68JyAatgF
GlSxKnBXIGaOLOxuUr1Fz5+wQcxnBhPQvDE9WGoVgzFGo4i5b9CHV9kDHqyZ3AYfO2AkW/S4kUhZ
lmzI3UdEOadssiR5RGTa1QA+oSF/7Fg1nXO+Xw34Wi3zkKqv9/ylERA8IV7dluZqgoXdnSJn0iJF
iWEYwjL4xMJ7hsZ0TCMpNFNbrnpzyzS0pQ6B0+FFj2m2QTKNv7JbgssCD3tpUjyHWzIoJM12deLU
pFrge7sbEX/J/FrBCTSxI94UDrGWtkdkWUa1Q7j/8nUlgUke3UhkSjKv+LXxs63oysr3Fxx50ITZ
73dLdel947T5NA3wEXTUHXTLAZMMhDU8lsQgeYtkbeg7psf3KONRItK0xxbpWsVksdi21Omm9cnu
bjb7SpHYUggrv2DivQrkej3pUQ9hSw7IG6yXKY0k02bmdHgdv805TANcU3OtP4ozTnlVgLcilmph
8sP/dh9+kKzVk2yV/kKjlaMB+w0z2mpYDoKn6PObuc6TwyNdbpl0vq1F+a45I+HlHoruTakaL7AB
FZYIbgfTXY3yGLFDwykHgoc7u+NpNoxIP53sVtsPbSl3chHLi8S0EZ5SmSdyvQMIitehTi1eiaKw
r0jshjjdh5wW0oBwHHoEkUmqdb1RGjMgb96bZ0kKm+oYrRLa7dL9J9Wu0W7HKxDI3ngas/ky67r0
xlgystEqKrYy8HeJaahEyIjvMWvawBmDWsmRI8ayzfRxn31Y1scL0DUjyt92QYb0jVtGVY4k4Whi
eUh830YyLUn/irRogbaOl3Oppd8xI2KpeDtTKOzpxqy+DTwbZXuDObBztoJrkyFajMAhkhZHolw1
A9UAJ/K6Bb6s2OUFmQisWZ6KNuq6p4fDw6KsyjDL8Q5/35dvu1Sf72BVERdPGbr2cf78344rLcE7
iV7ga1d0cNq5yP5j7HxE+SS8wHIRE34UKKSvIujBPnjhzrP+a+AeZUlpMZmsszPrmbM65aY4pPFN
e/KJXMDeXn+wtSprbmkJ16voQVrAtgboMOuBmvTBZiWNIVMcXMAOYcVXt9deqNb7nzKvELnpzcfO
2Kszf0hr3m23Gx+Gc8QAh+r55wR03JK0xMGp+yRszJnUn73zm75PdJNKLtKSDUaASS50VlDZiyeh
3ZWOG77rkCMzVW/R33esjPczkfKbxXCxe1QcoJd096IYR7/MdDYqSFl2ELMLS4Zzax5sYgoT4b6K
Izi4IUpnTAvZi1MjsU58gK48beIVtmjC1y07u+SfPCFtLJlFXas6UKs5kjNEtC1CVVTYKGFWaX90
o/5wt9tQ7NlZd2sYxd/qPOJZCnx0C0pBJnt1rnc1NMHz3DKw46BtHBtkLnMjPFT1TeEDOCj4ZTwY
+fekobRyUfFHS7QDOoYO69lLZtB/wK9vudcfJA4JS40+mCjzWyD/7bDUJp03pZqzih3V0QASwXEQ
eC0EkIY2L+3BudMKyysqjsJMHFaspnsm8ALBDyEXeDw7+TvScPyb4cBSm2SMrPHaGXNPbhyZyJzW
YGNbw1clv/fOYsSuvYdzOjt+xMpVwr4kG6WTgbiN6tVnWOYcvq51sJjwx0N4IeTEudm1j21+d639
B6uadzAH+1ZDGwWwPZE2mJcnmpcnhplyu59HUgTN+mPawdAb9gCPjGBnHPNI97x48fSWR+XW8Kkr
DdtwABOPXoErk+qnvdLEVQ5Fy/2Htda2p+akAG2CCLbuUV5WfcPzCc2nzELuvP9zPDi6Dj/pGG6j
e1HnyJhgD1nBrozVbrEQEdQfJ5GEMXjHPzDv+6Nt2foXUczuk9Z2td6cKgX9I4DxzoBoPyByomKG
PkyNI09JJ6QGJJaryq+yej6TFJxkcyQtUFaSvoZWvbKNyU0uCchDLbKqgvAmTDakMcckbXvyJCxH
OpH+KQ+53Iop+U9hdJFuFRv/p1BTo0Qaiady/hirZLkQF8AwHrcNqek80VPnbZu5jgkx3y4eemnL
buQ8P5HJhur9FdgK6Bq/H6q2xPaJlepPITNLGirOUl6Dv4EOiN0MeozYXOiGDGlotwdXsvU4sbM5
pyRbzbokG6GJ8Pbj6QcHApKKzDvmDHB2qDCTsc8d8Kt/rNgrjoITkgKUOjdx224KmdyNtt+Hzldb
AFIW8hYAuCi5+NXNZLzDHJ5OwyW+48nEUR6dpQEzxCvaIbenyPaGIhUBhtW1KY4/phaZZZZTKp3v
AjIYO93iY8hl7bcXe7ThIfFeTxxqpM7ymNAWX/m8NklM3o3iRTAn9Pz9n2nig2NGzBDjLxd+i4jh
OjGYJO0zDfFp2scHcFDbFJnD7To4pESgBLyAYnU+p+4FcXb0utKEnl7WVfdLLCf+yO58TTY1zhkT
AgoElAP7UMQYH/n9lJqMSzufiR6h0ySgRd8WA6enn5sVqk5IePtAyaTNfuMm8fLW41czRHrYjy1L
oZLr16Wv0Bp2oz4A0gQXqjk8HKVMn4DeIqsLCCXvuU2PmE3e8WPadHWV3aPeU8CRcf87VDKBo6Pw
+D9leigQztQB8QlFioJb6h7HAwZFzpYLpITYyfqFgOQe84myrZ4fqc7DW0YUbmxhs1N1apYR05N1
nh2jdc0g48LJ/gEj3rGT3hceZ7LCuAKHHQ4pl0A68hFVD1QK/6whccdA/yr2JeoWnE90v4cZ4MdO
oLuj0+NbBeij7vvRRd+1YqofU5WCG7KcnU3HG9uE4dMJhMwGW35oBJTF9hcy15IH9X7mFZssvOAL
RBf5r3O8QN7soYl6q0vbWhe89FgUe3sdSTW2273948OWlqDafxs6RC1fYZKQef4Y64+IrbvHPedW
iz5WVHcIRva75vcCkiiUPoSs2vPGoGHCyXzLywWeYYQMkr0M29xtbTZo5V0n2x1UBAwfgZrhJmKA
Eq5gzFSvteWWvXTnLSParvkUCrNjfLio+Yk21XTF4hDHoI9JuZB8jdjzjG9/IzrpqrLGJH62CFRe
cd0u4SCizW7i/6sjhDzhDCBkrwEnhYy9dRIwje+VCBtU02PyZTIc8qa1A5UCgtchV6q06O/Ts9gQ
jt+NVvQ0SaSKV5FttZCqK++e0USh4AJVkZ0iYSzi30eyWbBLKEK2IblQxzK7gpPWhVO9lXnVqn59
KOvYvwOdrKU8ZDe/NenVaMZelXxQy7UVNjOOS3MRG/3ky/B3hjPPgV0rLrM/76XatjGkGiGX8mXE
BG4TUUZXnV7W/scICkqpRAcBHorhue1TXy3iXwQ9MLrCLl3lUFsXgQI6u9xkUrKrUJGhBjifA1Zl
1R5v4GoKSRmiZqZjzmr+Fzh9L1fpd/zbyoNEC5QGAJrWbfDtKS94XAfp+yfz/WrA1OIebQXxFuAn
+xxr46vhcqVtztALfJWppERWDltTfvUM5n32m5Y1ZxOR9zj9sX+3e0GeHdfxP1i1iVZPkGrm/up2
7yZ5UnWm8LauX76cgiO8sYeS6aCtgFkgxsjCdCNeBk7dTgUfWEm7ouQquoEzoe2xPeMLTzrAmabP
LyThR+i4h3j/psKqjboCn20jnZ1xVXUSJnzamPDtH/oHgLloPpARMKdXi0NTOSfuWnpWw035M7Og
o54mKfSA4teF9yBHgFuUEeNvVRILgdlEuydx1UHqCezvXjmtlmxzT9Yrq2MUMfshkE5gxPnwms9S
pePkIpT0nv1+J5gqpLNCVLRLAfxeCMwqvN8rCTW0W2nPsKoIQmrWW10x92gMgQ9LnkRwggPIlFqJ
b8hpZkw3Aithf8zPNpT9AUswWEzq0LXqPgyvUCbvGJjThUy0Q9BftkMaGeWO6hfMd3DKh8vqZAlf
ZihhQqlvbhgLVqDMbwL6E55/IMQeDnJYgozkpnPnpjN7Eso9A1AcT3hu7H1r14PTGPogEOK50hct
ado2NCMnrG7UR+6S3vuysPMRrHvxTAnnzpjBMtFjT6TLKrSTLnfFRn1pBI82ilfiH0YpSWAYiquq
xiDdlcf1HSCkiDGlu0WWqFYj1DydzbXGQkdUlHoAtAcKnIyKWefd1nw7Kxa54e/2qiRMUe79ssoZ
jQva2Cxftf3Gu5OuW/OjzIw9zynSG9SipqAKlsqC//wG/MaxSycCqFLky5oL5FSRfK1v5vNB51Bv
PbtUPbkStMfEhGgcNTS2ohvw0+KgcuHcFw+EyTz9ec67eclQsmrkPFnxj2j03Y20LGvvpoo4m8+W
ieJyPiTcELSFjZ8f2lBtUHBhmeEw4KO4aOJzMaLztskc0GppYsGmRKPFYs+4CcQDaAC/y6Nzvb2R
Rs1/weVJHqSjjZrWgkhqwLD0+0+Af08+1QBVmHVt9/U+9qdVYaynFttdBGoEnCYBwO4xz/QwCbND
DalBU+kKTJhrSWs0iUwPMgW5D8nruJscpZgeCt2Bw/UE1OfWZQkUVqjzyskJFq/QcZqYRMNnOdD8
RZFHMetvBtxH6nLAhLYZiWJE2e5vmORnGE9Rq1kTCeIiPFpr8D/hjKJqwfhG0dUv6bHH/USUjwHA
dUgbSCxQdzDApunP4trGEQ2Q6lwK7KLbyfXhCeat48BY5QiF24SA376uSRFFHftlp3IonA1H3sU1
McuJbQhQEmZbJ2i8aRRa8qmeyA1jfhGwejytmED11yu6x/bccC40oX6xHlgxJwPM63qtotYNTEca
O1F5kARzcgOiCgSwgPSyVxnmbyy/dKJZGovZZSnUNqX1q+d8zPfVTV1OIBA/ibwsS1idqts/yVF9
UVolNe7j9uy0jeo7pDOFtepTpOyJCOZZuC5K5l8GTT5bb8EiWOJqxtpDFNtuiu8ogFVp4dzOm1Cr
Cg4lLpXPtcuAolS/0f2mzEBXfMjPLYWIIjYXA7uAGnkT+BbtJESQ+wyiOTQyo2UGPk8nfzcv48T+
ajK0jo7suq3huoIkZzZVINngk+RIpByAZ1W76wwSgYgVKsqdPHCXvMPMWw6Z/oKWBlhW3tWhGDYB
BUZ6QntEUWyKvpTswnUORg1qSbJw8lrepMB+rSow8lhEX9a5nRevE7mor00X0kRRwjaMlnLRbwnH
i4KvpoZ29aGqGOCerRpOGYDNMi80tyPiXQqkLSHy5Bthnb9I/3m6pcJCt3Jdba6+gfveP+b6wI8E
OdF4TttT/hGEfQzOwuXrLzzFXt2SfGTerfnv1H75jL22otCpmKWAAHMFmV8//tMPxTzB1vvikzqR
lDz3/RUOIOlidDxlZeSP0ecaNXg+KEMu8vj/9GnK3EdStfc496+s/3HuJ83fSacGgxp1WlWQ+6bA
dIQ6beo6za8ehvN6QnkAKHE4rgbfOUJhN/PsrLaVNMg33iSARmxfNTWl4lOP+qMMizdYfXfjfXRd
0wZ/gzu7Pc0sX6/VLy6P49U/oqsEmLbQI7/y9ZmsU3sE0GfiFXNgBwZJ2z3WCytGXk9tphnv3N/o
CtB9iO5BFveMAde+rGE5m86fkj6HlXVZmKiQcrTOLD/s4levRffn12cLAkOhY4WyajDG3LThIaz9
Y8z33eY4NlEfnbWVia6q8rBlQc3uxLftzsrY+HCtt/nfVOZ/l0x2xWasSaGLkZuedYaxdqpoa+IF
YMYdFShjkhl9OqN6DjOyJZcTfHyfvZ4ElXIF/O20Ceavwr7UjqcaruZnTekQvuykoA/PrzOSR2r3
wh0S7aAsLyzLI7FkAQp0BAofcnTFD5Cnmbw25C7sskdws36fgUpbeFKqEo3L1CLQrTHnptuD1kHp
2R9aEXncPAkaLU3FetDmuORmvcffemQRCBLIIEIf7aE4d7WJ0e6PZeozCCh/0nmyL1fkrgduxi/a
/p7Qn9pVTRv+MjGf01M6hehHyV3M98W1xWcRNfVUU8ZWhb0a7b3EVcbvG6fFt/01M0pcHKyln9Q8
n6knolmR9qvlQCjXamVsLPy2X+lo7NgOYj4J6sTxuj222zKtjVTmDvaT77vVHC/MK8HniE+Om5ps
QaTBtuALnX/cTrC4um4pqAnKvHm7ADmAsYJpRn0qBpQq+Yc4wFi0CYBMUH1XX0yWgpcjr9lo2Hvz
abi/rp4WUZCjh87CllNFHgdyVZYDhPZrNpXkBrqS9mJitGou0o4j8hZ4MWM+D5LkdSUzu/s+dXYi
S+GdbFJsXNqRaY/YSMhMY4pqkZRusJjp9PSqmLxhN59xOCaEsi8ZkFy9VXb8dS3VciQQ2TJTPcPV
P7n4qU/06eva8L+jdX/4hOZcmLb/rTMqbfRGZBDfB3ga2LLDNROwrx0oAC+BeRNl/qydUK1zbv3t
tjtCn02h/ZpTIaa/e2mCMiMCOI4tNu205LSgmh7Is0jMrn1sP+OCIkKjfxhzYW8mo8PXAex9klEX
4e09pVoXTXUeQ9yq7oad71YxSrkkMHQve1Z4lWyoieeSelIG9yRJ5/1ycJ9beix7JCR9k1v0RL2M
loAmjfyx8tA4wJ8ieiGTPLagZgK37FTKLxAHlLy9XciMnw5Rmd78/fssR4O7w/WoImAb+BwwYgjT
RTiikwXvv0eXhvpi3XD9HmpcabMzBJ/fQSDL7JnuLAQno3Z+13LoxbX2R/exkNRXJ5B88c4jflLF
4YbjRpfuz3cqKIcC9kFeSk+1bRRZZGPayAQ2imbDKg6ZKZv+cAfNsiCW0JoulCNBUEDKWMcMCvsU
5ZvVIQklao0riGe7FZLkvPoBU5ED7zwVK7IZYEPkVQCDa2hFUWsFSp3PwBREMQMqFkVKDW0w7Rwj
jMStFhsMcQQd8fdjRurlv2nS/RkQ6MMSVP1joYrrPSj352gCJWNzNCkwqMMesQy+r2WqrA0cxuGs
WRUMRYLSyseB2itZutyMsDArArmtN8kH20Stm0VP716xUCN8FzfidG4VqHN58nMHWeb8BH9dnyY4
SIVEA6rxJdvXteH0lc2GefsWT8gGr0P/UuuvciDVjqV0i0gp59cEdzyVTp3IE9ur6E5seMynbIuN
01SEKMgU51CZI7fP8iVc0QRqKUQdGkJGMs4AQ/7wMe1SqwzmsAqnXOchyUUU/YMQws6g5rHmAx6K
p+Q4v1fD8NYNNmd2iDVt+yZtwXOp0jz7wt7P2cC4IN/DQGRAZ8xBISyk4vMfaZSdsFWXqtN/0CBl
BQQr1Jp6eeQPGfQV5cciS3JL3mf8Wt9/TkVm0tVdASveYD7eHhqHX3uMNjQe8uc3MeNaK59788oW
hg1ymz9IbR7XYisTWRQ+LwWG23/CG2BNyW9RsIVKTf2Cg4bLAWcWc+Rl6cAVMdo4NGvHXQ0X6QYA
idkZg5WOjbBZKOlFZeEssZy+ED1j2xNJuHX4cTq7hCLhEX0UlpfMbm/CJqmVWD/Wij6XLK4vYBcC
YuYC3F+JMMwOZPIHFbX1Ni1U3O7OcVYbwHZJPpYFVxPEavAn25ZbR4FuS8iLRy9OhGFGmy8FFhez
pgug5d0W/SMEnz+r96224WopYFipUXh1Wqi/rpHu5SfkprQsW18WdZC7gogGJjmUgG4EOQqUN7Rz
QghfJ1Cugk0F/cpl5HfZRSffCsgV6dW84O2F0grmt8KDljaXXSo4+eL004Ng0e7mQeqAbVVK6XCS
iaVadEfvf+uWaN7uPI4Krf1YjMhhVrfcWXYHPLELmJ14jfTbKy39JOGX07s68xPeq1D3YWHmd1wh
Kj5pPyU5OMVhpycAKHGd4tozscxNnXnxd8ia9lm5jT21tJUjj+3/OIXUg/5OAtOBJ9XluDndN7TF
9ktI1BG98JdXLiR6GAQwDBqvMBS6HBIXBzKqLXNz3mjgDz6KnWfaPCXrKtR1qU4GAzk3/clsXFQJ
S7fiWLE/deWAoSIXCx+E7az3yH1lQVAiJNtlsaQlvXwH9GvSAHmxN0MwMGDz+xTFl4SbBHPuhBig
8LHxsWQJWwDKxzzYa1CFxvm0AsmfyV6U2bfrihOPsuQR0oBs8kQDa7wf3fcYlK6hAgfn6qPGSGli
00koxtsEn24tQARl6C9G3SRT7KipPPHdWrlBRSXMKT8gSix5EWNXcTLtUXVynDcXjnacyJ7cyquT
zDeUW316X6Cc811bkWsrxu3GNVN+7SzR/9SNp5yc4RiNuIMwTY8h4HyThDibck/1hAhwNsTxH4SR
uQlZiXT50pJ9mqIc/jKOHsh8AQ2tV45gkdFX+DuEAGTeyxb7hgqAVmJPSQnOSWhd788XxkVZ3ihn
SreoRwC0jDrc4dRf2irGh31KnNWJotIE4GvB9mS+X+pVVHSydh1mX7WE9STNLV6vlx14iQkDY/PC
c8pEMel4hqTONVp7AUjnSGkGf2Rb8Cm9j8BnIQ7txx5lF0Fcx7NTlZUCGv8TIzi19ELfR+7ksTCB
L2pj+Gz2aLoT8jSjP41OSMm+NnlVHLxjylfoYkX9riKuj5j19+n+p7YJYoFqOVlQinvvqNnaxKxP
QKYMogOzs+qrNg+Hn0i/GMFBKbyMdpS7FjpK36NLUU1Nnohh+ujKBGN3KOliisZreI/d5Gr/v4eV
b72AeQ0r4YMlgjVtIPD8a7ZC7pYOxJQ6eLin7tk+p8hO2iTDpiM7JWuPrflg0/F0jEvKIcuzG3C7
5z0geOHG0NtHRMKgcPOTVsP/89szatqGHLko0sZwgN1LpWEUjsZWmYm6SuRCia60h6H5WNDfQ3V4
xS8vA+hJcHpDA2dfDwYQYOHJU9H6bQQj2kWlbLicEsL2jnSqC4fxPygmLRNR0/oxF/NOpkPvaV4U
RUBz9fckFrKzkvZvsQaMeNwwG1w83xz75h26vA0HQmrLGGqUr6h0p1GYdMkjNF6KwXTsgEICVham
uiHf88Iqd8cZXWVlVrJoQsncWC7qebzm2Bcq9dfb2psizK5IffnShokZeTSwSBLz6SxthCAcLa4A
XoZuK0QxOYRrBMPc3J7r4Po+hdqw3JsS90CXeGNQSfQdv+x3zyrM9nB4gVnBmbOhgr7bT3YTYRyD
2q4jXo206M4Dkn5jCx1Fi9pKuCZgFx6TX2xeDLJN9o1tv46TnDFF3dKoXhckohOGtWuycjr+yugH
4WhDk10+UcMza9Q4g2PVIC8z+Ok3DZ8EcsZ8RgYRI1VJy55JJ74BB24bMVsm2Z1++m5En5H9JDr0
Q+UGQox96XJYmnxyP9Vk5LKQ0In3fDmm+rnPzI3sH8m0abTLoX7kr/yVRu5us/gVl5iQbm3QtdHB
9ZyVpZ0m/MkhOinBI4aAxSwJpvq56pvkwZUw03uB383f1LJ1vJGGMmV5h118Ca0fymSW0Ah8HhUJ
vBZ5rAZIE6YmjkYnIUcHZlnUYj6fxlS/EGaXIKfh85+U0vvnsg0P4ydWJDYs2JxK1t84MYEy45qY
7t2RP0uyzgTIbLiFBFnBDyV0hcPgbwHv65xqeJFq7oAzCjM3HOexrHYfth7wut5Q+aHh2PdFzGI4
uR79vRlCKa6yVNEAZSszMzd4E6+paGu9FoqW6dv8Jf6wy3h1j3plLVAAmr5+8TPaBj8Tsm4Bi1Ba
ZSxkSM3CLYTPop2EDjRGosnET2gTOSpMFTeJQV1FsPmLOP9jVeRtfhcYxWDgMNZHUyk8ICPtfNEL
2k0F0FVWBfDdsXlpymSKB4cCDHnIHF7VyAlytrKlLB9zYB43h5vqMZ9I6bqOr8tgtqgQJpZxvmfZ
gy6zg7MQa+JLPYskE5vNBJvLpUw2RWcKlgb0BReJPfb3I1YGEA3ndy8Dq2jA2Sgz/uV0cIAxxZsP
1FEwebNVdmWsTjaXBHoWlhaovZCY/OKb/tQUgltXKqxZqJI7f+EcJlVHI9BLEbwp+kCmSXhG8jTp
1vre1DanqgEZ4o8YY1dLBye8ixMvh4Nbg6L3H5FNDi3vdft+MxqU2gsHFTrXSDzSOsI08tuVOOMK
lWZv4EPIcOVvSGaWM2YwZc7PLTJqRVcdiawXa5Ye8rVXit0lr04DOjwosRbNrOEUZ2oo1s0dnCM+
ueg8r4jFhPTrBvpiQT957tQxP4yyEaGTCcWld9iuTJWglfeuxYbd7ehi30Ft3+k/RNWPvTpAcVJk
dQwkOAkRei9YqU+otsh6l8fyKKBXnvtgIOoJ4z9xsL0efgL8yyFJbt8jP7HbS5SWqWClEBIoN2gf
qLBM51kn2p6wJtZwvsXBLmvlOeh2ZzoovCOF8w6wX1uko8MJLBI/fg4jX2ML0kJ+f7dpcXXFE0wG
iJz2Cfmeu96tW3jJuWd0klKymugY7J6XjSGP78sIQ6GnEASYEGMcSz+hmcfDsysaptzSCppomYRP
0m4N2nl/ZeHXe1ypHkR6ESYBhaQ4+ve9dhTQEvwFpUNCJzN2r8HFqd2GdZVh1SWnfu4PyMbBmdr0
Zhr1jIC1PiplLIOqdoGAd8j7Q19a4XoLQVDgoEsBfW8wTKISg2HTbYx+WUU9TyjSqeZ8C30WEiRi
Rh5HYYLByE36PUGTAe3vPzUfphC4Gv6PWZGr30hbphznby2gr0OSZyYpfpHASxRj5Kw8r4Q3G+VM
mxt5vrEzE5R5FTQCbjpCzVF7yEGJzs9BkjtPEuxt28NokpwzYTI/7ZB3be+E+YLFKfPhx5fTJJAB
v0DRlSrtll4frI19RZUVYJuJic9xGDWjcd+OKWzG3zseJsjh/yM4d03hq+huRp2S+ewuzhhE0b/B
KmMfcVhgS4/MrM58oPD6jxtTAjWdsoW6GjzvKEfnNCZWXuK7bjC1JPabbOGUjgemGt+Mw8vLPkNr
EvrxAZQBQlwcoWKw6xSHphItRDYkLODRMwVHxlXMTgrJYH6i1w9kRp2xaScQvTQtOTKtBe2E9ILS
LTXyMoaWfoN2EPG8faAXCn3FWjfH7Z6jTID0CLq0jQhEaWkV55FX3dGPweymX1YUj/Vdqq46eOmL
1h+nRejeWqeYuwUj7NVx30poi/RJBCow5ptqKEa8p2tFz0vslPCF0NNTURjS8Feus7L2lP9kmAMX
3UNHa2srU3tOPYjAmL5nSwX2CPn3Keia+9PJ++cByNUJ37/4ap57u4KQKNYNfwcI4q2C+cu6yED6
pK+eWVBNjk22rMGRduasb3s5bWSl9S3gi1H7AzI/wBTnjQl2GDdmIgszQ0KR6+CpOSZynf+U532j
cvXTqbCq52ZMROyYechW0rtEVRwXBTcQ6AplOIg1YJRZDemJT4zjlI7qbLBO7nc3sQbNLbIk8myi
RqwqjdDBJRdqNz0BmJnsybgPza6tI3r4x9T42fzw4SIEoSiAVWzR5fnaWrhDYJY3IzJIYhMgwC3+
CgPimisFt/ozTIQs1zgzALC7IU55NDI6DoVtZeRgJxhx9/7NnYGsbJJfFBmCdqm+s0qM7VBWXKPB
QWIvcbvjltPLKZ+b39RGNjp2RV3ybMVBeRzSZXjmlOcMR8JQCEQuVmMRY0NM8Z3h5g9vb1ze1chL
uhw+9wdPMoUyZR/Yg4Pcl3bZiFlfcoA5DJdWpF7QMqNRIM1n8vS4zu+Ntt4vZZjKjHpFwYtAJ4A8
3fyb8K2dNu5F44O5NyBLafANrXYn9nMAyaGaIENFVavTk8G25u7KPtc0/CUWYV+tsrn9Z2FOx3ze
Oz5J+EbIbLPg9JGkcf2FUpAYkysRTTGq4Qv0b5VxLYiHEtGis2qwzwLr3Q3wCDfUMi+oy2n6qsWe
CYXWTkXNQM5FXSP2iSAICqq0dtSunTplpn/gxv14xpNGFa3wFZ/QgY8Q+86Q9UFp22hdbXgpYAzP
35Yj4KztUDm+Nq65Ye1qS3RU43UEnmV85ztcYQI/kj0H6XNfCPz/nETGv5O88pC1Gu6iRF/L7KG4
VPL/NZEnHGG0+2ncqa3ouiSNVTean1HkU7A1r7qSIzmxbpcUjiUKi+/fSCnY1qlzVO0YRF0iNBKn
Ny4Jilc++R/1ZoW6ZA/cMnOyjibgS1+LgqyUuwGA/Vx8EdJ/xVB9CewyyiHWaWpngRSw/JgRO7Vo
tcaB+LFtJfO11QS0qLNRCyyNt6amgswJL9BWhynCIhaufL82l9TR3EAGuPRWaq3LAxVQpMO25cbd
/j4R7hLMpJlN6ViKJBltW7pEfewvqAtslRnMYHSR3g1emdLOIXg/aGZorUyJ+9sdNfowaq1G6HrW
vR2Tykl0xoQR2B7719TEkWaW9+lJtTVibnvE6i6Zuyu9enLWD9l77Ezd2y849spTYhh1pSLPbCvt
oiWn2cxmK/cQXUMrjgX5sUTMunw/h6nt2i7KzoJeZZbeGuXuu5UGnU5wqN+kOSMtCS11di8TNn/U
LnfzTOEw0LQtBUSVwJZcyxmRWlETRPAJ3zX7C9NfuWxsYALl8ujRGf248ie4Ebl60NAFgTq14Anz
AuFeC1+hnrSkbrUZFl4PFNmnk/ZzYboh91/EOCksOxA91yPCu1tuBPE8hmj1uVNbsgy9EV+H6+Ew
6/FpsO50rJVW8KvDzV28V9UKeNoXigJKrPrvuqKgZvDHEjF1t5IaR6khJmuyFVC6KZ/rqvGnmoxK
V7oHRAdZsbgulWYHHyeTS6SuM270+4flZ3Hi6/1sWA3LodEP8X6ytNrBc1H4moTovnP9pt8n5RFK
uUrXVf6hir7dUQLRGggCg2f9LKpOP/YSwmkbv/ksRCLI09pU9JMXr1WxJi8uEBOR3623VH59dimZ
IVS1tOPm9KpQ+SMcNKdh9eAkDoBU6t9edtN8apFk9Jm9IxOQUcqg8jhy2Klc5ZNC4WKxCsUUBGJ2
htEA/Kw3d0HNEupfhmabQB0ClTYo+oysfGA31c12ilewFG+j/MSyqIseI5dz2gINspTgktBVpe9g
As9Zfd2mFm2B+RMamRBf8bauaCTkuVWLpjnC5FShJB7oLgoST+0v4qfbyR8zOC3yGHg1UKRPVWQu
lXzznCGye58/GTLu4MbRGSeq4BGIC3yL3DiwW6mrrAxRFI9mM/KjWpGZlts5kHFTJlqG5CqI3lr1
3dOVj/KkLvIyvjxVB+OhX6d2chJk6IuBm85NHMsAkPPFmnr5cU2+8LJUJYmtEGu4JtOees/PWcCr
jL+Ajenu1OaPiynC0cJQgs6npwTFB6XW93zyVUBDGJUqzLMvtFpxipqqrrEqg3CFx5od/1JbcHdo
Ia+k2aEc6gfxIhqege1EKzNfu4bjwnXPsc/0R2hPfSZvzlkXJL9GcaexfKEy832qrdYe6dL249tx
F04od+vC9ZRUVQnTqiqYckqQi/+QL3xWWXmLEsGE0PQA3xjTkgOWnBWcI8yV+n+T0ZhG+wS2Mkk/
eyScdhiZPbRuaYzsmRYFIz6idPaTBza7wMN0mBh+JOEuAggexgSmrqjgVByjEIGWCw61yyqsUMK3
1pmag/tjQmT9vl0X1ZqtaFo1Ei/ywcHE9IqJ/vjahTf1Ma1eKyoozJGQA4pycJ2duekHhJp7Iu4c
9DweKXMnJUy9kKA8O1vgF8G7MpWn1NxFT/4LOWGuoEf9biPPJs/gfzzgXk/0JuNd5wjEPUIJT4mu
IlcE1IuhAJOqjKZuY0xcctSyJgJY3znSqRYsokHPhck2Y2joX9KLKr1pX40ji+hhAgFOLYbq60GC
DXsLRe5yEJL/27hEs/DBVstomoXPQimS9E9VvEpSosUVcDv6yRLUWy4PcOkF3Qask8Z4FWiBEDsW
B7+DQE+SdPcYGx+7koTOwVAaRFoeQ1OaPaIs9CJI+5N2KniHRQ9EVkz1vH14P8DRRogjy9ixr7hN
HA0IdoZhRKqBN1JzXFjhJLhMJKn+Nwo0teydzRQMPF2nTWP08FhF0BHqB9DpTmypD2uyMcx1o95x
Q6Xa6tH/w1iMcGEYle1aPAcDM8HE8cmuN82gxSU63rQIRibtRNj9Uf8VkWzg7ijZg8DxKk0wJP2p
Rgoif+OMAzy572nScWE9t4nECAEPdGpi1Q1o6jQ/GxGasa0JVAsgpCyvqNFC+8K3k0Z50CjH/M61
VF8krMtrznC2r0WqRPkckCAc+abQ0C7WagC5wS/NM1JeaA+DNrfCq+wVFv/ZkTlNtY5StD4uNYht
Dt1Qax+cGpHX/7d6IOvGXVlEijF5INeJKC4wu866W9lQShdVnyhrZfruBuVcNPlzPN7gB3YAqa1t
xLPoQqQEjWPIaNwUuwxy/g0TX8VNC0IZdp6VnoEqlGVTSCzg3Q9/w23ibMhgSkbEX+sb149pvivm
MLyw4YPiJnsPHjm4SAZX5OQ3+qpoZR7NgbOCNa1+ls3I1EG742yhV1NScuU/8dBGshivCknmnqYS
+NFQTl4udyuMb66Pbm5VVs0PIyz7Gj6/fFbeSRB+lEr+1ZuKw1Y5V6yeSUEz2hx+fNDn5aJGNfDv
j1OB5Pr9l9wMKKuIM9OVYsHvI9YwCZXxaqRDDbo1k89LxughIHgubpUX44QDmSUx+IVrPbODegMh
AikDl+E0uE1lsCg2YYNT8kT5/NziHLUWrGttdRUDv+SbLRrbpvNitX0CxuTF49k7NNlnLPKCOzgy
KRw01xYKguOO5d29KXyjd/IpgycdZthlLKvvobN7t6NNgBwQITuiGP20SL7wa2DEURIjzkhbARJy
yoGC0kyRCmSPfkq3d3MOqXPdJXRJjVfNFYlWmdBg3qlX/1MecwTYxJMPUFTsYxiMIzLr9L5MibTe
vW7mQy53Kic6YqGWSDpc47fsSspbZ3nQogg+gQ2k/GyGS39LTX3X1W8CgEh9vNJKuKncLy67YYEW
pYjJJcp2mSRVhI7xv9He2ka5RDSO7X9+vZLKd0IMc4m3yTpREHMJopjmL9fv+sSpXOXtNmqw7lai
jVW1tzwXmF9iAtSOi9J8OIyt1l7aRYGALDeltVWZtC02X7vYPjqo5gtqZXlvp9YUN4LcIz8YJuXp
yIcnyIDM9CjD0C43HfBsaaaRNI9XrAcnnrKBxuwT4QxDWEzicDyXqF346XQvF/DmHzPlQorE9F7w
Yu4w/shD7G8oHVKlUjIxfmYtJtD4BL8r40nGyx+kaJmX5E83WBiQA2fVF5QjmA+ZT7YnbB0leqa1
zTp6JAOkUO8u/LnBU6Icu+f49EUC343GUtV16+l7FSSCFxaIq3O/qiWun31G8KgUVd+YXDTXgjyK
IqS+9YYbLPLVBoism1UVkJOO6tTX1QGwsZi1icED5QyNniRg+41vs1V7RIGt4UvDifxkFU5mqkr4
s1MN89K75O+v90h2fvbmJZFd/j+9jtdhZFzn4zsLiWib5AC5kfmM6ijruKMeYfHH2KKfql2BXL3W
eBncBTGLg3c71bjM5V/zvOv/vlFxeCCsE84VGCvLSZ/KBIL+h4JeRierXHrlpO+Ycp6oVLhM3crE
RJ3MayYs+VubImyEY92J8xX41xt1DvVKJSTkwme0bwZjAVhKyrPOqs+b1KFAJLECNqpwdtj1AZW3
ZDzrilt8l8Vi+6wo/kvSUVy7nIutTFRMovEgLfBcEmP0KcUnSBPcnDvi52ihSPJURbCkDWFbl+1O
KHXnWPsLSXMlRhZ8YV6KdudjzXI3I4uiSMxkwkNkrKw7MR/xF1CzRZsB9aseZXrjjt3W6HULy2da
bsU7eDAFG83iJ2BMjykvXeNSukkZvRt1bMoLE06cZa6Yek288pAQGu+lT8s96DYodIJYutioShyo
sHMAEo2tnGHBTYe3KguZycrBcsejlOx85NbqkVhe2RcPkvvKILk6r6cZKNR4OrMQMSklCj3h2DNF
UV1rz7lfuslpqtN3HLEdEq0Tqpn0V9Rawvn3jiKx3AMrJE129XeLiHPqInWGZNW7G/jitl7IMkiO
ziKFXte3842BGf8OFBfl39ROMa76Vo3SIfLBU8l4Qb24t/wTJsrzoqq0dxjTt0jgq7cZ4aSiDPyg
pckHSmBe8Wlck7ZmEEA8fY1/R0Z5eM/7aUfX+dTduY4UC1TC8wWjTkU0clBc/L/yd5XMCbzRR8Fn
WdcZlfTtP6XqQlJdtbP94vxO8x3idhoaSKYiSnWagk5Oq78OALghAXPThICsopOOuJB8ycgCkRp+
uC0hSsynMhzGJYUd1A0DSxIsfsleGvlQIcLsCYOFu4xwTHhphU10j3JCfpG4i3jqJZj/pLkj2izi
6VsAARyAx7okCkvbVK7NslOCqgP5E878q66fWcJrDXvyXJGInG906pfp68TBSjPWD/R3cZcA8mnu
fO32EyC2Eu2BahC5FVZ0dvCQOhFWpb8Zg4wY/OHHhGbSk0tuK4WVxjd9KtY0Ln+ZMJbudFGDCb8Q
xXJeVwYnXv3q78flHEs1kmmFIEZNCQCRpJIM+e7mKD+DzX21xceQR4iaUU0ROQqEatSOS85t8Nbo
GTlKB60X8QYoGxeARUx1tKlMo9WSaj7PkufvxCuhTDIGIJDJlMqFKxhHVGSu0Gu1bqYRgTMOgjZO
So7wycTyQZhrxSY8+gIgyJZHLvHgbw7hreIO6DrGhFaeQChOp8iwYRpTvlnTqhYbnV7DqKmmV9DR
WJOkJO+BbiGO+uIz9RaJGUDSPTxOYQLu08XOGD+6u9GCW/2zJJ/+CVJzGpTFGIcQekvMyPHInMXO
+12MaA7mN4asIrEsph+zvkQ63EAOdrsakNkQ2+kEGjz/yNlUQPLgbYdGo0P/ttbPCY4S8cEMGSjc
0BpREcAIb30BWTJX6xrDxstZtAPQPvqvbuQGaNzfog/HvKiqfLDyHjXozoo6WSMYn+4um3WjcRAy
fmzavCSDhpzxofEcdRiH0QM1y6/IhnSdHEVl7ymBaWTZO0Ehv0x+nDEGJd+G/henzWzCX+yKfm2m
cuUA3p04tFO8zDsldj7GfB/8j491T2JBGCSvowGrU73qYSQ8aRNv1U4rxRPBUP7R/tfv99TTtsJn
lRQ18dd5Z0byjiLTijSjIy5WkGyB+pAGVraq56JIrxPjAlPaJNkIC5p1xctNGano7NLuzuygqdXo
fwdpon+ENXbQJmyatTK4CnYWmDbpMWUp0X8xkFb+ZrVo2aRY+5im4Omthc2xcv+ogn8vLsMvelNz
2GAEbkAR0MD0jSlK40T7GmxlJSuXBqaYvxMn4wVr6vZS2KOeKYWGuklD1HWFhXCg2uPkiPjNwJ4d
P7gWUTeyoM6Ynj0oeoHlkc5b8QeFYy3CMcw+oRhiRcs72gdtTz3SLbB+omJxI0ylBBSACKrNDBEY
1DJibDVMoM1QhcWumrPo/VAobIyirgqU4rEDnRHQUiVkJe6Gh+Hd2HyHf0rfPu5EdkqLnIvhTAXw
X+XLdvmynTPkOC49FbfjCH/50LaxacoQBOq1mvXpuGcE6jJYaPy77TK2yTYKLEhAuT4FkPmdoKE3
GcYpXGHTxj+GcUSA8/nxO4QObw9NfDiihc8gtMk7yuKp76T8yD9JRI2YtEgluvqgCwTxOZlutsvg
AEMKcNyhN4zhKagbMDVXJz8lX+tFgO9bFxX+iDUvFJqXoCoU+3k9tnMGqCocOqe4gpx0o5/2KF5O
43JFsJ+EH/5mFejXFrNMKQun0RGVdeTaHRVMHxypCJz4+1/adm0Xz3a6MpFbmAo7o25XtFEWQjop
J6ebaDYTBp4WnHGtVQR+6HbZ+7EmTf+67uWWhlXsQCDk2KUhcBLAcwxUCVeLhcHgS+ezPweCOl56
mjeu0Am/CIGOIAKo7YjQB729PfBNxFl7+2Bu+KVW0Xzp+gqt+c624L3fNi+GZ+2Hlqmi5ZsVkplB
NyhyKjXyfeoyZZ9cnI9osPYJIVXG1BILqvC2w0PHK6SJrfLNjOgbyd+WKfwluD8E5nGScrkKB+l/
hlvc1EcrAGMWvwoWjeMF+/bbbhBR2jhgtfPn2ApFyE1Pgd3GtewUBXOGQUE5SSwYz1i47XCF6E6V
lW/KG98i+b4hAOIlHcy60/tay4DZk39Np78xq1URo/XkhgVwtx/+BqV3zDJ8PJ3Dkd5LE3uTE8It
+Ie82K209lzJJ0PsRRROEyqwVz2gIFDn/R3VLfGPYKGvMg5xFZnny0cOWnsj9GmcnqKSpFnkDG5Q
WvTXtH/fpfNWEMhCze2fePk7wJ8oBSskUZ1+tpE9faSEu60wraT43y70d41altpnfT5A14E841v8
aaKAf3nDuiRuzDorU9P7hyD7Wj2AYC1f7+kAWM89ZbsVBIKpWeDT3kbrBCPzKCkYHahW7DlA1a2R
/YWdDMbRJ4OKwmy24XyH128wb53wwSeAUdUw0xyknMmWGp8CwC9jJjbvcHew1TLGd1RJtA4zqLpF
Y3d259JhTHvMQVM9iFKKAEpVgBh252L0zni9PHqtHb9IkGpoVxa0IZVLHehlRFAZx5MPiCLpb3OX
M8OyAmXzOTHkdnhuph/iLfI+QfK5le6RpQep1BRM8gcBOweatSQtr/brFjkWEgGFmfeWvSD3DflK
plYUnQ0xqCzL+WlLPxH3Dzg8VZgF5jXd7Q3/78K9NemoZAY2D8tmyYt337/T0TM/B0mVVm31BsaH
8ASvgvbLXGSMzEP4nv6O3t5XUU3C5eK0ETmAlcjbl1Kgp4re0NOWNlL6v/lZ8kGk8NXgoS7sLtin
n0r0bnWlESsfMNVwHqQwKYK/jtW4QBF0TNxJSBZZqZvlEnxu8EApVYuZYlcJjaz5WmUBtv1DnQrT
a4h+2DLSuhuH+p1QLr5jweL7gKeWZV0hZaKL1YfAs10NcWLWshWJmFV8kRKEUSLteP/cDExCnYdW
EjENmp9ZwMZauf2/tfdX5YUMZZxSRWBcv9l6xC7GMsKvA/NXHjrQ2iWxe0KcJ8MEM7I4U2KCvk4W
S6DYYajrBZzj98X21SBZUYEXR0GkZq61xUMWVF+QEg+1ZvcwiFDeRzIU1w7Si7WE7C2IKjsI+55s
gVbhcq+TwxKWAn85S+JOmq4iK4R6c8sl4v0phqSIhoM9w3/qatGyFgB0L41FrFgBXTQKeRN2Pea8
Y0jdRpIa/A3WhKBGP0SqVSk119nB96ay/tV45xWZvMB6C/uyEfqdXeA6q3OjrGAegmkEgXFzHH4D
1x309wCUNZC8iYdi/XIgZpCq9Cb3ypTeIatEDvLHt70hulku+MoXV5RaVZEqcMWhBwScVTb7Yunr
zA0ewjQb1rQIvJvK7dmT3zKylIRLr2NuP2fG8YHD/YlcoQTGbVnM6nibERhKUc+B4PHwkCZ/lS1Q
e1Pge+wEJmOAyCi3YK/YIPiZYNj3ZeHhm9XzwOD3vvVzyurhX6eXJNrBKLx44ZBF2TTDBfSHYXqb
mQ6TpTBOOpp3CkV5uBEE35aez/LMY/qh3TqG0Y7uTOb3Dq9Lt73uWyAlj0JbY34/65/Lqjy4RAR+
QzgAIiMAg3ynjknzItY0mc/mdPpq3mHS/cV10QxLJh7F/tbXl2qLbnbjuNfVJXzr8ZTQjK5mDrAo
uXmmwxSw1gnhomyQV7MeAAHEbED0iQ0xmsC+6omnXN6xCgV+eqSB1LYp3miL+vx+MYLKqU0k3MEE
Snv8RHejTAmNtNBAvZBdQyyDbCCaAwg9UaP1bTDjFksq6tkIcvDmTfc12MEmuvE7uz7UnoA9+8qW
8PIsF0mmyqH2jOh7yuOE5lmukYRTf7Im6NUq017vDQvuctadZ5sHKfB1d+eTGriueqr4rgYNIB9c
Ru3zL2FGA5Tttz+4vk3WtRCxOFIK5lyhgHtSeEMZHnURh6eIR0a5pkE3FNdakEiLUXF9/m5xK1P2
jx3FlAv3/Di2QZ+mCBEuCBYDn/6YSEUt5wlK4qnGXO5cBRf7XftMWin9+bwdUsa2mmCMQDJTZ/v3
N3Q51UMvMXLz5DLGJMpJQEnTrIsz+jwuSL+4fVtpsQ92wNUkI7OdGH/aAhNxI8om9pMa1z48v4aF
m3WF16KkuHgTKJkGfDqbDN5vhKOmNcdGiFg9yCG/E4nJhSchlz6uQN+NhMQdqVvynEsI5e5I0M7H
cuqZuWBqhbfGmTeQBuX8d0PmVWy7pf8CyDZAVJGXHHKhk+jFFeS373V6sik9s7uQEJ/e1z+SaP7s
yC6AWUREsLrbJ4qt4NQaealHABJO0y+6pgpZCdk4Exh1neYrZkzva6hGf3Fqm9HhC9qV1Nl7IG+9
Be7FC07RqTRLAWnBLUC/zLvGk9qlLZJHXhHOBGjjloUyAGPXBEgX/jhIMaMXXIABNzg671aTw55C
S9jqRf+xflIiFwwHdpD3gi+qW727N8InRHe268uwVCvkWync0bCY72NkR2DUJLXOaSV9Czk5RMcc
A/MixLzdLCkWRlaY2nfVlKP1RA3DVFE6mYww1olcLv9jNirBb9kdwPQbYj/BzQ4bWI9IhvJq4jra
sjZxod5ebtvIITDVNYskpG0osX+u17mX2T1+mNCwQsZR3jsMGNnJdfOzw7DAMIvQa1jwFxzWejTq
/hFnx4B5bRaQt199H2ld7qZOyebk6zneylwDN7qHMd6lb0FptBrEyd7tNnOuhfWwBSmg6AoTQDN2
9EhYa7OkhdB0Tlfl/aKJqcK28YRUeg7bJyIMHXml0F4oE4u3CKTjeWL9bJW5Om7SoUjh6ZzogE+k
nsOkElr7qm0L7RZm69iSNvkjp1+exH94X3Gc7tNJcez6z2e34QDKt71I11yYgO8RiC8JhbUqyU09
rwMXvmN98s0M3sratHC9GuSF1erDOme9GBBS8dTf9yPR5x0P17cqJfwlTOfjA9RmogyVXZM572S3
5P4i4b/cW7PevwtEgxgNG0SYLJwsN//cEPdG5FXEf82WOlVkCsJUI3GJIqyX3op/yv7CuxjthZfH
n5Itvs/ygSrCc8YAooVE/kI18nv0uKueJZQVFnC1VD+dKqasvMaQZTjDhGkwjfVG3ar2cbAFdixJ
fVODotAPeydok/Z4bC8aRxLIFuV3HPSfg6S3RgP2s6HIOhWDbySf/8V6HVoO/L+twUz1WpjR6g/N
7JFjxGPiLGgimsIplqBmrg8q3Q+4g3VhvOGSdrZVVZK4FAkCpztDfQnbhyjXBzgDkQ1QbYWvpSw1
vOF96aBqkkCwY5iOSIfqR78DXLKOEVzQY3p7vg5p/AJBjnSfO4v0x3Nf5EIi2F+ZF+cEF98qnM80
AmV+BkdpkzTwzOvoALQQYPdt+j44ctrW509NoFCnpbtH09XyUV8WK5S2+3A6j3yOR4yqxGdD5dR8
lht6KPenXlGR//PAeR/pjzAwRI6lXNpguOuq0VF0WkDP8ugzI+JBQsItOKih9ZymKXOuD00+vJD3
N4ZH2KN80YSAeP/uWf/qxXXPFYyA3UISb0jY5qlBpCsg2rB2E8awLTSntPleHScBp+ZgVl9uT5Mf
z33p2gYBjJ0Xqwyxc2fiK8hw7X+5Bmw7QagYrHCbj20I4+zAZVFYg7zG0jzxWJFtMwlxn+71aCZk
m2k1e+6+faWu1kwuXInBzNTm09mCzuxZo5/NesikKjq994l3tE6T451At1T7n+LaYLKk04h9Ssp6
99RduUH55QrJkuTlsbnzMIBFAvOrKNgHNSx6Gq9V9Jyc02kKDx3xU+rjQwDca4161cHl24gUm6IO
vE0iSSq23zFuUhQu5X+JOB/us2IPDvjtkUyyyiYSDNSGMr4AwzXSOE/elXbfaSaC2qQvu9wJaLc+
RNkcIQaC6fI2lEYZg3zl/X0ac7mgz78H9r6eCU9VtF05zmzVYGijUTuDSB8bwSed1ThPsa8XSKOZ
rTUgG0XUzz8ELAKxn/uLpp+MLFvurib3gnGJVml8nFo+QWd9pYGHECYH7D/gSptWT1wFdHKN68Ma
ekKaKJVdLHE9nx8J1MkmUXw2K4U9/o/KlJ+jqXIkNhMT+5p54POMEV6OEzx8JzTJg6s/4nGTBXP5
cvKXBWqgkfQj+PkPkJaj/8aQVkxkOkSZ/93iU66iDEvSft2trmaNOFwA4n4ee/5iNztB0lSghYYM
FpNpk7okrkbPnOweYXS5qniDRxpIXAKHuDkmdO+obi4/hFEgVKPDXMl8JW04nKMQrurKvnTrnBYk
jy0iFb51bVmhQ3UQiCveTGkdWKiV90NMMWxtL1uai1Q4CdDtQS72Lc853j/iLWLjnJ20fOB+ggti
Tz0euqU29NDDswNON5cooj9fuwndgE9vBRbMuBTTbLjUi4xGH1DZOWkJryHvOli2hGjuSPrV+t8n
j1rm40KGF9e4g42eoX6oGRe66qf6JhNeALYBzqunaEMVATdBamRgplXDDF8zDr0D5CKkfAPLlGmM
+q1Enel1jdLka37cJQh5LwWqJ0ve4zZNio+k2WXwNPJM3jbacdOg689h9iU15jnDrW048tJq7SLd
/FXIviHb1xw1vczmkB8Um91ZhX0T+RSGgPta7TRfdUeHDPW7t5RP/E04HD9p/EqtPeSZq/ydB8Bv
K0flJBLyaSWJ4uWpBgWshI6m30J/bbdJl4ReF7d2OWhy2CLAXsG/XYDKidZEegHoPQRgevR99dn8
EuOq6TSMFsvFi62ugtaXdrfw84jka7nBsxhyZ0xHLOyoV5MLPp/VKyPdfkqTkPYskw4y36n5Za7D
zIMcNfccEIBsP29czn431mwNoaj0Ov7niibsuL1TAJ0/+TdGA/HY7ll5eLhhpk8VWNM0URf0v2nP
dIRZWgZbsywIwIqd1qpUwQQzJQTxY9Jm1HoM6rAoQF71n1H1nQDDKyHyw/PrSyIsMORvhTIsjxyX
9KDE888rf/oHn1lB3/R1rOdS2C1H3kcQM+a2CXCrMf02bA0atDeyU1Hb9sUpRju4Pq8GZQrYb6hi
aSLDMbZRELuneIC7q9/xnR1MUce26uIS05pmSB3R4JVGaQgN7NCvj7bc9bk0kW46RSd8fCygGk03
lukWAhmjFbkT/+GQXnEbXBeSo8jAQQVoU5psRyeJMiDxnG58032q5pMifjjrHdODJCrcZSYxg25S
3talx6lKfcM9fEajs4x8hcTVqX+8Px6/LXOBckjBRkxpmdYdbZzztBujdTUxm9ci5sX4CChNzh5F
MY9uis3hj8rb6kSzhJRb4MTdG9qqj28ZRqzNncWOLi47mZXJljpJefe9KXgROPtQ/1rlW50dxWSm
OMndK/Y/Ep+cgM69/gxg9dsuquGKKyp8cwaQ+NGzir31xuk9AohATMfKGE5pkbdjPfYp4hwFjUpW
1vxD/Ikk6GCkihE0GCOUsIyTBCTyWUcxCdcJbT0Kgtw8fJ/WYrACFtNZZFzU2sDy5LeiEG9OOhtP
YdGLe2TRPld0fbgPORk2SQcCMcK/aABloPmDKeZ8yz+w4b0wGfqURTfe+Git78I8UTeDVR7NIYmo
oqdmsWmkI3+F6MohGsDLBEpnjpmKLrSSoxzFWCxmGtQOHiJWrGube2TL4D3/DJMa/hf91zSYd0rx
MAw2x0ocHeIF1jtMyYAHlBnkb5kcvudqHKsaWwj3sq0EPwGO23wZ8gayCdAms/BUmea1KzE3N5/A
UJJBymVzu85gMm1AW5USYbYbTwUJ13CacUUrCbaypWzThsB00y7g9wYbZm1AZV9NM9IfA/NSBiLU
7OCo09h4o6KWyBbZjXhyEEXNHnaSXXTYtQHUi84J8y+fc0UTxTMtcZYRN+4XZhQmurliZxZLz4AQ
HxfQtKMBBpe2j3EZe8YsLBxRu0dxigkkRrdskL4WsSXjwDe4oAllo8SlqvhawdyZp5PNoXjdKl57
WnVzVtJc//PVLKoG3m3zc7Bz4r/Cvs8DaW2dc9etalSf2qxd7S+ZBnvEimKlub3F4CxRFohVWhk8
+NMg5RSjDxcHMrJYdgCgxjN74tugZ30X16qsm0CAngwxoOxjwuLB3qBQ/aDy51cdhnISf4eqoQey
GiXx8hIHIjiJ2Jz7KX+jaCx7xNV++eW+e8jMOs30IDP4TIqdGt3H4Uwg4FQUMO5Lr3j7Nj2ncO/i
/F92szm1TJNf8H5mOUg8AaTOnWCWE2YHAB6LRA/KebYbEg+6Na+Nfs4s58bU+pirOeZJI9FrGoYX
kkK5sc8Exmh9Qwb5K6WAGsvIlBKCFVBFFyjZ6QtdRq7Nis83mHEwO5pQtLr9RfBC4NsUcqQDni/Y
6JIXl9IXh8149MYZGUZgYgkvQViJz891H7sEUliaryBNsy6wnT7sTMXX3o7jj65iHNDg+Y0l1kwp
YKf+e6D5GDHmZlrKyre1etVloVmjdiXvKzhlykI3fVfQ1aE2gHj/ZgES/CLE3EMMKwwBsCG+6F1H
nwoz2/4Ugfp6RS4659GhETpCGnS+YbRfxyQRFQ7pRuLk2PrwJjHDAMJlDRRS6Us3q9POdWAZ9Lwe
2qtL//736Eq+Rv6B7ViL7QZaVrz7OWk23RMWlb0MbgTIuHk4VBWGBWn6Yi432qCkPnebWI4wRIqr
r2ZHBcsdD9g3RAmHqwEJRm+/S8uEAwycQUD3xt5ZybkhhLkL92L/NwAmSb/XrMHA4dBDF4SI37Gf
qpKBJxCyxxYmDXYv7bFgb3hGoD6kAqCxHDU6KJWOORBP+nmfnjHYDFoPF63v68JqoCONZmy6R8br
GNquLZXX34TKE0o9X2WzQgHyIKktgsZzZDEdhlbeVskb0a7TUCNd/z/qvyWW08E6EGg16r153The
Vy6pp87FS1psPxT3ofvmF6iUHdLpY5l4YRMKL30AcDdGTtYtZdV68Jhsz6CObqqohfXJs93ytNSm
mggsJmAXuUTfTw0E/d+qQeTWT0uuDMQKwpwuRcncxnE8QcNmlOBCowNGz3sEqWxAua0NRQaY5PKW
lrzjuv4B++dNEF6R2GOaYQz4433NHsKXYzMqxtCsWXloh2vKsBsXAYz4q6zN9I45AQFaZX+zbijs
/Onm8nsICLrIsrcM3/axbOl5UUeWWOXSNihxp+8JaKxnhxjVh9vxWRhmw+3fbAJ/ytxGbqMMZTwM
felHVUq54Ad1xtuM1bqL9KAQXbua1Ku5Xou+O/kwzoadj0nLlni0bQ39rCkObvAuH7jYFaXZxf/1
rnSTrG+Csn0xuQTg1KPMKTClgQxEi4aIvsDqKOlhjTUckX+j9I7CESOIR+72V1lhtt9cip+UsC9x
JMu79uaK1KUsHFPAhHL6wa+ntYayMdAmIkpjNWNRJqMt+9JjF8Oh2VEcuXVjauShrXhVmDrfPMqt
o5wAO2rflcIifzistDqn/2Crc+EuU7R92XkJeseaP32g2ZG2y9KaKv3yr6yC9DPAI5nGCv5yqEmx
Wc5zrCJC7BEUW4lqPi2OoooYgx+F0WoopCo9y6W84YF1NOuvyi6iRX02iWxKtMa5H8mFKIzpHC3m
cTJaMvV7kepXUITuJ01gWM545LvZ2uBr4ZYs+LbVVx/msxGzWvQbrlV9cN3nheCAnlfY0M8T+t2V
bj31qaLAzc63z1R8AzGzO6djivu60wHCMuszHykXCuKoL/TwPnYuKfhsGRSkDX/kVhLFCLGcvFGd
zGk/XA6GuFjiGJyoOrzW4U/oxN/LV3KslznD0RrGNlcEFCu6VU9BvdB25lGsYzuNqrIW4npro0Zi
ClA5TIMQiydk1z5+KtBgSBkkDYXiALh6uSJvpuTf+KP7zOB0My2DsmIacooFEFG9sQfeeYsXJRVv
wB8eE7hO9vd/CEWt1pjIduPl8cMJIvRh/klAySwchqpl8oJDb7pCa5M8JZ8imXqR7xizm5wbDCIt
WTm51I4eZCXz34aQwbj7gil0p0S0XQqv08HacTvA9bUjzbhxZvPq8dlb6OWmkvca8nGMLTHuGG+N
3i8fyDlM6396UZAhHIwbCf5PcOtUeqkMpQyAKE97TjQF6SNHsFc24p8OxdbARH5UR8FjAv7Oa4Os
XS8i6gl8E8/qhyRyD3UfsWRXuL2e0APY8pk+rdnL4lWJfuw6s4AR9kBxU3u4qB7NGqZu72XsnGn2
PyRuGmPsobVlhg8OMylArJQzmNoibD3pj1IjtBZJglWWO4jLt6YC4bvmHtkFBHwW8JfuEwNMnjMq
IwrPynoEHbgA+Glh+GCtwsecsEIl0UlK9E8Mr7y7w26YEvvuV20mj10EkrRi/iIgVyMoBw0o0RXY
aprz/VGv1pMxmOvhRGJBQwkezmN3XsjtEDcOPMxPM2tGXOFRJ2/iNZYvzZ/2qOkdCMYZHzok7OdV
QkQ5sdZrD4EfETMc0Mir8WUB0QIy8dtiJEyAyTFET3Dkqd9cMLYKBGyc1fdP5vczFGRSW+qqp0gh
K0RR0jL9Q/IOQTuQQttuLzuv8hTDnFrweFA/4FJrWypBLZALYjQexm8+5kO7WfEVcBolSl5vEKcE
MOf83f3ABqNtGgTdv48n9UtcVUtQBB2tCi04gW25wz9uEmNzkg+w9tUzZ8OON8AIeSvPXIGBWFzS
fJtFiYGmYm5e+dk3a7qyDzXYBwwaBIzrNQsFTP1KHD4CoCkkSoLUZeZu37yv9jISexhw4HrbnNTB
Fe47LWv4x08jRUPGDUY6PFrUhOUgomBwTCEU7MjRyr3ot0BMjC/E3uV+rW5owJ3gRY/uGiLi9/aW
lKaLDdefctF6MrZBeipE3TypQrK04UEtGx4A/m44itVmoQdCHQon38onhMio0u8i+fG/7CsW2gNg
adR8BAskLHWm1SeKcGzU6TcLDiSsS7blpmtziX1wmEFVTFaxOYohJG80igtOZczwVOWtidBTgZbo
yU7NoumC/7LiBEkmO/UKHxWRZhtAUFzz5AsKiQw488SyNpamEbIPwtTA+ymRfucCnZUAc3QC/dZG
k8TMy1yXHJ73/1oAL15Twv3ngUd3l1IrXk5dNrZx0hmZevX/hx/rklbsT5f4Ys1W5pfb+3HsMMZb
vwswrx2yRbPxOwgnN/s9ipZT9SRS4+ezT3sTG8gjkENPEJd/bK8rS6N1TP0vjAFtNVU0GWfd6lcE
nD0qLHNRt95rcru62HuRov9zKKArA1Og8iheqj1UJUpSAD3DG5WheDdZ1oL+/RaUpwyq+iKUbaLp
FxC/LiJ6L22b+xtcZ5GANwS7Cnhfwb7irbzxaXcE8RZUjudPb+iOQ1txKSocBM5ZtGhcaK/gMQOz
NagjDIUBFCgaVY/fzmR0a1e2tfJIE1MTYZ4K3Lp2AgZrKkXXwOLXJGpDypuELikc3a8Pv3x+MKKc
7GYf9YSs/d/Z00mCuBLIQjeHyGn3TJGGY6GNYRgC0s/UtUx/1qGYsAm14839kMH27HWnqJJvNV7k
w7Yan7Z9yYAhchGEj8t5HHoh/d5chOVHTgZJnGIKxNXlva81TqPpCxP21tGBHuGj678nfNnxZELC
fqmBAwSv4CcHD0JVQTihzOsk/TyahlLeejR6pnphjfjEppExoKHr/4uTks9fA/YeD2RDCOMO8+S7
gMSWtLVjdLSh27d1+4f0I5nXsaUsZei++udQ724YAIkAYlhTUmrrH8foKuY0OPF4cRHKJjGZZuyg
ENtFe0gpfGEfKICkQvUJOZ1oGwxidCbc7ToSTQld5Wg0uyAS7q2zS7L5UIEzKyOf0LwkYSn6kgyO
35UdWwL4HAHiiF8CAO4+dk8AZssPArhAKylyLR9hkq+O0NPIfCVsrCUqekxQtzuzKWB+vItQbLRP
pQ9eeBkR76gNrvO0kh22100QGFhBn4qHqqPiQM4qgXNVctSRA4P64upuMXlhT7s3vp3jmCKqAs+C
Vqky3fqtranDCQEd83UF0zhRpqTFyTNe60i64lOvgdM7AdNJ6TmwupMKvOgKSJDB+OKyfqNwrvE4
0jzNZMxIud9NeoaQiy1ru8uzw908VImmTzTNKWcXKIG1XT3aA3pSzhgiW9wBQS0zKCYesJmoEcyN
oaLmNkkiE5CyS862+n2SCuN/9yQa+oWP79MITRjTfL82zP2orj59IEJQ32hNOq8W1I98E0cTnJTo
1Iukb6gMCzzv18JzIE8ENh4zr5PKXWlKP1HvzxFMkiRVDrYymSLzT1gMcV9a7and5DrU365f4KvH
dyOmD0PTR3Che8fmXQPrsLiQX99UBd7iHe+J6afvl79RG8x6XoNXQLr2KaFZLZ1OS8ZMazNEbQdU
yqUXzNALpgcxLPeXzh5P28NNb0ZPFLi99Zr0XJKTpxJ0V0U4ka8qfCJ64h97fUrhsCwnEuZ555qd
GPAWEZG4qzUvat7NijW7o/uF0NnPiHJXMEfRFyEKh+jFBI2QfRa5ktZXM+kIYecZNZIJ9baIXfcy
OFAGqhsd3ErWgK1Y0IGm5uqM9AOtAborP9lp2fHKLuHAfP1clZqWQVySjl+oBKC9zjiD66bDNAMh
vpt5kHrjiFU+8cL2DWSOPn7/5muFv1RVcBykVx65faKv93kj00l9tMUjse0c6LzYf5tDtdhR9ZWv
LyM/3nbnAd88pqEHQQi9UBFEWoXjEsAVukdJoKfFosNaNucR/y2URi1fW2Ek0qjBQil0WM52JxWT
ytoEcnyXUPMmXHSs9lbBSCsrZdDueiW2cwML0iu0A1k8etodHYtzIlZ9xf1jGlYxsS1oG6SGIRMe
I8HI1vF+5F7jqxvCGE94g11nAFqDaFgRLtLma23pu1X9Favwg3HYzEAF86+ychDjo8aX1KOeFdZ2
02rjVvblq7MJXbHJesGpP2sqliSNzyLDSAIn1L7ojRafj2YTB/djJSbNFwbsOlg+MnLDh9u4XgQ/
8CWKpWqgadpYXhJj4rTR1Ehd+cyBg/uhp6w4YlAVbr0hGoyEUeVbPPDDjIdoFxc7roADSf6/172l
pnWvQW5fscZ4qZmAxAyLhtPq2K7Rm1Js+PDi+iNmSDdK+Jgn4xhfIsaq83jjyzw35JTPIaHkUhFo
ut34baiutyvlMIKYqR3B6EsB+eDiFTgYuDMeHPNWj+QK6mVgy6w7qkrVlDoHgcMYzVj4hFL9mhod
ySlyW5+KZ9o462r8CkTeXVGreHdFVAaq4yEgcw32hu1hrSyvYZSLYFUlNKWWk8eD7EIV1et9i7rc
o2r3t/8ECgkzkSZcCSMMn6goizrq4okRZouiroaW4KMCV4M3kTlH8OuKbknarwkFpOUPEDNmIJC2
uNkhPgBMVrACqpAPxHGqbN1CLmXbvQ4o8J20mh9JNypyKl7S82ndB6wmGnhia+hcxkn2Lfmw0b78
fcLsN0XNgcVrTTku4yta2xOxwRuKgMhvOqtGcgHWlIVIcJFNOAiYbSAC/KGstdKzlXtmmshe7Dbm
vpmNXNtj9bGTLqmVwiDzffkN5KfIZCuLxfwn2jawfrd5yfelSzW7WgA2Nwssa6dIJBeGhIDiDsnp
QRc2GCNFMbUnTR8HXtcCQEW4WHv8OLa6/iaKooW7GXtwGytYRXWsjqc6grIXiVG5HYbcWedPbtGc
XyvGZOGXkppsMvOnNXv34WapkxhooiS3JTftRVqsXWBvMaZjgNIpW3cPE5G4hPLDfOP/KOVRoxNP
u1buMrHuMu7S+yjDCyckCfcF3Dxlq+87MVS95UJvS3TbdDuVVC/5yrybjX4yOuck0YrfZtd65Gyy
7zaGvt3tkU4pEpo48cKaOk0x/pswIfb6eCEjPj1MMG7ZryzOg+RZ76sCUaKxJtH8nXG0T9WOHE8T
J2gsqHJdYgDgDm/ogn+xqYqqGMNiE2QrVAbKKXcc+sw2ZhzkR4ZB6r/lxqwLJGwWOKuoh+fCGHnM
XCL70O7sZq24sCBNfWiKC5y8Etef5OzN6kErY31Peln2v87QXi4IUVe0xcE7yINM/lgz74F9J3J9
KQBGLu2x7nw9YIIn/EucXsn/wd6yowte+mmhA0vUZbOUgySVUFliNoH7rSzDS9rWpMRN4Iw1vBmj
BjNmD++HlX95jY3a9L2u3bgZcUJwbMCz434MkuuAiVGRLLTelo7oJteFC5Z4WYh6qt+s6Uuw9Jbf
ac4wTgcNonGVhVCm3aqkdpOFmXPAd9u4ImeH4KoIIny/OTnYK6ndS4NM5PSZ7tzUvz+691pns31T
BzC0hF35ICUiP/TM/2u3xph6p4GVLRghq3/XXhhi7xkSg4qukygKL0IH491RQXwLhqAEaRxmCtQ4
h0JoLac2plLoj/0iyjEB71Q9tM8N3nSPJctZnemqPNtPa+UODp4iXHrTL0JahwA7v73PZ3hrRqFv
vbGjD+9a1Qg5Yea7a0z7rH2Wtn3zv1gB18mkgba/vbjme3Yb3WBpSoDrmn4J+kgG06nHg2f4A/Nn
bz5to2mVt/q1vroUKDAWNeri1fOe2PIHgR+Q8zqPsQy2jL1TeIOMbxfbkPAU5EXN/NELxbocqSQJ
x3IgXEqERx7FEcAtv/q0rAFJ9l1f5h7Zyenmxd6R17mKtUJGLHmtG4WeUzzTXoEt0K8sgvlzFBL2
w25WdJuM8apu/cSquyvFLPRkV3FUmuDuYH8c30J7scBeLQlPqUFtSwh7DFOErjlVj1kvBxgGQKur
t/oQg5NxFoUO12wtECWn0LG2hN7UcT3t7MDM0DDjq7q780VfzMQG7ckd3aPCRRvVaILraILQ0XiZ
oa/Hzq6v5oZ74Ivtgy6KEASswMm4Ub+voUTXcoSNyeLTzQlnonAhSu5fX5BTtqcMgIs6a6hLrzLA
o1jeq1Wf/qoYcRS+arZPO4irrDnb12LZuiqoGuypjoBAqi9jXiriyXilZgLF/x9LtABqScCCGQSo
qJPRD9OFKAqgxD2vTvmuEydUwjAeOlCyJiWhWzFnFHk4opi2q8O93+DO2CC015D8msAtBmHNgtI4
xn5TRLUAHFI/HRRAdBS+njxE6CeNThWGZSscWGp0XIWSRvI0si/YUDtZAPu/Tc9YqA6KIgriDYET
x1SsxuQEpzq3pEmu/XMcsHqyzBB8x40gOYGQ1noL9oMeMvA63KofCr2POaZpoJ+cNoB4WSXTg/ZX
7AaNYOVNmPU5yuA2DbySszo7EHLB1nhVESM2Alq60JrgGaz168TYyfjA64k7R1hXdJbrIxGIZmjO
w9GyVhunF/CFzrg9Ot6/hkz1tR4JkRO/S0ksMwrQjL0MYNjVzRqlv4f79JEu3OfeMG3eanEDQwXW
qXLICFBWLFgHuLAIvW46b2euEf8tmXoGtva14hEJZ3V3FyE6f4vgR461IpwaO7KY8oyGFHQb54xW
VID6OhrEwJ/r7joSLDCqJSsIN/oAT1tsK4A3kw2nn/v7OCVRXIwJg0Mvtal0XtwEHsN0CyNXbLmq
/BNic2imDyfCuemIKQo/AF3AwMh4zY+mKNYWCcb/Xz4Wp7926qXsrpAfxkE5QwIq1UD3W2K67V7T
Vllkm8erTaivobbZO2Xee64yWyEDG2ba0HR9aA8LUTkKs8/z8YL5yQVlKP3uWfJOXdWz0DSiBtmk
OoKB0QkHSwKwtk6Nhgupg8H9Qhdz9Cq6Q56Ep/lJf+3wq0Vbsm00Elw006Il7MBBeARPJ3eBd8OJ
4cAUvBL6mp2KDZDT38Ey1V137cZf6REfBQ1F/eAwfxo8kynegI4JEdM/CvyBfJH/dk+SyGMRJhr8
3dsoGQkejMm75sm3ynB/KuMj0vNl+pwlIyjQeFDcdsdOBqHMnYrgFv1uc2v313yABEei6mM/TM3D
bJ2Kny9qALtka8khEs4nUiaTrKlLews7WQizm8TDJ6uckOfxndU9oIHTksihrfQN0CEcuvty5oq1
mTxZuvkRHqhyARkeuZMGA4SzKtnPlq3DL+TD4tGnoY169kQ7W5SpZcyXUXGuMSvvQsLk6OM7Q5et
0V9p0RQtOkXxyMgz/rDyyO+blE4cOijPEBhxfuh3gUQ41GsbUUzw2VPy88FVvDvo7hfBuIP52Fmv
KzKyhzCslchF6cB8lA0ekunhVkGuBVIwePgFm18nrMgovS4utsZ9VhQVKL1V2ALQEYWkUEoFHR6G
grlt379LKQjjAZexauInFZxCWxY94s67kqIMG1yjQH9DlW33F3leXfCUw3E/rRjWWGjGIxwpWq5s
yXRmPgXCTirEfKmesmgFfgBw0j9MsXAj0fCxA4TcMR+dFUGhBzl7IfUqW3jOzfIAgwD12mVxXvlY
JxMlzvA6HbU25SMfZDaeZNj4rd8+VVOI1KgXLFPYxvEquLKunbD+iGHFK5xm7iGKXQULkw5zDHN+
0KRRD/fDqGKj/uqdrazeTyx/bY6g13nBKcVWRcLmK379ZVltUCy8OTgDGiXaKOQU1wcsrgSphPkf
XBu+dlTgVpK4ymDer6buCGAk7uEGJYS0hv2hENostpgo+2SrryoS8MvHX5bdroVMqZ6rygG2xNAG
E5BjghJM0n3HfvGRV+P6UZJhnw1q3jJHga1eVEdyb8l0EyfNVzV+9kk/M2yLDczwZ9kMMNEkKp6Y
+zT6brmUUqGbGs1aHXBtmg5kxku/6SyjmQi2qyuhVaqrMIyu7ZPShP61WCr82//yTOVOfUlWn/Ws
AZV7ilof7w+VdK0mo88DmQM0FOt4TvZq+qJHkqgLRon/4+qFABjZiwkeQwEDQDnvOHtD1vY3c8e9
JuCvB0FBoMXTIdn1hVz4wX8qebtkWxFQDL5cb4sN2PkXGtYctWNqlD9ZBDXo2d2glrzQuUWL03wT
viGi+d7/keQoTF42idNKDsnq2JL/yuwy9bDpDhsCult85iWhtepCl8tpg7umwz7GyqOOzEF5uQpN
iz4cas+9USrjE5E7mjbkKG5aLQS6ml/4UiW0ScvU0qRXiH3KFQZHa+9F5Op2pmHy/AP7jXa/IlIi
AQDRAHJSpkNn0CG78w94hqejBJYAhqSUiLSzTAE3TLsJmu//BhXGr2Mu1Cdu86aUmkRWei4lYUfO
tkr6Hp3YcHV7IOi8e5O0pr8kPBb7sVKFOdaW0wkriNR1sjTzjszp+7k4SGRk5GL40TAvOX84YvnS
UdXfiwW0Dl0s8I5/PG/Rbos6emuQ30Mfsx5MqVgIPYU/V98fcWsAo52igFbubQNAObphSZ8FlXhX
N8OweINDia+IcNdTmar3tApDjH8awrU3rqI9EGJkpxeuKCIAyagMwU85z8+FgNv2naISAX8y1GSD
IxXEBwgHZFskINqW5JWAfrf3wmnch3PlR/n4eB3Fv24EwIAKkyK0LBmQx6DG45GPu1A4kRcAJP2p
7f4hNBz9jyI2zPnq/Zcv1hjPtcmYhUK9x9H/I+CgjNTp25/acHZFv6zOfJDbkXkOEx/m8hfGO84x
j6HVvo8B8sQzVzpUze0uwDMUVVHoxxjAwluLM34+QJmywIGsBRDG2zVNlEIZvMVjm8ix2RQODh5Z
RYoib9K0AX1U1QTIoKy4E7jEuyXTPVIGRqHdSlyse3/ZdpXlLN2gZs8/0HIAOuQr8LtbgUqxoA1A
J/5jL73eBE0q+M24likPfG4yNGxC7GNwApqcUIbUqgX2ZV2ZEQoqCB+dhvShwZUyZo9WgO8arBHm
Oa+020p07Ks5BQDgt1yIuv2G6ZbWl+JIg7EsRTAUH59u4ncBLn1TZwByHtgdBkTz30DTaaSZq+Pq
C11yzmwz+uxK3TQT3rmSc4E8+Ovsk4lGnNubYklOE/GyJaGFKT35TEOqVyZD5q9f71ARTKe2ID+j
ifBz0C/ivQQX4OARuN3iZM20T03+DAlSLoVyBwljo+Xcbwt95SH4/HgJdZVXZJYAAMGTH09wylxE
pChMz2Qc/qAOsiaDr2nb6HT92rws/j4unQMiIgXHO7fM7zxaf2fCxouwJB8KcXs5XgQLGE4m4oeL
U/QixbPv4gST3dMmw5+Vk5q/+f23+2tWn+7/AQN8QX9NV9B5fTAiwQUXWud+0IiZKgswTpEe+lWa
CdbTwny323ZVZP+n6WQzAnfZzI8mGrSC/K9/MW50XFAJTdTi3/Eny9nr58oX5nTXJQHlOk34osFz
g6bfVz/WoPWki/36GlchGcuFn4sLfDDPULczZsaH4ttN8juH+pM13nFuSV60BbzdQwRWTBCMOIpS
wgXbqubecVEcZyov8/XmVa3/6yGR0p0aba1MO7cjBKrz6mj7ndkMBtlrn9ZvnqZjIz3hj0NVlxpV
sxQlzEdwfpjvxn2+tgbTD7BAhFj7590b3+jdRmBhA4pDHB2O+vghyE2eWTGuxpAvvNvXvDoTuI5u
AXKm4hv3/lhOHBWyOg8xUB56iAL7fs1TWyolb15uGf4JfQ5+c+JwGL4m2r0C7uUjQ5Mdc7AUpxhX
gvmxUqVe6jyhvQ6nfYWVQJk0tz0ixrt/1I/dDgNvoiPVr2TeBSM0ModQ03e7mnghX6XXBq4leGni
YMwsdbbgbNlwfQRCF29iRovSJXAamRnwj6eFEgij/r2XQ+giivA3GZ6grj49kPu1rgqk13Tf0aOy
e0OGnCGIQ06drEwZ//vEMfdTCEBhGGiDrg2FajcrnI6QJfp/AQ7/EVNoq+VmpfrpBBYnvpkXSGED
4MZA0UXX70dq/eWcuPMG9cfKHbXIX+9CpHWtDm/82FKROhTyQpy3whlk85nV4OHeO1MCmufoehAY
dmovBD2KV8cqmb2ENDOXWiHSTnC1/dMa/c9PE0b067mG9a2Haw9kPHmggTTRW0jgu4E7+ynKA/Bc
/HRpDvtlZHZ32opShhWNnUJjtSpjBRDQSRANP4ueV+Ao8SrshqnlTThMl3eLCPB3f9+jO/iD5lQ7
Gr54v65dmf+kSEltUCb+b82vwW+JRymXhUz/xEF6DNXIsmyFadNUrR9eKwS5YQ8BEv2XDnlDVH/V
BNfbW2YVEYq535fDNK+AtEQ5NKd1RCGCX8j+DVwNcSeh2fslBBY6Z2Nq4hXpvSMCaHLCsLeLIFPn
s4IC0jXD/iHcyBffmJwDvwxgteEyTnWInvQBLjwZ76RjZ4oA3nY3W+2q6TInn6AQM2O8C4Bu48Tg
F7RoNoIB9UgTBnVDFgPRtJ2CMjXycwd/MJhs7B5ta0Wi4tRlPvnXI1QOzUIjeVDW2GT4YbvbZtEX
ENSSY4n7w0IWpe4PfEyl/AwgvMqJq7zJc11nrewvP3oZYpAachU9uAyUe7kuzZh1kkxktVv0BNSx
tCLkLj75crtG/1K1g9F3YaWWQd1LhTOkZXhjpvZ6Hay6dKXWXg6/UeqT27UolIniFmQA19pSc5PL
ViDNsGcCRUhvqMpb3ZKsm57OMPkhXQ4U/5RrwWG0SXh9i8MCKnNqNP/MYeZmjv8pa9UWKlylWD05
TDS30qcZpJDvGgvPaBVOlXSpU+aKXoxk+N7M7bpizAgAItXU2NrEJCXAMjNXjS0zgvvK5p/hg2j0
q43c/kPxAiFXhjdQOYPeaqR2EMoWXcQzUFtHoHCCkK7+Gmh32cCdClKdY/wykoI9Dxdus8PtfNon
nSc+E0Ph3uwZ1pMwMp/GGwrnLV/wcUcHBs8NDp9jVphQtBNW3wiL116D94D9TnqcAw/B0vnzA3KW
qDoSWBaLSdZJRmkIzoQ5zUTQgLTRJjPTI4U3LLc1tm38e6XDgAIQB+l7Q7c8HofOxlIt/iwJP/Ie
XCRB/T8IbwiqbMl7DOReDaSDcSo7HQhJjwvbUo8M8DDTKM/79YUJmeBtV0BP7qXGAtFxs8w9C1e4
KwkOdxhS1s/IuAHhcGk0DWjrPye94qj+iskewTDWLcHnoUQi33vkjHFQcEiw9WWV32p+n15AIrLU
xdkIWDoL6hIh0c4aIT6O8bgVMr6bATwNAGzfUOVUBvBGNIWoY2nt0195DiBgdTcwGNgz5Mh6IkhK
R3k4V7H9PgxJc2e+F2vmr8mpMMjUm8oRp0jxqYqj4lZMFG/ngbEDPdncGr5xdLDnzt8kqamRGcuu
WburyhpuYRFwOtgoc6vOUzYuwsk2vR01WK7TZMQgvm6Axrz9BnLDiFIjvPsIxwv4SWzKKPe3HyZu
Tfz2Dv2zsNU/a9BC9o+CbqzWjH0B21NJGUcXjjFczF9w8zzcbNH/Ff/+Qu/0UXzvA5Eb75Sydusn
L5yzR2hFouoGqjMjp/visRT0qfBjx3ulzRh6jP/ZbnBMO7zfdP4SxKsJQ9kawAlQK6TwLbiswBf3
xA4xloI5tZyEysQu2Zh3YD1gMkcgfoN+/vpPgRAmwAtsXEhYt++SeNVPkXPFpmVgTbY4tCWY8GOP
OPNF2JoV60OJEzB3ogqJKxXbIqaxzpQmo7G4xBthX+Ee1bnmsvAoCu2Rh3vSCsvS/0VjtE/+gBdm
60mhSbE9P7uJRwmgGDuOGPEo0VeXKXvQlHSBZl4vLSv2OTWylI0gxOKSKYPGD01LrKi1VlzJC0CI
DoFZaL9tloIUQuRYBzlHU/hW0MBwsR6bW46bFBATWA8kRQ53KHxkxFMzK6K52pIuGKmH6qUtaXZP
vwCIvur8CF/Z6+hpbrp/Yspbk8/1NX0xWZ43Grftpz4YhBem+I69S+aI4bvN84W/omERdtNTXcYO
4ZaN4/et4tUdQzyv/wjQknlSep3KLtHWx2jE6iuo/VkslzPAqstgW9B1LQUQ5dcNPjDG4Uqlr9JA
DOz4uYmXjxx/07mQuowjiwNP90+mScNy6NfXEzTszFqYJoek6N8A1GkCxBd8WC7bfqYzHPQRUh5q
EyaCTEdG8DNEcSDhAULQjSyTSTHQnvHuT45XZGNnH6It3ruM/R50fbXRgBdJzvcGSaJ7iigYMR8V
vwwzNEVUogAm4PmOpxiwFWV0rZO9obovnmNMCFXaqpeqzf0URDPAc9cVF7V4tZGlmqoRm6XIW5up
CoEhWqXw6xcEZFCMyadWHih8APwJVfkmyh01u69uEiL7cRcjAV8BBLlU96HB9HoEHmJon6YdNgWr
uvFq+HPJwX9QRLr9zt5JgfD+qV3QeAg+jTuON0dRiJaeaKUY1FNSL1berHYbZmsMjZEF+1HbpT17
I4zgkKjhoMCgS7HbTTjeDGSlgACQB47G2SqHqHg5ltmNqixX/XE1S5UZle7kiv2vyWz9MEGoxtO0
f3jdlJenGW1hpwf5YYOnSz1Fu8crh3yudUZ6aQJaoJSMRY2yYIv7pvIyFPYM2hsKmCklMtLqEZO2
qnL1LqMYupZJtf1l6f3mM70kBqKFf59UiHf6LUKhgrLOO/N7y/Ot2ZqVDa+5pVaSRmNYi6JiOlmV
vRBTpqLdkLO8I3ZF+ssXNUx04FhPPJhYGKIgGwunEs83gCOslHqbO46VjR0FxNk5+QK09zsD6h6A
yVz/QRnS+3VsM0FFl4vktPkJOtxPC+uqCQw3kH7TbF16fXPQxHq2gw7lTksnDS8jh1DaLxX4dcij
Kc60zw8jeK/ylKbtSs7UgiDc6t/IE2yXm1g+o2cfAfqQnfZLX1afVWmN326ucRRMJsOzxqTNONDH
j3vLwsuDRRVfUC/A2quku78zf04/XS3rA1B/0joX9m5ErXS/82YRekH18AQ9/4FhlGUxIAaIvGHD
mtqni9nwboAmY9OPqUnMYVIe4YmA7EYpE3e3dElwl8dQBqlJDVu7HfVxZjzlfGIt75S42NH0N0y5
OqE6slbcBUdXdrrt3alvXr4uzdW36txNUGDhWecz8Dw+u+kiblo8/DpWLEfo6K2/buQKomOqznuS
SKz8ugxDmtosq1pWPVryrUKT6Gm9W7A6W5DwsRT0fx9FCxS+CEoHGJ15Xqf8vpJOuotM8qWlZUjK
OTbQNcqrVZZMRmKWJfejIY0jYQ4+ejQcesIkxwNL4VR76OthcE5GqvjUqkXUixAaZUjbaGO3n3CJ
MPv86yIIYeIpNzvzv342RT4yGwvYh3/S8sesREANwuLMawunZZymiR2DL2r4cx1xfyz9XGIUvW1g
hCRilYP8fYAVtH243e0F78gtA5O/tiG98gDCnmvv70bz0ZalqmImbMjTnp1dldKr5bU1fJR9dUiV
JoBxm8QM8eE8SPNzr7bNjzM+hCftIsS/e3NR+ztH+fwRplZEWWJnjXCv07q9hEc9qnHXa8aoAOHm
uZxjxfcTCr/x07U8tpdSBP/qNJ34V8S+cyO3dmeHRYj3kX7CKykKVxfRwyNAw44w9Q+wUKSvvJ4s
vL6Z6GcrU10tYQXnD+lUFaNOH4hKPvByYZ50wVeGGiunvSYvCYHR33itt30NPvRwEgo0QoIWPcnJ
+R4IuMvxFDTNsNnzHkdekmS7SWGhYZl4FNhYkwNQMJjrM+O1T6HQTIj1vzu5ooOTvLJYjWl4s658
VDqeXBgNwPhHmm4H6zXReaYKiV5OUiIe0j7w+EJMC7ajvsZYfEdrFSdaNm9kqO6mSsCNg6ahrPma
W17DSZ9J4pLboyVEh46oqw2pu+qEJRqdlCMXGCnwuepTC7X0ze3Cm1XYKDgmabDGr0o7obntw6Nl
7xR135O93wkcaoNw452QotVbAOUFBdfaUhjsfDpqk9coYcZj4qF0GWS0nGlW6BQhv57IEn5zos4f
hXrERC7Zwj1HK/TnUj6L1c/NebmsLECjaAgmkauWE1VUpCAMm/vrDQGfgyYD3MygPpozlUWBKKzR
r/bM41sr5lCa4ZVl3Sn5CEdE/pitLjeGuQWf5zIm8fal+B1vjeXqD0OWJxuXPvB0dTtNRR/+sdFe
IRiXukG+K/eX/Y7Mt3dmSjw8LwY/bzn14lcJwVv+t9vlaqUV18zJAwCf/oyGr/RAN7FM23pZzU/7
HVGboSK802bVEMCOtz/x+5/uBAZS45dIbBz24G63vjiEIP3RR1JJ5KOwIw6R3wnz0Kd4J/1BF8Dx
1+9XUBQFdd0lEICMUduqr5wt21/dmyOMZ7UtXI6x15poiclQ9CFSEfYc8hwNLYyQ2vr4eUryLyOH
UEjFs/LFfCbSc8GQB3XYjOS0TgGn0QqFkuV4BdB4laM+dWeG7lJuaaIWPRWaZvzQp8cO7F40yF1j
uLhe0X7kB4n7IP03pjHVdzIkLZ1zgS1g8wGIn9Fjq8ZT16xe2P02GkK6x2spU4W7Dc6imkFjR6+F
L2E7hd7EkYx7MNPWM3sVbniiXJmqWdTgsvX8lj5sjR7SqPlxFGXm4yTkCJwi6tb4KrEQw7X7rMDP
ZkppDlQxv8oRA9RI/QAo2VSSI0HQuwpOPpk41EZBKfnvRKCQy+u13kK87SILeGjSEcc+dcImVK3c
rNNBIHDkiulE2tIGZAIwiKkdLQ3JZQPnT8lYXeHMR98ssHfwKbxWL0jLE8JwksCqsnOqlLc7nd8d
1s1jWMiG+mOucT3DY6i0cL33gdMiHxCbxHXTZL5CROoyV8pndqBp29A6gyb9x7ULYW+l3ZjimgK0
Ac9O5rCn+hJS3KbAUk10+Hlo7O0smlW1yyUvtu3fq6605lnpERtMJQ4NPG34KKSLj+FSFRsZrmyD
KxiQc2KXyfDccHoNL7fQbeyitsDhw8xYGKPVidHy5WllQ+ktMZM7MkESBaIzQNDY1N9aH1ETwiar
9uFj6vP6UpaOojpM3ezChZIowcYCkk3KlQmTpPUiLp2X1O31p6umWuqmCGGJW7QDbWD8O56o5BML
gudgTqcHVxvSfRkSz7+Jn6D69lGF0M7oTkhNzIAx+uRB/UnYU4md93fluNdgX0k5sq/HSl9gM+4U
VvTDR6qKLnFZ1ysV/vuyr32d/XPBQn49WfdTDimrluKy/TAkRMv199oPvFWtsWNTQk3bjIvcXlDg
6QayPeghC/bRvCWJEi+PwEzYIrohF5YHuSf9W9FzTjjTQ3xZeJbrctQqszV1nL9oWn3TmT0YvGsH
FPW1sQgfYW1453bo69ILmlrLx71OwyZH27cEW4LetiSGkxmqL+k7mvao3NCfuCPqNWmeOGJz9+Q9
OS5rdNBBn9px0O+DrGqUDQzPzrnh3920Ma1Ws0ZY3me/ecidMPyvtBwXE5AlgVz99ZRFfzb1uve5
yGQeUPpWpQp7SeKNkPomcmi4BpUaLJqtGd8zeC7zdXJF19PpQuhQlY/89MKU0XkdQzel+v8ul3wF
50l5CsM8PWZFd1mKhGjGs+Po04JfajQbG7PkCq0ql3JJZaqiPBxQsFPfYsZ6rEVZHBCJOby6h1PN
FdgOXRC86fRwX0v5CTs0LYIhZHvvrKeqDsbX2NMAfvHvoq0uBmCukEVbPv0Az/9pN9cvuIzxm+br
pPTcH66qRLt6cAYL5+YoOtXlKLQEG7Wb9MzHm4nCmVqHQTehuQMXXG+u5NlJgsa2UXqbQgrBqRHm
IyWnUPrZY8W0TpAVffUoOrmPAv0ZPTrHJPC4AN5AuR2dFR0qQ9Hj+McbvFaN7n3LfIX77jabBmTv
rId4gZRuUtcbampn9pSfhSUThFcl3FHn8UdjMSPF5dfty2VmetKg0Sj/4QYj6pMmUNFrjK87X4bz
GqEfBeRBhSzu4QJL+j91jc7Crdz4x7dnDGXTMVuP7z/tl0rimMhqe3dbKb4D2fHms29lDErrauMz
s7b1JJ5UmTrDBAoBBrWgxDtLFFmuWmryXqu8ajKlCPr8OKQQQrqpGf0QUIlx6iirTCXdMUj0Jvtw
5UgTYRKDElSsSsDD8ERAPMH8T2b20Sq4a2R0RFKO94vuLkJzRrXSRd6PLm6WJ1z3Z5vvRpSYm6pc
2S5eWx+pKlBrF/mopxpoUV4SsTm8OPUUgJT2oihz8si3iNdvswfXKkNaRK5zsyPKPrXyJaWCCGpH
4JwdAgDoo94mgbR7SM5EmMnwnxLgSuG6oJmNUskVbylHCWQPfOwRewBIXO1L3I6zU0LLgbxQ+spD
2iRbjEYIM/Iocz5Bx2D/WdWcOcYMyHHuI0MugJZVCdJWHya9MbMrnGLoGSo5BoJG2T0o10tpUWdR
lBYO0BRENpjjVC1NJxFfIj0Pmr0LOy6ftrcheHhym7NdZlCr7D5oT1QQbLjlRINsBhLGZrqidOze
LVByhZBA/q3cp4e/N8W+90Cdsac3SssEdptm9gUIPnUrp+if1vKmiA/pYqCFmuuvkzWzzLa0KDx3
6MVrwcnO+xseUezTQZlOMjCdPVz72BIcdkYTPtRcZuDB/jZvXokgSM3Mie3yW2HNzCzModOvRAMI
/2zHvjU7NXk8JcbItiCcFAMOa17bJIS83QPMr+MlyPvACwui0pQXqLJt7lkNSo3wKfY9cH13EWjf
NFq/bdRN0XrUfyF94U42qwKOp/gfL6surxL+4XOmcUyy1EyRTze5FKFbTEyuyYkPJUiFsbDD2nNY
ynSpCBJa0Kf3ylRWq7ONB9d76BeosPmdj6lJBr6ks0ZBzgq2kELKP0v7n6sSOazFbmGPBXgoiN1d
lHt6yt+FIxq3j0vr/uMPYopSI8dm5SxFOMO1uW9JMkkpYZLMdsXy638jD6NkbBiDwTbxJYhJgEr7
e8m2YF6360lkCKV9FkZo5gJh1AMcKUk0tD9JrByURtOR9/iwTE3y8RVlCTfZp/IDea0GJCUG5+Ps
EeHSsJV5vI8wcArLS9j8cXDYe3HC7pKQf2FKTYfN6ZCUVb0b/FghFbK/HmcSNa6SeXo5cVedG7qF
79riG3t1odTfeLY3SDNM+gjAdWgSzeShSxDKBYO7F3SVcQf1bN+WgNFFy3guQwRjkfqHP9I+7TdV
W02LBw5czD6XVckURPMcVzECNrWK2mxu4QoMoCjlhlClpElA0p7FBf6DbmLcA2WsStOkUxVsRHXt
c7adqYP1ziyTlOp6g2v+JVGj4+omEfgrUaitW+kxrDBvJ1NfTCYCsrsVs/U/nB3GcgvcDmen72Tl
0fhrLI4xbEOz9fUu29d8MeLNIQdbX50CdsZcfiu5i1PpUskJvk/r0V0wmkBFm8uvXGvwwFyYQTmT
uhb+JkNZON2vAe+o+0zJb6UwBMBsIeyA/c0sNyC7Qc7ogp536aI9oENP4Vo4hjXH+hRePanpFItc
62Gal09X0HNP7FU/s6nv1q8PA/nh4+gmKR+rAjBTw2kmhBMctHFIDV1FsIFQWFpkmV5bMWXbOd0A
5QD+seSrtKcz+BvAd40heahh9zl2eh6eVRTpqtiNYfKY9+gy1jM7oOAbIyonEtroGkBNyuiEYrs6
+oxsi3MxMY1ORfb2UduPUz0ziLEuCGeH8qf3sKRhkNWZlV/KXpozDrg4cwhNhmOMpVQ5I4s4sQqs
cQJh5N3ZiWt5f0TBZ9IlQR6wJbQesjsnuZQsEWl+nN/K4So7H+tI0ePt3As/W4I59PBl+hYbeCNO
2BXiJV0+zwvP6PVh7tQhwc9fMJO+lyQJcgQhEpZIbtnPfUJN7Z5uzi66kmAWnBkMVOl113SDweKc
tApG0NUko4z4VLgy7oZtJ4GAWvt7Pa6fC9L0K6fEN7xfZrjp6auvlmAQMwg0okNaz3R54YqSMOr5
mKkX02JG3a5DmET9evCWPb6IaNXFzhYdP+o9KkdGv5q7kE1ekCmEV9spcMAJvJCWHQM42GRO7Fca
PQamQnN2JCmQ3ZuBQ7euB7FxV7OISx9tFPlqI/Xdq095jQeMrvmnAIOlKSWG4aEoVhAit7A2mk7I
K9lQ/NF3DIJoF/o4UcDsafPzwSDY2Wq6PdLhkvRBiXZNv1F5Wa9QDu1wP1u16eelMettgv6uw44e
nQKv2/uRGfy41c6lAwhtc8HlvC2/fwaX3F9KYpTfd6n3OwDxk3JQIgGYGd9bviUKdCgwimY+gYon
K6AvuEvINsjx0o2GS35jVngPVY9OZs50A5QI1hBNJC1mSyv3uWiDclxkGp5CRB9Wf5GoXpJA9rPs
tgeKKiDAbL1YtGRozS6DEQUVRN/d+3Ih+tNnYQ8fupNyIVqVYLaVUp0BEPsZuTEn82BXtugqP+lI
5dKjKIdoTXEX6lsnJN3X5gz8VHh2insoO5A/h/+qLLhCwdUMpcsU95/v1+Cwe4bbrNWP7Mll9Wgz
W8urireJeq0SgU2y51AbaFw/Sntl+2/0hfNrMRM+XLbLj9iTMwVlFc3azNaxjPMXTQC5LqJduNcm
tbBEUAMg1XylJfTK/G1l0N0dPWIAG1E7J4MKMqeB0aTAZ0PDoCb4XIW8g5M9hFvPptVfi3okSaS9
GKRPT6XfMiWH+rdiUm7A/lQXQ6HyfN51iWjmupG5n15eH/+dHUu+aF3mdvK/viPCfthi68muLHgW
p1/fxd1BF2kIqAOFxCdaA9YjYXvdW+EDFucU4+9asIIdRL2dnmpekdAoGobchlWK2dp9Z/ESTw9A
NLQlJkFI348J3nviOSHhCarBilih94MhPIv68ffa6oYV91sK7o0EIxKAJhrq9iSsgu3XCxNE7YuU
uO8w6S1GeumQs8NcGFP2zwUVWsnmIykhbXzUToo9FEBW9ap7WJcbdt3+7UxGxvEunKBfUnKoenZD
/slQtXYw1lMDn8AYRUd6ZkTEuOteBJz8yigFHLRhfy3MRjyLzUMqgA1oJdOM1Ur1FNXjKnG49xOT
RYFXr9F7NUnVzbw2hOuj34QlRLkgZ/5k2ifyIkCeGqFjRizihqXp07HiHr5vuqB104bcs3Xo+smL
Vm9Zp2wYkpYFmVPGoWjY47euFmkmVTojFJIvHVxU8zJ3waV6Nojye6zdI0elnhH7SWEDWjwizFKA
bLbI2gj4y8FmaNW+1OHSDRQXKG58Pacfj3WhntM87tfIvxCZGyasA28xkgh5JZrU1QRXmMLJ9Ond
CiIwuxPNcZh76MU0yBOSuykO+LfdIcXCkYLfT0ZxbNGd/PYhtZq6WM8IHiFgdd6SnoTcE5XyilNo
Gut0Zds6Gz91NKWVGMse2WtpT7TXbzV2QUTH4CC7DuFVR6l/oy3NUfMlfJgLTZnjH2dhxtRgNYdk
9O7srq4tr6hD7r6wqJ5CSL5KYL1ksbNv6V+3MMnVeIqOfrSgLTKlsOj5lCKE49UiDsarM5fkdi+s
DFSVj28kqgq02e/CqpdsyxKbI+7SkclC3QOpbhDgqyzy2O81kP0h75OpHw5RrW+5ZPeKchP4iTDM
BdUzU7UHBImiJbhbVOEmjIqtU3S5IiEMKhRGAgyHyOpecAKkkbuifg6+K6PgCCsEsXhqqijM+DmJ
qWMWE+rOEZ+jW+TAI9UP3vQ8A0Q9evilmqPDGV2/L/CJyVuFQJUfATM0ah/O6OF2DuGi8GlXuNaR
NNGmq6IrN5KLhXNYZvpFc7kcpftGDsOsBYhGTejfYbxbf4hKesET3e5lz6F85kXbHBT7Lcu9/4YV
F1HYlrRAxa3tKMVJrEEstUtHXvL7IEKEgh39WI3UnRTGft8V+F79hVJpjWzVwqHWcGpCtpQIUlzA
g7+4xs+2AQOWe3VYNMyS8HjYoYFFBewRkoBrCmjpWUXwrxUF6Bd7c4CIpdK+8UYoKm98qcVzTD1L
oikyQ85P8TJmor00ynuG5QPb674dXkJSXXb8HLovX0bQ/87Xfr/Ra6u6wpvIc+tq+3UHAFGP+pgs
QgoQxxJ953kRV3udPc+kLW2BuFOZkfMZbQjNzXGnMvr2oyWekj8rXrmOd1aIxokhBYpuiqzKkzhA
v4m7b/ZGoUC/ZkkiaQM52Xrbup8LXkFx5oR4wveISTeqAHjvey8TnKejDdecc9nkdM3JpauptQC8
x7+FkcYK6j3g8J8V9UaRSp8rkPU8jx7V00GFHvml0ZrzB1MdI7DAk4hRCXtJCjMtYdqTTPr+BS2F
XQQ3ziyPp6TbaReEBJ1pWHCJOIufeYm1IaBHOhmzXwFqazPdWiB/8/0AvzsBozToFULJnquOL1Ey
mNkS95vjq1yv36yM3f5syhzjksV/wA84dO8uUxNlaQp0+CApPDWiPF/CxHUcFzHUglBhIHrBGu0L
wu4iWlgcLpoYNKFDAVqEvD8+ZBNBjgOwoi2ksQ3nJJTeV2n31TBeiRg1ER6HV9z1HpVkoO0pvkzv
aUnH4EqydVVWP43xL2xr8V+5JtKoREofu4fWqPYbj6Bh88we8/zmhXWbQsp+XQCrwONlNoCkH00G
a2AdVicjGi0W7PT9Z28VDqiANUOF0TR6x0y/gtq5koTy+u0nTOqxFUKnh314j2KE5TTjHkXhZ+MF
fqoRq3C1KZm6YW1PfUbxNLKadsPg6JpdSnKc1J1lLziGf3uxK+gV7PQh+5zBN52q7dK+tJYnjfII
cAAgjjyx1oLtpeWGxNjNjdraTamdXzbXrNn4f4lkWqOvn92LEqHwUkBWAI3IiaHOXFz6gUemP8O0
ihWAwuCmAP3azxyD+0oKEyg8t1wh1PFcrxaUdXPNcnMX48uwMAa+Jkhpc9UrMCuDQtCthKlXlLZe
2jy2BfrR1jO7AwgglogWDpSnW4ZEI6l7Bp5EKgpatXkpuQJ08u1aqFtsn5sBuCe0MLTxDXwtNfK3
YyM0lD6NjT8Zvb335DJ6GX+maKjy5KOHcsN6qbc+D2SyQsUBelGb0bHN82eaDE0iHA/X6G8NcPNK
iGXFOphXTUmnS9ka7K6gON+2hU0KXbHcevE7a4dNKBJI5ya9lYC5Z8XKXnmkOTamavpuVmZ0lp54
TiWrpm3+5tcvhsM+nklROv1meGNPnEL88CoelgkPZ5mYRrvYfEbxDjo7cxOrAe8JbOinDTkhj6OH
+9wm+vkt1bTyXphTC8NhUEoUlDQso4AJ3T+BcYdutAaAxHmyp2UuyBn8A+5mEhfreaLjjg+oykDt
PWrg9nDCcOCmi2mtqSi02dbzsjuU5lXwyKpOoCJukFaNi9w+3XICns6+2KPGDgNEQ3/sdpSWlYKl
ZzQF+FKqTHjNoYq02wF0XmUY4EYVh/fO5VCL+51+9i5D8RXprsKEu6f8SJp0ExkgbGxDnbtN7woZ
M7W3UclptUctKbmETd60Xxh62RVcM26pC0IwPMuThp8ImU+U8I050F6mcvx0hzVRKe0k7GVx+1t5
9xynU2WXLQNlK+9es+tmO8ZR+kA1a3ODU6skeH4qXCZMSxOIuIhRwrgH6qsLKWTKMEQpKfIXIKiT
rLAxGD1nBBFpwW8zN5fT1yQKZ64Qq5JYxVqSA8aiYx5Lbl2Cawtj0VZA73UUn9iCYWGjdae5aPiL
SKLjl/VXWsZasTu/MNkoMAo2v73/kx2ZoaGjG7dYmARh4paHOvQ3jAR3FqFQuTO7yba1gzgLXCHY
AJ6FM8qmIM9dMELbB1RjOTPuIq4JQPjbj8PufodQ+hjb5pZBXkAP2jQsdTlRn8HFk3otbzhkrsJv
qcjKY1D8kuWqkkHsyCgTvdDi8nJW/xGAbhvpCGSxwTSXoqlFM+loz0TbusKcQXZcZa8qUIMzW2Bi
k1oK1HOxtavW3uCp+hLJ1ZplNvXY9nR4BKUcm/dLawf1pL7/l7OUDWAUcJEbwotm5Z3GnB/8xq8d
NOIhugyO30M7g4efy0NO1EBKFN0yS1XCqv/6X89RoM2KZZKiO16DflO7Fb6te7XpnbE6K1vSMlKe
Wmuu4Ha4KayfA2TV5HkhmzzLWONqUjbpjZTSzjphPjFOMVWJGDoF1fEb0jnMXHfbFvXjfLnEKJR/
Wj3xfHkjNOTk+apOFBPTz8XFqW+9BM94bNd89//nhO83whhAGgS21GoOSW3geHzeHwuti+yUvV+u
ZtUQR4hK+egKZiAo1B+yzViQlaBFm2UqB9CJxiJQE026/SCYnt5sC3bGKTycxvRmRhj6hXLchmDR
c9ro6VFMP54SF4W1fN5i5XxKjTAITg1lsHaJK7nwb6SnqQFLLNfPi7f+kUG4oxssXw5xUW90xNn1
6D3DCXyq2FAwlJVoRfO3SQ58LThxtNvd+7gTxm43w16KY+XGOANwyuu3yMenJ4E3L/HIv8dyZrez
J2Rr3+0VwzUjfpapjSs9FwCJk+dAT1jpOWOB79nt78uwLidAA2qgJ4xVTD//OepcfjElkL8wVtqs
RLBcv22sTB3OkLDah+XGHA7hQwIhQAX30BDZmXBq0KbtDmzsDu6fwAlM6k9r5gMx1Mq/O1qcnUfM
2fA/l52pTuku3+vb9pI81+Np0surOLD62U58xph6sg3djCJbldwFRrZyZN6+ZVtoySzbzafLOTd/
DNKpeJtOt4z1EOA4gp1cugJ+lCplOe6+Kta6UF4/VWX20pw7B+Dl6XLs2tyr3MMHow6CptEbqfpb
qzC+bW6qpRq2c5XprLiXK/mMdy4iBT2JN/C0wJ8EaX2UeLKg5+pX/NRjWKFXg1iiTZWxCHUN50qs
VYIQupu8H0ERQcPuB6HGQ7ehcWFX4Pgn0UVio7XbirjkcCaaj4P9h2rUbQlykom3ituw7/LPXD3M
HxuM4ygsjAgcCVy4szwuY6pznVQavE8fXbqO/Zx4/EDGRnN+tFPpy4Tyrxf8CO8dpQZVtTMNbKy4
3tlhOywJhdlZJmluebTlTTk/OhGvZ/O7ki6bYolKak4DTOY3tx4j9lHAEkUtL34i+V8gMTl3nkF+
y8Yf70x7NnyXJf0w4nsFEx6P7ZskNrlnzFJRE4Pn8thZMtSRcibwvAeQJkohRQ9tECdb9cytQmqQ
GBZK2xKqxMOsGJ96IvWXssrKbSwC1KzQQ6CbOt+hXolbPCmr9c4oW92EEywUAuQw/DAws9ZrnC6I
Yh6r5ZHAiqyt10L8RccUpdgTsR55SL23IJgcpojD7uylh0RI5EyMiiolTpPd8SEP+kCVnxkfrVxq
+E6WOC6ddekPB13nYL0DsJ12ge8Ik9Rl07pLDsK+KjH4mIPUNpKI3ifUk+6bdvzr177hflKFIQQa
f3RdRCWczLbc1WSRoX3XZqcA9UYafbYnskT+Hl2KroXkTJiih2jRKyrwON9eYBQbCeuvSPlLfe+W
ag3D+ZnuQ+eW7C7lamkAj+LQ97tlbxeZO95Wja0/fzaaG6nHo3rWTDjei5dLZqK/fZXXYvMYltEW
R8bTN/Svwh8ThCF9MGO9wNSG1aCtsgSBQ86Mv4l/yuTBxdXRA70wbql49fZiE6Jl9lto1u6vD/ye
lc6itr94YIYclqKgucjHVBSaaA0fd/biuwu6rCiRzhTJlat7L5qc9G6AQCfkrswuJCl3Gf3BPYRD
o7uKlOU1ZAreuTLdlXYzSHa+HdcsK1oRjgAuw+qmoz9oDibL0Z2qgpUW2nfnOF/3qQpMH2aFmbgV
jdzPkdRF2G9qyEeSurRRBF/+70lml7SKZo1Zmt/yUz0gfLcyjYNyJea5BqDCNJx1uv8YatOeEtbB
ibb30Lq87mSwCTSXNJTloiBFFRgu/f5Rx+ycz+2sm96Mys0HZFZ2nBSq7t5uAm2GI6llMkgRkQdz
rW6AxmTFxRlr7YjKXGXkUsxesPf6avlzO78FQcisXLiueMNZxLMDX3fMLGtqZaV+3rDjOHvCqmaN
fzQ0qPnZVlmI3riY5roaR7AOLvWqyQOu/3PVh1aG2JIM1WlquvRkuv0osX4Hyvn2OMy6OTvz6lTC
C48DcnzZ9ZLIejIJcSObIRTe84S/yIz51tRoMs0GSFywx2jf9jOorR5xLnHMMtHcp1cQ6HdTXmj+
ULcmNe9f895eGOKU7lJ3dZudm7wKAl83bo651S1H9/8pObJjHt0ehwkeKolKF0aytHgFkeqg7xqP
ufpdR+FgMgFTvfSfBCGffn9iKVyNp9OmOIY9oGT2Ncnbb09MpgaxF2uiJRneMuPq8nj53pdRtqrl
R/A6J/FmnGcl90NWPP6LBRJs3PbNWT0V9jK1V4TfuxPXOmhgy/pq+Vnp+f9ZigE9zfL/PzkEFduk
2NS0/LVLJT8/k5aOkfJcnUFceC7OWRk1ZkgYqPXXzv+Tzmz+mYkuTLyDlIBHCjrrpcG7WSPR/17k
QeaY/We0yKRAHTuVyhqFNYie73Lqhjmuima7SJCTSPkYz/HwYa+k9u5t0N8IoovUPTGPiM71lf4q
S1ps3SlU33BCl4dzpGF4cRgHjAEpkGGAo7XpEsQxs5d9O+f2kjmcvT3REqjlz7dcVVLov0Ytxnd0
FdjY6qyKdClR0bJBT44iyy7M1TN3hsTSflAWseEPaux5EL8oiOywsmi6XnJDyqg34nzX966TOFEg
lwSgyQuCDrSutPveXtHyXIVNUM+n1uPZcsOQHO+3WqF+9fJpObFGjZg/DGTF6P1Ubh+3g9cMlig6
/kTBdETKFARsud+D8tv47IN7wXCMrBBb8zZCLo12T9wvZDp2lhoUkzVuk8R0HAn5zrd16OFUyjjx
ztt7drIgr33t+mg7VsHXo2Hr8RoYUpAPyYM6wpbOXzhz9dSlPmIGd4qCvrXFNORoDJtoo+KwTHdi
3nzxznUTtiyqu9FMomxVSjfh9sQTEcAEp06yZEiWrlPDQp/Ad1UMeVFlPGyf/F5AgudV/CorVwHF
K4ovXnLD9ZW1/a7iWpGq/CUsBSxsgB4BQNRC87zBzkU5TGZ5n42dKlOsM9h1yVGU3NK4RRjRyXO7
SEo/9ddt5/9XXLZltwZPvM7seuqeZPv8zCetODbM+83Nh9rhkkaW6/DGSp8+ax8Xj35l+z8DSmtL
h11B/xaeshtYBYwG63nHI6Lw+1I9hmz4lL89OgeBV60hB9uHn/Jfy2eLNB9jXeFAOYgtCDE2wOP6
BRQQ3Sn7z7W/MqJ1PeOijRJkZFkuN9mz6pQCY/2dtcSgfc22Hp0i3ulolYu3kFOudNeoqKYEI2Lf
MtdH7lQ+EJvtH3lxGolYOkcUGbvRFBGG9nMK+vP1l+sUnxqfi1Gvy9sd/jqDVsLpklnQTtR6L6iZ
nrMclrrBPIOHdFCgtFp3iMFRqtx/ZUfKettanR7pBKeflYp2GOSsCzRhRAQPHwcOS0uE0IFTpy//
xcM0cGGXnb10hFu76qHzO7fVwGZdQ+jjFDX8eZHJ8lN6IKE/QkRCRvE5xOMYLne2INVj7UJbOzz9
AWLRClGe6lpUbMZNBP7YrJm3rUMI8Tz6Uh42ftgKmMSu8vclmoKXcVIM9xWzHDyGrWMmBOwipza3
tf01DDFRXlm6zdHbHqigMbq8UyJaiqeD3B8pDSJPsp/c7DEYvexaPpcwhwJyguKjkWwLCCsaSeG0
LMx5yA6+n8jThyfjsRFhb9S1eklr6cqbK1Z9XE657fFSzvYrgJZ/Gl1R69j5SySS91J4CGzNhV7s
jbnllzUAhbMEdkNRIQAFGfGmtH7s3xMArjfK+l4hJ3Gvjn2ZEm/FSn7hH+9I8c/6+jEoDbeMfHeE
1SwFcelL7m+z15DlTg3SRuU1SuzBl7kpYbZJhafGACB28YapE4k1mYJpCn1F22hKkZSYEY3mhEgm
+quibS/FpuDQz7y68HEoDam9Vfj9Hpv2GmqlNlFnd2IoMghgX0kksL34yYjm0sigKEadlLnvMX0m
O6VQ+6to9m6fFKvXOPemrPfXzAToIaqxn89pmSmzsFWWPPk8p+RrF+JZWZZ7aAg1TqsCmfbUdyHQ
MWtEKL80B+qdPbSdUL8CyjKZB5VkD+clVyJeDgLqadahKvxN9dCQSCdMgjxEaRqtMu7J+Hxz7b/D
pqe6mTk4S1GqYAmmvZLNFyW+Lban2GG8jUOUMqZPoPS+hZhJxE133zhz7uiAFcBs9+7k8B8H60vN
vRv9oMap9aJ6GcTDS/ixHf4+5MG3IsShPYFQJMMggtjQPgW3C9DB0fnRPVz2WTTMv4mC9LAZ+5BU
AaOin6ZZQgNgL2CBPKtOKaxJb6SMXJqSVy5AxloPMM0lSHlqWSla6NPDLIs6I+G5eihsMjGVGkNY
a4jmIarsF5IF9JUnGOGL6eIOgsaDWmYrth9pp2hvjToMsPh2X9lquYGDMW5Ka9tqvAcBpt3zurMA
sL3mVvofOKbI35L0HW1vRGvOconwqzVkIgXGCCfREz/vwGcG5DBowehtlRpoYV5dYqs9eNF4A01S
fDJ+s/5BvFjTB8Hegrg9MDF6FrqzrlcBt786RMZwglvCFSMoIvTaytSasv+XeunaO3ljFE+0JFV5
LgdeRs3A+P0nU4u2DL5nUuzscy86Y0kCmkjI1d9flB49FaA2gEA/uchrZwQoTxR6bK7GDpAbsXr/
kefHzy2i3+pxnOCPkUuzSvBgn4hKOvY9xCbwqBzmOL699m+Ff8Q8FXGVJ+/xVgfRegkownNKu2HN
kEO4vbpMZaHshn/ez04V6HO+8e50eeer3HqS6/RR4xQNtWqCK31ye2zZHXxPtbu3obqJwfVjzDzS
BmwFmLbEESR+h+m/ERILMx6iXpCqsFYD3MMvYwTv84OY7nIdUQWrGiaDBKb2544HSDwnVt/Qw+/M
w4FDtQDGSc/CXJjypdiOlZI8p1NnvjiVmcyU/JemrXlktyXbVDiPAAwKs71tCYB4ScC7gcw4Fs8Q
5itt84H3o6qbKU4sPAhhhgx7Uu0kaEJ2kTjJam+/D9JYpjq9v6CitIWdDil8EGAYlNxk9f1RbyRC
Z/1Elh/Nh3cG6eFrzUlGZE2loYjXdoHl2zCbU2JYwQLBAEnFdMUquMJOoMf5oM3iu4AKBX5xgmnp
czFL17PxGfb413QPgHYhZWhXtx20s7bcu14x/yyYFwdPJNSZxDKRASH8fn8MzP0eGnFufHqTy3RA
0t0xrEqy6wAFuFIWOlzD7c0smIx3lGFUqLTX00RGvxQWsFHXqs0FwCS26Qptr1O5L9/gKB7PqIXn
vn9zQjef9HT+Juo4etMNPXN9ji1QKyfg+I51KM7wc4S0dZaU/VUw0hAarBaklgMMJkUlQ47/UDk+
8PDxiT5SwlDHJ6ZDOM1WzKavrPmQQXONWWaPsuVFX3T/Nl87XmU8fhzS7jrq1iPk8JsRIM4ysx5/
/7ViNUDqq3GJpw+Shxa8IqGTChz1KWnyZCafpc9AtOqQYokqr+qAnEdSoUtkrsRdp5rWOobnokIu
geKM2V/uhF8fB+kDt/irYUZ1kj0Pin6hxLoUj4maxggjUQSbEk8T/NIehKLtdX4Yc0TtfJLlzFFp
kXXoiOyaFD9gNUdz0Vhx7cyfljlKtWxbXfQww/F9gfOTML1ybGf7BXEw1kHmibGqVgWk8bTTFu0y
CFnZQpRHHHltquLwwFqUov9lJJnVqjeJ2An80IFkQ2Q+tVxbNWpcIQQKS47CF2xiMCR2js9OihcR
7vJjihap+DqQK4AVlg/BVZtZXXPniMmlp8SWB/n4mfekGxxW5auRqW7YIYTfQvpZbBglv4TRAjNp
IQxkwL2RqFU20yOiZFPhFe4JOOzKl4VJzSgtTkaurNsdDdu05rjpjTK5pGnotl7jwiLRD2PEwM0j
Hkm6XMFDWz4TdSopoV9ETgvBmsoQU2i96PRd/Hb7P9kBfsFZIbWz68Aa20qTtgwKZIS+B9uX8ka6
7E9UlPFlasph17RtuutpERRlWHSS3WFXkyU44nkdPZKmVyTjlpXcnEL9k+H+17t9U51nJXhLmc3L
seke3waIoxszlRA2Z3pkcSq5vjZDfG+EpSC6uP1saNTW91lTFBsEbfdSr4MglcrXogWLHzVBcom+
hOp8Hv2iweMP4YK+a/ecl97hkse6hj3pbIf8HENIwa17wzcaKXLKmZusp9C7YEYgcy8zAMAGbYgb
CMetpTkrtrLfI0CquKistnnqTTgpB6xbwc1XlLWOmV0xHGEjGtNaIjY2IdRLyqPSeKCtMg1HF1aR
L4utSfToJ8wXQrKfoZwThXVJ6S4HFtfa/Mva4y4AnHUGJ9SlYQeZjNsLXq9fRzkcvyssLfjdGJjv
LhslZ4kRiFYBYykzEIDvIsFazw2m3rIM/3BgnLY5cP+GbIhXUveITQIqpOrCsEGezSdCjg/SQ9Xv
AC5PnmwUubxqh1HkTu9Qi2RQUlHOM/f0K9OVQG5xMH/i3HTdq5LkcGZtYXtQmWAUs3GhCk7Y5zwL
G/ry+NxWJ5yX469UYaHkHDPvTcWdUsgErs2ZJddmU3+91/ZK/GDm5NiJsy0eCICDedhSQEOE2zPi
3yixJ38DfFeWML0PJfimIDfd5dFwAXX/dv9BKes8Bl2nvv5XHnRulAdY8ID9mZDg4ZgqoktmgvcV
bwZxOZU4DRsrAKvj1q/xYOByHaoBt6vKqvi3ARbAoGaQktQZltmjXdgGYTpFIfySSfx2xyFdzMcc
6iuU/DoJ1I8cDbG3ERk6fZxqFUb7cWkQYENWIO/eh3Uh2Fws1sFMZEuZdSY0KCE0KvGtVzRSeA3f
fAvOvME/FSpsVxNonkLhIyxRUh/vXSbnraaCygXXixfkse62yaHYKxcq0PbKsxM/y9okUzZnFISh
fZisXcO7wEAerqqdiQBwCzfZpQQQ1kpxyEphUgWXvE46J9HOOF6KAcgcCjXRXk+nu1UG+T/X51uj
bPDxWgKC5IDpwvY8VWCQ9lg8RL5KkgQGEcqZch9Tpvvoqc0nbFq8TtojWroisnjd9qdtf/BZVO5E
qnHyBEz7nBXA3lRKJVDKijYVBy+tnMpMOFoCnM+eLz8vntbr9yV1JwJjJfobUWq2pamDgkpamIpZ
oIpSddvndscPeG10tja7gOzl5oXwOrud1TUVbQPupWQa2FZ7NjqNqizTNj2bnVsTOp1e+X8sjJoy
lfl8g1KdQp3cNXwUIHriPY/oca7xBUXXNEjmohVhEDaibwbzQ4fZGv2vuTVkS2CM9IR3wEAE/67V
Gra4RoBnYSJGilShKOmiDdagupYjCfdbcw8+1S0xo5PmwGH4uVToq8op2Qg7ZHGnycZrfZcKChXg
iHor2IXODkcgLfrr2/8mG1P2Haf9g9hGWUVi1breYLWHzoHekwIb2bWq6YoDPrSWUPoWhTUsrMfs
pCnp+iqt2KSqLTXBavFj4i8J8Qui4DlxnJ50KL5NUwSVA2BYooiMYJFbr0xeeNHm4iieWnYrkBka
W2dNO+x/WX6VaNfbEFhg2o9mguLJLSuUGlIJZoy9heSRGJCMmJktnwp6opmM5vSm/P85kOlfaZRu
5o3a/2tECbIBPyrAqcSQKf1CDiW6gzkcmfDGgRGpr4jj52uP3eep31VmilnaqNPEWnz28paqcoVq
hb/U3p7QAkjuDCaS2QwUsx7QWtiwwtkfdicNIJDKfsEAFSBV1WxZxKFfdspnaSwyj90Py4RjsJBL
3yQWqvoBsVoRWTGYymNHIWGOCH/9raEIACzboCKb/xMkJZyhdJPNV2GCR9VefrCw378ZMxormyko
ccDIFY37A7bX7ipMWfFK2hIBHVb7IOQDDWPspM9dyAKCf3MT2Uu3MON1de0rODi4Q9oz+Ab86iT3
+vGN8HFxYw/fwfpmP+mq50KTpzYR6x9eiODgwY0Y+vKYwCFzVZW+H+t/aMkIqE9jPpjzny7udRSw
dq0EoAiWWRTI4lKXfFR69G7rC0YtyFjiH3xPJD5gbFh+2Im2DOx2lHNpSwaK6t/N9+lKXMe0FpgT
/7aieQZ90ZE2KvPjqXm89VHHBsPVjt0865si3DizkjPzOy3cGXpJ7bfp6YMd8eGnNyf8PlglVMxO
9Ea0xehQGJpGqMtmcJ8SJ0Sat8ZMPdC1l/Yd0X7IAWGRT3vIv9TUOB593TxNBai7EVnxcENmydJ5
mrLCpf7HyGlhkVm1wZ/l80u1F7EI+pBLZXVdZtuyewV71qsIU3JQl5xNR2IjErgjMTc5gnQjwfye
HAhR6esUu+GAb5e3ql2oD/0LMMWUOLyuzFy2SXzyH7tthmKZmro1l+IFWrY33hPf0jlnXGneRCO2
xjV2o+NiwSMcr/qSWKavi3Wb2Ep8S4JjFWA/igPLeXWv3fshcKzx09NZA1WoZFyjgvLs1IY4ZNr/
HbyXI4IITchZ3jv6p8jhasDpRkfsSqOLb1FLCpUdhcZdN+aCofjTjtXxQKhExtu1n95gwRSpj9Hp
zzUqTlWcpRfY0y7wbtWxaI1ZP0KS8AHqyu8gNWUUfANJ9nISmuf6pLrlzQHc4MfYUBvw9Gt1DKc3
dLEOnGcCXtU8lBfsUxQy1jpdnJba0ZOxLAR//U1Wa9a6bZ5kuPaiCZNwvLXJ/lymYEXUWFu0QDTl
Ow7CL+OhqspzV0BbbfxXSH51HTIDgykxYR6HG/1eN9SwJrSTdsICK729Gk9+BQUNwIQyTff2wZIW
BnIaN8JYlRwM8M/8w6sB1COGKeXSj+KS3b+TwMjUkENSbmqrp9fUekvzZhQAv6AF+Csfgi9EWp6V
lhuDx0bb7SW2BO9J7WG5m7Pst834PJkWBajxcjY1Ef8eKcRUqWz9IL7MxxtyyyaPt8X1J9GBB4zB
/BpBpPGIL7n8eBk/F3msYghzm4wQBeIrRoZCNdRRFfT9fSatOl0tBiCXK+X7p/CBgt37fjHKrPsU
C0y9TEine61v0vF+KNgFHHDKHDu4qfSuepj13wwGm6uv0l1MX7PdzJnOCeBmJj2s6rOSCPXQ/7Do
PCxzD5H3ncgml/CiM6jLBBCPbn6fFSJ5bhIKgN+zOhTSCc7T2xF2MlvV+B+gbU2xil2m4a0jnS6k
4VuOAAst6IRGoHOrk890ThvTtBnBoS0feJQ2R/GhNuiBvEhq/dNDIwOVnNZsPuf0a5US5Ggef4w9
8FGGAzRNca42iAJJIAPqTqcVtaCw0KPtQ7eGy0lHUEGCCR4O5DwpDWXY1PH8CQg+LOEJ/XSzRNfa
sFDiLoh2vOPN1Abguu3MWwkOERea3XCDhF8z8ySL8uM5Mwlt1iiN6StI2U7lkBKkDS+T+jUMMVur
O1JaJejnhXnTBoNW8zTvaf67EVJ7nnRg+QNmH2vDOXUhF03Fia+pp4mQ5RwKHgtLBT/m6TM/O3gi
Su64oJZ1ZShJgrEI4g24D1yMzhW4HITIOCUIwm0b/eLvYFvOrGYcUusnINu3LP26CqrjITyEGr5e
LUJq35GHd+JZ9Lqi0yz682TSCp8RDwvK3Sekqi73d6FXTpieMQxYjMG/G3fa9gsDONkIFRd//iGV
1aH89KoFuuN2kQ/eycCUoL1yfayVGz6wG5h6Vihdv2s752Ux0fLddI5FKIau5hlbRRgEHSRJNRro
OlUVF4N/8vlYBRVnIoW/qnigXribAlNjh0aBe7RhtVDsJGBTXXeg0nS1vPlp9+JHNgE38L1k12um
qKFhwJrVnWPE1BYEzt8+ICJKhIwSg9rP4sWYF5qDxISFkxKHisvAPyLBY+29eY69lmyrrvH+s6KQ
hYEHzdXP8kKNMedfNWgpzUbf8URHb0VOpmlhrPqOGufEakU8h7qthspbS086N4d3fN4kOMTEjvAv
bR1KLqi4BN1TPjGAnx5WShq0gtKNtJRDIs50G6dQ251FudQvuiB1X9yYr5y2oe2FjbCIm5hZhJrR
gX/hgGNN4f0RdCkspCZIWNHJQSozll/16K1XwHNsW74W6I2XDhRXJ+I9E+ee8VJXIRzEa5AHCDPs
UytZFL1bqpHNofa9IYXMBLdG0+GmlD9bYl3lcyVABfoziXGNKKYOmyehHMQwH4OxrTXLBGwD5eSr
hngEsko3Pgti/NV/JLIpo1b0nOqUDJhjUTBGpF0O5kN9QTPdsrLUW/HkCOxTSjzN0HYom4tq2Lqg
l9NNIYwmgBMY1ir+3bXRqKRr1NoEz5Lqmy2XOVa6PSZm7UCJ6FiMb5DhkmfqI3FpyI7Z6psjzxjH
54N9L+0qqN4T8RO3vCb9TQTfJNboQjIpT6ZxFwa6a9ZhPr/6IeUIDKOGv9CC1NvtKlnJGvgbp77S
sZRDyZ/UNPWWQVaeAGrxcamTDZ0WwsbcRkCYNpizmP9Kb2nsWn8OTXiPrr/Gp+xFSiu6T/mKni86
/KgQFcG+fu/8CBLLalwYH0nktp6/kPuSAX7Uuo5WHoecuHRrrmztN3YmnFFzTySCufZP0CBLrobt
UbFHjDGAKjodYDFLa0l3fY4/e6HEynTx9YmuKC4V/u9BLhSvSEbZiueuyIPB7Gfq/o8Ou+g1lGmc
ykznynrwPoRRmXDAAqgePx8JVCUIdr0/rIlFssJJGurU/UUn6C4rKZ2JIltb4fL+I2iTzBc4ACZx
nCg/bdN38I7cNyU6QCnpfNixZKhG8CvbCj4ZicBGIZ40RaDStT2yYv5jY3dg1dUWe0ijPr4LjA1+
CUfMdF2A9jGVSfwgtLSeksNBUtPgomv4vZJGWLU307/plebKxblVxTDebXScmf3WB4JQIN169aQT
KyiBMuEyPf+73gcJZoQ0vWkElIYQPxmbuoIKL6V25zuKl/EvW0mqcmRc3pzWaG47rzMXZiBhMwAg
RvtiFLn/lRkPtH9RhUDuLyiP/rWtAdKQLK/gft2yH8U9C2A2dcP5of4MD/ef0k3G8UHgYDoB95Iw
j5EOMGf8H+Kq+CWsfjLByL1EgCelUbFWfGyyZvfjTBCreSv4d2jLcNB29BcUQ1CM5IpUp++0Xi0B
BtQtldZN/ivOm0xa72JbhHwSAKmrCmVRyKMNwgrjoz5Hp2ZaMzZ+D6QNpdJ5ospyLaYVQQHuRXbZ
BHKc8u4hhsoqvvGnWNBxcH70vs1wTC9hJNtUWSQW4ufRkxugMG/uPKzP1/EpHabUKzCJa1/0kOlN
PBxhIjcwe4799x8ky50mnkOktlBjR0TcpoPJP5N37GcDxRKiyX3izpqNSlIhqgFJ2903Iwx7bn9f
KVjfX2PXSyoXmNPz9wklxdjnKwV89TIekRTBFexr/wjhO0foe7kmiZJSMb29yQnBO2+z8HKssMnb
fEW8uaftJLpEwN/GOBeDWviNZjF1Zpj7RdoFuvBFbf+fEVUZjboTdcZH11YXYmYRnzFmRE1izUJ4
iTX9yPcFfhqPS8gN+nhwo8ucBooFRDbixXC8rfyoPSwH/R9xkRR5CQzAT650Ug2YzfMs51z42dln
ZAvFPllqTy8pZX77Bx8UVeM1bI2fEYpGekMFobdFffY474zJdSeNuR8ILp2+wxMio6KH0koKyI17
WVqdWtTkkilqhsqj62N+ZJ/y9FiIACKokD0j5/fevSoFk4vWeRQI0Ln5cV0O+6wJrn/U3BSR0VXM
1yysQulpY5v6xvQrl5xBy64hQr5ntxpyUNkF1oRNKd6Un1ZTgMsC1gaVp6n5NU5uGpJc1cCT9/Iw
d6RUSeCH+XI28+JC7FWsSMAmF+Zml7kxhIHZ395wpYqvPAXW22+XH2Fl8IXcGoT+fWqPF46PY6zs
PJUGTPlSRiRo24sCzVT+TtrWse6JkQhWkLSVAKyzpsfSSI0K9dafTA15Kdo9a/d5DFrUj56RELrm
faeuVPBHrVOSj/ee0iWrIy1CBmmxsHbu1vO/vpuLQC0gZrtXuD78i4hTmIyihmBRLdVUHspZQRuA
G2c7PdKhkvstSNNVN1H75Pko9MX36yUmqQMkssGitc9sD9aBKLfm3+oOLk9aLyWQbgwHe24ScZwX
RZSPZoUxQcV/W7v65Sav88eJE9WFJf9dagDH0JLeSvUDeQjE9CJjE9qE0948IaeLrLyziDqcHoZv
ljlnu7Cp+rw+tXUuvb13mwAOeQ5iTWhNyDOn/skijiwVvh0WjlaD2bMu2iVLfKyMP/KNj8kWP+bf
ho0VuxZDfv+pnrWwDljkR3zBphy2VY515W+17E1yvlHz4QKsjmpNEZ2qGyUuefn/WT/nfEO2q5Be
4gmAPQspYgcYsBO3AMsUJfi3wvq5rrsG41F0PVx+m/Uo6+OhIAxFbQMLC5a+WPjKK03IBDPlOpWy
4Ah7zLZ0qS89vYs28vxmdyTEWkGRP/Y/c5sCLC4loT6FUlcJ53gavBL50dtk7EsTxJFV927B5zig
aV/zqXU4SeyUx77M4K8nRXGLxoIpp91n6z0JJAm2rprLLmH/uNhK9ak08i+W3yDnw0mlBvE4MmRh
pZ09VEeI86mGvJagUOTygB9FDYeaBPWnaMSc5t387YTes8SuNXftjFAkkiCFxO7FB7+z6iYruNSr
Jb1BhlpLQj4OmA2x16xsW+2Mbv5ZuLVBpMBnKJpbcvqRB5VxFctDJkiJfIJWxGTIqMslxbV0v6Ce
OohdKlKvwmxY4HKeGlcSdJuDlyPTGVkyqR36hNFNuhfiQIBoaF6kqleTkiTJAclzwxXePl8Wnc2Y
iKGUwHbwaG9C+soJWc6uihVXTU3k+823ulv8LJMWtI61JCP4e1/DKkZHs8Oc69qtPGmCWz5E2Ofx
XrwlQEQFMUbVslqsWqtnu24Tz4P6//BuGbYOLsO52dqJKAKdcg7VWtwI9mOTsmhGqkEYufCOvVYy
hzPcKFHTMXqDLk7vMU3xcuANaexKi+3INak0ijBeBSrpAYTGToVz9Fk3Hni4PF3jsrNi0DQxsOhT
YLdUfKjIWrAbAKqDCkVBvubvU7ipxBQjaFt4wu1oaQVZKxeXNxoq55RA7qsqnXHlFAUUOqP+O4gc
WB+6qQHm/jjZaP5hR7J2VMv7GfYU6yY0DBMiv713y7jYrEciOlEZle5qF8xnKN4tAmoQm6o8sEkY
wzikIFXxo+Yz1CCkHi85OuAYw4RaY9UuNWsFnuBRP10CJrUdnMSRi2ZCkmYRZ5pOIiLioR/nJBw3
Q0OsH8YDbnt3NddPsY+hnGmI+9B3mfsSzXz4Wax6SDFQBRGJeRTD8QoV05L/s2/sfBcS2IWzctH9
pFrar7ZTa9g47y2yKk7YUkdws5OvIK1EE/YN8/sW0CCVTZN9KyI4TW7CTkQZtlLjP9H8b8f0UtGK
PKcl5WyErC/DrVSR5+nMKD42TB3hDsB3KeNw0E/1oJNC397mKi8zVMh27w9ZejwCE5e4n1E4Nfw6
xIHN+OLGnbnmBzmRRc8f373nM8gde57NDkQdktuwy8pUaE7X6fJYW7bvQu6ts84MUDpOfy+Y96yZ
DNP2VoCxs8qReJTziGXV3KR6R8T7tSLeIpqeoHo3vj6NljwtHSJ4YjjNMb+clZEjBGxb6lAZ1aKj
YJLGYCuvtyNLPcdg9Ts3B+72/gA5+CMFEL+K1zHM2IwLjxOQZhBGtohvc4CwEVr9yTbEKdcSafLB
x88EDB6ZeItP5VugT1Ytgvs8POqV1z+sa5YzJ3idF6OTb8lIna5i5L3dnvgDLOOxHNhgtJzFROuB
hAL91QtP2HL9owo0LG1c98IgX6lImQF0NditM3tAka/2iVbyYD9kyQoFP6yE6GbOdmEQ/Qo/MgDM
cr4wRXdYaaRwLkJtiDI2EMR+4g47lhnLXYnh8am7Av5ITlPbusJVDU16GVKUNQGQv9nAXdttKWIc
sEzPVl/Ck5aAw1zuG4i5e5vr+U0PMSRLTuzNNZNi+TnSzZ/xR6RPl1EDmjGTQo4vWqdRnMNpS1cS
exz9waAUzcqQag8umFq3w+KBHDW4Er+tQe4vF1vhKC9jYN9hQ8mTQHUfpnZ5S3qW6VFfc8GVGxZi
VBfvfD3rl3mlwMKZ7PXL+wb7jMZ4tDhTxXkqorWq0gocf7MtaBYGzJrHPjtE9Sw7Wrm0jIQNJTKE
1xf+3HVsctWGW3b/HqGSj/1DsUyv30wYuJbJ7XLLxUtAJYy6Vl3Sg7hOeN7O1oT0ps1I7YKYCyZS
x4uCcQ5+R76+zfoVMPUfFdH2ZESC+D68cjNxPjvnx/G6e/kaQSX5TQEF/dNej9YD/pLHdOX+aSxc
4lfTGewELm0aGGz+6DkbRuFQyIXStPCqUCiup14EfOMJetX1yqE1yaUNP2vpGkmUjstNrQTpldLm
p8CFiA7JXpaueQ2703T3NhKuvFyd07b80Q3hpkvU7hERNX0eZpKksPrS8Qx0oniyMHU44gxxAxEA
Gc3WZmAJMH/lEVIW7JVH0a3qGT67KmPLVS+oodXMbvWTdJQ/+1vOI+f5Xvffnq+ebYMq48SMvSvQ
Yta9z/NLrUnxqXTUjjrM6e3IhUjYvb/UdoAT3CdDqpJjqT1Yz0yTLt6QqJUlWHon2bHSsIj5IZTV
CNuB3EKgJPGespzEc0Tt3xolJDIQVFg/cRyeLT5Z1mALUSFqT6fsX/x4HYXFJwM95Q3qXHYnfpfF
6O5pwkTqhwo8KVMZ95Pbaf2kUIALDOvAJimdE8Jwdgopa8f7oWjFmOfx7kh9ToPwXnS3azbcVBF2
4muPlggRfJprGD5H9lUIztkGe8ixLvaQpLaqNrionVK+j1aNxp3Krne+c/iGG/b3C6XZqusLukB7
z2/9YqxvZdY3KqL7cp63HnXvOoBvtk1SdNyudQ1HEjZRzTdgmhirKG/Wlaur5MDZzUa5b2HqnWzl
NkkLZP6asVhT6LHxqUWzrJeHTPvCo2JMZ02ehjSFheV3zEl2pga4CMrsuGYMEwRDKfVwK99y1TcB
pQiBCci4mI8mHpejXoHKZ6DBWQ2AvgWrg1Zk1RZ9foVPlHRzNm4eVVd88NsbiFZmJqVoaMmv+Bci
WlKS95QpQDiv0hzV0A8Bl+GfR+7L34mZyNM8KXpYZJWhdFaQtTcahMTKSZHxu48JlIHNTPXuHiJA
zFFEkGAoP85T0mr8blUAwnU1KbL9/o3RpwGXlxsxRR773rENTxCeZxsVUBn28SExnWuDnF3QAt3p
KA8wLsSmqhXDQe+cLftXANDuMW8kmWDJHxr1SG+tn1X8bNd0uwWGcdNShz9iFUUDExySTWLxXVWC
zFg2RxsQ6XL4DoJysjVIKIhQUIuPGkacb45J06uD0ZIhhKnqW/Vf8F6ohrUXB5z2ZNedEgAV5j2X
ySz5Z1k3ONnevYMIUC4G64BFuMv73P0fo1OCff4NGp9ry7yNI4crrYu4enKOmMhKTi8PqJ1VqzOY
Na/nK6maV/qUL1fLInDtTtjX2XOk2VYt9XK0zvtSnv8xQlW4dZVXmYm3FLFkWJ3ozalmrhS/7M0W
uZtka1slOxrKdhMczvf5rekzvWpy96lCbA5C71IopsvBpm0BdbXsnX7yv0O0Y0x39XKMZ6TNoDGo
/5NX7Q/FQguyHGxFKlM7VLIyCr9WfLaCw8OsENahWJP1W9V9MVHVsr4TIJFe2CGDkRt9HPfu57nC
XI/fS8HqvexFDc3olQQERPWk3DbTeok19lCxqtMq3xZOObSk4DXg/+qCU9Hy8w6IGtaIhW1AXwLw
Zr2cTEh7jd7tTdK94UB1lm4u1R2NiP141vM8XpWlFi4RaX1rPrQ9R8SaxAnv1BKImcNflJAZ0pct
9/dp9sDmA9EUBZRs5Y+sL5KmZHKarsimSS/BZ/xIwrm6uwplGvr7phgFm+RcRTrUS6+UOEAkGbYY
icLY3adpnmBU/jG9D1ofaFhdf+jX+RK3gPSbNIKi9w5acGnrMkn6fvIA/w9nL9a5dkwfX/cOtw5w
TYt4RvVVJ0JPl1iR4wcqxpHHySPzQY/yND0UVJMcO9JDkAwNtuXXWehV+YeiVz9JZXww7vkk/Nll
vDOZtI1XEvC0dK9RFzFdaSn7i2vwkOdfmlEcQEXqDWHnvMOu+8ARlBan/iXq9fDnhD/2AN/b4th0
5seNn5dXNAGRW+J2pSXai0oTenzcdevrjM293JDoRByj4K8b8GAkVlitGFUfjjXR3fMbpywoiL/P
TPiaje1SZQwEhkrRKYM+QV2jpVRvdQwVh3cGZ2wJe94fN/RI06bH8c+OkKCcYJfXw4IvIhD0AoZ/
aQMNhIJH3y41iFc80QMkeNd9hlOf3YwtCymDZ+8G502cnVjoApU3cq3v+Q1VK65Rs50zjuaMoZqZ
KFGeqUgBikAzpePQwiF5WJSHmf2UtXVel0dJVDao9fyX5NGkb4El0/PM+cS9JJ5BtJ2569gklaE9
Wal6NDXS3z+O4msyIsEDnxcpyRhyH0mSgACnEgSiOyZDnMbeznLf262jOUw+cDrRV93oRWYnrM8C
UhOWhyMP6DsBAj1MggAToKjQxs6qjrgoUYnltmHcuRZeJTJ7wz8Vm6dbElVz7EpgDNUyWlMcUHKJ
vbhOgcrTzOhC17g96iKFqHPklh80Ufz+FajKsKC7Xrgmh0uq+TSPO0oI3/88KiRmaUa7zTpI2svf
rbWVtNbHlYTqp6tpaGqdcWOpR5j/9MUDJZSa848Gt/HFE8l6X6/jlHGqmlzHxphJwL6yfr9TTJxZ
ej1NR6hszpQIHXyMCLZMmlVydsmp4vyO7tfDUQNUx5wHfZdoM+f1DA9eVE88RLLrGq4I/wyoJ8+f
WN+/tBGq8t8eE59Sp/mmRluj6fHru7oU0uMecbsv5qrccOqef6wAyOcJCTc1DPx53wlZECromz/u
oc36FBmyzJaKBpBXB1grdJBIG1eFmUwyb9+juiBhUlg6vaLNhYuvKaL+rj+if3DkR0WYIhypD7vI
c9BfAPsizX7sK2PVBfAFXJUeOSScMSfQepg2Z5E7DcPP3/4+QubfuFcu5yhGeYO7UNndP6doK0hn
TSPD7x6G44e4KTmjjAon6FPb1A/bjmdwcBNJfDqRrNu0lyiNN6OTPdwomVwGStTktAwGGOUwRuQC
sr/sv6Yy1FL/mPMCNXz3NuXvOur11lE+U6bUiFYByiQ9yvYZh1ko6hWFPwZn6esZKY5sB08ti8hz
sVgNuQkFSrKFkhC7G9eQQ6lSxsyZzuij8MpJ42sSWnyFSktzNQRhakfc/0m8qhJS03p8V2QaBI9N
goBmbuJknR+Dcf/WyiJa4TPp6BvaASNkST6jLA7BqVHsQEjI2tRuO7ysTJ4ymN4gE44+jWNZn8MV
9fhaQrzX4UxbAeE0R/UXQt5ACWH1DemJy+JrgNKySb8gcCFSnk5MjCNySUP45BwPEannvgynqb4i
DOumxAIQWnNX/LQtVa9hpaH3iOI2rxHErqB9h9XW+SC80gbj6LLbEHp+eU61Ls+6VD6aWDtFHiiK
FsGYK5+GFyHLD6K+fpf9hOz9x6Qi3vwKWvZN49+i81ApS6P/4cMKo/sKgvmyFRliSz+AOHKTJ2L0
JbimdPeBUs94va9k382KdYxZfcghAhjJlbqfuwOhIPIGD86bj1H17l6Eoxq3ZHVVpulJHka1BagZ
gRdNR5U/3TzeGNK/nrq2nQDM5BTk2DOhtOBNy901LFP+5+1JUgmJB+snPEfx99AkyinxWACeT0o3
2iM2oPa8/ORvz4sL2hmF+qGYADDGEqq98dEs9MO6wi8uc0c9nbQGUItJ7LCFWeKg5C782cWncqY5
zeRV3OD3f5r2uUzniTo2uIB1nsFkLRInKy2Nq4C0bkA/QN+ikCPLFUtc96FzLehkZsOurh1JMzYg
qgKW1AcAiPjNQAf7X7UR0Dc2wMN7Iy3TCs1HdqL8enYmUpreBAEnUVg2X4dtUAAzh+Q9mPE2S9Vu
v3xkxJsp3lGwsDU/FzCBSrcqRQgp72Z3+ANxRBDT59gdUY6oFBDc4ilhJKpgnAqKGcEzcVZSLzQq
DV2cHI1IiRz6smU/gsPBH6oJonrPXTgOUaB7rDos2XAWwoL3OgVZCWh3YacZslyytqhFVhaIC5mS
nqJANsY7WgORo7E3NA1+IV8P02ijgeRZSBzNsw2k7dc3kJs/OJ3yhEAWvZFEdHUhBvplhRPmgEyR
3WvMtWsxTRTRTjLgWiXSCKc1fLKaKXcURARpYsTc1cPatmKhfdhbyAU3zS+JE1YroAQGtlwWbGBg
1RQ8kgrtxyElsFagLierTzT8WpCyVQAtPwRSVgiHJZgnQh6ZDyoj4kjGsUAftTqm+Ko4U7IodvJc
AZe44IY7g1PFyFZO481yYE6gHeJGSbTItLB4JQ9KnjIXODRC43BekfwUUQCG9lV+wZi1AL/GcZj+
5ko18KcdLBGGPyDNUt1QZOdODkAmVZnqfhfu5TfSYckKuGt0XISiJ0EzK8iYLtBBRZLR7F+2MaCS
mbQ3vTXYCoSCunBSlqfqYRlVlayBDfuxX7edV+5dIyrkF5CU5pom/gAJE18Pm8Vrms6QXAK8Xa5A
h04QVCnAiyp6af5yjmwZzGtZqitA3SJWxH0F1/iyMVXMLYUy9GOWZ54KJPHCUQ27Iq7Oo7nH8ZH5
2ey4OKby2ixBrN8OYbpQ0HWn4OY61/+ZwDvS5b92mN8oYzYljOveG7F+s3Mj5+yiy6jRYWkBrALH
KPVJuBU7TVy1rRPH50azcdVBhtPktQhDd49IXBdysDeKwGEOhQ3PqqQfiAF5FeZFJXXyGe1g8B5O
W/IvM44sR3aThDe2CwSAXiOtBzBKQRNyd3fW0sOsys+CYMZQ6LeDKX/sRuLUrdwaTSpGH06VP3kZ
+cdjI1ZLyhfdlH9BWlI2/HbzZnYaGrUwYbNvMQqhYw5flXwtiWXUUe1Cz/99SEe0NSO4cMcjV7FT
2TuALuiklt7RmG6usJQa6cTrrJqp5uMA/udG6KUZpvhwjBqBvEKazJTkp/luFam2nzQN/nQiTaNv
2F0Hc2bPbM16TB4Sy3EXXtCstZlfevxHQSnn5nYIpGLGW42akInTmvmoyUpRn+d/0tU+clVyYL8e
u1bjUAESOBPhDyxfgUi0iSbi246rLF3bsDSHRLB9c8j1ixnQvoT4ycT2Lcko21/8WBd6o5bfnok2
rUVvCTNL4DReUpM6rvt40aombloZtOYjWW0MHnKxcUW6NuAwUY5HGel0S+vSEpFkeCtpd9vwv4kd
DC0cfHD2q8kE8H+Dfi46icM0nP2WyYBlsyGCL8d47xrZAT9S4hxAAv1NFyQV1d9dx7mxQ7BJdADl
j5fgmpC0+oBgp3BUNMfv4kQWGjwK4KkFdjowgKHxzd/kKJDm7XiSimJhqCaCN17Q5SATcDQJdnLv
1D6gek5pltIuSfYMSRoZ1ZW3SDioAujIwpTxpmXky0IPN8yDJWmVDGmdQK0s8/Y2aBGOSa7DW/I2
mDyJwf2akpjlXy0Hm6aUX9d1kVprG6MFs6UFXyz6GbooB7NxienyIQ0rtFI1CVIeRTzh3CEVPSyH
i41l0UrMgp2YM8Jfqh/3xrdtaUSChBcMKXcjnTE3WWJnKgnkH3g9yY9TdtqaInP/RsDHEtNU5hBe
bsUNvqbyt03MXZav2WRsiB3VtF5xrPm+f4DPRJUoLcaqKkSK5SRHpypGphbrAgrqkrpjkjSVLeDX
cMFkCajBjSiv2TGS1erhxHwfhMcrnzb9GnIQ+BS2fxry9zlCzstCgTBxLQCF0s9ooxvz/rPkjkPS
cQbPZP6BmgFs2bC5P3J1IK8j7r+TRwhb66sNKgsuwd54Toe2sZyAABI+48HhY6V4ojpxvRgV4AIe
dzoh95ufpPE72IVa3FC4YeXmPeIGTXI5fiRi8rWrr5WDLHVifbwbo7ZvHW1sMNM8fEjByb5jUXmr
LOIajEBTSVLrouPewoXvqnr6TPDen2lPf95iLcGNf6TfI1b05hO8LXxWr+E58r4cRPkBTdJoLolO
t8nyejppD6UhE286cx7ElTyInc/6cCDWuYrpcXfHln0leR47caZWcGBsvPd60DWTs5yEzqBfgP8s
RndjgaVKomY5puoKaixobG0EoxNBxvmGKUjQ8lS5MYyf+OA5/K3tftvE78HaNSd+y6Z44+t5qEco
R9uHaA61FfKKFkHv73+FHa4VqY1k0CmYJ7Vf2c1rWwUGlZOkFbvrP0S1RMSW7IoLpBVftF5lSTbK
u2ksX3ZYwEG6Gl3VRlxNmXA/NpCYMKVu05VZe80Z1zobcqtsJi77qJ7B+jT6vSqFF8x2c7HiuSS7
eaqbkYM0GxLeCfSdiReRf2vzwMA3ENqVe+zSYklJdPMnpLJ1Vn3/HEZvI4hw2BWzZkJOMkP672iF
Edz4WV+GWwtTGwJFhP1B3xRsbwVepzf4kiru3AEkusEnxctw0uFKcnK87bSZot/o6GJw3L5wlKlQ
k8rXCR9ZPC+CH7q/hW6ymrU2sw2qzJg7VEo7ss2/yv7hQPo52jAq4BxdPZOc8UYUESNFmAiNzgWz
IBSHWg1SKKl3ZbQGspZcGHa8xGALyW7O+yHJyEwqkhXSLBKmsbVE8tdiDcImBeEr243yoPSczBna
aYibWiXZYCywedTzdsgFr6ygpIuBl+jNKSwUmXIxKzxgWhFq9kfkZhngCwM9/JoH/RlaqZqC0g44
cIYd2DfwLNjcBgnzsRHmrSIIf9JQ7lyOemR6CuZbnwktX2c619TOlXzM0jFGHodPLDX5qA7OZqiY
4HPLdAEGzKoKybFuLCcFIduKt/a+EUwp9f7AvYgnNFML8w5TB1tseNoHgBcmmWyQr9tx812G5gT0
dzPmMjzFiBeZG6pqUtumpIsAkbBKcw6+ThQGzyFTuYPGRUrR5IRHP7ANn5Bkpk8eUL6jGZwJUxTg
Xe/oE2aNGmoDTgoJY+2JmlTzkIevI1DHNbtCBddHhplvCSCX5i6mWANR97qCp7iDlcZnKhw/rwOk
MFAJQjYxEoAHeo+pJRbde8YOtO+6VXRJorKZMmgyMb5ZeCkEBFaGiDU+5YZjr/cqeTp8fupBdtHC
cgi4XwQ0ZfxaDD0fJICBhZu8ZTBIS7tC2yLXqQPeSE6z+LCJORZ/b0uqnaJhLGsXgMeVrqLruiSA
mjQP2IjEi8LW1mLmg9U9HrvvN6+ADlgrRFsvaKfSgvqDoArQdF/Fekc/PCh7NL8AwupZYIp16e1F
FYn0wNSa9VD6547M9juaxEAbkQARNiSpE2UDT1JOkopOzgArtJLKEb5GR1Cfb/skCRY1CytzkIM2
18jByNTV+JPMYQNIT8WpEAS6+gJl2J0G2vVn/bVfV/93Ihot8QPZrNqOQQapvfVUlQVsmJL9OkMT
5XV/hkGbJI/3l+Mp73GsohOiRuGVoFb9rKbWaf6VCOL+5nqo8qMygJGE7sx6T1aMZgJVkXVQjLE7
5E97HRPd5jEs99uSAjMgo9JFlZnau9SoeDJ8goAchb96NtQ2eTx6iOud7vzI8tAReJkI45XDHr7r
2RG8VxiPtrW/aJubC/bbYABiAZqD+DOxjPB4mUSC5+WuA15kvxh/UilYgDV5Ygd5CUnvsTuifa/4
klZHuJpcMAvgLbPqWe4SKGKBKn0K5poQK19uyih5pVS/hcoXDN2MEYiSWt7zq8BfdyUOFLenoKWK
+WgAnLyttlrVfHAV3m/S7HsGfHjH8ZBprma+kEk4ry855bG8VRmu57j/Ke9hEPRiLYX8Wmhj2mWz
FiSrfJQ1a2PxndC0zu89r58pcCCpXcu3RcrktqtYabYMDK7stOkn0xgGqHAkB/fJTWRFeZ2D5Ja6
9c8OYB1ka6Z+H9VRz01FNpW9yH2CQNwq22CBFZvgoXqY7bJAofGjS519X8m/UqOPr1YX/RXwoQF8
8Cqcyjw4XTqH5D9cKxOOvFQzYqiGjEkTlfCwq+UdERYap6sUQNsIroeCJX3ddoDYU/c1Ht8nSte1
OWPFgzOw4QVy7Mqy1Q05tP9UotxodmmRnkyv7GelFjJMvFqrv1MBumRVS71IMzS/31nzzzim9Wwp
8KqgJqnnYUVd8Lq5nbS+jXS4d2+dOisKx4kMt69l1AKnmbJ5bEmeH7KGBN8AgPHeTcqRFoyuCRBv
SW0kOKcqaewkyfojZGOwNTONBpM9RNkmfLVqZW8AADhnoOUId509oW9sFVPDiA8xsOkBuDiFK5qf
I9cyUztTTKPCAM39HZE++J4leuLP6PmI9LSApvgEC8mBxTwjOhfyVa0y4P6QQdc02rtIPm79b/R7
zCm9H4+3KN998pTsnpJazPKL6XpdEBumQ1ZSFOfsRHgZRa/jfcN+484MxMhbSZzWV+U4QwiKkzYJ
iRAisbd94ySLZyqYfEC+Lw+NqhVqKTpDyefoHFBD4k0U35d13lkq7NDHOzrYJBSNS20lE6EPvwsS
oBIcfkwbZZkr8IbxrJuFvgxGkY0cbSbcRtQY9E2mqBbqnmHDu8cWWcHAqRwairkJOdOnvU7qIML6
sMPKQbjGQ9OglskR9xD+okOVFmtmKKHBU0UDlHibUfFvuOuTpVzBROW3PPD1pzk0jBVg09cNcQFE
swmVs3iFJetbxzgu4Oe2LI/1Me6zCkfsvIt23CWGtmcmhhOR53iB6YTCaqcoOzd6naQKgQ1qSAKa
Ep94RT49vPfTj6tmE7ylsmngfoo8cRgMLgDOrItypdWUVHFfKpZCrnSeFWUW4Q8g2RNzIV+auhqY
2B5FmkOux3QD9Xg+JfIgvxVMvpm/To7bIFSc1u3VaakpM8ruj8khp+luFOShuLbGT9BWuyMrMWxf
CygBmcyD0+1UyvZ0sxR4ly4EJIt286fiNKvtcI2QxU4s0BfJrT9mH4W7I9bwAYdxCgoSX7O1H0iA
uFYkIkX8QQR7rBvxSmxR075liGiQ/H6XHH484F2YOpEafz/5cOUhBDLXBQyVUh6MLkk1tomVlxdz
gECMZK/DXC5qyrqMOR2b/Z2hGF+gcwXXHbV/XbTlCvDywWkbTTD1ogc49V7toYgt+2aCYNj7HrMx
KIYqh0i6txfqVtmPINUDiUokw+i+hYkedcLvZnDLQ8ViJhR7TbNS7tq4aV1rBCBsbsG1W0xFJ9bE
79OGhapwx69QDne4tvCMf7SNRWFPqR7jURGsond1MuFKD3RLQUF9Fqd3fd1Kcd19C9YtWwUEi4P7
T0dNAOUv/Slsbb6MgYbwwH1hU9mfWQ/MMq7vumDdjOGKeVQpGkaocLrGMpRETDoY6gXBmRQD/tjX
hL9NpfKur1jVs+rsdFJhGUiYA38FmHhnGeDVRmb933mZwbF77+oNYo2DvaHBJAnP1zY2oiFb/qMJ
uO0p5LvDm+Inf/ryoo2ySq2X1sE1gDQhNkkjWfHNM1yV1aqsLTNQuASWO3DwsegpqmdTp7jyBJCk
ja6SqYMQD+jIEtdMRC4SQUCaJ/8GDmM+AdcP6ESxDlvP79yyauyn7FSBaA6dso7cL2n9/OVM/Bk6
b2tx54g424uGtFYYxuU8G4lZHO3phpMhMH595XOQULRwEGbAfQP0yzJHAfRWcJfMSVFamUDkD8+H
jF7LaKQKj7U1QZSasGiEMaf8e+wngWXibnp72hXZ6D6GegurdhNIfPsR7xh6Y7TduLJ2TpZBUIyq
6rveVa/XMV6l0SFDHAalzpdwB3YFVufy6TarWmHBuCxfKnn0AakrsT4aik4YtFm6L0tz3YqwEXfd
iK+nhmiUsxoadGN4j3lP5Zo7kkNZN+2k5+K7SpV0O6jikxkqUP8W4jBBjvoswti1hWnkkwQHr8MA
RT8Fw7i7ZnL1T2zRCUd2b9hdUumuFkANIvE4pKCNHLh5dGsEzlYqyq1K0jUxvZ6ZU83wrafjNFQe
q3tYaZLuz2OnE6MFpoCPSeOf1pbbbQYWBuNWSDMm8HcsLPCcW7te70BOWHwar/fujj8M9MZM50+W
WER1qVq7rVcjhb9ORJRXBsA7WCXDTO4dTQw8uli1r5XGwSOU1BDxuOPwWq5NzTjJkdNQqeMLg+dE
Q9qoaCvHzTO/EByfH1c3SLsPYDgRhrp4Mzyz72L4vmodeV3gMa/3Cu2yCchGmLlEZcEl8xUVnaiM
nV97Iv0A128wRwzueSvCvC+oLnvF2027vuRFLbgsVcr9g6NHwdE2hJuCEA7QENqTeHits+jUqeYc
/72GX6uFI/6uEVJNYz2FOC08C5LYz9dMC5BhSG/DYerYuYFN2emp1TsxCKHxsZbar6cay6Jetz/D
6p9mPzmoigRDtdlYt8LosxznJkPFzPSdSjVrVrkAZF9hGEuhxJXZa6/k3Xgu/dBzsgfQeKi/2sAx
aB40dE29Q9csV1LnCxPCU3GqpmNmtb5Q9RLjVCg2TMblG4ZahfKybfxHmrZ/DUHWFBSG/VcZvLww
J5q8LUK6TVSvIW4PSmGEmG9bNyHgbf7BgoW5ern/NqvfSW5vx3AMnkBzJG8qMu6wtieoFggyC9Mk
y60ovgQv98RcUkiTTJ73Cfeuhq4CuVVjtGihhU1LwscVyNlXavyYA+EaCLhZTgfP8xT/wyPC6c/v
vq6TRs2wafFlcSHaj9rOuxtHCnE6I2yCif+v8kaoE8i6iyOps5obbjRQ0mw8i+HGkKq+cKt6FwSb
1jtEtPtENsQmtt+c4lnhOheBYJ3dz9ud8tjY90mu0uP1gnsT/Whjf1S1JC6ZQcbX2wkFkw2nQw+j
VRfg9Az+lIf8y/uMOEsoKZkz957+RwF6DDKbezNhwhN6ypYg5v61XP5XPF9/NDVzqxZf6cciD3lS
T/zX3YRGRxX6bLGcXVljBmUSXKAN26ZB31scLjRRjenjnfj3zzUKClLhjnTOBYenNDrjv5P/YuBa
I1R+4r1DBSSZaYC7WUDu2Zwugigqn81epRaqRmaroaYO2y8M38p9gBSd9oY/wYpv3B1X1sR7n1Bl
Q3Fo+Zc91CB6ghXxU1++GEEU2cI2S1jKLZI+uxa9/Ddnc6Piy8W4fvNQI9DhsJCd/ONjt90ql9oy
qh30jMvKlM5AJoL0eQrBu9cKdwz9SdFZthUYa5wcFM5T5cuyzCKnPHySSYL02vxPYDD5M17B7bJ1
dvd+HBnCsFLJK9RYCuZTOZjWnbkzayWzQpfnwLrMIAwnyspALZRauQGV+Saly852mFGD51+GbjMA
T8lVEoyJv9W5dPBx6iNiQRHlPnHiI2/tf3Wh8HfLGLRvMttgDarfYadXOXy7G79BxX/esyXGwyS7
Y7iEvRY+FoO/o5vLtLN3sIWC9gQ8GeEoGDFBTyJNsYnxDQpLMe8nMuO86OvdRuanVmXgcWKZyoA1
ouieSCnClCEVGFdhpQZfPgJF4djQrlBYsaPr2HGqn2jeHRd7+2n9ATufzS0imMBNpBc+zCjPAzSy
Df5dXHC5xYdTgN4CAqFysyPQZ2cI8ocfsA0b0+jminJbbc/24EUVOj3YgX6E2kCvnh9h79moJB2/
bBCIaJ7EKyznKF6pnW/+iweXQsu11By0KGLNLxRKXIhxdUdLgAy5yFgRYUuWRpqXR+rvYv2rCj7z
dFWS8BqNf4AcU8OMNFiOOqwV590clSTpJCHOnJ8944MgCG3ZuffazZZRyR8Z2ZTd2aMYLtCKSKgk
gARpc1M0nsXs7tFb5oRcQ0fmIDub4C0RNJELIXp3nJTe0ga6/B494jy+ppoClgacMOmc4PCCp5/2
mmCvnvxNmelP983wshMNunEfC3mHfCv5bwZEgF41FEeDkBmYxn3RpFsGRU5YNeAyrTk8KqdHu7dI
LcCfN4EE9MDD5yH9GgBUcO64JnF3nNpwp6tNx6X1O40PqewVn7RdBiYiZo8ks6OwXU8RHy63hbhJ
GbHc4KR6itWnSX+pCaqOslEA0d3+fPyD7HF/EtkUiUaVC1fQtzuNqQXC4YwG5egTlIjPUtYV+s5q
cAlfkt+bn+Nyswir50Jl0drja/qcQdxNiggk7fwiLQQQPgjd286NVCY0IfwG8KMK1DaqOLE/MvVT
eI/gF8aa4BS1WytXTUaQCgakfmCmusc6LeptKAeWI0tIV0A7fmXD/JIPS4Hu9vqIxxkSS1oP+i26
bKuraV8wdd8eBT5/kXJuhTI5HZReqsFAym0f1lUn1/lrTljAo+lGqNwZI0MtHOkVYevOp7GbyEgu
OsJ6t/bDoQ7cpq4oN8thrSXuC6CC+GCj8MvCBzDs1JIn065/lu6XrxEALT7HV22l9DYYX7W7NG6R
CXdte4lVaVqLT1Z/hd50tB1iAowBehxmNz/9EwIVh4YTfUjO39cQ/iHJElSMrNMJSAhXaR8xVZzg
pdRBU1DL4BqCdqB4DbBLDNszE7L9oMJOrxnBjRQ37CB51MWOEoTucxeigUA6DKftfreYxv6ZFasp
+hEuxra3azdlos/mWSo1Esjayw8Hb4zeC8ErtGkWtCsKPzy/Hc2MOJlgIwsj/HgiYolaufR1nYWy
TRGAGa4annW1hd0PfQCk+UjfRNhLbD715NK/PPDjL7h8cWfqhL0Ijd5Cz5r/QCefjMfyfioVPwwG
D6Giqd+jmLmCqCkLNaCmJn4GGFlfeOtkEglapFbOSeElwPYsWwcfcjfePFx3rGymxmhhyx5pa/RD
SbK9P18wpbiZbXO9PxAHTPzIXNj7NGtGjlkVtkVji5+nAfcKQeTNMRAY0CTpIC0Z8GOBah90h2JM
gkDiSZ+rdufZJ+rN51+aW5rqaFpL9FpcJ5q6iv+8zMvX1IXxb98IgNNvFzPKRVbNulW8zcLwuypv
kWc7QGEaGetfjiYiu+llwCkFuoa1HaTA9aApQxA1fTHx5m/vKLCpwyqF/LWKiczZh9cA6bif5aDd
/b55BjoRDr2mHESXDNeS2XeoPbob4AzsXDrbcQWe0lLUfAWZ+S+P+tFjXc1KsvQ8ttRsl0pEVAcf
5xCNNtNkwbzFWcvUdi4Z2mVAudENgWgjLD9WyYb04+XKvkmyiXMylygTyU+LO1GqwjBS2VjFYJv3
DsqY7UVYgguelsoZb74sVI62ssb95gk6TNnoorXQ2eJa7pwIrTX+dwNaFO1jW6lndkJMhD9M/jJB
wjI/EGy9nIt7rre419nAx84eOiHnp80ddM1JnnH7ZDNPqlSeWDJPuaLsCghdsoKF/AvPlB+R+Fkk
uEz91qCGvOw6JDrLD4yRNdcgU1s/RGAZA/QiQOlUUInWNG5YY6uZNzPDINuQOXIeN1IKO5+lHdMG
b/ofqLBW4tarx598N/wJX7BfqNBbZeDsC41oSshWELU6v3yTYtZx95Q1WpFS760e8qtnRTxNM7BX
0wyDgyg0iRrczwYiaMv4z1aEEsj3t4FzFn5pk58I1ZVmbEJfTRNhNinE+GfTAIYcDOeuRpUEmjln
+hjuDNVYAV37n7DXK+bwc+pSEjoMADDYycrBslnWTpELjcfMRu8N6xpDlr2Oyr0qpW7FZV4gmQDp
Acu5T6CXat6UmVbbmEHdnUypMoLsyIoWbc5eb8pHcdMRM1h+YtYq4EG673PnUm8QNm8+x14KD3pg
GV0Kyr1oPN0oofayTEcMFm/aLdYiyuFAj4VxpQa8GtvbWFBlMwbVcIKFgO8rOacaqJ9P7ZzZrn05
hPoW5Xqfi3iZaqVDCZ6/E0sv7wcXwE+nMItwztzZprLxWDCBRdN+T/A1+LlxO8nm0Gz0tNkO4Rjn
fdW8PrpfPtKpFSSIIPcxVr2thmmywRm3Vzd5m3vx/HIfQmGSbE99+LeViwQaa1ZPjZ1LI2DeItZN
fbjMxRLLEC05E48lpbjQ1yF8FucbAvmdw5FVgVkRUF7fEvcziCTK7xa6GOzdRPGsHui+/oPBeMLZ
uAhnzOP154dMpwZos4He150JSMILC8bNysg2Ohk5ht5cuIiub8eyJpgxD2xFCpkXSr4Hp+NPNsYW
DZnMogaIh/J+GbMg4f52LKoMCSGtW2pGMlcNlMDtI1Fm1dZmm0pYbRlt8qW7uahlPeuaizFW4ct4
7tDu5ztXCSmop3TyhxGADIWqDZSlIrJvHSEjuaVeRrzQEVupc2Vptv5MigNm426rUr3lQQ4RgE6J
ssr7eb7lpxZtybDcfxRUNV00WIMGvqvlLtM8b/7CcaV11HTd1mOjocHFouDDwWXyO6gJp8wtaYeJ
M1dDs2hoSXjlfWNLxlNKyDEJp5g2zGzbSDN9idlyMlqN5t+CakPtHu6cl1WZRhPbNClLnzG7bY0g
NPCN3L2kasZxnOrEWAST3D/2Icld14uep7lwctXI0dLx/voTEdOpdABuDBv0FpXMPDD0SlcR2Aij
/dC9g+krNhyLlrf8w4dZDMOLzXQ8pQFvCoLF+Y0TD1x7NFP8V1b8P6GhWj5rtank2FeK9FZbZgqX
FzoHFP2SB40BivcNO/EEXalrNFppE7mAFmoPs1r5QoN1aXDKvRMyMe6yJzQ6w5IATJo7HgEsQnJS
o7xQE5zV0W0j6UGsM5UAjNFDTXxAd6pGXO4H2mjc2TXCO5xvaZuWAjvh7P2UbEaqD/8aO9Gz/xgi
LRFLxRmwDpUyMi7VYAtbjiDqguV++H8xCvmOVfqIgKaUOyJeosahAUSG1FmL5KRnUjlMsMtpwSaF
3dcvvXeRF2KyOJqFQOXHn9yA+JcdJHOpkTkjiANu0PxstPoJ04rnd5ukEoNWokY+vF+AJ7a/YBRk
cvzaZJKNP/LcUgCNq7vE2Ej9gWHLZn9OC8Zuudp2z9ZJOblbJ2gldllDd+h065eOtdIME7hVoa45
lzQIr7xBPr/xVizkJOc+VLqdQYfPIkC63Mf57eS0wFHylvj1SnOIGzUkZHoX6u9dbOrnJ6GFp41/
j+362DvNwGl/ruLIPsFcH1tiXQ1gnkEoluDg+gVsC50mSbkLgn8DskBSvzXQjql1LTujS+aJ9zhO
fAjPm6vjeuf+OfB0npcbMiHHgLm6TTek0qxLXr1Dg7AHTrYJkxalWu+XNA9MaX6VNAnP6XfE3F0y
nOL6nG4+SLlIvqE7HBfZi1kgB0d8lBr2teQng+zNC8S2Q4cz2xFF08K9Xbb4dXG1RHeIMOTL/rsR
OnvSkaIkYZ8eJIejkwoE8bbpW0xpjJWtvDDVdytfuV05ylY+7rn2n0Q6bBpY8BPqSxNlf9NGNXOr
sEyWuG1H+XpPIcPXAjh28S7hjprI0G0UG0Smwt0R+HZcIERaFAYU7YAjLP7h/FGynlCA1JCjX/KC
rj6e01cfZldK8G3CHfxSkCq42G5N9YYwGoUosEFL7Ih5ixX+lJFY+THvNvcresUGwxdHZib58z7V
AuEwjiBsq8WJTFdLBPFhLDZUDIl7z3iZ1xbh+fCi9UiXAbHrTYcwrgDjDCEYj7ZAfWv/UDDCGXJ9
LePXTYDaapUej9G61/6vzZZoVnfFv8+mkzE1c2GhZVi0wabv9asoCnXOcSPIEnlASEykiyEyTwdq
T9pfBjQ+ADaNvUxix5bnyyBdQQKAQkgaIZU0CLKnwW1Ui7UdldHmHUs61tpnm7QPvLTDyN9KaOs8
vvQ3BzED+qfAedoqZfl+3aAh0itJEVs5/pioqTLKrqDT1oGBiK00BA2ChUzoG0kfNwli8SeJmLys
eOGlQ564bnjHzt17hooXAM1pkgRXm+VPfnmOtESb4EflKww51WeaBhNIPDeKE7vyvwYmpiPtJiJl
oHYMjLIEp3wIc2zPB4cMKxtT4vIodG+QOmtlZLgzOHOqfUQxbNElMcfrtJ3MXLe68kTHY3inyZsZ
bdhnCiFBN2Yx+arx2bHT7cAJz2eMbk/70yY3Lx9O+U1MPK4n8BZ7N5b5eUcfPwO7BbQJ64btV62E
0MDvogYWQrhaK0PzbB61YPCkERQDoSpH6OYFcXz783iGqnZu4TTyJ7KP1b4yjtj7jxfDb/cE6kvo
wa7Y+291AKmLqtmrNm+eI6zRZnHzC2vhQdBr8GWl0ety0pUFM19/VOTCgpx6GHGZH6HMjM4ia5AO
fFPx6ainA+xVcr5A/k7Poq02JgO/N7QhxGODpLH/wswxToRxizZldwz9+Cs5w4cK/qy5VbLYa53r
239Q+HnAs8Ff9Ip3TOjqT9IlCUJ3UNsNuqQJ7jpU+SlkghLEt4gK3jqodXWIurnONFA1jVtynuNO
hy9szbq1x83Baw14+MqRtXuqPGvsdC8pkQceP2FZWuRLIMzf+xM7PEZ0sSB7RruuLdg3IpM03w5D
6P2xsX6OokC4o0G8tnV+ydNjGa/Uhpn0zlj048ROqkkPGJl3bOmaxdeQvsCIYWfu9uebpVpkY6u9
pymL4hVDxhR12qC5zn7kIP0V1e0WntsZec97g98Vvjfv+5eJl3NI/B4yM5E/NbULW/TezCM94/XQ
d1CeIBdNz/CZTR7VoiUFBOWTmtKMOlf3F8BT2M75NFbYV9vMKhTZm0jE0t8kq27eJ4p/rKQGVyMr
VSLd3Z2YGc00sqyJNYogYh9jZJukRMAbjghKDe/7VZOKjzUZK6C42SLTRfgYmWQT52hbTX2VWmAo
zvYGLil7ZuzlNTz/d9otyzxfYviTs/qWQ02NFKGjausC/Pwspeg95yPM5//CzY39vsurki4O9PVH
GobJSIC1hENTDxACZQhR8lh67I3VYCHI2lUNlSJeUNTERsLt0FNmsClysbM/aegWoBOTXqf3O6/4
BEskiBChA6vMgRr0r607lSwW6jeGTz6BPvFpCIAo6z/n+HuORrhPw4UCpnndMtlQtgP8MrmOo3e1
g1Kvy8FF/9H3PPMNn8o3fm9eqPYAuKcybDq65zi3Sj67WqWxYVbBXrdNsC15VXbDG2i46oMG+OlS
9d95JYHGgnN8Dg4l9ferccokaLiTGhZU0VXbtsdrwudSDhv7SDqwLqdmJCzOSMcNmqO3I3uhzL5V
BcQKndBsy8bgl01K1V8KfG8/iiuDn24w5gvg275oVtK0MxY7uLND3GbvQIWEHs57G3fTIukTrpBO
pKRWCaDTRGTLwJde+bQq7YRHNwlOroLn3oudv3/Vbte+sms53lMFsm43pXlMqVR8aP5/VHXm7GRu
FqyXlZqbgg5OTgsxZTb+CU+Rn+DnG22Xff0lWsmDiq0socTt32ZdhH3k3FKymLKonCB8SDc3wGDE
8QhxuVv53z4Hjqu+4VGFshM1IvY52FwMQDpoedhtpMQcq2pK1oEXZaznhjfuLlcjmhhGVw+7tAuR
2ZAWB+UncJFTYmlrQXZXqVzIqn/vVMrTg1lFmB9tvgvZSkE/ZNfJ+pA6Kp4S6ijG98826cpi9FYt
v/+awMn/MTm0EiL+shx/iEw594F7QrwKQejgaQUMiLcIdT5cR78kNZqCY3E9lVTUD5YZbYCoCi69
1H/CiQLoOQgK33icDmvouSzdpoJxjZ9/5OJrBqayV90r6i8cSHzNxIlgbTf8vqjx1071mdCFXb6V
5GzWQmPgKor2v8mxJCJrDn/9wkI1IVlCB5k8UR/q2eKGrqVaFes+cjSLpDh2djHRiD1KEXNIpRuk
hlJDQrr1l0q/VFLF6BhopeRzguFDuUkn3fKF0R+J+Km0b0ZkgYv58S6EXBgLPpdgjFRQO+sQ/3+5
vTvA+X0Aml+3pvTmycPTSufkJOWtJWOJD8Mt9kvr5mJqfY0Dn6uYACbQRapmJ/go2AqssXSvW68O
rXHtG064rOaBtNBIzkzbvjj1aMyA8/OiXLH8UPum0LAzlXaJN1OxAOcuHwBBq0vFo4Z+peHFuf4M
4lSM3GukvbDObP8reSDh89bKeIg2ReTxlgYypsqC3+uUy84KuWPp16vrjjV3rAoaoHv1W+wGU3aY
Jw/saml1GPFdXg/jEqyloc/f3+YhVLGAogiLpJkDvi1F2ERY30E+9NdchvIVzRDV6TrgcWKgcQWE
Td+jsVKsH8ISvh1MnQ+ynd102m9v9cZxdshTv9d27n2iurxF/zPXkcLppcFkUzjK9d4S+EDsc63x
AIAtGV5cvfdFQSs6SB1iiuLMaGBO4/mw4jE/qFsOjDxZN3dGormXlw+XDXf5/cuSrmrFDwkVSD14
9LNEZbjc975FNK1YXLaDOhz00qhXeyvXv+jCsVvOPYi3/XuVXjq2ZTObmFR3BVOAX2MWTWDviXqB
7PM55/0gvObr5XIvwvadRULdnIsV4KbssRnxeFG1neoPSMCz73MrKf3KsVYmoGlwYAzdqRZrVdag
HLNCYqg2uyw+I9wb+N2x/9rnv08GuhOUnYsthTr2JOOd1NmSUXQx4j8MseED5M8TngW+3TjmUGJ5
GESktoudSkkkhXn5A0ByPWj4ITmON06vysiebNnGbue7g+DgD6YM7Ckci8F3Pfv8bDS2rCL/Lvla
wveYELp23elNUrHQG1roETNbiklAnJeNXPt5wT+cK+vCKik2jCwekq5BtKyNdqK8l/iEqq6bCp+G
AFErAW7GN59ChmVALnU+hVQEsSNK7GioNMNbATfimAixgYKZJU8Y4QPElA7XoQMNb9LVHR/Ml9Bw
fHLNpL/OS+3WJSeHcMTojaLWWvrUN+3Vhf3wsaUfeo37R0+9rJFf4k7wmX/x5Jo9SAOrI6oGsEU0
1vnDpOA628qnr8xtz4WR/pfphPovGzFCkAgSIdcpVwBo/JYomMfV6yTgJio3nwoGU5gyTkdMOjYz
LSKsxXdTjCx+gEO5NMI9CLk5/5yn3EKhY0eEP31pdJXUZ3iqZZm6tN8nwSKVZn73uCTlQcdj4XNW
d64PWq21nzDtT2BLgRzZcJuwRy4UJQRFnr5/1etYuZWq/zEtDZn9RqysQnSfuHwjP98Nf3+sBxex
lVy4/esrvIBjUknAoQOyFmc4reVV+hSRppyCJ9E8DwKgFjJjkSAoilmgjCknCYO/Vfgf9CGfjX/j
F59GhwiasOH+DgLlu1h6Khyw8cYiWLJ3NiJ3aDDs8MDWsjPIYgYNHWbmgMJK4nOh3syJrh5pmxai
kZYlpuL7tBMygCgkvQdv5R8vrI8bYpuwCn/INZzH7uhnnAeK1dqRTqNFgqmF02Q6hHfybrHS76hk
be7iP0gQ4c+orn/Ail9l3+cNAYJI1iAz2rwuyVN1hB9G/8jc0lRCKPYm3/xd+DuVD1YTU4tqxAnF
T2EybVcUC6D7UfBJzK93TpVm1rS+A3e2Mx50DPKbepSbg1qBjdO3E70YBBO2ilGhbFDMdh4Jdnd1
CQgydgt7fFdU6Ao/TXogx1faHcLVSBzzo2ilg71Vvvl22hp0s9HomXSYVhozElFRPc/MspVV68FF
ALQnbqBOJUIqaVjDehlAzUKLmqTQMIWrjocVL0VajCNtKHEfK8O7eAF2ui/7u27OJUKC+unmTJ8i
4RqHCQ/mJ3jrLYfsidNvmSTRyyAYe7HO3kktBdOwJEWfQMjrhqiUQWfapXMobIllcU0v35dSpAis
FLxAjPuaJqMHb01dzGo7F5inE+XEpQzlWx4pzi5D4KWTK2K4oGzFoX3SYxsTDxUBo91UjUwsUWAl
wpOV2wBfJi3EgWqDrZ6pW28zdTLe30sOBPbMzGwLcNCCNaaeCaIMpofpOeRg1/QnNpXUAaUSl+bJ
sUohq1n4QtL5UvkNERe3Hbh8BsKSr7jMwOJb6ldImSbpRzi8cM18fSNpbK7hvrgBIJrfg67Aqk56
PDnL9Di7JmpY4VNHdInmmf3J7Qh/AAHNrwiwxWUG72GR5Yzch0fCTFdeKisjvW0smEBtUg2jfHvX
GzEWomyYy5m2GbimlGjocj0lLEeq2P2fNpQ9rnUe5hq9RkqolJZdt+dmtsIibiObuZF+dbdvXtfM
UZOhsx0EvWZfWFhE0aCKWJcB9WDwc0VUavAX1I5BtQk3VKSmInz/F+liSgiML+xvkKusCOBukPWT
vrx+9YQ+MX7ubCskHzSC44ZdvXt0n9fccaHb/QC+MyHMzxpGiH6nKnHqSAF8ktSqhFN55XpfH0Ia
lohxvbtbLYhyEk7rCDGFb/x6/5mhmiE0+6m7y0DRe9XYrv5p1oKY65hYeDPXQ79EaaXCNYSaZwIO
93Y2rMnV8TmBgpZ+b2ek6nljxSEnQ34DnlHfeJQC4fO+aNVtGC2tTGK0tA8ATFRNL8XG1E2+4Y9d
zNuv4WUkTqVrhQ2w96w167BSK9U3OJiFqZ3+M6sKSsWffRSimDPz3MO2TZF6iT0G0ImpX+7/Wx0Y
B/lvEUkAKSNf8TJittuv1t4kZP5AYaqd2xmYAH+aUUxMFTfCF0R1rXrU7Yr8vG5wUq+osDTE4xmg
9A1NZAY1dY1kQgHCrZ8YBdEwQGMfCuLcWLLJFUMJO67tR2UVfVy4T4JjbrpyKFsBlXzvG0obhLoN
cgcOJJ5yz4O/QUb/aGXbX7kkgStfjPSNXH0uz+Gh/2hhH0As+QHdavZrRj30Ueqe7CUjwWGLJhS7
oLfZKzorwol03Ht5CkumUDDm17HLHoHmGJJ/rK7byh6dEgCQco9Rg5bRH6ZEwOk5Vbskk3UD4zTn
aWUS5cuK6xbrCnjVM0P3PLi6pmh+qUo2wZhZbgTF8QHYgNNAunLtvKvEojK8EU3u+qOIEYe37tZd
QS3Q5xOgBm4UiNMLudMPW5ks90FwKZ8bjV5Z6Ea1cjAZRzF2ivlgsb22lDgD4WP8IjyLGQMmc/KP
DyqdbNW6KPHeXS4DaoMFvcQd9AIOh58OAjI9XSFpM1ssV40Y8OITyyiBdFonSAakeKNVEP5Z4QsX
eXv1cUeSZT66CZYheG6nVoHxxnBOllDDwtPsF2o/aoqGLgjdk5DvFuWv/O+aDW6G8UO6LNWrwITV
06jH03+DlsA6PhoqHDPxaZrmEcsEi//XhhHD2XXdlDODijJpkddLDL6eKzsciXwo/Idx9MjaXnsM
8NfykNeQfOKKprj+k/XitaOjBZtzcD6KQVW0gpq1io47BCerB6zAv0LLeW1oCgIQaFQAusjQeTic
SmBAUbPB3oodZjZA1ONpI06usiqCyrXON272vqgtZCQLGbaunYdtCuYKmK7YxqBNOrj8kaSHvAlt
hiauDnMrCVzli7CClFnT5ahsE+B35EaTdw77v7RAH1PNVAVT0mpTCbZUL/X3Ag1DTpX/KZ8Xquhu
SBvaYboWAQkcuvEO5JPWVnjifk0/Lz9oiA2SjKYIbjBRk9JLCpfM7Dd46waHcw8s0WT7khVvUKWD
FxVEoVhmsZ3ZTnRY4Km5VpKT7Mr/ApYWWOCTWTnPjbEjPunZRlhe6HiedIwdT0Bti1r+YlxScl+j
AqQxrh2NsHCCh77IjXvJNw1GDaSOB7r3TYh46orCo6wS2YsaswqEgvtYDXIKXvJHh10ETyajx3TS
EQXjxAwrf7/ZSXGIewe2850o53g3lCR9cmUvU2IX7JmNCW4+vbZKxC8TVQyJfdaubMaPPsYwFoBX
w1IMFNE6u9gJZiyAdR9D10+4jcQHCChrINW66vJ70dAOXsJnVz3oxFww6XBVWndOJ0KCCBnXt3vq
++HFvqemS9EIEeLoUE/jSIgzXJ46Ojbn++pd2pABfwGrNQe2oGRdCv6fzY6u+i3Vvd2I/F8vHYsa
ebyH+oV19yLwpMth7oY02P2hW2f+M5bNa3+/lEuUXy/7DkCa9zH9MFeS7aJS/VjbtPNGv0wyHeXI
qLEIRH6qV4PWJndkzqajD5M7D3fwYEVIhXeOkeY+Ry9gfIhXft2jskCyo9QNZtoNZoJlDkpqV/Oj
JGShLlUXa0TZ0PbDHRxlK1datndaGte4/CW2UkyoJVFF1BttDNnAEsqt2/QQBn9VCtC/K++8KJHA
uR0YeqDlkxXwqXOy8j7nvDYW3aQmp2PujCVbSbRqU8L3GqcwDqUFs40jj35GCZFO6zgzOGcNbHmV
YS+EzlzluYejqpFeclhOwJrOdqMN4K9gkpGXgwQyoPp1mnoGE8wp0LmxMT0Kf12Gn+T9TMTaQqWX
e4cr85K/vtriAFylkBgrNj9zunxeL/WJ5iZ4B4B23OpngrYe0sZ6ukHZcHrXoy99cXxtnEG8+kCm
+iNvC31VszvSg4vLzStEB/l10YDGIH543qfeFEtLmeC+i7NahfHvSoIhyt22FIg+tb5gYbLSf6sl
KK/FzzMuIyBh9GqJRHKxJYkaehhwe0C5L7/bt+BquyR1fXNHQiAXk6S7sli2gGccL3eE6cSlp7fn
FzPwUgLPs24l7q9ta5TqhL3KKO395MwslUr6HmeiOdaMjp37Y+Vg8D03R6ZtOO2EaqylPAkXCU9u
l1gVk3wZoAekhZ9OjsUKT07hwoq86pK5K/UHsJF0MaIRvKuOpDN4Yxk3/YLOCwue1FCLF5fQeyJ4
hx24gm1Q2xdPyRr4bEzlKFbuN3C50zxxhsLGZ5QXPJsljxW5NfOVpE9aNZQ22F3CXHhAdYdtKACD
sdSKbZ5gKFOSq2Cvu3MCxqAJo6Li5KfqhO7eTn50jUAjr/Tr3pUcgxxu3MD4yfryiyZXKqQ03te0
w8w7LdvE20yw9CKdOvXebAk44EUiVjg4SD84Hi0AsAY3MGMQH79g/kKITvDf+iiw2sMUrob1Jc4G
VCdPlVOXoHreTQ7giI9hS1gnGEzJewFDJSfOz9PKVE3Uno01YmTZ/tbS3obXqZdE0f4GP+mklKl2
p9UEF/51HV7ugZFyOqorJm7njx1P1Dd4TxxaPSRKtIOVdJemz5a1RAGf3jUvwkpTW//SSODTjdr9
AtXjBQHsKtidSxgew7TTnt8RGIovkCr79F+LfdaYnzZbI88sczoYVB+MqeyHtUzwXcYzEPIjafVC
R2OQ+qPBTgm9dklp3ST+ZdLdn7dZEC051Xn10csfjXOWejncCbg5+YeCiSGzz6HLx94dGYtm8Tyk
f83GWsUzTsJ27SqlkMJud05tArlwQpdm15as94ncvoEo37PF47F7LrQLAXAySY1DzhFF/Sojy0eg
gIYv04E55Ibd/gFcXqj19J8f2OpHUrHybshcSpvSaWaenr/Yui6yHb3ClFhrcdHvAqjDc2JJLB1e
x6/Zw1ddSHlGAjR/t5mX2cgsqgCOSeGGlg0P5sXtHv+q5IzTNXgAl2OPIahrxpSkJoXToYqnHmHI
ajSXta2PEJVDsVOwFrl2yWBgkB9GDuy6pUqLdS+F0TPNe/uT0mWpkTJPJqQN+Y5GpMky2GslqA5c
niOowuh2NwV24epS2HscKduiY77qqO6CUcHJp8mOqejYfJ8z8mXQSiWBEf2pWg1tgUpGbP4C37ZD
dQSJqd/1NSK5ZOMMXj+lnOzQ+QWXzY32zEEl+JuB1ELXzcF/jOm6xxueHhIk13mesdhtiCmHwbl4
8GKMWxPr9Nj4Bfmgcrmd83fhWNJNSBszNfwe/ZHUTXRK+MCFwKVbAE6PojJiqw2XjGwiyIdZzJmr
pdBilTfLG0AtxgpftvCpIjaUDYXLv0Xi59rCOPOFZTRYqqJQgng4bwEvBboFHsISxKHm192GzJik
7EiXaYqBcfrGDTxWvU8fddG+XumHacHdSO2cZg8nM6P6n4lDJh95KcazTS49hqMbUlRFdORbhHfT
ZsEM6aMFbllaNJJye4SbeFM8fCiPaSnIkip6s/VmyZ1FWqYkIri78j5Yi07v4HutEcKfA+ublc2R
iqV3KLMD5+25X/PqEfl8YehOl3znEs7h6pMih8C9aIPNPLSNgRwP1eEg0uvWAyelrOJGBM/8bl0q
wv1rq3OPziJ08FonuEjex1Kkj62orPSOjuUPPPPzpWtV6JIVyGDZC/JspZMoerJveerXsf72aFVv
TSt51kt9rpgn7YijQ3E0PKK7RBDLvNo2LCVfqrFghDXZ7bCdXARqgzrcAvI7BV8Wi2doojKHUc7e
4/EAiE7fmKaI+ibIKl2/QDPmTh2gqxwSv89mUuCLBXMed0pxF9xlGAT6U2q9JwJPEFwOFK4yi9Xp
SyyitKb23IJu0JISrAHd10Ob8BAx2K6ZxNs8audWOnxq4FpeltSJ2yas/Hv7rAzm1HtGOqCq+p+8
yMe8sNQEf16+oJskdCABRQpBg59o4IaOzxg94gNV4Bx6vHHTxBmvBxF0oSW4etoPFWTJ+y6Fy2rG
FkTHii7hLMgDagatuJ2Xz3N2CmxYFfawXfj4SBxQFqu/kHC9l0cj0HV/pfDhvnddUlcEbmxWDpU9
mr95kaPFrefLyWnjdbJgVzb9GsblPx4jbbv00JDeul4tGx/83W/c0AZBMqtg813y6jifk8Q5JUSF
L7it19+K02/7+Ev1MfsjpXeE+wdo3p8g3XSkCAuYAEQg18Kt6QjBTri8YNLaHWFMEgXrZ8D3W0/G
iCNUOmLiZkUk/kQuUuHzS+TNxFgXboU457BS4E+RDrT9cJqmGKb0qmTfI+ANAGNvThzVu3H3xFWD
iwWM02OwdC5BBewuZvWiy6QgGDb9VqqeoA/V/qtZLGvVxOXTwxP4/wh+KhTbHXiXR5pvVeUp8nzD
bfYFyCZYIU1PrNrn57DfAJGLWJEAnbU/56bsf7mFNwotQrMCJArxvcz06QvdUeHntCoZEFsKt7QU
wryLho0hHCVW8xcPknUUy1HE4TZNLC7NubLmV4TGtXp8l/Dyo5RkvDiulO/AI5mkG3wdCNjtzPcW
bRSxQnt0NmVLy9mAQ8YyEr/+Q1ejj8bMKBfsA2rDxSDqiTRtem9C2niLlVpQr7ZY6V/J99L/IScw
er1t+XiIbLe6xtjjNCAiupcLSOGfJ4ahF28AXoABHCfxwXO/aJaAlkpf1qWYgBN+IQqX/lmjvdoB
OURRRuBYMTCVRnsMTy+CUZ+flhpGIbBctnbGrNZF9HIXpKq6GXWc+e0qPDhFLWSU5BiTSAkps94J
h+UGTehx9pjls47Toh5Bvnob/Gl215M6KH0iiOscmwfK0aVae+n3eW6N1Y1VXy0WufSxPIqwNXBT
IOkIw2VfGLxO2TSnLUs/0HfVf2NNRtp3zplqWxzyBPGUGZuoIdBSpYBdQB2A9Bv8omjK4qPuUHEr
7ctT/Ru/ZrTeiGONJjB5jWgAkEp68q0a77lMG4VQcOHJ5CFRHz0bxUtPpqX/HoVUhztFqiRWu3lf
JDeFdh74JptW1j8JLWyDbp2W31AqFRCQ7u0AgdTQ6T7S4XWJGWKgXuZHDNYavQDOZRsMwSH6u6CN
NRIa+hIxkSZg/az8GHzwInvdclYTH8fbwJKuLIl2q0sG+/uUGDRZZFY5Mm0Z4m/EXB2q9PWT5j6u
BcmQAc/o1ynxFb3yZ6LvPy77a7mdYlaFUVQic2Jzax/rkBb8g7AzKvcjPacldvNKGByQ5KFEe9b3
fYomQWGMhMgjf7r6CyI7GwVYoB8NWstOUZ5jxoOP2ooUAeDjiqvGmYMYmG1AQkMp3vH/JPknncw7
yDduZ5zuC946dqfivTNiMwuxYrOmS3QgSq5w+PDLvpbs+AOgtAShBpvkWKvpCN6qIfet6zSBlOYK
y295hHgZgIw46gBkLuvXIzL2CwEcTNcKvoc9vs84E8zTWLczwCXu+qdFYj2UAwZBNop+jnO1ZzAQ
p9gx4g5iG7iEb480nntMT52xDmwur6T1I/xTedC38kJ/xwojvC1RFZf731mZLwOmhSc2r9g1f1eR
tVbOLZxuN3YR7NgOFDxAVX9doKFMsS2C6VIoEJoTXlI4DeBFT0Xwc0etZ/0OpUzqamRs3zUe3bHS
3JcWTH87jDgX4/I7sV2nRwFqPIaU5+9X/Bk7uMPdMuQHkETLMT8W49VlBarkFW/JlByTl1FcQSnt
kwDJ9t+0/6io3XRR44MyIHwchvQnVX9A3PM9q7UDiz4pZxjVLcKqXIb39+gcxdEUFhKSzvraaIS4
qCcZbiVzjCS4Wgmaxm6jqgGmBdsSqBZYl4E07QJ5AzixxTBUqHO5Hgv0VIiCHJPkklWVc4qsl8vq
n8hZDgpIUgHAkDGFQVeGGzdGcQHBthnEx+HS/Tj8xsFxv9x879NP8fg7TjyD9uSfRFYWUNhXHntM
mAIvLcDJTzZD1/yFQEGb1s7VhQhclZa6K8iW2DerhrkaYuq3tSrFifwwxrwCiq7KSZOxuaD5ukn4
27Cqo1/06hMfKcfMg64l9MNrZTqXdZEAKTWf/9L4x9JCjqF5RGF5r7bAD6SL3W9q6O1XHx/q5axG
9LSb2+DB7B2m9b4GarymWlmDwGlPguzAz11cMz53gUMRLoU9Y4yShW+R6HGwxSbnw8jHa/SrO9dR
9rOsLtF/1Cw904PYh2sFoSNeqK2Ipok/m+LQTIq4anxe4pBZW1+IyqageB6zbVvyn8ia9ewJOdUE
zLmko23UTZT0cmhWL0lvJhV+qK/9Qmh1fEcMzjlmjGT2y/P7f07VVjWPrHmbIia/VM44DQrkUgwj
BmNlfRZYekOM66J+NnGlQGuGOOnylDi5yhrBf0NAoY9Gl6yUsBxp/zs34kZJ+PFhDNRGSeDR2sY7
Mx1SqrImLOxE22B5spqWVMxlDlXTuwumK6ZgsOJJB86DE1oJ4/VMUq1O6b6zQXJdyjAbQ2Be+zip
e4owaYFVKUCeo8KtI69pM6a5eVO32/ATu2EaSIUdyhQ4FvyIMO9CDsDzHfQ5rKwOXTHjdUCbY3YC
n6YC0cmElt2OnLjntxD9FiOY4vjkaHAb5lr+hY1g4C3rQYhuYJpEOfTjxxIdmRvKcBRXG8GqPGwf
ZlT73ukiXpYQ0qba6KDtqyURLAbvsF9uKQRkWhSWTSrN8d/7Ae5efmL/8ApOZeprtwnAs9A6e8UV
2C6ZyhHxo+ec+bVCLXD/c74D7LUkb3vGzjziTyf815vsLERoAX3HFl8Ywo9clI2xhBur7gkRMjlk
8cnQdSDVeph6L6u44uu1cN7WSJkKw8V9z+HfSKj7jUl7TYYkYqQI1wvB2Nuc8rC9Nu6/bM16hNi0
AQUgjBin/xqZSjGcZfT3kzJpxadjfuOKRNIH0QPtcf2uwcMPMPVVeSAQeXFIiySgf0uwUvosBKnx
Wk3GLEJfou3a98Wjola+Dc+OAxmgNuQPbKVppftmgdZGsMEyVOFqP3mhncGirf2dU+09Pbjjkg4R
vKv34QZprgP+9wetVnC0SQnM2nWXBbHzB4Ha6Ejqzua0KM9/uh3PrvkAH7y4GzWNPOEcZ32Xyiev
rFXtDln9y6R+lDdbO5uqeB02MhdnSO7b6AT6iaBgKF7NudL0rY+9ewQ3MCxZ/iaJH23ifToVSX83
IAnaWvqTMFWXCHzzdFrB8WLPRqGQT16B7nwFJBAfSqzmnTWY6x7aqT7+BXOuG8sDc/rf8/GIBXA8
B9M0ogH27qE50o1Plxov7YNtc5O2CJEeL3AAXd1G/h1qyOj+I9VJAH6Ftqe2XRMNVYYXMcKWgtd9
arJubE3+zhFFvlFoQ10MTNPy7B/yH9Kgl07WBZQZqiGyaQfNaK+5M5Bp8tXcHeAqYJYN4fZ48EIf
082DRTksjbHUOY437yDsULsa+EZEvq33Gzjt3BbdVhSeh9ZmpFtlkHJkHH1uOxuKCXReefHyfvMl
r+ZxB2JkbCo53UFkvklQXZQWp6BzIrh8Quxuxla4madRBy0dE8rXihPAWB0RKOFunLyNEefRlFXb
nRwuWG7gPXQUMgSN4daPD2pNTtfAIkf8hjX1tCWU/4EKkF4Ky22TgDC/kh0/QK6lBxXlcz7UJ/zA
0jIRF7FVy4BkBTD0Rgh3In0t55u5NJISl9YZf+xYuk/nQ96y2SDvAqWQBXIpdQZLB0vNcHkVvxCw
VqBX4y45VhHf0HaJASRZ7qzjKsnwM8GMozcSMfCDdlEBq4lCF/sxWbmxTzS6pOqlsW8unkbrhob4
Cl2N/SaHAoL8blEJwXgkTR96v/CL1JnwkaqfM9Ze4XTnM2aNxNil7qfpA/HkSnbG0hXmqhXXxm2t
bmUs7bN0oTfzsZk/HeGoGrSQKEqUFNEIYOaAOcoVCPvvXIU0MuPho1TimE3YuXDrHDmVEI4Dl38p
Tctj7P1HVcPyt/cLx+eOUB25NsWZclYVE1v0MiQIZW4/Nd4OiO4PDj+TXigUvFZ9HakQGYOn7jtn
ZG+HQDPDA3GTcNous2FDEZyscO4hQU/gWB3iJSZNZl67c2yWECwFiafTrhVznn/pbc8MRXU0RR+A
D0mJLmTJAC5KRIzkgBcHKnVK4PQ8lzKtN4MjcRVmqQ+mYA1MaACYqaxxLHgFCMkY6rYS/Zsx2vxw
pwH6iRO3GDmuz/tKd+4Qy2yt2QFnkuCvvNcIPPhve6HxJjVkSBUAffKobLW4BkE10lTizvwGf4Y7
BoOCgeNBS4NpXb4tKJPFg2C8zAaJY519XLDDq/P+g/rqqRwWI7Zy8Wk1e2MW4o2xaNlnanOTdKZS
97TRVW+KeevlMWD8s25yfDC/0Uf9kEQdQKZaGEOthM7nrm9CpcST4bx2e8fbiwgdhy8/b7UMK9gm
PMbAins++rnz9yIvKMq37SXgwIrkehufnE52y7OBy0ylLXKwb1U5lPt9kgUajWQhbCevhsAlGkx0
IgwU4rTGXwQm90k3XAZ4Qm1Vb0PBTjqWkJnZ4bY8GKHJUwL69Kf7EHYy6EZNzzi/SPx5drGI+WXU
Ow6g+Y9V6C7RBs5COuJH09XikLwTevRIETfuEwfZCw4UJdLVVlIF0jaOdpdzDsWA2XVjF64NtRGC
czBiE9qqgCo0SrvLYK13DsHJSGADJ7xJ+8Z1rOEAT6isHQi88xWOcEBRF8R9hbhQCSCcW1wbkTva
qlyoN/quwCJJHH/B1tyFTm8bXh+3rGtdkk5dlHndkSH2/XpwDUKWu1LMYRYfe6aYHiP/Mu+mw1Ob
yevgUx8VubZD9EkOesbQBsDgrisHMHya+Gn3o5Ft2GCHjvwbFBZQsVpIbZT5PcbzipW+lmkBpl5Q
i9ILweW2v3UiaztnL7XcZuRPFs6lIv3zQx5+5Gwji9+9Iwh5joTTtdlSuZ4MhWZlXLszUcqhvOA/
asi8veAIcsYc0NEBezXiX2ObzHuj/6cdYQxmH/MP8kz1UuKX6QwsJJxA2kLvf/K5ntK11jHhU0up
ICBBo0xmIr0Ez9U12XHLFcqKjs+eqS0cIFPIHRnsQk3zVLwh9BeQCgyI5MCBh+wMcWuQhgrfbHE+
3hJNTi/iT4wZAGR1Il8wizUroBSKOEs2L+tSKyoGH7uQ0NA2HA/1jamgmcXC5YOmm3Rm8YgVsRGt
NSk5pxzFNpe8CQLLF3EDZt+i8Slmnau2hi6p/t7OMGyVrPAbwY1RUnO7kmMrZ8ILOydb7YLjDogz
x6WUpIUnjqauD+wRvOEKKHTHYZ33WNzFehZFkYAvyx1MFlPYJkZtc8Xs2NObE8Oog5s4QqKnIoVp
pHM3cgGaJirfKM04IOfHR0ME4KtyomHgGgNahhzYqJjLFud5H1Aui+4fTxoxw66yRIhawZWT5tL+
IfrLEJe3+8AyP59wiYBw8I4Svr9xPkPtAo69VRR9niBMh7Ja6k4oawy0E6/au1/woptirgtZzqKb
yIOsNGpgvqTex4Z9irwXj/Q+5YbPmxNECj9dKZLXuUckDIMB8P1DSUSth/8ZrkDrVpNO7NRXgxaa
FU/8mYR1bLzezrQrNSJ4y094GbERri0evloj42Uhk0EPQx+Jg2GHSSwuybfHknoYs8g+fFjFtBHQ
3Oo3plMwZRQNFNqKugF1kl8jpjQQXtuAn2tZDPhc/9EG7gYa53+HE2ojkvluHtQTXTQC91XJHYz1
J/NKkiwnanVDeVNm68RvobDA5pAezSwe1GiaTvxKX0VrgyYXZruAV71h9CkVoASKeat4FLgwMqjE
nE3zoTc+mZd56gGJaRZqu+bq2cjEnaGP4JnewSFiWcf/0LcYinji5NWTxgwq8H8agepYvVaSUDc6
2Vu/dTbyS/6Ft/PsoZIxP6Z8PMb/EHT3pxsbEkO19u6KJf9LX5ma0qQ+2Gh6ovWYCDiHYCuKrC2Q
336i68xdBExHzGb+xDAGeeSfbz+olY+LCUvkD1KTAWe74sVR/cxp2jn/EB5lT2AvFdcbXmZHPN1s
o+S7RJ4k5pP7myX6jVP9XHV7pFpk33BzyQDz0OHC+DzcWxE3PUDYYwzwApd8p9cFY+msl2wNVf3+
GaIFeYKIOdE6ltUAGXzK1qJjPSBi1A8yy7dovF5HoaKB36xBdAYo4W7fkcm0m6jT+LL4nKs4BBWX
6yqi3FGgII5eGpLL2MxiVcl6SDZJUzhs3RZ8QW3S65S6kkviO5Rb8Ch8kuTHNe5cGElex3rGOUfJ
6NOwLfNG7F/JMpO7JizzT74epTCMsPZ6O5msumylNqOEFwo/cCgoqj5osVqtzicQNwJuvsHXasbc
83gTCYqdlM4sIxb5QF0hY8NE58xrFuoGABWU9hqEUTNRg60lByS2ILaitzf/cUhwnFJANQdwKinb
c2eaJfS716+vqIJvk3ECvzEiqqZUFn+fl5r+CwAxzmfSd+2PJre0hlVWhZlnHRPiGMTrOLn22Njp
z8kxHqh8cZIJR8AA5GKYm3ifXx0s/3vfvdoEfJmHicIqEvuUEUkXZXpPYmiXdJFBbjRTqGB9yPGR
cBQLSlTBZBMlP13yIu1Vm47367SE1i283HS68kS+H5H2sQpd8wwPyWY6WnE4AuofnBu3sYSBdKvI
ThhedTYJ0uPe/3/AIEMKxQOvEAiWcMMXU4DN0Li/mXJaUFaFVgdAZBiFgGbm5AcFv0WPV7HpOfW0
F1J1iOt4SE11LvVfs3Wlv/CsU6qFB6l8TAPwY9cio+kdjvvc/DxVekpzpAX18TBr1nrLKZYxW1dw
CjYXTrZS5kHd2OPW3LlCIEFOElZlkb3nTgNvv3MOm5qT5y/VfF2gz2TyRlTxLvMZnSBkK4nvhils
D02yp6Sfn34mXN27y+4U6TeyKe8ju6JW/trqIh5FLZFie7Pt6Eergr4OAV7WyWoUdCupczLdxyLq
OErltwvTpFjK3d9YOLqRhuH19iFjMU+O+ADAm0N5XwzmLpRa4TLQt5Dd8DkWIwC+g9E6flt5sds1
0/Eq7G9hDZbOx0u+MepnWqkKpgKp/l6URyafOMhLhYqrv7MUHTwI3b8qz+j95gReL6S9WL5eCPPE
EJPVuUDCQ3x+51FZGueG82ra6TwqhTRQyzzEGJYbfu5CLGBL98O4HtOO3H7ijQzD784sMRRyteXn
yyY80xQVwJC4GwSU4D9FrRiU9jFy6qbK9rC0OhDOgXbD09Xdc0+OIyUQPqpW5jAfVT+zUWZvJjPr
nvnPEo7Gse2G5taFQFBOoJCDCv5sBm76TZFhhTFlZCsFtpVqQqHAgXR+mRd8ykZija5S0Dv3OOEn
6orxy027GUJZUSuYbBEn1T2UxwfSNtzCmV77NjwBQJ8vHVnvzSf8Qu4oBqLOdsIN5rt04kpGzKPn
a0EIrrKVvvS3q3AKY4l2hfxzOZ8M7rh17Pi0ENQe6vcYezK7bpZmqE9xaQ41OxvVumSiVMCnPewK
hoh0T23VxP3Z06/f5fKDwY2Is9loaru61+h9MF6HHt4Q3rSneJNCFEc10lb4QISCJQxmShiO3Efn
BtrDh3qD0P3uMdCoL2JHpWihxtixHQAEosFxoHpdD7CtvUji6tNiSodM8+xDFPsRlJlmJgpJ181x
ypLC4jSHtAAkafxnbwctSCT1gc0qNXxAuLQ73Seb2b0polW2sYMtMV8+PBf4Ec2Bn4k0Lz7J7AEz
bUNHy0ffwM78o6iRkeCyE+M/vtxdRDlJ31uq9gi3x9sdrmllqVCtdWgW6nftFAa/BpR7vxRKTlId
z3RPBPlW36rxp5IDdtPP6wKac7Nu0JUk6IgSFiGD/IHvgizZ4v1Cpn1H8uT7/wPe7Pfwxag2LGbb
yGNCu9+oGlYFkZzCmSH6DHwq5tyQYohoMeBg6+oSEJYWhtfuqu++phwGhnbgo2nsCPktkrsNC4fJ
nqk32A4Hf4JgdtZLTqVd2SrWPziHp7//O6czpJDUXQq974x/FBwymmX8BPQsXGmH2Vr8WoTCNiMm
b4hZXK4MJatQu7EQOjvzpcdnTPFSEngorMtNKxUNJ0T1tJRmuoH0GYSAL0nk9jFfNNYCdULFwfId
F4jpUzFOwWdSVF053ohOYJSP37Ju1OysOQoZFnT/D+ZQfUvLMDwCzEC26a3u54HNlT+K5s6T+Laf
mChNJs/uAkU/x3HSwqVOenFxI2OEDbZOivDtBgG0cd9UDoHYXuSWKUegbM3/PkV48O3K4y1WnqiQ
5s6x4R1j3YOLhMt4OJdxAfdLqKxKvFWjLAMerQL+7Fdjuuy+uGn0cy6F3XY5Y5gWyEAjBB7M1T5X
V+TuF+hPDCgC3so5M24/HpgwE3j4MAJar8bt3EU72TrQ8HOfFYHO3eRmWHuYgtPgM8U2erN+JoAd
cyMAC/fwKjCXI1fpiLewICtSv+4BflkY8KuLpmdA5jVrcWth8cBfzX/YiElPsTahDvjbrGm+jtGb
gHGVY5lia+aVjWg9fvJwq6pCIARvGCBgiPOdDK/y5wiuKkbix7a9BxHVYZuufUdUI36imX/ayGrB
4xzr17NTfcf+8e6fu4aKQgRPheKesHkk9N9O7P3RTdpGj3VRFCf0X6Ro5DhE5aEWmPFeCaT7D2qj
iiHZ6y9al4lijmjdlH15TVLtfEnOCMXujXX/GezxOQcvIijsxKYiNpFbiln8N+GMxx58BscbIikJ
cqMkjOYFZcoBSVv8MBoYNzb244mcF92RFxB664y7xEXZl+2vhRD/BK5xkaSm6i2zwVTckJBcARJQ
cdt11FJL79qAC+UYlxMfGGcqT/AqU/gjr+VfcENjvZJZ0NP4Z+ro7udy948SxkxS4mmISBXRUqep
dWG1Q3FUzIEebeD1sn4ylPkNggLieLWCUwSTgCYn3gRgk+MJB6INQdUWwqf3sJx99zOEsEBr5mZo
WSajDD310ZT3dN6cu6mZiR6BVo2/Ny+UdGtyecF44SWWv7V4C8VDYq5eiF5yBlKDEyT3tpbLBAM1
25RDKWUS5HdRgeN9SpZbXhFXLqldOSOB7yGYd5wlBuSZYRh6g3x9Fy7UXMIaNUViSMIt1410nfG3
r+HhR12kPDiFMBr/Z0AGjl90aye7Tvcm69k2auCXkJIU8osJAofjcc0vXdGOcIi6tArB6ZIhAczk
DPTbNkkWXrb3BVuGAFEOOxiDs4NNcemyKRn0aO9AT+AQ5yuSFYoz1/GFTtZbtx2k6vvRLDP+XIMN
KaO+HFrv4vYqAg8+B4wkfbvUtnWPCQUaAuIYl10Ns8EXI4xSEVbLc3v6XlgBFkIaUW+lWObQRAvl
xgYv3GfLp1jNEeS4RiL3qXywZEu1jCjkijY3T65aZQJFGyGxJSMnG0IR/qWRH7UFK2Ftac19xj2l
DNi3XF/VmuKuswXIMYtm1WHtD6UrLZ/5s+bDn9eVSKa26OUuoz9qZicChKMlMyPWW0+Mbq+kH6Cc
fG77Sr9f8MypsjjhZfA1gm13R4aD0G+o42UDuugFyqXqa/720cWsgYI8SWj3AJLttmty3qDyrZ8i
9A5wexR3xuQgC5O5jZbIRzTL7SjMS6S+crGHaCmZVetkxDf+I7wGcsez3j9/NoF0tFY94bXGJyx6
eBrgOUD0/3WJ90wPblKBusycyAFi1lfCcDdOBFiqzM4sjYn5sEExa62FwWDUMGjiXBlLJw8dp+wi
m8Y+huUyhapscLk6ASU5ayIT8qnHdqbaJCNbEWq1RMmnJSCc4nmfX+CVc7eGTVZ+Mfi+OKJ3BZYs
1b9faYksGsaPz+HMi5XDqRrNb4SYPfprBG4t4SvhxgVuYs+vu1rkdN+AxlI3h253SdbyfGsc5VTe
c1aM9KNha9JyE7oUyYKdpghhIvo0+V7WIO/bkgg+W/2DyXY6h8/mHAKGTJb10k1hyJ+uNGalvbGw
zYfDyFYkVL5IPfd14rEb59UGAXl4Nu2TDldLlgomCVzSo0o24Eyy9Xd3ALyo4No3tOtgyL+IHkPV
XAMeloR5oRw+aeaI75Wc/VSK+DxfR506rdmCBt1ycmTsN18sPE9WXN1crnYJ79gNGt2bR5FUj2Ds
pdyeasT1kav9utl5HhVtbo4EZDEVVkHUU36lxNwM0PtqBTg++GxPrdbNZ773oB5031l89DyYyLj/
YBuqW3YoVMZKYEWIZTQhir0LBtnqrEpebvEbihM+vC9Mti9Jp/D0wQnsU7uJ2XE7/jYg6gyqBZBD
LEP070OqKXDSoMukMiaFjtXM4czXNHkMLYHr/Qdpvlmyh7Eq/kqmvQMm5ETfcKQn2UoHmLbEeejV
W41pe4/4o5BD6wfUXxq6odsZKM0gptCLot4Gwz8uMKmSMVmVUyYPLJ8liJEd06WkB3AQPq77mBcx
lpGkGg0bu4tXcIyaXQbPVewEMI7g0Ezhbfajwmx4VyVScISK6X/e+3tp6Y+zNKHmKUNIbFO27VFT
DHOn2BhdYYZf4YRx0S/W8RDs4oUK9CgDMrpDL9w5fKp1t8F/RBKT6efi6YubcG1l9YM7AX6gnQFl
Vg7szF7p10zeeJSObN4PPL1LvELUEouraVkbetT3g6bzNo+S0P6BbOK9vKj4oiZOHZPlyoG5UODC
rTUPaRoKBpMcKw6FhJU474gNShuSmGKiOmtachEDxWjjwfjJX2jxnGj/LewBGKug8gGo9xx3Mbdb
hqmsg3eJsBVq+9G2TYacq6EvkfOh6EnoS2sj9rzIe50Uv/Ms2R0abg8Yox6MYgpqDeW7r5c04v5x
6GEkKWpHf4ZTCzx29ZOkI3jn3X/pJloooV2tpb5wUO9lsxFfb7v6Us/kZLHZcOCOessMHFDkStp0
iKuliWzHmDJg4760YPh2kUcHw+6/cWPpBj5MjwfOzTJ2PuzSySrR/hJNYHpz3CaKhzf+RovALZFP
uJB7OH2sXaULbyR634sTdSueUqn4ZNIH2z19qsw9XLtUjhiu/EKsCXnZFyn3uH8E9e/U1nkSuKgy
eX2ktvLwU8Nwz4KGSdyRbs6LH/SYMQ19f+YQG3SlB9W8VwuxCs8aHoMrD0aF53Q3z91Fe37Ey0MW
XL6vcqyXkPc7FJgGH+2c47XlMrB3HjYH8T95gRFnphcl5mVAHysWPRD8cVEDrIWILA+2LYfRKO2t
ZR0TRqp3r/DUgqJmjxYgBJTD+rBpAWRpJprZ0RpBF4qCB5E5ngJcnySPced5RMxHBnffZCNxrpuC
m5tTIT3raD0xFaSpE/dAR2bVN2W8ifaspxwunU2T/w7VDEQ0jd53Ep/T3zMsvIT4K5W4PXecQ1b6
rbf9SZy5Jru7gcyGyCUTEk8qtK95BAumXBxrl5CpZbKXfCTmyWeGslqfRfjV0FnbBNf69HUpta8Z
ZTOClGceIISjjPSj+erBFTThYPVukmBVJnl4PgGPuCmoBtBTWzHzci7rwtkGVksvM8jSnBmeYqS/
OueSyGkApa+rk/8b4u7rqcQ14yFQGyuwsF/1V4YFxZtj/lCzE3uqUoJ68GLAEpFeToUqqhrzLoeG
6lb0XHqF+3r+JRqQpsmwn4srXGenFczxq3EYwrOjJCq7zEqgIPDwhIEu0vdRLoMubMIzQVHghtJh
KOyy8jkZGTvSkBP70lHcnm7oioZayT8lJeJ4IcoO10RxCbYPddPQCNfu4X7JMjMaozVoiMN8+Ib8
MoKJNbU9eA01sn/Be1ZF3DJAeVHrv31sT7Au2O1n3zgJ70uqDpR10QxaxERpUcpRyycCvb9PYW0Q
vQFWOF2UWYwlBvkIRnZE2UPtPW+HZOzfV16RxGoWnuE7GSciXuc6tBqqM0U+oedbYCy546J0at4v
5r8E5KGqYnRjx4Zl9elf+QXp3XwcCNkztRpYYq4kmQ0VACjWvcRSw0UMF25DEeuK7T6zLLNtKlZp
+d656OF/poLhCTN0bRaHNFMZv91kox7wcCNAfhlQLFT+tugikh9aVLYBtxvRyV+E/lh64olEq8Lm
cgHWQAFX0yHJwlMUjMYLmIa778QYZWIgGZ8+wpa0jjkr3LZt+35A32BKZZ/y/QL9KlEZK/GrBPf4
EO+seFidi49pQ14e+XTAsFZs8TwWPxYipwS1vF0KNZxl45krgP6mjeAWD7QGNb0rY06rn9LkruQ0
/kYIrteAZ8xXUCkCNJr2DDFElJF/duUqxBMApKlgiOsa/8TBJoGIZBuLJHgCW6odv/0AGhnKw+xK
UUFm4CyqwCZFz6cmIbhdpFBd1e0lhiCVIDvzCYwLMcU6q6GUbNx/NiiKnUlkx7zG0xJCA+ysIu5W
H2z53kTb9SSnLjOl7sDPcmimQIakRGguUw7iJ8hDkTOzd16j9gvCcHUaWUn1JvO763NNpijnSMqi
K738wlkxRa6TGCkMeeZ9WIxqubMyk9HC6G06WBs1U5N86Xg6rV0Qwo6yTaXTj9XOekXE4faSCsmz
PW0UobWJOMECpm02ZLVOS54+VuLfdRwMl4xoPXcv/WVfU0iwuFsPAbT5ZnrAf0fpLStSvD4uggHm
3W6Yf4YW7aVaWNHK6bGJGBd3EPUqI3BcFEcE3sEfdcsn+GnLH/lSVE8b+VM2OSVA4cpO+zpZeYS1
GgS94h5otHKZhojxvsSbMXeRgoO8eBbo3C7nGnqoEk4a3rHItDRc1fmbPwHnZzEBzeHtNQcfnB/v
5drq3fai0WPgKdichJD15qjtiBrSmqpMliFzT+5vyAjS/tyQGZGO5eIO5zp/Oq0AMisM2eMB328H
5tbTcVHCVWR1o17r869tTcY+ERfAl1TGGRjwfKdX4AohENurEL+x8cDpWUtYBVdqlD5fOEjBtY5w
EX4a7soIJYA5pgToSNp1rV1i87p15OpXYSakZK7y/WdKVaOkfBIj/kTOYWbXjnnkryHwQDyHFqya
9ht1kRAdTjo3a35OJ80Gmd0Mq4ghCtaD0SwOBJN0A3aHfhlDsMLGLC+6b9B/LO1WGgdiYprLKEaD
OXmXB4rTopHzvasVt6rWKyLwezjm4lPWfTLNuLbnz5SAdvejB1znVhecmCkPPt61LyNXzI1VQjI1
CsuIVQIS6B//sDhPgf9n2NudcWcbke/XQEeG4gQltmMMNUYMuUYW2LfIQnIoKQ4PUZr91uzU7giF
Wv3i/bUTh0XGXDmM6UQdwlPy79PZKh+Iq/oNmra0p5ioRHRjHTeuYeGYZHOtHJNsTTBrPaKS7b+h
Z7nDpJdXeoxXFS4FpVKwUCK3bHIO7nMJLJSUz7ROT0TW2/j0woodLBMqGdkYl38pbLJw1MdsfSlR
vYyINm1FNW7YGW0r8w4OLGDypgBK5+SVijExe/EIqDBidoqADiamUj8KQT7Fc1wUBRdInL2k+5e4
VMO5h/6/u7jye/2Nlf8OCyvi9xYGkIfJNn+WuZruVajuAA/iwX6P/bzLX2ht0t/ortM+oxXZBYl0
3jchKcMmt/bZUpW22fzywyx2n/2S673VMtZuqL4PQZnx4fSN/tvb4cvUw7Bq64qNolNnkpgwnlPQ
cLbaSJ0IDWuFOLIH6rlaWmLmCh6LAEpAuqgPI1ctRrkn3ovQJ1RXNJru+61TsNTbyemMlcjAQVcf
w+ybH+NdFeT8HoVv47d3u0YkRNMvV9KS3hshZ88YLYCXQJ26OHy3R3y2L8UJujtOFB/KvKsDnoOl
9V0ZahuY1phnqhXptRdcb659qGQVngrm6LNzZlcPDowi4rhVtL2lzTGqEErPQyb8d4E8Bd8dd0Ei
scvX7eDy9bSbkMmLa51FiL8lICXX9/HA52d23cBXnrdKnFyhX0P0cvZ5Fmggm1RFg6uWIpM7Sm5Z
yX6BD8HxtDWNOTaybfpUaxwUeONmxMoZfd1ZPyhRFdsMobS3kYz1DmSbzB3DzPteDTLM3QV89yTy
skPqGq9ILLcskI4Yb5c90rjjmXOpPiZY9sj+v1FEUq4BDEet3fDwmsycILMfPk2PGE0fgear5jqn
azHoqnzAL9zcjwp4rJ8CsFA/3zspAKtf1UT9l6BmBDScCuGhq+XTUBsnMSi+EHaIjwrspy6Rmz3u
2JKO0gaxIgzBzuwHwif+9anP+p9uy/mzDsM2AmhaYdNJAxZEZwyGwxHked1q/J36DyGm6+0kua07
fxRFek9qyl6yukm3cxWq7jLB71rAPUJLwWqL1zPdBwFLDyQIEkSDTLb0FJHVhKZj54XzscHhtyiR
88ZyX5R1pAGgiXEy7E/6tQvSHLTVDYEatdRLVw2+olmDIrTSXlI4zUM9SrAJwq1bBS5RNl0rwgcC
DWrEqSDJ9E8e3TqKoWKAa/5ua+YTIGEDqleCjAOped7Ncr+zcMeTKuG0HNtZHsGMtTA220dYS2iU
65mahj+SVvt+Xtqi1VoAhn8n17PEgpcU7aZEzkVpSQfR5AhiOwEL9ysHmO+YyA4K3o+bVLAtbdb7
Yv7EFSnF2Mq8AZUzQ3qbnjtFgiwGf4A+NWHELar53MVE76Kp1tJEejjLufpX0/SmoQ7zuO3h23bi
hgzhikOoc6OkCtoi48k6JQixHiDo/FI+09RG9PUFMdoPvHf4KlA8en8zU/jnfNaqTmHW14gBb1Yk
7bUqOmw5vQyb2SDpCsNpB/elzSAgK4d5bDxe+CZilDHF9wM7j9RCCMkGT1RcXlX+XAooOD+sai2m
A4i+/sv9imLih5jW8WEYmyvIWRHBYEVdl1aV/RF5DyLf2LRMJwC8V302e66H6PDQgdNfuvaQmtG1
b99Wsofhi5j8Pd83EjfgrtRWj5OFsBGWUQFvemx3f6aNeeqg5vdZkzz58/HBtjw0f/BBgvXGwpQu
lwGGaxNU3mssH+qKJxq3rD03igA5EIRdNQjWgUHSwOiaAmg4Ep52ialF9bu/+j3LAsSF5wQsBQIS
GTKzca976B8mh3Cmqbz5mPL/WStmL93QToO9mCK70RunedjdTyJ8VMP/FP34MnnB/2Gy3OyQIm4j
por/HirfORS6iF6+5hyydZVO0KYYHL0p3p0SxreXJDTP6TSSzSQC1mm4kcvQyNfgKLPNhbS4N9lZ
gIVv0CTprcZX2lHMnedO0yNMRoVLiPVkCj2g1RwAJ/EodwFYKXId7zFcWFGR3g+nV8iwg0ECt3+i
fobkc4+c2Z6AmepGCa22J4VZLJanzHV58+vOkXTBOpmNtopbA0ORYYcS1tn2BDFdvzcy4nfKy8mw
BQjlqnDQqh8TNtP7250kT3D7LmyR4+562xi9PSONCpDyfaxHpzuRafbSltU7lnlgmlf0GnOCGJ1Q
RudHIgc7UlQXjrtQTBMEoXZTmBp2he1UnuiJgeCicsa9uU1PRcZQW5s8BpKdnSTOuXJASIFGUy4u
7glJFTZMc9D2ikAU8bgDvcowQaDiC6rDtopn6C8i1/UZ/9YAKBYaOBkY0+yDIhZEt0nGVZdEJpae
pkE7mo3iSVOWFMUlgZdkyVLBXjruGfxr3Gg5nzQenWjKGVeYMDbCfxvj6P6hyxKeQr1F4cu2/Umc
KaaPxYfty+oEMmIExNf0gCaKyRE5x8YeVhxA8YqL4797weJvyRXRUHL3DvY6aMOy6Q8T/E7Y6bHH
8/EvnqLMFCF/Xw3Bw+RMML9aNBu8PCdtXpPLU8eRwyUeqL6+QB9ne+QVTv84jMB4nFAr+AyTo6dM
Pd/7Wn6KxqGbioG32gs1VmPsaPeLRgkaMWSjCp9aOp//pLy6afg8wsF+J6DLIw84TISiEimKi1g5
YbjFSZRHbsaiYNLbzMkIG/8y7aijf2rpNNlxXSxn4GluBRWYLCKrjppokD1fqBgYsq++TNxnqEHw
AbbA9p1wFTAxXIIWaSTNMY8ckbbB3WFro2RYZO4RPkIMWClQnaaRKKXnONe0deAnQMML4MunKk2n
ofe8ANfK1BvIK0LIX10QXnu4H7CJQKQvqq0nhVT60INZzBaGiJiPHq/TFUb9tYQBBYSxkC8HNe7o
unvMGusRB1SVuweN3uSGE+Es3FhKW6KA7QRgP334o83+GOUvPWf7MNsDJmQngKv1Th6S0f0ly/ZL
UnHURWGMOT5L91XNjxYrfJoyBApJMVJlOTWsROUeh5ENbVMKT3GMPl0TkvyStAj9RlDD/rL9KQ/u
Rn+Lu9UpvBPLv0bLGzc1rKjGUYEt0jrSrIJaeDYTedqocGGsXcD5iT+AZg1pv81lTYnFuGM2vT00
TCoJ4CGI8bGirdBMXsBT4MuL8chxtSKESJr68X8ujJq47HybrXSibs5/jwLIjvSPEG4Iaa9kjCuk
ZJcq5rQP3scUNSXSZvHfwNpkIYLvhyF/oU1toF2D19SBBFwgzoivw/CLA0opuhMpQXjntCrf47fW
+yI/l7PQ7lKg5uNj8eAoNWyxs4qVYT2PiCPslgzF60f16KEUbUw0+I30HtmH9i2yrGvON5A7I8cS
WLhQSCd2aPCRI5iROBLuy+73/Yb2sDhGjfd2nPAPm9vN241iggGQSc5KJe9KFL/wkOutxVXoYFOu
kgSuLb0feVBadQ8TZ7RTuEkeYnoUSCwgcfvrUMylVDLqQaTMuLi0wyYVP2quxVAXPerBdHz0krqY
C2jjJZ/h9+pW0m9cijG7/NyVAInveJfaf8gaQxQoia906i4FTK58mG/JOHXkmVNNXbYWYl7wgj9x
GFqbQC8NBgGuBxhP62cy+md+HYe2FOrojuS+EwL0wgRvJm0TSo7BtaXbVPOzycc/9KatOAgvMeWk
OW0fVCgbmRoKfZLFnbpOY/Fa9PMOc/xH/9oSIBibMvTASweaCevhMjZ1EdHCIBrUvbqXD8NoMIDo
qWVLxAXg2mmuWNCc31aYanPtN1SFVdnsX+0YFnTkzsX+Ur67rw/BjOaFDA7enVvmxWjfOjr+2S5c
fTxPFRaxLPin3ZHuWJs1f8X9VZX3501GyAksKjQ8lXpelihuqSMqF+q9NpOGXWzikjjzOK7o41g0
MYRLZWm5mcflgAdQaFMAgTV7rd0tEcGxy5ra3Z5cArEwtCOjUX+6HIGH/7a+r+ey7UMhd2NZT9F1
J6/+/ovgA8uRXpaVdBj5YiaBezWMSe7fqQ+kt4f2go+Y1Rsg1fN6ytcqGqKlzRJixIvH/Ih/Ux42
iGfOaEWkYwX+26sp3f28KAwiy9DgO6Hz01sHTpj01/rVFEZmzoFDsiB0znpAmo0TgGUmvRjQiSp7
s8PuuOChfvVxntYYZtlpTLPf35+wv1ClQJAXhv+ekOyHkgd3K4dHE5X2Qxz4V1hg+MrXgfoZ/0Z7
aZmKyqRXd5lloGF832Xd0HZSKlEPYzxG4ieynO1cbyJqUkxAwkQF83Rba5ZFBc7nJl3fq9llrvfQ
zZKdzlUT3Fbq9g/4FrICgZzP4wq1DcZ7jdFjtYpIhAJ6d/TAvbLtjuEoP4O/jL60SmZlanUwFMsJ
vkRvtw3Ggi0AYAjMMBoQ6FtBakVElmvQnGz+WmhEsWRPvtMYhVkbFhHY2CJBpPoZZNAI1FVH5J8U
f1t9eZ6ashSDmBaUgMEWy93o7h5Rg2z4S8oUYsnQpiiXRxN2k4gAmwVvvPVCQLfD0PslKZo7oDHU
lJUoLbWUGHcamkzk4tHKc7exen59KD2uCiijXZswFzU3i2H6yotqRFTgw3Ssu/RcnCVP+9Ui6OLk
XiUII9MHm5A+Jt8k1mElQD2W+cpiwpNntSZ2MkZeBddhjgrvJKSYwBvzAxTm+FdZMju5N84l03PG
Hrpd57U5jSIwNDpAATnrPC0UXBSUPQBP4oyvfwFwrWTbPZi5+nPo5ihzTR0gK/lgftjrgkxure1s
QwZabhHIhttQ23E9QRFRZXllECL+3jIuTbcvx+7j5i17A6dq8TNYf9mLWvEBDuzybEn0xRG4XZh9
X8huhQz+Taicnc5301MD+UJ4v9imwxQEXsyPPw26npo+Blv9lUL1gVUfDBxvH6bz+p9pDRbAT/xk
fG+phQLkSRgZGbUXql6g3f3ykJpcbR51t/bZD4UugvTw+kckgPzx+EBmoolu07oNzltOOv18d8SE
DqGzRCBsxQnO+S/QMtsI0lLf2xr8s8Xzs57/6uWxQ5gWvPG6LQNFQVRo56JmmbBRITKvDHt7qEyQ
Z49J9Tf2/UFVcMuwO0aPYlrjXWSRlNB/nnN0ozGt6As3PhcQ0MYksncbFVI6zG5nbVy362wbntFu
2pyjTi3jZI4IlXUES32fKQZv7+3Qc0bQRyMmnByTp4n8swj1y1wuMoeh/ZIcq57pvxyIS8cf6RLc
80TN++WlVEhIW1ktpNP3vtW69jT+LIEuSJ7SagqLOmdmzbmQRpt/JTeeMp0TdxhLpc5m11oCWhQG
jCaIq0KUDscLRW6SnOj/iEEdA3LPlUOMNWW8oPWeeWM96YOXXCVUJoFe0gffgyGBYEk2nT7pjq9Y
usZidB/YFFhty9UjjDD+ylYL1Acfu8xSH7u3nkpxNGD5HpqAx8oy6uEdIfHBOWQPz2O7x8Bd1THa
ZcQLub9VUdOLMjB60sYsgR185fkUaTtaGVEeC+5R5f29wXx8Z+JF8i4C+JRbl2G2RXeVcFsrHnNf
VZuAOFB0eaRDUCiziZ6i2N16auNi09sr9yJD/aVfAKgTssR41ZcGmXKsc4xlCt4iInO+cTHAGtxD
ZIGb6wrgYOujbrEB3Pld9Mqk8Z5HiYLC1e5KPacNEOTf9UdFnLj4WqLTO7apJsQkl4PgodixlUzZ
4hMTZcflyrnAQWm9eQNFeurUAk7k8n6LBcx0Y+9qV7+y3IrF+8/9pu9BIHTpVaoDMEmJ56AQn6nu
PSY1b95hFU6V2uer3DYFbpfWjGnchUZPSkrk1/yzDuV+oYewZHy81ovxmMiaQK0U6ictoLO7SL/5
2WqLhnlJvh+I6XRRYs83HSMyJs9sFdjXe+R3NqvYwaLRWJVax6Z9DBua2US0bUoX4Y1R58SnPhQY
+761w/b2w+JdpSwq4EgSA+RXc1FmeOO6fo57IOMNhoBwyS9vbubbp+t1zlitZPfLR+I9Bhj1nK3M
liu6ujg5w02Jkf5UYTulT5JjgM8WxMuk34J6vDndHr9F5YtBm7JdKi4EzTFILEMlxY9K4APHz6LM
hneypHhvcSyRZmuDcUODWq2aSw5qM6WrfVCHsYhcYbSUQKL5j0ORePt2gAaBLaIvdk0cb7mk6z0x
Wej0dhX4IgopKqtS1qQcD3Zi8fuoZjHiU3FNf7J7rAZHar88fcgCe44YZWEHhYthb5s7To86cyq0
pBGZWnhVUqzq6Gr2nti2Qk0Ls8XaCAkbbHGU6LASelao4IR6sW/Y2dRpVH2s7welc0Qwor2GufR6
rhZeWnwEh2EsSCEbytKXLP6NccACMg0OKgL75Bd03Ru7sOmMqeSRt6F9yjFHWRzwRskvlvFUkk9w
695rrevZ4r4pl8yGgttdqHhUASjF8lKhCwOx7fjfo0JdHRHsqNGJNZyJ8bXuf/qX7gblJKeT6grE
kDhi1dxYfI7OLqraErWhfA3tZ5Jkql4sR3O8JdawFQz53xvl8AUVkQdGlsV+2RGs6xVeaDZj19NV
ENVhSLqKQCOHUnSatdGOGSeCmiFHxLKOznh/P5/OAXbBAztf2fLffacui+/mVkUzgmhHPWkkJqVy
+Ms+UElMnefdEbLBxegGvV0p+B2QwWhtzeU++PYJnjUi5na0lIFV5PbIqybYiOe76C7jVL6eT+Eo
d4dRbW9pedhXuK9zTlr7bkxhI8Ri3dZ2kjBCmj6vczuL0GPYSpfVNzeanyhJSI1zmRvJY2vJ7QQm
SD1kvelv6yuK2DLTeBsL98nfGlC5YmcO9+CAurSNH5xjByzebY2HzH+q72HpLPN+BHBBwIgIN177
lzPoX4znSQ2e1E4qjWZRZ1N8O2amwx8niY3jriycyYgaOAnMdKWSVLsjmtAfq7UHj8FApLH15Zkq
fCdPt5XlPnGnHlDsz6CawznnuvsqhzrwReS4wc3Gtr1jZidqoGavrzLEZI1TA5UED72YVtPvP6+A
hU0GhADSQf1sg73Du+Br74pfRVtej8N0sCdZq3upnMDkY0oSJ7AMn5fdBzTAGz6yz+5BfF/unYKi
LLj7AdlJ8PJLxCB6nOK5cWDtjTnu/qXTGLqbjITZQ0adS7ZxK4uH/a5BCmIDmxYjzWJraZs9bs6k
Fak4lO2jQijmCYQG93hHaXMUSyYDDJk2hAv3zRh02zlNOiEmqjrph/YhygNN4lkDI2RmOp2i1CSm
3sSuodcCuYRpivqzjSVbzRCIDHGhtphVuNSIOw0BclxilBZQL2NSEkDSuSQRFBhY3WAz84nWOvzf
Wx9OvkH79DYrfPefUqHNtNLUmXrkyaOgu/mBWp08N9snZlaQzx0HTYvUqDZlsEx2qKznijhYJNWe
XYWNW3yjK/oGdMNAuxXCGS7lbYPHfvtBJRs519J6bfYIR2fijf7KL42JTobpZMMY26UX7ThbjWlD
/wR0/VVXRj5I7/RPB7I5WVN3+ewYGn4yC3kt1yYG6VfavNLxmQjZbuVDc+M8GNvWGtrYTIjt7vza
ghtYB4TCD8lQqJ+xaGeQF3rZcsMpHcgrtp+d6SUBqq/TP31vP3S/5nM+oSgHwm0ljAWao0GaNfZx
fKqUPceBp2w4iU7JYhGoXXdmTaeQUIF7ctQBRNLnR6fOBRtkEH87KpYisxdW5GnkYmvCXn1Llq5z
skRv1x/1fE2vwkS8EtERoYWnITurR+ate1x+MDdc/X7+xA1hGBnMf3QJqBu19B9MCqBafzzYvO+n
QZr9/u7kODRRFHudCIO3cGo5WNLhgPxT6xDQqaDPf2z6rc5FeWJ7eEAvvmVTu4oq27DRuZVkXpWg
WDV9dFoYp7pPwfUbN5HIYUnH+/HmKNm0JChzSw9SncxG37CbJ60QC01JIzpFoTzFMh7lWJpUP7vY
jDr/bflXXbBplsFGPH4WKTmGycM+Na9ZVElj3hEek8QSDX533I6lyd2JRArhfVVlytqXvLEedOkA
mU5BynHbtOIFvr7NvWhgPjnX2hBLguK57Xmof6/bAVxp2VHifM5KVS43VEieqkPDv/3/SpDCtAz6
JY5uitowWztfPxNY9tLeWScWTznjJJsj2rjJ04HMJKjdalRYZ80aGp+DvdOfzGciEt7FIhqlThsY
+peG6F1RwukAbYqsXhA/2J31mF/X9g9fa5bH7JbcqaKINoXtEAuZckPy5/T1gQPNPcjYVOtHdx/z
uBlZYkBhsq/8Cqk3Pxu9LjyyHKjAGBdBMG/hN4qVSeMkdKbSZHRMcaem3XAY9QA/QqAzZKVW/4U/
2vbYUgHo74A6Y8J8CRrC9t/wwGHVWSeR+BcgtxrMeJ4CVViuCnJFzvwuhj0I5UXTZBJ7iZhl2uN1
Wx4OVNKgTR9U368umfUV0rnBBmRb8q2Z3uQsEUQPfqpXefFzbkMn321/r2Fo/C5QvouEx4/9Xkyb
YYvLRWH/AKOPSS7j37ACY6E/qnB0Nvdzm/VhK6ou9l+jfZrwXx5qT7uJsf4BVt6+iCfSyqgrxAKD
YEbf5GRRD6ZUY3uFTSaX5wVJQ5JgOetgSugQKfQJcbADoRfgJShb6QT1p0xhcSUk597+o0naAxgh
ghB/524dX/NYgzSLMVG7u7z50hY5W77huaqarxJQxzB3wTdOCpOu2A+MSx4KXEKvMAJCLv6I0z+D
YgyWd3L7F14YjwWQSSfLyvWhNndQfmq0BDOQZmITyfzR8t/S/2h01t6QNC54BOXma3twydsryMA5
hZkd+TQ/Xvxoqz+mzHI+DiQBrd05fVQCq0CbDvRRxgYFk4THTmthvUR4ByHmzFk9gnZEKOsoCwC8
no2dSuUqkw7x3oO4BToV9rfiruNrsgk9O46NTTbl207EnGY7FSmNp82/HuIo09q5R1lZmXutUqyu
9Sjc8Mk/SAs8qGHnXBQEBmte28wiFNX+aYDx4nt+eKtHlALu4E8NR+SGIaCXt1GeWNhsedPnmFl1
s0Nsi7fwVpsh+LYW43h8mD5qeX1C0yoCVrzIKbSImsxXMImIQkDHK9UUu0pCjJHs0clfZWONJZmg
HQtrX4jHlS757KXnxDMJYj/S3prconaxOlP4K6awVCGSvAruvo5DsM4b/s0wvGKiz07zSidoGRr9
Hny4/0fIEnKEc7wYdtFdcCSMbn3K0Ai990MQhA0pWaeYk5CsmHQj/oVXbNLM7RdhCqvNAbvfF5zM
vE+0dSe4PjvFV8fLVtW5Y+PDf+RmUrJ/58u4wgLl3KFvNN1LqR9hC2Av+ac2lF14Nuj7TAJDVXf0
JHIphWhPkKOACTsA6aBp+CIMaBf/GumR/FyL3C3yaoS3sVzyhL6U7Br8Bkcc7/780WEKjunHpIJb
vOPMQW0DxG6esE1EXrq4vE8kM0b4Fy7rGhbSgZTEjAIsN/bCwtNg8RuSpT4ZcKWk6i8mrxK+sRyZ
7FDef3jdEmGSRDX6cost6rWfQMhrB+zUc4w4+FXRQMHebq39xQu/6xY3jQINqbgk5v0s7A34OYJp
SepQLjAnHOx5CA2dzgkiousGoOMgwIOP4ZGknhiJ3kbZw9jXEizYOfl708+HrYoThNhC7jnkNlRA
H5nR2BxkXe6NWsAH4a/kB5N3xTfaopdbou3VvzbDBegdWb6JiGONiOIKt0gLoJUz/Kw9DQ7FFSWO
K3/WTIU9QgsPOemfcYpsNFBOxVTZAku7YvQ2ogOPtHkxqs/6PDu/iA+jGzexPF0F/2QWzp9SErZR
ovIJt+VEzboz2uznIyCwhKwOwUNuBByJ4mGtJ80maHGPd+iFnw8M6l7FXFRZ89DSWK9QeVKV+Gre
O+fR9w6rFS8RVpzFgxqFc2zJ6QKVkLQhpimw8F7B9HnJoZifKV6viS/58JfGPWNVs84aL70auzhJ
FwREeUkk10q0pdB3dJrAqH2IcIy2iDYDqFZgPzT97JF4a3aV2c15ITs/XUQf4kxPDW/5MEDzlsid
PV6RnJbGVK+GLsl8LkUfCwfwc+ZE5KvM+7DeWeykpwsqRHWke5cuTqKLxGK1MLMV08KCipeVya7A
CwP8yCzoWGYDAi3PuqDzr3Xto2Q5X5les30JOoRdg9S/BPr3wRmQNOBqWE4nJinecHg+vW01yQNv
FnLAAlWbHr0BCOvkIxz5GUBYRKwaOGRk/VLJ5TzIOzeo5/hWundmzOHJzk1Kg9qElksVZQZi/DKR
/AdIpkuTmFqb+SMluMoQTMMZH0QIAxi+CRVFJiRq8/rsLZkZ4NprGFcXm9RBq6CbE/UFURb+sZyp
VT53HlnhVzll48MtUi7jeQ8Em5sAfSWdsQ699a9sJLY468NDC8zsBmS86AZOFT9djUzcmyvY/3of
QfQ2ZOWcOqJWiOtDjEuM2HcB1Wk6p71gEBYh/M6D6E3pIGaBre6obbIf+av0fVa3E93QyMWdwIYm
UjFpFnmz0DFCtMAp1vsygeaLnKmeMrAjSnyV7GfyfNiR1RWESZKnSCKmF79WW8c8/4nvXCwaC/L8
J5SkEYYYeqZxsgIrQm/nrCbWhTKOCK176TL3rnfKPKpNUVwU5ObwR0Ih+pB2UKtw64CcK8DNJePs
22BbqJTWbdwKrrmLeJ37HF5sqZjxuV91uyfesi2l7lNkrb64n0KoAfSpSpYe/X3TvUE1UK+Mi9Fo
9WdgCaHIXketNMyS8xicCt//qorx7/p5kDY2SW43NgPCyuBtk3HovQAo0dMXec+UsBbS3doYAytl
0XrOdan1J/AzB+tBa6cpDG454Ben0DJrrBC/+Lvz1k+2VrkG9ZpA7pRBW+iuE3riW+cfIvYPrRQ/
Tz46lgu7HSwckSelSWxUpA4bZJWE9oLeDEkYDlneglR9pwNxGhqs1+1fT+hC9xa/2mDSMtOg0bkg
TxoAuY7v5K2i7JYzlQpBZCXpxw9P94WyJyz8upiZs8Qmgu8TyDXjZd/96Rbu5tZEpzFxCMoxAQgA
dOT/zTPwvhGUniZ5SNDDwmnc0k7IDZV7nQvmiPy/Cj6r6sckZS0hs2ViB8hRDC7d1PKxJrXeeTrp
zGA35qEcio6vrMJMxfHuyN6GRHSc8JmdGG/HdjxPPS9IIjQjz8XrtNO/hz1dgLq4iAOKTpnN5xNS
T1G7Xy81iEabXTBU6jNvnCrFVw4FY0awM2BZzl5RamkiGgnwNAvLqzga3HkYLyLLmBwV3tn9VLpt
wA/GZtVFnYQJRWK0rOVVikHTW9OSaEJxvYYwFDTrH+a1klsAy1SLApzasQyLx3l+JgwAbnkg95xw
kw6z2bEJ4ZzYddV9PlmuAzWIR6cQ4ld6KOQnoJu56OHpqTuRuO8RRcyR3k+ZuVRZZK1ETEV5RrFu
QEPEkocEFkxiioDKdSZXpJ41JYYZoxwOnhVuH0Lri1806BbNA5QPjqSCQlgS2tUzMFl6JwKP3uW3
6buodUm1wsnasjffjFnQefPkL8r8oA/iMGrlfkIjuzXhXb1wkci5ds180bHtXJ746+oau8QLt4Nz
R+SP+jXk7FKCRZAOKomtRAtcd/fUN/ilxVyphW6gKPAeCWNzuA42RG1xz7VWXpNDvVb1zM1Q9ndC
OH7To7uWMTTrpkrbUJrBXQUu9ljvOQ9ns/RXOfeX4z7hETp4wXvwa8d1MaTmeXihGnUHzacOnqkb
USmj51vko9FLTCm7Q/JcuOaXLUbyfHwVSqEd6XCxrn7VMeY/C3e0qbb4EldLrnSebl6AE0ooTb4h
HbsgxNaQAShuDGx90erVPVg4pV92I/M1NIYJyJK+225tGD4/3x/3x1u9M+4gz/MsG5WC0fGxO5QR
/e14VuZkM6IgH73gzqDCQXky/KjMbuxzWq3m+JucRTt2zfeZIfJswv5i3SPoCWX9uRanDszoG7K8
orR5nQSEx7cOYIlDnOZMT+CZkGM2BPLsz2k1ZdKZFVmHzAEB5TvpSQtuDlhVwd2nZvGekA252hhC
59yKNYP0JDrgGemI+2XPS/GeYrvlepky9hw/mNSpDg4dG2vmaCpoZvzWO4n7zXA6BybdmnuKT117
G/T0eMb09J96DVOFZHXxRiBEebyw3xBZt5x+Vv3WCfbPeQCYB8nHe0cKsuRbn1APQwIeGQR7UMnh
s9Sgnmr7IZcJmGhvt2XRd3tUTcvN60HR8gAt6erk+Ab5B2Mjg7wdhUFM57eFs0Q24LxG4VARfXUg
jRd1rT3KJi41Eoyw8p4aFaapcAoyj526QIUNlTILdnZPD+OFUOdMLoUG4MAo9fGQpsUH49qm55R9
aMmUeA6LKbduhY/noJO9SrcwOTDHPY619y7JjaXS8EM9MfkNt7WP26tIi8Hl+nqRY+Q+U2qPtdrN
UUNW7JDtmR808P+bZJzMa9IygoP7Cwe/OuR/vQy0NFtsWzNSqR+YoghinGq8j4+qmvBJ6WEL2Ytg
NiSyGI72vtoomSBw69hyGzjPtx7pOAOY614RHtsnpunEbyXdEB9y61/hKRSRr+9tBRScDrcJRISP
p2ETqp72ZReek1XSwarnK0FVEIlTTwPFIFz2RlrqqFg5qptrQY6210E0qMaOyD4sleu1Za2dDnPe
IjEEtdEv1mOIVQWE58e0syRuauSRUYWnkCJJbjtABEqI/OUGtxAepMGi8pnvZZZJD6aoh7EFW6tW
zFB5fF1nXbC2MnQRKmFBdl7KSXDKMhxXKFCpqPZa1yLJL0kKtuddgFMqSIg7JcZN0mIY5S9y/Fxd
EUa0v2ooxi0l3wVX1wav64pQWjZx2Kk1zY8XTT7MezPkEBp7vbp+qGsYbCoDfRiiFSoGUrT1aYfg
XzfEEDAwwtPalS9vvmVZ4pKc+sKBqgz5fwgljb2QSajuc0MdzIYyaSXeAfoeih4VVkIu+wOUNg4g
3kgpzIJY/QaAp53CtYxPxz4pr/bLuu2bCJ/xZFzW/1l4mZT0MdJx1yEYcizcbcW+zZMwlUryrTKf
Bp4EYnb0+1XCjl1rtbFKzUG3cRxT2BC5KcyPaDXbVHi2K/7lpBHXhGfU+u9DVAg9DkzDy/55cF1a
baBd8dzJPeOut6zfkQ82VEeJd7GDOecaKiSO5ExwcJ7uP/vAnIBLkjjLfR4haYXXnzHSo74SDgdP
7285rmR8akoLdGnZHXTbyyR7uYTm7IWbAGjX+ZscCAOE75p7XshS0NresX0TjQtWidyuCeenMxQt
xk0OmPY+YKa1JBEuZG1jFJx0n3uereT2kv8BFLCnLg1iI4C+VOuNyYW4ZrOfXVzNkgnGw2zqAwrl
LdKVzWQmVSRjBivDVePDajjON/tbrHiXUrIow+/iVhQNs9sbDYAAG4d4yWjgmripE55VZFEoenLF
FGpzzfcwfKY8loIJSgU0cQAMEiKV54EFpW/Ah8afDfHLTnQomQXQk3Ec9QTIN3nv+bW0/r+PWnOL
UoKX51vhxL7x9Klh6RF+kSMTuJ6eJar5W3iJddXGn8uZXe57ufmrQRau+jxy/j8YMjw5ZzOa0ij8
M+O5Sr8qtPoWt4MNq0lTnK+DmYRbldWfa1EX5H9Vxai0zb4dBxBuG8uB8uE0Ltnk6qIlhoPvvV3t
ttxHyLljFxM98TmSkoP6laMHyqtVQJ3Akwz4BFvFaLQGx8SA9Q6Md8EkUEg8xfW7XhfHGfQHbNQi
Ks+mXnAzceK5it41hqWo3+EMaqTtCu5kcqbJwmIru8Y1gRwhuuIcE0v6mEVJBUXksTgKRDI/kHXW
GUsEmrDbeddviYxum1Yv1OpFC3vZ/g7OW0TuiJ4qPQzLOT8Xi61u7QTd7agijq7z3v/BMWu59BMk
pkCkLDl37q0ZliTDmVT3cYdjQlBbL4y9GO4AiOouM5K3489Zv7TZMwSoyOVpZVZjeKXivAjpjBmv
HM53eHm7SIvrqY5slgn3zKBPkJpC6VRUnzB72N0yTDNdxIvezCPwcyI9ESe3ude7fRJJKLGfl2LL
XTgAKaU4cxCwmy+tfeeH4MMbnTN1aICDHdKNVADUWR9VapssC1An+UnFZWGoYWLVbzt8RPuyIaBG
0DsE1yRjgQRIHiZwMrxmpBmp04JbVoe1JLSDmgikSgVV7YDXBgfg0x5JFC4h4nbqsjZZGqCE2wTk
lB8tVLUwvxnnFglvNuU5SS3nVMrMdfrLz9GE4Fw/xoe4R32lBvVxEt08UAycKi6yRbcoj3uuP2/F
j4f/ppX1dWbTohzH2YTWwf/1fFqsg1dajC8fRCUEl9yO3fWaaoHtPq+rawA+JWhQk+qleadF/ozE
Nkj299uKy1LgSH3cudpwTh+YX7xQ4ww5A+b6xHx33fN/F+Le0raXzABRW5vIqNlN+SQo2TpuOxPf
JeIE0CJmvOI9igC3aGSMy/yLj7efUJE+e15jFVAry4In//FgiNVjZoQ+/+oxmKOSgimT7SuoItLG
XSVdGFQ2pAzU3ShTgaQ8KORvH0tTxnEp1oJYedaVdisehqZ8P4HCYwi3twlCZxTWmAhVNZoz3xaq
ZWDq8an+nT6SU13k6Cn2EBywF6FhRh/O6qGvPghrMVI7SVGKkWnhNGBbM1OBIBdjvkxFjrubJm3G
zWuHiPurCPQcsg75j5JemRuMp9TCGut8BH05JNfE+Vh3v16WMz733ER0yU8Rjcewa/Mymif44oIY
gtzOETz7UMI7999Z9mTqiZrn8MtoXkKm96Dlybo7PzfhyCMPuswDlRUU7OiVXNRf/+Nm5KoEA8vP
4XUiPELq8qO1M9tqBJrGHbq6cj14Wdm0VDHZFFj+0niWHR7TillOnLW/IKhSIeSm7sT1EfOF/igW
TmJmSztgKeeznG3c2vmS1i/H0BAsYr3+kOGV8qxK7qo6AVrFtrG3enXQECEH7vVXjPH3xoEzk+RR
Pg8TTLO2b+bfT9XceAWuj1llA7H0AQ6jrebpLyvyCgxBNOMhHhFm8WEsUUk8iIL2vM/hCs/2+4pZ
nIJYP3wFzt32gTh+oEBHnESXU9FKKbIO1MgqzPxmAADPw5Vy6bf+PpAyasFz+pe5ixKyg4V8mT4p
8Q1PxpRqEeEqJaMj6kuU0thfeJTEKBosnIxxLM1cXaOMQY9FkFdJKyi2xvF4E6vk8t8wPp3eBY0j
XyNQ4zj8MPvmvb8XpByvKmn7tqBYcdR3vtzmPgWCWmpCQ0zQ6wNFPcKLl9/qmsholqZBZxMRBj1+
PGSvEg6KMxjGXyMZjH8CX/K+ejNNDCe4tZ72HWFYFZ7Fjlk4IqoODI9stzT2PAIEbb9nuNp2C3/3
s4//lw6BxOgJoNjIELH9Hc/q5gY7ZhIQMmSTuErj6p9/VFbefDEsqUoVE1+lOC56+Dy7twN7Hv9T
0+0m22gDF0Micdrxox01taw/Kqkqiqc5zjPpkcnrcamPK5u4HSPZWoWPbuhIcWvJnLX5h+klfQWz
9SrBTvaFWoA4sIQloebISV9Z/1Q5wfZ6KGQCjwXx06US4vXAeLDQ7tnYm+7TWcI03IEuorFqU23E
NK4M374R/iklgsljMkcpJ4pBZq6uB9fRYK9Ln0TF99DL3solODuaZSWxNhY1UpZv4CkIcUmc30Cw
KF1fBJHcXoLdLOE7jojHRLtP8mati2rY4x/16nfADNT280VHVk+4Wnms1YeXVcYp/cp7XuppgRYn
T+l0fiNCrCtWnxSNe72rNU4NE+7rn8s2u+jqHmfFSch0Wzq/bDjLgFPbBWlhleuawWSEzuV+k3Vy
1OsBPc0g9jaEddkdp89Xh2F0gtMiRWk3vq64lQJiGfeJCTT1/pNuTxMMhERtbMDf0Q5rK8BrZQkx
E3wt2FrkoFcIK0ePXeuGCX7t0U1vg6FQ58bn3g6JlgFj4e3ihM4BYl3a8Sa3BAe+6SDUhpMxtD1O
buZ5BCp2ECRcNfyfDp3Q02Te7dXG1+KzmyV/D4KqBbaI6ZOk7EIHoZPT7l6eOtXn5UZOz62aExYw
SSrIYp+4GKzZZASaaPEztIypOb1r/q+1MT6K4SBEB8SsEDKKNtLHu8dSmi9fsJq4QxeS/DHpkYYz
SKiBbgNRxhiD45oO3io27gBWZXscs1xWXEVWUWgnXE3bV8FZvPcEeYaEwzslAagy5ad5InY7zHkQ
7UTqvsjLSoNsPUOjCVxfCzJefGmebML52QZsTQzf+DAlwnGDTXAwVkiOxkdwiNe6E3LMi3Zex2/p
x7aBGv5DVPdmpPTllTr4n2HW77o7Jqxc71Z/k/HUhos98eqtht/qCruB3MO429kmJ65Otnm+xm3w
ZFsPzgTDD+0PLM5ZpBUs1e3wmpjkOQSiKSwCy85GfPd7vkvxKbauqavyBAZokWivhfq9ZYA6eS1X
Z+yMmDv4KhVf0hE2AK0rL5RnAyiSsJjPzdwT+/Gi6wG9uxa9BfRBKlELkAq+GzO3mj/gZO7+bklG
qHfPcfTEdKQ8dWURo/aG59M9jN6N9yP4bfkas67SWkDakQXttA/acryFX+WfNtwz7JLdEpb0LDk2
JNeRcMbOf/4foOaBasKuS0uHVIpFX58DO1HD6bpbNNQFp3O4LvCpEIxVwkh5nKp/Y9p/vx51bPCC
Sz83Cwh1pDqY392hqDTHDgtzuVaFbuqS4ugJbNwFfiziL25nQol3/xeVPzz//aoivAUKg3yJ+qNn
Azz+yB9Ji9SUx6q51lJRzUQN6HRE+nE7OJ/46nP3ADzEzQ65k9sRujQPRzofTLrh0b/7om8S6d9O
QnXB5HQtTQ4yknyGpOlTGJ+aS/wKr+UPsFtKDMyRmQhlwhH/jPRLxG06XI/apjZIgHQn1LngWE3m
vmKdvEk2GQg1h7SUtzn0t/q01DZM6xg6kr4q7Uav8XQ9vAlxdj3npVT7mKbUq2DM7JTU9bhd2WgY
DpuBRRDG74LPtaQzjcg8S9j9Co5DtxQreVViQ9in+yc3d0Ja8IC16sWu6kbVe8c5DBE87CxmOCuk
pxH0u73X91L0L33gxCsSQXLcMneWDsiDDuHm8I3/UnZQ2uWRZ6p0eC/pkdXBtndlVIkcpDwvrQVr
s3pfrA+zqBIw2uB1J/STS+72ZVMTfZQeCq32HQdOgH65sWeaY0gKcYCel2pdWve1ZBIvTSqLcDFU
DrVFw3gJhOxRrWLDCJua9FrwgfhZ0f5veRH5Td63HEr6XHFz31ENeca9ZKGmdiqupSJBac/oddM0
AYHez2fJpEp1PENY8xytEyNczR0bSo4fME4BhCW0RQIIAFxtQyQDq+bbccUZ3IwbJYd3a1DxZnpC
ghURc36Y4dxHTB7fFw/NY1EVn8SbY5QL8XtQfosLoAitX/5GmtU5OFgsW/FOB6NCGHGMjbumQrNI
hcSjIKM+m0IrtQJqByovRa+kKpteb5k3BpB5W9ZJsus/A+WWEqJR3knQ8YVfpdx+WXdj0zXVkdaG
ButU2xH96qihqkzW+Y2Zzdi5CBb7z8B5x9W9bmBWwF0I0LGBZ3lBWRko0/4zJ8HZQzkX5rMkkAoK
8MXSwjfS1mgOPt0yg7FE3j/IpW3Z2on0GTWGVS8cEU9ODf7p5GAV7e0pQivnLiSYQkiSoZ7tvU1V
VIII7aW5u2/ZrNrWBLk/pgTKSyIkt77rCmP6/IIA6gn5lRLNO5vGzM3T0a548x85222fk3JADlKQ
3j8RahAYIqF0rWxkoET1H0nCSW2UZR/4N1VggIfSEp1AGFene2WCNqLFotNxYP47y/ox4/KDIRsj
mDSoNmnmA4IPeb+T5b56RoS/XKczvwac7uFtnj0EZ2Mabp6q+2AJO1Qp7cupa3BhzT81kftsC43R
bWtGIjU0ksy+Xs5onGbUD63tyuawb4f9YFZ2mf/WHG+XpkImJ4aj/40nUoQdL3bknUwzINQ9ccQZ
n/3dHE72T+Qu8p1q25lKGzjDdn4hbWv9gRB+kbcK2LSu1KNFa9TULUYpiei9DUfiLwz3qDH7/ApS
BPt+/MlWYjurISoUJLBZkuS388IXjq7K0fiwhZ93Jlg2seXv8tqmAPXbcbz8Zqjh20nYH/L3VdnA
crgRdlAzIaxn6+B0ZPD8p1OCelRXPzQcpnVdRbclHOv2qr+csXDjLLhOVwa76IVIy53Pnp5ywkoO
bBzaCkS9z7lVfRSUfwKJQJukL/c2YdDxBKDp/04FZOLp1rKCuCk1cHFXPajrDh/S2p9e4avRBuFw
qwHjfSba3yxYze5priiqoq/1zUIFRCMwZNu9eFWOEFkxn2icNkSGo64h43uyiDcm8XefgOomEJ6N
AiFD+JA0XWZGgxWmkUqQEoT2KBTbXbS7zsRGH4Lh6mp/SO6kcS06LhO+BEYZZsPpB6IchPTWD7K6
/5UpiIKiWODy3TRlrFhWl2nzWspJiLiikRXE8its210rMdU2yviWyOw2PakRVxlkdbJx5C/4uvys
AcQqq40xso1/2cdIozB6dt4sjsn0lcMi9h+Gc1rWj3ivX2X+Siw4XC/8+/1TkLKrEteMDr+5sNCf
7U77+EwPCblw1fy4S4oIt8RBvWmf1eUEjwx69rm9P9CiFB2Tg5ZaBxktxYRmxX+oBsuKmzO6yXzZ
AQssF6neZxeoZTMQG6IgbOdmVbS7qFmIWVpLb+ZTDqFx/N1xtj0+iAcKtvli/ue+tJG77EdBKbB9
QcJkOMPsd6lOgOpotmfOjpPJF9RerYE7TkOTlebRNuG6Wibcme4R/mRZ6IFzxZYtmd5hyX3N1TQz
Wj+7gWv+/XH/nXSgAVbkTz/mE/frUrWhIa3UrT+ESy4S0d5NiJVbm0c57XeQEmcH54JpJdWDGao9
TkZoHGmFm1/+cqcCbsqbcEjUZ9+3cfdDmYPXt62QBBcGyAqcsfPBiv7/4HIHBhH68qYmDrzjuB7L
CrkCZ5jEMWtCUMdIiaErH5/gVE8TmGFSnBwZKAvij5TgiLC3XSvtnHklzhoAzKfKSW2CfYtiWF+f
5a8cFJl5j8GVt37aY//RIcdECnCiUIv6A3Y9gj86xigmkUhCUsadEFwBTnL7ePf5PWjkvHd8RBuk
+BgNkEp+P63c11EeEW0kLTl2CKk8IIw0bekP1k05WL+hO49HcIudUGsf3NJ02YgNto84BKn/QA2x
wN0Zl5U/LrUx6C1j3iwePqfEdr/QK2muPPbB9R/ZK4qQDt7BtOU6DhWHl4KWqncJn7OIUeJJjEzU
utWhWdXlRkT7sZa9/M8sAkSpsrcGic5zrnW3EdkIYfY00CW+puyoxz+It6aIZUjvRG2sQRDtbYz9
TB7P9nip1KggctSU4KLbqGFSpV5Cg44CgcyRMBpMKKmD1P0XiUSaSYvuCnGzJq+X3BnlsjCqKhKX
USG0mLp97fURr4HlcXF+HssQUPmD6/0DTkTtkSSAvOnVMKR/e9mp3fbS2kvaInX8Ba6tqCmstvt5
SpgHl//wV+dROpv5FOrVZShnQGZv9SQVdhdkIQd+u7qRLJIy4QvUAbmvtUwmo1pl5QFQMKAJh60N
T5yqN/5Fb0Yep6iGnlLjFlmAeoxTPgGaj/Z+snc/Kk++hdPqPZY6vtDiMO++MmDhD9sqQonPdIu5
QOC/NusqslrSNnEJ8yQkwZi4LjXevXqgQD2ybxUZ3n2jIa56G1z4WC9qANFW1V4NqNFOzQOPVy0m
t/mLfeCE9GPeemPwFfyPEDDuRCVtMeT9Uo8fI4PPUoDvcGLJD/vj6RF07rhCU0JzZhtf8zXuLXTQ
h85aVzWTcHaqWqM8/fGznPykzPL25PhLo9NHFqIIcXCPSQBE3gVsU49wmy82c4qwmhUMBD9iFg8u
xpZhLhfg90o0Y1uPVsIUToEBcTbe0WFEsNNhmvgW7Xo/OYXpt5xfAvt3lsamhZI+sO27fMsRaFRe
nl2v3QaVkvJV9WVf78pzKOFWVgXSadkL7j/D3AiVx5DlNCwv/cLNY8oUipH+qiQE8Eb1/tCKMYd0
+NSTXxFjJQoXiaTuZ2wVdMlOOFwxb5Nfy8WLnPptNzLj672dsIkOBgdY985tXNqVE9TgyvIZVUsU
Y75aZ/9kF/RLpZv9XD6Kwznt01lySOvYcdPrZX5LWfoXHGb/BiMyzKAJm8r/LMrky+DBBpdosl4r
VcBScm1WajuAc0xy07NO2aDj0y5AXi62yLwmVXv7NlOIKHzjaQ+OPD/wdtsiSyPHATbJ0av4+O0d
w/nCZIaufnUF56vkQ9t8pWTKJ4FfZyFCdV0uHyvmCgi0sHoAzibzPJjun1AwIc5x2Sb3HGKSrX22
9w2dx2/3f0pIRkCUM/NlFgsv5B10ggoBW2pe7AVzCgdm6MCXSZ3dEoVRpAT1NDoV74VIU1I5W7DU
rT96mZKFuXZv0/4nKRot7QS+DsZ/S/Jn6+fYZh5gBHp3Ykx0wa3fF2QwZXAL9BjtIVN3bfmVf2Lk
/jVXny36LMoTmY8tMyHb/YIcKgvMgzkJVnm166X6t72puvwduFXii4RtewFJPY9obtL0H/9coMVk
tssd9ZnfGKt9grul8LkOVETMSq4Da7/Wqa5zWabja9GvF4Hs3E/vtESDx7d3dwOHBxqKpL/B2Cs5
DrFkC3oaGg9beKo6IPamTOCvBQe9pf0w3HCLZ4FQxv5XOwMeCegrSjjb0u3Upx41zi9oNFU05hki
j9p8ia4mtLfbbfN0obzOmkxBPEbME7jLZ6JWh+stO7QiU4+dDAbZCHBqzZ/q0RsfgJv9/+RQFbun
QLByTSyi/myMG68TnthfJwFC8gx/qAGinCa9S+mEDpWYJ+pP8SIvaAbpRJcn3f36HdSpLf4gdo8A
65tRHB00t+yBDVxbQN7G67QMrsdUNLU67e77C5vEBq0BRh/voKA/J5ztvj7fVUa8BAVJ4jvVW/hr
GUbjX2UiET9RZwq3G2ef0/GP/lEW+JvkBVF9Wsykv9e1nZGV8NN29zG0/MNfoiPkEPR6sCauVKAZ
k5u7yZpwAOJrFXDv0GEsHtCZLX6JkheaWQmjL/TjCOg21Fv2w8tZuOtAjcmt46vRr6Yyy+OeuxU+
1L5PL6XU3xxm32t30IKx34R2FnQ9fbxAg0auw9QWvjXP6iJGC2xOJsjAC3M4X1UyaG2dO03IVBvk
d1lR5AlemxjBHA9amuEQ4U0CPzkQyus/oEwSS+agN2CA7WWAm28ULkVTblxGKPoUd3lidiS/i+Os
isop7+QzwSh9+GZl/ReiAPnbFUshLIEyamXTIQ006Yf25rFzM25gWC4wrM3w5ngDEVlVzfsx6COu
hFzCMxLMH5zIIikBf7iE3eroMInj9sByLGqCpAuATSUoK8hdLkPgks1MN/8ERz2IkjNx73cBcEkn
ytxPxWoaOQToWCuqld7jQu/NFPcUaMSWcRybm9Aa64uqbxz0eGxsrE2B7ncyfJF4eSidYc11jeyH
cJqDAqiY7vlKvaPYdnhP9NKQNVe9XL4ZPmzOJ74xkRxX4U5TAkz4w3Wj8XDBDhc8jYv44FEFqoI8
Zm7C9cqXhD+yadjxbD3mkh2VWQufcfs+SRF3kZv47rLtGaC4TpZ4d4zqA+8ka6xKyGGwoHUfvsbD
+bOVW0MqEQynlXrnbQNJ8REkv06+IpCxfybJ621stit5QWXGB+u1SqBRPcAoO7RdSBvjjxN2Os87
tmvohL1nsjBdJMB+kWsaRhDk1Yu1e6dv82atuuzaJR5WP4RwlOHUIp6GCO0KQPyBrl97WyKK+p8o
2iP+bSHV4w2bhhgjNimIv9cC0akT0ERNgoBL+9L9eCV9wGVprgMz/l5uGhPCkDo5Sk87zC5H6K3a
Oxcq9VIKH7NhcFP1mLZhxzNimPLoFZTaLfUHeMtCOE3rn5DSTYAKoW/mIs+yDQ5ucclfrSnHl1ci
grdc8kPJ00Rh6WtDoYUi+SqF6F+o+bHzlaD/h9IGUT9cdRKfSLEro5lUTJY6wtn9OFPz10TOVcIp
23D8nJ6F/Qfm2Hpj6kWnYh/j+tu99Q9WTBE4UBNan2cpuvdkG3i0g0SjU7x1TUIOfOSlpbtOHa0u
RD7kC/B3ajEhdDZGzFW/dhRAbIU0sTlB84WzRHLddTRuJyidyTefvwUG/VqpwSnLy22lJp9zuw8f
5PE9xSYLXIah5P8qeCkeRkK9YYZRzuWLysdxCizh5YXcui3MuFDgbuQjVoOssR1XMmqcfSFUFr7N
KRrNhF3k3AkI0IcXeQQeI/UO6SgdRlH0zFX1VsrNinmhb7whIKkcG+ZowZw0JlpVrR4wN+lapVId
ylauC7Y5yhv8+oOgtrEW2tJL2/3tHyIBu1sLnHOHJwO/5081NOoMze2JqKI8QuaMJmMkaspWQ2b3
aU+6u1kHP8QBrjkCKPXV602F+6Q7WoXS/S7F/On4oQWLzoG1uIrsxF2UN198/1AYTh686OBqu0VV
XLJK1iDvdXWCMjDJwq/SFpHw7BnBa9iQl4bO5py71PeoEOrol8UcxFHY2DevRjIS9VAkyaHcupFX
KT0ZXxCAkDEYyFpwUf5P8Je10NeJyka/yLXfE2lBP/q7RjiBI0rCHZZngc/PDJ3Eu2DjDqgfk4v2
+GIc4PSpTwIFEh5WHH7EFuX+WvwCO+bju2udDDU8km+wz03FyrKcLaGHPtZ+HkNEzDrizf8u/IDy
/yH5s2Ob5I2c5Yy5IMXPkZ9TvDSL3muW68ZNFU18rCCThz4EiRJU3JARBFPLObZusjQ3LWsgRDOe
3uyh5n/vZRXZXgHccRl/jlL4xmcwT7JhsPAPbSEYLM1X+SiIpn89dwZZc+zqa1QoaBfzDCM/Athi
D3ZRgI9xtbt9GCnA190lb3gVdXjxQ0h9XqHrfRhTvUA5pdK6mWeoJMYtEe3kRh5Jeqa47aEIFaNy
r4/FQw/BOiJBvQx3tqm6lF0M+L0abkUzMk+3gc2p10vKllEJ+UrQYsH0ICpiTdqfKNotVwpSBrS/
YYsA/Skcss2h/J57+3YwRTqOV0ARxkCP58G+epIQjpPcQXHVGEdBX/+tWVs2UjuYy9RIrAAH+VMK
emk2iLfneCesVSFcADEnu5MKdHvfO9k1lgynQWS2mrKy3UVBQwBZvKe8d3qyaAsctuF7TERl028h
AMNo9mvCA/vKriOBkgb/642AyTRwetPVP0kNpMk/aBiYUtwlPsISkjDo6R0jnSVwipiSs2rIQkfP
tD/SMV2E/ekUl5EeG6/P0emv52rjSQ0787aJA+rqXmjFW9298G+pBc9uT0SBB1okEDqRuT5Z/l16
wyN2iRguPNbvYQVJka1TfDE71FycpApUJ/BqZPuqy7tqC2O52qFn3FpyD95y7iJbD+W3tKhti0we
bweFLEkeRqF7Gt1C0USNsDinZS/f+HiTXzK0A06M8qvSUQZR/ym/dmOl9x34CoKnIE5nQ+C/Ohk0
9IS6qzENo+YrkVk1i5oczjPTQBnpWbm+wiNkY8SpLZ2jAMWxFwWXafYaOXarRo7w3ApQU4NUDpY7
DIRMPbt+4fOPTVRto7WPX8b0SSiDUru1OZc92qR6BkDvY8oHPc8MbdpEcoxkJ1Q0OaZlFa0oVj9K
rEyFlSzx6LoYlYGdmJfPwxRlGbeTYJE3146boMh4HBarjMOK8qVy8ZUjelMwNPwla167JLduK7Yu
vwgaV6GeKSLZkcGR5y0ROyyEAtho5juvHyEDEQAhkCCU62RXCskiT0KPGl6+KN28F9cf5vl8C14H
CJ6A2dzFFPcVhtSh1uaSLqK3Uo8W2wnFx8tY/ATJvYLztkKuVjdEdmOK/TcGEkvIZNAa4By8hiOX
sBO4fLo1PR2/eNFRcWNoypojPbpDWS1ggTtxs1iNZuJM/Ws3K9ydGx53i9ixjZlWIfihGLPsOcV9
pzXWSQvh98LQ3eklYpkHsj2stEERD2mQq3MOHXIgAIwkyDwTGOo9tI4rjwMlCd/T2f/lI3VGHZhP
Egj+TDjf/47iCj0OdOGkF9kmmMTNCY0lw1aFnoF6luvFgB6gjSAiFXVncOdCJvwnzbeBmLAbxOYd
00T3SK2CIGsnRnc6zuh0ZaBIr4WhfpNMrIoYkucvvG3N1CpBDkU4lfdttno3xvYtWyujr9YYedSh
ePVhahUbnSXXpUz859GUgKgxa8pXMjFUbX8BnDvtbjx4rgmnFbaSv/fgMkxNqvOYpXmmxkV9wS21
O3zGsRGzrKmRPhx+FQopcB+B8NzUATH07BSBGB2p3sr1AJiqPlMJmhdlvUrumFyVe/3AqxqaLeRz
eBfpzppHoHL1zeJVMkA78rLRxN44MzV7Lw/R10Vc9NDBWFf8fyDrbVq1ylipwE2k644q3/jvRbyl
lgU+t2ulrbsPtwRYngSGmRfVbr2BlAP7fVBcaerxBxG7Zt+vs6SJhWzdF7tVe5gjvGlbalqu6g+z
Sktef/lnwn9U4t97TgxuMbT52oavfvLHEvko6LffHfiXXFe6COVOgrVxU1LeIFiJVP3K3sgD8luA
skuIbMfyaUwrvyV8p/jD4MX8n/19Ku+M4ACvY/BjVRcPjovsgRz5vQ8YYNjUiK9TuiYso7cvL6XN
lSGeWZPtV0i9ZZgWKmxXzxuX7gICfxVBzY66x+apQd3MN0yDz7rfgfg3/MQ8p/dRmvsbhIQJ7Pp4
9YAUZYh+llnjsRcHHTIyE2Q66STqlTmLn2rb6qP8fQCtwYmewwvcQyNNbvuteaq/NFsHu/ogm3LI
mLAaEO3RUwWIvUW8Yx93kFN7HK07MJQ6FfrJJRcVEPCCExHbPoF2Rh43cU2jrehXYC6TUWCTS7FW
fHl8f2+jEaHXx+CUjJJAmKXbBtLDu92qIcvWvCK6Z4s6wZaMuw53YoaanupNyf8ClC5jabMypeP1
EwE5kvyBVunjHcAcsN5j26V0HzkAB60GoGTfIkB2lpjfNM0DFHsfAsTQ7qdDdEO1cSidgYy/mVUQ
10iJn5ZPC6dDz759WkBPbiI8GceyEgvXMYGDTRwDKYzuKvmzJy2EMWGhMqRd0bvh9DkCXKX1AEbo
7GkTPF9JoVCChWkFbnEFCE13c2KFb7dVxrJ75+XAqxGW64rHTPc5olqHQN+EzsS9aa2OsHyWBZp/
5CK0BkuaN3tIVIpWV4fNrNKe+5SyAAz9P+Tc6oMBkirUJ6kNfQ2wpbWSRHS3TSs7xhtO95got3MV
zlbCLqByO7xLp10stenXne8jXociC7arxY8qw/WAoiOm8QL1PD0m5S2Mc5Mksl1JrSg8lM1JMtEY
eUx8G1sK9tJXQdvTOKI3fAcu/ZvHqI2AFhv0nz5t67bDRo9dgPgne/7LzvYsoApmNgOQ11Pnorrd
HjnhsVZU6uZ81QiVdv846NBtscLf46t8e16eSAGrV4Z0h+3qy2J7rL8AjYDgzYeJ64gt5323HU2F
6ovccuY7k9nB680hg1rJnNvrW+QF1DMOhQRk02s2S4LF+wq89L2XAAhTQFVRNnp/9yIbdkZ+Q98i
wFsWJB3P+IHpzXo7N2cfPgUXPuC/GRYLvUZB4TBY9SuhFmuxnVAGfR2nzm09VFFqAPH687q9LTnN
TwzmnitTbE/apHZmkJDIWpRu2cY1Fjw5X1ctg2NLND45eLvkYPjApcexjQAE7wtzbD3CYq2aVDkd
/jIRHe6RXhaBVSjWd579gpfDYMH2hG6otKSDPd5b156+Esr3Jg2O7ho9GG+zId1Ym6tJTCo29dXV
xKkK+hOW3ERj4wV22BWX1vwYDPhu7gEMgCzSUPJAfWoJbXv/pvUjh0e41kATQtiEDW9x+kAUcGNG
B8tU0vdV0e3K8zQJMWCd3UxE8BYqQIpRy5Y0S01MulEugrjfs5sbLKm5fbNqBd8q5ezWYbWnd41p
YXfJkNl/y7HUCI9HSIFguLcQemcteI60+gasq4DV4Qqc13HO3/lEp+lLH7BPU8EGhvQ+Ox1j5y/T
Ix6oW8wMm6pX8EgyOuHy2//CvztX7aPob6U0vbI1hwnrlmLhSTEQ7cb9NpAAxchDt2Xf7UXwO6ba
dj5+MWs5z11sMHbNA5TSdqzElZF8f3E6lWlpUCBuPe8or5fZK3w8wp5ZCdQ7q7JJyH18ZyHB69wd
e+95RZ/sHCbSWN6ViZeCPEMQFXAzvpctjmZ59bWlD9BBMBDqkjwN//7p4I0WlpWutXF01i6Evl07
hk64hOA0ZY9GAJDO7VTQsz7tYQBzL5h4kRx9TLAWmuGyZj0TaNYH5JNNOFuFfoJvHnwo/nYwyDe+
F7RkN1vkO/S4DhtxBhEDXCIzlvYXHS8wL0lvKCVvx9B9SQ58pmzaZNvUVdMkPgIPMDz9znPWcj7A
jxbdAF/RgjIsm3eFX8shNHFxRveDOSvMxs51mVSgEFdyjofecs+pOTFCjaqK2zqvlPTOFbD/r79F
GgoK+KSAaHOf5+bpQ+sf1P+PdZE7oDGKpgG4nI0o7wSFHRiSxd+Z0PpVHEgxFjKNOEOuTlS9aJ7D
maHXfW3fipW0FolX0t3WoSiqlEP9xRqellm570xwdELKSxCFAM3o6R3rpUn7p9BnsL5ei+XTx6MZ
9lgaUE7sF7gSD2IBL0qSpLBMcCB4L1cYQ858Sw0aa/pQ4bIjz7US6TegK48kqjG6BPqfH1sjmbnS
m3Neyo+c+zeg8uCvlSNSKTCzGssr+AFr5EbInOYxjRYL6zLuStZ9WTpBbAKTOX7IK14vh+0V7uTP
/v8uZ69kFHiBk66USCkvuq2Wh4h1Xv1kSee+/DCwSiHK3khZx02sTteT+r3YUQZf+IrDOFGXjXBW
MCIsmRqnt8lPCusUw1UMr3BnnGCFZoHXhPA4pZwyorosrnyeCi/TwHzDdXchtMvY7NSu5jWNHEJD
MFerb+2NtILAbwQDr0gZ3i8HelFUFFGIS4Fq6WEboUIZriydUOND70dVU3PdfQYbW20cb7NZamZU
sUhmgflXRnZbXCwqJA1qTkmaZm3nwsDRtPmePBtDTZIs0jnDzndKvu2vfBaYGW8X7HL/pbDGvgLl
gNHEBEA2kzeZK5iRFG35M0npkwNDn2Eg1UCt8Zpr5sj8gM2MAhUubMB0uyAnC6bvQc1qJUaop1uU
boO+ZWyV8YpIp8P3RBn6l2tw7ECrokwNCS5Pu/cqBDFHZKlBA4VXKUI8Spg29p331o8/MYaTc5Sn
UGs8tuK8pqVlrUiinE5rppx9VF5AP7/8TjxfRvn70gEjjBl3brYGSe1rClskUfyfbXFVVvQF1Bdt
e9nJkTKtKUGtQufDRFGgcJpdd6s8k4QcxypJPMH6o38zmlawTNUCUyDLSbBj5WYm5MHqLS/MqlyF
QdLUKEsIrjbLDnpDE8QmqjJ6O6ARx+GRioCpyy273y87Yl2Gcl/dypBFRsuxdQF/wZntnmOxsVpr
fbzzjPPDXW7WMZ6dt+XR4N2BTmCTfp70Qsmx8NnkVgdiX47l2EJR9n/cwIoAkH6GcNpsmYqtShlF
rf/xANM1vifNaBw/bb/k6iTlO/ewNDJ+X5EJagF4BHVZIIEieD5ykUaM5GawDdRdAf0vgwHtccyE
f1EepQ6cUlTt1b0RvlGRixqPnCF4xJ9TdfzTCIa3yp5dtI4P96/5HoXYfvz39/OsrO7GdTTT2n8m
79WwQYy91rSUn/3YvE4dCyZITpQL89RkXpZQM/pLSORkN/SYvUpJlC524yhFvZEBkAWrxj7d+ztu
wxwDKSl2Wl1vkAw9AtC8wBAHbJEoxg/gZcfmHJ1ds4ysDrUseKBrwKMKbGxhn+ebHTDZrq1Y/JkX
mPLj+FyeSG7hME04t5FwEdn8ync/91ePA1w56odFWadQtFJGNs5m0URmOiWgPCYawEy1Mo67Ld8X
cMbk+wKJxhCyd3lpNLiO87fF8FCp6QmH7W2SzH2ys42Gqt36Ur/NB0FrZtQZvIyq/DssHwtMPM79
LEHPmueroh76TGqZHOFNQzdFOpDW11GUQZRAERIXT5CaKxTnJUz/ffzm+WQtyC6FVih0kANs/+oz
tUP5iQONKNBjX5uqf9jIN31bntxdLxTJ1W5qgDEmVYhdMqfCeEyLpBnW0vykGxb/TgL+A6Yjkqii
N/OurWwqOEBKxSKpimAph9RC72l2FW3OuaG86jHtT6ga+Eh0VHVpnnolMAu30UKheGgx8hqoRRML
B8RD+blezqifQnxpGZ3q+tcy34gOAjWWMb5kdDz95JhlcMq9Qq6OgfW2ONMOZaOJj7qLN/qm5ExA
xB3SSUNseFXUMmJK1JjBwg+4/SbibrOKTrZ7hh755cTC4gKQQKi9ig2/9sBjrRtaKxUEilqeI+60
6bbSDfRXLoVoNV90KfOUnRNRGoqHrxgOWhVFwGJPDMt6t27PimnB/olIpeSJcX+DxFjERAuIItjx
WTFfXiURYUtMv/B6Whr4LCkeJQRmNIsEv6UbbN/XuyxjApc8R6IyiP4jeMHpJfqk/oDUukioVg1x
pS2alA5V9pr32R6hEy0BemRcKrvjfCffiIUPzpoT45SV1cAIlBKiVd03Sc4KNj648gaq2BMPqYdX
17lC9wlKcQmiA13kZZ8gWheUSeyL5DS18rHAhCFGYSh183C2/9fPwpcdftUCS6tY2mFVrufHCRsZ
dIYABuvVg83FRnmaCF3EfHyGJJVpaEMAq+/hg2mSfhomP00Zz9hScLtJ6/mGZu5Isj6cadNI3Hz4
3k96qap6z68+mIV2NXoIcEshWFwwMpu+F9WOxdo4xnb83uzoxQvtCvzC6i/QLKamJqm+iyda3++N
MXUbXXU+fGD/YIgtgsjq9hsbeXmB/Mr0sUeMy8wlPADj5swKudi4p+jMOKFlcMIj12xdb4X1Ywz+
0o3mo+WITAOFwZZMC2iBDYGJ6ZdR1PGPVy7x7fRemMFs5J8if7bfzRwGmiD3XpG+2amULyCyIFr6
f+5Ac4tOOIoGSPyvVJ214gSfpQyKk1sV3jiHFsacvrvQHGZTYD1HffWXbN4J8hMoM+OErDvyYgxv
pE6qxnNT7/l7OTub9J2jD/knDjN7qUY3hAoWytG1VC70pBTneIRNfr9UFsCbM3R30PsKyS67XcFc
eygj6So6YTQ6Ov9IGv2/cZT21u5uFq99+kiNsrxYkbZtCTKX/dMbkUDpn+fU9bxtRj2oUPb3lvfq
L4vcnoHL8m32IDg+F16xMIrKAkPq2CKpAKP0u5t+yLjb1KY5gTD1ETmf3vkkVXHg3FC3zzBAGQ30
B8N/XCSIdZ+Kvh8ghQ0uJQaAbWn4kej8fONWvbLI1C+q3b4Gd2RG8aI79KG5CMwxSQwb/ukPfvfl
n4X0GaBt9l6UKSabuYAUAuxmM5xf/AqC0QnCe+6hZLXOz/EVs4wAoQHdatMo52KzIh1D6cf+BSBZ
axu1WVzIyGj2PfgkOEkf4EtMZHQZg+lEdk2xDzNNHPeOaQbeTMJvUx8EFc5z2MCYRYbaKAhNFqil
kMkQ56lvs0Slgt7bzZIgUBgTES15WqnxwOId3Ce2RomRWZ9ONC7Xg1SK+EG9P1hJENIOAiE5JrZ9
+eKuNPEtFKMa4c3fd2AO/cC5AoRpCou6tjA9zMC/h2XtRHMsDNj/+2PsHdZR4nY8XPdf0WQ/wUuk
Mky5brfMc9Ey7GaXamGiFqkbwJNPW+UaLVDkGrIX3wZCRqeAigtBfUuje7CbRd4ky94Xiw3PNXqZ
WvEwsDlUy1gpyPedD1Hhrd0WaFvUCCc/Cdcyx3gNHxvN8IwSmD7UCjKbLgWG7cZrrfhUw068X3Sk
1PrsQEVysKRSn9JRZRSYk0yTZnOlZi6xxzZd2w3jv5n8zVUW38rt1nsoIIzsmiadeSQiaYsw1ZE7
x8qa8y4UobSEztqPssq4Q2pZ1T5iLa9PFO9xh5EJiEzaExTxCAwhZstK8TBERLyVPe2TNfqlmhCY
ZESbml42bXApJtSEBL62zDY7NtT+xforXbXmIvr/Lia2KiDPWKt/+2KohLFfn7Nzyo6UbIJyEdb6
b2f1S0LbEiuHiKuAO1RENHdiZYmlIIVvpyFz3HKN3nR12vfbo+8KtMaCXfP94srXtZdhHSCalKuM
cnA0Bnxcu9OXvKE5qTPVPRZ3fZzgElTs/YmbLl7MlTibD79tDnPwlUKsupiWry++n3hmZ56Tx5GJ
ADDqVSZzndddWxKvvQVyyx7NITZB4SmXoB7HLLf5+o/77Rb9IZCfsuTukV0OJmypESjy82HvHCCM
pC8omPvNw/oNQWjtYS7GIYIz6H3m4lkm1TVVqyOAVpOQv7yVSni6ENowXmwVBfSyYMSpHg2fLiWA
eP+xNBYd/N/EX2w52a0GRsQ3KQTzv5lV1clge8roaxZiIzXKhtD5haOZTXEnAX6IMoXdKEbBarYf
TnV+GAg5Wj3fEoUp1Vm5K5BrYuqxUlMaG6SnG6D+vspuig5XIiyFUdQcZ6ttmvCKs22GFhAwYOV2
+YKsLpnnmxE+NBtyfu55EK8RNOetIIWl4VqFcu+BUF8OnYbR+mb84rcOdnMcfifYsB/MVLcXQpl9
xe0tAyxsGJBvBcutGylBd3JmwJ7zZi4EdVK57IY33GQNhOR4uNka0NSmEsCqMFqijKJe4pa8cgWX
X1IJN5OTigIgCFT5fQ/ackiB/CU2su/PAkhRfXsKCbquKGDw/M9wX53cXO3MwMO3gU87S5xJcbvJ
QHchxEXgFcDqeo7VdI0rX2QJxc1eaO+/ZdLXQ9Q6i8dtLpOS3bl9/Q6j/imGXpnhccAD+l+gSTIH
ORwbtAA72PiiHqWVifW8P9smeTlto/1iE6SpkzkN4k5UR9waWn5ikBXep8uiVkLPVjJvsylp4uYI
JlNjiBKD+wDPvkKt5VKYFEJLYxa6uORAq6ZTE8VbqLe9ZZF4jx3gO5nU+g/eWHgS4DJxzObLbpUR
AJfsA03Cqyw98GQpBIsl7RArqDRTD9CiG5lIWa/JTqU2zQxTaqq9VKrLhSplWZiRAeEAbMvnA/xH
/Az0t+rREyCY8KjMx/fG22MUuTVQnllUFl8HonZvEV33gEdzxDjiaLnSYJn1M65QBVMDqyzVqoFP
Hhu+0PgENVxu72WdK56uu9KQUgr6tWaQVyHzNbf9vKum3Hyk1NYv/Nj/g9MQGqeS3UnbKqZg5tHC
CwH7O3n3dvXPNGnu4XfUy8FUIXrPin84SX7JjN/GbFGrmd/8e81QsLi2qjDBrO6YPpKakEsEsH1W
m2Vd3PBpNavp734C/u4YJqs0fGGfz/SUFBlw44GcqzygIvvN/NMkLm1Bo44dLULtdyXxchn5mn7A
pw2WfarMYRJfQtWQ4eTgfztK8u2BgoqlGSA6Jh3vb9StMb10QRGDSNaaCZ5X3wsUYMd/eCsBe4TB
YTAd3VsBJweT08cDPV8IIlqSjp+yzt49md4kufeZGnD/etUAN22PGzLAdmSu0KZu1hDlWJ8OvrqW
eSnJjFvKD3FLzhhdr6Xu5fJ5f/M7oRLWvKXhvDaNb2wdQk2wWw2kPmhkX91t18F7b8a+L6FGkJUr
AGwII7vpRxBYc4M5Z6Qn0avxrswsZIAGq2jTWlhFQO8kb9e4ZgWkPosjoMy4cUPvQGPCw89JmoLO
VgojoQ+FQcIdVe/pOA2SjAJFWjkUJnfgkfwnEfsIEvmNjAg9YaSFPw2GYjobClwWbDm2v4LZ1G5M
BNKr7dHg62aKXNoNaG5H4wkv+7P11ivCLWz5ZfIC6CDuVjcIn5KztVixGciGsULu0hXpe3Unx7Mf
oiqSQVR+AMtmLDWOFFuAy0m01dnv+50Pcy6zbwL0oZFR+Dqkh4IhPRrucCiDnEFb8JupCJVYM7D8
fAWFDfrMczUqyuHgiyafeKlymqG3R2BQr33zS5uk83L/iryYeRzmo8SHTCEX9cV44kfZycszmP/K
LSIodFo7wKtw/s4tO/fX2peJMtlenV5DhRIRGH6uzFAc5GAfQLDvozw/9FPPOu7hQk0C+u1De7J2
uUUWYwZQ+UcbL0RBPlqjo4DvNtz+Ak/cV59J0TRQaqNG5qac+kIrlpzJBLQJUfYzE5kegoSJQfxp
3Go8bl0Iuw/re3L68bdYXy5GacQVPrwqBWGGAqmEvKMNUwEpqp28DFE3kZSFvDVQXVF8y8o/Pkdv
gMPnTOwAHVDtnyFYQ8OxiXw3QUd4sUhIeGKLhNiJ7VTVBurkwQtTghlAWx388zxCGBaSi4RO9dWG
J3Dvw1an5shib3zS60xJblcP+5pNTQXyA09OZvilLJUQHBBVb511OJocmNZ/X2KB9hTVh1YuHpNY
HgXzuS08XgnOh3rd1+jyzylUl430yywpLlhZwQx96zjUUXH4cCwCQr9oxIaInmuE5QNAyAr6p4hE
1LrCtvoNkrpDCYqI6KkwrNC19vxts2EkqUCQXB0cHOSEkAyr++L7DjwZrchgb/LfhUVnSs698DeL
EDZmaQzjYFq5t0bAmXaWWiTczrO81vwKNb+JWpmPSjPsgzvzzBrSaRQBUHjHak1HpaDrPX6QSJov
gerE/Bdp4TOJcKYrBwlT16ji33DYT/+M9unJEWkpE3Sy+8lFcKB+Lfxq0FR5rCtWPrbuUX0gq3ri
IjyFO4QzvMYexrZBpLji7+qyfZaDTpHHDEmVRV1OSSmBDsezl12ATFdoHPiac4j4N1dCLcj1Mvkb
W19SZELKoFjr9XoZihxwIjNo1Z4gpFiGko6BN1Tbb898eCOB5G9k6UYC10mnLXZCl5ffPa9YM6RB
k4of+A4jfHkrI0+mKKn1qu7l8gWz6ipWiZmNuyDaE3PmdsY4Esct/2f0V6wFz2ke5yhrj56ghK1u
kvPODlaiJo0TAcoK+Lr386HSMe9nlUp3ifex0Ji5lFYOpkYJWuaUbNHftmPgrSZEN/M71X70XiuU
TH5REc3FgI/CRzCOBb3YVdXgqvc7vZnVzwdwPqVH/g2Yn3hQ3d4S5KXO8tHFtaBXhrsz9g23NrBy
M1tZ0K9hNosMIZIm4Fg4TZs9QH9MG2VhF+lsUZOqBBn4/ascfh/ySDursuXqsO3FL7WbQQIjB2cG
aMLbNhlwDvLTi41SK2oG1/QUxcVQK3B9/7z+RRSzT6NS/qzxqRWYU08n1m+enLsX/uiinUWzXN6C
xBZvbAgvIySmjyJTK1oZ/2fDzDxX5OxjeuqzqNV3v4Uh4F90VJsfBOkGv7JI+Q8Mua80pNo2dLKy
b06RTgUD2YVZkQ4Ba7NxW2qFgRyMF81myr7QNYpybZoFGtxuoFFesxYMWfSa99E1PP3K36jupsSr
kvcj+tDTuwZqHKY7AucgHkCs/6ZqIuwsFdoGbh7ulCm5Pp9aE3rVKliZBjir4dOav1jA+A+L7qvn
2oZUaKmbjYU8aIfQVbrB6A9ma2hFSYsAOsSoxl0eLOnzxFvxgU7hV3EGPS/UFl+MOZd4fQ+GS9V/
tgbXO0TjCmRisepa2j9BcCXScdVaJgcWH2IMsSMoodwe9tm73xpOa1LfUjCjDA572o2AcyBk3Btq
c05vg549iyvxC0t5LGZMEOljyB073/3CQlwEJAN9gYf9TCLqi3NtgfYuR8rUvNZCOANq55rkEHpF
0Uzf1M1lwAja5mUEsHYuGQwiVLkP1I+C39C92irfSWdqYbimEWbO1pEW9NvOPxtkmPZjMJp6orPg
nVaC/y42+gcUA2Z/UHL12CFkjYJp+LNpIn0cTH2mhnuUsszU4wUwJeXF4Zywm11WN0R1Jmo5BSF2
wdd1XYdKWg+ujcno0X2wyW+B2d0MwXNoPi7tj3UmUYkxNSk10DI5nAFQQhS29eZBAxzKR6fZFPG0
lnIfOP/F+YhjJKFe2FNiNv8BQAkW8rvLFW7yN63aT7mbDFqVS2PX5k419HwTOTit8Q1CqrACVfGY
BsXnGp4sKm4sVr8IP35bZTG4mkcg1m48as5Iim53NlRbdgjQJixpNNbk9ISXwbRrUSe2UI6ttDFA
c6VsmxaWyVQmBQmClvw0WaZ3CIgwMLaFbpkTYIzrPwb+9cKUNKouumtTreqkmidVCGlgLfJW2O/n
B4xWs/23W6ts/OmRK9L1PKoVTM4EhYriQ9EmN8u1K42PTPQ2giTegmBlwy7xK9fg7PlBERmP8+w1
pfbcD0W5NQeUsWqYO+RM2zo1RKn+X88549fXH5IZsjQZ69dSSE20LozYiYZVKIReHVUKi6GItVEq
HukYOORBI7+zziJtc1sNCY8MzU2yY17JZ88h48ehLDmLZt9ETXvWw9fFDkBwnD7xcq9Y4XPnvtyA
6zRU/GdENomaKkaKOblsJT7Eqz98ZtXxP6t8FvJ6pIsVQdPoK6kJc0CaH5y/MoGoOHn+PTygYb35
b9kAGFJ5G4fiHx7aG26pNl+pPhi9/j2bKmjuoqQz2qrwVDIQWcuWul1lMog2fEAs3Wqh7VmBaAbv
K4ENc7WF44/J9FmmjybMoLbWE625h7357uxkZKOfRPgRqWxOkE7+Cc5qIV7hD17lc1jeff4GS4QD
d7zUyGAtbqE/rzilzppGKqKeAQ/1Ih4iEu4x9er99sWUNGwfIrdccBmH+YE2wkGCLfUq/cKK+uUj
oa7PlxO28YOQfr9OeS5/+BsnILOD2Xm8fBbaYdpRlYZG33to3lP4Ul2XFv0uQfUhYWi3cZSrbTH9
xhIVJCuA2AYh61QjDjTbT6Rwmth+kXc+0KbJftLZjDaefJZ28dhPNOZOykXtrUEGFAHysvD9T3c0
WxIl5otp7hgZIvB+G6rv8n/XfFrlo4Qa5cghlc05hw2Od0ChMKIDATlohLvs2t9tru0DYnGL7NcM
HnRSfCeqt1o9OvHGuxkolNsTRrBEDFQn1GJNE3U70sMAbSr4h8acE5FV4vv+/NItHwaVJ7ezblBf
L1PC6gMxVKARCaSNBAbL8fnO9hLTZCF37knurgI/SVZakS5fs8744Hwzq66UHX8Kxvz4ORtxxaHR
uTCA61L6uhVLfTUms+VCi9Q4HrwKGD34MzbVUduh8ypXV7RV0yrXigpmdnr3DZtX5vZxudJRO8Q6
CvMGLLjlU3FLnlbYmtl9ZZtNFq5oAT7Lu7FN5VFjtGjvEVgMdyUz434CzY9h/1IwLlL99MZwHs0q
XogWJVfIaIcVHJJAm5Kg09odvVgKEJTrqL7FqI5aM88VkLxMs6D4WWuUcXiVpfexuyb+Vcft1eNF
Y4D8pFZJGGSjfUKsCk6ePzC4UKTKJI7WBdeCapS8v9edMxznSzBqwdov6WZv7waMIDEw+Bu9y3sP
bX+sKx3wdcnEMycr3+nIajWuLgMnno3ECVl7nV/hnYgReZ+0BrFrC7GuTtJSJA60rrkooY+xGPNw
1n4BJnvpA2PqcdgpcuTkqVlYlfYDQZu1s70NgHBzM/Mi84GMgZZ4/AYmHc0LePQTBQKXKvLCwl5R
r3ooQ6Et24Y/Peg3WdQe5C3YR1WMjeV6w5YFDFGyCGSlw9ix5et4Djy4fMIIabwMm+qqTrYwcscH
2pfs/uxl8IogKRA4PkMtOtuP6K9MQWjTVM5MclB27u5UmjObmPFqa+YaLZkGKvl/yz88uvH7uVQk
F5Q0bK3Kpv3cEDyqXRNHPqYFVAhezoDrYaINSgJ82E/+aalSIc1F91DoHLSrF7MgTZG45+9yZDeo
jd6hEGpnu2G4S4VGLrhK1kDUPQU/6QG4+NsdUMvfq4zsmhqHz6J69LVaaSVlVf+taDFqKelEzXp8
+7BLs1n0XSN7MBqsu8lPw273UAJuCg9aRqt3IbTzf/+1OuvhbSYdh1OZkbHnEWuMEJw+e+y5h+wJ
g/zFSAtzK8rbD1L1ufR4yyTo1X5fe9owgc/7HALOyphecd5IeNrHptrToklPP7srZd7tAp1ld3+o
v7VU8powu90EbEnUWhS5L6SbFi/2WNASUYrPUB0VU4EYjPzYzNTLj9SBAuB0u9boBVt0Cq1jYlSl
jfMadn2W020ZNiWniL44d9Cmict8ud3vjbN08ONnLvLvKXogdf8P7JtkofpXarvY++hQ+AM7lMqu
7FoM1AKkg4+quXsuotHQFNjBvXHnvBWYlEe0vbc1RbNki87YNvcpXz/XhjMd3ymeZaRuLWEUFgCS
no07F6NpR4ypSOKkHK22xt1E0xJWhnhbZ2iBeIpnZCbJjocct1pvV/RJk5Y/Lfly35U5lLLRDJRi
+TMd6skuR2+eNpyHBUaNiDvVcz8my+FQBZGeQiC3YSBYHsuAFlo3p2q17jWb3Lac0JZPlqqDprsw
MjVkWwuxADeMOCXEgf77h2VdTKZheGu/Msz+xx+cbdSEr0Izho1eXxhbl8LSSOU8eINBCO0YSX2z
h+aRQbLCm6+IUN/N+uMpBR63y8K47Uzbn5tQP6HC25fkjKzzZkRH30sYAYCk0UpMxmVuennLv8wG
lsVUJ4phd4FavKi68WocX0I6aSV/10mM1nwMpSbKa0G1FkxQo3MmdBs3IPKabU22nzEUfP96KE7g
XkeLrXXLdK6MH0oAW+a/sJC+xiMEelzrjVI7vBbLW4nu0LuvDPJoRLM9krvTD5lZ4af4Ll78oeNl
kwQgjSAXJB7l7ikr9bs4SG4F2wxyTGLcOwJWpvjgLXX0JkxX7MhWkZP2MirqYVT0RtkglAdM9UfK
mlqBf+1OsNOobUiHjsY6tzVJxEvZrb9/jflJdcqmkmzwdJB3BL1T858hwlPcTAOl32/LbQ7YE7Kt
l9AnmN8fsrVfb8fPThzA9tDIlblbuLUBL1Xm/CtpLwQ8aDu6MPJyL7WK37VPWWKAvLmoOvRUPnxX
l6ndeFSLKQ3LvDRK5/o14Ok5eirdIpExYwIlSslihY8QyuFe7o92bOG4yQ43oxotvcl1wFEchmQ3
L0Ko7A/2n2/5WqnviLdpp/7etumJpt+cxtaWxqxOWaQDT8s4ENB0ipBsLf3VdHBhNd2Bs/iHVJuU
92Kjt/+w3gC2NgPmnzDbwoH6bYNZe/5sH724+wOzivd4WaHN2g7aKRdIm7GcT0bhhQOUbDO87P14
7aV57iXeu1GTQY8tCyGqILXrGhFO4nfGrCDo8/l6oCVRvaX3qG1ohdK86FSiadT4PyxvwxDJrz8k
BUVAcaGPi6bnofeoiY4WZ9u623JJAkWlUuE4y4NxUnharjeH771qd7muC3Tui5MtMopJuMVsS8hT
xxkW+eqLUGiRbqi5vjKbqkvCkmZYnjcM6tqvRQR19iKoD3U2X9EtoavnnupoW3WWCoEZZ7qOFQyy
45qwAzqKmqOSj0dbQGgip5lOhLHcl0hApjUv22snstYSjUauKWbLHAoBIUmXhoKFL5/sBbJHKAbL
EDLQDgtvnbRVZfPAdE4q0wNw8OkCYc5o3LRbhMN/tlBhNNx1YOFNeMa3Rq8RKZQXxW3glPJpw1Zi
NO0aEfdpHs3qS0iHlYEOj8umA7abBIXhAVFwT9w6HH2J5luPB3msPWe8oHOfGvfuzy8d4BOt93os
6Md+B7sLl5HdNZgnKmUYecYFN6rP4V6PwST0XcK0+PfYc3tpU2N/IMDUEK2pdrPqn7j9kxA96i1M
7DUTs5isJ8H1tO5J6CJTRunNV6IbrAN0nCYCkrgip9ofK7tO4GORpz30AE6wHlhQUbHzsvlQksqz
4RnZzVvGk/1IN0xW/qX1zLYEd+nj5ooQrIIK6ydL9x67IWplQ3MPDX4kfmlfEorTQ/35xOUVNdi2
Ex84A9UEF2BFMaF+/k0dfkLy4Xaln6HNLezBrfVB8IEgiSjdNdOgP06Idj3K/L2mbBeQcog9NoAb
Eh+2HGQQ1GXXSb1ynmMdZm+QNH0o+me36CxnFTyRkaipuj/0q3cLrz4xTrFzD9GfEf/xpD01mBnD
AyOshMd+4z6Mc5BOC1D14h+J+mDCXT1dPIVlRu2KbEbkcEMgAfN/Ig38yA15jsEnP1dyhL5KRqc2
9bsJKghsLOUcq3EWfrsuoYOswDo6OFnjwcZyhcBpqZYGQ4dqDSF7obRz+18STeXtnNh/v+4ion1C
PjGg86OcGuPpbg9CmVZUuorZ9w3h9NprdhEhxCTquzxkL5JglW2v5nt8omq7dXMSn101dgPwwY0S
nDXeZ18MVOsJ+d/pUow7JUooP2dnCfRnTIYKYYu7TI+34nhFeB8Uz5kUhk/UDUuq8ycXXTnuVE07
ybTZzfA4pD/tQ56R/OxJsIcZuZ5Nf+IiWo86pbkKCPnHYFG92RAtnKZmrcG2k/Ib2SqvbXNJ/JbA
aU4KYinM5ycsEcncLmPqfBawph3Fk7H0MF2CQ3C+hjdexpp5oBF/JYELj8B+DoFtlnFu5PmIT0mx
pTDBvAtF8N0Zy8w8dBuMURCWWvmz3rfOzRAvVeXHjcI/WZ3ecy7Z5I3tZQkDIQXRl7btzMiiBt8D
8tRgg/p0ykZs8BIOEAwPVQa9ZUodAezCcPyM+EypssTovxXEr3XZXFHDfyDSShXJkPJnHTVUhqcA
SEtiBqY2a9r1ABKWnYfHRSfh6XCumIJeKFPKphqV8pehBhhOa6GKnSJprXKnq0oTQcWwH38yeiPg
SfAMA0T7ATdT38E9Gv5L4/5Htq+AXPi2nwxVD02kFa/vaez2gV6tveq6u7ERiqk42HdvAN6XoPL2
Z+gqeAU4v6iuVOnV+4CLS/2Dh95R4dGhAKzXj4rMqEu1qTRtWjdxJgQ/uYrXw36OW+ARjSKKzhC3
pIQ4Pyz+viEvLfrXqVyONJ6iYDj5jBONfAwY/uZJXFlf1aRLhHEwkeSYPnICseDTxkLxPhzXeeKB
BKdr/dZ3J9IjEGk8QQl17VmcooE9JKsFIICrQYfZ/SPPmaUMjINfGgvOmiQV3vbE4r2v/55N+y8W
mMkSuE1Yn7tncI6B2sxBpq6NQ+BnbFfrcj9FOLVNXdOVvABJmxK3JfMJGiT/tZQmeRhdjewupV3k
d5a+obzd8eswnyYGu/fNjBUFCmeA6SVc91GZU5QZmRACJ8+3B6qrNGhT/Wpa/uKv4G4aqZOKQ9bV
iMilRrfnkNNI7yGKXb0jLTqNOTpLYrIxf90tXzkf0LT6Xm3N7gbimd4VcAc3ZN1o3PXJBKlE4iWh
Jfqclu27wASW27yKyAN45IDVhRXvZTb8D0K1mTz5+GOFLznRaylcLDSygmnhuo5nRZ948HApmFCj
Eo1XDxMxAYcjltaBi8KiOKQWIutZTD2CAogDC5GSIEaAeF5D5gnPgaDCXBgQomeptn3YePqTzKmJ
L2zwr5cQeRegsigstBzhLHCORMGOQeaUUojydMIPsyWiqRblzrZ0IjO3i6TwjeHcNJ4wCYhK6jdA
8AEvdmZUgfZISwNtuQ+U0rBFCPhX1U31EYRUBKQX7Sui6TARjCjTAcVW392a5DwGirImX5wPEcDg
w2WonF93QVh9dXe0rZjJEG4mPNeatlPmCl13bUZmHk0RZJaWGczbV+oFuqN1uqm0dw6ZrJLFcXA3
2TqySl8N9dk0vFz5b9uaAtMQCxgzxSbqm8f01Mpcln/ewBuVhjls1N2vMimkVoTsShwpGx3H5Zcm
h/JZdjvnSNtWh3vwMDo7FfoUOCpK6NbNGgMjD8IS9Ec88A74XM15RM3cH4LevKc8DO4C+eTyWas6
4xaeTCeSNQqcdwkDuJOSwvkZ8ecroBc+sX9DmzEHYNwrPVER5PGN94Q6fPs6W3Ean7aPOds2cm1k
Cju6BqvrLDgkZmyppXDvCGxyHoG47ilFdzDUF7sOk5Hr6ps6BP83e5kudTLZEsPN7TWrrFvj952Q
yU0xCR7Biei0fv+a3dVy+MLXysUfbMMzF8tQxgFMXjXDyjcZTxC/WyfVVjjkagKzbHJ4Tr5qY5wF
xpPdEDTLnzH0h+gP8gG6Ge7bRC6NpG/pTXyl1eUgaEQjBREdXjBMNAeO+ET01xpm0uvQzF/6hNK/
HVEJ/Fx+WWgQ/mLEjSZ+BFQ5nnWIN2u7PB0hUAJgFQ1nUrM/KZF9R0j9RGGCJZCTd3BZtcjVaQrQ
nlO8UMxqW1qA+30dc0KLoZeatPrGBJ0+qlKGUD57kIaOfHScBWBVKqn5m/lXOllN9FT36VaJtYBE
aOGH/cNJPZ+TbYkoukJQLzzv3UA09GDQMjqYl+rv9fKXg4iipSUGax6+S/ralkdn9AkV1HcU9uQa
QRpglegkyVA47kRAr15j/YtAZDmu2Ts0/66yI4/DYh5rqtvOhOWwmoHbeUwua5OI1+XbXYf/itfX
UsStaRmyuE3jRAAp7Tut16v/HsF1rJ317Qmr0Ev7gkjJaOsVgJ6RRJo+U7trGBkj/RZQ8mkcSguQ
jk34ioIkD73ycpQaRe2Xgc//kl8m7dz2o4gi8QsWfoMk3RQJCJWxEBCvfb3QTXTY2aMQPEl2yWVL
Up0TxwN/OxTYHHyLyz69ozCSuoHRDKg6HYiw9qstjA9QZinUZ+Z+uTtKjCbqZUN6j7VmfH/a2WAT
mOFuegc+suMuZmCMDsw//dbUYQg23VG+6X2h4eboHIrpr3aTDanXUh+GrsdTP4o1yBKatwmh3vVP
5YPAidk9cegU5THLzFlJSClkqOopMX09d6uIZfr9VnJNf/zqUeftmQgLtgxYbaVUdf0QW3B/Dn9J
Jlx1rUc2rBZabE5C/IZYHMbeOQfnV/2Za/5uNbScXHgHzvKEkPUVjKLweP5lMY8cGqcRtwhDLeLn
zoXZEXSqe2XgCy1w7JePkoibpZCFTSUvkiY/oaC37Om+mUqtGXu1aNMb1TOgVf9wkvmiGzjTXwyq
aq0iQbj79DfC2yr5m5O6eVLeJ3ohAtLQ9rhSMSS37vhsgFNTMPQiZ1AYzhwEym2aQ9wovFbDuPle
SVJbYEu58Z4qm73MHmSfewG66yI5IyC12FUCPu5HM87wL0C4kngQ/i+J3gTFN1jTvJWm/SHLPzW2
/2IyeFVvGS1Jkz3SzaMiJIy1SD4Zckzbf+X+rZp37nNUcZVphOyL7iRI7Qm3pstRumuQBY2u2VdQ
3Dj3OZsEsoWIG/MUYwX6gk79qVySOYjhCh+Qp5iBWCahww6/naq4HvH6oXjB6boEAj0zOM4xGsFJ
r7MMZp6cKUg3787Fjul1mZBzBiR8Z+5b241A7dgFm8gucNWU8RiGn+EZOVLpot0rpleVZDnFwrOQ
DIaF9ZH6yT4Y/4KJsAM+yQ6xiZWDne8aHq7tW4ak5QPhL/QPVPz18YPrHjhM5E0lOj5jHm1lq3xg
yHyiwASXkatPDU2BBiYyHLgCW88LN4E8npjeUyFwvecgXng48PTyTs7zIPjXL275iUP7ALa6PEdG
JcAVwQgjFTTUCf12eRhCeIrigk4pR2ZuV3wnBGNtE7GUUozq9B63bnS2pVaPomEWT/gv7+6CJA8D
RjtkC/jwE4i/Z8TH2EuPPacH47xEUg691RPzw152/WOe7sx6Mn/KN+nXArbrCawnlp2jcT6f1BIC
8/HOYggVq7U8wRtW0b8KLX5BUAUU8flaOuJDHFSHznsuc1/0UwiCN9Mpswd1+3o2kux8O+/6fDIk
07bgpz10IPWaEyLWqhQtnATF2kDgEuKc2R0+IeNFk2O55397G2vVuTLTQi0JbrkVWfoYJQkVLi+M
/uhVXdO/fLgqDQO+1OWNCWMuXwbGw0n1k1t4NkqrSaR2h/dUR3sN7+FT1NCX+pWtExwLklt5pVTt
NDchDGLW9PNjGmoPSVG1Maw5ORm/bf6WCqrsU1aRN/p7m1NJFvARujJbaiPtNiRLTfr0agHfnfP5
1Xz8IBK95u8b6UrbwwHKKWIJ/K1vNhWr6UG5dTxSzerqthiq6JPr00ZOFsAtC92cUccZrnEEHsgd
9uTHqQEZJuC9cOpmg1HDI7M/NWhJXFtM1rWii9mUatGMi35e8bkT+vbWxAUwIbxfjt/7BRpeyxNA
5rxr3jRzG6KV0Oxq8/WnsGfmLZwYQhqn9CPpXWKXWwD7AgGl6iHrWs1VbjYPp3tcW4fU/1ToVK22
kxz2PBN0sktLezU3Lhxgr7Igz96zTIYUXKykCQdZfgJNy/Kwo6DzEushRdq2yEHbF824gS5R2RN9
CSUSaeVedpagBLFMkRmpu/u6Szxgael4NPG+HiOhOxtC4m3QvkH6I/OHoFIXXiZhhG0b10DkMaP6
KS4ItU31frmLPVYZVMbLjjZQ62A3U9JMBtk/Ss4iE/EbJRTQ8Ny/7SL5jmJxLcFdO/hbQXFaSvxX
ynSCApzZ2dIV9059oTk8r7IqIvBn8MLZrv+5nXRMNrkp/IgkHPHRr88/WSHsbu16M0ahhsjWmP/S
ZAwmLudUc77dB5D75wovE77fLrvGpgYdAJQgdyO/4FoYs3OHmAJwFRud5dmxulXeOuP0SVRkxyAI
QIoYNV+F9292biIvNHTEjDGG5hMawiWlA39S7ibtO6qfj1PDc0OSn9HPxb1pAuYxnHSeNtDeO4+6
UeNcd776LEfjfb1693bhOE7YhHszKGqD2QTlZpeFlkq2hyc7xygJ5te5LVd/LeRHwv7CgSvbqJ9W
dU3LwngLOn6oYAX2tusX3NBGImH9GK+1zje7E8Vcidj58HRKFYIR2/b5/9EsWX461CG3h68XloW3
VWTEAfeCGewc7Cl6U+KTK9k7a56nBRzbT57gvZ8K1ZPo05NXVJQwv3htYCm2tAkMPNSeViEqjkK5
v0L671e2TrqFIYtXbpbZRZZS8/+Bk/g9yxKAQgMnEOQuJUobSlx1KZOMo6xQwftpHUifADytr/Jq
/DUKzU+XjRBxlFUsVpT4QI3nuBucJFlRICOflmYKLPZkK8WWWxFWqIPxFhGLWbbhbZki9Uq6lHlJ
zLvquCbKDd2iH1LtZVbY/aZdvVhZ/XImwu2+5r+OYy0+f69L76gzBbcYrCaM/TIyf1CGxAWlb0jw
zg7jg4d6Xu3IcW4tI45lWQ78wGtl7rs8pcFIEdH02p7LHB2mZ/3TWfCoOHFUuea6pSsfYQIgUzf+
8tCS/Usk5PYcD53jqY3WP2qyRloW8HCpSTZQ2IrH50RNcUUkm0dhtRbF5z2baY1xmIyHx/NWA7Fq
qGG628tsP87z8QeQ0j5R6eHWnLYWQzdDyMJcDCc6DoixVfBb/lfzYvs+L5QlTiIgilBba3nBqru3
UmBz+RahmLj6bLn4VrKuLyGLxEDmXnj0d/H9FK+KAXUkIYu5DzLXgp2DvzmyuK5aLLOtsS4p7nCb
2Li3WYFUyjR7EAsc3Wir3tDCVZN725w9hw29t9yRBBZ6wS6YqKg38i3R7tsg3DswEl9M+GSqN57d
xAxy0CLv9ujboYznWJGsBmXBpyVC2kKbxd6/wnOXeoNQj3E7FOYys04C6hABy6zQgT66HvHliTaa
fz5dZIjzj0cbZM44EWGOX4lYkBa2LA7obuPHCbN5Z6eLs9vF++qcPdeTZ3groFKNpFPNP2Wfk4cS
n3kaDMrHz10K8VI0wyz0xyBdXRTcpY4N2xziwgjwtPVV/Qb1zVAZJNxNPgxA5J2gZ1bfcU+Mg2lN
mj2lU1gOdl0BtPKDgK0VXJh1lNy4jvwmdb+GntRlVR8JSqwHoFrIJUu2cI62NbVt0E7D57uE3/7j
9yMLiJ5zJhOKIY737HwdSjXoCbXUkJeV2r2dfa2PCcVReUZc7/sHodFrjcava6xHUYZWbqhpzjJ8
6cgXnkvGHHJM35KFpzZYxy6YB0wgXnjL3Jrl0W27iHPyEHWg/oYTirm+iMASsLMUzGo57oOa5nf/
2etu4Oat0VyZSd4UmINYZbNxXcKTONQyw38qDED1GYxSzaARyj+127M69zkc47+bzdQY/mPdhZ+5
UNSWveDKh51uKw/m0DkthZBnuGAGjs7E4lOTEaCELr+3WxTtNE7gbfB7dK8JRyuC5B53zOhMPtv6
NMFf5tvx2gOxiNjZThkAWg4ZB5N+M8illXf+9mSuKmYY6n0bU4llyYevJOOkFDY2P06ehjLHxdCG
K6PsudCBvSc59Tq9jRnc8npXsKVgLPdo13w9OTOGlZJxOegCBQl9JAMdUerzRcSGL2XOIXs9P/WC
o/UOaWnpZapRVdN+7yIX1wDgoKLeem4tW3oRJ9QEbKuWO84BnyGccy9FpAcX8etlNYighBerH1G9
9lkA/gGHZk2+zEhJ7GJUVGOq3C07A8if2AUjlFG9aC4hDTrpG9sbUVZCJ6eP2YW+rjx8iIdVjvng
r8WyHLll3CT+ligycvUHeMALXeVjXqerGIH26pD7s+LsL9s6MMK8kwWvnixIe/IdhYNpH0ySA1AU
D4xjM8LAop9EQR2vnruNpO83iULAtAysoeNzwkkp1J8u6LSczZBE6/wP+3eq1UWVEI0oRbS2VGue
K6lRVa3uV0dQZX+z3WadCYGqGHioLyJ+0uXvlV0iJzaJ2Qw1saC8kaApL0+bo5hY4UxP+w9H71rB
j9wfYYln5krb+BHTb4xso0uYlzeSi9dASS7wiX2XgKb9JDGQGvE8CNa7DJqL+uVeTRwnZg+ktn4C
jGuFIv8QWYAmYTsp036urm8iqKNih7H/xOxfVPgueyx79sfUNAtvyurCq3QMtFepKsr6yiIikK8G
1zNQn8jxdqIkrvDjyZQHNjAu2UcUzKUuB1dx3Uhy+/xA0ty42don4u2D3f/2i9FSM1hYWMiFEuX4
ToWDKCsPVOFn3jY44UvZ6nbd8ylUATLzBrrqblwNOg+JiEF3VXPz+sCMSyRpEjm85yYqwb9MHz3G
jo8sO+wTqCCmMBS1ubkYEs4RrV4P2p5DX0nXrWmy3lvCX6Gz31/jwPnjZt15syH9qSIukQNSZ5lI
BSkijQI7Shw62J+8yIHbr0+n3Iyb1ys8tPpv4FmMa7Pe5fOo6xKU6qFwSgzSwWOvYkQDYIceTvT4
uhnxlVxzxpO13I/PXFXs075MCvJCpjk5SbW4a+QOCfWrJegJYRnPPkTnuVCmIcdd4A3s2eIQuUjy
mFLLvuowWheDPQckxHanZuMGrgu0OVByw147F2udhjQ8exdCcDYfUkVDiplmDQlsaBsxR0X+XnVK
ePtfACNXu8NiPqSyYfpQsuiX53InIVee3dmDgRmVKbRI4IHb5Gym3Bsvj7r446S1UkPt77idJJkc
6txeVzjkNqzxdFFFEnHrR8CLJNBgdmr/eQvcn13dfH8AWYeftNP0o9rTSqrloDrv+IGqQiq7Llh5
V3RZF6DJ3XxNDE0Pyau4lK0otqi7a7ax60EoyeFrdXlHdHwM2DdTnATJFjGhTU84Goff0d6wy7HT
8IHDCjRI9jjnbd9RoGtNA3VaJhB4oldqNwK5CNc0NVXIz3u7lN7hdtFHoYFjvTidQAC16/fkbd7r
RXAMuNZ6GJUOH+iqvWVGIGzQxwhTPY9i0ZKsuP84jUthiT8RvfFMZq0TiqhdI48vjRKctJrbY/OU
VZ28N/qngtItQ2GIIuxJrrlNmiD+/sIVb7uQ8fhpi7NPHvBxZudS+6xGQatL7JT2Lce2+AS+H5Pn
tQAEp54XuycdqXYpJVKIUJn0CO242DElAuuiOlSkUy9/xAqywIaa/h9UYmNSPlQJHB/zoLJZrpa4
2Kd7tDaWP3n22fjsxOin9aWzL7Dgk2qA4Yz8lNrLB+Byoa9GfH6ysh+EMjWfAf6pVpRDGdfnB/YE
iMA4iczDWS2CSih4tPlr9PPXWjOmjvb/ScI4t1KXFtHJH8ses4iyQm7RPPrF5IXiLxqi5btM2n9F
fEWOUtAfQQmBrfnCBONfGs8Uelbjs091ECjXIr6KAyeKyQfRQ7d6o6YQMqfefQuLCUbyoKtjBNSr
gyylB9Y1jQ8pAjFfDXtAyJ5fgSpRpeg0TqplqbCLiNKef6jmMzUOxtdnjlOO1n/TlkwSrJFj3qdH
eI02dAM6eAqI/J7lQgMzNiJIjMLiw2NeNskZgnHlKtpt1AmCMKh0DKosap3aeiK4H9GNG2O5Uwqx
nu5z0krvYd2YsewKudjVSls6V1PWMES16IV0GsatPZVwvFIFm3j41ZpFq+lZ3EHct6gkvIWVvCZl
8I9yCMeQgvGg9RvqZMVGKfUz60quRpG1sY4oQahH+Wjlnaak1nnaUtS6pCkf5uU6DpI2M8S0nQqB
nZX/Iuo5buBy2g5QXJltmHBrRUKulJDCmQWp/ELfgiIkcRlfnwp5FTzmdwYuUSgXCNDlh7iWLUka
WOCJYySRbG7uxQPBSZWZxFcRoozNpZKHrIWGBjvVrkSLw1xdzPnwXtpu41PLd5T4ZegVWJQr4RKz
sY+8654DNHyghRWIBcyb7b9dVMk0aQGcfxOS+9q5L/NZ3QaAypsWEU+jWjE1pdQUSeef03JST3Uw
s6maNPUfUjAXvgKDQwlUr4deyT639oSlMtsOsxCoNNf/UrVKvX3WbpzFCCZAqetkVV1S59mvWZ/s
ZcrqDaUskKAUT0cOwTU6Jpco09JUuCekfUrTDsvQKT06Ncf/+SipzClrtitLVx2AlMDk2XbupjCM
41D0LovWptkKPihcyjePwJOKLxNlLML8oy3p+A2jbfpA9ZgJKWD/8gkzk1gPwWs0z3IVMr8JQD+3
fMQUDybgGl+83+kqUBgOXJvnakW1W3avZuWI6aglyy/7y5qnjfKvOZG0tFUY0CAtDi/iBqgnibYu
57amLAPnxl/8cE9BgXUMpmJUIa6enTBXicvCqOc9+gzP37Hap+Ig4tQygxcl02DXZGDJ55JbSd90
VOYlak4CgiRWkzku8TXJhZdP7jq8WN5EDKNNTgxGPiFOBN0rEFNIs43CGkC8JtiM/rDqwTk4aTK1
CIKRCr0l4oyLQ8IDmLgTekhgrrd5iGgiXgUktDV74DeV+bYVCmkrY5pi5W1mtyxprvDKBzs36WDQ
BBC8iEhrTc1bIpTBoQFqPSzggZ8lLHsItz+ewz55N8ttbony8FNfBax7R2Nlqby/+djrAmB/50LQ
++gWij5ryL0J/3LdpY3zzgssi/nLdz9KGTadNoPV6tS2ZI19whoVo8caFfhD3UUY86eQbLIsSnND
OM5xsP2bj2k5KxWNNV48JsOi7VQ5V/kxsAx5kBrESUTGU1R5cRYciwi7nmLLxn2idiXTwC/6F4Ik
Bm40ha6y92EjOHGFKKI8ScMUBO/WABPy74iZImIQTIfLs86zy+dRbJx/jcn/E+u0ufNowYbch2Mt
E0hv+sQA9QNj0vgFkCRtCPt9W2m19XBMAVjW2FCf37Jduhn6AYg4LIprixKNgdLSnYHWAoLY0CcN
S7Ckv3lJaSLG+aSyuT25SS6+9J45JJgnqQXpE5JqcTuFz4Cnyd/+GMAbJxI44iK2faFBEypkoi/P
Gc0UWbQBeYiKFBjGjO/cR+FUJANUUjw+LruJ+FPf7LMvtQQeeKGkTV8P0UL0jlbLWIfWmtPG0Tsb
jGhAQ9loRtdwTIeB+Ij10+iVsRHHAwjDAmm1EHI1krZ3JrTh8QLTHDuRNWtV/idZDz/RwVtrByNh
nhmgpRmo0M+j6/frJ4E0heClCIoQVHRMvEMfQIfUw5y0TB8KAnsyE3Bm7Rj/AugvbXyHAEHk8Ar2
NJGPCGfDuMz9OkUY+0i0ZPDs45Xcbrl7K08ngO3yqu7gvD0x5VWOygK8fVOQ4AjV4gEHch7ohW4Z
mfTWRLUlP9NoidssNpuISIMEiOYok+nZ+opopG9Vdc18IEm3AQarXcuf/Pf9e15SNKDY6VIMeaTd
J2/CA7Yx3OP2TVY/tFu+whSJxUS9WXfZmodkPoLpphMcIAgPnpIxx6lmAg/GXDaLxXfv8q/Um3B9
VQX4mtsKIQsIuAQM9G63+XNhD1pA+cY6Az+DP3izFL3gL47YfyXT1K/rsJBwhEqL7zYBiuNIDiLe
8o4AsJqrG9AJ0icpY7D9qMVngb7Ub5TdJLs59XK4jnm9DLkpngj2IbMmkvaDc5ZiGxOKPikW4D78
jl1dTONDE/TqKF0XJAmrBer6ufwecch++CTUpKD2JjuchBzhOL2inbjae3Coqlik6A/ws6hDamx2
kfMSnIsnuO55T0SKo27O848/zbYexmGg0N6mPwwKQMH7cEjOyfLL7n0nc7O+F+i9zWOKFMkuGXgk
9gFVL8Kv+vr8hta7qMsptcRqTkOmcy7Pwym+Mcq9+Wr8lId95hBxCitVaRPZbAS2DdINcycmeO9H
fNVRbgjH4I0Fh8btCtGnw2PEaw+kOobXMEwaXjoUWKaa3gnX1FBrT29Mg0pAUuFzUnF3bnK8N86f
+bhPTsDzUfKrqk6G/EyyoVU5l+ap/cQh9a7ojEQZa8YjSq/iCSbwTvN0wAgf10geDlJ8rmRHJTVp
MQmVCg467hXf1wnsXn7TKEgNT6kfqEIihtnJzhRqDQNiV3hcrekzDAoMwu1+4MPfYvJMcRDclI3N
wDzWfACprH00iWGOMZA2MJgizn+ZI1l27L8EB5r4HS7pluZ7M5g1ahblz01MwfDhm998edaPS9rZ
Eqgei3YoQGciQQJMqDNxQfaigzpEkcorJiDF3C32OeLweDaJbC8nhpBHlYmWX+otNi+aSFz0ieSb
uC4NS2Bkg3n+nL/uEHDkLAKR/6/v4MG6pgAP7dpVCHOm/0w/AaeKzTYjOrFvkvaWUB6HMVmBIZG7
kiMd7A/r8JOeqJVXDc7qgVlUtsNlYFOCCVqj/h7VXDodmNzVrCBa0Sx78YgqEOqT9WpX+4HemHZ9
yFu00FHwcyieOB7oEcaHZKjPlz7vIUopGEnTxdic00yLjygGa/LfN7fLOjCD9eB4/W4iPkzET4J/
yxqQu/LYiebP97INYoBpWuPdtPflzl4L1vpy+YiYNG1KOThUyh80iuj7E0Cj2kjkKGMemtUM9gGm
VU/tpN+bRtjNNavMSIJDck3NjldNC1sCabf21YpAAUBtAUAMJfCSgYb0ya2s/K9BdstROG15ACfp
1Ybc2Rddx72zten8rFRgFMJC1DCsSU6/GtGVjfCZ3gVDPBFnP1iLZ20VIy/+8HOfzlHZI2i9ZhyW
ddZHwMwhWARFb/0RjnbK2Pd67opziImgW1HXNADW7GluWLc22db0rxHHnBeixpAuzZHOK3QRedZl
VyF6D1fdsyZXjCvmMVH9hRXhfiLBfS0v0uRz/qEoCL8LgHknoHjQwZ5HUkxiqRGbx4sCVrLrjCZl
Yp3Eie78ydVNjgKG2NL6R43UJQiCNVry/oXNOOtvCQvIgFwCDgESHBHMDTw41o7wbpMZ2t5W1HQC
muJgLgSteh3ZzSX24CWdtT47NpHAiDFxt4bqYjari9DS0uNvvrlAWe3R75HvFQwMLE56+yottBml
jehfWGz/PNR5K6jBh9Fd5UTKwpLOl+2JzgFVJ/jD6yQC/qhutJ6gcSAXF8GdVUGgQwDWCZnUSseH
fe7QPgTWwZRwLsVefnh9MOt4UFpjUORlpsqiMqzCkC5A5+eHTN7spa2fU3mZ5cyv8IH3EzOWGdkn
JfigefzCSW7NpocFrPKaQEjCok5lsadmWrlkhJbUmDWtiO2NU8wqkoT5hOn5WXemtstkkyvuNBcT
wqvM6BWN24MOSYgkIWRse7VZhlPaIrFbfo37ZTgFZfNIBlFo1SYoYeI35dc6qp3j4t9BEzRwvNBc
pP365lWlbuGDgQHQ4cYMXl7fqjw3aEIdRqNbiz5BOXV9leWwo6odqh+v8CiVWFDlWnaGkMXK/EJh
4zH0z3H9c+ySt7edOn0exyZc29MFwfJ3STimI4IyxjGuMxloTcFJUlnfJnArubI55YqGi2IGWu04
0BYusLjCIgHMgaeFl95XEnka4rx/nblPUFpe4NWjWR4ooQd4hGbYfQd+FL38h5Yl3yTsalkj6Cjt
hS2gL3wfWrGCqtP08dbD4l2rCGMmPYWU53BieB6dYSiyeMSxPZRLrMTmQLkrW7XG+BgMzicsEB+q
IfWir4oYBpko5wQOgfuuPTnFUommDA2Ue/G7qWLbN9CGUrU9p1BYVXHecfDF/0qox9/ux3IVPnaL
KJo7fJ2/vy1LDmszULY5hJ2AYnjPkiJbUWx0g5/Ku7AsVHPbQy3cfLlUSJ8hkBO/9VxVQt1H4Z7N
AacJo4SYL94JHLaOcWgTzLzvaZTtnBSFdTbaq7W67ovNQ2JFcTnRpODSxbhXM9vIMPRD3YjS1ABU
bqCX/pLeurQQforpxshHSBq40hh4AnrqSsMYR4hImN2xaRv3UToD+Q4T3J0t5yWFs6DN/TMn/zFL
PzTCAPeTPuAmIiFBwuIm8miiIt/vi+VmehdAckh72EjRFvRbIXzwY8mQJAUPML0Z+POxuY2hmfLI
2zHtWvncsSRsSc3UUDDp695KXT6IhFlt9YnT2Hh90u3ZrmwWIipTjAkoXMWo3PwI42gfmS41G3ey
BoMuIujs32iiTrFNADyNLhaaJDo+Sw4a4SBJ8Hc+FW54Ol9vw7qdEbgzrXlMigEkxMEQfDA91rYy
VlFlcmx6rpTjs97+LDX4G6DxKyTLVUbIqZ+Cpnn8geALNeWymbMaGHpnsBBYfHgwNvIPCeSrrhe8
sO//BJCYPUNcp07iLZHSp6EZ27AbzW1pREHpWF2lJHWH8j9tURX796pLFZW1Tzyax0xOfnACTBor
/+1nKoudI5P7IO3MVyNf9uPuLXxgj6uORDXdD3/6Hg5OeHt6uWvxpteR2GheBloZ80inh64grXTq
1a0JD7B0vssMyFcJvkrLPSkSwjjvjYSa94jZUGk9HnR9cTt6lxyD0s0d384e3TmdaLrlHwIYwl8i
PSNjSQVKjBxyDj7evRyhi0ppNTQuLLjB3vu4byI5Q4gPZs1UPdpnOqMTSQoPgUgBIvpn5hCfcRzt
Jig/2tNmXKZ2aUyqmZ3oHlGJJjUFcUPX7cJARhxCSyrkUnvIOI35bePBh88V8rOfHpv6dDJfhr5N
tU81EUBmUkn6vPAtq2Pew9/lRAoZxSg/oMVEAo/rB+gZRe/Lh1T66HOap9jhUlwkP/nC2PGJJ4Bi
1Vg539xXnvDRy0SVGXjHLpDHuYxwTIHoCV/ztPTLWWMckiQkWdzU+pbieet31INcT8ibWVGtod5C
bxlMIWn154zuJ2M9+HGuPFMpo9Z/335MWAvVHLiEQzmxl6fmQsZb7HCYDokZ+pR0oqqCVgVXYhhi
Cijmr68xPB8Ux0bVMaty4yQF2sIa5N6yGusXmJzVSl4rEUq0kllyVXyEIdfQzHZuCXpLOt3wNnJO
kkroJFuAEwgpybKE6w5y1EXIKB0oh/Vq75EA3NYysY8SRITy/52NH99IDzOPKytkrXL6kDvZmHC7
WlLzQnUlg982TJgaAssUUQHxPFfexMGW6WJGJryqEOrRtmA+jQMkQft7gXOip9jb82EKcPGQLFYY
rBHDne3z4pON3iwbwblusPWMC6z2KREeb1YHObTYSynqVMySQkLLHwA1NFqbcnjJfZAcmbZut8gk
3rCs0BF45S5OrisBhUzDPsU5fDzFGuN/BuQfoOKh/m5k7E4NPppjYf+n3T55ssF97s7ZnYEA9OAp
Yo1QgIMKzNL6NN/H3HKpmIYzRA0tEbbuVDJcW5KnFFWIZso6xHV8AyIjdHykD4Wxwg8RDV9jCX0u
SB5PgRUuRtEjm/irVGu8FgJ3ci4BgcDYnVy0rRoG9ME/rZTbRo6wsO7RkrflGPnTw5jMzO5364PR
x1LkBrXNgnRnkq8Zz0d2oRK6gZyFOrZKahBnK297fyR5zd9hEeNzL9yYr0qoLe3cQMqUMWaz87lg
4pL8kj7AjcjS4b/lgpZAdr5Hmg8FKLeH9hfkV+p2zr6iipTTQAMWcpQYkaHbntyeYLhDD+ApaA1O
vRBPBuuThVweMaEpTPdYJoRK4VLwv7IUE/2WJsgt0HNDgiEmS+7DEbTqRm4SURYMfkr65Ia9m+bA
xb1FPddQT0oj08aYccZZTw7+zj+z6LQf7k205RKjtODSIbp1HZwapeGGGYJDzO1AgyjBuf2Chpd5
+GByXJoaqERDOUsZAjS8X+3NOoOvYLw0QmnB2Qil9NtrCkc/9SachN//whhQRrL/DvVflJ8r+7PX
/XLQcvQfOTwFLQ7bOE+8t+TZby1qWhyFWq2+lA5VAuisLfZ6GH7e5ci2gVJVSnP1YMzMG6LO47/6
aRNZ3L3CcNKEBt+YoPg/HBs58FyqMrU6nY9e9FtJ3rwvkaO6sZAOzfGuopYgZwaNciNTSh7id/7e
gSZV5+woHvZNNMn4p5F4vKixGHOju2fWKNNQeeE+r22T5x3WBzdoTGZBX/GQbrvlO7PyHfkxqvse
lMmbTHxqQzD972U6D4t+Y9fFdWL2W1o3dJ3JbP5qulC29s2XkU0HVaMWkphtG8cu7eu0asfRalik
PELClb4AlLqdIF6JVniMpQm1rQbVp+4AT8Vfjy/TvNOerQXenTgx+90eVHHTcuG/RXcSVdv2q965
cPQXs6EMTegwskGVEimD6F1RezmmhwD30gbAkT46CRqqR00tVUFiQQQVwiKKZJGfQBaq5/S1POlO
MwHwkkjZ0q79VOCgioP3+yxsbWGoBzmB+84Zfk8Vhm6gW9skqjFOx/rqpO4KkvEydxoft5jZbPyJ
qzGU1nmo3bortkft7G1zmhagOrPp9HJld39kyuZRa0VNRIEDCAhlarwhIppFvA/brs3WMUEHPXgv
Dw7B/ftDlh9Lc4EZEMTecu6Tg2btC7A65VulgGpXI+deY6Gnr73tp2kozVT/XXDdd+CXXPYXX6HH
R6HVv5q8pZlSQGIjqnLJJ6iS9Ego0AAQx0RhKa0vDZYD9FzArwdJli0pJxB8X+axJZdg3dgs4Kro
RgpL0/9bnfpfZQj1ZcW2q7tkw1RZJfl0mg3P7nALgAHq8PgecBrhTnitDASw5m1od4ypgr/+dGXL
WDpXGsRwCIPHGxhSYCuaGWbY3sKb6tkEt6tdK05/Hhj33YTbkXKwahTQXzPqx7LqzT3zvNjjSiuq
N5MlQ3PxHGg4u4UPED7OeCGVtESyiCZt++JISJCZRsclWW1PyTA8Whdc3bp7QvcY038gFC9KVjqR
6E1xN8+DmTSRwAZH6GGpMmEXEe3RnaxjNeOKK+SR6Vdrfgw+38TmN9DMdP1oCUHD8PpMr6WWaptR
uO1hKVocSh/HithwoLw0psXFLHd/nzHZlqRTfHr10SgBdQwF/zEtaBb42zoflhr76u0Ov9b83Sxq
Yjset9tjlwLRtmu+uMU/naI861ryLBlU2t0R+yW2mjzBpwPgs9wVTns7oVhVV16D8nUn6LZ0RWFR
opRTGGChWd7enNTmbod40XouCeCnUZcxMZ1obAYGYwaeuPWG/gA4SHbM3gRQTpdjcffsdrSsDmCF
jRLzkRrYkMURa2WZbIPKSnZrGKwL2SNmUuy1uuiXVd2KmpilCkezpcO47kV89SD6ZPBbJ+NKppsM
lTK0wLkHG7YsTe9t9XYP1TGF+6ayZL8xcyGbkyJBavsC7iW0YD3L7zGkytt6X3F6kb3+iCFpshkd
+fl6A+lTUzJzBXk31cB8guHn6lbssTYMjmVQ8HmLNtkjBH7i0wlLNzzeyNh2Z37r7KOlJHlI+Dqe
r+jLyZec67LAOHY9My520peYAv21N06OPD2rkiLlE0vhfMoxCfXQKaMl3KFOlQTDTy9PuGKqg0RV
tsiU8JLXcIbzFR/6D72EDzhB7PRhYQWbUOgR9BwYS/WFjnwRe5XwYr9iKJ+eCQJ7trkU62v9L7pW
q5RaGbb6znXWkFe6EiM7YpFcUGLwAlyMEyrifBI/6//4YeOxbOTDjAv6Rri3tQBYFLw8XhajAsd2
dbikOjON7GlYH9OldtdcdA/nRc/c3jrSbY5SInA2VwBeUctnUGjNau4GOVWC2WVxifVFjCNlQaqi
+hzNXydzUZAkKl5YM+AO+og8UgGVma/379wOB1KRwUKa5kL1DBJnIQxKNMaYnV538q7VJoyDLv75
yDaCADfRZ/oLFcIYznfZBz0wqjwIxjEcy9l2bot2QSA4Ia0PZyq8rDUx2r1FhfJy4zn95hKFGwd/
MNo7nrsbJ+JKz9s9LMDIia4fmx8CyiuT2WzezozKjNM5bblOJ0z6yPNNHkj8WTCHVVj4cJOraP32
727faIBfn0tp6+zcBRFePgU1j3eRaQ1KKMQQkVjrer5UTCT0v04XtlVFJCH3O3E77PzBFAZvLowZ
ypQl+LQ7fYEjLvfqB8ZFwUBsXQjYzHU7Igdqqx+R0eiQpj50n0WqenNTJSp5XmK9TaitpnfT0GOg
ESVVDpYguipzRFL2u5uh1/Rbgor3GJOOIRZ/YTpuQxp8RGhUdJtcQWr2LFCDjefwr+/7KRqh1V6s
OqIcM5bw018969E1w7qJ9pp6ewQ7yjmrGAIyzM2uZlnTU0HzpFdNzrgyAkFlYiRC9P5TAPJ7pfsT
b7ne+YQxVqIznjJeh04zlcwYSM1yPa3rP28cXz21G+/8TM++7502ULcpnx7MhjgRHqUzCfdAqnyN
HooJFbscm89R1gP/lV8qxIKWhlHKk8xa/vYSNS22WrX3YuGlr+MEKmC2E5JYnbOIAuiHO4wuapwm
39kJJIlZlYGT3ord91uJw6/zmhTHbSgZMDfhx2ls8jPCIKFe8ilkfbBMVXCiNyUNSTAHdmCNObK/
39nWW5zmVcM0TohVn8NlC7AY9tJAXYtZInMymcl2Ho+cpyaYFQjNFmmgFmSoRN/FK7B5iUaxUZth
e93mUuREVJP4CXtxBQgpJ8agcCD3cNZT3bY4YIEin+D4pRDGuTiFDPkEZiv6ZRKXoWXxRdPQXYvF
iDyODC+BtZ/l1oNp55VU+kCsKYU0kb/Pl4D+b736kfKuKqB7Tp8us8dM/VLeLoZ2WqYAobb20z22
Xi0eQ1QxGLEe2JQOGHe83ifdj25LmiNE6CUOoSrfTGpB//mJqHB/o2ep1UnGz/OwC21mKOmBzp0K
j1LL2/oxt+vANcqyY4y4dop4+Wml1CGy4fhAIUoM58ZJxQT5+LN66wX76oV5s+spuWhrwTAifxIu
QR6awDVTpMvOVsoTbb9lzMXyePztoSNtguyZfeVTEJR1cVFPOxoPvsX4rjsgojXPDacKc1qmMm70
/QF70OCpXT7zYdE8SGoI8rR4KUW/v0ozUMeGl01QMw+R07388In98/WiaewinzzPN7pNkenfQpsg
IdCOCRhWrGqHmLMZ/IxKto4Jr2t/W+Yl663/mo2L9lVizM8kCOBjF2RJMsLifYyLICatYulQTEn4
QMNsLjgxRR1iDTWA4Bnm3BFqeDvSxbMTJH22xtTTllDXPA3fBq1MpLseT1wsnwZq4042JMzkC0EL
S4JGR7oxqFSJgha2EWU05cGtBsyTLFiNJ1CYxWnVSNL0SNzEUWB49aqZUK2jfhXQPtQYZDPHpg9Y
1VOvZZrh0SCjzMDcviZX5TDBbb6RmH8r9d7qzRVHAPRKtzSbfcpaou7VBSez9gT2W+BMKo9RW3Sd
r7OzyuLI7iUvJQB1QQD/st6HSIZvN1J4flNbs6jfZhQcg9kt3XiY1jssZ2UnxazWlChcIA9Nn4MO
Nc4ROpnGBksqVL6G5FTk1i7M4zFJp6Y7n4MTZQjrAobNS7GRzntTghfvoL8kUM3tSZ+FybfMzcBm
ul0+K4ICLmruhN2RVB/QpgiLZTCodx5pCHUGqJA0+mmGnJnvaZyCtohsOjEHBSVSoR6jQIibPyXq
4YhKF9cNrWXfFopXsf85hri/hoYTqoBomHj6X8xiyQfKoXL4sOJsujpDJbjYyAQlifkgF/pdObcP
i95roYiPR7SR7bh8wFoDnnqghCHwpZrHlC3SgSkKI0KmV57QHa31gVJuF9tPl3usWy1UImhJDJ0L
rGVfXY9UCs0pNzjk98vF3Jw17VZVT5eTyAgM992orfpuLvGZuvXJtuX4AUPRXWI4we0nU9mZhzEV
ADvUDtfJCiDaBeE8MsK1YH7qIqlaRoqrkZ1ctbpAEHK9SVR2uBx3aR0we9q0xB8NU9S1bnckOGmG
RNrpx17lSoH7SBiKZUOn96awZivnXXWYs+KgS6RizpTThTybR4VThJzvqo47LcZ+TrmLwPEM2x4q
5jZehcmavlG0rwksp7gOihuySjHyCWTkdpAceWoQcB0MsJjAxn/h3HFTMnOegaUaWT7zKKjgxTNM
iLsee59HPCGHaemCS88efwU5INOJDvVqnz0wDXZraTcDoSBbfzZcRehDrpmwYlCgedC2KfdCUihf
Xg6Q6lhaJsgCvJkneHCWuGTMa/X0sAky0xsJmyc3cxHonVHLvbcrwMyAOom1A5Zli7Ldg6lPKFui
/OB51b8Hks+eCxFZk+RyDYBMl/O1wt5Tf11Ifi47wExvffoYe/eErNGe83Mp6ROPIcoFC135zli8
7vk9bPbBRKIRfGNyVYYN/lrR1ph0iXX2QIYcL946pmyPkjYucih9PAeOqSgmnVZJpUiqqZKImwcl
1ErLTk5rtdJaSGnUOHmElF8AQgCLHQsIqW+hiL/xYhDIpFtjKLir1F2DVFv98VqpvrVbp0exFLX9
VWR6M0TwYarjt4ay8wjL0tTVxvASAiAp+4ZVFFFoV3zYrm90Sf1N+etKb+mND/2y4pWW1Mk97xJs
athwQtG8VRtKxNf0Z5pW6knt95Yk3vhQYUBolqVD7W7FoAI1QD9UaCr1DrD09QXFRTfyMckajz8H
E4qB6fSFgguRpOFu5WI43w1Qi9I+k6D387N3lG99ysQ4htBPpjDTflGK8GYeSqAiC9eQyLsklS+t
YLoMJHpgq23fXVTZx4JbIOxJGJKe9NNn4LIk/jDd87fhbNmXkNsJ82X+kW+cbDJnGiqEXHeza+6K
rqP33CImHJ6Qe41xMzjZFbcVcyl9ZjAwzbbdogoeVtMGKEedubMu2vgvLekGcvuOlwiURyhrIshz
FlWgzLYHJa43di272VbMHnXtOkdKl3P/p/2VURPTZJhqNBORpxOWeeJmEzQpFMphSvY9I6K/8ulS
O0SywqksMNinv7WvUJyD0gCbty2aE17NKtADFxLyxArrP47nCuXRatQNB/atXJTUa51phDjpfEvu
cU7MBXK9u5guyQ6MYsOSka2lVirn22MAZ3cj7FSgxIdP7JMLJ6pJO2zh/i/uD42GxFl4A8l8o4Ef
GQNEo/OjHSCjQORKTeU3Au1ps78DD2Q9p0DgpOgCPHgZYjixKmAyio+LfWvcAN2GQ+hpcOH3KXNN
cOlPL/SPcfudhMLnUtRtu8+57WhJeSfifNDn46gxeDghV8G3GxMpE1U+6qG/AsP7DQT4Cszy20nI
XkJCJaUtU1KtyYyjwDCjc5kQh92bhX43t+VxnyWp313n4bZEnUwJOegp8YTAx5OXQiu/YEZFA8O0
UmtU5j1o8idlUeZwSNj4Xzb5MgPRFVWRDeffIObMPsknbvdqCJjq+veKXOOxoU9GmRJnCcDOZEIU
LSYlNlK1lIYQ5KDS3VSFwIr1MGba5O2aVx2kLC4Y44mQVeLcbOrqfiMbGVsHN7R8IbBYlJkjh/kn
YipjkOD02SdKiEpQ5DFzT8YOVXljqXCTqD2ivzw6R9OVFUL64a09MPFuLlUNPYZW6jhQXdp37RFZ
NWf1qjCD9w4Frb//Pd0yQoq1U6KtRpx7P7kpSqaWRPrAkhpV1H9Qarnmb+WREEHSJdeGuamtzaJR
aHAYW8pfuotp5sOwnNC9yB5E+sGw9n7MKI1dRSVQ+Kh3UiAVxyPF/ln27tawz6mef0q+jRYIS4Ms
0GLPA+wROcEGUQYuGnfl18EMNSvosSzT+ohmKosPrIjRJnf8TGj/9gW3HC/0/rsBsaMo0bZ/PNm9
nnWMkF7eqkcmiRINncZIsQie7vO5oljYg+NFlDiU8ouH7aOCHKwQCkAUibuQA2vtnWj5WXSVTvD3
a36RHxr2P8H4J2fEQYdRKrlOhvUiUr1QvNwS1UhhbHh/wS3yiDdOxE4cXp0391qz9VJu3LeV1dF6
tB6x0RnspuXaxOWgpfgmLe92XDpcAX7zLy4p5lYim5c3P4vGDZohpTTz4c3+j82uW0tsA/Zz0ksa
tUrsj9fia+of4Gpjd6ZL6odj6D5tX1XnAvELCdPoqU278XdtEdOYy6Hkjjnw6FE4lUFuPFIKyMqg
mBcgQs7eiNpPZKEPOCNl+4fy0GkVqKZ/1b/RyzNv0L21opHM33BuyzAlL4H0TT7CnHq/HCZT3JJm
GkD1URKW/o5Da/gCfSpSZGick+Vvpf+F2GLxxGX45H9xAJ3sQpYYTX1Sj4MTwlxJJ+plWF8irYMK
ZobUaG4eFU95Nk50h3Cgr0d2FO6EohKVBTArzfYPfr8qRqU3BhdhC+V1vTWt8E5hW+nF6xOkIIjB
ueusPYaC0uqgfn03sm/C31PyDlWdf9j1h5FaHtdwm6ojIuMFCpTi29i/9tJj8hWK2aQNTNmIjJn9
igWvHTVqU4HBn4TnT6bCuznD1sZdoWS7fWnj/SmkFUGVUV7cSzU0Q+SjBT3yJ4nDFQZs71hRD/gv
YKcJ/Ts2hzxDNlNbUWTMzxCDhmNh7ojbTEnXSn33YQK0OPtpUptnoC7NB4YYB6LwZ/9k5AF+oysc
cUFEgu4RLoXC4nVx7SmHxcUN1kq1CVJ4lfYHFwi1gYK/0vdcE/OmfJDh/4WGXtE9ejWVuB5/Imku
ipA59QkIYx+gfECNCrq+GvZ/IIG0AuyNQB/tVdmy/g5EZvRPSbAxs18R76+nyQmFOHRD37khCFGP
K1RLaspRG+qBIAinMe3MLDKhrXbfzU3J51aBqrhKEknu8i5BmkU10HTpJXqIIaUVfX+pbuymu4+7
BxrolYCwCIb59DB915BDpj+IA7u97fBpTBXTG7tCCGp/Fr6oPBSe9oG5YAyU9kDSKMKjV+dKfcQ3
JT/xuf4m3hmYE376004aksrByn8lFjlfCHQZuv9kW1884rcIzoLIo9K7YNw+Hpj9PvFq2E5IedOP
BENITZGkoxN0v2QKwxYnOrDvCOJMA0ogHOYOn0/4GUTv4exXaYVmlOeDrSUtDlZroD+jb7f6dThL
UQQ6qX09zt5z19TOR/iwuzZ1OuF55Nfy3aaZGOvPaBdgTfoYqF/yV3+kYjh8+5uDDrnCHv0ZM+N9
MFTGQ3rhVPogDV36YAyGFFTKTvazuwLt/1EcapPUJGCrOy0XbNM9SAov8QPJd+tgzlwCKbjLYLdH
dqIZos7VSPrdGUD80x7TnKuY65ctaxlLD6IpYTLSyhT8aQJHJpufLMdL/QSseYBXCnshDekXLzIL
FUjTZQlXRzSKgME8ojWja8GvTK9fiEk4Sg4KmmUxcTigDNvbbCd1VOpoP+6glpMzPQXWdLzCCfdv
GtWzTlp3e/ASWu7+oOKwoATBOLKTGryAsq7PY8CPkQ8ljsMg/gqg/rt3UAl2HERxRE82aC72+FgI
EkAo98VNNxGfgowmm0+phshLXqBdFtxxGwsEM3oXfW9d+6182x9QIM5UQGItmyXPbJb0fi9QhuXC
c+fkOGhTWHd3sUkUl3gl73SDCczAY8wTL1/v5CVFaUPcd2cjqpTQV1Lztnd42l9fXM9IlVdjltCL
Pz3fAgCfwss82cWEu4S1pZsGL2q4xx3yLbDDCUadbKpLPth9YpaQapmUryX1J8vbn1UlVmGWGwzl
VzsDsvcyjtylJyNuXJ+14Wworb+zDKpRLDhU/6HXq7u7XNIIOkWT3Va1gml+VOhIUsmytidNFRIn
iWUqtGjVrHYjh8cdyoi1cCLsuZrIRH930FWlNd5zFcc6mzHGsHS7h8LS2unYr19R+D6te49D9+RS
H/JYQXp1Y/b4TW2fYebxYUCEiZdHIDnePTBuracQ8c9PDiugWVNJPv42a4AEPoi1I9UE0fArmume
8Foqljl4uixYgQVjcbdKLt+xnKaIFkYQInNuELGd0uTEJPpIety5fSbNCfst2EZtVqcv4M4x326W
Ta0eakBfPzMIBGQziWTyvrnqbeOm4BTw2qimTKS1cLE3ylCBOviBx02BBXwK5gN7mNTKIzuGvw6O
ovjI3qmrMLorREnPiI1IxrAZECzVZaWwjZ1vwBLt9jhrakWIezX4j6lux/dMtfZ14lDCgaTj9xwA
K0Kl1SSb8yVFvIhZugTDPhTFTHJRe5un3XVBKFulcARhq3AulaBsFhW/RTGr0nHUhNVaF87r60Mj
x3Q384HXtvmORKipT9w4yyb6ZbjA45UuqsvSLfC3gKSQd8KgQzJpL5gIm5Gze7Jcpe99Vm3oXBu4
OMiZ6yDrql5p6QDkk8CZs7ZZZBbtua4nYqpdXMF+cGIdNT/AYOCtEerIhZLaUqySwXT4GPmagCxu
O9vthaM+94YVUkVlLQd+272XmNFecZEPOSLT3vCzV1LAPNRKjHobt8LW1FcWom14iijiAUxskzpX
O75w5kP/wQeazpEOAF8Azpe/jaOaqzogrPUMHeonC+aFmHZu7wSIl7Gid89EIGNzDN7xb2nXtkQk
68+i5wIV3ICnGE5cZM614UoDxcMgFkx3zLiKdfO4i3CFXER4USyE5rUmcANSrko7GgQzU9CXLCTy
Pe5y1N0bl/0CTI1hZNv5cP+WHoQlwSxfgtYK6VkfbNO8byjdxVmHmx69y7dQQ+YpBw8+Ewc5ypIs
TxEX5AZzPsuEAUEAIeHA1rw5l/I09pSgVhbvalWUmkNBHmhv3D/pFJQyJpOZY+ri+Nr45xujWVsC
raHsRz+y4g/JCh9PPXxvZiDCF0wYpne2IM1a2HbXn3rHCCWr5F/gye64pQ6nghi0vMo01Xbq90wj
TYJd0TKl3Ebe4kAbeYHMT+ha79yjS0cE1tnww+2DCdrvvrB0+0AAQ8cvEdUl7TKz89HCNQ7bKu9i
OJLWBdOqMZv5noIsA0mqdBfm6V4VkkQHzaKVTzQXrLhSu0hj+ZJ3vcMiEppECEsltyJhJI6Um1ol
PL6aA2vmqSgakq5mplVqDeo/G7gmWEzkaQWaMtWkvWzSBXZM8IvJVR/KVExpuiXNw/4uCY4HX7BZ
lshS5t29rsiQWBVIVFu9USI70hnfFn/5zaO63w9GEEZKHbxmPnj8VkPFw79/+ZEflRAStJmcJxAW
vRv3Rs0w+D6z1SnNRT1b10cYXvfJujOc/IXvYcALqI963yFE0UnehZkj+sOqZ++qhCQcXubqDjm0
zjyyafuW/HBT1BxsesGIUdH+7op0ocSh+nM9zCe2RSNBaJJ1PL9wpFrWC7MYLfva4AFjF3QnHor6
8R1B+w2LbUjagfeLeshaQwQUyLL/Lzi+liK4/z/lEkT5o3J8hbOk/HcshAHziyAzN5x6l7+uCxp7
atGivayBDeIqAnDwuamj2IO9nlsjoo6+8S+06ua2KuyeiRj6b4XUAtcHfIJEKJuF2pFShAFoEl0R
nbpWVNKvoGb0SdegtEAabNvmlfNNFXPkrCe28GwQr//hDX49xvlLGCyLEaMbfv53QhK0IjZbCMvL
8ZS9xuM5hLsvMG8NuqmKwI4cYt0z/UgDVBmvWQC8nJQPIQY4I/thRX8CYli7hcemWC8cQAdrNjCn
BOhdPWt6/wRb9YBEGMVVvYhOvLUquFgh9pY0i+oiSKpigts5evGNByi/kKcoA9vzgNBVPmxthcnV
lvsXiNBuwY8iTtxEnIZgJcaU4Pwd8j0w+JTHkjWbdKu4KQDhUtJeQLjoCH0KHHyVmHgaPcNQi/G2
pRmUQLiV1WBFqOij0s1ItwBpEtbbmPQ59tC5dSToBFg8u71sWeum9XYBErugN9juLe34G94KsAZ+
a/Dk2fPFcfDB4gqdwgMdrFuID+tAiXlw3E4kkQhalMtgDrxB8S3Hq46ZTT32Fo3FwzMPmrhEowHU
x2JpdcqaKYolhN/S9xdFKql81+J9Ozg93MM3aWyYIOzHkQpQLXP65nN7HYHxiglA+j5x5p8Mf8nU
kPNyI0Adl8nMwxRvsGEJiUkA/zpjaESD4g5iYENPqxKz7IOQhPgvVjzKdvuXRnvkcGYjFBALWfVo
7k+DUHy0rYdbfYZXvoWfOxATTnHhgblb5YUWfkFGGq8g7gZIbSyi8xSOOZ5FE6DMoKEkgNBWTjDu
GIRjPp1OI9u+bzJ8a4blP3e97L+r30d5iuslDdWEbV2lWGoAeqRprQWrdl58ZLdyX5QAR+6oye2p
45JkkYODXbUyGxgvQJVU3mveLDn2dDDf7cvT4bql9PhazedegHRSO51RjKUFKGSsBU22cpAujOS8
8YIswStGoxVT2pbB5S3Culds7KTf/a7D+f23glytgvkGqMvAxSq+OwGzvdHsCmk0TgwBUu2CQ/Z/
PDwmY9tGSllzW1ygRm7/RGzblPmaxk4g//ZJO7D+lkELPhNKouxPauzPqFsbmYoX+apn3ZsXCJpK
3nLRxG4KXPHjyrpoAFs6pR1F9SHayPYezFyc7FXgTaj7v5t9cmP6ov+YxzamS+LNplEXSeSYaxyx
C1GheMvt5gkms0DSfceUzYgraFak8/MQ3KqhRkMqe/1dGqrxLIvdsHxiCgC6xMd/+VSfT7k5hLBy
KbxFskS5n5Tgny4bmtMsfSbufYDzJB1nB/IZ4N/Hpp8ghDPk0lJTpF/vAIzuhwlH5mgEtr7h9MbK
7KdKDN/hEpcVxqpLJmKAcpLjhKc3C85WeCjuBm70rSJ5TpP63je27LPIIKxRP0dqn8+qN5i01Oby
KSehgcF8GHFyoASu4/5uiwBVSwV6cFjDsplO+oNNJur52gmjsGuSOuDHu1e7uShsKFcgrH90JED3
gXaGvd5gKD7BwVD4QgCWet3z8F8eTn/LK3snStTB5ByxYsjA5OD1pSGODzw1iW0y57V/w90FsPgF
SblSuBrOT4iVXq+atHvGdeARbkSI1gP14mKlaadcIgAn/OTNu4NAgR86iY8H/dH37k97P/VBaMP8
56Eo0ALR/Bc6FIHMpP7SUAp8B+MqxuIF+HpaRD0+kqy5IEac6sirDYHNjxFz2z2iBNknF2BdMi1G
0I89lvP30dL7s7dRAvpMPXMigXUqpkGaKARMnrgCGZZBLOKCGf8i1kOZNI4a+8T5s8xmewqvwysn
6uaCPSltI7UqiNmzDOXgdFrHQAUarDB0MHVhWNHuogMtPTHoVIRfL0daYWyQoeVpR71IICs1E9GX
fobZjscBsE5M9YEh6cHqkqYgf45cXjrRQ9Ql6ZKl7N3vafWg/pjQDfZ7oGSBMJbmrdciBxwAP2TG
rSmGuSFRD6EwURkha96YOA+K0Njobr1NaYlVlBCXGo3csqLPKnz2hdavDqPTJiaGO0YUrTpJfajI
9urXqwwgMIoMkSdOc0b1aIhS7NUH9xhmwc1mMtr+GqFngFUITAnaSp/6iL+f3p5ShSf2+BrTexfD
r4/6HnbDAyWwbi/tfIU/rG0+W+Aaj4eEgy3zVzzyykP6/GwCx4GgWYItKfZqFStipkikxKBrLOj3
38LiVTtpFsYDolyvWnBWxBmzqXHU0A5L05I2PYtInEoCTykpkfCh+r4zx1qvYqWgRLxjUQ5gfulQ
//lx6EJkN2PxkRnJxggc7joX9LKiTIWoe9g3jAsfNoivio9dcAoz1PYIz81kLeT6FFzOik1tjlad
TyjZf0Qt42CK9Ce9lHtxbdqWNMeWBBqQEtmviB43JTRC2/3OR3t6gwJlTjMhDTD3/ijZ7yQLh1ss
aKwpUd77ZnkIewhgXNHkWkX4Xxkltw8c8nd4K/TxTgbWxDMe7lp2i/ruTLxrR+5DpP37jR25BamJ
dpVP7Uy6Om/YawN1HRZ3VqHCKITuVectFk1JBH+15ZBhhoB05Fd6oR9fjrzKNp2Y9ObRdAsVGFSI
lkf+rA4rfUmzBoncKVAvlgczs9yc5bfkaAqey0Op+J6o28wYdxY2xENj6dW660hdFcstxRYubhxv
4NN1JQFPFtWNd/Rp39dbk9DTFwW9ijq3po2Gz/wiAAHdiiGUt+gsrBQc3Gy6VAWazuFpxo7LnupU
73MSpJ3wowOxoL1WsG+KgeIINdIDZXMTK2rkpIHju1Fk9zwO8fJV5S4vvAqVv7EVjYOnJzW2uNVG
t5IZV/k0sDkmuW37q8WVSnMpPTflaDWIv5qmr/z8EFAojJ7JhCRYCGYjoaY25wesv6NpBqbIAoLK
AQgU+MPKgkAYJseT2cRPuhHHdlNgLl1j4EDQieA7H79JyYep+RorSs9MRqPd9Ffr92rk54NmhWOm
9V/4GtMrdoCusz/gyPV6fQeJ5/ILnxmS389qNc3pZQGr/w25SrqUpRHl0oRGG+4FyFCLXoy2cZ+f
sbXnPeHK/gaCiOxLV5t25ijKAoWvpWAo1unQ6WdEoAt9MXnr3wSXDVH6dIkxwkRhIJw85ezMVqRX
Ixf3P8cmsqA6S1jvqdPWVEARbS/qgshWsl6slwTJP1gn8PtkNaHM0dQeQEcJfbQLtU3lz7v8MOE7
II1dLURfD+kSBsVvtU3GGQVmSrlFSo23OhYCdEfy+V0h8/D28cMV+dMEnsQsg0eeY4O1qrcYprbv
06PI8x2RzhgzH+L0WRC4w2mw4gYgGzlgi18kiDS1nB+UEHd8dhC0kaX/rJZ/kONR6XgKfBd5nviI
/h4oHMJKWoes3XFngToHJXFpPGzOSjQWt+az7ducEfHMcRtHC/Rpeweqgt/JIau9yoQu+aYyQ3MK
W+uI7R43nz08XEcSi9evlquI/W8GwRLyFFVGtXHUx0UDvi5M8VE4lNtqWYIojtQNspF5vdYP9P8b
dvz/K5CJq1CFHLMvZ4YbRuMYdd0RKqnJ3JuCm7FNaNtgWkIv+4mNgqppQHFfAstQA2teJVunfyX3
WhMFQxrH0iY1hEaO5UPdS9Zv07Bfg7dP5n0+w7CfpJhpL0/nm0HAmFw3focumQV42u/63UYl/BGV
K28UZ5VUAn5VLeykPe+Whxye+TiYRVr+I8mWDyoKf4YHqBlALpDbh4H3DWQi+7zidE1irPkg0gM0
FztOTFJqizVH7T5xijjH9v+93ZXeoTIzsMKDriFbVUu5YtHIhvexdGGsTITJWdSkTFwQevZTnSHZ
lFq7Ew3mvyl78htO5jcCCgn0e4Fedcv6DD9ddrEoqVutpF6RT2ww9cgu4jBSNVgCzff+X4XAFYqF
yTWyCW6cm0IIIx3hl2+cJeCDkAtkfVZzhhCbzGhqS05BpP2xj8rUAYVbSw5jPoDlVv2YEv//pMGM
Cggp/V1O2J5drTpvLDGUV+bpWp1VXtNNcyEwsR4z7MkTm9qlwvVlkodxiS8hbaG/vANL6a0UZwQl
wvBkWk4/08fooQeGD8gag5LRNLnlIn2saLS5e2VIM1nX/tMc3WAaxRTc0EpuuRBCVg491BZOWj8G
fxVI2tnopqmvrosRicVg4+NLfTT1sXDXXSTfs7/1+l9tvCXzAP4AWzTL0wIgSiW2oJH7+Oemxtee
SVFgmnZMPJz3B7G+y/cWJ7CRHGHUx2/52mqfY+PdpbSNl/q1fNu+mYWVnJKooAPCeojGslNOcEmF
Zdxb0CXnWEEKwAnXjOOfITolKH6OLRBHM2K4DNF5F2N9coN6pntxCbTIqwiJfM1o7yNarVooROS1
nouzMHva5AhGZG/wmUoSa8VaBxh++y4V3ch3bmaVC186ZcXXKuQI4l3dvdZo4SkoOMbZ9gR7FJAS
DBLOL7fMadFJG70m9J3dLlhEdbdfj2DZDNgwAl79JjyYn2wpJ5zF8kWf1tDq6L4Op0x+BVNe6C30
SUHt9/0E8x0SYdo6QWw4uZOmT1WKnLjJjpDNAWB8g/isVxPXIsAaIG9aty+fuBBf89uMHDqF/5zY
zrGeEBIwA0GAJsBONd5F5WZR3Tws0jy4tyxpURqWrJ6AZ82+XzhM+Ve+8H1h90DlcLXlBILCfvfH
sEdPZAsFSeqQLqfrR29ceQZP6SaB0A+j1km/6j6NKLUm8J/kOyui78w3KRzb+QSpnVDd0vYkAGjZ
RZcf8lDdeyJebBGyEfKyRHGwLPq00sfa6Bm/S9xm0BEGyWAEKsn04MJUDWXRJHk4yaF4urItUgLS
KDjT4Zmey9InqpGxw7jacCB4bzJt4wBmG7sC1r8ahHmmBQrI+1VXO18t0dVUQrngemmzJqHTlTFj
8nJc/dg+ZBkiLpRxBxjxYqItTSAOQnWpF9Vt7tzWaeyhXSXlaksDzlJTr9rtNZhCKKgbc66K0t9d
LVwDb143bEliMEpn2g2GtCLHm1bXqESGz5t7H4lt14zjletkf/SYT0NvYAI87658yvstgRGsnpQ/
ARIwzz7YXmUaQxoY+G1CjjGLRtd5DDqpjM3CvQzc3Due5VkGUswr8GWB17hhwXseJdUrgpj6Wapj
vQvwdNgmHZYmUIr5oTa2i9ro7uQmpOymuIH2timuaKAmzhTvoI4rclYNe6fK40/UzVBUvpcW8uuJ
uvWHh2DOIpo628ltwfVtnP8dkJ70I9BNdFaXG4f0GltN8pwRJ38rtD+ZfjlQbs2iBzR4jAJF1kBe
7+YrZm2ZDETfJLdGfNuyt4/YRXOLnO/x7VEzQIg/eBNuCO20xenvrAYZZIowxM5kDaXTIzDONCqj
w1gylbf+auVbpFF9XbZ/vN/DIlXZCOk9WWdBZqTrXok+Ji0RLzOSC4WCUkM2yJObVwBU3Qab9bIN
aGzGwEUa/2Jwz6hhcyEHl4HK/rJsOV6yQyOzTuvRp9aMFLMh82UZd9haDwpFKpiwYB3lnrPC+azR
Fx1iHKL6tG+VGgkDjUg4PvDFFmGejZIZa63PZk/xkFxRDTrDCKCiTjr1eDArtpytrCf+lZLDouPM
Sj5WqondAL0vocis1w1Hmz4oVjcJLV6x2PYDZXUfO0p8+XJBGo2lNbVGTAqyvECe1+9SZ+fzLStf
HkfIsc6iD4yD9CzJfSKGP+Zdmq+bHcHTBfDhH14P0D0saoBIjmDUUD30ny8Kwe6mRs8QklAdzQUh
uepeoypHZTRTeQ/i1I/cOmp8xdXj1wTnG3IR8R/bnNFYzh5AAQeCMdhvfww9OomdA9HPFaZyRKcq
CVa80hSkfgCc4z4SAPlBgTCS+A6hGQAbjhCWUBFBlv76Edw8dbGT9NQl8NIgn0pXx8issi909eX8
W2Wk+aDKGuvaP9f1Av4GsIs2ftWosF5zq7G7dD+TmwZwdLOA14NFXR4+hhvFM/AvT4H+tVGlWGRn
hLBusjiYp5chmmRZiHaNL8QeqTy+7Td5Gkp1BGCpCelX+kQ0tLFvL9q9MLKNd85HUiDWZGgmiRj2
tOsfO2Y/ygAzT/JPn6dpgyaOOj791rMlKQrU2eReP5ZHbMME+mIbR27mLkkKlAfYOh6/eE1708La
MCCdmNtuVuZY2N69I8sL8C5KFJxhfs8h91oY9P/41r57ZgwFuqq8P6Qi1nbT9TUwHufqom7MMCPN
yL1M9ZISiyciQ6rTCxzi5PuDpk7ilqHvjy+aSbGozJB8V4bMupjddxFB4hwX8ROVfPJ0jPdQGwNY
VNn1uHu837Sh0z0qhvATmh0K0Ltj0ELgcjNdBeQd3FWqZA3GoMEBWF7prsuoURoZo/sNIVPKA2U+
YfcSaO5+2frYDX/CYKl+VvFhRrLoZaizmZg7S1cAkJ7inC6moi9mw2aEWTOV74X/70+KLwD+WgzM
Y0VCo9+9mJ8T+5+gz8NNHtH906spyg4BS6zwytcvu0xaeS2J9E+U+DnSs6sZyWfu3QISdUmN7WTQ
Hdl0wQJLGoAXA2dIQlxE9r3DcHZBcGH/p/VtR48tKGpgroHQxgiffVt2gxDaE7qsbnaJRpq48EM3
sZGqzQ+mhnuV9HqArBJfm8VfY3oYAkco27c8ZIiNgsdxWVvc62JsdY3oFvW/8pSKD3S6oxMieteQ
jvMCe24UQuGjEF/jBa2MsFhknWV78B8/NAiVAHiuqgYLMn8hSkxLoscZpa1GEIGl3+mkDORSMKc+
972FbZAfrWd1wK3I/cBVjveiYFDd/CWtwNmBiuz5f/c5Q7oIf6JYpeOVuq2ovzzgSaLhzDs1hLZm
Q2tTKOkmi5c361OZCOSdhdYRB6nNsSb/gGD8IG//6jsB/xgerwy2WGnj8yyx63kv1Kp05/Zw4mb1
3C+/2podI5M9i7aVi97ujG7ogFpCrBlTQ6VK5e6eF1Dz+vJJl50n8k17lShQ00sQT7PIr1/PLrgK
k8BOY3ZWR5Bpqb7202YL+7WTGnSHxexbTsc4AMDeRTrAuUulvAIRipqE3+hebMUyyFOjrf3oEsXd
NuF+RtMIb21XimsXNzzvkoqVSBk/G9aTLtMhyGBv0xdLXuONOibnMbSMeckuRpDyKJzyMX7it7DN
NtRlPfHk0nlJREFcSdnCipofPhzfrtkybL3j8cCi+iuP4n9qX4EAz8XsAqj6rVJcMEvLvSv4yagV
rsA/YR5z/nUuhDhnB6uJnT58vybdvJG5no0HPwIYbT54v/dlacMJ5/NescHIIiWKhKDAQzgPkRbY
TC4qbQ5tPiRvPk99ZkuVMehFcsc2eVzOZazBpF852GOmdzd48MHu7ocylTfIokcXx5t4iCmXnAzV
KztCopM9YpxOQ25rvh7TbzTK9TDLtCmIfe+6AeWE/PSak5MfboAdDMe/+z4j00A+Xjg38lYZPgRQ
ExsOFoyDdtjmeSbRzyicBl/A+zfExI6DjQXP2eDfzg7CT4RX5buc82vcXKRdP41oZdd33GcL5STf
5T30/1c4ZfAsTIX3d6FXSLqYwU0T55LcqFGkfo+vUVKNFj/NAa+DuEVJ0EPLVURWEf9xEEjbFrKa
boACra5CdGzDpizVdggLPNmZuKLIw7DmrjeOP111tDa9SecPYW2Tda8DEUDwY7xWKg6ao7Tume8Y
wtwLOmuzSsBpqSJq8okkKQ2Z6peqK+8zx4BfXpIERK/50uMnLWmnkivOlDhhXKDzce961h0HvELp
5+7AVRSluWeugr0Pf1I+KrDj8YY96zkVmSqFnY9PV0SLU/XJJGqEcwUY+/+2XTb6AB49puyNnU+e
su4ZYkNswxNN945suei5in5BQlIViGJ9YIS5CvTip8ZQy/rKj5hPClXWmF9EZZzeFmvpv6mjiZgt
PEeMCQ+O+oh+ZtnwJfJY//E0rOJOq35X6zMgFJo9oQhjazI2JEG6wITHCSuCPZZ9ctN7yTP3itJe
sOFjkmovdAOKDt443GEhCV2rpkqwf5xWmcMbv/xPFaRXQe/fv8LLTIPV7F4frUmOFAMhNoKSva9s
RuFF/YANJRz/IubSENbN500YQgVaMOTj6TvHrbHQ/+vfNiBSwBoXFy27JVfWqdZwMdUV4vfEeAi2
8JgTyGaxfeCDIzlRqjvPvXIbn9EadPzZ/pUJBtc+Q0bmfe2fdSguLHF0tRjaHD00/9h1ypbnzluv
VSZM6yS3bS22jHoq9PgnVYVOa2/zK0gxtgjRvsTEXJqzspj5KfDOop5r4VO4unMg/CPuFvyZkYKM
T3zQEIORGD2EixDaGu4ZLcU0XbTZ5zjYgssgFRC/gLNIXHEnNJQGgx2m7wlfDLb6LtVMIXGvBCif
hrF2/oCJQXLRGg4iJewTQSs29QkP4zpB9aIREVhXUvL9kb+edpfT+HaxZZK/uwK4JpJhlEDb9A/i
bmy1o+rFcMY3t9ItReOam76rLLzo1od0WBa/CMH/5HgXWnUE37FYnvu1K9VTt8wdZwUZXXNxsqIw
hup48xDXObMFZVP0MoBxOQy0LAn/itpW/wzueLXlMqKNBxRvNZPE66ZAe8Odpnl/BZnoI5EtfNHW
w0O00l1eCs29mZkMXRNra0GejwqXLTqwigX31P42KwBreGldDf6KL+1cNsZTkPD3qLwt14+0LbWY
GofVRTpfUtm7x7KvlHdWaJJ1lhdpVsdIGZsxgpoLhuYMJwgkrmdQZVHezzl+sblze/EWeArBaFSi
nAbo0AtHPhSA+TrRi3KcBlEUdGXY+JPKpAXxJkC+44LQHtVODE4ouZYfKbmODVlGRv6gR/ijdBrd
Js2lQY+l5plgIAoDb9nLFcpZwX4iYYt9KdVjbzA5Of6/StS83NLW7/dXVs6kDKOyRbni6vaJ3dyG
eh/EckwL2Bk3Hs9xgk0Hss5JKMafOa+M3tPxmWFQ8s30eLcKxKGmBCnZ/oDdtaJjdRaBO9+UIG2i
1m4iy70FN4Vz+N7hR+KyrAVi4kO7mXzShALOVNOJt5FmD1OIubL/xrSZrxOUc6fs40zCKRI/HQio
aOdnt0Les1YBJnRx9Sfkzs+G/mdLn5ujaiq+dZAX2SBy4yqBUmBP3Ai3wdKefwumBOG5YlSVAt8B
pKSuih2vsCpxiAzCy15QG0H5vI9MmBoR/3RIesT2SE1umx4qc7sc+BJh6D3wGOZfg+j/z5Tc3olg
nwsHeR79+WTJf1apsO0b5W6BtLBImmPit+ASTyj/lemHIDaRBcmZQCMS/qpMODlNDvk4cfPIvTDV
pBSppWFo8HczO8UQnzJDbQR42nvoPySlPr7es54YKDnROKeIrEj1deN/pQHLrvDFO6CHGewaF8yy
sRNdqJFD0nJa2ue98BpZhlo+6gXR2OR+sU/L6vmqtTJxqM2Q5WhTah5PDAHmDyam8P9FIZWInWSI
R0Bf+VneERe8xKsEE0x2RiBLDqDKuChcLRM1SbEJBRQUDRsf5Cw3GUH2nFeZzfkP1RWxuXYWx1bx
dyeGxQTKnyX1kYkWjsbgCo9s3c+E6VuA9nJfEmyGgJQNQ2dfserZa/T25yHIBofCcDQbhbfWyx2Y
aUK0s5VoduXbenNq8E96BwFgGGVnwe++kW7ecwrd6ehp/2j4/G5PgjpSvHuufAu06UWpZFpf8/Fd
AkzT/jlT1vL8viJkBVxIwdVIfOLIjc3ZT/0LOfoAvCIjf6DsOkJRAS2aT2ZNrKXsuWgC7Q812DSP
YYSoftoWDPVUZjF3g8KXXpM/suBMYtsqLI3i/7xJWzrZsTGuW59jp42r8ruV+/RhSrBqgS2co9Mv
DFjr4XS8TJ2roxeZ9DGvlswr7r4YOoNU2CbjHbrhTY58ZPlPA4RhtZW+dSEjcvz0btLBQoE2D4+l
Cw609qRxkDR1An0rxuXqVhBe+z/e4RhH1FbEro0ME/CwZ8ANuolp+6Y9BAjs2aNW5CwNrlEgVSkW
ZO8Q6dt/BV1XIoQFY8kqRCYHvfD4MwvGyLMYgENeEPFQNwagKZthLWGoqqbHmWHhkCWgbTQKXbhw
r+fKFtKq+G969cIGw6WTx69QcEKhweQ+701MTPz6LrbEbCyIgRGpC5LYAqZqDrvccn5s7/LAV6Se
yZRqpZyA3y27+HpNtKTZSMLS1yavlzj3gEWwr/fXc2cVv8mU9W3ZveQ36xSqQUc30PlnL14dKkcY
tJM2bX3TRODAepHI7zadCTba5M0i/PxZB6A4gdV7xu5MtEy3p+rdsGU27osIEVj/RFJmeCFqi74p
DC15pUo3Mgxeth7pBymVM0J5ip21XeXSuVy722mmS6MfQOxjUGy6OeraK944R+U6E+XjCXOaqjOB
j9ulhPq1qvfKkVjB/Flhv+0gy+USCMCFhCrJnnHCeODTl0O3XXs2yDJf4lrs1we7LFkBaRL5flAY
zdkPRsS5pumqZLY4t72UhLvtSpM0OHI9nYgMT5+6agdTTrbF6s6T8Ey9mzWhiZ/z/zUtCRY6IzSB
Spoaq+8YkcbG3cwBGlBu3TxiiGPBpjjHuIf+q3Ly/RjjN+J0qmxBOhQ2HYE3y0Tv76GFMV9uaNBC
S+q4D5OnvbG2L0PR7X+zZUxwUsJsIl+3+36NhSuetQWtn5nmUeyyOmSUmfatKrcTHEM6AAd9jlm4
0l4vQyliNHJ4PXC6QEoBFkkGl5CO/IaBI22MvJ5tOHesTWC9RlQpBW9kVbmreeYucVs1kR9J/sIP
Ti+wOtvBaJfOMQMlHP+JZQ45pCyjs//WSlM7snCnHV7Bd2VT7T4NeMdNeleD5KJ+93Rvo5b36Bpd
NdZHo4bySTbNvdNMjUGth8YzrqNFevZkkInODYxUFIQbJTIIPbGzRu/nyoQUDmyP8bzGvpPB4Bn1
EqjsRkR00c8UyUzGGYuEgqi4jBe083SA1kOS8/omwVqNB8Fn2u5lQVga6Gzq6uQcuxXr3FK1WEWZ
VD9dfGutu7oO+SzZMKehemU3/9PFEUfGFbuhC7kHF+4ulUUYof1TMNN8mH4d+v3VtwT9+ZdjOx/E
se6cIOjBkR8xBvHeQq4tMhvMMtw4lstBDViDDQyvkZCDnVFKFpbEpsMo/JkYVxQr4LZHYchkEVyr
CStWZubjIYKtYc9RAi8zSHGK9/8djchwIfjq8IVsxh+Dhid6VrDAKwmzSW2ABg9p76xYmT1YkSkP
niVf3c3PCbK0i4v9aTNaARsshL0WzFBaKRdvgRQYVwWX7/Ebpt4KHkTwoKN5pJcX2DvfbXAvRVI8
S+maE62iPsf/vnKtVX8YMNwVL7ug6vudOyBvzXFtgLaQsbbQR7g8/NqCtPEH5xOWSLvqOjseRTZW
M8X17/NWbShYHfwOiNI9fwXM9sN0mG+tYGAieIkixJfPvmJTHVkBI1vP58BlXHks6g5U9/xTlcJm
NsYPrC2aZYZFYFkMX+2EjdtOkgnJ5TDnPeQsFoyPPuDDMcJ3m6EtQ9DPOO8A8RX1DNQscdhAOMhh
dXZJfg7ox5epqk+mBEwbIjSXTEuXLi/eL0wPoJQuKsUE1yFtR0UtcoyKq3HV7EY8t3J7076ny1eX
CzsGW68/kdphjOimEomDK1LMxvpXiC99nNmlBbXhpChBbxIFhQTe73pedR9GbGMcT1DYu4aibcdH
laXOtCsvRNZTLjaKwwn2o/j1EKGFbNn+JnWE2zE/0tGoIxQsiEtWCDs1lTVfaJpL/7pJ0M/wj0ay
zLGwbZ7aBsGXH89pA3m40+f3Dha6zeZ4B1xcOSoWicwc3pgdHWqHZSc43saqALbIvLRjmxZCyet0
y1cjZ5I8Dx9vLjiBvc8LXdtUkyr7H5TOFn3D+Oa/n+kzcWl1OlvF21zUAQiEQkGjhB0krnKJ1Zpr
mwZnPRFA3lfKB4IY1GBE58aQ3h3TfXYHYT0hJV3W5MTW8zqPa/EdVQQP6qUwmb1brmCMUx74RM83
DP45dL4Kvyy+xQUzC7ResOeKN65tXUkhxpWm4Bq2HNr80fNTthkvzu5COxv9uFfpL6ZRcG/LtMrN
xdy1E+LcUZboIUmAzmC5A962EAEGSQCQnnrHGlIl3WAo/3B4tpnv4r3it65sp2qcyTghlqO4lnAO
J2r3RZtuTz5VLoZQQuCodYw1zXPNSnKAm/kimzAob5aWgbH7Nd4hmoRVuW0LtwopDogXRaZ4Myp3
XOo85cBzOlufZVqqUtaK5tYJpBouKgMsQIie/yZcM7yo8iVyR2ZHNyO1P3YPtpsGGBfac0kgga15
eb8NC/oDrLTZovIyVv4Nwp2tqAkA04YINjYEj3fYezCiB1TMipLp8DZQTm46Tl9FKCiL8KTsqwd1
plDzPWaLE853+F9V4B/aNISTXBLXUrPIePdWGKv0/VbEwu52D+Odb3ho342enlxXm2RcruWAisoQ
yX6O6y9zkrzmB6s2SEYmXxnHQfB/rUjscigTPzJQkZ7SmNAI4Gt3X0raP2Nj+McKEBeyAa5Iin5g
gqeHXwl8cbdguiHCh5Bo1xsDRe2rcapvhoI3rn1sIbHKjKqCheNuuvfOb+2jEvKVjq52ZNQQ1Nn3
Ho94OVr1cSk8UcTkh/38eHea15sO9NnoMQ0fy2dsGsgVdxfsEE/0K27ZZF12VlNLGaTp5TLDbPru
MM4SQ05CLsHOjJQS+g8N0rLvBGfMVM6F5HBNLsmAWnWj/dtK1vP3WvOenBIoXAZWA0ptgEjs3dRz
rTAyVTy2wlpPiqahM0ZvEoyrTLSzE5pQYazCc4xysQcYWqrOStAOQ8IEDY+i7SJRJaNZINqWgThJ
SnshWP2Dc0n+jMdWQdfzAqcishKDKNlzk+coUl9AxDZdY5p/X7auBG9o5PHj7paD3UZbqDdQj6C2
ddbmOPgs+iMR+oQfig+2DIMeVBhjmnRHUZijdQnigXiyObeJ1GQUq4a5iJOXzC/ZZBIBM4IHrvNm
aOTXl3L4HKxmkC7kjqKSJZAdJSY3Iy2Kiqgx/9A1R4JO7xA8IZ2/mVc6KwpnNRfGFTOyJtno1qvL
DgVTZlX7a81i5RGSjy8x4fMajaeivAwyYLCg8Eqy9nBrG59nyS49LyBAMLAdw1ILy38DdDEBQUgO
GJ+LN3d536y2PksSIhgQXN0IkWispj+kRY0atr3Q8xbVDjMS9EdX0CZJ5uQYSTl0+6czVEb+SgJR
JDvdjxFfEV+3/TXG50Ts2upZNvfbAnKnzQdMl80wDGKDd9NfGGHyKR23/ct4yWCKLh6Ub2Tse4uc
OfcMYVSoxgjmwJJhMOWbTevbBSDgxvDlBYWfyp+F5FQnB7elK4fFaKvk+YC+L++Y9lRbMD8sk6WH
dAWw6GlJttTESaPK0vGtrUqg5yP8n9oovSqJMFW7i2hIAAES48yvpKKo7kbQ9kcu+nrL4mnTGpm2
SIM26Z6jYHSKGeI+/Q4i9hPwnHItyR6gtdLR8pbjFSYbfGA/qDZrXZNd600FpGHGETPAggESLeMF
2d93B3RxTtLMi2sISZTbzMVhIYIe+Z9x+ktSGTMHbvOMfAYoctmXjnO9pyVH1zQ8VnDymH4eeTSF
6Mth7RsKuv3fW5ZYzYQKoAT0tsNLVbJ8qRWwe2tl42caTSLs/jkfqw9dYjC5redD37jHga2ffZbG
w85T/MKK0CfxhpG4jFdfCAO/UYBfnng0x0U/hbUUMBTAiDLD3vGh97YSDAz89YzeVd2nuI/Eog8B
UGeFTsG4cgavU9tBbRhP27ea6jsPgcIqDrdN5+ZBCnondGPRyCycsR99pmV4ZST4yjPBCQurCGph
RusRCyNtRvjC/h36eOxVc+LvPDjjFZ4P4WBhWNug6iGFx9/PJ2mZ/WgNlkiImHCSDW8Bmsf3QBmr
CCyNa0Q70k19N/6yzej8lnAYWH5Lo44Awt4KstYT+kfWjwn7EBL7jtp6iLnCt2oIxiM60OEVkkkP
BUcSi4H0w4D57z/sLWyK3x3zlEYXj1qJk9S4p44yKp5P6RSFWXX0nd4nzRsdko/3IM2rCL7GA/yv
n4DWYxyiFBMCpmjh6GFi0fwWB0BzBRTyfM9bCS+UNeymmqGDjF47zutmzDC2iWMvcyrHe6pDF2Py
BAXZxrKbwer+LqNHMrEPomoWhcGxJxhVePj61hNXk9jzGrEJEynYG6sAURxCQ5y0N9ldhAJVKv43
FYcRcAERuXkVY8lk16Y1wGmp+OGPU1gtIPPOUaRxbcmZjBXjBQmWCcU6vn951mfux7LCBR+IFyD6
DzrgVNTs06WH+qOaW0V3zzDcwKv7gR/aPr4yE7fLQa52dbN7kbASO7YcRiH4DjFfqPOEripjfCHX
U/CsChvAQAvRIglr3KbDObGWVuRZ+iEzEPYZH8vNHKugJ2KOL9QKgEIy0ziT4Qvyz7UlJnj0T69/
ITv7oFs5ZRbfUreiRh9m55LD53VG7HWmFTnIdCkURxIZCP77rLiBc64lJVTKR0h/voeIKLZZ9d1q
0FXjLfnB+GZshsmQAJYdEtQhQg78C5JftvaeCLMW5bIFKkQZ0c2mcEunbmKYaWcwQh4CvTrAsAUj
fgcKf1capeTj8BL5ZQniJy5Glf9Tnil9YXiysmDNKPcKhnl/0zko9gzHrYeIVksykJ5HKlGVNJ29
DxkXFKRp+q1C3aZhuF/vx/q1FYgDqqAZkxC5g7wRMxhEM5DdzCYi23/8g+28FUdgsIBfsYWX8KO2
yaqDqEmX6qnR6hwddxHRICwpFq8jaAFlR/DJNG7gpTo6Bi5dIdqmH1oqE7r5+3dCG93N1+UCewuF
IRN90f/hFGRnOncgPjX/+qTPWaEW2b1fCC93t97nDqpmlqRAVpRjAlcHSQ+pCs1Xn6mUrV67pHp2
c/VCDGx8Zx+xUQXJ0KfsUbxeu5iExj9M2BLZH9oY5ZyQeaDn6tX1kIyi8Uqr0NClWM5nLO1z7vLt
E0hBGlSrXVPrRyIlqPw+CXpm1GY/DLIfiNS11LbwXI6CsNRhr74IOj1lrlbGY4lkElCFbsrDuyd2
0oldAfQqa1DH4HfnZi5OgU2Cror0KXKItsnjGJEoyuy1gTJgU71tEftWShgpXgfEIvpQ6aaf0a7n
L36IaMmtjWXT4SeK93Bug3Gm2WnaSBkV2VdYF9kmpvaHC/tiQqDW+Upe+z7WMvo0/kbty7UZ9gj4
rUVheM5aEAZTxNWgXkh8vwViYPWZbfjRf/6u749vfpcHnEpWoD4XxnrefyZWSgdoESQLsfb9ImrF
LrJTHH+sN9r64WHe7SH1C2ZSZV44SbzEvXmS4r0DYy/fSHVBpHQ75LYOU88gjONICazQSvcWxSqL
iTD/RdorFYn5PJE+k8h/wHsEf47nacq1Gf4CbUzCpPJryUf+jBLFpd6glM07lVFc1pJCmbvD7dpc
/KJmvMQZAJSm8/4l4uVcGgCr0kWadBu8EzAgXxDSpykFP88KmJoX3u7BJ0+uHhTbbU7SC/B0h7yT
c+cxTbyrJpsT2GfmBzmCQDGjlXwRJTI9XlVHXyGLRfAuPPzksmdVzWBs/EnWKE863gjPpX4524fp
UTnTvlBt3L0kIdYQxFu6ZId92n8KYFb7aHyPR26F+USHZP+j0gwHhW6/SqSApCjxnA27/DZxoZcE
zXOgVi4Edqq7AQ6c9d4CQ6Wxfwk+qH3PQkn5cls/P2IGPZLVa3xsTgMaplT0AvXkjQ8SMbpu6vNs
jI31zSghwCifWDlKytuODRkY05FOP83NXiLBBKm4+oY2sSedXpogfXk5ZFR0iCwjX1TcCm9LMqLD
F0uLvPM4QHkeoZWvsP12P7gIAWAiqz/F5h+VGCaUb3U78u4GWQF79F9b9bRpGPMrSGUmKCLjeLHn
7uYXs5fwH8TFc63HhNMjQoxj8bd5BVdc7NwAO+oqH+NLoUiUfaPJtQhgfvfBrOotc0YHaN+V/byT
PiYXvs+Bz+YjRquWheFCwCfJzAGVz+ydB7cyS5S/9mJdwTh3nWbMQggz20nEFkuAGdDV4YsHv9kR
0MjXviDkbVEZSVIqBaOZJX7tjzIPiorAC6tfhWIKa1zoVHUL1lgXbL4NJ7tq98RMlIdNdZ0ACusU
sNxIY9C4X+cYlWTQm6JnB5O1Rw5TSRqRuiHLB+RyJIjC46sILD4VGPwmLel+TQJFFMl/mbWaIruF
J2M5+7u7pPIC/m/XDjxix3nFz3cgIooQAy7LvqykaaWYH6EMULBG0K8RizG9vcS0ZCUhwBaFRGus
ceDP2O3e0HdTurl7OivwA49Nd/rrSQpgI5NQVRuLY+8MNuxBqCYkdr7vDBpA7yEDMwC5whc/YLd+
jjC3VBzD9ZtqEx70g5rlX4TuAqut64RAiOB2GxAaft0HOBjEPY8c/vE+jM5+++xSrgM5Ux/opO7D
oPvZ6tpozCT4zjqGjtnxEYSDv/h2kk+pmWukBZyhQ4sKXllzuZk1XKmKLV0dcp7qNMCWANo3q5dg
YMld5CE1IMKO3KVaOhV+FkWL97Rxg3lrOZersIWT5O1tqNDsJkDF/HMRSl+prgnEn7O2E1t9V0IU
kYN3kcTk3ZsoDDfTmYD6C4QGB7sf/6MvZbtCmvcO7ENLXRy35dcM+rJUXdw7L0WIa59LmPH4zjbw
+f6Fu7+zdj3GuUHgFhrFn1EWZM6Z4AIHjpPkX9Aaor2zwN9xowW9sLKdPlVz5s9ZsbbvFu9I94d9
6f7Af5D5lw4hH+HupBWiacwO+kGqf6sPwuVkabpJPpW0M2p/qVq/F+xrNutG4O6shaV8qvtgafo6
NxcOoqXKUB0a7e9gWWTrnRtbyFsAFhMPigCredpf4oLaBPZ7T98hW38vDXX5N6ILur6kVqBCCW9Q
km/BEo0+8VP1Tr5EhWqIWGhCze5KWmCkNfVgqCioK1Lik9Z+H2BJDxdhLC/xrgrjF+hR1JiYwmRd
OezKrI8LAEgK1Uv5dUpr0CudObhRn3D355zSzLDZI2UKyvjtz2SqHm81d2XhScCiDCYWlswE6m7a
Uz36UAQcmbmmCkLSeDlEATEA1lreqPmbAm+nsAU+AED6N9pqw9PiBHYx/tzWr0TMX+71a8SAwPiH
7Y4ii6Hcz50msf0biZ2vk8qybUF6eh16YeI6sejiZHUN+5chyiSygrL0Ok8niEe2LUARckSATpvk
RLdT/6bU/4mKnEu749bk7X9AGq9dvz1VDYJ46EYf6WDrO6cjRTinoVI5O1hCWVWcaZeHA3ZxHZcF
6kguO7Z3Jezo5nxXfJdBweWdlijfebf4Z+v90VLYlVjBperxxdqIFotFjFlldcZnikWKqmz0LCmM
2ykelkSW8GZEit6JrBzQZJhjNzPHHtLSeW7aNX2V7sINF1WIp8yyyZt9FFn/taJXAvw6HnFvWDgV
Hi9oJnkA0BB5WW3Cqv3aUTFA5hdtWvYmVa9UcCWub/9nyG9Qs2aREoTW4bIc8vaKgOQv2NpD2RrB
oCJDxaTc+bkeCqwdl3vrXhfPE+7qGFXZtTIOGplDLKUUqJMhXHWyjEDLpfKeHGAw+5+2x8+tG51P
2aw1pUbfddNej3IHZzh99mG4WF/4UD8IqkkgSN4ANYAygZmfvqB2uv91FRzdNAAZkhOlzvZ9TSpD
52E0aj55Pmjg/2+Nisk+nq1D3LkdTRSdIWPMHXEslu02j/eck0DTIIbcDIzs6IzntQPJ8HsD4F2U
zQikF3EmTIijm63nf75KJcbKHJPCnVq1d83Y4jcrmxWlwewD6VrbzESk/XRjR02dx7Di4DCM00pl
amoyHJs3bU64Apmpzfn9AZP8M/VHj0qEZhf2w5Qe1hEogj9niD8NEtMBET5GZQx8XoMDgw9UiTDo
bnvlKfjrZeHPuZoVyWDTLDy0ZuLcFeOFnongWGyJ4nK2MZW1RTRfLWsr8nqIFwwLFZei1sbI2z9R
bHyxQz74xpdzc3lupIga9FtD3VyOHbrYR9dytCkYm44ur9wHkd9IUeKG7jAcvmShNEj1ksRjwgPF
vumZhpAfjv0X48+p26s3AyksA/TxKfPNr3JiMaVobYM/1ZLcOD8lu7QpxUEGMkU5G9k2G1rxg+w7
nsEUU1zThBYXBHYsFBJULpGly2zlgLQ2Cs8lJjzq4rcN7rkzG66aNuJhs7y57g+JUvSRoDkVanJu
HCEi+vw7nArB54TqL9L8acV23bt2FnGeeluv7DwUS7Ipjpb5yF2Kzo/lKXZeeISdAEaoP7R3Enyq
BS7xpgUe74yzfrANcnJHS66DWlSm4DRs5y9o+kY1QrF/lt1Dr/ZLpX0VZdXnzJbQlF3oRrtOB/H6
ccuphlPKO17teBiioADB84VSR3kc2MDukYgIh8g0OfpmS/TGHs82JY9eP+tuHZCOpk44nJsqWfQ6
V5UYoJQDOQdjN8BE29wEcsFQFNtWY7DIZEUQ1NIuaMp9r7jWVpSvKtfKmEEx7l/H827YanmjcVri
yuRGICnw/18/8BmHpbJY7I4Bmvbq7m2iIo2E+fcOOrzhFmr5IFQAEg0FOwaQJbZi0liad2QFV/Ys
uz1zhpYprx0uLQnYwHk+WXPXveeJ2ggKg5613okHo1jM2sv7lsw/R/Jv6rNnNuC6aQh8QYUU1FUr
WqZpUU4WKfwCbBeL64dBFj3HiSMUo1u4ZoLw84/JhiTZ+t2jcNE4THo/H+AtGLysQHE2NyOlo/H7
igj4yMvGXQsBZPpBw5/uP9ajYBuJuklAxNZhPCKe7dq/FOVFwF+ZHnhdKXA8U+LtYpji7/u/dQ9y
U3Nync/Sgxs9+G3fqeCeytQnfVQHc3h/mDAc6tYWnXqJa3pwPgeg2SwnIA1ae08fTkbz7ZBVETTo
GTlMC2Dxn+I9NObQ9yIGW+sTnMqQmPzQP/Fgh8Imcg/ipIFnoo2gj4PTfLMzm0x2OeVejOByJY7Q
CcC3XR7vp5nH/1R7dy8QjlvLilMxkd4ctJFBmd7BDP04ZNLH8S4gKK76Acc5+EwnPyQ0L1GEgFdX
DiJtt/gZqPRaiT+5EDp2OYMGQ+w1cYFRAt5pG7/DBGpx6upgJRGLIsIZwQmrYlh6MGxPTTNGdZhY
DdcpFLUtOvHGsA4K6mUdzpLGdpl8CNYitfRLsWPMdnq5gGA8LIchkQz0+YBRx+D5Bg0pjihKIlbk
0ewEQwDzqdiv72W4nT7mmh+KOLtwgA7QUpAmRFx/RDnirILhARnxZCw9BRoss35aNUUyFjBFbAeT
P83JfZ62vMrwb6qy0U1rY8ne05PYQMODOA1eUq8f4kZivqTnmh09D0k1yADEMeb6C1TMlne75/P5
30tZN1PsKR84GbFDxGZt+aei44yBuQKMflUNFzQOUgnu/gFdAz085M7q8wkkORwP6n1QkW8Jia+O
sugxMOz14hhWZ1giNQQX5C3oSc5pHkfxwmQSzo7Rp4182hBk8M9gRoRGPHaCSnnq2CPbnZFyrxbe
Pd9qQaZDnwgsdn6xLKoZPaqnNs5pmXKy73f22LqTm1Uy567uUMZK7xIUbvGxCDahEHciZ4b6Decp
WmmVUw3ucWAlDpv15cB/zvYdIdRqoac2oCzAQFFRYJg6OtpxYRzi2Ra52NH1FKEgzxX3Wm/VnaOf
bEoEhW59v3fXnV2OfLjo0lFYNnhQgKtgg9DrW1sEpqprpEmA/OPPM+ogmrGtSMK3QFmJ2u8xhADE
V7Al4ptjIsNgi3MtGcOnn58sq32JiF3j4q7aI58i7/m+qKQcC3MzLoq/Vk6w0QKiVqr2VvVE8teA
lWtUXdygADgjwtJmh8B4ZAggI15f0ioQq0HhYs/41JTKkFM/VDhdTPT69k5pliXwu5m4lxybM90T
mdrBbQNRKkYNOn7BtpHcABVhqK+snDMUCarQcflMCsoquS0o2x04RRugBsteyX72XjsI8KzwB403
pqXXX5ZhyWWXdAQ7qo2pgsewpIWc5LV6IhHcoi98jmDB7oY+QO3HNgS/pBYCcdtN1NNmzQQ+uAak
jAunp2HpJBd51NrtL4UdkN9GQbxfuHe+z8KmdzK1uOelacFy/Yf/+6o/VRUPqJ3DsnzIEL8h12Nc
NNPYDTddbSGR9RUOZ9n8qCD50Jv4J2pbVY+Ypa1Gb3418+X0G2zYZLioheQmIsiNTq2dCYUyEBcA
XAvpjKJWjrS2hq6RP0Cvuco0AAwzBcl+e3/OAGG7qLB6lTAv4A+cUDnP4sKbv+5nXJpHsywc1TIT
rCZYKd1Pv2jBSbcuPJzXFek9qE6ACgvjLQa4SadnDR1uS/7uzEz+QTvutIb/3Hb9npHBmj1+MxH9
qtUzZYij50C+T2aioq7uVxyhvcTKovtr/ccsw8p5KboARwDnJIToDpN3CbmGd4qsILnW9YcGd4Au
T9KwBDeiPbbyqL7JEv61u7M+PFQN5QdzfjlClpKlJzh58e4nkYJrRFtNcto5z7ZF0ZGQRC8OoJo8
GfW9Hg24VAhqIYUlhrLbaG6bAekpj8CI48iXKMLwf71TT4JfT4P9Q/omiVEHpf6gmQpzJHNcw+DK
TmgqOiUKMfFJ/xzovxVzhP1e6bK6l2MZiRIjLaoffL4DxPJvTe1m+lGI1V7SCED1bllzlLYNxy3V
YZnSIupZ0/04Woc4XED5YaF33xTH8xryxdQJdGvlpo1lVyOs3MLWo/x/mhPOVk0Fdz9GAWOKuxjE
LBhrmu15SO4MLuGFegooIZ9mIXooAtHBm2+zmdXqxDcBZxQ79NyJqrbHGZeAmKh8nVmgd+Dew9UT
8BvD3IPJZgpLzIrI/vSdorC2duJ/ZHWefXAAFEujBVhm0fchD0Q1Hg1f965ydAjITqk+iQrPgNz9
WNrlV5R4I0XNAjDLaV0L4YmC1fUhJvnTg9Hk2lJqt8iTE2OeA/9mVd9xqd+5onTJQRZgsnGq49T+
Eta83YnU1k7tYhgLHGoSs8KjwSsh3wgATOENZ8m1WI2E8A+Q7+bVZ21YyoHxei/YNwKdO4rWuiQE
sCEDdy8jvo6AIEgqnPVJDBKEeq9UDOJMx22mJw/x8QIp4MZts0JMbkg6aaWfLqZDuSWh3S69uQy6
KHjefi7ny7bvxAOAVpSwYGSloBRwpPByx+xofO2n+MNwiiMoQJ9D8XLS4GO/6CLdrONSVg27ixpr
NA62BF76BdNjAym8kr79pge6V1xK78xFsqqEEpueE3u8V9+9SRjQZ03f8WXYCqfoZpErn9q6KWTU
5QYYYFAUBEBlDk8ZFbxoiweqmN7LkDfKo8Ax3c0HFD1so0L1B5NfiaWCbvbN/a3HMEOzSHzZyA2Z
qcT4VlxOmOCIdTFWM1tKKuC69n0F+tTcWMUIyYJT2AA+GVesl7LLas/CBcol1mhVY6HgVzIm44fX
QMdUaG4/dMnXX+/3FD/1QkB5eUvv2XbVqhavQ+lzqDaaoIHLqpSElLC6x3RfFAGuRjHolxob9nTy
QAVKLzFvGGvwCC5aLjHP/aNh+kkf0DnsD9FmKz6sCl7iRw27L+KgszgNyWinH+teeY0p6QrpgE78
ZJ2iB7n87t6DhTxCZwnsF+JywEBsptbGatAv+Yp2m10hFWWZcR7+H+kuMYV/4dyYBQWMh17wU9EI
O/2P2ruHe4gwbKVsHyIqLRJXiClpKy7GdCRfieybIwd0LaRmkaqTO6HNAVxjYQrDbEj9ZuztWZNS
Gg3CBE+3LAT0etSFSqllIwTms3CDRXzEgdTltYF6xr6GfFtZVg016C7XuvDKrBSOBwVdnSMCxrUn
3IrIuHotxwybh3mmNPbAZJKudBttDQ+ZvPaFKqPiJOZv7wvE+dzmFML0IuP+75ZRB7ZjERidhExX
PkJWLmTW8k372RIthVVyq7KOA4qaduqqHAxlPq8EvJCYe43wyBWaTtaSgtkuQqiiSqrMurvTpEPd
+unIpjKJGMmqPIct7VXuQotkyu4GpcD7FqXeAQzfHl1gSOpEl/ScN/V8o9hB+MVSTiHNt9A1J1Vz
S4VhTjM00PXIoiPHw1vaG+qt4lYlnhllb6VCSvew4mYgXed7aS82ELpB49V2FGNk+Na4/W4+Wxln
sZQUgoMRo9kAZGII/2HGJtmfolTN+80GUxt97kWbP4LLhrj30mtRuK6dT4P/YvW9BWgv4Lkq4sig
2CCuGc7DQE0CXe0vIVsnIzLRHtOzsS4CgXrAO1NPzoZIPiFeu9XqjMXSUrO4is5KGeeNJXegln5h
g0XfL2axzNI4XNbs4ECgP4n2TRSQy7hRHV30QmbjEJ2wHNW42gS5cZjOdgIQl+VbZ80/EQQ4S97h
YlmGZCP8xvu1gy6g9h2vr3kyX7BmVpr+rWyDjFZ5OTtI6z0/neQw1BVTOax37mHDvvXJGCV3GQMR
F7yD4qndYbudAqq4OgwX0yNaDsKfOb3L9/Cw4piRF2+GN9EDntHni/msxFT2aWeTEtHXRpwUOOil
NRgMzbSPBOuwg3AZoxfI/UHmpVkwhBwz58UvesvHReMfFrIPFvOlDDVbN3qxrEfXJDo4QIXMJ4Jx
93y33oD6Y3gx0Xtm98vTGE77DukjZFa5Gk6XEhDq4SnTTzo4EcToJmVAFi/Bas5VAd/ICouzyBtJ
MbMs2wKvmLGCIQzrCgLkxcC2Q50MIWpsBjqWft5olRZ8AthI8u+BaPTH7/FLM+fB3jdc3s+bD82K
MHn0Rej5YX3dvAE6OrfGiH/UEndpypRcK4aih6xyNJxqp8MkD8sdojrEHocHt3LRXKFTqRFSFsnI
reoudPhmAvZH+Mcgs7G/18EKsGa/rUbbWtlBaMDGcOBuc89gjepzD9jfl8mO2vB1q+jI+iFUu1hK
6JjPogS8z5q9mnMsZpajqVQd54Yg9hktQfOw6sp7cQvhk/bvWuxdxoCJmxdLcnwp+9D9p2smN0//
y1IrTufhUPWS3riJpDNCVqSlgXxUOQtjMG6ooJ80SN7S1KSGIzb04SvFD+5lCED1Nqta1Gx7XA3k
fE1Xu3Or0CttIuHmc8RrOb4ZheizcWHMAtGGdMHtiF+Y6G+ksXcXv2X1VgdeA9N0VMZwCz7oSuB9
itz/L+UyZhxXuhXu5HPiKS9K0aYox36XwVWWhrLbJen9bM2HI8BEAqKkDz+Y+IPJanKOSOzhV6WS
6C9McyP/x6VYjG88vPqKFdJ6KdiIWIRY37n5SWNLJPv7Fv5cnmJ312oALy+BMptK7TZFoLbsa+7E
PpXbaqP7U7y4lYxQq4pFuRv5BgBc166FviEvKfV9e+qI8CR1dv4jud8pNkjrl1vFqTTgx/NM40lu
1YW+Y6dx823ulED1GPDbFp58cC43hu3LEhZ3euoheHp6db5yirN/gFT+9ooEmWk2KWiRrNCC+R42
3yWgMfV6LGKA4u2diO5UfaXQ3Gc0PX3CUTx4+8+W2TWYz1EtEw6eICYh1wUI6ulrdCjbrLPvUePT
u6uJGlcGiYHvwnYRhBo3F+wlqeruXjXwB/NjQ6nTht5YXJ4NjyUiMfVYaTlAAANDdTd7j2rLa3K3
RGzo2ELWolF+kFZbQw888Zs49vGUFz5LmDGWbGanvbzC+zb0ROhe7Zi4u1sQfL3eI0SWnzPyP6yz
mEnn79pwbOpO24tm/ptSyT/JnXHPAl7LhSvrkItR6TFKAa76YKhIZSSLU19qZQlsP62LVu/dvSdM
54ERsriISoYCXMsmJvJuRq5LQTtYFLDUPIivA1FRPVBSMzdinkeZog/zmwLS+c+aOuP064VO3aHr
0lYsFkyApbYMZ38SctG9foXYXlX2yMDhK4lWjcScOZk2SVbazIZQ/8X1ARMirCBxfxyC011EN4nV
H+w5PpEX7d1aKJufos21HMp1xJNk+q3ya3rV0pMJPPuNe4A/ylzNAy42XCDdJAUAnEofOYa1rXCq
PrW1qJDvi+ZeO/RjlbmsdvwrHbR1nhdATJ9V/DRWHCXtUO5j0ENmhoM2uawuSBB/rXV3TzZwqLEE
FmnHLUXjNFRrHDpKq5bK2TU0gaSR7ptk3SimOPoNg0p/SCZb8tWqDqXr6MCjmSgtalLO+j2icjXW
qmmW+TcI3BVCRm2Ckf1G8qesWxkRPn1xCYd618RzJlkNEm59gESGeqsVvS3u8GhQqjgIpUQYlWkf
XE/NnU0UPg0NiH29BK1g1K2P4FD0G7TjbRiytInn3xqgH2FPmhty5gpVbJGQJ8lqZQUZQIgO81Qd
l7Zwud/treNpKvKSJwRRQPfB2l/1LXG44RPPWNLCE9wY5vwSCDl2MnYJbIK1/LV7lPYpx6v87KIY
vH0VJyZ3kLNbYwT6MoxA7I6MVz3abAoCSHa5uCHGVin2C3FwQ9Op7XvTHC/FGGHbb1gQVxg/YLTr
YFLjO+8eqM+TfjY5eo4lZ3Zlwo4VNH7xd546fNrhWh6bPFi4ycIaKCU4NxL8FJmuQGhqpSC4zRNo
1QaRzZtfnKsGmnmk/ajtUsID2etUaq16YxTRJbNf+8R4hiX9RPHUfrHxKR9OrGJgC71PiCCPHdw7
rkaamRWZ5B08AsB+pq474cdiWeTSIv+Tg37di4mD/AE/QSp3EohSakm6YyEmHclzTykT0Uf+d1OP
o1EQqPlzcXrhPW3CqXvKySwJe7fMSGnYY8sqRwWlc4elv8tZAi9LaHJdl3UiiLp0TjZFBC417smb
Hs2tLpbmObg65VcuoB0j/jgEaRozjW7t+FIecuuMM07h9QbjLHAd95DzVs4D+FE4DymypMt9uvyy
0U3hKOggyhguwu/KBoCS2djxHr0Cv8ePG+N53OU/pXKYHCniMFFsEnE7S99tqFjkLvlhTaMwX1xj
2XjWYrzCRFw9n1TEbgayGZpkOE9qpU8c1y0yG/vSs5HzclJ4pih5CdNq7iaqjBh2jYoVllD3OOLX
Gc5yKe974rDkbJUJRrHyEZiiURBD1iCDCUo5JSYyPB4Xz3BIEI5ITDVUnK+Qti5xEJOhd+tTj1G7
dvXG8fVINtVuNAb4rISyIQoPMnGaLL2QdL+1D8osePiMqzN/d7BTd7bvYurB8LXskwvYpovGtyo3
PjOSNXhCoPipjgvQ5SVOjDTiFO7TtQVwJ+77XdXwYo6Jek0y5unEdSZPUPy4tDbLq4oUuMSiveYY
e/mwopXHxmU/B+wwHtc907N7acftBjULgokV9A0JLEqRq4HMieMcbkwnPOP/MXBXXnvQPrF1xGKM
1g2KKy19zarQsgIx/bdFUblKTY2N3DPPmNnuaMA38EYO/6XOwp8VsW9Ivwj19y67LCQkSdOpJ3B3
wsF9Z+28mYjJqO7vCk+Z8f/6H+XJrw4fnbJBc8B+UsW+fjZkAwPTI4AZ0vGehfB2HPbux7xZ5zs3
7fSNZriBOwtUQuwXYZlp0XDpQOYWn/piFCAgu70o/I9J/VdRUz/tAfKeVO++fPySESwlz+eaew8v
6ZAIUWeU08b0ySInz/711L0sIYV9S35jMqE8YX+Hr0PgYptM5MstXd2GjqoC0JN8JC2tDQYQfY3D
8aKO9+4z+wQOc5fsEpIdiNlr6i6KRlHgot2wAXgZSHbGI4DaGowLUw4BJlt2be/ddZVjGKULDpST
rW3XrnShyJg7Gn9WOodG0U0ENudTJHzl6fm8KplZZ4OAAKD77b2hnCa2jXX7O4eM1OQLEAPY4t5B
eicAX8dP2uJDcZjJ1frDbM4z9D/p96gE2WcvGyAaue3KPOEHVwsaKu5RGSJkJyfLTXdIPBBUFPAw
hlTHKPSUoazzGsOFgxDCka4Jvs1y7J3ntB2i+VhtBds5w3rHjIxdwZlxPKbuJcNWP6ce7MUBNsYU
+covNmnA9zZ5I8PI/UvN/RKxIKbgv35105t4wZlecoPvHO/S70hjRdtscmHiy4JbeffRjLmQ7lkO
ovKMVqmc6GLFC9MnPoss08dDFITWm6m+yQWR+Lr4gXPyn7zJ2NNs9jiOZo3tpPtqtdGQxmRA1D5d
Jjkyqpdqk4g1sfvx4mpw+W6PXWVKU09fGkpPXXRLs9YU1htpo3FbH6h/NE10rDS/tHqwVL3L66Yn
GptQNXOFeidNT0mggGachMjeQM7IgKYqKzvcuBVk7b+TckgLJejRllNU8ouSlzRWmRY/HynaZqo2
oWSs0V6pmTKHUDyiM26siQC71CEmEAMnay8OPPZbSynn/aVV+SITWMAXr6qwmfA6L0eyyBwZBLEF
P2d3pe0cMsxpcGebp3BshJOOl/VJ0Mm1seIqp1Cc8dhJgs/oyHXmmwufqJmd6MzySz1fEXStk1BB
xT594MCITy486iqlAKGgubkosOi3ZFQkqfk1Y0LToj4xphUzOK6QEg/PYWWsZVjTdhpDqZcF2n1s
7Jnsc83UJ1ovg1ewztxHPOOLKZxK8yEY6WS9fvSY8wLKxjiBYGxdCoqa/g9c0798iGSBfs4wjMFr
zyvljGfY1EtugHEwnN6jbKmspBM6kUPgnooe9dhlCopOgRAEP3N3OqaBf+DNthp0z37Y6H/TQ5Wt
7jcsNbgr5BxFUUlbBYGhGiCcpTptyOlPztdBLv6JfMiG/cT9VrL7nEWfV/cIL2W78PDzUFgFJDp8
JjBbjuFqLVyP3h5wRz+YGdu2s+fMf+l3fJulxrvOM9B6Jy+kGHUmcaLkiiWGgniVVCY+S5V4ws6s
/6z/k0bgx5M8knACDv+OajhRJmQp6UMJ5Hip9T+8gQ4RZxcnuFDyyXnfH4Q/n6gI7WG1ITHszDpU
dIdZsPUm2+KBLA4Z+Koz9fVGx1BG4fHLmv//bexnzFq8zSpPrJ57CUO25TxFysJNWjFJoWOsB7D0
8h7NQWecf3H67oqum9mHBvFto/lL7JNtrkJW6+f6FCw9UuC1RuLO/FsLhTM9lo+2vZCt9Ul40l+l
31iP3JjJ8HrjXaYR3RaB3wMZlvPJz10kBTKwgipX+4+Wo5Km7kbFFGWZz/kOOGh4aPg4+yowP2u9
8eRpTOiQga9kutRuRTuCGPGHTj5LiygM8DhtP2mx93Y4iQcN58OpjHAjYVFcNEHI4Y/8Xnj0xw2b
4+vNnTCxMeFONqkCesJBTXhA5R5d78dHyOGICArpjSQdhpW29KVqX1PQkhWcsWm26q6x4J8EHM0q
vRbI/WiDnQeMkA/+55Uktm3VhyByyBO131xG3SQX9weAcc+CB/riumSGb6WJODekGCTXtioCI8Mm
fngwPV7YPF4g+aCrphSY+RQ8DIuDcIFM3kkacXitD4md/lryuuBVfxtjx0nVP/i2CoUnPkDEO3mU
QCdSlah2Jys9FJR+9eqMqTh1JQFTa71g8z7n0BF79jyCSGMJEHaPRJmwI32Mvois9DhVLIKz3XlB
qRbtaVFpXaIzFp4HY9tsjmWUhv3JUUtNSSRUahqU/fNI6IoAYwvXAptXKuCbT3SoyUwpvFhbp/Xq
v9hwgu6yckcLY+icQ43F+QTJtwK5bdKLfMEolzJRY9VSRatpeFoAMlK46iM+rn0Jt6AK86X5HPYU
8JHBTN9l/MUpMsFkr5JTWky/FNSaOPUbO3+oNcLYVtJEVQrp9Spcwq+aVYp28aWY3XrHC5FdIV9E
c16UZYLr3tJL1DVgKR4lRZZpbrBzO5xMQpWKutmIPvuJeGgAJyx71D0PGm0WRoXm0V62UnBNo4Ld
iFJHBoIdxAyH+ol6CdEB6126abE2JYkTaR5LD19J/vv2WtniNTy/UJ4EigABG+BDKXMARw8OV4sk
V4AcX9sQT01y/7PTGaG6cCXK1A8jAdC4vRazaDcEjgesdGo4dPFYzbjexThS9dfUbR/RrKw++vcG
wrzk6i+xomdGEf+s1FqfX7hvCvF1EiumqgFJMH1KvTCQZV+rm3XVGEKB2+DbyrBioYwVFIad0RHo
qDjnEZzCC0IGdiRKcdUvqF1F4UlrP8Ks8bTXeASOqpFoFBhd2R9Cp5c4U3pQoE8fvCPX6XhvQVVV
ZmecMJ38CQRv9psbzOkpPf+VFI3PudO6YPPCR2lPyoRRiyhfeqIr/INja3UoMy7LnFrQdHaAcueM
IX59nINjk4+0dewF3XNKXMVa6hPPUHUB8MIMo8Vb07GfoOBt3Js82UjJaXE8zHkFqVnZ6iN6ihg0
X1GJUBWqs0lc6xSAUfihyYv2Mb+VtKOxwk+nOVWw/6VZIn436TrIcyj8+ci+cU0Seg5mpb9CJtu2
/9S+GAcuiLTY7QWnNxqpvTPs0KF8h3SNSVVcGIBN6e3d7Y+16AB9CNsZHJ1cH4uZQlY6bx/GUCzH
MJ+bY7NpWmdz/0br/LsNNeRoJZ8kYjKUACRTOiZXraRXcrZlaEnZYdLcS8XATF2PdDhCIjMinOQH
TM8ittqJK8gW6KKq9WAHXrRRu+y64nSEfAiX43eVxpybBVAT6mRngQYwT/pv9fcjh2fJMcOTRS0E
GLrNRAzclCQvGc7hqPr6F9t3sQnfJk4lQ1cne8eNUWX4VkBovROo7fTNKwVlxBUgT+IGK7rlwC4F
XT09O52/7U7h5NUiAs0Ta0zigsCbuoGQ0mMBA9BNWI1QN0aP505+4TN0pya+PCHnx0o72M5DaB6r
eRio0C1P/JSigrLZw9QZp1abJpsUXVP71TKQ7WSO49xBSZbrXO6up3T0uU98emqCckOInBaGthy6
NEwyaqOJFy3irF4qdDQ7QZqw4YvTrk2uoVQLjiiDKIeZvw3/xmZ7dV56ozTiC61PK80QvGYohSao
842VRCFNqZqb7yQeoP/fs2q5uPZ2ngKfZ1WI36VoAih8P/a2g6Zdqfx2zT9uPD391zuJPniYPrjB
wDQPT14MasTHjXEN2H1w3/+ey3HqaB7o1A+IQIlThozSeq0xdojYEy42V54tRj4oSf5pgkAfRIQ2
CQw8Xqrt9aqQubRjYaL2IsZ/Q6LLPYGgOOdtLDcF3lN1UiKnZ072JFDf7wQY5wYHM6x0+plxQbBO
yZCteRl1o+fOM2IGSLvtxCDrlK7QcxsSrfpmy8fypgC6DfM3aUATk4VuZ5ue/BWIn93ClQ91MJbB
zFRD5Pjmj8uJqgsVoqLUtyPw+ClkLUwGf4y3Cm2MTC81Ie1RjnkXpfPHLqEgLiacpT7HyKjsVhu9
u4e0+KSY1dZzStV6ybR3CorJu8CwJgjhdl0Y0y5tcAMI90WSI9DeOZbeXxkcLzpGDtgIx57fvFwy
Of2571/78id2YU9XUUfo04O3Bds64NCTVg8Iq2fyiwwLOSynwDv6bVth6qh+qI/mycpidbR/cLwj
E4AWrRAOT2muNUfH9cG5p9Vnw72/ZXaBaCEzMkWOLmY6ljo63iF1X6Hn3kveaRYy6ZIi1yLhyCtg
OtYFGqymxRvEMrb4tmP1kjA/7Fzk2Ahz5NwwDp88Vi2wBlOmSwG31malgjT8OhKIrue1fD/CMU30
BMnobs85sSSNuLvGD7N3HprfMFXXRaO0SIUcBdT/gF5i96oix9BwJhJSn3EvPxgyQOIlA1paP/Ro
RLuiSXzlE8lak2aPgB6ovSnJZ6c3Rxz1DYC+aif3eThbNXe+I/7qjdsKGjxzdXGcklZ2YVFT8IGK
uo0YsiEXuDk7g34wV1ljYCvZ0x9JsBUBszS9BxpagiY4G/0UEFsu+ABLmgU2kJPTNztAYbMxbG9C
yb7Zyv3/l56dOFcE3l6/45/1zF/Zsaz9KMw9AGoyhHqEqutsWJFFCQlon94/V+e9XrU3x9ik0d1V
Za9Nx/1SwuYieX3g+Bhv5eXLIAXl9G+ThwZy8fz4LQjTly3jcoNIahThCWi9iCfHb+WXGoHJIOOM
fRg6I3EVBdZwr/hana/Xd0cWcdK0YJMVyjOJ6n6XT4bS9K+IRFl6psAbkyEWYvnaIxucez4YcGXp
aQ6zJDxN40Ej+UgNgD4AqUGwdrNYNwHA4OZ2Bkkoj5G9/TZ7NSiGsiKz3ditJnsHIf10xGG06O5L
3h7p/rj6c2/M/+xYWaZYSLAiudZhQ51uY0qpaA5TdAjA2lk6qSKMu77uNPxmhUJqF7auHZ6gWLWl
5I8XxD2DciCHLK5jjvh2Tz4mNjE8muyyfCnbg0ve8xhFH78U1aI9GMGXjamBQzR6+PkU2m8T1dPC
thRagg4cPtj5+rMFmCr4+rKkAWo7o4hBjQu3M1BUQQpv4DzFSmzorRkY7t6wahCQVFvK51qRGi7g
R284vXbC0UIwSUPivSiVgkcDilINcGgodJE73TWhcmsNz4LRfpB3MPNQi7BjZK3FAUCn4XNdEahK
z5kJ4KpvDlQ0roj/SWlRDCIfOUH1YqMz7qU29q1CoWpUEIRNYmrqQ3jj/7cwVZMH98jyT6pFFIzC
LbdHXNsIMF8SkfAeCVQY2iATef3azDAoPdWzBXKkmI7kMvtIRLp2k7JKJLGZV/DHwbeRPY2D9evu
8pj/GrEcbH6v3Zt/aerRMR3z6aRmGrMwyykL3Eo5Tj4QPzXp6KPl6c19yjIxGhZw5GGs2Eu1hNi3
yeqGpAyqAjtS7f5bgknue7wh6iGjXx9k/PdK8Hfc7OK+3jUHV/gUrIK4UZ/RuC2YxXyc1ghJsmKg
ErK8f7/zQUGagFolE7fFjQrnap16sSavbKx/viqH7qHomw8oQUUs75ri+QowuUcrNGJ2gkBFm728
Pz1GQvdF0gi6HG4vXm34mekkloB/UJIDVUfka3Agbxn/D0xnzjLnreCsBtRVloV4DwxuXlckNeAy
aEjBkiXWlb9RrsPbFSR/97KVwKUrg/8cxtEQ6eg7JiLY7uhNe54PMTW5aP7PyhF9ihiAOGvtFGbk
IKIo1hCLzKeBwzoaDNG2n+GkqO50CeTjePL7OeF3L95+RtchrB7l3foL93N2wGmR6V9g1HOY7Hhp
DHVyN3i6kmEfXvNbp4ZuNC24m2Z3jysXfY3eV5XT7d+QRf2upYZHHF0/ZzXOqyO59aUQNGGUGv21
6IUED9ACeOmuu8CSsxblvWDs7VEhOAK3ZHzqueocXrIZFF43m1l/n2W1zF1rPFO8zwCoOirFLmfG
9lpdzaEIw2wC14303i7rlYrrFRlEBX/b25wc+0BU00HKf36VWXVS22jZsTKJQxFv5U7OU+Ko0K/K
9Kw8FqFXAxxncK0qUEPZ7G5+gwMtG12yBxt858KJhJGQwfTvtaZ+xosCD30cq7HJsVc2tC4auAY1
1lRoeHVNd94chqhjLXveqtfB/s3ibfsbdggTW26aO53xZtW+JgWXmCObsL+udnVzFrhKDHMS2VH2
u7CUFzpIuDf1pw6eN+0zznX3q6TwK9oIuf7xfemFJ7gE9HUHjs/ytZqGVb65MDSptaBkwf/Xr87n
IJL4f7A1so+smJwJZNp9I1lvqo5xkn244JeGUCooZTv9KqFFgnzDEvdPu6erP3Akzqr7qmqMvX8u
yPw2WhF7V/O6LTzp6f6e9Y6wc6DkiRrS8hlA8Ujxv/P3+YOgcaHhkO9AfTvIAoHUOHMLXAyx4yKr
NlzvZZ/qXaO4ViYgp51UPn0/4ulGdmFLHIG0bswIkTllaGyluguQ/Xp/q5x631U0qrsCNBsL2B8T
KhjK6NabHE0Dy3JzFD2WF5n/T/Yj0TV7wLEuYLaVry9eppxM6kTo3eUde1ANz62tvi5Q+JxPxGtY
VEwXr7M4ibX51crBQB0K/ikuRcGFqSwQ17H7g/qfReTZcIfWAOWFPSixjjinaDweMHtNM5klphJB
meNmJBVj2VTgODeQ+tamE9R7O+YASlFYSBnGeWk5aMyWC45zqVjECADRqPBO9Cdi/FALT3g6p4YZ
Bq7MkjIMq5RL6I4DSg42DMbkEknuMyBgpHRYVTl0Lpd1DF/bA5yHo+xd3hl7c5KbHUNzavT5rFBH
DA+NBEqSpDHhtQjF174VFAMlsaX9pqqoaroB1GiOF7WD4ad/Miau4MB/E/VtT/7+SMSmPDp5+Tun
opsKgx/gpqaOgnuiovPDIj6sb5Hz0VsCU7laYp5jEkRw/aTdLPOlNwh7WzNFaV/cr+Sq/4jv6anW
3SBEsKPJOFXbEMQXOJeqtrT/vsTl98EaqDwlBSvdIuwP6SiE0AycfgCqsD2fa9eUeHfSpADdqv++
2Z9X5h5FcZXzudJs1DLMwahk/D1uTCpBQVj4rGcLUDvAD7GSgu8DhcgRb9WObM5D/Y4rGSO+otrG
NKHaW8GhAfSroFI2n/rRh8SDShVxa6HuiUzVHujkjqGWT79FZwVcxxmL0ZJPwugDykLiwnMUYXVv
FlMbDydLQQD+pJk7N6eOg9JzrpMSfD7SYwe/GE8oNevtvSl9P85+XzZpKc2QLD4KnmEvRP6ksqic
bdPKRRdIQJ7mNGDGwnZowOibFIoWQfLehZMZ6xRAtgJold9NaeBg0qb4jUa7BDcnIiJeW0vJwE5l
HsacqZgyWplhvlrTe9o6jwuCiVswqUynGwPx9DGQqQapfEH5u0HLKOppUZjo1YP5EuCMZCAbfy8I
yX1gHuIfeYNf2FrcP96YFHz32XZhCiTwSvbMed4pGmcNUUd4QsdkSTg3C1MxDNFQUakttaxv4lRm
YOuUMPo+vSGetjcv8SHvACUtz+5+ZN+lMRFYliyLFMX9IZGwmZihJeNyO8jQDFpVcgggOUS+5sxS
dlSBCmp3UCF3KdKsWT1KCSTMghNlnpVb1RmBCcsLbgJXhBgoCKZ2KDwCpyv9EOjs74Mt5TzvNVyl
myqW66VdZ4Tzr9lSDSrF8EifyeoOxP/uuw00J8Smy3WzEZbEuEHLG1Y35YXMk9NPDpcQlLIu+bee
HnbKMqzvH+87Pf0H7E8Rt74HidKivqjLSbCUcB/gUJwyqXG90wdp/3qYXoQC1zZHhjQmvMIPgy0M
JKSnk6Fj6rwgTb0/bctnq/9+MhN+zUD2umQr0fGr/ORKEVlPEubmY23nz8sT/eFYRotWuCc43tF2
9T3Z4/GwwLbHYujc7cff53x+DAtLsz6awoiMkFinHuI69oWqwpcWz280PYoS2lLncvlAwn9+tLUW
4s4ogz4vWpkqdAKiu/mwNJvXSGwp4m/P/I7zt/pD808KYTlAM721/G/mi53pq9+6SREzW2/et18w
kgdnGk0lJevONK6ea8sYtDdxCXATsMdvUUZrQn+Q2qwgBrs7/bo3fDpCl3jzVILRgIqHNs5IvInq
0ROef3ZWHQ1tNnp+n3/bIHKDdU3ixTsnsM3T/sGXwiiAkVNCxn8e3aWQP4CISr3lurNrJQlYrKgj
yJx8AN9QapdKxdWh05AIr0dmPgP8Id4p9kYDIc/kT3a3x9dQCj3g8n57CUV249JP4ZMyCTns8+1t
ccdwRc6pux8kdN7LqSSLGnB5nz3J/fL7GNlS85AAoSVePpXInlNL3SVhFRW0H+RrIExPIE9MU8PW
+o4FLmyriJJ4weR6n4cTOd47OfBb1nVDc8jZU7fiFWVPuICkVQ4epRNh1nOWNkZv7MGJLuwpfDUP
prTGhl9fN2aOMPqBjQ29sam4cvcfRFKbubGaxKWWNi7jGCUMQgZoxBhVyxmPvMIQv1IE1AG0zVjp
e6dVzfyVOx9t8IOXh1lcwIwTuhkGD0TKNP4+SC46U0FD3SCwAmJPk7kMoQguew/2oHbhOJGffmwY
azNdW168oESeEAhN4n1Y18F+hrKQ1e+43UCy7Bw6MRtIY4c8zJER/WuB3UT4upbgUM2h69LlVeiH
Swa0tVQldxarBJ4ax88X1ssdhGtmSF4bex75lPt6pvcsWyZX6HR77zzKvp2sJDOMDmwbS9OhGeYr
VqJV0dsT+7QrudiqTKcwpaek3YL9mnHpM2bgBT7awIGAF66L71xr29LDcxQZm8C8j4g4t8CPJx5o
/pJFRsjTvlqibnOiVbeub034RYO2nSIRfvMI31EsBpMRwAJ/jqDPl2SWV7VczIU8eG0qsYJGoqo4
eyYdTF6RRDQy+Wp+ia9FMdt6vm3CEkVJCOdHBVQJQJ1Gp9NcBAElSRJicstk7MZf5srLO3wqYydR
1f9K9W3lW9VUcsAv9JzWoXIdEpu031dEgvb6B5qZJKcrKKzboLKcM/YLIw0VvmU8UV6SR2nghXPY
sxfQpP7JQXEjmfjAFI+13ovAeflYJ/ABkyeCTLiYPWIXbpRIRlVxQ8Q+g3PXiKqHVLRStli5965o
omooyk/sMCrKvzhHdSLj4qmDH+QRBNtQPUA+e2ZACbdNOsrOD0AVkMDHci2Ee9X5LcMQEPyEPTne
6d2Ek3CBOKhK+obpIPzN7dyUody4Qw8iSS1Dlwio1aC23z33hKRcVMVswvGE7lGmrLNp/DuRhKJS
z8MtxB+SACwb8y9rCpXZKnSS11Pt5cybR7eoEjqWO19TrMl4Y7fcLA41rPkxbFXgQOC1SOHt/Pp2
ysWyalgyRtIlZuYhtylYEMRezkWiD4GWelu7MfpGq89+MzhzaMtC1Suc5PU/hqxi70XeTCAF24z0
WSzhlzI42HTv6ZhR54yCCCa0zPals1lkrh9jLiHBakfLCmO2s/wEcUQj3NHi2k+XEn6Cp3CIJR67
PopZjiz3LEuyDwdnpJhlYBuRwX7yin7hwOeDp3jru/9WlvufpxConEhnXHtdavEICilcHzdyZMsn
FUbey2XtZkFFYr6P9urJhKtl9IaJXCAoWf2cicOGGophswXDJW425BbbCltDCGz/3eK0ZcIiPMT6
+yaR8PJNQEbgW+C1tJ79WV7nb9OBDZ9JRDZNM4RmHwXmmm4Rgkho/CM1H07pEVKu00B7r4Pgmr4F
Ocn2UUH1Wn5vQjJRLx5+O1r91z2YkbfJbguQuxy0NbfL8PT0qTnTBtu5jXB31k/esYHv624/pll2
0sPIwM9KQjbu30d31y3v8PzsZanlR7PFlBwS9e0jSa66NIvBlBjAhCrR2rBWMvLfsxf53r2WPgVe
9GUIqXcbabU9m6nlJDhmZoqQGzuo0FFKDK5NI3Mz5Mdcb52WiCy8VDy6WdSqWCziayNmnJ4Cg9cZ
HdPHqqMVoVAvlT6QuKd2K7J6NBUA+rhHVuSEjPK3IhVwRerVfDW7wVc/XvmUJZQ+iy+T84/kkBc+
wdbJHqIh0CeB3C1qb2uQ0DoSP/PysVSuOXgH/l7JNGGsR9dfoVpBecDkwn/oS/TcD4dTxID2tNxO
+OmFDoWqzi6P8UDNcLCGNt982tgN/EZuZyC8tPEiLh1xEGlzEaU7m1W/0WUXLPtcNXGUnfAcj11y
VWds4eiLQokU7e0ZKLfQlyIUunLj8mabqHsYCLCNI7qbOY2vzKdV0l+eI3VvAdRK/QNKcF8JQ3cl
9sVc4B2rl6VXQKQBD9uOcU6DVRi4VUXv0w4uwfb8pIBIxH8YOESEHi7eWbXvyceN1THZQeTh+EMf
N2gtyy24A1ElBXw/G2gVr4/KdwfucJ+Kk19/EukOSqUGtBcVh8iOkroSswJEpYPlP+vzAWL2d5d6
ok9wI5WLS4csrFuE2j7Y91oOqwqilFmYARY75uPr8//SZtNZ3vG+9ZkpnG5IwqKv657llUnbSj3/
ZROGlj6fTS6IGUZ6TxExVEoUCUnHV4GPwvKKTjXGGQ+dDUKH+/Nf2TKElKa7+K6D2fOaU6rOBR7d
8y3vCO8BxCafRINvIc9OBrHXvYIx3LlN2iudfNyDSYK1K3fXW0w9QRY1XpiUYwkYQomtkCdNL4ob
H+p17W9gYXKXwwNyzIxILpf9N06QWtutS+PlZSijpeykXEettXSGOUZBtpYYsmw5TGh4El3EoGVG
JarWIR83C12D+jiYxI1xIBgnFAA+YMJJ9wNlyqMlhLI4s4GmlU97x9u7wl/5A+dIOddYqTcavSen
D9/8JwOCL4BSaiabH9QRWsap+ye/oCDZgSD7kng4s5fQAbh9Ts9YNXoeZykn7xQsj11imOq5b8Ys
2RlvcSJZx10KF5ILvDv7KHsfzPkVpJru8TSqBpadE52a2NM/jMcsYQ28q9GDMiTs+jXcrtcE6V7B
T7rFRQEGhH4NdLnaO2b9RAJMd7fCm5DtWP4bVhpqpzGyR1sYuFaBJtBM7btky4NGbxJC3fALDVjb
ZQ8GX6aIi2qCALZ18eMkGvODwGKhz8nXwbawoXb+C43Uh2NoqR+YQcqLn+2qrBVtf2Wp3nNjdCCD
++We1gFO1MzdHMLVpmxUfWLyfR/PF7169Tdnn9yXlFmhvsspjtSWFhQFs8BQFnjUo6FtP2e7PoS6
13hr1dJgNpeTzDcfcvCJ8b1VrBdzC+vRpOPJ9YD2dZs8s257E8Bc91KXFoyFv3tiryoVt/UCG2gP
x9CzKwy95K4oqSj+NNuksiyE5trIb4uwJxkbOe7IFkvTZfqDHtYi5Y4G/nHYMsMsVp0Yt1c5EQ4t
z3tVeciCXrRoY8S7n1oDjQWkY4nr/03H3J3J03Di7s5aG8GDgnBwOQOh8+f7XWfnXsGm2myNbXBD
NyEEoChOTWybRCzAPEBpvF0js+YJ92I0eSqFJ0UN4KajFvMpk4JsMSKqLJJ6+7QeTqG+gYbl36bm
Uvzi+U4hJ5AygOTpw+i5E28WHbUVI4J/HYcnZExUfvUvngEMyH04PNDToK90RDtZ3cUcf1Vrv2Og
DnfFaibwgkCAiik2neVGBtVCxaEfmPE1AoCcmPZn3SzuziPzeL1cXmmCtwNKLKkKAQvV/suvudF1
Yl8JzD5nERVdHnItcc9nPqif9FEwg8V2BFLlSuqrNS2dbLlBdqFg2KkydJ/WMewCeONtIvZzIICC
lt+SAqe1gFvMhBaMGL1juTlj0P7szWWkHxuODnQqvi3RYXNE8UWlyqYBu7E07LG+Kho+m+qmVrmG
HMDt935OvoKVRSK2PK0QQn9TutO+HDvjEaHuShkXwKgbpiJ4boPHHXnaXCUS84bKB1WOdc4V+FGK
XTkuBYq62FBfRHD/tQwG/+pgyZrOuBfIfslCLOpzocenRXK1TgSYu7UIw6oV/XTHhTodjgTKoDHV
J+tqQJTmZkJxlnTsfOCDzRKyRS+JUs2Uw0etv9XR9G3SMxEttsrm+x97rzvx4tPa10AhankHXMzo
7TkvbyvgBMasU5SmRhQ60UAqD1FTsvoAaqGWazkr0DN3r3AqSdf54zO/Wl2o6KaVkQatKom2ICj2
VW4CncdEbIJHRraba+H0r3a/4uDbfXCd/wNuGC5cRP6LzkDj/W38AaLGUPAmLwSlwWdyEgn0Yc+U
Pcu01Tk8qmYewIPkGju7pJe8MNawDkss1hKHvAevnxlBAHcLX1b7muEnIz/+F0JukamHMdd/1uGj
gBnM29wIhKfJ9FuZBsk/KfyrBSS2QEkrmLL55IHyCuObOlnXpeFeXvOdeeJafrHbkmXMsZoXXojp
3ziWVREOOeDvoUjlsFJeNUICf7nw/SpstpeLoreRppsTRga0xadH3OrYNGRE7pcLbB1k9bLkpCSP
HyZauMbt64rC/y0EvO0OTfMjwbC7+DmUaSNLkLoyixQ7EpdP4Pjg6fsPaol+nqZEiOCbud7Az6Zs
QfsoEPjqxT0ze68x8f2k0NRzt+oCC9IsAO8VdXdUYItQrYLiEMXpOxip33xl+vlqgsh28+7YMVHm
OVF2IT3BCSM4TDAbgF0tMe6nOVtus2nJMRScAcWexwAHEC74pPk4mHYaFnnob5QTjrCFtCXSjskF
aIMNPI+/bI3eHiGoWWshOHCbkmkgFh2vvok00Dvd5Fy6xzuStLkqIcC91F1F2rVY6ct9W8xwvVln
ZjNtTmxp8I/u8aKSLa0omFaiMJ33LUpVj+Z8/sOsqWGOOF1MaEJ7Yoc6rgzKfAa1TTL0aZIZ3AIA
4oIMrnjL+GOGblVYyK6BBXgUSTqlFvU49iPLDtaG0rfcBpbhSJZU7UbyGDTObWHIzHphtBm6Hu81
Mzz9oDCPpQu58ttZVerxL72tfNAAt3EAERIwJi5+uwoqe/h2e2pfg0bZCUwcWWXD6ubcx4vZbsvm
BIcv8qryXFjOacCsdc5eYB8TUKRdvOG4jT2Ub8rnK/4YWYQ9xvst5X0m2u5AerWLIjJ/dgim43+a
o31ALxqLjtwky0pXxjHOi4qbunNFi7VoqqZq0UWCpGfCcLvi0p8FfYYJStUlFOzoUKPWCk2qTJvs
ujKDbK8X/MRN1+Tq9vsk1lTDDVxhwlFymtbR7NorZSDoAVf9Ex9SNdeBFtzV/Zwqa0XTSwMthxxN
y260CnwhpivOjsYDT9+kIbS0OaL4sXXj/HBYc1y+i/1Wf2/wTnoXftwCo42y4jNy1vXdaVSDmJiI
dfYGk0AnToMbOO85bIyFrYwDNxUK0mmqLW6ic1I8HqczIRCxc9ZsuHxlfDdH+qiWhdzqSgIXoQvW
kKbPxgh31btrvKgBmR/bLgZfDP48lmxk1OwEV1BcNNWwnhhPqmVFD53PV3k3CXL/bejAV+7ajS8D
iinpQ8J93lTCOYzQ0ojOdVVJcBXv3Xtm4opzYAmJmmjTo0RGQElK/lBN+Ft6wfrxmsD4axLi2U9F
qRctFMyxhnyyhFj8u84JCe49loI/M9WNWsLv9JMM2Zh5GEev1dCDEPtD+FzfcIadTktPG1Rr4VFN
2Vow0YsZj7UeWdfyiZvTrqGqmjp2Pis2QX9QXqYbpG5BQmXas6HH4Hs0J89dJa42tZg7BI0WArsu
HNf3X7Yuf5rg8VE/RgOvyKbNl3AqYT0nhl7VucmcM85PPTZsHz/lPCC4VqMaRIfbvoFB9R+uakXI
1BM/xX9AS49LUKW2cPxNKjrbE+vz0lzWk5uWG/Rn7Jke49Av3yYPNo7yqw8LqtGVZmZa0yG9JeM3
vKpyEHs3CMEUhPUSpQJtB88tX3cbMjR5VeITV4Oe+SDUoPUM05HWjTbgNhthGuHKZxvJqKwUyKj+
aJ5K0Nji/BScT7HCePzVUuXEzR7a1o8oGkJaaSwKDN74fFViumrV4lTH812S1thynJrdwX+46lvE
1AseTgUX8ppy1vkBaUjqKnZ3mt9yer00XNSkjUkxlWn+qcqrUEujzp+9/LdaAA03+S6SgyG+x7cd
rv2mMVmezDEgkqgnYYP8iqQDPS/bjAvPHkHu0nQm5G7BMMIsD0+C4piAFxnY7hneUpXXDTmQkcBQ
lzfMp4n9jBTlfTl5tsLjd8vg4127AiVQbqgLFBPdJpnwPkUx4NZcXFoJ5kFYPg6aJDc/x8t15Ma+
vKevPlVoEi02rJhbJmkw1o6h2IReAm1E+dh3wvE6nFmUs3Gg7wPHWqgWONlyODNorU4Ia4sLr+kL
fkLI+xfcmgy6uoGu+8/YMzHHXJ3CgsuUdXixyRZI3w9j9triiSxpiMlUpwMcWRl7CZgglPxq5cNL
TYKzG7KLQeBJCrRzQi2K8Nbu+YLIjnzKTfs+W81y7COqUgnhz13vH4jB2tZHmJrmX89gjoGmyEZP
I65Alr17G9N4lGfZFBmwk+JjHrM3M6dlfpoLDfJGFv5Edhuua83X9aOdS3l0IiphYX/O22/N9+3m
ScCkZ9Hq2XEGvb6AJwXVRascZgSrcrG/ZwEcJDcIqGfbHzfSLyDLAdZPSKHrMnohoS/kT7O4tSUJ
GUwiPbprCp2V+EpeS4WfJtd8G4IXpsL50JPQ0E/HsR8dxySQdiuaBRzL1+/Yk4/GWj1B4SN3Otqz
bLApmkkMIrtkyylz7CQeqyRVtfwLjIojGh2lhCH+135/isBjtWfYTZMQk0mjSycpTRugh/fFsryU
mK4oyRqMXzc78Ga0+opOrCsE+OCaOeA4Tc9SMvjazbs5CBQjFO2eM7bVYkUIjy/5oxEG/g9d5pdX
gt8Zc4HXvKi0tVj6ygcJnSaJXIbgO72t5/Dx89wWlDJKoA4c3ZGBcD3pbWNIpV3AsoJcQnCx4Vta
erCpSKsMjJSJNthMrAmW8R1d1C7SNbFeYJCeP1WC0Ob1ksB4FB7tbjNpMsqNzcA5ZuHWirZoICtI
F6xE5qfLQ/snZ+nHH2kQxODMdCrGozbfhte0aoVv2phQiUrvcB2UjOdt96R4q9ggMWQA0+ivyaUw
LT9RAdpuoiVX+nCgC9BVD2WsrrNAr+d9peQqsHb084rK+dGmExWFvhtZi5RtahNYRt7ZOdMdH0yU
QCVuhXJgHpyk9L7ut/7AVfJCreIg/6FQj1keNbgT8ypwznfXwpllEWFvou3rDhPOL3pk8EZjSL3q
2569hwhJKzLgjKmOvQVoYEkF2fPO+UNJeJC++IXXQoVtSDwgKeJfNi69WvroCb9W2tSiRj1dBmC7
lBoLh14a4TDF21wHwpKyK06vlFZqsJE/chXSHH/pFu6yF1eWi0J9SOsI2ptcgjT0IplBc3HqYaW2
mvzCfsvhWRmAHBgredAQZx8BdyXtgaGMWmpS48mIzriExfpxwHxbIrjjzJ+oxLfVVqG86wEgRGRL
Gmbl2gBkT01THnROpK2qZ5PhD79PHZ0BkAltyRUaYO5J8J/pyRD+L0/67l09JiiYBvmyMfqNTm/4
+lZCGkerFOv036i8XdbQ2+xmXZV0MVwcWhfgBsnzE6gjlBGgSr3508GBzglfbvAyxgN5ANdO+Ye5
XJOYTBtFHZ2eqzh+lRdUH8iwJpYRhDQF91JOIQSfZg9M6cGyhbJrmNyVZ1G4f2Ao0c/S5BWmilLL
u7muCR0oQnGWUn2d0a1AuI+iqclTkgbF/tPsfXE63bJyPSa5QN883L3HyRhy8rFYXylut9gKuB37
PJXxUPBxwZMQUt+mS1iWP4gpchfltNziqAcaZjPIOc6wZtX7yvS05OfWCY7HhQ0+WAHmgEf+nYlp
r9F+IMNOyZzGSeaLwWdMw1QDQ82710011F5oWadBPiUx58pnUIC/3xCmlxnHfumeHwK8vqzz0fBo
op/PWHxIpMS5V9YIA/rg2iqZ3rMJj+CJoiG2DOctVyS4+/k/HXnwfYslaGC3L7q62xgDRSqMtadj
CjjGE37qZ16I3CfLTZrp0PSCXzknJXAxLtgRgPv0sSlq4qO6eCkkEWvcp60S0pK8LbHl8rAF4JAM
U5SwXAvs8riesxlivM1uDriHnG6uusgOPFgm5MJRwu5uerIXdDL9A/vJ9Szlg3hKM9grr836CKPb
o7BNI6XHGYFTrJWmcYTPgxO16pHBImwjhLgqzLAf7JqpbSZifSZUisJPAPkRjsJkl/Qn6I8XON1I
inhowotATyWfFLxkFgMaORaP10hfEMLAETR7JplczTyxao2oMmoBzGhVQHY9XDRNltx5d5KZbU0e
eBqUrjLMJpoXqnKW/ICTlRZ0o1HqPS6t84FCbgV4h6FfyMfm8Tcqn4Wk82GJDcl5P+1+6WBXwgbx
NCMs0h3CqbKPVP65YUbNmR4I0gsmWhJZbDXEG+FZKaLwrE8J5bd0GXScsgdaQ4t5LVx1lOAajpq5
oMrCZ7xdThJceuDGaq3Def+chkMZ3JB0NiiGNkbRbX3iAeqYLlQMw2NgMYBZlF1ZYQh6qLgDgA0f
ABG7iNKQUoMpPLfuSTAaPftZt072wYpy4SAXxQcSMA4Xi1xQhIplswYG3TwA0KqU9SCAEN4Z582i
ss+ft+XuCoU7p2VBcqTHUIk+N6/PekDEa5RypV7PLKCHDSQsPP+uPdisMo3xdKv1eiw9d0Xjbexr
FAGesHgwmQel92vJMxzXznFzATVifYhSaXpsG4bfNZ5IVIg3fd3FCkMmqgSPhQE9kdV95fyVvP2x
hu1IWPsHU/LDu08eE0rtrDIiwwLZdWkna+M5EMAT/9LVvI/0XJX7sZnuO4n/aDU+0WCdbzebn/JT
h3VXkCBL1P+68zlfxIqe20D2ulox7zwsPUUB/ya+DK0IAJGWWwEe6OmCp5kdEapLe1ryWicRpuui
FwGOmZuLA82/cUavhSzhEqcOsLoV+mxSXtFygrO6uUKA10/yUQNjiaf1q+wdCqMgUlr/oDHexrZg
YQ7FV0ZgVMeImUFdx0PJx0beQUw1LeZIZmiWUMwCPPFqPVEuXD4QssB1770G+Qcne8mHwfGWkHf/
8NAkS4Wt6txz+bWCfpWuZd7BJFrkLN5fvp8f5/jZ629jYh7ArpkiHmm2W8RC+RPoXyjQshCDASKE
YlFVfbVEyC5Jc1JQHjzEZmsX4TFnG1P74n787p43VJyFFl0IdpFmvEWUM1DVAvcH9h/7l4/EFvHv
dzLTGUetHkWY/vLfcyMyr2+XXdx2m5koyEnkuW9TErV/kDR8hYtMF02e8Mhgia76+PiGm19liq5L
Ui348pEVw3P3O4MetCHXFQdue8DmHuxSHKIVLspFT4Kxp1gA+fYh3MxfrMlBukIU18FNabCaYoCl
1zqt/bq8D2kA9ckvJv6TxSlQqxMMYpGpBX2fw1dKv6IU/ZJHc1dA40yyvi1NeI39/Kz0fc6AMhpM
R0Pkm78pcrOEhqyD/BWbwy+mnA3pV6cjkkSfOs7BEtgDmd9hK90wc9K+YGKb+ZPjp+PkTRX1+DlU
GnGm+cGM7O76kY8EEEUfz3nPbu3SmGcB3TSj+NcwB6+ET9Ycuel3HRgAMS9l/VOm/PR/bKSBipXq
MapcD9Sbp4Fxjq5IdGmJhMcoWf3AVye5s2P9Z913JkXLkr4F2TmPTmH1r47Fq1x0uzW4bm2P+I+J
wEu+/ygalsnWLywKgzAi+M1i4rSWnHDFwkVIFdzcA2SOwq+Wvyugd9d61BH1p/wFxh5yk864054R
5wX/RRE+XwTovufUOiPZgGRRGCIp3dlFttFfDfvXgpEgAhsiSScz3rr5lAOzcBbWkjKqQu4fjMEK
6lLqUc3NwrbTpd4LCXTaYKkRKqdLpfvkNZHM6pXEMUNFYAY3f+2WYyH5Q9mif+nEl/eWH6omJmKR
L1zD6oNFK3xiOszLjYHRipY61jizralEQeeWHj973GYDfz+ts+UTn1N1VKZhgkOUH/z2izDDnheS
MohAWAAaJ/YYggnx/c1/M/CPOrD2URHO1K4nOrYwwnC4gejONuEkewCF5GD9c2T5Si8NBaMyUsy4
y6ec+APFeG2gVFwlsCR2sTfW+wlhk+KkXJlZIL2f5RlzyYQoryT6Xt8KHgvQr0XX2ZUamiH8O8fn
walqNu3rb2916yTNFIdy2PbzN8X7/fAHnmQk2FNVyqQz/52ter5Rhf0jwbZYkjenhvYkXDV566lq
rsAyZscHyCWmWo0BfgGTRWqAuWebe6MH6OUNiquaF+pkzvVizPXYR1e/UTz5PfGSddryWxDnxWz9
3xlrRvT6oilYiDotPiQ+DarvxYqFTEflr3Uwl4ZinPRRXSGYyzewV6ewqO9D34QDK3btWCYu3UQT
iLo4MTly2DXDXvZc2n4cphukEWZdkiBUeuWFx947RP2wORdHkBY8OYo0phBLmPMmPw806Q8QHPsb
C8WdbTuRlQHPFzKiNnqFZfsTf+X+mSgkBLSqr3ZAmO2//no5VvPfDEvSX4GBhpJnTzu38cmbfimG
ki6498Kq20j6GFE723k8bSvWTwFdW4640AIIpv/3SdO2yj00LNX8GByYfR2WKOB07GCT59itbydM
uPO/r0LyAFCuqpkuwev4gW6NQ2hWucNRm8ddts8wb9y19l9EWDYubOTNETlZo2qY4VjxmEaTMzPj
+1z/ZWxhI8yXDAVn67xXX9mINAmDueTXiCKnqSeSUw+5/vaBUmSRH8rJPp/qKjp9fu9H193wXEis
grvY299gsxtWkYjccxdm3i4GalGZ010co0JtVvF43gmdPfe0IQEa+MqgK0cPZ2Ff+1mg5BPk2LZm
AiUfKlrtm2iD1fJzj1bhYSNvgFcdM+E3/UUrKjujJGhxNdwiZcN4sjSx8oXi79EYBLvxr130Lf/7
g/bKyPtmOdXVdiCdGCodFBmggVJuxCey+THre2ryriOFnwBIPrzGv63EXab8fcMOUfUiTIUAinSc
F1EWK+aJDG6H7znUTvr5kUkFgEwpq1HinZQC0ulNISu5kgz1uze3nwnM2X9rmn7VPG2SFaQaL/RW
XfAOnQr+U6GQ+XJ07LI9xt1gnFpx6RaDqZSIsHWedg1Tt5hrwKMTIvbcuVC3SoF4/P8NhPAUv3Wn
ssctdcNccN4ZP6ooyGfDNX0IOmQ60I03op19jPJqzSFJH4bm+5l6HtwVhDOWi6sVLMmpxD6ibco9
Q+qCJ7Gnjep4iNsOeh2mEL1sHuc2H0xDKbyXmSfBk3hgPBuYq8dYSKxdJzvLo3JPAPIUryfWbaSk
tuyC9Rs3KEcpU09B/91v/4pGbJl2XNKdcQVX0ymaBbid8VZ7UleWXfEedibfJSvHJFxgdePdmehD
ahM08W4u2zFwIardSZcBIonYNpcLD+VEuiyplm9Svpebt3Qcjww3BO+aVcD/0yF/28udUrWrJhVK
HsCA6RQXlxITpnHytdwZufpd5NP+1zFcjGhCJDMO/gdk2FixfFQWhQ6vjnqr9JyirIobx3dh6kAd
wRVcm7BPWUft6AWW5BUbHSeWONp09rmdIMylwxSq3WQGoZJlyz4hiVdsGu8PppWVtbnbkckn/ywS
7m19ovkTv3oPVQmcnP5FoQVd+GsqEhv75IX7eXVXPNAE3IXCQlbphWfObt6NlKSucjoR+/PXHjcA
i7kN3SrQIE0GfyPK7fRkCKW4c6zY1mDg/iC9Bo3OtwjJmXiT3geBSZQpvxMDnTVtBsh9gvqwP6rN
4bDvPa4LtlFIGDuhuNfsM1R//NHRm9mEche9ClG42rkZ78Uzm/e5+2mlO+9aG5weYDGNukQBksmM
M5UkFOsc3b3QhN4Wt6/kSP1ZxvFtR6tN8ZYyoBobQIqX2U91VRrZjTxylJ54bAeno1/RhjNhevtx
KdkTonDzA45p5nKbU7N3X65uUt7VwZlomNLh/RqPOqMunm9+JSqaNSpZ10sigJPcoPvekZS4zkUp
pDz+gV6jN/Cw078ua5Rz2XTJqMj+QX56eJxQPWB7Kx6WlDlZPBrjh96OApzZxIrxgmozjrwmBiR/
74pFLSOxrzSH1wfzt3/9mdnFVHy6kfksTTp5mnpXG6G4n0W3N8x4HMRE0/DfIKpNrQj8bj8IjY99
h40k9F+M8mmvRfuOUVC6gO/2s9en45Ds2KIsLyAGJGAyzSFQyxLaejN5Hio0o+N7gVOniOaKIp96
n2YA6tbgh3MsZ0bVBJ82bdoHbyLJrhkcFaaWUnvmGNZstXvkmiF/8HCOqgJdVARAzTLoFo+eqh5N
5aykrqh+JfMv9aNmWSL37NXM7jTfkj1GtnBgNLZL/7T+MFG66X/UfIUnUsWcSfrdUjRd9J9vFSmT
gb9J6pETljgU0/Crno5gXkL5jU7ET4tHQPotIzfOEWUwgvrUstNqqbhmeXwUTh9WfLSxeBbDTXyI
t05jpREcsne489jD1q7eVE6TaBDejlt5PavPgJ/Z7RC8ZYsUfbAphykWHtItfqjOlCOL9Dg6bPEE
lnIymT26/1a15ah3TskRTNtJ8e4lu3OTRSphHXIIk7RZMGX/dcazIwDsH2XHkWKF+f9pxbVhIvWM
aRqUw1q7YHmNSdT0E/7VMCUUHl4+4PY1If7Ggcd9xFVmDhidPnNg6yWF6lO+n+zpioNTHNZeu+Ab
0nckpF/IUFg5dRbidhmK5M2NeEUSJH/iAXbV7lkZfqVvw4ur89/3K3EtoGAbXt2AI2tGPQd2HPzg
l0Pvt0cpf2st9qNrNXYSVBBJKEFeInjeVpmlJY79MN7XPWN9qiRs9NUjUyeYfUCTnIK5qgdjnfMW
dPzJHv88SbwcYuaWlO9QPrMs0xi/BQg13KM67QnXhD1iJ/l5WZbPU6sXgUI61/WbY4rpP1DsPRh7
0UOmcezL+vkdiJ+H52RqgTBuPK9a/hNm58zAjtRHG/2UH3C1HQ2MoDXjFVoVjVamSWsyXIiGRlwv
WRIWhGylrwi8Gt89Yb6y+i+SQrhh3RCXsuB9WlRcFdpNjTniG5jDH0A0ZiNRIlWHgOJuJJEAG0ho
5YnrB4Y0YQSF8dspjHcL1eYL+J/nELxhYwHpzAaGgF6xvl+LckgIPiYbLpdaHT0OIx4JWSO/xwLQ
fBrXbcQ5zcdKxVAETd9CPh5MsEQ5bhFC6HArgalrzdJM7bpu8rfcjNNSJh6T6q5GOxwJOz3UiL+v
BG93GGI3bSRuu8DHRYOKov4NMC3pap/BBeSomtvLUVfHZtacpgeseymclc5lFk6cnujulvcaaI9i
jbD1Jccoh8ySdo1Sqv8UsfEWTjyR5AY/K8gMAybZSqv6S58gPNUkZ6Fz+SbjQHDWEETR4vp/HLJk
WU10oQ/TaHkH9+1MC4gqk+TKWwfoaouy/56+PgQqcVocJ0bgQQ0gvc2pT/WbsH41zxZIdLgmpBIS
+uz63sCEm97KL5j36WriVGQ5eBwJRei8l4CgjvqNrjZjl8tJmwnZTZdnBNGYA7PxhQzN54WzDMTT
byMWogxYAf39L2+B0v6T7hgurOh2tH8h7jJUVa6/othzAF46F0Ri52g4PP1WMwEaIdIY6gZQqbGt
AdGgcnip79r94s6+PXQAjl/AcZVGTzIRBFVGAQR2b45oVE8Q+WLjyGYN171Q65zCUD0wLEtwR9c3
01zsiBapE8UkXoHhPTS3qHHtp9qA+gP2IN4kORy8XTeVA/TPnSp2litYJb9f5ztRkpAxPXRnD3G+
cXMe0IHA3oDGJ16QlNY3QTKzSTf9mIzumN7NyRjF1vzM9JdrII1FnSbYpvmwYFIA+An0aOzFFg73
xDEKmiswtWUlzsPwKlSAXKmiyli0eVrKXj+KgLYA8Msqd/tdsI0R7qH3VfK8ihOyr1AsSpSlHuFo
7kSjYqnvKEUamWMCyUOxC1pzL/6H1QbNTj5ekRp5jhtbJcl/VuMobygB7aS21SGnsYB2q2NTJO/y
ULuqQ7pYD6NoloH+K2mdrCEyZyMx/CjQScrnoA95x1Z0OsmdD5NrRDgPm219hUrA4oXh0frhjC8r
KmqyRwxXpwsFRzLtZjOr+tI06iBSX24MGq7FqmVFETNvKyQNmqudIeG9R+v7MLVdC+wzmrphnWtW
PMjmbuziJOY270mdimLfduaiLSCWdRFLgpzUD0IVjdVnmiJ3aiMNX5+eIjelWIcMZRPSWSuo498l
iMcgiu/nRembpOYAcZq7m2JXTMU9bGCRf/9Xe82szta4Pl9ZL0yE9AM6/hjT5S16TptweVvE7nmB
ddlxoPhL4A/8UkeCxGXbaRMKtqux/EJOHZq45QG0FnFgRWt+sgycUhLaYKKIRmPjbtVtjNt13dN2
EuAu/Rklrbnlb8XID5OrNGN7kOZLCKEv0i966sdO00fZ4NhgJcLWiu0bgwXEwfajnVh3R4zFLn0b
bKZZEBcwuAePKMi2NoBMokdUj6Ei1s4GGQ6pGxUpGoMuN+ygQfIaJwT6pohqIN4tT7GP65Mqv0+n
0irP53fAYF56aQ5A4lvfl24RkqvQfJXS/b2qdzQrnL/GCyTx4YJwgGqTlFYdmSLwXHxq25j//q1B
rH/fjwXUnqGkB/yr6AwCBfBnrglsoSq+DfRKVmzBJR95hQi1m/3pB7GJMnHHmpehYyngTniTqRbB
AQyn8LKCFGLXy22byddhjPTBU27XmaS17WV3m+130fx2bwGwJEPLa591KqAvVC0VYBew8phhf0CP
MUnAqmYFuCwhfOYraPCwOogawiXZ4Xiqa8IxKIYcWLQlE55ub5PRpOXPNdEYG7buN/GHZR3Fqnk2
6uni6Cv8Cbc0AOOyU41uyvDN9236J6H11VrY+BQQg404J2X+rpQkzAeNgHrOYnwECqW1t0f+/kIo
BXMtcjLj8dQZYHHQAjlTG7zDLeSxV/R5CgOYJVMH1USX5DKf7jzI4jPkZg6pBTEB8IfPxfYqmAXZ
HpN23t8Nh0PyAb9tijZEw0fAjVujkPkcTvyWVF0FShFrGxoJCfbHbHb3tMmDd03nbWdAkGt8J9Zk
nxDWmy8vUgh5Jml9C5M0kbWcZFCGyMJNKEggP7x1Ki4FdgZRysRz6Mn5bUtU+B1QhZJeLkWl/KSJ
P/lyFf4Z9TM5aGXERHS4cLcGjn9rlI4SWnq9SOH0jj9L+T6d0IlqufvWgIvP7SNcZIvTdKiJrwHl
NIDrexSxzjAKZo5M5tk9SvID3YiNpTnblhwN0gR1G43CNfJwCgsdL6i1IbqWs7VMH0kjDwLIcvVW
ABgTXHFCm+/Y/J+suiDY11iz3D2ksBXkBhDom9+QXQ8TbLl209f/wIUKlqzAOqGjS+UWCTfJovxD
83QaBlHVJ30/63GJowBQgTmUXIXb7jIaA4Pe+VS70o945mEDH0aEsFxFwuz4smQwnk7YMiUU6XCl
mJAYFshqmSi83EzWs+uS3Od3o3C3LHSAhqBc11w73bCik29/dS2QkI2+UdlNQi+kGsZ2TgujlNOS
AvsWncM+ZIfPNFcSA2u8T9VBhyOpdxDqK+AFjznkNYACY5XKvURTSrJ4X1wLXw1+SBQc9QCZ1qfj
c7TugtzX+/k2t00InlM6fJ20uQUorcvx/djP/ldmg40ubx3Ws0AqMhLETrjd/5qqGasAg8I4SvmA
APa/JSZOf59Bv+eCdgrnYIZobNbLEy8Y8kkTD+97jshkDQ8gijNl1SQKaYf5fWVFAEFMZC/Ls54m
Yhul4Fv5COgeICaxL0OQrAiYulPY8EiyVYZOVuL9ajxyAGWCzvH/Cy5W0I5/vCBsE0TQDT3UMisv
RhqHSLrNsg2/SNwyCNxQ2RHGuIlN9Sdhk4BXXjyPjIzcf87UV/C8+OQSQaGb4U8GRIbXB/1omqMF
aO2cMm89FXMPx5bV+wXWxVFDdJ9UEG9vohaYz1cJ02hnHxi38sHByuIMycqw6goOH+ImaJfGXk3u
QSdh84hOoxCCXSA3F0N8qBZYW7aERElH+SN/xLVuvWAr6PeIePtG7toulNog31fNq+ZqVWnINsnF
12khl4qPef84CHA/i2KidEqVDSDSGYOAzCb5b99bx6U45SZoM8mxCfwLSYJmGYl7gp+k62IGPISY
UYCU5asbuqoc39meZ1c+CkBMl6jox4EGhzLmaDGe5D5+a8kiLAl+lrTt7EBTOWkdG4FSVeVB1aCC
42VnTgphH7kzRKErDAg/wR/UEWFsft1MzOp3zXfTgG+hxTfAgHbYsm26GolAOk01HEVZr9yxEcsN
TtYBLGxdcC01IxPcxmwV/ovqVwDaeKNmO5iG/AsLzwuX+lRVvWtoB626T/DyorlmQe4GZ7Nuqab+
A4VYlmt+JHSxvdWajgiDTvAFQqDw0HeWvpuQ12GhnfkyKBbXlRnrGKfOR4ekImcxwedqRqCCSJBz
GlRQZiH8HIfV4qG+os/o0hE8k/v4S1VBCV4Mz21mG9nv8mLZV1hRZyaxyPHnmAcOTtTSMX1Pu7pr
UIzK7/b8UuSwqQtbPqj899EQ5Ww4HCrW3UN4Q7QuxeWXlgMCoK6gKgobMRzktB8d0OA2qOdl6zxg
ITtRp8+MyF0uKL41L2Dz9PBGI28fM9l1DZvPogFcf1R+KuFvHC5cJdXcCgyROjEpzlPImKAYcPTW
vxF3FaDXXlolXH76nD2SLVQ0qTRpigH8OY5AHY0pMRcCuKmh0dEW4vneaoOWS6QnHkGWOSRLu+JO
OFVjGh05a/YqckP+Jbc2NU00fOEXBNqUCwuk4um/lVM4vCpRbCJ9ZO2rlf0dKCJJ7oyNoqtBBIvG
QWBDYojZkAOHv9agTGKrYWJqd6bIHZMeti55QFrkWPyT+KslCJojk1/1NkcV/2nYrkVCYbRtUEao
Wd5YDkduZTNOoTFDq0wYG8RuXeaO9bShLJqVLScsKQ0SUmkAKn8cdGcyyOy65+Yf9552imv30XKr
OKlDBBJ8rbAranivVJrauW5MehI9+YV+Rk89w0+nD2AAhqKZMem6AOD5mXf7DBB4RFJcVNJCBUNh
liWLBvnytk1uFF5yWKNOqIjI7z26XmmhUExHMA6rhvVeOgV2NvH3FNTp0fUj4tNKIrW0CVaHG8bm
IzMT9Afsjq955vaRQFl71ZePQR+owzFAMdptVrEGPA67Qol6/Z3xrpsTAXmo7VzUbPAX2Nwq6yKi
vpakRolnR2/JEbrdfxyJj/Zjcy19m7PHVRV9kKzldRQQT4tC2ca3cKhJ5J/m69Nlp7Lx6KcEY/RQ
G+yWp75t5ZXtCznoSPFVDqoxFKtZSHT4ueBJiH238PMLKdX89anKBQd7v54sZtLjiDz0p/HpcULM
zyaSH4hvlpgII/BCrExcrjpQQfXAIJWPE5NySIjSZW8dyd1OTznjpqpIAeK56kCLRjrTJmqPpDSc
GI0XljfQ2WQm6cDPcqydUvEKAon/tof69XIYIBCWnAWleUJKg17MTdDOrabQ4tNo0b/gG5r9+6RY
9JlnXSSuLhzBpQpvsYabfjwEBGIsxcTKccZx4TvmMrovoYtSv/uB+sHgwXnygKiRmN0OVcEANdI8
NJsSOTiLHL7p0S5KNWInCbV6i+MjK2/NryT/pJ1zBZBvuxVIpZWOOOlyWBazBuK2hVTYdZLiaPQU
l9k9eEmC4czgvJpTiGQDoFg9GRsVQXWsaw3FMnliG95e2IJn1aNKWLCXl7prfEKMtlYf4i9QJOCv
5AbmtUYsBrCEyviv1rrlDNfhEC8wbJdbMd38spDgH9lc0kyM+Uqq3wBJzKVtbbEaE9cjb77n1sCy
SVCGVw93BFgldhaLzTWGNVYol0CMLz2tNI/YnCamwbP8BkJOcLpDoSlZDpEPPHO9/enf7E2ZCk1F
fPL3w6gclrOH2gNv+GLAJBXgIgzdxqKO6UNAfFDDlg9UplMQfCcMZNx1HRSgoAtqiE1n6/g6LEIh
grmHVMKO7DjAs9DA5JwGgk1k+M+f/VMC9plxmg+i/f/M1LuWsETTgy8zgEhxBAd6nHt0HTuUe/ls
C9K3yU2hoci7FNQet0bA9+uBKFzx2hsRfi3lsmPcdKkPhS7JgpYQt+SEeZQyShZxHqVQJGOc1jA3
1TfgYQyriZ54+3oVGyhXd4Dtkygg7unG0V608mASx8+rxYlqqjOYiyfOlqhUdoI5XQsFDGITU/VY
7P3QK/WzKNfzaZ7Z23CUuVSTsBnepTnyUJ5TAlTnkYMBinMiJWnRs34vWWn6PimYwpQVeLkGoS9H
n/N3AfF/qvJtwuvOm1B95cqAo7tpgLhFo3dVL0biD9cMLgaBTSxw/rzXn3cy5i7eJ+giyEArHTsp
rfB2poXFn+JPzOCAiOjo7+BGaQQRJ/cgKmpiuvHRvWxV8NPS5qVJk9sIiX74fpCkgXia2BoJSY66
sOXcO9LhTek7+bMD3KX81F05eWhiHf7ZILNfktmLtu5+yUJeWcfbin+1Rj7kzuNIcxof6Ohopdm0
6ZPxZngSOxnzPO6gWyUDvE+CDQlEGwfq+o4UUsRByD1srTKrxAvcKC6ZxV7FlBavimGiZL2IJ2Fg
M/79cnrIpHEB5Rnu9Gg7dt3RRL5YXYlgQY4tKfMM+jPZJ8QsHD7dGxQ4x/w6qFcTCQlFkPVzIDKc
IiZALO+4KxXaYxaskhrSaQy8wUKu1d18IDBQKjdT2Ci1/n6J8pwzAvNRl61cr+1bTPmpmcCRXsFj
7vlS6XParAcNKbznJ4ICpzGaaXyCbWzp53QsnnzjeMRbPOjrHyo7dxr3uA5avLuTc0qlGhXvEFIQ
k/pXvUx3h+7IDx+tpLX+OHqWg2QMMgKS9cxi9a9rQ50P/BcxhpOTF3iIynZG/eLi8O+f3Zlb4gg0
RAxnxprnCHo9XTUqK/gZI1XrUBnwwyMhYpoIrNxN9Eq87iIwO8LmJJkz4OcwzHusL+euMO1e+xZT
YZYYIyEeVBJ0A85AC4DbnhJdcHOLIykLCEe9HPtD2ALgEh4yEP5lFNJw26QF9VjKOxpgSheCjo0N
OgYBwy65iAw8H4allaWM/c17nj0hAwa68jzN4me2B+h61WsVVmezxAfnbx8p1EsI24KOPCG+IuWZ
IM2Ac0XrtRCkUO3qDGWIlBNWcwsF01xRmKE4BMQJFmb61ICP4vjZfCvWRkhP/snLXi8pVnUsfBGJ
zaaoVS8pobSnpMqxomk9LANa84TpCZOEJa2BIxG/l5T7ubENla/AIIt8Ty1gLxEQXxUBeoEQ29km
pMIpYfPeUQtc3SUuQ83dPxmeR2giZZJTxI8NLuoL3w98XW0xG/rfaV9u5iFmY2bhBMJqVdnBzE/C
z/BoJjQncaJDh9w+FVXYIfw9bh07M62Fq8gF12txtuOuIC4AsnvckUQ1sbWbn1Sw7qiFcTZ+yOIH
UcuC4ZfUzRYEk6dMJjDFRqvGzorrW/yO2qHsX1kvAXOpqo3BZ77TULOS2g1XDy2llnYlNb62S58s
JAizBYukLVn5caGiI0YZM1LsLkOcnnVCZX0gZSrO5o5bzmOysoZDW1FolwSzc80XXUo0F720VRs5
ocoXbRkFbyIFkgV5TRlE7WEWFAS+7eT5SvnZYRg7wgGW+AedmjWjbwTJvtOKdqe9o/Z3jCxBPd9G
CCR7C0nmRHxf8F2vgAYSP82P9zZrTC2ImCPXw2DY9hkNZ0m0NliKFSO8PK3DwHOmSz1GJyBIGxbe
ERThR52/SmS38dgnNxkjZ6vak7P1d0NzWkJXbM/BRXfi4eOdICr35QFcDtgxBncrqfnX9XvdBySc
t5v+EYqvBcbx5iT5/ZS9Vu1VGBR3cOsC+RpowY0niatrJWhsgEye+JregR/9iDmuQdOHkjUqz27E
M3xfJbApknUjdWwHBoIkKa0K3VQPmluIhi8WgOejrjdBS76pRiUCscAm7KFw8eM/p3c1o52Zx8a5
sa9Xpq0tbVjq9p+Xvtv9jDDxIjAFkjDZ7Oz6lADc752tLaRfe/C8VMQS17kJynFLUYGYfiiTaEE3
1DNeQZJpSFEWxCA8iflzuK7652re7RLSOF/E5GyGSaFxMyCGHA5orymQOxa/4TA/IefQeIdMdu21
49j47yGcvHCMLnsV8aTXSyXoBMHCynCohXFQ/hwTR5fyq8eUQ63fZU3ppI7KOMJlBUKzIlP+Eaty
aOskZZe+J7ByU2ACNMZ+E6OOpdKf//YY1BYVUrpM+8hSWtEDih+C7252bEScGDtVmgSjtJ4yQtUC
DSRd85W/35iM/SeSIzEd2m5IoZW8Ir4zhOvy+TnMJtMNv5RCypuO/rQbOzkwieTqpUl1sStwJ82H
sIRYD3dVDfKtrMOFvJoxvfEfbBIvu7CPomQZR3VpP88Ia06nT7MKX9dPh+qTw81/A33ClReha5LT
yhZhjxrcWEz5rPkqHoCaWmMDWeU93xL7xmkoXXYDxB4EIujA95sH0k3Aq3VHfZezSZKxrI+jX31A
x82VXK6Vxma1lnte81wPgOP0NgnqmzU4hcpMjPOMcGDaz83jWL/LqkwLCr3I+ssJ62oQ1bcWq4F3
omthLAl7IVKTEKYfgVUdA19A5Tmo4A4ZkRQDRMsA+J1gyzqG1uThueJRDVHfgbQ4pDBa0YxjLP7p
HjxU3kUOIH4SkBC3ArmPNyJr5tgb9yWuaFX3r7JEP8ViJAudIOPHRP1t29mCtkgknMDzBGkbDrab
n7Ll1YFB4bAlzbUsgXoQe9JdpYgtoZyH7uniMqi+U7hd6ePlRqDLyvLQ+Tkc1STv9zIPEBY+uvjf
MAt5YNgAIsktBev3ANZe/0qQabhxlqUoZiqsfufIoAns8PnW7FBuEiVqlY+TXQhjL1E5AHb1bQwc
pix0w9+mpF72ACgrbXTYHy9T7GA2Ny1lkwUc4J78zfb92CW5o8tXaRp7Io5FwVVE84KdLIUymUMB
CyYvB+dcMpu/DBCNL0/vU7ocmqpX9m28dNmA5KV7FwzBxhP+kTBc8+MvubdNLeERoiewMSwT6ui5
yhr0l94SKxSCw2QqW6eSIO4y9SLRh+yiDgTzMRaMEmm3aHMiTmhQ4o+DUZTHQP0vfNlQXyScyytQ
DqyNvRVGpGlePVABJMrHgWHUKCTuTHGyo12adN8ZT2Cv1p1hp4sTx/RxXoevUtyyjqUwM8deee2O
sKcsTPZHbHUVltXpJl9ndRU5L0roSB9CZ897TJX4YWly2kQ1o8eBwNaKgLYllX+6OH5THfrqKdif
JJ3hB7SudnJ8ZHNW4BXBXwZ8Sf1vsRg0yous4vkoxAKTCObk/I6kn/Zk8e7j+Y6+/RH1qzniYsKu
Bsbv+B/E3R6gA8zGVbp0E/DWMD15sYQgzuVAFXVXiFBC16Csi80n36LJSmydZzofP4Q28M3/dMvI
97mShOOUcYlG2QTjEq5ERwfEFlESB3nBdPYYftFjtuR0w1MJfVGaPSWLWmQ4G4AOAOR/YdKaQnLF
8IHy2PVLdHNp2y//v1masZZ8FDKr/vgxYb0pLhyDuJBJTtSxes9pMWw7QlHRe+50IZVFhzTnIfuZ
MG8gNbhqJnVp1Y/O9XtVBjU4fUiz3tPeI+vCVkLdUEkslMOvmG0rsbQwaL9gqd24Yyz6Un1qD4iK
gEWSUASxhgf0cczqTETJWrpKwZOkpsS80Wf1rguxNZcE8OvnBcmz8JaF46DlbLhe7YAnEvfgfJ58
6AWpz4jg1lhlJjpcsfTXXr7bNjZIzByjX8Iyqn2qgk0SDnUp3rIxhn9kimHFmFaWgIASd1K15IeH
2V7QIm1ZxUrcnQZwax/6x20y7iu+p6HgdNccvKdR1wtO4uJgdr09mKBn2GPJkqsyx/yR9ZmgvHKL
jlJ6ReJ2BzX8CJ9dpe630McW7jJH58uXXw/9Bfm2ENYmnjzExqQ/RvAUeXEOmBiao4C7Yz8WLD0z
S+8a0Pv++7HBVFbcZChrIDPQYxksltTgsOHHKO/b0to6dzX7u5VLvr55y3AZAigdWT/6qknSE2S1
wcgWq/8Iu30df0f7WA1HSakvB/P5lvLsUnus8L4eNWDQ4QO1ORpCdSFaWGuYYkeapDh+eaqHqPml
VO+4zLplxtjV0jAQ4vQZqRVg2t5BOvJu+A1t7E3jlLSQoOdtoaG0B4R9H77gjZx1CLGcXTu3BB4h
j5zrgS9iOOvw2sL782s4hcniPfdnzF3gBVkK6dFi4Y/cyiR+jsyTFZ3+L54tIIQsaWokaZqV+SM1
l82/MXYyKsxXRnRpbVN+MmatmayJlR1F1yCpNQNiWEVEKx1kiKKH/CHAAeWxeoYv8rt2FCBEDhqT
NVeXOSbRM1XeyCcJtrDLzdL2dBJqunabPgVyPhBqqsriucreAC2CIrh31omOcVxBh81cYcjCqvLB
jF61k1AviBb0B1+S62eeSNYcBvY4HN93OKpleLTxlxZjHgtr9dw0HOKlfuc4Jc0Imbr4UEgmMuhu
6iXcoUanMHSDGiCN8dM7ZH0WWa8HcdUGlXP+Lp050qIbkrcSe1BVNkGeVJwRZb63aTB/GRF0kYBq
MtvHdjteTGaoyOThleA6ZCeT9Ay0Vioj9wr+y3F9WMbWYGwY8muzi9mWE5kb2oist12KNXyTHffq
mqBZfiUUgp952QTvI1U1hhWryAMnshPtxbNtxxB7IODa8ntj23OGSI9EzvHcWBhX96S2qbgtqQj8
L4BcQ6fvHRazcGpQjEY81Jf9GHPZU6MbGR2um9vykjBycR0kynuG69278vfFRmtgnWw2fmWZdv4Q
N5RhA6JPqQwrRYqjJefELIirB+uowgHp9eCs+P+rFUEnibyiQHsNcHXd/qHpHGEVFz9zu/r/xtqk
JwMbb9QWXkIHKQa6+iRF4G1TiePhaaeGXOp/5rdFiF0b2AFLW7AX2PLL5ueeIAo8is1qAwwKGw1r
jhzWKJtQUEhq7cx8b27jBlyIlaNEOamD5cZqHQNV6cfd7QlSGgYEeyNgCDmHDxpKORsU5y3rFOhn
73Mi4PVv+lccMZXX/FKIYvLARkD7SNa2DOWAqS1gRMlemPSMZ5aGJ8/RAt/jstXIUj8RhGW1S5I2
8HzIZsxosR5SmcFyr5Ygz7PUdjYmMZUAUNPDOPYx7pQVSW3pvNCDzA3yIYgmDq8BHGLT6GAk0u0v
ahS/oFFhry4ALDqzp3az5+zn8qTDZVHlmP18dIrO1wVYZDETDqRl5qaNhaIXOR5qOQkBNQ/nJkrn
4hIv1Rdz0esqEZw5iY0nFiOQez3NQpK+LfO/IYGRnIdeNSvfx1UJgJizVrXIzbJSuBJZm07eNOA6
NlgdJq4GZGgDccx/CoAwMQLeVkCA8nnngHZ4AnywU1qQ0B0PH/TYC6KWx7WOM0OCCv2hZsyu00T7
aUw/6wQ7K1mrlTWrXLHO5stPvnhSJqMgHI/D6dTb0g7IRR5MIsb9BWNA44iiqlCDfFnJXJTMYj5j
Dsk6rXdvevBvMJWRxHLUnidVCZgQz4/EfKXi43RIzPuzLSMSyHZ35y4rP6O2+Jpsx6/BA6JmdPnh
iOIoXUjK5+tI2mNK7SKT43x2Lsz57HWWqbcWRzLjOSJJKRn5+RPehbnfFo4ml5pOcr8PxFdMGpJB
ebC6nIx5TnU8du0ibX5n8GyI36xFBDQQeHwq08WdWJ0rOt+luKnPP4bqfnoccRb00ZgrHuMNfzSO
Cj//IpcfXe5kA3UR7FPrCPU+z1u2Xm6B+ga1VpxSTmRbBYHRKRn749zXtZPBK+0QdXvBFeL+dlCw
MtwRX+8aL7kftpjBaM4pemczcLSLKVSuPOMMSDUUYEFD8ZeT5HbDNYgj8zVPuXnfsYT3G1v042qu
OsPgtNTEQ7CFtt0Qw5rY8icSdiWjdK0hLNBFTNRpIeUXS1MHAVuMGm8DpFyBDQqpQa2tcXdM2tyU
3GwAslZTFalwUG13X0zieSYDgqfOnQ6fCxRHjFipuc89EL4aiSLB8Y8qs7F4ZOYc1+d3EFne/xGR
tF+Os+AVVy5pS03dya/I4PlDvQNaLHYN/g3jPKj7y3yM6IW1sKw/lA/eM/W5QJesp2Pg2uwSp7+Q
BwbJwBDthtDs+PenCCZzvWtK6wb5J8+JCESd5JzWCRd7IYZvK6EeysdSGyhK9tTz4dDcgc5aiulV
AI8rl0/DzlCwfCPu3t7LJhaIMT+5pAgicWrihMqJSpB1+E6pmCNkmFSQzHXO8nvIuy1OWaL6D2gU
ElLDu3gIffgF1HXqsyElojfLZxh3qDmEavzbCNAKxPH+HNhGi57J1BER9ltPA8avDQAYsQHEdSSb
HF+5pZhCRbfO6Rk+RzFibED+eMn5cHpI0bqQTR688o/CDGmfcuYu9cvcmwAy5elWk3BolyYUb7RZ
KcbAZ3eNENdowrz7KBG7JWH8QLElEIeM3Y60foY/hp1q9OFIJMwxrfk/8C6sUNHixI7waJ9j5pty
tyTd+IhcM6p/+NF9AIK9WcWKka1DhW9HikYjLG9xoypV7KpxXUVm+GqE9uGujZL3X3UV73snD78v
riJOf5oxPqqSdKkcVCNYDOKuJZkzrBdDF5GEB4tHjGRu5Ppv4oAppxGlMh/zI3IRQCZvYGjMm2R4
ND4FGh4rgoPYLpBZgoIhnv3m23VMRGMdcS6aFGq4458W8jtMdY5EdWeutGmfbxNNph3cf5+jNHrp
DJwBOxQadV+k/cADUdroWD7/wnCyUvrtpgnMf4f2FHBFnFGou2hSVNQ0v3LW53+kQ1NbHBvkt6+U
OYRIiDmmVp8XiRwYBg2+f3cOug30026985qSM/PqGgy0CDOgQaqDZUp2fnaacXUYzmgYbV9XC31D
2Z55kWVqwozuBXwiGBK4TeTzqfsvPOSpZv+/MNkT0lF94m5Gy1Ac4434mSnbaY9lBqVgbvZCUgEr
imG+wyNGeUvMD61115/BO4hw1G2mVThrveTvmsnXQ1XksMt9UMFhNWcuXXjCCWM4zZh++CXoKMTg
GGrY00pGi1Q448xNe0wAESYv41/n1FdFU0iPVoNoo/8YktOYcNGx0SCHomH92vxzOtEty8UsCygC
ifkxX7P/9s1oXGFai/nVSBFBO31uTqeekqTq56AyA25g7zFTrY3BStGlPj4f70b+Utb9WRMOapY/
a9wOG7m94DHH7gTlXwVzTsvrBTxxvUeoxB85NS56kuS/xuthT4bkdmIJ2XU4iFPMyXqM9WqgUPYg
36GuQBMXGGt2K1AMIO+wRle6pfnw9cGj/xO5oTxlqvBNrsHVNIgo1lpUCsUINWyOtctoviJ0ELsN
OmIxpEnYU5nZKx8a5K/dOjQoiDCY/btOYU3f3/AhRxkmyWIiAy5Pu6iWmO14pc9JPtbSxAAYL84q
Pf8DZsMc7lcMZz0NKZSjeRHqL6YDxcjsyC4kIGYHf5V+qCDtRemMA306CNabWyU949DJ1aaVNPHJ
RzTFpqIdlMcmoMydWm/aaili/D/Dd9EbA7vR/exxR0Xh950qlyWQ/FRnK3edIN1bIU+ocEPCF1cg
oIo4JLmsckrPEFsNv2V2+U34cUHvWr2W3TwlwtzQifaNfePfw02Q6N1/KsyCzTw1Cbr3BW+r8Wic
1CRy1J/K9kSzlh+Ao9NsCAtQ2z7hUT7ic3vDcWZkUjJxRCkelOANUvxNdeMynkBbcmO0BwRRGjzC
XIzLFNVwCDJD3XJINseR03/EiNb0iU/e+WuKPBYNtKkyeVCwICtW4o89zyUFQZAQZknZoDWWu1zB
C9F49g3NVZsEegrXuF1AXMUOds7kqRaUY+I2lCHuQ8opN5MrdkOyvVKKAaLxBCs+h76eet2pccas
V89pIxzv+aAN2/uZr4GTp9vueOuCfcX9XoBgYJsHuwy12H0xM809wXPiOyDbPZRb6sUVtreDOkLU
cVBTnSxsS9LOIEgTk2DXKsLCF8TeucLsaXmHra7DHrisdUMK5YnbUIcjVgPrspqMpT0hAAE9m5Hz
PGTzY7IJEGALajJ+8POPdCP2gc/X+dhUY/LbXhe4warSqTgLYOkCDt2xhejqUIxLsN/WRSesfdb+
kQG3ErgOjnxqF2kLm2oxQTJPn5S2SgvJN61dGS6SrJ0Yvy8N8XXimZ66lzEykDVxDCPiey9YrTEM
f05GAVEhzlC1zf5XFtIyFtSnka8eGZ9hdd3RNJEAzTVTfUv8eDveFn2G+qgBJAR0zH5AyFsKfnYu
qnVL84NPKJ3v4t8DOvkDSjcXDMbINIDeuinCMKGav9tEZN4/cMmGvjfxLOpwpDfft8PJB6rPyznG
yt5aQ0WLAMPHlfHKd01rbhrdfDVQTSW6s/Y7ICnlVIud1PtF/JymS0Xfu2mrn9F9bhb8rbPDhEq/
1JvlJRcrP7dLZC4SJ1B0yheZnVhPW2UZicjmlOLGKxHM3OMjaG+g6TT8yitU35Qd+CgwDVFyISo/
eqj3HKUPynZggVPTfxtupMQEmOCj2HTxnditogiVa1WAQb9pBw6kkcgt7494D1ws7R6vTc9W/V4a
UdpZZaLOTkDHUCKsLgZeTDhtapGUD0rIeBg5LfLYl7Q6cx+5oEBePORXOpltYdB5Oqjj3WPNHBBU
DqA8EJ4KwMepiChmvZqVRIBmaSmbUmAW3QyzTKdQUnQ072ITD+kGk2W9RhGijCOlFgraI3BUcgaS
8EeS5LNvxS+VNBxdmqnKrU705S3N8CP92nxzQqnfQwaf9M9xFAs9G4EVtHuFeVvMiwWc9pdj5QUG
dEmQe8cTwwhcX8mXdE184F3jNb34ns/PUjSlbJskM47U9zpXUut21oIgFm0lF4IZxiRqiuHiZYry
01/OLDtnIo8ydlyOnC2NqzbeLd5yKCb3ujrWqOKK+sH+HReBNAlnaurpMugsj4lPVJa3TxD0OL8b
31Zupklcfx26rFGPM0kECJBxrWKETCG5ePeDel1LRlhDZEQVZ9/WGzQlkq0bRfzCkqKuQBLElZJ/
FYkvaBlFg04evSmeUbe+dUOvWmqBpe+455fX40NXbaHGRV2FgMuhaYhZ4scjA0tp3wShJ3GXBlcb
7aSdglVt3APMU1SLak4ysQXbzZYURourG+YlSIsgQqRz7VWdHYBrSuQmDMi93LBmlO/3/5elshUc
IxxOF9FSBpcztQnyVxq70zsgCtyv/tSNcYa5QT8x3Z55pX9cswS/ThHhQ64DQto09em6DrAA0l+A
wYgVmQLDjIKYah/xPZd7VdefataCY1NaBZXksdDXkADYeyP75cO1mchCukHgN+m35RtjO3hGPca6
B+vqYdKHNKfw/exEsDigEWQCyRw66jEEgNrgtkVITCbypptHhATWWfKzPiZsqEJLj/s9mKU9z0Pd
vpBxZaEpo4SAgfZ7iGBRRUMzHE+prpsQ2zn+q1FtGh3sm8xIcsAtnEGQNPF+j0kuLHSmoVsVcjfZ
WYjldpQHXptJNiDBCYkC9zKSqUJCF1ojPE+b/Rxc87aiZq8ZSAxHGcVHT6SgWvwYdmPbUTmpcbym
tjdEqimNWu5jxekfql5ZZ6gB0r4wqbw7JYzduXxBpqz0xDTWgpP5yIq522Yohfxc5X+oKnvGnyPv
xgdcsZAjO4MHZnccZQqa1Hrzabd8xZpSNLsN78A19b9xWqhO2dL8kHmURMql9ietgtwNP0P8MjNA
jfkaxaoe7riN9yCB4swgjPNxhzPPr1zbv4upmIbuPKQhmf2F/2b21mctyBulQbBnGoKyLONKgcx8
qYBMhTcpnigb2j202oUdqu0iMhg9DZMvitIsyV4VOONYfEnnsqErb/nU7a3fLWBcNR71I4DcBwJv
SWyYgNXF0QUCvqgqxgLrXUTjkPjoxxFZf8aKgZlEG8Ux7J8zOadQwJrLaS5OpYu/1Mk0cGvR/Ed9
WFWV5pdwGxmkyZXCG7Tx+Oa87Ctok0PVatfRIM0YwSy1Q/v2xOVE+N65lDsag0x3mWXCluhsqUqQ
9RSOVn58xc/fZLBh9Uk+9KIsSTPF67V/A2exq3KRVTMDdZGfMKDz2BdLWCXlBFVUDzJ6/i1mD6s0
yGiEE7U5bA6VlXDgo4Tb0fbD0rDq/W38ReFQczsnLlRSAChwmhnHvAJmAI/VEWZ+KjKyDvgECKzj
UngUSWEtTpGWvvy7opU4IMrPrtMGG9WNMvCHjYNS+sB6lapF7fkS2cKRziZgUqMwQYLMhFtBAPqZ
Wr+jRblG6m/7EXcN4RBIvwfdx2sU9PFk9v5cQEiasdMNCThyRmwe4QARu1gjubfM5PQqGHlB7JqM
pIZ37e634E2LaQ5518BQL6WkVSTQ5NTrG5MCvqtrAaLcpEvQyqtS8Dem+wIXGZhTAjfz4oHPuzEq
tjeMz04nwSjQwLCnm+X+qBc6/jqDMdzzIkfxFTzv2Xa4Xi63q7r2ylQMgdIZXROjbcrLfxNfPKgq
edjW4oGYl4/5gG9DH5HaZHKU2hIcpZAIorRYlGkwtRghiyosCqIZSpG13DIpyBx8Kl4/KRrNyQ4J
AO4YadDqpibfppvZYO+5cy770nRcIyofXKwk3Ih/VV5WG8UXDqcs8MKBnBHAvJFxkxfc0l0Tatdd
8JRMczwiJd9xDJpSE3XX/7TwlAu+9PprLuuT0loCSdHMNrobI0nplJym7mitH11H2KppJ5Wm37T4
0c8zLmOYCUWDf9kgp4hAP41qbHVTNwY+sQvotxz8xDix52RodhYfnLNwLb0Z2ooJbW9lFa2UOc7O
ZSBdKwlLKUeycDbHXRn997iyRT3+ipb5PkXlW0c8p0SwAPVPzefXrllTkPB6XZWfg7UadMyPP7RC
aPuPzCrMd9e/QVSa+VaBSnN1wB2cZWsT9bzb1CewG4EQcZnUe3WUG9ZYt0WvFF+/WoXND2YtJQ7f
4WaCGv/h33TSpMTUXSh1VHWmRUfCC9Pi+ph7bnTWO/fz4MCl70vlh5qzUQeqwh+JA2e1B3MLpiu4
rof53J/bsaJFD5JzM/WBbxeIcUTJQEzBcpObXcs6s2QmByqlrBQXg7hzYsNdJtntpv1dZzTEfm3G
qDog+4yQ7ytFmuBEC+0MLMHIklWUHOS84m0nbgMcaCQs9Dwd3YuDn4T2HPqLjo4HXarLQbqGFJUF
AQjuayo91iml3EtOvDpiWcTSHSq/RaQLOzlOE4X5ggTREt7cKiSh6RO2LfzK1Mg8XIpXUPpn7w/a
ZJmWXXaD8JiqYkjvaxwLZ+TNyjYyFYG29EUtxz28tlKQXEySf44A1qr1M99o1luwMoMbzC/+mDE2
ftBQ+eYqV0kozzyA4RMGPx+7LdmeVJfT7KA8glOxlEKl91JSUZIerDzipP6I/YtpESpBm3v+cJ88
9ojJUH8XOGRNsNa0GlSrDBo34jSZ9r5caoRF69ZWV1wC6OmOMXyL/qCS3D7gF00FheOb2i/8YIEZ
F8fmDSQVOK/NhJ1UrQN53qrWl+QNKRqMUi5oYAbQ+06brlpsACc//YoJW+srQ3KLkn3kImAQwTTY
U6b1G3Kk2kIkfvu9QNFsyU7qG+nwPHGDZ0+S+VDA8QcnhYT/Vu5k7ybiD5ByyIn2nH+mOkqmG6rS
wjEoAseIvzcqGxApwuwM9IcF4zhaqbtqHEMe2PODGI+i0gDQeV7CBP4PZofOod3EfP4IxuVl92D1
AYyjNuZ3iOvOqR/5grPeS1OWekdl3A7mI5p/EWmhK32EZeyuThsA9a6QH9gj4tJJW7RHtwwcI4N3
jzhiVoUKhj1mJAs+brctr7svLwx+VBF14s2rRILCGNPBZCprQWkjmjmPKQyUcUoktMR3sjT7SnzE
YyX7XAESdoop4SwgU3hn2DuhHOzeALQQcwowrEBPMo4n5or9n/MAi0pt5bg+9WcIxUaSEyyIgCmV
b90Ig/yuk269o9qQedwzEERG7bTUBmUp7bSK4Ldg3N/tiv/ieatT1umkyMIWKtym5ESnJrFhwKt8
SzlXlLClDYqtXzehBZT4p7vghDbYQ3Y5wu+fDQodyJCUsQcaZtDYD9FoWoaUwAAr2lrqe5zm+zmw
7F88+x4BbEhG0R7FRWQbehl8JGso5ktYHQV+WDMkQdVD4ZqgaMlTmJLKGiNc/43CqNPkA+3+1MlJ
NPRX1kBWh1Bq0shpT2xNdl5o0NlVIVqo9mg2hLaRy6Jv7ByWLkLCfdEcUQpkhtRuuIGegyZlFMJi
EJSVVeCZxPua55VdlQi5R5ZP6VecSXio1epe/MXpHmJlYdBN1am4q0/ZZwAA9FSbKtPuYcAP69Yd
o3Ur5KvwMgLH56zWQKTmTF3KmF7EYJb2tOOMJ6NCN5NZqtR6NikWUjannizyrRWziI57/ZSQ5QS5
KVtUuj0HkcICrH2uJryX7HZ1hckgi5rJgqJiBq3GFszAHO6FpaF0ey9jMEgj4C3Lu1DR9racIX3V
asmOjrVWGmMbyx7cResdseupz5B+Uo4egQbWwYGZggm4JErcYMrXBYfbvg2zOK7pGaTmB4cnJirH
LBjM2fHNAMfdH/02rSaThBkPgx353OnN+7kGsfeSbaq8YY3Px/cj3WMGUGnLB887gmLmq3pruEaP
PW03JxTaPz1pl4PnU6shHqFiJ8kyjYong8RKVJsEov6NPJK8rHJbxDjSnLfQRt2N7KBzTrfnzYwP
JGPe/qhD84trQGFOEWX+kab4uaj1p0zQOlkviNEhAapMZjk8bmDNoOig8fabLXY4z7F5WA1rUd/O
pVGSeCtNQXWC6ue6ztEoKyv/zoCHHeCFCqckfz3I0evQf7mdqbs6qcDWUG0Hafe78DTHvo9J+jk8
+ev/HYxT5t4iaCHPfYc0eV2zUpxOqK3BY7dadqFYPLyTATgQwAGrLw4+lAD5cd76swCwCjx6XZOG
aZ5xvPhwMEzb6wgdYLJR9jRmgS9otba3HKcwZ31elzmzhEF8SqOIIqHa5on6i8MgiAvMc8luyNgq
R2uuGZFhJzHcNIszOnk/46luAP5JJNgbtmYrceq3IX+crlQmuf9i70tUi8PvtvozTcsEUcG09HTJ
QS0z5WWZE23LN7kyeM3PvSRRajKGtOs7a1eJvPuIwMIk9FDkuJ70+e8gFxvKgtwS7nFnW5OcHSSd
K/78Und8lqpGIfSThgmVumexvq8ixJJfjAh/uHR5swxNYNxmbvajfHjkGAhkFL7ULKO6kDGmZn7l
T1ufVkN1aifMk5sVr9gkvQS3O3QLA1BQQqV1vTUQf8XeW281Ei4no5tHFHb5F8Nojabr37SKPz98
93Kom7Dj1OpNDgz/NaBA/xpYLTlOIjGgIjvL3GaPkr1sDU98iDxhPael43pjP3ZmlvGCNpmmH87s
ZcqdoC9csSNGbDVwFzvZ+zydMBddN/pmBtNYanvOSPo8FyuaKzdU5E7eizJMYmVgZMN1whtvVP5q
pMrcj6L1nMTNWsBjaqNpMdR8FW3eyAc9vn6c20W3uglyzTCGHOuesmQKIpx8HfP7ZAt+IWOsPoPr
A/T0OdDC7Qbgdk5c9qwWYM/eyX2jWkCGi/O1rbEgLGLkWVzK8KCaopDaLzlg+JMHxXhDKV21RuBt
Xb8VPfU+Vfv5T9HWI2iYSzVPHTbHNJtT1jwzIsNu8FlafMOrjyRknN1qP9ps7+NiRU1MJjt40+iG
5MzDVKmsL3dB3KzUDCiJulwEZ06yVn+CwdeTMmy7nv66Sp22yJmqZbs5+DjBZzdHu0zjEbccuFeM
49+hP1NRyNdB7meLMjuLq1+T1+6/KApYtZmGt0BpE4R4YJGrYUWNYaV2BqZbCyfIX+tsPoJSropx
Rjx5m6hjQqRDUd4D2XJcr9DM3uEMT5ImtafQMgk+NakNoGlBdXIdIbnWTM0vxNU6GiLqQFiVXdiw
B8lVb8qVGY+Uvx4UGIR3ZUJ6V1Qi1DwAJiGCmBnqSsAMKnMHq6jrYlk2/HJhSdKV68JxrMz5qsQK
ceDsrJLMs1OTnP0y84QzcOONW2YWGgPjlzkWBjFXFe8D7nKaWBj1Q/15kyy8vNZGix+UlnY5pqd5
kuge66RWPGXzoBOXo0+qgqFPwbOx7cDHfBpNTtbBVsODBYC015VDMUvnjIOkIpOv8z0MAwOO9x+O
XDKbRoSXomn39oZWp5JSl2dB9McWd1xzPIpzXhBCUDuVktLDe2ke6nvXxmMvzsVvNS8fnHmfU31D
M7dgxBFuZ2xEDnC4eNY4c8JsnAZ9xvjmpgE5z/VEkDCW8syvorFBr5iYzNSB2dDkAVltZWaP4dem
6VuU+MCg4G3sYx5GurgScCjwRPnfLVqxLB+VnLT6ImQmTScFgs7H03Gje+hblGTbk2drdwJDxxed
5YMBw2Ur8BHzrxASuRRhUUFkZjTG4OmQ7jjdblzn0AWrtt9Kb+Sw7wQq/RlHBh8oxlXluFCb1pA/
zuWWOzu3IgE7SJ31p6Wl8WciobJSHswJOxQeiZrrP4d5pM/isXsH83eDf3UlM4JkHJeY5koORuNB
nZSLGzm7/GUXrC3LZoXZXsMBoq6CeZU87JtwHsbvzLcYGAxXZodHK6CHOsKtJT27ZRbO6Dfh1QXR
XxJA/4x2XBn0/h5yD9uIs/2MYz1GGOfp0BR8y+nJjIqyDhbeRYEzgi/j12E8Y2deAzDTja8gXaOz
SuUkzDNPoXG67c58/YkrZ+mjMW99k4g+QEWIMZRIbRxGO8ftzKLwZRWIvJUdgH3E5goyP844sJOJ
xs7rcjKKVL/dzSXnrsq324gQWrzOhioX2viAyiQHFBG0JObdCb0fZHyAgyfkZtj5FDol4reONMDn
iKgWjsPV9jMCQ1BUxd9Z6dAy1mk5aHJ2VuRxq/80mXwFcG602wkyoklb8170R4E58Vq5dcG3Gc1/
TJsq7RH3Ku9t0gNuOXbyaa/z4CJRTr8LuqQrSZ9qYlbO85C7YbZEYXox+h4FngZIdZpLBdBsOAo4
7EmDz4ZxPH3ZqSBRhAVc9Xi97TS2m/yUnvaDnb5QAE8FcAWMCxtHrWtVWqfmGMTacktYJdyFqmut
+z2oEgZyZ6RRv0mdFDrfTvkRV+7HoBoAMpikJJpL9Eg+lczefxMi+oVhzBnpmjmpP99yOhpjMIT7
QNpDfJfGWgo74hMJ6EwM/pXn25U6Yr4jU+t9uNQk8n5DkkTWuv4iIlNLZp75CiMJRXOySakWzwTO
sCZgDWquZ1fHd2kF4MGEQsdP6hcutlVf1jAB442QWJfV/shcgiDfS95PjZGaZo/8+9DletMMbFjK
HaYZODR/RmJw0R3Mevc85gEpNHPN5OZb7MbUdDA2wYYwwadfY/pe2PcVkJThPiQZnH7WdljU5s/k
Kt/tJmIzrET0EHHISYoo0m0g+UGVclFeFzSrOFGwdW4qD5XSDLOUAt5sWMrfurTnblZtHdGb0glu
g7qNnIodhXeiTe/8YommYHzHkuZLS7Z3nq54MxzUdyvsoKYi4miwQCgcAhofuUbPRya3MmbH8nId
Iyab9KJ8MhwSNrm15YYiz/l+AY7p2K377Pad+p/thxXNSo+PZv1t2ZDlB3QifrHL1SnL7HKD8Olt
QhyslTxlrPyhNqDjIP9DHPoCWjU6kAkrPRRScFMU3a+Fa/F/KtYJ5CbW6w0Gz4kBnixkbBJc40PW
fk7uMjiFukvcJkeSa+o1XraQkyt23Zmd6Pj5f7tgKSZ4fDmSBHmBS7cs/bWyQIlqUNBofdrvzMtQ
ZHUscnQtNDG+NxSv3/qU/LcZKy0X35tVfA3e7IsnVDNnQ2G/aqhKm32FHZLj+rkhWVeHv85WBUQV
rivwtBdf9KTZC3ke7zm5UMBQ7ZNU8SU6vSCv3ezP40yeQUD+k/3u4Euyc57DTMPCSVR4eRCSv+qp
XBpVND4AHwNL4BPeEwdfD1sUk5a1YTixl1vp5FzJMkxYYtZUbn0TxUOouWYwCyOEptXnF3vmoVHz
sak2mMblOP5qcmYM1+ac8udkWs7lQZLrcPswcqPAVDFO3i9ZLHzm8MSb43RSvyZDmcIWEr6Yt751
HnoujyFtYzO/OjU4Q7XxQGACJ2Bvav+/sIY66oJ+7f0YAQVLnSVnYnd7j4OWrnYIrnCNY9i8wfrw
OkGfkyf6h7L2tZ413WUbdC9WqzEmRjdzHT370Tu0o+pUqVP8lwGx/s+MoG+ya0je1OU8bTZkYK4v
cvQwRr8wtK2Fgs0x7wRus+KHNfRMs5auwIPh/o4KswFgfRO2fg/7dvEemdXCKhcpA6xgBAvwZ16P
atNEQbHGdcrQYQem526Zq0M4IDD87KD0cR95Ihj+pveytqSOWy4jdc4771kd9mfutVGvIJmob84n
2G07+UaLguBfk6CwGJDBInI14fa/KT2ATo5W8nU/aukpRDJa98tYBaXwPSIl9cAAV4AiMYcFR/un
TfXIwPPtC59FGOF5lFGIZzzrqACRa2qd7bvHthEdhD1yeseQ5oFhYWhIWqmZkfWmRIPLEMyhi+X3
jDZUZ0JZTGUyUAQ2uL1Yx8odOnclGHwxSsmqXv3taE6vVWOaG7W6YNl9+buCxdHWT0ITdOnCsOZs
mutOY800mehUdBOLONcg/chbDGDO77iHygvCjOSTUU2ljjKbn6yugDXi0kUwlRcHtywLBlvb/Qv8
np94GEivJbHaXxFaYF7L6k9S9tx/KQyqlZoU3Y2kIBtvP8hwPFvMqMIs+eiV6ZaVFYGTzrQgeY/Y
UQaA6Wj4hAh4nxJ5oLaYBX9S6XB+ISkAhUMx49DMYRWTUPIi0TAOiogGoBA4DxOKYD6dxv2mS81N
6pRLIsqHMFyMxiOQrK0O2XMgPIwhHijAtx+ku885T3bdleKMwLfEqX17JSEAMMwQUKa5uT6XrNpp
jsBfeLHfKCzwtsDH4W4N8scVX1exqdZEDU99zPHnma7C3QS6+ovQTGq0w3f524qgmDXvAK0Lt9L3
xku+ZLqUCfFBv4xJ6N3vUFMOSwKQjmdUanolmzJT6ZKO++etBIZ/IFpFy1v4P2kFbdAFtWaOXoft
UH+xpaXyL3fEHjb2GOzTBf0EBMIZ7l2LS/jeeP2giBhzeIG+RViXqO8ZuEpnh8FppiEfGiULaPM7
wdyN1ZNovURvDJq4+8bKScfcJRkccHV8dcIhH9SbukHTXkI4Fr7YWWsTIcMPVTDJ4bXmblDPDYpL
ElYWB8kNXd2jFI4JXkbqI4ohwWjIogxhgWQsgTjQaXsFNJ22U4UT3s3ixvuiuT/fcKfoU40DvTxw
65GIq0eTMzvWY8WgNia5V3oy+fw8ch9oSNz7nqyJ/M5+GQbggYrirIV6Ktn28/DV7UkhVxPCGzps
8Y09yufmgU6Aa70N5xF8i8Hos3RKwbS2Kmr/RRqry56eHgAzn7p1ihFwaOVVayiGFEUXhKT+pzfe
HgBPIpUzm8l0cuyJZAf4kt002Boqvozw2BBGA0wxYT7HGLsNscrWwOs88037THYZ3qQBN0EQkRkv
hipQ36ra4UkS4KTn5we6Tn/ODO943vk2eeUnCi7RPCqimRS6DHfG19Oe1pO0sO9Vd5ti1VhFvFwT
uyCgsjeQaTczkk8scS8JPs9WPoeNS5TzDkcQ5PmOTslCgsWFJib/n3XNEKreRYTWO5tAGImS5NpS
iQvmYMx+8YUP9Kr5LuxHv5p8AEvlOxsN2f0Fadh368qjZHN4fJJx+JRJoACu8x1wAZWs7djzTgwx
6YFf4erbh7Xglwi7WqBrUAAbnA+3BI4hyLuTBvQx3Jt6je6QiFQm4rusxrSEC78LM9FqyEo++8CP
dsFba3q4ba5Swco9zxcdUyVQQ6SbF5JT1+PKzaFj0KR/gjSCrHoV9SxZrEiHX4ifsOFvSLV5/1h+
Qs/OjAavVcNwmJQbjD/sdIOK7nRNzhh/1OXkp1AAjpYB5wr4nAcDFsn7k6/NbzZ8S8J1yfIiW/72
XdfnbdnfPIppcP3f0DRKUNM1+9I1WiqrrDB4fwLwBBypL0j9gc1IMBk4377nhlt3u8dZPSo4NIjA
Vq93t3P4zmGhYbNMPGZweUqAze7/6UtuMi1tohvtiUHWvzduybP8BRCyeqEh2F1LvtuwZJoaOaq0
aw3UsdfwPsfXo/X0tw0vEnbwhDmZ+St5Eg3AlQC/ODgoxgZECRWELgpnkRuR/TMHuGoajaCl6oQq
JEFYLJnbD4NJPICK9gicQi7LbdrrVZIfC0JkWFTtpn8isDYdza6qvb/g67nGMoyxH8geiJdxAZl1
fJYXyPs1xuaADaj/2s8C7trLilhbf3iWYyqPSO9caCl0yt/szpHRRSw30jbWCuhJzvnQiMAKoW4L
LBr7RBjLoXqEwCfB5N6qyAVZs6YXdCvd8a90Qzxvf5CawHixUp88Nb8ullZihYkzO1R0Lh6oGOVz
xrWJN1hSjtHyTJP6l2rzRkhr6GU4yJhZA9XzMhz1xzQjqitOXWGoWHLeWBNtAfh4ghr/ssg5ggX8
xlt4o7ixJDfLFfpplkKdIeiE17csNU0Qd19+RLRIS25Yv8uWNkdvm9e2LF9LcC+vZznFZCQfeDVz
/+aUIVlHqmTNIWJsqf9nqHYGrfpqFSl9zJFZ3vySLLWGNE7IzlR8mdkj76a/mPsa5Vl1ckpXWc/c
kKa/yotuIadNgdUamguvMEh34YUe+T7Mk+vO3K2/9FYSJi0NfKT52KKsdrHSBrO0twWtpGTlmSXm
v2HOtPvOfhELUezUE0BtqULeB183+ULiaXisjgreLF7YFNyjDjbr2LLItanE2A498tUAjAHaLBG3
Yd99atmr2HjKVheGSyasAh2l19NcjV11AP8nDZlLZdX1QsNGsISWBvD0xfm7/iSqdM3OsESxYNBb
PS3soaYFWgu3L9+O7smfN2MW02uPLm9n7wakyJpQGLw3Ea5CQ1Kf3moPTRW1ax7IwS4Ncxddp/tz
LdguDHy5kknA6xduq1fcdNstir3sY9sIgbHOSMyQKy6vgDi2wCxu5TSwTriP8vopv8bxf0IwmRlZ
rZbUyjfVGbmcuWatiJ3QL2qeh1/eYAv3PaD9o9rFHv5XMjtTyNas5Cy2+n+SpbiMlrMLe3ellW27
ZldWTkW+LeCZFg52LLJoHOa205qrOUWOdJX+J96FwfXTP8rMGEVDwLFPJS2tPtKKuT+dSj9yvwqZ
RbuaBnmuxur4wSjFLLTkDk7yBO5swil+YELG/JKzqJnZ1Q0VP6abdt04GmbVMVyWMsZ1hkrKb1rU
NMrh1BXLiZ47AKxCl/fY75g3XoHsO/SzNjWUDaoQntek+F4qW7Etvz+sqrLShnCBB4DPxgxgC9rU
Ag8uk0SufTX9vPWGIimd6DUXzjFR6wcO+mQG82HtQy1+V4SLeC8iXPe0RFN2C2CpUg/TXrrXeo2I
tz1E7nRRR6K6UMu53KY6IEtMY9PV2TYuOaCHR3F83m4ApbAgJWucBm8aU+/ErWSB07YYlpPQqZFW
xY8kb9Zc9YbohYVzezJhDYuQFvuZRc8m2cI9PWWS87uSqiNEZzdNfevYCCgHwJ/4XWhJomBUaFPs
4n3oM9OBHTNuvf9XuV8UxX4260B3fzq6MWGjQosuau6pg4jzqttmkzLCwY/QzqSto/W6amRoY2/M
SEBYgBn+8ozziX1Hn/p+U0QnlkTv9vlzu/+8AXk4vdg2hcKDcJp3HHuhSPKVVHZJFL2A0H8qs0Ys
py2J966oWAshm7MDosjW2Z+InqhzGhkrSdXvyQKFZukVZz2o0fa2KAEP5VHlhYBud3R0Va4hX6Im
MCdycVHHPAmJC/QLqq4BAyDDQM8V0ljrsHwpYJJJ/gJGmCXAQpaAZOiyldTXH+PJt62P3vg98cTY
vvtA9jV/FnEc58/pgMX4TTGqQBRg3WZvlz95pGM2rP2YZT5iq/1QXPYglXIGlPcz6M7dab0vM0Dj
ngvXwrHirvTRJ6L38IVYPNm6CUUvWeSAF8BHsm4Z43PepE2ND8Zc2iUTlSrAt3zDGdBckfVppXJQ
j7pvyvMLCs9WpyRoOSQgctwd61RykT9utUIhuw/KA5knPfDRhdJmMwwPn8VuCrc8sg9ktpISQlCh
0FdsYm6rzuRQXgn9FTh1WIxIfqpexZnTOtvQdfTtggAZgGm4LMWNA+e2B6yappGWrNd7upLzkWkR
X+HrLj13skhjifzjhJKbIZBiji/e8olC4rnw21HkUVPahMjssdIyAPwx53T5HQNHXC1mWXN3JIWj
NpWBk1P4r5IBCRYOhzI82nG23SeuXzbKZ8MRZO9571WDsh75oBKXMnuf0MDudNwGoSC4/0N/aKV9
VPggFWuGwu5DSwLhH2M7fUOYduy/D4lAQ4pcOUmLEzLaL+stiSBEXUOGSq2siyELQWjCQSa0ehoO
r86NNCs7HAEHau3OzNf/Gq09BrFtnJGOhKV77yXx6KOdFxBSCJnfON4k0vSfDr457r8xajVuuRF7
dCmo5fzOpAHlJfbGXDHHUAaPA0ndvySw9DFWdJe7SOPVmpOhqZ21l5ox2q1fZw2UwV3uOfuL98lm
qMnQmv6g6kpP+QaULiJT9OpChLyG8YZL0VH6W5ApUCHDEcIpItUTU+XHBh+FGuyISb8ljCgt9Mgi
7LubtumJw8bb6WSfqXGQnPd6hx+hWKgqA4L+Ly5JyJ9mNVqgL0f2yrNL/tW3vSZ2tzRgZDz/5hlI
vjXw6wn3tiiSFfNL22RDQq4VWkSisTX9tzp0jJvUwEM8tfmSi4Ydspv6z70cNA9v/mR47GXzXhJh
+LEJSURtPtW6FMOKFwSpnAwBKqNm3MS35KqHFCRiMc9Q5sQPUCQOIqJ3eV5JoS9dbybRlHRKQdKA
fQUoJtVS9xRwGlv1JwaI2JC7o0ymJtaFyrLBQDd3OoZv1rs6qjGy/cegB3SYa8S2RuwkqM3KMw+d
pEaDolF0XUk1U2eXBHzIEXRyGxKU7tCgjhM+rfWYMxlYdubdBvli0wgT/QgmN+ohF2mrNuu7/yVq
b3NWZ4Ia26Ca1p4Y8LdjTop3UxlU6tSpZvqqJnXJa+TBC9LCZSkkr042wh1hv/62OX78aJ5hVpPA
GsvjOs211T+WcKBfyzWZgGkr56SK2Ip4ir5A+4fp9+Y4Dy3wJb4Yi4MDNeOpJyLEr7CbJJGhxF//
KaByzV3N7fRiqpG7lGqnFlt50cK7gZNP9a7dfZ5Paq4ged2saCwsgmMPwc8vtIlu+ysMC7+JSNoW
WIEcWqgSgXplygCrRqOa4Vqm/au8tC/c1WLaeFYh7dVMb67OKtnqHlad2TuFV5fHNEfephRkb918
KaqxWhTZ/2WqwSLw+v7SGee8QArLfCQZRTnpljFmZbrJiV88VttJVZurYNoDo/jX5fTiNzqamwP0
MzEQKjgc3rqQnKgaex9DdbIHWzTaQgDK/+3GqCsEKNejZQ/vYXcjCt3MCtloOjxxlw8MBoxL0gKZ
iNADNlnw282GfoH+pyQMIw6K9EtBTardMiJGgimGtpSHL5jzSazoTBKIt10DV7PQfOPR8+RC7P+Z
LR9T3dPdKrK/B7vOJOdjOeuknjIaXhV82korrnpLlR1Im1AYVXcLlDhiAFNmSzT+pDqFpWQqwQNy
igASkNqSsfe5payJfkGLN3ZAcZ75Xdwj3/hSI0zGYF664gBQnRbXHiaHyAbEKEDj4fmuDzdFNvqD
UHkawt2s8UhwrHfpqvmxDpJ1BVMQv89I9PspxF/YLkfu9ffS2L9q6kzLUwrQmrtpgV29sKYX5Lw6
Fo4G6r+ETJYLuScmUrbw24VeCZyR+CPKEl6fuwIkZU+AEyXUl/XjXikcyLBx8eQ5lSU64lfpH7cq
FDN4GnMtKMXnbd8RcHvG/fIsre8e8Oil8SC9fpcHUuADorbDDBiFtTQ4ncUbpyxQ/Seb9tvZA37y
s1mHyn57XRTvXckbAkxmDhRNO9UQMccXCIiIZ1R7QIZrICQaXRMJanb2X2e2kaqjYX6VKte2owkb
wkUA0Wi57thgRPACQozIYKaBWJbNDwSn9I/vSBMdTjV1mhYO1DoAiL65cKM7P2O0Qt0q8r/yHfg0
zj1yWJmTR2pbA491zzx1oQcIYZaTARa2/xWfDQ3JrBchb9vahJOL+Z4fiRa8caJTE6t+ZV8C5eNV
vIFXOzAETwdZpcROstFa/80f0D10ciXDTd7EoCDI0YKZnZdB8kgiAmZB5+GspkgXO2bDm+dAKo6Y
aRCNTwl+W2RcAwAQsnjNfhMiz9zGIgZohzmn3ZRft/h6Vf2exX394XK/JbUIpOtJsppt0JXVe7t+
yXFTwmlJy/Sv7oFxl+Q1X0jaOSdLPJxaUUdrtLQGp5grinowfLVPTbDjYPVlzyL6JK9TdQyDF19F
8kPSJQof3OeMSxNWragp0uE/PYBaLTzq75GS6GK1yi2Zf92sa5YtG6KSR6yOwO81IBHQ2xJd9Vnj
w8tuo8JHaNKvvPWbngAqwQIDx/8B233nICEZttvV1EO5LnYRRkaSDhsKAjZbIMm7tCoDJlWZ9ZAW
TuAKF5AGoIdQewbHi3BAay5cTLnsC9+iAXmhbow4lm/Jl5X1+jJFAm3MFWPNxs3DQ4Kb5RpfIha1
MH+IwkYmV6sZR0OshKX0ts5T+vs2AKs0/dCz2Nc05O3ZQaNjzrz6nD66XLbgWEcoL+BS2QpxE+T0
h2hh0Ip6//neiQqflVq99Zd5c7TWP1kUCmMmXnzkrBrkiwvnjWrm+bKOPvnxOO+KOaIcnHDglz9g
hVW0tNe+dlgYRei50wjRvWCIv5F/fF1WGscvCvz63P7+fzi4zrwbqFdXah0zBPRTR7k7sMQRU+Gx
uXG1PTVdl8yZhPdhfHIzXWFIAMAb5VzGPTwryFeVPGMh0/lWg0VDXatwoPog0uSr49XgJyTsyq59
pO2J4DoWKTJ7Q3/5/o7N3wg03Npr0W5FylgTmvqPnt9gfSrdV5UrBfmL0POaE4Au8hEwCNDvHY3q
UPfZYIBRmU/bKrREfyd5j0w4tHYsLt6TkP0WPiEUYIEviNbqgP0ifPhXWqz2JHNjPCV0SfoncabE
2LTzWsVogfjfPM2gT4TsTv2m1AArHzTA/iWZPllzPNbV46P29hQPV5VaULuSnjjilGo1aVD4QExS
YBb/YkHW5ghuvRk+kgI01DMkseYBoLShuPv9kUbs2b31WUvp+tjeaJrv5jNo3UJFrnX9G+1XvBe2
mqv3ppzrQ19856KeG2oa8W3F717ooPQSsExvh9gCDcHOAWP0hjfygPR5nWp4xfUMSAP84L0A5nbE
n2d/ZrMjkI8dCsvO4wuAfHyoFxvjpwZBFl6pvIl9qs7foWebhLSWDTQBSML8AkOD8F9pcpdOe57+
Cjx1WV1zXzd8NK70WZP1K+It+M/voYoBb8vvbV/GrDHiXkJgTGNfH6LdoL7RloEoNWwzMEdWL45T
X/Xl7wTezs+OZqd1uoDJZjrolNylhjLrK9xA1DZSm9YCvExzNC/rk6USY+UuHmm/BUp6PV+uiy2j
mpwoAMUiRu2BB7jp6x87DXFjYYbOwiHuJXN1Oa1HfNwUmioJzZsV77V5tZ0qFzJr/2ORwX1COUUS
qqCl4Yf+SqAfLXPlwo30XktcZEwhxPNaX2ERlTHPkVKQ8zzWe8nV8xEwqrOoEV6pM+5hAjjQskFv
9PiiJ2faIE7BQfdCjUWnwheACG9MaMXGfs7KkdqhPbnmcW2XYeQSF0OJbtdpAsKae+oMuT145Sus
uBLfEdCz6wvLr3WdHzgSwXDxtTfM3bthLnWju3rVRD4jZGMRvg7AJhCA/Ssgx1RXwmTZsFnELsa6
UIPOF/cSyBYPLBXTGbmePLtguMAbAoguezygcFPbKUYMcpMdyLUgu6jXMAeezDFrKzR9mXQ3oB3A
LmKF9cCBd+2tfZVuRXmANKE1esO5cmxiZA+fvRwO3lYGb1TEg/zsM3KySiviGiydaQZKyn2mKr7G
nI4BY+RwS8yK/PT8maSHEGLyKHimqzN3HSRJcLxJtVdubJNGEo/gpiG5TyHLRhbGJv7STVbX73pP
iHZns5M7l/+VsCNdhJQkhrJ1TaejwEJvLgstghppWgOGHQFGvnnDi/FQSYrsweSekSvG4FKfQ8mI
OjdEZ/S8VG+nqa+qdVx9kAZFG6vnRnD5AjB6rxo5kH19IexNsjitJJ782+d0Lgplx4IKFpeyOTyA
IiN0p4iaZGDHC4aVa5t3/oJHMaKVKBVnUWo7bPH0JITnVXH/l0Htpdyz0WivXm7fNiAfr4xDjrfa
sx5IZVlXka2H50/VGXo+IYiNGxw3bllan0bbhpi4G4FBbpw/O6ItB8aL2+G/73TQ78B4w5/5dQFP
W5Sx7CeAS3jlIIAY+WkLD6Z6H0Sh1eiK/Iv7BV6m3OnrHW+FmmCyWBdInF7a+ePoqSTsYVzOSIC1
Tal7Sb5PHHzVIzbBU9xwzHZjT04oysm2ctfQ32PySb2X+JiWl6JukmipkoudvXZwZGEu5cZI8Db8
/1524mdXrd1C5bm5MbZ6nTJiKCmDGpf05DK1gpEf/buO6ePnlrq/Fb2Fiw4sOYnAATI7UHODw2MV
JOqVVWBix+f1goBeibM/5U8lTu7up8t8VQji7/hAI1od4P0l5eym32P7oFXXeBI/e0YTRi3iEVQm
cClxVfhfgFXgBjNST0lDLmPYEgiRQSXibQAKdqZcLpPxRTS51dTwQ0eNzIIA67hyIg4y2XTVlopm
QKmxnQ+gwPI6ZA/2yEJuWeMOAmJRfHZmaTfMXUa2YLNnJYYlXYZ4+NVqXrVXqZBRsR1Jjj4mKVny
x9XpVEv0nF7mY4mih8lzDNYa9SK8XUUzV0xEDMqs3sGaxq6dmdMcBfCkCtPmcXaAvpIxABHZf6XO
JyyCxDPLagH9r6qTc5uvzhQFcFgeCDGvRjEpCJqKs3/FdXjoUXqXfKySFbWaYrGpFWBIfIsGAXxv
TB+m7IynFk0/bewcvzXSi9bWY4C8MOHaBDUmhXyF2kQerpjjeU8gZ/8C56b2c8UM8wuElj4YJATN
HAtHwTOk7EEGyR/x+6OUEow88y9R8lW5r4Nl5IyDAPOEpqsPWFaDncJ71WoXFpIb9MdV4vxNImnY
Ku5BrxSGgLcvw8AJtNBzCwjO8I0CrM6atVklzo9aL73KEgllPwwdFW56r/xPOvS0VaYWhQfGJntr
k8ZeA/pIsBdk3bWqEZUDFk0BNsfAI34XYg/ugcj8Mmw9SjaF6HRd1xiOMWv8QJpRm3zbkUIMpsMU
v8cRvW3hJbgKVJ0etJDRgIdqxgDMHhCPnqKDeFAdBgIMkvi5fc6BX7r1BwHMlg3dVY7WJ1TJE8Sg
xz0EVE/NXTt0NdWwF3JTaegtU/mJUBNbbSHFbWtavZWotgdLi/a0n3AlO5p8dBJBTVezbNQL9rkq
scbeih9ej/8c4VHhWq5NXIJg5cigcW/SlS15PDI1YJPd5evbVt3qGCktpb9tWRL9fh4zVacIJ7PI
sWbjdSR4Unb4uLJ9mCRq3Yi/dtg60Wg9rWZn8SmP+Tv9XCOJl6uERd3rPEXwn+2+mK0XGRRbE1wZ
s7WBNGqTPJAbZ9ggV5ud0Mt0qDobTebh5JgDDuOu+BmLdYVg8IwvHOBmgMY3AUUQftwbB1UMNJ0J
S2QRIYE84xMJSdsOuOMcQlJ3d55B3W+7Tq3R07wzxCqoVa4Rmp9wtHcKxa0rC0rpufLt9cJV9Uga
inW4iSFgUV6KKf1U38H5j+h+N/luLrQk7zlMp06pq2dHIt4+LBx8Y6i+NmNZ+nigbuUajk0a610S
keRcq2sPYAICi186G5hlxD6jS+ARVtRgHqOyk6zCiPQyZHp7tZRyAX++yVzh2+ePyoJs2pShnRod
W8uIWTIhVjTMUlwKi91r7rOa2tnRIoa8HOfVF+zoanyOnw+LOdP9yE+G5oNc86eoZ1RaFrA1pb1H
Xs6g9RtdiFr9/zNDIVZSBERBxXdRyXMUWv6nFX4qV/C+uxPKq3A4zB+UY0Zda7FkvGDIGtATm8hR
0YtHNKlQIlDo/ieLgVbjiAo85RAD18Qk5uLEHGF6kHH98ipRayR9icmf/tVUM3kYiMjAPjLekTRm
uWZu5XTKxmY9YUE0Oz9tftsStcWqRUiWLH9ZDKGPLPCzlLrklDlwKX2NPXy76rDWBLIGpSe5cRsR
85DWhiix9VczkhBkVbffUdT+QF/4MKJ34FBPgCBAbLSpSkZigHISa3u7srb/Hy26o1Hfrp8ZbS1i
pccVU82DMVIldmvtiip8J8NviWJH6aZYdJxgwqWNK1o4J1LVfLJywPywlrrIjBCQZ7b2cmned/hz
sa73bJdRbltXtKA69Cqm/7xINBH7FoCcmNzlNR/dwnyBnMr/2IjrP/O1VXf/UKFimXIUMEnujHBM
dJ/Pgv63QgLbZpfEJcqAIW3Pp/KOj/AZ3WCqFeGiLCBjfs4XMZ9a2aRVWUH3aW8qZpMb5YiF4qyB
sRflP1ZR/73C02tajhQwrROF9r4iylECaPwsrkJ7mWlKShKR7ny+JVuoJEbIwQQx8all6CjEtRwO
0kK4mwSwx7zE/vUoZLCHOv1CT4m+3+gdJgX9YWKYkIyA5ITEqldk+f6M8alyQpHJZH6NLKAKMhtP
tkc6rZCA3PWbxLYktYoNvGigVf7EsSknnhjF9Ih/MzVFZ6qxoLffHouBRpPYWYBORb/fQZ3BMoIY
kiKZMOS8s3e+D93bEPhtxv3JZ7Ie+fB92N4vDqQNHy1po136+Yaekrs1beeL2jy8kUVnBxBBM+jQ
05bnl7IwieJklQiL2JvxB6qfRUgWzJ8nEhvy0IMWslNNmTx1GdfG1fEywkic6vYZ9gaikorsQDIQ
85JnjepYvAZ4XxPgpPaTxZhYNc557kCQ/114zT4K0tSpAeZOPnjJXCEDS0TRyLfNTAmNtDBZFkt1
WQpzeqcq2hMBHWq1byr01raIvkioy7OQaFBTr61flhH2SM0YS6Ng1IiDMrqWRXMtkavuV9P5KEZj
ebLTLwJiFZp37chrRHGlEg8l63NDrPDX6Z5iTkVxYlubD1cfTrKfd+yy08bFu6lmw91Hb474FUlk
0p8Zvn0+0ScOQ3HSwUIEs+oSmjX9S5gn+yCoNMTLNlcyt3GIHda/3b6GhFPTPHvngirRSK0ayTtw
MGTOc419IhFR9Vn93wUFO9MxRNfYwE20o+PkZXv0rrKw35PQhS7C7wkKRIh0pf1fGK7TrMpKJkad
vldDuHjgcvTn3HZu0/C5vKUJ53/XJadQhU0pKoavUfESfZb8ZMMbgkltfAkwqIx7zTrHG4tvY3FC
EuG6pbdb7pL7C6Gh3XOHAd/+1sBH114XjpoIlZ952LQniKC0Rg2eNQvf6smsbrIClrwQ/qPJVzOI
qxUYUD1+Uv4kAFEFZgApmbCaUh9XJkpCfLWYwADdwkYwk3FmYPRC/elE2Nhblt5ay0TjcHsuW98M
Tic2c0CdyyCL03v/E2sE91f+xzmWH8GMj9btBlIhaDU1yfVRgzc6Q0NfIuRtPp/rOpNbuZCGEhnp
x7ZBfKdp7y8lZXNmS+9GbI2BYsro0bsNaQuZneww0F80T8IYU2kw7/3gBRZS7T1aVNjXes7sLFyt
sSCUNs9LIElZBYVO1JI5auIhZiwJQB/yJjztCDHI440t8xNqqPVnwSa1zWhKrs7Dp1VxN9EmOT42
Iz1tUv7IIbdIHvyeEqQ0vi9bqsAp+mTOuduzZCm2xfX79KNkj3uHQdyft72PULdvIuDyeh4xMkrh
+4WKmBm0y8Ml/a5/l/l/vfb6qcDK9CBacT1+Wc9gfnuuKeOufdQjd45ETgps6Qp+NKgjevd9FN1q
AagmMomc9P+SA6oWJApB/N9owijogUSLWRWAtnvhRTWsLnk8+BPkLkDCkgR7sfotnnfdv4Vg7+qL
XOwblhBlA1eWmjYeXBbQkxPnz3wuHfhvY6Y338V9ynjUC2KuamZDS1P6v/JMkwtPd2aF2rG6bmGU
lz8dvGxZ9ghIbmdUIOSPwsgGjartP7H4Jpn3ZpuHqSv3Khp74lfMOmpBPuQtk5HuW75ijHnkQj+G
5K8L/yPJZblOetXrfABGImInJK5KBPd9cMR958nTTPEx9xjapD4zfN1+aKItp4pLfRtYXRv2ZpaW
1c7HdEMm9TGfCFT6LjGWGVsiVSl0Fv3UAhnPuwTBJX6A1TwFAxBEDY6r8pAPOgTSgEN6XE59yXJW
Y1iPx8uTBs/4csySH5l1oeloh9+uSgMCsvhR4lYQnBv7V23KgHLoeEegpkiPBF9QVc8xj7g1JZn5
aeFp6E6CJ87NeMDS8yxd8vEALwZ3Bb1sU/BqLAqUkMoIuJFfzYIwRVea0F3gA+GzMAes0XA58AZD
c91Q/ZOi4cVVb1gtgXq3TANVVRqHG4qmn4Pw2kBJ7QON6ZIIS8YmACjXwCr6GUBy9ZkS/JoTpc2k
ZA3BvtzaiPDlDRlSpq3sVN+77RHp5j5Oot9pVGY/2glBz0UUCFlQR1mOtl1fTPE32EXqHvk8U6+V
XirN+sPhSuuMs8u7CTSHeIPeynyek71JgdrohNFHiOTEx/c1mOLccUJ3f2VypHFXQ8q2jh9K9uSx
w00DSUUQFBsWcRf1U5VHLmDrq8lBb2vvoef3GxvPpbEjUYhA3mamZEmupwqT3G4uFpobFJVRKES8
bhYoCy0RC4yovkj+5MKNr33odqAKYXQY1DgMlIbxwfwCLTae8n9Sqxhs8kUANww2cUpcTPhZH8QF
sW5tJpxA7bZbHoSS5zzMSr9dYrM5dDu7dq275UAjpW4w2eFp33DwJsK/+c8ZM8zRxwxevbmbjyby
XZ7Ge858JnKNUbWNtRbcgd1LIwI+gvqmjIZfFbdBYD0BZsjH2IFhVU6DJtr/Efxl26RD78HsQHJ5
+M3MErbJCeK/Dw9sBvUF+3xEaWyBTvtVhsxPj6AvS6XB6i6TgyIz/S+MR1Qw2onlJtMpHFJK1e/1
+vYHru5OW4ooIOig7dJhvjjrqv1NsdZhjgtSGZLcCgCbKb1LShO3KT6fwkNaLulaFDNjtFl3HYJa
1UffzaWoh5WCxQKGFRoFmIsjkC9bzHvDJxxfo27tna03vwnw9ksD1dfxvdZNgqdXeScENNp4b1KW
iLL0Z3YTH6yUU1w5dtCQtKJ3HLlt2X42LREsfHPoeauFvZIMI8aeeTi4FYwGdCKM0AXOq2ge0p4O
Wjd/FR+dqkvbHc98ls3aouz1BRTF+OZyYGJyalrw9LbIvj0unNvc+AejJPpZLY43d07e1XIiGinz
iKtDRh9yaGhbWYyjc89CuzlOD6lNLhld1IJ8C8yNqBb+6WQqAqPDnYs5id+ZMBt2nFJb68jkpHvK
W852cZKQG+/IT1uUGZ2NlWkPtFIr+eJZiix67Uru0YDWT2m/bthSGHJfxEQIeS7gXdEoCEY451Q9
HHTGX4W7o2Muh79UMHnAWtQuJcF6AOQ7ZfJOx3r7hmyQWCncUmxQ//jwjbGu65VOJr8ejizGNA7x
tyQoYHeEFGVX9bIMyLcYZEs+UeQ9fzpaFodPxdXnp5KBpL67TVlKGQdvclfOiRpUsrskQk4LpK35
u1IQvTVu36xmniQY/3hfpbsVwW8/HbKma13W6skazhjTiHRuyZIjp6aSa4DbfODm6T3+wWe/JUCP
b6hiJQemnLynnOtrsoI7aL5upWnlexnxxU+t2yqoIIdqBo0QCyU6/hvdch6BhEPJuCtqMGSLZ46P
JuJbfdPLnjjVWHToLwxop5Ueu9mfkYeTGaHyub1pOR8r3/sD74xSrkX4ILJcjaoa7oU4KsGanv9W
297pi2kDUuI3oCTVh2jD37+dc/0zNZ4JXpH37NTu+kAGvxC+rbG8UJJ4W3ZpTb22l6rLUOhAEqbg
JnwKD8n1bHrFh/4vdBka4bWB0+wyHgqV9cQAz5NHFttOwP02tHIXwVM7T3ueO7FPFDFiVgtRYmj4
hkCir24tXaZ+x0FxLwJoGjRtnXfA6zegZM63yxA6kOSCdiVsdIzWTWVdVUyOYKuJMQE3WTfSLBOA
+E6+33KU14opBNuIGFL0EFAWqR9tQxFVpG9l/QvAfibAXDFfpHH9gHmX1jjCgRAZdzhJj04Lti6v
vebGj5j0hjm2+v6kfNiC9YU3gP0cTRyFwDi5O5MVMudB0KvGEdRsK3vMRIgVrkDU53kHHAbwxICo
67K1VoJtDW8tVcroPcjFJ4uH3jK10DLKIhb1aAwqs3yYNWHNzE85x6OfoM3Ikga3wk3hOi+E1Y3S
IE3aLCVRpqHY+nNYxudPy+AG+EmxIgqgfKZ02RPidYWF5atsis6cQexFKa3vVqiEnvXlrw7tHizt
0o4ayBIQvx3/ZG0v9jd7FQ2CHJYBpL0faDZh5ymzVZFau9zZtJ5WU3OfTTV75YOsQTDughGdKico
C4SCMOQOGpEXAIkaErxpKfht0lqPUSDPveST4d+7YU7GHGU5hms8Z8hTGcJinPdmEpj8j6iBW/XF
FFeL91J5Wdg1YzwxDTYVflrkXvTiYhqC1SwPcEhdGgzI1ftRI7ji90g2icTFbYC+5Sxqkoma/Gkh
s7X6lmKKIJUfwAx5Spr7LEz8DMu6p1SD5IcMKXQB3TTyDNos1Bjehncj1udm7IN4C4x91Mo7z+nF
mgB0m+V4TSXy/34aYqT0CJVKcgI3twnLhNPFnEcefEhkTkxLqCVBV93W/J0v9kWbyVz0a65xqvE4
5L4JaFbyhrg1zF3yvgxrQVuvchwMETjpSJa9sn4zewGrjkAQt+A4VpBXFGPl9ZHdT9Yn29KcC1JY
CF859zue/cAbs2NQngbNidoISxYjHAZEYRtIZtxjAHqqnQJJq6Y6JTT2ijJW4QzqC2dcVqUyUL7x
KDq9GLGOVA+JCtFYYuw2AcF4gHTx7XO5MB8Nih40lI7GUSsz3u9+K087C6ldR6d2scVzeYidmnjm
vS0WypXGjF2jAbNFYL5AIm8YxBWsU8Kn0doolDTTNTZk+TebTj69F3HvVO4UiWlRQlEr17hUieTO
8cwt9VRhL8i0Sr76eHd5iDNLBoisRVLjC2mZ+z9HdXWAUy2SPVm+lacpcywLLNFppGjuD6Mvnrn9
8ZPCUx26wbOaiI6j6Fo0i1mj5G5Gc/Kw3rRFgTBss46oUU4/2XGnc9dejJ3rIoC/a+rBGsJIOa7v
b9X4/8PNtYn3gSKRUHQ0BB+8FEZxaF53zsRjJSDRR7RBIYTupmueA8ZD4P5+gB7fd28rIqbWTbRg
yJoZVsT53KHTcybAPgtsFJrcMsWI9nWsfH//KPOMVbJmwnU+r6cMBWs8SMaEvLBI1nZj3BYh8IEY
TP2I/w30R/ksOrdWD6DhChbJKbZzsg+MWy9ZzfBvNiurnCxQ4DM1vzQkx8rEh8u/dFDiyhPhYg2P
792K38GRYPZYwONuU84Ugo0D4n45FbmsTWJUhylH5uFkDW3q0MloLr8hnFoGtN2wqg7dr8ZyAL2/
kZCTHnmjBdR1Anx7zwq1a9KakMgrJh1YRrDaA3CeAM1M9EoJqYSfgnkADoukyfIDf8CesZb3VvJF
otLyUJTr/U4JX5714enM4JNT6jNS6jhk/is+zOUp2D7hIPQ2uvQ2TVWKdSy7XdC+i6R/Yr+sjKJy
NV5iMqlRd7D5auGp6Y5euYSqcA9qfOTmdkpZDCzTY8LRtYfD4cba4KqfyyaVjgNdqLh+HvaAkFU9
DJgz/n/9BVWheecPbJvcmz0e4tl1LiwQMCTFuPLXXsxkYNVwYrn9iMO6oQxziR8kZ5x10BwWteY0
EBpiE+smtvEYYKSWuCmBIOrP93ndWyjk4ywfOONpsYtUqBDdbftP2mnku/J/AZ/ujzWpg9TeCQlr
SaOLgRdJK4BkNkd+jRmQSTb53uUsw+OJ/AlAaZAmPXHUMtJP1BVMjBUu3RagNFkNpfLxrJinyyQy
X2jyHjpwtFCpojk+4cYnSH0H8AmIhOSsoDoRetlhwby5qrfAltdEzXLwySbeXIZDCXkbkBsBPCyF
jmc1UmEbl5nUh10mmBMneHX4nS/voLv1ShLy+u92Bueqf0HBlwRQCTENZR8R3eQl2lBkD5EmOHDw
i1bPbhI8hLMXXVZHx4HHOmPW0ysipmf56YwU+w+5ro6mhM06kSdzRlgjOpkpao47bGtUColwJrGN
qmLYVNyTrIGWOO6w/CvHoitguBk5/lIlaXoj7LX8zFHeK1uGiZ6bS0mlxmwZkHB9g91njrXnkPU7
C/qivpLOjwoj3YbVFYjcVsz8nvQGnr+uAY/yZVCnst45RGH5donrVdUTudfHSjmDizBAif1PHVi3
knW8pqX/YBIccK9Yy3o/XM7OfWoxZd/1h02bwrmnMfCKJWW7WpgX5TX7/iiWYvkM9rmhnm+rhv1H
YwaNAos7hUL/zC4XfovqRbFSz2JfhyZdq6anK4wckzfjvRv90kM3L6dmDyFLLfZEFH77/984oXIl
FGtvrL430lvT2pX0c0o4cN3hOg13o+sfuNf6mXB1CgpqVb7koU7TXmAY1HTuT6kkgkf7ekxoBp89
+REuXUepyas3+NDMcvojKUpYxWn+ofIGIaAtS8O2RT4oar/bdkmqgHwibTqYJG7Mw26UUZm4/rBG
p4Bg6J3D3kHVM8MUMkPfBSUn3qlvIV+b8P3Y9UYeQz520IvXxsSqnWL5ySpBzE/H1wJYcjco/JXp
9wVgya/OWRLt54hm5o0QgNQc52hqPnjk9A+0htOYRDPllLgwFtjVnktiJ82h358b0V+MbmPYvbLe
GHHis1japDNUzZ8Tb4dQuPyAev+f7ycrF3iF/dSUkssq5rsp8G/HHSCTEiH8pCxbMLefXb7AGBT4
Q8fLU7P9ygdPedF9+P2FJi5IWMSxXrs3wiBUmsVVX42hAJLZtkVP+627Z5rd9rlKB8MIqqUKD/wc
1LdmtONfKqa8Q+gr+dFwMBZK9ylf2WpZLhCWyrnvg/IIgC5VkxVrynRT7EShRzktv1WkF1JjeCao
jHYDGymYnxEhLbkaGKRV9HOHkUY284zetUB6uLHAS12iA02YAoP51vuelxB5bM9ctT9UfHZ1K432
LYgXDLFhJC8LJIlscVJmF1eowPYc/v3c0tDkO11K5TJot3ghvDkbleyy1A3hJdIYV7gzy4hyXHRS
w+d8+uIpgrR7pucXlrrLhrEIkmOtg+QToi4M/J8E4phk+bv34RlfpItKX/tLz47SkOC2IZQgOEG4
Sqeba8FOl3FF23VimLGncB2wk3fq0DebAAqi1XQ52wOYWs3NZ0mgo/UI6qDalx0Y6Dcbwx9xpXO4
BGimroxAGetSyqGsDU7Zby4EOAfPpsTYBbu6CAQUjd5nikYvZm7AZsoJer4FaM8FGFLueteLozDD
qLe0xR8PvF/jtuC/eqXlWlOwrMzDyq4pO0Tr5RZ/9FlG+3ErjCWTSYNVz6lHnHCkXvitKyj37u4X
USmok8BdcUV6mB4I6ocEhLybY184Ta8QF8AP8OnLruHO158X4Ar0naoyZJEnNfyhvTs7Q3ep8nZ6
bTSs0YkYyjvijQpTbZgUEWSg9CRcPMm0xzpirGg5Iwkg+gSH0fZ/jLZpzJJ92M0oiyvo+1fFMGoi
yEeDrVNTNRQtb4auHzrPRUpq0UZV7zrJG0u5yunTVotduvgC/tlSdECWyauVpG4mglTBC2JDrW/M
imgxQk3ePfcqMmLpf73dfGRenPUaGBCMliVYCufwi91K5JX63yORQAlREjmOtNmdQcx0c9jfR9iG
YlvZOT9z1w25JCZD+zmYcnnZd3Unyk7+/xdRr17Ovsx/qbT4Awx4YElgffzwJPOls6pYEziGT6N7
VnP7IQ6Btdj/YXsc4wldDunPAfDFOPM1xvgVyLwfBbUhoiXzFpgJelokQBcGtvTfteyBq0TCPcqo
XnKa1gtnflEScuiV89so51jXNObATdUQ7H0DNXNxaqdOPV/lrnBDxmV2sdsVnYedRs8T4mhj3VZ7
VqtZLIY2SyspXK2Wuj32b9TwY/IjHiBDG9yE3olYpJ2jMT9ct3HS330EGQpmSrrXSeqZIo4EntBc
S1wVWrEDtSmM20+R4Vfw9Gmdxm1xEWktfsMWbHyMPq0fBn2y00A7TFBE6YpqiTBgIV4x7DARSWwx
MED21czVQ6fdI0IZYXjgeDsj0v60jgA1hPmHjenQPLv4xTys5i3x9ZYOH26VMULF7Si6m3kY+Jfq
UoiwT6pi7y94Tq2KvF77kSLa0dnN0/nZY7j3rH/r0H/cynM1Rbz41gKZEaFFwAo7RV5GcOSLk+Sn
w/6/0PPG08V06gvJ2/tWLDjgwrjgREWRGSvHkKwSj+cvJwYKFnrHNGkM2R+tdHZrowwTnTk/dpgf
FxT0io8Hgxi/MVX96ntJbI443t2QlWsg/pAwj0GZ/E5NaSbPkIoT78UVNTWSAVc6uUzczGvq5KZh
r4uxAuSdeYip6GjciqVeqZxACSnI2dwRnyXBi08yv7y4JkCP9goBWPJLtwG34evGf+Dx7iNld2k6
g5IjjeiNQZoXTztAbK3UnlIMMkZctsQkcr//2T6ZGKR6ZQNjrXhF1yYwX8QRGSbjgilnBT3VoSFN
wtX6e3I+HwJRRzQeE4FpL8ybst/obGTYsL35tkuztDTAlxSVJnu1vKVqgZGbtlSrw5Az62cguTt+
zPu2V7kViR644NAI3f4paPXmSLQHB5kdVUXsX6gXLFt3t4UgK7N/Bgv5mmF90dkLn/2fpTPbsSIa
CigiXY/2a1DMfQuIlyq+SO2N68xqqBOAUfJPJ650IpxQfVXaIRVgJ3YlCQmuhDtpcuqfi8cYTFX8
AE2K2dovPfXuk9Y4SzMckiU0J02lfPjfu7DNkgP7SwXSQtdgkD76p+zp81bS7Sy2OAYGVLYLf/q4
QmkaUDL3/1CxZeS4StPHRvcG4v3llmH6yR7RazcAhbUgTiMl81pDoNvWpuu9qqs+S3ac0wdDcSSp
sqy5Xtabh3EafP47s41qcdPrwWqVx00Y/b0Q3jgTVtpcDo28MFroz4nJM5kU9JKEy1mJCAaI6Yvu
/70taq8zpEZIO6L6ZMq+gXVecpzsqQJ//IDQY9p2RPr+7lihmhzN4BZ9FYshRqfyxVl8tpk/ylBY
XfIO7iRjypnFzpO64O/OHAb+eCXfA2ZS9i550WCUJr4uDAeUC9pGUR7pKKruW9rMdwHzyRRFXR1M
ST258zLwmeViM8owJUau0nKLuNMqtqHmCbAGaNJY2x2qnvsyKhozN6W88qs48zNLHtvQv/mCtxsa
lYYgtlhCpKY59dimGXy6acFK3vYmE2/nqRMIQyxuZl1EsMfAvD+BQuYa5VzWORM9sqOvsmh1NBQT
GXvfOoW+pIGnjB+3swUwwVRQcn2alkrPRTKJiMaK0LnC49YzVNSUs5gM7Ln+s+bAo9O4PxEud3M/
k1oj4bBz8LGx111NHz0NpjKqgjqtTvXTM1hktL3x59vDY+UsJ603+WND/4ygwtvoBkGlEMYiXxE+
tIdGb3f9UbXuBwh6dkUtWYOQpz9xGTcYI9xT4fyzAb48h0j+oUs1MauQZ+1UUjXV+zw8MEfRpj34
tYqXZpH3CP1UMg4sgPzTVXr04uTP1F1rACbNmERNljVtBUOcfT4l6gaK7pBLygYAh+qQhzMBCZaX
NjzU0P0zSjN60ni9v+1lUriKFGETS+1An8K8ZnTgwpSWfdyJZU5MNFhGfiDjTcOEqInMIgHNNKse
QRyttmJtHABnt1ubm3z5JXW7TyjEaDFbqTovtw5ByCaCCsHgyqz+t20b9hmc46iTMALYTCPak5V/
uKRrmJUByuBRFCS8lMdJyoagYdnbbq+dSgqoHUGqrKQ9NoQF0+0+qTK27+yRs0dbnYKZdjyF5Vf3
qc5fkSfXe/BF5aAYWn6MwadjhN5OGF1+yX0on4B3hDI7G79u0usBuBatAekjjvcvt0e6bhC4yfue
yEDcfm1e5NGGXOXUgX+7+8M26jO14XdUfZ9BIqVycg+mFBK8aBFvGlNZNzGJ4Bdv9O5fOyeQdF8Z
iin7wsSumARYh/po0mp+sIEbNKPR4xceDH3EOxpgqzR7XrxyBs64zfT/C+y4/jcIu7mWvtEJCMqF
7yjrLkBaxUx4K5KmF9qRkxb6QBE9WMfN4TdxxmFsi7FhOMiY2nCr64qVTai4B83GI8GK4Ad+pEyk
Ji8E62BJ6WwbqoChj16/6bhyPlVPUXkLdwDQCjK8u8S+coao0oG3mVNeAecjCxlj/abByGYl3HSO
RB4GvwJfUV4aFVEjKxk7+BlWyJMu7ru2QKIr0w+Jv/iQaefTaYjIe7syMQpFWNUK+gO3aQqcPEDD
eMpVIfgco/Qz83Y9TlMjgGeGDp21Cmg3ZOmyOXYJ8FnW4fTqTqozUdcGTmbNnEhJeb3zrJ9adUu/
B82a3aqj4AiLQDFC1NJgDipbVWqNx3yDwfiwNG1LT9SJBNonolg47jI8Fl0Md5RJ7GPLgdmul4Xv
JnwkncuZkQ7F+lBgp8UNEB0mFx5QIqHzzPxIbzxpIlwkFHzxd6iV1L/RCDvcZv5CnSB6fbT3dNuq
49PpJNvsqQH5oLeUwcsfqcyrEmyGH/O1TS6hgbWrdboH8KSycfll996yQxhADG4W1wBgqB9daiSc
3ZRRrs3Q35YdAGMbwTnb8xj7kdVGoIeoSDp7A5UN+d0fP/fvkuH+64zg/YG9KlKJkBcTpmN3aUFd
ZShK+j2MzfI2h8mEAo67I9UiETChifl7JXsFTMOeHiNpFN7vU3hCmT2QBsMwTQgl5v1Qaj4yaO87
cBqnz6db0IlMI/v1jkynHrXY+gU8WwlclrrG1sNzESY3VO1gT0n4pHIDNpRAIUlc+RToH/gTSYln
OFJkWQrVSQFAioyrPdVnqmg7FFe4kuoSea6pmqalxy+3WGQLq6YtaggC/BxgOGfrGQCtfVu+fXDn
gzUBMNfHdR6jSBtIXYcpyRRJYut3ktLdLydUxz9RfIGCd9OomnQ7JHpkMi0WbSXJXOJOdcJtj+8i
UZm+pJcSN+bH7rA3qjb1pkeqsKn69Omo81fSfZFdehhbE+owaDknhcbIK/spekxxJ/o4OnvXVbsf
MVG0SDeafznk8U9d2VeXpOO6HgnwfvppuRxzwVPJK4grVQmnH9+qxSgEXt7UpTZI3hwivjV9uxUh
yceuaKg+BJk1abcvBWlV0P6J86mTpkKQC4x/8ZMgy2DHh0zJaDWk1VciggdcNMf40jNnZu3M59UZ
aOg2aCvKPq12FvyY+iVJKNQJ0OBUOz7u/+i5J/8p0Db8IdFRTPaeoHu/SuaV3gV9UJIIxLSHV9uT
WzBgY8DWG1lDNaHly4pcQHv4WSlrIRemJNn8kkV3o97W0AS2RhS3yyzN/aeVdui6wIc42OAnCovt
caoILLv7x8M6bbUpCo2Ykrkx6GCi9DXck9A9yLSUMAmfXdXItJmczN/Uin8xJX36oRQX1Pm2n4Nc
byv/1x4SO6NFqluMdSa/c8cNY+1xmUkmKfKFYRL9l5+skeR5TDyRaUPDc7A4PV+yP8c51EHrW4+f
zIPGsb+IsyWxVs4lRGBNMfHToW3m3SY7BO4zU7Hg5qM8/6CKxWLp6M6od3z0TXzDe4lTYUTbT237
J/Hm2tZbkE75bfoPXEhspH596s2x036xt4+oZXYmNl9eQra8ntbmNwrRyt60LYSt62hHTCuqhOdD
LGp0BcCfujsI3Px5nZ5XfT449fFjWZDoPebVOA8EdS5WzzUmu6Bxvz0Evpl/FfqenXuffNcpdejd
FlonOVkoTWOU+DC954tH/BpnHBxNyGcFXOPtSOgpFpDxlKPSHlDGURpeXJ/H7/lByMU8tNZCZKFX
LOu35Iz12pFIuV59JmtLLgB8uZeeP/mAeIjTfnTRjj1yrHkUPaMfbmq34MGA3BpOjE63CbEpwxsm
CvKxGW2ASaYNJpvZw4DZSdZw1VbVk8l+cg/yApBL8qY9t99mRph/+xgCL2y6s1YXY5I5BNCxD7nZ
ckiw3J9ybHiAIkxiwDy7imtfzFn/wQY7NOvjk2ubwwBLm9EZ72g7B6FVOXm1CF1v1C1b915GwDVU
dSzjuZBowoU1hupkuKhPsDsLmPXzoqN1o0d7caCn39OlpZJg47HYw24NxiK5jOuOiTLGqNc19wO+
ZBcYYsyO6QI2X6TP7/Iv28LPhn1HASVkRVVDE9YQacLGON5jd2Wbp9bOVgY246RRiJOiaE86swyI
x1nx/RLmWw3W95v50tyG3bYpTs+4e8B1nTqO+M+kjucNbXg8gePgPYhynmSY1vO/pCvgwmKTg6+L
7XR5XPdgODSCenIfPusG9saaC60/CqGi/Fhd5xRaeg3AssuauKOt6Ex1FzLIT7Uwf5F6U8eRNLz6
T1dHulNOA07djjt6pfx4jr4VQbyQdwbxlCRa6YDBzCSwVfoVpITYNA2AsZB7cQNY8kwtOSxpfU//
oX2GeuUcqJBeMN5cdlbMasPiSiQgXn+ZMTydO+4jasmz04By7XkO9uUrYSMOEMi4Wr7a6iXfgkOX
qr5dCp8aCHEbkpp/xFN30kEa7S0C1WXMHQ7Fx2leHGI2RtiglGqzcGh6FKAVtQ8hRsl9GiWMAM7E
ksO1kALtuigmyTHEnkTh1x0oQqn47q9OldjJj9ERl0fPFHgYR56bB7osEiv/n6qpCuSaoDy0qS5t
/mp4E3gHYjwzrs1jyIlbOqQ6nPpZ4xOh9qkc2McpSV6MEW6xrIqaClM1EhSDGy84erhpkvwSUR9b
NuBzhgFgNKYYVLYjAX9U+FMUCX31dBcqnDwUvOljjy+a/bCYn48Jz1tkrsN4+6+EUSS7gA3SmWSp
gKbGEeC7SN56LmiD3ssXVTCkEKGCVoc32rN9Zc1de02ALTec6jSMCLvxvVb7iFYfyA0VhSWJEdu9
oWVhN9NEk6oIanfAyDr0xS9MgeIRNcQ3cepmssfXnRjKu332Tqk+w/7MlQGbAUO0if5mbhNQNBHN
owqXYP0Ejh0zRPgR5BmWIJd/lQ2aSsCDqqHZfbgLywwZHeV9nJy98iD4mLUYgNmSmeY6XJPNr//z
oeqR01QmaoiXxVsjZ/ltcuqAiKv1inKfSEJrru/b4d1f+cDeF2DHiFY1DtzNnQxkK6YY4+iAIEQi
6qWpDidmNTqIawe+ZBVmPtqV1eww+lU4DtpA9zjaazfS08zvHeYJ0M7AfnG6cpZN0FTLlNiq+sFx
8mRWwg2aIKKvZxqAISdxKHiYGHZy6YF+AfztaD97Q2dl3sLyEy1Nvfkstl92kuwiddFa6DTgJQJQ
zQbPah1D9Zhbx51589ADF5fkgEYC/D/9jZ+fEXPFuRW8TuXvrFU0VgQ7KQI7bl96EcRmzv0Qryan
w71u76iWLeRdz/eV64HFyQ5VYjJKGJtRnAmyy5asHU4VT+DC7rUx2O0IVKaOjQB9XvfwVoudMkWY
t/Kwp+U1wtEVwzCMG6YwhYrw2Fv2WZkZS9XlTWOy6TU7AkDwl6amninSBkBHexiK0U3cH4tqcaJz
8CNVcLnN1Id5ONuEWo6LM/KKVOLZ9Ha87GJR1oC0lI0Bq5rCaUbrej6efBxa4ntHaYvvlSO1F94J
mDFvGFpxceW4LfwI50WGQ1p54uAgNtcF48HvXNTyrH6EZcqPwi8jtLwKvRgPOQWmSkTCu7ZGAWqg
Q8JvhF+gKjSN5OcB8cHcd6hKh2tlchpPBc1oky7xKc6zWLln+nlrvq6zjJv2g7Ktx2yVA4/A1Ljh
lj55fQz0FuMmmchJ7VhY54DD1LfIyrhaK751MdeTNhMEtkqQUlZ1MiIFbH6YOI7QbrllZaSt/S6a
DxYK2bAPt11PmAEddCzPTr11j7iV1Oh6Ei5bjrHvG5I+Y6Asvw5i8mVh4J1WoBUAHnnWq4NsWJdY
BPekUa7JmfgqcgqJGljC6cTNtWvJfFR7CVI23+z4135loXd11Nd1FMqVfvWVr79vtzT34KSuyWkF
FfM7DK7Sb3EHzOVMe1x7StLnxiHTfQD2N+jgN8+SKNbf7zBsDUueEDbKpDQFii9DQklUK9i2LdVP
+xcNQw/TWX3hkLNjk0mGGgDTFODQgqASE7YPysTPOD3N2P5YZEGIXlLTHCzkOJotQQS9XAQALk/S
A7OQvoTXoZoaH7bSh+/d7irocFamel3ta2TpNGqhI67IBAGYNEPnkGlEm834fYC33CIYe5/01ShX
y469xVQd/myhlEXz7mLU/E3pG+gtLOWPRNaInUwdsfHv2zTkvO87gWYntVJmqTHrj83LrJRpvqws
+EFDu054Qx+NaBc+VCEt34H9dOPy3gJ708mEDUPrXia9MwTpadkRo4P77nqiwNuftazCDjuFdhp9
OJUvwSztEog0FwsCMOB6aWOWEAf8DYeNensDGpxuAbqSyYhOfMKf2+Xl5y/+bKYVab0y+EUl0Ns9
aFNncWqimoeg554QNHzAqiszCbrRwTuXZaEPuv6g7PCJ7tbogxndxUzyMmTo66OLlKtfcWjfGjil
WSRZIv7mNFb/H5jUA+5VemdqUwp06Os8uGY/f/vgkVT8+UyJYL39Dh/TZkxlECIdaH/BZOIvO/0i
EWBoLSAYVYztvmqihyIl4pNFXL3dAeLGvvn8pMfHD+NWbE8dMpK3QJvLOBoptz+TBw4Y6jm5Ww9r
BuzLxMO+hzIKErzlqQKv/7VKRLFnsqdhRgP5tmnhFDTf7OoWQCkHNPEHd3wt0PZFYUySNkEV497x
w8Xjx6LUrvtMS0DTLfgWAOm7NZjavJqAgUkosN24xeQAVT0U7mK2rcTpxaR8LqTI2LAWvODY/Oy7
s3L4yk3UD0NIonAZRqneKW8BhM261EOV8H7Wcn5BhGJIrPzvpqfgPeGOX8AA8fjhObVQ7X480yKX
LiWJ/UfIDz+gTeUmI5SMX9TyYiXB60/lTDMIuibJfrVould6QztVNxjWTbXpkl+GN1czzu/rY2Lt
1ENmLLPQxO0MkQQGi1tSwVUEc40cNSY6Kshej59NjsVCWckIX2KOCg4cE3oQPvz4LTUiLlJDaGBO
ZJRcBV0JaDQDdztGtbFZTv50KM6ynpOaTKKEdmkbxOw/ocwi7tG6UhPNmhhD+OVoZVxepjbkzKcd
bvqrhrlf+fJ3fhvjDrLFCZcX5OwLVYwfd1ci8YzmfzEn5GLFMCuhuX6kxG1yeLVNtFPBFK4NKoaI
gSz+CIN9Bolx3aVmjeZgESVPesLkj9nAUfpUt3r+TG2E2V+EAEEHd7mlvrJ8O/J+6hC6f/pyiXLn
cc9JNQldwE1rG0Rqkllcgf++QuEbcJtRam/TS9pLL1LAGZZ41ZhWEVQDYoflOZvQTkHxu29h5YRT
pAelZg/QgqS0u/KPVczxgsfF/rH7cGcpCcPql/iGD1ez4nKx8FH7c2z5PlVuwLflwMB3Ui3YXQd6
Yrs318qa3lQwtSJ0hmdTM+mjxZlwRlQKtE2tCYySP7aNtl8WU1cpg2PHGMHGeCEJitzRda7TILzo
VlJYZuu0xrQTb/lymTWmd4wWrx2S1bm9jwYBdwnL5SJpZGTgHeF+monOh08mg/94wKwhcO1C4qAV
OfhxFiLTqzFHz414IIx/VntE1hvQIXgKoBbJv0J5R2Qx3hm/D7Ly2X3E+ucnne/c9PDe8GMk5vMA
heZ3Spu1yc7ydxtUQGbDjPMwbGA6fuwC0cg9zm3XCNgpgs46AdJOiF6wFnkzmT1WH7Kutq36mZRA
I3HqD7OJDXIkjr5ZjBqlnDvCtPq7a5U6N3eP3ZUx3DBLzHtcn+g8E5fXvVxjjjSsEQLKUWj4K9E8
M9jHlbDNNJUvmwRPIBIWcQp++ZAg0zUe/HWM/H+gYo4qD5wV+roqj8podqNybYodA3oTClfSlCdd
YlDKXAxCsqqtyy4mTXTWwcqmRPrMKsENzWLRC1RlD3lxq2DV0/rX0QyOyxheVWsX3sy3/OYbv144
xrNaWACabbpHly8XawShBFHO6IsZETda1SCkvAl6zLJvtsV/jchWaGdr7bj/6QkidlyG6QAkIhTm
1gAW3JkETLS7YOu6tq4geF6D+Is9UsUAsnD0JiIjnSDjyDQKeST4b/ZDU88iASo0Fg2tHH8/f1np
EXV6T9aYNIOs5JGMsy0bTgGxa6ipNdY1yx6NIpUa433PcAuFkBIx03SYR4DMAAKWwwbiDgOWVGRq
TyxDsE223xqXL3J17bCM0BFMt5o4TFdzvSQDHQ1XdY2Ajzp7q31xwRiwWoRKmqjcYQFZ1tkxc/fj
meF38bhoi7HWHlWBfn99LWZ7AWXuFZNRjM7mvKjq8MqYytOFVBuJNKcW3hqYNf7b31q8q8vv3zQ3
wcelONioC50uOED/1fbDhuIHoXvkVFjyyq3P6xjy2pJvFPiIh6xkb6a+0LB6B++euk6qZh3HeEao
x1wSiQRfYVDQf/jKVklgw4vOqSAToxerqLYFx5okpkctBcm9oGctCUSxrpu2XVCnOkbvSdHWuhaO
9MLJqT979mlkJwXKuVKkgUKXSOHTpdLhiotAwEpoYSLy+qVT74eyKVe2SyRe/0r/ZJ6ch2hRYMq/
1CnA62b1Ftcxc5TFQuPEYMza8FzfPZ2h9s60NhJVw20FyGxalc3+PUiPdnn0ToOxwa7rsuI86qUD
hLA0o6hutJrDd2YjZfz5J9pxG4HHnhXJwrCxa+Xhm+qh/Yg0AsZ4KsLsNC1QsQw21+emSMri/CHg
ZnGTSwqyVP/1ej8Jre9Gz1+iNNbwJmJECGE6itIAN39MeCL48/yKo38pkHFpL3VpTNTkIRDYmpLM
oliCoNrdy3WaqutMebKVm+VABidlzG5PLgOTKxJ+XSg3QShocnRmkPgnJ213rpFyw5q9zmhpNNw0
GVgaZnkcpHEoTvlrExiqivULrrC8eeS2mLjvF4lB/+nrHfrPTFatJh0KUnxKnWWAgdCjaM/CS0dj
dT2LYATiYLJQTmYLFfdntOHxRuatfVEkiWb2Hieop5pmNdG3Um5cHwt2mo66PNyK0NYDFczHW4fc
LV1OYB1Glq08+UoY+6Wc3tB5zYsEBWYRcfD0kPVFvOoYj+Z5dY0vngIQ4mbmzW6OGFpnPHfNBa7q
hcAyczHnTqboTamTCe/tJ60ttW/k4Ez8j3pEQ+YUjkxApa8nXJYwl266U2wnQsTWsEUk2RiFVmo+
i7V8SxxTSZxFCgfGtb8eQnNlmN2V6ERwFUW/z0MPl5tUXtmDHPDEnYdWiv9RbOIVBxTGTiGdDoU/
t7egunaiFKGZuODs7G8blLhjkD9iG4OlPtLOfJtcuInwBJ+t0UP+xROVT/GiryOF6zCVCxoqEQOd
/YNNuJxj7muXLRhFMH96b74u6wDsBhn8WnuA3I0AqF7P5p7Vl2qf1/A15SI0KnS/tfiscFc+Fotq
9DfpcIj3Ce4jaRCNJJV7iEqHnaZmFSaUvpBT7z14ibLbaqk/qensJOCads7tXuPK8+lZgmHU8Ywa
oG/yrBuI9ZFb57W3ijrYpJhbJtzz3kGAZFTlbLeNgK4w7EFekRod57CSY5oVKdvpKE0sYYqqgUJh
HVkCOXvXbxok+OLXab5Jl6kE1crpCBwZEbTw7LXVZTHwlcgsqd1IvS6xvfj/qUxavDIxwLsRl42h
7BWMpytCEh1Z3joiykHpAfUR87GMWVkm8nkLV3lH04B+aSUXyw9U4sUIFtSJEzTLtdwjGDJFELjU
CGb36LJTbNDOy76UHb4F3XUmmczC1yyp8nff5zETmthHsvgoUi06LXN77ktgoZwybeJql2YeiFhA
wRLon9Jo2ThOQkJ6mF+rbfphWDiWDBn7DZK7VLNyFUROXwx3+pASP6/uWQ66g8YacqjjOSz4vmgR
1dSpm7AEaKS9CdDuHnsF7+ThoOiP9VNCoqrcG5XgYn5y8/xEtsD5e4Ygfhtv8sAkFrsXX3xvr7Gx
X/g+EO9y5nLjGjgz5jWq+M5l3U4BdxAjLHaxTwV74lP0OkRxi7oFU4EJ7eJNF0HkS4J6VhwBcNch
74/od8ov/AlcSX57H9+ZC310zHdoiVYjVEm5nLUYWiWEXrnt2J2KI7VoPQU5ZNG682CEiBzh65th
4g0X2qjwFDQG6UwZjy2ctpI0n8i0gqTrJyDBzcm1cVYzqT2IFm54NDSyA/ayL+pc6+solXfbE6Ss
Gev6yWOX2idW6cyJ0dRdpz+Kxg/11tEVP0bgCFHcLX9HDasC3VopFO6Uy7jCDccFC3QItpxjDwLE
3Uzv35Ismt8jkRggJ3Xx78hNiXjrSjmOhMOOcxz39eFQAu7A+YLtBP0nLP4a4wPDhe/f8aSQ8ZxS
N9M1wcP4Klt9Nyn1i2Q+BlDUQ2YdPzFtfQnoKC1vHhm+T//S4wo0+Gb+Z3YCyjt54ejaaQL03I8X
ELJs0sozqffptU6tA4yUVhloTwL9ksDYY3IjlqQtlPVsDx+tGLkFMAV4iLIKHYCZG5B8eg71BHbv
v1wB78i6dm++hxcoCd8CMuSYH1g0sRaXqCghI9LUEVvkyo01BZrb8SJkdeAvSozGo6zNYPDd8uzM
uVu835HrN4Tjl4NzOiqRwTVRjlcTaLq4J6hTMq2LNFZvYSLgm9rh8U6tMUEiDiwh5OMHO9Cu6hQ4
yjRR69Xa1n8hJhNn99sucHCcQCWq3N2jaj2w8VAYNdZVIgRnE5kj/SKRFYA6njLjn4+KVHAP2tuQ
57x+wAX+7H4qJrbXTLYURGyK8bSHMbfM9vORmMuLQ5upN9nnivbmQOW9Grg2ATPi4mlaqTCXDg/0
iSaTG4WmBhISxOfppMaaQt/RK8m+Zc9dq81yEx09B/Fc2l82WZTvd7nFAELtzrs2lK+gUnrVZ778
ha/nx2X7u3n/XqERZSxVw7VZYHQZCPrtLz7/2Z7ktnzRTHvXSVThMqkaoNofWF4lEyrAOzWrW9Op
b72QCfabPEPzbS8arOjlo+o0vkKBxvSJ9jSDSKyqexYsq7xA6zfTzSRmbRWDTRbJyFpiap1DB5hw
h5f/UXLoN5YtBx2901uJNpt1Sb8++S6jWsIxyZe3eJW+EIq3iCRhlXPDmGujw5kITjkhpNX8T8Uq
bLNe7FgIf07sSJ8f23R1GUQJK4xqX2hUQ7u9rPsq4pJ3pfit4xaAiUnMMEPjQQlmtSTlZc/tDJPQ
a5MJln2i2SKeKAbnPR19rdx9Srk80ZklsCRq1Klv26cUrCtgTQwAkokK1/vTgPwQzOVsr18m+g/d
ArNa1VbusLEzUCcbZyBoDf0uXxFd98h2sWmuNa1uBbUsHzZr+rMRlNPHWkjx8ra0DL6iY9gsFC5l
pxi6MiNGnDAktgG8BEUnVeXmwIKmgdtcKRCaxMtfbBit26tNuQoYvGBnLBB9lZ0jqd2FMfWrO7NL
I8d/ejT8Dqce83EReA2LOkkHSuqJ5Xiuu/u0wFZNktyko1SFzVY6Oi/eaT2wwJO4u/ZwGwHHPIgs
CoTdkzEe8/stQCWzNhBTW/L2n1iy9wHVZD+DBj4DtixYCazgy3lWiXn4GxAg5CHnq82XzXY7wgJY
GqmuP1ERWKu3IBpE/f6LdJ380BaZT0Jxr07ogJuoTAhuetougSIcOr9s05aBuUaDyuc53Av0Evjl
9uh1pwZjiYug9ifyga2eBs1whTpfUF/d7Mbhg60tiQxi9jT6+nPGoDc1U3br2TZXKRmAF7nhi7fH
EWckQd5TXNgWHOOC6etiVpsSEFrtBZBpABtRYvO2ndBppi0VfCgnRLhHKg8jGUCT7Kc3NJqJ+Gtp
qA/gv4dPmCd/aM5XuE3YaZylxIE5Ryx90i3kUvVacXWL/JF1FEPhDMqWj6SyxJOBmzuOzbfNX2jm
fxQyXuUkn10wlpXocyUI7xeuA2cqWWnWG0H3Yk4cQYoqbjBb9XwQwcmmYLSY5I5I/l2hSzmo8fgZ
yG4YpoWpWBQoHiUd6CrEQldppj0qT8TSd8y3zJQYL3AePrY6T7vcs+iLOUFnw6ENOqBIDa30eJj/
iGfix8KipOBzMZIhCfH4oZV0kTSl8m7hQWpY2CIrw4VAOvDum7f06sPO++ZE0gR4grbCLgGycs4f
lXYZzZdpoYMo33CbdRS7KZbpS1SkJEhN93sRO7h1l8LpcTGr8AFNA6y12pQu1BU2O52q9tbx4u9L
2F3R56Sg/z3ztkr1gIE0avCVhuek3eV8xhUyefcnoMTRz0UcJgk2zSOV03u2te8Z3Deaufpde2k8
kuNjZ5uVmbRWUOW0IBParlc9ndN9glEpOfEwCcMQrct6sLZYq1a8SqtGj7tsSeJZBHytAEYGJ+Su
+50mT6hskpUQZm1H78C8T+G/uGMJi+YP6IStNyC++9HdldRcyuvRZKTt419S6dhss1bFovzjbk8m
LvRvL2dgXiQ2n8S+2L/nFoCjf44/CqK79ZDEgZs6IJBiw8S+79nhcLnPn3qEWT34Pgbfwe8OMY4k
p29eqa3x4q4rIUacX1FNjzfiB3JFsxOZa9gfYYjEveDoKaen1PaloGbd6H24XC2cVkgIaUksKGT7
irUj/+hDM6Q9bmxOyrzUNTeQ8p8V7oISIOrqazirX2zR86/UNW8S3qD4hlJqzrpB5kg7SNtKrHm8
TDcrXl9Iaz0GJKs3UFIA0SRcjIoxhmm3QegUGeErgQrvJcB5cEoO5rnCIQoRm8x1R8uQHmEvZcbO
W5Ku91EBmUXZODjolN4tC/Yd2cE6lohe2TYfY72Vltchg5gfYT/wb7k6Kk0Nb0Vlyk7998K4P7Q4
2LKEjndfPg0ACbk4Q3GPLCmY1Ui4jPVR+OePHJnz1Y8doOKnjFCL6JgHjokN763VVXpPhpQcZG7e
UnJE2Bafg4aUfO2fwSnAEE6pS4Np1a3jolampN/7R5ChMlHZl9T6LvfJ/oSM8VzKGkJI/QrAbgJR
R9bUt0hx+BGSWQm8ikGk0e/0xWANUSW/2IonOLvyLdcKat09VOvR3xzyFDkP4mu6xA7Hcl17QCcE
7J8EavmK4uTtIs7hgCn0vP11JamZ87z/aT+9T878YoEO/bN6L9musPfvM7mZ/6qWXaWE2msRDaDE
qMsi46aNOti38PHco9r0l38+KX8p5YqMVFakT+OYRBoDG/KU3HP3toeeX8hWAxCHD+ejbwLetv4K
NAb5M6MP+U715AXYLaAfSqR9qYAyUnu+fx3Smkj/5Yumg9ph7Qvu/hvOuZXd8aFUaZ1MUqGoJ4tA
BUAx/OhomiYx10N41RD+0idw0U0TZm8n/cdS0lVhq9DvACv8Oa6AADfx6H7m5WD/cGiqUn+Q40+j
LvOT3IQxJ43WFyrY50QqgTONKQhaHaGYImc8mdj7uo45viulIBoq8HDs6JjZ022sqghFUtcKaSN8
pJV62jTfU6gOutro4g6/3mQuEGUZIgWZibX2Bj1MjdCcx9oH7shNxDlU09fXi8zg67t3Hq0I98Lb
YFBXar2WTTWH0SflrscQKLeja16blh793haNJTx0vAZ94V+x1UrL5afe0VUi/7oN6i7fOe9PNyod
Ff4Yioh1Kf9rRPxgQAJGkXuK87u5eKhebb9ep7lh4/mCTgkEV6DUI8j2aSab/7T3kV7VqDMqv8FN
dMmBswhQfc5sU6nHZzBR4soaUQc/7MKUfRc+PZe9gE52Si3E0+spfYWjtfSr0X3MGFXZlEdc+zn8
ZEfisDTo0MAHR7CsRUD/tBIwqpXlOUnBn1CNaipnwVqrCfI6UXay/ZhPpAJWDv1r109qZUQvGzli
oz6hpet3ryjw4OmtF4quMn/AdwDBe5EAqARqPmF/UDT0/Hrk9uEzRAQp9QAunzBOxvYXll4f92fD
bvb05eWwJGxl/dArBwuP+uWm4diFrtc2UDDHNrV3ZW8ZOzSp9+EV587iME5xWzkJUchYoDXTDsDk
5F+FUL5usTO5OeFb/fA7JnL9BPZ+smsbIBH56cVl6U23/dXKaTXEMne1uPN3Io05INkuXZyuxb8z
BVKJT+9CWlukd/tNu95+pIyujg9ALniLfL53GZGI/NUprl4dt6x1BWRj+tOO+90BAuO0qSD0MHkC
0p0jFamcyq8aQMMC11OMehOgODIO33ql9KlJB6fBa3WectiYPNEYpXvG0mc6hPxKfUajDfG9E4Lc
aydzsWo/nKgN4oLt97SVFSj7IsWE83ObI+7xrZ/fjQlb2cUujN3E/lFhREKyFbck7BW1pG4/3WTq
YdDJNBcujEclSzBU2m1/oJi/p7+M/pIZJLX28ghqzZ2lG9yTzfzbdxzVlpeIsZrfS0NYZaipNZrX
M2LfmIrLvOZ8eXE/gEBwnaGR4qDP/kzNO2rgDMH6IssE0Fe/9gxejzIAyLxTc3If3o1vUZoQ8tp5
GoRnOMbPMGVEvvnCScti0oyC0HWFSz8vBdfeEipaCeGF96p4pd/2uAvCynF2VKretfDyxvA1VGVw
YqIx3wojeEC6lsjeBNVvxstmV58h5fUkw6UcCt9IE1jRNqguKXyZgcjhJS00+CPRe2Hi2uAnvyYL
BjCWhP4moyoOF76MsGq05rPgFeoth/n713CIYBLNskjljJqZbOb4PhDarKeD3iG9RO8iLnTBVUwn
K1da1hl5aioz0m3FA8wV6mHi5LyLTBpvQAxQuFyWDL1vFMhIt+C9TByLlShTQakhIN6uonsnFkEc
uzkVpavNcKyvJ8yrvrkX8eeZ/6Iu02Vs0Sy10Kebl3Ff/vtuf5KCwan6fdBCPqKV+cMDf6U4G7Q8
Clm/NB/Zexgx/TMjYZqYU+z8k2JWvRRYhOHgObXEb5LNu/Vcujaz6FtPAmYMqI5po+aEeJIHegSm
0/EnL+8ErLt7nLQYt1YC4E9MCIfHE0E4KGR1V5mRycpxeTXHkfylUgs03OQsjfhZ20gXHR/yWcF9
bVDpiV1GFzJPiOsSrZLIToiXkLqmL3jbDyJv2xXrso4vrJpvM1WPyxEzxT1Btg7cxslL1u63p0RA
usb5MynY4e2I1xYI2yGNL4K6ucQn4KqNuA4lhTbj7ZsAfprNGAhk7oq43LNL04ZHdU0S25M5lOLx
u0zUH9Pepl95CWeh4GJDMaXQaK5xPzJOUycpEhE6ZVvyadvVzeSBbANpeuJRjp6eanURbF4S2wzM
hv88wiLmkfbW4oHyBX07bwmlN5qncsdC2PbVU7OM9xaim6CGqoFPx5nA9qq/Z6+C0x/4ueDTYb2C
Y1Tqq9dYEEnczwXQa02ombQtLbt9BxGeKL1AjDqboR8vh+j5/2nV891bKaJ/oW/D1Ykgy8BsptjR
UOK5kQoM0RXC6JMCi6/Z9faQAJYDcwhVDlRCFdcS8Id+PZT4puXWc0APjuAOQf4G7hO/F1eG+4aA
OCH04uf+C2y9Qv84rqYf8HkC8gmxjk0LmSI4Y14X4PIy0kBjfebzQO0O2mPeQw2Kud2O2Bj0NADv
WWKRVI2z90UGNowzBztSx8uW0NSIVlPiQW9Ikb3t3qT8n/ynx6VlKzKRvx+MvSZxfy/9yaECR+Y9
jNtWCGgC48BevvIZX9lP0tyfEHVBPHEI2TLtb4K5nP1v4vm8e1Si0T07lcLJzKYcHVl84xIpwkPD
l16JIlWwUiPg6Nkey1TPdTmV8aTX3aPPk685XEO8LHrERbsABsIx1zbubzl9FNhZUUkNO8FxM9ir
0teZeT8J4KzMA3gIWqZ/CVrsAErUySzKjOIHBWRfUmH8jFmqxt5fYaa4emXxcF4F+sIPNk/fmgsN
iCE+8ZqI01TC+WYJ459T1VeQP3/5wpXP9g759Qa2nSUNzndDdL8UJj5Sm6iQpxL/bbwkeWs1wtnF
cTodRDY3WEaZ3wPdED7nLImxa2qwaXyM0v/yds7Zvz9o1n/kdqchYLvorn5xTD2x5AWTsj+Hir5L
8A7jaU2UOKBrN0KRsMiO0ahB+R6ggz3rdCgSi1ODBRS47En8VsPcg89lYtvjSS78e40gzH10NHkj
xjX2CrrYrhhPefvt23P/LD7xwjoztpSsaNCk08Pl4qdw8ZxsicDXnzjuJ7l0DfP/5tsSvP3TFB9B
9sPaNfKA5FpzvsjuGAxXOCZQ6EAcDWZ4Qidw9qBfLUhe+hQFfuufYFY/o4d7E5tuJVhvV5mtxJwC
LM9jmXZ/0JMctSxhYEwhUEgY3zcrunN+G1gkZiywZ2Q9B2UnCEKm/km4KI4JEl7QNRuI+rOW1Pxj
KG8P8f9Th3QsdhVJWRung0ZXFdfxxRqCiBhnfGJ4ybrLxiBJkT3oK1mHGj8tjjLHZgILpI3QPkcc
oapQK8pUHYAz6NMIXS9CPWB0dO621vRdNQky1FThysNZCL7SF7M5PF90WaRdImX9ESBlXHZsQnW9
yxLlE9ZBX7YpizbnU+Fm75LSZuNO6EgoXTFcIHCncqZ077LHKKmDNRZBO+4VWl4/Qmj2JMJusLJT
6g3V6u9KCZTfW6wbl2yBkMF23mzEGFxcXoSFN1XD00N44uPVA/UAEYHvVyfylkdN4vtn/QWvOz/K
pIsAUhPtYvnwOfzbKia8DgCDVzMgUnLjKb3OiOVqtZVhv291jpVu/Ow390k3UaRQj7i8N7M2pBD6
2niMaBtBPIVfAfkepIok6icZNqpF7Wx4ISXxBC38jVFDAwOFgtqeQ4apCtePfmIJRglik/8pjxh6
tf599Jkee8athaAcFZiPax5+B6TaVPDIhlsiRo1HsKrGkNfdsQicC8zv4fyuKAa+44iEc2nXvyla
TM6OKyaRYy+X2q2yWf5AeIDG3fQsPsPEXbZFX1RN8iYbYqbmjs+6Vk3qvD/h83+OErUATF8q5gtw
YSQkUnee6Pktg10SLcgZpg4iVqu/JV8ddLAJfouX5x4v011OcPw/7ZhIVKxyDrJoAD3mXmQuuRDX
xCesCD9BbhftmzX5MvrbSPltoK7uaXPXIY1Z98/WhDhLhaWaOB0SzBvWN10+gOOHFSWhf2RvS8vl
wTPaWxcVDkT8V/dbG/BxcQsLtw+en00aOZI2YBKvMOBijKtJRqCtFLc2f0wkz93Klyjzw78IFicv
U+dz73e/HpoUYJOgQSxDyvozp3rz/i3dti7dEaLL1/HBs9UqEor2CYzrodQ6ueveQ1jOLDCixoJF
jg4+sMk8uqm9gqI/2gPn4MMVE0f2t90KIKVn3BF7R0Qh6e8Me2sO1n6M8ezBu/v+3mXxkPw0hpJo
rGg/O8VnjVDkcQ+ia4YKpWegkq5SnKW1kiomTQEpDbMdIb6hUUr1YcaxEGkig7FMvwTKyfzWQ10g
lMZ6VNNINJhVykfi/3H+z6mFFJoDhIbuPZcFHCBNsrX1o6VqwCkCqyBI1nbFFC69IXr6Yr6K5iS2
OIKtIwLekbnfCWDLSh8ZvP5XoGvvUY5i3jaaT6hNFeRIB/jPtFHbNBDoXZ4oCCnU0BE/5qTft/Sd
LsTQ1hipO50CLf27zCaiQeUyp7/XifEbed+QkbN5+oee3KK/S51P4tTOpDqtrxjZs2iAJIcdJF/B
3bLnZM+/F/OjWbQEMhTwPOi6WPPawUL8XtPASKbR5eIpQQG/niqa2Wvv+m6NXHhNHJTrSxFjuL7k
R2lzXjYOxyP1GeJlno3NttnVlBKZroSAZEVtXQbmuSy4HxLz8vn0rKl+QcJZNvIeQWQx/KQhlxGb
MSC3qOHMhXq2HTBCwCXvf0cQWMVu8bxpMVNjY9PlNOkbuCCngRcYWRWMDwbQSlv5y6W2kmrgM/Me
jBMpDPGHlgU11dOFBRVesRGNo5LVeHbwnj503/Tgf2DNnHBZvC96ZX4U0rrPYCC9D7rSTH9f+Jgu
+EsrB31gjJ56FHuWTNOpENBMAT2yYBDNKG+ArQLI7f4ZNiKkDsO1GKLFO4LfXh/Vs+UEOKZF2PCQ
agEaSuQlp8Z2+99KFh0fAjYNlNfv/LxFb/U6R6Lru53RM72IDhbLcsPrGS2J9qP1ZCZbWgs5/XS2
D5GbOCJERhY3XWelERFQwOhE18aVbsBBoeb+IpUFYdElMoMWv0X0wp8tbqYiJI9NHT7J8uN6DM2v
8n6/H7+5aSRYXqJpyCz8Ztr9fR4vqBK2GuvUbGg9bvQje8TpBqp2RtUktsqOcbUfB9XPQykpzY62
SL0FPdPctoUjUepCzlojteDYHI9hNVHKdEu6D+6792GW2eTgkfbsg9CrOSu2O55H7rPc63SP9s0+
ShEpi+3/nKISW6ZigPFBEaeHv6XR0NeYK6SDfCtVYUOsXXzikjVn2HU2f2iQaj0PgiHAEgHgMwP8
GpHrdr5RDO18A+zHKYGwSJuUinsov1Dm6Q42gksw65kPej0YQA/MD0x24s5Kai/deWNFy9Eq0WaU
Ry3EN0AMMlhMa5lfO+6uZRziaqjBy/c5cXU+IkjD6VIeV50aPkiWFPlyyKy/CQelZVibaT45RyxA
yDGe+QEHs4XNbCKHakTydOjHLjN2ocgWkyycFV/Haa9MVi4ZEKxLTpNafZM1z2eHJRizrsb+XZ0R
Qw1ff/2Jk5eAmwjvpEArsdK6JlMnNaJlGqUt1YLJrRO6MHbMDvrAyHP0O5DM2YioiYk8m0RgT+lj
cDdkgDSfHnfJHDHbsEdp0W7IJ3tjAvG03kbx2i3fBNUqhkw3WiuZ3NZQ4I2T7pfm7bkhr5/Btf8V
0HFYDj6O/+mZEAohkc47+PIMqq0lu80lbydyTs34ytfZXvvCWJMaKWNPLPgp+QvW11r0HZvLBubt
vfNZdR/4lxOen2t0Ms045FwyWQB/PzrekBEWUHdUaaerGYC3kulafTuDNW4a8iR3FhbTASYbEPgW
WMw/K+Akq9IyqAxexWVnDj6NcJDeURaSgXvJOLMAsrr9XXp/1vlOdaJ3DyMwF1JFNI7hKm1heQel
DD3HuZehhfw9uuBR19V2pWXgvOpT6G5DulNdhjqp1UeHvGrlf8yiceWVNAonu2F68G7sHJy8gUQD
vv/ykUYk5NLegFm+1AaJDR1Uu+GV1LBtJ8mMbk8KQnh2YgfxI4zpy/nKjDwEO9w9mkulEVkhU5j0
Ew0pCfhue5WSPvATedfbOzZUbT04lzO8Fyr2UL9mPZ7ESInmZji38kdwd5hP9fm+JXvoVLtbb0mZ
jookbKSsYLmUY/l/cmQuNEighTJrVxMWkicZejbA/KVSZAlA0m9NeoBCEFMoj42A68kbpWv6mElS
xzJr+oD6Fqw3rfP/dSVlhe34jpXYXPCquD2/UtIQHr+k5JJdSXZkQzq+LsxPyp8W33TQc0K8PWrw
UuXJeqexQx2ATyKMPXEzhXcaKhgFkF0sEBqird+4PFpPGAc5B0r1vrJ++d4dcXymnx/9izMoXKG3
Cz2W/wUijygF9/IhrNB9IoVTPQF857mWAa3ReoAU62E21Y1sTn3knHBg5cXIO2tnU1t4HfoWgApV
MJWRv0UNMQVKRPdha66Vr85CIfPeswsQZ6YPcBZL/USClrJeMNi8tQAqC1fjotFmHBXUgIayHI+e
yPVhj/wr4hpREBSg55Dc4AvAZVvpM2b5Ay4qpgwo2avBT2ZpabOFeVgCFPq5XcvLN83y9dQLzpEf
S1q4LdcuCl00VH8FZIcouydiMq4ryCCXgJLiMfrpre1bmrEIB2TFM/XUFiQIDekFj2crXGVw/bO0
H1c1Id2rOQ6G0CKz95KMgD3A/I49YEhjRzwGjLbfY+hInuqAQIjHgxfgBoLimEuY7Qi2jnK+Yu4b
R2pRpb73hKK/avmDKYf2Gwsih+c9It/l0ne+4hw2PhDSvlA+A9Ko4eJlgjDoWdmfxiA4pGVJhH4F
rHd9+ScPWV1YAupe+iOMWCIOood78VPdGXqlqCyufr9lTSUyqlUUcJmsTaFrzoflemk8YbA1uWok
hfL6NSF5++lracN8bh6spTM+3IjQUy+KqhZY/QlfJNjJ5PFK06zSNDg5gGffSfg1muzBznY2i7pV
9Q3xdmHaVZIMUVRz+JFiWNlfzZx56RZ2WS1mD9dU8Sb0keVnWLNUXLFt0MgZqdp2ML8hiOyAMsF2
HOuGcAx5LvizEAd5jhwVPP2DYdU0l33Rn1Yszfd0Tgy3DY3djPYM7I0N8ZGcZpHmdMXrhx0vAvN5
//FKiv4NA5gPFiaAbCgwjpKhnIbLRkUmLReQcxmKZ+k/KU1dzcn/K8jCKw7by4LFgyVTb+1FNJOt
1NW1dcvwLbSFyCK0EHelG//eHx3YktTLdKjkUBYbe71BvKslpn4dZ5DxtWyeICkprVOdy3p3t3ve
Q56JvGy4WibpC9nUcP4ZA04PbU2wtX49VTFisdcHsNSwPe6bYYu75BIdfwbpxcDoUC70SN0SdIVu
BiswnCrN4d7MlF+loAyLliBbkWKJXiYX8MVNFAeebaBvM4IhCI2t431IRS9rPG+AyK7yLJ+PmtNz
1wC5nUtlTNG4XhLera+3O4yM5IuB01q5TC0VmwavhpKpedkAu4ayHlsbblcJGpx6+aBHfr1NPUel
2lc4W7MNCqeW/SbraQ+w/xl1VQzhE5Iz6+yb3gh36dHpeQLZBbh3PMiQrVUxgKkr38WYK67B+h+/
ZEJG8dPOcZObWMmDO0sP+0yybpZMkUGy9hNWbAppIgULZQFD22ljrLhMA/NXK/hosh8Vb/K1Zfyo
C7fbMYgzpBs6PP7UA93EzxlybGwhtN/SfqSWkU7SlS9G5Fg5LJLyv0AI8rfe1+uJEDHLnt2tZc3r
WEFuWOK1RsSPq56h7l8siY/HpE+7zCZMYtjU1WLQ9i3U/ewDCjBKO+uMwi15oCDYbmJbRok2ZidC
SAG/jG9sOOLTHa17wZyHNm8tcVkLX55xtg92R1bVV/hbigI30gJm2I8pUk96I8gtKL/4GRVeKv0p
Gjg8ppAniLG3RWEgll631aqYrjNuDlsJhdWzJgeksAglbzoZo3lP9BfKzI+NhTrWyeQ9sGqDy0y4
j09RmoAURt6ZEINT+J171UY1s0XUH4NaoDbsnHgr32k7gKRTd97BRprs6zfEWkTjoZrmhnTpQJMZ
VBBVbK/S5yngbgIVqxZSfh6X7KZd+N3sAV0HRDATECW3aH2y2BV3/8Ux6fUUrqkhqzz+R4Qlv+ss
hc0t8fbZcD0Qe8RZpPpat2k7S+Ww959aMNM9OzMqvcJ4hrQKGsIpc59oAcr3XIh+mnWJFT6k4cGR
w5ta8wRQFbpixH0URtINRgVtRSaQgIh7u3bZxj7VDkJE/qlGI8G/Vm6WfUmWkkyHKymF5bOniNX/
gDAtn27uItlcSw2ozzrj1iCOp3DWxCSU17Y+VVFMLoYHQd8SSXUFGdFj7DWw5VtGpjg31M2BiXuV
5+vZ5lihPaCWFR0P8ZMmEtxz0e0gBgzftd5r7i9YkPAHifXLprChoAPg1NUPMeBfca7KQwBNPB8d
mjZ3XoaKoRT1zXQuQk+ofuZ5CGVgXAIm4beVllmhLwlO5n7iYs5N/09WleYpbLXnTxXNH5DYjl5P
fSJqX8A3+mpeasjBnAPRxj+RLis42Vp2NU6ehAaCV59fTB9nRJV6gKlgBZu6Fmtu/kIxfpu8k1Dg
Sg528htDn/KeopAuDRDQbY6hfqb/I0eZgzyWxZskWaxpiBu6UxwTWGTTp52v/n7isRjLspb1t/wN
qDx0FWsqtnOS78DsKMDQ10zK/mbxSpeTH6Ugm7Zr6riMD9L1Pbl9UapNpG4vwqHnvD/sBO0+Ar6o
fJFVHpmUqa3yURAjfPCV5S0eqwHXWRkZciXzIyPGHQkfqIXQGtBRMMK7zg4FRZm1Iwz9fP/hfJN8
3fwTz7HS88ff3NfipPwCPIyg3tMgt9J9cjuojLdK6zkm1+8AbXRC8icHFopvMfh53sgm0MBRX9r0
z7TaG2reoK58lz86pFA3jibCC2bI8otTofl1/78pN4FMyThfL1D1LFY1WR71VjnFXJsOTTAM4/oL
9pYoKrLR5ZNO3igw/8DchPkecUY2urZi9jyDITSCWhR4Q2noDXfRilWLmbundGxvkJh0QOnG8Tv9
U95sCA3PYCMH005wxj1b8k961qiT6btnkX8+yZaHLlqX51Mji5FoX8RjnRbeDx4ClkUmD7hReYvj
E8jFG6Tiej4/hDj5dR5QWkSC4SR2y/dQm0fkbYiE+hsfSwmEoajrdpCyt1xeF7HOrFK/1TXlBDip
fah8/YackO+GpNvZKgrBIgwLojbhpseU4cQDywOGLfcTKYbURessEBYzakirIIqiF50JvAY5G60v
ByAtJmVKl7rXmkMFtPnr+TNyxy3AmpkEwqZc2mIZjg+xThmoQbwXWlImyYIBz+m+njp17FH/YqVb
3dO1P22Cp0Gb0hLXKhK558KvZ9FPOVqL/7ERKDIQtaG4uN7IVquwRbtHkFTgU6rD/cgBCoUXTuvI
es5LPyujuHpgvVV+yGVsGblwwAk9S88HyftPTES6M5wWltSF4v93PRgzx944JzPyxcOTHX+d/Zdr
ArQIDZdTWdTDqoAo2EEWS1Bp5DKdiEVJciZGBfSf9RJVOVswfCzR33QXpfWAmBGOAEaUS1RuzqbQ
Lx03vLoRQPXwSInGNu3g1pGyz9zCjlzX9d36zpMeGehSAwOmTMPulOpiDvDUltcKQwvLwdVJAf7q
RKIzxZ/eJlFSn+qMemtOJbujpUaWGzULEKqY87xNMUw7ZsV6jY/3nO/eMlA4EkxlQSkgA6XODeRF
4ETwIQK+LhPbLts8QV4zC7s3HR73rg4lDiOJkGNfpTbyxQPBepF4dPimrjaCYiu+4hUjQ8NCjDz3
82ZHQwkqsUNFSSV9xuCVKuaZOFQADXf6h4dknbX0SbLtgI4EgxXbvaeqRH9IURESMZRjDFJo7g3h
uSajHwK7by+sRCudOTZ9TwyRhHjW01nEveSJt84+sL3c66zoQAv0cIZ+mASHAwcy/ln16VRUlos1
7I+tUcveNEqjvsmKGmc24g3Sep3uwf+SlXkLkSdaT5+qMERp9hxrrDH6oBfS/yavla+zE+HboeEg
zMqR68LbIIm0So8lNAMK587ybNKy/7eF3/Wrtrz1ZuOvDR3oelntWo8lehQ1pEvRGEZXGleW+ZdJ
avNu+ze3uiH4GV6GL3bk1qhqFghnZiKvNIVPUL1Jemqpn0rExTxHxDO27avj88J9t4gygdWEXqWf
hKoOcFNS0GAfreBHWSagjPlGQRUdYSpHzQFetFQ7wRnRqrKxfaOYG1UC8K7wxHguh3a1Nfw3JPZj
wBXohvQswH3YaSAsw6nBAus3BK0Gp7l7Yqwlr4uFsd1dXVwoMA0X2kB7RlEz7p2d71dtjknOr4Ms
nMPydQOipwSP3tSN2y/WZS34XSAQqaQkPpoqrq+ciqqhs6T4+dDFQQAW0Enag26awTfvykRSXH4M
mIAtc3+AgY8ix6DBtK+wd274To+HCp+MuKPwBtGgEYz2Dn8w7+M8fnv+Vq178bIESp1M3aueGcIk
C0CfvhlI6Aa57/HYVyncNqpt0ifgvD+o3MIPu3XSjjjfm/UstoaxeUP6jopMg92vjGlW+9C6cdG7
R9Uq3EwOJo+qncxKljjsMxzDv0Zm4eTq2nQ5aXMZtYZDanByc2VxVdLl07heLgjD8SJX5Bz9GEJp
ekbDHVmizC2a6lgBhDMVw/uBwZHrqxoxrexEUNqbvJ1zuo79tzoZ9IFBe1ZiBTceB48JNYhfoB9R
nXx9/AwKqlh73RS1K+ff8KDxvyP4gGjfhQv3yRS3PisD125W/p9P+14ZxC9k82q+dR01mflbJb2Y
CHTt2cFFPYNLVDb1Aax/ePPJEgXowO8XnxerWrgGIOhoChRX/hXJCWY+B9i86j438o0bSqlYNGpL
5Svm5QARfEK36Takdy54XU/eAGN7Aww1OpMva2iKLiHO9odtJ/Cl9W+9pWyjqC4i7+Fsa4VoASPi
ekbW4WJq68053n+7jP48OeewCkvvl6HwxUzvxfjAZ3l0P9ccvKjKlmr7XtAogkA3l7JvI1taUrqa
rC+I9uIALsmxbpUC9+NCAEq37rI5OdCcCMnlg1M5Nt6nh43NfYs3LlH0GJKvmaSL49YWtoYOKxfQ
SQln8WqczoCInTON4kDl75nH0VUdbSyNK++AkbrNgs57XEc3vbBa//LHVRFylBI4fuZc7i0wpK9g
gkNxQU6Zgf7evmjnjoWE8O1Gz3rxK526MjnAoqY85mnnxi8VgPC4uzqZxSY3cXCLRE7zwNsjQWEj
EsxJslcYG0U6CyHRCFm6952n6HkhomNSaysuBnzPeDS0CeF/1Yj2AwE98oto89Bk0jKE4NkFJBVX
nvsDKZOJ48d9u4sNw8RG9UVws84sw7MbZMmXbYloULXKIY755AseTpDTkk6sw17EDWJgAiV13wBA
z8KJniksE29fkkUrbgZqrT1J7kOQmB4MLRwDcCqMjtcnBIFKz1Ka7Ac0a0YUAJ8knVA+Fwq4roX2
ErQRZkaQvihZEMxM+5rlTEA77lop1v+FIlH9GWw/GfBxzKRMWa8mHtW/dpAo1ZYlEV1BF4R++SHY
cU9jzaJabSl7bwVhVbDZHEihkSxtsm4xImZ/r3WsCLEWcQ64t49AX/zr9woX3NGDsPbrL4lTrsMD
uA4nC9c+AUBB3zB/G0xl2zDfhilhKbRuCcZpMyiypzf8X/YFsTVTQemcHJEzekIhF5PJDAi4Qipy
7IwpQokyMfeKOmTqwfPnURGbt5Q0ulUJPucSnY1M2h155lH+4vRWNJe1nv2xRUwmpnheKXYGcV/H
gDNO0i2kM4FaQKpIu/m2pjW67CMRFPBKEwegzNDVJoVeaeAzDwjQJGl0gk3X8B0gJoM1BCnWH+yW
AKPRPcDGcqj2S9umQysetAXArA10fOsIdw6FyZtEt3ug466EQgjS67y/+DC2rYsiGpLYWHOz43ON
dkXl8sQifPPR2z++pXPAtUx85GQFw7revf3pTLErWhzVO7AXRpyUPKWxOqEKcEN8I60B/wTqiXd7
d12C8Xn/94qhZWiWSOHV2yWYq8rRlV7UDAn5HxOiZKQYFJCpgZIEeeQ7IRdNeEGuEh8Brff6KY0Z
buPi+NCki85P74odbdXL+H5VuKUiaJUAXuhne/S98Ho/TAEHPcrw5tbuWjpOWkTGgkUvl9+1CzQ3
O8h0od6NNtBIu0VmiKLtJHnLhauiOaAE4pDEveHSXQ0Pamby3fyO+OPtFkiq+HER/fvH0IlPNhoQ
1tqvPoZrjTpHRqghlNt3Pwp/MH9/T55q62DVA7GwpQR1SbqdJjcpaUxk5GLgQdPsp118aklqm+yG
Pbm5LA2TvtF1oLMPcwWYbecmZRSB9jIqUot5Fw1PFIeKrvh1xppNxEYZGPWtAWlLrk5rYo2DkJId
Jt98VV1z+5MbQsXlvr5U0Lj1/RDDR67wywJxFDl2ukn0DCAGu16ku8YN1RnSxoJBJBFGupM4oOkZ
xwKTZjsPGM95fviqroBd9pEYwDkFDQ1hTFEMQEY3M5WI9AwU302YyIrYYtSiFiYHNZZ5+bxfBHKY
ZWaImmcUg+Q9wyvW8gvqKHSvis0+Mj3wOqKKTeVknRUey3tnlk8mIdJEQMexb8ZH5U6SVvfZW0+1
NP9B8xhHJVsfsG5WtN0wRORQFj2Hb+N6zOS2MaUhPmowEipCTp8pppSKqLMMV0mdc3AGfScIQ6ZA
mJZrWo6WhaaLTwRTGxpiztEqoDNu2SO7ZbJLdiVMegq8fY82nqFYXI+CI6QKqbubglCwQ9qf1Ofc
7NJ2CfRnDMgMfT2yqaZfI75SarTLNrQ6PRU+avaGMtU4ztQJ9KenPma5sTTsp/qEWeToPvjlksI/
jKRpR3/wgLM8KAg2XOUgkuR7Wn8EKqZWgBTyjpne0rQbulZxVa4zUx+EkcXUn+EfgRd5vwdsY7tH
RXqQi9IU2oc8JabA3pYRqFX9qf0xKn0cJei/SzGCYRrI7gWf+aBP3zKILVWvywEQcXJFVUS34UuQ
gJmApOaVUlrtbRcHyq67riLmOzVPDRurDf6ySkmltDLpd/UPKiZph1PuAUQt2mq2FcN3eq25aEZz
J9ayTVFNFSEQkAtIjsg5b2hoqWamHzyoDW8xVf8UBBLVsQd8XDVWNpoLsmxqKNARFrQqkxPSZLVt
YXFHrUJzNcOe0zuNkSaw1wl1+t8B4fbxuRekOfyqliaqEDLa2wwxcFHA/eNsl+v4ned0tLS0M6aG
REqX+vdJr9rXhsiH1lZ4is5nW7ZlUl7XASj3kpSXdE6Zza/hXpYa2HVIDK3hcGJ3yORadmukSE/x
Cc2ke6EvkoWvBpdhNFxthxJyGqMg6NIDaTJWbZTpRrOWhE8vbpMqTVecdxCM3N8gFugjagjjGIsk
8q4CeADU82MppjTKLyvREOPVlZnSR+wJRJnZGIke6gm0w3jvnIbfLR4FiwKOjCJRRe+0e6Kb12ng
OCxtTpIcmgrR9lQFdiDUy5QbRuCMOtZfaShMi3CnI3HjNCO0YUdnmkPxsaynP5aMX3U0VgVwj1Lw
lLOo4x9I6EQuWA5r4evS1cb7afhEic19Y0+rZtVZ226RIa1di4nMreNwxwHbD/C2Py3V+Y/LV/OB
78XiOyekMue3TxvkzzEqCpUUqtZDIAgEDaLen46Q8H3R/WLsAc+rz1nthB40DNDn3Sdk60e7L8Yt
vZsN7Q+yUye8MGZASLCjDIV4GNwbxY8l94xKXDqb0kqhuCRDUzPW3m8751HbZ0Z2QimrrDxSFs1V
ZDSPt8PCKw0h2oIkFviXkgLKcvP0OfIei9w0WGDB3qL6uEwBYoeyF4AeZtMy0rDb+4QFzwlBFvvD
G8OzSs5mNdYpqHcV7n2nTyh7KxR2Xu5taxvScJicVomPOJ/JyK/jmzcQpAT6UVrbgnLltHY562sL
D9yD8zYqPidYLNVcUh9K6FcsswBXyDQgnbbx4qeKfpPgwNt3hzEbeprJtH5LdpqvYWm0DsbA11wz
iwU6T0G05LXsayk4oHVciMeTsRS3TBbKU4wO3rwTKcNiqr9iiLMia1cr2Rh93Ic2WTzed9UMx8lz
xymCeijYvVHRochC59QsKDK0+5Iq/Apm90zLFbuuoL+MN3hlaUqNIM2s0RqjPoLV0zyQlMy16qhc
awClGLxkxrxxWyaVA8ErnPrZKe+NCcROxj9A4LNDPBPclTgdbFO1OyhcdpcL8x7mf4r0RF3VXRMq
11J9LjluYUykhLeg6uFmZpar6QtD7bTrtXxtZx5O0jVSHqvzD5JrMlo8zwxKsXGGbb8AXQSJJrT4
pqyT429GcaR09ru/scWbGht3eeZnTQngxDQVw/XpGmCWihChUR2F08KWhMv7YFMn96mefIwncgA+
VdMm6jpsHh42+fOkivWo+KwP8Au1JatAr0zEJtNt/wsSgm8hpPm7cspgIne9pa99X4K+yBy6TRTo
TbiDDZqiXJkKqiuCJOKQnmG85//mkHZquWLPe8Y2q4Q8qavAzhZepHcEapeFCFvMKSZBx6h831FH
yET8WMvL4QMi/WUmPuZzVYD9k4RZ+qf743ULxhJFOoCFpjTqpPk1MJPh9ZdRgT64YHv8I9EV2L4G
BwA07G9OoBqiyQRM2hKHhRKuJwvyUst5fvUbe+bpPGlP3tEd5Yw0a7M4F0L2hMTNNDV/8LV8Ra5p
ThawqOQxIXHpGne9bsEm0wluJLjLx6okTFr2AfsVwF9EGnSOzSUrR/Ya3lOWuVcYI44L/GsOQ+it
F2T1GA/yMsw/qBETvsv8IDvfOw2VzDxxEwBL6ZSubW2VIYe4uVrB+fql6HSoWFR6IgLGtkR65YxQ
DlBv+NupJz5gBZr6mp0b/XUDJF34Xu2BmNJfrhv/J/1Y00JsiTx6K5Ar5UudUijzQskLaYIdj0v/
xC4f8O7jkIswTRNwtq62fqkUy/l3tYyxBP7BVnOzATmaQa0sGr8xBVFFF0TC8+wGlzA4wuaiSIuy
6EB1oltPj6qj/z9cMBoZvTrTuHHUsl64TVbMReC4Uy6wtMA01EP2+Wi+QAyPKNTULN/vBlIXfs//
jPHZhpVn4br1+7sC8QM0MDxriEjCO6mfxupHWnVcIDjWnf9ZfSQIfhuCLQ7VQ5a1pcLKxbs1/qgU
zA/+fBNzARSRMfHoQiRyrhmoIejyDEBpWzxBokVdL0kxZOvgTW97M0VdvqsOxv0gG0S9UwLbSSBZ
9i8pymf2us5Sec+GklBQH+fDi2hTgJNxsE9yM4QoJ853vMpYJB41EwrNq7Wgr5dZUPDGM+6d6ysc
ke/1MJcB9szbnOR4Q88gRvCUkxt6YV91S55l02zPCPpzIVKktyBuTDrnOqUuBzUGI0rlMDtwpgwm
OCBwWj8OMYku5iUAI4ixyIDHiFbW2Knr9HFgK3t0iWfkqGfzWkfSovyRx8WshM2gCeLpe3mlwXFw
wBAdwM73utsHZlT35bq5QGFlIhbOMhvdRb4NmDkNm0v1eVRNTZso+657WL3YvGPXMznJUi9bwhmo
j+IeBpXmdm2hTbx2wUme0LI6M4s3jEmoWZLzsj+WqwvdzemmQ3PzbKGex4V3owgbG+KpwDKwrZwf
QQmlpKmOdFuJt+JIj1Pe4wKTV5kpcGsTdMVRih/60ylAqcUzqEGv4UkgBssAEP2mTQcLCh0MzS6/
QPmNWIfPBEZBwXz+gmAwDeGCrWf3r8IzS1/VpeKyseCxqXtHxpHBA5LLaxdMeIJQ0KmS8mjO4ixo
R7Qc+AA33vGy/+9fU7WVaw8KmD7fsQ2HxgJCAlv4ggVcmwVdknQbYdwu7Drc7+NdbtU2L+ZhJ+Cn
vl//g3Nfdoz38fHD2XpLE0jsf6hCvvvERyJGWj01ftYTNd6cya3AvmFYxKcIBgnNk04L9w7Qe+5Q
61wPej/7CEx4WWoRRwl96u+pBppojK5LAAF91dMFKqm4NATQPxoy9qrHABaD6XMPQwXbOHmvO9lK
5dJJU0fRNq+p5RtdKZvM3fF96A4HDCd0XvpIAqLwAg+dOBIGpHDEVT34U+SrdApvo9ClODAHdk/f
EtcQyTrMTCpMZM9NqknKmS/2mbSsFLSyNI+VAulSgQsFHbjF3vJ9umqx0tkkZzyTroIs0wtyxj/8
0VYm6xkHVjGO5EDJsClPiIfHaWVqMrDQHHhXnIaLbcQJrWkClQoF9CH7iTQ143dtYzy2mR0mGo0P
jUijjM3DeVjEdZmGgMq0YVjPbGSxgRo7sX4a8IVGQZ/joFNiM2twnOHcSgxutPDSqw76LVlIvU4B
ETA3kz0iCk99qvBrKo0W5CQTKceS/NVUxf4V94UYOc1WRZqhcQw99j/anDOGa4yaWghu86Eqlfa4
/IaEhdgIULrPlvTUB5x7Oxpheo+f2pWI/32NLkmkzYfKNRCSsGOHV3CTUHkGkayqUqBjJKyhTsR6
xJ/XkGaZ9kw6divlBjxHuvHGp00CZo5E/oJTaDcTt/gfoip9d/AMn0RBTuO6ASPgjhqI34mnQA8D
TrrmlpLRtoe3YKuMOdWz+jWdH5eM9MeCLKtjZ6bPV12ykDiTTf5kbd6TCFFKYIkynRPm4hmA/Tr/
uZsjhuI2PAm4g/8192KrBswzZJGucSFiN5hwbxnm6XTSwMZB6srmsdeLXJpUWjiTXGs1HTs84KUr
vQQcfxiMjkuRtDHh89Cm0fyr9pXVmpvvC5iZt2qGQgFOhsK+27Wtnc8hGtTBlCygpMvCdsktZT9L
2osqzfesY8tyLTkd/c8ml+36JcnxYhr9Cum5o2vpzzp8LDx9vDHZMo3zwnKSPX0MRsPA8gjK9F9r
n/1kxhGO9uvNiMH2TES/txH8WAqTR71lV7M6DMrno0xX178F+/XE/7M5oLtGCJ2zWbNw42JLNE4W
VUnHdQDtN+jUkIvTh7pf+xmMMUmFo65X+PyXxAB22959NziXCwJsfaisyL+tK8jGVDOVBnS4JyR9
Ewp5WU33d/B9Ig3JFTsKMXdMwOjGI+2zDizzyGVUXsw8/Yd4tzWPtzErzjzZTR5c1As0MoC4m88b
/WOqMBWIHxbTSYmFjnR4NFNajb1G8KhR4tDDC2/5SGNa3gQMc78FRvXONuMTyOcBNF3WlRnGJnkp
HkBdbZKghcg9h4hK/IW3ROvGyiandD10mpYI5WDZQke2G5m55kmOKUxFJvNLmXpvrND4dT7gSQBZ
garzZSRb36WmHGdhJncsxfXKtNpEquWnaB0gUDDccOz/cMmCMFNySr7K/IaXzIY1y5TMc482ZVB9
KJcgh6jfoU2yE2bX3KIkOHO8OP+fe3d79YhV0m+2QJmhwVKGPplth/k9cWTEOjOuHY9E5IAHG91e
0TTxZHWhDoPv91+L9cDPV7qTa2lLGRXA//xKViyQn8SmkUSqbZ+N5+k2GLD+hPAlrI2i4MGbf9V+
K9QHKd4MNGrMwp23DZmZORGbWNYl4u2vPMgA9VaEepGqIIjfwLrTe49zV4BSbpAFzLw6U7TqWFNk
M3dc5KFLYVsGJKUyH6j3u7rXuY6qOjVgF2iuYi8lsrynAm/8M+povIRBC/P4ElBSaSLKh3m5f/XR
Ii6qGx7+5adZYwjBc63AuCij9nUJr8q9PWZcCt838xpD93rIrd2veD6tJyGvEsrkQH4Uy6Lq+bDW
QGc9h0W0r74KMV6eH84ZtY71D15vUyALKXzpeshRMPnkuJwOvj2vdK6p0ZyRZYEHZYED3m09X69u
fEqE4mOVsa7xQExdnfkHyGeGfd2ioyg7fPuJ+jmYTnJEubVcqW6tf+1OqLdCg99ryToA8uj30DlA
d8xA4TODmW0EP7fctVfCjDBwJeqlXtY598RcDa6abIKDymBtNXBROfV18XmRa8ydyR3bcwmtEBiM
KnAOQurDUNGtxRrdgL9JNQZgbth8wj+Xb3VUTtumfD1jLof9IjJNzBXeFb9cFyee6qdZNZ88ZB3u
VLmr+2JxVLFG0kSUKt+Z1ZX4k2frKaON5nKC7T4ipqGglAhWPYDsEc8EgimimDPvmnFoMDAoH8Zj
9siLpZHCOAG+yeXQFHK9tgRH1RfNwo0ZcK4p1BXRuWmHxypbEyxrFaQnqujxNQu3Pv4XdN8TL1h8
oDBhKUbbVL+fcNkE+YRSwrv04s8y47ltxC6wAMdUyK8KXCO9SARd7CYx3CTPk/XTOC7hRymkzc2v
Mm9Q2QeZqlSJNOSdMU8R6S788Ub21K6TbVo3TztJiz/AtE++2XB18C4fEfNWdv5oBvJcm0jmVeIW
KP9lCrMEkHDnL6Y5n3tOxwhApP0aR5FChj/gFikaoEZ7NYXD0GL+IEBdJgqdx3lU92J6sgvOqGDJ
EVLxwN9gpnOA7fB+nTKHZ/esjd8ePb9nVa+wirDULuIBhL8HpoNOLGGM6EM2WoDsSVBLM1mHuONl
/8WG/P6CvHpNwcMV7kAfcx5rKahbRPUfWBCGic8sVllZoqZhSD0ZmHKbdceCSJkPu4uBf4J4Ldga
WfTebIDrAVbxJWO77/LIncSfxGOvDgpbHUx4P/WbGgnz90a7w1C90KQ1AzxjJ6xDdtQHgrQKXd6V
iHPIubtZLvP6815VpqBtXPQnjj2gdzxLvnP8N2MNzSomhQb/8pBNyQzvE0TDrikXWX0ftvZJE7TY
DuWI2WRbBqM/RqTXlSE0G7gfhewRUJO8wLdWMzZ8s1zpWLSdpoeq9f5PJunj+HxoGxpBqCa4WTeT
H89nE/ZmuBklQ+DOnigd+NdJcIiEH+9Ach3En+iHREmWkN2/Qty9vIkMl7KFnr7x3nL51I8dcAC2
1cxZJw+sa6CBhvc3CjXePa/RYnJtdPc4FBkDuXskIxn6LFINq5dr5kSXVqnjqxKzDV8Cwi9GdjLC
pVsus0ShTUv49JmeKh93sU7X/FWLFsujhmS0mtK28xL57Q3VPBBjqidkgLzgD3EbYs3Jz2lokz43
/fpgicM5bQT+NydqC+LYoaiSTP4FLFTXjSwlGWNJEeKwWZJphXqozwAfn6ESpdieTWkMdHQXKRKa
Pah6qdUL+5HXxsqcOpIA6EP1KKOEGTj1lp4K0VsZqWa+Lx6OyUSIdK6UYEAg5w0/hxbQ0tXYacVK
NS7KCM7DnzJ6HONCij4McKMiYmKM58+jhHMxgbdjbUiA2DuWgSmx3H2zd4iWb3O3KbeG049+ObFO
wY5bzeZlkcA504X2rD8YpxUGYS/kSF69jGI7cB1hAk6yF7j9fZt/Qo0J0MXLs2RMciTr1LGQ4nu7
M/gtiJ0GBEyn9OaCr4Uqb6tUxmJaOjeGSofGWsOHE0ApdEuyyhuYRHmu0+luGFeajWwUAIvE+G1C
1o8h/DTNPwiBzTHPOvxFHkDXEa9rkxYcGF0fta02f8e7trvVwfVIjbO/WfvSuNO3lF51KjUglUbF
Fl7U9ztk/DpLUYKhhtLFCAFLh5vicAseXkpH5OTz3I12AGrZey/r6j9TgVLH8VYstdkA54MSlGNs
Xqi8zVDkZ39XObfhpb+pDoXvB49q877A2fmYnBnbEsz02vksJePnfeBfrVnv2CGqczI4f2xCXWIV
YPQgEEZZvJNsyA1gfoigErEue8KH2CNUUzMYJ/Ids7GNSSZWiTPSC02KGTKCIz2/yWqQhXAyn6hO
fsUoei2m3Xu2QEYOzGwja4R4jUFbw2W4Gw9zfyiCDt38K8wj8pYO6pjGZoudtc+a0/OqM2GVpNyc
hf3rxH2LkDDdADxmbf3k2r17Jc2O4j5AaKd11vMFzeYQcksAdKUxtsMevE4s5RfyHB60bHFnCO0S
jwvSt5xTxLhuFCbriOvlpyf0zq0PzWscQjePbl8EpmWOoMFho+ukMliwPX9vWBjhbhOx5W4PlCv1
TYJb13Qzn7u5zZ9bxIlGW1aeN4BvDRphghX0NAO1CIJ86gbXlVG8jD7FU3rDBe0WSye7Pd/rK6g0
QvM4PIzqN3lhi8+UmpI+/N6bjHnvEDZpDeUyD+ZNctXHQE91bVn75UiNF6JxdEnDLtgOzgAsq1Nz
F0aCmfsXt6uFh5Eafw1w8YDojLVU0fgldG0Tp7qTyuyEPGDes0odijsm3Wpo+Om3L6V8Iq2z6i4l
hv/wTm2K9g8zTWygwfETQmGlp/Q//IuzRjmTr4e94cBUK5grKoEWmbn+kV1jJ9wejSUAdXvLE+TM
nbvPVgfDEijuIMWKd3LGG07PgRCTmuzm6aj9L2qV/XIawhNqC2GqgXKVmDP9OpIMfYUce5jCKwZB
LFzC1ZTVDwKrtUgcRggVaOdUe58/mxBfhixdlVjLe6zuCTYVq6Tpyo6njTAjaVcLaBO0RJRbmqi+
E7mwdvL84YFPDuvft7mxjsjmDBNVR5y01+CNIk3NrPe7zYiC84klSb0RsPR0xm98svGiWyDhVCEX
nQjstByy0ce0D5OZS44DV0llysTJZ66oGG1mj+SuJEe4h2AyhGl8+cdFzZbdT4c0r4t71XYRXz+Q
0vGLjcm+tfXsGEKX1z/Kyche5oV/S68/X/4P9BKZpkiQrgt4THYuM4rr4J95OrNgLb4pe4ujVmlm
bjFqtVIKMp1WJflxNioVN5yidUVT7lolb/Dv2SFHPBsHgKdv1GagrkXZ0Ima+clpksF6zFj/C/l8
NcIPdHw8LWwuQuvphbWiHQWfJNXYt5ENgC5yEVrjZFe2o+xhEswgBDWFgSOrg5opL5g4HUTD9Umm
DCvcCebx/b+Ql+Aa+mJOFaYDHHrCzf54lexFNzSCuNmtkdQ3yIW//m5Ndv/vMkUao5JWM6OOBJ70
jfE9FG6I7rxOkbqapynDbjHqldPVCHSxLI/rNFEUcXteVGMhIcnyBZIeOEOdRqrtM30hgSAcs1eY
h0QEaLnsjB7X0BOhBGpJT7RqYGOvkM9jmM56lvnzFsFhseXjlLwuss/4btyifUwZ/iPoniNAwogV
Htz6v3UwAFWbG5/ydNfZUopSSrfVK9yhWyWlm2Mjw1Q7JtAWWSDMilXVk3Z++6tCWBUuHsfB99Pd
NirFwcrU1o6jZVoY2/ALnFENUCbgGTYUiwhCLXJvx/YpL+ieiI9CWwzUnQqHGHlHKQGx7QqO+n0o
QGea/3sPbuBKlJmj/8MUr+98yOAcgDtnBqk1HsJnVBi+aQR8I+BxW9vZLsUDSBVacxHW0TKiRc7l
OEqaMJLgiSdVqSSKItDcmx13fHw+hB4Kd6zj8XfY6+VNo0JQfYEN46NTrFWy5oxo48b5sENMWgj/
96n4u5Ts+m30pXtTBns2jxIF4wHC7bTUiKRZWsC+rxmFwMdJCpl86gEEvKDsgiCzL517wxU881oM
N88Ph+aKiEusQMx944l3fF2Q22AouQoyXoIXsR5WQsdcIoDPOAwztZ+mDL22pE20kKZ5QsW8MwLr
aYMukYKlYnSuBH7Hbx1/Nrkb40wC7VGnT7P1Pt8tELPBKhpQs/Bn4HDMQB2/29m8H1EAQUargL3f
kPwn7nRW2fkx8wtUq6hq5qSkUnmN6OGv6sRcMNSf+tbvNtew8T5yD3EiIC9ytEo9fkFUGFplcnzU
ZWXqTvXVJkhWVfdJ7N922qoHOw0jSBg4XCur1KihpWuja+gdhiJPh74GhCMOojDyggpOAICElX2A
zSS+5p1R5AsMWhcoyAIKveELYv3ZDogRTzbbY7PbhCKG5bZT4j+9GBz/cZwE2NorGxPD9T0WEmU+
O2HxIbwWkP0QZagdDIsS9+Uc3vwvjwA7rFrZOpOSAmlmtTab8+DLlMy3oIy687uW4sW124wmeqWV
FzNRUnegNcUPL5x1IVc8gtCU+JANjVuICdjcA9gSjYRi43Whm29xauLp3Td4AfyJJ16SRam0v5rP
9FlOxvbo46a66Um8wfexV1ivOOk2Bl3SPAy+/UKEp7PakJFaNqKQ+f8qgvoGVbvXgTx0PPMNFaSB
wrgAZan5rZa+a3+aE6HLTb2xZYLcnWUj5huxk+4DLWJwG7SUTg+ye8CCYBcUCAYjVbttOjblPCBR
Uu4BlLs1pOUoRA+DyjnUsJM8I3a7NmSLQycDRXBG0ndG2VrJsJ6zamnqvCTkPiPgG32KO4gqpY47
AWGRyUUCiCfauJzXOmylFC+J8pqa1eXgI3TxEIXaHWU3mNeYbXL4OpxcL5kL93SDFoTGb3uji92V
Eu0Kmeh+EDz38yPSx1ofRO5gCdOlX2l8uGHJCOo6hI9aVnU555JXOrH9CqhCRjuxU0y+TgZkLH94
451+dOgYLenG0GuS3InJuRfiMuVMU3FOeom8mlmp+FRuvGPKEygJmaCtmJ2rkUfI4McnG5ckr7y5
GaV+wgWevYGsFLaBErZCmzZ9eGCBizxZDELQ1hb94Oa7YtyXF3AFCkmd7FjYKVopVOAYUq/FfJpj
OoTJK5UnF8JkTbGEe2zRLtTLDFF3WVzI1qxlVLStlx3EI6oBlVIV4luBsOlbsKW7bwwDHK0f1tI9
7FeTtr6uqqzEbmAw6Om6iK/mvrdtJ3DRAK749jyetO1FijDb8brmPmHaJI8a2TM9Szi7c+9cJg0q
3zbkkgBh+qR+N1C9gZ00NuZcyaJ3u3WJVTTRUUjxLyYgIiiFajXWNZFzY81ZYl3w1sVGwrlR5UCR
kpz04xrR1wJebiGBLubxsLbD5Aw+8yscGEnKCXORBc2xd0M6sQOO9L8/WdX8tqBQbK/a44Zm3x7B
AMphCxwduP1RhIoQXxZZCww113X7eZBOpvKWuH0tdD4Py0WryC4ri6O7pKyaEtGtTVECQ59e7KI4
/l1hsivqOpjy2Ifas+F5ySR6dE7bFUVl8j/3xjikIOEdk5BvV5B9VGzCntcbrQtBJVDmaFdi2MyW
4XeNaXkqlnEGjWOr8pg9YcZm/iZYXpLEd/qEmXOiwX4BveZT1fIA0Nhx/PbgRMzdHxR/fS7spgkh
Qu0OCVPPRWraqHFaf1H8ZKveKb44C5pBVf36yxqbqBDUfxn/jRTqeYHiWBX0BHYmXQ0G7n1NZGK5
dTLSVhRX03LFH/Jm8wB1qhnjcmmTAycorArwBiUYiWicuKwh6haq84h3+pypEhoT2FM4DBmV7XYB
h2Twa1TSjUie+vK+nOu/nIhcGGWa6VnPgn2Lsdqsk9w4As4ZnJ0u6LfCxIFZCsCXtbTnKQMWMjiL
QUZRQ7blnMkF6B6kD93iHx+LS9AeH35P4rBjISIYEWLCYgaDx+5zLwhiTlpZodwLGSkIlFrHy8EO
Ge/3cVlIt63heMfpbVAlTQ/HA/u6wluf7EbuFawQRf/7u/vD3DMoLtktF1u4W160UP9+JVnidi73
5p7VJTb2TYObu2Vw5CmXwTVrL0SOc7zbCzAl4YiDq2sTP8O3GRMMeu8w0cTdPIr+Bp/PELPhrjY9
2WGvPFUQTZ5UZd13Yd+82MJRbBA87nO6wp8iCuJo/lYcp0LmHRwMslG7bdlUk1ISW2MAWK3ik+6e
Yct6PlDOC4Ewyqwk8m5aejzLlj6LKH5093IWeplAGhUt387kKTXxAE7fAbqEGDUxWwVheJiJwH/k
kTq8yLLgCYbB5IKYWD2UNk1e4dq2LUbRAz3+eSfQZndDXr0WvbxJbsPwKDjhRGWxBPC1h5xPETxM
2jgjK8DPi7eML7tVbXaZ5BmSmU7OhTPUuUvVOoQaxEdJA8CIy+iHGFkLmhp6q67kJtF46nMzCIHJ
YyRsga2RKRtJX/v0ubJJsF9HCh9L/y2soAKPq8n3ku8MawwTsvYqOXfvcD0xZcr3OY1EQE2/G73S
s7/KIyPP1siImn10nvqMag8GUybdMFfbpkaoNYsbGlDMAGRp5OQEk/59C+VxlaQu+b2qHaJpkUN6
shpnH5aFgUt1vOwTvTic+aSv15lzX5l8Zriqdib2G3NZ5TPAiZCr8tj2vqo+4CG5hyBOrxRE/Pic
2Pusv7a1bU9Uy9oKU9+17Xgj7QctxcVV3aiB9TIuPlP65QvdN21nZ7FEMzRrGZl08E35NxNm3V/8
yx3kGfxNaad6HplDUkGpm4SUskiKFNARbEsyGWuMSpCxOOWUnmYCkhNCaGY09qK3BvcBqzqZGp8+
srQcob7YFi9XRiW+fLfHWCxb0gpKikBYhbJ5Df/bScnSWrTQJYo/pB1/Yp+3OUomYAVj+vRYGpFG
Qc5QfXN3NrnrUNtjbeSiPuk9oqHuU0+szhZI6PiCPCnz/zT6FMH9Ko5RGprF6I37rpmCinKXUqff
g8YZVj6ZseUAUb9AVj89PJqT0CmONxZ93SiKvK5epKCuAeQDVdP8A2Oh9/LH7GYBb3s2qsbIuTP7
3oYMtn9bDx6SPKm5CyDS9GuiALULv8qUcVqJjBEVYnBYJDPJK83RTCtzX4t0Rm43WXqx0AchRw/i
SCZumHXq/ik1CJGmzrQ4l4tAfZlkIf5U4vSInr5l9nWkfsNuozTbOpShmB2DdR32lFd64lHDPh6T
gzYjrurHi0U6plkfIfagP9375LW2ATAWFgo2Dk+xAN+eKW0lxgLDaU9A18hYIrouNMNl+8Rqggvj
grW8CKswddRvXdLqSxLLK9ptzBjiHO4sRFRlyu7DRvMkuK7oEqWaVaRhYaRbN9VugbB4KTtBU9Lq
OMewW6V6Xb5cjCr+18KQHKqBNXTrOC8KVOa95QFpIGEneocNTLxAJ0aagrKtbxnwjQFlg9+kZUdF
dWdAZrse9TvsSl05Lr3PmvsLlKgBcO8xmfJE36mXe3yw5VAMGe7QzCzDGX9PWi28FUXTKzPoVOw7
egNIesKvlOiqRanb/XlRGeQp9VQPayvLaobLEBTnQJUNeY0g1DH1d0Blltc/gOvz8KQnnjCBSuhX
cBNJqniO/bUkg2cg6mTSp6p+xE1GbJsccSscGEhe0s/McysumpQlL07mronZMJMKtAYza0cEvZnB
qU3/kh2WVSz03mIAi1ex6XkpAsI/DoH5UPRkZpvA56NB3nCM82NSP4EqQzD8QOC6yH0HwYMeGmDo
ZHqqdg5ZvYH1sE9ATlBxFGznDPFMguLSQWQfOV7HjUCte+wogJuanfnE5kiXw2A9zWkfBfecgM51
c/cc0GyNLbWhfm81m0aT2j0g0rgSXf/evPJt56moYWOilKVoLWkg3f5M34ZKbXMgMWQm7kPK/k1X
3NhoiFlW2lMeqsWXsNmKzqpch8x/pXCSGHz2ahNk7vlGsGMjFiYk8kyyFm7Idu2aSieug7FWEYAx
G0nohm8W5AGfqZRyEHHPcFDJn2S42bwCJdCIZK9bmH6hWYsXIQuomrR9sz63OdhmwXyJHJPnSeDu
+D/2VtcmhP4XQF3iuPfoPQZ2BBhCN6dVPq3I8ogrvDLrZYDgPsYiZceyf88VglKwJUKpBql/NgaA
RBxQ9drvUbBSOZTsRiZvc/W/eYYX1raWhry+mBo9lls4GoksgXLeGNEAN642N4DRMqM+NZO+/I6J
WryK51tSkIc14oglgSTxVwFMdhPZsTTVjOfa2tuB522VEPIlxtaot4h6P66SJgeCgrI7KqBw2yHh
i5X2xIF7mdhM9L3gz+BUiYjyJ3oyWA8SKjtj/3lyNY+I38royMTudC+zRhKWSjahN2GE3aPEnYHR
bxpfLGW8HL3NB6nIeN0EaOcvTZdWwFI/K677aRlKhw98bPQ2jR4wysvomoIwn06t78mKUURg9ZOt
ClVcJUXm87zgut8e+sVK3W+yO/BRHSiTkG0ed5VYQylatpNxSoS195Yev8KsNWh9nMZvyz00vZIJ
qZKHpR7KnziYEpZOYNj5Nh+8noDnJdkNdsivoNVDgwQMfEOgcKXQQnY0pPfVkzrcu1UkYNA80Jqz
WYO8O+/EAgwWpMmTTqNHx5Fa+KlglyrTCKlpZ5GeIzTTPssX3tTv3d1oXLRt1Ew+FNhWuUBW4RqP
Z5rcHMs7z+eqMv+JBFW/UDmnxMF15qHpAQzpPKix1ONL95mPjA2sdP++tKAVvlq9s2Hn2Q5OpZAR
RZm6hgwMAiS0LQmEmM7H2nTgosPwcxnK1RMOt8rbQxIjOBjc1NEklmcbbc+CV4YYBN/+Y03Fh4Tj
TMw+LD6PZKYwqHpXll/UdMKl3XXFV8wjMhvyIH7ubUjv9GS0m8SRvNVX6OQmWBenaQ4LVZuQSSXO
W9tIJTnqd9uKUBPsZddB7UBvw87Z8gmuyc3eh1p2BUFV6gwG7yejDXZw0VazBWQq+s67qSMoMkXA
0ShYfKv9BDRpSh09s5vby2AyY78kLfikHbDmZcRQPKrV/lwGMdeEVNpbcuz9V9OHE6JLajqHtfec
+xaKUoIhXPswHQl70sqI4WScW73KfQaOLjdeAnJ51M3p/2vi23iBUdqBtsJr/WI6mBnB4XxnPaXR
e3CBnRl7L7cMOVs9N6KlZP3F9sNbb0HCL1phsnkY86jpu2FtaBRubHAFtn4uWQPXA8mTOzV+qUym
uS5Zua54zILUHlLMD9RR7Hmed8/vy410GQaXXWLAy7FK+05/xyY5ezmy8D9LRmVErT53Tm2eRYMu
r5iwTJRK0Cu7IrbZLCx8SXaJ1SgQiBC+ilcxaaIVNcVNqE5dkKJAQS8ZuM8jM8AU+7qXc6+B835S
oqwyuqM5jx6anZit9OBEhyrF9bCqU94QBW/pMHyBxLpNxt2qTcggJCvVZJOF13p8n94ogCgG/iJq
b3c4mwvrnWKtZGbdJfq+L06jhgFUaXnB9EGbKlscYjiHXL8hT0F9PReUTMa4Sg5EXs3F4LVofkhO
i+nPhR5CWtbku4cXDBik989E/9/Hqq/3ydrfTmu0RW126ZpO72iT46uWPYr24xloelahkcZ/zrG8
EpkjK7hE5OxYjVTbr/NIVur+G5rEzYIN/HQdbMAPA9bGOSsshIu+QKhHKciXGhNmPtN2Ak7TpJbc
KG8ngshWRv8v9agN46iD9IlCPZ1p7bp8UXpajyM51zeWLmfXvrFQ+nkiffMDrx+VQKeMiLTvmAB3
UAvhLtytcxHAkNMvVgqhHh78cM9wKaZ/rKM+7FHe0dgktSh4NyaByB8o/Bcf0/fJFuL9xr3eoTQ1
GviiNKSLxE5mByHWG6+/LyE4O5hXBZUd06frDggH93WtnacwTKWOTa83FgzTZSrxWQzO66aHcOBr
ph/oZoEN1nAKE35cgG1OizZDWHBBtL4C4WfKMTnOK9l4uTr/Q7kGrKmi8XcqmsyeYgZrNZI1oEQ4
VXS7cVrgvCatM/8I5TGUd4529oAWMfcBoycXOwEWHYUmNgVnoM0UHbh0Vl4lHCzbBOq6R/EIKEW2
EpqlQyQnlKReAa/Nad4NBrMs88MjgCXoIwNWB6sKIfQwpIC9nreMCbwE7FkYgWy6GkUiMWpQVCfK
em64cZVudzIC7+cvP1qnqrcAx67qO1y70IxZ5qcA+np+0df72o42EP5QbKFbyaJ0c/+YIXq4WTuH
4+ESodTne8qSepwcDuozcoNLVFVwiIf+cOyd9n6afpetBwH8xB+54IC5ZUK6PXYTxc7o4qzPYqBa
LkIA5t/XmvfbkML0J7hZrNMcU+W5fuOKOKZlg1q8Oj9zVO2il7uG5kVfRS2r9EqRsGrS9rO7F3Zr
bn4ozo6JLynzJTwmUAC4H1rHX+TDAUbYOt7RMv0hFFtUaWXPNPMCF5zDgUiP1qvBZdTLO3bY40LG
yEWQGrZjJ6SX6zvmX11UDFe41bc5Yi6sM/a1vdjpSeTeFuwxVeajxEMtUQlW58cv+v8u2IFUW+/q
O+hf18NrA8z2uty1uZIhOWygEmbd2UPQt14AKHyynomYl0trphkczdk56sVzTZXIJPKuvr0A30eK
FINsVmF+W15iwjsIaZu2cUaai7WgahywAcEdq14Eky3Sl4/9PtZ6d67J8voUHU+qCR8coZv85MZo
4DGteuJVqjbw/9ykP/LgFXQhRXf+NbLc6aHmPaKT/Hc9kVip2j1MLkx/9ee/oWMr3GJ0KSPw87SP
hu7j8iJhqLqkC2KNkVvQKjs5df9j1twUeapYDvO6FnIik7Afylvgu8oQkZPbxbLOEFUSqJZvx3AM
5Nvyd21ElXLir6u1t8iRLnrjT7MvTrHL+ch+03qTAwLCM/WkZwFc1bib/1+9dGwIaZN4NlDflfxr
lMBxRJCVXBZfpsKsCV8SfMiBMitXjj2LuH80QJuT36PLOpXzd+hyDowQBAfNflmxWPEwmzxagCXS
2YFuitUVhdDhniM/m27MYEIWHGBnp97cOQTUZx+IW+ChmLRUQ/LE17/Uya9Mhvjh27+zVjcz8f/2
qazNMMcCASZ1gk10vRdM5vpNrvmApKUv4MVNz3TJhVah+jiJFMmdI4lBdpS20EeEHMM6w9wRsjDr
E+qhgO/2+sW4xMLemflKEahda/kFFMTKJrRjbvEMjo09/91RyVruwqwAsl7UBFQsebGvgCt1z8Rq
agXp2U5n1vBavR5L6KFY11FYyXl0rcuJGf87evrj4cn8fWOyzTxzh4XEQlTf+bSmZQLL7xmkHVQA
/5Vbn6rYd0sACG2uYC0SK5GLjpFcc0VYOs6/4yYrMSecSiqqLoqwDlebzYPfdwmvrgruM1UgpUJ2
14tOVm6AfLfS6ODcGpNmhOIUX8d0shYkAdnwy6zMyVMceUFsslCBr6mx59HKe5urAVB/RSZ3aZz2
dWFLJs2TzyMK8lSWwU/PG0QiJQ6RIwRS8FgVvDOU89JgpUoJ+SDnnzu2tzTUFzPH1xMWas3fMTLL
4YXUlX5RVmMz47esa1tDwtX9da+ePCQhFOTFAgwayQ5K0ifDVhRnX1wzWDv8QKzjLD3+j0LLnlFB
+HeG+ygxSuVmuArJI/Xx5qQJvadhFfy/ITwv4PIxT2i1r+i4LB/1ki0Xsvs6wvj3ZjPjNRo9typP
cCqNggWxbVLSqtJT4BXHjsSseYbwxG1g3xczqr1wjjG2xyy78jR9nP4LtoVdYp03kGLougW78ksi
94GSQPihpcy/VM1FBR0fMeEjDMtxRrM1w0Po5FG1pMwVJEB0Po0cv6jGZZFs9Nt8PLPvqqfJ6083
E1MOBM7yE5uMb8UJ473QerqaOvLkxP2NiPN+nQjcZNhc/poeiKsryb1xVLuM3rFOxLT6c9fL+MzX
8QDC4BF0sntmwe09wpdr7ox9NEeRZCbP6u4c/92Sb10lcB3Oxg4OlJUI6melxKG8RnjE5cqR4qZY
dDabwMkFCRl2BDtJ6y2KYkO9FbXeklNIuf0R1A6w/Z6fg3yvJMPJozlPp3jwRH6H4WpOh3LNiQrv
A96HbL7dQFTxC5uVmI0Ct/h9RbWBoO8MABD6tfVXeHPjjki4nfEq/GAwoXACPQFFfdHyCE2ZRThS
ae2GdlSgLtJRxw5y8kzVO+KW+mBM9dRbe5lj1D5bpHbepY1tS6b0uaGtTitJHnXgeYcsiZiooGJS
3D/NYrC8VUJLMm+Zo9qZZdbcyGUaB+MPoHpag0WjDaCXRQgdLGeekE6wF+FtYysiLe+ozpSfj+9R
OE4Ny4fp7v4uhzYd1/BBBWmBf3gf/NHqAcU8WVkz1Rd371c631MEP1twKLza4jP9yYV3xWxZZScA
ORFaf93o/CrmzKvxtELM7qumsmFlReN/Zjlvh+U+QFQbY2M60/q7AkaVEZU7UOSFlZbRmA2e9Kji
2yaViB+GeCkTVCIAMfunlj9Fe+shiJb2zDQJQNBLSwfvkMPsSlqfxXWBKTa2Qcrf0vqJFboXxcKQ
m1s8pocQu6LnA8A4h2W+ZPC5fxyCJ+iudSRRSA74PSabPjegm4x1dI6BjBcIb1VWAeC0qp0EP+7d
ZDVJ/7w/TpEhIBwa3Pjm09riiusaNNbgclWtHEYcKxSes8ZtrFBOo5U4S1O13pswzoiYknaZ9V5m
qWz5TlYGCJGTlB/tC/8PzrVoNwNqC2Misx0lNextsUnnpNJxCUBda3GxjRpa+sVdfJl27Jo0OU9j
Ob1H1C7r6wC52CCBHHpWubHwmU537uDO0pxTNFCFJurIGC6m9zfcYCIeVyeeHCYZrJtqSsUNll/a
RgwA56WfgGBNMpiJDgB6euSmyPzwk3eVWpyMEgA3cFBAGym0aPfuB+PGd2RSnQkaRAAPBy2N9+6/
KvJn6Kr12QLS2WDU7w0ZJ23mqUZ4vU0Rw7bfUgfwj7DvaHlplkywM2jFv0B/eFHo8RkYIUynSe1o
LD03qmZ0pzGJuaTKrnC38ypJfst+1uIQeF5b2e6eucqtv8WTlAs48BgPXqG6qADI/DeYEuRmaRU9
43mzfeCjTGL6CW0budt6KCVeA3PxwAy+0PSAVleHPx+GBoO3TQOynBKWJ2OhBUTkCcGj5VyjZYn9
jYM3vBUA8mmh6mKMYTCMfNqSRFL4zVM19IyRADz2hD9INAp0WQSuTdRRF5xpG6FHNpYdlgtCu8sE
H2gKUn0fwIAl5qAOaUriDCb+Amoig2dJgPoFwbnrJdIFOrOfCNw3mLJX/B/j+99Y6jL+Nf1ouKS8
5GjjGEqFM2Q4GW5Njtu59jALTW+Gasqqz7KssG4iz7Ly0Nplin5K0Xoedvhn2p3Mhx671jkjNcH4
9OQsISjTDpq8SER/FSCwvdAI6NP2228lmmUigx7whZkuPIiBShxTPbB/8UxUrpSe0XzKWpjOGm9W
1KJrD/MaD0QF8paPAUvOgWUNAECs0Ca9jupqgnZBbhOLNQObanUXXcmt6BMV/jU4wHnYMSxYWGE0
XgEq4U5XGGsPV/Fm1aVcNjKrCgEjzzCKDWD6QSibqZg2xOMx5r4Oz3ck+4mkpCfWQt/umrHQD1sC
mzMhOlGi5tHQH4YTwtRJTAsPN5xho1I3jiG3s+AtJfs7orcSgP74851biiGmKfkAdRQ2maIPNiIg
zwuRRw+vXLo+wBGCwYj3xnxYSScHlExOGpHwtz8cbS/Qh/8LIjyFZZ1ES8RdlEagS2qet4lwYlj0
NVJWE5bt7/sJujAl+quvWZOsVTpA/LEgF4zDzq6Glqcwh4v0LXKBRpncstKhNf+s07I3LIBqimsT
DzwBGZwi/v5tfs2I1ALstQTnGKqGPckjGL3BHS8YRyU8nn0VOEOhB37QVoGPZYmEsoex+WVRR47U
Kygy0iEQdFfTNgkOq4WiLVwylcBbxyFiQBnzs0Ye+FXqVlkT47q+kc50gd109uzxMWr5gimdxVZE
r3Ewop2V3s3LpE85Ptkz7Lq2auNL8fqziMBEjFQr8rmoPJ7qoMTy4ZhbqhYLpSGhQdygQwcu7cMM
oG1bSm9bzaleCAr/6Tt4wPWnrOsIZ9C5my5NAzQYeFPAG1X9cIhqQb3mwlA7qPoRUdElunfYiFcN
pQ2JqzBU8/icnpLdAp6o5pY2PwL8Q4qnuIDg82FNknk4jC2T/bYW7z0FXdfk9MV6OvaZdykC048g
8FONYVAOeh12eCn9Q7DJgiMsRVtZfqkokNnXObOnPSPqim70+viOh75Sbvt1gqgYF+FBNXvK1WS/
Xlnn/FUSCMAtde3sgBztaPtlzcCTgXPZ+N87Xyo2hGkM9RNnbuNtwmoaSVhNzvJn4yfBsBBF61FR
8BwTX8A3oNu1lgpOySNZihhvFUz42IASXDHEvGJamgalTWu8IZOehzBWD3Kg1QALO8soOrgfR6io
t5iALBMj8T9uOY38RdxhXdp1pgU45ukkaO5Tob+r68/a7PZ+mWQFufkeh4QF3nUWS9ao0PuCPq4b
Wd7HnAarcNYnJDA4uYEXtrqHE+StBVQG5XIuWbTEzrkrKMEjXuEq230HKjP6H1Fx/SzsSvT1eJU5
1jPmNLbXg2ud8/59dUQKcLU3xPcLkVOlJ8/Cs+tsf6e8g13fSjegnbJh9VS1v8yRAPnr1txcehrA
crYF//+s8H6ur0d0+Luhxz3dwlT8is+RjJ97m1cMLnCMgQGeEXJAZKRjeKpgnT5pskNOlzb5ZOhh
+4BmAexGPh5kzEHJEC6IweHLKARy8bHVDVHyxoggNzhXqkFb4JehxdOrl6GUmXQNlvK2uzeGF2P1
ssODXCwC0U5DnEVdVE83GfoXepKi9gwENzhSCeNX+HYn3ikxVzKR1FUz9wD2yMW3MLoGPu/qbyf+
2CLA2DqOUVHx85iOG8N0hTc3ja956BQ6sGjEB0VYndx0uAAlxSNqfwjCbKpQgar8K0I7g8lfPSJz
eFB45zKBmQa5k7PnZdYun9oDtF1Pi1R/xee2DMRUQ1fjPvYiu6h9yS/dTGuVs83mrSnvkvPNLRvq
gGPM/6TjCg0FInSbjG6zZAK/mYYaw5uLOR0RzWM0ghJQP9oKXC9guNtTLN0elXunBJeRO1EaqcUP
kpxSzv/UKhhmSSVMGMGXJ9szN6ShIuRRIYocJFMSHStnenTx5OyXhb9o8Zx36Uwd81BcriJi3EYT
shRbnv/L2+gsm7hU73sE/Mpa2FS817mR1xcgcSjvdITKQf0IxOv7hdnQHMXsit+VibCzEsAi4DU3
BXAXWeMdh9FxPS/ERgDFbHcQzNRO2HOqiKqJSaVHZxhQmuqSXX/jjsH5/LR7b7J5vk9MnD47Qx6D
HceOS265F0JD7hWUiaadP4+ieWm8mW1IBXPvr/QvIxxq2U2mQKRveETwqey3MbmVXKedb/2X+fsv
uT7YuKjw/G0QDdf/95Os/HQ8Kopcb4IYtiJYIcDtxrw2VsstSml+UCNevQWPNX97wXsY1ADuPhVG
mJwTaVIRQCvwD2JYFmzl7rwwBXF2ICVvqRG9i6iLnFbxL68BUMB4cY9duHzdcK3cBid2wNkxQV6N
t4s1S0cUHB3oaU9xcnd5IdVWoguNitiKpyENvMl1OGx1oHFQDxpYUNSBFbWinsGflIXCVQ4qGZrt
4TFe0WgZtshmjufGcqH7vwZKc7EqoOV2HBBG8DfLFApF0p/86XlPfRuY0XGr1QSLliVSZLVlMA1A
WrK3PhornzlLRhpYB4nkVS3L5yRKSzoI5F5a25B41zhunC7dvpr4r8cg1onzuVLmCRGYUXfFk0M9
ixtK3nJw+PCnbpIcNCI09z0db+tEa5hnBb8jnWBrNJv/1kOsUEQix0cNQ5zGirWJ8vSXN6U2l/Qx
Vu1Eb00qTBKC6TogNZSXifrUvLvEfJQW4kMwvzloQkzK8BoZRp9XmNHdBF3HWeFnMc0lXcsPM4IF
WMHQI2NmJG//3zR3orFBfK57Q/O9jqi3Lk2Hn1GydsbfngD7WA5DnbAVt1Q0BzqxR60S4CfQBR59
fjD6B0zKbP6n3rDfqDn5+6Lnvjl4G2sk4zAsYb5XlXFHJ/DKBxrGCsT+igo2XK0+FiglgqfXGyl+
jSwPwwrPnpvoEhuHWOgOmRSKP+CAR+/AWA3ex0md9/97ag5ursLS1jbaBhuYvKrXZEIo5waoQwKr
+RSwEbdYIOGnq+4ycIS1i6kkK/aa3+2qX6AtkvIsAJelWg86u00Llo7DA8KKXxt2cQY6DoBoeG6H
odZXVYcJuUWqervTAgpv6kuYCuugLHrztJ8jwqqSqMqvsL4M1nDe7s7fY8KTtLM3d13d5M7snXXI
6xz05Hy/ftqb71D3Pt5zfeTBpCIm3PZWTUuNzZGIjV3/ir54lHj1rwinJr7E9FwPnU7BGqRtVIGv
2Vb97Wh0V7cLKhuDClAuOZiM2l8ehBuzm0r99zmdPmoEEnkdqYY3QMdpMJsJpp+Wz7uSvIFfNiis
6shudTtV1mBgmH5i7sqularwgYOQXKrMPf3onGlH9W5VklFDOJBWyjpADbGLd9FbWAzndDR3s2ue
JtNl1u/H9Xv7JfzLFKKDvA6DQy3/GoJ9a9U6MtYDP+BQMjHkX8UotgEjl4SR0/PwPAhjJewLPuEq
BHq6CcIBfkQ9X/9x2IBHRfwA6Wg4W/iv9D/p68w3b6srnoBU972xtaf/C5YX3RZBZqs9RRROcrcH
46tbsEWJ0+SAavHSgyYYXlVgEFTCAA/iAJgjTSmVDvjnLHTIlI7qO4qNRQzDfLgqjOpbRvdddIwl
PSLKj59FNQxkpQX7Pac28AJGICfsOLmBNhuVqcSWq1BIMVOZoM45NLQ6jB32heInDchb/sO+rSYF
FX4t9b4Jik0SEbfu+EmICvGdBbJpYOUGo2DRIqvI5R7d95yrBwArsJ7wl0oJ/AvqdiKm1x+8kHUc
fcaKaeb1B2LJREEFohYQ2hJ/m0ILr4FlifR09QVH5ADqvxHg7bldiGjywZrjuMuBlm7C+IXE5m16
UrzCeSRULn6slIFTl/VBJXdMT+5n2We4Wl+Zjwv8MM6BovaAcHpLHkJt97gi5bNHDSR60pA2HITO
xim0FPjjzbjXZwtu47OjGCsGOvzP78vofBo7/1n/D5QPuQQ2j+9uFvN44P1YlQTZwllHsbnHa8Hf
o1NWU6kDfetn9AcD0H+ezkis3Dtst5xv0vRzy8us7UjpwkHya6hqy5HeNB2A8hBzWBcRZATdqbyE
rIF+Z/9qndePOFYfhaRxPLvhcFUA/LsMsgmIuJ32OPJpp+6+k9QMCqZjcO9xr2wYS8kOwqrxvLTb
xWAWRbT39osfd5kVrUpR52eDVTI9VR2USpy4WnAiUfDY+I0lKF1u8AvFB5uGhJX6qCuLAhbXV/Mt
Mx3xhLycLUA+wJel8jIJBMOKXHlF8hUF3G8DysTbYWXgkrnSNS2Z6ptawmCZ9Gb3KYu2PCcjCLyv
8llkSAR+mAFCGB6w91guISWg2QuXmMyxfiBARwBcjXeshKRfTemP/G0o5Fz3Q9EW+c9s9HPQALA/
AZzJgAS5/EGXQI8c7PO6fffkJLP8f2W0hn98V12TP4V4kkxiZvB2yFwZxV7K6weTtLZsihQDWKN4
nc6BabpKjx4Thc8KOm0esGi1Vc9xxMIIfBjnmIqkZHN78xVzJoA8x2jW83mYEW2uyLo2RIKeiJuT
yqaJh5N5WOpX6mBn3mHZ+xzewK9F+NXLqG5RCjCJrnfa5mFHXMfEephIULuo57ZG4tqHG8x1kDjO
2SRC/eqh+V0VQqZmDW3q/uto8H8nsBqsT5A+DwLKWKe8ta7DBhhxFJF1fjTHRi0gmLhIYovqSMY9
JlOEthHk0Xjv8pngI/VPW2q3TTCTgKD89ZEVHwtz5hWIyRmiug76CbjBFAgwCt1AK5IheFWDCnlf
dYLYpdjq60B2ozWQ1jyTqlgWGhIskp0cTnN+W+hSfOF6G1gUGP6A2VGaNcwQ7ThuQ+dTI+SyV2Je
B/v8u2KUxmlRELkB4GAvcDJ1qGL1dnwWGQ9xFzuqhZ37JqvoqTNOR5ZUvL2bv3ncYXcT3V9REBkJ
z4PCNlKzyFSRjcIU/yrKaGHReUgnrF4jifLn2/6j/DlaC+KnLR4pbiOmsDFtfAfkht/SEwdIcsrb
fb09pGLm7yCgkiJPLPkF9uY6fsefHiaqLzbwmyEfL0IHfAnHVPsdU1m6e4w77O8JgV7nIeva9slO
qMOzI9tc6aRnSPU2aTDVKXQHZbO6COA+poo9SKJBidM7uQRokB+WwkUuApdtcgRucPowTXbhraTO
eRZ8/GYHMznNagjyy6OpmJv6AG3Jbtxp3FTviv/6yqPnCsoh54G1mUH4DpRpNQ13oTKphZnb+myO
xuKV4UxfY+u9+JkrA30wUTldTBMyDw+xAba5bPOhU6m1hiA4zLqpiZRBgG5TSD28FTH1g3CWtcMr
jPvLkQt859vw2vFq8avsqiJQmkAw2RMFPCZ36xBjcKCltUBb+9K8ER6wEiymuKhVLTc0UR9QU7d0
v5a67CBGKAvE5chLuYRb6NCFtv9EhlaDXlGz4IxAqNB5XVMoKjLCMW1zgxjK7roU559AMBFmBqNj
P6SIMJ/Co+DWGDJ28g1qRmOj/GlIY8LEwzTreZT330dBoba4AUnOe1svcSRz8LTWE1//jC3gy69R
9dpMtPZ73zn0LT/xptv9Um94uNH3vFUiroRyITvzigZ1Xcq20Y1A6u9qOchDMPLlGVhM+TCz4gWX
G/SMTFD6nlaYeQNZzwTotVXY5pFR37m8RbuM893j1ZgXwAbc/jUPHkFR+fe+z8y+B7KGJPS+ON1D
+KSVxjW9LDBUte+36ntR+BSUJ8I8k6jnmHbfMNPS/HhLpBfH4xbeORLyMq7kNxs60maOSYa5bbRq
UnBzbVy3cgk4iXRJ2/PZFyBMueOjUKwX+lhKc1PvWjVHUrL1gFev+7zehpSMCildRUzxlaM1K5my
wnOv8DOSCyQWdKp6YVxApxbpJs3aV+3nhJjXpt+lmU0LIrE15asLjIzGT7jJToDFMvC9fLeNaB/x
j6pG24NccwNycKU+2Dcw7LhmF/rbNrKV6qsqC56X2D2x2F4JnJDvHZiDNTaENI9MCiBPguXSKYA7
Rr02hGm+jUekJHSdpbwx3W6lAenYrieXGrFcaviBbqJHDLaPzDvrRzwqb4rT0UOCOdedJdQlCngb
1PZG/l6MjqpQuSVOoIjuW5Wq7V5WtvfG3vsnDy3DyMzUjy8UVkPlRmL5wNgFNi2jQUe16yoSdZW6
7B3RhELyGTAbsa+2prU0+DU/PBXB5Fxi5upeX2WU9i1O98btl0QU64xIdLNqy6FOu8vw2e9wphwx
AGSrNWHB3b7eOuzUAmQ4ieXpBfbKeFOcplkmEH+q0iuhXKcmjofW7jZxI2cQml/zsk+BLB6DffaX
uoUKkxinSKiGd/WE1u0DECTYxFO9QtlYSXsdFiRIXRUTFvAcQMw2TS3jdokfhPYy0m9ekRtyxSlz
RnD7MbwnTL5qAlr7jAFRL/pInBbL62XNllpGQu2LoWw2rbnukoN0IenugWCboRm3Wt4lqWU0edU8
irIMGUuo9p3soFIPk86+bn5yLGjqCjBUUagyZFXzU2jjaimsSWhw2+5STSHTtrDH3OBfW/naKIFo
uXKMuZRT7eGQ1QLyhWR8GPlWq67L9G1YlrVG2F9UocAwUtqn13LXI+5sPDJar4w02IWvpOVgAlVl
/ap9mgGCONqOHP11flDLFTDks3f2gXm4Y98vcccsMDY92FUb1V6Rda7/YKsqFHZ5eFuZ7+93QTi3
DPKpOXWpOy7P4KvU9rSHEm/nduOOrzUTxNkLtxVCwPnPFQ0vCs1sjaU9mIeqeYf04rZuKc0xWe+V
quvlGzwcUm4OqW3jJYn8qzecoMAXOw5fjtNYlfX3I+XzpEyddVQKr5m2/XQEsuDOqvDW3F3fNYyX
luuJLpCCrW4oLWmGjYCDgxc8rKUGPlvFAhh07DDp8mV2l/Gy0uVU5XmJsvqy7a7svEblYNxoFLuA
vSQ8r2W+OHIeeRTtU03VRa93ndLXd57MeMYFJGd0X/43WIAjPfiw+r676JGlmI8qZGGDyDCRe6QZ
QBcAeHKjaIfh0vUfq08AvRDNtCeV379vzSO54JHRwHLww7OS7v5D8tAL/xWYxeLPrRDT2MlpM9Hy
TLYMz8nEREVHzzagpFi1A99lk3ENgBknY3mDfNKrslx8GgdQ8ko+iftHVAyr8aHZa7e9WNBHTY+j
iKPkEEqoa0a4JzfCqArlv9gTICVJE4CN2ocFvtb5mRpZrcKTOWB5RFEIiWSwNA1GEmz+PulrYESB
6qUGnRNyQ4M0aFJJq7788vHHTl5mDhI3KuqaaYhvTqNa17ehD/wWD4vipziCviPERiAwovtTKphP
sEVD0LHpZ1LdIfZ7Yy2XUWMnXxIc+zrYlaeS7aXvBMGeeZsX9tcovYFDDSwoNpRK3mpGZEkHFTj7
CAESBSEQRqyY7FOQrNvBr8f+93K4liIS6aEK0gnmY4g8LJlPl7ixqx28Qoa3k7YBBy/huj3G0Dvq
4nc/QbbHKC7YQobL59ZfDyAc2lPk6wVU3/aIJOBmB7DcOZ+/W+8aF9xTgR+OacszqfygKf5r+Gjg
yQ1BPasRyFpq1LVjH8xhGUut1rkEkLMm4dXE5vwMC/FR+sDaLQ0PBdpemDBmoLUVJnkSUq6osjyd
0TyZVdiwYd+MvW+VhGTNWYD7o+t63c72asdHDhpUlohZaF7/ppbJQWVPYMgsEAFCkP1U1nX8UuoZ
vu+RPy08MvDVSfloYAjD8f/wVdBPU8GSfr02EsO/1WnI2MgHkATQ0GwpxfXXxQJ5TAHHAON1Ia61
Ep9vp8/ewGYg1KWWgUX8QrVra9JAF8NanXhfrJj797p95H/m2pod6gqw6c6CvA3qexZN/m8EmcHc
662Mw7Y4mjl2a2zSZwDUDcZgM+xpyiU+WUf6VdhYwFh9e8rb/9ZwUS/1eF8aK6vcW/g4AJatb/R0
KwVdBs0VOWJbDxXgXda+VHODGQ0GbDuHqNs5ANW/QNRR95jAj3WcUvDBJ6kKUM4xklDowz37tQz5
uvId80NTMLLruHtRx/6Lxor5w6MHQljadyVeirUB9Xu96m2UddUhDwWuEnhS2DE4FmdZzQ+a1t9v
I40MQtPL1grpyk/M/wW3xB/A7HRGYIyhNednNPbUk88uOOCgirinYk8Hn5NwwMDQwBS1TY0cV0I6
e1LqJc+xzFsPckTRB02MJBhL7zNUkgo6VAyRUblTR+zIzdE686J+A3rwc3HxNVvX5UQjG9HE4Xvy
5v5lx9SXuD2dYl1P9EGDAg7G1S3DNSToxCaswsXbskCdukPZ76Nw0unjlDm7iHgn6cJ8HuTlEKCY
1UA2X59SXKpRfoRPk+CcNTULomUrXCXTt+nvyMl3Qiu68U1PPPcWNpt2IdEcmjpKVdj0E0Bv9mMy
ikxT6lJZDUzGoxNWb5NLfp7OoEtzUqv7E272kPAnNJEuAOmso5u+jNMQ3IVAT0dsteVSM5kGY1m7
pjyqarr6IrjSx7IjADwSgQYPmLgSt2I7UcP4jd69Zj/d5t5pZ72hoFPyu+n5sP/psluT/VdixErS
5wN2HI3z+aOxl1Qz1DWfyKYjRhmQmzFHfw8OGGnv9dSDQEhorsizRv+VOadUwrwZadN3MmFZPKzS
QpvLsRSrA4jm2IBne0F/1dk34sKhpqThZSeUujP+P1qxLamgr6qgpQ1abVRzOdJh9bKOUlu1N4gw
epJR/ZZ7ncCmVXBYpjjPisYROM5nLmhvKtFRyb2xnSP46VO/Sz38Eof+7x/WEMtNc+q1Cy3qLACo
5ZqtDghaZyGGc+jfMB32ASBChFDtw5P6jAaGX2k1V/eBBDBBtowcy0LqF3JQVzV4iFwW16/Ul/oZ
R3+MFsgvpUfMerWCvF7H5A+7RR7Igcsu1zaGFwYrDD07Spi3mCEDzH5k719mkOGiZryT8YnGOerf
iY0HUSPDOO8VNNbyUJbXexWcPa4xyYoF1djcUKI9wdvQSF7EirsISw+Tw/BpPidniKFlQUpVY203
MwAbIIxUBzkFQGiBMWbe9zTphgqfNWM9etn8v7PL1pAB/pl/iP5EU2KkVWiCXZp7GfC//uotLnIk
Zes6KADQPXteLEYrXtLQEK2hzcW+SLrc/F69o8TIRuo1bWUOc8kzBkiyEcu1hdB/kZPZihc/enWs
4SIx1sMkxl/Lp0EckQVr1p+a8RPw/MmAXi+SSC1Fu1mb2aRbZLlEFQmG+5lR5ly6PWlQLz31EpjD
edcwBCjnMHihUI59R3olwWN6BfPkuBohup4D4+YLJCruo1F/BHWSuQrs6uKCtbH1NJalJAq7DX2d
UdDQrMNVGx1b0mZ/gYoipRKp+HIIxKqkzKhz8Yt0dQJkQ0A7x6mv8xB/f6IztQomB0G42IL8PBuN
aFRZeuboPnhvHijgnKX3HK+UXexxtVa4edFNgpf5ZmdHT/wzxPD+pm5nh4qyesEhWhzFWZyEYZOt
yny1g7xhp3K9lVnm+hlCGaSk5hp6rcrfMNSaIySopQUbj/Cr4oo6JZdYt9VhCx+qdZnni8hmMkIS
GpThIBrbXRFwF7mUA4hZbm7RNUkGr1Gd4RkRVym7bCmbjR5r9ZX42Pr//y2R79wXkygMif/SH/gx
NX+GD+N0kBqIJgO7O3T4ko4AiQvZPTxAlLdSRb5V8BJIsN9bdmFHkuouZYyETdUjC+jEnbqbfrxG
m5/1Y1Ih96eeauZfZ3KvNqXH0KdcncgFnOxDQ8QrPeDUMrRVCX4pjbqsJzGm91U6ktkkRowl7+Rt
yOlbI4ZlzgFWOvbuJoXblDDiVrDtLUrtT5mrJNcLvEBIAShUvETeCT6PsNorwoSdu/nli3uUDT5e
A5daK9h5/i6MYWkJLQ3G+O2yu2/wI1VE6kzznQu2asn6/pXunpO2dklII7v/MImGzvILORAf6VSj
rCejci8vh+XG3q6MR95gPJViWAVfsJiKxMMAwGgKrKy/1rBOZmUDF59+VKWLR3XflD/bdMalqr8X
4nUHM2NC84N/nBZ37RXFOe8wkByqZGXyDVa+M82+OnwQi0YXAOv47LW0db0aqXSddjBz1a9/Lb8Y
MGkyey2xCpSKuEVszsTtVgjPUs55yi5v7onMnoiKwUgm6YYeax5HG2pnmHfgM55wvDDEPEU/SmDP
rm41E2PEtMDx6xcg5BW6R/Sxmj0ySMTfBcYgGs1DaiWSbLjkH9CTl1/VxvM4ZU/+XkF90H8N/7GT
Qu1kni4jyaqOnFpY6tm//7AOfvC6f83PX/pESHILdXLRuWDMozThkzuBpZ+2nlPcdMzNQojibMQx
cynvdVXypiZZP0NgYNYzp8FBzb5uhIdFnaavOur/wCQHx+Hefz5nl/mrjfjGRBM736IuJdosDFLV
OJ6T9vHVuetv/b7J1uUBfHD3My5TCJ9lMPTJ37IN8N1cIjFxV9qFsWwAMl+09iL2tOJF4N2Vv2RK
YuUT7qzLJYNHJ0wKfET1ilATpNxjmUcgflSeqZXVhHdzWzyho3fbmRUbWZ+qW+OMHqrciKMMBZZG
u+Y1P7519RKCmpVVGQf+MV0WsmXh8zmKRTAhUiBS0T71WgWcJ7noRhLek8VQ9OgnIXKwBxZx23B3
pcNgQeI7tC1m+PeqNDUpWfzGNlNCX5T7zw5sSPlPlP9W30hZnNgyFXODSNtRV729mph6Q3eFuYmo
yQqOqlBaL+bAunEPyCcFrWoeRRaC8DvPS0d6mJZpiqt0G9CaGC24JT1lsPV9Qb9LJHlklUnkvEZN
yYBriV5smLSpAdR0DGtOTJmlZ9WsgKgEUPzEm4QrLFkZ9hy4VITuPamdHWtZRycMFI5R7hFUxLf1
CrM6TWCva1BjFQ/Beu8CALX0RbbGAztcrJxyLxwM1TCyHc9Av2Wi/439vhWpDK9/XNqTh4xZBYmz
haxtKTEdH7n6bcPmZY5jUBfQfAHaAoVcsOLLxrlcB8z5x1NTP1bnAB9sYOYeAQ9aJs9CkI0OTjY5
yT4XdUhPA8PlInKz6bycXZMLS3Q1IHtCnTsisHu6LGq06HfVpEq1/Ef+T2YByrMRDiXx2Rw0EVTK
it9r2TB3sAo89hwBcRUCg9QYogf0D4bxAo1qpo8jN2lCQyZ8V/PWHpCGResYukoaxHaPRB2BpM2T
QfklP2yglvg7oOo2sg1ntBRtg7Whevz1pHIuYYR63XkQeo1qe/DnmzZC3MfrHbOBZ4SGJKl8z+Nk
UDXK0CO21tmsmpxe9CCwBQgzG4z/s47KnkVaEvbK2aVQfNuNUupc3joelptrwplIzONNDaWkkfVX
CVNQ63acgiMC/PpfTA9hMtm91UtasAR0v1zVIoaOLqvegautBLtYxQ2SU7GC+GCowMXc4tEzfxN6
zaxaqMOacK+f1tCxk9aXoG0NLbaUQVbDnis/iQjA12xF3/4pbEKF4X3HeSdXyvOu0BEmB4yWL0sd
B36a0js/MbBGqlgB5GigBEC2xhhW/pUt7Cb80axMo0XiSe8/Q8BAH7Im3Ae0kIyzH72TPHykr/8K
7M0XJwo76KTAxzqxjL67wkMiDh2m99YjJKN0tx1kndfOioHRO3ufVwOngGLzCsXL9EZBZh0997mw
I4gfxtffeBX2ntnSbV2QXYJwfB4paxOr54jGDLIVQTwO7/Nwsk70jd7/yJSmYR8nV1Yo12D8Q2ih
ZN+9H/568t+HOC1KijsR+sTH9u72mt1KN1bS/LsJATK2oOXNfxc94aSnM2vtZ0bxE5T6NcOiFQma
XY2Sco3JKIhjsK6+Q7o1+mntiiPEw2pggfoZN1cpuVVYBJSCGHQcfPGhwthdkdlPXJNic1zWqwRv
XEY+Du3voXzL1kJqW5cysaez7mQN7Y1Xtfr6EQ7XGAy6kNuUnujMoJsluQSqBm6MlLAlX2OuplB0
8oZpl9JXQ2V04TDhZibpDuBj+Qi+/6ASbkZyWj9PXF1aM8hwouMSpNFw04InHLlG0TNXOmxM6iA0
s8LIHoaoOu60QA49tGaBTCsvicincaiSt2f5P6W/duli1RsfkZ5r6I/6/TXjQ+oH1oWll+pC8VJC
dUsxzXYOQrRBedjp1hzE6bURkOtUxrbTvZcaXMWdxtQEJieL8mi2A6+yllKp9lIIvc7UVVCV+2D7
psaYk1h7WErdbTBga8A9nQq4QiyQA3OWHOdRJOGGwXxWly/vU0NUeWAZLUpdPEsB7JEAkRYm1y6s
tg0sBrsxbsMot39d20ZHVs5RaZuBeJZIww7EgwJde4VFkIJCYGgGPv02RZvfGsUHhqEDKk49UBK/
2qDfjCPt7d/V+Vj3adn5w83c4bkTBCSvwmUOlDMt+4NokhkWjTmgdfF/raXE2dNlBSWHivkJvWLn
hbaNstxXNOp5PSinY2LDK/fhOW//VxhsuGf2L5lh6GWPlfsr4qdxxEdYakDg70uESviaDCalO3A4
U6MV4DKS4EYqW+dJO2emHgLGRASWNVZRcZLJ0MrB7Mfw48EGdAt1xlEGh5ibOOGki0k38ZcBGNb5
2ou6fGz5iLKBsU/Dl6N4wDsJaMNk3orLSxsBFfB1AfPzhXY0mR+wJrGFVXc81g06CgvpACpXHN+Y
0MPLhUXsxS9JRZcwdHYluYvw40UHS7hxg0vCJqI4EA6iUMTerpbCDJhCjNnYkqmVTHAa0zuL5nzx
s5nLdGDMBUcp1MREz5CgT7NjpICBdll8uD42qdGK0IDxYAKdf4Z+C1fvaTJksE+VgI8fE4fVJQog
H4GRpXioszO213Uq5EM4O/na6xIwMDECRo0gyylZKPgEH46w1IyW44lk8iec/YIO7BvZWuYGavZq
0LR4arWp8ygfoS6GtmMrBU+a20qP29TAdJYbJftRI1DR5Qs7gPZrT3C9lSF3efqHgKe2VcexrRMa
F9EytVf7DgXcwbYZCYKJa3RYdukeZ1bZ6aRsdAX9fHpMi0kn39aAhMR2TVhHH05xIXbO6VOAgGsd
ZLQyx/2h8bVG8I7lWHUPI04kyu0AcGsCiOX3hFG6tkbQzD3gF2F723N9F8lglmwmmJSIxU/ppFnU
UdkyAPq0L2rVCMl4opCyC9YATcHzwHFJLknO0H2FgyGPoiP2DpKX2nteHAdLoZ+5+0ceahtw95Z4
NZOAmtDSHVDV7NDv46WzIHxqf3LR4iu4MYznIwSBRd5ghUUUpd7h7ufJ+xWeb46y464XS0Pynx4/
ubEvSYj1JnPS2hmU5aeuaHIp7i6SCRT2T4fWu4lk4PWKnCOiEwlAFoIcXZVyNDTX31ZHlyKqDr6t
BJE1jvnskNOOAhh1B4wz+ZSb6Mu0v0BwxRMr3mwuy7ScaZj+UuxbWm9mHHSsf064u7CW0ixPErOq
KVEiaIPGKQpN34arCYnS3bxd+YZTUMoWwO1MEMc+4uuPSDg9/P1yb0UpfDEFP7V+wNc8Oy2Rprcc
b4+TxHiDNsIxgfM31Q3yAIID3/wiV2S/bOx8fgIpUePvhYjA4BESCjL6YlAh6sWPoTFf3wmwi0fK
cCgK09Cu/rywHeQnHaandG9vraUktUr2/M+3iUgnaYbfHWw7e24JepIVcC8p5LHX+ndWWSzYN6uu
P/PJCMnSzsqTb/jc/MP8198xUf9ve2nxSrytdf7KZVt83SkyOpfs1JLUiOP8nWPN7YJUE88n900H
s2e+on2ytcQKWB072+6CAw6z0L33lET4+FCHLawr97sjg2+8tzGHZrumoCr6ah3L/i70fU6GydUG
c2275qwJnH5VWU8vfk5M3mvFbI0S7rXKdkTfpvjbKZIQqK/bXE8JGySDWiIQ49iPkETT4w5C8hUx
r5lyO4/gi2yMZerBsgs7wq7kie8HPEXJdybnFWSiynXGmotdMRb6AqUlvpa2TkmCLHGXa/2cxu+I
QhlYr0kcjj8+mSvl8n2UeLa15erxb81OcDtaUXgytArxtOasD3GssAkvXbTbaoHOfMQRbs50Mx+Z
6BD/n+oeYD3Tq+4c21gWASnJCpZCGQETFCo7kqq/wJZvZ+TZ5fzXNLI2OZwPqAkmjAmH4Ppyi2Wx
M2RbHVuoTyCxBU+8/JpiDtDxs1wTT5pybT4+dmBrWI+mPErMgBQ06DYnRIO5btGhg1Udv+rFnDvm
3kPtURGWYqBkN4ajw/NWRp73MXN+OMlkc6hfEoGzW9pRhkJn2RMiOuqA6UhC4fYYcC4nwPbhacOX
GxuBFSAV2Ngd2WDuTrXBGXJSDJ9gurUPu5tXSy0BFxIwQoWVgBY7GAB+drQaQghr+JPTYAPBHLSs
XJavs5Rliz6tx25ntA8dV2J+zdFk/mglq0XKyJcI7OXthZqG3xBl4wG3NgUQUZGoGQg0GVyyTS6H
7TQPTGuLpMqHQIsoqFRxzLsRVbXOmXqsn5lhA3/88ZTPgxsPE7NkeaGpX4DhP+Yjw9fTl4lVwVex
yizY1ai/eagHv+b2fscCubJAmIZH4hpgusWXENrphWHdWgFQKGdFBPZsnl+F4nT8xd/oS/faI8Lj
bMVs+T2oegyRk5Z38vjkm/ngKvts8noEjpCfN7W7jeGXNzrgSCItlFlDjH3haPOPZhOleia1vzg+
7gYcxuZHpovwh78tx9UQXEW5ZUogqiNCNIehG0lJyPd2WYXb20DjO4OmrDyKL0yMDJWy706GwI9K
a7MvLvVwWKvMfxQbuf96pcWOVeezUMsANMJAV6lMulf8ra/7+YOoaNWceAIdWS//cnEFrlo34rU9
3EroPMGX9vOXCMJfJVMWw2hfqomvxqTl0pPMWdpNHZ3tJFVjasWhuPFIePc8q+d5y0SN6XgSXosV
r9wdGGOTdyTsa4OoBbruSIA9W3sKfSNedzQoekFrjh3u+c5P83hmN8tqJt2L3Qc0bpVUVLlIzehH
pdnaifW1NdH6xj6bZsdz342gpymx4qsfYNIX7TcTKOWYRHknszq+xY+sgZ56m21tzBDhD1ujp7pF
Knv5x87IskM6GaP46gjKDcYlqjKrAtMN9W/9YNnOO5Dgg7ySQCOGyWoRhizSiVl/ouY+GaLzUtGS
TB679SofKX93zBiQfqWGieHaZOp0y2zpwKEIXC82Gx0KkD3nlNFXInKXIxQ9iApRcQzn4YP2wkLj
TovgS55jHJ+cMo6pUo1YBfKp2hEwY+0cK0TVQaZ8rLCtpktCf9+h1Wc3xU+JPoZqpOScfFTbrQpe
BLaM+1G54Nsrm1ujudEUc2C9KlCPHrqDgtHL0EoTlw3WoNGI+7EFKTAXterqb8lg+5q9RU0wm1KD
z58SZJa3EIZlPECB0Mi6EX1Rva0yFcjMmuO5UPv46cdldK+UVqM3JPITbHTkzS0BGir4zCuCX6N5
QT0c/gbtuL2h1ls3n6UAfIITE2wM3z8UUiVD45bs3rfui2+k2jUnOpf4iuje9l3ZJM4aFG34Ucg7
NH14S1plBg4RstIzD2tnuajTt/jU/RWenqKzh88UnHmXIg6Zxs+ujPB533d1gmVjyp3bjMaVYcjF
PKm/6QNzgi0dEZl1UKMqekKB3Tk4J1Jw9QkeZn8qrqirKsuKP+zycuULM3fQJSBwEzTIhYSg0/nW
GebhnGBs2T3bHiqxLFOu/qDPGbFbK6O0+yJsQcAkfhqHkN9mn0SQ5IhEyTsN0a69GY8GO/wjhtZT
LSkI/kUnUrMOa3IuA9K2b2j9csoPLiu5cfJRzzLtwM31k9JD7BfYGvW/JDIvVbaSm+Rw1AGUPI5p
mi31P7jQgXXk7dDKLQYh7bKJtXHootm9jJJwxbrd4V8EI57hFr1QDZjx/wT7Fq46Q+4riQy3VGdX
9iQTBDoUfKcdkoePwPkOmxjsZoPX2+cgpLBesPE0g1xOdyDh87ambul0qgzKhCLY1lJ2o7xqstty
CYd+jLY4tAFhCs9J3y4MTJg7S0rCAGWCboe1DmkxGGaT14x8FlODx4+rU9E1DFoqPRfq2Qx9vFRG
Mt9b1yfiWQ6F9b0O6ogq/TM5yz+fkH6WL/JsDxHevcFN2B217U8MflMDU0liyB2kRMv4yD5+8lFc
hOT2B6dPMyAbxOJlPwr05BFkM6wKPvE4MICdCb6hCVaYJbsSu/IPAp1tenmisp6oH9yix4EBLx0O
P7cZSV7m+2vudN+VMtiJZegeorTNAv0qIO6EPENfwcW3agvra6evCo8busXsDMOqH4B2OQKoqE3J
bq+PZq92wyw/5c2IC5F4yWDdyU8+sQVjWuAKGyiQK2hzsPYaogdvMrAAGflu1opCEoa3avHqAGKF
DFDCyCyzDQhTr5m7+iInLNoEUaTkU8B11Ld7kpE1EW51uedFXiOri9usdxnOtetIpaRN2XziBBht
gXn/gGqvcyKtouJ+fwR6Fbh2LjeEiyJZWizOFwCyiQ+3AW6BeLQZwdPZhtcGpD35UjTM9uC+hyux
rBKetTd62hIB/McBjIZ/nxxrz70JPxeky/UCfcnda7h8GCFb7wahMV8Bz5j/TqasEeBH4LbiIqyt
DEfbk93dx8SORaMijbwGRmfVTLnKfteeVo2IUeKiaI0jsVv9R3rqt1hRwfy4jGBd/CHyEZ7Qruz4
qDVEwx+Ool9WxVgvQRwt8aZUSG4MxZxaNg8zSRaHXw1eVd2pzuqWCGiM1idAMb6NaWTid9tZvA6B
ThvQxP8iOp1bxiTEzQftqkO/cfZhdtSQdb5ngN0qO0TVyM7pcSwwyzuqamsGhnndMt32MkAnGYbH
a26uDqQHG6293pev6KOHqvXXbsk8mO2K+ltFoZFuhpOTIf465RCsj+CNI8pcuDCfZ/WarftO2SET
wh0LNOG7vV7QPOB8oHXcxRAW9haPLBQ9Pn70B+1jgPbtwCgKMyuTuZ8qtBcwmcQV0IMDtoZBRI+Q
lqsV2PjMpSDM2dyufSRYO3yJCNaVVZYB6Xl48J1tuV4Igiky6LXpvOEeC/Cc1G+zNiaxQDQg/4Z+
pI7W+WvSxCL9Mpocqdjhk0neDJJzyj/H54PqfGyqTbIIBly+XVJLdpqGLoKM3Ze+OtTNBrvwgcl3
Lm9/fu9a9uJ3WRDQnJHQbFB8Sz5fTBN0cTJhYRjXIclJG0+CV4Q7/f9MLqcyM2Trzc1OZnaACtDV
jQQ1hoPJfKdSihzqGpaATuR9NUCO/DZjC7gHKX2Bd9mjVL9UmQdHNfY2Y/ndjlttsFYrgPIxheNT
FfhdHM+e5iMUoBVcLfLsz4HOnwaRAHOrjuqi6I8+wXzYhm5hYjV/7lEFxClPfGLy24A6Qs8+IrhN
Urrc1tLaeyWrWNfeYKAgHvv5HCRTbwfrTSHv7RDy87kDWsHtFrAhAsbYh8/OldihnfnzG8X3qUgF
mZCSjBjiDMbJkaz8DQU25eFK+HoJh6NGWrTVYOPGXQcf2k7T+x1tYcGvkjwbwNW988keLjxyVptV
gCYnpzeIgjvsrXC7sypLbmcPEnEzDNDAn1JfNT5uHmAw+xC7dtvOuaetGTh/rcBapK/1QhD+Nfd2
m68fmMbSNhjq7jiD5RdMjjE7Sj3Z7DoxzdRALZwNqpR2HKgMarFqQWW+4ylYJdFPl7DXzXEYNX0z
/sOSVPlIHBmmeVS0t5by/gS/yYlo2h8omf/qt3gsw4TTjtrKU9kB/6RqLRVts45CzWke4YaB4xPv
aKj+omQclIP67+lzsmWdtZTLu/HWjh6ffTq7Ps9Z9/bNAau1XynmLP71Pa1jLQUpDF7xBmCeUnGd
JyNpquXWXmHNhq4vYf4jWbodUyqretOmPIy10TRwhCFAeMJcoB6wH0jLgj8/vqiRdtl8S/P2yLjz
hUHqeiqxbYsEOXGe0Ilge1L4UefdTzKZG2Er4iiYXEG9o80JBagADL23O0YiQvNIWnTc2Kse47RQ
jyCaD1zpNhAf7xAOIKjn0JmE5pCxPWuY1q7pohOk3/btXKQj55tuTVwos6TkS0/YVgGTutljSL1E
pvlRoYcR+aVRPurJZ/hOGSJnnKgKJTMvPUijBn6f6xif2cyxIxljl0L0csQYws4s94A5AjjaeKAM
leYt4dnfDQd2u3Jhh7J4/2aCfFUrSZapQPdIVNeo6beXNtdGbp//FnrnfbDWrA9x2kSm4uAzJQjR
ryUHJYt0K6Cfe+WVCVIDXCA9MXyJr/dt7L8JRF9XY2yEhSTobCR8mkdSEJyCCWcPQNmGJNyAQCZc
kHmQbzSTcnjF2CPES8pQ+RgcrGdogxfMYA+aRR77g1+bOLEY7k5tr7oL29KioI/yS27xrrYruaim
bbK3mDrWTRV0cKbfGV/WssH4vB6+v5gOwH5kgcbAIlqT4cvd2iEf3lNcwRzouJ9OnWrKu614okKb
dUVVWldqaYLk0/1lbNsCmtIcRadFSizjhY9s2tLQyyqn+je5qJ0vgZP23JQD5jl7IrlRIQV4KFFJ
w/Z4qxaQDYWze/9DeLmCKvtQRgeB/scI93rNaErIzDKVpnNT2j+FWNZagYAGv8ZCVy9FtrGXS3aO
ov2fL9L12YrwtjiBTq+T4K4fE2WlBFDYqFzBDYqkELgApRrG/OtohT7YOrrjwIVR29Y51T1WtDlR
SXjVJL897+c6di+nyRQGix0XrE1+ZPhbQh69f5rdfMFW+24m/IL8+4PGRMzkKriHTMG0DwA8SAAB
uKH6xV87GYNuAZmmNRPUbP/eY0SilM4Hybspec2VfbDoqi2r9BSjM2MQZE0veDAfw+neFa894G22
BzmUw2qupOLHj8GzKIYE3+CSBGWeM92lapuN4tnnvdihZgUQcTmN74ta5xcLeIt87LJP6mEqMpQn
JwyaWL/+uF1Bwa7GQY38WGwpfNwpTlDm5VSdTpLodyYAPAeWkTdfY7ZuAksvMBYmBzuLFLG75tP1
XTfjFNYMe/vVg+GMh4T+3M6txA9p7MN2MwQy5prnt4MzAOrh4+liG6ZaZ8KIP8TLSZWlbLQwIYNS
105o+FA3VSug5uhW05ApYCd1yMYqeJ1jrYv3oeVT97D9FRcaYytnR3opf/cXhxSE6dDMU/S+eW5g
MVI57zjWeneGIEaE1Gf5MSr23rGJyKYMICZBETzjh+Up60vlSdz0g3p5pf+9EguzUEk/oj4fArp5
fE3GZLbSoRbGgPr2fZ0YRk/1o9Uj1P4pc7YSspfKlFsWoM6fwfZAIqekU38hv15vBl5wFRk8Y6xj
HJz6ogsXa94vEn5SB0EeYn1n4VjUabS54EQZrReoDbhQNV7UQHFQwsHxBa7huT7uk9M01psqNQWa
lUXtBSbABvMlVnfkrlQY4qkt0sSfRNGNUUg1UV0G6pE2NUC1YfKw4izCvCI6CK/8jMaThfGkcfD8
lcp+J1+E/oEtE+b+BkzPOgGX3uXRF+uzMCHr+bGakegrruvKBVpAu+steSbG/MGAOt2/9QbW/0Fy
pzjzAKyK9JDMuvggrHxcPllcLR+ZzblXjqV7RE1tEOLCchiO3WRi1/Z4+yoRC32Icetph+o1VPVl
N5t3YoYG/5V4pce1usIjXl2gaQiKcQeuvJVMsDP2/z+Xn+7PYdbyeyGjrvgt+an9EkkWu3yzuiKO
H9GWERRl8l+66nnzW5voTAWaM/r1VdxEUts3x59rfQtxWEd0tSn4DcZFaJtaJvPZizOkk3SxfIFX
fmZoP74Pr1wA7WY+tHGfW0pPQxRTKg8EjTB+vAOO80o4RYQY3pTuS3sNbjdMiHNb2xpgqyUF+2xH
l5O+E1W/dtvkH9eNN+MK+CcKuGHq8+V8+1bFeE5DhyaOjmgnDCKZkBM0HCReXCyPoIn9QqCtdagr
4gq+yAGX/8PRJJHkgk/S0xGCp8awwAxToOFtRGx2rhKbYhR2Dn7zMl419z2Fx4hCaHabCA2DWDnq
pe+/Omv8UB9mZVCIm45rRBwAgY1ktMDfNjE/MnErzzOrB3EajsNBEZVaWElRWrXqSSu0+za75Jpw
N1QmRQnfHJo0Cgu/Kdbb1aSqW0PYcfYN/zQ7xUnFwm/GX+ORophAolZqfTEIqUNAlaG02SSbCeLM
ILGQqK2OhwJTuoGct2Pk7UKZC7uk5vH1Z3iCharbihD5mo/AWVKFwyoX4F2+QE/rsyORdZP5Q8pl
fAhs4W7/+tb9gA6Tey88NvhkocOGTNri8Y890/ErEqlVgMjKObRDw/3pOLPVDOg1pDI6uIvysCSo
2NkabZ4uIhyTpjKEoFe7RRA3/q6JyQwt5b28djEVFgHkfQUDUV34qHDpkXualfTacrDt9Gh5fXEB
3l0gRt1c+XiSTzHVVePhKNXS0KT4Xf6MN3Vioj+TKJysrcIJpuYppwTgahgzmhJxK7j8a/eOxD6/
1WcyNkG18FYwT17Iw4zKCZYT8fxhBU8Jct1X/NGCY6eC0fTs/guelGu7sTS1iiSadXUR5nRYP2/I
SYTeb9oEI9P+PJr1kRMT2eRVnOawpMUJLef/Rc+h6YJ3366i6UCpyWkaVHQSI4Dg5AqXg3jUJYXP
oCMKzjW3MYlh2Iiw6EA/MbjPnMzwV46g5Utxzp2HjXxCnzvYuw36uZpSvEdkI4wOmrdKM3HSpKCf
uQAazDhcSWgGlm+ym78OrkjFD6FkjIjPJR39tzm2ELninGp88L9J3cr87FMI0KfiU8pp94+SaD07
JpJPmveeMydjoMJ71gDahJqo+N15MSNmp3nlljfX33X5VO35Ef29fHv3pOjlnbeki9FND67vIscq
+eSe1fmk/kv6JoUiddcmW7Hbo/xOFWEDSO5bgn5ICIKl12t2Mrfhtpci38ccNp/i69UJe9OjxOf3
sR8NKFPqmGzNkDMwZt7lH1h1jRKagxlY8fd3on0kTxE2wW99KqbPULbjOIrrdI5pE2wvIF7qaRmf
oydzro7S5MdA/Ta48PgsPHP5kdmjnkYQLi81QZa8GTNyqi7ZC+uAkj0Zppxv+f1PldDJ0L5zKsfR
m3olNu1/XfwKpUcV3tKI51XWUpjbJZL+EAL1zkVRb9HMFQSWxdrqUghxvOTL4Lxx86uBx+fzHOY+
1Q8ysll0YtKWqoMpm2rvX2Jc9HBOYOVeklj3uYJQBF6KvaonIUMy82qrjad/CiwNC4mMfjtbTHD8
vfEfebsiELICabA96COaJ+SXQXSLVW8rneVlydYQnavxv7KRcwvTirM5ING8C26PxqhALMKP4kA1
jYivbEth/nVLANeHBSFXKUadVptUhNNKpydthRzdbc41Xh7KSjj3dqMZU8UzFy9u5CKQ9kvGOIWC
vggPabCNVmhqHPWH97UBo5SzyTUt3ztlXNzxhsuQAkd6Nnxt4cE/6fpbDK8tjG43zJRKm2JHgMk9
vuWL7cI8T8fgOBS8OpdzpqCDPBtfBlBKWIR1mcliHz0+7GpLGWQbVJEMzeQj+vo6Ktwzub8CeKbM
lD2syAdArs8HrejK0iZBcQ6i33XLytWG6t0uIpxR6HDsy3bS4K08VSjNP7FMFqULY/JVMfR7ykII
K76798+0SV7d20ZwVZz+MLhP+rJebLmZr4sEtia2MyDzbrQIC97Zf5+WWidHAV4dlImBmHCueyux
1MznO+Wq0sYZxQfU5QQJF5F4kfJ/zus/qXGn+kbHEsUnU0EzMWv8AfKGXew9g/Iw2gxv94ddwGlD
b16GMcOOEDZ+r6zPlQgkY+wdUU7CPTALLWZE7u3CVM2YDJMP5rbTJNXRhiWb/hsUfD7Q1UeW9GL3
9RJx95qWNCo9+0HVBdKRLiQOJHMZ2YVcyu/VV4abyzaA3ZiEUT5LmTCkv+Py49RJ1JJWkiGPmZhl
CVz9YTKoGRwFSghak0bwZo/f/j4IEWdMIoRbHk00a0t9YelWu/+2A4VHKEHfxyd3BVIHalVRBkTw
NroYL3uZbTvzTeMZBLCtdQL5n7uGm7KmFKE6PsFF/0dtJTknJ6Gi3JX67Mrlcs/RFD4bOxmjS4oe
fMB+7xSxbLIYJ31xWZRIc+EQTlyQXN4FA0gKPTh7NC2rE5b4/DPJm+k2qLbaMGBsryBGEj2TzgIu
wqfd2QUkjgpn1ePg9S2k03sGHjDhPp0ctHH9KCu9kwN5rRFgreT7YG2397u73i1MUzIKCpyEcosF
zV2FjcIBswdNtulB4Gi02S51OO95Xl+VF33oHMYL5psgce6nOZ4Q+XX2SZpnacqnWzgK31QVPeFi
XXWJO1ei4ltyfTxTq+9zOV3YAq+HT7fKM2avKHyZA1CEn/Dl0M10QiD7XsVe7no3gKbP8X/TEi6E
Qn5+jh7lUXG24M8VoMgCCw/Ork/pImlVgfYguNvOpfSWBke4X9agHBUeG7F8pDy8mEjuST2NGoY9
vM4BEgcbLrDhWsDncXV7+bW1m3j+4EELoSe7+oTjvpYTd9X8pkuL3h7FQLExVaU9adtqH6F44/a4
RWrhj01d1IKeL5sNTrXpRP3eZCMQY5sLt9eAjdSi4WNdrp91LNWyncAYqLIElS4ZMObYJB4h0QM6
f27ABfdwen/crX4NzpRGkUT/EJ7fQ9V+FnmSd+zcIkLoE0MfrG/SP1GHSr1IsQvwS9chgIPs5eAp
tWE/m0X8Y6wSzvWXo1ZIyLoqP82A8nWNlnPI20HjBkhpiSgtPgBhomTxEaDWY1j/+/fn3xQRU7Ie
lEI0PamIWB/QMrfdrRjX8o/J7xmEoZawQ+JBwgjUt/d4sEM9ykmYfFUM+skzO48S2uNZbIty3xQ8
GxSO7h6SnRBPjdJhuoubsS/XmDf6K3aC5BMP/6ewY93DYQ8a0MNDt8XuEIRZYgHZfTA6V9cD1qVH
qMDOS6GknLeI1bHBbAuTTgKM8VunpH7z/hPdSZ2W8K8SzGNlBfUeq8e/DWKDlCxhWHeZG03Pf4WB
/Kph8Mh5QG0X7ySlo9SrpydqSKWVTdZhyyeI7jyOl3SIlIncYYb6cOGgazVYqtazzrJKMbqXgOVT
JnN5tXv8eJ0Y85WaCUKvUV9yQgTZ2vhoYbG+BDC4vgKlKQWe9mG/7kbdnwhBWar+lrAQZJ1Y2lLZ
TaAGuW0tqdOJlqZ5OpJWiKeMaAIC9VdFLPjGfWNDCAZ80oeio/yvWgHC2+ztSTCQwRPf4YGW+d72
h6lKpQiOha5DkNySduDXhSZZhCvKA3w46wGXwYTPag8enqdv1FOajzJ3TMhLtzDjt+2+uCq5ovDT
Fx9xUdoUCZSBWMX6pDbiSvhpX7Bk9TvM/yANjw3ZuDlO+Y+uSzIpsTu7i2sKPfu+y4/Yu6onxx7i
ZYityXDW8cmZVL59Lves7uejefychMdNzq4lPYSz9FuiZ9rPdcNkztcKFq/QgdCYE8gZuNdUKbSI
ZUUH75NwXZWyDw9qR9ralvUDFkQ6ZusZINgIii9z9QMk7MB+/HlGhBRv+AYMyJK//jYx6xVWbmhW
FFt3jmRcHqkFjAMGIR4RBgoCJX7gfqcjSxSEmLBz62L7vN2SPbdG30zdqHwjsOFmrUdB+DP8t1Mz
8YSsachKxVdAjsGD7+gg2TdD+NDRo3tsUomR77VToKPbOR5a8mULHrcxLh5X+vjGhaU5+LwqQHin
ph/CuBNgIw18C747DEgeON0UXzkUwETlsLr2O+Uu5MlFQiBZGaNAZP7mELF+KlfGce428C/FCAA5
rBawjtsxdTnWlyaDZfBHB+RjfqEr2sc8ZYKG1eZhtg/NXZy/gJJgFWuZxP3uietwpvH8q+IIf8SR
azPmwH/4LvF/lQMrAFwfhHg1xk8tj+Gyl0+GUMPteyB5SUX1zyBf4uT9u9wOYBravsH4xfIWuBBP
eLzMK46pQj/ydnNg0IrWbQxKNo6Eh7oGFkkwd3W/nLvTW0Sy1JJrcor9gdeGuv+ixUzKS2ZDxueG
1v41bFEdnqxKG9A5Jqvk/bbStZi4EaWGt6hLclwarM5xk2z9SeIc753TtWqASjxSFzn63NwFra8Z
Hv7p6a4PSYq9z+Bi0RpIMgXYngr9gtdIX3RrlJkP9H4bqyLSrjcLunCkQYBA6d6VrCCcbE90VZe+
PxoDgdEo3eHglIo0w6vfR02xpq92QQpLdY+b5AwUpuE2lyuooSUaxVVNHhIGxdWSkMIu1nlACxTJ
pqHbAGcmmm1UOUaGYmNqQ4jtVB97ylGAH+FNIC6diJgsCThxq9bT6k4LiuC2Jw0SzqO7Yvq2ckP0
CmsfhTYDEpgA7Xb8as5tz+5X/JGlUrSa9G4XfENbat5jlpMHIDgRQCAKcxv4PTNJYIPB2SXyYVVa
J4S/VJ2u4yg7fOhjcA1h1klbkMVWPpn+AH2aR+nsyMzw08ozabMdoc7hy2KsaTelfU6/UC7VzUl3
595taFTnx3r7wJ7IUBMhU7FuM9GxJFAtoivw3oU4yIfTarTdGyeLNSrnDUR4A6JINr8XfnHh6juv
Uym5KJXcWQmgbD9dVCy3vFXetmBlUD4QDd3tlaf7M+Cg5BbGzle37sEla8kyJs+oii1vZlDEtg61
NW7kVDGu0QxLb3GSQ/wIRYfWSxexbbQCoGh/YwFZoZwkpEGBoBlKr3eOs4zx4VvTvgI6J9b6hoEM
D6blHsEKlru4mjbL8QzDjweH0OzJtVR7SBDVh7n8cq3c2Q5srRLjawrH0dCY+U2FQjJ/LEhPoNdj
yD/eoWavNXuyKAbYKo9OX8wFpjesbkrzewacnbElnL80kdlNyd8gElUbqXbyJ7F75RDddGMwgDAP
0LdRbvtcqgIvkto5AMWmbLq6gad+hjaTZNeHf5Ofz5ZbLDC2j+qNtHXPJmeT70NkUnaG0vlu1igx
BHhKWodEl4nYBsalEM7nrXbJ5arRHhdTBd7h2dg58LCKOhoHOYXjKPt6yDUH4tvaZfviXhF8WFYn
xSva0Pr1PL0GcAbs9L525e6G+g5YfLb1QkBLFsbAEyvaxx5To1R3i/uZS2A+FHdpAwauPgBxTmWi
axwLlXnJ05Be1A4xYZ4QYH7TSpW5bdYemy8/IyrW0ZquUqHCtGfW3E7+wvqdSL0W0QszKDsnsAlz
uRj6rhp2aYHB/Bc7tKF0fnSC99uwasG8RCRw9415uJGD9XlRGw/D9B01svkCxX/3lZHBLr5LI4Jp
0zIwRd9oQCwne+vS6tAkbz4ElPwXb3wYnD9sQ3pEenyVmedXctWq9a+guppgft8dfxFuOD20AGux
v2D+HwdS2zdDAdu6QPms/xMq+M2RyILQofCIzKwgcoFpijmyBzCg8oLGNY3vUHIbvb1xYmlMAGzb
jOiz/+acnvHqnq+BUD/d++V++AHXZYykA51rCgLRQxeENSvTMyrF7zs5mceUJ8FcFKcUh76stlP4
6eHq7xu0oLtrd770sor/hRD9Fp8k2XOUWYH6HbjaMGorJE20g5kV0U2N62uddc7LVuwCTOcU0WJP
hfK1qtldqjHhCfTeWm0aWrt4tAQNtfe24jg2ahi/iTpaXGFnWqDf8d63JU7gFso7jzypUYIzn5J7
5HJWzgFaIqrmFpDaN1p/8kVKbnkrqH5Fgi5GT/m6M5plzBfnUzhRtcyMRYviaHqBvY/la1Z2SNyi
uwpbQ1u0kHy4pJF2oES9o1lhMyIaKDntKRgGLul9NOkmOo1HJy1TcWoDOJtFUJX+oxHyO0BWCUwy
3MGsYeXkRnjTyqPPj2vfrx/QGPUGsLDSAW7it4rHycEjvHF/J6YiAFV3R23rQcg1EWKb8ZfgaVUe
SvXbC5dMn3edZc26/gFUyDUG7m0cBhBqBj4HsaDTHVg7SM/+gqRGoieLe+gPYp26huV37qXkPM3z
m0i+feggFrwIi7HT2sO17OL8Hrx5lASOaLkEyA3rdUfl5sfpHYQezWelc6IphMcYADmdb26LYmOE
h8PRIGZthi9Ujs+JTfQBhjFhZeVuLfBt2WtjBE2ELBJiqXVIVqKmOuE/HZGR731aRMwf8Be4IQJ0
U0Jx9Lz6+JPnh5vjYAdvEYrsO1GgTXD/SZy1ijFTQdS8pp2SPOR09mYpPE0dEJt+vU8zy6+kq0y3
9bVuJwfAmses14sw0AftgkhmCB0cowdKkPkB/fP/CInr+PoBLq155i8ig8Kqj3uAgQJHsrHms8tC
QpqKiOX2nYRn/21c+vaETv5T8S+mgI053bl3Kg5T4L1E3jloy2NH/2hjF+P0ZpM4SYEGO+3y1yT7
teRFkIlcGH430VCxrZ5xLokrS69nNLN3h3JdrXi95b38XEtfl7YO6huzu7Taazsit8AodxegO+Q6
mv4wK4a5KdEs7WTtUkpztR/PzUXUQPLiFbkRAjdnHRAEK6f2POwUFDtLaIo5zWGYx/L47sTqymHu
mUpNkc/N06MTbsM/0QoKDAPq6N9o5Rgaapvj+JUBwS/Bu5rqdL1cl8amRj1YKKMvUG/OzNKANkx6
DNqP7s5RsCZxXvLtq1ybIKygUUdr5uH9crQ9mUNe3QTyx9L9HAP1UYKwmFYMU7BuY+NuOogKFjzR
7ZBadzkvnFK+W1iME5p9UZdm3ZS1rH7ivy8VSD3ZNfvPE2rXY0KVOi/HI9IbvWDujGmwoAXta2rO
9+jRNQN0YIIWC16nAc3eR4MV/kiBMKIk0F/4p9IwKCH57mwC1Gxb/ZnDjlMD7OkmxHCdHeGGsD4t
LJU7POsgtvtJdCfBdLzGoUxUWXGCg94zHZapmG3N6qyIA6zpVdhbefDRjYTI1m3vQjmByFpuDGlB
P0F91F9kBCt7ScjKgn5p+JbBP3UETHF8JSnNKX896CS6oqsXUp/UqGp6fk5lz4r/EcFApbeSGSBX
drbek4vfXqlJoz4NXCjs2dd8o6MX6XLLO5tgzFF6n7fEKWpyD2T4BtSFQlfqxELuDTNA/jYzVo+G
EWryaeVZQKk/WqoV7SYcfo7Z1sKh33cWmecGDq9yWfsOWNixLTf+dSG1dMYbsKTUavaggZQl8Fb3
olxX0xtv+eMHYLRfhgHMCpeJlTgS760ZvhPE1LAHWWcAcXs242UVMG0ygwus3Pc7eglpmlBZLwI3
QuYZjSiIi3wOMUScoqWuKOtFB8wt2Me+ZzNQxfdTxpdCO0W9gBT7oESgQGVi4b89ZvlAWUP4CvyR
mSLf0+42JM1ielqqU0GMYeTvL3UQsEiRUPOZJthUBaFJ8Fww8FalMdOgw52JKb7Kn2bkCDKAyDQw
xl8pAib4lc8NM/hvQE+2V8/dChRH5aII5ydFwnEG2Mbkjk8PuMf+pOukXg6BpsvqqvNMlaXocYG+
7BLgkL1mVA17liJs+RbKSTsRgj+bbQEgI4YnwfzaDGjSUPbUmvC9NJA9Pe/KPY035aaIALtIAmfr
UwBn1BGGb61pmOI34aZRazu8meVNxDM73q9+Lh/qMBxgSh5U5CMuynU8kHLxHfWUEwdISJoRqZIM
BOxVFS4OrukOlbbN2Rde1QzZp7bCUhONLBSxVabW6WR1zn0Dw//5XONWCYlTie/5gH56H50TZNmH
gIHqdwWeNX5fxJ4Z5JKDi5RosYGh+eqTmxfOSPRn4S5C14qPOYCj2os0NugDy6xaLJExZsF7yP3d
BFlOi6gBooLDFRb0Gg0bzduyzdT/DnRP+It24ITVWw2izOWuLDuz1vziBt9e9DhjTR+1Gp6yv9Tj
MFlQRNwUPnbHzWVecXoBnN5AkKfwbF5ofH349StVjV7Mh4NOzLv/YHTwgE1kob47vzxypY1ZvMUx
gFMswQQs3GdWvW3U3hWwQ/y8d7Yu9qTfQdSlCpeXvAPTackLqfTkQ0oq2VFw/xBzMqcWhbo+QWDK
slDjgvli9/vR3F6WqCUN2A/O+KkayaAFRvfMa8a8mevEm/rAToY1w4Gtkbe0lNKDmyNGJ30WvDrV
ForAES5XQjhBWdwPfzJP0MZLqX7uZPiuBlkkGQAUAQvLV+tAX8BEDcc4b4Xe9XDRz6S/2aOzzX0K
Xt9Tqu6YJLcvOUUHTgVohkj5WX7pUiOD6VLD7L+pzMilMAcQBTPNNH1Y7uxuoPDYGFMjUafGpDHu
KV0BbF8JNubAZ2UAjtcqVe3irNWlnyOJ+AgeFL0L80ve3BOUzVJ8/buc8aVHxvaIynfgZVZp8RlU
fgE3LNwW8VbuZvsBC0JncLrwJg4ZUFCUMcgGsx39xQAZoqXCBpISKEyfM/+Ol4Cv/WqjnHcdNkQl
Un6bKjmeR6aAs01CpXAqjpVHXnecapt6zp4Wr4++X8rNKJlooHiTu0QONAjsl5XPsM0fOGDvzC1A
P80tDVVcDaQN5VEY6kaa+lUsL10V71ld5Rq3o8zKMr/SGtt5SL7ghxOB0Dr/0IT+ULQqGrz6n/lf
FBq53uUz+V9PqJRLk2AavDbXUoNWScLKA3rUj9BjraR4mriD11cUjNZrsS52RtHAiGzYJ6Ej+Nos
WVZnJImvkEPGXq2yhndBnIeiLpPPYeQ/0ucA3s3lxkhbKW+3W4GudQHxXJFsfi6iCoMzoE97rbDH
rn4WKzsbO8CV+8vDUSnNzc4RyFCOK5ENu862E0/b2pduiY0mjrTV+S94lPW/j5N+8fE6p0MJuQUk
QYH8ZhaRHtStlJl+QeWnVvE4P/Ns2s0a57AnDj/JYcINHdNYyhp/0L4JQxUJkTgVQkxlal6lR07D
1EDzD1n8/YsVk/fcEndpgXwTbQ05piovwbN4/tIDpz1u+sX+81grZYmViL/46hn/NQ6BDJ2g4ChH
EVblCvHVx67eTut85axal81E8c65HXte8ujsCKA9wPTunn8an1xFRspWDMmoSLN4AHwBqzob2uU2
XY/dtDyRM+ExEXNm/DU0QC85NYwm/qarSQDnpltoF7uxXnachshXCOLYcrC4Zx2qDxBubRhx7PUK
FCsYbz47vAzFdE5t0TW7EoE7cFsGvbkwm3G8vDu3PKHZct8E/LZThjZy5CUfKrZ7FGmVhP4+5hK6
bOVDGHfbTAnEvr+c78+aEA+8yfKiovNMNbS0PczTsw5JEIGea+CQegyQhEJiP86fv/X1vJogky0K
iMrV/1IFjTw7N0m4RLBmMwHFPlt26UHmVML/O7O1Zzd0t54JhOU6AXkPNKiD0wcS7emPUekCcl1u
O6BtNFVX+ZT/6sVDLWTRc/4STsHlDYo9zkfOTzHlY7b8MhpS2vlp628R55hezfsNizsvdyt8AU4Y
rSGRlWqUqvgKAuHiUBy/GhhQcuV8aGQX9eNfRyVWGCTdWcBodYkCX19mbpf0cz/28QERgBD23tNo
7Xg+YFiyg4P2Wo4torPbVyDoHxmHQn5cgHp++OPy5FHM74y9vh26zmQuExDw/OcRHarpuxTInqdm
1/sd8681ir/oxxFXuifmq/W01QMu7yIM/boXhb7QVK9EP2lxq80/LFiAgczYIJYwlUE3omZ8NcYk
fjEfXJhbFzJ88JZumbI0nzEWZcrlPgV0r4afgdTCkBTEP31qQ7bSJljxAx1JkVvDsQsp0pnqtgYO
dn6wyIbYL9JUHxiPGK2DpCLn0ALO2Yk62w9jLTLdI6OmE0MhLEOeMWqnn8L3NSb5+3Wiq3tKCcUQ
adr7r9GTjBQgxhVRiejl4KZVoLJTtREkTqS1tpxGJdkAYLVs/cByl1qRXuARoe8Z7oKLuRJ1rWrp
PYkeoUllkfg7sDFMbFWTqSmRsw8CVGHhHIIv+j7K3k2s0S1UJI53EHKV8K8EmDudTeeBQLSw0541
V+781RlCwr86CjjpI6UIRWP2rs0upzOJMuSuUIIsNG22tij6idY8jYOnP07uJuwtlfqsv76oVitw
x/F3pWDBb3QDeKlAS8XbksIdvxOCN1GeohQ7lqTX00mvYW3/WQig9iUBeac+eA/avwhgb66o5lFu
7+xspbjIQBBVYwDm8dDdr00vvhrdV6wOCyVkCcx2VWfTVaJPVRoTihJL+VZoC4UQZnu8CtAO3ZfZ
tsVQ5X8ibOVgyd8T3mrGVplHE4etOd4Uiq8b7lbFEV/KLi9SZV/N4leTijIaMK3Q6PJDCdI8+4nA
vgWlonAW8Cpzki6OI6JQQgPurjWPspsXavtw6GIC1vXnOtJ7jRBnGWTCdCRAaFEfwAHU34rfmH78
Hf8psOsgMl2nKsbl8g3qfW40I7pxlLQDtYeh7Bs3cjNFJyYVw7L5519pyh/jqe8TYD7rG2PVe6Gk
lkZn8Db1pvrhO1Bw8Dwy2clji2byzyuJlczO2f5vburFxMo1TXr1SB0gWnd10jMyX+UGT1xGk4zq
Hglyoe5WZuh+uXROQRaFYiHKkisLxnTKVVXle5Rx0HpNG4Z+cgzFKlCYdn2+yC1Qoli8/N23FdJO
WlQT6+s4m2stLPGHKFJFQXRwwXX0w0uegsd96meHzwxOowukQN4bd4OtRWpKpKXPe9dAHFUIegGb
KiigOIRxKNrk/eV/O02Lhe2bxOsuNuyIdY4PUaWuM5SRlZR8MXezVPL+56ShCmdBmX+4+pSYNfw1
bbjRc2EwQwYAhGryGbjx0hx7XD0TOoR2bhCl8QBFcpISsCbQEjGbXxA52XxNcyFexK1mdfD/DDGa
+MAs5uyZrJkQkuRhftUPA4RW1BZIUqKVjXwCxowiHlSyS/RFjErQ3nNejmV5oAh3CktXFjkqPzjU
WWYGMGMHXecrsNM4wVlbnG/KtjdhNv9IqmqTKg8w+I2RK1FWIC0yRJKxu/C30Dl0DsOhfU7FN26A
e72ePLvj+LhlZgco9kISpp8XnwQfbH/fRYHJp5xQZTkCA/xH5vQPKzfarmeuvHqQud0B+p24p6FP
3sF/AMBgE2LJzKJm9tNw4RqXTyi7grcRu0z+QeYU04gBwsP5Cy4IAJb1IvwtT6b2PGwuKztv6hMH
jqFn8wqr3fvR4YjqCsZ02jXXLo4jkMFZcJBKTDgX4AsIpt516WIbSdN0GcHJcuA4AWkGI2w6jUQG
dtoJxvNpA7smNko1JnGJYK3DqO+jj9m1alCi95+9u76ysDR6qrPlvXZFoKMQODv88L1PwqYvCTPe
/PY4WGcnO+vWreu2fbBvpE2hEcqM8jL9QcCefOi6sU7sqAW0YslSktI+usRJuu9VrJbzVcY5LMKG
Af3tntPyY1RTJARsK5ruOlLKsZugDhNcJU4lDc4DXH1xvjqYPMstg8kHfHOlXcZY7v+uOEaOFF00
WM10Ys8rn1mPRSh39keJPJM5zZeLvX7ppboKSno8mAmjfvlKA7OQ3naJ6qmEMyff1GHfQkIrO3Ig
cbAxwzJEH0DWP6xEQQanZTxI3OtqHhaObGhZnK/hl5i5rC0H61QBoBKaXJ2SeLJU+YuPx6qVOwZj
M0QSxnUgS48sXIMLKMjoF8dDSGn7itx8zq5Slqq748rSc46iSyVKJ6gMuqh0eTs7i2jEy6zov2KS
HDAq/6xJmo/N36z9CrYwIuFGLGfM71+oWFHZW3x7XDlDuxP/jpWxvwEK9CbR/XHghkB4HsMbhzgM
nh0eq+vKGmNiWib1Uu1IwTq5L8/s8Rng7yNfqFOGGGknBy8VPTKDnFM298apt5/cuqAPNj+rewzv
h7gnyySk2k1FtVuMVP2Kko8oWV4+JUDn3jsl2nyZ+6dbY7n6FSQkbGBoxX9JgIXr3G82iPdJqdEK
W3TJsSH9rH0nL/TxqYh1AqlE223KRZ521J1wDMDFsEfYIkXIqU4GX014AuI8YIUfH/x5m0fRL6Tv
YmxaBL4BiotwmqG4IWfVZIZmZo33g7OgNn4lKoVYwboqFxw5ltb+BbOe4LqpvMnaU2cGZi3NSlK5
kJXH9ZWjsmhlTOMSyiz9vcBCg9WO4hyM0xXtedBfAVlbUClWnScQVHIe1jKa1untBGfAJvFTewRn
S1qiKmOIcNVF4aaNlvJrsNvAeyeF0EEIT5+5AVFGskS0JoQKr/LYnd23YpYvEkPFH1rRJtGz58pz
45bY7EgP8HNBuJFLPvN52LeySMVGZbtheLy21nGJNaEDwOrgmx9Mm5F6Ncg8YehdyPWzLQ+3zQJ4
Wf0jt94ZI30gnLpeHWvd4As8u+DFDkhLRGPAVJIYbX8LzZ5ksq+S68v1m0vrikb8Q7+3OYULYPCO
IMly5wP9L3Q8B09n5Z9hl5FiP7KuciqET7YfvvVbtB9OoVuxAI2z5WPufgUsV6p1AvoJWfDV1GYQ
nSPxsg8fCR4NcI6gCd0cfITpTaF0NJnQ/NXbbGli8HKkGT0P8GDOb+ix6sHr7LT+cpGquRxgUimW
l+/FAfItPUDT0kPfPLYeFC3NXiFxVIZkGjM0MNG1M7YU7iOwRVOEtimy6etk1UXpxeVy4A+1fW9o
3APtiK6R5UbGdo4bx7AD2w/M1asnSBSzJhVEM9Zj2hMENGr5oqSMpfWQ72EautY9FALs+sZdUmxh
dnjiiEfI2NoxxIJGtdPqS28wgRkkdmJdaXIUFWcVPqhM+4n8HwxK632ePk2uojn+utfqY2L1w7TH
IOO6dn2pvfEusb1ZS31W4tW/Ed1DH62/1fG7+gRjzgdaOowmvPKGQN6nPL6NAklFxmuxxpDboiZY
8wtzi0q966oYXmbD6kmXN/8btJkb41McLkVwP+oD5anxZB6AscPdCcAz6ZExe8S72g5Eu4ReKPZ8
owgayXeb3UYJU7zA2U6Zad1RMqytQQBZ5C5fTkL1belYu6giR00v9zD5sLAS2IxiGeRK+NNIXsR3
a18Z2EZ+6+lTs49V2jZ4iE42z0s3ZLwYL4CsqF1mdxdJQkM/ni6tIYaxzyucxo+wxg3zcWSrPXJH
fJxyLJjP5E2MggPwKLVMQFJvzpN7ZMjMkAtLf0AxCYdB27aNfoQudVy0YV+ze4V39SB5d3n+bY3t
0srKz/sslfsOWQQFtNK2wt9atq22GDfjVZAUToLOQI3dvGYdZL3ymkgv8opTZEtN18yfnM9s3ULH
CWT0qswpgGWFxg3V4NZEPYThNJCZHmlM9uGNkh1sqBQconXRgo5Z+Ty0UXOPD7yTDyimTMFuLFqY
KcVvOENkjQFwxgDOaZwA6Cl8K+KoJKhS2LuQR9hqZjAZXalYFMoNfjRBGDhumxoL000395UsSUPW
v4cL4ipMxsnbTSHvNOeedPve7Nl5KIkFAh+ywDdQgKXqxG8Fu0coUE6b3LFy0XrOeZY4S7T2yveL
9OuxGkp4PMbwpGaI41XJoLfGd41h5pLqA47U4XwRaYE7eU7PeysZ9Wpzuv8YQiC+f+ZoWACpJ5Z5
JKqSPTLQRGmRN+q+iBhqa20nxQfnVrjEL79UGj5Sqw1KY+VAw2vL7x0NRq8ViZvvaUvdN5e92OHu
4TYTu71qXVkvKpl5dlMOVCLHewvpQTTa1C1XlXNcisDJJd5iMjfH6b1+ytBuR0D8QGbS8oollNLZ
kSZGpVeHqp2jxpFdMvCHiCSHA+gcDlGQHSccqIqA9BI8cSlYRCZxMs2y3osrbnhNwjb96+2ZFKGD
iOXpLzSAyPoJcy46eXeUvu+b5lgh3C3U9olCT1OiP1LUVkOLsjPHhIwInKNfJCMlHGBBeea+2kmE
HmmMdWXi9tY2x1qmrc8TJEFPHS5/cgaWLc8LCOclnnjhdHnpjvQKMufBpgCR+lnASC3X1bRLiFWX
5qu/3zrbuzhlTliIZaL5pb5aauL0jvY3BKHW+S4d2Hx3E2jGqRxpmtWKhj8kI/Zg/Mke5CeUzdnG
3cNxSKjhrkJsf+KtEHkoNT2wGVfY5m+BHLrzzU451o5D2Pgx8WpxGPDDGJ0Om62nkMi/3comkskf
Hri1DHo1u62ozp8y5bWvJeqdPg/7gEExj9D7zwmlyT2Gv6Ux0uy9fjcSef/coJfdnlYKhv8rkjQv
sDO3+fNe/dqFRsA/yIChG0FOX2ecY3CajFT42uMVtdHmJEqK8ujp8ZsO2r7udSznkhCQ8SdhFE14
zXYNNLv/kN8M3hLRmKGitG+SKGuwooSCiYfYElbmuzpU1Q+m9sKkQDlMAAIzMja4ukzHilkuyhmu
XAvCzfFC9IVu+BjemsY1LxNQqyrR4wH3KMmPX0IlbHED3A7RYGx978sGf/VRBzT3EOoxJCtwq0pT
dCfss9GMnByxxEQC3lyzMdltmmJRSCAMSDRG/yRvCD/xtqamUkz2skMxohZdzINrRHm8HS7t5+qa
6a5rIUj7n3hMjfcbA2q634/GbGzXzcjWuko8PtKnAibIxVIlc2IVOo8fMEyKX6NojA+WlWs9b7T5
x/SoFYQPI+ewBNWhhrghYdX/OLBYXW3GmqfJ/yEbqhthQSnDM/U2YYnz+EA6nZlDdnPLLAUDXhe6
ezafR8sQjOqZYkNAnzrIK+6xAeJrRYkpBkydmHXIzqfy8FQiT/U1ywO4H3gwsgvR5yoV6tmCcXH7
G8LOJ+5RjQ4KAcFjq5utq8sYOhCcHfOSRveqeCX+DAtoVTSRTO0QobftVDIEdELOIG+MPKYrPm2+
3D75PggxC8UObjWFpwKi4/uB4RJagEYv2lG81h/d5JBtFLscZNRx1Yd+TLeCdVZkfNtFtw9J1iZN
7R03YAFi5x1TsGUQEmJ53wKC6mglZr1QbL1GgaBH/Y33GUdGZe9rtmY5O5PDdii34zjgf1fexfDr
pU0Kf992RKtWP7/a1enjNFhuHqgoH6w/SMPHleVBcDhM8O6HNToK2YhtfQLKxV7Xg/6z/hKnO/zF
IXwgx11S7xM3emHF2h1tsy6aedwwpfntJvJo2e7S1ElCFq6dyoCPiNxdDtr9PTGlHMharWk3JVVe
Be6IWRB04mRDFHWSen0IdQvubwzwNnsYcltzNSxkZEpSqTpNPIYBMYwDXx+Rc1VhcVSpHbB+LKpi
XcVPlkm3SIj9WJbcVJkk9Co+snGD5+YeE3YCVsZX226xw2BxmPX2TMvaV9OIWCk6dFy0rv+q7GdV
Mp1bN4KG2RsFAO00nFQb4P/2hbwFnxbHPb/LECOCT3GKF8ried8jJ4g76NYUk0x2WG6QDi+uprzF
w+r2oDx1z7tYjHTBTOjGILqJL8LFZBb16FMD/fj1vntDMtNQ/Y6aSQbxTsS5n7jNQzhjFpVdNvQo
8F0neEYH0uS83kXTdnIAdftVq3xXRP0AF1VauLTQXOGCuUkVante/KwE8x0ZR5XllkXaonaks5TA
Uxi9/iA9veUqLgfwIPOsTSpdMbDtHY+zBbIK3EjAjw20vfQ90Jm5ZF6S+zq0OLB8GbI76FvZBYoV
g3psbPuQ6ciZe4OMk2XjhjUj9EauAF2TmecAeY9+wc9d7zQYeVHgB3NzI/U8ZUXSZ0EB7B3ehYbv
W9SZLS0hvqEFbJ8x/D9QwsiqiF5odoUIbUtIWU4f7N0LNN0Ed5lN8PDKoMQeKgi7c1BdBgHOsQ1m
+Il/kVImouo5SzVATNSYvt/rg455FGIKLoOMx8CV+Exna4t5lLgeE6c65fpIgO1BjTzw11x5ovpj
/hi3SP67R9MCVowqZwXUEK/CyxprmTlOC6iTwnsLsG2IVSJOPQnBLsztkrNy8xrhBan8E+wHRCt3
SH5vizUcYMIpsZHHY0L4c6seLOL6e7f6luS+yE7XR7fsVfib5rL5lxuqo4/DxdzR8cJJw1VSZG+C
9g0w24U2la1QonLBBnJH8Tz2tpF8TIXQKxK2emow9yzNzsKwR6zXKzLCGK7NlNaog8OCtk076Gud
+Y8p7gQ4K0Sv1B4fvsdHhIPo/41vhhYktxwXGXLVfD5x8U87jnjfdZz9ZcWuhpKZyMt2m4+cgdJf
dx/n0BuHZ3YSGZiL6JPMRw4zZVG9/E1rFEIc57vuZAk6045lupWsxFEUweGcbfV5sxDErOJfpMsO
9JOidmvck/VBGHwt2aHgMUZ2suPzNMoyrVXDl4SR/CJB6p0dji0tL/HtWulL4AEHtecLkC250WMF
zw3dyEq2yend/G0M5tvroJNAZR5oeKY6sBlxoEWlSFx7SCcCAKvxznoOQmf/EUaGjfC9Ue6qeLXy
a+z89SuBAVDaZ5yJmVTkkyg8ADVWkcblr3mgiUjyNnOjMgNyPVumyK5jWEOPiD8c4ebO7Xt35mHi
h2QRC5/NBxoVK0erldPQrlFqyH8plvac3eVxBg7lwd8j52/bSyCwT28ZWBUo1o8DrgjEXFTbJYaL
Wf3qxGgnbFQkGNy97B0aasnG0CE+tf1pyYDKEytERjlbpXBn4vmFXRVwb0gI/nISEyWo4/W6Apiu
WR8LM2LKUc5cR4slHG9n5ONuiBuCID+cwnet1TCph9cGIJjtBS+twwLwBwpIQEpCnZ9h98RZMtDH
JKkSuJ5hZiAjUf4RXGZ4SwlTVY5A3cR3e1bjXe/3c0OaY5VMAzSiFE9R/q1QG8DPIBVaQJED0o73
aYu2sitsEIwtvoFwB4LiMQIVnmmhYG7JBOinqBoeLBl8qw0JybEZHzPgC+nQyBMXpVXb0H9p1P4X
eqzNg/6lPoJP4330cpUZ4s0y1ktF1Yqanz/eWaA+PscvbF4ZWtyqqoZtSbduPRIyAkdQAhqp8f1z
645Irx2UpN51a83h37wki9V6zthhzzn3eH5YjOOTlfReEn2QUtUeL7DSdmoYO3hPqSAHUO4P8DHa
xWA1cLtyiGc9aZUp4K7encBUeSRmDq4W19YshL7xRyDzt+HawduyjIID1shqVRSH47pLryGQ4MoT
yRYl/gahHQ+9If/7vJs3BtY5O9yeCfhnE+JN2q70IhaMDcfpI+oUrdMuqP09xl1k1g+4nlGGjJQ2
T46sdXNKDzEQE9tTyJJ37MfyM7vGg/YQpDiORC90+Tul6FBrJYoKQpyx2xP2qv+0ytvEHQAcXEAj
5jg0CFJ2aKizogPZORz+WdaQoEAmM8xVA5pcvgvnw7NY9OOAPhG5Vf+eOa47SBebZwJIzEaw3/YD
aFcIO8VNER8787xLcS3uSx8iNYTMOtoHnfYgPAbam7VfNrTxy2R3Ohlr6WOdbCB+Fcnnfsfa7DXE
5rfJjoQClz3WZNY4uf+b7D/e0vV0V+ZfDb7M1XoY+rgzyCBJ2rT4BT7KUz9FBmdbedTHeh1Tpc0L
uhoTctS0LdBbU/3axKVCd5lAeT26oF5cv0uj0wHoT+t783hjMSeKnLl3u1AoyQ6C0FCYdwSy4Wg+
qNn2Bjk83AiN3kV/tZDojwj3ZfPiIHckCN6NcCbQlWAoahola+FSIXbOYBSohpmU+bgVjly2HDKI
/7EggOUOzVHLI69poK/PCFXzaaHxg+fU+vxyBtym7sC2Z7gHIlJY3KqdoMOVzD2Pty0aY0hi7iC6
zYSCQr6BJ87lQmJiZVKjdye6/7BxMV8PqC+kh3wZHckcaCzJu2Ls96DjsewT5AZ3d3oJ3E5EKMA1
kajvIHPfQqPgIzCN620lqCXokgKLCD2CzAWFgoyg/sJCHWADZ4Yu8wumGOGVqyxQj3PPUxvIzxne
YypOQtcnTbpqt94WOEHOkTPEH/xP5E7reIqBZx6SF/Y1sD6ZD/a7LwkTdmToXsHGv4WXWr+2HQKY
RjoY1GkQ7QvunCI0+bSQ1uqJbJlTGVsjq6Xn+LLUOsBswpybLK8mgyVFngspwIncjEjJYCws5xrb
NaI5yrLakeW9/C4VpIIT/GVA6eBkirbWPUXt0SON9syhZrzF6SDJgb7OU1opMFzIcvOfSHJtwHUL
J1eoPAT8GhGOn1dntuWGuxO3C+6WybTvxyfFXgt9JOBkF/M13tbXMY2eiawdGrooKuvgNiOZA+ic
4PAEe15fqYOcu/hhDrGDl2Wrva+6sfLds4Yyx80Q0PyiJaPvrjSgbQM3G9fEJSvy81SB2rB8O/S+
92Wl1bFmwHLAOp7rA+o1+8HrdZrWMVbjm+o9gXyJ99R0QIemiY2MtfUXaa3hvjawA8pFp2EyBKJr
DZhxHxBFujB2WLBe/Pp0gkJBkXso8O17ia05ENlKoTqmeb3bo+jX3LdNURFZ3gr3/ktxQBdnyNpe
Z/tRaum9Yxjhtycr+Bope6sYvHtWpt5fJgVaYuTpuz7DGn4XRv/g3j/2zBka5U1+PoMsKGtN2HpK
LhLtPgozW0CuTb0N4dceVvejIXNUo5+m5R4iyQnzobpqmex9rA5fZkF0OzviapZroEGcFoNhy/DR
k3NK7orICOSQnr48W/JHWdIc98473ZYmiP3W+A0g05gc+UoLxpirLp0gr2WiIAJNk5uWeQ4vBXgR
rFtuQmF9kQkE2CPcuJgzJCrKwCstZfLwg7A0eEAKWzCDlmawa/jyWkQkHlYvJGkHTFaAAt+je6Q+
155nog5MBdXnQ7xx5JjhAMxOVnK8J6nN7kUxcCxPDtoO0w4aLf+UqMXX4LlW2rLhHEKJPCGW+qLC
SX8HHixMFCLlBQj3y5fHCTVJLfjsiKiKwGEKD8fmXBHH1qkj3Z1CNFgBWqgAxmJXF5RMyf8NtIzp
14mAmnIDc/qblI03tSXbleKlALhrX/26BjbAA7zmeLgUIqJu4iJdzGgw9WA2lez0BgSNJXdQw3ry
on8mgP2jR0UWbpouMmckBAAqNQNIB/+ozwi/HwKygTWyKrKofuzTrkVA3thefBvHRtrhZMVkuRKg
VVhbtuninQwiDfwWjv6xsZVch8JsyRIQkGx7F4i5QyGPgDkWsNWWcPeUdO7NQ50MVwXxIdOZzcCq
5mZgNDy+hVpE1jm14F/VAJ+vRSeM5DMRCwrv91rUxFJaAPJjLPuqi4zmZaA4CagBs5xGanBEitwz
txmY5+/CfZfjUjIuv7lE0mIqgxb/VPVaoFiEMUu7r8kCqB17FczPueGMQ35ImlHXx95W7L5Q4poj
cSKwuBGYNfmMIRx0BqqpHgQpgIxoAj7PfCVvKdUeRY3ZfDNLooMYSMKyotczFdI+zrGfZ5wdwxXt
f/01wjYifZZFI4tiCtkmwwZRCzhxC0g19Ekx4JzoNGBMZqJGUYlRww134vqNHtuzsmxMK2zHRoFM
ou/1Ln/0bGzZ8lfqXgL2zI61sWHv0/NW2+WKNA8TdebSKZm5+c3Bd/XCbuxdlU2REjxJAOAUpusx
7Mk9i75NwBWYUDKsbJRUGcBz5XU95tC4qPHijJLj6c9bMyW+rVM2+BBMrdiTjy3VUtDCDFU8xjZb
WYW8WCOi2J9Wd+n2Tlu16VE4NnBbo5ehYzt+r10PGjcy5F2IQFihl7JPurMrEtZTX6utiX/5MLu2
jSpXftJKzfkCiA1+b4curs0IBVu8/UcsEiCykj2OgIL37hzG2sJWtKnMRE93z9DZAQHJL0NzymhG
oxi8pqs3XEo/dZn9+np26J6vAGxs3n9nIt8ljBnxVGzJDdznphugIHrcnSUMM1dAVfc0ltp2rD0o
Snhj/HHrNYa5Ml5rB0/KZBqjNtvkWH3rsSdA3eo+TRsm+9XKkCQQydVcapLk0A7uQI9i+eWzGcVO
lKOgSw41np/HN9s53n4IhnGssu9qYPaZktGLHJNWFwsgLOT86LAHxkf59oMDOxXU3IFnThXUQgjc
R0gxUah8JiGaAqR+TVTR1clernLSL/NTU/vrIhIrE5RJxiwN1bdTvxLFj5I236e80c8+JmLaeRs0
PMOPj4bm1HpwUBjF9yBHn8PIqXD+qOTb2X0XSYoomXQVIcg1UyJ6fvaAn9c5uarGZsop4R11RxaW
/STekQBCvkILbki7lcz/KoBrE6L7rn5O4Mg+XTMWjtEJGPs2Gcc8TnzBhYYvyiK4FihUOuY+DHqb
4NuFNu7JClMo7OdlmXPxbE+R1gnYDuqeLaORozsEmaQRPZfPBdnUiy6Yu1nU4fFdR6RBYxt8/vQJ
yqViHqE/1oG3MvFeLwFm6p+d5XvHxaf8a8YWt/f8qxupqr+a74zOXk4W7MQzfgcG+M1roxvAI+Tg
mOX6dsteoAiXekx3W+InRxuEnOzR4JN/epyt6DtRo5Vd9U2Np87jOW9eFz/O5IfkVnWv1Bnv6gRq
bfxTNW1YuAI/nf11fliF8t/AlwzasRxkXSjfWHd/alAuhamZcvulbf8RAGMhvSG99XK+1gYkJJw3
RaQhZOlRASCJnwaW5S1mX8iI61TCvapEM7XEu2bFQl+Xw2Ez1qVnKMVku56U3BAJY5hw8w0U+G8A
8FhCJzkxcCT+8ExFpWzqlfaqG4igiGwB2YJ6bKhQsMj4Vt3TZmZ/m4IaijCcH4XPSD2z5NhLyVo1
bEVvDodEQCwRzn+5ou+cc1dWAUiQMJDRHBRibTC+x9aW29j/3iDU3PIXBJfPcbF+SvT8rKsY5iNC
gOYRAmrzfkEG+WTtixycwuaoTC9baDC9jczad7S9vDHrvildlVtnwPQ6zxnPH/6zC2TosuledrXV
b90L4UDy8XagInnnCK6lN2W8uCM0+CdijSCKQNMgWzfA3uWm2i+/HkfOT756h6pvtx7sTX047WlS
JiInhxrNfz2iBTsZGi6N/P7YikoR3OQ8VCCSC3aYZ9oZ24FQ4HWjx5gY1PH8dfYooZrl0tahBttH
tAifi5sh3fgZvEG6CVyb/fAj2uRbxaD3+q2S0f3M1jj22QdUs0j8R3uU/c8wldnfFi9TSgYmlgeE
qUvAA0U7tzil3XXEk7EGBZYO8ZJBHJDdbzwa0hVomJ1IbYy4ZY0jbfEBtXXq7zUHciviv2S/4YNL
08Me06S8yDac0cE4m2cHtzqZR22IuSBXV7Ub3OHSpf9fLiBA6ZljkBe3Dit5hqvR52x4xlZlJSNn
mFHIhPEe8IMsTttPkxAguWkI5Gyxe7AZk7PylUrwDFUKldGRurzawsr3o/s+Okt8wzDQFsnocBXT
vygXES5WgxemVxNnLWxL3Sle23Q57BJZIqYkpOKzkQ6s5TjJb02uP31QMvp0/Yl/e9eSEFCLN4kK
70jjEYSlHCwC7G7Ow9N5r3hD4LqYZRQEjZs8gE9N0kRW7sljAwUFnOn0dLRJJvfZuuXeAsqAFYTp
Wfi5TyvCOc69CLjdcLVkD4kgZkSTdIHlD1hLt2QSne2uI3o6AoFwU/IiYTBl7oWnuqhji2m1bn4R
5YXnVkEC7CFK8ihkMk5dYv+uHHd/YfmYbOKhi4NaotsyKj0Thqj4QPje99PotZDlHLPY+SD/0Epa
y2RXZkJeigDR63iJOtZ0DZ5OI+alFlW2clttr/1+qD+4qOBT8954gfakQDVy7jrayl6kTdHkQDeM
MjDqFFDF+2r0hB7rGgrXQ4R86bOLi4qvqMchSfg3uT3LZOf3AYgzMmRqClc/hlyEs/731G1bl/Bx
LcwiDNgBNM9xl68af4E3s+cLL+vkNuFIjDlV5VCzGeprD+Vcn7uaN+y2eIamfPEqLjnwXpOeVCrZ
sfM4gUJWKwnnCT5/GM6GbM8AL5X3w17PdLd5ExXMIrgdoNMNhOjfCu8VDFi6oVTkBNiaUh0zDaCw
aIMlvK1ad0lqol6tY1gKC2nGp3lDnP8ulMtcfd88ffHdQMzJZ+ETZtIIgEvJFuLo5JlwJlrN6NW3
ztqjoRV5ljs/ZuxeZfdS4uAky2qEkaPCSTK18lmDiHtOm3sg6dTgRHVMz/g7NrMkTB+vF5KGXKkM
9r+xsuHbBICD6ZH80q73Qh6aVtsaQMwLcJ/cIYVntgjxEXOdvla4WIkbQRXNWthvgqtyhEf1Jihu
SYWCpoHVQPZ+nB5LeJPXD86+biJ9wtrnxJsqBAWhg1jgj9wgqAtE2UWHOQN2NEGxSGGqYdTAPioa
05wN8HEF/serWT+P9lLZwJvmC5474Hqcb/BOWB4eDa4OG2Dm+fyisblkpoMoBcYS4CV7MTF3q4Aa
fRq/ezPSl5r2YJRhbBD5AW4KqBmLw/YHdyuQRHy2cQ4m0LHaqlQmF1hghK/2/QylgfX50X8GBpua
uPxmgzaMjkKW/tt5VQ52fBSIEsc84pUUi/a5tV0N2/EIdIHLs2AApSefDP8tYMhjMg7wPdA/2BI7
BkC5ncMbLrw4RufeuQI8JBe9WtecOr+dmmXsuNwfYUCLPPhg0UMeaMoTkL4hMN+Nwm7wvf7UxjZz
E/U2iI76pSrnrjnDNV1Mf29rD6x45TO0sLaL+LXvcwiacgnQH0aqEfjKXGhWtxcX9ZFty4GZT4kr
LbN/EVw8xg6CGNFVJpGfxwJ/usqO+5zPLGDthXKlJhHY27IbrNIr4pWAFaQTccZOTjvFGsBcd/9G
oCrYUQZAJFvxmVP/QEY3cECkHzi6ZYsKAuAC0M1LNxZy0xTekp2Q/nPotZeOrGfNPcB1DsSW/H4O
FQcl6Ld1V7u/ztuvFrCH5iHZMj6eQ8pSW3pjIdtJonzFazPfGHfrI/XA0J9LROiElHrVry88nrg/
YK0FfpcvHcnnpeKwgojD5tAIDdSHXrKIiU/AuCOvA7sc8U32Bt0fVJF1ByeAmH4hGMi9Pm4no1bE
OjagA+kJWF/+JjAatE1XPLnvlF46HVUtExRqZuW4+/ni1Ib92Kd/hZ0VCnznSFxeVo+aMe2Majmt
nKi2folj06gsBqRwx+ybGR1tTl9g2bCqt/yivBSND/HgMjTPPnCE027znsLFVrUNDm++ws9VOqLu
NAeE2Tf/N0XaYK7qLz0R3JryXctx7+XSF0VzuYLIjuGkVouXcGQCZFctqnaCwqJZV28bXKeNzIGs
P0s1Oahe3hXCjTrhkFbHqjyVqB4T4MHk0r7akhD8E03a5O+KAK1mDO8U9j5Wjkvqs0qyD/bJuX6O
dq6P5gHAXp4aeX5PHAAd6sFcMAnXK/6XFHv7nZHQqQtd4a9II2iS08Syyplj8YIxEndmF0XJ8efk
108FmrayZHR9ni5x2/xLP9+VsT3uoFxOXqtFZd7cCMqFN9fVuRM386fG01cq2wAvYFBHvIdY7xwj
akwinn5mOoyBla5M84LDh+phcmy/BV9srKmBNiDBgz4JsJW32eY1/6g5F1b5lwWEJGFubJfzR+zr
cvK35MeMGvoACajAVy1YfBS3zD9I5iRz9XDyAvn2nUZsq1kJhXPrdp7LWTEo0KHfUiXrkqNWUU5s
cjLSUYlhthF5q8+fKc7nGYzCoqjyz0soW4aTDyibFw4rVy3qy6Z7YRXXn+QMSGuOBN9YInbs7+x7
jAtWSGUM1y3nFC1TFVYYRmMA2lRKqi2lrV/XplPZ1vDDNDoNiLRJboTHsxogq5RQ0vJ6f91ZGsL2
zYQXpnnid/WAba+h+V12rkYaC5j4mTBjeIVJcTV/AtPB/6e/2Am0YR9WY3OhdJAjB/23uwpHnhj6
b5yezKEDnai1a2vuWGb2hoM0dt4VKMasNFxq22ZsB13F5RobfIYN3LxIA2ySwNM2hLjgMtbTe2nG
rKe7ZseyACCnEp5so2nBKBXUaMohIrqvFX0NzTCKll+jYLlPypjGR9JgQL6EUEnnt2os+m8cLwrK
uZNBXI2+9FF+2pSIIZPqtO9cWOZRsif85F6zP2IjZ0Kqm/l1LbjGNHntOfTv19ZQurVmobhi9F01
iNnP1PdOSZ8fZHICietEbxfKG0yBVmwQ6+qs9vqAtA4s8EJ+05052FZ/DtY017Z4QmCV1vFmY7B3
ifXcLRW/Bi6f7mwp/0B0SjK2BEcnHJ9ozfWLX6JeB/oYSrMTN9NLdZqKEeINjuDDmATvBKuA4Bug
JYKxc9O3Fvcq+v6npTR9yoUJMSeX198Ef8cMcCRcHbHUHcLH4adJrpG2AYJLeqiKI18ZEpT/JBiL
zL3OaRAKStYUnjB8564CQtZXr5Soz/Kdx6V9B8Dg7vaLACiyOvvzI2cQ6HochmIHYyqlP5aFPF74
qhpdMSsIitBJQvlHmJDjw44TaVkHt7LbTk6zip5FgFn6sXgiYZ8vhr1XOjTg08ofqzTtR+Zl76Km
sYDDw5ORGRlZWZVhyuHKeWtyU6rAHStpCskHECUNe/+gIKgTXtqttv7ofsduyj6fjqJU9wBAij+2
xREqbYlUZJ70OQWKfAcFtsHwsaWPE4r5N1F0YPnBAyKuaV2i+OF3lKw8RLFRfJdL6FjcA0WvxI+k
0TzJoJ+Ickm+T0zv8otaRqYTJRnVREGEqiP59f9uqX7G9diO5VkZxYnwNkFTTMwT0+DRIY5r5tKZ
dunEHfBvoPRmueyFM5Rd1x4YjhUbhl1uPatbawhcZji/cOyxLnaJYj+HZOl8Jr2n3WkN4Vkt/gzC
fHrwfW233++5WfMa4zzHQzi6Dm0+DwsKObenTF+6DEZ5PCklwGrDPMNuiis4f9HiRjHN8LWpkLVy
NRaPeSO2UI1k4gFlFAL8YJHVsFgytyubJ43t2Sm+PXrU48fFlHTpGnJ+K/G6Q+ekkWoM+HmMnjKg
UvQ9l24re8iEKlOwXpBiAYzEk86S6wJA/K6JQu12ZwWDU10g6WmhimYY86DfPB1Plh++xNw2uSkS
rBV9q4CXtHDt+dD9qk6KStmJ4mYgqT9Amm/rg19p/X32SvdjwiCfdQsCOzUu2/FYbrPbweGdxTVV
h4ebUkHR6gCK6mDbI0EY3/Z+B5j/YG2Uu1GK8kYMN2BmeMEQfjm4DSxqjwg2+ssK6Gk+R5HGYTQJ
1IBrOTZ4ACksrIOjMr9vOqL683EmqnzVYCkNOm+ekeFRsVXC/gLxNu3iP32FJNDE4i6bgQZ2yP6k
6Khff/nluqmidx/6CKwRegCY1/82WEYcs4ZSJHfH8sEgUOxhvWjr3VtKE/i99ub3xb890tu56Qvv
4vXmIu09ov0xcU5j4RaBPZ0JSl3fuJVu2c5GVvrTcIf6E/MhwyHQOVC5SgrLtfdczrt6B9mYWVCU
dvM1L2D2qrTf67Lf7ZPwFPff+UKnALZYmYhX1Qp5m+KaUSCk0lrk6f7ET599rrPWr0S46v96NcgD
4G/CTuzmtLjfUeLbMExmXCFh7Nugh7K70Sf640cPEtEAsOyqoXWCFhmxZTk6KGENAA05v17CI6LT
B2nmOOVFbnzAsJ6Mopx7HFZqzG4++BF1ubXVx74RvmgpRpCtES8OOIWWS8mqhO14AfGtLDk9czCK
lvdASg0g1Yw2M7xZlNNtdPrWm/m13qq0vvrDiby6GHfGVPh7isLPxO6ws5RONdbu1i807pwCyh6Z
0SBnS+9LhtIXepnM+nV6LPRENPeJS8Necah8+P9BtVgmD2JOriTM9LUSzQMTZ+c2Nk6ILhF3gk33
VH6mCaCpnXlKiM8fte8mSLgqxFOEy6FQBXuMvsmK0pjgPMERGq4lxk6W/rd4CnZ1xkTVz6bScfcx
skWEqIRwj7Z9wSKSiH1jhF1XaHfT1ZUHg9jG5qxuSdwppxHjHChBcjdez9UAvUV0T01spugAjpsH
cukKtinaZTIhV103oC7BA5o3dsfYWkEAmZ5QKTGQFIFetVrM8N5i8rrWtRsHhenEqJO1hIF53VQ8
eDb/p6RmpCGK362YZk+fBTY32vx4qurXfxMvUbY70aMjfasP8SgRLghdBa7qMVJkHjnVRkpDqjiH
uXpiK3GMmA66RBbWEb9BxhTK3+NNkwxgn6GuVzTy+Oy8X5pcFQ1zjZyTsGHdXfhsZibwjujT7iwt
mg1cEAU0W2Ed5dHwmS8qc/wE6mG5zoIJZM8MdFjNOO7x0VTRpZyCxzH+VT1XNgU+U0nIyVr/X6qN
+IYEZQANCUyIKMkB+EMPKJOHm8Ri1A0BzkQRMCgs0Mv+Z953MBcaQRIgU+UdURmR0SRdLdP2sEP2
2Bw8GKbhY7KTm/WKZSGiSwVpu1a8dHPVEa7Yo8DsY3V/IAeZoBp3/MV8IfByI1dilLCb67+xDZ/D
JUupMP9dlaj3XL+REgE9TJSSUwqSc3aCLGE0FbWiatCQT/TZ6TFUYPJNnYHvGpSTcfFmj39W92Pf
KxjPL1/jktTXA5OcwpqR2bOqW3e+8VnhMqffmBZCG21BcpYAlV2nBr7rOIpqU+UnCnQvweDlTfj5
tnYr+taOqZO+OXLnhOgBTHPsqQkoofNG8WP3tkt/5xxvdN0yQffLMyx0m1XintQMMMGVcwgGnrWJ
mZPJlQ0OI1FQEnRuFFEcziZf9XD2LA60NJyBTxKYF4WLrDg+toI1yjC9oZP4Sfv4sDcfc6iNPEys
GIju6vrToROURISodifuIpYlUkTd3DSi+VGdSVzGHeaaUuQed6r1ZPHxpWJsTxV/q99Hu50/DNfI
ToZ1kl5EJke2ywzahL2pGglCY3zEoD3J+PgLSLSciatTY8uGYiOvgaohrGcnZxO0KpYW6FJlIZhb
GEr1a+2dT8rY6u4yrPU+WswYjjN4/MflYwK/diPmZp0xnxM6RsdVQzdHlavJQxtx/NFrHB+laj0W
r8FaPSb8hjVTmUEBYn0ffS7EXSJMcOj/8sSLFtjEQvwR2jN7wHqYm7rcPX186CbAja+ucWRo6OMH
5s33oEpezoNlJmzUOzIXgayKOl+PV6yKZiHmtenz6gRPunEBXQR8tcUw3zW+bFnt7upK91anntuc
THXqGLVG8NcoV4msVOeFgjEcU71PkhfBUCY+Oz/RC8/QoqwVdMq/8V176F47O97jDvdCyxsjz2dk
iXVpN1K/Rjl5X4q/+1jkU/hlCy3EOZoYVdCWNoxuRvBBsxfBUymUfykGHXq8rSe/73oVm37xea6x
XDbhuDiJl99xhHZkFNeC2LNpL/TaX/p/eAT4MD2o8yN3uecmGgz5wJGcgZMEf6lKBoZIr39SjgCx
vCAUoH6fIVHPJvHQnW9LZ59clxPDWk09HBn3KJHRwrVd1oJeaQWHTm9Unf0AxgyW0I7FA4PITA3s
+VuAEPjYB8eOT43u4P8raS2SDeHgKcqAgO5yNrAweZhP8kGNpoGwTFVc6/Pt4Fid3pETWaK7qGnS
A4uwte0KbX0jt/5EwaOCsYBeWkd75aV/dHUT3611Lw8Ozp4251NGgwITU7LtLi7uBih7enELtofK
dD4rycx05E0rx/Hwj5eDeYzm+iITtBS7Eyf1jCW5regri3JIFy0VSm+IeGsNyVmyc1bzIeg/yoYD
I6LYxjTN8DuhqUFugANwTviB4inevcjSu+rKl0tchWSxsuv0P6GnqaMfsjqg9qggiHZlwu2t3CEw
bVTkM+w+ZzWO0JKnPoPu0eepddz1qOLv5PbaDW+UoHtmVqQxpdxT37yAkAWaKPXkRZ/4g3GgmZSn
g82vQWx8HYui6e6sk4i0NZBJvVgOn8tacuOVwZNZM4D3uMns15S0SWwH/NmcHupoK/XKGii5KJ0x
okDtko9xuBQ63Y7eFV36X3sy2UecsJMuyFCZwnS8GVd0T9Grx2VN0YJm6A9Fa/v4TQBRhCyFo6ex
9qtXfE96dUrS3N+GqOBBp9vJt1F4U1DHxa7YzLjoTRuMZKAWjjvW8V4++jpqO8+aRmxW3cyV5h0f
IkwhWwgfRSH8ybbP9+hpU/Jmkj21U/fJlIiuB9ChMwVMzX2urPMCho1czy9aMQ6FM899V3zJeyiy
Eq+S7qRIql3N+cO/79GIklOjQ1jp/kVRA7iapHyfjTjq6NnfKQ/3jN0FPkxq29+ysiiht74aCdI/
0oSsfouunO0YTThcTOaG9Serl2vKoXBDQ7JcWDUZIhcsvLgUcUOagId/MRvifKl8putXJ62kVAHo
8RqlCf/NKFakxg6Q8uMOp0k/hwBsCrj0PBn6ETB84bT4MCVGERsmMPcdNpnbBPjaVCJrBwIaqDjH
WYjgSKvwRdoAc8sBg99tx3d7Orav0FV8MD02EePw5KnmMp+EGFAtW8PI7fpyB/sh9uEHChFVspro
E5GCh3PlXL6R59JJFYdw6mDyAiXx8bPIo8i0Jy69P9oBrJjuQZnrrs+2bvX2i7+zCLbjhogBmZO8
BB4//0cEVt48xIHFjrlnfVXDrVfflxaiJ9aWoxy3VQbr7EwYwZdXmeOSy7FiLQz3igB2M1SmOrCi
m2+jH3QNINXc5//JProkTg3x/c4VldGd6ePrcRsmEYpOSLpwqcoyCz1kCg+g2WwiXlFSjkbjuRvx
dG47gIafTmqzol45Ygckb60BI7hnoqVwDgFn6dd+/o4qiGMPJPR+i0/VsVfzhhwffsqm2z6wWcyw
32BtmEDuRZroT1AAvWqT4y9qSr3DFr/bTqWozVcISoMHODPY4StNzoAjlqhG8PwgOxnqJFeiNPyg
7y3D5+Pc1caG2+fdpddkw8Sun83ukUh8aidXQxt/WGFljMKouXDcyHoN+Lbqxgwbk4HRg/BQCj+7
SFC3XlLpdpw/qfLQ++2JtY6FwsoC19H9jbXKOel4qq6tBchOLP0fZ5VjCBWKX5kR5NkUrVdpGY9H
4DPpON39hZcjOWo7MnbVTGx5EG8m94ApgMZa77p0yn6DD/OrpnAHYO0MKsvV4RO6Vbv5qhWJIMEc
c52KSZ0224n40yCfOwH1eU+tv6vVNLA17x/7TzM04IQ+0XYNIxRM94RdOLxW21+Gt6CoOsmWrkxv
07mVD7g08hi2tbMhYA/cxbevNZC5Y8A/HMm7Uh483uFhBIKEmrf7t3QDVpPKDEZ/ujcYdXUBtqat
XhHIVfUUfG4Eb92DJTWCMfUTl4AnL5ltceigFdnh1mzjF3haa2zUmyrFdeADKl0Eew3j1namwj+C
SNECJGeWTeYe1lA6LzEZHj2qOzu/J0DxEgVg/LvlMGAuZCOpAblXZIQl239G1jiAmRLghBKRP9jA
b3U/Wlw6yVMy/2Kwpgqr51nTDnA5bnNmHvcMQTQrawAF2ongniweng+tjtmSq6T9+frnIGco9xmf
L68WCrNMYwY2oINlAJIysCv0jpvgxZIO3nsbPJ5jUyX/hGg8jTOU3lWHWX/MBHBT52zdFHAU9CkS
3ZwO9bUGNXeoMU+m84fIAIQHLA4h65iP+zYKOwo9zCw6e2qDWmQc3aifxFSp35B2qRMUC2qsrvN8
kHuEIfYqfTbkHXxYHlcb/dAsLfSBzNVMimcSyW9eHrfmw/QD0Xh8vzMzDwkKYr+E8Q9g+Peej0W1
gj0uebjKhKRgnyN7o1Dhx4Zt6dW1NeFBD/4Ls3RQcj2KZR3DMpOgTEQwbnAPSpe4rBWxoI6gQGBB
HjkHhWSYdZW1Raa19M05NtZWq0uCBVxnkV76WGC2Iff9hPXP2oss+q4hDonadIF3TwZFlmubk4p0
BR0Dq+yPWbVcZLC9Bg0lK4BCy1H3GDJsY8hWEiipOMo23WFNdRZXscRmCoW/4bVGvvsgPlU18Uh3
ebXeOVmAY97uUKh4MciOvsH/6jKB3oaxWNQ7LN/YjP5CzRfgA9IHFPGmx9z79VNfnFRzjgeE9FmH
+nQOYw2UhqfrWgK7rGA/5mjHTtMgXNPMJOFOoO+aAVcH6zxq9Al9/8tD5CHh1pWYOMPMwGTzeDZZ
HPIQzlrjlzpMONiPsck+zpd8kYI2JSTNACyui0/cGCJLv3ZqWf38htD+gICl9UUrFfolOybIhEX3
/N642fuutaHZrFGL026VwKXK7Zi7iUwrPejPUvE4VggIWrIXeZNZHgLrBRygxuCPDLPmhi97Qfxy
mjpyxCj1yuXUcUmdZs0dt/Eqc1Jm+ZchjWgXGSYuaqxCsF6Q9+xFsyF9kYPCfqs6yCOlwG6tJ3ou
qYOjsHFLf0MjSHmM5EC0YrxWqWfnee+okw97WRSIl+mu1p/k7K+taHRVg4PrEkCqp6s0hJxg8thV
U49eE97GsfVZo4WQoMKhGdOePeEE+xBvwnvoStS/nFKVAYf06hTB8Rjxfx7aym9ABw4rrEdNOKf2
AfSPA9RR0tLUaTZ+w7PQjVp+cRAF8iLBS9EalggIiFrJL8TX5qY7qS79bwO29uqcksVm7Mb7iYea
gyZ9vqk9NsbjdWwsGZeHQsSOOflhLq97qWRJgcUmSGpElhnx+4MWVW8G5vE6e41E5xNHuh3XQoX9
ue5cnPrJ03ZO9s+WfpNjLa9A+RFClx3mnb5OcuntkJwZLuZIsRZGhxmqAAboaNMH78dRt7jyT/pF
oI+W1hh0O2XrD7jzVj3Pq22DMIDIbGpwfSlHRYr4Y30e5GMfhhDQ8ToR4i40b+DgBXdfsNKT0WC/
xBr/fXd7UemJiFm2UF3bxK7Yjn71Up8VmEjvygRovfrcNy66hpUoB0TGcy0PnDgkhHjTklSpWWE8
/mKTwxhA2hTwXCKV+JQcE99aYEeSnb3jA/3jitpveADEwbvg1YMAsBfxJRKDWdLtq2hvakraxKiM
uWT6Hcf4m6QrGDPPkTLB02B+yfvVce/EMtGnCjdJWkRvwX+/qNGLDg9Z762ocL2FOc99Mfwy+zvH
MCjwSnc+RbVbvYBTnVOvLxEnboHF/VN6f26E3zeIK2RMhuqZdTMKOS4HRnCGLBB2KY4X/0QdedWH
T0LgB5NOSh+sl3cPuqPbTqSYDxSDwoj0YjmjNaFrUzKvecEtuc4vp4oiNiPhkszP1rpvMdqWBZDf
59O+hvbYhq4eZinEdcRW0A5lotFb6fD9Ui1rCHXQf0Oi3bEKSub+lVjM6vcC6GLg9DBs3heCtaNk
VSUImukzbmJAQNe0GEANtalhLwreCXVhj+yIa6KhJywRRGDW8R3lfv/SyVcOj1yYg0K0JKSu63i4
ce2fVQMcdkimZHWAPCagjeNEvjO/OYjIOwTIO//XEQbdH05o1q0ebfN4GAr+LWmzJCEK7Lcu25wr
pFc2JMSokPyYN7yVdhtLq7N/9Gf1kd4gsRciBgdHHoRs3mo6gNDctSvtz07ADz/sextmYswnydjN
784UInCc5merIqSVT/Xfr84VjeQ9VDVO+RoYJCtoL7gdUksQCQCWEhYucJmLe2gbsMox92rtEvJ4
jMyM6JLBDugYLvboZLzpp5Y9QCKh421qkTVHrFbyz0BabWLwAD4T46VdXopL2Ughq2pmdWriCyet
Tt0NbmjeNF+ajMhmMckm4Aqbphcq4sNDExWTedmogadnK16IUnfj9tMP5P/1h8i2J9W8snbM7VME
TW23oYJfDuTyYVgmm7uPFkkeLZY1w9eIhYSRu3CaQOEKM/aSu8dDZVjJzlRrArkK+4DnW+vakWYV
d0yTCe0NvCNZaN2ymrH7cR1vZ/AbdgETNZNa4tB3CfMEoPtZoWYtqe5x9G/w0w/DTE0ToAIzf/d0
hYQ0w+VoB6qMZDhNYeqdr+2lyxbFxhdyLvbx6RW3NCRG6YZmOkANbeCVFCMdOJHrtiR4q0b/yMbC
Rwuj9OdwCFX9DtGSJJw0BG19mMnQ8ib8PUp5nS559PocgGmwerBLFWJZdlvBf90dwE7iRZojZNlJ
YNkIojAC0LJra8geZagMv/CG1hE0yuOeEi1CfFW2cEtt3axJpqv+o8q3ip16Zig5x4lwFxlqzFqq
pFTz8R5dGlk8FZVF0eP7oWD5wxJwbD+XLdQsdI4DXVFA4IvboHbIJ0LrqUgcSc/99oMvd86ud4jc
wB4Z0zfy8HfM54dHzf1Zo8ORYjJSl0T9Pq/UjJuAupJzponzSkvF1V/AfExHEpderbkcHPuyFeoF
z2IJVypXpbBkmR61B7WS7jZ3es0HhwMNOYaamuvmHWLhaEBv+lbztE5maG4n8/j5pLAcQqP9If40
8IYJNumrtz+tU/VTQyQA//HhTgd4NnGxy/YRPqcFsXynhmlRciKtZB1R9MPXosxVuSD5tkuFLtX8
tMjJV2LKMzZgE1Xv9uYTP5/VDHeF4EudtefyQVjfWzCgeXxPq3p7HzCdSpIXYzpLtS7yg4IgdDpX
MWnx3FY85KrZEwkNK/P8An+ZYaZh0Onn2snpfE+UgZ7D+FkXDoTrUiP4ljDccIXNfacIQzYjkqCl
zaRFz/5eQKwYLZ8lGJwXjCv15PMsJuZ0FaFiGBJLO9Yb7SO6ss5KLxq4NiSa8AhCbmZ2hm2LiPs3
dTDjKOO9J1EINyeICQ1xe7jf1rV18ydyXppa2AFNMhPQF3wIC5bipriAEUwJgiAK6AIFUfG4lOmH
HVMbHVtLno2NQHSsWkBwmJVVoixL6HQrAhOkS9Qq+zge6U9AnzODSHVfKiJMRPPwTTwFvYcBcsQs
QTv5aBuOsjbtbV4VwCsx8C9lfRCXONUqoZD4QntD3bh+bxPS+8bdZaVQuJRkB5Z72/ub3LaKhCDa
6GyzUfEtyp10vps+REOdg9vFeP2CItiCHWEmKTZ2MgJlvyXDYkRIIsGgbfe5MxsPe+inHVIQg6cl
w4urp+2UbDohLypBNf8yvcxhfptSCMqYRkXCTEyQSJj6BBXJ5WXYS2REdTCkaedPb0uLUVVZ6p1f
RBHo3jdV4RqdDvT+K3wzXeODr3AXrRDB+cCjNm8cIC8JpY9K3cQvsa+xFSRag1MOoInuIIjeM/3M
eR9YLF/iLoTIccmkd45CJJJCZrXUIo0a/pR2Epws5U/iF8EFiSXIrxnGe+DyqIMsa2rXCACCSvc5
mmZ4CPQWGG4dbMNvFudU5SMPpTA0VnegpYFS5GXWpRdSCxDAMIG4kXCB93v1NGWVO3qYGHJgllhi
eYZd/GnbMTare/vI6mbYpLqDuBR4LojnlvGe5fKpdSRT01LFcWrenUFb0+E/jjnPgTFLGe30JFgI
OlTQVCQMIvytSXuKP4orHEozsV9Xa4NsmgDVpc8ps/0+lONUisLh1Y56JwWCRo7zmEv1JooeXm/h
aCN+7zN8afzGAn6dbGeBuZFwIRKmTny//9hzhCTcXPUIcZeti4SEm7DK3fsrrs6kSqMqCkt5Etn7
Y+9tJMopbLEHDw+Q+bfWIW1hfrVNf2AoIecYyhxphJA/oiZ/7JqnC6gq1BWzL5olhywPQUXaXWyy
RgRA9fss4QqOdFBf+zcjRVguobPMLEM2JWqbqMnDKSHGpi+CzO3+Dc82DyVHUOWi1mR1Ak35D1sf
F+vXI2eY0q2LSy7I+Xj7YhnxY8Bm0LRWiNG7JmVDo+UvHoNw7yAQNG7xsGsKQdSM1JY0W3oSw6Q3
4cFw2fOnp6F3cx1JNNXo1RecJ63wF6fAd2sHbB5BPqBFXukWeKcW0mYrbanVxIZBziG1iwvddpDL
DGnWC5a3y2OPDww6GtaBfpx9a3eM31XL+iwGfBChUJU4/OuZUgnJcp4lbZScgzFqMWxnUxUqnJdK
uLwjkp/OM+gOIlPnoVDzaWaHQNKvasQ52UZIKg4eFlvVmw8IYYJNEKi3UW9nWhplbh2riOGZ7PJg
B5VJMiWkA3f3CnkrYDZk9FejPB/UCJiFXXvik3OunlmnHhM9gEVkgtpYolkDaroUZ84JNtdEUUR4
Y01RRF5L6+BOtdLCHluEx3tKvqjPXG/MCrpV6N+vfJC+6tirOrzpcxS9EXVGQU3zNr+sZiL3uVSP
uQmnAJCqIqPlfEBgkNBqAnAxRxodslW6ALm1YqK9nbNOK0/Xy9BRYRm6jCN8wbCpzp1SSFB6l7pO
78uDMpbSaE6jCRnhDLMtdbMWQQbT232FwiD9ysCrn/RWo+Ce/2bIBKMfH8pRz+vhAtof7/dYa+JI
g+zdJeYjtDK4HTLCHiSjsdemM9bwu1tjdxapJ+1rn2e/5VajXkQc6YHie34QhYNI6Pw7CMkOJI66
6knC0tOdmD488aUPiFYCsygEgWp59VeQLQJumFvMDmdKtBhbS0m6goLxDwi3aA27RfXwquOqldEH
SzUML13gWavuJV6vTnDQKpBvuyMt2/HqXL5+e3QmmSUrB8UrW2mSZ0ecNEpd+7NfiCS1X8gtZGwa
4cuVe0w/wD28SQVHthtKfDhI5X4mGeoTef5BMharcenEIMAI8wh1GWPOhuanDZf9jFsM3PworK5n
3bUnuNhySIwTTI3CcVENW+wDKq5mxvgV3EPS0mwKP0glib3wOUO50H0/IUSR0rEzx3i3jY8zLbKa
IgFxOVJ48S8abhxGe8zSLQz7TvSAPna7qP4PuBdr5mKGUmknsexXwY6Xa5POzLRSfC9j4eWCwRCK
cZYjHChjXi3kWrCoPlSsmL6NOLcSYr91yZyM6DjvCm8Pe/K9ndFxlfIi1Li0JkNxkvB6EfYxsRTY
WOTb8xHIc3sBg8IBYtgYlPXMDPRcf3WjK50LY/n+qgrhdSZU9/1l1oPsr7XWKbgQJFMPa6sKS75M
1Lv8HFVdWauhY2oIlpAHIBqjDk5sw7sXFR8S+vhdnDb5aW8RofWGhbvaPeOXGP8hvXjbVpgDboFO
TnDdHyzUM4OK2lT2Qj9GozLJb1/2LOWQfzcNqKFGoRuOhg4QgEZIDcsngv+Y0+OJe63euKkPbR+N
m7omXDd/BFKijw/0MdU8DsKPznLjHxCxJU7MY2Tk9zuN0BXVgYpAg0MA+4/HTwb1WxA10grZM6+U
aDLIQyU1GvxN32RrjZdNPciVeFVRqwjLc0zv/cCLTInsIH6JwRv6P9yzQpOwOa6MDJJ2fcG7Gpqt
8TlTuidVL3CYM4KGLmHf5RMw9eyjSJb6afMrjNNDuUGV1UkI7eN4C/H4Tc9Leaan6vGTndty1K7m
F/aNq0yndZ0JthiPtWhr5AMp3VWhRsT+V9tfhHN6ra/Xfa0DMmpb8u7SmIQi3mbaswu3TAkm5x8P
svCoxR9ZQUOp3TYqpektMPQI1aAJysX+eTrxfe3Q8Jb33aDVJynTTBUUazEkV/KRGJRnn6j7JZgr
57f9Jih+/lhKYD/bxRrE9AQUxk7GQK5UHqjClW4Id1CeBscAPHjCIMeA7Xipt8vSP3xspPcgGv1J
a3ePinNaEAfGx9//XbygtjyssTLfh6iN84tU6I19cC8rhnPNY6KajL9LwRMeS5vuTcqXN5DdImlF
fibQK9OFSj7D5ZZEtpF10L+AI7vv4cawpTuIpZk/MH9v9wPIpxvdGqrS9Ngkb+fpgL/3ERkx5LFX
NCZ6HiQ3Kf2mtZAk2KxuHA16kTfmU3xv0bHwyJ/BsaUSFoCNG2YC9q548dUb5YICa4nQE7D+mSyQ
HZ6hz/O7ceKdARpCUKqeqLWGTEID8AKBRgN6Ikh0nUOlslpw5YaFgzKLAmLBxBLHOelYSmyWjmR3
U09sFuWgWrfKtgxE6jeu66ToHSZO6nLogA/J7e3BAw/hYcko1UyvcHsDsIbJXT9VT0lAyotkArCv
A9RYgALI2XDPQQz86jKFbsM/Sms/4EIAwaouldMM3qvADUjJcZIXH5Gw4lbftrdLjxRj3VxTrd6s
kC4xmpG3QBqEvLh/wK3x4mq1BvBh5JMF1OP1FNl9MfjPnibFvZtYcPxbqlKVIRSVWyPNOtkWOCRR
NRLslMgvttDPVp1hOd0k2tIq4KgcodCL8e51tk1vR+4EP4XrR1PXpFnYH5TRp/ZaYw5iFFpZZADl
FkQA95RLMtzZSyphrijDBeyB6GvQGFee320e1b8Lw8R0BPCEFrcoHMF7kAWuBpyllIYX+NIgKRLU
EamtA6EbJCIMHSv2D6tfNX1iZ5cFf/gkc9+x0VQAhuGqtFE7CPOCrmksGvJN7Fbjk+EZTyF+mZ9B
RaYXsNUQmknWOqJgVYUB1ZoFyO6cdDe869u6JF3vw2RP/hXsX6TaSpZPsuNL7XghwbM3Bs7DuPih
8DmsyXE1OAO8/H4Sns49vHJgM+poiK1HaulPd6wKAYRUn5Pw1e53wCxZfgIxG5hh+SMGR8Gx9bdY
z1sf83bTdnssmzN0j8EGIUny5Rx4201YtZcemg7MsOuOXWmIceKlgloNB0iW5tg/z1IzbskNjXNl
xzk25ZUKEG1SvYUwp2rFtka4TDWKGw/2Zi65RYXTGy3GxMmijfNjeiJLxw2Z4e8bWNkGIDjOvCAQ
WDhgXniS+q8Tnj+JgyD3j5zGkYyLm6e4lNkCMQrQjrGEzxSoC/ZyrISe9ZWhLX5XbVapnEU0Ht4K
H2B691Hha8FofhDWy3+RI70gUlLpM+eTppSl8YA3/n+unOcFHKkijTHunZccen3mDr67Ean9lBGH
xiBAI2M44ZcU5TKqpI6Vz+uthzNAd6f5Fui4b2BV/zezs0xKiveueAV1U7c3BXE49VyNqN65flab
zaGao/ADXnG95AMIPrXpZbJR1A7v9n/HvQrXm9hmdA3dtckxeCus2cw+qQAzSjObbaTPU2f9gSYF
q5XB2QbQvJg8AWgcIUwgIialjGb0E04ORTPXk4TZPTDIFLGbiiytxGJ1KQwe46YPKm7+wJT6JXEQ
PzBTYW7W8JcS0JwvEdDzKZDz3VsyzMbJWyeRP9HZVz+fh9UKd36/H39W6YP7rgMg/0G7L6S44X/T
9hMwdTukF07s7euXIbI+RoWJI4qApSA0OLKINmDz1vS8tvFRNaaj4mevMN5t7QhwasW7jdIT6suP
C8y+Q76iDbqlSsKd3UI3FeZZjHFr9ISSBHUO1+3UjIv8gb9JK9YtDJPyAUty+1F2PxNi2h09RtQj
q/xvQ2tS1+RGfP366RYu2m1ngldK8LD8FhrP4Lj8VbJIKP3fGIFa4J/vFiXmehDJuO/fIMPrH3GT
2+ZTiScdB9ogWK6eV5EBssTRS5H40p0TY8gbyDquOHrB/6G2hOYFVCwbI+ZztPaTMdv7dICbP1rN
774jEkhA8PymVgLF6P8YKk5TIHuRAJaZOdOoJkGh1sB0KMWblU6s38LGaoUDm1anl+CaQSM9VrIy
DNfUu5Az80j2oTPdag1YwKFc64x/WEmddZR+Jyeykh+lGLA7ZiTRM9qvanu5MuINcKdUCehJiwWb
cml1BGNN6pa8MzWHJN9mYlWNtbsQDGyu1xrDPX9ii7lXF5u12hURcus8uX2qQqiNzaEepYSeWI1x
FoVQWUSjjMvhBxx5LbVg6539Q/bRgjTL96FQZozAdNimfkjdSmH3Mk8s7HXTidVmPuhwAwQxzcZR
dWavGIWi9BLFCEc5CZYTsaWUm+pSQRGByhwTEhm5ZZ3+1fcfGJmku9ZKOjcy75AowILgjdUXTbu+
e408Mi6oH/IFXroSsHA+cbA+UiGWQ80pm+CBnQYbQl/5ZbfhOFyTQ62hvT8nKiYULsXu6t7FCovN
7A0dwN0yWEEPj3G+VhXbr05535t6MkJRMEMcUhIyoAQLEM6hZ0Hhc0CzYtksf5Zh6Xi8jTehjttt
nXvP3/3TvKxm1huEr0pqOs8J3Tis93mLukIMJRmuvSGIIHWvZwFqGOYnCGOqJTZnPRcgCpJ/mDIr
/Nw+PhogHGWSzd3x1I+eZWC/ODqEhGa5lxq9o+YzRuOm4hT+9Lr4yj6G+ipUPli69t8SW3FvmX8Q
Qsqy/7PA5oKJZCPxE4CbNZJe+f6F6xUCsOutPFnX4KfFOX04DyP07jtv9vZa2HEDv6kAT+6sk0Kb
3eUC/jxucKeMFCoC2knMuDp+HWSHUcYWH0H38O/tQeLNpyTI/adJc3qwo6xgzCm4rmUjwyCCmSa0
399wsJ0vPacpdnLdoYPMDP6J5wiGFnrmw6w4mTkx/YPoJLSrNVzBOha+jJD3YSYIN5xBqQd5ym9r
7MaTgY4H5vOX9Y7RBgcU51tjKRyKyREUanmJdc3v642NagS06U3UbVVBnOkDc0D1ZPFNRcp9Aqoa
1tZhmcS4miY+mK85jcc+9njUeU9M8ZvTeMhhDY1zc7TtZbIOpQ4WwyKQ+w3+9YOL9GTS6Q/5aDLd
R0C3JJr1z/ycX/db90n+d9IkGqteQkXkUWkgGbSn3/fa9eLk+D1X2E+zkWIxgYGPZMqiZF8c8XaM
BIhDti/l5A3XK81i4BECDaCSLkZa1wxwh+ohKbyEQ+0cW4wZRb8oJQ7zN9Muv69WuoN7FqjxHBsH
W27i0+xujRGnqDAbZLe5ucOExUDBdPAJc6ed/8ETIWY2LmM3OOb5dFInHpe/flDB2qeyoQp+rSkk
UJSfPqAdsVP0CBxQMq9EmecNPKf/aGGrmm75G/JMYOpKYA5vs+8h1/lOM2GRtUzWzjoSwTt4Q/Wh
nZ8IvVCayeXuAPcQwt456Yos3qt88v5TralpFzbZNKSQASGhWjHKJTSO1662Zw1865hS1LVEa3uf
inlCLObCz33XUaW40elbIJ6tVAsyTnCmKQRwP2CWD43YNRWJo75Q0WbIfbEY8syJ04AdkYBJdeOS
0Hfa/wgF9PIEmW+CH+Dr72SMyj215Sg5wwavlQM9p3GV5hPYWlp2jaY6YEOQSLbNGR7UVCKree9x
QcTm/t4goKiXrrlfvJsLr65qt8252SPOap4PLXNhSl4TPSdjgafmHSY7xBKmVFhrpfWd4Z84v18l
sF94lo0NBXw7FkYwzTDrfuPAde4dNO6/DjS7c2we/bT7L9H1h/hBti3sC6QrKwgXhsjL0MSEPfdP
YMGXV5dQMM3ne28d7RjTiiDnLTv0Zd0bIpG909uSsmEoYBYh3GM3lCff+wJK8D9ARwVp7tVWXyD2
4SMkw8mha7t3gRNSoOyd+/wKA0DM7KtZ6XExp6VEM5xgAI6jYDBGI6OHsFmOhDyL6cIShOSc6TXo
DFPO6ab0FuL9b5JCKk9CeqQNItgP6g0obzjifYBQArtfnifhsP8KPL2RpITrK+Go+ApKHZqQUcD+
ErMpioCxMnSYS9Dpd6VBiR9vbjcP7UdpaKGIdTLiVwl6koKTsUl4s9BZJ80SxcXUw86stGVA7NFZ
jqxejO5goXbyaeL0LJImt7I04To/9eYPGzsS0thxaBTE2kjAslp4ZZCP4pXtLO8ypi3uLndqjfzw
bzv2nDC5qOUsms7jM7vQnH5xWIp3QG0OyJp/rbjlRcyBlTDL6oMp2RxB0KLiwNdy6gPt58VSPYpO
Y7xIx3QO1vnvjhwAokkag/ye6Ijn0YU/Zq1Ro12XVEwoVWDkydvs7OwaPKRUnODr+5Vs+/M4HZ3Q
G5lVbRO9l/qvkkc7yO+WH130SNbCcrYlFlUjlA0JxaAgAnKCe9VgM4gpT/cg7RXNvGFwfWsESu6p
sMYufjMB3EKnTlIe2+0KzGg2QuCOO2FaKn1ip92IclkxnHdJQeWtZqpDjK/S3pxkmSVm/K1HdyM4
+WY+jtzo4j1YNiGTob6ihJHRo75P8sqyx/ZcWRrCIs60bjQq8kARW/DE8Ruiq4G1kzoPU0BKkNEK
ke0tkVoeYHqUOMBsEoiJNH6GZV7oYHDU7HNaQq1O9s/bLBdbU7Sl9S4xbrEjqtia+3fWOABzusPi
HeK3HWXNBDKJ0iq+Bt2jM/5ibYAi4KhqevD4Qb8wZGSZamn8UxCXsfBfyf1FDxWTdRO5C5OKAhvb
oP/SHS14IF5wmwTakwavJS5S2tet9GGnM1khSNDPaaTD0RiecZ+lh62CX5jmpDBFH9YMphnTSYoe
KnezWPcYdi+D/NrojEhXlu+bRpP9khLQ/87xcv7+37P4o9sKgvISwCujsnvPhusXIXGl6GHvg7KY
27Ptf79ddSX2BUwza0KwqdEnlsTzwJzRf7x8j2hN8UVF7FTAChooFFVkgYJ6YJfcDm/bPwf95qoP
XlHI80k7te6vxO1c/mRJDZ1S64Mj2xDhUD5b7ug7mOjGXNSUczCF33ezWD87ZJO2bt/AByGfIGZq
9OvdDQrY8Oyx6uFnCK5TAiUCaRc4VIN+WKoqikOvdh2G50OkGxnZFjaI5SWEc4lpWtWL/d0sIBIi
BlYw+A2VO20tjEvDCbYkUalthpap5WYVdPebe4kmpd//N6iPJcOx1ahZtD+JtpBeQQAlWza7Q5Na
VbVwwFFE3LvwhVk6iiCBsfWUV0BBkY438NxKk/vf8Vs5o3Aip2OAC7W8LKVehztpj01vtz5u9Poq
7LVGy7PcWxtA5w8HP4uCGNxl8xaj8Uba9/oH2bBW05nCB09/sNJBexzvmqLRLsI+tKFnwLlG3zVe
Vyixy7G/hrir05KZJ+3czVjYFZOKdzxMvApNa8HQl3F5+hDYqWYLZmdERqJV65umYdRt2GUj+kXp
RXHt0YDHIA6vCvGPc3BuTw4pWc2wydPxQGyil38iMSYQVaWK9sc9CgoIDroGU97b3bHC0R8TSZCC
7I41KA2u155zYJyuj2r50Y2JEKicKpwwZyaCOO1W6Oxg8zH2Z7BJD0iLHmb6i1/z35cymgvAfWts
G2FxAXxGZp485yt94DV77DO9E39Bia5phJE7MmK8/y1PAL4eSZY+VJ/BtKix/14JkSYzWhooSzYf
gOnLFHdop1+ir0LVtjMCAj566MF9z0jhuYjfkDZ/JmvOpGF8Shy7oBv7VgptbljjFlV38tVB+4NG
2tsB8EpwO/VeYRZZsMQapa8JBrQAFagT8FGgQp+McCmIRezE1Ln5y1f/zLLXcJuC+Ix5rmGvKnIF
NNv3ReUmjYP59qEBNUQOfDnktymRh1WjFz/5g3fq1uDEBzg+L6LOIzynhi8HpN0RBYXVQgXgBFxh
raN2Mg0WscohQyV+woU2TtGoT2lQuVxzl5P30v/C/wzejSmuEYYWwn1w/8E+psX4gtlzNo4u32/Z
r9Tux5X8JxTwrhJx9ncRF4jBkxZgAnTgvirlGmuhrT0qLN8zEmw+/pSPzN1Bj8K4I1Npt09vBVQv
ILFmSNJaZiMgMwn/vT+SxY2JMZta8js9VFrV4b150TCe9YRQZXs8JWrgfjoqDU6ZfvAWVTmItd38
c+o+/tXWYA3C+HPbzNp0kR6g7CGTPpec2lhrP1juuj9YgA5FmZFD1UDnvBTUzHYvztRhpfbPlH+r
80OUhERJ2GCmMkHTxATBimNlQvUmQZMZEiDoRgnf4o3kZIo1Xw+QklL4nbJrtNo4/1odydDAipKn
xfs+FK0zun4C7ypGzl67qodb8CgYpufmkUrISBvV0wX1H0uANCFH7ydsq3MzSWY04aeQQaXTc88u
AeBqk4czo7/NAOgeq2OF7G+jZf/m57IdB3gvF7qQ+rapm8aDN2705g2aecexcJhl4mI2YDf9u4Zv
mevWQNTS+b33u0ZTgYA/v8SrY+OSCFlT1JiG2yp6+u01ondnYi0qK1WuwztaKtJcOQ5o16+hr6Ko
ught7l8LVa1AtH3Dwy9ckrk7ZNefeG8VvNzgOyTpYgQiZf5mKmhbndhKBciQHms0A61FJIoBgSmM
4YkKVvE0cEZQfuwj0o8Clkz80VwAcvDoT7D82uTc0xd9iKz+4ZbLEEvvClgEOP3SINx9ZtrAOdwN
u9gaj3KoaRPBsapDC73xZmaPdvhZH1THSYpe4fhq4KumxtbO+6N7dw4kIqiMGHdQ1uXWtKUa5zer
5GjBEluxh5pQDxT65/NqB9yb0xZJqXBQiax+7H0KePBJOOewbRUEpW0yLQi5xFTkG2pZU6vho5SQ
gj9mBt6Jp0PlYTmEdHmBHCVR2j+kIkzv3XDYkEpbCjbQEwwVoqEMVzsfNDjTdiXT5HWj3CvKdQhv
fTL5dpJhHaWZsKcezU82zYwJPgEeWmKbedjvkj39bANsC3eYT5UC9ZF5vnWIVMtWCNWA7dcp9D3K
zt4wENsCLiqvwYNW0/mOj0OjALFA1dL5LsKJjB6YTZaEImzscaokEPJ0EN1NkynTmO7gvxgTe7lS
nqllte8ZcO9KTM3Sjlzk1vW3QGj8J1qRJIKF+wl7vfwp+d4fzJTR9MrP45i/0vZHLjK71j5KMkde
fqAQwnIVBtUR7oyGSTjNMaCYAOzogI+Q1EHB6mkXDoGLPSUs6Ub+3445HnAtVMwdl08B5wADW0ZC
p3579Jvyj67PnPKz0sFQr4yad81b/w4LXlYk+8EZvJ27tw5UimtLJ7ZiKNgvNIg394BoXFOk+mqt
z6ijkE6nqQl8OEWN328pRSVODnGPlA5Jx4dPl8+7ABJxZ9FAO27kwAzNX1wTxvwgTvaipZA8OfGv
GSSRpi/pSWlouplq4sf2MPQxXjwkHemXRawybXwMUJOuYZc3zY4U9eUgDas3jhucDvRqOr/moMTE
dgMtsNPC3+Z3ltpzVLz0KgEDE9EvsjcDwaWdTb97dCq2DxAsBZH1a3cQOuntjiDqd+0Doqvvr9u7
Fl+nMVuGv0pA0wuAsLTsZpnaQUXC2HuOJEUZMTkRI0fQwS3sVVWswsx/KXpbJMjCWM5RzhAz/82o
ZCwUAlqROAi64Xe58rI6W3CEONdnm0gmKBBHaLcF0F+mHnWq/oIZWp3ChuA3QMimWUs+UhseG773
LyzR2+1WZfmEakYn9pbvtPRyzgQx9aePhYalp0pSej8cXl67oONqGpIXnzp6ZApEXD2/LRU5/0gc
ppJrJL4QDvvweTv2rvZtA1bzRuLi/CJ9cucVJ/R16Lfnw5Ge/f3H8DXS2B8fVqxwokpZrV38FJMg
CR6D2ub6Hfv0+7aMuub/Lr2fu54bXaMgWMliLCd2bDSJEXNdac9kypGIG7RN5bJ7NOaw/ZyHG6s3
SZ1ywuD5ABcHv23fCy07h2u9EwEgWB3gCRQjggASMW1ZekW70Ew0s6RVxG4ygNk2fpWOjLFEkqgU
u5/SZen3VO6yfgKo7a4ZLinLyb3OxGNRGzT3H4FjyMXaL2N3wEe+AEcJiZJ74cGHm16PxwMQrqGv
e1RAIYBIniu5NeraySWv6iy79mMiHXZpWxJSZvycaqZMkl49f54DHkm8hOfhhNnSwGB/JnYDXrM1
hMC+kgnwjw/JaRAv/FZz+3U1j9uxNxbXD4RY3ISLtOsXhsERcByE81qKNDtREyQH/Sw4/moh4WHj
NQNvXIJ5Gy4t46B0HHhKJD8pmUHZJ/5sarUrqKXQ2MBQmpiKoL6It+HXp5S90kj6YEUti9J2Wiea
ALrV+1XFPSojSPvdUgnS9DUjimiLU5Y31ft3fqFP3cq5V88fWJAkrx4UmMehNnPryDJHwn+U+de/
R+Hl9UKMEbgT9vLgPEtZmAx/XliUk40BQw3LmDC+zeyZxO5vJ2y8yHuN/8yYEVTmW9G4fjYLpq/i
FpLtVcXCNcrX6UmBoMapQ540QoYhe7FrWZ3MiKIzDHSMNOug8RD5cd/RgFgLsEtPZh7+bXH/DRl/
8OYayL0qgEom9Kt9uTcfFEIBdBlB7B2CCBUkVxVJkpqtXTdrPuOxnDapZXuoyg1diDID74dfTmjx
5+K/oflM1xrHZ6Zo7Kn0SWxq7ng9aKeJQNe4L6gdkFrFZ5O9HHvY7ouacUI6KHRFjZGJkJq6j021
Dyx7i4EFp9+BdQjCZ6wNFYRLLIPJY9XffhaIs8+YEmzCfGLpZO4TvyHw/3ktqE2GXccPvI1sVes3
iof4SY4J+pP8udvSVblW1cGo7+IiJsOcPNDRyqw8g/hFvLlDrp8FXvJdWL1ZfWcgAl/jbhVGj7En
9Q02lmB7gFcFayoIOPifksZiXRwSV3GV8UGaflW7sca4dMibRIfm3zzel1B0ZZ+Uy9GaZp2e3CtD
9zFSU51uPUmcmnmlHw537q8QFWHKz4vw7yhTEtvX4tmHgTxIZYvheft6E2N+A/lVZBRE5x58L/Pj
U/U8wg7BpvaAabCaCuN0o4IRnlWgQjBaNRWfo+HRUNqQCFQ6rAJjxPNXtVV69moblzWfEzG/kiCN
ES49IAnp8qJkMY0uy8DZC2MII+UYWDowUwGEeQaXl2jpPTNdY9OjeGNLaR/4aFoWxpQsSCQBFk1W
8P7uvIJC6KsQManmNrTFm7SxxszXdmdsmFXw/3kV4+9HJELHgUSaWWG0OcYqEjJpEU5Zz3Fj2h5Z
AKKKQWjAFKn2cNTojT54C2aQYiOPRgCp0+PnghleKkqxgcz9U5amlZSInWXBttGJ9tmyFrSSHtQj
2jzk3o84iI3behvOGvs2BK/a2OGVFceo7tKQLEshTi45hAq5O/yNuVRoR7+hhljJNcPNW/sdBH4/
EW55YZiG9KGx7NUc4ExoyJ1cv8SW9jAhnK1UK28AUAbamBpYJhDp6RgcuyjBk9KevK5HZOd4bK0s
giwWvGn8zPTnu+NSaOUCmbNaF3FKI3HSdDoSRXacP7A0NlJNgp8hJn9u5BZUrcM2ilIOsckaFbUB
nA9/rB3YY7tRlWrcjI9K0MnlH05+T9oSprAgrXcsGfeRdOu0Ktn56XSAeouJYqRpEr4fbY2++OvI
Efm2MpkzimFmmyOxzorydlV/kpezhFQ/0y3g4gzrMQsHQl+pHtNLM08jC9Q6bnI6Csdq+8ncqABz
zLxqO2v4dbxdFi14HcOGD2wWrW4hOpMxgTNipYXcxvX9DjbYCqohPZ3yhQ+BlK8vzd6l7h0Zcar7
OKRvhusHKyzEiDOQAbUHSMi/L+E9T+pWJGNoqNqu02FOzo+IaGtnezsU82ugKkV3Ia6hqolKKlDb
EULkDlM3rBOy4Dm2upjOu7TVM0xy50sWrK3VrISIXkGA8mVZzA2AglHj7zt9PQv94U3Dd6aoinQb
MNhZY3WOcpl85Spr9zIC7Ooj6hvyd2qOXcDfwD7cRdTGgvQc867cjtRpcqi83ivxnVbb7FyOXDdz
sIyiaijgSv90yYZZBHDQV8p7l0QvbWbfM9YyWOyGOVvxbAYfuj7u2Uy/dBgIPpG8rf3sAsOykxcS
t/KkyKqZ2iU85LD2DeloSaqKjMtaszeCZ+3hwCT2dbyAc/IE7T6kwoLwMxkjuoGyjNpVaYtvRmkR
p4V6YoX8OVchgOmwgREOxAja6YJpm8md+sLzfEl2b1GhFhK9ltHvtAKi1vvz4zmwyWMnBNbLGSLK
dX5Ai00Kw5+wmM8PF530SJapbROKgZ8GSjXeSjJUBXkPnJ0HfKTiB9eFH2bRcuMPZIOF4bx2r9/n
/2DNEybT80jqoI1DFStOKFPHmnz89qPPw8cxBX0SPBmL72BHI2UjZEtz7W1DzsJEn2asNx9rbFnM
wxRlO9b9w4Jjf+1wZPd0e6dnvhy8D8ND1CUwzAlI4Oc0Tp6eNY+3rYM3jQEfqgf5sE7NuBmce/RM
6v1D6F6hkrm1zYd/Vad2+GBgxldN5eLhhfXLXH4Jo/Gmxz5Hjk4ykl7eViduCqdDRG4MMR5nsrHM
TfdFltru/+PABdGQ1y5nkYbLtyGYWEuz0nifUm9BQjS675MC3BrAfDB+GSBtqmHDDIHuB6PxHEwf
fUyjhNR1Wx7t6b7FgS3UwV56vrnb/QQW73YdFUJTJ76TRlbg2Oy9pIadYGP9g0QO6daD7UDdNhs2
NBoUrJfbZ+uoz9U9ZkMnos09rmtUa5XO4cSBLiRxORNUvlOTr3feO7ta+cg17vxSKfA5WMHvmXJ6
XBWqI3MSGbU1yh3wWqvXAkD+2nVddH6MTV9pMzhJG+BoyPlbzah/GgXnbr/EVLKyiertPNWL7JdJ
/zgbhDnX8rqeo0ZzfVGxDBya9/5VbxgnzUVaM4V+Ba/UwTj77exFQY/Up1DxDHrTpS7nB0eV4tlH
e4Y34Yqq+J9ntg/LMC3bEYW4Ax/4zLQuuErauilZHzEz0+LbWDgMNDmEF8zd9vhTKnodzegYGBQT
Br+R3M+N3TGvoZaRzdqf3ZrdaeB8WtKGR42FrwbKvUdw0A2FyF9pJd0WmnTQ/5IzgIIv/SFQXX23
wHA2pF66ucr8DnznE1lEPJf3rIORgKefZEE4AbvMBCrVt2zFpSxOlP1FhQOUsLKSx2i7NL3OPdRy
V/sjestJr6UsnY78L+58Nf7dcCGvL+fimoJWg8scJCQLT9JeC6CJ8EZSXOBqAw5Y7o74o16zFWv2
8Mcq6bRrJ2jQUHbgW9f5uOMPZU1Z6s5ppiAzQHnrWMZk4RT1aKVWfjM7t34EHgJ6plWlmb41dXL8
IVy2oKkYwsuZDqgj94my1tS/iYz18auiPTGcVAbonmbZ3eUFFTHvODP0RNNEbOEBTj1KQEcvFG3a
qa4HJH5wRrbeXUdaZ92JdgRWSSuGOO50nDMoYNVR6uwdi3PBCIKJYVDMyDmDIpjuo/YjbZW65Zfs
2JTuoP2C6anbwFiThCuE+ZToTH4pt4PtuxVF1/C7WndbaXRrSyhob1A1oACrAlwC+FTO8sSv2BtG
JHOXtjkxVr5zrjbvVNgZiFJ+KJXijIBmommy26B59tIYwcrZa9qsa7jQ3xd+Ifn+zKAWwnCFYek/
uKXwzjIhMLT8/GCeCmAhpkoAnqVwwJA/XTyWAPphprw3SKX6bZtW5I5FWFyfzEHwKkLl9CIoUIZ4
C8nex2idVbf0xVG117o8XyPuVeG16TXnI4TEEKENtI0XKZ+8Mve16UWKnfd+etwcv1TYYQKdN1sx
IArN/0Dea7rC+BXsjB4bLyb6qaLhX2AlxdblCJ+LsevGJPkzkGjZ8fQCGg5UmhmwnGOzZddzgKDI
iAe4YV7U2crSWFVJ3689iFJkHmlyPfl6BE+6n7WfqIwAotLf/qNe4V2CA4n5Wv5THPkbeyW+lf1K
+YHPTRLrwSdiwtMVddk56b2YM3GP2vHiIGOsTzgtsVCwmZ/6vNxzgkrqxBRoVOtCg0kTekN2fP65
tJ9ka2bwmNTfKYJZhJ8QUCK+uOAGX0Epcf16fm2q/G12oWnvFcpsviQsaOyQXIHl3LEOLMKp+9rE
4/HW68EfsDGCrxSrg1NDHq9GalYu62dFNUeKybg4t0HjJ8xy49GTjEOEZ5/l6aLU5jGr/bgpeBs/
bEy5QBIV4dW2A1tll189S4EnyGBo8Q9LLwn3WquJmiYybDGerztnIyfiTfDAgY3b8hI5+wpgnOId
mrkQL8fnd42N9VY5uSf29snAaqY4UXyU1GlV07vA5HGvtU9nXqqPoHpmy6yTs4Nkhks+voP8K/aB
Vic3R9ZGgaAz4DUd2Fq3sImJlSmTVIti4tIJ8XTZ17u8YlXMOWxKPpTSI9ehl89ZT3SaHPqUvE6t
WVE8HDFgGPprPLtak+6NdQ4wl8ouGnj7CLvQWFim7HAPNl0IvjGK7RN2bGY4rBIzPdURO5Iw8P/y
OhDICJBMe/IyI8W7vSRJwEQhTUx8oAu2MXDdWgjEFE7Z2Wq27ewPrvBcgS6AY/Oql/jvu/63xB1y
8MireFuTBYu7/FFUs2STkveaxCROG5zMhoO26pPmU/baW5MDeZ/G3x1x8I8/V9q9UxB7d8uM0Web
rMlF+99PwaSkpimIKAHKKprzk/CpFEhb7umDCl6fxMaSEM3RpTp1HYF/7sCrjOcATbcRpYN0J50m
5jZ12x+z5m8V7O/XxZ+UN+KOazyPAfC8ES0cwwrri2pFxNdeP/bZqhqtzkRG/Ek0nTq5KFc+9Aw+
AJMQXkTzHdckVp2M7PJWIsvx8kKfvXiE32P9JJIhERzbikIvUEsm46FxiImtIR+kkZydMW1wv3oM
0XTFjAOsucD2lv4t7JNcSNB01NzlTqNtf4iDriswl9BkicPCQmxY4pnA4DRrYg9rEak8OGtbuqaJ
GSasiki0FqoBb4+nSLvLo0poTRNMrDht70f1d1FdSC5EdOi/qCgJvQKlkSdOz6ZjBa4xkN0aMtkl
QDO+WfxlwKPgD7QHs/W1Z4m21/Z5dA0cg1bI28Zyqqpkzri4hH6GR8XeekkNXVILNDaLF1HKlKEL
bB4UKKStzgTHnvJiRtmXoebC2+tSU2s2VwEF1cACiZJ8tXsYF2ZukqjGm2Ni39g+pbyjVZdKj/Ij
m34UuVF15ROG9VRESfk93AvBsPFhT00Fjt+JzYa7iVQR0d9qXIgsL7jQnDt/28+8/kCLrDroSS/k
wXnjd8gdicX3ap2TxcRgJFXbjYmzBr8NTjU1+vu/K7aejiJ0vRBlAEyU7jbWcyHyGGPFui5EeLs5
hZ6CMN0Db93anYfxUEP72WfhvmpJRoYbjO2rX0eL8X/NTRXHp6wOFC/DfRnq8Z+q8+NxmzJm6xyv
eRukw2V5pyc3QDt/ScXT0uesQtaGXpe2wRwYzyrzDWwztBUwL7OkmVlWLWzTgVtXsRoXkXGosMVA
IU4Fzcu5dE8jPoX9OmsViHH9R/7ue8y2Z+flZqqw+IpiFjHCkRD+VD1bP9HxMlciLtzGWE5tNTJG
oTzdlaI8lIhvszuDyXJo86j49FvYVUzhqRx1HEc733CEU5/4dJlqDfEFg9Y4iJ4gV2qM/SecNP8f
9jFlFc8nxU5gDCZQdFjZpXwbuUBXUWsoy3wAqxKqMnGn2WHG6m1WgzwloS+GeS+QtYFY3OPHbTMW
lwDpKks+YK+nWCkskHFby1iSKE26XEznjKB4MwehYsoendct0ioSh3cnbZQCA8Gkf8ADMIqHrksa
4Ykof5lmLdyKmYwsU8sJdi0ppzCjEu/D+zmMsyB9oSpkP6yjq2wqkoscYTugokaUWoE73PONFknu
Oq5HYWTPaTWgL2Y/E2IqUdEtfCqZmT7pbEyfSYSYRO+5Fursjr/UsQWYlPESQGZjh787WgudrC7r
yFMgny+bpsZtr46sq/LcYBJI+THmI1OVgOJJ9SZDz5BIsQz/rurxdalU8fQE5KOUx4I3s54VfZYd
F0FQpjjwuxyKyF9gn+CAo+C1TsIFWcQubQ7fkSKp66v7TuIUPTicFyrqrMhx2KWgWb4iHR1MfUXC
gEFCwJtQrrbKIjk9SjdUhReRnr1ajNGer/QnTZYRTT/v0xIoEOBkbiX74mh6C73LGMo/cmsfQMk9
F7x9TunMp48dOmFWuvpxI3xm4dKJg2gt8YfSy17eMklARS86ggEnn562XNzIqVp9RLck5Sqr+dVc
Z/LO+l7Do7WNCMcApqLnPzsBeFcqbdtlT2tG+SQ89igA1PuJY+D7p5Wb7jjQZEFv2UIhls5YNChV
xxPXDWQhlUlnQ0vTOs5FXfSCBBSfJt0w1Ts8LgdxJN6MfyuFRQeM3PGXNNN7tLuiawsCNHZptWck
aw2K9Pe5C3mcc4u8f0YHP5YMFBtjPcUV0AzKB+mBhlRNFXEZa0eXEVBSKYSXJ3hD7f33pZxPuUcR
OOzgJQYyZy/VOq9mH1wlgUlYXIgSWYUZF82oq3TmF3V9Z7LmoBd4QhY4wNS1mUJfKaMtDx3Capv6
nI+7Oc9GJKTQU1e9y4OJ5vM98PCpJOFBdigtBLnhY3vBTNsUOvgPZDkYHVhwqP8tfqgFFvk2Oktw
j1FYROTzDuL+V/r9xahYuTzsBvz9e2ZrmFo7kth545ZRPkLlj9wBR+YtV5Eu8ixLM6Ol/EfhcqZe
66103zRYIX9lG8uJQqdtFpJbQ2rQn7W5p1H5JAOjUQfpjo3rPfew6iKcTgU2SsjwgH8AMEH4YMay
ZA5jr5NHqcfKhGK9nZ68VHNGUgL50ufQyOSpPSVyg3lTr5FPGiwwn0zbDERW1NK1YD54hJDke87r
m9PDoXRWSaoAB5UUlgUX9DZElexP7yTmIURnOy6XjzhbWvQz+rsystcTO7JqnHMbJsPQfC/nnCcl
OtgUBmgl/GDOgr7KbFd3jdzOLMApDZstuh5RmfqL9pEqu0PA+xjXFExIEB/mJY4EYyk0M1OSnGFo
rx5RLcsajmGtxdPCszBLetqetqKq+8dN2bVgOmu9v61BRKKvZYz56dPVbxmmNBLtOfoM90S0QplF
DoXh8IQOr2XG9mFoXPL1XJBVSAz5fFauVQrne2qasomLKC+rRkfNG3rONfjak2TDhTi9/YcxOVsF
IzQ3BgGedRAzZNiaykkAYwtAbaTR9NHYjLTw6wdoS2w2QWeJmsbueiAnQ1PdpTL5lTS7VziztZ5/
zf6qz5iQmqgMWlnLpTPQu5ySaigSczbHD4bL0itj/xA/P+B2RRn6TRbuDhwpk1Z49GVT+pWkOcGN
MZW9j4qUCmdxkFRtNeuoW9xilc/Ar0FTlqgLDQV20i7HAGIWEZ2sVqI422TtmOZONF8aK2AtoFVZ
0tFCCH+1sBUgQ2TxCwhHJaBFrleaQuRIQKTeJLjnK0GPcoUgQl8ZPSZ5KFOMuvmOzfUy+1yU6gzv
rdyiY/plrUWkkNqkeJhpbLIz+XsbqevpIRdP9VqKkQrcZ0KBsDpV8fDsgP6+gT1Eqqys6c23fpeQ
ae6hEaPR/2ucSgakn/BWbYpbYHiHcFH76vkCktW2OLXYk/rtnv4CIsF0e8hAEL8aSlzD2dMT3Vyd
sfBe3OgQ6RqJdE/bKcMTiMLvuNVTClzC24R8BKdfHq/0U/Beb6xWRlQ09Mpa+bGWyXV2y5Y2AqKW
0h+MldSID1idB8gH0UpOjfdhBFbgcAxyzYIL81bxhRYf++fvVP5Rym6cyEVAqctdqgW98KW3tbel
F1l3KSv1L1N5gmUIHO6HdOtga53tyM+7DyINlnWbx1csRuoZAno3O3IUErY5Dc/ZYk8/yZgXk4f2
bEgMXW892vX1TI7+c5Y6DpmY/NjqHiPrIdaSJ+Nl07uuQ6TPxKW/8HgweNQZkaKJDXR40i++SCyE
/3X01L8dAx9L2/dGegsdFFXP/F48BLaoknYHLpyijscjnlRzvmPzW3o7fYQyjIKQcfXNfg2r0KzH
cuN/TA22xp8LTksEzwz9choLnBJnHHDtp5BpR6l9ZbCaHpUDUZPlfRukAfALdmH100QupNgny+XL
50kYRqVbvXh0K0mD58C9LhqzAzoBiM1K3Ti/B0Zm6ZXqvQo89B+F8eDVjkYU9ZJizwW5zm2h6bSZ
/o9PB8zlM0rMl8QZhY+j7Km8K/F4BTB/J318raTL41YJ+2OIfLKZ5ch8Spxvv3Na1ZFNS/+yGIQi
uebNPokl4rmxm2wjp3BnVr6ea06MOduH21LKTIHKpZFTxtd5iI+MbfJlklsM1JrZK2SuSWZE9RJ+
tJUpDmzl62fselJGcgKQbZNZEU99g5MYODrLd4SmCYhavqMUahjXWVMpcRuAVw4miQPECG4dnBVi
XoRZN8Qp7DlMuiee+L0FOtR0U0mbf+WpC5Qvuve0Ha8nUDbR6kT9Qg7GsBqglyqlipovGUKgoguO
PtPE2QMOziiyqHYnYkcvVj7RUWtbWiNYWkAM7BMMWGJjap4XE1C5O1b+gBgJ2AyZPmT9UwZZFwYZ
ByqJHehc3AmHzqpYkgocRgjaMtktN07m8in9X3YONh1cJXRzfwWf8rkk040PVjGJkiNrvu7RRrcS
vEqU6ica9iZr6L7iGkrDIic4gqpoJyM8Uw/RE60+Pe058GDTVp4RRSCKujzaR/VdR4s/N0VY5M1a
RZwZsaq/4saHV8ovGZa6M6MpkTorSsIwpt4lJgZqeCdiWmqI3HDTUqZIbpBUBVH4is2OUAlk8D4s
jlp5MqpCMBaSBftf3ahAGrTdWkBcrrXWZIlVYfdHn1a8aJAMU4Q00GTWjd/0iRRZEvAKSfKsRcIy
JCtANRcoAf+/y7Sr2htLzMY9PbsZc+m/S72KXUPVKbecmiwlRzEoOL9M3DI96oetqlh9OCB9g9IC
Z4a7/vfyid2/uMb9p21/CuFpTBCAeuO7ItTTJIQ1rJJ++8+rlSI79v9jnfc9qiZ5oxInskt32Hqo
yx6jfWKJPXTrR6bb2u1RwbCxkPeuFvaDh85UZa5Yn0iTl/c9VUbD9LeqZ8Q3surmh7TWe4F7hKFx
MQgAm4LzrAekH9CSHO5rNH6XB6RgVACSSN89s8HLA6N5IBQJXDI/dWZleqNqXHcZnNXG36ihI24a
J3vp3dPzLsgrKqw3mXA7WVsaCvvbUweCCbqCMxFPM8IlNw7v/u4/ow1YMCHkvl6mjC2Xjv+bXaMY
aLcTjU7vRL/CYJ1xHt/UCW2W7aqJQ1TfRe0TMwVRvLtI3jghs4MLlkKOyUiJNhw3EqvCLcJpTWD3
RZ5OFTSyJlR71pucKksdR6mejN6CJsJG3C4NlFGHWWy8NLZ1IlWsWvD+wvAEtyYny6J//Q/ZwUs/
IbakE4pg5gd59RDn7fhd86x+KZ/AZ21VLy+ycbdcHEhyoNKEyfq43p9n6Fu6ktACq/+aNyk2XDu7
NcmKNulMliXhZ9Ye+x6ExdGkkFYOpDpv3lfJULAqh+HRLQ6mqDg8ld20/EEU1nwaafKhjQOVNhO1
sbMvWnhsyGwUG6EE9Q7FzpTv8cFFN+z5O3tHR8pWJfXQlPfZpZW8beg0yBUWyfGuiIHeaartR+Ht
B9pkcDZYpEoDWE/1KdNNt/Z9f7FMi2V5zGc2+IlYhjO4xGEXXB30noEns/UIhvCrSE4k5nbp7YYg
9Eub8k4v2pGjTBWXXZLPe6WQ9kHaPS4ghWC+upxoZSjk9poXmOWSTjAZpS1SOnS1x0CbsLN+Mpy1
7Lw6z2LRDMIIgAjwQCppQdlYHzmTqWHnJOxuP5AHqDPDZfQ7IpkpLPjcKZEEoN0g/SYPacBrz2C/
W3AGTCsR3uzzYriIlSYiuh3jkB8FDE+wwLQvqhrt2hoDK4vRI77GW5Xj89yCVfMr87u+UivX5ey0
65MW2F43WdPQFcpQTkqp8u0c72KXJmdOK163kTvOfRRxgE0I9ED/d1NKYeN3Xz2R1Ciq9ujjQqWp
PEOEJqyFIewS7L5+5oOI3f8x4qmkqZlVNgtvVn9B2YbrnWqUl7DJJXFMEE04g/nvPRFzMBBhp8V9
3yYTsRI+SpXSA6EIKXo9TEpexSwxj87DZ3M53yLLV3ITBUr0fPX13Iv+p/mY9xtLcwTOwTImP65c
Gfa5o2+DXcfBJ6mdfjw3M94pWVMD3UpsrBnMo3HBCfsBjKx1URUHvRg+kn5G48dB4KaYg0Atq+Zk
r9aYrGKscPEULtif5b8YX3yaUYp7SBw/JEiUK+CRNT6R3qmRU60oD6KxRG+wVH6XTBJcHLNRFAOc
eIaPmTOZEe2DpoksEVVPhXazU7fTT1tu3td8Na8xeOjRwuKBiDnc+mF/WV9mjoey1rfm267X+zpu
8UBbijsepYOWcagvfTCZ1TQnC0HTJYNN+v4zrww9ruE8uAQb+gTDt2cWdKGYCQ8Y3wdsI7UJLdOq
+MjXQh/5uG/OmiXG8RRZ1qGSU2FkBWLqveQpn/NUHnHab5L/WfOAlOiRp4DxEA6fthmFTud9xJ4W
pwIZI3vv6+Elu/CBb9yuQpGZ1aqwsQLFj+Vj+D9DoE4LMSzXBYH8PgfYZeyOiZKBTn7SablvfnJB
hg1MoBtg6Emyd8pXRSNRtBG9F/UApgQIgfy2xui4FnSKYkYaagBrWbebb5iXYu2HZ5AOHxUU7TiU
QEiU2cbMqmzN4u0EzkvmxsWpJVPCk3sjh1Gi64dEXLwKusDYVir8nOE/RIq2GHSMObqU+amDWATF
2sUTMUHRr4CrEb2YxGspsvimYWX4a/60gqr3xFzOPXkcc96/VoG56zeZLBXUGlcA+KflIcYc8ZTg
6ac4dtgKkmn5ZvEattBQPkhKgKUfgx74rxvnIN0uh7/vJ/h6mguBAviS1t3LpMr70lJ4uTVGg6tW
ClEx7LkWcCPeo2qR6Cet16NFo/4KpEdVIN9nAkNBihQTLDA+GiLc8lOgxu9rEGAQWdmGSqBtIkUE
Peix0i11P3j3f7vMRzb3efxJDoU6kHyVaIv6HXPk6ql3k5yG1ktFK/5GwgDh0f2ySh415act7OVm
tRQr1/Psx5YfbtYL/YH/5kk9lxwv6jme12JAkVXULabsNTEYqEuEw4KX24nPaWJvGAO0I86aztG8
RZdFMINJppkFIOawP/kw7QWl4y9jWsk17NWj+UfVQg86EG4M1sMX/6L0cRMl3PG9h2HlN0JXvXe1
e63aALg7ez1hExJuQ4FV8cku9f8I8HarkeqgGTfNWKyw59YqUItsbbPnbNk7YcGMbW8hrYj4khqK
U0aYbpQydcW/MWJKZ+6q90kvlwXKVJn/3/+Zt0b45MUcsWuE0z/Onnwxlyp8c/EPKtXsRfs4jHK9
JQS8R9XWFsaQOb41tkMSbiF/RIkbFj7osZR4F5tkXrHowkSCZ5Kf2UH/W+ehYFdAp+keHSuHaBYC
jsGfJjR0cQjyjHYO8smyUcAA0WeXcaINdH1Qw3Jcovr5/iiXNMNEFvVvhpjfERHc6U/7M2MIuEn5
SzOo0ljwT0ndd9iU9wtBJtVVM30fJ85ihncSFRCNNozwPnN/nD5cNFZCLYxGKcrX3xpydCAjpr4w
BIkSKAnDER3AJrAIK6lgFtEzYLLH3a5yIaUHM6Xd6sZbFj1FRNTtQ2xUxD/vbUBczCRBurjzKm3n
sLFvfhanyZlKbkwW/Wov5fZRiBIduf8dxXiDSwEzE8T5OdJhVc3NKDwFHzXm9mrLS13mh/MjF2qW
jKbIempNDsS/65nBJC5fFm3av3jvAXuUNKDUwCednLgpm2DW41ZIofXzz/qD/UBBzffHfPGwBL4N
fZuvdOdgt7r/RIau5ku15F/AvmCWZwJslIulbyQzm7bnBSt88eqkx6xxUP1Uz80sQGYWp3IAtpBF
4mVkEZxTmGn0AVW6+fO7DtI5YhQNqTqmoLZZ701Y5E+oM7zt6wsXW3UrmkBYpRcRtm17iiKgOuIy
Huuo9XSg28R//lUvvWNusnASpD43WNy0Hgkgr2k5GbqNtnDehU6RANWRpV206N1gLXQv5xKPdj4l
7dHlGtFwbWUYUKxienncUUPPG9iTw3zsHgv6tQ+q81YXfa71t/mKHE5t1nla/o7qwb/oflj20QRy
buwWcC9OeiiLw1J4s77tuUS9Ln77G/+4N49miXZAQ7Jr+4wTX8y6DKNCqH3hjHdCcD9zYDzsaSqW
VHx9qrH02bOMWFVPSb02wlC1VgxXLLIRE+mY6Q2Z7FWRFVZoTnRPcKfpXNfvJT0s2XN11UA6+tqE
R4tCSNMMK9X0DxTR7/r7S8eAjHHdZ+uzptL94lYDML8AAUgcRm7aofldsi8twAcbyNVlq3xNeZzh
Fp5M+GxRUmPw54Yf4+FzqW75No2IvXf0K4xEoQDZfiT/wR2GqpdOgZyWc6GHEioHwmMsPxxBeOlM
TY+O+IXD35IvEmIi3BP6/dwvEHZpe94XNjqCWNbyJKZEIqiSdzMYqOgCa3UF7mNdWbZjRjn+N8Bz
Ll+Lq5tWyqhCftcz+I3NYWGjPv2EqjXGZ40jZi/1aWTWN3ixfBtTmxgUPE1A/BmqflsTGHX59xlF
P2fZL82qClCBpmc2HK16rcHu+/SnAKQn9K6h8kDCHs3VqDtaT43RrPBJqloGYFj319WTxopAqylm
pGmqafYCAVOrFncLw4HlPYLEvdh8LYYUhwfcTkaaavuyIJ3GqoCqo6awRbw3ZClY1kkEgokBoQlL
DwzMvUb1W+pGAELHLJYRjXDn6jR3C1ymk1RM8P65VM7ejOyVTURIv7w7Pt/gXdLz3yi8ZXmxIMKF
okBACPPmIte4qCBjnIWyKXTbgtcKoZFJIfacU95qghFGRQb5FEVat5FTMVNgLfguHn7iJ+eFGX9/
Rgwjxp925W7LQ1YYstcnXgPhq4+Pm+0IRC56DXRao7sqfCTvaykGqgeifNh88B9psYOjNA+LZ4Uy
5MnUg9zaHv7bG8wUC3vT1eH2iGoEvss+gSJK+kZoU7NWP26KZKYh3tj8tcjzmnZH6pJGjaYdVgBc
6S08X3kbr0a10HCBfYtawoUI0hKiORdpk7vbcp0Pl6swmzbgFGxH9O0Cc4nBtGYuV9MMeHy0Nuqo
e3iejqfb7RmZ/CHECHzqfEZVz4WMhYs+fpiGtHJaOIOKtHA+8yosfLrn7Hi/+HvPugAB10GQ2uL9
Zh1SGUy3LeF7Wpk6fv3ceWTFg3GdZtOdJlucDkznha+8XomngAFOC29j2gnHxCqQ59WmIVqWmV91
k4mQSajotYFMAsgkkMFVPxWiMqwzM/7x0D8JZ/bpiCuF3tVnHmzGaesfAG9lVozm1ND0F/aHSdMY
HcgrUGFjg38+OPRFwIrycC2po2MBzdKZC8fJaMV2AQRPB+psOtU2KQsX8+9YHQLJoSCiQ+kKk7wf
llxluIZ6nkhTxXwQsLQs9GO+aTEy05caSo138AIkbAboCLZJJCLUmFIcYFAr5d/v1q3HMgshUvjq
Awl6jgQqVesmkoTvI7KC0D6oddzRwI47VPfhZfOKhbn5keGokjLKwKssPO3pEGv2PhQoqUuN1+L+
aYLzYqqd+mLdBCFfR5fCJGOodl3oYNOv0Mb2zJcneydr8KPpL6tWZ/Sgx3ahitb7SLxdKisccSdH
oTw01AZPfLVmS/3LoSzmzG1eOJyGrCP8jtgzr/Q7TmJEIMxaJ4nKCwjL4dX8P1kt7+QjRsx6/YUK
fFZaTNIhUt9VgMkeFT4iMeWtlCbWPHHtvwvolpqUTWg6EWEuNc4sWOdhXEadRJsF36tNCwSD0KDH
NeT7gqs/okQ9zL7xZMeN5uEH0PDO8xv6NskOLxClR/quxVc4xd0Hv/8bvEUmh5Bodx0KSApMcEJ8
sWdMIQSyWVguH0cS52e/HGKKTxjoA5UDtA+f0+02AIHUi4nWPhWKRG2Q3Mxo6I22ikktbdxK21y1
przMFdH/LvIw72LfF7Z4mBA0Zwn9j5dEgvr/05PvCuzQnoyzdQCfAad0FaNlEtRGKKu2iVbCmluv
T4l+POJkftsxrXkR9OPkl4Hczcb+Y56DnVY21ppYK3HdyYSZR9l9VRbVcphp14t8sGihFm/7Qyh6
JsHiii7BGusImfAPKJrVS9lA2SR+BaJNF0/Ctpa1cSH1x8+BuzAtV4y17pBr6xYqmTYa2xEYXosj
PO/877O4Y1eP7VDn0Qp+NCDyGjN7aGP1bzv7HQ2ryzBvh/A1emnwBTop5cgxNmeGss8X83UiXAcJ
PyBEpi45uFbgWv7hFsYenQCfI0DBHaoUvjhXrL8lYNhKBRLRRr2Z4nZtHpPOpCvhvr4n5Ws5Edjm
aXsM+5By58fy2c60fCJG2ieO3C2Kd0RpTRd5OFaxqKaA32h+SmrdN2+YHqHtr2L586QnuuIutbNg
6e4K2uWNuFmFOn0WwVBp/y29dUCwBV+OdSliBTDDVzZYXM76L+7gt0xdi7O5g2McAsArzORoKLrH
ajyfZhws20RNUS98lTplTgACqTDZhEGf5H9r32oxBU8eqyB+q10MWLdxpbAVKpuMRUnHwZ4NHnU1
qWXp2F+fs9M4kY137QYpF6z06llFQLTjRAKvwthkfrIhLyaN9mWv6JLStPk+GlYXWFT0I5TWKd+X
LhlBcAxWMTJbXU2dMx9bJ/TllWr4WZCTMBCw1QhoOZ62ITIFEiDWzqD8bXdM3xRq2Mt3yN017Piu
AmjGP0nG03//cFPN6n926TjliOpk92QyEBLyMYftnzp1twX95r8wPupQGfk5AOyg8+9NWRjAdv7k
AFkBAA4SzL2WDKfJPigslKAJXU+FDwMxNzE0jh+jMGlQUyimzh0jK23ljQOxt6Yx1Ea2n9T7Gcvb
DEpHPAPv+J84n9iykVs9mxUCMIV031Cda8IMRARjTLFp91+mbyTiuX9jXFMvjq3/I0ZP5m3VBRSF
HchDmf7hriUubfQA8+yTl7SuNS+QtzIgCKuQzicT6nKihtJGan/4ldGlKXStyC5EhxTLTtIoHwSN
8zqsjnGiIbhBKsJlQm5BOalMrm3LvuDLffKOPjXuHxvXLCzkrYKBoWImFI6looh6Qs4hLhUIvXLW
bQ17eQasHiorrd7DRN/KLgOQ/Xn1eDfl92r/DUjhvM5gDuflnM/onEOpBSMBXqRdZtuPfyEt5B4U
puqbuBMVsc+2p+x6CAekN5wihoaxp6tG11ne3WIBNWHYhJWwX5ZH9JIv80p4Qt8qnC5wJbZM2Mow
PLRMF9Mm31JNGpakbFwWqDxKOrP6cpA1rza2PZl2jj1htpYWSgrEtsMSiRi9GHqaa4cvC7obxzSf
wNRmQoRVTulXihkI0k06ZLZIz1I0w2VzFSDzi4wMXIgN9ZxYP5o/RcQdR4ZaYBsEWIGKUJ0iwOTr
Tj0LY+T3gSfR2jdMOTJWrUxPw5BncBLsnU8yTI5L8ArKhDCCCcbIawSc26PebmavaN/wPJBe1xW5
KvPVdolhxNFu9H8TOsk2VUCHCAFVbTmaHw9t2tn0XKDF4RHkRzX4Ko78jrb3/VDcCx5/yNyqpX/Q
ITeoWN/92NJivXW+gHoB6RkKNO0sR6HATOFbZRCnm54FbfJ4skMkt+dvg8Gravm8jgyR5kIXAxIt
NbuvinhQGaHyLrzec7QVf0SI2uu4ecTT/IZBQOxmpPbXs9k3Ta6RwVCGPBv/Ki4Qqkluyeq/rBwv
IET4GEPHfKNBuIhzwkurFCgKMOLYaOA4LCtNT0XrM5XPXw1G9jNSxy8vbu3Ym2/1JDqC5Kl+ZHlt
uekooE1ZXsD/nWJQuie0RjL8y8VeS6qtIQkujfOcrX+bYQZCd0PbOASbDGssFr4qDKBWFSXB2+67
FvS0jDfzH3woYH65ZB/6r3rqvifU8xktmjA8/RpjUCwMAz6HUQ8U7LMrlGIcFZ3uIfQwTJexIQzh
B7mDL8G0e1O/2hdQKcd0jBtULX1LrBvQ+bEM4dsUcqIwv+zLoUUM914EgIzAmMgv4NZPjdo9ob9f
1adtOBDVvLzUwW4lu+U29OOQc+s08LNrTxvaEupiwleTB7Cdjq4bs/j9AW+C4dhi0jicn39YsAQi
L9KIVTOqM8rUAAyvi5AUoCIh2wLKS5NP3bIlFcamf4Z21X7iOZGgnF6qBtvVBGemJkvZklRlMDq6
hKNBzJiCNHdktfqFA05AzHXRgZCkxokjFUc3e+R07pghe1+ZR7yiPZbUBftZQJfurFu6xbups2k1
0Co70pgcEKjuG2l8Bl0Rp3KkYASMBEr+PNoy+1U8PtSZCDPNg9JL+A/CGhAKrm9AfOht/JEy7FwF
/aHRYy4MUH73bKm8LjLr0RgW//br716jSkUAfdXXJDUJTgRKqRnPuc5gKCPABoM0UeUje0MEsShE
ZViknvqhj7o9nmbesvz0qUHKfLpcqAn663+adCNskP9N0vMpVLHuSgP2LX4PxpD01GZ243SDx0AH
g77d7rId/Kob8H5ajXERXNMNsn2xuxsXWTpzqL8+UxODNKjneX1ETH9dhcREJNjJ0w2ZxBWdCJ+g
hLM3ERfs3d490ySfJlZXbQF26gcfUV2qs74C84LGPCOQCuZ/MlIGknfQE3jRv5BQabNgQL1Z6/E7
s0PcAPr3kGSmOQjhQrinoZ2BSQ+aVuoByCUkijaZph5BNQ81L4DQsZHK2AaHSBB9vbzql6V09sso
PAuQ+uFY4XQoFP+3Blw11pu8noZ1rvWqYU8WwfpIfxt7Q+9zEGW662GluNXvnA0Ikf+htwszJTgl
5EVCHUlzWRgSCXmQBtgrnb1D3h9U6tHBqOv6xPLVigeljqco66/ZO9KQIKDdtDeVThfdhD26Odhl
xW4KrQY7g4T9KVAE3QzkSp66PrCkd3qjaKvrnwr5Pbie5c8CfUrR/t7DJ1/IrMkpDVqpSrcbbX6O
MxQk12y9FCll+KjVuPFW/4s4+jEbUQcS2B8ZfMpp3y8jXP2NZrcYBGWFTgaXQV0rOhu2LxvzH0eq
We61/TvxGK0688ZWs+3fwXoKCgWItmvo/uaTkBu2cnM9ImCIypbT5mGKM10UcZvljdN23VdnIuw2
4Je23Icxv22rQK4p9SFMpaGFEZlakL0aVY2gTrZThCZ5tF9Ne8Z9EEIFAArv1kxCMmtijJlqNdkV
R8M5fz3tjTO9YqrWuRL/wju3qHDpQ3m8Af7BaarPMzq+iPQhdCvkftMc47mrbxeIZm31Z+uo19+F
pQd3TL01BZAESKNR/ezrlIU0jVPDWrMzol6YUjxNg9WyM+z7Zq9QzmA/K0RnCdGKAC0ADHiM4aQq
sXX+UKqDCKlsCxzgW807dDmb7mu/00ib5z9aEBxIo6CTp2B6eI48QvmBB4oyXb+OekqU4w2riKo+
s9YdXNfCMM6Ws4+WpiRhNFK8h67TziOPQatypB8wZJks4GaZ9ke26PHTcJxKIEeC6fnB00ogTkTn
egww8HLoQydZ1v5VRtMKSkM96aFydX+I9uKlgInbA1x6bfkgljVKvt8AEE36d/56pZFmvSzdCsC8
hvZqitfH7jRxePKG9ls/aOwyHSH5LgFzcia/1C5JGSknAUb6CDRpzi6mMVU8GotfcCPiPB09jH3G
Vawl0vaycQQheQhxh5DbLqsO3+p6wvelTs+h0Q/bpzUkwzcfau2XxozgoO4e0qJ0mLFayQr2hU2K
OQy7qGI/o92EqtmSBGdioPbQkZaX3lNkgD0J7ht99q8uA6GTAvMgrooRrVbuH9an+hkF4u0jayEQ
tzD9dmwAZIT900kXxT6UqdJFTVn2U6dNf4DrqbysJQ8jubHTzLArv1677EDxnt4OoggDV0mzeFEG
rNDhlwFWmFluVtGhTB39prQNNRv+mBda06RJgQOolmSaKhTOr0gALB2QxCG43bFJFItpXnglpaD8
Cq/fOEYQaS6U7Qls8ASrS7BbVbZjptXUfIXLE133AgFAmL0EecmRwxVBKLb+JYvHwz0xGrq7qfjs
zFi1zBvOaX9Wyy9mzMKczVWWZ2V564Bfb7JMW6aoyukFaJ6PuSPxBAOeIoPVtmJdp4bhbeSNmBRJ
QE1SUUaANKUFjts81w/gMBimv4Xj415T5kMR/NMwIAXTyK5EpkZpTVSBNnWOYbfLCZdh7isssO/W
4xisfCHSopuB+uuJN1fZ1HGo9KYvP0WwlRsTjtd7e6a2GOlrSekM8qyGtWi6iqTKbwggbGnOF4DG
MQcyk73l3NPjv0kfooaCFSIVRmOIzXw/Gv1F0Vt8vyytZJxpZzC9+Klv4HnZ5dcPSS3pHsfbQE8a
6bNzoXedHVk7kFoyvPtDEI/xOVWJEr82JC+ESOcqcBb6nMmqeYnCY0KkapHhMk5ZWspIzLFjX5nF
FvHn0WORGbpNfjBiIlR8+Y6E6TiARiO1hZoUrbZUb4hLD2C6I/bf888ONT/ahFGM+mavhlokhoet
ld5NmIKrMeL8NzvfTRgvWympEepuSWMgkO9tfLfHT+YZzM8dIXQ0Ub0o3AZ68xbIxQAFtKXLltcF
QKkTXn84FT3tUWKHfoR3bD5Kg2aqXL/eRrCYM9hfZbl7ruIH4uyoOZmlrhrSk4pvnt95hZOTlobw
h2EO6CEFO/05EDyA1BLfbGA5pP6hQCwlX1Iz1vPClvwJPHbnorqysRPkb5cGGDwFddiagU586mss
+crr9+We7wzfsF0gcT8FPqtG/RJ1UD0NWq+zMDE/++KOlUwvcFofdi7wNQ5zlm1dFlPCupG+tF/L
cZhSYZnCwIP92L+UIwcU0K4ENqDx2Fo9F2A88RVtHv1MrsnpxatyZLkgUmDNd9a1TnXvLM+LcOT5
I8BNE+mJDmebyADZd8FlGMtwdngwxPsUrfvb2KsqzyQ07qEDLnZUQ7R+asl+/epI6hIJXxX/vjGq
SM+uvk+WA3atq7YmO3T/xRxKfIn07VKPu4UeQbgtPYbd72nP5Zjbr6Rh9fkaDRVzEJdxg1wmK+W6
hU092GGE+tpP9+o/sLv7RLLn39LxUqb+ZAR1/5xgIR0shY5bTMGQPC0Gbe1SD+VGZN8/QmvNd9UK
XfpRGjZnxgwIaAMx3pECeK206+IBzEcueAujQZY36/YqVJoXTR9BGPm6gL9GeO/JtaRYI604D4bI
QyLjRBKEfJEr1oiTqPHDYvFMC1q9txczzRZocydRKMUmgF3L5jSMvLcVyI5WRgzTKl9ixGc6VNKy
JZ+P2h72RKIb/6bVtnsLZn04KbSsdsUvGmEbI0MoJyUrf6MYrGf9lljkkNcQh4b/ieWiT11lhg4+
CBNdKeh5eoyZISz2uy2LRIQRrIJlD/w1mdBUxWMWsFXDMbdhFUa2+SciF/PnPqPRiYXu2ZaUvYKa
KU9SiRQA5zLquJ6lpTfY0hUzjm2f2BZ0iWMCPAMSb3DN++QjQiLOUtcrXHO9aR5dmlCLk2hSP9tD
ncm6Klo6mkVCfeJsmBwbSFQ8KDW0+OxCTfPrq0wBLgFtcf52UB3OqX2dEINXoChXny2LEOwXDcBw
MNwkbcvZ5DPQrLOC/2Cj7m6QxD5waHtbuD4jIZxO8bSjIPXpFoXKYQhCnJGUHia5+B4ti0Y1gQoB
9bMmzGRXbNu7WBF3wGxC2j5MEf5QHy8+ePPLv3x4vjQmozcZSSDinPkVq/mUDM/QbemC0IJALMLS
mGvcSzcSZcMp5ul39NVHSkOIqGAJ1kwF9YK5Hp2VBrE5Nk8cV9PX8NKsvTi7gorTUfM6OEwf3lqy
vFozdLlxsvbbf7FpLif2y7xveSoWpH7a3iOyUJCAUlo40UU7y8MlUsrCzFGRMD5QfOs2GPReMWqo
K/q+OdJnQ0bkz40V4dVhsgJ2NX8dbaRpLDNORetPX4C5QQBRyr+bzqn/JYk5ufr4O5EH8xY918gm
10KR5J4ive4m5lUVRDgMoVimDzg7mPsDsQ4AkTJiNuzS9YHicBs5gcyWm+DWC+sKnLl4MwCZp7da
LfKa/eXRY1EZRElnjEZpG68KQmMCYt/KXk3glhVsVmDQbyH1w58iy5YWbbYNE4Wp1yRXUDg6ZKgq
y4yVa4L0pmOr12eGZ8WR+PoedEnOGc3bLnWjK2rbg+uSYvYAMC3HYzFDS0ypcrseSmNgAg7m5OGo
BKhFC0tg9d71VI+nn8Unsus3MdsV3s+ZdbYle+QF4yYTGv0mG6b77I6FfoQh2Mp3dm1l8nnc5Xqb
lQhx6iZ6nEtS5XidIxKA+uGwITkIiKfuCor0FuP8xXonXSoq9FLLOLkF57NMAU5qgpgf70GmfVH9
FYbYNSnq/MKe3zIhrNzOeOXU+U8XcEJ9Po05SwDB/Odys1aJbpxLJkPr8jjOpXxDKgmkAtoLnM71
ArpsG/4x5LtsEQa4/MMCyj0n4ZJ7H/xO1MV99U0A2LsoUjobA8Wn8yzvwxYiGRh4rZrMfDXbIvLH
v6se3R++pIBGtu0278JoXKGC9HLW/QYVWPV1nibPrlLSsc1GpmQfpPeccnGOAxnIRI43SkRBvuxz
FtZUTtlybJIchqP05K98DDH170UqZ7V0WL/vfufVFxRRcubNzAYIqyVUwwgP3wwGw6icwLcwYGU3
hHn7EA4XN36aHYGM1j5bXn4haXiNp/f5FC8OlkCqEuFcB//U/Rt3xAvy5Le21Q2gOzjBKAqbPdNf
WTX6Ai/T/jYHr25yxwJafpq5lISvqAy5uJY3mnhHa81KwT1SOUm3DqotLMAI8Y//+F3CBZtmFlO0
taeZsq5XBhQlqxiOThiv28d4OZ9339mpazLuwwySvm1xvNejzxbFbCxNvOKLccN46ZDBJHsjhxFc
fZxmasZZhZ5rjMQUDoz7oLSaULBcyahdxh1YA5VdEwCbIPw75bb8JSZMNkTFseLfMK/O6THqqzF3
HnMrWvizBg0DqzhlchhP84kp+5O1HfQwRlS1zxZOqUeKLivgERYzU6MqQ39yByeJcPp4lhwbKJN/
m6LprLP1QnXm4YbstwhE+lbUP4+E05hXUuI2esMSAlkFn5EtFGnmAgPBbj0gvRm+Qf5jawDIIkeD
ofmLK0EZvwog1YUyp8MouRibgpYoUK0fKreSn6ZVIoxhV2eP8uew5Fc9eSgbvhE6LhuEs6gQmbTH
oumfujuB5hLBxLtSPROTAUWi+i+QpLKWp3nBjVVZOuDz34UkN+V1bD8Pj9O9JmS9Dvqb9BdTXphn
goQyM0mf7Tx4GZWlOlY/9YN04PjclD6pzhh3cQOGVLU4IugmD/eME1V2ddOk9ewE5R329rlYdlae
xIdssv9uhrxpAIwBBaG0J/+U56gm0IoXiiIv9orlPrU3F1TVfwRGvpFBgBoA3tEpFoO3sSZnk799
WliHsOj0Ra5zhndCyNOiIsiDMK60XuKIbQDcl9obh45Pj6Tbmo0KmhvF8KwAXHLprKQgLCENQvFR
rD55UN/fXf7Yd8XLCrityahWPKSsycqJ4zBnjzM4UGyi6M48vsWLKLCCFYNLWkWNPt43UUUus9nU
at5R9n/7hqG6nZTJgPylNTZ4alh9oiiGl558UUYqqopRvaVSgyeYJ5iVOeEC2dyl0eEWeILGqxOW
p947pEhiewNs5pBigrOSDwa5bP+07fz/uZ46mTOC2hVc6YDki2bzVZSKou4qg+WzWqNV0W7wCpHz
lS1S1tCFYWhfpcINgw2MmGAsj4qP+qq+OegHp/hrq4ezk1qc0p3+faEn/NhXOczsbTgVnMn233Hb
Cc9LEZ7lEBqBCnwDbi3aOtfzfHtEmpCKofCtQ9pbcAomWdy9vlgB1BeIHB1yeKSbNSm/nP27bqK9
qQL8cwES3lv+G0W9Hv2WQXIQ4ydTc7l4Xc+K9K+5uW1Y3BvJO4ehnOgate23t6Yg6+iFUxQ1P05A
34gPKJ7As9aLcou0B+lXzT/JwQZSWdfVifLmYi+pg1UZfFw+MHWOt6afdLjusw4qSBpMuJ/v67+Q
qbDmxxmqVL0L5yqqmYYUyW8ShbjlIYHPFesSuk58aeaOmsCDhdWdcgM5lZq2Gr61GxS4YIr8yv50
Lme0cFwWP8KxlVLRJYMM63iyRWJG4W1h0f+SFDuirmQAlz5myr8GqlrGn003RWLGJW7PuDfCUkPk
wqQy4/sPelcp4/kCqZOMxbS762K2UDpK9gjy9RGv2er78OBy+XaeLKAt4PUNS49NbcfTCoEUs9vY
mUlfDtzLTlAx5GMd+p3oJN8sITM+59zPVjNSn7GiYq5zbmyCJBTB1q4WjxfxWKIwANDuqhhnNEDb
uYE9JchCTnmD3FpM7XfS9PzQsRWOorLcqNoJQSBBGEn+KT4jLc9re8bqa609Q4ROg3CdlARyvrKe
9+TWJ3w3G6fbzXH++mTgaMLnZHIzAWd0HvDDgoxGrql+89ALBrTSb+NNgrvxjeiu0nvxaUq8AAv7
W1+LC77JEqoUI4Ao9oug7O7mdERnKUX0jf1qpQ39o97gpffQoRJiz8rBmYTCOdK+U/9jDvq3KH88
mz60+NonvL5vOg9yzbndMIeuMRoxPoluEgEjT4+RoVN/q50r4uUmvW8fggZfpJTSjujWD7LPpIhy
bcUF6OTfsxAJSxQ964j0XIrIU7g5YZ47XQc1sWKcKRLpPbxjr2hJKeNMaUwVbMY5vkM99vjZDZr2
2dRlvb0SLqYLEUFUXMAEosT0W02Jw9RGLeZFtC6W8Vc78bV9KQwwn00FquL7a+/pGX51u/+oebVN
VxRLZxuaY+1rvHxf5CTQccs0Zg76j1kP0wImzPuqhE8NUFR1MBpmpN3h1JAqYFvn85S7bm5URZMY
/K+XydjrHbokHT3aQaujnHkoLHOCJnc/6czbhdPvssah8m8q6NhXr33neku4jxtmqLmex9ukhGPe
BZo+EP70c3h+wXdJTYO/NktzXMWBL79YzZz9S/L1J7ahhNdg323631kO6O0L7wHImHxQs7ysB22X
nDNmS16zgHpRXJcWgd4+kcrxcBtRdi98UAy6i/Cc0GOE2QKOJG5ec34TVBPpSjVqeCelZhE87yie
kNqj6hA0QRDPgqOqgu0ZQr0dRhQqYW/0pVMHCVfDipuw4xhjQ+PeOhOQGURzvoauch8GA0X5X07e
shMPQErxTZrNmBCfVnAvEo0a/p17nXltkq/hK2TO/U4Ixh2/SgVOaPLzMfZ4XpwKrDVhpBmdvJNZ
6/mAG1bdRV6JxUm/kmt35Exz4mK4RrcG1fHpyPnQ2WW+DqE/qv7Cw5FL65OLQDNRiLU+Q1uRuyNm
VRctzcLBSP/1+OOZNrSEyVJcEdIwLDX3w0LaxwblgcumKIj7h9gIsDoZjOSVTsJ7Th9c0s4MM4El
BeZPcv4WraVkRUYXzoizlogCBVVNoJY2RJHODEapDkmGoeTo6L2+RwM1vxXbaLAZI4NVv0snRUT7
CjUiP/baxzUSE/rW7wd3wgFrXPPO/1kuOa8zCxzugu6/HrniwaBz5NrosjDQFrkmoxVOyXs39uXL
vznRRx7NPD7KgIbHS7GnTbs9JRSS+NVqCTkl0FvE3KGZJtlE2z8CpoBOgCUilh41947wKgq8qW43
EOpa51ShJJo8hCukniEq9BqYFLRLQCZ/8mHCqwkT9FDnYqzT30khs5owSkEbZ+46diRXMMqzI6Qw
1SZiEAgsxvD/WSqvn8mmiPnScM7dMWENogeNKEBGey+UIKSWjFj+bzHuPKmX2twqJaxH/GxzfUSB
rkGy11AX5MEcnettPVgbSBpfF2K2W3eIlaDdkmPagvB789WmATVMLO8YGCMdI5xfFeZ6vR9YcTkH
UHoYDea3ogoq2FBnnFck4LqwkgT/UruRGpA+zph57YuWv8e0cQ4nlEuD4pNQGWJK4yxp/k4DILvs
WBSWBT7RtP77XIZqb9JMu/DN+OGzB+cwoRUeXLZuzWohJGZleWTSbPr0zavKHFlbuWZ5lDGheit9
ywi6XHU0wsHtJov4ZZYa0aHjI+WEVESDk/wbFSH7cLqsS4d1UEyq/yg4jdqs17OAA6wo/VMdfFCm
jlONgXXQsusxKYfE9pzsdMn6uvmh29KWqdUEuD8i2gQIHyuHGNpORrv6yF4E6n1zOikIWVs9oQbM
IDjKBMA4HsqiCUz0U/mn4wBUDcd4ozJu+HorvSKLD3B6PdZNH6WTLDnQJ7t23ndMGSe35quEm0d/
Mw8kmVOB0qnd5TWPTHRIbnokGysw2snG93dIgTETKkX0IN+SfIpWVGnZ5DPa/q6GQ7tYzoByS6XH
9139DKJVMfujgoNowQajQVH6JAIcVzLECNc9AKdjs3p2zwMKie40raF/IiwLLLubzWl5QpZR//ID
/yj7IdRwPgjz+ZA/Y7nsTrc2ctSaXGOPiFM32rYg94XU5uHkI+JgAhAf9GzFIqotEi6miPmXE0sf
uZUGqIw54jknvIrXsj7gFPMCw5xscrso7x+g3pc9m9SFAcPmJ77o5Tf3RmBOxoy58ncZhQAyS7d0
ec9kdEoDJG4k0/RJ0510+p/kBHg4pT/lSB3/pn7Q0CE2bvUTxtW+BEssRLVhitE5daJLMZ03/yeF
BIi5SsZ+b1DWY9VPffAvafwkAXVGv1tbOfrL6B12ryWvmzGLbF0DciC3kDRMiku65je5k2FvySw/
/VU5GRDnrk633s1cSdAqPp8lcE3GKHI3Rcgyb6zNxsRiz4WGjJkCeC3QPJfHTRMir6SJ6E6fmVeZ
DJmdvP+kAfMssHTTfAx/UL0Muh7LsTJ0GtfYMuqlapmneV2DybFp4ujYM/cjo9j3423NmbtjNLpr
A5zl/uwpBrkRIbBk+HV1AJmFmSDz0w5/eNJj26yCz7Q+mjheQgA8wxC3ReTB+JBF0AzYTDEOdH0a
lslzMgBKnM3CfbGOekJyBKWw+JL/TLcuvR8Ipn4OlRbORAsaHGpDvbNUZB2sq2xg6i7+JGDzgAzG
z34OR7kJzrBFuSX48yb4Ha69gakuGTSKcuyMaPGBQp6f+YfOy/pclgfZoff8khqNvZqf9jAZrL1i
10UTijeniMX3wPRettCXlg76t7N8nWIojkCndWtktkhIF6BokarOkVHVks1/VZKfRFIA1dZcVoBi
MdUWskkHwUDraHxRxTvE1WnsADz/a7ESye2WdsfkAQgya/t4YruIQGYXGrLsFTixc2OmuBmcHnFZ
XR0Kw/7zf1mWmlNiaUP7Bd/jUGQPgqz9zM5pFtTOsfYej1R6xIVh5yqD1jy8qoyBtqNwZ1UGlknN
LjlBlvJiJ/GaQXpf94QwWu7TOKjJnr8iyS8wT2JbgnvsXj4ASX4ON1SAx2aLUF+ghF2+y8Vaii3X
0X7ahKtj31cVScviHARU6AyKFQ+lSpgO+S8Ikfw9jSJn4xW5+Xq/uwu3M4g9eM9pNkRChe5OvsHb
NDdKDZOtTQgM3mA823fZMZn40xTFWHC3we96609IHRm9UJQcTcYPDUO1/wBuHdIRhbOmpBc1Kjby
Un3wEt457p4O5JwXUHO1OFcOU6eEmk+L2PyHDmORBtIl6kpw/IkjICMjmrgsxuQ7ptToHFCb8kdI
43JRje7bl4CArN5C8UFvDiAlk94/NqwM5rcpOa4nXu4ey95gahEnM/DjlxcBnHM/EMT3BxcoERZa
NHQGcvtXmtsLEodYQieZQJED1jOddCx/GDVRApwGRIOMe32PCoOZvm7EOyE+3VlS/jMQor+d+4TS
UtkJYlH1w1cmhpTq4brxpozH3p/xjaIiJtEhJzxKk8SVHzOMbfTAocZT5/irsU2FZuFbwYi232AV
8jAffZzYl4Oz3Sdw+M6Y6Zb9NuSU500BMecnoxXJMLz6zQTSDPJpV/69Lkv2lnqJWRKkyVMhiV9w
Auz+DzTDlCtBDzQdy4Hig7+5v3p6Vu+VF7wEB07trTj/+OdFJ6RsEOUa6qWpOls/6y6z1jtm2kxD
N7x0vO+oXGMYNmhRZUr4WcNSQ+ofDuy2MSrkFe0Nr6DwvS0z5zEFoIiwEeaHS/QG5tfgZtKH+mEO
pD1RYc8JLZnIaq8jdy9EHFGaFv06PMOLepnee1UM9ENTp90ntk1wZhblC/gjzgN3fdvau+1uCAdo
sv0JJfvnHcYCQB2OF+JuSTlcG4yN5U8sjWagxtUI651vKXoKEel8HVIa+tREb4SgbEDhD/toQZ51
lvA6DhCswxZOQ3iHlzORiS8UbmWc/y3HVFs92y5StmlU5TZccRlD2YvxTSfEWi4ORYUEbUdwhIbe
nyhldJmZdH5vUb9SQQSH0qnkYMsC4I3mnOaCaiIWmM/CIBAxQ1hAN25R1oO2lz5s5muBBbZ8pP9z
O551ju2cW6gU7SqbXf0KsPtis7slNJiFYTxdxTvS+NGdqu1kEqLCYpAWtj/AuZPbXxoX6lOCH0mI
J537AY/rAi34MRTg/xXSVJz0ZVoFQ2uGGroG7wRZanolc/PrXXOt2kARKvZt+6PcbX4EkWPt75xQ
UzdS2Isnt3M7WFXXLt8OSCnTGII28hVEl72nJUHDvswCoDsrDATGCkTE/qCCp7EmSJpHemD9KSb0
dgTdue+30wts+Fj1rDBS5zHnzx0Wp5/TRjCQvzw9t38It8K9I8lqUjc2kevxSI3eq4xNTRW2kief
+dZce5gD1WARRVZkZvoxvjoCmsAH4+V+patNfKsvtKGmMDO2i0jM8MGmIxsP2BeXKC9ZqJDhjQHZ
SdazfmyXmrmtcHEKnu6sroGDA/y0Z50/3xedW7bIzdi8P1xsESqyNCvNDBFcDdRfSaFdDPLGogrO
txiyg0hp757ZLzNlRaSEq4sauGzY+m5wBlFY9d0fsrV1PTEad/Pl94zIuISx9+sryT+nyi/7IvTV
CrDmB7aW45FhfTnY5kyiOObVRMXykZRxSF2IpCMZIj1CNtJg21PAIdjxihVfCaeVUIP7vlpXoP2q
w1V9FVGe4u8Zu7BeJ6qm5C1T6AeqVXvbi/KEQVfzmD6Odzv8N4LQaD3Oh/BTw/wzoQvDRyR4r9c+
IJelCc5Hy8rYD+7Xf5gT8ij4ANGvBbBc2XHgYWP21SaQbIQDjNFCxcISdypp+FmnsT/pi4wJE+PO
xBgTmEEPeGfNtuWVar8ioqFHQNbDdDC1Yz/T1ztUyvI4zCZEqalegmgePyJqArAiZszod55oUcMT
GasH1A+4nzhC27gtXovfB8KlzTmwBWK0WLGD4C+jFoymdiYG2McS3NuSPaQujlosolnVDdVmw21X
ycGb6baJYdVXbaSNMFp1NfbbM0LXE1nd/e5k1VojPQ4nAPpJxlxxMljaHn64ONmKb6tcWO+2ESni
8erjEYsbNX7+F6whbrDbeJV7V+s9XkovXZfq69AFK61yUp9JsVIYZzbXEC65Nl5HfhHBa21onW/A
M/NEq6BMmrfx6X994vsWFnwO/rXslp6ur4siftXtFtOBIDACfNuCE+c9yqKdVPHVct3KT4hnB9b3
3J29Bn8gXY2233gR4w9vd0VNpgQmoJdg95hQENjYFcEczNcQRj3WkuBsK4nNo/kjlFI5q2ZJQuuT
9m8H7YVLXa5iqvUChwXUfP8Qyhx8S1j3Q6uEPxnZmw6VsGVpxv5UJdhu50KJMKeTv+GqT+Y/N4d8
VY9t277h6Urkz6t8VR7//C8Waz8euk1gR4j7L1WAjqvk8xlukF1IQkDKcAMkiZwQl3Nytjm2yJZb
p+ubJWlHH4fNinld8ChvgSnJHbzdGd+seg2UK81Cy0+q4/R9EpKnCB3mjf5IL0drzWM5ii3BsTZI
lBqiqEcG5dzZasx0nge5Bk4jNfoweSozRHC9YLosUnINi2nM5uwGDgqU3CXYT3fgfjJDUg2Hb9C/
DCMmcHOzlAREL3GrpPwvToEN286kP8yHECa3DAO+Gd2/jtCqOMmKSU0EsiVmV0CVCL5Orf2jSdwf
Rj9g1nIs/x5EuUBc3uoWYx5uDS2/O2NmRvLqqE5gMBTlYvyuV8oQIWsxmc9NYEyGqNinRF0t7inI
seW1MNKtd3c2LLuon7/016eCVG2RZdnnaSDG+IMGsxtQoYT/x7kATrgspdxDXgtvaSXOxciSwijH
pRreMLqQQJUxRTlAfXDebC6Qdv69F05iEeeGgWiKHBATZjVx+/67ZWX1ziEMLlPkQzxeajkJHDdh
h9ISODR15CXtebqn9Nv0vFT9JBSTZDGYUeagimy6cfbc+WHPsAThlqWhiAVckFpbsg9KQLrmYSDS
ATQq68TkG49kfLrs2HIr9kMmJmcqLMwiceGahnmv+RsihFRQ+OgRs2kpRixpT1R6dZtKKOvvgh6h
m3Ua/yAFb2rvdiS3XdOfGRvuK3s54lxfc8NTUNhjQNJOis6aNtHLVzApOnB3Ql1RVj9DCcw7C01m
IX06l+rARnK5PYj9vBLMhfVCxLZ0lniA6TSOxPV/tnrulY6B6EvtwpHgYlsDKzfjZoXY4ZKQMpdA
390NcjtOInmkUKd63EXv1mLHV7M0QKXE8oKhPKFyc+phNcZeWcOUy5lBeobWASI6Hk+nzYhRd8Yv
B1DX3Jb5o17irBpSzP7MlpqJORYBT7KKsXjdUSrNrUuXonI5CfLv1zUfg5t9DFQDV6VFmYDInrde
JLIyckjhJmyW3vSvqd5+t3kkeln18no7NY0fPBSYFp8aPTUaR4Lp83zs8COFgyRm4Hf2fjAm0lXN
RYj7hpCDlkVf4DGnIzYNL2vsi6ndDLimRw2T98sXaeClnMRm/Uw0HZmpSvpFqBNMePX9KJYZ3YH9
pLUV6jXQlqKzP6o9/ATtEReld1P5JmNzxDhDH1nSxUyqwtAawhVI/YCD0EDsonYfexlMuB89B+MK
zG0m5fs344yQUoOHsJJAfrsDnN3+MHnkyQxGaEo5ckpk8b427gjhvhYRbRx2ELRoEjbDJ4AJHSc0
PpOuEKh9UjAffTbgqx5so4mke1+LRzBpv4shs0zL60qpYOu+9uPz6vhcUotkEV/hNnx3rbZIsmW0
nzPr5r9NhhY5+QBL0NoHByc35rg7yZhicKkgMpeJ2t43ueSjYm53qd+aNaL2dNsGQwRrzVkKkIlH
8mIdar/Fnf/2m/IxWk4sNjH21IKyS1w++INjXO1RL02/lM5Jfb8yvBUsL3agitfWPfw+Z5D2wvAL
BFjeQ6aO3OhlDI2Xj72yzMrGjUEy1TH13vpJHazhKN13Iq1y07cIRPLw145ugr3Q5SNHbNXp1izb
YyWaHFbTiEa7TRcBEHBxqYjsPtqhgSF+/UtDDl8gUYKjeCuG1EHP2eXtVdUmJ0wAsp9AVAxs8H4T
4RrfgToAyq0DIMfSP7JE+cwpi5FLiEd6aXtTeeNNzMIdLDzAFy3xpEZP1hlkXMo4ztFutrjrJfs2
4mnkFw5pij8j/O35nqdHIsdPhGBFxGERGSCjzBy0gwmFwj9/OKIZUv6E2WuHQV+iLFs9pSItcLZd
3G3ZoDyOFnNGN+UFh51k7b+v7J6sMT9cUKcvp+1PIuahLY8bciApabe8DegtQDePQ7pgCGLW9LRY
IcJG/4L3ut8A9Pv5TdqDAwtYeURwvpxCJWiRZEegLLOApYGjONarT5dQgEVVRwiUXrfdS4Cow/N2
Q32OPXygl8mPOxFdHrAm+SEY9HmSkYJuecLfB4AJf7f22WKwNK5dWu7p/zolseJWRIFW+1ipdwhE
nqNUj4njyjWmjT/rz7+XYVZuy65DoL3m9nhZvJZ+MeYrG5R67i7OsNoxZIslmNyMu4vvjJUlWkdh
ZODxDZJKCyhSkK/5LdzAkI8lGo000xuEKU3K6cJw6w1u/pQAinHXs3bPTkb+I5m7dVXRMm+Ulla+
63F/XR+LkjEZeGlM/mUxu7p7GESDWeQk7rYKRTOkxPhBO5VDyFzrj/UltyxbM0BDSD+Tr1r2Cs/5
/BqEr904Spxe68tixy3ZFWIciOGqSYZBL/WJS7aNYV53sIM805Sty+uItY8Q8CFsQ18dMtbVdhGN
Mp8W0cqxMNXG1N9FkBf6FpT5kIjGue+u1yW4aBZO3kJ/dlBsSA9WfwBGjZtonwBsJaJsBs3Rjjyx
58vbm+KBNCVvJYLDLFD3IpLOpmE/k6x5Xgao+gQ6dG/F9GKcjz3if4rjBbALOJv6zRcOxh+tvbmp
3V57Yyxy92eq1HRJFRLDxerY/bEvUhcWdt+McHUUJ8/fOXHRivAhdNSyKv1ysnQ89NhVNWccSl2M
BWaB/oI5EIYGA+lC62kpT9ZuTlePBtCQIUwtrhzYbtdQ+j4KivT3DROMF7BhZDIrqSJECsDuX/7L
zoQTDRrcGKO6gCAC6pax1QdeBnFpIS9mPPKStZhDNHi/d475MzvarSq0Wwasio0ehhPVVlxeLx1b
WpUocusUgZqnKI5HYdRnTXXMpEw99hjMzScuWh3Luxs6DKkxaxQm8SKgVrYVk8X5DhmW7DHBVbJW
59O4Zi7MO+L1m36lh45aL9zRa5Gl01bafm1hhV/Ybqp1AxeseFaTU9AwThuGJy1k0R/DnUb9bYff
f12fyXZpwxxygvlNJep8JhMi5smcwR4abi32YcQWmwcug+yD8+0jpQjf+C3IZjEa2pzhifJ0CWyd
3nMWI982RdbGhSBxlVvlhwQgd9vr8hxgmbdzcgiKmguejtp6jz5uzBXZmN4cKDudq8++UzUKDxoh
uAPUqJs2qemeU7AfsaES+xmib5EHEJvdmjZDtPxv6nBXVxX88XkfMsvtqLqlYLy9q7cGKfK84yRt
wAD6MdUF9yhcz6gOGjbQjZ1Hj74amIwS9QgBNYLxyfKTVEEoCKrp+BPYFBjVwQ26qGiFjlZkgxf8
3D0s6I5p+Cn/BvTiaBcqOJzt9GBtGRY7+tU1X+yUyxx0SEqHopxcaJXPJF3rkci+VwLfVKYbwpto
kHjyc7WN1F02HpdaKnbItPlXtNvWByAFZCCbY8A++ojl78yhqh5RN5BCf9INfeCtGhZETGaPW495
mB4O594uuyyq0ag8i2GRU9WHPmjKa+S7MxS9KqYAZoyzKcw4N+MWFROd6Np/8+85uyi3WMehaj8e
YzYsmFgnOJe45WuJB+2BYquzs+M8Xbv3aDKIe7JLXFErvQk5kXMLp3kR1iBbDGk+hnHHIAhqvKh9
lmBKuKHhYecn/L6bJZYVxStySYA1fWfAadHsuMLPc47ew+8kRc7OSV3fgj93HafYgQf0q+cLiMAM
z7kFY/KQl0qe5CMd8I8/DnmNtRAsnszlPdxm2ofnhoc63vfvHYeYztNt7IuzyCpBA8saOOR8RCrr
78RsDhqdX+elhlRyqPUquC1PkJ5jFMBUowBEkifHWYMpU5cqgwoIFMbGh3wYbiNz1QaAaj9q7tlw
gyl6ZUQOB7UrqMuSShNxe8DiMk9Smo5WqsC/KDU+t7Djycg1c+5OCM+Sf+ndlkEmxhNbclFHO3fA
9L6lzMufoJbeQPpyUUiLEgXlDmN4v06fgTohJ0RpDIGdqlNzgUGbZeN3ny/Tj6ZAeWqywrpZwsqH
m0kFmYz948t5Z7VHJ+GbjU1CoZ4d8HOiDObiK4VV7YBxT84oPJ/LLlXeSJ+ZiqmZAM3cY9G1/h3f
XXK/Bi6wZqvoaQhHo/Vz+3ZBYz1Vfom2RMUNlBR1sP331e6OOAC+B3upbrDHnf91A1yfUFzYIF6r
Bj2C+VFsPOKklyYrYAgIxQlUg+Mb+6JVRNvKfdNO9ErO3tK7mvqVt3GFbQZxSgT343buWI632lt9
Za7NOIee9ZqVFgII/qmm/PT1PFp69eywkwBTauQyuVvgILBA8pxn7AudEToVgaOruVMA4tgbfkWw
co4iYcY7zWoqwJxkrtCKhpdokBIsbr6Nd8oPIOG1995ARe7LNAvjUF5EeMtRQe7QzwALbyCmLTHq
9vIxOYZt2YrcekCeKtsUQb6Pjs8KeeXYnjm4rTX1HDL6p4/lvY6rehuvAzvnnYDnH9R8puKRNJxc
8jB3Ve4R82zqHf/HsvJbgkByYd77e5tTKnFwpFIDdEYioHS0SmaxMbX8u/6caDPLMtc98WkKRO7b
rLtRXnU2h4elQZtuv+cAAm8caq3KXiJn0nHJx+rFmsGq9knEmjPFJXvSlLmj39wGr93CeujpLnbJ
i5/xeKOS05whbXeFgL9jRnkPwip2JwNTlU5wWUfcu7415WhNjKSWhpGGP0sozL+wKtBM/Bd2xIKn
1GDipcjD6Xd7lc8D+3WhjEpc+gqrRz7prSzAdxSSWpscycZdV1INugCeqroBVYuETY9y3LkpfmB+
0ulbZoWzkQcQ5H5ZsbJalST88Ycoo0ypGmodS03ZGuWukzP8pAjvlqWXv1ehhXDhqRMlTp+r+Uav
vLiKzLXLA4eX8FZZ/IS51BsE5LFwyZAjRz69moF+ny0FGhJ8h6EbOhw5g2R8IZoGMbGq9ABsWiBI
iSihLqiYvEmiMW0+K0wdyx0EAdLpt6KVPf8eNZb1MOexLWrDVT1o93R00U1t8oRnQitJFD7O3sDf
N9X6CgVEKaRtZ9zaw7XCgRPJEwwh0aUyVFb2q9/FTuo3F3xAHDoU16hpvr1rm1+aYHXyA450eHWR
lbGZdz6e1aLWFPagG0MowJ5d/fuUAJ/v7iWW6PpxoxwokmhZIj1JRSoBlmUODfpU87JaZ8HZYlgj
sEwDo/Hye74cY2xYVC7LAjKHp2z5Saicy9sAzFwLaMFXx3SrScHd01sw5zsCBSsOU7c0HJ1XCyJj
Zzhmpp5DbXcDqJclhsTsoGHtuvyQvrYIprkTIWlO/JtEJJgPvsbFQtLuikbJ4Fs4XcUcfnUrygYG
ovig/IylaCKbekcIS4t0rDcuam8L8I8ajoyUNwQfbXvewAKVSdZ/lK06mVYyMn2A+ZHwfQcVqhel
aGxC5xY8lsZHmPNJMg9c7HE8WU1oLZlBy6k1qgoImc77QgVjOG0knuZWtAlFHvoyobvpJDEw4Y/5
2Vdj7OXssMAnjWd4cJhIok6mroJr9sDhEUTwcnBqc7B0xppXV9VM5Ut8Azf/kLzb1MuqhwM3A/lE
zW16uU7Y9QJRVq4sDh5byvedkPX7QeXMrKwjl3i5iQegrrOulJxZhNVhwIR6pIGOpqASEwsvtL1E
x9vCZxaUII12WBs1qitRKQL62pd8ilXQNUvB/nU+ruxR7BzvQtkoaBJxvLxiDzR+fktuyYx37GtI
LEbTR7DEOO0g/1x0VthMzEzVA0qhtql6DnT3KoLkbaACR7grVLU5v1YCe5eP1onOZ1JI99xagJkY
/SGPDS734+hk51CyN7e3Wakra8VtDdRGSzg+/Ypkne56DmY4KRWyu79pCMv6yw0pKQF8L6pa1PJi
8AB7DoxhG3kwPFUJs+FnArU4HCzPyiUyEwrKfm3nwJCPRL/v9/X5iVUgYO5c5NKs1O+DczoURIzl
ueC74Zpk9dmNs6tRkYZtXcR8Q3bBfdRXCLPHr2KnsfZeLl9IHRKRaW1o7QwuNTld71T1cz9bbsXL
wcwtN2r5SXGeypUQFk1DgeBKBxwVHp/BahU/qH3yFPr1AUyWxt9QqPWTAuRbaVJC664/c52HvCVd
X3S+y5UTl080I0+8Lvn5Rcc+d9SMwqR+c5Rg+VIcVcK5ZXH1kc9s7Mycg08hrpXQGeHc2nisGhlx
CyOp1z5RaParsei/pZo6tY+MYuv6K0zg1yrW2XMmeT11N+VkR7rvNlLSRR0WnYJyVzONSgj2xWnq
49tmvukvnOuXkoAbv1adc5IJpMypGh1+w47zA9Ysjmsv10f9ML4XRybriNPSIXt0r/YWoFUSfONt
E6HPIKMEmftHZbhMczR7BeXNP4gcHqpHp2gx7/qwpL608F/h5wuxIj0dUyiTRpZMO+5FFnmRG9+x
l+eF83Vf4M8zIOkW64v1Lk9C8ztuAK8PYsKLFFEhZK/XKwLEVRQGjrLDD1D1en/2fv6bac6jMZ8s
F0mx78a19xhUYbFzIBLqVt0FSKPwkCiT0/LJO6V6SUXq1NozVVOyC2dwbG5LPFdgS2wfSSyg6mwS
UtCwCtle93SeseDel0F3Y1/jF6ykOiBa/ferOK6ckYJPb23xsSTlZWZRQdrYUb2T9sDUi2TYYD82
GxjtdrKoEkyCJCNq/x+OMFuEpPEddoaPsSQXyzkgHMpndiMTmjdZNlpTZGSEp6kpQMWcEkhNMDgp
HMYliFEzs5mHWEfQLQpvNrWd/UJsqppBXrfS+at+TL2pozwEukJHwZ3dncwCJrkAycKEEY36VAlE
PgIQMasmWDDd6VX/6ZKYMoIKXv0uqqbHQIuAOIkycN1v9A0UK+6NBkrWuhv/YRJq7PDvlzFnqdLF
UXTveXTgOy/BObUTLnJqulDhSTG7Zj2+TwzTzGfnTABeTbBqdmSsMFTQUW1wr+DQP/pjq1gTCl/h
gV69yKFyNOOUF4KQA87HWzPY73uQJWBie34QvNwWejzy4IhQ9W4xfuEgtoDrY1PMZlmr10AzaaoI
N0xaSvSjRF2mG3QoUMcQsGCmScmoeKthswHvNwSdb8Gw91shX9l+Dr29l8rHt5AnHRI1hNbnU7xV
Mp3+Pw/dXmCLomuwTUvuuOGuIXxcKd/q6hgNdBJj4fYaDViqGgqRLywSSvS1/f7L6uqWukQrLtif
6DUHEffbnxNKL+utVb/D+IfL4BFkVfF3NvN97uNpLZKUY42orppESIK/q55rYjShFL7o5Wrh+R5O
zrmODA2o/ilHdNhcW+cmFnjBm/8AcnsqH5hZIKXO/2fXGLmdOxu24Fz3vg/GvM1HkJ+ZDV9v/73Q
cEXBnCtuTgs1UKqLCp8uRQhH75vUSP/10Ye+zHyP/xKqCHi9X+EZiFeLSOgrYFAelVGHWATjMlRe
j6D89T1tx6XGmAo78Oda1f51mb19e5QJabgsrW7T3WcyLhYeUqtVt2cBiHYCiiZdzneEzZvBXyMR
QPK65tOAvzhlWjypsg5s/OqpCG4sYWHwAgSFO02LCXCcGjoEPk9nHyUY5+xrak49Qp1cOgKIy85H
ZiL+CXWKaNYnNU+UroREhELQZo+aJHOsvmO9FXa02PCmBPfGn2dRag7IDyIEAKvKVPKUN4AvGo3O
bsgmWZhEUxrzakZcwDe01kIokUS8z4cb1bhae7TQ3QZZOUSYei/sOCs9qvlCrlK8KICUJUcCOg0P
JrfeP0DtZYcaJFchtIy5Vi34in3mMg5FF+qQwqrZWjs/GblhOforF42PeAYXdWdvVPoEwyTvbGOo
Mj9MQFJb3/1V+0j+15lujGagcEKYBc+Kfv3FMwkNFjc9wOGLNqTpFu3Vdk25NcL8d0hojYntXfLD
sOkbEyXvMPEefSR1mMRLJ5+PemE79OmxhsYLZuSMfopbbuqL9TEIPzMuqkjBFRhLnX51vDrV9TPU
7oz2GDTCPyVPrSU/5e0v0I11nYL8ByNvy4OfW67drFbP0ZxlwK7jU6ZEnjnzEWiwXcbc29Tnd6uN
CkNtiZJud+0VTPc4L41f7PKfNtNxeNAjLkZDnzud7Rxkza3ZZuvmsAT70GnVwVqTdUGLKlV2WpME
6gIii5q4vXSmXIPtR7GCR8mF/YEMg1ZDge8rp1lKOIiJPQxjGEVAkNZvyhcKHZia6Mm+DOhRSMlv
3LoJrIYETutdFFfLqzlTeLCJ1I45YryGm5ub8IoJZ+E7mr5VEGfJBwjUWyJZmf2ahY0J69g77ulY
qmmVSQIXxkcW6aULBobV9ZL+TZR3FPEN3ojMLvR+bjWxx7DWCB2JO+JVA3q3yh1iTRheMv489FM/
GtCu+8kzJOHf6BQ16I0VgArnmy5cryBTPxMRiVXLq2eKOExPLpsAdmv1SSTM/Inb/9RLqK2Y/W40
ggVcHV7g9NcpOQbVvdBC6OYzvOxADU7ptzAt6370x3/ILvNnxUUNz7mOnIuIY0GaaobwehQ8DvJC
txqMjbVpnL/527lfvsunupvWAzeFL4d33wTWRZ5dkxDzAWb3ElVBI1Py0caxTEcSLmobt+/GQK6k
dKQP/smXaFVoaHricrHW3MmOuWvFDbY5nds6VXADS2tVucbZSuuACGD/MHjvAdzlYKW09F/6/Tz0
M1kqhGM1bHQ/rS/cGoCZ5HHx2jF6mIG5Qg4CXgNR0MDOAPfS75ejpgDBUMSmWO3qZy09eDzpLIPA
j1jIu9R4r6TNpzMRELaqq03EnVd/+3j4N4PaDqeZsTL/1aXlek1SaOZY9uTv8nisC44gvShl33SG
tkDJykwjbZp2l0V2wYUFoPFtLCJHoewvaf3Vf/GAC4tpDnL782WgQhoAUxZVKtkrbi8huDObfbpz
xOaBVtrGS/FU2g7wgqvaeGJlz78/L9AEzzJtcf092xwiT1yQbUDFhAF8OVDAUj2Qyq9LDNGKZNKY
RbpMRYc7hzMM3LNT1g0iXUk0fi2/E9u/p//v9bzVVw78whycZSGO2ods4+EG3WCtXbz8sxpsaoox
N5URGqQcCroktHsyS4BGPpZ8bsqoPW1KIOTeJYIZKt/MfO9UzNvlQUNwLf6dgUQRaXvVwFPFNs3h
k/JtsWPO4HOb2WxKSpqujQ201aR/7bkiACYXe0T/lZVUGz691mFX3jOxUf9529A3H49ZvMchxdpY
3Dx91b77+EV811R9/7drtgR+PL5XM+ihv2Y+cX0Axjf1D+KoT0qe6YKvQ7LwpeyK9VoyJ/gqXv/e
sU2svUxfEX7Wp6FWszIydfvRlhL19IyoB8mMfPMl4FTG7m/ujpT37qxzfqE9DsnRz76XfvvY5yco
HT46d/+5sbBrWg3jTI0ezPaw4fa8CAByygBq+6OR/ZgDjMafOM5XOPxdjXWr8jMnhj6ApuN6Zyub
YAvBCsZNWoid03mML4fI59X7yDJ4bBcc7CQZM7tupwv7s2HNLrgBUxqrFhhEqoNyLhoRbnzqIvTM
rfX2F0Sns9zYmTQjcY/Gff+x63jbRhnkskYrvbXzu/gauV5sV8ReXqiG3kuVG3it1hHfK6gVc9jk
mmO7FlBfphb/LLX9AgAHoZy2YuUrcWlkChVNpz4B/39wjHBtzE8/XXvEJIf9EuJ9LqN0hxv4++2D
Q+HI/XkAGSTc7tHYS2GvQeb6Q4PDmvldbpfeqMR9Dhen+70yam0apZetSDAZvzPDloPoKpr9uJtI
cferZ5xgW0SwxHONosMfImwkgNsJXcu3vPmFtHjsd5fyODECFxzXCa+rCUsz6SpRVXMCXZUyHtUS
lIBTFta55oAk23Mz0NDKo26gLyO7E4fz73xRA9VCwDexZLJgpBDKlqRjnKoO891qRtOfk04Yg4PR
8PvXqWwBlnwQ0NwXeaP+IykLCHQHo75Rv7pNe/bqsurLtCJ8auaS5PXP2rM+JvKTtB/qSzWe+rBG
400Ae4/fsn/yRytQJgpWdqHnrND2Rc9UaEztt0Nhn5+KmCeLfHzN7xXRf+kYiBXBg5i+GBKViRuG
X/D82T0Rx9rvwLFSneeVPllYqTXW3ze44apNpzH/s2LbGNgXSaaP5WDzMKyMU1oRrusSymVOL+2Z
GYtNwfZo9VX7qDUzVe//4ZPlgCbWdEtybilc6aIhmbg+dudKO8kqQXjYZExaB48fSQ3r7LHi/IDI
QRFUjKGxtITL7eap0/KDBB+U6wkcCyt3ugR5T45D94UbN4x7yAmyrbnHPY2gmXOSuxof8fbdOBMy
3GGYdhPwKx7MIC5KdKgZ2DJwn7UltwjkrWgUZpYKCr8N+6tog56hK+cyr5cSzvyI7TxuuqbergQV
+mWcgvNjBUIPGvwNTq6pWzj8KW4urepSw6n3JEjDskjksgU10K/Go5fleRVDpxWGFT4c07KabVgk
jA8JSrEYcCpVHSNQbVHxcaOjewzZvERDyB4j+cJJaPFKnOfPPuJu2HlrW3IW7SFcynoXkM4us9Xi
C4ZjXHu0eBERfxD0RMJcOY8MkXTRb3zphokWazGn1l7qBc3BzGffkNJft4ecLdGc3cVVI91FK3hm
mDO1Sgf3uFInwbEXYtt8fZhO44KzKKvpkvfpxd5e76IifYWe39Cgc74hlu/nAQeQ2CfP7Na5iq1D
h8Di9sfOx2owcd5atusoaZt/+hP55mgbl2nIglXH2KBlWJp0snyYGpK9Glk2w53etTp2/8I8SYvc
VefNgtj8NaxJ2/iMo4z7/Lk8udynPjvdiJ4LavTqObu2a/XAemIZkNYZaloTcd20qivBmGCX0u5r
GySITwFEN4fiKJ2b/y9EqxfnjTpb+B+AjbcN5o2KuV8WhpxZ6PZBhAnHxMUWjWzZp3sNc9aEup7G
aK9o3Fwxfn6jTXL6IUQe1xTACJQ4ylXWnH5XPdOjx7BAIMcjGU21c39kUbvqO5K44CvRz306AGMB
GTctk4/bD9Ib9oyPIrNo0y8LyeehXvXPlnMY2FiRKQbIiWDrks9M9qFzQ1WpHcnhuAiEOasnYH8a
45E6dgdGrYvsbTpbMMX3igiyvwtuEPTm70Warzm85Wz9KLHEE7hwdRwTQRUqOcIuxailzhLRJPm3
sBsIXpdC48vYCkRnqYJQAnrg4DEBRUe5OuS7e8LIUC5p+2hy1NtwOejTNokXv1Q5HbhCuz/UfM4S
T1LBk2B713mtFTjzP7Tj4Xno9Z+28dF1eV8SrhqHutu5JAPYgXWJAc5PGAWP5MqJdHHPUYIldF6t
yjWzcRBjzgFJk03W2S+D1jLoqXAtM3xq/zQsqYgEXlT9UWlKQnQ/XuFt7QEhLcsIjyzxhJSvHw9Q
0D2/iBdE+9xaW+9pFjQ4xgpbPvQJgc9RwBBr+hARyRznSKQ5aU/uPcoM1C3ssQUokSduiZO8/orA
errEVJRmDXfkbWLLrda5ntxFkodsZD0ZiyuGahizF4/LHZnWl3zVF4CJ3kyzO+psJfHwra+UkdV1
MgAGr2EAiWqpiniq03I2Tyki5OQ2y7aW1ibhkQ55LfryITcf2zdKYA8d1MmtAXiXidH3coLo7Btv
vFs5RVZBeK42egndbSj5Z2LovoiJTbJtC8k0vmP5mQmM39yoSKwGxE5TmLaE98qu2kPAPFZNQ0IK
E/hYLUOBwJAaqG5pB0gAx4BdwdkpSbvJZi99V27HhIU6jzniBo7PaUWTup/eWRVt7EpJl980Je+q
KOFxwAJUfq9lSPWv7lchvVcK6ZEyEi+iW0Iza+Mxw6tUkLYCw8DWSaFpsQ6aXOA71DTk48W0J8XJ
rFFEGDksp78hQVS/lzrJHikR/TGDDLg59lmHd0GISp1/9c0xvrmYDOHO5GkJG1+2ErfxdBFhKGj0
iFOka3EvubawDfcEZNI04MK6zE1PLY6CD5mWr+/5a53OuNy3q1TgA+YmT+h3AZYxOWCC+zGUfWq3
Fz29m4kOVN9IZPBEj9kLGfmuraKTuTRvDGEp+8pLcY+pxoeKVd5tAH7Yv7kQJeSac6knppe0dYgp
QwQMlr71xyVawbru6yQZFvWMzfaW7ZdVx/NOz371RuZmvdy8L7voRe+qpsoxWeARJC/grbdThwoA
hLIoC0NxhnU+U/yl+cRObtCFdXrz+os3rKPZoUdTDsIsVU14wKtfFX6O0pPzkEw+lPtWBCr+4nhj
RoeEllhIXV7mzhDTf02jFnSuchsstPoDqVsv11Exg+0rcb/uHvrt+uDd+tfdRZFV+584o2Yi3qRl
8x1dOaUieSQ447rEzr72SVveJF7T2u2cZQxeQ2prKuxXMjsEPtCi0a+uJT3om0YDriEoaDcgeKLS
tknfMkFudiAtZpgwb8rXb3b4hZ2zESjjQSXlYcJEUXEyrZtzrmXiC3sGGljRj5ScY+bg7YhA1zWn
jFvv6O26Shc+uDaQ4zUgDsCJ6zXdrwCd+9w2zSu6g9NzQm0zf2gU534ws8l9nBWznePRaJKxktzw
0ZoaTa7TVpSe4SX6nDogkmnxcS409xo3feZwp7FP8aa5+Eb5MyWY2rvRhu9Sz3SS271BAy9E1C3c
P5aX40IcjYl9U2VGyi0TKXUmsY61XH8NWmuIkChz0nRUSlQbkg6SuPr3lNCKD0KBQMELyLXhw0kV
U4gBuM64/tDMggRqAitUaelqDTRKfTAsqMbkL7WTgwl7ci5zn8gQ0RCehbAAW/osvfgq5GzyZGqo
J3VvatAlORNOokncHv6vh8fqhCeOU/FOX5tF7B7bfgLaSWEDOYlJT6Bpdl6XEzoYugQQn614XZsY
IwUX0CcT0z5ofCmodcISP7RGv6RWbksJOh2OB6bgD5GdZp4YwHvHbcy/0NMa+X6W5ge8aGaMnDLL
pZ44y0duzmRPfgbtarXNybfXKBiL7z+vDV2aFsyoahTSqGMebZzVe7LYYbfG1iHfXdJtjqNRSP74
G5g3OGifXPStutjmflq10t3olCmuntb1j65drG3QIaudCuiw9C/3uISA7X1jzyiHDQNCmFJuLlic
F5hVudYlvkXHUCFRAh812LHXOSW9Q9uvnuKrufRcVtWjshUaxJBQl3XjgwsaM/p3gUT9eE6NSwFT
YfOG3IXNIoZktHkp1jO42KDGGHDzA7ph7C72o5Ck4CckoYC4jBLrZZkkTFRC5fbzkdaBpshh+coe
wfBJOwhxLd1uLDGD1wqiUiRDvR32zvW3j2CHtzYB3XOripqPWHQqTxXALHUZHuhbMtPa8+0wdxsY
eJFobDB+fGTubhw2iQWBVIpIw/vNPVVFzoRC/Q/hQGniT/y9rlu28ORCsPPzckOsMDHTTD4T8y/E
AusbLiYIG1d38X4GedXLeaHpa3sxekM6igXIg6x/7E6gKGYEBwyI5ffGKV+IbjBj740YUdfEHMg2
V2mdLQ30vquRFIK+wmPB9Gu2e5MqAdqfbGFdpo/GLOBDhIqcP0CDpXUeAbrUH0LXtN1MjWtI30G8
XpvOYZqEEzrYRyy89ni9FS7Qlx1PgvTuJxmug+EwzC8RA9YLuf0dvZb5V8OknGWilhHvbpl3+cEP
3vAz/DxYAZbxb8Ic2LLXwHqaIo9H35yGRmQYzGG9HPS2On+Rt+D1Ol8E1lKIsRq8ku3GpCBtbsKs
lbvuVIuD+UamNvYjn75I8hFb936nWlNSn8G7/Dhx19soIemEqPrwXGxsD0zIJO74Bc00idaB1rdp
9jN2Nnw6QJ3lGaUtCxX0XVhb+bpfYx8cKvX5fjXOxN5q2/J1I/QbUTqxx/ayyD19rbZkovI+7N2+
QrxKjh2FIqoLUjVuHaBgk4wom/nZlMJUpuDDqABntdXlBnVp5/Nwc4rylZyqS0zKaAhhzAIb/qUK
mZjlpFx8+mVGolZ1DBYG6xXn6LxxgaUyPTL4CIIT7PYTCAjWE9BKX6OMyzjhg+OOlcsjoFiOFA/2
QeVNkq09HOTSD4EBDsb6zGPIWcGypre4iN7HXUC5/3ySPOO9ZDjQKNw39GGiUIJVPrQgLcLO3p7G
P8mNUUlSm0eA1a74GBC3Kv3Jb5oStX9JIm5p4p7uzOO6pciGyxs7vB6Jl+8uDWe4yf2sU1+LrLsJ
2GomChlPYRudQlFrsKJkP9VFwSG5pueW+Zz8vPrjgNL6tJWKsQS9dnHgnPK+c/w6t1oipa6oNpFx
OwR10bRWe0b6biO/spwdFAxuL/jGNn7pA/yvJHumWVKB/2VwJwNOTdc8VQFPW27oPQixjRqLJyF6
VtHW8Ur6V3xNShkQhpIr+B01OMRVJHM5u6TjqZwNCqrpU1UrVe9R7DdpjHKYrsMcK99ubIUt4Woe
ItDocWe6LRAEZozcFm2cftyzx7QE7Ou7I22+FGhL1EeYTvQlCUvyaWb5LpRIXSHYXGvs5Y5O6ZY0
T2jFFpfkY+WlkJhQH+YWytF7Uf5rebQKda2GaosKua3UWnuXNMsv3xd+o6n+97vNo//8RJbeFxCM
VHUCkigJZ/Rv+GityTbBdMSNFYLoBdX072DTOnbwd5dTTGnTjEW+ddqB07tufJT6+O+wMhVh7kdW
eGX50ACz5+hkYLtgNuPq2UG5ZI8jLsoaN28wio666lWvGUsckwJOe3WX/uKxDEtAmRm1n2qOQVk1
g+RcQFzQ7ByjRSA6PrSJOSxhNf3akv0TmZc2v01qx+/F9N4WzydACLrqgTqabuD9gUtDzvBh2/D5
JMny1FS2p3ZQ5K4Y00Nz8/2lzC1wG9yZM8PzDu1v0rE1gJ+iBMC3c6qtpSnYsgHb6Y/AN6CH8S2E
Q0mXlXjbYvSfjusGV1L0BzFfI8/B4lbmSABL2Ge9G7yWynXQiVjjUVdvmUKkxCnYSn8aIJ+44f9u
AuUqwPRuFeHb2uk9vn9f9EtakBNZ4YCTLw3J+OZU/2lWTdF3ajWclHWGjPjiOqHNBeeIt615T7/4
nXDISuyvyzMKSNC/TddZMjRIz5gRzcxwZBXd7aRBnOGFffhmKUsVl+eAvABGbxw9+3FXU6iU84q3
E8OwQ1u5Qo5wqIIV5dJ83RItQ0X7TFpdiSw1zBvXnwp0GTTaCR07U/AEHjhNGVzsIudU/fnYNvlK
a+7F2pxkfO9krFkh6lb/aCuQzimNOOIShgkIZ+hpXEWgJO/OTgZNTNF4sShUdATQDF+NwH22YOi1
5iKttWASPMquzmSUcT+kwP91k08g3c/8oDVhliKu9Pz7B5c2dkR/ffmd577MrF0Q4pKQqvEuHQLp
WEDNrNqXUICyy3KvALHT/vmjnD6ExCiIJxsF17jOSQmTYMataq4ArqQv9oPypWnBGAEROuxKkWyQ
Eoy0fKXMxLIvDFfQMKyjOcLBKj5XIFP3Z1TbxQ3h1v4aJe/Mjp5ph37XRA4Uw8x1GgLK5RuI2Eup
LMaHBQK9lnv1FSmu12jqPFQdavo/r8ygR9j2cU8Xl460adtYxueW89y1gEhl7Dl5j7QtWJ5nOThC
oLwzhNPy7PODaFmpg+LT/tt3SLWNj29vpYHV+h3CKREnhQccj2pDcfkkVwSKgidSWbreTfINyi+o
xdRzI/PRE8Inhxfxu686Df/Dv+CuVFwsiW6PXtzkDsJ/alAVrEjZcsovizPrgflafL2/7yMRxuFz
bhR/atUjts8J8Xql0jdzZvJKVaRnvr/NnnApkHl79utuI/MOKObZe37Nv0aatTsZrqWXF/P+B40s
o19wNHsXhbc/c0VJYu434goXzyIpshhKCnFa4qLM669Q/Igra0tzjBh7DNGL807/DxJJEZulccUB
Kyib7j8YBuPdSnsbx1i9DZQMm4GjV4DPN8jINHhSn/2TY3wUh4zYEUidgCKDFZfXf2vlbf5dDEV+
EbgaYRnaKgRHkmXeAhWSJxjEXaFX2VGvq/xkwPt2oTQgOO8UsRguybtEHp9xMUVC0FwJw1hVzttO
TC3RuItS8w6qT6n+nRIOvevZ4IxJOeig+V3gOAHZX5EHPpi0P0mb296o2bcBfGIC+zqxuRNbzaTQ
7Vi69RpZuzY7Wx4SrLmB2yB1Zs2ryMyoHhvkRF/UHRJsueODslYBA/bbLjm6MQf4z8xZgn3Pyup4
7Xzfl4TpepLW694eT+r+UJ6AIld9ioGMY25ZKMqG9qkGGOessZXrLDuX4X3QV/i6NHn0b8W0C/5I
cunStRdnCAjfjw/bMp2GpAhuhh4XiStcj4j4C9jRIF3fWutGBz+t//5H79uOe+9+IW5rSdi9iOM6
+07najKJniUXb1wLpeHfiMVuGZzjxf4Sw9kQ46JHH/ASd0L7mgZ9K6Z0HuAsEokCP7y0Btiyk1DO
a78jx6Ml4Y0und3WP13KzS2dA/vLeFROBwnq2TVPyr7PScd4Mc6beIeTFz8AVftdymjiaJc2jU9X
dNjIz5N7KqeMyusDkAFqZ9VL5rcSxQPiNj6fVyiO98Ptv+9egwyZ8iGBBPGmyx0nXgpum8DxAUiu
XEC82ARxVWcsrUxBlz1vXtyjTocprLzjkA/DkNOAGh9bXWd80AnW99eVs7DzSKSl2cm7McMIrBAF
QG8Oftb2t+83HMgTVaKy0bK1Go0fr4nJvUN2+xAh3CJCtefyjosykVfv4YYLEW3QU1V4TxcxS5YB
XJ6sAZM5SS2BjHeDbT6ob+m0zgWxdtRupvJ63fwaufaNv9x+O5uhXal0wwyPcbDC6/3S6jfp3hXy
jSXY2kUNBvcOeU50bAxqEdRqbwUrZYjOwrhpD0bJi0hT0yyCkPrRMw6rLutrQnwyiLu+c5UgJwx6
FBpn49c4zRmjIX8XRgv77CCIpnxTrxQWDDfk/9Sr4lUAds6lhuo+air86lMBb53h8eRp3+Ysccm8
7tb2nKd0jBjDtNNCnXMVqEsnbUZah//d3OFYRH7YFU9ree3+FlPHnVRZ9mysOycSCbhv2NK47p9I
TPDPFijErF1CMX9KInyk98/0ZKNQPwC18vy9YJFnDI1OOcwomI0CszTXGroXazwZL+glSEEIvnjJ
uQefGgwffaMdkDbJibMUN/gEkfzyvES+K0pbya42gsy7g4PN83q/3x8PKn69xkYXK6D3OswQm8pO
NavAlVvsxur0EHTJbbf0/q9ZEXyrfOZQJh4w+EzNI37vlGJwNFlmOtXOYrzFMim5iddkK8Hn/o/U
JZk+JoduLAA8DG3JLu18v3sHrdTpmRfP4P0iVdJNfETtc5609u2rFND1D6B+QfVkzA/iHIvGVmIe
PBdl0fXh7QQksT6hcRyv7wCkqfZQqPNf8KUg+F3am+3PD5kKWFBc9ScfAZX/bzFogXrIB1A6a6pf
2azmzeA3AzkPXX86f/t2mgsJOO5STtNxcGzkP2+sMW2gGK382UZjpKCB2kvsfIBP5skS2lFSKfLe
D9Nz6aV1tcYlaT5KsmBpnigRTnhXkyoIxcmyfVxPsv/Da6WD3bD7JMdDEQt8h8SqN9FGdl6aEDkZ
Yx41Bjb3CNiMg8ZmbUv/Gc1xABZzWRhOrZf/tTTasKFqo+HzfwO6O77P9jWkJTv4m4mI7clONyZ2
POQBhj5V3EUasgno+hbG3aUxrHnulRXupx2XhpuDlZ8hViYYN1a2krGEDOZ/UuNWoM12h/3gYhMF
1YqOFoiO33D+IX/82SPoUpk3cJILoTEjDrwr0sLmSnYQc3Xz0XkcXfhSf7kYugdp+9u0g97bP7/4
py43Bmg78/tGfOgO9ewgCGeVikIlm6htX7ewDqKqrzFdxy1cWkAEl+FwmvS2hO/LeaT4+1VmUkJE
Jjh+xO9Gl+DSZSXC9jN7iDD4mCYBs51ktEFvbiE08QdhJTHHd89rUnjkMGNZYkyd0TyePYYRNAB/
QBunumUGKJkhMtbIO6qfJLlxoR7Fq8uUIV/Z4nmzWMVXOZ3F29EhcXsToxNCg/uZPJkF6kpwbsO7
gOvyqd+AQvGNCcQ2EEXUlcAvBUjoCE33hp4YqA9CqZYOz78Kkr5lL6rF0MG6/PaW9OghuS9YosZs
F/Z5Vi5knOTQgsKde+NrbH3HxGR15/VSu6PEjMgHaRtFpePFXW8SQLS2CMrwZRCY/3L6BcdFHlnw
Q0V7OoTTc+3zk1o5UaUxbJjFOFNgPwsguOQSeMTK2LCFIlR6ISuDtpF/0TzAlRQ3ZcARcc+b/Ich
yLc50geaFgEjKHE/eYtG/b74uNVlldc7VxnTlMg5knq5v1woN1rxJmYTFg6SBDK0Jwm8EkCLgV+Q
MNjmMbCIZcFPqgpOSl5fnFpH2Jae/oZTY8USM/+OCpBdoaiaWQBE/Nc79SF1yh7bnuCzdePPRXJL
hm/06j99Hu6LIb3WTtuNwn6JqVCg3E95qSEMpT7BM4HFIkRvHRvGR2HYhNMYhmPukL6FtdjO+azm
Twb1wygo+YvzQyoptTnAmC0eptMazSgbqmSQPDycEiszAY/wx7bfeAtogqfKzUSgS8xsV8SaoWm0
KphD2SHvwyRmhfr9Z0/IpZMn0W6iXYcyeS8lLr1m/7fgmPUNL1XxMqgJOvI067BxrCbmnvbwvyvy
v/Qq0B3AEkSiuFIrUVOxzZ1J/6egzOLn8pacecMDAlgKCggYXQimmMJM/lg+Tu0zb5CVG5OSfyVS
QpwRT4AO4j/KF2yM5Cbqq+2KIXat011Y1gDGl3JqORX9iHHLGCRewv7NhaSkt+tSqM9EDHQtD38r
NxeS6wIoyURpMQ0bC+LLRZ3/EhhUcOljlDDSViHjaZY7rPdxPOBVWQBxC5OCDtxOjaw5uIBc9TQD
FWkiqYLp0OkwjkyBQG9A4zqyrHR/yZ7C0nyPmoI0ShrUK+Ew2vjOaapm9G1za+R1WZksWmYoS9Ux
M8rQ3+DK7Trp6PUhmWCwJ+xRg3jgjQFL5J7reYtSnSB/hMTFgGbx9Yrhw3GuJ3FgQ6enyqOq9Gfa
7lMyXq6JYKoh0xWTw/mhEggM7ioq7rgCwu9WE/f1/uBnf/SL+Uxg8uJMRSxAJG5DtVlA01ULWIEM
vlqylzt2m6CNaKb4905sedtZpecWKSZjB27HwucbPB3476b6cOyceSxDvGE0lsmIG5odCX7aThj5
Avn8GkQCGCY2ZcIwxqgNWeYAZGn0V5EFZZYDvJoKcsN1SoM3fTErBn8AcVBTlxKDhk7bYA9c6Nvb
nFgQu9XwOSQF+CRn6infFB8jOp7HvG5kB0ZxqBnjma+oTOrtkmUPQUdQJCMhv4CfVE2Srjb7P74U
z90opVp396QgJUstpaC4xEizp0cUhST+nUEnXUAFWsAeCrWux7M+Lxi6B2P/S8RpQcWwzxZzCATR
3MfgX61+aECU34vgPeAVMfnPJvUIsHJ4RIukAYRj8s+NvZW8YhxCYrq4DQxbtqHFDm1r2adY8ioj
gU/KGIRfYOFmaDKBdos7jVbnU6+nRlaLaW37gqtYyx5BEiAwQVfQOEjp0nM0TpnjDw/axwEv4h22
m3MsWgE6sjS0P2Zqeq+rm4lrmBTrlob+bMsAS4MIbRjmB8AK05ga3ib/C1y5pEJY3fdcpjdXWOQ8
JN9DGYEVwFTx3kMh0yRr5UohuNOOToh+CcRH1RIasunhQSn3Iwj24y+/Gn3UdIo6F7pEmQC9uqlh
SkTBK/yfRLHSb3ONHFr7nmGN73OZZBj0Wl8+r0LEeLlYVZ82UhdywdTBwmSAPF6eAzt56QWgZdPL
r+T9IiOEfQjC9tejn5uWeamXEicHjZJ+qowg49KPd+RJDDohew1Qu71MXf5CKJhfZTJhSuTpPBm6
kggm2OON3A4TDZNR6vB7HQXqkSvQYLd0HTJ/JBVktqNjLVBIWazCGrn2TUJqks5uXXXEY/aCwL6L
zvkXMSbyEE++8c+J06nJ2OPyYGqfy0SqaXvNCPeFmi+h4m0gfjgGwtNOzitXeOg2ASCGryOIUCVI
uXguTaCWB1BIp+1R30NHyEAbWeP2QIIRSQjAdyq13mqpPfk7evncryhH5vW1VO92Crn3Js8BjOQd
ZcuOyoemgHayn5xXRVVp38I151boh8P3m42ze+m3TIFmbj/fGmiRbJfQ5owo4zlgkE6qYta+CxEk
MP2/bh7bv74Ql75u24Gm3Zjh5fSnnbNxnHtF7ZLDS7qJo8rmOAOeD2VKSgJsnJQAqNGerqFftcXa
vEFJuUj34kiRPuiSwGaPkbJFPWks9W46OBExtkPRd5q7jAmo+0Z0h/1nSO1NQfOKkI/3g8os1Lqn
DsZB/noP/8vq+2hNFsR340kSS4DJr93guFVOfaQNq6OcpGgr3/2iepcsH+zXlnuz30NbQ/fyq8O/
z5U95w1AhCp7nwKaVXXD3zCC6ndkTtvbYgUSsyAE0E5fVtksA2Fb+mYMw7M1xqMfP1Lcot8XGzRE
4C7sm7HtaiTtm4Vm7Es1LK4Su1PSSVnHHATa/1pHZJyEgU303X05QFbwyYvp21B6e4Vh/lRKdIZ/
BHGVrvpYODRE9/EqlUfjtTcsPStSF0tIKG92nyAE360SmHdKsLl/LcrdH7VLgJVTPQdIYfYFlcqt
CwnIzzx6b+g5pE302STUpYZkAznzNxqyLLA22lXOX+lrxxrDEVT8cjf1dxCCQkerunrLTIjfjjDb
NI9h8cjWiMzOSnhQT9tMKphrjjiK262qRXI4rxyEpqJ8THrXfTAwcoob6sl/GH7dtZCL5ed9mM6T
ja380rCoKV7ag1meR67aonJHcOAMg6tpAFniawBNwULQ2bK+Qb5cThGtbPR+kmmgbs+oXX3tGHGN
CBhRd+iUXk/6Em+PPW8TBX65Jk4nytDj7su6jxiEjLdTDkOUS6aTYOhcBJy/17RG9pXpMsl45UUl
8CNMXxLhJhGhtaQF4yoS5NMljvEJKqseuaRJ2BkMtEMtolqnbP/3mReh4Ztb0/kQQcLSU/y8sDc/
bMwlZiUkzhDjrZy8AObBjvGySmKXywfIehzLM2G4K5nS6uFX/muqS521sdZ1izAeaI96vnEQZIPS
fO60Yzt7FMPI5XI3Q4thtVmbtMfwFB76TJFFbVeW96p5Y5NWiNPKbHR+ZKWnpE5AAiKmCCTvJDYz
mxUYYNPRRge0RenHQ5XHBTAYAzDKEtOjH7MiYqgHRkxslrwevQOfxN8xwJQNxcMQ+oWkFEubg1YH
qqAsjwVTjVmmXSK9bK2/QVT1nkbDi2ez7w84ptJN39+yRQ0vAVni4ZCB/JPa34alAhB9kyZshMeP
SUfh2/iJwqH230ANDgp85VBxzHsaeE1uaoQJB4BDDHOqM7UuHqgQ3XETveB5i4ym/iD2Q+MSC9KH
Ukn1zbeE8jWEQmLOLNDFapyIjjJEcZkLFNHUscVJLTC3mzDgDtaO2Ucn0JME9OnT2hLwjxO+C3xO
LKQfhbRkLBYb9W3egjvF7qcUuZjqYZ8k8FbN9+W2NPn8OP3TWkGgfy4Y4RIRGOr+Ggh2ZLuwRmOE
HsfmNRhNWM7SG9ezNOM9LJiN/nzuQ9xWVdKRI0784RnsconmzFRQLYQPvHP7IMbpqT7GR4f2iTYO
grd5MjACEwX18Y6wHjSUmAdEzKaE5GpLr9B4u3h214eUfmSvou/j9+JeRLYTFGJAIbH+GK8pxy4E
ELBpGJKfGZbRs9qKH5lnxsJj5ZFHY971in6h/WL9Tll06N3s61lMH0E6KFZhjTFN8332wNejxPQl
00y8vMDP6wYsv3YyBgx372Rcmpmbg2D6gRV6/W/Lr3dw+BqwZ3vAX2Eq/raO9tlVNEvkRv5eX8zg
qSWk3m92Ea6RS/i+Agiki3tUN8bExqEu94pxUm7A8AFcovU7Yysx03D4IfP4gmIC8A11JT5Yvhdt
FL4GnM1c1HpOfNSvor+dQ3ZnJ+wklCze9F0NmymKn1BYSk7pnA6mTmBUgEa2ZqCQQ57UjxaC2T1d
gl3QY7KUsh4/cZ0Mym+jdoQGSam/QPNUqchbbKRjAIJ3ErzNhEHSs8mI1UmOPHnyPrDQ7BFneVTg
2Zk9JJ16fRZBoPLNrdA2Cc3k9DoWnp0BDLivapazMtpow10y8SlMGOewV22bsNdJJIfGRnYPZLPg
2DKMW1l92ZVrBWYBT9qPzumFJ6KdiXuYFZLySva+Ll/PE10nAEHGOTjOeDv/q4bXE7kjc0fygYJe
TdudGJen0eXVnbPg6O/V1xc1tJUOS7egpHcrsyqexX3Pq3srvd8o3oNI3Qfq7jcN5H32ebmJN1Mi
9jarPSXdOGlV3EDw8md/iUTo0qbFYYFaIfZfwBqdbm7B3uOrhJ/acMURIEKMacpvM+uUSBqxgrnT
9ZE/Foudufv9w/jLI/bFy7pIL98QhOGEGwizrm5qL4yiSJVhv93B69ub2CtwmzJK7ShgA3LvXJwt
ATAfftaeI3xn2mHqD403gdKtR8adV8S5Vdn2chxdO1Sr+m3fmQNdgULeSW+CaZNBZneXW7X1ebrJ
LlLKPFCRieMjZp3IG21bPoaFe1eJdo1JyoVeyg7/gGQ9uwiPP/vglzzTSWT+ilZDfHzCSjEXUUDV
Qum4DcHUW8k2c5WjFC+k1/A8oqESZWe6QrChmaIRN1o9FRW6uspvRQcw0Ily6jyJR4jF0owThgC7
OWzLxQTO6gl3fKCfcwvYZg0d6qPJsuIehzRGFtEAgv/CMMsfYrzzNkpooezBsBIIhawjVG9TpXBL
AZH4jJPDCbICH0H/p2xu1uyjP7g/v43mxP00wRp0BUs5dtNlNvRstDPF66IVn0I5gwL7IfadHXkE
uFD4rQToojqig0x/+vWKI0IE7cXVyAhbiYPiNhg3USilB27Mo58kWyI1A7xwJDX5gt6WhjCqhQym
9eYUWByGCMakyi4Y2w+Qs1XoIpgpK5umO+oRBb68JYrbfwjzuECS9/CMcYnOJJ4eVAN+OhHT1zhb
KwHnYrMrf0XMJzxZ7yT3tysTQ3rCywwtXaNCQq7qt9//eozMflDtKklUw8p6pHrtVdJZ6mbOXmeM
sgi0UUrn/3RzubydUqdb+Fr14Rw21SHRDaJew+J+l2sLZKOvtkti9ol+mr5Rzss6mz9ofKGuU0rk
lZp+0FXd0krwbfv92eQ6WiriBXp75f0Tl2HPlR6F1ucKDq1lMuFjsLlmConbeVoKBnCpOXZv+xmO
DNeurNNxo1PUlVaJrkTLHws6D5/a737zP7hg+4i9iDGatPx72cE3+piyJgYyr7cMsWCXkdluBunv
lJTZt/YgKo/un33ctSi+lUwR1p8l1HTq987HahK/+mmd3w3HHJiNYSWPMKNh2emYbV/A0ZE/tYya
EfSPiG+Yj8NPpE78N/L2mlQywBC9yJrB1aPyth4xyGzdzglCOxbSkMeG3OKvPYKaMk46k7Sbza2t
mOTABILfBtVMCsAtdxg2UYCrnD9T8qjGcu0k+VVQB5VIY+NXe5tOFIzGfSOUzugAUjOjBK/HnjlB
nZRBfS3btJxp8bR5UVfCcKjhHOeLZ/vIGlzmY6I8mencYYnBneWHit8LOD2KwXeMELlI5IdGCwMu
QbxK7j+PVREgTLsqLX1jkfcurp85WqvkmZBUcHfkW8168ONUlnwvS9jKtAM1EVByrwq+OBINYif9
gvbO7qs+nOJve8zMVvcqBD5bwtmQmYzrrVZc35dl+yJTPBOKRMlUhXkO/OIUPW6R0lINn9i3oZGY
d0sz4+itiheGlrAhPW0e6R9FZZyIEOD1+Lr8pGCTjVM3t+XJWmJTuUXd9sklI19OSf2ENZ7af9R0
dnq2KaU0hOeA25m5eel+e0p6Yrj6cvZEgUWapMUrV1cmR9n7JBh+g1HtdjEGvZst40ZbOQe1GBGd
WXVU5UtgXuVn2zMnAvYu/AKmqpthtQzvq4ttjpIpikGsANYg35/oyj3RjLmFSfjKJGjuxkvmB3Y1
zuxmHsWmW/HKWXaNAQT1cciIjCFl5PCX7PF/lROnI6y/R0rEYNGPBcqb0Gt9pAx5tiPEI+DiZqI+
5bxV/48m49YMQpf2W6hkGU2ewBf2OIHZUW3OrkWas6sCaHzzatovIo4UBfmKCvBgk0vQ+H9HLWfQ
nh6g8keIWKcPCb1Ax9r+ntOYhqu4UZfind7KK4KX2wWNMaVMnXxf4htYpY77khX/GBPBvDdTK814
rv46DZ7OrpFvT9Tt1jOF58CQBGXqqJrLNOOw0G3t43KXEoVcCn5l/tdyIrYax3k4uAAATFqA033L
2XyUT12aVHBbCXDfoXUFz/8KCQH4Ss1S9iHzptHeaGjSiAX0xGoEPwPGKadbMBED9XRoYrGwTbUC
ZXmUeEK8ZEmsoNxG5uW63sgNlYhlUvb6TRHWuLQzQA3oKwk7RYPMoxO0tbQhh2pc/xQ1TOZR61op
aGAj0NTWCNCOrXgrmOnQtKAvfFDn9bDGO1fP8UqRh+B9YckhraVCIhTm4sbdujYyByQx+jK99F9R
7hcodRNpbuYUmLxdR3T+dgEUrpjD+qpSAVPd4cgub4mD3MX68BDq2MMX72n0qLeAngrfZ9wKVZjk
P3ALxwaugegldz+fcehQ5QufNFZ6Kl+Ztyl3BbrkOaeWUhCqFCBF4Zzw7+ev5KOthScjjMdyP+ES
RTQieovc+kmWfikZMa4IooRgCjLkH6tYjKAyi68eiqR1B0GJt8u3OiD0eQxDWYq6BR9YSqeINSlp
r5x9oluszPyFygM7c2RKaMl4SMsysyjJQ2pyIghlRt3EHR1maASJdAsthqrOSRHPB/ipMRxgws1J
zoa2RZfXcmCACJug67VfzmdRBDTV32VPmXslAwAT7+adrArA2EJ70+wIn411hcLj/R36XLEOXnpH
qZKDLNhAc35VWoBRRU4YtAmTVl4wWSI821/RJBfEMdfbuzE8syQxXNr9qwAR28V9zdIi2aEGLqHw
Ig0Q8iRKCwFVjfyySS8tZ0l/VOxRl2azDvps1+bNF9XripDkFUiAspULw5ntU+NsbptPBV6ypDBb
x0SQx/wvh4kW+P614jyHJQi2vIo31hwivo5AHQAqHRligPTSU+l3To4a6hPTk+d7FXCOtBD4e+wO
USs70tGCtFyn/OCunZ4/94o6H7d5Vj9OtSjKn5SAKkl3RoMNjMiq83lLN1qA1fh6bX4y7Jd1EWJ+
g/0dvPZ+BvigwQxXclWuAZbf56E7/1za4L4HL8LYi9ewXNSWI+TvUsRxxVTh3IRl/WzTJNgZLDx8
YQD1Gxndz4hgqYhda/mKV7/mTc4KE5QMhCiglvl8BHC8/qgQ6rvMVVt3JtwTlv+smXqPfGroPYkS
GUwc4C1sFz0PPbekAgDG9u+9uintrUUqT6VvEXWgN0pxDycG0SBY7gz/GmYu1xdyioDFDC/VRHJI
ldhJ2mS7SvTjUMIH01Pe2ZupCnwCbrTJO4y5NDQeVBS1N9kKDWgLbOJkoVmZFfR5BoiFqXShguJa
IWaDwtKCecPvuNgh9jlADJLKFY4g8Dmjmw3wn7ulP0poqrE8DwWnkkDhKlIihDo7mOO/MfVVh4Kl
7pzLNgQt0P3nlKkMhTeYYhvlMQ2in2dIPs+EFSmfFPFGTMD7Idm83u6fU+noV5PamfTivsNe0fTi
a1LQx59CLab3DmiW3SolxIwHMtYFGsjjnqSh+K0w3c6z/KckfQd5TWbuuXIUsN6dMtLImemzpKiK
09XqYXgqaXAtkBT1eac09L4hYK5wTTjTg1Dcejls3tRksdGusjPEjx4VOKMTAQzThlceRrqJxWBX
mkGGr80aHjLkYCFbsHPMQdmfMWzSrgpVU5dSt/Vepcivk5wzzv9jN6zp6AHJs1g4NLX3CcQgl8ma
IeFvOeAmiug6Vj/cWK/oyhG6wuM0rUh8TtLg5qxMalnZMTCQGCOsbhuFYdbXX11oiOIKbJ7a/75O
NMJSr90V5vScFCLgInMUNpZ6z+TYtSarWAy2aIDzz1w4iwFmwiQnCjZGvq8EC2IHO/mEWZ4VDzzm
tXZW8dgd58H+4IpMGmFVQfsFVmt7e55Zl2Z44Ci55lFrFcDULPWXA7+VTlWL+8PVmgXgk3BKrr3L
WsLrzIeOK3EN92fe/YL0xnh4kguPI2pMU9gMYJ2p9Zhaxd72+R/tVWFBeU3eSbvgR7zo5GBPZ8M7
CKDCvsFvSLQR1eaTjA+4GVoTURn5nVWR1GItM24Gxd8zodoat/Lp6kSrHGohR/lonf/Hy8iDHUro
9Zygyui7UYs/BSbuXuADRmUM8CV0yC7GBVkmqTJG+VTABwDUoNz2DMdSYKvAH7qkMXy3u7YZyyZh
HKrQm9XjgeO55qeiF1mbpkaRelnbkAkuSZRbLoCC3Nbsbk0woHRlIDdmVWjVPvOlS7W/22G0tSYg
cHNAh5lwKfSYGyL5EaIqGdYEur9L/70VQoX3qHZ78xSie5dITnKBgJG/Lwa+ZMQs65Ma4kSDy4w0
bVa8ypqRgwkBc8uhTRILcCYPMytfmCCDJDlM3m8W78Wk74/T3BA+hg/RS+wt7iC9uw2L9HWJBoBk
tRflXNm1vCtW+fhfO4mwz0jZplsIi86PGwO4+CzJdPTXQKPePDW6yumYLhENoAF6leLdnGuEt/4d
rpUiVo/L+9u2qdQCw6nSlYsLCrk6GCKKOikxL6Ku3uezf7KPqLi0Qepgnqh0Gq20NP1CYioXu2lT
bTDhuto3QnEDKejqXSEAlFxe8M3tYrGaYqJYoWCEcim3qZfXgOJ1tAyHP+Mt6stfF9hEdmhxoFmC
6DjJ1kvq3CqkVRFPxNa+fRBVWuakE1NRA7uw1YEvdZ1znDTVqMqklZ4j8dkh+8wfSqT0rISqrQnV
+OOzhp6yQXYKK5BPlP5DEuWfEF52cBmj0b+Mu6gpApmSrvlc0tzdNgpN7tFsvefDXpJyCInhneQD
L0Nv1j414MJ2ukO2G7mc2T7z/rB2mKbK/to/ZbQDNEoQDDGoAnkrm8dyC+20ahSU+/KnpXoHb5s+
y+qSoJVv0SqccE58CvWVm+4bQbDVjZ5CB01R2gbXnEs9DOSX26QCWwMLSHxLWQv54IcHHps+/MNc
YJu/tM6j67iqV9rmEUybNfv7H2DTkvXqSAK//oWUjFHzYFSKZGD0mvrK4nDIJkzluc5utyuQTw18
N1jLCJSMSQ8KBsav8KNW1pi9BAbkjgsB213rT8iBJ76SdRtrrlJmqr2wbvsVhh3KbHvTY6+JbHMA
WDVos9wuJfJbrw1RAoGHH6MnJRQ13ISUzHQNCFlrOci19j1TSaebZMnih93cTY71Oo96rG/WTF2v
mlNDbNmMIl4cd8l7S4lgtLxn9Ilgfj1Y5FHxCBqVWMNsdQYfZh/iROYaApDaiVSgSLleilfszMEG
UEqAhF3AMvam3ZxplUwToZ+BtRycCEE682iqiydHs90X7iRVvFcyNBMxPyJPSdsrrm8GVlCyUALi
cxR66O3YuqyHtFJ7FJpU0JfPAbNpawWIMpqyMFqVfbrFJbPBVaUGcaEVWSB8lJumO9BQmaSQ0C2k
MqoMOzcygI6tWgTpSt+105AAEqbuMTaOJtuMLFu5XIOPHOJf1/y+s6ogbpjIWTBifb0qq4ZNkCmV
/sCNZXxOI8tc4XnqMLvVAfE2TjZQ+j735LrbMwFWoW0umF4MibMSkEy/Lw+W54H+/pfpqLeXkai0
s51h1upnuuFlpBcA0pY0tNzy2esZlj/7qXY6AzKBCK6eZksKE+ZWAA/kXn+W0V64SYKAj4gwi9Wf
4OVtKkjbrdlejJOx6RPul6WlK13N4IpvQcPiOu7gbPgsdsdaHGtJ+ege0IUWKqMtfrSxPSadgm24
LKiLl98b6oMzhRZq9/DzAkeShGcJQZB133i3VqdR+kIZJurPmxdASzEkMyZE8chahMpYQb1tW2fL
AwhP3QsY12eqh3xwm2GpIFlkc4T1k4QmfbiJ4hdc3vzUpFdkNXx+3aFVqv4dRvrY0Zb6P0pOz9l3
Ut21x8hAdxSEISLW2xW7EFUYmgGoeFxTTv8tdhSL4QJpQkPfLxqd8S0Fm0l97T6+jeJYfEXWxQPJ
DOL29/XbNhebyFRGpVBfGSUGNjhRRxskHygpiiYO80qnZcby9ILsnHlS/4QDAhQSoYpUodF23GFg
42y0h/ju3GnzhEkFSK44m7wowLbHNt43vEbkhldSQ2RJoTFNsslVXloczyRi6VMqr8Ctc+pkWqtz
Z12iOxzLiXw9JBmVKMO4D8Md6ZB3GGQdxCbuAyV5kZxsTY1js0EUdNj//SGPIMsu9+fIc+v7LVsF
By3veCZjorsHI8582fqg/BNbhNbYjHExRi7vEaQ6ErWLk8FU/00TKDHCoA4Fz2BJ4xTlRXL/uGyG
RYSW96NC11gdfDFksOKOmIp35eHP/Fy3StXRD9b4aehdpj/fFEq2rN3PuupTPflUn6ZqI9pYBM1y
7KDFFveGgJB+MyX0TUhr1wMK8tgiSeeEFhkdQg3HObHkl4VayyJOdkJAnyYMDNnco8Xe6Z/xsF7R
A2v22obiAzsS6vRiOvduGBnmrAo5861D0tdP2KCB0ZzzKqEUCu1Yw98ox/hAFVskBn1q6TXdZtRi
55uEkP7a696WMPdvYh951tLhF55I+CpANBKMMUH8pbgWU+nbTQliLUhk62PjhTuJSWUlTm6fr164
cSKthsIqqGOLXVIAEhU0iYMss5wbVJJ9SRVJlGDvCf/S/ACvRxsxHuWbyCY6fR7HLTgy3CJgX5fe
+r1cVhUXHZzj/wgYVOo0Ts0foN2xIkN4zNK+M8+2dQRMbA5U9rTmrUs6Ww0SHk+X68Ak0IAj+S2g
9XZ0Tb34W+Qsyk9TERTTc4Vz++eSoq7Sl9FIWyafpcwrvsi7QokMDjfFwOaSSOrQ2O+VrTcWze+2
NB8bw5efw1qqAN63p2hZzp5TxpBvx1zJvd/CICM2aqBrbnPPDfPMZ6+RdVntvR9iRHwYSU3jOvh4
8TVW0jUjX2ifR0xuc622Cp8890mxSmGMmZnOeeHgQ6IowmsqILL84ne4axjlUp5xJbtGRt05rrPa
X3i+3Ey/KP0ZrIBIJhM4Xeo5FUq5I5NGi0yocFpMSNB6IgFXVuVSI3z3NmY/q5q/aYx0+WEN1D9i
5z82UiOcmy+2Qd0iUVcNMQaJ7Ugtr9Rjs+tTzZXEBkFUKnefdZZymoUg7rgiaCOQ33lEEpo2/a27
dBOV8z/6NQZsbjeDU+UVizhaXWd7j78NITjhm7XL0/UTswNulYK1siZaYdty0GMHjsAoE0/xqoqq
BONQLFdkk0dXIMVaYsguqTy5gCNZYH3oJAlpVHzAB7BFGVXCGALzxd5JzHSWL3SRLZbe0XLVmCH5
grGrfpQCF773rpv7+IBJl+BpFZcd9JsqriaihXwT0I1YYmWxWEuFbu2Xg1DxWrpQd+D1IUhQlswJ
wsOJxjR8EkaAZVxszZFCn39MUXccg5V53sjkqGjesob0FVUrAhcRodk+pCo0xUr19RhniNF0F5lY
gg4p4QroBl0LmAsg9z/byyuvxx8SWoe3sJmhCb/CoP7S0DHznI5J9C7BpwBL1kD57C3Vxpv0+r8y
ve4NtV7KViENkGelrweKJRd+gtV/fR9R+HUcEe6tpW1+MwK2tA70ZhucVUP6QBizRIpa+gYzmIVl
GZEJkA9e/qDh6n+7Pxoynn8fqoVKmx1lrQ/uP4ShyJG2g937oMWBkiwPmOQfFHKuVok73FUUBHqo
+BTC34hri3abQAfet6XAgCgsqZ9gpvdqeII2bD13lyTCCyOKc5TsuSefcB3t6vLD7C0dHrHtMulF
36FndTyrYlmDsPb81tHw6Qs93QypQvJ6cLsAg9ba/nM9MeZvhP1bI1jhwpfHTNMdaGdL6IoI7N9K
EeMqaELm/L3e/uImvLocRrkG+7K3MavmSwtgEk0gOui+Sf/3zgPqd3Tw28lZCl0y4ipwTy8N29gc
BghiT98ZzRp11AWJVKfkonppPGoDVKcPBRrOlVS3UkpiJUD08hhL33DfXv+OwbQalxVH4IwpJCRG
Yh1n75dDpc88pDZDExwBFcrsIoDNBsxl9uNCEEhNrsyXydbXC2m6iAqnvYAs1GrMcWujNx55P/J4
HTlOtEPwFiAOQZRnlEQ2kXAv0m3aLIjHKzIGelfqasiYlqUhUmlxqISAK4UARoz+5Mgvtjmpp9AY
tkxmNdkGh6Gm3fpfCrsX41eQEkbEP7Y78Pgr6woEAHueUVzV4gNB9ET6h4kNNpFILhA8OJWs0SSt
ad0XFgsTl5WT+0yyEH9blDOF0dTPtfpBu8/YZq56MdauNlotL9ZriZM6z7CV9kDDje3zlcvgrxqs
XEjCwsPEPp+SJ0HQ6ZhcUx2GZDULRVmaxSZ+zcc/yYBmy+cVdQzmgRBdIWavTnSOtAggM8Lk5Vbs
Axgm9hwezhFa76Nwn4GosAMpOzlkiTSbSLqwpOs0/+qge+CjUgkwQn8nFDz4EVrl4Xuh977/OuyL
IXJhVH7NAfq3RvzqSQnFEYHYuncvCTfP0BIJi6cxATSC2QEIo5IJR3NDeu1nAEitdxXPXpXVYhnM
bKY8ZG8YQM7srO3AsEhO4mkL44qWDHoawby/t9sCIAHRovd4wr3RiMgfKLEp5VmaM6q3JLrD0Z3t
30VX5g3BNMmEQS7Na7J6fCLU/Gy1WtYXAsTk4dHaafTXTWN26iFMAPhiMLaGX6ViiYMSLhrdOgyN
YSrDOvYrgGrUMFgQnwErcqSQvMmHnkNFj/W7LHMh8d5tk5u2WABIrADE2NY/K+OtgJLCBsr3B7z8
A1vPLkU+AvxOeR+R1/G9/p7/LwUjOhrnbvHMAgrBtv7p2+Lnhqb3R9vkscj0VLGA3GZBEma/fwoG
C8uoM/ALvHNY9jqza+AX23LdAlK2D2UwdBOr0ah2GYBBmCeLYU16RPc3goBh1Sc/MFqE7eKPQyVj
8HJjA8sHIy8lOVigrYMLVM0bv0eqHqt89gD0/wrjB7zGJiESVPlT/vjVCjnu6JVIKXhnqUCOLBP7
XPWvXXZ0UkMifjWFtREE5O2BdP8bDQWoZq4EVAGHkvQGkZwqxvI5p9hOc9n16/DcP9/UVI7apZeU
Mqs9Ue5kOavQQ+KtujxR203GtvOOHpXJnPhy0MwqklvdDj/FN7QGDaqSKk7DeBx+YgsefOBpNKxD
bXHN5xRzygvmltfOFxHCZjyqef3r9GYXb0GzRPBTtUDXJDuUKVvkikssQFaQrBjIBh5H/6Gw4XN1
5wShIcwx3oV81fXuW3MssdCM3OvUtDL7Lk+Fsa1LzIzHbOSrS7QyBag5CMkcpLQiIkxQ7nFsm/GR
jj0xaWiy70pBxCqypgWuBeZuKFB2XMlzBqM5OQ43kMJhHTf5gsLIm+Npfvlrmm23a4jvXznXY4Uh
52WIKng3D3HdY1rSWVCs9kfZ8CIGjOmMoxuKKOlRGXkaUGJGdwjxyxaeNYFashQV4uHmBa4Be37y
yz+KJYNES340PJuz0Zbby/yfAuaXap7iPC/yAGKbH/P2YxMVt/nv/CfQlmIYvZaTjoHKxNDsqEbN
ghyLdbunFoK3KirUmxLbvu1qfuMFiEcNJmv8eDg3CvcwLsQD+NIHaQonvPCdctxXdRwPEMs6MJow
5M8Bb5OLO9vrvvcXkACBBpl0lvagyM1aUhHkmD6kk+Uh08T4xcaBzNZCpPQ9XUMiYnrnEryd3qiP
lvZA+o8BLkOj/cR+axpKliVnD9aWTBdSpzLCeRIkCyhEmmPfXZ13d2HSbLMpomO1KKTiEpn2YGxT
E7rtUOkN+2/raXHEHj1ESS7ALkh8duMCB1khYSA+TQStP0Jk/9MegvgPeyK53wgbznCgGQu5nxsw
fIdoeXdTEy90tfI9SQY5WoYqkahyQgB+xfkqpdbZ6Ha5/72CdmJthcCyr6WKS5c2C8Ivy6+SW94D
RRxt81PQXfJ2bz0R5QTHtxCOZWXh10zyRhB5Pl01hC/8fRr2x6UFcJkz5mjTGzkVhVwwsfmXRCUw
iol914VT63+7fQNovnv2a82jcYaKT82J5rqvWWehATU9AE795/0HAFU3r3jkNzBwGvnvWJLQVm5L
6WzKVvyG73Vq24wBUzu3zLLgv+2x6uni9I/Yan4FMf3NnZnFjVR2z4t5zrRfWoWTHpjhlaS6vliO
HcJSZ5xmLhKATuWSXeRxCllr6qp/2yL3sppVwaqdw6BXjWZv0nMNW2FwLxBaI4v6RRBjYjsqQ4S4
Pu3YgF+u8zf9H1D1XKiEjNpptyS12pOQaMy2JCD4EVMzq626GPPY+KvH8HH2L2cOqRkp0+kK9LnP
oM9q1ym1mB+DkIoDAckkjOiZr3ehS6Fe/0yZGXfr0Vsi0TA1SXn+S8JHsqUte7sr0M76PGz/pvRh
m0sg4zcBOHY2bnqCC5JC/uYtrl/6Fuf2DD7CXWPsPh3b6RB7ydFGgsIfOtlu2PsNlFgOCOwOSC4Y
VxkV9GlSW9SNueo73f42EDAt57FjSdR87E64jaXCADeDgtxNEErSKwFMEgvQfku1DYVfADiDU4QM
lnsptdnqnxzMffzwJbvuXpxn0yRPgbQuzipsItP1LlsuWekyvzZJA36NWPb+mCLbJxA7uq+u12Qi
a0uMwWRMJhjfwUXXqAzaGO/sDhP4uP6RzKgQG2U+OOa0z3AzwkwmMIZUgknif4zbEU+WErlAUbWG
yI7hig/ZK7a2K4BAj3EIH/eHrMzq9bIOYJW+0CJn9z8pSw2NNTVqC3PBvm4Z2/nTFggV9HzJuAsA
Abbex3JkmBXMw49yGtSHz1oS7pSQAd6P0HQLJdaZprEIqMAVTfl8s4Io0L6B1rumc+s6Ha7Mxwni
8I6z3H6LtLn8tOwTLw1kYsjtHFDEXamNigqdUAV2yrQh2WBtBjLAfOCPhFIZvsAGMHm8rcHZG6+g
8Kw4EZybs3fc6DSsyD8GhF03LSdmwVaQ08MQ7+EUvp/h6bXO/KsaeVBTRGiB0DFaZYrjEGF0wTGj
YTMp9p0K0RLoz6cR2s/UeBZxq5ZGEjtTvorf54XbkAx3CGEvYj5s6TfzdOukEZ1tx3dg7GAi7TIN
pcsAJkX0SfEH5Et+1nzwyzvKjf+E+8XnQWKdb0xb/7hHiOTggYrd093d/1fAYe5F7EG+ZlBllTl8
TluFLSDTl1o+yUHbMNj9I/g/CWdsnhlMBCG5qSSzs9T2HubxSYR+ZU0/k7UrfpNpciCAMdDmBl+E
ppu+tIXATeaf7csZrWme5r1DDmTKVCiSb5h3gLmaPINojpnylIf4cqjAhS777p6VWL7qg/ITMdZ2
c7bia7HYfN6jrO7Jmhla/+wjtu/6MG8tATUt6JuTj6pKTXZCOKHqn+x1mJ4iNfgE0eTeTciCZFLl
HHaERx6AvCrGBladszLhVDLzK9oj8AVgZZUMoGoZLsUd5nZInjWin3DRBJAhF4mMomU+xUQaXWZG
YAww9IYwhhM5BMzad/zgO05lwCGzzTyGRSM7Akbfn1ifSjjr9dbUnc76GAy1AeWYBq6cTWXDhwD8
a8FBuOxCMQBuIOA+EvaltYWArloTSefNTOaRDAiroButrYUSogdEWNoLyukDIb9t9UQEhuR9vsBK
qxHFMurG306Q92Zmi7IgWqG3IY0ru7G6X6hDKSnW3i9u0PFLe9Iux8kYh06AdlH9Dz1RZ/1Y1TDW
FS1LP4BM7Nv1jWkRR/sqX1pHF3duYcBrCopdS83JPHnXBrfKM/6AbXYYrH4exblycADsoEuyuuyG
LgoVWBez5dT2ejPMrgxckMTPlkhDceI7hYRFqip9ds3H8tg9+ewfVhtmc+FH7xEJE+Gr8vu2sk+C
5W9S+HCn7YO4BGJwOKh/RbeflO8FIMLzH4Fg6P86ossNNZJSNGPm86qytUEx1xyW5NeP63MZRDjw
iMs2fA/0Q0rBHwWO4QhdikyQHO4izQOscKFnVTcV5CnPvleMr6bjCQ//Ia515tFBqSltI+TFVWAv
rehz7xy9gkBRExwBO8Amwvc9rR2SalkAE9KHlvX6UhRfT3EkkuZqeIHW98Ga6cJY7I8f4YJ/ffi7
DHR7AHKjDdefBrPoXdjG8ewX4pMXmGDIoPsvz1Pt0biZ1iNAw6kv9wVUJU9V0HzMIrs/CBuC/827
tymaPIUpDRj1Hm/JOR+l5R+POwzD3mFG5MYZW5hFAlNCgMgR5egWBSUgWlRvb1r4XkxE3EWrU6ec
z14/GXCPfsvOD49V01Kva5cck2jnnaLdf3Z3DcWnxYyQU85wkAnHM6yWN0UqUTBRQwC1M9pvuDpP
KlNjkzk2EhDASgHd5IHuyvwBwI095mCGL8tMG9deYtb5s+uDtbIN4WQqlgJNntKLKiDkGtMdzs2c
eIaJEGKVpJOfL8mBraNAqDRIA3bFo5K3flm4M8hVwdy+iQVK0ZXQr9QHHicDB6urJlgldSYZ2UeA
hbSar/cVYqNlJIMkx/zv/W1qs99AqIRDgznIXDsJKM2KEWsvp6FgVRU+Pp0xW4MwnzBWhxfbQWxq
jUe78pe1aL1hDBOD9aWIO8wXH1ZKVU6+BojcE3TOAts/oeRkf9nkDAwietEcg5yLUv95ngcXh8sP
IcfXjK9xumnSng0aVn/PFM7NdJY4FxuJM3DubeofcOz1QGTEo9E7wXlQLLVqoA06fRjx1x9xCCsn
A3MYqupLzC6jwUHKqM3Pd0ELi8+R/OldtNXdkJ8l/6z5PUcqgG/FUjETxP0EkXXaYzQ3nLgt/dC4
h928X8DcKNCA46mjQm/FnCmOIzSb2LysU+AvwaajVfyG7ITPTfljuyZIUgiJr4pdTgyIOrpgssZT
tbGgjG829Gs2Nh37sQWdsGFhCM8bx640RGymssN1ETH+tgfs2Vg7KycXTNrIRHKaOYUKKGgjpa2U
Ksv3/y76p6DF7S/FKz67b71OqKYl33mvwL7BGXJNJmxKJ0zvPUAaO1OTIxq8JS6HVq8nb2Z9eT5N
oIi64jPiG3cZBU/JZJFQYFtGptfbtB4sWNnfskUMsg2JfObaGccNgCj5c3H0iNOxdPV9pfG0/5ed
8mEPYt3ZB5JldNiWuFTZrR0f7DVS79gSWJ9TrcoNukhX0q5JZWkSXuZPK8DX/X/GyrocY7P3sutA
XmoyKiFg5LZXO8Qsucgk2l/EIh+CSmLgA4x8tO3w6FhawNu/r4CuhGZJcHhj1GSq9mp9741+oOMD
RCxa/9V/gjdD2z7O+/vNVixlph+XbRJ4KZf8puCN0qC2vB9TirMO+7BE4syQyuXzaQp6C3qoRJ3A
6Z6sE7Ctn84l41esZx/KodhiWOdcwFUEi0uTi24hIxGZ0JHkp5/dJxMVzX9+bvfWgHE//eJGwOSQ
NwVfYO281+AW3quzZCbHH1eDLcYe4mSjJa9VVslpQ7o+qpMvtU4yFkigOc02h4dJuIwkeGiZHvSQ
BhBjXooSVs0Yh8rkDDx3wMc/CY4rwap0Z30zxm75cU3IKqBYDWwXss8wlhOg6N6XkrWIf9gnw4J4
8Ley+lV7zXciv+tJ0ABrS8m3CaDJUpKgZj9my4ME3WNrJdAvNkuh/Qnoqv+NJDKLFq5DkjHX0EzD
JSHAqZaDlAnLvq+XeBhStSQ5m+r/lRmGN7AkUjtRvzy/04ghL5YoNhhXQDwGAuS7FR0UQw8d+u5S
i80KqD+2kmfFwoz0KCY5q9ySQa6NYSeKDJ6oUzjf3VmnkTvCD1mvdLeEtrNJkdD9dLzX1/ZtAfSj
JO60u6NQnoj64BUkCyMfnyArBgHHWNluaK5ZKzfQhk2bHX1jFWdlQYZNxeRc9QIpSQId8+/2nGjZ
1RyqaiY7ey7naXTemQEnkjOUPEuGqJoP6uykO9O9Pfv+IPTSoIj6I7ZpZL3e9LTSuapN4oPRU3Om
mByMhEoUe2/mqpniWxvkj6YfuYn/VsTgOfFQtmNTnRexzx6+Tm6ZBKy3yOtH0rnbAt6lz2n4CPfc
z8c/DuMm+qNnG25p9Ixpj/jJHWqRuJtWR4amW4y1p3d9u3nwsdgK/6sQLPXTsgnTsZSAYCpA6LtF
u0sUKboQlzDFZgKWM0afw3wXKQ9uqt52Pf3envInNL8MOQAhz+FLGeI5HSf3AsgMHBaITUDLqAKb
ctv53fq8iKnW3NyliRBRFM2b6GD/Vh/9nX+Qxq/I4eFIKUoIIa9cHgWqX7BJFDTU8QyBQ3dqUxig
7DsUklrT4toKg/89l8Lxlso3rA9Qf7GC/CDvQKnQTI3PRiw9NrB3pW9ayZno1oANVqOvbNOpqpmw
eRXx3atkLPBJI72dF2pvRdXbo286THTVQ1p9Ay7Q7cngKyn7UZLakUPntD8pzlUvsJCgoKsOdM0m
xIycRidVBS/FpS5kE9OXF91r2dsQtF/fDCUuOfxcNiiJdhJwnlDYKz2H2T3P3FHFJEEn8rJJ15uV
0gCcCuyLEHI8JW9jLmuF2HhT37EzuU+EqUKnJP/sG7E95ZHlMorTsU+r31GBDtTsY0+yCWcYuqMZ
ZCVJ/ta+F9DwPnBy60UDzYan1ci450fyNps1ErEpgKIR1IgxNjvpAqh1fUc9sGxm6RN+qD05XR/I
1wd9BKbOe2XZP7BUqTOiQjdKdzOErV5SNUi0Vj4dTGouCuqkM+niGjdEybnPMHLR3Tp8ngYUjWvj
6BsdclWnoca2hML+UorOIHwfBX4xorDSMNLluqAeQDg2JJLB/SfhFN3StSAVYmcZmI9Pp1+gpyRL
m2m936Se6m6Jw17epT4ca5AeKinpVSeGL27WzqoqqeIQBmOuvzBOeklKr/THl05DAeNOppC029qs
j/rStOrr4oOCfm7WJpY3i84TR9dKZHeTpKXz918D2fLiz7C4ynm0MKAtiPuuggqCb4QrEIoxiORw
xuZhXGZEfMlxUxn/VIwvMdet3TxW5bTA4pvBo2KJINZbbtQO/KIPn9OkFThEcjpNe4i7P5xIeJkM
mMvRBCvpLMi4DIzQsYfNfxnZ3LcVDY+J01OUX6JX7eA7C80i4Ly7ztyBaiNCO8BY4rytGIHI+JYo
U6FINpRez97XEM0g9yv3swEbkr6SdbRIgqBi6OTOBhT2vxpMNIlX2earU4TKKIEcz5QWJyMCpETL
LG9M0EVPMskC6EZo69ARzSGsOY/Ze4xfmbR73QXaOsGuMcg1KuIUOVFc7kQ3NuDJbNQLOnOWOsca
srm5NCFIibW+d4tiHr765OudQiGW+TjNhoCxRgyWrwXjncapMJ8ZXKpp6BlDsYLSFh36ZJSR5Y6A
U/JiMvLdc+h0cAkxYbRJ9+ufYbRIPKbfKFrljinDLuU+dMgeUlR1l0cq9VM09Ufz6qua+py0S/mC
Atvz0XznbBSVbzAqik94YR3VttAg7MYaYpo61f+24FyYf1HprOk45V0/wzUM0yE40QUFciBjiaCb
qeoYT2TyeV7iPJWPn4PKQb48CIDAonuHDottAgk/vjVT3caZfjnU7AcTdBoMGioIDbKQOmgwbytk
Up/ku6ShUX3JBPo5qXfu2tGVdLymHJumdnelxkmKh5ednNGb5tkl07RRiV34uE4V88A5gmDbwngd
8j67PACte1b0NGRDLbzneUCyoFhEP1cHQ1Dkxg1qetTh7XQODeyvlgPxtnUxfoUGG0NyNn9c1oFS
rxBtXbiHRSQkX+SODWb7FRlwhMveUqQ2LiXyOBQESs9Aw+2FVBLJq6Llp4psfNZk8v+nOgUqQ4fn
sE1p8TQkXwFO+Veenb0PIet/wn9Ro1Ho7MC69KILW0Xh+jzI91XYzNA/2ee7OUXHvMmZx/ap0+dj
IhJuLiuDLwvdb2hcjUGH0+ffSVQ+NSBM1VcXrhJyBUtrRl2FWzb5/5O631Fgh5VTsOPE8f/zHHG2
dk1ZSYxf55WlfC4efJfjsLheRvmgeBJXFQLmvMKDfKtbWqQ4mEfBA7gEMeQ0ZSe7mV4D8Wy2S6eY
i3ONblUgT84snrKAtUnSSLIRwW/UrytlDeezC3Vla8+ZucaQ88M2C5rGV3t7+7gb+wapfIR5o3Dl
wgB0ddoOLqVf4+rrd0MLLltHy+L0qY+dJ943GFa9fwA6bnHL1gyAatzGqqmBBQKPO6fSfAnzvfcS
EkTTIReA3akOOYoJskWSZxCo/Y0wJX8rylx0C0cQOqQxwzeaNL0UBnQ8e3IU7vTKOEVe3FdRKv7m
Xf/cBM8URo6AArW3pPpiIwNEqNvUz9bIOUb3ZxdkH5S+QdgLr7QzGFb/td7Q5qhkVsDnDn2945iE
N8363MTS6sWl5ZlT6GY5+mvqyelHFb14LfCbefFwLCQfKCacYoL/8kShunSSimi1rpHi4VWjLe1P
33G+3/quXJy/QCb5A/5ztvAKS2l+MAhSInK6mG0v6QNwn4bkXgQJPsBUy+aWbjXUsnoOIMklnKFr
oVKIvs5B1pTsxQA7XC3Zh0wZjAAM9oXBXdlmIuPp8lL4AgqtG58M4DFmpDYnKipHhLTOzIyKnid9
6d1YLq0yqqDPfjdWEwYPORfiHa4Hcz0OchrPoHJwHRjVt+JGkvN9cX2rPsjpFXIRqNAejOmWX3cm
5xSWntvMfcNIv2Arm7e56Z655eGW1hoMup+mpBVmpGBcSJuC7yI/HLxbE3fwS6psK98M571qpHPh
bdoU09oxpO08hg2MDSqpzoiW7gbqVVb5emMK4w/4Vvw6w1tm6tG72s23nFtDBz7CxRl81YpsZVUQ
eHwngzTJZ1GQudOHTbWyBjXU9S1LXzqZxeeEXY/ZpBUxAGveyldk069MpArz8okGCKQvVYG3YZhI
pHGKq2tjs/Ov3EVyL7/z7ht7/B+/KrL+x9QZRgb1ebYiu8s4louY8BpMhchq3sclZqX5mWkUpmTm
0thsNauH/SpUe8RRsSvJKAM44TS48JeXl3pYDSqPRNDQlQpxnRAPtvF6kPgEeBrxWBf5dDeYJCJy
41wXih7Z/wnTsoq5407JbaYkj9oCqxuNCAhvmGiElQNppXu9s2npy4K9zmjU31FzcUM7A4+PsuQf
hugiJndMYdSUVpsqkiizzkyA5TDXouQi1Xt2EfHzygIDvXmnfceSKzPBYjg2toH5RZTcvIN1jiBM
/tgipR5LcFfqS2Ksj4YDGEj5InnIgGgwTCzzUtKFA9TGtctX/Egv7NBfH3AucsEyx3BtXszb3CTl
K7n8zeWcFfIJ+wUbwXv9wm4ITeKlADU+qQYd14KzfPYgSgvB+19AtFodWdG854oF+jcyp0YG1z+L
49ztHCUSW3R3fR60wCXvJekI59qtZvjWF881Tvg0Dj7hUMshKfXB6rQuDVQJf5msa/19wMPgsshI
RkXEdePzH0gM8DJQSYoICGHBRZwJLlQJ6ID23CvHJVMBvH+SgYjoSA5z+MdWNd+TI/7WXGvX4oQj
/jZOTDbYZO07LUJMESQgbQFxySQD8IDhat4F1Hijpc+h0HyS3B6IhdEZfXSDdwoyFegQ+8gW03Jb
OEPEAO4ili1J0KA5FUVbzKFRI4sZUxj/HElLIsNAuVRvzXWGknAL3YRiL7TQjq+7t6MVP2u7FaCL
UUslj/ckcrkJfcfYVhf/+U+KuDEIw6TCheExjv7nI0hh3MW60/q5Gsw011vPICcEoGjw6GnbtdF+
INuLiQGEaxS8N9l7bcxdVvATS1Lzj4IcBRMD7Lsg/JvZ40BFTdCvYy+BZIYpux3v2aaYkf+Skkpl
EpBzVqkadrV+t8ARE860NiQxrH/a25n0K9vFDchILGp3toss5X/NyCgg6XL7grgFUr4THiTzfpNq
jgOIIVGo9SMSdAvxrdbDrPac/+hd2YkRweXFOLd/ibxVn475WFsQD0z6QjSSevUoisX4qSDcZ8lV
/yF/ucRIvYlBbhVStQ1Y7d/Se1QK4P2HUsoU5EUJoJHIBqa+cCzV31wCwx13g8nauQDw/c7JlRxR
rG6LNDBMFFVNd2yLElJAhqLZ0BHDt/1kDwl2eFtoDKb7wS0/F9QXdysSiHB4E6UsXagomo9Tqg+e
JFfcaumj8I4S1kVrBrO0mo31sqghbvlAD0xzatm1tZq8IG/FslovfcTmuQAyESu+D0DsY287GH9G
zTNHUoAz2me2h6AfTNpw97Jr1x57TZL8hVrVp0UQwJivXrKYO83cYTPzAzJmEQEteT7rItraACWy
pUzZcbVQFQQ49jvy5t2DZXiHgbd10LYz1IZBxgS9+zaSG48WIwNgFeE9sRu1ITZPQb36/5/GajLm
mgCFQ22oTxN//Wh2TncpQRZ+TT3dlvskGVsPjyDl6jydyquaMD5M1pzcKjpsZgkonASQZxEBABv2
p3xRooTDbbUbWVnuHaZnI0j15jYj+8yQv8SylALiB+CcRR0A4z/s7aWALE1981gyS12fLZcE15Ux
2D6zGcrTA7JlFSoieUbh/w+9sy6B02QOMpbKsrwfBidEvM2OLbb+WOGcilRjyFW1nqA5dDuhea2b
oyWHssoNyM/VWBIHLQvDB4Yg4qIkKwelkGjc+G+x8l69kW/d+n85Q8If27oZLhQhM0FZTZeQNAhc
74kkZb/nkdRWnX18HSAB9BgA2rd/Ao323P/GayE0hls0KPbqjeWgzlxYfi2Ayizx4Vyp9aiJ5xPj
opDa/It7kJawkfFFzMfoYKZFjkEG8oOgANhb6pHIlgYHsWzp0vHhWgcCDDOshKGmKuFkb0PFMvcX
mx5WQfOwsiWgp5+Z3eZ7puxqiZMDUaIidt/s+QjUG73lZLNAURgdae6qIsFs7r9ma7HJj0wpLgMN
0tXk1alizpslrePfJSauo0V0xyk3LEbt4Ub2lrIiO51xnjTJLLolVhNA8vyw3K7X48dQb8XU8sxK
g//TE/EuMJTFV6+YACYcGBVOnPREyPM7FMLzPoViBPfsHA3kX6zL3JkQ9V7sEOTQNi+DQVyBOtei
aEGOgZyGUOiB+zH4baJDNObwLSTwHYyqIh47l4MEijocn3dmKbocfFTzoYHqEW58ghP8noSFKHi9
XNwLGrJ5r6xn6WnEPCzuoed+nux8Hb2t6sjzy8sE6J4weIMWIP86btj0dZ2R1ikmCjdyMylFW681
7RBeJewPnwEzl5x8C4uJf3bhCd1G2eDKnOJg02pcsh8VLFZw/Q4hJRAji7Psr7HF1+esYPLTJjf2
Q0VCLRFLZdF3lEUcg3qPkP3R76YJv2ZfjlXZILkVEhxy0ArRstOY5DqEnL7sqhodeaUXTjn2NFlj
bM2rIkMzbIIWstq8bavTWRizjDOsnoZqyQcC7FLmwoUwcI4yH/sKxWHIHomu+MYJ26/3Yx9hiGT5
9Ktv0F5JNJcCUQQ313MvknaI0ou21nBBiXehaYpYGXmP9IvKSgu7nKZRmwVez9VMn2IgxDsjQUjJ
3CBAyagDc1y+sQKbb9F2Oqt9uIokclcJiKXNq5JPRnA4qj9Tq750GZWgQSUeIbTcsvpdIsXaGDah
uDPYnvBahwQ49CkIDTxTr5AhcyE4rbPBdQ9ieMS1hK/8hCHHqDMQJJSQxoZIzv2Q5My/vZeUU/gs
X83Vp6gRymmuwdnLenK9xDDBRzXTx//mfNuP8Ztl9qalIjrknlgbKu5av40zBzb1fYWo28u5rn64
pwVgP6Y+nhjxpcGoKqCYRKdsmkC6A/n+l+XBxd7QikX3LdWWt1YC5b9V+LWz7SzizsJr9Si+f1Qe
OlZsNMtv0NOMBux4FQfkRjLNZYdWNhLVf7V6nnuCeEVVs1zw2UT4J1vOwEPgWkJzlGHAVB72hvvD
a5YlgAPyVrq1/dIfBMtjc/4TjdR7AoCtgBHPyPe4noo10Cds4vSmj2qUViGwfrrwZwEqLkmJfeh3
F8taDYGUzTtLHQH3MS4220dHFcxGMGR3sWrGaFY1dEbK6B7r74QRwnfUOQIzki62u/z9rmGKAmdw
383nM/tw0C46zTDQQFVCzfqfxcNx2BwvElPQeoQn0Es2/Tzs/6ML5hY0df3Wd6GE52MBL7BvhMsX
dDAghjYoQLyFTFzNY3KjBk35A9q3qxY9KfbTvB4BCIHz53gJ67gWHJJRCi61HpkSlvafMbP7K0dO
Q6KZvcLgyz9VTHtr2J+nJqWz2fhxLrxrEGvT5Qpx6/OvqyyAK3tS50bKfh0ZY2Z9w6I9x9c6guAf
dZnEf8/uCUKh9o5mxdcBaWDQis8zzNPvcmP2ZR3HNd6i+5qWzniM+u77tZbF1BjRsa4ksNJdwaEs
fllmkKyznGtLKdv+BdWJmR8OQreYzmumH4UGUqmnm0EGjW2MR929YvX5WV5DtMmU1j+YPaOXVbTi
7OMHGO0a8KO0lJ6PBfKFMkZMWcMfXeSRmHaGlAKopG3pSGmeapdQIZqi6wgNTrB4hSZrE69ccWd2
IAdwSZ/oKHRmr0tHJH10YPvznGAV+j6OlW+RwMNfB4mDV2/GawNog1TzRAHvdg3b0jepI+jQPT3e
p1of/5XuQyXLBasO1R3TzFvYtQIJglo9lIReoD6/v0oM6dO/mafPla02oUgh9UXTEjwteylG9J+e
eyDQGEwQM3AVcfjf1eisQbrXxwEasz7eun2tTtUFAXEkCexz04l6mvRZjg//bZBNvn4cyn9tyqZO
aQFbJFqL6Pub2WPTFJutxxDn2Q8VtIA0KyCYgeWgAw4BRXq1UFPDCbDisTLNTItdoWQ5vqcSO0XI
x0glGk/4OcLTF633xNb8dOFcvclnqXAAIdVHGUrUD+zfrPlMEWoIFvwB+w05ucvUWGCMNWZPGcYz
MKKUJkpQ+HEMRCjn7tFgPHp7G6xozbewLy05YN5WE6jHYs07iu9IdiGUCktWf0bDV9F03PV7ERG5
2gPSd5YtdihYj4mEF73fwK7YW1kZt5SMhzz6oRLoaHa6wnyiPZ5AVJFukiswoA2US6foDiHtYl9M
TFHXbXJGJWyZHrFMxY2tp9sC5oI/IcItjVUvOdJxIDhl4OFUBaW7HVmf2BpchA9OiFoJM38cap8y
Fv1eNjsdjw7UxUODYFb9deKRHiQvbN4c07ohE5m4Awo6EvavOx582Mm2PnK+RDx72vFcg4caJIc7
e9w8S5Kqx8rGDReCgZCAVxymrTtoZueFbBV9FM5PUrkjAE7VbPv8ixbF0C3lY6pwFv4vEqliHL9b
j3ArOlzTY58iKBXr4GovB6AGpnwKZXQXeq4/i+v6R8yKx+GTdnj6kEiUgCSCTSTcYfnLnm/FIIU9
1vGBd+8lAKzUUQ2qKkFfi1elbVLKLTiiqlPaRTZNCvtYLLzvmjsADV85KSvIgLoNHOU7xvE6J09T
mtGTCu8ji2U/sldSve9srZ31UmwtKkelAGMMC5C/+9tyPqKd0EF2g9Vlna/5ebgqFSocLusuUBhY
FSP5yHsif1urSYuxChZrB+svtArZbdUEs69TPJNM4zJ6Y8+2YkGmnKjtKZmTbCmtWfwWRs1hxUyS
uaLdYNPfp1bsc0ILYlIsPDAeeca80Ta9NCcRObymK8i4gtQv45cWMVIlU3rIxKSe/4cK9j4ZwoYR
zW4oG8Bn7QHzkhq/3u2j4olbYWjc8RrAUfOTyhnglCmaGdhBO/1iK9mXv1y+Q4oUWXLbo2zmIORp
RC4bKFDM6KwKxC63jE+sFdaq7Qdq2c2Xw8bRviOld1EmYCAKQSymiJUYD3cyVar2AR03mb/ydQdt
nApeGyOui9Wf7PBnVBReifcDBRw/jVP+IzPlGOhMV/eHd2ziS/L+ffsw0LwrUkIqEcjt8AKZ+m2v
NLn1t8vw9dxG8KoTB8Yf4AWm2LuFoVX8CnSMk9GbgnSTQyNUC3M9B2/U+E4IooAgGCQk359qhjrH
TZmuWZSRMUGyvOPjW5X7s5EDX5Q3g/aKVAa8zjTXv23LGuZ4+qDK1VZfVq4iGq4mNwX0u6XRzrz1
8kPHo6AW1Gptb8ljRT8iuPwtcZduSbTWfl8Q5MsmrEcDVRt0Z09C+vXcUz29vMjXV0510TkEdeAI
OalJM4Q4zZshCKGqznu5m6J7r38yFWKk7686l6ffCClbCR8qtFq4gtwPAjLMUh6Pwfg+OcklW2XS
lRUL0EFhtGH4jsdK4R4L7zn6Gry0acS4ksxV2E7xSeAEhtAeTqaawdNq3vNr21fdaUbTQwZimOUi
P8QuLbhF5zOl2zktyXzFdLNorWNlQm+l0OQPZprZjKHZZYAEqncIoecj5fJUTH4HdY+v4i9tFiY+
Ik/+RvxyK+4hznWh26Yk/AE1H/ckXRKHmoolxmEGZ/G/zxf4mscqq60jjqgUOy5dwGPePa6vKvLz
fpPJR2JRzwqm8UTZZmZqpZj95CSYNBFqq8T0kx7sqoSTCSTiJ51QDK5XkiMqqfRIKxdkeX9ilhl7
Qsl1zbbOKAx7uvXj4i6LukWl/f9ebIj26gZp3gk7EbLNoJ4JD4RqFqLf37NSqCzgd1/a5rdVz1Ge
ADNm0p6wUqjZ+F4bwE9uafMheBUA4/e6JRlWWFwCb0giXoEclNvII+lRdNdcGG2cya3dXLfPYnG/
kEUoA1mLIUdoMBnxqKAKzoMuimzPMA0xi+Vgx22xqtSd5NbQ7JfmdaNqW6WZ9Wekd60gTUZn4qby
nb0PaWrHvWLxSBKfYgk5oVhD6UdlPwQBI1nvvd7yyDEuanN6XdLiFHRmcsOpJ1/VzSHQL+Zg8c9m
uNIemWQg8p5xfD2vBnWSEu4v1L/bQ2JS3lUazaDLToUhbtHGZ9dpy0SHrYoIIZFvs03CR66IZp/Z
2yN9jNQsJk1r/vXJJoBMH1/3G6HVvWOYBgB6Fcdw2XoR9ppyu+ZB99+MbtvWWWKy2q7ATvkGvoo7
4TDMTbYUoDIiKRhtGoXNdSqKFGAHdUa4XsxPEYJ1MpZvmE+8opvBm6vpmRgQhhNfsyHcvFtv1PXd
7xZ9hp6hzUrsbZkr8oq7Y4mMFbFd4OVmm3jewBcnbGFVDDAsfOhJQqSoqbhoGsNCJ/4bnYvDJKk7
gqcFROdx4/ulewAF2pu1A7PBV/aiKPJVkZNRh7akeyq5vUQIFoErrNpHMGoCbuncfa3KnFBDqbJL
AeYS+sT6C5zdufjXd+SHy2C8w3NYGP+zNRkhy1IJnBtRii9YZegB5r4YIMp3XTHw74LAdRYLY6xh
3pH7NLtASeiK01q7PPGsCmXypFGq6SxhahJBhE6axdnvZdGIixjT2QWQPkDMH5FQEduB+hdhZieW
Lypgcpfql0hAVmlAay2e9FafUHw/OqAglTB6p+pLKkxHK98iGuSRDHCMzRB4qh2jttWT9EmRtGfS
7XG8PqUksCxVSwFrFt5aIuk54+DaE2sWfZKKLG6zzG9MW7O0k3jG731h4Mfw4FbuXt7ue6iDJFrb
YbbPk3CF4CruMaYrbLA4rXjg/6CF7irA2a5zX5Ew4X12oCqva+65OQCMn48C51LevmI9cDeo1gAB
3XxyeWAjZ3IBFgq7NIztqW5mOnbJ14KSJWxjwQBT0XusfXy8w5czuMkGD7N/l/KC8A1cBz3y7wJp
oceh1nCt06+eqOygd7xCbQBAZYwuPDMCB6MQaRi817HEaDeO91CKdhrbTE1dH5dtAiqkWjWMJano
AMyvq6gXseKc3NJTsuvRQGGHNGWA48/xwUKg+508aURWdgcsxOSEQxitJcQllV3jOf8mt97ZjApo
FDiz48832aDqsn3FvvkupYseMuiRyHC/JaXCKsK973WA0z42OkIUfUMlz1iV/gqiLVod0IUhabwF
vE3Huyf2VlZMIW0J6eftQphESPtt480jrnDm/fxXi6t27uZrod7spIa/xYaRAeuR1scACVqAiOY6
Ei2zaSEoJHPUL1TY7yW3QUiXyXXYRdcvfYBkxcQJDkJaq4Mc/62zRtm/Q2cUI71M3FcnkMOyNjzr
zrPmeCJeLfUSMS0DJ0lFwhQDa25hB1jMZ9/1vcLW+OHr7SOsWdEgzS+jqXmJB0xQvI/zW1kKzMnn
ITg2sSup2fHuee8h15ClF4kl4LUJDYR9h4aCWsjzIDWzbNspNtoM3w+WvFobMYaWtj0asKM7Lbuz
uqt1K7PjDvDpECk49uzkhAKTyqa24YmJBxhA4tAZ04gN/HPqcff6Q//bSz+CMejca9ECI/MP4hPm
UzUBkgXGfO97ObeYgxUAmtg/6Egta0HrEGY7VEpBNFPWJ5rr253fzm5QsUTbmYHL16dDvb2C9sMl
If5WLc/MqMslPyXL2u8HBrODalNh48LscqPVVEe4+awSj/xAM8auZxMucOfDy67QF3hVYhacmTKe
AfkOvdwVCcL3f/qWQg1LxtMtGQewZBPtGHfzrVaqb/3d1Cs/vIq3FhQHw8xuhcqjvxPiMo4oF0L6
7CjWr5kX0Ocl9YoeleQdLec4cv9EWa3sWrp0f4UPu1w3SHtujHV8dUdjvy3RkUJpqeetxSEp0J83
SL2F0we3pHSMbZrdjKHV6S9Wj/hNz7HEKI1SASZb2Ye9d4g6nCgGnNzy+xAg93RXVxKDBrCMfjCU
Sdi74kctgCHdsVrhEhvc/UhWxk4GDVhNV/tYe3bsXo83obmSeQy74oH30iRpNL/z90/+fix4g3jK
KCMWGsRnl0kWMjF/k+PGUpiAqNuoO6WOtLD1MGTtdjDxbfOS82db9x0LTtetK5aJ8Olymf7ciZgp
Rnd5lsGiShdYlquz85lfMBkmzT407bdTTU/r9p+zaDwY8QA5zSFzOkb6XUdrL3WHCfIe5elEy4Rx
w/YkbgM0s67wIwusHWaXj0P7nkudlz1i6N2PUKnOPB9CUUY3rgtCM4Ue4H5inOaObtKKXWiPntMf
CHM+BkV/vZPLG0yb3QFmP0CxDm1EcMUTqlAHZAbfpE20AL86UPwBweRI8n9ud4EjD2M008opLaUa
05grEr456RtbYGBA6+AKmkQnF5HX4dASWqVTh35ChCWA2NUj03v7f8JMoiKXiYFC8Ib5klFDiK+k
uHl3xO6qVVJz1YrmvvX8PN6fE2QNVzY8/tCjrYyS8Z25JZfUX5tMbRSGUi+9oIoqZDow0vFMFeXe
JQjCJ+fYWNLtv3PIn/B1HF83qVBDlS93eN2Ee2Lq8fScXllfT5uJzzW1+Siul3YwGtYShaLOuPtM
h+ttPbT5eYIDvB7pBP8327BgceVaz5MDV0zJRmWx6g9g5+vr1ppMJvtuINwINpCgSm+6JQl0p8SA
elP+gG1d91ApwWG5ac0xa3imgMYaNXlrsu7Jw64R7u7VEccP7tcVSj8Oj4+eazOCXHbi5LIXEoP2
aru5Pra6IjUQ/AyKeF+ujmi1QAN/GQOtDmNBm3Sq7BXG9+w9rsuNVjHR4FmzmH+qsU0SIzNVf8L2
Fi8O3wEQpS+85fmW5sCiGiVb9skNow3tFxtlqzY9jA3OUqbkJCwsRleB8KTYOc2BXxBUcbQMwy68
zpA7b3CEBcepHlTjF2FYm19nuT1zKu+13tjQ2MrKHf7J+gJCqcA2orIfb0diw0b5wUPMubuXId5N
HNWpZx5pdvu/DD3eOyS+Y+7Z+pNb+vBY3Yl/nhrQLgxPshVGuNId93/R3waySBb9GESkINaX0ur8
I2GGskwQPcL9zfCRA6PHBUeK0sai+kD8T2YYW52nXEGUmwO4mfxFfy7fszvBz9hbq8VNORjsW9Nr
FsxdRjpPmgOcDHD6FTPnATWQLkRl1Q6zzmWa6QqSTtov7FOYRD38Ue6g4GF499uxJxiGwDuIyx/s
xOtXK7IYoMh+3pWhz2WgkqV6tAsLSILN/qRUpFEPdz0PZvjAcM8lc3BhDah9Mb/3AOKnVhYnCgjm
TBKpl2bwtQMDy/q5Zqn66k50YtNdzscRNF7z8HuCs1vawNul+kQ8u++rOI3StfP9qVSa+i0GW0em
8/KgDrf6xXm3W3O+UEr46cfniRaHBomXBtlpSYlgY9t8Kc9W/p+aNPx82KBbrsv2Z+8EnwjvvARa
+QVffo6MPPB7tuPUfwBc/dBXFduwkF8hZWYWw1IRQmax2xBi4oN4om5OKnsgY+HZ9rZSlcpQ+r5p
rAbYTpVulh+3mtV/3XP/orByKwZX90jxZAwBszoJMyf4jx1oPLlfZldEXUYNfcJ0SkNACyNh+6hh
TR9jLbhfiV+Pv8jLzgUCXFmyLXF5TzEsaye9JqPeInP4+/r5aMOaZtxbzx+e5u411o8VPUJYQPaE
3nFyjozPE6/kYsSyYGPNx4FnyM1kYqNPSr/EB75RyH1O8Hi++/RjUpFner34M4HD5CJrgjG/CaWj
vTR9ywMKZWEdwwdlRwtG9eXtnMXjTEGycAG/nrq9pnD8CGslaWGZlcHt6BjPG1/mDaw2dTEr4U6Y
u8yU6Dm4Hl3FM5/LpyMt3u9LWU8pAElJ5tpMwGNqzC087blnLC/J6cjAAyVpt9EZbRxRSuetDFY1
gBwKR+WaPL+fJJJo416p6yUUpEhmr0/7uNkkZyjuyvDjvv5//18PUmp/nR3Fe7F1dDM4/y4UlYab
q7zJf3VRL3PWjtOBl1skehKzIfIE2ruJLXf/NBMz7NmQW1PH+T8yIDuA10UGsnH2uSEWHSpeLM3C
X1dK3dzOedyXggLs6n1Fo2cXY658iFn1nKP8qc7aOUQzpPWLxUJusJ3hqoQQGqskWSDHFSKqFIwL
pZQi27LiqU+bwvsV8wmOkgvNE/U5B+6gU1/8tNMK4nucpE1xQpdb2vwVbIJEeCEb7gPHVoKdTDKx
+/GslSqouRhFd20trtjtaYgeDcjxteG6//ntLvwJb8AtQz2x/2neqnXnOLV6U8lyGKp2TC+0+BvZ
nxP6r6cATQ7a1V7yDRy/nTpwaAU95hmUoxKe8rXAsvTYmHFETqgmLU9wYPzgPEMQO25QkHn59fBW
5+hhYRv2Y5bq+SEF5/wN3t8MiZYFDsqy4JusYvJwGPwvCJlmZ3oHkEWIe/qv8rlxNr8hW7GsSVis
0x+jgcPDQrpoOU0HD2/Met2Fx8LvtF7AqBRvhNRFs7XWUMFnI9BeoaZ6mePevb8sniNf0JfHIbV1
PTLpjY2j3FIZESROnM72KILGj4Xg+2f56R0z+WN3wYTvBpMba95olQSnnEZymGJs1ypytGGHOeNW
6e6Z1Rr9wOFLGgjApgF8OujMntFSZVWXV27us8QZUTOstL5ViT8qmyLOlBwQPX9+tialyxmXPPE+
Rjxx4qS/zeZ5LmT98NuSKHL8wKq8wCoX5rrZL5TZesZxKNlnybx8ddvLPijWSLwBn0JOci5qvvO+
BXFGQCny5nO1GmO/6iU8a+9m9dvWqK76PL2g2VYjX9TKR7LnzTWMcJgp041ouvh7xCdDxYIp83jZ
Nhb3HLZaZXoCH83fk+2Ia9y+zMVviRi8l9pv+ZTJURTcRRVBQwmNKpTFzAn4IvN/B5PWN8qx4Wmi
BQl2t8c8Qu9jdhyv9tHX0mCR3LaHGTz5LNxEElepvjD+/ULQOqP7wmERVNygGfX4J+Fp51oHKXB+
ERubNNfakB291ZYDv1+ovI2P+rXeY1PpLpAVEQsHtIn0M44MrAd56J0D1eLamoD5AQHPCyVsaOBn
Zt9Qaesrilom4l+TaAfoPWKA9hNAaDVKKh6XErokFKTSfy82KS33FV0SwgoKsJ4CvkjwGYzt9SGb
ZaKCsnb0EFAr3enpGJPTd7VPtf9UV3jmF8uH7miLsawuMAd9Pg1XvHH4Y7guQ6gut5TPCY0PWuMc
52ZL48sPNBnEqjb4d43ZSJwBy9ZO1v1B6Z37y5X5obPLnCzIsrceK5mHhU9JF4zDt50asNWbOh9U
eSV4ywen9pRiPvs5S5Ft5ljwcP2lAskcC2M6QUp10AlTLE8oithZr4hlMOiQOu5AyBs6kz6sSC3H
aSTbKw1OUFfeIDdGRKwFFvMJzCcnlxNgEuxH6d/n6twaxnG+bwUzli2yqksujE7d2pHHp+b5/D6i
X02VWWnxqdJ0VWyGz+v6CUFN26V3XGdrB8DJUM7u80+Mh5dQsYgVzad+eNzajGv0uWHWHLsIESWY
uxZ8ZePNWYMebT/uaTsPm7/gR6D3nxHmyy1oc+4wVq7j/sXr0hatbyJBIJFGtJ0nYi5h+sTJh6QA
T8VoLft4Vx6c5MRsqMgPG1YrSK6bL6vC8Gs3M9SsGs2CkMuStZqU0FpWHMEXjsA8SSTuu70wsbkS
OwWqQc1JyhjOasWjbTRf9IWDD4YME6KZhHZKKIogj+QYvchSP/tH9F9JjkNKpgGsLjdylWy4b4oS
i7QMXjZFYMnwdBlNjp00UarfkOlb+3O9ReNBqBhZon/R6c/yflMCzOzZTZNl5lbogz/MRBES1jZX
iKOwIFOsX1RVJu3+Foa3k09ZazaxgtlDmnut0W9e6+vZkY5LP2QB4EWSjMSCAMcKEoHoqvo7tyNr
Fifom2/w8qbaKfUohX5PEI+3qVWD9rGy5qOOTOXqjtQWaalqvqYpCroPLVzZSi3dqv02sZPzrE/C
Oo5i1W7QOoYjOcqXshXHlFv8ses2zHUjHuYWxbIhGoLWQyvlMP7eekqraF1NiMCUl5y+lAk0n0wh
JP0gJAysIooDZOOTNMe8NSTwEjVvK3oQm85BZC/VgyL1QUS3tdLhuiOjwhUXdzjYTCZjaCI1i35Y
Amubh0DzN1Q5E2hwBhaWzbzVAipzE2o0Kr+EfJwplJgm+i+URVekTFCpSQm0nI5YM+i63fY188ld
0YxwBPs5OcNNrAFKEvMK2TWIVTy9tkokqEh9uVWCY+VtuQ2QCzsi62OPFs+66yUa3llaQH0z0zRB
EilN5XGqAoisom9EzIqawqdWJDKgWe67DKOVrXuKox35IcbdwIQKZjh53FkF1v/6R/IOYUwyvF+z
S9/i+kZRGRJmqvVpphVwVXMJKyBDTtdN++dwNO70EZorW5p32ij5nsztHBbs/rpm4gh3Yww2UHDL
0nz4zMtcoIJiUCXqqiLok/w3Igz2/jnoaMn9LEbzO1pXursvv31moB79FQaIcOW01Ynz4tzkKbKj
Bh2Fx5rL81vTfx/8Rme+GFHyc1Xamm70SnQbM/y431dKpOPKLaRMtDit+pC1sdVWChWEFil2hivd
HdNbjvAePM4Bj7WebjxvsSseggzS8h1U0OAfuM4DWOF4n5Ao+PCTi9m7DZ53inaRv7JOiGfjH68M
GgRCGtGKeF2NGYC7aEe70rWkrz+lzmxedXtT7fNhfk7B+wxvrY5uvvmxoin1R6DgpmuCsH5Ebqlg
t1E1YYWP4fR5UjcgdRWxZvLzRyx7N2J5fTT01fEfxlXOMkIEp8+JuqTeEDxywhdgnrMInzTNNI6N
o1qDnFfjnKodV7sqbZzfJdbQZirT4ea5t3Y1/z4IFVnTFgv9podov3iur0bYsMvKOQ2gYyc9/Mn8
ZbjCiAxLz5/KmIeHEDTeQyidCph3y63r6J76DRVMOVljYGpkAwWrBCpezWGx1HaI+2mWnol6H0TP
gb/wL4uqMCEcridbncVdCZ2fZujcqZyhhGEJeiBMVRsr3A3up9cPh4ddqgo5PvmDvlVIs4LucjUg
VwxRepximXAR+CsmRjGn3m28owobfn/w4Yigp1dz9kP7WguzdbFHi/yzslRIt91pOXnSI0EOhy3x
J+yFwRBi1EPcikTwICEJ03Zx2U2DpV4Z3+4anFyK2dk7MkimDu9xGBBcP6NbUviQeeToRPcWiizM
uwKYbU8mfpwD3cfAjMQ4mbfpFrZhAw+G0QlfzmnPf6QAeXObpE4h7elfWuVB4ID5jMoUvi+/M69G
0b9H0nXZBHMiBEX5PPczaxZ2vvZanm8aMOOorXDb3WjxRgPGSMe7puNMC6SwqrqEVT428IwcbDdA
vYdSfPKiUkj3/R1VY09RfDGkrJLixpfVWzZ0s/UY7rkCRp2hnJZgOqrDR+y68FDD6+R4xLRqjop1
xzJqIuQov9JZazDCkwA13HnaJnGKkz55IJaTAdPbI0EF6Sz2oIjHHTYsiWgWlRr2sswcABumBr+v
pBH94Bdt/b0qjFY2RhOib+ParxpS4Xpvr6Sr04wjT12XNXky8A0nJ+rDNmAMp9jSYdpqA7bFbhJ3
jDsjmnB3o3l4i5kKzwPgBn3JsDaP0pxOSp8g332qAkh6LLTiZ/sqERzHZp5JRI5pRwhREs8VJrk+
ufqwYD/M8ssFuXGxlqB1HaKaW58b+/19B7VFKnRWMmDzixJu6wGAKYnmdmF6VhJHDhLSqcIZGMBd
BOH9CfRkFGoJnOjiOdl8t352ys82dVoGZmKGShyHbcxj2ZvDpBNPgMDLSL5nKkeQwVYyZDL59inb
/MEGWyhgrvEX+3JMVflnFHaNkSMZ37Zy8T6uxWwHRKBnY8gzhQofrWBUh/s2SKRGlxURb4szsd6q
BlzTiDl8Mu5Xxs81rd4+7DUwP+HV5SbU3ii6ujygi/sLeixJA75GXHNhT/88v4Vc/pyUOTQgrKD9
8cjGBJRQmeBqJETfVVRXdiiO29EzePq8B741b3Msi3DJcnD+/VM2l6CY4U1087Dp3MhE1f4+MFnY
GmmFx8kqHVCdl6tp3oeAMYF8bdrp3fLCIuNDq6EOaUIvaCIOYdeMdQNIVxBOZ/j2DUEBxMExb8LF
9hBtpmH4u2l3ANrObkNxuiZZTClPgD2juWnUpL4Y4rziLt+dxzf7V6zlmG2KF9hVjgW5zD958Srl
4Hhp2c6VyLNGANhb5CTEpP9VQA1Psv66z5UhMI50oo85FATVKPaW50XQXIsNNUin7qGRLRbSuHJu
6eE3nSH5AZErWP4JOez/B3cr/Es4aitc3F/0AOAnrl3YAJzYY+W6O/kSGDHjZn/4AzY0ySQBjhFd
21kEpEzCDyH2E6BLcZD2Q88jSkQWTdZGIMLp8w+yDu04+HqOPeUaXGIvPoVcylwTCXoAuW0Xd7pa
fYnFzGJlv8+FdM/QiMacroMX8DeS2Jrw7qjFseTBiKE49lTtzZZy9dd6DEkEw6NqBwpMS7zTKDd3
Czw9CKEmmd0JY7qfxr6sJhR35WYyUFEplW8sKZlABXJVn2i19Ec/T6WRKoo82JXV1n2ktuyljTvi
yVl88bxZLBoDLSDeYp1VN8Jc1PKljy1seSNgXtR9Kwgi00PjQTfU4yUULfIyowuWog//N9OQWA/8
dxHuighh0RghdIMcTqVNEb8XOiYOO/12qYWr6M2lPn9D+pmKxLUI82nv0KCAaEvs816q7tKdOwRc
4bRVYv6Duw7Rc5Blrst6q/Jlpykk/XNs7h8qDPuR0Kdk3cGC1lO3Oc965q/20XjTpOsKtlYgYWVk
GS74PtQrjjFIxBfzUzIBlj+tDicWMz2YaLeTESuluS6ANBUaXY387u9agCkXpWqXcZe30NbE0nC2
hb6okYPOD9fmmf9uMcp+8d5+xwijoVX2kphi7bhHHXPGoxpC8uAj/fyAsmkTuOf126SiB2bJgEHK
Kq0BC2tU7gNwVnNfACcD+Td0TqC36+3r/HIYgdwFXrPAHiUib2Inq4Sf8QphN2P8vwj5oTCCkSgT
2efDMEVdvUJUsz3HYsNLEscoibcrUOGpgEzIAEHYcmw0EA6/zsPib19rcHAZ28OABlM4Wz2yB7G8
pbmFp7jZ+cws+PeUC61AKZgWqd5o3bUYwzQ8GuV6w2dsTaW6AGGREsYvZxs/CIybrWMp8Y5iNIQO
C8WkWyxaTlJzT4uptqoNWppbd9Zd4GdJR7GLhPGy6+U/xoDWSAx8o9LTVhBIw/k4n7otKlapR6w8
AbbqYRTyeqsGGo0wntr7xhDItovSFI4aYhrwJWi0LH7sfFHB29SdyBYJSSewvQFEoGe597wFABjd
b2HpUfmmjnQ0jIbmJAAwMw4Xg1rjmAd4gwOnzN0OwN/F1DzK4k1eSeib2qx+TGBudBVNR5IXVMW8
sD/G7PzmX+iInFBTHUzRkQqp/3fijCbGiZiHPm9Z6Lv2tElE9NDqDjwPKMlmRGCDaak4oNlCtP+g
ePkfl0gcCQ0/GQdhRhF34QpG919EOaEpbDCVVxdb6NBI3bIJKPGS6pgPT4U19pR+7gJRCIS+WGxk
el9oxMUR/BQt+lh24Gg5EQWIMVH1kgnEpUnbYFS7I+urJ1fKJ91oMvI4NJhmLGLKKrAWLf63sveF
vh04i72O+ET6y7UoqIC47gvtT7bVddn+6CR9o7DXJPk2iTVaJb+hY7xoIL/Vgv3EoJqwrt80ucif
nrsXdCTkUZyHkbafS1TDoDqR2RvqdDnAb8+P/vXtjqxLouPiJbMgPwTpHeuDUFz8iAmBMrblFLdP
n8i+s47vgbnOSH9KUB2B9rsnXN40LD+i4mgfYM9BdBVu243xHjZ/RDfBuYOheEAmFq0FJq/elCZ8
9sMEjmpz6yCXpmAT1/hFpvK+3JHGI7dWo643XNxiToaGzW8670cQE5Wm2LLrtxr2z6L/An/XMq7X
XSKlXo7Zo9iPXHU7EzQ96110ALM4LHNIrtkN84lWpPKIqxfXZIQ9qgJ5P208PIslDV3csCJ1Ysd9
Z08y4BfcLCP+D3XuSqpIYxTJNpPhWSWMFqQS0e9OyFfxwICEC2UAMoZt6ai3wS6G99WsJs3WORA7
7Jk9esG46A2LRqEJG15sWH6GLq0vKUMaI6pZ7+i1D7mu+Y1L64gIi2/tB+HycQXSFeNCQ/GFXd08
yVjSDiBsM03AU/vwvClhRlGeN307F40dhxleW9jqjK/UbgvwRT2wEMBl7MGm1mPQEaAxw8GV7EHh
D8Ki4PNdLygm0zqVS2vVOuUBL85SAfGNvW1jB7BILuQi9WcMIp3dsAGjRNu8F71MQTELKbJv3zR1
9Je9WRl7hxBh9B2oxAb0n27+vBaInBcVi1OWs4PARThFx84V3TALZDE9ncMW9FihY/EbkdcglIKu
LSyEOdAvEONhYfhcyDVkXn+Vu2vmbc2P0veOL7lULwDsFMF0D7y4swkRiXQzVl/oN2MZgHRg5jIM
oshZTS0ip9wbUa/3la5wQyoliAplxCh3v2nSmM3mCA9QadaI2B6TqYHn2IOZp5DUBt0Msh6ovL2s
NnZiKsYYSJTPlIGaSGep3zESE5FfjS0m91mTr4J+5dS+gKSzqthqGSYC8Tic63bvwrXds8AH6nee
wr/qWTRRPDFjxeFpRt8YKBmb2+UfPyd73KKVLNuzv/Tr7J7YcQJhVpKlP4xlMAlI+HyN0p20webv
x8z/eE7OzZ/Jlc59EdVzoTQtDHh3Lms5zuBuIUlt/WsaAf0DezilRcltSbOxYAGYt7GupifaJPM7
stvJ4S6OAV+xlpvZVcUyGabL7AkPOX1mjSj3HbjtKsJvDzN0NJRMRqQEw6HKZfpmtDCaLUOZP9l5
01A32ZDt/GY3TNW/n0MP7zsoMmoWf659aSucoGuYQ6caop+l0egRe7e7fGNO0YbqqhbzijzdmOgf
QtFLiqNgCjasJI3ai8RZ8LhauG03qgVhd0z5HdtVVEZ1Gwrc6zegMTlLLa1OV/QZtB1/l+XPByGe
irrxydDiv0I81YTpLmH+bbrbBlxssQ+OsDzi0fx60V+40y5GlSZFgZrDcWSP1oPQpUiVeykD4t+H
2RJg7r/IoNQmIrPW9diQwet/+4Efmv9+dCzNLxSqS8ugNOzejJiUZYORSqi4NThL+p0+NbQ+m1n8
gowFaHyBgzoqJxodeeGYyMt+6x1ZwoBmr4gZRokwmOOUaYT+dadpaQJK61PooB4Y61cWdvPw7JE6
tuGrV8dIt/Hwb9xwwYn9IZKxOpFxuOTlhRVXjNNcUMDXcyY9q2O6Asj4QswVjLiPY1L3zxrtIXNi
rr1gOimffGVHMeI1KEAAQdl7NcvZHgQeZ+bV4oL9ExWRb2F6lDeeYdVU8ND5ZYquFgDe6HWqlVXx
+hFFuLln+8N+fXUsOpUxJyANUMDvlJm40S06cJiCajQnl9L0t5bHh76gGAOaTRNwab8uMRMjJj1j
n5vEpoF9U98zSJQCQPJ6O3pczH6eA95qL9pMMmisLzFX0hzrMu6Gji0MBlhu04b7VMMJblj9ZgyB
WzkHHVILT5mMWb9SDeZ0CNIbW8avaU22op5ornwHQNZLLZKoeYD6lqXB/7Z1U5Qmz0o+ysp8BiNr
0b60LaXAsX8AcCSi63wy3B+ef9xh6kW5pMQiVePGCYulF8bsZ8NDz6gXx26w9loIezzFW0rlKpPV
VOV36pPtgLFAbv6yqxD60LMhDkFfexvE2vdGtovW1xWAvzN83PMIVmKzbmXG2UJ65CU5uaf/qbsS
M3Zk+QxdJUyHwdvjS1syt/ByenyGLFkoCydiQYSTFqxHzGkjG0UDyEJGZzDmhkFsPUVsLOq20SJ2
sV7SXcSrXDEfu5Bi0esZvuZIGTSePbXfZR5AdzlzKEQm+Xs9LPGy7lGgKXW1k5olFmayaXxmInRf
9/eFXSvI8Bsuy/XX132ojCtbm9s/re2RjWmHzCek8jSUBgYPRMsqrLnf1t9rxBnfXdvYPTZ5iBuq
MN852Av2dLXPSEfnTg5HbXU8SuiF0MDWlGPvn6emFP3N4L1KXmuGfKWLVZjOIVbRcqJHYTrgb9KV
+nGZxW5x8ol3J+yDfgQZU4cB7L37kfQysU9OVvtgAJMmqF/vL+lS0tYmYlkuMfng3Wfi4AesIr5K
C7XacIuiJfiHg5aQ2XKIbwTvTsyG8aqjyh0XXK3Sd/WHRfKLF7C1rJMuWqJk0IZ0yM0UDJrNDugC
OXZtS+pUji6REiZaZ5WBEtsntjHH9OLgcy52guyyi/1SGCEKV3/pOdYTwG6WO7SSjhoMLsAcDVGt
r5GV0VlfGdeklT9OO54f8LY6FpAtl0VhzOgbCsaunwpMojz9sNReti8GSkZFmMbXgTBAxVdIMNQ4
UKZZERslZY0kMb/8WY7KGNrkPaoteQonnYQc3dj3rvksoyUAF7LlSac7mOR1rUHKaaP5E5E+TJPS
EDUi9Bkh8XSlVsyKDqX69GVK8VrSBRrhibUjHwgH5QJc5TGzm//RS+x3y8lj5Bk6L5tx6+9q1SEl
WW0Bk4WEiEp9+6FYrzkIck+/AIzxEDRdmX954ajryhSgK0yMK1xcvQjI9ryQyeDVIW+zYqWcJAFk
k4yZFisTc6+mEyT3Vv6Zs5sqAdknoLReFViEH5RVkk8Do32RJY+xF5sKcSc1rOluGGCTBYqeqcs9
n8ByDcib1zTW7oaxe0NpLs1Y1hYvvHujFZyfkWpFwigCqCZz9pwhbOrkRUWYXc5wBwMlNJrvw9Ke
4Q+FjABl+E1Ce7vKr+LhL9Wd4Q3y1qQSdULoZsg4hkBuJ4Jzh7S1/VE/SRN7jvQ5aMK387Dp8wKa
f43TAGiBfJW7sOJsNW9HEzUqScdYpYOp23UmDcSc7HKR59X6omLlxcz3EIFA0pDBS8QuTnYxljpS
c7WcWwYcYtgG98M+HyqJ4AoT5qkgjB+pSPaF88ww2AX6TuUX8OxOEhhefKTjpJZA4A/hBEDxlq2N
jtbLif9HniUlgUkvfV9KuedDDM5dR+8tNXbIPlr88sRTt29kFCYC7zQxL2tXySk3+B5MoRuno4yr
06M4SfPgw+lnUSMT1P1KsmYQT5bzfKxgEQjO9xkNn1vIR1CRI3fMqUmSnKcu8ggyBf+GKG94MOXr
Ac9w+r41nbtRRdAbnv0Wg5KqaqFOo+k0qYTbdJyQKc8uNB2VaG4EH5KN2Vc0ZLaebU8xRJtDapnK
o9retGhpKRdGByS7Ikp4mSbqUz18I57x2GHMhYZdKShdv6giGanzetpSxIlnYK8dyZXO1+m/ODjM
gf5UrBNu0BWH+2k1BcQw0O88HjbScK2MkdCZf+bDbOrdqVTElo4IwY2GIs8mSaJsXxj9qMydQtya
4GeiybvNNrRY2iEZG4FDiDU/OU2qN9709M2R7tkuASubFHW6Jrxd6st2UHiVtoKV2XfcOXPRtBNK
WENTZzcj5UGj7CuiuIyovyNrElObJr1fkcxTUTrXWbpvwNSMhRw2vNe0LV41cVpkxKqg5dOlAno1
zkgDHEh9ZtpcuzyeEe43Myiyxs12LamkTs5GL8booZOLFCRf3z8nyGN4hfuH4wxqylSCQ74P27KT
dtXEUMeuhg+UmKdnKq8bM0eJH/HAfdaiRKGrK5zXu1BFU5ZZ2eHqS7sRqCIyOZHLOTYn7QwQmIYk
VK9fBW6RjQLyFAx5kHL5EzA7WeHqK3g7Xbt7dMRT+U6hTg14jfcGxDEPYT+wVgAJ2GoPasvwPH60
nsbEJqfbUYKSfOri56n1VzL6YMT9K6KYsJ9jC38q+OutZdIJzBqNwMJ5v5wAsbBWmCJhP32ROc5H
n2W0ZuFLt2TrGGY9vxQrj5e4uOVqovKsA72z3P2ApgC8MvLQyVEhDuRlcCH0UoCsbnp7R49HS+MS
Yhewo95l3EPnz/9oVRLHQ0ip5LW9vhXWixdzDkRKoFxE/ektHsgLxpJWWKEViLsRqVK78OqzXF3f
d3a87PMmVqm+akIlEAD30yXyU7sScwtco2ZkyU5UHxhFWkqXuiJ0qMZlxDND0++z5PzUK84eoN2a
+pQxaQdl4WPxJpr9H6vptSPe38bL252shtfXKDNO/cuen7TMcND2R53FrJdKfrcO/XNNfbt7ZMcC
+sVs6fpOxMC20C4gc27VHNXfYxh0qOgwJYnudlpcdEgC9HgfV0ZVs+Fy72i7uDWo8pki/qSbYPYB
161S1XKfvcvBtpKBb5NA12F4kjiv02jSl/dB9Y0JcSCojh+53nm3U6vAuiwITmWw6G354bWeoTQN
FFwpgqjNmTIBR2dWiD7Z8ktxgtcUyJSSQ17M6xQ9OQJAn04y6XHfPJrcthB6NheOHEbvwzfJhztd
s11dBA0nqdW5y2eTK19rLcTMgCEhz4yENoh1H4sxSw03FV1DAEMcEL0VoNhclD8LeVk3WCgKkBUJ
2BW7XHvHnlpO2Guo2KjiWlE23F7zFJCgG82mkGgVHmEQ0AVuMxha+nqO2/Mz5NLGysJ+jiQYIQs0
gzmA8fKMp/iwhznOfdU+Z4ljsxnZ/t3FKi5Bo3ka776dbfLcI68VOjVpORPeWHi8BHWaIp0dmuFP
I+OnFQN8IcaYeJeFKFVdN/GltP9GMbmTFwLdgpZSVlq5uvtKSFiGje/i5uTreGSoRJPYBpNY8mm8
1in1TPmgG8uf1utPTL5JxyMhLKb7aeyMTFOasyBZY7VGJPsgeqoEc0R4CauUKG9U7N8H1i5B3K67
LnSOsSz4CEZsjyu8yP3YTsQPZ/NqRZKVmH8xpcVG03P4QQUeg7qAm1pJwDHvR+MQto7tXAY0aB5e
h8yrmZVNOmrn7yd4IQ8O+xDUSaEO0od23lGLF0jhKwY/fwUCe8xZ4Fjj9XcvRYJdVufoVj9nmi/t
EtMBaB0+d1UnPDVRV7xUnzrGSRSeGA42z4KXEUUiYx+pItXNPOgUJyGIJtYydvWVmAjugolHXOkF
8KIZtuqRQAsbPuMJsy0IwW1Me03pKc0qCIbhrC/tZimV4g+hnWIJE8a6PFmFKZRc4Wq94aVa2HeW
LE8TTQWzxo/Uv33Rmz5i0WtWmtLlmp32AmiFM+L8S+/z3osnmZSRYvQph3LGvyKUPtmFtQ4r97pf
Fit4KXxooyBHKbvsyims5RnjAs7WA++yXyu8Bgh4/oQQ1wz/EAd1CKj6+JOlXyL44Lw9NPQTzPrk
TKx2mQUaXK2x8TtZyPhrwq13ELSsYGvRn6wRYnHhoEvXffhZ8TG7b+BxgJFCJSHgCGJZBpcjewED
XNGtETq38orKzhd+aYUzLuattOqRwM7FnTamY7Gy3BJu9REV3E3az8e4Wy3lV+Vzzd4ngKbxwYm0
wckAdFp72XV5NITT3IDJWXMJsqJ/F2XJezpcgaVn9SkX2Jrr2qGorbeC1pUQYzQe5qdLff8f7e5H
DdKenVGc6qJUg15mCngfbVTz8wOlSKvQSEPV1OayXjcnaHYN1XA3FfxM1yNA1eplj2dx+jOgPyXy
C5ZfIQCgCACm1nu/ChzOcrNKztHTj/Kji7x3Eiyk3uX1t3ANFYFPBgm9qn8ndG6AxsBY6uk/87WO
k06OyEeim9ZbNTERAVemSpprKAXXouGe5EI8KFxFy9SI/p95bWVMqgrcD+HT+j/zBhbvFx7fDThg
ChObJPWwgOkRBMgyiKYOEPw0llQ9k3m44aDOt6yz8phrB+zVvbkAPq5cRN4aiu2VebfaYtHFN48o
8ygGKdc1pPx8DBPv8Vz/AydEsyM56NGGOjV+FPINGiY4CeCoHi2mvaDAET/EB4YK4zHVAu1TpBIS
LmtgHSJ/+qINnNCNCFAhJYEmzGq/JxDe8FEo+WPvQQh/wGGxEUPL+rLXGFChV/JtvGb6dYw8E9Fj
I+JbxLXcSIo4ofKHQPPlSggEax5uFAm0yAALEH5cPUrsrl5V1PWELDQTije7J6x9E0vzEO53+ymm
z2tCwnip/pGOnVGnQM77h3XddIsS0TJObG97VF10vuKBfPGrnUgKSbFWHmp05gKEplCWgEA4QjvO
B0mssxMnocQqatY44eXgnoaFiW7vfSiW8wXeKSuu8iadmUNq4tG3eah/89mDf/ZVn0Saqhp9RomU
EIn+ePywTKRRDCEND69oWPNJV2nOcjl+He2k0zzHnzU0xhI6+3yAkTyIf+IM+QulBLt1BoK3MIz/
G/u/gTcQHhDVuQVHnoq3E6B3qpAW7QBrsA4deM+vvv/O74Is4FkNfIYn4H6GxiJgfIcWXwAkwgS+
mO2uMCw09JF48NMl0vCzHDZrMNHtI2BnfrrtYyWom3EvMRIyVGf/YLGtzJBP58v+TofTkuQvniz5
9VhYgzZKiWmqFPIu+BSuuMleXAS1u7t+zgLr+dAPZ5Mw63kYyN3FFNdfQDA6QEDk8ulN5yPldiP1
rs9SxC0z0JURn64okqWdHx/GpE9dGp8+Jx0ENbKmk9gnbMDhS3i8X/1H3krCbvZrGtX7Jx70gsi3
EbUZ01xvT+lQ6/CJLQZn0neBhOuCzkkOSAIV5oq2FxrRFDz57qJJvFSqhsfm3G6UN13ofy1vduHD
RBaVMB0bz4WNpdEgMvnGjU+1iQ1H9PorHK7tPXHV3bibX289zKgYRTyA1hbGI4eNxe4edNDQ2XlI
TwhO0uO4fZcclTwCgoHyNApaYslpBhThzypJSqvWXQywj4un8QAbKXQF5QS9+qHSYwGDOHmDGvgZ
NXZefB5Hwn9tpZmZv8OB4VoC9N/7hQB3UBXHHu86FwBnyrOhD5Fdek/Uz2qyUAfYerj7m7Y7Wawf
ygL7pdCkmUvcRaS3XEEjK4wFLoILy/wjHYojDNRWBo6m8zteR4EGKck84a8WMqOBfdf+sFBdXZOn
Hknw2OclTzlN4hofq3GZoEyK2Zo0N2vNSXftt5tL7pHPEL8kjNNac48uqbBB/GXsCXPxXuKrag4P
6W/97q0o7CILVK+Ot55szdqP5MRKjQJ7Qgx1Agew7+L4iBFOCKfIrCHfKxmbFxDRd8jzlFIAkmnW
GNxnpQ3NUACUrkfg5oyUjjGO1hoDPLns/kytLF3yLy+l9MX0mKZh1sWt0L1aCSABr2LGzBzJaoZ6
sF1y+tk4WMMcXXAoh3C0YgtYgQNiUQE2v+1JpLap87aYar0vBNPkWZPyViS98ttWyW1ywpHOnOzF
4kEd1a7jh6r+9at424ab7V0peN5MqwjygHhQmVjB46NKqSH5r1GQ9Yl74a/Og8AUXDyzXkXETh6q
e3zx3sWxEqZLZFY7lcaIUNAzZz6AzZbUl/252Z6TTniorhAFSVohWn5NFgsjBdFNx0oH4AfV797R
Qk84wMchSF21C1i5KyJUk/lygPpp/MnCaSrAFe+K6dqSeoTNMOicjPBQeviQkc2v1SowfCY7MAYN
9YAshRAG9gR9vJkEhjvgfcmJjyTL2kSjt7Hw7iWlg8dyZFg+/OxD+P7t9opz9ujc17QO8xflRgof
4rlW9znhBVNOmeJkfbr1NdfqK0SuRfwLG495PMnLN04aJeclHSfvo6c/zbs3Tl/MwQ11i4LuI/77
ibNUAcAJVOy8M0nsulRG3AzgawvWy0R2WsyCPv+4cz82bVO5PyVVLg7WvmYKNehElWD/Xw43imc+
d3Conj9MQwF7sxkpO3kDacsgQKE6q8a4M16lKNXD1dGN7xyzVm1ktWet1TxSsjyZbYl5o1mHaPZR
Tz02b72BuiP6XBe6r3zjHJMpgbO3B1C8i6dOQwFs53MpK59R7hdCrEue5E3BAJSB3rePndLrI1Js
ysmRZ4WwBGL1sHpwsai9jQL3J4pZl0e1KjzoFM2qHfAUkrypIeNQ9X6N3j0JZ1TDq1YkkWT1mdQj
llKDw5MN5l5hflReeh2EAVN77zanBoNj5HkWJpQ5ljRG/gkDrrk2dltYflFgQswB7tDiEAFhHEFt
wOURMqYrHjZZ7xMt9tTnYOdhwFe3L+b7Kiv8d08k38ql9gz7GdzxBzr8w/4yiGm7kePaQVymFOLM
uadaje3fnUGrPoxNRv0k/ghfcJS1ehbh3Smn6Wtj9DiIp985mX8IEr2vds96P+FdGKa1AXyBxGuk
m7QHX2bKj6y2t7I5yV8gysfGr6sb+x9hmY5TT8UCmQxbAbzmRUsV6mSmPro4EMIPJBJq1aaya2sV
DUvInAMCapBdgR1NreegQmEj8U9nN7klSOSJGTqDMdQPTbTwEfsq3XQw28pyCfroRU6SOQf2IhNJ
s2WbqoDxWeXkOMYMc0ahxlrWDXPpcmCEQtyllhSysWmanc0teqAXBMfab+77JH3RnwnRXUJ97Mia
gxubnAxdJPg1s2CVpPawZIraMH3V2AntjXcGUVXkHKIyI4IJFlK5D0tE37xFXnTSa+Mxk3vAlPgQ
gxx//yUEhjyq0mB0Xc4QBUTVhURzUM1tqoaEzbBTTe1pn/9HZwWSn6TV9tfxWgS65uQuLHiWDMDy
X7QxbOKFWmWdsqEplCucNpSZY8ghjKsQGC9l9SKhJP6341tlOu/m5m5/tUkdHnhWMzIQAczHc+oE
EFulP50k0j7Dchs/GoEw/4952Gr0jGyEB/AWQp9xgExKZmLK5oYS6nqMurrK5eOlv+gnvTb+q+y1
4JjDas+BtRKErtEQOXASmbiyNIJMCgy3ty3rUP//tstyVNqZ04/CkmXOm99h9KqXcsYA8R6xBuKd
zce7DejCZrRkN7lAlGKgRGk0ufzROjL9XUv+ybdgFzReWzxfgEyROvTPp5ZJJGjGkHIv6L58NUYV
/fvmdggxjhlR7/MxflgluIiLynR7RrdxCvOLMcDXl7VqQ5SEbXR4euIpM9C5gbxUyDJPYXFzjlwl
xaosFZx2Sdd14MlNCyNSulGzf+EQC07BbSN5BxJ4AokbSdQWL0e9OrcBziT00w5AdOoGS2wXeSU7
UTWNuUdranYesAuyCpWu0vaDK+pPwhrbJjsuyu7YUTIs5CDaamdVgiBQAk5fE4evWYOL1FBHAy7c
Xb44KO+6T8KOLW4BBAw0bBftt9NOGgEjcKCb3WgmHvcQ/zHizH42wjIq43BvRbWsOTbMg+Snw1DY
EYDUGocFLD3GULT5e+EfUnSleH7TxlHftfx3bLpay6woWaQfSCkx9c5+m7q4jL6PsLusO9B0zqQ1
EIMknuyEC9PS2XRGqhFPldvouDtk4mYuZgrAqrvJiDwoljmhWLvpL8bpoVFdqebPDJLUJqz3kEPr
ougVv0t2S1XrW8zG0O+PTSw3NPanp5VsdEFXwxQM9O+w1s1WBIYaDKGDV+vKrerwqIw7bgYDdfSB
n6cZc0D0rnamUtoE7aSk92m/ovCYbghPHCXsDFRkNVN3VM9dQYjiaZw2VZr6Dn+nOiubbTvYJSut
8jPZH71fBV9D7y5EDbyuotNW7GmQtAxKz/yVsoclpAK64P7PTPkG8E7MrwtwPAHqDG/kcwU6Ic5S
oZua7o37qVpJ4n7mUPiggpomEzN1lDcFkSwzVWEz14F/YAlTcVEpT0+Uap8p5fuXdZggWJ9/MsJ5
kyfGhryVQ/JM5SiIbbUzomjQgx8kRzyCzdz+p01sXYSygt6+9MJUZiWuHinPQvCvQlSM1zD02HlM
ZXyVBvvOrOCX9wbWvtA6yac3jBf3W55nqGyi6xuEs2lM0GJldB7oTyRO0UibOuTk0wzHy8angpTe
O/Xtl+Wz64nnN5H0t0t/dG28voqZ24oFffRq36+/fIGi/sdBWmoLefEC2w1VQ5f5qmq5ctKVGTp2
U1Abqs3BBo7+iOQGGb1aas3kej8XUiQ44RWBToEGGwH6SRN4Bv0+XnGAXleJpgoD1FJikJtvPBo5
bKJdf76G5182YZ0ftmb7mvSIQkSTfp1/WuKyYI6z1ry9SWHade2f/nrp2IkqLnzcvgIJZ39V8MiE
47ZClDyEJZoqU7xEfB+tgkdVCoI1sUKQoSmhNKxKXYtKdZWg4XhYPpKKjgRayMzKF4wc0d2GbO5a
+ZKtWut+XjqDeXF0BoMlX7ZGdIGeCWSaNYhKkL1xkFlMrE9k0SQ8DhHYTXGfldqTbSAhzqN8qC3j
9bxPxkmcM2K/TfCGyTufC4sCiVAOe+4LUv42gq6DpwOBA4s1MO/Lht6A0zddPXIfEAJoTFALjiHs
41no2wlFoDriwTi6+v+p0Op/HyuoPBnwmXp/v7FQyJVTbUX1GgN6nT35Oa2/UhPLpomDgIoPpz7j
oVZO4eRllseclevUSu40/v/wRsnMvXNPlbS+j8MBrKedNUfFgR6KwptVEot3h3UMCREu6hPNITx4
1gyLjGdjVgkyQbkpmA0BM6+phGmhBjVUWdLwxgL9Qr7Jtv+A+MnVqIy6A+pCFUOmoieoH3LEWbl0
eOkz60u6qYcYyI8HelokKZT9gUEP82rVGG97qQLTiej23onuL2ehIokk7b6GUJGaEdM+ss1RNv00
xkZM9qcq2bAagx8LMNNWo2lfibEts5OWNrPYQ6yx3QLzfwhTf8rnUFrv8PQodYYnorFMbo+8pm9m
Sv7ZAok//NLD+AdTFckkv4dfjUG5FX2sB/AP3lfveVfC6MFl4LqdTbGaewj5S+dpuJA+7Sia+GxJ
INEHyp6wuKbDqsoH5Uic2njXhF6ndCWfVx8SdpbYhSAess958BPUQ419CgeLnSmQNZ58RlSJdizv
HIRkIhuloMZWgjKwznS/0rCbocLP0XEqxpRbGr5c/H9oFCl3NQvSdI134WEtdGgXxraCTEOeU+y9
eQ301AGLRBrHDDsmV4ROIi0nmmZBGTfqnbbeERqCvioRLts9wjWsp/LTZWGpqPxKrMtEe4vgceVu
MdmyMD0wmqvoIQPhv/O7DrFsOXZ3/Dr63mN/x+gVm41NjUfh9YIKmCwCem8hGDw6hHPjoDNwef6W
ICqpUGSgSPnyuxUEvuCR0kwobLTVhC7/ZOja4msbns04YDIR6RUINU06Kr/+oYQKaku+B+34+gtm
TAK/8UeTvH80hsbTTnwj5YjtgG56K8IT8tKLhye969AcYakcNpRpd71G43Hboh3QU01rdcjBtO9M
1h6jBtdFyx+t+FxFmrDRpOjZKQTMhpFaDDktQinChdG4XuTC+ojHp4IrsEcO3AAn2EycEHCF9KUy
c8PieAwVi0ABIyBL5WfCmTCpkTKNmd2bhWHZx/YQimWsf47LZ38zhbzQrantEEZo6BurOagT/EcA
SAjEnmMMm+OMYuTUHZvzr4oZN9nACs3SWkDVPibR3z0gtcT4LN8exlmrHOTXkgJSUxHlKEYsUPwT
CR/ZJLqjMvXz/MIQ0ocTLUvQQozfy0GJFgajKvnb0WObUuKco75WYkfUrkZNjhizn917TRERStAF
XrHMDUgBjVj8cuKs8nWvbY9HtreOqi5PvaNtVEjMXU3vWEMuqihBUQwq+SBeRiWGyLZCottc2lW4
MfYyEPLKyBl/LQwyyYq4ZfPUrDtNa0M7ea3frPrRjO7oRQFIgpxgcSoKBGOZioyqnzLpKUzOaVcM
0bUooaGXSKOMh+MiHwLKgB+HMfzLD6Se42keV848YxcplYrxcqE/4nYsrzMq37lCPpcxJnZYFDFR
CezTWG6Gi223iq5vHBM8XlpbXy8n5RSkLT88H6JOV2zJyfWZL3ayCbeh7vZ9gPzrACzDBcXHlXy/
Kp3U72VnSm0nyTLKWz1eJMgBj9Nbow5ryXzJue0L5Cwyr8t/gtkcPPdUH05/4jsXSBDSC+uCM29T
Cs9wRk27jlPEYmlGZrobNwb5dgbawLy7UyQBTKdNj5BTsV/BJphn+RwcZdqCSpUxyUVWKBJprgzb
WZdWFx4tJuQSS4QGjj0fTS5+qGisQVuTHSLbID3M1iUyrhlYw0/aUiBlT279Tzq7mPwymPOoOepB
sVHtmfBIC0xvjVMOJWOON4Ljo89F2J1U7s8XwBSGkqtqTMTpsNN82ZCZp3msTHbH6yEJtLkW20py
r1DhKHl3wfxeFXnJHeyF+ch8Fh6yYRhtn1EaPaatr7NjfcjhYSK5D2gdPX9cqa9OtmCqbDitXAvt
cb1xUgODSNuejUtr8wYdlRRYAEz7JCe1zgQqRB1FieLjZGwsx4GAQJpgieQOsqfwz/UrUyaCbvZe
HIer6ro1AfhM9MYHqvOjM2rkHNGTx3R/9ef+/ganzCqd+vXHM7/eLPDoFI5jKmx9MUTDQVSQ3LrK
Dfqz2+MjsolknExM7uWYudgYJLNlYUbu09lOJMv3ohGhx5Udr/bBtJTWNPbHmtbNTZASXeeCYUkh
S2bzBBMZeCOfu5M0FPD8yK0QsBaapxgksJ8D1fyro96TI/YMzMH7fy/Ws7ZcrjRswjdw6CSwbYXI
9CNZ6EW1q/4pNEE+7/pDTC4kvlUVX9ixGXd7Q+dpwnCdVlCv15xWQcHFsGhnIGgbRNL2fzLd9ShK
KRRRUa1SMbDSVYJvZQlR4TIcjcSy3elrSdSFSeT2RvZoYpSZkrouVgqF//TASecWqWAryXNXXr4R
zCDjRyQvuT8sRAnERRS/oiY045MU024IyLoK63Lb+NkjVd61R7EGH1LWchaGXDUhd6ovhsl/FELi
43bYRUo88R4ltCGPuG0bkY+Hb8cA7aHYPB2XnOk+ffLT36JrsinbYl9c24N4xqOJTVVCUOuz1Psh
rWf2e6yPM8znzp7VzzbY/cDGB9T5IswKYoduEJ9XppQLVeBPoblIG50rxL5anIP1mwItZXZgBxrk
WWjHz+Xs/Kk/CsrhnKQYhrAVYhqlkpMkrE/YkQXFDsLWiqU8H567bsz6TPUJX5tMwKwWJiDfUTkm
NGNN/CecYOXnyGYSJy4V3NUnANRQdOEaJivQhl7nkVfWoRcpFk1nkN/iZ5NcdeJ1KLwCZrqV/CnG
xF3in9wFrbjWKUwZ6F8WzOx3wJDPD2OtRO91SXMZOuCMTZMOhQMRtwUbSOoDQa5paj8sVrfOR4za
3R34ewm763GTorw4H+2A1bVg7BR+mQrVIz79Dp5t/fe+6ozbGm4RljtT2zLfhFgw/uN0JJoI4toz
VG3DSTIqviL9rAOxgYhDNIEGHes6jn6zAYiPUP4DRSGbUDCich/oNiVeFzPq2uCpJlVivUL2XEvu
hqGpAxPX/VkSrlSc4+Rw5pZq/fGHRzjs9Q7zNIR1g1EUJl6jnVn6Xs8UxzcouqSMHNs6+DoxUndS
kyQTp7aptPxjzqARh6iuiq3jp+Si7yus9E1ee5J8z3a11emrl8+Xycac6oIfKrGKjVoIAP7Q50ue
kG2/zCPlHOM3oHBWFLq29IaZGCItAz+j/p6WiwGN1Po4wkoB1GJ1FtFPxfqIska6zCBxSDAAzrsV
tnjOTpTtNIXS32md5XUKXRo/BEx6RKgm2R7QXivVPwQ3D+W6kPtKfwbSGM7o2jixAeHW+sqr4gb7
8BKABc54mV9H9KPIW8LT2o9ADAI45CSU+TFCXN/yPhjxlnFsHzXX02INfsecAZuhJ8yl2jamo//T
ncsiJlnRp966MCCTMLMVSXCSZG4zIStYyqwIBEWLQ1lBY8fFN+fkVNVr3s3A+If43v+crdvdVcjp
ZGPBruDn4PKHUxMqUX5KbsY33RuCIFxA8KFrLwbf2Q1Tky6Af3zA7Og4Hv451j/hg8Z/6f9Bmu0u
UdJ4wjyr0tctIaNh7xS3ff9mryffbcaGJhefXfUUuPKVzzQ4fGV1WLQO22SF4oa8zc/K7GomzbA5
wzSuiH74zEt5E4pJVgzdTixYgetdJW0ceQa//7pp2ZyfUlbnrWQnVwhTksspI5sigmQQfRDCLF7Q
H5ysciVd5Wo9LhLXCk/cEVrw+VZwiMewad6xcXhVMGExRu8weNvv6LQ0MeYIE5aZnEgK6ku4YhLD
3z1xk3+qib6iQyeHARd80yz/VMC9P6/BnjGz683BsJ4PoDQTEgftv5Vje8VQPtYQrdx1t8tU9eXo
T3LwseVHIdeTQRgqGxAi4dRFggw6AInmo/J2hvprMfAgdTpSPyzuDy1WqQ6xOQjd1DUyKiTgFyEg
oGgOwTpz5gXv8Q/saShAx7D2sKp8VEooFM54IiTgDUuEnpPsXaix9e0cm9kdQY++ODL4oHS+wpDQ
BJQEi3BEmvYzqMEmffFiTQj4oQ1GXHJUQxpu3QU8h+IzMRwh/KQ6/tHcdVuiqM2dVUF5cfCxoYni
zffqbK/cgX3O9SeEtynQdn5ozm7vJ3dNX2rehxO2U+9g4c7DmTR3uVyzJewp19r8Ht1xbXFGl5sM
2RGqEZvz0svPpQB5MYqpzzhVcfdWll6o6O9NMxnO7KJB+u9SbVgMSiXQqUcbQd5yNGnYt9n9kGHA
I1Dwr/e0Iodmpbd1YunsN0yHglcK97zdQ0D2iwofOI93Azo/VqVqsp5axuyqDjWGSOXSKfR7YkUY
uuTuYok7IT6SVcRHx27WjcDcbEZnZDPRYVqe3+U/9EtveG272WMOpkcnxYSH99ROav6YMk+sivtU
QbR+SPfto2q0hQyWlthGJRWxmSkGNp6krJLyuapiq1B2D3PzYbCROqo8qAsaInPiTg+O1lrNhm6u
nWbprE9tTaaXgmugcdzD1p1N0fa8VA7BwBLJCRgeUi7kHbvONtfnKchESeIVPiKthChxBlq6KQFq
BXGZEjhzH/EfIrQQMUvMOd6VAOQYFeELLRZd4Y3IIs8AOul/6zNWAdptJTs2J0C5tcRQDduezI8/
bVnpO4GrFcN2LgcpeyKliM60OnBSFg5eiG2p97ePIlmcH2BStefehlGV8sZwbijXvJfPc1rgAAtx
ZOUE0xE9/PYw0df9jRD8sRn5tO8CoezFh2vPjxLTKXM8VXAIRSJD+AqVLMK+LGa3doL7KapxQ+CB
4lGJ/qHtLJha+fLi7cqyZKd+HAUCEaj55o87YE/Ev4BFZzWq9k7kFcJFowvkqCPYwLX8lo6aZJ86
vlXf/2NOgvSujKKqbze5K9LA0tLpuVkVzjAYoCdDfRx2FHUEdTyI4PSUvMRVGGdOWbtPTtUo35UJ
Y6SNHJU3+CWPhv6QGJTZHwjm/OXvQ4Jyq/+dahvdXaaH25gC8+m60KAhSJrYkFJyLs1bv/v50CSO
qayAJ8gBS2YjuDx1lCHD+qmuXvzOAF29gIaKj1J9j+vQ+iDmDott6fdTYXWykX1RS2L84oZKVYx2
zrFrEi1+P3lBpEWd7oYSJ0ISGL66x8aXheRJmFS7JKbUWysE/JPqcvLi/QN2RuH3AbqIXeufiY/U
c8JoYQYFRFT0gR75f/IPxKAG0iOlu4xMf4dRXMvG99jX3S6eyPhjWGH1VOhbdjMNb+qPeJ0M+Vrs
yX7NFPYp181bD4hrNgCH1e2b7LdiXveZSIhscn0VGocRDilGY9wAmoHNrM/LMFyKd5AkmP0dQd2k
LjxrCWwgrohSXWgBGnXZW6/5XNo2p2UsGCtHQqeH74ZWceBplsFAXgCF35o+KyOLOADjLlICf2A3
jJb9ZHy1jMfeNjSDw/hnxK/7ldR3CnMVGGmnigtlGst0LY49F43bM+11FPcTqjDoRfXS/a/Stc/0
5f6ca5BHwcfFD1m9MNMitpMjEkSH+Ivm1LgOnFCigHxX++YbbByJvBLozr001tk/EFgKR9isPMoz
6mUZF5tPA1YS5XIA0M23sx4RmbBySHIED1frfxK9rnf7o14oip90E/3ta/DW81fnFyfv4IW8Esnu
JRXSYIFhTuCpM6uQ0civmQ/Pt5sCNCogfyxxwhum+yeu/38xnxzac2KhDKTYLA1mKj5VhD7p5bDy
Mbs/Kfa9cbWjlluIZorg8Vxh4dA+mmJIKhyjgX7tsWhAYsWw3+I7YB07PghLUTNN4s0J+lAAu9nz
tLlucRLtDRTMxHDxyVYbpLJNGv5qXU5Y4rN5Xlsi1g5L2uH4HOM3RebrvUgYI5p0d6UqmvZCNRiy
pPrIVSS6KZstReh7P4anw7W0YGF5cn7Qkn6NN7aUw7HbGv7fDDe8PdP3mELMROCNjk38ba6pUz9s
JIX8O/ZMzkI6wdRZXm5hleSjjxLV9f/6f7FSi3Gj/SoI2vqfFBvBj4TiHdafvf0XIuSVEzA0qNHd
73N/mZPHt5xCN4BqcMAyp6+gFHOcAn0rBqPEmr7mKQnjed0f+mzuSpiLqvuEbAZ58xVUCDzXtDhE
ZdCe8UaFa6A4pFxigmqTox7Q+/0FDH0EsTjqGVRl+gz2NhnEvib2uItz4Q1GCI1+IgOhUda1Lzuz
DcFL7YVzA7kCqhhHDQsKjBddih0vmQMUbp/2HnHpncdtT2fVNaima2NCFndI1m314FXiJrPh5Cml
etLRI0So6Xm5byKSr9m+HUfyp2EgxxYjIzjI2L1K6zfSO38zPL81EkQ992ocXUDF7weP9cdM8wVe
oBnJQQf5lGmDNk+4E+cwAV7IHvKuTG2/lp3e1qvBJIEE3KsC39qvGl1zVyTPUIjwRkZpKJ1sF+df
9lVQRUmi5rC/9GzP2BsvUSZKU1MA+JDKPyboDQ48mBXTDlc0f+1nWKqAV5ba3/hZarvoITkygvI3
A3rb9zXE/qwwCy3+NqUmpHvisOmIbTVMZTf9yYNfb0lac0PhCOiBbI6IdfMb5AAVkwVO9AMdpjYc
NGJaJOGoOgBFGRZVPOUk1JzGurHNdk9FRwVXQJuV/S2laKCLIFXIv9VfVgyd3VvtIlAXwiAgz9P5
pnD2hwVWbrPK5wXvzkjqz9wv+nmHUycgwBHdbVigS5q5ilYLNkcpBiZM3FHdBU6fv5znnfFEU637
O/TCyT7Wl+fKZbhlIDiC7aClRjdnEMZHItQCYgjQU4fW+YyIA040dfqbf9j/XripAiKNngFS77b9
d+vW4XQm2XIBwUSMaGa8oIykTqxzrzdfeMK1KC1A7na7/3i3fljgKHyEtFoWM5ciE78Xd6H5pHn9
+ht+zP+uyCdCme9A8z5tkzy7Dv/bTwVFIRR3ZVgoSpBWdKy035NfuNgRVWqsNTkQR9IB9B5IKK+p
pAkTZNysNpGEtmmBSyPNZs7fdPSHZkozXDh0vs9OW3KiyWLJxptYQJ03nGLlnVSapOwcYKk/Aumk
DgKaU3X0Bv2Lfw8tWheu8BPkFFNpJzpIkwwgoruMWMcNpXdpHCqdeRhfImFKBKeLonrhrFmf5Bpx
lTHCkMATQI/KNxS84/F789gunMtlStVtBK3JlFFXkemuJMFqble2RffuVK4O9xJJiyFUWkXi41Vq
cS9MIIwhS6CR0yG1BxW9CdquiDHJe15YWoqV3QIcrCGZbjQ0afiEVKndvf2OgLjPHZ1nwDyws5GR
vE2dvnzS03+09jnxzqsNEyGE7PhGzYrdhBCbygOnt1wJxCNBpVewu+bkaj7f82y/etgTIIdtDmx8
RZbD5tyFLBWv++DVPzXFz2XJeChWhiQDU//KsxMxq+Gzg+01kR14x/lba0WJDHb3UcU1d2q7y2aT
tuvmpZYK9E+ksXCoDOvn+Y3y7mXx+SmKq5abs7rFHD38whuVBcVCv5kS0/zZ5ZLIdkwKg9zgrZJ7
xH65q8LvSPPgQ3jI4UHtFesNlzOFh5f4EeEFh1eZ4GjSwAwJKlF/ZY+A5nVFQtJBZE9q8jDXa+WX
nl4jykWvDIeC/guVJApHy6STv5EsgmVn/PJiQloQrgDjDh/+QZlIhrzZ0WiwVdAx1AzRaZrJ3cei
Kvucush7M/Whvdg8vK/K5bf/P1dWHqKbBVBliYceLh1zwCmVZYXJxc93ex+/mv4h+SwjvAokFiyG
chac9rBJA3mZHg5mz7kiI4jmdLDuVemxJrrNtscumTONJoTqqrnd7QNLMIEPaIE6WSZLbjDpajuI
dGF7YBhs9lyJfvHUQjTfgd9ILZgHY2stfsxJdyblrky8Wrn0qc6ZDgIzh1u657l7pFzgdyXdKgIb
L8mlOcnIdt9XGp7WNYaF8/ECrDMeG/kPNaPMu2ELbxXr3YexHoXcBNc4Xkrxl/hfZ6fTN59nBTy9
Y51RbiJhj5L3WB+XAwdhXx9ZjMoSaaQCapjakNxgdPnXc8qAuNX8M9M124FpPNzboCfb3FTCWQuS
KL1z8ZT3MEK3+v9qCXyPg2IkYjdRSUQPw1bfU89QZziU7tKccehf+2+3gZL0z8+thQr+4yyxeP34
wQfQQg2IIPrk5+v03kvFBtvU3zBGQGRD9P2hbmEKzmLBf6kQ+m7cq+5FvrBoO5yZDG0pomw2BpG/
89dvmEf35A+C6OX34bfE0pjPNwiN1S59pqSu9wtQJdms4z6pUKo2zGCS5iI3i4eVJHKaRAqS2BM7
UPuSGn0DXutoPZT2z1/TYspojc4I5Uvxwmw/2NYaCyHbutBK5+YY6MOp0QyeYecfPn4FjReM5BFF
C4wQpymPCy867A4PcaHpdpwOIXBoCVbz0B8iWkvsIxQgUX4EMhfZd0wQkGej+qVMpyhGUPkiuY7g
VekYzoZI8cGnYxOWFi1BuQ8bL5kU0UwE2lSshFTTNJAvGrGCEXkWatzKG8Pkh5VgKZzG0ka4CfNP
h0wheb/PpmgugN2N8JrqQNgZu3PNPCViuOcljrFKKh7Y8u252WU9sulT1WkC9nCD39SGd+DzT8Xu
lWbkpGjGPIpalthRwlr6uJlKctTMnx1gD2m+lc6HHL5xux40JajEDLePhoqWUbK+NxUuKq9ZTyjU
jik3UhCPvTtgypCwFSzOzOLe7yeRKCVbUe40GeBfhwOMWjw3aeGK7ZI8Vi6H1sPOb6X1KUyOe4YE
4abjkObhwx1L+ecprEZYDDyyizuTN3KWisS1JBqREvR7g9xjbOI2UeWFZoo7J2hSa2CZ9tlYZ3SU
997mA7YQt/d1FcRnLydPruWbrcDvg/G65aBGHq0cNegAQYWGdFi6Sgx8h/QBY1KqNvkhlTFAuuWO
qGWhbfmlKBg21jm0oWPugObkk+KytTe99OSKqZxkH0yx2xlrtt4smj4x8b9+v/6+ZAKUejTCtdeH
L72oh8e5o/GwoHIRTxT6VApL6r2olVJgc0dQJZJJtKK8yr4LPFRmk/EWPvMUReXPek9+YqKDRtLN
dPKOfqiNZEbL1JJn/CaL92KCposdCXJDz9AEDCMbtE5Vi4H9i0nfL1GlNE+/NrZaY9CKVNFz74e1
wttXoqyQ7kxR1+OJccT5bOl/YWOzpi/ODBp0BFvwcEby3I2X16hslNhrBjvcnUHL/YqT7E5/w1Pn
6LpmQ1ubRWm3CGrrVyNYcvi0Tf1C1rr8dRSDAhcBzWPR4mvuG02fRRWeUuT8oG6sQdp4nGTpnzO6
d8bOkay2yk4NNLRLX9Gjabu6+l06aB96SZgK8IEu7EcOb3EP0bPICYxtg51rSCmkcPMngx7sDfdT
qiFjc6F6QzBwH9viwhkw3+28rzgEmADDLpe6s0dvjCuqcPh08j+p0tmOLxFfHu7BhVYOy7j0OVG6
P63kZEhILumSdyBiWIaDC/TJNE5gBc0d9hDpTbdm/sCeCpO+6w59EANw0sQBC4kpoKdKWoTb2iJu
5IeTDxTQt+ePcOLXdfygmX6WNLXZl04J6LeI0aurIe+ZSSdVWobLplaztGnYm9hfLTlN1pD800OD
NJoZpTAcfyG1DQeptYSc7yneX/FuTWcOM7JNT5dUtIvHS/XGiLFjLoEYrz5k0yYy5nQuQvpoDFWr
irNNcCiAgcNXQ2sPmr0Mi9muBqEVFZM5tN8D3i2du40Vh+0gny54H+PyK6/euhHukBpYC+GXW56F
X+Q6tkk0Al5+6kis6bno8WjgIl9Q2kIPT2+1staIlz9+Q62ns4jZls5L23YocLqVkob9Tt3MpBs1
wwU3fyIZWGlU58SxJPs49PBlzPQSQhzyGhbur+h3cWn4HqEgsalbihb5hHT/HGfxJeFIlLiNqKVV
BlepeTluWnKiIKoBP6SCj0c77MRRX0L7z8E3N0b/HMtNoRGJUFIaCBCFYocVIbINwOrA27SlTbpa
TEnKON4mk9Slmc8U2DwpxP+V4lJWuGncKDEAn79trN5PJVHK/eqGRV3CJhLz+0T1cnfTh7Oo7y30
H1mJRlKnSQeMfyf2jxjt0/M4hMuZ/29275nkLR+NG6K6NCm5YRbCWHcDVpH3i1L5tFm509h0DPBV
w8Q5yF6Ecg361gbhh3GiIbH3ExA6G+bAkUzGXoLFDwfQbTVNvCOASK1tYXyVSyt7x8eO7ivKgaXP
aclUq9UYpOsj7MF02fiM11BWb0jFNO2OaYDOEMaES7X+F3YSJpcZG3tx6JdZdfd4Tl7eqBrw5ll6
695RbNrblVTuCxNaKd0+1RwhY4DUi29UnLZxlC/JbePLUVgfJWT00DZy2Z1F3BQKK7MDmfugBZS9
IPPtg5UxwfVl4qq28btza2EDgYnemyEtj9mvJK/6npOu4mxUH/qZhSbQxsMGvDBVSETG6RLi7pd5
mXLWW9a9qcuhgerSI4umKu5CVAqlWZDw5BLoj73IghPPnovN9YghKFjdavwIp9wdlobRA5SJvLdB
QsN8iESarr8ZbF0nUIXfXKrmRkrqSVqWqww7j3MP/Jh08s6edMX5huyOsBcHuNeaqBKZZm9EtZ9A
v8sxEX38/6rtmPY7PCKiPLvGShYbafYAh8tsTr8MVHxlKnpBlI+XVy/QQWqycXnnlR2Ve+YCf9++
FrEcj8vcHOJvamyeaavJHjOs/N6x2AQ9pFK8UyOceadxsYfZ0chYiRHqJS5E5401fFq6TSessiwp
Mk9dGr9X2zOaJ8S0eYMMxOa2vqzwwxLcoA44K1mfXt41s3hJ2hZnxiN2kY+P8l3ihtOI3PVjz0qD
db45auc5KD7ptJ+YYgOWm4bJ0umYPwUbEZzmYYSVyNyiN7bYH4NfSIs/cshpVUstMQr8OMS8sZ55
j2OOutfLExdqt13bMcT2EDdqUVNwaG4ueGszRGUteg5Omo57MT7hPC3blA/A97XFQ6pFQydhKXW4
LjuxnKy7eRGRDVi5aIsE3CD9sQmZNt+PfpyDXV2eAf00Tnxsx/59VYBr3pBLpMsbld8c1b06wxW0
+ZxYgH9RbHrmu+prBslCsKMyghUC/luqLPehOWXlYhYRKBseYs3BhC7nfbUTzZuy8SX5iGQoLP/d
Gca6ZPYTfcwUJi75Y694PeTEnnLhNqHAhHH4H6iI/xj5aJKImU3O2vctkKuT28/KbpO6aX1TCaSX
8aQydNIsc6DCu5STpDXI4fkuWGZvZ3+nLFusQ2oLPcS0eA0h8doc4DS82doDs98kFPxI4FEuGcgi
EYUoZ44h7iHIU3tZ53u3+Op4QSbR0oWrKxp2x+hWBhCy0NkQeYpQnU16X+NzijLZ+5aHo/HMkCtG
mjCIy1ksSNimEmLcq8furHNnuQlFw0P1TOOtollDVi+0FEUafXy5zjCD7sThu2gyKl8LWDNXIlnO
ff51/TSF0N4gwOyqi9c7djK8WPGI+nl2XP+HZ+Aa8W97S0LaICofuHhwd8RsCnuM3Wc9m+FidCre
5zPhOcMVfKuv92tXOm0MpPWiPgBdP/6MVbzm8uv6OrMUIqAShnr4r1MHMEF8KiRVKtbDDIx0he6n
enpKOiSOpxxvcxc5/8Oda8sez5yoi97//w62mHChjTP7Zs4QN42bJ5F6Rsk9iaR7sqFJ22FVSojL
Kv5f1Z7WCNRBL4tt1KZoGPl0wfM3oDu0cb+V654bvx8zzw1W/xOpvQtiBhlfhnGGHTNlyQr/xqhw
SkqdyJlQF6ja86kjoY76/1Y3+e4PkyWWtKeEXwwYRVGfdfXOizt0jX07OuGemrsHFC0/SB87/OiH
YLpSba1Sc+GTdP4e6ZKsRXfiflywo2a4CZ0ZvNGauRUZVnqh/ersCBQ9yPvMvK0Z/PzSwpHA+GRZ
gqyKCA8A6tjNNepVXT8ikykYZmUqjPRx5MnOyk+xFueHtaFC+rcuMLnqgaADN5VgTemZaOWUOqkc
H3nOkvlORn4BgMHRpvvfR7tdCHU6P/8eJHllnBCJvMrhE7BqB9jbdru+Hk4K2Y880lB2rMEHP8iJ
1cuB8Q9H0DEPYx9/MIdgGBiR3P4C0VsFerWgp9jOs5cApjVuZfvujtjafM58zXqZn/d0janiLlua
yDEqupVRqP4Su1lTBuak6D4xx6bxF5e2Yo6BgO5QiAoj4JPNhPL/1zV/iJOgK1nVqRDXac99mX65
/eqkZ88SMnFQc9r+1tUyxvmBc7fprGZF5/2BruxogfcVQEUcDCBrYi5Wj6VgyaGv/1wNvUTHa+aq
vdj4YSCDcK+oCoVumBAeIYUsPkslRnXbstMd/68CcpjEeJE3L2beWkfDxXaCTjgYw5HRCbUL6Q6x
11rP/FPzsF740NXPWQFFkFHl7+fNyQSnUbKB6XzbSIoisfkkdcUxjVjLNvC9/yUwGN6Bkfr5bDgF
BEx/UuvcQY033FHljL+PlJfdtqGojbVN1BWMMT5dALEvr/cHInHN3tjDJok5pNJihIZSBPeQMwZG
/QD5cnQLr/anPajyT+OZkBg6OuaRCtEbUxZ7XNHBUO4fzBvGC0RXrdjf2kIaphG9JnW6U+Y4Evj8
hlrFfn/DSJKrzsnTMKRqwnCYl//M0tjL0PPt+41BD46VjTx3yRwPGhf9MLWEgXMySUgP7D2rkp5W
0igIf8jMnenj+UX7bT8RMpfTIZtrYUr2q3mrnbEV3uk64rXFtb/A6snlaxpLDd6lHPl3B6ybtw+m
qerXTlOKA7wdG5nXRizr9OYIn836agDMhon6+bmkQNPT28L/wRdSu38hVbAdWxjUIIUhNmmRvAu8
ca9zeioHPSLo9jSnVF60HKjXzNS8dqQw5r03wzU7qLH6keGDYUBclkkK+lYMpV6TDFgswuq9rOfp
SzvNYxfOj0xF+aCf0t8A2VAuPSTddSciMy0p9hjzII20lLHoJ0ldbVDe+1I97lp92iEbEAPLvfPA
oSC9igXMZ3kErz/pta9uR8OT7d2HE1mlm+zn5qjjMxaw4Sy+7jIjOtLV08ewF+d19d2bzCOhQbgc
7DyqKCbrNFx71A8IeIAVhUtb4P/xZdh0ar2N/fuuLfp3f53SB0V5I+0MxnJJ8Csic9JoruL/15U2
J6Zeno3ha7giuGE1wKTDu7c4xgAUUAbcLMTU8bphN9TWDM4WKnERkhM8iiOP8fiw87EDnPw/gOoI
Yt+O0fSMVHzp209yUU0PVdJoZyi2/OIWUU+2pKlqTq6DeSgnRYENoESRSyieLx1yDuQhJw7x8kor
F6PWE7JQ7BkJfEhW4S/Npj3DNMdEr3gU9BDa/OA0c0j59oDIQ7Y9mLqMNgBQP51Af1Ew53vT98q/
g8x5p0DG9WRFVRic9QABFUKdcc7Dzac6a4AXBvsD0VmT+uOocZAPUkCb0JdTfB0TNTgb+aJdmdFT
l3as1qYWXFIdg8e3wbOKBU4ogH2XVU0AS44zaFqK9DIDd+OcA/TD+BMYy8UaOBfI5UDD/d3IaUH1
6Rx9R6J0kIflUhHxra8LkL8diYJ8IB/eBw44TTGqd6yDWQ8BCCAU/lzqYzNWp0Bl4CDll2Hl9tH/
C5Ld3u0+QKi5KiLtG98k5ZsOOU2ZVVDJUDqqWF/s+wuIdQQ27Bk8m9Fv7Uf5Q7O6vA+k2IUjK0od
rsligC/5fIO4a13ssaF2mDTVz4pSHuCXdKpGS5+YDEG9x4GXAeFVnVTVeDmcr2fZxLa7Dg7YSUzD
acgYJOo//mL+5PLbJ4XpFruomLWYw8qUVVMVjvTjjTylxWj/ElQiWI3hG6VfBiiA5R4he11sDRrz
5WsnUZ1BTLZab4QhuHQSoS8bIJdOheWVegLzWza4qT47iJMyKaBE/MWvPU+N/q3AKIT2jF+e657W
MqPGV5dOjfJisEtav3dm3xkcC3DgyTqizoPbo4HtfGhrTXBMT5aUW/u2BUA+RXxYZ1YI8rq0anMt
k+Rg9ARwOI6RIf4fw9e5nXmcA8M0OnsL7Zrc12pJlO3kGfL4/dph5WL0ci836/NR5pXzCEalVxjp
Dvq0pPF+XWewIhnNsKE+YYl3wkQld9D066mqf9wBmhKc9937uFwlCGRR7gAC5kXt+QyxUN3qzaBX
KzDagNdBnyY3Vz2j31XZdMiK6ylMJmwhWPsEEMG3SqW49sY5uaiykkLmHx1QyVmDvBOzA82xblVX
tUGIZCvIxzrHd1KjQQr95xI/alcSTjUwtXNpmbs/NIQ8NzlewKRSVhz3Kyg4Ko8qQ1fC1XYFi+6p
4HGghDJklQMVxrhvDfAWCnEOZaud1FfnmmYa4vF8/JkA8Ijz8piQa/3pHlbUwCuVUb3xU9uNAYwc
LCsGwiPJiCSGSnbwnWnpK5YMwj41GrGBHxNRY2HB2whq2T1NCDE7tzZ0TItt7Jr/tJeK8QAFMR7H
4JxTHgGjOnDlYEQoGVxQ65DC7T+sBMfOwRZsr0XzOQO82g9m3LxKjhFwanlt+MelA3/YrSHTQRx/
7Ijhqd6etfhjWBCFYyat/zF2+e2EGep8rwaibNyY8P4BKwJynAgZZBYS6QCHC4Za/diGoeVUBeay
1FXTdivRncZoCYieC7Bn/j6EEwXIx99r5/vijHWDmUD8pUkVT6o35+uPObLadRmbR4XnZ+YJcT+n
lsqK7vqQ1r7GpyERManGfeeh+bfIZbDqWPEnDg+cLRX+LNUoD4jQC4PhYQuS4a3p4hGC0OcsXdhk
E4LDIi4x2r1J2awVP6IOtSKCN+9RK1/QlS0agJMBhdeC0D/pofdBLg3NgnCGYXuV3qHs28w2GY0N
aCznU8ZNSGFonqAu+hC85klotQn/KlJ6A6c/NFg0zuguYajHQKjN6FYsjp7YPfzYZaveFdvrW+BJ
N4yPe92KIHU7tKoRa9gVbnbk0B6d8OD/waPr+FsJ29rwCHpPqFeab19nw/rKjyOQwSH17/MF+h0m
bYXaDsY7/pt0BNS1stzN9axmKKVSXVzExRQHaZo+lTVW/Z75AaMHjIRm7oCNcUEz+PDjsN5BlYk9
5q1ZJ7RSlVxnSyLPlHkDWFY8+VsPmZNgUPrL14aCAcFS27MrwOaOsvAz0uI2h2WB3+YIFxeM5CI4
nSQJCQy4h+7kjDG0RG/4AP4mUC61AetcsJ6Zda7SlbSVuq9MKrNLkec/lUvUdVyzKW5Oun+Guwl2
9E9+VO9l8rWH9YJrhfqE1EbINsG2zBmmk4tAX8dQfHvwFVIt7i30SRk885SNWB8ZjcBX7wH7CTxB
86Ej1MmO+NwK9bLWOyR7+CByzmIpYfFhxaaVRdUbVJHL6fRMOkMSQ+fMOyVkH9/t4sZwnzJ2UpML
GnvQzOo7G9sZiMs25xASPuwIRCTPgNotUdF7iGmyU9wttKyt/fQJ+OEoAs4Iorwo2zvfYnWxhXLl
EK1KoRfBO3T4vY8YUxB1hlF61mDU2dPfeLPMui9cCfJncxJiTsZSNw5KLgxq0SYx7MQJfybD7Y9P
7vrH50h3ucNkXUzjEH9s5V+FBThW335CmL839GxB/WlWBWRTMet3W1dasCdQuj/DcACVEIh0NCQ6
iJX9B79RCXZL5VD6Y47BkXjFA4+ieQqSASgZOfTNc/bMZtF8yQ++9u417uxh3UpUV4L7zboHVPBr
AVBa3twHPpS3V9sIFt1sL236EwvhBwfc/51vlv0W2z70lQDfWac+E2i6GbvmhWkjTWQvENw5ZvS9
WqeT3WZUGGp8H8Igcc9ZpWGbDhDBgTMHbsLl6eGaDVy3M406DoZN3fOC5fcsroPAXESnm6Gyn2i8
0V2bbOOkL0hBGVtD9DZGUCsv4PeXgIbKVcNiQWoWTmwB2ozXZ5FWA9KWT8GZ+d3SPFsunoeMfA3m
6CMVAx+VEVx2m2lucN3DRLrCkHGUPMSJeTTj+sJwors9f5UZLujA05yFh6PCeQ1DNQsjPITHi0+4
eabRl6Hib63qA1TmihtOCriIu4oGsWe7gXKMFnDEzDxej70AKfa0hVifKEjWoGNePU2PQxMKnURr
g5AD070agpKoBNUHP50aTJPB47/05CBUX79DzosaPPUbA7qhhw+wsy5IJFO67idESoBUVrZwx5jZ
VjbRDMKR15lpY6EP/Auv+2Gfm9MPJnjDF+VohnRdRgBWJZc/yaagNtb6pIx2PlLk+oFx2GP4pfJW
qRDR7C63yg/FV9Lf71jklY31DCQIQVqscLs45Urdh9Bly6sN2ezZ87r0hQ/iUhU55c+NYBsQm7Sf
oMDQndvIgNPMNqw+2ceav2dY/1spjq2QnCwXPujdOMnkqEPt62HbGukmBuHLnmngCFNsDwtrxomE
icGqj2A69OgkQnZ2KHtDu+WMOxbhYwV2v4EqhfgytJFHK6/CuVhUKle0WuZmt/8rsxYjEmtazZpU
I34sfW2AmjOfqy4pSq5eqHaIhToJkJltm01pNkex07QGzs9h12iEZu2OcK/qRZ9/vuZEiVJ4eP4R
HSl735j2WgewlANEHxLtl59tWWwEKKzYmzvlbi7ST1qUwvTGYFK44bdSkaNGsA0vO+5nXsXxFO+S
nu43SnRcUhzXP1hQSv8UTp+9jr63Oj/D6j5hLYQvqTG/6Ar7YTeMJgIAvz/1auQA0OB7nRCUTsZ3
00GS9PhCX8ilGlbLqtG13efKv7PiGyf1xbAFJfyy4EqIseCrA0X++/+nasY6uZIuw8diWn+YC+tZ
PlMlcapwD+LDtRqDapuUpUf4ey//stGWj+KW17Q1m6BCtZhs74fA+arBZXnPQz9sgfQWBw7seEIw
LfTxeFRGJgqyRSxghqdYqksEny7M7K1ngc0NRd1y5ill09MmADHSb4IYOgzx7rdzpA70y/0RHNfa
SR2e3Iah0fnGeOwgSzglcgWuuUTN/yykGSYAjRSjY6Gha8hjzG8OimcTf0sxKjhPtt0cvrP9iJZk
yTQI2VEckBJMA5wcE8nV+ZtescBmKEmniEsea9bRP2lh6hqC4hMWWoq/rqH/KrH/incTmjfYghZT
Gqds9s6Vq0gNfrCMgnjq/VTGFEpoowasbKHyVq+WcS1nrULWHO3cqyIMe2xVvK4r903/ImuSgA2s
JfJ5TkbnzXC4kCNEWAiMRQRvJWe3BgLuApEYuwTJpVYOndUDILL1ffUcOstW0zL0I64hMD8ArAC3
P6GjQn7ZLH87UBCzDcGSoczEEkicdD6J51hkFVhkPnWRSyL2u810UgB4kazIEeCDV4WJwLL3bKlo
W8X3Op8hhHo2fO0lFw/QKt1iafpENbUVXCfCwSBwl9Pjyq4rsfh8vnH9IyuPGujJ0YlmFJVNcpWb
7GYIZejk39naQlVWCfrjKO7NeVRwfrAadXe69jps7fk47aqSuwCU4/B7EWTJsghHeVBzBtL+U2cC
WutWaDFozqyKYT4sTD0P6RGE2FDMV2GtTOXRg0jKvMYnfwpcT+5ZINoWdOK0uO+RLPnPctv7B86n
EXtHlpBzsxOYoi+pic6MPmC+Ig131y8DQTn7xy9js8GyeCgN9egUUuIf4QWGukmwETk9Z5pe3x9Z
0/kRbYluGo68rmF9K/XTZkvWA/eQuiYSyqpn3O8IeLOdX6wSaNaf2+4d2LA7FqrWiwu30bsy8uxZ
C035rwrK3sx/ajP2oXW/BcMmWstrH0SGNC3NGXYarnHQmyW6vaUee5t6+X2Kbgmijp2FylQisLSG
vKbCa2p+m90SeCQkmrXqGirxs1im4wqkqS7z3VDTBPL86vz89959u5qL/Er1C6hJQCMwcjLylCbE
qDVkho9TWlgF+37FLK/SFtxpUlwhudrv3X7aqK53uZP8RWrShxW2v9B8877ycHmcw5aO03cj2QEZ
8gvNSKXwdOEGWVKdM/zzPeYb3+BtTJTji8XYnZ0hO9xAcI3Nn5inZk/2E1CDiS+BweKsvybBfc3z
16F1VYUcKskFtusjS/tBjGUWDBgQLxfCrHap3FT09nmrXCjkUH61MnRHUYcNFHRHq8WGVgjNI552
a4muMZWQqadPNJ8Gub6zLjlANyFyJI5pMlJHbNHPPO5NeUkvKWtEjUvs73hvs1j6vZno7tRx7JtV
Il6tdQEvs8AH159w3i8FFeUHeDwpD02OX/ROOHNx1uW3FcWwaOJx/vC1zEo/TvOIQT7I/Du/3fRc
w8xLGUG8ZQSvOtr3IPMqFe4KQtf1BY1UyJgSyHq2yyHARqAB435K6/v8QVPCU3Qzn6i+0Of1byTV
t1Klni5VvA9HoA/UGwXeQ+hkMeM3QLXhb5rVbWHWNyN86cZ2a//BlWWTGcZT8NcthwmGucXWZNJQ
q0e+XrbynKtEqUfKL6WbOSJEJU3K7p3JcEs8v9aiLCr/qTpFF7iziuPyVlt0xUEpslg3KHjvRf/Y
GKhdNPmIzf+mfwiiS9Z+4Iofij47Y/hGQyw8XObiv/7RQUvNJedMoFEvwhzpNKKqfe02ySL5jz85
OH+LOlM/yOAlZ//fI0nLeNilAw/H9+KWpsXDyM6teIipb3itTQzJWe2Xzr7PyuSNfQaDoirtdliw
1dbXmmgEqqIfBDnyfK4PFoXrUuURGVfBwrsg8SMP7PQJqA9UL9PhN4eGU0CABm0jLO9wNwHoJG2b
9af5lF1B+EOZlH8S0BZNMOF5jqzXB9R/Kpy9qN4KfsVAz2Q8pN66E+G9sfmrjdqgEDahfU1d1v6o
wko8vO/htA2iDyUuN4gnI26V638PATf030rWcbOvhwiGcgtLbF4fAXTSjmzbm3/309iWAGIkssm3
6bC9b8My8ZgG/p9vaRA0kaPsIgNRS6eq7VbaVnVPa0HJoG/5XLbnbZe3QlhGsmZyg9ZGihisg/1P
ipSQ+tX01YCVuzU61USFlT34tgHLf3D7DXrNGiF16U+cfbzq2v2zO44EgUVxdb/Hq2i4STCgpVfP
InGicyAXgLxcI66zQsIGX5xuDmfhIxHCx0Jy4fsvb+H3AJW/hZTBKNj+E8CYsIz+s5QjGXbbSToM
dBDGNwQefmToSZbqQA8Z6swDAgtPpfDrVJA951NmZvQ0KryD0biX/O5EG25/t6oRjfFmjAmgbQsz
mHp0f+cqSqFSmKKeUH/6eUkq40/PrYByGRWH6TspexiqIC1rsTxfdQLwGbKwcjI4b8Zb2AER45rf
UPz4/CoUGDLdozZd5DDLQm7oxMCIHISzLfFH/rjhuS5t9B9rLh6rrJTpegxXwZUdI2t9/eaHW600
ejLj7XCOFxFj1JqgkFj32W92eWB1EnSWTBuviweCjRDjUTGuvWECx/CWUS1C2cZiZz0JNuhsihk6
lMwMqU5uRmNHNs6F6TD3b7FLBPXWjt16BM09AeFH5+k5xWz1ZD0jHNg0ghXe7qNa1MnCsf9UflNt
GrBoTB5X+87NgGO4enRtfrlVl3MQetN7CHc8XcOsx+ubHY4RiakbXwQItdfqF9N5Z1Z01MGZsglZ
yY7bt11mYCxLrUcmC+99OpqB6T1m41wdTfbiF1o7FOSqp/yPUU86YRQjZIpjp//bjFKY7DXr4JBp
DtCEvQkDn233PLZWnZfnZUXp7I1KQFgYbXVdBed8ELmduEYUpdxkauZExteml2W8w5F+/Dub9q31
RSovH2jlUAFcmYx8uKccmk8ahrJNEjHNwcxmAI/+XV3VH2B+H+cp04g2V1SS+eGL8jgI5Ue8Fezd
jQ91ZYOSgfK2j0lVrJQ0jq/x5LiINSWRcL/7MGwa4UjR/y7QFC3jVupvDYVa7C/1LSJof7mFAH27
K0tDC11pbjRPzQoCAGXa/I0VZwlh1V50+AP98Ivny1pquLG6gWVWEUKEoKMgDSCToswc+d22fsz3
y/eykE0qPrZ9EHmLUas1ETqm6JW5WU/3WFVwHYeFUAoy0fNh9tld+numt3YRoYxTjHI0/KkBMq2v
xcn5di0IQiuvIE9mwTy9JJIJwtsXwIAqIMyNteDxds9Yz20qzUgV8NxvRzwDv8NeaBM0JqHLDYpD
CdowV4lUAwjPuZzw6p5jtPYWYieukSO0DB7zbmY1H3d9Qk3H6AZSAPIfEyziNp7gyISA2iE6S6UN
jvz/w7goA+YYEj5kyRQwzB9c7ZAJLpXKwJAk4OAacc1B1Mgc1bJe+tJvLQCRxzlR5nbaSOOxLepZ
34VRVS7sOO4Z9LPVV4BXd1GY1SVgQbNArXCoI1qxC7/QgS1bNnN/1nMID8WWY6LNPkS9RzKqE8o/
ItPFhmOJwRuQ1RQEloedb/XSYtTS24t3YlsGVBN/cxpxfeT7WiwbOuxJ8joMOuEIvjRPKPoaALCF
B0MqHQDO0lw6H3K4XoEHEjwbH60oPW5EWgoVu/EcVUxslgGiTqQ1FSDCqdFxNguDvQoLV34npWME
JIKsXGO5s23226Etaj39aUS2xKhC+K5T2paDV8scOY7VWChCsNcf2qtgxThsefVhZz4MkYDXeFP5
1d+d6DBLZKivB2ii2qBLnWOixu3fC8+hRVhQ+wrMUYq8JkCI737M4c4Q2rEfWHmDE0SrjxlGgc5I
n+2Y+wW2R+/eHtQxRO3ekyBuoC058x03XegXwb2B30vkVbSRaU7Avxms34qHcaKlbLE0NWhO6qwt
0l86h6diyRXtT8ugi9zLm6aCxA6WKNV9badNdxEWLwMY2nnlRd0Z7C6UOro0x+HO5n2+iLe7HppT
FB3FY/X/XBk7zlLco1h7eduM+HwHacfJ3NHL5gpxWsQydcUUGLb+gx4hS0+oydnL24f5m3geQ17e
qQJQxQzAMXGhv/uax+0k091fRLKhZWUtg2ZDHS3KfeQrHlkESzF9gtatILKObORg8OHiN3pMCxzM
Q/EHAxzkh/fskHjR8ah2u2zK0SEK10xchiT7P9vG4DZ9zxUS88eQMCeugV3QNq5IHlpCl8BsOC3H
wdEYmJTlLhtOKnRDqHvlQ4+XnD9JbRd8lwMVzDG7qG9xkln9MMY6tDuCWls6MtnqC2wMorrQsaUj
vIqv0c+2UqttWKr4DiKjNfjg4aJv+MA8EHoHuB4RnmWSfCjBGDSTCSL+Z5JOXgFYO4ad7vqAGFZK
ZVQQGrszzXt8Y+FZl9z5hoKm1gZZ8ri2cHYdbZRtFgndFBkYxdCX/FF+RQ2VQ1fReQoCy6kssHuz
NLTzPBF78PAT8RuwaVugNgMUkEjQa8ZwjbT2TcrHrkl2O8l6ucBo5SSqrBNYL03ksGcre09cvUSq
yl656el5PAWuqxhj2iBOzA9EbjcJ7WMdXs/b5XEO6UILK+2+eJkON0Mbx0cajf14EpSrVcWIBGiZ
7XQWdV/q3JGKH1XNuC2ojQ0kp5bnX6yee5brP4daMbsVvIBZiI68i8e8Nw/KlSwFw9mY4GbNZCnU
jCACFfhFrG7q741H0GH+IizxAyZ7SpXEnlEhktPq2IqggQ0lUgkr95yDCshMf01Thex6+81tueKA
lbzevg4E9UH+T767gWkVKx/c9Ct1RBU6lWMumLGUEWKFd5bGV8p2Xk5MxlSvPMr8BLMuIw7nBn7f
hglC5V6HxkRxU7KK4Ep29uH6HYMIVGv0PZRYNYHNzMfqxClkULeHSlwzX8wF2Clwn6Ean2UmKNVS
ld/tLWdRRHQI5DRL71pr4/60rDJ9C33rKEx3NEl3Nj5MjXxq1wUdyNtUSxl0Wf+l6YyvAuAnJ/gL
94NIB1z03UX77QxOU+XgLw65m8IPNMflqa/GJApm72mBN0d7qOME3BVT3Z1aGE5q1R6fdEzoiEPc
6LmGoKhC91z4V1rK86ldLkj/xIrm59hPPoCsMR1YqKtPeKL6fYDHHR0eiKdbb9YAuO10OgOiO1Zn
APM/N7ufRzc2ynX2jHmV0WaWvetPAzHnT5fKM5QpY4JkDrO7S5i8wrZw0BzCgW3mJenakKh2g4rU
A+UoBVVR9QMah09btaQ34IjWHndDnM6Bqw0SK/+wMhl74Um9xyD+CDVvwifN3FSSfbek6VQ/CUA4
FDo6z6/mmW14zm+WuIx9aqF3dG+zDu3trirkJ0xMr+/CYQX9pfyv01Q2ifRzIUVXyMidr0QJRMZ8
g7TeqxNHMAm4tNuPHq20iK5KEfv1eMwZ2wBUxIM7tFCCwIGfxWyU04bV+r8JVRXjYip7mnijulFV
F/5MwBxHEBSSu4AJCveF2eXDuK08DnOoda9DTBKWzAJztXcLeyEZLb6REfeAfmn8M2mYxCaXdHNE
c5cGv8yJDoTRGZx7xvwq/NdhGfRoP+I7kt5fe2eZgCZ1wtrU8kI99RDHGCd6TmIXQGbx+/yL0wvN
yZmQU5L6Wsv8dE3JaxGqyRcgwERdv63GzGCiMpkqJyiB1GZ8Dtdn20NvCdoDkzCBkJdKS+tSV6KQ
UYtokcWd5r7ctK2ooXwHoGaAvc10mB/yTc6a8pYEfJTI38f9pqnhtjneYTSifE6F0sc3i3V2jVNj
6pyjrHuPRJ3t6jlFhNTckN4VlL6u6OI+tC/p7yreblCF1sGxLn6NElpCkY6ea5cJ+xB6hviRHgAa
4xZnlABC8zfT5BIBX11Y4cMbXwS027GJjgTdsjZxLd3E97K6tYLXV9CQgtWkm6xdvkZVn8o6m+6i
bY9dE2JgkhNc8NWpo9beVPya/gJgOWpcu5iyPfUWTXXr/0NDrD9WCCOKwxeUuIW6p6ut9FLBE99B
B6cW53A9FlX5ohSpI3ikB7M4h6MBm/4UdntN8On3pY5IyKL+3Pm3ScaknMEp6PTDKgikYD6LmuEG
M8rS8AMQ7QTlHYL2Ogbp3QuFv9E2SdAQ6TC9xoPs2NINy5L1ffITT+wYFeA7n4u0MKkKpPAvlfbO
ITqF+Nwa0Ps4jxV/eZ8INEZSUMZzx/Zwrk22WgeLy+AsT4hveFj3S6sICcIExHqI7cqpzWZtgJgX
4atquKS+vGwYh2Q1MDfTPPqqzwbqluYl4/z/mQrKuyDstslQqFDD9uyIasoJFZ9J+Q4xRxTa6RBQ
jrW3BLMBe//E5SanZnb0D5MSYS56WLq1ZFh/ppacHJ0ssBxnDyHIDiZno41BZoi0vuukkwqX8wAE
R/YbGAaM6geJchpsEvWi3YwLQiWhxh+nMl0j0YvLHUp3+fFLwl8qRgPJ050e1w84ssNuQOFDnGPM
myAb8vNSXfXuXIlLWxivCC7OEiBalWxwXDVBh3RZczCmkIFPSxYISt/K+okjBwB7OlhjqVPtU3Cu
G1vvGbbhuvLtUgEtk0f3GhbouoAySi+n3Q6uKfYSOWvEBrkf39o4fJxv5HyIO04/1iutOWFjMrsT
B2LbFr2ovJSURj+T6ZmhC1OmDNveIisYYJ+qwTl5eCuNHTQJNCoFvcdJgyEUEcvpxTKK58gZz6ni
FcgPz1tTLj4H782iaj3vQzNyBzTT2a9xKxnTrhQufEJkPieQ/0zSKkHcVqscdGjEgcNqD1djVKuY
xy6UjRWGn242JILhnzkxY/PwU8uAgPv9xTnjWhEBk/DJdX5aEzmdgEc7ZV7Ikt2OMSL6IzjGtVhV
jxkbPohst2PK2plCEcUZn8jURh1aOg4kqd75j1bwQ2VYgUIjsqlDGXf6psTQ8S7pk4O6D74qiVwv
XTjOUTyMy21/JAYmXfCtlYIl7rbcT+gQqzmY4RrukiQUY/ZKqZkVvbM8FCkls4Tw0+6tGJZP6O3p
xJ6KYVIkNCXWhuFx4z+71I6jowpken8IWybUxSr7wbOePMB9E+lyf7+2oPTWKeMbv17ql+A1doMl
hq1VgeWLWYlVZ4k+R2BQjKRLXIwfaqsZQsA0HYC6L4/+7dfbaK+dnCAOXq+edli8xJO2Cu1PDYaV
TCAsH6g++P+M1x3OzOtZRJ26hFKhoRGGPlPxyk867W25Ec7xAlpxdn9wA2DWo4Lp7EQx4hj5nGDq
bFHmUIGF7ZQMPAaIHjbnQGSlVUgRd8qVLvt3u4K/oeS3dADbRtPP5D7EZhre5q840cx7EMsFagc7
TETCqhPdcJ8+wqpUP8Hs+r+MPla6952blL77qlG5DkkMXC2UH0Wk8XeGM/TAIvugQTZGeLgCGn+x
zsQJBtcyv9G/U7Bo4LRHUOVBp2OvqkJ5DKdQM3KLUyxuTYKbqEuIjRU1UubprApLGx3Nnbza4vYx
VGQJMXLiiBxv9BRnuRv/fK593Is7kEH8rAzMr2lqMkt0x4kbQfRAc48kkEPrSkepX6y1i4tol3uV
PASmSah+hrvepdi6DXzQfr3dd7fXPZNIv3Ntw8TW4iCiYPBNVM3K+bG6QpH4JWg7DbQzC/cPMEcw
Iq5dVOt/lbqrAVejvg2CvKVBx+TnsHitQcZCN9ubvSBEFcGs/PXv2MjOm9pNd4RrZR5SEv/ccH5Z
ku4aeBHphJZLhG58ylnt6RIwEwgTv+i55bG2QZ0D8+JD6wiZT+rD4+/KSacWDAQKNZNZ3OkgGEKm
xO6n+fXQ4QOpL8fCgn8f9ABBSRXSyOQAusi5umq7tS3tI3KyIHmfZvgZn2q74JchgH1cK4fhku2Z
/lKXeCgGeHWGC7CFj/lPUlrLTWkMsrps5aJCxtyxTkQbN6WkAJvxi4GqEsoj394l9YIm1nPboCTR
d0kUuuHBUDlR/ZLYssuV2mzImHWgIrJtMNbCHrLIFQdn6p8bFXhFx5deoVeuCE5yZxQ7DqDXeVpv
dKKUs9H6h1cgh0La+nHQEgtG5VILGwfikqyEU6EQ0OS3lMyJwTj5dDmWrIL/5Ghijg31Jtt9k7/S
m1kLZ8R2cQ7uiEjf0a5oy/QUKQsEeIl8fMdyPNu7cseD4n3GFjQl2jqsv0nS7062uDo8vMf9FRjA
LiLOvTFmBH1tXr66fUAlKK3U15/a2U8e24MZ0UpRHGME8UakDWNYhD0VRvxC89TlV6Iz7qKjbt7G
KP1z6r344MpejVQGWQeH99bmCklWOi++gix3p6CURermqQn7yfHIpr9lbL0+GfWsQ/1r9uZVPz6d
3Ep0I+ryM1B86N2hmd3dTnLFK0+H96RVX0QAL7YzTx+PG5yeGGYfgBjzFY7hXszPPOrW7LJO+RcU
gBBV5t/L1wFd0oDuSa9hCcMExQopNGU+pkFjTKT0RZSrYvZEegz2GD7Pf3+zHVKt2dZnM158+lZk
rczTyJKTmp78BGvsB+WvnUfZesjFouo2OTLmf/oa7MH2SOSI0/GoM1+6N+NkoFQyu9QkLaLS+/gx
YbM/S4sYYfWCxbAWvvoYfYHnr64USw4gV7smRbhVFIXYAEELO9TL4DeHwW2kPLuuOuq/MEZBoXGs
4gsUSljSsbbuM7yqKp7L94U2zrya35yeTfgzrLPUsJuaQ5e13/A95lFD8hVIgJX/cKDreDGhyT70
bRMf4wpiyGF7fG7RMSxcm+uXmNcPR1vxx3OVk5G5lmjiXW0iFqBzph0MQgNKfjjsMg3MWy82UWG7
QOM4HLi3ZxlJovaPZIJm+uLHxnoNHXn4WZuxPYuDuCb21yJDDrWeg+m/b/nZ7Ydwu1TSx168JkfT
99Q6nPwuZrWNmouG3vUAKKmLLRYhyUInarzHQxgRdrvRlPGQyeGMi8XznidGUtSsV9gghBhT1DQR
6N1fsUcVXQaqkT++bsbNIIo8M6wHGMdAEs767pA3NscFKTgo5+l6K4J9ESnDcgB2AHOtUHCiGX2E
2UP/vXTIhf53tr6xrdbw7rX/evtd0zqApdB915h8EOSR7rBv603xOyVmG0XBjdjujwAkiNGE0QZr
liMEjhr4GAAAN7hyxEAURJ3RjyRddvYmPFAo3GM10nwINgy8VSPuAKRovV4kKY2ubD4mK9WpKNTz
E4Ps2FM3b1OkVypuYC8hBlvxHoXltTXWWUJXo1bDzsdwcD9+CMUpUst14Toayw7CmPm9ED0saWMG
XpBzhYTF+TNT9jbjwCBWJSHwACO9fv+Jr0UTg9BANNLLw9e+1nyLKIl4foJw7SZZ8wP+JfauTYJD
XK6dRA5q5Pi4lwl8FpI1l4xgQBBo9KoI3IXk7cx+OoFZ7ubz/sJo2ErP8H0TV8bhSvw0DS/gzAl1
zvcURypLRSLkOXusXpet0kIwjtzveJApJeKrnzwOIEClK8n7BsoYs8j8OKUt6PtdzTkQ1i+Amq1C
B6hm6EmTLPS2WDXyFOlBfd+qYLhuDQWVUG/qTAWIvtRsr3TJaqZlrPADT1EeSU0qX8GmFTpXcwb5
dvePZFyKxbE1X5Tu1bbUiWnK0bba9HLU32TfBWiAw7CjL+pnHV/2DDZLJiBronsBQZpNyzCWxaDm
LaseGMNWKMmjmaBS8opW/QcloEEe1XcMT5CcRgui5Ab8j8+eLSFNqM5uzsKm4BBy+8V926FpoYB8
QgUMlMu+6R9EeO+BHiBNTBOCRhnj/o9pFk+ArFxF/yCdCvwrpQ9Lqf+41rQl+UV4vYtAMNQIcBtv
02Lgz2OAW5gHS/SFUNQhgfUnj6n/Pr9z1vFzfIimpfFH1nzc96z0gnaJ4hiQ9lpFwO9nfW8Ujou9
+673F7GlFiOZ7XgVhU1KQjfvdvmsHPQpacyvAdF2gHF5qI6pgwhFx3Ce+Cq82LQDCosrPzWbRc+6
egnAj/w8yKaOrVMTWV+i2Eo3k0A3N3areW3v4zU/bQ1ITFk3r22AeN2EAAPnlWjRizichSDHVfID
iH7P5Tma7aMTORjy19foLR0Kzk8Ou6xx6zKGfEs05xrP13iRJrVj/9eLMnNjtsn0rXEiFURzTqOy
zeDbcHg3q7iqbE3Hdra6PUckhfFMlowdD5SohpXlQEck3b4vducS4MQZJ5S5JZ4elTQLCaBB8m/p
UGXaY+TSnHc/Wh5qJoKAZMG9xUXDvyRC1Hvv2p35efxgO9pFC3Z1nKWQ8dnmU2PYVfJbXeKP9GjX
QkCqwsntyk7lG4rTZUONb7lO1Dg1VLKerxNacbuVABsjN26CowuL3+07VkFvUGrJtrxzIQATr0Xw
fa0CQ/TjYUvqDsMZE7RHkztRTYLvB59b5YZZtiq9k6q4PI4q1+VC9bdfj1mmy7zhhGzXwVoIla2D
gYaNmRc2PxD93l89QCYKLOr4u08H1crXEvPEoSSTP5u3XDBfQwyPkjdzHoC04FEOo/8+CrPMJQg6
4TMwXj5gSVOKd4Lr7shRpX6tKCkTVfZFwOTY7zxWNMAaXQPKoEV3gOQWCJfgwnELI+8SMT5XemUg
OBD8yOZizwoOFg0xqc2HuBMcxk2RvKNS/TJZU2yVPvvzUvw1sIVLTRGS7RmW9T3zl2lmsijiqE7S
zqSAXGpxTxHkXeHTPNgmP1fUPHJuGXGuFFYZSzNz0KMGX/kE16KpTAG9X7G5f+34QR4OIW+SIqyX
fyK3BS3cfj0CRALjzhx/KbWgu4a9Wken9Ad1j9AT6KaGMogIiLz8TWh/6IMGCg4bE15HyMTZ73zA
nS4bW8fUzWuqvuAyOCGAfTbPY+fw63dwBMGqsTsyZcYKdyXPPmZHjHncqwq7zgxkexO/h/9R+ye2
CeknYW6woPqAuIrgxeAmRFjjKNQDeDG6+0jsU6E4EBp2mTM1gP9haKJe9sMxLg4Quz4QpRKGWIK7
LjVG9AS9vvxZ6AYv3oxKo+fNhTgwhAS64Ru7nQRBAEvR9KbVV/QTGctDwKHPy9Iyo9sSyzpX6opC
SncgDEX5rTlwot8K0TfYZ7V+1j9lM/iyxSw9BiAS7NLtlvGH95tQtqjp1fISXpG7HEpEOuSaj9Bd
f3Ux0N0h6dh4OU6vWpUrHJ+6tA0rWqqtvXWPNWshZIMnvKrrqSCJhHRXQcCP2Lfl9zImr514WBwm
/rtx9nW66OH5jx1qdNKtlXv6XhDM3NHxlH4H6UwT3PZzcMGRXWIdJdHsW8T75MUM9gr9fDmNJ36g
zNHpz7DBlp4RSSV1qABuCXuPCnIAObfvZbhgJ1xPZ83FqAjx42cgCT6as2kBzFYiL9yrLhrsvv7z
yWpnYirLrfu8CYh/Sk2DDLDql+FmADGoBm2ORAcCE+8FkSi4cngnQdl1IOBE506GuCzksxZkGPoU
ebg76k6DXLj67ZkXOoHjr+VsWIPzQMEMxKzG3lmCbM84QFc6hWG6gb7ACM06c1w4QtvWb4tRXY3K
mLOrYceWt3gnG9ymVwCv+bBMQ/p1bqXv1A4ufP0yTTAD+pMo35dpZmY56oS350mW+W+l27/DQ+rd
tvm3PaFIyh8GEHb8yNN07HsZrkTX8lIH/tV0ksH8wuIGhg+XC3yWd4W9F8dw8BpMQtAOMY8ACBSk
D24tdFEfh2auTFu1zryWQQ5/0exkvaeyz9UWYzaIJK1m4ToTgv2ea30zLol1xvrGvPs0H6p76EU2
oK35UdQ8kKcaJsm6kbaHiRdhVDPGZ/6wjLt54epy+daOc61cPZcTLq+tRXrbCnKxnroSfcuD26Dd
vZ+Rt/5v9l2SFNi5EerUzDqzUC9yQ/2WOktMBm+CANr0T0McjKbGzRiL7kJTjUsC1k8x9LHMTpbF
IETrbmggZituSkkYGsAqsFnE4K3OgrbMR4ncBGRgR0zqRjt/D01yJr+iQuAknmQ44MTXf41kTupf
7nP17IaU27q9mKvuDIsKyLy2pcP4HbTLwzxMxz8tyLLlr+3BExBNorGaWYqtIDHR0L387jDGgIkc
/WsvTbIPRVJctk+NogIgJFph/2JyHeRi3kDchTISm29K3jKMHEKrAvGPO/9IbKc5bfti4nc5MdoJ
GYNSEqHLyqb0yWsTgrCeYbRwsVOnCm7PfepggrXYg6aRkPl06Hv9vPH1OoI1vZ3Z5Bag/lxa6y4V
Hz+jCqAQJsKTq/2u3EdBQ5D5FbnnTi+BYgS0j2PdpOzdGkn8teXhz8iknLh7P/YTD6b7SjIFYf5t
m4awqE0qqe5axo4NhT3ePpvJF3wtX62SOcUBRAbCUlEPBaJ535fY+R/w8snJrK8c4KdaoFiakv1S
gIcFwTKTB20W3ZplCFTVDlZuvvm73Gg1PPlyWt0JzBlWwDJoDwoqS3QWgk59VdHRXtYZPQf9/4zZ
Tlb64XORIji8YXJ/FH+qTpj3mPPHh1/WyniJm6zi9igHvAprMTl2TQhQbzW+re1ZRkK40m7W7oFr
aB3Nd6igZ51uR0PjLONjQ1/gHekNmfMTLj9VDVmvsmy80Mjzg2oq2RUx924HSYrfVBDeA5QW7NHq
HG0Y7kP6OBal7O0NWwUq8T4pTJ+zP/dVvN039Td7Jl3NdbXxqUAqHqGrffH4TCVIlltJ4LjFR8XD
FjGeVEU0JKS5UOdsIxuan/NJixzswWQwkIeL2l0zZFWkLCn0tAsDahRwu7gR0QqxnCx3VwZWXGft
I2dFcWClo8AHB2fvGxhCb7U2Fm3SeLUvZ2gfpl/ZjAyNjD29CxGNyr3h9O9fVoRNYVA59KmExgfB
3Y+juZE6y21FUxKLpD3lrPLnB1Fl5cNo9aYu0FHXkO8KXegkdI3ajG7PvXnHc/L+N4Mjhf3pCIfD
MYbI9CKpNB2TmbFlIID3VpckZEe4fKsW4mHy1tULbC4NbdXtWqF2XvyRRdubMGVCflcCjJKhHNdj
8JSAVGxE8kbK9D7WwJHg7yLUg8SmOdAAs5HX5FsM2oUycdEzBC39zNq+dgxEb+61Y/c7NHpnmrrs
mw+kgf1rosZ+GqxK5HLI9IJbqzVsw9lTERhoUGqSTZOe3jaUACbduNNare30uJsvbkYJCQtytNKv
8+hDhOA4YE6ZQeTWRrJkVuaLXu5cqF9mGV9Cjtzt9GV2xOTwldWZyMFBpGiNMVPgVEzNfJqQJBh0
zedDdKJSPWGdq2mZZjSlqOfjEYpwy0MuActlc+Obv1Y93FhSCwWNDLnQzow/7iY6O/u9ITGLGcWp
loQPz8mj/MILEun5GGh7TCxCwyaiVvmW5nUqaYxj0WkilP2H7vdjIGuusi7B3YXGiWSUNsU1d+Vj
srjBkJhEB9gVn/mDujY5a6ZOMZJqeTsUphAIOr1xMTJ0v/Vih+FwAyC4Rs9Vg++7ZKAZAwOUqY6r
8vqhK3fDfgN5KJ2UHEt61/t7R3QO5RVNq6I5ewuxzmqvFplOXkrpBflDLudetPdtys9nLcrUnR7d
wCEDYbGQfAAVXjAw27rh2qF2FAyQAoQjotIPQT1jP9lpR/eXZdEEEXrRoYdoTNWOzEVU75+EMa0o
BUEZ2S3sPOSME2F1IltbvJh5n/g3GQDEjnqKHPe86vn7Lx2u8V2lyez7Cv4VBYCeV3VRQnTSz3y2
6mVqOsYZrccAiRxIu0J1/eEbtMkPN+4OHOJfW+sKvKssh+XUb5Jj43pmpy80sNAiG8agHsLtDjQy
HWEXmWdBiNIV7v8evTI+LlEo/TAqKrA/Eh1M7Kh6OeTwQTyy0qXXtxadLIEASOcoH6yVZZydVbwM
0PXj6QeWmXE3vjMHjS3oWLxL3N3lnyWNFnoy1qnpPdiJXLGuQdseH+gIeGJhf5p/lcvT/IVcNAIv
PSyty1jMsyj8+8TCJ0BmtFiVz/LSZB2R/Si51RyYvFiY/EYfuI3N7OWofY8AEoh+ugSq6bHKePAL
u+pMzzL1sOHEwCiGDViQ/dr5EhOu8jKGZfaqiQJxK642rhG+f2X+jKaVDXJ318Ehz2qyibaQ8QKv
jkHN8aOydwPO7tPhk0Sr5iZ709Z9i+qS5u8Gin69ysjqJElAY/A3egM/KVSPjWHhgmdCjRvh8Tnj
c2BUNA5zbWlN3hr0IyfHaVhDl0wAtdt31RFNONKaBkDtr/JVips0UkuB/vB0jkmW6NpuoJxsj/mq
tQyqexectTTHxYb3U5n3STn95mwshRY8b3V4ZV7um8DBNUwxnnoqjEgND4tGJlpx5zX0y6tzqQyn
qQbd4iLcDXNcpG30RmJcRf0uRIEKRkaQ5caK4cQa+grCgs8gUiUZh13l+0r6wtgjIFXRGBZG/YDa
GkQJ336CoScUbrUbw2iyRricR34gc+M8xy1c0JQZW8d41U7Ul28P25nFIWX6BzwV+2Y0dMO0PpJr
ldVQ4pTpUaZ1Z2/bwSe8Pu5xY+kC1jk5HPu4/UGFEvU2sfW1cYJaIrsvmFTYLcuUq8Y6bohz/NAG
AHGFnEEebvPs4syqKbX76oPLgnFj2qhRHUzvr9aZd206uQQOuMiLsIB78gdEfgm54bAQ+1NwF6ca
0D/XbAI712kiZUY61B3uYKybWpsIPiZ43ZYz/RkM4BZ2AIioa+w58KggGfluYCPUWB2FW5u9ebX0
+HMPwzBMHRl4I5GU4yG4IRmLuL1vY4nb5NMoJHUK1HcstRudjVJZCYcWOzOCAmEoIRUdu1s2lKOq
Tx5MuDfbbZjQyhTFCRozRRNfalxtqe2StMlw4gnkAmJs5jp2NN12c9SAa5lw2wPN0jZD0Ki6Y3lZ
zY5z6hMGkQRYT7Thav00HVnvsyL/DH7UQKb8Q04bcojHq2Sk4mmTJ5AKOA3IVoMAwXcMe6ebtTZf
B26Orr6RqLWtOy1ko4YDs/SLWaWBERPYZ6+07Vx4/keARIgxwqpN38NjpP1zvzSlBWzfV5JH4Nt8
M4pT/RKYdNBbyX72OBvYOrfK600yryRn31mNB0C5UwoGfQHsK3RnZ3cIXJK5Ppaqo93JqQZQQxAN
lP4+EqogsllGc4LcD8e4LKMn8Qxqxn2FiP1kvOAmz6i3Lax+rVFco9SpYaq5M7pEgtGr+gDHyaaL
UB784gXviw/pfv15vL6OVjTkF4QzHcIL5AfjiVOsdzxx5c0/9Stm3UkP9MyU1TdfqxwfpEgwiwxF
HM5P/SQ9kx6t/a2HrPEvMD0Dt3WzG3+yhukF4fBJAdMmRrjnOiLwW/4iEM9e10dZzBb04PE9a6ya
AfTmD9Be6lpu2Qhlt7J+ZnOPU1lR61NkWEvOFOxoRCXZKbtiAYkh4F6nMKbxxGMyjHTm3PEorpmb
bdahmOMzzfLRknkaX+w8f146jYy60QoJ7aUdJmK7GlYbvw4dGhfv2lgdPYu307aa596rWNr+AAro
xS7AFGSuPTAbsvlDQ9iOYNb2aJRBFar7/KjV7RRBJDsRjQFZ0KaUTbVIu71VplEuZfidNqIMevgC
TRcG6jZZ6+laiGuJ/9YTm67K+JOb2SgqT8eSbd59aMsPrlO4VOSR4PEKLbb9o8AXehj2Ztruq/sA
kuuZvqq4KRrp/YBFSEFx79o/JBo/qJCgWEI/TdaKYyw6Up5rEl4rl/egVY4MadOah2UgpfBwI16c
4g/y6tV0NJYfg22GD8JPrkNmgb1F9Nxgi4bfbYrqZj85kR3B0mryhPO0KJrpyi/C3wqL8zllgdn0
Syv83yFoGT0g8iQkcFfPOnejneHg4743c9RNhl7sBAZEMYyz7EWIDTC1NsIYVAkf/4VDpQwhasBO
2h68Wne4lpuhcWuYh2HEjHmiiT+vQ69anO40e/G9FgettSRReTL3lcVC4MIfvHiMFSDRx+XWJzy7
oZ1QZWIEHbXOUqzJ1EkJTh6XMIN7Asld9sCi6Y945lVgRdxO+3jB/bsyC9e7y2IwZRSH5a3Xizx9
bDZPLGtfxWOsVbScwbjAF5ctm3edZglzPzIYzNFWJgv86LYntu+n36qrH5IlKsAn0E2OEkZr4xrt
b4r7rrKm37uP+cQ/yl3+pvF0EvLCg6ntwMQziffQDyfxWiwZ/jIOZeubPTvoefY+HW0288rQK/eC
/2Wh2ksDZnl88PEBae2gfZohbJnYuLWq/QTMUPbgOCZihXBk3illJq/XmgJ1iEce2mCwe1TFSK7l
tPFCr3qqRa+ZA25Cn/SHgSmLGzyCzdXdVRY1vSnUaGPxxbE2gCXbHq4ceAKyN9fJ7wLiZ3GCbZZ3
S9Oc5ktgjEwgVw0LL52lDDqH/Na00NrM66hGtuswhf+kJZOOqbDBCbA4QAAA7y+ZTCQMvO9s+g+n
JVf3Otymgo228QeJaA6Z+2YhEptdDrKf4emYQGlQ8Kz07SvURYuSGKdPDg9MXnBwyn1Tpw1q3KqK
ALv7OmKTiVJO8P6lLrKxAcJYi/AZ8YPbVq2r+FiH0u2I+TZV082Bu16JXsp6o5ZXcN7GrI9b8kD7
vIcOVz8zK/Ybjav98BzLFu5g8444T4aYhKHYuiDaLfmtIkUrzv+06AN+eD9WQhY8XQ/fdcS8im1I
HMujRcQrayxV2s64fCzN6ONMzMUKavGzq9v1DOclqhlturkWnlEID9bNdO7jS/UsslBZCwz4wwLh
l0QcH6faHYLlzxfknWlJcFCDt3/qPhcGw4Wrq9CYcwR1HTy9stWkJiKDdsM9KceP6Qoxl+LYGATG
FitAB5AgC/Wn/8/22ahnGUZ7aKETn14vJ6GlbnIp5B6V7E/d0eITs3R9Rr4WvPI7HI2vrx2JkS5k
VDZejrwOVG1rK6pSuGDD+gpaCbTkW6pVSTFv6kbgAIPdj9nnqYMh7XEDoY2plseo5l8Z8JoXnwUk
54d/hdtcR5TYPdFpu8CK6wMGdkJjM+b0SjUNj8WhLZYHcnikLlpGszEIngxgUoAWso7g3e5nQM3N
hNyyTHn8vR0YvpVYbvyrg2SuL8keQ3tnK/kBgTaAnx3HI2WmdzxKanj3Oybp07QMDRcby7pXNa8s
RtuG2V1v0amKbKyxK1Cxjb4cmvJMSZ14+fS9wlVOeo6XEFxPdyOPqsJpG7GrFNkQ5ZOwjqRlwPP/
/9PNKkn9M3CTpIcVJo91zPisW/mCPYKjVA/WG0w3S5lOqVCLBFJpWFF28JKAB8SMx883lfjd9LXk
ioZDMs3Tn1RiaDdDDgd+CnvslsYeLFVhCphgbM1Hxh8SHkmkOk4OCMvS6/ZMhHuBp1ZQm/0poVub
C3NgubTEYC+Pq+F4SOJ8zkSjEYrL42u0AXPAzw6CLq8ruoxYb/6q+IlcQ01HVAXMSOG/hZnBLfFv
arbDIicoIdBtAKju52S6XT23+GmIEjZQ3WxT7G14ORA3Zc+SHrgAXceYV7DbwbFyhGz6S6oE3rNY
nKg7uDZR+g/8uX5l/LTdW0hMDYBZCJYKoypnmDYdRpmQ4kqfzkMQSLIkCp13zru794PfnphzbGw4
Ut8cIbgHiz9PFvE1paZW7xwHP9RQMW23nhqlUQ7dWTf9FxuDFXtOzaxVYtuWMbSB0BHeeAfCyoep
J5Clkw13HAGFEL02cKX/ReTOFoCBflEcoKHDg+3pastWYDUblwttyPNhatr/0ZEpQHH5NUQjR0fR
JG+udAb612Ymy0zTa5J1SWoPGOJJ72bHju6HFpSzekqZwbziX5HAEyJfAtkh+zhIzuxD6wUEJEPz
f/c4xb1cIv2cpIAuFHUpr8/AQGyQ//7difZ7u2qPO1ZeH0EL9bapewlRQgxIm5pKEwaJqiWwOB5D
+5rTPtsZ1oiKj4NvnnCukBPXO6GjlCWmBXEpJzXZrnkMdgw6qpxnwYDShqeNNJSV2QSLSKWHLx2m
IegVQELYnA0ndW4G5l/RoZzYM1g6u9un2qVL70NVohUDbJkWJfUV9sx0+LsGzzTXtaXxWkcfWZw5
iAoohWQR4tAdV8NJ2yeH5IKxHWbdfI3h/taL+7xVig8VE3waAo4r9N9VPpDCpk+Ri3ZVLlT1SEZe
A7rAfz7F2hLtap2fv8urwy8y3K9lBxxE2A4FEn5CHkw6pQxq0tlhW6irrKoIWUoA+X/HZDMCnT1s
0RMNW9YJLs2I0Byf46huKlIfSaN+dqr9nv9hq4011GPWd6iV/oP260cDjjpIKM4D8qs9GdqRqz3e
DSBVJb01DsjCR1DPmFc5Bx0exG5OMFc9WsQsuA67drUuPvCNZJqcngJzx/peDBdW50UdsHFofVAM
248mhZAzJfErcYOZsjmmbhz9gPd8bNTQyYjlSyBwu0wWZMURkOrEtBdG7G3zUKrx11wj+GuwNSwS
4Qf0dJSJb1nFSU5QkD0yIFYq1LU6XqOveZiAxX9MD528huj18rXtu14kngyzdx4R7/A7ttYnEuM+
c5p0zaeceDLNTvZds/uD4U7ZfomV0RDic/1vqm5j57NlXubLcICviYJnw1xGX+M3TJdVqgvDlUUR
F/cvVO2wXZab+GmaKsB5jz4nUaSJNHp8s1cRyv1vdLg9aeSe/9ic6ExJ2HgBABjkEH8eq/c6fOLC
jLEScapevU+DLCihkewNS1o+Qtq09D1O4IGVbc9dr3Ax/Ckui3Z1UmSVgJUK14CgvDA96MDrOyo7
3P+d81si0i0vDpOxXrH8Npc0kH9O4SyO1ivgGaP01OXDA/Qq5WWIalmXQXQpaZ/jbcY9u4FLp2nf
HH+QzCE65vUCnNVNAF7w8QaXeagjx6KSLtQv9uCAE+wuIzsAlEe+i0yxililuFhjM79BoWZpZGmP
jgvCuhOa8yFxuvofMwNdO/JbXikZ7RKdLXp2CzBeHeKy0OKOQ/p+qM6tHvHfmMTK8phaUyxnyanc
ixBDke51Sv+v1rmJeIjlVKZQNVRlYaEbu27CMaSHMX45/Ym8nUnzEYeHZcezYohQtAjhVNrhUpD+
qLc3bryMUHuMb+V5gi8J7LvJEvBrRm10ubzgi9GLPv+x9n9Hf8LgXR/60RLa67/3RFxrcqF1auwc
50chFjTPnvEYvDtSOrAwHdHLYVESKWs76I3QFWIlrUWYlKfEAbg02QNTQSLIuhtTq/5UO7o64pJ1
Wz+LHKP5BbeHs8qKueMyw2XvW72Zh01xLTwlFgPJPKpbQ5rBBRowMOvnciHRaoB6xyiMLG4B4q/p
YCULlhoivJt2iKmIPI1ZyaNN2+0SbePqqD9JInU9YeUs2zLjUKnfX80FDiq2BjSNODLPiD8mC+HO
Vr8YpkKk4ef6ApA2F+sxaDnh5/qjoDJz4vls/q/n0c/7ruWuHVcFrtAK7/8us80WryZEjPmL814N
bK2DY2Jv/LjWjswvB+KKsmKg7aBhIuBwEUwAoZ3Syq4J0Q+S0ZMWEl3qsPkt4IHPY0J4QaedMv1J
xFyYmlfi/VUAirXuMO1ajeQIVawgEvCbyaCnksNra84m4mCwPZoTM8rgxI9Gnip+LHGK/AFN0xo+
eV0UgKl/OD8Nmwfi35P80CTyIyd7iEuLEFgkUGosR8Vt4vrIuUT10QL/GQmxuw5cQq1jaRrRq9Ri
LbtD6jeSIMQQikymhEyqjfVHoUjoWRLp89yEApLHJ/tP+8g/R7OqaNERKpMwJg6Bw/x8vtMypKYf
NFA4c9wCivHN2TDwH0mxZnPVn9HpFr88OpDghY6MUDpCVSqrsR/3hK/fU2Inhp32u5+AH3q/jjda
g+40wDX2Wejo9+bk1Hn4DjtBagYNMqoPoTP9tLWTW4kDUSSsn18u2OhfaTusG8YAJPIpl9RFG3DJ
kyciLvqkfj6xs8cffNomAnV0szw2/a6Ct/GSUzX1xkBLBB41yiEK58F84rnxoLqn19gfEKQalzUV
64L7bgogFaHeJCDvi9LQEXoVP2H0eiNTKPwO0P5UNs4BbfROQjCBw/BOWXLZz8+aSP1nhLaFSh4x
tTX5nyVwhoQ2iQ0otmTGOzMSIzbg8tDWJESwdDScNhmpxHJ6aionN2xpE81HL2jljLZZ3/xAtySi
XJpOP0UYSSCchPjttMDn77OslpIBQfsjpCcvCe+CfyG02jJRIuQOWAKFGubwtNqCoV6kUrCf2DmZ
wyf+S+CC3HSLYr6yYTCrUet445OoqdVJOv6pZZKeQhT40JiCNRZY3EZR5r0H2+ZAI292mAl+J5C+
kFPO9PkL47UyU1bVZV0mUyROW37A6zxQkUGKT7twKqRHMcXBcBboNajNaqAjvyUeBr2Y+t3UiP/y
tIRjkDV2BIGainYc4aP6hR5Xp4dxAICiyhdAPMv/KXqgYXLyWnUtGJXWp90NK/FuPZ8NAc9UcQoF
8mTAtMaPW2B6EstZL1zQt09E42yjPrAMgH2uLeiDGkT1/4+eUKdteFnEiBIqRcTWAHk1mLIn5cBf
TC1TNemuy6U32KfTdqHv+c1ZaZCkGfTGX588FzL5UL7sH+JEg5/m2UGE/WvPHKg5q2aCi2MErBtA
K2NXpoluCdMtqymWCqdsSBN682a5Ap68+cSYCy9M69EmHx9sJQkfqLaw1JBEDMr+ETBMA5PBJPhq
KDka89/rawgDfFzaZUb4vZ5aGP4eWfInGZxQScBdYh8Lq75Z4/s/t2/kdtaMv9S6vVc8f+SXt+cJ
O36EBUgxyXonhqXdU2uYySkQ8B1xMWdoGrLlYYjNZcQaCcGYVhbo9LkjKrcVMyFXS6GKGix/BUxX
s3QqkGefw4tqTJtVlYmBxF+z4WDUtIKN5ZC/42VoTgvejrFwmaI1871EiF51DChQsTXeOmCHDG5m
YXisD5bTOoxlSLqx92kJiZHS4AUivgJczIS8V/UC3ETxrs1eUV2/O7CMIXpEGz+/pE9wEKKJEAce
IaxqCGAAaIUJoSBD9VEm/bETmhfoNC9h4e//QuZJq8oObthjIiW8xGw6pWRlSk+KI4VJhgZblCsq
85R/34WmiyIAzq6n8mm8YIKOKpvwDTsjdMY7T0X8OCsXCVocXj0wBfmQu8KDE2vGWX4qDdv55twp
JSJkjJFNqDQRTlvv6jrwexe7oRdvdipk5S3GSEqYtxnYnMxT0KLSm7HJhV3mADH3TMTCeSbVkd0X
I6FkgHaPE01tCX9IaCZf7eCmojTFKlwJ4tNkFQGeuXIUfN7DdD9ZN1JxiYQ7JRkQdQb4agrwfnMO
efZkCcs6moELQgaC2JbgZC+QKL6TBOUzv+s6OtvDL3CsBH2+beLi6Pbm/fn339lY1mVEdyjk0Qb5
nzWShbqx+3T+oaXOw3flj3zqI1WCr6Wf4CHy4+UfZUuGGU7rcxnCk0D0d8jwKCgUZlzq6DipNZ+i
802cb/kRWitZerRI4XHaEgIiwk3KVEZixGsT+6Of7qGxsFvawuDHpZgPiymlTAIecOCACZ0X8uGJ
RwomPNDIbQHHssPMNHH4W50Z8UZkTzgl2ODVO7DD1ttXujL2t2nIbufV4YheZtGN1tkqdPunj+YO
FvuYTgdefBqJoVm7nA09cax5BCA2HubJpgwKQw+TsszsAgAAUGKWbn8pDzw5bktj2yBP/vit8z0c
B6Y0OlFtmpw2Qfpx6zp5i8YYMqZkvg0x8MP430hAFFDNTR/sHeoyk3FNRF8Z2H2HSFbVj88o5oFu
4fFz47ApjSNWBVno6OELPVjdSxfxA4naEHyYyln+nwvJUz9XdE8QMIRnNiOtPPuhMb6X4io8Oqbg
N4iLeLYKykfKvLrUTRQPKqljTlfJXm3GOtX3is2Nr/tOw++j+tTTHcBIPFmhggw+mvhV1wjvxMMC
pCsHZWpN9hvvrgsCdtWElkC/7KtIgmvBwla07+krE/SmD3BgqJ/UKVcSzqQmiAs1I8/1ziq4fwXn
AxmVFK5c4gswTVlpRhDuitFiFQLlhfQ2idRbiuWCXOfEySUIw9+y7fKd1nOTHBLto522zNkT1d84
+kA6xjZrNbiUDUv++4KmJBsn/OoPgHTb7Qvjdkso9mkIFqKw68xiuIV0zu0G4Z3rMcPoVuOKtgDO
UXyuQekzZdLyqKJ4BBgSrknlsS1bL/1kzHZ063w3pLT88Kk9UJgcJ7sbf5aG5W/gGIKmtINOQMcA
2ze2ggWh5DxXW+uE/RA7MBPu1kVv3D3Bwa1xyNk74yHLk6A+U4wkjUImCGkBr8bNBah2w23dyd/h
1ga768fxWvxJKiodIPmvtT4RlKl8cfzYYUMRuQIMnu5V5RobdLhbtRp6oYEN4lW0TzZbQbO64Y3k
ci5gGZkGD542/47kthJz2EWqgZCjELGFsH0LPFGakmqHIs/8JmjqeYi3PucpjZwJ8eF5jzxqIXgW
oU/+yZoP43TRuhtBJ2kahWFMFhLGWCXGdXld9xQQ4i7ns2HABuCJScBxQNEIjHVNlyONujwFxrfS
wP+acZ5QXxI8oFUD3U5uB477jmWPVqbcF+p3rgwdsX2Hh/HzFVmiMCdlDlmAkt3xvEanC+NvsNyb
ka6+t0cVAeXeJp+bDIWfrU33BIqTRiR2tHheXVY/2oX4lzYtCyfwgC9osZogFi6ERObzIxdWnCe3
Wtn+mTJ6XbysPZaDUeFoPYGhMHKi8rEcx0cFfdsI28QEXYVUgM1zzh5hIbg4mAI5CbohwkJKCNjz
gGOaFphqg5yKVh6oFkI/lP6VIeRU/dD2koj0eN82bqaVBZuUd2SuQu0KM8T1r2JAp5SVY0IoDi8k
8NVfOYAoP61/98z8RTu/BxTC7MSyyGI6hCmgXbKcnHKa3oS1Egl512yEP3FMyzoITDwufuP3JIIG
WG2L2tTUC+Km+34aC6qARPTf+rtiedd9ptpK5FUJK15EPTmR/Q4SW8w3ypSYLO+wan7kr9nm+0op
j87yFLWMw21cST7Hhv8k1H37hT2FPHnC5/VHN+RvFTrod5spArPTPvu8wsUFi+HBIGJwdQWQWX++
/XoH1Hx2+i+M1lq9xcZHXKvq1oR3kB4T7JeMt1CtEVqSGw5ivudMmc5KXpPsVV6Fn7hdrrxdFTtI
gTB+eS2azGF1PL+FmcPI0sbWh8A0KpjcVwgS1YBQEDK26KvfG3Zhulu+IKQm7awwbjGYtBgva4xG
p7CRj89wbipcQ5D8gSsj+uWGGhaiEhRNPYMFNcd+i+VwyDPtpkM5ndBxSq58R9hEb2x867nsyefK
2qwf9hB+MdUAXqhKPJrexXwmNPBuaKghwUhvr4cuV27bivlWvi1oFXxji8f7wQWMhu8qzSvmTcvU
IIimmVhbG+Klug9s3i9wbF/zj9TjB1Bt5955g6mhb5Qx8NTPIbWzdXvpCQmEISeMSxvCyXEKNhqh
ttMhkZy1ORQiWEJv96sJqKCVgA0RTlAapFUEAUmlVMbKobuzkCA1vnz8c2Jf5Jy69iruYeH486W4
+PmA9uX2ELA/0UbuQFFXlH2V3dvoRMETAlR9R0P4lwYVjAcYST12VsDObKGdnL7iqNFXa86xRn1b
9SQOiaAynJXZxaDRjsNCWjoMqm96xVi4YcosDHW8/xu/ms1a5bGOkbo03oe7AovWe12BDVYITBkP
HYfIl9TihbzPnX4mkC0Cwo2AzW6nFULyNCF/UaYAbfjjdNn2h/aLTEjBLvqn1qHJ03BmAQA79TuF
MZ5PzTZZ5J85XYZqIKau+G7YNYD0vH2Ele3ACq5Dde503BSA/VBGc2RlzzsMjc8/wy3m4Wod+y5y
A3xK4D4Ehrl3+44XFSiGurKCGCoG2b5mgN8GeK4P4htLY5H3zZTDZDZlfU6jUfNOu/QjIEHkurMT
x2EMdYoTkPRbi/5itQJTnsZVQWHwwxplDJ2/AzT2EDso2jCOHk+vyQv2twH2hgVwAqBlTeslxJ8c
/TLVU3iLpNYZfjdtqcNRnrnnVNtiosvs32LNJGFUdFVH54mNSCiIcsy/27Is/UHf+NV9MfRc3q41
JX8hrlq58/Q7N4yyuwV5qWvyhAI46UHbxbE4GP6DNkqWDFYVpRfZegfHRa5MUMYq8xZYyqb8cRJZ
aM9pp99Ynen7l7bBY1n+XYQJZqhJo1ROwIjP9o44PIiSXqBxiby1iidcaovBCq42SFfju+pDJCrL
xkskyRi0H9NHQT4CthNkzIb4mtw9cTR3usAGNl10X03xWJyWPimxC6OeIbDIuTl7XAlBIEcuPKiG
oTs6khbtI2Jqw9gQ14ex/nscqWaPKpSNSYR4I14jTh0OBdLES4dM2mNoPn4MTZx6dGWbbRhAQwo9
2ZBRQizORdrfoKllS0gVhuodT4lAZz3r2ODY+tOcZY2cmKAFGNXzk9dlNZ8/lGXosoPmcguwQf+b
L1AnDfmW7kUeKh5YuUXBPFqYAovaXJgwzny+PP1WpPfJtO6pRJBYj9KCQi8R51QkSJNmm8+k7OEw
DcLATr1wp4oxDWfTQd0ZtQrWm91yJOJ+8Yxrg4TjMJbjfypL3honJ6cX1sBO5KWEKmxXlK7YgngB
X8NJsMG11oq1a6aCo3QmI1o2leJ4xPbMrIfe1iW/CVvtIBg0OzX+606Tu/3AMef0ECbLDjX4uj6L
8JIe+p199nEJxmFBJs9qAUjvolCdy0F7i++rf9/IGc0soliWbVTgUnAQhTBe/K2umMfXVMEgXbJa
qq6wN5GVqFHtCaXBz8jhTBbR34N+qIpQ6scJLwuRg8D3P2y4vwLy1HuNIwlB33HdmKHsN8zHTWdH
P+4cLsPMya1/6xh3LMcKHWukW1aOHysWzhpryFngQs3LJFSN4rbzqeI87hLorSCQamYaOx0y9L6p
DweTRTotMnr6rA+4RQvarLna/Y4ECn5I8Rhm19AeKd/PRpHb00twTJiqBwOQFxbfhwIfk6UZQdGF
iqCtXBIViECWag9eotJL9/0J3W9mAGYGpUCmi5/hBBNT8qqVspKM/pogtRqOzCwFfv/H5iDXHcV5
VKC9EKBOOZOo3QiDl5/RDqYbRGj5wfXJAbf2GYyw6cl2h4cixJaw3Wkf1wqpvTWV9SECtk+TI1Na
MyS/TLZgvqArduGwM0VKZzKnH0VovD62G0Vyk77O00wyWMKWuubGAtZU3IikVHKNyi01Q0X7hv7K
hNDCLIVfIEcOUUJctB00i3mqNy54bFuuSKryrUqwjLuN9dZT32qU/sRPZ2TzFEk+wjoJhmoSrn/X
EHpX5u3RM96ri9jGCOUoUdeUac2P7eW9DjrvLGK0SwtQrVTsZYRzNvRpsyPNxvFkeNa4dTKRU4wG
c/UxnE02z2LUW+ADq/mTNkgQqxeCktZYqZz+6UFVHckQ5o6CXk9gaCd24xGF0UthgP0SkQxIlCwj
tf2c7q0dDcd5qwDHesyOG+cgA3HCCx+K5YVAXTHvhEwM9lhg4LXDWyZUKlJe7dCND0CtaCXtB/rd
/LzomZ9XZv4QsLdB9KyCRBKsRzmZroaACCdvdoO0xKp5dbOk8wzTLMApe3h+/K7vbRedwDLtYzoh
UnWSQQshstk//EX/vbUg5x5I7R5tmhMDRMnAkbMB26is6cMcLNSWXXGwRNFLvXd639mwe375Wd3H
5W0jUtfBKXgq6pN4meJz5b195K9ROtb4Ou/1WndX2hpb04lG2lyZq0ci491Wt0exaIDtnWsK/CjA
1qHLdYc5ls5/KVNkUaCjhiR1xs/odP+OffJD7MBNvtk2sDDfsERmusoMWrUO2Ng8ZpBi9oGi3I/R
9/6v9U4aPQ/D1PRJkgX6GJo8Ofdmqxa+rUzrRbO9ON/biQSh09tJ26Ezgaa7g7+94Hmakyb51Irv
M+Di4S3nI15qDzFe62GwfWVfW+aAznEHJKlKJ7xCd8nVpiAfeQ7Kidb4+K0sukbLc5HbxMTEu93D
KjsIrkcA5DQAj8OW/pszp+534ChoAOOxYFTsYw63orKWHlsj0Li+tKHJe8aqK3HKECpt8E0FXhmA
3NzO/XOmKDPtCiZiQHSmVxcc505j96nf4r5QcFtrWID4CYH2SUpSda71WNC/G38WsSBapBjYaWAH
TVYXS50bDIoYkr5J1HgBaybDrHbWWRodGjbdz+QO7HL1yOdjVy4dqTVWy1LspLEgfU2KTvaHGlic
O5Cs4v16xvW3FivORVClJpg1LbmUKJV6SV+UoDLgusm+bwLQ283/a2sZwFw7OX2NOEJR/19tXy9p
DTx5FxrIIPOsLxZEbtaEYD7jVa0P/ZxDWmB7lDmH/FTNsfi4ZHleLDkL4av+QzOUK92Q4XpiNKlU
VWBQTuQCznIvhaSjyOoVmPOIuNXbiYYNDvRl0pxjH3vL+kZGNLALgANh4pQmLBtCRM02PA1Zwoz/
+KsuxPnCtackDtjOoQnWH3LOkCIfWv0okH23HMnOqdY08uC7Dyyr0LhJeKn4JuzpKFGfjlWAwSKL
i0xav1B2pCZ5yFyTmcxUAa8tMiutErtL3a9fRHgXVCNzzJZE9MP2dV2JZXqcx2DlywTKMaaXLufK
thyOZ1e9PSCp7jv/4Kk/REN/hbtF3nN3Z85vLlI3RMdPPSVOJV1W2i1eNhqlAik0nLN0Kr4Xkwii
Z8z5LHBSkiyHER2NOz5J8yG6Saa7Hmw74CrfL2ijITK5Ogfx1+2I3vXbDw4EDpeFGHnj3znHCkIN
1eXf/kNpZy4VantTk0c5ADRaNFfY4qlU7D/Nbei1bDkD2udrN6XSJGLZGPK00Ooggee+lXLoPpgI
I/jv9FsuaYUqzdbL7zQbIKnaJgmd8FIU+nc8LE0loGfLj2djKO9Whaqz06DjAVfokqzidmRwrm/b
TPcWt8kIDz2NmKa+FDo0/uzxt5G4ZVRGqRZGnbQm8YVAk11KKTzbN+kG5a9kiHTkjr2hhmnZ2LEQ
B3LKIkR34v5YA0LHfvgXJTM/FT6yXGg4K6tuD+3h1QhGEjC6UEQej0th5v9rejRRJZOZfXKuOAxC
AlwKKv4yjknfyvw/KXvrNqilLrErgHqNFZ0QKiGbcjhqZXBbkUGm8LzZgfxYCCXwFFX8yj/0WY+e
3XM7AP9Avb9xS2REj73kamrzGlUj7xSs1+LpYvJOZ2f21KHBiC2Lc3g3admFBe1Qw1AyYkuClRoL
OHW1im/JdoOi48yjNQDqVZr/FNsIVy/kGzMsvS89TfiZG6Notczo2EdX4jeBBYrYoOlheqqHmhBA
zWvBHIfwqhNQu3X3imL9CDvaq2rkQeNjuwpa98E3Hg7vkgtYpAYRWpbONsKm7btsXArpTC4sgGLj
psscX2c3ThcwE8awfFNtqcsa5GnvdKEqGoDmHiYPP7PRDVMl0D1AkaX73uUlYKt57l1U/jUbz023
ID447UC8R+KLB+c+Fs+VVfHZhhxQHsHoqRuu3FbTbRN0xbaBudZ64An2cywqb913C+tsgY8W3pay
2hQiOIusJEtv7Qx55cQvRLI4Peu/B99hEeG7Jx5i6iAkOEDtyEMdCFkiSoVbXB1oRzPUlddxP2Bd
YoPB0rk2kcguDJWNSBC54KHJiSxf+baXHqaLklUsmp0HUxK7ldI8YGg0ktk5WLaommPSXOn1sZX6
6qaQLPmvkWf7jLGt6azjTqKwke5JQaZdW9fwljru+UK9+umJQWrWfyr9nm/TPKiXAolu7d/A89Ih
amyFtZTI/sgQ5RgOSn5VnuIjKVjY7Cc4RBR4DR4HF+i0ym6snwVj7RI4OxWsJHMKBCezDBze8rKc
vngtm/07nMUw/sY2EsUvCqSj8xguXN0hY1H5NPV9uALJnfUCdwRMCMPjL8j4wdamdvxvT17EPZEg
QDUFGnXUSW/8Quu9onhuWqKru306EffkoIASCZE3VpgGL293+5UiexTcWoiC+EM4PQdfRbqHOD/F
xEApnbbAGR2A4wrFm/8D8H5BB7sd+b39JwcLVM0Ms64WMWcy+veQS7pa6vpnzX7RAA95A+Sz9weB
DCKVHMPLmNiwu9AaTocfA6b5MlW/9Zg+qxLD98myvaakiQAP2UwU+BSvIP4oi0C5+sKLaoodMrM3
uMbQhh1Yi/HtqfSlr82UffKuW1M7KirHiwquTs7wDpdK2vPMnW6ioF9C0ZJH+3LB+uIbQwEvhFtj
/vbR0cCkwoUfqnOXjoO2eWAfMtSbD5gonyre2R1oir/0PlXQdMH/KNeGL48IIoyD94mCs48i5shS
4NMju7YCHyNLt2fhSjVbLX/QWK0lKxuIt1gos1lECiCKbjwjsEl11hIf4+MPNrlCBj5gV7v/RYMZ
D39jMlbJjTJFL8BEDH37xZzWHScIg8q8OxdWKzrJb/b+diJB5nl2LV8Q8pHbf2eP2uRpnVGZEEjY
fcZ0LNsdvI5kwh2Q/Ry2UtPx/WyJTvhtT319mh070DqBzVa4yaGAZjl6uWAz07jDE6Z1t/XZXh5Q
O3KqEN/711+tRmMaYhhurHgWZxWT5F7k7wk8OS5pERPBgk4G8qfaysL0T1vljiInpupd8Fz74MHE
ic7OsbYcEHgU8vldsQzvxIiqJkrerQI7f3VA4J1TvQEMepqnSl6P4Ui4yGNZEjvE9Aky9myrgBcG
jFqlOd1Y6pZq3F6BuFYMQjLnBarDCS/NVIoEgGzVbw9zpJL1wdAi7I+3hlmfDyPYCjzCXGJtG+Wy
xTabngRE60zD3isNEu4SkCMTqNA8Odukgcn4HV+dKC13/t5eb9lgDcs2hqVYKOFNUoGXoqGlWxHg
INv2NGtHdVrP3XrHg/7UAMAeHG/klBphZLb2uPb1Lzm8mzkSR/XOfEVQ/9KtRmAJ4nw4anwwSMxW
VDePsvX4kkt4F8AWzfQlSkb4usm9V7Hz87NNCFOfKJk/iwCuyzuUftd+te96fx1tMwRur9I1OI6Y
ON1KdNbOn13IzLGYh24qGAnNhP9G4ir/FDmT9r8J+qIAImxIUYxAW9DeM4IG50kaZ9OdeCVtrpk6
sLClp/WRWuaS8yW+0BV+TOPaE9xavrGTx+5D7xN0cL7//bBQiIKein4irnvbfkMC2VvoJk9qiAdX
9TsytjgZbmiyCCkz5A0HAcIkHMqjAecB6zdzEHn8PhS3Knz4Nv8wky4lcFY8eXwZVF3jAgXQtDyV
0s0lM7epPxi31PrSaCBH71o6Z8R6RhZ24CQlJU8nlC+4G530iepQqP1sVfSDsufeX5LTE4/1TGPN
SxbI+Ltf4rv+4K8PP8z2ciDYx1aMpE6re5Xgt/iVRzi2DWW6pieXYVrwNZDXJWwAs+SeVIFJkePc
HjTOTQz7rd4NvY1KAhgWQsi/XEwvhjqWmDHW4MDBO8xb5O4flxhlXE6dQ1Qi5P8bdUn8+OqDo7Y9
3xzEkMwJRZ5UiouL9r80fxR1HJhl8r1PDFc4L84CRd0kdmcZyxpv0UEW/mUlXmwDCGkqB84ppS0F
+aUidTX5B4vzKYf4c15jSTWNHStFjqPOgZ4B5MPicS+2Z4m3XWoMO/F445eunui/Wu4fNkHg7b/s
GxRnTT+WzXxe6noHrLy5FTb1wNlIu3llot0fXa/4uJHT/zEWo7wpwpTRttJDFQ19JeuKlqEOUkdn
KNE/ak65GtpgK+EWJ5RyRdMWULO6EDwgwpodHgpU5k9r1NtseTY7K8YX1pyC6pIpUC8wLxhC1aGO
9ULR/S611AiTLrWTsBqv2J2YC5Qn+Rrc7P2F60FyVJkDghSJmqDqirXUxZ9Z87+1c30+RJrlJxee
nWPnUCDQTAv+oDcXAc+oCe9kpOMd82q6VonSTvFbm5+xnJYRN+ooFoNzcBn3RJI7y41o30cmeoht
YotoLUly7ylAwGM2iTRoXNHbkFhNDgN6D+MK7s0yLqqNjFf3gRN1sfNF6fQXOE8UwUBD1rMWhHm0
7Ntvx3KpgvG0u3YYXHucTymRTGIXRhZ9eJDfk10vm+t8v41t8HdyEysKlMvqh3YjBLDrlRUbDfAZ
Fk1gS8lbojAayYH64SWqQuZn5+QziREAIFkhka8vXk0/lO2yi9W3xiVaHfebRso0lc+OgY0N4xEj
QqI13faeiPwY5lAk3ouaGCgcWP0rP3U5ubqBs4d5579UEKt21GNhtmJe1hQcyNobSB7Y4dAdA0DG
lVkbILTFFqtG7cg8MuI8prZ3aMqBJPub6L8UwwvHFTx/8B9WV0P2RFNYMSeOd6HvX6FC35Cof9/U
CmQ1h22ytOtuhQDCR4HPChVi/CujJvf2O76vBQCb96Fn2xniJAUfTMuBFud5AqP/1VirVqI8aG1T
J9Putm68+Ka/zp0g0w0Ha/jpTdWJc1sgOr+JhGyR61N1vktdZ7boZHhkqdDufKE9rTgePWhLHFvI
QvwLedVzawbFacwGlK2ImzSCLJqfF5eEeuHNLtD+n7FvdEJL5/B/z6bicOGdpv4/mcAxSku9ob6L
TS16htVNSzqCrLxmQmv4x6tPekeL0ZLHtdVfcL9HAipNtdrvEp3CkwK9WxLXgR4FedSNJDmC9pzh
SyqtwaSDh1NvuCqi71m94lq7HFxcuougLNOyF8nk7JA73M71QplsQ9jYNuxThno0lDRnMUi1n2iE
f8WZ+7qGeu7qkXYWEFQWyKT6RczNJVvy7R7WN488e6pptZAWO7rxtbqVuMeRCsICpM/5exapgYcD
ufr6QklTGpWRACxUM0QY7J0/pCDG+jTzqvS5tTImy6aeslByl+vaWTC1ChYANAwEE4PyjRhRGPeV
yOSlgpVIlnxMYIKA7g/k2gaVUGF3xVO0ODsZph371h0yEtUyehCnV0lRRpBuFXDsaVGzsjH5k0Zn
6Hkih8NuyvoZVJtkescdWou5qQP3eSJAYeujs9tn6ORaIlqK5G/NdZXuJlGfe5uNzaBaSCLcz8Rt
sM4bbQlROxVcdXzKtiWIHmc8H8D0yHGw6bV2vbH8WYmq4reykU2wz7+S931+38Ct8GZlqYGWmd0+
2FdVvIzcjzEKROOeBPzohnisKLOdSWb4/EMdPaTzik3srMRF3suCxuMsExbvMEaIY9lAtS2dRsoJ
HJRoyyRTtjmxB5uypj49xTO/rPKPw6Fcazo1XhKPtJfekJO2s86qWQ2MWaBiElG8OHAXAwJrJ0Qv
eNztPZS87rExIgjW51uSShau/qmBV66IUbYd72zZHSA3oZzuYyXYowzmEIgD5HHJtya3QaAcX6gX
Rb5lU/iRCPNiWTs+onZIVSrWeAct0aOuyFzNR3jAwx04+h+qgQMnVTQmBciA30q/2B8EJN6fLLAY
GXA0rGzyZ7VSt2MpXna3bnJ9SIxe7KnPrjsvXchEEQQCENhyuX8q13q4xk3HmzKAF54VdlWvvljr
oMfWx2eP9vWKUdGz/VEpkC+qV6oQNm2zoSAHeBpqGW/VKLBCultsPhIyXILA9nc3OR1jJFOYI5S8
broO2fvUrfH8tqJIxNCqD/beBSc7/eug//TniporFZsZSjLEWHmXZFELxc9mIA+TKoWcPPdYhXQg
LjxXZ2u8RlYPYnoHPVyOcCQhbZo76GZ8yVFOFHbua4rhzwurkL5LYgxzreDej0OCdjctwDz5GkjJ
q3HH61AuBVHZV4xs8lFc/jT8uTVH/Ic6OyvFtEjARW3swb1rvXse9cioau4KHSWPYGFPV8MC9pJC
8ADhmSRHZRGsRBSp2OSzNSg/IR147tioEXsPwH9Up/vZjxDTEztATwidAj9A1kAgPkk4q7rhp824
ZzBW4kPjFeBp39DsEJW2kbm8jOplzDgnF5aI1vsWRgbm36OkIJlexuDQ/wC10jE27V27ZgnT3+UL
1gWZQguSJhZseMFqXyOy9c7jdLbJz8zMK1WwSu9hPjExGlLwyOlnDNkIgVw1iSUG5LZTUnj94Cg4
EJrx47yHPj6G4/WutUa1NSo1Pih/Drs91rUIO2/0285PidoMJQ5wEnaOFQZK2FVXkizpIXe1ugU1
DllyavUNew0ZR8o6GujiOqV+oM221nB6gixcKqGqs0ZQi+k8qFSDc83Ohw/72Y8ksbFS8katHJjd
Gc6lIXH4gv0Ok1JkEdfQCqx2EmiBbzSeOfgSsPGG6xeVQBsIumH1chxC22Kfn1CXY26K+zrQTZtG
CIBbSSmHRZOv382YkA8K4WJ0Rzk48TxDT/3G58w1RZitAwV09GmctOIOic88sdlIquB3wlyY8+6C
jGA0B+Z9sIreWrxgEJFw030AnlZZZ2kjBF2RWw27sZz9974YLc9zl0Z+VlrDlm+6Z/WhsjVD4TPa
VJq4LCy8QtFm2bM9k+EXCQCgZBG4pB0OUpLj2APQB3TpUdt2mfwBF2unfmqowODCtydUHnlHyYr8
0O09rijzWSY8Wx7txmLPp8owjMf9r5KWRjaIOIuSZw2LxGN/fWMdxxn2zcnJjV97V5tEuEp9Z8dH
VdY0mFX75aT1FXAMaQKr26Hp4BjEmOB/aSntlHEtnhfMRVWiKFcYD/OYzwtfk/VdwByC9zbBtPKe
BMVs77uZ8CTLv/Wtd9Lgq7UqjzeTtw8f4v6mbwFJpO74l41T9TcwxOu0y5Ho8xpNNYgkq71LpChL
WJ96n1C9cGbNfsZCFD8W6Zh8Oy/1qkcZXNAFfHyFYcLUBV68q1y3cFtwtEQB5yaMwgPL14u1HrFc
d14vzbatP/eDaveE8O7MYa5Q+0mtLmqRRdkBYVxs88irZi0vCjTD5Ai0cYQy1FN/cZhobDPX0569
+EE+q8z/6T+71A926fMwGkZ57l0Ru58bvqdhGsUOy3dn5W47eSy7zym1z9pMayWyAmXrb8M+uGfU
3pQ03UleP1c7oMXNFQnzhB+r7867rC3wfluNqjYnpesxDrNBlb2pSNmb4RwnLiQQNeVD7lEXucLK
c74b9UkFDppF02N12D6ptWSgSRkX2D4r/JZy/GaEkSUixILEFrYQ00nLG0nrSnOP4wNPbiUXDKJr
nTM2HtaB5bvvYWkb8J8TpqsS3MNbEEstQjeszhE+FyJaqAlQ45zgl87gluTuv6ePCJIN2Mg4rAXj
eCObE4ZHJLMfayRJGMW24JXMrCsoX0R3tLtQe0hdVzYTtAr8J3rIDuclov7N0K42jXA72xjc9Dbx
QMZ2mpiEyo30I21VnFWAeBeLBlPtzIxdwPmdXuck+GCT0IjIK9vuTiwfYXEjz/8SehQEBx+Q1asT
PTxsYOPSBpOqjffiBBwbuCYPPzChstrCuGugG3hFnkOHh22pB17ymFdpa/hfzcaJRZqo1MDJjx45
foQVwRU4R3Lf7kD6Hv/qDIo0+fps9jZDn6CyfEsGHXRaYAXkalral7VpKrIWco2qavfPVqVpIxqF
V77waiKYnwyzBC8pUDBE0kkUEkE6xCFRZP/AIXXZiOgLtLQoble76w22wiU4eAaGSo1NF9eFfb6l
hIkixJGGkHflqTXUOkEY4EdhdLUc9hf6NSH/YFzp0jyJJvmkRc+zOeA91VAMCtUWXxvNuQX2QQS/
ZeYPDf7V3NrZKSi6vp0XPGT3iUNwJKRppVAzwoAHB3OQ1Q84VSWxrmp/H9LdxJRS/bRSbb36Xx8Y
Hm9PbUBRiipMBLwE+9TD0Zi5kSd0Nk7m73xV62gBPAeHcWEIovQQ/jx9bDDDwGSx0Oc16cIAHwjQ
pdHYG1QRiY12BdblWDqeSdkeaZm53Ij8aRGA8+VtwJgayf+AZlJd4KTau8ZtuJWu2lDpbOweEKKi
vWAOqUgILfR7W82w5OsM1s/mKJZjAeswS8dbayu1rFzRJ+4fzEtDUT/NTazF2vU1bs5PnacMPSHQ
cDvkKhpg8+4yZR8f00Df2w+BaT5eAAVQjbhHW4H5dqFz5dhXHa7fNhfK//imobnRQxi+Jk2KZQDP
EVCM8v1xwAmRGMED3ENX5+IkIS8fGeItQmcZXp4n4Qc10iP3WH6ZlyW2u5/HjdLjiRRqJqYP7B6S
KWKp7H+/9SYF/i7P09RxQNhIUxf2FWjGriM6cMsMWTpsHQ7NuoOXWZmkf6sR99J2ryBoNcMxxdW4
dJZIgkcZdLHOM86r6zkJEBO1UmWiz33XnmEOPZ5PfEmpHgUqP9j6zeTF4MuwaLeASyEpv7B2bApj
Ano8TYZFhAO4h/Ny7zyEOqLWzaq02MGJyrBaSves4kP95PjqRfFIHCrFqWDXNgxfqt9EYsmWnxfF
+YsMgPP1KxK+C1Jekr8O6goEPXEYrKQw8rjS7RjW5/HSu/0QNXup6FoYwv0coXyI8mwYBRaEXaEg
J4cHXDMBV+KzYpqXqA9oqaOezUA3vaIg7K1BuKlhXDVd2sl6E+DuC+fqqC4dHF9aQ1gpUPB9CsD+
fyPrNZxessA5qGf2HYlzClNFTKeOCWSF9chSBmq/ik8SngF/UY4R8nQMTnM+FRE5qEAG+yIIJLnA
1pOIo4hKSIHStiGnsuApjO3u9UpsYbgMDPhh5E1JUD+cEILLE6O4IDb9TWv06p6+L6DZ8XrPyCBO
R2LHJ9qDmKkkpnHICZDa8WB7OuKIorC1AvHR10sPm6lPYkbllQ+x4sPRG3zAbzcnanwDgoYVHW3O
3KCOKvS0DTEYbWx3vlXkIjA/DVpQQfIv0fCWu3kxAM7nnnHjesirscu5YJFUVsbhgWHaFQZDkSVp
ozdOPOhDHXKpxfYYwER3mRmJvhKzuw7CjThGOIvaV89lIxUVfj22UYrYDg+kBH6unwhfue5Ei1/Y
p3YvUNKQUMQ5qMmPDoXVQrysycd+ojFhxLHCekWNfeKKQ93aHKQ0uxBhMQl8U+GH1Kq44MJ5IL2w
iBYhZkkr0+1/KStOcqxQW8zyMTLzoiJwD7AyWlmIdchueNRLunpAp84wxeCEfg6BiibWPXNNwmmR
BvbjyMAJmsGCV3vom96XgEBZw/h3XpWfWX0lYMAUhJgaUSS2gHsNhQhJ9bHEzXNLf3oh+bcPGhu5
g+S8xhBYjJ+UeDoh6v6arbI9+x7Cslv1cn9531WD+BJJLVoT+qcqDXPCSWcMxrFG4gw0P+Tl6hrG
slqD3fN6Ra6xGlM/qHUMK36IUORHhSGLznqVN/mRjXtT8BcT2B2AtGbNH6u7Kxg0rmwI0Kn3+lZQ
AnAyj2OfN/e8SDS0CFamnAqYi06fdEQ2tq0HAoXPIWtVk+38pFIH3uvlHrVBtKcYas2k+PIgR7ut
FvZcLvC0hH7UwL74H1+CJq6FXDQYeaQD39JI3X1tqOP5vZERr9bsaljZsKTlK+yrz27HKpQVxJ+m
9xE+/GVGNHj53mZxV7x4nOoJ7v61NkOf7D3xgVlnNAzfL5WXgk4mOOhtH4zPj4t5pAgiqGO1JmGF
Nxnav/JMeVThItXD0VNGOjK0ZEeDE1/TIiQ5CWQ4PPzGJmkTHx1NOgyqzoPBlEdgYAcUqDo3U/q0
mIa+lmYtxTws+Rga6j6AKDuAXjJ3nXEe+uD6fLADAPFJa4gG4oL5LUYEYFc1aOO3qTAeAO8XTtEW
UpO0X2Y/dR4eFRcxHwJM7jrH3bxdBORRQ0GzK7SWthr7gM5Ee8FBnDJVNN9cklnjan/q6/2tpYDC
ib3DEGVt0qwjWW3qhDj5t37mT+W1626PqxqTQUDptpx82cAuFM9e6pOmKvSwzTRIijT3IEWI+tDI
HdkaJ4Rq7IG39WAEXBQAylDH0lH0ZyJbSTs7oN06KuZ6MRKKETr1Xu8CRvDB4mi1KKiyiCHJJss9
EYCl7/Nuv3W1KXd9sHWVqaAX1uVuY4oWX4EL0c3HTimyYf2g8Q3tbmkTU3n3jHZKqabuQPrWdnwK
oTkHYJJW6La2S2skwwMBfWo/+yXhsRWJjZ2R1wiI8fGAYiSw7X0aRI//wvRKlSYKDHMl16NNj19g
88t+jKGMaDLM9jlTCtZy95PmJhM7TbwKpIEpKyy18MzQ/njB+L8lN3CO5DffjSW2GCyDMIpSIfhb
bM9xHMngbai6T9LdBc8/doow4iQtEghU6VbIAK7Du/9uXa7g3UojIPlqaCzgYeBf6C4rpZYL46Vq
KFKB7jXgK6JfYfBQfEeQv/0ucSCxYQq/5rTbDrL6VM37WyZVUUkzQOfxXkdZhVdJbSXSyfDf+FD2
qodFqD5XypDKQ6B4KdoiCMcV+yWUIswu1pIa945PoQvufSm1OoRttyBaHbIINwQ/JYNTHh8qOB0V
n6e4jx5b87/ptI2Zzt3t05/O8LmsWox84rAHh5dPBXa2UGVA3ReGdWAYeoFlIXnuiFlWKYUTwxah
DsSJ0us2eKyNzLa5Mlu/T/dp8egoUdRfgT4U+FXc39w3tifKaW4+5kqJym//MORE8DxnVpCY8Yd+
ShhGZkxfE4QUq4oOzTXNanrJ4ig2gjMkyiWUH8LUqkkSM4u+b5SBOtB/QAEGjWMoG1WHMJgVAiMD
h7P1YXqYF998TbpH8vrtl3NkZhlru76/p+qHclRe7fFq3ltG4og5fLM0Lrbn0jjSG5VnWUl4P2ke
NYOeXmQn8hokhcraebp7PtiQduc0oTOJVBD+HykGBRS9A4130t6EdPQmj8fiSgG4OcbqRL9BZC5A
u4vuWpDu/yU86PKfqoDE2y8ezsWXidYGoju+/fCl8N+Ag/a0RD07vBl5taTw0qQrQoazhhB5tHAm
fI1tsSGySX6oU/uIthdL/yIF9SAjHmDcUkCX1Cgi5A5zO3K7DLWzYwnUajSxQ4Y2Zsx8l1aI0ijO
enkuyXLW9lx8ZrUPruJFLBYfvEs20Iz08fWFciMhIW7Breg8uLtB7BUkAYy2Z0y/JXQIWgb3gLtP
E7qVaexoAsBm41VOIkb0yAccGVOrV1AxPmzkbZMlh2jZ1KEXTEnIz66wI5UNdy/jek1c8GgGmQfn
oyvtxP+Cj4l/nDhoO3Q8etNcGi/Xtti0JEy0waS08QNyO0N2xUiwWYxDUC4p7gc0D4vj7kAa26PU
wEC0PM44V1e43GpJJIVHIIW03n9O0ZfFbw9Bmlah4nffJCQx04UEnK98blFaUDJ0h1OWH3lM19QF
U1haD1xxLRCcl0rCzYrqRQWC+M06lf7nrC8l0tbqkaIrSo7eOhEyZ63N8tb6ANdsLhM2b5GzVhEK
i42FB8NE8NfwSWcO9aPUHTcUVZEHZP7fvw15gINAqZHamLztGFj6oQTMyAg2PPtAWX3hWJS0oLtf
CXIYetNK5y1/RgC13WoDCEQhIFdhKF4jyA/WW1R2EJnRtrYj2zHnqE7/eJHSg0XO8UqeRUvaMBXy
LEqIS09tAsRkgOR5UGz3G9LtYw+tyLxqXbAU7v8tNUoDueGKVlooi0CePhWlH6XChF3YbwY3HU+R
DtfPoOfhXBuwnanEFr9Gyr1mS0H6SdYdms0CyfNQNA7qAwjclGya2czmGQWs5GbEXxfpn+zOUIgx
FCCpdYu751Er9xTRZ2cJbeiLkhda6iX2b1kTUIJyyOxOLC3nbBkcXSnY8CgAI3O2aI5fPdRd3Ye2
BIzXYMOAa5D69sye+FGR0Tx7GGo/zyACnMN7Yy0fNEq7oirOkYHomrkhr6bWTpzlZ7/93YWI8+za
XtxWl0dvsGL1E3/yNceRAJ+ybiFYXm1LYUZiyFa3CD03+nRxlhT8I62dBWGfg79osYq6wyBlzz5w
QC0kx0Ejpxu5HGvbFFPWoAXeQHIPEz7JGu3vPQzOzhBawoJleXsIemEot1NyQgXcZrRr6cAr8dXI
yEkic0UZZMwsom5JKUFMuh1GRI6tA6fyX+IXIA57CHZepNkUnL8pgLCNhnanztDa6Wb8c4PGtKoF
nM0dwifpaGsgnPuKlVR/P2LXrPJOOaa6syIwI5MSPmUY97lH9jaIazCIw52aBRPIYdQpLzbKHt2u
lsec48OtfZoipgIoH9/D63j/oBP7fYvEe6+aNckqVXcco9QET69Jh2ElyxiVWIeN6L1gNqXEh5/k
khGzK6wF2ACIaZoPtTKcwgLxoQyTuGzGpuxpZrOsZPnQf5rwMCy03PWp8745Va2P5Kn/B25wqr41
WnqR635fqQNl2rj/TuN+OthgNhqjgDra04vp52gUuhb2ZIJjttHtNNKFQ8V9/UnFh1nacBWOJx/R
T0aAcOfjwgsvxrnYPiUY6bIvhcuVIHlTM8K8AuZV4WllAEO9hsTRLBdgwV0auE00fSawKI+N0YCd
khQxo8/KtpspD6L/wSIX40Bd1WgUhjSq6Wacj/4eeXWSpAzT1qrTBKlVQcL9GkUnt+JFPdIsGEE0
8JETGYZGCqFtiM/9Fm6r9dP/LhmrhpIbCVXgjBxsDz5ro9jZvAgGkXpB5qFL0rCGJZ38vH+jvYsJ
C/RSJq65epW+2X9hd3/rSDXvyhPj4B1eBpHVZVdBIf0hvPEyDKv3JB3KUqMmM1+DMly5XdAcB78p
tBmP6zMconbC0uQaL2U570/hVsGvReOlwOMHEwjID5q7MGLkdGwQo22id0PoWdEFne3/I8arhlCf
PFbnIpa61HyqAW9zdSJDIgM6E4qC/tJD8/2BPS16g85OS6F8zBbjFoxjIDg7DJwbpSgl5SOFFBDB
tGOen0SS3odhSRBnZtd7fyrZutyY161oPy6bW7f3azfX3nJLfFO2N776MNqBMD5jhOaRDTY3a/dM
6tZq0MZVQ5S8/wKA6qFYH5EkJkPaUJ147MInfGGA/zkVlDolyqV5hk/GIbGKI0slHWzBBJVcvYhm
h52RcPsmFtgmZgJrkpcZxE09XChhnkPMn70Er0JsYShM4Qzs5Z5zIZMX10NT7tfiYxEi3TR+Q+PU
rs7aNkbO9B13wXRwS8IfILI0GXecYkpNjXlKWhMaXXV8N/V8lpTJUvynVotUqEKpbIIyRLILww/V
lnDi0iQQ8xhqlhLbjtM+c/1rkDBuC3JCqXu6K3a5Bg2APeDsDdvirdnohK6G+iqtT4sZfOaYGti+
sPNoj6IcA9em7tqVFgaWAee3G0pQmxyINi3p66vgWgrcdTf8PskUrYdKC1Z/2rmdw5b9DY09xQSh
YMy6UrUq6S3UnScwrzDQJkECiLQOYFDSKkLcGw43kC6ES2zITlEyr+A94umeswz6Hi1JTcYOcbzh
W9yr3WOl+FVPBaVgkDijEH1fEosvLU7lVDnE98PcqRKr5LndnWZJkDciWOK45uvmSPAYH+XHX+QU
ijMm5a7CdoR1M4f/7w3CKpiKq9m6kgZ9hMH3+m99+VsPo7ujdwE9/5feRndHqGEGXpiv+E+/Pk4+
ba+lqbQjMElxGGZCMYkCsYDdClrHbnG6TTb+eFl3EWvQuAysdJ25X8q62RwNqjDrp64AhEltKMvr
Epyn550qunc4IVlTxAZJiZhgr8uu4992VfFhY9UqchPLXq4ytIDeRvciOkLQ2gKURKvnJAHQ77zd
y+EHG1GQZiVCP2A+uWLDOsMeXmg6HEmdaty02ws5Y5D2OQPtzvZSOKVXCHCyk8erH+e/uK2hfgFr
yn3zvuqBK9yS5xYaK0ngjEBxfD5k1wouig7LWbMTaIHrI6cU8hw2lQ+kJCdsL5PdUqbIgDVuUi9a
rHuiT7ZFsNNACqQvQza4wCYrDTRLpaQbsdWRkbJaZncuhBxWxSo7Pg2syYN/6UOa/t4yccFmoQUI
7ExUj5mzev9Z0qRBak9v0zgrCGvSgR2fC8FyHkf4s2Q/HyVoscERqKB9LSfBl487OnkZBgKuqN2i
3baC7Qc6EMTjEX1tuXhdGweD/QnCwCr650Q1qCgPwXiTzjhYgVFPXMw+fn3iNFnJKkCUqblOFz94
A3zGHCkzk8DNlEPRXY13hYRwqMMFSnYJPP+jKqFJwxWWGJ8Jx907OOUQusqXmebtXft6etKx65/h
sVKE1qi+99GTtHObEoZQ0xVrfrOrwKDY1OpkCjCsQYCES3lZ3EURbp8Fc3uLGv1DqY86waSvlNt7
1JVS4X6QWmyZw4pFZQx/6DZZyzUNJBZbHVagLFmMmr1lqLrziQLaUSGzfcpvmviU2dwZNhrlhCly
k5C9zoPo1e1xRvRjQS7jNtMgl6s+WHUt6nJFbl8oR/tN57zdGSHGVDSb6xTOMOMIbJrA3BHchBtg
B7QlV4bfMGp0RFsxxQPHMXnUzXFq+4ES3ogmNExByjNagnUOMT2t1YitaI90VAvGYSUJI3AiaULf
JtaXDSwFdlpEZ3HUvm+mV8/r+KtU6RcMaq8xkQF1N/r29xwYCeMEKfZjvPpl1eeiVkMuDTKsMhSt
LsC+5AbkU6yrPFi4LA7JNmSBPxS8kOEI7VIYBKmhNQcvxURorCw02oRwlyu7ECCqJdWb7760XcVV
M4z4QycWkejoTswLmFibEDqJfas1aaES5i7/lCkOKyldKKjmsYLuSl8FOyQFI1aMkMw8KYX/EMb4
JtAjkXCWLbGySWjjop0YvoRl9D+qKon2FTc7qZblQ3wx4mvLg0UA0zZQfcXST0wbd8X7V+Yqrbr/
s1xE4vW29Nx0pRnfq28wblRMd/FIwVnPYd2GnJg1g9l4AdcwVV3k1xXEoLQD34fjxzSsNuNSDEW3
TyRBMpRHUhp/5F0W7+zQhvCdwS9EhABcupwR/NqmjlaM658GcDxd+XIHJAGGX+xX/cf9Bf6XlsCn
NLbKRNu2So2BTjsiLCNuppxDj+078lkPph+K7U3ivSr31uUNNVpd2M7O13jG+L1jbR0YA0XRQTLK
lnTO+8iTFknJXTKBrXyAG5C3lfcfxcn0rqzxIvyKjRJ3h/LlxP0kcEYMlVVTl8/PX+Z1uVlwFap4
EveORj1QBq4d74eCGnm0OmFjdNCJK5HzcixQlGy4dNFzCnA1LkDDgUFN9JqCk0lyI1ugvNvxiU3S
WPHHSwypqO0njcySww4TsVn3ZHDmEZf2b/n9SoYyR4Dx0dwM78fMEOORqDsn8dNxYhlBn3Sxetjl
BugIUH6UEGP8qVxsJf2hYnpoUsQbGye5+h4LQVad+ytZJ0Qgy08UQlgAwu0CUbiJHB4QTvFOAYQc
kyZ9X5ppyEYzxjM5n4SFXBYgjqWdhjkZP6ZQrN3dvhsZIOLWfmwErx6/Miv/8/26OhiSR4bFu4yB
uddPjVeCemZHUQt1J97pd1GcuOXIIbisVuTC4bDWJTBYKKjoSxN6RcQaExdzsuQBsPkvC30H2zLb
gOW3bVo5FSonRlldKQj8kRUii+VrbL+i4p4gJVsTvR8JjQEhQcWmwmioBzFrdrCn7kOMoqHCOcnO
SDg1Vg32jMXiH661dNKR/RfXWpfGtm0QyuSdWJjWij6OIlnsOxi+d9BxFiqD07dnIrnoTt3Aa4TK
CG9955jg5w4VnbtZBNqN9y1tF4+cP/k9mAbIqDqekW+QaH65qbLALg+Thnm5sg/8XxMbG4yD0S2B
KnZnXFK4TjisrhkeDYR89DtAxP3i1oVr4UNBOnJX3cTluCLiea3uBRdhPM5G9JkDoj+F4WJGLsou
8zrAjQrRAy+S+LP1iIuhleOrnwJI7Kit1uCmvpuAOSvos4aEtE0mEy5xne9+XUUa3ms+qBmQWsob
q6Gq+5ImXzEoiHPMVW/gXrIRhDomx+soQDxNABamltxJ0bzVgSwL22i+PQI2YLr6PhVTACyc6WPM
B7re2sJfSy/aljcpHBJbaDlfdngVkzIyt/2fbbgEQmsaWGtdhJaLvh8gFr+DByasnDX7DcMBNPFS
7Pp+eZXU3EQ7hc7x7Z0xge2XL/C1RIZx29FXzEYeD1H7U1zOu7dyNf/J+Cm8kRi46+VI0o5FSj7j
Jq26b8T7ssJIKpItlRpZW8rFcMAJlYtoTKMqzKgYTE2z/BjhvlhuQMubrNa/aQ3LSVtQD1yxl2Ty
eG7VYQlctLywSJVKI5Qp3rprpAifgNNG6FsPoyFqtoPcW/ad4mg+cis5JF2+LUr1x+dYUXrSELwH
JMHnVf8FTFcxz5jdRu1lnunzRZqU9BbK1cXF9TyVWBueIf7XNj2NMdvVAvHdmv9LrYEPGmoNoZqc
BCFHPg6yqH5KinKjHRzFKpu6k7Cnl/DXK6ZvJohvPu/cgtRx66D8KBKJN12bH8arzGTMxSMPkm6u
9AGOxfMUwl5KiEHG+kPlT0FvHZMwROfxxTx61k3YEksdylctYN5tLlWAfdNta6DQc3qltv+T53Cs
Pa8HgzLbIpcir0HAMuDwCEOKP0KBdHfyg3bGn8rb04icyhf7NTCWihdUPnGTGVZ2NXqOlh9m6yZ/
u85SDAeMkqzEkWyoxRGEjdMYFdlhEmm0YlRHwbdTDSPZ41seP05BMHwkdRdG8T1GILxlG8oHPR9S
R9sjPJQcP9OnfK/jmrknF+mO26N9rFK29b1GjaYgwFWO1gN33INp28RRoj897JU/ZtLctbU0r/P/
+4VaMj5dym3mBIRP0r2/9DZbk9zxvjceGC+r6VknahLUoFkdPEdC7MShgP387qQQ27zQiOnaotKu
FbfXY/jpCw6rMhGxMAQnuUYgtWeeHtqULf4+bhxXEuq0hmJL1r3ZFYYiFfkz6Mh1vqDdhwYphYg/
fybugAHS0XqUw15BI4YihHsfgL0HoCjnWMG/o+PCWaUOprfmL1rvjyKAlVsHCzLICwDQJT9fDSvz
kOQ0gKAMbNtcCndlgWBe3KdamCFEdprCneco5unFAaiGwp6cPoW9wUKKNxd6r9LzAMvAvAz/7dtB
+K9Q2xaFP9ic+A8hsKzQ0fUBQ8KWNHHiFA2Tyv6PjSyUH3HFP/agUFNHZ5dgs01EGVSuX8tvR9Ff
GxeZhmq2vrlpuZk566IHj8NDx4TcE+UDh87L3Q2RCw6KTp+2/gNE9yfTdC4LoiK+8AMWWPwYJOjO
XkFix1NdvkH3UyRDrCt/k8TtqFFR4rQ57E5jKFCmdafH0Bo3yyQbClmn7DuzvHLRgnGe67i1nQ65
ej3Y+A9G4pI+kIdmaig95id21gAQ+V7mHavvQMjyGAEYjsb/e0POiT5o/mCr7hDjyez3mLU8EeJG
9OCDwUU1j9qo5D31V+Hf9lSQxoRv0/6ki/rsN178/i5hMWwEgZKUCsFXhe+8gm3QSJpZUZaN7AIS
XRUzSHeKXaDj3gtQSmN+6Zgk8H1yYY1aoPK76iKtXpvE2KrAqo4xAHtcCRDRgEiJ3QL9KPumAzjl
9nvmB4hnBXwWOd5HEgnKvRFslasoJlNM0OQRe2fQHCDvvh/L2FOP2iX4WBbs69gSsLXXznvwQ5Mh
U7KuA1wmtDqK67EMe7HYJTrT68pGNrD0Mtq487DR0uepYtttVsdpLI7Qu8WNZwoJSf/RztBpPlW6
o2kUAVWn6VlIGskplZn6O+H21NGh45bD46T1u9GqZJUCJ4LmdHVkf8CpN2D535VftvPKWhfaWGqy
aXKSJJ9zbNvI25gdSnkOJ6wvOZSzftA1U6Sh5T+GtoZD737Ycdy9qW5fGKrE6AebKtKLGArqc1zt
BYY8hr8SIc0TwvR3F99NtHUkG4gwAa3luPu8nq5npZwZrPnJ177xd8yDYJT+w8umAAUb46p7pyft
qmi+pOGxznqyzhzErd34+B8YXCwh9eAXlOrEMlsl4dhd4BKXyWXWD+Dc9V/sqBLve7E4AY6PGluI
iVwBv/MkBsj/+go7atpcL0UOGTO3xLJpBdc6TynrsgdALWc8ic+gkjzkf9FpNuGLDjeCNck8Ry+N
nUyJGWyeHI6hNMJ/x7FRDkxgoyKs0PPfnOfy0SKe1ycFWFtTX80KH/7eq82CEAfb1mSKK1PGvlJi
w9HogKGrLGUATgsZOGPgz0WowKsOLgRckoQKfCUdaKT2HR72qTw8Jq/bIZh5bpjnwf7ZT77COOFN
ZDmI32GSt8FebF0782fYZhKd3OBWr+zBzlU2VlCvHtML1oFM8/ODLK6wgs4Cp3Nfp5b+0jNGVJxc
w6UAxBjHY42O1sWsgLiK7CzB+xbR8Yro7w6MD55hnpPdqu4aM8DYfd2ON90Nyr49q6MHtsoDBLIV
x1nVJO8gPRYpimWCPDW3sR2bqmXN260HfnKHJnf9gWXAJogFdQ0MNT+F76fyZZnapUYv4yDpFY21
S3M6YPKkpj5xV5O0SQDfWtc0DYlemOoI3NxSwUJv/is/jX7nkGksozze9JopclYUjvhslgOImZ3S
ukYe4v3HC0d/Wr6zcnnbypvLVliybLXOAjKhXH5MqAzY+Iq/ayltlBbn/6pbDkFEyYtxsLZ7TQZ2
tol0Rr34FjO3e8GFE89B9XYFBbUJDPSvSaZIIVjyl5L6jCQvWHXWXt7AaeIdz9PmTuaPKuwBpZM7
nIg1uUt1tvE3nJOcOnV3m7Z0glPLevEmNkgQ6yOGmnci3t8sOrjwAQJMSYDcaVcBBrSrg0PB5ZJ2
Df5RU2glGLKlPdmf+z4kOZsm5/2qjj16nc18zl7chREhDe/9DhpDoR48KR1TLWwdmkM0mSUfQr19
AzvweDmFYkvb59Ip3IewiEk/c0AC8pkC7C7QzxVG4SVC4nHeOy6NSBpmBAs+Q0eknVnHKNCP01Mv
Mhx6DrZmm/hTa5aW4/2JehRCHEus3OdMEJQT3neM+Uq9Nd9UDgVB8BDCcXSv+O0MbDdPJ1pHp2z/
prAogGdW4caZIKCYLoglhaxcvb8E/g+w0KjqIpGsKaUBMzj4cCwvo+hPYPBfjnjuMw2qQeYd/a9z
EtmcKB2P4g0+sLPEMyYxD01pw/Onx/ornb+rq9hYUFdkfk+Mlv0JKs3P1o5iLQHAVQbZS6vNWf6E
uQ2GGFtdjtK3o9AeMnCVhW/8knU1P1SSOYxH4PsblJe4iOT+oWNd6kQomdn9IycuR9qlwHVAsIKo
EYlKmjaiL/8dvGFatkmpY2jTJbnzXXraCnrITXDQHSivw12uQyOByNX3s3uS+UnFlnir1oQddTS+
aWsu5866jL6xIZ4W1Fh7B6PV2kYEuH6t7evjiAY2ukSlZq+Jkf+Pe6UgCVMoJXomeJ9itK/glB1R
TqY/TZVukgCuPRXVAcr94oAprYvI+azVD+L/bT189gWpSa8GcfXOJDAWBVstplYRI5L3I3NerNLA
6T4AujoGgCIylM1MmSALTpmSAcStVyXUDFyMhqiuo3RwY+0qeZEvIzr68HI2PQZ+bxjbR3tGfEBk
AH68Sf2EmHAoQ3TXuK8SUF2Kz8tVdKNHGHOHx7jOZUFYby4kBigjm6yTZ/y5suRi8DQVRgnjbhHP
K23rmQ0k0G4+9WWXDB+3P2V3khy1liIUeC//M1c+kjdiKHWhuhStOgJ7mXMDdk2yQdchRXWXY1XP
EaSW7esYFjrG65gFkuEjbFVXd5BnVgLIUr6df8P+xuzb0Mfga0+80RWF6KQSdyuUWLS4R1J5lOX/
sgqPwd/9tuXMaj7VRNTICrsYVIeGejlHTZjF7mR/f47U9OKeeJDlmlfaLXoMbLRM4bs8XOGWiMb0
XoyRz6Xr92n7iXG9XC6pqNqpi04tSQR13VIvu3LXDNFvnX58PU04vg+eODHpNgofdqDi/yh+8z9e
Ki7Qr/yRLjMInIFPq5FSP+p/C/LN5lbpxd5KiMoHCUFIQfO6tFt2gZ9q4KWntQ3KSRRNqJk/CZ9H
n2d29PQLXGpoKs0UyByf2VPxtQDte8WFu67SWJiKgJFm3O/XrwRbaDAsnNrKv6DEKjUOIWQv7jxr
6NnVKBv1Cvncrrf8DomR8NWtl/5YO7E8m1dBJz1p0/4+gh5nq7SWXjZQUx2qD99Y6TmaQGH2Jh01
gznSZVjiQRyTT7B78cGSh4PWYlNeutfz2y+h3682eaaxmSji0y8l2LBD1vlR3A/rgcvTAOLq6dfp
LSeRyEngLg5MV4JXPX9B2HLjvqtYtDWt3sOO3pA/8I1ryXKzlWJGNxgdQHk/C1U/oEpcUPi5RZpB
SEbMXAkIvcx0xPmR1Mvr5sgnoPizDscqApL0TcHeqiWzmXuQw7oHe9DHNHfuBCLjlauTsAtnZlxl
o77vjPvaWPY/BccpHq4+8PcoDQlg6wgAbRF7K0lZ2fzCCt+ozNnpRxLpinM6MSifS3BsN+xjVpTR
Jiw0ihNMXHmHYtCHcMThU51SVBcssNOmFIOvbFpLFN/UyTPa05spLDlOMo+okAUkmL1q2QM1Xgw1
x7Qt4FTFdXGlIeYN7XxaSu/HhmsspIVfHX+rz1TCv7y7wd4K+vaousOyDc/sw7Uld9k2sx3RB80K
wnv0FcQc4R+bP/2WWoA4KzKxxQ9+diaP4DNe3v6cLzhqyXJkuAtnqmRi/ExVhao2HywgX6g0SEqO
oEX3ifkI7xoWO01GExE7QyObrvvIYH71MBabEfRU9wi79SbyzlCB9NO24abiuz4bqYhl/oTOx4hv
xcnpyS8pWZP8+gf4QrwgoM7KGtE6zkQ3dTQhkqWTkercaYMQwn2d0DQI1a3tIFjqaHqbYzA9P7/a
NH5sSykrohuK6rfZLF73/WeKvGlleRl+E8CGc+8lFykfC6NzWafWDZopCkXkxncHjN2dbJcG0p/B
q93C4BfGxvcx885ieUSk0OieDImj/naAi4Q6Gt+u9GlTdjOt3lE0xqSRHq4G4z4caQiVNfRTgvar
wRJT8xwcM5tuMlWE+X5XThWD88wNDSEJMgLcJv+WbalabfjiIf9YWZOXv+ETRFSntrr9B8zgCDui
8i2Hw9HOF+sQOojtPAIlYS0jfLpJXsQd38DTcq8TEfhP1M1xIgCpSt41WyrqhHMDEson6jQ5m0TW
3y5uuq/vx8p72rGEzrgpQ+KZ9yJ0d7QmTbWLRePfUR2WQd1LUST9wXSBHCCzroQ5n7b9BhFixh9j
Xoke2/Z111lFGeC8hMQW5+MwtoPl80vmt2GfYI8dx1/XVC/JDRyNlfHiA1zucmuCJDnNdeIFcrg6
X00TvRXMTTrgDyUnugq+qt8YJsoh2vCjadISSFAO0rPYkrgQfTaq8+HlcwCWehnGBrv4sRm6LGKe
OdkRb1bNqRhUdhF2jiC9m+MLXcLMO9gxV1TkQIV4GyFjuLWAPAeb5qUormww95l8YAXloMasq5xo
R8VjuQfEGSmFKBRo/wGqFhm51tZw3t77gXqVBp9nRnFwoJuJYgzRo7FsS7I0xk1Ls2GtMHW/Xp1I
rn24n9HY0gyWSUhi8YoV8m+LAJrUHoyjGZ6dHL2gSV2CWNnj9/R7+0YZ//cgNj5UcPt2sh5PfAMt
Mq6J8Vi1MOla7+c3ls7dZTEQowoPZNu8xa0lCd5gdlpMuFMT3b3s5N59QyV7EpNQLeFdV4/h+0XH
sXWvAoL/tKZVB58esZ/Ibf4/fcpPA7j8kr9Fm3840akFJK2IMjV6OiW+LDwvfqYy4/aW6pSSIPz2
AyaAIzxampdGAQq5c8/yN4z8cic3jrKNJBCndiRTqpasCBCQ+9OYD0Oh0E8lYoPnZiGsVKEFp45h
gQLVmQlRLf3sS72A9lEFPq5qNojK//zOUPDPAYvyawzjepKMOqeU1X38GIubrAFz7LeHgPShvuYm
INLVeunAidXLZzRBb3qDbGIkGL3KCySvjyUz+6y8MJooXUlDd4EQHhsL1LN39EO/nUfipyYOPJE2
2ugxZ00gxs07F5WYF+mRb3ai0/qwoOchBVuRyqdkDXHo+yrutHpx0pJZ50HdQfPDTnXVRuZxYjMF
U7uhIyXyTGQrkl9KH1TgzGz2ZoKB3y5oxHKeLn5rrfYBfrIEdFVUPtGa5rJU8SdAV3J0VzM5wUCt
aawl/ehqPieWnxfj4lzwL5HjHf7C6kcHAy1jc8I2fEkVQ2MWUQC4DHWsWVXSvb85tcAFnybxuEKK
cPcBVL5FSoaeXj638MC20kp/42WRyuzCmUwre1X3JMtDoScWfCo+uoV2AAzL1WlhVulCt/7TBrZQ
YMIz1zQNAE+v2UaJCgdrIgr56tiEnBYhe61JlV9HOcnuRj3Iwc4P1wIDxgWG5wfDNRIt31oCZ+Uu
s6JG7v0Rz7rNh/pwKve0Vxmvzkv48xubeXdfOKA2GVjQsfugC6D1ub87Hg6obYLZ3pqSzMml1fOT
1tSfKbw9s5PZa304C1TdwbAy/QsCgTLVSDCDMR2G3uBYMj/SPN7TBPkqhhY/ewfqS00F4MsHz7S4
girctfABFxVe1V9c5C6OdYkmxG8zKEIEWqvMo2phVnwceanzR6t/jXfZw9noY4LBgDRKJQYt11CO
qCcgIYWsknagpirFNdDZj+ySbTYTDa0UcyezN5aVfhSUziZG5QONwoA/bDRJOC0Jm8UNrITCaNNP
2Xz55swdHecoLCp6rqTl/zerL8AN6pa0p+PU7s0D5XTK1oEkO6adTa3I3rD/ovrdAY0+2sxnPh6F
iTVlzW1oixN1J6bRF0qBO0MlNAOZvyVpnDgA6mmeUItluvcp9CO5bMAZTd2VRvGjsyuJyZaB306v
Wxd8sE2xsw5MVrkR90oXhRHl5xu8X+WCGSvsTLt/EYPw2ePZCpIzV6+gRzV15+c/0LmLZP9KDJSW
LhdbUk99U2W/dgn/G9MbxPGAxr7t74B+zpS/vcDY0gTXa1QxrSHp3dzf2l6fVeBHnSJXhssvmbJO
6eaNtr8PcMVkxN0RJDCi3K5F4T0WhwrqW/uIJtSZekTYd2E+tHqZJObg+rxKXIwXF0TsBSRC+NAE
I71sLT1Cz+O9m0G4uC1wS5Tq0mxoBWs4ETY+WIiAceiOJvzMiVH+K/b83oK4DM7JJWjZ+4f5qDME
OVq2EuKAQ5C3DD7+R8JNQ5CtzuHPPWdZxZDJA/CJqvC45HGGVIywJWOjGyOZHwfstZB+W6fyPWM1
4CZB0Ca2isP6ysc0ud6YUHsCRYvjxh6xbbFygwW5AWA4P4v4Cyba3rPWTcEB7/JuD/H5xcpt9HVZ
gxpgA5KTK6YUHZyICQLxUW9seVqimGhQHja0vqN0G2YbGoY4fmf5aD/8tVqsKTfHZatNeXFJSdRA
obOEMAoROyEtVNajy2wlmKd8D3uCkgKpteqsgBy80h0+4JdFyVyGCVD+MpkPY8VoGeVM766WTo7p
iSFTfMRvaZLilJElv8ZEO5eLR8pR2oj3JF5S77bt7USrI9xN3gC3d8iVasdMBSYW06PV9Uq/1KYP
SVhikEgmWDXIg35ZLhJassRge4T6rFN4KSA3Vlp3L4bCtNstzekGB6mu2JxK6v5+qBMc3RpOCvYS
FzbayHuPtMitveBp54TJGMZtjmPHZfK9u7fT7jMWy3gUO6hb3OyxFno/Fua8YDb7VQZbEWjbGoz2
7YPPu9B1ibg/rzIETukEiDci4vmfHnwPYRxwsvrIag+7Gap0h9L0GTHzxsGfa7FXkEg9aVEP2kZd
47R78Snb2J9YlGF7Nst5urMoGHHRswktmQ9WQ2CJICIPuMpnoi7kQ7g0dTM3nB5K6WBPOtnKy3Uc
iL3cAMVyVjbENHhEp7qRuInCV6bvLeyMd3l9VC+AJJgbcmPC/U/bPrIBQCmMqvftjK01qhfz0hKw
oS1Bo6Tg3G26aXoJtv/cJraEUctYDIQsdHz2+Wi8la4VgJc3AUmgCKMQ0A46/seE6OO6sh5n2IFr
e+l1AAeethkz4tAS9oXMTABwoSkOSWKH3Jw/J4/Ye02vabFmeX/grfzuWqTml3Wft5sWkz7trSn/
PRJQ/0SKeZJ5ZrXq9xanPIyYxKuwbT3smVU1SxNQwy4GSyQ3nIeegzaLI4rsf6vrf7anRcY1K95+
Zo9N6TW8OL1OPd0bK/j8TthlFj0wkTAy7FTd+e5IXKyFu6KQ18QFNhfJDUY4s8ESkc1O/2dXUmoR
VAieO35JrIWd3Ouuv28YdQaARxRzprkzNzSU/7r8o3OqBZjjRcESeBCz3DtuUwcSNd9LNcTFLpMB
eVGxBDKASE/YvsiM76p+CihF3Ygzj+hkfdSWHD87b/X0QZJu+Epko149lt5pEGlkLquKcsIORsym
RsIL8zWTSIjGwEEzqb3paUfyGCabGgFV0c/vOY013mIByApGFlABM8ZyH/BVb5MlNf8z+uPYKCgK
WfGCx2TVmzL/TZEn8WGZM38//nvpYD6IVJ4vqPlHCFx6HcLFsKy62m0xaL7h1HhMrNkoZgNwt8+I
ZX6hnAbbyVOxxV6tm3nR6pvNYhdi15IghQButVXUfO2zetQPdhU4uUNuqatmsTA7jdpEZnsUq0Px
NDxtKcgfiTXQESq0i3MYbcs/P/vydKJARb6kKGJLrBDHKtAtW2jvOeSJsHnib301ViS+3uQTONjz
qpDqTRRQoH+r0hLqXuumqGryntNpe7/8Hq9REnKDHUXlPn6+3OY+khSghPgJLP10/We/QAZWoHYG
5qoLLxuwAkl23Yw8FH+m013GQ1k0ckhfwGIWv2TG3DNaL1++ACicThH3JNtrYsjnzLhwEd/E0Psy
VzLZUka2khMCFDNR6iObvcdw5KEXj4YFSHCK8uEN+6rGgKan8ifOc5PCGe6LKswVDVNkZjNW1r0Y
x6WzKIz+Rj9zWFHtScvXhT0fFDh8q1+bqytqgkTgM9qBGDcob8sDmzVuF0Q/GNRqbIatRz+hOxqb
F65LxIhH4Dk3tb+s3vvAVDRl6SS0/SQx+5Q4z5/mxGsSeikEwpDPnZFzHkBGlnehBuawfMVNtFPs
VWPb9qN2wZ48fgOksmcPI3R0Thzq3jO/BcUY1iJjbdGFIQhkhwopteASKOWvhF/Ip8I5EQz3CW9m
AlicXlyizb3mq18YXhhJ/ytuBEFLEc05qw0hPYmurTKPoHWSOYMqGv97oYoesaNjKiAk1VCHgH14
alMUTveo+i2EvNd7MqQCfAv4yFOP+q8VgmE2bo8l7CUb5MfPN4yjRHL6jGXrVUFlrfqebUucm9yM
pu2jCWTMmb0WRh6PC1dRQAWyZebdNr76NhmXlhj74c9Mdt2/qm95FiIGKJs5MjgMLrwda8QSIwkx
Zx75TgL7mEj0qZwRAl8mhQzLsDGYCx1+vWDVFxSXHUW2y1zTHLl/bbRgbt9V2osptCA792ZvbRrl
HTbxwCwibcV/6ZS7n13SspLh1Bgqskj/AMyRJPo4jPGoXGde2Ii/3Z8Gn9xNRd/cEMykkOZkqLjn
YZR4Z/lvhoa/e1YR9d12JfCZyyMZ6obrOL337KOlflg2J/S31NMTkHWFdLolJHmb+CfpJtGL8xCy
eXoOqPA7ij2hUJ4/G8UOmIb0yRfyatWnPsak6TeabPRuagKU3xbJV0jeYyFiiJa2UyELPpQ8Npf+
CC7Fe0L6WzgehGzo4M4CSRvcIOnE3+dbf1IdX3sSETNtvVpD2/Pp+g+iwRoZV2Ya4g3SUAVnCFCp
xlMSL0+lDZNLWsFeb8X6F21NeRVyqgNnigSw01suZaRwDhuK+Y4+7EzuH5KHZptTcf01iahfFyhQ
AgCh2RNSvBhlBps4P1y3Rfj+pAf8eF/eScCxRKvGH2oUp7GaN/x59NAsW4H1vGkBhnsSufS4vghC
U+t3eJLTN/sPqedq6E2ZoLbiqAUEdT0RMi0AKaaR2N4tU7ImcyRkz+LHINwGGdaFTRMEC0gCgLNj
8ks3z67UZsBe+wW1qgwk49Fb5YCjAVV2e3zh5FC8eKyUW8tV3yrIX9g4GSi0n1a4W3QwM0I5JIRM
VbQjAwGtdFrRVAeI9RIvNir0EeiyNvN3pnnv3NMZU9XVNdqTD6BmBrHMj64CrJu/4muWWtRNaVzA
ckae+BB2d71YhbMtilA4qTuY6QLMIj7BfnTMTvsgSBD3FhApN/YIiqfImY+sEV24NJI26IEX08ud
28uEapDsYfcJkT0sIrKnrFMNy9COL3Nit/AbPRgC7dKQ5xFthYCRM3Fvq2HulPZbfKdz4Iip3k+y
9NT+WhlrK0EZJmI/CqV6e6pDHlJxDsFlV6sHbA4X7lNGilHQFlHqHdukHs2+K317DF/lurOd6b3P
K3gspO59fXZJUsLkCCYbWLfaiOH2vPfA8sFKUK9aCwuHXiWZ8/wieDHIYvb7+UVGxiSUhAdGCP70
HZ4O8TqecvhOxuKVpX8/2G5068VDxAlfv3R42ZyufSzwvgyryB9IppnSfWASnTf0VS2uSfU/RLF2
i5DzxHBBziKs2tmoUAYnPCzaQ21Xld/8qtT/5YSDk2MffSrPUHmThf30k4Z/bPirgOjKMkHQ0Xyx
gwsBertB5Z1oETHQuCe6Y4FNOI7ZDcc2iYqc52CjuiTca41DHusdmBjACcKSn3wh7KogF6MbP4WF
U6d8NHlvJrHCdxI8HMsrNakj2YrW8BV1oqMoL+jFSBWHlBslndnxG2zP+U9BReCrruYsq1Q2kfEE
dLIRo2pPG0jP4kbSdZIiDoTq5/h1k+1ndw7tBCAxXudzsFuCcKe1VGw6sIHm5Njr4zhfcuJVkgsR
KyBBvjU/p+6GA17lEp1NH8nNLdZE/+pS1mmCEiBjFL1D3zgXV7PuZ2lWrd2+lzLvUaa6kU8bsXNE
cAt8//1iLO+UsAug/uJvo9ERNa/PuPvlwFtocrX4s/Wk44Zy3u9BenNQScsWMft3jCrkN77CykTl
pH2CgzHMoJmJAfqzs4xcwLjpsvhlzxSTg/JANIEb6nU4uuBdK1FOpuxwvun+LEHqewccNMIcAtts
P1gbtXAj0qUtkcbPjSkV6KA6cAvOGRVedJWWnU4YhqG8zSeOZ7JGI7nAiJjR15/0W4fv1nyrBuEz
+gksQ8jEqwaYS1XanOU8n7/N/5NLiK1FpfwqDrWeHOYDQO0u5bF5pLIfu+qoEyuzwOImPy0UcS2z
RChxCIdeGbIO5aFu0R3LZ1g9xdEjG/EsW5VxU4GDbmH2k7s0uPoRzheMUl6SpmTP6tmlib/CFwgW
b1uAWOfuVm/XOa4rhxXJxlBuHoe/5M9dcoaOszLhlisgeJvHkH88+5W+Weel4fM5O63tAGFP1C9t
cqhJRuDm/i3SzdoAS8T44GpKVBEbD+GRmLFVwq5knNbGUztf9WUjs8iDsSMglIgnASeLPFnhRllY
J2yKS48ZeY06iGCiXy3TphK27p5qMxACrVzxtpUeI+Y4PxJ9FVNBW7LnXHxng367FWRJ5DGvfe5d
PaZ/495EOwnHlHhoHNKHmcVFWbGZTycx7cnLg0+F20z3JTxeYhj7sXvYTh+c7yb1VsMwvSS3O8CB
ND1t/vswvBw0yAYoj+Wg8gOYFgU3m3v3EcroBpM5rj7z1z/pnLd2+M5zxvz3AgGS18GFcyDjsS5I
bmUH7RLPnkC42N4TrNTEgKZGOr5jIEGdgcBXIB8vBk4CFCT9mtEvCe5lwTFRnJUgzpNl07i6+mV7
uyrrwHiASfFTkLaAgK2Eo3XYgEbeme3fVcNNu4M+XZYCqyqZ7z/aohOCO4vdj2AUGbRbIWKqL/yS
kFI6rIthXCC0gYOBgTwwCACBIn+BzHoYaX2+52g5njuRz613+E2drUBRT8WF2YopGoyn/+SPLZeT
cpyVQJfNpllEidinYAF0UJjlL9LwDajNIadX/263L6CHCNAyCs2V8zaizqnKsxyKXeSh4DnA+Ecl
tLu2q1xAzHBAKLUKCXjEuqexyLvcqlGgsruTS1zDZOyRkH8H+F4qyNMwkWp+ZibEi5LFFgj9VuR3
LuKx5absUrjATLuJnFh4mWVUqLvhgGKvPcbnmvbX7DAoNkAnMQmLV6ETNli/5ckmvEkj/bXHKYU6
22AFl3cR3vcY5TsJew/WbWdWJ+rxFRJNk800AQrzP6d5qDS27VPTd1NaXw/kQC+OeXSYOBkDmsGz
66nKm/F5YCo+U1fRtFvxFBc5hCuo+wPqk6ogkGCv6o2JWqDLHHYPZRzokXhqo/5Bktfe11kTQJMP
Z7BK2LkMW4gtzIeCT3BsDg6V8hCHncBkXAbfQav3siHa579yiGMoF3GpZyu2/r5eVegg5UlXoP4B
34GVDPO4KCdXCvc5o755cvwdHyGm6TJnYPOSCA9pTr8wM3je11xa/x7ESPxSfyHdfVxuGKxi10gs
34rqJaoS1ovTjEgKP56wmPCaneqTl0tihA5/HLKFd9wAaoVZCnZJyVKmanVdnhoioAUzUzfWZY7d
sTfpTVctUrEMl5fHu4eBire8tkv8YxtlQDYJdlBcT5yjT5J6tPwnHc0eLlA5fvYUpla8MBKZZbLo
gsrTCyxNEFg5h/sbh3xUt1PSIR2l5wcaDidmDU/sWgdYQLM6y79fYUPfaHKuih6cxJODanynrXIG
UH9/rp6Dt03RQ7IXdyVcKyzvsw3rhZzxp5SX8uqcil8rVgQBd7S5MYwXxjBZt+E9jCzqjqiRy7dg
b0GwRXFD0XsYBSI2IEH2Yj1tZoEr09mT3cSg553R0ZVk1IgdpPs5WdYuDzvKL0TkyoYPgweerCvB
Ki5PIgJ8h5iSzASwFsJ1uwfC46S0g2z54AVOzPTqVZG7cqKX95l07ej9bt3Mqma/Z9mDTsg7HN9O
ain66Lu0tV6eivhhnOXqPFpcjCWjgJ9zHz4AFrHOlVs8RT7152LM1nAqrG7gfkm9Arf7b927/wSq
PnKYsYsWGlumkaXUZylpOtVl9VCqoLdgi1hRfzhZ6edixlE5vyXsSJL6h+C33Tm3GWWIIn4kUapA
lBbKhfXGZ50k6RkUWhrrAK5Fytst89gHm62YPs00EHh9LDw55ZVpQXwgypVqEFkJoGjEnhPhryFM
6S6c9/sNO1f0E5ugZ58AEDjnT3XR5R1sk5d76nyIPUxQAg38eZ4ew7NNoepBtYPS/7o8hCfpcsia
Jkv9op2td66dj0PQS8fadfwlaI9m2mv+o2NTa8Ve+yZiUWMFjRwvo8BYVICuSKlQCX2D3tXcA5dm
2XLWVnSVLmPQY/mESLlYw0Lp8lXkKoixScryXf2FWKZ7w6w45Q+FgMVgCccirGIajRPXV9g6M3US
KleAY+p6IBO2JiMVwHCfiJGPEgZm673peGTig+MoNO035DK1PnVCHUU9QjJMHZ+P7OfIP3ssMyEz
kwkKF/trRKGynR1YDSTwPJ02CvAkjRR3ex48cMQJz1jzrWp1rCpfd9IRPoaV69znIEoaYX0acAW/
/aBdXKGmMUMN3UK9a6HuUVrCpnybZZ9QXqsCyereHCf5j3nkThTGqm/c2fIZF9N9I+gAR0nC8HTR
dRzuLHCPyzGdSNK4LLLs8XV1VqkCB5HRb9WxaM5AiLeKFbvaLcbbPFY/L8UpB+oqcE/FLMZxyX5U
xTmZD4YjWziSzs2xWsfbUzmX19pvqE3ldJNL9eEF41mt7m/VsYogjjoFVtOSxz84+ItMdrCLOPCC
SL7j2WoMToFPIzOZIMUrMmuTiCPyfxXGQyoPtns6DsmABULlcB6KdYd3ttXPoK1tGr5h0S63sJsZ
VTln0mnjfcYhjY1dALClmDyyZz6gTSorVtRlMbD/DKG58HnYx1JDpdV4KqfgleVabtyJVMctBgNJ
EWlq5NW7TGojO8Z0WskWkOKSShl5ZnDqlXY+ITOf4qVye474i9eBwFy2tCeWnAs6u7PaSaNBsvN/
YbZzbHsZ32WC8LNfLwY/P317I0a/iCLAvWRgV6ICGk3aRUZcfM7qa5nv2sdhlZOIVMwim+3Vj89w
l9cd7MTI8N9eR+KnEvjSVvWvUnHBefMCE4ZLKOcFEDk3ZvgtuY1fndu440eBw0frHejiCaGEaSFc
JWOnYzrbyU3Pdm4tHVeNUBTtwmTK7MriE3JgKzCJwUjlBQ82DgbEt43U2uwV/+04aCKmj32t+niX
yMbK2CGIx9wZn4FrrxTsnip6E8x9REID0CNj2zj3MFrpgGqVJOh7P+8pz8wciI6OLOf6e54IuEVt
yNKU0Fod/AeISUozcFc43h03dp0b6HRD539iEdLM+gZH9fUUQPzrHz++4bC04ceDGtSgTemXszN/
ip/hDQpqYwL+QDr0jkGyozoqiMwM+mrEXa/dStSXP3qIq2UlUe8gLplToYjoMrnY9SQaxcGucx28
eZRZ9WsSNOu94F7217uZ0vhEaW186sbV8nRfzPgh4+XcyMolD2gDegbmWX98r8UQmboyMw2Q9uDv
XTgK3DzzsOwI2K4UKqqLl44JaWZ/KIWPjvASEFeKKHM2iCoLv5RbzKmVD3WvXbQuqXyu/9ZX/XIk
KzghJ/6rwjYG6du2TbVxly454Z6E0fOMUJjw/KCDXm9zUBr8bMSE7+HZaC/Fgeh5XMynEqWk+sd2
RiMsyi+qinJ2hSozjgf+v2GoLrrSHQPbKYBbwO+0i7ApDYB0NKPCslhB4Qboc8J4EYcjGUMOjSpi
Kuxd/Z0HdwKW5nwYILY4eJx6HZh7Br76Xl85Im0PI3XgpECE1GCB3Des2see7XwDWKyDhA+ghGU3
DeS1K2eYOsmUk6gTvjaDylagb7F+9/JKTQsMbukSjAodJ65zlLcYCSUZSajw+lcDECrrzX/CHH9d
nzNQzMdZc5UQFgxMxwjeYOTySUroonv9CVYxWCFBR18lw8PnEf7/NpagdAayW533aVNFongArngX
KamXU92qXZWlBwsZXVoaoYa4WsiqgvKOQfJR6I2tN5rjlhKppc/NcrMc5+DYOpVfaIr+2wzuNE0E
ShnG+/z6GGHP5UsolnfB8ilv0GAOWyWMUi3hUNEbx857A6aRqScETYhhzYdhX6vcG1GQKtPgRqbO
ndZh9YHYncxObiAy6IOVXnF/bwk0bTpNjQxinieKm5k5ObSqvanaUjUgXQaTPLhtzbRlt4PT/T+Z
FbLR1BVhP0vjNvwEuu51oMF14PYKsvwWJ5Mos0FhMebVzelRxxJ1pK9jgwY8kOi4C8SgXO6YbJiV
LDUPD9GmA1lFNpSl9H1G/W8aynGiGS+wHL4PTzdM8M2kSQobiN/vXGmopnhLO6Kae7K3fJtwZ9Kt
yFOnEpMsoBNmeBjFSyiMLEGnm3Ning7lU7yLRv9SKBL0gDF5fqq7RcBJcOoPJAn4BZLCWtizfm+d
SsK5V3KaVsTNREWDt9/Z2HJJjE1kn1z/+R7WzNmOm4fBYZpIciiGdnVQvoyf84G+/7hN+R0alBVQ
Fef4uHejnFHQy7GPGGDDoQsMjGFYcgoa7X1TvxB8GKv+xlPuY3ilQnOWlN180cfj3W+XzbXp4DNi
iJQ1OCNHAeDTM6eWs3Pl7C9pv6DwyV1YN+q05MziLbV8CJb7QCiJgBViW3pkMb0DbnpRJjTaehRK
k/c3SAJzSSkNXHi/IgIQUqmtgClOArLBYZCNsZEyjdkQbfLn4wzcV0+JUR/IqA6gWMpBIsk0kvDI
0sCZG3WjBm9tHffDr4G7RkVsDmjJ8JtzGs+E9c3Kq/7eyPtVAryC3xT8bA/0EGC++NaHEBQEvnpQ
1upva2W1DjOelsrsWj1GoS9GbIj7leVtHyaSU4FsVEKXoNj1LVlmisvDHzq9NTCkQ86GpA/StmJw
EA0ecgkDSdEVBFh0elV9HxItle5la2/Cij1gJI7Gtzg3IlgaUlnf53YV7tXblKVS45ek/vN1yWPB
V9S9iXvpj+kSyel/1eASNFiy1Mxccg5GKZzlyHTRE3fQj+KcRzbe1lnC50GvaYPwkXkUQqNtiC/A
qDFAL0XXJ9+wSy2gPqjDPliELyLwBo0gHb7BEsxAfo7H7aeM7+UKGDf0i+gRMNkxyxr1QH66Hcpy
nxum/gKe/PP9CsbAJKRnexZUvTWikc/vPHZJ/ZfkXbFwgsRb8CGGarbd0PRoNKab55sZITbbwZDr
uUuYQuwOkkMPK73HW6Lq12UeSLplemeY2I3TzE3Vyh6jF4zGOejx++Su1MBOG02ywJCw3ChM2IQq
UQYTwjLw/tbrOa/TJosM647JuG6DgBYSJDuOyvmGpa5TIPVCU55eB75YrGpvayZMgCkFXefP8stf
DjAlRsJxDkv98+0gNth77Qm9yzey07LxTihAFcaxL7l7aUm5v0unDhCgYkMyKFVIqQOrkoS4c8fD
2xYE80jWzLwzsE++Cenp3y/eP3J/qHA6eZkPA+GUiuhFq9yHmKLZRcznPHL/WUZoHP7LzN2uIcZc
OAyBZTZ9mtRZ+0mPbkrwZ6MeQ3LSI/kA2VH8/5y7FyZRoo0f+BVCKGvEwA6OvIDy4F2OkmvhH6Hl
vobo8J1Vfx+pF+WV4LI0vv6HhvaMIjfEwGC40qs5zPfxYD6JxycSeZg03LyxKk5f2kggobqF4bdL
dQsuW3ngdzQyyuLPCNTmmV5IrL5Lq2yMHVkziplLojft83ubOdrCVbek8rdIYMnuj7FNGkeJAPZ2
O+77VBBCPWSDbLhHPgVCjg0MxDMiKhQGmULK8CVMe4MadjmZbMArNmHAJdwDczj5dZtBTzPCoMre
LD2Yjg4x8qKxGCL7BDyzUusFOEjYHBcm8mrfLU0641O1xLt2alrkYKu8WuCUgVPqXQQBtxH3ra53
xFogComtPA+8vB9jRTRAsFyCoOKbKnNl9MfM3vQguLjuGLUllLKj+HBUwLM37ySfUHMmy2BXrkzT
ELLvpkpQO8Vu4JSnqmSEyM4Se+zi704JsELCMuR5O+XazBZHgDgcTc5HdQjCx4uzX6DlSG/YKx9A
8QylCpiKu8jLJRSxpEBMaDK+8t2PwFIBJKNO3huC01u/xhXErHx9E9NBRfi7OM/b8PLxhoLtiSH5
BWj434yH/S+xJGb/xu/1PbuOcK9bCPupBBaFylv3L+DIeNuE+lK0C31Ppjytnv5le7GQpPQ69eYT
BDiXj+jfv5ZaX+2oTJaYsdWdxCWBwCHfieUVgnsLHq53leYO0CmigT/X9bGjA/LBMv4q1sY7lQkm
M+6ddkwynq+FI+Iix83xyrf1EZI68mm6/57QT0fof+01Vl9chUssTScLlwm/R98CDaC2INBFpOpf
E9UgfhG5kN+vQ2LCviK/3jqfratcWNLkNLBP9JXkBHZlGdV93OMxpb2yg906MPPG0UlxRfxpOFt0
qPBWXSHDfsH7WluxOoZDxXiDNYycyn/cXaqIUjv6MLDeaAdpJTq66qfoHOV3w7/yut+mv/ysT41A
/4UyvcvhmY/w6JApaVhUFcFwXwXYLLLhaI5lDlLkCp4/ficNi+NaFa2ha3lxg0Yf9qEuY2STLznk
fH4+LNuJVCMfZubLupSgaMLnJb7+eyL4P/SAs6IX30tE99+G1t6X72FbcNi7xBhYCrR1cXKxre+P
/Loodg4RfH84ESyNqJb22K/S9xY4upk4KLm3O0DJx2nsK5Ut1uMJcAQLnW8WK6GTsSEXlDLljFRv
oCBypOxh6GRIDutiRxvqMnhAEtKY3hU9AsGA/nGkZSpdAnWgIBKwgdeAKSldNsH9OlU+m/5Lgbpq
YwHYzkqfCijZqrGdJccebxDfCYwnNcVVQXidnCXU8FrCsGkgFlO/7FiuCz+d7z2NUHzWjrtQ06Tr
oLZsNsSZlGUhkWQUsZn/f0hKKkuU5J38KK8qeoNt6bfyjgSS4quvL3ls50/OG3T/PVFag5ILS/uE
xNPv60cLxB/FcL7H3h/ZjnrfpJeD/4dGFS/bBGSs9yYNXrab3fvppI7/Z35KJu46T+/i3G8ek1l8
rXkJe0K/NRLPFm3qB694Q5TCxn0njoJrJqsS01J+EaddQfKOygIPG/jdsEkKKMREIKTK4x/uI4Av
TFQVKT7w/CpeIjxTQmNh55cxM2WGieY4Qdi6jv1fwM+9H0ZZ75n6zjbMK/mI3VHks7t8/gKE7bSh
G42mVBup9Bi0nzZFLimcRQogDocIuvdirMD0ZaKTby74R2WJflZzSYwUCTXQh8B0qzW9SucnPRjA
QzwgR+Xk86Pq4ZgJ08hAcVXkfwDJHmsu3j/HquO/OAFx3Mr3Ws6ws+wQCUY39A09/6JQRCffV5sX
I3VNH/n++9trxFfoAnVHp0rjqKE9Iskwo9rYrmWJ1BSziIhNkBse5QLeiCN7bb3jD5k8k0MS73Sk
c5ATI3Q2x+qaY2xiU7S/4edP6M7s2eD9PDosD96RDahC60aQQ4kEYJ//jaX0wsYVHwMfHTWq7Suu
zdg6DdqLCJKAFv1WQPw1LcA5wQr8hlqUooKfJP5ioroM9JCSQrwk/+ku7FvScgAAAl/l4PuPcm8V
1NLz3d7wKU1qUCn7m1AowWFH+AnYoy/Lx3vAqTp3QBtho67hDwR1sH/xGiM7XtSHGrtDgUyyhKEp
pZKzavuoCNzgguKQ6FDB1yjDVqJTj1YBojloVgIQl0z63zq8t8NuC4Dbigcp/fh70lumwylXrYn3
4K7MmtrYiZv3txT7tFRpAZuKqbanbOVSQT99ftanlMr0tR6yV/pa5SmNNJHQ7yV4feP3s3n7aqHi
pGV64YSeK6ZzxYcvfQRoclAswFaEieQXSP5I62/ccmD/DtIJdi4uXOm8MuQxjJYDh0A5ZCc+38V6
26s5baAMzjKebGxqbKM/UpTq9vOxN36BtUrFCtWovDEHtJzRno2eVYG1MRS/2mfpxdibWYSHZxCa
25QTnRVgkqQJpdJhKNDyS7NIxBeUGEg/fPSrsH/1H+nboAEIbGIKuwi7oYRAuFOVlHYsSca5i3cZ
VZjRKBskY/y52yqO/v6xkWFVxcQK9n40LcGOv4N9ZXlRaPrisyHTRJ2lBxsln/s0PwqRiKlJqlLZ
U/sf5M1TvZIL8MwEP8qouJzjQmAYPFu1JRykYRTrXJRAp5MsGvjrO97Om4k3zi6er1Rhrn/GcpoE
86ZfzNx+5kOfNvihybGFvnBoCRYABDoKvA8buhWbyG/rlj4HzObX+DcuD4zfNp5rg/qNW4d+H3kB
E2y/Ovzz7hqFG24m/uAi1H1uBbb8n5Qw6v4Dt4/l8brVgTnbrVcyNmAL3D4cebZr2FzSxIb+IRNQ
fU+Cmy691jW4TjwPUr5JvZBDs69mne6p37SVcKFmF4Rb5qpKHYqSnS0txU1mf7I40D+D4hEznGRF
2M/Vnfc7CHDG1TPa6gSa36NW9YO8icPjw7MfI/CbYvaaxSSY50jX/5KeMaz2ssFm6cK4YTxQiwkx
ofJFA5BSGozty5W1Jj9U3pz5YVX+d6CyKPqeXFOWxUWVuIp/LHUFwKz5QaXhHnGPpJrGPHeBfzdb
J1pfo39eZjXRT2hylZJSHLCz9hMZehVf/qxeLxNHCK24vunPNtjUJmRj6JqnZiJS091HEASDpae1
YAnuCTmFTuiKh/6B1q7PmLIHehxV7lhDcM5dzPb0ewQVzzEx3W0Sb5Cd24Cb1P12gCsZAJF/dmy1
fP4FM6NDmWMu80yVpOiLTfbtdCUe6ErplDXmkyIhlCD/TEB8t5nu577t0bUkez7FBGuKLzXzIy3/
o5a4l5Tes0LT0RatCA0Hzhhc8rClJ9lPqyRvy0peMBZXA4BIftDfaiEXT4r0E8rdIgqubc/3qIDw
nWGvhP5RlfZcvIGn9IHYtMbt45K9xTo/GxN3+Op7Vxb7VnJcg1J3NnqfNelFzMfJ8MDs+HLXe+04
jqoFZLPFRDb/jNnTqWt9UR/pHombvaQ+BAdlIRfcnfMZZQCzN8eS6hcW0dX7B6RD/ORaplKfBOwE
B4Wo+NlS/QZLXpMifF+ME0rhcxIAccQXxwcv8oIDyTLEpC6kkx3WdYbE4p4oS5H1A7g5F33VW1BB
E0RNnhI0sD688kXKJdTd/dRJIVCH+jlnDxW6Dnvbp4ISgl4B3AF6wIxxWyN0LzwJ2Kq77z0c2jUI
C/FlX7o40xDJJ8dq/O/JxdeGxheUAUqWcWyyTPQqzuhvokWKdaTBjaOQ4aGPigPo9JQtIrY4svcS
gNHMS6QwJRTFNi1qroxB+6Rbl7lBUIFE3dMY4uU8brVR+jls/eekK2rGJdJE/7LDIknDBtyL7FZ2
lS9ZWF41qeHq98nMnojjDfU5KjPCsCNwq+tn7BJ08E9vC1Ji8+f+VHi86hsMaGWeSEgPGQQeqPfz
smMbBG5w4WJbcskdciGSVgZUpu6/3Cx7KgcyjOtZ8U5jlFRHXOPwvMDMYM53CH6cqNmWtLnukilO
jTEOxey3P3yc2epi/WmpAliVy/adr+i4HYLWzzS0aDUtMX2LAhVi0Oa4OJvFsCfbu8eFE719oPhY
1mhtjIx/D8WzmFiD090nmbfR/7mmPnyfyGxC+qAb5tosdXSixZXXbeJaWAAQmIyYoA2Y+MX7Cs2H
DK8ozD2SgofY3SHbnPkJywzUkxhR6Ye58ZFF1lOwbX7FkIuGpM7FnePj7+48REKBYp29TFQ+dKlv
3FnyGKmVhWVLm5b/F0Xu98baeWYK3DfGhlZ2ojsqiIAFzYhDreQ+cShOYY6t29yovcCx4TgDID+V
J+Hv6wUK0qx8SXZsXaSgaLFrr0DPgHZSAsOJkPhOhVszHJiIQ9j6Gb2LItYTsaGSEJtBtN7tFlh6
q9xS/w5uMcAFcRkPj6dGS3nKv2eoJVCQuPNYU+84H0/EAl/fO+FY8P37T2dhNyLKu+CWHkH5qLo0
jMXZa40MXOrtwVPvMEAHY+KwF+R4VXMfRsD9v4RkA9sRMHTTYwpGd3Ryf5Uc+Hw2wMJqQPx09TH+
cWcOQBe98UfJQEeCQReNHQ0wmqYd37FvVihhd438egSIyCBa0r95hweGRyY8bMLfunr36kbEFusV
lH+nsVN8quiNJ2TKHcF2KVD48OAgpwGpgWHtHZUfcbTuHxeFKhdGLyYdl5SlPzYufwHfa+k9+mcf
mh8GgXbnoqaSwTz7vJ0DkN5p5p50uN0TTuES//Oe+tu8VThHAbmgjnCduo8UgNJHtv51Hy7Zvn7C
pmycZ7kDEI8dvX8nzjt+PCdCKlYT8L5jv4h+fNX9x8/jRl4+PmlJ7hs8coipSNkD6XozJIyWkn/c
ka/C77puzwJLA7xgpPtkduz0XIfj2pkZSiNoJQA7aNylF7sjh8J2QL3neWzIikQcwzBMG7E0kLEn
4XNNNyZDHVkem7B8z8AmUgqPBZTj+J5TXpqZ52FUkVLaqhHg72XJ9YrS9cDX81TRrfWbciiv015J
RpzA+SF1Mnvnzo4upIyTm/cxuP0Y2J09KQ9Ckr0ny5xtRVGGnYZAe2qendc3Myy7Ak2XBCMtiLsb
TfHs/aTqT+DxigbfXxH8wndc25xlfT1fkbiFbplO+DDTjg+pH5NJOPTnKAKTPWydN565S+bM5TXt
xUyegLbrY4vmj/SFL0MqCzKAoyGVRCcQhElJ0mIl6/z69B4mMB2scJcJf9xbhMNI3970OWF5CoYa
l3NpZhyYfPcSoylokTMYVd9na4nZ9Pc8+0gNmdFukVu+QWlqp7NGixO+PSKAoA7KbrbsOpSY1Eif
RxmI0gJUQKVccqQL4zYoRmBhWju4hNt/eESrHKcsvRAoSPUilSJtEj4AO61SzyTk9UYky3ivEOqQ
04N+8kEe9ywQMLLADJBDYjCmB0zIjDPTip5ohfz/3Cd2F5pQssNnu3FozrlEpQw7ISH8nuoNbWsX
AxQb8DuGY4FjK/HmbEkBSz2ThhcYpdS1ADhfKMD8l6N6+J2vPvqLp63CjWAXiya+A1N/5r2VBFSE
RW77klxqCnslKX2Tokw/wyv3lMMzWXTwR6anESbV28EkQg9Lv6wyVwcyqKdpBk/mqpyyewMpymwu
IjsaVDZYNbXd9BTJiMcqMP8TVKVA243aIvMu10nQNmot6dUNgI9w4kJuCIreg6WFyP89qv6A0082
w5QW2yTsAd350xvFSyJh/17QpBDgkH1GJBtW/GVmK8Jt2XJPlwkkz7ubBnixvnw+QYbPq2JgLOBa
e8x8PKqThykDSxiY8nuHDHXWwpi7azix9efHI7CzCOZDAH+ONkr9KTqpyMTQL0KR79UrZdiKq4b1
PjoHgOx43VEnlO2hcyyoCLAOD1/L9BFRbYe4Imlh4YS+AWYUx6B1kVBFz6o83HGwvBujZkCbpf3y
UChb0Dc/C9CPEBuVo5tVC3G6jXIBGNlEKaiGqNaiJuUv40JN+JpFFo/Mk0jxLnuz5Ssig8hU0CHL
6714VheDwHgQVGa4QbQAAfBLcl2+NIVNGsV7B/YrC2+evOyrG63jEGvZvSE7Sf99c2oWS4CFFYtT
mnEStMKUo+uXpNN99jp7gCbI23NpmHqMAUaBdHCnbA2YJxTKPg68f5DI0ZSSyHxp6IoQeCYJ5Uam
zONanNHyKZjuaoCRQGxL+mUqHUPWkyG443tscTyY/CEm8+OqjHY5WUJgycnemNMV802KpEL8fvS6
NxyTzm3dBoahkSpe/NIOUxxHKcYSt7gHjdtJFAEI/pkPsicBFcsTl834fT0+aBYQIFu18W2U4FEZ
AQCG3bO3YPzk/+FMVNVkIxULj2KWVIsOyG5172ncXEkZPLQQB4pgSLihZc7Gi0otAldf191k4nTG
0W4peexnIcTxGvXdiDbIV6HdpSV/9BJ76bNdGQhifmpaN8PMt9ZOxT0ysOUA+9TKKS9IrJsnbPD7
m5C13KYJeQ2TBKPDUltuHb+72hTd8kEAjF1H5uMj4Fb1MSOJoJ98WNP1m5P/LmBwwomNxLjBDBxo
7EbaE4pyHnlpGt34e17YaTmbyzT2RL+AfJUvGdL2BJ1BsP6UYj/pE+RsX877tnxhW1VR7r5JyC/J
5Y2PJvPly9D1bp6QNjL3WplYSt3WjZ6jZ3KDa4ReS3OOhknlY5kJ1RK3QEfrdhUQRYAhzfJZf3qS
UvqpvmwkITbVRV6Q5xRiV8jTLGyFeyYL1ob165vkpOw5UtKLFPpYxIUiEkg1665GAViqWBTN2Db5
5vGu61tf5GeHhv69ns8BGg+EUtZUnRQKYY9W90v0NlJmiew8tIg3mKoP8dBEXNrLVCHufz7T7TJu
jjGJn9Zlu6xcBIYnIgV3gm0xQXGupt7HUt7Ry5RTx+9dFMLY3IviBzpmRxnGglH63jMGIXjyKykR
zKb7tTwdZa1niJTgcO2ODa6OponWYGYjIX/RK7S7G+ur5+36SXbsqK4/j1RkYFxGlENqybKhnrda
B/7/LwnfDDsK2ZcQuRyfoTsA2qrB0/ynXdP6AzjJ4VHN+9HnZqolKB+e2rBGgsb1cv8owRXcEykX
quiHOQGlUjpMeGBTmJ3zj+XZ3ynJPlrTnXRM+W6bNk77EUdtUmjxhjxaeZ/QZVl840sxN8SznbOG
K94oUutBxQ2DZprLlOlzMA0MisJTUFc8T0XtXHJwU9RGmr8KRbw95Zu5txuFs+DBdjDv2AyZU1f6
t9XBhhk9k14cBsHsBgXrcr5P5LX+t8sjis+7U/LNNMXmYVOQ7CqyHygloLR8cqRVnWjWZwxT2bSa
ogmTw3la378/3SODLh8vDLF+9h1XKdIp5jxtoWB7p8H3VynvfAVv8nx8sVmZwlrept4uUto4Yius
gX1tPZRz7nzBvvXiPMStUqYDAq46qLT+K6QeAcqlJnXTdqk3rjdUX837+7JPyOyybyIFipwaz8W/
1zLLwjXO759lqUNqQCP47xkqA1Y0lJaTN0QdmBiC7yNKEYnRW6sD6qhRuvWpHCFzdLJjv5cngU1V
DxYqtN5Qz/uPEIjyrI49ix/tipOzh0d8ferSjbwYU4ONik/QJblOgMUITYwxiaD8hxnsBtLWJr3/
g8potQ9eJaylLiE54cTfP701WxJoaY/qTv+RkQljUJhwKpHZc+zKM8VaLGRpxlDBqIjLrB+ENqku
WoxbiWWj6xZGmhXe+oR4PaoQVJUsdKKCGeu0dJAI2SJ+dQb/+RX0+lkajJlUCrdVMO2vJw4X8P3X
fKdQJS0GBTgE+N2//eiENsdNxIZtjZe+V3Je8wZVu9gS+RI7T85O42Py1pIQEauIb8R/mo4whoEr
rN0jmfpJcClQJmmNt1uH1ZsdNwzyEJV+Q+gr31ocbtLJH1tgDYaonFDee4d28kTH2C77jhoIO2fE
m6L/JFLmbZa6rgB11D/aZ+9z36/63TghYXCdLz5eH/gpPop577wl6TeTEX7weMzNLFLUrtYqUFnU
nRAVgVxPj8mJfo+yzEeSl5aXBOI9CIM7X+7MftUN4Ef3kV38FWCSTUotPdhHzDnr9mRHNavMhmwz
KOwKxM8pYfzCbUyAPE2oCyN5w1Axs70Fp0UvUYqwx1xJCJfT2pNh50POMpo4i78+a5T9crjVay2h
dJeDTB5vGs+Bzr9bzeWxDaxps012hUV6FwHvbBg91jAS2RmEWHO6PI5jQ6XI2jYwG2RphdMmzQFi
69EmWJMLc6IC6qzLJH9EsEmc+Cf1NV3xDQ9BtQFR482SkUaKRIt8McQu8n+KmzHbDEBP99q10qND
n6zvlv3bNhIYAQHyLNOnTeD2cnQZRn221mUyi396ath3ZqV2fKFmy0FcYgUAYoU2t/OSqj5hH0ti
PCtZuztSeYPso7HWX6ngfG2WEW61ysx6fJ/LUx+Yd7VO+eJeslXEj+uKEolFwMDvI2XXLcIwn/nm
F2C4MbXPGw3pIkvtg/B8cw+hu3s6SExSrtRuq2nLT2WYt3/3+MPaMmeG0KnHvzickiYC6ivEHxwK
47e1R58xGpwBUoNTnJ6EHIRIplROsKVxkQOxoTjwRS4hPYvqzZnaEGv0zqbEjbms7JSQwO9oITM5
g1veesgZ2frsFP5O61T4ui6ept21z+WNP0S79RWmXpRgA6BMv+EZ8TpzUH5W2auSHkdm9redkmY1
SbrtwOZWCFO9smvHh7UkvRutzH17r2xi/mHQXGwEfSl6JppgHf3kH3tzTJbcxGbJJhIpmxRAde1N
Jg1uEfKDeuXNqggU+RysyR2JdAe34H0P/j0cVSGu+pVej5zn2Lcb52WQ4zMFvI6aYwf9jrRScd2+
+YBQC9LrIxoiAs5nE3iWAFvrFsdrUG7ioZYobT8jQp1HWyjl5RPKDi4tcEf5dwGCxr/r3G/CDiHq
yPEcDvMvrxX66ulIbjf49u7TVsLX2FjCgKbgKoYKHTYX+SYGt4nbKfwF/RyRzveWWe0UStXnvvf2
IY10VVnj9+vvgDQYWTKo3kQF/CccynW0mDZBsAhhM4McSWJ9emTE1+H5W1zZLHC78yfXD+u31wWE
JuT33e1IdYjrdI60w6hacdSdNUclvA5VbFo0M5MOpg7AA0O4XmlA4PuSLyfGF1cOZhe5k2anC9r0
6hKPg7pr4q0ywEfCv1L6XjdGJSRfsiMPQfcTV4BAUTTZG+webPhS2OJAqz+EJ2YNOeJUTX6aJIZ9
EnYcOnSlYT/ZkjT5Asc7IAOzPopYu+np+5Ju8ThF0Pd30CXzm4s2N0tq7DldMhzSmSnUAj5KunNH
NYzdq3f2MlOg3tXUibcMnpTHhxzziUeaEbEertV7Jir95X3TNPq0592zDQxwOh/0IKsj6hUE/ESw
4Jf6Gy1tXIPg47hoj095HhrPqq74X68Wlb3JnuuuBV0Sksg9CFCf3SRvD4//EEgWbYTP82hFuvaN
R+aV7dTEZULFbfvDKdw9gFCnTxfzqe5xaqmEGh8YhrFw0MjdCzYBsI0U2YAN0ZUJVSY7po2Ohit6
dSpD6kG7/Segw4lSzOwJ0JG8G68c0ABU/txkipBvC9iNWUpXUpJ6XWdnzwq9EXVa7UxazloHEtzA
blvqEJMwO4zv49bCVRFyhqM8cCBNL7IOJ9aZMoa8TVeHsMRQNT4+8DtJBWy76kAW5BTxdYJSd8Kw
2u4168DS5hvFVxEa5fAW0N6M65vKSOYkLR6HSbjx0VpDfkpud7GW/stU51H8Fl5GeYpH/wHCbP+8
C5aF/ARKWdODL8i1kiVjjSum/GCTWGfRJZfrvTshvoRjWrpAApzy3uL7ldch27zKOor9vpJQpM14
hjznx2JzALl6jlKe3QfxXloOJNn0anGu+jesm7Rq0w/7vwZeNflZUEtg94tmMj6h+mD5RRC451lc
ZPLWs72PtsKL2Qsw08WQAwg9Rq7DtPa63XZXTyb9crUIU2zleTAPdYVmrdRYUMnCDYYWjE0K/S8O
NEW/ZazjiOSXJBDFP+hFzF0Y8XWAR+ba2yaNFymvV2eBhr82a2NnpF37STfvNFqw078Wy+6tnjWB
qLiPbvlfqPYZo0uGd45sOfIrxNFupohXPzZ9ZDa9ZaFE/AUSlLQNtOfg2bqcCd7rYUNnxs2Hjyer
4JGbGsyWNyAUJl7rpQMQHCsOnycsvfWgaBPlPZLbVS4LkS/lJkcigIvt7MSpl5RFoDGow8rL5Ve+
dib0U16o252H8Qpgz6g15YuJPw2/1PL8ut47Z4RrA7Fsysn1HF7HpdC5b7K1Q0fsfZt3aa6oYZb0
nKv6XrY0hnPLvofiOeP7POYtolz9aoCxg0JPKICL9izHuhHvCmH2n36AgmZkM6rP55VQgLAjo1jn
E1hEmclMeYW+ZYHPuLHAOgvtcWTwm8C2kr1PSynJn4LDEUUHikaB53ML28qmEDXmsbfY+W34p7BH
vEEN8D27y6d1ZOhC64isLaB3CzrwPkAXAJoq25LNIMIm9hcdSw7y+xdj201wqEuciGpGAnTUqJeA
oV13N8nvRnDzbsNz9jSS/AMMAZrzH5z0CzwyUuzUVw4F+SI6YbU+wRmA8VTlIOXW/AsicViLs73D
5hKDoW6uwDSbSfcKk1+drfzCk0o/A5E8WDLD6o1TVhlRjGCW/bx/SyeikeMv+r6bBTUDrk2yW3qk
Uk0ixkrc4ph9dei2TuJ5dgnwHe52P6dC3n3ZZUPs8IfOU4Cn8eVVKtCHqUtNpaYbg2L3i/5NFTJT
RzRLIgq7TYIBkBXGk/iJWMso14yFLWGuPvJDiec+7RVwjulPW7qOCs13b6HVbuIInBvVud5/DqzG
LeBkAFZ7vW47rLHUH2uEriQCi/YoWt1j6AzQmcN5AXMYbIpAARvHasczqMWshtqKTV0oCKRmCXO9
+tIeos1Ceixb7ZPOXpS1JOXMoh7Eemot+ztjmfOqBB6euCUEYsraQ+7nVmQlv++nwSsInB6W52CJ
Oc6UfGpFIeGXIjV7XchjVU7V2areY7tsvGTmbZwFRdfe8g1iwI625ABOw+ey4lYwkKDnxNsIHtR/
BuigDINlf74sA6Y8QASb76zB2VeFH1plP1MjltLTY58dJah0P2HKnpqVTWTiDKrcoKdxnE0Qy4RE
IQCMIC2re0fnc3axGKvhAu33T1C8ht1duNmkBP/PNMFTDC5oUGuhxlPwAusNi9rW1hHsmcSNpZnx
lf20HWUkt00YYIIyXmDi349cdi+Jscz2A/xfQvdy8tBpfxAyEaBKDW1z9cCD+TbAC9nkkTsB0w5e
T6kGoLPw5A1TBJf2ATWY5GYHK5IJYJqjjur5gU2sGAr7KG1ErvRxHj1pKaaXMiPJ+1uH2FtjHb7u
U47YsVlsriDjlOmB+pB8BtkTLSS1mDBy6zhmbU9i/PE0pAzbVgyoZrp010BKhMs8R92yWUTMXV9m
hRxhdxqjvGZUpqToHOOUfYfVUXG/jIi1jjKlauIRY45gdrtwCRcif6sQnJa2cZOT7ZO0JjAWY3Et
0SrQ9B8yyeViyV3pLEcCZFFQWvlVnW/bl4qdauZcmzVwFRI5farfDWvO6cPW+Xhhp5JFBKSikoGf
+OinNRRkbHgFdsU8Hahdukh1Je7Pn7OyT1G5JUDNidlbVfqmLt9XfhwKc16yDsA1xTbMmWGrdth0
4MiIQzkMjXZChDIOvspM2hNqrw2t/C9X7+YZ04DsUzbjEKmEhmnBxbyntAUJvbcx9quJG4+GBP37
oG3IxAy/SwDfXHPTvqXQ9dnhAwnALUsoRTWMYU23DgNee0CMZeDFrB3HX0z93tDl6mrBUUMeY9EI
UQNPqPxb+pRSuk4FwwQ7iFNx/t3vh3mmJPAHA5JKD0QpfpJFF3WJ1FmULyrE9ZD/TWwFHr9tnM5v
udGKhNGIw8tUeqBl6uYxiG22tbylXIaY+cjR3IVq7MFTsnP30ICsHtQkbE1hGYPvrXz6gr4R3Nac
nZWcYQSKdqNaM8i8sjmWLxFwUIkbK3119v8ga1ZXxHawiJzkS64I8oSNQv7U5fVasYP5qqLQY3xR
czTZafuDiADEPIIIwnMN2D5iVhHPjvRxgYYraTHZDMnS0p33PqrifBhMqvxrBr2IzIiL4qGvNkaV
WYesSa9vyfltFdvejKq7Ly3DqFFZN4Pzk5Hsh4rCCevoMPI6vqxV/uHCMm02AS2lxS4MRi7Yhs3U
HSmW03r/zwmw+0Fcxs5Rn3YP8OxE0RIQw4hZEkd/1i+etglniVvG9FR3fgmqrN5qNCDGIdrv6fFT
uWtn+IKIfl1EfpziNXMq+QcLTtmckZqIKb6jyUXdylYrN8v9p55F1wSszA7OtHQVQde8zGsE3XjT
z3sWbf2ymQ0OkkfO5rX9b79Y1QkIYvG7T/BVRJvoare5nrpfCdAiKmKTrrZ1mFlVpC2a3HbHrVRY
2ggggpHDDbKoEbvhsGeZbKyn0krVfrWWQ5EApDAjSVy6xT6kPBXq86YVM7YFvfzVpK/s0mFB++vN
nOSwLz+Lze2uTCOD1+dzisLf30qFPeqe8y2KNeecbfaj5Dc4Lq2U+5OXKmXX9/2k6/iAn51RaZ8m
quLWeSdLhnUs2MCG/uUSthrsikeC+KdrF5Fpm6IwE4kj7+Z3obxXxyTOEMptlmvie0NNbpBqOGkN
hdjkAdcLRaH1DscfHIRHgylXeN2HDWmVH3Wrp3cK9Qc6B0VzwLAtGWEePBeHYgBm0+GnCyjgvo1X
djWZtUJTIztHImTUe3EWYIhBLnWpDy0xImWQZXVi6+B1+w5taQzbQH0enidBTwXaPXne/3GVrj5h
GlfSKjZ6TEtmCbtzERpob7UDXhLgjDeDyDHeYMSgPf5jLOgTKj4BRCA7bA6XVn/Vl5EuWpq7yQSc
C0oX6rYs8fz2atLKG3u6n5dy+LltYHCBx+vmFixhCiSbGAGVMeebyTLZxREOCpm/zg1bWtal9A1+
MX2aeOxyLLPOHQn07nJIGhFvsRIfzAMziCmbfP2MVR9MDG9GBzIyj5Y1G/YAXe5jLLcIJB4QDHf9
LTST97ERHwffEURPpgCXAowup09K4ti7kkfMJmyVK4Ye9Y7MzGGV1miDm3EVVKSD9b3v25D2GTGy
w4+x/VlYQCT/OWpiFqPaUnMKjVp7/Em6C7u0Ap9ImvxjcvFOrcXXWKV5hM6vjXbENXPZAC7oXm3z
6QVDNI1J17aY0WTf7HGneuClxlk4ZdQ2IYFnj4N2ELYDymqJVTtIJa8UK1Yo5vcWj3KJDinbmLVJ
IAlEDNPZUvd5XU3863rFDJjV0vs5sHOI57n4fv+fk0ylX/EzXSVSwi4er2C/ql88Q1cElHqecng1
i4LzKJttMRhPUVH1CyMBo7Ro/TyxZi+8IGtt4fSb4PC94p2kEXTOE7kKWR6dqHUxLiVpoqx5iM0J
YekBLTJK2YjrJo+W+ufgsQJ7d7VrTG2q1IEb3Xt0cc1eBbVdvuPMv+mJItuxQ6pr79wQA0fm7VvH
za3D/i5GK75tqkGVqLvZD6/2lf6Zj6iQ6ZaYy/L4SW7ziM6AJieTtaxMc3NT7hVLHdtg7YVuChwI
IyymvatH30VSvcQq06j9IxkQMssa5zJfXhoTtBWCceq7krxgRaIi3pChVOx1lRuMLxmoQ6sjdwmr
3TPfu0jxpARwNorhVkjSC2BBFHMm26+mmja/2Ba3B5YdEwykFkwofbP+e4dN8XH8oXTDZR0ZVX2C
TMW3jMS0s+1xrMrEl5LrptHgsjpzLyVSLj1OxbL48cpG8zTjjH6NOPwncVhJY7r7B6w0Jcli86l7
s1EoM4phYOSpYVCKKmkM9N1mW2leI/4agIdcPbElRhka0w0eQ25ixgH7agnFtnm5TwDBFzByWwrt
fL0ggdFDkx64bF+EO8/vFstkgg0IF1iNnMnzUjCgcfUjxXOdPc73u3Q4oIndzQPBmyTpxPIl6uow
aDS+rCOORdV/3//LJ2jpRRcZrBhWYrwgATQS5YP+qyMZFBtj4S1tSbeMHdzuDCcziLvZ4hqOX0mV
A8yQzQUc6+oYp/DLEqt5m3NuIplrpQVDsaDSv0SB1ANWDG1zFw8+TBAYWrnBdAL/H4sRI5UHCNsm
BPoilg4oj82v2i4IMsCTEfz2pvUq3LoRSMBdM+oWUKek/QWbD9kx1/Mn0sH1igDFR82RD95o2fAI
kIJNPBGJg9PXr1dUPWwxvpWnvXDaPa9aIL6It5nQrnl/wbchDXw4NAKLxs4FINXVQjP8ldBGdmVr
i/Ox5SUVE2T/XwtzMXgmRGjhIfcup9VWfz1hSTLN0r2A4ww84roOkwE3g88AbBUtAk+sx2XF56AI
Ih7kUnyO1UOHf4Mnslpp77g9Hi13ikKyO5PnaSgU/ybslPKOEJIkK6RegMSVDw1tjFXMmQvkA2Qh
9C+p1aDw6PVvqpZhnNv9UM8xHDd+OH107l5tbLvJGOhlxIkyFhzKmSdIQh/bix3Ed4DSzOJ08Bg5
V9P90DyCm7BFr7SzcRpkedRAMA6vpjtqrRJNvlixung5pBJ1JDhb/gkfk52k7muL4paWt48B2LVe
gEOpa+jF7oCniZ9wfpZT+WnYjebtz6lwE1/rzwj1uqLg11II4WfyrXKxixxresLmjH8/uVyqV29T
9G3aFROfg0Oi5PbWWxdP/RdkRkNWiOdQRPHVZH2v7n/dovXW6GY9ZBMBYHcMA2+pHPtLzEVDXmLV
IL0aoih6+gG5F34EHlj2ti4lsRwgywBB+Xe5f6qhZAwkuEVGbXZAvyxMIGRsglxX9DykKs4afXAH
vgxpcexh6brM4EJ1Prqz6+cLjWc2gzCe+wkmNAQkhm3Jvgtk8JpVIrBqhIzPQlPjNPy9ukuG2MEm
XjFfSX/z00U1PFU1QhlgxV95gNYHo1Ol1zWrO0Vc7pmeHgqhi7DO7SGuvBtRoucFQcGcIXhnKc/e
18ewyPU7qbWbmJ0zqK2OR29x2pkTe0dtR7GsyVLwfLIku0irUbiJ/6oML0XSFg39CfHz1r0kI86d
QpdxasF9ZpjUn/idr1y5QmteX9LYvHYxJwUb+u0AZo9MazidVA/I3A98KTzOl3Lid9OPKXU3ks17
0y83LCMsL8T/aodInt0YB29Q13pb+gry15LvxkJ38GOTmotKXD7NMdSAAxD2+P4duyAuTjpt71gx
uNrR19i6/FSJtX+MVC/2gZY7Q5JdYs6liDg1OhubUUXdPMwBzs53PDBk3bGswbfi2VgfP1jZV1pq
UX4H73nO5WKlOnL3XVBPeKgAkJZtsndtSYY4iqv8BFGImZ50z4JCKqSFtF0iCOXfCCqXut6GFh58
fw094/v/4IcLgTxYReRbfNmqBcY/Gnu7jfo06it90r2jIRP3YBEZjpeAMlTdoeKjTiFb0JL2TigI
aDmw3lSCWtR2innw3qUJOJ98ZS7P7sRArNUrZohAHNfO4IZ+xyOsbtETsxo5lr+3+myCXyT/jLvG
YGmYtWRTe2jFrDjgs+XfpavlhE6ffFB4iGN/3nBYOSi2AKyXPwRRO2NuVoEnIehZOaSDd0z1x3yF
rmhSgzeh+trjNLd4gWrSxV7jKC7pAtdr9nzG7+9j6gWAluw9zzP48/Yx5naTr0LtMp6A9o+FnNdt
FBWrVuXW77y5+yPTH8mdEFjlhs2l2ImgUZ8cvaPcGWp1Cb8WRIsLz31lCmGtbisgFbr9c8xVp7OO
ak+TGIn6ur02McVX3uCVno2KyWzoqlpNWGYSmsndyx2MRjnP1cCpuIDo8ndkg1g9Tw6d7j7JHztr
u6hrV/98Vi6ljp4qLSxC0NjlJOp/exbnoICsF+JlGQCnukUnmIxCgT1oP4825Tsa/cewCBFoIMrs
P4r6x9EUiHwQl29etdJxxJyBkurWOwV5ZxhPcCyXXVUXR8yQj8AUMYJz4wnWZNMJhvdmH1r6mAwd
2fGBoGy0s3LxfKr3AHz1fTrjNmPxtPAnz5J60KREJ/JRrUa3VeZB45A2rq1n92+d910nk/Rzu0pW
RZLHeSv9Or98lDuHNquPPYSz5EtQZ9ItSdTC+zNwPCmycdvckQ9yGmH+DD4WV2neZasAMwWplaEt
5TzKXWAaVqHV2qo48eTmacG2JXnJwQB8ZV28NwwZLm0ke37r4cAfCO2RBP861GZuYPHlgk7tJl5f
Gx/+G+aaSUiomfgJx9fNqx2WTYtUKPQ1AJuvwcF5wZ1BLHIrhIH/TB/BuJo79ZuxcG52n3mIkXxc
cTxhNcWGa7yYD/QYuRqLU0RqkEJInkZ+8GaWwf/tv9PT+dlecxu95VPubfzGeHhxUj34qjpRQzVL
hXQjcwiDZIXjhr2tr2kNCY4v4KOucizH9HJ0KrsOT7qGWUa1hj3myHRDs8EXT/5Bsy4HqpOY+gYK
34am2qw/Doec9i/9RHKIhDcbnfq0gFCK0UsDIxHOvSnDNbfF7nfJ8GwFiAq3ThxAeKnXtC8/su9R
dLPBgiezmowIAPhMfcU+AX37mrbm2tVBOmbQI0sbB5X/hwBo1LbQaTrTBs219latoqGzX4zGqeBv
UH/3Zbk7fg/rWJQAMzFCW8He+/mFNoAApz3C61mWaAEkdRgXyD0Y3qwjEgin6LWDBzC3EKUxKA1x
JwHn4b/hM4jlaQzC+ky+bJYKD5WaS1NAJuQA71x1FpiRsrK2MuaEZznEUh5tsQGK9Oo35UqJSI51
0+TjSOYfY5biWjKIB63h1JZ+mT58JQ1T5YhlwJ4218MZkfTxfMTWW4Y3SuDq6tOk0SlSbpf4eg2o
yj+rje4Pb+aOINzCqGzXVhFZqQhQw4eK7ShcrFRBGnMh4oXAAR9q9hkKK5Y+onJB1J/39BTzACTW
FrfET1IlCdJyxPzONZ+QGSEmSmDzFnm3yKLnm5+mYFNX75ZWF/m+cRnZS8g7Kk3DWt1HYaKCjZRl
/bVds86DN0/P4M/ZaiiwExVsEIBiwppjd2cyOe144gh0DCDc7njWSh5Kwf1+Hq3qXzEQ+TJ99FSE
zK2/pJlkEvnPTJXUgSYR/c2tOYIxjpEADp0Ry9Fb15bLMho7XyF7DGuZ8kRgM0+O+piab2eg9pSG
T4tc7wG1otmZK/kGwzf6SaaWzECc67g+yGBlOb6RLZDcE7kW9/DRHWEmBS2mb4/J++5OjlirDPkz
EWSEQQupGsmLp+eTY+t2DOVLO7P48E88oiPcbmNgAp0lHVjecbs9ko7jdDfZihxTGz3SHHPp1Lh7
momU1XabhjwjUlb6r9dn7420gNgG6adgPBgNcfaG/Z+h32png+AjwrmAA3mfHRSgZc5rOnp5Nbru
5VW0F3sEzGXT4jJocEhQtU+Ah3wzzVOiPq2lCGfzNmKfQ1by+owWjIJau6JdNTP6IlFB/IigOgFd
nrHBfIt0q2jol1DyOR4LJNumT35u6b3QLViI5/XHPXXFade2rpOifH0W9vfiickt0wfBBjByYv5h
6VAuS55uEUSKf3Hk0dEe1ma8ye7kaOOSlJRej1CUA0l/TaWSQZNRod/YZmY8I7ZtQyc0ndeA1Njq
drkMKveFSgEhoKkQM4STyWHpz5UwDB7j5YYZWQaS0hL/Ds8xWFOpcKgdQD4VtB9qz+1czEOl4sRC
pSHpfXTiwIewiJesU9Im74wPmEtjcWpwJp+yv0edGCD4D7XK73p8BkTIs90OODHPzkMTt2+hEqri
n7vsH/PutFMuVnRspns+Fvfr9lXicb3+gSp6OHq3uMpsc8hxa+YNmsV160Xdv4Q3A9rBDyugLofp
gZGgC1Am29YIGnEzq9e7XM4fwIOe8gDr/MAfk6y1eqlndu2+Vg+ubHDtZn59j7HZd8HtTa0XxGgJ
kzDQkRrgO/DehipH25MMjDPFuEipHMnnjQG624GUaqyB0NNsKYb70C19ZX/QLR1/SrRhzk3EQfuA
tawKHQRPX5Nek+avHqeLWusA0V6EP/2tMAhxCu0Qp5KWhtOSBpneAJVaMdRyHRLvJwB/AzWP9SdD
MvE0YTdqAipXaowOowkHFM8/B+w9nLhSE8vX4BIR8x7iCW1gx8BLjkU/7IY5cyNVW/Sv2Fz+wWAD
Xp39wyElE8+b3n3XW+1eFmxiYhso1JrYY0Cf16qBMVbslm9xK54zj/t6mWQskBoItdeLbkQ7Bn3c
78glG9urH14YhwUYm+vNUolaeFg9+a0+P8WJH/Hs5wXRNhc1HBiBFn0z58Y1T5rjuAGXzs2Pmwae
OoohjlpAgPyhzPDvkZZ+hGcVFfF8jjBL/uQTJbaLDpNq5I7OdJU87BEI+iWtcj/1G1eH7qrQQ1Bh
N0puQ6U1YQMzQAYY4fREq65HsHNmQqILr6PCwd81flvIVUzwuoYI7XEWUPR10IgUTN3CQmG2zwyV
DCfbOUR/WwTe82k5hTG4PlJome4CdIDh1n4IBtpHeemY0hXLKa9YxanlNKbDwWroY6tZkggaqgGU
BS8JAoQINbYZW/8XTa7bmhUeYhIdVcg2M0vpcDq991/QqIAx0b7XreQfQvjY2dNUld9hu53ymPMX
oeO8NLfmbd8faicPRYsOxFItQcBz3BPIGApZT+eoDuydUhqa3eF5SduPLEsqzc7P0yOF9MWwvSAS
ETiICzm3etPCa2ByJkbv62xtLQSm7pKqENj7DLiDGK0XZnGGKJkz/KPIItlBWXOZWSIqn7rL7g8R
+5iHZq9HgyGEZG65GjVR+uZhwIlrOfhRlltWTOMRjuZJTi3lvFi5hCMvkBwelb/u6ZGvWqCOsGTt
gC2Gl+7Bs3Q9JNX8Dz1g6nIi47D4QPH3KzYLPfDUCo+wNAJbVSrSqIm1VWqF6DQqVNdH79+5C2jj
069YaJfQs7SSI/V5g+Te73sGqyCEBIzpz8lpHRZo49lvTzwRljhqWAXASwS2w8Tlal0KYAUOBK9n
DpJcO5o711h1EAqhjXXEyn0xXkZ7EB+Rat22bTFNgmXw02h/6adhqWE3TI7rST01hm6LNESmRMTT
fDk1+jDaHER2fEvnqDHtRjsor6w99MfCg2uoWXRkThRK3jhg0r3MWtkrQW4dMIzwwMgE+btHVB4n
pUP8T0kusXp/2gQAWcLv/BnZxEYwtWHVUdAKHTmEhl0AgpMHn9KgpAQjnIytNHtzu9dEHWe6ZoYR
bf5bpZyVBJT1pkSJsaLB6FvFClB0fq0jp+tEkNUViI3DAapdxkmT/e3IOzl4jcyfGwhGjlFXVz3b
wN2zDSJ6ywr0KsZoQy/l/mT5X8ZqBTGtYCn5rrZhGmYNpaNLOyFwB4kbMLCEbHuAgRm77afPEtfJ
EBhGKmh3/RPl1DNzUIKARfjn3VdlWGc1SciJ/d6IQBs/Ln7sJMSk8dnauDGc9FEt65qg5ShLyrX5
3Pgic4R4FkDDNR8gGGUpOcZ73NIx/Gh7ZnOrLJj7K9rWxHMOVwQA5ar6LmYsSYHT6+eq+Ut+OmyJ
djRpbQnYMTNd07K6q9yBmOVjmAR2kaFowsWBYjizXPUmNyOEbN2hHCCKdv/o+Ah4ScnZXnxT8PRK
Wxr9GwLKU13ijGiB+uXn+zZkW73L2r62fxsSrFtHBIZapfRz3OqxmVMBNC8JuXC93PjvnPa7092i
L0NlPnS3Q7ZziJVahFGmlJuQ/5LDJF+W9dd5/kQnPo0r/7VLrVKU+DGbilIj1VDVg9/KvpRXF2eI
bKfixrRYd3H1bLSHiOvYHgbmuR5gNmW3YJDrqwQ5SkIYNrZwVIuIxJEaIabukyvJtbuUYi/LLf+V
TxAX2Te/dmpc6jNHZtbOlm8Pyx8h0XddK0KqKCf1xVkYfYupuOsoytRUYrIJsoVaZINYvZDpFegZ
tGPKHTSejJ+xb+d9UzbTJyHNZWqAmmQV7xYgrZN2jJLur7ffjEBJE7sIPsDdESLz2A+qlqq5qV1w
2v9/Y5Td8U5Kv1/nz9BykWGsHy6GI0poGhFTM5dDsNuaqRUDjhrJNhz3GNMsK83lgcaAXJZIm+0q
V/AN2t1l+JhvRiTFRyeqIjSQzTeRPZATTpX3ifgm4tfJ9jf+kWAYtXYJhXvZwSqLu4AKGuiwksWf
rffa2m9zIGY1mKGtlhBL9FqVMIjqfW7Z4Vw0rnjRQBM3yBtjpiKFEpcGaX1Zq2K9tfW/v60t0Dnu
voehZCy8ncING76LolFOB1IcsljCmeoB6tDQghFa0dfquAg1QSP7TDBBa6TOugusILe9bkKn6GU2
/PVW2nlB8P20VbuE/HK3W9kPKlsT6Lm27I35nTq8FjQt1QjTntsoi/ufnnpdt49QfOZ6ttZGiIIk
EScT/egpPEeUSU1UTvs0Myi0zQqoiI8WlRKBD3jRM2/bF4vOUmUiKUKqoY2lAfaydohI0MF9AEXZ
aX+PRHMdLKe2jdrvyqNgFSdw3+Ch5yCOr/acin3LNoMNhipojEM+QvWuGHxUY/J3jaaN7oSTOUkF
v8THVj7un19NPCr345GvLTgyMvHWHAtCtt0UD//PAD4v8qvG5wvTcQg9yuouvbyF1yzevqfiBpig
LgToDM5/Ubn1k0793uaiXnldQ22ZjfgwZVXvtYkd2z7FNiCIDTjnuYdhsWMTKv3dqxlybCn24WMQ
SGyOb/KqF7JP9AYnCdRTlSLzM+Vqg9r1JLeuHKB5eh5yFC0bZvva/zR0G+CXBj8lkQnjWScY3MYd
B4FN0gssVFTxvBDCRDjsIftG8waBa5FLVip8ecoblETEhBbNQhhSBLWZHu+4jaAwAyMlRbjX8Gfl
LNfTNEZf5cQYpVtQANfyZjKYYY/fyG32S2MMg/XxndLyAgCCGN4GScO6i8C9CB1RvYqzdAeE2/3J
Sds5exirFt3eRs/OY4LHbhM8H7MzDyWWuO8QQfJSWNBCEb9wUnTF6CO7JDraOUik9noXKG2Jm0Al
UYFvFC4G2BB+E+InD73TWx/taoTY2Nf9bmnP2Rhob/ktu1Cq4krt3f5BWq22bVv41oC823+OcwRu
b9pWB6SM/cEF4HERlGAQQw7zvydJro0bx0sq8xXPZ9r2daJnsSIW8ZeKs3RsIt8GQUgBYWSMrw2k
Osa+ReqiXYYTTyNynB1LlbwwvNRblV08ww8IFEjjCOF7h97pa8O5gaq20Ym8Bo6jNW3dEHvDx2ol
LvYlfL05Q5bH9Ksm3Q1VgmXwj4ba/nefq7eZreJSrNdT66N35lCvWITDRWlTFd3dQGhQuQyn0cbI
sOPv3f32pOcTflhwybEibTXFhwxMgyQdjwVHetsF83fo7qplxVMR5qJLw4Lxxbq4yvaloWvYBD7L
Ut5olHhvVmSK3xIUJcZyuT6UFhOSoWx4R0kmJ8zd7IGucAUQWlQmuHRbr02ITyiDS0y8CSfoxJwC
RLYcz53gaU0Hw8VuFCuf1vA40fecJJMZUC8I6/ExQbLj4DBJzpAkCGq+OFzCePPJdNf6n3+NDiZz
wHy5HVrBuQOaTy27qds5EoIv37xjFuRlBXoW26ZuRNUQ+Gt2kyGPD6rWm4yxPjCJEeUggHgeYauQ
VBIKFf7N15NqVbZLB3tEe1B55M56F4omeONC8KBXbl9WkTyVSLZtB8fGaBGERPfJ/va79x1w3B3K
pTsBiAfs++EK1JEEbRs+pfP/x2rzjKUq5cLZBpwz12zCYEMKRR9oPxJ3bLmm5FbwmiffaTJCt6cO
R4MbqC8sRYhkZ9YaGfuMxyY5TYbHKQtKHxgF5QSyiqH+uHBTZeyd6EQhJrYV8S05x6OlGMgOdd1W
GwMDZzMv83/y/5et9hoj9qLrAq+rboH/PuBWJdXG8M/3ft/GFsDzlkloT9C1rpz9Temaize1n/Cg
hoOgz6rl2qLZ7N/uGY5dwSVGsuAt7gJe0N2kijXF0k8zsJFjYFdqXELbmSpJHAzr1aqn1VxSjFpf
q5vmLgLKqCjwiY+0qhS0ik1xF5JLyjVsEBpq7aD6/e8QL3kdlBEmRsaekYTPRHDtTljFEyIYLoUf
WvNc77CPLpz0h6D8s507p1f8Hi/XJYYSVxSWGp4ee8KNZ9+O2NUL55paOQBDKRmqcGEIt4T2AB25
p8CaETj/D3FhtHFPjvRcYqDma/txwU246zBZmWt39b7mpOkrE5LoxTDph1jwkHzBSQVDWdaW1qDi
3O/7MEuCUB5jqySwbj27KzLbV/Ixsp7+R7LMxeaoekRbQs7BhYf3vqLfI15rLoc52x/7jH7LrYMI
s4zv5YM+KTsq1mB+ztWu12KM99iDpcvWD881QfSAh0yHdiWvoXd1RF153cx+v9hDf8QpgzdMoFtd
2c5vDC0vQTmsZ7RvmPzhf28Pp0Mu5lIy3XPh3Z6qDjL2wNMuY9v9vU2Veerd8oeUbKFv3ySEkl4k
ccf0C6N+86WhvxtBspXvSkY3hQ1dFsRu24U+KG+TKu4p/90qMHDAGWeZ6Q0mjN/d106Cbgqben5c
4T7KvunCoHMz//j4XTp0N2UAALPomSBrL/hHcwi8oouotAbLFVPxr75KkmtTZ20V7FGEt9qTZ3gC
VM3Pnl4HrVY815ii5Agoruy+BwT0ITvmRwSbdaJMwu8/EPdqDwlTNu70VyNeS3CbkUMD3U6rKae0
0R0ZZvAKC2bw9eMtPLy+SEfMu4u0FEI9t6a4CWTZaVg1jnDyblzrapcij3JDt0AqWAtQH+GxFtwO
FZ9Sbyf4fKseZMXWlXRZ4YyeS+I30cabAfVRGSycMvD53cTtkh2EMRHKf63xCJeNnriPm/bei1Ql
vPutVGf0ZqTRYIl2aAERrO0UegtHUAVzVzjNktUiUL5wAhIia+sDWz8rGAnsXEzBwIOiSNfvzdJ9
8xk4kmWbmDZ55AD01JM1L/9ifoW+1Pspbr6If8b96GMhHuAWV7Wr5zs0ZOVK2PcvwTZMeomLE3L1
y+Wu1JP9WQaVxrBB7W52LiDn+dPSKXISHVBARqPcSasVDtiMZaI+kQsDsfmZohVvMVRJ9JKa9uz/
e/MQNtKBe9R/uAszNud5LLpo08NR/sQmy2keiaTblGySHAsBoVWlYQi7pXk4Qtl8cLQ6ggCXQDH8
WJUPSH7qPDCbQeNgVIWUz94egzvYS20t++tUiCemtoAqC/q8JcH9HBOmNUZKdxXgNOT9v/e2E+xf
XwMBv8JMUtWjSy4mWeNZnw6BoVWKZyLGbtRuSpopN2guA+C3qcdcKLqfkUBB2BwbB/6inZY9gx8e
zJpyXpbSRALWrsnL3HsdbXv6lQ/YQl//+94STaze5PktXvT55c8YL+qj6XADUQK0PDgo1uRNuV51
B+qcCDi1EsErRicDFzCUaQKz0PrU3r0acAS3/vZnq4jflJseMQ88iUM+KYNd/X7HldjigtjCjP84
gKPTpyczN4NGWPVgNnCRh5JBGI8e2QgRcTNvpct2gq2d9gpTEqvOns11sAiI9RsKgeud36KHA7nY
9swpca4fYChXAsTN1YC99mQW+9v/H1T5UaIE1z2FgXsMdstdMMPkUA1Y9XJ+sO5TpD0cTOxN8AiF
+DgR0qyA7dQvAAr/8TTrwRSzBWafjWIrxNcTgzgSApoZDhctfN09MSD+QdPyo3CiTatPAoqiKKTU
90HXTBUUFly5aUGgqZL4zsggiDXmx+ObkK88BP5rlrqBj1N1g8izWOi5ClnJksiFofw/Ya6mko5l
3sUFASZbn1wXu3Ih3VeY3sDn4L0NXfdtM+UCHPOu67/Qns+ah30p6D4UOChW3+xGmYi1yICCYmWr
Q9yCOcGBlmHANXa/83KgRqCfL8xyx2z57T+4RMi3VlST3fdUTiawv9xBTNsgfwkdahB32iq+0vgK
MYCQqpoTPpG5lO5E6RqaJ3J6O6x8+M+4KJMVcIxvMW0vUpoYAle2ulfb4fCOiG7FkNUfh9YMcNBJ
xLuW4qBneqt5loZ0BvXsKq08NVEItpVdtMl3+CgeNxAQ19xc0KBcML6FNUXjTGX05V9Cec573Mtl
3pWQv9lZoS/TO1TDyFxO325HRtSXMamDs1A0BsG/IBE49SvImccdA+zsILbF/2cCXrh8l2D8fm2z
PcPynNffth6EW0hPfp6sOPpd9lAZOumLwdjpG9NZg8s2kGkatErbRLZni4zgOKE28nGeFsLgHRPG
kJbgDdVyCFaQTAB3HBMpD2Q+8ZjmGOqvmGo2QF9J0kZcyGvGXjWgYNoMiYiQDyVnBY57b9r+PFAs
dtFgnZYowNHU9qZn7jqQhjVwZBrj/s9EOZ9gg2c2jLhlTzAm1etBltZkf7X0rbEXwUdeZi55wOCw
x4v0SFn0Ixy+zYkwvw6k4W41+skqgqG4X6AB4xlz+gFqHkbQAlushjVOZxtiCvB9bP/hvGvBCEeJ
/STTVuRyMIkx1g5vL+ffsRJrPnIZHadqgj1Ywbpnu+X5JnUtOGQQHbSvudf+A2uN1GmGwWTnJhLE
lMqXWrOO3bRWZVMj33KSwSDileXEOwI1y7aiZY2pZhrTNjE3xTG/x3t/w6/hh77qwiP0xRRLVqtp
OZsUukA0nZ8jjR6NQyZATU6LxWoqw9ssm0nXXED8z6q6xj/m6c3psLVm9diXrni2IhupmtirqSSz
H9XFc/H/wqbmLHuBynfDhrx9Amzqvbvh8m4W8ieIMn46SKL3Daw1mure/R7T96n/xhpOg5CDDgZh
WF0u8v+T4Luou02RAtZZkamPuGs5Qli1pZw3ytaIse/55Tvb3TeFy6KDyj4WRObBBGADu7Y4alPV
fsFxCalX86EUq/uzFf1wYtS40LwxvqQ3fcAZTxJ03V/qWn5MqAF2QtwFb8gpEegN0GRoyQSqXT+2
ufRy23b+C27roqI9zoG8I53dLOy+a8RfxGp5MmI9GcRpT0f5MxNUp90X8Wz9o/SM2yny3YiplL0h
KM4wWsR0h8P6SGCKTBOg8zms+MHait2l9mC2aMbPvrflcVyf8qpq1h1ZrEzBqq/K8eeHqUxcdUkP
ZUs0jYXrifd+XSDG2BJNyw66eGXQO2OJKAiI7YCYC3T49O+m3Gn0dyethVHxanpVu0X1TEXmljpc
mzilPRGZjhxmDXROvr1lIfsXHc5fJgf544cQT38VdhK3khgHUmOttaT6hdNKd3tSMShCmHPTj96F
TQS2BnNl7ANIEXacmKt69MHFBt6OioijRCXwAkiaTfj1u+KGAtcLXMuiCjGzrv9m0Ne3IneYmxua
fO4UozFGF3jznwEOzFtebKtp8Y0EKw9XTt5hQRJrqQjW4ug+GmTQ4USbVmEkKDN0bFnhcylJl5ne
IJXbJBuU8au2LmMN2EhqPFrF4J4LG+xKPSN5XkaDOOvGZAWQQIf0BIS/zao795ppjsMnnN9Chj3f
ABF3tJz/whQDktGerZhB32kIUkInTREbfIRKB77Ll0QL89r95hviefqIDKVjvcMpt0lfZ3CSqoEV
CobBHUvCWQoFLsrMn5ou3VYHEcahRf0657BkttsxycEXrbNOsNqwO5f++fZmKA+mLmLnSANaqX1b
tlmDGa81d+d8eNbNBjL0nlPX+KCVYQF4ovnZ7aosCkb4YpCvn2OBJVxVv1CCrw0qyHZJIiLKFRfe
aG9VSL/6T2p0tTpIlCPpyZ7+e2CzFr/M9zmLbQe4zgkFsUdGKT7YjZ/eWl3ikE3yN/tEWA/mGEph
ANs++s0jWmbectACwreO+JzqF0rOGFqJajgqxLDve9oY8QO52P+GsYqXtOcwccc4wzmMq2ZNz/Rp
reLWWDJ6TPWSwQ8HVBVM7ewgwYhcVXSZb75z2U8GjeEXL+pE5tMfLzS3V6JYxCsT4rG/ieMkBunC
Z5g5FhOT7Dc9rsb8lBcghBZ5f5PWKYL8ibTwQY23BysubRcav3SxIwAwozI+Znq1pSKaxaPA0NBJ
7Lak+zBNHgENfeB/oqShvdrBCnshy8v7LfDnN+LBdjI6Kki12MFp5YJYQZV4Re1WcCr/+sPEuRH3
a4GcIYUgj6JYEEvQDSuwk0lcil0LYqcgMOh1m2AbBrd2GyfT/ToBpAl5ML5TPiNBHQq0yyrRlaAW
0ycsTgCS5jUrFJL264oXoKxUIm1ko+C6Ey+lvzGGRnk6uROQ277uhy/9OpG+jleViWztHR/rjb+X
jxFLKoSDn2Y1GKjZTIc2/FpgZYnilzEPFmIduDPrXJwSNUSpRtLlHkcK+A1R9wtfcsbKRYQQoAuP
pq7q5s5AjdSns63bUK6H0vFHkOJ7rnuv0aqfUYIjw6fRXSVL0Rci1jRJssX+Yw4tF4aUH5s+TXe+
VfoifdGggA53CR8BWn8bCMIJTLRPi7kveY0sBooU5bhsh0kYk2UuT4c1ICOfo0jyFK71COU3nTrB
1eYUSeVUpdXQJb7a2BozvyNZRwFlGLiI44HcZKSkLr+3HIGRXkiMNIdxmC7E++/0NkyOBGd6/kpf
4f89ZCejHfF3Kk8W33OWVKrGeIzZwENIGek1e/zPLiPmiVUcUUa6DvHSD/5Av29lrvAzNe2z5jR5
bPISX9chYadFrYMfjLnPCvIIXxF510Y3bqayWDyZfxlRGnelvzhnMdqCuUL2640i4RXaGfspavlF
G4y0k3QqfQa9j49fPmvvuh8KTAh7g48B8Rj6Lc93kVLjoBwYeA4WxZT8XrwoP3WXyDpjQFL8lK+k
TdllkKmIyP+kagqPl6v/B10bqfjK1ukyo/Al7tDzrkNlbb8pXIlQUNvEYq6BU/nNRXmCao6h8zKX
avlLPRX/NMHK/YTfSn32tDwotAn/G6/sa5BuOw4TmrfWCkH/uYCpAoGDmcQ4j7YDTBFOXT4SMwZm
QgDPsFX0jve32049HfMSN0PjwEE2HCuKm0CPCDbkd/swC4NVx+reBLGUGBpleGWdMIVJMDNn/bIZ
UjE2nvGNmBj/FYEZf4MvhG4S1+GhxcXvR224mmo9RnnBQnaFsb9AGTaM9dPcghddKYtpXgUNn3+a
ruHC6bon9/tIya8ibrHgl17xh4h1ZHRha72H9GugWwV1Tgo812jNiEqnvEr32kdhRGGOwSEGldg3
PblIeGp5pOZPRx1jMhZT+8wmN54fokKrAgk+ojVZukvXBK+44o+oIhqUx+1NF9uIU1yoWhZ5yFy8
8nyLkvNAldoSGLdTH3mh59WGMjh5zf98/9kRdfdNK5Z0Jg+0B8r9Jp8Hxg8IkCXyIYfszFXUIVGR
ZORoMfCpxLcZW1sTcujJT1H2PBAvoQO5dFVlLYGnz9zAp5WNMhpy2mymSSw0/2iRnlSSV0mcPPcu
hH18/K9jE1fUk173fEI/ZT2hfIKMUynIk0gOQCPqyzw0pWSf6mzGWS/PT+XgCCa1SCE22W+n8z5T
v899a1rWfE5pwr4GA+7UE9DI0bXHYlp1I7BZ/4M9D8sCHKRp9VKtUPoDcvdqo56ysxOZaW+wDoN9
SX+LQCEhAcnFQa5IAQa2Lx6ZvX+VLHVoc1R1XRWYtg6yFEg7mhdAmcImHyFUQ05xwmPvx5iEOVgY
3ZgDY3HEhPSSgmQHjbaC9EVpWrZyVrxYzIZHE98UrSfkyp5wHocHEFE5bM9rqFOMGJ9D/yu2rHd1
PVjxG8E3OjQzOtHfYwytcqCNvm2UWN57g8dkUwinyazlO21qzNWpG9q96N4NuUZaJuPZc6QZfYrR
UzC9EhCy3yD3jX6aefAcxZA8O+bMKNWxcOSHWyvQq35aM47p3imWNfA9/iLtlgq1yxiK6nJo5sxd
ebrPyCFxc6J2+i41+kGFr2b//Y7fK7YEyjiSi9JFAC2Ji4+NbJButcc7g2V7qO3FRZI9/8UWy+Pv
UWhGRNVKjbXqAFYhD4MnBk4uzvvAm7X6BV3vhcJCwYCRHIx7L5+xHJ2nSsWY6RHFHWx4LLlZ9HKR
nJNy4pN5MlGAGmggc7PsxCKPFiCtL8If9TbhX6klhDkn7hxl0SeThD44bLuoBl0VNh/PaWdZS7nM
eA65U1N/QI1g/GzI+H9ztLADDk5axJ7bY7z3q1aBAbhwwYuOzacYbkl/Qb0cGImR1SCgvkKcZkEH
eSNTKr3or+Pg67llMHolCVZX7pPZkkyc0ZfDb6wfzduLGGy1X/fo0mwcEPJvU7SuoM2KZ5E9mvl1
kkG/NSCup4is3123RC1VpLFNn61ijjcZFWXjCGxDb9Y9+wpw4or8lTU1NVl+qwsG37kFbKxFsiFn
pTU1RrMdgRAb+5vLOpr0v4ixVn7durbRSIgY0F5MXoir3ciZEe+C/W700GNB8uEc7Ovh7IPpDqzU
LjYEzh1IY9XFrIgK4OARL/SrObGnJv8GvCiVio2EPOGkKOlD8V8LD0sISEFDRcWZkdv2BNd4BT9U
ojcq/pHJVFuF+J/RgTJYurOXFybfqVVTMP22VMG3AVH3Vn2eG4YqaLhC3FzlqTH7JCitpPA1elcT
+aJell4HAgrc9D7udaoRL3OImodSWyzky46H5NsYG3WhNZE9blKZMcblTudBnr/YKmcqET8flQze
x1A2ELoGphPywDZUnhdiXHo4q1CBphkPoTguA7aBnd87BQQAV7E1fKSD+g2mmE94U57MCHaS+bY7
IHuCwSADQUPCCK6MAfzosDgdPcPCBzXxRtntt/Le3y0rQJ/+5fSxzo7XENvbf03ffNLF4//+X2Nc
rAJgIwDY3owgLPXr1FY/y0Eb/ONqfdTpdqN761UuYxa/5/a4btyVRM4z2IPRTG4lk1oDubA/VovR
Eu2YN1BadMnuAh0AS+MLqUEtEbwBMvl7AwrJWj3YD273SbARzHckNCogX0pSCeQlWmSfEv3Yy70l
Oi9rf2DO6DGlK5Mp+UB6CL4PinEaUAaMUYH9SacLfNltjP2WC+XTPEMp0Tpjs/gAxIW0ZGlWRZS9
8eNSAlytywwEggX4k4/LdCB7vOciIU/hpB1PCLVgvNFVDP+yLuYYbLysJUE5FQ3hF7O98VmYofM4
EZBIHyEVGerEQ1ta2Srlob+oqYwCADGgmzZBbRXsEqJBthduftG13M0oIW/cEPmyZ9lMeNendhCd
Fc7QWqfytG7wmBkAhyBoNezCpAfxp0ukIrPYDCkWSlhgcWQJFKahE96h23pDncgQTukywB/ARuKS
k88Iq+ZZXJHTquWGQBMnpaSprPOhL4Ff+ycoIkJHXz8EEYLRsJX6vhgcIJLhBI0mGHFi/4JlK/Zi
ddRV+vMsQaQIHAWbrFLWWni7zdHYYCDyIP2OLsXWZncakcpAsU/Uez42KSuCZ40TKAKu6lVmFpBZ
TrGfirLP2UkDx9WhVbhPfX4LPZGpaGF/OTp8g6emK7DC3ElyqR1LXL+CJbQJKnuPR2UfmcobUjzl
lYu0LRatxgLsgkpxP3hYZQWdpDYXIJdhzMFMhNS79oQR7JT8SafhzupikEYByo99GfLN0twAMIZf
ebRp0B8anlcM3qaSkd5mEz0ZJpsOWfT45JuCxiWTDm5AK0SEgzNxA1FTk3ckljTUDEOQWH14Yuwd
FeYx16OTOexswfmPIXkLDBvXmxb4pPLbkH52N2PxunsswCRm/5QSIzLenn89qHCk1C2HwtfJMpxg
i0YStKZJ4EaTuqLRsXsCf28cy1wM23RfrICGBkcfz2ZHYVzPYH2tHzObZDHrMj1ZJ7jUp1GvnzIJ
wJzP9N7XjWTTNBOk6hmON1pYIXuQiLIHNfFF3ON+HWIUT7kATTdSH9D0+hqPMfRbhjljZD919QDl
zMR930Ts9ZoyjYpydbp8aG/1FQCpfqWpMUbdOmnomlW4Up5n8A+VLOf86SUFq3agIhzTsUQpCVr3
KRN+urQ+942S2sIsmIZa+LV9Pj8v4cAFYZQHh0yxDD/whgA+AVogZYs6ScZqsbcpOyxpE+nSRnFe
dBY1AdyD/lLta8k3PFPNK/pWJygf3OJKlma4r1RGYXlydUavHYYoIVCD3JHsUe8cFHDIF80bWH7v
wVm2BU4fS1jKeMW4KZD3zeujmjnVSSUmlhugc4c6UqgO0sT+EqwoA7gyNasp+3bAXSOeLrLzUcEv
aXckW0zKWy14pVXWJ/1M8SZ+0xQx+BJf8+xkvUwYFhcphL1WCtMMHGkHFTLZp+0S2pu2cwckWprH
SV2rMdCFNhRhfyjLqLA8J6mlCod13tB1DbKWnL0dpWI2H2FGG2aJ91qeVra7LlsDp7Bs4NOU4nPO
dsBGoQtUboDsRRZvupMUtEG/Im1My1l49ZqyBpO3nW2Jxh18g0GO7+e/FbDbALBPHze9r2CfnND4
Ffslu6HIAkFzIddtcMhR1j2wN+PAFgb25LQZ3V2VHQeLFjOEKHf5rxUfYDiOAwhF7OXhoWlMuU27
x7zSTf6j9wGsoruf3mIfPqFE0YhIfxmCqIQY3eEYSzdIaxPac1OMka7Qg9M2fKIlglNZ8PPFUAn5
uUFwrRsYtqxCXRzY5saB1Em73JIH7LkPS8wn/7DTUSBXsshjLSMkc6lfj43KufrVtL9b94rmLU3F
YWhDMLvUJlvpOLDUNWOw60EfyDc7tnAG5y6WsqN/V/KyyS2JsPpLRxO6vlA5ToPIVBKent3fM2mP
K26Pz9/kUVXwNkEZ9JMfzYqjJ13buo7FCl0LoX0OQAHfqpWPRwvrbI7asIOhw7Lld85M+imiD8wg
/ACg7uFCrEYGyK5Rf4Sft4jsaFrJMzUce/LojHqYiN2Qc2b8MqVD8vslZXCNz85hfqMBKmb2UHL+
O4xn436b7EOYL9NcONDJgPtT0ucjCv5FmlZoA+lYepiQRaEI5h+E8cRSkmL+GTIczMMSY/clfa9Q
2UYFjDXK25WPjKLi+Jmp1BNUjIevsV5AZ+4dqWIzwRAak0tPgdJsbnTWTRCy08ts6I/ksPcn3uPO
TB+ddJi1aKCMN+3An/L7ChoNuowXMi31cPBXuLwCrYuDXRDo+wRMR1LHeC53eqZgiMbbUn2pQcCB
JOCOVPYqS0YS2JiN/rLwlFQH6xUNYN+fuxjjmv2k4pOmTemmvonsGCcl1nRDihJq+pptI4Aa8kAh
gu3gjk8KCxReAJfqm911A+70aXj4zYqkbQx9rNjELMnwMMoSKJFU2DuSdmVg4FHpIROO3IpKpaYS
6PkueM0YJOIF6QGADeRJ+xwnnGrmaU+/Gd5rNvs7i7TTNPahQ8mU72Z3uqCjFSWa/au5nXE+libz
ZrePkXstZ88f5LimocvZb/PzsslMqs2ThYbLcIaXs1GCSvnljhboUa1AVX2Y/syFZCW7ntwNliyF
gpD7RKFnAx5KimuUygR3q/bZAO0tJQGYt7GUoYYnIrxeUPXaNF5o1B+b+Zqn6tk0aZ0fRBJ6ciTK
+0Xl86jBgFxX0kFRP7xDb9YBTrxvQ5V7TKH2O2CaLVXVJbTojSSsx1/wLE3JzD7qqadUbUGa2jR5
sY8WTbH7gO/PcmbIJ8es8llh0CGTlSeJ9loC9RG6ubxvrqU9l4Z4LywAx8c4z3pphJe/ybYjSDGs
825l11MRBKETT7WP263+c8DLqASGqKwlLkxpo/NHYTBeJGh0I4fkO7Os3lS9CtzcIHsGmZmnPbJt
FA6/yKFAoXDh6v0rosjokeQfoHgimAiFF63cE1yi/rchQ9eO9isBI59DZ5zNMk5CY/lOMIkk2pph
yNAZe0T6IfAKPv4YO/n3g8cOrxDuDfRdmFHIVncR/uDzfrk4rfH4F2ywx4UDcaS3OrFjw6Fmcx1l
PwgAEhzYLc60Ry3vqnKb8La6d2nZk1nBMtBCD+fy2mgbzzkbouVJA++1sGSrBehvxLe+bU7M5Krh
cptG+Di088XDSciahhxLLUVzdhzdg7qpZLwRhTnmjDm6B86DVVxqpQDFpfUmmmyZXfBTQNfaXiq7
LES4aJb9wnqxlCHzQ4+ggpZ64D9Jjkn5/orpZ6MQLMLYXUOTD4wl/Z8ZrroQrVvQfSh91kEfwDnI
uAfsIYQqwPTvK/qnHOxblKD1AkAUIEMfo0qPpSo5nZ+cpvsahffbCGIFnfcMiGYZuQp1JE+vMF8n
OxukitCFY6yXmRNrXW0/MfwW9uBvgHIhwhN3uvqGkOwKXNO25toC99e6YNCQ6MSTNV+h+F4CSqHs
rRnShKo9T3K/5P7tN1c2nK/PuQhkULbQX+4+aH7QpYgR/mxple5va9/4XoY1DLY2IPepZUwFZ9On
QhvL5nIHMwQx13HwHTSKNLpW85HlcF+rX0QiuxaexSz/wmSFO6pGQwo8yr4CezAt2pAghKCr7N28
7hl2YZwi4LaNfYLh0R+hfo2x+R9WoKwm4MCMRjEFjFxPM80X/40em43DcTrhT+DEPhwoe3AfPBtR
6DCSzMrquJFQ0eZ6uuoXChspeuk3+XisSRLEZTGQACLxanlAJwam+twF6cCdolGDidWsuTHBiIJS
2UH758s2klOrefydZzTVVOErhkay+xv/uoJVMW3tfGIOUem5S0auwWNRCoQbE0v8b9F03XWs2+71
ND8/ybqFWectz5BgymhGzsw5UC5K/W/VpiXiRXLVgw2o4+MllVFurm2W2j8pGAT7Ne47t66UD/Lr
lCvJe5Y96rDywXRkBdeP8PPsBl1VU6NZrkGudcTc51M1Ob22i8PPVxo+eKkz9GVpU8pAA6Ch8bAm
OlIkekJ/TitFGNLomnz68wfq6R6GdDdtvd0jpUFs2Tdk+MB+TVJ8KwaHc2iinnOtUpBpo6BwFIO4
pqADZJdwYG56QW515rm4gY6DwSaiZWa6LbWYJ4MgFQMRNXZXGY7KEAQTd+4VtvYAUCFZ6Yt06cBe
Iaji+kcKkYXOHnR64myStr4yWFmAKKJAu81KxSVCANDco3SE8qTJuqywwSys3PqPrWTDlXGhdrBV
7Fwo65I5ztQ4AlRvAZ93mZ86rimFqf2089vwXny+cEXji86TwjOQ0dMNHbTHznNlprJGxdCEmq/j
n82vDlgQIllHfq3FxvCCMnsvxPsaCO3d+VgX01NPMWt2s8/6DL7IOFc858GhFtV6Fmoq7OsoHw9k
OxB1PHuf7thzTO8toB7V1X8xafOZcM9tOlbaDJyYlB9ujd4lA6LM0qfkXWOz2V1v1dmyi02QuS6g
Wk3G8gjD+KJUMiWdCkGu3HHl/enoMwygGxpFkGSKm921TGfuO/2a0xOk6ur+mwf7palMwrJudj4K
pAus3JZBkVVT6fr2f2pqGPhyXn6KFxpKZ6vz+5RTtPOArE68HgUj6500Px9FrcGDIA5+efkVj3ML
K7WxidRJj0d0vbUwHfVaILr+nYXCVCPfkbNg1WZ+g1Egp8wwRxwUrum7YH2wGf7ovVkk8uw4zklI
sW3zqsTDkrZH2SHLqxhnODh5TqLJ2Dgg9Y01KutAvIYNZ008ixG3akOiyTtexWMbkzZV+Kb+ygsS
yoU23PNTNGd6PezJRIT/Tui8r8tuEZ/UNw2Zwc10Cu6P0lqZaflDiNXXe0eNoDZOk+rrCOPwGovp
oBTtvXpKHOIk8b+5zDC0zQnjyMLO/dpuv2MgPWoVlZTT60+p9duHkglXmfA9ODJS6MKakkrHue1w
bF0vRq5KOcpkvk+b7JZzGoNDVXGP9UqLxz8Hu9yzwSNVuh8kFPkgYM8gwoU/CG4sCwx8xKaZvjRJ
f0YBOH5gYXgsn00ZgLSjmnD98+fDwxSHLtVoZuTjbfciZ3Rm0g5qzC7Y31HMoinNMRY8Yy+TwMlw
L1woJA5HTtwT3C8ml8bWoRbFggxTqAAoHqWWNtHD/ozy1iXzbvjZ35w163UdNMSqh8NAFcTPnQI6
PqhBuo24nViK3ce+S95hgNQBIWCqVqvhIheR/ViUxWGcRTGPfvHMMS/9M+d9wIvH3TAspBo64tPX
Yi09cEOng2HOf+srxoEQQG2QzYCKb36MGmOMe8S9/opStqD9vLQbq0jHx91WqKCzKJ5UvQReYIdK
oZ6rTz9G7OiYBC38iiNsEFCiNP0xRaSqHZGf2DCXYfwuTiLMXrIFODsS9XpYmK6VvBEKp/uZpaAZ
saN4TZevzjR2FsgSUF2iawun15dApqFWkTnZJrbFo6XQCTPJwpzU2eT8eWctFSZDvsEdGsKr4Fne
oyzG2KFGNcZq6HkTsYSPLRIayJJPi1np/1mkup/U/JYng1bRB9+EZJ3A+HrtfoZQ0QzcQ27iz45f
U9rPBMiY3k2qBrqtCejDZRBV7sB4KsMXxvQKsc1dxst18TrbfnzSy6eNvnPUJk83jyCHL7FmsbqH
t/QTnnIgpGTNeQkY5+OEPP6hsOtIoTNbshR49z0+wsdI9XNZIF5FWQ1HHUrIz0JB3N7pe7t+5J42
QOoRLICFWMkJscCUTE7F8nRSBy8O0bG6TvDJ4sH1XF15/ng01q/znmImn57ULR6v4CCWKBpQTPfr
g3OxdotJ6LIYLDr9p+KXAE+fv5pmLB4ILOpxENpbmmrhcASL2x2LmucqXCzuMxC7wXRfoZY9d93O
vOc5/c4vE1mVPjv4S9lLrK1fWD4MhdbORDNO25hhpVtS9y6vFs5C8MR0zkFqbclnIJnFxuapmgHo
nuRlrJcVmZTqI7eqBVnFqpfZfmoYVBqo1UzWvT+enwjegsv1wH2/dRbk/9dQAzoVcpToFDkbFLnD
9rnxbp2YuxOY+ofwNx8cSz0RGt8fxLc1Oezb3NwqadgTDTfx/zMlE24/h1ofnb4whTfJurFy1Dkf
RW8eFAZGTWx9KAkT0LomsstQk/2Olc1MK3pA4S5Cv+xkOKmzFD/dkDLRR6LZ19v+BGyGcAXH2u1U
HxA8ey78/DaKF89QkcwSxgAxuADvWrnRJxaqXLT4K9y/3ARPOUZp+SLHr2CoA+JBML/uOieaYdGp
mOmkBMmcMsCFeIEW0lzN0DIWTyfQAXcC9z7/JdvYJC6UDoOD+XxKYn1egTinz3iOtk527PTD2zGU
+lAXGOzJkxcYOakha813FYvLqETLZj7STvQvb/5I6WRGgDn1AIdR6vQr3jI7FR6Kkwe7qmdbQNNF
15A+h+Nh9xuwURi4uxCNUELbUpyG8ZpaOJ0lzQS/v4uY/5lu7EQKmm24WxDnm68MdgHkx3TQ5SL4
FhEnAx72fvOrPMsNDssveRFNZrEIHlVSFHJzBGdJj5BkEq4x2aQ+LPfIrpomTQ858uPSwkFY5JX4
yaLE9uiQmdiyHQoh0gRcJcZjBm08Aw6j86jIISNySNI33dNQ4qYCMU8X3RyQJQ9BsfRCyC5EzQUr
U/S0Wb5V+Q5TIgj50l1Vx5NYbXkkQ66PHF1ror8OcfToTdaYfWwwmskViUENfkv3cdwq3YKz1rLl
+qI0FTr3X2u3UuapRMFJMxLM2v3RkqePPAyeI8EhxtDqlEesklcC3zfHWxbxFn4n+QWKNfDsKFGW
1n9+eBoOZA7xkNAKKasZ4UXaP485txz+0U2xMtiNXWPa//GoO6CFlfbBxmQcba/DGFU9Vp+OPHkW
AtmWDGhhNyMdxnrNpM2eFgnKlq8LfmujgbBZIwGXBoW0V7yddqSir97XH++S1FyIGRifbeDRp134
5ux/PxIpF5UaIU1AvlkTKlOSNraMNHNKN0t3xSFeCZSVa11G3eJo5b/Ya0u5S0BiGchue3hppG1S
gvSo1A1zEPfiDh4/naKvsQnq8YpzV9BlxEB6BhdCkrDfPvTHckv7vP6Cu8iePIsskRjSd+wATImg
9H+Vz68dFvQIYOhruNgiRyYl5lLPEHRoHTOQ0JnvVs1owV0jDL8ZiZzBe1VoYiB2ax0wDT2860hS
t0orBhG6ebHJxN12BNTKfmsONZ9IuQuchYNpNz8IgOo2tHpeogq0KgUhlPuSfMMqqeXt0kNErBlz
X3dU/XteLO5265nFFa3sgciIeWWepcRSj0/MKjQKOWAwYrJiPLVNOMvLfTQDJ8GVZsvUPjIByL2K
VAN0PqqHECAAApZouAgtu/M1qR0Y4U6LE2kp1+UKSlQ/azOqoKbpqrftleihmaHHoYO91fIQNXLN
3n/rX28v/TTXL8VyT37mJClBV+NUjCxTnJeA6tr63CSsqqZGgD9hwom8EjirgeyzqYzjIFpexc8k
COuHzjkD+oFz4aYyg6YPz32XN0uo8b8KpvSEXwvqGs+Df5Ni4jrzhShC/hSZo9JbEsMLSQddYNFM
7JuJjBzWcqpD05ehbFvm33y/jXLZ422w/XA8TVV1QPmZqzcYG9XYnphOlJ4/rO2JDolH7WGSXa3D
GsDmUqKlmTShmilN0lbMyQC82tZCBotRGjTJBhy8E01g8DwwyCP/HClVwS+PYjr8jbTv64HXWn3+
CxZ4xUafGNiUd+4uBncHAAJ+CtYtDN+ZUo31tj37/pTRgwhPCAgEd+Gx5Dbe83yB7hU0s2PCeOz+
i9rf3BgYyPLz9kaW95B6Elh4jI82EWWq737bbfXM6bMvuES0pwvSOLm6JObv4siYNLphJ53Kt2+/
e+rzgUTGp+n/Yxv8jtKhGcCCJKlUm63b1MrgxuYSP+WLD0qfQhi11QyhYWZen9hlh+r9SMxsNHmj
DzZHzNF2ukndSd0NSfnnBDKAD9UW8lJAywZMJwiQ7+bzeri5DjoN985HIROTmeYI7qAwGMHEdx/D
QCBNnC0IbuYNUYLXxrLhRB1Us6r0AI6Jnw0wfD/9ETg3ZC/J/8ejhrknSe4M2fVMWKx3zM9GFz9E
yUJvH5rlpzZwloguCJo0dnDG+0ESFDOcnhvGBaEg4Pd8oxlFImMbzn7UdqgfjB6YlTj74KzIy0By
slERdmB/l0GCeyypPiy8E9uMC/xI5ELl0/2pvNhqPYhebfjutRDrdKKkqeYA7YK8ABtSuVNnmRm3
FjmlL2NfUDPUE6qqBWRfWG08Ys0ed/W9AVNJURw2W+kWvbc54AY3P+MD0bRe9Nd2bdQFsYx1L67D
fV+j437iWkJFHoSYc3seuqCVJYznLOOJ7XOus9iSOluDDdsQpCpp3UvTmYwVzDUmuwBGUjXjj96D
q2GQfeLGlHoEFv9A8o6lkPoES1vXwnjHBqrBR/wCCBnbc/P5mgvzKEBLtipuv54JwRj3gM0whteE
HE7nI0aAzysU5Q3uLD6K20OXPOBx81TQ3MDGi/nYvDOuv2X+5v36i+jey9MsXTuP8iFO8hCNFuQX
BiDsezKaIgSL/Y2GGNVjzeWGI24qK/Hpm19eiGNvK7GOZ5uuKiPgXOyqnAsUfaT4Oea5CuhckUJo
JA4QOCEKfaYwdbRClUGNcX+qh4PzCBI/CkuPT4FtDFxlbesE8F7zGkvLEshLuIIRY7lFP30EHYbN
1CVbTtv85rpbC08qTgLWP72BvExpy9BO6FfhRHrcix9ogGQR/KkQrlNONYTTlOyXQeDmHW8V/gCq
KLzHQEdzwpouF/8KmR44Lw6N7IesgfyrUpY9dBhQ4f0VfcXgLC0xuGVvZqVmb7GJilG8LM2GwqqJ
g2xBvp9B90k9TKi8vuZhuWSsE7HvftHfz2GzhpyVoFwXN3uhRm4c3KnWmwvoC5GyavaqLt7se/Ef
7JBz8uH3NgBwdaKypP6QK3xPiCZ0EpPnz/DLfVBn0PifcAXqi+7Sf+i8BxZs579B+zNiwlXOetiP
eDHlzaBoe/k23SmixyS3wI93kzzewF7Orws8kFV0/ARpC9yG4TwfhN1W+fPYCNJpr7PT2XWsj5gO
JZIkf8wmp0wVnL2Lb/UA3yjuP/Q9/MWvQfkZV0LJUKmGV3rPRpgM0o8mDq4DTZJ4Z9fx7xchU8Rx
V9VC5+K3rlGma4ejjrg6dT9Wl3j82yV5oPdhWLAdFUI4B09I5CS2JcKO3qN+PmX+a6oFKPTswwqt
vogeEbCgus+KPh/XIK5VK6NYviatQT7dqJH0uDWooN+iM/2EVRld/eJWK+jm4eLhUgEOOCycrOu1
hBuKA/dChkOM9mwEMuimpQbdP0E13xdTXWaV82nC5XolHyZDrrzLXirSYkQexUhCj6Wgo9x9lCfA
45i8whHqZIJGPB2oDs1aPQ9koKFBX1LG5sekCK7DKiyYWj8uVW3OvzCkcuHsq6dZUKVh00Fw0rAO
kdpiexteWi+DWq/uNaNIVKpk5WoEZ4RmhVY37jcSNVUnpeByFopttIrByq71e32VPjcp/Yaf3oMB
AKyThNqWDXVBcBeagqy0ZZTCzgU2FwmfMYlELoFCSXnwZqsMgORYiwnaYQRdI55/jUETl9wwkSJo
JSfZieOMhZANC0w5FxRjWED3EEQA1ZfFTgkAKfGADF1kGxr7jas8rZ1Cp5mrLMHH45rl0ZiJNzdq
wW/YA6TEcieaJo9kcF/oQftkgk7tkh07uEUgLyJTLjmcXNSEtHT65hY9lk2r/QjWW/iVx0kQmTBB
K3XmAfhU6MDyx9zpULuuxNC9mlPfAXAYAspIPMF+p3mS1+fMOKrw+BYf4TgDvJprhDlzqnqf1mx7
vFdjX9Q9kYy3anmLDZ17h4Vsa8EcOZe0hXwPr/McUjVareu8miiXn0bTWT8K+x4i/6YpCyzp2fWa
QBVl1MPbbi9OiPgMAVLXEi4ElrijPt4X5Qj+LnksTjvGpt07hvky2S6HLlYb9uNAZ7ATbWd2SFmd
Pbijd9NOndY0e5g7TL+gLeJvJD5qUxvHkaSLcqhQJbCk8fY3ss1D07qvqSotTBaJRW4H6KdgNjoL
pwLNq4HZg+ju6BR3rzSLMih5xS2suEPixH6iX+81y55jDJgyNahZMWREpjPLelD3blRyFyuhpGBZ
U9h2m9g3WxhGvDSaiU7sZseVeu8wv/0zPaWF0BOGA7/GqciCfo4drO8oo7FYOgwvVIn+K260p7WV
d5Q83mhmyEnrAUPyoh9Es/LTF2Sy2jV1z3LW+DVzBXD218ILk+P18MfG3kus33ZDfERijE2rpKtM
eHy+mKmCyHUGKr5JN5BcVhmvaMx2k5mB8sP8EW5BXZotbVTgr4pa9mdAVbZgb5qQXFtN1DTuufz/
vpmXpbQf7KVoNSf0xDxQ9kU5NgbWCtESGBHaeRYH/R0r0t6IOV8ub9bfNkYw5junZDMDsqiqIMVe
CGpSJ24vF3V/fogKEG0b4ag0D7+gGCFNPGDMVtgOFntXeVH+AvjMP0tUNgwV0puiJInn5HBiHT+h
NmHsu7iuLCDKe+509wZeDyP3PjKMJqbmWMVxGZske04LMwyMwqrc0bq/0AQADgXnQVanxtiXFDxL
+tWQsfbq4yGKE/IfKd4h+ZUM/DzpKBj1D8Ts10gv7GoSC2un5kOVcC/jPDI/uYQPZ7+GbE8QYkt7
Y3lfLtC6PpPRlfstQiIVnvnnuhKz3sqzLopj9P80fB9W6kM4CCcsKfEJjidRk1kAwUhl93IwME3w
Xai8kYFeAx7iqNnpM8EhT6/hdIWr9UnKsFtwn/Z93ilwsEY33tdfcCeIrqVxi/gbZwtWOdJq74P4
EyFgme8EC9O9I6PgGaeK/lhZ0l3X28lmA2s+Bgqoc8LkOYq5FyyOBnrN+fOvcopNS17FC+e9pcsC
n33WjRnAkFtUIv4wlyhMRDqsRedGzb7aWYAw6lJmrP/K7fYAaqsYo/xWmV8+WjEGwEQLC57Y+x1y
PQA3OG2YTpdfZyzUKvXtyiYsc+PFPbtzgdMjVua/78PTROELyDkqRzX1loJGqN6sT9WnKFUjc3Zw
JPoTB+mDMiE+YfblhVnVz89MpnGKnq6u1y1P5sbhygmRnjaLIVoX+EPya2MxwfZNShZQ5fvgJLf2
mtTVHGTiHKIERsZZ4Cilc5M4RQjtqst+exXCrHULoVeXxxlniioa3U1ksjhxdORQ6tacXpVidGQ8
IBUQV7/gXVOvsTZRJOGM1pt+1Amt4xkm8QfFrfMpnKuybH0EkrzVhjUah7r40tSjxcpAfQKhF+iA
+IiLyftmo9t+oF/Dy9eSzIYf7F7bhAZChgminf1VfJ1FHw1gMsPh1Y2k/gvCOWtmL7UReDs3J7og
zTTI2yjxoUYBUZyU2PvO59nmkJlyiUSv7QeSNRO1k0Xa2soq+A1tD7k/Q4J3vPyeO983UPNuQsHQ
hJCTNoDjdGp3VLLDN3bNrAbUv5k1yFHD+TwJVU621aajJCrub8BfBGSZwg3aAdh1+haRKLCBseP5
AAtithOfc+0plKpm6WTj/72vh5+3y4Av7810kKgzya5ZItplnJmXUdB6oHlWU+l6K5FnG/959tMj
TYn2J66T1ni1pbVtXdunnNS+esAoRmfy1yQknGis7nqEOBGp1EwG8aJIgpyhQrmchtz1HZnVwUfv
TVrXrqhEnah83hzzvgQCPKC4FOCzqffvN51LxnF9AhDZhl2LlqB9/d7wMvxTDfLBZm5AIRfUbMZ2
IXh1gH30I44v8dRiJFjOr6NiQJWdoNyPYFPwsbYALoH0eAhZmY56Wrb1gCjGkHyKRJkwOsQDdjI2
Tdfy4eRG3IzoE6HW6F9dDbYOoSa7sj3aj8bI0dRwA8J+t6D2/drpYtX5TFREnBxUD1tFnEPyS1MY
39XSrbz2aFbNg7wzPUcziNtWtcqjk45r4GHml6tHlbUEWDLniys0FltaOkX1uxWJVMHl32Br84nX
IVid2rzG/RoosfS33w94f/jChjIvYMXM1mJr1vPhlhjn64pEBWglZHBVYnd248jf5Yl5nYYoqRQc
p4hS8sH43j3RzbgjHZH35U1xcLwiznNFcx68C/GXv5ZOQYkc8H6E78GPICWFisRiWhawXKtomqcK
OvpFdh24PQn+uuytkm6XdXtZ8+5MHeN+1Qrxogz45tm3BYPJ73SyGZj2Tj/mJ0foD6zg9asU9pNk
dMZbI9Eb8AtF5quEf947hu99S8RcDqu1uaqMgv8yogb5gX0doJQ5iIJNLnAiESWg1SMQos8Bsn4D
NM5fwPTkvDcFsxuBjSYkeqthiBYTAl+/6kO7D7FLZy6+1sj+2rPipvewVI30QjU4qZ/sO4IeUrHN
SKjYEZBP6APVmVNFj3a3mzwTzMhZ00yleT9zjXjX84t+QqprMAceLXMyJdTXuFsdWEiTAEyiYEFE
vHrwXx1Pg3xi9CLIphofsQEX+VavDu4pFqtdo71BnYec1C9uEFRK8olYfP72LYw3ozC8lRyRKrXT
6V2WURBae/Vt7D5li3cs9wSoVjakhnFmyCl9AHfq+uZzD0vCpUO/RmVd552dUNgwpJlV5/VuSDDQ
3ESKXaeoCbKgRD1GuqfgpqrsCkAyYQNdP/haxnJ83LsgQdOxdwzJufyfVOlUG8P1XOOxiqHY4QUU
3IhZ/itdco483WobXeY2rn7cO+dfggIG4qzDMVfKDGP6veWUNw2GarT5r98YnSa8S9Z+GEnm7p+r
TciXugmp532MpBXyy09f8aQxIqvxDlEQr0Zm2dhembBh+mleY7t/EKESC0X5sWnpQ5KNFrr9/Aqg
vDeB7EwBETYyzHYDFCo1GqCL7vtMJySTnv+t3NuEgkAwJtlvTGbZDMeFmCfqBiDe875pw94jN1M8
Lp9DRej0D5xQJMa0z2ggs9Cz/W8mL6zoQjvJBqHqpl9apmsiaHpLQ3n+5ROy/SVvJ2s3tbjGpklp
I639xvGx47rHpXg2TyZjjIt+cIn80AyjzRLvaVuEk+2OH64tExYb17cRsC1HWRrOxJzRQfTl1cqh
xZZoLRa0xIos8ZYgPyE0+xDdBfGH8Dx2YMxGJw3d+t68X640ULhqFa2iJoFovQ3WF/9g6eFTK4Ka
TstYaGTDhZeMgjgzy+lBvuJtpyhXkfIrbY0eGytOEWjJVlUDDJvHvD+JJzyhcBDdCTL+bGHREkT4
KfnlcHsde4KuuQYFmUexz/Hgs1hzKDF6xJlhM+5nXG574x/Th6fe3J3ntGIyp339FVEkQKAXRh0c
2FwVMNHV9fje2IOKsaNKDV6djtYzlkZzzrpREdsrqRpOfn210KUVlW0lwGGOVqGaFK3pHrj3W42E
kRmhvpP8VpHOSK71osiHEFBQDMi9QYI2VqI7qoQeQWdjoAGJFNmuifJRxPwapmPK+8HX0HSA2RgM
955p/dRM9hb6d9nd00BG6fi/72rCppgpr1K39iO8QvDgLFVfzBnzb4qw4T9KjzyPgfKiDA7BwWGl
E+tR0niHuwtGDiaJA3KC9y79hOspDbFA5LzLZEFav28UFmQkJx3rmyZwOWgyvrFDoXpElqLelv6o
wsodK8P9Z+VGknVIeO3XziL8rIIs+kSfdGDWBNV79VZXSWb0xjuzRXGQkFmQ7FHXq7QCLeIC+bhY
4Z5/3Th8GZzNJoKPKBB8Opp30IrN1VBD8IBjUdhJTYZmt1tUpS0ek7MqunJf1HVukm1v3gacEttu
pQOFglaToCyJY1DBcusvoyb7JY/tLY5W0zEBc6TJTxLBTYW2o43uq5Gj0IMMNXQF0rxTwrj3EvWe
+J3LqKg1AN6f3CQSg0uhnKsgbKfMFx36w5XqIZzuW5OU+qgRtI3b6nYf1pscQ7v2c579Xz1U2do7
z63j4nRNgqHOpHSa0zF7InDOmZvXurRPnb9XDtqYaXiEv2lMOR9EXimy3EY9zfan+aGm399PB4jn
PEf16Hix3K0ntN/ptNLKXxt1uy0yqRl12gVAP2OfrgftIQMYZLlegSTa8eBtlWniXnJiuyte/b/H
dgoHUFtLcsa49IOWF5qoefoC0atyp0GxGIYzch3vlBS08ZGqYp46/scLdMZkF6KAJ+6Xpn8i0IJp
a8RJMSf87MubAx6iOyljzii5vhbwyhwZdlPCp0qOG6iyyVCSkRLjEApBF28XRXJ3zNbbE9pjmESf
T3RqhIJbVZYwPnSZ9J7cpo0sj6bBjZeKuIm/1WXvWCw60s1DRpiiXrXZPsjqpOxGSoyCCJ7W47u6
IXZ7kZSmwsRBL5bw46cY0Of4gfnkEo0DXjNChNZ3LTm2A9vW62ADTH59JSGGIOwUf5bQ5CyD8uOL
dOT+uiOL27gOMqyiV8KXOzvXTnE8VG096t30hcnU7PvxjQhfsHkcb1FcIrT+tOU0SIq54auMYU2X
lSCsq27MqC3ccd6l04qClobVuAC45UmHL+Ba6fgK6a7Dps5DOeP7Khm4QlnHKStljTWCr8ZfYrtJ
3YfPwPc2IzcjkyOOF9RcZv+mQofoQTD8aSihmlSTpqcv7vTUBEUOPxSWlix7bhC/PX9LKmrp6a9p
ph62c7wwMSWah+Bl4lxbaE7IpWK0qoGF1MnZskrp7VB4Yssul4vk/jJH8AiDyngopSXYrcZbUcp1
A5FyaQJQGJUJi0KCHL4KxDR3G36GKOnkcFYJozY9FS+sOzUitvk1sVLgMCazz+GlHPdvETIRKu6k
k+c6J9NBAVtLY3cZ/kiOiKtvei0Wvkaon3FSC+62NU1jHQQG7Mw+85aTEcSgV56Sr3clAaytQIRS
gioeT7B+lvjMZKfQInRt9IZPDdOyPqNTnW7ExCGbLskqojCZa3Ll7VBP7yhzdWiNQ5HJrRUAj+bX
VdLFyoGujHrR4qPskOYXYD1ezhVWuAekGcTIb+Dq6fGvWjsJWkQa54qMwQA2R9hTGATbzB5Cdat9
yGy+oS4bugVZqU13Yn7w3mHwaNC+jtaOJJzSKKMLuyANDQQqZC8mXh/jE5ubrwonPVTNeQf70EvD
vRj2zl+CrsvqkP0qA1p3SIFv8FSZ9PzGQYSaohpEX/UaXv2H0r5sGFzIn6GwoPtC/+TUY6rI/aQ0
mx/VS/s9ApdJc72j0pmVo9esQtaUG5Gk2WC7bJceoi5go0rHqn4y7dm/qPs3k+/UJDXoP3lCLsbh
RAb35ptGE37pXvXeA8K+iwiERcmWRX4MwSOxwr133vVHzRw47qeqchc5a5Pdl97Gur9cfL3icIhE
b7sfaz1itBa3KF/gD++rssCPeFt8eCN7m+yMUdK90MMWyh3eSSt4xi1d5Y7HaFCwEy+jTLVW4vHx
bmijg9yxGIX2uFaIfi+OFwRannaY1SwXsz2Nd72J/tgt/Rla8MGhFzaFzHVaL8nNZBwQuqQtfy+X
6Ug1cnCWiS9WNlA5nxJ5e+yWfSWVpwwOIsC9bGk5gLJvOzYIhUWpv1IB+o0i9m9dP+vRasF7CYVF
ZidEFEaMulu9Ka8p4dNnb2KCf1Qcz5gKkz9Xsc69Rjf4LgNvtl/6HkPxGcQ1/BeRkmxaBmqE8PnS
aSBpArLm9wTEebwRcb4LuSHg7yVK+LAG5BVyttQXk97m8Dbitg4IwD0QlKUHbKs5hMrpq0BlnKwo
XLWe/06lV6lt5+ruFcmd3pxh3GueOKgHV6TXaGZvxbfmZygMUENj76Z6Fy77NSStMAKs0p9EnCWo
Gfk7PLN8DPVe/qTL0RHyJP+uooxv1M95mLX9kUZ/AmZ+jOMBYcYmA5DMk/WNAAeHrhn2f5aetajv
n86g7gYBbo20z8BGFY/J6/PvXYLPwQImkv666MVpVIrpkbmUR8aYPxa27hknDtUnAhrK7Ck3+ast
ANhAEcfSKn2OvmtbsLPnKxhWUF9ydAW1esuN0dHGkYxsAqeF5tQHs/h78//jJVg+zIslYZfkrrdi
SwUbuPvBGNdKq2YRQDBEV+cPOeHb2u4n8B4HNH4zx4DUw/+ADYSkQRwDAYRYhIO1NLWb6sxgU671
ZBImpetVPsj3XZrhOlPdIrhPF7dApjK1MLfqoKmJlJiD5w8O0Eo0T7Wk7CXJkrBTs7PPq85s2Ejc
uv5McRXdw0X48bApz1knBZOvXXwNuvtJYMImkXUvvP5U7BrRyLDquIgHVO8HzC133dMrGqK4kRBi
b4lqqfMnAp9uT9Y2TD/n8tH8f/pLuR6gQZ+5orgaMvfywDo4v19IiNlYzTzMlPhZjaarpJqj6jT1
ITs6fVGke0tJpyrAAEbh65e1rDDuG1h3yW3DUYzcB9oqKacnJRnzYAAhB/Yi8XkPb7ul++IjV89R
YJDldrZt9XINqFXO12jf6cnktMvWviYj43DV6nElNU1XGzBYoB1wIIpumdI6bAvultR8mJNyPgJ+
YdnV04EqGlRolYKbLmDhkSUUXegG/umIrMZ1LRd+GqS5T2xe/eWHfu2qPc37/r08lW9borhCqWZe
LVassf4azN/5DmDIB6e+nLSo9/X1qnyzcr2Xet9RXzFDJydUcAvkbqwNJ9P79hz/mSUCudmEoOT9
FpdwwVdDO4To4IpU9GMBZIxKC+wMvweuJGnMWlQGYg3RRn1gd+qKlxUE4hBlIkc2gySPt62RkuQl
lkxyuJDjsKGN0rEX7mj6h2mDxWqRSzoPyaoUaxcICszVgFGcL3qMlegnG+2JTuQXh+zV5308Z3SL
pSmTyO60JqRsbBfpFwoBVYrv7zdtoKINjGArjU8LUWCt1QTUMtt8TROeoWa7Auj4cOcrxs4keFNF
2txWQrdu3/wbaaQ+dV09XK3VCxekE810yR+d2zrKLIzXhf4AQPw+y3FWm5xRVcLPDSoSDlTbn1Yr
ixSQb7K9aZPNtDOqdTYrjG9R2GLtr8g/qmPHnfsmZWsyq0CbiPPNDdgJx1NYrfuY8uANE44RGR7e
fKqbdd8SdAP1oRCDkU3H4nxm0ohWo+8WOmlWaZHPrWapQffWOjvdzc0sHxP2Yyqu96+b2y8VHjC7
Bv9YjipJuMCnJUooc8/81e4TW4i1mAEu5TbKgVX8U8Nipz+86H/ygMoE5JPBkuEHUQrN1I6y81zn
1QYEnjiPQDpO02Rw/y5slJQp964k2WpcaRvC0Rv1umnM6v+fDCqj8DmEO206v3YOK/NVp+YNsivu
lVn6d3Gx+cR8L/Kmi2O0PvJfcnX+6Xtjp+E2vqycFqgfOlCSnZxAU/P51GI9x2Frsq7LmIyXIOzL
9kBGuqS/MWeeueKQk71pPy46sy/adGhYigFoBpOqv3EeAGqx7Y0GqJrike6ZsGJ6OtRwUWh6zDMp
0EjXVXIF7kJ1Utb5YdjLooxX6tWHR2++1zyi9AtSyOXAG8cUnjk38eOxz93Dia+CRPGdZznxhuq0
/wRA8p/5MwTgeruzNYVdExdz7dnZVu6SNa4KIkUgqQcpq7MaTPnwp/xSq6ZzJ22UlxsbxZY4HGCY
skDYPTdZ6gEM3vUgxaTpuWEUPRVORAk3lM5U7Zek+HlblyjIJNboBbmICLH2SV0w5tkvjS6F4jsk
IGjss1YJ5M0JC/ecgzQ7bLX5qbDDy2vUIFzHykgoM8G0H5ubpuoogI0eaIhTq495ql1hYy4D9Xjx
4StStLMVqllmNfyG6lynFEtTt7ojgV39XtsqKcPTz8lNkRghI/c1VkQ3+j/lCCtrm44eMe2omhzL
KRSLppaXuFoJmsCtd2sPlhUo60fJc0GaBA0mKVZp9/bY5tFZsta0sdd9PLYUmq/dmWKSpWwua9a0
x0j7jNxcr1YLqOhrvy8rMeMQtzC/pCysIUYkGZrN86f1N0OD1ZLZgO96Yw4utr+9hkEQCqhS4JoI
t96udXp7eJQVROeWnQzTmYQFZ67CasuJnLbDeie9Ts2QWuHC3PovAbX/+FM8QWLb4JFtX0CWMHQ9
JPZgZthjr+K8PbcO4ZndKJAHgCEFAnPKxQj18Xy/OQnOvE1j4F3Ts7Z8cngsMTsJUNOKrWO/M8nE
UuVlr1x0t8runi88d55M0KOcpb2UgYJOhHkV4xFr5BEEdXdA3z+EJTR6Rq2zf0xa0BLg5X6b5w9y
gMptqmNKvYbjFXiP/pcpzwJJmZJkgpu9LcmXRTYs6hkSP88utdiFcj5VYWCgwNVPleViUksM7jkC
yCt4wT61urKPL60cETM4HTVWX2bYhOC8cBopodMmdZfl8pYU8WQLOmEjIuvv7bTtW4HCuHLB1M9U
6Wpi1CmUrYg0X96Pz1MR43eDeetQfcro5d2HJxpYdGzSvC9M8r2NydsDEGHSPSLfaD1upYksbPnF
Oxn7EVdTNfNmKBJL8i3/U7KAPOWh6EHH0OmZiC3pfKnudoftxPMT76NU1kegYHJsQjWOh/Ek81o0
PteayrG9vVSP0NS5GJLXrVsnIRzrwYwg1+G3lJI78ChBfDlQ3461+yPkqiH5C96hVP1cqz1zc6Hq
XgPI0lRfaliOWBifE1UKfGUMu+Nz4kCb12nzwfVWSPIG9JT/z2NnXIgoIxBmxmVSMyVR7fKvlnG+
Ov/X9i8BAY1GJOFwEces7UyJW8EWfDZ1ug7hoq5xZ2X+xSSWcB4Em1cThMYS2APn0ZT+2wbhYwBJ
vjx7M45S6gB7JZf0c8ogW3cDPpd/RjrIaVRoFd3O6WZ4Be/RGJE0n5Z5v1st18wVj+aYS6N6plT7
cKMNXE9GM3PnlvwfKZqXEgX79EI7VGhfg479iJBQWbkcxgACdQycXcBvyWET4ELUZSm/hDL7Hu6I
knQ4Yy7pMf7/YUIwu29UdUGNd9mNFKFp3MVn82T5Nm9l6eGbLAo5/KYntYGMhXGmeudV/wGTYha5
dIPWDYws+FR0RFAnvA7Lp/bRHExZtnf46x4HjNUYcdvYkTAejKquWLj3/a3eLRuVQ7wM1WBsyo4U
uobTx70hSkkjpZ7Uoez+pHjmC6vSZ90C6BgraGmT9hbTyom12ejAhGJDx2wvbB44ZiaimghX4mpc
oWm1q8R13dIcvxkWH+cQhoIs0Vr+IJ48WiHOXZUAB3Hwvh808sHnDMB/c4AqQj4tkoNFyiWzrpn1
lrWHC1iLEz/2FLenmfPR2zf9t5aA9u1VlYkM09DCj4KVSb/L2A01I7SWwC5BGYPNkPhAPxP7YDfL
sXBBvDJp8ixb5sx8qEDdKBXarR7AiAxT+ME4lMx9E+Pe/7k3cW4cx/qscftqPYfiWTqtHoVX8b5h
Od5HKLkyCsafey07Fmhv8IVeMztVl0ZN2yxfMHCRRPdc2CXJtm5PCc/r1Kww9Gw+vrs/03wVNNe+
i0f7p+jggDq9VonP/rmZRcI82QR96bmiT4EuHbC4S2bPVICgXBrGraj/DlJ27k526AUb2/KLKIqU
FouYSqkR5IBwd/wjrP4KJff47KWSMKOD7R0wg/Qoksz3j7ryjeLcplK+Q/tlFWIaAK3RuwOH/+vF
T/sI4ahXsk5ig0jogUrYhYVH7mBnycNfW9VplVN/HiOmjmlvkFjLzoksYtzveebwlW9i0on9Tfm3
rCZdWDCDPX/xGUtg82qgmFboKYPcrclsPxSXLafEun+Z2frtbLmRiqis5qOT1qfYCQfUKU6JY6gy
0DvNsJncZPuKT6DsPOxqgQ23PNp8tI5x7hCWokpv2dHTDl8ryv6W7NhAxUorIJoY4JlFDd1MbYGe
7SXbCGM3ApPJxS5p5O3sfTQ3Xhu3TnU5h+8Ne6etNv5IXp64aQdHDf8N2c20eUakmMoUM4rB2vjs
IFb1p8kgAE28oYk/7o5qCVYwZ1kYDzmbEc6H4N8/k1jxDs2b77N1s/NIxpNAckLo5oecltc7tKNJ
AkLq1QW/jnhQQqaoydqlaLH9Y+X2mkr7/unYDIhAFoj3ez/pRebJjfbbCSxDS638JzUN05/HUmnn
H7QT1TovcKM2vCeo9whdEm332kXH3dve+5nFZeAFq8WwhDPD3zVCGygpBBe9YA4b6lx4yz5Ozlj5
jNoEPUliu3a3VAk2/hlbBgGV+CLy4IdPTDufVftyQ6dB8PEIEflfoHLVmv3BainXMaHQNFWeiMCA
cksag+UMNVLb/UgWLFKPBg9X38GKm8lVXF0hYXINnNvyRtGZnO6O9wcUhlVzLKFac41OgBAEjfHv
51v3Lotc7ZdGwjILgsQ9Z5iMOUmlu010XvA7JcUHn8SRAxqiKxlcs7md1D7+b9xzINO/lV6M4sB8
GsMujGL+cN8Dz2ku9ZNIfJPZ6UuKUuFWZ7mtK9AtirxbWtz1kycT3+08qVTFFO/zADyAv/euLHf+
T6+foRa7dw7HsT5zeA2E6yu4YWpvyoYqndZB8GesLZIfcIPGd4yOjQ/RWeeYXW1tx6IPCM1dMCe4
YXisPrUfxbESc0fgnrOz6XWnF1WOSPUQVPfVuYz36220Gi17NXeFossywcfSdc0K9N9FGA9DsuW3
0oiOznXwDyxAKtr7THXcy/eTNh5s5MFYr8yd3TJ+AQy7zc8olU6qRdefyC2dS29Dg6DWG1q+1V8A
2o8qjPzr09UFFupceTgDBKKHkhI8hQ7A4H9RaTZv48oRxai2xrCp0xbvR8eQkL+GcwCaWzbp9J3M
+xObHK+xNckBL6cV377OS7RZCnXYe0HjJs131cEh6e1YPARbKJOwPLc9tDY/6IC55TwUPq45UgTQ
pHbEbQC9N0kchZ4E7HyU+y5cD85DThlVMKErdSVHf/ghwSv+KgZpl/8hDkde50QH3/ilE69y6yKZ
lg4j1dpgfJC1i2zUwTfKpi23KemMw1Rscf5n9n0o9i3TZRKMW9clFtnz67oDQYETumTbdQdv5P4U
r51uDI9mmGmYvNFp1M/xR6eq2CDZlv2yXjniSWRSk4W/QbNFWTmqOvFetxtQlwMgCXbRDW+Dc0X6
eB9yu41UP+BC3WesbKUWQRSZifOAjzHfadzUJbQGNbdXRuxasryUY8Te9Xkbzz/JApS51Ofbn6xd
pC6eL5D6mHnonJDV2wmBKy9gJfUfbyen1dkF8KIf64foGpguAZR0wkcjQJd7hwCVm3h8j+3U6BCr
k2ro2JcVV9cwTJGb0hNBoPY7uezGrfIA2TGUjA88s6nrgcZ/gcQF2+wFTzgUUEHKEH7EFW2X3Ay0
LSuD8dOVGTgOrJZHJjaStHPnRbs4GH4awI8jso7hGIy7XrWJfWKbtp6qX5Zf5vG60iXtZ7ZCYqnW
jsKU8rfYkkUUZ1sYsm8qiBfXKdmcOM2wb7rqkWkI1Zwf02seKjTzGNrMYYvfcW6qEIdeSiAjJqSu
UwoCS4cmTE0Tpd8HhZKJ2LGUrCMu4DQ0HtRy8/Sky3PJQZNL+LnhhSApCRMb8RfpT6YtVlRbB5ZJ
hOXdWG4bDO0FUmrOX7XgspDGM7YblC90YkGozsSEHtYvBz7vkTl/6R+CFfj7viWChfzf0jzftT/Q
EHijDg9KndpNTsIKpDUdkrc8oyGr1UK8qxU0oT1aNK1OQ3InZPIu/VTrXPdhYUNVj4VjyVG9poRE
JlEEozhYv+If84oeQOT2GN0uSqehEc6w/FVi7gKqSAuNPCfWQu+YaHAdYl9lJ1MXIlusSRvCskn1
BTWWAFwuhC1HEHufjPjWhFvip13Sr4m9eTaYSuhMSwkJpng4QNrg8uk1CP0B6l8DYmCg5MvXGDmv
nDCu0ed9iS2yvbw/FuVXFmw/eQC1HwBYGyau/HGe9VRrVUWJUJKuBKilN0Mepc9UuTC9tCJ34vw1
OaKb+18IDL0rlkla9qXnnCuCMyZuAiRTqiaWl44R/prEFA8q7b7LwcEdODN2x7NTGD+WqGGfh2hL
EkEie0tzX1j3KFeIoaUPvA8nJF3JUA/M/AYS9gslbVoM5yZadW67/PGLXAKn1ABC2gHD05gAYryI
IBKnJIHIZO+qk0kATLqoJK+AV/2ktuEqZVeAeqQBSKZ8nn1yzfXz1eSi1KNdt8FXo6KoLYcszWaa
Q423Pt2s/s8ETmv4tzOn03Esv6F/HBJuSBj4lbi4eiSqXA2g3akQpvu75QJ1ZT8WgH/31xDs3DpZ
6lh2/JRW0OHcpTIhWFQWo60PFMNqTcDFBhPLMqC+vKpx4Rc6MGEO4pLzjobclLG52IQbYb79QQWG
myn4Cs8v3r/M1B4bwoXvLuCZ9SsxD/vHG6NhqU5ArQBINPncYJAYpsDTozHSbk00diQrxoHRUCph
1hw5bqsNEkGkmJGji3kySmX5+Jw6JHx7U8yzJqp55s4+9hfBWuA03XHoCArcBvuUlfi060MN8tMb
0BcT8eICL2scKeKEokXzKWFLJOjYq7wRG9v9l85BQk2cuWbYf+y1YAQlgM/Q9stW3YejKYcfWdfb
xRLDDCAUR6hhvP+IVAhJYZmZ76E2qtQzuTMBZS0eVb99GI7CxnPs09LFv0vb1idoDJvlDqrI65n9
Akkb72VCFBb0kGjwRApKFYt5xXaUJBFWCH1yXHA9YiHWjJ6rt6BF6pw0lzUZxBGNcV6lYhrEgsmE
ySOoGvWIqQdCe+eoLFX9hkow1vB9QUSZyEJDwgC7PpMsxD8tBk41C8Z/Q/88msrDZIykZ2TZGse3
o5JSO4Q4cCMQj4y3mDne05g20NrPJ4oR/3bSAs/27HQmgwG1Azb/vRy7udDUeEFW9ciCYOwMOLXc
4StkddXJDMnZxNmD8NEukAyhsHsEhiywqGaJ94X2zRPvSluKXm35Adrcn8A2z1HKz9JUua12Kdi/
FRvfCoW+UDkDjtfdsW2ZodCsLha1ajAN+7Rn3bgf1LEIAMPe2Sb0X8vP1/ax2fUL4mwcFZimwPMN
yhwrylxEziXd2SpryA1p+oAG+F1YPhgmDl8MVF04GwXzSED8WkAVIpes0GBL1o8+Jxgx5hBbkSKG
709EDYWzAIK7SURvdRSnn7sWHf9OGrh3SHwt8C2UGEuI5lhRqx6DSYJCkRyLNjWNQm/SSI+zMZJR
htSR7rj4cJgsqRSqOpVc8jHjhKL+IHjld8j3rZdexX7r2qcs1fqz68fsrkWB7vXNEBT6HtqVz4rl
DYtEfDjyGlNPq+mQ6OOq0BB9A3F0UrGh82M/bs5q9NygEz44RrAXY+qvHEKj57GVjLo4o3iPK4XP
QOLJo274rct0k3xntM45C1A9U8qZWJNZB1Wd0mk0tq16lDXzEhlhlmaTmyVMEU+fHnid5EIBGFtu
kdrddWHazMr8q/UPc/89FMz8q5pwHRWak1dv028VmXbPxWoUQmip+7q+UwQmtB4c56vZwHLxslMP
+FuGc0k/MIzaPfP5XfR+vudXT+ZZlai8eHFk4xobIE5jzERTqVbPBivKI6zdW5AUMqImmGAM0vN3
XDy4da80dCt+85OdqhcBQ8Vggfbbt+JRmtBBBWNdbTcrBfzRPnFWk+acAQocjinFMZjcGT2RkFxZ
0BALxr9NFG3Qn+/yUHeUsyAAl0Q9ZiUo8og0CFFy86tffLAECJbbTBljKwwhoVNi2gW+IIf5jzW5
ZJamT31oM8weA8InC2+cj6PDsqHnYkbTLpScvjJq0z2tvLcGnA8vSkIhd/J4HOB4Pxnkzlxmtap4
haogYEU6VWP7dkHQa2m7LH39SnXLKixFT1qjHa8z14fqeTK4YBdhWLlvdPCjawm39bLh5e9pUmOw
XVpas0lMoodyC/XuG7DMKTUy2WMbGTVYixClNVEraiQCN5LwUsI40HmTc8KYjedgmfeyEH9HdQVg
v4O86xArsmAf9Rw0qFtC+PioGeieGo3s91wKnlI8G7b8QigfI5KCCLQ5mMQeC5qxBT7seUNF+Kt7
I7LvOkbwieyduaDWeodFyN/HTkSaDqM7SwrNXg2fuH455V3X97Gl+0n2AiceJJlGRpOJs/s2TDqy
oIKuzuyC3p5EYvp+pt7Brq2H2qYLDm65X50nygx3X5bVsg/MKtO1ELh358Zg/kIrB4urrVnkCb7E
sxVyf+tfc2xxD86p01tlt4vRyvkU5y/coeVq3G+ETFv3YdzaoPoM4TeVIwYWmbZ2HPzP44ZjmzGi
V6VqMgm/y8d8OKlSfWjqw3zHr9r/2pBrbT/j6VNKz3JF4aBUBlJcj5yLq5w+ajntR+X8e2kHC/MW
kMgMn1OYTXzKS/NKvsz6hUKDOGsQ28Eb2IgKT3GGbVLTZVsh/iO+JRbAD+LbL32Zpf8WOo93sw+l
zLsGwnjsz4opPOJfF36cdRNKgrEOXkQFErN2WWwKxmgbzjqHfMSYYpI+EgOOpsbK/j6FJkEaz1e2
8zZYG7G1w9XYL2GGHdhggVU5CcWRSgSzJMVDZJniNmsjxvl1tnQ4bbniyIeAA8oPPOh/W4A3N6+B
I8chf+MONVI+sxrRc0RKs+ljq/HuzojG0zDxU53bqLaruJ37+kGiVNW4N0988+fM1DoDfZMtjJyz
Gn0EmFrX8OBj/nXgEwjbXuXUhMLY4eUgWSYmvOFxcXAT/UxuuDZ9xyfY4zMaGj34zdUA2DDJSNWB
FOS1FQHfrz6hVaRrXZFMgnePpfpEXswJDfxo4hmlGBPU3huN/4gA8J3+hQb2R873KZxKyRLrMHOj
LoCaQTw3b9FxJjq+B4DukTjiyFfcLk8tDttpaDoTgtKqFWrCgDpN8Viben6wFT6jR+CNQqcvE37Q
dvd7bxZEVnT4pFGzyCihpoIrHjK3S4kqck+DZduYx9CYG9QhAHbLrkfeNIUZtNCLvpTlrMTdx82f
rh+7YAL5CZGXzTwFV6FdZeDVr2IQ4ggCrr6++NppYKcCwEkxJBgEOrUuNRzzy0o7aWDi9sJkFIiy
HKqAD7/TZmiR5lHG8pj0udyKbTY0eOjgzNTE7nwCy27RjUoyOacWJW2JNdWxgakZa6kjQiWTvZ6j
GhlTvPl94MdnyImCWB1JY2RXYT30ygpVfIJSQqsCQ+VCjPFnTZgKjZBt5mScbyDZSWmoSfOgXMoN
AhJWjtKF1O6eHnP7pBNSLJinh/B9V5uup1v5y1ynA7KuqNgHR/BX3ey/Qt8kVPd+15c81vQYRgvY
wgTaI0cf/+HkZeATdTLREFixsD06wiqlF1IgEKKPHlFmuxHErXhbOkiEFyv2E1PxzOFxYoRexYcC
k01DJh46UhBWd3Kxa5uA9a2wtIPnG3IrTr8CFoxRHhb6SNamDUcoY6+0EQWJ9XjnDhtT5R4pMkdw
E/eqdVjZSAAbemIu6A8D+Sqvolis8nvRSHlrJHzXE4rA/Pr2N2blHSlQuOnpfaFGtTC7VvwAjyJr
pTkmQ5Bub3mF7dPRdFxxLTC46lKicL5yYFxU56B5EN5WZgZFD0ptaBhItco0fECfSCBCiUZu+HFc
l/58yacgUUCwHjSMh4GBBtCduFYz22Y2OWjyRfNjM0lUXoWCPPhL0GdhUCNfShS/6SoQY33zjsny
LIZL67Yq/B8z1oxYVMuIYGoDpbXJyaY6+FbOauehABpm2hTEJQdz/AJuoc69uj1Tk5Ww/zNXfF67
v5LST+8MBd/HNfFEi+vqr1gb+F5XAUK2jCupNPz4pqgBfoOqmW9GcTuJ8CEKnyx9uZftKbPybCFR
uXMzxhYZj36dbCLp3aQ0TP30pOfcvcQ+fMRS7V27P1+e0CC5Yd04IXHaJL9+5E7tvtNHeRrp0DmP
fMkLtwqZITCw/VYKuhrP0HVu54MAZi/KVvgHWnHothi4nh33ugZHtJqUVVGG9DjqRB6YVYY3CBkV
ZIH3Qb8sB9qtq6UD4NhdB6PGuRkHM0TVj9CDnY3KJLjjnoXpB6WeXJ+/GhdVQVpBB6sN60DvexNW
tg4lhO8K/gSpie2XINns1YmiB5Gwv3BK0Zi/6DqQGFa9o4DQBiV40Pkj//tyEXesxqli1MJzwD88
hlsRP+YDXy9T94mVS+WkR8JR3EJxIn/bcSKXIbMmeVDL/IL6NQlK+cFNYWEADxkFTv5z0pXqkjaa
6MzJ3VlCKb/2KvGhtcNW184GxtFn+ARMWJxgzA85W1iUYuJ0HRHqGr07BjS9C455XPFfRvqSmoe3
lC7QSfP3Sl0XwHkRQ4bVokI9YwFy092ltbyV/2bFSzb8P09fojl10815X8uA4hpoeiEa9Wg4BN4g
H2qd77KF1BgyH8vc9um5EroHmPZDWEQdHsCj+viV28wAZEzt96Udxt5gWHdhpAMaFxRMKUojyueA
BUwjNBQLL4KpgqyUCrheUqEtb2wrPshQKs4zBxVwyuomaJp8RFyQx62Mdu1DcvIYME5XIhx5Jexo
fMLfnNoGbJDI+AXtolez86KTumTOFpH6vraQPXVsOr7gm63EpehuTWbW2Qu82UjSBOyx1RIksWe8
MxWSDIa6xwKqKXjhpcNRY6Ikj3dLGcJnmRa4LvFx2hzFYp3+lfJwu6pZFhD43UdJuBCw7WD5YvuN
WH4kvabx1b9ehYUTRLmnl7g5p7pGcapvYHdnxR483hycyNY1W7mO9z91MEzdNlUESIyBxs1rzk0l
tUx/pvRjCQpvyQy0GvIH1mm+zo0SWXO/mVYr3H+JE0csjTlOQoo0E1yy7aWEYoIV9dhvEHQyDuuT
+nFyJGbIzk+mEm/Q1UaU5Nc/sUP7dtxMsPooDYrtxLJ/CI7Z9bsvPeeSOWd9XvPOZ52wvUzSRq0U
2E5u/VmGtv4HIc3rq+JEH8XpfP6ZoSjpESUl2nQHIwM0KWagTIG1vwAFgQ3YUFX+9/K6yoLgSzUQ
85ZrG1iqR1vEqkMimf4nfNNfp4uytgg7zGfxUv6NEhM4hQ1uv0DJ5vAWblJ1bzOaHnzQ7S6z4GRa
DZcK7ROORoMttucE99gB9+ZAhs6zUiQx+0KghN+zf7u7+Z9GPY9kf9g8S6dZchUDdeYI+XFBUA2K
LCoWx5SlC7dFz98otMfZNk6xiWOuUQeFNE5nrFBZRnAkuIeeUZ5SYgM2rGdUMdycovd3mFfjcbhW
AmPZx49ofbIR2nGCa6K8HjsZkb4BqQcaj6nSFnbnaiN8hA6UAmT3HFCXKOnNovhJF4WR7kW2kgMM
fhhllE7KDX1JLu6ri9y8bZ9gZ8o42mVeBquTjTWBTYIx2wpFt1G3U7He+/cpDkW6C2mdssEEOe7n
hcfihEhb2j+heb7ySLocilbml5MUrKhugiYDY4h7CU8cRJLgw+cimfGcLSobc4lyEtRpNJ/V98DJ
W8uI9bvuvNam9IJMgtdRcGq1vUGau1vAAF+G8TQKxDksaae5xfXURl2gnBd/pEOGpT8ngVGb0bNg
cDm879LP5y0PEt/zy52Gm5NkH+9/acn+8DeYl8IToMc+IIVqGIRMqEdJSYSslj9+MSmZ5xifAoxr
0Zw0dhrXaGKfgmfsMDAGjLeAh7Fq1h8VcJIDlcryRaOknoPeSwHy05uFt8lGVqe2YNSyVPe6he2o
mbkoYyF3tjRACbWSoeo8lmEEhRme1vzCmOFtvqUX6grhHbz3p9xWE2wIZhLE0Ew+deyyGD/4vsM7
0O5IpKwIqeYG6t9aj2dCYbn08qUFKAz6+sWDDIOYRmIm9W3y4FNHYRtjL2zcd6++QQlmUaPOW76q
PfYVGA0XEJJVzY5qcuVU7AlpX9vIx2RdvXvSLS1VoGrfyAsvMNq2kK3chfvbM0AzQAfBBtskn1U8
ego3vwWxMTte+WW4vzy8UXHXeDsJH5GAHypD8bl9DUpaWabEopnBt7F+gzyVDDNyNz+s7eejOPus
2VT7AUZXkKnm08Q5ZnHyC2UEPT5t7n0hFT6nEYzijiot5aDL77r5lZAR0vZBOwrKdYeAlGlqeYxU
nHHw4hHJrby/xpDwJ2U5m3Z8yOaA1z5PtV3mznim5X4PsXlzANIhetfKEwKTqZjD5vd6YgDTLBPZ
Vv0rVEh2kr8vzCuHGK+wD21wm1kroetLnc5HL+5bp8PhSibNNBtZpKqlYm0cbmJ0NBlWcbs0e+DM
KcdS6TF2IMYX8s2pYVCF8Lujjzk11o4BEMpysJuMHrRs5H41ztnuabhsOw8EH4pnsdKrBzvmxtZ6
SoIRZ3YJPLEMSLg4uk7jXVk9v+CGRSh4f7+vEXzMFCGMRo6OBWwtGmXHdeD2AJqyAFSe8YxciZKE
z16Ur65ztZ+h62NpfupXqNF9YKXippmFRVbDfQZ78xVamdF4YkHo6dhlFC5NvWgviSNY8Dqb3T7o
sxdvIGLGHfVfgFYq9oXLTW5+9aU3ieJhnJvGO+J0ANbTDIMDuPeY42mOuxdQjqmBhvBcA97RhTrS
XHNyiTj0wBfCHAdKpmNF1gwyRKiEMdwgHr2c2jrU71PMJi1Kwl+Njml+XJ19aRuQZOl2wA/fhb6L
RVUVYPz4F6YJzQecsBaOWl4+RgERcvPDLwt8rSimQePn2r18yDSt1U6NIFrKHf0OKtdfQp7bpG7C
dNgXUPT5Tz36/yuTmAgOwo3YBNZn2HRs3Ejb2KSV1FLtJm+0SZXKe5TGnemz2RvUNYfOai1nstyu
91mDiL4Ejl2vX8m9ShgYKZI4gGD1EloTApJC8Q+Xo9YryIBzuynPBRgZSAyx53toSCGEBzTmFHH7
SKvD6cx8DvurKSsCl8/l1Uq33COzH9zUhgJIGzmYGM/VicCeEdbRMNpRKJ+iQYtpXwzZ2U5JwYLX
zki5+o49xLSal9uSJdkiPYDixkuEG80y+lDHZup7Ow9Hi46TtllchEEEVwNuHphROJNa6tJqAGIL
9BJ3t28bjdLxrdH2niNZcjyal/l1xZclL99PLDe8p7X2ww1MPHelzBPUs3RQD/o920TfGm/pvka9
hjEjx7r7KQjs1sKZgNQw42TE+dx/jgB4Gl7jwGzbGUU3k6nMq8Em4majNV0XrYeq8vdUWAtRj8nY
SzI4hrrVIoOuvL1TiMGsPqNvoglJGgyZCTiCfTaNAMcea6yEWYu60bZfmCqNBRf1niYBjXqo0w/X
Lr+b8H55SotJZTS6yH9HzxpioConaJs1NZR26Nl05WwxzDl8BbFCP02I3zjgEpObOjelcbS5nqPi
yi3p6JQESV46Lrn5L/WpjMq90rodunP/Q8lp2NhWmCjzPU6YCV0PTpLT/Jbf47nze2Z0eymLPqg1
dk4Jkbd+ITP0zSCwRNjpnT9CaOcli0k/SWQdTMLUz2BFyvk6sBR01CcazOUbZSiCpVxWr9Gj8p94
wNWPgUU9qYNI9n3nUuF2JYZbJZjrOBuuPXIojz75WcrQl5oo51N5HZ+364edldKP6GL4xPfPYNTu
+Imjam6XyC0FgJvaVNheb8cFgiahYTeAvvytbKyz5v3b8qy0HxrxWxNQqZu/h2acbeNWvB4EmwI/
TYrYb7cDNjZtyc3QPAno67DS68Dmiyqdh/UqvP43+RfgB/hYLf8B0bYdWAXpTX3tWXSDe5A7ybhA
YhPSzyQ/8elH+vTkiRWQKdaBIgSTVy+oqMi4Q1JdKf1J1OS3LAADyDW3GhHH/fPK8tcCkSjU/Or+
+dj42qG6iHE+EjK93jyjk/GlvDjSLHUQbSgjbeZ5QrySZfEp7/bZvyqv2zc+UfUXzDYM/nr6uWKi
SNyrKXqzH6SC1Mhu2FMydZEpUW/Nza9iiKkahZJHKA7s5TF8ge2mtVt1JOJwD4pGEySnOWj0dS2c
eiFVlHP2TQQU4jpxXNuJvnXXYnfxdOMsUUaq/wgzmE5SgxtG2E0iceyM9i8605W6Tsr4oAU9Gkto
/QU6tU97BFAYfyMnEjSg6DUEurosteTj0igACjrCp5OD6a2QT2QycJEjmO6BO08SVaOYU8eFaukO
HwOvMaacSlilpwFn9FD6ssYPkdoa9FCN5u+AFKvuvlRgWDX5A1Isk7wyxiqWc5qI+rLKhDxETCJj
f8DLZSNV3AcMVl3l9a2bfO+uYOabFgjW9aec6NhE5nNq2FdAKyv4ZAl4Ca4MYeCvHElRI7OB72Uz
v9TMJiqXPieeQPvWZJlSCLDXo3VlrRpnEEOik5XXx/ftFV+fr64w8YzpMOMsH3SOLdMFH81dUw+D
9SaveTuwNsRdf2PSaJdxx1fyZFPcf+rr2FEVmoS3Ys3oIUAGXlpQjbXM7e3baunSaa96WWJB6r/2
7m9WCbqXU+2lADJ6/yIyT3qgWwcFLziH6wnlHNDTIgK2F3MDwMsHijgR9yWVP9b4FzVcnow5/f/3
kqDQDK18DtFz3vCxvcHZIyZgtg2x51zBUtxvuAS11VJUHkChL7nIOrilXOGgi46lmfeVtI9qHbkk
SVbEkft3FMPh+OwOpRRkh6dgC91Jsp+sHn7ZePTPUVLd6qVPDCXjbpj6mRS7e5VzlnH3AJHp7nHD
qnrXhAdqJWNqZRsyLh1vrNXwdRNndoxovzcMJV0KRmAdxUVD30LTRqx48xs2+GWy/oz44kdgc3ev
rGF0u7Ik6SkYavCcg+If8B1QkIMX7eKMDqLwc3KBwAuxtzvyTDko90Fj9F5oZi75QLChl1A4i0cW
lA4fid7kLUOvWK5tXeurKWOVNkcE2trZ+zzzBofmT8KwDBelvkmkpO2gzdKQsR2zjijsYme2nMFH
S3XdpAWUz4HCgE4VxwXfvuh5VKfs2E9nB3IuGl/faoYwoOegZZzdiNt6m3sN/EE1Do3RKwWYQCQ8
8h0tWJxmX2iP7eTkhKd2aKQM7CPHosoD5GB8EB0fYU36xmnkdMnXO5w2hCQm/YJBCJaE8rw3jz3P
I/Dog/lMYqUDrOcG2KDZbGkldxjlYfyn9D4OOAO2MLQL1z042RikuB/52yZ+KloOy+JPtds7vB4l
5hGZqnwzE5j8xlW5F9SBvRTuxycR8X/k5rq5WA6c/VX06n64EeBsJ2P1j1e+idjm6lQQCmUg1Uyp
RNpn1ho0qrhleXB7/GbG1n95Xcu6F4KY4SRuIZo18MCHCDUKTL801yD2HZ0IEFFwzi/0nAu1GLTx
ij17V7HUfqoU7MCmaz8p8abYTmb1KqgE3xLJfeuREQZNPMiooSigrFuXlvDzTTK2ZuppVmd6qPpZ
6ZUye8184L00iV64kDMzjCMHpV3kRTjVpcK/IoFot2PNE1wLDv91qfppkRFSZ/Itmy0b/NU8GRFP
7ovUI2+BkhhlJ8E5iphfb5bOibR4FHFPYDHJUXGi2j9fpTsbL0I6HtZUWRyFHT4IGzToT+3wCwlU
4eU089iF6KyHb7Rgiz+Hd3W0B0SX7HBcEmCiz5eMmwbYs5vBRKniFyMMp/SKPLay/NZ5QLRXQFek
y1iEuVT3HWEuQIsvED6z7K16aotJ1TOlUGv+DV7SnLZoIvdUFFhQP8uJjVs3intI1PMUlRZuxyTv
YXtFF2iyy4Yp6xoYFt3zXZMkxPu4Gp3Re3YYc+fMRlJ+YRmWjRqsTrQEvroBoStrOCyZZI8GvhDF
sFNJ882zRDZ95cOt66k7mgpvlqWdIZDXzvJRgDzjlfuEVrrxHVDD80yQp4jyYRD/J6gUqeajU3x6
ZtBukIiNGYQfshfm9J7pZCun083PFcB+KorLmoei2sMBf/CNAlCdMAKQKSn7+hS+Mc7K20iRCNQi
7ZrWekWBjcG7gfjYKAZ6lE2/2/ooP2A2PVvbZLU+OmxzkWYjyY5wDnz8si5rolNyBUIFYVkjuPmX
cb2JFYTuwF6L9VIoR5YRAE6cW4tMzcm46IDjkTTQ0xTqvriNamwq7ZoZnF5cwFyP82yj5Ia4CMHS
lJNYc6TeWqlvpcw1vq3izfax1fkDbNFZtYYwLFyd0B+NQ8JgPJNW09VqbOFetxrVkg9zOhd+G8nC
0M4GUZf6HFtlY2G7XDxU5WSue+/267ZYUToL9vmdNKnltHS5QTqNQv7R2zrGub4zXgVBcIWaPm6Q
tBYu5C4lIcx/B4vJsB1/oCcSTm/BU7Tta3R/+uJ2xKqJ6ufTgZf9vAxFVfJaL8lXgK8I8IbsQRH9
/Us3DQCaAx3I1hXbB7ZpOJPoc5TEpHhzltft2VPSlxf5WUvc6m8btClCU1DrQTDdy3YI7PjjH/la
MWFP1Y3QDmCG5ei/gTE+SAzXJ+N6/MY6V9sWNQDa7fpGkDnvEV+FmwGIxl2uosFVGhswQoo0oDPT
YxO5PWSISKCjkHDlnOxYortwPpP82rpJeTQfFz/a9Vi+qlUnicDzU+fBylkAWtWC22R8q3D0a7ZY
A+GoYiYwacWJ4rPc0hwtRoR8VSsHyeiVru4TWfaXlhrcXS7diVHlVgSUgKLp8AaZAEVgbzvMigr0
f8xE4LkW0gbc4cvygPabGu+gQUgMdcqXhdsTDnZ7Wt/dX0CSApxrtf9sX9q/9Ek56qKnijgLklyQ
o0fPvkE+TQ+WhKcbbkB+XUexnLLsxhy06GsMsSKzyTeJzKLQeVUDk+cggfdSGx7v9qddKEW1FQBu
8vhgsziaTEwLhbve3tHQOtiu+L7UANhAXXJ2F3RriwA/u83BkerCg2B2veIEGG02IyvKqAMjcScs
EYqX2skOljwrhRJCVBFS8qjwRrof/3M+DusECvIz2ZsQUqRZseApOk6Nb+Dy5ovPtVn0LenIsglU
PYOpLMxYKtITJPfVj8tu0Jnc7Gs43U3/BXIkXIB5MNnfkjqUx6t63UT95QE+WF6pEgAYHL9gcAbf
SEC5mu/0NlerELy+PFan8ityPdmfLpmadxdRi6/sgEhnH2H0JyUN4IRSC7r+nFroEK0JT1XI97G0
J53HdyhT0dARAZ4fldaERiJn4daenjToX3fIx1/FGyNSqqhaGQ44OUSzAM9980lqkNMc1WwklMMm
AdKgdmAoZ15luABQyc8a+q9btVDMojdejJbGzxl7or3St3bLRiHKyKcVjoUuyINOSI7A0L9V1BRw
lB3NrD1OkhI3C3fN1IjfK1vV6gb37OG+dwmN9GCPtBvTNlOBTPjgchgQALjHG4mZVGlC2wzPnbyk
eomPS/VO+TSaxwz8dYgm8vo7ZmHdCbldiZzddl458YaiHEY2/6wNQSanAJKSYkS0cXNqrunTpd2V
TCH3cv4Dpzwb5YoGFMa7YZEYR15/walLQwH0SJwpuqt7a0BqcdpA7As7HtQlPOVlRwe819NYXaAd
XZmDjAzVa9ZJ7B7MwCe/EyvxFrRD/ef8+794/ZUSTUvm7Fff56jzrYYR1aGgj99nfpb4MCHPZ+lz
/3ZkxUTlB8BtAPv8syUmx0hWSMyttZok53Fv2qrEHdCWOGK77ciqUzJ3HvAsSZpCOvy7S11ntCvh
xa8EAzJYTUo2/Wp75LqHg5+kkVjgmTMaO/VyYfrmnXLTqw4XyuAUPMoC7fJUq+V99RsU4PabYQX8
3IZ9F6LddJrY5YHsxAK7R0glL3hKu2rda2XQIUHYuVJN+36JP15n/ZXfG45YAFIHvudNuIzYPYUH
qG/n87nLiqzgpc8XmkovkEU3RDxKArY1s+/2ifjq4irdYI9jBhEerpYTBRtxCM1th3AwaFHqYVkH
3LC/bo4Yi21nL6PGu9k4AZxxL72r5rtTZAmE9LUxvavmTZ9i1yF6bUzPO6IdcWQ9ExFDkjnpnHXN
S8pBeJ3QwCeFYweN8fd+esXp8J+yNzLGg0BvSPKAF5OVRZWpf6VYFJFpSfCHVzQUoFgATNKJVWTm
tc15Z9u/Q/YssyOJMvDvHNuAE2XwLhsLgnLTRS6dnSCbpHqIZHfW+2m9dH7rJG/2MykWGqtMLXxa
QI7op5C8o3IeYlc8vEwwxELaxKgv7rx0ywW9NfvpvazI7i01CPyHRAFRVfWMtV+7WN9MziTHSrCY
/Mra1WCa/V16J5USrw3TXh8P3JOddeHeWnlTr6NV+vMbSbsicizWiQWm626mlka1WuR3wW7iQv4T
iBqh5jwbm2rXtZx6bFigSPeFb+TXu6VR0Z+b8ySSdnGzpyAoKjq5CuKuxchjFyak8S7/r7e4+qcU
sAWty4uXUZomva8jEibQ5xBe3ZV6ONFDXFqOwF2198Ga9kjXvuz1Kspx8w0A8VNm1psQuZwTMQj6
GRrz3FKFd7PJxdiCqNfdRxZHWmnYHg9RimCdkEEIeh8mv9BQeARdJXOGh6lEZ0wmWDDhuTZ/cl9t
pRkzMCC/Wa7D4jbWLwos38rsXa68jSxkq2jNHsLHLF6B8NaahSyfayRT4V1FX5v9yXbsNPWmHIj5
haUJ5shiygLq7sEwn1zXpXSk3LwxYsUwrCZYsu36n2B7K8bgmBTP5c/DzzC8+4Fj9Oz+iLEXi2iO
dJjy6i5pB7KJcBTevJ9NASUHobCnnz6o77DgTd44Odt2D6HQHBhrijT0qIsaVWvI/vUO1HAqXFzh
DPZYjCEP/11xlaE2ZHL/sRSexGcvb9LcHx4GFadBa2K9/hUh0yvXHJUeXed89oIW6Yqlc0b9RFOh
PBlJoENXcFbRtNY7TkPx9INa6wOu+j/jLpSoBopqcO8LtKjovAdyJHpEYjdYqMb2ip+/uom1FREk
i6Vny/WneEN4llLFqgmyUaf7QPvwH3RbfuJMziASQqqAtzYvbkaOl01oTFonPkWMzLHJz//LF4p7
4lLbr5SFLnomMHz0PLTAoGdDwlkZqA4jZXSXraf/bucMG8XcVvnZi2k+shXhbO5ccfdJ0gQGr2wp
3kFLBBVk5xTZq39jH+TndEQnjtWlGzOLtPRULV8LYBZpGA9dtZhfw2DZjTp1jmOEu2xl/uZLAXrw
bAXv8VHrJIzSVLdspZIlEL7tSTD0j9y7gLDbFCPOPLxnjuG/8vnpJ6GCQE1MmKqagP/M5qfolNZt
O14bhLgYpzd+uaUUM8PnzNVk6DVRceDSlQTBX9WUYyrhZECtT0ndnC1gfJaY313ArjxeRDUQWhNO
bF1JajrjoGbh5mnTDo5zKq0/wf10rg0AQ4CwCqg5eG1ieBuuUADONOARIKSYut+dPN8+dZcTHaWN
P2TrhGsaZzePGyHlGUYKCIyZpR26YRR2CejG/Eh/dOup8+yCYldnK8VG2CsMH9eqVFxB2RbQ09sC
sWcSpvqAznkoeZY57jmQH2SnDDm/QfR/JSI39TPaWsV8f9ng40Glqe36xkQvv0FkOs5tfy3r3/oq
ELhS8cBNPMiNuXjOzYs1dCXBRrAZt7mI2t0+QltoUxCHqNzdV3agKXFqPxy9bUiizQLaOvjPmBVe
R2xcnps5pCdRrZMyt90g+kV4gkzYNM+etUKjlTWX14DxNZuCXwq4biPOb1BPLcrNUWoMjNTudu+y
1qN46KwRzYsT+v1Wdz6rhdc6giXq/31IFAH2cbyBPoeuMaoTmqjlWsp3Jmvv8P6gmXl5Jr/Kg6t1
z/qYsy1U8lQCudybzSu97yI5ALPG2bNGjITPs20GbvGFsodWIX/WEy9/Daaus2pyr03mPlPbH8wK
XN8k5fSsxDh4kfQWyldGMSHLPqr1s4QhQhJPje4KqAEsIv5jw2Cz5o7HMZetoE8CVqbLRToI/JKn
m5bH0YViNFxtkyoDGqcxosVD1UwAPxSwrlxkbXhJJ19Rr0JZvpRmV8ExC50mIzLkP7hF2XPENpm+
hWf0ktdWfnZl1YRjothH6KXMI9qmHFURcHwCIySScQMkPjQ0IzuxAjQgyt3iMLW7bhJKTIQk/DD/
gTc+HDEc4ZQAhwFUhZFpcGfBmCXEcX5yw+lEIf4AQmpqe5M+yntyN9BY1zjY9t6hqoUpA7kD1EaP
I7iMyn9moXPzk6aGMfCcwVnSbm0d6ff5P30wInIB+8U93Fnt6OMf4onxoxMG4US8vMk7zPjpyTNv
wurYeGx9nEhj8qblrGxXB5/zrJTySnLmzVygfQI1UQKLt6E8ssDOIc3BgpN+XTfFkWgHSuBJSWM/
qFv0tF2UwFc20mAVveoZS6TDzJ6aht19m+29qJyBuxJWsQYfsCgoXwPQEiFQC6XP851sMm9dSzgm
x7sBy6Qt2qBZH9i1IcFlvgAXMCeWKfgvqJl7cuzkD6gWAyZMi4O+ZXcYtWNnf8BIR5q92jGRVAY9
TOMRM+q7lzJhROZ/Q+qjSAI6+jabM/SAQ0w5QWDWjz/GlKXpsvtC5i5CPH1Di4yx5rwhbPPcSG5p
MRS8atVP2zW5hAPJ7CSNyqfmVfKMb6sUUoRzWOkBQBeRBryEmnADCtuR+tzZv15jMYB5hBHbjet5
DqBkq/sWLjjYXQEDPWr8UAxWbqF+NkSG79xSuhHofeoxu7FhFYMz3R+wb3PNLBwDX8zAaZdaEcFn
TByZAMSvtc8CXNS11pqrU5nI63l9ie2D57mkxl6Q857JCPc6tL9QHxc6P/uAAMWWCKGjZZVzBoTw
+bvzktVeG17tpRwK80jymCMpQdWDTH8SPqUlrxr5K2E/pdhCQrk8FU4UHZlyFdtg/Xsc97n9D8+K
FzF49g1HEkyl0M8zMR1hZJ17ylWSXyzWXylfXMmsshS6KUswDA1kqChUSgUZ+Es6i1rD8jTXSrlH
n5FyylY7i8SyfxywmQoKg4zROV4CbejwWK2l5Mnht3AEl23AHVLptmAsS7slVTYQ01wRz5EPiycJ
rT0dfdrKXV6qzgWtV4DxSleGBNPA/+JITgCEtdNh25QAtrVDJfC25fzzb4gmtK9LK9UkNU7jkpKY
sSS8AUESRoOK32ADozryqNw4v1dnlPvld5e28GGA6D08CWBpKFERehH+BzdT5NdrQuKm5JxgwDFh
saLxtLHZBNycwJnwbV255Z1R5Z6Tfhotsu/HrGvPXVxocUb1P6+TeKcN2D71AUGnGUucyKiiGXZB
6oifSy1zUrQRTXKHltal8hjqNr0eLp4bz5xL1tjS0LS57LAHgou+IzAo4nzBCgiG58XWXzRLAFXx
2EHsAzbnfwwX9/EcU0bFzbTdq4CSssHafAxk/FQNIDxhpVKYmbfgdHE6kEvvMju+2ipK2P8Ac9a+
aJOcMw+xlVEQppxZycBgB4a0NugSTM3JYS499FdZi1GBiZbD7vcTrjr2tKGay2UuvvK+d6sQoj5J
fvGYwbwP+wxNImpASVLhvkWphPnKx22OdC/T8DsQw00gpHyU+/+9gny4mtte2ic13X6IZKYxrXw8
EAYA9HJFLJs4ZcCL3mtQ6GG3ubzgPN30cb0Pv6kncE1TcuJ21sFbFENR8skNV7Y20ZXbu2ykVlMU
9UUKrmCeznck+MGrw/jA1w8NNnM6QK2iGOWUDY/+Apf/eLIvfR4PrSgcEe5Fe/SXXwdZuvQIJ1At
/yMxgipYAaglW4Hb6UySk8Tx9GHJ1hBFlqbWT8cX2zHQTV2wqvPm9E9M4Aef8yj3f4lgvVnHUYBb
eFk61mVswjMve3Yicmt88ZuEACeQRh0JAktABTH9/7q4wbL2USuyoP/lDiyp9F2DUXkb9NN8p4KT
x+X+1QE/EmCk1aj3IP+D99jGPqVojbF2KoP1rRwKs4A0qRf/zX5Loov4i85HtYZzWjo5yCJHOiAG
CVR3ze/oLaJ1cknvlBnpev1ZZsSE9UyBMV07hfls1AV2k5TNug0NhuNwYlLO1E9ypkG/EzsqsA24
S9emkgOfp90CA9WTRyfMIK0PF1YVz9b9d/TVxV1x8sSNz1MIM0iLwFXH6j7hEBcN+as4AXqpCPmH
f5cAQY+FVcyY5tVuFV0+26Ka6nCu2YXPy+qSMgAI2Gc/A8EI8HH22K+TrZvwI2E+1Xq3WSRuRdQn
4XIahRooSw+tcwVswXCyg6jtC1A6ytPthGby4BR0iKaSr+VzgbZnRK/Dy4cIeKvEBWgcz8v5XM4/
CgkyhR1Zr1oCKx7819aDdIbY4pr/pRh5OCjVFbunZSCxVNeKkZuoKV6YlV+5fX/trm9twauBuzNv
G5mtcHTquVJXwmcmLnuBP1IS48Wom93OihQKZbvWq/IAR8pY1GL80yUvEuFD1xstQTtsqX3MYO2h
sMzItzEUZGx/x5O5hfaenmQQWXlFCni2ArX2fglPbiknvWdxqmuDOEv+KPhJ/yeGPhR+OZf6Fiqn
o0xr5YdeFbvGe4kWx5Rsjx5B+xyN73Sng8Mgolp1rvjN8IdoaL950gBqOEOLS46k/h7NYwLh19kM
yLEYXIZr2rbA1j/O9XxBMw2kkGPlc6Mml/oelUXW5qK/Nxlfc2QW1JUvtGBsd7i0gUifJZO99Zdx
hlsZGiL3D2jwp6Hx2fvyEZrEErWbRwzTUlEZH9q7jbRRraRb7+XSKeY/JeZ0coZUZMe7BgmtCl7w
0SBcQyBEo5/8ye16wVcnjTEy9uMZFrRntWKo3lcMQcITjsVmZLnu2L3sA75h75hWPc6DZUEn75Aq
gIPw1EEpANADxzO4q/47rD/gHG/Vzp35q0qzEw/smMsnwnq3qLhu47I8giKx51I5veEdPABbKKcI
FJ0KS6sajMzILzqi6Z6GQzWcOnks5v6oIviKsovs8sIWT4+xD/9ojk2eNr3uepey+2SlQn7c+a+P
aasyG95rouaImjIzArJsOG2xCNz02RVB8pq2W/rgAtgOi+MSiWwV5Q96rytQpvdxaqeHgistCUML
1r2/pEYNQYCzuT4KTOieJ260DWEK2ROcK4EdgYuhJNcrckTo6tE7tAYaJEQKYKuxxxRJhTKGZvap
3elXM6Ze/VNDGUJ3SknVQVevWmisPvFRrQ/wMMpjR71lPeMfCADHHutj/WbiMkfVfkohk/3D4uAd
dqwXCIXwnJN9hstfvUWTydBqLmrC51G+zy5iE2KnRjUkuatc8TW6UCwcpfX1KeCoIlMbf6v77Kn/
MaxswbwWJLRmb1Qyl5PxY0ji3+dlPIE0blgkEpdT/zdHfA+JZlnWNSAWBg1CMxXu0OFUScaUbDWJ
seL1XYn6ImTGH7YyNSB4rejypDcoehARqHDfmHtrAAHSwnh1xtazfm1c2nx8PeVCqoKbFTdT3gbG
y4whUtezZwT7DA0I0yBm2Ye1DYZNCLy2W3a4Hw04PjmkfP2vN0+6OYkvDGHxuCsH8hlcJrHoG8z4
XSHDpPlO7Hj+P4z8g2+H+uM/6+Fue1DOFQ8Cs+n6L7m17ZHRWWUc0SFQ9/dpBe9C2X6HGRb8BIho
vyceiVQ7qwbz16mkwHnOC3PWdvMls2K74XpR/bESoNZreR6vO8C+GDdpS59301RRUi7+0hINa2+m
6g7WCudOz1GS0Z4H4n2Vtn8Wos1QdPBC23ElpOVddNMjikJn+8xUKB85y6yV3+65ddgUrU0wYQhI
fsLh4EJc2GkJ3nCefYy6Da+dP9AFaHkWIfe46Q9Qnob8wzXAcKK3hExOyVNKBUc13rWi6QznN6y4
mxAqqnhabdOKK/xCFQdRZ9WNKRTzYYAEkTh8C2+qJcRTKzA1us1rOtmEF5Kkzlsb15IdMqEUktTH
K92z4+zyX6S1UCusJRZs15gj65oC/e8urf1zpGaWcWRuZNjT1GR0QjvArRRmr7EqAvykLaCJ8xq+
YPF+dajH57RmIl40KfRTypJJbvUs1gc3AKM4la48Ye4Z2l9nJfMiWJUGK9OGzdH8c6MXu8LZSjRc
LsoFau9wj9HB7JwUfsnuk1yKLQfNm8wREmTyxL8NovUSIi9YoH6wmh/lWV3jnypWDlAf5IaJm6VZ
N7X+gqWblbOazKtHv9cJUL1gba5C4i42It3F1kVSTD7Xj70OPCtyKEWOlo1ilABvg0gYi6TuFcJl
oZHFCpXaao1NXOVZTagYy0bnLCIz+wxsgHVDlW84bUPF4l3yBkmgXNxZd41beU7q7DuRKjBeEaoR
YIXh40WgNS1rs9cj/75Pi1dr52PIPkDyzPXk1MS1xF6e8m9/cp3X/CskDw8HumnKKGPBhtKnfIrq
KKNIfPP/vSB4tlcBK9Z8aP21tHEOMSKkvaUWXvef2dqlM83xhTirj6jXs7T+bnDYQmkfdtoqDYi+
/+EybrVR8/U7NAf+s+c5CUuCyHQ1MJh8aCkoAKZ8x5fb/d8RYC7vr/sBKERcU2GyRseqGbPl7Aw/
3dZ61v48g4qfF3gLvL4ZY8yOLM3MvrDcqBL03/gqhRLDgPrYt0WXKBL99SK/v+eVnH3Gk5rov3Dz
2vL19MibpQ25AliKqo5R6pReZn+hi1uBpmKBRMcM9Uuc8q4uHdxg5+HTvqIYYURtUuAXoVGtdFZV
Ye0tZPXPyU1oKw+gNtyteYSAge+th4X8JwZ07TXEWju+l3AJeABl4CPscdPItEq+XUglRiqgCrrG
F4ruf7G8aiTE3iJb4bPRufQ14UEwrQlIv++lGyLg0DWE59YTXCz3sVAwzEj895kqawJl9HCJGP8q
5X64xXGm0/ACGMGHR7DzyeCKHn3kIQHb6v0FM+YmPc3lpJ5B1ULZMSgL67SQ/a0OxNrW18dN0U9r
4APOXOC9aE5k/Bi0JPU5xN4x00U+g5oyy/prY9hejxoUZ7E2NOLVH6I+PQtFo2KMAJQqM3WVL5rR
J4FQpL/rLynbKEp3fPq7/6scFhRsUHwbzBVDwjeWLgjHtZkIbZhF0Xa4YRNFCrW/8A7P+jd+OAXW
JDlbd+6rHx+k3DqvGD1HyIWtNqnmUcjHe8slsTIoZYQ4Kn4yryv3KlLn8ehUUE035XTuflNmFbWE
Yuodmu/gB0qH5uYsbmkpWNHFTgF3xdxForlkEkJNPZZyd/ojHlYNjO55d6VoQEWHgIN/83w12H5o
9uMpwZmRSfs0tvN5IIgF8/qNC06+UOhQdE4bP3VHzFAGOTGsiirHz9ZCGpjy61vwAiw8EvUdPTP5
NbK5Sk203XoTYLr1JSisCA9nzbg0C++Tjyk728y6OHPg5wMr9D83IDxbDdzrDwUwjGdw4uINr24x
IXhVi/lbABDXAthiY9inVq3xzF1FgT/+//eYNQery5kR3dgMSUxvMSVvm37IiIKAwzXLt0ieR8yh
d1whE1hMt2yPXcCAfn2mvdssfkBOWfwMr+Y74tZYaI033jtnBPLi0ZMdT2uLHvuxAyLB+9Ai4M7Q
tbf/5tChXeKM70gZF0c+YYNbedRIFwD82NK1gj1azLheqJUmDXHuV5sjlSNIfRURMcrDFRlTYh4F
rQ+SBLrQLwHLqsp6LMDnXId6MEb6TDdpBFd7oFj6AW6ZBnua/Ws/0KP1fZydtci0sjsN0Dkrm76m
iKz0wKdakVFH9qAzL7gXXDT9oJoeZ4sW96mQW/cHk6yA1sK3saQcMyyVazVhqFmosAW+p9WXxbPI
jC97EOnEYpHdpYbUKXJVOxfmac+yIXN9gHR8likXc/Ys2LYZ7PENm1S7dpC2+Mrs+zzYDgDNBOAo
p4XTEmlZph9kZRYkUh/fdQ4d2/Q3UjQuM4Uxyk8uApg/n4GCE+oatRLcBhAZuBmlZsEcQY4XE9sY
ThWq9xlohY3LiPFCUnK7HZzQtMAtz+A3JoVMDcI60ilOtj2I1F7EtE4deFVvh0EJUjQWGkjCnbNm
+tSBCsl7DjnPolOl2flJjrWkMa9ND+NZpny8aNen/rqpIw+Q6XExkz5UuEYapCXSWq6qEmkkPopE
y3dk1BBQ18VL5xv0sFWz6WeZnROgFWtuNqj8MdXk5joEyQD8yH5ept3oWvoXe2fbHVV3tmGv6C8v
h3j6jiB2HntoYWqNvucuFFBN3zJ8Jo+6FnY/PVdYTAEU2+VJ/wLPcnyKr6/d7wKVU99GmxcI/7Y7
gStA7DsmxEUK9wX1ttGT30oE3RPfLeadylFzbXH2LPnnW3bo8glJcc84SNg6YX6WApCHJsrS51+s
TPqW0tgs7lCcg0+cfkw2bfW/8p7bFFvF4yTbaqqgpcbq2pg2x//xq7ntHwheFkTqe5Z7jvKrnVKQ
SPHq79/U1UQuqBjUKPzCvjcHn4NmpkPY6G58XReozv1P6I9d1PKW5x0TP/ybJ1Ur3DScNPuKmQWr
vu5N08mkKHblaC00XhxGwEQOfjMbvWJScbk/qeyZ3Iw61Xe62yjafyTwsrzEpzL2BkPgsnt74IRu
0YVlKbpdagXvgmUtaN7Gx5W9CcFALoWQcwVPUo6Pap6pZ9Ps2Od0HEdwM6nX6Nx8U3tlcc8bLPpn
1WLiysY8/NryjjNYxuKH3LFQVdssfd04eKmdZjuueXWXF5meGcoUlx6j0jV7HYWNb/vDqc7VHjBm
Ew2xSxrKSpXW449vt2Z0f4+tsiqSNGO0aJW1D1P8IrDpgJHkT7KGHZBUem1qmSBCGS5q8v0fl0fM
hWA0XMWsYDIU3Gyo/BNhsWQMhuhNAnH1dKg/5N/hrMV5oHOxJQUQsZlXWucV91XCPp+HexxGnhz/
1x2gDjyEH59vShKjN+VBF0oo7yobhWqaihEM0uEh1JqyAP0mUsrLaRevVjN6en6LpIezjzSkzsuw
I1X1tucJy3+mvSJd2+YpeRWQdYD4bs3u/nR1YL/j+2DiC9qu9pU7yHqWwZ9XrXzH/9rc8imctbAq
oKm14CsMhLgpbtDR15MpaJFeXfeBxRGIPTkXQ2rb6dTUwOzu1fz4sPcDhrE5ENVUYJOBUHMbxSnn
vNesCoQOAIJd1LBzQFcI1JhJ+kICcVebymmSJ5LDXcKU2FXfEiV0/o+A5ldA50nNVYZTxqDk4qHD
HjHDvpOHDLdSqBVQOfoNCkJsoUecdJBbzoX3kUEIh543/LjabhVeHipvoETU9nvwc2X064q7Cfsu
r4A3VhSDnSd9uCHsxyYSnf9fLpH9bYjTvbfqMTsc2rPranJwcEEUyzcr4zkDbDGGXpFeacwC8mMc
MnQX9VnsmaJqQYfWw4lT4oGFdZeY3ImpoExyBNob9VPVCLIBGHZY2E/LgE4cRERe39tmIfTD2I5T
4MRMGz5YuoONRaFNrvb9LKSN3XRyHa8ta05lCal4v40sdQug5q9UeDujVuY/me+DsHjppWho/dIM
AKmzghaN/KRS+pNrq/fzpQIZxMaI9BORLd2099eQlBfLVeg6yekkIzmDp1fY5BJAV/Wjt5VNPk/w
1W3XTvcv4hZHl3k44eiPaU5XdzBz1qTvFHR81XqIxmd6un7+VHodOSECGwDK61nb1PlBTFLx4AmZ
+gG2wNp9OG2AgVLjSdnJaBJAc5V/TJ7ghmafbdiGfASkDDrzFeRpHkOrW8yN2isSfVJHIC0Zvt1z
9okOpOnhvh3deSmcSTgdhhVVSkZ80p8yWqWkww0X4nSGbZdJBdZCkW8ml2qLOWsDYAzSb5wuDnJP
kFNJgOKTrVpKo8EDzmfDAhVasMPQQACWBlD9iIxaPVJbeMVigg+LqyDdmQf82AHs/mfuVPPwmUdW
q3uFtfw7nd+sCcBO3PlEsvVbogJNl3S6DioA/K/GFKqvhi7ASw+UCdUwPaew20fCHJA5hcHfTfyJ
2RcR8WsalaYvtP2RZF9H5Pzr/wi2f5q+sxFBu8f4VdivfFnp5xsjVhLdxdeXbp6VnIhrvRcADqGJ
nksKvoS0WeR2QZBw5sAQPGPVgdpG8/qlUfShTr7AppHZqOpVA9eDgRUfv907n2DcbymruvDbtiCy
h7fsCdzKZILy/cwGLifZ7b5y+yexrKo5tKHkOlT3y8YrUJJOa2QPOM/NkZqWGtyCIHpTDXDHPswe
1FDtuplqguWwH14bN6nftw8J2QcqXA/S3OoonF6ytoWMZTe2fPg91hc1CErzYtIHXPXNS72YjKtz
zURRp6pTvCZvM3r8HIxPHXVKlK00tYiUNzepQhyoleXvytc2tBAPJwLbCcJa6c1NSTDH8M7sT1Xd
1d7Zj1wD9p2u1ECcxRNrNxF7FtVwZatuGyqzvzA50mzd8Vmbg4rMEfRpQCVvaxra6WrwIAQzKu4t
+N6/2NtDYXSFTLPDv2mSrhOrx40rXIRdVtd0uONmNbwJGkaNLjN/AnwJBM0aCpZbbw0DNHQBkfa5
XLa86aPfwfU3Zx6MPcylCbq70lGo8tOvYhti3mSFtaw1l3THH+Z/bhsTXwEq1nvZ8xnnCnM+ieDV
RrYyDyKfSR6m3uUHlRIWuCHkRrmzxV1qapli81195Hd0stPqFcnuacUw04xvzAwP/cV7OWhldwDv
j2WiAl21W+v6BDGX1lLOXd+Tkm1tK5x0qjgsH3C1sIwv7ebaFaeVegUIo1AEIrIACx4braUnoCRB
Rsb2b5Z72kNPGA7oETLEOLeWAbqGzBJng7QZv2bOSQMTTYD3Qe+0lrWeGFDyhin0ivD/SKaPdTcm
7rszql1xl6kkJBh+htFVdQA1KCnio8kFMzVEuS8j9hsTUJDGsCskwKmtwDGx32XOefY/iz4xsg3I
UOjU3k0vy3O58K6twJORYoTYgtgp3IonX1xWG8vIi4hbX8IKU8/b0tN9pYa2ReOWtJC+GT1RZ5Gz
OW1SKfXF7a3xxTZtgjh7yw311l+BOJiRLZTOTQl4IsI1mKgZMvnZPQ9tR0WcHVcgD5Z07xcasabO
S4SLjZP+nHkKX+mKNJt4OMM1I4bsRTXJoKtsrJeBSPtIqMOtMTPa1XNcr6qOrYbWqf0meudDCER6
TBq1bRyn2mSsJRFmWylyYRkRF1RjTq9UNa3kCi+fn8lrn1wvUdSZa9sxM+/5MBbvtR1/+ZZe4A/G
CQl2KFfHxyCIahUNa/PbpemIVWWCLoa74az9U6l4sSBGYm+JYVsbmfbCbV1K2Ud+OxGnlITIL6+Z
402PzMTHBMiFBzyftNgLCXCxosI+nsCMjXEAnOZ0ut9VOBaiA/wVYIp7QnBDUwWIjz/t2GJVf+hD
Uzwz+fpj5KzMTzH7HbzQu/Im8woLI9a3VhSJ/wr6GYf4plc9AaAqieMM09wxStYqabeY9X6XDdp/
UQYuc+6/LLYvCTk5xs7CRYoNsFsYs/PVPP+KJERHpHVfuT05fKHNyrhgbo/jI29s9VTLmIQKpKzj
lzx4Q+7pOblYHAPC8mqQpccoZfPB7ReMoZ67vrVG9bOs/kJWmCMtW1ZyqDyGcyAEVkTw1G+XyYtn
trhOucnWlLXX/1LlpLp8Kme7kSla9lLoDGsVVCP4QX45OjtltKIc987cr7HgnwTknzDgk72TJAjE
pdSFUUL2/ZBsUpicPGHmwUF8McSDfa4BNx9wcRy1a92+6KP3VbwLEN3bQgx4itXEcVOOdgDWTCUt
tuCgPLcyfyeNryeo6coQPF9gI4/SKiVjISQs2Na81koH0UcR1ULJVDmESSHDBSC/XyWwt0xmORiS
grFVDTOxLbP7M29cGoZwW54lSK3aR+9N/suTGc2/QPAdA9ZhBnbEEBIfbZ91D2UgTIbkBwfzs427
2Kzr4yiW0quhHylOiajToDiMDd4ZDTULQmTFKcQfPkMxn2v+E1IFesxPa/FU8Entb1tFSTcPFBST
q+udCNrozVwMjc7+dscUO6wWi/FE8x5PaamGKiOqqjG+pTOawOGWVDlSFIG8s3mR3rnNm6gvYOJ7
91iKCsFi9diIWRTIm4orjCuoQXqBYtKtImnbW5rhmy/c9lWKpb121d0oefIM6qHBOaMfd7iPn9UH
FQRKa2VTajm9KRejoVPsIZCzABsFn4qoikmZnQpji7poRxg9pQ7z6AzcOhZHQWiQHnPRXblOkBs5
2wZw5bfeffVO0QHBEQ74kQ3PLoIBpKk461YOwvJ81wPBS47G1wLmOSYyMhflxJdLpUQA1RpQsAiU
atDyFLhzPatvLCNn5WbwHA8D4JTva+Rif5lJVqsVBtgAo0PwS49ie7E0ufzGpomezxmFDSryof5K
0En3bcrWUKn2VFJ1YHr6Nro3b/LCFFoQuNXshtksonkkKCa5Bgg0bxGt1R627tchgnK8EzhYbXAS
HAYTRMvwgLPGvVpWzEjR9691mieT0WnUnj6Tm0ycJ5eWypLhtXkods0+lnxZu5dd5pm1zDF3kaWu
PxGffXkUljmhL+o6pAzCZ081uoScmhGMUlwIsukdSUIbzh+xqFrTBGrwzaZVWHsu+ioB8xGdbXao
HxYMTBQOwHXyUgYEWJXoy9t5trrbwBTUpj5Bs8XhScGHiAHlevd7PP/77cctBYeiGHZL+IH7ZC1a
Vzofj/a/z/LxM6Ie+SjiLj7w9wzOaBpa6k5EafUWhzAU9wdDLRSa02N04dxDn4VErKHtxAnveZSo
lHQvIcPibgPzEsc+QiFS4svFhtyI4rsYwC86WNM853H8+aS11WLNCPd8SIwNiqDjTcXD+nP8G5C3
sFZr1tX3LeqZqz56MYbcqe9R9+vD1isspn4GdHMnMVbmCo8Y7eX8+Mvhrl8jYot+/SmlvZ3NgzN/
dKdYL7vr8Vhw2Ku9XR6+lJQA1LQgB/vhfj3fj1y/7akEVTnAT3WQQBO9T1kFauWLTjQQLvLK0S5h
Of9itGuRjeJaSMO13RmPXsqaipOHHeizu7lgyTsBSC28fDqDZNHFtoea/BO3a/KctrCt98EkWe1K
kl3xbNk0A03A7FpgJnXSuoVICsxfZxH+orCEfTNAgK1GxC/ckkRGvcgrN8Wz6QCGLTFeHiz5Fitj
vnOgNkJcyw6lOEeMdHgmwvPcNCW6JpYAdehi9ys+t3zr74MXaWGlCr9yyyzKJDhSldBD0ua+9p13
85B+LDC3bo8udsrHZlYmbba23aeq8Xpp0XFfAQo5JpTjDii7uNc065yNLlwPiBi/aufP3l4F1HZ4
Q9xVP7VJPBRKgdC0MX6WuCcFI8F+burE0APAN5vg+HcKjm76ksQEMzl2ZxlVl/EIVVCVH+esrkQE
opzX5MoHqLgeYiJP66cT1d4PUfzpZnheytfPTbCQkxpe+usPrFWCEAIm5QdYpUKIPDbkr4db+MhS
qNhKBXSW2P96Do/qO/bV2SQlHOKOzTPqTBMARUYsOvF7QESoJTDKaj7dEKdT498Z8xiNeE7F7n15
raJf1nLWp8cf2o8Sq0RYpsi3+ccWzdsHMlfLrtkmTu3Yz/wb0bIEPK6Sym1CKjLux5CjHUVlmso1
Ahre4tB5sQgysDQUMs2sYSeF8xf5IT4gFk+qMibVebq3LlTPOB7R/5H43Mq9GEpumJaMDQgdzBoF
6glXsGsCg1wwosSwlCi7LBBOkkvhqYA2tYFBISWwvotFK74aQOU3qwxXQXmd5fn2o+XDYJdfgVQM
gHXtIESTqmGJZAyLJpcZU5f5vltKGRGMDz850v4A6A231l6JGI8b4tTQwFr5B9LQVE29p1sic4Uw
lcTWBy9Qr2tyiiz8f1YJyJ6gUPKmLUIf8BZZ90X6l7j3YhItThI1vP1vbjZa1/TgblFtI3FqVDqq
7yUQqkJ7Uy4TqYg2ZtmPs7bEThNgvjL+d9SCTzDdm/IHU0dO99DDefYQuGzTz1wBw0iYzzbqaZWA
3b3j/RvOxsBQEFsE1XaNgtu4xNP/53VU4mcTp6QVEuCV0vDCqEkjdlGmLmKdtjFcrzlcvuKdCPa6
zt5xJJdtrCkcpZYCtHc01Y+d2SXKXCX5uIi3GR5AkgHT0J4FKAZW2MwF+ZJTGVDEhSUVqYx98jV+
oy6234SgD4Yc/Q/Q6hd/UpcatPwcRn77ch0mkd9nwkwMJE+0hk0eV3eEPaM070/CQ87GwKhNfEk+
KdyytF0yLPBLAl7OAtC4Z/P0Pi32AVt30ZssmxIhRaxk7rOUN0b3SQnfJEAiPejsY0AFGUTVWKui
UxWDMPo9Xu9+nlUg75Hi48gan/A7xS99Gpln0n3610pJLiK1RcAgProzPf/NJCi61qQWKguyZFyG
QPR/ixm7AxlOyeq1mGxX8SQd/INZcR+ZEuQ79UvpFhEFGV1y6qSi4B6P0aLtGfr77t5qR9m23vRq
JI4AkcR12YttJ0YeaipKgtkAkshfLP6D451F6pTZEA100gmcbnMxILt/mbnlTSC5Pq/QBK9vn8Qh
DNpuZ6kEXGwQiYyyg8sJqWfBo0QEluW280LAjVScS0oRA5ZJUIV4W2wkxtUjJA64CkYgBNphKG89
rhRIjx4g5ewCcwxb4Pr9JCC66wxzX8YwHyvzC6muxTSKJCOQTrPP6/nIIwPw4MKy1iwn+r/qHR98
3St09BHPBxjKbMOC62c/XtEWoY9FDCsUHRlkK0mIFw4PhMqx3MXgekBOboD3Lh5OVToJj/MA1YVx
r6lsr0sIkjHQw09QXKFzbl7kBp11k+l4XWCLtkgKgHC51VhZ4NksuyDBpzFUKFI/b5coTajEcIUf
WqbDvYAo96tOakTen51VnBerPgC1WlGAqAI37T4kifxjpd9vLrT4a5U5jSdLZjJDkBnMZJwFKOKv
SCSlzMONFNxOglbOAts8OYmU5dNS5+zAenMDg3x7C5A/kU79cJljYpnjf1B4ah/51q/wPAy2VzHL
TvjutoUceK7FgHAJ2owYe00AlvHM2F6pjMMdBNlCQLUfY5GyeLOy1LDlAgsGOUmpr/jmkaVotFgc
AddftbIEM2jZRzMzt/qxVBaHRfVw4la+ClkvgIISXpE1103gq5WMcxqScShnnUIaSibq9g0Gb993
AORHRxKnGS29F51VlwolPWeNLVmeyqaAuxQZ8Z1T1dekXDKNx20XsLaiHBGanHBYfHcR3j0TSrV/
b5c4MDNs9rV2hJfaZUrrX1NbQEu91+NNvdV809QiFF7YhaHMim5/4JXP416olC3BvFLlCY3TnaML
px8TJFnSYAg7mD57wEs9iqa09cd1VwWAOGYeGa7nHqLfHeqlCGBXHalH0zr5CYfYtBR4+uDxOs1w
06bC1urHumEykbXZuE/MoglFp09zsigVSff2g+u7PC7BW+nR8UGsQyzLwzexc1ubibmeOBBxMeFT
4ICgWpVlrqZ2ROZ9IEZ8UfXNtX7etz2e0ql7OR9MnUhJ3rZxTNOuHKbq9n/7Vk920SYQ63fr2bUt
MxZ5crUk54PVIu5Q4Jz9UAwxZ+moqiAS6Jn5sNrmohb9xyfKZEWgNLG1k7Ixur6S1XugwOZNl3BM
5LWn5S5XH63PaoilKyICStHoEDVaNPZYKjm0ltHbCFHjlIW3iGq9SGpS7zTkghkGs76eibiJ/GXK
tKPZhvV3sn1d1HwqQVH5Fh9d5CYJqYGvGbUuMT861Bs0ALJgbwqKoMWjFzFwqZZcEj4UlwKPnNDz
57z4lVYXjA/bne9OTsIIuv9eco+K3f/pIXvU2I7+HdPGXS19D3cs6RTCtMmhoxpy8wml87Nm5FBR
a5UWtinjDzARsrZewz4xDe0TRsQdM0hBywZXrGLTOEjx2ZPiByqieTB6JiXnOdvmvInQx/B90d3Z
5F4TgeBn8UZZy+6ltYcwNVUFlZogiVYCzrtz+MKQYBCssoFRoHnrhXsavazvo4Ds4uvmTHPa1jXG
uaVHhh5M6Yuq+kzUh0pxUqTHS7LOg8lpJMh6p8TvvxaoyJi6nh0Ip2epcJlbA6zOurdhq2X6hlga
pjhNO+B/Ul1Hb2sBnGurdRuowRlxwiXcC3CYRD0PdyNevvPRLDz9/QtfrCCcg4kOh+tED54P68i0
eFKnfeoCFXlt2VDGTYv2GWY7K4KZvfAhcvRdo8SnUgpsH2plzl02oRm0XWTOeL82OzFr6nbO+HqN
7a8NR51fIkHBlyvajoWkjOOWDtGHZgKu76VWIZX2sAZihpUevWANpsielNS/3j+0jZ8gUnrdttwR
62JA8+Fuq/ZIVO5JGrqZOw/+5SgXBJ6lTXLWIPk5Okz+KT5U80hSCnzLl5TpZDwnGFOgzvAEtI6z
5HSRR3IdDvgeohYqqBpncdodsVLVekhXDS8KLez2xiYQG6pLpfbf6+lWd0NlWKyOyCB4v38Alc34
nH0O4iFfPDsBXLiE92tqz9dyKaPSMyDLXvHYcU27o4cl7PxcXB5mBFV2VI1yRERb50EThjXMy02E
gHGoecdWnT1BgaVjGQeb+VFKa/KNNg4lbUtuk+tpsGPlLIsDPhnYVBK7fooc3JrJTxKnKjKvksts
VvPKG8guFVCqXQL00iP87uDDo+sVo7jzYPAlheRPCeWrFAdiZd3O60dw/DkQrG+M5szeRdNJzYap
HBjyzhgxuytwN3ZQW3rc1L98LMefO+3Fzgt1g4OMh31ZXL+hqDXUAVOTx5RZ9pwfWesStHbYCqxZ
Tds2UrEMGuGQ0Obi479/VMiO6q4iLwwxfZ2anY9fc3DIIvoHSpNiQIDgXHZYIa/qUU/d6MTq/22b
KsP3jkIP5+wXVcyQR/TJkX0rbWFXIIZovLpCjdnZsZ4dpzqNhv50VrXMoOeM/aM+hcm4yI4LP0bc
i/FqLV8RGIrG/mVCVp/wH55/kIAkKsUCk0hL1hsnIW8wqW0hwlJa8V6ASmWm40PBiqwF22w+g8k8
teYbyljSUlgr0kG6TXfn5keTlg0o+cCfhdEQeC4S5jziGvBCXsfBIWFLePB04zSkXSUdTDDRNXr4
0kk5N7d8K80WXp+eeN7GiF4gbjOAc1QECix0XpvRP93m5qfypxsqcTK/hv0hKgdZNDSbr3oyCwyX
wkEIkhyF65c91w6kFP+PlAdKYmpoZ/+j3KW22sm9jsHDS86qKuIUNLFOYywxPUInVdm44bxrCRkW
GSqWbAbjlMMTsknxtJPfcK81yB288KmESGfxO0+6COKQ0ZFfSBynTb1Z4I/HPu8TeI9z0TJryrT7
KvYjms55kAL1b9l+Pt1VvqJDGyjuUE7p6IS2g5hvxxZEBUEX1eoh6kE/6qvLClcpm36UYW4YrJs0
aHDs61Ib1Wyc8L5MBoQW6vu0YZPp1RpmjcfCMIprVes6OQURD1Th1k1qQuLV0MCPGtH11e4hwQ7T
Lpi/CKIfUJJwQGjgkvxBudNAAEMB2VxUvnqRQZro4+cr3AJOz8HMy6YtL30prx+FtSTgEaDeVikN
7U+3K3r6iCvFh2VdAtB9kCdfy3SevlS1y6CzBmj2NLpVUF/D4H7zT9I6NAS1/tDW61jiLN3YrXDK
05M0NRHVdH26jQPfytQzyewtHba5OE18rIGkYDnJMGoIV2Ve0XpSg+t/W708oj8RejATQCfrj722
pBs+p93fcW7vgCMf7VfNvAZXg4XJImre7lSFzxqxuTCnodBnlKMMLldwR6rTCj08G8qRRHGhxWD8
a9GIFu2sym+Q0vHNO3W4RDz7aiCgvxK5eSswezWU5JDHLGJavLUxtSKXkDOA7CRlGoBB2LFEyYv9
G1cAIudVV00T4xAmL5UJR65dac0YjAFMvQOA7l4r3t37M2y8daAA7MhlAmF7QIcFS3pkwcqzaFMy
8LRqMVVLE8NpiQU+KPI6jBr3jWDlEXNTbR8ZnbksT6AqhyTGS3kJAZ8pXsvo+IuxmLN4GBQLOJ+S
4M7sZAb1UTyCo/j1tPr9mn6hckNbg38YnYUbVEU/E4ZIqDCa0nm0nBTgdsCabhCwcXRpoMNzmu2H
5unlwugVv+sAGV4RaqLrXX8suFu00buQnR9fTJOUywbjxxynkLWydubVRS5ZOQJ3YrFb87tFylQt
t8Hh74fyWYCRlq3fwx4BpjkTV/ADpIk6mBXIvFH8YBPkm3SsNwU+GGJOJmsGtCJ5yQYyFhCfU+eb
FB0POWfTUHkpTw+tjCDdrHENPRZhRRXVIrCDNWjQOGCrnRCP2WqdTF3CymaDpdz8vpgDvk8vWVrK
OvFTTddUwWAJzzAlBCeXzPcA0gngwtIk7ni5zHnhEfyS7Men9zYXrdg7RmCeHooB6jLp/nILEEr6
54Cg75D1G8/u7Pzd+3GsTRbwwm2zre/GXFe0XB4jddumWC9wqVIlzkaWQa7p1LQ4OXPS3DPu35fL
PMK1JeK48rzdVs+D3IEftgGtvB97BrjBwSLjymlqKvjQywdejq8rEdquhNH3LAqcm3Z6bQfR8qIr
u7kJjwn7VfYohkWWuiVcxcUWukGuzAgHdtpd09WaJC4q4s6U8a2lAX9Tw4BObChb3v/Sp6QLo2if
r8vcVAGaTj6YGlc48nyEaG7nMJ6k2WAbqsXNPlaUjVGoSTSHtGGyK8P/UM/qRqcTsbUXmRH7m2Xm
ihiKozHAefJdtgPueh3swd3/NI35RC5ZibOUu4r6ncZMGQApmxyDwDTYPa2LRbND3Fkc3l/vi8At
9uKUnVAO7Ah3r+i0iT8WrYuKQ4W3CP8f1JMdcZ/dBoFtGurFpiX31tAWpCLlqxeff6yXXVNi66/N
Qhymw/q9CvOfuz6+mnuHzRJIvTZDLplOyMEOTR1QPEQifsl+hagbYBJUObmNBfe4DGyjM+5RB032
OgkUx/r1V1qH+cUQGPcvqdVfLdKpzLxgJkhEOGVB/zcmG7Hf+ggB8mBg8JbEoJ/zzlzAPe2IBEyD
GWkEsdU7RrHglX9Ul8lFkaeNkORWTzuEKHkcb7VH9doCqA5lU8IfnjmbUB2m4HdD8n3VSMwH9td2
DnVFM4GDry6pzzx46wz921ha+dc8nJIMlb3Qt/Xx939c5Fl7jolYVMikJNUEcv8+k9yXVu+75LD7
mZbDCcqKfvTNinZSqC+jugTaTzhxN9N9jYBuo2zvbtufOLfuLeiEIUEU6U0teXj4lXRRj4NIpS2k
3WOGDR6Plo/k5AAnY5jGe7ckTHGMBAiXdKpZIKrh96vG1qs4DlHPxilPPW+2c9PkEkGZ8V5luk9Z
b032etPWFcVGUXtCmi2Zqb/4Nf5IPKLAKuiqWCwAq54pzK7nZN0Q2ntGrKGs7k90tb6FfdMePfwW
/aIb4pNgbjMphsOsTQAvlRgf2tVOgjCr2QwoJBTPrI8ZmWdGxvA1eNfCWnzm+jFcp5OaxE13uP2W
8zZcADsSrpL8TiEXrd970XFxJH6a1kPoJ0leNBPAEGYwBHUF56KY79wD6RZc4WftFIZ5jdcz5ovf
7Kes3/r+EKE94LEs6kZqj7BwywH1P6I2dZm48QP2L38nviBhSu9QSaL5iQZ6Xp3Sft3X5wdJDZiy
ENosQHN72+HHWD8TOGTWR/+f4LKwvvov83mPQFW7mYRlgtlqTtPqKDQ3XdxqIFAICP/6R/YUjSz9
5R9RaKNjyI2xRbFfJ4yfiBttfe7T+Y4F7Jn/Jxl+RbW89OyCa3riWh2m7Dy9YvJ4gINM6XSRn8TK
bpNRR3iUd8JfsdYWs7k5cR/U+B1AP96X4I9ZkNSCFzd+zphgtqTi7p0fCypYMdbHyfmk42aPsbSZ
63ZAElIMp3nvQSO0lcjIcGiEt1vrIg/uLq0c8SgPgR9NLTi4QOOjxonPzTRoUslDyGeYRGBNRFd1
H/8Cb2Ohhqp6RQprEZ93hgja+ogTvO0Ae3DTFUsNYsZ8puBHhP3ILY4sskb9U7ZyKY1KGMEWfuwl
zJ3D+tpVRXPyvlXVY1/ZivDbDekU59omufDj6xKLfudBqU4hn/VwwrD+ouRp3mCGSBuLvSw0swG8
u9h2FBBdm0HWO8gYO/oahWanUSzI/zAoLm15HSExMODL7t/CYV1IwoJ6mGoTk1m9AbUnAWL0hYbm
f3tkVin0ytBK9TNtopPwzXBGtvYB3e50WuL6mOfoCta22lqeMr34/X5eFdBFghD6NHyrICSOX+ig
kQ7TioOvMJvGlrbTDf8ijZ4XG+IzdgV0FfF98TZ+ybOvZBQOD6uLXIR0ExR0CQijUNga1Sbxx8WZ
3fpIWWKttHblGXCQjNKAY+CpH+YZfX9pSdQOIS3YlXoMIwCDMWr6RsfGcRdfcZbUk8j6HHzhdE+F
aM2x5dLm3zYovpfMzU5mGC2ovtgE1amork0biEwCAEX3X8pXPwPrWYN+x4EWAI4MF7iNi644AGSq
9ByvRv5/LAmFU1phywpAxcMTYW/uYDnhAna2LWZw31F3av3YZHQFGL03h8XPWbIzCwrzfjH2StT9
degwuPgJobKZli9QcNMgu+HL+8MkZ7n/rY7H1eUXR0AOD9kfFT8Q9kiAlwYlQJRrKM+T0ApdzuVM
rZ1k/G9/HLcxMm4GOPR7T+AZibcEdax0HXkOqqMxGLxgBbOmtcHsGvf7dJrv7fS0wboo9GsVlo0e
znyRyIJFe5N+7ZSALpigpwWik+3mUd0qv2kLAn4dS+xq1sM1aigbWeU7bMcEDoN3KJmeQ3EG4FFP
PNqwiejm8cSns6tINMUZ17eexE+W9FnMny072zYlYqyhpWQjeewynBpEY4jfHdTy9uK7uBPg7HUQ
9fTa0sJa6X+8a92RNyAbpFmSDCPcCkltmvPYr/TUQSFaM+0M9h9YBR25AxlGWuYiTFOQksYiHMa3
dlpuGRMfzdtV0WVVABOwwYyyajPIIm2A6AHxTG5lATdb+zwWSjEiVqXDm8qbQjtxqLcGPwuDJzyM
ER4povRV7cQyArBjSi8zUg7VS+etNWP7994YSzdB3BUMpYpy/vNUuHfHWnNELNHEqgx1fp80U/jC
xN6WD9IbUq7MxbeF2oVXEirWhtpgIbb8trfvFjr0FBKcVQ2pPHJ76OwyLhqlmKfiZ/R2NwLpbRuO
VsS8O8zVoIErL1y8JudEcoPD2uAU6VsPb0phiKuK2EBQ8tuMaLNh3V4/mldDvFMHxY4qulGi5Dsl
l5Fj4DF62W2EtSLVoB5yPcpOgsfqw+0Gwx/X/nKAn1pz32fjsRzKctjA57JuGr81M69cPMIFDDiL
F8sBQ0zFlijHx5PkhuEv8XvsBksWxeG8TB/4lFPkSsV/+k0wRGwQT0b9riSMfyc3fnKZd7T2QqY5
YM7Zz3ffowEttY1TDebJPk/vDBN8jgSzy/y+5zOTQxHXGrB/S/yhnumnCSqrP8c2d3COXqgN3d1n
URAKnr07pFRD5Ux4gtuC7ccwEad6ZHLYlZPIvQCMmH3MV4Wg+E43WhKVoOUj76tXFOaLFShcXCWm
bJrfJgforjOFmC1nMTLN9JPJrVa/JKy1DZeUKC9dih/rd8SC0kNK0CqXRUeAfdskxiQfVX2vAWqy
RGVI55PqtwfTjSwkTDTIV3r2MgaPGzEWo5tIN+o0bjSlq1QEp3TBiQkGtHZISxUfQkbPfkKWyTHf
nr+mJKxntuoD+74xFw8jfX9fEEKsyKyXf9CysBcPoBp/4ETY6zxkmB4I6I0Zp/mPyan5E5m53jX9
/HRsSJSN3CEDmH20aiAuE8wPW93ylxhlMDaVWE/JfI30aKHf0IVtlFbruQqXLOYGSHGk9dy7LjW8
+ebfrzXLnEgCt6lVfRlI8PcRSpUwTtdamOG8gHP4ujpX7cmyCnWRe6Wi94FpimT3V1ciZiWtAg1b
nKCiOyIa5SFtsGCeqHjpIm20eyYmFJu+2NDyDcu5zvD3oxXK3X+E25RrHWv9xFjAfo0MqxVul70y
i7uZIZfQaomo7Ned18ehMH1WkjyfcJ9YOu83ZDr7Bm3mdH7Yj0ZjmqgLcsKhrA22GJnmfK1g1vA0
XdahxZ7WqyUo90au7R1EIDlAo6XLKLH5iZu38ugNeN/LNgoqYT8l7VbsDqXOQXrNa1gJPrxwh10D
mmUUmpCZ6ny3hzvwa2c//XQ8qNfyJJZ0uD85AEJleFFgc4xs3R/PatwXraU7ez+zk0feQh9XElet
fxmefWDW5dh7o2nqeWZeakGWssPlKA3r6L+kKvUvhKQ6JdDoEcalU9aiqKs9gqJzoweFH1XG9jie
ID/09cJwM4t3NVpLxWG9QwziVotWn7hYvxRyAtIZUjCfU02U27tuSFmUvXt959BtHFzZyhnAHomJ
c6mr/xFHPvG2kXkAFulJDLk5dj2kkosboE6ul1UncLzSh65Ygb2CoOWVN4gctVk6pl8AQuyQms9w
GB8NB85/w9dwTSw5FkvL1Um1ouCpjyQ6PIMOL8bbT3flA1i5hH2d3HCHJhp0dqI8CjMQKIj28PHS
/xyFxwngVX08pKnCfeNnP+zm0m302Bh0bUhat/HkvAYuPQsrVi3mOQlGBzCe1bixy3efmjN7sQRp
6Vpy/9+U0+mcYeBscJs5C+/TBlQLp9KKsATMweQpsesArpDy28TiNOiqtg10n1wpkT4fFUQqkK5Y
7EufOplFNFvUlvxsmf2pf0/7id5KAYNHYIVqA6i2WswkVAIj+p+sVVDN+ihD4iF0v3STMj7udUOn
7biy1ikpDlUCuwPx0NNukyF+Rint3HJCDdHOET7jJKL16nMDv/sySLBB9oyNtZl/Q1XSKgm+OY/u
8r6p3u6Q8HCvi8r19lMp1b8eLeTZg9gibLGrELqVt7ZiLFEEwqTHnUvzO37dBBy09+uP7YfR+z3O
37MjFx0mdUNz1DFbJd417lg+NJRpl6Bpg9XRfvhK1TOWYfa7vDMtBW19FqYXoa9vBPCUPB8rsdCs
I/qrv+OLLQAQ7JyWhH1LL5sVUd7MhLgvCm1LBfz+X0qSRs1sDudSaU8nIHpZF96RnbPc8sfbUDrl
PvJi3y0Uihk8KxaAYLuZFuPeQMDxikG//JUn7p1RxSts6cMkdCNf5/rMRKTA4qS2m1J3X+U1cVb5
LMTjzuOjJv9mHZ07L+KXtFxELDot8b8TB5ihBRuPOvH6HC5BQ+XZzz8yH1EqY9/tckG7EpFGVU5k
RKGPCv5v2MOl8T9B2pVXF/Pa+9vMQsf7yU2UlJccJwn6IKyGaBMe3UYdIcCJ2z2wWZod+sOc4Lyn
EpB4Mw17/mGM7nUyJIf2nIV6l2bq9k9YNtilVCEq3jVG883zsxQXOB/Pgz/zpo9UFAgqnXXhANjN
mxdLJidBKi5vXE9s5WxFmwbje+kKh5gdhAfr04+KzIGZwjC8pCuZfwFvmYDHWRa37Jg+MCPrNeGu
0WR6RDHxKQTsps2fG6hpfWyS449re1DPJsddCxbi2xakOIZcRSUGzNc7XsCApIWs+QuFPcV0PDjy
g+7JaOytZDpZztI6YOz+UBa0BIqpOrcIWijUHrtD5ybdaSf56aHBVCLARpi6e1a+i5hA+y7NDt2K
b3l2XyKwVlYcXzK8Mq1TyP01j9FyAMI7pNHHzJdQ+hN4+dL+CHnzL5nHGzdhJOEqFGZw5lH9jkj7
J7lFZaFm6IG+9HfVa1YhsoOQ64P334oeCSA1r3Vy/ossAkpz2VT/xjFEBL2k0+tL2j6nobdP8h0V
3EuWr0Nre0e/BeKQ5bKpw1RKElkFb4aHOYf24fwx8EYbFVowV3I/bzI6vknNNz4Bc6Qbh23cA+oT
1J7BeZRdxp/H77NdajOjkCSBWRYr0IBhkk33eZl0Ch0XNFkHZSiy+gZvd16dZBTfCavN+yAodFv7
TUMZdZKcQbz41XcL6SSXGSOsuuMLn60303b3S0LzzcwRjPG6589bzJ5a3vKWvjSG8rsc+1zz8Fnl
ISTM8EDrU9nDTMjP0Xzc/VvlzfPw7xi/7zj8WA0Re7OVKmaPY2mvCtRTeo6+Q6eBqrWndPMqRAPT
OWOSFnPVc3QGJGirWo6LUEcPVMKpcm1/AONSemSPSALv6MecL2dwJlphylXfD8tFUKvkBsnxLxOy
NtwPidEv60iIx3vpMkZluMZ6Ar+akWFUkBUShwGO10FJ7ofXosaN0tlato7xkvs21RCxSZILOPm0
OGZm7AcLxdG52fF9k3nPnIKbq8WxrVvkdunB7Z24cMpMj83V/yB4zdFhMuclCueGWE0wJKF73SeN
8YmXaxHt/oAto4Fh0wUdnjIfyHuh4KqR+YmMh/JuyFWsKBT/STaeBIXpbT8I71HDKCVM1+lnhm4N
ib0ggByFPWKoeDcZKI28/+ikqc61j1BtFu/QtL+IvHYs7jyAmyO50bYOOv5UtiiU/Z6070v8Sz4l
zhZRp6LG8i9cIYc9zxauh8PtE1JvEuwIfKVIqHvIvrLRgmCK1WWmqEJIH4+ZbAWoZHVfCJQOqySm
3EL5FoFR93WLe6I9zpLNsXQ5bAlcNdSW1hQcVFtpY2XRUkzznmslvpNQ1M0JKv9PE+QLLDHLO0fN
S8SbmiNhDEmwMy+1tLhDADciZB143f5NLxfX00assdxZLeExeMtRqp4P+sIg5P5AyE7Lpd59Fzt7
8HhezRIYsmZESXrpsxDL+Ydx7hnyy+2uEG0YZUsooiPq/RV99EA/uKxObV/c8C6BQpykiU7TByod
g8ro+ZHIypCrHm5WWziTNG4KgsPkOUqdcEONMTTK23P622f+dE15e0SSWzUYuSoKqq2DJb/oaI2c
vT1Vi28rDxZglyzkSq+FhJXj2k3Z1uWupnZMBxhf1hEIJzbpkNkSizreyucnzEgVwVG3VeCzmxWv
EZ3UeLtsyHhRME/QF5ZQ7ct+qFq4sOcQ0WJ+WveDXD7xZ2ZU7VK9XlEp+KAWCyvVl6+h4/+1fthk
X7pYb0GiHFAzj9NCVGGvq+SJv5JSYqftz/HMS4mgyRT5qZO0RTmGvT2uYdsRyVZuSS3G+EAbVJrA
D6jXEiig5oy8e5ReH4Wk7jXQ8RZXYDuVyBlOFO/fWVVsQuU/ZSFZcv4AhJHdhh62vytyJnG4es3n
yXEg6I3BtwV4MJ6Ee2WkpbcFCdwGyVApJwNqf32cocM7/i78wYy07UzvqkIAV7I9La+ZAfqmwv35
5wtghek22xoVUx4/zfBWBl2Vt1p3NFPToAFUhiZnx8cJHk5sRvsyjpq3oKl79huJ5+r7mp5ihyZ3
bl6rBvo/GLMm8SgeTgENlGOZl4V2ujhBhAOmzA6k2oxXepaFShfWDqLlZ5RkS66/P8MmCtAfpD9E
thmjxTxoVZWAChiTZD3OS46qqRLcHRyZlldcHerepN07DaP8so2mRM89sirO5CDPJBrmx8YoYBEM
Tt3fpQHttRA14zxCvVgrzRig40dBjAzE4Y3QtI0kjqebSwXiyCjfFz80dIPIoQUH+U8bVATFBtb4
kF1f5TJYFAxLR808nNebcDZAASaF305v7uta16WeDwRZD4h47KKLkeJzt03gi6TGrzNQGVe4/Z2W
yzk36cLLo/F/uWW9rVZlFcIRNa0rfa4z2TwbfJGGMP+nCTlahbD7IijivNG3x/h1hx/sTInmq4Dd
0elLUZAOSQikxwKsBjeLv177UhC01IMJ+I8Ef9IAlnf5uNfhUJ511A5QIi6LGKH8ew0E14Ork5Mr
742/FmPJM9X91M/i636hVaZITyYTHTQ9QUoyIpb9qHdSBVoZugrGvg6Jy/ReIMT3qodGhNO6KOPF
wxBve3bDQZO+wRPtEmiqIN+TKMOjEbjJ3HZ948YKVQSBA3AVycfCfsmRiieBCN5Dffg0B0qfy730
HzpvvKlGcc9rLei7NHepPLzLYN+WHM9ZcStqJpIT7Djf3v+PgdpwiP8FjbP+skUJjFoItoubOoHL
o5QRAMLdMJ5+MuyZEby0cj3Qlr7pzlfiVJdViDglNe6AX0MHsZtfyGkfETODMjAXsT6Usj3CE7Dt
5xGkIzEhiAD/2ml4ockXPTeXVCfWjbP+UIszkQrVuysGD4A2tk2wDkqD2PyB2wtZE7IQybSNewzw
xoF79nDOSHgKLokzbj42UwINxaIhN3Rf4llQ5d+x/jvM+GwDpbb0lNLevjTsW7QgLIgqSN+OmLOT
XRVy62gAsEVxD+PIJBy93sPqmKC9Gu09HgnfIEf8NmHn0jvXdhrR7+uFyNf9GGnJS0oPEKu8YD4W
cI/gMFeciM23c3Tpd2fUUpgtbxBZPW3hBDm0HnyHobVWCoP3bGVlc+d/GJKsbKq03M4GNSbZ6jAM
XGmCspVGjT+XwMtu80RJDxxjQW7DkpIumh4emJTdDEg2GHZzYvYcx+UY1L1Q64G4ebQCNTDe0qi4
oh0R+NDCX4BwYDRB6A86D16I+tD7Vl90MrARUVKyAijwqiN8aoSvzMClQaf+lZAa1qDyKPKKY9dq
tgas+ip013tirwCHeHNN5jr/xpEwiUyI0eCtzQ5kLxwjMwmpltXN+J3UfXm1kXMG7fI6Au7PZazq
gesx7/WN8sGcmg0x7fVvqE6kiwHSdo0O50oSRQRFQhMMJv1pyI3qHjNVwZsc3/pyM2XnNg1+wYfV
YJqqn1TnUiEkwHO46GGvy8wE3e2mJEOCWSoHMd899k8JzeekzrZnXkw1CiGVel31bX9XJy6kF2Pz
57j5sLl8Hml+WAVs5/u6OSOb4SgGHwSvSSem8IFnbR7OmWhOyNgQfFlnWCZEUrPY/92FhJz1EE/q
SHgknqNH9rCN5dnfD+R6npU1pu4VBsDNsdhTjBTxoTxJYTIedIpUeENc38GRCY13E+AYPQmn9+B8
bcyyCY3VrA35WK/nd4nVp5+ZLaXtXESRe88kmjCd5DVAHKXikFI7Rd6DJVqRt66UB4lk+P8boARD
o/3hwR0NyAYLPUsyqbRPI6dVn/XTNjaJa3pcAFK32/jFZow8JPkja64Q3h+hB90JmNrjPP6sTehU
lVzIzEiuE5M4mBOw919lAro4+X/p2wqdWMMlgd1EwxVGeojzsJBbSg1c2FKJNYSPkgHd3aXjWmJv
t0z6/AmZNG3GpobtercyFJgvcn6V7r7L/1JZlpo4X0itcrJPhw6wpPK6LPeB3UMP6/yydZJlPhBf
HVzN6vqh3eGRSISwkiAwBi/bWxV393BvmRIPWYxKh6ntlX7NihzXSOOmZB3xWG+9AZt72gpMyBs1
39518fAAHunCjsdJGKMwRnZV4b+v03HWMWVAaLXuvxggJkPCGf0ZsxUc+lZeaLG5KXMig4quhHSU
tp7CML7WIt6+hBzyqJYY30G052armFHBSflSMdiU4ScYwTmjIHdvE98BHDvaJcu1CiyhpFFQU2Lx
7u3/gB86t2BDc8V+Rn/3cjzllEbssE3kr/49l20jg/wO/oWmlMxECR99/VpHPCZ6xmCpVFB3Wi6G
+lU9ewUIY9thZr6BjuTlo/ZtQfFmXwNoNr1nZTpX2Lp4GgWYlW8idvMbRFVZDQFUl8blhf9vEye5
ist3+537rjk2/zhUJZ+UfTiBFaLuMwhgD0PE7M4fcUPsjuxFDlly2whkPIOk/Qx8e3FozwaLZGad
UUcdavZ/NyEy0kTRtE2FQMNs/Ed6u3/gqY5a1Qj1+7CBpjKt5w81M4ekHdyhWaA44ssq0bAFzEi5
EQlcNjnoztj9bgY+Vfc9HZY1apVy80Mr46kT9zkSiDCVxwXEIDbfm9MPVezgNyYEK13r8+Seh12g
Hv4nkz7z1MkljKT+qw5Zo15pXWxDm3ffka9YwQlXPpuiKSrtvp+DM6rED3spDL7WHqDCc5cpPfoz
Kg64rWr4blMEcjwSy1tPh+0216xs608A9jDx292FBToc8dCA61PsJiZbuH9Q5NZ5WVKXOWJPqUbn
+MWWedsr9AdLvJuaLOZ0HtEAAvd/R1J2eXfBGM3fgg2basCeeudprpseLu+aHJDXcA+GWmEJoO7W
TzyZgAMUb07/TSZlUrxphNyx32B8F/YKazSEHepMn/pLCouAGlW7m+ReNzy/VWT8uLq+lp8Dv4yv
WPia2YIg0j1xmlxZM4aFH22LU5ABoui+P/bw67AzMmQQ6m+V8OWNewKvAtPFsNy+qM51/nx7gRF9
2Y1D0mMDIuW5AMGEW5c24b73H+IpR8aR9SeI7m0zW76/ZV+XypunAbG9SSj0/qcVYkMio6J7J3xZ
CjSm5vfzRS2ITQUp97dZCtyV1RMFWIAu5YjsOK4dAT6RNmoRDGrmPN2TKbllh6P5LIpLfixV+PTB
0RUTGs07R1foM/wzSxhTx4EL098V0Jkil45MP9/tJ9Mod/4OsrmbNCepj0nvjHUShbjqDczB/bWP
ynFWzGJDgCerMP9r7RvaTpbOvA1I/oMjCM/F5QQGqLF4R2ozeDa66BGGuWytjr1v12O+ch1458jW
BHbOTed8B1fsH9gjWv4bZbYGfDh7tNQHEb7zAjpjMGvmMJndC4FinlnICIMk4DoJURE8zVJG4R35
cSxmlgnS6bw0tfcz+okKAKkl4PkKkirLfVJxuSy27CdmiyFU96Fxkr0g+5S7PAaHHlhFGxii9mnM
uD9kULRtuZAC7R76WB7Rb7WrY5JVDV/dxLwELD2G0g+E+y+V5WIhgI+HP3BF6Gmk5v5P0HKgDPNq
huJvM+KT4GAavdIEuGErHzW5ndbczNrL/HV7J8QSvPDxwksQWLcXZ1fR/RA+kXXTjcxsMhPeHwPH
RqcXXqEmEv/55IAYa/IoSy9chxQ0xWdWFIEU0ukXVgE44988nYLYnEc5x/eWJ1AoJ3qyxeTd9RoJ
+E9JOcrpTxViKUd++yQjFjbh8zv55/DVliCc/+NlpB+vM5LDaZBRXVfY3q/a8lMEeNKT7rRLI4Aw
dwueBxBqhKa6Fj00WS3wyuTSHhDjLWaTRzhq2Zt+/wyRzobVjpAbzk69jf8OnMZWQql1P5fWF6Iz
JVVbF1rHzyuc8IJh/fsv2w6+MGT/+RXZ6SFeTbFQy6/3RckLqnWh50CSbnaIKBZ1bO0E2LzSkC7e
bcqhRqaBrgRDbR/f490TgJMv10K+RfI/3kKnD796j+CZCmqPkZKE5joWONIpZV/ic66BDB8pVYmy
EqsjhIByssEWBoogv4roco4PoQJzxRViYxGsb9gCa1LdhS6Ia+JKquhyuFTx4hBSD1+oSgTU8fzi
OejXMUmbZvBcE1Pjk65xid2t3Ebz9N+6p9JAM7Shqs+L6td87w2KcdZoLCs6w+dbg3eEUgvARm6i
9md+wo8Xvlx9pmR9Jsl1n9bqKx/p6K1CZsXB917ko6F9cFAV6srZB5ICLuAcj7wr926uJhilAFXq
IUqRvKXbgRBnXjzzq7NFvP7AZl5UZ+KqWy5ZzDqQmcJ+nLiWsa2QbvMlQqERMsCSiFrLWU5zkg/7
mPeWep1GefHjj56FOcNfqI9PQ6+9mGeXjaunwEVUOhjbNnB/mcsStP0SJmsK1lioT75yefx7wRdH
BnlxhTLTCYRVJsGybOYK94an5wWQhJn6LbmxFIothFzLas0zTlKsOOezV44KMVGK91BS/VIO38iF
ZhRWetZJMFibfliAVjm82MzTy8z19QcXKTVqMZVXEbx7Yv4dcrPfcIZ7PGETSdWA+vEfg1Sle5Dg
kBqSQ6qSMxgkrALsUcdpaEyQH5+kSxqUjdwFsS7xWhved6qT+xFxPe2mqqsrOCp8mk5ueGY/9Te7
RTQPCxj+ZiJP1s2/s4kTcDJAJ1CdNSNCn4ly9ZxeusTyFyr7HV2uU23j+coqSXxTulses5qi4l/U
RihhpbNIAqYRwrNbVmm6eBx0IGJxJEsg8BJeMHNMdocg51+/XFrN9sW9HtL6NtKB7W1nxEE5JQ5i
ANL49+4YCL81y+S/lrmAobi4s6IyF/w4qOJpmN9yDf+m4AIRurr03tNk+mOynMQntZ7GjPmuMuXJ
EVAoSYRapCWOUFoWkNHUYt19t33X+chbidncGsxo27zte+pfJBeaBZc41VDDmI87G2w4w4kDJRnj
hTFCA53kLvLPRPxZMqrsCWCMoTOekFBGGhnHVF9Kes3nP7EuU90z4aQXkKdsxhauJB5zXppo8P15
vih6uB9v40bllbpuyRpaO9byFYcZFD8dRs2sAq9bzKDMwCIZLKgKnGPC2g8pSCUx2KRXSQ6CznWK
knX4KZFjpi/XqiXoQiPXoQmDsnGeRzjthmXKVAMOxVfq0o1QzlOoSBhqgaYtVdK8bmeHEXZgJt2A
xQtupxE6QR2UysDPUdNEjX8BEWaCqVwBrUk8Kba3jYoVdvYrPiTHGg45xbMX96bGSQYhj9dxkyTr
HwYoRP9/Is+/Mzm7SJJjbCqh6FB+X6WdE40E9sMt0LiM1E3b97B7mTYeWlcDkmIl8UQkmh/XKsLQ
/chSsSFJwjlRsJ370TLX5K1X9DQ2T+eRJSO1+l/Jnit1pMR3saV3hVH0NzAUplOjrfrv6HJpTT7c
7Vpsil4CyhmrMeqF4EL5fHJ3f/sJlQ0JlST39AzismmB4oQi2NWN9jdTwTIZ1IoDjaJ2HasfVcgs
a/shXTEe7xBsCQAXxB7oweS81TymC8t28pCAcZymGGMv1l1qpAxNf8qI1B8Sgybvye/s6QN05w4l
AOUgQm+l1XkyYCYCMtUISgRJ7dFUj7Uuj0KN6dTaA3pGr/5vyRjTwZW2lRwKUTLCMJE3fw4VCmR2
rZV8Goh5bC5Sn635saumjBc4BmJMI+hAhycOG1jq4tv1wtX54dT1S+YBzKV5g/szRiKJRPQZ6Woi
cLuHBZG38nY4qUB+aQZB/ikPw+qUdqTaf2c/jWddJWmiB+3GNZEDOmSlGmrnbDzxqgRn/aDVC8oP
5p6lhxXeol2PI4mkit0J/oqKAwDv6QdlQEuMjn/51Xab3dnmLI9CGcEWED4j7dm7sk/uhjQLfk3F
Ra6mlyhtoQfFrCUFr7IrDg1KLFIBn35P9qe5GsOjqjLfiJ1v4Hb5dyRYqtc7YR+82lsnEMsz5Tkm
TWbxUg8dQS/GH3/4ayOYtpu3JZyA4UB8oDlVHm3TTUVPBYLHCsDxr/QWW6I5fcfAHb68D8B03Zey
GaFjJQRskYmGM9TkuNmOO+PJ+e4WjU7Ovgekvsr846aJCcDnY5ACl8K/KS62N8nbRHajCWrmE27r
9S89gMfkx8UkePc6IQlF3nCZzSu9Yd3RjCB0/RU+BSpHg4J5wy3Kflut5dHuij9FxoKsLGvwf9vE
KFnfOClLDItEhDThZKZsUPaGk9KsleKWMReHARO69QUa29yNMbtnjeSGt93Rr2dIKet2sa2aDHpX
YP8CnwtmTCzTgCghkC25+ZeyYkrh5l/Sdl2R+PbQnn0WDzRs6KD274mOG8ild23EgdkLZWGQQVPs
VurlhPdeK8SLGjcfmNumX8o9KlyEp3G1i1CHH/4QxgeKyAdptzG8fclcN/2NrMXf0KYl1l1I+eId
uifrngQbs860zZHBbqr3GhVZKjsmlyEuuux4hppBgkHk+QO5QAeRxMwpmqtRHItpagP9A34bL4YX
HtYr8f00+qyYq6ykmq4TBvZyy5E1xGlQbt0dUOOvNNKzwgqJ+p9FrC9QE5kN/6x+WxgExpyLJUz6
Bf/5pQ1uwz5pvX4H7zN8LUXxWnx3NpSQOzP0JDSZ9Px85c9oPbzdFjrK5bzhx6vpLwYpegM5X/Li
r4EMJrYwpG+YxXy5l8VF0T8LCC/K+Q0H/O6z43LR1yy0Klgp3EUrsxBcvk3TgZOhQNCLduj4odVq
wXEaotkZNC+Zuqk75U8GGq5HeX7rBk0DSJdIMhL3DWBhxMw12hIawmPZJzAuPTAnsCAEoruc2bIm
TMrYdkUweHcKdi1G98SRj4HbJAaibo3Z1Vknmt+NBHexleJ0HgTuhqmdxjzGcKVRXmMZ9Vu8Mb1S
KA5m9l3NkHzrJidUjMRLsq+KRgHHiMy8h56EfpjsJLE7A2zeWivReSx3nKRJjPLWu69GWM8WMZDy
AZxPFFt25RrbXNJuHHzs4byFcGWmzszqaGWAEOmhsLKS+OhYP4RzIv+lIYZXyOYH/TFE7LVEu1XK
h1aiZHfZnI7Fj6wpiBKZoTQG+Dtw5iuwK+1a/aXiKyWOLZ3mccuFPunXp0PAtvidTqDIy081nTWL
LWP8yqVY7NZBIC85Z9/KV/DrH9NLpYEnZvAIIFY2qsrXop5YDyLUShneX9wxNaUfIATLKqUaeUZq
slCQF5LUL/CSiGS1fWUNFbozVk00U3NYboEEERCs6o3VU/XZeiuZE2vzy5Qy5+SSYaSI24lup8gk
AGDTbyaTO431/qmn4xDdK5x8lR1NYpMfZYygZNAqV2dzNLoqlGl2jrX/qw0QpKVLhFPUgk6neTLP
Px5J9Zm8Z9NJ3vTsjLt4TBh2umNBgXd8lUcc0pvL5PzrZOrcPe2SeoJNSOFSCI4T+f0Yh8PGBSWA
/BOIDTmmWKBTy+VxeOsZxqTs/RLds/oDugxHFzB3G4cdAJxQGAPrg+EJAKRxPjUAP/+0JdkIqgmu
aNWyAPF5tPNy8kcMb36MVWQtTTcIChKnVZYM3CrfVF081IUipZu8WDfnxtHBR68ahpzj/ppQDZsI
daklUeaiigbXd5Co3lhSytIbHCilWAMDMREPekzgEVrooIDsypcsMGp9g4JA1GghqsUdt176sYOQ
sniphGJd+K5dtxkj1qJ6ymQjbi3uRhfeJEzJ/qAQ6fvSn4S6/Fy9sn+2Qh50w3uHmk5RjnHohR+e
h+NVuW7aQFW95TzlYN2qp51ZSH6Fr0vcigsSiECfXdDPnXY3BE/M3VymqcJkBNM4P0CA2IjeuaZL
yaIpvEYXUnd4TQKGnvgM1XeRNuytdPv6VWZw4GwOTOwN58w15lTPz7FsVwzWl1BehDIEMQ31Ubxb
ga66hqHOgG9BEUexUGYLAezUc8PQoCsmo2r3bpAAxjETGgWa02Jv6vnknbD6NafcL7UOMawvBRaX
iw/gssKbIqgfQJSXS6dTbeZbj5rD/Bw0s/8TtDNbzmchnfqHP8RetWbhkv0XWS3vn6j7ycQrEVmR
4YPY1np/N846DaBa4uW/obptIz7AZJYRen8UNXh15EBRer6hDnRjgCKrbcKKhVn1Mnak4JFH2Rlc
t2VLuJUSF7WOPXXWygpa4Rh10pe019uF/sQDn6crkp1RjBu0qgZzXKJC9PTPM2HALNgObaCgJTkh
eI1LWnx/MNsrvfxTLMuraHHsDErEvRYrr+op20BVFgGwHoG8XS51Uy3Z8pe/uBl0mSaQS6iMl8/W
YTjCgRcOoHOJ4jtaIQ72+VaKdqISwH0W6ejsvTi4MJh0ZIfpChz02T7LzElx7COHtflz53SnyRE0
1qrn4jyAjguLRofPbz6SLfK9HGoUUJ2Uzw+tXWrjZbU4OhNhg+TiffeC+OWQGKgf1fp2ezkWxcrS
aM4T8ZNHmdLBr2T/A+LIwGqs4/iQgtHrfvRip7+3/5l4OrCcYk3BPMBHGDzJ4m0nLk3OvqJYq2B6
30MAmrG8+VDwhhi6/+DgErL54pkx5Vsv4drw56aRa1cdkRJP/onkegRlfBbSJxU30bHkfRXyMSqo
gGS/uBodw/rlGaC80lHirtPR50/DiYblzDxacUcDIWyVHdlrnLdgn91Oq1zvNVkAbm53k6kr5vJr
+KemPWH2dtCwDA2WyNns7tZPPTC2sfwDKPVdALsqKaHH9BM8bQ3oLqF1YqLmkcM6axyRh5QPaJ6I
J285b1m/xJ4wbRnJZ/geoNrJw+gyPJN3PsANlxMtNgj0jg4MWAcB4PgqKJH6IxeU7hKayQdwYJZo
ov6G9JtNYchWWei5RiwDicxKP0ZzJHO+wa2MgeXOmI3519wYDQzieKSG8fuz/SF79d3OOtefEu6x
cIdpBSVs73kwHAe6uQl/E2WEEU8ouRpxW3ACoJWEfGCaQwmyPolR24SOplFZ2BWOKjhkO7AW+JEA
0KGdMFNCDnlN6JyLuVozWxhweIgqKi9PJ/59feOZENm5BusyTOrNczPLROqHFOOGhegmuTXMM5QY
CoqDdk7pDVMPADHxHulTxgBB4En6+NJ+LEQU5l2LnULNawpSVCHIhfu0YXDmT28c3iZFAQ780d+8
3AXOnW183M2JDjVgMu69BPY9flsuri62Fsg0Ddvk5VeI7e6PNyjcZXRbr6RVeBZSz50wFAziNo00
BNH+bRegqCSURSmLtNFpWUSuPh0H+b8zLdnJYQerSFCOgQk7xqErSzemKmCq/+oP4UqbXTis+cLv
36Hz51Z5EPzK3PTyMEBzWwQk/7y1dHuRAomsUNEtzoqXsmOSPd1PmDTLol3SAyn0SslG2V/09lAk
105NxraUOxWTBdJc4EshW/T+53WMBFSH/wZroiNalf45OHnh8vVY7cOqshlZdfHwe77gLpij2OD3
dTfVV7UE/uAzQ26YXAAGUnWlZ/6g+Wt7yZWqsnEGslbdLxHT394paQ0Mb2hix+yr4RTsmT62o8he
vUWPXS6kneFikN69LanzVtyjTaAmRONVIoMYqeQ4zAs+t/OzMQcHu3QXVPcY3wPFpyDuQDORteew
JLzx1QZGaxwLWiqSc7Ej4WBIwUeHiFBL/gkmsiS7CzOC8mJyLJjqO3SePoyw7SkOmofKkLqNwsdK
IA9BT2ZKib3G+dZc0rAtzhLOlARgWhkURTDtEh6m4akCtNSUJi4KxcZhoA96fjpK85QHGgfZRFiR
q5K+lHUjxdIat8aIKETN2VdEJF4Ux4ZfXmfH+FORSSuCeZkisQ442uXP7Q3LPlDGB00QQAvbnFfB
t9VuFi2iWwOvJdItb7Ll4MANAHSp/waIa1MM6v3gv9xSFQUD/q6enBtOU/HfKC2tvLszHIRYYSOK
KqJ1td3x2wX93s5vH55vzCJSqLaipLYLFNlGxXbpn4PErLitX3gdONzbYcFMSNLR+o5m0bmkyTi8
F0g2Fqs/mM/TWpjoCIV3UjBIJRzI2sIwiC5id5ws/ifBcYt/eBIQtmog3WHVmIJHnMGKwL1z17eY
NRIKxFPrT9h93vp4t2TOi1Vsd9zGDejZDrS4I5MsWYC6AGixMlruwd34KDBR+X1wjW7cSl8VUb7b
8Rt1cxEZkqlvTGg6hW/JrcWNlXurXay2KwnQ2EkXIAmG8DyNlwKLv+0PvQ2/dHmsmPgFvyvlybml
YTfFP2O5BawoG4CHg6Uzk2o5JNWppcZgpXGhC/ICxDBfpVk55CQuZilmXwTN0baNiuGOwxP07dqP
H2dnRcjmge0rNXDLEITUUxT80d0N3G0TEAOHTvs8F8lrjfZFZKyyWqp7KFz/pinau6PX6xhBz2Pz
+spt/6J0FFN+JQSAYWLqBNPb6xl4o/nvnDV8pjIL7rUKTXeNwg6PixZL9FJih1jOCg1BMFwHE3yx
uklsY63o1KwXozal0mpNMZtRUnynUhPHhffc2/Kd8sv4DL5Qh95CAAYZHWI6vYIojho0t4exSpvY
ox+uAJ74nRJbRcau5mNptNtV+JYEdXv7gJZjeU2me01jxUaEEwBYG0PL+GnrI1qtnJtrWtFMDuZK
ODUOSt5PgYylOQbYqW9VV1Snt1mN497mpSvkb4T5IgWaPo+xjRxsnx3Hcuj+EHOl8MAjt+acFksZ
FJunjo/fGeGHN8ZVvPMr6vpW45fpE/lcY9h/lRxxELFL1O4QdXesnFz8nKHtJAuCSa2Zi6+rVGTm
XS8jOHiBhqWoeXmwynO+Vcwjv5Xo7/KxaSSKprbD1oguTNPNfaZ7EcnnGylOR92z02SQJTxpGoM2
w0sIhLeid+JLCLCAgR+Nxpuo6VOGDgAqCFRPnG4nFM/N3wDzY8YE/PLbqKfUs4manpcJcvWlJRH9
bwg8+9fKONOvsOuDNoicck7ljH1AUMaRZfugjtvnCCTes+q6RiGSSSkTpqAkxkY3bjTkvm07y/5L
C/rwvpi+U75GdWJJC3trMB5R98gTUsyajEwCa7M6/prHeNYmLEOdz+Sbvtvm9j60RAAuGkibR82t
s4njQuLKER+SH2TCzIdBwYoIi6ImShsILQdwihKjl6ohV4vh4Z76Tcwl+Yu+I6OukMdZIf30hckH
t5SVZ+pnkqkM5SJsczTzm7AZGXihEANGZcxdvWEmYJU5BaHm09IavyzIY/sQxcIAPGMJZgD7euq4
YrXUUOUP2JcqxhTE+WkkwLhnKgL0karzlZNSN+4+aNIa3lWxh+SKfMkf09ol+qw3h0UHTDXbqaxa
7U/Ek18MZUmZVbe6/EYs4klOMiPTk4XOgEmht7QonQ4/U+UEtSQezOebAdUsMw6THv4+5LJpVNX6
SZKFK5nB2emQ7OrMBP2Q3sE0HkDtAj2IUsh3YeA61zVhDV/T4ZlbmVj2y39hk46SjXX9H3/BPu6g
rqqIDkWgWIiaEyN1RdyHZ4q4R54WsXxUBJJKi2v0/YKTVXNrpgwHVYGI93yckAC4L7oujhjOIT9r
+n4xwObXiqu5gqprar3WFKKBsDQAPqSOg8pXZaJ0zX5Aeydh0XbYfEarTVxdgSzglbYEbDGsr1Nh
upaw5dhQW0W6IbbM80IQQr1kdOTKr6zjVrhi3r3cTmlIXKSA0fdP9NAskZ2tBpL6BjK6ZE7eAWKQ
uepi163lI1dv2xDWy2lit+dYTyK11FcrhnbLtjcyNnI9F6ZcOJYMgF8MAHU1zpjC2joN57enzFwB
R2Uy8Dfj2JdDxz3mBeRcDYM8OR8ElgX6Q39gN2bgf4XWsFlZTDlvwXWey8IWa/EqLCAPrOTolHO3
fbZtmYzGDY65AsfaVWZGwSZfdL7dEcfSmIqRNLwka7daazkxcIlVR1xCnWyzh1wcXQy4aeDRwid+
87XQBQaZzg8ZfqVHAnC3jet0w20IQ13CsjIG3czPZTN/dIRffM3hP/hRi+UZlSt6AA/d8KayWt5y
9yvuaLHB6ZH5EOD2HTVPll+nEbyof5Xw1eznhsXIHw1Shhg34SA/OybhnKnoDT3UJYwBoQF5jUYh
GUHAnTetHTaTffnhjJWR7QsZb/zyb3G3SYiealawVjFJVv+9zKhEZvq94xK7oLIDlOESXsQ0phTx
uewYEXS8tVT+RpY7SLiQ84lxv9SGCQvwVlX2PStmdCV/yhgEdbVmO//bvtZ9Bt6PU/VuTjSGZh/0
4pyQwZSfjR6engFAEczGjmKkNexOdjohWE3DAUeqEbHo+F1K2gIKKVeOAplYz+BdOOMaDQDCFdOv
pZDDQL1I8sQMDZY2+Gh/GFQ+G8oK/IybTZsStyamIafuGMJpNY26GAKsmOAVfxuuW24MIIsW2tke
QhidWfJuydsA+X4a0/YaTMdsYmjeaSgI9RoraCnAczjd8fR11N8EgE34uL9z0lXcZ0sw43awK7G3
q5Rw8M2prtL1IZBRhwKGRm+t1mrQLSQXb1MjsCFR9xbXN6WAbdeI+EK56BpptLgMScyN0PM06NZK
FvAfBmXdE+JQq4RbJXUQ3CgsmSaeQMMpbX3rzewqX18nPYRex9yiJ18Vc4RzzCXzjV5T9Zr22NmN
UCtu7OLUWAQ9dCq9twnY2rHlLxhtHodVQ39gkIVKcsKYXLsWqD7o1s0hCHZLzTrquRKu3LNjlVw5
7KY2f3UCSG/5GWBi/iRN3OP6OTruLlWSrCg4yqM2kROc3A6t1NFcRflxI9OY+IOU4LcYnT+JycHr
dSxj+8pyXhXbulennF5trHH5nz210dGKW1Xqh/8nmxVyfUtlkITcueTy+4Lq44MuYswbmZjsznHk
y06BrFXnTnIbf24CAQ+x4NDhr2iyYARsQdQN9etCTnw79Xq+csJYZfoGbKyqMw3M5OKqkJL2+dJe
jJeRhNW7H+78+ocwrsi+mod98oGRp4Akhifh1CcXeFtQkdha0jRYCMiBr3YpLMKnMACzC11barlT
V6YqCz/PEzAZ4PHWy/IQPVtyRXAjHmfLazmHMKrBZ4TPuTnWNeNM3g4SIkiN8Nl8zwhQLyHDz0pq
+/NQVmNzDjvXnEDl+Yn8L2j8F6zsxptYzwN6D8wpLqBaN/7+qszQ5BrTBagJSdgO1I07c5fCC1cS
TS2+7nd2nciC/5qlhjU3Rq0QI2+9IA6s7S/4JihTbDHC1VO6IvIP2VYo1q2VqCzb38LiPH7KT4W4
Jp/goOUkRyLEDUHi+3Tz1OP5FAFZf+vj89CRFqLS7rzNFFk1jxWLXOF0CZuwSah8MvC0xHcqqQHT
u9caoIgx/VpZPCUDiftzn75/LxgMSEY8Bl+uJrBseARVj8Wwo1pQ6ZCUMf3hgbJdm+Hap71Nphk+
ry1B6/EzO5WrkWT9cs6Fz+QpOg7tble30KdejCM2QZTKF58/n7bEgz3FRrAZ8HpBWqTj5Ifq+Kr6
sjJj0UDpkpIwfuU0HJUxIhLcZp98NRtY/VcQZu6X/VSN7cklFGrulWyWtXQFME8Gwr+GHmE7gNLV
j25GYWY7hATfG/wf8C6CSLJ5uxXmtiLE8Us2zrOZvrUwKd7CZayM//V37J2GwXu/Ge+fCVmbt5y6
bQsqQZ/BozNkUgQVQCKLNPKLVvBbv7SpjZXV9GwIbGURYPrZ9Iu4O0O18K9iyCzE+/1drjoFOJ3B
z6TfEpTecZqrWmqhjk8ou2569fAsYkMxqgPJvdvdiQ5tjgJAmp6LrL77esN+GK1ma5wuOCKJsaIh
C1qwPMpOpD4fShqG4YyXnBljRN5v8zjzU+E0toqdRbrVV3H6ul3kw4J6IK/DSHk5l0IY2XvlPsp+
k6inj4A/ku66ERpFIXOiNzbusFsTCq0EBfHwznri9pks9R3X0XDj6QrfIvMShfHc5CE0BHdcl3f8
JLwn9gsCaAXG/v4JBNuHgLTdF5odrsMeQ7mKtfkcIo3DkAaNRaI6VwcNxvJtTi/5iwZ0n3j4ZrrH
QiOxy5OFkuGZAUsbBUhwPlhW6Sc8ytqwZKh+sKZfNb5owUGg5h4Y1VO4c5QWY3PREeaS6DlWEiQ7
L0B2ugzF72J7LMQYb/YadRfIdC+dKo5Vizg1aQTgZnbU9h2c7bkU+wKW9aWJYEeE15TfBA7X/IRP
tz7OIS+V4EJY9IRkuSZjTT94Bnn7pdTgKnrQgtKH0CgeT8r/LC+eT7mYT4Z5v93Uhdz+/anhVui9
tTvOGQ5PsJ99dBWZG4ONRbYetZgZ3clVutC12HBig8Lx1rrjxSgmo1kT4HfHEcuXZF7DHfojbeta
vHMzRIKlkBZn6L6+P+jzG11KLoQVrMNNOQczCJC7eFPtsk/E/kcSPs4N+X4l5dtyq0/viu/XDad3
IkqvfN2fK1xs9DAJ7basxdioE0fgDYxbx3Hd7w4dx425dDtYh/F8zi8aobFM51nDA6b3rpQ6gkfp
Va1Wll3dgKnXmm3feUh8UuLX93cwq8FpWaaxrU0h7LVMQtjxn4DlWAdSeHMXBnYulAetoHSkTeKw
frb9W6mNB5Z3OTUeMxzJVqRaaKWXF1aSMgJBagLlfiyR8RiBWEb0UJmQ0Ia9I5N/CGejMwiJwuT8
sgACw+LDLqjI9viJ/5tK31zqif9yRhxFwZZD+qKMSITdGF+cilb6bBY9fxwLhaubyxF05G+f1aP2
O5CoV4L7837yA9otJlaWo9bTde3hI1xtSvgDKhaHgct7cptOOa7Ef6KO4tmryxzcJdUesJKkVB18
2bZUvdCfF450Dli/MM+FqaVHUrknXxVDPp6D1JPmeHzIsvfX07UKNo9/5sdtpAbzQ1ecJfPjiWeR
r2E6pHJ3EHY30//qbIvUd6BKSNB5s41MUpJeyRL95wXCa4ER8LmLWd1B7rfE0mCw2HF+KtjulP1g
9hK8W1OAW+QOwDN8kXNiAC/Tt8xdGLf4N0RGha+pRDX43oct9sALYpjYIi7xR742esF5zHqIJOID
NKLFcQ6p1qlw8/bXs1YhyRY265juBhcRXHjpUv0MVq2fj/UHGA0l/jCBSDatS64/ul1v56dlx8y/
tnnqpyS9zgQarqYek+qyWvDxGh0qkp1Xaw2A83OKhJwR3ArsUyUymddqWaYvbSEpBKVaryZ/FlZT
BhUts6RAKZAWJo+MFOsnBhkK2ptAYu2h6kueqQUWZjt5Ydto7TcZ1JMRiiR5IBenrwS+Hx67dHBC
7Gsk7Pyj1CxaqDPTALdvFCPGKXzv0HwamSjCPYEXgNXhLvOCbwgHQ262GQLgk8QK9GntWAT2djz/
wFnT0LkyuQ+RFUCyijVOVdGGSBcV9ZIqkjBI6T0jLjTnSyC+0Bkf07Fmj0dpAQlLCHpouJhUK/c/
NrWIGG+tUl1/lb4NgLBmCjriWlvi+FZ/cr6jmHMWOFm27NJYG/2D2CzEdgmFLkVH6YAjxqOTAXhy
bJdI3QYhPEwsGcRMEj6LcNVDEA8uzzlvb8cd0SyA88eTgxT2wL7l5F16jfkpqYzn/6UCvWn/dd1c
L/RNA8peoWPw4QoeEhkU6ezLveNROKTPmxmGfrAevbjkdQ16/9Y3xKfJM+PzENgJM4n3rlC1VSJB
FxUKTUoVvK7ZDCuZie+HzsSDKQrt9fvCU7KSsEHoznjORm7QvIMcBoIlIScxMBImpTZQdfgl+bFO
BIKz5JZ9E3APG4V/iDZ/0MY/1cssxBPwhAtBkbyDPQyqSb3wqTDbWGq39hx6Wlz2XwPyrwh/di6f
Ncpl7aVKoWS0SXWZvJuGTuHuQYCeTzzPSnlYZz/SxlJEh+yUnxJe40cVZEMVBf9hbEkyUV6i4MZG
WCv9XzFdE4wZBg5WMsnrX5mtzLGccZCp3IFVEhrXg4oQhw3OsiaG9dVOqukfdwV95Emp60ox8SNw
SRlRj41G2U9LYVZo9NKfASOqd6UGe0p98e2PPYMavW29KWUJDruXVg7BroqUU+kSiWGVBq+eY1Ya
xWDIjfKQO3kbZ6OyjxioQNAWSROWyza3tL+FW0YXu97FZiApPYSZUVcAB2Io/kC4gG2veiw7H7Yw
u1vZLziMoHcQpKTe2TynqrrpHSlewFZW6HkvXeip4ptaF0wLpgoinzrZ6zVV2gcHYUdbPsbZ3iX4
UdwhxiIo1ojFotLhIw9KypGTA8Oc3tNiw0tkLCPrDpp5duXoq0iXf9xphed3Kw6rB/Sn7nBMDP6P
olQskVWmeFmPYGt/24grXmu0ckTQIGmYV4n98sy7ip80a7BWBJGLAlnW/tgLg8MoFbUNz5LVxnAb
ROlOpNTca3I86BGkPYpCOC8lXLlt9UdYIDV+OekPu2qCXv6GsxIEWX/uigoBVFDtLfzPuuD67AWB
ScbK2g4kDM9/mOwn/nj22CLMcWq5dbS8K6lgm/MxTvaNA4tOMwyDyKn80MnKBSFn3lUDBJOfQ1fT
BqmdHTkeLfSkQei6KxohnNw8lCSZITolsB6/nCRbCoYxW8ZhWZKS5Ucsfajv/ePyaFRv0Pe2v/8o
dPXLc1lIxaEiCrGqPBTGowOcIlA1MGJ8ldg7ZNd172vF0pg0Rp1Vi9PPTCJEL+aXP5/GhbBbnAfQ
pW2oCG8RLLXNE1krQiXtODVo6w/t/6LIDG4nFwJGpVpRx/vjdQZ5xWMan8r4CozRMSClxPvX1C6H
/zvpLUELzG6M57P3GGvrF0oZxYx5fGbiQwM4WkiCEvsjGgPW0+MDlKVpZxAmOLSuCfZApzLGgZIl
vrNGL5i0VOgh0FGIOA90PVOmfp7tczer8oWgVzzMq3MYsAOy3MwOgP8fiYXDLmRsVC286lf36QCG
Nkk+3/geqBlFYzFLOiiQ9NFSixO+RPTgvnhEtAZgxC83jnu0Ij8S6NrQRW14rgzqkMuz+1kJ/tgS
7ihmY2fQy8zYX/DMht/YhEfVBAOv1I0MFHmXoMHK5HgoeYAuSmLoyIW+NeowE5hKcbBGLa/tP62c
sf3z5lgjenqEZZx6X81h9Vlzm3NktlGuRf14BGlYux6SLyQtNaD56z9Jj2JqiURbvbblY4J+q87Q
7E5FfuDc1xOeUc6/qzQSPo3pSEYtGA7Qr3A6tfmmZ+aOfum4cqyOf3rqlyS5MoPhMfNJj/7b+uG9
9yeI0haId622j9iGUu/Hda+8nF/wB6VeTr00UYkK5R4/9vlfkejKdz2GDRLURZg0IvfcYNoq9ZMZ
wZvNR7pTN8h1AqRa6bpKrr18zLcIdoWTw8WnUB9r8GOuvD0d3Jfkgg9J2925O6gHFwS+QW/+7D1Y
3Wdo1OUzaU6JEdQ63q+g+F2wjkzkXmnSZu50uk6VlExrg6tQIaDdJN/GW6KI768Css5buNny55xP
qm8haE0HzhIoj4bJHwXJSXDHx1VB/H6POJEvuVaGuuEfaP8/EGLEjCLmGdsquWgA3R+z+t5GrbYO
TqYUPNnElUvx98eV1p3uCpDjeZnvk774Vno5ZuA1DMrGJt3+KEPNCTFZgtflCcScQnyrn2iR3J/S
ivIHel4Fo+7H2+naPP0shw4p2m6ulNziMrcwqZdzjs/30OdghRMv2n8dNiOHqqtf1eJtuYpJvZiM
/sl2QaIfKwwcWnNA5mWCMJk+nW6oUzLnXguYJGpDvkSIrjZYymcyzksi/eseNgJg8Ogg4ZI6Aaxe
oFKqxoABuqq3aDqTV67JjHMnBTcMsfmxsr1HOpBWDHXzIxTqxT5Gmaw0UxXmbQ/divKrHeUq76Rt
s7rfKS/FdIYXA5iyBaHmEu+0MQNhsSTJmsrumSvFnJQSYXV+HI0YnBloj9ZSBXVz0Hj/hWFTnVZo
wdd/gXtD0FYZxdUfwFWu/6xjp5h4Vr0iu4OdS4pIEiLHP5CSOIcZcgjAMRYGXhXSe68HL92v8rdO
PXNiz4FVQ5T5egLL5ULScVjPbTBw1o1Rbxoy1KCic7NjzfWbDFY/pUO9+n8sanH2ILTEiny8jCdD
Im2vDdP154Vxg8B228Hnz4XrTieLIKVwHymxWA4IwArRjeL99rIiIstEWE4UBmyqkKyvg1QemhT6
prYUQ6PQt/PYrZMB+L76ihXB4hfAiawNUog2zu5g7iuag1kKvUEslIWSIsntDIDtDCDY29t4MCrw
0BEDRad9hjp/tFXOLFBmDQTf5fRt0dKPebFULmHKkxvnqoz3j8Wug3oham567X99+I+ALfFuJsn+
++KKlUu29/X1JIi1NYRoQvgE0oPoi9odL1n92Nflygv7npsRFQ0JcV8g3x/vbdhgdNarDJ4+y7dT
lbDdjzVAyIkZEPkUqF/100GtwBKSKlmlVKEXURrizDMjSrcG/BZxB+0K1+0/0ZKEHM3NFa7qCPV5
UuERHDcqp8XqklIWmgEuCCpzo5a/qzDvO11z+ITCV7qFXNt7NqwTyEP5hQ3so1Lync5b2yiu+/XK
3elons0x46p1oOycwOq2+CpUKDKnfkdEDOHjguC09XKR01dFq02vOvNH4vGVvxuL7MUWV0+aSGQl
Tlq2+dr3cyXNbhW65Krpz4qENaxCcjaQcCOXvGWxj3K7oL8lXg4gx6LhNNeChvoSNJOoB9OBb/ke
l7MK72llciT0QqIIMpQbjXxXjmcU930BcAbKHXmVIuL2U0eQQosbL6Xdh5IjMHGUYNCd3sTYnshS
YPjns5ztz/FZjjwcyf4shB9h9gey9bNVoEvfjB02LezWdAvAtORDNhV3E0BmQmMUh+E4JdCMIT65
BlVSIE7WfnbW8x7FmpH80kcSwHbO7rQydbjGhP2snWhsfVhXtXmYw1tuF3DiJZjX/H9b/Gtd1r0o
C+RhFZu1U6opSdQwu7sSKjNZfVnj2k8HDxKjbAJZFdxI7IXhR/GTqnTeF0+5uThm5rKnzOsGzeHW
Hr3oetA7enogPWcvJyupmdtB73o8xXZY47UPjO+IZY6IckkHZ6sg5MekPnEwjV+xnpzEJoErur21
FmTpglX4J1BXxcyKfoFBtl/EZFxU3oU9r2+6ePP+UmoL9Jempa3yV7Pac1bJdfX/p1C9A+G1MuaX
smb9WPE2PRHwX0cAn4TDGnCKJPfjffaA4BkTqRjeCgg205/bpNkpqYR/RASejOixaCuwUQKZKGEy
TiD4X32Vg6afer/BFT8c++IrsJfxTut5Swv6tkOVjzoudyXo/4Pv/mW9fzcqD/Ba28fqutGRXdN3
/B+mhVefg6hKBUuPVeqSzEjDsOxFqfJ5oepy0NHcb3QjnqF/A5VuG34S8HbT7aQKPv/Qy8f53hDu
FjoiFBhDhlIbKWyxujwL5stdEyVxoe37KPG0bnE93GHx3t++3k0rcrHlGAv05M/Fn88idllKG551
PCPz0+PlgBfZZ4UMr8jim8VCL9gx5gFFKEO46AWsH9tkg9sDYyfUoilDNvDW5sXpxWzFWCmtdZ0O
awqfjjKXJf5SLCEQH2zCbMo6tmP0OnPidiIM/P8ZHMcy2sibdVG8TKIKUFHjCe//KGajT3l3Hzmc
ynjgZxzN4D90flBupaS0GTPgkir6tvoUUOjG8zCT/d2c/dIM3ZOlHHmLy4VswsuW+fVT2Pjfw0Yv
bRTIuQN0FEPt4RyVhzAAyYAnYzqY43Q3NjMHXWGTSjx+iWIgPoNi9X08vN+OkVyGGxHUMDXk4iaE
Ai6jnhsGGDOWywhkSMRXQc1F4op6h9hNdzqatILqPNyjwIVq8j9X3yuXIaQzTUeOsHTStx4811F3
bGPzxP0NX8e5gy70Q9zhbBXGLjn3ojDyGwzlzRHOk33omMjdJC8hSW+pqdTAOV51Y9w7lma4GP1k
YQJhinSQNUCXnPs1syXXST5f32GHbOa4V0/yGkqTh6xDIf6aGVkuFa3oqSExt9KMuW6yz2w+g18T
/UjPXAKXaNIV4IPDrLPvKWVa5X1Kz4kLxRp9DqOuv46BSKyOC2DCubnzCtkY0m8DG2cPI63neVED
8TlCj5g5TOclf31Hii/TOjbE8H2KN87g+4PWGcdNkQptauwgOpm89iNR7IYEpoV0XvwVKw2cjfr2
wlUw4yf7QVw4ruAUGhhQFidRqaP4ieNcIECc8aPWj3gjHjDFIugVo13yuZwLC7sZgtlln/Xenm4q
DpLPKg3JcNHrQt8WLJLIzGhuXqOgAULioDAuD2MfGQfvlV27mERbw0T31j0/PgVfYF5Ei7gSChQC
wTEHNxOmqeKBYWMrmXwRLUTvnYz0XL/nRJNoR0gvugPhAiyEmv3P4+ZDetKmVoPvzfqs5v3JjV94
ITwmbZ7rF8LuNwYUHz3VuVvye9MNpdEnf2Sc9qlpqM3igLHpxs5L/EE9U6J/VGU3azAOndqu7waa
1aR+nXiEhxOducldUG9t4Z3OCcWIWFBjuzxo/kJ+lrFJchNsvdGgBfnxuQrohWb7nQgqac2+HcNq
mg3yxj8HJVUtuRJhwxgrqTE16CHTsJHQlzteBi5ylX/yey+G3keQOerq8g/gQ1nKhvhGUg7xthCn
pekgulwuIclAbg5OMCnwrNKezC5gFzLN0+tmpOO9PuRDx9YJj416/A3r4PJHpUigzUR9rm5iseH1
eoPDCrF4ZgP3i9D7ynBHsDKnZ0drdeHVezVEpJuKg0i7qlHCO9XErCpz1CPkI2FiUmfyVQq6utnq
gQejqg3n/TbNfvyndPDNyN5vLZBclEtvWwHtlVeYNlL5IFgCVE8zkdIT5qFob5zDYVM0C7fcN8TI
cDktoAVD1My2kBcdpcYpiwMKbFHZZlDu6VUVeKSkot5yLabAyVE8NvzI7dduqTi5LtOWTTpz5bc7
XNQzmpSX0d/NVPvATn/MZLys6FDd8oVdAOa7byuYkC8P3dsbWGuEl2CEOOACxX3QDAXcKUVEGLMu
tDltLIffNyIfLoWVyQuqqFU7l3FReaMT1s3tFLSVR9XvgPb4JFZD1oR2dlOdtm7d65JeUNm+Kqsd
djGyyFkGmwEKCR46Qkx1yqJh9XDXLCMepRV6ldu6YPtz2h7Uy7cx2wOt5/6MFVfsQVp9Xk/MsmVc
o4UHihqEqtOr/N1dnv1Gu4lR094cyQtcvl9Wur0qwK3F8GHofn472x4unP+LcZuOtdTUL6GY/RZu
IsNShWg6oXQTHiV2GvftzLxDStd+7u4PhXe1RpuFyANNphm/TCXPiXi3/sbC6MHOWPJpxAlSIWsD
ZxGXlRy1Rwe9oGMrikvQ+4TWxfMhNsOFBTLcJevngul1rIozlBsgLdXRKvG5IANxa/Hyg1WDp6ZT
1DiHunlM1coNaJRGyAP3bv2LIU7Xc1dl4O+OXd6nUWfhagorBbh8Ney3vGUY8jMOjM28cBgmrvlx
BXeChAJwt98VLnHiVK3aRlA2NLtwYT7/nut6QoyYJ8PVCmCceZyeDTN5jFO/kHbkUdZ6qOBL8wPn
jsZ7MHT0ocTWnmXY/iTEk4AqoufVWd/V1qR2i/MWSg99J/UfgrHIbTWM2WUD8BOZvP3UFR91gkt7
nNacCvzPhfDhUJYhwmsc2CnN0bsxSLXRGAPJ2uwfZgIRdiKHNfAhNHBDrWApb8V3G3QguQ+Ves3l
wI4lOOBA0Sn2j/lUcoePBsr5Wt/mVxzf8NagpXQVRMnS46EIPYBPwPmZn/E5asfxEaIok6CjYbwW
Cxi4rxR6OWQL86ErxRwY7sneuCx1i5bQ1+vSf5u/46O2l/btJXYzuIZMv6lDJ36Ppaxra4NiaGMX
24AbQgh7vn5RRK1Vxc10plMvXBs/7/h76a36tHELuWkG1D/2E+hNKb80dgbuwTEoOcVZgo3IgkuE
WaeQhI7EP7a8zLrQR7ANVi+cqJGtMMj/hYkmAd5I8TKyzuzNtnI91pdeJHFj5j4LQPv5oK5HSMBA
xIWf0VF/kJJMfUEs/2sKigvfVSkxwFNV8a+2dUAMduePzXrRzQg8THCqZZvlI4EFAbVFqjRlL8p0
3rctr9nhSzwIprdndZnXwfZf0lXGDaGfWHV/MUM0pHXNi1BV0uDYJNB4HHGwjprh1P7EVeVNm0td
nCEkpPxvlfn3LSiaP0NCoRRsJpbXR56Tun6iDykj8qUjF/fkPtvHoy7KaH421pZQRge18Zsbrrrx
nInPY8B6At4EOpMIANPkIK2/MlGYKN4Z4mIC+CIvZdAkDVlF5VvOrapOYovcr6YGZLflC3E8V4sL
aUBDddscCBkDeomWdq2/9qJdd7mfOnGGik8GQYT5dRl2Z4G8XS36fnx6oeaG0j0K+Xsc51XxZZ4B
O1JFghkkpZ2hK0lwDSy5Xt1C2prh76MLZdP47Ql2EeZkuWbTSDDJMgfK6veCByseol/QIdGBWpjK
5P8LlXYO+0JYfICVzWYo3vbafZBV2nZgDJR+jZ7GJMyM+SoDQSnDBAgwle5uZXftDdImpetSmXAj
83q+lclU2ASi3S2KwFQz2vpdCKa31RdM+jFnOJrWvxmEVlEJUMTpKsMKGFqnsWs/KhCdA3XiJLL7
mxsehw9IjYUSTAfaP6ZDN5wlTgCsCN5IxbxRr5+z7vDLZvcIOlvXE9AJF5G15BXHwDNSpeAFROsb
xmA0ZiUI+s214soNdQ+9IBLoSoyMxIQpKSL9yIK5okifmkvcUlOvlNLcvEY284mhLYaJa+6N6KQG
WPHk+8cffnxLI87Wu/mdLNxsXWwD7zx7MgXTjf7eK8jQ0hs4OKwVU3ht9cCU7/YlRR9K75kBgBR8
xeB+LKjCNlBq+imA6WP55aMIslMeQpxa6Sexab1g6ZZV43bMTOXpA5YHcoiR/O2dFh4dorFHEzTe
Q9b3yIaxQ8utPMZF9wCvSgHEVvP322SrCwkluAi3IlLlG0M3x57T87RsLmVr8bPRSBpQpH7WMoLY
N9JjB4h3dSLKo+w2L6EvEH5tiWHEWJqAeJKQTHk91wjpx7qtmKNs5uxaL5r1/ZT4vnEKlUlyDDYo
r/t8o0xIKIVHdHJA/dggTXGUAYKagLQZZb47ta3UWKAqs4Ra4nmSe5sKPbFnSjliqT0EMDscN3nF
lGgW69FJFcsPnUBVgQds7w9XA9R9h39+wJuyMLqVyS9ayIPveweIcY0oi6JLohQIZfs2vY1qcxCA
qI+eUjuSjImNeQUro1iKvVZ9jejZN33VwHL08rSffE9DChePaN/YQaKbKOLkPYAkLXmVEjUwyB08
GupGVput3/HogG2XgKJ1UVeAiry/dl8X4ciO7vw/0KXVkPOjWyo049dkoFmNjVl0pLv58BvttHNn
Mwmscj09f8legJ4oInnDMXRsKXbJ7K7RNiTeQrSSt3nppHQABy6VzPpz4a/jjgzIixlDrhDmfryt
vZ2pI3jNrArUR8QwSHRps4YjoYa63kkqMM975oNAf8jm3WEwRK9eWzDgUE/QFBvAjm/8yYJJ8EF3
cvnxS43BA6L6m4zgUKAxoZFaB4gWo+WJWzyRNijmk9qfZ1n488nrlO8gjR7t2T+6Baxj9JrVdZwh
lNs3zE+YRgpSlsDXE6zmQsj8VWPNhBHNa5SZf28sYLPjY6Ox2oz26gyyAlumTIa8s0AhLjPR3vtZ
kJSi1Cs0Fce3IYy9qZz5k6Vvbi84d9/FOtEcj756reDVyL/HIJhGUyMZj6fMxKtlmCfge54OyK0L
e7o16s7yUDIbSa1RxOfftR55E4W4c6h7gbVvtbWlNBD9qEnJT/4535jP+iVyfYJzpDqZd2DONpKx
iLhws9MwCGOfp1b54ytWHiLqvJ3n2eSkxsU32LueFKsPo5U6lD2MwtGqMNh+3IkmlwJWHXzr6wGY
ikp0YVT9cfydHdbYO32odmZXB60ZfP3qJwR2v+zRYeGncGK5nZdPfSxQttyiBtAOp3ED6XI/UlRr
7SYk9hhlqWjbi++ZArtuknXuN3Nl5h3UDOTJEy7ZC34iJyjbEZjiI7VvkZrq3OR87cgVRgRIQ7i6
4RKtpMGUUbEaB6EQIwcGe/EII5y45QHstTM8rW8oR4JPMOlhCvSfJEMOH9KCg+8EtXFw7oqdoe66
QthCbjbcEI0AEcvpsn+0Nss115hWaar6SeE6WKvgfEBUXcza3TeAcZilBWoBeZrcFh9WaJDp/AiX
fKtv/ErKORTYTR4bSz5tjOW0Xi7IBySQFuSfqK/L7cerkUS+0xkz4bzGkLgkVI5myAgo1Mw5nLjC
xaYpo7NSi2s4WtjLa5GSa/sCQKTcf+qdyHJIQEiPUJ0Pf09hbdpGErCvQC0A/xmLmedABZPgP7Q3
Glmu8EvGyxLKvNZELpVJxkUNFMw0dwebLHrooQi/xsAP7CCsR9mly7umYzCk5osVIgzkc3fGEFbk
ib1Zut45skHZeYPhM1LLCFsX554+xf+Non8t6f7AhqUSKcrCGIqoJ5pIz/bVsTAPYx1I/6oRSUUp
JpLgbeMLWYT19YRfsP8jHoy1Ud25BnCCynJ7mNXF8eRvofhe/mX8zGrY67g0zqoIzU+QW0us1HGi
vFg2UO4hXntG+Rz3fEo8ILpgiZ5Zy9hMVrh1bT9YCyDOTaFEqpLssKlD0CmiRAftsonUR011Aein
6wsZqW1xNUx5Hs0urpXRj5TYNvKdJm7WBFaaJTXHxroQrbuEQ2S+1J+RTEu68X3agxfRDPGFJMbs
qMEPcTa+t3jD1zMXx9pD18NMgot0DJiyQXdnxEINTtC6jA0+yDyu5FDATFjQnPCic95OmAT4qg6H
LuJvNCvCOwpZF1ZTr81WsynD9/b5z4skjCxU+7CXuOVDKVns2FXpvKWaL3EDelrdy+IECkcYGf/q
8KpRLUzHmAL9puT65T5btmXqPW5nU4CZI+kPBzmObdgYugGWfinPNVIQwLhlh7ZgS2xHw/fs5xNw
fGeGJeaskwqz02Q9is9cIefNUFLjNLOFNcAKK7i2zStDJjZiXnCcCQu/JYsL27q3k4fFJP3JApDK
2rz+fHq3PJn9qWXyRUqd9cItHtyHqzTIAfOKdSijjiO330SWqcqIu1to1z4R/CIp5VIjf9D34PrC
4el1dtPno8HS4uDI1crm6wrirEEJ+joFm0hxBk7NtGkKfSjajs6rH/ppB4FXWb4MD8LaQatouR6h
UBIAVr82Zq7RAfe5ifvkH8/xI/wjTU15mchUXyXg1+vZBGzfYMN1GFg4kx8i2g7oT2gG6h+LHt7n
Wx8nuSXKoCL+V4Oj/t4M/ANx4S8QtZVnVvA92X5mzCOS0z5k/H5cCRM2JPaNGvcSi7easnQwHWDv
myk4gNOThMmAlqpYbRWCpXTkq277ChVDZzkK6DOe03+3GQKJEZjDvrgW1YaAP6BFXRJQZA9ItYuL
LHiho5epkbTJC5SB9U/0sbamM+2m3ETYGrgpNerMYOCzzi2X6AApbhYFEae6eIVAAe6Ff4bDaAFZ
5neD9LULj6zzLkAyfegcphv0u95Y67KuP+6/aVSdniV0yWSdkv89ynU4X2/eW7eMYF65o1mYUXsJ
x1+J2oqHd0UpV/fSu7JFpXhSka0bwJ9oCGIKXWCwen9ai50F/fil1FXcPlVW0UxObsqcWkVMGwAC
ThgrQwYIFAK59L0XrW+T0IPjKChZ9RWYk8jl9U+vAq5cvBYabYMrO7xWM4Nb1zCh7o6g26qM1ugx
6RLw+erT7NJQQVBJfqHqEoXFNGjA9P+phUppPZWNTUsAI1c2seGHYlZ+Whd1WbFzMkr25ym/0vc7
0AkSdEdhunM+dvOQBQO78Ke+oTz8m9SU005FATjuvHh7ZzZgSKUU9shwcFnc2c5u+tzZMZxU1CIr
jkdJf5KOg5lXk5fT0dv2i+DhR4W5U90INj7fTFljExpCjb8wXiLzr+V25ZagvCnf6wQRW9kYYF18
EEpCPPovwjQdqXZgUA1qbWQcOaZVWMevD7pzYIoGjhRXAExWnnkzqWJU/qlj8455E/ahcNbMjy1e
2F8jgCQ8F3rB1jchWOks8I5JozmpFrVY03UlQK0VQs3ImmrlYWPxaFySXWV/3vHBgn328LX/LjZ2
bA1dlx7pztALmrNCZnz3Q7ezghAp5xnkv8M6Gt1bBDp/6AQe70x8HhsCwX4FoRCbzrGzj/z6lGuV
ptgHOoWGyg64Sk32JqbqQuxY2S/qx10P8o5FAfWsX+R8IXCzMBj8arEM0QDrL1W+5MkLua7X5f9x
MqSs08Uf1oQUWHYpEJJcxL9+39/wzcG/MQoXfdPxLh7tQTpmnHYV9wUpONpnCtzecXVkb6+Fyylx
rZAFZ6FJEO2QJ9RTItsf9OPnZ1FYxSMQt7TJ7J6ozNoP1rRw1GHDYiRonH+15mAPofOchKHOys6X
aRk4et8KAAuDFYcFM5PBajDqS9LXFFLB3VotF12Qb+inyhxn+buUg6i8h/k5lacjh32lGu9j6uKG
wxdOvI2o9Zpra9Ye/Y3JDtRHymaA411W3QXmc2pKbt/Po5n8rkumxLfv36XpH6DcG+5X3QKuflGq
GO1fZO0scGntSlpMlFnq2ZMFevrewvp8kUZVv/q5XIaneflJ3oFP6QMj0+HakiZLO+8S2hMOORud
qS+DN7a1BZQiJW28KvAYPlhijcRFUrBoxXGST2kELTGGVaAD2q236dVhRgA5BMPIHTcJJ5AOJeU3
R1VvDhVs2S0qMRGhVAQzDz0577Cl4CUs/FEuZMfxRObq+UqQnZGzcw2FszT1TBojDPIxu8mwN5aa
e9ekOjhEh9Nex2ps30uGUbVXlfy7fguWC+VirXLzsH0O6agOGMu71RRkVxy3oT+lHbIM7KvaMol3
KmbHA1Qneit8sHCK/3YCx759X+Ue9ZQx2pouq3XT+hQ61c3+6d5p+spvT5I2Z93Uhd2MsHiUhOA1
JjFWQouCPArohLojG62uU8JeA0nrs+j1kHo0FELxsdik1aBW9RgsAwsF2KkaqubiFjBcOCkwQS80
hWTl0opLmdCAjdik04KQRKDB7W4IV+2Wn4Gf2oXOd/hZeQtnIRASS2Q4AHtu9YsVvECG/VdNi0Tz
SkyKjBbPHhAG91MrHQ+T3b+cTWJOAx/0JHM6JywYbTtLtVnh5wbdXRp6ExVcCfUjBdnBmbfDfFtX
gtaJt2/w8+ISzj84VDFD7GWOk1apLiwjdhXjvmm/6/L75owAp1fBTNrrGuO12+iFfpHa9U8cluLm
NZfRKj6jp5SkQ8tarQqV4+rCks6l+tbA2WkD0SbGzKHhQkV0C1rQLd6jlHD/Bs72uw5SKhaSA6jC
PWeywUC5VvmsrXI2neDBbax1zWIVg45XOKYOm4fee3VCKuWpn4DbOgeddfkVnnxwIrD2JenLyXRq
5eHRiuRxc8K/rEu50/qR+mk0r/z51VNON40UHiEk0Q5uY4ZPSvEjA+GdoQk48QaswOmV7w9NvxrL
yreUF1xYHAvUm1ZId87p5OVKe7IRxqeEfJo/dJiGDwwESKCXfnzHrD5XKDvf5OjLmqPrsLu1bAHu
J4+wb6iRFWfYXEKMC02BaFycnqfxcwqeaT5ZNqeVZKKtoLB+RPZmbKU5wWhVuHevY+58p7yYIoOy
fUpFQ+6hfirvFSvo3YB5zxOL9J6OBjNyYIDBGr9EK8k16a7WmPpJCyNTHFVwUtOvu4y1mgrVeK7Z
Wb9ZWyk0Kw0oqGL5y8fmKaCke15RKt0hoPB/rQoi67bOqSXo398HKXl2rRnAEDWRNCHjwfJHYfAf
uboTg3JT2SoXleTu8avwO+aSz6RqHh1hptqO/ltl+CH91Z4LiOg1OSp6DPvMUQmgQIqXl7v8UUgc
cZV1VC5n0Ju0WMVCwPafQeebG6J6X2zq04d8iodZSFV7DBeK0Bzkl1g2K9Wwy+U8dYhm0BDO9I6M
yoqdaPbKeJaVkdiIEX6CIXQFoUHtUW5a6O6gx5u7juen9Mgg9rDjEgHTcyleemnXXPMJjcMjAX//
kV7tdw8UFsQ7pUvgo0biSJtu37shNxfgom5WF0GCS6pEOQ0pYv81j30IQ84YfTsXtgMhBD8zSBlW
ASzmDRdc31toyUa+AvUFjauYNGrpp83bEE3BDDf5JoMCM7rcCsvW9GHtG5RsWIl9uzvJdEoRHt7w
EiHiIroNhvpL4JIuj4VtqwszNCVQXf0M5opix9Df0kZ6AElI5Si0E9BWFUxt45AD3GibiF+iV1pk
0+OI4kMaNXeg6vGrTFXYcsIf80ZaUpDNv2fe1zrdxT6ZFYMzmqR6y10pIJYWmwQo5GBQ6UFd1cx+
O3wcsO3FFmA53SHtYo6JksBEBopHYcdgqdOkBvCf3mpoIW7UL23HRXfvwGWhGjDkg0Wyo/+MWa1J
1O39UTtIe6OsVtBAASaSVFWnwtquyfKHwh4j5PfXcYPlYaQxeUaUuINKUnUJ8U8kNRTRkvuJUek9
ApvXg6uZsVMF94lQq6f6RVqeN/lP97plZF2uyol1jhG71KtHoZI1FrqVXM8QXVxZPynv5bSCHNu8
uSNE4wBjnJDX/efI3Qie8Vo9L2VzoptX/6zGKOQM5yAQLPWDewTnt8ZA0UkeMXj+cHtXd0aDeFfj
cli/UQ1wxq1q1lD/fhYf3ZMNh1hXy1mT8JTkdMDZDKcq7FQV+vZtl0dgQAEUDnIXNgXMMlKpZJXn
tIvg8ksStVu12q1T7PAzUrSPU2C+gx1j7o5NzUFKQ8WwixTJa5/FizHhhm7OmnK87MfNoE2ySC+H
S7Pgra7XrKdMCWAg6VhzaqznkbXxcVNQl+YoKXIln2jqEj7BLgmr1qynASi01JML0f/dQgrZ2LHw
kCghiEpy03TbUmhYMbGQb601jZFn2+jAEgS4j6hQ2lUXo5MPAlFF3/SKQzS8ud3vgWQSBNxvnBv4
o1W3pgjfX1hjBdxh09EBFifGGp85+QM33KCToM0isM8wJvdxnmYoLBJGCwIIkl+2juaTNl/Ndxzc
/1v5dpHEL438dO1n4NyEyQS9/AFd7QxfkS3JVoNU+FPW9jh5/TWnBClW0c4WbxncE8tnp+g6T7d3
sNTDkYWVvfT5nsbDf8o6PZgm0FoYEPSS7hzyEdRMKBbfpwq95+D0N0SIWuDDh25ECdcpzzpAuMbS
QTEYNLwF311m5oCvGGDzrwqQubYW80kCi1IkjionjG+pudnPHk83GitN5Uwfrwpq/CGjoJ7GuxYl
t+8lUfXs3Ry318oMmtatDsVdS857J/y+yHI0ui5oPIx5pet/ZjbajTr5sm/1PbYdVjXhFuSgQ8rW
uggv0kD+PdPw7WBGYQwaaE9QkfrQRUjz1YKLbrl3QXvNubnn4utro982q5O0kUvLbb2mc6l/a/Co
iHCd3STpge2WVqyCc+N4I3iSWYVDcjRWV3IKQOANFVvkUeeYaHKSd7NFmq4otILp7qZQZv0lkoZa
yfkTC7HaoiQCaO4yJaBlnRbzvvrSSSj+rWlEbEpk/eSa8lHeaxrqC1weGOrbDcY4Yzp0UFVKl4KR
hc9Ur4j4Q2VE/rBIpKuKn46yYYG4ro/7YpKfJW3g+OSlbZqQbJleO5FI2lGDfBKjKOoSszellFaA
n05kfvWeQIFl9DV+QEIAQnJdiA7LV8h9GD0p76V5TvDGipgjHfW1s7tokXefsOx1gZQbyMaqLDGF
Ufjp8JXt9rB9nbpmeRdhYED2AEiPOkyoujMKSBrGPSzqJzqLllSkzRxUEOi4SZpVYwxowjEM3mRQ
Wa6jdnHi1PIXF6g4fap6UuNupj7hLxPWlzKYLqZBbL9CorcSiQ7ss9Z9XJ0UAbGRlmTOFj/8yxYY
tY3Ct09IS71xnY1/VqTzlL84olMIRB0aX21n1q8NBS3w4AffwPI0Xijd4PA+E/Yjac5EpRMG93g4
LDjpNq+eEji4a6Pykh1py1RenrVyrWIKnudFT2zG3BpoXKMzHffHY3nuX3CjI8pkMWOrlgJZl1C1
PnagxvRnefahpYUqgkkqqePSwQdpfC2+FtP6FmtQxt4okh8CZz5lXq6EBQV23hhODWDY58Qow/VX
cKTzXR2o6p2w/4E3YhKgl5aDyJLOYK0GuBa8gSgQBj3jnqwQTmuxBJedF/DAtfFqrssa7Xol1LB2
L/RE+7YDULA/xbP/Ff9RPHH9rsfny5eTdHVXhhSuPhhtWBiGQfd4jtQiMexweMB/7pPN7TKJPZnn
ZFPzRxBue2ZGopi7AxEs/+8xnbCpr2eu6sU4UXpX/RvP3KxThLSPWrSfsGkGaQXBrgyeGKMQk7E0
owp+dMX7cD1ZSNBCnXQB9ulcl3IOqkTsZG4IoF4V8bxfOrnC7EsAfrQ6Dvr2ZrhYrp4MOTyPJWBT
Y/38B+Ff+N6UEj3Kf6WRs4Z8VOeDj+rzNILihiZxLHfHt6JvSqJI0NKl3/6b4xQDe5Fcmcg1gHQn
1PTI/pjdzZnaazEx730JuVTvHD10BfMJaeiHToTJkpY8i81OUu7NQBTq3uyDHSogSl5hBu7r+bwj
q9BUi9xZmlp2K4b2YjyUQBtNGzT5lT7Xk9Uc5XRaD0E0Rj8gwwMjXHqrus4NHL4iisZ5kDeaxrzi
eamo/iVU9X4Q5b5XjBwzUBM9tW0a6bEyDWzGyETWUSkygRZnB3Qo5hz90Z8ClGf1qwoNlGHix7xc
yOGlPLs98UfXe4oZpslz/Bm/MVapmBsJ5BX+4ks/qtEszTtlrewvxwr1AIRHrLlkxJ5GPnkvriA3
R092+mgQiaf7xvQqHsveucsxsSp2yuuOz8RldOO/f/J/PqXLMIjdaNjY87o/iaJFz5Tp0cf+O48J
+AGUpnwBJz+ju94UqhScrAApV84oyEvy5H4gwoM0Njn1Ls3mnLhE98l5FthwtalMaaGko5AJ1adO
Z4tGy7OycctZfGK0xKvsKzQeW1+b0mi4RTscN4KD4hYQ/v8oEGigdgsSyn3Ja/4wGTaGd2XY3jcH
KJ6EvH31tfGAWSTg5hNzFwkSADhGE1wG6nPT1q7S92SNOHYgfMZHc9RSbhOsFcDWGFEPh1NFcF/2
5e1ozXlUn4nt7sGXQ5VE143a/Hu+sgkrsKNYhvzDfakBTkIM90tet1xhZXKLiVrP8f9Gp2eA6Pta
RUJ73y7U8WfmnqZLeySQxxzZwKzeL/gPD9kxVSWwf7UOOhhU8hQNnksvJhVr63eAI7bFpihBVHz5
nuhq5qFLrsLNV3M7BBtFTlDdp4LKd8biWCqHZKx2W8WhlkvvRGEyHFzhU8USpxQ7MckvrMcy4b0o
sjU57oo2OgfBg9zf05vPotB9o07DN5UKZzkr8RMj9R234QZ6+3TLDBp1LXk1ivFWD+CSesE4j50F
qRoDt3TsKmFWp2A7W4LDFzRScoZL7yaMbQsnR7TidVEvIIplOq+Sc3SyQSYG+6phuzZxbn1efLuH
F+cG6P4fkXmUTX4VpSqJWg+MgFRkHqnwv1cA48J/Wika7TNIuz79CeW/2OV+/avQX1g4rEDGk/Dj
I2s98ghAXTHezf7YKzkY6oDN8ZglN1VL/tJo6qiQEym40XmDcQKLHZpWdAEbbKp29QSOlbogM25N
r28f38hmO+ecw3QweYmRQtd81Oo9bzTDWgIdNNElx2WD1ewqv3r5npE78peHQtuYuI+aocx0zsjf
BieGX0W10T+JfpSxcXxtdG5hR3afYFSfJLf3yoLyU2zwtZ4E8yyK2CRtG0M0FH2+o0Oh4L2kkaN/
AArS7KH0J4B4ZHnzeyOPIsgI/9nsic+R1gwfgnESP6enggOE/VeWKZ+Wn9AEHQolvxif+mJPzzck
96g5xz6GaDPokcNgdW7c2HjE63WHkEsKAdAlaHEVacu0N+zn99+CXV+9DYHEUkyFrXMwdfIepXmk
98i5AObyMjNSH3o9LexyqHJOuXcIh+yBB/NjA0ZGiW2x39ZOe6VBwQEryqBZkQFeK9lI5+KJMuvI
IddBLho0WmyUTUbgatp6R2QSTjNvEYZjIwzDC1jWKDYz9oQRUwXfwdhkT7JwkDcoqF0chv4qoNXt
k7f1ReAdg713enCru0ZjxnU8Gw8KhqU8ZiOIenPqJNVUS/VBx+NfrNSh7R1YSB/HLgOfPumpvnhR
T01v2LmujNOG2jBACduBZYbIax79LmNY5vqMn5sXo4uE2eEg9i/oF35J8ExHZx9I2DkzwfcE1jei
3XTvPN5IwgbEbrmVCd523fBR0eP+c7sBGIWH5O9KyaaNDwcgpy8vF3esOrPKfMQ4Twug2Md/4X0l
0KUbE56FPFT1Ue00PsMOgfE5itxk2BMy4+65KOCc8Jo/Y7/ANNIEPP2EsGxTLKsvXLq5EXfNKFMs
ywqztFKOTDA9cIPWpc/1qjoSoalvYjCUmHPhufgMxfA8p4BDsW8b0PwLIxAKiDlyTeGeoVS8ApO0
4Nzi1D9SFkTsqqolk22nZfUaoCuHbVc3S8Ol1r4rI1VrA/e+pWmhJyjeAbi0FiUtax6DmbHNDGvn
fTi2biBuRzeONMtx+TqUlBQjGHrTnz95tIrSxW63SZFuMf2TsnAPduPMxuutNElw0wvWyURGfcJk
nNaaKkMSjTOQVNxAmQMfust5Zup3PdUuCCsSqUwdXJ2xSbJoS0QTppL/PKTQWbySyw3R3WXvQG6y
9p+zPLwjdBSouQStA0vv5woNkmjYwJi0WFyHtO+c/OeLv64HOOpC/QoifwFsFNJNb8QqD0u2Q3/W
yrw6Q+Uer09mm/wbRvGfmeLCEgj0pp1GFF7eDXFQ25X8xlaPZl2126CH/6bFLn1FEZa5c3K1shi8
oOilGmu/7jnBP4mf3ACkJgGAqW6gYBPdycmn1Wuj0UMJ/UoFNBlTqUzclRdjDT88AYxTjzjJoIFg
2KSm8qm0j3E+J0ci8zZ0xVD5Z4IfyzpBfNi7na+mTeCRF/TsfqZ+2XtX4DL/FQOpSQHSOe1tZwX6
zBGq0FeZjtr/rg3cW2NqTCbGdOknJROs2BxVkslG8UkG+3rc7cPx4ZB7hq9ocAk5bfXj9us6UB8m
9MDzFaks2vdlrzTgAo6lIRf4QzQZRMpOOOiJo6eAn0VCCurH4PCjFD8MnNkFU8BhB9whBfVZxV04
WG9LK3VPJLH474qgp21jAV1w273/xOTGEHOyNGov3xH4sBcrmvycqDqx8xBaH1ltJexm7IzN2XBh
pIzD5aqcuvBL7R7SKjfXyyeQtCeIdfOmqByYYyb1S0AlLNEjMck1oGdSTpLQOIVPP5FNIBq4tgLS
Yp6vFWBm09tw6x9SJuR4op1nVD3FDoStEdL5m7YVd8Ts3EdPaaW4ROmTQufW7kQU1gCsMCCt2mod
lJo20sndUkskXcJcomz5xOgVvSU2rAgg1cVsBaERq3ref+rYY6hofqEvoDCnXrNx0IQ2HJXD1yKA
EHPzTFWw3/v51GklXxjt3UV4tF4oiHGqczQjnlGzgt87hezqPmZVRH2OB5KhpyB5i/SO53iW6yCy
clKDUmm7QiDRw8YNZt5BDNhT4uoF7H1XMRk9TMkBIwXyo1iuz+qiVl6Hz6ys0ZTEM/bCkC6n4M5t
m2JkJMh86wtp2W2+0DeMrimafmUj0Eeg0LNismIxzyr9WVL71BWCVtrw6W7hN3mqc8DeiXY4bUij
NBjspeyldCOLSmjFp0Lx/+egK3lb5T4EisqNZMbG/Nlwy5zWc1ttGZBHvPLcDxdN8xSwawDgEGGk
4N6lsLppDb/d5XST4TbaCGvuq+PZClRJHOdYnw9luB5OyqE0ttEVimpvZGf77ER5QTu2Ui6vXEB9
P/wz8xtEVkEKqRKwTqjbhJ00shga2c+av6IbsIvEaAdi4n61JICJb5hZszGoM6jRFaMAQRflvtK7
3gSanxnqm5aUrc/ZUlPc6M+ztTogSZcGEBIG8k8ZloR1p8rphudfI/6hddSHLWmIQbWYJD0uePuH
UfvvNiEklR7+vRJyvIV3cACLmdI6DO1gYji73vvPS4iNj6Ydstnvrto+AauxsPsDSOBleNpnHl0e
BZomeb2m+RUTW+t1yOW2j0Kv/tZ/vlrHy0tW45Os3eJyx48x9g61s/mKbvFrrylFjau9aVj9DeB9
Bnjpd2SD6EshdIRiK1DYVEba8tnX31+z3cOqGQKDqq3DNKNY6hCKQUSqqfT8wdvyVFQ8ka9H9MqG
paalyDE8coapnDq8atex8MOxLDJYZociZOANiEz1kF7SmE2+B8VRkrLk9y4ymR2L4rz6HPiaeKJW
C7iQPxoWMObTT+llmfy27MTc9X3LjqA4NUp0OpqggN2XrkpMuZD+0XURjEjtYj+4wkJfSLDs8eq8
/lOhAL8HQY+Kth6B8Uumm0Y9lDlAZugXtFiWAsqOFApWeZN25NJ53zTKI/T+E2+1/bd4s/D8focA
we7evpHovQTplKiF/LgrGXtL1NlV7Ikz63SZlDNJL6K2caFAHPRuxXKo8BSE5LGjfC3ds2R+ctam
WYS9ZT7e93AOZQk0i2Dh/0BBm98P5ocBUuaYGiceTfYG/3EGHWP4RTfiQ0w8DU7Nj8GlSNRJQ6yJ
DztNAJ5Io0Nzn76qAXGlJkCb3225gF6z+Mk5Pfi4dXKKHQo8zN8Q5Ar+rmsnX1/IzNyHRwjlCSFy
Hm2HlGuC0luFWx6wKQRMcR8fNqt9bLcea/xnW2XLNK220bE9HnTKrxlZQIDzdpUwjTBYG7h8OQp7
lTm23y21BndSPnZss4//iD7IFI7D/fMeN0OFo7kT1HAWsvUyGSfgZ16jH3ql0CKPUPpJPbpZdQ81
7SKQi6WeHkao4YfUSIq3wPf7OCZjj0M4lnXeVBDzCerT1G2j7j1fnePbsNdy2syFhGRvE9up8LLa
c6hR5UEjPmV5Vd6g9k8fs8k/vdC0GokGjj1e5u8hqgjKmQ10fcFQiDif6Kn3JprrCGtpxiiHw6ah
pa1oqReId7xA9LrtdJLyApktN9ADAsUH6EJwxHyISogQZ/xpXw8EXalmCebWQDXoeg3XJLMXPgjG
HhNdMVrmXTvsa2cFqZKCKjxxAE2/iCy7zW0XoRzGWWGpq7o5HWT85neHPNbp2RhM+vs454aiQeJZ
7abPfxtCSovisXCUonBo5peQBxY2RO9JQRPthTSAD8VSqCxVPAeTt/E6U9Q42q7FdIa8iu5PEz0z
CwcnAGsrrKosDfUTfIer8F3H7RxDkjF2DuWHCozXxPLD4EwECAwHrhmaSsmN/kK7a9c6i9Lbn4U+
TPANuYRedssBpCplE1cqOehymRjlQ6rHAc01mWydKtCZATWyMNuzur14fQPQkAxBkmST6jAqcS+J
mazVmhGLF4/5exD8e9p2u0Kgm4HIILEui6WhsQSR6CfbYgCVTDSFSr1hcASx48Ad4T3RMIZGZmbe
t+Kxlp86MmmEER8xHIbThPD6u4Fh/KOpQBrJkxNpzqwBaN0SDs29KAGZYBeUnUKGsaHY740Egnpq
onWF64jT+7KKBlCDyIOFFrKPHzottobeqrN1DO5tQ5hmNIZlSEc37QUQgZSJ1bGEx1E/wttJXdGe
dAd0WiCAvQNTfXQjvrZOsZ9GP5p8ful4mmYQEV9IozXAyisfMHTtnEa+0rSEKhMiZeleo3wWxEI3
1BsQQXnuNKUhTZ2c+0lTHF9GVJmsbv0AZJ+3MvDO6xnNMEJsXX6Ufa2lb7X29H14TF5mfBMJnthM
z/N2kMPHKLgtHgUwz5sqz0KZfQYX4ip0imvZ9ybzACwEP9VzfC2WZ8sjriDR90qWN2Y8d7odtWRK
FZUvrZ0mOSqnMBzjcN2M6yTFhVxGRuCMBxkm03EIg1pXvTSAaOA5jGYwT1cogj9sU7vzhwyMPBdL
03+b79Ponq/Tf/CeOHQcosc8anVdxb0hXfhFHLrXZ4BRDnJriExEgQIxO176mwgUtltE7zhOKz6i
Ttspgnk8YyVCHgYvlaclOI6HoW49swpnFpwnB/3gNLSKEJYd9W1dhM80USngSUNNHlu9UPyd1S2c
MggAC8+4qoM7QSlgpFiClu/TmQc/EvjfJHGLdLHBTAAeTsBwQXa8M1TSd4u1rtzKIDWS5ZnfGD40
F0aXlifJ01NJrOS3OP9ZqR7LhXeXmkUMNV/rpKFZwodF3tTnLPqufR1vtZd/SxGAOTJtHMrezInY
ZIEUeSHRLvbQuzpqq3ldQ8OiWah3ocwkksaEF5Ro0YS5LzCERVlYwCs+2rsqJICOCBF8Jf1BwjII
KKHkFy3rsb9EwCproxNhprvql9KvakzXdkCAz5nJLXiompyC5Y+8fOyvv7xMUAGh/4JBxoshcq20
LWyM336QHrWIqIa8eXQ8CAKVe8uqRfLwV2yKMAu1Y4JXhuLZ/383XeySoOytIaeYNvv/V56vw2fI
uMEfHEV0GD6TyoEsR7S1JNHVe1NzzRrd2WBbwJmw97v1ybIGbmdCevlOuFD5CeNMBn7N7Pq3tn8V
BqJr9e1O16inXZnHbgGlUgLkBdTO1w/Dn0OYUI41dZVrPX7tdn7JRRaJ8mXuOvyJDPuIa+VIBrpT
os/BiEWnvG9wMMgujnzavoZ18jCUxzkFsN7yKgQOE7v7zqD52oV3J7k58Mn8EYtJD5U+Gn5o4LTq
sQmTP9b6+j8ZBBHZcZbaiFNbXZ7JeRIHGOKdpLwsql6oqj7f8SlmXHxTS6ssgUez5XqQxIDwgQMZ
RLDN/ucJ5sqmj97L1MAj4KZtY4Y/Cms/yuq8ywHCDNrOrPBfn69EbeXcSk4hlb9crd6N8XE0Go2O
v6QaWhF48wEK48kwPIHw/VKsb0tDlH/zjeujyU7BpcXSBjo7sSOz3NcAcNJ4IMX69L+McoTVF8oh
VzI5WnuW56Nf1enWym0toZzhT2+Z3utjHFawpFaeFYiDoBsYcQDx5dw/mtruDZG3UhOfBxyp27V8
P9s1pSvZhB/T1LlKqpY77LZyHFN/fCjLP3dXxibk09epT5fdIS3O3RJsAP5LGcfnRlC6RZayN0h+
kMCKm20Dtmp7hgOXRZhT8Qq88vDrSkXi+EmXFwxVITDSqK1/vwbs4taOOITyNnpb+W9nv1sIpyav
s07JefovoZiz81Iy2ou0/W6ftUEUu/Bw1kEvUTU2elAdYF0VsBGGRY8OzNFvBSaxKqX+6Q1gs3wP
ieGr/B9clcVqjQX+2uGEvQwBcMmjLVDdJx63KiUotEVbatwTZytquGGs5FotTp6rJTECP+cgsnEZ
Li1becxwUQc2shxFDIBXKTNQEnE9JBFbsgZ1hk6SMEfbuCAXgx2P5+ouB9lZyI4GxhfUI/5hRZkd
ZeKFakFaBvjFvam/Q9Ch2tFURop9atbVf6YZeaBu3oZA1UVctrXc11rnaY6VI/SAL3m8jUR+GhxW
EMDqV0weSoCOsxMwbsKIDvM6Q7bcc8OsZPFdgilrYFpz/hxXzjgQKdFVPzgRR0TxUhKh1B0C353L
QdJVz0XiFwDryceqlO0Hom+Opt9Z+815JitmWKSQinoTqgXiXGtl0Y/Eyq+hdS8SjUYoHO+lSmjL
n/FvM7AJmVheTHOOdmg/Hh/WslmhrhdwwdbjlFDpsvxxnvovV0a9f8j4DpvRWNlkqpD1a3gpvQ63
RfQL6mo4opVhRN5bUPKmjuIFM276EHf3jTR9dMzjReyZLnCaeSjqXUeDTOCb507ynjLMcW0FCJM2
Y2tlqdbTBBWcm1KG98KxAqSBG5Q2brafPs0V6IGyH/FdEX9JUlZlFQC+EIIKM39xg7Xb9YBwy9Zh
4/criCU/+rZru4sOwpINHyN5Lb2HuiKCc3vBKUzDs+YYKnRH0oji/TllWY5tTlGosFkcOiMKC/+n
gSuWEh2h6OKsLyGhaGmDWnVmkqakyNCByXnmBIaPykxjMSbPqRb6nFnWJnv/lDNGxPwygmRV+W1x
49zwR+0mdZCf1KOd6MalQqfNpD8nkVbDgh/H/srm2CeylU4kBUbDph2vr9/wMC+VvCakWuTJTqGG
sCSDkUwa6VyBWS5vzVPRSq75gkPEvMxv0OzkKD81YF8WSB6JaWDGO/wOLWK9Ub29T+Cd4y69Ai3V
nmSq0qd8gGhUbAASX4lWjnpy90fSCChHpH6GuOxCNXuVXQKKcONsZR8+s18ufiOkUUD3x4Zc02dr
H0RbkzsVZtlIB4rhapbKp8ZijwCe++gqtUN/wyBTXT3jRZr3vj20mIIN0+a5Moti0JDoae+FN1N4
Z424m3GWqvRFWovIZW17Wd/9Sb3Z7JK3DmA0iZ61IeqZ77YLYXNWMXIIlDm01aL966Odr8L2kiAD
vHl8wSDaio/tDACdaSI6oDkBqZjWilvIiL5MzHm2s7/n24NUztJ1zDUoNFUuwu+ZW0k8BzMaThYh
nL8sKqpcIStW8UcKT38pJMUy2TO/ZSboteAZoNxT9HL6kxIMMuPunvXrCPfs5UqL9fPtjJmQza+b
CX66oiLhN/qmp5AGtPR2vNNse3URSA7w2eA/7ovLMilT8HkQULIX9DirGU7aq+Pgp/TNDsUUunap
1yLCLZq2/ugLxON1SO+RTrmj2NChgYM+cS98c22M8VowekVuCV4nghzAbj+acLrdE6BRlEYdogTN
CDSmdZidgmIjaW7wxrjd5NIddBG4mrf9Fa9mHiRLLqVKYpJDSwRBz0KdrP4mFMNlUfTuEaSY53Xg
SVowk2BHBuy0ERGcf/uY1RAKdRwrqUSZFctSW67+W6Tt4L30gd1+Z13Jlul0r5XFRrdQIeEjCHem
H2+tKZ8GaLzT1JQZ3UU5H4tPZM7HcS6XyxqfXgXgreFGSigXOIelxhcJSeOp0vbsrN1/TapehLcQ
jMAC5OM4/TVjsTkyJfR3fZPt+FusGNTcw1uW3xtY0ezN8/97GNbkSsNs+FrKw4TDFSvkDEWMFWaN
64+pM78w1u+w18kL5RDyeeIjslljDU9Ihz0DfjH7y13USDHqMX9ENgrFBAcRxaGchI8uauSbug2K
WVWA9Z+td9GF2KJAjFodfVGUgh5KP7iuugP4tfuHIA3vL/b+DjVKLhXiiWlwLzfUmwOU4jCCHFvh
E0ofQZojGPdflH01iNCcIao1etGOuJK7cPGOMJfekQjrXK9O/MwKK+zjZPkadnXTGRzslqFXQYNS
gIW+dGjbuPu4mFjGARm7y9AT01wfwlMgchChcQmFn0Xy8yt9iAr8Aq2df4OPK7C1MXJNPkjOrbZp
VfsfJ9JPcM1AAZgZHBR7KjM6f/Cm8Auz9DLXUS7zGQgr/+y7gEUvHaTh2UxIL/vg+csYzylByozY
ijVOowGDv5+GvlF2mNdytNsJwowPM0l/mPqDtnh7zNflMfN3aLY8NC+Bgo7+2l2WOUqp4t4AC+mG
b66CIhcsC6X7tip8kZsc6xsCYY3Mffz5WRG5KXk50UJlIPFGU4/h60ZS0k0aIEUftcRCdEjb2Pu1
4VZJ5KB6HWz8KmrTOy5JIo2CrDw7GxjCPtwmzp1g4D8gQpOauvf1oCXv8bGYFq7u0nHQLeKkHIri
YEEP+GTM4qH+Mil8OlhQgNT9virENcOdQKu2tnWkFitBlN3DU7DhzqAOeHhcJpYh76U5O7HWDUgH
7v7Y+CLrvhYE97z90SqIGVjYJXkrTwKu+0XPxGE07imcvK0wFMb9aPmy5eyfWfB9zJa30orhfM24
T9ANTkwIu+zi2i5IfMhOXdhRkWEdP5HvzqTAhqPdaph9Z5rL/kAlbyzPntTU7kJadbHoEjyjahL9
u1IU3jwgQd/AgN62XKiA/79rKXA1YicZ+kIgBxF87510FDfdri2v/8PcZg6gMwn/vZXWSob8ykgp
GSH/FPJNN3+nueMtSpCM6yD/m0godO2Fsjz6WmxEgtjdENoew8HLQ5af96/1XHXtQSqpu88vFzyX
XReV6w1TCOyrRGWFUHztEFWlk1n2im6D8xrHV2tUfxjO3t/hlI/kJNTiSEJxSJp9nNd67O4+0C5L
x3v6uUPscmkCvycdqqEKxbgZbd4qcGgGehHCz2z9u9RCZpnBWp6BAsF8ImTKIecc4g+4gx8P6OT+
GfZOdzMkm3FlvHGxszQEaQYqLYloPzO0zBSlxg20PqAAiLgDljDIY+3BcXzCNxyxZJxPKq0mzmBy
BpSaqDeRuCgtLB9j9xmpD6xg+eRT0VVMHKGHmFiUjZc0Ivwo1LE9KW6VE66pivmEDkhZYuONSoRE
kq2z7nSKhfQU9fxBH1CQrsh0yj5xHAR7Vn3t9sj3KcpO3vg5Rg/h0YlsQZUX9JLCv5VdxZN1LuV/
NorlKA63AFJ0rhBnPfyzR2oINTpLgjRIHYg7WqxG0QG3kGzcuKzpkBFC1Yjx0zTZbq5MAc8oD6zS
jS82b4vtRWIp90EZg9iqD3XcGWjnxPbqS1dGCiDMhT+WwXXRu/EASDgfa+iu+vCephPBLURSjdpd
krzcaMnsgOs5vX3eaziA1gq2YMAMZikXcKcaPtjLHr2ekc/ak1904pbqmH4iW9HH46xjT4Ni3gCz
lPQxmWgo9KBQ/3QsKbWBYkKwOR6vip5oqrrDa7D8YSwNUMcHSY2/wsg0sjmmAlOOiB57o/8VvgD4
LqRi3SzTbyrWsNWEpQhj9SVFJVCHVuBcF3Ufl2ITNa7MjYEZhFRVMfCxsL2g3xZo+7wiT5eUUGQw
pfwvms++X1wxajy2OnN15j4YHjXIt/NNDsFEDWwqvNnRlWpbM5NvI6tr7zGTLVPzUPSjVjfyvtLv
mZbHW2AMJNSULXrEqibMgNRJyhH/VejFF85naUXgJeAvRg3IYeFEwTY2fUx3Ss3nsNHdWqtgZMHz
ZeDhTsSg1oRcAq6zCVqM3ozoGZaAY30obTt8IplMIyytFgUS9KRyXV7UxWpW5qTAvS7/K+9Z3AwT
zGGNq/0vv/jsRRJuI9pOg1g/C94+eyGnvOeY444CVGPiX3C5CYWm/atCpK+Sr2bt5DgE5TbQ46FN
bUQtWP99p7jAb7XakTx742ZlLMO6lxpuobaH8cyZMNfIWb7wWalTeWe5hb5r5meE4onVNBqx5BK2
YzIpmoQdmzgymu7WxGjfvrnaD+271tjKHW58UoL4/pfv3ilwdxg2ijlcssIC1GlJKGZ0jrVbGuJ3
KAqdnHc1lZWkfN5AJO3gteG79DyT9Mild7Wus5+5rQtBcFDiLZHrHoIzbFA10CKemRC8OPrFoIql
5uSiU1Lm94aP2X2fowEMt1pYWPa8d2M21P019Ps/CJ6wr6FFAY1G1Gqv0FEqD59wsHrQzltungBX
VL8WmpPz2dOIbKAZ3HkO4mgoyHDoEO2O0d8ur/tnEciYU0N80W2iV4yKk6EFc1riJUe7rotBUzM6
ey9yW2nfxYvGcu288szNzsFHFZ5VTUYR+k1knDoLQQjxGVgKcOKMPFxIjK4NKfUKsQKtxDEuQtD0
Svq+g1JNP9amEjoLGutULaDuZVBxBA74YzW2p7P7Sabl7dev5AomYO7X2/ekpyqcJdiIc9E4Qfyx
sSdrjrxApmtZf0MnxVp99v6okuejQf6SZlGIaoQHZKrCkNeIAJxyhpBzHEtBm3AgfV7qhQ7LCRxD
vQ4IvclaLt7IblZ/3qBl6yfD+8QKEQNVblEGBHODlgqd43cHf30oChaLCpIqy4JBS31nchKXnPD5
jxRCURkn+6Pd6EW3rxaELilE66h3ooHjtE739/QqSWiyNobeYSjzRDZa+mpiDvEgvNEsp3aBeOBf
JxnUvOaCNbSn/mZtInFewdtiEBnhjdky1Kx56vq6+sarHdI9v7UTNTioTV45pDsf249jmvHfZ/u8
Z2KrDf43UQjp19nIJsv9Dq7YKNrrkg8uaToOCKxeLohcR5cxkDj/ozDDSJ9Z2kvz3wzosJ3f+Ii9
XiSw8wLcNvehIC1ggYl4tA/UeuChZckscj8Xrf4/lD86n10o3o9wA171IDyC2t/8jkaSJa/aFtCj
EneMGFcoiz5saoCLgbFaQYDE+rE8DKUEXIoeaIf7F4cTB042rTnE1hr0I/b0cc8sg/pviUOQdlNh
ZLKF8g733EOiMTxcB0XkmJOA2lH4BFXcSvm3DLjmU7tw7aUC0u5VTC4IOR+CtewnXU0JzqK8821u
oXejqVn1CU10vHZeOW9NR7/Kyp3jfLyu1wJSFy0QvCp3jYkL8u91etwMaNA+MxmbvQkd+3+kurkS
Z5qhG2FS9MzjJ9HPSR7ebkb0o6BT4kWfZ8sURU6nAjNuqUzfnVmJ/mwpW4dSDan/zYrgSIw/Gz1x
dkRSYyTAlsA98pXTyT5JObo3YNGLgUcm9HbXRNBFx86tRYZ1O/HY0Ab0qwKZ/ZdpfQAxoAQGtkkx
+csc5vh2SKlkA4QEbsdkVLA8PmVraNTcpLnBBaoEtmFPD41I5VWi85mi6notpj8APEkZN00ojtK6
xNFeXh3mZKvtsGimn0Sg7GvRhlYEfxVoHNycCMMkIzbxHnu+sPdRHcwWyYALr0+vLqlPvM9U3awy
wWrjSJF2ED9q8lqWQmiUmpfbSMSFuS1OoPcAofC4S5Dkp0a4mr2zVn0iuBRYU3VjDr6Ed5awbUmL
HfH8fkz5TKCnE/rrNM2RvqHvxgIKxW3d7Yq9ydGxQ2qb7EX0o4buMFxSTCJXKzqJBBnRd7zBVhTJ
gq7F+XpZdq97pxWs6YlurGbTrPw5PVUPmMPsFUuVSTvhgcWkV8idvT1jz25Id7oq13mPkDes+9h3
cFQDAnTYNZhM7gJL4aJpJW/r9Xxdfw7+yYBXbn7CypxY5ZR1A6kbyVXQZClp7yUd/DY2JkVgYkjz
WDUt7NLQHb1V2kU+nlekP9APQ/IiuadU3bE6XFQHIYBpcn2oSEt2XZaIlEA2uSZSw6N/vZT3NW/n
nbdAzham0+z3Hmh7Rf+kZ4eSNxwS8KNMYo2usMCu8bONlG5ItL2CnrBnH/BcCenMwxK5kIFPYzuS
DzrWQGIr70fruo7C0RQFrs1JA2S8D0F4S1NhxsGnxbQDh4lkSg/y5CS3lrgsEARkOmiHSAr9v9HK
JVtD/5f69Ux6KwwoQJrKdBycVwomELWVWQNjAZ6eR0j05xyntCStNJHvqzVMUjzFbugzsj0YYYrC
JlPwjH+okyUEh/ipByQmjAmTVt/s32dad+rj+Mo8vDim8ah+CC1gEghmMETdCxywdR6xHBpPG1BY
dVihNF0XpdqoUSfLbe0oMcGUjp/RWh98VY9/A0QxphLsWo4j45Tr0i+zWmOupCBFhQk5pEKd0mHt
e6CxSG/VOJsLMHnGWr1RAbW7k2+EhL0Mup8CBTWwwjLiFY0HcyktFTrDrt6/O/twS3cx+OquJzAN
iVgUdc18HHhS00M5T3S1ML6TfnTml5NNVHWD006FlAAW1yPmr3vdVWSuT23oZRvzlTKEf+FLeve0
8oA5qEbsLs+zsdWvGgxMdkjxd+PU9U1DfCtAsLDpowJtAtq9OzRCNsPXAdyfHiVt9ToS0kSJJ1jU
3MqwPFBYDeE/mnPm3W18hCGhdX6T5JidazVo/zN2Snd3VFhVAKhR7R6EAjMSS/y3NtyjGEIU1h8M
DkIfclrkgPCS479WpFyjwLT7iuuG00Sbu9iSydKMDXydLGziX6kXZZBj2KzK8poIMTIhHr1T+gXc
C19wMeX9hgkv5Xrts1wg8p7Y5OOfrrVkRZNd1kQReGre4eEWnSdy7HMCI3cA6aoyk6fsqWzBGZA7
csDslBm6oxIB6GKga03v7kFB8QJyi7APhc2Q10MaLUXGWU0j9n9k3UdjOGVM7wS893SWiGGgCA7l
MrJVivMxfoJhoFRROXU7Ck/sijIBL7VVN+VSYthwYXtyEiVhIP7Sb+98HdwLwf+VmMuSvWkvB+bi
6aVvJheX9unj3DgWnJ015X6BTHE16kSEVCN1SbZu4X2BHfC9SDjcwKDTwng0N+lKH/MXj99HNWGT
1RFDoFLMIaUPNmesUOA0QDlxeOa51+DSZgednTmuqLY/u0JGfa4VyNAj3IKE5iGXinP4rhsCUqc9
XZZTcYVeY9GKFM7bFpSPcR719ZgRrDEUqm8wxGLRa2AzvxoVRAk0oWQOyUsj+O/1jlm2BX9Julbz
7eBmTyOdZXZnnfjWgVzMPZvtjyQLEOQ7gtn7HKDbZNeM2yaXKJ6cyUukSOPjA2sUjQrTdsgw58KD
dzr2K4pvIk4jCwwKPKUXvr29BJ7mfZAKTD0g5JHetXr8R7QhAFuFn7xnWS+pR9KO14mOopjCNHzH
ZplQwq3tcYrvplfxW1lH+g09Vn8JFaPGTiLL2Xp/l4fS13A4PhJz1/CL869UQqIoVAaHbhDWKNOJ
UlKJZE+tjP41BUveFSvuIH6SvxrwLs3GrJxpvVTqV+HxkVCfx8HxaGho0x04qJmpJ8AlxWu8DiYH
PXwNVLVileKosVgU10JQF6fHUfVJCN1If0/8jPy6a2PGPZsNBlFTYntxaVwN64aXiGZaxCnKVBAC
jHwL46hcX9b8gLWFTHBlALPcsj509vgq9/H4wGaDG7o48b5kVfqyIoUSXxFb42JU05ui43o0AqZ6
O+/9zMmj/Hib8gVaMraXB7dBWyOT2q9Zyh496gi3HPC6wbqfd71dbudg2DWy2N3I0m5+4PdHTcAB
ybT4WGluWhUvvlPgntLmsOhnCD/7J3AN2RZUOxsGUHKrj1bcMhErPAyUQUubytBLGvJLw8RMUFFB
1jYVzfZ7YDUYumKmidQZhcOgPTnuX4dcAxYMxa+i7oOCZGqNAezN8TnTDPNMS0DthVEnO1XUYWvD
vL89LHWq7rfNK5sqGcVVSllql8lgm45zEDmv1KwgHT1SAAFo39QzYn/gFhb2BWgvb91TouuSvFQA
yol9Bt0t3kJL0uS7kMuusfBDvsncEeZBWLWlW8b3hisGvL3DSjUd3rYCJmIcCH5TRmS7wG7dJl0L
JJINPb/bxEXlNZ21Q3R0XUO0B2RHeDQe3IHEbHWnBgGZPX24R7VpTZ1/IA38TmyeQRoAu69+u5+V
5JvRQPWbkR1tgNu1rwb7l0cYZY/mRPGsYJDnG3jXL0RJfyw4vWX+WzwKksHq+cYrJ5H5r4sprpdf
hf1p1LxKzOErzfUGY3Km3gWsDfF0YI4UbsOLeQVBrmH9U65UNgd9nLy1ifKXYiiG7+qP764zBNGG
tdPtbNdI3dBTxItzCGGXlpa5e1UGDLhmXmAP8A7vhsGoekjM5kq9xOHIhhvDOVWPnYmAaOefldQQ
7oMkQioYp8cWf+/X1Mk73aoqlShNeUq6QV8MbLMtZDKJ+VglmRLevZ1+k8zh8jLSD186qSBzVYjC
gf81hX/fqwmIdqgxHWbXnrlChwuvC3GkHqSqzd984DOHNWqLF3yVOA4bXxGYBG/wwB7q6Yyp70Xc
nbtX0d/n1KDlJK1WEQoKuEWv7H4sKuTxMDFhzmrJhB+qPbpiXs/Gaxl8SQcA6+TLxi0Qjd4au+H0
ygfkKI27QMxZrkhebTMIgYU/PkSQe6LgB1lO+CmxxGLykhM2wmTZw2QUoTaweELqGsNCXBTYthDX
pmOZRQfpSls7NNWBgdEWn/13DnUAUKEq+qS5rdsIuWKtkPASWDV3LBYuxk/J34zHuDClSgHEkWHG
+tHbe+WhWHkylDtksLPjTxKp6ehwAhdm0tWGQFp1HXUtpVU8g3c0T1Zu5ImEgFBA+YbiphglQqq+
VEVh9uvZG0KPL157MALCRsZLNB/9EMMhGdM5a9/d4IaB1jxzkwds1e25qX2DFub5LBC1bi+psF8r
LWJM35XIhg5wJdO0jPaqIj9yiYnNXzq2jED7qVHvScINWSClyP7Q27f01Siz06eSCno63ka6OQFj
FjG9PMstXK3/DLj0mH0COljIIfNpqut2gt5ngdoWs577vuU3HvqD0tmdZ9R297u/nMRz45bPTDdH
dwf6AQ6CrLrv66JDoTGZ889KuSyb55oxaNVxHAQBNm7JjzxKbQdZyMt+hkBzeIpIcFa0iQhH4FUp
khccKJHZHsljfKwBs3Y2FqyacR47wUDHl6VGyiP6mJDdoA/TgQ+AU6cLMkBywA8bqgp3QR2esiXl
dO9Hz3P0MGzhPcErZDtO3k4fRln/h0ckwF8kwbHNGZ7xt2fQwuDrB6fSg3OJ7ILvvvUfFvxIvHms
chLdrX+CgLoEpnKgL7nFhpegsCp4IVjTZlWmzpAep6OIPBICKNXz6mhZdtU0O4ILGfEDr3KN2nPr
5Zh220CLTtNSAn6GXAElE+8hDuQ6PbHtNRvoB41D+elCCOI1j4TOyYg55IoWzuiMjuvSetHbepaw
LwN7w13w9y0TngFllqg434cbEDRSdKpLWhQXmWeW7VDajQ9Yyl6Nmf4QRxIeQ7vXSANjTpdlNF/c
4kbF43U5FFFhjpfMQVJiZ7x0SViMB2hPLySN8eAFjAbBiZyT3OGvxqUuTK02Pb/+AWq6iYDs6NdT
0ZppWrq9LpFP/KcZuqaETQ/Ecq6PB3opCSUWev+oRWFDxUMTvKNf4z0EBt67tbNLtQeQ8l7OGImE
+ztaXVYVYhhvPUpnPk0H068F6PKttPGer9syMB7fJql9EveV6BbjgBXwfEtttxB3CEfjVBEkrGU6
Mj0yf60LtsFNja3OmirfUzrTXtVM52OGOFrLwcu6+OZ7hqCfPoFae9YrwkBkpEE5fPX+tKORJQoP
v6afh/Q6u0PfZBsy7VIHCJWlqP1Aor1wJBoL1ZHd0IRujUDWzbnimzOHKUYI+D32dxdF1D7B4ef1
wmt/5lEH2aR4yFCCNIg+DQvuahX3hwWa2zh3B4mBBT80VUyOY7+ogiWH17qrXhidTufWSwtBe/vW
SsnvJPGNG5BStJSGMbocnxyXTFpVslFptDGdfP9BYy6aDnWcB9pWKWIE8UBKEDTiXX1TXLMdIOSR
7Yl7pMdX2vcD2PnNLSyiDjRxkTXo+xEk1idFMpjOBe7WcgED0H1vRqY1jrk9Ss3lnvLgutDRqhPo
U+wYmvkdOf2fT50ZRCEL1o5GGLmeTJyddgyv88pKHt59xWQ5w4PGTrpVIM8XkXf/hTbMgqUn+Lxp
2sFjjXW5ZyzrMkjOOQYSqWyvZ2Z6SieQNYxRiKO1WVjXG9UEQyfUE4G6S17moRBkUkZkn9kXZoHY
5DN2cktYA37cB0ZIH6zIGxHimt6AjVX64BH6CMHZ92Q9nfHewUZvk4kSQFg92sE4DlS8Do3Zv34w
TsvGtkBJ8l5WP8Reqzdk6nIRYHZDnlan6rVoi5QeTFuOJ9Yzds0eOxWUTFuJec9kEqjzADOmnFyU
tCT2pISGW/xeGgz5tQCIB1Ebab6LT01DuSIKLjzLwQXtGzJdM8Ez9vu2z2oqHhVO1t/NnCapz5om
rwJYUgDw5/NZTP+1CwH57cGIp6V6PopmOYYvJ4Q7v9wWU3yIGo3u3g9jtc6og+MDcVDZapahA38w
FrBs7ShrXaXOzdxLDdIPs50Pl5tcFLekmHacnnDvHeOgA5wg3vif8Q53OjNEZGppKvTqNvZVkc7f
rU50qsVrSXVhpQFR9ZASNfLfP2CHQyoc/xN9qVprRRiPL57+nwoAyw8ay7Bl/YfvFl5+nc/tGaav
DFE5mS75VnMctsnsSPhCB9SkfYVEV6MKW664T0hmDoStpUsIFwGBQEWEz393O2JUz0gPnn/E/I/2
cMwLYwewuiF199AMa7ocJWZ0j58dZHFBW5AGl31DvuK8qVUb3Q38eC/t+dP5tKku+VTgx0swy0rM
AOPf/O7rItxYdfwVOqRRG61tKJzYHgFc2M52cUR39N4iXWXUjH/R+ZgCbgK8bhhHFFWYNcyZLU+m
VPfu+KviQHrCin7TQ/9kWBdpwGRv536/k7TY1fggXbdt6BNFi4vM30TnZem0L4PmKq7socThBa0o
4VzBxqOErk42KIGiqaJNeWL5ZNpgy06sOMLcWN6oIfyaqpevTDPMLnFVYEfKg796clLG+TEI8yMT
V7dOdajtB6eXVM+g/DHGj9/Qt1X7FczZoXp78ijfbJpS4AwBCC+BuOAPY9gAKHpPya6uKETg68QV
Tc8st0IrTJFyvKyrXDK/a2qni4J+EMlsbkpuZQ1Q80WEzOKVFFLDoHJh94xRaqbBIuyaI3PZg7Wo
5lRdDmRkPgz0+6g+q1MzuXxVWZsQMQfGFvJU+MdNtl4fn6SrWbfIMYpehOIU5jTkxJKrHXYaxuC3
BqINfNHLB/AiwjAVOuzkKhFFudospgAxxzA7mTIMhQqjWezmTKVJok1fNG0hlOUH8lWE92LCTFkc
h6wZNE+q63aacVcMZHewZyMwYfSe6HvmxzUZ39a439EJEwyLTlI7luc/hrwcFHQ3zhhebpgFvXA/
cys+s6ipdyIpWkCySNWZRUkTpU60lgVAEk+SlDILw7TaG+cYZNmls0HBmF1rVw8eDgv4GsQfwBOL
tGYfQigpeCLObRflQSRtZagDPNA+AfVSG9lVDReNfm3v8vezFEXJPUuqSlozt2DpfXF+FUulGLjs
7+XbC7WK2ohtbP8LmFzUYOrHnJdb1BS5dUlCtpyXEbu7SaDCk47laBqEify2JXBV0/WYrw62s5AP
zUuXYJUg5uVBZzSxHVMhbxKTPsrDrcE1rzLiyKLJhM8Tp9BHIV0dnvSTTo1+wZLkWe2zozAmZQOx
rijnAbord1cqlLo48lkKDztBxRR3GZXgoo8mid4ziXIkhg4QwqbB2zFXoAzSCFPvLZI8MR5ISz76
Ovut8o8108PjZM+1TB3W5iij6ormRut7MWCVYqcq+fx93t5X2Sb08riSXj19R+g+1de3nuw5pKmT
waCm7ZEcHClplKhh7ITHPrRE77/MFhJfExeZz0qOJeDho0k3D1BWuBZ+UQejmKXScvnSgmqsLGLU
GMbHDEX9kkl4g4QGCuIF6/dv/DFeer2R7A7EXWJkhcyptGzAFEfEB2NuvDsd2xFIG/aY0DdMdAg7
vsW4UoiZM/B6cwA6+H/FGuttc4wernXBfYqam68Yzt5epymku2OoawErfAQNM01RnkJkFesxskh8
8k7Gh0Av5cE/PzmVdm+F1Hn6oO6nbxzVfmVz3lPr0QJEcndLFNFUJM9fSWgwSeG0lVMRouvNcQae
7ONwLpPyeSBGnVeLBENsvJcHGJ8C2wECWPeiQLAahRsf5gZKLUPV7HLnn6x2jQjATlq9bQBC70MI
au+O5etg1ZfiTkYvyUIiY8zSE0mKtiYihJSYsuO38OKyyAv1xBLMgZW5y2+6jTWpqMawUnE/uH6V
ORsgh5ipBwX+PdZbDBim8XVX6YsFB/5rqEBvFMXl5Ke0K1AsgVtJoOrPWu1zekJ8we6SdJn3Y6Rs
zrv9aaEnNpHX2bd9wrXhIgUlfTnT8DkEo57LxKKfp3g6kpsPK3c6rHwqgNIFfPtt7eK4IZJKE2Cy
R0PEPSdrLCr/mf2immYA8uOe7Z7Yw80r7Jqv37OLcuCr7fQ+K7lPuYfYaIspCnIDCzCw1zbWhe10
vWgETS8lDqhNhFIWtTnTbsvI6JRUptyyzlduwDInLGbYf30vCfhoBCb3x8KeQ/m+oz4nmRjyoLY3
6wGSMJBJE8ws5vags5IUEVE+HN80MQx1r48zIYB4u+W99YgfpX3cEJPgP2FGimu55qYKcp8BHHj4
4oXmSdHKJcV2hghHaFxiZEIYhSIhBnLf2t6CtVs3aqWlxsRGCVpFP/8Rzjtm91VfPwhvuUp5Oh3u
B/V8a0zr47nA/Nsyehg+5j2lwVd8y7148vXNslKxltMn/8jBYEDG6ZLY0xzJPpriRoz8XI9vy3+q
4jdB0vWsSNSTWMWdg+aNs5RVI/M16sKOoW0pJeTRfmR7FpHuyveg6tDCG5aS50VL4By5yg4i/LZu
pmN79SIzu3+PY81uGJS30MXDJfvSM/jT1mRDcPUh5PPDjzCA8z527WQyeBGXC6MvahgEVWMyFa4H
UOoPG3PkZWjbSRAWsyNpwl/Rhr7/UWKUzCsnBzGCkaA1lPQRZBNvjh6b545zRvHeJKeexEHfNS1b
zIqR5mfByDLXbniHSKzYw7F/ppgms1QSEjC5tIZ4Q5QH7Mt5ZH/TwGQvMMD2ht8dqIMVHaw1OG+E
1iNWj8RzBqzSbA5yvItv9KpH1vq0ZC9Ryf3fSbSNdbGTXFdTnxb821T+CZciy8x3uPxuOYsRThS7
k4BTS/7Od8KspT+Syb/CNEqAKKVpPdtG2hGag/TCzPPq7r68UDjCMatyhdcwP2cgHX+QOvNOGRws
5Tjixp7qf62rFstuq1of5lwOWsGvUpWIyG5Ahinw1j90QOykVvQBodjRmRCzoM2YDmJew/XWvClE
GbROhdtwYCJXZwVjDs5LlFJYPY6LIirLeqoSMPXkN0mROn4JHGMHqdsQzfomvzHLp9DtV1FyQuuu
n02gVetiLS4sA1XolZB4xgwC5n17GngjTxyaE7ZOJETPHNHnmITM7/W0SR772uWYHElM06Oju/AC
PHQUESWnqyHSr+FW8WNn2fCSTvj8FB3Xsi4mJrY5k+yHzNQYpnq/FhscIo/06yGukTnWI32Pvj2B
G4ArQXrNqcdoDX7fjVBC61O24ktZoAlcGWzm6ItXYOvsmDaFxo82ndffLfG4cZFtAfreWtJ5qrIa
MzHNc5QjEsBbzRVty2BADF8we01fG9xRf7oZ4wgOZAXeJD4BHUqn0X1L4TpxVH1Wj32Nxda4Thfi
MMtpvC0msorg5OsidP5Wpvx3EGiYXRref8KbHP59Tw+bRYBwVKgrUuBZKJPuMOMoXvRFdeZcC8pC
EDoY9RbH2OItZyd/oRAvmPKaCLsxhVYjimBH7i3kuLwHB0Va8NWcZkg22Rw2ysnVC4wgjdVLG3CT
x6RL96hvHDxD6oNBpk7Kaz4v2vjLgIjIioFo2ILcpt+kEhXxRmxtxFIwBZUqp6ZoaoTLfaBntwwU
WPXm7zwR4jHTpkVcvLUQp5EDwKY7ywh5HkTYCXiC1ygHysi86LllqnUojsSlTp3FbBzIgSt773rp
WX4SVNMbKQQPilLH1hjxHBSMb2uCBcQ/CHIdkno6NVxyt6R5E1H1Tpulvs4qnrAvWtZ8jji/z2nQ
BI3fg90h4kyOS+MTGuApvuaCFmsrUoP8jqJsprm2tYPw5IeBF2s8iqJ5Me7kMPbHUtOdUSq9U7Hn
a8iNtgjvcl2juCNNz53oj3TW1/dzwJHy/Je0hwkSS+q/Cz9A0Dm690oazTYBR/idvNW50SJrc9HL
2B2L1pBHGvmeTqStvOiY0j1nHWazunRsCJbKF4nEpCzmbztbr/xVQalmuajAKCRUikGEDqeNJGUI
KnfxDnpHdrwiWJPtpFzUAS4UoEAbxw8wQUbDq17SCYLHEqQQ4Uc/59itJrzqTkNAndZVcZ8nG9bl
MbXKMfNhsu4HGNDmDm4JLCNnxT8fRq0Ehmf/OU4ZEB9rOAmZrBMjG3J2YNuYbwfaFPIiI4d/VOkJ
SHz+/umd8G4Bv6gYyDbIrV3xeV/vzuxcdY4QlqYUuMmSJ2DVGWiD/onLDZuqzenMIGwsCNKDDTcZ
ynyWLbWrPh6LImv3UG0Rh+Y3kT3P7sVWYfeE4k0r0vrg7RiU8/7jlRbygHQzhCyH7ozeSuWhNS6W
LEkUJDBFNZbQ8EASHglPa6rOimbsKGjXNcRQAis1YziiuwSsxBRRM4s71hpyPe3MYUR3MiUdJpqO
dVrbHSqpbru2WwSmVBmlINr9ZcUE+2tMrbr17WL2M18omQBgG5oVHlEzFLMaQvVTcQEy0H7PGOW+
ijh6EdWOHi+2Oe4+VZowzsIcrVjTlGK+bvBF7NN/FzCw9272T1cRGyeFTrqJ020WtpYJtnMgAn1i
GUOt+5/1eh3mbK2DbRyRERSgbAdooK82loAjoYxSMmxY4L8/+Qs7mYAj68oC/OXZaVgr1TeVLmGV
/BLkngZ4LoQiG3QqFJmN4YbGR36fTjet8Ill0OcwXAuZ8GL+LBq/1t7UipNWfPLBMwTtq3Wzfowk
9NUWfwBFiG/4RxyoSuCR0S5AWy89gyqAq5N2sszOWsIRBIdoi5GLwFLj9OxRX+A2meMJwZx7WZxN
WugI5BqUWjq8Dtl/8HCw+AOBfVt0JGkbv1kS3eKnYpUeHAtqSMqUSQiC96CCEV8YOJ1HmMjt4+Zp
DkxPJJmd3JhFHCU9nnTSe3y1za0YPorbXL+GzdL9UmHLpIysegsfhk+5zKMwfkQvO5zkNuVsODNj
c2BcNf0SGSkUUcAj6IbKctRo6n79jFN3SSzPuF+bKuZ8ooScYfv2KsA3bjFYfDDb+huGsVRm9UqB
kMhBq78Zn6rNql25kl0KzjIGzcbv+9B2M+25p9tk3/DD2UX80A3g/X11f+DQe9NpBP2SpORpn+uu
HU2Ne3nZW8SoKw2fk2D1mMiVmrGoEzefvdoJtMaqj5rw+wM3rljF/lh1xBQEVoc0X+HYggMrFsKj
qOXr89EXtNXX3J0n3fOopMHAkowOfL0sxKHVPWpLzMfxTJ/D8u925/7s3ZhPk1KuKdAyw4TIoFU7
e73Iep3JdTNbHBaVTTMHWe7MsbhowmJt+ydJjYSNmOLngD+/MoVPQrMLqfaKukNAnXbUIw35HmVQ
6zfTshZ4dKUWoxENIreLy2OusOZt0adEE86Nx20gY1EXGqATbXHFnH6qByPmA+MK5JND3td8NX54
cyKHpKBDPkmJzuZUQjPVnKXtl0swzH/gCErxc+G7olwGBaO38fmM6aHlZgq6B3HK9D353dyH4vpk
6vzUcoHpcoyCTyk95XOG91IIR/pZPux3r0sWmcPoAnGmEKBCzQEa79fjC3w8xDxvY4jCcla3DOPv
rx9jsidW/emC+Jn33MRL2mEFuTLHILrdvzU3rd3WNT3AgVzKGHd69/2oCG6iAtCPw79c0bOpbRsh
/9CqlWFsZ9b8Cbb4M7N04DUHnzW3yNwrd4xXzUgsLNmE1vTqb6HYbpDUWeaYSt4ejAhqIX2pDL72
oT2l9x9ZJbRtK+ytM5+/KnPX10UcJwHpC1ccmDap2wF0ge05uTfPOkwtuFLQeX96/MK6K4tIqkxH
xilHbqJ1dOYtb7uoJVpTLUKJI7IiFugp02kqkKUzGEaO+2ZbQ6caQlIJSJZS4VHm+ovwUAuRzSoy
WSqZl4ay57bDFmXYfVo9D+zqWu+ZKZIVgnpLen5V3+1KefOvo618biCqlWr7FbzRYLu/ugZ39dlI
Y5HUZwIa6+pk1F+jBx/Tmh31qH5zh5dAl7B2h4ytpUGNbN+Wi1wENDbZOlIlZvuaBzVNtj6kD2OR
E+vsqpMojQxkgA/h3DHTl1fVMsXJdCj/nZVV/Ul2RhIghQsIW8VtLQ91kUmL6lOYi0dzQB+Hxw5b
BZIXY0b3jzdvnS8+ttWjEHomhEc85i9EoVg18SjayfVvOVvyOzHuNpJ24Sq9crFCBSz6pKKK+5xD
7nWuvuKBE/LuBrccmZakgS5X7SWP5NrNLJdZbgq145be/QyF84MDadrLVoVxdBKavzl/9hPtZW17
q7YBzPhFVNtKLaKBZSzkYcpzEdwnFpLUFQy+d6xbxstcEQ8YGdPChQgptKfSXKAcbS5YzKMzMrIc
VQqDhEESVJY/HMPuDzMBj3PZac28uwTUis0AtJbqdwxNtQnonyCSkxqR0r/UDF5GhxX+fUNGJ+Z3
hyXhccXMAVPYO3+c0OrrI5ggEyrn4NAVYzXP+x16BYcz4q/3pym+AcFGSTWygMEUOv2VoW5ngmH5
CKoHRrIpnXu2SxysE3T8wils6aTfEzqk1O2ufQfh3Y6vAhXqCMGB4kUcW28U7GYneYcztSiTvz2J
uPcrfERvUIjqKr4hBGcO3ztqsLZRDlDg3MsIO1wA3GfG9+TnxIcVak6VDZJsIJqaecyMfjicghN2
UmWWH/bA+cqnBKZeGK6nCa2r8tmIPf1PB6f0aV4FHrcuQN8sDUjc5A/vvNMqxo2cBR/lMiHUY7uP
NqMCp0tm4ZveB+vcfag6ZzBLW05t/X510NR7n4Zu+wmM9PfPU9Zm9j1NuOBxbI+O5NSE8WMQqryW
7pIvVEw4bWeA708S3rBsQLEqbQXHw5YlSy4ZZ3zOaf468g5hGlnLXB1sdAi8XMxJ/bzgY1kee4Bt
8Czdf71WK3GU48r0yB/uFdvq5zRc83GkM7uNO5fPZVH2Fb0eJ3zARb6ZqG5+Zf1Lx4zH2tN3LPwY
Bihw/lgohMH2g4MnbEfBHEKlrNIAQV6ZtT4j5cab80bAkiHwct6eHoCIniefI7CVqQoPwp2j9mV/
TXchlXqxE/e4vFiWZVuhk3HMxEqcUZjtLIWVX8FhFcsvXEegsSQD78NmOH9YxoFbyH3lAvOfc40h
eGIH0gWKyZjGMO91fVi7nkD9VUOSDaK6RPva8wCRTcv00RQaiKngBBJ7vflZVCRWX9r060SSIIiu
R7dZ5ROzvtRlDzbHq4nuKA0TGY8RDRoCFet02NyUcmyy8wodYIf6JvxvI8mP/1xL4CQDin8Dhex8
/XeVuoas62tFuITsIuhYPJXs/j22VUTFPDSL6xgxFIqCih67rK1cDRo6YmLUfzL1jFJUKVqENiN/
e7wLjxvmvj99NK1fx3j60TMRn28wyIfZhH7r5Pm6YkeQHv4VswBHrzTPqijT6NV0kSOAOq283ecU
U5wm1fZP1CsGFVavJjmjJC8DcgjloRx3Wx46AWFUqKm0ffMGhAFk0jeNKdmgOuEcjOijGM+dcZqe
2EV8BFAj3AFzJ2yzRfXTna6rEe4ninT6uqfoVlrV1P3D37SyuIQTaZwax43StjOtb6PGkhXsBsco
8M9XgR38rdo1j/wDRAI9NIwtk2c4dF/IzHHdRk1mZ81/ibJkiPP0bxSAQ27nA6a+OQ87m/+eLvu1
dwq7s0mbiTyB42RD7OlSROgZ9AK/rmAcfAG3k6J/Mvk6zh0nncFCrl76VMsZl4i3ODQ0plDuz58w
MG9seZSR5ATrp2EwDZyYGrV4wGu7ulZxkdoKd6INNKValTUS2SNV+BilvFJEfwt0F10cXQ3vEGiD
r+jLJtB7Si2qwBiXOB+Dx4UFOKIBhpIWHrZKoj70yv2Hl4UPmaxP0v2hwy3BZH1wmZmVEMuBxY9L
nlLZrTMktZn3hWybpNX0s1Br3dpe8kZFdd35UMLQewV+coL8xnzN2j2oyQlTVjbRmLDP9f+7EXT9
JBln3Ua0f7LwcRxaDcEy3atVcyvfjxAfINWZ6cZVJLspNl8dVAxhSUThscM3K/lUcTDDhOzjZB2U
UTfEQm39rJCNoVKoQ5MHBncGfYvJ2U3uImza3YOBkmMwxj10AKxOiOcskw5fErs34u8MxIe02kQA
N0rSkt7Ct1k77OR5YQwmPJ6ccxDQ/w26wMfQuj44N+ACBFtkzavHYeYNdQ3YZ4/yzHHr+v7SkYaE
53OgOCG9LPOT8TUfyEWzUTsq6rCKtWuNQAUUIvuchegOmx1rmNtEQ5PnIsvUVX4bTZ9OybA7ApJt
7n0OD+B1YF73sXK7S9BFLw3tXDqL7O+y8T1H/IIVPfxskPmI8k36BAVBJ7qEI/EHP4iPWqE3+9GR
RyC3PNy05JlhiHLChpsVHjX7qRomCAigNOMynAFeY9Bccf1eyMDvOM1/2GHnQ7dLEqTxfxL9rrXK
MVWQbIBwuqf0BX+l/3QTRG/JPfg6GAxGoN9eErohK6hnLBq9y/bqwLadICpHGUD6VAchTfGBG/cd
8ObVPKbP1fydXXeX4egnF9y+o1H41AdDlkenEnnhfR8mufk9ut8OCo63bRZfTmY0Q7kRnf7ALiMj
p/MuzYCDFrdb+EMPaGblV1L5BhXYgXv6jzKpOGVJzwGcSdGyIITRA4dK30FIBoSRlMqzWL5KhPFZ
n8cLs9ZaFc7WA4Lqn65bB5KTcdML1aAH69VW/ZxKwhCb0TpB2A1pLzhLjiWjKjhbrwfH3KIVGHGX
GB77/1LcDz/FzSaoq8q5WVdHcTxyJ7tMMPYZLh2OK6RW8zxPqdSNGIDw8dqzjIOjFfr8phA777E7
u4MyIGRgUy+5yt2fWykDGspsDxf1sLwXzfLDNEcu7S4xunGmVanLhKGqfR9ikUObZUaiYDTXSHlm
+S+uRxG/mei9U/oCLxm/w24wX0sm+gURkvNjSAQxK8Dv9URp8quWkZKSCaISPBnBrXL4WDVF5cER
t4fvcJ94ueaayJiuMybkja40J67gZY1nlFXuYjUjWJB7/u3kR2CS+GJa4lccwoLUquZiV0QFPi7b
JVBNQ8HILtcT9PfpJg4wgUI8a42gaaj8jSltjhviLvwEXNNjBGwFmg2aUiNMSVG0F6QMRqcI6sfH
3PTkFNhqRzdswbDWZazkKu/2oqoMuEfX5PIqCto28boDdUCHE6283299Jz3ga5MKTXcPTNTc0J6d
zogBHLI87OgPZcphwn8xW9RxmoEgh6upE3qqLDtPZOaeaeNguCEpS4eJEmQp/uB4lNwSyl1C0+fR
7vTH2rubYYQZNDYev9OLWzTZrXMM2QXnhsj/w5XTrLErqd2k1SvJJBnn4g71O8lbAKQsbpt3imE5
+zjOhxSNi422jfLbhQCvs5LCocNQ4/usuBgQWk2V70RPg+JEVX5n7VkKAz31izXjJdZyeNUFTyya
c/oTbU4Hu6Q0M8v/uyqrD410hcchtbtOatONryAKBZv1Lm2XrFovJE/CpurYFveHkKQ+GGoPtzdU
x2XCknDyYI+wy9RH/IiLExaEbEItmp+0HWP2iLcS2kpQ9vCUj1gXhAG9rV3gh6807sVIICXykdSr
0iW9/mMErv+7FtbAIN5F2kyFxSmSF08OgRwXntmptpyU1sEYBSLmtg31mrht1a+niP/deWkVm0Nr
I81N0Hd7e3/GYzVRfOAPz2XMC+gLj/s+FG2gxHm9XSvfxXBZKUcAHEPhCGjNXik1Zq5jJRFNbuVJ
w0Ab7VMXJuEEz2QjCBU9bMXnC5KdollyUpQCDoQCeOx8fvpX+pbEXgqxCjmV0FFa6H0u3tiZ9W3P
DAyvSAoEyETxglC+VcYodKCw+r5GnBOlOhSyC0+rjwtECgyL8ZG7dPJ5PBdDMg4us63/P1C56DlP
QMEzhw9f8tDxkW8GgWVb5sCvvW42Mrumy5tYTpidhdlCMH/8KAgBMl4x6aUQFQkTLCYGsM7shSHL
2UNuXnq+7zc8OEtBLjMShLl5fppVtDToOKopP0FLWiIuzY6+82M9A+tiyJdlHuXPuCVEa9u1fwhf
1t08NSqzSBykaQ2py+ys6mkNdUm1I/ssA+JQJHBjEGLLaTYD0oFUFdAZU6yUYnu3RF4u0tcxn+F2
QUXy3Zf3QlI4qKo9FMZlq5Eec9/TstiLQK/+pdpzLZ4XFD/+cVBS6gBat9L7gUBSDQT9n7HHDCdW
9og/WhPscUazi4PZ05Y4tOi08oSFSnlh9L9DRR7PZCHYUZZEAfVomAsG+Odw9J3CkBCAf2enqkxf
Jar5p863r1H/D10bI5ENjakx7kCiJ++9uGdJAWNenS1rvGOtC6V/ScWY2/wr09uw2Z61qB1Jpxgr
C6Klc6mj0IkdPn3uAFKgeMv8WK3WfPeS7Jqcz2fLgHNf/JiOhEMteN/b4/2QNzbdOCKzDWadSXDx
h5uQ/ejsKAOIDc2oFVQ+sVZ2LdNpqdWqy0nz7hrpaBraFHzl0CsDmkk/zi/BrvO/Ef5ob3WZm4DQ
D9HFIYgTEGTL+SGRftW8jbxwW61StPWpaJfj0MDBYHyH3HmNovWl2LRbcQT84OJrFUcr/1yMGxH7
vhy5ZV9pV2PzqYhGpSpeB+farGEt3fE0WLpTxmIKyy4oGBNU8SIiNaypKw1hwBGseBvByFVLPHkI
Ns3Xw0pd2ijSScfTrItjGe8BjrGWOx+7nj+xwXLys6hLlvSFP5+2kh1PQq6fHynnFe4E8FbAT6Ce
mYqdQYYw/l6ediIRxeltbCOup9Z9En3vuy3bkVJc/4LuBh3iNa1hLaktf9gvSttqU1VxS9W5n5bW
La6Hl/I9Kf8X94b//qV2Qpmh9XmPmYIWK40sj7hgB3ES0PFX4pR1Gd6YkO9H2jN6aCjZKgptUtXE
YGbuawH7PkW9MYZSGa9N4Re4njsUz6xrFbAah807lJ6EftX5eUmcPxweb0S6y7vFBMpAMPZyfmCG
xwEob7tbJbBqMKvoRnrC6cDJp1HKqO0Ml9+la6U5cQlIVM6UjorLs2V+cmH6RVMlQxPUayQHZDOA
/Xj9/acSNwy3Dl7NJp1xq/tQE4Mrj9fyt/acRlVLCjMXLmayMpLlsQJIlU5cPmEdJIUTzn+7noJz
7RxWU8RY71bjAb6skdqCH4tp8MCdOhRZRBK45sH1ZB78oWb6fXqd8oL4fEHo9/hxnegNBHsdf/p0
89arxoBpnYfJs0+MEvXBFKidFqeomqz5o7qbViJ9JpgOzcTAZpReut5GhU1MW8pnq84iWh5Aiay2
h9rMb0htUUdqzRq9RP4BdfkpvVHHB29OID7WD4cahBfFyjq2aFEDjZh4w6ZEnlLw7qVMFz+yGZa+
Qstw1P4cdPgaMOYyRcGOmzJScoQOb03XR6Kg4um0eIdUf3FNKFObtNlv9NL4AwFuk2KDM+CxlvXW
ojxrKc7U9wqHIwyoe/zUQHx7dz1QJkswMhrKYMKcn45afaKaWNxI+/eoVN1RYXnrtSNfZOwtFKoI
CA/Ibm33rV3flkun7880S4JlfTzsOCJv6ti1O5sBz8dpY8fbS1zRZQ5NbgAKBI+oAGwuKIAcOjcv
vqzqjYGBqw/GfT8Wno3i+7IWE4uIwapvgxMxhguRImujwJKNmCT8EiTOn6QMcIo2VH8AHMujGRy0
GWnvLfbjZAvysrkAVv9bSHUfEdJc9EzroE1SL9ft97/Ju2j+Vok8+4DtlzUNTyXTRBQrVbj0Za8Q
aOSWHN3RoqeFruQ+E/LEEKHzFEEV2iMSNkGRzBYzqPdetjg68dWVeim5UJ7Y5cNPyHbJ/ATVR+Gh
rv7U0x29JISMLV83uNhunWQVKZDsr4j6/Lp7vWtbD5oR7qBL+DBzQjI3Jy1jAXRwTguXO+R/teU4
jAXlwaKj7SklEY3FJt0kAH5VvmglCqT8jyE4D5X4ZXm2NhdLzOIO/yqfWIwRB6WBk+qtI4/sigof
IbXCusZQjBrU8gwhFQdvq46sSR1Tp6+7i/U0yp4+1n5ag27xLkynhL+wbuBxog1sKX6kNAl00hv1
EL6DDAQiwvrsJK5pQQKcZgadnaXZjL3GzMIjq6O8JkFdWh6XD2iJkIHl1YHcTf4Wm/kqgQLaC6+y
lRM8iE6jdNcNb5Pbww/fIuBNMV4GQFrpcqhdht1COXceN5MiM1S5OMIBnbda+b241iBX8shWOd1K
6fgm3by/hcd1XHabHXX/AE8HwWcg39SaoFu4hKIZndZA1lmt391ycmdKLOFo4z2auoj9GxQh1wDw
gnzRO989DM5m3/bibQcoW8BRYHO1LTep2yHjh5dH7woYmx3aMvM81Hbzf3yWWoIWFKZQCm+FSrYn
me05rQ2LLDMm6U6+uegaHwb/FuG1E5I8R0RF6ebROMVrwlXySXyiQ11lBZRZSxgBImupjQaD8ise
CbQFuJBg/k0WHnVhrQOFJo/AT6fFhxVOsHHdtHycboK1cpa1mlak642VXOGC0so5ZqGg6zAeR1rj
srsfM4Sn7PbSRcyelHPU9iWAWaUervF+bw5IlM4k1yj50YeD+LOPCgvztKnHV2UQERVozA/knlah
rHOtH5VmfnO8seJpuUsuxRrSA1VYaXeWFI38ZkqRY5tf3encZMJs8cUXDiwKpsz3M+xAQkjk4sjt
ad/YH8U6Y1ryTxH19DTNkRS2zBPUc6LR2cIabcG1Tg5J6G/ocQum4sW9tdT6bS3fKt5C/55XpfHH
8wO9PZeOrdOHGFtPeYatbu+wIv7CdMJBe6dyZA1H1NPO5vKr6wNUGnxTBbza2yxSFaM5O2ZapNS9
7B842v7dyEJoTFqzYsv3E/G+kckf09Ef2WT9Mk4O1fX6Mnmjnoex8x7KATtfLHDiQSXHxhesKfvk
MbIEym50fLkCvhVEnQazOuvi6GILskAQOS55FS881NGBpIgMNuxXS3oWEXSUw6dnxsH4CWher37j
cN8Gngz4jp7+boLiNKiZiaQg7swt1h0QTFwuczTv+Hm/WIGlANMqSLmXKHXKwMiWosuqg2sELVY1
KlLoxU3/3FUqCJnYbRtGKb4An8ZCQRHIb0WwWhQLItcI5a4EeD4nuSO7T8zFMgQWWGZ7a7CCkzQL
WirRbZ2eb6ihHJ/Xr5pDviaeriqxRlE0g4tAQ0SvwfOIy3PrKmTdJIkF5tucDu74IJzZ/Ot8z9CJ
Nx702H33+nLJPmftH3h2fgzTm51qfkzY0LkCipzyJQahaQrP1mBhNU2hI7TuYscouaA1AxD5Zgvk
WCC7nuWoA6pv6GUA5jTqUU6XMREr06I10uy/cOAZrR/GSz2Ub4MXIHhyrk7J7ipU4Bi84LUbl2Fj
6ujg7w1E22ivXYczAkLRNIVWokufT7wTOD4/MVaMFXeXfS4tAPWA/PhEwgEjK7muxSAXUho0Lo6U
xQo85MjZAfoXmR34Y7S3lTYNJt4nFAbyuyVivw+leK9IZa95caSRl0jnDD88ZKRzaVOILWq/yCxY
R0DIPPPW3KWL4O+/y+C13uygIBzgeeer4IWsgwYLqEuxir/kM2v4TiEtmNnwh9bQiSEj9hkmspMZ
2KddeF6UEBLML+ix1CFwu18Yc/EN/YuuwOmQdE5ZVOdtgoVbIyp2hDpTY6yg/K2qg9DX+FG3TrtC
n8mHyUWtIKOxOqtq56aZa+U8zUBBIt2XWP3uYqLjWlJu/fUYRRJydbPeuKeBIDN7dKDIP56lTW26
XeR4Yhu9Nv3T2N12th1huQVopffboi3BD1fD8929ecilxDYl0h2lV2Yqx6Uz9oVuDKsBTIrBhx7a
2vEWHUhn2PZ98HEPeV++uZPiLEADktCt9fw6q/a/zvaYvXmX/ihDOGfFF2bzHk5nl/1KIZskSdMv
eyTsbAQBoomvqg2/u+OjMO+k97gfBvhcYSc9CWYhkWTSXm/4SULD5TCBejbj63qUjCgj9Gjygw9V
kV6sP1NekTLmQ672StEGfXRW4JI9/DjOgaVZwWTvQF0zJCcMhx9zN3RLOvTl1g7jzaij7dlGHVon
myCmkErNTiFDul/1+OtppWOasZ1uCPQTIj9EaVs6potR+CepfiWdo8cvgLrBD/zPBgUIGaXnEiT+
3MdisNLL7fETbxbL69j6Gp4+cmQUEfAXLd4PDGSl5Ih6HGuJTcRW6ihG+iop8fsUo8z3eXs+Xx//
Yh8YsUzr8DypD9S6yd2dXK3RTHW6LS5RI/TT24/giusVnG51blsHBtA9HDyviPHZmoFYgjPi73mM
1yiGRkMlnGvkEruwrGu/y6tMNiiWUDj+VWWzts179VA6/V35GEOQbnoebI1zOLnQbugn5Kqqa3tH
EgP5B/2ggfq+/I178sdxANQ8rkCdOlhWQhT/WDdoy0ymCNPYBo5oWXIzYaEqEOPcPf8mGxRjWIuh
+OF7BslrMh8KDftAV/QVqV+CM8vdbwiVUF/PYOfMCkALCCFPGqMvwZbKlI0OthRXsTYACfv5x18l
RZ43cE/tPd2IWinxPMS2UZz21ChsIs6JJRI5RrkvnbhuFP6z5ATN9KQio2ypSp9SQGTgeXZvUJvr
yu6R8O6mkdGrmMDtvvMXMY9YZLSs1H1oaWFNRnLO/hrdsX5PO++OhRoaQpFfRidyJP/N7cK6CLue
SKJp5kkjaCm7SaENnHsrR8OiDbTli/DwAaFKUM+O9ED3FFmRiGJtFLHdiqaDzrizp81PDIgo4ek5
acw3mhj9QvCC7H1mSYhvnbEhOYxYvp1O5xV2cEm3OAGagK/XjfDYBhEBPNbkIK01gWNHIsbm3PHt
89IAtk6nqfF/tV6YsBWCL8QP3EoYqMjHD7yRe7Aj5rKNKL9iG6G8KIfJspZsW2WpF3xIPI6bgCuo
DcECSib9bauiPNoUwB5g0sBt32vkSDYS2oQ0STqMoHaESU7Vwx4d03WGGUSYZGMV5sY0XlWO4A/L
BmlLmzTrev1Mp9Wb0gyHnrjL0KGvKorqFY106YgLzh+7Qy/lUkBvryAjX6U7Mos50lOP4hGCTSFG
hk2cqAN99WnEDBWNgWae/UmMuXh439URB8PzKu54Rccx7UbA0qiumMkoZvpFF6sCV3joNqnvZYWC
cG05HPcnjwoBQZxOh5SBhd5P2gVjVj6fMilfXCra1BmKqUnjOf3ZbRbGgMnlm/jMtDhrBiQCtIYF
VTpB5b0egBYn23zmGdPCRFzp9y+kl7pVFRrXPfwWovM922s0P4CdmKhbrjCRt06HaOAPbxaAUjAW
vQwPqgdin5Ay6vfD7RuPOsaaAZdXs1/6fLcxHtb1YCOShd+MfuGGpej9Cccgo4gXfDhZsWXGSH52
lvtbtZ0ymwDaHOWeexy3aPnIEf69OH1O9JM9o9SMzd/AtKdHsBM89jsx1BZDtZaURXiuuedDte+M
uQfINFfyGRNBO7x9qU6YipkBaPCuot0pvghSxveDIcNmJ6MuXtt9v/7fUeq0zaxWNlrSvT4zhY8R
tSQEnoBQ/MUP3Xzh7upxWZ5hbp01eoaDJA6+rLwrIv0+kYIroU9KjID6K4zMUv6HESwyX4c87HAg
m9cw9tLKm44sSkSGWNzzWDy/nYh3jOXEBSf5kozcW5IScdZqXvIT7wEwFE71SbJ5J6aI0pNxo5aq
Z1mLNIVvGK/UQyxXNQv2rE8of1LqxnXSjpW7mnP2qlXzi8fcnDdrA+/7dzHg+Nd2q0U3cK076hyT
wbhfjQiJ38P9+otpfUkjHyqxWZmh10FYtqHeHyzpsj1xKmjUOfARmEsu2UJEJ9w7RbQgrCUoiLo9
0qqExxqhcj9Lj38S9vowjDI7xQ733AHPnPZaEDu1Qd2no1+2xZu9QgGRxnsZS7BmeW74uUQWDMeF
kBqIaHbRE4qsGINjnkvUHgEjZHcUNhP0AT/yn4KvmW9y2JUhvkaehVW+CGfCYyqO4NDx8lz7KLC6
PIIlx9L6mg4VWmO8c0/Hm8pqcFcFt77cTjzlXf5HxC+SQZW3V1i0An1GmkxFRGZnp6Ssk/RsvfNT
cNu+2y2z8T6MR69wFl5GBIQTcDHXnpMsPWcG4Ok8Lom3U7y6p85VHqBcF6Vm2qg1p9BrGcfevKhN
BbhBce40rSGU4gZRhHdTvXq/6BeF2sb1PPqHa1df+j0D09EQkh1gXUfQHHe0rOkhuedd4vPIgCjf
KaUpPKEiqsgO1yHN069kYYhS5a7spj2Y/ccffm/hnMccSjy2pnGm+P8y2fs1qbWOsntlSeYJ3Noz
uxqarLh1scmuT0+CdlFjgjjFYTKMk6pQnHQVNyZDZasoUHrPezNK3PCTcwt5Z4BRA9b2P/26cQoh
Cn6yxpxRgKoSVecVwp5o1PH9p+1h6wNXk9ovq6B2p8ckMBM2nlPiNYlVVxd7SqXZRJ+7yc34jFpt
65gLqAteVyPzk19bM94teDW57MXBFOAK1H/phKACvkOVxAIFT/A8QmdyMApiaenAG9DiwMGsXQIb
ZU+zuMukp92w8c4DcDxzzYo5sQn4qKWE472zU8FYna9RgWKcm8ZY8iVVDRbWhBGRkNFgX7q7GRtd
vuO2x5oogYRjG5w38NCb2gxCQgBCNpXazpq49N3/QMVsLylXL9/lkRU9QRNlGlWQ3/693gV9b5Vf
tHoJEuyOLKWrm/mRPqKdULOY/CN00tUUtNyogPz4x220kdGdRUANsrlVSRaaLhVSli8LhGEiZd5x
1pushPk4YbW5c14qRk/QHvd/Y9toyulsJWluGOO+z/JPJFeBoSgdg8msVuNAth5TUwIAJ+K7QmUz
rsutAbJ8UmG/2WWrJDRm3tgXaQsbtYh/SkaxW50xgCoRiyD+iQALwHOTCiJVKbNdqMjnt5qWxj3j
MeeQJeAlp0XTJb9H8F7EL4Hq9+oBPAxg8C+CsjT95547M91B3Tu3Sd9hks0rBwO0eEyq4XymV39T
FauDHJfhPcPcbtM9wyHwB8C43Dlw+564QV9ndUOv4JmtUHIIHyxcWNZ+5Aim0AizAYqvb8ldpVUq
KalArGxFQBlet+dbnxWjAXrQ+9hpx68A2IuEGyGFxlujBFlLWcdVaUuD/s4KU/Xz1qfqwXraaOuh
DhrlnPIjip+0YMVpKVNSVWjnCoDkHRfc4UT19q1Sfzi/ZUav8LBObDPkVkOACCFJHq9gBfJy3DN+
QaCrq+rVzhcW9FL1bx+9Mr4XHZOlYuUoKu3iBxE0nQuDogzQf/CtV10LVS4E4n+VwLRMgkn4UBzf
HUfvspCigf4qC7mOvshbQlf+OWg95DMd5dukn5Gttl4FkBIH5cNf6V4+1FQvB3nnMOTGSTxb1kNK
YNsoXcKldQeNNPg/86/A5kH+LqUEJt09XyBT10wsMO28RpjjZa4u0Ox2aZqneZVHCE+ZpIYf55z4
cKDKMmfA5s2cAMmAiaJOmbAZmpJfe2zOo+11nS+yNLwLGI4evxVs/XH1wJFRLptvqap9hS+mcqUM
zgRC1rkOQi/VDt00tGKYZ1J58QqyZL79gDx7jH1+hNx4Zr9wBfZh+hoBgU+L8wMpndkkJeSO2blw
9oFAEcyDoeGISqqW/C5fvz8ibc3Y4XY0AmxdDyehJgV/hVHk7mC8TWYfxOWutRmBArG0Qe7JS7Ly
jaDZKgxV68risEd0toeTnGCdU4CYJokcfIRlyU9T35HU6uRhk/1GFJ9l7kwsjc3tjLRub4iNEnmL
lwAj+d1JgJYExLRQr/jQLGdA8uAOfOWnMomfk/sZaxTZd43gLNbghfGrVApb4A+7BA0LTU4IS48q
pmYe+X0+ymC5usmZPwYkRkBqwoK01lnbhFSmNAf4WSLJDM2murJpEP4zsX0qupRSLRMT6lAYkERA
nDoU94qe7oN3RO8HhZKFyBLNYreZwRCbfaH4FN2NlaH+4vdcszVbonJ1KH0+rdJIN3Gm4LvIbSgI
jt7D3LVA/HriPkB/jEsazT7IpfVtURZKhE0k3FfFQNOXNYA0sfs1+4+T6BGvwvpTzDhsdXp3KBCd
sBLit29dg+0h3oq2+Wz2mxGKjWojDbtyUJdJQN7J+zQD4M31dSmkGrjxIdGDYjtuWTlnPLDKZFcW
8q1H/NHMgf7PGm9UIdkT+szy40YDCIglE35/gRQWmnmpRzegS/hpyFuhvFREzyz8MoOZSgkpqwMx
dErXcE9GLUmPiBMp8+Bn3DSeib4YXttjyRZYlFOJ5FHk+dnr/qfkab80mOpmWZJwta7AmykDQ7Fn
2DIEM2AcCR2pJF4V6ySAxTHfsfvGv25H0U994KSlsfiEPA2rzAymY3GKJatpvfzTRqM+aMuGszK0
2vt5lMoRfieLquvoP5hH/jZBaIewXaFEUqCKiuJUUr/x308IKr5Uo83VPSmefuyL/KVWFfQwuhgP
dVjYe9GytVOfn2NdhCVnm7cme+dADdlVYE8GggfEBE8ekwz7+xSByLRLngDgF3HrFGKoazx7TZgY
wIScCUKpJn/d7UEamrRa5qJNDvE3+QhhJPdK/MsrIwTgN0G6zLp7Y6DJLp6nedesgMqsye6CL2T4
zEiYNLC3UBocfGK0xcRmRA6tH8a2yzs6r58a0hdbJi3O4kpQhx0FditzJLTszRvnYSCu/Popfy0t
jPU8/uT7O3RuHB6z7Qmsoz8fLJDnp8wKb42xUaNDPdPcfkSBtflw6+29YM5qg1bzUix9K+qCwPXF
PeLmIdS4tdKGY1IajCPifaOyvuUOlHm8iZrQQmwclp+tXFoqdk3X4We8HSZtL1fQDVqShEd9jmyv
z0VWCPKrhe5FsxBDUrXWvjYnuKKU8uS8DnC+iJhQ5+3oaDM8bC8rVv2bZYbAOZEkWfcqfOg/PNdu
vSr14fvVHZa9mQP9IbLG7UBUNjHjnR9tV2ajRnC5F0Z9uHzjXS5vIJ4IlprGyBlgU87oPFT+0epi
PmeRdtF5GQs1m1FXkFfG3SQloMX10FKTaaKMQorqo0dJ/w+qU8/2q7rvi5+LB/vhNMUloWg5KpVz
hI/beyx3J1jIU4nRolbA8y+PmVdTCkP2pzsCEvolpI3V8Xb0RzKY3GEFpDRJ2IjFaBM0tg+nrS0u
crzki+uDSwrqDKdbtrJM8kpOhIXGGlDEwzldKIYL471Jg4zxhWy6Jq+U7s/gMBboXpQoLILtHn2V
TyIEtq9EXZZUpTM3KYyvXig3nc4d5ck+kaNE/Vf/q+AWIpRLP1p70vcPRgYU6Yz78HnEX46dID1X
qOIlJv8AuTv+eCCf1HxzRILc4b0w/TVsxzwxY7dEB98q4fsEr8vpcaSMQtqjClWnJoOthBbx6Y/e
LlNOvhAS9wyUSSAofHIVFuV6ATKWMRPEqGRMZcMaNVTnnv5Lo84zZ7he0bjuFs3/TVJixGTHS2df
f7Cpdrm5+uvfxnxAGLXxbNvnw2VYUlGx8u6+GSyC3w6wH0WlWo4hdtlLJSTGDNGVTIvkWtxeX7sY
B2d/m7XRHKeA51apTLOJdhlHS1m2SnuBq775w681qoinQLgZyj/Fh+/S+xmKcw4BWpu/bFQSxRID
EzUqkp/HsbTOCvNhV7uTTX5I67P5vv4t3Yj8P1Tv9V0O2mI8LmzRvKW4O1+YWRg5Q0ilzrhA9D4i
bdFMIh3DDz/+eVy9Ke5YJQ51u247Ksq9zhufsnaJaOptpbpJ5BYJDZMbYKSkXYio67OFxtnK4ZUv
NXIjy0Je1r2lpYM9Tmu/esdFyUfgAplXvTmEER4s6z028E2xEXPyjo3z+g8Du6ZDybN34Nc+Ip12
iW7RgM+gh35upCkeZufEhJjpkzAaPNuEtZG687vUk3/kKUErxjZsNp8xM4sZFSJj07PuQl/e3104
NFrJx6u3T0bBztdfqfg+wd3Gm08I407riY7FB5KriFMh9JSbSX7RUzmWacifDfDi3mDn/NUesD5k
CnBL8bj+UFTjBMmo4NaVhLhV93AatUNXoI2vzY3muFAQoO6KYOgnJe0PrCnC6c5N/GPskgbqhVop
f+t0YS/jtb+1n3akevAnYXQz/TQP7b9D9t40lWxJnUIHtol5Q5MIU9O77Ln7ta1KKwpXMAX68F0I
FhRCrXP4w3ucnqaS9a8npUs6/BK480jPhZhOMnRlnuU1riFVyrgoTC314wiDpXsNsMuNcpeg0v+u
Ryx3ov4SnBsooD/NPIkra9IEvJxmIJCzNIZO/5L5Y0mtlz2AhEETH8hNTgFHtuWOD2cABBGzemIn
dZ/PqQTYbDWjKaey9B+3mK45EWx6dv+3wp4dIcNq27tAMB8HyO+vyBvADN/K2DML78GHNSyN/cGB
5aoV0SGtTLJ3MUMRcagAakJPD2cpFsXYjRmkpQH7zOl0/DDTXvOH1LdbYxjZlTKFin9J7vT4wbVE
acgS7oj5Ycf5XuBGU000eJIbp4yeLwRHm1EDm0NFegwMp2YKX76aZVsKWAsMzVpyMeNxDoXhY33F
e3St+FU9lqnIyjNlHnpx5raALCnWiRAN2P1TzKH1wJLRX7sCtOB0agmZc76LLJb7KeiZSB9KAO5X
NflT0VmtE7LzurOOXF/Cw/J9640iZYFaFEPpps3JehbxQnU/uPoZUTOrGmGvbMPU04GETzUxxd+w
glcsdCTo5KCVedVvkE5vulb1IpHuGx4Ilxp8jVahJEEe/4JE/DRIhJ7ilswHbQEUrHiSw3TG5YMU
UBS4EtTJ8aZPGLxPKaj1cabj3HITx3iGixYdYcohB0pmpz4SADt9FvleTM9bUYQEx88TcwV7NoTe
AT+swH9a0WH5bu2LySEQp6bhvZPzCPMN413/VTM9b/Ei2RseNc31EIgqlyNZF3RQqzCjW/y/UuJ5
IF2nnHBOQ9e3g3pQyVdE0GakVjyvbyNTb5bojK+33EOKO3FK6SDsrHfkrSywZ4L3G6HRml+JVjg3
vL90/2DBphlOO0601SQb0mCG4KyNNdiKfxe4dwsgooyeEE9e0zSsqeWOtM4Fh1cL0ITCtnRy/Ikd
EKXlrmEoM3oWTo9KXQ/IZlacahSR16ixmxiOOpSc1maoWO5Nls7rcS4/8iuQwhQhSq98haUVnQpA
QHundG9powZ2jqYNpxzhkcXrdh4GbR/XCpkXi+sleaDqpzosI1d7NDmMMyyRmY0Rl51VCFeBVRXE
HEYv5RHeNDboMf7sU73uaTpFGv0bRD0+O9AJaJ2uc+FPiT4w+G+F+U170/MHqtm6qxG6JMMjRoe5
8LFmtqSA52+UuWjVxTWkuXVFFwTPyk3QgrOJa4Si+rBDbUBdHNQDm6f/d0jl0ldyuqi5+OIPbgrS
p3e5jKhVYctlSSr4EuQtsW0WyptM5EUyql4P4hu/5vFfG9tfy5a7CE2XBwh9q3NzLa8VBNo8Hcya
fPOMkgjjAEmQOan/7Tl9nVVB1fhqvJv1fz7wFu+ZSvQHg5NHtxVdj+aRJR0zWed9ixsE4VTYYIXI
+ec1j/yTh6SJYpr1hQWnxCagEPwZsqMNEYZRNF6bk+L4fPFr5SE6TeaMUbFNt6Q5eve71AtrodGT
EeF3QuZuBKgQXKOvrb7NQbnhRQ+BIzJXGE5ozhn1+Zoj+jky0xpYVde9UF4jn98pfDf1jxoMxaOR
0YTt5khBkFWv8H0rKiGLYk+Jy7nJbscIUgR8Mfv6s4pzMx8r7D0xw/Mip00+2ra3F498N3kYhicC
5qkADjHYOycQD3cxLgyglHGKBWr2+2NStf8xEXOjyKn4hlcCnuCPfLV+Qm3HP6JJAjyBczaeG3XX
mmDlYBfUEzuBfsfU1KqDQYXKXJ/Q5EiTd4srSh143E1dvyN1oo3dCNkucTKcbUV/qmcaZFhNTtjC
YMX3PGwxev+hjgANhV4PGQgqbyONAJJGrBAdmGmOxllVid9+yZc1ArD8ZupBErvtJUWnS5J9wg8F
3K3m+NLgwJ5U11jFXRQW0m9pPmmfZM/9QY3vDzVN88tLF7LItU2a/MGcuYZB5uQly8gxi6hbBOh0
RIMknxK7awrr7USh8IPgLwpMQ+Hr/5GyM1ayPr9I4P/X3eLtYVLmqAPaYGBnICt8j8Q/0DfQKToC
zBXlzKlveWXK4+SyBh52zKAcBR8JCbRnPS+6SJWxC1ZPcFW23Y6ufOcFTo5Jygx5gQ3s/zgZXkMU
32xQTHJMdUs9efxKifcF+bstI12nwatHFLi4KmxUyTgIVoNuGMFX78rbpGdZjG0QMWZ7W+6wDwrs
AZnE29foTodbHWObm3CJzx6Z6ZyfERMJXv54LLT3sEkw2JAFXG7bOI7/yWCsNic68hDyZijUrMVK
4wXYMJqro0ZtnjJGi2G2NF78fK/DzDFaroobqwtjsRq1SPDkJm/Gg6ha7jdbAdthBQt4KBUwzAo7
YWtsayvGTF7LWz8hzl1PM/bw2QJfFbxZMB3gYBlHtX0zbRGa0VQBcye2GtWgB9XSuTFf4PWhgND5
uThqFoLwn1B6ebTFTRfY1KH2jD+ZlXI/7dNTfM5rL0WLrW/gAP4ql2t1kIWc5NlveSqeR5OzSLXs
NGEpnlli/BJKQXdvDlGuvjRtmbKLlvqDPBCpI9Tf525pIUbDljjGqfLUUomCP+CTU1SJVRxffFto
hwjjip0lAl6SOmUj17cqCYglhfMLZdXcqu6ApPGUsF9zltUxTfyh2hBfzIBH/Tp3ZT/8OiYqLga2
YpZzC0wu79373iXn0v+x/R2TOTQQwCKYjpYyxZ2VmRQEeRrNUkUPQBH3QB3q6i4gbLMkzsw9Dx/o
1aFYDkF+3TgComOMjTRl8CfSmjiiowXt6zgXCroO4dQjyV2bup0nN+66/Sm3NkENsnAXqrRt2pvE
ChuGznun8lGP62Cz35lOuDopkCZbCgJgK6/Urqxd8hwpP/Y+Hzc4B37YTja02W/BWWlKyiH/FC+T
l6tUFyquI4pNnd3zyeA5/86qb1g+lSCKVGEiIPaqIuwOg6Xx6RV7+iu8038XnY67ka2fU9DJnrG0
N9n6diY0hMaCjq4Q5GoLxvToxyC/8AWS+NeI0nwcOz05M9dpZo2xIY8BqRQ30Bi6rTfwoXcfvkKF
O6Qx0VPLqWgw45/5e5HPt7Ov7/BwvQ8PFwDCyhzG9nWe7AMoVqKYHjGf/OgttcWjj65dE+2+5g7+
8bPLlRAFo9rROG+QyDZpbB1vN6iCbDCJXtMd7U9Sf0aBaO/4sBrfqpF0o6eOHMSn5wxfKyc3AJ2x
nEILvZJaJILzLKF1KlrrfOiqVABqIQg58epY+xjyyR7eBGVXksVIhrJzAhJPY0on33ag+L4dngqT
sE4EqxM7bTWylZx0IUy5ybL5UYKT8LzFc0cYPl9HIeijed5zGtWiMa6vY9KHduPiv/hNSxqVj7Ha
OuOTbqypTHVDzVV7WZVzojiHkcPDPpY+Vgl8DPj6GzWYrLZ+aQ3ZqFiOogglmhyNrAJXTPWkVYq6
xBdpSwLTlB1nPYiEgagdlmuZtSJ2dZAKrLoZWgI0BOrb4SmUlWw7HwtnIPs98wB9XWKiNZcC+X9N
y9ey51g1cY3eM58L9bNmo7l7GXDQH0JRm52ORtnvHbf5CHi1xEaUIoBHctsBGFbtUxQdyi79pWAI
zftJbNvLoBPE4UryzUOh2ZqSgOZ4Jh7lNIbBQ1zI3wKBc/AjrYsEtbRke7TDOqgkhxyWkHNLOI5M
NcpwsrZUO/xhYnvm+FTf/RIb7yfEFIeAgV9CcUTbdG/lZ2BPHRPipUOgeV3QTpZJa+pTZ8Mgg35I
oHqYYkzZ/nq1okqsFRPMZ+m868vHwVR/Im0a89ThSyBgQ027ycWGaV4dyKOdd7q3tCNp4pS2/Ouu
MurFro5zmQb2s6oc3219gJjhggTTGpN3GvO5gx5nCl4MvEYfrL1ozfnvByao2iRD9ZAV/ISin/MT
Z/JH+91+qR6+Q+FD4/nxvL0G24zsq603QwovT1Zdd1vOiscx6qkMpkW4MO2JexEKddDfxBngbuHX
pJB2hyeWb2G004Qd7hTv4JHO66tH0bj7bMcGGcyWmfwsjeDNFLsxRr4PKF9OENwrH9R18iAAKTAx
74ismZCfvBDpp5S9sLaljA4iDTBFMCt0oOLvHJnEfT54DMWvdUomHB6fArBaNxaHV9yzaMYND+9j
/RpDs2jd5ZSbhhU7N46IvlbDlTMy9KWRvVKWN0w2gEwbVB9YnRfWsz+IDUet3cWgoscQyHWZ0NUA
aXHpK5jfhKSqvQBN8yiH9DIVJKOT3QG+koxeHYPLae9ukidWuOLx1BdIhl//sv7Ji3o8wGG7M1+W
rtsc0y0BOhiLQkArRaMsQyd+S5+Ejblg2LbZ33pRFdLakQ0j+RTNbJEhwAARzjUEZl14n4vXvcjw
djHKTM0JCPeHRVgV96+Bv8Enqi0omjAzee6VoIy2qkTCaWw1QujHL4mShm58Zf+UfBE9Iq+JsxCt
SM2e1f8Ac5RcTlfgO2+UQhdvnR5A+ebopf162PsCJ02qNqG+nP3GcjZo1P1idG6oIekVUEb4NDGR
1u6oUzp90GRfcefGr/VUQtFZMIT62u8qlt/Hu09gTYm5TucEEd+oxvSDI7ouna1yjEg65xwgka5L
duU7I3+ieTbKdyqPyNmJ+AtCWhpUa4f014lZguGikwZlVElsai1QLqSr+WOUyeZkO0yPdzEmY1cC
QXv2tWpR80ZjqvlmrsLH09RDAxfC9Lks0uvDPUwVBo1qLgh2EFPjT6778hJ8AEZNpwzxS9OHS203
RS+usz1J8tj6MSGkva2KV3kLjCd/JqXcDg5JUYdVGx8timetB6X4bUIOf4RUZ4PjMwz51tTdJGY6
nPBRULLxziQhZdbuLAlfKiDg7dUX4DejeNPuBT/NNu5M6MREHHebHB98+PP9FH90c/FU6APDdnSA
4PLH9Qsla+UZMGP0Kbn4/G5Y/ltq7Fg5IBKskZAYUYhZYNg0tvo9NHdtiRbLtnubr5MyY2+bDjIw
frRdHentlZ41XZAJMRVvjRfOLCrqXYXyd6qFqtL8DkXmUJp5sYUHeqF7wEUCZMQvkYb49Uti8m7B
C/6xBZ/DF7Mhlp83TdPKbVaqOYjRL0T66rDgP12UTU4o3P1Ea3t5VMfWNJtEXhA7rZ3d+32aACSI
va0s7uMb/B0d+2UFz8ZI25jPJyJKvIF9yBNwsafEXU9kAPrjOieXH8OgYUNaZr+gDDC20w1viLGQ
VgTTgX3Ro9rSeM8kzzl75l8zZK4j/J3lV34i+o3C1NVSnu6XmeuWb6YOL2ySXeazzzgRf70nfWet
YYPpGCr6nswp8REY8jeMheGFpRYEDtBz6RBbilHC6Ea4giD77mxDFMM8L6lYpraGmWMpWCXpIRhb
LyjJJ7jKB9LCXMYriwr++JX3sbVAPKhLSnxW1K2vdVpNKkAGqrpMQRuut+Oxt8UC06fT5UgKtEN3
EE0PU3yD8KHIaQPRP2zSOvj74ot/sEuatasseiyK8L4FenzFrzVbIqGW19sq0ZJDlrWlhGNi+HQ5
vUhT7zSxXk8dtJOwE4C6FgLUx2wWNkK9Yk29TA2YV4uQCKuJ+YzZ/bIGSdleQD4OryyqSqA48Wih
LEbiP4WYeMaK2OkgRIeIKRUpx4pFYlAoy6OFRMgtOlJGiAiR58dNnrNiFFOG2nsyA47tDVzIRBer
zwLMbdYb6Ykh0xmHxagnyn6JZvD6EhEaiXQFYVsXGs9x/sMSfRqharX0GmrKrzTDHWU76EhGhDb3
9m6035GLGB8Wq3T7/4sOUcs26VS03UQCWJYAHQAkAF/9uPFVKhbySX/aZYRcNpNEvyJhpP0TKK5A
z8aWBLNEIjjwy1VIz/sE532fcAcJBEJOPEh/jGHBVA8bWfTg1b5sNdFVbrGAbFzduuWWQsfAO9nB
zQJjs8172JdIGB1iUwl0AO2Hu0yox/UODxQPFmQ6JoJc4kxs63lOkb6d0svYOXnQbJBlO1Z/xTNl
/Ry/GNngCSlxsBSTwal9mKj58eiVZ6sD46hAcfx7G8UKiKwQDpwaHN/mFKVOPxEIOp/FdNSE1XDj
yVnppCwwfhwxGpXek+upjKHsA49B5uh5xlzUaShxnaqVMfemeORtvKJPPJuV/Qx+4J0T65Opk0HY
zklh+u54WScyoie6Oa309lf0UC7o3b5PjdFZUgQAHOVRcSCh2PQTIWSbETEj0TXLv6pnMypxTHKv
5thH4vJs5bOKwILqQYNOzZTlWo9N3Z2xhqX+oKRLCTUgSSTh99xNeDiKmjP++p7+Ba3xkIu25Pai
MPJFbYHZrvni044ftEE8RcHHiO6OCpKsJlQlWxUogDwE0U66iiDadcrVTroxAGjIN1R0tE8QtNcv
Nv2HpN6TB5nOXpmav/xHZfCvLqwfLrX1Va6F+YspsvapWzrVKV7CBuUnbmHDxi2HTsWYxKtBDHgY
jEJQ56lBsc1c8z0Upm6Tg9/tD0tPjoMseTXwu3YQ4TJIj6rzFlPsyMuD2tc1JnQbC3gJcp4bISAp
raJ2lhgK3T/Gt1SDKFkG5l0sYWTNcCmE1Y5lavkerRe0vmRJkWfleS+CpO0sP5Iq29rIoikCNTjC
sy8z9Dl07HuIzIGlOYHuqgKMKeEY7HH8TaJx/5xxMc3wbpld8LbtdtO8UTAe+eOxe/C9YrbpKaJ2
i3Wd5NLeItM78pcWr4oCSEsYBgjAlVdDnrQKi60TgHyqSf5wiy7B9YxAlYLoLYwcsOGwxWKG/6Og
pTP5ZChMw0Xff+DaRXucei9gGclxA3e4KghHayEEwQDN0Q+VKL4c++WAZScfxYKzdVaAk5Kh6jaC
IT9TqXzixDLwFsY8KekAzcLaQoVTbon8LvZYNUBmulgaMNz8FrC6eWMfFsyVT5YMgQyU+6OvhM/g
bxTS9u7ruPx8/qzlwqvf07XSSQVtE7zOgqyLv4HYLkB1pbJDR2ySp5/Z4rqoLtFchTL5qoU6U2GL
tGWPZq6frhlUrNaEoghwteARHiM83mp1DuKHZJMJ7iaU71mjq3Ky/cHlM3e4LXhK7bSwZMfq8Sdu
vIEYvCOf23DT+PwjVB6DufXr3BCCG8JLMGSHIk1/ywDeyoJ9GRX4fYjB5P6k2ggoe8jyl0jgPVvJ
lrdxvU7F5g6BJiS/4P/Pr5O2Wyp8IsvC4pLeNYxKBbQuZ0mUp27QuTUMIhhFo7m5oLQ1PDj0NLhS
+L6uO9XWF9ULLtm5FEu3gMKPmVKOG+vaD7dFhJuvt/kPoXe92QnADv2acIt3DdPBDaWzOf4NGfys
UdrR0aFVRvZajRIORyA+btixjk2kAMHmmKejcs537cYtOTH8ExXrc0eKTOCYpVF26mbkOsv/pJD+
Ik5hxATZ05wlwmGxRLDzjQR7UZ8HK5RJwwOh+8E5K97bOQMrjsIhhkPMAagFs23g3j9LzTP9Zmv7
fEJC7lcy6EpucUHSdZm8adHYeIrWiowOKB4gYksOWUjVnzTmxEyn9z+9d0ngM3dqBkQRm6ujrmVd
RJ6tk/fd5BLpVdvnU0ldgqHTF3O4FWxNL17aNKEIuCbJcWnOybah29jlgLhBGSFNlcOCF870SCWj
yNg4RpMr7KCl3oNoLiD77NqkigORdzn2giX1DuzvJpwSvVNLv+Qcf5UCgHIQySPkQK6wx81BnPDl
f46A1Xb74S3n47tOSZXYCFi9k/AdapYyk/OjkVwks+Itw1DwGJzx7IC60wMqgjY2R6NvCbud+1wd
aIV6Mnb+HrsIw57EMATjt9tWV123rIzmjaBOVSUt3aQgEKX8ffwBWYQOP0m3rWZiNgq0OKam4JKd
ootbtPepTbX4fAWtCv2kjIZLq8nibduQnzZrNyt6fOqIVgNjgbUMc0DXBdeyCkMgew+T4hd3lNz6
JkQtxV+3Me9224B04Jn4jQg5Rl/c927gHftm3akT7bjtBASFkCN/KkPsR2nvHxAUCjai4JuyVvSM
qNueqSFVofydHknRN2XjPakShrHRjxSuSVyMzWk8yrlf2I3LhFmVVYSATbnTfDPl1A3UJcOMarTt
osuQPLIVe5jRwczdDfEnIKHrYalquEeVbGstYfNIchPtYvqkhau2S3k2Z9VW6Z19JKmkObQnNtdv
khCzCbSjuCT9ZnVXVKqMFcYl2RuAQOoApQhveNlxw0PoucjaLfv5Ct1DLQDveiLAzsQxQXqFpa2X
I6dQD15sJIJLKFDQE/CLSEIuEODCy2MAXYGTq16hhSt23DPUKlWvOgI6bceRuBMH8uGjGYpz10o1
AmqvzQPZQi2EsJS8Dfp+9LxeXgs4/b8KZ4wkQ6qUv+pKuz37Fb7P9lgR6vWGN4x64qEjHmvG+bkU
JVbfsrGxCOFsTJ8qVAqdKKZLP7u/xPJtKyv0qy/9Q7antWbrS8CMJ0v55K1Ey4VAGg2PA2lW6bPn
T8jO8Qu/yYG0kBfDXvpMDU0mM0a3Y64OOm8Hfv5Cpk3WacmvblAqEAeKIjHhn25Ij/fjkOQQjBy6
ANooROriNZWyv8P24iT/ilDfIm+0QvY4Qkqr3j1Hwee4QuFEhwN0u7N9Mld77WJFCsvSS74ft6gy
Li5Gg1NllAitVHoRP+SEuBboIWBfdMws88y/BRrRyrR6tJKvkjcqVl3l7q9iLmYAjm5QU7Mtrlud
1IhZ84Z5YuSicHBi/5nusTKotVpt4zBLX95YiRubhVVjRNk5QO3YbLtSioLlmluVwYGC2PVqflnU
GYZqtjmSPpvPyN9ywDmcqJu/LVusmG1ensu/oOGnqZ/S/i9eezL1ZSXiZh0Jq1Oa1wRkqI57n2rI
CRY57FWWXGR+1r4n4GltLvnbN4FXZ33VtFpRiJyBkGNKymFIFrqaP2NDSqDD3lSzZH5Xc0v4PYJX
x/uzyWsDdE7AA/ddO4KZUrlQxPcUJ87HTvkeUVyDctvhWZ4/xreXw6jD0Z034VfqHcD/ubhqXaB2
9MBf610YecXvc4AuXKaYk3k0H1OzIh6rGVl0lmgrPeXgngGlYsV2eSYWHqAkKG/xoc4JQke3nbl5
opTqyw0FQc3ZHrz6HPqQvW975ytL+yNOfYcaHLpptrTWEsuA3qbtfbvohhlW0O5c8ZGttXcYH+0n
fY4mIquFlJSQJYzLyqAA3xbXXo0iJoHlOzCg5U3DxqOdDlyl0z3ZaN6gbp/+UqheMgTKZIQLRLc5
vBVw414em0CbfLnKYW9Y+yPqoBMFna8pos0UcQSzmV/WLHWebTDgsDQOfgb+bNY9J/gnMI2yT6oh
Qdl3HaVKJd9I4YrD7tLZF7sn+/GvYaOLYm1pSyW2LqcP0eanZlXd2Se8VKKiKjbHbHoavMsl9I3w
kZiTm+XgbTknIrnKp7Ci+Sud3ACZox+7kkJSSzXN89+urz64jNLCp52hRzw6wlwZ0tlolygPCdIF
pC2/0IbH9yFnIOBG5wXv2OA8+xFJcvqwdr5IYsb/Rfqmo1VDAQXkWV1VZZ1XHGoBsSp0gVXo5uls
tr+zwx6Iw4gVPQ49nERwxsbY1S3wOIT4BYAcOC5mzcHDALGH1g6ofnBcDX3wmSbN8js45vOz/Jq+
i/e0bXszLc/wrhxVme4J2KOzQ6Tb4rb2gwgAXhdhiYeuPFDSOhWMuLKIzc/43R7Kbw94I/qy847H
4eVPpyjjBEmeYD/odq6DwWzbsxcbXLSZYKK/VrtGAaq9mB40/dgZanAm2KLOZiMwxYib8m3Zvw39
iq51buy06z8BwNge7A3kMQW4tE0hj7qfQKe+K9WTWV8EwfVTG2JvjOxUGqW9WpQKVG9aEzi8ZgXJ
iRTkHwy1iGHGU5YScQPZAhLFz7TDvDYAAO2hldi2XQOby2wDznFyys/+/2sTq9jIqb43jdVO7/TL
6eotHBRDSZzZX2KB8uB5Iy1srdQruQQSP8X5xruswSGcdWSI6N7A1VfyqjcwjmFQ06gk7paMJUKr
zmijAnYyj5WK/xjgIjVifbpMoJb7FzCc3/BZG2zKyLVWDHMbdQqR8rd4PF6zI9XL0O+NXYgT4e3y
jkbqwZNSIKZFVr277kKIyFb/gXd4zdgnAxEq7YA2RxWlZAJy4laiuk6cgVm8k9fNouXk0kyVlvr1
Wa6eJpLrvXYFBjZnRb72KjVviF2bPdfk3at9yH5mV8y8GNV6HE3iBlDhdVOMY55PQ+tyLzh3ZmK4
mZx21/BqBDoD3NRGvN0tIQ1Bm2ESo5FZ/h0zBMAaUJP0PpfChxQEK/6BjmUNQCXdUBbnAZe+e6De
vUJI2VDBjZuZxZZmbAja2f/4CEbrskC/CVKJEKyJCBdXoqro97kVbVlxutnyuFVcD6A4ZJuqrgz3
w1Ou+LedIbCCvAQ5SpdYhUggGr/7gaKl9W99gS7XDg8PAfx+ThQo60IiIAplKQx9nIm7RZ8nhMBa
NzhLHOwcp7A4B1NDaSSxSZ2znhmMcBb6hrGdUySvXTM7/yxCe7ePqlfDdhGYKq3Pk/QIV/Zvp+T8
9qrTXfkS0DaMdVHjLacvlk5wpf+Kw+DpONsJv/ZO71lceMKS1/F2ZphrGt0/1vQyDMSl+5CZqWRI
r8DWAV1WzTVVoNbILRoRl7v2XUezUFJXoyUq8pbn01kSMftT3bxDD9iC0G526AZ+ol/zilecYrbF
HiL4WQhT+6xYc8OvndmcQMqs5xI4F+I+iPxdjREh9RwWrxzvdcj78/R2z0VZOfarTgfrPhRp/Xlv
Dgen1lboM5jM5WLKQH+EQ7BJz+z+W84pFqWVDF7xR6s+vrxPob38CleezBZTiuLvHSiL8X6nmoyX
FJmEEETNeHBml8FFVG4nO3zO2FFLgJasYiYFgg9LhhkpzS8hJqp8DbVikbQ0EIhfRJq3nBQMuTWd
uuymAtEfHZczlM9ztW9awUqx4b3SDtP1vS/FFq72alVfEUOLYSCX8XE9XU5xjgp6dNg81JH0Z0Ur
3SDSAo1iQ0836E0f1JnyrR93Pw5ADg3tKtZPFyViJfTQA1Wuu/+WNwdKF8Oj6f7ykOqdWEIaZeO7
ecrnQBHjrEpaom7sNfQDnnd51qGF1M3RHHRl+kadv2vgOeS+RGYk/1sXFJJ8EeWMGvIVIbUOijGF
eChWr8Z0DZi7YYgAfeLQKseL0qCjbRzOK+7BT+vieoJ4t2p1U2y6lUt2TUmKogpoia9sxFmqYdGx
s1LhCn6rid+EFXXmjsSIV4YwuTNywFZCfPQJG31uD8dQ+Wr8thuudIXywh2TIQsjiQxLpMnV0KJU
TeEwqE/Lzn+2jRBs+D//Q4o0p+d8n4Q5XH1CQQks1eSVBQBlhSFop3Yq0s7l0+aroooixL2JfDlD
ZPJtkNqCAhz4FCse0AhrpmHtK/K541ShFKWScfIE+n9RCQ4kBNMjdTB77vY0PNeMDv3VPzXRSWQB
xbDA5yjfOUJw77fKgp5XbatWHLyhLpvWhII0noHQ/aMV6bDM1HW7Tveun/LpMvSFPNhjV3iGjv3X
nC2HDvAn4nicrZtb0yHxd4cmTcFcPHsx7AZe5wzdPzpMa9f9tVVIOS+mKlrT8xQfApijGaotLe8r
OyCDEPyAPV3zqT1fE4Ya9Ipg6AJ8/YlGz1tnMOh7/HMJZTjWrZAAeaoPaQH2qX2HWiZvy7eYn5VA
nhODNR57Y1TLPaFGnDsYsN/fi6iiEAELXcrOklmcm41XnXJiHQV58sjyzAy5hGyrJX2/stEXVxTY
DEslF6klT1m3nONM3m41s0IVPHqWBC7ebNeWOqNdwBJ2zHNRbQ5fwqh+XHOXbRERbvMsbRhfXc6f
vypOWF4VexUUpVC72V0UslF9irgUayHbP8KQmoc4FV/Eu6jXFW9MXg+xlzjWPmseq0WNe0fiYmBb
iOZENJylAAmbOosaRTopDyzUemh8wCBDZwAMDXcBL0jSUAgcGygGtwgizPlra5oVqInRt1hwXML3
MlrQDrveV17EsWTokHGVJ0RYi6/jMkxo/csC0cNvpqt2L2y1EfLOUeasl5Lm220lfHH7PPimGS1M
WTWtF2ONoNnDuWESPRfUWpg89eA8DwvJFga/arVl2gJu9pJQG7MW515sSkCeX8BXo+U5Db987HUX
UuQjt29b0MY5/wAohSiyAnIrMX7vm4fDf5PYNjUO3yXbtgDt15sRH1kgsRV9Hlm3jzsKv3VcV6h/
4OjekwZC4W8waEHWv5TrKZny3/9aDeqyUy5MooSyuUpXtx2C1pNthXvHvyRD0YQXbycPg++wp0Be
xKWtBwKVxJ9eLST+X61NVKmkEf3isEaYZbY/soTVTMf0UDyvEzKoE/PtBz67KFIYqtg5GDMT/ops
ydoQHmaBZgCRiCEYrejm6+0XwsMMXW5IJLgnmScV/RIgM43L6qoDkWsL/8tUSaoLu2pb+TLe53O9
dW+byvWp7oPApghp37lKb8zvjD025mN0DFkJwBU3sPS6VNYDeRWDCuBz0glM1HIFlOyxMstdM8Aj
gNmd3AhzfjadoPKmjR4WvTvHIorcW/mZ/ITH4nCiBDcDCPLFgpW83bSGeJV8h/wCaGfLlN2h4x4j
JT3z/DethNR3IsT/Tcv25libNrjJQGQV4m441p0ZoWswlBuFQWo0YGyaZGAGGvwMufZPtzPwLlf7
YLW3yHUIVNV58y+l2sG1CnPLwqoag1CYuKHXvUXQx83hFhlq/2s43lmz5pkXUuyKOiALQlqeXOv9
UHOUnMLnugvRO80rsH7NFOm9WmPL1G4o5v2rMcitYm1K+IAcuXIee2xYj/ta9wR/NaP6qzLxTlBX
HhdFN+826w4Ya5ILULLHl9HZ9e5D+YTW/kWYxdah1f0JvAXS6T51nM6wRJwqg7wdDq4qZn1Gbznb
VrDXyyzugGU9/M4sGv6gnyl0jZtzs4wVKOa+bAUm8yDAQ2Bwms6SvrA+DvYKIJWCySwDOUZlP1sz
PYN6D0guBLdjW1pNSxZikChVjcuVpoWPEY5pgibAg5xvZWC5s6H4STxm6N+CelRfHo2tMNT8Zps/
S5/kPr8AlnFYbn1leTHBUHe7uqiWXJe47prz0qkuJTl8Q7QXo24DPHXI3CpFGR7NT1znlTrCaM0X
fGHSd99pZwZ0z/phNC50iiSOgx3OuyFkOBcwaXvOpB6FFluxqlp5Wth1+08B6I/+Ar1LnAbeseT0
mB7WC7Rl77SFeqjBLf3uiPgIcntpzjYfuvhPJSu2QVMYl7UNjVLgZKemfQk/ZCqiqN5QzFsEH8wa
rhFjCBW0EswxUmIOJuLDMYvSIXUhmzV5D4QRk9WLUAARqcrGNDv44bBDzBHvyKWy6fafZVKXwAXE
ckAIXyBl4vvdQ6s19Z7QRirRAv3YuMG+TgrOUr+DKZ1LhMo7lzjYHBpAVW3P3WzgjKo4zs7EZf8v
jZQ3utBKBrTeTHGFjTP3u4XzJ7eh6t3nMclkvgTsEskzNdFP3iMlVT5Df9vTFOe8P1eOVDX5lNIP
rqbKxLMxNG5aFVUeJSPxbJ/7jVNxUE4TpEqk5bxEGQOb8WIEvIqnYRv182qnz1J5CFYCiP4vNkdl
5xsKjVWoHnl5A0wndM7PzzNy5hoTOQVObMWqDRo5Wjn0M2ZIrQu8NFPBxADoPbHlvyJWJu2dCzwV
cDLFEipWbN5lYcG4D6wUYbCMcoKFtv6CkSIXIqxIFWNJouO8AagQxvk9NsASKR2TRwP3Fo4I/u5W
tY92WztFolShD6fUQsH1FxzdrgBlH+vQv4kl/Hd9G0LkbubeD+HpwwMjPVBPSeD88Nc/Snp3+1Nj
BpIVbQMe5O2Fo5wI6HDMv6PUvTd7R8Z8qIfgD1y3T2hdDyhZa65Mr+7ago3m8rpbhQPukJ84DJE8
KeBTT0F+5KmVabEZmpOKmxyCWVzvt1jiSF/ypVFaw+Zl62gDX0j79eCbRV9XuhtiGbSyKzCJrN9p
qsP+0pBoWr39lU4lncliSYry5DQk5Odh41Kv823Za2XwHv6hKCGQOg0V8xcc1XNeiCly8vgrUx1n
xVeNTGwuIW+D4ORJctiL1M9R66LabRs0ke329sraoktfabC4aCkTJeKMtNcXoy8EVmGtj/mfDl0C
3vffnqVb0hWS+lYL6kAzRuvuD7Oi7ld6WlqkwTd0St4agM78L/8qNKwDU8Q/rrzRR71Nr50+94ZA
umHKn2TDkOLADk2PCLgN4BY0uctRJrUhwO46r0qRDTZ83xa95lwOWnl2u81n07e69cH7dxf+6zZ3
jo6RVxLokGcEKA/hkodfMfG3P2cDb2rjbh8ndMZqXF57MYQPZL96OdB1J8XTCghcLqxGcr2Y/Arb
ypDpyCsBbr3T5yuvh/vg7D33RxeHIU6jmeA+oqcTppJmYAfSTX6TOxIjcpwK11/SVlB2hZnPi9GN
Gm0GbPy5gpsaG5V7RSsXIgIUb84imSlDGldZzbazrOwaJ6vfOTNFhESrg8OsQyyovFSj4/cYmvXN
1bUbsavoYrIJB2z7uUyiKqkeHeixt78INFL/slD8nePVATG80NROZhQaidzlP3FBWkI/vG55JNcm
TS9EzD7RSZVZDijG0ajuj8Nocc//S96O5sgaPirEqe7Jznr/uUoES95aXYvUHQrFWY0/8AoFXmAc
a1coLf5b06GvCng5PWvvx1Hcg3lnIOYzkkfg1U1h42igUhu0TfAg+vIFwjQGOUSvWyhwWkugJPvb
BNgl/pG2jIsOUxBj07waPBtfV5gtdP/7pGgziOtur91BdoW3m09hwj76kh6lVVp3NbpmXUY6ZtQm
S+uoG+XhZ1FFDsyeo082QpaQQUMRS/DB8zm7yBe4vT5JKeLM/sC/trvDy+fDDLudC4zWuUeVf+DK
oSP7PfplSR+48wsKuS3Xtzx4SlAnAiVgQBPxgzPBy3s7VtHWidoy71hKC1H9a7efrOPIM6fLkj/H
T6G+L9XTXFD13Cku/ISOIJi4aHFslSYHFdNTBWsZ417e4+mj8zQGGmW8Tz3HkuurrSW5L14VUjbm
vwfLjLLSbGrEf8AVO7Ik7LbYJ0ZO0lSTA+IAORDHJM25ZqenQk7cXJWyaHDhFOz1VC3n9WBikOoJ
QFxmi05EYLZJsIXpENXG80R+s10CCZ37vhz5/WWrYMkLkNcqKvWtVhWILOUKznPvtW+Pm72TzqH/
u3tiep8+Zip5imCPelpJE2i+4QFgipq1Lw+cQYKATXCZW+e3Exgy+pdfRidtjts5xBz8My+O87I2
YI+Gyc8i86G7pkC/smcIBsJVROPd4VmXNSWIlIiRQJ5upG4y3C6rgCqk6WodRUMc6vaBlKCH3AIF
jrxEfUJ9vUFat1hGp5/ARLMpfSGa0WaJNUhc6LOGmk8aZZitWDvXrudXegvqBk8st9zL16i0WuEw
KbT6cnR9GBF79Sl4qr1pvEVgglfMyN2oQLKVN3QDQDeYBba+aiitn0ox1z+8okj72RRthQfNNwN6
lgLDwsfMAcwpyOR+M2YmITjxiSdXKFZ4xUL6vwvxduOrOWZt9FcBlUMXL17MGKyhvl9LgqqfmcGR
T5CZhM1L6pRW7SQ9jiVcehaV9iJoK6h5SfYicVC/X3OJJIMHQQQBJ9HQGJCkz0OVbbFbmU5oY8o1
F41UoQDd91QAI4RbxaO4Wp9LWky39kOasxhD4z+wCPztU9M0t4fjaKPjIrEzdyz+huo8dmprrkHY
C2PEkvRw8dJ5UzLp6pNybOZb2lcyipi6Eb8nX8K90wb/JWs+y08gZHyIY0dYgH3OCIs1bmQYl2za
uGq5lNI5orDuyFp6IPg9Wnd9xAMb8Xa2wPOMJeKycBy/HpN5GwTNdcxsPJPFsombjKRns2T6wulj
Ulj1pPYm/2DWrSD6utDxQSWrRcfMhN6d6h+UY/FRZx8XV+FQY2MxLp8bWQRYfBDThOOppIz5AQ48
vNXzSwQIKEoiHk3Toc/Kt4kBUh7zUbygGTe3xX56mcNwcZS5xJZRZFVmYin23P5Om8JRRq9rIPTZ
xJssqKwBxr+a7Ik7FlFtXb339FnPuBN4OlZknG+CUjbhgk5h08h871U03ecUwmS9EO1WBZtbPlc7
kiDxOtdIqO0cLVCeIAbRKt73OTtlKd7AKvoBFr3DFj5xJC5WULcmrnGoW7pgbLgVL6lLZPVtMJ0Q
R/49iXeQ9gDQABEkVNyYF7n/JYmqo1DJfgU4eEQLDihfUrq9WlocztbKpfJPDor0/8avdy6Ra/tt
AEHotiXO3L//YXsx3GBAt4tCKUgkkCJ3pmLrY0vskYdSJvka+s93Ulg0GRFH35Vk2rUe8DKzOviU
Ir6W9sV0uAEUMkuwH79EEn6TLHOu6D/eQVW+ONJxkFu1hp8eC67T1bu9xfinkiFFbGUO5S3QpQ7T
nL9B+UDRuhaFkZb4EpaaJbvgVIiuCYUf6GjmDXCd0mMHmOQzj6cEhgFNRrru6KebcPzA4HxQJSTh
Q8kENwMn3scBrTreyDltoYqrzxTX/n7JqkjJjB8WmCeWFLdNeM1gIhyzaalxZh4mleDcqgYqlTm6
D2absdFShnLQ+pJ72Kuu885jGvvx8AsU2fGFWxkrG8GKdQyfRGgPH1mViNbqMvKdoWzLBBtyk1Pp
x3J59N2IAAiWxcU+KKB+PA80hcemX7u6NFZJZMR4gFxyfhKlPlz5WezRxzhZSBdjv7YGNC68i8SJ
DZUVL3P61WVm0UqsVXbd8sLe2cO4jrX+Nd0KlqeJ7UmWPTGJfcC+9gYaylcnYX1zIbZDkGcsgDvc
VHNXWiFIMyD9acQOanj0kvh/TgpJXD/3Xv1miBLYO5LD5RjXOMV6v/fIFH8Df0reQhihrigreIY2
2EJtcnpev8mGlk39x4RuRkZZIUR9a+wYIp2XHpMafhRHGWEynQIt9PuR4sLaursp3tAD+16flswD
HJ0iu1/Cwj2aVpei6/QysD6Rjs4wS7i+Ac/zxvnqNhqZB2zxShBSXRgEcAGm++gCRvgN9szIjJIL
SGl7JgKQpq9iJweJ32Ldg0HYpXzSS4ViFr1iEIHGbFWuizMCyTWolVC53SBbVJhv4Vsumlo53jMa
zyVqaMYbmykwFyN/EQ6Hg4pfivItKaxBFSSamLYbvG65ZJg8nOvmMIUr3rgWdW+Ihl5/tUCHOXzM
b/yLC8Fa6BFA6TaOtnDQDbS/eHXTKlWbuKuGFDTAVydiN2VLYdGMqOF0SS7C1zkmHHoPH3jVoCeY
arD4becJmfUXItf+NlYtCOUe/G5KeSMnktAZomDCTJUsC+Ii1L70+dKL0k/3+ubwZky+Wzv7us0q
TEwvqK8YAL/ee2jnNysywlk32fBGoKM7yisdrL0VKCNzSvAtrF+7Wc88KXW8/skzOniFh9Vo+fWB
jc/AJ+BEO6yaM5uKZ79ASnfM2AaBP37pl0yjS3n/vYrWJ5unSbPK3g7xoBaxb8Aax44We9Q2JVwI
w7iKRuBG7J+mmdr3nGGvz4VE5+Pi0oHWzaCtChBv1DQeZJ64+F/CUQE5NBuJSrRksaEAMFVpPgcz
kReDeQccj+UoDA6RjOjiJYwClRSmQChFCGnHh12giqWNrmuRv9m5m6DcvCrm0esMaJfmLp9uoLeX
nZEBsk1XRrjkCz7u3lEh6eNVsItk8FHNb74fadkKNKqnqvkXvv3LYanJBDHdFgnPG2xfu8qgxCJa
yTUgYaa6OVqwCmPLwWB85n0WI2pnBkKEjpwtoCaznrEXAAWJq3UlUtfvzpg7/i9skW4A3CPXuHE9
9kmMOoTGi3I+UvLnEf51GpXJPWMZEbSahV6eZMhbB1Yp/G+TXzZL38hEpfcKUNSzppA7/RSEizjB
BoUu2qTL6tuid8rhD7tqu17KSza52RvCsjGBCHusvC4XA3GPPTDGPFEY14jzQos1L2lgcoLx+2yO
Q4qIRc+WhKUa0H1/sxCKtlOpccc+qqLDXz2QDdXwBcCxNsbVZMVVbyYeUORDATOttFYPCVc+B/aH
3uSxoKbHZbUj/RxCh97n2JKAWvII9na7dwatIzC1bnw4uRdpp5hLIHuli3Nl8OyBcO5YGtUWeFpS
G+9CUQT+JODeuQwrNZMT2kTK1u0gYnubSp/TAfNjOow7LQOxxZQSUXoxEWxdmnMHA5uWgguNzzdI
xC8fsum+QLv0knC8M8pNAGwrHqPSmGldPh+hK0R8bUrNKm6lbLFv15danY3F0D51sXmIbhJLWCnJ
jPf+xv/kfWB3cOdrXBCsg/H0IXVohbYh6O0U0ceez+JqqJpsy4qWFcYz4qh758lYG1pCYZCFCMcz
IA+VWXPDtH84re9OftNndBL4SZQZDOZzStVBhSKrMdmBC24pf0ia71XqckPySShGAmEZ9E7aqQ0m
MD9wpNnI1y5qKZPVBcvdEggGjQ/FaJ76oq7BdUPcPg19Z7KQ7y7q/TTR4+Yg1/bDkdHGL3jr4k7P
/OpEu+hKnaNWPo7qdZp0OmihkP+y4Ig77TkEerwbTLaFqswjTYP3KD+u/LqrqsVISZTrUExNRgOl
zktKI3aE0SABsu4b8UhKls10If0oUSkod1nuMXxZXsgH6Q1L7Zi2PbFcXA9bmmNhf9L1G17DcB3t
6ILFMxc/hkm0Bh1kYLiy+1sicx1zVgj8GTwpBO162OJ0mZgiSzzdq4DSdcPe3V3nlpbwCLpdB8uA
TGjAmoDTgxErd5+KtWU+SeTvsKn1+ldZf7ZI9wUDvUNUEV3o2zz53hJKt+pdxBeFAR0buPoaYGdm
1gWPQA6+E+6EZbduyZklAzd1T9L/o7r89ZElmsEzgjrqTVK5s+1Bu2CJvchFpxxCeBAK7f0Uu2PT
6BqEH3xpyDa+9WjnGaDPpRLfz4kwYl8lBBWwTCVQmH8w50AC1SmRJGT6AmhtAfwYtxpG+fq6zDny
+qsIM4gwMNffOy4nokDQHNSfZIvX1OUZagKd43cZVV/hgKDm5SFvfcj1sUHvlXZOizUVrMupPVvH
W7hU1rPf2g95r2vvK6O0yYN77bbOCCA59mE3Rpcmiu0Tclh1Jx3MBAH7juUmdLsqFsFSonz5t38j
R4+oCFfbksEo40Y1zN81o1fQqoRNmE0hiPEyKJsPHbQnWVLDSPzBnprwRkkIZDoSLAQJy5vX8HA7
VaipXlZsaffl0SDvs2dbn8SQZS+7N0Idj/GuU3+QPdRTj46k+c/ThND/P+7TEdzwnSn7TLW0T+R6
ZZkqc/qBKqC4YsHAG+C7a3CgXpKs02uu50aVu8zwV3KIULsvi4wuh+K8SvITaPtpIIHJ9s3Zc0N3
p3P2GEJGjWZ5GzqrGNKaEBiAdg9mXKWtl53/08VhGONnk1VuYVZj24UOc/CZAoUXVMs38buDwwo8
SGh6dkyDqJN14fv6lCjNF+WlBUOt655fF3WyepCdHUeOZxuloFy8nNsrDTVVS3BRLHtdjHPvIiOe
O1ECUkqaXtqHwVBJEe9EWEOd4IlyksDeiLKgWgO3uJMPKtXMz2zfrEL/apd4Nm5ofFMyBtIHTIyl
tKoo65na2eV3MrRkFhf7aiCbWf0/VjyI5QQfgbsnifdMmR5y4cVsDhSvLCEiND5sFIj1sWe8IyRf
NcqwVZVDJMrUVLLHtKlfPG32WTv56bUxkaGaAj9hiePPFjmjzPZJkb/b3ZcVgvL6i96oFemags7+
mpcnispA2tXohzCkkxgjG/hwEtOWO6de/DleYU7qOkN0QD2MsfUMDlFMwncojIIHmvBMS6C6bmrL
tjmbgIm/gtHHGqWvhF+uN8ZAUg+oLqbkioE1F3ZkhedzYZ/V3l4JLFlNLsQDHSPyVWbvjwrUqjrR
d2c4hMPJsXFJL3mx2ajxZlyeX3K5QRBS1wts8o56X6WzeTTFHu/SJl4FsmXY1Yc2GQKiQEC6pkrm
gjc5VnR9vdwIMQchI2VnDgxgZHody7kz08B/0EwTSJSZa/Y0h9uMF+OAlta8EtyJxjdxlb9F2kXk
b5ouQhyBwYH4Jp69Hwm3RYu3L7ur90pSxlVQ7KfK/pddv9gNBXfJNYl9EvPPgcePfVmfgibpr8uP
ykaxxNreieqOsyn2qzTyyCsmXCjDq77c7VaCX+WuYN8mLc18ZQm+inu4e7Jb4jEj5/Wix7cDe/V2
dzViNnKE0oQqfkyOkfcVsKvB3tiweZaVksn6vV9u5ODYkCM+FSnawk/xg5Eqsme4fG1SKFMCwR3T
DU0gWmAnZ1Kv6exvOCqDdqrUmS095bpAn0tOSoNJQ4lU9hW5pmeff4MjjLLeyVGFGuXldO5mTevX
vDdVmmMmQWzX5eTMNd6OqEaNjcExYacxd6bQ8KHs9VtlJrYzAq2o9nd8LlOufnczBwfQDTKWwWyN
F7u+CjAxfBu5sJGRvXd/7A5YSfJ6E3KXTpMKid5Xmq/UZFpluhDIdkip7WjB2OKOt7mWToBTv6TU
nrXqepTKsjLGetrY3PfQ6bM7KvpPQmjjKXrFKhCMXijgprFiI+Owda4W8zqvOrwMOVFreR85tjab
XyYPn+rgcd93e0qL5dKBYvlQhxjeOAHq2AtlURveoJtwp3+u0DDWGnS0lHewqnh+qW9Nbwa1VaUb
POxeATAiNnSLGJPwLhYLz1qY58oH+3pZqspvWACQMmUqZjdVFEeR9qZ33dq24cvtoiKJ72gGU67v
45OK/AWKBD7wy+31e5+DgsDLl2ernL6u/QpgogfjA489dbTvBNCjT/calHIMXWv+QrZ+bSeB5MrR
1GEkO2SS/8mFw/+aeFjlYTepZHsI3DBWL0ZQLoB/d+Hno2XOZSCAjokNFGAYMMGX89q7JC9lE6xw
NQmMXtNqkdj36pHW+h3nAPIEWYw5ZpmE7cgGXN81eonyGa45lD4lBkEbJd1sc26Qk2CawIfwXmhS
bh1owggF1zVVdjnp/GyrW5yVvsQLU2kQ0jflprLGYz3hKLwEHRlJWP2A6m/NMOzeHKhVI4IX4dI5
54tOuxhiuDNAGDBYJCpXi1SYpVhEz50J/B8Ta0HswPtkPR3wpV334ZE2y6k89vVZiXbZ8R4qD0+t
xEmIBM9coxZyf4LZeHXuRz6DO/qwzcLuyxf24uAZsvmNaqTvVpfFiH1YLsRGpM2jvxMVhUSWnLdR
N/bcS4zsj2eC6LNkW8Zm/T3w6nVcOt2c2fSmlW7ljFN35EVtYAVgQh7iDZy4S/AmoYpYFrU77YI4
nBguRjYR4yVxxR9hLbzwdCwKKfDBtElZUPgCEceVDpQ8feHdi3fIyJZ/fmDsoVedfJtiW70TkaRg
dvoqssdtoNII1dnTay6sdU24hmYusvSdmqNXkoMgBLbrQFe117FykHnarNoTsLKCEakBKgBSJFUJ
x1dygma4V2pQ3kTvYz8+cZJTfOCDAZODRLNVBdA/isv2ofx5UK/v9ka7I/UtBgib9q6SdHFoCOc1
e/ijMB2gBbPqv4sonIVu46eAG2Qq3O8dKU8PT/3xYu24FAEpGXx3ImO51IbEKLnA/ovFZjGAb29a
vCxJZnijMz8BrKwp/mYO9RH8tAQaU6qHltKYZva/qTE0kOKZh63PdegLuqBeirdv1XukYz98v4La
266rlWF5AiPC4c3SEoOjkBUJjzbIdvpwRJmDe8pzm9InXuBI8kGZbyeC2oQBomb4ima3gLS+qpqm
uJYVGfUvi900flo/+uZuzGy+Wu7xDYoP4VGUKsIZltSiX93UmrbntrkifcFjXKzgA8BbnWGRoRdK
I0Gl6CWuej+V+ZXw03LNbb0ePGCQIKd7zhGEAMFKJsiqape8T2QnTOLLImP8VlkBoy/d2ZYr0WgP
Fp96AMxQZi0dNwvl71XsoxrawTIHdnw9eGBlaaKveCLngg47a+ocnSbLtF6M9MSwTEl0CqxxAyt4
ZkYpe9YYOwqC3Q5PPH5w/U8caJDtaOkTmDhRDsldnHMqaUONWg8oxWzGeXJMo5sEm+wVuujLUosu
W2HtnJRNwdIADxefKRLTM7kpvh1mip86SWN83sCh253WB/ytCGJrq1+P5XZiaSuUC7xxLKkZMkF5
yIgankKXDgTeZSTsIke/t3bPA957j2OM967sTnUPHz94HHGxk46tcy4w1YeCu2TeqF6QF9MsGA5f
vgx8o97t2IqjT27k4juQN6WL9oET8mKePXo2gb0+r0xrw/IQ14DdOzVRNEYJ2iq9ih4udy8BXQyf
B0v3zwUJVj8/8WY4KOIs3WNTYWq8y5/oC+JWacIPFIIKlSubjM7PODrBbdyxHZZ2yyVyfj0ouG+f
/XGVouSqf4Lk6Yg19nMjtX5wY0xuoFKEyNTfWafNAEeLMjgJpKLpztgyLUZtHbn2rFdgWjp3G68f
YvAM73O62iAHMdXfENsqN5oLvCnBPmv6nwyiEt/XAH8pNJv1bFASqJQJm0CKEeqCM8DS0ztxbun/
9UNR7imftbF+VvjbH+n8eIwn6soSigoF1plqFCQFtSApXVZCa3oivYTFrF+5/C1M2XArTKmp9cFo
JB7UrdD1emilwnR+UASGh0vA8xf3LyPhq+SF/sSu7WUTIhbtgQuwMa0Ikm/GOa3xioCj0roQ6ECU
WkCYcfAT2+dbqAnOe8YRnfDQDNHnvECD4klZmfyvsPEqerCzhlDW1FaFlNQJjLaeqdNmJh2HD3BF
mRlJWmIg5pb4Y7mInv1QbhaRSrm1Pn5btWTGzpT2ae0Cj9HyRQAF7v8tTLDvdyU4wGIrXuUkprp9
Wfa604niNLFc3+a8N2RTGieXDLGHXqMNu8IhsJWMZQdYNm+5+GTDtniHVIRXKvBtCUUSfriiV3bk
swfkpbouj4YBiAizAvXu9ZyAOAZLyS6MslS28RVyXUjq6Cat8baJxEJYgWPM6XVBB4HntvYZA7Bl
k+B2JZkZ5AMbKiclg3jH0ZYmEfWNYLR/7I9UmicxdIa9+pi91z/8rqYWxWt7vbEjxiMPtetd7SXA
52P4Zf5ZMTYOdNHzWr7gd4Hbvabi6fhR2RemKwlmUzYR2MW9TVMyx1FH62hyQZ0q1vfJnvcVJzzE
WcSsf68vOVt1VbSc9KLx7pY78K0cHj1rSqkWyskPMm7Amx7IS6h6kZUKNsDR/Ruig/tp6PeEBjN1
H6jW3loVCXG1rQd4SI6GLeqVd8eKLaZHub92/d2GKsOjlUU8yKhq/ZjyLE8z6du791FEmSTygN/s
001P3owQ+zyArS6H4838XCtNK0bf0osRSGEvBjPHVaFo+BLEx5aKSrOro2H/cnwVbztY7HSLe8vd
XfdnXkmoUaOKoXBcCBu2lxvKNdZKMqQsP/C+H91KTLcBXrNrM3UGM8UUWZ4GVm4YWd5OLocDYpWY
qBPJ2X5MFG60d0OT/rBLqmXgkY5+0F/vSq3QgXINtngJi55p7ZVH7Va4edYBGZcLlH5l54nW10/P
QrFZFjukC0j7HnKd9AQkjFWuPl1D5wTReoZ8v8uba26KLmQtt4gRMlVwTHn25MFngJ7BfDa9fgu7
35E8GZA69ubOAF0Sm2IsAvSgJ3iJRbgb+XOp8pKiXpq+T3Lz0ESmQwgtObiBTD4rcw7GvZ/pNIEw
8jIgdP+vbw2nfgTQuyc7ZT2xpxzSJMz9w9cLtpBCWDV++9/9M6vFmiKOBufXavW+Dh22SMvcAl3h
X6rG9RQK7ZfVlxL6QFMaQxQRCq0vVmBW88kd4FhjMvqLAzuZDSH3o2xZxZpJN3VJ7TIIFVUDcWII
VYStgFcraY+1Ir1szUrDjdUafBzEPeGBhmKuP2HCcwJvQbqPwOxJvepR2yOyLQJJKRZpFheG5C8Q
F/QtYBfTAIKkJe/QllvoNgUisokqNAkFOPYc4e91qIfb9FJGisg/aPPnhVf0Y+tokZaVXr1VrBXL
QbgoPj+gfmlOjk5lci8AOK9aVyeJZkSbwooX0/8aGGc93IgyHrRDQPizXpC8WZtoHkv8xigzU15F
nJ8sQOLhOy0CaiTAiamL0vKfR7FrVNAwlj2ZUAOm04IU5lhvJKsOPo3COo0OJuM1GxFbanN5qMwH
KWrVsP4RaqUALkvmNK0WgmOfo0ZTudnfFSa2XD9YqtYogiFpjRUtXSUiLCRZa/6SKjcy+OmxraL6
h6xzJlAdlAYGd2Ikib2WF66il0aa6mkQ4s4YyAGCz45Hv4ExU4oVBA39mGot3P378oCn83qCARU5
G56mUlbHc+2s/l1Wdo/DGLtCO/IymG8e/g5cUmmjcTBYISHUui52ofbbVbM8y2kTsKZmb7rUOyZd
W7dFCbnA1glU/PrA9EMgpyzI0kJe5dDmL6is3kyimcbBdAArhX7Z8QvPevY1wiWyBWpmBYfEhGdz
jBw4/STiDdCwfh7IRYVENbAceJAUeHtdiM7ZHzDm1DU++K2VY1v7fw9TJBkPBuOlgsQwvNpsBeE6
IyHdGebNoK2Wj1cbk12nuuK4DDpSaatXEaV3o7wa8ClRhAsoIx0zsk0TztsQ9vVmSAgb121dgS7W
zxfRexdkWlRmmUUDvbm0zvvn2qrU7dxq8FnT/0JTkeS0riJX+Zv1xI/kCCUhY25Zf3Wxcv8ckpUD
OktcLv3f3w2Qqy4G1AecvrkYF1A3nFgWr7lq9VZlmyknQbKwPonlrjqBg2UOAgS/8vEFZ3SjIxZw
O35WJK7LNE/LSexCPSD/qex3nwuZ6g/2bz9+oNaykLxkOpizO9goyk2QoxAUAy5mbG5eJOD/HqhE
KTQIYv3CvSZh5QMFhLYj/DGJv79GQ+GRGYd2Lw+cnNrnAb6OLALVEdyRwWyR0KJ2yn39/jvD9Yy8
k6/qQnzd+57HlM1n1SPkbBc3KdGlZfIL3gWQD6gsKv+xJqC5HiJabvFMHbuNOugUTpz40LiWkTaI
G9c7UpO0NjGUyvreipJTpoAvzqe3R6tfrb531qsb6vX9aLjtQC5QZz6pCC+C12Qzrc8UcdD2BD9v
ru4d0WHaf2c84jziKDNRAxHM6e9aa6oOvxSgL7Z7NcM/flh2jZenFhmHpZ+/daKrX5HIw6b/EbIw
FU0bO6TT5LR+SkkGbwhFOb1DZ5xGg16bNulm0K7YwxN1NvCaLG7/jucIa9ciTIKL3VQtyBvN6Uo9
JEjI+xZoOAbDUgElnnmLn0e0bssukdAJVH5zESBuEonhxiYgNmv/Bt6I1dcQ54iB2wZoXhxxqeLA
QtKFMAK50ntq6jmlTDsG57KWxIsMJefZHm1f1d2e6KFiO/g1HTSYsYoKaByENozb59TOaPk6S8VT
plKfE0pte+sKdlNoEZYjJDYEqHo0ejbWX6MbBWjjZdRxx2tEpd7u7MoCe/rq5RHeWm5To2BYHxUz
8WXTxYDBwELUkxaRCVm0p2QhBJDFwvS8f0w2isKcLAo7WZ3YtWw1gc8V6H4XVKZnBGVnNAd2+Pd8
GTySmJ9N2zPul94eHzX7wu/87oPiIaSSUfwayIsAFSfEJX+uE5QeNBuCyDGL/Ikk0CdhkJVbZ9E5
oT35vWHWomRPLneobouO0wbKNvW8jX8P49ZMCnjFn4bfTN0ul35dqfMB3Da6FGrEUi9kC7ND+Kqh
5gD7hVjdHLQQRZewbe/cwXhl4SOkKeghNYA462rpyJWVyyYUNdq7c+lDZid/VIUTOjATXs7uT6yI
lD9BNDBrmIew+a60HlC71pkVzyav46JDDpBzoAtPlKejCIT16Ica/7Dt6C93M3esZ9Xe0wb6/3nY
jjOJx2h4OA1oqBl9NUFMt7kiM53GGgGsi2Gh7xRmeFNHi9Xa29zhJka/Rfru8pJLOKoF0PfN9vxj
+qjtZzsLA5q7zwzicfN+1OuKsYiBS/voD5+Vye5elX7ms4y4BAhfnWLdV4VZRyIiXpUzQIQcNAdo
X2wbRjVA3wm9Xbw7q1oLNTt2D+2Ag2sQ5YD16rImsEMPduBlbElfY0h1lJOV7l2UjTYhndwR1JRK
scGuqMOJxhTxRwSad9E3CJTgBEhdKQdUeah9vy/hMM19NENg0XvFOJrbaeLoexEILhSSmI+E16bi
mt/BzqtRcnY6oFMMguT9UjOlDvjF/s8CY7WiTVYe8dorySfYmmGvpmt6Ll8oAEjvIgBTGSODZ1My
2K/qnL2GtKaeWC6+A6PHimDSkukXXD6Vvqg0bLmlkO3wF3ilmrIJFmkyMVzEdT0nLbxqkEUQExje
x8F2TEXojHMl8O+0iYvdJ3a3Mr7fkt9cFQ/nPAtCKCamiC6jq9bTXJ2CyTt1M8gGGSlSvPLs190l
t4Rv6v0Y+H6s5ABCkKp4R1IZtznwH7OhY81RmHqRZyxNflJQp0fXpwIvC00zyPGgkHnhGPR33ayp
y1CD8WtU3/E1k4v3J1yHFUnEsF0hG4NQXhE4CWhh58SzXjPbkMDDQBAhRB/KBzCQnjFoO4GJmHxB
wVaNIZC2MkTSgt2iV7XwPVILgfrbTILN2D/8xp8rlSg3swKIeMtpZcXsNUbV0M3AvcshSXlikFSE
EIXRe2eOGRALBjbadEa8jpJI7xaGM7bL0dXmMd7q1YfzGbe+2TPgVqz6X8beLOrXYA0a2GEE2CKa
D7BR0rxIByERp/OQw4XDzbVzgHscFi/mPPXv033tKmQfTs/1BDEbXziUrnMFcyxVcUx01FtAGjry
O9SEDoWgjaOlILwkgxiILk5pC1hp8EmoOtFzRGQfkZR0J6PT4rP20NtjiAfp5VgtX55UtrUP++ZB
k7FhPt+RYXEFrdpirdEADebf1zQT6UflZ0uTIdbL8rCIVGFSq9sSkG6pWZZPoktWvrETk2c5Rxga
BbihbGEMjMv/KdsmaCLhlkHOdsRNkXDvWkxTstJ4SLifjnZ0+f8BkjS7gmaQLCeIP6Ehw2HbS/Rw
wDdDo7qcdXdB9SOONfbRRG6H4QNObsodZ0q8lnFXSkx27NHAcDlN0oOY7JaJYS4qSvhnlf+Eyqtr
SgaxCzVkEunYqzZsgaOGG9BjdgBFp3VKaCCo6b4tb5RaSG9/3zijgaomjMpFIn/nqC7JFFfVdNVI
qFSIbutW2Hl42ystTgzP5DlwudII78UKjQO1zPlhH930UbRTYgWT/wKfndW9tNfJkDX82uzcSRmG
M5QlgRKWg8MZkFyjr+Cim/r+Zt0FC8XDuD4W/A/4rpLSNcxk6AQz7VeIFgK8zs9rFJ8pYJwBe3N6
KkS/V6c74EXzW2B6+JfTrhGkkgL29ycQWDCkc91TKkGa997r6uCrA7sNYhWtvwrLrDqipZbC6yps
X1IwCcgI3+klDUlI2ASDmlXT197xe2BGXhbDlb1QJ9oF4L1fH/8l0Gp+Oa+mwLMq4KT3w3zyG/OB
JDF8PBtp53jEaZuOzplLqC+YK/LYIdohZ843w6D81xKy+LSRvuFfz1jD2LTQ/NhvFz4G+ME1yv1l
VYRw2N8HTOb2ZlhsdHfUm+QSpC/LpPuVu2Ke8Fvien6hP8p6IxKZY14IfJaEI+ZbObepi+XLZOXe
FO7wSDaSxInOEXxCYac8dGwPOp5jwVtmEAhd5HOOVDGLDpInhuDHKM1kujUO+tZZutZUNDYjS0LS
P9p9vuH22/31ohkjEkS6XdHoFbxv1SLd9XNr/GVmgXGeZS/nhIwtOFuYrGZZDpTX/ObMpFCM85z/
ldG4/XChalHmdCYo8HVCtSdMfPGde+dkOu6fiot5pfU23Djq8PAAC0zpCfF5cJrEb7zCicQU9KTO
ZxES+Xh03rXY7IuzJWK84jEwu4LBXSgzPW1yNO9KOKVrRZbns8ZcH7lDTbB8IJMhh9fiFOhF8lnf
ybkhjq6j+gT6S8+vss0o3v0qFxgiHIoiTM99WcIIz42jJ4ISxB3SZFlLdsKT+rp2pbflFa1bzGHs
hGgLoYzxhvnQVDW6MbzIepl7xOpeaWzaDRXFxMZoA1tbBylSmGo91iOJ5tAxjygFYI7zXa1YMpRE
2TxRXVcyrMc8RQMQsfbXigTIdmZ8/Ph+nGGaH3S+03DiHN4G8YzahLwP7XN/aBEhQmpfhAX8kYnP
x5VG5v4XO5yEdf58f6Yei2ERoitOYFAGVLst0ppnBoqs5X47mypEREZxHQbLf8+crOUHOgF44hTp
eZWJdHF5Afbqx68BzYVWIQoMcyE276faD/vgomYQ2wTPjsQQsNiMH9l678lpJtKhOwnFbWXylvWn
xoVl2WlYtHesBATKAwiKGlfom/zuKV1+ww6s77v2LOcE0ty53x4IjIYBJsJ/IIwdvHoJM3iIeAVJ
D6cd537sTxNOL+G13MWFZqZljWWPRzxujptN/OpLdFOJ/RQvNr2cEb1WM/TRORtzfo/vU7L5caII
6nMf06LrARSo7buWBh8BY5S2QcVDvWxH2qous0hhFBF9DAMEwtsRhZeqY6BuO6ySL+faWeuyDVDv
wNuFaymP5ApmDDqbBKEOIelMhV+Zy4FTm1KqL+sFRDocEurDbh1WfNkUvRxDytPdjfIf17BYxkng
tL1Yj3/nYDgdsl7OP9+gdZPf8dZPojZV3mU0PlZrazKw+8+MJSRFxtSG1ISoVu0KmLLAfafjqpow
Vm6yaVdv7gvxPnSgu5eqh/OaFHQODv4FDtEAW9zFULbJjWAKngG5SsqDAliyevYm20BD5jMKrTJu
6GUh5dPCDSip7PwfIrSLDnA1flKZ9P52t8pOzUteyDL4CoxArUwmvEQEO7Ct7NH1ImZ7yr/NzT1v
9PH6a0sGFuChP5VDHdOk2fbp1yb0cErrOKOnO440/OAD39vH41VRXu+BFut7E+zg0/F1CSnlXCme
fZ9VYe2hJg4Hj3jRiFtECTEtY3pf6tHGYldkZ58eVdoPK9SZfYCFQ3cASR/vZc/C006EXAo0wZUT
qbgSrVxmQ6mwd7oUobLHfSshNV+CKOXpbJEYm4X1CNW8DGqhxCko87Ufs7KdYKwnjQT2ZJ0+mycJ
eoiiAryvghPj5tCXbU0QAcihjC4mGb9kIKeTnOpqCFxgCTSuCBNAPkv7kbDi1CE0qrMsHvni3Gt7
8pqU9bUullIgmuWa9f4UoA+pySRo3sgV2CEHSRk7gyRnEULA/ImQIlyeaYJUdysvtB6eaibPDxjM
C9dn+AD8CXOumx0AYxmanDSJA9fTRr+PpmTZ7Zjs55WkiwtwvROZvqOyrJQBZCkbWELJJCHp6Sq2
1Gp5mmG3H94t7uWifcmgd8HrI8CqFb0BkfhmLLKEIZgAJTxRrvJdjBb0UefC+cxQbTeoXiTQP9Aa
y+at5lGInfKxKXEurhZ58anDZfTT2TRjS/Yi+Hx0HwbaBXIBhupHr7H/QU1xmD9YbXpepYnispH4
bF3nejrEjEcdoKj4P0DhtUB7tDOzFEoKGb1Vkg9a5UVFRL+NcjVjlkxjh7X5aOvxDAlKvsi+07Ou
2jC4syvJ/U7qaL2nHZuddFdY9nFT6jvlk6C3w5J4sCItDJ+5CXn/znJnQIZ08jHtjthXwicWcab+
ScNO4hgfaWot17mo/y8fkYhXbUuEJTgieB1O607krE6yHl/5KumeP0MWlbxbtegUTp7BwNRZtDUw
Lh7o4LHD2X3mST7onJ4fjklaitWRy/0jYyExkViudScReIKHW99aWLNLSMskhFOnOCmkfx6lMjK3
SSSWD3BEBRFa88oMyKuvR2QbeUxNg4LnjYg653ZVQ9PPiSVsUD8MwdG/NeB3XzB93yfvHduSkTPK
23MQe6IsNoHkM7XxeTe6BESZPxjmmdDo20R04mrMvBpJZNherKd2rlnYQIJC4TpL+fsd5Ve6R5iY
3lIxF4CCJjgEWxvhcrXRviJOdjaiJJ2sUe+fKljuCEL4h5y676QvG4slgoKuzDum0FusGZJ2vl0j
unk9hYlI+fve8hkE+CgRx2M553Phl8fnd3fnOQrF5WNRIeNRiws5ZhHBnHj4guXBXXqp/uDxBTU+
/8QzkJ91CUoqaIjZdRPnZ2WZFrESB53r7gTguayXs2L6qkIMiVXIcSwz1//2AsIATyI95lkmedZl
QSqTHjPrthomyHebUl2dYspeoSsOM+9x9fwo0TqAipMcXvb+seIoG6ICO7UlhDjXwEVOIOrFIZau
epB6VE+PtB62ahVrpUQ7aX/4s0NaOSV1ADalwT7pDfNSGqj7sRqYIAsQPgqaidW24Pagu9o4wRSx
7i9Rowv33uRMs/oXxH0RALhEbVAmNbQO7lGm6pfCvXhnEUEkV8ww5AGcvHrF4m/AqS10Mzk/CSrv
Cp8CoQrDlmZ98rIzl0uThzp0yylwsoyGdjLAfXavRuSmJog15bVN6ID0H+C2LWOoRTn2P7q0+41Y
rWvxSGTmj6pd5xJDF01WT+LTgPg196pAbYIOkeQep/DqWvxvWvW8Zf+FS0o6NcR1CnVeF3Tbo90g
q4q7a6rEbfiS0DLjh6LlJQ1nQktZdsilP93PN4Eo3/rRZ5TDfkjUos+wM8TTRG4+0YBwj6BWRdL5
UqsA5qCQrQI+yan7KIy+X+J1jH56CFzeHnLgK+pOXvhut0jSOkHCzktvsc7GeVEhydJ1PXa05ZkX
LwoyVJejkd14A798RlAwJ2QKvdVu9SF+cj5ISCsW9kHhT+MPT9McAsDwnIm7nVjG8yYUSGyq9Wbo
VPxM/7E5dGZ95d0/EiVU4uGUMob1QockStRAAcS2rYztrPERUEyZZrwsUoKPu61AemuhSdAtLVfG
GkxzxduUJaFC2eWd3zeYu2L0z9KA4Ml++bp9yccB9T74otsVH1ztl/AgV7XPJ2irBCac2rp8cF9y
SFYrNOyElAsndNnqcetQx1QDNZ5l52XoBX/pRWUkFvErPxxbsZE+6fQvY7JKMeVGbupJXmJJ9k+R
RnNFzqfmAgUPvIYROw0Rn1qJokBy+pgwNIK9xxh6SeRBsDxIJI2o+gRbZImkrodmVhsKeXA0nRxj
CGTbRArdWsnTd5sKrvjPhf6L8+Nz5vwC/1FQ/PmFjNuVoIrHB3s+7aQOPIKwleBA8psWQBICXjAB
pQdhVJ8nODue0szfaNIt0Lu436VPXhq+Vr0T9V0Cveo/3e7XrKluPOPVIwhbPnR7ssYO+YXx575t
bnJ+WsPTcryJkBDn5bw9uEpcuDI87IX9OnK11Z6QEISulu06xYGVsK7mOJRnjT88dT6NpOT8Vnoo
h0jN/wiemOF9appthbnDi2Ebzhp+KIDMrsSwkM5JqeVsN/bO5nYruOQP8J2gDgWZGmUQWboFyg9P
35EZuTHGwN49VrEDeSGJZT/lBeGM8fi3ttjG8ZPtUGF67xZtz08ak+WMtXkaZ9JZpJ3VFWf/5vP7
Cp7e2DtBLSxWMKEDThkwoKKCrk6yyE9c0tuXoMU19JZyipeH1A7GMg4Dag4SFckX1Z9qFydPw/Bx
GGttvcuEBsFRtkqdxzLXQ2SbQf0/rD2/ZR86ch+UdNAmITD0hNxL73OO1kULw3RniOhe/bVg9K+C
wPl/+unqO/vC73qoqc/Smo1Txv/suTPChR1hGzPyhgoeb8pGjgf4o0KbdFMI5aGpHdfAfMeXE3y7
Km00bUlRHSPGAW3lAflrty9EadpK0/c89/j/8osg7cKEsSjShvAYz5OjsVRZK+v9ub6MnJ13BOEa
0tv8kyB7L6Z6rhOm/mcfZ1+aWcUCckYsmsZCXdK55ulBoLkonFGinW/Rs2kzn5Y2gvBVWPbKgFF3
i/dodAUqM+ATal+6QK1+0AsAN0cPQy6TexDZitzYKaxacyDdeSyrPG834H+mHkcXc1UN7CT57dKY
5FmYFAe3GHEOf7jPQc8YZXXSbUb4xwnm0qMwUAIsyNv3G94BT3ZMaaMjulhET6kLkeWZ/G0vgB9L
G4Vm2lFxfCWkAPFFviXhu/4QPk7CEPrGZRgeLqxmsDMayvixdwGgYvB1vobD8fOwB3T3uzh0MRVc
7i2yPZaLGm+42Ml7/jB+9O2Afm3VSvR9GYdaH2oRngulEMcG4ydiCfLxHEFWJDA/Hv9DNGvXlqk9
CKdQ78iuW54f4AMN/aRI0vHhaK7Y71KHKIbOKYEEYiGfExFOQDE41zXvjoSI3pVkaYoPG2CEW5ql
6GmxzWwMfmL/Thod2V9nRuqTOHCSsP4pHaoMONhmBjbGeWHZeaqkHSopgBFRD8fAaAh+DLawDTTt
xitH/sUqVh3N1cQy3D1vAO3d/n8T/XlqzbJbRT2aZAPNk2cEQ3DnPWcZXJ8/x0ktdBgQ4QTBfw0K
vWIM/Jqq4XBga+wrBxaNHVhPysXsrSQO/p+/ERyKpBoiVH/1zER9bExqCpm+l92tDNlM/oZFraHW
+6rJDU00LBK++avLmGljyUchaKSgeyhXKVNZKd6sm5N35HktChJ5BNJ2w/aAkKNN9q90V9PQrbdb
K1kaBpxhr98FMVm0ml6xJ0Pr+TRb5pkIEfgKQwXmjAWVQJ5b5RjWETFprbDqf8Qm+u+iQOs0k2jO
xQ23UZUVsUhTzJDzfvfRxzysAXwc1coSF/1XlsyW6Pd9jFtkxQmuRQpuSDia5g0nugqAJIVDq2Jo
nbS/x1UUB5hkM2Mp2DeL2UfBgDC86V6m3gLM2sdpqT4TjRF4oHHgB916Nri/ynt3Uv6PHR8xTW/n
OM+3w/yolzqLlvxHQf7bwO61RuegKtZ4yHo7aXQY+nWkLgNwT3hbh/A8SHcyDDSyw9zmC7Y1OR8h
y+zg+7GQZFumD06hyVjVCZRwTpORa2Jugfhu9P3lu1jz7hanz8/yw7gZ7rxcRr2VsGTN6pstktpo
n6f3FNTxssf/U1OLW05s9ByAq0Am1OGO2YhD/bpj2K8SQvTu6Qo+EUNAymxVjjZfp7EDaAcepTqf
5TsR7hNfnfgQrorMpq1PqvfgKA8G4iSgZl8JaYWPEWn3wnQn3ZcPJcmDBhz7kQ8jQvjHGu1LpnXc
4UBmg2AgKlYgfwenOMLucXz/yR5S5Qlm0yjK6VDaS6trVYWGEnMApuN9dg/mTmk54/KZfMw8nGhY
n4bM162j4AzQfDb/OnPG5sNa8zSMShsQZRoEP0W/6wMSXvNdNCKg6kEMnS3fZRGwrewYSP6KwLPG
McOAEUfvWz99hHfAtv+Aapf2kLwY/IrGrulW2pfZd3PFGFUe818bQk8/hOcysBxOiOjHzxPpjJ2U
FN95s/FmHk53ALO2uDj6H5W2kSbhUEe1TVHGd1ndt7I+wFCs6gJpTvPF+cE2q3w7frMJHw8IHE5o
MZt26d3qyeJ2fl0XkmW03NfK0mKg4cJNEpeQVr9qyYyAjL6plcqkjpJkSEQ200DemCjO8Jf1X0us
/e/ka2K1XaoQUcBzpfz/ZJ7Mq/47b11oPlfZIhhops7L8AZGaeisKiSPv6bF9N2k2GuQWqfxb++f
6nl7oaNVPowPI2e6b/mkMbqXlqAjVpJTWLo+KF8wNfxErkJBcT25hmwszE4hPcLli+nExrLOTlSy
tq2di65jjmTwm4ex9LsLefQ6253yXi3U6K35ZmMMCJWJHsNwFsi2UOhLWXOYARaEjL78bhoKWs9K
1X7S/s98maOmO3+T8wGco4iKZ8VGT5NcNYxclcEe6x5RaBZVOhVv8wWtBJKXO7mYCVZXN/Nn3Hi2
pMDF/F75hKF2KdSmCjQpESdbtmPEenyMWjnzVdNJLIrlBXrPF1k4gnQjZ2JrmFFCX7qIQJARtAvy
suQnlw+NYo0+Ym//tbUJyeIdoCqsvr3OmbQmFSLMG792Z4ROqFWXHbBk/oDMcuhpTi+ws/CSUxhq
2ox/LPVP1nfXHzBn8P6SIg+JM5IB1r5rD+TVnSSUSiomXlGIyZ8adn6kSnLjY9H9rsset+9PgHRj
MjYzaQ2v7aTcj6/Bif9MBQD8RXfjexFxJUdcnBKaft6czNFTuBBnRIG6c3rCTwX64zLZZy6bI6Wp
73EHU6h6m86mT1VvFt4Irxb5tTktVoClpAVtW5qEHsM98Y2pX6eizJ94HmdfexJI9in+RpKpHSZg
x9r57G3334oA5OtZbe/fH0T6rsVe2hQM7I3vAyq2MtZaA6BbvUhfk78nzYOLPaBkIMHYbfSIKqM3
FJbsJ7Up6Tu6aaNbLoK8BGhnpDzXQttBnt48fnXkchHLDzz8e5vQ04klLIw6ngZafdRhTSWeG/uE
1BvX1HnwjtHi/+TwxmsNNm2TuFbw7L+odSBNe8qElW3Uc7Q6ScmmFAqxRhxnEIGdtGiCjxmzhgul
nLwawRAUpKOyXLQOZ9CX7F1uNJf9Qx7a9VDTbOgZ27YPkweKHPSiMXYNnHIRsYqNYCtuQ7pKRP7e
uCjNd8iJkS0BU19ZA1Ty9yjoij130eEm6ZaUoNYIcjYXkE150MhSTXNL2/GNF7p2WQIgy96vuslx
CghA+fGafbqc1HWI6vztA45vEGQumCnBOdvA/8ebw9hnfSKuq9XblHijfuTdNvwdDO35prpN37gA
Nro/9NCiNMKJSE2N8JWN78HTLW3buncOhO0ft5QtZB0ZYBzDWu1dZghf+m0lBJPiLcHFruju/K3y
P8VrzwX4pbbpq7f7pc7oYkw8NygykleD2gMDL20CZrn/6PKU+azIetFYIxq8eYOvl9RpO7PCGW2l
+YybFaw6k4ZhOHu+XJnXAapNSHOLAzl3Y3lfEzl/Re1EEYRW9EwJ8jY4tnkcGahFsv+vjUahevzc
8rnZH/3bFRlOLG87iv7nfF6TvQ95FnB8apMtSP1DDqv7/QbWU6iaAr1t9H0+PAeOG1igvULRMNzo
8zn6ljGT/vdv5LAZr7FvR1qS9/eJl74xkj2oXY+zHZSPFzkoE8DBX7KcuHR7d46Gn2d9MRKhznim
ADcO1AFnrpUFLIVEiRopY067XWyvsuL7w4g+rAVL+dN3kgphn4tpqEwpAwPZtey7ZC+KuTmdPbm5
0asF0VVsbbX4m3AhsPBMNAc8H4wxJ+yEBQ5Ayswij3BUk47pR2dBuRdA+cxnm+b6z78LGqaMfjNp
elfkFqCjmhFjZZBwRe7SoZIkVV7FHQNR5oDoP/NIi7W9iTWQ9KRizfG4k4KtjD0I4sxFRqyKuKMG
uKc49riTJjmTi2x9JkRy+PABbc1P1I09R4XxaeAOzBQeW1Tkc9wr/jCfk5/nm7YkGZKilaFzi6jv
UfloHqNsEk4ghTXGkJsT7XU4K2DIMtl6SThtM0N82/ippO30f28qIhyYlArie7mimHebFlCVN8Qv
oKmF/basBUqKPBd/gtUPhMusRfje81RajlQSPHWFMpVVb45/RpWRrFcroEghId/gG+JSirWRRvLr
E7YvIP09VhDHdxVFh4wm1hT49gJ/js2OHvGGh6Tc6A3H4zNu9UoCekPegk8vCP8UBKCU4CaEJv3J
rBUquQJVVfROlyAQnkFbJa6BjpkhkYSM93MNFVZcjkeKzLonY7x/3gbMVQbm2cc8Sqks0DSaxKaE
4zZy/XLpBEwICsp3KwQN7Pv5MyylbdNz0KZxkVLFNCs+aBVEKgCk9mp4UMtShd19T5Y+DM1rCfPz
LWgb0sOiKdWFcC49jHYs+6TOz1EkcbDlLY+aPw0Jx8C9h2yup+s00mAcui58NYe3KYVj60sO5kLE
R6A0Jr95JUJhFeFStt4NJpNwAVggTbrWCMjdeGwywQjHGRx6q/clX+js5Mxu2UyYMhkuwbGo53uJ
3/5gzqVPAvk5u/jSXbePXN4dpeMRlKxsGg27hIteOSsZG75rfoE9Q2gHelVAQxliF6+14naGqUkK
qTbjlUF2nPCLXIAPiX4Vw6FzCpdjO3t8YHFOBcuPQT0Oa8C5y/WI2QlQBKdaDfaWbzM2Ih/UoKwE
I+eUxk9pc8NPC6/Nr1YK2Kpmq5WB4RnoMl+6RzDx3yMY8olqSU89t38RZzinSvHh7U2wdHqoZMwm
5wA/ErD4Svrsxkgg09vaGY0pISOY4uND0nsLUQf4r5hKve/RkLCVgTXIoyHEXWzTCr83AmOvuQKY
DSAQbsy0JdFJkgPbWmfVFT2cTibBmMnn+7Ppd6/Kz/zINMoge57WXF0ne0hN2ohLAGtGe1qTi15f
ESAEHRIqVcTqxvaG05+Qs+rfAy0U93eCQ/jA3hIOVoJla9FheJmABc+g6se2fidUCjcKQB2BF4VI
YuOKu2M6Hv2UlmRzv35QodSK43wMz9TC97BuRXz4b+5NWR2Uk8WN8GwSvccYJyhiuWNLqpxa3Tnc
3wzuTu3UJtPjqG950fYR5/6C4ob6xJgMq9+aIljZBhlosl0Rp5vePR/e3p+y9HE7VgXGuTpnS23H
eISAZUVEISEl6zJcAnZGhv4mkG2FEVVIUoe+Sc+pDqLBBdB27qDhE0q6Qqn7jSZVvhfihvLxs4xj
R0JmGPNPIIfhaIoMezrlttBcPn+MZWjMgs4qLmfuWqdBX2+u7aFUdPiE/lmCJIVSnyMT0/fOn3GM
suZHTtLJEiJn3uJjpe5zL4r5Pq8Xoqd7PV3IwmHNSun43ge3awQt/CTvCqTnFRsuv7UQq1hnPAY+
f/F64sxJpwnZVEr8gamygkjdd00nEJo5bmqBHuJSd4o/L2hYtlthoOupeP4yERoC5682d4N4EFGd
OzqD95Vg36f/VWHKE7AKQol/c4kdwl1iItdO33tKi4yI29WqjOsNNPs4zaBJ4XYxaafEVkcPqgRr
RrI5cKBHScfQGxKnrf2z+Gxz1Q8C8/M9+c977ted1evOqh2aZn5Ry1w7TMhzOPsoIGYZvBvwMkX/
GYnRhvZr9f6wVp7xNV1NbDyxB+7YZ9iW9v1X83K/QM3MXty0RxIV6feIS8B2h0DuvzdbWHqBWlhI
bhHfpfbcyIwirwNKCZ0+dRTmwyQLbbpZASi/BdTeoJ2tIDaP26tU+RfLWDQfnMBsFdSHdsjApdEe
rz2Em5po1GghtViGICAKZk3sA4W7NV9eQKGOo2C4dymJbfHz6IluQkqsNmKtlT6ecG2gEe1X0e7X
p7a+x0SkJUXh85rxwXJzANGqJAZQUq1Mt3Nc/KYE2x7OTIdyH0DMYsVk16QveoexrlT3YhhI4CMr
qVk9mVSOc/vR+B3IlwDqmZHX8HSS7xTdwJIOHC8ZUc72OJjWlVjUWElU/QnuDlvyfrEhkK4dEVpT
Ex56x8ZAObl3E1Oaqw2EfKph8CSjupl1OEEs93uYXVLa1ZkRxxpNo5bdhjsTlkJGyPAZRdl8ttY1
O7m+zPyRx+k40swCQlXSF7/IJxYL2efvyB0vlSPIDVbwhFp9hqlyW+hNuJwqcvsg9D6xpnJ37ea8
rJY7ZY5AFjnnvtD+3ozMNqhfHR7YN4VSHEQYk1g0IOn2oGfZy/1xR63nhf9QHngFpb9ebewYf27A
2EZ0Dwbi+mjLp/kF/nPgTxtRR0lBBpVAwFj1TNK2B2XvEtW2h/nD14MKpfZdiaoBKnXiw0jFc8NC
+XeLhO+fQFnHt6P/Bd7JxpDkpqXc55Dx6zU46E+6yjMUtrE80YW6Gonc7fsiXOrblt6xJAREVne9
Cf9eBeF3VTmDeMDkCMOpGv6TQyW0LDR0azxD/UfncnN+K7UtpeB6OFOv+kXG+OIq1Oh2iEqzPr0t
IENwgKk52QkhKaYDwfuwPE92lae6oei0DwkZAUh/ALiq4DCGiQ7uxiuQeBFhNochngDl0BUw1i25
nY7sZXdB+3Hk3QjaGEVUATgBv3nMb5QSU5A4F9S8JL0H2R9vtznq6urX7G3qj4q68+KxGVUdoBbu
g1eScrci6Uwvp4SKh/d9vUuk3XbhxJYxP/vJb5vLAwreUQkvMy98AyK/2f+yH9fYgGfiaSrAfd/F
BQGAp9rABETjgyf0/NfZ1X+wgpA9GTDLtOsmyjqlupqNWZmw0TFbp5ZlijMlB5u53dAN9ayVapn4
J6iOsLqzDNeYA9afVq7wViZGb6wVlogKZUlk8sbYgxcVLrw/A27gWw+3FsE47weAXK570Q343pXS
G0b82kfeRWS8GJBo1s1T/aAcuXS/uwzwbhWs7JY0rlgGwo5fKHIoQQJwoNqUiuwLX+MDJKjx1odS
gQSxskBKNAl5VW/j26XwZI1v8fXWmXCf1vVBBFRLkG7rzWuirHj5IQpm/Nw10TQ93Y8w6pMYbqzw
VJKa8DNMEQmAuLX8qlJ2NAdmG2tzpzDrW8OrQZg0bZK5dFMIGj4VktBnpCbB5DjBSwPUEWUwPIci
fvwvpIG7qrP8p+Nu2f+UavspPdEOjeorwZp6Co9kvQmLAfKnaJVZHDwl5QpV6VW460qbCflmjEYE
N/lkfdwqeI1lYnhqFBWJG0+5PgCL+6otshgHnN/IZLAj95E8TWWGfkZ4Zgb7KSbzViCeKPR7j1x7
wxjWoHMLhCv+zPpz41iGz5BJEpRzRdu68wf+auJOfCyZ4tBqZi69X1YKRkDGEcueY6eCr3UTa5Zz
bchf/87LhqITv+SJCt10/mdZsjYDMgAHlzgwCdeAnW5xTFEk4WpMnW5RuIs5lNxBQdRwua7s+593
7CQ28zzma5lPRLKpSE3DzffM5xg/UCjxVJ2GH3/09+FkIYvZJZDlY/OkZYN4bNN+he2LZdzjgbN+
8i+YpUwLhuBdpH7Rqnfl5MnRwV7keIfJoaGK0qDKsQs+nhjPt1fSTdHKpoIwE+FB63ksArBsOm9s
p8MEK6lu4rGYKhcw49KLNnqwoIibxP+RKFGzBc3scxPAXKNYYcEnuDdVGZ72mHhNku8/N5fG9ILV
3FzHfxayC7yxzVhA/QK+RPB1xZE42PH1zaLvHBhWR+1jE3bbOI31KuvvffsI47tzIoXv3i38g6yW
RfvWLgq7TtT/LykDlTSj/fCcU/vAsNR24VkWq7jAujhNAnmwLVuhqdn9c9cdOX1IxSHw4WfJMHS/
OGe7E61n2kikOjGUFUBsFdpCWmFbx1ddIDO0TGoZ2kAJLHUm9MP8PClaUtRXAftbdjJc6maCOd/e
OvanS96Jt/IojrCkNOJNQ05kN8nk+Su4Efu4zWrRyGDDt4Zw4JNx8dYdgpzv/kJQeIctzgZ153lA
6kd9vb1TosdEq6OMPVEm2Z57RcQch4RafHMeb9J4chyBc2gcGVLMSnjeSdncN5ptsXM7jvJhmoFG
O93mO9RHz4yjiocVIgU1RYPugjiFGZd7xjBHWIER3WUvdTTDx1b6uffq9GDERHf3qzjiF7cM8lXq
tWxxuElBjDgnIeT1lG+g7NCFem00Uo3KNPnXvAU0B1FWux4s3Eamga5xthhyxvbkAW25ULVtuJCF
hUzFxmt+/UtxrIcsN81RCSGIBONRgH84oQI2l/WK0T2stXOpMOmAegnfLDqKmGDWRiH8LWusbTDP
7C74NudhGdp38X96jzcw5ua2L36eK2Pb0qIYJBFZAqOPkt7R1Z45CZwmKF24v2n+8xsSmsy+itl2
utdxAwY66SfZiIaPw1P3jki5ulLWShMTNtSAAb4/MgmCZdybT1t6wZPJrgYxFGxD0jY19cZl2El/
7pEx8HQBuYCwa7aHTs0d+XqDN/qsIZS0n+zKFgSAdnKTiozdu/S0XR5H4ngjOvmTwIGwg4lfgt/S
9Z2r0DtwPumLA1MqG0efIo7yjNafAl0nHwOsQydpNdH/rBHcDEGqwb06gssMo8H9GIggL9dVB/TP
o9U02ewkpxfZe7bU5QBJAW7qylze+t7XnZiO0aVFJllcLBt1uxWSF9LBFk6F4NtCuX00ARNUkJ5i
Z+WlSEhznYvx/VxyT8cjF29b/U8tiGpXmcEc4YPC5llw1SOvuen2BqerZmdcjepIh+uCo3rAWyn7
6gY7/z50MMlI595TCBYYMEi63zfLqS2iyY9287HritpXGazKGfe39nvXP3r89Uhrtj8IjhoVQBlb
WbdL2Yup45L4mFu65FNtGJ2SQJzceAeVwXEeP0nTnYCIqk+UG0VYY/yxZ+n+hewqY/ANkH2eQgeJ
VCPhr1YTS0DjjJhD1EHQ2eV0ngqu3SdfD1z+GeYkV2Ruo+Uh+Js6jJqUmMwvCT4eR58Xfuim6hKp
l17QHIwg3q407GsGJPh0pHccl7ufPJLCI5v22rRHFBOlXnZw20V6Ymck8nnfjFqYeWNbyVZqLixQ
419i/oS3p3yWDyM/I7iFqgZkYTXPndjCZQ7CxzQXcKcXlAR/Me0f9EWjzyTo/dJ3Le6nVVts90TW
2LQ/6PWjmGxx5IOhEjMq229KsAG/RA3G+YZCZJRvujB6WrDArGP2NkuEXyJt7/AIKFBbopTiIPY/
IBYQPoPtFgPAno6sPmSn+Sub0oRAReuReJdTqnKvi4SnL5EZsKilI1/a6srMcWL85RhT4tPMvZDr
DJ1RcXRmsnQQRFYqaaM2j0wS3dToE3XmyRuQrEAUg0ftMV4c237kJ25GHwDTQYAE9qZ9gcQ3zHQF
V55uWbHZT3LzyRjC+ZNHcYhYATdKkQKAMtxEknZojgKzD+K5QgyYbro9M5fOqZ/dOdhylw4V+Lk8
uPCQAAC0/wJxu0l0TVZEeaHt8ekSSV2kT8KbCX2S5PB//cFAx4wd1MtTHkHFpR3CXX8JGTgaIX8X
3VvstGIdKux7DBUHcchmr+DYcn/zrGP4t/ZhE7Xe31gaA1QDOposIqa2v18wfOb/P1XJrmpma2z1
NYWuLs6BlKXA/lQCzDivPQfIIrCbs91tahIXk9REFNnpypVrub56bneFEeMZq1Ow/3vOD9BLyVdK
3ZEWheTUclykl171EQYCpoD28gsIZdcFqKBtKVMnvBIIo3WJAyo7LUyLThdmD32ThNT71ravhHGf
ZcyyYGH+CwdZcGgc2kQfjQtNxLqnFo3zu26TWUPa3Ak5FrsYmbbhSoOkBCw7KikJwxBsu5YqT6TZ
41vm7JBaF1jhasWLBxI5dgzRC9nOuc5rMZGKV19EB21c4O2KAk4BS4xFRZfZbLL/istdS+Ny0zaG
iNo8ygnmAxLEhRh2mutanNt9mA97RiC1unUvqueuNfm3BH4+7Ctve0G8YsJC2q+Hj+g62eweXkLJ
JTexJKzBzIYh/BPhicTOxLm2XJQ3lUUsc660DP/NJkMUzfM/KPHpfjk/VipqmcF5i85zXlkTyBfy
JrRXMMN4lR1mtmb3lRhga97ljH0OCxQXDaSrroZidGjIiNK8b8sRFe2o/jLXo0DaTjvln/IOdWgR
5MOWycH3wKN+PrOoERchuhBGT/VxScQWDei4iyVFzGYrXlWwmOdZiJ2zwC8phiOF6WNHFZwNnqpg
ysepfWicvCjcPA4+pX245oZ1simpPBkI4OS1eGSeqQQkYDnLTZ77UILqamK4gCvhV7TN1KeK964T
dn9G1LXUwhfoCKveWEaD8kcQHxNsXy3gyvOOpOw3sWad/xADunTQTfIbYavdFADxvYoikSeUcd9U
+/mLNfCKDEO64D73Cv1LhDvtTcIW4xZX8SYD1f3sSAY8bWXD9Qo/jZD5iYle5Lx7rGruet5shXV8
GdpcMruTX7AfG0XWL6zA6HlC5NDQ+x9rFEdQgiBg/SRc6/yHTnrfRP1wUdqg7n9UvuiQL3T7B3I3
TkClyPJheNO05KmWEELKuY9ctjDzJrR1mYSTcxR2ru+9+tFARIWNcz3gdN2Z8/a/uiAwmtTlIsrj
pt294t7Jb9JJDzWcog1xtbejAYl8ojQYdq08HpBSnjDkfsuUH/R9eEbeoypHYllW7GWkU5vYQuuE
HXZiY8WDI/ZcwRkgQvI0rg3hyxJ9t7Eehj4BPIrEmy+C/VUkB1UgbFsYphjtFIfTicd43huuT+MC
2Ejcu52b6iAf1aClU9O1btDdsqtjuqW8ZgwShiiQ6R6LlrA6HmNReudmEA2Q2+iNYxSHFQNKxTF1
xvX64/Gb90tnRts4vkpuFASydeu6UYWwzRWi4E363Mp0VkfewZA8QWYPmZ/XyIbC4vIpyMSJLWtb
MYPTv2waOA9I006dY06v503sXnXMRp5IST924y/NA3w3aNypgeuSOxAHVR6FhtJwWbMBghtybU9s
B914sQJq6W0SZXR7uwr1Wdlh+74OhGVgVrJg2EiUyd4wqtBPksI/GU3JJJsqiH+6HB7KNOEbErVe
orwvo0o0xDfWcBeohmHgQezWu49Oa552ktEZbwiWPdcKdafu5eZlW8nMJE86eR2uyHVrK/2bpVgZ
8uh5We2sWR7f/5W+KWc4kF7++Vs3fhe0t3mxpiLPuKrATlgycu4zHs47GtuLlfRD1lURA9HK5KQg
uwrx8u/j+WMXiy0MLGbcc/UO0wyIQI+54efG1zcufCWyb6TzDi0VKYjw4BaWPId6MM5JcgD8301r
TU7/mWL6JFJJWZeojkbDFxMbrQOt4DdewJrfxa/gTynfWeZpYBT5+Re3TCoGGCJObKz5zPjbYf9K
3dObTRIg+TUW8r+E6Un+ZL6SLbDuuHhVHiQ56BvvxX3HV/3wz40Mo6ncDHucvv2m66fiRuleLeaz
nwWVGj3P/fgn4GYo+JFCGNoKMUact0wa9SGAgEPTknD9VzaRv+e+0XLJ+961X6RBceoEeuyflICZ
AmyEDiHHratGBcBetfThbhpbwImMZjqGSbfx8ey+MZHNZyFYXhNhadjv+WQo3oY8mgPBZgUfWGVQ
MvsutxGYTWn8MIusBB0RiKHBAg2C9sVMzbaZEfJrq8roqrBFOQoGDCO/DtFS447S071FXmFmNF6v
gWB9cTapK2in6/91ofFnNiK6nocdMHfMG4Za1KDr4FBlZN/CjFY/DPvwnz9sbRfchb+1o4Gvq78a
mn9M2tgUtIq+WeUajqx/2j9sRMmgk89wDPWM37sieDARqyrjvFrSDz/mhfh4xuU8r+dRtPSxoqwe
+yV2YzV+BJyMo7xViZWvQq98/zvKaFr7u0EKKszMpSICVjUZ9LEWwl1YsMErb7CkXcjZFk2aHii+
KuKVV4/mdisGdDoyPWrYz+9iMGhOkFOufrQl/d6cyTep9eqAm/kx1tTEqCTuNSwXWnCX4lwaoGlx
OqHnqiXhZNyY03XpUoFWrNbHC4b399KQ9g16vwRpF8nezDg3xhJQA1HsNwn9uMBN3oY7GyLWA3ei
J/OzIyR7uxH0YewY76Hjpe6KBxx2rCLsDWnZUmmdumvAd8mSltKCmtzYz0nFQ9h2TCPaXI5FSINv
Owl5kbi/M5wFb+rRevi+5ZleIkfa9RueLc3PaU5ldsYOBktdGdSXl0idF66hl9J9FFBq6teH5iJ4
3nXti0RnQWk7/776JRZqUsz9LVc1H5ZXNF4YUBu8m+d7Sc6RPMq4yKQYzIMJDkiubOMC2u4Z64sR
c5hqOqCy0iiYO8CwQfFBg4SYxMO7kPjmay/SXd55RK/VOcp0KHyvAYg/URFkp7IUC7Hoh2IlYqJN
hYOVNUxir1/sNqNAd9s7R1ExiHZblYIRPc+kPaXEWZpJCyCAFOPiAaXeFVRAbEVpaObIbFUZX/Uq
rt3XLwPvsG06/HyvQPKI+4LZxc0EfQ312iGKcwlS9m+DLkGamA37eJMma/tBEhb2lg9/xmm6vm54
jTJcg3wF1fePT/giNnaKS9ViVmyN5B8CUYv1ib54py6qtVn3w3yUlvtCA2zN/4LHDsVWUG8rAIN9
n3hW5ZFgW/G1MJUuTmDPD1KBlBEXiTG397VTKfWNQ7qthIxsSBbdT94k78b2FmGed2lhDPzvG5Xd
Y2krc0Mbt6mBgfkkZsdCeQkKsIMkbUrtlWHJTe3Zo+5p5xsS48vYc/hd1tUUg1zbzi8ygF8XS9iI
e2TJVKD0in3SsxaCmxszONihv1tWledqbKJzH7IeIik6lQioqZ9MxoUcbbnw2J0yT4J/BN8iJMo2
FW67FQxts5zayb3cVTE91XqwWr2rIOCGYA6UopqvC7eCeBwFDiqSJ+9nKQGLIzhvFtdXa3sXPk8M
mmoGcmQTXWrNOs/K5FB9tsgahnrg0y0s2LJhw0LtNaysOQ1GjC0tmrCAZtPNuGSKjL1EY8J/Hag3
hGqo6numaI6zg1zWWPB3+FTguHU+Uvg5+M3BnGi4Aq5dRsIjFBzmrCNV5P9FKRKWZZIO4tUhd9Cg
Znk8IAFjPzJL5qs9i8N5EPvrlCkUGGX/bI44rAYJLWDnHbXini4HaHDIEYNSD2Qvg53T9aNVa6NS
v61Adn1g5f55A63yChIoN2HHuAC0FjiiETjb3EQjiA4sQ+bweMmpZeSGgxAULNZdSqaNiTH3L+/O
aKrkvgqTB0JE6utErSsSoxYyO8ixeS4SqapgS4g4GNq1LpnOv5lYWd0yq/XhGjJ/oD1iQ98/Qtp0
qATaljPZjxg1IIhQM2mH8kLuEtt7m3MvBtm5w7PGV/tmQ5aBfH0aPqueaIgL8xuNssa79KAnA0la
IcXaycDUM+GsgLdjlE89GfiInKGkv7c5QmeWuKqBlrCNwxz29/eFKhAYoh6oSTN+XriFQrsXTBJR
pvDOtp7oHMaH68w7Dl+o6xr6FhMfhbdDu3eXibkjFyXBWfpMEZX0iIxOb3Kt3n7J9VKocPNfKA1J
DONogg3k5P97rTYc5x/2IUVjDpd02cmJpbuBeT/8Z4YW5PsM6AvyuIhQWFjPFlDgS/q4hLqGnaz9
IWjxUysdX/sX1qFbTlviXf2naGiSFw9VvPkUbN7nvHxrKkRvUVO4Ars0VXy9vIR7nxHA1n3v2dtS
JZ9mTZ7/YwatGfIHNx4E+D4bHS9wkG76lxxWZSgVmnDQmM78PJJIOyNP/EMytQ1/TD1ZIt0Lp9lM
T5sIUKwFm6gsT0LxFpaWI2TDwNx++Z5oOJOwt1d2IDRKASmU5m9gQsvdwlkYDkbRa1PU9MtjunON
WPTWHit0JI1Vwql2UPrPBD0a0kI8hbr3q0RNrvXxEYDYpaWklcUsZRvvqdZtkYbzYfyjm/twrN8h
frBD3g4sx1bDVuA3Lk0lcNMrf21WFdRQVF9YwdVhsXc6Ux75vNg98uPqDS+chW5KOGHvCXFJgbuv
bv2dyhDcQYEl821xhwU5G/5aiSlcaz0Tf70f4BTSwUZ7MTlHtgbDWF5x5NV1UHIdR3JazPXwDf7L
ATRIe0rHW8kgAhDlsHbpcJeLqgpGdKMNr8uQFM8dpCfokIozbzWgQ+BVMkUna4vo3lGepozPGiIN
LKKSrFbhpxntPrgjGDyE2pQ/CqSkmyFXF32LpFV7nqzxsFOG0eKnihxvGqmXLsTIRa93ZH+6M+/Z
amp8rddIP6J5XCDaJbrcaZsBM2FpfS4KWltRkEvvVikXMYY4gTP0AXa2Na7ZUKMFQTcu/vaXrJiD
T6uMwUUI6IitZ4iZzIakhm6DOfLM94zRqArQxY2/YB6GtFqp5IkSSAmshy5fSe4AuKhAZn9cvpmO
faJ6s0DOO25PQWkU9RtNRf8jDh9YD4CSjIAUODVpv9EpyXw1+9oQHusTnXW41sOun3yHTP0KCx4F
j75ekTd43pun/Ll05kcIf3FeYDfOSUJTuhVDFJc8o2ljD0sXpU2Ir82IthqZqefnwTwBNYbaq0E4
i76x8gpWvPsbb7RG/lAvHbmEXZIPs08x5cpCXHvfyPLl8zxvDan/0rSVkcWcIF9kYjMjGyCiHYdY
MF6wYNHLMpeGZlk2jGE05OYGS1cAjXHVi7+fswwS93GzvOZI2nwC+pxLGNm+Yg8x8q1TZBNedqxq
Zu5YtJW/uaCeCQsAQ6Xi2M7kXsMqXN0iC+2kmEZKECa+sdcgMEbdnLbqFUeXSp3C6bMPaIrbbAbH
zhWWOBRNxapMgtdvzyfjCFcxanp6Ge+dnuihPI9aimV+5eybwZkoBBeq9CJLuCOUQaPRvelWsZ26
NaLO8W/ZBBDCM13WSa8aTt5/3lrSU4JlCgvyUAq9bY/ZPrYUjr6dMECGHn/A8R8uyqxXsH47vvzb
xkMaR7RXQ/oeFUlciQvszsZ2lf8Nzq+U3xsU61SSYHH8WEnVzIznkS5kAJya1oDsJvM9VjcDzJbL
aY2IqjLoBnDse2d5+UmAUdNX1bqMt3zgzLPzC8mDEUeqWbqH395iQFngHTkd/yNXKqn80niT03ZR
dUwLgZMXWL35w1tzE+EbLXa47F9/WzQWmFYaBC5uHWHGGBLm3ssBiZlWR/YeKTyqGTAMMuFXUgua
VIb9afSslzvB2BiOd306vS2U6pediueGfvhkt936Qc0IBMdRf3KBFSrBz/1gFa5LUhbCP33VHhoC
YFpFus3XMttIih5gLo3ICSCCoMuOMwmMOrcmXjj1DoEhaytDw1mWm18AYc2FA7+3ldrtoRrlNGCP
n/BI3Yd6qnZae4jvUHakA4wNOsRsRc7FS0wm004FKxzlB7nKOzfMHRAVaYDVuGaSUcKdxDsWX1an
NGFqc36ZTbw9XIr3rfX7Cfuv2HscLF40VOLVE4SsgfJv2AKrCbB3YrV9NN/uEXhzIT2CV1YuxIe+
MmGenA8kxONFxuvuQJ0fpybG9IxMqciDHn2U9J0+at2bMr+78fYOTA4SjczoAfGaWWHlzA01U5B9
tfFNhstqF8jmXw0srvBapJ80LYJuDxNbkG2kpbFRslbR/0TO6y+YGrtBFnFr7v7TnYF33qfCEcT6
i6lAg9kTCKa9KsnJnxnARmyOanXF5t9EhXE9QLToxst+OMp/8YDSf+3qPDi4T3IiCnHC9SNAy9fb
Yx59PXIQolboIf5gRJkCcXYkiFgbwDAwgSHAYiL83cvRCeSIrGxSc2Z9Wccc+7rHPA3xV6e+vood
LR6SttcqEgsb0IlHBNFCs58bNXRvKeAerxiRp5lrxOFWKaqByklsCwDNCfBg1FFWfFRyuD1AyZqw
gOR/KaEbVlQA+THlm4j9eTcsSaUFQH+WduG84nNlDjvX0HVuF/nMRgr+52GWYFex8a9kSZIKa5lG
78KOGgrKd1+Y1utTbCsIy3wy5npWu5nEJAcm13ma87+sS4m4RTGgbfRz0kZ3kzgD/nfRB2wgWGuj
ZXJv8yspTd7hPTY24sWhsaTUj9aFiUISfdA8C3z+jH9a4oVMaZe/XRBcFHTXwYN06EWEy70t4guk
bI5upBULRWVQQYOEysGWEnndyqTq5nFdpcHjTNQu+J4OMyLm8Y2J9MOO8L2ex2mN7z6QZO/FBngz
d2OnMIsgK2caPF4pknULXGAEfcgKzkeSTxVLh03HF9NWn0tZ1q2kHGogUoYb0jQk2+Ehs5yvYTOQ
uFJUJfOPdVFi7F21/NoFYeqFSXWUioM7noGDLHKno6X35ZgERhcq8j501+lwXmTSZdrstZz9yxqV
D42vcWiWKJi3fZ5vUmFHnTGFkwK8EW66ETev8DlKSmmK0oF5A2t3terNjCkn84nuaii8fDRBQ9Wk
S5jRr5K4NW1KGjjbnpheV80+bWj7kWwP3pBsELMmfj9vauYgU8PFG4YKAIlvlfm5B16OIdjhOzIU
fY/SqGh/RMx3FqQ3+wz0ra+IqSVds+Hcjw/O0/LQ0FHybAhlYx32zH6uHjvaUPaITwfGjyXsHAR9
BG5bjgVwK1RrbGY659SX0+WKNrJdMZ49pTk7y2p2gL75JAAFX2gc3Ok2rooSl7ghFb8yCaXpdDl7
nFy3KtC77RmNReQ6KmBwklh9ub/x3zxGGJQNMMPuwzITeVR9ZUGj4sI/7S8CDukwqGN6AtwhJlG1
Ck9glAX2CCjZQS2Odrkysah7el8QI1lFBKxFaqXJgfz3N8v7LiObs+SJG9f44e6YM0vPDijkHN/A
CWq/DcAojjw8U/a6T9c3x1nYJlQYVfXMpXDlH0F94xUjUjZsrfte2Q52vPtlH4Jac0i1/dPczMmQ
Ntb8VQckFRGDnBHNyAXBAI2kJ/gPLKmn5pXPgc0kdy8gEx1nfiLtfDFk4fKWT8nsva7LXdhg9Rvt
cQL0v6i3WAPEHObkRr7M08ElyIQPunfkkz8HV/anr8pnXlN0tKe2JFjhJyLgwGM+C0OYFF9ciJFA
G+iGNP/BEuGnUJy/9Gq2hrkkytURQqadCrY6qFl8kZehk9HLwwLmOSbHg1W3kHO+jd6p3meD3tK6
B+bIjTX0bfHRquTICIu4YjPn9lae4MRinwvyWa8UXed6M/sBJJ0YQTY4axLoNxqAQQhOOFvNiQxV
SumUnLRzuCND3r+GIbDS2k6qXCf48634QIWhwneMrpsQhyW01BokdhN/0za1iizm5jSGeuyeZJBB
O/v4B/i4iABYXowH3vPYOk6Mbm0pGSkhAqNn81CCWsI6ONQSkCksJjy7HdbHO4ibUlU1BbDVyHFd
bXdYMLneLB3aV9sOPVHgQiHRivpHNxnsvJL6afqLl64+s3JM8MtSr/JV/SwyB+UQrHO5TxOshF/a
cnWoSeqzfR881xMeTYvlKSmmcyZFCCAWVTIDrt7BQtJMXIzBsrzKbGgyzSlzFxg+O2wT9mY5Pcp9
+z9fAAhmWPiP7O2OtM+kjIYqgQBlFZ2zEGKiWMd5yk8fXvL3BxfKtfIgDK1Ac8hAn46EqwWcYpNL
nSGjh9i2ch0u+/LfGk4OX3ZJ1H5Z6NsjCItCwwgILg0LHCnuWcRbnTkf72xPO7RaAWaAXCQUgH5O
unXAXpyMS1uzdUwUbe5r9t89McqiAswkthVhx+1yMjb5LYeRijGHTD4z3eytohRLZqNdIL4piR1W
CjDz5PQMzy9X1FHjjsSOmEqAM1n0BwxwkdADyhdp3lghXUoe2S75W3Fn73AvhcDWp0t1e3FKuN1g
LHD1Aq9CIvrGBKbYpWwZ+e4oTIQwNzUl+BxcLRqSGbIue0W7tqHf6M/y/WgHKNUZ1m3bafa1ULvj
qN9H0eU1ezbK7p3TlthtDDvDvp1T54se2uQOi+2wW2Ya1X9/QcVHx3u7hxUNkjTS0N4Y2d/PkSGB
13Br0gpWWgecWZwqafQRboHT3fJhhuiyJM1C2Y7UdLxdf1dbdCO3lhClaaaj/E1+VPAK3jERfdTU
CjRrKlsWNJhb/W1jUsd7+AvdNEgIrfVa1wNkx1IUqVo6I2R0bxKmIVh1G3+DIG2LlZT6NhMU3UDy
a2/IR2vbRR+rp3q7Aos7pA09wU3l/v9572ROsNluLaOj7zh8rke6aAP63YLJxfTH7JehKW0pfZox
/asSloH6BlTzeIcfy2N+ajHHUoPVchR50F6tiU3H/Kr0/dYWjJb+FHLizhH/Hn8ljMbTEP0tWvRx
QX5QZyoQfPj1ZykuCQ1kJcBRQsjVW2TbFfOrWCf5wGmY7319RM0N3ecGt2q35yQakwzlwCK8tdD6
wFSZ/tYtQosbOflAclwTx9Ast4pI+0MAbSYpgnHymNmPe8WsNaz8nCe3Z+YZZeG5R3ZpZrejKD/+
GUBpNmlcJ0RQbZBPos2uBdBhsKLELnJAqx86Z3n/BxdrYEMNyyabDAWlydvW1pEX//k6GXkn7as6
FS7ty+QwBLFQDy8riHQBNfSVbVesjpI3RbPqxDz1ZfX1AiyWJFlwJC3UhYyUrMfP28XyD8FfNch5
EUsBgkUTS1qMKBNtWji65DKUbm85zg6IRZmU9I0UhxvDbRlkC71ATpuoWC/0/TNveePqCDf+r6fm
zGirdLcH5/8Je3vjWhwAX/dhrE0U7AWhFsDEfnL6qTjvQJj9hQFhcKh2Okb4oxaw+GMJCqxX5lU9
EmmSLjn8sj9wcc2GkXgnIByra34rQrgg9OeXivj7AgmeKTmz4FM4cOK1UeuREixHly8l7xYMHEdb
6M90Ya/SSFl0JLM/boMIDKhrUeb4XWjODmu8RkeI/YsOijlkPOsEGQ61ZL9WpZ/ol6OSmN4r6V/N
7LcAHnI1ZuvqAXWLToqMkkbch1vcIMNa9Xck/GrDLyJAr82fEY8P0WRvr2yna3oMoeYw49oFlvCp
kAPHxXZtclIAK9+6lGeUeM53FBCt0rRk6E8DbcjyLXC8g4ZWelv4zWQrKH2jL5Yz3Rb2cQ+6Xspx
+qEXv1cxZAWI4MUqmah4HurxQhc0CthC/agKr+ZVIEXgqkoegAb1jbWTF9NpepH+bTFz01XHX/1X
6kSnXszviy495UHdgqVToTg1MAzl4UExTt46umqEo6lFO/1l580c96nQGYX3GjwmHGze0rKje/Wb
kCt1dSEmoxzBNGXZGkCEz6FqQtefSrDGoEeBL2W5qJ9AL1fQUuslBfmjvllZ3KmWdrYfAK8Q28V6
wCwwCJEi7QB4fb1bhNmzAL+0oUmEoWTK5u7dl3WQWE1qqBUOd2K5PTSX+z6FW8EgarrR8Xyc/ZGk
hdvgtV3HJnGzNLI4RmzqtROy0u8cYdskmUx0RpvJ+7fhY8/34oZFKc1K1hFUHFjMy/a3rx1A7Lng
MlYDZZrzUQaPVkUjlX7UxVh+JVsTUYy2xk5tycs4Y4lNETGu14ZFHSgXmr6rn6LvcaGWA275LGJj
bKO2hqPnovO3YVRr/QmHq6TKkqnVG3fLYfgxKMZp8+U8VsKryLloOIBabxSsfxUaSohZ/nvJxT1A
nSU/ewNyYGpkpi39t5HjxEL7Fk8lYn9nHHXKju4wz5xCw32aGAGeS9r+EFqS2ysVyWHPpKV/TZW0
/Qn+fmMYuwjqgVNgzT6zycJo9Ni7npfC/w+7/M7p8nYp8ohvMZGVN0h4jUCmtB+NeUXtHacseVb0
baXqevnF5tQXJmxvsR1GjznEcOJY+A548Xgz/VJ0J7AsCtAZtCGzbv8+6a/+ttOp8PWGktGYKd01
s8P8+Mx4JOze2vizOHTaffCBB3q9eqemD6cs+y4lPtTjrGjLz9qGo9viP8O+Mpwq5ohOdLBJLjdl
SOfvwFek+3QYds/fDI908AlhFc/5TaGFtqCK5VD2HoTHWVFDkmVk/HPsXl0bAoiTpQjy81lGIfvZ
q5ArltQjGXJ5WANayFb1/qvDKerraoh7P1LuphENarCL66dc4ep+OD29KDQzudQXjMFUkKnFWHb0
u4yaOzdBUUZmVP9YSPjoBT4eb95PFky5C5TR2Rvo3vpgFwatGJq8MZkndxiCxxAMuF5Zoco7JeH0
jk9f8oOIOVumVtT0UvZu2oEeJWzaiRwO51STry47R7fZjAAq1p8AaM+/tgSUdo+IoqL5G1nEs+P7
5mVMMrc0w5yTNtwtivWBusNglBzy0i2SpGA/zjqL8B8VWNLNPECFloRMqNimSFcrgJp5KC/Vb2vB
yN08b5YJzAS+3/AcGB23mnCJJ97ApV4YkuNCy+JjaffW2xc1C4smbA7G5CmMS8eGxUWRzEmI2BX9
uVVD/okRVjXxGparsVo3Wga16hwgZWE7mAevfVZZvSD8B5jgTZ/VeJaJNIOMw1t6TGD7O6L9682h
DLAQrWQ3idSrXGQ4eXJLGuy87RH9TLUpcL2ZAn/NTmT9zj86mlsxAuy3z38X8Xsp0/DsK+BcMqoF
QQ0TxtntJ2SIAaYnccarOlGJ4mKaWc3jil5fPxMySlx+fipvgyuNp7ZymoATDEgWjTc2IKFTtrhZ
gkVFj6pLrWvCckpdD1WUq0bn6AgoDPDFbCPAvPqIrYTxztR1j++utvbhODe5ih/PNRAhVFg6N8pT
727TVfbf26L3snbpcRoQnzdw5Y9wM4vvXLu+uAy1RmqyNNx2IpnyJPQ2U77AfE/gUgeH+2E0IgXY
+cbfbwFRtydai2JyXN2djGrDmp4LRLM+jwRVJ4CfecpaCdGut+QHAb2LWUC1OYBN1JpOOXG7H3kF
2g5vVp87iQx4dV7DDshE5Z3v5ac/JfOIhocBVcItmIoW6qXnNqpL57zi4jKWsdzTq8wpgxxc/xGN
kphsvrU0sc3cW5Y6vzYgr+V+uSwF0Hd+wx4Xj3jzGjKkl2fRwnmy+FGNVle9bBZkchKCUy2x9qHu
Fk/RQbBUWev7L1JgHYODkCM59utwJDVmYShS97xKGOQL4eanE6HfjqdUzLgSlJfyqNeykbpIx3Ot
zBEfKcHNVKUBGHa3f+QIMfefKYB6ENUeQi0sQ2LGASkB6XgwZ86nfLuPsfdanqePLOxzZJbB0rwK
kf0H8VXkG4zeuhW1pzcrLsNkIahQkPVppohFbGu6+cJOyB+8/YRdRmkHOAjkCIT+Q9aIsJLB0aca
7fbtwWwVwXsp/l7pLrAOmuK3oR5XrqF3cB//AFxz8Z5fcAlvqyFzCzQZOGQe0PoUSDyTdE8XReUi
pWrF6Gab62ow9MkMCn9v+Q63Ye/s+2ZQ6q22xWdq0p5WUtGRURFH4B4qaG18xTQeKZXHVpnQ/d6w
Ok/l5ce69xRZsqf0C2sYTG1ZkFlRMh7K9/xhpWaY6A4f846+WGhQ/MMNYXhjEeM8C2J2S95fbDK0
KiK4G1O4m7iYAaXihtNUOZ/w/Tq2w+RcdWcNxRdRc/UzYtD+Ps/0y1rQsnRAmQyRyuSh/S2hfjkB
IiIJHO8nmdScYSy+Xg22tjdmWwE5Ud/xNnWLm261S8qnor0V5ce1VHZStN5BCjPlr39UTiHVPzqT
L65zwX65ArvVTUzQX0aMUPFEEr7/i36oSFjlJiARWvBof6Z6GDyIBmxUVBodBe2oOsbpkRc/ww+i
g9VlwwpLA6gFlYONRLkPYevVVh4gom7Df4PVxjR/550Yrepp2w/MyGM8WfLOqPUmBsvHvNmkSZuq
cLgvoyOr96sueOt1LmoKLQe7mXkdCizHfz079O22WNx0XGg8X/LTRB6h/37K7kkNfa0Uo2GQHRCo
3zV8/7Bvt9GBmFyMEzr5j55TOOm53sh/8vbsWDFNlMIQ30n96J8fVOUjvS1UnUGD0Bfdj9WmCjIs
7/tMrlVU0s854QCfLeNhrH8VYF7zxN58+IxygKtiGFTxQx190vBrOkZiMPQKoLsZeYDSWoYK5cye
GAoqnKVeEdVpNoRzDW3iULCyabePbdpbxfZFi2x5NX3pgvjMprEGoz0WuJOjrmGimr2du/XcHF84
nY6vLCPI6uRZcoo0q7Mg4JdqGcFLWORCC4mmlvAcw/dokUJ1wEuBtTB9n1EZoC7ZqSjHdsRZD7zE
1KZapmK5jR2LxFz5Tb+OufCr/NOlj7hRNzCZQ6L1E55Gm3MUYKw3bDJuDfRAee1dsMJF6N7b+sl3
iMKqJGWmOS4RgqonkQ3fcsX4sfjaO6HIYT4TRG2CG8xxaiBHzzNtb8cnp3yObsQFLpuWwbaeU6/g
iTY+SvZ2COxtuA5pPve7n1NdyrS9ITbYtAqvtjjBINd8yvCIg8g/7ZwVxqOS6QH2es8ftms7vuLG
90J+Gxkd74mxBBLA1Mx0lJp/87a7dnbxuEWwJ3YwRpOU/bPAgLn6ObMab7arC1BCM9gnMsevQF58
aw1ZpuvjfzOH07qeRltXfoBB/2t+A/DxM7V52Kg3j/FJDrST4wB9lGRVWLoGk390YE0836acC9pI
Xv/Nhb79m+Aw75M4M0cwV8qoJ7tJ1EaqeX4gNc2xTkwE+nmIKfNOMBmOeczIhzeUMPCdtsQPAV+N
41LXfMbZhaGDnrs6lFy9elptuKKQIAnaX8k6jieYIycRUuQ2CEM+8VQzKJ80OM9Y3SZ7DfFsvPtF
HieuMm3b03QLD0QxMlPoiDmvIzQqb5bP54yodTV8OyXk/eBZihFcKECocyPXBsn5K4Z1hK2OmX/I
QBYjVvegBAVv3/5NCj7gTIdEXoieFhgyQCIA6ZvfuMrtBR1xjxBEz1zmAqzDsok11VL27aLZ/PQN
sCtY3cag1KeDtv/26qSlGB8GdgoJT/HSkVDtw4S3Fl0AogAr9R56FybohA4nUmNhOQ5Hp0xtgVjQ
iK6HzpnLuaCS1w/uWAXI11Sy0ZbwcexJA5k3/JRaYCVWksQ8WYU2OT7ILzqNPjTNimjrU7Oss42e
GRupsVf+qHIYHn0XJYWdX42OsLxn378IvlVu0Je5t3JU9vxyGjHpn8GXsZtqTTWf5/QgRZbzx0RS
AGtDetdEJOsS2lO6ctxLIuqfjDpyMZTv1NqSTeFEtlKEI5eKw8cXKLsuggtMGe3rA7PERy6zzVs5
gUBndztjadj6rUewQBEEjcb0OPO6HCbLddo/pkyc70deRnPHDnwiPrz60avCGw7z04YffWB6F8kj
OOJZlvZzzPb0EFY3oK2W5j1pjPrrWzs7KKhDzhoJ3M4fToo7gWWaWYPMUZkx1o5OtZg/bhhGPrnK
MHuaHjILIYnKdU6F1ugameL8IF64J4n2LGdRizTDU6yN9edBQ2IAKek7aJlNQya2BvcRhNMIIZeX
ymdVtVajDn9Fx9druYaSK4GBwPpY5eD7QT/R55alIxrHaOQJkEGWNlQtXsp8kjAzQ6Hs71yoBnY0
wMsVjR1IySQGsZxpwlKryJrb8wdvpi2tR0vfOsfI2oGHFz09TH/MSQsBxzdYrGGw77+xJYHcHP9J
pSIIwgn1nS+457qYOkVW+MIeZ1HdsZWleW1fGdVj+fnl6pivgbDgohOvkEIdBFruxOHdwgsEufsN
mB5Bp8ZpNXqp4lvK37f8tGm354uZrPPEe/hcOjJnLVewfYGBolFmk2rwPmwApqyoSCiYaeu0wzio
aGb2+Rr4hJ7kW5j0C4q+wfZzQcTKOjrMLakz4ACXf4CkQCwFMGkQlpdZRYdouijeFOaOjfx6Xip6
Ll7mh3/qq0t6LrPtwmGoui+A8ewvz8sG4li3ua1Tbb71uVRYJjeKHvoSKmpvhmi6g4z4KZux33av
4l4PgzA3isOQidwNhG2WqVOKbWJguIhw3L1yO5LhMNWXxtjk8/1uTvcO6cy5b+c9aV34pVJgCJMi
kIQnKZM6A3bjx61WpZt8pxFTaGRIfU+9pEWVTP5TphWlniBhcoImDgMi+vuzP6+t8zuHlGI9ZaJn
lnjXnZfrPGESQSr0RPZtIGq3qSEAMICgsM8ueuZrXw7U7uHsEha3ELIdrsvadkw8db4DJ0ERMHvh
idVvw5fzXuRM0tYkLub65lfqIxxInDApznI+K4Bl+PC7i1WXdtG5zmU9bGCN5/Awa1FjwXGBzQLY
LXMvOZZSyRVR3wnoyYrI7kb9qxgtkr7FVXmUMP7iKj90B3WbwHa6rMR/tlTFNXcs19F13c3x4h4U
oQo+lURqNL2GsURkMQ0oJJ+TWPOntxtbMLteZFcLfjgSJyQ5ai+STFwUdd9kBZD2SNXiDR9cVNMb
343z+LvlpvN9CokcCIiEZHcBtNxJaVDuoCDTUheqJUYEhjizKMWHBgjaM1+qF9XL9nfb5E8xWGUs
xX8DHeHX2/0MXAXUQI5bpPomORfZIDHUh/5LOJm3mbZklK/sV9B/Xudg2esKp/UrYf5Tp9oEcOuu
YCY+7BIC7yuTuJBOSBwcKdNbfdvpRPwbLMUFwHXZvnADs4v37MmNd3LmptWaEbQBnMgTNLEDqqwj
iWhvJvkhsyuSsUG3dkNJTZHq/6gx0kquwKdmmtifVfJUqU7nkFAGvBUq/rdGP11yNio1MCVifEJN
9x7wC0GnrCHvcN62jGntOpv2kSBHTsgCpEHlRPZOeT4gUJxsnv5RuzQ0c1UYT0jvyLbrm6fiZdOj
8nvOpKyDPCeGN2iIOV0PHMeJ+HEIBEznOeuat/24hbhuyAk/7qw2fe67OJmXgWCNfyYpcONkj0Je
EZCAYWAxwCD7ymohQafIPyXMkctQ98PoxIAQ5gIhkkQh/QvJXIuuxd4rDg4r3MJ5UtbaBanHL8wI
IRz6bsYUAtN0GQgWT5ar0bFk1trzK2Zi0enWUrfi2BgiBLJeoaSkWPMzayxMlFAceYKCi69BhCQ0
/tAtjn2a8Xmj3XXxZH1l/HvR8N2GTShH8yRTn5UlcpBz3imDstlDuo599fP4SrvgtOVeCN4CgPRg
ba1W02gpo1Cq/9uboRXreYUFHbhC+PA53b3vlhxt3EmWrMLaRYk/bMrRiG2+2EzFg31+UCLSxZ2y
xbK7DcjD07zYUtdCI432ptwl4Dx7e1u+saJf107z5es9CNt04TynfOdOb9M9/Na0eYKdWIPY6J0c
lKqayjXRFr1EMPdj+zNLTSsCIdaoLVrcGZxNiTlas1CcUJA1iCXeIokUBCzve7j59R4WCjZwTf48
7Ofnsm/Ry+HX3ssYZHInbCWirgGTMWFvANVEVsZfXXzHEBPZI3yfQh8c/KTk6wS5Ez+DmdjGDhAY
jGaamLBQgPzKFS2ABjWt7H38yidGNAUAftH9SHU6He2AtkxAeijwbrv0Ut64ItxBb7RkzjVAt0B/
+hK4jjjEMVYG/AtvwUaCYEQ0HNiHqooWUEqT4TMfiQxtcQ5Mst1C8FH2SHnijs7o4+j/XbgGoje7
9MRbjuyLFFMMnXOUaKCVrwMbFdV8DZYUTYFCk/k7MM2uXf+6sk715G0YcvthunMSjI9Exd9816TC
ooQ9KCsy6ENgohr2qGJunIIKjXTWzcTiMQoA5Mb1pShUMvTFdf735r6HvdIYLDuhaKSzor+dceCz
5M+OspoPiwu8QD1cC5rJrUkozvQapcCAIoPfgVyKGeRwPMuiuQs4R0RGPbhlNLedGpgBd3t/0mqC
beXUztb079jXgJxKreA/IC8Ytzt7NULv+h50EPl5txhljwxQLTUh99L2UrKPmEC9cIgcPZbIGOLe
Baa+KecMvdaYMRrrvdbMIdKnpH+KO75q1C2zMCu//aOZTuohRNJ4UyuBNUt+iEEAbJ3LAFZGzMcb
3v9ZV0cOiv6x2x7DPNTSY2vW6Swid7WcXifXeeKO9Ctp9bGOSzsP8tdoOQ/eYzf1i5R/owQk9nBz
kuFSkiJkuTMS1IPIbXBvdoSr+PnACXDth1FRNtWkHvO2D23QCYzr7VN0jDa8vCvRVndI12cbeMe5
A4lV4S+1eA1ImuzIq16qkB3gxn1XU3O7fbwP72/Dxmfo+KHOEOIpSYR/PbKtxR9vFQuM0EOaD36c
EjpHZHJnGqJLyspoEtVN3OTTHApeuEHf42TtW29vsED4qwawhfXotqZLT5tp/zTCPp53ol0hikrt
dE4HbYQ5yhAIXkBkQ2bsConjKhjtEjVkFr5C7TyUNTAZhzwT30blKBBm/59TUdjeuwVumlzgYSUW
389RqRo2yjZvC0C+BBcWwoC99/qLXEoW8Po0IgVo6hRJRqUupjZJqQxvauqtLCZeu3KJ3MUPhnP8
pgAupbtaY+cLuK8LigpRgXLV1P+3aQNeXsYUSsR8sxpFgfEoUKbWwbqxugJFT0NTZbHSwjqrhA5M
KQVezl3Jrm7NVvmga4SM7DdRhk8NxUyNAoqVbzFvG6J0vjAyFlW4iSNFesiWACMxwzsx+cnwmFch
LmFmONcxAyW55lVSb/0PhF4D2ecRAdcL6xqUkteHbrBtz0zwB2PQRng5u9iTaNY08tsKz29fiZ11
fgGtPhMBqJ6AjJJQem3fTgRTZYn+WPefDKyq5l/nyN9dGXLewAPGTE0a2SJ0z2rKAupOOEpLWtvS
kCIqng7YL70ts/RUcccofx741zqBBEaY38r7+meadMBgoJyDyU63piNGn8n4en1II+0/L1+H+UnD
qRY8A9Zm9hDerXmbu+xTtFYRSjFj5Vy1rMO/Y+eI0vS8WW+gP+itVC9IrAM6KLi6uRFcCPQr6Ehj
2mLY3wvHUB2SDLAE1UvOuK/d+zpTt5EnBzAgztMBM4wSF/oURLlHnhg00lBMHuyBsluF5/KhxRYp
3RTqMiavHoKMjzi5KgSzB0M1HkWsGWsqajnofQi4motiLF8FM1yCckCVB3agganfyRltkRvxII7Y
JGOrahy1HVZNMj4hQQ1BINJpYuaAOTKXaF2qRDSb3rh2J+E+8bOy/HBT5JZCDsIss1/F8pU2wYMq
Zn8lsmsWZulIUjcWBsDudXwsVB/kVV6UdE8s30V5ibJg+M+ixLvX8BpomBzdRT0QrJR3Q+WfiMhz
fVQ5ASMe9rYml3ZFC9yeewCUSHLnLGXStpj+WjLTxK5ZVcPNorgCG7vMi07lMpC0ljOOz226ppGq
PanEYLXvDbjUcXujW8EcK51ewsFnICf5cdNtA3rYWeS6IOu5eRtnay65yqe56GQBSq0a8X2YL4V+
ySQYnVyJcM9kL9VuVd94yyRPOyoyxBmdqhzzxUuS8NPa+6x/PepRgTqE9Us09KUsfAykA79C0R7k
fQwlnT7QGXr/MHWKlV8UiMDB9/ULH8ETScX4wyoEw8RR+KJ3kSNxXm5AGXfmp0Mau+6Utcgwg2DN
OBHtHXOuWazmK2VwZO/40Na5UADUCAhoVnbRo2OkWuu/LBBossHx3Nm7HNlG3IEHyAbyz08L1rVq
6fF3NpOzc18hhbZnLJhBuad1H5DtkUngc72vxjuD79hrnzZAm3iRAxRpHTcDqkdS7+ZPqgEmdbXI
qRp7cYZvetRXQ/5e9MsYh8GN+sIX2Mljuzrl3mAfmVyspq43s4Ffcybt+oFS1WzlHHTvA8s2tSRC
4RBGcDHsVwhz9BUUaWCFEdsRH+eVJDA/hMgeyN6V0qYDOM4/hv5re3omj/Uald7ukUqtHnQhUWtv
UMeltJj5KFN1WBxx+m3/nZuWF9pm11ad49eMIudGGfNe3sCwPtck+BvE40PodBiwP1rQfsaPpc5q
WBdkAB7vvCf5KWSMQ33HpL1hOKsV3SP2ADiqfdeW+ATgv0+JoamizocbrvlWYdiKmjot+Qxe7Fx9
p+jUtn5M1rjlpJ4JgwL0WMTJsV+IJjejh1vAMncNosKfQMopt15U2Eh808X8s/ImMNIBrGThVWlv
0EMB1avOiopiLiY2+0tRfgmOTuW+pTYQq8UMRluUY7MAlRRKIOFg4Kkp0fg2sjafkc1e8hE996GN
UtliKjMvp/X5fS6BUyhlyUGkq5nAksRR60tfqnQVRxiFasQvE+6iIUqsmjEEza5ZFkfLJbHKNG9l
oyIqmvm10v0xMhZOZcn8ARl8O9LH1etTpvZijcw8o1owdw6mj112mVm4/B61TJoFwYLL6iepiE5w
G5TQARDafsuEQx2WJKcuhQhIBYSOn2iGUYdFWbyAqyNMQz5/2ZNzW7rTHRDC45mtyOM80NlDXr07
2t8qDjUYaQ2Bl7KecgxD9czlo1p3ZdSKsaJ+/XzmPOjRfGCTC5Gj4W2UeeowDmf2glvRdMTUR7W1
7RDvskJmtU0S9kIwkfe40NJnarlQvrBoP511AfUfGffEGVXhGgDCnvkOQYFJ12uJNFHr32ufPUgh
nP7vFdqyPhoA9lPB67JBfzMrtgpejBqNXjfWiljaLKCzsUf4WPubwIg0ma7++biIlnJjldeQPFF5
K5JPFa2Fk2OVr8YZqTmSI+VTDnx0mcg3sAPlYjN2O0oV4IcU1+5BZ6ZtDegnHmScRFItZhqEif/k
VYd5uHXUJtZijXV2SC6lCmMIUXILyoK5wRTU+96DFE1TplX68HiJcOBShUZe9oLqRfYB5jBqJxzg
8JJCDyRK2yklhWrTyz7Szd+BZ7Vq6Aj28xhcgo73gbAwKQ88f+8FKhiiAfwhan8VU/g2xABMc1GD
jvnVcF44LO1WGE4Tib+FM/VfIOHLtvGv2x8LmN95KoF8AoMrH5uwDkK9tS/1OYqMesc3nCb7LuGE
HZSBmGEjf45tV/vUCihtSjn3hs9zirpuukfhXlUHubii9g1ieeWejBuI6wPi+MNkLtNXG0F4hS8X
s5UUZWQlB7MGhMXAplEMI/oUUtTVbvCM7vn4pOx3cfJeMwEelAbJIISxs2fBmR3Vp7Em/fqB6YyR
MSnblHPuGe/semH+hfbaEcL+ALdIXkv6P6NJyQsDUihpdWTTOAjt5P9wCSwERPsmcAdR1tAPkCN5
Pe7LjGiteVJAUHm1BU/MojeiFIk08bza5m4D6DZXL2H/jJYd4ingONgSgBUYiwLSYo7uzNgpl+AW
2JFBFoWhnCbZu5IPnVMInw4StCtVixZ8DLDWgcSTlf7nCuFsRdBglMLgZ+SQf+XkqYkMqbYiBFP2
pKBRSA4CzfBUK9kGM+X8XM4Xl7C9JkBJo2euroO0Jt6CnEcVpy2UhCiK0rzsocmRqhywXXyfT0Sn
Kwgt6t7U6/jY1kUYh/H8aHbC0TlkaO1Y4JYOi9gJP46G/mYZF+8RiTjs2TWDBej6c7ni1LNiaI5d
XcER7dwHAviOIPfq+bXj+vod+27s6T0bLr7lSGo0qk8tSQE5UlbLUMdw7c71QLfn1wBADcp9wH4E
TAV6NPNhdxlDs1NRXuAh8gg2NSd2jsOPn4+iyH8OChQMnzeFIrxDsCKJJVT03hypytqk0Ey8csSU
TKLrLHuAbGJrk2wI4V9HDH0we/YqrYTINUQjNOHEZ2s/7+J0/mRyyMM8AYYqJ9BJckGjsHQ5ezqN
v3n1EhllO46qJIdN3Luo8cirbkUXPt6UI0rku3yjgryxSV58gBZlPMiG9hX6Uj1SDE4RBDD5tSl2
5zz5tm8UtBpkgoHD5IKO++9R0AJEKzhNqTXQ722QY3PIMk9sOB8jWPgyCX6aXFHls1J8vBu4on+B
iyPbW+k8jM7Mf8aCyJEl6R2Gxn7dK+r1TFGrPAfE6L/lb2np5WMDYAhbJ6JqCcg4ecZMbeLoisen
WkP86W4m9er2r39O2H9wzne3cj5Box9+9lXvhYAyJmnRuMxqh+YLmSXbHDvm4gs4mxMkLMt5HYbT
ugAEtf35B1NPIfaP0mOk85WHoVmPH6r2LrQ8+aRQwPlfyGl25RiivxtTKW5maKUtsy/zUve5u8o/
PhuPC0C3iLt9l6baxO+B0f4kM3OIL0j371rbGLPk782nMN7ZdhF8bAtiUMRO/4CvyzpRZPvkRsEv
sXIE/JqAkc99iENrSYMCeTjFHGZ8pmsJLHkIKI2n6Ass4LLmto1Ix9lPKAncxhd/YUat3EU4adGT
WQIjtwyZi31HRPRg6SQSt85pL1NUNkCp8HvcIO6l8wTDqSqFeaDbMS/MhQMxV6pKOYsgexTjmOZ1
NPn41jkAF9u1j75nr7tSvBKhDUCHkK+1wZeJ8CUe4MgUEkI6MNiX/9cUWCHttDiPg/eeVJyXnh4W
zCIW83cyPRi0yrQpnnmqaQX6B4uKEZwFyLHop8SzsJ6eW6xVM0T+7LWbmgGZdu+gGP0GDD1PTRdE
b+oy1BtWO3qiQEMfOQh7hZqpc6lxmY7bi7wCye2kwUef2pNpVuBZa+Imb8Nmthym9Vo4bVsacQ4X
vM+KIxWoAfksTJ25UnElejX10WBaD6cIV/VzOzarL5vmy2HG9vFVTp4RLWi5ShHYlNIxmqnVhft3
duexo2r+jVI+yVmGIyBz7xNIwa8H/Z2dSgaR2jDwajJfGtklUPf+IskYLqTcNo5ln4uRIoz5CFSD
mtj/ZXfHei15uYO5Ug5Q0dSU8HOZFdmozg08CkaFK+74RJ0FaC3nPl9WwDE/j6hXU8OuiwJySH4b
Gcs5aQ4bN5dNS9+9YLQfO4G5FLsSmSVf+ze3JLmLszTdK6TfR0Bi0zg5K3JiBwgrW2hykdAmCmhe
xu1ws7cIy7CshCQ+3OeutcXrndxbXk8zCdHB2NAOgc0IsBtYWPTBxZPmHrFdPmmSczUcYXdakkzh
vuBgnN2v4tpMbaGbNdkiPQm73AoDTCCzXNFYwW8oDhpsnqMfmSmj8A3aAcVsbHnSlMjC8aZkE3Zj
JcOHgUv2XG+B/F6sS6d6C8kcFMlcA6j6vMvNtpD7xTNEWoY4f7J0BiS2Q0BK+Y4NRmnILDFHggoo
TXoCDX/8E1Z16SodaxFN3KrdbR0KSstnOzw0TkC8jZTs/1lDMiaKgPRbjEEZqtz8+1uTKsi7WUrT
lk6xbPfmxayZ5wqQmd/DZIfHywjVUXsKY3Dcs4v3HD42hCNV5J1GsINwF1wkA7QoZNTEqt7CWIG2
/J54W9ponF+42RyYKJDcPswraWhBVB6M3vm8d1OmC6OkQ15I9C7a+7vDrKypf8lEtrPu4RrtDN5P
IDbRCGuwttyG8I+isGayr4Nz4D5f+D8pSsQKSi6Am2ImbRyJIYu/3RYI1Jm2H5GIZFYeq552nLfJ
YuBKv8Ag/CPZpvjcAb6655MXyh/DmyGbNT8o1BcHQ6ZwsyEkz3n29GswwmFhGwi/bBuJEeGrjEQI
KSgpV5ZiMxzWxZf52NyIM8FL/O7GJVOwKD1dCA+F3F4HHbCQh6tdmVpTZZFq2Ms2Ajg8ZQFbABYd
kAHpvDmgw86OJNyHCVlGGAwotE8/ywEXGM2O174AUIUxGZ8SVRhSSRTgi9wEXHMYeysaJPDh4sua
0w9Ib2mjpygUclut64/cUUJvwkTenDGTxh6B2W9GcocxpXZ3aBSIijxq9OuuSx1T0xAOt4imQtHL
GoAQHbhl/ZQWw52ttwfdwjNxvuQLRdaQ0y9dS1iWP8T1GmG3VZdQPKktMhZQPMArv7jRxUF73W3w
QTbQpo8902/DeWeQtQWiP4/CjkrdJIfuUJbmsqhnc7xcgN4/4heWQteEE4lRQIHUhdrlgI+ufQPk
CiNxb1vZ1yBQQG1wqxkKfmfJPinXbxrdxZM+9rM1aU2lxRrqxSX+3zUIhEGQQ8DHytFebJhFgjEx
Fpfvf9BI4zr3GXkt7JGLdsmxRSHJRruAEME4xX3eLyx2ZUgISNP2MC0e1uOMsZEpadVQVDIOKMP2
kFNvs10u20xxeMd1KEi/mroEbRarWWAEhmUgT2cQ61U23adBi3qzF4PsZ22XR5wtrtJGxShFv1Lm
Cr4driWk5r6aVVlEV3MxFm9KrD26LAD7C6Y6RoS8LAZT9yVqFZC2zRxrf/HDfZX4HvlBwr1PXqew
VncukZ/dYyrdOomH3R90PzkOAj+wVeFf168CQfHI96yV67UchpkiwWo2v0snk3HBfeyOqjsIXJt8
8DzDX6MQgQ4P1gNnvplf2A1HHSa4dVNlpPK9VsZXkOSKXo9UPzCRRS044N7MtwpDyUtK7DS5qNii
ocPnmwv+HDaU52Fp29/KVUgII6O9iajdp+gto799ynDB5IlSbC7mey3J6/EcBiqvP/FCtQHmN9Kk
2uULL5keRQXQVernsIcc3q/Ap4KRoh5/uyMXXPdR4UFNHYJhvzV6XNnbegdB+nRlilo1C5b4rILg
5oEOKj8cuBAzZgZl9ywSiiWqUw2Abw5APp5tWwTNQZ/GMfKyqIvySXD/7odW9tSXn2Jus75lacQm
GLuifviWJo/DBccOt8kmWWxXsJHXerXZjNo0O7FHWCfBptqlPg6uQ4CQiAaQyrk7aIlWLg8izh9V
/xl8mV5E2eptJicvmAC3oAcZUz0yARJDEC5UUjoe/EGQkTx4ra6qf7+kwFhJxTS5gkG1VLixz4Dp
SO7JWv9v6Ybw3idGdexHQDM6/PfASk/Vz6N2FbwCOef9PVGNcbdnz323QDurjg3LcbxoitOtIWxW
hmW22tu9PJSZMeQa+J5wo65pI+aHY1AZgmaucRVhdC0UVC5fMulyA552bxIhGO0eAQq4erL0u2sQ
zOJXckF4OLiyw2R9TjtFo9kXJPvsQ7mBu8havd9cJZ0498Dvgih/L/lpSf5yIwvTURKXH8m/so4Z
CjWecl/+84JN6UZrWdb5G0ftmAZS+PQCDiaRfoX0VXao5ojcvxkBDyJEEVA5m+UwBv9yuk61hFGT
cmfV0j+8joh2E5id433nYtVXHF8x2Zmz2gOljGNAmiQLQ8Yk0vJ5WXkQt0SMEHQgmySTRPhhl6NX
71odXvj8totIJcaDzbdaD7qHiJXuwERwMafIR4WqKmBTLFmYIvvjx5xQi/qIatrJSf+3RR7Pm8LO
v5OvcAT4Wj0/PInUam79MGHcjjqD4tK7ZwFOc4gDSJGU/vK094nfnbBrnbMTAxsv67sezH7L8HlX
Xupz0vdMroHct3naHx7rBrmOEyqEpFJkADoqIvWER12AcWG3SMO6QvdJasSFCzegdHsJ9LhWlzar
ck5cEh0WVuonNthMMqQ2TjkSEBwHSQ5T016u9z31Lf6ImjypkCaQEdMIAhzxD2+7TB/1pEzojLHr
zMuvI8rCgx8aU1ZrZI17BTPNv5zdvlt3PQJA/POxSpbcL7RYKht6swG//aBm2shi4jL+bpq8IOhq
eTG1nGgeGRFU+UjU74IeNamBwp5A94DJcToDjQ8h6io9jUx69WZanNn2tjz3Xlh64fmHmI4eAsac
ubi7DAy2YJ5uzqZB7hAJKWIHSzm4MnRwOIxt6BsfEN0HkjVr9Hfk7Lsb1k9dfuok4vpsO1/JEC04
YQEXmxfiQVKn7z28nNZaslDRU37VfoskhcxacuDddBiwmjjAsqHstIQsIC8jUu+JTs6+dN/0g3SP
t3+EpFYtLn3NU42Svq+EkH4M1gttuQkDNmsChwTrEi3zcnPxcQ4prqR741IF4rWwJwUHD1zVp6D1
X4XB+6lmL4RC1ItpeyssA4j53kGmxnQX5uLCuSY0EaNqha9dhHEQIbWHAfy5B6ambsVzgUAmLrK+
cv+CaX9UKhGWUoWcYNI7twfbP2j4otmegbenYjrvOBHP8eJEe9Qa4cBm6kFHOSXRfzqHzzSDPm+Y
a1ibmdmXGal2IUM953Tkj3ubBhNTru4PwL4w+dWcYYNcElnOqdpfcc+URx01whJCznitgcjv40mr
A21pI7Bqhcncw6kSMubaX92YALXS2y3T0TRyTf8VG6s15vQokOCkvd5HEPIO5EltHnpcZm9139KY
xIM3aMzfHLigjgOlWdeGFCRtin6+Oku3Gvz4b1+6LPs1UQNckE6YooLlc27awtkDEfPAudEVF28y
C5IpeC4OaM4wVusR6NlMiz2AFWJv/FmeTJQrjMezl6QaKiJyeTSpW1ntRxo9cW153l405SyOW8aI
SKMLZtQ/FgmAI1YGMRPEceAEaSl2iKrvpjDPUXpyKO4im0aet+hDRyBWmw7DAw86R6stOQ7omdTC
U24e3LXushl+p4upXypz1+jHR/QKlTGLHU1tMuez4QeDxP4Fz3WXJOetS7z1aIhlsPMwL3mT1yhB
bxk5vvQ+uqStfr457mSrmSSSMA3wlwMMk/IJaVd62QOiLnbMka+GBOPelMueqsp/SBNd6M/+6lUW
0GGPLCWqND0Aruunp3dJSgwyvVKiK4vW14XIvqd2d4w8w16JE5zVR/CCItqyip73VJhCK4Vj5Nhy
luj8yvJevegh+h+sVVoj209QZfaDAzVTgDP7v2DnN2YnXyZhBcS26vx9eYdBA12U93sWItRXnHvi
gSxBLfUdIp91GTNce9EFIr4R9gwLDGNBeQLvVS8GSu+gidEYWg/Bb8mm+Iykgavv5OyKuBJQOFp8
YsTm67tXXKr8dweSDFSzL/Hr1WrE4YA43z8tn30UIwrDczXnuZVQ5Ea357oPdGMEi5Hc1V/uvgtz
A4iXE9Cvq/HB9QKRuNMZMSnj5Wel28YgGffuKkzsEifZbTIIEX5xAsHT5/Aiy39PPz4uCTc+PNyt
eyDPXNDy1TuO5LN8ixm+e5+zElwXkdeKU+PUNjiFIAqXtuLF83W/gQJU54TVZNis4/NrUVwlbkMz
31Z4bOUu8CIqFBPGVDykvtHh+LxOS8OsCPdS1eLtgB6Xn1DRunint1hI2WxcnRTDH8y7PQHxjfgZ
f0BFjh1DGXipOqFhEL9cDR6GE4yhHCrlzvptW10fvIZTp00vMycTGqHF0+lPY/elcgj9Po1qxrJh
BL1Bc8nOQANtiJJ0sHOgs6qH5yVMMNwVz5zPCOxo+FHo/nuRuAfrsNMGn8Zrzh2jm5B8CzHWHUMC
RPnfonxBZ0m3bWHx6RazKbdMLeZwaV7cZ3LnCmp/JLBuuocZJqCD31+JvVRMJNjwZMGKS299yKWl
liqBlL0KQpG2EQtvg+vQZWWLntPcV+sEPpks5idTechLdWmauRcjQcrjtD/ro4xBeuwAMDDq20FN
KB/LiNpxNE5cJudIZDIo+zaeZovmGK2xcdfo6Xuv5BqJKHXCBKf2G/ZifpZFnpG9X6dC4HKfG2dy
0vgW4Wio3eaQPoVttsk8cNbxb2haVyYgwqYEYNd7iyOMz7dIqcxszpuMRMuZr4gYu7VFtBhWn+Qg
yRxWS1cFOV0bjgmD6e5RiBa6+RXrVW3+uJpnR0TYXQiSHJ9k+F/2yTxEGTplt7FxEJYSJ5aIXfDa
NNo72/bU/es2LKTjo/X/nZ0KfunuwKe+y+1Wa+qdYwLOY26nKEyIXJTxEpqJ4bgY9mgNFZ+g6V6K
c4b4mMj5LunoO35ZOtm0VT78iehwa7GEbTwRrT11j7W99x9B43zfEZfy9FOxQfHpc7cUq+XqSCuW
H3MLt5pq2bIMPt4d3Lu2iU3dz+GQXralmGgAJSZ6YiV6zRU1fu0iQwYkdUAQ2OyGz2Pi/qwL5hXj
VkFuFicxI2li7Ylt1gLwxDHU/AIK6Z/dG+CGUKN4qeuccMEXZKjPhwBkq/Wn+f2TvxG7EtLtzZ54
+iH2kaElK54u8nx/0R2vdbhANuLX2uadGl8f2sW+yZTCgpMWpGOzHUmANZpXOWY9vnrFSun2iGJy
LfM49atHiB/hjiVVAZw30kUo9CQrJBtRilCAzj2sQAYoE/dnQHpE6FjauTMGdAH9K638t/lMLak1
jZR0QoJtZ9xU9vsKW+IKfPEQpHc+YI8Zs4QSe2Ko3lTbhbEuYvrqws6MqV56rZdEjx0Y5lukYf6T
626ue1S/u6TTf5UOaQAQrGTR5hW/WNMXBQ3Q5Z6y5sitzigj8VS3CFBxiP4OxZFvF9ulPbwGjDC/
rP06F4S609ZhGz3cBGfw0Vp8mvnPw4tAuTum3XYSkL4gzZheZfylXYSc+CNSRUDEoow05VhP0wev
ia2eZAJtlZPWXWQ7+gq7fAfRVpVMhv0Zvr1Hy0qfcxkgkxKIoYbqK8NYSns+7g7maV1IN/fnj4Pf
T7fiJsQ5WXRj3tPKDPD+QR04Eq/mkewosUQ84hRYDlDlXjQLTkmJNrDbQtVz/9SLO/+r71mAitnJ
ErNmNJHaeAfPpUsaZ8/9Nkr7F5Cs/QNMbtHLc/3t8IkxU+PXOsjqvuB1JqnNyqhsgIBGYdm+2gl3
CXhPCgB5QIZ/MOtbCM5pMI9qdkDROG+BQtnBFIWlPTGT3W/KCjAXgJMGZGdXek+2zvKDSjf2GT7T
SfSXS1BKJlyQWTG1ztrXCyEHe0eHQvaJ4zFuo7Si5x/eRGIf7tz4Yo0+fEXOt/eFUfcPnkrBBRTK
JK8uH8lcGmnobr8gIpvkFUbJidzoovy2ShKRrt1PQggIzyrt1iwHIF3nJ+k4gQFBPHsX23xsEXSM
MjwRULGb/4gJS4lr4HJjNe/O3+8T+zlK4RrdhNvAvkmm1vrTjZkY9+WZ4GGbL0yN6V4W1a95MQ1e
9NMZAHoskTCTQ+Pu5S17G0iQNG2pDOV+voqoTnNnpVgotqi/rOxcix8jKbQF+hs5L4zN9xrGojCN
p9kG+0SykcxW7x/6vC5pHo/yZ8erODQsT/ahkK8L2ABMJLWOmy6XwLh84xji/7iCIJHLIGKMARI0
ffyW+PqC0r9KRaPoO2tzHa2e76zaGqFfAB0E8RqiUktt6CW1t+WSq2NAVxN5FIAdyz3KkeJokdSM
BMQ410BfplfqpZOyCHYp07+GE8VjaCLjkCNXaAtm0Q5jfUrDHU2SyiJ+F50+1yw9U958HJKIY/tR
6gtqkh5bnL6+BVfEJwcwIWQQInrsMrRc0GXAjWz6bDt/1Oizh/dUx6EInsuCbWXas1eRcQUDsX1B
xWuHJyWsaTGRmGO052ZaOAOc6EYzZfUAxDXimdcpLGRGq+3GaxmJ42sg4u8nFsrAlpSbEtc2MAjU
1ljLo5o00SjljiE/ozd1i/yiaHGb4gawksCe1n0MZVH0xjGeBSYMHPNr/+8Fn5fy6je82eWfq+BX
ub143A6kpnY+jlXT+Z8obZjXdm+Gl56CHawTs6NYmXHakTPLE3Edfcef0E6Syu9LdWPeWput0qFu
/XgH1VLSOaO09C546TaXRtrwYPjjhCIog6r/U9q4DZCR70vRFyoRBnZ+nQOj/RSDhpQXFPcwHVsG
WpUu4NG7I3u8DtOoRLvoWJuz2oo89zTU1kpzWfTLJzwNLV63zBOn3IjcpafYhobpuIaQFsFOKvX2
haLl4h0NoderPs09e0X7NH8RY5GHLEfBA7wkrn4zqYAYnPzBlxCK0HEkU9fCGVooT6K1XIenp7iD
ezscwLBqQKrgOhSxMeqObqhLBW9MhzGMnKM4DTIUtq1mC//lwnzgqf52rba4nSRaZj+cBStZh7fQ
l+CSr8Kgr5dLuLOvn7M4EZNuSBbuh784/CSW1VtB01RugE4AtVoNFIGOFx1o/wUnEPsn6ovIhvS4
qkmJaHeTxR0Xmz8lqzv3VVj3S2dl4nAly2yYAEjyNivzK1jdOk7kpm1Mk3uMV5sz8EAvWuBWJ4Ct
RxdjknbH6VCiwo2aB1KLiOHjVWzGTHj6Fk5Z9ZJ++I2/YBqx8bialran4OJTMQph6QfnRln8NuHo
mH5qnSFXelY+UBHnDox0R5ltLpRwwh9uhLlWtwJPV5glrTo+Z+iKEWZb5gfvVSwt8VwzUXdrB0dc
3IGBiWlTRFlA55FySb2et2IndSsW7Hp9CvWqijTw9D5bFR6scTc7wJehDvwB+BFcNwbEqX1Ksbze
ThraD12GtydU6OWKBxWrNoxyphzIHlWgYXFzAhhqEFQzVBJojxhypUvWwcmhbu1kCcQ9Nul2Gy71
iqPuzWDjZGrZ+6Vo2/dxVrcY0uIrdkftcKBvVyVcmkxxnCVZJLK3+/BD4cG4iz8DSL4cOQ3cTPdu
iLj4fjbHOPDRQ0sX/SZUANA4jvEXS664OETVmV/UGryXcBILQ0MHwSCKJVrfcaPgL2tyHdHfz2uq
DsufWr5ZfqpwdnXGzAG7m9ePNya1kT9sXBDTE6qtLYt4rN/l4vQRLOUcqYzCMlTBICF6KPvkb9ap
Eh7jUaK1mnOTK+3WxtZWJI2OzlPp16GfoGiCkSiH87uV3uhwa0x+6JsHV2D+RrfUvBb54YVdl+oU
nX7J4PD0mgTZe/xrEes1C9WucBhZ+76SlDAZHCD0TGO0+v0Gxu1n6jWjE3x7MeFuz+hfECSBf9lt
oVII81A5wndO6LhQzgsbfN5tcbhRWHdo3ILavGpl49pf1x7PogGsf9CU98QFMNMJk39C74SSld1n
IxryWWeoBvw2dTaeHJsVGkRtMzXcqw6+hiJQ9MfTBo2AuupOiQfpUx2u4zdqb4T3ACxgxQUfuLgy
hsEBVBkZldYmkyXb+tntmcs6qxyUb1GhkotkqXGJB+wrgKSrlQOPhgtzAwLYDtaNm3oOaJtE9c9c
mwMN+zU7+9PQVRDqdA2CpPASxdi/TRZq2jNfCdW83KBCu5yUCLu8UO51VC1+awXfbXLhO2RHbLJ6
fLiFFFN8oM5X0SimHeA/PGphK7gBmYr4EIoD7CqbV1ncT1KuDVURPtfR3FFu4Sg5DIPnWIw3ArC6
v/BnijHBVNoXvDO5TzibtRQPTr2Qrc8NRUb580W1S2ul/0zyRV3ppQdPcwMLqUVRW7d2h/ZDcVCz
eZ/PKivA+2uHoYxXmyw7soExKV4ul+u72OQ9wJD6HBJjhBejuTZViOgwdTcePZ0+t04TTu597nlj
MLnIuA5sjapQ0Wp85XquJrb96ZZ9nRaX2iNSS3262WYguvh9b+hA1tHG/dlnhjJ+uiopjFNuy2GJ
uUw69rj70MQi7bQxpsGA/6vBYBA3CpfcGOdgJkAXuAyVQjnOtlmhtENKyvu/mua3yIeBAaQjn+ly
oY2v2nqgy2WRKGYA/dvzxXA5bfTA1LPdmyq3BcWpeNVbxXXd5d+lmCHYYLi0pKbznQ9MxV5TW7rg
jHxoxQHCaIVmqwd7EbsQwosGMUMOGDZPf5JFORPytewvy4P4wk75KRSPaEyHQ6BDyhMN7jOAaf8e
eysrDL06nh6Qc2v6qCD5DTA4UZNpFGcaol1XxX1F3jFrtcRoA/UYWPnN8/pdp/M/ofqcLl5wJR8k
xHnFK+PPOQkWfJBGfu2xoZ4Uq9igLe8Qy99EsYr6Uir0A/YSgo9xB8h/kiXM1qT9sryte0ZMfnE7
tAeEd+2x2U7mq0j/3UTHpVrJyTrZSa6xkHZL421S6JMHtV16AaPeSNKfrSfTHXutxcDy+4HvHGck
s7fLhfZjPx40xM1rU5lo9WKbV0xJrZqFbnQqSgINqPrZc6No3c9qixwB3M+V7ifA9kt5yAEoBgJd
Q8dBBmRczTKtooIvDFVarYlNEEU6FIIsMto8WeoqQzUY1i12kuF97ULOGQnLfZQ7T6TKS78w/CpX
j1rPYuIwxorAYTdfj0tV3SKVHyC9igTgn6nntx3OPcsaH3ShXQoqk0+VusoJm/r/EFNZKSj1/ere
IN0WmGIz10EBtUcyvWHwAnPDX94C4pULNzuEf5QP8dOFsptruRx3Oq/vfFq/l1snM6oZSXgrTwS5
A07MxCx2sSn+1Z2DQkZLSnWfAYs0coqFXbbNVwn0AdoBwZNTHXuzwz7MnimbcQRUYVZBgaylhU82
XKTMtRRLOL5oV5VVx20EsCPj5CvBXKYVHxQ83eia56+rmQFNneyrdEyTri4uvFuIwkoc7Gn1h1Vb
l5WdXNVZPK05P6JT2JNCwA9WOfhNA2zBUeGtZFYmMxU7mQdqsrtRfXwMfESgtEzRgxp0APsCWEyO
WUd8PLpwBTiP8H0NOqKoXEL4wggR/HbFp/cux42gkGtAWoHqUx5FX2fGorG8l0JHdVKzZXeRyqIn
vLmoUl9qFJJ5detlP9iZFg/f2/JkwQf26TaoXTuM0O8zEpLeJIvfX7L+BLhNIgZHWfSEGu/Dgxf3
UQgn55VYDXw2CttRci7Yp1YyGORBszecnyGUUpbeTQS9df22fHTWnTOwW70s3vfoelX+7/V9OUF9
GdNhZb/7Up5k1fa0tDILXym/ZzQKNRUJtBVy49s7cEfwsUE35nLjB99cpOu6ds2283wOqtoGsIVn
YNBPr77+TDh+8zbsXpq+3wjgOxBlVaOdNj0Dcszeek4To8giLPuGCbkMWSZ3nyLkXYVX8W2sB4lG
9/lA0llUI5O7le1mTFmoshVxzSuubZJ1+JZCfYlAyEdS7irgwnC+X6rCsOIKf1Ve5UGu+HQMdkIH
P4lQ2kU7ARNh4XMTbMjEjbNWBIPy1kRxGAYvokn3nB0hvUzrWysCw+uG5tQt7KraYiFskI6UAw0w
dTWFZPeAU4fpzJ/ICuvm8pTv5wzGLK0VmI0Lbh4anXF6MkVI99p2QGvICbcvsBhtPGWs8OgPP6ae
ciEIzEQFoBaTxcYaAYbT45GSQq3kwEsAMVxpXk9F7AC2Unz+wwVc32JRJZoi8VcUQ92XMT6mT4Lv
0WdnmRpzu5YszeN0dm44W0FwyRW5H0PfEZMJ3iK/ixzKy8Tr64JGcj5F57+5ZP7PrnXYVfdJdEgc
Upj63z2Ic6bitKDYqm02710jGJ4XnrUPhP5/xvNtftbwBxvFfEQVb33lOWJgv48ppRMnEaVND1f9
RCooHxEMikZRK04E2hFRW2tsrEGwKdkfTwaIBUYuxxrxbSzQ3K6XfNjesx+mdNDEVg78DFphhF0e
oXHPNEdsxgWBXy/WesO3Lhj2HOTSgeR9Nwqn0L3ABINYzJDcdoOdWNu4BZa2/87R5btvyzsCx7FF
MvuIXp1hJi6Af1i9RAAw+9rnCT5jpjvwdrtaKs2AhkTwNwWpf9ym+Bot0PRTNYUlPddgS0yC+Wqf
NSJJim1mwgnbb0mczFaoZYYVZTr4O8nvv4FreOMSMjnO/x5O3kUC+kYlkp3u45t4k+/0Eaw4f+JM
mcGxyZ9lYmadk0lPzjImwciL5DZrShiaDxPNIE9+Pq23/Mxji0Vb+CyvC9omvrn3e1P3+ZBbZP+T
3XqJkq5DrLhdI8CuifCHxfH4ipwpPMAk/A9/R6Mca1VIQ/obrWJ8A1E3lTCf7ey8MM9qLM20pem1
q42JcdrO3SA6Dyp7NurWbVJDWT2sCA3pBPcFhh8d5W7RyC5NtQ5YXQWFgQMxe6aP7lKXbzvl9rwD
NZI9WYMrUx+Kl/1oqTAD8HT0XnIIvDd4moKh5L90oY8j15SnRnpFpBkyYqHHfUNyrA6BQqAlVwbg
IwL/N/ik+g4QyTn7djFsHJjjfwKnJDCYjbcbtm9nguKusFzW84Sl/AJYh0DrB1Tk8cBkrdIJ+OqB
nJD4jqwZp0oQjm/V5z7LdB607D3Seb2nIN1OtXWK9TiLXxvG/SR+/0N2Mn502qPgaJTlo+dZgoXk
VNtDPELbebKO11KJJou7W0XcF8vMzEOvBsNckMSpYgg3BcnhyWdLM7h+NYi4W4DWjznSxeH0cUqh
k6fH1XsPgj1GNQdC8OHWypqNDYefGv8+6gukcwpqC8JvKpIBu79910zbCrcZezFqQsOT3nv5eqXv
iBYGWC7zcrWoN8s353QUB7D+CT/XD1tsYuco9MP+UeqCZPZeKNtWglZiB1cKFnw1FiUgzk0aqw8K
qAS2TOg+GrNON/RN6bBa3tGt1qEE5BfkKBQAHSydlaNbuSEMXvek8lXqGWxXD2enqMP8WvLmWBh0
89Lw3UJVZvhUmpsYr7m62OlZ58sSHhUvbuRfozMaXp+syATKYZM5Nim/Q+Z8YIZ3Pm0bG8RePnmy
rRiLhR8w64Ytikpiq1SPiOzOQtEzASKeoqHzs2o3qBnCjA648va3X1FxTWCnatXQKr4v/efK8npV
ItEwXznAzIzoWWrAgvLLEf7qiKxul61e49DkT4UXSDeHIoKPuJBTiBZ9uXDsa+trz1okzCtYIss6
f7iFxoISVZo2pzDbZSrw8YvCoiMTBGMkbhbz9fzIQI2ofSlrzzm4TiurPSZb9n2bOd12gpEzivLt
yksV8627vvCff5P2rgnePgd3/3jKhIxsmjm8FhMMPf84N10UgNWAqI4gg2XVyWKoT4taFufbT6xN
1LhWr4GENfkZfjFWzyJSWuzTEqUNzIawyzln1JbG5fxk7KRh5RNPLXCMADgn9wuORiYsgt6NbwD3
Gd5J6gjFPWl4dS6QWIjXycqb+oeDbaiyUkpR8Ugw0lqUkv6CLFkGhbApkSecQsPonCzHDD+U5H/6
KMyKwTr6kTUTjelH0920MNvQ+TsttRVIO5HvBTQgon9Trwuyy/FRLxwa37ZyJDEqBUv4QgHvORLq
I2pF1Try2BgIJs2pYoEdo6lFENzOMFBiN+0poXzkeyfiNR68wlxn/+wjuvyERuthgCLS3MRGcbT2
3/s5BqGNKihvHM0E4CG8JUE7YL7v7NBvC7+FYNu9Z8e/rXPJDDBLRATC6+zJFDth+khZoFtID7zj
ycR637u7GgX/aLKlHGkGJp7dXWSoex70DBaaY/opSl8Gn7j+bBGzpL9tm0q1sab+MMuZlzgK2Di8
qrer/aTXWYGE1dBPi2dJ4e6FlNcfL+rviVWWiPUG/gMGwOa7uZnsObJSr/jIb7ndDKkTPuNptIpk
LbJorv7YX8kofPikSqEObRSKvZ6xyfrNf45vpLerZ6jYQX+wc3fiVLEnnOzfue9DSLTdqax8D1Yd
TKd0aY8OpSuKcrx/AiPc/kedamYZve1ZUPsaYAgF/mkBWzjsoBrrYc7zmP1TrwyCt7CEL/znsvI9
FaOX1Y6eV0NeeVQSO7c5RGZgyFGus7txnWIPsR9FW7StKueaCcNyaUZh8H05PhZGEnQBbjO3zMOm
3icGNGeKfpS+Xxsg07hfsKnHibKOO7eKwEHxTLVYsEwRXN7pr4lkYs9wAAHQd1QBrRh15Me8wGiL
+BsGqCyVWJ0cH9sn1RKNyv1pSgPmmLJ96aqHxdulsRDnsk3wBLrF1jk9C/mR1Ct1GP2p858+E3WO
GMuxeKCvwaO4+Ai+Ot1HYwAr5oHkxI1NCj6dh5XdulgTKGU2X+V9msuv668z5ZA/0hqnr7i7QNEq
Tdf5rz7LR1ECZMjLqyb5eDeCHkdI83/vvtLKfV/K5mJM30XYrTdqQCxMZZxVu+b9t2iZULoVww2c
qvgnxGdMAWrWujEf4QSm2KuQqt7sUibvcyV4chg2CpCyKoF7D+k9cR/c2FGSY7kP/3/GTAEZBqdr
J6wNaoIErvwbJMSdd32rhmBThfOhXY459Ba3J434JkuCji+cNezmykneNBgHMYuEmaeDtN7GaMjL
djGkkhLy/HecgEQvRUxCDDr4uS5uLh1UjrRyHJgjIiGjXMcNcX+EdwBYWyRIEkjBeUBCHvnl1VZ6
Eus5cEpe9+uMtmjQWQLo3A+LdMKhFbkQA+TjzLGVrWxzf0/XzOa9J00RtoL+Zopq5tkwZ58WTRYT
G2FNM2+tPHRe5TeOtg0+qd4QoV4eoi8xLb0dNYPRdMKKCJKTDnQ9Oq3mpVg0SpZWsoD18+/wBWgK
Q4H5lifSU1j694bgds50x9ZZUUTLWWcHCTCNJpNEQxYpZLWbtS7/vRU4ZicHYELUB8xMkoKjtkFO
FB559QS6e+0yTXH4Qzp3Fel8YbMApxHMM6LD5JHWy83XEAcKkc0FJndR7TSlPFUhp90h2nhqFKxs
Z94WFnB90uvz8U44pI7FiQgAIs6gHfmMSlYwMQ22pwviQF8j+uxSGQoHcyTaB/IgA0AXvrWqf1rU
YxQ57RzDiA3BGcdTmlvJ9Hn6Ieh361AZ2sEjSFbifSBBomFDZUqcMHB9RmalzbA0YUyw5oNNTxQo
yf+mgz1Ps4miIE3aWDbUUjyjf0ST32VGugVFAFlRrrJFrgZMDfPnfUIT1AInafREuwPRNa8Mh2zF
EA1BF9gitvyg8E58w2YG9vPM8mTp6xGdOFzG4GosyUdf7ivMs7nw/jLnqas+RezhnnUg7CiRkvFJ
mpfq4iAW4ZngvCB8iW2dsfS+6Xo8dNL3v7wf5mKUARC+7gYrQJ4kTPkBhzwme5Yg2mX/h1bSeCxq
j72o9ORyRMmrQvaGpJRjzF8KPWO3v3DFn4NbCXipFwHrS3Zm0V1lqRr/mza1cfwO0GPto18h390n
V3MvYYo+dQCIiMCJ0zUY6xTRLeTlzpirapSuxeU5LAGBcc5m4qDSgKQyOgLep4l8SYup6K3q9xd2
oY835c0VdUrsSiWjt+pRqpBlN7UG7oPuj4veZPYNZop7pjQwM3BYuG1FWP53vUdw2ZuiZU8ffK+2
QVGjWRGhzggq1I46c3ANhdozByBAqrv0jEKO2wHDjPC9Iadlz/vSPoEhseE7JfahVvk/jcU7jnpe
EeFon3L+QcZ514mshXeox03iqh5domSLlK3DSZ7uk1Z4rSGi1PJ79QuqHCfAZbXMO9cMY9+VEn+k
zVqd9GAjsVHjJkEKPW4DN7+iE5jHZDOOUIYmqMOhsY0uqtlZJ4RcvW+zIuzdk6+xkZaVLFqJXz1S
bXG4RLoPSNS6L5ilUJwjkcyuut91CA8lPhbnQPVZLxAratMLROK0wAKdaeJnbGw4GsLJCbaZVP/F
e6Cg8zg+1AHCdL4qPROKvqgvNj5pVm6Kic5Ae4bNCocPPfqCgouOsAIHp7aFJ40ujhz6ScJ5awFb
hPxA4GmZf6qHxYza/BfanGSv0PZTn70xeeuMBENlFZ0IU41bAfvTv0oA3UIPeb1eebtyoeJ65u/o
146/JWhGdPQp8YVRUrziUwXQ0l2zBCHtMQPNOZGCxVYAVS+Z3aLX1Pwlj9r9mjw1U77zsIvrhwrz
fiqQ6a1shMb5CyQaUOj6PS4PBGUJwPamEWJwwPtH8XQH4nyefMn3W7WwUR3l108tPhmhLSWIk8jm
1y3VOtgupUzlkugONsOesIduKj87BEXA7UwyPt6MiGJSZsrYwBNCjuJVQ4wo27r0f47F6A2T/FLt
DAL1/nyBT1GlKaE95ylFbs0JY3VOnCmoYRzh1DQWWsCY6NbnXaZEXrbQAjRS6dBl3PSpamCpnnj1
SRObYnrVcApGCXwm1N8ioV1RxsxWoVmS5dWI8tieQAZT4SDj/37p1XQgIF6YZ559T4BTqaf/5N8s
UWcq8erRGix8liADHDISVonbhvFdEGn5Di4kBzjq5CyJBI91cCEywpy39n+/u/7ny+d615XvCQi3
svif/XGfnx4blz/fJ/WGNGMdhqTqe3GoRssqBHm171KvebvxsAYZGxD6bOVvQYc4DvSnEfSPT5gy
rVjQ8reSlPwtaLeQ2v/UXJiMDkkg8/Pv6JsZUR8DqLdvdLF+bma5w+9befHJidVfotyMTf7WyDO0
5KfUJqHylYDJeHqbKiJbPXBKZdZkw80dtQvHW75vjw/FrSFTXwfhHXRhM9vykb+zbIhX3q0oFvqj
wCZ6+TGj2VQLT8zDZ+9rxUafnoe/KcFtMQLC4z2miDIeBjR83GP4XVEyf3DEfehBdHyjz7Lvedol
bN0QIPpXoBkkuXK3hTnJD9+LwqUp9BVimFCrEjT9Ge1CELhJQ/Apu5ukFfC+vZjf7vzxcCfQdOJX
BmEnOwnhQQ4Hfb7hzev9KaTs/GGrmLJfVyGT6By7HFSyizQoBPDDceicZIv1gmWNHRNCsqlpOCKJ
hfxNPu+/etK07+f+DaoaJPLqdU61dgxjPCQCXSRAtSnZTXl3hn4cttXuwyPOzACS03nGIr3jVt1o
dxvHEN8XYs6fLa7m+XbQO5Ohz2m5btCm1DeWbO/KxMJeFXFkA6nCunqN2UvdmO0iZAGKnPXIuuS8
N1zqykvfSg5s71eCM3bTiTeY4CrWGTPv2Lj/CL2M6kNuNBV+KL1mUA/tInEn4dGSannLt3wtAW6m
DlcE6righGRshK3vD74fIWsfU3sbd9Ow+miMCaX9SmUZt3cV1jb3y3C8LyPcrVcg3XmjLRhInwRh
+P4PkGLp77zV/ISApVYYyjyDEIrH5D1typyf7sEVCh1LnUr3Mf2nLG+zFWVEIUcMWID/oRDoJkFe
I5UFp58YD0no2dNoRHgnG4U6goie+s/cB1DfchsEy4rCECwsHujfguTzW7AVWzKrudMwhxg55FIK
e+dTPs247HGEbZ1nAeAJ6feOPrFzjGwOGg5kcSKpRprDDUeFrW9kf4Zd7/xZxHa56DqxEEat/OBx
gFNjhTyi3/zAGRSYmc9btb6BDXBaRHxz7lAQr0aSG7XXeXX+EpSahMpY7JOQ/UFtw502ynKLVGW0
KTANng7z9kQhYiPVPGhUx+7FV2AonnazAMn9WcSMzNHU7XiAqFUOrNI83Rj52p72kZyQ78Q4jwxo
rVhM32uzaHbhREt1YHpH9BSwbqpg7lzbDZ+LYq9sBPvs/6s8IP0+Z9Sa7BClO86HAJtkJ6LkqXui
X+O9nM5HRefYK8ZYbvE8ailY1nN+c0EL98bpH607rZZlqD9SJjNSpHqW135L3StMzReotRFHpi/e
uz3DxZYZklIpzxTCYMr8M3kJ4190HKtpkiW6BpVZmMOYakY6s1+TRaR7Az4sm32ErgtXoXZbI0RQ
407Iy3rozZRInpN6ilkcQGZE8kxc+7EqxTWO5QYYPOmrAj/YEcLsiKB5qJ5VjByKG4jotEHA25GD
ZzWP+xKd3vIb6SGRiykha61/56E2p6gG72hCp80FnDjXAZO5jBZIhyz8mM76s7p9LLb7s2sd8+O1
hHbB1ltM7luDUT02IbArhm7P2ibjNIQNDuDm15DR2KrI1PMsWKx8KGkJebI16KtCU86ZrqBtYyjz
G6lPVPAAiEytemhiGAzQ9vIWrXBIP4tFlBDXWzPnqFKTp2ZByuWtKNHwcFCIqchEJFpccgqh55hn
r16g6CqCjFddCLR5BafZrwY1KF6V1o7Rfl+jBimjqTZMNhNhYMHP/U+pWuWjL/uuACCbqgprK4O2
967d3okBMBaGjjbRtlyZvY2Y9wBhnnG9D4uz4dXFrnQfNJUcsXwfRiy1SMvbGMvBTOmDBcOJGxv2
qUwIqg/CRR7jpN7RUGRI6xLgxnxKLNIhRG3SJph6wEUg0htOAm+t2jV+oljcLkojF5PuMrRIxsxT
5INHSaiU6IUor5rDfQE+rEUvVBgjrAtetzxmbveeEYOMEaWKKE/ES6m3Ne7m7/sLenuOtNqTbrXv
HakTb6XZqAzQb2Nsr2SZnrJZxJYMqu/y6zkRn+uW00NJ4xCcmP1WiWzyHY1DOCid9tDVnTgKmz1f
+7ITvj6eoETl3lj0lpiDrC9leoyIw8aI4AQ/6fthQBHd2EGVs4K/yPHK0S2tfS16eRgjksBWmqR5
Y4mTDQmUtlcwp5LIQ1DzZXKXT63yLEW/Fu9J9U0ngMvK6CynPQ+IkwklzCJy1UCAaxXgIwqbhW0b
yM9okzLEd58pHKqJOOvgwv9uWsGU+uzWgABVbpE1DR7TdA+99D3s5PvQsQshaI64Hig40gsuPo3V
NVgRnM0XUg8Ccju0g/xG+ljtniL+HkBINJJBPjFbaggY/pfJLWk2kESZa3bDNicxbfoEmxvQR4/r
JfGL+DyGnvi3OIjQYfuN5WFtOynl4h9dzMW4+RSot4GWFnhQ2dwR9iscd/pNPLTFRl/6S3+yyeTf
v/dv+TbYQrtlQXS0a82/sh6EmJEX98stIuh7WPW9YEnpwwfv3dvfCMnRxU6sB2x+AOvSZEeDU9wh
BmwRJ17KcWiZOG5suJBO+78RUdpzcdS2gKcvvE80eYRt73iGYKQmeZmqV8HA+mPEVp+mlad+CWhk
TLkLBAwmPcaSyjA5wpqSlQ6eWmBgwrekULnzjVGONZ5/GxtjxvnLMcfjoAvHEvuNvrVHOkxdMfp/
Qif22+OHNzlIc/m+94PTpvL7kwndaG4XYia45TOVssGUoSmeCFWcFIQZsxpPqzo+84Xpzp4HLBpI
FKEb6Ale97kmBvsfraqL+z6o3akvH4jVTM9h/X84kg6hYeVuwmlHgalk144avqKNSjyS9dMII5st
hSd3mBPCzpK61LyqQgF+0L1V4ndizxut0VSFNQ3GEH6EOYtJN9tsbfQtDZybryRaUJZCb/xtPCg5
s/d34eNVojLwKiHkMgDMd7Rmp9Hu3Rzvi2hLlbHLT6Bhxe/PTMr3+2SeYDRkY5xMccjIgG8r8oJw
xxjcQHG6A890AbHswWoQp6onzk3091svo9mMYufbRbCnuWNmyNzOWyGibmT/bWbjM142WNsfG/3M
1/WHzUhcP+nnqGix9vQtOGD7XC0zqi5Lhrq6IQLy1i0t6gGqhOyeie4MFL60G0ozDpbnkYEBBA42
4NWeiBhBjFRRatrrU+WMRsLqoTsTFSNEt2VvKjLLoPCVNuS6AvLMOsPTD90k8qGnqhcmcNWsALRx
1DsGgzl/uX53HPbJlmaypyxCtbLcomuOWjRKkHAE55YGpdnrufOewqLKZTvxU9ApBzWMS7ZLznZb
gdCcsIHSIQ8UB+NT6hCbsK3vBG/2LaXKcndBqWgrycksu/1Y4ymtSW8eKdLAXDFV6639+1TiKv0G
DZ62G9Y1ILXXhNTvpL0sRe3a8M4PQPLJqcLcg6ElyCLbwEa/9EMvLUR6cg7/m1pJbHWq9bh0Eke1
Vawlj6f6/I79St6EpycrJ1yBD3RDEWXTZZL4VdPV+ETMll80BpcxejBEI/m1e+D0XJhGfcAiFMlI
XhtaXis9Scubz3KJUbRvojLeD6eejVrjFjCMtSpLt9tpkolWL7VZwj/C1eUjPc0yTkzPpz3Qtp1j
vdC6BDxUryvPwcPY3foUhD8tPoMOXb5Fho9/ZdW9hYhXdsZdw3K3kJR2Ma/6Tlz2zUFRXsOfgqgf
WMTQ/iCu6To7pyCgaQAU+iHJWSC9MaSi6QFKcZkGEDcUgv2szX8jiUNDek3r/oROjFdcdsnw4Lsf
vtXS4NljiwvDgrury06Bg5uekrRXZYZGr/itffmpn1hftWfIJgPguY6fnkITZiIZRmMLgY7RibMt
eeh8KnYZtbjB7I+PONiExkSlevAFBMAT7r65f25sf8ypN1+aPHiGKIbAEaztD+5U04FGSEAPx5YJ
ORydW2TXuEdb2SZrYCPwzwTrzqGkyf2NH/A+FlayzTli8ktQ5hs6umiX1zIVuMIwyXw1/p+9t0Sl
NNZsL8lS/jWMziPOO2l/RJHtZyMKCla+QrTRf4/WghNREYZ7TVCFKA1TQEBuDpeBinvVfc3kJI3j
IzOB/c/+02DknlxRgk6v/9cRgxGLMnqnKFa8LgAbA/s3OYShqZ+Y0P+k/D93toBgDhO30NLLJXnL
jD2RsEnH1yq+WNbRnL+Hsu0Khs/7AyDbEmTMWfZu9HITov94q3/m+GcUQMeT6S3KCsIYvRuR4MqZ
1hPB/WkFEeR0AmkF6wKlcgo7rnUdf71hwsKRnVX4uR88rgsSM8cavh22N9DGcwjSmY1zbc1ioWtn
KCT7A01ri5O62hyv82rb6yv8fa7snOt3zy8OWZeQVAByt7Z5AMg7a4PXFq9ptyZK2jAxOZhyIEm5
cYhPwS/RjJRXTDPqx6TvhNU2YGpfc38MssTa0nUKlRGKKTcHrIOC/m+E1zqQ3T3C3KCHzCMy+h3W
nAZCqicOjUDPuzTRhVrdYtzQ6UHTM4+RyohjZvjE6iI1sApMyY/HO2MfUzD3ejX38JLSOrytmQ08
lmnwDUhYVrpNSYQIkv5JhteuZ4QwUcbPBSUO4/mIl09fH2Uhw8HQ247qSlrFYC1oiJCqes6sO6kH
lNr0dDAJcLrfJ6cLuIA6YIeOJ1mnjkmq0CdCZ6oKvr0eIIb2p46mAL9mH6Ullx8yHM6RZknmynly
3wkttnh//pStMyIuBtmPXM3awEyL1kCG+hIau7XW8lV0bABIzngF/EwPHqnrQy1zo6VUWoZ+ebMh
BRX/nE9+xhkOHfDGIOuzSxo2C0b2VFNOZ6s/KLWqbcuFuJM2vVTFbxpI0iEOo0DGcZ+LaXjDrfbd
r1/69hbC7vD0RVQ8w/jxCJYQsQxMRhvnSVPJnC9EJUjbjkAcsW2i6s/P2fZbhZ7mUYy+44cLLhVy
0Pl1985OroUwlFrh8+8WQK6v6u5Cdf3fkEg8lH1P4kS5ZyBJOq76isTR2GuLjMrjMCJ5D8GvgFRZ
MzIwgxgr3hXo3VunsImT/K2IEXaKk+TUNVtQRRS1W6fXCey+99ehjT4TOmHQdXfTGnrhDZKcPWNk
0aOAH8WbVYiudIrb2fIUrJ3T/Ot/xCWUDUrhXjYLrblBK44SPOnJupT0w3ppnEYVgH9oaaWTOrMy
r1hagl4CmibvEsItXeh+xc/XZ2RHZea04hH8cyU25DMmnuw3VjMH+xJx0rQBG2dsXQ5ImyRH0wHx
BoefSeqfU2eMlsf/4mFuQmQPYT55wvKAfY5iXbm48O5QHzpUbk9jI2s3CnKU35EpVwquwPz7vFIA
HsgxKsP7TXyR3koyAuQn9NMF0FGgO47HTBw9DB7tYTW7fj0dJSlPc6j1NHPZDC/Zixxpvr53gUjU
VFab5uX+IIggXQnZgZC3Qtn3gOidje5ComdKZfHazO4pm/T52Qx+sEle74sm1iSmXnNjA2bjjplk
p5bAzJQ4R1rUOwtytfOo8lyQGz9m3VKYbIj4Bu5oeW/J/xSiqyMIxUYIx+2C6QMWFPwEP2Mz8UQ1
0nazZNpBjKNid3voxii1Szlq/PsLATNey5hsy7Qb1ka8C4NJ4361bA8qJPKKDaDsHEcgdvGHuDJZ
YJ5dgW4zb2laD6NNcihpJlUFI5vSADdIJcwXMY7c+joJnHGlzdgptfcU804aJyZ15y+cesYlaWPw
grdXr7AjZUcRVNoKLWAZI5thjlp3fh81UbfJjTCviTFVzY6xVazobLBq5dNjKszeKE6QB9jjD5HL
/zKWuM0yoghGXo9kiCppbNaGF7xM1gyKMx7v+eHMlPq4CDWM3K4Z0BHzv11ULgex8NZ7HHV2TvEY
XeE+u1G+l7BgIX5F/nVN3vpgjbq2PJKs3pUSDXGbJAw7iZ5926+SmLuKzBB16Pkpo05QiZJTHIf4
Md+5Gs2jZ+mIAx+LUGfj2lpPbpF8YysDxHtSW7gdwD3dvXEjovoLCSUdQfkDI29s9QrFKwpM+g1U
ZMcqxWLC+74mf2hsYZ76Q6JfYFCQapgotVKA2LjLo4rPMWk3s49ei9qVe8dboKhFAoN9ielO8HEE
1MUL+OzipQJdytiWCnWU5yjVpZvq/sMFQv7w/IGvdt4woCdR1nmovOnyZN0JmnzSFaNxiiaEy78V
21/hjoFvk6M+2NiBiPop1JvixxpwXpTLurajiMUh5miLkpr/qAznfHnaXKiepUO+JXEpExVb40do
MiRQHwTNsaPHtIjHqTAWFdf2rTO1hC4GWYJ+dyMQsFuV03uABJMamoe9SnODDI7O044Xx04FMocn
APLknVtxOdcNcAPawe4+QY2m1nIctKhbbjL90VeO1otzJshQm+jIiJaMJyVyeE/MEildU65wjdGQ
jXOX2CbjduDcmtKES8A7UhPzO+dP+MCWXjxq33qpKdY2h9XBvB3Ysm1rdr3bOLitbGohlLRHf2is
XtFDT/DLYgfiQp4nuUVz/nEei5wLyVLKjmUmqAfdOjiKGkfWJHBDhdB9oJsIp6oUyYc/rkAnEUtJ
Wshj7Ds/OOJlVTqa+tE7R6yMFuDJwtTKge7xMqTWWyw8JStlmefPjRdf56xND4IVhwzgZey5Q4Vk
6/ztvbqG/w48GM2aMnca7DJ3bapNN/0k2yJC5TKmK4YWSRFswuYhh/SJDRo5mtIUKuH5HvnA3o9R
24rWB2IseIGV6f7c5DXGbufHeCCZX8ioXQ1JdjHDzm7bqkumNzAhV7CF3LFdr2UcD0woQ8rneR2k
Mh+uLaYZP5JXZyb+QA287uSRY7t7EpasmF2l9gY8PJlhXTB2fHK6lQSRHFuxVstb0qXxOezjiYJH
hmaBxYhtpW6KkGWD4ZcxBBhXcPxFRDZ0aw0TL2q7oTb0vOQ85fVnhaq4iAkaQk8kWX0pO4vrFQPU
W0sqIPUGJl0d9NsQH96heTnX9gjwbPGo9MxDzsUbMCSalz+/Su7OkAUAkfX8zBeN5XcGCHO6vjHS
sPq072iotWHMqAm0Gq0+7gBWtyZCkFurFKVyA2YiigbXAs/fGssc2kLlClU+Cq3+eDruA6ZuBWLJ
9L+5u4FLohFv++w4XjQQ6xKF2c6NDAKS28Zxj8OnlOSLACIpNb6OMPeTK/3X9DNNQlxtJA1J6dam
ZKDJXNrkOeVC7/SHumSxU7S4iO34mh4H5Fco3CoFlx1jD8hl+Y+TdbBxb8F/7P6ArrVI97DtPKkN
sQw6KPGsD94R6rv7dMy1c01Ayzy0EZOJ0gkdgOArQ03qtFeU1bSIGHXbE3cNCLClRZrfQH6bVzPH
baLGICjpNQWQ4rx7A0M43cvqV2l8kBPEwQTF4uatHsNJIR8YG+g3qf+h3mt9Nkq0pXD3Ms5+FkjO
blDy3+FnBqHnwMq7Fa4JAevZgjo2JEMJuZZoRH+U/7+5hmxKzLPLHT9fcue5TWBv7ZGOhk8EmeGx
xwUakRFD1fKE3bmCGcldLpPmUNNKvDhqVKTPA5rJfoUD/E5tC31tnE+AP3NzNniQHhC+42qYLyB/
Q+PHf9gcMMMn/X2/Va3g1sHi70nOZXJf8iL/ys5Z1CNALEoiLuQu/IGmMsLe89a6y/gEgLtlXZq7
fmbA2IbMm+k3tNo5EbQhA30F3rDd2xEyozskXq2tux8GOXsqtZOKLDdN6gG4UbWNnOE0w0TnnTRU
aP6YyqTEZhXw2jehqKoLyzkJzo+tADT7VMetOViReeceHe8WqRiLbZcOg406BGAgYxMqjsft1mOy
n6sO9NIaox8YG8XIDGeIlhiyvhlcmIVtjjizQrFkhW4JUn7SO5YYYP2fk9l/49qqH/SuGHUqhovv
txaSHWZhae1q2n42OX3if6oQ6if0UbY/VPU26L8nuNV7sHG7rzRvAzsj8vyzBOitVIQWd+3SEs2x
y5+dBwe6CD/xGyevrolVJFgW/uXlg0gMEg5bbrq7tfLEhgvqpXFvs5dc1JKoEMGPu11BM9RI7THt
Gsyvn3EiFI+jJLxHD99xpu6etFIHCiBG4hJe/+W02tokaVkpq/oki1PEaNcDPMr538wdIKU4LBGg
0g658VLNbQl7BZjsFF04onv/hvMayumQoPiHxi8qXJp7C3jrnWyRQWn5FG4JXVUc7LI0LRRWofub
CjgLO7yYEjzufIQDxE2igNQE+vTP/AnGl3z1TTfzzsPAODt0ZGMtl1m/xbaErbMnnyV/xhtsJIqv
vQNqzIjKeZNgtHt8t0bOjiYtXDpLxj9sqbrsDOA+YeqT+AopmVrjpG+iEfLL5sVjvXxWJuvQO7dD
eaB2lzHWXTIZCURkT2bzbVK8IlThgWfuEKsPwXUcv1EhcBZOE5BXWqeFUJMg2AmRfleL5xMwJvrD
mHaI/PSW43K29xd+hrE7ET+s/oCRPF9akzWZzNaW/frWqlkHhIU18dVjd3IV6BiegGgvgLVfviCp
qhgCv5pdd682ss2szC73btf/KyM7eamtOG3adfkoPn4KB0fZM19uMiCRsV4AYTqcYKlZHDU0OCYw
wNMd1xCGdlUT17sLS3gXp1MxQpDVkNkHVocdu5HmCkmZOLMnHgOa7ot4vLYtCuTfbyrWRsUBIIMd
Wj0SXNZjhvOpwUHvLSWdFuJpW3T0DkLQP4VdgoBZA+XYb7NqrinTBfX9dgmOxIcnDiZsP1Wijd7j
WcGQ03r5pPsCI3dyke+MCzx30F5XtTUsoP8E1nL8Zawed5fgS6aWL/RHNdX4MQ5JKrM8ZMfSIEU9
7MZbjRj7Fr6bEnVQkhRftoPzmxTRYLnjOrIk3mXXmgf4PJbe67x5bxETZ1qDMW/9W9sWclyp5ftO
UP2X5CCqpVyxPBxc6ZQBuMWEn14cavLu48OxkovJwOjcXJVeZYf4cZ7w3LI1YFLj13qcxesXbsh5
7VbcJiFX1g3gvu2NBb4oMukFzLjOIY5dYR5eYdpc9fExXPL1Hbw/1P+O9EbjM2GYGURDhekWxVpP
TI+WF8RqHxlX9jHwv8oCZ0Fq3+JcfA8uORiNvKQYA27AfTLxwIsKRUIE12GkdPHj6y02KcZw+ksj
kYNqs1/YVhkQnMY7kpa9bG2SxTigrWztOmIjLJJNmdx6uVrWKSmvhnYRen/JdB4eABDIjH8GetUQ
q5gtNSvpiZPe1OXbL6et26BFDNi/D2qSJU01j/P5/Kf30z43KWxSyJFP763JNjFxx0uXXcr3pefr
uzCNqtsEjPxZW7k1HxCwZZ2O/69Qnr/yt9FmBCTIZaF8Kizx6V+kLR4bY8h2jUoF96P+iyumv9Ec
mALX6W87efths1QBn1FlGodFd3jQ1Pw0bZQ1LyRMnZ7OV/HMqcxhVTZtBfP+YnFEBMguqmv9mvzz
H3hvr7xPNNddUXOg/pVaEI4NuHHf317PBJOFamEbjiKMEv8zD2OnsiT2Grjkv8heOHI/RefqMRTR
ZDGo895pkk/DdUhRe7Uubf2H5vVRNpQn1dPScxg1jhqbNpvMuX4TQVnhBfLKphw6eeVsHP1SePup
fvtrAZhvv/+Fz3mMzWIHHRa8ihP3CcoV7SaFf3YdlXTEemURbd9Q9KZ34rJT9Ci45bX+4B4Q2Ab2
Pmz6QswvH+VzE3Gp1D235LWMrv6zPlYcjCwcfI55VtKtdY2W1HubtOYoWIaWFGEPAtwwtP8KWu2u
MreIYAslc6VAdNDJIcAe3/vFVS3GJgpm9QHzAVMCSgyNljPBi3VJKJXMfWU6fnNpykN1sh0FsGwy
Zyb3JAOyXnOdIJH9wS8NrIMEQEoL1r/h5L1lVeLByl3ph/6k+ItciiGoWjN9k6ujoYtXUDkQ1zs2
EFbH0xxhBYaFd7n49sVw7XvIgr5vLhPYTGpq1YK7zkwf9yNwGTa3J/lHsR8NvsTbpv2FepVix2lC
JzDW4blNr63GUko+O4s3IMUHf0nGqP87vP1IUVZfM4XNwr28NzPzJfPEKb7yVDKRI99jemZOf7Si
bQDsjowoUxHvzGVXlyDEYO3HprRMbS0ZxT/bEG3c/G0ELrtfTnILi5MA27orZ4TS0bH8YlgOmgXG
0Owtfbx3UIpCMbnU+FPm/XWS7xzNLz33tlS5OS8mdZcDm9+xiddIUPWf8hcjeoewjyXtxtevfmT0
IBSArB2Gwb7Lm5sX5PzLtEQFNpZv7mgy8QtOWCFDE4TC74IcCF0pl9u0c3RvaeKdWUkCqEwh1yTU
j0JlDkEQkdrP9rUvc2i0ydpjLy+NPSFN1n+zwGINYkRVmb49t3kU77bNYDJSo9PZ2uPFq7iLsBC9
emz6DT/c/xHotur+zblVT9I3Hd1ojAX+nhpVyEZ+R383PVD6+wslKtsmanGWGrKWseeH4UVO8VMk
KcxA6VIyWYc21Sf86XpbSXrd0vswysm8hGv7O8b298VP4ZYeolthHNmNRpXuWH1H2gKf+fGo/J15
AajCpN8AZwWiZcjadb6W1ZlLkLBfxGTYZXVfm/6QH0MleL/JJkRBnoYarkfw8EottwRsBI7qNF8O
EaHPvAZPG7w4X/Q0lBbZWQRpgnJ+K2z6sAQbH3q68ciqDxCKK3eJfyZlB7B5hNFeOiGy36e1bZty
HL5L85HIZ0lrNErLiEVV3hU9f8fAifHhf2Jauex/yG5AzhqFN3qEwt6XCHFNiLxY1Ms+/jsnjJLd
gl4U8cOoCCbPwGRzWcs2JjXk6EKRGstibchQyT0k9OTM5fH/z3HOqBBqhfPt4D71UJ2uqragyrOJ
e464SEGoolEbPRDRdjdYizbYM7FEFuQkdbS/QCJ9A7tPl/6SlDSuNLcKBWg6fDc4DpuS5rAyI0qN
VTe99cfvueBncmO+i9PVygX4qBquIElnpemL2sJ+D3qP9phNSDKmDptOx58t9N06+gc6LPdDTcl0
ms/MfVIMhBLACcvrQLcVqduMZY2+WXWYLrmAklm0EZUwbI0xcsuHIWkqkn3FWO0HN4YQjd4GfUT9
Tnmdq4VDv4YqE3pns8C+diq2n3QJXgQdVOQlADyVsQMC/UH3xhXOeabtv2xqBSA2g5PnL/GhFM3I
4UA+xnh8eilIHvtd1xbNwICnct0XtUhzqO7nagv66HiIFO6nMQXbor/DeRMCMvxM6Kz+Hx8XbrzU
mcmlGKsUzyeVEjz+MYctP+qxrMOoW9CC/QHUz1D067/ept+45B09yT0F2aQdszVjDtOuvXoEvSkV
R8glEsEZXxNJ7VMPZm2MdvICGZH5C6P4dbU0QTEWhqvGRXGlC3f3oTV539AzmEy31Z4AIyVzGzpn
5X7+UAhgQ2FVd+wTAfbnxJJ2oyz7SCpDPPe2ysTQ642JO/tbSWI2lAdu2FHKgbXagLh2dj8ngfaY
jxB8WLMqqzLglRXAE/OvVhOPZB+/F+nI9TwQo8kcOHsOMdowB6fpGwrNs3l5ZHB+4im+no2+Yue5
si45dSI6wPcrUBUSULHcZo53UKqSA2Bjd8JNWSt7y/Nlu3HN1wKdbDhMEV5hagJFexkVe1X7d0t4
Hw6T7NQDUrVSRyAv9LEox/5riff2iZh2U8HtJv9lTkKx78eddFCaOpkuS2aXDUQBkXpP39WbIWVT
poJ/9TocfisM3QgPNJTsfLbDJKyxYT+Mjq6UhnD9P0Qi+/XuxN/seFZ7xK5EiKJUP0cuzrHqeNMl
iwczmRsX1Uk8p8HLgkmP1s97Ki1hheR5hM1lKCJcIZtilD6lQT7v5mm6bYHB+3JtKXb3pvyNYcZW
8YnUMr+IFJmGustk6DNW1CU9kaD5Flm9VWx5CEraQ4tjnarzCQQwSb28O1QNbpFxZb2MAiUKjbJU
X9SkFPDWLyTkaeZOQXTZLt8HrGC4SFt7qS/QFzK0zoGzgUiLfkcImyqCtFd1g1AsoLjATnSJFXy9
vek3WeVGriAM9/aBKx53Sy9umsboDRujUX9dv5JcS8UuMhgo+qDBRmA2qpi8JzeQ9CSWIy1FWxOf
PfAUogX3xmy+7+oUgLwjhYCMUIzCr6l/Ye7cd1zu52u0CP4x4KwBLY8ebY+xTKyg9HeTia9lYoQ/
s25SzoADqAqUMVKrVSCCMYia2NhvtKXjokXuuRU69AqdnmeE29q/eyjfUJSevJSaJTMjIv+IGKhf
w7laDB+jTqw0F3nCcQusvmu4OLBYjCMN0uZYJPeoFFGlpIGATYhmz9m/jDOGSR3LujRXJ2kePBX8
l5OK0KeBPnoQJ0GRxxKgAlVh+PAYuJ0lJbATcEXe/A21vcY75Bt1JBrKP2lKHSN3JXCEhzyOn69X
5JUzluTx95W7CGK+pTwVar/6ErpzHUvFvLfNNS3etEC1DGi/AAadfkRvzgwNwdGxvZijlUdlFwVb
M1kr/jBJnwyxFaJQtLpKdenLgCQJv/jeC6RCfxc3mySAM3wQmL2MkfvDSi9zpLmul6m4PIXDamVy
tgEx4gjH4ZYzKlmwFxEZvqFwdDX+/do/sN9sF7sGkiw8C6BI0h4eavU1KUOG05lU3ucvrL9bxaMU
U2SNc+wAUo4BMk1GERjADCtKoAwHuwJ7U1IXRSgnItxztrAyxna62UkeYAUgibTJh84AEpV6H79m
COu0/r7wgrBExG74dL0YZWBXLtX6S79yBrKsRkHWNw0VZFpr52l0CwHAiSFqi08WbtlGQQFhiSJS
6vrJdLYrcOU9qeG8zoIHqvaO9XnW3lZBk+jLp8tkgSow6tT/xWeSriVaziUhBRdCnCNlRUUVZIT7
MWmP9X4ZPz0AUNe90agAZ9cgZpQ6HJT1/qDPyQCq7p9eXKiSsVc51BeYuE8GlJuxs8tlwU5mK9BQ
fJLok+hUCVSrISK14Ewk65s7zpExZGaFQiG6T1LWAyHdhdTtyLiyVRZe+4Zrw3xLZ1VFbeyrOlfL
n0hEuGhv+5EVl18YCEeOBmxN+I+7ULhag+n7NyhRmSVFrzzS8ECFUviOf7ifd1ZM+Nb6T/9d4ax3
Da8ZLxe1k7gqi5VlNO/Cs3G1nLlpZP+89DlFNRcnZmLTo8kZWhnCQajLTTd2BinAoezp/BH2VfLI
klgOr5mK4BxDE6JVc7YPs62SKJIsjnHDQVS/R8KDq/fAr7S6oKak2VeBDZ8LboWkiOd9ArLNKzZp
anRSbmxaIlOxz6dHGqwDBo/ZhpK/wPlaVouwu0AFi+56l3rtrBmCBhG3h5ua7eT+gSumhktoXIJm
GWpJuPOny7nYPuK7dgPV4gSsV3YDn5qjASknQRwo5NxF2XltxQdBs7451Des5JRR9GNKMmU85Lp4
H9DGLfvPhqaTzjiMPMMjFf3wim0dfbi9ZMuU9wQ1IVVjJfPmJh8k7BXgG6XXKaBWiPGIKEEltW3s
23WYJM95UOGRVIejkFeePI1ZqT93mLkbKSdN07MBzbbRz5mmXVoUa78Sg101F08fDOqizPckpehH
nXsr2kamNhp2YpMAO89hS4Oh5TuAoabuyJffymiGuYpElALI4TgTLb0Wnt5tRdBDhr0iT4UDajjP
qpcr1GKyhrCs9BabLo+sTF9BwMCOFqOx7Mwyju3cXfyEHI5Qw0Wz3gCvlEYaIE3Gcvgnho0ikCsN
D3WO2jSRE8ZK1SkAXgHnNF53wh6dR4O1U1mmJZx1rIZRtB+cZPBWG61ctiLxzLDPTsSQZU4GjpU+
sthZ5aZqKZJm9i4eY9EXRpnkOBKyF9jryA8pWi2m/xlLNMSplDGXdm3tWFtyiOJZEkwBp4oOsG0R
+kvv5kryhkWRqy8/Nwg2Wb1obpb5gkWc4uGFzHdeLtDPWqAHhpzzKN8s98rjpSkH3UfVk6Zyr8A9
Kdtfgz5zy0xQq2gQSLb6AOWXyW6cXDDD6XYmWHxWoOP9VfyZ4SvcOpD9omb51AAIVrpy9yEu0h4e
KrfEE4Qpi/I8ZyUV0cj6bmGEzqNQ6HSWpaZ9AaGtOOg4GZltfaITm3GIRkBsAglZUu8MpzyqcMwZ
UEx/WglBxcU0eIP6L2lgiP9dsV3SFkHmHH4p0kXXYbKPNZ5eXybJVqRfVjmdwWQug44B4GZOrT3K
j8MytcSQvmAQ67CB0sG5BGmKuLCZTtiX4ZJovkeo0XUFphuXWsUF2wTbhydBVo3uRhik7XBOqLYS
cmC4g/8NFlQzakG+je8picVvtlmAjrcw7h+Go607Czp6+jSQzAXINHLZvMzAHQX6U/ffOQtCB50v
HYoph3s2ZRfVGbjeiBDUAffly5uvGoMLKq/yt+UEyahoChfV2/kk1u1I9okKDFG4FAEZv/0+YptB
N3+Y6Lcfk50rH4N8MYWed6yHLHbpCJtlzzSZRN0X5lBUswAwfa8LmRUVlF8KU58WTytp70A6HTJf
kvNjGpu+OfJF9ThOGGV7nf1Z4Nec83eQ4Jx7t+LcdMI6rnlHx6pxk+ityDP9b6V/jvqEFdZqd2oo
azkInXO/BjGTomY0LSM4Fn+NCg6xDm5c82DcYMrmzYXo5s04jkm4S8Hj6IM/EpF6OvzatanFCXco
LU50F++b9D9ssOTE4McPl29ApatdRay4uTiAP2IjQ6/hGjdRdD4TlrowOoBeGdp9S+xDYjpuGOJ+
obG3MoWLD3Hiz5EwGfRHhQmb798wSqfSjqf0RmyS8QtJde1p5ue/FJ6STjTnZOONIqNjhJw8vx2u
95UqiHvnFtVtK810nOBXT1P+af9ChEg/71jBPWDYvQQuah/5VCQVojoyYYiGI78o1R+Ge5RB/2Z4
DudvMzuYj7jiQVVgOhBBziaMeCmoUhohozZrPvFXNezZ6MYl7auhmkbxxEECOZHD3zZgOAPcMlYW
jZG/nbm1YGf7Ry2T561GFobWkAOouMoJZz/xXI/JPArnr+MRxL/YzScGaZLUgOAkL3RdDtYny9TM
cTW7hyPjIxvBrTvE5lb5uNmJ4W1II6kvmB8pCn0gjV16l6x9D+Mu6r2e41vA/BVu2P4N/8E49Wn4
tZZ6ANthr92o4p1ecX/cSX0g5JOWaHMEz6caO1O9KIPE9ZXnU6/1pfbZi8GnsSB/zgFYlEE8yveK
TXvPhiM2T2XCCloqyL/Tfy4ZBC/TiQ8CVUtdUx4DBzTFRiqGipBJgPM+JSLGXGMbudxWtCtkMXOG
C+8V/osDQ6RBxlwvi411ML4PJ0cJis0S1cwc769bzCxa8f4VpYz7an964pmkAjfQ9gibB8PJp2vT
2oA60aBXmSpGdP781MDRmOUN5I9GwcmjDxPrPYTGLrtBt0dBcCPq94IFvUJn7/JYU21UqkIwUh3w
MVnVUPbPD0NI1H5FkgDFp6lI7VwZEx2aJ/t4TFsLB5CPyrgDqrFGYAUIBJi/T3koBItX/lkBtapB
XPm/cWdNVmZZQDS1LVgsjRtp0W0POZEp9hg4fsGIBsq05I8HTDouSixjEUOeVPp9KbLzkk0vrPsO
k8S1OFzq8mNNHfLI32b91k9ovr10dWTEv7P+DCCIlFzIAm+0EeVwZaA5XTjqFlmJt07uOGfACmkg
R+D8VpRdf+tknWKaDC/iJVocQnv6ZGm80QSF7YNr35hyYm1MlSAto8jCOCAMfjjaGQ6G20HPGcme
TZdNJL4Bxpu30WDHbi42l5LhNAqbSMVHLlRJgu+vZByN/D6nwGpqNdFPT50XDetwmvW6XTe3Y1/s
9VA3VrA04ZBPEyePXRpEB6ICvjofcX4J6VgVPIAMvSpDjQPnclFQeyv3t10bmRHuMELo6JDUGxjU
VxX+C7xOUrKMxPQfUdVNBlxCWZxu/G+cK4GfbluNNG6yEQz7nFw8EPfkoRSwEI8i6XCRotux7/wc
Keoa/+2D81iHB3oICvDWGFjIKPV8jjAccJUVPSr8QNgAH2ikTRcA3EaRoZXdMFHEWbn9U0T0lUU5
s3scqsTfFr09McTTVFmD3IgKmriEIlg18BrO9TymYk0wMJh1cyjWO+/IAva4ccRTh7+Sw7SrB4Rt
TVsbldbU3wJE8QZO04yqpG/6QzsL++aa+qorbzfKGJaedyHNDZjTGJwG3bgEZdS9Cma4+Poahd1P
+KLH230V3ycNWPWK/WGQxOFTQmdy6aD82LpDo+ZMJfhM8FzX0dnjgdoWfDXwQFCQDQrAMarAVa4I
ac6LnuRxV39pSjtKbYA4jtCn7XGohgLTeyKJgb6HtD7F5Y3Dvj80KXULMHlPUIe19ZyK93Xrw51E
s+IuT6levbc0MguhjT3I576nvSYwdSQyAi9ZDixFPuaxvrVSWDqiNtP+YkDjHC5ja9ytVsYLoQXS
IbhnJPMkzVJHXcQzlG2s9+HgZaFUyC+JNHDYVLIcwl2IN96ZUgyr6BlR361ijskZVq+uXz5K0BKT
FCmynyw2ZdJQ8UzNBLu8s4dwwxSGc2HsDHiomSSwuY+z1S7ZRa9t5H5+0jAfXhEStl1DwqvjPgL1
XVbipWmfiuYqsYdQ1LVqFP2Y66NLxYqWDH/lAlN1yqsZGIs7YKE7H6qBLe6ta4plxSvU9sLKtseK
h6cvOj38+bAa6Mm6y81nGjlXF/VruYJOA59RaMSmxoSGv0muXFs9y0MUJgBIAmmA/aDn24zTkimg
YHNctKfBWC+mgd2Wvh8opGMLR3ChC5GJBplPJsQS4jXenBGHN98S9AURP0DRmvZIIfWGDf2N1X3z
hE3lvWvYuOmAdU74DnG+oOHu5H8mDJMtFlyB87jpdVQ8phK67b959PGO/Dak7/cQvt+q8vXAGgI8
lZcN5RW+WGMbR+vcwh2GLXxCcdNrr1oCgBS5sEt8Otx9j/nXK+/4N5ZCaTWAxFaPsiK9YsJnA3J1
7bGBvkRnDy1XceB/BMmGSJkoSF9R4yRCoEmqrlKCN7Lbm5DRgCINEPd2lIF48s4tzW7IleHlwAND
vhp0gfFIDcFDDtnEbm9KlSEa33m3SYwe9WQp2rvxntgK6VOZWSQCnVozjeIHj9gQl0YALJE8+liX
rNUevnZI4lRjlBclaYheSG2u5BJ/HYx3T3YiNTWvrt6Q+egMEEl++G1CGvGi78kOqCQmhEGDru81
FgNwQgeu6kFuNVXkJ18FvycPdgRaMf0qKq8Ob3qRRGbVrc4D95QCqubvLgeOBDcKmIaDevOiOQOW
TRQRxkyXBpLhjAe+d9gl5H08JFcg7uPLaTYV4p6M2/OQxdNSO+Yo4pbxncUCPtsJGetrmelsTeJa
ija3lxgbF+ib+Gbj6m+E/QpMXZSPDsYBIP5cDLaqRnj+s17C5R7Pwp8ABRx5xrkLQ9Hg5Lz34UX6
VKHrOew8ANWNfBY77Ua8GyGlWt9/OcIgmnz0oPq5FJCbqUA+mLMafqIo3kAx5v2WdA3CzHtUHqT+
NqDIqFcxFDDEDe8aQLlJdG9BmJr7VOXupSQm4yLM3STibGFiKs4p9SFjihkOeuDQlsUGrkFinNit
6Cet8Ugiz27Ja3iafu0gRZlvD84+4C2ubcVjTcB0vHHk+I3uGRp6EgwAtd1VZ6hD77o+skv7oz+T
TyEj2ZX6iicdtAvFSDRtfFwQ4vUDXViwAAazOJ8ap23wH+tU2qpcstyHvk8olB5IEw/AiNLvfC2H
/9HHODeFQXeDLe2wBiwG/obaNPWnmKJKTtoqyooot0urPC3BbeUDP9Z5XDbWbVyXLVwz0JRCidE3
ALOwIn6JuKRYMRBYMAE3s6IgDdafVUgPL2O6v/nmNDYZbzA4JurUlpj92nuRIog28uOoNTTuixAx
jIy3Rds6MT2Xcpvxox//mmfw4yieEmFcX+B9UiusjtXuTsNaQItAqTniSb5tvMXzKs9HYojCvlDK
6SkFowL9VMlmtXSdtB38HhRi78FoFs65eunJNG40zq/kQquNabvOGyeTeIhHpsAO59XN5VXC+m14
SoA7KtvjSvdLfWmb+BKTodgN/GIYr+qyJLOJlidNlp9mQWlVCXRyZuXv+F6U06dBwcK5Abjvo+6W
SXHlVld+wUFgD/9bmZ532vQEVK3vUmyD+QomXURcE+RTg26vpa4+BWG4u/9u0d4QExqGHO86Xv7y
4mw4Xkgf+gJFg7zviexfK1fXUwfabN8YCANoEnnKMqd5y7qmbl+R6xrF+2Ovtf6c7OIu72icfEhg
8gfb4iB+qNd+suYvs9373wLr67FHwHiNDMTS094EgpqxE5RB3vYmpe8Osycn433QkimQAff8fBui
0WdQNqhWP/D027lYo7fKE4yCsrURRkLxVCxysYT6Xa3NXBja9K0H6FlyGmLkxMHoAFQAgweRwY7z
heiWi2jFNXKeU6Hahal0UdCf7QkHnNQ/2T5VqQN5wzziCi3LjgZXalhlk2z3+YuW1ZrJH7QpDxsP
UE1KKG/c4WCKdR6iE6o4w5RuVwniZ7WeUHQhs9uHWQ4GRgFaToYTIJ3YxaRF5hnXDVnDKHZKu/uU
eg0bUdJjtV7ldacckjcH5XkAqI4keXRcklVWrWF8C4u7xFH6ufUb7qpb5NPLPOj7EFuCr9NYCE4X
yhyg103HGcwJutLRrSgERvuyMfRJV0YtAhj/EccN2cJRh3KrrPEswJgZfHIkxOx3RJBQhTplwCeL
8s1UKpqu4C1C4urRUdoSwInH/ldzPBUBEmLqv7V1zXB5OPdiqYjklHPU8oJR6bdU6+wLlccvayzn
Zcuot/ikzM36enhbhNu3Jen3JILkag0/xTS1A9wBKAOxzMxxcLmIHDPbPj3HdCMp7G6E9M5XVgPR
QhYmD6MsE7sOL70pVORA0+sbMQpOgzlJWC+Cjn6iscRiw4ul+vEgm6HgNtHk5qJsE2BvMC5zu47S
NHPx+tCl8CNaAEl18jVzRnFBe/uNlPiq7hFWAthS7s1o/Anzvc6XG/x9CvLO/YFlsT+biEdR+8Ft
YoFAAYggD0peG6s5KYke/nmU6xwFCY139KXG2AimBPGT6mI4AewBGKGK2098uFoJrro0u9soXXeH
76qIJBXRo1TPYgxv2FV5lJ/VTM0ZQoeTgLku4y0xBTG5Br4vFSBAzffmWNBQ8l0rFcdQdUTmVlPy
bt5IQKvBOvK0n0NiC1RJq5riR0rNUa1lQ+VLAGfjnNRVmg1iuswXoT5/LV+zzlyl+oFHVRzUd4BF
vy93fBStfflG7BbYv+MakKBqdONIc7aHpWEku7Z3bS1I7Si/KOwfxG/4Jb38c3TWMUlr9kX+0r14
M+1fFS+3ETAIQJ/XwS9Rgs0XFhvp2PHZJ/xUhLVuSdS0neuSdIVAgetRqkqL5d89u9nbfzsIHCCn
pV4HddUzPab9udmUFIAJIg/qB5lm/SZ9olxFwpubPbzd/2yrqY/ftL5shoguxsp0NFRgfdw+AIm0
1Bn2tZIiIOVsZn7mzPtFlr1l+aoYtoaSSYWHQL9pM18h+5GQMhgbVdlS4i9tG9r3C1SOEqaQPu9Q
XWeEiC6SaiGCpRE2i2nqV+xWsYy8HVvWDV3Zf4o6p9J+A0stQSTDEsXN1UoLq/6HUG7azR1lkZdb
VLsmV+hBwiMjXjRcp8rgDYzaI7UYOqPKRp/Hh8g7DtunCGcgfIOoNaxKjwMiAoFW+GOOgOv+A37n
S2NEzVlzgCRf6Edu+ToPJR1w2Pulc5wJQ0wqKZ4GLV2WyyN4bNvIOTn5hoN2kuRF0FTHYPl0NWSP
ziOqUuo5LQcYgYA8vgxeoMgKuxda3k/agK6nWdQoZwuDOnWeRzyUBF04pMMFDbkGhioZQw80y/0y
/INPr0QARd0O8BIIc7AsVRq6p1/USIA/ypXzDi9PTSE7NbnlWS+AhPQYO/Y41psNC6frzkkiWHNH
Syi8mc1KVl6mxV6HDDX9NIA0YadyIcTnDpi+L2eu1hkMV99P2mKcIp2NRLQSl1H2YYjnfFl0E8J3
jZDfmwQpHKGLG5xJbS4xY/Ypg8EQwhag0sN2xcR6hfoAENGHhd+2UG0F+zeYfw7LqPIuKDoFgFeZ
pCyJfLzSbzYPq8SQIAZDQMoa/fOdIv30TcAoR7QOlXNHzglgYy787dboOQ6pODNIzDt5Vfb2t/4h
YCMDBIKiSqWNMQ5y4WeUF04GZsXNzfAoQyq37qRv3RWoyHhjOlgD6Uz/EkQozx6/xf9nXpf3q8oH
PfYTwR3EnZQ4D6OHb4UwMfpZnBCOwisrmKXyOsfo5G0Wp3pME5UI7HmrypL6FVRXM9FKu7z+SWVd
biTmA9/geS0ca0pnz60Jd3icPDBviNaKVLi3jpFuV6GGI8/MD19d1BTw5i7VJiPucu/5BV4VWDnc
xJ7988NgfpxcnIWcAzZwnOMIdG/4dhLMkQssgEhIzWjqg2HOWiyHqeDr0L1XCfTSQkmd5XmdnpY9
QtCFmTe7mM11SLODmGrWoVYAOuvvWKZGwTbkrzX7Fd9M/lf2QR/MPr9RKNS0HU8VhPx2UR8Hng9r
gSKXyF5aNdQciFpabWMUmTnSN6VjfT+Gv79w31RtDPT/X8lNVkoNViu3OCKaQpY8Ttl6It6KcZiL
M4zIlb57egwm+ESHjJLdEmo7i1clHeWhQE15/3PMebF8mjBkW3IXhWZkJXaCsXAEOmHt7cg7MK1F
/VN7tMRfbVjwPiPRDiqeBfhWQpqv9l9vEEohqdSlumw1S6mko2Ez+rzUDt0Zww7LwPgdIrl9LjYs
KRS4J7L7UMB4iCL1F0hTLR60CdByqeaZnscMt2tayJXGcmg7X865TshkIapbXbf+CY6j5oA7jm78
u9dBg/oauXYKJRH1xe12cfa/OA8L4+c/4lez8wyeFxVkZe95JBrXktmE3EoHcC47xYpiLySubx13
zYRtIa/q6VrTS5OemsYdN5YSWD4gUyxHVmhf7sRZbcnN4Sodi+Ed5ccIZ5OQblL+eWVu322oY48l
0fslXm17pR+/Gl6Tos6tgGPW4QNbZk2FrDZlxjRAzgkRaxFDOS+FhRHOZatX4wd6o5c7hSpQKrsf
U/dxkwiVkPvOEEejuu1pKyAnhoURpS7O+1S7LpACL0HK/hv7AhvCagKLyXVt1p6DedOgGBIfUdnC
zqajH6qS54WlsZ5XYdUQFPdPky80AwtV4O6PVDXF7869CowAc77raE274Z6LSbL8TVnhshpPMPtJ
bn5iRO8eI4Da4pgM7yMqm6Bexl3iYEKo8VdcW5SoR26E/fC6hLX5ewoylqwv9ZLjEMy6NRpI7JKl
Q1W3PSn7oZd5v3YrqeSWehkK4X8XdIPBRYG612lzl+pZ/IT+6Ev2ingSP3RYlYeNAE5gBdR51Dqz
VSs+8APvQZNgYJuTMsqIcNU0S5fhLqzf/ZLkbmMRuS/y0Jnv16SjM/AL7YiGm539m2p/aI92IV8n
pq/jkDBnLPNEn/X8dGANyoDgw/lqzCnE5/Hv40MOFEn1xI+wmF4rZTaDITlIbx2GTMHcQvYP3GrT
ywin+Y44TYUbVgprtxUcksj45TQpqMHoQJXiVxSxir4iZJdQFMQpt7rBH+qMsa7bq4NRizKGGWLi
r/puWViAMeYGZT9ig62+cmyOLQCk2jZHVFTjaGJmJBUJx25xhkdWnFW3pDU/L5xJh9CgmHSlUZHw
eD0f8uSOcDMkMHFlZ3RRf08i7S9lh/CWlMdq10aLpfblzHJzS8lXnQ86/ueHTswQsummwy+K/R9/
Jzqs+iDCwfPy7hXAfPvg3P1D2tlIXcaCu56a08Fw8HMP0nh+RoTlTA5W1VwZeR+xiyoKVHtRr8mn
wR9fGwY+I29yooLKhM4e7KiWufXP7yBDEoOHvEZ24ejiQWbML4UWrX+9n48leAGhtAv978l2Z3qT
TPTi/xdAOvgE4i6WKe0M5IZLG2uZo/G10ECsYMZ9yjhu9cUaQd9y7SHcbQFMjLyICc+36SNEKAkn
KdmReFDptBNJaC61Bujjj7pbn3pt1EHr3SPH44zjNvx1kSjApFFPi/gNp/DkZvFGhN1SGE/XsBV0
hxx+N48TU6Ckcp8WHxdx88Xb03uZkXJ/qdTMBZMA1GQgpDqr1z81E3dXR0PAyv4nutLQEiS3QE3Y
aHw/glHi8l9k8slsA3Y2mXG2ZqcOJw/K9kYVD8+M99wwMkcdDJGRQ7/Kc4x6wDIS+cvFQA/qOH0T
/aPqwBhd3LgrnAIeAmXumZhyFciRkIvYv+4/wZEqkMedrb/+Dy+pwXxa4P/Cr3gUUZly5ZQfTiN3
0jwPTzf5CS5y/gYgOY4SOw/2Pcdv+qNbAuDg0xy/HNi1AzgeODKBqJDDr8m5zTDrtscEJvyBbY4j
s7VKH9mhhGyTLBdDfOGO3K0wCPfJbrYcJ2J0jn1zQLIGsxey/XAEalRJfaH2z9T0aj7vjIWeF4Pz
la91vWFnBhpC4Unijbz1fwmY1pyHugVAi/yEg41vBL4PXYacSn66t1GnSuAvCQYjadKYC1prsh8y
mSugZ1Dk0F1q99b7K1eai2wrVCmNWY3U1JEp33aqXX57dteUYD3FkSs2hoAcm63rUFZ1lDRAPu9o
0YiANbPXf8btD/lPWr8WFIEDMHLSQG7l3iy2DM6eTKtrLeMO95dSd1anTNqwdM+NHqPKnDqrqpT4
R3+ibWIt+Ejl/NZC7vBBYOsQNAl1GXL9D6EeMMqM6FA4rZ2jXkYluCJ3ZB0J2XbjFaIPu+PRE9iW
2kYhJdJlpbGm5wWvsApzzhlE6CnKC82bUakQ6XElMCs4i5FG0F5/ozLOdOq+ogQsxtaDbRTj1YpY
7SGgRr5Df+A9aWFhYZWP5YkBv5tjVjDL5HHH8x2pg0a475zgFYJ7vn4rwMTWz7/YvjGpmYhExlnP
vSYy9S5TlQHDbYJ3a0W6e9iGul81m4SZurbg/zqLLAvdHLEvLxc+4OiY4ER78r36wV7olwOM7Ftj
bpun5qeLdmecZaYiJgazdIP1SilNm1aTlosgLPQTK3aKL8c0c9oHTZmPc/unCwsc0WraNwHh04rI
oypkroJHY504UY3Fcm+B0DlKReBduT3vUeUS0EEmUWmlu2xpPBiNBekywByqtSM8DEvH6gDC/PI/
Tvkf7VMR2JAZVip9JJLCb8PYLWg/2yYi5C9hptDSBEja9wlB97/RK1ZlEcoyWjKYKJKH2pntDMwN
4Vv4q3/9/7l1YbmEh09BuGKINqvjdQoeTCo9G9wGZMsia0Y6ub+FvE1yYWLMSzk3pqAzRrlaGEBW
6EtZojkwBaTph0/iQR2LuNDnWn1IGN+4aN2URjrYC5Fhz4kI44sOa2s+iUwlnHDPnS2m4QyJW2CN
y+ZEoVntv95FVkgqdMvdFdL6r2rKApG3NTvhTg9A3ThGMMP6BjYJB5d3VnWR+Z4jwU5c3u3HNG6H
IEhad0WaiDcAceDKXL8QM6O9HAyE+wC9sET7zMH+dNXbMHn9R6OUBbZbNYqJ1U4w+xZbhXUiaBnt
CZaRL2kLsPv2+ddqK8PX5QYogtKfjsTL6y+j9to1BwHZCLrnJq9D9Xo7x5Yvu2T60veh+2rsXR4K
RjUffHS2zzhfQIeejJxX8vEg5knZkllF4Yf73JoOcnwoqYjutUinxEy8Aa42Lym8Hrfdd+zCO1IY
PqHMvgFunLZO1ej5DdkOYZsFTl7WPG/rv0BqIMiXRcJssTm0KkrO2fkKFJdbnLOjUsdV9zmGV+Ag
UcVqvfPZuKoevTsbjlseDKU8tEyKVezWWnFwA1vYt10onZ9+KNY8mmZDKp4BWlvX1FdSjQNvPWAc
lsiCscFLvadkKXsDAlPtQCPN0hyOoTpEXhPADJqvpH1+MYMtcsjycTdCGLlSiW1CglEdvmoVOVGL
cs46GshyXmw5X9F6ziKSAkUxFfaRJGuhvvkvmkef08kVg4CgaDgtqurWOd39m8dtzk1XYx1jj49u
N6YWzHTP7sIu5i8jd5RfoLVRIgempqHtBF8t2G7/kZmkPuVsCnbn/knfHD+ljf6xj3lHhMwQaot6
Wijx+DdCrj4dn1p+tZbAnNGbeBW9xYwoIXZxl+eLp9LIqYXVBp67jDjVZBkj7q3BQx11t+CAGlSJ
uzFKPEhQvqjCag1DjJ1Y6AuJqFN3Iek+bXSdUhw5NaGRjqMiyT5KfLEi/+RafB2+10ZPNUDineA5
S6HCBugimrovYUkUQRUaZMzD/Up6iD7AaG0k/Pjl1tM+SvQ0yBONwanAwbGrG0hEl2PD7dSrJzV6
QKDJx+JkjYlsSXtOLvXn6j/x2Lb58Twfn7EYsg8R3MwnC6J7HKaD05/h+5WPoPdxYibCkTeknapD
1m9Kij2lcpsoHO8T+hnkSa5iWdgKyWs9a2UzIfFflAVCGVKI/i98FczLmK7BSa2rXEkXMo5H9sMn
UT2TJORbrNU1nQdS3IWzqRFAEdHPAb4+0S29MCesBaP1yzbNeI3cGRbRL1WGmLLA50NzrPCdIhnZ
7GDoXmjDDQuT2Db/trC+BqlSJHXSNg66rEagsuBJ9WNTMxPewoqpPbeU2qNgj5qPtCocm0QxijKZ
PXg+tHqmZ95Pi0gfsOBRfBDKYXIMN59DgfkfEQ5zWhnXbhp3TxpJ4PIRT4gUxUR4fUJDLLeWJWh0
VoAz0kLiJ6I22O0Nem472RtfmVuLrG0AyRSJe73YssfqH1NFKsoQ8XV3Iv/XQF0r+88d5kxS4qJK
SSNNjNfTWvUvB2ZclV0D0nhufxMia5VHIqgK6pn3pCBSvhT9MkxtueJQVlGTi5kYuoxve2+tGpTY
Oy2iv7SgO5XUX/w6/HrosvWysoyNqfbOFoe1qdsDtPkz/hMLyzfJsOBrR0v7LMngsAvWRgjB47Ol
s0iCjlt8SsEpiUwmNJIndpzxMP2SxW4nhoHvM1hgulz3s46huRZI2h4Wbo6QtVEOBCr0y9+SrWco
iJa6pp71FjoRJDF4NANHwlV/GfkitB0p/fmPwSaDXEm42mI5GXfrVq/NZjjWjQiI1wzrLYmAmWD+
R8vLL+gkp8H25rC/pLspjYARILrbeXxKukDTuS/QySxnAWGWGuSz7Btiz4IFKALhEjfl+YWjAGu8
90w2uMMJYU33TtpigPQSVD6ekSjeRPt/nH04hO56JCWISUOSlNLGNPrJZbRHcfhEJeaCbah/lI2N
SRStFObbS4tIUx6Gi5LLRcJzuvkukHv7c3Gol9l5o8z17vWNnrUc0K4xGS9ABHmWgwRwXPiKeahh
P0SZIqv5c6dqB1XnR3DcCTgriv59ZYJ+MDjPWxHwYT+/Y2CQGiP6mwzWP27ccRzthMeygr6Bidzi
TihQPNb+Z7l6PJA9bDxdUSZEJlcj0OqbLfrA2XN3a5VXOmIrvLXTLx45cOhcnaX7FndskNmkH+zP
naST6PF4UKOLk7fKMUhhMZXoJP8+GoQ7b0BOktQA7OPCeE+btusX6Zae2qgAzJXTg1YRkTEnlC3s
23fip7AaNWhC9q2Mv/Ua6qd7bYqN+7JiL4+GKEqviSuWYP1E/TngmlAULbGgRlSflMJi+5xXqH6j
2Blv+ya5mb0y2BLIQdm7W1xsydkbl6/jNyu/WOi4PSPTt+mGjH0mJ9Jvplbt/xb4vTJhWi3mai1z
Q/W/izbOAb1ro2oFPGaKlp9DrAClrSoxSZuH8O1cWLwDvVOTU2p9IBdPz4jukj2jrT5hMgZ3/iyV
UmP9+0GY9r29pTiuiQ67VWHp5enbmpkosQs59QnjbnndOD5xURAyybiX49OYGqlZygKNbpW/7TSW
UVNocZ0o0JZYiwzYnwPmN6l11hF9IytixhzGOG2RumOVk+3Bxq6iZ+bfqG0cg2gNZSv5dXsTy7fr
bhvSDGanzIp5rukKSBZ9JdFmBaHaMzfG5jkzoZ28kP4Y6UBfy+zyoBVui2ExhubYlGXJDLFvFNQU
xFJNbi5HswKzKu1+EPoA6X2seczAWz0c6iZWfse7OTwmcVpgj9BoxviWxh9txpUN3n3Hhz7rmWDy
MJcxJeg7beJdwXuvUzo7dQj6LpwxSsPoiTpCcXiEjsDNuquD4DmoEcwq06njgGzesDKEv/KVEq6Z
BWxhHApMUnA/dFw1jHn5cHaKjX5n1rjB3pcQR6UqCQB2gygQduVxU5jcLi8wlkpJH+eUvKyVhTFu
IuMdLcu1yC4F0hZG26iE7u70foln+2GSe9x+1Ee5B4mR+7sN4615VCklMliP754J68uYW2mbVoTa
jGSTYNjlUNgmffWZWijgcoawI/AitIolFLVhua4p7Ous0YNSgeJFjOE21BYmcruBRAGYMMUwmHXa
T7Vy9Ej55+zVaLuYrGKVO9aqOJB9LOXknE+1tVgryk/f4dv4XfUDRkdVqgiQ25Eqja8MHtWtRX04
Nuumo6U2eml8s6hmVD/R3cF2W/mLpm/0tOpArYyzZGkZjwe0ylBZ/SUtliU+pWUnU13oFG9Iw9n/
0+Cj92pYhcvU3UNsQVaIG15yA5COWSdDFTQiCjXc/EAD+rJSPD4OSeiTJ7oaOnTX62osZos/Gu1A
3QjhocXM+pl/Tc3eLvut1L33kDinWytvOw99LsEuP1WShGePCFcgVypmTWKoMTptIgvA37tupq93
MP7evW+STGLbhxGVS8xqwvdMbrV63gujLRWvznhflqfXU47YP59cHTzfk1mwFeSqvOxLn3vIAkZf
utiCQtT2UBaaUEmpMzV0rjEILWFXRE3lnJ8hOo1xcEZj9PFv0fMy0ElT0F6z5O6FyDbfI0p5Wk+j
gnVr0TfbxbRKGGv40rSTomCIEDlD+9aFNS69ROuCH4sCmmADn2CMu7BBtJcD+dcv+UPSvY9f+kth
agUDYPVs3VWI93PpcLo7RRg2SdSSMWQQGbCL1lQOM5+ibUJGsSUvW7E4Jin1m7UZY4hxoUX4xZGH
ZFDPPZ8g2sc7LlNrweult1oqfa73wG/3JrnO1kQxRNIj41MgOVA3Z7PXQb6LYepRg+kpCcSDLRVT
EiFm07fNdpQweZUFhFL0pl9nF0QFF+cdzCR0O+Fv2RqgltIxrANsNCYUCjfP9nswwJwHfXCYInQu
VjZVhEemoun0kwnhhxPmvx7m8Z/zuAcRVTZLEa+tlnkCpIWrYAzRYkBWKFZPBemQX62c+irV12Qo
EUxbbS5/rBvH6g9Z/c8XKSrM2zDg5uuxUeJ2Xa4+9JAef6M9oFdPz4R4Ufzobd5NWmd1BjSvtEFf
p/OH09svPgtTpe37t8A8yDssdNs6iUTfM/T+vtOZGXKffGEJ91cauBmDRK/XzhwZloSuZkLuX/yT
6wRcSTQAM5T+hlGZYvoDOhYwb5Pdo+VAfdU2bLxUtTRSWyBs4KtCFHeUtUpKkVEJtQCTn28JsWS2
+RKxYtiM3r6PSghGlWA6fC+1anyKXwl5CUh91PCGVvhzWVXrh4RFkPhYd9B8STLhJh6XkHQxKxqL
xumTdTs0MqXl5X4B5uLhqw7vO1a3evQrf7IW/L4NOQKKRpvvWJ5LjgC6igIQDoDfl1zEnDZBS/To
yqm0oDlDWudOFGy1aKKVcfrvXGImmwlsuY1sp3HGfj13BbfZjDdzigDY6N/vnoOcGZ+xFKLfgxSq
l4mKcuxBJOxto1PfFM62nh/z5QAFpxCgfxmEwd4CbCiBsfUNoaT9uusno59NXXny6SM5h8o3w4vX
hdf4p49W+Z+HFich6OZwlyEF8fFc1e9cG8HJYZV9cnk62cUiScrBgvLK+GSDuDUUH1iwG7SQuxWX
5aHRPwleNWstNccFGHlEXDt5Jo/A0lc+jIY0cjxznILErbWaa3K9dw/VQNbFdmLn+0gJlVipmJRK
YYrKM+06IDzjvlT0RUIEv1G7Qzq77IGyarhxsazkgUyyVExX85y/c9MQv8Ajzl/kDfbayb7S3Ji0
mOicRzfyc8+UAzYqtXH7qG4BV1qSP4qS62DYxomqBhVCwrFSEygXtvb8oQHp6kYDUXV3cFWBclHP
k3LGhRrSRz3zwzcvU55cMQJMxaDnVCX+VxRux3jNm+Df4U/r+2nQeyjKq0FLUfItdXTU8ssWSTcH
l8NdUjTgPoyjCBEfx7tCoqc4DaFyemLSImQoErRVR7Fpi/oad8Z48imiT09qp509sUeVo4kymgrA
9DNAnpF2ooISZBajxM0iKZX/YW6yvZJ6cwZidmFkJ/5q6tx8kNDQToRvaqWUeSvOOzOXVzxjgvMp
0gggOE4AXeZZLxLv8x6gEWJNqOnYgcUEZK1i7yhqEBvM1UWzLk3x+K3ghMhTRuHXNy6pyUO5NHuV
W6a3qsdAc0OgqD4DNtjruIAdsQGCtq5NlLgWEhl13QrFypqjec3XY/3R1mSIPbwuvpyxExkHqPTU
n2A3LeJgzTPgPDsNZhRkkQWZwjRhrFi0VQCDNCVQs6T08jJ6/3g3ndo49wLdL2Y07/6Iw3z42ZT3
5+vZDUM17o9Sv7c5YH5Abws9O6cMt1voMKf/KyWIP2gUVhBNF7sna58klDF3gh8Cv0v7Rq/zDqv1
YdoT+k9P/NVidyxCBxkBPGxyqgjazv/n33oNWTzQJgcQ/l3vhrWtpuhj9oCJpe+MxkmvSDIYso2n
gM/JSw4DoklcDCwPjBXiQPYUw4gKpl2VdxdET7EAjl1/WBfGEbZBNLAHEz41Rmn0Pg2aMzTJHmYZ
qiMFlxUmngZRdaI643n6xgbMd8PsZ31AWwZw+21WpYpHqJ56vWMfXVaINdBf4mHEFikL6LuQUTZv
QAAM8feHJ3iuf+s14YC796XuqshwSJTp0n9o73ej2ayVjbf3iMB0xcm+VZyxEOFOhBCImw3dHJzA
Bo5kxgnaYAgny+KWv3cN+Ck7BgeqXnrQclXaoo9TPUpYY08+Y9Yms00cxpbpRi0B2ZFUfKc2U54O
/si6BPDOlnXiGYbhr+bPDL7Ie0jH1PCnGBoOOKV/2prIvxrWwZcUESX6qT6Bzq2y+yoepjw17M15
giUTcWdyiFwiV5bq21cXUFeoyWsruMIEQ+nUvHjxYMVHyzPh4vzTXRh6yKTThguEz92FQNsOi/M3
ILqN3wCRRHjcSn5Rf8S/P0NDs0lq7JSeGQ/vuhauQTv/Ke/l4CeBhaDBLrG3NJu6LkQ2b1EE25ST
u9CFMWCoPOssBHdWgAsbnSsDw9VsgbXR6FCNTCUnJ+G2H+6yg0KcHbHX2rS5SOuWkDHuIEV50FsK
h6VrvJ7vhPKPyEQlX3VM/TXXmJOVG1+sJtJQZAzabk0HdwnPbTHQ7njs2pDW0DXgcb1s+jtWrZET
5EH7M+Oxf/8n9LX/l8I6kO5BQXUZE1qXIop9jt+PELsj2Y3sYewE29lXlzEBKQaYGX/OnpLIPxUZ
tqyNRXWO9fOZzAPRpLLFYfiPydFjqDboNgt833tXlQ5Gq07R3f7bAUdZmOZYWU1Vzao7kz7xpvPD
n9KFUYGnPP0d7wQ0WMToklSiOuK9LTLlqfBdqqAvLxk/a3P4oPM+I7MCSI7o4HTsUriAhFWJPjTC
etXh+L7YJIVRc/+REDa0S4z41btEC2nWhK3sOYFaWm7yGtk9mScmMRpCvgFnj/FJdZBHiCOYQLVj
Ha9Ei4eeywddVrAFiYek0Ob9VA+1v5GqxOsjCgHgASWJzWRyLRKEJUpGkuRCPOmOaYCRE46GyA4I
k/VauP/ILh7KmFIgcU3lK6J29KWA307wGeel0tv8sp+9nFgftYszOpPxJJoOtd1JhbNgnF+pOM7k
N77lc1IvaTN30IUr1w+jmZytaGk0yeViL84vpXSBV+mXCL5au78pV1biQfNShtDwgLNh4SJPjOvh
Je6w1dUGse409rtq97i0bzmlm6pqh3/2OBHBvlltJrt0AOQeOM3S2PyXbzg0+3zL3DH6SLMcPNRb
rwZtH9LUYAb82OR/DSJ6FJzDVr1yR7pHyp3AGS1VwvzE5Xpaev0i6nMONYh1c1pJ3m3QEAS+D0+5
mPeCIqNEEjH9QIyGvWdTdM0N+mg18qPExWYvRy0Pi6T9H9Rrvsiccz3/I3/ZnEhohFt6wXevt0A5
oLG+6vUE9Ih3v04SNmGCem5e0MsrK6UXhWt821iZ9KSxVkfu+vTEwI19GZVLeeZgnSRVkxmMUKY1
Lsyx2A0fw/iWC/+Y/ruiEjqrvABwjZJMM43n6FrU1Mvn/TtpUjZD+vk6NwacrY0nPmmAXOrwwMZ5
GIq796Jp5lgnXVz2hMbAuVYefQaLwoqhBWkXf6T4j1ntLgQiLpcihP9t4HuPestsmceMS49zcd9P
i+pk9wjhbo00wggExDcPyOa+OAuXLpMTm9Cbg8xvx1U2YySX4ic0ZdsDVg4zTDKWnsfwQLcWGEbs
+gjfaQs5LEjPE3j5uIL4467FLql0YrJmSQSGtdPVv/z79UL7yoMjQ3LjcpRFvb7ER4A9S5ZOwYCO
4D4WvW6S42GC5uecHFiuk2+LefjWpxtGCHdvufYa5bfsa3Vdk3K6a6K33qViWAJF7mW8+fdt6VbV
RJPHea6t8pUMYe7O8opg5FqII3PTr6lw5PPOxeaMc6QSku4Y2t7vK6rsjCoGk+s5UNA+jz50TUH8
DBkZ3SEALJX7OkUU3MY7InkhXC4YXII2wLp9Vc2MWis0nKfj/gkC0KFsQz/0gHY/cj3eKgwf+IeN
uZ21h1qqMkbPtmGWIb2EwGNkp9guWe/HBDGUSwdJXKVpIWJ+xRyUqDhkAQrvA9ulovmzKk3irjjh
oHKvHqHF97sspBDgtub5hEBynuVpN/4iU6KOsn7tvqriYwxkzMqNz1to2T5H+9UPvSJgqJF1jfbQ
ZxNybhYFSafTQkLfVLNLPzRfwVGM95RICdQUeYu0yEWbgsDuPdnwVK5etU/rEa+N+6Rb6pKHnrMO
f6zcF0soWN+9QzQtcRujT+uXgxo4LdJcbS6XvPnzqPO60/nHbNUrJE8vputXIbsyD9h6Hqq+aBpM
JJy4KZqwOncE3dovF/oNAMDvTfXg+6XdxRp5S54wtNNVIPeibzmqv21Yhianxo82yYGjGpAO1JGX
cqkQWFkYjd9YKfOjTx6YLVlauWVcuvdBH/ErVg6Tus8s9tSdPfO30VPhXtlhAVJrY7nfI2K6qWuz
Wc3TDGUEnwdTg1ps1fkt8wAOv0DtqHoXKtsLidv+8vocRE8Ya7nouXKBOwVR/3CQbPx3tn9EuV7t
c4l23Z0u1HoV9oQpBnDFMDfgKvT3eF8U/TZ6JG+NxCOfEAQSZzJl2Mq7wHPoFlHpF5/q58n7GpcE
pOyPuRRACp1W2mP6h7BRoLle25SsV8IJ6VnwXmKZ6xylylNwFi+6+D89hxQ2lohJqq7gRnLdv/2j
kpLe6uTdG6cU86fdz7Bp2fYxBHZlJiVOvNx4YY8v/Ryx2G4Htf2+GHR4do2zf+uTxs3LjW8ahiww
GwfZfguiUEnkarviqNWSFf8KjbA7J2MpM89iqez6Q/tL6lETkLXkt7UyGJe9t1r6RcJiuEpOZ8fg
TcxqBfpqi5Ib5qH7gNHjDLGNfByZtf56BwDUzF4DO2zU6WwxP9ctN0V9Z24KUkD7llbws9N62BYN
HrUbcEyqDj76nd1PiT165aodNWqtNL9tsq5LjrSVFEbXuJc7iYYGjuixcQUxvN6jdjv3KYfjL9ok
TPB+vVpYkZMEzJFSUCO1eBlFwSauZqccYwWfWOa2OrKW5y33dteuC5Lq7ym6aCgzSQYYuEz+q9pF
W0HJPhYSt8K2zT8RHK3t5JIInE6VA0GG8aTJ6wdQhUZ8VlrWpCkhcz95Q+y4NDWUVJzjGVADIzSa
lVn6CAOrWKLRDdhUgyAzPuDzsE5WoaCzEKbK/zvvrk8ISTstvmY/ODTvuOf6k/04C+4CuL7kcdm/
+mu1c8FfF6ouJQjp+xXIXzT7OWJcW6BmmvjFjLqs7y9bMfuPwAOxmDpFI43BVDvTJAjW1CL2QDTe
tJ5cyx68B15w+/exuTqLwbXUa8+oKuV9mNv/EZ33Vh6jiXpKV9cFXnQ6u3gNXu90oagjSLj2GLVf
OjdjVr/IF6MluTGa66LN1epE75HqVoNQU+EhpyeFUL05Ez3FUHN639pnjqrrOKhdxfWe6jVmegxx
Ze/GnfyW0xkWTR/pQho5Nmb+yCRqhUpEtrKZJgsamrj9LaHbdtqtNJEmXaZlwA1dzZAw3QoNCyYP
MS78KjSXA+hgKBFGZC/sIi2S7ydO3J7zAcTb18Bn2pzIYu6iQaSZpH27M48YKy68Fy1WuA7X+2MZ
YYEr7DSZVUY23V+fa9ZFDv7BJTqdT1Tc5KYPWNWXbR0x8T68nbAMANPyC3u4tWiK7lzRvmn0Fobq
rGtefG2kEnl3rTHDzUtXWfdI6CLWuXqMos3IRxCLAHAGnsiR+OASjgfVzYZ/z2YUsjuMt1iV+uSq
UtRklUWpP0JMqwoaVtIZ+Fv1PyfsR8odaAxI6n3JRGkw+ANX5+Rnqt3v8nIfP1Pf06IFZtEXVYgz
6op9yuQwkRHN9Iq328Kyhl61Qu8zrGrUblLm2I0QVzdeXefHGccrG4ZVmIlHb14s1oo218g3xXK8
yRdHVDsnkBl+AWfR9YEbTUMvILsjUHFrzY1R7w09G6kG+5b684dFQi/LldhWmPsN8eP/0/h654PN
fUKaLYsoqlKbnjcpvUS8vHPlgZVC5K4e3CPOtHiJLmJ9zHKtuIk1TbsHFMYgKMWPkjv81Wu1efg1
dfJ3saRGQEPVovdfgMkgOoOHCFZ0jMg+FLchQ+LVAyvZ7MIQ4A5vmaLHM4ho9Lwknp7GL4id3/u8
Ls7aVGDOkKSZG1IITexkxGuLLsjycEEenptiWWGKgWqQxvZseqAufm4Op1pVc2jHsKrzgxGkbF49
34PY93iayIxRvasjXZ5Tw/QIhlPgfVJ3m1r9vJDktlMps6v/Od4xYXDFXaB77N8P/qLKqqPQIxTy
sPsZeknk4bMscBNoLBHOGaHOa1T2QBYoqoEpZvZdgnAVWyFaxglaRv84zA98aY4EGiDD4DHzT2dA
hM80HxSzt2FTB+68v9GEZ59UDmu8pNMpwTjdqnlttXmKNFbWZwfZvB+FhmJ7oPtjWUTmYmd3+kLW
BuIZu96CwhsQz2qrd6KOCtT8/vrZ5J6wWO8IvqHSzxedOzzCj+LVrHax8p/1Y7gLz82gIzP2VNfh
K0iS2dqqQitd0YAbMbV1bhTeFhsWh3QiLqLV3iy50Thag0OW0aJpBPzs7VWQP+GxEuCuiKVkwcX2
uE9/7dG0WGdJMvWeiK8QzjbTcy85HZEltjsE1PJPaveki16wlzLrnhaLkI7mdN+gnBhuy92Qbx1v
19qta3RlKSvNUZvG/3Ssmg3pXsLnPEQtMS+sBciM84hGUhNoYbt6xO+gBxq0uSUsfv6wiRQxsRDc
PDJsc7A6daZuZ/l+QK4fxj//W9a8USrOWFrlqZ6du3YVMjagFe7UyzWulGIO6Cg4oXK2csSHPwJd
FxHLBldYbCjrYOOX/DPjh7zaqkFBQa4P1OA0hbTegT0T7leL0ahT6qOsIeXgQaMqrs3Uyam8SKjf
VKUzAKe1MJp27StmKFHRf5Vxm/Cd3YoTps65hn+o6cZJX8sGnznsm5GzNNJUL63iH1WkBuQuO0Nn
EpvUYVMAsZ9tE2fpVONUKMIfubxCxFCecMZu57usjngMFPnNEXp6rnmyWmTEEhi0E8ZAvzeFBUBh
NSBZSkstwDmqy7+9jO7ZCvMAPGwc04BGMqe82ym0wWjfh2ZOeS1WNJn469IwQUDE0ubbvedWZ5bO
Y7Aih8OVF2+LEEGBnke2lAgrmh1LJkgbZvR8DVxqxJd3Iih5x/jwmPtsYkW0opWISxA9GT+A556K
pS4q2nafHdDMfzi+1s5GIe8UeakgLB9xsKYs5wYiMO/t7aPypo0i2ezcGT6ZN/koc+Lwh5t4GjIh
KvEFN7Ih19DvtCXREW5Mha8em0skZPetYqdF3eyVfRqxHa+2n737OBwWdITlXp2Uea3oxc7JVw6Z
KW+XuRWy9WPC0pvSubzpYkuGZ8tnpmdh95gI/eJbcLf50ugHQxGb7QanIMLsfexcmtjEej3ED8TL
Z+yDRtUmb1rnhlBykxYQAdYDAzIt6PlGDXBUZhSvwiKHjPloiq8Z8Q7Qs66K9l364ugWd6X7Joks
3nZisY00F/b08xUOcXnD1v0ulxT+Hrs7PGAeFmFntJzV6MWa0J4f5u3Lmh98iobsKuMu8qIKUVDd
6mwxfK0FLpfwob7z1w8t2CQkEc+daLvTIBzYDZFto5jyOQWasaEBpgy/rtPZBJ6B5JnsodS8dsle
qPo8p/zE5yudOzh3koFITvFUTYDmIlQ9GXkIkUh1rQwChXfeL+UNnicHOMRATZ7npFDgC7dEBb9J
Pm8o+mfVyao6uSeUajr+pt537d7pObmBWJFstN2WeLfdlwsOKiXlxZgkMGEec2eD1TsuFUX/OjJp
Cib8vH4uyXXr4vSW10VLXqqYnMbMEaFSAyKX13eeZAsQHROd9pSfNC0MyXtPWiUsm0YsboqhwAID
di/L9cf+SJVfN06A6E7aEhQUz1Yse2yEFKFGIk3UHdZnPu/C0nd4hyyxIcJwHOxvf/TFWuhcl6CY
DyB6TvswBhL+9pok9ZxiDv2akUNxjYwV0AHzCC0IA3NeMyLX9X2vJLCm1QEg77dR4M+o+zIyryDk
s1ZUuBj9H6wRB4jP+gFNk7VRD9yGrFeMfBsyIShwg2qHQWLs6458krsBqtKjGamBIeZUTQqyU9JV
eiGN/lhkdpuzmsOmlvGuhRpfKPFKw6MrVj+ahU6CQeyMPsOITU2pcY96/L7OLdIaQ6CRsJH4S3Mp
W3PMCcpZPc9KW5F3QVqBMHJeWNVTuo17XV5UhfYzc5RxBcajBYpaFj1HtElG6WPAn6+60nGnKbwy
cWp2QRsinv/8y/5bjG7klmLMgib82teo8ILNl28tgP+DO8PzhujrAXugynvECRyReNoTx+LzQZdW
XE1TDwt6dYNMqpSIFqZbqoOrQAMEcb0xjevQhHeIQg0hyVQwpm/zQShAvE6HdQJiOCMqzQ0/lSCe
F7g3qaX2ujgaA4WU9zGHu+sN+uSeyHZGuBcc+qPgHmXiI2S1aIAHwH03mGhtKbFqGrx0y4KNX12C
8zZPVJjRN0Xaj2BsC6WncQuhF++1bN3GczB8PG4wkS2yapalIF4Fa3ep+2Sk+pogvnStcDvG+uVc
riRs80XZvzBgz0h0OeYHf++sy1sszf3d51vihdHxLP8HNPCrjMUCYmFsnSfMKYogB26WnWKAIo3m
occcC+V5JohUMjlrpedu/r3Xk60PpKrVfjbZH/gFTbq0ZobJaC8ZP47Sn+kEf8gaNzD4LQmR/Ii7
he4Ng5e3rtH4F2P6pRQqkW1C4xKtwEOVl+aluln5DSvfp5WUGLRne3ev24fdkDE8+bB4CP8ERvXi
rRV/QCb9Y7L8QbhTRXQYSOrJJxuU+exd5WgH19u6up1XWBOfLmuFIWlxLlqUQHcgfb/bknwHhC4y
3p/lDBvDfbPJ5KCyC31lIs/yySbfwbF9wcID57KtzkKpOMZyzss6K7MwPbTzithh4z3rBrRxsrJ6
dUhhXeXOAiGxaGpAUfjhFsKQY9OPPJC8gFK6PC+qGlFAwOCb/4KCN28UDBarCx8zTnGdbglFH862
CsAzQmVhOQlgS8uSIGzwMx+YH5RfLWpEvTPQcbXJF7PUG+xLbj6qdJK9P4KjyC0HVedcZP0CGax5
bRjL3TBIecB5vGaQdEhxZJe6vIOs/nDPezBH3xFX7kK3f4MhkSLjxPnFmCtLDfgXNS4vngh0SwfI
Acq9FI+tW2+xPNkrMSU6clrCy4xokrjdmP/eBNvKWtIVo/UCtpgQHe471Y7Pgozmt5CXOS9uX/a+
c2PCxgd26CXEsbvBYdg6rKC2EqqzLYgq9GyA1yq6HDyJ5PuODS/lRSIHkBgaT7cGWoffHqVSzy6R
VnXcprEeArQ+MwCvrw0AACtQle3X9Diq/YIH5hfyIWQ8NM+0vQ3DU+/whecSTQCrZkqD+Gx46Udo
OZoFXq0VDMkP5uURoY/z1QZmYM0OLXT5cqC3vfPq84yN9Ca8n3YDE8ubirq/Zbvhb8PqgH1RH+0z
LXyZM1bVh8SgfqRJyuZW3pNK7hTjcZUlISnqqAMzqxBDfMt2OLdwyhAjm9svBa7BEYgiZ+0v+1C8
YHGTsc+Hp3D23/s2RdCKdaOvIFND4DeQ792wwfZCQTyrBmsdO+VPT8ywJ/mgEa8R97Mer70/TI1u
WjHuzIn5XvD44RaeO4ky410GlLkb0DIswgugeV4ebASGgqVfL051l5IWLMlF7Wqz6QvjM9VrJPnH
bDN6R0GhvWcrmC+VPfwrQFz9ZTlucM/lT8MUTpaixIr7GRuhG8IYlbnMxRpwx+JmH/z4wxKHA4Nd
Z369Y/yBnvwk7VZ5DclAVGk+FxjhHLA9bK+8nqrNaOjwNNbnqPG4Fq+or+li91wX7zIWetJ65XVd
QgT65ngONILbS+ZKgEXLVb1Iq2hYlrLp4bh4K6AukpS6ZLC5wcM347KZIK1qdVm+VfjcmQSAvF9v
1R36WSySupC5l6GzfY5W2wS7y9N2+hA1muYk+grPFSF8jYM6ikEvQBKeW+8qDixGIDBZHs9/yPBG
KcA0MyAUtzW6tOr6t1ZMEUOKddezaLir4COTCjwRIYomlnQOkpmHIgY1ZRxJe6jGPA/uRNC8iMrV
oHHIkfWxagSorSC2FDnZh8gIuBRYLl85ra2BjbKBH5OjgEcCt6lh6UJ3O6Fu6c5mS7IKjksTpQMu
mbnvnTzC8UESHpozZ5a4NcL1/i5H19PrufbpP68RD1GH5o2RmNptyrcNqg6IQbkNCX8wYEN/jHo+
Yk3T2cgl6J8BxyYH88W9pX051d1PpsxQ1gdWGLmg5fqal4Btl84jZQ/vgBnPU6q4NcImlDNu9jZZ
T27UDu/Ahu7yjlIW1WQ9pnCny43eT/Y5opGQfZZHoVQrS1vJefvuI2H9HnW47yq5ANcieMYrIjCj
AfTNAsaWrvyZczOncrHFYK6G/u9eETbmsjj4Mz7KjPmxGJXsdEqT0K+UHpFAGOCmovsxiibfYijG
YTzFTv/yVB/rmQvRp6W/06iqqCQIxt6bRA4+K1kl0eYjjV3BxrGDct8UHuyBeNaGAWSfsAtMZJHn
QOFQvca/yM1yR+X9RK6m4rUPbsMWKiUUjKUMtzwLyPq1Qd9n4qPWUdiG1PNfDUrp//PHsUkOMEWC
R1Ej136Dy01xeTpFFPCzxiQchJYSD6Oadic3mVXv/lUaDZYulrtWyEnEcBsBhgQJgbOrGAd5Mdkc
BxXAihUGjgKG8dO5yEKY/cApr/Gr28RYSsi+FHpe/CYYf+VjM9p08H4K89+rrXYURCLGxHAecaLx
ndJ45GrORwuTMbwfey5ZnFwYZDNbn3PbabrciCNyEqcPgG0EvmkWwQ4sdVLjapGulWn5Q5w/mWIu
1nx0SlLuy2oosC0THbNB1NLgrHUWMo8ECkbMA1I/5/X03/LyzNPFxjawRDF9YBCUvcmoGWKeeF/D
CPQBnmzdlX7OGoUpmI2tFJUIzWseMbunt8LE0fd8XuMMDhO4pa6CLd99A3EnZNloqsaNOJ8GBd8l
2rZV1glE2PZkbrVE/Hceei0O/P0E5U2fqu+UNlMyNbUb9yv8ORcD9L61mp6yfaFWEoimOWimv81s
C2I0qupbmCGuwt0f3y4jv9V1/FTTk3eL2bD6JOOUW/3Gqyk6CskoKxzpn8lWVF9WTIOCg8LbvCjJ
nxEfXeXA/MIeFGin9hkei5Sij4Ldamh/wAfKLFNeh04uL9UFpU6I/Sb+02Hx0CVSTcgK1Hk3u+ct
1XXjvd9c2+QdGKNOo2F7igVca+C/HIrGnOKySbnqScTY4BqweBmWTZ8nY9Km291CXPMt0UyM+JC5
u1x+9qRRaLJatbnOpSrPmjzox069Nf6zVEKK2qdtsoaL4ISoCGQ7pI6lV7PymzsREagzXdEHV7VW
YXk4xgRHvY5rLPik42nKLVKpPAtyKkL5UjzXb5vP627EjZbz7PLcwHNBBIa9RpEeQinc4wKb++Pf
SnYR6tCKASs0yMsvjcmnA6rrTMaRvUtJYm87dhurqsWbO3RLHsiNlL/9RiXfQM8UedVGCSlvXqMV
gfXiZ3RdUzEKFgxQLT38aRsJ3/eEzZSRGg4u8P+JsxZ85ya/LcyZtGwKeiCXUle09HXqtku5j8CI
2DiL9cb1rrYMr+eKwvVtXKUQH2vc+zU4F0gzSbruQZ+plq5KnhIEn2gfy40OwY7GwhLReAZ7dqpd
FGF25t8E20TUm0Unl9ZQNPa951nYrhKaSNY+b03L3NY++XwHXXC8Ps3DAGBr3BpwVR0PpvtsmWRA
Uc7HAHkWCh893D1dwJRieCTRXYJgOx2Rx2btpiFR9XAHeZxXqgXRxFubd2YnfhcZarmLJxDhWy1L
DrpRakGM03B76GKa9MhCu6auZhXiCjRCM20tx95K07sKKBaLHacmcKhvmd5jzHr9RJTahnRQySho
lV47o+deRImK6UC+VMIDoa/Zgh+4NfltzDmAQ0k6FbuVrFUmEtEbAniuxnAOeMSk8NEvF2VaUinE
Q6X4jB25AP9JRA7VwtrNYmDzh/VuRsDW4ph78QEjBS2loQ4zxIZ/6Dv6nrjdOn/d+jagLzcHcPWa
uke0r82t5T+L7P1s1qMinFoIHqOGyPJqE4jZn0u68at0R3vs77A7LYJPxG7t080p9G5zVdheG7cj
cECtKYWpvmWHrhJuVvwLAhx1vkGtJKIh1nuh/ZXxeEPHlfqSai1KtHESxEcdetxBDuJGF00LvRDM
WBcZA2nMCqMZWE8N8ZkGkmBQQCvSKRWQNSPcs27ALwixCPT0pLWGUBC6TuXTjeb6JFE1ryn7pkNs
aRMH2TWb8wGajRLVAbdmWYEIqmguz476g1GBJYI2DWUXilbky2aOg+YOSrObRKL2HecVzN88xcQk
IbYSNTL9/LdNz1BGFAamdaZ7+TwsIwJ+ipkDNzeJebDvv0nAi0uBnn2QndSHwZB3vdQlM7EVuTTS
OwnrTP/1rXgz39FoBzElIDzQj7j8Qt9Obn8BOqfY9CNKMSerfIfHl5+ztEeVM05bY5eZNzboX6zP
a3ez3hFU9ebFaPzn4J56tm/sAhVCrBMOl1DIFjDaceQe9mXKgDuYzoZ9DaXG9h9pe5YM/+hrQco2
bsELjXvzugf919GJSatQ5sRGhi+nVN/RhfglqfvNltdeck/seLsDvL0Sfy7VYeDmx9zNPp3EmQAe
pWkHtmvyL4b9Mjj9yMlJbIqIS2Iip5966jMQc1dr37go0mt+//Pdqw7/y/oYzfi68pruOZ1fM1Ge
Vo/TWsLtzSV2DFc5UAiU09w7XFmm7FsEsFgRcAS2Mo26w5YAFYKK/SQI1Zo3FJlLHFGrIKD7NHq7
LQqyJEOcUnN+6MusM7vorwukrLEzj3z5Tc4UNOE/9JayTjLv5gEiWezRHxz5fAEqNuyGmiky+wWo
gI3517WD18pIGSrSYrs/SFR/XjK+yAiGwKTST3XSeH7TGWvfJPYrmouTgO30zLaix0ewXZ1VvZ7z
WkGss0iUZTkD9rCOpvnEoPvHFlZm21xCcePyEhkZPMOpRytlLiygpAbKgjgx/8ApbkpWFMhLv5CK
w3L9lHpwA6KuGujXs2Tgc99PnksfKfMfs1gEhql/nAwz2XMH2r6fA2nlrDRvMScH/tTuqnLdWXKJ
+OwBJxba3D/rkRHaI3uKlnA3lJdvYmzHO/W8/you71SCvef0rceyrYD6s6SjyRPnkS/LKcyCrMRO
JRM+9eUeNQrLnC4anHNNu4IByNkDaHZNABRgMC4MltEI+XJr2b95DL/YH+TsE16JCqBdxf7j0fST
Js21xa8R6HukEtBzYHs9Gt6EMECZbsGX3ceP2eEjPOshGt9eYe3Mca3kWw6INQsJ51HAoGEg0qZ2
G6caAPqDBaL+aQnwnfy23kr6nhM5ByLD4Ev2I8dC45A6lyx45kS/Ou6ROND4vWIcMjQaevKR7Iuf
aN+146PV5X2jL2d0xaBUl0cnbv9ogR1Rn0PF3SeV3TmGWqPVpG+uUz6Qiy10IuFGmyUMx4UlYj83
Wg/0emo/CK5lkFGVEX2N8SkT23K/KuE4beou6o+j7cvyPalEUozLbMLh4/2GIxNhj1vyQbMJmwIi
uARqOfnE5BLi0UNa+XxPSn5IPPpX7qSMqGwxiGRKZ6V3tGjzgnhsEy9r7uOR++GMI9nVJwBnq1zp
Jd+/eVI9x1LDZF0mn1lYcr5jCqQ5Qevz9OamNACDVDdGISf0FBdKI74S+cmgGfbKNGgTZztn2GT6
E6z76ayZ1kEZ3luXElMRyGjKc5ecC6UhpAqeLIK3B9dx+nwV8rOJniicQeXrlypq8cNASt8IX4MZ
8TmHvbIjcibF1StwEdpWIMd7o/gMCPVRxrn3l/F3yh+h8jQI2zOiO7qLFn0kxjzFK8hs/zpnHDNe
HVJawzTt497UvAoaTlUJwjxsgbtIpljwIOWQ3vEqAkxpLSkiDgYtmzFhKRI7WH0K5B9hgeFmwBp6
oYjTV+RHJClP60OZGwHgQzUnhSHF6nV+R4S9bv2xuWpHz7FpMesew7mGXvvBbVGegyJd/3TLn+7I
Iw8JmnSVP2dhELvpHZDaXPuXw4NP6y5xuX38bCpfVh4jGwKUD/4nek2yWFQ8NfT4yZ44115P6TK0
lhkRXycQ3Pd9AK6O2KuNUgp88QdFdDPm8O4ogH7dOb5QmXSBFXy8+EiezbmnFukNzjTmi9PLdXCA
afhPmgeuhtRREbs/u1luI3I8kzu+5JP8PqfIeugG/noZC6g6XI+Rpl1Ae0xhNJT9VYiFFhjclPsS
LruShkHD3KDU1svtIkfv3HPYnvdpmS6Pnz3L494QCX3SpAd13yKvczmcPy5Miir4wC+FWKIBdS9C
9vApNWjSfHNGblWHcdXmn7vAGjHa5yv6p79hYwdl+Kc4POb7v5Wh/vKc2+ZEmno/5rAKqSsMooGr
XAFVWHipVWzy9kYZ5RsrG7E2ZzSpUOjcXISoL++z2VSLflOeWQ4fvE00dBdd2XZZLPFi7JU8oz7w
Xu+XJUenH/EHlUqeYtHrVzzTB8srC6SEi8317neE/HB59PjoZ5ukjcYsrSuyL9YGzwS1if09ZG2N
KqvvCn/2W+Kyy7E2rW28AuirtFXjWOMC8VXCIOaUDE/9KkfkVkRDRip6WS+iJ+46dZYZxjXakwCC
bWXo0qMfx6GagLuHGfx7QdpfoXhyUpdIWKuB2ykOfdzA31FV+yrjnnjxKksHHSmRicG3p5Bl8lS/
s974Hc0nl4fS2dW4KhYdbvdo57Hed4ynMZBw6AMNVuK4XQ7ANOwPfbOmgHAIUgjnSGVobbtwueuZ
ONzvZy5fbyq0+7refNpYiCWoeYtiG8BfOrEBfYK/LGl0lIRl/XDfiLnaALufXUu4pR7HpAKxSfLI
MtMfqZPyJXv1+j1wTsF4VyAZ9+Q7Usr+4rr4y/uSX/QOJ4mEfgrllWPwzmv/6x5Z+6Ls8XsVLKeo
YFUojQrQ4dkJV4QLADbXm1A7jlli5lesc+4k3WjZ/xdYjHwSw5LwR4nZ+Pzzu8R/UULzFoKn7k9V
uvEhVQtjstz75DCn+57AXb1RUjZWyrtnVE53UbdzcrFDDToYmrpmwu6XnAGAORsHjQPoOR39WpEL
N7IsTC/0DskKD4y7KYgL07k8C0tIjta+imN3taA0hURy2SDVL5DIjZxTo20EDpsLFPRQ6Mz3l/or
kAmoMw/sEIuDJRgJAKMyQ/tRkTQxTzoH5IRNgU/s8KEx8twpaBFlAclIV+BvOqkXnwup46wDDxTc
drzbhlWNsUYMod9YlhZNFq7XemJ3WlIEjRn+5R2AJISpC1No6WJDh3q4nphmF03BqepSumy1ew5y
6EtrRzCAgZz6kf27++hbUh2MklIfLRqWkKeF77anqFzCVfXJssmz62EU+aAg7ppQGXCVDqfMtkZe
RAYJUcrVrkEK87IGzFJzTWRuFRxKlEt4j5gUO1NmyjeVRCUyLzVdFMdWnDdPFpHh/FCUVpMyla5Q
8VRsjwButdxy+AulnzLv4LAuG02Py8fo/nhTLUypUOiGVdcmV31CuvX+ABj2+2YR6G97vHAiIZvU
rquxaw9xjBKnPEQYl+JKdXjAaPpTx/5OzJAl7aFnwlsWjoePpmQtcTHv36kJLFXjLYN/kNeUrsGn
s/CQZ+cMQ6EIeM0Ykk2t4JpxvDCXxM0LYiCwZkrLUAsopTUjlc0LsJ0wuPBB8tL0OQGUPtOCULhg
tL/ZvuPGLajRXiTb9wZoKo3/OaXO+KyEiVyvcpo4umMOhsvPvawVs1JmwRXgVcFu2pZaQTRtqpCx
sDRQ9k+lgXENst4Kf72DHuHjVi5g9WW+YNRS6u1ygcNcmGcqMu28I/LYNNQ12ajq11NMwNdoMe4V
n7fBlzZjOJsWCk4efOqeP7O/UzOaMdTuAt+ECsK63z9sukAC19arhJWuNpjfSNfmveB+GWrgzqyO
8rYUU8844q5hKnrANIcvgS2YjM2i0u+Ip+6N+6CIBzNxK6TXIV3MN21dLXRqHdY8nKjdVPNm4AtP
uQz86bjSq+Y6chTZP5J5F3Uv6Tl1FfvZLKoI1R7bIqhck8jc5Wi+bBfE8kDczrcEbWWCZEGewgs0
0ANXIJQwRBRuSBnB9bpa1EwJhTscotjw40WwoGbWoCtOaEBlNCj4yEFedYM+RyQuFv4u13CdG/xi
s45hRor1i/k120HUNjfdRxtjNXCJZdEniQFnUZfinhsychcj0dTFkMR43psYg/eXWcmzChC36ISu
RxrEEsKGdTe58YvlZpr6zXqRxZiHZW8tnKIJcB7cu38ispFsiCG39by+D/tlRkWIcBWU9HXvVkXK
XkqbIaBhV/pnjBwESlRczj8vUGZfadtL613CAgYuoSdhZKc7LyG9Qf0caWY6zFwt1BS04OUDmlNR
l5I7lKjUrFkX6ynYPdGVCNYNMSkMBOm/ti0anEAOz3iTyZLLqVDb1asUs5Ri5r/OQuWq2kyk0DQu
sfGE39YkB9xOD+Wt+4H71sn9rhtx4QAFn6oBAXrtoGqHV/xLv2t8ciOIf+Qg+U45rlqz+9n/smyR
6PmQjO8AJvAWLgssKIvdgC4H3xdEAdJU72a071ZSsWgZDGIxAgOOYFVU9tRn0ond8fZ1eddWkSOR
oRS1Ja7PXzOO2nvxoMPdN35zk8uHcnfLlm/soVunbbdzxyheI9BJT9t+o08yNzbUVj5E1D4BKdI6
Q0TuGounoHqFM201tZjamjVLXlVytAjS6NcU7gtNxSRvxTf85kQOgmN0c7TQ+CVqGMIAxaHsPp6y
cQGEeqhvIOa/uGp8Ico5wseDc89OlUwYAI6kf9tZa2OwGicHF7MVnhyeHGqp85nR1J7MdJIwHRNw
lxVPFhLPjsYdn8PThuHeqVuS8YspyXD5D5ex9d6CPdxWlunAssWo4wCukINKEdrqlzHJQRUM7qFE
DBS/Ea4QzdNHna70yUz3fIl65hJU5yvOCL/FOso8qHIEij/j3tJUe4TRekuZGM3RVrt7vBkd9+L+
iOZyVa8bJXBoTretAQyd4YFfcLisp8M80IZv9D7jlUJu4oI4p1VB8aqvMQKYRMwgX/UCCe/LvpYR
1SjVdf6OWHnUjZx/98uiygH1GxCpfBF6+Ql9WNKeKKcXxxHPdEkqGOtgZftXW2Il8EzBLoSqmeBj
eTGSX5vgn1Uj8M+M8efvveTuU/bq3afguJpmboE3S1aSE9eplwxRbouZP6OtEmhQiHBgT5c0okIw
ZPRpKKiJPV5l637+F6Lsia8SAj7CrTEEwx8yPGOWKa/4SXtB6OwRWzzahUa6B/QNcXjBjtSazAmE
25YuPxvGGG/Br7K/1LYwsANKwGjmgczaM0Y+kUv2YkaFUy7UfnQDQ/6yfd9+JqnfOkg7sQSG2xsv
+S84qMKQkl5lM4Isd0WJxkFu4SHEMFR600J0dbDkTQOovIv0kNLvXbpVgj9v1X/IhwEYrcKATk1F
zeNmQyUjB+1y4AnTn4VR4uga9jMKCBpfahW3w3ADye0xTv6NgGn/gvzqjefQqlYiXwK7QF4jaggE
v8FJ6ih2aH3AXktRWx9Ct5KvoH3iNCrkVaZ6xV5IjsZEt/WVnu3GpF3Knmf6/qggFrnE6GdCQNF1
Xr9+fqj4Ou6C94OdOZV3wXpxnIUsxoJ/op5UdBbXbEtKNwK7WDA15M3MQ033pbvBTytJfAxHmUAo
hKq7tYBDZiMbaHttmc0U5sBzB0UXPtu53NkdSfhPv2Desasn14yY6nzt+4+n8FbOGXzF0N5+0N5H
o+5VLuCLDS4GhjkNAw/Wl1xyfimVxeYD6T5Nnxw1GVQQoXhCxjUs449p+G3qDEGSQ8ZIx6marVZX
53ttRAG8YhuTfQMQbsfeGyGj4jVJFHA+LcCC5NLmHi/WcbTzPvbVr3d1FQBT8xF5lK7faMcmyvYr
mRpADZnvJzEEBRaF5F2b1hLHNNed2V89cJNcGL+ALLcnzvyZLYf5n0RcCoUId36kZCoAjNj8ihFz
nJ8NW8AqLNnzS4OdqVqlVwgquJk58kZpbnOnLZxALYtgcqXFpDhcTsR8eCTIximXhyM6Pd0WeM0W
L6UVbQlnsrM+zIVVtalPXmNEszfiG2fdyKRIl/ucsN7XpjEOp/m0NCEBRmR/APwtyywQu8bbIt05
VMt7YsLa+kKyTRXZULNbHDFfmEi5WWde7aHWBVS3kWf9NBg9Junwa62/OenzOBWPGBXp9OevSmqW
j8ErdEqkurd4jUtdIdEyvO9L/pADmdAV57+BUPX9XPVXO4lWZtSqwiKdCFK6xwYbXqz2Az2/Fmzn
aQBh465zloQ35JAN5ER5pN/9XLfHOO2rUOuJKJy+RxEzPQJ8maih576x/7rPcLtN9UJNdjylbvC4
KXk5EYlvq1nhmAtIsTc9XOaQvseJ1N25HL3PXpQ7EDQ0QHGab+VV70UD841xMHpQhnaL9y18UeCo
nUWuQvh7ZNnbL35xJfE6CYWh74IxSyCZShnc7ERWvgcSmAgja/roD2Fslq4tepXo9lEhp5hIyLYz
xApvOal0TRXsiejQjjQYW2iBL7UBEGZhb8ZXKLNhkysmXIVTUi1Q7y1unEKLu9RqEPG+KeeCMPJn
Z7Bbci3X7hNS4U3mjWU6YdRP4tYiv+++nqs5MQ4Qh1GM92wkSQqyw3xiwJ3wuQejkOtPynkkhP/s
mLsLA6RGmYKGXmVWkLLgXu2e+ALHK9MnNYLNx9B2JFVJqqloDf8g4KVRAB5X23kkJ3ui9HN8+yJD
4HTupnVPXGQ/d9yhKt4RUE/OjENs9jJRpCvUac+QqHOhpsVEPqBeHQNQpEVeY3vrW8MF9wm+koGg
kCjcT4alm29dvExdVaNgYCOFZ1ghtCYdTb4WSKYvkOxdwpZnwaRs5pmJBALAIotIEGAi9ehUWN62
mEn2j98WRXHrKj20wy/XtVykzzJJaWPtOS9GflvZ37vyT0qf3n76SlxLxqEjzo8x6LgB1YC/q+TT
tLev4F2Dzw875curJ+khbF/2cR2K3NRKYHJUkE4rJDAu2tal/t0jmNZ0YC8MU3wv6SPnW0xPQ8AF
/y0FPhbUP/b7QtqGgkzHI8SwGJdpfOGvMp4SBnkVBZjoFZ9utUQcaQUpxhyXhfuJ+yp3mWJDdMB0
71e8lc5Hnoa5sOFQn2p9jxeWR7esHDKB34x/aMBk/GnHSrePMyMyJRDJ28JN/jxyVN6vSTwn6Tqu
/oB7bfhvlL+ss1oQMnsoMnFmPbkjBrjKXiYRHwtsTY/AyMVGAosUsUvHJZEL4ygexr3p43mZn1zG
41vQvDyY/FTa4qAb3g2EzfzFUp+bG5NbchCCqfw93lSmbRnp23RZ/G1Eb32DSVErnGW1pe2DvrCv
bkHmlOVGA6hupMUWxBu+MeMQOnPMXucLCx0MJnk661DzlP4wWn+b/ANH4SeKKLsO0tTu8UVhxgm4
BKLMKvFCcHMwOZaCgJuzoGINWgsjkFI+rSz5sUwvC5un/9x960uAfjArDK9u20jSwOdIiT715ApM
oC8hB0mRRTh1ZaPOjubbMw7FlFAO/N1EoHcNfgTDlMq3XVYfu3RvEbc2gjqvpPiKoUMwx2PWnYQp
xD+Ne1xzIXazPdk/iLc7ZIHYbbHlm7wUirKlhM4QU4TuBqXkYvoM/2OnFuaDAPCFeSLAZCtPjlnd
WyFYcKZc5vhlj/5SQ6hWGKcCOxiL/vE9soIUKs35c4pCFE0xWo4MLt919Dzun1nRpkb0tCThZlnn
crHpbErDW5JwSZKUchU5+JoUcqA7laBSRQWLk+xGS6qIY6bTRk8zoawAE+SWZOoS7AlLOUO55Nc/
Q0XS3UYiFMfEgS9QA9Cg7gXZTIaRRjTkdN7s6tzC3jnZQclozxh6EyoNtCXJMmN0Qg64mY5GaoW2
3qhXsVogIpfi1EjdOOCW1hwAk1uCJvspcZSsIEV/AFOQmvXAxyC4ARwuX1DeVAaXxakAOWzmLL2J
ul0w1eUI2+lOkNwKPSAvL2H3VHKuFRQzJFb2Wq88qR+wIZmThnd+FYyi4rOYK6R3CYlzVEpVQL1q
E4OV+1khppLcJdsuLcQPDLkk7dneo2e9nJ8Oe/OghzcvQ1M8dKMO8HTdK6T8ZfhGsrgJKZpkhzV6
mmdG/n8UUbGfh7nENYL9lacfwMl4DwfpwUj6Oj73WRVp9+Y+v+NuYLg8ln/5GO1Fk6piePko+eAr
hViCBIq7sbLBn1o7GaJ2lMcog5Jt+D2NxDeybTIxzw5E8/LIUIkUpXEz7sdkX8ePlz/iMQqtUcwE
4ehUdpgeDyPnz4b9x/2yTtr5JXmRBYXpTJJsqGxxe+m9T0FYnH5/8rwuHtWRPZ6Ht7P0O0nAAQbw
t3ZLoa4yJ+cAL7NjcN6ljyEUCleMmI7Msx11JtRtEUUOFt0Rd5zSSLL88H9DkyJWfT+GE6RrrA+p
eHI6GMyJ8dk/YtUFge7jZhQh9s1E6Hnlq1yVzfo0+zYHK2kUef4fsrgm67lAyMnPZXGp4qjRS3au
7p5KSTXzrmKCkvlICk26xpF05tUankMNv+mEhwBjYkpBlAs0OfifQNP4hAFmhaKfZwfRDbs0XfSf
Uxmjay9OpgqeFLwuPqt0nP9fsFby+ZWuCs555uwmU5pfBJRXFY8CuIy7gL0+9ePRo+cpNrynKCPe
xtYJB3W2eH2yf7jSgRnCy4+2mCr9Lo3A3IPRNnOykbwPkI9EONb+ld3YvdzyxAR+CUEzXFZcPnVB
lwRCKIoDd47UoBV9/JOo4wW8zppGEYrlXjG2hJQe/hUY2D41p3FXy9tlqdo/spAnb2Bp24ov/sbF
h+dTfwe33JPK5T89LMPZWm+Rx4NdAzkm5w1QVmReZFHqHSAmxCG5akBFPLaCfPu+XQ2VeTJjOYv1
FkBh7vgbZDpzeURSUVqJq0XYlDQ/m0mQBPgQwTmyVC95PjucsxGRZiOEKSHyqsgDLv427Xu8KsQ1
/ie4Q6R60TI9QECMeWoWH2fxHN436Dco5eoA+4jcEjqs0ZNQ36pLDP/0ZfLhj/QiWF5bpFxVbzhb
VI2sJPqScDTMxvRCIDseb2ntMtsi41T/fjMJs0R/g9R2ww3dU0A3zzAOgvaV7cxxC+Pkd5unQGQu
boEgJQJH53wm+LkFFaRZYWXcR5VMk5FowrfoGNUiw7+5RwKodMFoXrNug0mW3gk9UcXL7HweJYLf
YtTJauHVejJddiFD8sGMKYZ5kmTpG3NzO8e3QQTUw5T4wrkswUnsms5j7wgyBVeZdybza0oBrs0A
lqxEby9pRWpf7brjOWB/0wHxIqkZZhwjc+Fvc+mUO/DgOSZhwVTFwu2b11tRjwbsxDSPAMn2kZiL
xQYJMwg8Qm7h6AJJ0cGvHpqA/CfQ/lh55ydwpVGhU3rRQZeWIM2NFUtuNXTjkHqx/6JhFACn8IOW
SJZo1TJPUPYFXB1lXXg74BaeB/v+G2srTOj+7KOFRi1SbTBcMJ/ruVqL9MpHN2i4iyxAJ3zrlI9V
/sEpY0oBbtgq5XG0a25CUg+bZVT1AC8WXzMNvd1SMBWhPozC3R72pYlUYPbirkVQMRztFII62MOw
Rxbw2Zdw9Fkzu7xU7b/0+vnBI49a5rfRM2zHYrCssifDU/UYwe6B4d2PP6zbThdevoj18DsE2U5Q
D6kMKR8Z/OOWupH4th0jGRWb3Tlh+YzukpymRWX2vWBNnzJWHXk4mAmfCS6u9O3v9Ev/AAOFXr5J
4wPO4jsI9/ihxNo/uPJvLTLHISq650mVp1fq/10ciR9GqYmSXhGdhCBoebxyRt/++P73n5hrMQLQ
RnlD2S43VFBk6o8jJREAx7InKyTx5MvTXfSTeTPS64laIj9Fc2B50tFJ0rcOuV2kBdM8HDhY4Sic
zvJgLDqi1FzsqXZM0xNoecnyO1ZozGMwgnZ4fS6XU1gybWmEDz+EVBg0FE5Ai4HwZaTmtVC1tS3+
igrGVrIgVi+rQuei2FLagSy5a/vGkb8qQ/64JLbvB3HH83FNfapdiC4rgdJaZ4jB1bU8FgXRpGIG
H/i+F+db3M3pyi0XVlfuqCoL4EXNYiT88KR65ryObgWZsoAGL4nvUHeMO04iFPdn9CXIn4NyArcJ
7GKt3beDVC4dwmB9fk48kuaqzxQpujco9uV+rnsls85mjAsCGtILwpnP36leAcZJPN0Ezdx5VGis
X3OQc/Ag4OaQ95fz/8Bgx8f73X708eBfs9WwSXvlquDM5hLWHpSWtVAmHk0SgbV80sq1CFw3y6RG
4MAQuL1Z0axZSSD5An/dRB/XlWyCMgJNteVKA8AsCLm+2mTynfWrvkz5QbRGFXvJFwizMXxwZDTd
n7yM+x81/+I14PmWvpEk0Rq4JfLzxc4cn//ye/wE5+M3ynJ0GDX06+uUoFCTCr/RQO8J0DMELF5X
q5wG44yREmkM/3Bvj87R/XVVnxLctguOR777TWQfCpNC7BB6NCzGkJWzb5JVj959IJMPD7t1l8TS
tLGlmK2pjJOHbnGTCzCIr8aTQQpCububvjMgHxD5dt7ulj+2N9iZaU4cOeuQaG1AemUsR6cY3/Q0
RcgYJqZTfCFQEFoUuuHtvYPH/QOHIB6FAu/2dEbZ+S864NYwwzVA/1l4WY8gEB5ibwWXuIKFL1du
e6XPYgaynyNVfMLD9OKxrqI/6TtkiAEwKWoqWWxNZtzT13kC321mhmbqc1ilMp+YZJJahlKhQk0b
ksmYUVfb3BtD0WCm/Anpf4SzPHtUPkdtCACCbeZ8rrycVInHminyhMurBrgxwnDHldtpuXzYYtZU
/zU9b+0T/vdpG+nZ0e93SrdGMVzdJPomW133T42qNkLpE3QqF9F86+FOvxMbogwoQBdEM0H5IgdG
YO38g1awef74Gi78Ps/br/oSVqP9WVYFGkq96HxFx+ipJ7dl3HwNTvbefCm6kRflhAGF3SgiDfk0
f6/Ry4fKxuXZq504ic3KnKTNyVayL5BuRhqGHnZl/GQZmCuvIgs9vCqcbVRRIHAEx99d/BHI+XNl
DtvqzDw71WbIvgKdBsHfmC/6YszayBzZAVrveI4NQlU02hlAjb5OWzv/UfNVExHJl6Lr2rBJ+Gwg
t0HQVMfoOwoiH95yEIHG4o5LlpvYzVMaPYEo1nN22S/Ljt/AzlBTGumnTet31DJdZEFRbRrkBRPZ
ZIv8jKwFgWnZIM2DkL77Yk/itrGUFc284ZI3kWCEA9yi6KR6IuttwmV1n2/tpRPX1nouvXHieg5a
a67bljPjz98ZCHuXdANBu4Gp2s8oHo3QZpgAbNRRdIZ9CfQ8UdD0Pg6UhFjcs6bpOS2UL2/i5veu
/NSD3uP/+V1+ZFnegkRKyF2+CHbq7/wwI8FEQu9mpqGsuNM/IUEpd+VoAF2+kRQ73r9aaCS5ZId2
nhk7uaFxKQYq2XI0BMi2MxL0unlp8xK1DyqkpgupWnacPrrfWTH0CWPhZyZE7d//NK1oqwWi6Y5a
etzUJJftmmlEupWPrUoUWmUYeh7WsG4UEje5QzInWa2ZfTgYDWdYepQlZpldT29BT7Tc/tqAURgx
SoyqYgb838z8Ksvw39Q/xGPh+Y6iETZRr1Zb5tsJzNI9y89/HM5zvxQCcqRilvqEcn630px2tEwb
iV2ZtruBcPyMrQLQJO9S/DRr5/sLXRzDfywAEK6AzOQfcq8XzS/VqQbC0rOc/OIyS49bmd48o4IF
eLhslsfDHzNErzAYiD0DSsLwd78bn+0aT9FCcsIje0Z62bFUENxqWirtpu/m5NNASS/VFXbWIOtY
HwVsbO4/pcf88/w2f0M855qZ78YmkDO0SKEja18jNXggGH2kj6/XN0OghMw7aap27N8HHR6JOf9b
I9vBHlfqDHx40Msds9mSlM7XcLIbv64KBQGWqsrilaUR785ldTNYt9gKff9o9FU0dAJ3/ZmncUpz
R0RNHwFClOFgXbs8To/+FktvwsgcFxN0bSi3FKgwmd8vlgJymKcT9DrgFFeYozVO1l7wvti/d/9t
bf3/rbj1ch/YPkQaXelB+HIMz9wyzKHOQmiRzeX66sPs3N6tbMM6zKSrTlYqrABfBtMAaI5pwEW6
/ofJJ7fl4NCyhm0Yrgm4MliGVrTqPyDFM8kaRfKXQqyTQh41Jfd6WX5HRWZ+xnRKXNCuoZxSg9RC
DGil/e5azoOGGzfDm+31nxN3/V944kx0Spm9Ke2I6jGPzVWxGeptgJCPAPyGkVM9OMbeOMDjc3Qf
5XrF7fUHetsCWGNHoLd0KAOb8CDL8/O8iUqBo7K7a6P09Ig5IMGDRaiClWklcsBrdVc4x/Yf6+zc
gWmuhUqhkKEitNeRFL1uvqqLOIcPbAJbMz0Qw5Vcu4m+r7+TGxWK5CuNCPwQu7a9KCnz6pQmcipz
EYicddVaFt4Od9fImKb5/ms/+0Ix+KY4hqUarKsDSLocyG7CRiLUM+d3ZlIv0UgwneFjegaTm0Wp
MNQw1UTPEaWLwuME2/bmPAMC4yXRwX+4kbfNtvT8adAcLZxzLupg+JPYd3cqxYnbiLF8WV6D3sfn
Ogm3ycqF9sMr3NBsTpgPsI6lPPtybJzUXJ1Z3MBWePtZNcFG8nuLXJn3CWdhN5e2N8hXpnvfqIHh
7qB5pRw1JEilLKU3C3VkaJrKnlT6VPVbUeCCwrhk75mZ7ziU0oFiuOta64Jvs3ryWyhI93VwdLm8
E/Dc5nWPbM1tIAF8xKhbOwPmW64Kd477bwg233o59u/WJiUAArd819mGjfcglRYCuOnbo3eMDSbo
okoFvM8ZczKZTOnGshbdwhOvOrc1St7zx9j03SGM/ipEFgPPkfOmJa1SyoE+94/nUDKvSBzhF8bK
pyO9WU4AIzznSnf0mHoT1hl8i/xIcZd9RJnl0i1OGdUuaI4oV3LCAaQFGKA/EA/J28jcrJ9+ne6z
aMBv8HEv67nCm8g7/wTRaRsFaHtWX+xTvG7Enatw6SKK+t6MjKxIGqWuZxpdtyuGnWEP6I/jKpNp
EqFIWg1ksMVbE0pVEYqrXV0QO3CHRAKlCkV4GjqyNGLWl7iVKglwUrEp7/N/nBSuhaolxwb/JRvL
DYQRPVOyo6QdK2j3+KEAG1kZqn3YVFYTDQkUNCrh2V43rmXIHIF8IzrXRb8FdTF23h7TaT3wf9MP
4fvNr4EXm+FpiLEpIJsne4dwmsnhhzZ9pZqIYeb1093YDMVzK6+dM/b16DSq5NvuGqSrYDmQjl6O
tl+0xdIuyOEpx0DnbJhkLGXD2kFzv1fIvgufCad8lrLLvFgPyds28L+9HIcBLf9ehX+eZtQX8CS1
27iXTUtpn8dJ/m5XsjdyB7eMTZy9YIfI/koXvnPw6p7w2ra5l6WjxBUO7Y67ZVnZVqyS0IYt8D8w
OVf8dm04knXskPpD/Rvf/6RaJmXHVHcuI4czEF676RDfeCC/Y52hmShdyy3vY0ZaIZASX/D2ktEj
JY1PCFm9HDJgosG9guJBq7ljL2CUTRQ9VNx7JNyLnfk1Q3r9Afmp3X2PfAX0otqjh4zcwZ8DFGq8
Kkfaq6NKBTv+8h420XvtPV2oD3h3H/LgfGgZwI5eDmPZ1QnWO5C1OAvJHxR39ifdCrQdGfDkEcQm
sadAMnD7oxGCzjnqdO+tRS8yeIbWrm1kcv4kQrmLEH1sppQ2UtcCTIrMJ6UGVLijLSGUgDQCUsPj
ecdFfB/RjuYOiraQJUghGOZKXx2uwCnq8/Jf5LEIDNupQHVTzMLz2s6KH3tV10GrDVcFaAziYiOI
R/bJocL5haPgdD0kalU/9/GhqEevqky9qLXPK9nmYesoaaf5GmayXZGJRULdZfbxFD2onKF8GfKz
DBQVDfDS02m/3CW4C+vW2ErBbQ/+k8rktv4M1BuwGkWJKMQiRkD//xzphL3gM/6HOLCs+7EhUqEK
j2brv8JYuiXBULYR74RySRCoJUY0ova7MS+fQuwmATxiGiswvJqC02kOHzPQSClRU70BVN8CsSEq
bZJOQdRzd7Dmc7UyA9kgroLX7BSvdueuhd9CKDLxeC9gEU5i1f7xnG0vqGSRgNuQVOxOYnbhxT/m
xXEZyF+nZcqOQoUgbl4kqjLNcKiISjvlsgEnNyWXTiuTyQ8giA81V6C8IdtJhTYmH7FDLes70Mpv
V0spdtHMCdRTC8ksbAApAoxO9Ojm47nySKzWuh1A5HOMB9i76PlHS3Gbsup88EBF6Tx5Iw84ID3g
yRbMg275R7cjVS83bcDpMpdLwLjAGG6qxAilw02vIqF4ZC5473WwzG4KUs1GyyWUzfSLWXwZ+Ogu
6E2jXNzwZ4Oc9jeBeB2SKINGWaIV6cH9kvbbnKC38aypvS5EAeCn/k5MJdcaURL1tqYteBs49uvj
0R600q4+CeQooYycHx5US9fzrne4QjbyfR1WY2NwJWAkFBogLJLk3DmBv3j1Llh3vtefzOZKQo5f
oz8kUVtMnALdmXOEG6qiGufyjEmE+U3pggEkWl5t5LN1WzuniPhQJoqNhwtCY5uGlLR3Apq3L1rP
SfTmTXrmv9JqLtqiYhmja0KM5WFfYsjnxF6cLN7DkPXnYUFDi9FFG8mnnzz2uClFFXbIEJfU5ZzT
db+3fZXRmpFlgZoDDQbrcJ26lMW2e/Qr7FJ9yRx14mUjqISa4UjGTwHjNxck+RcNGvO+PdV5hft1
Lr2WVIN6/LD2dqFljhHMJQaEsQYIal4QTcKlmRMLpb3/nlZlEKorioAN+pGQ5H8aZgFakya4vUAm
/7vUMEcz/KVnvj2rGD7ndHbgyG3zUGDMszcCnJcrhFFjGMkd8QvW+q1VBzFQ7BdzZbEfUEwWid0d
isHqLoOKp1tDyTZJGnrRrpF1Wa6JH3bFIlDXnZ8l/3qa3nTRc03uAHPc0BBL46jxoLBRdanX8dbu
pycH6ncEYUzUnlcC1vkGOzqp1fGHVDFVIIuje0MGczhk+paohrCD8KdUaO5L+GvinUEeQNLkYkRA
zDb71vAXdsYNSrOXwioqcYrAMHuhW3CBLpkv6rc4GCKsrnZi7i5K8Yd/TL+SH2ohFdaSDqiCh0v0
7tWJAitZbBKgSxrHXYFJ1gbn3m+Sztdo93I+sDQ+h4CSF2XIdIybdQwOKHdZkj1bcdaHQQTxjenr
WN6J5kTdYQca7XsLQ0J82qankifRgaihJWqnkPWvUH5tEqM0vpAMF0c35Cgepe1nac4+scIHmRAF
HcHx/SMzLGtnuCDQwX6zktD+0qsCybW8ZCG5Y/w3RHod7FMZVy2Ke1GmNZePSNocu3wwaI4Z8UfK
dGNcPTubUhCM8R+SnRYD4j/01kFYPr7x2zjefK8aizyYw+UBTx+fB5kQ3Uigg0lAQE997CStof8o
Wlv8Mp7jhsxwBtRPqAQUWMV5PxxzojA3eLAVa0kW5mjKt+8vR26p5u8cPIoB34g59LSBsfuRryN6
38IrQ2OBK5bgDjNxwHSgLCWe4CR5gpVdQj5cy1s8UONW3MmnydW7yDSRuqJAWe//9QHgTPIZzLq2
/UBYTAreJ/kpBSRETjqwDotizonsUCIXC+2I+b1gkwALvKOihHSZvmw5lTu0igevvzfQ0SuW7XdV
rXNov/oiTLrVRL9pnVHozVGt5wMBY5fq2M4+Xbp3w9z6zRFgzURvW0iFcGv+2UwBBakpnd5SqrQW
Tl9F+5F/D2Vwk2niwLuKDrE2EAHkigKTPX4FA59rA8Qm910ytsAuCSsNtqOnmLRmbH/nIEQsbBP8
1J2d87olSKDryIYGE38z0KM0hg0oXr5AOIjrzR4t7gqf1U5Ku/v8fE8WD7O2h+bUHDjAkSQHssZO
jUBhWT3zThbqZO3H9rUl9eF/YTWFRA4BPR9xBZLotu/buBljZrNxmUFo8fDR496n02i/dzNXGjow
VAhiij8xD6Qs8HZYOWx1/ncb/iMKX5wyLKXyXedUYkYKQheixIY2rIJwoDq3LLLjh2yZxeVrzlTX
qk+WmWoYJh2vO8yL13zmpjkOW5LFJguSupv5mhT+bDJN3lTExTv0XPq+VR7+/KCE48gckJImTDYZ
z1AyqXufrN9kSF6eqoAJiawqzQeu10QRTs5syKvgVaEDQ9wEiKKQfrOxJVGkE9xhib3JhSXNwJbp
waNJD0gAhKYe1KSxoQZ732g98M/0gdjFYmGIm5Vl5sb3mq1HIjxTK1VFCX9R/ZqEJP299WkBRNrN
h8LU3WU6Q3x1rJ2yg4GHYLA8Pwo8tUKM9MwEiKY1KEE2D8sl3ydkYgZCye0cq6cIWHZNaYZjYbsq
hf6BGOjP1I06aOhWnFEVEJcCqIcJrQ8Ag5UtWdb4QVi2zq/4nb7fd/4mR7sKfnMzBdnGh4YcuIYY
587AtMJLtYzFp53Gt6l6vVhgv/DSLxlaCOPgVIzUNLAdXoiq4Kz22ZFdZ4TdM0UFH4nXNJecE1Vk
fFQkLXtGwTyMR4wCg/Fjh556jjcoqV9or+PsyDQDdcOspPSLa2xhX65RbcpJR4qh6OFRPbYTFvY9
EvCnhZi+xdHjZX4eDWIW1vM0yVsTv5GUmHprCwM7efY7p5KTK9ZWMdlk4HMud/ADfyRtuUgmblvK
7wJbeUoMjXBuNCX0xyb5UtEA408ELDr6rdvw1E7WTO3z+7aDRwj3uT78v217pHtG4SHFqOyLjew5
rJ0gQ+glGfHkrkrQCXaqxitXSTuez54ZvR9KXv+l4oit1PxDXHLHFfoqfkJWGYYpLtcel5jLwfFM
gg0D1UdeFDvdmL/D6PSQuPzg+q5l80YhYSt2Cf/SvHfyRcQjJ9M5pf5UEL9SXyacd74l+2V1hKSm
hIlVFxyfFGr7p9U+1UGc0Jb1FGN9BIt+Ao2kXnV2+/GsNt8QvJm4uHwbr8Fa2o/FxEM9WR/na3IN
nwY6ku+DxHsVpPpPzkTIkqT1Ef+mQ1pRJlDoK49Y9f1y9p15drjo69D0UMlSu45yP0Sz7Fy/2hv6
d0PSRBKivGvfzo5nimDH0ObV48dxVmU1rWOSMVED4M7i/6QN9LfswzWfnlRnlELbvKW475kLNo/Z
bwNzV66EgSqjHR2xq9n6Ej1r5COm+gkAb45ez0Poe1mScOfPoDRd5i0B9mywe+Ik+nbGhax839Gi
G6+ZH0EeCF2xKXQ2gIBAYAzzhTzDLLpqxMneshx+AgM/jhTrDCTCid0DU92z7uCgEfa5uN69TyMR
7WPDG+l9EHD2Zac0VXun7sU2nFT0k4CRNMLxzj6uUB0Hwtb0ywKP8h8x6bOUxUH6tsPm+s7P51Zy
iWkPQJzucm0WJrHE1TZxO9oca434d7bR9I7v3n2Nb+5R482152VgaSpv986pMWL1EaZmoxy62etJ
oQMi3OEN3hP+6lj7GAlbbvyjVwr5zGDKkk+UqGT1cSxVff1jdh1+qLElEDW5P9UPYtXuMeHY4Jmz
Ro1MGF/785c0sW88YM7i/cj+IE4abU+80VCj4tCvPJtPo+cJ3+lcrRfbWnq/9+7g8oDkCvcvi5un
d+/0AvQTGHSSYAUZQlyZgj9cAZMWQjw8bJ2MERu/MmtmnqL8oMMH/8boO0mbvlL9/rfVegRMp7sP
oRBj0AzKUkYceBxmwrGUdfR2L5bcT2GW5O9oZ47UEilQAHcC+POF7pcYMlW3uUfcR1f/WvWlmrvH
41V5hG2bYzS64HSfVL82R6L9wQzQP/DRgqGjwp4bUxEOhHHOTsqQQv54ue5k7aXo+8+J4AB3GPI0
hnBx9jtXwrWkMwTmjkQDgF5E+zGxm/0AibmGdFa4CaOApv6ICM8TJdRSz/lOvImSv60S+GKaxYP/
osleCYCxe7xLg6fTFoymT6z6GipglKSI63rvTFiRhTS6YqP52xHnvEGAos3ohyT6ERtm2aUwr99l
EigRG6xsMrsE1GkpCmWerZ1pl3PwzzryAdloTjhfh/h04JW+pEG4gxodDztmoZmxu1Cg/8MFTmFr
yd5hMKftl3wZi3RagFJJrQZP+2LPJsOyqqH3vcy7TC2aSuXgJaUqrYgjEoyhUCN1B8LAMcw+2o/D
aop5lhjkSR4sWPekuBcAxhDXejqVlkxZiu4QZqylSaE3zozZURIKEq1Md2wgZRyfyxQYZUTCjlAs
1c1ZIxRR0UlRpZDApiaszcDzk6E7WzhLlQn32teCtL8/jZxcdGjEH9xyViNoCmxLxU7LBF+0XPyk
QfulagmST9heanlwTzE5XkyCGoCPcaXJKLPclUIhFA9haTsTFEYQNzqLv0Wv77gnByfzpfWbs2oy
iCV0J5VCjRNz5vOTWa684qTekg/GAls+KpO1hYfdTVqbN2LQeEJ+SW8uvu320E3652Vm6ZQPtE2t
6qWaMUqNImWPNxewtAn7tE8o1F2Oz+fRLD1+nQ/ejjoXrBPpW8GlHnjefS1KNCaoKVVOZepshP0v
bxSXjFHOuK31tiPOVivbyPb1/TaGBex9D9GC00napncZ3xd5h5MDFjmrLIQ+0aCK4EANQBxVKJr6
hSL0/Byc++5BuUaulW7fGYfwJT9YlEbmHbcJKO7oEs44uBBPxtgbskgmM0Tg+Rw/XOvG3t+NXsdK
ngfN/ncM55NtiSY9tJKN5ZKhkZoSsuem/C0BrXXt4Cz9h9ydDugBsvP/yIVBpvyefUe1Hwqb5kjq
CBbaPvXC+6CpcpCBSiqvMYp+YlDro1KpZj4GRRUMklGutXF13I1LFpKXJ/GH7ef4XsgO/npuIr8B
feiI4hqzszKctQIkyk2WQnsgS2GaiaN10/E5XFxxarTp1SYghjArotIcBgQJSWtzb6OVMs6oSos0
8sDYDbQgfIbLMSgkv8ll2u1DRGC0sAZSApBj8CVhczP9obyVYKNNzF4r83IMv934o0LS0mtywL3q
BOzMDt5pXG6MAJ2b6hY/X0rdP+jeN2VbQ7ZiNy+2RPxt7H9kcOjtm3LnARI4mojAU0TbZt9ec+xN
LE3hfPT4t7nwjaLAmG7d34BD9c6YYeehvAlJkRf70a/c01SrZZqp4Dhf258+wZVdFVIHX2bpk/4D
mlZ/VTUNykDsLLk5cEBGjqPsYYWXPkbj05YxRMRORLrkj9ALaiObKiot3MDanU+c40VRQ4AY9+Ky
Akh54NX0IEwRBDqtZTExAiAHR5dkMuYy513s9WgJIxpGwV079UK0JxNbP575r/jB8LwaEhEVHwbL
VGElK069uNK+QB7n2l8P2oxOuKwJhySS83xxYzBXby/T/L+/GM2gA+wnyZB+YvfgTDOI4NPDpBHL
b7eFlL1aFHX+VXCYxhZp1jrD4J2UvG17MO4/Ln8MupjGfgYIKkZ8qY+qXVMOlYLDNjNpG6tgAwbU
A9/8PjRrU940op65iCvXsyXbvIfcSM5QQ+diMPaMTaCMC+70trCQYq2s281jj39bAfjjykTi3xqe
HyLsIJS3chHsEdN5i0usDywjg9pAkCsvMgPBb1BGshjv6aIWtjOdrnjGaIA92SBHfO25tZ6HnlaU
ojKBVZVg6tZmrqbckYtdJB0uKWSLlxMelRccut3VWI13CsHQoGpYHZZcZyjKR2mDIq4lR4ZxJByx
9HDVduoRCSWzI119rf950XaefBRQmyrXz8Ji0VBqy+1N51hEqMF6SXgrc2BcTnYoFCqZSbpBKZYk
hBt5Z1b4hOyzNY3IyIaNBCdwvxH7PVkSuDGsP++rmHAqLzPbwwlnXQ4qDfZCjlQGQsN6tOtut/Vs
7OvWHN3VFylIawLeb09mEYXzS6JF9pbdSCygR7GwiaUEoGWVu1z3iREzkOpnlQOw3V+nAeZ/Pq+p
YvJrfJbMW95NrejjiSszRRXJbZooWlt0MwsnO/q2cXin4uMnOZRLLDJ6X5KM/myeQgsAwQlcNUU2
C4orkT+uCuLQRUhYhGzbdA9VPOlEBTYtzTM4YPYTEl8qd/eYa0Eq6HpFRMAa/W+p6f6dyZJ4oZQx
FPTMbQI3joAvQluRH1bccrnFVXLb55gu/rwehsWjcoI1CaNx7ueuMFeSB7HzjOvZ/CSyQzUd7AOv
7c5wHQNF4dfiL2JpvwpMu9C0kCyk2Iir9NNcfCoTwtxWflA68+cAIVCBwUCjejnQ+uDPxVVWbpR5
G1cUWntw2EenWqX1ojb/oyBDK69+m8INxoZkWPpRpSqAijThtX0EEgSa0BO7tG/B/duY3KTbpEKw
mg+ZMyBakGopxQngyhmHZxKLTZk+HTXgei49lT0nZEss4EdFF2GSxOj1uAGSZVv4werqpdYKtIqx
cCjn5lyqwUPRucW2KVfXWnPoeOQ7QNOdRWcbtqEwLdizWtfuDNMxH6xcKRVsFfHfh9MMhuLlK4n8
Nm+W+6z9muC6p+R0ZC3ONH2S0m+uNIN0KNC+DPE27y/mr1D+veaJST6quilWyCkaeHAToDkJagEZ
5L15E2GtPE7XOKnUV5u5f9i/42qQlfC8Gt0sEsFxUHR5VcwadEXzzFCjVu9aLoJZuR41LtKsgn+t
VhcJRmKS8h3+7Y1XnoNhnHZG86ax4GLZ10YUw+7y6fVcz5F8IucvNix8lPhld5ihPWQAJReZc4PK
QQRAqJt9Ky1+yb1Vi5aVlBj1LqlceLldfgo5gyNrIQnKlkJfPT5VPt0aC2zHA5RCUtIeQk67wCun
LBAdP+R+b1crimDnJd4V6XSmrrrwgFWufUP5vxtL0VtFiDqn8kXcomxb1L6xFnVyAW+re5JYI+67
aUb2ku/H5ozYji+WbE764pu/71cCrlELWOVFNJwVkcd/mpFePT1wKDZY7uv+FwlHIN/5uwbNELyF
+a9520KnF0/otihYRWJmNn6tZczaB+nJGpNczB/BR9qQNyDEyJI5f2O/NVEUbCkzoRvq4jooNIT7
Z5PHxdTbAIAQ1FlVklZRR6+I8+uJ3X5ZNG9TBWyGOdqiaov2pkZr9Vnaqug5sbXPiPR7WpJMvcVM
5A+FQq8ZG9z2s4E/xgcY4wzPBWRQ7x6KqX/eGaQRVHzIXcKLp9xgaUJPsI11s31tIDsLT41elQII
5aHhllCMgq1yjAujLzDWnurVoaqeAvOzrGaO6u0rp7NMIkrtQ+SKOE9xoPM6J38xeWAJAuhhP2Fs
U8V7SY9lPOrTCeTHIltu0iBIyGOH1IwwjNJMzZQtf8Wp6634NvZg0tEjakJ36zzzLj2flMVKCFH3
17WlsnLe2i570KI9L7tGRSKg8Q0V0hwK+/haueNenwFYQg2pPfdMtmTpnek14vQqX2CigGbm99pf
SJX2UWM4qawEZcPI8GU8gG/sZMM4dmEyD8dBVv0ViihC90Y4u+FN48k8Y69LxQ5fhn+Vzw7mBzmA
Jq1ZwSqcJIZ8fPZnWf7ICN8ZWdUiGEp8vjw1dTIwYjI7hrfuonN15ioWbTKf2flScIIhT9lnP+Jh
IW4CTjegNz8DRBSe6xvlCGWnprYWWogwfGYbSbk36SNJn1ZSgQoVt6spmjjznB9lNjICeW62ldZW
h6E6r7qQWqw5sSHJEXku3b3/va3JOuR5Sol7jS9XGL+mfdVkALCOivOq5oKf8P6Po+DGdVF2kMEi
4J7Zug0/w3ys0lrCluWJfNRC/bgj/P7nL4WJ+ZHxhdlZ+80HT6EbLf27clrDdx8t0MyW/5qQqv4G
Js0C/p5ojLhA0pL51IHk+cAjbwsUFbGgQvRnmdo9EDSMYu8bbGKrJfvWeP8jrTANk8B1MB2dskNE
QFnoD+uj3RgMaYc2Wd0oPuwT9q9Pkx3wQ7LTk4tmFS1GlKIxZBIXC4scx/RmEMGLrkyqftardvPf
eTShmlfozh44/beHr+l2Y+E/4wE9k3n2MYUll8xFAGwzmL3aDzLHLYU478v0qhJxciDE6O8SwuGk
y9yThyLHme/KyqTnROWH15FbPbfxdFCmRxIUlWKqXF8ffuprH3U7+L43U82i8nk5ytNYWG+TZfYl
9ek/ex9pzARCnLaegziHjewHL11rmUkzCTX9//YlFsIx2aHgw2dhIIi33AdSFUzLiy4D1Du4aCCA
9xeebbVQUNk9wCNKNH/cI8ScLJhz8tQR7C8q8JziJDjIkI2mbocJNERDTaeFWZyLbn2vNZdQEghl
EjqQyO8BXw7k3IQcnS7qrotXOnjl98yoCvwOs3t3v+Wg/ljUX4pyz6qpdewX0RMYizK9ne8hUIUs
iUlgU7j2gJeCRcW0cKbp7OBzy/Qwb9PVcMnOc07S2tpE7qx/CUq7hCMccRQTAjU1IN5dmQnsQbFE
dF0NTKxFZ5F5gf113rSOB5/2BaNoYQkrmptLT/10kEI4G+kNzO64wV2FUxFpC7sfeMpunf8bIpbN
dwlb487/VJFxmCyif0CHuwx5WRgiwH4tGZ6HPDDtrsDjyBpXgJBOfzZcVuYlqplwL4CBBacy6wg7
Q2VoYv0ydsJ2qPkkgM7kQ/dOzLhMyFIlLwEOAYB0DJkA3ad0wWxGGAwoN89xvvkqaYQ+MtEwWyGX
xYwdmvbUx/CBNjisgJcf1Zv3bxXf9FqrzSS5nQkdF60sS6/5MymkPvAOeJ2OkQYXerY45on5FDou
U/v6el42LIgG/0X7ksApMrznK8ZBz5ih0vfduSY4Aa/cV/A1fYhNugW5ELauG3kictKxBmQqszhL
IOvBrqayY0bGOOLjaaZQc4yVZ+JEeLugfAXd17Hx5SK85DCZDGiTs7mc1zhlVVCNucp6UPij1LsT
vjhxFqaOK8S/cKKW2sFsXPlHgTJfWq7PSrF7GO75j1Lw8CAu5D165oTjRpuf+SuDg1ycY6dqLilm
AK2LR4N4kqPF1N0ZVfenLugtSaP8SC0kkE77owKVOTdfuAe5nMRKkh5kY+uoRi/QUvtsz0JfWrpc
a/SeJ1P+q3NNYFlDkCRb1oZ/N75YVacTKwhTwTjN0QKoomfOaclOo6VrQ+E5dqWM1qJSEmMhZFm6
jNz32qdwvXAgJjEGjiraBbwaUjb8I/GGIFLedYPLaY6PP2ou707m6JUClAnfPsX8oO5NQ749QRJK
ePjQ74Pg5XW4jwWGNy+1KUMlSvNoKoLKvA+FxIv2jd/TA+7LlGswDJ2tbpp31MXzChJMs4o/MB2w
DL2YQeS3fwA5LxIA4TKcySLQKFrFahUP6O9fJiVAxB0ZBtWF0Fn+YxhZTdv55XI2LjRep9JOcE+8
nU92Qo8adg8rtpghrMOb3Jfkwp6dw+h8CyPEVKLQxWNxjiegAQE1q5LEkMI10FpviG2o3Jx49/KZ
GgtNqq64bE21leV/fHxPTXHiN/BFP+9zhAcDwpHu0QxkgK04J/Un/eKIibmg1jdHlgAPuI8uFodj
hp5JNILFht3OhfFDp/p9QF2icn5roeJ3qedTJzrgAkT+FlqnQkanmOPc0VKBD8OhhPXdjpL5XdBv
+AYA3e/JHKfKbzGb1TV3KElF9o0yTE0wmwohufxNfAbM8eyEXeOrfqP6E2vJvPECz5MAcbFrhnhP
4AxPKoHqICK2RkyOS1qXGCD2CsEI3BiQs5ejhHtsmZrdBXV8YHu4oFye/wKE07/IvoJG/UHz4r3o
9JV5lK5TmrM+f7WSGAnyN9PCum7JSFfNG7/ptHDeYBML+HmO3kkxltD5bYOyqRrrE2qqZhMZNH//
4AO9zwDBLp54GVfIW729w4aWq07ldqO+s+Nl40yxTy8Hku2YoW+q+sIzvjc5cFKZNQApW5fnOaD9
+8nfyMBC6uF4bn26Z1BcuGUPhXijjGpOR5vMyxd1iI67ve5ELswkCcpcmlc0pmVKn8Y17JvF8OQi
2bsE9+cc+nvD7Wy2oGyyjm3G6nhvPv+TmGqYlGuKohstarJzZsDKKLBhp36acy3HNrtKc0E/uDTc
tWHa0ypOj3PdcyJ/O/OWe92AftsrM3TebGDbPLPmb4rt4KUW6d2nFbjDSkFfJQBcG+6yuh/gnEN9
MIh/Gpl6chKm5JL267S/UcGN34os/ID0sdQzvki5jnUxaHDVVm0BQZAJBXWGEWyH9+h4pEEZuKv/
IlFrbt6sO2yplG3nljGxyWgeczNFkT6XdDtuN9aHcnS/NZ6eF2r4PQGz8W7JEIpGaXrPqTEg2I5/
qwc7gfcqAaa9TbWP5FX9HKKznNlxmn9lUh9JAjclVCp/7Vk5jbSfqvEo1q+ApWngQJoyccZByDHs
7HTQUR76Ve/KmFBXSxgFiNC1FsQ4eUL0eLKWQ6qbsdKuVeWSqYJIiZFQ+rx+obOPBgwmYe1leN8Y
i1nYK6UepmEmbo2rrK3yRnuRKC5ECVXJPh2xC46aSi+b4BtDYHl5YhfeYjrNkZB7NV207EMyff12
Ghk6nOSGfR88N/QN10ewgY3ERt9+JY9Td7wqIDVrCW5TUTF3Pjl3wWTj7CDh6K5ewrORlupzxudt
aNBhr8rzA8wsvk900CY7YcPiozdJKMHu7L978n4OCN+T4ROLsIf9J/DLKQneVod+iu5b2wRAD4QV
Yl8zSAksgbfG5C75MRmBzNOlCRal0tmL4DL/R79C2Qs8B8b7TFk+Q0Fsbu6sTToSTSiWmGaFMfYu
Hs/+KdDEoPHExe8w7BW51MokrlELgoLBAOpoQ8fAsBbRZZ8eYBdGDHQ/Jhttc214xYFtZhPt7aJF
RWb7VSymqrRFrmUIhXC5U6PaU+EIfbYZT7zbjSk06Fnlh0+9Z5YYnOdf+0keXIpXvbUw6BHJTnfJ
U82mjbQMNgJnmkIQCUzqEGqajtr99prqpd5YgjrQaHx3Hp6/tRdd4TyRvSI/NAP4Dt+Ts49XUqRj
DPRuEBs7ibqo9p4Fvh5t68TJ3rFWTwc+EYhPMpIXNPaEG9NKk/kJoWKIyaXzlpzIuwvxTXBiYmTH
Y+mIbbtF+YGgyLBXQ+LtK2Sf8vu3u2bQqmepDCsM8ulBVgQGQ3NUNNg7xZogdYna+bo7zY1+8SAW
2kmbnqzefNbabqMILRHgQx2T6GE/oPYRanlNNW39Oh0fJ7nAnYGV6MZwGxBN9pGCnQUKlf4wkgLy
0ZS7jN+wDToHNFRkGel+cqoBuh05BE6kizO4GQJW841PpUhNTGNdBrdddQx9Zi+2eSF8sE0q+x/c
0jKrEi4UU5PEE0uHJy7taKeX6xOOyuliSayCZYSflt+KPnvTyev6yLqSgX7SgXwi1HfyTyh8hp5C
NX2KV4tMbnP++jJpQzM4/zQEDr6/Not/ZaRLOGAsT5L06Bacl7/ODvU+mtnRIz0uZXNgkdFfEBLx
ca+Yu6bBAFOIwwrsbx7bRIgidzRfWW/RFh9H4dWK2+qsZI6OFqQ17J0LQcBXFYWX6AkLPYmHV67t
SegzJS1cSTWqiwaq1zITq7DdEA1HnOvzmBm/AAARP/SELMXc0NFGhRbHoOm0xzE3JKVgpErKgSW/
6QrT3fZnkHI5ce4H5RDfWLJBe2hzfoqKMXc8SJdtxUHDjYKfCr/HsJ9K48CElW9V1hg14nwiQ4u+
RG5V7wAekxVYpZ0XlBVqjNStUfuhXg/IqA4cZxe+MmOeTQRbqZ3S50piRb9mxCKSDe02ZkYInSZt
TirrI/z6LU6Yh9q6jQUs8VaVvO7sJCfc01qwl8CgJhAPoOaqLPkzPk0L3bktyhdCY+tm3v6Y8o4X
3M+uIez/t7zN5kURJKKtxHbB36v4/tPL1boZuE24phbYiBn/BL7UuERl/ANRwq2ymelUV35YRr1h
ZKeUExQO5a+4LUSoQje9lHAZZsNvSUBfIxIsbfPerRpKMj0GDfJWll8AJWLje5ndh3TEj3iEtz8I
5YL1lL/NwWAQVvhiUw1lLsNL6XoPI4bp4DRJ/TzyG2CKxpl8Ncy/0nKB/CyCzJoKdopcGRTEk3AY
B9ipeFMxQtJLaUJt7QafB1DnJpPAmLIqFJ62KZG8JJ/Pk7gVRD+VDI3dnijI4OhJBkKRt07mml1U
1yBhmYqq9HqKFc9fFhfDkyfWzgaiSFBybwTHIU5i2jasCfBrfwXzmawI4GCrR7yUJ/k68Sz+y4D8
NJDjw32MqDdsrx9obUg7gBHFYYKjyL10UQwYstOz9PDbqrRDKOtDLipeKF93ZIn7Q9H5UIsazoXK
Rb+TixNH2dpuFPxkwNM/N19AYcJcQb5/7N3IysWKmxsl0xNPXI6EK2vOrVq4iY+fyJNyrzvw5Mg5
g8Bcfj6viKVm4Lnqk8Pd2vKokK2wlIYEfRdfNe87G7rztBrHBz66pwap9l62L/jUkYsLGdbYOu+l
lxR3O6+01paHp3Iy87Dy7Ge9quw0TxEkI6qT+mq0On2Nu4riwDbLZEhs+p5NSZBJlbxb5l5FsD47
EEZPa91HlBo153Xmwb/0ykx0JzpoBMQy43z0UtQ+LYyjcXo59Zh3sMPGzWS8ZMnpNFXmyqpQxRhl
WdQY6LjGrb/OI99Wo428fe+eZrqHvW9oKfGQc8hFvvclsHXAw5iu0VEWHc/CgtxgJbnxVrBQIcG/
WVX4LskuafCWkQcBNxcT7rhEFIieeYdpmzNrtx8LvgKztM0tEZf8oXKzHDKsdLnWSCCDDvQez7Lb
RSdDE+0UVAdNpEvKbQkbrvIH5dJ9B7c9ExgOfLgUL62AADdkgfed2fo9eedsIt0jsoqkk2MmnXXY
++kA8NzQjxqTY/xaNnuB6ZTIzDlYfnHo6BrEgYmgnQbLw24BR/P2Vn0k3h9EnwX/QYBMGDM8qtUf
oc2kPxEk7/bmt/053u/DXyAKAvq3apEDAGQcJJkpIv47F9r81xyxk71YT3K6i7Cie2lUCBkKMuPW
KKOKmi/IG0I94C1Oct3vQ+NERxHfqfO0WdNNXdcd7UR9r6AGiwqX9uwCRD+SV0cPrerM2n5mbcxD
qR5qbOpkJOE43Ytp+ngh23OUSZbwTlO5k7V5TLv+JzBXezyVnbeJKgWZYm76YF4gUf0lQGmGZjY3
8YqGI93FFU5nKA4hLQ5QYCmpNWrhv8mQbDyKNr53xMMwUbvaSWgZ/mwUAAbPVJJaUUcqHDOu01aA
+0Boq23eDRiJNFqNVxE7neWDb7lw9XL4DHm/YP/zj+edzT+xR/x9a2a8OXe2IFnXmSZrgrH+rfgS
nAAl/xI/YEteXgCQq91CESGwCxfDqGZP+K4WVypKOR6FRHesStDh8BHCVYsgsu7jONMi4X6tgNeK
sB2dhQUJJaK9hMdRX/U2xei3FD3RTXhOsm7/0wq+E5o6G0LIAu5DvuN3wT62JuoGS8JEhBTQSdQu
yHmX8JgOwIa05odiwqpfNgf5fUJxIE618e1NqYFTxpxQzU+0HNKVYtyOMfdasp21n688nIqwbcff
QUHonOb0fa32l+Sygrv4+KXUkBWruJSn/WuCP8pDx2GVhXZjnG1ASuljjtkAZQQYYtEObk70bE4F
gyb7PVvYQaHgfavob2BXbBd1VmaH4Lz3QjzqunAQyzaN63j4uRcvLGLxNsJBR3odgfFXgFfZnbmP
rFRPl9aCDudtIowA1JDgxnJst3JWh//rZoY7WKB9R0Kd0JibRsjs3rTO4GovHAeR0QUojS1YH+Pv
1MzoRYZICIFO/gA+G134VnaYVr9LFmoy+uCoSMwCWiyVRg4+deHMsoMCL5WMOmYJrxoS9YMP61AX
+ZunW0q5+FcQeBnAwLcYgsBiRdxLhAO1yX9C1rNdMLpl1b4g8AgNq44NiHPbU+1CVpLGfRErr9wE
C2DJCnLiErSoLFps75viFeJEHRtCnVtpHAnM0TaXq5z5P5xzVPx/qkgDvxkquIbYMDkfTbwsdqB6
iPvIZyI39ksh95wP8Y5J4EWfUTXQ77Xr8V+JivXqbwnAw7iNXMb4egiP9nCS/1qNJi4Zw3c8rCRe
q+qjatOXVDMKbnfdoS35uxYsWqB0h2TZm8CPMTyMvgHoQ6d2sZnYiSQ5cDreumyWzExuNHTEgzMV
NkPSCrRgIffyt0ecRrcO7/ljPifjPVOey+jlGRuzxV0wvwR80AphdJ5HqvKqG88IhX/LUeNKY5L5
u9MgemVV/Ex+tmzMCf9WGgbdLGcP3rcP56kWph3uplH8dW+QYXgbm+8c2JIVvSfOPk2F8qrag7df
Gv5lp7c7SU28BPKfSnzvl1fiOzlVMEt1rzbXu62TSzkIwrle3XiNbLkqcu/uqvux0w5x1pDIRWrW
WjpChSFgyEjEz/i9eMlK0zxzY79YlcagcXexJOEfEK/fwythKnxjLZfR52jMaS0YWeAdmdKopF7v
WFFVn5LKBDLV4jmh70QyGWhmGTYPU44wX/GrGZRuPOJYG9mmFhv4xAKFU7UpTqv5EErKQP4dQ5yg
c4qXqZFENZ5XztMmi0fZ4iv7HIwDGsX+rQ81vxZh3JKpllKFxx4ZSM+O70UuD5nfSjp8CzwD0oc5
RBf91u50Uzs5NOmTH4BAIasT5+e6y0Skd1W8lOTld19Vc/R/pSEcmvvQFKgDYoPI+rzb80l+Pg9s
P4IddzqkxwuoPjvCKQgxMlLLqU6cvrVXlLbF+NqdXvzfV16+S8hPohb7fTqdfW9+EmH7Nze7qRNu
6SorQf/EGApFYAu7JvCw7+rA6pEoC5szP9NPTKp6Xm1eSKXC68kWy7X5PfT13agT/ye9CFA+iYXr
fgvsxbsOcpo7gs7KxWtvFaZHIzT0T65ObJN4xyY6Lm5yJX5WGR/+KSPI34TxREclMM7ltWCeZYgp
H4PboXuUaJrRqgIbUvAn31/y42GFT7uvmGWOCe5hjwokR7fCso62oOGsm8A778jtqppsFceM81rV
zzMHSGY8ai1IPi0YfSPkdgcUHs/QXw5s5oa/gMkY9rZG2x+jKpgGmMZOqBsVYP+IjjJQtMgcYVve
iLe9eK3xLqG6K/GSqOeXP2Sskp/2ptXX3Zdd3OimFPWDOQtVKQTzH+pmefVXa4b/H7g/AelXV2So
sk0ms5tTclufKfkZoBctUh5GzswT4jB0SqKhVFwzc66dW0OInVIp9RKoCsBEEL7RkvryEschTHbf
ZBAESK3PuH4QUVkkN0xuz+z0hau0vM3byPbTD8qg/X26lN3vO1MpS0aD+/lky5Y5D/MCGGE9WE0I
iotPbWMT7WJ0mczTFMPfFSmQ8sN5pqiXTFkqDGsRWj7kBhy0NCvUDZWUaLHnI9RcY4Wje0KHhAeX
y8GrgYR+O8Iq/q5w6sP/YM2PuOp/dboJdURXNqsLEn9d0tmSvuSb2cmZuh0b8R7IFojfUH8wYc0r
JxNYTsJU9TQham1BkVmMVbhyc6KOwIIGKNG4a8Ia+WnvqN5+TnOheCs8qzDNB3wK2yTPZ1fRChLC
u4H4sLYdJ8vDlfF0mcmWu4jDFjqr4PHF8+t3vfndfhUkvNWgqUmjGMxMmGkyiDHYdbOIOZyvmQH9
iIbzDajrTs3oQ9WkAzGuqBhnP49Ju/CM5PMgSuPr1GJQFlG/PFicWxwjjafw1I+QpZ9LR7pYGqsP
cAptrIdjyd1UwImfFYitnQJQgu8S5RMP4xLzYcwigV7xdIX3iYed51wl/foUtEcBt4u8qcVraF2w
lE5cENVWW3bIc6qIihwKwcW7eHgONIdD7375moo0Ek5nimeLvU3bAESZJPTrn+EdJbHqWJrygpmR
q6NY/IVLTDxREj+Ve0DSYTQRRHoXT6ibLtnvZrToiBSknAbUBGVqQ7q4ro8Fwo0ztWq+G/MgYzYv
cx0N+be9rytAjQc2RPYWvrJnVlslf4yQaf1RavrjrBOl91GbmJC6kC2jiwYVA1r1K79JesQKH5mB
P3q+ZKy6LA6674A0vW8At1ti7no5jfao1px9R9H90Mj7/rXz2EpGe1VL5BAFCAxwBNEXvU0JksMp
yi7BrMTDVI1adfWER7ZPNqxZ9Os73umoP14TRxldVBcwgwz3hfeVazwTripe353XIZ2Xcir8oZ8A
rnrZbphGaFf7ZIjD8zAYWyG/OXgtlfMArjDEevAg3oEFI5QGTXtYk8ekrrqxPuGOE8Td6kg5jHl2
GHOSTO9025LRQwXsVWdlvR4Uk05xMdGr+2cTBUeyszpkFKp39mGwh9kggwro+ucVBxWlG+WDrurl
W1CKoj6WogxvycQMUZEbc8ATuE32idoXPAhjaXH5V7u79AURQ/wvaZ+gXlnaS1H0Nj2P5sR5VvwH
qogyqKVXgDQ0SSqEaQOGpw4URq5FVg9GHt7iagGqbwowK6JjfgSE3W7pb+2SpIo+UWo3SsE2DwJP
Ug8Z9R/mDCgaO+0wuFYceArjzxU6afmUljImjN+foUKtylifT0draV14rE4C3wqoWpoUDO7q+NzQ
JXU8R+HmbaBHHWA7VRhinW9SymJ6TGezyryPVmWAnWBTENAcZJJwWkz+9z5VnFI7aYgsctZbN0Uk
mFk0+DO7tQPvLeJpjWiCqxn6ryORjNtppJloLjSuynl2q+FlTYNKK0Fj2OD01vSQvROPq7e3x2Ox
5SBkOneiHPudIw7wHIN9eGwvntSybjpEYeBk+2K/a5UzUH18GHxx+RxfWwytYEFSexqJ69rWTEEG
wReYvP7/KtoYV90/I3hEiUBWGR6IRepwlEDhtWOMM4hRTvfC2ffa1SbI0pKGVoclWTURqQImWffL
VNQyJ0YIjhM4HL6NixUkVSgTSvcccyRB/3hvEDi76CM4qWL4NE3sqR6Zqd8CAVveHrLgIf9puE8A
0L23tCfz+Z7/ULzvdstZBYnIXGx21fY7rsoT9pQCvbLaNVSsBUSUU+KzSXiTjN3wRic1xROgRFOr
asYWogGGWGkctKE8XnZnMcLJfJPhccNZglcbY1BhAqF3D7q/5CCxcBb2vv7lWZ6vMQ3XrdkY7SVW
NfQWBykyaOYHb/eGq7roAzKoN12QqkIqM/Bcquzr4sDGsSurknNUEAo/zooy7c45CPxgUq7xDhjc
X7G2I3sgaAQYDPbZaFlpL3gKQzkmvrR7YZWyjLOJosq/zkGiVYKDg2HN7AG8f59xpB1p0C6NJSzW
eif9ySX1qJfBXOn8ex+6Yb5ovmzDrJJ3q64pP7T8+zesc4FpnY1zctOmsOjuAn4IOmRmM++UWVf8
xTWxT3+axDJzbZxNkVKNTJGs1/YmZE6Ux90LuUbA8ox08yHyCrrxTfkKWfJRE+xx2FmCFFvQDFZM
P1Cc9gZDN/6xYW0/9qk3E3HFg5TXdWDg47Aezn9p0UBLgu01ykaQa/NNBW2j/k2sHQRxqNb/rR1b
EGS2/56lfrgUcemJIlvK3wpxleFfdqNe+2wMWP76NqfE2rvTna4af2y/hXWNEr4uJxu/n1Xup7/a
H5UDNYLeBiGVGnkVtc683290tuZCCu5E6tfOQvZobS3npnwojHA85oIwlpEA53Tu4UqlPYsYSQE1
9rnbqE06HCtnR8imvz/Vvv0Atazgka8gAz2mBn98MgThUx4/m1ofWR7sb3013PJHB6lSJC33GUGZ
XMKSjGihbkHM+ZEjdidpF/U1PMgeSN8Y4g4PdpuK+Yx4FiffY4Dbp9w/aj8Ywh61+3DrpBEz1AHd
wCGULeILTnGRS0LM01TdyBc0mfOz5wX4MtIkiWLSUvCZ07b8RXv99td9MgWwq2KtBaYmkiEy7uWu
0Ri9olupJs1R/H/GHN4X3/gIz6jMgE07/4jNGFRfcCm8IwkfSKx7qvmomtoqOtzmtlFVwN61vLzZ
ZV6HP2Ic7Ndj+IVTAFJYCj/4boOm8ZXn53W399veel1uwzAiWa04EeF+F0rmcA+dhBE+dd/lDi2P
jKHxRejPkVEI7Fm+cu5x2wFwaU+kxIpKRGrWj1V1b5Ym+cJ0HMVe31WBq5XrCagj3d55w0NQiyPV
2Y+VsH+J5cFuwkD+AsHbKJA/6cmjQRwxDElwCHTjEwRxMbi/HYlGB10mj6nBiHWT09XFpwlmaRIX
gWZrAPcceyCDOFkYNR3BKDQS/lSpgB3O+Pp5cPI2CH/wFgSxIUWx7SOm+KO68DjZF+FBGjYLW86j
jSbuIkNapihRoB2g8KIO4YtNi4rqCg8/RR18dQ8yzwwTyxWFJHByLoISpnJ+nhOPMcmwfkDbJZvw
LYfa28arwYAWxfv4qobUzgRR+0Z23UZw7fuTr7ZGsJvLGmhOOOv3LFY1Z1+dfTNZizsLiuBTHdFw
l7gsc2+qoZQX6mbRZ3USsx30BuZGsS0+A/wJM+AMJf2R+fb8hrXAm+DrqjsHXlFLeNJ7uZrhYEex
Q80PSPaHhQ7t4sqc7OjAn7hpTmR/ohZg7uRtE9eA7To+tdDvQSykjxYtyti+ZzHvcDzgi1X3K78Z
pxUtBnc71Cy3Gwqgo8ARea1mqeHfxC1djWW9bQC+zX253/n359WhRjEcufANGDCnmQf2QA8XHDDj
fa5ZgD+tQcLnDzico2Wnyaq0RfujDSNYbakXlvmYNkqvZnxwk5yNSeQzu4tYo0uI+PnLFhwztmrR
I4mnwESvP9t5QK939nIGdOFeyaeCRrXVXC/1BppScs4IiKrtx54MebxWmFMBkGtDSi1dFEG7tKP2
pyChft/bTEp8KipNk3MUi2c1c4+LLiE/KeuPA8FWiCUMvQdWiwLeQwpVYnCNCm1Eib+6Zek93F9S
9tBu7mYXce+v1x4Riw60EPBYCcws41OP4dd2XPX+Mu1nOp6ezVdaDzMQD2Gwb1lEbMBYeO4xjR7O
IuXLOf03FOEJYMsUid7z+B3tcZPk19LZQCPlSzoqe/H19Nyds9RCSfncSNNtmnb2a/QF9JIrblRi
5pzcHG1uKe+wUzghw64qBlaA194oRqwUdSwjsvFutH9fwYVlLQmWIsz4swlLWzRD1SCjaevx6P7+
k4RCSEFXQnqsG1kFCmA7DZfkPvNpTh6iisiUZsA+gcFB1RWqdhodMoXjR+Fr7ZLuQsnPIg7yVlzH
ssVjVGDolx4Vxo5ZG/1fpuiLQ62qN847mDBD0GJ76Kh9mHlHo4Q3VOjmd1dPRu+zSPYL3CfneUvf
Cmxd//EybUXZ5+ZI4G26qmFZuT1NeP82LRWO1XALmUk+kx0mrWjZnguJIxTbonos9MdGr/uJefjY
iB42DJJumk7gi6EvemFNXG1bnInvzc9OcPJyya7AAFDv/Zlgxdd3FhbvsxzbPXrOcRaKFB/LfYL/
spAbZe8HF6TpdF77jsYN72muKHb0pIcIjoHDmxe0Bn0s5Qncus7aTUaZRSKPN+6fvtl6l2WsbnKf
WXJqx77I0dBUqgr+xEOKjRs5m4oXUnXIkXk1LfeZ6XETGuA2c22xOUabxVGSg5Gg8jzowRl0Pdoo
IpN+cmFXwsKn4bZZTKi3YPxMK9aAx7QwIsR1MVADfL9ABfLK1M+IQfpeuzvZFbrSZmzpMJsLE/AM
pPoXYehedP5sxyWpG7+KpjcTz33CHAYYCQ2TtpAYlwf1SS1gk6aDdWoqHxb/KQW9dps4hxPifIrm
MJ5qTD6k1JnzZtcfZNwi93at21eZk19DBhEoU4DcN8ojMQcqYNvvG2JqytysSrCxUWrfjCdIRFFe
y6B0gzyx0zPM71LpRoBCgckAmEgXWe6PwcsILDAuyA8hWiPzkHo7ManrWuSPtOjGwRgMvOh8uSxi
usOhm1klAC/t+XU7Nt2Qu0H26tEUEYUdy6MwX2jKCu5d7MTkP/gEp6/KAoCRVkaLTbALfuBIg3wl
GbkNl8PwZ4pHzPBC/ACakgScKLREkdJDg7a6ArqvrmTyN2HlG4eWs6lcsnwb+oCoQi4LuAo48aZa
vInlopTicQe7abEDTty6vVJaPTtW32CkssUH57NyNgGVnwDBTTpz1tisWPr6j22yQIlW9htmCOXU
ZSoCYjOjk7Uo+CAERLL6CeQbh6G6neK+mClMpF0OHiquGENzYuL8jEtdzd0mgs9HZsdhl/3BEXWZ
cwhxWvqwpgjatO1jp2dYD+MNuw4aOcMJZLN4yVvqcpW1DDkqGFO7sQuFdpcougtB6/LrHShpha8G
0vNMUSolKG+BEOskzpXOExl3KRwHqd35PqUJjHYrxRVpyuLTEXMMFhDy6zmmkuIWyFWy62BIVOfp
sOtNSL3yvxQiukvsryuU6t/H2jmrWOs+ybM9TZdSmmMVLvtHPBD45L60L+AF9BYgmGGdqQ7MGvJu
tCGwCEkJb/Qqq8NxbvFpeKjsJfu9BxyV1UqLtp5kGVks5KcJjac5GlP2gbkq4I7Ac5b/IOBsZc7q
Xow5KyF5k6VyFZ8B5VEID69n4K8svSGRZsnjWr+MxClSSO7bEs648fUH3fiSBylkwOv0X4CPf074
HGGDkvRP3iGWMD3f0Y+tkeJGhwAy2ixanOtu2q37BmILHJvn7CnbJ/mfrO8p9k3a04l0uOvPD3tD
PB7TMR39DTiHAj6mD1Dx1+Z/yDtLSeRJeehepcdxFe6AqZ0WwId8zDl/iev7n6W81YA3IyfDRj3V
rkcdSJFi34aGC1aKNRxyrL+38e+ot88PIpjx3YDH5CBG7l2BNN8tQFttG5eG4N6/RCB0PKGg1fRE
ZGQLA7GwzQXBwvLsKK+JXmmVJCm0jlJSBUnNfI2BxnQ0ie6PpHloI2Ghx30HMzbxTvqQSOsz8+1L
dUnrYuCazxsQBiLanmIPdPn3WZkluYm0F6AAAsf3djdrPkge5xI0zWOT3q6Pil96sennZ5kyWqE5
dxVHCOuFxOBrnKnlfOCiw1eU7Q3TRw7/DFquTprj8cWn0FtK2YDWAQf0mkOpXMhGHUSqsKdz7sEu
HEmFVqIYxD+nzMkvEbe/yIptN1F8ZVBy2Q00ZwR2pHT+y0UtFMPp8d7TKe9Fq/5CMLkxkk+UIHIS
AYAMHQsH9g9Mc/3U6tpsvysb0311xGjud6TiTw5zk8NzmLlgodMIpFsOlsvxqOqmVS9kU73u4e1B
JngpeA61c3dn/X4qCvEAw1iJVh6nkqvr281RBbKo1sWCl4ITeyfwRIeaFoQDpn2aH1PWiS9Td5yp
1+MVZAH5i8PYqy9LLCJBeIF2d9X4NZQMq7JzUF5hDtoh1bzaYtnGxZwjErU6jQPvRXv2E8xN1HRE
n8IQi8HLyL5XFcRVwJjwn37f9bT9mIVnRfzPf5d3fZlg2SgfMCZe66auzL7FQHEO/UqkYk+xfsOq
KE9jFxkVMqRSHPFsqFUOlhcPir6unm1YJBjcvJbSzTTTE2CRoIM2+++rhl0KmCzGSG6W5gvg6LKA
SOo/vVA9OsqCgKMW32myuOujzyd/N9wvIvePYHpOk7ZIJBa8HoSd9CgLhghTc0hpi6xWOmnmV8Ej
qSjDWt/NYEvvoYJ7HCELAe5MPyWg35ppfjaT4uimU60kTKIPsllbrX9b5m6FoEXTY2suygeifRZm
+fwLxdw9Irztg97603EsJxLBvyIZwIdAN46AcCcVSmZ+s/kd7NsErLQHA4kfC6krW+bJsSzRyMLp
NtR0JJup5Hz7Di48uDDm0nAlBH1Pu0rSZnQPwqPFMte0sAc9Tn7oigTpidpaddyOZecIZaeI67eA
vQ2Kakn1lWfR74VSGg8EAFA2OeBWKS5GQcXtyJAg2BgaphqXh4u4sH/HXuDt5loIFp84RvW6nNdz
jiX5SbNshEF+xNC+xmMTgDRWDAbuJDsWxTNCEGXCeSwiKQlJj37sURS25bjv1BeKEnSZzUgtzgau
emg/BnFEsPuc6R3vAwNCWlPm5U7sXq4TYb9mhFw2gXZhIC9HJ85Y3Vp5VDDCsK4xaKgOiiWa6IuJ
KOzmalc7FNFPrFUwODE+STUqcLzEcSSOnvRNIFBjndxNpTT+DsNxwU/+xgNLEetsmFH2dpjRwfTr
Y067aBDmxuDVhvjOc1R6RfFvWKT4bHukqhM1qENu5vOiFJmQMF5+WITKrcB6npICqdeRLrcCpFNT
l9zfjEwLBQevS72npgnkFO7M5O204J97dHWYaBesMYvexl5JO3yoj32QDymCfDks6Q4vMiGM1dzb
jkzfEQ1VMHqHBZvKKzh/uqr3yjm3Q3wRpw1KhwR6OzVo8nm1R/f1q6yJDs7jMcPPgwRppXBC4bcA
6v8pfIO7AJAZaIe5nwPhRCR6nTLYIe5b3TW1s+o6lf/1lx6KZNuoZv8AiSdMnb/btHHW/EvZc7Du
l2qBHGVXVNlWIq5rPLBvyCVGwdCR3hAeGCLn4auBlq88w5MVnXNTZNhlp2m14CC3WuwzU+RYtdCy
S7lpsPN7618BU8VJDdBe1YXSl+guFKCUefYS2Y7jRlDvXNvpOvlPRu6XzLXda3OWnH9UHsfTyu0g
WkecM5Mjxpae1kXY2T7s82wcPqJUkrr+m4GG5s+SI1xjIJKjJhkGyeQNrObMN/WBSkOvXRXA9bII
f5eoc0i9Qw5psFwXNrKwkrb5h2CTWAUTRl2QBND2/vmyp1NCkyE038g1d7BeVr+H0PekjgyhPLda
QmzBU0IpZF9lMI0S6pqpHdwN/FituHH3MIQ6Ua3EQWYOxgHFLeFGjs+V9KIfWRycPykYkobAqG4t
REDTDsD90K7p97oy82gwG8BZ936UvAYiKksXj/GAigD6VSZvI516/4GRRcL4A8/aKWjUS42PjhBO
3bEX7siMm1UsRJO7ccu5nVh1FhAitkSKBWb1fYCfdVFt2BNG9BDoUc1c66kl8DDsl4tqk8StpPzR
WjcvQ3oqLveVDrP4SexW5mU2ziaiyQnLD2MfGQZQlMxRrPMNOboz9YCc7Ol3iY/HcQf+E45ZIAVW
JK/VK602QXwNSCgcdsXRNHYkPUyzqP9Z49FdIwfXRv6I6bAV3aaNvL9uX3gtB7llvBejZzk0ESVW
w+BX5CH0+YwqPDMWuZBWe5u7c6nTwA+2mFB+xSDuomzP0U1xL172LbOuAXuU5i/aoUXRl+KgsKBf
tVIRaYNY5xn/VD7KO+T8LFVMOat3GkNF+thtZ6rSie1Lemu+zUvMAgtE7vo1g7MWlrdUUGvXbruq
likrrvkpGz0uGkeX5NGJVGSTKvqjbi/91Or4V5RYGzx6Y7rUdmZK9lRa4aYyoePFoLPsan3/Mz03
hd6tnVtB+k8ha40hNazWXwAYSwEgykLtAwm3id7U5m3jQcE0BF6iO7VNCKpyZdUY0AhUri4/mA9O
gdglFy6WNMvzYFCyqntH7DNICa6za/kL2Sy71xYH/Ji8rVXCtJau/ZbKmFrVfQp0RuLZD7Yn+saH
TaRwJpRaslhjpAyisGDXmOsESA7dla5f+dsles0p34EO5pf2uO44BVaYSPGfY9zMPL8HrhFwxeXY
KFqND8t6vnAb8x3S1UQyQNTGvt3ELEnXgGFGxUJygk1GDXx434cUHl2qIwi2vyGNNN+iNIUA1qAn
H9AGSW2FA5SITFpwaD3ZEmWvvCLO1ciDXmDGa2yxVV6IhLE5JfPz2HO1kfLHBroJsvsZYHeiSEuo
Gjc145+gfGNts3vyS1DMTReW2Bs2Qn2kDoQZrmKKQa9Or5lTslNdrQcNB6twvUdio6XY5336W0Ci
bKS/WqKKw6UyRldam7MyAMCUvXWrxM349GW1xcb6j5ukwBKU71qb7BauwBCec5d79miOzKiNVFJI
V6YyWeuYq1bAqAAqkvVCh4PHc7gXQDPJTFO4EHoohXh3iL3LXDZk+QBLdWnznY9p/JGD3XmwG2Uw
U2q6HUgNTdBefnXu4tSluvOio1IECsYMPKuTdHLMli6wx74LK3j0K6VCmOcF6Rv0nh5ctd4baxyT
6atG07Zak4QAbbq1wfnOOKPo/YKNPGDZAi1YxhaDRFI2kmAHl3Fz4z+NlikAaWxNCGXY/5YaYMd1
p9z2bIcbG4NAYY0+z0u9uWE2DK2N0Hsb76u/e0gP80f6xieavzFqwGf4nmcKh9lI67Ys6DQ1gC9m
ndRAwNCytXDupFsels4PxtRkxL2vQYz3l02tDciJpp5RzxHLQZeygDOsLa7srnjC+4CItCOcWhHs
PQ89EFinMDxxYV4NJRfHW6UrdLo9HiE3BAV3eHS0WVEPUznC0MpcWX4N0NGOtUg+58jrdOKGJmTD
Ninz+FskL/cOnYdVuKHISFWDKe2DC3Tic+bIdiH22EYRJuNVJ217lRXoLNVTRLudpXfEqKFqB7gW
lzFqmKccfYeh1v05KlvEV1kS2YCCpaD/9XdnrosNOohLxUgofrMuLVAZH73Nd7ar+Xvg8Qf2ARB3
NyCJ77k1EkjujvzZzYCA3z/LJJWMCM7YAU5Wvs2d6szerV1jjMLfvQnP1NJcYoX+xH/gvpnk1OKN
SCYxMtt6IEFwYwhPowaFKpz9rHf2kRaMR/0idPVLWxYqy3rp65KY8Bhpnzn6wfVcb9r1tNvsFxjv
cgNvPB4x6Bkm5uD0AqU1J0wx0JIuknbGFbHHXiTUoB+4d1R7kxNk/k0WI+Fl1YWwkRDQARQOPX5q
bXRBBHrMTH43bYJoH10ToxG9vdDtW8WBzy9pckBVDSrGlfplaCXldA38EOZJlbL12GhJuTKNTtH5
OTSIIzOKrJIrS2uZs6mfuzX7FYe6HbPv9omRAfRp43fac2wXc8cQ9YJePjpr9X8HkbPebukwX0+N
lgvmFcNDqp2ksgEzSNnjxml3izjZYW1212pQgC8BRRPJyibTQvV1zZrkkoJbZusZmUFQuIvPD6xL
gQY/efTWnGsFhj6AcFd0qYSFjpfKW8ts1Dzvk6pQkHZX0oeODxRXsGojpiMiKb5VbbTMIP6ZoBrK
z89X7O2d45TtU+c4rkhZnBLo2o3enoOeQabq5RRVRFbdsYotDAV16p0EqawV4TectnhmcAMufgE8
PoScFTqAE9OP1CmBQZVfS28kLGDcsD5RoBf19M8G/VlbM5Qhz/Ou26vu+kcXgKvzDfzhR4ltWDl9
FqjQhUKa12kphxJ0Qrmp+PCTjZU2/AWpvAcPSFo0P9SPjPU45bSC96qM3R7smtSMtv7PpJgrxHLN
QqkmZfwgZdo+gRnyxvn0G2Y39v+yf4aX8rQBVXwEjhXjNxEdbSrz4tipMKWNED4YGGsJmJCyyYSZ
yWB+5I2q64t6Pu3YNXgsX2z4LnyGoaqK+AHmBvrPOfudy3evvziBiYA57cDLOMOgJUzP7l1l/U15
jOvA5fg9nZp4mUbPvOuUrkoGUn7BxefEazPXxsr8pFpOA2b1JCcC0kAH5+mf4vNbk1QYNS6AGSDU
6l1Mi8KAwS88luOWHRe2sNcAkT1RFoYfzwTT341ll6vByXMf5O1CdRIeHSc05+mfyfGlWC1a/bER
RkRFnUIFHcaDdk2GDnCAqv8RcmhsVEclkpL18DZRDCDbOrKyJUflLOeX4HdLdweJV7bYWKkZOilC
mSnNTHQ/7MX7EV6VHUwzvGXzZUn0G9kIDhlxNf63s7vSEx3nnEW3tgOIiEdbITNO3g6Ujhd8jyUU
x3Sta6WUBZoA8WIy2G1/q0INqbmGMynwX98oe9S8gHREWlK0S5iCfJLLizYkzf5M6kIey9LC5z6y
/Q95OiD/jvnNc6Q+X5dkvQ+ZdYnIddr/h3b1uYhX5uCp2acQ6FplKj1vNNQ3ZeE9dnSO0cfy0hbg
V6p8riCD88GubOJ92ZnrNFgYCWjeyiv+xE435dUAGovwrYcUPRhA/+x43RP9I5mmvzNO2At12rvg
TyIDI2XmNVghqT6r8KXNJ6oa15+RY8nvlsk2p/3EJsrqKx9STlBKzF0gkn2vbX/hRMkoswB94Gic
XeD5ZK6syeJ3raE/xr16DpzHcRWEZW+S2TLrgxBkodEqcEYM3tdOehs8OZBxsmVy9KKF1qDR1sg4
2BDngev3UcbtN7WcbzYZAYM8EsdyTiLEg3qg7JZeILh0fwnClA2Yy9pck4PueoJAZEgf+mlUXp4S
jkDCKngrWwP+udTQcZRBH7MhlS0ujDzwI2FQruOkUWwgSYO89mxVTOqlW7Wzm4rlrB4l1GvMB2/9
9eLXH62o+eVzboKfpnuqsNaIWiqwVQhvPWd/p2w1/vXCAWn/jUbwjjLOvwLQouk64QDg6v9ZaGDB
Vf5ndCl4xRAdHM7AsfLlTlfZ0HUT1euHDxvhyisdWaKyQ6Am4QQEPKPXqQ7QxKLD7U8hnSnc0Ti8
NQIF55M2gbdiWfh3eYUH1lqYOiA3rYm3n5N1/fu1JrFP8lpx7WyyvTkBnC4d4HJAxhNwLe40fZfS
ygaKYxNyg7AuVMrjebWeOHuAg0MtwapEk1TIfuWL43keoJQ4e8eicZ9fqJ34AB8X7lZbO0ocXt6f
MkVMBjR1TLobp/42s1sXHf6p++NZr+2GEP4RMdgA7gRwi73nVzKgWTvkALUT9U+2ZOF87CrOCio/
SeG1quHGxuOyCr7MSZDYl31amQGkA+PzQF/esx9YPZBthZBQNEwvLXLUpEA0kfVZBnBRPpGDMcOo
tV2aOi/OVWQMUS/6lMEF0knlLFlUqxU7J2yHkQSN1u44FwsO7ja00aj9QNI5QsWgyKpl4lwIhYs4
8SnuhCGOwLqf5yofPQxWQZ6XWP1fditiMYEYOHCrgGc4CmGhuqIs/HlJsSJGa1B6/mubVBMZoedK
a28Ednku8ACe/dNd6uEDopJEc1zbtdsLJGs66QSdB9n+Gz2L8TBNQj4tvG8icrzQIrxFYGwObZQB
olae9VTx3+diK7+1qWZaf+6pGg4712I4aZgMf0j6N6hv1nfmbB64pjYl/z3gh2wT96bmt01AaGKz
NOU3lorEJWVHiWSqy6AlCFr9BE4Go4MFce0e4CnNLDlNOQKv1tnTW0vhJZks+F1jZ4mJNi9gFzEY
tvcdKQ/8tVfadvRljoIY5FTwLWFRJvKaTW0x9JcHJiK9B++nEJD/2d3uERGURG3EeozRvEpzn0is
AWgoiKo+1et5/N1P9uh6oyY8CgZmSASQ6AVj41t/YAuGQbqRNzV28SM1jeYTfLVGYN6tj3EJp7ef
lRtzypkL06ZsyYDGp4mVlPtoG8Q6ZiFVFioHLdttp44kzoWzaoacyrRSGKZsPiF/NMJ9xdaH4Ixq
+mWPgythVdPxbQGC4OYMMdLy+KJqXvu8TO7j4lyfJaVJK/Fvpfta2C6YgdPqUtFosofk0+iwv6P7
daRHkhZfVKKnXfOTkuXoUXe/v485XCkjXXmPT6fV9rvLzekbVIe5uRZafWZWdrNapcOAzUIgYfD2
PIv/76djHg34KY6CaQ/dhOHDJ6dBicUSUb/NmaecGa+soFH9oPxWjMb+k6vsBRm0j3CxlZeTh9vu
/I+Au3RyF0Qjr4oB1EbVM1yvMVycOu4bXsNpBhS8OlTjZha7ZQmb5LA43ejiUdvA8zLU+h+tlVZq
Ms4VwAjT2CQRgfLacBCADtmqPlpybpcYHHLT/ckCHr7S6Bp4FZnqDBzskRz7FODYJimtvZvv+7Ux
gHF7dxXiI0gv3IxcfJx7f2BDLsoJIF/NY5rWI3+Bv5iueyblkn0qYzlLM7g2upQoXf75TdeyvL9C
cSqbKOMonmqDjCxfY3Ab3bCzYCGFLISG5Qy8nK0reGHvtjdJKUf8b8PgPMnXHx2sfbq82GutZglY
mieFYGG6jLIkr44KvQMWlK8mowW1mDjIB6rvd/PK3vyJh+SsZZMkWi6ah8Le8GMSlFzkIcCyL3va
6/7PYWIE02LHYZUmdyyEiVBtVrY4W+XlG+b7LhmDUfh0/yAn52g+jQSxgRWej++ZN0HZnvSScnA/
1tmP97t6hKoa/6e0cacMM2OdMy9jyFi7o6VXVPPEbjhQ6dMiirgRwgolpaM/bWNGUFyFoxCeHxre
00lPsEp/vbGMbKS2NKhtjdrcYAY+WgAy7BeFGIkXSuNpe9NGGcWBhTgliHrSwZqo25Rg8DCD8Ybw
4V4CIGsz11/ws/wlEQw1UYIo6CcxO1GZYYhwo5GRwsi4T+XJA+8+69faUPSDR0hCMySSjY8NQqGO
76rPAAAgOwYPFoZWOjRDhr0yMyyrUHrpZrIhqgnv92r3Gn4Sz95AApHbEyBmDmV2OpTsLEAR0x2d
AzSSb+6nbDtLUxaijK4JxZ87W5ECog2bhEXtns4BA7FNz+HCacsx8STs9LIp6Ll2AbHC/Uo6Fq9i
mH17pL/uXXV+fnNbioXAMbaLk0PmK+xN3fNeTdJtatU4gESVSKXeBkcOCERFbIiiCgj2VuUojeih
hu5XcCmzXSNr2fq1I2rFBPo9obmRyRCMVwPy5RQiUH66unKkls4wlxq7NMzUZIBynhHwjoyIY31T
dGbeig1jRtpsItxaoVjsf7KSxuCqU3DHopEWCrkkgE+FZATH3NDF6Ywde+Z01lrYvxCAd2xaxGp9
c0KbmCp2ZooEEvMyVC3skQracI1jw3LqeEc6cROETVAP3Jzb2AoSGoy9jrM2RE5MyJ3iq096tmGO
cqAQJ5R5QAjZRtHyp2XbRnvFclOHl9B6EqfiVyGR5NrFsQml5hA0ecfzGRdhhq8jSkUMQoszvkbN
R4NIdV77fnZI1k1CdFs/spbpXXL4g6eoQeyEhZBZ1LuVzANfAJ53Qw0JWYiLQZHZzr8w31p4tyXq
AL5s4Tl5vsM7w1G95H7m83ClD7Q+6zhfWMSKg06bUz192onMrFahefULvegR1/UOcnLtauWMYZbp
m50zU9c9Z4E1Au6hw8ku+UuLPkrgQNxIDwVQ8pTlOthV+WRlFlPvI51S+377qaHlKoSanN78vntP
LunkAtO9tXEt+uMDuHDi2YKX3JjHZttElVFFCOtqXaSBoE3C0AhCxt3ib5cpKJ/F0bHgC9Sbjj7a
Ve6yZ3lsl7oa2AXQJT7dUASW7fSglwL2xH275/yBmtZXrknHsXo+1tIhRhHm3TE049BSsfkI0HLQ
1ZAHIKzOObu2ptYEYqWtn22fFi0fRK9Nk+2y9mBep1OdiH+UkyM3cDyZ3MmwjLi46IMH2/nOFek3
/pjt/rroTI2tTn++UgC2GhpuFf2b5c1durK3xHIRxDnVjWrsHiyWZ6NKYju+rxu/Bmsx7Xu6Vug9
za/2AhScUo7FYHkvJBPIxYxb5krfADZOi0Leynl9ER96g3FJdt65BK3rWXVLOHOMQNqhwNwr6Rrg
/lO1lm499Kb85Ju79kF7eDR8ec8NBboMMLZDqTLvncKOSbSsZ1h+BxNwbVL6tsrUNJ05V0k3mFE5
jRJXHeSKTn/Eua6fIhWT3HmCPNfeTbcDyYrVLCX2/eUgx6oNSytOM/gb8xHjgbOtwb7nCYo0GbVe
ezjxknGFJ110OQBmAX9VRzm9EGEIHaKk0S3hai1AYl/pyzCIP9ViUKufiBv7laaZGjxQHQWtUzRL
uMW/MkoGJ6rKtjppr7dNHxXiJDyq5rBhSwvGLmmPyAmKGhlPw+PSMRJB3Re4e7RPwD/+jQXG4DOp
AfAwY+3ffu76Jqv+S0QTlR8+LRT4NTlL+ARFNBeC7Xn1THJWcPvtDFP2BIACiZqndhBRqIgF1ILl
c5Nzw+b6JZ4FMMmmn3oq72PQfHB4/UbPrlS5Bld2nHNXWOG4CRyx9uqvpWz7C8q0G1SfJ//HPcq+
LgNGYAF4u7AZ0BEwBdfTVx9Nx5pBQHLbJ2lilc+k8c67uiWZ1OVMAQSFpbWcI8mAbPCFROX8J9jI
2hKpbC8s8uameaXA5OKatKqxs3HU9wR45dhLa/nx/UJn/pl0k8CMO3xe8tZhf3+OlfXOnNm9nYrs
L76Rebo20wvktGbauqTuqnjepPeg10zr0vqWKwr4aU5bWk6/xUkix2zxJxwv58jB4TyvmJ/QJUWZ
MGXGBESXLT2qAFt4EmLGanH8qmPDXZ4cnOQ52VyUXUe4QGqGr0LQd/K1mWFdSKyFFb/kCwbGhWE6
TN84CFUDFdHG2OAB+JGhnXvbQzVXwFM/7ikqNCe1YgYxs7UCm4lqns2cZKRlMPN9QJuNLuZ1EqTl
KM+KBe61FYagSppzwsBjgtVAG/kjZ3KMumUJVj9A3gMEfNZMHWc2SY2v7vjlLNMp/hX+CPCmCREx
FW12HUJ16qb9eZLFXK8IE7qdkTQq0q5Zl2HN630UMHZzjLHvrsO3IZmYqDrNpr56mvSX38gcwvBr
SsbLcL9f9E8LyipHAfVxPM6kkIA6MZd9twhWnrpONkyMMUwVirQOj2R6mO8wmhfnZh2M79YqPcJK
YsLEdfVOFhaZu/hjefMqsuoOJ+Xtc99clD6oSu59untrg6OsyjQ3wUN6lXDayODIQRBveuyP2Ua4
pEtI2ba5iGz7gXblJcpoWgd0QiJzLLC9ZelcN3RTnF8l0/U63WfNtYoTE6SL6jZn8t8pxna54o10
tDgNXdPoerOxxFvNpu61PdRjQH+8iGjyERyxQ0xMrE0/at/KtaDS20dzAAwtUcvzwY19YFIbOVLk
qOdX2IKmS2rmekYdm7p7wWQt4ZlEqp7l6mCwYSGYNgezXCrPZtkIKlzNxTTZpnkWaFFfX5e6fXnU
NkmNvPA2d9fhKA9dsL1Tz7BKbvvZqIe95S6N6tg5fO76F1rsId9cVLegY7zGQ7gZwFP5DBDRrqJ2
utoFI79zE879lkSMKA1Xa5MBNT8Xi2xe6hdbOtZpjgmL1DacE6giHY7CtN8X2yfns6iaIeEKWm0o
aRFnSoGCpnUdWRp2N54HvKyHK9d2bbWXMIjuppV922kj7fR72y01wJ92JhNVDdvCs3Z9p/EkBtVL
60XEBccsHaz797Uxs5MTtKkioaiRmuDWJ8hyXvDO/liMAPuQ5hs7hhPMQgugkNPqRnn8XAOGQ68Y
m/iSThqebDsjx8C5cq5YS3OQ7ybH0scRhND4ZV7mipfsmtHOFvCtlUKYnwUBgowmigbPybW/e5Er
oH0mfhxMo7tRJjkhe/xL89Mam/ewHQlZ1KUzqhFP6GXB/9mkYlrEohdQGLbXF5m/AyEsBIGbow41
VPLMAtHqnLW3PXoEgFdQBUkTjl5zdRJ7FqlFu+bfIWGNdZBeHXPHCOhsQC9YPdhva0bRyG3vxPM2
p4ha4vc/Sns2cHZGvBu5z3gEvo0DBuP7vzlRc1F+fYmOpgm+p+zotYAX7IZOWe67SGoXCCM9zb+5
o/5oH++cXpOal1Gqh7AfvMOIb/Rl1/kqqackFwzreblutWLm83WdZK2crcD+c+CNsi3+cymWlNCK
iE3/9kW2FZTGHZiaaldBYPHCCakczGYQPfsDxySLmNnbZV0dXw4UgIg2+tc5h/jgJFCKJ/LP5QWo
JQFmdLTlnvh9yAOl9benSoSV0zYKBNyz4QZ/SdLM83vIDaeQSLOWrfNuzzeXdEjpP8YjVIzYhDKJ
UOGQSsZvCSwIUc9SamvAklHTp26GsOnw6SFgch9q6SI7eV702nta7lYqZidCf3yR+oKtqrTukMNY
w7BdYa76GLnd+vKTkmvp/lNIC2RHqGfFcXAPCkIS0fzPQEs5x1NuOOYIxiPi0vsfNXaJltP0iAEr
1dPRASrzOOROa/8ON9sY+RpNJoC15kme5DKnN+IZHNlVar/qFRdIAgHJEyDyz9p6Vd4u+C/qXis2
8k/efXaM0f1y/XRxWcud5Ge9KutnTy99/L7bZFi04vHJhtQirlOFnBiPaPxDnXF3eXkNrXkJ06sP
xVfJX8SZUBSMGoMS6K/sDmmCiAs4tOWkbHfu0W53cXxRxQBG27JIhkY0dG2L6ErcIJ6wZSpIMfo7
fr15/sUTM4CpKbTd8ThMODbunB8xRuiahXY7vB2GhPZxi7IOa2Z8e0uD/TCW+lk8ja6dhz7vt/p7
kEP68HlfNqvWKSwJ5S3snAIGhT+2L19Rhu7Ay1jG+KNBNlap+MHnrTokp5yJpWZfctBtQYWBLGa5
Kd6V8oltw2RSCssEqHH0qK6v8FR9QqgM2Plug7gVlXkoZrwMkLAoG73Iq/ceqZcc6gyXjKne+WBe
XpxR+/Ar4iWj8NepKL4e+u27yHt1xfNlRnJeOnXuGbWqiabzK+DSLLAlGZ+yLcHxOZ7tUBZ5Z831
N37uhc8GbHtalNGUNs6TMtrXlvCqRftYSCaacTr4wnIefgNYPU9OC5irWNcmKveYKAT7MI6lOr/O
ww0bjvlF581Rrr2ETaXyTrkdv9GhwBvO5dPwS0EK/hKjZ4gxAEipUtqY3UCF6YpyRFPUGZsNIQeb
445kF3523iqoR9hDXCPjbhNTvxCeZWZCU439mm5RIh7PJRL+mzyyoI44ixJLJgBae9uKekAzYmvf
cQbcCZfsKZKTE4fEkw75Hr4kYBTnJJ8U2MEScWGKGeDXuVDfY9Pdn2BqG3ZAt/qMVTrZelEC1Lq+
yvVKnd1eGXrtLI/2XLA4FcIXKh/Tkk5E5Vyn9Zs8CeyhXy7CUzEN0/kLPJPMnwmLnQ5oATjE03Ms
tmOHc0t48Dso+/RbfZoioXfbSzgZPkrFDP2QzP7l9OCMwMF+pk3tw729L3C54ptMLUv3lA1WwbFX
WsJM63F2wJ26N3Enw4Y4r1xIWlhEknymSJ24dNMooYwt90DmG3aj2ML93K3o7B02uXgdJCKQewEf
R6r7uUaPHp1XTcLnrOqP3yUmvZySSBZlIk4nrVkWEQw15xNlKeXsSFm4SNXLNloNHWJqU5iFt6aX
mH09ipxIicygjj36f0M9InFk0OCh2xkiXGAa/OOSHZLbFMp/HiBSUyUAEhous/x7u8QalwKEJChS
DMoUb0beDuUeqWabVXSEfSNhcQwAF8rqLXQVoSUgsatNfS5GFn+pjz8/wATyN+/7Lif9hWCdpzXf
Qe9WDfB4lmNDncIFMMAgL/W9al2AMFkDi97yadnDhi4MNU8yZ+BUf3TC6c+Rxl8RzhPKW6gj6tXO
GQgn3QDEt7MrZbHg1XLbnbrT74lRpWYx4cHjVX2pUaGYyP8PwYJXah787q7HYp4eT758vwkfVT/W
UDLJAa4l/EOOKGYg7vn+/VJiexv9LZWq8Squiianw1xA8IzBAj8H2z8z4tMp8GmwV8CH1D/a00KF
r9goMVxZxNcZRow3tjdQ6DYCXSOBFo2FEirBDah/aZ3fv4rUqe6i9moJqT9owQ5GnKAsJMF5HCAm
iFZmFezec9aCAKQWP4P7PSDtBPDFRcbzAxTzUtxWTpYXOIcewjtBPP0DV16STN1JARIZD5f1Uv4C
aos2vkoVRzHmAMebYuQezWfPEVz07PkjLtVLmmPRiM5oyLbT4RN7EoHTO7GJ5pQUAumNZjksFG8w
YAs/rLsgn/a27YTVtWgqImSOvpRbGsXRt+/wSCnujCdr7FuCvpSO6MzVH+Va2/p3ZjggLoMRMOh7
hNrzJ4jd4MYDHF1BgKt6ZCDBKvD5v1IA08IHGxDqWkU7LKCXE7NlWrpNPu5PsKxv0wjE7zXDC4X1
EC+cCZPVWKnJ1Do6l4nyyvah8FxDHsvlY3lABDjgWm71mwpz9U1AU8UIETXstnw3juHVcAwplGP6
wYrH0zm9mwkAGXMQT9nhV+0yzDdAiyKVjF/4rnmWKUKYojDGjrbRI/jzs0LT+GvzAoh7YBOYF8bw
XMdTTIS3mnUjqYUjb3lpTV2C4UNgscsHNPa0jeER4gcvvfE5Q7Ezvk/r835pf4uXaTh3YT0ldGi0
ry8WJRa1RLPqGGDVDRGTECaB0qU8LvjozMVOiMFPNvq2Y1S/1W0zceU4QeEiyVFXlix6N+oaZ2Zf
vA2f/7QLmKDkpGMM0DH+JWm9xxgh+aoCijdKugSt5iuiluKx24UNTN557GsExsVIcyJGNu8RTrXm
Rl6RkdprkeneFXI/fvgJF/PrcFsFpfpvmKg5gfQAPhbqkPG4+k2F0nUmTN/oYtA2TV74dosSpplp
ZjjsjgiGoYqi3kcnjQQ9gvFblYo4pbIKAur6DbW+97GtiAnd3EKes/0jZYD4Y/+MM4Z3IsBPg4Vq
A7ZRJHYM5b7C5NniL5XKuJpdf1Oi/ShOjVj0iPe1ZSjdiY+769AFNP7fM9zYdTekabVnJNpQzxGN
EDLWn0rDn35lcfjAAyakvYU1wKk5tjaGjV9g0O44o/gK+gRVT7mP5JywnlpRxl4Mxa2jQT/5MHDQ
BmE/jxsOq0pMtJiejex2TsQDOsiFTKrT5ue1vBjNReweMVYe+VLkLoxCMOTa+PB7XiW3Lfea7HZ7
HUKN0wqHK340Hp8d3VXiQ6E9Su45W+RK2Yx0izDA3orbIMiHxPhJQsc2vmrPRTE5fGSMHAIRSmlU
aaAXf0QW8CJ8fxGeZJUlLqQyraYHQj1AyaVCpjBUV1gzdx9C14oAR0sZ9pcJpVivaElGwTOjal+I
mEbuVW/oP2Y4nsX/HmysSymJVCSGkexk0DSDNLyW/g916wCRTbIMeQo+NDDbnVN7bRGITOhhTSbi
V+9QmrQukDpp3weMNgP4MZ5Uv6xxipcG0bZScj8VAhT0/6OFIj/npN+2iJnt1H26HWeTC3gbC7Tj
J16P/PyNjfGErR51xMoOVukgDMPCoQ4t6RLzl94dh5VU/lxFKmvObmxV5FSY/l3vXpI3dq6qrcwG
NO0N61IdxtaVLvNIxw7Pvik1LAQs0Pr6tIXqXWNxhSYDw6KYhdLNmkA/dNSokbiZ0fuWE43+hMzz
jlGGY2MPq+4Z5+uHpkp1Vo/jKi0ctzIkhusAoqBdka8m13WR0cdw36ahDt6oakApEGIRLtxEryQD
q5M11IqlotrHeDs3cPQ80W9MnIa1BYgTAWjMJMC2QX6DeGv2Zp03xBA3U/1uqIOhkEnX+V1wbrgz
Tdno28Ahr1Lq+AzDxlhPq6eCOmkRXUrOMvIB4kayJAzKE/g3bqTuA4pA5EltVT9eUMdhFLAfyI/r
k9v0aicTSXK2mprTXOVaqg3zcr/ZMgRlXgqTPVTphhl5J28ybFwjwjV+8cpI3GKCfZZvcJUqUXbU
zupM/lgGHHjPKA1MhHcz+8ciH3QLBsGnvjwBzTBKQuJhK9L7ACFMyez41NCCkiTWABHKzYdtuYix
XHnaCw1NLpSQY0LYGHfe5M69r6YLNVPyDEIDtLPWoqKrg/LsKV+UhrkRYlY4Kpndc6UPCvEZVOM1
Dy9MEZT+MYncdV0+IyOH9D07WzAaOrLDbUu9KsCIVC+/bjJnf0ovyE6GJg7ADnuM+FBO5J4/rgfR
c5Pi+0xQOcH5DM2GRRqA5B8BINwoT8g2FZYxCZldcbI8FcNvT+8FHkLj3hv8Jg5WjGuwmo0y6clo
UUTdg/wSin+ZAgljPlPo2QzvH0vp1jf0wNZQ+ESmUAhlLqPFi2c5y7sFAKFKWNBgHQ623fl8cFts
hX1ungKheF3IuX5VcKErk3n24g1nEEn43+7z3nNhjYVph6///JiSqFac5DDUFXZ+MivZJE/znWse
rhs3yf/zZ9/nne2VtYZOPeq+qfTrUG7ba0YPcatVn8ll+eDiMNUVfEp3Jp//vdk81132NRuDk7fg
inDytS7K1BlR989t4/JPaq1EcA6RRyniHxmxGZRTBlSZnmxDJqnNmnkGS2KsTnf6MF3N7mNWrj41
KbNtqnl8CI+RifjIev29NfPTObcHcgwNwuidfjiNYPJ2CKqYLcb42nw9wSOELlT6RaKz2ZPK15Sa
2YFTJysU1eoL+NE5cOcrXmnbIk6WP1pOykHYi/vPFv3MTIjOOrY4jjrqqIIg7kyVoT/Kiw3tKQH8
iJvT6O05IjlbqepEtMA8PPCgxGzqJjDOgqNoVhJZB7aYh0yV7U2u2LYvYgq7MpOWxeB7fwXIOHq5
tMtobqB7nr3HuA+nbZI0Mk3bXh2xghzrSXJJX3hM96b8vRlDKLGyBSp8xmDbkeAEp6DcAt5sa0lH
hWAmLut36b5ChHJOlIH339nQ4tMQA8nesVSQy5EeB5FLbMLpcs8+vXT9dVItFuMr0tvJLKFZwAGe
Q0iWl1iRUota4dEgW13qO3yvWPNmC3zg8NLxwq0eYl4Pele9dKO7gCdvs+JRbeqAYze9WjiQQC8q
pK9Hj8Qq14QB7I1CCRdsqj8Jd+EFN1yaKplee5XTmBjs7hlEy8gIEv3XuoZ8aUQ0aBkwreHvHuin
mxacwHa16h8RgjI3gg6rk5BdZLIkQJC0c6Qzg3CuhSp9xwFGVY4iOnlwpIdzFuzP5tzZi7qZwB/4
fCBd7i52YU4oaZkPmJeW2/nrDXXiKX0iBUD/7PXBPc6Sqn05oNABqcB6atUH/IlyP1I5V11p3CRE
DuHRjxs2F4PmImmokREp7X9vyWsLrRHvHK7njWY6Gjskf5FDnB8sijgdzxuba4Z47ABGFpmOsbzg
It6HNr3xfljMUW1l0QknYIRkShjxBlK7bCeXr5RN9Vcpfrdt619MYBe7RTFc8VuEeEO5K+AHnZF4
WdTNp0qMUodDJPUd7v/5q7Wpdzlm1YOSwAiX45OaL+sK0KN1n/wBHIYBz91PKMOJM546ZM5rvI/H
MZFYQCBqJRYYJidlEJMqGFzw6VFapn63PksEhIGZlVYd5qRsfdV+C7hsvxwhv0hmiPf+gIwaqT2h
PhpT4lVI8106v4E9gfzPoJ9CpHZj7FrjaN1skjHf5JXecdcMEccX9MpE734ImKWvkpTfDGIyRKkD
3lKJz6reG0QQ4pll3gnj4JJ+eox62YkHn7g4wIfAACJ7ZdTAoTad7zPWxLatN2IBmcxldEYIR5P7
+K2zkceJZwzM1TK25DxvXrEzIU+hcawzc1sWg+h6oAUscf/ARhgzNCj2I1CUtcY/peQkyAqVVAaG
sKOpEApIbW+E+wxPW8sF+ajkruXC6Z4Ke4iPAKhqdinrRA+RmPWaMURvS0j3o1FOn5d1ay8aW9JE
rB9md6c/x/wgpvzOAy49qmbDgd9697YXnTcu/jzD3u9OuVqMCduBvCJgk5ApoGB3PebSH5fZIqIq
rMR+GN1RaDnYu1qzgcudTlMvb+HuqVOKwsNi2GGPsNGw7Q2/4bkzEy2TVOpBpI65dTYvHhyzR/l/
WNVa8bbP9ETn0Zgj+3rzoXCYbCsTLatSTKVQVEWm66ZW+y4j9SoeC2IUOfGCpznYsCUj9uGJ7w1K
GFGv2oeTNFfpFtA396W/usKb8bQ8mEQgC3COgYEZhDdO6SLt3U0aZYHYUiH2WTX+a5I2jurwv61W
IJ+ckwjS2jIroNQfL5SRZ0tlDXIENlGL65a/nfOonOj8N1VNCoKllrn14C753F7u6lFKehpoDJK3
My19CA/tRSND4zIBOtv4E4e4zLOa+1tTJ69T8z5pLFnKrKIO1/LvY78LH2oLcwmKGSihdIU0JMaw
OCB63YkG0yLhs2AcKbhr0bnUpeEjRxfJ/PVeh+pzPnQ0JBdzFwBQeVMx2dc7kZTrN/9VBiSWLXDX
VaSNaQSkLGhmsiL6SjXELyCY6y3vyVWYZm4qtIxxIUOUvdkErmbUJGmujMI2t1RrAmXr5UxyMuaC
0G58ZyeTYudlfL4xb2Xvra3fs5c15BmYTUvQLqjQ2lT2DxteycoAd4RJ9YlfOC6Bqoz0RWB0yqMR
oYJv9eMrrqm82bDi+/NC2HZLBa1luzvMlesDc+tkE7SuhLl0z71H3yAZPYBDHKKvNBHUev8w5Y2A
m4Ws+dyElaQqLESQAD4rdNx2813IDZPoXSnpDJRRVswIu5eShM3SuTWIUj+VwTFerCXmZmvJRJ+d
IR0kHu0bZdEnfwZONKzZfQ/4QyO6fXVoeodiydCnaprZlfT7TVbEhaaz8WuyO/0z+lZbAGhhxw5N
VN6DL2lo5I/FWaOczFa77u6l92NZfpgGlxYGk70stOQS15m4XuK+gtwUCOKCK1+CtTW6358HIUvM
gb6FXWiEAjVRXjYU/kiAYH1ROwy4OFtLj/eGDdII3F+7YIjcGaJ+/XMXsb29QS1anmF30NWw1rJh
557I/00j0NuKy89Vr3tAkPXC6WBuX2iHvk5i1YDlIw7YfrjHHA2qcCAVDaBq1sKLG4rJm5QO75p9
fRq3WzO5tbBI2bB/iZVvrFbYe59iXj8OlIoGbyE4VwIePsmrbJJjZMZbDA1iyzMhWME8KbQTWjOc
OvcT8/jIFS5Qzd8l3eldUsOZKbxPpk/bbImgzRiTTE4mE99Anx+z1rSfioL+NpXfyH2zS3yXkbr1
E2oM+DFmFBqGTsTAE5M33fCIqKt6SOPz5yuEGkkaRgyngbQlPQa4r/GDuCPyiYzKkOv5jiDvV55g
GgwdJizEsZulWdyX3THu2OLc/QAYgFr1dGr1pURqoSUpw6O9KaQZwn1N17SSzWpZr5ZFhtAdeiLl
4sj/qp08wC3a4HgllRO3NIB/Y7kA46PrYiyB2BFQTFOYt9Si5/oCl0GC2v/FVZ4k2UQA9rFc6wQu
ZKy/Ukxq0Lr2QX2uoHBMKAR4RX1bAfscSX18LHg0C9hP603FewqTSkfm3kbc6co0p63aVS72DKpC
lu62teMz7IwTX41wVapVdIm/2wFlbtlkrrqVykASRQDEAamqsxC7OdufBFbDcaEWZhh4ym/0cKo7
y3FUGeG2y7XhCyBmESEjQxFhHkkvivfrgVk/WPVk64iu6Y1jcBam0rI5o+Zd/OqKtXXLRrIQZjpT
4/WatfaAqWTxo9HxZGS7ZamQBUCIdpTdg/X2J2NV29Eiu0yQM6HYRQSFE8RzV0rcKIGgiUop/XT7
cuHX+f6UvQxPScpGg5hfyFiI4Us7nFSTk9ssErSGxr6uRZFOkUwaAORvaD/EWQUUHm8sZyYmTd+8
SJqd36N4ScrIsLPTOVuY5y+mt7ITKrzDKgCaeYRduXj8ZxbBzCMgaa2xm9wVmKOAd0rt0zmPLvUB
GdS5aWGPWxlJbWslxAF9jP2wAX79jkVheMP25/o3befZBPsIhZbr+BsRANa9czX/sge06sWYMi3R
q6tAahzfGmyduPUCC5l1/0CZf2T2s5AZETwoZH6t7Mo8KvMHK16+NrjaU7wllWOGVLDzm4PRpTcC
+djONjwu1MZrC4buBPYurAuFNMu5V6WxVUG3a5D70EDUy+zFES6JcCgYsKNh8JHHJdntYMzN3YXS
0cqVw0lHzqo5Xi096oob6PLcXks2mdVJ9mUjyght1VFlN7H3JFB92hFidHCtGspbcNSsWYmUBCXC
3Q22igLB7NBZefh/VOLodvHfiig5cEHqmG1wCwRthZmoqA/17UyvR0pBkZ7tQSVdCjMMVeIbQa9S
4PvxrVXBU8jeu/mBxyZlI0wdHMFRR8ggRWOzfKxm9tuTMjTqS+V9CoPc1mTnv9HBi8UxwQMMJyP2
lB2LlPcT1Tk2vXbzGcsj2EZCSx2pitIUv8w0ahL1q9Ms9jNxucfAdmDaMpdYYQPJgZO1RWwEL75z
bBUYNO0+XaM43cDRETVClDJlJN9Ojh7BPptuSbvRNQijRMrHUD3pGazH9+KEGj6ZWjYlTyhcr+L2
fS/Tkf1X6f3yeW5fTD4rFfjQtNa6tzZ/QJsXId+3NPX6qPsXOagtwkGujFF3BMj0gVcg4gU9GOD3
0MBxqL3KLOK9bK7pUqw2lrvZSFfaxrqSi1bciePHuzrfQgW/QoF4LvdrwcbQLU2deNQ7zVey+IBm
StUuH7FlSx5LgYgx87syKuAdhrICyXLHslyTqMdUqG6xe/DWuhwZWVPLFmzrhL6FMvOmu5LxYJYR
05E8IFyHcRwREMuv3k83GDL1pmY5HdTqc/wLqYt+grXXyi3A3TzrAZWJjx6Me+JJBSWnYNToZGM4
0qHm3/lowvAIMSB1m5me5qG3XC0lhjrq7TnU/UpFVZdvlV72E+s5lbkAnIbToLWBpiUpEl1nWCue
zY8Ve5V6JEdTgKLnGV42JD3GN3KfM4l4fWtkZKpUj0mmQeYqFuzIJlHQDD4kXbp7J73h5w/EFlqo
bf59gTDWhmQ8yh8pfzsa+OaAuAqltjBFG3+Vy9uSMRewa/jKuaOD8UcdZgPW3LlkLwayXiCe0MX3
EOZu7g+yyQ82qa4NO9WNqTLRgQgn0mW9v4qrTn2/ZMzL20fkGLWy0qM9DltBF20tem7NRP3HEauX
CsfNyZbCs8MGx8wP67DyAVVNlPgx+ymEbeVbuSmwvNUP1cl8ts8pyw7RGuqcv6/D2BNt9uwV+CWM
SaaR1H6qUfNV0vT6C58Yb7/YT6mUIO4s1md5IBKf0iKPAdGOksKh0D29ZQL/1aafSyv4d6ZPdMSk
jqOtjH25fipE1I2IWmGylbmJGuVIJKwMMt5WnJDHfw9nzJQl4Mf5dITYScFv6agzWk0uxZx5MbB/
aIey2L0pvzU1sYMiQIgCdvsHCWKO4bzS3v1tTGeZV2yruIz/+f8msanSgfT684ppqX+mb8saa02s
XPNJJIZ0ivHlibkoniYdxdLXNq7mt7pZrtXNLYR64J9rA+WmW8Zwv5lCCVQYqo9fkNb6PjtmknQD
cqreXgMKsVwAINUqCqzu5K/0l9v6nzod9IjgoVTIHB+TAM0Xyl5yvOxbtn8RayBX3ox75YY2VxbC
aaZIU8VwzJpLnMnT42RFmVXB6DMYd8M8yVFYln52P8IoTBqcfkxiLXlbcNDKBtb4Jt99i7CBl+4D
bThHxjlIuq35IuYTw2qCYpRqTYd/pzfLH7VtNmSg8qXA0bj+Xx00977GC4AKCNPCLC0aVVvsEy5A
Cd4sckzytWikW4yqfr1jcXyYjmoJP3NvhNYdl6nfcSgvg6SLXMIVYv/nEoyPs8GlgYtPaKRnhQg4
X94HCKPzH1d4jy1fm/un1YAy16ymAuPLKdM6oUn8xoSSrnptdhmg0QfpXYKpVa68uBlTUXicQH+p
KR8TBOw5A9Po4nYFwrf2Y7DbG5AtMgXl0ETHLFlG2Dh/7n3Xj5S1e7Fmb5R2dzkF9W2cFDDp+0pS
Oza88aRmOnYgMQ3TNRf+HEo8rjfIDTPyjwPMrCb5ugI9ye055cix+TzSR4KuCALI5E/OE1rsT+wh
+8FED9pZ4sOc56Xl1SMsIklCzgGXAD7EMApTf6381ozqydytT+x8+H8xxksknNcT5J4pkfaUoI5b
OtFFecYnke6KxumR/TwO3+wuEIc4XPP2buxEcN/CPa+JTwRvIwgH49D2yvoN/gsvcViZY8AG3iJj
HjKrqIzBgooMcjn7HYpUYp/K5yPrB6bAOSuwdOCZqHWw57i/OKjwNQg0P4NelPR/MmX7iwqQ12ta
KFPtuPfn5/Ja1EphsxdJSPl4wCcZRpQLGPSs+UjV7FkpUHX65q5A456Mo+l8uNj8qtc5SmAOYDlv
padOzqa4wL+9akYoaxlxcn+ykfzQh+tnPuvEhmpHykedilrbWk6ke5erK5cp63p5WhOfAXhahD3M
RRIyge+oPqEGA1LN8vc6vDExr3+NOgLZtjRuAuQtoe9bvcJHmIZIAklfLnimkqE5r69REe+9MrMz
r0nv2bx2szUrfnn3uncrypI2sc+QrjkD43LWtwpKtjnGPQ3e6aL8qZBn98kYmZb0hS4xO7Zzf0td
iX6WkL2iGMlk0qdTj4vmold2jgtkeOyeYRqRsb116w3AvbDV8JaFYILJLhp5e9KzsTS/iVDGIAtz
h1Caq8eQUMAxvhneFiw292Me/pmvwghnaI3BzgBMduMpGI+PK7bGNTKjVs6t/kb6rdG1/bRXaams
6fg6fZEs69HMQcM69AdYQnENCLG6OosIkbq/WQgbf7TD3bIK+hAcfq5EIL/hjhdR082zF3h77Wr+
JhmkmsnjLHI6dkSLpKOwk/+nmkTANFAHTofHGUJAEE1dL/aV/ZVaKjPl7wNFik+JCx2lIR8tBJA/
ELSXinN+rexKB9OFZ1Xrqw9RkWf+tt+9yKxp+VFgC933mVwS6jzzbMyt/uQpEIkeGdwIIAld7Xa7
uu00N4TnhCZ9gfbwxVr+J6gRdYISSyd5YNPqDtVDzolqAsZhAujln9FrJPrDf1AENZJRsxlYqCl9
NhAqAhXj5Kt8Lyd6d2qjnhUNx0bPP5h0LqlLYallLiiszygO8Tl/T2zX+20v5MD4bl1r0ew9uvKv
MKrMdLGjlrcWcf1VBYo6Sv1MkV/JlKlVVfdCFtyJyUAKjNP9iqd9/wSwow3vuD9NxSnfQFi1RZ3b
RNNtzNFbKiaO6/YGT0Hlvc5cs5reth7aIc3TxdywlobQmmYv1m2wjJ4llB9DJRlyft0TuLnNBWLA
8HM0SZt0TNl+3tCL+cxhsZfq3V1Dv4hH6NnUwb2+yCD8Ifnm8p8TelNaYj2w66IWQLwn3JQKqw5f
65oiV/Ho4Z/3ExcoCMNAtyDWPhnQi+aiGus2UxE94xg8DJg2Wc3h3bFyjX90yD32RvxEecTPu4R9
1zH8yQyNBS2AB8HAeHDJ0+jEIna3EjyuBG2Yt2gA+b4fQV5q2hQoHsYT0vOF7RZ8e1tt+wU1wDic
mUn6z3FwDWR6C+WNQtIf2d8G3zYvF/hcaon+KrdiG1CR5b9/dMUzvmoDT0vAQbGosKGvv/VvdgNE
db+8Ihtcd7ggcFH7TlwJlFzVcrk+xd8epNwiTiF8hG0HTaGtHJ1RN/LYUWvZmWmZ6tZv8wIErZNA
bdMZHrP878q1yzmZcMB1wA7fyvMk94rgQpscpG7oQD+RAV35ohuFFzCR4worQGRk/e2ta/RNeYMb
o41hbOIMeF1p5JEOY6hICRv9LZMkSfk7yqCfwC/oSvdqwFhdLKFhiLnG+bTt9cI3LtM778MP7xcP
QDB7SCQueYWM44wBUaoECfkGc9oflUIsd4thuajpEq/Jdg2+NkUyCTxRE07m6YYLps1GjeVom02Z
y477YifGTjoAQBwmGSY5cJxBubihUFZUe/WWFPszyGUqbEP47rpVDvK/BlPtG7fGLTsggELRM5cq
hDdogt1xJqtlFW353H4spAKg/5/ledUv46TRMuRbIokvyD+cUGERub6aWXkPN7vghkskM8HPus+Q
TpoHO18NolSRTPuU6MPJZAqwv2ahrfIp9fBp0CFlwY0/qb7OVlklG6sVRCFQhA95+BMDMzSbhMtE
mFVTU7EK/SBYxmlKndOydGOqvbWgu8RJi5WVnpWkgyJ3gavhgZkveu0mSfbrOVs42dclXi6I1JsG
igljua0IhKlOv8htDYLBaQyysUIFo8E2O27DqOA+VHHnZ99/CPQupVUBJ2qdU0lehxptlwi8EjVa
wtqH69d+l+frtcOvYarh2WrwNQ9ExcJUN9U+2iO9kn9cp/7RxaYLLqI5OrEfQi/sFBkDP8qysl3k
zIXPZjys2/DkcPJQElX/ndRFIgCUXHybbF83L4UJFdCQVSs5zaMgjYjM/FTTDSK9uHfwEMyGUvd/
7TFzoR5GGnkZf4SpMtogoqg8ALimgOqIrxOGodljsACD8Zjyjwbwg3oiS1eUeyfz4qJi31Ahfeu9
PMWhTj1XLTMVtxxDvg3UyvUyO93EhvHGj0UVqE1t1+4qNRTRl9mR6rhnvwRA8Gn8bctDtrM9c/oc
KgWZQuZ9M2X8MCrGcrtA8r59aGtd6rn9TMUOZRanuN9ywetkO1sDHKFIqUg/ITGY9AaddyqxIutM
cnrOYwY8kSeoE12hoexQHhEcwfahrPWRWm5oBrUXtD9Z9M80Ll9REVVWC0OkOVR61rpNc1FIPbK1
4roguc40eHBwiSy1/g/atvITa0TBks4vHzswXI6kLsIIkI6EO/kXhYo5M07pd5l4eDtpy5ek05LL
a8D/qcj7OK9/P2ftgYP3boejta2YN88fHKc9SVgH4j2lDWX3iUbcDlYUPOfu9OhDlQTOmXPyoWI+
FjFTz0NTFSmGfPw+65gWLKKVtL7iIASseowS00Yw8nT/8azEjBC6BBLTmdqCU7tjZbbPgMbNVzhs
76Jjin1XBH1I1DSq7Wd41hrO93NWpKZw5o9iE8EJJDcGiYVqOrAfUJpQXJY5BTR6y+aOobcl/msz
FteF5nu8AIvn4SBrVSwz0BZY324PFDCrBdzdyzjtOqEKhlPIpdZn8i4opyPN1EtfBfo825o8s/hu
uRj1jozQyHHHtOod+asnrWXmeuT7OCI2tZl98nY7WYvjdCyiW3eMUiOpxgSg6DD17mQlhjeGTpKc
JJ6apHWXCNRShByinUhFXN/jvcTtGTvYyr0EtxrMo5u0mAGJuTI/f5qSlirgw3Ez6PU42/RXb8h2
rOISILkzOf/ioyxuudjgUp0dwX6cY64h1i0qy4cTte66ottqK7ldExMRrNFjhW0nENJWCKymToFV
eCzXPd77wTJSdFs85OibZKsmEARy7s2d3o0RBgnKsBI4I5MBKWhizgylPw/BnLN1qrPVTeCcI7a0
AeFiuqw87LdnZqwXLjvKUhbBdtDcSnVF2jn6rY5hTiLfILpCdviYBnG8qpFoWk8L2z/CM1k+vI/d
RStjbrN3Khwci4DYJGmJ0KbcZXGb0vdQO/+86c8f+G2m+uQMAHZTJZHJ+perJigJGGr92eXxxWCM
p3TqmX9QA9e4I0xOoLSMreDLnFIHKdMOx+8/Hgj8aP+5ysC97EvIdsSb0mGC7UfZJY+tJoginn1A
qccx/flfB8wqsT1Or+YfsljuaMgfiVbLfkpsGpS7Nxp+STEYUTFueC9kzQ6e5Z1enILkTEJNotNj
eDGHjs74hx56kZAi3NyXMxXRTRldtmIXoS+R1bgQt5q329vPKZK8tP5wzdhxpaIreAmI3K+dMu8e
e9zmLFcR6xY7RdFNlf83yw80ulAx02iHhBIg5VuUrqQGGEbDd8P501aPaKOSavWeO3ZA9X3MUv7a
7EVKIiKFi2Xj4iFhUfA7dNtebPkPZCw+8ULXNvSFjEzzbcjqoqqCawHiKwPQnodVFEbvgOyJorxh
sUzw4O7O8RsmjtVts5RYIVWRb9//ZukR3m/1AS3SiJvoYipnTpfLzwk8YSR/qmqfKoDHTpqhhhOU
NRr56lYbmVnM1Z2yb6eVwOYbh/IRjK5Lr+MuFYYlHygdRKQW03fpqoOTEn/npohXW6N2GQS+n8kP
MX0lbwszrAKnstm+gtRpOYGQL+t/h9Bv8f4nhHuCmq2Ul+D5FaiG5n362/9pBuGDzcWpwISLCM7F
lnOBVJzgoDRCzMwWsgjKuAvNI6EqlejHi9il5RGZ38I3WQ5Q6dGmpvKPPAzV7wg7vx0smTB3HRVz
X0p2efTwKHJESMplPIlmawcXAWcYfyhCFZxdLRAQHbnS4NwD9eOY2CbIPHjtjdPrpSCoQD2Cx85E
teS+CLaIcGgjTgnndzA9oW+ctLe96LFiy8ikre1tBU3fBMe9Bl+l75EVs/luL+v5FfrA4pI/QDEI
29P5+WwXTx8JEWe6lJUPyUfuitwfu1FPgfgF9fUCNGFjAE1HKXlIaVxqRDClqa6BheNuhWuy/kMT
VjWQil8eMe6gl3+vCH508BbXwyIijK43SlXJrpmaDhWyb1fTZNtOqJs7B/BqqwjMTy0Lxvaxjy+3
uPeYKJF51qpNcZ7o4tYZSkWkCeiYWMgiGV1SLrO9vT+votBywNrKjYnRRGq55H07LeRcLYTA+vmo
Kp8fbEtPY0JOQf1w6wdianG0S2h/7uRbeVwCPGdHxufQuAo8mTx6qBjnQCi3RRQaqHngiWkPHG5o
Fl+0kIRv24UhDtpGx0V0RsYN+5LSdWi0QjblVAcFR3Rd/516ainyS0F9FuwporBI588UUn3Iscuc
QGLtkU5ih9S7BgMeP63biQFRxQkxLYiSs6jUdcXRBDTGtr9OvuJdAg0MU4+B8F+cFpNO36UQ2XgN
i41WysNkeP7lGW5Fj908n+oDECsmlte2Hjy+JIrVTfD2a4DqqpQkBGdoiJD7k7o5oqJXl6v5hwVx
EqhWC2sb+UUD9Ryfeh4YZTY55SVw4R+EgSe/cY1KXwrJNfAa7lVYDpFt+8GjyzFQNNMF1ya/YEsS
iXSDoPsWCibI+aYLK8NSdz5mLG9Wv8tWgtuNwygAFpA+8Qd2TqXKBrbHno5xKENSUsl3sD/Q2HKS
6rty2xznqcFCFtjj9RZXDDb+2yP1PYch92nfEpKLc+1ceXWmR706X7UQGZU0xJsrtEXU8cYFp+Ut
RZ+OvqFOserbAQNLFQ6iHDBweg5ZnQg4GSDApSXkrAErmlPiD0Jjaj1GIIdXKHc9pCIIpH5zNkYX
2uZzLHlp+GFFRHLjKy7p6pabjeh5dhIuVVH66JaMsG05VfyTS02HCsv/jmjmw3hTV9dNQcHmF0Hq
yFzaWurkxS6ftXnAb0NW5RC1dDm7YyaSQtX6CVev0dpGSpS0LY/pHgBOPBNeOSPZPsbriBv2koGa
E9lH4FG9Gt87pFEyXzZUWjjJM6+b/z/kWLlHmFLkufEMvP/nobPNVIvDFtADJruke7ETOrw3qUN3
hacVBbsQNSpSNI3pxw0ZlwCy8wNoyMH5p2EXXMrZ6Qo5yfPoOXf5RXZC8/iwS9rg/4CgQXLqvYOu
aHgThVz1+5/WmemduewprFwg/Xwzo3DhWzZRbdgnkrO83L01kXohtjt1Fj8WnyCheTOZMpv4eo2w
IMeJMraUiW1+9Gozu8IZPqpZdCVYZkMqkkHzd9nG58oFH1p4TgyubufbbB7sx8TosDW7iZvefj5S
J5scjSSwiUEcX6+2fFUvt8nQ+FiJcRgvMjiZm99Gzp8hQNUYtVYqaKQHjohel3YkaIwSS/T5ryfF
5wNvJlN21a/aWrVlwtBVLokXA1pRdRr7SQ1Oo0P58MLfPFxEDPESRKsTCku9353U+rB5hYr0CUa1
itBxlWtiNTBn4C3RksPJ3vzNTHtAP4R2jd1+MHpJYF5TWxXr+eTbIuXb4MRfhRVdAl6TFH9bQ/RC
RNeJ5LUNIBMgGB2PTClpUaSpMJgqHeao6aNtxxunNvRQ7JSmgkgPTzdoSlZ7naWTQthKd3IHWH/Z
cZBtaSmRiYlC6Cf66+X2j/ORnPn+F6nVKPk1BySqX3i2Pz5fQMKijS7bq+StlFwhTwqBNTQYv1fV
xNfK5oPhxA8UvZ2xcOm3p6WLdf92Gagr3uORAQ08jdX3FPzSCkI0GuAKwM9L3z+D2opB7QsJ71TH
f9wxhj4tkcrSyiYcAtp21O3s6djBHVeFHkQzfneVfvmuV8sjH+tFrS9eWlEsMxV6x2/ev3vWrAPi
5CbgN/EjMwkfcbZeJ3gNO+HUrw/5HdVWTJrEmhzbik6SFizGdP74l7rcpguQxQgMi//CQiOWrPq1
lARU60WMaQB0fvdOGrRNsHeqsWN2OUiXr2EhJ/GKzhq53Hz+beN1YmoOUXREfurhIXWZYukFcuGU
VdR1mVfWD44w+t+HnQPurjrtr7KS2+5f0znAfFjSgK84O03Y4OgzRFidQIVHLSOz822FDuRGI6RL
QXLo7XWzE74vgua1nHp0R4vqvB/dbw+7hsKPmYU7/4D9sIawuRdlZmqeujpyB+WLwAVuxDLKiDNr
HMlKjIsbMeKh5azdloIW9PvGDaf3QLACtxUFFLP/Sl8c9HwxQoY9IT3sACCe2ivgzaYJyavZf22F
Tr/Q7B9EAxD9IBMv8SEG8aNpLIfRESLW7eBkylhNqcEPOT1RFCvwU+1R+JxMQOzrNrjV45zaQ01Z
FO2bhY2koppdVqbRjv4JRSbv5CeY7BB6rlWN93P9K0KKKITjiMO8/sA0gabZmzsxtE0Y54pWiQn5
TQnblObWWKDoHIlS0MQY9tD9B0Eg7ab8r71esFGFeMZDm635nKA/J9CC6Uda0Dd8W939PSvHBOzE
rJInpbGnzQz0S3a1AKZA4/+aokvRBtoVANaqarlLpRrVh1xSi/8Cqm/ePyECCMjH8Vs5rAe8SZ9O
WkSBP5DxuYLQA+wcPGkN5gORE5C/4YtJARurtBUBxrO4SP1mRwmTROuDFwyvfkYFLrUjxg9KqSBH
ACcfLBxT2XxpGnfoBwc62AeVUt4d5FmKO+PGUj/zG3jqOrDl9aCvRKkamWhzn/hd0+oQRCuLE43v
YrCgJU+qa53dLDFgkr/3QvbMhYSQNM1SilUxZlEBDdlTKt7CRKfSmq8jSNT1lDNeLUV1Wyd/pVgE
AN/OLM/5tF1r7gtU/ZKJXVGipccw5MxwN1MzDANaK7mj0edlxYyyO73z+7kU6nGo0kHzpnNnJ9Xu
NcC8T9aQ94fpJqAht8ARUhS45sVnb+4+UCTq2Yz0jwSm3SYXENvvh15mR694n4gjW4pyfeMVd37N
7ggvIRbsoYQipy57jn88dJQUnA2ieH5xl7SQoRBBaUu+TDLD759UVC+x9mQWsi3kF+Mtz5xyFhTP
QXoKLLjpiCLnocVDyuxcvD40BK8NbR7A5EkQl8mDJZ9tA7/Orb13/izfRoM3Z2lxZKY3uG5s7N+g
HvKNRPE+kIa9l0Px6ACoX4Jqm/ItwLJYSygXthMPkO1bCYCyztkGookxZk+9x+LwE/HjOsWNOfVE
LfpVMYQdKaFB8eKVF6XvKMQuaqXvyCoCAXRnVm7e3yY/i+CfuMCXyFYs2jbYukA5AZNEQhZSv9wQ
jnev9B6MuiSVfC/XyhZie6whxmZD0a5vC9qg6Y+fymWjQzBPOqOpXCrs511QP6h6qVSE6s/pDNAz
lbG9exFumKR0f3k3yYAksMowzZEbQg4t9NG8WXtIVePF+lceQHyJUTpYBIRZ9388R6m+WV6BlHWg
Uxg1WvC4jQ69nOIlnpS3j4sSd/vmYH2EfRWz+Za2qUrrYo0biS4uST0dkmgvW2NKLRrNl9g6CeJF
Pt9eArxpU4EKRFkQJJVNen7kTsfbIg2WsnY86GW6/jLXidqZPhdEdJWrmkH3NhX0y1pmEHG3p6NQ
JKm3aW6DCZ20F3HgInFgS4lLRY8XExu6t/Mi8Wd0DGvOO5XWTymAAg8H2+ckPpPKh3hmsmgEGqM0
stVcAPWfLVO1KfMoDhmrH9QsqRRnyTgFDhqOvQrB7jBjwbieXeQ8knRlQSZ4hbYOLVkrt8Xwv0eF
2kYVSAdNVKVZk5z/izEUs50VTS5wZcYwPau0Cit1y9IOVbOV8PjEmXVsjUF7T7tHPKU29MZSLN+1
6FoEXPS+HKxVsLvE3nKLYR84igsWlyA5vqDTaxgMcxXB1axfM5zxmZuvi1gtMDzxNeDpKLp+2RQq
BbpcHsLD4Pdo2BFAoj/0z//hyQe4wWrZ0gS5al4IaURxbOgK+ePVvG5lebgUCSO/bhTZRv3z5gm0
aj3S1Nomn6VNldM2mxkwlfcXTMC33yzmI/PNtbf9QA6kuziptj2foH8/ZkbHzhB0Nb7u73pUW6cP
vZ4Hx8VxfggaxPYW2WdaBz/MWOw0+ATpT69R2653QdxXFZ0QpNRDrtbHzPMI7Klz2lemoyIytMFr
LAjdU55ffsflsjluDjREfg7fmIpjZ9P/SNrzaDv5uSUPCAXB8E2j7SAUh6v+0VTXUksfRh/bSd0+
NhuL5PkUYqeZtXV943ilNBhajGmCOjedRGl0ZejjlXqUaZqrjcbafE+nTXWGJAbBYLLfIC68dvpv
2WzMPDVBEsL/tC4fWc1jCNSb1+HM0YHB43isMKoxtcaOZBqLHnUnNwagIlM8mgWAG8PrfRUmX8g+
khg5isNBn8vaNk6DO0JY3XktCu1Wu4pLc531YsxGzoBHdmBZXVtC0cdRqCIfG0C/iX+QqPNPJLJQ
3pFvd0D7tSGLK/Gc1MXIBGTSFaBG/O+o+VRV3OxcNt45Mp4/su57YeJ0n7g6r/SsGuDttFWD3ZU5
xeXguYPHParH3mqIXiYo6yJMSQjiuo4eFFxUV/m87YDXCxhBlcpUG7QEAH2zRTUbZuEy7ruE3czN
nfTmCAZY+DpPmnBI2jZW6FQTT73u5OTzMOCO9M3Qsq5RTp3+6ofueMXi8w8zNdg3E+0nHk1ld0ag
/Y7mNG/lf3+KggzY8ouZZJ1DEUOjEHx8h3Evq3PF82M29pYFe9CdFpkqgbsC2mSMJYMjgm2i+BIQ
2JPB7CsDOOIyI1S856d+odHyvH7UoizkXUa9afWlJKd5ofQosUsAb+AVQ3qOhs6916e6kjM+WzWO
8ke0ZXTsbIG/i9Zb2Jc9961WrNepELyxOaL9M5PYGP6/KBcQE2RebGjZZCdTeBv0JWHhpdO/3b98
au13TDPHp6NhVWysYgoi6pbyH4oPZ1PAWjOCI6YhLnlGeCxeHxFXsyiZ2PgjBc/PQHV4abtYU74y
ZqQSZzh9xqz07E0yAeFfES+T0+EBxdLWGra/FwAXDBjHzx4AMhSEDu91MMs+1j4fxC4vuxaH9AbG
vw3LFUPNqAL4O32ZuFBYodUFT6XR9n80t5ahVn9YCEMCmjZ4d+aYOB6rakxyaBj10qCsIZthcw18
UHLkN8fuT74IYkpVsQQfNVUedgoCx2qlmlA69w/pGYKRnZHo1IXoQW3GSR1x71TkAF5LMe81NIIc
TKYoDLyBP32dY5b0bmfssd61gaoNVvTsiqWpBWV+gSxr+UO88cwD6JuhCf8miI+yiwrZ1JoRumcf
O1+cS9NokJyWAPE9PrnRQ1pq08fICgkofo6Naue/8n5YzFk4of5pymYuewSrmm9gE1Fq1gp31o9E
z1u0UjgRKhfHXaZgq92munHrc12o7Rh04RM2kdtS2HTjbuiSm93tLyyF9Yl/g7Lyw58N6lLnC2M9
fDtLjlqCBrkU5ugRI2bwEAThur2p3nvO0Hq8Cqh+5bFB5tbPNN7U8sTD5h9K+5iHdX9Sc+Gk11pA
oclCu7kzHGbjTACJ4lXNvQMdU6bieaP8opzWdOHHk3kydlMaXPK7UqVNcGL4co7fAMa+bCUWcfRD
kHAzoI73kwNUzVsyAIdVAUGanMy+YJ/2R5OWBekh2TP2smdYi44wCIHukI833/UjA5epe17xOs9v
hp9G1LyF7bhMsr8M4DE5iw8ib1Ew9Rru+3apTyQQ5KVQI9h9thu4fXipfwl6S+10/qzl3fSnrdE/
2XCYcprE+uTM+8JsTWkUX5hjairAoDQ+6A8nRmvlZ9kpzPICmzH0kU6yBP/ZVCeik8KvzfqdVlhA
TKRSYgPDb4rwj84uT9rGhRftaCANurpYwjjs+ag1963r8wtc+Pfy4fOS27Ig9hnAw6DXt+NcPsp2
COUHt8pq86HGR6jDALtkRPvNgNPAe+SGf+Lh5B4d193h4IvAYHb6smd/gbLu5W0A6aMBXlALGFzu
81QqkPbGQXL4soSoD7rxEofBkRo/TdygPZkFcPMXZJbAiqhg9nOJ1GaL+7VPKFA+q5bss5NR4E+D
ai0KgSBDtSA+g4eNcytgaGic/d3MUYMHxPlUTyLWIR0LwYZr2TvMMXFoWYGGboAuUtFxOds+PQvD
gMr3AuizK5yLgmc+9lbfKXOYyAVA7gbG06hLvWq54s646B4Al8gCuQ4eC/D3SRwgMoxIa/sWNYt0
6ovv7AwFzc28s/omEfWvsjpFxJmAPhiXcgwaxijvPfXAtWgbgzXDexcXtWQXWKsZ8aSlefqagihV
qrg4PL/TfzVO3Em5Zad3dHjkL7tMMCBliDvpGomMICSG/GfZGfFAnAAKHld40zvrYuJMfLXXPuO3
g5XRvItBLVUpTza0EU+bizjkHpnF0PlT2i6xxo20/Wui3jB8l9914ZsjsUQvR2BBp57MFzjt8jJA
OnOfWxF25DFFbi+nsGgsLfpCB8+cfQPwb3Bwxrf9jtJnOD7TROnSNPIacAwTMSuq5WqCwG+84zHz
k/W+sC+tkuNMMcP36BP4sQ+eP1fxIwqshY/FdfMc/eUbATDFSg7XrLeWjdo4BLEg7rvJNrP5HbZH
JCr3w5WpCJh96TKIpFMM1Hq6vEorZnzj2hFvSFlQkLQJvE10NtlZaTxgzCh3JcSbLNspDdlMvGfd
WYT6n/Q+hvqgwal3ajEgkJVVUG640ICOn+VR3CY6nykWSmh+mPeEOX66s96vZKrgCW9a4UVvshg9
UZ2ni8fKwoHdwFobjvrx/PUwyJZRQQeCy9Y8xNjA6MKASrOE6Z5KK98mJ9Kzdznd0KYSQSBdFDcP
KYD9sxvN1/I9vK9f7p5y1lJrdlSPZgrdTN8jvWHFpXc1v1k3pVEUvv61/uxeiUyaUjhONwNlD8KD
fus0/ZC8KuR6mR5sZhPcZKYFV4hhDX6tPgEnGLR11MXdxe57W7UWgrImFBSDAknCLxTOQkvBSitO
1pdxrkI3iZ7d7Y5KXruOwv38Dr/gyWZenvBlwWwVbATnRRcqMz2D1EYFSvUiUw8ENNPbgyDT4ST+
z8U32YVYMjf2Y7QRM8vCcQbN/V78frazXSRiQ9V9ZeW9TYZ6LPb2RpRtclBdxYgfkc40BzUD2lwq
o3JuV9Tm7inzTLnXjtDBcuCTeH021tNvhkcrxtxzvKTBS2gL2SGBQMzapRWpm5THHxxKeix6yv/V
xLjm+b66gABHBWa50AlihpatIhNUnrmHskLnEBzmdqV8VXpLKbPZDeB2rBAFwKEi+kig1/ou5oGE
W31mo7RSeYq4jbqnyAAyt5L/0RArtLS64HgI8Yt3y5BtekfyUIzIlODfn4PTmZG5dBI3ZQ8lYGpo
MmZ7N91F4HD7CifExQxoUwiDgYHE3eW0V9+EjNWtHs3p6970/TzRoDHcxJm9BwoRaEEBUiL5NKRj
9ISs9DJbnkqrpoDqc8EbxP/i65mVhLk7XM91mtWic9P6IrZsY/9IlaMm/of/V7GMfup/cWVC/x9a
zLdWVeI95j9nYRbmipiahnATrB17zVTqqgo8N1g+7QWke/FD/cPNiQoLo7pVR1jBOl10QMIWMG4/
XqFpHpaR9udQh96uG76mex0o5CwG2Z7l3YlrmE9r19KBzOQk3nwARqPgwv1VmOm9IltvZTxGGRUp
lvuQx2uKJv0OwmTQHJkcYWHOZwOhMaUVwVDk4jDQ/5XN4sfEU5TLpNwFEdZCHqSHT7rKrz1uBZR5
n4Ej/gKEmVFv9r5V//NbhXG1wyaAHNT0rvoDXfWnYzE/+Ag+Pd7eObjGkr44unoDevt/8IxByFxc
X8mJopEQWKT8pdQlTWZCrjb18JNrxj6Yr3EnaIEjSPJ/lDTmRKs/YpJKhURTab4CtBE4x03tzoJm
M3YrF9bWZ7KyPbnmDHAubuDR6IyEznWlzsYuQLwNpuzE+TTuFl23Orj3kMjlLxDwIiKWml3Ubhon
uXgzVZJD1ELME4RzRJPfceav6U/sTiQF19Y+kQ+qcVuDyQfCEC0yErDMk40Q3ATPPkGH5Hm2pAp4
07pjCEVe23RkyE4T3z+1RqZnSXlt0UAvFKYzM+WzjCpczrRWj1C6eyxCP2BZ+CzMcBCSMqVjgRzD
V/ybDDr+F3Vsc9MyXCmrQj67fbt/8v0vKNNt93o8+NxDGjFK0qQ7opFB7tBwo6AhkrQSBKPR5dqM
3rdmB5d/6Ev3Ivy1eUBhCdMteBnVi2J8NYPRraH5IBzde8eJKUTrlsGtLzfy0Zc0H7pPMHDhsj2l
e8b50GGuQ9dkx1kKsDykjY6Tgfad3p38CPmvA2Sxtschmnxn8ytyOpI5NUYuCj/qEk8P3Uue7FGZ
uiOxue0M0Em+HCSktKhSWqAtj+/p3CW6qfqXIpyh7mMo5is3TpQfRIJ8zbOun/MtXknBSGHhC+y0
yXxyXxNP0jjx794sLrTzvqCkwSzL+E7TT3fteqD2nZPywbJ0ElxmyKvEEA1DUmbhH5arJP4wKYkc
S5gC/vwJs+Gl1vkXMOub7Twb/sf4+uOPbe3EavgBTKce1YLd6tvNhBnuKpjr4bhGb3P6lIuG9JOe
GMqZ+IuafCPhPnnVRIxyLM1VvgaOhMqGmq1moAn+qb3SztQN3HVzDQigeGyCevwEAXJ3eC0tM+jp
Hp9VqfUCgHwOCZqYzNGJGplHNw6NjS2wR0KCxuLj1JB+qs2BXLKqlUUUucirYlzzyHv4n0QJvyVH
j9zjDhn9LNfh478gOSUJS9jr6ZJx3NuSPjDIkDkBJCbzK0Vz85azpQc9/qcD4vfA5oB4nVKVJUry
f+tpLGGVstSAAVV2vbVgOv331xDPATU+sExVCyDp+2dVC4KieIbXAutBB0NzASDVxYdR/BsQwVT0
lFi7deG0v1K+9yAdPDvxN+Rh+cCFBf7H9Tb4xgOrDAsqQzxk/QRtRehENH8sdSVmj06r5zEgYYfL
EoF2W2V0OePCR3KVbOX0fjkvumwldE6ODRyhtp58Z9oPBiTZt5EXf7xE0h9Pf+AhC/ECG88cRCgu
tieFSwttIDhSODZPo67wKkw9zH4oRTeUouo5gcnSNmnnxGLK3aZYMDMYv2x+j0wil4JRSsbixgkt
6SKGo90j679Vkcw7mJ9iX7ezs8Ecq/qilk8sd7XicNtgMZCuw76YDGrw+N1u4snJWduCqoUpRU+i
mHwoWqKsOZJkYYumJxoYLASzZ9zsNBIpc01wBMxKr2sT0zBWGc47jctG5T3KTTFYE0J8r1VVy70I
MvACrJ6D0EjbAd/tp0Itd/8iTDgPVcyxvWT4xsegF3aLCEQp/kpEw+k0oN5msWLyW6XXRQBx1jbx
hLfQQgYPzcm1eiZenFFrnoidjPaAERhK8aJjWVn2zQC+BMuGYO+55J88aojs3fB7peL2zKWPkY/u
JylqdwsUbOTTZwlT9Dpmk7zscCF6Z9GH2ayy5ZAS6fYZef1sHdSBT/4DJKXyI+mhhwV4hty/QsKi
0dC+hAi5hZ3ndM0vfOO3vFcqRb2u5YMj/ckQf5yVepUIflT5XX0xL/S8E6o8zJY8a3W6Of+U9yYt
9xwJf0wngv0KqaS5J84PvmDUYnaove6TSi2y6YPcyu6a2NfcTWM++kMwkhGGGHZiAcNtI34OasCX
7MLa3X7hfile8n/M5u8piiZibJ2rfkv8ilYWE2oRQ72rqsEuM5RxDUQjPAQ1SIO522GaDqSJGGYX
wLi5XPNERWd95lQiK7lugt2Q5Mpuc8uwnCUl0vfhDvlvydQUWFieBCq6C9+TlGdXGImBXH3yXdVI
9Vs9GpfvFQaRx/xvHUjxi8UKgKSnVGRkqcccmOx2wsu4pyaow4FZtqMvXgzDt4dikjOgmnB+2qdE
hKn0RCkp7DQGqrD1N+g6T4JyVhgVtxZpsWvh9Da2XEbnO9/IyaFHnOEKM6cq6psXqsdxtl1/hnp7
f9SULjHW3/BO7Kb5VszTG5BbZx2tDhdYiXMJWEmekEHjJQCj2XA58IBhWoD2s/62NJjp1EjAOD0H
DWRPj2EdwYPDNAvqRZZOegrTNJfsol9NWYgN+VLxktbNjg6Z9Tx+R8+ppSdRVRI2d+EwqUFPV+xs
TY8OfGXnZomt0MmeXjP2QEM6Zctx6ieb2TCHI08b5oe4qopRG+lOFvOJEnU6VswfJRXMMwRhU2ve
D+LRCamc9jpkrp/1IwubzTo1I/ERaCl5vMOFfCYUb0UhJQ1eyJztFyYpX27C2vovy/cz5PCk1Eyp
7YmYLEs2B0IgDccKOz91bGrI1X08Ip1ErEqGkfA1D81WOiyzC3plDRW0XE2DCOyKzPV0XOSSL3Fx
VC+m7+VYrTf7ZWubNN9tYsTnHmHRGE5taDMIZZpwB1NWlH4kTv9+cGDJ6lP/kQb05SI33kPCM12h
STkBSDHcMll7UfgdymrDNAc8pykGR5XwvuHPtHFnClolDmv4t3UjkJ2GdFQLPGGRazqVw/jtwuyG
XXLwLwO9qSiVVNld8ARQT0mBWV2NesXqhzLD9tCn4EREoeWiIx6trTCTbbn1FHdPFTnwSie8eKDx
V1K4Ubxk3mUv65ZwW6mzi3e5di2EmiLPFk9rQqD39vKwCHcVEIA/Ej9sdqTSeSgryw7HqxTUaVfp
7BhZJX5823eaXlwtghW3AbMTjbLUOOeDRg3jg1Q0L829YZHUv/ZDW+06ipIFTcPUlmHSnvTQOWzt
Dy3oka1H7BrBz8z4njP8AKVI3+MC5GpEhvjX2zLFiepu9KSSHBY22YsMi8JQC8uQ6Te1RyBwI9CG
NRl0jscMXwmSBdbYbFgMvO87ohSYaaN0hWvPz/1JRouweuQmWIC0LHg+NrznKIUwrm2feNfEirnZ
BhijsvTlbCrOaO/MK0rkXqBGL9ZAGjbOOxE1SXworae2MNqdpCOvKkAih7zMB63yQBmTh/pl1Mpk
nrC/ORNTiQCww9jiixp3ytJ3QLWJi3qXvnDeqa2WtA6IciKHHwpuIHZj+Q6TUYUoMyJNvgAktGOv
4wB33QY5Y83h9SzNc03BzdNqGx8NkFL9WOychCAncm9obhbxhDB/3ZQXUfEH4DnYHMkQ2VzphT91
LTH7i8XYm0i04tyki7b4GBScViSwBMBtgX/j9qxQFeIp+RrW2yGfhntiRuaUXZsRoFhrIwQC2IOS
IArwzidjMQpaCdnkfjrnMZqmkiHFF6HN1dDtZwMI8Rjh8unHeko9W+40mxhBSuMJMmSRXFxjyvCj
/P9VfDH7WXLQ8WAcl8qAWnfV7ysiiRrOck5IDfn5vH+wVgW66PNqEbzIclmWKIucJNYRYxQP2vug
TC27999HnaSCC/f1uF1Y5jAioH4QzKawU0WJumiZkHOidwXio6ygwz6VpiW9hMZUYAAiRrK6X3TV
AIImLeV99CXDW3RVEl4Zl5q3IKxswcwg/JSBeJmCdyvV9wGaWGC6sj1DxEHOiLFJZRlNfIvzwDf4
B+0b4eRpsBJoWKx6UsqB1nVU9nV9o7HoC3Ht6y6Db+eu6pfML3wwrMJ4e/LvUhkNqx3u8BEPPvNH
Rda+m2c5+fq5o0DtX7ZVgRLi/M+1LYfo5oNixjn9Jam8KtuiU4BmTY8/aElxigx6uk18DCaoazmw
9Lz2DCZSMztDt22RqRGKdqJNh3wP7SqwsijI5fdfHQnSZxJPwp7Vb8nVkOjibY4CF2PzL5ZCAZ4x
L0niSJc9YNo+rqtmAN57dpO8pOekT899Pc0ms/2LsV5fcKyemQExMENxD1aI9jIe4Rdkon5TjP7R
5qQOIEMaZjOpDtwluyT+DUTvP3mzT3YgPB1p6BI89vm0zLlCucgbtm8K8YL46+Y1+h0+H7+bNtBn
eqRBkksF8S9UFWzjiCs3UCgiURmmZd3d45F+aFENS+6uNWm3FL8xmuAdzr/zWQvppcmsKBDvwawP
oHeT9TOZnRORDY0+eFcisY15AoZOoJk9yU2rr7gAFKRyVZz5Be6cKedsu4xUzTzp490v9UhmOJTG
8Zsf1tK06Ev2e+qPUzFTlyqIM3GZ8f6XNTrbREs2gxw/FV7PgZn90ydPDQeCpDKPCjWARkbm7rdj
25jIpQOFkahjW3iJKX1mAA5Tk0h8BUz59RIiE94sQ7xDX0vR7BdKi2jKiYZPS5P3lBngdnnw5hdv
6oSBJx/btK6lbK5fsbrKEE5Othuo1XbBJTghBzq4SwhEJq8kvM6JLLuv5i/BGim8WjigKFNfsYRu
wM6TUNvcFEEwwQX/MbLXq9Tqm8VNMeubOurnXKWiKjuuXGgTUiRm62qysgJr0UvT/qHIHQ+FF2Q8
KOvzO8IkwNJ/rZS3uCtb+2LKdUE1DhJeIr/x/uzN3UuS7726CvB/BTncguGU+GbqXZb1Y99kM3GG
5sW23jtCsgDzu4jpBPwrQ+HzeOnjlQT9yyMf88c6pJUjfdcb81WEO5Feg2RXGsil2iYlhJeCHFPp
nWr+1Ef5tR+4WEyrkkGLuNwUs7OhKc8gJczyc9Be9Ckk3ZOyhHPvEc4qPnExnHr2tEqhREikJfJz
OloyJn1JNtOZCLgcZEL+Ko+67vpAgSeRCNyO8BJgC0BZsFTXc0fKMGrRucx5kaHlTgrcptizBHjT
mW5hK4n+jpYjlFyy6ItrTVJ3OhE4J0v7dc8Q6/Ir5CEFOX3U5j0PZNQ3dzcUZrNiymiuFSYuN0oT
1d036Ac7EwOmFDZzI/9E9vJyKeKHXNmVnb2E3LnQogut5Z3+y95kMWUlDtx/UMDxvkBh0Dy9CAAW
+7U35YjFgzMMLiVvDBO50jpYxOAuBH6hOgsFe7Q39J6aRSqQAYp2ccsPDSJKnZUXfQkXFRjPee5+
mi0YT2pQL+cENTI7Wt4K3V5IfA5TV0N+Wgr+NEQK/Ch2SwJMJDIifb1SE23wFMMAXcc251ANSa2P
0WINNYHbpvVTmlz2ijR6bN+uyfDFCu5L+opRYnz/UV8YMHa5arRmA3nqcjxgzVggW5gJU1V1wq6j
u0q4q/vrbzgU5tuVdsAk1bV3fiONUqqraRgIyMvyPrSNwrDW0G1j2DJBu6t2zaHHr2DwWf6Z7DyN
REMLTutMd7inN+TQojGQd9Sv6PLlWj4HUQuOURwaeF/ozGhrZGeoEn7O9L+sKjxp6VbH4uuX6JWz
KDL3EUDEsQPQ2ZhHpU1sEHIKbWt3Ugy8BsKYTLuYGtpbcQh6P1rlYa+Q32wUOJC59lqCdKSsyo/p
wjaTABIydqXGoSWV5INpdH5CZFSm0TRhE4iwwmFQPiTN/lHhBY6SgxDWHk2/GHQ3NCEXfPfd/BPH
eTmOHccEgZiVi07LjoQVpRDv2eE5Dbk6axBqzN+cbC9YV8jYFwJBVnhnA5nhm+1j7gJxPGcpA47F
ZkHn9Sn99ndL2yoLi6AcPmgkr585R3CUQVIOT/qriwUFVcXN/wwrj6pUS+b5f/78RVGv7adWVO/f
Ar3zd71fDea1YUiwHMxNj2cozyeuJiDKiKZGm1lrwHEMl2/MvG78Wr+W2bK43OcnmAOKR8+O9PEj
omiadVPjQSz8Wsdk0CNvp6OjHby+D2pO0w9b8Xs7gZ3wwJwe/ZmrHNMaSAu6zbCoYqcfrffBKwlQ
buNA4REfYG+q58WB53WTkR/+Cj73GBKzrugoveTBYI+iXw+INMD73n97PuhZI05iK78oL9gkzr9T
grtCCfnsp8ceD/kJoWbwyeIVzDdk5QlOwgrTE0XvMaYco2MZYwBxf4U+NI3IYEXJaALxWihPyFhB
xhcyOtFUMRNaUaymologR4rmKA5Sdrd2i4KOJGM6HoTanhFoQwoYK1GMxCRtsdR/xR3rQJFEkqnJ
/gLJAlznSBWGVPf1G2zInH5RE81W2c+SYpOCv/BRdDmfGE+FtPQMMY/VdFx4WvOwZFjdw0rjYXzP
Fu75XiA0aWKtIzI5on7F4oBdof0i7j+7zAROc8qo2+yaVk2hZbfLNZ60DXWm4aVlpoBtHikDMHUD
aV6jAlH1/osjO+/zkAj4FfoN0PgNM+N+0Ywu2ww3U3w+YFNINybPyyJUteS8nNq/7CkNjm8F5mxV
fKCHGu8LhYzbiJvT7H7UwUBoBIcaf/FHsVFAxDFkW7Sdo3dRiJMlypxamAAEZEIkbCE7xTE1/h0/
Ds3UJ/zJ2ETzKIl7qiH20eIEq2DcoT1rDK8ENv5XYyr9VFl6OeJPZdmh4IBOo6p7WlweOrnVbt8K
QNKBdQoAUQEFfkQP+X+06xSagkJuDa4P/htw5CZ/IQIefPfbcPBwZX77lvLG9KRdYonZPBJE0wr8
VqCzbbLiI2J38r0iKfkzLoAKxRrFdghLx3WNMsQgJT8Yli1Ss/Wy27kvKAT5XnmUKDl6UcxEfsEh
vKRskQnURI/+NyyC/X9OQwlTdjJQUl7xHPS8Z6E4MxIpylrSw+K51Klg6IcSEhNcKcfykpnQg/vZ
5e4UspEGzjDgy3KRI2wPkWIElZLyqoCizWUGhGq7RaAgCReDQBroJQ9f7qFFoobiWMItUDibV9wh
z4xrjR8O4/vRqpZ7J1MAQbvh9na/kBdS05NJ+JzINcNdIZemYVuZLb9E/BtFvC1mcXf8xbw2MjIz
l2ddKN95p/G7iXlm3qFrIpQoroM7XhjyTsHq6/kMVBVOqLtecpTGQUe3DbgzCi5cBjkqL4mWZZ1l
yeaWee3WgEBITaJToSL7lixFGu8qEj0R6t300PL6CCtn/TLlELEK9XFyk4EJJ4UED5piTcPMNNI3
B8dUWs1KYvy8xMg7i7yQsZFrBz4yqh/eIbNM1FbA7IB5uf/woRjUnjR5r02jr0FoVsoq4px7GdST
x6lB17vKSIRqAah7oTfeTHoJHeBR3x/JdUzKr3U9dGIWikffdRjegZVFBGtwrMK5McjPsVczdZw+
vXrMSgIckSGk46d3L6U8jg+cGKhFxdvlL7O7j12wPWl8IOODUI7hanGp4QAzDdtCP4blUiGT1bno
dV3E0yRmssJlUykPH5HaKiqbc9iFMbidupuYhaBQ3/F4DDtWijhTDsjsU9NoPd3bAFq4+cap9zQ0
5RaZPbam19z9Jm/c48tMKbft6/lVsK+ocopR+ZnseVKX8r0pMWDBkIClIzAAASOZRAkb+6pkzvPH
nWkNJA0vcDz7CCaVSsmhBbfwnBXIh1wfBp1GWrfQIuz0l+vVUH2jjt1YuGFemDf4jzqaaT0/yjL0
uKJoba0WXduXLOgpdO0En6H2qsDgvzk1kOW6ADE3l3eIHbiMS+XVU5rghBIsQF4agi20Du9nSh+h
k7fFjqBNWJJX/w3ENqfZHOx9Pa1sb+oeXt/3f+zWf1qsNXKBMPl655DCh3RIXBceNYMpnkKpno7S
vLFRb0MfT5ZEN8XQEshoqUxfzi1grVj+fzRmxdUbpVsaXdV9t5KX+cNtPRCyfbGI+HJQbBbw03Jz
thv9pgyNWapJaiJi4ARFYFNzYMmQnv32+l6Cs/2KO8ucJeteR0k0UZcf2bDEFg+OIQ6Nf7GeSTue
QdmdtnC/q62O2m4JNpihI1+gZ7PUtEX9T4t2fD4C6zIydmaO73Blvzva0AsDvjCFKGwBT9fZE1Ac
X8uisT/BQ62ClwgJPpUKFQhcON2vz3pmhM8ve93Nyh/7QyWyNvMyY/prIiyj+8jEipsXC/UxqTUI
yzMtpRzHROf2mvMMGlNlTaL8I4/qqDutERz7y7qtJ0kWizqwSR41M02wfs2awrXQHqmIvXvMUfXT
Vq0nmyDgbtbZpSfDyJCaZe5ft3thZidE9pLvJp38Xs9JB38rx/F26Tdb4Y+eCVN8rem5uYQVKnTX
91DiKadjae7M9Jc6LNr/C6Z6h5yTba4GGK1Vw1DVScUTbl2SDx6SyIlcbS41CGv/v5RHvr0eXicH
mQ7lfTVe2ka7xMQzu1+7V2eDbIKgcvJxVEsmLjqTHDjUguJxbbEqMofcAsusgTze5vEhm8l8YJWZ
LkK+CG9voBk8dyRo1UzkGP0AmDZQUMpMyjusyf0CBSzNNhrIEJeuivpbnlB3qmzPT1GY92AV1mPK
clYrM2P+/f2XXLxWYGTB/kBN6WWJBXd3E5PQOTmNgaBHYWy9QAezNaIL2dXCysFzYSrMRf6+HJ9x
DQrOcRvzay2rGsBDLoWkgXnFCz5zjaKwVwWLq6LIO9KuDbNKNqxf8FY4OP1pm3HmTjVgI+aWIePE
7qDjfIx9J5l/YsMZipoyIUhg9rQVyzTCW5GOd67lCbGH/8JsOVinI6B2313CimjfowPQSrMO3y11
Mi2CnQCo/XvU3xRbp5m6mZQ1xhlRR3JT8slF+MJijyXCnauQL33YxCdDVN6xQIoGQNQg4kUNXEw0
zJDX0GySa0hR9nzFbFJ5NpUTXCqkvUD6p/NP05AdNtdtTwBJoKiQ09upu1ilQfONUEtw4NMadush
1hf44zLTJ3C4gah3xv1dWsouryx+78jBxHs2Sc5hwERSCupKXpzAJs3M5LLNAhe801p5um/Lx3mr
X8KDAoyjqxl4f+Is0iJWSqDKJawYjjJ/QrocmuI3IG/+Gg/6UQndcUTozqqV7WVTmkZXobh8q3jQ
YFfGuJZpH+h3hljuO2f9rbPkebopklPrHxLPtO9ayi5l4vqnGG1mGKUNysbLjbc49G+4cy9CDV8H
zmnsfks0FUd/wUTjM8WYafrgjs0xT4YpgTYKgQ2hmKcto59QmwYXNIgmKTkpMk3IiQUNbWgDdlEx
EL5Lwo47uHlPD9RFALbpG3b24B5C949q7g7crneFVm4cJS0AxEvHtqUYeUnvTcmaB3pUYT/PxNmv
LLbhIFPwpRpPpEyCLxVL+kebceIJnAyktnjkteP5Ct9WlvUw2hD/1kEYa75dzk5R5YiGJD3AYlPn
BsjzVzQw7mgKRlIA42kp1Gdyzl6uKDh5D0gxSO4ajHpLPqvaaIfJzmnr+3W+GGEcjfyNjF6bXqYq
aSwC/hdI0S1omRFKU+FXd2By//CntDpwvRT7UEv082Nu5SdL4IVcP5w26v3CDZELGLoAQ7JrNjUW
GI6JAfaCSRu2IoWNbgnbw760r/vzNybn4TmXLX0wEWtvx18PxnFSSWP6Rb17ejQq/ZjroPlQidj8
R44t2VPjmO9WZUUPOrC6b8K1n/AYDhhnNonIZNpK+QazsJCM9nB0CDjf0N6xDhYLy3MySgJvgd/+
g9B7NjDw+6W9raLB+2wnxc3i8RVucKrlO7vdSJIWQy0vXHAJl3566PxTAhcXTl2Gde0if34EZV27
iMDoAb6oYeiVoBmB01J6WrV29ydPle3U1V0nGtezstORFr2PHIwLDLKIkD0fNXHAvPpM7adOVfvl
Erm+nbKqBDR+dy314h1fnOufoshIBa1Vno048+Zg1WhWFBdpbya1Qn1v8tdZ5zeUrHyc/7O25gJ7
RqXTBWJ+u8zWtZw+ZXFrHzbBZxBSHO9wlRZQZECslm6DhdKLmpq8PasS4NkoJZgxNh8t0vJNdeUJ
4OVcPO4S/oVDbX5qFAynXEgaGFytinT3pJJwZKFWzMn04mImqJjFHL5u8Tx+EA1VbMgwfkETj7UC
Ff0H/hVudBXbyY9x4b07bMo95kzx9BuVEzZhkKYSMXD4u0N3Jxu0lm9fBh4hKAJIfYfEUI7bNSFE
fWx/CNKwenuLFAtmywJiX6phhtpyBtmO5jkUlwfh7YmYjTChvpA4HwzcH5X81XYpBJE1DIfmiuw0
OcWjq4TSqJoPS6jTy4oOgQgcIzIV8lUX1IBPZTCJIN9oGzfj8pviulKp8j6LFppsgj7C0jRRkZzp
g+zdXoEq2ZzrMjlED3ATEbieLwYMJAJKv/lVicD5mGI1kiurbCKurDi+dpmPMfsjZ+a2M5GnyQrK
HA2nrAnxRdSHglB1z2+mI5Lr7/3Rkp5I/Mp9pUWn72Y8Y+jqWHE3C3CBjT0jwci4Lw20NMsOOIil
geZsPO6fJI8dZMn8FcptWYroL3hBI404KRh6Tu7QX3msmryPHzRY1MAkdQiEi7VPrcN7gcCvH+7k
ni6ijsPI7cuWeoctemClklZ2SKFq4V3l8WsIlbm1bDo2nvHyDtW3y/vEFlpwRQP3rLAE4q2Gvv4P
+3GOc/Wu0yLCsMefJSoqH5/cRA9f2mT+h5vwXt2lr8OGxMHrZS3/iA0JfxZFk/f+r2JFZk7NiiRo
70/LLzVkW+CpQMZ573YehlYN7gJTnU1Nbdp+LZJ+0YCj5FcGlTE7pRUo2dxPofzP7GEPwqo1duf+
Ob/jPCDWqcDjnhLGblacr8NUeTf5RVzwF511gO7TiX7BaMPaYiOYjpDMvm4cw20/c24eGhsWPlqK
eMABkNNBuhaw++oyl4FfGMGBzFDsU78MQVl6pyjITRh7X+yyatYe432cy84VI8eU/kIOZSULKO2W
GERrT2P2Zz3Y0NESYiogGsc870aOYOnKswHdE9T+rdhaqRJ6x8TkZMu0zjWBdeMP5dG9JUH8ImB8
VkTF7ZCVrdpooAEsMwIsWhctclTkEXt42jPVOeYGtoF54WdxgVdBWk+IOkH1bNm4kr+nLKDt8hIY
QF2GU9r3D83gDDRCPw5r3C8t5vKN9JzYs3K2Sn/hsevj5ikRyy23DSmuhiAcC/JLFhQpLs1XPmgu
s+Me5zBVILVEbvenjh5zGWxurkvETcFtq8R8wF/rQVTmF2zsHmUESnk9XFLuj0UI76oHknACuC+D
06XB9ibd9/tauswZVl/NEpM4GtOXfXh10GURBOP4FkJ0AtzUofVyY6JqAIUZJ45lkkyBkAOsd6iP
rcbtdd25fJFeh14w2bOvSiZQt+9IIQHuyOtzGtqtKCfvvffvfeWRxhtYpFDf/MNVUGZkNyTD8IBN
EmpYVUEBuVVGpj/RRDzTLdvaZvBy6RRELUwiByFxdLJko4dchhNYkM3n4qOt5w3x7PTWEz4pqaHn
icHX7Q/aS5Xqn5XXaFMnnEoq7yRbIS9axTuU0SezmOI5YiOyxIaQCgf9u0xbT5HsFslcWS6ExDF2
0HWt41txaPqTqKtGkuuSZ3Q3GgJr+r9UvdVgqRO/cxkSYZiaM6krbzN/QPHcvi74ObwLfIqz0xnV
9SP3Q+s431EzVS4d7wRyzgzZX3kFgqA3unA+uaqV2qfwO5PQarLzJv2HSXjS3L7KooWCsDKRIZMd
iyRgy0uO4VRoaloYUJzLAZtGo3w3VRO60o5E6bETDeMTvQciXyZyObDqYdf6LuXJS2yNwXfu1oKJ
wfwnPb0rNcsrITv1pR2Ok+XoOq50ZXr7s1xENGabuKFbJuOn4LGah0nAq6xu15Y6GpHT1WL2EOIf
SR8aqMqo+YM8aJh402Uu7rbADQIKAKi/M2Q0n6B+wGcd5kGUhbXqPWZb1O/Dk3R54BqZ+Sbl1I4q
q5ANMQOYK+ra5yxbtwXKlpp3SEe9ghAG0qwOXtrjTNSeIskVlg/vdOfzfOinDyKyd0N9A7mT9xkx
+e6DqPadfJ3YlatvDNyNgZIFH95296SU/Gq8KqOSd2VjzMI/0TTXGAHCK4OwSpaU7+RRsJX6w9Am
5Y46AJUeKBjaFica7Y82U7uGJqq12J535qeoWspJ7dTU3evcVx3vvhOwzxrfZBn2Ct6hk5rxIPZ7
CDRkqegD6+G/j5JoSuZ7r0Kh7E2NsO8nJUv3IpqUbPYpv33F1/W0C/j3k3Z1ockCd+qi6dqRUSR8
8rBgmxkLalSMtS2lvlTzvZZoU9nEHpZTR7Dl5k5JXZeG+G1LT7DIKAO+khxAsq10KcP1TW9jThsB
+Q/l2xWKmuzr4SLIhdOEnPsqISkybeO0yE1Yzzw+vawzVizWIfaeM3Uyg3S8E2JvXeX+cE9D+7Mq
Sj8DWwhI6301wHzaH6JKNx1Hx1zskgfXUCJaEOgDKzVeHOFq8djxgXjztzmFssj7IQcCF6m1LzEh
5wDjVPExiiaH1xRxVI4NwbhYMJAiOYuAo9XJAUMxtTT3j8BhzlK9hdUCItnQYd26dFPHDmSngCNE
t7/Qj4d7pDZP7CqprdizjeRThh7G073QwYs3QHgQ+JrjhaXx+C3wOU5/WbeNF0CZ3gy2l2Aw1jPF
RD+K/jW1Kj6mI1u8RzXOvS+kAU8lWKSLcrelPvKianre0LOybGkBvZctM4tjW+hxYXRvtG4DArX2
gA2LAmcrGtqrRA4bpVKBFp/govuKxUjt3Oa/3AkTXPFuQZpcB6Aoy0B9RGB1/9puSOTk1mJ40IAF
xUITSS9DhpeRNoxC3bird8iEZC1b1lUUzDZDgc/jdn9IjCD4kxDPcK2y2Q2fV49re8ADFpsClJU6
7jB4OxeG59ScLqN8Qn4mPGFy+Q9iiVwShPm9OEm76BZcfdKA50csRiElZd8Db7KX6PTJOW2KAVAf
0kz50E3aEH+N2V3+rXOOOuZy7SwSVfHYr2BXklUjIovFqVAkP9zvARsP+FmF5dQbptOQyMm+yjFX
fCkIPNZ67Tuo5DfgFLGFxyxbs9XwXpumNr+4y6W/kbjabO3lpF5HLFHm8RqjtLyYWjgYDZkGNo8x
OIkGTB3snpNHIvUTLxk2dnvPn4rwaQxi7trgLOUhrAsPjjNVkKf5xG79SXfgd5h69FyaDK4FBspv
TcM9Bu5zSTvonbyASkEj5edQZu52+GA4ji82BmHgzwYflsUPpU85FRJ4Gn+n9Sm4O2XF7yS9lzYp
GADyxrU8gTBnLyZqbH81xWojxStuy4l8tzwSiuYh5xTe8viH0wfAOiPPu4Bpuoo4kDKRXQC/tJAA
38sGNlHwwtoBwL0VsbNwhVpbyyHRLtqvGub4i0LgmWWvRvZeOu53haS49uZL5C8bB3N1RTFx28J7
76rOwD8oGYxg+dPA0gtT7O+PLPOs19J93a9uZHV0DhF7RJK9SMLsrXKXssqheeau4UGd+52P3hHe
yW8761Vp63RB32JGgfY8nVJs6bfFSKVlF5HcIQ1UD7kib3yFBsWpeWwYOtP3Cas171ljf+jNbzIU
NjdqmmDPhQE3FfZ8Z6ow7CyG4fq86hVzpNYNPyskx0YrIaJZNDvVgYj97guiSPsPpYgYptKjCdDs
PbSFZNW6mzUWIbon7f7vQu6cYw5f91x8hdgWV3I6HwjBu473wIbZNc1SxhZLWS/3dgE4fRJw6Sdc
OGXdy+k7lXx4uMr5XgXcd6fI6VTsaIAse7Euz+6NBWNOvaYpv/VkCYZf/h4KHVnRG/p+vCBkFNzK
/JqvhLr7ox2glhNwAil1yvryNKBLJLee1B45vIthndEiVC4wLHIZqORCAl20pnPa/UkFAOaXlXIn
oKLLfjXJ9WHluHxVTxvsy0Dgc3bTAl1d3UeT1sypLLhfuMsUHuteuXFKWDz8RhDoEFx5d6WQGJ2f
Se5LogoHny7eAMFXTcReTA2l88ckVWrD7f4buldshvvhKF2h/I8lFTFyqtY2oPwAhlGanWVVZEHP
QQjjC0spKBTTmrx6HXMnLQyPnuAK1PzDwdJ2dxxwAHMr9UyBUXCjJfw8tV/6ywgDVuPf8hGhTAhS
jUvxMTNDngf7U4Pz8IhVWE3agCeToZUCVL4M0K4ZAmKghQoIgv5L/YVABduAuRmGBkL8H2BwCRo+
Un0TjP8PeXNtSUmyaew0kAaIJYxZiCZ6M5EowR3aKYSRsLWW8G/sTMH4cE3uDAoCbjWuQfkPZHVF
c8ZFo8gSHYa2aSMn1kOcyy1ZcxSN1ryuxDDll13+FDCPx6nRDRaYS0SuK3TaXmho/949S9cTeJRL
/9V3nwYXlOybMHKb1a082mX24IQTawjX0xvUrrE68DPuQWtpUT713rDl5gNtq2LZBYTR9d0b9eA5
F6lJ/eWYquaK7paf2CaiSVLo/CzM+P8gDAnsv3RiLFPs0QpTgy87Zjpoa/WPSUbyq7T8B7Cffjf1
GS5tn+hFjTY57A6M1D3UY+w1jiBSPzriLBMJMk7unymXjHgmEuTesgEUOqI/P7DmJEsnGieWfoo4
rCARiGdwCG0hyIrSBCYf82n23nvqrocytJegaRVwxlHpXkNYCqwfdWgQ8jPn19GPbjz9BL1DYXa3
m9xJxF1KrUFOgEs55NhehooPsNSJT8QUaw9nzT8cYHXRBg3QWR6IL5QNrNKc03Gs0IQyOQ1uqFj8
hkCzxDYMxCXie568ORj/dpOVNFWiEjXJ9mmhmYCc+YvsHC/w6JpGlVbOVYqgAEmTtgsmiaZcYjqJ
YcwlxMhb5D5MwAzkrBjTBfRQLiOA5SJNK4tHlFtQkIcOuFWUexOiGsZFC1q7FDR0s/qBYZoYT50K
5zALGSp1CbyTI1OqKOWajdUZcE/cv6Crk2rgj/26ZLGKYGFQKVVu8/tyZ2+QmrU4nHe+SFzRfVeL
d+zsRh61Jaen1skwb8KgKcEE9pLiAT39bB74OIClu0b0as6Wc5enL27Ppwz9vh5CRSS0uI4/gT4T
/108WxsDUeugLb2CTv1+SzdGZxKiAxpctOaVgohcTVP9ZKq8HXPGjg5Ha4dZy/mB/+MykubtwtDC
4RwPY0L24CT9GKNG+yTREGi1w4EzDmgq3bbF3ScphBGDXQkj9jF5f4nbOakKyjnw6MuBOeWHCQ4D
WsdcksGVIBlm6PZ7Q0dvlyr/no/Rb8XMi0gxqDFadWfAzr93fKrSITGF5kWHc3eYqsuEZYN/ja3P
JOZZjo4yC/3+RxaspMBBah04bliLojpque2TtiSi5spsn1W4eHspTnT9739/UWUChsMnyvRAdp6C
DEVhxAYTSWKsAY99rP8IsVdE8ez6wLKX8CO3vb5h4vz6Dy1eTSMFyH7yoXLVBLgKn8l15naUOEXR
ixRap2pFak7Ayt3/YrEwe2uW++fgZj+gwueQzU835yzbtMZhYwDWZPugKJZ0MjrUGaKpFbti9opv
biz3tZlr8QfRpmq1Ao6GYKFAisWjzFEykApdjMcRHQ6cB6lwHOs1Xw3EjEtzKb5vXDKx0J9fktgL
FrRLLAH6jcKg7vnRRCwwAMvdu3sqslKPmfszXcZDy33hRTVBasE81SiRNVWaIfcLaKk6Z1LaCvs9
bhp+7klmlqX9M+Hf7XVODqBOZ8XKnXiQqzyNRWBcj15JaESW0KYEH7CHBCUDEiX3ghl86vW7w552
X27OPCEpt3JuI10y0+TRLG0d/O8wHPEBFh0at8wyzK1Y4NFTc7LJaAz9UxuOG1spRhoDIHK7fy6C
0QEhQdaWvbDn1OhXXQtbNENivuKAGY9BwkGVrPJtX7O22xPE7cVUeKRjL9mUIOcofZoxgpLPf2Kz
KT9emmJaAmc/VyQJJ/NTucwXwYd7mT8FInjcjAYm7+pXqi3UZHRTQAZmLryuhXIcnfkHQTgU8Kyc
WZzGOqxY3PHndyZWhHsuZmVqmSHNHRfay+LXOz3bON83B53VHbQm2WpQK0zpHBLBQM+CdbRWyi2J
8BxrRd9xJlRL9a/1P+Cdz/bW0lfdJlVo2nfBVsUy3uFBV4nmS/1z1QKgVJMfj6PEdjuq8w6LK2D2
Al3IJ8IG8O0I1TzVxhQBs3C4VpCELlk3xx5G7oNUdPt9pgHX8CvAEhxqlqhQ6pGaFvO1hApwYVml
apgCK0lsuXskkg40j+TS3A/Bc6mbqVS14RB2ymHyj6+2AOAZvCN4kYNsXIB8hu5OF/aU6soS4mII
eb1803x3yZzhzInq0qjbHw6JWZCACwI8oTI+d1YAPieH7D/icyhTRcROOlcfA4L/rPTaU8yvj4mc
ErBNf/pkhcu63e8zs+n2uBgebmNcJ6Hb/96NXc53FKjnyOWvh1AE8tVVyZwdrsc9GGQTXI30QQL8
Al666wquYnq9WPcCSij07UyNYLmL8Yln1NEh8S+dIQ2yc7eToRQoqgvDGT3WkJI6D/baFl9DAOro
q1s7wyM8207EKH3RQNfQL0MP7DRtxJR09SM7Is8LE9HMtw7EFq9/VYp6h/QQ2uNJRCrjcwqWnTAh
Um6tqV2zcRDa2MniO6BvdjtspwamDlvfFc+CbmVEhJ8DoJujSYwhCviUAcTNaR6ocbiyw0SyOmkO
B2Aw7kUgNHw6qouD+vfDOstDu5vs55BgAMtUeIf1dGbCcYuC54TCzZ29Us7StXOkScXCCf3ZKRZ2
JVjpWGINx4kdpKR/iRRC0DPMhLKzeCnx97W0zu4g5LpoKjfgSSKxBa/4iqum1+Z3KcmlMve8tErL
WLi1UXlowYY+wBqn80UhflAeopV+G4z/zyDU6Liq2H/Dsx9qo+611Fdp7G5ggrkPq+4w6p4iZcT4
7ACM5DQ2Gix37iq9AFkGTn6u3THLFZBjny2e1mZ+jKt64ri0dkDCJ3lUzHx9/e0XzlafmfpzqHwu
6vuFohSKEL7ZUf1i0+85L+jzHLT4kIq+2OOVg1q+HTfqhEMUN8mAkNRBovDmLGTxXg5IuJnqWLMU
WYR6dP5iWa6k7s37SLJrTRsrJcEGJTnDbzqnlaBWFIM0eVGfl+cGlrwdTVdb7RwBAB9DZuqiKY4O
rJ/EAlYLUQ8b5lMeXw5ZxQMkNwyeUL9jQgKjDHVkDOzURp6BEq5sRPjc+kNizrC/+wuwPpNbWNl8
E75xs2laxmpyruSx32/8SK8uM/5QAyCCfxo6kuBUPF7Rr9OzBKGy11UixlCIRICGa1YL36cjuze6
TX3LJ5QMsAa8Hn62BSFD+tMln2GsTTDNN0adX0vGSjgh37tpkFbf9dB2iJjvzL7bEpuC64kZtZK9
ZlzEa36vtCI1HJBIlh54/y/HSaWZB2lw2SDvC6NvxNFAafh9CPdkvYr527Mp7Oe1+9nlLqwNoihf
Zc0bCm3WdtNEmtxT1PUpezduD52yBSYj024C7jGqEmGgHdSrJb5hii3wCem66RS6w/jaK+Qeb1b0
llDPU9peVL8m/jyV3BnwME7E1PxJwh+bCiwUevs+e21rL0LLTBg6O+TfPduqNXA6TNjvfuY549IW
IPdrkWKAr5jkFjtTSMWO9r6B4pQ6mjDn7cyB8xSwif/sTSfedXbDyjL0XAeEvVcYcRsaYhxGpJR9
ZQVwhtoh56/eFsykKluvIgp5Y1YGagG45PTh/eAVAnItOf4sVh8VZ+6X5EUyeh3NNd5DvnQ85kIC
wZlSwPBWoWGDSuCiGtBejh7WhlIfIJHD0lL5Mv/wrZ9zc52bXApLAChoH1Pdy4Zkuq0WzD+DGOVs
BcFE3uIn/HzCPId00avWPJkfLQlWzbNa2dZvqACntiGN7Ejge3b6gSE4+aqcV4fwORu8ZjW6cyrF
SZGYD+tz1JYFQXzwURF0lA2BwN1RLrYcTlncVqgT1Q/fQgRkb0NvQ22injmSWFUu9qXEiT1JEoJ+
2ZwyBr6dtE0/VMLu3IQGTRZv/MSH+UfOyG0Hxa9AazXq2GlRJQ2cfNrv2I2kyoREofNBB0f7WwL5
EhE2l/T2FjtAA6SQOISu6/N4CHIL9XYV5Z2Bb18FoGu3wur49yN5Pil8t+OWUI4J9MZFXvwFbOsV
iVEax2IULuPmqgd6aEQpeI8taufPVwT3jyzjrytx8tSpdg1SOvvrrVm7hHkWf/3ILEUDd2ys6Tpj
x3kBn1PlvqToqIKNfdGLplSCYjSH3e8NiytQMe46XWi27UE26yZw4uOTTuSUXDGmEQLGBzUYBfgk
7Td99YU7Uu/Fzw0DyDEV5tza1REY77/slOONH4qL4IhAvsSHCrCB/3GLVBmuFhqo95iQt4ZyV0oU
prpg7Zj8pQa0A5fFqHjWLqVYXoZXOjyh0YeXtI4TOdUf4RjJmucIqyulFuxY4e8LioYI9p9CIZf5
6SB+gPsTJ6/oGVli+qxyRb7c/JoTSzmm3RX05sRhFkC6YvxpmZYxuxCvjCBN2gaEQsDIVB8eIVBT
r+aNcqbiT2qPkAfki9FbqOS8h54jPf4oxekQWGpfhXLhJm/2TQ+k9OC+fiaX17ME0GKjPztQD6dv
WisgDdeR4LUH0XQ6fb6ZnQ1XwBCNuYHfz1Oe9+gEyU8YRKahmR9soTijYV085bDz7bX39XKh1e/G
YOVkHWg5j0WRiHjHKDisdDW5+WcDPGEJf8EADY5F95+AeHv2jbDaRjaMkVVj+i80/ajDaAxXa+q+
gZDm7Wr0HYojBTAMokNzggnAtbCbUf3mgskRS30SCkjTRY9+Ze9Tde/w3ppCNhBZzs1VxQiql2bB
H4wJyWu8zoLy716nAOVTr8JnhqP2QR9EyXc2ZfTOFbJGLoLaaCCVwx4f9RuzZ/ehrWmajy2A+8yv
hFPhddzfozhfdItH8fnDxOkqOCjDRPxGYTwBb07kznXcMusV7qa2jUW6qDjKJtzAKw3OynLAPtvh
JNdptumhfgzClMzIeZ+qd0WbUiMMX8vW4yY2DZMTzoK+zwdK8pJOfGIiDrHVnplIM21ubLSSSHHb
EDKTUlsbQd2Ko07dhEM62etSeZMzA8FmO4nV3PPsC8bsWIMvJG35TbeqCOA8C8PiyMrq60TMHQth
ZBAsXU7MEz8+hV5628R3DFhkbmkO8sKRpBpLrZLxfuWMULStsffdYoAdRAdyKLLf8D2wtYxCZU3O
9zg0gwgb2x2W0yI+cdbm2F4+pTdV4QHx0KVL3iEFx/WEsEjqxUDLaS9/9kFIMyWJ0+2uZwYM5gnO
nTxw/WMwoPR7+Bnk5z5KIt483Naa+vnMbkwZf+MxPprntQ0KCPfmX7eZur6PbWGCEa8U7PeNeFUf
UM/v/u7wK5J9wfrp3f2JGUa0Uv8f2ENBVHGfP/TgMAvCkEi1QT+ufwZRl8nrCjL7Tx5OG/1WcHTe
g1Xg91mnRKeSh4zIGqJ3sIL3LSnsxP4JiBSx5vG88GTZcmjru0S4xge84K21fCuFvtiRJG6msQE0
Cu8Cr1c4X0vKvt89atADIpnjQn+wtMz29sSpg2mEgB9u6HPj9d7JDARPBKpy1rmg5nuuJkDpI2+4
XD/yxmDU/P5O8FKMp50+gNda/Voz7TqNov6FhJMYYbzs0NHyDRN21MnjjqXgkKDLHlENGoygOBFe
SH8es7VovkHi4wd7Q5aOB2eJYTwMw9bGG/fEGuGSAhFW16HDrKvuaTd4USLWOvaH6WqG6ZzvtWCc
Ef4XGynZE3N35192O5u5WJUmaKFNzbT+GL2dvu4eY/9tFdw0HMFAk3ctJhnLByfU+bJi7eMWQ2PX
AcOLk5folJemUB3CnlneU+vO5L17n2wNmcGsRdImwlIM5rIiM0u4WfAU48an+b6Dkde3L/vTsR4W
+jof3T4B/N0APgchMv1gbd+lMD48S+1LmfhiwO4Yf03UQqgMO4QVhhczQgSPImJDLHGQMgmXfhzC
BHOyxH0qwCoeIb3yWHgMEJxkA7cPOS/y0QuSXfJ735yIsAou2psOZBkM+aM9FcjPJRPeViN29g6Y
cGMS++U0ClxaZnG6kywAmHSIDwRUEQl/diTUK0u92T/GrEVqTc1KSN94WNUtXjVUgKi6RJrQaa27
RHJsnNSyyxaDS1HO59ekwdQi1t4kH5lkaSmmZi2LCRxGkXcqEoOtC9r1vrkNZbtV2G5+vYZmfKiS
D58IqFfufzecesHGuxpvHUzpoLb8/j4GVpmM5+hoLwYE6eDJlofyaLBRbTF5t8Ra/SMusPIOfiMn
NSQFlhCB5CIr1lb7GPFJqkMVzzMQ3X+89RfjvyxcB8JPzNvi/OIZJQ/KV09Cy4ChHAyzRZZa5npa
CHO3W4FPoE0Wb6DnDkv0xFWTjW/rFOfLIZCqlGP+TWg510td2DtI/2L1YboKV0qD7dXBaAueYrvm
BQZBK3IEBTqhqrnSFQZATeDbDvmMC5xY2Bxd7tpluvgXkHXU0bvl7g2MQD9ROoYRQodMnrEM9CZR
gcxKr86Fb07S1PepoxEZ9JboX41KOV1FX1zwvP6rAT9F1fBrOtNSOjZi4bpkyWU3PBzzvN1g0Iyu
7MOx0TuZx0bOjM4Ao6fuNGHsoZXEfRi/o1xNixM1A/eqCKGefsU4KzLDXV7N64tV0ZjHNHgiCudh
QgmJd9Mj6NJ4PncwtcDVhZ2tS+jSLjXeQcaqEYbx+w/o7q0XuuSFSVn7TzW2BPM77qb7LDR3URwy
w1lmuZDhio+nZhwQu8jDfFGTQkavA6Cfhqh1uTQwjfJ4TdPK+qp42PsPO602iNGyBvjVgNxYA+AJ
YetSzRmuA4YLIFt67GzeR0a1x955xkZMEkuvgkbzXAVnWelFuaLgkDyB0jm9pwx6twvax8S5mI2L
mC7z9lprq1SHMDPmeYlMUC249Km0tBdDReCaTSXOBSfc3WVmm4jJwDSQi6SAj8okwbMYYxSgtjxj
KOrlINyYYQGgrRDbGM+l1Y5SmpVRUpiOgVPM0fmx1rWP+KauCyqKV8Hd9SNWjUOK/eg1tGP9GqaF
mNF0jzw4eFdCfV3zZY+rJ3rdGViTI5CWl+QjkAgWQfjfcEK18PufnavZB30u8NjhEWDja31GtSqs
2Jh5zOs4XPRkjijf59DAviVopUUZ3J3mwTn7OY4ZnKjt3RSqtJCn2Z93KQmPv5FBM8F2+pxYPTVV
0aBoRyJ92UPT4FhBmaAlflqQH/lF+xO0HFyara6lwmKlNoTMU1mS712dHVYDzS9LzNZl5zv2y4/n
MlmMAZh2Y8f6Tmn6GNfyPV1ErH/KfSlywwchbcf8TjzEFdUz7iFeLDFQapjuZwdDapao7UO77iKp
4pdi6/UxzyWi+mOfZWMjfUaddcu4CnG0qzeGairTABIxT6ABYVOWnmudjPVyHDxIFRUDWLNIb5/V
xNxKOWWNlmBFDSKgytMZjLRFJqyvpxxi5otAgD208IAUa9V2fpJ5v2bBIOfBlMEGh3I+bA2E3bWd
OSWLgyl/pda8+zX0nH8rtCh3nMQjdzEWSEsTAAjwYizGb80ZTDsm+4U3Xj3KQqOI7VQkmQdDCFZ+
MSFaJSNmsR4+N/qUGEJ9UUzt904hnHTDdi5Hvb0yKRLs0/kFIk4RdjqNar9rf4mbNKV48MBL8Ewf
YsHHQIQzDUPFdb/AuBMfJv0WBSbi7psqOHuqFOqsx1Q1heULwysnTNJ+TW4Oc5/CVIdpGSt/ni4W
R95K+3L8LybuGg4z/hfd71wIDy7pu7k1AYBC0oLlRmi3YA61aWtEMev116bWiJTJhxJZjZLqhd4a
6+/kg3b4I0g4fNszE06w6PLitCQD/0MsD70bye6jfmmBlf+POpvJEm92ugP7DDu17av07isI0cK5
dd6YGehZOr8X2/jIwu/9uiyb82ryP5jav5oUfUJ5I+1w2UgdKqXHVc3yBTn3KukHsvMsObVFW4CT
2V4sJsSvtK17iNSWIFm5YDxw7xWaNO9FerkZJvqsrZQYVAEr2GbzeLNTwT7O4jOO5Z1fJ02fJ8Yz
sQtJ6zv4XG4TICWxXPG/0j9VvVYRJc1ppdXlzttlk6LIjyMWOUuJQAh+D8kSCuxwsLwWX8NqfenY
HooKKa+AV0KtSqdsI8y2EPqjhOUYx7wr8Q9T93WEMEweXM5mIN7PtoJTtyyI85hfZIeM2dOZb4Tw
f1BCWI9jMRuZo5zEnNKcizd8reyQ7tSryxIHv8ETDqFZMiQnl7Nhe2a+imfUyeuFCbTdHDuhBuoB
oteT/K5j+XXDEfhApIS0yyyDsV2EfV1lrXV6L/sY9R4r3R2ipURZlbRQm8IAMw0xe/kcYqJT0V7r
EjUjV770ktuYPelcRLvallcVQ8WxOEJQn29sMCnUlE7RzL0rIDx+yONuQWJXbEvDFaNgWADjmA5O
7JsCBUi8S0bF6qsgOTmF72Es2LbLASD7YYnHOgvSCieA9/jhuStWjJ+b4hxAb9W69/oi47CRYMBU
HXbk1nDO9j2npzu35VcOAu3fFV9/7zT6Ucbap71muqMnchhb6krp61R8+H/dHQmag/8yq43mZHgL
UKgpd5qxu0hHqneJDuglJPnv9U5avaV+MPpbKrs8il8TK0yVAQxe4/hX6+3GjrFhfnavegTj0gw8
Txx4x6sXsyRYb0qkZGtB18ZYYH7QQ3Bc4vBoeJEO3z3k9PEVJ4ZMYqPmJPGGTfcTh6zeE29N4Pqo
7E4kpBt9tQ6Q6wS4JpVdSBPNhtuZ0BAhu+sd5Jq0AAsgSCW7NIuglduvJL6el69nMLz/jxAgdeaT
AAr8ERGoWbSVTvWQ6SpQ3Wl3q0w+0cXcaBfkTimqshArghdDEiSrebgzJmZhg53Ml0ELyArV3cSa
rKV18EN/h5WmcwJg8O2q80T7GJ1KNNY8T8H2XkqAsBUTJyEdI46dYAWUAPeOXgL0/cWsp7IUTKT/
kcwYuk9AvXw/Zb224YkRgcbZz41l394kOc9aLC96bX/C2eXnDFWxbvp4lA/+PjGQeP84L9pYrdAg
cbzQ+HZvy7wFc68/NAQfoF01LHdat1ADfXbiT2F4D812eiKbNLTQIiCdss2JCbO4d94vB3RcM2RZ
KW7HkX4D1shr6q7EVjnEBQcAi64FwvyLe7pJphcUO/OgFywK5qrkreaSovWBizmp5/3hQSPTrAAH
IKS0JY3hDJyEC2W/04LMHcxhoAPlL11Rg1sVyL7+8pgfWKMlDrMzYsgbPdIsD0b3+Es9rTE2EDX6
p2b2T/QtZRcPj03FFwOD/R8euYcjxyJBLrg05wEF07v8prmFdmCvVuKZ8YSVC4H1YUZjNKYbYavs
WwEsGsBMQrqYe+6Z2ErUGPrD5eUcke+UwHqBMqQhxb/V0lvNw+Qal8GwupmUG2GE4Ub2E0Gtj6zO
zyKA1/WknCNgaZewMRAMDNkKmzMe3rwUbaz+SAkFZERtO19v4nYDcizDUYH4WkM1P3eG2Y5dSu5R
JNOa2amLPQxszasjHJ0uJrsUC4GYhzDFvxYixFcq+wy/Xpn3QNLsl1z26utO5FtzLWxaGCf2kIRD
wVibm/dZX3LuqYIdKrLICariuenzaTtAVe4Y8eJLuVd8UZOsPq0HDKjexhsP8mw9kc77Cft26Xls
cEELpSLToOM5/iyMw4YPkiue+pQgs+s1eYchad2s6gOKKZku7uPKUtyPc3rficEACs8QbuCNHkza
ic0zunr57WxxhI4lFH2G857HUnhUsdBMKK6O5cZjiZnfSDK/9DUQJQnl5Mufm0EWE1KVj930ER+k
vf04rZtIz3JFEpjXj+q3GILdz667XqMOeBzOlhAb++aJPxhyIBbr7IBpp9BnPhkqjqTqTghGp/g9
PnfYk4RKEdL0F77EZmftN6x2RAUBknG/ddR5oyT98RjBZA8JL1GQSY+Js3W20KGqyQ0NCOzGtaox
ijGLI5sRHpCA+hHV9We4rGHKVwnIUxX8BZbITQxbjIm1rE5NCGLLP/19YN91bqXci7LCmznfh4O/
6m3V+tbv2VRjqluW1y8JgPrq/8tYl+pfKf6TSg6EA74ipBW6vousNggtmJZ4qQV6vA/hDNviZO0T
4bi2DFXT5QEanTxM/gccb494iXE4T0ruR9CJyCVQsFBnJz3biFBaPQmFKk2fsJMYDdvwdC9zjXU5
ahnsP9ZSu12ZMYiv05Cgi0MswShssC832o55j5sQHUb34i0qSX2RS+AdKfxvKYtxrmJJZlNPWn7z
2w1W4D5E7szXnvi3YEulA4L9Z71B+4p8LX1pxZchQk7/M9Vv/gAi4CipO2gR4fBwcHAOVzXC/BJf
Uwo6gaSY16xS1RC4vvGcGULVR9xx+CW5rLC90LASquCwFE97G/NsnmhIuubP1lM8DYBf/pZqgB3+
H5BY5I80DUTuQh4/qNB+v1HcImZYZzxN/DKt/AY1VvxJW0s9HkbaAbtDyhcoUPT3JyGsz63gLroz
yr8mNdUR99aOx1ZWPRiafeGab1Cmpfn9q1P1bICPQyOO5+9IEutwOVYUKdWmw8OJj7J7G8ZrGFdt
mry9req3K2EVv1RVZN0ObRdcf/c/1Olq5tLNPejaA0s9Ws+AUK3Kih0Xz5ZfzYCniKaD7krE2Mt6
KFk9Ra/pedWSaZ98JV1atPDfoBGG+WHsPCrr+qK33Y/KCPGkLm7Ta5hv++jb1zIvmH/aE0XBONLr
zEFN1XIXKlMZSq54y/q3gHZd3t2+yZe5LEmRbOLCuIFtTo31Vma7FeYjn+pF8/5o9cfqZSKvSv4h
929zaxTO2L69olBm1VlLOqeUxhxi9KZwkTzVDR/D2d8n+GHg0KMUXY5WITGhPpIl6iX12tVdfwbF
+7ZqBdIhBKidVMaklpmr3oO/wWOHzX0nKLNuEtW1y5mKcg4Yq+ElNE0Kpnb/dmYKMx1AFj6xBY9q
xLeEGxblzYZrq382Hxe+hV+pSopYTi5s1G268SjE/efxENDiDvvixoDwwLkfG6SU+OXKipOcknrl
+ev3J3FJ6uZ1fxMJ2ecR26OQOmkHa4pZHfPz8VXWT2uppRrbvNSRFPecEdJAo/4A5RZS16pMUrq8
a2OL+05kLSevGj8+SuZDi0fxSLQ5k/dMgXO/hjc1o0+MREdY+Jl/7wCQPEG7ffTxBoUouSPxdmnY
F0Dc/fs7VTIC0oYMuRzL2wXGifQfvXdbbDKVQXFrRLMWVpSeZN7p7TIDVcy0bkpcEHHnIpKxXRRv
rbMUJNe0xpub0FTLe06ObKW+O4xn1041GdhJB2FthbN2Ol5ObFNfp7MWSwkPxJXZin4YzqvmOvb5
Wgv5mD25X5qwOiOZdQCoq0Ul89P75QTFcrBRzg1P1pJmjfc+UE6STpWgcmX5X6/2jYRlG55CMg25
VA87AE0dSQKwq5L3INDa4Tm+SnpBwFfSU/XRClm1ABUe3rxZ80DkgHxI+cS6jpH/KGeQ4qYSzyA7
IaKikc4k/KkunhzHhufE3+p1VieJcu1Z+Ba65upNJfbHg7adoyGW2gTCCQuf8+GO6dMYjPvZmGhr
VL6B4Ug2t/9Hnv0HCgZiL6DsrorfNurW050Ph0xyMLb10nccl7IBHRUkJ0kQH9OATyPa9Kg1ELws
Ftq8wMDO/w4NFz3KxumAmlW3bpxp8kIA0Ow+E1CHoFx1OQ9pkm8FbIuR4JAmk9+H25NE2wFcabSe
V8sqt5s82XfPSFbIjiQYCJG1BuUr3jJ8uYsvuPYBR9AvxQugCVjzqBYb0bu3suEA2j4fsTy8tZ4U
o0UKiJalvSwevaDpueFcbXPVeNjyd/av1AaWGH/Cgf8z3zqVHdjz0WRdGiHSrniCzPtHg0CPSxkH
pESWQefn9CD7waiX+IcU1aoGhGbB94TXUiDZKXOwuCnN8v75KZjx0fJR9AjcZDDQYhQBJtA03mol
OqT+JlaX2iueEZDYulfWp/r19qwdBXlhhwLQw966lu5JuQnVzOd/LdfBM4y1iCq0blOANxC4d6bb
H0Y5CHCE6R/+efeauD4EKtve9EqMoxZ8hBsMeYQFruTyzEAKxsjb//tBxRo92h0Z6GdI447qg2Ob
rGIcU63FthkJEnrBwV1k4q75HUbRkDD9W+h+tKt7nxEjc8F+K8JomWGSg1l21CAnJCjhAOV7R8LQ
6l/M/HK30qa/rmmlWu/jxvo3tWfunIjI0Envr/lq+SlVZQ6HmZR9ngkxjOscEF4Kg8BOKMjGvBFl
sGmOnP0NenVWw2kPitRTmLziyvXVerOwVKdpbLGytvbYcqvneSyeiIS17yMEhavTJb4yCZOLuzxs
dQBtsIqdZ2ZDby6ybZlV8YvjlP89GhSkOpbXwSPl75qqlp83KuifsWQ1Fh71LQSL2zeh0I+u9KHX
KCh1BGxo3CKbymO9a2ul9Xzxy8TG4z3HFtXV4VsvGhCYVYLD9jFsQOBRrMXKqJyD8UPBnVqLPsKQ
Buk2vNnCVeZ/i8uFavwFayV1xLxQZBxiTiJuDRc3UxecUMmeeTaX6r76HGhzIXFmM2USYmPAN7Cr
yT1mpjztZpluf3PpVwhl0DdbN8jwu1T5gAdHToR8GVFxKLVl+NgC/RjxhQ3zDng3WaOGTYPOFeV2
gEIDn1o0rXaw8SD1zibr9hWualUkMkXapmROW5s+dTZZQ5BMZw3Wryz1BoEV2m5FgfHThcHY4a/8
5NGBRiX+4YzbDohlsP9gQYSy8uxcFyfLq8veeId+zJPAKYlI+ORs4vG0cWmCVkaxBDFoBEBpHZEK
NmNPjaY2IGAMHvomeKBEwQkF7BZFXU61IZJfBnM3i1ZRBW0VL9Mf4G9PvmnkegmkuMUqfu/Kvs7h
syPMzZ7tvlBomBWSHgchvBsBguLQli5jqK4p3wu2pavkDGdKRI79iKHg+lJDMg6Z3432hHwqaCNH
trGN/2wg/W55zB7ZpmJe3pJ+EN6G5A2p90bvfkBmGQo5y+9FTK2L1CIpa8oS4/kYZbgJBAhszTzI
MF8MgVOjEw2/N2NdTsRurTcJkVljswoC28m4rtGFhySKt2gmBqyzb7r8LmFZdSb3bKIc4CPcmISt
IW5hUYQtf8hGmy8zFNNu5nf2KxNOUQ7gGnqRkywBS+lQnWMYN9ImsWUJ6qlKQy/gC6LEytCdd4Et
zsOuPRgaolOJDcxjAequqelzho2zR+513t6PiLFvsocZMV2B+rlBCfl8d67fBbUEr2/TgQS0Q1sx
PoL9eewaeQLXmRtlfpr/s8vusoh9c3DcFievfQwgiKLj1Miq0bRtm0FcGy1PHJxIbV7lAtA6JbYY
VQLZIADApxDatHs+G/GaS2lH5jNwLdx3HcrukWLcJlhAFlanZIq19q8V/klAtWSIOuH/efEtbQVn
sVJhDlRmXt32snsB6PvtQhM61AHkZgPjgNKRhZvOkjQR5xTsCCH3clfbu8ueMkIFMzBpuXPdlIlB
NALcSq/vy9WZiwE3PVIytL0xDvLwfcvm6mk7wYqxwUzZ+/OB95RsdejWhizXyd2L/6yvQDMt5Trb
ls+2QnMldU/JEK0+pMkUWfTTGIkULJMH8YUfqqhkpTtG1W4bFjvK2Rz/9ZMIgkPiTXkCss9qdfE9
yJ5MXto62gBzTJ612YHtFqJw13fxBCCpy98Ee6N8XB4Q2+VSaXu2rv2V24vfXfTlHhHZkvwWyeYn
W55aP6Fi9rj7j0AA18wrnopUJ1+SwZ3I4zmMJw+9x5hQYJzuA0XMqs0ogGuUBF4H6YxmSmlm2CUW
C5dMlJPPO410m+BAL/mjzwch5Ai2mOraWhtKslPex4xgpTZExzWoGi3Vr2FDrfDi7V5vsPF0DAGr
FdUhEVsQtbJDpGyjpPh3RxwwhbCLoHtj1O9nEvDrNyZKH6e/tQnuezoOikziRYRLhlpXQmTh8Cfx
WtwVtyv3SROY1EBMTUVJZz3XYDH51k+4FxIqw6QEtNTnsY8XPjjtDy/OYWVdnOH8JXu/15C4Y1b0
+gblc9M4j4Rr29H1VXvNSeerJa9lPWikQY74GvrlBSLWpskvxDpx+xTVoViROZMNR9UZnz9bQ3Kd
w94EKCIHOQGaisEWtmJe03Dnd0qUjgw+xCt3bdOOd//w7uR2g+pJt3VQR9GRQTRnPr6A1v/ikY/y
QaqRHP2xRy/KgIPP7ia2ojD0kjVhd49n9K/dhBLj7jvu4DDpOp5hdLva6XtgmP81EioRtHTV9WNQ
Nkh971w+vqrL3QCvW9jB+Ho0603UiMjxjSkRTIgehpepKvUYOgRWZrPj6P48R/CkDCrnzZJLKtur
FI0C8+ApsJy2XqyUXYgQd6Ev9YdoD5LdhGN01QBVTe4EleEOHaKFnjhgI/JBPEkTB4botzlmdXZV
hcXai5UbRKrje7CPX9Y+Z2h+XP/ENLzQMViBHpYcn1TFdTngof6JTPJb4/PgWazVaF6V7oDKG8QO
N60bdmUnX1j8rbpcjXzdAu3lyEdapOU90FjNKoa6Bn/Cr4dF2yVic2Ku0CztEzTVLRtqMc9GxgAL
HzBznZThPAeFvydu5I194t+J51GrH9cJtaRYXulXcu1mB452xKAdmXEMzHLN2CwDMLcKjb06cLUe
eMJ6+vT6MrkpD9AV937Jl0jJ6OA8M3XdVK5wP28wbtiNNRmvS1YLYeyYMqS/aqCO+UDAo+QAQRCD
q+nieGlTR1CG8AMaWncWKhC4HbChLuPp6neTLVKA2FFu5YmGAxkQu+HRZ8jYnMVMQ3PpTJzWmILJ
0CRviFAfssdnbJObf8pSN18dL6s+LH/MzlOeHLE/+BDI3GuPkWDfSf6c4VaStxDZ/NXvl4wK8Tk5
R3z5A9n8QJPleth757r42TDPkFAeSUx2g82LzUdH9eKL6KsAGaRCdezit08NeL7zNrri162Fu6d2
k2QkVcW53T94TTEEOx3O6FB4iDJ+V3ts6DbmX0/qeAee+5P5J2NGUXyCNQ87BJMlfMUHZ26eIDjS
Is9XxB4w4ONlqAZssC4hUBVxOY+c3fpLA2UX/I+OAJ089Mxi1iS9g2P0B+SEHeni5XAn8nEs6LcI
GFV+O4o/iHhwuQgbHNGordkAeitfkgCs9/yT/8B7EuUpCnIS7cw+qmKisgZSAL2c513QU1y9W5pC
c8NAmZKs04vWNHTGIJ/vLBWiI5FpxrlAzaINr+zI1slLIejPld92PsLPSfFP2niYw0U872uEl649
CYH91pPFt3AfByQXmCFxpvHGsMOvxqU5eLq1yt3sicGMK0k1lJ5VY5s2jNh3glxfRxI0BTuoI1l+
WV8s8jQxolbS4orrbCjQNOJ+3MMD02fd4E0/7eWYUSH6Zhqv7Th6yGifABMHWH96FzaiLFqS9A7V
BeWMIXOxyYB8K74LSzlJi4zl3vWPlkdj8nRAKQSNq8YtFS7ohfsZclCY6ok+sxfuUIlKzN6rF+WS
Mfod3UtpJSLAlnCFMM8It3UNdUdsiNoDD8ZRMrOpMQ/BVuC/skuQJsT0KQ0vekomW9YJ4rySOW9B
7iaMl2QgzklhOU1NRrHqYuLh8eLH4Lcnrrb8qXOPFMhjL/5pUYvQt+g8bS/hhsGy1beLrghq1+T8
sUmIbUjx1LvTaFMbXhnDHB7V3cO++KpZGWoMXwPyIOjcFD0AapZA7PBUR200IqZehCzbC+aChtBc
jESbp1r8cqqBDR5vYj0TbauSr4p2a3OMgjxrYtqK7Zc028h9vEjR3FU2qqhhdebqkGSytonn8/lF
ujfMnqP5ntOF4zmQ6Yo0LMXGonKJvHeClv4wj8s9djgaWolkh1HSBYDjUzvezpuZYdGxTEcS/eE+
sFzjyVlDIjgAQ6Z4lAptxNaOdoaBipiSka7ioHjvxknqrG4v1Yf8ZRN4VZWXYpOz3GtY7rZmmjgJ
WJo5wO6YA3rRY4vMc/hojCCOcZwHz44osL/CP8a0SJNvGnFzNVAW9jZd894UJveF4RZHqOJ4bkCW
+kqEhVjk8NwGAcgPq9a0qf0MB54HucvVIutpN/13AHJE5x0Aq9/P4Fy0OVAw1wKuMSQ5NZ7rg5uW
yFsYh7pm1gILc0MWBO1AChBixgX+uvv6aquUtUtFmNnWtP2BPRmqr4fM2359XeuKPNKneN6+Nxc+
EyovOXfoxt5c2rmgM69MIvCdkCmM3BHOY+SNSbtdvUcrXpFz3osKBPVlfAggUz3Px3G1+jsoJFjK
JVBZn7ME+ajK65ZvRlwKLIYt11tVfFqQrGgw5/sVgCAGZ/hZbFC2wSuFWFWgGQvpxjwNk5eBoLvT
9zk1paazj7q2xQZJd9PTBGMBZfKOIM+sSzNMCfTVztkrYnf0rwwmMAIS0ZEbK6ldLTx2mN0cSQoZ
M/CbFlBCMeyLRloXOryGCHzFVPt+nX54mG2gJtD1KUfTDRye0yStw+JffJNE4e4zP+M31NAvJAGG
oSFDIXxWtkbWW3RbXvVwI4oAkW+Me9B8/f3bBruSh8zT141NslZTOHimio4FqbFEBNep+v2h5daj
/md1BRMm1P68UDW8hpmjq6GNCsyjhnH2QY718rGYf4F0Js7APoxU1yJw/ceWmUiXf4u6ftDzJc6z
OIp1RsZRMaLB61ja3rgc5GuYwg6bvA9IYpmWzg1qxTnwscXwK+wq/JZ42To+3g5p1ASjqefGzrfD
PSxODmKeXas8vOVi6dkPHr3ua06679+Klq2Xg4NWMySoY8sbSPV1atl8m0oD074oFtHNSye2PraT
pmcg4/ZzjFEmZtf+3r8qYgp8eoWmbx1kcq+6+6/x+fDdfVmk+ng3KEBRHdPkjEcLqt7jDq2msPd+
bwwBYauU/8IH7FOeWeH2EdwPwRWarkXvJjMBt3G8kmGQDm3v5bEa8NOYQr+HENiw/CJ2fL/EOao6
xTi6EExLpw+Bwkba7/uMCnsF9/lwj/bbisfmx8A+HVOwEukkWr9Y4fueXxkoY7y6AvDi/5mkMDF9
Q+riYtHVQkW+mKc67tchcgLX28y/VNFHCcghfN+Q2i3+6/++o2UBDo6UQuhCQGomjhwP94DOsV8+
w/XOQ36bdCRSqBfom9alx1TVEz+AQmblDmpugCmpptsD5ODoB4jsY96KA4UANph4QyEucnXuqp0h
IUWp2bytxuCEQ24dK455rpFm040zEBkxuHUKgJULi0ayit06GtFgP+y37mqvJ1S6UfvkLdkYho57
r+PvEC0g8sNBUtZR9TnGhycOMbAtiYjMQ/iC+cJqhfnYH3U4oAEmDpK/7sf87JJNj5B5pqc/vRJq
Ikoz04AksRXFpwlHLth9CuE2k1J6PDXyM+M0TjuHVXWkTCM6yOqNsJ+c6cdh9S7crszMuzpSITm0
FT6dSlGBXVStwsSBmYrNVZ5CFDlDjZAJSsF5IkkWW+hrNyuUQN86Vl8Aw59oH7eBbFrhXjJm+l1C
c6wi4tj2TPu8Xup7jElbfjKYp9gmvoC1VwSZ5D8ObxX8D3T5qCqWccVZvz19QSy0BWIqmubVdZ41
4AeDTol570U1TDC70Nh+u8JlB0Az8IaBxH6xS+2uEOwTPJnmInrh4HaQ+Y2TlfoKSnd27fsxFQMs
GAeNt7NZ5+GeUDwHn/gMSVIGvz/yYDUkxnD/bOaPENQYDEE42DZJ1d6uLl92wOBIHjGm7WDLSRqg
sUEQWPqHl+sPd7UV7LTYfxcR7RZDXWuiGzCPVAmskOJiYPvbgDUMXQGnhsJE3SWDwykdTjsuN8UX
PEPcB8sMqDeRgjhW2UJBATJnQB2Nzb7NYsjgg8ubtcsHzACxfCdn0UyF3QZ15URe0p1ZuuE3IrXF
us5yrjg9rWph+WwxCFHSJX7ROorkQNmwGNAn50Cfzf7qRWXjc24eIravnVLdHUL+wUGNXYoYhBRS
FhHlaMGr5iPOgLGja57IFAmEviZ4QSyA2Qta/9qmqIp/oiQDdH1PJyXnEs4KKuNzVRyNat2QG05X
fL+l2nQrHegR/bxfu30SgOw63S1TUjjZKzN2R1jGlWJJDM9BOQRaJKDKkYvefdsEpWdi+Pv50yMp
8TO0+nqP2QKTqJzjWWybVy4Di5BL6uMY+otwOvgbnbR/GrFEioBawNEFYpHsty8a/cCx/cNGniSD
qZwG67yo1g+QjZvMV/4p0bYPSPW7D/OgASxaRu8LOG4TVOD8YNLj/S3Sc/vahn+sN0kiAzN9J1rd
GBZ05Uv5D6If3gVpPs1xW3pzAKXMRM2i4fki11MGjaqFMkaZUFOfb6/Ps3AUoWnYSKKH16yi/rss
1G+4CEwrb0+t1JaXgbveyBFPGAlpZv3hKwhLDBL7kL4lpLE66KMyL+Cfu8oVj3w8EYfX85zaH0aj
0ypsEe06P/XjrZz6i0+OWYVTaDQCLNSV+6dG7OicNC1LsrnTYUr/RSwLaQhpjDvr+wnAjlMK6HFy
6RsuneWDu7s3aRJJuB43jDjeIdgyXvNM+RRnKyIN5oEipjDuszNV4uLbu6ybXW7FpTKfVK+g7cgl
Fg0Crf1ROZ51v76xefz+b/lzBYS2p75jC8vB6e7HU81XN7Wqg1y/9YPyN0Ln1pkfU7MZSwJtoQxr
Qbir5y7EVM85as1ykVFXb/W8nwijiRjWtaVD45MSFR1RArG+MRJ38jmwtI+XMvaQkIyuSyJlyKRM
JeeX0RSWj70D7FXleRPXj/5QXDEHX/KlUmvziBO8Dm/AAjq1Wq2Ykalok1HNJfRZyWSe+ok+1/b3
KBTeBsicJd1l6SD6YCCMlxp2OGfkQPopevo0yL1C2tmndKrOJ8wBLTHhYgjPFMd644JjDxMAlZs1
iLkJrw4uiGc8jH12RxrfQ4/2guOyPl5cXOaRZsLw61EN7yljAC9dp9HkUnl+3CHluR4YvP6WGUX/
bopLHCO9JNukhxHrbcIKiRh1rUqeOQkzoj0TDyzbz6xuj3RuK1Dvyh+O3FixlHS39XJX2du1pllN
OqIMrzvfVK/gtGcGuNSEnqbZAL7nUyYd2vnjha0weienaOsHmlaREsK++qt1V4iqZ/ZcKPgQMM5X
D6lVWTMbWj33cvakidxsSaMlKayyu8i7aWCTFlcCFJfDm+vE898/eYfs0ubbz1vL2PWFs+lRbU7p
G3VmiRg4MInvSs2mQmfvUFUoxmR4BvwXES2HDu5udi0g9exEGjJb64Gul2Vg9sOfb/fC23tRDf/k
lSktyI5uIiQM5ZMnLjtJA4N5jDTqBGcH9TMFXe0wukLKNjL61XCvKmBVUfaqqsUH3kXT6ah/Htmk
EAeAbJ7H9TL1oe0a8JKxUZfRKPjGOZT1lvJ6P62t0q7aaQDegxjQcVASrSTLC5u59qMLT30WfMUn
71Iwmik4hcZ4RnMWhcEo1vnXxjoCSh0PBL5ckULvFrST/sBdanHjuJiB8lA4UH1kQOfuyvDXyZqN
SO/AtcJQao7c1092lSAHQcAsIawJYkyy2tzTIKycvI5VdjRWc1WrpivdwajQf/mvoHoIzV9Y4ZE8
0sJW6wnZ8lUTaJ7/gb0DqOw4m7cuNl/Gv6F42GswmeFqmfBtfKgtNcl8bOy4aJcdTNY3JAZkE+Ng
F3BqA+pUMg7dkYMgLFTZmwZbwWGVkIVnZ0va4IJL4jqOabZPYvmfLdr0I3ujXb0Qir8KtBe84wqb
HHXI66d+TsU/XHBwmadBY0f/ia310oDMYnQuuPPmSpC/iRWcERLfwBVedaXGyy1bGSU8f3UoJzwg
od8vrhQfD8YMlKa2FGqvp1SF/QN1DkESCr42cNsRUgml4WTHf/GNFgtTzMsOmYpzjwESUsLFwpq9
ow1ZxWmbRqeamnFXgCm8COGZ1qClXJAIXXal/gz/ko6R+zUCL6CrEtgdOTLwyEK5tJYJuEuFIf6U
WqsaMUM7wQx15ofmuFt3N3P43zq9jWvB00Fs8WbnM2zQ7Nx6YopKAqzY/gCdvZL/1Lr2iCZJtl+0
ktNwM+CkzWwiqksuw+D6BH6sxEEXDUbvvmfMvpex3+N6pbBIWlG8OAGA5Rzmw4WA5kv3Tnc+SqmW
6JaIP1p9knBO8/Er7kcr7dlpTWyqTL7zcYsOTFmDj7IN4npPeZBEDw35Xa8LzlkrIbSy3AwZYOZP
k3kGHlcjpgfnYEE+S5o7GbTugcLVnTBh7LNW/NA9Br6ClfihlWGMgpHFu10bAvdo3chvCiUbPND5
xVMmrWdEwt7gvCS8RIWPDmcT2/rmJd89PsR2rMjEIxCBQw+vQOMD2TRy6w2nMUbUpzIX7O95OS8e
vM7Shms6smUhTLWIZWEv3wyZppRkQngDdcNl+1bZ89DdUynCYwuUDHm/SZ82c85XM1tcS0t0zRAq
7VEb0KFwHIslNQHJ34tViVwdyDFUCdB0IQHZjSp7XFsYewxOLkQfREitN9YV/s63P0Mrq2aUEuL9
ffKq3CL0x/1FVcQ5RkYIPeSMLJBmqMBQpdyg/PM4HWGfhUiCkuRt8M/QabeRg29ABE+FX2Gtzjhs
VYnu70DyUlgeyJr2XhljTuSlgh42H1+BEGAqyxa62LHZrAqgTqyR8pZBGXb28EbqypHyLUcy3r1Q
4Hh3tTwwhCrHcOlefYZhlMO5gqAdL2Kap6jt10+c0DCrGExwGfduBVmcQPT6jHpcxHXa19b6k6u2
OWsxohaotQuTDbjK/+sarUKp4RrYgggFayuXUlixLS5EuF3NwKcs5zWb9qSnLtnTNmJNa6IZMAP0
pDZ3WqHcf8gsDZrot5KsJLTRsl0kpz8wycjd5meDGeBigpJOp33CqJic9LccFfzlRabDK6pwVm/K
PsvgWg52s5lya2BS4qyDmFejMXP17Oz887JolVLNeZHWhPnbOWl4Bh1sfPy+NSm2re0gHnovZH2p
DgDUDTZ9dO0dZ8OtSgl+MDa/OcY8Q+H3g0qN5NHZbZfu4huicEkAjRUf1/akLeJQOptcMs9MxgTk
5bHjlIOiZWkXRJfbyJ3Cn+10trRXMzUdVOtGkyIqn9Sji8xKgltCSwGrKB6WCJfFPIXySf4asVRM
+G5l4GIP12oBABHs7TkP3MMG4vnK30f3fMOGpl2hVLOH1esXkwYtrMmcVe9gUK2hZsxvdX0cziB1
GBg5fMVjbWnKT419kzxbB/UCAwred1ThHY6w2YRHL5LtAwQiQa4lqsa7DZFJu9j/tIi8I4M72/Ut
0kabs4n+c3Fze33cu3A2LOCq2qfydWANSu/msD7EcpU8jkJ7smpfV1eInZwfkqBwhZgwNyp22WDI
KsMclc3h+q41rEYX8ocXiEDURgMq5OKzJKQCjUf8cWJC8YmLJ7nk92C4QhSRjTDMCcvW/JHJuAJ1
VGdhkHQQVrhZ5kZcgrdIhT0jlBjKcgolq3Hto3IPLas6yQD2D/aLJjFZhjdYdU6Fv/DXYCzJp2kn
TDSd2+NXvSO5qRHvCIEORJ1oqfiyNQLxatpGZPYO+W7Asb/3BF22ooAqGSKjQukH2wdjTDahdq6u
hoBHgFMsaR1ER82T3rCffmKfXX4rm1O45glBswS76DlPRQ2CG/brfZyKAknVhGApsPObhXOodzsj
Yc5HIYAY5ekn4EgMLPSZ4C5SOJ0I6y8xu03Yk49yOKiKJ8wNR3/73B+UniKM2rV2ZtDFt3ZJGrlq
0FTmHrrdddKJb9px0bTcfst0LDh5Zt/66hQsWJgt3ycedqGmy/ONPQNQUVpWumZsCkCU/lVnBPhz
U8H3ppC+kfVgFiexIaEfFQ2WJ9XnDXpSguMJND3baBnIBGTK22IQiV4QSYB4u52G8/wZvYGNfpRy
ZWObIJFLLXAgbw+bGCcP+/uvH/VM4mDMXFIyvUZcO5zRjFXt+B/7IdhUtMtC2FVfgC6CqZcgmznC
DBaRXcboSM0LlMFZ2r1waVzZYYmAHe+yf1Hvi4IUPyQ+QOaKq/1E6i0ZFq9u9+ZIM0cnqjS4vIx1
0Y9VZG9e27iVY6GfIVhy4vGxbHAABn4+D8asv53tcn2UiCCwbYsCgP2/KrIZYptmwy3RCK6E8XCF
ywr/+iY1ktT0UjQ+EfAERqcwxSvECCgw+ttm3ClAnVAaCarV4wF3xaGiGDSYbx/Xh3aM3Wg3Bq6G
VLngPLdPm3/lNz119jrnIvbJN5PbEfD4bm9AIzi13ZvJ5P9uhnLWSJ6a9GYxiFeykvojwoYKNSNy
vOQ47aSrmcJUdjrY+29C5KPgl90EZPelH3VNXIS/bywa6a5Ikq0tFpWANOJ+kL6h77T1uszdCz+/
DOCTHvND7J6U2tRodu540WM8MYnYNPIw/qoP0qnywK3Vrcl4sPeSk1T6pqE/tKDwlUmuwSXzZiiC
MfzMYnI1B5PLFCNbfOakZ0FbR4QfiDFKQ46RQZzCP/QrldEB1HWiRI9tBUyEQjMtYP6SQdqbeGQk
5gOcZGWAHMVn3OHU8FVvjKLZFbZMFxDmvVxh7EwKZQhXO/2uEqf+gyicCvM52g6FMgIk4ULxGUXN
0Rxvj6LAUie6I0ZVUgCosbC4mX0kzQPQ1KWAh4nj9IvQnwZ24m8jqQiM1NU+6aKtq0lL/n9GH176
+G81682/CaFw10BQoXhNGjqH4QqQO9BksN5jc2IerldZN4HmNGzn4/QoVAZMLoS9xhmTxNwpx6ml
gy4CZG/A8Lc7p0tl+TCFmeRu9RFHKmB3GsnOi9a3O4dS3mvmgOHlnEYbBygMRLR0ci3GX2ImKggN
vng/e8QfiuL91483B6HJ+8OJAxhTfmxLPbeajQokP1b7sfeGUpysuQz7dgTYng2Qbl/EiFe82zk7
Pexbo/PWfMU/A0XqwTXtQPj1SEtGnskp4WlKC8kpytBFBWJb7tzvaLUmt27T64z1RdIsETPtwz7o
uV8NN758i7sLWyDoMYketU1oTlFY9/CyUBaqQwNXTe5A2eSO502IEmaoRpgCPMkakmncKS9rhD9x
yZ5dwVF3rMY96fvf5qhaKwtbCtl3h+sYOr3h0Rw2nPxfmEraiPCLVx6H+1zqxk76zSitNweYEqmY
pDmV723Nm1Oht3d5QdVuy/c5PQMO3Wl+6w+AtLD8YcHP+xltLSQvPXCUUApFWcxjcGgAFBgOcmP5
3x69aJIvSkRZhIgrKHmXzvT+l1ng+zp69lz4D2vSmUNT12om4oegnC3PmhMxTy0cFLfblxTOOKqV
9Y8G2RRU8GkiKLOwAaBEF6ahkf48hKPkA3JCpoGQXOWV8v0OO5MYQ4sSWsGiIaRQjFx+ng4WlJmW
8dmZ1p1ao2OPv/6IjRQaDUJZqERkzpsbHJAjumFLroRFWA02wRCrJ0hHhKcCGI0C5GXMzXLloAm2
5GbTO8Td8OPYxOYGB2y4ldEyJI4/SnZRpCB5hdJSqTjpxPw1NIDmO69TDAHrseuWjk+h4k7uE5eA
ioXa37Tz3Lqq7z/yS7KbqQOhpNs0S2BKQ9a+YEQS5Em59IstUY4ba5XffWzrPYkE4hGzWR82x7e2
b0CQbIyGC3b2kpSYBa8Ic0LvapoOI9BedvuGo9p9kLbiuZClxCvirl3mooSHuQZQSRz02+EuXJcb
GqD6hQrChTfDc2Rj710rRDO/AhZ+muLEAUoS4vhBZx1hhxepC3Sxgyvzn759E+NNLUzIZASDWEaH
+XSB4pwYu6A6LwvOaDsKspowLLhgC242Se5Qts419RTZ2H+E5WpLmRpZknay5AYYcjtGIUCcLcbI
Bccfdkyh4/ntgARW+ZcpEYkbqlW4itAXY1OD4xiVoEf33BVas4+G8M9VdtYfHPOe2y7YN5p4o3tX
3WzaM4egA3EdMzFWHWkpyeWj78P+Es8WHxvkE5cTYGlVKVX5n7Y500z1Sjso0NxfEBxmp3KZmBp9
r/E6jKsW/qS1t86WbmO0Bu3bUws+9ASRg84qCBe23RYiEfusOAaFIvsRpjwhRGUSbWcbtn0K0D/M
/H4LTQ/oVPKLZw/cEz042/VcEs3B6QVe1KDIVmyTJofaOhnpTHljvQph92La2KvcowLwcGAllFaU
ger8Ekj5ljv3uojbOG00aMNA6wGhxv/+sjwmIVDjl0lNLbYXIqJEp/pTsbEBUGPLHNKIlbdx+qrG
kNs1dWhvu3+DKs6/e+ep3ZBEGlmyjc71yTLV+Q+fKxMQ61aReYFMiRQzsniu61Btg+AdtLE+g8LG
PuGT9PJmgHXj9azZKe852hTdaqwe8PgjccxMPNU0vGny2H7yLvCJBsc3vXXJvt8e5aS9bIdXLs5i
Zy1yfS9eEXdXXCg1NvdiehtZbsqo1lzNmwZTVsloUxuTK2RpVkJUZ3FT0+KSjC6z1GFUdG6gOjxu
iAAgXiVeHlZvQ1Io0oaF62mjZPoJzmbv5zNK0aOsSuajrC9JPvudzgweTQlrCCJzVBq+dWHQiXZn
hLK2Oi4yKageyyfccz7At7vIx/ypAEkAJekoWm76vsgTNv3RPqVsJyKtFfI9z9g6iyc9sxfJv9Pe
2cylcbwQvnsgxABe2tmLfg7NihIOOvHYvtlFP2eEFtRSWdB31QkTnP42A1QM35Pcox3F/t2lCNTU
BxnaI8rT/b6OElbbZl4Kc2+p9kCDwhPwLn0UD8OOfugcV7RBvEBTdSKBJhl72wNhuMhBEFxJARmp
2YL6hMIPFvlVexS5pjW3hQkGRKxmH0FegGNor+EhsVU/H1RNWUj/6ciA2b4c78IQuvHQMVE2r+LJ
id6k5hVbnSrY+cJ2QNfEraJ+sTjtM3EdjNCPFpwD4+6sAvIb4CiEMQRSBLCRU/EpM/PqexY2Ur0s
MmnG6PDNCNbE1tDDS4LwEuHJDLFGlzgApjWyMaQ6yz+Fhm4m0Rxj/n/QgU3jZwu2rcAAXBfHSjPC
SgfggvMSrm/DaAg56tO9/yIdkKjy2YZQ4IWy0OyLN5UhVFiNigp3jCW/nYUQHWFNWu13XHIt9xne
3FQHpxQfeJ0hPlSwQGkTeu2VwOWnCkgR4Vzh9JcOV9FyeRnkGVnPUtr7pVnvyx8DvB9/1qmhvQ9j
v1StLVN7Id+ddVE7bQAlIluXhk3rN1q3HOBybwBKiJpcgqpE4lck5dOIe6/F/sbceHENHXsAgqH0
V2AqBeRDoxVmbNiehDH6qdf1TPfMjs30pUs/aTw7KwMvdTr9ENwzzgquiRjwE6cXlRM9x6W6OttL
CrPy9NUW5jMTu0Y+31HY12vFm9mZW46+RMo5EavQjI9yGOEJgEx5wCuhbrytB7aCBuIldD4PUnsM
KZx9IYFwKdUpVIO32aB+y2I9dAOvJ88ZIMu0we8MVP/SdCLN2EdMS8CRBLupA5kfZ/VOqUjBx52P
VHmVYj2w9r1uHC8D9XyZd9FjVFtyxLtUgHsaP3p61WSanebdWqY8t9IB1+KmQeHiY9nCpQIsY0iU
NY2bL7of65TwjVbvdqsAhUf2SswOQiYpc6cEpKwcADjIHSkqK4ubOMVs4BCGwkU0ifFwfXcHthEn
deN2BnxUcuWkEKRd74aOnb2gkKWAOYGr1HeXMWXDyUHUBUtF90h9zHSMdYrrsZmu/bhHgIQjEavz
qtt8kZQTNkDlzI/Ddnq8qDyaij144cFSTqxJBaf9j/rI0dGNQwbgHLx6JMg4JBntvK+kJa+Zfxtr
LVp6OtwJqkWElxPdI8kaFFBO+bDHiBT/6/XcdConCmnKhNhpg09ORJNSPEZySrefj7LG0YM5eXSL
i+accXoyY0/w+xu4hkFpo8WZ9yCyLKZnI0kK5g5ulg8siJBgl6Hnhm60JlqSoNKifAVrmFlFUio0
HjWEJPqmiAy9tIJMMAbVRt73mnYLO3/b//DZHHfoPaEJ0v8Y7b4Ww3HzC3Ude6J8N7kvgPKpnJak
zfEX6hR5ku3ua1vBkxnZWgQIpoM4G6i00355WPYiwnMROi3Whj2QMmMQKaBmqAFx78Z6g19USuFs
3tI+sEDHPKZy/gobcR8ApWlXgUAlU+VBrc0wiXEHKwe0l11tbX6DXiCgKYxMGbZiO7KpvlvR0Yco
anYR//fL6KpMKRx9o4k9JABJxw14o6W7P065VVZK2F8hhv1ITnVsKmvdIdMycvYGOa39h2HxQHrF
9E0AuIugDX8/5Dh+zm7RM1gEZv1pllEA7Pk1qPdKabzyvJPS746G/xDIfbi27ArXfTatjt7tcK6v
1veMNXlkFzClhxYP975XVQdi4CtYqiRxM/VDerPK9wH18provdttwTbadRfd0fws6fKSo9OoMSZ2
VIqY25Z//wR43UUv/w3fpLTs9D99GxJrnG+VF1vT39HlGabX1PhbHnsDu/0oiH5Lf/xRcw2wQb7n
4RNxIdM2UbSF7YAXiU3FZkkEo/NIAEzMkyrLcJmdAcSlcyLVuTFA4wbCodTt2Q2xS+VW2DmnR9JQ
XIIp1HWzm1l8XKZfzVtInG1qpNQ+0DE0ucJl2WTBKPgLfLi/67lWpBsWbVvGRCZBhJaneaaJCOCJ
VqvqkvKTtjcW1EvH5hGZd5tLX9+JeYH/MxbePRFlVGXM36TslxxcKDGFT2+ImPjjRAMI3dU3Y7Hs
FIRvLLG3cjVK35yCnpI6YTCnUNrKelXapT3MTIxY4WI4/UNQPcwSL0ZtOtTE+JTUYnO5jG/1eBSx
Ycl66hBgg3IpRPheuPoZOFiOjxHAbE17gG2au+mml57h0OCJROVB1np6GFhByms02iHwEP1jAIBw
4g8qvDQ/wnlgUfcyJutuCOj/F7gBbDw5MNE2JXWU/zOaENZTjkpttReLHBFZL+3wHsbjCWuwbt7B
b1xUzvKyegzVyHtUl3W+j3kqiJxmP6ZjtmwV0t4dUzyvqeTZj7s1P+QTPZxQAfoVL2O8rEFAs3eW
FUudulSYIG0oso3r+K9dzKvBtGh/RD/dJ8gHf6gs583T4FObUSbT27Z5xHLyfkNbbYFp1Fgvo4Mw
N6D5fUxGjsOoPK198SKuqDynxN9gNUilEmtZau1t8gLW5mA5g0jSyjlFyFzbAd6ILam3+OycQstg
BpsrnDGsI/IiNDn/0L6sYvFfSjdC2WeQMAvaZ1P1IImEV2/RQ7TP9khypHTNpzoecr3o7UegpYiT
UWPmgFHkgAfgRIgpw/mDkijxpdsr9PiOFyGLaPvi2Pv92g+GXy0xSdt+EbN539BvUSgyEpZuc6go
RllXQl44GPda+dMo3Q5gCCtZlBHi2n10EGDYkBpumVOhPLgAzdzMlc8cN44rYlggwBjCyRGykQOP
s7djTG8czPc1EqggOIe5Zn5welnJ0YGujTHJBiPbACQKSxi66pEurRP+il279q5yIEdTmvM9H/8q
0dvzHHdl/7rHgc2RWN8IqoR2DLJWVPiEnN5juHNPvcMwK40WqoEsruRp+UVxHSID4Nqp95PbYcfi
QNaR5B3ylcVSQJDWsfvPVHGokOiwAHwmWyKUGEVWOYcusOZgqWDoH0jMjcc/IpOIb/fmvm5OUQT7
8Pv8c3L7ekb3BPizxmK8ENZghT9P73giEs9ScGUElFGP3H3VwOk85JRqpkf2lzLu0Qh3VjWEOTcS
0uPjvmOihsTFW/Ibvit/IN70fctfHlF3LbMnA2vmnAT7IbxHjwc/F5Ap5le+6XUR+evL1wjCNN7e
vF4aTrGkzRfgJbTT8YpMpmAt4BYjA7Q/K4RZf9M74RwcD/aISy5h+oRJ9WUScnOOCHa4IOWUMsK3
qY/HbaItcTBnjtcorwYp8ACG0tK0hPvl1Fe1/lIVQPB72oYzZHvwjNoHoji7n0SgXqe2VlYFHIYB
GRqNK5vLXBMuz0qkwJXxc0wiPmOJFRA7Foa4/thgp2TB/lNuMoHNrP8T7YwCBOuGNGjGqAoR1ReO
B1oN7862N5iwp0zU6KZq41aUIDA7CkT8RQc+yDnPx7vWjpCpdFvpVDX78biWnesXuo5Y4CZLHDeP
atHpK2oGr0NtNWc1fkg2KpwPu7ETDY7Ykynf91c90y8Z5toLqyzhXhYfZ78IVzcQxtjB2P4ASKj0
df0r+Z7xX18uD5wdziGQxntcfv3cFSIKAUVHLyL36uMkFd3IP7gn1SsVH9SbTEVL/OVAeshumte3
KLU9cHQNN49UcrayfBseweeAzzfLkR9agT2vahCLKm5G+fJfYAOpw1Gcghx8BcH4cbwPivC0aC1b
zHi10ts4sK7GRVNwcOWyHezRUJUFwfJVC232mK3HS/r8YR7TDrbeicH9kru3WqRAvf78bO4moSIM
bnkckJ9oRZoKsYyMQ2npImYRbHR9eZ1LnNxD8t19HGgddAEvDz13kEQORjv6LbmtcrBAq5605uTd
aByP8yJ8+d6PTR2BEgkJUir+wWtZX+xsmWmDD9AyfYUw5AXspgkdJ1U46zkold071qgNgwl8HqmC
ISrD5OTRoxY/U8jKIL/LvoN1pQWqLBeRjycz7KPuzv0seBRDAoKJvQhxrjgqDFo4GpMcFEi9c+Nv
MRrnKyfAl6fiUouXQUJbM78K2uSmK1SFF0I9iDECxUom+WK/JTybxRyBC5iE4Q1wc5DvPguows/D
6a7AW4FCN4+Z9JTqQX6+F5Dye4fPm7OCp1SuKkhk0YkSKUWmJzpKaL2Z9tNRBSv7tPRtfuRiYQbL
b4aJOpz9oqsiqi5L3EIa2MFpb9lHN7x10NZSALYMsPYk3bU8H+7wfSpQgm56n/8bFKKN70sSGTjI
FWWxnW9cZJRrdqwdLdl4VOpR7Yb9casnaiXSZPcb2KBGZkoLZw0oRpVEUSaOpjFD+W8osbu7kcyt
dbXUdcFYccelHUNIAFnXjeqSMhuSA+fndYkWi0KD1PwYmWlrr5Ej8pRtBqTBkpqlE7JlGFVTetll
4Qo443nyJHhwRogTPsLF0pFLG6wIaI5QFCTuphZJlSI9KkWuDIYRc2j1JPlsMqwiVBkTj2TOqfKB
Nxp8vX93N95sRYp/otxVMT2n50tWXrTg/W/LVUTR/RpN8HAWX804Bttz6QRMePvR4N+ofXZ2MftM
sMmORIHGw8z4mt5IulG5r7/5Idczp2XYaCGtvgg5bISR2Fs4djANaIqEisBfd6wJJu6n+B65394U
Qt5R5HyJp+R7POt+0EkrO1wzA0RIAi+QmFvnL7cpOoBCESR42ZJKsTCIFRKM13YEhCfDlKCWKjTx
0NdH/3w+O65wIW59UNY2MWY/VpRMgmrSIQYk14H9a+w86kwsg01L6SdyHagKwM7jD7nDpGe4SA1+
xgvr9hJBrColxZVR/1JVlkByC8oLU9cqZcjqR4YdpF2C6pfiLbG3BQe1eRrXJLNyCvo6Q16LVNpa
rQb0bHegihlC/TtgL2gSijzmw3VfcIIKZ/8GRGI3XsaKQjYNcCbv6hWRmAq8n+3ieFD1rKJMXH/B
hrNDUrOy/4FDMWu88HHwRaXjzHtEnX0kvRC2iJofk0cnQ7aXnG03qqvRTYAyv7msWOV7VQdfHHzP
08gWKiulQdbyBAso+zGsIZU8w5vxahoouiHLYgznZLWuZWRwbh54S+Twf3y/I5S5mjjoO4U/Fv3I
pv50h61EBCgHoh4/lzed8+qTiZXTVad1TbQkwRz4VaSlS2paVTA3KoLpkNf6lKHRMFZEuTUrAz9b
Ka4rSCppYVooY0P96Cv4NncgCtu9iDnOMvzDNQPRQAO1Wntviu21Y4hx5q7XtOsTyMONWVoIJr9i
H8CDepkyztGKF31LaX7RCW8/3fAWBQxUlOn7G0LNmHZTOqgAtCCdWIoexCIN9rM6GV7aFNRoJbvD
DF5fLKmk2o4qOLi05S7lWw+zboQ4z4xBfdk4v/ZDPHXZzIFejOo2FnvsfYlcDJPHSYXuIpprGoVB
1l2sMF9KCyysHu4sU5Hm5dGB/xDLcyytCI+zSsOpqHdBRbfHJ7X16RofhEmzsLmSYwR1esWSO012
7S0BvNsxHDgW57xxwDWS7MypjSwpjveNa++93VVXXsAFTxwWaL+aVcNB8t1saPOORWv2k2R7JFcs
FVO0TbrofNAs+oBnZMnLKfHJf03DsenAi6m0XF/BGOIUSma9exNVNQyIMn5/vkB8+6Rh3RCgnxv6
G/4iy7l6oXeboUs6p9XtA7gb4vPruUOo37LxGAU4c379rT2mIC2937lXEdjHQ0fMT5IT2YC1YajP
41ZIEeMATsE3RC0Gl5a81kAeUGDbzjwKxRBQIzmP0+gu6G/rzUVhhcKTW0B/PSgm+ymnoagMFv0f
w9MizZFLJ7RLlwydDlW+AZGahjBoDxyOizWuzyiSsmp6TkRQNw21DKaIRqbRsJ4baM/uAu/DXO3k
3SLo7tnV4yRMrj2zwo+32C0wsA2SVSKdJSc8PdVH1TS7ZxgoVW9MJ0jO9Temq4b18FlHXG7hOdZF
4YER66C1G+Q2lLU/J1S+EtsAH4Wcdl9bhoEEbIVP46ZCMnCy7N/vIsAeLlCuGufWlaemk+4tiFko
DBGs1r57mr4/paYegnkKB2vpA4b+xbatrmPrGNsPHtMmPWesLUjp0S+satyL7/3gUC2wl+GM1Oxk
vA+MUYaN/4yRPlvPi6Lk4bqV+5BGNDO7AJSDPxA++eACitpzqdgwKkEsylIdg8FtM35b3Z6zCVH5
qQagXBrziFLV9WrAV9OXCWb17OvlIVIShVP5M2KIBPP7ZJ5khh5VYxP/7ncj34Kaf16A1UfOsArL
BjymTQXcV7wyLnHG2ZY39CZp2EjEPyNwdxIFFttLQM86hqK9bm5ptYnCaS0keSoQx6e+5JLE7AUc
03cTZwhv4uyRz8Ex0m4vs6iPix60STK5YqlfOaYW+eVz6nA8+N82wCoANZco9l/ERdfYQqeiCVpW
szFZkhmpOY8kbe1tD3XIf3+c52UcaZ/aHERWxIVSgx6wyk4qDkVUohHRF0GkASVW28Yjxp4RWIF1
Wg2HqR5zGs7HXjBomkcyp+aB6go+nwl5LD1UJtWkxyQaddnCGbkJLWfaggj+qKDpeYGtDBBHshwC
/OiiJBYP370pud//ypyz0XOhacwPbsroPyuKrqijpU6cw7kYml6VTR7tsHL1mHSsnRi/q3zGsM0+
oXeuX2jhrmvbOvRywtxZhph3M0V3altAt+hdFIr/VdvHFwoz8cAP65y9GH0U0ziBwjc9sIg8yzas
yGp0vC80E+D9i/4t+6aEAgJ1xNbW/Q34DOHsdGPqeB8tKE9ujvsDb3+BZCBrA+4NUbd3pF2G7E7q
VvZMtQR5NocFM9fgZpdfQhLi9XYpNCeppZQCLCjMIDl9ISkcGha9tFr2aYCQvg1IhMIpHjQyFo3f
QhRwSP+Pldiw4spfB5hEFup9fYKzufq6YhFafJdn4ULfQ+mI5wvYiP09CUYjht5LoP/fZ9ArcaUi
K96dGT4KCxZAGtMYfeU09hg5V9l9IQTjlG3+K90j9C/TFfR2i3WMoZEXx2NZWE0YFwL6vSzwbIex
s2aWyxUJnZ6mxNjtVhb4nU2tuHOUNGY72cq9ELUvZssrp5gj1WOamnLFzpZi2oHImmPtojETzS2x
tpu8fdn3QBhpySsTAh5sVjdXDFCFfQBgLxw2nw2q1YEAoBULfXHGODhd6YNrMPA1lI+8hJMojlTl
1VJi26W1xGaS9gqwKcv/QdBFLffYKEok7r/C17HhenXNIYbkDFz5j03m7b6trdpeW4kwVhIgLcOH
LgAF7pPvB87ABw8SsS2BxvSOIwAIPK9bMfxCtFxwFuoepPkbNADslIda32ar0bk/qDDLfr4HWgcJ
MPc1Diq/YamhM7CF0q4LyiGb38zKYOFJx3nUmcDWbn9o/RvsJpJiCtVYd1AvLXDdWnSIlSozVdiz
tTU2f2rIxgpRTAwGyCUy8e7y9KmuBmuxuKYOop2Nido2iW614O3gzvOTqSggE00zPXri01cCfLy1
cYSHZrD78dQFNovWKeAnAa/ODbu4XrZYAVfLkvkncv7p8AvIv3/6SPDlrOoq2c6xiGKpok/b0UXc
sDC/eAfelCutQxtLWeF1MLnEmJO3qT06SJpNnq5gwMrY/4EZT5OrLNkib0xzV9zg5aSz7MomE5hd
KZ1U3Nxmyh5q+qSiGpCYvhD2+Kwm87zSCplvLsEBdL9Q1P5EzDT3E9wAf1KKM7kNiPBbvTtKlrXD
DKDS3EUlidZRZB99daQ/TNUzA0WsjrQHIDi01wpQUjOvJ/tQQpjeQUlLdsnhVTWFLXk8lxhXXYjQ
8y+QHt/qEI+eTW63NsoudsMrsUp0//54IHSa8UsMRCYpPz2wV+flOdkAq4yCn66XwHz4p3cZ3aGa
QbF7EaEasMJqTAMkxCJMt4mCeSjliLV4BwDV6sMqKo9PDha0ZGmEb6kkvCJDYjxShtCzVv35udlv
Hc49CtY7PQMJG8glEkDSUDULU6jSQUjd1sNniDiwkMtqsANyouIao8s7lT6c/9q87Lig4QsCjtw4
Na3kB/7SXWHCOopXVR/g0dCkNUq65F3jk5H1c5cKP/t7EXAHkSWyQRygtOsW4RHmv/VAT6ddqs8+
Lmbrh/mLWbF0HKabCIG00xSc4vAbenppfIboTu+q6WSWDFB2I2MoGOzfK/OnByKV0CL4OOG1itVA
aZZwumkW3uBiVH4yzIH+ctf2IVtgyLgnyyTFlnSs2gIrrHzQnxmUP0Rd04qA24eP4jjVnJGozd3e
I45atGxMWUuuzS6C9oHl7JTnsfdGbcWKOS0j3IWMINpXkCwjnUZH4HtN0OLNxPS4eKjbrSM4dypT
uZWn8LSaDvnVxFDh2HaS111I6WvGu7k+H07A9MP9iJhH1hUvzKV8g5eBC4mXNh0AyMxNlhPUmteg
c+RzLPHR47iIKSStfZ+fCCJZPaeb+YsOJn8W1WDYdyQ+GRFHs+kq8nD9c9r8zy4wG5YDjB6I+Qrk
rU0Za6M8hD5oeS1A+idtP2FkRZ25TJ0yv2tD5CPd3KYjlIVnv0PiIcNu+9bs+R3/oYVBvOxxhcBq
5mOYahLW2tVD46jXlX/4Uy8uBWuKivy2EmlSpozvKo7hmN3t2EX+55IaYINPy4z1yqAoj8oZl4wT
MUlK5jscVkCX2Kq3DbD69bMysO68Q6LAHZLYPU43uXAlD5Wwu0cuHDv1uIRnnDaBR1/54nWz1SSP
3W6pd7J7WpDaUr9KY5g78ALNmELRr95YmqS5ll88NLzu60p9f8ta/BP2si0zPwW1R6TAq2rt4LOk
SYkkluEKW0KFA+OG0+nNNtXfpiijGsusYZHlTO65MGD8RR04Xt+dq6ooh2p0yuouF3hEUhsndxYw
YuSjAtT1gGrrvRA19XBHi8kKs77UOw3jrIGBciEW2wp5I2LVOcrTkxR7SGwFQajr+W2cNOPtfKeO
7mgYQrQfgyyyFN5AfGIVNKZQUpkAC+hCrkpG6KfO9qMSFVTJhhfC32pB5yeSOsrnQoC10kuO1/XJ
EN9PTi4yiNr78O2DsTgpMlvsgBP4g6jFuOPRo0DYhhYzLdW+77jf8lI9+XOCbGEM/GEhyudITpgh
DpuJ3ubhhU178giQfbdXwMnr0AUOHmbkzKTX1a/slkT67KjnvaqRT6ZfyWiO1PVXTJ0DqMVtzydV
1mfu+m5sUZkNLR7tetc3Sgy2kuySoCnm5b19zDmq7EdpE3jMClffsQqokfJVV1hWCeGX3EXyTfDi
7/dtc67NQM3KAmwQXsQTe8HwygqDkTteKZRD4dS0MxrAt7zBJsyF2zI/lm1Ope9kEQaCJnewa+Zk
TIP1yTFSRLgnKuJPNPWIQSAz8F/0qpfN0uLjNORjZhRlVzam+ER/m2FEV68ryhRy7Owmc2HRMmhQ
x8YD13ZDo/5cVpiiexpR92ZTip1+rNknrwIpcX6YQplYsbpMtB5TPiUjDPj7gQLuEbIaCeKrJjIH
gKe4o7oaCscY2zhpuSpXbxffFkvAVh8OyADKUWOqyRHT18fWvEpbCRoCGJrki9uDc9GHBG42vnBJ
o8lCGBBnQdrNyu0LakPPA2OuT77ZsckdTIyYpRF+z2Kj3lI1Q5v5GiHi1/HxjAGAjt8WxybnKMD+
GC1Dr3Dkr/V5O+fdqf6vw3QqpLkDJ43DFSbX4pdvDQ24EDRGOxIB96noCzbGfQGIKG61bhgJLjIK
CVvtdvUKJb/QEkOZ+GlgWJSQEJ4XVVEwt234KPlbYaCssYo0A5Kq5n6PFJZnAvgUUaJUDZ5vmKxC
S4YPQO5uGXsNtjIyLRNwVOTM5SVqOm9NfVG59noRwIv6T8yD6074H/NcOenl/AOPIzVGqUAVJaLC
6blJTaxS8p1Hlzi3HmMgcalArFl5BoBwB7SSTRZ+upPmO9Fchm4TquLI108ZKPK5S0m4KivLDq6l
s2rNZdy9cMoY2T4TiQqbM5bg5zxc9bhNP4RPgWlBAxJeFKYcVS8SW2JowxctDYUmG/ku+aif6pIG
p60sjYrfMOdBym2tdM9UPCWEcbn1UJ2hzx3fVSs5HQxLQA33BIOsh2SyPeC1YnxizPEp0vZL1BfO
sfGnGyGvqi97RT1uycuVHA0S23hrdSBtDqWM27Pl8TElQ+B8kgMIm7Qgb0nQa1m0VNDARPbOk+lk
beAYN1JDnUYTMjh9OYEq7IipbuIeXRH6TwGtNjeldpGQAkK65p2ZPTUwa6ghsgPo3zrkm+xpTQ4i
b+DxUDkOf6zRsTKqiPK6R2F6tJEVEFXXssr4uxFuJ7aUdc15sDzq/LBvT/su4Pa8iPUMuc5JYKxd
RoC/v2eSdiOhGmsoGewKf2QilPqAQ0XXObSAAn8jyoKHY2O2J8StOlopEYJdrEydCmE9TQJYG9Zi
NdlffxN2IjhvULxxvbYkET/5otJfHzR13nssxQwNkapeKY0AbjAu3ROS05l5Y62HZWT1PlzGVu1z
nGejlKWPnNUa3R/ImAsCP1/GFyHckgUdnqxJysMuUq9iCfNPU0GoD7ZSk4JlSJu7/YlhIm5O4WnO
/X+hbhf864DwjvdqzXNJcNVRCnk2mpuG7HOTz5DlcDJBhPFfgv+PpEmmdwOS961F65hjRyYfif0s
JWLmm4Obvc/cszvzEPkiEHeZJpkCrKNGjLpgEraLCEaPsPKXo0bRTeWHHfoSz0R75gW9mHUMDosA
QJc7YUpwlyIBi6kQjMwS3B41BwJd2BOK9LP349AI79wzQwKTM4Lc1y528E/pXvhTQmx+7QBqeEGM
47WhAYwSWCS3hqyKy7/Dq1GaQdLtSUYIBnYtWY2q6ymqTBsIH1ffaj4IvgcFSdenzMvxwviNtrre
yh+Nwrm/hutEiDhDTwUW2pEJ/GE/D841UilkCXiqHyvO9FL4uGYhv5Ef8UCZGY4prjXE/GfWxGeF
tVQm+RpSyLw0ZtC8thSc5atYwCqgQv9znLOPrFztXjuNNT70zZdoT2owa+7DEPGIhvskTEbkbv3v
ZdZ7YAV9wozJIuODxVvQKGiC1SPDVeJ120YRstKl7/4v+b1/2VX5On3K+iMBkJ3HRHpNiwwOvswU
D1PGqzPY7dXbvpLGZiri2exy1o5e0V6xHxRdwyj24Nwlj731pDbiyrHQzqEsivlOogRzWQkIdzGj
pbQgLrQe/mJJ3xF3E98PzcJ3k0FcNfp94a9zupZcJW9MpsubQUFnWnLdVEJtMs1oWc//wOJKFoRe
emQ8BPng4iJ4hnRLOJEGmUlgTkj/fAxyzZFjiOJ1SfHTjoARgxQbH1p9fqYtcx+owdZTZuyJ+Nby
rTp0frbCWO9IpQCX6WizvPqkzCP5HTTjgYT7ZgbB2vZxdLYaan4zqb/5MkZh6TmeIKo2nF2NfJ6S
VkXcgZ1/uYj/wh5LbuoOpJyHaEfDCASFu8V03QjNY6U/n10qVxOM3L725Pmpf/ZAhSxNbBrHkUGU
FVkmPAggO0CUbei5q6QndRmkRlPz9FtA4nwLhXvko/2lLtAbEIZJQsfKd5KPvRvEJP7WfRZGf2wA
NxQQ7TFZhhijWXBb9/V3jVrr//OKGhvnu1Ct63MbI8CXeXF1DpB9ktb8+qP2Cbbkxqgb9A1FWPui
/iFAZyMW/WXl55HSpDz2dafNPEdmDm1OAe468Ja9UBDspam6ROVEXojDyvE+E53RL0o02PmfQxmA
TM+mUNHTikTA0S+Ee/xLjva8sMuZ7RroGhc8oeLFXERyLx7jjNq4x4pqriBY3iVU39CMmcyKlllI
WXW+3eWzdPVa9CZY4IOt9G4VsUruiKvG2I4dmhaGKpwNJ9Yd6i+vymxNHXRS88C1JQIoCLUFUdjx
PDP4Vn+kx/Jdvol4QrVWtMSnYfag/WAPfAeFGpLU6S4WwmG+d68+jQw8eJjnB0P9GeOO1p0sWyp+
XUow86UZxxYtENuyBJAsmT+WS1rG5uIFQcYFuec2GeSIjg87wJiB0v+mdE4pLkynQ/lKwAZd3DE3
2nZt3P7+yMMoZuq6EQPm3uH6/fjXZBTXQD0g6CR8CwR5+vKh9yWT94dwPd5s3HPYan1pVFoIP++J
48MfMo7h/uF0mCE5D2ZaE9Z1/z8ZdpY6pIqdQ30dNcrBABxt6HwUzCVqlOAthVvHXo+byJPfQp1Y
hDvk+jRWb8Xa6dNrsPvL9dKw/Dx7CMBaBK7XpcqdoXBPqSfP/YUXjofeiQ2sr+srsPcAXMbgKxzy
WR9A/PZtjrc28FCkvK86jQCVGP7PKKnSlOjFQDnN2RofjB8GNoXRDKeSFLxyAFpNhCss3EAbBHn5
Z84WMGN7JRAJgw375NELYwSPD7c7Rqrb/lNLbZrV+l+Int/aruYwR8knb/0BA9ak6ZLoEgGuXH0E
DDREKJBIDJixxhsqIq4INhf6P/lPs6oqsQULPCCX8CgcvWQBN2yH7XjCCpgbmBbkzdukuekV36li
6xo6EgIy0ecKjqApphgwIVjm7we9CQjTT9W5btC41WMl5CVafxFi1Qre9j8qpW3P+fjxAhAG9YoF
A33tgvl+ylt6dbs9+y7Fc9SDmeX7wBXlWf69kMjfsGgjVWfC7p8Zc7/o/rm+qCcSNcIHU67F8qaa
rCgWDhPVp7Dt9UUG3HCh6SDFhSOl+VIZJ4PFAlOp1I21XqOrU4x17RLf/sLpTBbqUwewr5snx96e
q155LrCfzFj945v8vDNd0OHUaNvHiMiDp0+b+0LRhQNBV+AZigTVRitLv7r8jfzAgU9Msl3O9XD2
8GC8f5Q2leJ1vA5MjqgoWx2kI+OWuMLIUyxxLy4PGWwXrFi858ygtSaeElPXCO5MKmQOpve/nRpZ
x+ZESeJzpskc0UhF3+4g5EG1/V8s6KCpqNyuxm7hG5BTCkqY2lk3CnUN5R3KHG0805sfTHuwDiKK
geudGtuQ+334kaacABniRGaEspryBiWmLDywNUW9DV0EdhN1tJpECAFin/veccNdqizU255sta7k
8va5FgYPaRgcpPfAPAqMmKwlQUWuXhq5CoXyKk2pSqMnQXqpnZHgvGrpNaVRE5O9VuVcKNLW/aX+
yJSnMgM0BwDt8UBZJRizyveAvM/K17Fpa4ZUd8YDnsQ+OBdHI4EldUWrN7GoJrHkpCDkZ43kh4gm
GgNBgtFyzMrXV8hI0QxMEvPnbJ/IfYiPkij0la+Eo6wKJm8sY715oT5lA71hWkpboiUB7rAO+RqF
JqKu1d5s86ygd9qxfNhNd6V84nEtprkSqtN+vdXPP8AyKWHMIqEKX6mjIDnxCxhEhsbYD9jXxdyL
p6XDXVXrZtw8Vimmg3lUgtZSKNSmq1nJQVBkEvm/yeQhi8u+0vbZvd3vcm0E02G8+mCogkc3jK07
B3LjlDJa6AvUS+I94lDwW05da5dfZGBbuO1VaqQvQLxGlSklLOGHPAEptKzsWAsW30qL7zTz3Bx7
ZNf7+Ha6lGNN9MzR6gZ60c3Yo9p6GBNc1ewCT5YinWigpCr2Y9wkCWilI+maxRCRaRoeIgxRNGkC
SfrmNvFNW/2PCVEWYfFEGEvLZodBQ3aMWM37pd0uBJP+8Adh06L+bVYOGTLpfdbIMPPfMHY75h1n
WGetv+4EdKBa2WqYvJ1x4hXMkjgTpN+J3zW714DcaeNaLqaw4e5BAyk8JT2K99HSAJJl9kByOjUz
50CwBEpCg1jvoYNAD+K7LBdlXSfTM+P2uttMhOifuX4IQLDNeUsg0RkZC0iQ0zUqPu/Jx08O6SLS
/h1k/Q0IpTubOnKnL6CW9UWmMI1M+MoX85AyWQ/BsNSvbqekdjTqJOPJI5za4Zt0cj2m2jigSZ9Y
S6Zd+2nCeA2rtSCZj1YiJC/pcfsC0YfNocMgEB+b1se9s8yDKuGCyTkOwxtIvDOl1S1lgmk/TzIi
2lamdmmgGdATlEASe95/fIkBmRm605yN5AQ0nQS+PByXi3aOsJ4qZkEi/+oEqefuY7h1RrBz9zGZ
CSQJ/eH+lMB9SFHGTqiF/YAwmukNnrIyRJanuLlaCTAG7zY3BZD0vlIUvaP8v6xNmnA5RHOJzvMs
b4SVwsfYfjRF3fwLgLlSbq4xY1bEiBH+k+/KWzvPshw78cYBvH/30hN6ky1yWbnzbSevULiDUwjC
cNIyyPOB1Z9qdUYn9I03/gqBL5jL0qOm3qE1moSBNseL5r6im40TdMPcY2OLoWxe9i7iEYE/P65z
ZQi0whi0g8jEu83is5k5tDQbNLeVB8ZCL9wCv2uYHD23cR36ylp55dSwjnZOdYYQQI+u35z2RIdI
qpX+KXr4IwmxzllihcQKZDXNpW7EXcde7tIrc4pYHhj0W+Jp5/7SdiMyywr4sYAVrSsdtuVwPnAi
eCw8U/f2NUjKf6hVsq3cWSlheFcEONtyjNWQEH9q8JDQc9u3GbfD4NORNyACD9TiLPCrq7lYamAa
gQLQi3ZUpcmqbXvB2h0IufIf0P6wQd2eX8SuqowU3pk7wytUCZrBHGXOD740bS6ZsmuWMeRU+jrV
cRTGECCcogumaj8T2Hq3Yv+01r/ci7FLmkhNEaXMQwPpsonvebusZZhLlHr/i843HUbujYspKFFO
EYpwTdmznZ0leug0sAlQjzcnQSRwuLtKyMU6r1r48hAkKb07pQMUVfI74HEu5BeMxFYF8PQBKhLR
JXGAYT2RI2lP00De/VusBll4JZZoamIkps+dkJEdYXer8VhjfV0Jb2A/08H/8QHPd2lKBZLGnabF
mHF7rP0kdb4f2dLH5M9iyeUE3jdaIPJZZeluGv5kXZskt6dDQKpvhxnry4nWjlAuBMylOvxO5cCZ
bvGaYoJSGt07LQ81kuf/aVePT3ixGkM8H1v4dsoyXF+j3qxTT7zdlO41skx4SJGiMiaRJqjrB3Pf
Qy6PN16SqdilHI1t4GFxS9LLGqNtdYFNdp1k2UNhLaRsC7QdprWcpvT9v41xu2Xh1JCf4CI6bJmh
DU/dw2DdO2ebxUSz1Hj7sl3y5zPvKyesZiclnbFC7GOGPxA5eAmcRhf35De2V4sWQBuZC8Wu6nlz
F/AmkrCXgmGp0tXeiaAoQYjnJVVKxfbySi1UwsdProFePILZXSPkUlxE3Fg9dqfEWBoVsW9CrV8/
FN+dXLqsEFe533r2eN2MfjutEro91WW1OuTk3IYwnM6bBPKIrPe0o7VPgFq/Apv1/fnGBG3f0Z6b
w3UtmcWsEC7fKIHSUnQyzKaQVLIHIIkBgXn4Cmrc+WHrGOj/N4TKJMhpzl0WNSn9EppFsSMPEgU+
9d4LZOA7xynv2T5SObrg0+o+tEU2fKDOTpP0uUwDQfKqhhTobYctmedOzhx5+1VUdWHsKUHptU3d
S+7tKCo9qyjMMbJo7amL0fUnmP+7IKllbjmwox4niZRRRwNkaOuXONMibw8a/PAFAKbmQEnu/c1W
WIwnNbo74XxPm9tGi4FLYuu+09dg5ghuY+BWaY8AI/K+GLowDJjv4jTlZxGmm/FMxmKrdOobvjuL
CzOb7vM/regiHDeRjuCEpFLeSD7C26XYpZPuqfdH3I+VPiepuIAn9OHpl31qQQ+OxPVPL87hbPjq
NXTCVK+usnfQo2SF2aQcoDmJAOEyp8FlSlC11lSRchEpSZkUFqpnIi56ONL609w4axO0LY7hdzNC
XEOVhTE/+pYPEuSk20pv3y8XtN2TWazcic6ixWxsunT0nCrXP+RaaPgfD9vZmkvb+MWoB1HHsljZ
dYdUzA7mSvgt1/xGzZWpzfP7k445j6o6HFelejsZFEOj2b+G7coQdeZS7EZjJ7RbOqWJvq7QahF6
selTQV/tYxRZdZg/WfukhPKjQymMiiIyY8WgAhPPHteMpcJLMbMQa3KJh2L0A90oougJZ3OGbLwt
q3B0KA9hKN8N+0GvlNrILzyHYVSIwxBlmfN95n3ib0x5AVC7/GFUmt7uT4zf1uZuVaYKk097h5zx
Sg3FCY1FCTgzODTfZIdfy92lcfgASdoXkwQt54/mvecBjo2CXMkDDez/5bbFSzZ0LPmRlDpDYiOZ
Z/80Yz5JMFEx5sbSLCkn1dqxZcbBvlMqe34N9LC7uuGc7izISb5IQuzIOgcGvHKLdRAAOfa1GUkV
qpbY9PsanwKHk9CawmaCUJn0D74Mk+m5AHVbRSgAyIGosu1hxG48x8bafae5pZ5Fhu6DC/RdKPvF
vRqqtBUi/6JaZst8/T5Q8pv2TvwI9AL3diEBt/6HvfL/8AsB68Mqd5PKvbv3RzEtGI0rj4kTwxDT
iG1YdESiNEGOME75b5zeu1r+XIUfwY9xwDZ8+swwwMM1vSnOd8jKgMjo+y24PzjxPuKYdpqWHrmK
6Q0wTT3LavYn0x5DAnP3DR3TXW7tbI0aYxEAYihaaGXa6g/sBUJ/Cac1dUBoWCZOfoBPOOeKv3Vf
GdhrcHB+fdIGGor+/34XHj7gYnoE2WZIp0ik+bryI/PfleIpymriyyEhkSzO3gqQkdwin8ZURA4V
8JeuMDVTTvPpfW6guskxSH32+zsReqwbuP2+vpKYGvVwRR4s7KEUzEL5kJiGR+Scs3fABTiRovu3
2Ja1LlSQDFZ1VcfWWvjZ374T0JxQ9UaelQrY/o6zsP2FozcCrN+IMMNHcmOUEn0hG0kg3BXF67rm
gWRsQ2g8SjG226LCahfJNhRKYTAv6WmLct8gu7Uhh8MBNCIQEA6tcix2tJ341GdcXFUMv6jUN02k
bwdnUBKwggNovkbFG4FudWe6oiVXSwAK68WnzHX1sKjtfzoxjgeZSp7RDv0PwXj/LV9lQ1ctBEyy
s/u5Nz+o0NVuyAoaFMK21mL6l4T+Gz+I1JsAWGalMbeLMjRL68PKVKybwVW/bLjOuxBf3Vc4SmXs
HzsMoCVsdqSG45Gu0+5ObGC+GB3mm83BPXEpeHZlxFHsyemOBnNaAdRDQgJxVWiyDRxuuITxNJtS
GtS8rkTtu5IjRxtw1vqSCa1ZbBzdoNgRHutb4KCNqTlJxjXTFtt+jqQZ8iJ/zw8mP5IwrZEL/syG
AR1nCYFgIyqbqI8T4mmY+zzDmon0n1Tj1HKfM4bbpWGqJiLfzIjjZbpml+sazWnNM+pc4q012ds2
9J7fRX73g9ajKXVxctboSrFjta95XZg1HElxztvLKIJoif/XYUV/wZftbPKMzJU+YSruj2fR7sad
YH4UEP+3Z4kXXVmxPHszeek+GeK4fgA0A1KYaSLVYQJSljvnka4ngee+QQXkG+JODAwtJtiubHCp
J2v05e9eXmBMasFM1lqzcuTNFQOlg6YK0Qm8nUTLqMOwQi/PIv54voP9PIbROsXWs3cN2nCzvBK6
pfbC7Sah0wqkPD9fbc00O/0/i3gYill922CIt4bRYkVV9kMnpKWDHLOLLMaXLdVIby41LNLVIDBr
kCvFutJQpwSWrHR5mtkXkbGvqZecues8fNVoxKlLxku08GQ2heXoYXtBrMN6w7MC7v2zyOUBtbtq
kQjRWFUANHkWAmUd8P4DU+GyMWr0cJH6Oj1rIpVfmoJgUyZAF1BZqpHeJlSuLs5pkNyoY3J4qtbH
8Bl7Orot7Cb+w7KNWX/EiEwl52JZCqrMXEk6Zfof2D4SxpNpbhSQnJcvE03435ZwuOE3aAaQXyiT
HlL4CSxeSTcAp1VzVT/7umgkMqiFhHMGbCyL0hEzkWNzeoFx9VMoq4tuGk6qSOpE6HUeyukeRHmQ
ZkEPEPsx9Kqfoos/9sQ56Cyj0mi2u2367yKftP9iuRAA/dwj2YjCp1f3F1w6FbEFpnrL94zx/gl9
4g15+e793DSINVnTbRQyEIpUOOBBbsYS7G0ziXFhfstQc+yNYoZhuBIsq5HbmdRd0BeP5dvbtNzL
8wJbMEJkiPDQCeJy8KSzAtyJJXWziAVCO08KCLoHYqauaX+i85sLIoRVAzCJwrknceB6iLrUDvN/
81D7a9udBBC4cntLqVqofYzLvgxgCCcaiteNUtsitF8QmJbeKF62zhSwBbjIR3Mi0sgtfmY1Fxta
rnn1RZKMV+rlcxNKzVWY8Te0MO8nya5knfb7b+XkGH/CIlPCuvrRhPFEFsayFWFUDcIvUSip5e92
J5AmsoJNfIOvvyky/pvbvueK7DQFergoK2i3wKnhETOQaJyHvqtO4QP3J9Sj5b36b71/0GaD8Aiz
Q2KvK80fziKvr3f5ezgQkp3yRCmL9UUUFby2bTg5rR2GrS0N3HaIgeJQMD3kwz4ESuYxpgcToEq+
m4Kc80pEbT5ewZA5TMuKJb80Bv6bm+0F+2Ap++6FSaYgmYmzVZ/zpZ6hEJ54kj6vdnxjWBcs45ye
3eBSjwxAb9O4ApHKwtWXrW8l36TmuCAtNnKhjRkQwyAempjuL7P4+PU6y8uF6C6ik8jhNyV+AIHb
hOQUOw1CjmkD3ZAuoaRIDT49i7+41BBzsU2Pdt1Z3PccO5sDXcB/91bUN5Ng/SUL9/RFpWod3KUl
vfmz5ovX/opN3wb+lYjsM/E7qWy6bH+3YeO/Cb+C7Ito4yg6RkoI/YiISMYc7sWkH6RT3ZWvCarZ
zKguPhfpnJaTlt0FhJlleO8FM+7kWOSAfuygqpaY1HSILShk2pyD7PXerBUayGQc2VOEn4ENjfE0
HQXrKuMplRfF0GvSbz9uxUAZS4M27QJNZjgqvQU+dcjueI82p+7eRIUIPgh6K2uT8YappL5lRkzs
UaNQ3fTs4CnNbA2Flv4pnqVHMuXmCKXcHnYipksfNr3Ww0GIxAJFTGrcT3FsiIKY8BuKGwCA4ZWi
eBgDPK8wU1i3E7caJX06mGQQd0VnfwEYeHfOuSRbm0KS8GrsLIkkedsDcy2MmP4d6lUn/twcuKj6
bFHn71zAnRy3YMTfbGUH5rTR8rDlsqzdIIAd8KfYo+YuM9ja4xHKd9vPcHAAqbE3alEOLXOMrk0j
5h27Vg91n5Ooh4T3IQnlKFqt+xaEamkua7lWu+yTYlGAM5ReF9Q/alYmXZSm5FXWz0jMzc+8fMEV
cSZOJyWcM/ET62ffugIqBWwNo7Mwa4KLg5k58dkosrpPHfHLTWB4ciGcfCXsKBrOzCcyxbN3WRTc
jVCVEnn4Zlz+kpK1Fvcd0+VrMsq3k1a8q/R3CFBf0Q0fycuQKGXzpsPP9COSQrgufCuJ5BxSn9hf
+sBXboPv6tPPJEvhNWLmkmuDTt2yjoNHWijaBeZ1YDFovRhigKIwmFmmC/xju9QVNOT+bphTgHeZ
LltTrmETBNlk7qma5OlAyXFUPvk+Dp3dgEQXOHxM/UgIGiwp/1rvCcDj1zbKe59JAaaXW4NNxqiP
cTnGQINHWIcTl9KdRmGSWuks86ArhH900aFbdOth/2hzRGq8RL4ZerqjLsZtdsgWap+EIawK5Erp
hZTjzds+XWLr4bExvcCzBTzjSk3G8Vu3ChedQC8bXqc+EoWCOXh1n9CaMCHBWkhLuE/aHw4PgpDA
19/StclV850ZWo+Vpo/vn4NNkRgRjuApScGXIkyWBvZK2yG60rNWpoTDQBxO63f9Wn95A+IKthg3
sCgZYmA9MlhfAKIgxwcjcB+3xcn1q3+0lmlxz+3BGXUI8TUten+8udNnXTfOdTeTqHclxqhop/u3
Cnr3UhZAm6FpPlhEFi8eG+509yoaxcDoMr1wijSXXD9qFwCyz98PQ3Vg3ro1jKuKp3QIKeUOZdgu
6rqMlowk9WbKrr/6wAHK1kt/Z3+6RWjWZJp4jJvtJkACP5bhIHon8yjBTNGL0haqleqzmB2coYJy
rx5zvU7W7o5LV33smD6yIpvDdDu6jYiC83EK5s/YlQ/YBdmfx163Thmc+RHrIh3AeDSM7jCh6pgV
m6tjV7IhxWFr6Ab3IxfGgEhBx54M1F2SfqY8vRD7YnUfP8bsdE5al5OgpUgNXoz1OgQhnrF7U/A0
21qaffI8wdf45klXXAC+yzVjDrSTHYzLU4h6kqlQgJuqzFgFYAJ5NN4pGqcaDCS2JAt1Vp30tO4h
0JkX2/kLX+MZ2DjChFezvLWZpRXarITCYnbmOzEDccXesiu2kcfBNEgXIyqzCFogosVn4bXrljE8
vETZvvPiUmmtdSVXv+CQK13mp+5yQUI9iOMkJ7TBDIvRDP1ntBXaYh3SJ/zEFD+q3PbeK7k8dmz2
zsg+FyQy5lW3SzXnntPhZ/Tmm9QEnsVoL436tTYmPoh1rg+5ftKQh7PEpcJJqWLdibAvSfeOjdJl
oqMs++3T8tdWZKnc3en3lrWJG24gJJLrU455aAX09Kwep7ESQGASU1KE+57BxDyTjPaIVXJmuVv7
iFWfeY/eeCahw5CgOvpQJscOoFMjTxhnr29yJrYkw3R8d1+vP7brsOf6v6hnytPzKukCje0/CxMc
KIYDCiC+H6kOKf1wDfLZ8jxketoysapjkRfYGvlk5ck8b1fzhZMXfVKrJuDELAr9nVDRkxMwLqAH
KVeLUTVeNOllj3iQNxH0uAftDogClXl/EaISrswpPLZNylpMF+OVvZE8yqapG9oIWY+nt69fHrmA
b181I+S7qRteMmltbi2Heqmk/+G4zn87ooXqIQUeJZ/LyCOv6jSdUMNB8oo3jlijxfb5vFM2tpph
BVIJHuYO7K1wNQd4MC2ukkR3vhdKBiqlwnezXKIXaPsCFrXDirQQWUkJi4ejEA9uSVZBT7dSn1lE
zHDakLuFBegZJW4QqqGV9ri+stfezE9dkFfIsXjop12AcSsMy2pRmxAw7M8YyC70ShQ3eful/v8N
OQVrQniG20uFJNtzP9czsKMJQU1WfkViSz5mQ434FdzWqXbmQkW8XzGeGA8znNqCyyDYQa7YUXQ+
GkfhXOzTAMGJRpEycLwe7QXchmrZHY/hWw60JH/WEwcgk2r5I4qSna3cReWcpfOPXIE8eJAbwEAA
iWUqxse0y91GN1ltA39HedMUiv9cyH8ezeMp0Hl4TZAKQkiVlMQ9KuzA82vjXYSiYT3TOMQZVE7y
BP/cQC3QvUo8Q8Uw00gDHFl6nOLWeROuLN48V0RRVVDNQDHondNavD+sJcEseRgATtFecMyTq1ej
S9+uafwnblOC2hiVDb/x1tWxYjwgnzIfJuVOMV5RfyleSiVi98MdsTyBT5vAXGTBxrqq2+N7udSR
sua58wOp49LI/nscz/mZG4X9e5+D2inPt3IWej+HvTdz6M2RnQ+iGMk78pmJW1A2SKrxVqMHooBU
PEXYHgfLba/2iZEzdv8dh25RHrkp/agYDeyn/1SWjyEHHjqxbOqZpSsiD+z22Ub+XIfIMoufkxAk
JB0BSG6EaMb0rrrqNMRq3M+frpk+VLCBxtQNUEFZZZaKpfgFkmk3EqnhIXozjdZwPhItweoKcmRb
9sOvWiTbzqNfXCbc79jyv5VlxZ6H4306IaIM2dim9gePtcUNm6yxYK3V3OvXqSBFL2CC6rhLKmPm
iDz6ggN8afFbWYR2eL7TPWtL1jQsKdnA8sqKZ8iOQyKOZwtS6sJfxgGu5arZ9mkDvZB4QxXeYz5G
A2YbTByqSpYDlsHaBo6IMh5QIWQz4duEAIvaA+fgxXN/4+hOyCojtaNwIeOAiGKEjkRkBlG7g5rR
3HEKloWdEXMGX9rZFOGZvt32/1OEAlcdhJbx6srgAUM+mdrYA9tqhwK92Y4960pfQYhbi4yGq/+E
cqszAX9JvPkmPkRmo02HySRR8ZqDVV9mx9ZQa4SGdvhpbydw0iSXXcKWPQo8wXTD3R6vPFqmf4hh
r1P7YqyXQoMIpOl/wjYtmGNeXhfeCl91aYDnp9eOzU33XfsUcRyfDlWkGtDhldipKog9VwlNE48Q
6CeB/muDjqQjGLi73e8S4F38W+ZhHfKbjHYwaA6gKMjGHePkMJkZBbUVMeDU2OckJS09gk02UWkJ
aIeQrsWySC+feQn+ar50VHSwI7I5R8UfBJ7sMdfi7Iym/p8UTATaaHhJkAp/5sdio3+SIbm/E7Lm
eQFau98UrMqfVgaug2nU2X4kcRc9+HklGOstXjr2YiRpVTmb3Q7drDXQo4cvg0aL8Qb3jOtHIoGM
aG2B8GTrpptf9VETq5Te03EUis5xBfoqq8b9rBrPwX0JjEU+1JOk9zxg/6jthlsprPD4b9k+vOkz
GykfTZ7OZPF4jvdxNVNP9Dt0MmTDn5rqgaMVvIFjhtVMdehHViWrmJFPSTMA8DTstah7CrfyDGzQ
MlKJEAs8cUQKfBggcQkUdnl6qWSc9Ayj59JfTWC3skVAaAyLvR4bndL5eMBM+MrG3iO1Q6VnJZle
FrSzdmGcB9QzpVxL/aqFQ439ljl2wXOhU2z2N0HSrne5std4SyqDMDvzPCiYfoXsWaQnHgSwS+vW
82NEvq1LwDVoRQr1VVIQ/LBeDkaiaCxpf4NwDofkgwyveycMEEoRTeXDtzy7p5kwT+LFzteSYcvp
qHuICKkq/Lfvejs7w8ZDxpSkMxqREWbWssbffZj4a8lsnb45E5gwlLZdULPmvCii3DneEbS7dh7G
UnaHzAaMh3jGKNHfhqo8Rb6Y6PN21UuA6aB3F4rF1XSq+Ts1Kiao+F2DppNbv8QXt9apgrkNdCDW
ou/oAWxpnx5x7TN23goT4CMzR+ASOJS+uq2mNyxC3PQ+DZVlt4Dc2pR37YhLwdEioxa8W3iX3bD3
LBUM1emYY78OlrllmzOexy8fQ5FoDWzESmI/AEUqWnFmUH5u2sW7NuF4QIeL42LimzfWyLPxwPxF
Jqm8S/otbrJCuehbXJpWgi2c8fG/Jw7+q5zAQAi9sFSf6cOfFjkk1T4Ge04q6+sDdr9G5IpRL17Z
DHmMtYbExceEbQJVCopSAVr/Jfx6xzgsqraTODEv8TAZIZ4oX3MHTZKTLM5DX4o+kUlUbGMCevD5
PL7CeibNw4qZFDp6UgNsNchPxch10qqAElWWJXI37iay38UjCEnf7K+P67pLiTfzr3sExs9Ayxn8
xADaEYRnr6yjKHVT6md88Ychk2f55KjJp74tUP4aKSz/h0VaEEjZRuZIVboowhg4jDOrtVtOaRXz
s1VmKfgTQ9RrsoreNuIL5GQ/sVAYyeYwPgEUMPReIN5jiKu96xnuez6b3xuej58aVYkknnAapwlP
bNzPBKWivhdv68QDsh0W7SJmcfYVMGIm/oLFZ04A3+p7RxQDm+S9HzqwTliNofinLWx60uLrTz9Q
Bocu88a8Ytf+Uqc96QnTfb5bI+Au1fFRcwLneLHC03BEbv9seZVXt3Y2kRyu5tnfcJSZpBJ1QFIB
oAErvKPuSLrNbFqLAHrG9yuHYrzF1IV0iJEKyQpWuc+nvL9JC/KfjFBIPvKbLJHLBPTeOhYNrQgU
3f5z7mFL+wPdr4h33xPcwhnwd8O2wcIHRjLlngazKyzO3j4NOwFfTZUKHREpcSJKxgvBilHh6jGG
nJ+gwLA2ycPvlT0miUNh805i/qxeC0uF+8mc3+AfxQcdkMulmbrK/xONaCmDetcxYEJPO1dJ0Zqg
sZjW8L4kpkAKoNgo+o6sReJz3sRvCzteONLPKOtEQB1QLIlGRlpdH28MEOZZdMQL8KUC0D1uGqJq
AMTmG7yXq3eN2T1TkUuL+WLs39KhTs3XMuAvWKcgKTFfK/dpi4g03q633XxDCnmAvyFIwGb5O39D
+iHKylz6HRq6Fv9D0h2BOUMM/F4OAh1JDLh8lKsoGgEnqF+iP1jMn1HI5Yk2CUhhf1ND8YAdRgM3
Ks/a8tmfbijHVYRh4plVQ7pyb57AKSJlszWqbpdrMWSKWr/d33ZFkBHcCvCmPsiZJmtwgxYH8bC3
ybtOfDMh7u04FZXX2SrHjbRWPy5j9k+xSy4P/XWlmGOmvR64Yv1UIV4c1tHPPTpcOCNBbvnAOFxa
DyOL5j1aCPcVdgjOcTWSdyROfDRlHwJ9W9YD9MppNk5XwkPc0jk7VQc4U0vBn0yUzfW2D/e2xpiW
xb6/18/CKhZIhGOP0YB3U03+CN/UagfOdCnEaz0txai+3+HFpDc/2DzrjtoFVRCdgQFxDjIIH6PD
WYbqDDIR1LwGrlqqJptbvo2On14uVs2J+932KTknQ6xsbTDEYgk+6sIs9FfTFddjeb+WSBrL8zkn
Ix63233VxKQOO5W4FtjVPqiZpVLnwx+1PY53yyWITuK6XygW/3alJtb0HjIHEu0Br8vTQEzqO1vz
VVpzpDomcFfXLC6OgSAD94FmpzAEJYcTTnEgkFZ7Cr76flUvXTKJEF3QW7vaj90XAmWq4Elqj/oP
8EQQCXSwWs7WuKDkBER8txzFSfOGqyCP4N6w8FtYV5ebOIwa/YPWt9GEXero6dWKyNyN7Npue/BF
+YdHr913BsMhEGpg+GbjSatFc0Zz+DiCVtwZ73+eVRI/JTB66AiBLhosMVBR/yjymOPBvnRZlGnN
Bbx+j7jawgtG/HJqKrmTIpKmMUt1MMhKCTIDOlE9PwYqwNWM77+C+gPgdaLFJJQTtxd/+/WEa+LM
LqrrOH4qI2Q99Pr4jqGjBwwBmgYKIQ2iTbH/lZ4JAnbI+lC0AXrNS9CgK+LcGdVccmpgVFo4m0B6
rThSLBme7uPuJyzAY8sViFWAad5GAqRtSTG7nwKSBLqBDf7pWiO5M3SJ0oThP49o+DemCXOUc93w
VNTf0KfnPinXt+0aSVPLywlqxLBzOTZ4R6HVGQxIKePU4Gzpv8ffjvWfTZ0BGkNB7V3VN9zSS3Qm
mzdt91Kz6thyQzuvPx7NqOKC/oArr13Q+TT5Woh6rozzkRQ8jzO6ybiyTuso7Yz2DTJvyCo7QFYQ
fZ0YBeypuqaYa44QVLDcfl2tNvZnVE/d5ztUsunzwqon2WSXU6SO+R4+z/MQCBSL1/V7KXxR4EGX
/HQao6Il6FyDSe0kUrJmMFkwDdXHpHy+OtnbM+jxdjhQfTd6D2Zo6nUfp767DEHZ99qSqa9uwxfN
n2kw1WVEoh2VUJUjGK/XU4iSi+AQAWUKxkWelMRThOYd4JvZXwRjPdtnOH8ARpL9mrwCPVD5HtNo
3IRaac05K5kfVa295/6fsupE4FvIx0e2meBOBeBNXa2/p9Z8hrbe8N8R/dES5oJmWmuOk4OhfIjC
ALg0Tu4v7SpeiOeb33mGSf/vORTXFg+8vtdedlIY+1giUdz5Qkl33BLxi+dldU02KiTD4sQLZcqC
d0Utl9w9Ij6XvZrx4SyqqssqbNW7MufeIUg/N17gsMGpyjUiJBVB+fBSW2tXfJYc/SIiOX/c+6if
WRLfg/Az13RsaAWsiYqBS9QIGDB0iHZpAsZChMIHJ5QGoFu+W0UQOn2Nl5arkud/8/Qixmvsa1rs
JsoYjlpHkNN9lfkbIWzHpHwEiCEMEfMq17lPfiTxvg6cu3q06QWHakabNkKkBoJOD9hGmfyXe3zq
xisN4gQcsnXOCKqGnrmaZ40sqpQDewRJEwlgOqFfuj1/m8weWv7aR2oH5tLjAQeChcNWryBSvyrV
ZGnJ+XltPt+xa4ba4YVLaj4tAzotdJ/Hqi+nBMqtP4qvpBhF3kVLTXMMNmD21EUApo3r1r7ZG78g
v0tUmSzzM3BpHBD8HzzQxrOp0bJIbJ6goJHJiOmIPd5khm1Lg/3rusFA3pZ1xaar0Hx3s1iAeImi
t/QyNtFMqbyWVSwoAFCe1iJT3BoajCOVNHKa0kJPf8MESYp8k4pi9BVo75DPajEUozgSr0OJRu7s
fwzJzoOrp381NQVZiaWCmwuzHbWpHtTOpTRPizqnbHfldnLdTADK2P/hBOAaw7OuQEMdqjMt+CwT
h14YvAYu64WscO72t/VQR1sEYLOjTI/aN6oS24lmFpEVopkBx3jH4XKp8UJdfRpo2HcpG/CO3pGC
ik/0hcozSq9JN/93C/B3EuNmLn1Vy4DfvfyxeGUCMnjPn/SpvDdiDcszwVfptYlCFJ6n9WM7oZVW
08XKn75r3oqRWHFH0Rx/y79dL2A59BzFnY9Sd6YrsOEurSubEHLseA8XqgCtPVa4nDP84JZHU3gJ
KmKfStxxp0MUD88tkGjXI1GZbmr+JJMIGAQ20ZNvtf3IZV6MDN9RY64bIZyTR7xKV4cvtJ2OEsbP
quK63ihrrdHz9GX/YtGuDKxjgHI8X9nLsdNlN0BXA7PGIiwDoqsCFAz9DvjjYiGpE7B9RGPLIu6w
6b5ZxJsJR/HZ1wsJ1eF9Rb1y6ONpzthjyIMf71B6Fg9cFqPNvj2067yI0PWnmVwxOMdU3knBKhfy
3HUpbOx+nKdAvhIToyCWlyI+tOGMo1yPtzmBtU8cusr7SZBiwqvQKYeXu1Hlyd9aJX+M4oOV8cf0
p4qWrLMLFzhH5EOy5nkLLR6IVCkRK8h/wWR1fky7MxGkPlmxnOEshz/sSdd5Gqtz4J3x3Qo+ihyX
kM25suEXdlcj4VGARyK2tIvlACIpEBo42DdGP2klf8PQdGyS+C4LWI/0g59SDpUZGodTox44xbti
oYuLFOgpzkJ879m1IYCPsqlKVsch6+DdIB7LdV6cJhvYapzyYfSnM8EUGLsjM/pNPx9RrQheBoqB
+1TjXuWPwy5yq+/ranR1SyXF9z0FyMz1UAX72Y/D7vDGdpD2QpLZsyQUij0peTu8lE2dgmHH+jRK
Sgz/4NwRZzfjI+oqHI53FLC1+GJakI9iUxheapmm53RUQUSXZMw47rTRnHRYWl3JXEBuNbVOLJP6
2+qWvuLLL7JsReJVHFoM2lWY65w5EBU3QfyEB+pfB5pXr1t2LXmgS78W+9f9tHYCJZWEd5W4jT24
Mfdi1lp1BOHFYYW+UXim4IraLkYslTwFVULYIMZ989f7gMwJca/Pe7dYI4g7G4T5/DJnfR7veTo7
Ti/eDu38CCTJAUwQfNI1b5Urt2QLrf38Yj5QgsV3aDThbHrgixKqKwAPPLN4JBlUbKjWYld6cV0E
7AXEWPcdMt+L62ToNkO6TpqGrmjfgNivUEgKplxZ6N1DTnVQuicyhYpo/a02kafKcrVVOJ1X8BmU
B7YoruqkYN97i7YQKHfrHa2uE5jypfqJalTAQ5E3X/90QqCauIOpSzy/dvM5Suvx6tHRujqBchWZ
wIwgDDxd5Bkf+thJ/CTWMJ7ndRT1L2KQ2dDVinYdemlF/EtyOtDTRRUcf0YU14Cp6QOCdzx3WZtP
lYfqoSsAQE/0BM8OPAdtLxZ2KBuMwFmC51IuVmKI93ZT5ULcqCP0wcD8tiPQOnAsR00Ag+72KQtR
PU5TKvMFP+ST9vwjcjnlQKpU88w3Trlh7dp5WEhGDc1TAD8nKpbI169mLVZG+iKL5mcZfndPd6CF
VKsTaSUoSbdxthGuky/MtclCfXJJfUxzynt3Mx6R1bRzAz42khYw+bpkNwLaLN7JyylM09nGTJoF
/e7ybSDWqF0VB7yGNP067j0+Rz5CIyY9nUqSd1O1v5TrJ2hWVhshu8on/JWC/J9fhXCyK02S2r8D
P3+2w0+6S14IFTOESu4H4sHMJQ9mQoC4mSwzfR1vdbGAa68fS5ZYcICVv5UZaktix2asLmqJGSjz
AKAWPXWTUlre/fMIfAhPykJtj0YiXKpmMMzoD1qkjFFX3J6pqrtXDuo0WIk4HCBvAbrj47s2selx
ju+z16tyJn76ViUNLgPkk/g3nFWm4Mi0l1+x5Gudm3LFa4MjnVdo+GyWRZW5oqU9lPauI5rQjagT
ip0X/+klks7zvW7fPJjS+rkCKOAh/1BykwXtwzySRHjTSGEnJo0Y5860kk37DLGxhewhbjZfWUOE
kPMPxn1tNqGf0bHzFBYLjbDMp4mQ/ETc91m0IH6yksVB9xG1Fg9Y093O1xr5RU3w2eiFzmguS49q
W//SIW3onipUqTCTQVtPvizNUuNCjbIFyzLxxj6U8KYunTvpc3zCPoP9u5YJFz7+z5tY1upAukJD
049gHVZAyHKT8JV3wtMBlrHCXgfn1XFAvLm+JK/ATA14sTvxD+QZs7Hrp8UqYbUhK699bsoia33n
eK1ryZfeil5T/ObuDOWUxUjlLwrqGdV5gkPeYiZ+WVnJAaakLmsL1FgAF9TT1bxMdy0tiRse4Hap
F4yjRpPPDpEwUlbLT8FJAUUo83+qlFlRsuEZ7rVcPZsdi5yDx3marJOalb2ISxS7cvaa6JVF/Fo1
qhk/lb8VLXP+EfgUQomlj/FUwVj3qDwGSjaYX7I0FK1dJyypdU32/nb3mPPffakj2hLUPS66wD7q
icKY9pnetL8NjqbTwTsQlU5wXm86WQcc0RxthQJGGaxaG5ByIOYnuUxW0FySshEa6A1E3bMkmAAq
rsOdNzD88mq5KqzXLBtf8oS1qlCpI31TPd1UF/I6aeSmsaH0VR0twmzyCfsT3i1sD6crwaa8tWIb
9seqJH1F8pe/CgX4YP4t4rEPlTieQVHlTkPPtUQhuZyx6o84BhLBwPVKi8VtPsMDs0w2Hwfy58Tn
ih1oshjuEUQSIe0HOgfWM8Cc9RYnIvsaU5gUTLbzVOnrImxK/TUsHZzOqfKpxMJHOuP9XRawqZei
x+hPgHwgMSRw0g5wuys0acC1gmeFjHsE51fdSRgMqMiuzCspZMtWP9wwrLo+TmrnVkoQd04GYWgt
4DorxxjYYykjX2L7Rf1kopT8iBtGViXH/+uwiN7wXpkEcVucfvtXLFrfaMhrMnta9WB+orRrKBCy
JMLDpBrLFAzbNjqnSro6gorbLJgfsj0xJSyF4W6xqlwxZPSzxMqzFNtkdI6Wdc4J+mNdQ8Ry+Gap
cX8IiFbFcfzhbakY9WaINyWta6qvB5/qbpcd+1Z93t8Gx3f33BcNM/ncwRKusIwawfJK6SADK5Qq
d5zs2mfy2I+wrkn9+4A89UcjHJSHhY1hjqm20i4/K8IyPUHloLZ6mVCdsxEpsJ6nQQ2aqqosZXvu
dmLdmHBnBLAhWHXLgT+c4NCu/t8BXFX6ZEbdF8PlxoastDJoMwvuInA82IV6pPOLAzcZDpjpsCsX
7P8uyUvR+eU70YSlqyEA78EbmNJoG32iKYWvfLhTFbK0XGIjr19VjtTttLz0capEZ+PpYMtaMpJY
sPb1ilT39fUcftnP6BqMn1NVLUARHV3bBxH0ZQc2jg9/fJCS6AycBHjqIqd3j7LdsXl8r9O9oUGi
Uv3mGcxlxB3YXktZ6Bmmr3qnB1TGNBJVF4OMOdVn+JdlEJe5JSSjwa7SstYcaoNnqqzBEkgLUJc7
hCZwHVI2FbcyTDza0+u//nhJH5TYlLfyPdDXl0hovbda4zr2k3gff3XcP8pjm920Eg/9lRowJLDs
SaBOCOAlZREGIqarKBqFL/fxi/rFWnPAyRPJ0MdNGuXhV9HMqlQvnkS4IKi+xjoe6SCJSbcNzVM7
XSVnvTmoCnsSYnCXVRKjHXq6arhNsuv6O6Cdvkh2dXJzjxYIdT33DXcyPqhxRsqXAFzqJ/o9Fkdu
Y+59piWOHWIRXQNDQiyVvMsEkrg9jqDRBzMgE5FLV4rxFYRhiICjShgIhl1JRpnCzqmnvd50o/Re
ZlOszIihCBwtyFlxKhtSVVfdgnzoRhXDVNaO/CF650zTyiztXB51yKfYgdwPN6rVlksfq0yAkJaT
bCod2ty/MvWhlWjM5UNQsdxC7YbEVwqelGp0OsyEipGXQWfU28QnVgZrMG2ubCDyPm8z3u31Wy8M
hmwkLNrtcB+osqEyoa2sP6i2XfAqqwI+FD3wmS1n7E3V2HuREY9eh00mDKJAIRj/AllQI6tJgjfb
EM3HgqlYLU/u2j0WxuLJTU6/uck4RYnme5+mbLpc/6YkRaEHtdlcGi3OkS07P5Fjn1VjE51oU6lX
1lEU9f579T+fLR07j72YpnNqUSUGwqOkJqTY88/+XpH+XdmVIFCpFWgKlTkCqLyqSLq/aw3A9e7a
ex+knkA4y0zKtpWg4aY9273xPkpoTCj6Byj7tzpNQ5qCzL95PAyAvePcU5uHRYjjH9XBPBE8X84p
8C7Kx5FmpYO3d93Xk2g2+qKa1BESAf47bpZ5vEOSXOAkT1HHgIdagXcGq73GJZICgxS1MhVgsUBh
rJAvXm0NhfBousLzNAbsMm1BGW9s82X3F4edF4sUwXoMh5OmkUGszpx0N/k1GJrPb5tQQ4DD46oq
SzGxiHOLfk0SoyP/IXM8s7B2l8LhVCNxDH32u8Zazp6DNMxR6YYNjh1z5dg0AQWj2wv3kzyPmU+t
OrmZ+b5HA0h0GP9dEmXgB+3V8KvDQKTG3I0J2ByXbs0JK1NrxGAILdz37l4TaAvbqq2g6sbkAOQn
dKrMdUezquQrs3APPWSmQJp7rIa3+M9flTyiW0BAV/LFTfRVuGA7E31NNFlk3UTsVMxadNQ35Bab
HJyY0jArPgLVQ7UoqnQspSRf9oUk8QyDdOsicL+FbiIWehxP3g8ClG8rxbCkYGOBjaatXNSn4FZ8
iLWkcrf/1wc9gZRaDuoW+HGQMpEujvbWYT2d2fcF0OmoFdOE86pTh0erAyc5u8sDWDtIslS2BxVm
Pf1l5j8ArecIzjsWsif1X8QAznKJN8PDmuYlj61F6a3keg+XqnR9+FugalHVqyiIlH95374nirzr
LidsT5lEDv0mzzMHjJAp9yN9nxoH9n025jaZh/ZyKRpvNsoAk6/13T8soDKTDM3gf5bVTAsQr18l
j0cCowEinDzLHOJ25PVYe1NC2jghCNef58Jcf+YaMbooNnmicLkxLCIQKje2TML45kxa2Uvm6ktJ
4HTUK+GDODOOl4Hri9aZImFvhblYDFEhdwj9sF5rYV16rC9VSfTlvZ7QqxkkSYKffyfwzVyMRDr4
5Kw3zc4391R8YmKntbhgNEgTSRyd6aunEBAIjV95YOK8I555Y/Hs1xcgCAjNg6bQxxmvuSo240r5
dz49RqVBZkPxVFLdkyifwD2dMk25YCbqv7HpK55Hzr4tOnc80zQHBFeK2RvLlMiXOztYCX28r76M
9IUL2QD6Z3QdFXeC7Ov1pcNKi2nb3qC6gVROJ4s+ycmgB/sBWQoZqKmfFFzGpiWiNq3w3xY3SGhh
t2NWpZlrWz3FmhgMmzSLVPB9xeCK5JAdqahzBOhXCGd+a4bfn5z2Q2pOBx0dX83tPhyI6k72pLfz
S5yCTaM5QMGZkYNwmsHT9akB0XP5NprUVAO1B2VxCVeGpBtP5on0gEyyTrIqQSlBB3tjOxb5596C
CUuDHG7RBfYBaklElVRuB5epOukTh+2QdRRzYXPUsshtQSt2qJmEypeql+nH9feUe1czoUgq1v6O
e79TMI7/PorRbxkvU8OUOtvLZTh1ZNmoLGyVCfYjJe6waqqPjCM98/pl0Bq7QZJavmJjlSaVIDVx
0qIKZWTB6UYFKqfstfG+Zj/JBklg0SNI3OSNrioZIMQlhJyhXj6fSPnPO66Tp3rjgnUOiR+45x43
cK38mHYm0bcahlbSF8XuwagGzyTs6DrRXnThoWpNBqJxuWIK8ruGgPErt7g+k0Y4Ffit3PWTR7d/
+d5invytPdtehemBYj3pGF2rTZMcv6O2/g9u2HZO4yESdQQc3X7pbA4S2wtMaQZh2Ba92EFWIkl5
MFs0LOt+mm2+l3UKiwNJpbTd7+GNP6qcTf5ca4cDqOMguGpVgqX6ogLrXduWRVfRyZVWPXjxRhkf
kJtbeHMQ3I55hM0z+2ZIJKkat/Id2r5kfiREfXsf8m+Io80ns+77XOjQLpJ+eNSbvZaJ6UTxQfz4
jknIOsgZmpfg6FfmF5gclCIOr2NJIfdKoD5/RXG9PsZ2z37VhQO78/2le9PYo5ieQuDwXvSuPWbR
0ck+wLBWwB+BHWDb94cOAFU0zWZO5GQKm0ixjd2JBdvWvYF/H5MVl0LYh9o5isgJ96gjWAxqPXRl
ychX5F6OxPGqhlsYzV2NP/UkJWFHrz87SquDi8WJvG4f6cLUbRg4D1kdMWdO1YxWVlzv0w/Lxier
vrb+evqw7gHP92FAKu6O4ZaXHJD001KzaqWG5nXYG08GV7mH/8kYwxUPIvHaDQVuh74zYnWXMMVy
M/5l5aU2LNmjysy7ho7ZwVxbKDrOcUpG0gSR3R5KLyh0V2ljNBR0DJb4nVaQUe5vH3tjn9t4MPEr
TAGc3d+MqIax8NHRFbGmBhvVZX5h90zwXDEv7J0mffatGiIn3iR+EACb8WQBpfFP5k/k8l1jhDx8
QbbAFy3b0xOD7oq0we9Mn33ex033s1vjtLDDuemkIgsafU/3uhJh19KX32APKM+aRcNUwxh/MSPn
ZaFX1M6kzq8e1BsqAnCQklS21oqtHkpDgO1g1c2c5ImsDwngapWVI06LhQNMVbWEVk37LsKMPB6x
UkmIdPQIQHbHRBNrDtoAinQp7VKwBFV7x8xpJ/1Iqhfk4r4Poku0jGwRDbbvRcC+jdgNfEyhujPi
n4eednyYd7sZVzu2x6mhHhPp5EfIb9FOawCLNgTrkYh60CKJ68DZ3u+8iszv3xVZR8OA4um3O34p
I56osNjDh603RxW3mYtGOg4HaDI8zRzFB6pgtEGOm2xpnh+Q7VkL2V8RTzF27wHlwJBAT8J3UtoH
YMHQ+xZP2JsReDMuKlGnAIY5EVUpUoZIv8hJrZrfBwnvG/dVwrxOrXUxGNBL9misYt1yhiSktXj5
GRrVI+vlVCkS/ny384aw8GxOMvKopYNN/yaohTTwkxJ8z51FWvYURyVtQCSuhl55+pQVX1yOJVo6
q0q4e0b9po/DCSpjwKrxl8RmStl0FfDJd9+H5v7jMp2alAIiLvQBJKfshz3Aeu833XeK0ew3zCGt
pS+7D+zsGHbJUfp8xvognfdqar9VODn+oV3dpL5kL9adk99cK0rny7ohY0e8Pu2wzmfcFDNDnxI8
1Sjtrx6xVFMjWOnipX5IB384RLrMRaUxPJzt83dVEUNWXVonuSFX/8vRrvc/mj31rYDY7xtm+5ui
MlFtYrGHXVXYNuD8z8UEDPFE7lBX2cCvZxfJ2PHAnE8KX4CSpCViGCxb80PvANsg2fbSF1gep8Ja
YxplNMkyP2KIQguplBYjlR5bp8NApqYnGDuP543P9dgpmBpsj4xy6/JFYyUgnJkp2SPin4k65rFe
iIYqK94ewQUI993hKujtoYIS2+ljo8kY+Df6A0hOm8ys3c64kdSwK+ntcJkI6OK+lUz32N9aDybp
4Zi55cxvE6XBloigjDd2nh3jf9gsVOUEY16LCxKbxcqUv2x47cQhrV7w6PMLk2m5oDcWp0X1k4h7
S2vgU3MnKADvyVC/Ls9ttBjF/V9UqouoI4mQE3oNEv2SM/L+EmtJK2bZ2Dw8TD6OyY/ruTJIzacj
SvbqJelYqLUvvfkq0G8x/LJUkHWVaqXe18Avosbqrsz8e6AqDr/jxd510GdMTM/Yf6BCt056pWyp
MSCWloivzTWjaVR7ZvdXpaQQfusZRRv8gdw1luqcl2c33eiGaz/mNXTF21U/njtbw1BkzFjMp2LZ
zYKvkuKMQ0r4yrkZTGxGXl741Va/j+HHdvWdouN/xg73+Q3M5yDmu/eLySj4C5xBUMLhf/pDoW/d
++OiToTPWDrRBMUzY1YvMEfNuW3FCtevrsncgyo+R5nTlXiD61rEsnitzISOivN0ZEZjQuKxCnbj
7jkjmGRBaGKm5cgWaMwBPsbNXbUjaU0M5e/0Tpc1IAW8xLHCU5AR1zoRtuFPDyTtrJt7aedCfLW5
sm7mOx4sSS8MLInpNnqVSjcllwtqqOmd4rc1+QkTiQ5T7DTYfT9RoBTSGtgR8Rt//mMVbqG2Rfb4
5YOftTimej5r4EShg8W701PBHn3SS+aaqhEDap85goRJY1U5eItOhueBcr9wl3DPzPsAyqUncXR6
E1OWOOPYdItHnT7X0EdmuRyS7IzELmST1oM6ovkVDdZ2ZJ+yd8TD8r/64z3dmnhaOg8GuITqeI6v
SWSNJDvnVBq/qaeMYT/bviP4aC9VIJFnpBnf2wM4meIosFT6tvO2xeiK22mESee+u0vMtIpQ0xYQ
T5tVukmXxh0mZvWenmp1dsJpU/FUgerwPXUb1MmfJSbzqBzK0fUHGzHILnxkysgZPDlUO2ZA9w94
KZrYKt+NcBLPpGWlZZTb0lmlvupTaxB54YkpPa0hYMfO/7reHLmb+PVxQmtX+1Icg8QAtBPEkoOf
CUH2dRcm2baKjlfsPj7LJ/wJq0pw2XfS0xw5W7gPjMxVe7hWz1qoaMlfdrjBYOP2YSiVb4/BFjx7
oQY2OZA7Z9qHuLdZ8U9p02Sjqs3LThbmbjeWcML4XeR2zGIUlk8Cw3Y7vsv3I7OWsuti949rJ401
UrfMxwmHxrNPCywA+/3Kg1Kfc/HuH+Dy+U9+eh8/mLowcHRtAxlIRlGGhnyppq7qWB75xhH85Iku
bM/GfL0p62S+d7ZXeLYj4dbwV1cWoKgdDXwD+q2maUawYtM26kU5R0muipMn/XmPljZwm9iUPS2S
AHsGA7jw32/4gQQkEiO9BlqimoR8mSm78vmfH9/yTK8ga2afvloKDlJIHpXwJpx9v/1LZtg8NgQL
Ddx1+aK4ppBcmpOq49i+2ZwsAe0u4RYV62VowdLP5LMNQuM6yEmk7exf5cMMjEZ+ehJ9lD0nMW9m
KM2HDnrAwSXf9BZQFBQ12lhO9rvLhpAiTno7HofGYusDWyAPHVc+yFF65SqhEEABLbqaJxx+LnsK
PpOQdGXJzg+b37kUmKinHTfBWEDB1zlLq6rErwE30hjtL2Wsp+gOkj1MY4LcVJr7EXn/IQJz0GD9
sz6UwJje9LqSFPruQXfCIK/tiSkjXpbcCMLhvPAw4P32an56Vm+8+7xz2wQi9OUfvO+4JyVWnEzc
R86ssu0LRBKoDw9E2snjFPXkEheOCtRL8//ziyRgIibMJj2pAdxZZVUV+fTy+7+IxKtsdxTvSDVr
1cujBf8uPVxEWpPI+E+kSE+LSgwKt1V03oir5XBWLluJfx4OTqBCW38UML0SB+2VAO/t01lmUN80
M3vxevN8/IROqtFCcJEn9FvY8/Ud2qXQO58KVKicJQfxh8je7db1z7tpsH6kMQnd36yzx2uwVahe
hVCpxWEA8o0dlx5zbcMrL4424pnzA3HkRim9Mt02xaRZI/zkbb3lyRuZZ8O0rm4LM0I537fw0JnD
ohimHYGLZuepUz6RHQpvA9acGqjtPSsnl6295w6hD6y1BxY2y8lLkd2D6SqHnX5nFtPkj36v3Yze
ceCLdFXYKPDKn578aSNAS3BOCSyD4g/l92sQG2oadvroMJVZAPsRdOzynSDrTQqPtlBeuA71t+n9
dI9h7cYRgmefD/kSf0uut8qvat+AeizJX2027xwXMAs547NAVg252j+aLMZpd8ge38JmW9zUzrIq
MXztpUwWgfHo0/GPVnn/Snv0yCg2GgbkVjZA+9RgfOx0xr5Hw4MzotUNtk0xLJtzujodpiOA8A7Z
XCNn66VNx+SSttMyKxWutNlUqUwJNwWjoWpK77ploM+1DKSH/Axzs/MHdvZYX9i4iIGL86TQY+/l
0r1Ut6hyQI4kTUXpzstYPpidrtY/RWMuw17u8I5kWwq9xNOjx2aRp/7ntqPPBl2v+XWhbFOrKQBB
si0fyuBOqqLf2YgvzV9r5OtC4onkNDB4vmOK1onESOaMJwhL+sondh0g7FCUeBiNkhZzbBW8uy2H
zjdz2j5qKeklLFknF/4biNqcYrdioO27ZlB+LHGTWilvSXbWiI1Bhsg3BcV26DMVLDX+fN6MrVxp
vytWYnqok4liAJVEHu9peKeW/I9c15jP0wLbM603hmy/z8IMT4n0Vwr1IfFLPaGrGQYqmSXGFWxR
H+8sKonh8Pwh2u38P0vCyKCNiYKnWn7j5e3ykB7Pss+ZGzLODjPAnEBcN0ZUS6CA1kuPB6q58RFS
2heqrcfjNjpO1uQhhrv396CcOSsomYJjVNu8sg92ao6HykBIjjhNVrY6neWpMmmH5CPTjoYIGKqB
uxdogJwj4ctDGULZhrsKRY13dFW3egwtWheQGPoNazecd05OjtO6EUGGLAEq/YwRoR3TCK74itit
/NiUB1iyOmWZhtq8g9ciZVLnBS2OcXvYGbv9GXqOiBcbuJ0J1tJi912JW1rvIctzBO4LtCFoR7z5
j2EuA4Sl1TS9Qw4ajTCiCtIcSMWVdmzVLX1Br0/WJlC6gLHjVUKr7xDsm78oNqvBn73z0Qq0xk8k
cqC3VjiPpopB0hh1VV1GMZ1srTiCLzCKaR+UMhdrJ5oFwh6fX8c3stAsxnZgUIdqLd/0HVumBsmq
OHlWf62uofmucLUnAZSXjrDZYcy0g9WH6Gk4urS3dzlvca5zfzK5IPvP0ESWGpDEPORIhBBE1i4b
Rc6dOIc1MqOXL1BZZ5dpfLiZIwElKt2a7g3WH6W9OUZX36BO0lPplJ6r3bcSjV1fwu+MqJk4LmJO
pkoEUJnCxNbpQGXXS9KZ3tYjWNLd/7oAFG9P+Grc6OMCQN3X9EJD4L6MXMWui/OnHmaxaMvyEyoX
oK/22Fv2MTsSvvDLbOe5CgDmwrqne+jGjyJFWMxajmUtw092wiPxlPz966h9acGQKYV49vVm2F8n
n5bsqIWaobhgrFi/TxE8aDrDxXYYJW5xComzsn7P+v+fDhx1ycyJDPyZJrtRmOajqy/zCMfhOBHp
WfGGf554JwB5hQmYu7EMejRp/olc2LNr475+r5r7qL9mjxlCwrRhmJvbUAQXbsBsrPlsKgju8wxp
x6AEUrpGJbX6GD6Qkx9qj0wZV6dXGUyaFb7TlU370sQhU5KMujMPtiIRS6FgbLnGJkj4aI8GBvhd
G2dXVZA0Sxikp6G9KhTdQkXt2dUxugYzuP3K7MFlIU5AaX/G2SqK/P6yYk+5168p2hNq3JbWefdA
RgHN9PWboU/MolUm5/Pez8lf/OwX7xvJV/vilDkwiHi/pwtuCcHn0vi+3+95Jiz1nfemlEFkIVss
1eIe/OJAAJq5PZvT/CETuZ0kktgKNlElbuQz5iXsOIVKIX/XKC20n9NKdiz/8LSrspl0aM2hQmIs
ggiAi7y0sbWkGiaI7d30nDxh8huXdC4YnniQYBfAdNDmEi4gYo02rzZdzqYZ/N4GZnHJxPqK7w9u
6eQKp7+KYTpXI/Ulg+T0tJaMMKSVHqlb75sPiySEu/nE2GE+5QNFcmwlLKYKlWukJZWvSQfHETsM
KSVEL6+h4gunXZMvUXVhbk/vO5i7kBV1EQrkdBsxrLQqXhNmTl7bZpbuEVxY9ApNEf6ROftrtspe
vUgOk5FAh6bPzcSTjc4OjjjIOkfjFtzbp+K5rcvwUEIcV7YOeMgY4lizGuHW1peMtRUCuoiog7s6
XBBdGY8MmMmqtLKZsI8OOoc9o7oiRdubNZnArFTYNsZTCKASoaOvO/PojFiDkxtujmWbYR4TCdPY
s8I5ndCxyQIdXr4rnzMaDMlEkevT70sAJqdlQRHYXJZgQ+IMllNgDiowyoz6ZyFMhfY1EWLXEvGr
D4uK502EubLgS8Sr1a7EeasgK9xfZVQH+o7D0l3jqAFVMnzP9msCW0MCntOWK2UlSvpZ6mgbXNT+
ZVD1d7GhJcmpWbfke03XImlHt6Yfrc4yIHHTXsI992jWuvhpQoaOrQCB0IqRCMHH5XuOyuWGnSWu
rAam8yB2e3ASXMN4hr2jZSAmaKi6JSQpRUDoAzMI606/XsTVaAk9K4EFv5vtyGhSYj9chMuqqUlm
+xOTLPxT34DKLygQbd/AEqAyVDRfBNJBdpRvbat8xbpmd8ezdZCUJmhQ+0Qzz9QDlUK7E20ASXWu
GqAgMRhpOfTnpkvXgyOka7X3KakvtxAtrVjQ61lB8EzihsQ3L8/Vj1siGiQJGrxUn5uLNJgO2Boh
mSQIrbcrktujYYST41cBgwK37CFlrLlBFStAepnVinVv451SViva/ZzzjKYl8sNNG4aWlEpjD0qY
Uex0b6jcDWN5GJeGUgdbAGixV0iDlkqtMxHCWCzcYmJ7/sFqPhPyn/sbWp56PjJ+PHWjfAjL4OhY
klpLMdtfj/NhHGWdCUa1iDH87i+uea2XGxR6btfnt4M9sWt7KP1GEsCen9zWrXhP/i/CK+hvf106
ePAGNYlzi6i0CpvenvwSppqFqj1e2xV9qT69xRd78z4btlJbmpy4ys6b62yU1VJV5snYzXs0hIkA
n0ToAVj3BZBA2JAUIw1CphVJRUnnpA9XNQHqeQkAzd6AQRSOegfidLjPnGQDSaNs6fthDhgTBzRR
tMRR48/IGcuA9vs4iZ5x/XFZmMPVXsvS9FKVw/Agkrm28fX9Ruh2FZM13yjOMGmIZmI9RkK7LnrX
O0LhiBHZBiK7mraeccfDlywABAbet1vS2E/jzCzs33g7XawJpTwx+Q8mDgqdiv8tjGOmS+KlkYUA
RY7phrjhgN4nVKALXj0duGBfflGlpIwVmjcb5pujPsllw5wPH5zs/JVcoQCTi34oqcYJ/0pH+6lF
L/9Zj1mRleSlRJBQs05/fMssV7Ratu4Owc914DiBfzn4riub5b/XB3JN+2lj5TFYH3+8xk210dIt
30AezPZW53u2AJHMrAZn18jHC2BouOFnZOVVKG25Y9px3I7bY0l3t9XIrv3t7ebGXraxsEpKt9mX
2JlMOjAMY9R+NW462YEGEAu5KkkJx/nd7tXOy0hRpHiuIJ1S4m7BO0qSVwdPx8/S1Kx9298h86e6
BMKzeyIFDgtJfBrsXVKcUlz3PlHaLQ4Cj7HLICc+aek/Ek5GnnXUJnbtNdM+/tCqEvm4dTlwud+J
ckDq2xT5cfFoIL98VRerlRIw2HL5OeK/LjjyUkc3En5u1EShu3RV1D1dIO6VxjzHeVy9iXg/AjOB
aKXwAwRTJ1j8EqNOXAJFtD9XExhAyO/mMYG3S5fUtkXvE8GrPppGEdmGvj+Cnh1JKrdix8p0CO9v
dKx2+8X27lpcZrNwFprwy02XI6W+x3jveE72osXyy1W0AHtq/ypQ+ltybvsgdjxjc4pMl0i5bvVj
Dh3WQFBRGqulA8OQzdH1L5OYMymq6lKe/+34cRR8Oh8qI7mmqZ9bvj607xLPBGS9/uQg/68YhDcu
NeXKAz4O97yE+n8r5egUBCNuTE1eL2+eeIGHcRmvgS1+ArmZD3fY2fD3NBy63FLIHJi4l9fhqi6U
puC7YxpUnOCvQAaoNSlYTfOY0S7uBh2ZdJewA8MTlfQeps5LL+QGgz132RFEf+Q5n/xUx1s3nI3P
cxX9gd6zPb4Q0XEJ+VgQcGe2r0drDZwFZi2e1PHB+q4cYCwNM1bAcrbWc5XAfrAQ2ROtefFJUMZt
nvd2bu5SPXZ0qQaRxMsN44qbcFYBQcOGCSLyOdpTJp5DKWC5BoIiVf2ObYamYVvr29RXN9s/VIDl
/zjIQFs64THNNCkQKL+RR0+rOilk3mA81b+juwJYU4ChwW4+ZdA6EkxYRLnit+yKVAZH08FEPMN8
SjD+HCyQa8LIzwEHe/4WpmU15nQRXmOvSeLMTCcF3rzDL9Ee7h3xezT340h0WVP1fFqY2oSRLbg/
Yg7j1VmI2VeYbfyJdzc1yavn2cwhxUNiQniOv4ufE0oquxtksMa6fLQCDY8jrZs8wMnDd9Q/EtxW
Tf2khJw1aGAxSXi6AEwO2ujHnqL9rdLZDHXC7kkfd80AUCgyRuL0mEdeD+dN2+5DWfrddTQyIzyv
7ooYLDY8rd5iCww+hnElCLMVFYZI2GVbGce5rLtVJQuNtb5xrn325d6g160dZljSgOmbucEEnT/r
Ss/gq2wr3+pimLRwiFowu6lO8gU8QN4pyFKfTqrytzSd6pldSzDKbk5Psdq4OnXXpoSLKVmol1ut
67ZSpNveYRd/egAqonwOP6i/z/hsV0A8D61PfNIyHwgv+2+Px9WgfI1yoVxFxC/Vi+ihYkw1AcYu
2AklObksfNm6AUbdWnhZvs+fqfa4nm5/TB2zhTmp89UFNa7waCWCveazcvgo19tt5mr1K3du1ZMZ
eXfvowNdOK+Cb4+0sSiuu36el2qgiCad0y4wQJPhG5aiSwyj2+uF67/Q+Cv3+D3mWWURbcbXgUEo
qymj9CEFOvXps/LMNYUjyxUMcGndAWgjIQZfalcEm8snBbxXjuFTB5BoKdv12pgWAmp9nIvPYKH6
7lEl5xg08XaoCnUSqQdRlgzrcQsk5m30ELUwD0YVcKjt854BIcBjOfJhTj54QCoKR0G2QOa4LsO3
SCk41hCaDV6Xk+AYt+YSJWbswlQWjkkVMn9IlP4F6ZFzJz5c1A598TsyD7MDPiay0v1Nednw1lG/
vwHvdpqmEaqq5qufEcR/EtoOE+aG7ftLsBayjPchx4taS045O9zaA8scu0Flm9xHgHhPQMABbWHm
L6DM/WjKJ5VNwYYpXL44Tzfd2bv5eJauiHPgY4kdt2i02WZZGJr4QmD0LArTtHqwyIZ4YPgmM2f3
RrVXrgTv0i/6MVpxdeEd+NOckML5F7WMXLMn+3hUq8XhXLQvZ9BH/OtFhfBFEN9lzH6Lh+pe3lkh
qfc+gQ15yICGVEJvDpC6uXLkAQ+vhZRcg5CbejFypxTeoPKnHtqZNo/m9QwbCj59a58uy2GzGXgG
GAbXU6UERpTq99RNC5gfnxhSLIY2/X7BzirmA1ZP2FZmqBMvjy20BjbN1rfdre7Ttbh34fy21jhU
+7nRcswAAdCYnF+nOqnZgxDRnjYxZCGbwcHFYZdsNFoNp6er5IXmz6YPSbIP0qzqF+zoGtVLEhfO
IE3AjhirryaIg1N86AQpxvK+E48aIEfozfF/8Q4jS2Q3HoOBmh/fp93ipsFQSeltgMis1g1bsuqo
QiWwdzvI7gSRMPMiXis04YlV14nQ97lGIu0OKNGF9IPULQYx+COss4RhnV3oru+DrHtCAnJ+IB8Q
yNiXm0eH7jJM8/CxfDQrKnLULMR/kvyTAswz6MGc3BdEYztuR0UaUHReJDkUaGNBf7NI161h1xd5
JwC5iYi1cDIuGX7fqYULUwyS5Jc6QlMPdzeI/V3XTMpPwmhFOQtO4sOnS8ixLjwIcvN05H0VmTT2
j5eu0KAr3iSnRYi1MYgPP42QgptNf5iKDIC/l0t6I/v0IGp9RjSbdB9AqzrmAwVqH819JwbP6OZV
LZO1GgeEA+t517ViEmwfxzk4vfobwbfzT36NmKmDxEIfB2wpGbb4Nb6W+wizb174JjwjprhgiWsD
Rura9Nz4eQosLPlp1JIv1YFrIKrSutaO0ghiW/9wJzPq5HUJljbPvynw0mSRQI9xfRHcgfPjoqIs
itd1y5tiGRznq8307n1ZWCatC8ODedIG2aRSy7gu5z0FlB0NwzFZR1skBi3O4owjXwxxF6giuti8
79np66oTZp9kDYojcHO6NAYKPFpRYbTdpourDYmDRZjVFVQqciAcfaim/fhpvGe88nGPoqv5lBpS
ARxW/i/+/x81ig7QhnQdgjZX/tO3obBiyXeAkPEPRDardfdaQXX7Naj3/Xj+Jb0Qfbu1uSIRrcaV
SjgisY9BBNYFdmzdGLUvFSxZKDT2Rg58yVyJ/XOyfu3RLVG2Z1eTHCGa6EyakrVjBbB+yOKqKw1l
8eoSGlcv41prb2LsHyvsCfjrBArQ25EZTkHHpXQyaAFHXG64pyddZBoXXZiwhObNvbSGNCbtktr4
ZxLGFy3/vjYwwh6/1AdrAPHKmao0IxrZA46Muf3NRp3r9gidpaCh28bJBs5kIUS8AxFPWHtkXkWi
fJgDIvlgIFMG3RKLR/sxzMt8doqAqY3np3il7vdd2M5Ot6Mo77cFa5AupYoDAzGm3dAFgEZvYClH
A4JzZZlyM7N5I2QfRC+REe3Dr4/qGcK/N8IKFPM+PI5Qagcwj7YpxTWnS1YBX/kqxpbzGSbQsx44
vPpKPx5/t8amXnMEY/Le4p9l9RPo2HHr/NGXlklHiEbZVXO7wja1+hCSu/hNG1xPRvmTEiRXvIOs
BNl9wfmHtcr2b2lKDNbr/z8AJQtqCZKn0lF51Wz9MvfVJiVQSqiYRz0CTly3Dxjls2ynhJzxMq3U
lH3eQxZ8LychtY5WHNoTmUNrdoZNnfkcojwIjxZGWztIHJtpcjdrkOq6Pm5CikIdXWm6diIVFPHa
F7yzYxT9n+xKIy4xqW32otX18aQYGsuPyhFFRk8eI2+a8m0NS3JKCUQ36kMPpofU05jsllKDfbZQ
SW8BJSk1MrCEV6ewcIlGDDkCP0fDmInj46RZ1QDmqu7ySm47Cy337FcypSoe0Z7q/urlzXmFst+U
0CIbjISFJN8WS34SLKnkxTkgP3YZsV+Nf40bBRzytS1fh8rgq0zYUnoC2+bu0pLmgxWDgY0VhhNL
4aA9mO2Oxj/JpxjCIsVevebL4m84TGTnpx50S6N2oY81Ica1PhjIFq6YgIpAuXw9aNEejLwbIqGR
6jV8nr29xm3t20LqMHP100gI4+1y95/AF90FKnlTnYjymxxqptf/+MB5oUuM+hNTVJLRYER+TSFb
cul5n4BlGjIvuCKPBWN46uiXd8NbM+5qAu8Hn+06qoStLtHKrGA2MivId2yRbdiO0h/gHUqvAele
De3Nfdm+mzNIldHQADTwrlbTFNVmHq+kD2obw6eQnA49i/JCrbVSvAkz3rIJSkRcPotB3Z3PXtqf
XdHFNhFWx3krOqtSFoR8xMjAQVxfVESeTtjPPI3f5i+lw/cOpC7FJNHRQLJYvIB3n8K4W/yqSiuG
ZjM8j1IeTxtyXvEbFg7uNo5MPVuH9QsE4Q9cv3PmBxy/Lm65vDiW/urmoxp1IjgwmQy2elbCH8M2
LfFuEVjDLVRoNn9qeD+KnY+GU90kPYaOsgfsYSTycrYjZb1rX6tMKtXM5Afj+OCqwrjEviDtIQY2
qte30qaesWBMuERVEv+n1ffAzdVsdjz9eoC9ubtTAm023BPFSqAm7xp+ZrHrHNWUDlBorMUsuxYr
oeYA9E2Gr20EfE+UGL3B66FixlBcOVXADlRhAc8SQXeDvTuZulyfk51ZiVeUwqvci/+DL9HqTdZW
i/jCckm/ID/AAhJUyiDYAm7g5AsnAf251RQToW9vGcXFIhmGnmgBqIWBzu0WkBtqrKCr8zMBkKZK
MbRBir3LDmnNtB5R+CpMPWjDcp6IJFe0b8Ct4NG6yXzYpTJ82WtH7YxettyWKcDKO2OjrXQGKyNn
OrpQ83ShbeO8E5plzi0CY2VDhqcTicmtpk4Duanf6CWBFPkkCM/hdREWPCSHohOnkDqeEjOCHSgr
yoqEtsBmJno/QlFM8dpgv4e6ty38yHqqP0UB+H7ZqHyVpl5tPst7Uf9SB040CNulJPUmRN5gVdlC
H9gWegG6YdXx/sAOsfk/yPiIhvVJUTEv2i3fiHKuWFg09mmgJJAsV7eXbOX1aPyXGWobSOgrx1u6
DVh46mMDxoqU38j6O3gSOKHwcMvcuaUM1ygnlKPXVcbYdYiiFiadGIt8Xwsx9HLzzPFeO6i1Ju7M
USz30qlxIRQvOuI/JNuQz5Vean3J5J/4QYz2BdXBTkGUoNuKWaklqwlAmTH9aZXCa9pobtu1ZaU9
/FSDst5y+DziWZkRlZCICbuKv0XZRKa9N8iLXa/x0fQBNBB8TfVk7P8ArvP48xw/QH8cAFIl76Q7
1nSeTXOjUp34OBCx9MtA0BXRY5nh6oVJzietIdmQcRp2Xbi1UpgurJ1N/X2OwC96sNubzhuvIKJf
6vMDdn4zPdKxCN6vFL9046OhMdm16ZagXI4QPIoBtLuKgMi04D00AT+w6keCw6gxE9tyrVKSfJDB
AenMO46WluddFtAhmjJqxOwD4qPYcVmaW4HAw8vNK++INvoldypPTEsTY+7v6NYKho5KKPYH3/8k
W7W2taDAMqBgLgCc8wOtq99aGVzzjo59vxuOI/NqHs8+C9Tirf4wUYLYwxCi7dekiuQhLmIN+FzD
ADcPWNWkwBkomO9RH+CYUIf1NkvkQGCYtvUP5unfvrZm+44DA8rZnt4iFy9vIs7T8Elqeo/qbv+I
uAU5sKKcGb4jzKTyD5m6FqfxzIm4pqTMPhXr2r5GXPdwuOhFDumYVCe2uB+M+PpVS9gMN09W/AFg
K+ax6Nq8BSzE7Nc+Kg2kjY8wXk3Yy6Q9jmTpPnxSRzvOGBm6Rb5Bejt21nv0d9p1ewi0WDvcuQkv
RRUSWfzuZ96aReI0wj6gqSotwzpHkLoiR59XoWXKLZVyRcoJTFh9raa1DiZXFR9GBogL6Re2Giud
7ldqwFiH6Oo+J0Zv6od9HBChtzyiAs1Em/hpjcZvJTknhJ9WoFkgRHeM/iM/3IpnfMRVwklE8pOb
XF1UKmNQWGqNAFSjYr7qT+98diHNZgP0D9OSYW/cqLDwrqkDOY4/Zl/oiBitVc/1UEWzBmRpFvnN
/UAjzKHzK71me3Uy8D49QSddX4XSw8/xjAgizVEYufKF6KUF1ZG8a5TdlobG3Y009wyk1mmRhq1e
5lH9IqI1A+On0t7gGlGxqeH6HlBlTMSG0CpGBiYH3x5bdfHo5QjxnIS0DdP40uoK3cnRoLZqwmgJ
+bCHJftCDR+sFnu1pHpw7e8kMmqMb12ILji4dlhfAXAFasvhGyYEWNr4+hSb9O5I/xuRfvjFqja/
kNW17Fh2hw9WpjOgGvwWvKkBs2u4ZUm34R36j5qOX3kpUU6iOSMS3ivtwCJGx7D2uHveURpJpG5G
tWrl5ZNUNkE+4DZAGihqllU88yTj0EhsRYEUVyNKyA9cW/fRCqQ+eWBY3MfyvkhB3aXTZ9QiJGJ/
+t8qgT/Ftptk0iBMN0qge1JdSeU/NR+D9UzVXv0p4afTU0RJscJqCEX3IV/6NA/ByKFArBzxShhU
yniqAcAI3Tmbj9LgbDjL9PpkdxH4JDr/vyL3dAYyq0JNxXO2YXQoMHQGBIwd23qEOw87SGKzdkh+
NyIIEu17b0Z3aspf0lAW3WOYxIkGcZWQCYof8nAFBDpE9AdqM1swgLRDF81H68pcbVDcR6a6jjau
mfPXDORdLg/C9CRYFcHOWPluh4EPfBnMqdcGxOrIDCdpsUCaDNECHrJA09E9eYStv1P/ormC1DzJ
AhTx3vH+LFNGXVJfDU0ObqLhzspOIiyCI5JuE9x9WMORFrpgTbifdCoh9EvUm3SUYsewKaDVJ3Nt
GgqGhNhtpe/1ReC2vAMEAez8HvWaQGZr2N1bkl8R6gdsHeCJ5zIuJz12Qgw/c7KBtXSzl2WmP/q/
SGPlrfZs4yWJTyV/sYbAgnGkNUqu2kaYoEtxFzTAAKNR7t2DwIx8bXH1vQ1JJ787Izflrog/sLHl
WtJXRZ86jZ0eYY7w+M4hkAGXQbMmO0+sSLkSfNm5cn1EBToo9OsfgFTlLOyYISHcg1pTTtWAoGDP
3lKcS+pRZtQc2DDwGzZJTmReK8eQ+xiAk7U0jp9s/bSP7dOB1zVQyN4l5UBNg4Lz+A/rJRAAJgDi
IyByVbtSbOcfW+wSA4181w0VtG+hS5MCzs8S/rO2moH5Txi0AB1dP64Yq8PLwh4sk0OmbX/P0Ute
s1M8eIOyyNz44E4XNJXqsGX4OykJ+C0jOwOwx7R/0BKrJV5IO6ThZ+qAoG1tfqsRVmNF2Wj5IxZi
eS8Nc+KMVt/TgNsAeuAPq3h67nPlZSfKZuZwUQtczeb7BYd6eLY3yH4fSOg0SJZWBNusbf58MQDs
L94keQfMKanQ6KnlnyUfCIP1Ca6Qto9oSlw6AKo91uw/gl6yFjBx/Y17/F61ypq+jm0IzF3Oqcr3
ue7J8SxHhZBovgOvEpBDQuX3sgojitApp4TMc83l9koZkiklPVZsDc2cAJEF9Y7g/T0gWd/gO3xc
yQKaln+l7pjicAi5IyCsRc6AvV8xn2NRzfIuzdVmqVpSw9PInn71IDJo771AJFQQHE0sI/g/1HvH
7tMv+manLtrrc0bNaD8tVoyjIofekmuUbnq6h+xxyI+1qI/j4LASeGEgx+COYPC31Nf1g2pKc6nL
BPuQLiXVIwgSKRi6vzDHgWvbw9OBOFp4HMdAME3cud4Zt6Wa5h2LxBklqVUztyIaXv8yJ7uZcDPY
hqlXpRbUv7is9+WaFSo6T5fs0Zo0qe84HDWlGQjIfJNmEcnRMe1KPQxe/Zgz4soMNy34WJ3B4ys/
oemooTDJrOVyK+QTFLJPNfrSsKEIfCd4TMTFksuMjTVgAiYNciYPnmUqtAKS0h792JCdPrEKSzxv
ktHJKUTdT3timb14+o1Bxm44w1TREOF21bQ4FxE82yZ3thCYf9qqDXnDm+0E4fD1CU21o5zYzT+q
gjzM3Un8lHzBVgTMyjaqv0grHxCUmgMmXOBoPnw3oU2UkYkbRxmiADyau5N+7rD92BJzBTOJk5cN
mRISXcK1jfOutTJJ9gJ54rYzBExPypjUzsDd+LJkn5PEBdTgj4uGxntXwFO6StUl5G+n3UF2kK4b
hENgn3edcBQuZgT6cmB04gRmEGksPb6nNZKFG9HbqKLjRMXk1ETGj4kfN03W+yO+0h9HCQ1IuMgE
5aS7HG8MwwqWS4wbDhQPM0HxyLzlMDmF1eP7FjJcS243kSJcTAvfW7pRmU0jglnks17ZAQ+4FaAC
+zOd3guOWTCAQGjkYhOkCl8FNo+6yyLmqCLndicQ07gBEsqKHhDaQoW3dvnhJGHmwIsbkz1bPvjm
rs7A6AY+5bV4zutwBVuhSt8KiIvt2cMzkN/Fk7EIANwYb9AdOSmO22pVe5B2AAqKjjym+WdYr8JY
yPnaWlXFmJo5XcCwtt5UJAqSxSldF78YEIeMLq9arCBOxS65pkTYCyIOB5mTu174Q8pPwLB+PJ0i
rzjH/Pzfz98kMgyWvnoqQ6kfCa6NE7J4BwktuDavoczC1ehZf2y74m8X7oe2qaIDZjaN6pwaQcBY
fl7r9t2sGxVuLElTSEAfBs8V7X5tV7KDEfwPw7o1GaJZMTY5z0JpD4VeTauGj89bu024mYIMgJFL
76nUx+k2nku4kKAhcIa91KAS/KrEi4vINm8nyRN4IRIb5NCoGZCBg58D2d6IgQFK8WpAU1zKH//v
0GD9mshHlI5nKDdGy6HgvPhbYOEOm6JNFdwp69ZvDe7pyPfm2tO4oJLjm76fnx/6Iy5NkQ9XR5gp
KMADfJwxXlzzg7Al2uUj0qyQTKZQA8zMARiN/VPrSbPJCKXEhLj7xqLa6fz6dxWMpAmy//KMyPGF
SL13ArE/ZhLsqhZ5Xa6/8cjYP7TGZAhJXa/7tLoXoE7dCqdZhMtuHKqzWqJcCbgDqNm6TrHVOYeW
GXcfte9C7GPbgIdivfBJS7t2uy3n4fruNmo6VKaeLcdcZdLq6j2+3IOGdEcMecXwrhk7AdWR2Q6t
R9KJoeyS9HM/SsICIlVl4+q+RxUp8PhhjDLSxzK2FqqK8GKrByQLW8rceL6JGpR9JyxtCsziRXZx
SzRgBlGn9l+tsSDn8Y9SQeMIr5Aj7kmvmKyLNTQ6/JwxnClpX4+pahUCP8SFJjBVUnGbJsBZcwQj
Cid0PdoA+9EeUb7c8jx+QrA5jGhRjY4bXi1mmgBVOjaknLBNc/5vZXV2miMb1B/iSpPhfVyaYz0U
aOuQrTg98FiFMLq6yAW2Q7G6/7GzKn5umwSMBvdBaQC+/nzGKZytZnzfIYyQbxoFml9MARaSmliA
h+bWuZc6ZfdecBNMwRGtxEQAxahzc44qasw8LgQhpjsNt5w5v44trdUrxCfZ78vKjn4kmc67pScv
GD9kWUWQ55YgkjjV6OhvHTJoxPKKLcSQ713TzNWs5iuMjZoceU8FyAdjUpzYrGqBSTNRcQdciLUw
8RMDGmFURYKa1KGJ8luv8e2r9LrwA6YZ7vBbOLdr2wDXRYyHwStDOt0nrhKhSin7vHfq1CU6ZvNC
uKdhD4nHtRFX77K00mQ7ERqY4fOJXa2X1fYBfnPVKwir1wWSU42LFxxE5f30oRRs9sWanm9t890M
CRW3oKV+cNMVNSVaupOfXtTkrWpwdRJkpnFv9yPt4Zj5FiLE+Uwe8ZCV1Tbq/EeixdMq+HPVoy6i
xwg3SVUA/eHdUwrXwcqJPVAT7oWjsyJpzzUM4gcBHWMfi97on0bTy86AoUVP8c4QjQPh3qn5y8E5
/ZAgx/VPX6aiWa7Cf227djiAWkErKpzN/dxGapRo37lDG2hOmsGRQv/dxsM9Ky3dhvm3pjHGqp+t
kRsKxVDIeOI8cHy3lj/uqZKv9Nq68BZr0P8m3mXyb/Aoo2ZWLZQzhZ8VTUP3tXjH6OHMZm/B3ufj
MqFW2mSuD5C3+pRKPtChKVUN0sN2p04ddyoyRa5QVIynm7ZKt8GaK9enOVYth3uRD9mgyKE7v//C
35eofA96UmIGm8oji2Z7csHqhCu3b2kX3Xkx5mpCDBJsa6+HWfZzMKut/+Td0MH9j/EFLy8fOOzH
qKAAo6w//b6R7VejDTeve3fXGVcHiOeKd7MiqhXNGdU+EFMjmLU6bJvddCfo8HuyjditOq/H/gmO
wy2N1e4Z0txjq/D9whz5PIE+kcFeLpjh2ydlKQaeS1sX9wzyyNlcrre6xrshwjbBFgIcNKnXZzqn
wGtYYkMJ4Nn+9031JeSgeCONU40/uMBPs9aGiPCSnt8Qtp9BmTs5UbXtfaZCiFIJlbtb14dQZ10i
IiViF3PnB6nDAwYUpBCW8129G8e768bPLlzyfIw+n3ORW919QW58fGgEwYbTfTwQNix5+X7l6qed
4BD7+t1oSvCmtGQo2OnWJF0/M62GwwthozhmBu42KbcH86g5Y9At+nEcEkdJNY8RhIoulSJOs6ev
4kX6Iz/AXwrx+bkbIPLQQomRp2fOkhNM+EMhJk8o9jnhC60G9rZrn1LMRuTeeJ+HiIPPz1Nmd8k2
1uzOkFkJW1t3RxF+Bn7LTODIMF8Kk4hSlJ0fqh5Y0shjkkGyl7fPSkggsoWzWeFbZgFgiqJEpJPh
Vnn8xA+2tpsPlbVXnMo7dTDXclN+a+FB6SQlRauses5ncDa7d92GHhVWlgG/mpXq63c/mx6EVHHR
9CBLkmkpUgyct8cq+ocpxsLz5Wt+wIlhWjZvATHkvSSYTlvgiiPaIpLHgxsviHhBtAQmkFWD41sM
ty2hHp+8Y2P+01EDW1Oy4xrjseftR6ohrxpBeqVtu0T1uPEOxKIpjFOy8zutkprqsJvDp3LLdw3N
C7LrC34Y7Yzsx6jRR+9ftfMKUob0GFDESGui2q1lUmvuywmAqe6U2zBdoTzjZSs2Ev7/WazsDrKp
gVwPmlhx1M8nldhLq71o+1F2Hlp+eBItOPsNVaSIbRbWmPhYpzc5HhJiJqNx434ENQ7o9ahkcoAT
NmActdbvd5jabLI+ifAklGijOKkoY6dtk2ZBfBmN5SCucs5vbqTLqIja7JO1M2GSa+ncNPRfOkuy
rAKxDPrxW3BJQbNi9XApGIvgzURRFNSjVW3smyNHvuKf+83bFz1nLQ8q/yuj9D4TVZVi5cOzD2rT
JEx2RJrafr4b9UYXDq6tTd7VPH914CULA0PcqR7HyU9xerH8M/LLRcmPt76uqHnLccCV8+B4oed3
27LAJCgvLtouMIx9a3vteG4/vqIAw8uonLkxRbnldH1Z12USMU/xeeoljKxbtaKa42O3ciGdRn/c
7UbNygxHf6UFyHRnc4sLa+afpuxhBIa8BZ1KICQKecdButykGOKFhhri7vJC8Bie0Q7UzeoCKQgQ
uwtMhViGkyTCgjFWzJH6Obfy9WKS65PYdMTiFEdvnVfZmcB8PKaSQc54qpUSVEzkkNrrdJgkG9n9
+vrpjVU5jRW5EEO4MrlWZRNzp0aNgAKR9VOg9pLO1Qz62R/cerRNtx69ZpScVowbvnkh8h3n1vcQ
fhynQ+3ZPTHd1Lpcz6QWrWYGWZZmL+w+mCzpg6qs0OgS4o1lYLqQbQg6jAMVTMRehr4nxRQzcfRQ
1R/i7KcnfTYkgxAKvmfpSmhnKKEpQFrhYpBpnYEDfSNrPl4wDNrtdKu4K8vJhxntE7ugjsZnpyFT
dUj/rvZkykFtbEPTp/N9G0MnmyZgLMXKImCQbd06mpBJug7SMfBZoC5afFCp25AH14IdjPZma2Hs
+JLGbuMi/JlKLjx50S3A2432rH2oQqIjAoBUBOzW+MmHuG0jT3hkVR3bcOva0FvWJP2tiFvh/Qt8
dLw+45MBgSO1hH61yTyxC45AukAM006HitUl7f2o1MP+CoMO/MB0lov9i/3pXVu/kEEj0aMX7t6n
QL+xhPs9JOr5ifyRvhXUXQKUyypjUPDWEFwlXjyvHIdiZfHCBeq+G2eJEbhXYCRDUMt5u4dhcXT0
NuUyo4kHxWfOQQOoEfMT6+vy+R0JjHOvB5R+lLjqQ4LH1jHxM4MPcMgkEp5r0Hrc9NLz56e0nNam
g04qWPoMiSHd/UGg12p+aFCQ+096StaLWxIZryOcDUyb3j1CwJdVEKMqi9T9TyL6l1bAHFVJID8A
dcQwLIx6GISycBPc5wYtQ5C2Wh5b+A17CpdB1j9No0bpwfa3XGgm/x9A4jCIE937t9eu0308VSUy
h0fXzmUJGIj93TuK1NuO5w2WPHOBsfQeVLnws+fJSepDPaMZIS4oibbxyvtMa7JNPmj61icRBoce
vYERlJcTolK6YK0WbLG0FdwGQ/P6Nzj6gANn0vztVMkp6JzM4bIBFl5dGPXvyClT413YCkwPEZq9
c42Hp3yZrHVYLMjpHb8/pCLOG0cfMXFTm8/+wtC1vTyLTwTKlEpFfKKFepFtgdCRP7WlbrDE7NGY
psLoJ/tXq+5TJumKxoRA4nJXLX0WadpY1jghxmfNVtEB4Od+mK4oraWnqZLRqYTdBhYI4YhfQkVl
p6e2nComEPe33yZPUEqNg1N629wXDCBuPce2Rej74tSRu9tIxUNxqRyPOT/fQ1R38efQ2PnuWZtp
BxpyR25SAI1P+h0B4LcH2US9Eb0/0Qrh91fQ/gqgnYE1Pb1xHeq3NJ6lGCa3dtK9mZyGuLqBCXbp
5NcT12gomRCiWNm+JP3BJLsXXgRHrI4oDaWOhCOJ8tFZDkWqVcA53MAxjq6hcOM+ZSfkVOWrQPM9
S5NvBgkVeqDSSVRVIjpZV1SPgsLSnL401qLEn1ULUbbbmMmcCddb09NmxfXKsnVYBD9JTC5AMLAk
IMsFjO0ZCSqWm9v6cf9YOdKHBiiLzNtu3HpCV1dE6W3yl2/djrmDf5guz3aspO4gvuUqzLOyZUk9
177nEYhWJ2UXVQySA1TdlBGmyN0t6Tbl6ygxTsYh5wfW5xYB+lS9pKnDwuDHU0eatjOxcewmmXF1
VmImqdZZbedwergMaYY05TxAW3DydT/GZxXMeSnuxOdfb0ydIshcMuqV0hQWzpw5gaqi2PoVpUBS
juf0qH6gjNr7dItd+MFMFvXrbcnLqVcEW5xh961TkLXZI/I+kmADFhJ3IBrAq6sQL+OM3whinypy
7OX/C8o2yn7wrXHi0TYKSJfPW3p1lmdDf1OPFxC7pwFURZiJ7LjA5np/MqL/GacRmVUhWrI7oBy+
MyZSZn8r13VH0JUqnEeakXsZfKnBpNYyK1yvFZ02kkidZeYyMagDHfBe1m7zZzI7JdeauKa7VHhf
sFwWodzvi21bbMwye1cTX7GQ0Yui4BRCmRgHyt5oUdVy5K23XjaW/yEuDL0KfDQLyWLpW4IowkOq
zyNbyidqk6IAauYJQiiiKsN0BG5qoUmJdEYn3QaUJQiOywy2Z9K1IzgZlqrv/EHN+ck1SZYYeYiS
M7PojrwVyiV/N6z8ZPPlx7Epnup4XH2hTzvfxa7d/XaR5hB/VMxO51i+bqqqg5HY/8TsAdYw2RVD
WTJeDcK50J+nu4MYKM4xreDaDcr4jH1UFXSB53IkXoPm5yBq14MwTH5cj2QsyNCFTJzNljfLyZzq
/U36lWBriUf4fst1tZFcWBPWvslIFVrqaE8P+E57qQWb2GS/a7LEPvQ2HaQSbkVjCt044IEhLe5v
cuIuhaxMUUUOM1vt7fUihs+FfNr/8tAfIVRuzwUWFeLQf3o7AEWmb+ILaiQfZewdOOThotc9YXGt
EFoCiHYcL7ZQxED5s/aX/5qjxLrmchatF650HmUtKLUwSB767ASry4Y+Vt9rbsMLpmigaK8hCKTP
/KP8RbhrEQKZuOAI0xCMVTzug/RvGQoRPJZKukMRxK0GJbBrbBk1xcaJnQrTPyYUUSFSicacHQCo
5RrEAPOuHYYdh4mmPOoahk5KrFl1iOKzxvT7OvWi27RsLtWL7HnXT93452KbsYh1ryPtH83StWoD
L5t0cJzdkY9GtKxR0vmOFErhXMIpEs7opjUlsk2AJGA9Ii30/xLNXJu2kOoWoZ5uoYQYmWiD8jU7
tCrm1B/JFEEBvDBN1MiiXYhSRA69ama/X/g6tvWsP6tKxQQtmYU0SwQcp9pvq7DYLCVqPd3AFUV0
A9RS9GCkSsNF5ou0OrB/rl7/OLNdw8pawt1evtdibpeGtUFv0IHssccyVz+7BPixB0+paPXinoqL
WXALh7sQwk6LkbdHPWcxvWGw8Umy19+ITw8YP0/kTgdw+ThcpTt7Gzt1RvwVlWhuiETwnnBpevf2
aGOkqe3UOCbHD7r4rmPLfbQBhs4UbMe+35x7mCXiMQCnayrfitwZ8Klls+DsHlDITFa8ryqqrlDR
+pQjvQdUxvNUT82mpmYNt6fgg+IceB9lHQhLTWsvnbvcov0CLi3RB4xmNtjrGsKZOMAPtXO46yVA
Gw/b39KI6Dwx5/JDqeghnT5qmkIxbckLw7CB7uJxseFlaSvaU1zJN0yiIUX5k4z1dSE6p791Kj7W
TI8j9Y6AwnQ3tMLsu3NPXyi6zxDi0YyLEwoPRmdbIMizkLca1JJXbU0R9wZz31MfZf+k2lFiQDwD
n7i67LmRYy4bL/+9KhWFXdPz5FtiL+yZMKPDmTwjauZkFJUWf4VtbGjBSu76G93FjhQKfrDx86Ws
Xs3g5Ry1vnTAkgC2zVgmCL/HevAd2/c2YT95BfVrjGK+qgHjSxUztXh1gxg5XjKRAFqCjnApiwdq
G4MSekUKhEiQFSdpXOMil4cbziABs0hiOF3dXQtpu+Ia7aCB5vU0cU1gpfaIRU2fLLRRa7t9RujU
SCTeJaHopXpb1ycHSwUQIBVrAK5AVamm5WKwUQLlCCJsKd0+2Inwrl0YmPWqp1WPIaQ23xeSu+N3
DsjDbklTw9AYwmhnZ1YQxKl9qAR9PoqyiZNNhpwtTs50ZyFGtLhEIAeUxa8+vH2fg0V25JxNTsQa
1I31mVf0Fn3Q2t4Xq9fzDDLR2oFQkiDetFlYa25wsxmFpXHDnGc5BlQgNxs5mso/mRPdptihQvBF
vMvajlaLOz1evXiMhP8FcJMy2yC36lCi9vI01FbV/rhSTDLe84yag4rinmP/qPmiCTRn3vqOS/F6
oI8Oyekimu8rvl6G/03f5aOFRtKTQWNbhqYMlOrn7G6vFhgH/gXGnZ/gI5JSgb67IN0CkZNsMQO2
sl7aUGs5YfcB2smLVtTQN+4vBnQwPiJWihT9k2K3h48UpodU/R+IreJtQT2jOrhaCqfzvpuLMmJB
A8RNK6l0+NhXIjpVjWvHxBuwikRFfOVAUKHkQIfDr3roK+dmIGWLDM52ZLqhrS6G1qmO6EDskHuL
X2KLrUw4gWgIsBoGpvuY0k3Ww58bUy0MuPDB0jdW1MB2dh2mYjePn91fQioJxcGry1/oseJOe8MN
Exhu4cafHenHFH/8kHXLQzRdADeJoKmTvek9gXs/WtcgNqCV9ffKADWtMbaqUHuK8Fh057YSujKL
SrRxF0NSTyEBTXl+Xx1Ij3bieFV4gtW5r1e7au/b9BVLQ+ezBWkNFkDwAYRmcl5oiLO2wj+grkd9
XW2LRTwwkNAquFWNq1nUeUlccGMBgSpy4245MAVe71EAyzWwDwdsxXQeiVOiG4RIJY0dK9Qs3uox
SE3A2z4bPh1at9qLAAYrqiI3Dt6a94l6SXUgAOdhiyqWI/+4VMxmTfJ8WYBNp83eC5k/5cYQLDDD
pTMxYX/pSMlX2J36tSwJZF2eFDKvuOMQQIEkMECQCUvYHM4JGx+kz7h7IFQib0kb3Wblz7Sc3zE6
Dk5LhbXvyRM5YRuea3hJbhPN7AgmzJZrZ+3555AXKdyEq1wEkzpyLWoafnS/CjPGW+VG8WbPZ/3J
dVtegN3ldfrtWolOc6cd+EGl81zkMa49fdhET+CUSQpmT8jDZt4rwnoBs02mj2ysQ4pT//EcEO+I
DNu97ySDwHBlEqOWhnrqubw9ey9rSF9kybtC15ik7BrXT0Ek4ejVSXWwD87aAAGGRnjDKLjCer9s
ovyEUtirsYKFcB0vSK3tdHegSfJ1kkYBFLh/OrK5wxJruA4xkzNm41TQnfKm49SPGzOpAdFbMJ39
yYeqt/mPOQ2Gd4EKqVP+LAQIOPz2RDk2A4tNUko7CwM1etVVYFwYC4B90ztmko1uRsHxsI8tHoS6
wC4Bzm4eIWzj54Z/FpjGB3ksQXNkoz0kVqOtDKZ7EM2FXqWyycByms4b1ayvPESurPyvxxPi34pt
qDvY+22STDcuRk3wL+3e3X0xeuW2Kv1CeitTrYfqsamTHGsJkRJTCG0YyaH5LxjLKcAaRqOyBu+B
5J8lvCa8pFl874aj5LiR0ysx8SPkx4wtDdQc0f0dUpNnMp0U1PhOu/+Qvdu+PfX8hHwlo2BAJwXW
+7Rxhzf0ideNaEi6IyTtzGIcVpFwaW04scLSP/gUcWeCRrlDACLI5wCHiSw8veBjtLRBKitPLb/1
xsUZ0iHBtLSr4gyIab2y0C16hGCTO+Pb+gO/OHQ+ANV4FuCTv/QZ3+7+TeyP1WmB7AjZw27EZQot
IDz3pOxgwXPXHK4VqZSkqVV+qPVNA6CuzCyc8R206iFFlMHs5DOCNw3NHNZ9GsLMr3e8dmS8EvC/
EiX+3jPLFGtEtirfM9LBSXUJE9nADApNP7358sDlJH6tA99ALzAi5GTS73qc72tt+VVvYSC6FKO4
vPqfCqa+xzVznPqg1XDXgGmesRlPm5PwggQYTVoCZFpGOuX6AOYmpJTZS8Cl6GaEswjQ1+bHSgMz
zY4qABsLqcQMzu4Bm0SfxzwEFo4B60QG9yPVXg0Jsi91diL0rpybbaUQAF4g6k8if7JDEUaKDt4z
CYLI8TxXwb305idciW6IMtOYgRvakrk7AdlLc57xhKTMUAFbSPGiItR3Ilh0F2h3nMR2QnCnB0jb
olRidHIh8GP6fKrUiTurwQg27z1+f5W96XlsrJUD1jXKBY4Znw2y41EjtBcWHGqJGb/YQEwO24cQ
/uL4iupWWkyTaTwovT7Jv/FCjjg4AYt8zdBCG38nyFusTqVMakKLuXgfb/rXUogXJJcVMYgm2Vb4
EM/MQsMLcoN1Kd3z2D6opapiQrzTfE2ztAHGLcddaMP6KWdDDzVwbZ05uK/8q4+WWC1INV44xkSP
GrHf+btMZqd9t2BP6MP1g5ltBlHhIdq4TK6LPqXlzE728F7ZfEBDoAMXw25RoTHjqHsj3DZ19HxG
4cJ5YHFjoy409FdYHXS3YHVaZWZHWSCxeLTJRfpYA6GKc6JCNFai6W5dfOAZjTskD76sQSK7IZhL
Yfo1Z3E3eQWyhIpUkDVY2zO1Aedl4e0YxQisX2p3YWiMiCZE6h274l3vbnTC16C2gfleDkUHTuI4
u0W7pNHo4uJuyRr63914uv/DzPmYcgF3zBncAj2iyoPRHjkZSYzeU3CdFgPvJzNWwOWJoDffS9mx
hMX1KbaZ/QjzRPIgotpNUtIE9yqW1PXivBHlQjVgeRh43Hf0KVn9xNKiUMNgqHj5m9kR1Kv6tVX+
Z3cAOUEGXsl9f2ddO0nYpKlsyCn9yZ4hk4kA4s67mBp7sgtYXjqr+Im/vPJcBiFzlkNAXlRDvuUI
WoGEJSuNMeQomnCDmUlUfiefIg9Q+p0n1VT1wzpM572SuaO5aZt5q89zJmbNODyGXwVRHQaXRcYh
FWdSQaTpzJF/u7wm69rjlWRNX9acjExQ9jdN6poW/BT2WxKg8VkqMe09ZRzsI9sgUZoHJe9+Lv0L
nhBkUDWlth/6HcBexhcKQaGruZfRh57YXQWm08nJbHLBlVKcz98Xx2juc8qejUqyX7q9GLTnI/Ae
VNNvDSOa3ooMWOpDyn03KPJe88A3kRySjlSFJ2NFjoSjMTxBJdTZ+IWAP4eEM9DiyJTPwBR6ut0k
KAt5hfSrZXX9wwJSslIPuLHTVVYT9apifIM4ctKETiKl3Ml5W+E+bfXa9famW4GeANMvCsHq83EL
0ZtpT0s2C0DsL3nFFA4UrNJLM+SlBADvqUKL5h82r7VwO7whkRszH4SKg21VVabIeTXgFYOQ64NA
aFeJDvI5n4j4yspqXCMXLoewWWP3WS9+AaaRl73+z/7fsjxWYIzZnG7LfG9M0+jOQo/pEVoShQhF
7by4geyIYgdUZnOQSJjfXeQYdO4SBuvvZ3bO41rkSFZoNIEQXAw4crayPUP3qw19NbauO8UCUI6Y
0dqrCxAIiradri4fbnxN8OsRHlidNH/U52bxc1Au2XjY8+u2TH++REC0H7xCASyqFKrxVUa0uMMd
Uv53PEsvwle3J7UozC3n9pj3pIG3ZD1TJNokGD8uUFVBbniWx3ysBD4gqQcTJaWRKZQS1UOc3sUK
dCefQUFaQX3TsRe9U5PsgZH8mowjtqIIRAPEpnMjSZLwGmA8KUBKgpHkf1ssZR57UOaEq1vUSl5T
JqWIAx0tcnAvVPbqeLE2zjfrZCsQ8FdweJ5kVlNivgGKnduzB7QjNLdmmSw4LA9ccW+wK7DPpjgV
rAly2K/YKNIysSw0vyv/8LQvQkVfDwproTjrYlBd2S8Hr2TebNlUx3LbNJed8+6bsIWiFDDm70L9
doJ/wr7HcMeNUCWQ+bCdU+pSnze0iO+rbu7k1YLdWMludSXLlXPnjDEDRYv0AGhvMtNPoVMgEX5x
NtxCgfqBWydPnluWbqp7bV28t4UEdzV3gW8m6BOY4LQrEixR8hZVoHQ1r51cStPkJ0Vh1N2Lru53
XpUV90aAUfMSnnWhOu3tpxwlyitR3Ywc6wWkSbE2yrEwynIWENhHgT9/aMb/9fxw5566R31r3TjX
wmnOYA0SnzCbOyVMyIRmWMOlf4D8N0eltyDIfxn4mSs3xDJWKVRL3dtmKJ38C9fJ3z/5uqAHwBn1
zC3/RhS+RYTj3ClGk4HmGzdaRiMgZhJwQnlvDHHhODYWYJgFfInUzkKkF6wUMWPMGajM1DOQhaoG
unZ8jYRYTfYpAGxdFost2zovg+Z9bIzNYcK0e4UttwehgfdIQoXy4MXydPJLNf97713cWGtc9yoQ
Ebn693dFUUG+oLmmZ4Jh4S+Wi5sGoV6sxnP4/KkP+VcIF+ChmIYJQc37TqoprG55Vkjnd2DtMs1e
WydfdDD+o3CtF8uIeaIxLAjiDx8h6EdfTpotUopHQuiPuBW8fzioBC4GqtOnptnNhI8tySbwnY2Y
wXV4FEEoopvddRd/q6OOYMEYarS4I3CugkDSPT2qAL5CjgDVb0+/8aXbzTPzRr/2qtbrsCXZUgHM
NP7n5I3OT1a5tl/c0kBF/yf+UggpGza5TES/LSfv6rlSQw9gwlhESiJCx77rhtZbcuLd3n4kchC8
jZtggIvSEun7rrv+eeiGGyRFkhB/qLPPo+klOtPmhK+B7MIC+PcZLwJ7QhXK6ccel97ieTymA4PK
ntjmYRaZg7SnulgECWynu4oOjrTkGMvxmDvZSWS0mWX8JF26C/7UFzXTWVgmb/mbjngXDsZsIrtD
ocs8rBw12tiOpVN3cEgL3K3QJCFy2FuSmrKbCjtFnvEAEZEw6vuQcxQEDr9ypMfYriB+E+6gb8q4
2D8PsMeWdAJ/M7wQaY1vepyQqstWuHXW1x9WuSSeGa8i9pYwsO6PYEEuULAlKKYfH+aLPDazrULd
lSyvnpt+xcjCgFsUSNGog8iqr4zno0T417SNkZlvNmybQqRsXi9RpS/YZlALramvNqyu33dzkuhC
DA6+zd002iOv3H8DOs2Ix+W/z5naYLUh2GLEF5XWOOLBB/buqDRoVkoTPnf0lhE4gJ2g1DHHvZhE
vaSuaHwscp/4dQv2gh5fFQrrDjzPyig2BxoZ9EL0Mt1x1SdnozMdQteEJrrbuyh7Yacqh7NIr2vc
8qCXNSKydBMA3S6qn/vhr9OAVJh+xWCGwB/FURF2jV/Wdp/iKxXenH1sItANahmDoXvX2YGDfw4O
C9r3yxBk4hcIlSIcGmuOTqG7mTJ3rHoH1FsQhlZ5/JHuhXtewUW379yRT9oPv1XIqZv7gGHPbekC
1oDNip0C90P/LWO5eRXSgL3g0CeCF9LbaNt5rMdmAhvPKP8ldqPKaEihD+VoVt79AQ5366O2+a/E
GSM2lqUu4l0O65Vm0A9/yDzBIfKURIrCeb21T9xG0lW3Oaeh6scBtJEpFpOo8V9OYLRwASFetwYX
xkrO+C6DtKvtWbm5uHEpL96ubrCJKkGn3OQKNV6l2k4dNJ9FYaT3RwCC3Qc6HQU25kIO4HfZ+kVu
PJKmTkQFlyuKeX3pVx5cceFR7Fiw+shM+SS0fT0XGYVk3o/G/zBmTCczwgOCI2Ku+1gG1+URnvnp
OQ+EuTm89nhT/EYJhXOHHng/ca0B07BIHRaNeJe8TtrOA0hhJoi8jq4BLqMgzfOzUdBV87kn9PNi
NmwSrN2cm/t2oinb1fXHxJ1/QEX9NUS54e1N6lG+C8EFWofHatGQ7SVRVvFYrA+i4bt1suP2pIFz
AfGVmlH+El5c7EwN/zpBidzo43VBwob3d9O5Khq0l8mIyNUj3OW36ztBffASIU60lePWhjVlSydH
+Dh9Li1GiCZZlpfiDPWOaARvYFt0wKShKKZFxcG8YzyjedPnWffVDmRDFaN5oWUE+9Wv97fVO0rj
qFi5ROuRjypQKKp66ZmqTVWnjlp6/DLzXOhr/sQOgrs01BFhTeDJBB2/yfskablrnfOCVhiMYBro
EtLPyi6OTz9yH8fTkd8qjqzflyaK9bWzN3FvbvTtsNL7mn0KXHwAJnRWnlSf31Q5a9lnicqb528Z
koQ9iHlYXtb1WhVNg1hv4j34syxq55+oIqI8eG7dMYvOBBlgyPmjsSnr2e2KiPB74ngOw5o71MfC
NPFclU2dTn0OumcaJ35KgG6rx6pdFDLOm5nIn2kSirESJt8KUXcERxaFm27elxtO8VxSYRiqukXT
/9bCIgxpwBI+BkZpP+yhFR1A5KhoDRhZ0FEq2UK92ya27Q8CqihQgatWj2jkqtRWbo4N5TFQVYzl
vFLZ4Ox6AvMYQXMGP2aC3xCdKkXFVxqkn3q3+iA0e0sv8QUarvXiOpk9Y1zYhhFPEkH38A+uUT5J
eRVAeMa8o1zPcCXpqmP4TVCPhcR9jZVqQVpLyewbWWb4bEkGTfADJZ6jG/c6B78KWZcji5EXRjin
5HIdMAWo0Sj/ABWD2aSVfBA8QKXYqAIl9lEEnTCLPbyCtcC0QpcNVg1JFMmt9D9H8ma5Dciblevb
ZnXGk3YCJxyuEH9qvMVZgJ82GSvlgXT2JoG02cEYgwY1G/N5DFjj2tWXh39b/b648AQ7nGu1qOu8
3JXxIii31NnyEiN+q9j18IXQHOuZXOZ2BCeB0nb6b88Q2ZeVqiATy84UbQv+zEsd4nSHTivqUVOB
sF+BYAcXwYz7QfyhH9u4Aj0LDO6Q1K5DmA/Oli4bCeGjt/7vA0kfnZrTHr7k5wD6UgTVc/rqp+PN
edSWG9djNSJ9eNszJjb/QTnYWVMEdgc5b8z1/SNvTZmE2gvq81oZ0zPIpCn2Vpboa7W9qf2FRkvt
orJdoEFBcNV+Mdz4vd28enjNjkYDMTDVAa6rnrOscknMhxWCUcVkvTdDBgZPU6a7TeqyQGL/6wpS
LQ8WeqOYtF2Gh/P8kD8TmSx9Gm40IRGscBzcuanoIDdjYBjJaIl6rG17FfZTcN28tnGCDT4BsHqI
OVWWrBg1orUTnKPgBLgnWMqs4q/RU7a6TQ4E2LCtQl+wtMYvrzBLgCc4cBlj9fkqW2ZsPmGkmTWO
KjVO5iJH6LwygtHlQBR/Qu9iwG0qqqv8IlmZRqOlhZymmUJUba9VG+xO30cJRKZDp4xuOjxYPhJE
kQJzZpeMqyD5N41KEo/pasQCMfNvjO5Iaqhe0+Ni2V1QxsI4nK30/ryfREeOSjI1uKA0NoBQc5ZM
CoDAHTaMytRR8FjYB87l6o4bicDucctTkdRBJxaKc67TVZHgyK+KhOFT4pdBFeBC3CIDWR/W0mSr
pc44aloHac2TbOp3xopEAzQnYBAdNjdEInBlcf0qNyBcoALDtIJ2wDnZh+1G+ZbEGFqA3Hbxprld
B7mjaM9ug+FtuM3lSw2fmTfiAU4PEzK34wtM3Ll0biq/SyllrbwhU/P6HAoHlG8B3Txoy41KHSTI
YxuVxoDZA8bRTdCly3ekrx89+jVYnBsSvgMFdtDOVhgNW9V0tVOKGcwOTOVOxX35fz8+swwP1Nvc
vgy/hdsbE/MHFkuS/k0f7NZaInIm1SJNSJIkSEoLYucn4j1QcEllwZmEUIje6I5JKL/dAP/0x4FG
4toz0D87s72+zjXjlAQmFbQiMa8VUmqP5XCqBIy+U9Jah2DUFBKIFuIpYuOBOlRLqWJ1eZaWCvaE
iVTR87rDBzHDUBrnQvkTSMvGi1LKsjogA90DY1EIQnvfqook4MkcAfjjid42msd1LmQQTazyowiW
dIqQWdFvTfHnErMHwIIwVIcngPuz31+WDrPBqmX4o94VP2rm008i4kuZR8DLWPlMFT5Tenym010k
mI6brlp2b1P2Uf8vviUlGXHTYSA5LSM84HejA5p+EbhLDwH9FyxnDGeR6ZChCm7ecPmOJN5G164z
Bb/zIFiJYVg7/1plvonA2r9ykBoY3eIISvNJIEVFmKcDVao6QmedASp8uatKl2wQR5M/bu/gEoS8
CmaGlEj1kCwTaUqI2e0XNfriaJp3KQN+F/xpwnBHoG46eEHQvRkOMIsh4LdweKAnX06vpaHnrECa
43bgaS4CY6jeLXXjdI8r0Cr2Kh+kHU4shf9ubf32hjjSsHEutwBWG28ftwufXbPGimLz9lpOcKic
z4ObPSShieEwKltc2WPDKRd12NpLhkwKw7e8atILNfE5IN1AqjEK6yi2CiyQHVkeAd8U1KkwWZnJ
kg0RB2Wk+MkOayI88dh3t0ucrCoC88adg3iY+lvg6fv8xoQFMP517LwBTeqhE83rj6A/9EFFMJS2
PJb3gXlCygxvHhBYPynt0tQ5e0alyauVvrDlnK9S8NGtMD7TbVp/fsasKjeKlkfXrPIGmgTh6va2
b8v3PE6ydwKhMBNCX/xsNAlXtkvUnNX3uKA66Kr+q7FF9ftManCK1hbc5JabPNHixMnR5vqVQj2Z
Vag8++qIBOvCCB2hf2niwt/qlsKWp7ChMX+9VqqMI+1fOKBEvy6tEakbjk2KwgTYETNeURONEZhb
Vf54LjxZPX9ZOi03zm+AWGj5uaVEMMHjCQxP8H96H/oWNz2X6xsPZLDvNEvl+56yu9BvP9CKSLWn
InyjzLm7+8MYVBpT9QfOe7pDczvC/yCZuZQGtyJWmtlOF2omuoSxCFvrbL1sN2IBMWEM0jkrv53v
7YB6EY5+vt0FA/Qe77vWLwlBI6M2BzbEfGo/EPbbA5vURqIAyizmnGLcGrqdSwTFHtytgKvmSkfD
ciyAhngElQmk3XI+iuL5zuQuDMIH15pUA5pgYz0rX4bgY5oXmHdWkurWAa0XZyKRUGgKmYAWEOl6
eKgT9lkGJ9ET9LJqdFJ5ktL0Nlk0V33SzPAF4zz3QwX7h7SBlgoqYCDKPcP886oyLE84qbV9QoGk
QbJOGyKlIvExAwFaoFNM9EFhhb52kmQb0lMqaV1129oItS/060Hls9qmoIvTbiYy4Sc0Is9f4q/E
1+SEcKXn3gRRV7U+gxI4HjroJmCWlQwOKkPcj15LqkWfP5w9ehqj7LmfRQXhKS6XKc70SleJXqi6
W0b2fkFj24j4CGNSqbLjdU6wkDKT5v3DcGSxTjaT35A5idscduLvPwXqAfl2LbCDM/bV5WOaSwb3
PJtaXKLBTLPFdmG7VHmY7cihO5ec2spyMyBhfgSuvLat7/HfUEK1am8DLhj/EoJC7SY8iiXTh1gS
oK3SM7NVsbNqYR+Xj6E5Uo33fJzIlTSIt1luN4ohLM7IiRFJXEpit+gB0V6vNU7tvDT7e7WMEjFw
+QB1pzzeRNIxjUaIQ4rRQzt0o/fSSdNLSCfCVTdFMfDNj1romwoexv3i1+6ZP+MtwBxB13WH7zT1
gqG+jgaeAIF/LwrnGYYR+SA/5aqjwHdRal0uGOYF+RvjEFVFXridVyQgu7wD/zodjRRLMlViMqxQ
iF3sQ73tHLKIRAYR/9sz85Cf/F2l5D1mzo8fo2RIcSuMNDFHhpmASQzsjE+lseYlgFoigNGAN0P7
Q3dnu8XnyFqqtgxRLhL+rzYPuJTDF4lGWjSYsbd8RGTKGtyGB4+EqZGWAQqWGT6ES4wGsBJYNWw5
d15gpatfMWlJVmtds7+Jf1tmPLG6zz8dgCFGFP7Yr9e8Rtcd/IESHmC0tSoOcJwLtt9YOLD5rKhj
ciyN7CN5/cBH1laoy8UPIfApzRQCkl77P46eFynHMWhwnMjjxUz/vxCymad1qFHfuffgZ+LF34N8
ru2C9ARlir2QlyBl2nVNAOkzvb9BjC2MqrvYQlFM645pvfzXE83OBYWyFtum3/haYAPa6D7JOJCF
Jp1zvOyg+7hG14Fze+iQaFFxr9lmH567i8Ggugm11vQBkKaidlGFSja9SUKtql3rGkJCB0FsapxJ
j2TbCfx0xUgl56Z1ubefr+uCzK60p2fvbmDfpkKUu0dlIE3avZvf6BJU6/pnOegYcke4jgsqXZX1
fjkVx70jnNZsvyPFAIbUJQizgICr2YvFpXpJaC+9fMvvdogJuhSloXb7QEN1xg1Rj+j41LjSlxiM
2JXs+8jeb78C0pqWJJ+K6R7lCB4M6wMwkRyM8cZ7Dnyl1m1YP4mj0FlhEbihecRAzurl5HmNXrPg
wY02YkcDsNZjiAs4M6v/A+8DOBOxqpK2yL5oo6gOGL65OFFK42AIldiBwm7X/QAQhwROvpgXLDD5
XVAhxY9IOYZU0Y2fpnZLxjL+dkTjDaTO7eH84HDXmjGo/w4EkQfFGXKrqyXOK/ZlaiqSpSWkqEdp
nOKfSLRK4HCclzswsqE6zZPBk1kfvx6r1lJvo6+ahcsCgpk4xuyDa3islkvaazGk1KAc53t8RQhx
O0XyaDb1dOnUMKctAK+EsLPLQzHXHl1X5rrvdipuXXy1Qo3zemVonrJxgTCaeIIxuZinyZ2NolR/
tWXkHyUswZP3wDA5QHDrK+GvNDF9YrWhYcYffQfhgndQ7OtdhgT5ad19kWfFEBcCs2qfXagWQKSK
8PqJVysGjWrqA6corw/JDiBs0rk89xb91Li8xL4+qIMR1ehzkMql44ZZDOIQQZuGXNhhOmxgm1Eo
7LhdyE4MLJo7x9N6/TemshLJVQzlwIyT9RDEVC7c6YKqr2f/7KBQgE0ZNS1oAPwshjSBj9IaWYBx
qSg/x9myS3edsUgqj2VFM2nknf9WRKxcsC2EduxYIV1XE9Quw6uFffAvlSSYxouTx3wwVl33ud4d
ssNcyuLVx0ceTNAEXUn05ZMS6B602VCSOnyiNbVghBHrDfkwcZ2UY9Zwgwk8ftMELfeGgGqFPrJa
YH8kQIIz+zh1rS3S2VmuXTM2dydnWth5zycGo0aFvosOw6M5U3+Vn5S/w3YOleawOIAkBVYNaz0g
mldjaFzPv11BFEgHcOQbbEQRmiIE9OgzjoHlJHi9QDu4ejPmDoX2Y76mTAAZ4AIK4LhjhEDAwESF
KkfnJ+4Opp7SCxoBZAEROFGs2vE3SAe3o6ZIpZFy17kENXv+DF8kwsIo9TL49t4f9ZkNi03eYN3q
B2kfHOjJu3pnMYAwckCKLfBoTqvkSLWrXq6mSGZuOiCLVrJq09gF5bPTdaZgC0Mc/NBMxDsvAzqS
upb3co6E3q+pk1Uq10CFFW8xKdN17fc9ZsmonX6ef1UgkNGAqHoCpthpUGlK4RQhzY95U21NBkia
lG7qb+CE6fda+1VwD1qSLr0GxNMnQM83czWIgMzwLVTy540tX4XGdpu0iHMGXYfpOcAVIxlU3lIj
CidXJArh0gbbq5ILMWQtz8ZAubWgvDoQOp+2PeTAlMfUIdF6ati6PHkLxNA2DfE/og7SVe1p1B2O
vP2aPlkVFL8rQtnMeX6e5Vl3B0kjO1Z5cNyneE+34tf28GDz2M4pBMsqfOieMNWfhINVd9TogalQ
chGZJjtnK/TeSibr3pl/yn2dJsAIIKpemybJCn/WqEVZCqtvKzyqPQR0NvOzgVRSp1K7Xn44alXZ
ccqfChUWfTRU5BueKAm7K1iogpSpHUQhKKwDA0207qVfxol3OoICYZWbaVmbrmXvQ8yPOQQ4A1D0
wUVbpimLZkE793SK6IHA/uL55f19e0qgVGAH3YuImCcxdVKwv6MfShXCDz3OSY6UtUhtF+kAewOi
XSXdwojU//9PwIVWtNuJwN/rKxHvcCoj0gR1mKfsBQ5gs97MkecQB1R4UkNb7TQstBzgviIMSO/K
9mABzn/T5dKFrmBeiImMkCsa9PLeLO4cLHbUzCCkw1/RjpNuHC1e/xDSzhYRJ69jnxNlGKeCd6Nr
UxrBmOGF2o8YV35s9icQ97AShkHtBM23cW20O0ESCsoDqKBTn/Qz+YlI1djo1v/4ochytiUMRYtD
ri1gMF3a1ldbjTAT+lX3wyZBJpd21HG330EFbVKwsJh1+H2qhL8DuTP6FtNdv3sjsgxJyAFuARxu
ETGX7sjkZST7HFzcxjWnBJMeXQZL2uDQpDhjyVvJO7SkWxm0RmEtAZwTbkgMnNZi4jKid6OCubzG
kVlH+0HHt6jYrPFnitjZ7ZputXgDe2e6xjttXlvD1QI75tkd1hbZOHpKWjPgHpxa4tZ0ifHbYIng
4n76CFGeiWP3GZ9TAsSCNEkB0OoxvCx3a8xccCZqdJwmzn8pJvqgjFW21e4hNxvVF5ggVMs6TXDn
4VgDe3DDKUII9Do1k2POCHR5G5Ga38RUIqEcxOmDU6xqeAysdaMVhvYSbW8U+TjZj7Jr8fCcWife
2qdZ1D1ZfrzaIST3DOewq5XAkExAt0Q9EmliSDFT0uf2b7e1a7IZtK1rv7HP9/Y5RjykgIuFAo6M
SLL95zp9noIrD/bBBchQATszGHwLUr9TxUpedLr/VKWfHyXXalMYlNDfa0KpC/Pw+RgeDA/zlLYD
tayBuYBGhx7O628Y7exZ/JR1EILyx7r+F4lKcOwvw3jz+qG6A3V/MZ6diu9KJ+gER7+6ukeN/c15
Y/oqVAOFAwsNzQqPLP7B+WeSsmJjTcIT9u1eSFM98NfZX5qDpFHS86Mn0R9ZscPveLhQ/tU6EFbd
XtKSR/VCwwKf7P6G5RBtGhh9t22GynLBAzjcRMElaA9T7iev+PXdZZysO3XTzKWLHPFMUdbMTkfn
O2D1jE3jSGv0+DyfZSPzLJL/70yqTJJHWqc/6b9YF75c1uoNPWShTA/zRcSfoJUJvxVkhN7pxDRc
OoMuPdba+9OtHBjOL/B7VYQ41a52c3eqRCAdpiSo93s2xusP5hiZaItYqjLjnpMqQs0i0QKA351w
E6YFYhiCiOcnoNdA81hH8cMM7sikzkLxtdjQKyAID77798ddm2933aYIw6bB1anc5jyL4r/EbdZt
InQXvZ/dsPE3nT/qBkw+0F/VhxKZgAdFzA452lJxu4kDJNOasxmpQo27Jo9JXOwycFf9qOFOy64+
LDhiiSY316MnF8zeBy+RwH7o+r9PBudorDBH0d1cIBMqiFWTQumxw89EKOPQQo9uw/s1i01G21jQ
+r+k6nZxi1FF3BBmq7w1/4m8jwL5XHhhz57KSuKC0ekaVx93fd5ZTQD9U2E5VE0jfYwxQSiLUV0O
Qa2Y2Zg9wGcKW84Cwv59NIzCXnDD1nT+XJoDodakCtWRtFtc1EGpEXl6ZDIsf+X8MmqIKQCOWZZk
PlYhpnMrmCOo9YmqO6LkykCWzuYbStU5g6PL538MNUKKAEpRD67ctwZGBQY66yqbRjXRYBhA88RX
M/Ts8vOFoaINpezfiDos6NGBMWi4lAYMkQDozffuvM7ccy2e5hCW0XifHASk1d0eV3f/6jsIzclp
LS7js1i6G9EmzUB7OTpdLoMTZ1JkfpZHiR6Pc63wakZgEHGqIbvpij04/GgpxYdWoGxGVlroshT3
d1KQIFmm8EQqW0mzQt+0m9sz7Sh2zJMpw6wc8qy0ab49/ptibxTg6setYDuHPReidT+SczHLxVff
6luGL+uf9SYJr0BeJ4+obdlr/EVYja7Nr05H+zFBZJmegyVtTxfV6HXOZqmxloE9tvK5uYsIDTmH
9gW7lYkMJwaVr8tkZvmoORMDVnnan+VPxa0hL3f/qbiyFWY6iLi4pbONzhKbMt0yMEfIOLBciG3i
gQrMSXkkjJc6VRIeuHz11MmnH5T4kbDoOh2/UlLtvKJ9w2PtY6jl4g6QBsRXlC7ndjD6vqg1nOxo
WRfVrcObpgQs88v/yWkkb3yfhOc7wGuoVBCcNkouynI0X8mYCqSzm/OzTUdHSoYrg8iVWsvx9Uyy
sv2FoLKSHYdphLRaXR9Yxj2qVoGTjRs5tVaTHHwg5Lj8lvoawsnctc5rttk10Wcbt+hfYc+S5Q/S
KxK5iiWtvUkxQmvTgv4vi90TMDO8csrYSQZpF8Oxx9tL4jEJLR50qAcOuXSavv/zLKHnKPtPi2Ro
X+jeqttb1mzyju77oK+pY2DGqWLPyePGn2C+b2fEoetLQolG62xbZd+m7f2AL4DyHwdRCPXQe5mJ
E7UykqIjMzqD4XTtSSMnw1U8hlDqzvjV+BAjX6rQWwMvlLLkWH5+WbcA7MVzdI50CDKBaAmIOSS5
EKwlwVU0/Rwm9wIxTj0TI5WYUP+QEu48iSwl88UNjNEjzQZnhMXv6FzBPCSYMnblw8DC0z0z4b5l
uWxDQXP4pqjJ/5pEP3jqcxzA4BprFdtWri9TTc5ukXbCZv/p9tp1fzfjP80Wscr/EWeh8QFndSm4
oKPK5u0kz1Db6z+DuiZN/vYKCJYYPadlwPbPnBVfy10xxY9+f+YhjTikbRAHc2D+CCKs10SPNmqZ
cjtQMo1IGwO7MKVws8dLdvh+cSLIEpQPL8asIRkZ9Vln6WGok4XZ28MqlPycZ8/VqpCmb/BNsX7z
i74iO/kIBPDreVmhdhwGTurtRECP03hnJky5lanP4fwevWZh4YgXpHaPujHbWWI7Th/gRCaA6s4L
fcG6kz4KaZbtNWLiv/34VTob5qegIXRiWImsIWuU64Lm2JYQ8sd2cD6vdkyN6lvHa0ZkFyQZsPUv
tU2zePZ/SWEZcpSeJFvHC+uYNVoPZ/zBWvQbCNZZlpJceTrYm26QBkhFo/+71PE3XhZSuEGq3Tm+
+9KHYBEFS8qmPqhbN4xr8haakLJm+kov/lsRQmxYtCGHgdIEu2vwRc4Ipa9g62VD7afEjtBUibdE
n3sqyz5On9mFAcSwbdo5+0kMgIfhnWRJuY7npn0UUIX6UO9v8CtCgrVPODA9ByxitRoizldbLdQ6
zqfNvBv6yrtESNSP0UVByL+WecOY0avLU/hcuG1x2HMSC0zrDtjXfOrj/ImieYbChyo+69i8EzWz
W5hHpbuOrn8PEidhNiaONYI70x8UGR4Z5v6XTS7VpQyH2kxb9MFMsafrkiqlKtoNp+yx5BW5TVf6
dhr++XfpgGxbfZ3CRALrGzoQgMKdnoqDFaEeXA6hhEdm0KCKRtt9po9JXpKw3Qn7ZSj0Cay+h+29
cZeBCX6cnU0A62f2Rz9HrCTYBCaB0Y6HGTWoRcjNLADxvEyKosBLrRLgfArUpWhmFu51qmq3g+YH
Hhjz6ryHfvbkSBJbJpaLhyXk/OBhj/HaVAZVAgTygTrw6Igwpfoqmg22/U1JhSLaUYgDaKcT9aK8
y370KN/8kjCKm0jFWU/Y/gmx2Hz2RC0Ve1Nb+iJYP/2r8HxGqmWHxuGlr8d3N5NuDWwQznq4/wWB
NevWGlWF79tJrXB0y3B+F2SlwQVND+L+qpDEmg5Tv6BfD03s+HLepbuHInE7keILPIfvOQNJvrTG
EGbmBmuTmcj+A3gVmvI1PkkuuI0B+VxqeC26+u/0wUeDGCKr/Nx7/+DPJvXPLncVDoKe5QS2JfE8
8rhaSQNzgolbfG5AmqXt4lDFZIz2vbwlnAYbxHRa/AEl3EKedFFIcxTzr91wFjCzBJlVERT/vxqp
4F7JdFitq66QNiVpLRc9cus3DeKYsxUMflU2naEXMQo1oH/znaNOSWouNqA/aUPsj8/vltU9LNK8
pkmnDJsw/jjkA+dbuk6/qITiCKeETchi7MWyqIMUE8uXicMr2nYU2I5QilFD1p0+z0C7on1ZJBE/
vGfpPldDDILm4ZuDVmw8sV+df1CXji4+cdb6s7XaBS2H1C08PfwZuTkWj/qhMLTZMWuHs11RpUxZ
2n1hDgjM2/6YGn27P0WZts5JQTtwfCBfKqB9l5r/JOGVhHsFPgeS3gtXjUZq8zDJNXcgY5IQWSKE
CV8qGedpJ0fTop5O51uCz0fR2/dFqmXeaM7oiLeLADs7GWIPjge72LGcGpqvxpCl5gLDGqgHNokz
3TKQaNk+a7paNjNe+GFXWXEt1XN6LELgBu42Sl4yCFW+hk42ZuO1ieAKRFqUdRE0rDzNCI6VHG3V
ru/2w5Kh4sB1Eri0i0gt5BUV7rWKaUY0iKVbI7KVp1aItRFATEtDBIy7sSDKDRKLPK6GPWaqDY3Z
5C9zFOoFATL36cKbWMwMetlm23tlaID64XtIhmtnfay6Xti6Z5TytuiNZjyVwecrZ5frt0kqQVej
MeQqAaubkc681UXjftrDlrU6Z+SPKqZrkWVbgi2A77jmvM6QRYRWiUoPwxQnltorsXGj8m8I+zTl
RExYTqNX0xAAChotlnY187XUHw+TrO7ixEy8ynZ8CHqqQRxUpcLj5t/PeqR7LHWdEhvBQs81nvfm
iAlMy8FnidJP4JKglSGTvzXtxa7nuCZZ1Kg0LPiikZNOK8iMBWmZhij3F5OWmmI3elwvPLIVzAqh
Xnvy5146q7mivihql4CzOfpotVWx0oreUCzuA9nhdtzAB9jVVLg9ORiPSyMLsHvHAaelkhESjEP2
wH/KppRYpnK04Dik+N6a7U5K6oyIhvu0kCtjOVHSzwDTK4P73pk6zrhKBIPZMIyB5VVTpG+NoMNB
7sb3L8Kacqsah0yhDcfnIadb3skuM9lMMiVmZKyT7JMfFgNjQnu2+IeDkvdxF4IGLJLcp3GnzLa9
VVfk/1coEnaFs7Kf88p1FNW3CKsmcNO8Ph2lKsTa3pU/eqyE22HZAmRT+feNVAtFBy88J2JQl4Al
CZEUxX22NDBlD2yxwTa0rG6Q53tu/vT0En4qe4wB+z+OyelNrFHLkbrozNEA9q6G8DVCH8VQzVGP
ZCxc9kklnZ1i1y2JqRWruzIl7A0j6Yw12Ge0ih0XYG0H13TAVSGyJ43R6BcNVvy+KgGbG+X3M+NS
cFJaSooyjVnuS1tXmeoy6SOYC//wkVLljzyzBBsMEEhUELrC4Ha9XQmNFyw9glYO/hkvNEL/FTmn
yre09aLPcT4Vrpjebxzs89XIOOS/xexV1GAO+QUbMd96/lS2LpP/BbDuHhFa4YBjI2KfWBw0Y0qz
tP+oIo+p6lPPDhUrcgzq8+TFJuUw0hH7lOR+Xr//m+Hx3t/miGlYDrrEiloO2R2aZHYHM7dNqvVY
ebsHMrh6NE+Mw8ka4aXfWdxhAxshoUNIccy7jl+dcMJp5/ee4VLiXjlg3x9V15Dw3RTgh6jab67m
MwqyzqKgvkvZxObBXXTnEmdTCRLuE2nXUzCAYB94TrZg6oWTqp0U7USJupYCFiVb41uMbxKcqVjs
HOnjpoiUEAJLnLOHHn87ACCwfoL1pIVwwaqPXd6w3l+zxK/LmnXjz84F0/lgqhP98aQbu69Ty3e9
bWH2FLgsTeMzS+5uwE8RichbxcBdmmFqbPq7eF38doXT08QDcW2A5FpvxaF6+fxldm6uldDSHQPP
wXAqJCLLX8pUu4sFWbEBvFSZdEGHe4f8AmHmJ5aCxNufl/bUsDNsbDu8w6DPbM5jG7WdhBG27+ql
p3o+zjg3FuKtJfRX7XaS9xdvGGKjennCBWHC3D/1m9sIdyU8oPMFfF7IxYKQXBZ2ZGQBK3sSqz+2
iRof3oqzwhUp6TQ+X+V1Z6rDG9/FDg9icBykmvQuh51xSoLCk7aJj6oOllrpxGcVs00z3Vb/UPae
wBnCUCdXeY5R07AodaQjVTzCL9zKoWYSFS40MsAxR1wmhhUe7/FABfGlAR3tb0AAfJIr54u7n8X+
c5hHcfxDV6AdrwAK4AH9XmA6p9Az4L50K8edDug20RDYlo+gE9VesuLM6XQM9pTFEEEmCQIBVc1d
Q0WMxxLtDSd0Gg8vR5JDLsJbFqdWRz6DNpp+MjBkvkuBvx9lCNyx3EwRK12/5oOM6qx7F+wl1j2A
sJ1jtvXJmE62nzD1xcHTbSd5rSBZWs5LAxi5orCG2CCyzZxrnTTptQWwniFKke9kNTtzk+A1+YeS
vEWzPe5eYCgZ2RVEPQjz078m9dDjy5U3aXeX9Ngeao6KXpBFbzWRodCf2TN/LLvW0RHnOIq0iAPa
/uqu2c+DCaG5MbP+2l5bWVgF3xvR/W448Juoe0fnbFo99+h143mqChQeQUnrIgQzQiP+x8CjnbvY
WmiU3MJquQT8maPVGP+Oy81CwBxMcbpUPT5nd8uR4gKzUG/mnXoJTiRzaP5CMQpAddvaBQqH9XKM
aH45Ue4tw5xcUJM+1aWIL3KwG99mzzGYgll6jgH87QFHYjuH6RksOvgtSlfNlIm05kXVNWSSXm6X
9Fhiptn6yLX53Uq82H5ceEczNDC08FE7XIu9kAz07/achIwQxUB+wMNaUFHzovfXXmXdEqD39vRg
MTUDMVr9MhD0y6AXcNk6I9QH/+uSsZC+P9oxVgfKsph37Nu3pcaxnLmRLSdRRTBAJfrl7IqLsQ4d
1ex4gMdORFA2w40IiK8mHascM+1VZ93A/HUC4LxCkEWV3Gc2XDeh6CT3plwbJdQ57DW7rcaRooa2
iXHAYnC9IvAEKi2z6D6DopAoFBGObE6Rju0j/zaVrMMBomZK/QbdA+F197hD65JTnTR4WuHvNrTW
/Ye5048LV96JjM7Eqp8I0xLgCaEYck+/yLn3LsJbKfOGmbZprM2OkeeIqzDGzqXaWMM5aDhFLS/Z
xilQcnB6xjEtnd/LRyElDb5NGe/BKVjxCv1t/bM7OykkuDC2RVMG5NUpoE/g3DVeebMfUh3ArVL/
OURdqOYD2DYKjbjmTi26FWP8Ljb3z1Gtz//BGcI5uzLR5VumUAsuRdN9Dn6PnDZ9mMHDLvjjqZN9
t4zWA+JORjHsBlJBezJp/fXS9KQKPpAkNHvqa0pDZyCWm0PUYUCrfjFxV4o78az6Mn8hOljck/MX
KLeYTOjmdTN0rP9YGTKaCMuevRjoweesw8D1lJmfkj2fv965WJcIqIGpAihbOFACNpKeLEQUPQo7
j2fifDTvwoFR3JosmgFY5UvPE8Fpt0+Or5cCvbyS8r6Ovd14hQKknc3gLH0bNeyATvMMEZidvqRn
oExNgdfxMl+aBalXTl0SgKZ/JE9M2f45IO4y78RJTmwjlSqo65+qCaLZxggp2to2fGx9ZxY/Q2qj
E7Fccmjf5K8YVL3Ebyf4S3KRB0D//UbiREMxTITFjG8PCjjOi/deGwMpM1olOTx+09efFQaiwmb7
T9qqMbY2G8PCnAAkLt3awadnJoAlv6wQLR4WldpYh0seb7FZILEm0KJnAAb37hnYyiA3xNsuQ78L
CMHDUFVgAa5I8PmFWKQg9jV2ObF5h+Mm9ZS91wc2IkVUK4BR/tU0Wpa6//lVzDZdxtSw9NkNECKk
Wx/taoQ3snXDJvnasgw31TvQWRdRtDCh2Ww3/gtEXaN6HDYd0pl8QNuvI1ztbw23jpr3zK0Z5QHS
bduXOPpFjFLUgCdTiWLkfv9AQF6KoZBU8hlVu5llW+KD2+LbH6Xs1GJKpXtmCE5ndAVENSrDMn3Q
NGXPfnnaEdOkXQPOCHQOcGBFAm4cErISK3wiZYTnPs18YqfAosWJKrRNjecqj9mFTemMISmSqLia
oKq35QoAZNa4CyXZRNuqfV5JhdyPbjGe1QAwUf4C8KmXsFczPOO72II4vmm5JgPiVStduYrph0PE
vcv1izXCTbNR8BPPW5XwOvPXgQIZUb6uuEE6Mm6moGPWnnqSZjQQknK6rAkRGCj5c3Z8ww2zXNsa
/1UDiBiEjz0BGSt+svF3cIywmQo8sjL9Z9bM1B4wmzaOCi8Lkh8evrIKLwXzzTNVoisOWpgxYOxY
bDi79OwfjFc5OT+fYsXT2Zfj0EGLR7/6PixBbsTsDFuO+0OLYtvMfuPlTYAfIYeu6sRXn6rMkrQa
odRowjs84dxN5G2YgURuj88lZnRQTvmI10XQHycFwTiJX6JF9Z00RL3qOkolBVckQA3y8mcuiSHy
zkAAz448fyA/l1lAsESip9vcyLXOidiWKcr8WqX0mMmlc9uyPNUS4hKo8uNYoHQPCnPBZh6yQY0u
PH9OvNmCaIh99JLRLKKV290OjbzQAZIp6Px6UpBT/0Mt5XTae88dGU6w6uK5KXXOgJvUasz9iXsQ
KWRf6AcVTqlEqQhSE0RXZPL01x/Yv5E/5+jThtOipxGhzS04Ent9ePW2JVyRJ0jH8O4CS/j23R5v
NQwB/Iw0xiPm9LQP8HpRP/HiD+hpn5FiPQeXsxv9dldgQNe1YWtZcZvGfl53h+ZIWyBNLEAx+t9N
B/Y48hHr3Cmrqpqz5FR0OOlXdAzMF/ieSKhbSy7/Nlg78iJ9cBWfCyjZR+3mqO5koX3uOUXWQSKb
h05daA8Fulzr0nObN2unT+UNXKYkrCHskvzefzGuWZDjRosMUADJ4TooVDFO4HCaROO/CCOwxwwO
PUVyNSaY+Y9CBnbXBvsZtVGJGcCb1Ah1B88KKRr8aBHHeSrGrkwouseNPO+Nvnr0puz7u+yzs63D
rHzpoCghEopuH/YReF3oUrLsI3RmJyC3U1G/jAZ5FHCIFDUOj4FMTLve+Y0/V19xjKUcwmGtmt4H
57CrXtmvv1BNyAYJR5BqbjfR5IMjCOoZ8k/DWdO2NyggSHPQoWO/XacuurtAyCLiaq4uRb6nCbzI
zWNX13nD5XMbsbsviN2nLmtmOrCISBENzVhAu6noemaBsMmWKz+YWIxx29l/XGJnz3V4i/p6QKcU
LvfKPjfyJavAYvxs38j+24s6Wu7pbPXQhR2a2eRNxxZGnsA82Kou1KLxxj/03zguxWxvBnExVnkr
hYv3Qr1SPl3+fRFGPdnzo6amC00JBfXY+xguAv/shMXAYpX0xJ8zRtoeSoYZkYwfGSTDum4Tx6Wk
lmTFknB4NKE/YFqePCVyERkHZVDEuWMbqrdtFhvdaSf3WBkYNi5+DrtjO11JiakhxPbiVO0TYQF3
Q3/dWdGMPFNMhmUwaBBjc18Pmomj9STjLwqfQevErLJT3SGfLKTR1vKH2RMl6S5OxfaQpvcSjibZ
RWj9I6eFyfc7VjBnC782KOvm/4nuxmHuzdU1Uk0WXglzEi3vYgfS+obu4/uW0OZX8fT5/+DMud6K
K+jrdXJVgbSfw3bjQ2D40btnoNdPG5rsGn9MFwFikRRVxW35JsavykzqdGaR+H15yfcJQUW2X6Ck
85NcMiNNUqIp/gRSn7GGqCCYExX+7rTIH7aHvm+SQhxKpgFB88Li+ohR47hZUKgkTeC+KfzD2D32
3MTulxzVd47i2QgqFq1vP6BgvOdP6wqzYpuKH4pGEmCJJw+o4q1FAmwaFcDA4z6rCxQleZNU/W3e
/7XPi4DNfURWqmMSylO+H9tfB1IecjkhCXVk1DMsxRqE9qOzKhGRUSQrUhsBGXMYpLGp6Gxv9xK5
CBySXCSciuU5AEyQvCM7UWMiTwQ4vM7MELIvNqoi8NH7QV6bQpD0I9Z1DnwK8tOGdX230PRq+EGS
+ECcO30XEoFytZk+QYogs0srLem9chTyQK0h4bZJAz2v1oitBr91RiBXmUlUzBFmDka6AZzum65v
tf/P1e9bX9+o5o0ZI+W4BQplY+PTLFGKWH3d7FZsCqSh5/kjwgqPJpMCMcN+NU3Hcq7vS6j0HarG
bjS/ChGhwQowy1K3Zc4v+dp1j04URtI15UE0GKCq0KM+ksA0H4HqRQXHkNqNdk6iO/r4R7p4Ah8R
s+8zF95h0ihGUyyLv4E5ZMqd7jaZQ39MRW+tHH3mw0S7tN9Xj7ytCvLRfxbVAdiolh+5MpR8cU2a
LeeIljnCRE+xuUe5Vvb2ZXMWetUZl/3vb3q7ZVHbWAGiAWBSCqYuU7Hb2qvEqlUrimxktkPOrli9
KV0V35OgpitZXS1Mc68g7KirJv0xjqhbs1Y+Qoh9SDbmGAqFgIz4oUnPT8Mjib4WOGAEZnA0l8LR
2MCM0ZGSI73iQ4wPfaqVK5OBfQ3jHs1sL1vLBiIUPjt7ZkuDg2UR30ezGNcqhDZHaBGEsvV+zJBw
rwiIZ92VMpcYHpWdYY4FrYo78SmyGWBFbeMnJI497DAd6HytOSklmwRKX2qlL2jTjTR6DsZfqpcE
7n8aWe8DFcU3BpFx3ijCI/wo0yCDXFfOJPawUdVj2CgUkhYSmZitv/P6Dal5ZPj5ACIk89beexOf
SGKhE5+L+uoGwceeHZdWRSajETBQAxOsnMWE/XegdUN0Jq0qJEib6MK5r7E5TIpxOo8pEdvCHeLA
QTOSh8og956MF5b6EllS+yJHF3rZ3P3BO2D91KWdqdwTU5KBiHFjsvPf+BFsDKG58jIur8RDO+66
NeQiFqL28EwwkT1G1imtda5ivqEhj2vBYIteWyk3BtuTKam/G04XR2HeVulxO4aPW+B+h98RVcFd
CNAw0kYyFEOFwjvO3hh2YU8oGXCzbcDtaIZLfpl4vHOYl7ejVav0+eibrATZ9XcigvW23PSkWunL
tOoQkrhOfe1b/AiGg0Pvdy/vU+tAF0TIE4ogs6tc4/yi7Ui38m/fS+8s1CfwOjNplX6xYBp/7eA5
xQdboLkOkt0Lx/hxznUsYK2sHQkN+IHDDw+F04NfOFZ8tcJCOUmkQCzzoQS2+TveiKt0T1rhQ53U
Jo0A6jEmkkUgtYcvnkOagiKKABJAbfuZIqHE74PubqiGahFfCbNgqyfBWAgXzVIyeRGSk+wn+ZA0
6oCshgVVuO5hC6VFsu5j9uJLeiel76ayliuF5hnU9JZmkb/HBNH9ZKZ6qFPTlUvRGc04gl2yUnvN
iccVctQcv2JXFp4aIzeTqfNxqOzJJJIJld28oiQ0GCx/Ns1CW72OYumHI7N3ibT4oQAecTLM6FbW
bnk77Xr4v5i02i/s0lN/YedHPV333J7mSvSnMg/KC2pOIw/vQ5jZybhyVBdGwIVCtWU0480TyBrz
gqGE2IrybqFi34Pn4POf/1kgB0Re6Xar2qkOPzR9yv06rQHrcbpXraX7MUNvbtZI9W64G78ZHj87
/hjZDODCvn3qdmMXT+oL4jVvsuheJazt2tddJlAQrg4FbfEHSDb2GeseIBL/BuSjIjCnT3/1L5Bl
Ga7VBEhucu+fiVHWTioXzDIwkmjK48drLTY/MSIzgJnKbYTjdQz8N4cQI0JsMp/wlxiegH5KyBwo
BPjUigKXEIOQp+KdgrnDlN7JFcn2HWIdxnyM9zTnTNi/KHUhThbUM1rIXUjp2mhwC0H3RxGednBc
9A456Sv5blbGioNe4Tn8SnLU3KRnXtBHsVd6gcdomIwIjCSr0PnPDLpXAHDrqfdJInNuZQqtJVAK
Kr4GcC7LzVQooOv08cwxjDzTuyBTQ8gJe+Nu+Z2rOpT3rpZSNxtdQGDtfx/RXyJ49VrxFMJxX0Oz
YxxcBqDwhRKHyKvyoBa+FNrspvCSd3l1qjE/QcnQuK6m9m4b/5udtWlSB4ZYHITi2jH32TaCGpJP
nfVjNhAE6acm6g3q1edqwnrPji6YVeaKSjbsvOeXlgTe/Mf1A1L+ryhF2oZunU5lxDPHb9PWqNos
TU3N9bCN4aFC25NfWOG0YqRB4wqWNE0XFrMawtCW37O0gFukP0Cejw4wiS0xd4Qby4n9QH8RwuUF
bucp8uhsd5YYlklZCtZcCH0UpQvgIoSu+HA/lxvmooHsGdp90ae49cugTOmy35mAw4feqW4FQvXJ
P5P8pFx7yp8bnlaHMD6tBo1A/1WCzjN4WMz2R4KnEQV8PqJvz09r93Se2Lmhr5A8AZZUAWyEvDEB
QBf8B8Rd81TE3vKQdhpp0eEKnRjp6A2w4xdbeVo9VPJ+Gyvny83ZsNQ1AYPDxPEOivMFovHG1SGA
ogWyGTRGDv3fYdhq/AeKFRAKTp3rtJ/Y7gGq+rDzzcv8BG8kvK3n3qsqXcu2O/P5c4UHyXyZfOA6
t3KGryAM6LEzJgt15GYypIJn/AGddRZS/KMPfhcnPmc2AG0q+LvQ+rsY4HBUloME7aYMFiTwmzNt
ALpR+sJKX5Z402E6yX3gi6013gN8DUd/9pV/dHdZsi66sSFyrv9iM2NK+j9MLOaYB+Y1SXlTtyKy
xosqmVOzZGCOeZxrnE9QC5NaeXoNOj9j1CLZ0kI7QKprrKQWWNZLs5skB+F5JOcICE5TSBdYNnTa
KtB63vRXhFp4KCAJ0qtm26oH/F+BmxeVwnQSyjwnSp7XIqiKmnX+1sucXKu+u73joArJp9WNzmu+
CRo1tp0U4QDEQ7dzfr+85MqH+JbrvPfcrYFUA+UCKY4i6QxAhKPqZwhxJ2shxJ6+GKXJg/HQDERI
tGK0gA+FUGp+T+jBzb87lOKiFjE4ZTjG3KL05+fpCjA3HKTq0YvQjtadP6dc0gYrAxKKq97xkBEZ
onvtazJOrr64nNoJIHPpZiee4PiK1VuE80uGU+pJcvFeS6lLUi1OdGMzyF7ALpZhNA+YYl7p0g+X
UNEr919MED8JRiPBUXK1AscG7mMmqdZdrP3xQ5hyHgDcm2zfQwGnTuXbPjBHBQv4cgs0rls2itew
WEtzALwI9Bqyut9F11flblCUmE9XuqzsSmTeS6pIoASh/6ZMUdlLFlw1WGBbPfujpuCF9dMK/Jfw
XB6BZf0N/7Wa1iTU7/21dKxKK/2FiyE/MPpSAxpquJQnbf/zNVay51AcR/oK6KNNswyXEnzUtjHd
QHiGGZl7otQcKmpNfwUHJOfqCAXc+msyBpvKssILqb4sf4/V8iiTcukrsWMJj4m9+x/wYFe3t19w
xXB11/QolBtgQTFDe52ahUuw2OCG2z1Eo5hosdcTqbs847PuB+Tzx5FEgFjmnCqnZBKApxUP8eJ0
tuRdAuWwZMhRHpB7IhjLeRbdw0Scz+kDO7B3iuDx+/253YZzLDeNVmXxueMcenllgwu+JahNhdFj
uqh61VE7sb7G/ir0JE4iprRiRwZ5oSLH0Fx7ciX0NkHkN/8+wfTwy9tglvAWMM97PtavbqlA1cPs
OAYHBd8p+cYIHKQy8YvhVVHr61TXdit1/4Rbg2tGYoxNNfstZ/ZXsnbJy7uTqzgMkEXwcWCvqgby
eEPsgYH7MYCH+rkOq+nIu4dq/scoS6pygVNHEZHZS3z5Pbc9qHrbCcTZlT4WJ87ASdxdphHFUX0j
ZcA19ZWWXkoCfIhTUD8Ang4m9/+YNUGPvOGQPWzHRV5dWscMtwT50pJHQD/2iC00b2oE3SRJRhRP
c/WYGot5DiyNcivJgjnS0PDyccx+w1eywiUmk5Hvmuj0c9kWlBCabPCEwbQAnJSBfYGNRZbkBF+V
mRKXrTOJTIK6EeeeYTC00+GW86WE5rurGl2t8eu7sD73mRgpULUSdT0gD7JOV8YrHHO7bWp+JBr7
8ZUQhjJ2swoAEhO/WTh0kmCfnsjT71XDxUnfDTKX+Qou8iQhdKmNyitquMLqmH/5Jij397ltMvJz
Fgqf0FRj/4ledivzpXMWrfSOtO1U9v1EFhuS9RW/CO+xvUQmZJiMTbLW8LmRSRZ4m6vFIjNulld8
Zg/Tt2hXSnox6DYHvD30YOFpJkB0nwlKmaUR7oTBaFFJgzOm+pgVngAG7v+DYqlhT2EIpieYr3Fe
2fx/+YdW6u55tMblFUxWlOFiT/Ga1ZR5DVzfBRjKcnqhwV3GNKgpc06PrlU4C97vFpRnG/mqgPK8
0bonlhjZYwrYpsDvnT8q8RhyhVmSRhzg8vLjuux/rw0tC82h/OmS3uogL3eapnKame6cI2oB3iZO
oliz29Q/owefp1Mqc4W+ADoai3Hz+8/No96DkIR/HNJTeiO6Ax3cuEluJWBnYoRP7b5dGMUNY/OM
iAznxZhY/14oTuv8rk2Uoy+oQC4+AZ80zWqmhYkwa1S0dVlHzeGOaB1+l3+HGBjVKAyj0OWkSF9v
cSJKmAVn4pJdhTuSS5nGJn2QR4pUb0VzFti4oxfN0aXFfGB0pH3ruUBOGENnDwVykXKfWNsyk+NY
xMqDIOjmKlsKCogWx2/0JIB+8M8xQuXzIJfF0nRPdBnFp54Y+eLX+5YZ/3QjMVIESCblgBGXAm3z
sgaQNLcdMx5cCoun4KC2S9zX4MjjVLcHiL5X1SJauuy4Opnmh1CVLu5uL85XeW1GB3ieG8UObKBm
Jx49S2HRau5Xa6h/2RqpeDBnOW+NrOlkt0dQMkvoxEuRysRPs4U0PgDWx/aG0PvDzAiZDPXEXW4A
R+95nc7Iyn/u0hautV5SGsJcG/kKfz3WO/S4HW2VuUZ8FvTBvU37X8QWW2mw8arePVWrB3CTxprP
9bM2gg5fReCdFt4a1eBWuwwEZX+Tp3PY9szX1e8Wf9VWm17RxIjyIW+yALDw6uukq/iqBc+O5LYb
MAfP205szzi9uXKeR1NA7ghdU4FTH5JE9E+jz1frbUrhVDAvkY7HHWbNFG5FQN75G+3Moe/hoJ1g
tfFhwgN+Yd4+GmIkgthPX/QuvRlKUiHEvmyKqcMszOqLbyA16iVK8r1D7W8bVs5keGSZYsNK5A1b
kkapqQAe54EjPattEI5rtht9OsxLR0hWUjBC+BH8Gn1BJNk/IYoynzUIVDtT8vaJrIgFjSGJZRT6
3rBIP/BJecNxjefpdQSINDgN0orghVHjzdUDwM7kqfcdJZy594OcNjFQINYav1zC/TbpVVcPtqTo
tLl5pyTD1WL5n6i8WKqYPgbCAfhU6rB3AEAn9U/WtpaW5b/++ueSUIXSFKaJTJE2Yotr52viJI9i
c8KB2x2h9VsZKtxXLJWhY1GVboAe7fMZsZa74Q2bVpI4Ib/PuXWS/iS8fHbpeBzOTrU0yudcyI7a
TIWNzWBRav1Dz1utYvUUEOtYE6xKFN4lJtNaxT1HTCVYWkq44OcbWfwju/sfBPu1dgiJBnrTamDv
ZXgBImKnJeJwWU4GVJKx2maCSLUcuPVgU1XwlJGSp1wOhU2g2IeeVVlpX3XeGqHkAX9dufqlsWPW
s47yaodTv1og3dSCYzyq654Js/vv5xnmpGVf4lEJX2fW86oMAqlUS0pWD2Cxs4IBxYUAqCf07gqi
CthakfmuZrStKLRBu8gCmuyaqdndQM9IehRVIKTKdmUBJVrDHarHNo6eBUMos+65elSkkcAuK2KN
A0iTJU3h8cGqhazQrfme3gSb3RwJ5Ky4hqVzRIBmEq6t9nMy18YRsTtIDRR6AlutD0Uwz/u60IGp
LYbhbHvFHLXon7F9ZCSuDdHRUnVQVtGOI62s1eDqu9lFoorwMN0XEAF5xJ3hAPdgP0JZHXxlTA3Q
UzdcgS10dNgC6lIp8eoDrZeElL6gX0vLE/A+12cFHm+gaW/88wAbY9xRqZrRUzZY6N2C2X9QdzFf
yMvDNv0p3Paj+kyZ/LPJUF71wdzGszi/0F40ePysFgINFpOrSUctx1GRjtHT/tybTjkGKV2iCudB
W63NRinsh6KkFsTXqd0CFgyFmC2MVNvx51TMMSHqB80ze6S8++E5rEHcDMiEW4yyPe9tmYTY6U5a
y6H+B8YjnQjOBcYCFJHcKIvVJjDrno/7fYKhRhDPB9PDSDMg+cMQ+Bt+xlwX3pEw6jLYoa7cg07u
kCBi2iezKbKndWPdFg0vj4wYckbjXWfRbecBShBQ3hpEU5KyfBOr276Nrny9iZf0VQd3tio7paLH
KkZ3J+RCf87Q5h1YLwIygPoSq4ieTjPolVGh6hRaYf59AJI1dMmB4oTTHSGYMk18dXx6yWYAql4q
7Z0B0UWk1yyw51hagvklzcW5C2yxgmQ8gzN7jO+hpOL1XiMSHnyNr5dCHR7Ljdze+6WymZ/nJEgv
pZ+CAkr7nSDZVHFoWweZmV49AehcXY10i18PlyIbwjXl6BYXfYO66ALyl2Um9AmWcOuhnHqqjpMX
Y+Z06g8tJBmCEo+x09YK2coFbvz7b49Qm/16uzZQsVKMNckMcAJEdmQ1MenzNZKZ10J+6XGeT/oL
Iq7FbRKeo+1v5EDOZz9Nd7hzXGURa7+1KgEd2IPaP8fVqNaAENCGk6LBWWrO0HisX3zyZHB8WUN3
oHNSIDgOPMLqPXCSwCr4xyHdCgZ/sjMGmRQ0vgLf1aNn+qadSIM+MgcXtVk9YjBz5oHNJdAynFvQ
gjF6yJ8uESsNz78ksJCf2fbp/nmJlfvDR6oNuMSaqZ196rGraBCTSUGx/OQsDPsvPGtKDjW0N0Ms
HFuHjUQewfMN84V4LpYUb4RaiXilIRBf6lNTr9Uua8N455yzuCiMz3etnwy5KGgWxH0o2cWyabzc
WwSw6n14ezsrVfQJcrJUNa9ZLRcD4KSxwAVOsgEz3j8/LYUGcPZGHeOHVWpI35tbEI6YdPHVPBcI
nvlMM+1IJL/GOZKkAQYIH4vMlCoodXjVllUprdzmCQ7g7sJlOYfbMx/FnyPWMA30v6MgrjIF4lvc
+ra90tYlpi86nC9ugKSkjstUuOS7lyMx619PjwicXF/7kOsi2S/8ZPvo3JLhcSPddISz/CSijFF9
b5Ynx8ZnTpSmH+qfNsaAyhAW2Ml7p0ZYTt9XTj9TzuYPLA+/4Y8Mc5l5TnXvTnU/jcNMi2MDVxKl
Gdjh4h4rdm/l7lyleKs4k9MI3jfrCqngBWfluUOiZPOn2otkpejx0tQMW5ZSqGzQXLP6E3eiYPJ7
4hXpUMU35HEMeSAKwOL+tS6f+nsz/lHrlQBTm8ADsrdDpYIjLJNBHLZGr0FDDkkTwEq0DK/525NZ
gU8c8R2jNr73y9Ed3/L3JQqmXv9MjJdictp8HGDTGabSciezrzPlW41P3CZ7w5ZC6ANwsl7miDSq
cO7XjPPivZ0TkfGP4oy0J6tXJXLjxTEkDod3brWcOpdm+D8Mcc5FZtGYtfnlXkpLSzYCV5+DBcAX
sC7x+nmlwWFX7efaQk9bW0MBdlLg9fBexXrdq4LhYP26iBCEn4p4O0wSaoUEBLozC4YPTB/tc3vR
JCT2zVeyaXeC/Y/VxSUqwuG5GDBFYWV58saTVHxlqQLl4BbM1hM99m9MsUwb8R4xcW0YXbymFwwB
RcdrtQArPxyvn5fi0Ea8RfloQW8prdLh8qLgHHB0Rl0fARGsaqoIVNZxz5u6pwFqFSoKGNYR4YEd
sfyjAIzdXLf/gEQ4xCs1LyIT9mTU3GY+cn3+U2P7R/MvPj+yy4DkHfuhxtKtJIhaeYm+gnCreyHd
4+Nu7TviIASeaMPelvdY7XQuKPdHAgHSgtmMi7ahp/tiUT8L68uymzPodjHgrVXizebRZZdYGXlb
v46qHutAv6xN8dY5dj9NWUWP21MsNulcyy1hGQ+OefEB8VX3eVCqAmbGOc7th0yGVfra1EdS06Vg
1nHwhlanMA0ldvUkhNy7T4s7vpUPZQtP9WT5fxN22qSgHYOebSxxn4Gi5s0SZYOVHefVr2YYE2Uq
lvsXR6zJbzI62HYQzT1dE6vnDBExeFiw6cxxF+deg/zJIRnBcqVKxzVWs5VxMgJKsUyrSN2HBZ6S
D/gPiLDf1gu8FoxZF5dZqniiFw/KdzPTY1+fRWLimfKvCcFrvKNAU2PrPjBYLpEY8q1K6FtLvWor
IpW1RMLXZL17GnTFIoY+/BOYfUjYxeF2Gg6g7i0syVPqmD9VNk85StmEpOLFr3OWaEdetHhDyOcP
ofh4GcsTEjGAffd8barNP6TmTHSR2wP5pL1NNgBqil/HKeYoEt1fldNnKD7F2PTQH1HAdmiihqMC
rS1XjWae7JSe/Ipt5uLgt6Cs19fYTGzvII95Wd1aC/tuViSlofqiFQ+4LEgNuN3xwUPZ12r+hqsr
iAbEPlX0JoxTG4Wkt3J23e4wtJvpbjfPI9yWzW7EjjbdhWXppSo20T1FRGzTjguSTrBwGix1Ultz
i4UhZB68lIc+LBVjwQkUoXRre6qbxdOmnPSQHTO28OlNGBNv/RHSvVeohJT+tXdazNDHwYS7/UQ1
WGgmbCqTpaZZPrHdPulmWvNFezYUIJt6IsKxileEx4t5KcU7wftCLzPbOfHgJnE6H9oHgTkNmFEG
DdfddqDvo73N9nrVQPiJTL0xWqFg/bKZ6VUp+49Bo6YRGVCMpQrn0YayjCnpZz/I1U/2j5Ax+fdQ
Ziz4xmJV0vd145QdviiLXrevnpJpcJNBlJGM6zq65AEvL+SvIjRePI6UT7oHA9up7czXkAYLdQJq
YBFq3OV/41sAr+XgDYzDcRdD2kWlL+E7GMlXgQk5El4ih3k9ZO7tzwV7HilENlJeAK/sFxeGTIlz
nowZfcyaJ/jPlMrpoKEUW2ySeTf0iaYNzfoc1sFxbkP3Smy7JkAYgj5kj0Aec57vE+DsCufN2g97
J0H2HK2gSZ/NIudHbdm2+O2OzOSiPYlmbwcfccVD4EhHMnKfSGx6cmMFAWHahMfabjqRen9XWZgx
e8In5sOu/l7jmme8diTAirOA/Pt7jPJSk3z421FjEKLzyTA6ucc/j664k0eG4KhqEg7i2vY7mxWS
8i+VCshnha8sGWyDWaoF0WHChop9WOopIKR1XYmHwnBt7lpOlOnBgboaKzqMKwo0c/+a502wY9/X
/lTAfZAFrCP1Q//nzd5MHx2f3MqcoOr2J9zZT0Y6Xk5IHa/6CgqguFqKBt7rKsAd1k3q8MtZS7mL
pCxRJh6ADEyZVOP1q11TOcZzaW4mzEDP2g01jom3FRV2Sa60X5pvjzjuuK6gd36vJDowuZlSFIp+
IOu/hSryHDIiKPzyDWQeDzZyZlA6N8cli7M23rjGmZ4QkTP5WKCAZlJZKGUrT+mLXVj6oc/ptVzp
8M7hLtVh60wt6TTtd8NVQyOV2MaBvBorihnwhAOYKVC7sOPjtvJxe96U3IheX2VUEvnaryXgJYb3
2qy8cTrp5fKVyL5VJ/U9cFGrdO2cRIxysiLOUsUXlUOO9A4ZYEU4JYRwd0KJVephEyEPYToDBsol
2IxKKXWPM+1yRirTTZZDdYgS6AD8MGiSCZ+NfVA5cSJOi6yKDmm1REMA3uTcQ2H/vIT0fRYJ/esW
ERWD9rFCnFAnCVLJYMglRQw7+LruMm9Pli2cFdX9RcozrUSishPRxUrJcritjlcgcUcls65QiAYj
6UY4uFgZZgSwh/dzqshxrGYQTpZOtojNtcciQZ3/EWqXwiZD7C4KQ9ZsxweuTOjhihlDN3VimcKe
tpKSYGxntH/S7d9l6p9HVQm2UZl99uMoBPy3Dk7zry4YdbvVkbf5YRmiafk5Cb/XPh1Kx6Aglc/m
xPifPp2s9Waz6UOLlR6tl8+mF9XsNUk6fSJRKPySPKcxXrMb/nt7lucU1oL+S5VecqkxQ2PiMMLr
8+QEZ9VFPV6vYKRJABb/VCoIuwEs/xj/MP2XER5KmkMjNwXHmj3JWr5CXpVKnlTV9Be1JetIaSiG
5Kv/pBPbbluVmc+X/833oWUbtFnpENiD/HFHYsimeixq5ZCSLSgTzBYjBgXLEHwuwrC86u6RfXXq
+vgJzMDDbjfHB3mjvYYkU6lCV637Rlh8BnhRQzih98ygG5ym6A9NSiLIA/nc0LHlhgySJ3fnJFkr
ZlQIsSEUstrhnY49f4gMGG8aBwxi+XlZqrd+2bLYO7V09xS35/Qenjj8rU2I0FYhNeLpQmmMy9Lg
Dg7YHorCdSgg2LZ2st5b1z/zsEUnEU4mm5SCSq3lbkIonYG5zllGl1YG/c2a7Z7AHPRQ1oy8s0Cf
CaHAy7Ar/FCF5K54JOdnGP26SfVACGvIyt7cEGt+sVPB6Eg1qwxDQTIgN+vg6vXZzaxx15N5djyf
D4KWqmT+18vrCgZECwP8IrB0M7G0xxcxL1ITNmM8yZckQsf+1ZPoKfUI07vqSJUCrDMqHVGJrBrP
b0HT+3JgDULHwR9SRTpbQFtLRLIsF+FZf8wM4rFvlVkOmWYpdKnfywgnTW4Ayz26NX+djMVPxJJE
ie8nW9WVUhnkQOaiyIj+E4dVvH82OWd305AqtG2+RyjOkjldly4NBLvvQviYb7uRm7SUJVbT3YMk
VJDoyAAVcpNsL0nv19THC9FAharM228wgML0s6o0YRa4UimQcTvf8M2PK5x2DMnaoowmAga7l6+/
vE6q0KtGRgTt8EYb1smYdCgLUjv9Y6AmR++MI+7zgx8wTaHOIy09CE560pUWHtTwEwsfmAoyukI6
4AVe8aIHgDOWwu+ZRzZKeltu6HfO4MnJcxvEhHhCxfTlUnVTj65xYTtj/6gfGdXtK8OBP7//twxY
RzeBaAy5giX61pezkPYs3nHwZCAssGNEaRSHGn27EQN1HCOQFPyt3OH2yQvS1p74KYUBHF8/NMls
9fJUa8vRIc5U6YZV+h/+VW7RpqU8DhNL+q7wQdu7coWiHfiQFEEK2Q0jhXjT+IZ0jgFFqwftCdTb
wnEfP1j8dMCsyfCr7Y9LvCl4ERrIg4akJ3wcNvGXImNQXQ0CGIOHpUIvwrcFCs9ilSFaMPmA0Vxs
FQ/CjEpaGC4PdBw/hyQ4Hyqw0LOfb1jxvdoPjqztR5mBSmhERtoYfuQjAhMdbsGoEd7f1GEOVBAA
vXSLuSmu3Rbm/OnMkrI78kc0TZaL/ouYzYC15vBuVcZtwEeePVUGa+Dtpjls52Bj/Npbb6N1ALuo
mF4AApBebfzQs5ynYFjLdtZCHSROdo3fIGMtQqjfVAY1PNwZc4Ws8vmrZah9AG2Zo3XTNiDTRnzh
Y+WpErS0/GxyydghpamNudmncGKS8SzRIsGx0Pn01aqCzlBcCqjkCJp/Jt3APYR7s1nedU+47WBP
9XRecdvNNYPeY2QQQY2GDDVmoyDrBTpPAlb0oVNDgAGgHlP0vtvlZ06B3OKiGHxXaQIe4w/CFTYw
aYxOgLwNdTjyI8GvN9yLndrn1AmH2E0gTBdGHJ5FhpNpR8c9SRK2LIa6CCRq8G3ri/ZkgdrvC/Q8
e7ZGjL8AjyO8aMIFWSQw0X/xxRoaTIlZejgRtrbXvuhkvikwKEtGrcN0n3l8eZXilrXvy5FSeq1r
uhAxafxk92hDIPasQ3ss1b/RyYze+c5gDIj4q8dGak9NL4/QewWBVzcVcs8CJeoGgo7rKTGP9Q5u
zQ+tv45UbOKoVNHuRMrc/Q3UCcT25K/d3yU+hgh0n7xZ8d1TM9YfTiV0sAzPXggzmWCTdEfJCF9n
++pyUx2lplyBQ5yjRb2aS7PXi5hnVeiKCl+7U2AkBab2WdmCSY5Yq37SqUzH/+YUTSChkDRgbNYJ
L7CiUrs/vtmcLFVI7ph/xt/Bp5baEWIPvHgTKn8fJUOHTaLqzN+TPmgN7/t1OsaQrMYner+UgrU/
OojarhxhIOA61AzBTrIVbQdcBdhbv1ooA/ZSZTynseOtm7i8x57z1jfRWsCSeHOJcvXUsF5HKMaq
vmKV/f7zoCCBeu+m0rIs9oPeZRFLWLSnDn0+s9JKIOPg/FfayntebhBbqv5I9DBnoS1vw1kwHFN0
d+obatPEGDPOnGqSDPmxNTXw1L+6MK28DESeRwoVBhgaORgaQ3VMzhm/Ud8al9KVnpja+rxxqdNE
2m9sZG6WRKNwSjNZnGP6MY5HXnRoqa8ORJFpIXlxGjOSYtx+PFl95dVX36wEYsL9EMaEPCtx11W/
rXXjEwa54s6hU9E8XByjVHRP8ruw56RNycv+5Lhez+uvWEUl3umVEGyxUPMYd/E8G39W+ppNP1Un
gkB6SpA3ccwRO2OTf6WAfo9juomRMLKSkNd/Mi+Wjl19jKgNgeDxMR8LPqNJq3SrSwXJoDH+PsnA
msU/EfL8Yq9vlIjR+0GPiT0peiQy1n5PiycoYoj/ngUb859CQwJ4RpOpr3eg9gKEt9A72+ETqaov
KuPuiztW5SmCZiHYWgXZJFuFVwd7FZve67adWjWWU4FjdD/5faXDg/m2GTnT5R+sPCm9KeDXTMv5
cVhXiwr7pCal3aE0VFA7LEnOkD0ZmZjK4M45fYLAabp3exxRPncPHZJKPPz0PNrigPjmeRSxzmdA
L8q8jicixdu+1I6cpXeVld9rMUQmoyF0ToGvWDWhqDX370ZvJ5RJnP0uWhapMNJAOCWXQkbi6c0t
JlKPVRG7xokYtaEJVG33ZplFgXv4shMWxGzP07/ACnP8ua+xtYcZarR576mwtRYOVRNmlzClxXi+
bktl5R7iOZJI+0JfOBZz6iWLata6VwR0BRT6P/Y26S2BgK1ZKTvKEKjiQDuli98WF8DhaOTDJM6R
Hvq2e2bZ3bFw/rYNLhQGTN5KWYp1Z7j0JKUFZ8046mDFFLqZGjSwh21RBQpESc3UTdqarX+9kcg2
uraWKa18+h0sY29XyvPKAqE/i9qrzTLp7IKTIUFT5fzVQG2DBFzv3UwpqlSOmnfdl+NGJ1Kdmd6f
vBB0vM/Qxkf9kKSxnjX2ZmnHy6TrRNITij1sLGzckbTwJctUzmsUKQ8WuwxIEP0dYvXliocHB5LM
l9SKsFSpVvG9vRJzF0lLL9OCjbXt4Nz8nUMvHtc9uIYWQz2GUCPcMwhQ3nXFHHZubojl+e9rfYMA
miRYNJLu1jS0JBa5JICTKxG1JgsWD9ZrbBtCVm6fS6fWYL2Cq9pi7vOax0wRatmlubP0AOPnGOyk
EI1s1Fpb4hw2Q0dHGIbdTj7T3tFeBvbnQX5TW1swkA6Ohj1tVwkO2pOcGJWPW8wg2kKk9+HyXrgn
MwkMWc5qezVy6khbq1dzVAfrcJPdCWguH31IZy8yBMjcY9pGGKUKTso+DuCnlHwH7cCa9Bi4W0gT
aGtepf7kTp58fOUYF6sCzSroY1kGer8/YYDdmR3jLy+gCnztmh/3yOjRnEsnnfxhdR8rZqbXHFMI
DGrVKODt6/sLfvS1rcBaogyJnmN/7lsvCHLrg6F13lTNWp0a5awYQ9He4GAQ4f8vELpb/ko2bW5J
AsS0rj7KYuzS2qHszvoY5sFLNC9OxvJUoD3xqNmgKlJrX44wJ8ja5/9gO/0TG/cQpjTyAesgPssr
I1BTHQgy8f8EtDqTQf09f0999fJg1bZaG8BHFNb1cuyk5vCZjRSXvyYtpS87zCCCsNTJjwIlt6Ky
u3vQqkqMmgjGrml0k3rMluOCqBxIMWmFjDKZ8tghE5CGMJr15gusSkUpJT++tI2hUGex+CX+9g66
LcwGfcZIOfbz4Djt/Yd5/QMohaXl88iHo9fTXVze/x7HlwA83v/XZwczxiB/aegt4O93rJDgHCUg
akTNkUNGPKSkU20sYV88EVt+a+6nhpgcMXBwFkD1WzIqEnRK3hLTVFdR3r4DB1gYKnZE4PcTM+ok
BtokEWtc4ZhZYJ6JvE0MuCiQcSpJjkvy0JO1xi0wEgzMax3gaLaQ8CIbxMGiuQmaWuZgdDczUCpN
Vkc7lLIx7x0KWltrRaAFWVQ1tGusY+SvRp7vmX+r/uuROoY7MAiWeFwe3MJqekO67HkozdnLkYk0
lAISnJgEtk3KmYtfhl0aQGbAK2PNW8NSS83f86RDNlhqdE3PlcRQYCyAITbgD47wJVldBmEXS1hf
erX/gBTUuT9HCEAlsHxY1+MleL0jI5QRQz+ZmdlGrNMDjYEOT4zmHuZBz9Raq8S6l4wE5vQpc+a8
xTUzu2c/B773lB1aeVfXYayhvGdP0IdtZ+Ut+VGvLUf5rJ5AbiEuYe4ySVmTRad2MwsaEaX5q/cn
xDpCnwO38zlUStMhGsgxt1d6toOhQK1rEjbd55JEsd14g6QR/QqD+los1pVGe8EzCn9sQVgdoxIY
RD7qwayIbZoI91wVZi7Q1qFAk835yqV9mCrmqA8H/hBCAn3alwZZ851HUO9CAd03Vxd17QBWzS+6
v0dqmRGUVxX0rXBOwQLxnXN6QKYdfLYrQpu722J0h1qNJVNtQhu2Dh+201ZcGKwyvVvqKCbUIvHE
8c1bgnBm8PNJL4/AZhlURUBe5L0To3el5RjGr2qkDicQAFokuoWaN2TGoVKTrFcp/uwjdpLV4EiD
t56fBkgTB9JukG0q5pYzNlFrOEoERpAddpCU7SrLn2FkesyIvi70LZQYFDYLGzWeXcQgBhY9vF1R
ZjNDjmZgTQ/VO18/or5TYlNfYLAFRx2DpoM70pbMfUILbfYdxXl4gy9XVvfblvpLga8U5c3URt8D
V/akTYsAqBPepN/yf7+O6zFsDPPayvSlkwyUZReDICW2RNRxEVhL2EJ5gI9i59I7/8m+e6a2P/zV
nG6zfJRnUflAVTHo/108nGVWs3h9ZHAjVsAt/79yZFiLn9arare5mJ/Zy/XOgvujwt3zSKNEyvb8
KZ/mFmr9NQKj/ZIJL50jHmeIjcM/jorjvE9dTsZNrUKpJdtycINoM6zuW/NmdxFEWS1Ycu91huZ8
+AC3TLIAdpzPHffFwWoLeAlih+zSeuyQRty5SwrY7aJWBc8IlZf6UhfY6eSC0ie23N6XZkOa3MFk
kYr7s9lM0shOX9d/b0WX7HxcHvVNMD8l9g+5+0nTbBkbX2QoTPd0Aoorq27d1F0ecAWn/7STvQNu
gI38q55o1gRbbQKgXdT+DZxP4eJ/tLWsXdK2DF6JpMoB+t73SEwe2OM5maZmzgvRh6SkjWIDA1dn
ac1s+6TtNhcCDWKHpv0LplHq2oWGxw9wolabJQ/1pVQGOKknZN87aoGMCZ/Gn/xzo6JUebkf6mWD
0lu9JWTayle1vOH/dudylSO2s5w0X4lGzp1KBTu4LkJ9qkztlg9bpsDWVUtNjE/FZDZ2BbbjC+/3
Hp+saSaCmc8oxer0ubLxwbVsdrkudos2Bgdlbt+GRhEOzxCXolPujfV1mYv21tTLj4Hlz+0V4aY+
lzdRY715khnYBwlD98Pq/OiRBkq8Y0yHlypaBySWT33hnA3XYdDi0afofSUEkttLgJyIShkg+8UL
y5TGJtRqAOR6/ozc1VPk5HX2o7WgeubvcG97TmSpjH5z6tAoRoAdMY4KoBsIfAR8zGTUrYG6/e/c
UWA46RGDp2yKHWdGY/+BNBWkL5ckmWAZXUUYoglWk3PEIbrdIvoqnZ0lZLDWIxCqSWHD7lQ4dYKD
1kGcnCAhTOHym55zssdh5HZSL+FCfphJRmLf5POj+1+dmo4QQmW9TSkFB0aHuyZjXNyIqtM2JEoC
gcOUQFdxaLv8S4tVGEFYWPhZkr/8UpFus/2ufMUH/WnPnimxRAnY5meIH2c3MAhZ/EVuuUoRG3kB
ICoHM0yaMu+OwZxxem0R5C+WVdZN/rcm/Rz0nLKaj86bPtsrWeYbOytOniXJpiFDfHflbgilBWFv
H2YWfvXVouybfZYONyPtN3vMLwvwU3eGyVrzAkrVYoakCC8zmMDQSKcmRnK/vHje4ZbjLdkM/Kow
Evs6jRPpUX/Hu8O6jnPgiLMN1lEb7N00qkMw0zzz5aGtNmNaUDwVn/9vSyO+xzCaQavD/lkr33w+
YZ1kYnrBaf2HnsIUMU+t+8cvaEeWpGdPVKlKpwnjGfiKEPEJWWTUrrj5I22y5oegFjsVgLh1bhlJ
RSKnPuoyhUVMua+boQ2zgl6pSsRvhTQayJtgJU0YdXfWn533P9RkpIAKpA8fV9BKn479mAGo/kCi
UNdftgETadwZkCK1x6XMSlLwC5UnPns5R6vW2ISrf6oo4dI7dC/nBZ2YXRynqVB4bHfcRCHsLh/3
Mc92Dqoi84F6V4y2ZXp7D0FJ5Cv8QfyQaoH/FYxmUuI+9x507nMiYVtezETo19bbnDHkeLQVdgDW
LZ8uBmrlBb+YRLt3iRucbqPFYjxaVMKGknoQFywT7zo3HXDChbGj96VQX0Lh8rXObXUflYSZpV98
tjX9TDyAoD9lO5+WLNaG07pLtBZtc9TnJpPKIn3CciR6tSnsoz/uBN7LOlsVao/9p98OA6Wb5eRE
rqWRnOfEhsWqdj7fI9FzKGZrzmSa6ed+4Di4fVs3DCPPRuMft/GsQkbDG0JnADjGbxHDcbwPD21o
xm6DkmhYEg74lYZ/p3jCiuuAksjE5qWng94IROLpiEjpZSYbPf1/IK4tyNcl+Ft6R6g80o2/1zfm
t+0Sirej8ljFXhmQRdq4LZh7lUDfKO+Af9m7XZ6wnQlOIIK4Y9t4lxQwTP610tEwvS1WDAbnfQ2X
5Ufl5syeVKr8mgFlkgps4nZcPY+d3TFF8jF3yXzDRDXcp4xknLormvjHn75Nn1V5HJ42HtaDF6j4
PmyT7GaPjrpEd0UKyUmipuUhJZ2e3Bj6FoAFhGXx6cqOwVnDcIsWZcZksUFZ+lpHEJeyf5/NTYdG
ptelnSeul3U1DDHF4vM08qk7T2HU4+HPxjWJkb1nLl9h5KHDUml1+ec054BlmIhpGzV43u9Jp9EW
xIvF9BOEiB/eZfDsCSskoHRSRo5AznUr8GAAFqFsgHX8V20BUOIRXrSfz6YGcsxPyOPo3qNm9wGe
cazwzGzFoONZuSblPjmL0dLIwxp/wZZFO306dkfOdrh+FsXIZ0fPYAzi5b7pWffLAcrwJNtHRar2
qrz3qb6meUzxK3qmmnGdvSQmPjSrDjEqUaQVdwBc5j9DvzNfz3T5yUhFgMPTnHW4ajiWMlPaAu6o
v0YQHZJ8EEp1qns9pgNl+URfKJN3hb0EznalpXD4KCrZnvneu9KHdAfaRQyB+cFg/kYEYcGIWSmZ
lYrBxhsNpfGn7mjUU3kLEbY8qhqW8U8fQ/aBalZyE6EqY0v9VO3FZKsp/pJaybRi3VykIM5VJzEk
Ad5cS7t86PTiXJBWhgloalQHGmAunhpeH+/7Jk/dcA/BnTDrU38qfsYIPyKuYOHCuk13IKbAxQbT
fP9EVdj14iANpO+BnhhGuvAVsIUf1bYwb9wUcvxIWkSHlZncbVUuj5u+OcUZMAWzmw6lM9R7Rq0y
a5pQOpEIN/Fgllm3E6p+zxN1wi3vG51WAeVO4VZngTLa9zijPOoTDp+VP/Nn5CtWnuUuYVHPeo8G
vYz0DQ+Db/qNUMdjew1CqfW1MVzlnhmOG+598yUGxj/7caJvT4hyHu6NRCfxjWMT/Eg2IrUrECKd
eDLh3yTwKdzZacfo6yQAA1rDTeWP5gPOni3sVWvdEKdCw189E6KLJo1tQkFbNdDr+Dy8ynBO2+AO
ypYWPdvCzFTK/fmouq0cCtgJtk8XxWqu9/YZ9clHFKpn1YZrs5UCc8fIz7rSNBOH/jHKR/P+XXgv
TZ5VoradfD0W6NpmYlOCkS530/85xawT2LFf0xAP+Q4WA7jCH9ZxjbcshX2/EiDvqXTDCZOmjaUI
97/DHGAKOKE1MbyD1AwTiJqGp0H90qFNDoZJIXHSeKjtFmZIgd0m6Qa2Tim5qOZnXeNunf0KuhUa
7cGVCcmsJrVClYcnXkQgP8rjC7hjwm6eRGbArAqqS22hCAZOWruFrGXUvLgoNouZ4tzWu5XtIg9e
jVOpdCaf3YjApQp3Hn4/fJxhVQU6if0euG4ZQmuWSL5nEdZMw9oGJacp/n5rfSNtovygGi+yFFUT
lC2ebku0q/TxxQHt5Lk2vYm46UcDGWktkh+MoZQNPgJllrkx0gBV7Kfm2GwguyAcfWDkpD+Ot1w2
VPjAnzkOb4jbnUjBN1Lf3eIYoiIhKdjmEhCKWbHDxAKTGJi9/uU2VX7RXSn9CjowVWCJrKBJ1dh8
/m0pZaqlnx096ysCv4QfBml9TUKY7t/kjROzh+dNELo4f5db2uw8qsD26I/PROzLcrWR4cSud9PM
ExbHlO3LA33C7p+TI2QIi2Q+uPIwOw5T/Au79CtWIn5SV2NmcWyMExAN/Cju+Z1T4i38KX3E+yAk
Z7v5fFtporK4BlgOGfjX3SxmnZO7DaGeu5fjtLb+QYw4qEJnwOaDiGgpByXZL4Pk1/vAifzL/S6M
coJby4CBKGzD1oOzv2kmd86+lQMfcB/7mQHT299FOI09dYW7GghNcvhvKxz0pgyKJmZWa4I3rDMN
b0TUV4E16ZOtt01/OFpqauKML+8vSYbmnxsAuLYGlrOzzjwaIfhM8zXV1oOxRkxORAK5zgTze8su
vbCmF/NG8D0P2TjIUnSUhar4lOC3+OuDnQl1knqi9xOIQY5WezmKdZkiCS1M25VQsBgz3aELwrE6
r1sJejJzaawwLga3UK6veHiLbsMh0PeHjISu95KFG80qeqIrOpm5tmtJSCTyBZGi4WvkylXfib25
KskXtsxIO+TZQt42jx9YZ0Vh2WOpY4sTj4laBTHjWixmVvrpOBQTxt794lidZGTmVEBmFrz/EHJy
royeBOo3lYpvh2WEkNnOC9vFz1f1CO6x3iURL7yH19u9VUOwEh/mnVehBEqlZq/nrwgA3RcGaeOA
hSWP8P7jQ94Hf2RU8TPPJyVyNQnGFkSI81sVxCInwjU2KS8nZA1rmFG5XP4LWRcjTTZ50UOZsnxK
tieBWaB55KVzNNBksLA8mZcy6VUwxLYI51kDMUqJBrvIUGOF4gx7sjxlfGITCWAWR4spRitkvi0J
HKVZAY1GdrnLXsoZjn65mQ5c5fyNrq8oZT27ca1BhucUJQdMnSdSj6RXueIJYF5VNKek5Dy3b7wT
yrQvvydlbHRvgT1fhzQUlZCPassL3tzuuEC1y514jqpdtROYTJxkuucE1cmDksbFMj8W2GlNHqlg
h3KoR7xFcC4xGNXTrGUC8MoI1+cLNo7S5y8A8i8chy42G6i6uuE1CjHLDyYL/o2jFFwViiuambJ2
qZTrrnnqbTkC3vpEIl/rDg5T0CgiJhuMYSpzU0QroEo8R9lXrTmAsfqgi7yYsQUz6XQmpRg6jgNI
sxm5AHPdofWv47FDEZz2aG6flaijH3ej3EBdmY4ovyo5h7XfkAGHotis7K/sUMJG8ReN1esKiGUa
7u2ZTLU4Hb1zMGgGRsVbFIAA1hHk42Tnjh3dgyviCLuOffYxvU1CnzEOZ8ihVI/ylKSnAn+HvnoJ
kjhBAV/HRdOnfh6zVo6cG/tyV7KMXiQTCAgKRXEgDFi6GyvBXMPDZjnoA6D8MqclRQWd54Q6q02q
4Wcfe4T4aYZfH2WaKW1/RfoAymLiJQhDEd71qj+TZeBqie9Bu+TtBywHLdGX8dtVIKEG6k055tx1
AnbCC2SsjdeoWHythH4dvRGg7kd/Wghi1QTZAm0cKZHHta2wAtt5zcdcDakbpkyApENprip/qJo8
gYHT05oFeqVvDrDKUfAe2koM8QO+bBA+fmLELXz1AoS57x/UBUNTT7Y8dkvN1AlrEbGx2MwiIUZn
mlR6esU38vedJZWbmLdX89lLbDRWfdieUiEQ2UPgJvjdYjSzXJvRXbpqig6/QZmSTYBgoDyfzV48
GafWqGYgH7Oqpcbl3f5vZR4ZlNl1d1fz1q49HMdCIiSm0kbrgBa/YimBwGyn72RaCNh7q/ZcF3aw
JjK4KIg4OY9fc+0HSnCgm6D/9mAHw0ZsX6tVRmdUdpWZnc/YzL6vV0bAny7elRra2dRCmc42/eZV
+MfrDRfSvg26I82Y/Wb5fHzaicw2ZKry+hvIS14RDqDHkLlRBrfJgqr46mONvuJ3riKzv2Ami3bd
X9Dl9/8d6JkNLsg44SB6ihdIr+RDaMfDcnuiLeHMO0NKC6x2jRKLHhNFof2Z/EaZQwZMJxJkdkSC
jnKu1IkF9Vklhef5LDzOb0yayQ8tOIeDx0sfJRMso+iuLrvROGWq5E6ZCUMPiIo+jctCAHa79ckU
/SfYxJWbmNG6Hlhe+on5Qjw9i+V45sO35UpFgJkU7X/iYunrK+Ys530zcnUffEyGrw2V7Z15wV3Q
+T47VJY9V1nnE9IOZNcNL57FOFzOSDCx7E1XRxsQnpegJE9X2TC7DpeJNzPL2OWYXoFK0MRc8h2T
xd3TZVw6uR6AgUMpQNVdVrxl2MjVM7llF8m2exv0XolEoVDfOansP/RZ7RuXMmvnJ52N2v1Sx/Kh
ANWWTXC/u+foRzpzrVIWmovm63vFmFxo7A2dSNt2A3nwHjwyZWxzaptNsJLtpMQc5X5zmW5Qc4UK
MvmVenHtebMRaEfmtJCupmYQ95MDhYgp6O4988VMn8ssfPhQHiunXqppTVCkGVHiyOxdMgMZwRHM
GVQC2FiVVmQqkXAK0Qf5UbJQQRhlI+EuGrEwyGiPXzq9cwKk2bWFLPLO+GVlTRS7VOO72F4ZP6kV
PI7EPLCJIRTlxzfjdqHvrqQ2qvsijAxIHdtuZpPA85L+D/a1bxOAuQOT2FYmlKBWGG1kHAR3XOQ3
28XbPG3VxOikyRaoh4u1KgAjArFMAnacauk6YdY1wRRpjwoNcLyWLFPozmxPM5d6pWajaPJ4UoFo
CK4XCDBNT9ZvVOnImfyVGt1w589WU0dPKi/hSw6/NkpCE/g178zWztYI/4vAxwx71ClB2ITBqEee
IKeDqIjI/8798/C7ajzvfZURnY9B1d10eofy27ew0FVF5yonCR99kciMP8sSRFU6W8uXv0h6e78i
P0GoqpKteCrtnQ2f8Zg5keDuJ5mp/d3yeTpcL9nauESWjGSt1t7hqTawq5Z2L9uzwONlAb0C+vN/
jdW6shSThHIKB+J85XS2m5504cuTdRBNZ0zqwdr3L0gTQ4dzBFfFmamDZpe4Ss2Q0fZUFuLMK/2W
UJ1VB1ZfpnWw676zdsJXanvWJ2kowoBV10H3aK1s5aDShfxMPpKbyzvh2rXv24nFUENIMrMX4I4B
1vyLDg9RqBm712fRmKPMXeZmRqt+HFYsph+nu7oI12Hy5yll7RSJSemvCs5Ymf8zNI2G6Fv02Jcq
AWZev5WKQxg4rR1y95BOXA4zG/5CobRUSQQ5U+9tlLWfoZFbzAX0N0PG0F4BepP8Qwe8ld16/5QC
UzXqcmg71HtdyyEj++/C7nbvwSfcl1G5vmhQgRjy1im1I8iMjL6bbn2pnszJhprZFODXMj2sne8d
9ml6Yph+0eo8he7qVti3Es4e3c1UxeCK+0PmBSSSSFXNF0LE0f2jaWRbtbpFd8ebWIKnd+6HkIwk
UK08XSISFOX2W0hXNwzAvH/NbuxzicqzdS2xOIPWrUPNZrlFJLEdqEG4P7nLsWx5qetWK2KlXJSF
lBfh4M8l7nJzVgI273X5a842BuLAnr/AcEZkBVvASYJiogzWe+gpLMeGRY4wueqH6av/yBxrPsjz
wflGVoq89VXzH/4nZn19sqWyVT22z/0kDF9sGJpCaLibPJdGBRCCZVm8P4TitprH2CKpJE4cUK3j
W+SErVBDw4RlaBOR4QgCZpgn9sj5LAIKAP5YiOwKfHDrBv4Pi/JHCzLJKiL9jIbKFG/FeK3n74BU
a/x/sYh31VDTJSxO2HcUr/EvVnKKVILgrXnEKkoARI0rnt3Fcs3rXrl/vVFQJx6TmmnoqRABfGIl
A/nY5pVNEHV3Sm83Fitr/M7ucFvmHMs0nZzP2VEswRN5+6c867Qr7dPakgrjGwHfEQCaWnnwnThu
SJ6MWTwaPT/gwQEMzyBVEjJhp3PnuJOE0GovzEmpSDqRAJOtR9n2TcykYe9DvmJpLL7DgY8rSYGf
vzkSh0Vj6HtElwpUsqmYkRPsQv/A96YE/LLH4ymlAaPIrRDOZXAIJc4Ds6RKSli0os5a5Epb4mOT
/kbbbTyOXgufXTD+qmAgwrk+YPUnp0XU2SndTRS9K2fbqrDhZ1AoABJ8BZXivg8gT4cYbYDdYf9E
FAPa/G6FhZiCAV172xMrv/lh/Jb6g6IJeZmOcs5QsA8vuZjKpntZbYAWR0CMcgMh5mCJs0yWdvJ/
vxeNcr7xbGZ7YFyWSVnU4G9k+isGRbz19I11UUN30L4o/+3/LNYNlrGmIY+wUhSDy5oH2u0XT1R4
hAD/NxkEE1GhMnjo6wN6JTVeXVjOFaaRTNv1wWqJUhpZ1mnWsshAS6qWy0e3ep7MbYt5UNA0p6cS
2HcJD+fFIMBheFokFfH7NvOrv6FMzvcyfYxaDDU4HIFr2Q8o9/LpfTg8NSx3107lwkKls6DIxk9B
1T6NArNuRXKKeQrmQmcQUzkcPtUIhl+u5731tmqGTo/+WokT+tjd/7GWf8Q4GOOOkVVWpMvS6Vd7
BPfKw5NkiYkx9kdKCjGABnosbN/PwO1LRmraFJkpDV9/D9vtXQh+5vJCQlowKfmkfLukywT8z3gk
wxFXHnmciTVlB78j/0QPO6BcAEo7DHXRzrPP3Hx4Mn4tw4V9Wkyc94hezf7Q7L+CkvYlLCnDfKcN
YEae97E3D5pRtkpJJ5671xgY9wC1TWlkRvHuxbq1ura5xOoVA+KfzxYjW2xvWmgRUm7/zpyJCZwh
vN+CrgZGk6Og2obj0S5IoFVemg/PGlAUDkrq4F9rXZW5LSl77KKdeoWkBT2oYVP3ds4syeErOBdx
FlQvVRpGjnUFgqTkxUColwVYi23v3dabWVJUf22ShwKXqIvHCxCTdnGAuMe6+OSN3ICkZYw5Y9T8
r8NPrmHJ7vytoXAR2qdpjeFHtzSugmjxXrSnrEux+9y8HFI49DVVQ3ri3G8EMBWssRjc04UjLc4b
6YzfTHlzI6f1mogL8IP0mU/JlD1Opq06chAHq6IucGDQO9s+AABHnoGDxtkfwFDr/urclGFk0SRN
nHpinNrm93t42GSiriR4R/9HR4f2dfVlritFpztwbN8L4Y66EsL9GFeX7D8hzC/Zwmie0aURj/+/
vJNHDDxzMZPRO1xwJzcstgAHvMuHd3gTamKxu/inRuvu56lyidUeBq7rQIFlw8iIWmgEbbr2JlKX
o0t8ZYl8xtV98K4dUrTSGxUWUHEv2O+UUN+ypWm3dqamO96XXhUEKNHE0ZYF0N4LKeQcSNlvzbcA
2ksmJ/bOrqbnZSLHtqDglhrE/P5KuDbrmI+MdNeLZ93I6A2fm5GlW0vKx+iz9pLz4sSqdsog6wlR
0YyZ/qv9X6s3MRYTuJQBQodplFYfgkOuz0MeARxcVEc+kp1akTo17x/qPIUShuw2nXZfZCIVEq/D
VLRnDR+Jmv9pUVM4Bzk3CPoHadnVUuDhfzwNzTxi7RSyBvCTXOJorvgqmClyQKxKyeSC9NzEK/wz
8OJt90qtVNjJSTeZLNt96Lmq60o17t9CEohBJChpRJijs+JZnGURBP9J0RbhMisg/FtOsgpbun+/
ppNM0o8aID9+VDkHwoZs6F82L7v9CavzPSiHwb2wTdDKjO1orzYXrSUjcHFuhoTGbsjsT9PAKCNX
OQO/7kP+2MdaEHUsfwJ2kkhQcK0UCf+wUyHwfXcqch/beiQrXzix4azBLxbcI9Nn6iZnM7ABSxnX
jHtJKEsZ9tZKsCL4ftSkAtMq1zhqZ/6zsvYqe58SqTkyPG1O9eHr3pxN3Qi9tRoHQXaO5SkKoZWV
BT5x8RwOy64O+50LWJYCGFNluIZUmMX00V3Z+BfYkXNb1aKuZK5HGdZFJTX4fiEe6dMH5yIciKQh
vn4UDMRs1h3fW3kXuUgFNT1h5tET4p37OPfuyJ3dFyL+XNt4FsFuzrhYUJgRzrvVfFrjEYINqZYs
ZoE4N0pKIkyQg3xj1IoQHlw47zsvdPhRxtrMiBqkm22wfDnPueDVumtgd5d3mPXGjDhCEuGtuVOS
IfR4/yKld4zXxf0FKhk07RAHafz34VdHqdy6VFZcDQj6g/JT9q2Cf55lEyIWY3hBV1KaU+b5REZH
JCYo5rqclIKfQUG8Z7CAmqP0/2WUy7bvWDFnrgudufUAWf16c/P3PitE/myWCZE7EAon9pRx6uOY
4V430/CgPxiXyMHR8fWB3fWVhaQk7lnHXclvFqG2WfS7XRTOttdtaMF5bqEyCxPcf/gJYCz0FMpX
/MnZjlWN17ulIpxUvEplW1RF8ScIs0pbOqL1+SCuVYZc+YYvZRry3rkH/mPJN5fzs9UyAcqpFTVe
15B3bN5jTp40iwgeE56xSZJScY+DKI4qRAK/LZl+Af+1QakjwGy/on4aNXVEOJPJ1i2wGGCCgV6t
MIJebE2rkcZfgrDXB8Vw53WKnAXkZVI/1ASFG2AtQAKTlEPPcsZypTFJS+EbcewX6MNgcvf4OINQ
oXfSVFQCNYdP2gK6AiAAWjGtm/T2lyCuktQwCqZJErsM+bFsiPWIHVuA49bliOiDzzsdppjQwOlG
YR8aXhQ8kcMtaj86E566xxyFFBVYf0TdrKZPOGatnvUMszdCmxcYdPUL9PsN5wnJ/Lhxo/xUjtEF
ZJmOERoJJLChC6WihCRwI2f4bx+soDul7K0se7CXDblUlH5Z9A0z6E2bh8BPRUJINVifvbvbxmSD
WAInmXeg/EDzQFSl0hYqNWaAEcr1F9pa+hAs455fO/7cL/4aGaxYf/G9rDaOj8nxJr2JFkeIjv0W
YEslAYH7Mj3MKtwKI/mf2f1BUmqnrbIsTDwJJ1U59VJYVtqo0v7lzNBdS5XUH4RVFR/mWLLI4cx/
U1zLpYyZBTzy4F0ladXVVhCIbbL0a5r/XXyD3DyOP5PX8pdHFXQW8jHNOLfdOpDpZMHP9DzOoJzV
OqFK9+wNDwy9iLhN4oS3gYPJr4AIz/2C+9+jHU+UEVnAPjIEmB7TvcjgxY9FlYNCsWNG1vOPvbJp
9cgqx62biEg5I+BtEOxQeAojrEGqBwI/4BSt+8VT1zraVZhVXyEI08xqiD6OkHmESozJ/RjM3hdZ
P7DFIXJs0EE8v9vjXioQE51nP3JrZNpmfvlAhYCE3VylCII92f9oXTOCI+3bUS6pwb2wtYEgBXgC
OMzY0APBSZHPQkeOOVAJnum23HBoEhayaqy39ZM4ofJGd1yDt2vDDTN3AOn6Qhf6TmhzfmEX2LG3
6EGNamD0qIjsb9L8D7YhLYDSPjjWzchKkTJiKXN1DfdFl6j8OhlqHFfkL+xDnkuGDk1ck/vB8UAy
cdIqqZT8AICLbNxOIvgIWBq3ttGjKIefKq3+0qMaT7dI+KxfoyogicR6tGq7aPZf44jKGESG3QX2
2AK1KUygB+NJ7H7UEtG3V6VCTQJXnuJxMMj6G3HiqDk2uubwXf9lJvkfDkEQPxvXBpuL9csKTFB7
XsAShbRG9PoEsCDOrr3Y6uhoHW3edxLA457UlivP4bdbtgQqtVquPVWdLaSE460rdoQ+RN0sLP1s
R22CzPs5NKBHRaIJgMYqaK3V7w6wyMOjd6lKnyAIEn+lPKuG1WqbiL7WpmbcT+QOLXMA7WT+JgEu
ppRq8DCPyFRY1yF18gDaFFOJQd5t5UhQ6CTAfXK6ZCeZHyTXJjQgvWZhAemLyxAjJWl4oZyiCfMN
cbFQEdkusEALQwCRG/AgubthEPAK7+HA0gdK264J8AiPWns9SSAMWr8feWz14dqVWRGcVHHpZmjs
IPrbKKc4C5PnKv9/OBBW8nL/Wver0XsBhbfF2MI1HFrnjfNa3sBSL7UTOHwLxe+KVQiAwlW/My6J
y8ThcazStNdte0DfK7xvSW04oc/SPV37W1D6he8cqJbtqzo2YlU1SFgcID0yDrPLZVeKdNFY2h8L
kW4HLLjWQIiIFLm/JyZyZbbwxi3dd7TmawC3FMoAUJoz4/kYhBaIdpdGu/yGqQyxI8A6PXydTzOs
MWpeN/IKM0MCC1/Lpir8Vk+zF16GvC1OfViIu6td4kFiFlas1joFt+NoZJBqDod8S/vTFOR5JzNK
HiAqqr0kRBf1HzcA/TPU93h5Bdk/n5Fw4ZMen2ZeNYsOMYHO5lGkH5u/cYHNUgb3RDP4kLVjLZvw
w/AWwnaZ3zSjKxdB4/jyAUo+d/hApuBghDa1fFFJ+qbKcAaYqxadLFpXaQ6Bb90H3lYSXbpYNFep
10+88nESt3saR2318OgVqExyzgViLUcfPC6zUzWv/fHiVI+wgmDHG4RDOGt+VTdhdstQqYAqMZGt
X9YME+iz4/0F3vxhyJkN6t7DDLJnWbHlfQNAONCbq/mFIMZ4OJ0k0OYqZmo+waUTqCSvJpDy79x5
MgqG/vBRIdtZAgYEcexg7VWSzfWY8Dyn1MmpY9D2ibI3YjyYFBL3LNSOyaAl+lUHLujKe2MHE4rd
oAMQPCxofQkyPg7rlzvcO+QuuJzjCtx18EvNVAPvf41hEoKnoiBCbX+hnYVgagcvA0lCnl7xukG7
iQ2slUakP301TIjafxJJNAR7mVhVu6+seCN6/5cr6TyNbx14aqpC163Dzib0hQz4jx4SWG7iVpw8
T2gxJGsyoW8WGZC/FoIfM1D+nbR40Gbslq3gMJBrbJuL18PF7sVp50J/GPACpHpo1XtQR39fIlW+
naGt0rieZngfvnz6ljtXHa8SQmFEiOtbCRspdCDFevmMSDInEZe3gMJzoYvsKaEnvogtiMgYD2kL
spupM13y2ZUZxolfQUF9af5En6NDopIsou4UKHb98DRB7kOizyx78Rr5jveUkGDBaVMpSRrD3QtZ
HrKLrz3Zycm7sLxlz5oxzPblrkzXB1E22ABKz9GvnTCABCJ9sYesuTTbqrRI9vJZN05Y+FYKT7iB
h2zzpFWtx/tdOAZltGc4JaeaZQmhDNMo0XigQGA9zUKI10x+hgSziKHK5Bdxa1SvFor6S5opE6SB
M+vb7V98iHE+dyKCQofkPW8cX/pAtBSmuQUDZt174FJWXOCuiP6Epp9wHKe2GgjATNbNVRwzz7Sb
N14GLQYNa22gr3O4NEp9NKWOZnU7wdvaaJNwJVUouy/2AWlK7IEdVdw+aUWHFxM6fdRZFUF9Tp12
cR481aC1tOH3GkSf88re90VoOFKiIzV0ie39uiphKZV5fUPCO/qc4sxkDN6MGT5yM6ZQI6pKqS+Q
8apiu26AojhD79fSF4FZyCkVzc6FASYH/NJX+9/YYhLcJuZyV4mhBHN7vB35RhRPqegq63XHVZDW
8axt5Rk+g0U9yNKgMmiCLNd8VrjhxkIlzTY2iQIVlP+v748EyNz7lEd8diTUCZ3WjZJncbNtIU2J
4O/RmKGbIGPvl5/wD5lBaYFZNezuYMEHqV6fYWvlF4U1xIjLmDZuNOGI4rOY9CzcHfxsMwG8wFAL
w3IEEhS7mVXak9ty8CMnW1KtliH/8mGpEdhxZL2uA+4JYm24Kwdnxs4jjBr5wVHKm5oYBiMGWlmQ
89HgOX3+hJ/PXWWviyr65v+bsPq1b9ihAhs128JDqjGF6xtDEtQMEmfNcDzoQ0P+CSTVdgP88VKz
vGq6q41W/B8ahbaSqRutqirkyS16t5/uJPT+F8dF0rAix4DF3WA5TLI1FwfvyWfcuuW32g82m4k8
klknK4BCXvg+PkOpDR9aRzYUspaaVH3V4z+3h98wN5vBpCc8E4hp1w//mKOKVOw/p+E+GIWsu97F
L0lOdOXI03cR60b0ipNeIN96tEPJfUldmHSoe5Gk8SHsOHyD7bsaRM01ynC+6IxeWQksQzf6K0/E
3Fp6c9aw2Rh4WlAj61OV7yMLusLQoclS+lsXSutJkA6HH0kwDzyl/HImkghS7zgxltACylID4kEA
uEgcLh2RfzRMH3rXt7UOLMnVGb3WCnejZbQV9w3BE2WEXhafPjROXdjGllChWBiR58AyPfcYrjcC
z+z4XmOjMeu7fOIWe+ttLpEZT6PllgFxWKGDKvfDJ6VwuJ9jYziHesnOiKQgxz/OOfDTjl3xz+Am
elE0/JqtcuJ88TRRKpiYzxB0hfLrsWGAQUaQY/FosvKcwlqLEwzoOi4GFI0zlgv+JswOBkDjEKEP
yBgEFs5vC3wSwtC/2HwkYdpCRNi94FghCw6asgm6fzC5nuM/94W36PTkBvY3C+XHYxLntDX0FyAK
92ADrijOkp/Tx+lqBOyh45oJcMyHtZSs/6W+DpC2XBu0deESowtD+UTURB1c9Gznn+GRaibKYJbp
vl6un25ET0BWfWwS5TXQart+uQTBgpM8y5WlpUeO6qMw2Y2Gfzz7KAGVUkE6vW4RnLf9VXev+i4+
eRLDm+u2TQXV4NM7ynDEsywEuKa/gC3hXV0x8BbVh7QmkYX9h8sGMDQq4n9Fct3Hn2TIw7ucTaYM
LTYRTEUi9OeEUvynoqoW4eAusVEk3uXyFKdvKvGJ1vigX+/8A0r0dQIc82Yy90GrPkUF/HgMJVgx
NbMg8SyR8MkppIJaIJCqF0xlQW2OI48LX2uMhcC1V/Kj4tXeyZbLkgA1IUKQK4aOsSsc3ciSCIQ8
0B6P9+iXOMNKH+LmDYER4UUJUI1wcnby4M6kRWfbTHhVfe02hiAO5s3oeFN04aobPM+XrwgrTZg9
RjUo4WYkdbdlaGNZ6GwhWAAnL0X3RFmU1ceNdseCbUUTZXMRzMCF4USCaJb57cV67QZ4SyLFKDrd
5VxCOQi2qVkQ+EUK/Mv42GIsuO6heoFlnaUuEmlMJNC5ro0MNd9Vg3oXBPFU8IS8lGMImhhpOL+B
S3m7uFC46riPLJv37GkDxfCBNehYtKsZMCn3xclXoYfDydYilqFeYZbL6V7eEnIk5ckxPByxg9wo
IJvu76E/55V83YuNF357jxEPPwm/f1CGKr6YUBqiEWQqyksFuYfxErfcRYbTJbrTFMw/g0pUv/3b
Wd2PvzlomcGstzsfRAiB+62QLJ9Pu5RioaFJELh4iQIN+HyNIQDGMFS5uoR7Src7iEeA+4ypI+Sx
gDJDXXYnxVuWUYWjwGCs92WAHm2g7c+RMsFO0eMG675PqS4sI1pxJXt3zEdsm8bbQWbDMS7QLCFJ
DwsGUCtYSz1qCk+2W9FlWLQeu7PYdrTIALLVXriHXvkddXP0GDzLy4zOSqh/WT3FzZq6bXJi7/Vi
z8l9SoaB6s/u0LTeJlzRSze7dUYTUjLnlPgV34IOkzxXIIy7v6JnoRCedUvv6imP+k3wp/+zMu7A
3lJMky4R2MRXdYvCcFSMMpeVp7/h0zNbCztflUEv1E6bkmNHLWDR9UxqZfOMAQfDpk8W3OiNMLyI
iJPr4GeXme0TBPI4ZxW7k57kT06EOLgexQN4MGH21+fALlKwOb4Eo510nD5UT8QHM71lvBd0tE8i
eLAU1APN1Ow0UIatinwCqFJ5uzQ/dVqOA8WS5DWRih3fPBhu5yBCR+lnNWNp0Koxy2Zt4O30gb2q
VDLeRjbZbkAd4LUNbgHOpUAph+E+MJY1B0VJvjlJWYrXl54KU7CHtTGHDplwJcz148scHZI7QSe0
sbUbmijW0YSXEqV/QnbzcVSrxq+APWq0Opo1wCuOfPEb3kfhF1Ma3coIPmVT+i5hf3aVCvy6kcGV
MOPA6wHsXmjxlh1Ms/+vR8D4mPutRykGGKgeC8CgbAjIu4tmR70kipdl2hOmuGOa59LwKuZjI/94
sbv8Cl7UPjonzNzWCwHuH3tCVi2EseRqvgZXF6L5EUcvqZJNuh+AUZA6RThUmVUpLw+ofts1uPpl
w+gsYuu7BZL+IFVj9QkqXBzt+evLMWQrQT0VH21q9MaEwLT/K8EaRTGX4/qCLBuQLUEfKagJ1+8z
0Ocpv4NkdrfJGw0gSk7Ul8jGG37hnolO9yzGzv72EFlHRDVvtuBe2B481s8MzujWNrDfgX752uDD
+gog/T4ZM0htuBNz2UAChqJ16Q/c7hbUnG7tOV5DfFMJZvwdBV3jpu/t9eUt0/hdpdfesdGMxgGZ
Dl4vqZBl0ru9OYPVnPJXHJt7Jvy5F44XuKEtr0iqLelmhD90ky5pBUXswd265Nj0b29oNUYQvnxC
RA9dvv1qxdziUP7TDjVcVyccGiLX50dHcSN5BPOFU9EQ48BoHMSzDPPToDcXROXp2D5aA9zHF+b8
/NjjUgy3/Gh9yfQrxH/ovO0LuyG2wHJQpvRFs6jI79WaCyqPMt5X3W1gGKTyB61WGqXJpCJ76HMm
AZy+gqM9x1omNBxdUB9zsWEYiJPoX4sWuwCqGOlJvrBmKLkOUXZU/RZ8r+d0asO8yltfofMChwDf
j15cqjd50v8hO9F8XEAomEsjhkg0DBLTSOXeJMawNcrHw7hMBvadoEZvxhnz2wlWw91xjFxftDFu
KQ+xCb6NmwRfZhERj4zFxDgUc5lNRaoDiVb/aUav/SBvKDgwYR0nNF0VezSvAN5441kVxs/tPOm3
GAA5qnh+vLou8KRs788Y021y31REdCUmfIe7BNE8G5T1A38BhxPB4qTi6KG6AJWy/EcqWKQotpEi
VxWdBcOthZqJACd6Ga6St9pA9XXXxmd5fnrv1ndXSMZi/asTyyOr6WkWLuKdj++3iIltEBkrrp1+
rypzulH4xYIVEWskwP0MZBQGYTc6m6alZU0SujXtQnEX7HRG6hKfwI3psop0vfOVJpFwtZFyhH4P
nT8xdU4uQT8/8r1b+bIIf0s6H3YHyUyszbTUMzkFHlmfEd0FP9ZRIAxIglYO9XGgSUy6GA5wleW5
hdlWhTmnxq6IPJcso5uKUJCILlOqRMuIGk8G3aWJopsr7LcojFHf8/qyd8YllXuYnfEPNCM/02pp
d4GnoBlV8ixwRv2muwJv83xOIaT5TIZt87aYs7ISWXoagSV0eRXYlPZg55WRd1FOaDS5jYfpzDvO
mlqwKGOR49AbUKoL1ddwhefYh5pFP2lA8U07jJGBpaKmQ9idnOmLFe7L26Y6pYKQtmnEteIQhYkO
UKwq1jVkfMpO1GTUZphJqgfWSG8uSfnFRB5XHUcGjGADQ4t8NdzdMaZcp+3Jy75pgPMEnNeZQCWs
RFKV9ZAFI5mec0RS8NNOnSHyzwrLfLTkVOGVovMA0ZNL5rnaeg1BeO3ri+2HFFshdGQxoTtt7V4j
cnAsMwbX3TDQNJ4uBpEmjIidxc0D5qVOuQnQk+gilW9nzS0LgNRepTOIStB91u5Yx5t/Uf6KsabC
9Gbspuf1enXc9dqMNh6Bbmre7+0X4uF14ep3ky/i0wF+9A7vCxkJ/HsnUbBX65NiNz/rBaSAYwE+
nuddvZRbNdoyDGTSW8WEHhi9SNSPm1YvozwKqmIO1w1FnfjDEfpG0VBecLcXdJV0PLCHiEXUQiFz
ZJApqHJrlRE4SnWBrrJ4UuOHkwgigey9R9E3mHku14iSwFJPdO7SJfJ/BrNXIqMY0DsU+B0TMTIq
DV6BiHx15vFi+LM6v+UflxUykuedaM3pCrmDkQJsaUnGmSikHF5+9rZc/DEfDp3xe5fcAUBN4lnW
GoE/4YvDK0kNaj7xnfmM1khdG300IuqLEUyflhb2YXat714aBOZ1YWVvvyEjXBNVYp4h2/6P2c+G
DC4uCuI6GkRu0j64NfvHJIjpQkEc89OU93JBk6WDx/aEtqYgEAmrjiKA8CUNkYE93JsA/48KAuTZ
eGLLw9H8AbmCrUFQTse9Iyk7f3f4ltggFNJ8nEKoJY/8tNIE/5ajuzbqN9GpETzz2JUo1r7LXQs1
0X2JRBOy9UY0zqOgseI1opRTMBU2LZYpkCgrGLyPrmR2PTpvgFh9vNWkQKgMf/5HNh0skeeS5sZ2
b/+cmoTql/WE1+R4+re5qIXFuBA8rZPluCNLajdIHYDum/opqlwrZ6NJ0pq402OA+6IOoq6UIYWH
dk43BGGHHW0CYHQ87QjypuBXm9WeH3Zq2fBCwWqnJVVlT+Sxyl74VR0h+LDUaWykTsQKODwLVgvm
tyqXav3RDiCF8+67pCH55VSvo21cmPQGSC1gYrAzGwqN3AQdRyhYwPj602HwLHkCdPwiaA6FbeNR
0Y3m1uVruIRMjKgAK2KTppycOFeO016tk8EV1roAnnbHjSqlFvqDNhlgeLGKZtNzy/moG+caozLH
+TLesYokAt9jn6+ZqnVmJwDWsoQoZo7siRitmbOllF96qt8DCwlYtIyhle+FQEdf8ToORCyicUWt
LlpV9hNHFsgyRv+Pi5iod0p/8uD0jFqnlN9llqUQSsUE1inAXstVSRbUKrCnpu8h04TBJXF7X6+v
5xWmOB8XyO0yU2C/+7dqz7VdIVdLoCdsP40TL92uYxvvJTXV6Xw84BYe1104q12c76XfoJL7czFP
54mIXS55uVUfhlYO9u+dB1C88Eihg/hOC3ZbaH6Dsy3cV9nrdOZsmPNh681Gp7l2EJhx5+Nb1ZCj
S+0MRx22xtJLhWxarcvRRqlyy0AG/B1Hk8m+673bQNGlb8D3avGmEYxnZ+32pKyYHGAubGJYhzoU
PIIUA5j7w3ijHmfGkbyZg1FBimhC0YT+JNRFO+rmBnkDFU1F12rrhHftX+YYb2b2lgUuW1vrhVao
y62eWAg3SwVR3/jwgICo7oUnawU6uShEQk4NEXkJKfGDwv1LAijAA2BJhTKHfsd3RrYc7u4xuSia
F0LcMJdea7LcuRVtIc1cU3blkyq6J9fx7d0BO9wRna5QpNg1Ttui+C2Gd8duYSIuTC49XafemVJ1
+Zi6GF2kzcsuRAPcxR215wsZ51drLHl56rraBHLHGqYAvcfa9ikmrOb8WNveaqS0h/xvqppgm7xI
wo3/U24O9pVm+b2ghKJmGdujiWi9OPYCFzYKmbXpfy1eFfAjORqqi4SyPQgft98LhBTmZ38tvuwd
igi3Q4jfhBjM4QZg3+sBxHqz9i0n5SfWgf3ifLRh+n2hx6Fk6LqTlGjt97+pV173J6b9SCFxi6tk
NfrVXOnZI36GZk4onmDdN2DZvuIoaQ7JyVEoyJyoQyB5WnYwn2qdC1Cuz5K1cgjxkyTVU36a+UES
9zUSOmQNG7m94KfjlZREMwJH2B178jjXUhpApSr9lB82mim/bmyqwet69InnsTyfnFDay0Oc8RnR
oXbb10WWtWWokJJxyniEN2ZBgsh5szztz0I1vJcde/mSxTToW6cMNBLos2n9ao7tqQ7Rn2/AOh3e
6JTu7OSylIyC8yakF3rbeUjIppoTPeybVipS6LQaHnX0cc8f6YkKYYIeyyREsGwVt0Rlxp+LvOnx
D9XXFiA9LmRf24tyelKT8MWIKG2RBskjTnJTeg2N4rWgKyXhDLkOdrQHvkBzD47a7uHPbMXc/aiy
AVIsoZPOS2OXjphp18m/uuP+FjqwyfA0L5UCo7YSWyhDY2gtm9wwHh1CDW5GRh3nYwZxFNh6ndpQ
rCVCvLsQqQerw4qPzztpvU1u1rduYd01v+LCwrf8J6Va2LxtNRNlDCSb+Q+oTqOcmxP4Jtgr2hBg
AkRbVE+0QT63u7B9OOevTdy+PjTRFlqLqvP0TTgYx9sOsRWMagEazSsvNjp31PhmTJ5bP8x3s5PG
LK4sOiYuzlvcr+yvpNWryMo66Y7SkpQk9GH8ttEAOlHK9xqu0rJsYgSrpWftSFqcpQ54QcaMNfw5
DPau44L31hRXCmV0faOQxyqVw0cDbON7nXy59znl2M3OC95C6jXRwJ1rI1m1Z++Ye30fD3z0ZNyN
hid29zhn+yszwH7fWT+AuYMr0KSMDxMATH5Ov2CHP/NQG0eN6LkHDHSdUjOYIpcJ0Ve5x0tT0+L+
gSxLEEwnie6whaPZhn45ENC52g+uwAUfdl78+G3dUZqxHA/vquiClVSfE0/cyk6nzrRPd57hQxMF
DFwls99TUkxbVtpb3cDG6zV+JupmdvTZ0Rh6Z8SPkiTEv5UHfhzKn2m7ZttRGu8ZWMaWcb6R93sI
BD/8i6m9clsdMYAP+x1RFkZ66GHZb+GFQZEFnPw1QQgZgMh1jrMryC6moMBijp6zqOh5z9gVuCfs
CzurmlmJkCi1zzgDj7j9PxN6gs+Zb4G6wo0PRTmk68weIwtxYjExkXjIQTnPzchlggKw/5pZyq7S
Tq9M8HH4VrgPl2sY5rUztlNS4ivjuQr+p8niB6YHlc3PGdyEX/K3EewV6e2rcd2lBYOl/wNBOv5z
68Xvg2DaMS7olxjHVVQARKqzKGXaeAvxGvbDJdwvGcW/yH7JaQ8RnL+QZCGqkqZgoQ5Ey1lNCG2r
gcXuvkLjAVnUhreTZx+WyTFpE4MP89qi2eeri3AOjBUvypgJS1nMVmXa6kg0nOggnKANeere8b8H
LmcNZAq/9CBwkAwMaLngrHzCOIbyv7wr7jUz+cHEBq0t0fuq546qf26i3Uz8xW2kgKU7ecv8SFQr
DxuZm35dNrWGzz1gqWVy5pKEYj1WWvvdWDzmQMB9aNGRM1UFZqcrHhHff3T9vibIeIw47EZAO3Ad
BepVfGe9JBHCuiZfMsVe1Ye1VE33d/xO2uAdjtBMOnR8wc8u9pfNawF3fpMdGvOkEWD22UZDqKOW
rGaU1qOZ0gex0p5VrpalLM1uMqsG24zJWLL3BaWHfFyGC/wTG1A+I9BR1gsAUpM+2oz8qZ8W4SwM
h+nzxBJMzD3CI5RdtB1YyqC1U63ljLYo/uvpoUo3KluKCVLHG7FK8MSE9lhGfgI539gVO6OX3y/S
9wxJmlAGB9qk1gMiJ+WHS1AQn81VF3yP1nPmIYIKHTBYh5/gXj64WHmQI+PD/iSPhr0vykfOCSyo
Tt8NrCFXei/Jcfp1ENUFBGcoUpMdBzGsaA+42JcX4PriA3az4WTWVaAeessCqs21d5Bi8lkBiDYt
wkD3w2ry1d+lRaYSYZ6UPqIKWq2EQBmuTpifUt6SzlDW7rGV9bzDPefkZ5op9ebCWMPExHXi8CPy
gJciSKk9SZsnNF7txFNe1zGZnS96Aa3TrQ5NdsgvJOti236xb5+6SCqJ/qPjwbr9llU89A0xpAwj
ET/KeykZXRHGipDsokv1P4iB9bhKcKpZPypLY9Qiqc26evnUeF3eYtxKCy2Ha7VWXV9KPBGDU7p1
w2xVwBhSkXsOv12SZq5MUJe1+lvNaVgWmZTa8NlMumeoXiwlI7GNLtxY8i6TPmcxZgPgbuEbwEG1
kth7a+wMBVJxvGAXZu7wVR6rszCQEdBWku68P4miHN8tyrWRpkuZweamDOgb6tEr14lxmyAlI2T9
Nk8wMD947aONZz2Tlawf78uBwowxVnA+N4pw9nS9XgRcQABVtSbu3cjb5jvY+FSZBTjIsmJTvBON
IJYlIs8v9T8FfKhAtRBzwvTQbVJEk+I5KzjD0HXt0+4SdUTuH6CnaNwRECrlqe998VKdA/frpVWT
vc+gJWmYsMqWVP7OK2Kjxv8V3QfMG1vGUVujemhLtI3fYeRLmo7cRfmq68Xcs6g8EKpEEt6lJ+uP
74d+631QmHBYZNvrKMRi88R8PuDbL97Iota+BRGuZQh8iHl/jf7B4PeDvXLQIp+EfXFb4CJszz4z
8XFtIWg7+iheOVp458tMYltNbFMxIAVjMxWocUsBnycdCV0WmkF4bOSVCV7+a5hVPggd7sUJMn8T
0IYlYeeihUVuKW821zOeTPv2kmRg2zWGZyAAWfiVfAcXGkvyVHnznj1uXWTvmJ/UVLNJw4ZbEJIa
aQ7yu0jXNsMxNKubBTKV6dxnw++T0/3rpmnPB7IcHo8NDM3bjmfUsw3zQxfFH7St7q7iR9eP3yRj
ueTayDkpSwZc9nz3StIRotP3cXRC65mi+Lk7fLvU54wizloDK4mJlD61nvu4tToIlc9kBeOXxrRd
90Ax/nFJla1HBQOacMtq1C8Tj5W7no/9Ge025ysjFXgoaOHpc5s7bRGTplMdbI+YoSE1pKDksRx9
iHhCpoX1qCd6LEm1jpxUA9aATpjz/6EtJbXAtyzaas6B9UCMP/5oCdAj9dAEh2kGVgIgWO9lAcRX
n2GpODFuKVGjV3mNnuuSRcGVYBtpTvnlHA4p5IhStzhUuUUewEvBv/pXhJnp0A01z1eDESxFC/aG
HtqZJo7bKsM2rs0sIva/A4dxccXA4XRVDmYsOY34iZgAhgqbDitm2voPIpF4fjEieeRlKa4L1yuX
onLn2HZAovIujP7PdGZfm6cM0l38AC51UXpym388bFScZJ6V5mbgirVToUj4bq8NrGxFXA5eBcQm
KAP4sElXbFPZoDvk2YKT1aJqt5F58qpam7Ky5aEDdAiQrbQv6agjW8XTHx3H4k9mY5sAF0sqaaxD
tUQr0HQ255s7yImh8g5eG8U53NG/2fdzT0hFFclet/kTL8pcHHmWNq+2Crp5hqnhnnWVwUbwBQ7D
aRqTnWejVN1A6y0M8M1OghR7uXp53+xb5jfi/KeebwFQ14YX/kmI8vC18ymKcXADamZ9wM//Isdk
Jvqy32KweS0DJ0EcSZvja1KVsgZaJZ12daciM9I4d5q6IePxYWgSeqkHhc21YrazjN9yCHjrqiOM
oBtf7P8K/pmpwpSMTKBn4py0gvP0J3SY4/F3d0wHXEnQpqkc+WY8kqdP0zbN3tjp17GuRp/YHqnF
pO8HphhBFnR61p3Odn6lGepMDOSwIRaQRakoywhhcydco3Mf+PUBJ3rBNP159Js9AGwwc4U6tY+Q
f3o5E+A34kndtTBVGu9yM51aaqStEF5HA08qoDNh8Hn7cjxohTqeHcsEN2f0OWxZ0oSASHOVVcdU
WVnaqjCheiHj0p7WtIRRSJoF2QEk2ZCFzhw7pKsL+c3e4/zWpp5UlMb34DJ/IW39zK0gjCm/wiNR
DK5zGYA4H9ontZRYxhVKfncn9bfu/pfSPMM5NM3QOqGDB9D4MEutNjeWQohAKmPclVX32Y/NRn4L
P80QuTYlQgGRSm/mo37N1umsi4igSbnE072fI+kCDordqEm5L0o2fIU2R7DLu+OIdNBDov6f+h/P
0o9Xw/kxpmV6Q1WNzOnJuu+pE4hd3PKY3b9zjhHVwpuzK8cWbHA8nuAWujPMNKrKbLjNL3n+ZrMB
Z/Kc2vcnumgIS/+npVRm+9Fnc841a5E59/f3LHlnPjaMyA0cY2PIwos626M9qDhPs+O1iBlSkxjf
2oxxeEthX7fwfFW3iDId28SUFfn3xjvOou+5UDDFiXZ+RcEzK1ULpRqlQ/rbipJZEyTbY1ed1F3T
qNz8ijG7W6Y2gy9nbB4LH16rl8hFdKMOgP7IId1SRhIe9LGT4nxOCyhZSG8F8Gj1w0uCb8Xs1lLH
fT20u5JC2oP9pqLKfXZI4Myfziust09E36+Qci1Svygz82IN6cglaiGXClLqRDqfz83ftCPLUTyL
GjkTU1BTZT4PXoRDzQU9/zU7kiHb1sC9OKDc/STal9+AG6rUkfZ/Nrue6GHGS9tgG3HY8a8/vAMW
4/Jms8Lex72tVCCPdbxAGYuyXBQ0kv07u6kSOOtDXOx+Zadec5qklGM5alqvL5d0Ahxcs3+g117I
Xu+2y41MP/MQnKW8C/5pZx6dA1nydiNTDxpt/wP3wPVAM9xuo+/+7UdbWoVSbvM1GfVtPixHElmF
yF58nIZDH/aPnr2/wYu0ydylqFUb1KEJkDxftx/v3NCQST/d+BuxM7FY15HrkWb4WrQuRsFEs8Bc
JK0I7wvanQnE1+QnQ8yqlJkaCP80TOe3Qx7gRKiQwLpfxK6MxrAA3lHt9FBdclOxOc/IKFgWUPxb
uFbx/0KL/ft/LlKHpUabdjQDbJl7HRKmX2kof6oryf/mlm/wSJ3V+UVM9PNmicUVqoPodAEOsOWT
gG5/ds+aMAyikGyyiC5Wv2q0eVw87Jf+N6fa58FbkRSHoDJ/+H+hrnDHZETJ3/636fibTHEDNB4t
FQlqmbnwpYyRIp/gl27etZFXi/cY/DsNZKx44O17f6rdE4jnrDmxK+rdd8UGvabXSd0+cXh91bi/
Z88bY8+eGhl9/QL9jXEl30qbQdpPBk39hYiMNv4TsGkVso+Xc9bZK0ZC6PlQsYbtODNTeFrmRq2E
xGG+6w9Uzjo5X1p+ZTz07Lypb4nVEw1C68EjDV1fROCoVxc5ElptjTYXz2Kg3j2OzSHJr2ByTkNS
+bgOvNnR9Bd1x3iazy9Lus/qYE9YeVU+COSWOuYUEdCzXv0uqIKyTPeILHRpWmxL3qAI+VLcaTrj
8jk4JlV/pJKHVb2RldccAO3QaCjTWlkCdisk39Q2dWbWKPqGVwueqwhrT5HYURN5d26fbdruodK/
tZSwBpYh9nt7Axz0y5MTtoc7Dg2ivHdu3Ron29hyIzhXQnCe20cDTyPn3kltk6FGMRIIRyWE+sI4
4rlrY00/OASZKn+xBCqJrqt8yXxwZSc0+pMAjyXvd85rcnFJqFvwNRH2Qv2kffJ0TG037bE3j03i
QxgcDILHdfPPynDNqd6DnHBBHr9DJmS3BiQ3uq7/j/0xoAwvo4W9B54e0nfFyXu8nmPsWlmJY9BW
KB0tVoH7pwPq+4Fan7dob3thwLgOJ+vzkgAij8du9xGk1/jvV3rWHmQzDKNODPBESz6GWMuvxuei
ikjInJTKIsLo9kKSi0Qr4EhxtTft8eXrl/tkN1xC+s7PpGE19xPFZl4caOt2MNKexy/CD7o9i6lQ
l+aikbk/yNqA9CaO7gPFWOWN+SxSG+ymsSDAeC0NDJNaUcZ+NiugR3u/OcRGBLeFTOhb7PpxkaM9
Wuh/fW8Wf862JoD/fMkYkdiJ6mGaibfh/nOZwEg4ukn1yrCOFrDHKYJ2HWvXrIR97xY+tqiR1mBR
xDtuLLp6PiXDYw6IGJq9Dv8adIrEgkaenVE4LTOYSrV/cGCqU2mjC8RvKRMeIcfoFQK/R8l/I3rz
gZrYqD6vEhDv6U9Km+raHhslhNKkN5xJplBXcpcWUEox9HST8Zq+fc1pdzUyZ8jVR1DMpQrpZY/B
ddqgdHNYqE4lm/M7xTLL1GwbquuMigHbf5DAcuX1UDTcOFLmC5J0/N08B6So+1GVF2UfkiqTdStg
TrkT7IXeWMBllx9cj1/TyFL3pAEzpsmq3GqsjMN17Ooju6vSg4W4EbTbRwN3B3gaz8z2e5Ux+Qym
qSl/gA43nVG3CZLG2Czr8XEx/Jj26+TYKusIkyuNMzx391EYgNwJ3QnxM9mNdkiBA+ZPoEb4bhXc
j7vFgV7kBTlDKmgqdVA7DGQVGHV1+A3YzjZ/aVayAQI31sni0kPIdQMKcpx/8tbod0yDxwaSDZ+4
ZuI5Fhve9WM/kZLBqoYO0UK/shblVup7yJopfrtyYKb6UBOWaCrGz+6BbHMYwNkHWZEU2/xcyDZy
CKONAjMJ7U8LfejFOzJLJnrat0R9n4FFH+7xlJMw4HhfNmyahT+jZ1zVBYRG1AnNB/KcR65/ifVk
bFdN/+ahlqecBeKHETDLXFZ7m9GOA7+45eVcG2Y7lOrQq2ti2xNP136gNjhG6VJcJUwmh+MWsIF5
SNJq2QpyH1G2W1qH4nJByzfagEb/Y2RGHq++hVluTG1A2TCCQbazaBaMCODpZTS3hHDLGJ2zWrH+
UFBp8tEn6UGSUMU5L8CyaPTpH34rmthP3+w8KZjiqFGZ7QXf/R7z/56+uixw6AJLchzNpnRlP82x
uG4Q5rhMovj2A7UzPPFCO2CW3GPxnnXa9Nh4a/brorNScMwTirqTMuyC6XdAWuCfGdA0QpsrxWTy
VdXREZ8N7RAcQFOVYYXntbKmeR84Z7UQLjDm6v5uxhN4wFHmDhFyD6saIh4Uz133LOfWNc/U62EA
7fEeb2rNOumn90dLaa0sV4YCC19slZXhEJirdVlhmWsPSIWiqae4ulZ015QNV7ImHifPxZylQmLN
TyvGZPR+9ioPcqWIdi4cQQQ6os1FaHIuH7mRe/5c4zBaHJo/a12j39lq3Ipehsz/VMjHIie5x2Z8
x/DsqFeIdpG5uv7DRAsTH7tSpJAWzmzvM8ryTTGdsRgHW9hJbrJOkg6ybIHJmNqKH/OIUsZiL6vn
XMLuuHr+XTb6Rcrmz5b32kiqM7OVbeFj9RgPVp8qOw8C0zdbkzqKBogs+OAgf6P8dfNMVV9VPGkf
nAIlm2km6+o/AM3CHu/Q4kbWQnl4WQJcV/XMT9sFeJjNCWxKcgARsIqpf5w+qQ6Vx9kkI9SmYZua
kMWV3D/csgwbGcsbqbkRuZeWpNttM8Mta9tRX4BsoA+lPew54Qp3IrwPxtwYkQEFnB2EvayxowkN
RXe200c5bqEB03qH5AXBBRUN+jNSdxbRzhE4tZAahTLiAezohBVlPTG2jPpiWk3Ou3bfi2DamuQk
iub6yRae9yzFerNjKXRpwNHXYYUOLgkZJDMexCQ3bar07VTkkicERaKLaG6iQUmnHSz2p3/o0Hi9
HRpe/pkGlQr/IHBFtxRC9NY4FGJ+RBQl6Mn98+k9E2RORjhHSS1swKHosmMHQWrL7njQI8SOr7n7
h6bUauJyXFaPpFnRnDh+iDRGgMJBbPl8f2z6Lw6jk4OsUbu6G5AeTBHd0x7+xugZULDNwrpgh8mo
j3FBvXYZqOhc5DJKfCWvGMXgn6f40H2cAplYaIPCNeTFZenb8Rvcl1xD420xgVxDuewofsuQ0qjs
AZ+MIcjBqDAe2v72Pex0MXXDRGOv54cFLQ4CN5wXrilT+nH2rZnUpBW9T04H5l85YWUEVqOMSNfs
jOwSVm3jCCChMLUQlFSWYyiHjTs43EDr+t7dgxcV5OosbPjpsdQVpIj/4xvPXQIcH3FPZ/AAnn+y
ge1cWaZfOZBTclhQgKut24N+84gSKmCSuCuxDUWrMTVmEZDGmqAmT7MzyBfgOGvICfU1AADKGYt3
Ontza4OQFvzgKvuNAeSq8KJfBF92QTfohrD59Jf7AVFZngAhESxv66jL7GsB/HruXRPHq3ONbfSy
XSfjTX1NsfaRz5oDPHuftAu1sJD3dkioHCnKVht+feCHldkmkqxVFJUEbuzKkLgQjFwsdnfzInu8
cm//53HuFcSVd32D5KbbBUVXVW5a90mue4t7SdzPDryPSd9BkPGIbycnWPGWE4mNGJXq/dbC3nff
Xjd9y+snt6oYlD5G9f5UOaiPcxrDFzNdRswhajlbv9enRFE0iDQnDpsA7xfPf8xckYVZ+0EsYxlC
EideZoZXiWmr11kEkhqrD/qdK+TKF2/SB3xb179pmW883Gm7850mCB5obX/dZEbZDncwQQe2QOoB
f8XE0Wi6znacZYkDtWL/pI+G1Z917DA9jGmRqmtjfYfS05Kh86KiH+5VAFI6l0QdK1EbTvbrMDVP
gTtLXLZjaxT6oc9E8Pw3HQfwFzlKww5kdRcCEz951qgS8wFP6O3GAMO53cRzpE1e7hN+gvBd4Xtx
zNSyynkauQNFUJHa4aR4moIo0l3YaFJZPOTIuOM1lb1GhttT+nWCaaico0KR79uWlenuI0zat7ne
SUP4m4k6eRXFwkaT6VYQxkWvMecn2FqN6dpOPpZSjH/XXFHJvZzXjUtvlzxO0iUy5HHlx0UlcPcH
UpoId+sIgcHR2RxxQDv8maZFdViFKpyXxIu5FXD4DBRIigVCxHc9DjgDleKRqa6GTwo6JTwhNZEg
QAjlnQ32cDDEHtS836GdSHit1d7YGImoWiddtdwylvW1Yasq8I2S8TbvmgSLpulw2N82zHgxmYht
PTsoj3BO3Ad5KxG9RH16p37+sMfq1xcOukjczk+OGC+KFPg2v0hLTPUmsbX4tlT2xImRn9o2fFLk
1+f8iE743xfD/A+TAjxw2mOqUnOE2PvPTz138Ks9+QC/C8EsuYi4UFWuOwz+mw229r2eDQSGJAaH
mJctXEMWGTWfn3C4LUoB5+7//6e8R0GMznM/Xwiexvm3B90v/n0tslPGd1J0qvcbdzOEyifLAwn5
3UnaoivPgXMHqBZkIBx9l6Z9Rn0NEkAMXM3MuaydD9rYA+cZunzyO2KyaDsRBRv02aVJHfJe/sfh
unmSq71vJRCbeVjQCqKItY/xdRanM9XgITizBndhNouLHsJmH9swcFOVzImQCWBFWLeYNptz/ewn
trGYz8I3WaOaigFKCZvcNGZGfU1aQEVww6Hr4RPfGRPD6ij9YnqGU7NIqXBnvLSmVAqEm7ovWyNI
y8dVfNj3lqE7Enwxu+KGKEHM75z3cJNZT4MQaoAYycfQUbbnwMbaRxhXp7R51r1K1lzoQhCgzQ7C
avpYKQdFRso4XUZlJbWQqP1eKLJ1U2GmdcWPfKxAH10fS+C96IrTHrcrNuRIeKia7OAerwipE8tQ
YUmLt7rrDoqRQz+trfwCiLKlGJsPwWlM3uSSM5OyJIuUupcsLKz31BAYyph2pcj551mqb4Kar6Yc
Oe9wEiT3cUvcIbXCRL6A/nd8dCXlVpDFpfVVlwiOI36dID2o3O4a3NBg/ZxU0mnHbf26wmAIgsfl
Y2FFePKgA61qj0lufiyJZu9fHb1twU/b7fBz2QMcX8Cg02c5Jbg8mzSbBOMmrDc/MWiJdR3547T9
kuenOtUo/IonAzyLB6B4rELMByu+Ss6gmeUeGPspw5KZIgxMHXyqCWl0Yt7kxGxstZLVhcSX4xLN
17kpf1AeXcY44BDUbLr1+PqMY18ipZhz8/u8wkP9nN0sV80GaRkQEJ/az+g8Ak4j7cDQYARNlOKA
Pkcupk61lVYEeNQ2FaPAyJgS7oBsawgUjazMRgdn1izm6cAtP++oFOBZfh15R6EhB40l4uBPqUNC
HzatXnfl700VkHdcDmOA09ihHYXYWg9txGgO+lv+ulwmmRkCJPUKs8h+Ej4+PQbhriFBAJzh4pnn
VmcDQ8PXHsYN7+qq61yJP9AI/kzMTG/mSbYGwEWvbwz6aeM7eXrqbeH0MGLFEDmmoeGOmyKa3KIy
BJSlfmTu0nrUpyT9DOaLGgSw8k/5WAmdLX9Z9W1oW7+LgZXMDO5CCbW4jHUkCkggSm9nE9fZavyq
5KmDCCk/koy/1I9LAm9OZguI9QNj6H2HVG0VeRm1wHO42ZSgEBiKYPNSnZlgHzoQeyQS5QLZpts8
01voOZ20m//cVCPUGUARI5B7Q/aW6tk3BCxZWEUmlfDcrgZscACj2TmSOEKgX9mD2OKyVlN8F/YT
x0TV/BGcaob/wYCIsSsNf3KXxPvz/yJlmChp/nwX74OiJ+XmUmKagLP9rQSXx+FlXE2YLyUX7N43
w0qJuxjeYSaCqp3bRna55rNqPJr8IAaB/Ppm79R0w6mDkeufzLFsnqopxGP21i6H/HRCQlHUczGk
91MbTjnWb9ic7t/LMSnbDw+T43NSEcDTSvVfpHLwaKT/MQxJMv1BOjpkHcldZonEvH8umED7gFA6
oZ1CmA7fZnJpZxulVyEVHy8gnOJQZ7u26hAcpl17gcnhQYBGtWYdRsu5JBQUhzSXEcGd2eQO3Oyp
12QyRpJltP1JaWhGQLFDo9TStGrpWDZAz4MR35ncyhGMdI+mzsErXerGBqWyDYgXIeV+WU4OKqTa
0Ma1m8/MwcwZBjqsAE0+n7VCCcD6Ne+SS0gqw9PiWNkbtvFKeK0/ajWlOwZWKFLdYfSxOHu5ygA3
RXEjd+opiMYYJbK3WhezE4kAAYYkyGfysM1rriPoETKU0CWtiIXGEfauDy+3OW73gr+Ulp7QWVhn
0ttfTAaq9wnqSn5+ezO0V0sLpXh2M1jmS/YSK/4xbe4j6sdOknN2VMh5iLmM/B/ddfKKXQbitCGJ
Scg5c1cZ1fppoAHxDklIO7vdKgPmNxxpsoYtxuLKjbo665t5jvU7VcFmJTvVFeDswq/2TJVfF+aW
uK635n93YFHfF8RlwxfwjQ+xTe3WnLap5GhqB7FHQLYphuRJpUoVgrXriskPe/bvRRtZLDtNWzwE
Llor2mY1ZZK4UKUEfBOooVz14gPHsgCb203jvPRlFgk2tM4F9Vse/JNeCxtftC0S1ly7qFOxaiY9
4cYi68XuhcC4PFqjHJjoirAQ8rPa4metqsCibWy+KUlh48dUgSGEW+WwkpGlzx1se6ops3QNk4Ga
44V+QQBUZ/pnvRSZvFH3N0IkVIzk81riNK4QHm9gXKlIc5mBUFBNd+WcAGklW3F5ne36q8NC3fzG
iv3+/VN8615c9EQerCwHWR89yhEqXLizOPKe/yZ4cEa27AX477QhKvsVMK+0SsL+pUYSzQxCoYBc
0j9BXjc7fiwS/5vsjiobmsMnUy5irSZAIpXyUCYQ4aC05w7iwWE2UcOqkTH7zwmnJ3lQTNBJBRoL
NWLp6gMwMOZgGL8oFFp0XEh02PhrmvhSwCvNEq8C5JRnTRWs/jA4cbOuEzPELft2w31bPdJ4uTXD
i/qR0K6bEhgtZkV9AebEBHRqxOOLdl278XZa4pO0hSF1NCQ9QP+R87o2SUUfCpWsweibT8ItKmr3
aBfAzeHSqLo8ssf9mjhm8KbCMCVCewjCWpg1VRx5dBxoIU9TgiBcKzQjgZLI3FhQMkHJCEV8tWiC
ZFQXF19z27fHpK28T2f0LFokOgUx4SNz4+CFO/GSKSDEvxtqpP8Of3tdo69lvAkqEpMFwVj8aKFn
ykU1fSC55hrtYrqkq2vVShuGonM2c/Lafa0a8B8UHCLIEIBUNBhucDKam+mu8erls9Tge3kKmlaj
ALLgx0V9SWcncm25NVRjgYFELsCpIGLPGJ/oM5RWEmZCpYAM4pBENPvUNjLWtp79TAQGJsBNjCgL
7CVKyz51XQgyQSYOq+UiYT/mRkkPvd6W5Bo1yx87RSsD7Za4Ee6xAQLQoEu+zogLSgKgaMfvUyk/
pYsMpsmSICTgIorRxNoYaJSTxcIbgqxCE5eC9t9gTfam34NmQqhohggHNixM3+p9euMSPYg8Cat6
al5XxaUi/wCIFiSisGlPimrwWB+x3m2wwoOx5OCENUSgahhcF5v5xMIY22RX4OIPq2gB/qlz5gll
cPWI1/4/lGDuc096WCWDzST+IdaBhRTpE5VObLQAjDT9pgxCTEAMkxAr2UIfLzo+6ETuNPeUsRQO
dZXjfpDWFZN4w8Hi/tu5mL4EA8464i/DPU1fXeSnehUyQrsudhRms9yOJyg3PIY/ZdoqY78GU9v8
mRFQYpyO3DyTxooAtYOLAoGkx4Y1TSCe8qd6oc7PX0CkUFdDZjCAX3ijH/g7YnoZ+RjdsVzeEWqF
Sh8NkypzXMypia+qoQYJFlI5JKPXyWW8BnTDOL1v4RJR2ja69W4MXQPjwn1/dXE2HeYPypAGdbHp
lTjl0L2lGgOp/jMqyf669v8Za91dH2PHqntGtqFTXxDP492Ch0tBbmX6zCk73/PRuYU9H5awkYiR
T+atdgh92dZYPDom09TxjAAqsgVkbArEgwVx6gqPzAJ69IwNpzSmapI05do6MNYbeLUuPQoZaHY8
4zrnVrnBSddq5FRDdUwCtD+5nn9++R0TaLqiGBsdX1spT6NKlznUiM0PLPhWu8AQDyfP9+9Ymep3
dQIPB2bR85wajenJAtYQJLvJtD6p9L6M4toA4SaR5/KGAEinDVyvyQPXowYj8m+Lk8cVsUqYgOy5
Kc0BvKH4ZBAKsRttccsn7L1Sz5N8stH2A+M1vc6JmZjJrgjotCxbW+XLWjGrglFxkLCJ6o3ZKBRI
6y8LnT/hen/q6i4kYwZfzSTB7hRQsfi4ucbh6ik77xLkPh60tlIeuIeqZ28oCCEZsW+ys4SoXHFQ
B1gZr0nAc/lGHmX0L8dgQMPTKOfOeNTn9PgmtCbwGbJO8i9sgRwCseqzh4H6e6HNp7rQDBNSWPfi
nZuGXmMXw3CNJS1AxIOqnn4hqXN6U1unth5XckRUu3YaV7p1vMmcuc3uApv4OBB2zQ4mYSl7yoX+
fhk6W260PdquN2/XenrAqTpH+7y6lEdQkg0Kqxl3ZCW0DGSUfp5E35UkexpttZe5Gl+HU59SAKK/
LJ25e6iiZA/vFVuUM1DsZDF0BIOTtBKAD7CLf16XwoS28lQtwmMQTDjQXWP6I9XT3ci4D5A6xZAZ
y09iMCjm826+ZkxIN3l3mirXZ3riVnwSlxysrJpOOoXSaQ2fU52XrRS29v5IkB7Fk+BMpXOuGR77
R91v7wk5mqw9EplMfUwQAuP4Kmnsszc8q5EqzFyjCITg4Xs0MWpbDEhg1KiX7pP2w+64bGYDet2m
YqJn+0ePCqhZL44S6CaOeYXCZCZXWN+YclUbSHndJUwsqMJtWTWrU0AxXkTsI+HGWHz/c6aJyXmp
o0W7KLPjbdunMmimbcCpQcImUtKRTtSjFLgifxG9HhgCRCo4JSRSXjrIV6jNSTSLHN7QEkdF/RJG
Plhvle3hv5vOFsCx3Kuxt7LswNYCjHkRLDdw73C6iOPC2coEO1vYPSIa5DGRzDtyGmigAs0oFJdh
V4dIPhv6gv3fx42Zveu7AMNczEDIXxQRpBCiXVjcxBA5Y+D346z9TTU+J4/Uc07tAWUWSO1Yp8/0
hZ2N0ljuk63MquUUqfgtyxVNbZIbxaAcKuNVZhBwS2C/GTI8FhUpSollEOd61rDba+/hCDTPKs5D
nySfMLjOUNR4KYpdrM2Jcu/eirUq8zdVb7v0KMymC/uvX9bxBGso4ALKwzYIhBnYRhSZUdKJ/PZy
4nghl8kz57XyX8KAvdJYH/TE5A1oTF/vO5vYsBkNn8r+JSu4RA8UtGnKnf1Kc3AeeEdgxJNL85H3
WXA5pjaRHbNQmzZU3ppTatYxGOICth0LqNapKq6HckS2YU8Jx/+eOR02aXcGcWWCQ12+Ln2cXnnT
DX9vmZGVpnGauc/jqojhDrRauudq9sZCrsUCeORICbSQcjGpi3DIaD0os5hW1r+WtHOgWdg1wf6w
jwrGBLCA7gChDR2By+HOP1ZLRvTMtl4jwqOpvx8/mhXEPASsEiK9BxBcTiI7Ar1oVQg0G4Nwl28g
nTbCLSqNBpdiU+fWK8DHukB9OflQ6UV5XpiUsVuPCr82yL7GVU3zg1XKRKWjayKSNCEt1XmxP/hT
vnGqjjY5QNHhdVLmkg8JAF5L+nbT9AoyUyQBR4IRpITlvs/MZeDNal1yZg9MErJuc+kzKFaQkX0c
hRHtObXZwBqeGUOcjKr5m+0bq23r4Bb78S700QnOu2410HmWNqRoQQupYBaOMT9W0fTrFyI6ROGC
roJNhAWxqoiMeCGUKEewXXuHmUOEGPvA3aX56LA+pv6odyFO5fDMlR7qxplwBvKcR5/6zQIiFPmk
JyqCqadGYgdpLAeOQuH50MHrRxdeNlmdYJkr3CSHuc+ZC46MLAPd54wXzYbERi8ySxAstllG7ExA
0pSsd7dS0tpt2wdcg0s8UVra0Sa1woy+T0ZM3nyEGotMxdjH6oPTrIyo7sq2WdKImz/HkAnGpP6L
gy8kq9Lhkt7TDprlCgEWmWHZahZqaxLXUqlpazvBCaWWqPUD4ulyRE/d2Cavm/+W3cy5NrjJjYSg
OueP22zfFU1V3nCmRF/gBtrW4Xiah1bHTuyZyyE3gfNYX4Ii/i/VoGM9Yg0ddnjv6HfsxMtjxxlK
CM9DjVeipDNt/ALErnUuP27wVIi557QXxLleGB4EG7Uea0sXn+BPVF/q6NV8SbZkpJPRBVImC16x
LVbTFMeilveQsmG0w1Ty2KMoPPL7OPGwiQFyP3a60YFPHUqJbYQCRqlV75Ia0Nq7RqzoxRUAbfwN
j8R1kDHyVCvokWtUJXtHmU0Ddu1BB5FkNP0LSglvxIyu19ycSFAsVNby+3WWxaZoB3RMmv4XM4jt
yXQBXzxlpJu+ZgZilyOyKVZ1uS3fNjXIkXBEYkkDSXOPGfpNGasfojh8dnb0VNZ/GyWtygaobr6v
iKWNxrCt1/z0Hb0TggpiOx1MfOreP4dntNagmMXSaX2yo3wwKhoqkwVhCQWAQ8VeyaF0qr8YCE3/
WMEQXIy00LMURs1BW9aswjWk+xadauuYJM+JfnxHU/8F+nqocTIJC41SpJztt3pTFl3QN46jZZW9
n1Wz4nmfSkOL64z9d4KLftkKnYHZ1Z8+IcPDBJSmJC0Tr/0SuTqrx4gkJlU2IsZuJ5+xvLrwXP+g
o7tazhwiGvmwl+qvN5S9DDGrVwxZC0rj0GRzD7+duXw7B1vnQNZyVJ2Cd0XSlRQ7kkct7cy9AJUe
fOdQIosxBsMTG0/KlfnEr1OB24HWPQvmp6ISRfDNRYhAEQ650lc9MYiMwBDEi5nqeROxzHy/MZS/
e1WDlaxFgFG3nlL/1jMBfhFNjf5xifibXbRMJ1hhPEUaVoZQWuhbU2HcvOnLWusxGXzpAlDeUWXX
yTsen3RTwzjf9npQ2oy7QehuzaMjD9JrsIkBQLmFt2H1fqe/XGfzu32vZXcx8+AvASuCwxv7QkRO
q+ddAsqAvDzYfEDIoJG6Fp74wtwfrL7ZF0WIds3J4nwx+VcL+8o+4EwvyvidmAV9JxzFNry9flI/
ES5ucIipZpyIF69y9eEGtzjj5wWRwziZpkDVcNOjv9hqlFE6eXGN+xLC/18KVCGQsH5YPp3zx3zn
1dOMF6O7jsALgO/B1a10JiF3gCggmxZyJ9MrjJLrygwwMq5UbjiljmdggI5wrSaKlOjvgkGSrCYt
onpCmerKK9EC2/L8yKzAEgtz/YSB7GJAjPEwU0mz9rEk2JksFfo0Z9Jaferk5AI7/viGH5vgoe2/
305SqvNTj6gCseJXC3FyEzF//G1lyOEddECGGsjZgiQIThvsjCC/kpu71QDEQ5BSRqZqeQq4utLK
QszggxG1JE3098Jjwdqz3NMYqi3KVhTOLhcMoH+5eDv5D9zhPLqZTKYw1pKbvKaWyzCp3GYhiXVE
J56hBV8B6v5Vbc9O375zhu9+AMUKVkXhjar+Vikg6x9WltO7sAR3rqhQHGrnQjcB0rYjlgMIc4g3
lywCOkdWJJMTjqKsiTQvE1pr661yUngMVNQcVMqgGIsdLSa08Nl+JkrkksLO7YRPZFpoNTQSNtfK
svvpd0EqaocD3gshkxT/CCHN9ivlozJXcb1v1Y5FbyUi2eui2wmBtf7OpgegqYq0TD5whlnAr3bH
LYCZ7XucElfVRQrA+a5ti4PyT9zZric6cCuIBimzKIS+Dv8aVONRzeY7VCGbdEK9VT2iv0AxtsT7
0AYrkDzxzCMWUFcPikpIrBMyWhS/21jZVBtPMEPGyhSAqrhaeony0W6/0x9S1RXfuaRNiV2UEQ/K
ZGE8PuX1kE4yLZspnEosKvJHwHcWBoHQ1/PLDtFzPubCPIQ851/G1O4TnLjp18CodfDHCyhK15wL
CqUDvZK/gMvJAaP7YRB7qiNvE4JA4GqKwr1wp+Hd5jE/3psU6QK34ILfhDw3PlHXP/hrgmEWBfUG
eyDrIKzjPxp8WOcngBi/G8E0ZfYB2KJZZsydrgVCggiwmiBnxJ6azUhK1E0dTfI7AOhlJYd7V3DO
8FO19DiSJhEvBHWl5J8c4+RDq4II/541V7tUeZJC0G/tyoHsNZT5a+/CSZZKN7A2HfwIsFLxGxwb
oPxe/3RtYXEMJm0vdey4tgvbdAMCK/0kJCgu+QbJomF/BqWx3TjPwoKUWID1wQpZ5m/14LCLr0FJ
ZZUnlnhtr18GMBrCKph+m9LKxkV2YC5TtnIrwaPe3dVNAw6GQ5h4+TkT4DsvPbCLSrE6WdMKgaQ+
RoP/ArnLRpPwWBHv9ikPRcSGyuAxHnw+ByKzG0/WHjiKZ4s7szHY2JBvPapOVW3xkuOiFQBUsr1o
dMrH5yIHkfVpsq04W7q6cW4W9x6xYOJDdOD4/F/QHPFE1fDSklxoNlRLZMNmY1m5AZxplXntM7xR
2PnnUOPP5rNuB7PSwD8sGnn2OKKizzOQnzwpx913jjH+s4TaAgjEaqx575wVNKuVV2aKhm5mqrg+
WV1g+o155fIIaEdWQmQ93CJTrzMy0hFaRnwV1GqXpk5O+U6+RSuuJ8+N3pMrK4oelv+gcpYsgAnl
VIQ6Tzd21dbmWYVHJWl3QZip38htbRdVHEaW//7IUCouLFylflkBvEZ4x75qD8U3EuujYa7itsFH
RCtQYyQNjbvOpy0gGyakW3z0YNk5t4n/WkfiaEb+EFRRSIWWL2gzlkbE2XSP38aIU0EmEkJFj58b
ZJjs/AlVZCflnr+a2yxjgjDc29hvqIhePNwVa4ulOJdn6cLHv8qLVM8DyRw/Fi3lTCAqMOZ86GVk
GFES2WbdVY3chsHEmHDN6Y07RB+M9IeSna++5obAAyIhJA1uu+wXJC/8hheg1kcAZFgrXVe4V/8u
0ODQboYP4a9B+Or8Xpz7koz1FFpbexmypZUkvrpoAlDZIPwwnyODlIiTVH59RaLUq3jNc4auOgmy
Ep4lUBSmuC1twAp7ro9qUyqMtodHy5algXs4TNjLvqzhWisXtRgrcZnVoC0Y1joAzXlMjXqOnKwU
GkEduJDT2LFP+HIcTZBprlg3kqNIlK97W9aVlnpTURC+cqSRHRYL0rbH5IFke8eljNCLELU3txV+
wHzxs3wuj4EifPrVuMkO7+r1xsAJF7SCHGv10arJAZF5OUfeqMYhBdH7u885kHB0b/1VIvxhBNzI
m1exudq7NcWpWlrDkdEZylmdbWgTDnKIM2iLmXqI1N4K41TYKt/CbvQr/R0W+7XmR0pM8ygDzk7k
PZ0hYRsS0S74JBnSa1Z5B9Ke8GkvugiIbwienQAjyEvMoHCNoEm3wpNuZ34rJTSOifKyryE5Cid3
NrJJ2CfQtQ85VfkREhDFx+PrBUVjeVoJCL7SXiHp94Auf6cTmPVmyPSxjzqFw4kNqwkBfSLl8LxP
i/Z4A1KsLyOpzUhWi+AmAatM9p24jq81G9BKj5K09PiYoLCA4BXdo/Oa+5YD2yKyMOsw2J0ebDOJ
vp/yHNq892fOVuwk5dEItmazXuO3kRgo9vLcwYp15mUvwYuDm0Bw6fX0hSASDL2HdY06GE5Gz+F+
UZdomAa9pk+s8EC0F+JkRGi+41nTp1ANw4TbQJzcpNA84AnoWdc40fiE5zJyLjP4HeB4++O1/87t
kR5GoGVEL4/slcnd949JBnN+4hRy4qQiQGOUtHUHgU2fhB98fHoEMxWEaxPDfsoyjGCVhJZ9s8Oc
YQ6Jo2jkewrkKtbMixliKqRHdbXFDnjAdltnMb4c79mmuFjtHdqNhRV+fXKLZjyvf8WRt6JlbQKw
KFOaYqoW9v7bLpxnqN2Td5pLlE6MUfangmQg20DnPxCKim1cTgaH8DrevKqkMnD1E5tIJ8qSCYUG
PIj9fluB69eQk2QEBUxy5DDEdEf+zpGOwjfUU9DsjkhwBkhQaTS6rh0R/yBhtIr+0Os93E5oIlgk
5H0ioTyMl+r7UT8eMxpdrCWIA9oElqXEltTXQpmVy044cG/KuM97eIJJHtx810ifaqwkbsk4/1og
3AnNyPF7YQXQM1PwgvWdpWAV2xaoML4WQDH33AyG4bHPXWWWWnktGtffvqxez0LdLKodXCqqHiSs
RxNtmhm8jzKRkErhEKi6XLtblL/pMOUDFYyP3uD2Cio79MNPSSWcw4VClVdUnUn6jrl1jnPfaF0L
eX2rOuL5NSi3rDpUL7WVLfAfaingLkJLQp8CthAFv/oovRmrgmxPg/Xw5ChCTuOV/o0Pggy8c8Lg
tqwIw0TnJBE8Ah+SySMXzGGfVtofKVwJbiAJoEu6xENnDJl1qTB5l6pPONOjOsMuQR5jucyDFgYV
IqEF2c1bWK4nrnSm/w723D+8Q3SimjWFQrMTEtEr+MuH5SBTVe5WMNqtw8DXOBSJKfNeEZWHcbcL
/vEVTTdywcoCVQfkDvYbjKaBfo4sJTBEgkggx8NV0awOsPlv9Up8rSDbHEt0JPTjaSo6DTBJG/dn
0vFOhCd4OGBRbAl5N8DSbVSis2vyQ9X0xECNMtiVz+ePl0NDvpe0mu7LZnSsgRHqFQrRF5KhK3PH
HElk+s2auIM+G6twikFfq/LmLUrcE/OhqYZp54rYzhPCoTZAKYm7msdyVPwtX5xapTcvchw/Dgmo
6oFt9o4uo+GBtQK00vidUwBKyORBFK0wNA/BLbXojtofOdgVKoTxFU7YrFf+zWfA7etG5ffGA9Uv
FBqNIabs6cIL1VQDA4w1Ygh58lguksLTWCmOKOHPPDMjiFF8U1FfF1l03ExBSUc66v+tydpi47XA
mkQ2eX+8qdn9Hh/OYqYHIeWviAQlao9wSbHlSnPTHmJEvMmIV/oaCwWN+8Oh8lo33ZbLRQxuDk66
mev1V1CL5SANCr15Fm6H0jSipW5NoguEASgpsZN6WUzKBuAbu1p2X4Nr8Fkjw2nsLSvYFlXgSuqa
2OpKpUkwZYOe7ftslG7e7R1OsGXViIKjrsXKU2WtfHBZwJAbNKJnGOxY2uXXJjBxASwFaTlMVpUr
sQ/VkA1ycAQ79PzTPNpFj4PEzgoKqGoPKUK7kqwCwodvDn1b8ukddd1tMPTkojyFNS7Pc66xJJp2
Ji1eezs37TLW87U4Tx/yO7VobVSZSckhxj5lEgDIaB2LpfkgbcbZOBHPnsG0kEKI70Ef6vJhbJ55
sQTnHRu6reZcDBM7BvuLrck4ikfI5yGHSjO2UZarzioqvuLizb7Sc6sM//GzdhpzRKmQqJZIazvu
CPMwPABTYrmFr0Y4ObsbWOhYbFeBCfX1qyy6Q+CdJ208HDMA8R7itIOvXzuuI+Vi+JBvPKFGcAFD
M6UNHqRM31Z23Ew86Iz+94oLWYGjOe3Zlbg4zz9b5hKICqw8itCZmK6/atVrwRctrVIvtqczEmZD
ewHOt097WgqxBQOVWtx8NnNTpkPAxHCHv0v14Kaqa945djMx4wLKT9yZnpH9Gyo8snjb3/EXbGip
DdnPU1bb1MP0yNT/CqpHchEhKSnsIe/ZkB494JstE++m5N9MwrhDnevipFJ5yhTa5GsSEEzdSCZ+
63JcCDuigLZuBJNzI5+cAh7URnaQ0lqae6gsuq4fZ0rzPs+MwgmOlk9thNdNwQMeQhpCvpwsk/O3
wUs9GJ2BbSHdR38PJhaVw4sRuxkW7dy2eR8ykTWQmpYzC/8/Qv0uk553W0RxzKTxioZ1dPjfJLKp
B955E+1badS6W7WPSg38ikbVKgJEOQdWH91KsZGuvse5TFspef12EDbbmQbFKHCSmf44UmRC7Pqc
qiLEl0aB8LCuRQH5wrcYhAEU0amwczb2GSvJoq8R++VJAuVUCrCNerCl40KJu2t6gjNcZSoUT9wt
nyG8z1zV5jvnzzpOlfrMgG5HFXGTMG3RuKgWkaBHhnaa4iGngHxHW69qShL1hj7lcFwtn65c8NbW
9OpDpFUEJd3BXecXitweT3KpfO98U+DFlRSudyTSrhO5c3XhECom7GjSa5LO2EmIdR+H16UEGejY
0Qn6M5W3wgwb+IVIKd1fgDbtL5RZ0iktArklcEI94RHDhg7IjNIWVeKkzDMWSo5maTcZvnHOwmeF
MKt4OMx/KKVfF5CHzTu2MSheB+6gieHdw07Puww/gJOhjagbc6OaYxIGgKqO+jOalcRyg8+Umxd0
rN18tm613OSdaj1lRWpuhzMAWr4VsZRurPnx4ja+EoUlLqJWpNjwqOMEhbfUkMP7msdGlv/f0hxj
Lh+CHgEdPUt9UGQlTkrgjpPpp6h1DccL23spNeLTsHM9F4aWdCT7YgQwyjfVXFaybrM7U5xDz0SG
MDCjX87wfb/JLtKp7Nj768oM9h1XxrbA0VHttuP+a/7zWSGUh7xPEscWwus+MmpIEvHre2nBbu3V
/sQIq9q6CQE6IwgwXmizKxHDNVw04LWe8XOl6cY4rFr0v+238FrTVDIXwofEiHCf8JzMOm+VsYuJ
Oxgxe2wGlxbr0QcVe0FGDRK1WLZuUmu/PN4ga3IA5XmD0tKJNttrk39NmBiOAd6mHaVWP0MbtPxr
G/PUlCdyO1cPw7CvLU0dsm4/b3GlwQS59q/UgBr+iv4hH5WY3yjXLzUapqr6HCkhlKlyQFKJD6az
zgfZKlN0OPbQEf/y2VpnzsjWHp6MNIm/MZWc5V4wXD1aa05Ta5eQ51NVEn72PY3bRc25SfzIXEWJ
dOHAUIh9biZWJ6snU/pRiRMO5paNAYdl8MRvWmK5485pmpsHQx0LV+v8X0Xcf1M0UEgQSsadzahY
Ck22JBgEodQ3FVaq+M7cZ0lm6A5zOrFrKQuD2mZeuYQWvwNEKytpDj7ldUEuCmggwkJg6CMljl/G
raz7VYoKcxydZ1utQ8TB1Qe6b9we9XT/9rVNTycFw7wIylQGbUXOL2/MUvJzjjKLFqI0rqYZDBFJ
v9aSK4bfYXvBv5OOeQcVMy2ucyxhKygVV4O/dszuACU6ytAs3pNEyMa/vsGC4Rg0fvwvO5dwQYJ1
ojLJoLlNOw1qOajV5dzhKl+EJyhxrPnrRIpLNFaBDOn/c2w3CbjZpzWrqkgColbGyn/4Q8sxS3rf
DnqywZ9tUrSB3Y6dgZ1hn0UVzUgn0dYd2/VmLQ+diWQjEGPgjYcmWzvyDBw6/S+PzII4gUzgnrOF
d/b8m9iNglsEnyqPcwW1nQVehAsI992YO2gsbdaUP6AqJnQ8UN1tPYBh55z9m/sBcelLmjKIaeGD
qzbPB7cAOeAA56GrZFWq5/LKyxH1JdfixwCEiee29clcMtyOUrhXZc5McUEI6dn6FAeC3K2PkJ+X
UKPtiFbbsFUP2m4bM5U4i8jAn+DMngmY9GSdSpMi34ysIFIgYojctC2ug/Z1wtNeZ751+DSRA//N
SinZKuCvbC6lfl2hM6jwu1P8CKj/eAe6URF6XbvyBOjDhRJiD9FNR/aYYVwTa6G9kTTm1LfzcNS8
OwVc05VTv5IF5l3q7xVfUoPM69WG4DwgYwvzjCqwMq18heKIsN+NTEup/PB+r/uhE3DKvfsSJ/y5
egAcRN46ZRph+gL74x14ZWy1Mlihr8k/5lnM9t4ACvmYIfJD2MAlsoSQOPU/1AXhkijUfYayFGxC
CCsPF6ZaTe3M7zx2EGNZo9Wk4pRclzk3EZvVqaT+Rm6A2/pv0KgavLrIvVCneIvQ1ku+j9wbZ34z
6VpCmnr6xIJHkiOAZVmMpagZTZLY1Jv4b6oTF1DAKFO1M6+S6MyMqZxqtZMcF7+zHGvEWoTxECbR
ogt5iW/MvX9NlvD1FpFXUWTmoTH2j7HnvBkw8fiVMVCZe00VFCN7FUbjSzvJ6pRAZLkYPvBs3Cwa
imS6xAQhjPM9fDQWi5d4daPuQ14YLtgzMKrm0QlJYANKQKQLUcJFSeq6SJHuU9uy33dfGGMnlqr0
vZ0XkfqCyxEk3QbogMDlO6p2OzIHUCtROVSwppMGBnVBBUlc4laoeH27qaX3EIJ8qAOQyTbRrKjB
UaBfo7m1fNsg3zThnBKzG/51lvsbuNschxFCUKfVWVHEKPn/1u7Uh4ErjXiIdQlUQ8eozv0vUPjH
r+Su7h1LdaLhHVNZLsEwXGCPE7ZoanKb6fCbI+mCLJrZ1xvK+sGHMG5WTwqIOps9MiPr1UtjwgW3
ivzPsb9Rexq17UkPvwlfv+oOYNwzwb3dNNWc/BRimm1fPOJzkEwApi5UDaQkwh6ffCH7cwAzHwGM
3tUU/yZgozFirNhl9DvepMu+E/eB4kEL9LGtuayt7xllL6kQNEYQ076DnmMNH0T4xX4PnqS9mP4N
L/qZ8qQCDDTDY60VnO15avxYVrfzDwv3HkaZ2USkwrhK2LUSs0NNVrewsY+xZPYmSInbHYBy8ZNT
rO2K7kddENb2Scb4pHff8OFU2H4Lea+mo9vOkkDwG/qoQ5nLI5SYmaH/2OrxSGGS/2v/zyz0WJlM
21j58sqd3hFxOFuMWbbNcdiFMkngHKEOjBNBRlIb1ugkUAMh/G9IjSniBjZmC/h8ZKBZnfyrPxyo
5yz8DKFkn9PqNkLvzaqSBoJNg5jMTGT9r3NzXJd9ZXCRgKITuzKSufMwLyQBbZ3bbOsfl/MQnSpo
+oMbdzLnFVeGENvVqNz6cawQY6qJrlSewqErNecGBpT67VQhv8k/tv8UUrpUXpjxljJo7teyX+Gc
hT8LVWMp/QtK/M6p6cLJBnUVp+Yu7uvyGlXof3mORBYNUv2Zs82nqIbLB4g0aGAyG22UvuA7teaR
SgOuXYmNslXgNR/h99wu6xpjGRpH4nShZW59xOZLEhYyDwG52U/hwGlVxabarYQDefGLnYcS38QA
QyBW1B87bC2yGB4N2wgR7M5wV69EFAWcZfUZlJ0bdCxORG2mWLBvVh6RGojYcPlLHEtc06ROsR6m
DZp+WBznVL7zbZv0oeTKgEuu4lpU1zgGgBK2p7u38EtNawM8AzHgGf5z+zA7mcqbvnRqxl/Zg7Fi
hCz2eG9CrmwpXJYeERVIQ7idKKtM4NgTbdLaHYzSPiVjAewkDF0c01Sam4cNsOlcBuNQ64St2dYX
HVK5zlUzEFi10SQIW5G4l0JbVDTr4ywXgGFdHRmBhgE4xFBJTqAPqvjDpcYSIfB+3UzFG7zWNccH
U7j4rbAYhANDz8i19OTR1Fow/kKhE/edZdoIvHziqwkUk/XBorLJCDxLd3mgdXTsyrl+r3u+VzUt
AkoAzFCjGwiOKlYgS5oDpY+6ulxj/eqEE5ZQChJtYDRiQnLkUH5wfGe/SZNv4swhaXjO+35C7ved
5JEDBidjnU8Yi2r+gySuRcImO3WxNDVdu6jsAKq8/t3XuCpo0FEUxeTiSZj3jIIwpV34n0cxYxaG
jtn+83rjA54cSKkkm/CVEw3lM5Svo08RrY4RzogEjkzHh5FUWmQ0riyjBxqUpYSdjf9rImrSaanw
ewbRvr/ovtgXFhaMoD2zixu5t10fcvEc58x6rnyb/O6nTIG47hsu0sZ5QRUxVG7l/O5i3oofSxLk
sq8Jg3WaruoDQnnA/XuqQh0tqaLIRtB5JCcnaqIt4iYDcRo2JwRgKHOILqs9C2hPa1SWmWosQkq7
xF3T4cbDGpquOGhAlh/7OvBEmsJRPvqwZKBCMKnlfneL1QEq+fItfE3+lLtfCSOEIla+OoJBM10c
koFGmPDDP4ILSS1s3xNAlXxPF8o7+pwq4sR4VMWV4ZsNUlTOLCZezOq5Xzj+/Y36YkptrPhIfFGm
wGKXmrCcpEavnbd4T7E7m5A7bEesd6mPuu4F1CtwFOGeQxLn34Z9i25BVH91CfasNRgR7BEjX1qf
8ucuuAjvKjQSK14t7JqV5xkTnuGWxOZImCDy8TQV4fJP/ysjEMs7YT7l4iG/jZmXIzjn/LcBTxeA
oDcpsSF2WTpYJioan0jrcY26v6cvOhSCZKYuE8sauDiyCr3lBNkYgivZci5kQa9NvsA66uFCVInc
2fl6hO2FcfpBCs10VD9/6VZG/iR46w1uBZx3TK8KiYY2yG9W3KxqHGjBgoApyomIBf8lrDnEf0p8
Kex5cSrs9Sc43HQg1kpgGZUmVBy5LEPVmOJFE/RvJUsGjJMoMnhMeXrb7Zfo+Gk1wYTUl2ksd8r3
iAUmWbdOLHxvQ6e+6vnMNuOT5ZQllNp9DZB1VBdIGv1vfMP5djaJPOves/14dKqgctUvtuPN6DgW
qertC8xdQSumSjBHu0VR7sDu35keSkbEJTXZzFEetb8AEsy6ACZoGfM+zRI76r4CMhJj/cwAR7eU
leZQt7SR1mHSPV3bBJ2bw0n+2OjgPU6aOuHaUpwG7atr/6Qv6nONqcnqr5BwJQzCbJMe5kiZTfoX
FL4WeYgpZ6QIl8nE4TjRR4vlw8oqd1+Ux56l/acV8I0ZnUoCbGls03vDpveGeEqUWzLEzYPiCu2H
utM+aGWANMCm+hwYx0d+0ldkacCUAqeOiPrGP5h+8wCUnapJUAf2EbAdCa0V0AwRJLLfDNvvxeaW
T9Kl12Vn6E2tFlI5X0BIzERG+TdjwoBc4xoIuinwEi7PvahSrgRI/+CYvhqc+KD6yM4oin1dyYPE
HUWbE0vZYsmSSi9sIVA+GN4+2Ikz65276pB80TEumGW4zk0S9o796h9t9IFcTLXyYauDA4zDxAxg
2KTKFT8n4nECRGe9RloIEVRaAeA4POExxbf01B/1hs9Fp7V5n6+w/47bR0eFUxnFVFVOsJ4bdTMD
BXWy4JrUOK5VFq3RDCTDf51VhsGPgpTDIcecem4QI66aM1PKx8umsZzG/Eptli0fx/UrcDY1KfFW
1hkeyImsiYS6uHWwcAkfFA1sTeqJ35EinaZrlFJEHDASLW8EAXbP4PdhQtNTNe6i1Xy/D3lGcfCi
kw1v0x0+f7V8oB5CQfsi+9dHhLxgbxRHc/4K5xwBalb30fkODDWzZ8tTLgZu2afhLR4PmdvEXwhM
G/JixYRTHyqrtWDcmhpAs60TWocVslqpcqBaF6wiR3GDdHT7hgsEpYE8N3J+zO39JDS5StPt/FNT
7dTRDg0hPww35U08sZrWw0AcewHN5Q4adiQmIOcqD1aNV+ofFcNFeCHu4tgZshUpL/FBQFy/wBxR
IRfvQjBzHe+36MJTpiYYwoBh7syAQ/Yh5Ti97hr7v7Thgl5sLEmBTvWxUKirJWhEMHhUJbQqdo9K
sHzHGO3r8xA+08EVGVnMwPtW0KwY+vyARt5Wia7Q3G5EaGt3eVCEEcFnu+65EV5iZ1VbZ/9eDmdP
UDVEF+5xuu8LuXaU+7ddQWMFnDBm5ihPO429UN2xR925xhujZANcXDi9ctFq9ChItG2Naza9mkO+
Ry5HDmOVwkZGjvRbOW3UcCfcWVz+5UPJ17wtUFuc8ADjuXdQX+ygsz+EcJRL9sn+FQwq0BYy1txW
ghxvO9ngxgXBzRfQsJxl0fOIhO3K8gYKzntP4w3y9dL20sb6WzzB6M950qAo7hZ448pv9M44ZeFj
7a1+VlkGY/Up3BIPwTYXt2etsc8QeKVy1PPAFCoeMmTHRHXPr3vWXMR79xrPYFwyVL7Mhkt/DI3Y
+eYGTZOdYIxFunaip1yNH0qIwWFX3SmfZN+pl5rtsSgdkrygAy9K8XS4DtUFVrc+kLfC78Pd7Lyg
e73nUHp/kz3oddEmIsvMEpeWu56OBwbxHM6zuqS7IovOQK3Kee4ZsaUS3Ws3Yzod4mkyzbb10n5B
j4EchPGUYPhRel/MyZa2f5AJKpkdzT/ducQ0K/wdczRY4RLqQj9laRg4qccmUVBYk9ZqSMcY0zOI
5aYg7AVoQfNGvInb9jrhAdlr2WU95a824FAkvTcfl3H97juRbUmBRn3+wIr4VDpDZp11oMo/ypt2
nJoDjhwDyZv0uyiz4DicTubk7ZAEvw5wTUiQIi6nmZvAbeVT1+XM/NtdPiwDQ2td2TjMJV5AjdZ+
2tf447He1nK47WbGC0ZOLNaQBKBNjoPyN0E7C6s86D2LjS33Mf8CZr8e7Bdupxx/gqHCfaCX4agD
rKzBBvnVX5vnpbnr454hDoo6+SVrjOibnLvqlGiaU7GKvCgxbFiCJp6WJGBoY1fgfmbtP1AwSCkG
036sdtWyZUY6LmzGWlykJ6NU3fshPPL4gRK6KS02UifZK/U0MLjH0T5TgC/eYgTJ5PLfVR+BRHid
LBg84eP1GFibWZL55FMMGneaM3jCUO2sbW80NlBjkuwbYNsifbC4C9cYLTri4aYnQRIDbZgU3lur
k41l2j3L1Sq/u1Qy0RpzIFd8Kk7+KMaGu8sw4gpLW/Ls+snWJdqBdwvH2+TiG+rWTXFgjv4r+ffg
jQ4rW6mLy3ppWRBE3BFx6bMeiBQa8nZ0GmnaCL5WlwQLf/H5kQNAw9VTdONtn1EYUaGA+JmNXY+6
JbUGSxEWqU9QwMfdm1zF7/l5cS9CF4yOXW98SvmQIrnjE1lgScenBx9Y975YjMxCz8qsKByYELvo
XMninOWhXinN7/+sOZGUecMDegAF+rq1ytflnZ0GDgSCDxiQk6MDf4cDk7eFNapgTCHFyH4wtdj6
puw3v2SsZHVy/scvGzqIuI0u3d1OsR6zy2QhDmqTrnGZqg/t2eywUlOggPjEhe/LZQvExfMjxCKM
7IJ0X0JMUrWUoJUPuAqcqBRbhYkEwCXx2bOdmPW5iDcHq+WijAkyUUWuDHwn7ch5ygycMWo5sMJc
iE52ErHJCmHUfLh4J7ghHMQxRq+mLm6TBufGJ/zDXuqvWqDzEeLWcdkYxNIsLamZfZl7NufcNwzk
kQniJpvNc4rNyo7iw6r5VUM2BS0B5qx/mPktX8LB8i028kwIPwTqeIk+tx5CnBlNaRyuxbNr2lSJ
4YLMxgd0nbD+jJ8eKNAfOX2gABJbSUlFYbx8Zitf1Yqvc+oIDLhBMlPb+1b5xNU9JGs1v42X0caY
89y1Z6Tl+GZcHwph7c+eHDsSRMtZRRGJzZRI108WrVX9qinc7CgQuEHML21An6wExhTtzy7j/Y4o
IzCu9QPGPar96F2mgl7R2sPyEf6It5ilbNN5RZCGcLgHRWIg59zt6CnOXqHdkiaBsiuWBjy4Ls85
rdWk1Gx3VSE3qqH5IVv2mvVpCl8d34uEd2Za3lez2HS2Nwtx5535ZwHT7Suvld77cgZhLldbno1Z
xRS8WDHrLEDhK+hN2uxMTM3BBsqAnjMnuOv2CvZa7Is9iNJqwS+jPw44M9gN2k5KkHTZVxli6hLH
0tGFcDWrCwpub3bR57oQMIijDJVRxz4ZsoZ4ujjpwbdA6V6rqoErNsJjWvNnXUAJ56oBAzfp7lGM
fANAWPDVzLxU4ofvS6FcmswWGLEc5PooRVBq2jCerRA9qzXVRyFLyj3fMH+xzZhTxpzAn1OAUn25
MCpq/tzKVcLngZY3uAYaCVrLzCVbBQYlRE2NdvvACgF7yRZDb4rsZKf/Jvya+OjL2yK4XCO6h7vQ
q5XcBExE6I5cnXIK8BFHl7XHlQ+pcXF3AOSmQXIBJwxbYlnwJMM98n8359ZZoJAzP3nKq/AZypYb
hDkAGoMwLeJuMOJlBL+jNXpB/uG1C05fiKjhQsIJdjucGZcqStRMcDv0+3RB8GkGazXVMxwVg8cZ
xcLuxR0IQf18mRvoBGps8/gvbFSfAZubtV1yjtCtm0vZK1NkLcQAQHnPHgJo7mfUrg3dqQteJC5S
iDijFxCu2ELH3JCHSmgEf1GI30uGfaztEAos5Yam7Ti/t/FVb+HETqvoCYkBrxhKgMcRfBf+ZHt1
4KLU/X6Lf1NLYB2nYP5ztoNpuuxuMJevgtLZiU2dNJa8hmHK+3ip0iHyObRLkSsBmpArf176xsyC
j//qPSrfYAdS9jBjSP5pT9Atc60kbPme+i2ojUrn5LWfN88NcURcX0n7pA10XxPW8Ma+8qJMHfqJ
RD4BZJCU6nMvjA/oC7GaUYZmxmy8OZPYee1d8dt8CbUMnaf0BhHCjmoDefYAWHXgFt20mZbUj76c
m3E0xIHg3H/AIfWR22wQFX8Xpy7bhueM9+IWBWK+XhirrWRHTzZTEcm3RGSIDsDf1UkJ3mimmD8o
cfqz4fFSNFUYA4ShzgGc3Dq8pYh5lXEbYQ8AHpuypxrn+K0wlkDDPZJfGGfcAgTcDjox9MXApmnb
p4syi6uT8lVtzRHm1ZgwlJsLOqnUSjRB07iY35WsyC76zGgfjfjI0PLjs+2gs3xogx5XX5FLW0ee
jQBp8IEG50fwAL63NeUhQNnRanQYIj6RyMz9067g1q6SaNt2ZnohCN2tKCj9/Ed/74pUx2OMJBfH
OxqwC9yXklgTyP3WtHTTONkfyxP2aO1MTTWi/HaqTPa7zCjMpluMaIgiyRUIYNZ8oang7e8Wqfug
FtgcyjclM4AfLmkAnpPon4Zg4S/zA+9jeXJj7SAHurKhNeSThLwsyX5LqyraAHdZcr9C2/Jjypo1
wjG6V8qOn0UjwySwUIcRFs/RseDT01Af0E1s8zRK2HfPljKYkde9iLKnwCEXjea68XpirnkVoE5j
Hiwcplt2zDIA/qqFwsxFRrWMrb+In9cIW9ss8fPn51U8fRAiNliWdDoGKCCBhixErJJxcgn4C7wn
ngUn4TiAqCj089swA23YKvu+/dMXyDd+5B4ogWfkDhLMhSxc7fZNqTzJPvzLN81iXdVnAb5ngxta
JNB3/WKwFh1S0RRrLuDwLcTe5/LDjfXIgKpGjkpMJkTMPY06HcFf1UWhwm/2WvHu1ERddTMUuOvM
M1idr8/7CJmXetnQeBF6LegvPwcJ00wwO0Zil6cD3ZW/SvKvU2yWcPHo+yP2S3Q3MaF/51GH6Vii
7Cy3QhYZIJP86aFc1G4JchJi1G6jm0Hi4yaCSvFAF3WsortYb3jVHJleXDK5MiGxeZnPrwc34fb5
O97ZkErhTr87wXZQVHz0FASquHPcwJC0TsMrwcQXlAiw72G4BlgBz7eyCfo2mKFz3vmjOycLryBY
yUzuj4RnjL1KG2+gWSLaZUrn+PhI3Sl35IvQa9zUxkLEqT8H137c6N1Ku1QSSXCYGvg7qip4ys8a
khfyfQckDEmtYXS+46CwnghUICXicZK3ILHT7s+i7K97LtIf7SYTCUtdfu1o0NTLN4O8yi/NJ2Dh
tpytH4kp2tlZ6e+8A7T8NHDimPAOJ/GlIQImLauCy7OxueTdSkq1jnMqwhQv+ImhnIYysRakX557
I6s8i8cRIZ+oDssTSADYQGgBx04GfdpaicxJw4SoSYKCJtTtxM1tRegicncUq0sbBjzQFU2qZ/U8
ntXJb/UzCXJnir1h/czl/fyJUnG+qHhttvqxrFccKQCeOk5J2xrq4AnyLV3DazWmXesQHSAvMlhx
mBdD2UCRxjoGktHegzUcl/MrDnRWKQplR1lRVwWZ7ppmjLsByBeF4tES5cQDz6W2SbEebjLVkabU
3jUOPWE6h8OyW/1uuuxKgWg/9BKf7jh49GpxmDZdsA725fgMNP/zaV5j9CU8llJbqrmln3xD73uP
hm7TpiN1NDGXbomVVOguTvzXh7+nRPikEt3Vb4E3LRwgXpaUZZ5nMTEGaPgGpD0JHMFXRQ8VNYJv
n/wP5ifW9L+rpe+iMcVoqxPIkM2jMoztggFjEANuxEYksRLgaWpdVBbgF9ujWQ0yGDKgqGDhR7b4
as/SvEX1uf1F7VsjNXscmMaiea44JfGHQ17Y6I9AZv2d4nVJeadz9+KWAeNvHXuWzDjcowqL6KkC
VTcU3mt875PuMkOp3/qhtbI56dcgXzWg9yOnOkohjGDzdHNEr5Ri79ClZoYyhfX/mJ2hyZ3hJ8nB
YtwWusR96IGyAfdzRMvtwzJbDQM4Op0C3hkfRnFF6P+s7vFiWGv4HOqzSUQ9dWh6HhA5JSOci8MD
iJPU2j72FebFcMktpjDykmaeVCyjYHGi+NYRtYSnPOng2Dbkzuzkf/t+cnOrcYKhoKoaZtLc++aA
fuePvpgEAkg0csNBHGYcY8+kByN/YbCATJGeQZsuoRNja1IwsWcMbyVZl3ZmCzXvgQ6jPwmLTTo6
2fq8c4qEGudj2kVxFRXqKxEwATp+sSVLHwZQ3JNTwy8dJMd4eQquvnu9fuJWufYBeEEwWq3rrgNu
Kp9uF+tZIpOK52nj8FBT0TavYkyOZqIaW0QABgnuHDNosC3BzyHoRkQL7m4BcEePBCUgb3rDb1dh
pj+PTiQFy+6zzBpGynt8iJltIaPhUmSeBM7mFcFrcS4Htfb43Hs9bdkN9Bwu6C+/ql5+yMTg6qRd
F2XkpAgwz2YhAA3dziq8MqdBUlc12k3LyeLl6VB1Je2wXZg6KWkUwbyrfHNPQc+ThYzccBzAEkSP
PBlEWGmLrC50qumQ8Ex0epDEWE+plif7i8CmZpe8usmT5iWCjscRvXDXaMXK2MqWRVFkMxIVcSKK
duYPGT/zeqdBiBq+FVSFcZIGl2VGBQQIRvm833aU9/3aeWjQ4YuB1KvY8Lhyqmc2AT21Bi6CTzvD
ezavYmNYwoTD7ydMHRw5fa84loRmugKmD72l2PwXiWxPiwYfLKKD4H74qJ0/QNU/mMbW6fq92oFi
jb4Z01ccS4+yv5doQm1Lh0mlrPSpGiJGxx/GsQxFJj8dFyGckkkPhB2FlHf2TNXeCJJWzp2vZSFn
MANBrFx/5NrrV+7vTyZ2YGjH5KMj6FDNbcayBRkX20nR4eGD+74On83AsIvw70a5i1fxBBF6sZ8x
rayJ/IyJIdsB54CzqsnZDMf6/ZufTC6NPnPB9f1fRK1wzlBaasIaRrCgPLdoCKBpIAa7O9BUI6hR
mC5YMRmGeV1kQO6sh9Ojv3Ro0RsnvfpTYhxAe7VG0XMMdxch2+G0oL1psj2/0Nv//wEt+mrsIGst
uWP2fKqMbfoEhSCpOXaAGGbqwNUxKG7kiglzD4dVWN5YEqABdIL7RCnVjNvrzG2A5ibhzbvHyxEk
7kVP/ZtaHWIW/MMMLcP+ycpIxmEiDBNwVyiD13BxyEjlkXL8fKHBbBbxDcIBDgeUFPTbzqpuMqx8
+Gp53tJdftd1DB3BPgN/Z8/0SiwVOlhUe35alWorlEi5NknqSnRDgdL6/UOMNDXdqaZHABs8Oo/Q
GGjdnOoDGjQ8pC81E+y/nDSlKpYx6OdYFxYgia9uIjPGO3URt0SQ2PdIJo0weGyVGPSN3b2X9JtC
rXyUe/S+Z5ZgwosYE0qwL6FbKxolK9k93s9Lzs5CT1iJGuWqjuAV9l0sv8vMbH6C+bUdlJEGPgZ3
asLL9yG3+Mi280HiVHQeYXcefEHSb32nRoSpNYkafQkJLSiVCR8djpflL6djjjdyR1rUj8Y0pZd0
dL6Xi4lwnutajQsAtphKYbXw1kC4esVwisIwYwVYmOp5oNKJP+NXmwMzZ5AAiI7CSD7DTk+MFJDr
FEvbHkxwGH5gZIqesbW135luph5hgo3XFWhAz+nI6nE8ZDMc6i1fZEurti1J+5ovcvj/wRflgaGo
gkbgrtZF7on14SolXxCfhUWTYy2X8oIsOUqlipv1kq+ylWDiJJq9WfY0ltsnX60vNA3NkIprQ1ai
0vm8lYaviVDkegjbcD+xGiioKxVbWYFF5mjXy2tpW/ePkymcyMKthJuaMLBEwffdFtzP2uD3KhoE
NmlcCDDduV4ZV6CJNu7lCluJ9i0Misqdax5n0F0hY6OC+au7crR1QZmlHwjKDrFKr1BP6IFXQ8aX
/GXLWnXAIsipVpZd5HEf+KZlwPKMyKI5IJoCKDdw3iGg7CNxZMZMNbj1OICZ4mbnU54VvMtgzlnr
ERjsLE+coUIXBOj1yv06iJLCqyT07oZ9xyXzUfp24T+x8GFyVjm1vxmbh+gKdLN061OfU6LWfJfc
FA35hzsz9KXOrlurbVj3Pf11/s1xXVnLX9MgeasHU+bHzkjKvGfw/KWo0/skhyLoNdjGugbIDliU
XptNfDqyq6VzhJJjwCP5KESrzWN0dVVCGE+UlZ8KXSMLpg44lKqBSiKMdTw64SSpH2CeUUczElIQ
ejtjzoCVmgku0dqOF9u0F3U15GGquoMqA/+ntUiIYU4mgdz8G9Y3A10QZRYlMLQg63CB0m9k+MY8
NaEIz8SSkIaH4S10egqFWirAwZIPZvEpzMXdgWfUfq8Trn9eS9OTOb9rgVSfjYL9LrK7Y1v8ZAQ/
SDF79IEFEef4bHTJ4PLrkz/Cj4HjCT7KIqqw4dTHDHPsfiho2oUwp18V6kX6VhIDezhDSFecHO/q
jIbtGNN7psoeRBV0iRJTVYlO8tcHSUpNvwpzizJu7PWnf9V3pGYKlWNxyhM/ALlRcvVkZ7YFFe6+
LhsS0v7n6NuMmrMoN1Ew311jkpB8YivteXRr0K4spBvaTJJWVePL8d9nKEcB+yJ5c/VnrJ/Ck311
8oXrLJhgpGoRNlG9PjpPYwyOBUiuU4yfKjoB/5ijqcahS29WaOj/6oskNWVGG5593RHcWx0WHJCf
5Nl6rtt/FN0JvzwRn+LA7TyaSApWfjWNHvl+CK3DCMealOQg4aP9e8CEANdNpv5uNna73XZkF6o3
9EcIQC8YzsGEIOFM8MWy6lSCYcRbx5MfEAqSM5lzWKyvkEQNRjGHM6AdE+oi3t7J0cSTmND4zA1f
u32vMFuh8+iFoj+QwDuINcddnC/VKfzTCcfbrJSf+fP3gxeKtFbzTjoXFAU3AHoifBpvAaBimPIx
eExDPIzaoJzcK9A210O52RQ4ZTw9jLs7Y3AFWTV3l12Uu3Mu+lH9JbpmSY9qzsDeRljRUJythSvp
9cQaAhwfKjYiHxrLkfRXppuuX8G4DxLAWWjZFeGiH73VdXeALu196ZeHukCIPhFxJUdGFZRjUtDQ
knxQgl39nTfuaVjWlFHpJjWjw92YsWz3iTtDYnBpGGK7n0OUMTUgrudUF/QMQQnwG/wXKAPsOh64
U6E+2z1/F7OoaA0OW295G9m7HQ2kBmRSbD6qPT++5T9CsTHMNNK1ehzpTJiAMUI44Fj/yyZkzgOZ
LJEyzHwJNCEBISottm/qQCsTh8fjPzW5YEy8Yl3ghUObJG64iW51q3tTWWU7mq8es3RgtnuYenNv
X/CNg86y3dlSe2mO+oPTztTH+AGxssDXGms3smhuP19A1XgJ8lsT1f4jl7P4eFkzuxb8eRkULY1u
zcBrDGRuteiR/6ArRgnE4AU9vdNGkA1C7m87WY9UVlYvpevDJwJt0ZHZnQzf3GpOmC894+5uDLpi
+nO8s6dCQeAjcJZoFHYOQTaNW/GhEaM//CjtzWGK3O8QS1S9bvKc/a3k8Nwi6MallGsSEHTTTY2U
hvXh/2noXN+AQdM7xhc2UnD2beBlq/VFHEUDt+XPi3uyRDue3iO+hf1/xzCW+1Ykf/u24ruQwMp3
EMqGZYeHY1poqbblVGyawA3jIpMRVxnGeBtQwAeHxiYpNSPH1g3mXJ/RYpDuWS0j77RPPsrcnA+X
cjKO8jPVTeWBJmBzK+eazHesG0uvBe78/nSO0mBBi5uON0WW9RgnMLxuqWNFj5Kif541ZwUANSNV
ALZiTf3QpVZJXtaff01wcPCBokZxmlIZCCHB/uFO2Cy2e5DTUHJLINxEYFsDniEjlZESWRUycANA
cekY8C+6GZS1MSDX9d92og0BwAUI1/eWB6t8MvSAeWfIdbE1p5ujmVGS2O67dczBPnZ1WpomDMAz
Egcz+OirjuVpLxFACE6HEJjruJ26FguInkxSItHb8yWCEALzPDJhXrCu0wK++w5Zl7xypfHp8sf/
yWuWopUi75yND1UyXfPq9b0S+/W88oZa4y29XgijWCviQmjH1MPAiTB2d03YFG2UUYkvFSWsM3iM
QeRRogYZ/h0OSmobfSgYqRIBG6cwXZjrRdDm4b/VmrDjUw9PU3nHtwXuZ4qi2jz26emNXCOgSmcB
Bz/lrcz+fq16sDFnTgIeIMkEQEXBbPhLggz+KB7TCdIcgfYa669EvyDviPh37kfNT6OB1fo8qj4p
O6aJEA58RnqXlLJuIXrEEUqZHJUdNCOD5n6KNjnbHaW6s2HfcLWSzB2tD8K6UDM7ilp8pj0656yr
WkXc0mlYCSv/72U/UTms7wSK7pAna9mvW0OdFYaLL4yA9p/7OepJ/2f1FtqMLvXIRa+3u2jm2+0O
TvQwThRbEaN6+8f5NpwMGcrbwULWWEntRypep/NQmBRHTTGlTzBNyEk2osL4Sxh4WzjPOAa8fkMd
tkufUOuqA2wV/nhod3D7f5/1t+3cb9GepjNk8681YkmFV5iGYmC96OUZ+7mU9CftNgbfqAXzLmVV
b1nYGMLKkwthlKGABsi+O2LlG/2HhMKLp/Ye4PzoBI2jnepfMgtpI8uwLKv6sO1wWNSPuzv4wrdb
S+WyYkBAJZrbnsZvtR1Ax0XpCYjTdjEW5DRpvcmREpsdEIxwEGjRMtzf2FpWCIzaO9UxgYrX1pOx
LWlr+JKLoohzSBejKMHhmrCwYQ9NFHSkUmBLHPw6uE6WglX5YOtUSpqZlEkQQ5Bm15eILt4TvRdS
M6JgNZzu1lMzc2Hc0TEqx+1lwqq4sqx6jcsymZOkhpDXavRueC39TQB7ukcUboVMARrHSctoZUGL
y6mtIbALqnm9J5Mih94ooN5vHfrKNVhx6g5Y9dgk0HlArnNfC56lac0BHgVwC5AMFp686mxE8xh7
4FrLhMpRaSaOzPk7EuaJMfAGfWNL9xbd/5tVwA9n0IKzGSusVm6Eom3ZhT7/Ktw+TH28PQWFchvT
4eLXdKEWGOeETrU2D0iaw8BnJEAWMOq8hn2ALi7TMz53vzrGhGE+Psl4L8Db/S8LZM5h9mtlAUbK
BpfnYWG5l8ELvwQye9XD87xehDvdS8n/7ffuAv6Ks6RVaAAfNkLEyfCkPODzgwZP9mHEpcSAkQBe
3V0Ud/kw1fAgOYX926i/0qIuaIrRI773hPKo9Er1+FDIg3G6BdbLT2J/qq1nrs5q/t1gEatI+If1
ROKDk/BySbL51I+Jf545A6tkYFQdaqdHlo9yf/7b7DQya1A+zIWGJgMD/xzcTCRpKgwJcPcmwCI/
e3x9dvtf/j6yWs6FjV+Mu+5Cr1tsMNGIydsvN+Gh1Ai/HmJoHyCEURsZ3NJEt3sS92ZjMl5zlbqH
hzFTvi+HErCSlv71cgHqe2kgjdmY7ue+kZvhrDzpuBv/9g44PY51Ih81GYW5FJmGYfp8CMDCn3ZA
rqLK//7NrhlCc5OC4mq9blu+VudfyoUfTxUysx8yomkxy+o45BoVdJ4YYqrwptoF68oOUjbIn5pa
6Fheta4Oy2kcMT2UIy/RI9hnOYW2PX9vgnqZykEs0/M88LErmEjovI5KDp3z/SCnbYnTAFBNMjh2
QdxULdVQOfXr7tZ86nWJxZywjUpaCxk/SA3YiPWNR4qonizjHH9WqMWeQ+ZYkFhsUk8mLUG6ig3o
dlBX33oNYcKAmDZfKmq6qORKCHfGYuO9+OsSOXcA58Cy6lYHCLj6rKJNi5w7+eqQcYm/YfaHvJGW
oAbhyYwWcmzRrILieBU64De1U3AnHdYVM0nDaPfm/HuZbDY53yLlerknXOq/E3ptfFdljxduK4R6
BMe4mk8Wr1K0+gAbxIjr1o8MaGsGmqVr+eHRNuT0qDffIb59QH09zorXryITmsvcimTOuLYelELy
StSwPSXJI00tkkbspqGZ724ErRlujrGFIqH0f2vuawHkyzWzhNE7Qc0pG3Xl2FxbCtMbbE4w/BMK
pn9sMRqYO/Qle+E2uaVQiB3PVGCcqPtbHc2j+qDEwTlcCqcO5FGTWL0zvUoduE7fQiAbWj8RJ29T
SSj6Fb8kKFWk38jlP+MS9/m/4ia1H56SuwQII4AN0053nIICmz7Z7rKQCq3OT/G4pi9qfBXnV36p
zjj9WT3vkpqbRn2zTUTv8tNMdjg5zEzZ+kADOItNbU6qYi+RgLeUSC5VslSTPLCAp7+bw0EsjjKv
halw3vW1TKx5BCffiN+2z4oDA2dMMSEk3itwuBkFzmU6h8k0p/k2F7LCckU3xetdkXKexcsRuQ8i
BTXMShQnrF4DYSpUCZ2F+H4cWUeqVw3198a12TazNnlN1+O+cRTicFS0/tH38JEmcJTBq1Cnx38P
SIjdEaI6CuHHnP76p9CfWiY3yY5Tqme5RkEih3iE5stcLO7LnitbLF6Jqi0fjS3KxAvf96Fus+b+
mhKHFEiZ1PUtnIF+vgXKwTX4yIG+J+63axq+aibu1XKzXl2ULXh+oNWiVB9flz6byTl8MHItKb2j
IH3cHrr/L2l22/KExrgqPQC3Um/0dKxWUXfxpjrFIx3lmaTy9Vw0/qsoFAlYXdfwL6Vn5BsJguSq
SX/wc7lmX+ZZYSqFES0+WfgZQqsIvAfnmdfTviPJa18RBKf9adVoxGewit5Sd4IYWeocPN16qyZp
ZafebZ2VXlzuN4UGmQeh7/ncJU54gKlmw+IUep0irqlubC2LfjYwf7dz2+h8+oVs+DwZMQ3v2VyD
cAaCMRMfZguXtD3+VFoFU1Ulxx88PU+96jGPm1ofDTHqRGCQE57Zv8BvFQkX0HIb4Kxgo7qWSkop
V3rYtxlnfuzvkIUYlvpl5a2577nlty2Dt4+hQ/j2Ui/p6snCUDFdDCvXd1Jpok3kQE+kmfArQDue
eFDIWaBCHlD/qDk62YSei0ZPucr2c81K8u4flbqAsBf98RNjhMxBALi2pbRuHK9/3zNO8ByN/uZz
rGewp96fi4CjDIZu1ztCDUPXBD4cEjoqmLHrVpUEbeSZPytv8w59WjuGtIzMZwsYyhJJa68hLr/T
aFnaVLCN7tAnda0+aB2Gc3LP37+J9R5HI/mADSKo3qtUHsfiNvFhsnZT7xbcWcHSfg8En45HJE/N
yztnLUJV34pB8ESNaODchaSxW0MyNUNXW37TD1bgko+SrZAZPk760m17ShUWqlsI4EBVB7ADmhks
2GUCbfy3MYoTmol7k56ll/xibF8diRz/iDiXKZfDtQ+KGW1HQEsG1tMW+awm/gK27EN0ljI6LoP5
g4GUt/6l6Oo2mXWLGh3hobKMo6tJGFlEUMSWCKuWgmOfqkMnwom6oJtsTAvEJfVhF3GAeUdjlZkP
CreYrP7VqLrOD5ZcIHVmrzbX73NF3AfH8y5UlnUn9+142KdG73sT3LoUiXxHZqf8GDhFhlxvaGQg
s9j0IgI4TZAyqn7RHddNAkMB78HC+X4flyDqiRZO38XX7d9L27KcIYFury+OUuICcTP43VoEwEPB
YkHfBFrr7iHWehRLkw/cWyB4aaRc7tBaX/3U06jnCpOj2QW7KrZyOKkK5Cz2TVAqSUL3E93+0+5w
wjitttZSHuanVPw1CBOO4hz599t0im1Cu6PEPi4wkdg5xmONjp2uCQrYss7vvDG9hnjow90SD76A
LqCd1ggQheMuidLHtLn/sG12GQ9+4jkOxLKxsXjf6QrNULO5rS0AxwyzYGmnlv/4Czg/XHzry0wK
/BgacWOU+7CsP2+0gYiffd/UBmoRE7hWsETtvhtBQYFoaCB93YYj4uBF4DsinXgUzlL0cPp9wGzV
Bnca3tbXuI9RcvdvP0biRoxoxym66AlMejypgmldxWBe2pBcTQqe9Gx6Uyi9cb38pNBsEYNix5Ly
a6BRtyTROOrXmzRDvdloM4Saya7vgPblHAGK5NV2UGr7n/Qxpli1JwFpGnYbNpd2lLJKyb6HZSeF
t1ve/jMxmGfshUKZmJJnptB+rAYyIfXjEd+gk7uLfEeU2W3kbED13CTyCdxMmlKAXuiJAI860xHU
ysqmJkMtxP728maSIKfCtyqxt7GoB2+zmkRifwb2AbHoy0ITmXEuwr3dUkWbqp3FsAQrN4KiEC9g
GbDrlhuedlsiktKTy9EuAzqdONay5Wv1cHmMhYpQCdjBTrxZ6K9Cz5D4KBHkg2KPDcm7B6rV7N8T
VWnXWxQ/+pafDL1Lek0hEmVUqktgxhkAzSQEBojtyVmgLU/xkzFzFJjFlwKTQUc2iW3vEQGg6na0
6edpKzX+mFPO8cwA/KCKDpk/CWvXeXCwj8npQdvZ03CKb3l2wJUEt+6HXYTZqKiHO8FeyzXSlZDg
m+Rd1zNvKWGr1H83r2192aaOYXC6t2Iv1Bo16l3IdAFhFM6lqJa8GmreTI5xZdwyvnKXzwu0Zzj3
7GN39MI65C4+PSDMM9/0WHVK5mOZ0FiyfwuJkX6h3BYD4ol8O6i2w98TjycKZry200s1GY9DsiKF
ytCFOkM+QTJrnfklZewNHP+DDwk4G0FsqnSGLsvnpO8PGO7PnBeP5BvWvFrGeS6esIEr2hcYbKvV
BzB5SpfeCC0ubdLo8HKsz+vIuQNJ836rrPViT7+Y7hnyFy5XGFQGNKhffcl7YCulXVg59mOzUtmw
L+FbQrpJLyn1QC834Ha2Hu6lGyGA56v/GWbnPAPXllBWbZ5+7IggiKaA3MCCkaUYpBPor+/ZZ1J7
3P0BDNruD51JQlC2HxDAPUENdkjaORJME390Jkv0uPf3KLmR02BruqgCbk9uqXdNmqj9/7gn1K/6
H7VvkZZ0xdhLVTCmIUXk0I1+i7iJkm6dyekqWtCnJ0v3goEECWtn2lVpj9JY229nEIAAQsVZypeD
ahfimpfk7GeQXogBa/1ftzMAon6lSrMItGWI4pTZ+xgS6fazuobTaYNkPjQzBiHIrtU6O1EyrTAf
5q8uFT/i+UkOJw6cT7VSxoKehwYwDgpokae8BAPJtRx/MM3q6GO/RvO7k/mlGlSX5oa6T8ybOjxR
Td0q4we78DZadgUZFkDTicdQP5pdHu38QQZspnvAcBdpj+KeuhaLLRnP3oxgv1u5L2CTu/cx/jI7
9VZtqokGD105jzjHs8ecNUMFKa6lZdKfpewJD7ct6VYLHWb0QuxIQVocZX71FjZFyy0yB+kdEvoO
v4magetcDYBvecWrjQFitVsoDv7NHQ4PimKrBAK4vsj3ag3EceTOxdF4LdSrw9cWj5fbQgFKH8JU
3Xx9OAQuYCU1NajP1E+yACiYg5xZgRIuvLttYTMRkP3Od8Wq8IxnT4W75QG9ndsITLt6qTnbS7TZ
P2Yk43iWm7a7FO/mLjmnkcqjTaVY1DFCvt6dVGUN6PqMudqg2mtTPEW/GLO4Cdp4+xed+HtIIlZ3
aCliOidszn2ATabOhm6+b0bTaKHHcQb7lZiKT0dF+Gv4Aw4SVXuHZ5IUnVuqktfLuf7GAXNGAr4i
2SRG5qOii9+P1x2NJ9XdoeeX94DJkEVPZbmRxe1WYeuaZUzYPnPABg6kwcxyUU3rnKwBeil/ihVK
boJ02bpAZCgggLM49E7m1vNbeNSikJGyqUwE58nQ1fVCo8clRuHyKcUvfUCSa3KGOfvW6jEPQKvT
QP7N/cqK3TL8vF1OEU3RA7VWiB7R6Ib+8rSdHkvfHYXUG9otOXqxPtUTaPPftX0HEaf95lbD0920
W9T5y69HWF+W4AVKQldQvkuQN9fVCduFzJqCsanvU7n0M15YLCKEoLJ8brNW9yDAbCstZyPxU5ph
E1dki5z1VlG4MhFu9ZYHP1qn2x2qpvUcKcCKUchEpRIWlgK4MYFlwgHRmGgUMwLeO+KBbkZDOebz
yeEAkHu66p5lBXH9eyR7mD8cIJWrTsr1q5YPcOJJLTkozrYUmGEgD8vU8MtzbuC1WMVemR4dqiTK
sviLGVjcSl5PU1TtmGF5DxSz12PhAYvh511UO59wazyRpmDKzxLT80bAuIxc/LOT32RoBWMdJ0Q+
xZrG4v55o+Z/p1psGD6pE14NwnxL1R2NJzReRV5BvzAHvtxMyRb93QGBrgm1028ZJh1UAGoD+QRz
zczrhuiA18J9PeTHJtIPryMFpa5cnTyr0pSxDmA3Oxd3mcUVgJPrD3lqX0GwEUeAKki1cfjoRtAX
Xb8zgRLJd1x1ZT3MFkQuQg382t/GCWkfjdYjX5faHLYpGsXcKf08k4Nq0T2f9wDeWJ6i35XTkKAL
51ksQwN6m1/pSIhZt6kOAl8eNTvvm+ZDEZEoHCZZbHGd4uWZglBKeDyUtDqbTb63RpVPnUJ+BbYz
scGeh/fy6fuy+GH+DVL4NZeqVTGMDQL4JgCxI4utuqhL0vob1nxR6M07nwp3OU5Le6Fnw26KVlJb
l6YMZN0LxuonEKRijpZWNJ1q7hQy/CE3EVuoQw6MiMOo7jGMcDd2Wh6YbUPr7rjOAnMt23DcQcag
65aamisMyIgn/fz5KyFoBXndTSrPen/s+QzFf8Ob/rQ7f2GdU/t2+ptxl0zda2Gy7+L7swhOGDE4
GSVHo7MhlP8cp4PqP/DktAPLEdAWOjBnbRYv+bujxS79FZu+L5wZ//LI1Mk6lNQfa8PBQMU5LT9n
PU8mTnSkomz6f3R9us17deUkDXIAlPAuIIu3CtIZNW29SRYt71gJ/0nh3ZF6SOxx7q+dbRRMomZ0
T0fLCwEbLQ03UWbr5VfSeBMa/mz+ao3fHyY2blB2OYQJUNWpY3+mOA47YVQxBfZkfMcJkqbeds8n
fAwH8YYBxrh+lY6oZc8NRhD7nPEjZDCaH2Dc4shkEuBDy5jNfhttG2KL0nkfS1Psk8ru3plgnOrC
3MqQTKrnzBrFDYCFZnK3AGYs0bpgsQkqb0EgYI+LK1OjQgCoFphtj4WyWZPFQkdPtu/8myYyYtsQ
tMLUHBaqYl2wZF02g2+KRhQEP0wK/+qBH/T7IIjtJvEPnDzULxzTnLIUUwVPT+cy4CD4CITkPUf1
vfRcP0Obl0s/9mPsoI802wqDVDy/kJrshPswc9pk/8WjIqdeN17IpxggvKzwD3+4jma5XGCr2Bsq
iqVNyMHmr44RzntEPIruE8tVcH631hOYaGtLRSzkJh9rW6epW4P6b/J5uun8Vm5+V2ZPytekrmuP
biILO6MgrDdGOR0TfLRU+3V9cBPsOBXa8M0qZC9o+Kc7+4UD4zX4rkYC9ewcHNyBIgZVf2IOVRjK
w23EWZnDqveG/2Ejyb97YCR4cZ9++sYUacqLDJhgbwnbaSxex2PK9mjhbvKqmDjSu6pnDrbUP8YT
9NUbwEON3XJe6Gz+bjdM6Lxk+ANde+LOKJclzjV07/pj8MgQ44bYnSm5BaTfNb4z+6/JDQ9UfxoA
pD5eysdRwlFzLEqFrJOq5YGfzMMbZy4Zi326WitYLfznn2DYU+kLbMaGIVCDKgzpYNo0aaXLW6Zc
ca28FdcuytkafohD6Kw/2loJFbMtmcIpatulFE2eRsBHhj7QjG85KTpKl2gADxxZIHLl2Lyh1DEn
iF4D98YsyMMfQaNZ3xPlTeMqL/OR5ZQ9lw5xBP9y16eNey110JC+wxHbr4s3Gt9iRYXJKmnJPeP+
lYQDoLK+vL22jmM0rqrDVVMNZLlS6IN4Xrmsm414fa151j5zcN08h/brkFkFNFQ2evJ80Uywj7u5
NK03cFxCgzTXFXBzd//ga0krHxarSi7w4LwiHJsmzPoJQVjXFRIlM8G7e93c4D+7SE+DzDxaQRxr
Wb2Ta1H/QvikPgxrQDH5TkNfKcJor9s33S7UgT564FSFq7lFUV2dHGjyCYomHTxOLC16JV8yjm87
TBMNwNHB3mY+kh4cZcdqaQ9+3C3VbepYDR9GKFOfxx/+ixjHY2GM8uARl1JkgV2pdLt+emT/6DCo
GFNTAUToB6hyaXSfAxggHZrY+B6uBtbLm/ZnYF+5HiIX0P3NIPNGEQkopNrwQPysbdMfFXYNUMCh
xtQUrSFlk8Hbuu8ilyPA/atwlvP7SFdwQdDyvjVlLImZrnBcowYZydjtEciKWGDlozCFbOhd4ckP
LvtIBO9f3adqtPUjQh0fZl3Ef/6x+FOpiT+OChW6Rqyk5YJEUAK/asbhxPaxe/upaoroNyV+wLOF
+0we8Et8ojups4yP7KwUwKW8CMGotjEuH3aT4dWjqlKdDkxzlPN9ZKBWGAG70oNlCefuhdcQSVIn
YWkW3QhshI3Tzl6tmw0/bwscjQojzXRyzRDBdU6HDEZjHp2Rlo0o1MAtekosYssS8bW8mjxs1d7G
ZRnKY91yinr966PuY2yqgefqPOl6+G9UFlE1waQH2nJdVPIHUSwZ8LaLYLyKlKZijNH31cfiY1dW
euGmdMzlWBTR+qWtnn0ocojat98b1rxMqSB3Ui3tV1tl6zYSM8xYIfQYrAE+rIQQMDdDoI0cvVkL
6eLaFFJ+dPt0alCvwHyMDhwGVzLM6Z0lXkox14QE5WnGcktJMxIF3QoNrdnnGD/io8/95tjefKfu
lzzN7sU6ZtXLR0hd4LHvzzZ7VW2LeVPsL6t381yX8Q9uDLzsj/ER4lFVNjV0uVlJK7+jHtDGt8LN
OL9MV6KuYLME7STA/7/Z70DwL9Fozh8KiDaaQ6PfZ2oTdzeZWOdgJcG3X+LNntg2a0bwy6Iq1uQN
PDKetsq6UIdJkJX478KWdUzH3tktdzyP4LH0qauR7Ef7KGaCjkFI/ncDcS7wWIM9OZ124p1mZX1O
uwqpuFLYUthmMnoZXS8jeV0M6bTsX9wDVcdUD7DtMVls2Al3VBIP+TCu4wqJAfiMsP68ZEy9UM3X
IkM9AWfcHPp/e4lWcZbuvF/xEHT0298UGGoH+wCnkn/23HVjx3F76IHzWyzGtaeQ0XPysBt0jTVD
9shrPA35+ub9zO/dCD2lkp5D54gCUgws9jLwsSIOsdFrEaqVzW9wnEQc/gzDVtwC81pAQbJdWu4+
8JrWy+vcZBhmzABUCE5Zoz7vW3D6YTJ92Lt2a4P90rdsaIOUv4LfXwfqplFfiBwNaGa9C6GRoP8c
7kDinxzFuk9VJhnCW4HRp0kkjdklNexAq+yBsg+t9o/Sbj/vEmYp+c4ecwV/kyH2CojeFSBLKTYk
auxws4eZ8kxv83XZ0oM6za8gxw0MEEV4wRJis8Bv2L/sL7t0tQE2KUsPiuUGoE0QUyTezSwNpTLr
iXZgoJ5JiYjkZ2NtwxNoacB/EGzWHpJ/9zn0Pgmi2DMin99o8P2IXiU3v1+tJOuTJjpqqOVnqsrk
gjhWtiK7o0tI1AE8wsHmFM7b3/4ku3YxjXhlapZC85XBJiNeb275Zo1QMr1dlxRnlgAubA/c2GBj
UzFNrbBIWnofU+uTw8LhCp35JaiMAcGAVF6DuZGT2x9kbVvPB4ZLYqTKVZlqewr3DZQ5H4gbnXEW
8gb4bFUQfGMw4u4fpOVKWMtAqg3VYJDh4kUYtgf8dasXak37lF79RlXVZSnEgeKvGe7NZx7MgWrL
DxfYbFBcjeMkFFCxl1ivmK+XVEoBDjb0a4mZEiLcj2zDJsnPcvsvqxHDAs1jOvW13T1Da5nFg322
JX4pEtC7PqIDUJHMuLyrtfM/hKT+HAKqHbo2x2Vu5gcWhNW4hArar2rYiCcPTkc3SzvhkyMfeXMQ
mM4biZ4nX/+GYPwQDYWUR4ro5uqpUn5pz6N6aU0SsHRc/eB+/K8EfwqJJmNQV2v2A7jvNxkm8Xrk
t5zY5gI+AmlbwH9zmYGs5ZmOnb3Y7CM2TUM5DDiElCEXGOW7sqTt45c43KLLMHIO0Re3sCONQfTy
25qkK7eR6KqdKGCg8Q13COhvJ3Sf4g1RRA7SY+wM9AzycduPcpIoLkOY51BzyPN3aYHiOfc3wg7j
2Zh/87/QMeHiX41HDzLj2rKGHdCHkWVKwczzUwDQUWw4hgwaUtXMF8UAVl4Y5QC0uvDPh4LnbENv
5qCOd1MV6BNdhcIhRK58dNQHiYtdduiLW3ETUBMtOe90ErGTOaGlJENvIo0gSm0/sfiurTM+VRPV
HNwpXhS080yFGAKS9YavMT/vqKypw5N3tRh6E/nJDygMap49e1EXiswjCrElsBPesrXgIHd7YYeh
XfuAGfBIMFvBIkGRhZguMYGNwZ6yOdX38Sr3I21vuNVgcgcbvyVeJR2qntsRRK/g2UGK3mRdTfwH
ldyNWxfDJUxwuwHcAaflXQkfNfjnMzH4phdXKJus8PvhshHjqX/1QMwElMlQjF+M+FgV4U9Mzo2z
Brp7QTL8Mdu7C13vvlOSGML93XvFq3BR9IivfTPUCULasF7yPZ+fNZ53b2CP/bf5BoNsMhvEC2sO
6/WvccCBO9miKva85I9GoYRSblNaidKeP/Ym/l6pgKyOl1w1QcZaH7QYUvmkpVoKnRR6ejkhMlK6
exMnLQLZBO7yYKcJRO6Pf7/C0f88mK3wH1DScRnVOg9/AtODVfD30L3phO0TUVcJInqmkYu5sWZV
XE9MH3BiJT/xvsBWpgDKpHGzhNKfYyOW0YB92D14mUWcNbG351bmhOINE+55USdHyvkkekCe1VI6
ydVR6XkSt9fQdmoOW33LoOhayyqqUA8+2VexPLcBw/l1pF4fs6nLfR8UiqCGc/lmxtSQJXfEPQzP
my8251qQno/fRvgTkz+XP2oUdwSRiSX0meCDv3sPUUNX54/bS/L2PFrwBhxs0W558rV7DnewKEAp
ARIwJhaB/Azzk8uA7YVxyGLMPW+oyNv5f2fgOtMe9dZlI9DCKMezk3BsDscvfcUBHzMFHgqM4wR0
UxSkpSXDMO+Kkw1nnsKJtzs3VO/khB0TNlstCWVAyLd71inK9tNojMl1MHHCphZhI+IeeBm26OrH
B3UA7PLLjeUJrSRB9jEqWxYDJVNJQR8CpQ9ncKJC9SZys1uQ7cQeXDoaLTGEwknrAWohToT8b1Wk
AeY0eGPRcEUYhN1Ji5xRtaqrjmPZtTfseiPiN5h5sUh+9l26BESVSOj+d8wBNVQo/8SvIK84cz+Y
JBM8nHH+6Q82RhtILHTD/TW/VfbktZze0hIBqmt5jzExk4UbsZSmPKzl4H01KKz6ZVnPk8lYmGhL
GWlQ/CqfX+ljnLCQ3Uo210JOTN0JI+aCjfmiASSCrC9tJRsMMeEWHYEYGNicyyyRoaN9AFosceyV
klILU4EzheHfBApGk2IINJzGCgoVMO06VDtIrDu3YyOap64WeC36CP73Klcv4sqFdvux3XCF3uRE
k9vybP8bgm8y6wAnsh3YBUCL2TKo/TBKX9urnkkMhtPEgXsnbHku5iulY3eNQTeT9qQhZr988IrI
GToFN+tL8Z5IIJBYptfHq8ifeE6M8Gz2ZVKNRa4S/GJS8AK+G4kkkGignZe+386bLHGBH8rLYOsT
aaMfcvTfcpAmebHSUZV0fJupwzqt5bMgpynqUkoeiNw5JWd59v2fEQ5uE7/fEW6LJrt+a+uZNX+b
ZafUqqORlJHkHCrEg7RmZXdrFjnOhWqrTrjU/f1tsXXKRbRi1HD7AQwygFrj83x04kFWHfgR6vzL
X7PIC0TW78gogoK68JPsYgg8LXUkaXMMqwV8/RIo0QW1VS8rick3y166Z7FI90M+qFCKpGpjwuvG
haQHgxkX5wBsn6FMYdV2YEIVRBHPGOwJb2beExVrfzF60GUz9lU9SswVYFrw4r3HtDkzTRUBR1Uv
snGN9/LQXrWLv3ujg+07I04aF3RvqeWuHEuok4sCLJq2R49JYsNeEDOXJhICFluEdao6ZL8ll+x3
O1Jz1dY5OlDA/TqVT+hmdYShUyzpvVOuQdW7VxAe59edzpI8WIYw0U+3AwX7SIIlRQoXST9QJeDS
KHSelxs2in9GBBNHIgtm1thUcAr0tIvU/AZoVF1mOpFV9mtg71nzfnwzz6bNQIg9A9SsLBbdgLhn
H4HT4IujzAz2lPXvj8U6t7xeNwVeZQgpIQsLYnY9xWeYBX1kKMy0k//kZ+mfn0sRsWSyLoT3W8uu
dKM/qrOOzF2f9TSR/mYtOxMmjsCTLYcnzkSwwWBBOnixOOmJ98w8DbR1Gw/f2ZexAIL7zL2E+6bJ
+Qy43DbeA3Qi9AC5Shm+IQt7TAkHxYtN2GIypMyE8oKv8KRQkW8o+SVbgiL+bo/pVibwsXLZ24S6
itVlN3TKvt0l93QbMIvhel0wvnTL81nnZUwjeYYJ525ctRh0XVLA/uECP47SLwMk7I6u23Ja/jZi
3Zkg17ygMz6fYvjk3aTL4qBLoiCO3jQl0CKuOcHGlyS+jLEvI3J61t6rTHUJKX27GlwV0EKLIuh6
YwGPLc3WfvlAqHvPXsoeNa97zc+JBawUKI0c8KyBJAMkUUzvdVrP5O56EBNlqtLoIUCP/EijvwN9
ihgdbLZVME6Y2CkVX6RGX0mL5a58tt9bT59We8VE/VXXO0oLcdudU/sWet0v9E+DFUPosDMbJDxB
zXmYBIiIb91M6UFm1wKu/pas1UYF+C2aII2bs0X9mtxeAltSRY9HdGzfcMItBeSWeuweeHzkVToA
khcYbs11w0SB0AwxUK8DE+iAZYBOLrRDELBF6Nw6W8Len9Dy9oSQDPX1/Bd6pBfcZkC53/9ZSHiH
wakLmAP+HNfRqfY0X2IflLLSsoEu311tADi3xUlNXsHC3HyyChNxanHGWM+5E4CYaJphkzF41CRa
3wMY7NwiQewvrTHQdyziZB2SXrjz6NmEDeofTU4O0zfoy0h1vL/CAYYuS9H2pp2KhOCCbACJYyga
kTxgDi1Kv1+STGB5R88gYgPaORo5RXTNUDuqEnR9++81CgwXdvXu3gy/02XE+HVDnM/PkKVIuPtJ
QkeoEiSm5R1+6dnpIP7kJTpUEQeH3Ec2LpoiG8hONiFvXXSZDdcUPhhubfh9AMsvSjRKQT7Vcpb7
35k/jiq55jvUAouzIBRpqkCysjyvvl0psGILSnNrI1u+hte/CYxhRmO4AihYj+US96KJtoPc327Y
PjPRGHdfT+OEeSoFQML65N/ZkWwqYH8v9ZgTi4t4o77/+3UPw4CzsZfrmO+2aH8IQDMWyp4ecwMT
njTy/bZKZ9n5PcaS+SU0mmPQ4VwAx4+ORYAXPla+0CKOdSxhxtq6eppD6EcSKfvmz4toc7BxLu2z
kNkyJl/lkZUiqSG28oZgbuAdtRYRMZelZ/2SRTHOM4RDbhbRARyq4+TsHxhZRzXKHG7GV5as1bk+
L6VuixCxwXtcQ+Hu1FOU9vYdMHTxpzu2+nNLbyqLxXRgewVjmJTwopUOovyErhbyXgZkxtG/g34l
+S5/FEJgwuhNW/57oTDqYfleU1GGWAVIxbVt4x2Ln9G2fQ55HEEKUZE83kKVU+MlFSkkGxjxb2fP
e1gqkRBPsN/OMXS6ukVvDwV3yp86l1IFyY55Y1BkzvUJ1GOBaqzdWrECpOuIIOoJrq2dNFpNl96P
k1wPvDulHMLNn4S4hJe3xLjWysUiaiQf6EO6KkCkHI3s14WcYiafg3nhOAJCni/NjY7slKuT2NgH
5L+1mxlJcFJAeQkYSjJEfcAFXn4+pfbUTTjT1UyxtqoxPCpsukfxE1+KuQ69F8ZH/8QbKj4IBOWJ
TL7VAgakd3KLbRGMv6T3ls8Quxg/ufIWXx9nBR/jcp/VIEiR1NkBxs+Sak0yvnLFVGyHPr/PqQ80
h/CTRro2jzfsUTRQHDHBDcD0XFfPa7gflbSkPz2hTxj06bADC6j16F2GrK9lVPc0aiZd4WGbjDg1
4db9WNFR8xLn2ddcbNkd7i6yuntH4O4PnMIWpGMbOL2mav1vJ/SOXrf1k5jSgDUysAi69JLQ5ZZv
foNlsFjBRfyij5BMEzaFUHXmISi21fycaBtxqx5pr34Wx4U2MCQU0pjOYGEW2mmwfO7eEhlNd6rJ
i94xwx5CSwGHYdeZE6QYbMs6ZyxPDgiSorkslirTj1ETMy9nqg8ym89u0p90GnaIsHLC8lJvN6YW
R7qWJza+QftTOyYzdnw+z4h1CXdAUsOBll3o8IKJLG77wUH9kyXrDLT6c3QpvZu898YnC03q76G3
F9pKMCm/8SzipA8etQZ5Z/GCxxMOwfufCjMkifFRKx/Pach+UircT/XqNvnLEEHLsOhwSZNevdgT
uqaV5HxAo3RZf8XCSrzyqa0QchbHo863zNG1Wk8ql8SPrTBqqvAjR4mcd8a4JeDtlJRS7HFjrIe1
5uogKuMyRxUQ0hTuvYYxvyQ9aOAtivDWh7sUUiPLNApYiDBogZlCrKs02K4uY7h/+wbCygULMol2
am7GFj+NWG4Zno0DFFMM4vX1XPAs+r7KY0AogG1taSuh4tIzEdAsKiEZeZk8X+Q5JgzNivhdZzOF
NiBVVhc6pqNUua660K7XIHZqT1lG6Hdog5B+ReDsHo4A/Ta8Cos7BUZrk/KblXazLPvUWmnlvRWd
5FGZeWeIqUeBI62O8g44rAhStpwJ7UhuFlQmJz1N00whHeYbFvqjetUn+u+KvLtszV20xOzmPpMd
ChKcuWXDE5vuSpj9uVs1KHbHMy1o3RQpl7GKnqMPwT5QPhptlcdJGJOEXl8+gwqCAmwj2euF6U3Z
x2l0DNXtTb00NgKFXrpFWuHL2G6pUuNdW6EO6c0lO9geCyxSnnSp6CCUpvhmkNq0y5ymg8dIgFjm
nG7ZI9VxLmWI98J3mCUDRUbNR1ZaN3LZZpXS+pLgPxsPtjoSER6ihY38kTHxWDcHx9rSVy3a5o4N
Ws+quogGzgnWHPXCFHxMnoyHSnXhQFLq5YTztkhjQ1pvPHi+9NklRvR24J9moQiOKcTWvUqD3kwl
3VEuEfM8PFSZoJKNG/6y8ySE+nNp2uagY3FDOut4VpjmnIByxo73/IdBVnmv2t1sXe+l6Rky1ykv
jtA7g98nCB//AZb6PifrhAxY8q/zZnrVrlgnBnCyWx1qVF8ASgCYBKTXJt+ntgFqI3fcuyn15Ivt
zfRe596z1o6hiK/0PGYW5PwDECQMpzXrWMzrNtWhuKxmAHT5hYQvw2b5Llw3iJwgeD0TK3h2RKPw
hwgvVzbRKP6ZulVEerkL3P6QPUwKoAbg5m6OZW6kbboLvd7XaRUoJqK68r2CHXktbozTYm6Bp1x8
K2vvLw4+feWOQceW23mO8UZSljtnt9If/vHw9mLHBcro/jdjf8iZFMAB9b94L4RnBiCNcIqap/EZ
Qiu5UXCs2RR/t6p0cRkyfVGeR7ANsRf/6B0moWNUmNItB2SWIceRe0AoTC4lxZKKEUkzD9g/gIWt
j0pdcPwL8NEofbc4ORO0uPKti2ZSsdq6qi56G8/bJZeNIfHYXKqtCu959m66E6ZUJ7Y3H4nv9y7A
BOu7Ly3CQ1fCHlcVXUse8CDrL+TxRNtHPf0ptT1sQxpPVyrMFSIK/RG68Tk3lVHw6KkcNxvQ0aJ/
nCXChya3ypD3hb8vMNj98JN5LMWHHXRCr3HEiE8i2HRosycAWKZx/eyGcd7eZsyB6ig0vpJWlGvO
61JgOBcVPhhc28iCG3t8YbbHxXkGSk+g/Fs1mha9/a7PHjp+SjF7F3MskFEXV5ELKljnnddJ4im0
DWLOfy4SyY1jN3cAa30xvR8YBZSTX3L08/gx8/70r7wt7E0dvrtyv2Wnl1Emc+lrBwaeyL3/kpy9
3bx++voVgZGRyXgp+uLICSZR+9RIz5ZhiAt18UpDvGqRwB38oCKcTWoP8V5Q3JsOWspU9dK6Xq7H
jY9VSX0ZN3IUoROt6XubL6L3dgpE2bVCJWgiWTazgLcct1aDZUHj4ILw9UhIPchzzHmMydivvdgh
luzdez8BB4rM06G6CcLlASeWyv7oW+4h4WwhOR41woEZeERkKprhC7I9haE+tLrk55s0HjFeh+Rd
2S967xGG35oAp1NieaQPtI2PkbxqSNhBSCR2cw0TXReSdGQLTk8zQho68d6LQkxwdHfmPqlpqVES
5rFA8TdNmXarZKwCEIHQ9NLzrVH9YRcL90NfjIMlk5QD/inQ4xBY4islaCavhd3FJylyi8p20y0G
zA1w5B9XUI6XpMXW0s+F+goJWVJZSe6TwEwUWMHVQFKfzEJijAIq6MDEjm/uhMd19Ws6oceAW9nZ
dAeoxsAtKMsKQHOEoeo9I2qF7+ikTiz09nVmjGT035v8HxBHGyhQdYg83vh0aK5BKElvxORNt6Cg
spK4QCNAZBKzur1IX5yU/Jz6Qjni3BME48y6PHTUJoDpmuzkLx9O/4MUcC0NcUJop0SHTcUCL/TC
c+K+Yces7yPJ22dlBTixEhIxaxEZ1LEa9+1UERzHqLYLDjnYaY3YwDjtMFY68fJYrbBe9OSCI42y
UkYIvmRZb3n592qDY7bU4w1GGcgjtqbWDKLLHymhrf9ZQpuMJmZcoqWWJPONEjyIUg/N/1TZ25Lk
W9KDJW1kR6QyJG7GyEUGmNITUDbKad6taLNIGcQxnIJopg3PUKsC1h5vDFnbsM5TL/uxgid1PbmL
hnWpJqJbtt4Y1Ww3eI8tOQIPhA0EygT3lGuExt0YPoBUKPjnx1u4jnZ/+zQeKt9HdkCb4h92XcQa
QcyoXL8iW/qYq0K5It4/IQjPh8gtZ3BxDinBsJM6CbpXnYxy+U5LW/r+xzenFHhSaH4QG4Js/Xww
0D/9RLSHPMOJdId5hv557wZemKLs60X4rRTEKiMU1X2NDTvI7Lk4E8ZdrP5GeeupmQAdqON9YQym
GX3ykHQ9etlcj9g50PTsI6wJSu4lzy0FdPitzccD2U9zxnbT4agYIEcshoGFurdoRiExprtUad8C
ITK9OEcshHe/0m5ab/LkiSST7BypjZuDgxPe/hO3pYf8ZuVONvR66lqOPBAqip9fiZ6ovoKOGq/Y
itMiLC1db8E04tHzlFKIiqo+A+YsuCdF+dOCINZcQFt4EMhQtPnHPeA9kESA4WksHDt0AKhsyCFK
8fcubjZu8TpqpvbsdW8FYZRMowafn8cmPewF7Jnsr3i6aWmRvQ9srKLVxHhEDvdT2iUvtpZjV7pU
Xfu4ShRIBoGnXOLsZxATEHr1Xk72QQrr7ogHc2G8JdSxQAQJJzTuxQ+44iklS1wJLeRAxWkuNvmM
sbXirXXzRKdv99nKIeV678h17XVXBtWLLx4k56bQ3odBX1aRVeJvkHf4LwhhkmcWXiKMgV7a9Dcz
13e+gqtkzAJc2frfnpvWWb0zars5UDxMEEQK9FVvm+RyfWaCrgy9W/PzRC4SVpXARKMCTjhkoftG
hqlFj0fom4jL/bXlow5xoyjD8tFm/5pBl3YUpOKX8DNoLu71DQH1SPyfs9Pl319J0FQiqR9LdUzp
niMP3y2R8Ni7s+V43KCrslX2fJ5ockxxOMIu8Q7ZnAwLgzb+yA4RhNr28FhHPuQwNXpotbrddlmz
ZC3wdsNbtPaHRZB07CjnhwcgVT4r58JyD0n9AmMID2c31Wg5feaeZeXy3kzwmQyNR5+0rOf39sV1
Y8SZ261Rz2KL7QP39gf8XW4mpUG+907nO69/RCPWqb2mox829CSdF0qfXdfNuFvzYLx3ZGMlD0I/
ObcVrGF2E+5RvwdCNdZ5GyXKnJpHSA2DC3iUqauhWeAtDXLcXOmMNytauwycaYwqmq3IL6ZtjfT+
6HgtBb21gbEeuvHyvXu3jjPouvikegrOiLubFZirZQbFnXNoISKkOBaOprf6ThEkUlpruPwNQM03
e0IjxfC+kEjPpjH3tAtV/l4siSIalKOChtPOLzrYPAwvtdOikTJ88jO766E5BV4js5q/AbyT4BTa
h1SyPkIPj1k39Apu2zXMFLnHjwZJaP3dpb0G3GEEbA4izCLwWUjovu3rrs5m4sPd8qmjQ1t6WRdj
Ik66BmN+4PkN4fDufYTHYjRnJx0HtoUJ9hp2hOcVk3d3PTMgFgIPgNnKn8jWi3z4M0lWdiqxd74M
kP+o/Kgw6mhBR67f+hyILX+ci/9f/Vq8z5MIPYWbZGRZXOoFJEo/kBO4UUI1QgT8746BK+lo7V3K
Da6szG7U0ezwWvMCexRO6joel+GnEwwCuWRNwNPxeNjy1XNee7ASP2fRPNdsi6hOAI6koChJ1yqS
4HYUp44AxZBVWKOt7BOXzmRaIgjpLrbpzJq/Warh4zeC/OYHciriL6Mu50RHCUJ0CLQjTtvJ24lt
n+JTMH3mm6WBMayl1ceA6SJWLJWHw5Xy8cVAPZi05LD45nkXjzDV1C3bv2mOZ9tZB2eU82UmXnH0
adrbNhZLKpgg2rtZtUZrvlPpb12+tW9pCBoZpO+8dsx2jkiB4MnPClaklJ5QAnGP+NMAW47Zo3Xg
V9ZVejJxx+zZXYL8KIzp/YzuVkfNiu5TdKb2xWOAzY3oGF0h91rZ7QVRW4F5DgxwSvCgPWwlXTAU
NgXBFvSBP4WAhV+p0Z5CuFnihBfAiC/MWOvZPdv/XiYjBpik5oZM1dsJ9SZhJufQ1fQ8JgHOWLyc
z0mhc+4B6zGjWC7D0Zyh8m6c570gfNtwA/mMuDgXW9JSSG1xHX0cjHBGKwuE0WluxDa514Oc5N1a
FhdRIhXcwIUCPHbtPGWIeijNobLtdJPxirMCr79ZjouZFh6JYibQYeWbCCs/+sGVADRxFg9LK0Z6
05zrJjQRXBE+Fk+0k4u4x7L3AEVxbz61/iYkPJA2zdT5TWf+ACSaG5AuHhEYKaio6hcVxaJwikcv
QbEZ3RvpiNTQcbUX6w6T9I4uVednUPYM35yEe414H/K5nxTErQTYt4ieRibbGxzOH4ZdYBBwqNDG
/k0CEdjBZ7Lsvg/dJr8EKH6tbYnwD4wm9mULtI1z97NR4GS2h6fz2mdtafg35HZ94DV6rL5+2lnh
tkW89lnZzs7GBZ8YWszbWGpvS/Cx7tuDb8Gj9M6mNtCRnqi0TyUnGhoU4qVCnNMbsuI/RrJ+UyJo
IX0WJn9AZyrDMgK4grdB56So9iD8lZUiIoOwNpMmwmigvD3WafnM9ZIee+nBf+AcVdMruLez9kYO
RptYXNAM421GV9cmWD6UmuNXjUAJkuReI/PJkCoiQDmTwO/A8EmHI7+GDsAwzFxPOEUDo4n66vtq
EG2jwMn3Apt6KERcJdyicnqI7Oqy9xI8xcjNxSsnv2vJSRHy0cWNSH05L1PXOHKP/CeDUxy8StBU
3jJWz1IdLt516eWyA+oCkqIzAaXG7pn0ktJkCJpCtAInX/nO3C1oH1wwj3+rPBOQ0P+GtKQhw+jI
M5FvRIaOWRUhlH2bA8sAyRihGhFQVQFe0MDJl/PlmgRI+vOp/nLNNGyW3AejyRuU6y4PKlaU/4Yj
0vFWyUbm1XDrUtJ6H9zm9XFyAYbzgtQIAQa6/+E2OsdGX9m8+jZS84+ttirZfXJPk85juE7B12c7
32D3QWIBjrYb1LNepeOVi5Vy4OsZ4sRV2aFQJEfVy2XJbFJhhZz1/pmn3umXsptvNl+t3vxl2aIE
3qkmLTICAHNEBIHg8n5gR5jxF8itfHzPXHVEz6FddWZVQX7yVqXqz7T0SfJct3pROT8qBpLVZdaL
MKJWlTB2MRFxsT3g70ERbqbTbG+9HiE5YK7hOdM3J5DKAd8GLDUZ3SWzIutSyEbemwDHeGpkT7uG
YokHtm8Tj1L9YDVVFMv4akGEma3rmEdkLBlE/XTAKWWl3ptZHzS52gUOQI7mR9ZeSkGETG3Wg7MM
jEef4c4xIWkQk3UC8/+qUSybdZH3w8C59zfIFRcBEal7+MaTglMr1Kkk0ExIRHP6eSvN2Eyt5/bX
GJ7Vy5qgGx0tZx1Jzf/G1Xzob9racZe7BJbFbFvM3tI/HljIaeWAZt2k5PCmG/itVyjq8uJZAAUF
RjKZDcVRrclkMyPz66jcJuBH7zu/fYzeeD2z3KwvQFwmagcqOchrnPjyWnLf8xWbQW1KO+7NUb/B
0S4pcCvpojE3D0ho1X9VcqmVkphsG1JbxAeQNdwyixqPBJ/RZzZszz/PfPtALTTMGqbNN1zKcaJQ
6O92qeL8g3eo42yirr9doP3D50bLPKv606NfOAyMEu+rvwfI1QDU/4WbcLdI8kCC1dp2upSE/dEZ
lsHzDtGEfVQ+isGeUc3RjfGhSa/nW8j2AqtnTLBth/9+F6JBxtmmahcjKFEu5abfUzDVf2Dtivxz
3bqKVaGveEDHV/Z6GvwWbpKjlihPVyCMJYIHqupslufvavAB2go9TUPCUwEtfehPhebHx6goGLSk
iDxtsDv72Bega0OqYjJVCDwyqCOW6JYvQp46NSVRqD9OZ6R2fC0KF9haNwmzWOxtBOCRveHrYw1B
bFEGtkdm6Zw8L9t+gZ3qXs5xIunroq9iHQ+VG9nelyKVGlztFsvaqwSEbEVrx59OlmexaKn3HKdY
Lo3SX7vLxoAFlL2d/OSR4jZ+U5OlCNXc5P+TWeeFJGjHhkUyZBJPGJvhr9nY/LA6EgWy1YPw8iOX
PEUXkiMbN7m0Z+CztZHP4ko3QrztmTYwAcYb1IfyrWZcxQfDPqyrnmeSQ9CeokEtWV70NdX8KyZ1
+SVOEfVxgkrt5Rvq1tUTPJBcUbj3L0arcs2ihUBSiTHrbNnMFjZ2JMNVPAhXa2zuY4WAvBGPl36j
GKAgJH/XcXEw9aGh/ES05ySVUDjOGjNGet1N6/sQSfHqJGjA6/gDyPe5c0wdQRtnOy3e/oZ5AfL4
QVoZRPZv51FsFKZfnuGdqdq5jM3/0APdtfYHWjd7mvj5BlTl7szlGG25PGqIuIvCNy4W2UnmbqFD
bpxC7IOFv/MYK736lOF9nV7RkqZEFHMKpovBwwW78J3164TJirJCjFvbPrOulUosDKcA/cd8qI51
8fRStFY5rLCH5TFIAOm3IbQ5ko5ir8xzd2d7EhFydQUPXPRr0F7vKEMibmgujtxhvbqL+doywMXk
qXCKJZrTy50cJIK8JEpUnFajVM9AW/ZD2IozA/O0O+OZWkcLnpDXmnVVoqUj79BQWcAErkfB2TpY
8xiAuTphsk6kp2Z+Baq/tlwEGTouIpuSrirooh970CDT3xMVS2qUloHuAJe0uUD0hRWISGiNZQNP
afse9luQWytBqfa6NqzIyICY1jOiMf41mbvpwKxyQE43DYi8Vww6skJ5+OYw0vrysyzQjv3ToKWx
t6g2ER/9cv+NEIEdN9sR36gkFdzVExGYPjLLCXdm4i3L5aprqzZ7XhXTsF8KXKEGndH9cl5AyszZ
W6QJRDUshcOv4X/fjZPffKPPpNHxXeTt0waWY/R7ugz0pR6tLQ7OMRFWh4tXMzetbISrSHyi+4vC
enUzCpjkSGdjfJgDwQBUB9G94keCSKSZ5h8hd0fJjvIrw6z4qKmJoK1SLuq9jlwXMLuoXLyxI941
yMLUG7MqThU6xjXjtCIYBr2qOjEGUxgQfQBE4YZQ7Y3MIs9NWcW2Qp9klAx03wtFqtnE4iefOOVP
YoTG/FyTFg3T6RaqQ1Y0mNl+d0Yyk9yD6DsNsi9M/AxEJGS/bM9134BtTXreaJXUbs5Twx0ZsJKe
6GKvnBI59Ind03Ev07voK3hmpSB8HRiUhwopX7xg5stv23hxlA5SNm3hgUZ23PgFk2KIrIbaBAGm
KDW4ZHkdoHbgG4Onkvc161FcMmNAhgJ3uYu8aMofrLgKKS5mu+LNAWACdGqwJflXhEi/5g2PJR1k
uPh20ra4c+qRYSs8bLPkltTLo5Cbc16vR5a471tylnZ7f6q9hUh/Js0If65NCImDeWY41iwwck9o
ly3+OWJvCKaD0tq7QzvgtTsfF9Jap3L+Z9K4bAE2UU/4Ef/uj4PiM++U4ko46n30eYz/ApGuvtaL
Yg/3x9Ue5DFiSABwDxK+xshJhObnqKeIsVdD24eKip+CVgfdyE1cHdlFS2Z8CdY9s3Go5W2WKJSw
8OGDLA2PphQOrfFxOhCZBZpPTCyIyD+o3oxHXo++rvta1DtGnuEREcocuRD2950ZY0OG4cjL56f/
QJx0T+QffEbQ63p2M0mEk6jMtSMtDqOczdSNHCniSsB86syqg+sRbPHxR7jFaezjKlY/OVGwdvnT
fWz4SL6Z/7+qZ1FoJuPsiCx9eYgIZ/wchGztl0TxCo+8uEgCaDKF0Scr7sbfiZXpTwk7NWifLKTF
PcoQMo8fPMrcQhLDIQ/oVhfMg6c0zl09xfLG6GX/eUAQimCV4eUE4aLkVhCYIQTpDETBWAFx1BaR
MdrqP/9tKP9M9stC3qxIZiUxgmnKgkfeQ8RGUxtTsea4+PLo/TXAr5PMnGUo+PCiHxAWNBo+Mspj
SNINjt0Q3U2mT08IEjTpGAmtb2y25WD3/clSOOoZr5xj8Amd0qErB+5pucyma9qP9tH1snXepctL
2EXDMq/SzjJ0cR/7AamO9uoK6ts/j4JSvl01vvRmlxY78H7pXhWjpzWgdg/ckwkYJKsQ9N/knvZQ
bLYRa8AA7AU1jz4YB/4uTu6RCEcvP24WIVihMIcX1edOknDERUOK1edfjikF059n65ABqOU18cV7
fxqzvVGda7PnmU8Cu48bfj9vDnFQbQa7L7X4d1GSXNwWg50sL6nO6IYPJAIgqEY2wRiTWRCQrc3W
ThrDB/JNox+LOeb2KUdRmt4mh1wlZcSYl/LOFn400kQMUuygqAQOBfW7L30wBiEji4/F5JJ0TsMz
eOpNNXPzJhgPQ9AoxjdK4sBrHvTlLkBu/b0Pcf8I6e8rdeUhR+YL9mnfu0xSy9aH5Yg9y6tUtA/R
1PJlNL/uv+WgqhDpRvoEFOFOi+/GKifnILkBOJ9S7Y5ZBlqZ0U09hQojgSJYdOEi0tPYGOPfzLWz
ByFTweC4VUCTA49ObkkCqTJb+fKgmVbmzsuE7NWYpDZ3FCJkKEQeHZCltDt4gy+FDLi8cafjKtDf
AhwPT+irWCW6zd9iRzhhE9RODUP/K0HifRpc3NoBVZxEhCd1a1gb4izZGnakGFs0QQ3gnGT4GvaC
ylPP7LPuO93XfI1ckfN0Odt0kSu7U8KzAAy1w02v1ZxOlFuUaW5bJW0gI5idv48WMo67YROl+sYk
t80RijLLiq+bkYEbmdWIJW0nNstIT2dnSkEWCpA3XQtRUxH88oEvd/H/QCPq+vbfet51xSHnSjfg
SvjIQ0jk0tWVsjEFh+h6AlK6hnOFOEChlHgZNiLt0FNnj5d5ZVv23UXZxeqJJz49UcszdMZufBEa
mjErYu+O0sfEY72QQ5f5XExQ79XNcp5rBbYgS6RIp6HUK/P7hDl6aM89NoZzrIQJ49h53Kn0Nr7e
bGo/DJZFZ36pQZYjrmOsSCZDJzEbw6o0fx2w6FAlvgZbylMqytqv4eYfyaVhGoBqD49m3ak/ugV+
LHPR7hqf0BmM6BSrEku8mtwrTzOrng3uB2L5TJuuWR3R0RTlW1lU064OszsSIE2/f5A9rR7goiLM
zWh0rCaWAbvHvz5uaVBsk6FYSdrHB5t5v0uxFPVmaP0/moBTnntPSS82X6b38UEE667JS2qjKWuy
7Lz7m232EMa0b5t6P5wrTEffJwOqKY5PuS5wId6wGFULdheHsCPUJ3c9I8R3XyPEArxpVXxQBH9T
LDKlkDz8S3PwH1OLJzcOgy1gqyEC7b0Y6jv6l8kfUA07+ZYZ9I2OkcKx1yZRp4xzRAx49Y/c43+B
e2riXc8W3KGxJ8yAmRysMq7qhusHGg/GVKgp/fn8wspTUlGvN9JKYeJbRz1q3J5LxZf2A3Fk8KYi
ulSOMZngAzVKUwvuRPk9deDhHtsh7m1ad0nvCW0YKlCcaXs8aMeofwEvvLd9X323ZRPWaUd5n7Vc
u90mfnDvYYTXuXjDQXs8mDi9JzgZ0hyqY2XhbsGEHD7bzc0OOWxuWv9Aook2wN4pFsVLLDjAV0R5
yuT74cIBycSnKYWXecZEXH6Sux23Jo8YWo++Hi3cN1NOUUsncKALzxQFjLYIxim/idNBdr5WfxvR
+tSBfNb+D6g//lPhPIoteY45jEVbmF5mqnLx0wU734tETKbhKJ/mlhWiReXNXfGvAK/KXfVUtUtI
lNlYnzCH6FYsdS4d5zKm9yPB96TAMfxwUzcT8+tiCU23nmqlIxkuFETh4kLoETx8tV09H1Bbt6zW
/+UsWgDMku3ypmdD3EKnxlmaYSZ4XKV4zH2XzkwtJyZiCEpNePgYFJEFtKk4WzIgzA/b3lOEdqo1
vH2eQ5sW5dD3CePmh1BwfB75WVfMyXO/G6VLYHSAligDGsYlbEciPMHRdY/KHw9UKQsheysGTG1r
sg+H1fzpkHDtD+vDpjOFa8jmL/hH5sTJ+l6anyn7/ZmFKbSlE8T7ipZ/7FLwozN4qKc4W6A14tz+
GMJTsqV+f89fmNGJvRSPMouQka5qLcarchuM4gXgWqF9+neXI2D/6MPa3SE9sOyALJMq5wDq1GFv
2m3XJ94f1GpxQyEYBVwimUdh01hUrrWp1Blu6t14DH1Lej1igpOirmZvukB/tCdm//TsTMH7vj+6
vS8FkDWxBfopn5IYtkWodnBLMDSBBfqqudBpFIiXGEg54/LJB1bD0Xh+5dTDxOgjJGJBz/8SRIRo
DZyNsL6mNGtDLnzaXHH0i9SmaVJLRaw+oG+TrgWlpfb1P0ctOZ0t8kLt+YCAAf710p31mulkimRw
OhVzQCBJOVUhxYn8eG/GJDb5+gHUQjSyPS2tID+BK/9+wkRB/cK8UehHEq6YJOEO9Uvl1kEl6ix7
sZs++1S4+j5w/8T9s9iHnI09y7otdozm7AVoguGWDcYtDZ82/Lv3kDHvg9nZU4C6hDRsQzlHGrIr
JtWL5hoF7eBbnlTvoCbH1QcLxGYfq6pyDtUDoApHJ5IklBcLZnPG7jxLmFwIWvilq0Y+vaFbISoE
DXQslx/C3hmjjRzKEt9bF5UYqloiNzUSGTEvIrjc1QTvQ2pDcSL/IjfNoWb685GdY2afrMdYM+Om
BFGeL2XJb/qmBX1MxNEOphZHODnqF3zKottUPAdW4SgroXjQNl1dDlSqedkJrNnCiuOjBIBan7n0
WWA5W0ooebncjJ/c3BSi9Nswn1WbhPVvuJiXviHJb0Qe/TxiUGke4dLjHscE9GuvzTrKYdS75r0t
i87Zzht4qOie2JeRlkitDjYbnbG+qvqhyo5GOF/imHg3Wop+uvdBn2Duy3rOvDSojoMPpvCheHcF
cNAce6rIx+Si0uLmqF2fibxh3h7ei3Y2VCjS33F6ZmsoGOrprhdIYPiFvi4ctltlOfSABNZ2gbp8
sP+yjT7ynXwC7L7XN7wkf5NdWb4Bsgoxf98CFDRBkCIJtEhGCxFlvH0WnDuxjoAlPVA8Z1E1DR+9
9F1sRI9UZ0qRMTnS5hseX44T01UlPt16Au1OaAd1WQHb6cc8j5CumOSkwdc9Y2LbB2v0aDQ9mVcB
+WCd7JfUdhJ0WJaEw/3c5MM0mlgAS6TimoWDtdh07Hnz8PTpw4eWwpMxCLVqqWsrQycAVjLn4zw6
paj0apdDkByczAf4+B9nfsBdiLWq0ikXyYCrgCvvs9bP0P4uk4KKVGnmu3jy5qmMKLvIC4OoL5mS
Mlor59XClpbASYcaxV9uz0TPD5QzuVEwgGF+LgQsmFqLj5roSFU8ZhXc1GBPqp76cVRMoTvJeoyo
kFfd6qHUAOtlPyebPAANb6pU8m9y8c7n+HTbFW4rjcNYEcLD8cvGoKpS7XtBlzHb1pbCaRdxeQao
WMdcFFoQ7cuAEt+GabmEarnZI9duqceArHhYtyOI0+Ide43lcrGGENnHqTZngZYWRtU2yiwNPu7m
KOaHWjIbGUvlP2Xg0OO+9PLPKg2MLRbh6DPLneAPPol4OpudjHgFdhnJ7jXcrQyfHl/WLAI4dYif
77F9C5PvfuhLJ2WVsJoreDmctExC56pB/iZLm1YC24LvernrgVbUF9X9fXjY9CvW/OKJ0EgTUYkX
AxHsOAssfWG3QARvCRWR6kTeSw/JtvtlsnfS6iz3YQrAiNAaaimfqqCDYvrozg5//26YAhBjoNwA
6CrfPeiVGhkJqkH5Wae/wGiL2xD5oHlEFNBCzzdmgjWhkAFjD18am0GD8XucyiwnjkE38qMvDM1e
RpDbVH4XkIU8ZgT5guhJ4V37znS3Sj9DUtJ+vmWUphUXqnB4wq9oRF9N0HA3rlGllJ7ahnostDRG
oL0vQaLrzK28/sGolJsGSJUIRg8moCJnz/R3yw1qKhGZ0SQ/147Thd37odvdaxSLz5pZShzZVaC8
WDkWzrVRAEIJkASHmrP15bOPlUeawA26+8NRx4DmHeTecbhEkOiMg7QdQbLlF+BdCZFuFdm4i6FP
A/sRsxbKEbAFcN4Ysw1aYbE8Vc4DGrayBWnkqFSMk9v83M3bWKog2JYPXb1rL26Ljy63fpyrdmFF
8ttO9jSDLlRHTJjd8ZL7jXaut+ghqHDZgYsbwh9qqWHO6B0DZqCkrT3WUs0Sbs+ZCf7wzvr3C4B1
kK1Le88RKuT4i7OfIGyp1+7Wq4N5HmNn2V+xTa/SzQuL9a6MrRVzqlTp4utI1FKhYzqrg6qtoLYy
2a6dxfEMTfXLXmBcNoZO9LnTC3++RVqivsDbU3asaIlVB2wtitO5dEy6jIJRBYvYrVGJAKwHkySZ
l0wqs7jP8Aa4503IjDCVuFhv8J2aenzl9WLPcDM2WT9a+IUXMcV94aF8mncH3A/KyNj32x9zTbis
PB3YImXVmLT0STFSy72OYZDhqVj1qxCgq0Y4wPYQSFDhinI1F0xe6650jW3DAKZSEasCgi5P1cby
PxoC9NQrPFDVdn81bdTjdYMyeraC+dDnsS1oFAv0f9ri6KEgcpb24vdPgFWVs3vT2e1kbIVfleKy
KnBsJeVZyb5hRZJNaXWtGJJSUEDfm/yOFb3WXKAcvfxKbsjsQQQlCYkYVvAqAlgJbjC1WRoEEVOa
g7u7CAbe9dLnt9MOPRjtUZSy80TVapPn1wwMF8jJNj4s/X/Yn0bi2m1LE2jHC4wBE+RhN/7Ohkxh
0+FFqwDqhhNthtOBKE3mdLDYSGBFgTDGGhPCiZCcFwMN/9kQUy4gBGBZjUugN2OPqpftZ7kzrERm
hhRzC9IobIUUbOrakquCysJN0MxLMKCPQy3wRKMC7yO6DVxk+Me9QrVkreOk7UiNwX8FmCSNH3y0
pbR0CBPq5+gZljmffASAja6m0YC7MEWqPV79+KNDP6SdeRFXqPAf4heEUlD3lUCfhA0289TqSoiQ
2CjH9mBq8i3hqDDLGCQ2LVYhwek1m6CsR0RT4ZRenG0c72m/6bXjAVT6qOzb7PqR5FINuzZ/wHw6
mF+7iczifZymr6a4eNPqG1vccvbTsyeOE6MqGKCoJySekdVckzrmEZjhcM2eJHmLvQRjyFA4sTsz
C6UyogUYPX4KNUaDBUOoyNOGiE8139/JGmmsns7KV2aedFhEHTAgA3EOLnd8ocujRcaYft5YxqKs
1W+fC6NXvieFcZ/7VYMOOifxBuX77xhNKYSkGk1m8oq0OsPzucMFcX7VHuMbHuumrBZ8XN0v8FH7
wK3p3TCeXV6feuVE76B8yw9njIlMoAZKwxLZQ1mqRhE3iPe2LPK4OAV+unp73Osj3OxsOhBjH0iQ
1hHYEIwyKD9YPSRBu5CXzRCNjbMDfubK93Cj7J/93J4OxPy/xiEHeBK/D7tRrMv3Yff6On59D3Zi
/jO4nOz1PXj4nZCf3MQT924QqfsgUBntg5J1Tg8sQ0c253soHKYT6UJ213+2Gm7zG+hIHNYnTc/l
o3KICR0bOa6tCeBHef7/x1ggA3+1qXjxtyxxkCGQMQHdKFc3sorMwSXoAXvhZmkKH9l49HmuaA3K
ymK9sARN71LogCL8tyuoRhC/2UfGb7JU7T6HXv1KZjng8yabtvY+vc2DyR3MutO27kyVGIxNEm+/
RDEk/jfLrsRF1B/lteQWEL2INnHOPONe7AvRScsVrUj0/tRM92QrApjBayCxHM84OgqAQTDnEj0N
kj3LVFXzkYONRVTPvEWWa2nDmB97kUP0zHK99vuO6xPKQXG1lTngHh+9yR05s3s0CX6yCErOkaG0
yECIWAl2ci2+f7AbTN54Gu22WSnbDQjOFBvEfYhLTQ0bxo8dFcQIRW5LgVr2W8EUxUELgmwtXW8R
zHEyoPAoCFJuLgTllV5wx16M88CA44CrTu3dQoVGv/8El/hcvKe/amtD0x3DFMw9BB2HqDmISEg+
dwF8e8sFa2rR111u0MsFOQ5CiJEyG4ktogUU2eXeUf977ml7V19WYvhjw3nhXnHJwL8ui539OkpC
qIIpSjdfL+UbBxgJFEfpIomu9ChD3e5Pl1YIK062ue8A1m/+jbftm7SyYI5TVTI0pS+JTwXDO7JJ
dOcB6prca243okKgooERw1PQyUxkRVib4aniE64QmuEF8mvVOcRgf80+IvgAYlLj/hnkU6ZwG9xJ
2KY2b7O8rNBaxv9NkBwO5ouGyNkHWkPhaxyCSUzswVrWNAz3SMNLPKQA39GgCC3tGm2+C+vYrQdq
xDjmwMk+354GI14T4AF2S53U3J80ea57rh8tQEFABtmzLfPvAUL/rOQPI4HLl+ksIMSU5VFRKUiY
1MlEBLqw4dOvsBkTWNVBo3zW41nmXnx3VeT9HFMNmClqDeVmqAesWQeMJisA+hDn1CF5elWCZ6aa
3SUSlzADQXBktPL1FeoAX9U98lgf5RK/fF5Neh0guIiGcmG5qJewGXLziu3/hVcAEwI6RN3M9VM/
/8CM3tGHsJlvf5T6WmfOSkm7dGLcGv2ZN/2mVp+WedIRZghylaHA9K03f77CyebWdQu9aSzzoChP
yy1yqlgxlZadQNz0gwCV9f4GpBiUoUc4xjiMy3J+ifekHiJWTVlLYLkpWRq7Gnbz/LOUGhEixXGP
6dMiqr5s03cBhfbVIM03qiFM2nUIqQpuMbwVlNLfkNDNpHseqMh/KeghMFziAlZDqyJHAqa2Eaju
YRWGhoyyH6r4CFKaeSycBEFg3Fc8g6Get86XCQKla/Aq0Mi4BbtS3d9TT/MOSNx+WNzX78RtCejv
bTGSHfHePRAsDX04z6wD28t+tSBJ79aSpjltFvTFbGSE72S86zN2yDyhjlTXhuhbW4znbTfqs+v1
XR4Xkk6w56FDKDqUGYRynDXHouLbyllnwCQr+nRtNsrnSZ++FLfNifw1dP8VYiWUJSu1tHV8NEog
01n4YJ548uAzbidsBn70Up/1x/cEA01XskyaDIgbRQplMBkVdKEFuzsn4uPkCyQoobiUIPy6q5nj
I9L8ctanjYQCPlDCVuEXSA6YH7PH6VrFc1MdjNDi07qK5zbMe6sh41HcrrkbZ2j2gO7GYxAFtYKB
9c5RJ168jRjaT5aK3yY2UVMtIFM/ra1JGRpE2MHogj/5s7ynKJKjCLV/Ffy4CEr8Bjtl0VQk3g+X
vZSvyE1C6sCLdW4MBWuOwJiNu1LhvZNpuDFP7d8Qjs8sRqVwDqtroYTDpe4IMdd7BU+Q4k6mDujb
rhylgKHpbhl3EYPAta+yobdyUIX+GScx4f1se1b27RMJeOkRN57exRe5JvtWgRjppe5W/sW43ibb
jJItt1uOtwXFcWQuGPgTtM7a/FVM3PG+AgjK14jRkc1TrlhzUPOS77LgT8fsa3vc8c60tN0tkOD7
1PeN+aKa93nGEcoQvgYo+8+ww78AdH/Fxf7oJt1SHJHhakFVhubvVYrHKLGx6G2DseiW57s0gL+b
cp7mVVVUYMEKYLdrji7JCZsBdd6u8gxMy3JLYbBwke9nMm1uUz0vFfVDaSNkT43x4GRU6TMTlOL1
rZez3c1X3gWpXio+dwcWKX1YFzFi7z/OQh6hQ/MIu1xibvjd82pbElYto++VOU7vp9Nu4HqyH62h
0JDuWw+bs+Wz6tpSnkWbvWEi4QI500RLM/SGLqTnhAPKEZ8YRBHDb+qd/9myGwAFXHgfQ++CPwF4
984R+SqO2pyYdmmQ8fSX1971ZNNFNtaoqx+aty3Y3s5Dv5enerpk2IMnETIy5iBRj1fB6rA1KKeD
xDgd4pqx5MgY54g5fvk6f0WStPsfdxBx1PjnG9zOPJ/65tMYXDppM5TUlHqdAb+OsEZrEpuyUNiB
oczQMWGPEyZVHmIAW8zHcO1S4lzmXg5F/B6Y1oR+D1qZkFvxSsRI9G4wzLsPVRnrB+mOAPLI2/xc
SgOYIKCOQySrvF0YX8sJlpWY2f51MPWVH6eCXllTTosgboR4Nm3Xc8gPXI3YYcvT2TfD4SI9qq27
I48Yei/GdoaDxbQURxhduaHJcZhgARrcO0KKsutMAns6jKgMdHN7IfPz7y5NWBy0s677kE6Tie3N
YvoIV+WvxbIsCSqk+NyfljuHNvW8sUOEstsIYeDjA3ByiVo7jac8YV8EenUZHwa0Dm6fTWb+tVtP
19kPu2duA8DrTaL4Jbl5DiS8UaTSvlGBMf0jowIvVExvt0lbi5o9VD9RxzXCkoBMlcVPSbksZyTO
jOHbzAl8beJJuWMjE3CUv0rPK5vye4uVrhHxr3DBU8Y9fksOlsYzJzRvhb1C2Z1JVExn5OYMdYvH
IEenGu27a3Tho9nK9a4cDSaio30gHv8+fcxL1sMdve/voy5jFBJJOZkT9FBU95TSHFBAHg6kuJlk
vmyvcRSlTemROfvZRGt5GcA2QiaT/DwlkiIG9lWUX0eTCKhTIfy/lk1Yd01VYhzNu+C+mZT/FbZz
IuJUG8l728Fvq6CTH9oY+OuXAVc7h+5vo8BuSeUhU5rWruvSqbHSTMeS469ICji6kuoxXx7gvvcB
i/7MV9yqG/DEqAZ5lvR1AfnumKtoLmsgELGSpiHDnWEW2nnM0RY8LyIqKBwFQRnf9Q/sCfMk1E1G
wFF8hAUjoEKYCN1RhLthf+ykz4cM3KP7e4XaRl4iFInQBfpRM/LbmvzuY4VtGQXNwdJ3PxP6Qy6C
9WQMEXBlr5htI+Bq0pIrQN1sWWspTjUut1F8n3NItaxIEf4dqIH7RhFHimy+E2TAXaNg1x4aJbeA
GKvRXmARQxoBtWO9gt6r3e7ZjMSsJymvWHRo1o6buYNoqkVxU51/jjsdxkIhnTzloINoi2IE9d7K
AhZBE1aSDpxzo5sPGMm+EtWC2q74uwJdXHju6QowAjXOQRtGNQqcf9G5mRR2BDN860dT2s+9sxvO
xB8L6JlOG5Lp8e4QVZ6wj8BLV3wLuSfO2Po3+/7cIVTfFri3epX6UqpEHZfDI4EjK0M9tRVlmjkp
lhY5VvXjlgSMJOI+FudE9HMVbHdTQiWGDAJMEtkkRoCHsMYb2ZLUsEyxzgpvk1mPzKzug0yI8RcL
1yL6e/4FmhA5UL53vL2a5sgcAullZmVKZbPwl+vOW1dJ0mKsXszumii5DZrVRsVCxM36SOucNoTE
9K9C2AlO3ZbCY8gWDVmsYpZ1wqk6KfHJTZh4LmR2g5w3tz3yvQODc+wo3lyxZ+iZ/3I+iBLJqRq4
ZIdS1uomJMil3nRdt4i9/jOkl9EuHSDLJa5c0n/CGrRZAA0BaxLaeU/76myCTlnltQxYtc5vuUMB
+UeGhIFFEN5b5DHj4brLaN4iT2BJKA3WqKZUHDEoMVsNEt1us935azW2HiyznO2aoGr9JZpm2sTW
nCArXyr7581hhLcHuOgcT7HwaQ+Pr1msXk0nbFs8p17bsBBZZHQMzuSlfsRWH2fm77eQtr4zN0UY
6DHCzbxOnPmYNfApwY40MVt3js78mTcXsstON2/KnLosKHHgnZLiinl0woJ2NhHlLNP1EMTYIgfZ
NmoO9WwZQRd0l7ndGxAiDT8lgZ2JDA108F8kiP7QBgbeIzS7ylq0MqE6ze6omCJxNJRbQYgplJq4
54pBznCIeVeMSkpYPGN24CULLGRh3dIP8R0pzJ2R6Z5sm4LqQvLrOxeEKH30ohfpNeiJCKKgdnSv
1HrSz55MwsaAYZQj8Zp6gKgHzWUjT/gT59oqjQwt6gvkdKawE57CmXjRdm1YtzNa1oEDrFQIKEzY
z8kBfYXuUnf/lbl4+r8vFPyP9aW9uDE/CR+Qvu6pUX5+JjdfY30oQ3fh82cTO2gMu1E5RS8vinNW
91LQWG1bYhHpdyp41KdgVzCtxt2xPtsx6SsmBRXWdysQZWeZv4BlsIpFOiXqwaBfaXnGzqkFAvq7
Xi93vsd33+fPiUsTxZ8fUa8l+dEl6+U4kOV2fal14LQKARRPLVpRjGggIKR19Qy7CeM1kL3iJxAd
XjJUolPj//q9t3ROA3WczC1ieNAG4kxrF4znDDFBtZkeP1jbiSk1D6ym5oFuQ1YR1hITefVzzOEx
7sLhDRcQ2sAXjdmlm6ST6I9Ag91Sw5aJAZL1OntCAMKpbIvTL+hHmE8lHvif0Vx2+F0JdgJTlYix
1HMacyusICSlsfXRHrKSKt4qySQsNHopVnw2jtIk3RFaZm+QxD4P4uNd3xPgdjx/+tKNj55Y7smZ
T6idmNzmzAB0mo6hsYr8sE3A2FpQUv5dVvuYkggrEyC8ldRt7YtL4TJ+lcRy8pEUJHn1xs2tBH7B
Kc5/4mq+ZBlMyBW2fw3b2kyyYomL7AzMSZeZ+H0vMfgiIM+3cvYxccTnUYCkhT3VqznP656J7lzB
wX0jE11A8rkR2muFYwgWlbhocUP+/cXp9r/Bj2vO24nmrDCNK6O4Ozm2qMl0kTuBZNMGqSSBqxiA
ZQDuDFDrgmYSeMEw1YSs9ivFIgLpBE/ZGo/sOeX/r/js1hA5+Kol4XgWWFsJ5V2AJ5NVP8yllsKI
vuM78VO2e2C2sbLFd/e3asrL23trjSUyxqH4NBWlU53Eu+KEH1nRvsT8ttdAioGvE4n6NB44wJ1D
nV3pIYraq5d0mPkqu5K0ktVmZrPDdc/VKeSw56HF+CFZcjCCoCJG9pzUU9sV5eik0fJaCb45oKZr
Nf2MOdBIPNv41vN3c5oQFxsqwQsxOQ/3avwvQoiaAUmTLruOzN7fBIxG+clMr3HXOzwbSO3danzQ
vAtzgQlMI6I0f7wq6Nhztf/+uttxQ1bKZmZcOkrbxpr7F0+QNO8KdtksCdfr/RlaYI3u1eJ9UxWS
geV9el6+4EZKFrZ/ZAIdzuXCConoUvKIDndors4Ggbqs8WnItVbnpnK5E5ktfQGNEDQi9vhySTYz
R5Ci4nyYC9VqxcGNbIVBYa+IFF2i4+BIvTI1ryCEN/kQMpM4cadlYMI6oGXiAUAF9dBEW4MqNubl
PCFpJCu+69UR18O7bhpxeVMXgPYURE86IOrmMZ7XqzmKBJGN1/Nk3fY21EG5B+gIHmd46m6ApE0w
J+QdRw0kXQUGdL+JgL08Z15kqGPw9A2/NlGCwuASV8SNfu3pqJFPbEiwf64whb73njFxhq15uSkF
MlGEOpGmEDX/ZC4N0Qn5SPfbGOZaZqZFztsoInHwDUo4sqr/7ps71brnfXl1zTeckUnF4hZpNVbO
wjZQb3gMEseWjtCUL3mEcD4d7cqm6+8VJBNylXZyvdUVircB66yoYcAUVj2824EYoLbxQSbcSHro
8AYEnayCVl3p82UY1iZ/QlV/smc36u41zNxacI8ZE0x2Z1JWXcaZ2vZ6vep5t4QwyZgQK+bTIQno
zksjmbsRwsozsfoqmTbrhSR9hJAZVL08GJaSu5cqSiG6T4hukVYUGGX5PrM87+zSKyUUTipqqxpk
XQOkaCqG7aqoPm7XC7i948bkkI4CXvuIH9Braf2czydCAmvY+7ZroTIiBRxLFZDTDnX9GCuIYkW6
KGvgoh6iQV1aumm8IQeP636lvXo66FW9/Zh2wPCnSnF6M9yyaaUDBsJRFSDHvZNX8gAVVqoEf9Xn
zLbedDqC1lr+K9OJ3gnDtd58Zx9u1caNCeOEOy5LBLsxleccGe/4SR+3x6wZyX4HUQ0DXRNQDC14
4LCXMT2GYMP/RQc0HjMOIj48VM2SovMCkqyBFQdi/424lS20nnFox12r3rfraZfxuIPpRGJ+AfM7
Bk43w46Z8UrBEv78hHv7WlD3O33yF+ulUxyKgCv9zD/zko7XnYu0Sitx09YbJGyf2cVojaPyHoPr
O+n37ysTIkB5gJ+wGeFR5zZD1HMS4eEUrP3KyD+33Yg2sfSQG3Fwf3hO1EP7366E1fQeoWFYcbEI
T3bpeTlvzqri5gGc7fpBUhFM/Nw/j4WuZ8mEgd6V2fBXz2g//DiHVmbVOoo/xn4HObPqw+7kDWVC
pOWfHNDqaIuCNCsq38+bbQFL4KkWQckiatWETER0YqFkFL5NMC35CU/lhtg4VtvyKXz+5+99h5xU
c9RA/KOe231/KH81zwUx53pRC3CWkXKYWjxZ2tMWBEQG/iDQG43sFKryBML2fCRnvtCpvDw3KGrM
RWMM3HhuFhTX4jyrwr/xFYccyD0QN+ti5epk0YeWNZVY/YAXpBCKBprGbKzFekGgGoLkbHOL63hR
7RYQF0zM/h0oQR8eANtLHkgc3fU2tCF9EDbbvPdgqbtn4dqaWp52QPBuHKFrZKsyUkuD6uTeTAeT
/tq8QYdaGh428zJyYPMjg9qvehJrcUry+pn7gtYXhn3z4AsFLzP/tbr8yjgW+oT5ub9F/iJa6vpN
fbzE3bP0CjD8A86AM8g7/pCGs/Jo1RXq9eKoUw775QOC8Xkb4lVdbSaAKoEA2vWqcjsh9m2wrqPW
Dusp8zMNQ4yZP5mg/ArrbjZV5z/hHcZpAXfEh+3yKcKhVum497plyXhxkMbJf84iSI93Cf1xYOcI
p5uR/BUDCGCn9IDWmEdn725DkYuckcR7sDoYC8pHdx1eN5DbGXm9Th34LRRMXiS+dV/rJAPI1swo
+i0MUKUKcS1x48ph7NPJE6sTH24J1bkQp148kveK4JIIxFaKq0sPg2oZNfkjpVTqQFdIUpLwGnjU
yT3mSL9LJO923IVXvzcwWBDXZtKdVwQ4MvlwkJEa/hh0ob00tqyptu9FTzu5gc02F/QdwAOFxkIt
J2AvGIYsH+FtlrRTykgPbothfb9jZsL5yuRdEgBoXFv+LjiOJaAhg5n7fMqUrCrmq+ydzODwRry6
4b/KpNRtrCSN6t7nFvJTQA9mHTs4tVJV0UlpAIzpqC6iGlXT2+xxPZzKv8s8DtGarof+oeu/ndwi
n30Sydu1vBixfPTnEEfgsPpyWR2aOXDoPoqeg/hKt9M57uf/aWAVEw66ZyDS/0JAdMGPV6OvbB3f
V3LSwwIr95vd5YwpNH9VKYMPNOsYu8QU/A5G/iJR0fNiPf7kvad834cVAn/2hRuXHNBj3POXwHGZ
ikJUVwLIdVqwFaOBjbLzPGPXLHSWVd5Oo3TlLqkbG86vYh2lUthB3dUDd+a31l8V5mEpgHmz+8FY
Obg9RGs83FAXZ7Aqh2/HOwsUEWZa3YJhrCSgtOTyhKJVksverRliZgeerZK3GiW/dS6zXVK9GT0s
6DCpK67C2OYK+Mc5Yfzj9pMg2S/uveKqORFAphBKsM8QKWhKllB0m5SVgCCZeAxxBQfoAAYJX1Cr
X/OesnpF22kgGR5tV5KTTjHqWW+jxTe9WXL2NMsc//hXbTYxoKflPqTpyqAwJQpm+qcsihALOnZS
Tiry06k8VzP8WndthAU6+NZ2m3DC47s/7p5amDi6kb8SOoeN0R0w24RI7Lwt2zsejT9dOOpDfsCU
cAIcIDvICLQ0DqciKCpOtKXzqJJ8RmDzo/kq12WSWp12L/XA/YCWOCqS7CA9kYMg9Hipc1QqAQAh
6mVY++9JctpwMbhOrnWVDRtc1IK4puah7Q0Ed5qkaUO+eGCZBI8eX71gWS+UT2aDz2HdjZwUV+th
8qm4OTzW2oX4O57DGc8ST3jbw+47tOYp0qJd5Yc0QweKmHlPApmQzXBqIe/ybwpCkRhMu5jWty6C
EDOdWfskBfqdaVTN+PtUvf9snb8Xkw31rbIdeOP6qj0a5rXf+mC+xyHpcwvkJVWlaOuqFDPZjpM9
Ij5UCD68/fqzEqPinaQd8keil54Pbbanq6CGoasReIYhq+CZiR7IgC34TuY8jtfcn0YMLAPpd3RJ
odydsqx+fKjPBQSMpl1N0fSkQ+0rrI/b2YN0w7na4sL3NL5d9fp/qeFEH6dky2cCZXsg9+qyOMIf
24QO1nspjtZWMsq81d3Q3PmfA/zCdl4Uoa+VbuffVAGOAiK0uSDIcC0QvZyrFwfmCQKFxO5cJZOb
P4eUZF0JFxTT2sitOrZpx4c/gURNwlaN4Mo42xsBWUwyLfM0/x5TRVSSCpTBwZNxM2EVsSgaf/DW
5HD/iNrdZDZnfOB+Z5FQQ2xrDPZY6FJF2oFaPoCb2dPp3Ej0/dIScOfKZWuinygwxYwgighBccch
la+LNocb0b281YWazNZ3LsCBdwCLUxzd4ws9rH6fESVOda02Rca6w+cubVFNz9ALr5BSrzK7Dx83
hZhSGGvy6ON8kcQ4euKJCLRET+YJrZcvZW2tqCuQaUtPLjEjxJpSloT32VBD8jpRCCioXXYsU52E
EFLmiE58CDdVV+9az49DPd8uirzhYqJ8EM8gyC1yj6xa+2zIIabowvn+gVtmH9tWOdg8piB4MKPF
ACjoNVwY87lcsfnZkxWzj5EiSiKfeNQ3CCLTfjuiBsjkkvm8wJ0iHTAyELaGc6FZrHGLg5Fo6exo
tiRNZYb02DsnrCnY1R+uPU4vOXZK6c11tVmdyKcokWX0drRussL+G8+EPuoxVN9DgqIrYLpxK5V1
a8vs25XzoTe8S+nktho0PMhYpNcuJpHT6PeX/5xMqiTbmoKsPseR83b3QU2Lq/qK3I7u7S5CUI5U
8UApm7um3k4uKaYM5msLOOLDSwobypXWHyobA+DI6OOD99ieNhy2OkHrY3VX2g7rmv94XD7uDJze
8npBtQSt3iyipn7dxjan8b5aZ90oMIT5yCznfs9taKCzlwWDHfxW7Pz8qej/Pffwsphj306zZqzb
PhmNryHzOtIdS0QiPUExgwRO6lZcvRXF3ygE+6bZHmPWjGn9fLifPODvk2ucqpD3i/VqrtenXTbb
iBqqg6U3RAKiBJpE3ARy1X5jiU4D+7bVecD+zO7nk4BBDEGmoniBLvH2VVTll6LEQFwTILAdc5+b
iGP/qNAnM0p+XpyGiJXiRJGgidtAYmWaB/HMkUYLfD+5uFLmcPvtiSNyfEZxCZcHw8w0vnTDDCwV
SWjrPlJ+NhCpxKTiEsiPGHZm/ah75OsGSg54aMnipXlswKes98/RL1BcURL9WDyyUPq0x5UW7cGd
PrlPcu1VzZyBjBbytG6gRd9BU0i4CRZ79yaZPX70R7rU9jTyW78eozSgHXJKjwTtpOvB2q0D6+61
yBrKIZ4DjEgmYTsFsDRk0yDfoCLxGDWPEu6jrh3jb93Pw/fv+XJh722FaMlIgn9SRerzEak3sSwW
xE+38uE0FGtyZ+tg2hjcGLHbokzMs5Bu6zrcTppZymXOe1jN4vprT9Lm4/+h5XNsgaxMA+zgQTcQ
YauEp/KBagoaS2Q+EE+TFGrmXmNBMBhwO8/Thc9X8hOrLaxTiSa7ED+XZotaD5A2XNTvYUsnNndA
+RH9Y31LugSDp3cXg/ZsqfzsK4w1TQeWYYva4X4aHWImApYjGTR5jYfcUULcnChNMT5uFmFI6NXm
p5zISU3MZdWaa/EChM0bwz57kxOav6a/hAWVaLutnaA6SPr0cn0ZpVj5USd/JLooVCYs92hyJ4CD
0HQKVHK6dA4z/6GvNVq7wTZQVtbNYGTjkziq+ng06QGKz8Hey4CykxAK1sx/th+OowGVrdFkKucI
G/qAhmfwqs/g1kxjpeIPhPYV4pLEB5y5G6459L3mh8Pa60Jszcp9IzTbvsBWsnp0fHq7fjpTjf9m
h6xbZcp9Q6V2xS6cZVjDGn/GyIjJ21vzS8AIDLDWy1ejESCGogkDsEB22HKSjBf/W2LvcZbxLQmG
G+WgHqZV9pcbDtYEhHmLrVKGnt1Gmn1z3YrrF9Q95fLHEohKHhL01im6DrLoN0OdVIKsrVAwP9Ru
IbEUWgk/RzO8QgIEJf/Lv2aSXiFvsjM/cui3z7AlGX91Ye1a8KN9ueKnda1i0uctRfCXOn04gXVk
bJsNl+TCLFrWHHu1QN+8UDmINZlM0xh8YO/G8ioh+hLYOaelOLl6re8Mp3ks1HV6s/a50vzZgKD9
DbNZ1ax94QADyGe9awZixCxCwBedUdfEcgkkRpnH5f8QuekA0QqODZe2ZhyJx5f22gErSA4Vid30
fx3Lmc/KfZS8z+s6xTf4EFP2aDD3pfuCLZIhKkMBW+un3Sf2kvXWkgHPsVlXvgdkhz2nC5QcxhlK
VeMPO88h/7ReA5mBMyV6PAv2u15nj3UzBRLsOwUKujlQOwa6FzggVfdBgMclpEPKeNeRzUSZXzBy
HsFA472eG00KV2C1CBBj08A+rAZ9wn9JJey+fmZ/BkdIdi2nAy8H02wc/GMaxKmrDPfFM2zUUKPn
D8brYjg0nnoah/u0ExxKjowtYzDedZskcLMKRqSKCPDl4RRZ52ON++s+gEGMlwOQwLizi9H43KEQ
NqajHSGNxcYQoz6tA1WJZ+TDTzCeNbyf9YeT0kemg+naNlaSv25/l6Ob/yNDy07BpHpiX87Yw9HJ
Wb4reniE8Cy9abklAISR2vz4Y4wJpunKPaC73Rhdv49ZHrTCkr0Y+L/67c11Sdt7gW6oBK22T2yq
TXD7Sfdnq6CA3s3/bBVNpg3q7WpQMk0nlxe4G8/Hc02ltr7FNGjJJwiSF2Oft01igENf87vD08Yf
tUagJiTJpm4Ywhb8swJKwEks3Oikja/BpH4yO9tvMR6+bYpAU/PTyXWozb1CiI+GB0Ax46v8Tjg9
m048Ur9/JYx6YrBHtdnECc4l/G2CykgKSQ1mzjJCecviHAoc9JVNkH43zRv+sJZZyqPh/mlVAKo2
E6DOFLNTdH7cuqsCU5xRktPSF/xO1fN4Ve1lcTVc9llo5/3moRIpjXPRmlCNzF17/Q2ZZAyK9XLM
c7C2vy1328ItI6tEbDVXoQHTywuFbQ9Bb/eN8PSWDk8ZeZJoy9HXgaQcbr+mx2ItWPsBWR+oVM0H
AfzYV/UpbQxUH2OG0q7Em7qnU4xu5WnAd5pb3OTg3n1BVqXuWthscBJz4o6kKkVkTcFBcnJAM4Gl
4vkwQbv3zfVnW6YeZD+pE7J1oBNqaE0txCWLcmFCCd5L1F7BWeti3oH5HYMbRDHEgSoKAPO+vZNI
19tf7Tz/UTbGjkMNgfRpQmyjBt7PAmQAhyGjE7kgWBgVl+/QyKYTa0rKr7aLzfszDC/9rtyjlavB
sVxGGn1n88pFsO/wEAnSNZ0scYdo+bZy5ErfKpZixp0Rl7Tw1okTLR/77erqLPDolCBVTWHaZDlH
bZVs0OqnzEkNZTjs7YWafphRBzb0LVptuwxMWUVoGaahsnPK+Y0BK09HtD/gbaV6KstREIljUzhw
o1BBihX02DLXX2M/Nr3eeG7gUvuhFld7KKHRThqZ/madhcw0rfsRyZvfs5YPuyX4juMZgoYVtfdo
54IUr4ulYtlGwUe7zsHhj921tnv6JqXwbIZnRXCoi8lI8ZqqiYSjwg5YeHtAir/H1aCDiDrNnFnA
4f4gLWngxCYOad90QtNuyVANbTfX73EV46dg/W6OmEaLvcBdpKl2lZTTQayuarG1q3aLigNdIqQu
/c90ESUHPLIOfBetVfl8tyInhbJ3JmlJfWdAc45vDdvRw9Dcls7khdAZkcWkekcxlO4nLSbkWVkZ
X/rXqF9Yx8isVwUlvqLwKCn8UTMccYUqSQ0HHyJGzvEdlYnbgfEdEVea0yNlwHPMyWI3N/1yjXqF
B07Po7E+yxNIVu8k7377ZuVgT//WhZqzjrCWtlC2FTTW2NSEC32opAt8ecV/1XEIk3GLg5PAZPnv
noTnzN4XkEsfpuFyLAxUoHeX11rguF63ADKDvel0xJSZx7Q455G+0LGrd5c+FEiJ1f7r2BJKjpi9
KcK4rNZL3cA90rHVdAc5sQEafrLml/pK33UOknkoaVSTHnZBLYuU2eD8YUF7bDutjG0h+rU+xfQI
gWH659Ucxo/nfclZPHbdz3BGoU2AVxKXZD9b8erUdopOdrx44oCN8Lp31PAQpQ8D0f4M+ID4Y/Bo
yt/kk+ugbr8lo6wvzGl2jPFUafaeFOV/Y4DorH4hGQqO97xySRpZIeCsPtvk+DnnKCvjiXTYg8Kn
hlehMsxZS8tatmQ4k0rzI9+XljoSSr7Bo78gq4EhGUDPmQSZSXX3VArHEkDmuZFz79BJ/NC/4hGN
DXz37qpH93yyl9sHNfVpRFYIKkCRzAhoOOg91SrjcG+gMNrN9EIBQVVGWiTUFPWaT7xyLAWspaCj
Kn6u6U9LbvhdC7BTlElrbDUnF0JHQNhOwz5NVSCrWtGRNs/VrrKibXH9n8NL65AT5PeT4pkfGf+6
G3mt6mhiSAIaOFOvBsugHJzurvkwSZ2bfigo199XuQmG5dDmeQ4y7dpNmpU2nj5De68HlfgyZ66D
6rrDd4fynIj/BjGEyGM7figS+P1fwLm+3uzVuTAMyr3w7HZxIIQOKTtOrzVYcFb7/a56jkPavWox
rAbYTBoP8Uto2WsHPYtTt/V0nPAm4Ecg9YW8i6scPYmt4OaDq0xfhf+aock8AryG0x6BKc1zlZqP
Gebe26j4eQwyAfwQ0+Iqmxl3MT4GY8/OSMAbxnU51OkXSbXfe8oELeu2qmzIUecV4t2M46Wl2BwO
8p5YytjNvN0geImcOG3i7OlUucakMWuaOmz2m7p8Hv3i9RvkOziBLXCzKZJjcEyZC1CcSPchp54I
bOPy9OD7YJvhBHPc48Ym5QX+/JhDW25I6CciwiSZ9UqV2AjPmh+kZARfw2WakDSfF56fNRStl5GN
n52b+r+kpwYq6n1jqyjutdNiPOO5gWL2bld6eV2ei6DzZaVwFIlANSSOf1tJjanZaqfjV/+wnTpB
r9FJE7ln3YwrwPoFmGz6yq3lBo8jv6h6zg6UHnj3wD/7+k/rlbBTTQ4oeRrikgyIfrWLCx+rnd3a
NXt7faXIx8lxMTyylqqG7d0cijX7xEhLQ4j3yZZaKgLW9BapnxpP/ZssAWyejqKG91xOjCsWyvXM
hJrkF4c07u9bjBWj7FfikbYWwpLf+MDvbqquU/VWwWIfG1Cqs/jDHRlyVlkyMQWlqm76iL0NpGXX
TMh9WB5oZTMttHOm/xB6bXkyyKFAf3QRccoMfDLskVfjdPInQ3alA+QrZ3iqLxQrPc4aemRMqgs7
mTY5UHK5/z5nk1bg7B66rhYyxiZoX4WznL98pSuCFXM18TAQyaU5ahkxKMxtU35VeK29hdr+KlhF
QvPvbqcvEyrMtb2zaH2i6AYqtIGFhwpCHNx3l+ikpGBjfgDVpHKjCMQDo9UintG3e91dqrkconVB
HTU9wwfL07RLw6SIE01NKD58MKliDT6NgVilW0DA5aS4YwakWT6+KXpTfCN83gZX5/lgZa+T1hOF
GedIUElN9QJmg1ttgr/q7mw3r+4JL1m3DJYQ+l65YytvNLrc3Xxs1pPD67MeSMf5RDrNJCAtfH7d
AQ+6cIeOJpiMs7LbC3zYQBy61TQC5D8JOey4fqfXjsqJCSH2lGxCRFgEMLWQrhPKragQHfM0+MV+
M7R7LWjUq+bzPHaGDTlSOoIm9Ev9jaXSknI4eapTyHiSvVqRc+lm++oDSksf8MIFjqRa0y/IGbkY
cip+cyTWiUpbwozgH3WkniLxdWsbo1krDbppWrmDhalfq298maDBbC+oNpBILXDVzowLO3+SUcW8
f2FF6LBl0soFutQ0tfWkoBLYmCwKxXgMyU2Ue7V3aNl9WCSjKSo6VnlTT0/EIy36omwK0Zl15XG9
tf3F4HLrCEr6ZBq68L4n5ai1F2eS78aVejD/t/quq38ly7AJwmCCSx2+EA4Bqq9LbHXdy2/d3XJk
mySUClaZpOdnozBWUlZOrV9BfpBcg2XUxMNyWCU0OSZTWSdlF/wA+iyXg8izrU8rm5hxkcEg/7DJ
txbtW+UKbvYH268zFEiYEhBvVhLyb5oa6GOrogFcpHHJY82q+Kll5ZaPPkxC/hqG9rpZbM5gZOpK
YaRdCeWmaC6lJGNz0hq/aZ8ffpeulVX5jZLyUlQl4Zt/PW1AcNYIme+GJKnvcqnolK45HtmmjyPQ
5jlXXm+RlqpYASYSOkoUddztwTWE/gyoxmjPXF/PSBrKLGJ8xini2o3O1M/klI8hdticgGktZvJ8
JsJjHxi28cBzeaqAWPtmk6W/4HS1vZzBZDNFvLW4dye0PJRnWb9vYMIi4iOzlR6yj+zAng+jhr2F
mVb1DTn1HUjY+fndxaPe/sgrj4UCsed+fwMIf6mkt8OC2GJB2Rs+JGdzK8WiUxN7QQPUhdLry1hu
xn9de7SmgJnRr5oSmrGlOczqgN6kOzZ8obN8g5Emv/Ip1toHopq7flT2DZoHLh3N83Zueg0ZIf6g
NFLF65O69RPaVqXn6IKtTJqXMQeIXUP2rhfXJEaEJFSg730YSvR+mkv6S7VlYVAIxuqYxfx1YKpZ
9tZVMeijHdx8ZvfoL4zp8LJcKZxoPJUdnO4fdnEPsFsK/mKIhp4BGeAMb9jUimklyfG47SqALVS9
m1297MCfmyRFnvMvYT7ahKfgnsixr5XmHjZCEI0CZcerc7O33f0k/x8xzpWLatmrK2cwAmUSpwez
QvTIaRnVdkIkgq56f04ayOhYIKxZRAw79ZCrm2kUX4yvRjrebLG6iPpNornN1NT0MvEENQRXnBSr
MqXQykXDItWsNrOJE/dz4mcShr0/qvrXGc1+I0+Tj/shEvvCUNp5j9rWHYnmPNWIcfse308A8OIX
YZXhzoft/zxQ7dyAcNEl3lR6TIVpewkc0gfqCEwR4gdXG8bkVyd2iAfxLvpMNBq4TLehtQE1kF19
Irc1WlZPJYobPu95tFkrofSk5Kuu3Bn3glimsTsRApgT3JcMoaa3l/K+dNYUYzI0Ynpa1Rrf/IKP
zRi+lqJKwpbk71iQ7T5CWhL8jy+K7p7PX1mHQrJ6TPEXHs6ZXG3+TkvE8fFw37qXSsONYRTvyMYy
d6RCnHfbsmeCl2Vvjwb/9EeG5PZddnGUSJxoySwURzxzt2QjHrRKjhdLRIncaECdIn+9u8Tm5tur
kcS/ZPzyzk0exnT/Vicd8xlSGrB97dxVEGn0Ues0VqHoN93iWxUgxvEPSXBSGymGegZKzjlwykZY
ftJwDRrWKimFPG68SXbL4ypXl94oyFo728Swod+qtMvSPljhylkMO4CsTPfMJA99UX/1SlpZqw55
ZlgL00mn3SuBe22U0CFrWxRNsJpa9IcNioCVqay3QdFCcdPxuvodvHHZTVOLc7m+9NiDOYHgRNtd
Mxdz+ZMofwLOUySE1QtyNG+82r1gAlHNmsktDrTvtSmA+KI1OsjBqHA1tRcSY/2xxHuGEJaHgqud
khoP5SSvcdmWixxdTZT+ORehcJjcbRO499KgEcNt82UEC3DrUKHCuFkNuUdE7BolGP3XK4N4AnTe
zYr/3CjdxrPyDl20jPfjsCzFZY3qrXIerFOzWuRXRHpo840t6wdcNZs46bS3bn9A7B4pkSiAY8IR
4cj+JBvZkUNzvhvHK7TkxlvaCeMtlLbfhGzwiTGenf5uVY5z32mnrZN8Y744E5jVwQ8z8U1m0XEt
joaqmFC8iKgIVsgdRVkuYSIBGqB5tUMN+Hmsip4KrbEOpdK9utSzWFb+gLP/2XG5KACRj44FCOHz
5JiRgeTEYbkDloxr59KRtVedDGluf2vaQIzSgNP50KuypZxvJXzLVHDyV4vldK6kZ7xeFEzj1dVa
BuLN0j0o/VBEL4Mogvywf+uZMjwfL35eJLSoWu4RlARcGgLu25Nrp3TlIwk6bNlm27VIXKEXM896
56nRMJM8Ow9Re+qAa5w1cJX1+ust7I3iRzhynXnhL1J5gUI+Pfse1LpWf9LmsYe8CnmA/2TPec4k
fDCvs2XpMcUPpyscJPkmnagMJ62nxoP+AKoTL5hVsjM5qXoExQHIrxvVEtELqECm2qHWNFna1PZq
Hm+IXTJMUJxDigHJu5LyKXVxbwWASuec/hJ4neZRpkOWzkg4+quepcwmFanmbWmR20wDER6A8idK
vSnIdsCBve5g8r9zPdWVW1FXvyTVbhzlrBms+qJ6sq/2+7Q/HKv3zAQQgVkrwsjudeOB4wF/RlZH
EA2dggTUrX5PtjYJ632ebYYwtHHM6/aCfIsDL6SZhOtry1TENzjYdwdJI41wbBvGSut4zhRi3/Wj
TRsX2C3s9jVxeYKQeqpi0KrZfk7Ac30aCnpYDdbXlcuSvKWMQDT1dkBizaRsvigoDLxU6F3n/ktg
G/RuAN7UC5dpeb5zo3YBNSkOl/X2baPIdkxD2cQnyNUvDbeh0DjoHh1YT7xIhGNdzbD7SBRvtKdJ
RAZ/VSO/cDokWH1xODujmRGFgUccoa1Q0mN6SiNr4i1ADGd0iAmmIbFixDqkdQP+G3gnDpz3D3dI
rEqEj01ZJYl4uMq14uOCRe5Y8oOMAtpmK7h9CrrrDLHSnbN7X5NB2XGw07T3KX1ENHOBCg7ngk5c
9Mrb2qRbQaAILm7UeR4c6pn5/SKT+6mYtK/DN79KRzr4EeviphQzM1lxqQcoRRaNBGPt2y3/0b5j
jRztnKT9b0vo30gLbpeoc+H2u50D3AmfHE5deJZFwm/4FLEQ8CQGGKfi+Han7VhFFIZGJSAcsyga
Ax3yUi+kzxdCm4LMoYuhXcXW3FXvvifyXPHNksYTtOFRSREdPdzxYDMznoaP6tlhLWR5wsbupnRD
VwdqyMXrTrDYR+C5urgOxcTnBfLSGQg3C6k4mZPGzLfDgGLyCUEP9DwP+ma0TVsal9Wt1i/IExU1
VjmuA6lzwLOl+M4q7gjKjKgruF85YE0duNz4izqYM/6lRvErXo5+LHyOFkjdJfKixjTgUvsIaSm3
W7M7tNuB/AxiRja6hu5FXtYSpd6yHkscI96OkJQugrD6u4RtSrKCTqXF7jgi/H7OA843HF0iHRdV
qT9UBEtNI5dmnT/LE77yQri3PP12apYVaXzjMAYDeSdcJBI2ox+JVlhNGJwFxaHn7JhR8ZfYqD64
XQ36dU2gpo6SJbGSfw1xIGhicqbJ4sC0FtOSU+1nwMPhuDubLAc9ctyOj+OyOpEmnWrdjHoCbIZt
lUHNzOq1E2FBe4VoXID1ibdftoRBOskDNY9vufxXVnFmtjlnNn+gXo4CQ9eYb35ue8EL9orxlbzG
v8yIsUcd2oyXIfh7aLFJ6rgHJfQaCM97QI+AwMK6Plmg84OSE041V3JNltY42J9a7lYIatCbNDpV
BoUnt7DwI0WYyQuNC7IL9oYqdBDkU0icVSha+NXJZ4gLUchuP25KVq+MYYswXoSTh29of39iu6ov
uzJYNpvXxVdXbdZdC3k7D0lT9sZJhul2HtvVS58u0Q8WS2YQwghNRRohTw+i4YXgPtBXVMw0GeUa
friQI8KK54Z2wxjIQZ03Yz8oYpEQoZgW/8XefSCm1T0fo5iAppIoGU7abfrA08M2Rr5pcbPOF868
7TdPmtZ0bXolgmQEQ8+9PSDNEQ6QyXQCgoi5cz/knXTQgVDnviZcc1LfNHJYNMOa3ez5mqz0PdTa
1Re788dVC4Fioa0pHnQgTfC179WxzgCINcEK8sp0VN6vSVczgVFXIUwytoMoZDX8COXW5qDVuX8/
UCPBXg5Les8ZNB0cIWeZX6cePiVqG1dJNKmMj3VpXTviHg3x4zW40zOO3E8JN/5uaoVFS1SLt+bm
XUizM76XhtkyrzmdSDdbWTWd5oMSx3/yVjPp1BCDq8GaDsIQoFfR/z6cMSFUt0DL5OL0Peg0i1tj
KIJp1dmojhVhiVDAToDogQI2kdm1zW+gMz5u6N5RUqS5Dzlp0HzEHv6TAzQkgxXQ1peT6MaEqap1
WNYLDLtREWbYnuhJ8H4v61NyAl1PNOqhIf0k08ODIHT6GcC+Jta+JpyrM/ouivFqt88Zq4oU50sc
gXEqaRM4fQNLisIFCKmdvJJIEZEiSYzvHq2vJRzFwDWPWxop3hWRILtCJsIra4JpTux1ZkOKIDEr
27mqxnrQy2J1v/2UQupCG2LItprro0QwYuUSdfTYS5TurmMcxp9/0Tx4btp5IUNFTzZQt3FBvooJ
s9E88NZB4OsFf72IGP9btrJ2N0vaMqTXV+J3VYjO0d25M4Bxcr4YA7iKkpCpoRkhPcNyp1qh4GlL
8f0KhndhHE+7FfSvOZhtG7lHcuPD9rFb0i7iI5dN2nEnd/V32j7B2t+nBzmNUmZS4erA5ZqpToUh
+zvbc21BBRZxByCEUOyVw4Dx09SHMK8DJ/NHNxAaOLqkD6scu+ZnBxWKXxookrceb2BlhnEO4kg8
a9eMQCERG82BmIswr2BlNxpLtuDU+Uysl/c6AR/oS/+FQfCu9lPbvow9XSJhJL4mc2e3a6fproLN
IBRfFQuF3/aPGI0oVp6Et/iZadPIBGhN4R2JkR6ncHBSZaE3NABH4Qj/q2UX7Lvq835uZ/ZKnpxj
/1f+EP3XUx8Hnf5NVymg7j1UkbL2U6J4r19sN2ilCLSRYYI5375Fk+1Hdyxd9uNVELY760W/KwGV
Qr3Bbwi3Bv6gHTZDL9xm40OJPaF0CNS/SI3g4Mm9VFSWgQWM5YZBMjLtNJGIJCjN7TNdhjP9J/Rw
Q7X7+9sJJKRnWshki/xZvBurtglvPvGFJxe42t1Z+nYJmWK0N0QrKXiZ6Z3belK7PU9nQgwXv5Wj
mfXg7UOUCfFzApxmX7V0eC+rp/Wl9dFKipG+Dt8rTWTH/Ot3CxFs9enIsTS8ZPajuFyIucJsYYOZ
YbrAftJc5HTnf1evtCyjxpw229nhEiY7DLecIorVwRDau0MKgknF2Vd6V/Hs6BvqWlsvaaQlXT5b
icgK2q0O6jXoO440j9ytsoKOWUsTS3vZjQRLSD7UTjDN50PgdLC8bYAsRx+ckQ0bTK+jTeABN8G2
jlpcxa15Q1sygLp8BLO+wXeku21VuXMxdZrnA9slLK7/mK8QlYv87hLpXgQofL/c30oubYoDb6Je
GNmY1OVDhNJqz6MkRFAuYF4lYhvTIOdbP1x/G9bZQLJZp+c3uhAG7zcRaKC2ZPmBmdVGggPz2tGZ
SOCjpYdS3hGyFe91g7Y+HJdaRkW+QYWYeanWyr5cQFEC0XsvZJRfGwTxzW3EeFdpfEtpZtdkf0G3
2zGJqnmEU/OdIV9MXBDorsOJupDOqBjfEljfHwu3oam5kDIW9KhbIOZal2+to2v/T/uyMbSD1jqa
X6Lnfkgc0ZpbX5V9OiR/7M+q/hnTHyth4t4P60to0SVNdmogkCC3ij4u4GwRV+lsOtdWfglYbtGl
zNzxwpZakSYg2Vf3clCriSBmdXKZeP8gkaAjb01PGm+SgLcXNqZNunpDvo4OQ6q9gPmO2hZupUvX
USUXPFvQp21Z/FVlrfHX0arvQyN734srvFZW6TCks0wQsLCNxkNGOtAeqaZHkmQVbxhLovYcs6QE
QtnRwkvQPzMH/QMZEg9G4pbkvIGXF8XLG1MhMYErqiVxpbe0A0D9ol/ZVH5xGVkA+SJxhDrnd2g9
9aXIV4LLtpPxwxC4KvrPWZNa//5mzVIM+5H+cKMHdYNtOPab+pItubkL1Yn7M4AV98h3eyFdePWy
4WYaQpljDidOvwO0ZEKLxrDtNC2HJr3qPK3Y/AzovkgdsEO5+wZaPfhgBBmVbSkjpBbY4zLPbPjK
QQF89pwGZkH6GZh0a0qm8bobHNKfkr1P5hAchfN6oo1ZZmwU85bRXpPDPT7e0RiogYbdLd0bggWo
kzdGzr3sRFSrfNw1Vs2sttf0dclmu76rEu908oahD3mZP6tMVcSoWyDklY8c9VjxD/jFNAEA6feD
66BW9XYmqIEprdeDNur4s631vFsx+dGB8EtMkyxPIcJdGZvOHWFxlU6NLxQUxB03IBjYcnRPLEQr
ui1FeugEwn1h1QYg94+ihpb/JdUqUpHvLZEBHLgsgrEI0gck3ew6Pnu9t8qqiu6vFshYfaYGQAzd
BwUJOlpg3xxrzf9ipALYcnA1oKbOzeAq0DYt4Bg1Ou/HvsipGZWmVAw7US2vcHgVvXxbIZdN7hrC
Glc8zzhTO+PKsVRPuSid9nqE1bjtAPHN1Vhs2R/IcsUpUG3mfzC05Km56PYLWMDtNcsmpNlIYH6I
aYv4OqSzEVEanN3vGD2ioSTtMKusPNED8dB8bYlGaHsYetjiH+23gt3dVyUotH9f3dRSP2xzV1dM
jj6M3S/u8ILJkMF0cDEW+SrM4nGNeMfJtCOZ7lFbZykNobN6sOqY5JBeYhJ1nMEKjvswHAgeXaRh
3xjEng396CgeZWDSlgNuCfd9bMIlEVz1kkEcv4G57t0q9UoZ6pKOjIh3PiF3viYY1Voe671VGysc
4kQs3kPwCHzVxvFdQ5kl4PhIAq+06Jo3Zj3siQN+7DNXN1X4eR+uhJ2ZHqq7bp2rEoYCCI+7MHFe
3Tm1lyj1vqRRccFHI/ZqcpoullX+t88tKPs3BlkLzmgNE89eQ+9yTWrMvhKpQ7086Xh/dn+qdp1c
MLazCdl29Kl01YBI/bDI4sAjOlEuy7l8KU4fR3Bo/ckQ0ufmEGJzttNQansChsvHmjmSRYY0d4z3
AGI1HnLW1UbBZ/14HbVjep2aVj63MUTEan2q688UYbEvNm6s5dDR1nOd+TZoJp0eY8pGTYnpIq/J
BYwrHz9pStKgtBGdmhBHh0WGRt//OC9fO1yW4lmzDp1jCds2Qvqwm1vhIVPcJKyLtRwqKdiuq6wM
fQPd6hBvlvl4xk/yg1SEYhpPdEdmjy4G19TbOWb4bHl5cboblH8/i6jw0tTuwINAVU36/csb44TK
sU2tkdygeiDVmbG4IOyyLxOvo+2+DCjKGXOdn7nrxL6vzmsn34GsI3GXqW+L40HzInUWE71ehVQc
DMgmsfC3ClXxIJdQwZu5FJsWo//nlr/+ARTPrfr8g3Gn0mbEzmWYQjXK9okRC/kDhCG6i7QaLJyf
+4mM5qQUqnq8WFG24zEbJTML4SVwXexJAHOj8lFQSEZBuxKQmMtbJRlRZo54dELp8nemA/5dRyiN
EzH7Lm4CvhV1MUjpnz+zkip90tzKZepTQiTHyH7nkXVipsQAyh3sZ02hS7g+sFMPe0dp3pCS346O
ptU1geNz4IL4gFPp5qG05xmXe+yOrGLM/6EyZKx4T+AlOswqOqjRgi4368KBeSG29fz3jYn88C5B
9sYuQ9dv/LrtjpZXevUHgUmEr8miH0arTcAD1DhDcW9k0YOFDfgR5KRDfNc8wUq51P5kCnVrCJuk
6kZYTnTHTWcManLmc3EdXJCkqPlDoDzHUU7ZPTWyOcsZ7k7OU6oVqR+iGhl8k1uN6jB0jOwlPbaE
k50iB3Z9pmntAle4kykkOnhYDlTFRFwV4cMjc7fymTTWrXGLej+Niqz9Vv7CMO4dgYRX+uL2Nx5X
uF9eGp9oHD03ZLN0yZ5qbakXHTDkdJ3KDMbYgEZP8MIJexchAuu5kyIY7r+/Zo9zMvYTTzJh4H+k
ZDr6/NfNGD+SvcU/3NMPQGPNIQG+p+6gz0fBUlWxa26tE+sLSirFnq02nKkey2hzDlGrxdHW5AYW
T8xQBlIJM+ZxhrXfwg6Vu/14Ks41fT3kkGePPQQI+0Hvcs0VvEqibcqFrwaAwTusPkvWl85Vy3Q5
/GJuD1J73xQWQtRU1G7GR84jkPzfy/q68Mg2m7gujVi7HGjbJH0PlK/kxX4jkVCVNgjD863ywvhL
S9G2CPK8qPlwFUbaZHnc++RpIG4cTzcesSRhE0QuG+uKuU9ucaFkd+j6rGEI2I0e8UN6mnMzQ1xp
WGamS4lq085giSUWCOLvfP9V4Kg515lin6LmosKFxAZ+dfuTGygvgqaxK9Wz9cJidXwEusK56Dpp
5ohHs6zk5n1IHjktSmiixlYQIXOCyF8+SV6pVoHkUSBAfpyIaeHaJ10tPlDhvJdUE7duz2HEXeWo
VQ+vevjdLali6R+IDScvcFD95CFadlN8pQdwEAcnzw+0ofmxdPo3OBv9DaIFSKGl5NsCVmdS3A40
Tkntf1jRQi4mEWKTfl1bk5UXWbr9Teent4Oi5wkP3q78HTegSbXAKbueG3xHzzX37qdc4auA1MAJ
rg09uUqd+3Q77GtVEbLPK/4AUpBshJccvS7A9Tb9RKlADnAnvvIeF/VbBhSFPyIzDOVb0Fbp1+Nz
G15EYMgIxjx+eDhzZzg0Ruy9RFbzTOOHLnZ+2tzMCzBMUxApBffeWH/SH4grkhN9Vr/ek372HwNS
HiilRDnI5wH5eFLbRbh2nTrQHWLzlJ1ZRmnI03ijYIB45SScDnkxVlZmcPCDQg0zA0wRqzWExJc/
K7EUYFsKySDukqqiiuVPC6fWOI6hglYuWen4KuTztwtpzXYNmPWSWymJnywcuXgIH7nhx08qU7z4
49/VvelmMtZc1SaokpBYWb6VhEuMSHMJEUv3TlbJUnmn5Zn7RM2BMAidfduK4hbXoqgT+1u+G/VM
Lkj7ckdC4SAdApqWA5oUSrTd8AU2pqCwMC5qha6jhpTdbJsqRkVajuixSnN52bj4m7AjTJYEOBaZ
lE7d12rr+KJwINJaxzg5cmRT0zf4XM1jQzqf09mofx6oSfpdQzU48gaybdgCLnKUjpilcVmJsuAI
O7PJfNjVG/NErmXYUrVFhjB0AE6c9wLt3zJ6T7DydttjNayCc3GVPv4sAqtm86dxZFDSYIcP4SXP
ggR52OAz9eBjCADIIGfd8iptTjwIsLeh1CZ87QLRl/O9DRMfg927fR246cSBnGqt7rVSJqU2EvP6
F6fHxK9PyFxTH3itF8yl19AglBABlh86xPThCh24ZbZ6eJiv7PVMF6dXaYfiwdV5oY1wKg2p1OOE
eoBTXsw7sz6SJ9vKh916LQq7n/KtXryQF9Wtl5AIHJJw3mhBjUYmWmrjMbRgLvJ+v3LAQQu/wJC1
DskLTvhnyN6wLPwG9WQlAEG2b4JbKHmccrz5RF4k/PnafBXDO7J3bRyBSZBo1bu3hjxqd2W9ow2B
M4JRK/kEiS6sgEaffEFttNCj788pvxB+RZoJ2yPoPRvoWuUwY67pddIrkduQSIW0bPekpoYWgzbg
LGjXpd0skTqkRUgy8aqafzm9O1LLUZw0nZvmt+l3pdTI0JaAZMKAsTfODmJhcRi+jDeJu7cAck+B
XewSzpzGsuKrH7uEU2Jh9H+ig2gFmpM16u+YaT3C39PYZwqe7il8gDy9AvmV8srj3OddwOxef8Fr
5FRNJnUWZ6uS5z/fUHk8GSFNVtvbBqgQ0xj/ILJJpcJhuqGuPi3eYtXaeL5B+MADbJwSmLMShI8k
xGaxZ/FjK5HVTF4NuNMS0dzH7tWpYvFV3YWh1s9PfoZZuX7PEaSyCY5wp9YsfFkqrzkSwQzR7wbz
qiFHyQTJgjImOQNrxcv+I6H8u9TqUo1aqZ/V3DoQZAsT6LkJLL/12Rb23kOnNTlv28YJ0hSc0lQ3
JRke3JXy363V4zP3lTIlYxHh94P5VctrDxwYH24RT0ZZN75X30XsRpaUJmulUttX3hVBe0Uotox3
OVNut1uReAVsIRcXGIlsVwCx8rUR70k7RcOMP13x7E5wvOPTlKVl+PNkFfvVM752mMGVymDH1DYY
WxvYOzjtn6rZNkBIWh13V5gipLb0O49t0dkkNXPp148oaevrXtzzZAEo1TEaQfYn6iVeNCCPrSTE
qAVHUyfZajWGLp2AHwoEaB+NYY/hipc0v5LFtSEG2xzVBnYmgUUe0vG/dbXd+yM1E0kTgJ3sR/7p
btIE8lEC/evqhlspWTFo33wWDeyNqOh9VdqkOt9q/tnODOV//qEepQE8mGQ5jFDpi7w3dJZ9oKXo
siwpD+Iq6M4XAfIH343hSh7RwN5AJuonbHdJuQWrah8FZoj4u5ILO05SQr8fTPQNoAvmoKdzcPFh
vsYVlTVR5yITvw5Z9WlSZL4sGvZstV28mjcPwY+ULtTE8IX7L9bf+vPMfZMOj5NWf1zikqumGQLL
nKL2elwqKuIZxQYKnm2EjzBgxwM9ZTZVn53fnpgAwT1uVxQQMkm+U/mSCb4ah5ih2jTFKbilx2Sq
MTQjw5vhgtZ6ex9njeoYqF4Y6TCXUvdo1GQB2naL5Za4Zb9M3HMHOY6ZQyrahnh3gkG6I3IssJf6
PoSWp5aMeDcFdaDsVSjPGAGs/KYlhUHicdT8EgnYhYQsMHDZfx39L6hbmALPItxkShJ6HsXVeD+f
ARPLVilfeX7lxOr4yAHczhPOU0DJlbTXqcPWOL1IV3Isj5OYUU64UecqHSr1IP5S7EycYvA0STqV
HKitIGImKIuRKtsy7+4Cz6fcBivl15nmfdTOONmby91vBzCPnKWFOOSlG/t9Xl/1LJITeKyc5J/L
xmD8bFEXUahMP4vkpWftUW06deIYAKDjbgyeFWlTp1TR7IWsS2+Pl7Xz6nTTkGeEjwEF1VcHnKcM
1pFe3+ENTzHWO7R259zDtJDnyAqLAtveHrIUwK3O29rDymtyEiIt6bqzVNs9LAaRCRTUj+I7jCK6
5mZhnazZzgP7inmEf5ain39Zq8+K93TGtFVbaCmb5iQIDnZj5VRauwyGqgFN1EmjCuR4BkjPLwUl
QjGc9/OIdmsXR1TrijMGsdyxFSAiMfafwevCm69wkSEkyAiXMA9Wz+uyI9j8x6ET3ZYFvzZ/Oe6c
rgQ7NwdnaBbHsVeTVmz220vU3Q755KB93KJhAXn8eoR0THeSgTvgfKVtQ4GeNkPKszNU5gA5LoFw
uLzMdU9bWDm/Fb4QkC0/apFGR4r180Fsd7LgBLvuCxkgPKmxqi8b/SwGP4R+T2VtI2T65vGIT54U
mpWovmiEv9oRGKAUowFGqcGSO/7pozaUwTHWlFJwmQAYY9gqda8MUroTmkGYLOwOjewQao9tg9+S
VWyVXeQLpbWqTMRY2V4FdrnDZFZA26Lapv9a2heKkCe/TVK+v40Ds7geiZ2gvXlyty41IqoY6dM2
3lniboPpv34Lfx2abxTNqJxE6mkHceRjMoX1V2XsM2OScYqCZ5xeC6mDkogPRp5Cg6zhrTsPOokU
ydOGQL57bGtkibpWJYeWsJu7OjH5C4x3ULQ5zEvPTquHhl2DXi4KFHiac6a0u0FmfsB0YFjy2X0r
JCcdbwKwFs8BWBK9dBpJY2Bf5ARz8Q4GhKFyOYtEON0NuII3g6O9Db3T3ysAGAB+w+Fv9X/Id5NQ
w7sMtVY/KrAiord72CxljoCwYh4XD6kMJGrLkV9N29aIpTEH2I8DTQB6gLzlsncqgbcSCaYKjZpe
ToE1mjlXIDDwKrdZtaCjdfki4bTp8AaSmiZ/kZKbcLVCpyxxyarF0x8dsHPCYJ0AbpPydEABKf2j
Q1Db3aCfvoN5UmnxRGtv/dxnuWqGucydFnbm0wYZjYk8jJtoq6V8kJzzWwvo6sTFvYUCjpaA6Dc0
ur30ZVxhYGNRGaVFEuRZqonG48awJf3ShNX3mZAxN/x/q3VNVQinaDlYjmNR5yRdTSxXikAt46kz
dsHn6ND2VxKuLNrm3SLH3A2nZDkKJkqSn/RU7KzOh2Rxa7un2Z+g8/6hYx0RuMY9A6Ta/co1WmV8
lAbpZy9DOx33nBqnzjYvkwJiQGzgep24sp49xYdWK0znTtRGbf1TOJD+jM3+oiRyU94EdCnuitS3
3cW35FpsEikiMAkjQbK/1b/ZuqrBzzyc52WRbkzOJ9pKlE0/hLSidilQvsib2WqYDzehwBiXdRd+
DWHZwkniLjmE1ByAD47usl8XmuopV8wydZauPzkkLCY0EfkC/2EmxCnNSrGQ2YaPil53Bx7obwHs
nMvESh+voxUZVPzY2YMexo90UZXDdK196EuZxCo8M1qpUeN1/mMEIikfUZbMVlbFGpcJxE3etJ1M
MVRw4uXY3OL1PPGMbxktXLTc6B7ghzVX0IvmndzxibHtWuoNN5hfiandbbN7jMfufMTq+Y5hNE8i
0ZVKhuf8HEi9AnJOd7YLJhIJNpIugDMZwj1aGYFgKZxDolChXB13CIRq/XCx9qMu+sJgnfZW5vEq
E+XkqC9c6SLxw30KLil+jQbTpMAaWs0526v6lcvBpmwFVHxlvztcr7fmnRmJ+PT8MHJ2s5xbKzqw
cQQS1vi8vUIcGAei0bBtH1XojeX1cxgy2DudaGK6ZKllnKmjgH6DkJDlJos+Ze1cQMd7z+61q6W8
ZDRF0oDGdUrNpwGzCMwdrk0UH0T6q3zmGRlTOdjE8CaQIzH8O2tmgqanw3zJ42bu7Vsx4BNBjSbn
QSu8kD2NInT+Lya1hg80dEH0mzWn+7s1HcwceJk0bwTaya1paxqUPSrZeryvdqWSPOun4pw5V3kf
xD5fY1kiHsHBMmyUgjsb9Up9s+mqvSs1l9vClZ4Bkr6TIwJsQicAkVYzoIUdiTaYu1i88m+CEdXO
8BLd+Aa5t8QwYmY65wQ7YTJrVY13T0x9QNq2IiQXAQtzPBPCLHAdzskXYxSrLyNaXoL8eSF5nDQQ
m73ZOxjptmO0miRb5KmHdAPKYZU9a1obSINiueAV/LPjRcEf9dABPr0eery4lmlfKquB+H/ISQU7
4xkslQD/vitJxfk9rUDgGJibPYOSW38N73zqfnRTekkdL8DZYgmxq/5vwmfuWuU1DlBM1FXz68Os
9jjf0R/yN6Nkhway1lchcXlE2L42NWcp6UqCzC5Q5id61SrrW45JapKUtitxIOQ6KTqt3c5J6Xb8
mttFxbTxqFFB6mEl1At5KpVbqzryn9KWW0MPdPaqaneeEe9kIEEGIV3zcj03vsT3OYvwh5J0W0z9
FCYvfnf6V0dBBlCxoOZJmC5PCzJL3v43lY5Z/ALJjJa/2JPVNazrGyRnFM6bXxgvYU+9PMBpYRbB
r9nU3qwWGSFUM5WpFA76uscPfk7s64Uijj4kPJYc9wbJWyJlwHX3HQejF6yg+96auyOpI4WIp3u7
sJAIUZp00z7TWCne5z2aSOhzF0oG8ZmmcGbarlzaOYnJCnzMSQ/GGQP6//guMlnhUy5Ps8MQIJ9X
oJusEuhpyMFuLhsVjY6D8SnNUB1XMz/hcsU8fngJXuTeJbRtuzwoavwNUgp3eO2l0xCUbcWOPD2A
I/Vdi4OfYC1POw4xjgvtofOWaGrd0xmIRS7GJSbltVEW/pqqKx2Hj/txwy+8tlAhMLOlU5d/VVge
AlvjyguvJWcRu2l1ppAgsoqdzNSAkrUhMIoByjD1KUND9E5UIHUK0OmxB2f3wvkfOZOcOozwEzw/
Z4vohWP+rKdOulst+spn4xHT9NnV76AsIvkwT8TjIZE+9zQ870J+sNH21nu3ezk4KV0hnlOrqBvC
ZLG9OhKkL6eT+YDU1K7kk046CLPh8L/EAIGVtRVEuuaU4sS2RlnJZplblxCsi+KYUoKyjE/pfcOu
Y2QQDxSacAxOJuylPJZ5u4eIWIDSD/I2zUWURXy9byJHq8YbPSof7s9mPt4rRdzTNLRvHCz0NJg8
DipLkU26RiNAtlOq+SDQxSnGHx673HkCPsTAOrVITOcn/eJT4C3XPEjodgvOUc+dRuBCOXHZryBv
OY6bxiLR577pQyvQ+/k5TQaH3EC/6ufDWA/+WpKJluQhUtBbMcxWmxG2YI2xZRWHB3akdFb/E7Te
OHYwfuEnwBCxlB7Aq/gd0o8zp9FHwDdQDV9fyRkydt+KBKapJVk2MWbCGBOZQCtyRC6Z4hny5k9+
Nu4Ub8FoD1vropM3K/HuzYF4Rqez3S0FSGI30tH2p0juBxGBbfoGfPlm21KCluLPUr2/iuFCA1sB
SMKWNcJ3s94Srn4+FE9lcJNxXtiQ5OWNlX/FEATj/2rZhXEG3tu281SX1Yj4Imvs+YkWFLAxns+T
X/OIp98nrT0jEF1+pv/xiMN47yCr+GR3Vf0i3qRmNwyHuWN3K1c7hSnaHuY1pL6VC8YHRmj0Tq4W
JbW9ZkLSpo4lZgL7XlRofjmjv+G9DNK9eDLiIJzb8NV2LIz97E7rPN7kgEJHEyNPW40LOUf0xTJa
3u6Uc5AsO4JL0Hceiu2ibUnLyLgNyyhNZBoqkAnV5AAE+kcOIWLXOl+z/ffTrJBi8bbOvuoIr3dN
FV9w5n+FR6vIUTEVdg8l1xkWe0ENavIKXFTc0QQnb42YYt1ulJEmQogVw87Q+bRZx5u8gjY3wW+I
qaoxoNCOsjG6VPyUWjNPh9vgpm1o8N4WXfEPm8ptfgfbhXoV3svOCoSL0dp8sEwfA82FoLSvIm2m
VOKbtVwqPcBwAXCF8wOJClc9Mn8Lb0CX0+2ZSq2uyDn3bGj951K569jfM+G/1+ELxKEGLAcEjwsI
VODe6vP68rZwLkyz5XAu/W6NriTG4ZUgvEdGAkfw6/tMJuv0qHwofmT4+YK1UtqKFhJfXlM0pR/w
Q8f2Ot546BE7ACha6UtlACehNNUZ/MivISxVh/lJfg+trHdUtlvOZHxvWyucGqIrdU2p/gPl0xiC
b6jCPYiOB5MshaS63f5vKuyo8e6doZqDmn6w64ivkoZMvesJuzSnB1YF+wb9tB8Uzlfl1siwODQG
2KbAEsXuI2Z68OQGRdDD8QWQqYF6++D0pO2EXx7LfIsKl9nL7Aus2gEW0YMGSAJFB5xn5S/AwYnX
ct6+hcSP6O0W4k5nPw72Wu9fHU54S3I0Jn033p1DQZwu316vMJ/8bT3wBSxesid9rrRTCgCh08bP
HW2Mf5Kmo+pcg6jKT6p/sR0+4FBEGqcjJGAGNoL4jsjJ99CklJm3avMOqegdY3nptUUeysDR0B3e
RP91y4T7BjfaJj961QpLhAvebS/JlFHKlfiCBd0IBezZe3go57k1ZB3W5YKYu+V77N9KfZgZuY3j
Xh/bzJRVtJSb39xyBqK87kpUO3nsYhnAwNCATaui+8CDnPRZtTeIbiszIvgFW3IzsogSN7HPQLJG
97oaqpeed/j5g6USJEBh7dZOOrY8RZHF7D2xO3Lo2mM3iP7hKEhRR6J77ZR/61O6+Ubyc3yK5Gwr
vNsmz81oPcRfnPltaF1Xv5wmJQ55H3yYKX3765KUwFSZQFCF7INab6An3cRPUcmVI35HAugEh6Nf
CkkvnS9BWUufGMdrqUgyenzciFG5f/5Sm6qjzpD7zCWfkN/XKr1KHHkM1PPwwfR8K8/H5uWUanIB
WbOOWQLjYE6XY9llqTC8rEky19aYAckfuOIHCYSZoXr1b2/PVFgD+3IpEgV1zAeJSqwkAnS/b+Vn
YTZwTRNUaWEfB0doSpkLicvMkwLI4MhxIH1X+TLdIyyJsEEtaEL7/53VtrjrQjqLlUd1ALb+aCzz
w1tsHpZGZsTX36EQCoHfSvEpMSUgs+1aE9MpiupjioiJDJY6ZaDZv8rrwLgXhWgoFHQivxz8VloT
PkqoXKAO4nHz5bsSySTShnPeQJx6tCMg//qfTbq3agH6TAsKSuZsVhVvOTMu95kDAjXtWJw1l0Px
LUFBCzinBR07b5ZDhBL+KbnHV4GtNLIGcjZBegadgu/N3+Wv4ICgUarmwZ+2zzbq2rgIu1T9Oxa0
KCiT0c7YfgVdeUbxGxS0xQQ+77xy12LG2/pJMCGui2FzlJCG+5jRuRYZ1e3KosJEX1tQ3fJZ1Ucx
6ujGAY2RxBtkXwuD84bnx7VriywctDSlLG8BePVByapOnxfTfKezxmyoJFuZwskLR+W8vsSarREd
dBZJpO1ZJ20rvP/LhAs8Tq+rJR5Nrt0TTa/CR2fFMyeQ7YdlVDk+TxcQZGf390UIRRrRtp9KcfTC
KTKOKqlkMCllNt1ruf6RSLm8zhxZrshVgfYEaOsTQZb4uX7vqC56VgT9FZZeORdKClMozyRPtse4
hjDZHvYytkjES3Lg2uBDI7OjBaGqMm9Re8SE3yAJ02ZgBv3fPXQ+c0NeMJmm/DqfwZBfYXC+LVzL
j5GtC6bXB2fiOHDDo7F+Wj1F5sbiOYoVyRS7/Pfk7NI8Xt70olWqAlpnblWE54AjwVsEtainYoCr
8aKRfujwv/rS5+GdSPcnJk/ivGf4Gz3MIetw8IQESoR1to3oMBqJR78PMWRSY0T3JBm/Aa5xvClb
/KpP37GDNtefVAZJ75V3QkFxc0++rpglVqjetA+zBNxa90v757jDwcqx89knMFnBQ+iyF7ThcGCo
NGfp/p3phdHVeToOLe3dbW4SM4/QuYOUIZvjhwtOQsurI9ZlFkXc0ZHBSG2R4dqqnC/4iVuFcFl6
AKzkRi/s/L+taEIxdrcw4wS+KYKU0yEISrM2zSVA8Bq3qw81H2IqJ2CnJvFrY/5GgcXz0SG6ghSo
LdaW7fHlsLDLzw7xDCZhIrLvP98Zu1EmVKgdZ5SfTy1bju3S6HNo6nHGuV4sUj07LdMU8Tk6Yehw
IE8cYZBYt6gGGboM54Ei0yYBn8Sjc0ucnWOurXM32Cgwl1vP3JguWGy0hDJxw9IJI9Pj/AGypCrO
v1tzlA9sw++4RxVBMDzFe/XOxYthL8wpa8n3oxxDTmeqyoexEio/AzPBDE+OUM8KFInnKeX0QrFM
+QjKd/hMG2lhFOHug0MsingsvX31S/NMx1ACNT5XU49O8OJWwCvzgONy72LyJRh456zmR2xchg8G
GPI6G2y6uOv3WiVfQpX+iacgeIhshdVcZVVB7Fd7ulEqePKG01rc7i6XMeGjbSNp2mJ7/E+mk5x9
GxNxRRc5peeI0+XE5ZLxR+ggHryfbktzQ3Afo3+DsPxHlZh15UPS73v6qDp5BPRPrrHKTUIfmY6w
fdqH1JJ58CkjpZIYeZjL1+dMhAukc0hAtl4wFS6B9XoCrlpCNuqOyVTgytJN2XWyNnmkzg9hfSH2
TQn9JGAt7UBlw0zTWciuOLtfTLOgUt09Cat3ejsYfBXjs/3N0Juihww0RH2cB9X+eC989yloF9wk
Y+Y2bLKU/QLNzmEc+nzts773lx8on7+SEDARdW4+znR1MZSeNW2DtKBQsMny3HtXT+P5ACP1Fezp
2SEPn1NieEaemPJNV3q9ZOCLhjusZ4f+AyuqIYOXnz0OCjBeXhF6ZHwDB5WB7088UJkRnqYACalM
Venvn9txmlt9I7VHyBIy4OaaAVWoz/hucS0lKPlrCrCfjvWi2dKsYnl+gyqVrmlbbTANPvn3Iz0y
XcyoIqDr72zStaT/b3yht6jT8Yi0OS+a/HnZqOzmRwOmeI4YzGlYoUpnlEMOpJWmoP/p4iFJJfu7
FbvSqhIeqVFI6jrjBveOP2ot1QToPRLBGHtAnX89m3HIQbJlMuyLtwiRZzbV0zcDHdkwtjm31Reu
FKyT7hlIH/Hx72w84MiIMBjhTlyYpCisCfVFm8YzpkJc/pCeHxkiOWbKKg5svrgbznpIAMNCvKHQ
SSIbZcoZUipPF35k+C3kQtZmAxcTX3YwObFXhHDdfdjEHnlQAKTZWUaXgIIAKhwKLjBZ76OSUZWn
6gwRKbR3WvWa7POX6aG9cpKT9Xf73FI/17bzwp4d+ewcPihw0p4SWjRLxAy41i1sKuqRmZfpY22U
PLMaz7bq+/mw5VSnESzXCLyQeTswsGBbgCe4eWrwdjnPepHBi2hfbqJ7TeLKPXhkMmCHk+HmomJV
jymyAUNo6TOXJ4YzS3ZvKQW8BTAGUq1EliM4CoK4yQzxCMY8ma6/Klifkx4tniN6qfswYRx2IFaV
oM9e0qnDVfLWbWqylIyGD+j9YzjiPmc6MVx9sXExEIWA8vR8VdUG/2eVtK1b/KKwwU3Qw8yZauoD
LZ7fJIjS1VyswF2PB6Wj0g/oM0GrkzK/DWvutob6Q9/aYguHdqil8V6YuZeKURofET6o/BMyS70J
epEEHTQrLUBT+OPGB3XTr4tmuEkbIMJLqed44in8O91kDVM63LNmxkf7xoQWVBYuBhEgysz3SVfN
sHeNCQgAGTxk/fpzsJNrNYt7bvr9hU5O7DQ1JQFqJGyePV3r+JTKXyiOmZ75zepY8lJfubz4vLg5
SV+8A4s/Ts+XBXWP6L/5VDyIRj6THSG2aDTyRGn21RPByIpjbz4b9KX23XAHrzw78JfXS01vEoIO
SKVrBhqpHohSyacQ84H56yqRVic120Q6DpWyqDZCL+DC8BETs2NjFRKCHKmfsfZaagXhV4aCOB63
seodaAyGrji6N2L3AW/2xL7SJcHIYqQOsIHE45F/TIsl5bJwg98D736I6tw8aKwHgrRNxf35oNbU
7ak4yCofb3br+irWdiA4jEq5pU1dRLg51PcwzRm9qqqdbDaXFDhmybar3BVAd5ZMMrpULM2OLAjN
K+OSKOdzvfXBJaUFL5I74MqJv9YIYkiAa7GE9LBi6TnF6w0vYiG3bioB8r4P1hdDF7+qn/RDum1y
9Xo4ymGNxcoLiiKwUqooaSNNcspWao9lw15zIf/I+vw7KrvmQfro4OA8nd5RUk/fnUzEa3x5NYU6
gGKbnt8yEibbKkayeUI43e0E0cCv9ojgTUf1RDka+bUsVu82Cd9CE0/e39JW73+A79Pf7K4HsqC+
E+NP/cTx9Tv1w3zRYMjJsj0erDuMwRQOrTDwhlCJgv2+4SYg1wMmegDFpHLoVfKbgDMp4TLaKjuk
mZDTrhXAgqIohNP1viaqOyUHq9qzqmQq125JYTVBT5/DY86gNTVtVxSWP+HcqRQjT8P8hng5LZM1
mBDVfPMt8L1RFnihYPYVKn74MMwIfittzA7MnDShTK8zWChCtA0Rq/vAW19PNA78MvNuQpVK5Iap
QXVIrKOy+wBDKHmZznWuR7BK0zmERX8zcEjBJVjd2dr3+0Ab8WhGutbo5McI3wi7LFGzxh8i+CLv
abA2CYG+hlzkkojifZAkxLiKczsVo9YO7eS3r1Pozxg24B7LhaAKubJnVOx52ZnB8aCe67Mmzz7O
Iy9rh++nJK2syJsIckOPjwyoHoYWaA2u222UusDlBG0Ranm+lJBEYFGmqH4mxzl0ceYSyqGQ8lur
942J6jEtp10p796Ra4ZiqtWSuiEH5Veqbw5msaM5Nh91kXhlBAitMGGHA5pohRRKwwQDGt9L4jaE
uhRHO+eBsSIRZxRj8o1vAdtfw7UxeOZ1uOBoLw3pyt+axi94cJnJyfheqKyKB7J1QtgFtCkd5ne/
WA/BquZcA9xYQqFiOnNt8sLEpmM/ZQAvdZrGY+AzOyTCmAsKm4yvm1Zctz3GPrMTat27n9xVFdI3
4IvM7/m0dKJAci8eHMqPgGVAg9s8midBs5VQgxFTTHOz6N32IBSTThAoB7jk+KBX2EvqeQjDCfNN
j8a14Po0d53oNZm+6xex1l6qTOMaQqyhZhLNk01u7Vp3CU5EK5449IRq7tuFsPz3Z0W01IoJ+kYK
j/mAfEdoAZT9jR8Vg9j/aS37Exzdpj6BwXzocGsVEFPp3UMc9IksNcqCGMnUhgSXOey6jGxUxF8H
f+poXueLIMlKS2Jsa1xIaD0uZA7U1vcIcSjum7rd4hUur0ivhytqbdUQw2Cv7jvj5sKmelpDeA/7
WAU831xphqgZ3XcVvp1dYxiBjqvrK09icEB8XrZ1kkvaKqCKffT0RFUzKeojH2kjrcuhbpfbLw67
53EpHmno38mgOgcrk+myyfabThTjcRhiGIDZTrf4S9WCPFJdiwFI0ezSmf0kOWGRuVXc279bUkbV
LRDwSs1gpIx42RBGYknFFPP+rIeszvIikUB8OGWSBuloijBm7v7JCTRcMSfB0jTtStV/ioc88tQs
zCaZxx7sbtTp5kCiCieKZ3Sbt9UUSqt+cVl/DCma6C3htw6iqV0wvS9d8atx1YxLCtq06Tw+EKlA
CFAy9/kBkinLrVaPboipz5p/Nmwqzq20+Qvfyk2hgWmO0YaMPUMfsPtSd2ZzNiOf+gGLzUuD4bpD
78jmz+3HHs1cBPMX2u/MPkmZyaslxjciQkbHTEJTUaQJcBo5kFim9UEjL7rHPYaKKr98pgsS4gxr
uFByRLalWh65Dey/Ho83ar3b2GlCw4ZRIx86uiiU0OuVp51/4lRrIq7EybJ+c/2Gt+ZSdLBNi4cD
nRB92MJN53G4b2BQk6uqmf4+i/JZXl3ZLNdNk4SpNX48PnDc9SSXW/kHNXWGrcuEGSVdB61618rK
PxDEsbvJzwk//xKNB3EVu/bfx6h6ZzeaX/mONHMrCax8ji5u2m4tNz66Kx/xwhkTGYTUFd/aFyE7
9CrleYk6mg2pXTxgBnOekPH0no7WImW0AN1UVEvazt2rOFki/dIWX/ix4y6qZR7cj1+IQwBar9cM
SC4hwf+tTkqBBUBSwHZUQER6bcbXnEkNonrclSsa0PyVN+ftrLT1VxuKjp+uAE6TTxEH8aP9rvof
T2A7rTMqBby0dtZ3ZVp9ZcHArKIWVAEJhVfeIY+IUe2faxmIYqI+08na2rz+DpMVbVwGaNID7fyT
ry3jpJiBe2Pw5HgxPcy7R/Vo/yZHvG1RgpaUiIKJq+d1tqpJi394YPagC3B+P5H2aueumx3GOiOU
SU6Rkm0xlADb2tCUmcXp8zQMzFkm6bZa5XTnp9LojgvB2WAkFETFmO+J6XJtiQfmyJf3hBE34xY4
ll0e5gjD4vLXGmdmduFxdc7wrIcE/7bK6X5K4ASUGs0wgPSBWahTfbG9JcZ+YwZbaWyg2TG7rBku
0w+IPtm/+Bebb/SENSDBFXXMIQw1zQY7G94hNAwqershciiejd88CzKKPw3vqLiVvfioa8qnhpup
pt16Os3rlHoOePfc5AxTe1zfYoiME5anXWDhaq2ynK7m1g1Z+2/f1eKoiQsDD+EtQgFmNDw1NyDb
2H/7mrqflcPvAiFYN0uKtxohe8EWNEwpLvKSCwMmlOS33ypsr+U1h4WG8UOMIeZaMG1XKo03qdv8
PAu4Q6Z3/m3SNso4vu/9mEC/6JEDEFDvZcGbipEjVcjdZrLtLpMn98T1KpJolpGEE5HHZ1efA4ou
J9us6cMTKtuWd+xnE9YZ0tYa3AScfFdguu19SyJLzK7/F6d21OJm+TdjwuSsUqtts/HK3Up3VSSr
DzgOcPvVc1glSY+8jV9nyFpGDXdmf9ZsTHkPvQo5f0f3nmE7zooZq10/UlY0ZVzpYaXIBVzeInBJ
skKYSwqsrtV7075mRZVLFCRkvG/r9CMgw/QlUHF3Nv5ioOwmfK7meF6+1vEtsDQn1DOgrhInFOKr
q13W66RpOrpmFM+yDlcMNc1oEWIGBVsUNV/w3+BBJsy/X/DDbIoDfK9XX3dQ8bFW5TLVe21h51xh
/oh8ANDJgScxTHYz7pt2VNPJux7kuPYeuHtZVKzDRC7HgrDr+ITYaC0YexjQiM7SUyQhLYJUabiS
3lplTDQEnd1U1BM1Ekf1C+iTYJw+gaOQ9w57asQarPOE44EOsrwskPdy4cNRYcdoWlT/rVcVo6n1
gYCIJlN+m57lMfKeBZH2E00NAidBifTPdaE4Xf+YwO1V7e/1MJ10Hyp94vU9JjTgqAZumL64ywmL
NNBU+ZvOccVtKexJMuciCWlYPZPWtT6mC8UY0kRqqhqL/Mm1NFp5HdSPsO4hSN6py8iCFrf5Ff5r
eFgjh9RSKBamqoNNOxf2vb9WaXm0fzsQ4b1y85tVaLVGLKj9mHtHXAiR+e5xDtOBNka85IB+Oapz
v3jxODyfkBtP/EcEmOZW+998l+X8uN5UFvlPuGlbuxjDZTumrx3CN2sNv8Vm8ejYrf9IYTwmtgaW
TYHaxlxb+dcbwBClUqy15dvQDf5tsO/kUHd+tuafyo7JpIu2+1nkLSOoPJ7zlVju3ifDtjaM9iwu
gXv9cR/jJZx+J+CEDNL6w7PfTYeKoHGUvq8UUmiVTPPoTgUnUlbCDbtIj2WGfO54JqwBAOwBhchM
OgN+4oZBxcpR/En7jilr0G/0q1IQ7SAzim9ZU2HeNyyb3WJFrciQ1FHu87PBcVlVNUWrH98ohgE4
Fdoi+c/ExzqUexojZat1AchodbD6xLMZ4EgnlhgvF/KKZQB60Ygtb4zyQtC4oq6VZlp8GManRe6I
OMl29ZRd1hkHm+oqq4GzyG4LmvLe1FxCz8iOtUdJPEg3/l3r8AOLp4VIAqD4ob/KklCIhilsQlPa
8/H7JkEMmjQ926CPqTNgwp+RJUpwYWptp4EaPd4Zi11TXGz+2FZBnEIQ1eOla5wftgKpJd+qNpEA
4TFM/KnsddYRk30sVOr9YgNtrEnh1DTKxNQtThEgcI+Vk08XF2XqKXFOhjjeTZeaaKOqAq2yz1h/
OskbezcpBN01juseF5KVE0zEvo2fhoChAAkinvUXdR/jJ/hWT+8k1YQXHTaX47ENy0nlvPrDYbyJ
9OS5Yb9MUqPKi5r5JCrm0gGlNac76m1qEgm0OGzx0TGkQyJZI6LFaLAHyfMITb6c48O9ZOAApFP3
Mm20cAKjI7tBYAN+keRvNIKjkAEz8XYxULPSyrJ3JSKpaPsx+oUYOY/UeaQbom3C31sXWLfLgILJ
6M/8YQWRmLC2pz9lvdEoiFMHn5MFUnAzZHZX76ufhb8c/HJ/QtyQq13vtmlUlSZLqoWENpW8Y54e
Q0spE5eRABbxcY7OjzBHwlktzCajLJlEdbb3t11HHZJqmyTczVB5QEpqxzpilrIJji+I6vc9YegP
Z4qrizt4hLap7u8TGhwrxb4hwh5VMQ71vMIDDQ9OfRirSUzaN39d+GGk6+9I/vLNTh+ieBAKwMoa
ad5kwO+oWi9VKOnjmE5T26cGuclUnTz/ow07W9PWXp3NHSsVO0//EL8l/vG/6JlHuAQSiGBVk10R
0WVVcne+yNB7puQSvpqM4JS9lSWldRJcWjaok+W6ZMzO5yQQ8//GEEbr/SeRu2BZX3NVd8qV7y1C
xBIzyiOi1vd5FTWzSNyJ0WRAEyFywh+4ZvKIKk/cfSOTnxmMnlWk1c8uHb2g+3po5cfJBGaq3YXM
47JiADyFi8fqXnSK49nA6KYxnyRubrZWiZRpbwVH2U5akXLd3FoEA6cwd24Lxv/vMXt4ng/IT0st
+7snaVoa6fJZ5l7AMfbY/BpdGz8gl/txIwdnJu5SUzlqEYIajz/gwasEu5ZF+xJwLxM4I8cKrHQW
ute71XAtpH3A8TOhkErvbKdyc5mEPiSgPjvh+hDkgf9nDwJTzymfBxF9cNjIt/US+R0znJ9mnlOU
OH/wJZqyVb6TOJNjZ6fqIByj43k1AVLvXSzuJDZDbIoCe2k8eb6hj8Q1w898vww5T5jAVFPpkmij
mP4cUt9wk+eTvYBY4pmLYqSGEWdzL+DQoutlNuN8NfMHmHe8xdNrbuRaTRc47DyDzUMMxjCYv2me
qavlCBQB94FoOIY+BC+/kGs1HARxI1OCfcFE/n/P9hxtMy6KPxZsGRCgNxh2355OPyIX2kZj9HjO
2/NwR8KogPw8mkjTRAFPxUqkcpHYsF3e/MWQzIW/KMTmMhdlWSVGlF1HSXcUNtP1lfCVY/6WVdKu
RS4Ppnnpe9AUeNhq+IlXtO0LTcI9PKpa/UzHfh4Mpk2Gx5Lk0O0C1WFTO9xVM2QlPJECv1M3++Z+
G7cXZ0cYfm9jdYMeOuC4VhNrkPNqqm6HL7ZUU4aW/n4mOtN02MMb1ttkidy0wJ3Xf47YwQnRwoYd
myKvL4xqj9D4mKjvLeOwsu3qAktkXcle0EHmfPpCjxr7IMRaIIQbFKVfoxsesA01tPJGTDXdZ+Fl
91CQ+1VWIq2LAu2MxyUoVFiA0sX+zp6p4J83cn+A5RQPQCSO/K33lqw6qas6dirrqCkP8XWvJ4Pe
5nzVT2z4WrRlHNbUyPSlIxLrwO2dDFmulIDr0XFhRthcUdJEr0ORGHni0Ug8mOOrITaq4Gz5QDd1
5x5O9bnS24Gj9yJmyc9r44wLy0NPGQyKrEAs+tSSsAmRHy04DwQkwy3U+w0sRaJPF5WjlZkDLCSt
sxQDy8tjzXsnLUa/80hB7Q1Eiql57UmEfWND/X7BPqzETXk8FxOOYuoz+HwI8Z2G57xVibMgWwFN
5kI4lCZJQog/DJ9RzDpaQP4fNxLqTTKmlEGP4xFMwDBZr6rnLXSiKOX+PhLzi1kH9td/mZLPERpM
W2CBjp8AQKGWU4wlvqLKl1YeFwNk9n/Nqu+XrgdFcF0AeDIGhEM4B9GgEdzIqJl7pW/NmDzEL7/L
31ojz1G+M7DprwnxQv+1zAys9oiArl5knR5CNZZsxhAm+SLcD6ssIJDWJuty1ZqrpFGTmPZpijGg
Or0VevPG1KUW341LF+1LCtLBnwR6EN0W81atz4s3p5lULCSkLx0ZbPLnm+gTZIV9XuTLLI0qoLp4
TfND+4j8CmlP4n/5RPNL3ZGwPcyS9GxLxwjZrEQSTz5qoFtSsGbUFYUVe6bephrwlIhTxsoIapII
xrQlpYSqsDUHknkiOn1tf4zXew1GJ6OJUQMLJbtdNBwfZDP/NgH7TywXxfC7GU4Kc2g3FNeOazkv
cRR8kQq63+njd8keXQEzQHrqTQG2Wy5HtmIYJjcR47w8J0thXV6bHaKxc0TgBIJBBU3Es7ln6keG
/aK/vgKtCp5b9lOplJfU0Iwqm4yhH6dwL5A/Tmps8csnX8VNiCLAY/3esTsovDP9zVVnpOvrwFv+
bHV24e3gxz2oZ6qksrXWQI0CD9/gLOuUgrxwyiVy1wCPuTRKGQkwllW6Mo+a/141IYk5M7i8e690
Gqj/7+saV1OoG+XfagV+t4tFE4mHer5tpJNPfDjPGFEjlcdfKBBZSt51t1CQ28PZ9lnhZdWh+3Wp
0pqtMJcuwHCFGQKU2o7X6LqUS71PtGPMNTGhmItAgNrOm/FCAnBdE7K15+MObr+/XmJu5vWsKH0I
d2z5IA2I5k0DPMOCYlT4HLVdLQdEkPC1neeXIVgysBMK/1iNwhYctSIDCwHHXz4RO1VerORJwWpf
CJKFuOkWVOy/Jn3li0Uj4ykD/h8fRmthLm779c7gS/XaPT2imBo1Sr1GNWwqWhObJcgmW8JachV8
ZQiXgmVIbPo6yBoCTbt6z8Ark1YoqEvL2bvHOZWEFQ20P010AfrU0QkELX5h4hLdZzD3PscSnTMV
SxDaH8iHSTZZ3af8ywzqxtJvDpGLCWvMGVSB59xJuM6oWjfgzN4z60VwIrVJqy65OZzSe3BOBAbR
nONUt4p1GnuIeEZIwnYivgQR3Ukpet2fJoobfHEbpBp4TgAALm0neSkfiPbnFRkUl1YVOZM6nqM5
zNH1gAdawj/+vV915fM8yrkRfBGlLhHcvPK5nr8FHXzYPJR4z+UNDGwmlOzLY5WSMQzr5fwGimWd
DlX3UEQeb6WoSqXWKHQqUvkwY34bIYYaSx6FqfJTQLtGk1bv61gn/sASU95r0eeyVb5KdaU/Un4M
yF323rXcXeF6wsVnoAWNAvuMUr2YUnNoZcelsaPeaIui1pGlAVAe3VlOfdPCDnlLQcTODsmWm0nH
SHdMrfPQQQv/Lc1bzmFfi3pFdTVc936Ozay6Nw2fWaaxXXrhpEfXnBXxcad3bvmuzIznPAW3MUAt
JOoOS21kcHKLBxorjb7GfeQxoYrRtFKug8MFqidGN1Ry+MQc/9Gw4GgrZbxgn0U5dlaeTbkbgBtp
4Ov5omgFU1rLb5h0wXgymMxSrhyr+HP/CDJPSvbjKhHCrX/xovq9iZ7Iv7Ten19sFfkjm04TiBtl
MM2RVPdIg7Votvq9iwNxrGg7LVSskODb1UqtXFPgdcadYK9jDur55R/HBKSN2BFKdGybULkUrViA
DDnmX43umbpcqySYdk08VrjTfm420D7Xardc96OMba77OWW0cGxNiDZtPArTSAM7hZmYVwa7gFi6
DmdUgDdgq35qIoJcobg9chh/NenKBoLw5rRSu/rqhDv4xXp+QFERua+EefUDPfofeownRDLOuOKt
gmmL0tLY64qKwHAktcyLqPsqs4MH6YMVWqvrxQcQdy95H6eHoLZnlLa1hTUOD5cz3tVYzfGicT+6
t90UBbD4EsGPuCdbaqq2K3S4vbPXeAhAufR2dbHLgiTt11AFEgsUVjwN7+UN/P9DgUG4mZYsuPX+
FuW3v0yhEB2F453Q1xnou5B3Q151A9S4ibDgphgFAWiOVHs10SXwVM8PSpcwO+ENBgyfnuqRuntt
uuHEwOx84IDMWOACO5y1aDttGSE/aNwws/kj4lsuBXbTWCRjgUmyxcLz9bZmni4fd1S/R1KGVHdp
/AHoFA586J9rbeuBVrMtkNYrwOVwI/1TZ0KSyEgdMk5v+YCNqqPE+lDe+ei3Re5e5ThV+taqLfGn
Hrbk0p2UWqmojdAMFJmIcHKuEeaNUdr7SiXTnY7JCN8b4IH0x++RLnEbfmp6VbXAaxtJ/7rWZqhm
9HLcTTWuNwBR0gn/gGZyNFkRNwGyn7C/io4wqAL0NY5JIIX8Lbc7YXqVXzJh1ofQJheO7NOePTNf
VEr2bZmICImBpH37+pp2ox/wBGiRC655iKnbR3eV8xmOsUf/VmAvHNt0lRs65EjYWHh7JDAKsRPW
YNNXx8k7zBbCFk9SH1cFmrmi5QI0iijOHk07UoEr45lsLxxoIJOsBlNkHlpx/eu5c/WFveHACM1x
xmHsmL/IIuSC0BMiE0KgwGpZ8ZeQJXpfque8KPmr5b5g5HjNC/uLnvRwvKIdcA+/AULRc1TWEpMf
NpF2sDHD7Fh1W+a4VCmk4SSr7OewELLUlAi/MtCsG1ZkVeCiNUTDwwNWTgPptWszafXxfWrZdn8a
5ufX26EkltRO5+qxP1OcF9khb6Y4CMqIkNSVyHJ5T5IDfK7TbINhZQo86YM6g0ePygE75WjwTcVb
qiGtCe7TAWHZss0ebwFAl/hnaTaHWTjnLnS2EwU26HKgc8lca500T7jGoorEvam/rquUiKUjUCHr
DHAqa0s+zbA9roXVUgIvbPjo2q/CHAfhQ3pfHhe2vcDjVaCsCTGX5lJpty+7JJrkNCOlM3gdN4xw
TkDxOWBWGXA4hnzzsksvsoaqShXzC6sROhITfZMQE5FgIWR7iMr0pydaNr8TgxIWhJ8uDDmGIWCU
ALb/bC45131yqrD+5LjGKS1yyinAv8XloingNloWSduCQyVkjxFaA9vGFJ6gNNIHXzscuqIN7Vhv
9czauaOT/3tv0dSRMZC86XTn9Rz9NTcvlQvTe6Vkuz2DchfLV4LE19zA57hH4ezqG7r+fh/uhtHy
SHF2FFB0Bh1T6/ZcfDW0MTMnIqc3UltsJG+kJ/46zdbPw0SMzEZCssszcxlHM0B37EIq+lhKIK7v
xlxs6T1dRFkDeX1HyH0hRrU+oCgtTS9iGQ/qfJQmKXkPh64IjxIcKeRSTj3+RccQlBtC24Sdkfym
hhbbEwrKCZVwtnv2QcuFteUe9s5+egCTo7grzvLMy+JLxDQJHg5yPSRxHlpdCTW4/fg2CRIBNt5T
w8hW045pUhU8Rvd5Ac7ozylUOds5zZYQ6XoAIa3InMIQbBWHgPevj3YWPoI05rkLqJGDyzR1pZQ4
JMbNE2m2CFzC2xJV0OwmbQCH2YQvlxNLcWKlwJmS6tvM753GIvHYYC/mxJUWvaTzZ59507D+75Og
/z+cdFZLcwVxrzpSM9R0qWGBrkfYTO4RGb40SynPK0bCnwKSooqKoBBsIo+2LhCr2/YwarTlnTNu
7eYYBw5MSDFUJFsYWRwnKtywQpb+o0VdtUm5CpkbMh/ICYiwqhnr6/FXIcH/bqowlqGMfEee9lwC
n/i31xqnUe8be50plaUluUe9nV5F9GrDZH/YecD5MsHx+lWq+U3J64y7L8y1tGmrTQuhP4UniR4T
YcsFOr9av8t0dvewkx26kUet0hg2gNZ9LPKo4lZSfxzWW8r1Y7GPA3OEd7fy8sE9BPAr7YrqvXFd
YVcqrjyxQ5a1oK2KvLUMU4TiB9g3RsvzDUQDYHENns9FOglGuvVfqOkQrlxtVDkx9ZzGTLcLlB8y
OBR5XOOeop33PGtSenOfvAVhPFjZmwLXP4dOHQ4NPa7tAtTp/u1S7xYVZRDX90sEDYjf670dzPR0
km6j1Y1zTkUZ6BqQGEkR0IyLupKcsZk02qW3LUn8UlSZ5vPkYqa/9XX2J8Q/kr+hNZ5c72Su0UNp
PCKzDVhKVaz2VpD3CddaCc2Yh3lQ/cajvQnQUczRDxnzSkyG+n+QX+d5KobMgcupr1TZCoDYlHn0
mPJJuGUECMlneL62sqpeg/VR3UFKfM8jkKM2Bd8dJsYJXJ8btE+pzlk/bHSOmdv5q89ypUmJVZJC
v4JjbhHN+0QjJKdm3uNg2/E+LTUb9wAcP2MUwcJPfEyBczccipkwJItVA837Tjzf0aADrgUR5ph4
aVoBywKmlXSGyomWkYjDePk9Rb4UI0AxiBVvF25DMk4P4WneW9dKjNB31Xv/MJ2GOBNesmKRESA4
77R7M6Ycx6FUIhHelwx72UHapqy1mOAhXYMLgdczXy2mbz4YSFBvFIq33YwGMqbbtAmOO1H28Gw9
6Vu0pjE333O8+GnAixgIyA8yVAAhbXgGtzWc09PjkfTFew+ru0bSQc1hHJy0z5HX2Rq19mhOq4f9
ZuunQcCRnS/4pxN2T5yv715I47vZYhZNoNdTXR7J/0SDvBHQhkVs4+Al/TMCbH97T3eJ31HaUc/x
T3ewEml1M7X7zvJRTmBDSyBON0RUCnHiySlfUeLwl6Kgy+VmCntm09CykfFLbiyTP+vxeYLFtYqA
9HDnLe2PY5phenp9dc9SeD+cTCo4CLRmefMQKMPifye9yJ11badt20afRZxDe+MfhxjqvVUq1Zc+
ZgZXCW53kfN8rEvr0pACewPIxQ3T5Kwa3wVGM3wt/2bC+w1yKLe9tAsLAXQMXKQHYi26FXNfowd7
deKX3TfK6xmNpPKGBXwcM52y6myOuBeNxaz4UchXNxY7J0EgloEFSF1PiYN1oVUgp5ljX7+A/gpy
iH2GWqQuv4/w9ku4IVpe/0jp3vozrIewBEPZNj2pqs1N7YhAtgrIjwy8gWa8L72pj3GVC3jFW6iw
wclFULBieuEGJZO+c0Zrw8TQZQH50AUf++OIH1ozhjNruQV4WuPsBc3TRKMb4vyvvl+wsdhPbuC2
Qun9Jjs4OuvIDmgUSV/awZzv50LZZcDwgydmUvWEsWCtfDHBSj3fx8VFZc+BcNwUVqeThO9L90me
RS+thlpbU99EAq/do9wUqzRJ0/xy/VOuhR5O7NyNfXgxmKfBxL+Ew9ZQ5d8H5kiIIrh7nLD/g9An
fKgQe9wkDY4k7rNf+bOxEC4uB1o9ZQ3dCDQRqha8zn4HzElUCP0DvrHDnA5NjTmUhy6O5fES54TT
S/Tr98Q3XCvI5lDMQwTMvuMG2iZc1FC/B7EMsFaVeDooUMfu2wvUSSt7v3bGGj7Zd45s8QANy/ml
18fTlyhVbT4JwDVvGGqtN9KzungeRJm+pDL11zh5ZoARq+hwWPISg7fMykq887o9yE72jrUKVtsm
ptWawUpV9XXy15Bu0VXTtaBI7eM2rjHEjCpF8ZCs4+7kGloFvwTbaWxj0RgW4UHkfTm7qGrHx7HP
27BcmfixppNzsBQhOZFDoCIyJYlI5ZeVloNJzm6nSb0tlE5nwFX3y7BNnpAYGhghwztCaUmFmxpY
UMZvgOlkFn8IsLiiXt6WZFD0H783ojMpcTbBhocliZYNREGWPlE/XsapXVnbZrmsaU2JZZTHu12D
YbOTC/AuzoEv4sjkzPqymGe3+ONvy2ScizTIHR8wTu46f/NFT3wXgrVuQlR3XwB8Wvm5N05iZPPu
nKGOKZUxb/WCPZGcJO2pHEZmrGBKQQRTORdvR1BxYqX8UJah15r6IB4VxI0zNE9LUUDP4922t7f/
tgN58zGU2a6oUD5EYWOrRY7OXj1GfuZpp3pEVme19UExZSzOws7bxDTZbyxNo9/zfHNLV8vTuPhY
RUNpgGpTP/Wj0qy6qsVyZwl6jyL9cQVcJtl5bypCk9XfKUu55/0f1CcRCUn/k/H0Y70olZSHkOTZ
EyJ5ClmtPxRRHF/GomryOkXPm2X/HgfXYcZAtTCqxPSAoVTFQ2SB6mhYgvNB1ZYWg1mDzBu3fKUD
3D8nkwuGgYgQz+EAlDVNcPAck4y8Rz5grDO3X0UhCoe0bGukhwF8j15xMVTKuycaQLf6gr2fQJq7
1K6lubCM165EpNWoMIUB7HwDPbNythbc5EJiA/0FeLh4hFV7h3ETpdBu0uBdKD355PqYAyFcVckh
P45OjU9leP6EBxTbyoP3NfezjvsfqqnUmk6vy8ykO2FZpZ9Ud8SAq8bLUSXl+0aRlZFzTDvh5r6Q
/IqMzMWYEV4CXtPtHFRrJoA2pWJtDAhH1BEJgFn5i/QZk89Xtq0QyUNDusyfM3swBzkKEfMPOBq4
+ojED+qdqvh4xGmOwfRSWW65Vd256zDXA0xvq7DW59QDtce9Yrmg3/EcupxqHD/1oCATaZnQARDg
rAwD/cPpyZWEQANSXlYJRgZNfpS7kcfBLTHIyhgvnpWgR2IBR1vPGs0zfN2utAbMWMywfddzIMqx
lPlfM3UF/XZxDOJ+eUnNYAY/xOTcRpySXJYx6mTx7uQCuEFuh9rkPaT+LJMaFdNJKSZ4cvW+0Jct
VZsL3nd7RM250buoBdNZQ75wN+7ea5JFC8TOxxlLfELL2UdnR3YyRWt/2tQmth+d0kzbwf0NkJVS
PGlq1a6YcZVC5iDeUcArgHYd25Kjtkvg44q5PIh8fsw9eLD7zVHahM6mMvjH3tuvbIQ2obX2+M6M
12RR963Ovl9Ksabi+gvX0l5UsSko5RHZGoYwTxDKFxYgN5KjL+pTOuFIAhDE2kkIjUbr8lX/83ID
n5m3ReVHHuu9zIjrlE8XqenBqOS3HZd6bHEVpS0uTOVnOXyVXXBr8Tgtq1QAXaqdxjlbtFmZ9+Ii
5C4nHYOFmiypZT207/7D8dZaGxUyt/NejZWIqwXMtvM1mAUpVrMw06X3Jcj8rdrpT9GRaj2NvXg8
+ErQe7re32zfFbyGvExvi4OCZEga7CweTcjPwvt5gjFVooz34tns2AQtQWBdZe+nePzZGIQ6HahX
xOfmK8i77XkuzK35u7Z3gpnzUDwb4TH8jm5sH2NuVMqV4aSrsDoAC7C8QhINv2I++/BymYzOaW9W
8yKupbOKuyg8n3X8fj3PlSHKGPBRJ5HDitjF+349Zi6hI44Jc4lQfHSt7wTqbDlSkjwirEg0aQCv
2TgVOpKas4klI3SMWNcOrtXh4+N2AQBHduQ08lKsAqaGaCpf068KQgEReWlhFZFYfFxpQjDtApNM
mS/2VkX1ACdqV1wVFzNVf85NK6erKehSnTGx+FZxS++ycP1TD7KrPnXTxKq1B6rr8MyG1i63osFL
SiJMSiq6wOqj5wFF7hZ9gKti8BJvLyrNosNNRjJr/5IbSFuCW4wwJkQ7eIjCillSUyEJSMi8cgJj
KeKexNRhaTMKfRv3CIMOgduDPht9yCAO8KfSAY1iWyPra4kJka/4ZfM6RC+FigMaeNpH+ZGcjjvB
hLCQ4Cd14sa+IRD2fgt9v7rhoVtRyvd0+iwFWpRLyYsb+ZfSZl0ZNVn0MG5MfIl5Czeal6Queesi
lwqvxLKjX5uVstCheShP6wt55b96/XaAlgt0RkDcVfXfVS/RtYxmlYrLTugfWCgayfxhCrZ7Nmh4
Inbf3TjZOZqf3rYCdOLSwzxA0MUp2C2/ZLi1ug2jQTOoqBaM5lU0YZiGr58vZfQ8zl3IyeNvQSi4
/wndf44QJ7VQh6LdZeuYBZ+bYRErWvBaNnvveE9CDbAntHrac6/UV8f6pM4M/6jMQ94brI1M+nyY
tRmMIHI0WtP51SGbYv1/VRKrBKfAQz8qKEmRe/F8QDv4/+Y+3+fmfK2JEt82HWYXbBBsMqVH2ucq
DfWOZChxJvOyt94vaCW5LqrQGNm90De58BHqWrEjhuGC1vwHbC9mHKyULlKO8bx8yEpS1U46xTgk
61MbXIeHv6PAcKfls1eQNNGkeYvEDUWQJ5TBgGwE0DMia8qUGmc9xkxEYomWgRRiCrf5PgDU6B+X
mtmGHPecbMvFw8TaySWGJ9kQLapCRgzS4sRI4tlZllH53O+uz3GZ2BEvA/IMcCW86Qx2c7PfNvRW
WrisGp7O4kSgwtaZMAE/16F92glIQb3PZmKCc/+VlU6KAa3+2mZzSw4Usrb6cJEs1xMoanRaAfms
DGAngeL5gy8Pg3l7TX563xvrsRnpK6E1xYC3d1NeZtUEnMDHjJhlWDPOJij5QcX1KSSF0/mHtlU0
k9UdGfquTvKBcsJASSQ9nXTx3whMWG2B88G86ePas0gZDe1WZhZ6IkyU9NWFGfgHnyowQO5apaKA
04ZLCqDZQzIkv0ZlBGa72U+Td47bjzx5cSg1q4x9GXWnjVnQ9vS+nLxK3PQ5E8XX+59KllQiZy/o
+3rFSohARsnnMIesqHwLdFNqadcKdUaatGWd9FUZSlq7l5vvjsCqdgix7C4JokafMIOo2rGHGT+l
60iOk54B/bM8s0Q7ZM+TVQ0G4fMiwzWOH55MNbdVTpCzFZW4ZUqSIpAt4rvP6hsyWrppkS//os/j
CAQifXbvsov8RRefwWl1hbcgr3SFwtcE8sUY8WEznugS83pkp8q3sCIMbup3uv9A30S6iEtPED3V
RXwndDLwRZci4fXRDPy8Tnk5rEAbPV03T9yqzj59GJ7unkGb9yXm7PCG34CTUOigBpBQ4vPCk8iq
HlW2lT61PcXZjEBuGgklDLmTRdGpY0Gq7SnZRJuZJURBQHsk+PeqfLDEuTskuaVDz/yxIUzawlu2
4FTFleFeBhB62c328Wmf+S5wDCOJC6f2gpBY8Pid8+Ma9njqiy3s6VF9oSkL09HJ9vt3AiH5zInV
Hdp2U90OnoKIs7WN6A8YEArPPoi/oVk2q5vJtf3n9Jmsgdngl+VY71XSATav79RHZ8OAMaQ1+2LS
2dEp0DI1BZO/F/QSTqBOSVd8c8XYvzmAtszV81VXsAhXhOvF6RMArFiKmh7P27/H8UeTRD06bKqe
r8dhyAJPR2j5EHForbEiH00BzRbGqIthK5yMwRwpZuj0uwDhRm/SyROl3uwy1LCLXwlyxmBOyWVM
GxgDDoTp3YnIJARgo+m1VPRQIJ4jRveSI3L5YObf+L3AIpcyOQnw1bgK8v3N5tv2aAjNxnlZAba1
rwkng+v6qEWzpGoYDPrID72Yv4hxyDuwf/s7XnEYZ4WdA1ztKfBbGXZ+0KhTy4ysfzYaC85/uWe+
55IN6eyWIiFqBynk9fsn7CFvjOku1TtlXcI4V9pmQJX8mqr+CRNiD1qIU12eUT0dF1uV2FnfgySj
isJ3/ll1o+ZyPfB+rmq4szOtG4zXq97AY3wc4Jq/y+0mtck9Fyfpzzp4RI7uxkLEv9gvGXKXQYPo
svwuY9NP3waEvsqjNcwmfrfbP/ydq/dxF0I9LLAaqwg4ddanNMb30dq6YY3YKonaR1JJU/Z+kqb6
GkZIxYeRNEreHnzgfgRMsoEv+wIXYJLEBCLwp9jml4vbb40CqBqsfxIKjBLjPY1wL/M11FvQjrEY
din3hwPWpsEQhTXUnG/2WQOs/4vNl5mjsra3gCpMy0RNEktDFm3zxjJ5l8h5tRRE4lU/P2r4GrfE
XnU0LkdDgxc/puIy8LuNO8VcHKgl/EnhOjcfB1PoC55270b3focz4vb2MqdL/xActavJI/j63Qs7
s6g6S/TxjPF0yaOYy3eFVaT0Buh27Ba297CHbsMpDpKmEHhOwqwYE5+txs5G7eakSltRbM6xKlUp
8ch6K31GRN+ydzM8nYudn4IqHbEEeuScGJJmrcyUXp+uSJXI8tKU6Jp5q3MNuiLSSH7QU7sB2q7g
nJwMk1KSSWlo4GETuZNQFy9UmzVNxI3sHR6AvocE25FcbauMW6/w4f1+/0WxvJVJ1+wbfZnH2Zas
qTEQRLlHgmhFvjVXYc9zN8cUKneVnJIxQO7LdCJ9K0h1kY5gfAdd/Uv2okSIHn8O3kVguo/VhYD/
JOIgMzfApgSnhqMimaFWFbrfuRsHMe0Xs16KMsf3DEDzhNyPnMtUPu9xIp73J4MC7BBLoItF0ahN
g5Wz8QnO0bluP1YJn1UnTT6SHGPWycUC3E3lRq1657CyBAsy84cPkRLhQkaV3Hz1l1GwtibNRXhx
e85um/AeJAaM2Xzr1jX7ENQaZphOKfheC4IAFMj+UBZonZiyprNYJrKiqGgy0uMc8/NgvDMn9aqF
Xv56AQENgsn8iEE0o1UHgBL95CyVX44Og1IBFVAdk2sdlZSO+dkj4cnFTbyV1utRSfLlgIuMJeB2
Ka9fXwyC5tebvnlIGA98LJ70qsi+Q2mEdEmwt5jR/IX2gKeAypcGUSt87vN1OLpvBcLJakH5wOL2
rg+EoVjeOpDlivsLSHG8prwOfW/Bar87NJUNtDvTx4mLuTKVRxewoJFpvj9TmOERKbrBWtuVRL8H
5ih7B4Txp1eomBeJuBCcEhf2Cw+tSRHoOWpDop5msjbdcavoNsRSrSsch1ACrA2ipb/VKLxpg3Hg
pdvfKOjAWZ9yrvgRQQknbW/IxypuGyfaEdoJoW8BQygj0IMdxa3aIRPPLhycXBtLIRgiaYVtN9jN
JiwUGeyu08gPJUiw19V5il9cCaD5cTwfIyeIRb1NgFsiUOApAc2soA/ipkkxOjNhowYEz+ZTt3Sq
14EFKfrPvIeAIu6tLdcjYMJlRXjYeYdwJsmZAbNzcqCK00H/zqVu803mHe2JTlcHyVZcoVVl8/AO
Z6kpfNVBChdMYYJvssHiwau0gdbnHZ+fwe2arm+azyIGXz5ZsjXlnz+aublZPmcQvR6Kr4b6+jov
FR43DrWn0PMLljtRHuhIQiVDxWIVayj0d26ejygqfF+NwykawezSg8o7nhpJVa/84Jgz44K2+VCV
TkKA6K9gP0w8Vd5esxCvzNzqo1d7yrQKbEcS5eQOQ88IuYcR91+qRl6yys9vKSML0DAmNtNRGR+v
KbGwcZa5RZeFzaLEp4wzJ7jnpTMRFG22Az42B8SwHpTJHXFeaRC1yR+V+RAJQEIcJtlU1bHb+OFl
rUKGuvH9bB7BGbB1XpxFDVxjZqpiKdbiIzi85bZF6zf2YmBdRVHkeyszWyZONXPtjNC0E+m0na3a
uIPza0qF2S0as55NdM3hZcB6yy65jwEXSySu1mjRPkOboR0s/O0ixAWgoCVXiq5XSSXKftyyBt4q
1mafNNVLsUZ1oZiGA/gPo2JHHTnuF/I18kd/CIhbZn6FiM31FGrfvwYr3KWAGIwhee4bwQxpkNa6
DRnGQ8onD6tZtjVFcmCOQ3lx5X/YfoVW9kRBz/3GuZVEGO9x6K3ZejH1AK2Kre4Hy8G/QEe7PbVC
1W4suVjZm/odtqmkzExlduYSOcbWdo64HK/0DBjJ+vXKmTW3YmLjIPHxo16rAPQhR2zl64l1f9AI
1Tpjo3ObBZxSVhqsZcF8ZyHztOdpMrJCy3Olbvc2suiY3QvjyXdIGJmisVOkLKxcicstZN7DcHju
M5TYIHT0XHbWfq7Fm6rbZKkhjNP43ZNXP9pguCmErA7BPcIesoURWLAyNHNiCedTssq9Ml9L8b1G
ArUNIgApduh4HHAB5MCLcUgbFflHMABwVkW3CdKZDUZLLutTUBHJeKRRei8reVo4npwnTWd2WBrd
zTImAcP6MJyc6peru0yDWEP5WNkCgEL2vhSU3qOjNsdP9RTDItsb3zPo1BXqFmmcR6mm9neQdTxo
adfRkWvGXQxk5lqGRDxbNiXD1epa6MecAETkAF0RbrfPOqEiNy3I7N9g4ykI+6fI8454OMpgWSP4
w0go6Af2CHXXQuvrs52drHoet1jcZWmuDwzdfpcFDAiwGMh46w49ajeRvKpeDpt+SHvHDd/tAe3l
hhzp1M/M6RdeiaxqwdpLtD3Tkgo2pu/1RU3QzcpbzOB8IQKPDq/IZQv7yH7b2ld/OUAIK6AYC2SD
yR782PPws1s0rNqv7fY9o9PC4yRrMAR9Za2uCWLuiNOp8JwNzLHtuwOSt3mMg1pyOHAXRQ0+wCVD
l7lWm1WQ6T/0zrRcKbvlJFnZIYz1eRWmOqTmAic0cbDKBrouNcux4W9ndVCqyYZBwjNdqpjaQwEA
J23KqnbLOgWQDvJLnBKMeZbaOdjNiGfOFnY1Aava+yNc6PIXf4ekzIgH813flD7ndcjIe8cCPjTY
y/57s9hV+kVvWDjdQGxXuwDJRC7zEzhZ4BWmp6NE0+BaqDXTTb5ZKAhDWhAFuUj6VoN1oFYNKLGJ
XIotlLRyfIUUwIW9jc+TgnJfkzVUwIE7sO06hog8j4q569VcXPWXs7hXTvcTToCmIbXlhE/8V+D5
adVYJ8uOs6A5ccTfthfKyxrQvZZg0Emm45SrOojnjB7YqrJ3RypzAjSPXQuQR+Dx8i5vVn4yokBq
f1diCW/rK61qgh7jh33B+P13GqjnwbhXHmDjakfWvzW/FanfaT0y/H/Ez+QbVzrsX/m01DjPAazU
CVvke1XfMH70ZlUFExXdYX61A+TZVVzyEKgFmrVRfBcB8EqUK35Iuw3XKTFer1MaojIOuEO4LkJe
Af9/JisxZlMcAuTbWqJYwI0MWNhKAHxSgbLrJM6cZgVaMB0iRxEZ+WL48uBOqo1F64J+WOxWSGrb
hdz5L9BT3h2FQZs5cpE2P2faArvcyoE8VhzyZJK/vE9jQfDaDuftZ28Lo2qWME9MF+Hi0jXTNSs6
4VAmvstRWrpYjqAPnYFcrQC/Kc2kSSYV4vV1H1Ibh9DqH3qtZnDy9Dv+tibBCeELNeNtTy4qHUw2
Bj26GsEYouM1fpkeGLeIV33krIcaSJDGrd5pW7W6zmcj44UaioJ6v61ScIB80v1QNPxhclxYmZhP
L6QfcuRrr6sHbjaQ6mC3GmOBvX7AcxTp2nWaahnCFWOlpUlIn36VNAY7ZDPZuYRtTxzYL/XIUzd/
OURgyRr+2TttlzMGyrY1eyv+T0EbZiCfR7WlOJZq01oeDWeCLO2eTIqwCfyTGf2yqLEdz54fbefx
7rENK1HhawU2tR1kHvlDyx1wCWA/cZfxKzZaYyPyQ2dHV7xlmdtYXZDHvNtwf9vRoAXsCUeg4dR/
rW15Lhb98d/TH2QcCr/WEBkjFGpEXHYPYnZzMAKuTn9qqPcGupiOIfIL4OWvY2Ktu0V1y2MEVu1B
MSTTT5nWIAFzbKd+NTp9xY6zXqONVm/UmQWVylCzGP7/9x7Yh1XPzBwkOeXuhq402oYM86rH1JHw
t2bG4VKx7n7pVg++df95qhwVYwdvM/TZSTVd5pebsugBGBFMyUYXkyaD9pv6TFVTKaqrGqXEaXXD
yURYq+NE+M1uXpwie8SEBM7mtnnVaR8ca4dtV9ySmCoAwHl3ixna/DXEZxqHFxF5bkA0f3ybEiY9
3Zjjc7zY0t5oOMjIwIaSd6069USO3lEnhuol+66c+hL6TaRaGNpGFjFrz46tfB+Ra8iATD5Tu9Eg
/OPmXUspaaHNoiiN60GVzaYc3zqZCDqSN3Yp97XQICTej1jlhgh3T3H3x+Hq9VJKQoy2WwkukqH1
gmub2SDFfpdbfftZg2RX+C+D1u3zCcai956GjqPBBRdE0qN64+64mBxwS6/SxPWka9xlZ8spbI0h
BaZpzxxKuEd4rH6ORmW2T2uHAMtLNip82GcPsTMvuMHhf37IL2MWvB/tHdoMCo+Yj4D9mTsUFgVP
Hn9ySYPVyowOKy1U7m07AtGuZ49CXJHaf+tJVPRaCX+KYd6ehHZSd2GmZj6U/NwvVQXvPvi9Awlv
xjsK1GWTxC32qzZQ7QVgCa9Q//FZRRkylgIavqHQPupnI35lZsOQxrzJF4UwoJjS0fzXoKFDxT1o
ji5ot59oyUMZLv/bATYXsGR8f+0vcgr8knJN452AXu0DOV2JhuOKQyKqxxrRcdu6lS8wGKz2WSM+
PSITabLepXzO7DVrpYUbrXKGK8S7G0ajUZDe1TzSkE/M1NcK6LUp/pr61zZe3vbXyd5/ybCgZvxU
lxK+xrMnMtJtYtdekZ1TFOhqM7Gz6q3RTHIa6emtMQoLAQqBBdxfLUdhpxEFbVwglEZ7i2Qsx/M3
tTmet19TANuN2dPqkhSCZ+Q9+cDfRzkxMKm2We2RB6WK9Qp5WBO0ewkwffp0uqXH6SCg8p9xyEPE
0kSDPTIpVMfyWw7GOZ3VOM0YT3i6ov+Y+XWng8+02nAzMTynMnhgFff8UrcysNpcSLH57aBMor8v
IoiL4tJPiFgcqCz1KfpA3jbJo2y8prmv1POG7x2eUO7VnC5yp3hVxo4tqrbF2FCLdraDUbywV5DY
w42u201ZvAxQKhQy7DQ0H3oor8ebAcfQ89p0EckR1X2moLIaKw5LvbHTcFih3Pyq+BaGP5urvQEz
DpyvdZn3frfySY2JE50It0IMzAbeQI+vtx25Dy/dwdVZitrVgbnrR06T6btIENCFUapmSLjKEfyh
5QBP/qWHjBNHKcqeFiG+jVEcimr3ZqCOYZvNZnH1eUyT2fIEvoQHpGF2j/L/Gv5dKuhaJtXx+AeN
y1ZyQhCgszPks3kH/IlIjigyQRDNt4FpTmPuy3EjDema/BTNu+dPKJvWPVnSaw3Z4Yj6BJEZuJtD
kqeMzgWutv9z6NVBnBhwQ6YdkDruso/p7cIOcr+I48cYCbfP+rWU72C1Gy8SJGf5hLgbEkyUFzYf
HJY8egg8b+jz+t5GA2oOuQd2io9UhL2SDzaS12qlLXtrr08rVRvknowXftogTp10HKm7tWu6+FLf
Jx6ATPBxGi+a4sJscVeZ237lcOFX7MH1sxjGDrPZBQybdNib3ns2ZGISwJcJ2uqTbICkrntGBWlo
+kkikmEQjOb//M9mGZ7aMJVJLkUjUJOeIkB4DfUzYLkE53CgfymgYRpdvwFU9mpaEu+J4580Mv/r
Mw2bfravTJCzh3FgLl2DfzBmb2dG7aAimm8V1AB7HzkUJt4AD2NMsdChFy/ogHTmCCvfenOLNCTU
2tVYzcHD6jj0N1p9zUKUNtjevh5WQR3ezBCLjLCOmJTNF5p3wJ/IUmhdKqBelo4Os78qZxsMiZ2o
4Jt44bZH9f0YDSmz0bXFkoZKF2GRMBOywIET155NH0oH4UaIgnkgLSJb/CrgDNINV5cHcBktMJ90
9ANRoww86rHcGfyKEw9fF+h1BfkAAmvIAw02+D4HmE6TyqUedGVWX5kViJChD7SuQ6Pkdv/jSfGj
De5Fo5d9QAKVWFyBbEaEuPFhklectFjHR9WYAPWvCDyR46NKfkcj0Ht0QJko2ZjSL2+zhwDuwzt4
SK1MeWcJrg/CilZULp6msFG6VSyfwl5UPg13nJF6W3fXIr+mRMgBB3FlklkWD6njpc/eqpSiPnqk
TzLxbuMDUmmIXU/uwO//ClTayBLMyOaQP5NdLTMYo4rt1AqVAiLKEjvPmvXa0ZqCEB8sUTmVN/E/
24ciQ+DErwr47iZxBu2SLNo0k0vl7B0cV8Mx/8ER2MtfMpfz9zPxtE2WWcbD+A8GnUtnxvIi7CUt
0+pQoT9zoz25UGn7pb0SoeNH14VN3iP9ZMJzOBar/oxNsa2u0F3XtpwCAx3yRbetcwMhGFXr9wcM
WQ6+Fj4Z+b75oH40gAmld1PDKAtJOUkcodNgM8GHb/Ik613GTTLX2fxsYrQJQzVtNxheZLIVZBx3
tI08hL65uhnx2XPKpK4SLyN6YOFdaGGCKj+UelkqNoTsGfRtntwy1fUDHNC+yRdTaZE59nVdAeVp
byDt+kF5Y1wtRsHZ/QJmCAwJi2n0j6cfitgGotN/niQ6jODJVzvW/jDuRkQi3x8RXJ6rwrde1iXP
mLU8hf98YGNMkD0uUYv+pQGaL5g5qwL12a0gSbc0dm/xnKdnjIc3ZdL4/L1Fo2xWGLfX9pla+AD3
chFXUMv4vQrchy186PIIcM7qe2LdAa0aWABxNn2pcfWgRUMFMaJx7mTE+XQXdXSmcrwStpydnsqX
BAtTX51/qGGVoK0bZpBo3KnhWWYYqFxF8MKBYv/q4SVhfd1vMB5ox7fHKIz2ckKzJQWqsJvZsW1I
pns9a9e51FbX1mqTyZZ8atzb+5FTgGtZedEnDWP8zI2vHMK9+SjINAPDp2t1ta5BQM7HZJC6yw8i
rlOL6pIvZLGG2xDPGSURMelyVQ+PGDSjEa7W2YqblWqe6KgpmPyhGvYf9+kUDbJv62ezPmCsNTgM
3Odxdu+gur4PAGPNsW69XuGP+mau0u4Z74jQODPtRn46w6AI5Ua/v0jtsfKxgk/XJ0/pR6cJJoH4
XK84kVws9q8D4FkMgy3W6rG8NGUKVjsgSCQetiMJg9y9jpZCVJMqPxmjsh8Z6ffjKluf395FV3in
awvhCobnr2WII78OTW4G2MFbwNgW0Qo3nZ0mr4nqGeppKyOPAazmOL7FeGI5yDqgvyorDXV9BS85
SQ4nBSEXU68MoCSXErWbjdBdhkLkJHwf4qK3TdHueVDBYJ2aeknisi2+BcprZzQN+ztqtiWiTLKf
sZjHy4tHFDqEfmtYhjB5ZjGLzAYRnbdnc5RH0pppAfHpZDIULH9UwBeLdpwz9QueYiWM9T4fH4QE
+ogKvd2HaBT2mMO6FPvdONPbXYjdbKmfXF/POFwPxleSsWB4tXwifujlR2+y8us5V8Gt+FBjNve2
p8QHhNHFwxiLiVkHVShXaDdFzBrIEq32q/2NLPXlKWUzwYmFvGjIbDlO4Mx23+b+NPOJFdQjyegT
y7MxbfFO6Q1PklhhEiFid7fzj7R6I/EUjXmQtunzCbIzf+NQPZxl8O6hn8jo5AAP4HPbTlvOUPa5
qjRKVBC5hLl4acGjJHI9Z9P2mHxAShuLvR8tTOv8I2c+8eTyJQC5QGEH5xRpyPwFUNwsMIlPJFcl
dYlAj7s4CDJUfvLNdDRTpHSm2HbTmoaxaTTBDACTyIiK2dm2aFH2jVUTXdIflWwGXlI4e1iAqqVG
3R+9It2tzZ7Q/KsKcKt3wu74Iypdldk4l0sQwvlfsyW4jpa7ny7GimQRUwoVn7ZdQfzTQ1NhxwRx
rIxomEhrbHhsNv7nKaJkeUXBLDgZWfUpND18/aZ2UW1D/drYuAnW4a2YIuI8BAa3fK4C771sluzL
6sPO9S91hRD+s0StYxmw8AtUGtL6Lwtqh0gWy2eEWUKUO6WCAzhaVRWOqZc0lmQ2z4cF6pdnTeXk
B2oIQR9O6r4Wn9b1rn9KLUP4WZpfjWDB8pJiY3PpmivVhn8CMdLLJ1dLlyXJo67B6BrmnkKScD1v
E8niBbo6jssp9VkKzSwQvL1iKXGBxbXOYIT8/yQxZbHLOLyBAxsjoARBJBXFNAQ926KSpJkcddRT
LrxpwWZZkhwfMtYgR6QR95eBuXykKcE84gZNLgvgj9qJVAqLx7QaVQ7rXmuXYyssQQ9feWFdghlT
pS1jVikKA4ZTL3pwDmThpGnN7rO+V5WffexICQk6IJnxRjdIkE5ilSPj0XO0LVVtP3Z86RwTUVa0
5btg2L29R39R5LLzVlKMrf1EKWTxxksTMSqSgjo6RclWwvqnomhnhfEDPCQwxarwkUznSsTCiD6P
N69+EILCylK4R8i9YSTBZo4wSBra7vHcJFXkAJUILr3KRCck7U7wp8WZ07916Q7o84RyYN9LW5lb
JGjLNoRPKgso+uo3QyVlqOPBHeFv4fA+NgyawTJawfbug/LvgLUgz8bmzfKrYMPOGhxWC6KoLov9
4mc9hLpt9//wNYJlcndjmaofY1S2nJ5RH4gzGORAyYHL3ZAIBItZMTc71lMippadiR0uvWmNtsqx
c7KStcTqvwjZwVtAMh+I0QA2ybQVF5SDbHNwwtYqon5XQ+YVk4uz6ulaD9nHnnkaY2AhFrz7MDFy
su2UWsUHjz4mTM0CBQex6VbjIRh3u9zTGVJjwN75yWEParwKnsi0xRZzzdytl6mNDp4fkBS+xq9y
BFuWjPMDj14z3iudyzLcCuHtOfY0ocDxxYN4n+e1eQMuE+kHVT1bUpoBThU/QtgS1NXMdyuC3UAX
hT4GgbUUaFHJp+9ReVPhSlHKwZzvfi2VmJjvsNHDYTq71IFmscisZv31rm15k/6oduBHDWMWvKrj
DK+8FoYSRw6R9xLWUDi5fxWVm/Wi6E2GhA91SBvnQQuTyfkY03vkdOHqTxS9aIpch1JpxiH2HPvQ
iQjm3GkqtTRk2N7zno1zPikauV7e+BFLq/N6L3YWHaY4yQm36k6NIsa2hG4qxmjZINz9YcbwBUg6
HYkyP+G9TB1aedQarPllhaXoiLAwNSvT/TyiQAkXNoMYRYc5sngz0Z/9ozrJrG8rWKDbvxo/0RZH
ZjBA1chnLJnQqFPT9jvJv2hn6prZtp9oYgVDhi0zspt8k02qkZmGQ7xILSV5obqZ1/dsOJvFjVjP
K5Q6iGQrME1h3eDLvS6HxFxTIrBqRoZ0iwDjXHwfFsEjkw6UQIRy7PC+X1aE8BLz4iMfr3mpN5Cy
2IVlXR0x6xIz0rnk7UUYfKdLEhZ9N7QN8E6NuN7jitIZUl3dMsHk7R2IArpkl3ZLx9hGrix6+yHx
uV2iqGW8PZCnVjFjOTNhmIbpmelhzq5FG28B+cN2p9/HSE2dQufi7BKzPTvs+lOXT4ztfBxIIMnG
ZH/mma13r3Fw90DCefaASp+4RQq2WJa9kAfvmJLS5QjA5jITSKgoMK8gJggGNadfYQ6If+iiopgY
u/oei3ZXkWEse/3mYXJ1Jd1E/K5KY6S+C4bf1ceFGzr7yhSGY7rUfvVH/xIgazVqP5DZPaLC7sjB
MJbm4VWiDlWqtW6Gf+Czz2LCPQoMXOtBTOmTlGrpBZIgi9FLCa+S6lPyofySkH1g3y2QNbd/KFTk
S11vZTjDVd6qqP4oxn8SvCkWmK490LWXuGwP3AOuS+65ERn51FzJeeZmnr0iF0tJsAsga+03rj4r
y8oLhhxwBfkUanx5aQp8Tx3JsMPs7MN3H/Q2DCj4fXf6M50TBaBAiFOtnEW3zy8KOkjE1aKJqL5w
o13XdpsDSHZFnPkwKBEjb5p0dCk6WM9HWwUT+Vej30762NmqUofPv1biy1ck2Hl/VsNZp3NsXxAa
zR6+emJFIMMz/64abf6PNMAXJ1BOcwRtCo6OvSdeXCuHaZ4HHn0TkG6p4T1YZtpAkZTbkuESygW5
avI7HTdusAAB3lPpvp6L7fCd7CF8Bq4Hw3UZjb90qXNIeHSyf+AmHdw6I4bwCSFg0SkVUsa+KHL8
JWP/DBy+JsYTI7ODmGE63UGo7MxZ5P6OtG0HGjoTTP/L1CMjznbUOhFvwMyq6aWKYuSXaySvd1SB
Tg2cDrP36Ui7qmDgeQA0W6d3aSu8agZW9+bAYiyjV97VTVROdO3M7uSEsJ14AM5hmtfQTYqK4ivz
6D1N/uzI2MMRqZSZs2vHaxn0SKK3kFbxbsFRTO6esFWjdJLXXwFDVYm3aUQZhSGHcQi89+yQgOBm
CYR8obga4+QnKvWh9W6+9coT/4TLLTFxnc46Cm7sXZMxkyR+98GbfiR8nc8E0zIKiWKmeXl3JVMV
0ldzERiXJPDo5peI3IlyWMrbSBKJDOaDJ4QIyqvrKx4LWc4kpSYwsTqtDyLWrt8CsyRBxPqtmFZQ
JqDsxO8IPtEFc8eQwlE2ygjsEFkg5UZ0g5ftLka50JWHmMGFFvldDZSy9biHlWPOH4r6Fwu6yf1B
x15dJkN08NKLueyWkmazDl7AHFoXe7g2dsCeiS49UEzGMYzqxF7nIUG736P6nm62VP20gvBd2Jd+
DyxVM6h8iXiYrgf4kT6FsWyvs5X1MmsrVU8GqAbphxPlCRP104ChtAnKl6lesHF4nKhj0Y65CLei
sIiY3+sSHOCovBjSApxINdwxnRy4gzzjITSUPzi8OBQgUm33eq0eCkhXl+tvhcq6MHg0kyKlYli4
fs93K4rzoBa0Hyru+BOsFYfttgEPpsvEP0P+vLrdfB9fSVXshwnATki57PphdebKa22MHjb9r5SD
U/lg7amRSLipGdY9ZD3EP+7kIp59lYngDNgc4a7mihFdrvAA0jqp8Zzb2SR7yKa4ORbBAdqNsESt
c+5GZYktv/LlAeOyn6cjYFc5jA6S6jfzk/2ohYpa0VNHlnV2aiibmykkUnIU+VFN25IgepAU8uRV
12alNHmkqWJQ6Bp0ACwWrNTF7SUuTCWz1OyNg9JmT41xHWJ6WHWc6/Jyz2U50Zsp4XDxTRTi0f3c
CKYPbtvK2Gog158IcfwpE/rmbL79xNJPoWZqDXznI47N+lcv4/OcOqLG9Vp3PCTS7G8CjhADp1Rk
vQXBt707OpttJtoiKsY+Ngd7AGMWsA8vB2AZXOGTEBcCiCMSv83cjXmp1D5RxYIH20KAni72CMTN
H5sW2ewZTliYURJoKrUKFBP4img+SnG2ZCKsxaATc2kKGUG7yDrv37me3wd24E1IbmrCz/xz1ou1
+Jn7LvuxRsnY9T193JW+CbM44cfmpzvSm9mVEXjiwd0K7YGeIJQSTZ2zVV0wCsIWvXGbNn9b5rI+
OQvF1Ru9ZoghBonetA/lrvfJFvtb1x15I9gKYePpjDOgawi2K2JrrirCnXPDTRLxvz7vBkh4ZvpZ
zOlSBhDUAwPuhp9VjXRxGnVJ+vdbR5Zc/14RkUrYZZuooCDkXPCJ8yvgtrwLJQp3xd40w2voz0H2
htlAzzmlDLtPnaw8y+NthmupPlsUV7wK9y41PrOZC90uYBhoSHedc7rVbOn+zEv/MlG0Yk2vyRUj
ZKjk4hlM+nrCES1dOZlY7iwz46VLJ6i5V/J3SMsLiewzSycKdD8dh4fcmQqleBLAun5UhVVJBtQd
APpnTteSdik7rQbm8EsVxjOmRvvPLqNDsziX4MAbAoZtNTxWbtmqvUrmVMeFhWVezieWtJ55W+Zu
eO8lqTmOugAqzmOtqd45i0sYWVmlrdogmAGKJkRerO/kS8qlAqNvIQTTZV4KhF3tY5bLjMGktvlf
JaZDy3lyrnSCPIpcFTSbjuRiWAZJwQC2LMCmX8kS+QA6HgwKy1WB8GZJekBtLH4ltRB/VzpDk+pG
pAWQ7N0s/EiOYNpLkMIkzgXx5T+lepPiNemg3IOnvqhaaE2ULk44ohaUxro5Hpm0wCdsdbcWiB6j
2nybjna+D7KjEYCfV3p57sMFs2Vy/ViwUWr6dybxwie4pcQlkV7DqUmjLpDo3KMx+vYzRMp3v5fy
yuK+OZXlIR8OTRYlMzWWqYeVYFo6yx2Vj+wCarHuYvwUz73QWdDCq6jmbro5MVYjsiEi1XCdEYx4
DbtO1tDBv2YL4+mqfYBRQ2lpYWmPgKY65NpPUkS9KPHILcme7DQpXYCInWpajR6Tlux24U2vwmmb
U7lBVaEcAAhiyQDVBMwkuibwi980CCYaP5iuHHO4ZvtpeEJP59IB46SnxEcKZeVhomPiM3po6ZGj
LweehM7HsHw/0CZo8dxsKkE+5AYzQ1uuhivdf43Jf4QvQGNHTkiKQSe1i91BgJjN75csSfY47Csk
vy6t6KnwLf6wUAdWhvNHcvJnz6LOpF/kWAt8bE8nz7lX9XxMpftvrra72nUOq6t0MsT44turwM+l
ETm7v4j06wWaER5a5LfwEgMJvfK2dNCN0vNftrm2bwcLclQaNXwTL20uiBAdu4wKPzaqEjypoSfr
nfhBCTuXEaMmZE3FKqqtMcqoiww6z+DyVQqwLsDBFkKhGMHbMg/oLuVsbh4r5yjQHfmlJHabww93
kTriysSeKLxCrUVWA+8hAj97ja0wFgfuHk/MTmPXYK/B3WDNZ5O/dxEE1yPLjW4o0R28jPeaMHwh
mM7p7dJ16FSFz/3S0dTftn6TScLc5pEbDwZXw9apB+k6AQW4SHxbmd2cdinkoHScECLYZ1GYnGBa
siEzSFEO+5f+ZUYJClPxSedDT5KDMhgK7dJ0YWjXa0QDyQdETxZ2ibRCU0T8Q/SXegxPcIwdkU1F
nOU/ihOj1MLaBRS2apv5q/svaHjE7e5q3we0Revn2yrkM/qV1i68ZnWxgBc4IUfowQFyWJzVl0nB
55f+iaSPh33RO6NkI8qnlTp+H7OPwxb822HQGCcRn5v7Q7WrhT5vJvUybonr0VsehaaPnuNbukjc
Le69yBJMZmj2j6W3KqM2c80J2FK2peRdGvog9znP/FQt+yY8vPo6gsUcjvO+MMOfpBHaWsb5eDSO
thBXp5lGF1z7TvYoCUydlnNQRCe3zmOVEXgqXlx5ZrYOcY4hsgJ40wGvX69fzC8S/91PTwcjtxL1
UjONEdE0TzQAo6g7csA1gZqm4Il3pPagLkxGW9z6WA15iBmlksKEct7Slr5eh5s6VaTljju5qOBV
sL6nfKdAoPaltKiKCps50+k0+uB6zL8FmkUN+N/2++iaV6Imf4x8Ekoy3VSNjIoFBA6ZTo4GmdLt
j6lliajdf36Tkv5/fohXWB6bMN32n8n5M2ktaPRC0jU4Vrb9SuOicfTLn9WX/OKNhoV0PlKQhs7z
nK/SayBzN1Ha6ttmcrpGFPGyE5kn9vtcNALLuMLB0IYQS/+DGxvfdNErYd9Sn6ieMdkJCVFd5JuG
J+3S1bMxvHFq80mdCr677lnJoUkbqi1RHKB7mXg+1ZvocAk0ihXHa0xnje2X/CBVQ7XqXZuPi1/k
Mm7F0FgLUCiRirksSE3X/ab19i/6f5HuShNsllUBFNg7ou5aScIQ3TqXm+IO6sbNsg04L3xNhxwo
iIf/sYnha8bGHjL801jTf1VvmSSt95K7E++t0feuirmxf/R7PlYX5W7tcjNgOrBhjKquWer9sVTP
xNkzalUrVf3tbdmtkYDBBfsVU52mkiD5EB/YsM4cGRHt0dbXSjTcFvFEbA4cjq3AZlY1iJdeuAyL
3vFYTuDzvYX5bykhxlaqbO3HwwT7fznrPAiMchT6Q0NiEYANHzXOl86CJ1l2gGcOlylpO+w0Ou6V
bCPkNmqZPkhbae+fiZ34QuYRd7thcJ/IS4WHqixO2mZR0ZrgsQB8zoiXlsnTVQ4NviN5Fc/CB76L
kNxNRFlbmXZlwgbvLGz3Y3yqSvGDszPNgbgPJoZ4Sp5DVb3HlCn3c5CTmaVRwnTggKY5Jd6BhiC+
xWejRiQOodPtyyiJI3PFwxF7I2MNsZ5iSOtbchz7qPyNg8N/KP45ULrZkUEkiaNopUFMrZKeoEbs
GhjoFknt+5g83Qi25fpsCVOJRmcMvVb8oUirUeG26b1u1J1NxlSdgWZQphZ7zvWqGeboq0epYGcm
PTha5VjwjRKbJQL+NgTefbdDEe+3rRH0eC2uo9oNK2jzOuVSklwpOcdeUrKmctqa1D7Q4tohCW4n
ybpaFkbFnnxQsTtCcOVwx6ppryY+lYC5WMnhW5R2cGijHXXCYHf+DokvoYzTKgp2bLpYitfcpEKG
RVa/Pyl3clQJCTuqYpXYN/F04If/uUjHuUCG01QHwd+OMAzvj5zMJ4eaaIYvUc1j+CzxYHYaKGnf
xNlF4rl1a6Q7Ak1hcUH+bFtyJvvdN5kaSGoc4vBxYHlh4G0MghvKtKUvAw+R0qBY6B99Mzy2qykP
AvAHGLrKtr3i7NDHakjJJLBUxkkbAqqGdsnA6xed+7YGzLmDXvRA9Xh6TNvdhUliliIYgrcX6jq9
1CsTMYxuWULMo6e8L+DvujTRUkhR+0xChDBX64ETzNAl4xbaU6C3LPBEO5m83NeIMdM2X/UwdDLx
Lwp6ef7rnywgmyYD4cq3iziFzKF3wtMKwf2AhI3RcLt4CHy4vfxQ/dHA3CvyH7UcC82aUVMIhuRG
66pw6Ql8RJJb7Qy2MainRoGR3+8qENn3EG481kXxJ5g/T59656D7zHancVULOC09ezvOlLj6j5jX
poPRHVGmeorQbg5z0JOFulVVgmp28LKzOXo1hhzZQpTSaLw1PibGVhAveK1x/V+S1E7BJrsugSzj
v7hmp0nGY/oLgx16uAvjEfK0tJfNo+6wAW8G6odr3g2JjsjeqfBZtlY4YyAD9SIJG7OQxDbOhc80
+AOTT4z4D46SoxAUHz8mtMKz73KhLoKnR1Az6NmF4T+FVIVRQvh9apJG9N7aTREdjtpbAungrL/N
QznjaT8HdJ/z+WNdefe/4lgUzpxLHDi106fU+MDvsiHVmB1LxG7NSpjU/sAAIjznTmR8XHWch+OB
51F/N5nlhs0YSE3H9VthpPiXxJb0jcXhYKx6egBxCgGuF2A5RpXJDbo0GEuNIoJrIbhaRxc6Zkdk
I+M83rnzIlW0qlZLUC1Nl/6FlKHmAz3jDg2slJZ+/6V+D/dVkSfEtWQXyMZD1R21l3PGv0Chnnqx
TCQhR6oIIv1O4E+sUtYw8IiwSKN393JAlcXjhV8oXUi5YRwqF9VEFSeOrs2s0X5kFutZP3be5fAb
on6X1imnfVqr6DzgDgp2hgWqobh8jGwn+QBxOBVwg1ealpiXR+tvBGNkrWRW48ZDzjE9jL3mnsR+
KcT6QOx6kJc9av2z0ygeErSq+Vk91AAhZlwjlv1IWsNpw/NcaEM3vVcosCO2UndFJh6lczkycPfS
Dbq9sCWEKQE7bY2JhGW+BI5R/wQpF7Q2I32n2sFSIvlIEgY9oe4COZ35nVU0obPViZWuBMuua+ZO
YE5iBUb8KQmm7RsXNbs3Wcx6ONwMla6VkeQSsfklDA2g9HmxOWWY0Ih1cq79sRC6cTOEAXQXsE3m
sM5SoXmHkFo8cuvoqvN4gqstA5pUjsRwyY+3hhoaRPACirn2W9pQUFi0EmmqZzUNSS03k1ehYuZP
z//RwydR4dUiA3ni0YldQB5RSZUh9kfX9Tq8hTI0tHh9Ruscv7GOm93UlBEYkuQjxa9jcmyodxCE
4wRGzPlHWHT5wAc8OwYIHq34LPtdYFUqcJIyNBUJYM3RfAoq3NREUSudeGSadDO+6P3n7NM2uh4R
tGGRsrg0VbWwRo7FBvneSxGTRG4Y1JJLqBr3237PKFTiBdiMHiBgt64/ncIAR8wjhycEYM1ksf22
hvSIEC0T2gnDulTT7XDvTmH13OpTVF/x1/wN6MqBZVZlv8iwmRwE4q1UhMXToj70XCuOOOhyukZi
d9+7vaml+L6aYoijmVCV1Q8gW+/yCP/7xHmLA3NSdO8VAovT4RdLh72kPUWvdXlgI5oar/o2ueFO
yBNVn+yMSNABLVe1pEpLtmBNr98D3lDuHtj4eY6pabh1ev5UC8E8g8MK2p4P4xDhgqfA/D1Mzur1
i+uOKYD0O9umUykfkrPW6DSX00/dWlXq/DvyqnPazZF+58HdKfdKaijKPa+YRsrTT8Qves3t+lyj
5TjUMNu2CgjPQScBj+pF21osYf+TAcoOUV4Ah6yA4qnKNi2mMK+R2Di6FKChVEVonwjxKDL+mJOk
ktG8ZKrkzJ5HWsJ2shql2rSI1Z2cZgEGogaadLz/1MOtjXJ75u5gua78tot80WQtcun+as0ZVto2
H9q0uJPuLp1qNpjYA9M6xBDNXAkBxNrgZm7EsJxWbT3g6XpefMBpDpP7q0Sh40l+7V2wlla2m+28
S6LY1gGyXR9BDbXu+N44JROrbhdNw+R8QP5pLHAXh47U4YQdkBjaNSNb3lwmb9zzvTrMabTkONkI
mkt5N6f0v2z+R6DepUgMBDVG9emtH1Z5pPBaVt0dlq2gNb2KTm9wgJfqXWVvZw5u/DWqdenmdqdK
P0EFHdPyqi5MkQAeuvGUEgIkTue9GuMrV2hLM4UrNIQAgi2wAGGP0527X4zfpR2BlE9fiw8IsWlr
tsFVQvVTRSdpuLibQan1jfgn8ExxQs1sPErCFBEF0hY7fni2vhHMCtYp+ZcEwSVZBx+UoMzIw4UI
a2rSiwMPioSCf8mOV5xyOltvw9kau5DOPCvJP53J+VA7fUkLOmoQUL7HZCqsqWO0Qts1W8A+mFrr
Oc/R9k3Ou+tGGsdwhBvnJPQEZpYOyYG2kYsr73FWItCKIvyK8sXG1LqVf552bIGh/bDLS88vIPd+
16zcULGxsSo//TyCAeSOAOpxgqpKMr+qp43pCzkf34HMJxDxcMmAcc/PgNy/LKnDow/sZ7WTYuqg
N1cxyMU2LENJ0iFjvkCf+RMiCHb1CXXIdRn3CaMrlESI02Jvcdcl3L+g8lrjlrO9XkUpOa3Fzwvi
/paJGX+SpJbXuJjka+LP4FFHMPTz3Vs3gKEZD9UNYaBh32QkR5y1Q4OND9zvseis5+7fxdxGu/7e
XO2adXKAD1+1jnCwPrqbMU+x8b9Mec6G064Fby7j2tmU3YCBthEZ4VoStw9zh7Oha1eOfxfPeB/L
Zn2EhW99vFsVvYLwwsukdhbSzP/cfBoghMeS8ntURKS+A9Mhc0wMrDJILC+7GRhMI2PkzBWkDl5r
uQS5drWPvTfGRIoSUi7stX7tQSjQcnQHnEaHo6y2WUIYKIwI9TOOCGHOrIuT23kta/6Ac2UXNFpS
U3RsPr7ynYV7sqySlgzus8CSE1u0Vf100s/gSLV3Kk+WO/3UOpTDPjq/VT2S4O3HoYfgJnqM4pL9
JaKlDF2neCq3KUy+MtxlHx2tJxDliu8lZbJcrqbweOiNfS1w/jlfYWRidIguKLMs04MONU4TmE04
DzWeC50sVWtWOgrO1AO/jVV/ybbcEupMUpESPaIqCvpg7t9b/CgK6vxKUb+rsPSwp/n1jBLHST7o
yNLv+oRhKwAw37EEjUiLuIOjrFhzqqZjpU91FUDKZBaQY1PXbipWSUl0UrOGtv8MEDd1AawsjFU2
fJiwqIq0vTd6ebsgpRDUYiC24FUZBfk0/bswRvitXDYINq3TZ2IAVc6DZnB6B3n3GEy7yxHEWi/j
TBjQRQXQsKmS5yEVrHr+sIrG90wv8fgG6DNJBCyzL7ej1Pu2fzPu0abzc4N6W9OHuYAuCPs9mxe8
bF5G9H7Jj03eYvsRr7tRKUinkUbaKc+soh81/Fl2zi1gpreZXzbivufqq9P35u3wNZdk6AkEYrKC
W+AUkT4lcYr2YsJu/LOjpRedUzZJ0khNwITrmv0vvQkEVVy8vtx1zjzGrbUzPPpoOAZN2SYI3/u2
Xh3s+j8lx1QK6S14R1xQGrrkuj10e84AjoT+p4yxLFOCAg8+RZlzo1ODegfpV91jmhFqwW/g0Cbg
ZlTo5dLZeC6FhsZb75RtfnD21Gza1jXxG6yfaXTRIqFX2XYCymwnmkdffttCPsIs9v3ysjP/9jg8
cvvzqpyfRSvBUQbCBAhIAQ3Sp/6oflW9QVclu6d/c8c9sw0MtcsIUxmKnX+xMOS/kVTizpR1fRfp
OKqQ6iVLNx/3nz9J6ly8uI67LJL6EmVM5OBBKKZ+8zl44ZLcE8crMg+COKphIw70WobxRLoX5Kva
ub7iBStNn1Pn5dMnYzMgOhMFe5qLun2DlcURJIQkG8ow5k7kXBPbqae3tmqj2hmJ998+NvEMjbPY
wnUjtRpjOh6OnqQXe9n/4sXu3as1svTPi13K12zknUaSJLKvcAZh7wZ50jtuWi0RD1MqBtQe+F3d
hI+AV1wZVrlJAEYHEutIvffey3vdEctUJxj/m5tpheIfmJQybfYv0zK4FpyIk5Wu/O5cPWwRz4/m
EYl4wlZxmOWZZidbSO6SrCtme8N77JKpPW97YdTirGnO4fY8J0cZ/tXLzNUib79LNA1p2YsM0Rhj
rVltjr6oUvDiRq63+6wRycIx6En3QfUZX9dqUrp+U02BkGTJmLgktz/VmJVA4JhGaD12bKZ4VZCb
jDp2y3aC1zSVmZUYgk4KKe8xjeseYg0FXMr7ygyDUbW2Ry2F5ulRsAEOVU4gHgZmLddTYe4385Ik
Q9mxVSfqb+UCF6C86wqQ+VyPehc0kQUyfgVRqieL4qgrL59abc/C07RNqEj+bLeOm3N79D5VLmJt
JXOMhE/eFf8GZ/HJ7SNKHpeoWLMJG2U5cKX/j8iYdIDv0p7/FYQywhoTl3cXNG8VVTMEoxWfoMTo
kdv26zxWZrvfDKZoTCx/Wpdd5arAfadzjW6J3PtNsM3narejrVz91v73pHNxphMsxYLeycaTr7fX
BqRQwaS0j6tqeq3s8Z/BEWxnxEknhnBY0V/VRrRtZ0G/JJlUZLNAwai7pVWk4K1GtWhgi59LCqO0
4h6w2jJSJpj58dl6eO6g2DV4nEMc4bqFGZnLKzNkLSKvxEmfFAHViw5vG6jOLCpXcWLjNXAtkmTR
et92F8wHvfbVmlNsjU/H7exxEcVng91KBeJPRhLknxQmDaDPhkmTVTMFWudj0EYrPU112wY9UiB7
aGaoIZuKdj6HgVSGrO7g9HPh2Qy72uJ3DjS8RaT+w9Da2TnZiIFpcfNcflYEioBIxBjFFkT9qQPF
wjz51W80tfF4CoA7FFRNKZuOFiE3fYX5auZAf9vaGUQstRNzONDQEDIH4QrIP8KJPFS57JFHQJfv
6yk/X5duDksFzHNfAE2S5FqGpN5bsPALucXXhfFVd4Yv3WciW66d6v4JjlIYHSn5wvpxXpuZPxHB
2HR8Idwc9VpKmMTEnZqerXRO51lhw1oRc43nu8ZpDFDo1kA4l6shJHWjgN1dyD3p1tOup4nRaxvW
9g4x28Y37rk2D5wZKgf/uvn/cpSs7BPTXbSo/Y+kuiTZ6n2M/pTO17aPHkGkttrNVJyDqOY6+1OT
SZtrj5yt/XNarcuBlxXwpEmF1BAWy341hiIHeLkFyFyDCks4M/Ef0s/50bSV2rtP3e8O+hOhnaK/
PWnuSn2CegHaYqglVul6K1lkpobEk2AF5qN4BF4l0yuoxTQEovHS94BtNuZ+b9vk3UhKS1mf0shx
NzsAYiQTChUIidBx2VwfD6uFCBlqODhUFGJg29Y+azmgw1Uv1gX1VFXHh98wj6hi60TMKxQu9HFE
2hV91J2gJkyn6wDDTXZaxIGAUYkTs5GpLo2ewP6Tm2tYhGMCECmLLIvEy7v/v7lTUYBmU5Sfow/P
DSDgZFCZDvXEd5c7YBsSo+VH71HlkNJkXxl6jHASRWTBtZQAL2Z7Q7eW0dpiJT/CcfGXPi1PlxSx
9qCkRiloA1I4avgQlpwsMyts3bN9nTczM+FdO5heOHdwHjZ+DxsH05cMmEZnC9hahbrWq4ZlczyV
9M3kFqgQSLO17/o/ShYc3slFOW52ApJ7a3a5kk7DVYaHirVAFK7AVs++36s1UtO0yY9pP4ixK/yl
jPOLupDgVyL2GmRc+rGLLBVqL0A2fRqcmgNVu/eScKu8I2AA9kKR228rtuAUHNLU5rTmvs4ETEpI
l/3IMl3V4f01tWUUNcoOtcywvKkFKjSZdjlR4tmHHKt07J0xFZwyJqAK8pW9j1Kn1dNhqtactwWH
Ra8veL4rp50qvRHhmuRYUmmHH5iqEP500spi+TUtv4eVnNS94qqaPY+QRYhzWCOIqIh5sAjemAAS
t5syXB5SJd28ti3Ktw9O5MmCmad/8V8JAh2QCEPZH7QLIuYjaePpYH+/B6uAF3+YVabDBunfUhkj
yiJOV8Jkk8CNOdSAjj0u7SdbscyZQsnaUjqfo1maIsRlEeqrq5cveEUgUpbQAN/wkguMV+53RE1K
8bgQdg0IVYcEHPR2qhOSiqHWdzMyV73ico0svBdG/6vV8se2nMVfDHlfmxnrwOqTSHww2s7pJUNi
xIgzdCrRR6ZovMU1BiazvGULTcsR4IMBhcS/GfTpomUPyfWqmHF2vEDX3LoltPDCTjQ8B7wtWxh8
AH2D10OhnbM4Atv8UWrzZVD7hP2KNYeAMrK2MwA/HswqTzlW01ULGF8VRXns7Gp6uBK8uL+0lbsa
fmPKKElbduPK/IZ21CnCTx1QgzPfjrDeUF5rKTGHc0ID8ttQA/TIVj6BjEdb2G0XjSWi0h3PEOhb
OVDwFcaX9DjqfNGkJMikSt+83X/6b0bK/hKFvdN/WB6O4VHfdGGGGNypmf+a8jtgTmfOsq5qgqAH
9fzXHxtLgt0cr+r3wQ0iUQMzUqSfJydFp/mEuoyn2JJAMFkZI2XAVCGExEvQmhO+uV18i7eaXhHu
E4JqcXTydpRSHVpciaNAD3ETg7dqb2xkj3PS9nZpwUPOo73kTVSHwZyQ5YuJFvMTEMb9LCLseJzK
ylpa4rSrDER77n3nnTrWhyOj+ywSkmnZ7rVRmJt1TbP8hvSuH8EokYJxzRTbRapvVma4zM8NDgRL
mlZ67EGnimwl5Q3sO1pE5EVh5oPphwUvXvQUMiQF6zBsLNzc7LPJXmzpMO3kOukRgkc2oKeW9I+C
Yue0JCvmVRkUg/Thyb1VN7rG8Kj7mbobIcthEShtr6h2PQbBSoSn3lH8/oVpU1ScNNyMMAor0dG1
aHN5JmWeRuKUh+kQVlt7LnuGbfiydVh/sI8G1fMHY223Nl5Is/F8/LaKBMOIARzyzWzwXa7gYOk4
q72nIfIQ55POcyftt8XJFvrfqsGoTpH8J4Me48EffDbPQUqfgeF5dbAwnXBucl3RgVam1KGWmkq8
fvnzI5FAHY6nAVOVYGmsJewM11Xpx5QqmcIT6bESWHE2FyVoHycy4W4YXzOzHeutSbhId+TBWE9+
8SG+yrPDbA+mh51FFZ7Mve3Lz/idyY/qX69iF2EYDaiW5E48xaH2ZezjPSOdzz8H+vXcMjl0dlCv
ftEAULF0pmvHh7XKpVFi4z7uLwOUiuIrxByXPAN1V4iOqxr89yi0+WLYkPTKK2i0qSUkdjxdDawW
DCL76WEgW5clr+nkDviZf1e0hjxAyZzNpVbOBSvhiezhcEqa3n5RyzedgwyJnio3VgdMd+hKko5s
0d5u+eqNEgqs6QavvAyTQrUr1Q8u2QfecMMnvy2rrKoTHMq6sHPFtRKMsXsjQ9F6OhP1iO8Uu5J3
Jbny0kdtT5TPA/HZIv/wYFeoXJEiosb097JWgFIoz5QSN60bIxvCB3SftWusbTEqitngDVYctAnw
DRd8AXM+goKmzEqzihFXtS4QrWXLhuFIkE3ZH/aAwuwIQlGFQYEz2b9y9fMyv4xUriWMDL3HGt7x
6Qe9bo1CgVkT6PxMp+dpUoglYuDlhCZLgN9LRZU/yT0yIjGXLp/MK5GgpVER8nih+Jmw5pMhvnFC
IugS/LGLI7rmWFyy/TcJwKkU+yYXAdJPbV2Hm91TMiTIBe9hVJM5m2y+YjX2nRPJweMaS38IANQQ
/HBAWB12Hvw8WPp17Aoh/4mDLdxJoUlgymJ3iyoQdhkdIy0rGiqRzoTUsBOLSfqLE3bUFoDJ8jvE
U9bgHyPHMrD5P0ZlCwB4wjmgOOk63f89C1eYcZYEfjX6cA0wVkgu2RufvumROR7T5fefxvwsf1nI
pK4xAZkcmKO2F5Z6mlEdplkUmwxXMpmI2lm/plsmnGXCjVSpXDGNcVA/csV6pzTtRPH2JJegLJqq
AOdv6BqkoOF0yZqLKouKQP+20aevry/aaKwcRW+NkMWhIewA2oXMJEfb2aIfiMJsXLArXU5df8tH
ox3JY0MAwJ0LqKXDv6QlEDibc6dJmrpfm58AI3lkWhmybrt73pEYTxogJdkYHxxYGe55h8YylqH1
jZOG0g1+ZynHo8rOR1Ft4Kq2II77tOcCINZRRYcXLkRt2YnvMsijen9s4/0CKeF+7t09mLRqNuf5
+blQt567CLxKQl9bmihNiLXSguK6ZXV2TCz+7xQMhabPuWA8rpMkCNb2DXllZG39/xRdbnFJO9NQ
1ocTp+ihWSRMDnmrB/NJgF2B8TPBWTEkbwUr+8GalgwWDJ51AKzmx+3sflK8xCb3hF/pV3HCtB+R
u4zSgD/9Z+yd79yFCp6d4DXZq9ATG78penfhKG3kIAjGlgYwgu6f/48bUt5LW6iHNGqa6Yc+eknM
Y1caPrg3734fZ/Ht+1pMM1+63VomVaMQ8pq/uuYp3/jDtTV7e6tjc4NLdsnZ+UFvGcEaZydvVEXf
MS12uDer+A0n5FkPWWWAZWtD1UWN/8dbswBP0OgidjWgPyY0KM8wdrKAI4i/U/0mG061+OuM3xQR
7tijoGCkx+0BBxFabC6D511sTmIsC9Eupf1AeYttTW/LjHQE0J3ASJeoV7RUz1Fzjx2jWi5/xooG
TdQNpQPLkaRQy1GkC78PZoskXM/c5kBdHHSzoQdvBth0Qb8OE5XgBOQaa7PwDIijXNfSNKx6WE7Y
+nTdY5kBZ0nEc+M85/bgd9QzZVaSQaNKDP6yUoU+F4oRXgdIVQ9L3tvePX0Bv+Lro9DGBuEoct6M
OPkJck4UVAuU9mibfvmyD6C930SMcOy0mP2UATOAW4Zi9c6TyruDA788KE3zaPIcf1KfG6XZywHB
Vn8bvt3InswwFtzFwFL5nT6ZauoipPLBVwO9Vxg7whaHEFRnjBVzENRrBdR2tSLuBsOtFelEf9YU
LpkxcBMRLVegiX5RrS3W5UbdbJ1hNgJ8GK0qk/O8x45CbiJbWzrxSQXVMIh4RAMwa3XWzH8eX1ai
W0dqO2oywqJlEF5zMTHuj8hy3e97GFmvp0ZOc2GnAnINTCD62MyuVIFcvA42QT+JJ4UnydjNvBKR
n7hdf+Veytl1yAwfYkBlv37YN720Rn2NlHmx8LMWqu/v6ROczWcoiRRv+TIu2snUMXecshCOlv+N
ysqnEjl1hkXoahu3y4l3o6j6y7X3WTLCL0SH61koDk0ILcHhKL1XUQk2YNI7Vb1ObIwcf0b9WjOQ
QuXaf1teZ1FkUAFWLsCfyxBc3XeVn2Be3IfXh++4iHDLkJtZm6/RstnF+AHqT4UyRpuUVn66CRfi
V+a8VcLiCURBt5jPfAdp/Z+uIl5oYpZIos7HEggWdPiI9i8SYSt1LEiMZEUKoY1bG7PGe+YX9gUY
6cy906D+5Pk5l3pQ1auKeI/SIBD4530tcU5U73ASfzqmtZrZKV5UeS+tKVSKD4KaTqITCCnD8QDZ
GQijbiYLFzF1fjkSxlWR3x0yK93OfEiT9Iu+ClzdcG6gXEkSiGPZ2QXpuX1AhSvBJpm3WBr3aTh7
9Jd9lvHS+FQYUqwpa+iGqhUvzjFhPUsL+ddkEt+IGi7vxR58w/wyRCoqZavJ63FEL4wfFgasQkUe
/grYrvRdVxoIhVm49qez4fqrZw6sFWW1+B3V1F8tiGuEaDi4QWaYRcAgZLw0lUlCYebUOXo1z5Zo
Oo+uE08IBf3Vqvk4bSLm94cvR+SZkxo+Fz8zazHgpXxWIZl+d24Gk/r0X80rYsGapARLnouCFHrZ
ipWnN8eMu7uH9/QhZHHqwI7lnHq3Ls729ve040L9Be5M+loAg2a9azNMWttOkm5ZxOVXzLOfcLbJ
IYfdngrWVC0cUrdKTepVMCcIa3cI4HlrXutwlKH4uIWK02DE86fROe4Ttlhw+IQ3HbTFeB/aLf6l
kax23jC46DyJKKvPWvMGvt65UuY4It6QU7h554h3SOOs9SjQBllrWBzZUoB22ptPpI8bxrbdWgtZ
XdNXBcczPE9m9gCqXjILpcrp7KgB0XUsaPDVJhmjriRiPQ/9TxC5kzkjFER6k93d3mKoJa8bh2Fb
nA7aZLHR1WPkWeCCYbQgety5ZCXMSbQhXeQTXUfULK4mGGcJ876gbwyWGw9O0bcpuUOULHRwPMS4
rn/iJMC/42PAL1wdwSy5h9tGMj9fTlwGEwbYjRFQv/N7kPmijhdphbQev6ZpEmbkqDx2Qw/iEQj+
pshhqQEVWHHHW2Q96m9exgpjIkaGZwiJ16FN3pjkCVybuD5VMmVP4/ibl1cPKZ89yWROcZyItDBO
/6woC/H9oneC5i0cCDhos+fe9sZu4fpEnvCWMoq2IA5XlUh4DDhOXDxt2YzaUXGM8SmdqtFMZRet
FoGsIc9EZyy/v9TVxy1C3Xd+itGkNisAWwwy5BZpcfLK/Raik65xDc79FOhlgtiXrO9aFMuAxytw
6xFZOl+RE8ylsxU44LfSyLAVuaQbKjeOe4seEnEqhvdq3lvx/b+AF8U6EhrB2jF/2bxgvRZUyIu9
o+wHla082TtLspYI/kbYqpEra+hlQ2+WIYjzrMntivbFQmcmFoezsnJxdXXz6VLBQSizIs3X3myM
lgpDiEs1U4j5/ywSocQr09xODhjICog1qus6yniLYx1N52LCUWnIfnm8ACEe8ZBsgvM6Vgg8QV5K
soYZmuHrxrJR9BHTL53z8J+pSAP79HzIxln6xo+9ju6TQrKBItZyKw02QbVK4vdgFdMKg6UrW3Dn
qP6gd3un5DdhRjoNRqkhSNM9I9T6gsEvLUDfHziqvLmHhnRPF4RPL2O/yX4JTHWHA8xMzLNzDD8M
gvgF0HNXlK53CVR+Rvdn6uH62jsWntdA5O80baDYzdgajv1FQoIL8y/RqcUycG3jsl4huGFeHadF
Ntdm+vj7Uwz8zHVainpQatpkUpRovDANwSWBgro1Q5OIqGNQTJTxfOFl0qwTsveyYw6c+iw2TDCi
pAvoDYobQ4AxySk7B9dE7uqPk3GSK4q7Y1TOqmr8YdABPi1SJmOUigPQzZaBbqun7ZySGjizn+5K
1Z+XFO4WSBWjWtxtJW8D9AGcqSch2CdwhjUqLNRRjw+w5Kd1J1eAcZfgdtEOLSn6f5qEpx21nyPD
MAJ5MzJiuw88r2a7+xvGtjDeQ/XSblVd0Qxucj5bWJgKCzlBoUx9gxv6NOkh8oWzmVRtq4AQA5uA
e2hiAfa+oPV3KrV9E2jGkgp8TGEGyth2uCBQGtWT04JdFMB4xlUYPCZJ0/nwFpk8GbicYc+MWnnl
lU3Xdqv1du4uOQM6n//idxnk/6VYJpwrIpqwTpwQQkzie4Z2nOlJx6xXttL5eqvpakcNKj4mEgLe
WGvm6aYDBbh61/zJVJhKpJ7QIkvp2Z5InOLym2EqGJq9Mryu7GNe10u9jeLZF/2EdApV57LH8zhO
B/NiW5ZyEQqe1oIsWAltJ4M6znKtlCCMDBzVlsmSPCXcr4AUHq8dNyriNTfzO8Yv/OQxqg+yKfE4
v9UIeEFeQRsL8OYNu+ZzueuHY4e8JOE79bNrA9/8x0UCfo5qH8LEezs0NpqcEWNX1FcqpTlNzyhA
aMYHMFwIoTUTzfoEF6B8BfOXp7kthfl0D3nl38xrY5oPff9jmSoo96280l8fFF7SdvGw8HJLMFAm
yV1yodQ571M5kTLpsheKEml+niyLv/ivXJWSZfxgU22DPgv31RfeuYTnSCDA5gjW5UbxVCbW4VeS
zR0BGn62cvPrZnp+KQqrOr5FmuJaVnG/WQQpWDYunBhezktRMM0U9+BA/mJbtqu7Uc5AQwtc7VTl
GbPDOtgKn1tEv23d4mt7lPDtQ1H+KiJ0WNqfrxLrSabB0Uj6xCqdyXF3VR6CTuz4wTjgJ11xC8us
/TM5AalkzU968yaekR75SaTa8MGjJecJvkhDUyXWkTuh1GXlAe1X65Kx/lmq4XVPKbOx1mHKi4sL
/59c+2I62I/8NvxihmT1tgUp06YdeqjtCpoIjye1b1oq+YU/C+T45YEKY7X3V68TDBcTvzRaPjOa
6GDdIN+BHXBT+jNE5EHL/08Dh+m27gWnsgaIghPVDF6y3AGoGmM3llY2uRT73CwAHaH+OGZDCjDF
A5F4EA4tGCXC7iX7h3lggK0txfS06BQwZr8zjQkpwCWnbKHdjkZOcE/7x5Q/kefd2ugu7T+j8Iiw
4KHrmqqQlYdwXER1HnVtgUoBC/syGNkBfSzBP0/9eUpdteaTe+lrJByzeW4pW4cEJ9K5NpZO6gAd
fVVibrNSo5YJ8rSlQTHipbySMADMIBHNbY8YLMJQ4nCpzeAfHa6BVS09ENndkmXu8IyARBhhW+h9
9VLI8yxSrzylOyMIq/krvwFyfMLBg5BTzdo1t25vmOEfzcQ3oj7x6H2+mmKHIyq3DXBwRbyWLAI2
e8d5E0ixt2Orfi3g08LKt+0kwIKs1jmgRop3/0VrDxXLwX+Cu1ihDxF9ocIUKpkN9GIU95gAAfcs
q0WSMHf4eUKBRSIlywdFPUo/8ovzlbN437rzsRZp8eAXbOWgRHYWPzuGPMSnjwdp6A7Zi/lhQUln
ZUvu0S92+HNN8R6MJtkDGObmcP8bB9et1VkTv8fONxjqT0DVqdMVaceSfMDUDD19yh5mAibijB8v
ri3TzZvFzPPrCSbE8ThxrzyfjywVr7Vs9TpQJ4K9nJpGruO8TNVMjouwVLobxvNJic8gMm4Q3tt0
+CwQVSMIrbhRzdLInOT8i+7QsRzq0qF7NFKCXo3i1SNTy0xnzedDLZSfiGDsC14h56RTM6T8IfGd
o0poM2xRk+7QnmM8fvsZ/Yc2jgmazTbzQCEwOv9eV7+QUc4E48SxgFcPeQLs5BXk0CbQZUJo1A61
DVYLmauoU7xbQPmo31/znKl07z/SiqLtN4T8PswBhiYT75milnxphGewfMRcAUX8fljMdWvT9MU0
ZRaNVkmpn2iGhjPlMolhNkTKzKVpIsLBkP/PhLo9WUuSvJf1kmYYbEAxvzcicm5m1kr2Xte+iimI
GxjMeIcC21JOxuu82WaNa2GwMimuW26qqyz6k2eo0KPVFI2FuZmw/S4GIIfu2/DLWwRxmCmf8XXI
RY/dETKl5D0VRopXLCQ2CNOWp30hyDnbIXJNZociotXHDLA6MxuLc4nEyoFxq4UihqMntouiLjvx
TdNMb24JQ+jxxUz1Vi1XP+nEjo+RxyYRmFs/cEM4GCRhRORAxuRE3zdBv7Ir7QQ0+zshv0CCFVUR
a3+610iQhdcVRiHDYhSDFdATwKFpv7qpWsQpFcr/jlmDiWQfUcgBybxXkWXOZjOHJVKFEUsAy2Q9
FiipSm+sXs6eZObTj36AB8B27kdbLxVLhxPH1SmDFJQnZEYiugDeNVpv4Gt6DZDx3XeFPG9l9bTb
Dq1jDrDJcGL0EaHRRg3kpi3R3jYVSn8MayMAUySrVtsCzBEN7KWT6jW3+upEvFPZATfD3K9UMZCW
ZAKU7ac2AE5YdGuXd83YZq5oJVuoYnhEvileoAVhhr+ft+fnRrJPjWV5/I53rg5kBIPRREI3AIJn
CZ8BUe2ihaxboPGse7YKO4H5MmZ7kAyYNBfwmLoDWtB8FnjgxJ4MdCzz5wCLq8rw8966fv2GAvEn
z5g08UcmIRtAfttevdznY9QUeRU89kockV4B6MTy/TheAw9zuix12nKRwuJwSOA6kfxOBU2GOQ0x
PHxEd4QdHvxvd90PoFPuUX8riHRo9OtEoMWCG/tRrJtpIqyeXLSRP9TigrMEb97ZVStYLogWY+yP
y009pBS4US0mczWz7kqDrGnnjZikoaVSyH0tqfVZTfhiFvvpL+MzMehFyxGjB+LByGtMjBNVhRrx
zmo1ZoJc63NahGEJ5IIxYnXIh9GrMwkCHytFKY3LwzDpTzAHbT8qbYtc9a+NheVsaNKclRxPcSd/
TrOA1X4mS5QLbHTztm+OfVX5ZTpnCDfxdr/c3WKzW9S6bkRsZvISVwcvMhKCp9eLCNXQXcZEu5Os
jWsYxZ1j2/ZQMrMfgF9B4JvP6H/WQcGSgBMJgraefIVBdG+aIVJN97SUCV57ITShlo7W3W0+3cH9
m7oKzaqHbITOozpKj87jwIsKFLcAN05VRA9KrNU4tiD9B6hZiTvNdEh6uukLzfiLrm9Mu+8ve1K1
9radql6s8A2BGVtgHmIWHHwwN+cTukj9vibYY6CqUmI9ZzL9Zj4Cb2VLVhGYiaTDGJNEe7cpZ8f1
s4ryCirWvk9nkyhIJ7VGq3R0cnveMNX3qoC+v4a2rGBMQ+ZVjzDVPAaPOX2RIc2wuVJPGxrhC2yp
398WXG93kebk9uslIkiBEeu2wxaqZatHpd1iP3ir7FSGYv3/hy9abDGhmnB4gsm4UXNRa6ERK3D3
+RzVg6AXpSyBdI0LYna+gOUJMoYdASO6TOUTsYlfKcF4CXfoLqxeP+Y24PXXCoB9UAauwkH12fJz
5zEkmmtvQLg/+p9t9l1Vqb8A0VIzBB6uYQW4U3q7BW0mFdh02tBYjoxOj4gyMrABQOww6cOUmd8B
Loh9YVN6XxOiLLPMJC8DWhaj2+am0itu+q/mOof7y+Fc12MKO1Ds9pyxKPQdZTcWTAJR3flxkmAK
RgenhQIZFXncb9730Bmoh3b5biWGm/B3S7/k2TvOHrsR54F08X7MHhWZbussnhZwmSvUfd2dBaa3
SwsJecRM+my3szkYkT8+tjS8/ujRhZmkXuRqjmuK0pILHBAZAGiqc08wyq8TeEujVHLG/sZa543z
tcbI3GIur7Sk9UFVCrIi2xzqg9vqhbcmKWKXWqSDQJvB8E8AxxX5lkKinvQoI5pqPvRouyWzC0ij
Tp6/vnXUeQPF5TNA/MpNj41nd1SXXdjr0ZZrj1w7WsMMp+rcdw3SXJUu3Qm2f8ek/IiMrFEvLVgi
VCxDYL55LR1hwRBiyMggroIiw2mniSA3ic9gbDrI7Z03DaTfS1mZ0muowGPWP1oEKcDg+Zkk1Veg
eDGmGUfGPhbz+1J14odhwBKAVkgA2/iexgZ0oJC36ruDw6wc3aUjM4eXV19n023uY16tvXHu5Yg/
Qg4jJB9UVP1ymNTZt8m0QK68KieT1Srsakgi24LSLkkuFMHMb47mRgITNIpEIBJY7io0dTZGeq4d
VL8nTtp6qf7vLbqFh5IzaX2dDFLnEWzo1s3E7kJcuVW34ZCo1yNGNQQiWqRiB91jWkHA+daBbNKU
NJ+iY6hye/GKbPl5HXQ1U7RIS4mabKlREyq7nhkgDk5abpHYuKh0GxLW0eQV6SjOIH5thYSBAOkS
CStt6GsDMSXFacfLg2v+Lv7/JPRWEVLMNP9FNE1Oa/f95iO9WnFWkE/Wu51qn5UwVUCtmT9O/JsY
87AeUlaBLDTGUFW+jt27bLOoWgW2FBpHmP5aUOJgejwxzJ7uQbD0Yx+T85tN8RP5+u19q65zJNJz
1wVouwJSrDXbWXsVB7NHAcGFM5QRJ1QeHKJo3vA/MAiyQZdT/TC4jtvLGpoGbv9MHw96NRi2lvb0
w7cx/Y8+PuMjz/sifs+Gt8edcZRGxuJruhHa/r+cjfIDQCCIBvx5PmfFfsAl5kkTZIZ5ePsCxwDQ
5A/YKLAMNDKOANJ/e0I35WYR7dOXi2cr3QP/ET7XOon3hiYf315+DkBmXz51sG9d8J5sOGwhtHB4
s8q6AUQk0KCg3SiV2zdSsY4MbcZAb6g2s82GFpCccgy/zy5c+ngKW1SwhjyFKzU26oF9J6XAvNLu
qj38M5bpjQcZ8l9o71k7rCDl/KYvP1kxt/DAJ879uOtxIqcKRGGuUbMdToH2UCd5CJ+eJl/KFilH
I51gxeyo44LcgTm0xx1z9hHeVcpXK2o7Cyka8VvpVDjzpGnJBOXmdKKpfRmCkdAKTCk9EuDycYAu
SHssR/DiAlsgRBl4y9xDDfQCiIyxf6VnpgPNwDw1JW6nvJXHaTmcs8hdi9zFP/nxIKlaTi/70SYN
t9GZZiLEllqrVIkpPReZ9ViN9NqDIblxVaWfdyiPXqxpqm/nxspmWSQvjqcDuR9lEv0U9p1Rx8Mi
atMRdlBvLUjzkuhhG0E3ITiWs0E6dBn3LeQDi6ADdwjGtcCpPYOhF2heUKBWC4wFiG3LzbUbUeqL
mYOoyQERXrJfBcOo4oftEwSylviFJe+lze3hXK3chOnMf4AzpJ4O8uwqC+vx3kZLXY4tcVjAoi5k
fzgEpDL3DFMS4kMQyhBKKxjdTL/caH0rA+Iwz+RoiWIMm4eM9Sg1JUng1io5eDvTpyvQY2rnFyuK
E4JmR1c36AoBtk1nIwXqyik2kfRnC3HmyiVs6PyEAPwKc4LRHMxfTIWKDa1P07HxMHvSya1li1pa
TNtlcf+DFSO/ideq4gg4RJ8TUrfvPF4PRO7fFO0V1DOa2N35O1FjB1GIFEX1yFUKrVpyw1HOLUYe
W7b+B6Jl1SOGxRIpm04oT1WDcGOBdypzTgYJU2K9mC3wdkh8mvJLhj+tAwV0a0/Wxw8ngqvUMfHF
dOMhYNYFr1t5YlrVfOxqjm88Lkhz5rTyZbJukD8k6IAjOi3BFp8lHoufE8N6TPmGNB8w84ef5v4S
7zHv5Z094foGYWjaZjsPQvydKLrLFLmC98Lrcqp+j8qDbPx2+Ezx+AmwQaqnD+wHgtY2xUEqfxj/
VCs2vMqWJEUGzDENJgzMQ8kz+pOoo8fgsQnJ5IZubPNEQ4jJkU56UQRB+b5wdSPqSXLTfQjswoBg
7yJt2xPIFkZHihduC36mZrTmqZD8Nd+MfLYXTA4AlMnFZNhyHYkvCJPTY25TxKA/kJZx4bBFG9r1
TM9J9j08d6MOjrkg9pCHqjMNJIJngwr6TC1aaYRUbSewpP6xOG+pRyuK9IAXSCg61xs7YrCjR+uI
jbyoitZMxNWv7ctNBYjVljMDF8XKUVD3SpVcC7QWil1V1HUH3uF0tyZ4ZOiD+KY50XMWVHzqTPMq
D+34thfg97MaR9eGXjAYn+zHhOKF7YE2B2P8h64BWiyxyqaTt/BTXuiQQEDAnOzPorYd4hl29jQA
DizLm5BcwTcoWchgCu9G7CSdO9LRncwZa2FW03fZI6ftVe4agNCCCflNVdvkSktvBCYKeWIKml50
Uc71lVf1qPU7/MD/kY89V8Z6BplqqsdVX7Ydl1v30YuwIsTfaEzE9rbXpUcPZrEJk0vmiGVqNAgQ
/JVDAJVGxSb/+GszlNcuUrvJCYNbgrgqfjvqICnTMTWKU8q/R2BNhFVMIZFBf9GIHq7laHyIW2RW
+5PuMLBy5WPuN8ZAGuxqWMsfv/weVwJhIEU/ndLBXQJlY+3Mfr4gTkLmL8e4x4nV2fX0JgCyVWk4
5rhOMUwZKOEYb+TgUbgXMJetPt16FDKQ3mh+d7oGjxD2pa8XM7vMswghM5TVYL5L9IV/1GZ+uFuf
ZSKlQmBriAUhGYmLPBHW4NdzGYf2F5YIDfgeTU453iio9/TZrAXfCTB0QQjt0fJzCdvep2HKqR9C
iFmts7E+P8fEaIfAJALQ/1xufrmA3Ofpb3/a67qK9zn7kjilrREBypE/Nlw37amV395HZFZXvTAh
Vujifqgi8xuahA+s5KwvNH1sz2Ilq5xF0lhPZ1nAcUW/OpxI0OZq+/gIv93mY5mlP7tQ0yH1IZIL
Od7SJoj//QvEFLd+nT9VIf59jtPBSsZM5P+CZd3HNXI2ZIzyswPsne/h4BpGEXjQqqPMmgTrnPjK
L6iW740kqgimF6mZ5hIcDj6vPxRQ4BwiLQrZOa9QWoNaDBNk942KDw7/wuqW687bK21w2JuAAEBJ
/skCa8oQotgVgXr9rUCgP51UbGLUCQXREKaSsbcP4NjFhtJ657iYREUpObre/UZtOHexcOpDW8M4
1vmXZTL4F1VoqxUFnPs/oFfOTwMHgaDp+tDxzKLsP5qCI83QCa+YY2bK1xo0U66EaVJT5AWnQmB3
YGxo61Bsq8oXET9CcfryG5Ufgw9WIhYgshMgWf7R6bYcQ6jYBp7q2VXGO2lK9HZvy1PZ5l8q7Zaz
xMsvuBEpPSk6AEPBa9YQPjy2chikyyclIL3HCEyR4oDTYG7YDzWMERjZyK05B9OdOxXBQDelsCkO
tqc7wVoHASepkN3S/iSLk+6koyFZ6rbdP59d0RsMfMZiDr/6uaF7qRxMyJaV6/43QlMwKO+ASe8M
fuY4BysSjJRKTEsaEd6FKapngnVO8HhEQ4K/qFOUSUMHLviY3W6af7BWalF8/FYilA/3D76bukIC
T0QueOW8tP7KA9ffRBxKqL7mamJaiQ00qlitUn6PFrWKVARZppF1wo9IUbd68Fk1Fgz8xXM5ySt1
2ncI5dOSEnm40cK8KjQImGVa56LBSz134Ot/U2snzdLMXCclu2ZBo5OnXUDN9OUL2JdHE88JE/u7
wxnZjkcNFEHeU0jZ868lqUHwhOkKRUN1TPfV3SPoS/TDEveDftXRy7UMrjju7g2iTT/2/bEYZsjU
tLntqpkXUwApH2gwDHF9OD4OtLlUqG5hbjKwd0jdsy/+fZT7kPSFQTmlWgJWUzXQcazhsIitrzvc
hl768HmAXS/yA5L+3fJ9DXGHR8ECiHIaobbtrDBCHswVTOr6Z3itZzCzKcT4tuRkaRB07vZgNPgM
sauAxQeRuIzueU2GGaB2WLcNW9BEucO6YE/LcVzkAvLOXPfqmiRIdCzYgXefLwSUtBzLYM7ICm/i
Jj6y+/t2k0hB12t/Q+z+gdq2zZdAIE8BxnGD2n/ycltqzH6J/FXSXgStrcYWFP7HvoKaH8NFDq2D
HJQz1uuG+wLKJpMbdy08db8bL0cIxWw6FeKORqEQWPEGLBPCaGt0J31gGLFCLrH+ozvgrA7FuEwI
YVDPI2DwGN7nuXBk9esnjwgkw0pIlDTHwr8Fp1T5coH76a7e2jpskHfaRMcUTR4hrklg60ZupS14
gdDFb9SlaIXXcXvO8eu7zlZQ9NHdpr1xUi3ZusFV29YL7DzIPbgeoWtJ/YKG7NUgPCGoOGRzXU2W
e0HTC4jUcltK42Yj6L9JZ8EYGvkq05I8p1vVpGfttWcw8/MFvX5zld4UfAmquCKuyWC7KreN7Bac
3vOEHChxEpWI+gNo44e4wCVqlgV4q+aCuPvaFXUCLUYcSEnGc8wj+Xy1IUv1BIUapGakI1NPZixn
wxfhtVR7S6Egduu4UOEax8N1B6SkjW+/7jHK1gowi7bKvP5K2wKdX5nTW6SumdVVTWwvZG5fefNw
08oweeVp5zgNnv6OJy3kA0bsbBsVnKNWzZRCol0dy6y+6RT0lT03Pk+J4p99XnMXHH/FS3qj8wL1
pTvveiPisYw2P0utXsQ3KLtIfo0kx4Q4tbmQW+jjP/i6gxas4klDhtI9HKLEDODMHV8KekS+mmAS
9PrmbPMC59yuTwGgaFU1HGtBxXWkT8WMRhlsyQFhGxxX+QXLhnj3VuBuPZt2sts7n5Fx5y+uGEnm
TZyVJHk3xDsDILIMgNCktxDUYPu0RDeVSB+HQ409jrcnCvfRE68cCzEJgrJipD2U/mPqOLvdslqk
vbT4A0Wdlz72rA/FSagYYYLfhMNpFHVRsVNJpPgUVXEs2ja0HgmPlRzJ2xEjXBl2vSGpRIqzYzXR
QVZ8rrtNncN+uVhIihDsFIAPS1AdQZR41blJ/QO49NBz3FckGWOHYe557j5PaMxP7vCT8lzV0G6Y
pAFC1bGx67I9PiIskZTEfcVjQYySF+ziLgDM/f1cs6zue+xDhorExM3yJKSAWC/FQNeOF7+Ohmwu
WO74oQ/bNkEt6+d+9GdqtqLLKrHw4jd6p/O3P0tvVWOWPPjXc/EBH4qh71rBC5l5wBRpVWZwZQfr
Y7bl0cxGFScUTYONLCRUs6wRrc4N7NjlqkfgY+TUMS9hCv2npDpCnEZcY12zv8oP3oe8FVshoKYp
Q6Hi3zbTbDW1ZXPgXVpm3HjKMhkj+IIZQ8ZjOBD9MkeRjpYEYEzQLMEt7OF7BbrfJTMQu9edxIoL
vnypZlzD67ijuFM1EBkIFmnXU/VjmxfndqcrdiYflRXfk6EkYmruTQvwjaw8RrGiI327ueimwrsx
IZzOEFjGPzk9EAiI47P9g5zspZWOF9g++p2cG5e2yx09t8cgruuJz/A8XEWevdWRaExZUB9BPbkp
Uj5fCdECftSDoC1Ovn1bekEPaF28xEiAEQRK2ldJYe2vG5CTLX6A8I5yGvpRyGHEdZFiMtw1azUQ
vqxJyopHk2zY/onh6uR+hwp7ntndOfb4qsfXdC6Vhcmtq2nKa57g+l0C0hxZ/mJLAxU6sCYwlx1l
X2s1SnMXTUirxoJq/JOcE17ofd+KD1lI9nkXza7e3N3nALCB1i/RXclr/2HCE9+0mmH/7SvATP7x
j06+Mn0Qzuf8Vn0wyMxK+vTGPXN+Cu2yE0b+RnO4Bb5U/29QYXEGmWe6K2qCLpf/e9dpqyzougoo
7I10Eq8if1gzeMIfENnlnBheV57MfhKOrLtjTGAiSW3ivHomE5vH74L16yONQglk9Ov8+QkdLtKO
+hx9yAIM7AlOMN7MEdq5alVRzTrdxtsq1YgJw+TC6CCvDi1DNzGpfTJyqAepVwj44oIFbxX8oW9x
TtcbcDhIh2+mKGbFdcLA31c3Yq1TI7V5Ytmpa9B9Q3GWGK/1DNpuLbrSQH0NE+nWxuix7TI30ctm
DrhD3IsKAqx2CDVjUgL9UbOkL80cRSQFQcxkqv32KbGxEeu7zmbkYFmeKkYhkz/UvJNzKzmyJ8eS
ZQBfzDrLO1KuQkNbMU2q5H1mMKpL3c3HkfGbPGJsEA8/THem52ogc6dvcqPvGUwiQFZ9jcjsa48n
vS8KAsTa73g7u2rjXaAUbTIv1nywCezlI9Qozi4D+WXKIxjRyNI3wcCvQ/iue8GBtvl8EFhCRI1I
uV88ye03+a24iJs8OAJ/6c70FsVgF1dB7l88zEuJXV0tNSvgJ+C+/x0sH5gONGPcFRGR1UlQAHiy
09E6B/7Lj0Dl6Tc/g3JZ8lh6KSkrhKcdEGoxgDMNWp5x4bAXa1Ne05cu4HLp9rUbKh06nmAGhMJW
VMiW/qvMScj3l4NgzA277w1DBGGUE2wlxPUhMb2YlJkMiceZ1UzGY5kTn6Hi+dU+Eg74OJkETbf2
o3/wyZ9kbNe3PL01RVakrQtYdBaAfc8d+AJ+LneJF6v8zF22zdZU08peAAwLe74MKdCcI7XaV1tO
JKVjjjJFbn/vTgzkNAmXfOs8RK51YqTluLqOu96dUTJ3EqyGrg2JHrlpsJyRrAJdSIEKeI5YELhl
stUILSBxYsgWA7rSD+hvG47EWkIxS8yiVX87TVpwzq4Z3JwfwjMGPU2T7cF0IAfYr4OI4ccZKvpD
cJz9aBQuV9DvF7mq6VyDfETHB7W0ElcTGdlC2SOBMaLJYCJ4fByqgw/32cp9F75bTfERhs+VKGW/
t0Cmcz0B9+39RVaJ08H8wQAhNW1m90TI8EIn17zNbHdk/awmhxRhjAnxlRD3FCUA+OmeUmbC78Q2
ta4uTv6+09k6re0qfIoGb6pgr6nGe+DDThXwRKuyrJSNa2KbJuPkXm0pJqBasasNJJm02wh1Xpfe
vSEeYFkhwtlyBU1Iv0PkNNs1n/P62L8JPjbZ3VSJB0+ZTQLXT4TM9yA6wxIKHE5opwEekwF0emwU
O+/hHFvRLyOtM8lzEWdjvsNQio6Hh0YUKCNKkUgpyVvK/DUs04gvF9230NcAmddOu8s2Y9SUNFEC
wp31CeZdVw2e9H4edPJf0SfcNQBJ679oFhh1cDywi2F2Mz3UPMtZzQmZQd4DfqRtFaJf6Ew6+D6s
NZ8xo1YpbnguTQ5xvLWXS2nBU7gr5o91zEP1B13AMtLCfmZkvTBf86g+AIc736/CyDCN3YIYH3ht
XsXjBQtuqaEoUovCXUNJOsOgzfIopUI5CY0kzO+DMxaE33sC616htk1+Nybc0PkLMbxrgoLvuyDR
I4C6lnDkj+PiRxaUMp0UlmJ1ooYOiChnEKNAyYD8yqkb2p4SWGV9DeZYH38ISUpwDfHAUOrOVDT9
1+YxMMGM42XAYNZqJMO2eM78sNcHikAdy8Cndd/cgCaZLfqKkm5gZJjvj/G30g/tMtMrMdIjZc4L
DqLsFof3Hszzx+WT7RJniumXnF7dE2kdN+8DPNK6p7fV0107PHuxYQF8nYCXN5Cm6jpmpVxav7az
jhrCM+SO5WUdYjC7pxVhLZDgK54ZirrlyCZFBBDM2ajYeN8VufJFq8OHB4aTMrzdby8jciGdeGv1
sHuY5nnPF4UQ30ssUDbDOLLVVzSIsVdwiT1TLWGuONvzo3I26AWNfi3kveJI6VllhAsz3U0sZQ8s
6CjcB5VvYICigmXX1PG5xLi5uZf4pQK35NHfKpr0Oe96D0ZW2237IYNN+EBbkPdaRBWFDA1eYmeH
FpnFRYNvpXEiNb6Z9YM7oIpoj3eROUdNzKlc8zuysNLpK55/2pqxquChVKyYwhmBCdlNFlYClvCb
PO0e4seBpWDXgrtNCA9S+pG1sF4uvUwmnCDkp5INiI8/C2LrQnDq7BqKIep36sG0WCTspuCZfn/v
5GzAtulVyPv6mlBZtojUi1JxJD4qjEoNNSeGAt1ORZe5ABkxZGcVdzeWynEdOdBuSzcZiEGfl7hL
JykrhrZzinhyVPhPlH8/1dE2hGWgQZ0iWOJXXmRIUY5I3+OOkOCztwpbAGs9iagMC1ccMNi3uRIv
6MGVes+Kcfp4Zv5tPDkQBdY0mAuxo4RMLslHIMlQchIUTFy5c2Xcd7f9uQ5drnvG32r35vF702UD
j6QoaArGbmWwdMGnm92iGWFx2ElZk9F2q4j1hFkQOOTTwengrz1orJdC4qYLsYm9+z0XV4z2h5e8
eLLcit+FWvK8Aqdr0L0moZxQhUgsp1ygGS/TPlbLWQKNXhyzA1jQVDFQ8SrneSFcb8HFUcDeAMsV
6TFXOfH+K9iLXEypJjA8/h5TwdTbmRjBSMP+QCnXXw5SjezjR8cWC+BTc5OOxMA5pbChiJ1O+hhP
a6WIgkJgYW5RftW0P5/POf8S8s3Vk8wZa9PpFiW/9B6r7uGTLg/Jj1hoax35aO41SX4EV87u+f1l
2otUVk1Ln+EeCj36dvQFEZMUYUKs2dWfytHgfTNkc5KmONqyyDCjmNXO957VEF5ZWVkyvsXWkjVv
26YcDwWELnlTQfGTthpQ2B5Uqjeoes6j7vCiKKZZLPjXN2OwaOEQUrK11cs8fekHqUv8sroHFftg
JthRJn5bAQjAoTXNFrF9Th3Y0Xwb85G6UnZU7CgvetwUTSTiwJ23R0xRge8JgUZK4yMHSnHTeUjn
UuQI65DllA7l1+TwBmT9IDHP6VcbyCIRi4/+kcousjc01MGWlObhsatFQeS09+YXYFeLr0fnLI7s
1vfzUTfu98vmIAAqDpxZgM2B/Es+Tr1dK4ER3fM1uycwK918yhhk01QZaFJeRzJFimJWMMm59nEG
aihHNN8qRs53c7gOuIC8wdP46F6eyFU+t/ZnDhxWKPVNrjSHpzznHRy0zvfELpA5gbFqv+hjNB5d
IZrNenS1tRzmfCXfXL4gX46vJLOyq8ZERzEy7ImPY9TXswF3h6L3XC6NMrozs0PhGbfLWfCSbPno
rpnQOtCH4kDZLgocRUSLt43t8IjXU9m39AzbqAh+rQh/KYRUNE3BpyHCaA/l5tyjQX2/RlZZCGut
U0rFIsalg5tCLl9qn1/LLnAAEgrc7xpUUyQd2367Smx7g5mpTZAtPjZknePte80pfONxp0VIOHmt
PO/l9Qk+pVUsucFVEBTtSaL4i/62C0Nnhtm/CPXFdWVrus9cGRJt9NLCnvB781U9kJzpmR2HxReQ
kHwxZARxJn4trDspRj3ouqNpgU2j1de34PAvT/Jf/VoGi33j/hCh8oCOAz8cxxemjGpzKNWAtJBr
ZbqsGGgToAxfL77NpZhy88u1ucZJuCtcx6uaNZ1A+vveOSxE48m22ZaDeUK847PjZ9nzpVsRKiBm
Fuu2CkV1kpFCxJGnIddwVScc55DIjDbPVBQKQDbEAY7V8c6kN2Rr9J6vUq1AVqshmqToXJ1zXpnc
kdnpqg8XekuwXpWBrxCwnSnpM4lPclrQc6893+HRsH/Fyq3BbbihVufgXk+Xtx7ZuzZbhh3g4MKs
8DpO6eHnLSES21pOEizayTX4ELayiTq8frXpbfEcEk5p4ohFiL0Pv9+t+ec01eppyyl+DryN7KB4
V2AhAg0r0eg2ygQzhKSLwyv8As1Yv035fF7CVOmY73/RDrCGTUsjzsVOSXeTb7yOll23ifltee5m
9lHHnZQLN97WRu6p6iQmeCCS9bUyEq8TUl7SEZVQ5EQs42PEVmQ53u4QZ1akycnqrvTrWhx25S+1
mIqRCBo8pB0akr6/UFcGIYRtxYV/qoJkkKoPad/zZEDAb7vir2r1XNWO8z5hklh739Tl+8mwIlWg
T3S7b3T5Jo4GqK8Hoq55x3X/aQadwYZb2DJUmWl+6GK4AqxBT7K8XBe0UAh6bnrpzUxJPp1RiuKO
M9YPI/GQJzvCVc617uYz2zxquVx+A9fN2HgYLuxk1nxpfPhjzyWby4rh57FgjOc/6d0RjLZHCEIQ
kexSbp2M9AFh2Z8LYma5iJuwX1FbgzCkK0O4nVRgL23UEDJA1vnuCoPvmwa+ejQX+8YEPpSPAYnf
7z/+gIY3gDN/UnWUIO1oDyy3WwKSMHAXga3+2XoqITKkHr0t/QuIIyWaTp0RCsw+GPCeLEw3TXok
xd6RbTGm8DXeKiScxR+3AEpIabMMvvZfGf57MKUOgq1ajxwlnDrEFGM7Eyp8Mjx7vMevnQbm+1oh
J04nnh3R/2ZyRkmKnhuJpMyhMPMTNrTlbeqthxfiwxH4djWTDI2DPzPtvCDzbbd2aawLROvAAsLt
YrKeJTdZ8ZpB5WLn+6Ee9vFbr87+Bi2LsXtCn9NjLNe36TTES58NXJtQFCRnt1WT7S44BwtZHaYj
3plRhPZBr6fAIQvBAqRo1zPDsZRLKrgC+pxoNDLeqztGxLPWCEv075HK86+tyxXYrBTSNzL2Gp4H
anDwX+LKajH2/yEF3OSilLRH/Se8TCVOPn8Uq4dryad5+1wwzmWL4OckP6hiBvGBoA44xRUGQwDb
0/nOjru2qevPqkLcuTf/CI5iYTJy1FBBTy0W9B5CPvur1TVYoKFKMvnBq7psWkaiS1qAzUHH+U51
JmyvVg7L8ItR3zssAc5OlZv9vKl/GCxWB3mwblHJZJg+MN00Dh1nyRUZ8UaivAVRbyZcNpeCIOaS
YUp6Xz1W/lV+CaKGbB8hopM4ism6WN+bM51zrGeke3id/16G+UNBwxxfeK2IZXUzT5prOuoZdL8b
ZmefXpFDUGN88p7sTTPT9nFYdhQH26T6ecm1C8sJzrwGHCbG4r3ELYCqSSYkTXuBsFrowc6ZFcjZ
vOPoS6XdYWHb2hxYArGBh0BiVZH0BWvmEFV4WBeZr5oyQKl94suOvq9QgDpv/Z9fQhKEW0GaPu5V
6y4nMmULPgmf0wLjBcZ+UpJggCQu7ypGcHTxmkv5GMzUOjJvAgby+KhE5K5Te9qyEg5YSDPDg/af
LuytaA84Yxir+JDxyJLftCKsl7tBU7Xq+v31YFK/EnzbQq73V4y3C6NAEm9yu6cKdY66pGygVXfi
X2XdI+XH+XtO7CBGWNGHpckImJ4D9jXn1T/UTh8HcMmUJnR8A6mzdv/kcceWq7k1pMuzJZViIZBp
YYVmnCu5hBvAt9LHDT395LTU4uxFgVJHll4tcBdQizbtYErpW7nRJU7AXYnuYXllf9425pFJUhEH
7G0R1LMtPbrwcABlQ16HpYwszpPk2Gu9Fhay29ENEOYiGHgRcEMtnp02fX1gir/eGXmcUOmJkXpz
DYlfsOKAmh+ngaxBQ+6OyZQtco0LgjUijabawWSWIGrlewaQZ91tzbMI4RbWhTubLYwpRYM3Klsc
dTW7+eTiGLjWOAxwobWbE6qndENtM4OFCKjIhBWyKGG8857fMfGUP9iVLq21kRgwjYE+wTpuGMCH
mZi/NElDrsC43e842dD6L838Uhxanx4g1V0F3UXA4NrKRm3kXhfaLljGrXlTZ4KLv/CvgkVNl3aM
OexA743WN3ihDxW8McphWcFHXCeZB1xlFxhGKKEr1sof1ztxOxLuFY0T3NQs2s8OtQWc+Qh5wTsD
7ocfNpynA5jjzxUnOjSqvCYr4CZahVvkCK45NWIrUDNVXrsWqs9wI2ikjNDOonGBwg78XVP3inGR
nGTxI3VCyX3AjjnKzg6UjGvhsTwHQ+mUVieVa7ZhUVmt5qoeYLzcPo4eIkZxBhNCSP0fI3gYUlD6
bvJC+c0zogm92RcpCOVY9AVVv6SYzr1/s9VH3sH6aRDzMW3rs+73IYlqzQzhHArKxY15MkyhPEGp
R1vpZQ7mkGcyijQKrAP1psMblJAnqGBeuUejtL+1swrH2qlEiYhN13JRR0C1tW5Bde5TPfFFN5Bm
9rMfmeK+ER+efQtiUp++rshG36rFtB+w9IBubZdPEqFJHACJhFq2IuHrxprYTLQN9sqY7qlhom4X
3pP/AG80S4vQ8nDg3UvTwYB1QudU04SPm4/nWs7Lc28Btm8fG2MRn4hLZiVZcCI1bG2//a8yebIw
Jw9rb8CqThat+lM50p2DAEoTbsASscdf/SNq0gA5/9eFsO9OWKOsSYnYWDltHik0AUyE9BGixxae
KVamUjGQudc17tNnhLzNs6Y539fcmCd2ATj5UzBiiPm3ZLI7VoX+w0hRdoPd3akPGbO/1H6ygQzi
+E4Wkmk4MqUhxkxfSDUX7nMLZvvzV3PfVFEr9NzUqpXMuVptayye/ZugjQmDuJY6YRQiuLGtlrSZ
vDbYQWGtrGp1U/fuG2wfi8CUL1sGo4Odqi5MwpppimbrrTtjakN8qSoQ5Tp94KuhkUob/+Z0ix5r
uCWOoJovHj7AdFlOY+gEWlJpP9O4eV3kzTa6Y8Ed8kJzpnIXvCSp6hrY3MYUc3DVFXUlvSxnb0yU
P879/KQ3RXWoa8VHXjNgnaYf7cOxFeHE/V6yK1MoCnq1PiCN/baL1qo2vTeQ4bIAZn548PClwRe9
zXWRy8fnXSRf+zuMBWwXWom1xcwqJksnz1BDQ+oJ/Zsfh4bEN9mCs1zpY8fOvsKVgQoBTiwHCRJj
iJoHUixlO7Pq2+k1DlUsSoccwlZPWA9fHR7h5EVTen4tU3AAI0Y5N6nZUl0S6pSkcmXAdoCFB2bJ
0ehY/Fsfdln8K0abEq4qXUL6Gre0NOszM7j5UqBSEvMqUNvDaMgtMGSd1wNRyObMdPILF1UlYPB0
a1Jbeq6/xAuMvQ3F7f8jlvmybd+8HV4FQLZmjqV0o/KxEREMX1Rmcb1IcVxNSY++R4xgULU3QUya
PhUzjsuNpqcZuDhpAavKuywGb8J/fWhkJLF/KKbsqOT2RRfnvCCxjMcRKK6jHvCMeoGGObNGIaxb
5plRFVCyvTZf6dRNuS/1/JdIwxg6fbVHcJJ0iZ41sgHpKvAFeB/qSzIH7jHwaWAmVzHrUYJb6nJh
VTtKzau8huAQr205ArtQHUgvvV2ZQh3xxgxn3SaOu68G+yJrDott6m0PhepcQVNm113NApKci7zA
VyoCUat2Y1EdI9irLHHjtLOVK6KuqxIAzT13KG7Ynea1el/+NuZ1TMXX2X/Lm0EeCYvYbHexNE7w
PRvi5bszNE0QqoVvIIOj94+bIpOT8c/vJVN7dbxaMQ7iGwSymu5ouSDaYTeFaSr90o6MBf1pG2mS
vOjNho/7PX8RIeqq2V19mRjEPNzOYrQr0vyKHbSWL5ensc7jMUg6zVLmTX650+U/QIlaJ1D0fgr/
if4siQJkcZb51/8mvdmmqY4cMxqhveWnHsJGQI24qCpNO7QDy9lZbpXkrwX/7VgtfC1g5hsDYLNw
jeTHWuzXWGxvsyzYCeqCtSMPCIRUuf3qMO6QTImH1PXmLVt/3iFDPMKMdjSQKT3PtjJkPBSUEdt4
kwAADFcH20d3PkJDgy2L8aGscvvCQY85xZ9n4SSNbgNG9cB5T2SxObBbHWyeenBO5Z/TzeWSKvR9
3mL5XIkyABAg+PEZ+CW7HfdIM4GXE1BUZ41GHY+9mV0JkLjSaSC6tlJ99A3d+VHtxM1D4mBu+/bX
fxXB1gU+oqo041p9FT0EhrKR07RmW8BvlKwMekSuGHIN0h+JDUMqWBzsuOCmWUAEnZ/GgxobH437
MOj2eBEWcP8NdleE/Az0r9fyoFFIRvm8vqEM/3k3JJb7dA3nrGCUtieYEil9oSSXUyybennroyor
EAa0zxJUjInsiqupvcv8A++Y4VYxfO9G+SnQJXrGNhbskRNuNMGWVIVZV0ggziOcvGuaUXwp7Zax
Dt4BT5dkPT2xMDMnwqypoVal26mRXygm7/QXtpac27lTj17b8DzbwGN2gL4entaOW9V2z+S6+U31
oBN5cr2VsOtE7zUY1IjSg0DM1RZKp8DWYmWonEMxj0rcUAmAiTY5bGb7bSnviRIFems7iVLpTNkD
n52JUVncrGWsIjoL6wBlOEl7xgW/qxqIzvaNmDny8RHfR6vwL2w/tLrLmV9ar2AUV/23FxTanFoS
r42sd8OeWQdOvlZ5Opa16FFv4+vLXJfxgXHcoXUx2XyFWRuAspToYhesX//Ze4suQjX+5Ltgy8sH
u+yJhHbNCyrYaCq4em3A7FVd9KHMBPPtjVYwPhcumg80kSuV9fHxtWwEfqfAK6/wHYK6Z4N6k0Rg
SocYRBorDY3hqh2aQ5ucH+gUokEoaUqoMAfE8E6RB72MLmYk02dIpyQjzIyztEZTpBNH70E+ZjMg
xQKQVvCv3YjNm2munNEbouhm0Xd7kUffvk5ITB8XaG+tYHcuMM3YXgHJHhkniWPPRnBdEt6gylXn
fTaf4MKOHvBDL27Ux1NbtdR4MxEbJEEIMG+v/ZQqRiA6x08uIWa/afzO+htfNv/JGw0WawbhMN3S
uoBYZl7HWK/22nyAZlRKajdAU7jPpTS6px1QVkFdtbyhupTKlAY9an/hoNCRzTVfBzAXOBSR6acC
6k+i0gVt9Tc7g95pOvRyqOHqqHjLBlxN2cC6MYjkKvoOJXqIg3Pq95pxrJ5H69MdmMmlp9ukYxmJ
ZwIY66lvo/cM8xX5W8lcXB2sat0NNX8TDxtsvpqfN7F6ri46a2viJwL1Fq/9Fx5xA0bNapv6aSda
kF8RC+z5gw6LgSFT1WqY4pL5HkWUsYBSK4U3P5J5UK01FpO+oFGv3LuhbulbRQqw2otxvIl0wE/H
pL4s0sfY8JFu9sIQcDJ7Zmv9jDm/CAcTD2gdJhKd20cFaDVl+6jn3INf1yA6UVsK5pCz1Dj1y6Ku
JRjA67iH5eimrUul3Iy3+fxN7t2QZbeJgF9bFcJFXFzhueEm3eGtzxVw5ccMpe3NDqnlTpCwkOwd
PLwG5qXR2KyNzBhhnTY/9sxhqZmYlqJo7bqg/UrMFKvw2ClSaQCFfbX07Hb3Xf7GvAuNNatyCxfI
97Wu/7BCi0jtKMtXfVnQoiDjfPL0MIHlIsvR8e7Ft4oPk+NAIiMHW3WR6o4HEQe+whN1Bm/h0asD
YV4MoSRKOSjCdgT1nfeUVF+jO6dGwAPOpZ+wi4nIumEQ8XOhmltqsFvFmyAfeznlcsBn52mGUcNp
feicBZ98zB/qSRWlMbghkXdDp6C2ZM9EAMmzLbnqperFAevZaLneQvXogp9GGGAD3Ji+LJqJB/t2
FMYievWM+tVCOmQVwSrityn3dgSlS8ODkP8E9gxpclqo2fKcC2FctnAweRNUJIxnT6GVjuu81wz+
w2rJRtv549lry8DTI3WTwuM/eFQoXS/0skQg8u0Sylv9cJb6IqvR5dNUi7qWpCxcSEH4htABGq3D
7hbxI8NcxElJItIGpQv1WtrIB+eO1+U9xeaEWD0dOc+ZX5GTzl1kLCEQ3b4xEsCoLRpOLz9BYKlA
v2pCSbgV4FRXgB6Kw0HpAcvqfdUJonHAX+9TkVUgHwCSfiR3XDt12//jinArGskkA4Vf04hDkQpm
Nqb+ptr/YvsgeR6jiIvjJzr0UWF48b5xzdMRwURb3/8TVvTdusWOOIG9GsrGGzfQdn+pM1qLVf+c
nkD6+iomSeY89M7/9TmOXNUqbNbU7ZTlM4fny8xQujthB+z35YC9zQplGPkPybbplZgDJW5nrvCQ
joiJH+xf4IMuVT395L/U5Wf38uHllU0X4JJRaQusS1GIn//O3+Xj93EcVpkBKgxHdyLFCFzsAEe5
rS4zLxf4ZIbbSnDovueJFBOGWtMWE5Q6/dlJUsgLvO7ytxaswiCHGE3RlkBt4kUwc9A/XXaTlG9J
k88yVI7azDkDlHH7ARRa4JR+qFllOXsVVWx5gjIgqvgB5xf2WejswMTPkpvt75DMq+pwuEu80MUU
nZ254Lux2hJ4Akp+2v71iO2/sl8wly9j9NHLo//cs68E1Q19dG8CcSSjlJtBgr9pz5XvgxO8UBlT
2K6L6OIXJDgcOO+rKLcXujGQjPy7+I+Id8sdu840SItoU9Je4WVgmzsAYwj1tUbyc4onB4oPjhhh
NNBEKISrFgJ0BjvdpnqW+cEM9nC4NfuC8X2v7HxfEPqz5Ba4oZfOqCHmdMV2IbTlEytt13a/cB9W
ZJI6EE6qD0LNBEI/LmwSGkLeVpDq7txlGUDChKMloOBygw9vD5u3L3eWquV27/Bsi8MROVkfZZvI
4jX2D590vv3vK72Ot0oYkC0E15QyoDm/zl2LlYZNUgFXyNaOb/LPs+PXASxuwTtLkuIOPtbDGs5D
qApq1WiNYUjDbo3DM0D+tnN7w+BV3yDsLcPsWVudvBlK1OgIYl4tBRFK3DaGITpo6l/pPpTPk0BD
qODJsGdnYmEYCncS1Kon0kcybn3HVIUdwVZzRtCUN36giOEwiuPMa0pv1F+tMUgG1w93F+a45sWl
BRlt1VetDOCmWwWmaCUMlXIDqekDCXv0TW5FNz+/asKg8yHJ4dJzmQoBxDe4eceWrwVhT118t6Xz
wPeu//sI5R5cAhGseKH3Zh6ho2pVckh9iXo7wwf6tJwxsAJxZjs70IuDUj+zyjap3qWEuahX/5tH
KC44QH+hXvUNn9imfvnDE25zpcX9VoKcZRNycD6nRLfnM71yLkXRiYwc+alCSijPybAif0fnnyhf
sTZfCdJ2ZJoQGKOhgfpdCmPUnUNivhXcdjIgG8dW9lJFudaOFOHRvPkXmQOOThk486rYDGGlx3Ru
XLX6nF1nIFVyl1DwePRDLJBU2tLg17nYS7agy0B7Frh8F5XPNPHzFwX2MAk+CJKFIE2lmWPeaAxP
M6h1eMuudpf5U9Y58HOMytD9vOsq873znbYGCCMsUNW9X0f9U6hC6/r3PwvUrGYxJxAn3xBBWx1n
SbD6/syQCCJcMvnFAH4CsVSxKsgzrKVToMUxBQPp7s4ZXVRIJxOnWBo66xhgMiM6zyi+UwSclmKW
ht5dJ1UQ22Blv+GfuMM+qzTJ9zRCg/m1/M7LdrerkJFONc5pFPMndyK46RcvxDYUj3yTkowyzeBh
Rpk2qC5UE1pPW9mKu+QS/JheSEY1L0f3YK4mz6N9Wp+8ieZZ8CemRtV6ls2OFIss+Np0t3JOwn2D
cTUnWV9C4MBxgBTwsFX2gMEb/fRqdi6HivA409yhFrZcXWtXGQW83eODBiq8PBB8P1tW0XXFAQUL
3wQAACdWAWONcs/+F6X4Vm87il9CtVCMjOmUdtARTSU8w1RbGntvaCqegu8wlCu2h9C8CYm5b4NJ
3a5ra8KrRhsscy/3Ie9k6U+Iupjx+LPoy77fpzmCLihDG533xegJTro09uLKqCNCZS++tquq+sHb
5mzkp6/E238clmBVh4Jb7zVHxV1OmcuVZCLSODttU4k7tYqpjG7KbHmCK4xHQj5E80Mwjw+HYTo+
yj485nv2oiJCeZClp5lBAEw6H3s6F/GL0DyJH7O0RkMpblKktOQCoUTq1ZAYjN1IGZ9isPiYiVxL
gcrvlZZfSKpirM8yQd0iMe6Iqp04nXR+WI4HYHGmy00DIZJesUYAxCMRXzFh3dONa8DUCDwOW8eB
Mkmu/icT4XJNN7u/6vE8Qu7adVRn1EqUEG7JlmPGuXjfSbqYRe00hqT6XoK+PUaZfCvOU/GZRxVt
4BkGVvtN4kUxcl62mFaHWpspKkqC7BoUnsDrzFv1kfcWMwoyZC1hBPD/pPFJNETmtTjhOpRv9VP9
rEoqfT9cdw94UpHT94PkYeXwiU0wu2fCrcL4xWkzNgMwGha04KC+8K9vJv2NlTDKdSMbfT7yh0da
1Shmav3NecplyjVOI2UGGL9VLrgR9F0g9fgCcbWMAJ+AmFXEkCNCtMl0OiEOtk5cDpmWtdF3q0JE
e8jCh+i2z5WwmfauUVlbZRQcyobMSVKjUAXS4X//QcDRCc/v2AvHbkXN98AUa2zw8LRZqA4+/1Ws
RhB2hYt1mPn/DiqsT6GQNVP0EykYOf1hQNVvw/TU/+6RRQse+KxUx5HVuo3WSsqOE1Q6uAtQXehz
GvS3y8eH6ab/i9pzoHBpVMEoyzpSe0OzrWjg4xfveoA9CBMCp32e17tM5MToJ4988Dmu1AgAfXUS
3mdAL1wAhuSKYHZ0GwtVsfRtDaWcB5FFi5lN9/bYkq7r4a+v6Hb8znI7eu2gc5rYlOzRYsWW9mZk
1EPlyFApB24TAukmRSHK+KwhIvidNk4h6MUav7bgial8hoFTFLczUimMSVKFcKbhT9miSZgsw17E
pIUNlNfwBfvqaJXEOrNWeZJqH+VIOWIcJ2ZQ0R5GHNDrAwVQe7GUreWtfpCH6hPBKpMblqpOWgyx
JCQEUim9bwGWn/4DAdEz8BbdfxDRBrFiYVE2PQUd73uK7NVBBBzx77X//j7Tw91g02fCDfrNmrks
pgztuY1g6hgOS0azZ2/JrdygcEvqlhK0mUIEx/rZddrhua0x52eg0q2qPyRSGSRafAb3Cyhk06mu
KxOMfSw+6SLDk34mdMBpqO7vWLzt+smnbo8LeQRKtl0VAptwaRboX8Fo37uq9XkACHlcgikUENFo
vfzoe9vGWKIErauywnxFoZCDKm1iUwzFvPzEwd6F9BvFAWX8k30Cbk2WrjAwDTQdgZJRfOye8ZZV
zMStnb1blpfUxKQ5cTIzNmPsfUHeNEJtLrwEYG/k+8V5kGs22Gtml1mpHoOTSuc9cg2ROTFo/3lj
wc5BSakX8DNOYMhP/nKg+/13EGishUu9txpkdq1kSvXxEnIe8MDFymZU+G199w53SG7ideSfCiTk
+V/jveSMm7B7aKcktW+C7Cxmq7RDsXEex7te/YSApicOPEfNtwR9QB82HsFR7DMYHCitKIPUTTBM
+5IAvO95aohE6mmUGEmz7lAP3ZjmtLIY+4Hj/sQ9VMkWcoDeEe5ECsk4vCX8RF3oM7GLM+T1Qruk
hFO1VKdK8+PoBGw73EF76WSfxv7KS/O/tP5J5+F1SQVaRzIjS+n0C5BIKpWVi18XEcBAU98IbQHq
E8or4OBYbbzXpWEQe0E+uExMvpGXemXRe2Mb9gXr3R0uZby6iy+gX0r8OBeKixlYeTmO3X2mTgXG
JkpQxE8k/Qpk8xwGKz4sUkyrmLjOegoPB9vdc8TaZ9e4LDmORLW/Lba3zO8xHL+Kt32IrL+6otsi
sQ9+DZrIfZEV1jfBlsfOIYkBtyP6uFEp6ZNnPimXGxVcDmCMQZ8HAi8rNsR5eU4tb7kKHcA8D0Vf
E1fGFe8PZ1hWGIjBqmp9BaL1nTDf9jrY8fjSidl8+RhC5EOktM4UH9vN5qYHVnUeWe7UtPnL1S6y
OpNpuD3Le8NgJrbxnlhgLuHpQLoA9S3rUHtVZtRHj2tW10pQlFgAPvs3LGB2WcvMqV0ZJol0FsIt
rYQQxpjjEmKDCJ5T3dzhbmiaJyu9IRrfsg/ISIPwZLR75Yz++M/clDn7wMB0c/tPYb9LdCvW7Uuu
++HI8dhrtagcPNOHZTDPXWADmHMqDCF9a0HmICpIUtugnk7SFupMGb8HPORtHOY3PhYvizwd5umr
KLc5hWDIgSmT27GvO/aWGZAwbbzv9u5NBGUFH4rFjrkCwA/jbWoSaxXYVeX1g4Co6/DQdb7Acmxn
U7hY9DEbbJyeZECzbxwsYJFvxA3tkAgAaJy9ncNyxsLGn1BgJfiZe4DnSsTnk8RrPC0UzdhbufG3
Zp+PIETc2WsbWNZqv1lG1sWZWlLGFOsIHhveJbWx1E/gvCa9yTDXvG2U5ytCmieG5BQHKzEEgfeD
V17gZsT1M5lCbUbwRPOh8P4M65ymOUGF7/LQHRNtloj7B/IynejHmDfHYhDrSyI7sD9bRkI/2Hb9
3lW3tD9LI6pEqoYq3Cld+6LxKOkfSsMrtIR8P+6DHShtftaGvbM6nv0mkjzPsj7PH4Z2VKxyJQGB
prGBLLgGPncJ2c1R0icRU11FYFqcX6ZhBxBqSHDt0HNBGeogsPEFhxGr01MdvL5ISLE/y9GJk6nm
lkA0xYGjETuHx8kwpQW6CVDqx58bTrGONBZS7IgCN7egtIXmQtjNnX9ZZgKFujULHjqp9kf+VYOa
F93nFfDRLNMSL8ARZ8VnwFt1CvfNb4iqRwSUw/ssiS21Mgxa4v11XIow0JWDbgJ6kgW3zSl4XXJV
rTkWTKoU1z7juFOHX4tQ2kAIwfF+EUxaWstk12+kBlPXmhxEwnmgcf7MNdRH9tJIu5WVQv0dxAtk
DMU2R9z5a/2TxxvuPJ4x1KdejzC3H1TuuViJ9OHW0EuZakTioGgfYBQhrcVFVot0R6GrymEubnob
P0m1Pzpsbl6weYstF6vWuQist10nurtBIAJwQhlMNWW4LxCVgqBadKqex9dsZukHjtfb+7vAnAu5
UmI4KlcK5+Q5+xzfImDy86ru0NAUWZ4ZKXzlHWUNNrWk7xr5+Wfo42PywjDhf63GcfDteHgHdFAg
S5OQZoiiffsA2NHqTamYTAtYDvjwOWNfKHLD6NKTHZZmk4f9MWWwESBefTngg2X/agmnPg8gIDz+
tS70mOMa9dqz8ZulV4WhiV0W3sG8DAPZxiTulS2SnZx4uoUw3+BrETxxjWMtAiy4CsGQxe1oIpx/
4oFMrPV5qqgd2/qQgVPeqekSdQp1R6LwDezElvFwClyESBNKxd9pM3Mw1LiYKpGrqK7a+7Mc+cSv
0Mmavam4twnUqvxk9SEV0VT9dxbZzONhHQ1brsLoF6GTRKl6T1/LO7xxLPHkogKVuKJ/vap97m5b
90B6FDaaPfXAe2Vvou2VbpS5WYyuyKOcdpkj/R45pXBn0zcCf9x442UXEcblAoTGXvAVtWQd9Y3s
m98udlm74+pu35kKRtVnns3Y6iUB3ThSADU89xc0UkQhsjjZBXvFAR0be0JRyGSq1y0hOipyKhFk
xf7Jx7QkmKiGZeSMLFZtPfzSU4kVH/oaRcTk9YJ0ie2xzP8NpPwsyuHXAORsL+ywXL06XeWRBzE8
5lpJxWh792f5YkixV4n3nfMQZMWj5cyJx6ZbuOhu8d/WLh4VYxuWjoHk7GbdKn1HvI2c2qOCPI8n
E6vBsEpgwAyarlB40U7oFoSkpbCq22IGLYkpa3rEl2yzH+zwA92yfTLHXUudni2ZCErxjdGi3dXQ
eTIZYqz4mtYZBg8fiv8fZFeB79nEACIoe2wRGfLvodMVZ9TWATF95vUbyZGNNVGf1lDfveNDlgHX
vz2ZEppgDJR7it+7dUE/KRxPC5p9fSebpZ4bKr2JJY+yCxO9b9J0qlH0sqH49akXslwFJkxsrFaY
jYGDJkDBd29LdLxeOpdPZTpAPlFVGRX8pUzHgbdYJmtCLn57Xd+EInzW8P9fiybvTxgQ/nJARqj6
+7eHXissT5otw5wYBENukW2HM8xpfLsTVH0kFQZa+mFF7dyxKk5Nim8jvxmmJjnXahNIM04B80FC
EQSrALPSiqgces/8A7x3fSIA/Gd1dCjwp/wzHLsOwIKXt8Gqofx2DcXZPbVluLuklTx2GPXJYSP6
eDuCT8J2Gtu9sGJg+qxc4WurZnu+/f7YQselMnS13o8xXe/8DqMSgelPxg8YN0BBll4omH7l9xok
f55854r9GxDV8O0hzmTP1NgZK3v+gfHGdJlDC20WtUcnabmIkgndOJ24fehQW3u0mimk+7rS5qlD
cJMUr2dknO/PrYiGAgE9exWFlKMmLK8K37riCax9UtFxQVR0uJukCkY16STjAMCsougbPwQoUvqX
W/G7snxh2A98I7Wc923kctiJybgga641XqV0cUF55FYLmcsb480vi/DlticmS4BhtZLzmcId5sSz
lpurN3dNW+K8h6pMyj93knjasp1YSx4X07Mq6wgtcseOkYZIjpWV4z5D5Ldi0K/rPrxfzaYCbUUb
vVaD/CBsUvSA3velcasMe19DeyeMYQhpoWeNdzmKDlFakpeCvsINSNXMQKcJRwBTSpADCDh/LrA2
+OL1FQAEmVlcAwbOwSF/8m7zmFaUwg60nU89cKE5FvwI6yQ0E3OhRJk/Fzk7NSzjqP5u2YWk6oNf
hTPGrBXdVhxXu/BSJRaZQBMQwBHjUKtC3pIFAHURyjJz0AgZdRGWtApGhtHHSYvTYogCWVAwgbez
9DxCQ6ifK5emrG9fD77G2C4BcfKATO8EP7Eel/Zk/h1viVbX3jCbfLKS4335FTuoYiGdDOsx41cG
thGKNd2wpgHOB6EQ25meDRgGn5kI5bkteHJHlvGYcA5blNvrB+73iTzriOQdtZAtSuEHVgComggx
Wg2apch+kE899YzoK34QQiF+r74kuc6NHfNnMnBnhQyk/LkRJ3SFz7YdzCg+EoHCw3EqUH4WFuc/
7B6Ob7AvU3XfiLTJhy4hrKcmDiTcZsWiVSITSKy2m7BKSO1ziqQEfYb2kDt0c+8HPjs86fNWRlgj
rUSfM6wQjf47g+kh+b3r5aCaCvEQIG3S1GIBtESBfaeu5K3aTyltZIhC5HA4B1y5IC86lEksH3n1
tAWd2qDtI6mLGngirjPXitu2TaPfAHwwRrdeSCe54fo32mnp/OjsDuwgs10EoBtYCSnjqeBczwUb
LwEMP+ZPhnEPIBD4lOL7Gux4peSo3axu8ufeQUf/htL0rh7mSSHihCTLEbxvUbaa3uTH92KxWf5W
9nXAQMXWXitVAVOdxCgs8gnd9C4LqN/N974dliwOaFdhp/H+fKMTuIhn8oobaIE7YVLccRbTz6rf
skfZi9nBlc44yf74YzA9tlJfdQWt55ictu69hSJGyhcY/4K6Sgi2qZ0sTvQBBiNXjpZV+fzci2EM
HZBhVvHqCE4mH2N3GKKlmiY65hsP2cocj6PcSnIq+KpTiuXY+zD01mv9ZJObOOtbJnKv2AD/sVgG
JozAF5gX3aYkCiJMMU4O54izZW2K9QRHqlm2Jt1k0U9M73JE9sR3RE/jemyfmAE65LXar1LTmHhg
izbCrfyLeKzPAkOZWh+qtZOh069fSo9m2ys9P7EQk3tgXyPHVbJZ4Pmvf2EUxA4VDviibqEgckB6
hnTcBQ6iCxyrJs6M/SzUAEcVhwodWeo882+BDeTK+0Q19XqvrPnI5MyL3ORcVuCmu62txZq+IcnD
xkXoqpZE3WSKDAUNth1aavSPlYxWTvWuTM+rELKRsf83QxZotiMqnt0hGJWDFcBOJVOFp053MSEO
KKiUJ1uTFuYjTx6adM+0UOHF5YDZx4a1cK+QekiKWMkT2PTAgI70Eg6VkulwLMeICZC/rDfQSw6z
nbFg88bUwoy5qhuuFvRwq98Ppso6Ntci9J4OFjp8Alvp2j3ZFMswZ4lbi9oH1fk4p9gsrjkYkL3u
BNNb+BNP2efgsD3yk+Kl0lPttvkh/ZmbrWEpwCWukMV9tafqaaGgvUnG/hPI77u03jXfGJG17DRE
oe+SGr507ISp69MVJMMt6e2BN5Lj/1qrrySV3TaXlDzztgS/OCN4ETBdEJvSFhw9W4qT3YDSi2A6
cVpHRhwN0Cm770c2TjorB6GF9vio+5i7rcyVi0mHLPVZWIHJW+gDQR5BDIGmdmPWeP7Yx/sDzq1M
Q82UxH2eZKsyC88Oj2MmOMGAWdNFku89vmX3JYkBaGG14MZ/FbSBqDY0S2VIFXtwkI4InAI+5zpc
pa27aKy/AksDCH/8ibZ9dPovwzR20sxbx533jkrfaTIYhNh6HPbVaQNrtLjR79JyHW35Z6c53Jfy
0px2Zig0A8r/UDugbrpB+p3k36RFUseQNSZFGDkvwmUTPR+7HtX2hgHFCyh1Cw1DA84Qq4WOsJaH
5MiPqkgwL6f4LByFufYFXcJ6FnDc22Do12WYBrJMfAuRnGYZXFaO8rVKyDt459/soFZAq5bCfm6b
9Y3dhgdLDMKBePF+xE5SAt/YZQrCEP7snyZW/HWYhwVJPhOxux5R84+I7ZZN+Kwrbfe4mytIy5xg
98tgCCE6aPJUz1bA9JhyGSltrx6bzSnU3QIRt4tR9lMCJjs1s11jPRKTKonsMAnvYjFDR3uk+F3W
0WRWcHjMnJe4Dc5QwbiJ7gg8EO0WqhNJFFhnmlaO/g4ux4zuKej6ZVJMYaC1DMaRY3CagkF+LGnl
w3JM961Z7MVt2tIBShyhuDHYm+WonW+LWv/qe4a5F+yWR41uD/LHF0NT0gAhwkH4N2lEJ5Z6TVp3
mKmacJJKDZHtGxRo7OTvt6a1Xdk2sLmjjpdZ9VHthxUG5Ju+okYRDmecfnIUOdtM0mUouWcLSGkh
BSkn5U0y9xbWz2dSYsdRCm5x+TVZKT+3hrtlCegrAn1EZMH5aZt6+gYzO4sBwOqShdRyKPUjquwO
CQzi5//2LDI76IWxtGgCdxigx1DSRxBJSg2MXjdCiscvJi0Sk4XWgeV4rd2OzO7xW/qebeH2LGXc
9UeLl2uVU/yLFyUbETCFN7mstbiUSUqByDzPWpJw+m3K7kdY6ySl0Qmt6dFvb6zSZjbeG+NFExGK
1qJ92jQCODPzX898qgKca5s1mOrfe3q+ditC9cZexM7o7lVqXStG+tHpIbAZviuAfmhejmWfJWH6
PTKoyGPHPrJF4cqwaVuZ+Dr7qVznO/126wSH3dcg9lv9hU2gFzHK+AxXMWN8B3WndQNbSrxO1QqR
Lm1Ze2Tc5YHi4LmIo2L2jjOGIjzgp3GMCmUJ8p31ot45I9eWVZrz24vfBnwNzQ96UuwtmfjDJTYF
jKsu3OZldamplfHcnRX1aENv7NTp6AqNsWNhokp+FWDVPCPdkv8v8cwmxukKEarnuwnobm8/lf4f
sQiHBYTIzzlf5L2wOxxNw7gjdAdERIpvYqFrwAVM2eyMda4Uqps2PeZ+29PjjeJpOrkLg0cwElKd
QvGCDVr9wFmCtLDWzVdGXR6E9AT2gAXun8ZQc0hkdyFQ47Q7sQH1vgpRAm/2CLC5mxmPJnDVwJls
dmlSd0Qqd7znUxRXtgzE9mVAZ9YYB7hFtzITSv7iCfPJ6NHXa0jvrv2zfCElLvp5BmG9NTejd6sJ
mmpN1tfIKpECjgt9t2QiPb/vm39nFNJOANZbAwFjgRx8L4GNx8yI8Ol8gRkqH2M1Gi1awcySQbdS
5lQigiCe617ka05JXEYf0kGEb9uOgSKApIt7H1ch48skmM3PytDGl16Bhd5IdZiefCTptSAhmQFw
su4s8HBsUOcdxgwQewj6wCBa/CzYYq+ZxRaffGZG+GruO6QeI10z1CTkTyrJaPSZzZpUqgZbaT7J
5Fc56oaYi7wZCHUt+Q5FvakmbYCqMY70sQtxriMD5gn09NM05dQo0Vc+NTIO/JYZSfJCns3YU0Bl
puOhR0tkc8VSzw2A5Bs0ZeBD0oFGhqaGFvTkB/rrSuLhkSiTT0z3AXyTtXk0ycjvqm5hhHe2QRo/
+LrzaMhS1m/wDVhuGhaF104v7iiCqu9Wkj3nejDz47g1F7fP/E09LhMl326pyvCufEAbE+o2PGt6
dNGyju1vtR0ertH90rIQr7qRJI/iOd7CLX+C3tIBtCU/AMEbKW7IDoeDxF4B5uGNWIXnn8UL0m3r
Pu56rIYrS77B5UXLGMokzTSRDfkJWnSKR3rXsXTAohzLu8ffpghMUTNKQGgBUlSqUWy/ZsmDKK+f
fzho5lwzo77rECzB14SFt0d1TqkF1T8ZXrHAK1lNMABpmh6MvljWxnst5ZpnrwkOk+GWPJVUjeQs
rRCfbqvvvp5dceeE+sZ2yiCaWOlMSxVwzApo/USMikgSmzoTX/ENfQ5N480QzQ48U8Fu1B0Q/qXA
W+s7B2w3MixwIsA2ADvmjSsSoaQRMbgk/a4PIxE4BsOKHOiC6leT++KXpGF1N2P6lslyGlRYgqB1
L9xSGqaeNsSAjv+Gf4yXIpHfptKbW5WjaLBVV8dr26niypVMGopFCRKTUB552u48KaVUFhqhqW5+
fYNfEicWY+W31QqiB7A+TYJ3dJgH4BVgR+IzsR2fBLdbl5G5kHnsgARqFMQjtHjrLr1fKfqp2hTC
X124Xg9QAyJ0NMT5Xc1XKhV1oAFmQOV1eL42ImVl5T6idJDrzXA1MESJB2D0ywkwh0lXp7jbDZFt
rAdDBibRNS0hy7OuXaXtbfdjB883HQxmbA41Z1SmXBGsWikKgv3l0izBQf4MLlhJW1TLd+zcuO7J
wf+cxzn6xAWcLRl7eAETzaiN1JP66kmBSdmvw4Bk5NAVNF7zG80hAWsi5xvCoRHYe/tIv9Q9yaw2
z6+VylNE4CfFj7dgRcfUhfXTr5vzoLHa/TkAMc6P0h9X9qvUO/hFJ6xO8WmDRjGi2ZTjIwbxe40J
x/RNbDSI4Y0ta+WlijJkpzcfNpf1HRKO7XreBAsrAQN4Kef2zi7UBW7+BUR7fdtd+x4JiNPETHIF
IobgctcjMMJAW6sHM2UwAR+KhhS13MFKN4fKXU4XK/b2jXQmpopWI5zV3mzmGaryPX4z1fyWspIU
jcxOtOGQzlCMTcaCBrJ4aBXqIB/NueUnqvy4+IgY5mkMNCp48Qh5R4bXOuk52dUMvOLp3V/w9rpF
jcHdhnJms6C8/U3w4w8OoxDWWdwQxVZh8+jJmKtkYMd6Cpqa46LG2oU3Y6TSqzUk6KHayoHkHeJc
n3XQJb9HBhATWrNpkgutYS+tQA+Q11k9dSqjKiAjhsdQ+5O+43sxvoPJcUPBhBPz95zF+Cz7znyx
wxUbmBI/PWcskXTifq74FHEPTUByEqn5r6TInO4m09zlBJpCCtMOf5kSIcRW6zqyr9Y0mfUPcNtc
/0EXW+oigMY/JIB1FrDNyArYlTwf0aRbe1lXehk4OIrJOgmr+jjv/WFzlHtJJAw2zWLaNG1Gwbed
qmMDmQ7C0DYAkbCkDQFtBR2TvMj/qhmSv6TmbLRS1dUUPZvUi8UR8Ty72yiY35jlrUKom+rt81e1
R5sK6iz7mCs4jz33kAVhb9ILsrxTr01T+EFQ99SvQgna+6wEb9aUF9q4MZEpqHVdBVPTW3Vb3NeT
eHmWfnANfBFfhJGmtEI+a7Tk1OOQjxknAd+b8vlR2ptSiutkSTGU8Dih759h+8lYo+D/XokTB6jw
nQUWwUbqObTHjXzXr9lhINPSVBqW0EEBzhaq8DU3KZFUJ+cwtfoeZ7Q1o4U+9U2jrS1gMY11bfyY
nZdnsIL/bAeyAUz4PJ0VLkcPZbPcWDkzhC4wDkexziW1HUZ9LeRMjVTTEGIFm4IiwCQAKw1G8afE
hZE+YSSIf6O7DcwUtQbA0pmVytRaFSK9zkan/B6BdH8qSCFir48NeWNCdMH1vXKYo6noCqLaGaow
R1r8V2SLDXd0K+S2fgmLpNVkmCSths52AwdX9KAr/Mxf/zRuD2qeyuGDQub8dfdVdbOUk52vY+y3
I+c9C/vBJ6Dyfs+fR/7JlJ94M1aX2fU81xHG4mzBf8n8GNY7+l6wn1HKQgR8bzMm7eB2Epo5fNGH
5aRNJridjf+G+qnnvvjgfiQndS4pn+aSKabdkfy0/T4K38pYHW3TnojPKFvOajzuD1P9Fl9hWQNQ
k02Nyu+3rok1XhUePWfXK23J35n8+fZdQxzyuUGZWYQHdMKEFBr0sTJAEbZmaHJHB/ZGAx6yJNN0
KD7Wdncy4cK8cbbqOz7Z1FGoyO7M4xiH+YCdoaceuHUPyX8KGlXueyR2GO5ZMe6RfVzvhCCu+LKG
FodH04WBps1y5W+j3dLp8OEx6cjo4hr/aSW+SPwRk1aI/Pm7IFwXp5vbOig6ryVa87PNpWZ/rJrZ
N386fM/K50QNhTKhc0yEZlrUfdRMEwdRn7cVFu3hFH6BcokqflaPG+Y6bSGgczxGyQYw5NF1NLAj
2n8McxsEJKGaN3kr4zSD7tHeSXQjBoxem6o0ixNQOKyfJrCA5Dc/lkbAT8JsZycwmVKruQ4v8X7c
0GYrmX5C5c1loXLqzZjXBtHnWqb93pHDWzN3HHaweJivN3X3p2WMWv//Xw2nkdliSVhRsNntFbP9
J8jFJVvoPgHBiPn163FrDDsrV4oxbKWZCwfbGXtBRhxL+ktdqtlO30R9Y3Onpws/P0Nvl5LGdkXJ
d4N/x9fHcaO8RZcyECxle43SR9qdlWJ8lWrIN+2GHQgbiwsaBHc30XJkLVZyqNfcy5YN4OZzBpqf
obUlJ2CErr0ZdPecH9hmSZeYbTq0wEeSD+8vUa0WA/q5gF4JsSdBT6VAW5SYkUTDl6d3MB1LSk3S
o2850Ih/toisj2irP3WybYerdAwg1YvQAKXUBkyHTvWlDA02ng9/iPJM6fULxVlmQgRFi9U95oh2
V/9MyZR6iwsWb38mmzlIiAEKllrpCllqbWvgrdwK99Q8+TI+Y7Y3z95vpRPqUFWzvACFrsZ3ioMI
4PZX5FvWPY20wgK3VLG68mFQkiyVDxO2Wm17QFgO6Tg93tL/u/BOjMVVby3qgzOpw4NzqpUnyfku
nUaYzarPsCgnS7uBVEcI3/bbU8QYjz3miM4ktY0lr1bbLI4wqoVdSkyeO8GJkgBe7j2zbglEdKYC
602TFfHRRczLq2TiVM3TvO2Qj2gXKcS4tDlm8DtFr+KtuzhjYDCzgItHIKhojgHkEPX/QaVMx+xQ
gJ50ZKog+kXVHhz6TLmO8AtD4WNfq0iHGRryJ420T+W/670ss66CcfHx+DcmNMkId4S/7akVWgSR
JdoSR6EPVRkg8Ujro8bXOr9mymA68Bm3WTgvIe/0EyNgTp0NiHlJu2Py6zD0MGOCLBFWS7l45+Rq
BrQr413SPhSPwkJQc1DB2frYSqMy8Z6tlaQiHV2dvAEnGH1Yx7zrVqZ7yJ27O0+RQN16ORR39Q3x
MOjgSvQ009Huq4lJ1UYRuhDnw92nD0OA635qHllllzYPOVAkEoATtwDX/kbP8IbUY5oRtvnsDmPX
SMLnelpD6a3It3Hx3wrocUWZVm95KAwfbzovsnxzmyhsuZ6/UEbQlTnuEapkrOiPAt2t4H0i8sip
FbwxxbqpuLHrxrIB2U3k2+8ROgjg72asH9L2GBOASalLHs6Ns+at9K4aDluR7M+Pn8rE03AJ3anx
+BSj7HjjupcXA6jvg0u59qnYiru+wztviDY4SohE1HS7Gm3+ptyeLZRxroC+b4UQsB+lGI5ZPnTy
xsMNVeeI4pZhGOnCC5hfSzKwzZyQRotJDMRlTqJycatuJCXZJkNhLMmdCGuwWGX85mtaUkKB2v8D
p3BV423xFCS68Y/6628b6YWx8SXh2fUhwvTIywqqE2Dl+qlHPudiJQq8qfSEB6UmRXvJUFZe4sbr
NR5+SyQYmhAYgLpTvllez/vzmOmDjiR4XKaAWKmVTLkilKpvgyUTqRZ+W2D9kFtuUOfwX+o5QU1o
oINlPiN2CSCU7qcVrVgQRAOL+BTlUUkab2U6+TR/Seq8rG9/4Sumuu3sYbPTd4KsDfQ8VP53HFQt
H8Ztxw6i+tCJqUu2fabB4D7PMvUjGt8kUwkBmuNITZe/iap6Xbof9mcIL+1pC4+kGZ/nRosfVcab
tVGdq+DvnN0f7i4xkMJU2mTZWYIBPuHzgFj1ooPrGy3xUG/bRQWe3aYZbmqINUHvawKdjZb89RlY
boRS6iuSdNJHDKCISrxQLnTQ81luWJyGGB6TUhh8zrlNAL4FIhvuV4RCdh0UyEt87YJDB567Sk4J
7aAhJI+taads270CX4Da4LB+jFTolObfkZ2WLA8GHW+AVdhQXsaefugDA3/MKQbtd9jF71qKcqC6
tYL5njonbcwH1VmJpMQjIeO7hLCvEG61hS5TO0+95AOMA++w+gD7BzOTBcP8t1Tu1qwZXSjs+oo5
/yAZr+J0ZS5zMtDxZtvvRq4iR3ZF80zhCTMIO0lMVdoC4eWGXi+eWlaR/wjuQpQCy8sk5Qv3yziN
dQ3tVRQutbpyccTPOyAqkR/qr6PXrTWAm5k5wmNLlcNpflsnquwwsaV2NQUwohC1xPKqycCHIYQZ
RjnsoDTWQkatiso1padwW/B0fIr2h+0h/wPrn3giRFQKuc/SUVdvqvosOYj8KaU7uG3N/dQ0pfJR
exXLmAkdt/ZSiquL3GZaGuk+bOx2Y7cftNCLJ/qEqCwpwZpLuMXu8DfPqYbmTjRfM5/kKL09i93F
lidns0v+ufLkqq5ZqgRdyRLtyVT2kLOS4nvcdzMhi/cFzA7AxLraTAbypZPUeoSgyWczMJcTKoVh
WkT9QRDmrYL7R99grS834KuZM5UHLMQWd1NjPBfOnjHddIN/cHPTKECzxeomKsA6jw5xBueJOY5v
dQu6zhRrWZUrQ6PZ/u9Mh5kfY2GV2CNRJzlbq5oNGFGKtD34tkO5KGNAlPHAM/jyEJs0tElWXFRI
Wl5W6n2Fy2PPZBiMYXeq4gAY+jU/2uYguKtlxsJ52P08W+qQ1sq2wHzDObL5NKRCO02c68QfKZpi
Qg14nsEX4PjrNg+wLHw9CEKwhJrvWBtJH66AWiOwOy7G+Wx1qtKL2BMqx9sa47ZEcmmDjBWvSa+Z
dEm1uZ+SAcfSn2tYzTHyk8UOpUra4Bwf+c/PGQi/5HRB8UzA4cOKdwIiLgc+qnv2Vs4AzX+dak7a
rtCmuSy70DCnKaEilNiK3gqXSrJlCYZmbRRYlAlS7lnH9OLaqNWOKc1yUNAEyWkTnW3mM2hwHrKK
9sg+wwj6Juj3asJTKbeOl9v6nJB0ZcweHwASlNU1SR4LCkG+oqwY5gi0re4yea0zJrFCZL7JqYco
63ZdVpvW0Tivi9QhQnFEShMe8qSoUC2F8g6X1tU8jcmjFHCMFqULEYetLAERiE6Bg2iGK5Bo2G7u
sCaKVgw4FOHjXIEfUypH2gBP7Jr6dk6gdMbrn/wTxvK64QEBWPd8h9RVQiubR7RFIc7JDm3bUCAU
iP/PqulIUFF/G99FaV37Gx9MARR9Lk59HgEnLNkXENIkFKyYIiDGtI72QwCIElijKCVbL2EJOowB
SeOxeKlRJHNSeD6sjOez/f2xpnesW3+Y9h2sWBr7Qe7YuEaut6Qf2r8jj7EWTrnhgmJ+/39NBPFh
/c0JTaUDfRk+TtcrVnA0Zu5RVlfrs8yGiV1LoYf54ihQxZSyvrGBcIq0u0ZgBy2CjM8EO0xrOpgA
IcpM5fDqfwuagBtfEuqpSzw8CPvdR9LlyDIcXL6ok4Zue5G524wNmdrA/HaFmfbyrKbCDdAu0qhY
HNRSK0A0cxbt/DNNpPLWjbxOR/Ka4uQT6gU1HZbmzKWmIwiceQKjth8+gx0t94vefzzbILz9CaG6
HW2QxC110iAWhN5MBQTlSKAXgexGYqHp0q+81cyCFwsnU/OHSCsMfPJQeuyB7z4U4AC+GS/VfvMf
3BEFkP9dEphoujrnnBzZELBgwXam6Nvp7rFTnK8AUPinet63uxqLQQIfA71EaH9kiVrV+pssudru
zXBE6QUo9me4R9UIM92LotEOYLZ/6pFCo6FFIFY9ktzUaaD4TRvsYSVB+epwswQ3NoumkZkseCQq
u1/48QaJQVlOGwX7xYX3huDJuop58mGjxmUe+PzEPnzsr5/ibfCkjkSEJpXVGTayWtOi7K/st1+5
yxznAd2+/KNJSDgkrH51vBKZK6wuqw9lxaFuBXNHnBtHUl7tZwmoc5wtx0AxtDKT8IfrekZv6Ko8
sUlup09s9VGdYAZ+Tlig0422WLob7AGkhBAMKcOBvFDk/nf3BS0asoSakIVKtljFbU929qaFsXFE
TutbcC/iFPVoEZxmeWhwAkT5mYZl21kr+/vbOseVL9xunjujI/g1JarOTpbt7JqPOn/Vy6eDTu6A
uUpNCnreEsWXKp6K5WLUj0hC43buweIZIcXDFZJoEgZ9kqDaCKgRwoxHqS856d4q1hdUdzhhIrUu
AWBKcBrDVj/B9xxK0sYAKU+UHP3MqBy5UCjDL0qLL8YOMXVLM1t738YUtrja4kinAsXT+UtwO/HX
Lp+x+80JLakdn8rbtYl3Mt2RaCMgWEL4I266oHCheAA90ScynbLK1K2/VFRNF0MVfZJ5nAWZ3K60
Xtd4389Y48TgLRb1e46haQGK0x46C957gQC7b7J8AHoM51gEyiQSoXCDe9tXn07IHYHF8tRhRC9E
fS9ctvZwZyf4QCml90Dv4tMy5VxoZEYThE9Kc2X4rr5ndlsca042x1KAbjwQbgAcNmPRRGUV5Z2T
BfiJiskQzc4+H1avaeTGoS/VuTDMTO/TKog4Jr20rTKNb9c+LSCxV5uCKZzauuhq49+NwwOCflop
yx9JOvgPAlsxm8bNTTnJQOUMp4RxnVHMRuVVMxyrcjYV8d842MQ+0yacdCQoJ5q/hn0hlG+3jIBR
Xc+6lAe9MVBeHIndDhuAJTMMy9OH2B/pCSrm1/XQkpHGA2apQCbCMfHGKCdx6K1HnfO9agx8fuk3
wwAGK/qY2VQ49anuXVtYoHsLAIpI8N5MrXbKPgE98hvlkuftYGN1CtNiDbPlOWX5QQo/WLivEQv6
vGboXhrUVGqVlQt4IkrFRyB/wtw3Zk4ZiNgsIcKUqTE/6vgpE+9QH9SK+iWI1Z/uhVyE3aXY0WH5
FyXJ0KGRFRTEfXf5IZIgWDnSMQytHF/nYB49cmObB+z/46l79bawUu/YJGlCfhIS8aseFuqyrxt6
5hwg9Cm+AiA6oN9d4tRl5n1N5CuuL49NETsBwp9ZJqGEKaWdNoYGHlJQY4xtWrMx8VCRWsyCCABh
m7QZyOCD/NerbKMy5QMd9mHHRjQ2+xpPvBjY8YVhgHzD802vrxogSLYBji7pE55bvVa2Mmi392Zv
LSbRfYcbSec6J5e0lfmZQhCjhCF7Vv2RlK4eOHE/u/FdKfmrd93KPVWPfu9jK318i+R/h8nBEGod
UpHWjPYQmQBVOUQrSlGh++ZjrpEw3X8/voElL9V7nmidrU+dLxKt1ZkmTrY63lkSCAfjTkl7xcbE
FAF2OK/Ng83lDNDUusT6XQbsl+F4GYk7wooG1WYMoq9oSq5D8czhzSBWu7dFoLbPI8Whprqg8PJv
XSO+2wkDFLT5hJRdfM6u63LN4J3U57fjIWU/Xvf9w71RaqXnXipYVJYKK7DDDDqhwyjI5DmXkv+6
5IrEnBqW3WK861VLmlAL/Gl+genFErpmhUtEvQKoLz/82VSfm3oIkPab9QNX3L4LQ0z0ukinpy2X
ff9Y32vCHtF0ddceGbSoZih8X5ppZmYeRmJkHRXWkx9vC4lTVI+mie3qZ8UtcllfXfOXHVyhK6vp
78V6CdPaIsLCyN0x3bDI6RnJ/LAef5LNQpmPGb3zCFMBSci2gHMpWJNCLB5HrBacWcGxsiyibPfW
Vk0dwogCjh+OglLnG8TbLNshTzB/L1mL6fizYD4vFQaevPCHt9Ad5t2faDL00m/oYIjvBhihHH1j
vqmBLectIBPE+SbYl2/TuzoWYrjw6zqUjuc26fG1DTUOxZIxx+kxNgSJMdjcOi0xSV/ZvR9U3Ad6
clbM2/Kk9wR0FR1Nc0N9Zm9xZdDDqKoLaAA6jfdFagfIuVyP0YH+klpF5/KeTarDOgVtaLFK6bqb
eKUAN+2Ewq9mqEJ4orC/1o/yFkFkvSePplp1fctEw3tOShXsTwwFTdEqZNb3OwXSgQI/SpGpPav8
EGR081yGOtEMWqpkblRojDHXjWOlnrH4DxaeH61cP9Ce01PTrbImbOlMJXtSl6XdeJfv0OpjiJ27
rhvsVqYTKHt/393dhz/3Cjd9fd/VMSAe44tfS10dmt03/+VV3Ftoj5p1gZ1Lk0lqXP9qEq4UjCQX
rF4o3ZDikozOeD2ifq9uXK1GqSsAna0Cu+4YpSpD4MXNV0HwiqrMKw/hyk+1gd0MmYdFftXDV/z1
2bXcJ0HTHVQpMiUERbyjtvLAtLzlL1NcBsseLIS6hAjUEFjI91qAE8X669phCNVRtzhoZAVCfZ/T
xa0XU13YI55lwv2qy1WRz26+zHIUGbuGiC0K+GTrEmwdc83tHiuP7X2NRbCP5/gDdGrlhoWWaZmI
xC6Ogxs435Y75cYNMax8C0yvpt6BQDlvictkqTXGhsXV6eYFKEvpPKnG60lf7tTJwvTiGIbEBCmO
3KfwspKAFEVuzavvYjE1uLbLQ9r3Uqm+jp9d+BU+uvoiSp+eWMbFtNGT9a9QAu122shytgzZof/M
M2Z0FEvXxknTLryAvuA21HM3kKUXG7EZ9jihuobxY/mCY5IZTdOXXNRKsZWjcNGiPkB8iGaq0H03
pmZD1oID1/06wIfagvSuXi8vXlA8fNOrR1idsylnXk30/F5fOF1xMzDABUyE7b06k8BX4ZrcmPJn
wujmFSxFH7l6oRSMXEOGCf3FiHuudXHPKp4Y5qRcC5/1JIUtoFxaBKU60ElU2QeHqqxrpN21Zke4
GLhYeAsorNS1cgv9XMCZOf487EuLwfQ19Kco/oZjGzaw9kyBqcjVKmXYsYMwaX+GDhRB308xA2IW
sHTLnNSRVGjiVZ9NF7UypcjCyQPtTlQMhvchbA6y51128OVE0STBe8B+jlMJPD0Zq3EngL8UxcpJ
2/V41ByGO7kLuLBwuwo9QbgcLR2ST8MEGTKlqVgHrafU6Xbe8UUr781vM+Z2QL/gdnhVEATvAyWb
tvhK+T9MFTthVQambiFDXfT4xU5rPSRdk0QXnRDpojZlmQImQSYtQ997O3LcqMJWhK5MtQ9hHU66
nNARcQqMP4wUH2mSrRHFP8jE3b6DGocDwj/Fp/5t7ecLT/voi0StZ5kna76sehTU6EyBklv62qrc
kCJvh57gWPNx/xoXkWZ0qk9ySfOgqK4tv3Gu0fLLOLqQKOt21mJ3j4nz5eaqlhASFM4/aaQxtAb6
od2pqcdq+QKbzzB6qV7vsuNsr5NS7zHdIkGBQpIdehO0mXG0HUS8rcK0Viw+mzmeRW55t0NLX27c
XXHrhXhmJTu+BVt4z23WXjO0aV00FwVFud6XgI0LaGuWmiYr6iVitEJkU/EveIOtGdnrK9ndIoxI
ZwufUz2oZV890DyqvltXNq5p+ooxtUXNwScqXKVAp5BMgLWQWTgBoag4iJCDpJLx+m1CZufhn8tr
KFegERPGnIZwpd6TKdWiDGr342hRt+wnoUi6qAGaBvdZcvDo1SYJvF4WYt5nNNHAsCm3v8Gt3ljn
RPmVXta/i0fRxOI5uXkJPHge4DLlEUpQX/ANWIvii6PqoWXVjvmWt00kV3SAtS8Ct3bYRnrFqCKB
ECnvvB9TzXGsv56iQpoP0XK9I9V40yIpryJR//n0V6+FTrm0XcV1GJNoXbWypDbgnMoI47mha64c
QCyd1iyNfq/ciBEyeVTc+Wk/85Ge8Lw46xbk1tD+5A2mXg4rZG/8vNaWeJH6qIdRybDKM5tBOWrt
+6HFlshF35gEX9YLrpleZfKYVJoUEgc6+ZfZaW/FupyWSgyYfjGh3I+8kIpK2a6rfm2tjY3CRU5z
3ZftsKYrtgJwYi2+0EidmZ3a4vnZnOcb5/UIpU97oDeMAQhJ4l2X2XVjDa9J4xgJQhRwkIEmcjLN
KC3RPaBxqINHoJvmNv6VDr1hxcJcTjn/4lkU98FUMPY6m68GfVA3TV2QwUGv+qlwBo+Z+R0CfHrW
XF9oQ1bMF60EI4X9dW6i0vu2Gb/ZJVCb1M0FQWgEya8PgJaLfGlPX8GZU9t+R1baCMWJEWRz9N9D
x1MI/ZNYiJEnwoS7sg9N7rLQdyU7fycVIFkUCA1DB/fRKcO/t8d3tZ3vOS5andHj9yfIUReAXAnu
/W3/uwb/IREe8yVYVVivdRYIhXmDyPvulUUGVeqs9lh8kZNl7BGUU9Efb1UDun7okt78meCmBlLB
RnDa5vSA2mijk/WZyeuiLB00Pz9GLSQ6Hvmw8VBh3TKelJOdWdXDYgGZ8PrXh4f3b98XVvSZAV4H
mBjuKG1Ng9JtcOLKGHANx7qqLH96qil8XoEz3hvll8VwSI1Shvc3ZxRtJYXZq+z6XTg1hy4zEcB3
B7BLHPkd17I9nRUQ6tczqoW3DJ9gi5Gk/PWfq4ySeoc5JQf9bUiu8/ZPuhtmDXA/HOZ2nT7/uUI+
n50X7jKza2n+K0pG8rBhKvDItk4S7tnTOS37Tg9cSJMKDKdiYUg3UlkxwojSTsTX7YxbdEyeRjLr
tPEUl2DzC8J2QvIWjVvIYsz+dXsKT5NzNVCJaBct7+RP2eRGOOQ3JXkjj+v1oNzFnL5wvFObKjBv
lonitXpcPCI6vSVdyMqdLNnQNi1dA0RZdE6VxZMtKpNZ4WlOgh5M+L/hcsp0cFzCCJXZomv8KNdO
7gNxCA+hy1YgyIlPVYw4iecg7fSFnEqv90pooQ9kTuq8cBHGrJ4n96YynMJbKDaQAHendiP0+AdO
Q+yUAvIOVzfRcA1QlBohymbwQudWVtd/zwXG26rCPeP19yYkkUE5NvtDZ1mV4AlAcaFSeAZTeRRO
/JMarseC/0RCQTayqWogB+0Wp9eqQeme7TmxhKzvct5K+TXvwPw2cs+umjiCUD84FflXo0dl5ZI8
WasMcXNi1KHR/FnVUgHUZYzmDPYga9K+cmdgHVnQlRBu9G1Y1t35njzkV5zpli51Hqp2Z2ZHVsY/
/KertDUZbKbK4ZZCrar/yTN8JTzIrCNfU5etkneZrICWr90yQ/0udID6EZ506Dnu7iGf9/6AfuPp
Dv6GGOXOqMRTQniR+g9XsKXpq6d6FuBTmN8ZmRYgvB6VSCKt7gZ9ScBYd76763xc++Inj1bIRMPT
+gerfrjWrQ2iGwt+FJ6M+W6Cz9lSkumaAkRkxtwtaHeFrwAxMex4SteXjuN+0OSjHAD/U+MIrZwl
d9ufoi77MkKNSe3hHezBeoeOEHBojNs1aIAvLN/KVoJyWx24Y5pcmMkaEJE1dXKwVmHjRqylFSkl
1WJLfqq5hIfeohtBYNALIlyX9oT/0xf4pIusNIt4T/g4WGDEYTbnaKFgZi5Z6AiE4vVYeKgBA/H+
lpqy2SvWu6qY2PUrh0AtDyPUP8AeLRLKc1fssDE8M7uEtc8DQ4miwNp6mBKmpsvh2mvWBaIL6Cby
/5+rZ3svPY7qYmK4HnoroyEGwppLAWaJg2tPO/a8i+dxJde/ZXtjc5QOPj5R0Dz/VQ7JYUGmOOXM
ns0fLJjuehFyqaZ+t9oloZSWXW5k5ZQo3lZqxHiS3M0qifR4A+WxDAOIb1SUunDw9iowXpoIx13f
UMJzP2o5tRCbntapYeIyuY/BetAALxj6q7Uboiyo9+BHYYOnGTdlDM9TQHOrPflSBZug6AZuIJip
BE262OGUggLBIySq1UmhVpjchQk6g0UI5BgWyQgKKR4fNvxEw9t4tWC3e68dflW4m9RdAAxbQrgK
3ciy/nNw5w3EV15t7crz4906nkAJmn3ej/Hb66oMxNuZw2xRHcxuC7T9/CljmJer0LmdI9U0Hf31
cDlBZC2UCbzwyB0duCu+Uw7Nm+eNDx1guwybJGMoMKy9ykEAbHVjl7T4SUbksDnMIM7ajP7kTYdo
/y/plcGUARoHbZOf53GvqS1hw1t2ntkjQf94upr9vtarY9bc6AdhwphNjETwVPbskDaliMeaOoP4
tLEjd3ARVzzGvGXtf8FHgX3i84zDtLOQD0EONepEhzdrlkBQIcEFwKWMre5V9CrxC8WmSikuCiCj
GCswcJkmCXKRjoc//rUL+45o6VP/JeeB+8n7dZ+CIiJUlI21/sMFVZy1rwKRV2dmYlRPt04RnsQ2
jvPkq1HlTmBTedmNCPUNw5GqZASpgsv3hEgUa7Hs8CzncEnK+qiOTaC/9UAHhtjc+yXXId1/epo/
J5gL9csA+6AGwg+EUa90XZUdlSEkA+e8bVF20h9S4YRN0IG6SMwn7CQetzw+6jdFE/aTDpDhXWag
bmsOBe/3i5DOudhuVCwodsXajvAFDoCDWHozl2B7tM8hXHXqaJIPk8tOThmnVAqNaQK4Mfjk3j+K
MDwG/E0Toq60UyDwJVUer4Y3v0YXGyYcivnIzn96RG7vq0xKpnRraN0GFS2DD7+w8Flp1/oUrswS
VJdDdtPBgRxHI9+f/uE7jNxl55Fu2YjUsW2qulHw/Egtm2zV8w6R9b3CP4oDJXdeyCayPLymJtV4
MoiTbJORJiTgmZtNn5DAKTpYRYcCOe8PoKmsOyda2vuZpKmZzRiljWi5cBPkMRgBJTvjE585co/F
GjLwT6Jt0/YdprkIWYTchz893HGC7JsmFk5NamDdqaF4ISoTTuJXEA9xe0PAfpPz5gcmV+cFOlJC
pTmOsrIve1HQsK0td8vz5L/A03aMt7vKFTW8ICkWwNtofh2K0b0dlEauUgjmmDXD43N6SEsUAAdm
XtGm4Ofs9Rdg3TKNmd8jTiI2rGD9lLrpVAThOpvQRKjkU/y3aURIn28eTYlyagaUwT5z8r1ZALgw
KdZfpZhYvpQqHFJOaQJfB23z7AJA38SAjCsdfmoLNTQU+6aBWPBeJFqsfI6Srvp1UMaecte2DxOv
gGQVkPUkfB2/27lbZiTN3bENUUwT+pplWBk+GBf+b2V2itXcUeDSJYXsRYZn8lMtpCA/O/XSidqu
rjiuFvg7ewVmSbL+zVdAqRZfAv3P8VJF/2uYOhzxCje2LK6AWmBuuGpcMqQU/Nu3aEZcZ7QrqHxb
a6zbiKysqwf4Au8IwbFeq4CTdbemcSlXEBdSyhqndE9RzUz6wDV04smur2EOioqrS8VIrLDLyg0I
VJwG3eAUkHSUoK+SsVYbJVP42GUu1ldNM1oeVMW1+YoEyZzpqjqSoql5x2JvQTFR8g7KjKG7ift2
ZHg3VbggxxpWPoRHTm8DR/cRcIYDO3LStiMz5CFjkZU98RBpCQdxJtxn3gSd196Est9W4TO7ByKu
xm55MPQqUUOTY510ZAfUfL3B0MqCQ5tXT0TDaphz+tXEDQmfxTDQUKhLwX/IIafuM0Mrrsaw5z4z
nVkiVwuRHbAzmUFE3xAv6hSUCLy2Dwbp4jleibhQR8+7ky87b2VRFAaiF+FbmWmTkGQHVkcejsOy
gbLM4ipGhH0W7WxJr1wDfrFxXepzFGltNnyj+/PTn9vCewkKys/zkut5rrQGdx9etbRQRpspWeri
Kg37m5CLDjmTP7olT5RRfiVhf0OFUbKvYoHwSfjsWTYo08CnWB6D3Rg8Wmn2reMgCUM6gEta99Nn
3sUN9iuBU78dV8UfDr0X3vbOOkaqqfwx9k6MeMdCQRDYv56F4TLYi8FdrlBQAAjWD5vwN3ShtVFW
Hg+yGBY3GpneVgUQAbLtPdaf5D8SPkSQn0MTzD/5IEBqB+tmgMgHArU23PxlWe1H7eAqof6kkRjm
g16ri8sdCbHy0eH1oEEA3KOGX5musIXDk6WpzP0tPxZNQLGq8vIrGGRpi2kVS9k0R1Gcwgjw+vgs
pHh0GkLiSmWBNU1zh7Az2Z7oq8t5vsjGXgM1IuYEmhETen2Oz5E4b1B1aU5aVie8REgO9KHtC0rN
WKvJzCQkStYhO9UlbmihAaJE92VwUv8G1KxFXk3M+888ScOBF7Z+Sg9BM1ZeY5njSogrDCAnGxs3
CCZgKEjKeb9I63JcIItEZSwTDtQINcdk/SidCAbhl3IGdkLNaWxRxm3qtuMdbseAP5zW/QWUUuq7
z3z+KTLle5t1KNCpvEVe7whYke39v9w5nrxAO1e0fchTrWKEDE0JEUXSlu+wZdkIwcnll7Inr96j
yABiAiHFl0iGO/Dquz2jirr6lLNZRb+cKs0P0R+vH5XRRBfc4wsbszT/zLFaEC4x5I9Pk4OPEuqB
KblZQVo3JVud728KiVLurjXXttFizNdkPPM0mbAkdRkGHe0IonDO4ybFetGZSJ+SNtw40o7s1iGy
UQ2+JII2OX8rqeX5YlHUjNMTXTHZ1vXQ8sa1y9pY1yET00wXAiPwXy0AgpWnD1jpu/TOtqGgDhJa
sTFP0hHbC+ezoSvtzJCiC+IvsP8wTtSOq/Vy9MB7fIvYsoyuygBY6IEtSuj5HSTNIuNZG0xaA55c
GCiCF87BdGjpEODkQqBKgab9w2gd/Fsbt0Z7Kk2I7tPYDBZ6Ia4Wn3khKYee35dqOla0OTC8cCdX
KLaeIITDYChcayS7gWRspL4mox7GQL14rJ76+iQXPky+fW+Cf5a9sVX6lI8HKMtzIoNkJnOGPRiD
J1M9pC+hCcYg3RCaQLksxeR59qqhKXstZwCAo8ALunDcPJtXyY+7R+ApnFgPmMuD2Z5TLXjXE8xr
IeWSHW7OmSZTWmASVHQra6pygXQEq6X18djUyn3HV6m6gfqZU1RJOpsWzePOH1VAC76+8Lz/HpiM
KYKcrEfSUx7csjy9uUpJ/dPeWoUf6OOnO8lkZVE2e2QAs81blxwnMkvUXP3YxGH2DsRpXsFpOsFW
VZwNrWVD3Hu1m7RzabDw883pZ/Be/nnzWdSbfD2YZGZNwAthCgkHjTlqhRjX6PIZ5N0PXRq2R+q+
C37eim/6hV3QIwMBEusGw2venC1dw4xFDV0iz7vJrHmsdr3htCmGe8KJ5okTkI1UoScHzZdR0Cgo
bDto3UIwkMLXftBlQ5X2Y37S5oDGb0uHXfOnUrjuFBGIDCTVXGt2VNXg3M6KyZ3mZSE/9CJs/Gc4
EYx+xBsGmNkD8qqcTxaMAPehMh0xQmlXYh02TfSLlD/Qtuj7g2yIAgnmFSFvaTavRhCUBbHi50bi
H0VPoTTd5tjGNvmMf06bUp/vU7VIt6BIqtLDOVmcOEDI//01sVBAKipat+yqn4kuIs+f8UYe1YNY
egVYxxgwq1adb+1WDrs2W3oMyLoTdNzh1nXk1UJldMPbmIaDRj3XUj+JhYoH1axCa94BSM/gSfaD
XBp0hp5R+EKVEuhzy9uzjxGVK+8j/7UHzLgTiX9m/EuJM+/R2Sb3YfYybo4xjqZKQWI5wi90BRIO
ZDsAHm6/21og+XwIxi3tAIGl9NDsxdfVtY1LuGCBscUf7O3t4vspHTj4j33CH/wjl3Ga0K0kcf67
p80ktKLsRAnN8kQZSqLluSpkHuBEcYYjsPt0gtIfE25xM8CAQYFQhk1iwBoEZfHAJEavoIrAXBI+
/lJWEh4zrXXtO8R13Cx+0eT9hixMzXOFM8VHtXwTmD9Mpax8JOFcQAzebaf9oHwYy9tWP6Fg+9h+
W7K7+LXNGOMVBdXC9cNyCstwt+qUY885H6eI9wE8NiIL28XnR7UfHV/4rLk+0uUwDeD0UCSkhD4/
S/YXkx9+YKAPve48TOaXskKE2+bViNgIFOPQhE9jALDORgFrJuF3E3e3alpWMwr5Pn6UBfBjI3Zm
QzV+lO/VyqwDSpAp647Ba2rmrGDxjTdYMpiQXC/KmVIqRV/Z7dDBUxivwiri02DgOIXzk+62gwOe
BQ2PFDzLlM0ZCjJPqMtBXZG26vnGQLe4bBP2gbaD3cdVv6hwqXnXPuxslMpjqugCyp4oRHXqxHWN
J84k5eel1nL3/8CuwAdHKsRU9RsG0n0R192WKaKdbfQyRQtTWaNgtBxq7OSjeicBUnOtd8lOaAYt
CIv9iDQLZh3XXkc46AMqRH96PrOw0OmGxdKGV8Itb12HmJK5wTTK3mqrf+HZbPhIvzXKCRL9nqmp
BE2VXCIHfs4EoX2lnDKr397F+iLLIAKawWtQWED0wPXtdqHGMsUWDb2k/vuusV6EwFZAnRFvD+yZ
pPbHTtd7oCYwHWkipRxH7uJQSCt+PN6Zdks+0ZD4qDf2/wepoGaDG/3fXpk1AOcKVnWXLRWyPvZn
dHwNoMXsBz06oyQKM5/QWme8ATCxAQh11D1DVsyyWLsVtw6wTXZyfRix2Gg6BZ6+iqx+0LvD+5dV
xWy+cftg8t4f8he4VmDUD7qooH15lkWntICQwTXJN41g801zvctGlOR7hYW/ARRrtcLFYEB7v78N
Xk8t1VRotCU4xWzsjcZ/bdhRJnzapEF4lGRJF7xYT1qgjAAoExX2Uoeyu5LTkHMaXbJ+VO869cY+
dT/3bl07nbTRyy2bwwAq42e/AhGMorJWwdSBQaXi7UF0sIr/dn7e7jSVYSsOPzITKRXB51fuAkNQ
6ia0mqNUDhSreOz+dbdl6cBhnJy26wdKos7ApSAsI7e+v/YDxlqGXDD+ucxxYObn1kol9321Xfa7
We+UJYw/pKsQIIAD07a0ZuKiSc5VI7qS10QOiVb8aEGQMV5mN0CpB2G6D4lMW0nJrjaZZgjrsCBp
0z9fSOZUvT9qh/Nx0dVPImcENvHjtgKxCoodBpwBU31xfcMqsQlO1hT3MK1EgfOFUQFTIA4UYa7u
uUNRw9HVtuMN27m4GO85PdcfamY5o++/N0/g/zq0C1sBKz0DhZinFPh4zU1uvyNNAvpnHhgdXNyr
imyy7KpgQxahEvsi64vzo7NUeoNQYxedow/tXMGC/j7PCPB7cNL99qqB4KVQ83DIDdhzTr0ZHBey
FhBU7IYd3akJvI2O46d/IifeI+HF6YW1mMP1eBDx1wNLbwIBtp6irKF8ZX7DuEa8aB/+jnlpWlSC
MR0VxXs+NsOeFhNWMPygOKJVZzeIEiJX+kb9w7FhydviBvolZVP+/pF+znIXBQdoWRNcYCGnd/Bw
2QFWXz6ioon+8GpSG7okTUaYWYXMObJrHOet0l6pDpAYulOfTn1Z+CIMwtO3kUaSSIbSP0j3idrN
spZuyHmS7/cnHiNKJilsssRgRHX766jwi454qP1hLazHQUYJPDntbD/ypKan95R9l2/JpUMwXeNP
9cL3+6a9FN69Et/pbT5GnoIiB51IytKNBEuVT24kAz+WwsJ1osgnd7GwqjGkYNKEX8Ll5Q97AOXj
KNRceSSNHziyS7zNMUgUDQaYiL14TrckfhqYgzln+9QEQXwq61YfkxDiqDlIpsY575YRWu3buTLW
Dv57s6aIUzr4UW/O+yoXsmOE5S6B+p7eV+bF8xcIs8OoYeE5wkiEeBxoyKu6tPvwhMc+7nFqWSSg
hozAXPl0GSITNV/8YTxY7JdtvQ2UJNfrlTBq65euOsYLLgUOHC9qYCbm2/b1k7bzIjmyafr1yllB
bQh1qQe5CMu5D5f6hEcDJPadvjAIhsltcDvjbhThe+FKL3lCWiP6KTkRSUhBo6EwSye3XaT7dIQb
RHBWrIA5u4nfp+afqOBySLiwdBFkMhCYHsq87ToC76PxMJuXWV6QwLYmCVm7LjZ79zvf88ekPhuf
LqNnM0TK4d4yQTUwonO5tseCf13zEHvUl8fKgZvpz/uMHcdm4kAFK5TWV4p704MGjIk2pMfUyoUe
pPQ2egOCFqUaKtMvoMCqNMC4SFWtoKmLSByduTTmaX4UUumn6gnKYhGZNy0nBTfY/M20Vf/u3Ucj
kP+DSSBtbsVwxnpIUL/xSsALCcYM+bO7KyErTeOdRyaieXfbmil/gtVJ9qQ0BccG7jc+M4BblOYt
gwjsxO9tgyIA8Y8QnUr35CSYtl05Oybd06kfOF/6RD9ugZxiY/kpOiD1VgcA5DbjkmLJH9rUSL4L
dVtk7Zr3HZDLgdJJ6/69DiyNsnYl32yauA1bSI/ySPSn5dlHKsI1NnnBpQxL8yFdEYXsVah+Vp1N
gMzf7rfbwAV4lkc7hHUNnpt8aCpOgc8Koj3lwrDYzWFOWpL65JE9ccLpK4UWjMHGq0bwIX9lCrlJ
MXjOKjEHMPgFVpPBFu061zVTEw+rr9BXFkhlSq8PjJjv0giHnWj4OW5uZwgTx6ntLTLxwDQTDvfW
Zk+ECVc55xR17w+DJX5K9p4/UFRp/wqMpxLYQPISv85F8YG2jXtA1wJqJJ1JZ6du68hetupR6pw2
Tlma/KOBA62UmXW2dsuH97xe/lbUzndRq6zQ635j5nw9GYYWKwXejEqgHLFFVhBFwDc5ZZWwyV97
hib2O7UYQdm7MmLy0BTmHSvqSuTNPxIhWJ1MkJuFkzI5oP3wlPa2WLD4UUBO35LWr5y9cMTt3mDY
/QiAVkmYXewJgO1mI/rpk77I0Jgnxd6P2HeSjSi8mFCPQtWb6h5F+YDcBdhVg/qaTUARrNu9ONbx
lkg/U/ZB2Iti4i6Vh4plibRua9K0E52SNB3gx0ly3M1iYZeslCl0TYs62XPFLtj872d4HP2Vw47A
OS85v/xVBKIM1OKjkMkrVhh/XQA+wrC94NUW0kGBrrzqpUeN+OKktJJsv+DduTBMLFbnFHflW0ZZ
j481tV4Eetr2fFN5yOoTB+Wq6IeTXVTOL3HLAo+7tANTBdiOURHCqf7YZwc2I8Z34+BkrblKz2Wk
ltwT3ZJcJIlikpNWDgZHHRhfkvsyi0T8UeHisPIi4HBAB7IMV60aiaY/fTbNbenTshhGkgarafwf
2ycUy6Mbyo18hoG+NH0oUxS/Y/bAXNTqJkKCrGx7aOZyuDfgahuR2Wv9uvzcPHXPQYAMz3FAn7yr
BL5B0+O2T3YsgEDVYTQhn1zbbpR1UDmG6WdTpZimc9W/BFLFSvmUsPI1IvQUYhn2TbDskOivcZBd
cCEPMITybgB3tBm5sfVz11NNnl/CAaZXr6ceXNBAZTuzw3iOSpLD+jQ41XexqDdhjOdIwjeQM8HD
HFLbeeDQF5kYdaf+RpbPbhsfOB/KUyhcobEDI9sUq+ejlF98BTqahSQ2OA3OE1di35xygDWLAPkg
Lq/T69qEG//QRDPnSL258Q0YdXh669ABfi9fq5mBsauyC38tChJFVZiiefkBNWFWdFhIxLNLGKBZ
q/8Z2ZqGWMrJuCT5ipAuBT38TwOwkIG1gZRyAuX9lqlFh6Nudn8I7t3xzsDQ2OicqSc72M32iQt7
vXEdrVttFe1S7Wb5fKfsSFkIbdUz0Ffjlw6C7exun6KTmXmpqxbbaD/bcF6H1X7Kwdj86miox/g0
ER5psG0ypPek1kvShvBpHpBeYbsQg6YlDoK/+7xe3/M2PLMdIdpjU9zNm1vPWxfP5EZjlY9ySQbX
Ai1Z7AbBYBJ30Kap/rtTQWnK+8wXZW3wQ48QAENM0fVcOfmmnIEvteees97odFZrK6Ijy3PirsQI
m5cLAoxwpjKlDGWxtRnUmXPleoALD+uFc78SME+0j4mzO7ePD//c6m3IwH4dzoJFr022NQbFCzAM
egXLsEVdV/Fdpl0NKi73YtaQ0BIoOGSyOSCafMsXr+MAZ0TuBX74K/dVYFLR39nEG7SGr3k873ZR
qFrLauG8YicVY9dlrJ5k2Muwwux37vlgxekbwQ55NzzVjpkW74jEhMfK7YzMJVFv8To1iEN2HGb7
fTbLnfJ0M8DAlL2twlmkOQuq+X2PNSS5J4Kac6XOdvx5O53v/M1z0YQK1uMAZVHfcFoM7DiSPoCP
XqzP9RGVXWFwXfa/EuGDBc1o+fozbIH+PtbxBcCOeQsOMpNtbmpq4+QNzvSaMEBgpo1tVIk9eqpF
UXKubxcx6+wN1B2syM/siOH31nmLubwQNGjBMaWDx1pdu7OOG95OWqcnWuyeSFdyTmRPSTk9/9S6
AljAz9IWIWp3kHwggo51Z+PWrtJ/4EujiDddhr3iZRfY9D5s3cZJhr03sbaQhgLcpwofEZM/SU8A
rDxb54TdBHYAKIjghA1yRdhUjxsxvbiY2g9TrRF0jrqH74GDsOYXdxsAFyWPdMHnMuIi4l0/afRE
Lz1m6XGBQRvc9D4Tmo0LXbJkT7d6fSyN6+L8NgQemPwiLApDJTkOYWyEbrBe15KPpHumKUtoJ1P+
5MBu21HQm8uOYhX9YXdh06/UzfyCbCoW0VmTUt/6ZfCGnCO0i63iCalKR1rvfLLXPTIwReAP7ASs
lDkjAC1lxcegJ438uK3VebHdJJ2LNyOYIOD7/34iqyNSiTh7CFAapErRIlGbaDXrtk3INOPlplLs
zXtIif9bwqrZ/N5tQLL5FmTuwYy+TNwhqIeARV3UJRInfxy87ST6t2VvgUisUkdg8hz2BPP/ZFBD
A+aCxK5bpUs8G1gN7voyXlVMp40g9coD7WrxITrMxnpSP8OqLCzAImw5YCNI74vms+ZhckFkqVlC
zC6rlNP40FrDUKf9p0QKgtMWS+yAuOboduKuRWABnrP8LT38ae0+v7nnoqRSKuppeLwE9PNdWJFp
/efHfmDt2dMKeWHt/LlmaL9Jfw2UZ2ILIqGQNLzoE86KKB9o18cRflRh4hA4t6/PgcHKNK6LQRDI
Q/7JhF7wG/HFGLSL9tS1Q69bq2x0QuprLPw4rfR6kc3brMZQyGXoFakCNAAntiCecEkQJVY/HdnT
9Rb9I5+kcBXa5tz3T4abbvD0HFKVadd1WWuU+FWpAmxqgOWTR2nrTAQ9u8rPjyjgGPDqGix/MqOn
GffNmgNr1i4iwxk9pAYmjfDc33nZNH6QJ1utnJeKuJzCRg4fLsgXOsOUlwYlM8jGMQab1xVDZxe+
uD3MANT79M0f2BBbaHFjXSkkkmelW1GTG+hh9irCasi0wq72HJzuQc9tbbThRn+v5hFxwQCr363g
l9pBQtdgItxsGYZhNWfnTsmEEU1yJj8f1O2HUUr0OwEpM30AZKOp+SNTNKScoJOhlX+P3FNfugU2
hCSr05+lwtBNXDbUXeZRNj4n499hP+MDrKC3LYUBafSb2E7Yg3x92rdw1SQVoS11LdMMP7+B31p2
V4R2JYgeRYT20bKaKaeHIKx+2RwX9c/1ZtmbisrqDKOS8We7hoOPBh66CHjScyepLAS7Fkx84yU1
u2zzFz0TOd0Y+xx3+wqjcOHpAdRearA/FIWOl6n9uxJAS8KMaBm9jXw77na18BiuWmY7bQy3xZ8o
0hZVPLxT1KpP1Ui8Wm42X6mtSx8pzLd6WUsYVYXJXQggmEDCYuWtYom94QxRmjQwrroFA/egleR0
9WUWfBC8sHuu3e//NeZFtjQ0zOryJ58MMtAUNQ/gmaFeNWuMzunR9sNNOJV07tCfI5ETPm2AZ1C8
onmNsmJICbx9EqiVgqQcyHhMNtDA8TxKeU5nyoDQapWMWtOIMMDIvtns0kn0Y8WkXGCI/ZlXAJZC
zk4nD0opYLDox6+Fe8ncUN7THr+tPVY9/Q5wwM2PPhOahlH1Axc6MdcWmwOC1RQ8/6phTqdMeZiS
IgANuW/EUPecwQxVCdPqZV4iyrwaI4v/n/CmxUfN22TqEhF1QbxVtdogS6nE6qY1T4Q+mDAZ7uWM
0rfErXDZWC7kbeKPGp8gdF5TMN45KjsowJN6MdzhSPdGZttzDxdk2l++6fQZaPS0UcingvIpsW34
031j+ZvspRQCfUstj/d6UbsfPLcU88cWAAPHfTqYJwo/Uz+CX5y4/J3/0I8zH4S3COOq/3QiLa8L
ioFCQIUXcnuW9lleb9ft+0XvU1bz6cp2DDkA1VPcMFc+JdaYSc1hpSMr1j6D/DoCXCB/vOsjIBNY
RNGFjPk5iJf73nPwMH/dr9s1VmSOMSJJlXgTIqIQjLXTw/kjCIzqkFlb+dkRYzgDupZ4xFG3vNKq
WfV5LJVqXeXaHperD8Z64tPNYfG8zThXUzpEzItDwabCdokG0gd470nZbiycu4DeF/TVuq3MxJZg
gA41lMD5ZpH/4iD/pjMXeZoSjNQ77momNiMkdGlBGqFrcXSRsOaI3JZch0weS1L8FQGCd3APLk/f
HPs8C4OmKLh97UbCuHKcE0wKGmRWeBSME2OJyWeO0V3REuLFJP+a7IIlnY9aCszYMUbkJ2KwlNEY
m4oyHAEXrm5xKCJ7SS4oq+5j+m0RT/bM/bqs44ofG/z9Ex+hqokUxmieAbYCp0gARWH4fGSpwYlD
vZ36gsDAOiweZr0h4rR28TyAo1RZr1XVhMIct/0lTYawhA+usLBLoy9h5WQT+rl3qpEzJZEHyY0Y
nzkvxer2nXARUh07wAEE6O5uWIeZV1Ykja8Zexk8Hws0VtHLRTnFuPChLhuQItEz8gqwaFxNCy1O
XTZLL758zw3aI9LZbhdRzGtmUJbI3ik87+OZAAzgjCB4K7eYSOPf4j6kOeBTz/g3/pT4HESEML3C
gby+hTUSmlckirRpiwKT7zhLFFgiNsTfDSswGuKGIoEbpyeHSYKNGSOMaOv52zszq4wIhYibdZVw
0kTtJf+AfofGX+9VYAmypDB8HS3q7JJ+gWgC3+Xkasf+lGiWGmhxuNpyUCS02Dcpdg77ggtBQ6Lx
ftX6Il066HInHeK4gU68fi9h1ieqMuXU9sebEJG9onEkKCAb4s5RCleJUcOzrDtZPVdRzrMCgsUn
VuO9xNNbIP31m9pq0+I7hyYeLYNO1efFk86thzoiFa4V/5t/9fHn7U8Qdj0wtlVE1wkdT0SAKGAK
CLLrk0o3N7psC8Cn40uKKbhm/SJdvMpxmUidUIVoA3B9nfSiALAzV/5birAo7IJqxMH+oZGxj+YL
s6SygUs49p/R9YERBzVlws8V0FOXyVRDffDQyAhid3D8AbHSyjtPer91Pe7xB0/wdEcxkRNEIEnb
k26JPiuRsi8MItxnZTCsHIqBNCmmu6Os2ZJvYBHAAEaujelK5+wNf7+RaYKigYuRiUQiMCbOfBjh
sGCYM5Q6TJANRGagW6skLd2vI3y3UfxlM8e9uT0OqOiKktLVUf92dtmaavEtVFmfIVmWJozQn8p1
KmGroCjFC9s8SfowCbmoKoLn5BKiCaLeOc9gghZlvBaCUpX9PqldolBbRwH4rmhAXJFEAFVZ3Ut2
1pBeGGPM/bswPOZeunqzeDMRfLUvOSZtKe13XQeUSAUtfhfXgEsSEA4OTAvYdvSYEX2nZ0iNSxyD
64fOYrwJhDwMBoIKSJbYCA1iVVomJHoxR5mXeT/+knosyLg47pICW7nHIZIkuaz1NaZn6GxQYEuL
pCmoXDDJ4FulSwKpu7hzN0sQSoTrSq1SG0ir3dbax1hftdVwdzoWzvLCrnhNt0mn5zkzt0eV7qB9
qKURcR7EeUHPZYi8Eq71z1M+mKIjp688fNInozfB77rlmEA5TKnmiKqgkGUG5MEN51ep+/Kyu0uH
J8Zd9zCWXHsqyiB2iWRU0J4l7702CW/A7YqsSg3t2Al/hwUmX1/7++hIOiH2zI42zL72GvNAbFmo
jWSwSFNDK17swo9bPrCZ/G3rYkRXqZvU9fsrVJlDR8ZHBhpA54HkXXl1e0P5SW+OyE4bDDne9i/o
Z5g0T9hoqNoOMCbVJ0dN8E66b/Rk7O5JCHBYDj8B0CU+kzq+eKQ3+9Dzd5FhPGdf6gk2ctwI9DeD
jx4DZ3uLnNONO0Z8ZtaJJbn3CU9izJhRlcnZ8aPU/qyatgCN1BySkgppNNinkO8fjJ/ThAsmwLVk
UABO/T6Sks08chK6ziSS/5SxVwgCa6DbgRdktfykqC2C7PTT3t0z613XJq7byzhVoLuyGQDVOsIr
cXPlmg7VeHHbAyH0tkPi6I3xP1OZR1Rxh4Q6L1Iz8LU7IaqnZSoDqandvfSLNQo68C2EU0LTdEG9
tD1QXl01mVFS1v/R0aKsycyvjoSL5ooNM89JBSWw1m+IwH5+RtYdPo0ZF2wrzC9bQ/yCJNNcGb8Y
3tiAfpYL9OPO6ySU99jmV74xJF+iwc3oz6xc6gstFxyKtnQE23PWMjjUV32Dyo58u6SfloFjmp1j
WndkJvcb+YjAFQ0+Ao4rgeLCdOPhj5cx48ixs9eMbgdFO3BIsZhs9Fid8vAPyRo39R1biD80lAz1
vH1FwFiXrWzoTZgtUK7FhCCmpDh/xam5uSvVTkigX3SspVtS/YXO+AnUntNSlK8XuSQJnZB4LjvZ
OHG0Sc5/zEtuMkdtujVPtIp3xjQFeIknEWS20tELvJ7DiHV8U92WDtIqahwkSMYMHaXJEW1MTLIg
LnJKrjSuiMm8q+OjODgR6qNbDdPRb+xIY05cPRcc75p2qWoabO05wpYZ4y1jkbwlDpe0XOox1Mzk
wu1OJJVEPqiUkObG6VvP6/RbAo6/9OEt3PU9FkLuukzXl6K6JQ8uQ2QW6ZrgY1KDTp17e9ZeL8pO
ln+cgHTZItEeRVZhTYx8Y8Zv3f57ZfJRpmTkByRgJh+/11giI0w9vEVu0UHejdgzw/HxLtxFj1/P
qibTktWX8ijGHNP6AiM8wTYB1B/2Sya/shhVtsylKO9uNXuep906NDkGG6PhY+8IVUphgVJWBMGE
4qyTaKb0yPZ0rFME4ngc9ayXExcHU2aIqthV6Hg5u45Q09/pKovhO+k7fOyJ7EbfnXiGDh1IMca7
sbZcjRwKF7lmBTdP/z30OOEqBFnBBnu3lALyWXIc1d2akXfxmyDgR4Ng6aPUcvYvYPViymsxTTY4
5RJfHypVNgfB/5HZ51Cn+ojRQQoOZp+K/n1mKQOPZ12mpPwkr89C71CmO3FQFjxryGxOCEzbHZh6
DfvQ8Kz4IY6A3KJCaRM27VOnHBdJsI6so7GC/SGD2luOR/60lqbNKx0BeJ9pR/JoZQLtwjx5BG0m
JIGx0Jz6b+E216j4zEOd/jGp3hHiLYQnicOaUW3p7wjEv9Az/q48W7XrDjbcPjIT22qnvPsERlF3
3b84pCx0NmqcAMVfMAZXsUVYN2QCWt54G++hFWuhgjddq++jGqdqQ3YVRUyKeldMuSCsjBWCoQdT
czce4Y0gndLDo+5ZWMQjIRzxUUvW/GyBVLmuZzQlaa+NTWDnK9IwtgKz/KlrxlQL5vX+lWzw8LAC
+P26sbbcSy+xbqDtGDfQb7io+yNwgLbl1HHbP6FNLwPaiWSz4J5h7fonwGBK6wsKRgbsURyFZ9+B
i6pdmwpT4t1zaVfK3XbMfxEyNP48gHAutWgVemehwbYTeNXW2uaARMD51DmUeXDhdnWKWpA7kAJo
x+j5rPK4x9Smi1o0otxZ6ed265m4sJaAI4qZ9CcbBCPWH0diV+fiyVrOhX9b8c7Z5aG9fBRCNicw
5y05yGIP4cza4YEKJo2LuldcWrp7aoVdeWBzqveQpQ9nXpLCHL84wfdgSo2AKgqDONIGaCeJvQ5M
t4SPFpDHkMkQIsgeZ6ZgYgtD8CU1gTYeaX+rtBCDAbm5UiNaSdZBTsndl8JnCmWlksiWg6hpxR0k
0QUHIqcBqhwjBH8dxp6O0r/gw41T6u4vC1ZtN94Vr6wyjTi20AEuW7Sx8SZKcy/wjcVNBR9HAoJN
weWN8g4uST9OtijjWlDyC8z1RKJdY3s3vUFa06rln0EeJJev2snnE2I9CLBdEDhT0IEkpKcOrMAo
4ghyjUdty/HR9ErlDqRgFt/X4ippEu0xzPz0hQibUQjpR6ODcV6Lg5QajM2RD1XluqaRea2xk9Zn
h0MwWb5aC3CVcCzhepyI3dVeDLhqW/W6A+dO4SbPQfotwNk329uDH4RnKh/FOnlkNWZN5ZevZSQU
FpV7uLgwe016yYgD3Gp7//f2XbGwU28iHSj3lil+4HNTrtFzIiTV6CT2mEZfuOSS5BkMHmJ4gpPK
BVzlp0E2bAhTmfz1VXn7J1VkysuXLJRHMvLqsEDPO0tBbrLD4SEk7m7JUm7WuC13boaF7gfWZNaQ
uw0xRqhBMMYyoE3pF0F2eEU8r6jBndGH+saymBIJVpW//4wENFYXWV72ogiEuwHB3NPb1foqcNy/
K9yzcY44zfXSVobAuHhqj6POIys7V2g8x57roFL0zTqXk2g4uTAyMf1q5iX20HU6JA20+Jvu46Yb
hceYWmvzkPlPEDyU7yxu9zFBUlsXccwE3XnhJxAsEcVJHI9tGLFJHlGDJ/nv9RIycWuxrdhH7+6l
Dl4x0DiW9dldgXBPidI+UlsAmPCSetcNfR07SXUziqSkHZi7lpKLJWRlphqOuQ6VGbgSLrxK1VAT
Bt0wH+JTw1JvFzyMa0vt1rv3nlpyGC44fvyOe2pG3CGlbmzzbH5dHLzY61i82L99I/+rwUnEmvZz
fTKzqAQtxvanU3/69S25+mTejV3dOXKr2qFGrOvmrdFk4JjdKFYKtE4+zoHLcpN5zNARkH2THRdO
vM414c0YFmjdqZ+fB4Tkdmhtko7X2dOIDZ47eVbzokpTe8zRRBNT6t0OwjkGvAeB4wZbsVQeKt51
LzDlJI5iIBMzQvLcjpV3+ZD4+/vTIBjWPtlAwBtklzK+aIrZaQbR8BBa0zEa2Hk/ywFIIV3VNQZ3
gQyLZKg/0w0k8EQhkGPJ4onuGYbwfwN4oguxxqLdnkZiMMssC3sQR+Z72fB6im/5KCM49zAqehdu
mp68035a8+5kwddYhU4hXuctFhAjg5Smsz1jqnKDCvTC4VeHoEuk/VUutbOEhoJ0c4zikwnpreyX
adkna+zdwbKg+fRWh3LeTcz4oCN2p0XANlI0GTmn9U2yX3UaNij88UN+D4GGk7Ot508zZV9OKItE
mPNTo7Ht/R0Gh2yVfRnY/N5iDI0QrgvurcS6OXJTte7CGWwrsQtjhtFTF5HehDxM4YdnG2DQVYdN
FJTS1i3VdsFDm6IYynE1WJKiL19a0dBklrLvWfGUg1FpSKNAuH0E2bsJwniH1W0rHIJFv7u/MQKw
piCBeKoc/c0RRRGHQYlL9g+GAOi0dJLaM8g5hoDBOmxFVLXqOmin8skGTNqQ4nvfdmVZqvHymWjO
TtiORU9LtMVL/0b0j0pkNjP6mDKL0PbPeCGPh4MRl7n9R1KreL1LE4S7ox/8XC2HmSdMfrWI0BVU
0w12ImqjDLNXLZBCd5btEFqfSxu6BRbDVicscySYMEobkCLhbOz/MJLYbXNT2pFrsjdsHZ2N7xhr
rNLoEhmzGIOMxNEcGSd/Jwmu+kQZyYgU1YJpf6EeInAIV/we2TTfYQB1BxMKy55czdMBSkhCPmNN
99YW0St8QLUUWFyEWZNFfAokHGpPYNGZGBE7xdFq3fUXsK1XNEGgiPp+ExWSKPRzp2MohIDjHTP5
BZcbkz8nFOTSnVNOo87vO1eqKpZFaXgZYrC2gs6ED0Fl0M0rfJJZ7zAE9x3Q+6LN8b6tZyzmabFy
GEQTtCUJVOS8R1dqQuiv+Un6qznpQMmUTFxm1UtdnnmGLzd7lDg7k5enQmPZsDQBIOcELDVI7nYC
UOgB+Ce52OtW2PJEnoP03XQLYII+MsRk32SQSCIs4gSSgSL2W1wg6mm7uARSN8LczRA3muB6jQt1
xcuS9mZBqU7ROPzW6OQMyCFF1DvQAS1RXs3cGnNoRWdb0M4Qx590L1BGMUL4G4zaGLayobvEH2Bd
9f8zuKUF3QZfD6RbCd25fYMXEw29GQxj/y4wkOt5qvCUb9DFfUwCzq+iiIRYOpzzm0ycDFE70OUH
4XGqV4YEWkZG86JNH/XlEd7dt1AfL9i2QbN7y2aLKwCJZqgMXJqJPlEaixPItpF4pMdCuODxc5qI
JxJQERNUzpBZ4X3gFVWEy00g/TS7u1ZOxrlB6kWsmqSDZkJhZoP4cDMgEK4scYRloKdOY03ydpOP
r0LsQYQshthRwvNeLQlEsIE7WWKqpjWqDmZjxPbsFVWCP61b3gCqqopyKJ0b+X3+douH9+mDgr57
OoFXy9YAWOuUy9jVsHzFIV7RhYxsVZ+scP/KSF/UgT18cSOy8NRp3EW4WB4Yo6ACA0Jm+9OG6U6n
zYcOWrJdliJbnq0SEZaJTziUXnd0ww7lTzPUTuwatnwNA5JO3Lg5CKO51rwS+yYOmcAbfTBMhydh
DW2gJxqa3x2dkMrD8jAUzbvRfxd/KYs/RxE+wi+YiBo2p350SbKJNW7d+fqRvzaTxRRzT4CqDmr7
nQMqZriv0HXowZDzC3W10hiOPEj3Y9jJJXb7W1/y41kP07HehHpBxrZD2lYrLGoaRPyxkIXF69Jh
LMi7Ngv4L+uWE3T4mgDvvx/+K37Z9PRtZqFU/qKHX6NX5JVE6xc272KClVgonakVZXSswifDYdCn
mVA5YT4t4hzmWtLU0u55YzktZhPtm4hu/QQrG6K4MrdHeXeXvPZcyjNhHtQiH2x/JH8mMurjkumR
kUqXYCi7pzyCjnLwJAkAAEb8CF4kCxIKuiwlCbHxrufGoJypyBxO95J5UA+0F/EtW215gM5SUlee
7bn8fHhJ4qwEPJZaCXJKK6BIzn7lRcbx1gsMBTiMHeesRqc1he6UumDT5d8dD0pyOPY+oDoOND2T
eeoD+vHfQA+nYbSfy1O3tdgT6JkDddGe4IRUnITA5pxbEH21cBD/3rBvc5e4oJ6u7cvaAs0S6r6p
lAAG6hkDR/DaEc1Ymtx3VwNyjQJjPQL5W+B2hqEhsx3KVm7pX2XIo2cIAnAtPFqwVqq4HHBbOu3/
BqHMEc+fEw2At7hld+ehMmay1ScGRuSO5i8mWz+Bvhe33PJx+WCzcJKRmvNwXaIPfQS1TDLCf9zr
byR0uxXgjFKqBeZ7ZNmPq1VjuXbQ3Kr9cUmu+kv7hJanqqWr3FIxtJ5sMpy36Dfpu8r6UrulRL3x
8D8wUZlGuqHX8/J4OonOVGCvRrwbUOk6lnPbMEyByOqboFMhgXLgTWfc73RHD14HvJFhZfSE0pGl
b5lJIWYQSO9ZVer4u3g7bf/Z13y3faAa+H376fYhh6boRs2Vjx7YohAo5keXYich1cP2wiJgEfO3
JUDqkEOoLYYfEG87IQdOKlISgNC4xQQoMcE3CCwsKSs3nF0aactFzVzW4mhGg+8Y3dGc1/O1R4ar
xXbsPmrxpADm+IVXoq9osF435N584gyZJkUSXM9B1WNim6CAqI3wxU3JkfybytqHwMoHnQrglEKR
rIzB+24+tTMhAA1CSefLtFNEiBcz0Z+jE88vF+RLQjUXzqbL4TZz7/Fg0oSyoiY9i8RFB0zjdBM9
mBh1JXOFt9FqbEb2QEKGJahklFhDcU4eXaoQK+u45Uw/TKqZVwyA8XB9J+ZV+s0SoCMEeviLLMJT
I/v6aWg2zLfskyPIaQpMErRIjx+ONR19RG7jGgb7fSEDaAY3OqPG/1bfZvSfT0ean5ChO80Ak2vN
R7EYZ4rzniZBghAq/xHfm3ni6qSEAoriuSwrWDlZlshY1gQH+cSM1A6xlOak9NlQP3heB4QayDtg
HMNlqNB39H6SNrqTlsm9eboWSYrFkJAJwx5/+G2CxtBzFPGgiPmo2t8U1AOeyR0F2b+I31giQ9ka
GWVoTzDGrt6aBC44ie4Z/ndlJZ3rt4O+vjEUwPa/h7u9TOYmbn1/slOGKrMec5x+/mUU7PKblp9B
sQPv/F7JH7dSvsXzHXD8xV9HeLp8ShfELP/9Sm4KsCWK0wjD7OHfMKHKvfgnBe5sF7f9SA5Qg9ul
Ce4m89+rYjkEckIpzbmN9oSleol7KtjhJjmw6f1lz3SklZMfMjhPBMf+sFf4NX1SuYQVGy2vx7+H
lacT0vhTMWSnJm6Zf3U9yKesVCtjswQiPfyZR5yeXLEQsZ8yTAKCdl9LlZNqiOCw2wKGHl1vMCE0
I4lf2jlEAqZaVy4oyVa5sWAHR5cK7n/NlF0i30F/WUq4dLQ+t9kp3LGHcA/QHK0DL0inf2Zp+k05
o0pEhGnPului/grC4IAW8GkC9fyxAbRu/BWJx+AoPlAfFf51PaN0P3h98/n9aMdCxt6aDQ9gDX+t
3MfPA9jWD2g7c3WBVDObH3c8opmM5f0+4SPHXwqdoEhgVxqKG9F3r9VUtO1WQayAc1rAHju54w32
SJmQjYOgROGlMvQ+GC4fiHaumamFPGCJkOC729Gs9rHf3THMM1CSIvcSUw6sgT0XO78uh8r0JasK
hctVMqova0evr6Qo3YCy2uKeZabTrFadkteYFsAmoJ6EQaOs66wr8sGnqmF982hrF0lZXaWULBDn
qqqfBgZ9+GNF5+hZzxB1P0Mwceg1EKNcuv6wCd58Oq2IKzcCCuSRewDBl5lP6sZUldUMKnOUMt9T
bmXI4xjUXwDoI02LRUBT0Xd1yvsGucgilPlb23zLR1UAeSamqvX0dAp8dtR8GZir1NhA7J/JeWB4
amax5mYVxQarGl+DiBNsgqgm6Jo7RZJZ9vpqPFVM6obD8EchChwMGJEnDlzb2cK6MNuaXdQ7FVHy
53o8KnqhRsiNKPE8gWWaT/Hd1Pr01mTX3ngXMLZbaX6hdN9aiy/mbHSEqmfGIXFDBq9Ca9LvB56K
+trCgKdTiq2fc1d1B6AqxpFHMPho5nWuXbkL7+/q8IoFGF4l9UBh5BJcdWHE1WDR815dILQ5Vnkd
CMkmsri89FtytwF8U2gl+CG1XFJH4mlEPW9gcbrngcRrIToVXoVQYEFHmFIyiEE1nj6ttIgmqqg0
6A2Bcf+n+9oYWLOl/offY6+ROOfg3AbJHSPf7fsN8OYG+yU5toSP35byS2LD4jKX1P1QZWcj4BSM
vaOW2Zb/Y/D4aNa8R70Zt0T5/MMgZ9v62tXhMwL7KZ7jMXv93uWSY0XQ0c3NbLy0p/GRIMjXhTvH
/0xulwGmd+cSCNkg4z0ywP6ERj+wV5YGfbCkBI2ltt/voCfvGfdDCnavhJ3CXSVaaRG29AtmlsbC
PnpzNAIiQs5tfjeVhVfRATCjuCB2oZh2wvmIeoOJqGSUXOqK4yY/BW9Ojg7zMu4cPO4zWmZayR8u
sCkMoMirRor3Dpv3Wtam+3GvgOyZMfhBuNXXs6NUu85aTMKYttSECD0tZoeCqdjdshkf4bc7RGMf
6Iay0/E8yhanX/nVxwdsnSLgg9CHoahPk+whEN9nsIBl5Ye3WkeTyL+qJlTL5BnPcBe9XcFFgJfY
VvB/ndyXCkVcwTBHfdVYYegjCb+HSGMTlDcQnQaT70MbQhrV71fsXbS41tra/mDTcSEX/Q+36THt
0cJFFdb69y2+fZys1l6CfZvfGzKFfCOk+q+LtUdBKJISC27RB3V+aZ1AN/dS2tw9eOFaYxLT3Tvn
6k4OjfePP9f68XMU2O2et3AP/urPB6oKnwsyBPGOsQ5kBJVTuxaP0F890Zv1ByUlnuW2bwc6wwxj
fGMdat8gLBxtLr9vm+tM9m2ub0t+2eLrDo1Gh4SH67z1nBTAfSISCwI15MrwXm/b/9X1bP+YqHSc
Vyd7JmKh0HSw2TnTFeCQdBYcHK+en3Abf8UoDsEXhf3W67/FcWF9Jh/KbQX3Ey8hY2BU5DZF/TCs
Y4WI5FpEXlYtq1Z5l36OqKQQvlHOGo11uTTh+nrQCQWKj3vQ1yoSOhQu7SimDSeJo/ydgyOicKsN
ZFV/6EZ9wdPWJWWr192a1NMybrXgSfK4cnu4RfKFe6GaI0pBG2XydvBrg5nyQNhh+vWCu/4GAZpJ
6JFoO4rgdKyhCGXo0VA2D7OdyyRcVf0JoQySCe9P4I30KMqrapBfbZ4M14OrCOjHqbOVgr4GoTMq
d72AZOciVsTjCDhHNj6pGd64M3cw6+N+SZMtl9TuDSKMnNT55UnoGh71rYrNvp4nal3Qm5r+8Oo9
haq9CispxTsly6b8GgrlnPbdyT4kmMlqJpEdcSLSO2KJFOOtdW5Xu4Kdf7VDmkMoOpFl7igInqdD
3IKVGdZxUfc5uBMpWsw/o2gMLNbIUvKbSHD5ob8g4KNmcKW6KX7TH+DsrfAVlEjgtMN0OdVsbn8o
HqBRDFwT9rR6XJsZ4SECwH36TyGRfuwH0NtaE6jxG8IkIz6N6ji1MbtOgOZw2NegBngeJlTmqqK2
6/aKClLzV6A0xT68lEBnknMUINWd/w5sKw6K8OJ7edsgywEcy0XA3McKgbFhIzRkcUsNTwkoIPOo
o7VoUHYDFdWnCmGoN9YMcYrczTaIZmoYloCCveFUz7ZBAX+5/yGzB2S6aWC3iG3VxKE13diKHcNO
Ad6tDq1ne9yt1R04XHIjHwISTMmOK1oOo+Hapr0LSduej2tvv9+fWhDJZfiZ4Af1UlieNutf5er+
ZY9sY0cAATTDizTvses8ADfy3TPlj8J21KgN12XX7cI8fHRQbMDFwM16rxp5hwgDvPF5JCk8WDQT
6azTeBU3sVZc8cGtCyF8G6Ma4y95avWsFBdu9Z9zWfxZGRP8QMm0uEz6HXvKHWUR9gB+De/RMPDh
EwxA5mAdmBOCKx1eAswjAP2lQsfwZ4e+bhLM1oOzOatThB560MaYj236FJ0QegxPqw3//apcVNy6
IZlodLR0AO1iWmHLLQEblnR+srJXCP1gdwc8SUqkHnifozYZeA5fQ+qvgs2GEvx20GZiA7acDRkt
2Dy9SUX0DamK/qdXogjI15O4VYXU4r8uh9KK+blZEmCC3XH4Jd6hn8MNtalf+1OIBsGbGRJVLBo8
uy10jRglnkhDHCoic6mUhLwpEuuCU71MJmoFov0vZ2w6BnHu7UeIeWvRD3PTqgBGe9FEmSkawUH5
dlucLh2B5hC5fpsvlbcCmJwLFhULtfsQoJKU2uiBvtimOP7GirvmJIyuuz57tZQGnj5hmAvBCuMX
TGLXrSlln152e55YQHZERcZ5ATW2Ii1siwVZoj5xrAhsJ54+4+ra1YstIXIdrVMQ+GYrCmX+4JdD
NPVNXLPCWUW/03IQfavG1Vu9/W/GhlcRfn4VO2HX1KEVi23zKbfb7/NAcKuVgJbgzC3bA7tQ+4AG
6Cu/ltNozQx3Xq+VzmTvyvB7yIebxtiNn1OQPhV5N/VLgLzXWqNq4wRIBTFG4YG6c8GhHOM1RzS1
pGy3vYoVWlgDwVvdbjaWnFWcKgE/rqQNqC93/5KZrQRcLsEjn4dp5WmuUzBm8fHHCA56+t7xghF4
Nlcz8cNoFifUaHkjCsXfi0YqBBWmYMyvnG/uU8RwLHWtBOugv9UVoaOtr/pLHQr9AfQb6DDZRtNO
L4ly0a2NKmQKaUQXMsmtd9Q3TPrxW1phLbJZVoi7MQi1TTcZDrpwVJPH+y0v7QCISUbcDkO+lqgi
kPcdr/I6s6Vq7pVaFQPbjuEI7uZl+cxkJSr5Z+2UDHp12hX5xeU7YrXuSb25X/pLnXGj+yPpf9xg
57JS2QoNMiH701Bl08pBcmOOT0FULcj+SXR/kiboFBeynP0psi1Wh4nmOIzSaND8JntDIK6YXPII
a2EuDadRtkNk6YszWpwc5wLW/USRreQJR4EIXUuwTuXXZBHPQvJqqP9gGhFy0eDh3XNV6nAyoWqA
DvbLPFq5Wx6ul2aGME2G1sulTYpa8e6+8DkXXVW2J7Eu8YQAqp6RLwcheYIvUerAd1VFPdRD1LJf
Nmqhx5wrzmc5RyvjDRc8NKFfqokx+kCSWzM/0CnQeNrEEao6VSVr0B1gKxhRpy3NCn0q8nXyoIS1
nQXqWM5qHo6agrZH+SbncybuHJHdIyIWcX3ohPjdN49L+WuEPIrOnaILv/QK+EzRdEWfxb9OkmbU
UPaghoCKK5Ktnf/p/rfhgi8aTIoLMmWMfaUZpO8A6G5WmYMNXYh1JeE8brY30jsm71+Qh7QEzJ24
0Cfhfxc1WDH4R8L9Oz9Uy/OYn2n+AYIFG0ARDEOyEexKYMJDxghryG+bZUk31i74NQYz2Ep9yV05
BOqdTG3NQNSzKvyWtRPSAs4NgAOhPuJ2itdpDqFX49NH0ID9ZA32usNfgrCjXENjOrPe2MT9djUf
ZrFY4LZWASqR+8LPB9sOy+xjhYMZGLwEmXoWiEZzW4Wr4vFq6Mz5yxj9hQX7IxamCX65mb+DlrJK
2EOcbVyVFg7/ebSA7rfmOX0boEzTqH4p/tyssGX5HBoKSHogciWqquKtX3eiuDOiO6w2uTmMNbY6
BeB+PwGkJoViDkevS1FnZIz7qu2SPIO0AdwbOlPyozkPG+WiMnyuI6abFB/hkHHDjDzcvpbuMk8w
cFjhXxIKcBiZXr/Ebwa6WdrwnZuzWXqDLYcxrYSpmLWYnxNsHzmHD2EpzfFd8mSvMc2QFlGnUgHO
26nQTJJ+96VXDwzcCLdHTi5dkk64VN6DTia39c/4qe77BH6dRhfqCGMKgBA9rU/A043JT7km2aQr
pHQ9R34Kgr5wTBgLdVTAfM1AZHOVDN0Fmj92jyaPwRSRQKt7keXXTxFHbm010YntZ2GQqBJy9eiK
jCkKdHRDrHmSrrBSGHKnrD3wHbKGahpxy1lAsd1f/gYGBYIYAK4lwkk2ARSTd8eyD/VE51DItsTB
zKqghQ8LFKEnSLELT80t/xAUkFz4E6uy9CNssNG3vJzfaPf4mcIxH/blmV1JOJscedy73gWidcX1
620u0i8qgvYeUt6zfKHbLXSmrLHIn/PU8VcosaM9ZmSC9fMZL7AtyyRVZcKmJZAGMVKtUQ5y+MQa
q4VSCc7wQOM6qDMGc80L3uVoxkjHYhU9gTzE7rVNTUPHvyk7bkhlheF8E/D94ZGduOnYZiFdaWTG
GkTGy8leXJtP6aOGkkydGCZVC4+mUiXH9mrz7Tdj8YjuMkYZ53pUyfiKUzocUd5s6VT57YrAg8N3
rbwKDtYQjOJXvF/y8NptdxXa2t4DZPDVm1CIWpzYquduWCb7J44EC/tsDN3yO9sYvVBlAC4v7tgR
XTyhdNCGvHo3q3MhrwWucks+YtG2fyAizi4HM+Tg37coZeXOo1C+wwAPbyCdGthQ1mcOBhq87+wB
1MUYfGJaN7AetOfG/UNBlgfCqADI9P362kswwTPrFLkyNM/4bGz9h09WClYrgMy7H59vTSZdAMGm
rJSgfOPhdIHhctjPzSCTdkoTn8j2rHetWXMGKlFR+XaY1vuStU02XvQQBP22LCax7T8BAZ4tBg2h
s0kuhCdzT6H0VQpVydytnMnKds4/EoqrSlY+07xHsWiRIUlxQw56Yj/5LLks7L+HyfWzkRoeUH1Y
NoVZkwdhQAn9MOVophOU1T0ORSCxsHAyF4Gq/bTaeEpQoS7WznwFaQr9O5Pl3/lKjb3eb0SJooaI
rXZEYiREffLPId/4GCEBk9XSKCTXh8ggFV+d9mmPRxTYmOtpXO3lUtdxQ2BoM21/r0uJDqe4znI2
+1RySliQKb2yf2FPD664gZ+VSVgwGGiaBcD+ITNYHlPvegmqU0U2+/UF/93u99AbvqQc2pxglCBg
NwO814zujQfh4e2MFVKx8sid5nDCBGIl3Yf68V9O7hlNzotEWAwd+Qs/EgLooSLsM2Bvlj2rowlS
q1Xjki1FR1AcVIYwS0OYoqKvBVy1uhCTm1Iz/4BM89gfnfbMw71HzCaD3gpLcDY6jYXiD9atdSRr
0NFyJFv4qZY0P0ftVFMHkVKPHoHglDCCwyFn2bOERUHUwPiwieAz1yUFKn2PN9ka1ODmO4V41asC
9vlExsAQMpihxGYcKj84edyItsIkSOJs2SJNe0Fc5Ju2LCVgaeJdia2XxkjRvqDWS30R0Ers1P+d
bLNXubvL/4iYh1l4jkJnPxjnAbRuzq6z+ExRCC/bsXJ/cc30CtMbe3l2TYd4uAUZ/d6TPeaIfYnF
hQxutxTuKyuE1yXxKEPrBU5q8vXcpjuJfDv1tvkC9tdk5dR4OO91caWyjsH09Pf7CktTq+Mipw7W
Yc18r0BnaCrfL26H5CcadgQ/IZoF/uETYYkPYm2D1AQE2fLLzCOjTUMuhplzcazyKQyS2Cs3GMYc
+vVimmfJsCPXrj0fnGxql4WJh6L6T9yIPtUVs37E9UO2x48NBJrMgJJDPaHF61/LeE0OFBUw93n9
GMykfwr+/JrEB6LwTlCvDEJT63C6DgE43cqe9QzmwN/RM0bTTPWYd4iBU3JVyqEQG0U37purSp6T
yQG0xhA5YdXrsKZiR9v5sS2s2DFYjt5F9AaD2soEwDo3R4nCMk93FkOWF1JvnydPz4zqEb5oe/3J
vchma/QoQXp+im56DAG26D7uI9WbkbKzLFrnwlIV6JPR9QQuY947ZXPwMqi4NOaaLKXeRT87xon8
3xxGClYxQy0VZ8fdI9OYZhOF/W84XPQKmXRlpwANj8dOXkah/FK9CEOKNgpBs4pvf9aCz0q/wf8M
g2ymLcEHs6BVrmwFnFZYro42e6WI11aLzGoa5Tnhiiy3bgVocitjxaWSc54rMvGrGUTpJjShumHz
gThsqBajYn3WNbnY+DAol6UyowuelajN+BBvmHccyZ36OVXLQCZxj0JHZsKYVCMmIu65gSGGza5x
ZeUQrhizA7tOAjdobGEw6HDZVx9yfHv7IeabK1HkHoy0OL2pJC+OUdg8syweimyV7clUta6jkb0E
AIrJdstUxTmLtrU47Z2Xrk0r3tfQXtULVRhDckRMHnGO168A796ngVOEluRujcc7BhtOkBmnuX+H
sJ66U9CudnkQE9Iyp9oPS5wQ/g832MzKhW616dgsk+8zeNY0doVkQcbFCskJxeEkgVYt+h+f7hWR
puayHxCPFTJFdUy0WeTn3rkx0rqpf8zjt4ge8Pvl/OlSBliYr/WZEo4A+pg3bKbN2RFvJHv1yH5A
nHzbVtsSHU0cf9K9dEp+BcL5gnchcif6YgUynQwaGbk1iX8f5q7XK9JccpuRxDjngCDIqNdbBceq
UUeFwZ0XQdoNlo4G8qOZVlZudqOC0KHUMFj1CJkLYQJSJdrdzRW12gLaQrcEKu9ACWdeyCY0JJAN
Es758baWj5nZ+f7UyMaVTLQ5Fn5JmiAK9BrOczhzjQe4alHnAEhjsnyMF5CN1TND2YnvRQY7YaM+
FRv1IVzL7DIofyNkGo/gNVEjwW/Y/wEO6nIoVPokUCm8ZAswuAnzsflaeb0ePHQOEqlqPCzIFM59
p+1PaSXl2M+tjJ3puespJiiQiPK+hJYCJ2QBNrK/UeX4zIsZOkCDv3ocrm8tXUcIXuoQh07F6aKG
v07InzjIekS3+h0s3OwCSnqbDdKQNQkAxtwYDMBKnUGU0EoUbf/ua/90RFfgmUgoXYVibWZkoaqm
MSlgSw0hQf4CSseaRjbycSFD3JTrvKLPccUFkM2AYCowARREkynSYMmyARWPRPdESX+OvgpbOr9L
aknJzMIIimFXl9Pkok9jjPVyKoF9Oa/p8eJJoqiRluPr2NgySqxixjd8N8QnxnQHhbdbdZY9LuDS
Rc3bLBBdnOrRGfs7+y3mgtQvYCV4pu27n9avBpg6KfhK6wms27febzgbm81D1qxzDPl0geCmprgI
Kcu6IuOJRUUUtT+W9z/grGC9JCmRI+ZgeeVoBpZ+8YXnO6/e1LkGcAES+pQCdcg2qumjifX14yf+
zFYauTqNSOoHbk4wcdPLGmXAL1iXQbpPixLoZONJjmKKjeh29TfEN4ou1RFkinAXDr0hKbum7TXZ
w0wJOMIOa+AmR1jkRpyzGIPnBN5Bk63162pSFZnqvAq6nNxR9aZIYm8p0Nn205eoZm0pIND0xuP1
fqQ6qzjTFDhd9GZVa1LXlVUuKoPr2zb1V7qXxZ0DQ00hnuTKZi4A++CDSXi+P8MvSGQ4GoF88HeD
hpw8XQDqbPc1/ZG5xZQeZK2/r+q9hLm8DCMPScU9ezUZnr7nOTfRVI7DE8phE9a1KnNeJGu7JgRg
pA3jtFapUANXLaYpC9/j779byWzNM5rXdFjJANYTsUUsYIRZ+/0wlYA+PJbD22U7E8puOiyZO/6u
/h8wT0e3YIOCR9sKT3qNyQAjfzkP1jTM9cf3a02IYnFq6WPQhNu4P+XEYEOTYCr8JAbxyDJUkFPr
chfMNKfj4Osf4dnuox3Qzg5pt6aSYL5yFnHi9GGiNYObd0UnYO8SL/ahqij3HEXZ+hbe33c0p2yV
cDNYInAv6dKyvfVGh4LdetH6MmLSxHmoDMM0Ix+llJ271Gj0PnikHoD7WOZEWEPiniFpZnpri9E/
Yh1Vqx2ym6CnqDAW/Lh96EwZk4+m+oEWzdStcUOT/j7RtH8mSv9xmitmIQXCyT7hodN4ai/RFSuX
L/Xh7aKXVirASgZFk3pzJyJPK292OFOnHS/Thk91xiiySJHrxSnS8D67fVpuPm78p8HuNAdCFcJb
NNem4KcvPENQ/W0J0oIfDJoqTQoSYC0MjuwplSkxD2m5M6dKA3/zPNjiIAIT4FBbuQ7NpXd7QA9a
3C5xyjXFlzKwVTaxJfPWWWxX0BwHp6xsDS/NPp22QbZ96g1h2s0PNod7k1wNa/4SI22JDBhtBqDS
Y0vKFGeMzDm5MP7/GGFgAM3L1Vmwh051f2xgfiykB76Hak2CkGv7j0t/nZO3vx+/fyyg3LKPF26z
H1oBa500QLg0FAfOsg4cvjQtMR2KZjYo/suma7mAusvpyHq1bivEQr1vH40/vx9iOQtgno56jjyt
JdB5I0WcmeDEVNEJc72bfmR5orABmrfNf1dGy/Ue3OF+jUjgKRjakhFwmvXNuNgQnIpHD21x9Yd+
EpAiMCek7QIxriDy4MCoBw1CcRlgSDEidvjP89cG0q0kdFav6kYi3RV1Vkf9O2+rNdfpj/uOQAFD
BqkjM/PjUgRdof+l4WycdtvWwrsinYqXq/o8bGb2x2lYlH7YpooTYS0mdmUYDBeZDwKA9zHfYuK0
0bPM8WPCAlRe0Nvylkv1JC9kSIgil/ZGn5cgRhKtQ8F04p7blnDyDIkVaYBUQX0iZJBsQBqkiNh8
qVW9K3MTK97EVv4ate5QrkBhwoDcaNXe0Pi+RLPGUr2GSpsBVHv9OhpyRgwxTLvhvYL5oxo0CZFQ
VsI6/lpgRTMVuceJQGh2aMcz93IUBGC2F6XCruTSy3/uRONwHzBzrISAa6iBHXsIdoKSZV+GuZrq
ALoOf3Ifsrjt/2BVzYWn/t7kP6YZFsn4X74MVpaifhwiZ/j6f6erRR6dEeovwgmaOwX0N3U8uqOE
GqYlkGr+Cs26pHhIS/zBhwvh3hlZk/dyjItf43MB1UecIDuL3XfnJWi1rMpwPBjztAhe+vItWX55
cqDBAeWavpCA7nSZdMmQnEy82ivvIGSk7g47qlUbpNw+u8tp9YPB16yMN/ag0SudfEOzkE2ewWoW
jgysxCj6+7h3TkkKbzrySHxKiQthECKiMWL8GFKdvrSscBHmGqGeWqELP72yB0XkFMUI5GB4mNXB
IJ8+pVUt5As1PEOuZ0exEvFpE2G3FIHIkiShZuToykOpo7p2MpdcFOfpCFszKFpdHO3hdkjidl9O
mKEPwpyY5qml5IDiXwblGgcAVqCH3gKfEaeEI3fKXmNqT/vrZ6RjDy/xniHxjCPl56UEx0Esl+ut
YwpitQfzgpMflE4M+pQLm79Eucsa206ccPWEIuKxCoT40WKgW/n8vCoIEt3e83IInAAPtPsjjgpf
hEscjeqfEd3kcEWtzLHy2HU2HHxlBHxRhb3KCN4tfX1EHkL4LFM/D+YFzqxbWSW9ZotgXH64Q5Kf
kEUVGMNSk49roEufEUdcH1jEm045W+ybz7/0g2RHbUsLdDgTZI5l2yUFjUyGzXRNnkH77VWU0Gkk
iUHhXkJkmzZRHcM2zHwp1eE7MfH/kSTlFnssMajbERBCshg/kpwJNdkM6q1Ybj5i6rn0XV6Zx9M4
d/sWLfdZkHHsKjBhhmp3UvuhQNc2jDw3LYFYmKfB89FZh5zRX2mETF39J4KHe6A0BcD3qTvHSlOf
OgKAF9zmuOBIYIfRQcVWC0MMhc7KhdGHRG8tEhPxdcFvyRFSCNf4bEVz/+4h8jDGQGmKZXKrCCoI
Rfn6IrUem2Daizm5uu+r1XHYX4VV2BbL05ijDd04mHueKbPMoanDXzdU3vYxPbcR4Cp0TvnSa0Fc
3WkZ9ib2aeulr9cBprREBrMDI5av3kqD8WeY9xeoOT/53zG6n/fBEgSt4OD1V+WEahjcVD56m2EM
XwZkNShT1tw9GPs2FQQ/CyD9w8mddBIFTeQ74slKNPrtw/mj32nlQcEJYGRmNS2I+RnXiKs+F1Pc
G6lkZfORIdWtBvr9Tb/0KJhvSahw/hUrsDKPthJ4XLBirIYI+VeA7/ad0JYoX2E3KWgNG/GtCAMV
+8eCkW+cY3WI5W8+2IyRIrFGOatFaeR/TGzn2PKy5v7842eZ9ztQfWnhfPlLZDA2/OKCqjnD597x
ai8h72n+0DZnr1XmfLR2Itcmwpieohv3q+Bll0sY3TrsSO5yT96wF47KTS/MUKrM+imiz64BHNoX
dhK9u3ZuKv+lKKj190YfoP12aZm3VCmyKMOiLtWg3BsFzJ/rOx+fkUDt5rGtIT/+ZGNebOOmmJzA
Pe9TKNtB5PRasQFHNxE2geSgFEkKPgaXh6Ad85TBq3fgJ/TbdNOk6qjaAspg5N+YLzZV06mshoS6
T2XMBiHch33MEMz5fUkMYqE3QQIEfxZ4OvrhiD/ZsJUOyx6x9SyYSuLRv/y8CyIfJgby/3hnQtbC
7hBNSCkU5tCYih9cKztwz6q6jickdA2BpP+/ms2hJZNcaW5KcspOKa4ePKsf+6IE7eukMdo7bzpJ
scuNoMdx8odoOmgmEISJRDIuyFPguEnALkvacAJ3nMZ1NfKIEFi+dJG3mOuOD1fYl94CaRPIJ00L
/1+ucknrN8nRucm7WMY2CvFvP8ltQ270OvZBfcOYrX7r7iC9bHtQmwz7YQE23s4tVnEtHKwWqrmj
im6uoWzuiFMkWwt6OnqS/Oi38vlwBT9mx121JQoXZF1TBAvrqlortKoqV5wFYVn9BlEr0wTSzS/+
fxYbd3XP0yd9MCAA0zYqXY/khTzNtMN9JdMk3PYkGcydGi3ow+f4v3XupPIbBAx4II3Kmkt7VCiB
QjQu+4Yzq0+BYuh3a4Ah0II5IANpgMDCtYQSmLO2P7idn8BZLE/6Tx1I8LqAwFYXzqm4qkSZDqrn
qufoxUIaObHujosdcdblkxr3c7tQ1Os6Bh6sCu4OABRR2uatMP45BAhaWpIxhkFoQlfVidBuoJ17
0fRrHbfIfiRo/BlkcRJyK+qnWDXkizVtf6GFDSV5Ut1ebDWUu3MfBExtnUHbgi964/oU3SpyMLeG
cFy4RN78lF1pUd8QEborlOQGPUAkRpTrvGJw4mYiUKAix4m8VUnLa6z+YL1rWmFkZFsRCnXTEcBw
EIslZ8rz5qT5FOmpUEkEB1zRyVSljIJYYu5+QZZdTD2X5e94JdAuPruMHcxqgxvutY2byDZAN5hQ
dTmUh0NfQH369DPWtv78CezxcTFk/XyDutvzlJSiBq0S5x4BduocbZ3JbAbiOEdh4KgM532kTeKN
deKX8FlESjvnn1oFBx58R8hr1T2wS7L7R5UAbNDTPkoCpqWMYR82ia1dOy0Nlo90EQ4rUnmF1mxS
HapINQyTSfNGJXRipETN5FfTnJYsdvO9VCtHeDdStdcFXuKFPcaURsBSxtUCSGMoFVRm+zlnHZhy
ck+Sk5V1GQLG7XRxeqCIO4e54ppdDxDykxKf1tyOkPzF0maJn99/sRnU5S1sqrJ9xFFYEB6Gzggm
7LjqlhK0+UN5reCRUVw0R9auWLQQ5WVtcfrnDdOM12KicslFC9qLws8IBnM2s31ydSPll3sJwarc
EUsolvIjwwuhEDwHNQRMzTphWElt3F0jG/uRDRWXwnGEOrwlta7q0KbL3Yz8u1wG9HUHc/hKGXRy
P5nZM2tEc79iod5CS3PfOA8uNzkLpAQJSvnXs1bCw1kp5Vb3zvpb1tipKi8mKlCf3/4YgCCjW1V8
hPxJOIiswixTTluljNGTDW0ayZdt3H/2GJFDRV0gDp3+8HMHfWpBdztd6IQhmZh7li5QmyFyn6H3
c/tmyBAsFULPBy/D9afnL6BzMYANJyUX51Qgfim+b67TQGJnUdNCq5E8WVzI3cSCVLmDHUcbo8o0
tXKf7GJ++W60EXURwE/Rd0cr050l4/+SsYinhvLAZ5HYpO8XUz3RVx3FFNS2iQbTyRuV2Glmfqdf
/bT8l6NfAhWzvIeWF1bk/A8A1d/FMrIP4Ve4/f+nO9miI+LoKsnvq+i/tmi9JdEEnkfs5eFahkCE
4etoSmW3bnPPTc6CV1D+8oFQwfwSlX0Ev05HG5MxaM2msEHCyJtkh75XQa/5pFl7UgdBarzTHCou
YpSYgAM5/Hkxe3jvo0yfWXSUHSg4aCLyMFTzMyiJyTF8xKsIgNCY+tNscWSWNtRf114rrxKw/A6r
xLyg2t0JEeVC4V4mnu1GVbU0QvpwuKWGRQuKEOgAfeSs8AGuvdALRyGIgBir+Zmpqg7uOVjLFCHI
T9euzjo7DASTm9cxHJt2VYu5eQPoMxbbc+W2jWhcvCc5tmkE2XH+LOHn436JTgAhlVbfFPwwN8zm
9gXECsZ/W2k88Di0+scXzFc09xhUW63uXSLb78edgoBeopnIWl2liN3GcdhiIITMGalswHbcEoT5
ttOYtvR60cuBzfDE2ta297B/QTlwGKJpzFaZ/PA7eytqM6AU/Oli8D+oruL5L4U3Xgzf7DsEFgqe
eIh0s7v+EbVwlxuNoXVOXmgo/rXUS5lRaXNP+2fKVOpPeXgR6GNXdo/ZYAIiCiAc4p5SuZekawm6
by7fO2+BMJ4jGlVuAdpAxMqMn7v7nswlT2y4nUsOdSgkGFd7mxu/gx77tz7Yrasem3kWIt3EI7Cr
BVW0d3NFWjYPKskVzd0GP6cm1BJHNHGc7+DknQa/Tbn6YyQj6jyeT7vmmuqf7w3tHd+szxc9l7Qn
KbzuO2g4e7Eu5PYK6l8xNqpsRCAWihqdaMuQtuaWuUZnC1n8zrh+kNNmCQ8tyPsLRVPJxzRV4zMU
AehiJAibWscvKdCrdMafmiKjxq/g6ejmuXCGjxl6pd2M9tetqaOefaGaSgJ+36Jr6pIMW9mGF0cG
5axLzGbM9/F4Xxwda7PEfmOUH120T3ZghUemDebAHy+lHOOjFDXxHKgL5cfyD+17zwYBxS6gHnQl
GZkUmjMiuQOSkWW+aH2UdTQFPVcLf9cnzmDR0SUZ5ne/7lJ3lSmUk6Y/loTEt1eGu1rMVmQGoiax
IpSBEaDsnwOt1dBNDE7NMMEpqXHUDkhtNhohI0hMtW7AVjdtDXEG0Xl8DWVhoYIkEWcyZ7pdb7ri
HJu0/lY+B/Xvoz+l4E4edadIz2LONmf6R+ASVzQwM+jhXIPsjwnPUXYJ9O439YdzqB4vfEP6Ywzz
19hN4bt3BWwtGUxbtD+Qr68DDM9DAR1wzcFolnQb7+Gk9F9nt+4V5J0hk1N8vH0Wt/ZAWqclExNS
tzZHMRsQsQqHJaVdQQjCRkiIQWmgPcXwfVApN47rKEsMo4nXJxggLqqmi2V8yZbhGcgF2VQEXzPn
iNqk/OFneRIUezq2HkQ3lamLC6Lg1uF1qquZyMWQATzqLKbBQ/EIk6MMS0biSSYNmv7JTXMLLC5X
W74Aq/ZNQ43ZfaY7g0XLi9qIE84K4eS0hIlWqMIGhbExh8/af+w3y6+2eA7mn5+L+enfC8uwZNq5
5DDBydqL3axEqYBmGj2WlKw5z44xi1U29K+MmAkuHc7yDJi7FJi4FZFdVOzv8MwWCqdG+MvJPOuv
bKxU6w8dEuLoPinBRnpnBA7Mvlha4ufCly9vDZzxl2jWDdQ6ozAqeqTSp8+WE9WiRpFw33Fn55Cw
aVuknrPpWPCBAvsTfogPdBYD8hLrOWGcaISxU3BEl7Fr/atQjwIOU1sOM22l2cx/qhh4gfvy5bJ2
McS2f/TWs++aphbbtBEsBwG2tRctHYbzsRJcH4TymiG5Loe6IbYVVnrPGvTnNp4xbfL4IdY/aDwh
Y46UCY27eIyLX0NJy/26LmQw9CWnribRrM/Ud7Ii0/L4mZE+c+sDPuJMxGH3f7BHF1kUymsM6FzD
d+NyTPRu9vKu04cjKOD/eOqlW6TAR7p39OcbiVVq5JrXG/biEfSeM4Wk7HyyNc9CHOftrTWyXNAG
pljDtGqjLRdOWrC25ab0wcSFuWfVngtlhsGy42byCPm/vduaVV7lrmjz/WkgJUMY0BBWn/nFB4jd
K7icfmD4ovSwQm+wekiKrKEwqfz8hKfnYwVrXpkclvlNxpJY7GTIjYk5l1K0Ush2VaaZN6PY38LQ
49DH+RKXgA005Vjc5FEguhjdvPYzNAHrO2Bm/Zm2ub0F6fepNjvTa2SeseqEXREXrMJVJs9C6EjU
M3hZUj+Np+w4n2ZuPvtkbwXsFALnX5Kg6F4xkFXtZFceh7TR1/T01Bi2rzPJ7AjeVJhej/GmVYLa
UD31bwAtOgWYPda6J3rsa4GZBQi8J9fiXa7OJSCKSSWeZ1ozE7UIWE5S9rbelEOtUBKgP67/eoza
S5QAcmE44gqRNJxsFBFWCwhZg9R3QXXb1D7QLO49PpQDHaWKQxddFYGJvFF4WGPfOxomuM/3osTn
WyaDQDT2j1soy0f7CF5CnxfwyGIMF7uoDsESFri/iALvyOGPRknf3I3a0ZueG4WGiutvO5KUPNtD
r6yCVLEtR2069dCj8cmFLITIXzddVaGyYT+bWtSR01P+APUzkAVb+NLCNc1bv0OLlnc3YaPSQXzv
yrkspg6W63bqDGBQ+25zYWWjPhCSiAY7LFB+kgh2DPN3zMOngqxS7cd563aIQWjwHAMwHzKhv/8h
1VZrMVelaxa31jigTqFJlRqT82lyRNLf4TC2aXI+FRMtEkHxUXhYzZzDEat376ywKh12LsAXMfL5
xeZgMkviTZ9CfTFSYcvhVLX9wKI8DzfzJtorbLLHssrqpDwfDZw5btUl7uUxe7Y2Fxwu+uavc8B0
WDa3Uzz9PFRY/4iaQrY1rwV/oRRYGmDEF2GsIb6FJLpeWGUiXPTqoEHjHNRULzZ9FFih9CEb1H0y
F5kO89dcTnkJBjGa2V2kjTpWbJ6Cl64X7yrujWwvQsGh1Faq36sqfkyeyNx7/e9eLw3ox2wp6Vh+
SnSrP6m25612JkQNOLdxo4RXVZW0SyvfH4ntf7C/4m/O38o+6pqU5rrCdYMcYrDqHwbILxnwbZqd
HWGkmtcQstLVS2JbR2hTMWM3nn1cO1yX2s9q+CIdza5EmE0kD00oUCJbNIp7ewoajrY3gK3IvNc9
h27SUOoFrqmuI4JmISYqbx4dOPTFWD/bABijTk9ApCM502ytqm7ej3l9LJJALhXWTg/T7wBjyNAY
qsL6sMZluyQkq4W5T3MLItja811Rh21v0RcSTCKTefNnt29JafP/2C6eiHjbcYErDPd7h6ZZo6nI
8S8mzLhhNU/axyAOvuzMj0EXwKsjzxbjYh6K+tedJwsJXZQyD4Wpi664oKv9F9QRVt47FXN7Dip1
6IJiwp5xFITyPZPGDQX+wlCXODzBg5sh7/lM+RG2aH4nIt+9Jbncf54QjmwqU8gKHfH6oroikeYp
gXBRgXnOW0AWl58AKOCs9cb39fCk80RmIuJ+++pxfZzzxuS6B7XquX4hJ15ZDYyyGo0sw3HBlJC0
IlDmE4SQGSeNqlREIo82Jkw6CU33voDYONVA20kJVAYzUX4NSQ9qhYjEom7Ut7WxY7rI2SBn3RTS
1lycNa1KBTbRC5CYFlhznd/pgv8MM4Cj/3cexnMMUMuFJoQXPE0I3d0wVoLDvASgIjKCuzE+9B+o
f17Iy+8+6MmC1BIXtmvEbJMR8gmZ0hCaJ5p6v3ELYVambWiIwPv4U8JyGHUS2jAj9BmqqbG6+0RE
MxKXG0IFF+J7W9EctollHAP9KaASCe7y/PkKJQCKZNkpE1drI8kx2K3y2wjyp7PyZUOWTmaLUhyt
e38UGf6Cn8QLfZAOeU54Rku0RBI72Bck2DeK9xMfENBQXVtWVh02zO9br9vaolz1D6t/N1xVI4lj
upRvW9Skai077f3WVZmaoNAfPad9VtNvqg43BOy8qZ36ZQWHmihOQo/Td9Z3uCcLSba5PNXX3xim
qlCY0MO0vs8JU2P6nnR63wfng9vwEUP/Q5TarXD78VGZ5ZkhwEpzi5JExFPbiCFLC0qCsshuCGHw
tMpDcx3Is9cVFQ6NtZ9QeIpH4JV8EZx1dB4bUBtZcbzCBXyQU8uTgN55X42RptYrNQrWr4Hmkj8v
3mk5fX5ZBPKvxiUSalwRRDPzjFDJwfXo05lhqm75/bdjM/xJY6louZ/LfIO3e0no37SKvyWYjdfo
iK8GpyYm3IfauiEP00TK04N3QdzSIYGCB7FOXDedMd14S23xqJHY13zWBCFj49NvFNrIqqqZDDir
UxeJwej+iDJFDpFWhXFBnQjpM4QqfDe3SIdWpggqsWBDX4zaM4Y57PvdqucWAJ23KYOD18yYYQ1U
tvQZs7ChTRF63FttZggKfeJSAio5WFG58UdxYQMKijGJg7bE+kUYwtrtwuxNy5j5KFQDXyUU4Z8C
yIeiA5NWLYeUTI6dec6S1v4J78RONMTfCEUdw4egIRa8aRZaU7KHNRZIlW/lHd0viyoxvkdADst6
joxvlqB9ga68U664z2xVCSX4bP04ECLC0YBNCRFN8kr9k0sujPK66tdIiSzmsrtUrTYNxsY+I175
ozFXl6la6f2Glj4Tz+PwbfBDV8ZRVIp1yUosshvkekq6wK8EcwxHDhKQHX2odmNxcFc42v9RYqO+
K6VYzAJ42WUeACy6AclGMQk7pOGlWOpy4ul9+AmziVmwLWqR9Eo4tyWjY/M4yodvMxP6QRfxqN5H
SNVdBDhd6PJn10Neyt2j0shH+fF7GYNEDx5aQEONnLq/lJVadn7mMeps7bpWNHsEXtUvp7rZgbl+
YXsTys2F93BUsVfy7OrrsFD6W29Zc1NjQNtuxEoFWSv31HxHwTTOXO0YbzNABgltjcYo0e9X9dFh
jPWXi54HRH/FozAUM0xYWS9o8o5jKM7uekD3lhbSL3+BP4ps3lXYcSuTQLbruIasC+jYrHvnx5Ye
A1fMSpBs3GKMGZr/363hT2plXFSlorjYmUVixVHpkCXMY26LylEjYEgLKOVjB9mTIcGKHpC1SsFe
Q96O1xc0gzZnXidBTsLv6Jb3B6WjMZ4FfDPy5emVe2I6dDQe7lBRGTvdk4nv5v+So87Cb0kpWa7p
iyh7wIGnEHPwA64lg52bK7A9nwV4kOqzfbg2TbLyBYp3426gAibmY33kS0wVdJ9tYDBGW4maX9KX
95f3zx2cI3NcbNw59Y0dOXsNRomgRffcL2MpGzQNnvgeVyzJg6OdNFZFsEtrQSZu6+FM6fnu+Vi/
Cm3ZvMkcaWSIxcylXDBnoftzNVi1scKdh6ApZCT5ebvycGS21XVu277uO9yLZNwaxze7ElIp1t6g
E613NvX690RgoutZV1KR+a3Mkr1MeSDOC/DXoLAqm8W2CJpBt9bTVQ1i+l3zmefaegNz3crlm7af
fgHWDZCzSGeN89NkVqD0/ococKPkSH2eLwcFj1QlCWRcHcbakTVYLGLtGnfW2AGchOb0wzLoWkHo
6D6iZ6B2AV/QlX+Wkx9cP86/EzFMOaixHFQeSQoqCYH165aID/9FZOvhOAHoL/xE/AzVQHC4xuCm
YO3RLxBAbp9rFrqECCn+NCHeJ79OrOnCBSw/v2C0IZP48ge0ikG4+vVLhOUqesDHwBCEVeZ192Hm
E++WnOY9B8aU51D/4VfHnzGKWMjgwjfHtS4LnJKxUtkSK0sEB9cw9c4nADjKFwbFXfSAxywmYBU6
jqCSDOLRCquV4lPzVen838u3bJiMCFGPF+7NJlZ6GneHGa2otiBZuDrzwkzArhuFtqai5G96OWXu
24UxiRyiVdu9qYtd1dpfKjkFa1lAIJ3bZ1lK6ddoSU86prZu5mHrS/VHvSaTbhV68oWRNu5klR0S
gAvNl+Or4AH0DkQ4oo11WS0C/gwh/7QPRKlRJ0NYg6tIYTTjPuRRN31/NDKcbOXj3z6mdeFuFzv8
4dsZFf3bNa0UkS6l3/A/URDENYlGKKUvMhixp4KmEa310nu4/Ou3LVJJoPFDISJHvmkHwBhaJK7u
1QkApkxFaH8mZPGGtOmGw/k0snmDCK045iWrpkn9yXrELar9d0DTIIG1sTMKcD+wq1zESMMx3JsW
KCv4EKeOLN1//lppYp2Zc4Leh3TJkQBFZcbwo2EKs7ThalwYHWA+FWxhsXShE7Krvg8Ko2xN0yWE
Nw75dRUSr8aoFlZVu5q/HUXAr+mCszx+wDwsmHxbIzRo/Z4Mxf9rOFYmHNZA1uuwNKLcILmkdyi5
4jK3ghgdXB957FyyKCI0ybcFL9f47rH9UBDpPpY7pQpS3i15TFyKymVTsuOY643g8gEEbqCeiord
FXllzLHy6wpPVn3t2fsX4nZwymfdx7RRooNF4agRBZ00uS0ZWxeybDcQORe/N3lQKwQ5MkLLRE1N
HaqfDVGxsuKwoPh9T7bY3XhPoDU1O21leo1ZEIQLTYzWpOizTZDkOgm32sQhMxKaAP52GeXZYjpC
xnTZoNspiv0jvY+YNns8Px3MHXxMtcr3IWWNhqgehCLWAj8o62lEphx3J211+0XVp2WL7QLh89Rq
682ZIXXCOOMZ7EWqL3MyRg3udWWbK7lV5YWvg6d1Tu2Q5TsWimRYfPEl3uu+T3PNZJXkW68ErsZ9
hAbAWO+i6k1Wp7tjZ+gDqFIUdngch1cholI9ZwJsBaAeuGqRtL2qfT9gAT7y2g8bUtiIarSpJkCg
py0csLNxrcrQAQq5m9koGfSRQdJz9mSSr3UE3DonDxmnXKCxfvXNLPBlqcR5mA5wJ/osogtzpZAw
IjHlJFcgqFjHAfe4Hi+RP4H6UcM/2zH3476ZEfg/dSTV6CJKUdiSTRa5YCOWC8tXbp9SPDkb3MEi
Q5RCZD18n/d7BsGdXr7JNtHyvolNvkbmxr3pbTpuROs418+WeR3pXJeJUkZ3zODpdfSfiqNN/l4Y
zCMA7WOzhh4r7NjNqOMvit5E4N3yIHPcxXOTD/T4aj9LYZjbwbAGweM0ZD8or6XMeIXKMK08SWPd
asw1aL6aQ2/eIQriI1GgZfXJ63d3L1OhiBXBjqg/ixlubnukAwANcr8Whlbxbg7RePLaczwOaqgK
YykFG1C2Ym73IH7AcT1qf1Fu/t9ChQW7VVUEBUfshQDPUVIqEWweL2VDmuPkoRlZAPrHTVgeyLsZ
JTN74/nIE+JvRGWyoP/7InhsovA+F+kRMjge7RjqrInK10yiqQZ82VvtdMLJ98ZUv1oS9wmPyXcl
wSNhjupedcWsWCLQv2kD6YeQsJ6I2JuHplPBZ9PvwgAZbv75f8DOSmDOoCEkfwGy/eWDJnjJkTxA
tn2lfAWyJb6sp0jEAuT4Pzh1IUx1DLWfCBxize8Yk2239eIxPRSQ1DWmT5ygdXANlUD1qFm++vrl
SWvFuuk4A+k8dwcxrlDcirY/LHh1/PIRuohX5FPVaj36/qL07lYixCTiuTTLV0wHWkMCCo/auVoL
7RC99u9pZXg4OhpPqE2PiryoNmYRm02gPcFK9o2qmQl7HRmCMDYm/bQ2FzxARsdoIatngZRkcREt
5nRVATP1Z+f5v9KfIsyOP8ToN1eCUw9iEu4Wcj+mFAkyGPXryNmLgeEMqIA9AwqFXeIqlAwXwhGQ
CiDi/35HzfxO2jLb6vtZmgo1+z64BcQ8klKQr9gXD5+iSxZGxnViKt66oPUcM3nQjPh/11Dt/nZk
+M1ahtxXrFl1+hmocM68SI9klN02jJTu8ZZ70kI7Cr1H+vraclto/VSrsPQmr7tReCgsYTWdjI0a
WucJLMTxwcTouV7gWtZZ15X96xt1z35aCumnRIGYU1OU0SKW50dPLJIHmxkQVmjti7zK4hJWc/mh
xc3iv7nJN8nf+dTLbVesrEWwBy4kK2VaAslz1NRmwVMKZRLNO+h6bSkiu3fWCerS5wvukG+qg2rR
5OKMlzdApisktDI3gHafhwYi1lEMnV7aq5H+hl09vOdROPpOqR4dY92tw6f2x7yrnZ64ac8GVFAM
g3z86L8KdyZkaethbsouXaX5ODV1sCpZsbevJxxk0v2HWEnN7Khbw3OQHmiHe0E27Nr7FrjiGHCA
QamJNCQ5ZUXNr98dCsdHdmLGuc+oJzokLePZ22lGyInu6OrRpQ+tsU6pqPqsfB6S0A3QVgZrOeeU
y7012UYX/9K3z1ImhA1vQgo5fEZmwEctMB5B7tMzouoL8FmtjLbAQflSo7sHhMyUyXeJgNVpJTmM
lD8PHYpLbrntyr24sHrljQb/lPINmx417RfjDDq+TqwF0MK529WJbfmclxdCQek598S7pkZSCG1g
csoVaG3lkZlxN5l0JNvjbNpVARRZZv5TJfo7vvewkFX4bkeVGvLIUT4cigwzEIbJkrdgbi+X95dG
M619bPwNfLXPulrjEny17o4HmFaSRevxgOlhop4eqyWn2Gcn1Qk97Q4+xlKm2gQWqaWpK6xWvUCj
6MWHVkVvx7a4FJN8uNHGGNPt7ygRE+4XzVcXfWF7Mtxj3/wObPmNYMoqD2zr+DRuZqDd1PYm9TPJ
9UJoUY5tfiZwHd2uHFRGup1n8QO2ZzOSs3tXp/9vGfEAOhJqtq/SSB+PmBEzo7pximL9K80eqc8T
RU8uY3d1Arva0dXeCB4wYAGOTRiusi6+ipQxAXMLds0Mj8LURjnqItt9eSMePgsoLgKP4BQTiv9S
T1BUFUOGDCfdKfLQSBfNo0Hu14LXYzXpiRkeFleYv9mer1LnHVYNnIfPXdq/PRLmkUjSgrvkmV0j
gcTPgI9thp+Zxgw2Wr9Zx5WA8JavNQNvFm3k0fF13J8yfMI2lxZ0+RqQ61/hYAykfxHooFG4DGAX
p8/QwpoZqxgGpAQLPfTWP1p+98MhM6IDMzbjdYmDC0t+v5xK8HftjK3n6xElksU7h0p8krRxhZrK
zbaJsyWG0xdrWVth5sEEunNq8xA6gXvlXH2/3ToP8vrK5sBaLA1froKpgUL0vMa06HQInQaqqavU
OXwHM8PyjN5bsODt11Ei3qIoIz7KWNuS25b0Intk2iQA4P7gs9fwSTXJ/+Chmcjv1Q2wBfHBl9zf
T9eGvbTcvKCjiP9ei/dGOiVcljlFFtF7kcAeXB3jbIFuOLoaMF3HfSy4RaRM2OnIxiI4xJrOSanx
4qYYUyVVt2R+MKwKxf4Lxvst+IvOa9Ji+mxBdEEYUaisBGvFAJI16A4txEH5Rfh5iN6JihyHXAPt
XgQQtckF78UXNUHYbel3jeI0O+bFefClAyymKGeDKebP+WzM4UQ4BveCXYM78b2dy/MMOgOnJLAF
iCCpqGdI2TrJZ3Po/tcA6jn3Zg1U0Lg8h/rrehEeOOGLt9E9aUmZq1h10tAuewyfbei7VhxNxuIb
54a6UpiNdkk1wsaohp7LjmjQjdNCrKf/OJoi7ePFWpW44h3NHTMC9weZnpiBtAVeozFt1SI4L4bc
eQmRgkhFRGK2q3zxWjkMNAF+puGp35W2S38qfk77uc6mfvdwl9kutEHwmUU1YKGS7DSEsiFjEfPS
fGXRI6sIryjiW0bHDuv5syYIh1Zl805iMQlP3AsSc5QAcYasFct3C3bXUzjx5Gf7ilj0Vb487q/l
1L7x5XaSx4LsWKjwf/H63ibtKAK3vMA0E1bmUencNZHR225+Rs1jcNiObh2253kF65h5tzvjDMJr
69rFDqP0f4/4NCbxcf7ReAwo/jHwF7Non6Lq+dKc1Jr/hCTAu9GGSf+E6PfOfRNGcWCvcrm64xzb
9N2rPXh6sQgK5dJ7O9zNAs1t0+hHUHu+nkjVfTY0ViDrwv1JO896mIi7ZtNE36quJAZ81ELG+FuM
lBrR4oMgWBq3MXXnql0v9DZt/TaPoJpQoz/djw7p6HJwUV1GClbyAaMepZ4o8M4r6+dQsusFUDfW
Y70V/gDdDgW0XITk1+VXTfXY1kLHMLgYf0/WKdx+AWNneYcVjCSHpx7C0KoK5Ai+fcjiYIoTa6qr
iZZOp1XhPaQvGpaEnc8+/UjeZXBjYQKUJxBpkYX4yeu+QsN++MZjSFMYqrXYcrUGNqqybEIp7xBF
ZQbfZr4JfzCVFXC67xzjq5n6ZVU34daz3Ejzu5XJ/JP++a6fyO6883mJmtUP3bxOBXvOAwMLJy1N
ig1oDS3jHa/7fkci4NHP7/BmzCH89ziuxRr7tcYwcg/rgls8KJZ9attV8WRjxeKuu7xt0Eg8Glj8
HcBDAaQ++auuDhRnEizwyQ8X/UJXUhv08Qa3SzrHH2RylGpzXCWZ8+QZx7v/oUEZc4kJpWPA4YHL
j0ZVjVmBX1EnkzCbfdPUUStXHabIqFELrndP0TXeYkYBn/ytpiMuYV7KGAezjAcNoYEPbC749ssb
0f5Aj9ePTAKMajzOr6gAjpy6VvWzcoZShFNFvRky9YUS44/AtSAtjPt76e26HF7oAEq8HZZCGZwp
lygInuRgUtO+pPsCkwk25I2BufHZtP8gnEgE5K9FTyyKLQFpW8EqF5EIwDk5VpktfOzHC74bGDHU
+ZK9Ht4nGoLeqY5891vJsNAtP8sHqvTU1kDyhCRtoXuMy2WD+SAgjRiDOle8yfEPBIm7k+f1aXtp
SGnjdA6M+wo7F1HLZxPNQXYZ1QKe/WUwfahaTeCZ7Gi9Q3U4/N2ZmAlouSeziu3VqYVQ7+qbo/8z
+9cYoM279apFV1PyZMu27Fs5aHmELc+sJtf1Cr+42lmafqWXCrj+xWS5rPZG0U5RBhOtxa1WpKq1
KyLyvq933vT0+z+NwnPuBEGoFtdAw63U4mA3xYyvizl2S0JoOGPIsTah/JxIqXnv31HISZPftcdR
thvwXNxjGYt22oj1Rs5H1lBtU9MBj05ncaGiy4dfcEGaZVuHrlBDdBRdvdNQz7BKkODrWNZWgLQx
R8SnHaAkwmbag4imL67DiU+EkPOnrYeZcLAWgVa6a3QO01JgLc4/ZXrmXZLA+Zqux6P0SYojQBRx
mQz8+D0U4kRlftue+J/fXLwQm3DiOCVm5rbNZUdjKXC8lHAL+z1DLVVoEyGP0ux64RDoPvlx4waC
Q1tj1bBiBRlBhDZhlf7xYfihBTEeH+m0a0N0p3xU8AzSmaVqYjdeY/03dyNZ7lc2oLWxhAuaVvEF
Ia1DP1u2TP48OpLrpbDMnVftbY4tzm4XiRfiGnsa7cFS86HtXGSNjZlwmnXSR2ohe4bjO53SLgYT
SzZKQNu9gBQXnBFl2M09r+kCQG8f+PkOLUcAXe1TXqejmy16jEknHoB5/vPHdfC7cpwK5yaVV5Nt
z8FoEB4ss5LR8Px9cqdsqOZBRX7NrvH0jau1oi5wSDSluJ2SuggcEwniNLg1rqKQr9xEhxe07Z+U
3CySQBCtzKaU6UH7cBquz+yug1DcWN54LrOgir7mBfg3wb1tTqdBKHJXMivCfskngDuBO2p438+J
N6ZtSUNrDkMl/3UMZuyWhdnsXRyLw1ICaIFhFphs7YEZEgH2xVi7WgHzB6COYHRrd35YdTOlhjEW
f/rBwQ61mXTe86IsCfo1f4UUlY0aLHrtL9mGhIfEuFBuWoquMm2Gaf351Gaoh95mMw7QXgYUnbWt
mN9tYcM/Q1VtEc5CtmGoWTWzEivmObab5URV6r9Y1VUon1UwvzxnAT5IoFZ/DMr7oB8Td05IT4+O
y7k/ryQLt03KvavRkAR4wUsV8YK0I6zIQQslmwj7FGuym5ZD46ocqrQgpni/FPo2NngaowRMNrSp
SIXV5BnBduTGmT4lPfTfncATFfhis0hI4pRTmxd1qRnfL6r08NHTuoA3zvn7tb7dJtr63VxKhwba
aV8XhPZwUih3nyic5uFQJbmv4zLPbdQzBIy9xW1ugIONQYuaseZqSlQM3c+BF8ZUKQHndMwcAmE3
ohiuWcyzb/v6PBZhWnoBWSuqQ1f3f4MZonlYMawW6Uj3hH6aQtLwRo3l8nZ42m8Sv6GRbg/+DrrI
ijfRNY5QqGzdzwS4R478rRJtBBf3pRdrQg80z6kM+nl4itmOV8u673yyiSXfEJt/SIhUr0EN8VbG
siApBsMKHi2YW5qWpdqb6jugdhM0e39W/LRF3dXWsRhfa5zVhFNaKibiBPWUd0/ScTpDaza0+E/p
qpsMjajAJVUpfquEcYfga9GNn+HIav6xybsTKRlRP313eu2tLck4QdFAYYdXARxpHJnLXIJJx5No
tpkXPIMDuWerzUXm6i2gSm5hgEOemE55jZW+LnSGnbU+2uFcKE6Hu2853xBhVWlgxRjlqkryWTIh
QYrrFyDI99s/6duHv38YvHtvvKDrxj4PDConJrN0MZq6UQasBDxsSQK7fnDLQijvZiBfivyMMTks
QCmq8dZsOLKqGCCt/dSN1iAchQQ7AS+khOygXSiks9jLwCKrQcGz0bAIGUDbTj/9zn5/KjoqNPnT
ItsNoUKtjdqT29tU1hOznlqaLtJL3cSiEoAhNZVoDG+3Yz3zlO/L4VdOg+2Cf5fa6w4unAa4YqQq
cbBDPZyVqShr+jkmS7CQ0KHY+R1bo+Uzca2fLK8srzhNzoyCpo5GTIJox3QsDKKjfBmODkj3zBkW
s0Qf73V0QGhrhgZAx20sM2Is+b/nnRWcxD4dHd9f5/7MmLWJ2iHqP5faGNeCbzAY8lbZVXM8CqDl
IpKkxQtbVFDH02+QXREEZtdmukBGyUvqh4BEKFaq6uytgj/cSdRXQMDZ7/G2xUhohvTndGGz2BfE
ghQsx1j8UoowVzLdGwgtAFYQULerUykTsSWdfuHcTT8em9cTX4qvJ+64rMX+mbynwGSSEfXO4Fhs
KWy/zPn4+Ud049O35PHWgBVP28vIbpX1dW/gwBLl8xYEehdhR070G9ZJDhLwoMP5mY4xVZtvN79g
HqsbuCTBnObJI9ijMRefI+PIf+sYZZ7OfxNi4RX3F24Dersr1Sj0JEboBBbiDvI/VKSW0yI7VMpa
VfcJXP3w0t4Sm0OluBQaQkyftnI9vmtk2g1BYrlhWONbgBnQozy/+W0WHPlN3affnRue5bxl6zIJ
9lO/ksah/r05SN51TuwTten3CXiiE0Uu3xcN/nQ8itiR2HXEUFy3bzMXs5YWqGeeAcAhrA761sGf
Cpa2P6JkQq0Wi++aK3SgNRCF/thNmfd+5ghUYWlPecJOjdrATEKslyxs2p/o3a1rZnF4HjAOGuo1
w1pATRKouQMTUdEs7ZskOQIs11JvYfVFp9owUzEBE0bG/I2ETKhQp8hP/Mae+bdR4UJsZjmXPHU5
dQq6DEDq5YIMj1Od0IGqo8Bv9NthSHoR0yrl5/laFJxyyGE+3UhgKOsD3DzBrfr0bQFI0xM75CUy
YvXaUiFQzO+jT8x4s86eUticjD3VorEUAp/XxZdg55+NhxTbegGxBvE0R3ufZWJdoII4JIeJfRVx
+rzmIvnih9g01ySHpUUil8igdMrLCxoLyx51npw5OvxpKi1J+k5XoVkdOhwX0965nvjZwcoGS9jc
yH87LAhJ3YJh7kcmS6PWo9GkLHBoedI08HQ1zuSOI4m2PYjfJFG4OXkC8KqIovRNQdp2PxBDBZxj
/z3q2104ax6u6etSZe88DcvFvibMlJeSnKeMTrLvrPxrBnZwIoirC6qxnTWgPCS5ShCN+JmhaVTA
fabFy5TPcBRd3cZREAKDi9e50Cjy3ih48yweYdCwFhxGAz08IUEE5K5mQCAgk3qA0+Xrpw+2uMpE
HjwTEC4CJCNJ/BEc3alpcRoUyGaoIvLbkyRa8azkJh8viGz+9rUyeUxX+6g+ex6ZVV3ErKYJeHJG
klvl12kLaWk6jdpHL8MYWNlHuB/kmXRY4C/PP0ia26peJkw3FaNQxuP0lqk3swdo7qM9vCcGAjog
vLCy29hBwPXwokPSbdyzy4fuAJYMGR62kh3U759vD9I9qOcorbV2wCNPG2un5wo5XJ6xMW4lwumV
Gcv5+1xu7BaKyCYy8Tc7fhzZqfCEnAN+gggSPsO/y87FLFkEfdBIM5v726RkAJAAKqLsWNr6b5fW
nyrrAfOOm5qq3rNQqngbVHxPHl7f1R2avBz6Qwmxx0zX4Hvbs4/8RpUjZVck0s3xNaJMHz6xerKQ
32P/gL3RaKb/e0Szi46EYG2rH2BytD40Bc1g1eNPIUFoqzNwlFq21XeMDPcdmwRS3GZaT44UbBDF
/1nvhLEgVKcXMSPxLuw4onvVjRElI5dajJLAzHiXgyhD5dCMIOsylKutP44aXV4kOvNzcnrtBktr
FWCn961bt7KVijJZhmAh1MseFROeN6d1+fLSf0cbqndKv/E704PasNofj23UUl0Qxu1Ev+YjlfDg
Q3qZ+Mwc03aoZabiVZe0u3cI0GYuaINPwc2HOLUXKzN2MEaedbY/dKFHnyMuHgUC4ftXKbzplpEX
QutUQG8tK6yMu9LQeGDp1tOJZrhX4AcZA97AR2HFAAtkNTyVs2GdpsjgiKCHyrBXbscxkU1IhJWK
S1flDvm+3mgDGngHUJXrIs7kiCd3mt9Qoz2fVhyChl/4tMSruijjknFQDvLBA7DZLrWNFFCOV+Q/
xqaAhIFn4ZLhQqC/ycmNxt9MQmeygtezg32QKN1DneAGdpcbd4EH1IAWNnZz4kNadclu1PtchX6D
JuljjCfmNqbPadNUwwbZkh0ooE7elr1h5lVwMXbJ0Ir2wTSyHbJkkdvRBtZz1VCyRFXKdQVpeyyq
LROuoOjd5+wQWf2Tq+jVZnJxByFk/jPSZR3c4gFsIoP8LF2gO4gWjpqWDtLoCrOVJE44zcOGhVSb
yqNC2eKvxVU+PFrVXyR6l8JfWx/TVt7DL2eqh2aJDGbl9xUwcN77YxDmZ2UrPWNt43Qyelzexu4z
QAK60+P470p5tKqofMGZzbzF7iz8Oqy9A6St2Z8jTrEOIIaE3X7KSiAcIuLNNF661fpilgRzBpBM
Z5Z5lRUCPWBbP5IIyQGP+yiKHGsBRrDJoGKzBkoHQ6OpFxu8L2VMxzFZQGYS/Q1LVbEnPRYn2QZU
P5gggKGg1i+uaUsHTLTrn5cluEupklG+O0vviwfZM+m8VDt2YRzwbptRCyfgy+2FoZNtO0isNi/2
f+dSBdg6LKBIAxGvFmVpms7HJ1XXZjj5HJux8r+OA96T3PdH6f0hKGYmS7yudCOR6HOsNCNucRFc
LMMz3QuiqjLLA2NCLk+ldFtVwk8UdTVPHGh9Mvmw2yyOaUVzWUDj4sQG4AKtuTH+dSOpn+QXCWB2
oFrMIhn4f2E0+kH2xDFVwrcRwurWH1xxL5onJIqi0PWB7AcqsZ3lkmGYGAUEi8zeohmI2S1vpQDG
eV90p6lIsbFiRwrfxx905H6iHFz4qHj0d7xqyw7HS4WuAHg02aqGyv5TrrVwXo7Scl5hCn/2LgV6
aGibJhCw5ayHnVIeG3mkPf8jCNpktjysG+cRcolauSS3BdY+xa5Y5aVzYXvI1c6mQDPPTW5baFy9
F8z2Ty3MJpST4PPVyqOoM63AAlwqk8qi5NWGIBtCjliHAmfCoCSyZ6n9DGQfioAxbXip+nuiRmxB
anQaesjO3ENjGPIiH2Y49uThBan6Uy2DlupY0tZZbACMUgp69F97Saz8fMd8zoL12DuF6O2JxM3v
GvQ6/zgvvO5chhkug9JDFZZCQlaapW63FovqCaslSA1Je3OBRg1rl/1nSvOX69DbcHkGrA1fl2Cn
7IxcLG959P3rc7/VXG7On5z80XeRxf6tMgKZ6/IKFIUTTnY43e66z50j+Vm/OcGuZMNP5v8t9iM9
AxmwYMvywZncsdS+G9QVOW325JMouVAd22zQh2mKxvyT34uXpQ4Y8m99OBCdwctxg8sgDMRaB9eE
vc5PghInaraJILKQbSXHqj0c1gU2lj9pFT1ntsB/jn2047aXnqXlRtGxEGcRqZr11zvjDcJ5e8rZ
lowBcXu0ISwFUfm6F7PB3To93HZzygF1hbh5DakNU6eg6sT2ul6RGDficpOzDLNY9Yk0oWxrE5WI
uou/1NBeFUzhSH1JLFQSNpM1vNteoNy32hctfl84h+ykX7gQgN5iaFQdqZ1ie9KayQCWTva8mB4H
qPmpp7lFEznksk6L6PlpI3J0VLnqzwuZ0rO5dSEgSR50hvhQjnZn83xD6xU/xgSiaJg552zZefbQ
/hz8jKMVO2w7lwJeCFcoEMo8URO7aU0boqEqSltk5lB9FDm0bzbT8BRZ+oxSLN93jCkalf8c1TR+
OwczwCaATHbxuQ6Q71zqFE1kIemUy216t4EU2YjPRREiA7Qqs9nQgJvYBQpY6bfOedYWlar/ITe3
5MBx9j7iNkoFYwGBijPLzpTyr409aJJxi0+QW+STMoS5xBNKuERJLpzkUyU7P8jJPpXRS6zegYDg
rkMEPC8X7cwcs2PLkzKtPG9yYBd80WWKfa0jtywlztnWhktjo2fSJ7mrxXwSypKLtUtSb+DNlA2P
gG+91eeb4VJzOAdjDGjRlyoj6EKz9nFoc23s1Iednr0XIr5anIBZLnPQLv7KOY0vhOFRTFd7cjGN
wBUGwWzwSjDmyg6w4O4/HwlM6KiMKugNa5993zhj8sNZF60Cc5h+sK38N7zm8/+NZJ4CLF/NEJ7n
KKJZanTemGPnWdr+fQgBKGKDzaJnMwQR0DNNlAelwPELTx1LOWCpH54w4yDWDSjvT/I3sRoknxXr
cF+3ULK080jzEvXKMNPxVoQlX1Sp5x1piAMgqI/XBJgT8dPpAtBLgqn8K/PTCSAAIPlQjBY2Qasp
rBHYaz+mMQ4YJ6uxUXYceCtRpSfSXe3IH6pk1RKERF9lLd4F3IH1IQl3mOSyP6vdgzkPBlp9CIdp
ZiP4DbrGlVi1SCVWybeT6aBCp4pvKTWgD1OzKAov3oH0HWSQ63Td4koOc9ngvPVCisFRPiJZZ4p8
jmM4QVSXXeGnIn2ktf28rySe+16R+CWlE4wxEYYGzFYgIQ9PnFUGVB4IwvywFfJpMKfm4pK2Ow8n
3CxckyRCJX2N1SYg2d/mp7soZ25KE26RI4uRnfEBKGUJwiG6LZBxJB76QqNh2jhYq/xTRQ9X0o69
PA8gGjycvWTaujd3ajZPb40VjNFpoby84gWRuIVI3cpD7P0/ZxIIca7F79GnaHhHP3LjJZ6Ay/dF
37Fl1NEuRMTYSTIUPNpYsKGRqe5wR/jpufQL/UVPgAgyozoYYBCnpxLe+9uZGSqUxIrfgQg7kE54
jWThWP8mzPn9c3PDz4Y3O0A6Bjb8/ayYZYq1gcsDEF+BjLiK6QMuOnDJ+gYafR2ck2UsBCWglikz
j2a6QOkH5kViD+inzvzzwb8ZRQWddDthPDGkwOON1QV3lAwyKGCf/baldM1vMmdnojhLXH+3wpTy
dM58vJRKb/1jtz6umkVeWD5lsUNAoozRGCNSWUVUb/xRWb05FmXAM0l7MSohcxuWEX9PPEEV/LyT
eShyvzzyAKDVTwI+ZbukH+Bmta3P6ck5WiRrdXCnv7IhoS3Prb05eGTXY7pvnbDLF7L2ztNDRc4O
hpyX4VmroKs6pu7GXbcOJAUpKYawrsjEHaY+XS40LZ0hph02FVHyLjgNSxlH9UC09Ufnh8H72nhG
2lR4NEudll6o//kVd/C//IH3iWlBKTMbUknhMx526ziMocFlalXmHUcaEHPyTwaRO+OZmaVVsdsW
WQu6uhKiPgulQJYcFxBD4XF9z4pYER+AFg5sJO1oI3qZkd1tzMPQ57aHKEyqdzAIROyTOhj6JRAH
bK6vg+dk/lBqO0ztJG07p8MFYdYgsfqPsp2h/GlbcfpEa395s8XluldgXQsmabO01zVGSQZjEgFM
PVw4eU6WgSb0mwzqjASy5ilXYdNmMEubJoTYLs6PkT9ZmvQkiaPwaATyc7jbzNFhXRPgy94gEO6U
JaoWiRvivF5OJKRWHKXQzxFWeXM2zfr90irrtLBAr91/2qJlHP0N2+8iscCAzsnNc06pMuLiJptV
xxUsYNTCShVt2cO4t+P49f7Ee3/gihwGvgJDWmnCESo9A03jh6AjYFrQ1TXLbGzeqzs5D0jWsSov
0mQrkpoIbcJS72lk0Z1z+2wDIZC3MG/kyLnPr/GnVTgjaWkwN0m8EIEuL4dtegiTURfT6PX2Fz74
enmPO3nmn+zci8neMytN4fZCADL9FDYrfRRU4aLy6rcVdy/b6X0ZZXcRSdvyYLmtYQifUnrjq9tZ
T/tX3GU4CBRnaopJXKto0XUwqxTGYJ9T1WaXP7IbXTbCXvxNyfMjTIgIIBxh6kagaznbyQRw7JBS
HUSlIBjm8IMG3cR7EeStaW/BV52AYX+QUWhPqE/j6zdOls27Z1dUGS9NTxZmCbX8iXRj7RbchkoU
WjQoK7f7FE5PaL9rVYxhn/IstWS3ajtI+xU6NNJ+WMn8hlfPoYbhOwthvJuzRh+lxw9O1DWn5M3n
uj5wJJ0yxVeHCCTl3avwznK9+G5N/CLJMxXYFO16pP5ZYv6GY0OkqVwL58VJGZ+bK1MgxcyIvuxI
Gug+LWYIWUHARPRZ/59WCz17yX4eYHPBcdo13JReJYlSYLDnH8rTwF5TFL38uQWugHg/Zpb5cjuH
1JbVgVGiPXLtg250N0+XR92FAiL9AOaISGzYe+Nkdn2CI0bd0FdOFx5xsvA9rr8j+Su/W4/XLBc3
7ueWEmzekctOuOIUo57ZrHw2bPIaJKbUQAwJmcReoETHwEqc9etSBPau5j9tYPZllgebmmeqaCSH
cvLFHjux8vBUO5T32rjxQAK3P+mCI2L7zoW79WHiCrMnUXKlsoZ25lQwwWa1qKI221+gh/oYOm66
H5dqlRQ5BhshIEkRn2hUwEB3tzOkF0tPBJhKNfuWhC8E0JVnsBSwdnmXeJ9GwlQJXRi8gV80kWgE
cVdKEo+IaOngPagXoqRZk7uVbQcvq7wIctQJNQb520I6FhDtAsoi/bwPrN2fAJHZO7MFkikFXJrP
Ywh8xZ2jRzPQ9oPBJjV4ugN1TeyF5uWiv+d0rtnCrowQYHXYzFExwFLNMdwk+EC/sRpy6gL8jDh2
KDzFoSxRsy8nxFeTDvL42HQ1icDRuqi6UYMVssGcXJSkLyD/ZIwd7ymIfXvDBLvuXCRnvhYJWA3B
GhobK8brEt2TLB+uCy24Jmkw1/0wMbjogHPYMh+gn0pRuUHOWVpCWFZjJVMQiaB3SBddcm60cMwo
o1YR5lof+3sfqt2RvvPlLEn39tYpQthUFpS7cbhAz5FUSqJ6x1aRFwNdGC6c8GlUBerUtGkBnJbE
xI9ymS0i4ND7AWvljJS6a3me3fff33AImGf76WzRgl5rGAVEkpYLGt9KAH74Lu1hiY5843Ls6kkm
BtjCj77bDneIuDkVMMWw5OYQ6lHkjO5E7rRbTrF4mG9mWXsfZYlp4Pe4w8YQKOWrNmUDmfBJfrwe
vzeO+AT4AguuEc8t26PZp4hZuqIU3Fto+JpbzCzn1IMvdnbeDb01KKVNj7FWBeU/ez4Tp90hwWCG
BXC4o9yZEQz9YQOP23LWD4fOFsYpI2AlV3n1albo6WWjjKqUo4SGiiUDK+dmUUVy6k+wVAd9batP
5KSzcl9fAEO+BG5t34FeGNDOdu/x6XG5gBJ+Be6qrzOn7OB0ug68Evt/zqPYdVtTkAs5OhOuArvC
KImr9AM03cMRLG8W6Wyvhk5tIoqSlDeQ39shcq8XtuBXnSm2Nu8W9O2trzNTeeFLiDAoaXFOO0wD
tnCmyGYrsC/dpmDlNLSAh9Q2lI0ozmzUxfXjhigJa/YnYy09/+e0v6uJFlRzGofvoSbzsONaOzpG
xXes0dgd2Jym2aJmlEhuRXYYSXzooFPn2Hb6wXMfChqTu5QKm2WF0nI+xjLQO8Z2XLODc8Qbb5Zg
kbLrwDqvja8Pgiinhz0kGos42VTmQjlvhEbLIdKSObuUjGNJpqVcOeoh4vbIZpjGbrytEF04uHEJ
3XdXfpmAdh0zr5LJsystojlcABOShopPUTZBJxRNf1BXATGIjL5Qa11TtEobic9193IjBERAaicc
TEtBMT9FqVnk+X3ZAJcKowCzxlgZvp3IlpDgDXOjTk7pxPSwfLBtb0e0UlW2ObO+gFzsBLFRVGfk
J1ollxizoC9tK9l0JPJCPudDVLLert1nbXOMp1Vvu1uMWn+7U+a/M5Kn+6OuEbkDFUpt+BXAbF6z
3vUAVgwI/PpTmRUCSznRFUBK2Ps4XFeCcmEwAEkiI1+sr0Wmmx2aOZ38QsvYZk8fZRBOAX+Aodta
ixgwS/UKoD658yVe7vpyHowprSFx0qkfkTnukBxW24cOO34tu3oPjz3xBmPCLYJsrbc2a44xa8Hm
Hev6EBdVsgejthhzdNKh+CkHDqc9JnYnREf2awm5oV8Ta/tVH+ocUHv29YxOBSltSbzfbne0pV1f
/btsp6YDyOfGgTeJrSZbRVHdpsxRRpUzlGaMWE54+jGP8oANYMAPlA0W2fY+19u2WQAsNoLBRnuz
iQGaRIE6zdKoSeA0Pz9WJAj10Q1hkVVi5cCF1BLQ3bFzc/MketnYqfu8lq20ysiDmrCezkNp2ZOG
ykm250CzAdrnqLngqI8yV8+xhcKx379Q/dmAbYugk92mJnIwehC+wRKkybCc4KEaz+OrJXO0EaSE
cAnKP93gAJm18MoJt7fGAfnSb2XEhfCTf8nLXt5mlvnG4XX1aFE/MR6kcjgv0fwcZkAu8B5s5Ufe
25halToKgVMAM46HJo/YXa6Brm+t+5Ohrwe8pqQoKcc4TluAaerXIXIlEvBHKdHbnj6tkTbL52Ob
37OGL1+kBwaF1oMumdXChazirQ3uNe4AAbyGQIyMMqbVU0DAYrwSiMLV4saeDTqFCYG0EHryFFVF
qbgF6HBLfujM6q9jmTup+4BqpyvBCGBlZfQ6G4JAPNuxA3nB4F5IdIRq58GJ+3pIL4ZIVIvGAX/E
ynUmLWiCyDmaqHTKeYkRfcw6yA6v5BOTZVbj34Av7WfiZfmZvrtHLTYISZuI2DLGWOqXlkKWpdcy
ttfXY9yn/YpgPB7tMUdhB74r0dLCcbymnQTRU1Jk89QJOfIvI253TCeH5CIb4tBhKXU73D8lT5vN
8jQiKSIZoUPMDz9FxmM5n4kf34p9hL8QnMVMDjCk4Cnzw/w4eORWzGFbKzqdnugn9M4xAX7usyTG
EHnccfPJ5C1R7lsrKnvU7TAZVNIjR81Pmz0FRPSutSH60EKrZWmrtT11CuV+K0xR5+HalRXb9+Uf
Ew+Q/LxSlCK+S0NV6mCKZh18OXRRPHwcGOxUURLe1BN8sPOx8oYNwqFAVlJb9GNmDeznmg5Z6E3C
gJgiMzPnXHu3HCNn2nSoaUsYbYfz5oh8hhemGgiYk9aTZYK4juQrS8+X/sUvV281i0lDvczljcBN
xx3TYT849u3/qzeoWFIqGOsPhKJsITeKW1pp+fZYIei5VYKZXP96wES2bzA2+Anv/AQP/Su/IiSv
E7pH2ZHaxPpV1gulttyQE+qFUo25JtEGShmCl4r+Nfn36rmyQvwy0GL0aA7byYpW8ledz2Ufwdjx
zB6giRCWFUvowLbTp2IWhdKfxoAbcSavAjuLhuZmifsy0zIt/6RiVgN3560SO24SnrcqzUAoJa0A
HmWCNfJMDPey8RyjUInFhhBi7/qxEhn2X0bTW9N8TiKMOcVFBFXfHPEywNNFsiS13GZ4MP5rRTBc
uEPsfEzT+YijpIjufGLEv6GBTCbZ2i3COLCn8DM7VN0kS3hLgYJFUkJe12GgrqKzcMWiN+9lAy6k
EjImuFziBMnsRn5uGkHMGy1qSciJfP5vnYizGrDpPIYqrd4/SKTXNW8GNa8rFBmNVa0MzYrC81lM
hFogRTrA+5QFc/sF/HOq2Z0pmLtGYR7n7sgA7OBokuyrYWVJIzsTkD1HPwtnWF3dmS2NrSqpmy/b
sPyofslMOLrUinte9ELehQzFRuLmNKv/sFuA1QXx4ffcRDMxQEy1E6z0V58sUXeR2/FFnLGarQn6
m/i0/WH3WdQS6aaaZDV6JWjVw548evLx2sSMCdAc4YK1LhH0WboRi3ddEdgCj6j2mCUHwh7UF8Hi
leKTww5DmJRo4Dxjo6stj51dsvw8nWHgNW78bEp16yd9MnTyaQkhM+7kUZuazOz7B2VMcye8uqa0
uv8tflHkNUidLmANee18BAvjW2xuqBR/JkgpnxR2Vt9nhknztWYrDHtaZAIYn1knI/v6thohZDVi
u/gQHRQltwh5krOR+RNnDXQ6Q1wpWOrFib0PiKSj4plTZdSg8WlbK19gZS2bTtdqHPLfsaNL8oRI
N8mR3jOVYYrLz/Gi9Z4O2wr/VQcrdJ4++jlxxV2NI5o6Yw6EP+faP43OEPmuim49NBCVgURfXZj9
Rb4c7hUUVyTY2zkx8FsjO4TzlP1vb4mjBssF6vDWxzi01uzynOTAQsdmrABC/oizin2UJ/aCumTY
fEvEf9W7t2qaeykJb37KAJIwD9rW/NlRbI2S/+f93rU2PiOZJr7CyWo0s9tNVJBIYZzOvrsrkezy
2e36a2Rpfc9bjZkDd6yCoAUGPW9YCmesMcDjMOY4ZSXB5EOmoO38opxuTcNymvsf+OnLl9+q3A+o
cRHoqmm8n085Jzm2Q/Etod7QlgXxPhUC83W2sz3fZfv3FgeN7bVtBUfWnBoe7rq0NY3mMfqbVoz6
RMuTrGM/2lQZR0ZlMEteijTN7LyN9ukG6SUruwwVZ+zA2BZss1joGB9Tk9Smhnq8HLYyMJ5wbea/
Eo5TpfWbKX3HootQhFbzNYhEI6GZWmBNIEHFBuE6B8BcybAMhfIDlAEotfPfGzopPj2y1FTDF2bc
pw/t0k8VwICu1TclpvNi5NdgFjHMe4J3k3t7SxuoamdhA7YbUoVXN0DPqn6B7+EAZyZwRtWbqlg7
y2pB70Z06un+L9m/qQA5e42wXRnuhehjX7fddQeZD/AovZ+teSx0m8mCN1ZSwF3qu8QkaYXpugoZ
v7BcMlpfgmCfIJBCT0qeLSCKIZnNGEquDPYJ8T5f1YkmMakLZgJIOz2NDSVnKc3Qj/MAtjWSQ9QG
90SYw7qtcRw+kPdtj7hozB3fqxnlYmosEGeRssBTMPu6WRalGv89PZMrJ38B41fk4hQPj4MHOkfF
H5G6t+HqI5HG56MU6x0YwQVfQvpStlF5E1RKu/5THp/KTZhl3NvvrBGyV/mvfFj2EV12vnkVjMN+
d/oucm6qW5NTnCCLCbk3pZyUb9nYGE5QpVQpwoXQvyF1HVuNiFQ1Ng0+k2xWE8W8Pj/8GRTHtoci
/HqbZ8Zsu/H21YmnwQwN2SfoU7QcDm1AKIZLch5OuyHxPpAKiTu09xUqepWtlNbKUANsADEDbi1y
WzT2VCnowKDPhmuseCV6G2B49TJ83jlvBpn71j3+biw209y4byGjmqkQHrw2DUazmBOWndFlFWjJ
rRxn1Fn5xwz+fMrt4Sc20audAHZXu7xNgkhiabfD/wd0LXVPfPM6vzhVdb1hkP+9Wvz1UP6DtpG3
f8k3rsuUYfBBN+Oka6zfjL1wmd4Oyo2Ma1q4lWV8An/FmZuOo3bk4cVOsYMSRYHYfhClNYexVvJ4
iIF0cURePuvniQRLR44v+LoSlsmw2HdCS7IdJFaN+YuuXm1B7yXk2l7ozYPrfdXDMX8WtDAHNvBU
3hipB+p3yBXVPnqLyTSGUDf4cy1/lmvsTCquNEfW5iCPSNKOzVk/EW1NKCFQ+FBiA9Pz1Id3VUTe
eZQNWrCMYFS9/G2LntJ0DcnLi212ZiZzs1lG1hJHV6JcX+YYBmstatA+5kpmGBijI+XVjgRgSfIw
3pfMb+nSkHIoZiCyEHbvEIKlajZ5Hzmqh+ohzpVzWegEYIXMvcpSTA0sdsr4lDEHGGQKtwpnzo7l
CR7qgVC43mjB86BqpKOl3NqEV+guZG9JoaGQfgz8nIRS4s3op/ZWrGAVgs2cNgXpmwvV8uuxswQz
uy6LvfS8emZqTgpgQn46FIm6fHYII5jSILNRCH7GokioV9TAZQey4n6tKib3pj4YycSaMFGmwJQw
KBZpygxvHtIqcgXOmiKvFc2dKPhsMcNmPL/+SIdJBuYRcGQLFooUnDRweSaWUSXSzdYrO/OwF+m2
d+4h9mm8Nk+1Gyr5KxyMGV85sWsh8wkDqtfQJgu33aESAqppFKT81LTKjR/92U0TW8yWGAhgZF2o
yycrepMm0NiHSyAVbgb41CM95F6MJIGHsNQvoPnYsI+Zr6pbNBpFWJVSK8Gx3dtJN03lHU2lHdfD
wTFoE3q6A16wHjNLEmpCPidznh9tgAanvSpUe69o89Jy+bvSWo+KiPxbgwVqQNwrfccXOphvGjJ4
VmT7ZAw9g4F11AZgRfdpj55aIBTSJkyObNjDCRG6l03KeYNVBvlajFNvwy2gUn1a1hPwoi8jIzCn
ZfaN8iwe0ObU0tdQ1pMtidCigLHvpzf6CB2azG3AsDtgmBezrC4IAvmcdLriU9ynA1ddz2zuW2cb
/8/xneIFU6x87gN6EZZFLaoHmBUMzkqZFzEmUTEcR2UmfIRtsIbaQX1xTvNFKjn77w1v8MucO796
WtevOmmVEU2KdkK1afG1NAtplzyvEeR0D+wj4dg/yksYd06oDftFVa9tMKEXddOFnbj/gYY0XNlT
oofSqn9oOhfDghmLO7DWxn6qqEwjSy1FERrNUYBLde6JWRBSNBX2pMVzwtbNjyF211gwlri25q9w
dWTvnrgbF2K8ye6o8POOfVSOu5xF0m05vR8+wVsTjgFqXL17mmAVdHVdRv8SMGGV3T0D/t5RdcXT
OmGHh9kOqAFl2cTOkLGkdNwa8CRxyQAEtdSBNwLOn9+1KXwfs4Ga54P19LpSEYBqtND5UNWfK9nS
j+unwQtIssJjITUG/iDkCt4QYE3yDB7MNkr0Gx0fx9XrMVlah6slrjq4Cm1ltkJIwd5WK/9gyINL
Xhkww9RGJbtVTINK906gNvZsKFbxShQOUk+W8nCdwZ4yDkvSN2Tux6nlyLbnKNwZH/LO9RSqUkVU
TNXfP++0/ICnFip4k2IDRvWEbfVkSPhangSNL5/mp7kHw0z/WGYmibyVJp4HuJVoVBqcjfyEAviD
lXIESHYxT2hWXsBOGQXt3z1arc5iHIphZ6dO+XQDZzSdFZpI5jF3uL6JnL3fD/FNHmq80WtXmMfl
rZ81lK52yEym+dCiJXhHBGpbKIbvwODHQEScaRyUHDB8KFQnRYsh+hEf6fd97Q9AfN4Bw4PJZRhp
44tHI0PAGNOHzzl6bXuWaU5EQ0UsQB3XSf7O5r5qG7x720xj06cutNjiiCmFXBkHQ59eyr0l2Nes
Iie1A2v5HSh/YE23Yx9TxrpaDU8xrOuNY+Uq/JrK1JXB5ZUwTU7PQHM1nnRdFIiUt1kswQX5MT90
Jix16Jqet1Js4BaREl+4nr7wO/0DgXDjrAt5ms9uCuXnS7uJb5hM+Vv4nk3eCoki4oVJp0WO5lIc
7aaAmAPBV4tici9tz+vAW9p+i29wnRlIAIyNpLWKL0Krzz7hPd3TdUZoskL7hOryMJz1NEAoK6zt
5aRFaW6BKgtH/IBGf67Fd37aRv2aNyoPSqdPH1lj8q98UeoQ+yXUGNwK9+iKxA6zKM5r0uIid4zo
1Q0FSpnEjyztu5L0Sq1qqKsEm3UNtm2Rafr4xg+tVTSjRL0B8NoILpTGY438UEPuJA5owhN27HXd
EmNCA0xJQgJuCuhQ1cWYmpJHklxoNHc43xUfJYM17hsvPvoYJ+IV6RGsfYyVvp3bpl3MtuXBxKTB
kn9TBNNF9r1HOLibNwmJTWrkT+0YpZ7pnskmZab90115ziuPVHmG1RIvI+/lEnI7oQ014+j93vvj
4rrOXNoV62xIIAABNGJ2VaeoelthImm4F9uBGjWYpkmbIUPdrahIYnJNrjPHS0D0XnOGwQTDSllO
CxsHwj27C9KFj42yJkJePipgU+h5BAmAaKmgT/hyprIXSoXMwxPTJT4CO3lmrgI/qB5sJlCzRfQL
qj5atKn4tv3i+j3hTo2PhwvDu9EJZvYK4+BVPo35JrbfP6CUEP/oC2Gb5AeGt0rv66dbWVDTs48+
wj24VvvlCp1B9cZhc3rBUH249GRlxqU73GaKf+3sXsrgKPb64qMrbwsGtkHIJKMu7KUz9dKNmeuX
klH8yddMzY3yLbfw2t+5X7zYKNDLyf8toQ4U1/3uDbYIGrQRRGYoFwQjR0I/xVxuJjFF/HbWhNw3
WYS1jOXH9ABuD6/kifQdiP+BLgnCZ4qdNtqzYdOuCYvglXj+gMFObQNQCDTvajRSrS/+04VTFc9o
LjSWggAcosHx64mq2YqwpaNkthOC2I1I6gtBdodg7fZhlvjQf6FIMUfyEcA40hACAexhXS++quux
fxRntUCaPyfooilgoRfQ60+QzEjg7vBC9XgKym8cHPqn3BQXO2TYmBYKfWtnRt2KjqAB2OEvn/8p
3aHrkPYkUWfTNiq88iYDQ+tdGGotyY1PhZA8/3ADPyOUFaRUKFs/+XFO40JrTQCZT0Bsk2gBTL0a
Zoab4beQAZ+B9qcbaE6T0z2zJ8hCqj8w4fYzuxb7zFSMkZRLyB0MBjYSA5THUU6pHg8s6ZlUMper
2qqg0O0Dn1+sl9Y6M0as+rbyLQw3PK+zMxY/hsABmCo8mgloFq/Jm27O0A2oE8KM8g8+qOm1pNRb
IK4VFdtZGbxKIIZknnnSovakP6Wyi95zYYWj9iY5HRRtIudAduk5j58vfsReZ3nyfocGReOOjBzY
tYFI4i6VFdNxSQbUgPPbSURwzKh3q0bHPaoF4NQTq2npRMdmJqSFgHGJH/YknyUnon4nmg+ZaqSJ
o+D0n4L+s5IdZULS2KGRVivE7yM8O1HJbdJGGUpZXGQVjRCDAgdvPdizYlvAlbDHN+f7Dovvrp5U
waFungtxHJ5/1YBcpYMCW/XUaPm/aywc3T6ZscvlpBFCYTVzLCYhDwBd47nL7ZVv9lL2yVvXwdaY
jvJZCw8/O3ZEMnFG7aTm8PE51Fdl7hIPJKJKaYNFQoHr3xTrp+fYWxTmcaN/d9fqOcJGVoBPAUHs
Rjm64ziyicCVN7KizrTTr4CpGp9yOKU11uxGPPkVNceFHp3ivUS28RsZmzXJmfBOlYU2LDg/9W4v
L8W9s4gzMnQoW8NZRyJXY+D/ETiNvEAGQSGEpOUsbvRghxifzxQbXgV36RrNIZ9T3uJeoBTu+zwj
4P1mgh19R140qN8jvFKqiXQAErclCI4IIeaKSlOg3z3PMEBlO+RsuDIk8Ue2SHQseSOhe0OaJGjH
Vh/j/3hXp8NQEUGxc3ZN1XTY2ICmMXN+JbXg761zN1GC9dk0QdNHqthwUml+fvaDYjBPA9d+CXPA
y2RbgDlEG3BMsMCSGChjV7++cM6keKf8rjvA/gMs+e9OVHGqJBsu9ViX9vCcFiIfcrp1MY803k3o
yz6YiPXh174UdO3GXhwz39Wop8aycLRITqkNUJqQbCmqlTf1gjn7Y807rQONlwAGzliVtmPa6186
f/6E/G+84V102wyotvwQdN3MHRRW/WOV8odOsQfkuKWv8m8K4QM8thtxJl6s19tsEDse8AVEqUWO
0OXmUyS9sPXJMpP5kkbG+sXY6p6vJg6dZKcvgFFQ1IfNKLmpJgO66WBVmbUN+w54hxjzaPPOoFex
O/abNbFsqYZ7XFID34931Fb5nKTHmGcT70GsJyhSEWm/fqzmxFjl24wVRUrXkx+M+dMBji2/4Zzo
/w3hrTHg5xTk10f4To7Wg/oM3JmXNyUNA9Ze7NiB/VymNdtklf8KxtwnKlJxXXJfoKcuMvQWciZd
E1uHo41aUE7wKrcM8tC5/UDH1F0JvZ3d3FmdpXmq/WFeo0vLQGPaRFrSEoWXW6AfXSoqtbDgO4Pn
UxpF8XnBmouFX9wKlkNKjhaRyO9YC41dSa7I0A1xz6lS9fFQmoi48soMwdkmXA6Lh/Z5lc4jbDjg
yNSbMIkFoEFwFaaqD7p7BDSMhmJcKCNc5/1UTtc9rDsSXi6USRE/J5UIrLxdRONYH6TQy9oKSoHn
4ur0ux3UfevoGWVaWHVhsmrsOfk+56UNLNZf3ZW21xn82R0eSO8r6Kn6a6ToiQVFTv2mFwm1XBFN
BmsLGsh0fn7blXVLn5Bk161ZBUXn+ku7WPs5+6EtJItUEoySjWTvyo3Kri8HOTO5I8tHZub5fbwi
HYgZ2rNAIv62yM00bL2kNxBlqXlpVoubHawx1PJweo+rr48Q39jP0LWA9MZjGVephRO/JcLal8sq
kn0FLybxpd5Ot1ZUAbngCGYA0Khmqpu33Jpy8QJpGa2S20CF8sbRkblsEPKcjyXB7+ryWHGtDCXp
R7Y2mdSZJGGeUS3424xrTBWG1n849nLMkPZO+YwhxpxkIJ+iYI2DUR2c03Mbvg5+Q/5xLMblkUQz
eydhi8sg6dEGlOtdAMgHGmva0ZUzBOd/jQssUrdJcoeFZw3ND0EEJePl46M6kBoIxzLW6tEZzi94
mAHGN5aSXPkntf+A8aCnvCvrnCkbs4jt0t+gwjt7yBBumhsFWVhmWgXe8k5cpht913lctd3cAJsk
Z7UXTRGS4D9lKhFgL+POaL8Il7lTFTLPdnJX+tUrcpybZ919/TqfcQltne+vLHh8dj0DvHkAlkJD
EQo188L+USA+WSx1/v8YQ1ke/IsUDJpxp5e3FLFMYjpNBUQOBKZXkozDob1c1edZn8NdyloN7MRj
vZypR9PlBuRs1eYLbn+N+8XONrHz5gfEU48SkWZw/JRaVxg27xWS4j+kCqcB8ZBwUKO+YrR2tA7z
heTmAQGOmpc091k7yiOgNgruODTWZZYjuoX5hFOS+bJ1SrFuG3YdytuvvykN8jVPiz35vE5eqeUl
ildCauAy1/B/DCbYFIgX/9SuEve1KAe/Rz1IYTzHTwQ93l3TpmTNTlR1GDOnzDXqqzSXGnNng7VJ
g3Jks7wFbVvegkKacnUgen4cNO0wlxQgcG9+bIlSe5H0Yii6TjNrEp04K/+EWXbmnTGi6TMGARCh
RAQ8cfS33+rpqP1ifeUTP6iAMEOZDVzkIbi+8PxPqoRGu/7dMeAuUEZ7T2eWtzb6RRUb35spcXVg
6xChmK9UeQHtyGkr2duRz+R6Nu0BQ1A6UgsBWYXxmBHBb2lJ3HrhIg+82ubelOKIaoKwJlPk2Gkc
rkhTg7d9PYzu19qhQgKdrVe28u4zKXFFfTSmihZZBVyehpAZdv3+97W4M5ekkkU1XhNVmA+7BjDV
8xZ8IxRb463RS8MRnmEWGoijbNajCS2qQyqC0ntxlCuergWd/LWsYZoz7MWpRhwfmbm1W5+B4IF8
MTNugDOBpcGXbTlIAERGMC99Ik9432J+vzsy4tv6y/VXqcaPc9o3RwzTYrk/fSEqAOoaLb64q3NZ
3Z27v7IWBR9cG0KO3X7bChXQy69XbZdU/pxTfUe1QMZ2s8sNTgQAZsGq5OpdwgTu7U3Lzb+cl03q
Jdu53fzxICcxYapd7pePFkLt7/HPYUT/VtPh6arXAeNHtzeL9sd0ia3MWxHcJ9CrhJ3ztYl84qXd
q6An/wGPh5DmTuWuYQAnGbtr/j2blGggOAd5IKN2SuWGFBo/a21UNIgZL0IXizoh5j/uWqtyYMop
SDz5WYXG+1Be8W8/oD4ZKkK2nIAuNudc1bpuCtJfLLPIgdpr51tLO6MTX1pG7RafGBTNtd1H+pCO
6XG39JX+VrIPtszppHdJzL0Aed2xtzDyLDo6sbAebGJAkavDVWzRc4eH/VmajD9lQFPuaj/Noqs5
0s4lLwglgwMY+96AcVveuqVpI7g7IunJE/fyzIgpUvYOD1iIBYobLXVC9dTqtEQjF1wuo1mBC+3k
ILhYHEEM1nPA4UJUVWOpa58OKyNFq8uZUJc8KhVwNAgigwWzu3BdrLkMjrbb1dZJAEI9z+h/sWAt
qswePOAhs4yJHUlxSOoqGh4b6uGm8rsvnEDUTnB+ktQ9YYQIOzOgHXmYRRrwfmjNHG7klvh4K62L
s1eWyGh/V0GuIL7jNvl6I6GtfTuptCF5aVR6vC+1u8oAYpjBw+Vfa0SK6x6NkwiW13TzgBS9VHa5
ZO55sQldn8PjlvOATKoHHJa+L1TZucwU86agbjLvSLsyg/CqIZwuYXObshTBjE2p904H/UItrmtp
GnxH3iQb0cxa2hg5myX6/RgmIahpFfszeX35cpSV2Js/Z6c/8KMaz08TD8ej1hxzPitHiQwu18pO
4cm7z/bTPXTIL6C2kiTpNp/tLLZFOvx7ZddpnZMrNdhLMqz1XK0rA0/nf+2K4rmAQ1Mku/7w2DvU
9qUZVwi3agE9Lel83WT7y0wMxRpUTH7ENXKCdzAYa/nMiGoiZZntVXOHGuP3dyzt3v1xS34qP3do
bDWndJKJiywvH5/6mDwUQmgmFMWoGcAG3xtwFnehw45ncBmUmR2o+425E+RfxcS5et1D4njAbxfD
sh5t82ffpcJdRtg4GNE/HKSPyuIJmcq6w4Kb1s4w3AJl2zV6++vEVG6bgBE3pScHOdcODMprsT0N
NU6WtwmLzSC1jEZ+Ruo0eoqD7uPxpmyDZmsJ0qIfCMWpQ+2FbocKbBSKnTLAbgWdfQNrwy46RmHg
MNHp+4GvgL6Xt0mDzMIRL3ggrf3Q+SlZ20/EO0utASE+YLO9/GaXvdnv6V6L8F31Pg/tYtS4hJSZ
sZ33VCtuOk7VngCngsRgOgVoTtp9aewxvCh5ZIvLv+ppnYgfXTdN43D1cM+kmmUI4vXQ7Qk8uaX6
FHB6aJ9VyK7yPcg5bRd0OV8gpZHLnHbOZ5PqDYEBtPX1F4J1ZMIKRBveExJ0NNgVrFnY0rN7cuNH
DKN9XUQ2G8ugldC63PfReoN4jOYnkC6z0munYFrUbjyGV3/zI60y7DxNNew7gAyN7e2wBgvXi2QG
gz83yAdD99RJ5w4U/h655MS7mvHggP1T6N5FOs+u0a5gSU/JLBta0FmIdnPWhiNVl8HD2YpKqvqo
zMZfpiu3H+ITUk/RsXoSx3OQTESkd4XO9EqbOL39b6fP2Qh/0kq65iVHHrAqQ14gKndBfPgktMI2
btom+90Z1mlNHYJQrbxci0LWP+0CgJLQpMtJbHQ9n59L36OnUwKo8aft+vPME7jg1BFpArkoBiGc
H3vBD2/MCznIzd4s8JS9x49PWJg2T0aPvSP7qAJ62W9SQ7poCVyDr6RYaHayovRuhidqE3HH/meU
SHGmwB7xhNkUwCPcY6ZSP8sLrl0P9iAaVf8YUlgSoug4AdlXy0enPI2HHW7NdtdheHh0E3mXaWE0
WLy/r4ztlFx0jeth8CHY3cEO+V9W+q1IKMcHwDxGl0MCbc6iiCnP4CfybWgm3sWxKQ0Rud4/Ejxy
MX6QyYoGe38OSdQniVpeIcm12qGMufqx6MEdEC+c/0LxHH99yefkwrHxNr2U1xp9ylo0awAESQHa
y0PIcHvR6GT72NSAfa1nNLnB7oNBTzMADZiCJpgeYs4P60nnHyvWIkSPtEqoGryyUVWA34M8zf2m
OeeIF0Q3HiOZ5TMfhSvYq/Ln1oUSUFMk65+5mTt4upLdUrDAzYd1bbwWwsqf5d9qZ5Una+r0gE3c
seO6J+ioM41Mvg13qZjXLxjD/8XoI1+QgjPm2C+ZGJ/D++HwqK4HXIFx4JdXU36F9v0zAxMTBpva
hnLJa2SYva9exZtEDKhdBLO6nPu/wRyUtCe2UHY6fuO3waYI9tmTTbRoMPQqoJL7tYosqA7uDQLr
FHUUP1b+MprkgWfYdc1IVXE5DID1cNbnlTZ8QzYOe5agKtSN2tGpjkRDYGVWWyA2ma+YND+iAyMp
dr0mJvRU49IojiddPoiPt5Ads9pizAMe7B6CrUyJUaeHTCvRn9aDrQEpZdOK68li9tGJ7Sa0DLSy
wcbqH/7JiRcugT5UO9xKZcFRpHxSXVBFITpL+QwUDkmA0YhkwIlVHpo6+VN7PzyrP/GPf26SOn0w
Z9MhHqyn8jmCwOITPXw5dBnQ767T+/Kr2y3set+EZXQiLhHiLPcag7QmF6d2pn/ye/5wZwuVSWMp
fHSJTpwmt4ADYLQCNa8YRBStGTj6FwK1ZRiyjdDBKBwBu+IkORg4OtJqDIg5R62KCl2orG8BOd4n
pUpnG0OOxzu6sVkOon6sx4HL0NvGsLJDkoW88M9LOAYRmrf49sO/WdW4aR7gf6kZJVAPDSofYZiL
O/0UVypX3xS/Veqd2oq6FNJZ/LdNTiuPMzITMXCZqInXOj5+AB0ueNkJsfdaL/EIbOs2YBdTAgYp
e005NAANPKdFco2PwIYrEhGpeno0nxW3OMIo4uQHE4UQZ4vh8QDch9dkgNKm2pxlI/10rrrNaVoA
JZambzWxpC+5yAPzRj4Zd/h23P1meLo7XeTinH7/ocdZjH6+Sm8oB3FVOEXfxTpWZnhQ2+oJHfOh
BAbiIKozwFgn0fq4NskmqXcNvGH2WIqDgpbZkAda+flz0jzGTUSGCjSBCywxZSt7B11AkK0lOrLI
BJdXkVq0vIusZ6R0wZz5rOVyk4hUfTR3S4BvAFqqnKNeNTJddqYnNWYAnsDiyn3TOr27JYMSdgYj
73+N/ognoTofgVp7OgnAwtuUw321sabAkUF1knyCM/lQyAhmjmyMsFbOFHEFBucLsZFmFHRKEwHP
+9L6rJaudCUjR6aS2HuRRwt2mbbYaULRsiy73DcUpnU5eWHrCy1x7qZ1s7Lpn310fEZuOx6+JWXm
hWhVXSQc/igRazt2tINWTPldtQxhDT6YTyxFJCpOBwryV/Aiou3lS/YgEm1mrJbEYFXb9rHkUAzk
ElgMyQXgx0Yd71/Oi2cS6NfBZydOPEe3oeYQ0ngqwxCHf8rv5m+w8ZuvC6S4jT+HJOsDFOsPy56O
IeYmG1H7oHqrMtkl9N3Wkp63es3UZX61ABnigVswgfDnZIrJFEaHv1mYbNt2U2aohGr/DIQStMIi
lmo4KghVHU5iDj8d78mmspF0YlZ3mxUQ73O7vF32nhII7gNL5vn7sgu7P3h6TV+acZx5lBtQM515
W7AHKN8oo2T0Sdes8PWOHBiLMEr+H41dFh0frsf2wOb2nCeONX8MbcWfoT+y/CspLJpOOdyQRJmz
m5fZoXgAAR5qBXP6T8cMhRXMMkoWwfAVIjdvZueWl0dlx0M/TE+VCvgkMBlJpLE6T8/aFFh/ry6o
ZOqhIUGYvr06oWKmjQDQuApOq4aVqEEZoWGCGTej9S8uS5pIusB2CgvhZtIWCoUqU4bqeWC+zHz/
77nlOrOR3m0v+2+Vu5ayHIVPIPw+510A/n9yx1EsKYBdmFz2CpzBhv7ZJbrpKA/00QWHjOfIROzI
O5w3I8KwHPcginX9D1uL4O899923zXEINWGUpoTHXOO2qALSKKOMT5FlDwq9TBRjhtRyZzgeLUqT
lv7bc5JFdSVo8FCR1HxlkQXqi3WOxxjLInRp6sS+YFk9VkRQ7vGawpyOmPeOFi9xSufNSlLbrYMD
knKO7J7xt4K9oDnGXSlL8KyGwfeEYHXirl1r6qhKblku6BUUtXS2f1AxhiRIQqioCSqOER5Zt1kA
puHaeUqPJJXRwWVXD6Y1HiT4cESckOPeZ5GoAVH31vDy1AJhg44+NuqnlGkLjXvzfqzaJL78uYmh
mfwomzFa+Y3+5e9qtE4SjJPyhT+F6A6Mi84laoCRv4Zo8WVlgztj0jtIN69oEHkR+1DDwgZCEnG/
JX2844gC/mK5Ashwf9NSVPTEMggXjwqxcG3jRF0RRZh9gadUY/mJqnk4kdcSoWI+5dfy14p2850m
lSbr6G0iu7gWBevM7kVADtm3xg6VmVu+md5LHw3/4smcfFUXt6I9f5fR4GLQQeGuZ7Dkar/uXdfd
DfyaXUw+EhCWAd6yeVlkU3nIHD0WR9YMev7VaMJCH/qhwgEAqpQKTA6F+dUjy0+YMXM2CemmQw3P
U0yFk4cSlB2SRQYGdK71P+uy31GiXVjVQJpOH8sQbvmTbi4JeZ/yauBeppSJC1Q1dVY7CeQoZiTE
DIighvpzWeoo5mibLnkYhRnJeNC7fMM3z1UqDdJ9SdCKnXosgagcnNcrhTeXZx5apV5Mo5T1iu56
M8imPIDpVWdxlpmqifohdWcGVtcmke/nVQYrpWDWNKme7a023/uBmQYPNsayCFjTzd8+BNo/Y7ti
RZ7dm3p8TfukdSB1RzBc8quV2sD9gNar2lOvqGVYmNUQcV7/eeAUQ9XxdIaX6BpGQz8dUpu45X7E
skVAlr70W7WWvohuntL9dmPduL/0WMJtxFZ5ZPjwQWMXu8l11mXvlonScIcdAp5KVCqUufmZj5F3
Euj4pGe0pdi1KuYoNJamr/+dcG9Vz9aTPHcrAq5Wphtg97bcWIQqdLhXGUha8spDVC0LrajVFbB4
P4LHJgtxHb+d0hikxg+ZBOev9pZn/+1hTxbfZmT8cHocWkAYS3+AVaSJLVGV8E0iUlL7ui3dOqco
TUJPAS3cKILHcu4Gx0Ow9DOVqdEd0PvbvGyM+pz/viK/vXeXC5SN6+sa5wio7H8hZpTlf3tQ/gGk
7y4XRDTUOKpd8C+FMwwq5D+7CsJoPKOxGVTpqB4xcEmVAW9U+XQnODvtgCd2cPgc0VPGSmAz8QhX
x1s8KBg7H9VOHLHA3MguhU3J0fFLck0ZOY31MuZxRtBz27x8mrqxAra8HyCx71FI94nww0Akvts8
9+4nlSM+wAkmR39d0iEfBbQOGOTPECvM9AuHK2pmu8GER8jL3YrcbNm7OlO2lSbZNvtzySk2//Hm
PG4eu52u/FWcG++iHrqpERXo1Jq7ahYNyFEPoRm6XImfTcgPa8dd85MB5yi3I4Z1oWMBm5yYnbSJ
ENmMB+PCbMtoAt9nDfzCKOKXfeI+3z8+nV47fKbsKW2ScxJFP3yxA8dv9QGGoUZ+GkTu95vG3QBa
5DkGlDhJ5WwT2i8bO60RmvFRb03y+UcB1ryIR6YGVDj4ftWX8pSW/qW3nd0dZGjBimGo9ulFNH1j
Cxo1tJXq2Qjgcnn6knkvRHrC9M0fVkdUIP9fDqew9ZZeQJQyNPbxc+ZNpLWMTFcg2kQ4qnfQgAkI
X+sdfh1/ytDWUTZpFI5xDL4/CLQZEF+hTFBmJL0j/XL4ZeBGawuWhWM76o71xnHzAaG5o9PqKqZ7
cUQA+qzDOSu5ykMrt7xi8HFuZMVLNwBxI0LUVk/JZcE9rJI0NqoX/SxEb2n8srtMF0DFD7RbUjWf
/gg9Ersn1W2h/x/NsDKMAGIAtrqli2bGMx7v+dj4y3BmpPYd7b6y107OEaYuhJqfRuTC431Bw1vp
yNYpfY9i5cGLeXLB1Phmrrkn1aMRDSD3BfMeX5G1x70F2eOzcLidE8ftOVSCdMzhRL2POG2r871I
Vtk/u7daPbC4g34HKf0D4Qa14K1jJ+4R+XckbDbdE/uGuCpDhaI3ghDvDTIv9ndsit7vF5N89VZF
2c9H9OQl71B6w1IsWC59o1I4AhpnhH0Nqi3x/+ZnXOL93xDL4/Hqx2i5w3JQ8U7UZ/5O2laTXe64
xt8XemD0YwkZ0d8K5Qlf+FKoPR46HU+9yp5MNx/KHokUuKsthrumySS4iudmQDVmP6JQh2KIN4we
VqL0uL1hJNp5ABYemZ6UPGSYm+jpZDjURFN5b4D11iTcjm50NEleUWNE2KyaA20GyLp8/Z9UJ1y2
b2ls6peIqBXtfK4+WHJMh0tPLQTTQMypuTpZCf0iZa6BXINkBcxFS25gyyIzI4Uzc4Aw6Y5Dt6jI
/AwVD3pe21Bm45wRh/fJlkS888ccuxlcVWzjlBtwLzzfnu7onYcDrk5ktUS4tt+Pr54Z7DRYezfp
jRFWWOuHqqq5Ecg+k2w5hOfYxwcwdAso6f28k4FLk4f9n3CVbk2kumen/k5Y4iIaGbmxNyZhWGTR
HACqYLkWsgvmYs/BiUdhSOtGvL4TasqIBwnaX52inFvgs+kcVm8bKH8Z+or8hbzw6JsWbgHvWM9l
t1oAc1U0tOMClA/ATuMt413d044tjAj0r0I00tloezhfCYk7jr6mFfXMmdMJYuehVHI++Lg2SRru
cHKkcvYaCxYt5XTWoNysKFM2Zmk5fplNv+AxBf1mL+fiMpko+5odavoX4jPV4l/6IGxgIdPw50Rx
6cnGvSB2HCSAttKb8yBk/G3GJ1VDsMVAMzSFYUnfq+qPBrZhZKhtUL5cgHi6O0+xv/RG0sC3A0Z9
pQQ/cULuLItBflWsIk4XS+SkdQDGSNCQK/0ALCvU96U8sfhdAMOFO+Gms6i3MZztbs8UV0gYO32J
UQKhcg+2eymQ9vN+draQPho2NWS2HMMm9yKb9WHHKuhZIrMDhQINje/IwH9KleaWshXICVRPtKWI
1gO2q3IdU8pgOlq92Uz609RoRbuxtcZu9nrfgGsNwEpqYr1hqnYXWm90Gr8pZpoiJu8zhL9aEtXU
jAEmXQVZyNn7CvuRRBp52mGLfOY4uY1txezNFQupvMB5AZbSfJvSFqLaJRnh4kzwrUmgAN2uzqaE
cl/UchTmJj0JaHDP6bS5DZebPZzNzMXKIQ+EC8qQSBjjQ1YJMvaIqelHD3uWDenzdyWGIl54bl3U
SJIR/HwGY07OUOS6QPu2FYO/j5O9ST60tO2km+GG30ickoxn1F8QT8nQ5GKJOb3QzpGa6rWt12Jd
8Iq56hIl8+b0mRLZsbj0yRkURekcSozok9Qt2HLhHh8QdWkhiHCnmM4YE6nCkHKcefCz9dr5r3VU
bvdXnuWtdqSyrh+Sj0s8p2EWsGWi95iiPEVbSTya9MFnQ8zVW5F3AB2JQP7HyPGGeEj20IJeudmI
XcQksNlxu5L15+ENsbpWGtPLjBWtx73OaSBaI68tjPUql7a2WZxau4LTeHJ6B6eryHcjxZSUQpSF
5R5kgLwtn090pqA3xEboMwbARYpLanr2JVWiVT6R4c1MRNTYdovASR8GHI2YUDWqSR0v0taBUyqO
ROfQhw9HtBV+wyuMQlxmiciTWxN+AVJ1lRThR6HWiB6M7H0iW3OknbEFbMsR+fm/8kwd3+xHUWOZ
mdaKwMHFGO+SidnY80HPfHQXe3LQpAhFk9XlPvWZUQKTf33QQQ5VSDb6nU+dfgc+WUt767rty9D3
sTdqn20kWuEf7/QjnyfKofc6FD8MOY9J+jZeT+MwFno5oJR008xBhEfNYVJ1ACshPg6fMCKProsT
5clVgQvklpa24oUjxx9JcEh6hA2s0IeLS6ODVnbqarysOTSfiEmTs8jSS1DJYw26X3h/e7xD5bQP
gDIOPzejaTxMiQIF/O6jR4SFJgoUEUzGvCqrsAXfS5x5NfpOE4pWq0koOsCTJ3saeDt3dbnN2G+z
KhOaLe96Rk6BTVFShV/97Vut8DipoelHFc1FrB34XtS1IObiRUgpVBq5ue2KCf9szxwataxbBWcE
YUPpm7bMwmL6g3+fQmqsP7k4nJc810ZMIZCngSTHqVmReHOc/V24Ko4QqKoFWU0WCnFAFDnpgaYc
AJ6hpK8YRinfvqr0nCDeXG6GdW4VPfGW69IbxbOf+Qo53Nu/tImsyK0wDScaCtXTBfZF4d6QFQX/
9hfAXXLifNoijNPi9CJFPFc0i7pameS0Zx+qSbZKSTNDQB1xgunixyzQ+yOQyVPtIvlb/9ootI3s
L1cY5+kDB4b3ETazAU06L4dVCYwoZsO0+//HH4tBK358zNA3g1uf2eitYPBhUNy/fG7OxkiEmvQ0
4bhZyY7eD/muw5FJbv/seb4yXT2AIwD7yjqMt1E+oeGgp0D79q9NOOqpT7woK9kVzqFg1o1NsjCE
M53u+0RJhphCM8WS67l0bKhNd5TQA7JxJK2N3Hh1BPNyKks1wnCB0keeBy8roW95s2R2AHscl0aO
yagC5UbDUYKQTN7t2Whz0AnRuCSOwAuyAC1fDrBOZh5KQZrpTc82w2fd2rKodl2+rPpjqJwTagze
2NjOYp4FzgoZyW0nQez68WaG5Dz+MnCb+f9AlINLUU8nrgXGephqrGt1ThKW7zpkcDmi6l9yVNon
7bJJFG4BEMhjJ25MiAejS1yxySIFyoKG/soy8H858KhKZlP52M8mRp5I8tvTbluJhnhKpGfaCiwK
qI6RfRbhik0MDf+APXXHEPbh9BJeltihzQtVji901a1uFChJ/m+cJW7kboeVXtWphGv1V6oe4VVN
yCgnrDHVgZ9ZOFisICHvVi2932bmwemnax7na/ugE8x+Y1c4NnGwFiv6Wsr2YxvHaZSeSbIEbhsd
9kW2lriSpweZW6NP+4zi81zCBqX1WaR6OPYZ2gbsPEElJ/GTUoWcNXp9WtT7S2XTMTIc2Dv56MaY
AVtcpiJg66LOkkWXO+zImEo+1QHfBhGAsDxb2JNa+URqJ4U+TgDEcd69zKRDxXacgnMB+i/iahN4
MO+50LGWDjrgw82B05Zd3GHQzVERSGuA8xPJiEfllTaFCTFMQSYfFDNX3a0KQK4pykJ3MggAzbPW
+RrJf8F+hSC9bCec7i7Pc9c9s5OcSnaGkfgo2r5ZtHpAZIzGE2wog3RF6jdoGWswRP3juXip1Ep6
vEBB+V0k0pMMyP3JKZ0uDrTGdKo0xp35DZkw3qo9yjXtkFluDSW8vsP+IoThHGWEk/EUoDY4m5iW
KIAw9UcFhWvYDVQUJ++2dWWMEP9brWiymQE7NG9mr36RQS7og+yKQLyYfMZO7dZ6973piqIin1u0
qP8cWLaXwul63FKvVpD2FbQzv4ViCJ8gHBK1GwMb39je1tOhxoqLNEQg6YGVobcH0sHHIF/P95+S
rXkFRynaYPARAY+f0kTvOk9q1+w9OITKTCgjZDWvkJLZoaE5lutidZu8Dm6u861OfDeS8e2Twsq7
m4NW6qojUgto4S2RSQY6jEoNmD5MuDzjEwpnYRC4mQe0QgIs6MkWJyTCx+zGVCRYwkX8uBiv3CTF
hv4IgfvD8iNcZov8rFTYm3+0MMwT4uzs/pXIenZ1JjND16n1b7VyaYVYhsRUYZbDdisnHZ3uwkUO
PVQ5r+Xge5YqHLZeqtsnzLNjVK5yUbJYnohF+agtXqKmIKJ2qQjwFO3z6NUWdCa5HdDPUKasdOsP
6tN2o6gBt888tjHNnYp6koIoMzNOVa9Tq5albMiGd5GjmfTxqo7oR9SuDpWOCDo+9CxB/YEdmAmu
DniBfu6N8S8cMb1dNkNs2hsi3ntcCICgBUD0BkGyTJlDqEk2SWHfj6YClf0sDNDZlZxPTZtnc3Bz
oGJuKUl3g36OcDNm3rv1Esz9B8RY5/IRo1zqItv/3SHU2FlQeUA0eXoQc+iecPfvHrQMcDB4TWJy
nMngsu3vn3CogZ7TcPku0hAZRwIjdmuiTT1j3wxveeI0CCSpQuRYDufO8kBvbw+d3pXlhSvgWrJP
r8uqHnesGDpbkDVZXTSRr+pWUMH05+HSIsBxBNcgUXE+1t++CWZ1nzfrJ3ZM8MBUPaL444Pbh1RF
yJYgEsIsXCZXRMSwmnho6X1ZWazHwL9SmL48OwRC5X9OQHZu3/8Q/wmUxOAemfxroWR2ww8ywBb4
bwgsfbrEh7hNmLWbBB6/GWwma+7/urQ7i1s8u8gk0KxCGSC1cYH5j2VlTHf7HfvzE23MVCICY5sE
GE8AlUf3WDW7seyjfqhXIuZ1uiddOnNf6fMxX/RQ7w9mHki1Dio+qwB2oX/7nJJr2gfk0w1h28CQ
RL638b9lGHnwdjNx/vzw5uHwZjnUAoJG44PMB8k+PseYnw+j7okXkRaEsbDwiLV6jqdY61aUqDbp
WtkE80g3mdNRptcwRmx1ea9eHDQNVa5qTKFe7XUwpwusjaKd2r9FLPBM+noVVy5vxM3FYVvyIlL/
6E6ZKp+JOa42RBMfCFObiziAQvd/mXFH+Ba7po0SUD8RXLN38zgA/FZhWZbhY+LEO2D3ysLe0h49
QV2153FqgI3HEbhovRGOCDe64T16uwgOBjLuDfzah6Xy0oEr5QYNQ5djZdxhTJNy36tWHrWsnLgn
94ITaga5zAjgUCIj1e73S2h1eBQCrChOm73DRfqEiFpEAU9Zf9eLLc6h5BoMRSuBroylASF3mQK6
QgXilPLriUkrkSxg0PIy6bSTJAtACyBsCXPBWLaXYR584ypL58C1nblKkiwPQHLEOcwxM5fHoK8y
Ff0g7kq+bSoF0Z7KXbxGTrBcx8Dt1yxWyiTUUM0qkDG4Sas+qScO640vV8LRBMyjOwgecUzfVdeB
QbPJKxV8OpjLjBmZemK4DcDa2WAbioxcyNzHKQeuce+Dj92bDrxXzfY5liNNQRX9bK6RDZ//rkyt
YhvNkLWEG7ji25Wyf7Q+HaB+isErO5nZOt/4R7nk3gWMxPhGYM58WeDqLwS5ZX88vOmWDMFuHaYA
MNvPv0Lh87ro524zfA9x1EMq8n0xGoUzmtHGmD0S95kp3HIosyvwTT5fcfQVvD5gDzIZQX9iOJvW
O4oDWSkPXLjkccvqxE3O7difQVniRICaUdzCpLJSQtAKIVJbkRbJ9Ijd8WDQ6lOVAjAisMH+Fo/Q
rn8J9uhfWEuqYriUAFL0FbjNAJ8TXFY1GwIY3rXA/eWNccjTbwWsF4WhMxgDpbR+D+N1zuQeY38Z
q0pGGceLELUm9qpftVPbiUJ72vYu87IFX6Q8N8dxkRHK+/1U7pShILpIjUOvlIDVOLDgkBEMnDAS
ZP02lifXbobYRLmM0OrifFvfWvUX5JWV58C9pVAw0kXHVBl4KE16NamMUehWm8YsNFsfCEn4VYyl
Ew0SYR/P8ppqi6/JW61gqL5nhazGZcNVLJtNlb7jfx5gGXkZlDG13LEGeIC6WseA5YP66UKQlu7r
gpOTqHVeiTbEmOqY9lKDzr5Q340vysY2ajbSHBQZhhWm+V8MWVv/TlHBHyo9dalt/Obe+bsvvDFi
q9TtTtawL5+4mwotWkiiivM+824kTMgrqn64LSuDYpx5VL1oUtaEmpkEBZvunC/k9SBn93m19TPv
eMF60JwRDPc8XcQgHBxVNyveby98yn4BWvIkzPtls1Rt5HaHiOBVoo4t8sMnaTkMpq9YHMeufsCU
Rzc4U9wtKw7xxMWvYhh3IbM+QpB/93quwn5iuU/sq9tESY4Ry89avHWFYADDgJsHKx9s1RFnBhkK
7EK3pVG2UdF3L/4VJmt2iikJV5yq3luebCbKHdCR3A95k78ZYnEubAuuGhEVcj6WFTttsWrjvRxL
gSPZVOf2iqRYOcoANBCXsAfM9dd7rjlPntrt7f8vA146keaHGzkRl1U4rI3yUeYfiCTqwwN5B4/e
Di1FNhGsLX+GFDYb8dDQ91XHQg2SNHZRRx3XkKMVauQIr/tkdpo5kVKE5YvLOCnF3QgTfmeP4mFv
8vr/VruLUhgCWlglhGxbnQ1PjeATQqCi+QBUqJbe19SQWEgGYayTY1lm3eDBL+PYhrtvJr6FUwSl
IlfWUhIfo25QXmGZcJacCBdkWozWDgX1EDhAFwJud4IoeCim2LWvg2T1pxGUDr7W+1NwE+dlzbQI
PqXd7nH3l70o9vehGqUzQRjXWCgLYTZMEmexEQyVq5vaknCl/GjnOZxbBA4Pt4aBsoQppgbeU0SK
SS1IKz+KUUNDlBCVXKiMsl79nM9w2TIOdZiomdETqkNsKbaZhMHjiP1O2ECtUMw+NrAWXtGYe8wM
9ID9AEuzg37uEOCprlmvBPqxocjBlPYSYSVwoLelbfH3++Eg2sGN22IQha4OLISQWybhwzC3Y43d
n/ZF04Ne8GazKtGqdFVqo8Ab2K5GRcvSkr9TIa7LM1E9yvexqKIu5wKwhaJJehoGt8Ie+3Ep8FRT
vBc54fCGlsiyoOqEqLB/fBlUz7UlMGjKwt5cgaaynKmihpp+K7SlAw8o8PP8IHKKkzkI5rxxiPD7
ovsgby7RzchxBsKpNj3LU50bnuUTvmPH9FmEiVin7xhd9DOcK/HORSCUBDoXYZm43tw4pDNHpCLw
yFcYE6ambaSKiabV1DvEiRpTHONd916AUWnbgbMGPpyQsrh0cGeJXgjgyLPqdbgT/xAs6VQtyvsc
kRdPq7tnHqK6D4t0SG12rHg3XIrFdBPclNWELGPeyrccHC/wQ5e/dKaYWsHWiGPBKSNInRZh5+7V
EFIP3h8Ma/5+g20EFJ2hBlN1oBLoznGt/dVh2UAOa2xjg2a07ckEL2d1eKAcU5vshKDAyXDbhRy/
SEByCOirlKWZ7zPu2/Y04FcBO4NoqU6YyXmdXGwcvzISB40sM1S4Se3UfaSZV7eDB14QkLhDMZ4n
xhd8S6r6J77LwoyEbN5QC4ClH6UK9u0z3xWkqy4assUR1kHlpDnFz/0yEsaeEQt6NYxHXsoiLuL/
wwrflknJSuf2NA2iGZzyxDttZqApeyry+GhStp8t1VlLavtMtRvkENwwlQMAC7uBKaCpCmEnYtGp
GW6X/P+nTPC5bI73aFZ3ZHVmf2xB5r3I7nK0dOMcCNfvnnADvfQT2EJf9R8/AacWtAAGpudkzNDk
YAR+uYpsuHos6+mHVQVdKqvRe5lzhqaSHmPiXuBZ1ypQZQ9CAhkfOhjU1SVnmrcrAmInbAe/owPZ
cLSZnLL81f5XZfmoSadhrLCaowXHp7xp7POr7EBeDVjAOQw+EH6w1QUVIOHYqBRicSmPcOVjoqDn
6yRq48YeQfewHuQprs4RnZxxBKvrH92mmuNu6ghf5+3v7hbd5l3apDdKnn2tHW6u+6lUe7xKBBbJ
gyUTcmejrtkhZD3xaYT8478AYPR60c2FLujemCSy0iMLwFqW6eGFDJqRe58jHWk3b2z098Cr39kT
hgE+g3PikeVp00cWZB1zHeFnAlLkJPWteCCvTrfKSUPHw/CTB+j/rwMBsy00wKXf98Jr58ec13w9
8gvJTVsdG9fLd538BePsydJfEYrQOpaiJu1J8QiKPx4+dpGaa0eTngHUO/2LxSgI4GNe7q0K/N86
QVFf5GbxXO98OxORXO9mIKJDZpPUc5LnSbbYNJGc9HjZOTgDGznoqFQVpLLZfIcjF7fjuIecjLET
4j9kpeVUQLJet9BRmfXoqTbZbBbvif91HQU+GarBelLSaMAmzZz9jgBzmoufsiiZYC6yBRpEoOio
/pmDpxuR/eUzmTsiQlV83Tk/91UkpgCZdQ/DtuDFZ5vrzqqOmuxhjFiCcxMIziPqQ/PN7n47AWEI
jx9sdYK8YcYVmQpcZ1Sob0tU/PYBDZiIlTLq2MG1bDRaPIB59+qB45rNugb4fvrPPF4pBc2ytX2m
qFvRYadIZ3pOR92IUupKo2Xt0Y3IBqJip26+Yw2sKMShTGrfPq8J4A5TSkeYA0h/4o4YQAlScAWl
eUc6NHcZsU9HTt8nWNbAQLBcFMqJDNHzwQwV9lc6/JYqiKwX+qhFRwkrOxpqlTh2HudhsOC6aBFU
7iWOwp6YdCjjFRgCHNU2I4QzWXMk53vTgfWBBerZpcbzyny1e9XioGVc+zTLy396azG/CEpAsV7Y
CTUevqNftwnV/kVXTqEOp0OwLvqZ6CU28Mf2FkYv0twZmhfIG326kBKcBgpxh11XhHOO1X1NRSxf
GFshujwLiLuu0GFWZUHjh+zQ446oQxGZCJTztC8fM1ehtLpQW2ITCotCmd9cwV5DBUy9dP19uOei
sxHnLD7l3YJg2KhTuFFxCtR+lZObE10uqC+oyInabX5lKk0xD2YhWHHwLCZllm2qq40OEB2nAdZ4
B30rkj01j+GLaITJOUew9oLTVhAXJHJHtQ8F126/7Jnt4ZXfQrEA5Aqs6zkZV3p7WgeH74kehFEH
VzYXxf+N0k8PE5Fxu+uoFxJYdBg9nnjxku0WpVCluVY07zWpVcE4bBGae7fGWg59Vl3RLhowP2l0
qAW+egdJe1jkLXEFo59K7ArVJHZqkWymte3tO5JIoF4UoxPOSZtmYA1mxwhX0qj3+JMJ18Gc/Iwz
wpT0pve+1sUWbUsM8fEcvQrYtVwMUiWU1MCr8A/87bqoUJFwPEGbtP5BA0ahmLcE+LvTZwIdgrYR
0P7Yy6TsmBEIkSzBj7YllHqymklpXTLzSjGL3rKZUmuXSmKniK8Cd/krcd6ssFiVeSRZnNpsvEZg
0UccWS0nzI1W7CVSXmqWA1aHeV57ogS7rOPvYMtvH9aK6GnWAJ8a8AFFuvrmRGold1I5dvK6eAQg
uFihSvuupOZ/Mp0sNGkPR7MfhTZnlDV61c2DW75f7PG4BCHOHN3npbWAjKSpSkPFMxl0UujAPJL6
yp4OMJuGXDY+yVEX4femrlpRgLKToDm2yrrtICsqnVGLsWSZRbHodJF94AJ5OyJQSJK2pLdAePT8
MFKoU0KbK2gC1mTswOJHreonMw5TCar1WWQP7zDfWbDCreqKxyM2BcpXfhrxnCR+/qBE7EGnKyHF
tRDs31AI1fNR1iygOe2YdbwwMoo6bFIrYl8+2GqFGmdM8URXu/PWHfUBZr3yLvbAW0ppw4r+j6xt
sMycNqI5f8PdH0IufYX8FA4QeBPOpvKlbDoS6OKPL+WxOi/PT942dIOjh3zpVfLNEY0eqgSMypZF
ZSDocaAaXc8CCZwBSeXeXCw1rdyw5trWy1sUJzsBFEDtjLuVwQjLlpgHUrl/z6CSvCl8fJO2kXkq
tuhzVevAOpd79naVWxHnvmmOcMx4SJnL4LkXcQeRB6e/T44aG2JnYX2cx+Hb4m+yT0D5Yuwe+O/S
/9aEL5z81ljyp9cp9HH72vDYCixhQHKLBDg5+uq6dE8d3JiThUfPNR2X+U3t1mw76zRz8hEYyP9P
77vQ6OyBRAllUpyCKrnYQ5V585LnZcA5z/jF7nHia3a8tGzrGeakUSBn9pfis95ycPTcpDI5SpKK
WdeBl+B73MoGmd0+YySu46PbUUjRVJwIhIaeXLPClGMNKdbZ60WdQ22g5I/YerTgWg51S7Q6xqq0
dJrJgUKBuwDzT6EjOjCyetk0Vx7FtuWs7cYS232X6Xen6zKoKoLqFtP0pj4rSwNzLM//w8DJOC9t
vj0s3aETB5hTRBeBoxZhVMJcPvPnhsqyiKcdxcotfs5JywxSChfNU9Ff2oACRhlpxWPYA7xf/4Px
e7CtIW8EZyiWmOh27t+jeG7EkdzTRmgdThy0kT3IeYOYBqvmeTHdjTwu32tTW3wETkigfk6t2pqP
L5GGJSyllnI3HTBakvuWpSSVtCn6aT9jJbJ/pHykH1hoF8A+3J5Ccfoaq+lKUsy5Vbe5AkEVKr91
QghjEWHCk8G1HMSm6dBMebqYoc+CxOB7Vq8oJzz7UZsp9rHDBvAMq68ZcTUKMtY0rKUmmfF6ji9v
Q9pDERN8Hgk4kIo9xeolJNTFZfy/ZaKhXS8SGrxI1ZkwbhCkko/eJaAUcVJ8UiIMovF4g0ggfs61
U1G3//hasCHzfX8cmvrTnP0VyKrX8LUog3sQnQ9hMGKvmY8OcUfnYBmJ/YWSKWtDeCHUfSoz/P9l
smT2tsiiiuTkbKLyCnjLRr2eGyKcZ5c7HmIXitGPjfY63RwIo9AnBdMHFQGbZXg6CpKhSVEeNxyw
Hp6AqwvakO9EPU8GlQt6TkbtoSscNjDel6e31BFd2nVNS4sEZMnXvIqT74MYfAYOyrqO6vIaLMkd
vIojx5+ehkEDQWs+LYIGM/Bi8VP9Iv2NBJCmW30jOjFFf0GS7qMAakTB8Z6vtHN8iZ/pMFHofAew
fZPfzROH77JFPvj9QQ/N3I4uwVs52yI7F1MiKH3w9XFnC18Xjl+rjV8ldPvQTl5Fbjvtq6yTWKYm
FhBe/Wpbnb50x2RYPuz/NTew0qRzGRTT6r3ubBtRfSM/TStA3A0X4gfRHmU7b2w6f3F/zECVdWFH
umNFPpr0tAHEa4BdBmAltPcJAByHKAJJqDlChlWTxn+OqWu65NYDIwEaaBuLuESbaUn2AlgrqXjO
GDGj1crmN5eC7OWFQ7xT3y+5ht7sSerRP5YouN3tbTp05TSEqJfUukLPuioocjPdAM/liMBg+V7r
mqTBWxt5ME+Mf4CYeqHkaTXUswTc1xcH0IQPXI/DURbQmLJnfDp0YEUbGIVWUANzSZQUA6fDmJtn
9yNLnAIBcYzZbNPxfCW/dVKIpT6ZkE2SNpuNAZXzXE2eRNIRyRqkvbun9xOFcRN6jecN1ifO+ez4
VZFu01AzkvfniMRwwtn2rxqZaApT5nzh+ZBt2kOi9Gt9c9fXv3OEiNJDt1FYyQc2vuZeIDEJP4gy
1DK7IY9OsHcAXx/Sy/gN29dyvHYDSJzu2mXdyXIzOLEom2F8oAZuOn0ASMnyVhBOoWctu1YUn+9B
7kihw7ASVcwLSCsazO54cPa85QPeFP0dN11QKt9VtJj019DumBcj4ZQTbBdcr8e8JNVRbX7uJHrH
HOLClfjviY8AqcM1YmdCrr5JT5HQexbd+dqMcow48Pttqh89LVFLPVxsCdnvH2XJTjx2eb8XJ2xG
dG/SzhTf2sLsZ+gMtuuGBfVmVh7R1MxfOOqK7gLdBiUcXTR4jL4SYz8T8rrU0k8wAheF5nGO1LqK
AAA9kGi5WUOcv2M+8088rNtp2isS8+zHVnhKkHLNpqKl+Bds27Y8pzNCl3SmroBF/7jxhIQMlCCp
VTAMs9YI5coLjqcHnNq8Eu/SFZoUL3k40cnLqalV20sD/miQzZUk/Y+sC94BC3y4SBTByuKZJFqr
aE6u4I0l8iDLp/jMhuyDRumWI5lVacPQfPjh93hQmbuRMvCHiGFF+4M0XIDuTVF461f1ACN/XEea
3Zt7sfu7JhbehnK23rm40wFDmfnJFRRJNITJaYD/stJBT91azSuhQxr/CUvi9wWspNfb9YeuzIOQ
TqTmuHmYbp4Iyy/LXxBSMkf9IIfyM2uocBQcsVZkyHcGpZ+y01FwFFtwdOPHOgV6sQ2cAHUA9ed/
71UnbYI4PKU679haXqtOlLPO316YZ6MYIvom8nXFtn+sfjYX8ao29eRH4c68/eXoglHiVOdtoDy8
51XqJJQXxkgOumgcvGF9MYRXuaKSzPRqc3BflZPzkzKHas+PBo6Ej8xwQrZA3IvjCB/audOz4Ouu
eGGdyNjxJ5iMQw50vCHo+jZSMst3H+28nc7sBEGuCCcpHPEGGrG6fL0mbxS8XuJn+kbPDF+hpzUo
hmbkQHQk3jd79cimJ4IHtkweLt0idL/fSKlgKgNrrz1PK7lVqrXAtvAqPFgTNBTJhSNxcw78pQvS
ra3BHq8Tf49uFnykXmIoj9T41C0V5EB5BlAXr2eUuM4E+Ws3VTqFXypfKInVTiblNnBo1dbYBggd
6NFxWQknGpXQ22m3n/jehmekSitKKHOcGD0Z2NEIvCKT3MNL/G2lBipyl8RZcyxX9J3qJtMnz53O
tzHQDMOceb58BVNSs3qkRP8rEJ2xCUEMXge0TzvfuUttFyYKvgK9pIjdijmMJ5HAPbO3ovDLJ7Y4
UacAHdYFpqsU25KriYEtpI9DIPYkQrDbE+m4kB36d14ZyfaToeM+LKqDgH+oAXkZZq+s7g7NVcOz
LeK2Ht045fzfvgW89ii8CEHYi4LumjXUOQq3j80+hEL2faOPDg26W5do/sH9nMi9oLnda2GBI8DU
BioFe+VrTw0FAE3jugWpkSkArKDeAqjS/9GTNaCByqqYTtwsRlumQv/Nz4j6MJdkA15JG2dIVHo1
ZSxPRkiuM/cIeXSoU7wgWDCMUNnZk6neiE/+ABDz1o2D5vXJepii0He9UeJHkTyTQ7Qat95dgxxL
O5XFS+4ZoiSQhQ++AI38AAjCj1SK2SLpDkZRS/8pcdvJZ5CCucERwnyjthwUJqvtq9FE3rePXkU0
FRzDCtud3MacKpcugO9uN6+JTwFBfHoHcAezj9W6w6gfIvh6+T70+2c/Ua4aeSvtoIhKSnMp6y6s
isgoiRMoCRrAgyGDZaJtz/kfSk10VKSDTiIH72FuqIef92l1CMJPfOEnT9LRApDHi6IdfbkUEij5
fdOipxkKs5s7O3f8ZVZR03/1w554z6yACGg6loCf8/ADCj8FaLUJSehrBj1xeM72Pror9sfaiQLP
C3aMYh6AdMYwlyY0TbeYy7hrCCqQToFW4ZhnBHtJa/mDrTWQ43ez9UFEJ5AFsGNHIwk2NoVfcsS2
k6UHSQGfwxWLO7yVmkO1AM2K7TABcEZmWKAII6pJq29qK5p7O8TLbIm1u5KoVMQsj2+/mBI8uyh5
o7XD0riewERaVu0QuLtXaOS9nGouf/JzrZQOC2dSZT2YLZeHypwJIARadA3m+r+H7wb8KQw43bAu
NVBmcYvB08CmcSJGPASv53H0C3DzdBqpqWk9AYz+pazzIPRyYHycMhJXR+Y+fElum2QGEaQV1npg
mBjOEDmZkMY1dQiQ4aJn8C2SU9PtSLGwppKdQMUBgYLBCyFiYXdvattKtOcXdpccEtvf3zM+PYo3
5hzJss3Ts9KMcG3oLeHJz9/7YLIBG8n2Z6AtTqSW3qqBL+2m2DPRBhCAzpyWDO6OT5MRuTlxdIO3
TaLUqjYs7n9UbA3H/OvhopmhXBTnnIpgU9KdjwEojPmuX52Rxck8pEimEgCQvWEOkcvWWBfAzHR5
6dR1k1js1h10HScVp8g4r7CinDO6Z+arraBhMFAKTpletcMYrjrbbujOXKZhlC6g+EV5tRNWS6U/
sUv3hXAw1YN0VCU0nvACstG1GYaL1bi//kxyygyRyfe8AVqU8+rSgL3aeBMY6mxHoXDa7+5rYYoO
VoH/gk8oVvx7poSzncqE7vJXX368kgbmHSYrLNMb95ezuDkU3qZJFY8JZ2VWBAAAChg4WJQRrV/Q
Lik5NYQECQNoggFXxtrc+68WW9kIlUZZMKlnhhCcg5A1Ob+U8x0NwRtL2FrK+lLBjDS72B46enR5
v2N11XfU/Ll4OGzobnq1ZsjZ9G76aV1ZpaeAtJzQ0R77oGGD9FiqJ9CIBkz3gTqggm3mOsd3Vbt/
2IEOIEfgwJGn5R2hy2AGBTVWFeOAcDZCgjhQiBe5Co9McO07a3Ab+fT0Ng2W9KXifTBvn2l61W/X
6Lt91eyPjr9soIral+3wQRvbh3htkgmc1OQNNmo4WBTEIEQGgX8EUXYKcg6CtfxQDBW9xnTWe059
JLQCPQk+mJar+yKKMmByr0WtC/CzIVprLsiegXtbGrDeXQGDSmKdGo7RIHXFKp/CI3hxpu5ZXl/8
lca4gf2RP4D99CD87HzuByv9g6V8Ni7fDPrX9p3xVlqPON3B7ZYP5Qwye9wD++qLHPQzCmmqAd4E
WBM0ki+OKUk2+14iC7W9acs1B2DyqVyzk4DCzSZeCFbTIdhIEhylWRJEW0cmu5Xvfm9MXawDVo58
myPt33gK61keKJaF6cNZ1NfYdRmALvE+VA3j2jr5eMjGo+rXFsjdK0bId7WtHa01wojHPmPd4XJc
811KbMMCmLGKrKQrxjFEf9aHXbs/EmG3gVitWB5H8mT6eIKU4kQgMCQc9T5hKm35BhdVONl+cht0
XajP+/kSTW/++n9cott0bm5yYZDgoOFs4PS4zjp77Ao1SVcbpsVylSJUsRxmvKRNrQlVyBGn6wuj
APj97A2hTPCIYMI7QAyXO/BDl46SpxU/pCD1s36eXcdSJFaRJDRleV+jJt8U0T6AQXWSZtLNoaZF
ansgrPAvQpUOETgqOwkZts/FeUysAQ6S0+ol+Gm7l3peYTkjLmPLhfU+9ULSj8J64H3UGgsqD6XM
C5DM020OTG/S4gq0PYKqdh1p1uBj315XltP114awlILS5w7v47QJHUWDVKEjqJ0+OYWmRRJyNtje
V9zVRABiXxgs869qW8Mv3mxwLuY4QA8dqEdyrDcrwqxsZ28x5YJmi7g0uk4aWzaXaFFUzD71kxpz
Q4/V6fzAxIsbGj1fUDSUlF3bsViWI5M9kXXtEDk4vI/9AgrTPtfPrDU/tBYuOV/uFI6CiPJWoCsi
P/67L8OfcMrB/uMweZ85hXFfAOdsftrEevRR39+4/rO2UqtO0PvUZjCFcfvp0jcIKGVmmy9z9MCS
VvmRsLFxRE0FwyOQBRLEScBHJHdq9Z1lhQWKuf7tnHrpt1aIcaz15cNymdLWFOeVXO1PiKRCukk7
N/qu8ymLJ5ZueOFLD+qNbn1XBUIlIqAHqgFvMO+obyRZHwszWcVeRCyf/2VSKwOq4dNGGMi/eNX4
DVUBex2oZ1qdgP7WchlCp6pyLBwK3gn/ic1P/EW5/+K4dknegtOObm6vuHZE8AZivBLaxVGuEmby
SuBYBd4Znr71pTXeUsQEXwPj2RUJjspcMHsHTgi8LRSljbv10fXhmgGvEl3Cx2CUq2Kqd1bWfJ3n
vLdhe4DHQuoPq4qrtNvBbKbNodZw8vyy9SJPUox5DFew9dK4uiCZTEgoxt/saZKNXQD1tTFlegWH
sro/ENwPES46yV6Et29FIL5KUx9WLJcxqteHb3bH3Mcmhgh2HcOeeA6CBu2gUzYNNYI7zoEQQIB6
KYQScYJINiWpVET7HOjOERj4afzXM13kQ7UTBf7z2ap4vmWz7BbZ6qf7k5Ydz0T3qTEweT8g0wam
9M+3+ccJ10qsPYPf4E9ZpIF248avCk92uY+hJvfhrLrSFrXz4bhrE/i1HV7SOx4opSDNzar3m6T4
JZ5g1fpvVVwIT/X9PiFA3Hn7+wemVJpgaqauhzkNgvNwvYtaexviJuzKCneVpTYk8VFAzWy5P6Ww
2UcWu2laBEl69JawqwesdPDsgY/USE/wa+wmvr/OXTJofcqXAQP5VHBMNcW7CvZfgIwODf9sdwSw
78cd6NeZ1P1vHJMrqaHtvpD0HCXwvKfzu8JBWbKIisc+W0Fj4reH2/M8tRbq5cIxvFkrS6mgS/3V
8k0Jqbf2GixnVhmVYhuoP8gOeiy+tmpVcHfMMRT01joNOFHONxBXt5/2f25ZmCcchx7TzxePNDBA
O1E8NxKIS7ml3Nlv/pesvxUfEMHP4Qy0zvgt5k0cA8t/C/d7P9w8XS8JVQLSkK7zXqddcQ3SFL3Q
gZd/x3yMI1NCdoz/SXFbPj6waDHWgLHK1jKPJ5cZixUFSqQQrQKmcWYEnfuXnMcjLFhtom4VREba
YcsHulVoJ/GrRkS+BbD8JINBjo44A77rT2yY0OsFlpAYQQe+pVoLjOy+PxXTD1JumPHEKdTXiA+Z
wgw7+KDnLosgSrZSgkcoUBO+fP2W27if7tUIUrZ6M7VPmIV10HFyRYYLjPsFgZUd+8ZPTXzrc3hK
8O/3zFgM1kuSfGz0m5QAHO6pXosgAbA1AtMH4Y/W7bKdsfs7K8ai2OFgL/IAxOcc6IHittyUtc00
TqEGrGu8vZp2dGBC1EFjr2la5DXa5e0TyTANVfKjUXLIxuRxwwAzH15sv5fLEc6O3FCsUKijZrKr
LKw7st5xpwdA/FiSlT5Cf+rfS5/ve2Bk/YddbWzlM/KWXDeoIhnuZJ4PVwLkvqwsbxeC9jsRJbH2
Pi/SmoLXrvNKaYkFoxEetDKaqPiisyeGN6hgRphWLVvue6YlUs/f5meJd8k220yn15GXyjVhEW88
bIpKtiHPi0FFu94rgelVGSlaTdFRLZ9TIRWcAqKuMGbZJGlLnM7Vlmn5OL53uUm0Ixuf+GneuYry
RqOH0QGmMumK/XOVIzZ7mFg7o8CJDL9vJF6OZ41PcSJMYR6wSHhNp8P8LwZCFOa08gqVHRH/F7CK
BqThvtZqAKSwvR/yXC6dAE34EJd+1ORDJQIcNvyfu0ZRnsh9NNwL/gvnulkBgy18TGN5QZ6Qr7Pf
k+h2+1N2PVlGx2sD1CuL+NaqSeCf1GMhdLpte7DMe+FxTNxfSHq/Zw7E9CD0pkWqUp7FDF6Nbpnj
gPbHbJBhAsJ6pU1iKIkmzHzgkR65+bDSfrtbDPOHAqrZAXlR7vMNwIFHxGfni38eXVSZk8LCeHj7
BAz2MhBQ3OUnxEnJ0WMFLyPzgMCQqnKGsCDJs7Qz94RZhf23aez4+h28OW+pXQ3Qij4RqQmQezoO
rDjnWJ1JbKyLLjDKSuo6FXysz8qbRNV5q1VQYGJ6udtcy6v0lXcUoEUcCILEf+PrRsLX3SMkM1x/
jB3WiMHdVB2DJjdzNGI/IvYZX/nygJJ1E551mMMvnU36PEvJIj/1ToD5AHqizyeCIwUmdSJgkWA0
q1XihMaBdUhhgxqcqkbZKDNLKh1VIzlYvkTdV4/ARJ3EaE5k41D/5qqpyqaqVBbDOw8nE4v8cpte
h+yvH8yP1esr7gPKaZHf3SE/JuisM1YlUvMIw/uf9AKWLIINASH52P7n1rpwBaAw/ryCTc/NiEIP
B/KrCrMxBlZbWof10cT5UllFrM7CSTDPWnaPLl1KY5SNggDZzT6znZRdtkUeDNIET+wk307goBkH
vBCMcPxj427XlsRjwneJaq/C/wDprXz9N+NuQ/dsmI4EnK6qxfgtatUqrdwruHSLz4mB1HD7oZuW
FnA3nd8Wm2bqXWhlReH4cyCw0oSD3qhEDab/zPZ6Rvz2R/3a0wy/FA+OkJuQQu6uICDSTxraGQcY
KCHSzM7jfX4aZnj07uhZ6dtKfYT1JvW+nbtY6IYRQ2rUSS7EaKiCuu1a1cS0tr09qOPKYEfXw/Uw
3OGG06y9ukNqRTP7ZQYVAIVwFSJOuEN8X+MiDitsg75kYyldbPG/1jpH64RbyytvIQBt9CKs18tI
KoUcJ+Al2wJ4f2geAEd+iImL7WZpyCM9jDG+0LAkwofkDoESCDhX2ooMwAwF7odww7ilck7TImz7
ey8B0RlYX2SOvxbzU6BEE5Z4TT2t8MySVCXoU4C9n8YQLy8R1Ce6jrAx8oInpHfdvBa64EHxC0QR
bzoTH+DGeowiXYzu6RoVePAcJQhJZFvsWs2sjId7DpAVTcBlcKSGYnVEIacwEQ0LlrIX3L94On+b
r/nSjr2OxJ8fZHcDYozHLIGogB7H3hnahF7vXh+k+e0E/kgi/6/DL6LOKTQpBefgctQteUZyD/43
NN3rOLR8xkDoVatI+5/wJdlMgjn+xzqO3aVo7MyBo4FOVQKSreIvfSAEBZF8zQtOtybmSU69oyGf
K8ILDWmzp3ucNXtJZ3qW1/QiLfCv1wHfh71KcAirxwgaY6Fr1UR7R6brlYJQJBeObORw+O8rtdla
Xuejgbit8fZfxqfwjD5P5gtGnxRpjqDq3UL50o9fl+WrGO5zZttILy69pGXzcAT+C56w5s1wzehu
6WQ7p9y4H/jf++1GAzOUvNv0e090FdFRLovocoQ5aEst15Zr9i2sMi9Z2X0ZqfdfNudkJxoV70DF
ffgXGcfJe1hseUvJl+r9fZThXGa05Iupo+oBVzjZ0J0aVVFO5GN8fIuxMS+1GJlYcqqPsJD8Kr3E
v0nl3kyLtfIRBMYhkpCsJR6Ho7rSoYHCMxTr/xwXpBjG87+3UZztr9cpO6U+nUElNKuTLHVyOAkM
srYshtRZqcakUVCJv9XMvnBeEEhQZz8lZvW5K1NXjHd3byGq5o8xgHJDrnWyu5F6avZghqUKp2b4
b8Eo6TtI4g8BdnDhfDxSBzlgfw/6uNRe5hyYyKW+PF5z+A7YzZybtNwaOPKQhXUsPgoGykZ4juL5
wA/HJc92cvkdOFO0WqwAJGGnylA2fwCIEPfWecT8+5xcWReoaKeYqVqzSTDnFjHpPgxJycXNJgob
cMiOFP+GQ+pTHr3iRD2NDxU7F2ZHARMWhHZo7hTfrKOkFFqa5jroEu3FnJaXiE2mCF/SMqoBNJ5n
XL2F/wKZ+jlbUHARj9RR6WPv1hQ6BDkkWk+fbQtyKda/t1jV+9moAYS3Eafb8cPeKuFbyE2zBVKs
dUeCncyxpn8fOMj7w3vlygcumr9E7L//elrp1PX2XPCthYyCopZE/f6ew+hs/NDTB+q0s0779N3n
O0dtYw7GNddDDpxwZ5TceK9senU86xHuv5n/sUCJPVoJpoAu1DbOLBc/pq5UH5tn662dJf8OoZwi
lLhRI+jU2rymfNnqnsBg6gXYsnqD450sjYFaEDzM4jagVknDKou2HOghoNBQ45t/KLtGEn5k4Xld
p2X71iN9IbBF6FWg/vp5exSkBSLLMRbnLucYdB2yi2XS7wA6rJNYOjtck/i0O5n1w6ww223hchVg
Sj7c3Su6GnXoA76QsTa7Z46oQgepqEoC33elH7GzmqIf8382YddRWiPv4CSvqhSbAi9poEOjsOLg
mXKDRYd3Gym8J1rIsuCrJFU9fHZ3dGlaBvWUX5xZS/sbtUtyY1Eb4kXcas1VLZC8RvIy7/DH+PO8
dBlfY752k1mh3q5VV5yWU0qm3j95K99sUsE8bBt3dCiowJjSqaheBcXBFpxGfkLzLM/PLRDDEaTa
8YI8gKMvbTFDoJf9VIs83UgLtWghHLXUFfqSg0pYGuBCAgOk29C/+/BUmT5qPHfYE9CWo/Dk/7hH
bDYePDGnHiwQBOtumzwd+TEj8NdeLdliuXnZiw5OSNQbABH+H1PIMcHLRxC2BfP6/xbzoL0Z2sv4
guoygbf1/7wz4RV/bbPt5Smn0XkzkpeG/tFDssJS+qAjmFF4OjTDkbyfNdWIgtDOLABmaAsfTF5n
Gq7gyf5Eziqj8iOkKctMI2w2Ki/7fjIsQdwAd2JfTM1odC9pyg7zo2ZPDpjYuKwLFQ0zfXr6h1Gq
V5YFqAO5rzqyp7uFjSZ8HDpmBBbqett6Yh2DnQemszzodc64agqvOH4Hwsxj0jGAeVofvp4ozONq
gYprPIFz0KcX/fx3xl0a6siJ0AC248oF9p/+ZKbTspnKgl2Km+9nh6uGLCYSvmVuNdCUIn7D+sGM
QdPSE3fvOE+4R5C11OlEWkyKeFZQ+9KvdzoW8/Q+s4p733GR6skGAskt8kG2u7y4sqHpYqYUr68V
4GSxvRgTAVsXxKy4dkpY4YK16//6NeLVXMxVm/9knNk330ECUCPJPDGz1rnH8DrK4FAcMAUKW5i1
RjN9UBGQHYGVJ4gRaID26l28YuOVH65KoH1Wphj1yBdT5PPeJrvyxFbWWFI4Prwuzeu9Agn55h0e
mHqgzH8rfo1PJPySiPLzAbu3pkJkqy1nCCvcx08bDLrgHX0zN45N/AXBQ4b5+o0BhLnSb3ZQI6H0
R8ZsrXdDJ/o9WN1jd5H1Fkvk+AqPj/e310fEmcjYlbC6Nn31DxtQSOsMqK3fOkH/sc34TbT3EAQ0
L7sZm+yCoKuQlY9tXtwrWIHm9p6jssdetApVeeEHASwlTPXnHBA77dCuZ4r1diuAAHaOjjaIPPhM
0ydShro11W2hoacCBoO/f255XqGvUYxwm2wNwIHFbcYwk7x80Kjy/1PEyzgkeW9x/xbG2ggfle8h
6l7WLkVsGnPQs+HUn33ytNQDdcKNszkhxCmvE6hqvpFVpWrieIUxtLTn+Y2vh4NKfS99xK4Dh9Lj
JWY6HmUSjsadAe/dRy6yaur6Q/AKbvPejVxbEEm1a9QUbW4d61SWHxYWilVhQD+MqQqM81eadaXW
NuV6q7xoT++jyC09SCvBUrESNGbcwen1c232LLzhU90HQa7SftCxSlra/8SSASznHY7JeXtZmL6x
F0Y1Mxx1G/Mg1u+bgkaU0yMRx+8KfwAOko0dHnSmljEj6rCcdUCHqc9jaidgQ/QFYDWjiRQvWs5W
ti1Xg89JSZwQDQzHeSxzON0Fd59BWx6Feyf/MdVgjY4aQCCjbVbX/KuqcntaeHumfHeUncpWiM5n
jNXOfErJV981yLHWmvTGdT9imNanAKJREjoV3i9u2GCUj4DifP5GQSEzOMU3iiPuNzK3ixkQys4F
RfVR4WEFR+ozST1uLBJ5evEVF/Y1uAnwKWp0zH/rTg54Ms0yohcO/TAERp3DFweT5BxbTc/gamlV
p4KvPWQdZO/O5C7Z0ii7ZN9bPAVdl2zJQ3Cxn86khwi6loy4j9K8eV4P98GPOBUtQUvmVZBmYyVY
FmchFr5JV/TZF9+/KbupFjgrM9lH2MPxsbDNs6T130PaPZnduodso9f4MvN5RIOJZ2myoGEnBr3C
4aF66Ytkw/6V+xFIRePcSE6uz6qNJvXdRfu5NSGJmo2tcCGwcjjGMIECf8Q9Zh2p9zd0JOAmSYzM
UIWeuXPyxbriNapbFnbjaZAVn9eFvLFDZIfQZv2oEcAFHcsiUdpuybER4RtvqQtEg7nYvVlUA/tY
yWOCR1TMo6Q8HNXORAywsb+tji+ZJwoKQ6zyY6ayRxsEEA4DEzVulztapdIehBSqccxfBG7yoaHu
cfbwbgJ/oOMl85OrlTMPGJJ1RVIFx8fLRPdjyHkNeF0uz0a7z83dTXXRPoLM+WmDZTRdggQdn6h6
5i6iz2HmpmPXpND0vpxYShSAgOjFDaP8TfZ7UgkVwcLfJopDearsgKfOrJzvQDG76pI5MMsK1Mp0
aw2wSw1iHhGs80CsLVEi0Ft6LDallz28qi0tusw5Ib5s+N+UX7wJQ7RaU9zYboA/1XiKdFArgGPa
L35V07OHea6OB5UQF4uEmPvwqoCqY5F0CEChuIZFFowv9uCHY7i/925uyDmcKpSUVk7kZgxMUKho
aumxLuOY06N+QCN/FRpK6gtAcUdpcoScsZxoimtUAtNgWFivs80Tj7jyFBPQY+6ACtsoKdumqyIg
vV+RnJRTNiiiQP3aoQU9878X0GCg/f8B4qIR40pLhwjRP4aYp7NHGB5JXGCYCBvm9pY5tJHr2Etk
4hUE4KG4uLyv6+B9Vzpj/iUtCkI0Bi9KWlp4jds0T4RtiSJ/T5YHPlICZTI5Srp0aqZJFnUVLVeG
VnCWk5TFKGyv+ss7UIBfR9Kq8rEGwhyiSBqsJrvmH1Mhv6lgaxu224MtHbiVsplRCHXeL1MCsMz/
4WJvcIlmG5NnttiLJOuomSyB3lDBlvMklGs8vpLEmbmYsE+e86rbA/+WsFOu0pXzkM2soygUwR5b
OvxNqE/QxG0ScD6q7w4Y4SQp+xF5CuKNh1DT8PYwwYEdf2Z8ftIVw367rMFsefCCQpzTPzrTLiHu
w05t/YhWg/A1aIgiMuHFssO3rUdlt5f4rpUNqEmq73tY+fanpR0OVBZoIsYTKZ0N/JVEHhC0atIo
gXzxlpyRumqAFvcpx0jyu+Hr467Kakk9ulsCMgVYnK8sO32xIOZ1umNu5sSltaN2oQrSuYt7mk+F
do7jt2iJAmrSk4UYXhajTu6+yjqsq+2gmjDf7o/GrY/g6z0wzdFU14kpszC1LxY1iNBttM+BOC3C
KGS1Ulv2nDVQKkbH3aI/t9oJILxUxk/mD6hUZO914yY2Iuu3xZvZx3Zcn9XLkQN3pV5G09fuhi4H
Q0LTESjqfgFkq/1K2a3/kqkARoPXi/j5uIakf8LPw4fMXdW8nC4R+KVMyi9CA0QhXqZiavXeq694
UfuWhIl2tzys4QTeWuolurpiyEiHdAm9tGITjmXO3nUPqD3HVJF8TWzscBvNiz5Z7f2Yk0AdZsKv
hU2r7ejRJIMV5dIdwdfiE7VeCv7CKIz5AcKKxbLGzE4M8yXR345DANRWh+VZ0aYvyW5njc1Ik3q7
aFZ8j0rLYdWNZwbMhertTFCjPUUh7jufErpyh3Zkq4n+ft/CIwJeLkUFYVPw2wlFVhlGtYhtId1j
69gtvPdLCYCfxxMFa6+Nl7xItULgrHw+pv8SP7rKuvQBwFWv9ciKbMTfYMZZJpZU2pqmtvXHLf9/
Owg08WkBWarPC9pzAHCe7TktxlR4OUOhVuMd9D3nhoI7H5MrSc8ToW52EJPjyxD8BmLIDNDOKuc7
k/DpK10vLhjdsAq5WFhM4ab4lfLXqSba0oZU0Dy1smgpbDC2zSn9wI1B/OD0bDb/zbm786CNXKt4
/AaHRYlaf5PtnZyZDJ+aSvzEdMUfh1FlMaWzqbI6Ni+NaB67KfeIb4OvYV8RhUq/+NolglMIOmA/
bkdQ4jDGLC6fKxxHr366eSz1oIdehvpQzI6F3DXWk3RKuZUNXnPUQ3ssNqOAqMssby4zCngfdnju
oLLtBUJCyx6Sz+dq35edZoJeu7wZIy8lyadtIR1wCJs+xtk/6s6SOMhBw9mCBR3yTYV2mr5sLc/s
NgCpzmsjbo/88ANAh6J0HEG2sB6EqJgQK2J1F03JO/D0QDmPFM8h6sKsin9xLH2Y3kEsYS+P1MC5
Mcb4NLyuOHzKI10faZ5O37j49h5o6nGqn949ZBVuWvSUCozailZ5RKdTjWGuXSDUCe8eMCkHv6lL
71kRZF8407cLVa0Fy6GccRC2BMpLxM9IpBzYZt9eDxq6YXXlHA3Sg1PGgqBF+hzx6cJzl1Qs65x9
kDErUgNTnPaqiv07uv71wmg0G7ynWFNZkCf0X/P7Qu+rymUnRXtOI+P3aBLQ+IZKhHa8iPVzLVGU
cL/EOTvxd6/vX/64CamdZ3t+eFy+/FuQu7vCKMq7GHP3kYff0HHAaskvj47a6lrVH4WfXUQA2IOp
vDm+U6k2Ia5EfwO7pVfKB0beLLRTcmVS0s3T6PXhOiFvhakiEyj6tRyfUZFF6/ayoEECLCVmilNL
IHzsZmqygiKYvob5VzxvAi97Wvpz6rKyP8wQNpEbuz9bntf7Rhw42zrwEcxrkF5U/lYj8/OUR3mh
KXbjT7S9wRM7RIDTaRkrXX5jgDGkbtgKtwbMKnUeYXt4KaFWEkF8JSxTU1hIVkJ/n01gm7qZ+sFU
YOnEhMeRWVbpTUHx7SOfBU2+lKfdE2XCUkejguUdrWUJm96PeYgldVAgkM3g0EKYRpbjwCISFRFG
86kMk7uHIKURt7HnscW3ViYc7H8liOGMKznn3zZ3ZsiOGZdgOUoztXsw9eNZbKOnOHKp7bt/gd5A
VaKP3tvHBpUIpcsLK/Z+3hjNZqSS2UYvdc8f2oEgEUJ2TPj1cO5t4oLvei2kiOU7z2yhngsXWfAW
urFc3YTA4fwtMTsqkAq259QNJV+nLfXZ8afcHrckIh3xxEt3wk3jkLaocvndpOmYniTve4eQRZSF
od+pIS8kVL3N7KOMdnyRIAvM0yURvvO2F/dkDKP5KVYOClvPG1N7uAekAQW3oGeAPGA7PLU14lYo
sMEBcZQPrenrWZEHHEcpQogHt8gyOAjDV59iLonIGZrE/hcRTaUi7Vn94gHtElcHQJe9KO/fDXI7
A1GwpLuEiupH07yPU4E/txQisId1MNIQnxg5CQWtmHK1uO/3p8Bpr6jzbafsUQkxtU+jM/PfVyjK
G84CXqsXi1OoKjSpztzQsfQKmU2yZudeItcHE9NeW5RZlgUauNU9pj1PKwcqM3sjnMdS0sBU0xkL
X1dxduMvW9KSPv9HHNJNWmb9b3c7W+tSZK9OtjlwPOWg58pByXw9fkru0qhvPTm9H/BcqijrEPfT
Lsb+srJrksKEzOk7T8GLWz+4cUXlUo6T+XTwfAsPNCSWmgsaSH6hLLls/WEFW05peYbxCKQoi6NJ
LZU7V8eOZHY8GWRMkA7PtTJyJRigX3Hh3M3+OEiqV+TgNPj0mbJTVsbXBnh9yW5ljMlgLZZ8l+z0
SRd1EtH9xa2XHoeDhGfWqsBFurw2Uk3LMFkPdmosdqiHlBEnu68vguBEWHgAUT89VcPsycTE75lv
Wm4M51ghdzDaaQqXWLzLMsIlnKRI3O9PqBmma0KnFZrapzojHF0mn+yacOqS2BkEXmxkpDyDDmBh
RPzlRityvPOEksMxQLbtJzB/iQb3iyQ/1LCLYwQexMekUjOOYEUSwiloG9wru3BeP7YkmoROvmgp
SUtHoOFeyRBYzCSdTwxUXaZv3sjtYAY1qju4XiErKZhBELsLn1YXV+oXVNRq9TRzTSWk7+OGL2IR
XCyGpkbScQ4ybaxff7yAd2V+LJq89iV94h6jRMu7tRpcRqS6e6qSbEVIgPx/P8z/tE6czakzmZiF
9BeIPBVPVjBVxgRT22vmwL7oDk/J1GIQ2OZUlyFWJBDneJb1e0aBrHtY+qRpPiDyLwGNwIPO4Zzm
6kKsTUYTc+8NMCHUsbNPRS6SKpUXUsSYMbLp66t9RHd0GqtxRHipndLivdYTRpRObR9UR0zmF7VT
ukfC/mGFTLDBL8lmWM0QX3BBbfu6D8YWKEWeW0vQ1UHLnqNQmVXeDoQqcguwtzVt2/w0OprrOlEK
TrZRP7B2zxfOEzDPPa5joy8amZksgn80YR45jZhAP1d1ULWUXOdTpZW67byBX4MNbwc6+tKR66Mx
Du922rXKvzylulbe1U6dgP4uVQe+JmPnUnbFGSfQl/oint4ovzKCH42iFKFWKJ4zlQLnzsCXop+W
guDTdPpN9i8kuY3qdXrV7Xjz9tGXq/h1cMsUFExhNZnjK0c8uw0qb6onrSo1UDZZf+W8brwEHuCj
yOnqfADRDC6PXhO2IvMcDrOrE4dNehIkYtLPzZcfAdNikyMoC+nVtxO/2m5YedphfXAXMSRr9tRn
oKyCIs8jFaAI+n4xd8XHYC17Ygd4mpnhV0PZg2DASdJdHOlO7ZkHYn0sgECgIL60+yAASLR37l6j
ncLX9bOBLSNR+RwKe3RTFY42y1Qofl5VtedkJb/s/qab1qnoVeVpUvkuat5EsguNI/q8oUuoRFUM
9i4eY7TuYDmoGNe/aXzPfJHLRxkhfywrShiMk4Yxe+hboDu8cJIcNQ/MV8WA3bbsatvOcDiNxoSL
9lq/G3ffaJEFG5E+Cu88jfTJt6m4+poVFGdOzw/pkE39E2VqGaaTDV+ImEWSKGMu7g/LRl2Xm6Xr
DoS8FkwtAaztXt0L332aHDXglh21HBPQowvs3lkA5uaYQXMck8OAmnwGTE8WZW2iTqbQ/YUfSLBe
NOTt5g8P1n0iAmGq3u7ugfMK3CU0oUPZWRrwb2iDbKegcXR8XYsXQbDsnI4eHdgO0b/jMTYOq+D5
49FGbI33Y8dU8OHgVuP6jc7dPzKjncs0ZZJ9yzmaXIqe8zvZ5YqeNkKMXLi1VhxuUOSJ0NEZ+DJP
ZSexKJRZu77S1GHbauptdzXeymorMTr6SQtASa1cH5RKvkA3to3YK8y5JWo4urwTbrmXhaLWjCWu
sphnwG/q9ladsIUP1koSR5sMqKVNyOkV3MKPCcOvGu/FdL4p7vEGk4R+ARqho6UOAO9ocwRnR2Fn
w/UmoUlCmRBpYy8Z/1S48MtzMoh25rxX65g6mwPmcky1Ph7+8JXWFB+ZdcdtxgU26sFOkT5rWETA
Tztf7AO0J7zXFZ+BWm9TbYJBJUfiJXcKh1CuBImlq0zOjJAhCcz1eSwSN/I4r3DTWNyZgjrW9OMW
BJlSksaHfmnIGFMYJGMZBpt4+48XOLgzxgXw5XNnwQ3roKcvKODOg1EhcsT/P1mK506UfqXA8Z6Q
eHosnwYYooMZoRFWQUFwevbEA7u1JxV1RzH+5Mo3fOHMkB3uNhxb6OZaB0SnjqEXorO9YnvEYD3R
t/nheC2ITJLb+bA9VSHMHeh5njcWJUkzMdq/RpaiOha4q3imDLH+EY9ORbotXQCkf8KiOnJZ7YmI
a7JSmwgaGo2oWrqzHeon2DwuMI5sErc5nVx2DmX81QUVxa6s8K6VYj/s0WDT4RiA4vNKj4i7anue
GcrDRWyH3ui3LUTzp7XlLvLpR4GMjbbY6IHjTyfrKT5X09ln3SFEqXTwi+BzK/vsNf6EZ86YqCtd
DWMxc+TnMb3nR14ukRfEPjIbgkkQ/d/8uiJCPhJatp+Uu5HtyWGs5CByuVgKwYq/WfZv0WVFyQSM
eK2N+KjXs1PRk1ZSCaunlJZglz94DaNKW75U3YhMNSHcWM0IMb28hIEogE+tmUButskl/rOBDOHq
9EQBI6MG1NRSGYKBW2v1+VvrEDDCsX3TJ7V/hUp2ZYJwNMb09UjP3fo/8ef29emMvz4hn1y1Eo5p
rm31NKznZHLs+RBjQXZIoGHlnd6+xEUcutucI03AE+hfViX3ZtKoKY+k8unI6yqzPZe1EIkQ3ou+
tELqxR+CCyAW8Lxgf1V/nMa8igTYAqijC3RO4KXWmUszy+4We6AQxaBqZxhAMHytMfzVcdFhbhLv
RyVG8GsSQKUykPan6eJaTGUIcRKx8DVyF8dDcp3g6g+zg3zHclJ3uw1ejfBeKp96Z9cJgnzR6RFJ
PBGEB71ZQrmjjfWbPsD9N7rDMhM2iEJLcj408h1/+WCdVE983SxIkdgGRR9cHQaivsq7h1VBGUqp
ReeAqLzorOZaFKmOA4FzdMjJt7uHbKZ9eChRcQuNTx6OnyhZqkChzU8eVkB6JjZBC+ayDBk21wxV
uZyQSkZR3D+YweOCXkCWT7BLtVAAOkgmls3jatDtbHTXdJDdNq0h6ZDED0NnHCfIMB+TpCXOdIZJ
6qqJioKCiDwIjZnI6s4FpwFBk/2SJ6E17y/yCJCzzEdkxWyy1Yy5PmxmYQUCKZKZJjLZq1uzkNtY
S+VHH9wXrhPorWkPCMVGUfFO1bS7vOGtQmq2iuOkCuLtzYz4wfssY4rM8v+fvukTMnNNLl5ihHRD
jHvu9cxOpcvHyYEMlQeehFrzlcSHQZXiZIly6baNP0PDZymOgs9aYUsk5hGdMZ5atYKn1TUSBMPO
Vrsd+fVMEoKcb2eQgF77LpeyUBt5KIphwDHtNXbTOi/am/P00XJyYiaAfaTmbc3bMAw0JwSCtgiV
7BzB/YOhO8WHQFzKXcvgxD3uM+JFqrc4uRJhOxlBJs4s+IwDi5zeqTUa5ltsLEgHIZgFAUV77OfE
OZfbpKl09bKjt+3B2G/CiGfKn5DJnmFfYyJB9Thdlhrdr37rrnhMhGQj/cyEMsVj/pRGzU+ZNa8i
2Z7LLCx29tgGK5Dqu/DJYyueCVNzBbTCemS4vYNmf91BeS87LogVjlJYkxEBJhe/gCGzrj0ypAx8
WyZ6Feh+kzbumEjUNkEoDnDXiAl9900lwEkJw3LWvV2BzDE9JBzl6lx9CzDXLlmQFtb/T1KiBsvw
78IGBMKtJGsGABBM6M6/StUQD4ew0M0BwSxz0Y7hDtbpDIBC+mUj6ESJ7fiJpzjqnfTpfkwy+5OT
IrXsoM/E3KSSdBA8UKckXWUjDPObsOSyUYExcfJ00zY9kXMG1P8Fd1FlsGO3V+8CHFMXWK5LE9mb
gNblYoGTbMVCvSmQ8mIFZEOmQsewt3fH6ftty/OqFeIFWLRq83OZuCC/fviZOkfGiOJ0dwbmyCiI
V/PuyEAmaUgzxTovboivD9e8vtMvCy5QHo7TTHoB9SJDMQ51Lfs2N/40CtIYxofnsKWSsQAPIufE
SN9O65uz94OzA/BrDzwqXvB4w8bU2M1CS62uL4umE8kJePABBgRt7A20WUuvyOa2wfXhefP88Qjw
csLdDjRwBtUZNvGVZM8j3aQkgFerdweWfwGT/T1N7loMLyYQFi3SnxN81jICA+DtMpsRj86UZDK3
pywsuIuOYjLmkbMiw1tr1aeLmVv7DdpT/qnefXvsGhHTEoULKXfAWlisZO93kVP39twx88Hbn+uO
trT6TNeYHxVAm/HfKsLWs6ROo7qYCbHlWOGKRNj47Lb04CiZxXrLS2gCkuwkhVdtQ6PhuzcK+kn2
SkccMMeW42n3XCxIFHlq/z484q2NcUZVPiaHjRtj3qDnolr91eDnTun1NAM72fJI/Seb4bKljnyZ
5L6KvVQ85UVT4EgFiJ3ZnX/+rXls/LKmfu1wZJZDWyTPlA+dQXKgDZ/9tuxV92AkQoShaQgiuCck
0acAq/ZZgFcfw1y2Wk5CifPs3vc9zG2TZx+Hh64DzU+VwtW0pkEb1IsDzMGyOkeLpd1MlfsJ88p3
gOmpCc82W2NkXNkurJawYPTE4SOa/0QBFgsS85zwn7LHadQ2xJuGlhQcrZgLHUSkxfiHlHd9J9wA
PSSj7/MUftvDUQfd8haz5k/dNE7ZDgZuKZ2uQEmkvsrcCEOnAIjcK2QMjSr+U5xI+Ly23oaqIlct
R1C2rvcXLPiLShhcdSqu0UZ/p6twX3mmNPbTPdOrwBS8bA4OYn3XBwUrFm499ImWMpjdRvvIEPT+
5L77SH1uu0x0HquSGczAzZgyYk+2+Cgb+iPSDJXpNYOmW/S+ExMRor1d3Jk/YJrS1XO3VQ8v7hyF
nGE3z51UlVsYApeArD3iiRb0i1n9aNAwE01VWqNzAtPUSG5zEw9YhGfrQQH5Ba8gxkYl0yH+YZgw
sUApENQFDuPY181nSB3KjimZXRD0rrvWKZAXmpLMpm7K/DLTutFVww7/FZBCvnXVDmQ0R9/myv3+
TPeueQ3wr92HhlvNKrFKjagoicRhsxhkvl3++jR3V/GDqy9cRP0uacfSc1WA1f82Oo8C0sbsxQu0
WSte9KYbLGKvIuJUgruvIt5D3eLE2RYdY21bLeBcC+tJngAIBAjko6vpc7e2AHxwRZ4hZmjPWvPI
T1X1gjc/ed5MM1wamzHFzTzmd61d/cZnFNftjhqoAgW2IpT2EkvO+N7+Q9xhW5N6OWPtCVbS3egy
vu476qrzQ2KiVzup+IAwLflc0VONuNC6FaKYgCzumsp+h9ECmODnAqlB2W6eDwSdBjvTOCXZ6pP/
cSU0TE5XHABXax4jy1PLWnUoKGhGuwRT3UoYjQKEI4rW/UyvS4tPOzjA3b16Dy7yQcYO2GCmwdje
l3og2BPTdCiHkONrIFsqcPIW0G/HxOBKTynnpcj0dmYUz/Q6QZ7DUcbk0lOqQbQJzCkPdXoBhP/e
381hMTwtzKBDXBRaC7NSxiCfuCFjA1pGRjoAf7XIB3hHNXJnGQhAOl9hUOIx96YVRMLuzJlvFYv9
xJgWvc1v7xpEAGPfNaj0kvfafnWiFlCEFa7TL52d3yyEAQjycW1dsP4+1zFtScdv7DXgeKsEc1e6
b4Xy9/ULySwhSoSAOnZJnbelOXzT3kP7sUXXEhXCoRKueV+5cum35FhnUKbfLbLeXD6Cioc+90H+
p/gPCGJz4b2kdmZW3+5aBTEGHH4FZcsMryudmrD96knYy3nNbjktHyVhzGcShD1wolmVB2JmJPjP
YYfYXbmHBa4YycaGhDAFRlpENJ2BME0O5lHKXkFCIVjEPDOWUBx3H2O4XEr1HUrKap2CxJS0wNy4
S4RM5Ynzyn/8OwHHn9vSpx7wTVYg+puzM2D63xKiMcO64PQ2fYfNdZPOn8Jhe58K11skuUlZUUK8
RAlUX2/JEQ96euTc8xIcuZb5tZXQ0dqmyhnChQbQ/2vsMi0Zj9bI8+5TMcvTK13E8RBD+e2nCjTG
dhdTKm8+Mkv01AfBaSQFzWc4x0J7n8KBZWGX1xsq/w9KjeaIE7KRHTH+zPReLPrZawakRen8xJUY
N9QhZwKQ0aW17d2gHR0BRkwVlhRWeu1GswQnF09TQPnhjOeNb77uTSbzYkpV5HUeDDdqzn2KA966
l7A1O9mqv0jjk/5/2brcYqVMSu6AdFIJJ4/8QFHQGZa79vKJrtPVBhGTsOmdGIKLbmmW7kT5pkrS
girObKRpbTSWMyQdrJ+S9ZGUBkgR2gS2+l616XJPzE1qUJxoZNq9Klz55F+jnhvbD4y+Om20F+5/
Gu0XzcBCQCsi4qNee2QZGXlC2hQuR7t+OrZlCGMcL+IcQPyZyfzrEEqqxwjovnYn8Iw/ZutjWKO6
+4aNLfMtkaFFPLgW3+bzfq1bHdVnOYN6zowIdMchAyUUL1EXj4/rTThjmcLBqXO6iiM5fxmS0UIy
R5mbtyhRhJfONdprFfzJODeXXkvZgNGG14LlcLa/HzAzhCGrkVmMjVEcZDyucZtrxp0cLaCLjvJR
W0pB3zK6waKuTRIDJ2cA9AU09TH0d7FvKeOMy9rT/8pXNktXWSEym7gLpQKxPi3ldfu7MthkEmzI
Arhg+UCquCyHErxTnBhxiFdTO/K997TQ81sYxY5rMSqooMp5nF91A1cINMRB0xlZYk8UL8rXUjwj
9/yfQVBEEGR7PXGok78JVIfJx96+CXtXg0ip14o9bsXEd4FVGPlYNt5l6T2lch8ELWj5+Qahv7jP
MyJYwLulUSG9iX3qUA2gK6AIYwXQmW5wixXPOsdKVf8r1Hb5bvIDUajh4ou1vPGVUipx8IcPfz4L
Sw8FHxd59spTyw+MZDpSab9eD+CVdnfkT6YWgdY0zm1LhTTQ9Zlea5EPxCFj3JHu8XcVsvtLXkgd
wvSh7Xmz2GPr8GoVnChjIeEUo4D9TzmhvOwZNIHxslHapxODUuCjnzdRjtM7Bh3P88Dd9HjLzxlG
GB9EIp5qaOWWA94+JLO/NRHcLF+jzYfm5jTfVJMTY9iz4A4538XCPpueIO8ICNYeeDMvX/dxbLrL
ikc5Zcyj2mOvHE/JsZJ0/FxSjVAxsj9ydOEvFuFdSxySH+C/bv0JtCIyCANIvp6mLeHNu3nmkLwz
a6ceBX3O5fQAF32H4paLEI/P4Oe+xNQxVlFFPfCft5tDk1wYltjq6RDwZv+Y76cOSck/ZRvgnzVI
00AvqFwR6UPQewTIi7jjzWriB8NRimMozPIQCdMGmzBhHdarl7tR4Uq4yNgNf6H5n7qPecC2Qhs1
BIuNYc1asKG3zjXmPIdWVAdkmXcY/q7KNEjMQf5ZrYauHoQr3sWYlkxJmxRxxClol/TtYdoV7Kh1
D7Xfe8Lg8pEIeZDDnPGlSL7HFBNVlS+Jk72ge6xvfhyStEgsoP1dpQmgC/OrjmrKz7nx/qWu7+TX
qjT/qfbLz/9Xb8vFjf/zuczmR3qmczCz8nm0kjmjleBtthrM6T5Yzf0Ep++nRmsbX49cs4lP3DLE
U5LrJAc7oYoy9/+6C2m6px3Y10BUEOF6jK+oM7LjT6r4PUcGRcnXcoy+Wor5T3Eq81uKVxGVOXTA
IE8uhPCYqRs/LJgNVaAVx/NZi1FNeQpIFFNgzj5m0QzSCahuiV+WvuVa5/es7K55aym8D7D8i/r6
/VRqEdpuiTzAO03Li3ny7UjuVhA4Ga2EZl773aCtyhqE6mKRaARdCISBI97m7ZC3uYDtD6WO/SJf
MM2wAozxidea+aO4f8mnCOumpPzPwjjNIxd7D5Uqvxg5LRw2WGX6etOsEM4MxHTkZvBjmVgixg9s
whcsONHwhC/59AtEHHjBiAug81Q51YVHdRtb1z4li66NvyqhI8xDvSAoFGFMZt9XvDJXMbLQ+Y6L
YK1/tHEFndNe7aY21T2XFE1NQIeIKQJvjiATN2MkwebLoWs+G3FvHkaSLABCABMs62Cx7eBbo3Vh
djnleGxHrs0p4O6rXADDUovYF+JBfflrChblbNDm8VVljV/41iCD8y07nFEt/TSgzLDlVOoxPen/
exb2Yw7r23C+63wwuLGqj8TVhrgKFUx9TFeTuo+6nJpj+UvGNVFAqopiCDEG2LE/TNw2/OvyboTG
gZNvurp22WiiZJrpu+moz3LutPcPPoBHbTiwgfqh2BM3BWvDlrXyEzqlgoALv2I8BRcvFcLnUj23
tCYw4YOxYIm8taB+clC2ZtBT0mF/hSe6FjLIVPlbnHsrUO6kE48WOYmI+Exrp5xHENWReKajekGw
jo5W0xi4lQPbHJvuvrpSIjXUlMsjJ9JD/7tWGQDFsZ4cNTMeT428t4sJ0925bB0DZDois33E1Q16
jqP5oi0GOIBX/hs2jvlvhA+UYviL++IfG1ADwZ7s43gHSyeFq0Nx8+Qf9S8d4scDcyjbDsnQMqYe
dCbc0jktDBYIO9R2OkxB7tjYI7u28Mgt40JTjXIeg5qdvqaFNcygwlwOhwfbL8exqB44vHwHkikT
EiCG2fdWDvMqJV3I8Vv/JY6PhIyuBpCxvH6jHrFwpepdnIynz0HVHAdfLktp9R1TFcRj3Ih6qmep
RMoSCMKzMru8IKssUv/Y5MfcK2bTcutE0aa4ad/Iya0yxaakDs7cF3W1VqmCX+XKBodhat/BwL4+
xYnHGc4/HyiRnMdv/z292hUOAQc1CYzE811ysatueHUFE7iNZCkWs/scqxq0bGZOKUlM+P8sWgvW
HmgeuWIxXrrdkB8x6zmaz/13TVUgzH77KhFKK2YeQRSP9J7yKT+kzav+zagBjq/dXo/Ei6uwpcT1
5V1vuUKsC79EzwxXhRtF+kQ99QmdjCF2m9XzDyIUZeyd0kxA60GbwaISE1rTlN1EVx70+QQExudI
z/qOoYmDWfeWI/J+i1z45Iz0ciXVbAynGLl/lg1e7iWs6/n/27tXM1OQ/8oY5fdl+XoXbBPSVFv9
P2vdiVkqmGkKfegu3lFfGl4kTPaM409NQQ5/P505zjT4l1sBEePMgIk6cLk2+J8aLm5SnIijerB7
plY9v2DyXtHUbJ7PdS/wl25CbFe8XApYyGidxckHkjy5oquufIrISMWRtAvzcbC42Ki+SJL7T5On
a+Wbw1SY3wCuQA/c0+UElIzm5iAaGfNyqZF5A3o6QiTgLZnM4Pl6wqRzFMuCa+4dsF2vbW3flyiA
gNpJ/JuJSqSOGgZd3nEDxqPplF0tLCcOvhJDQLJPVuqmt0Ti1K6NzPLwJxstAUrT2TUM3e3KhSEH
pUiDUX0gg2TGhIbrKZUk+SKEz37J6n6o3fwARljMFzQb220H7eaZ04xwDX3cuORh7bxysEMirlt0
YrjJcM6y9EQC1CQyDdCLtr9vanKJuRNemqQ8ceGYOpm16BAj6+pbuSFrQsBFjJFwXqwG3MvdU7JK
SQfpjXzH4yi0gU45fIjlJ3yRgVL9Nx6D3mFpqrrpAcxF6pEaJ+zlzYnCscod78j8UC/pFUVqy8oY
A4iIospOjZuXWVNlTQydkz88uIyVCaWHAjJAGP8S6jXuGis/ZptKqi+UT6r94T4fPbbWBffGtape
YWBC+BhH3hua9//TLCvMkvNqLR1kQa9Ac8MKL8TOJ3HCEBWNqGNl/UwZVz9TKrCSvhm4gaQhV4hO
yFSq2RqxWv2onQ7Agy593bT6P1qHaPULGW6aqtiYsEpoPawTvDKytJKVnZHhHzO6Cdh5XyxAztyo
Iuet7/+wFNlGf8vhalOfYin5ki9cbqWybJZtoc4JDP4AYjiL9oj6CMpHK7o5twkdn/BF6TUh/Ebe
JOWxABpDVOEJvNN9ugpJE4O8SlEQqOqZSou9A1cO4/tjMdgxpN2crqKiPiyy64Zoz8YA2pDAbwFb
BcMlxYOXYDvIwpKxgdOKQz92WgTHyxVofL9KSQpXBIaifjWfcyC6zjNrtd2F0x99wVdvmr9V+Eoj
zoQL5kQx7z+4CTihjFljBfK1FrCsP4Na1uZ7tYt1FsXnvae1TLU2s8FpodejKAlBmkDfpzwVoVr8
8IF2q0tFgvPl51qgJQ+PbnexqP83N04xGXbkEQUMzgWTqo49Eivd2ReFzwB1VRoiDvdDa/TN02+O
FzDD9/CXIs2MN8usDouSXmhu7h3MfVZI2Ves5imPt5JgxRAz0u1wKmE/sYwwbroE2ux1SKYC5dmv
ZF+pWbmD5fAvJWDoEeYJ50XsxzD0lxBcuVzjeehDV1ryLb2DypStgQ/y52MXoW58/GUrOIRMITlo
nqj8X/UJXsWZHPafzz3TTCMa1olgCX1huMuAvuaL5ZSXxtC78vL2yflprTL7Loew1eiCOxAtGIxi
shxw9w7U2Yy/3HMue3EgTO54NsTMf2sdvpbCIuWl3O0ivSZNTSGoUKuHT1jLhZWVKXbsmsOzw1jV
GeqdQmFrRcYq/Ojmm8EC+Q3K5CoGdFw3r4ePwh3NmNZjlpAI+sq/dCz7VP33oSH1fYZxDLSOLFMr
umcQxx3lexdwN65/FCqC459OjYQolK6ETTOlQ9tpkLd4jBWjtRW1GznkzwenMiGzo7eX0dRdOt12
p+fyjfPqzhTGpdSN3/XR1A9w8M1O4KDvYlAixJtcDFobUBQuyn87MdQ1OSNkO2bCfnSgkk1HMKo2
HLloyUrLmMh/sKoZIJ925+MXcjk0tPdDxK2nuqBNtGEbKf8x/Bp4oNvrVaxeXkWK7UzQO5mevwF1
EVY187bIkopobCuO4ztptrJPhJlSVEjKBYCQJUUd4kr1yOqaytC1p+HuoWjOByFBN8EDwqtQOhOu
ViVql3X5oeLCFWvcFUtzSsvKAUqt7LfWED9C2AeERqCkqKrRXcugNfNbISNPqs4BoCWDuiSYEavB
JnW+IH2+4xJ12OhO3yHOza7bNd/dZ8pM55buW9cQ+2ZOEMAgSYfELk/BQpRsvOnR9Ym6UhzoZ1zV
NEnyUQ0mmswhx426e4SMukFlQ8islstwqza3Dw32Z2orgcC3nLgb5Cb+3H+8eh+LCrWlGyFSZIPy
3BSsSc6VHjBdIUtiGrjKziLdQU+gpKAxkJrgKZ65lFSf2SsacZ/7vnIl+3NjT5WYWt6RyXQnjnFQ
n57zPCPMdWN0iiwdib/T1m8KrckpU3IBsJnikxKaX7ulVvjtpQ/wiH9d5OLOmN0FowPcdRa5jafR
gBHMfidakvTY3dNlCVkR1R//JVwnuNEfEi/8xWnav58Zjems7yx9dzCxbxwDC9nA76jmgjHbIJd9
JDGrToXr5IGAWOxIpRnfrlQ/XfthrwpHmWDPuvSPZC7SSDXYR+7vSf2oAc4a1DqZG4TKMVdpCAG5
lKOS27h7XdBGh8FHZxxj6AMMaNsgTq61LRgaMXvcAjVm/dtfAUFNe3PYV0j/MWHEY8ACtmM91obP
TZDpkcVuw3F1gfDhHDdSdFFLe78+d6ylNea4on46EBOc6imOlv+2fYz2FdqWWSd95LoGcDle4msi
+8E8nn82bXG5oLswo5sd9l/qGn1SKwayVSef7HM5sLrh5O4dBJfw2rpEP4shhJ9oRzXdi9fyEd2Q
IbYeEyerOWANR1/aDS0Pyn6adYdc1ksGhpUVw4ZOPqItxsDWITPFvY0L+q8HvnBSxIaNJuvp7QNG
KH4yJyeF5kd8wuf5Zbvftv6nk36XRyEkNx1wrfQ7w0iNEMptxZevFczWVJbgmtcBjFTU/eT5MO/m
Y73dH2pmPhjj4pJydc/7Py8E1JUKVcPNVjzZcDT4U/bPgGcfv00rMH1UdE64d5m+CZH4T98gI+ge
HBN9XVvCpgeQues+XJLiKgRnkbwsjbs5WwndDG7eqkf5WdPUJwkydEIHO9M6bo1AazC0eiA2M0fS
ubq+fDZRseBgfK8TwXFrxUEMqm2s1ZGL12cOTjcDIA4JlrD5/inTovIkctNRuYObFVVg5nNaua4o
mnBBxxn2E0cNkFAlUkvVCaIAuif5mRZ3QXCOtc3hKsCcC21VzNY9tazIkp0IMI1B/8TpsFR/I12+
POm9MLpHaxqmdV4NVSYtHHjDULwU3SkWl7ZiDQOLzZw9wgONo6WmHhUZVLeDaLKc9KyKLWDWt6st
82WYcYnK16wuh342GLkIqH9U+6oc6m9AQdhFFwE6EUua10mANyYPn24i0RA/NfMwvcTEqCyt+0I+
hzlIaOq1xLMCs3OXab36qWn9I1hmflI2oLtMJWm9xUuAboaNIyvBEPIZ4lScxcgI7ExyVMRrptZi
+/upDmxLasWRju77d4h3qAykbKXaASNqwQVLRYfLl3tr9xSd30LGiqIpkf9auvE32xlTqK1ZGXfI
UKvXAf21PF6jm5GnsWkvz7oQZOcp8XqZMEIXeo3iBQxmP9MBCSLhNRNt0T7CH9MuM5wrGftXnzgq
RDRMybwbWYhTli7nfW9d4/+CzN9uLId5LqduC/jsJBHJ4AXUFW39UDLfLnGB1O0p4lnbD7QMK+lM
iBy9+JPFjjD35Sh3TV+hVoWLkwf+SKToeWvJq3CWLP47tCFyDZdKPorC5hkzBCejtIn6QxoINNJK
5evW3ACt8SveFt1IATFnA02N13/WFJSWzudWAjZWCwPqH9pGThmCY40+u5qBzOdpitxvJuetzM30
a2Ecl6jgw8DFepirTxgGx4igUcEli/wUcsRFNjY5iMHWh+PcGfLDlBCT8uSDCJojySwK3q5z4Ex6
Jtzc93nyqpbK4r4YY0wjYjGJXmv3C83LWyoMKZot0m5uVS2DS8hIrjaAH9y4cD2J2DhpWME15tZO
NwYPXNHN0PIgxB1WPWpbwlCXW5F3vxx04PsLLH1BEN62xdNypok9lbJmxLf8H4gAiJxmObgnvN0s
GMB9JoZGU+xV7Wx8HQO2bYa8FA8sYxwQk6mj/SDvDZ3pwn+2gApr6FLoxeJbosrZZRwwCG2zMJoL
Hvg8QS52vm1c8isCZh50AoYP76FjBBgs4LcLJGpG9w/VHPMN/2/mo8R1JP25RI7nfc9RNLhg05X8
YSkkDx66zL+gGt8fDjbwub9XNcKPGlZR0CGkga8vrK4JAbIbdN38GvxvehnBlq+bjpmrj72U2edq
Fiw6u7g7Ei2blX/kcyXnbpC/++cmWKkH7VyBLckAZb2+4EcHlpwScj9K9afkD3XgqnL1lcbCLhCJ
4FztlHcAeUlX9f2ae9Pb3DuVUSBo49W5mKYBw9kJdcGhFwmNIhWaxUUYloUAQ5gxZYGYqqQOH0QZ
IzSrnKF6q5Kmei8jip6IGiSWyA1WhI2Ka3FNf3d/dTCtr+Hx427pdJHIcuLv43nczwsuvpDogFGo
ArEPg25QZIUKsToLoY1VYmGh21PWBQQTLgJYzgjehUfbMX7d4j//TScOiSM00Db2+7nbuZ8yTymi
TcnyJV+KUKMipdIYvAi0bOk9vm46i59opg4R5rwoviOCbq1GyYYkbF3huGuEk4S9+ZEpLTd14y9X
KtOxMBCppqukqhlUutVZCwYMbhDyzS1S6qkZn2sTz9ynViT4Pw2L5IgmiORxJ90lHf3p0PvkDfyK
cWRrLiGtLYaf79qWwZCV9nHMalxM+V4K7HoSBmrwaOvILaUnk2XUyk+uZCl5f59CvS6A26/6rWr7
lnVt8DKaZaeQl0GlOzdQ+Ky467LgVu4o945HS7K0oO4/ybFd75QeDYlo58CQTDOL0zu2uN+hNVfy
UL8HDWP1Y5T/MmZiBHBkl+YHOKd7P0NDMnWyBxSLmgiJ3nBgyY6Z8K4jkD67XmAj6NVTMmXcK41c
61LZdPHrJKhRFfl0CutX2+Og/s8YZLBvxhyn+RlvFfkl3GzVe6ztiPt3Cm0S/fwqmbUsZ2B/iiZs
ROliajdMK8arH5Oym+2b4HhZgItwm+mepqH5KAIWhTfGPqKI/eWjW1Ms4uKid5464G4clcZ+8JyR
HEDd1+T5nt7n4nMmoKYvZ3S45Dv6Sd0Tzj+wVtBTo7FyCm8toVJNn4I4CXqe4DXKUd4jC120+e0Q
HGl14rSIyQ8HuREsMQBOttVLnfv9i2XqYLr6g52ySL/7aMi5CgqqPCA6aA+GkQSMW/C8B0vWzRhG
gbiscpMkdPL8tN6dHIwfr3nVeA+DsmKWKv3TDxCeUcjwGyxaB84bmzfemevRtKFMJjitX/elxOeE
qZi6ODZhpTmO+mHg5r/N0OqkUHSQi8DcB4znymGCseETMLqeOjB659ysCdZ6ZENLbZCGH1XxTKRR
MiOkm4AvJkkK7uf5a7PD+EnwEwi13W3k8IXVp4QoxFzo4apGMZQ32EyxZvufcQFVnac1tFAii22Z
UmLajo/3DI0y/RTooNQOz6EBlXT3VqD5KDiLcWuk59r7FnpTKCgqrbZRzLZpJnb/e7fUhldpYERC
3opdJ6ET/Cz/6lpM32vzCkLiKzZpN8uE+o45tpErmqRcmgk7OgzHN7ey+87WOSdlwdJHpxnT+3xI
LWWCcwQFqj3Eo6tr/mqMEX8y9EQ3iPimP1nrzT5FDoAyOnZRn3clmf1ZnMNoVo/2dRggnOJoDO+F
psdDmpImyF2kqjTvkEoQYJQddcc/IayFrbLrHEILn5hHyZPu6gqfUgJLSbI1YHQzlavH5+OwqPkJ
J9W7ScY5Cg08bjW4nFtEHuYC13C/+UgeMzZHbMGDVMBYUJfYAOJb4hG7ZKQ77wBvCW1ykz2H2qCt
zooQP0kYv8aaBomS6i+bl+oigqnsmCKSs4HmfF4zbnpg/+mkb97jaHwOjIUQvEM7brlxaU4N57qZ
qthjSbCx/R6fZcvBKIOTQ8iS4uW6H8n4Zrbu5Dw6sFjEb4dGOlPl0qWnWnBR01LPGzZFNCIBOm3U
2UkNvq8f8KyNZEZ2UuOpiEmY411r9SUkny22Kb4PHyTmPGhA5J8IGc5slwODkvdIq1UEPfyRdIol
LbgXKbVIt1ymxwkc0Y1ZTHyG+9RtVjygS1eluv1tkaKgavlaAapRSKvK1FRJRdSxDgtuv1+uDvdY
bhsNTgB7t2kR4MlFC54cYph4fr4U8MTWWlcVeb1t26q2Vrty2OMil9o5RgeHD0BXNFPWPo00JCRV
yUQJH+0gCjREvW5bLGogx/Pc6p05o1PtP6YrT4TVI0WmS6w8za8jYEgl5zGVtJo50hMTpRzOIjEV
vTw/mqjteq+UBNRdgUZVwvS5N/6El7jwliOSHDFToG6vqSWbEno19V90ey6XORCGNrTSS8YtYpOc
yADQzvISRQFYlxQHgZ9g43HHCavzNLqrd63qNe5Q36csXdzOZjMNAPIcVLN5UsS7Io5CAmLV8FTa
r7WgqloDiJ5jCMiw/yItzcWNHn6yTyO6uIfoYxqc2336iX9M61kj+nsqL1kDjeHTyF7a/ovC/WHL
MM0XQstA4J+CCGf1Y3wlhUjlLlI9uZossmQ5WX5smnH0H49yr01gD/mYfPfZfzKMcYEKmb78iJUK
Er2J801/RUEusBwaaVDJqIL1xiz0NTSEYVSUlFSVVOx/E+4wkVVh1YH+mCEkIE2KfUbCWpZ9DZDQ
H84pcF5Id3e5AE3cnrx8ulurYyWfuo5x8Lk5Qhxu2JHt/z8PcQqwmP47OS+BFMV4UKwyto4R8q7w
GF7diukTXHauzp5Orp0DGhQBttySDCFfVyBMpcyHZwpbBuUbfFZNWiKDreNtZl8Yrr/xzkzWCJnY
9vW3W7H2Ch7153eYtycuSq5XQq6BU24ej+kReLff6z2EGqFn0Cof12nEHCtlVKG5uqcmp0Q30XZ7
4O5s9hvOn9TuBIsGXK4JA4SfrSGpRvDz53193ff0oYXFocB/2Dp/bR5OtQw0OMrn2kVd+PkjykCS
R6VnwumBBC1gyo0SMYiCX72svmbN0hOwdbQ7lz4aNNUtqubMLH27qv+eBGx1N8gm55e4YgEtWxHY
mZJkOXHKKpaeztaOBJbXIe2rzX6ihvz5f02djxA6OpJtXal2/C5k9jw5mJ7mo+uGHV53B1XzZScB
tmGaP3sPqlWf83Ce5LPJvYjBQzMML+dYYCqKRgnDEs5vngTsL0Tfc6bZ1hoLl3UDg8X9znHo3oBo
nj9y4PNigS136swEMoisYBrHSP1MRE/MOn48oDK9g1WC80uqrBcqgENAyQ/sgWI85kqoPh1nYIU8
7ED1L1SI8MqkV+l4/Vml6Oy1WTcwawCrCrKsixsuStnz2FchWJH6nTxzdHYsIi/Qvy2S/yFZCONY
OoGOkgRd8RCVSqGU3ogjGVTgqiUv6Mz9DdEsiaUY+r+tJPnqA9SET0v3I5YMpKh54YptzZrEbpfj
HH8IPssQneVM+/pxzR00Jmw6H+LfQgfUAQ9jcYRFL2JXxORBk+xshYyVvmWQsYnTFWTMZ44QAN1z
UXD/PwM+S+7Kb/zDKFjnKleUKEV8yIlmFnVdDvEc+Dbj0ncfVnIjnx7oP9dKzXKWLicOaKTw+4me
wv7TID8+z9GFsgb3bnGt5uPgFlLTxcJc4tkpZQDCMij5ihc7XYaqOl/Lm9Yi9O9riBIxmssA1OOj
fppXFRuu3jYwOrjwVP2C2J2usZKCg78X0gJOymtFyJ8F5kGDrnVoM62h/GuA4eG0KMzmrKjOqv7+
FzJMlxzTDqqRxJio2U1KuKGkrCavaUQt19T4BdXO8dAfgjcwKYVbiggmRY/vdYLW9XZv135iGtOb
nr7ZRsBE7Uj344tcs3wE9gA7x5F353ubrJmqm+Nes4gBvA4siX+vfb3GiM+LJwEWCn9xT/Lz0Q5U
V0+FOHW+XsRoBcboQgtgQhSH0f88qtAgC/iTfFvOUSkPCkM+1tVCfUOMPsgezRRK8OHninRwcSkK
pEhhZ80Z/ZWBhsZ3QvEkt8+VBZGERRDgBaq3hmKfDp3DT5VCNzhEYi1z8w/pG3vOHxom+yd1FZjc
xSpsr6DV5u52Mkh0bgqKD1uxXbmS5udFpLnJ/jmpq8naFrX1gzeLa7yrE+BAB6cswDBVDcH/hKy0
2cWw6SSvtGkq/8AhHVk8F7WdOc88FNtF1rkTbVru3GcFk9+2ypnsxje6cJ0a1XzURLBwBhdPJM7E
992YnivMZR4zeEofco9k3oeVRPes/nXjTBTmcmXgSRNWhDzkPL/Gg+qu/No2ncfRxjUJqf3tyL/C
fFLQqoPLGe1HjDFmP1yw57tC8WCJwsWqUE0UhQ4eIfUOxo9ArzFSuJZAGuMISsnoBewK9lo/clQ3
Zr3KU3O3nOm9bzwMukXZENWLUh+aiwv7PnFAtpAKpuE899fbdBhMjoUD1LV0bYWQwShJVVESqNT6
GNs+HF0hzm1cJ25vKIbSAfuu/6IBY+qNJ9Unj7uwXhIcdxPLcGtzJ8bqNht8lQP7IesabA5twpTO
jaLbD/LfqqmlKfhbjj9Gl8lo2vGDWPsUFv+cLdtm6+35sqGBG+b4qh9a1ET4hlVAwKVBCZebbY85
/Gdtd7wtjH36QFs7s0nKKHMCdNqKc6aG62C4je2L9kWR1OpwqJ80tF7lz/8dHwY8mQ3af+MeNHkp
Oi23sY/Otk8ru2Njcfk0OXzUMuCKUEnwIAldoMiDvH394dejgVU/CXSATjsnCBMTxEeDlmtAaaBM
SFDUbpmC/MBk3y/aM+rQOj1EgPLPDdRLOeA0+D9UbV+uUjpVZYQVb+qMiLXCDjIlVxsJ3V5uVslb
vWAbuQMTtNvYAsMUZQWTe2PD7tnzKxRWb7EpXfru3NcKz1YQjdF2q1d94nZVbJUuQxQ7UYh5pgJZ
h3Q5DqtRVuMXvTZe4UMBY4artjHn2WHL3oLOcQaxAsJActmCgaZ+LmjKWTLrbMILukygZ/IqUdcF
jm3T3bmbpN65oNAXdoU1XdP2KdBIqu+CQ1G+krPdkrLbOIrXbEFrb4P/U9wLmztjWExMkosFELq9
spysPxCqv1m4/+qfzzH9sPKsqjYHHoqpBnU9LLmpFWIRkyUyya3OzG/44masX+zLPWA7KCJrjCDI
JktXrVbRmyKjsDFtXgH8EHdDa5bkFxNdSkDJ3DilY3liy6NRjw37wU9tVkqDEGVh5GZAGuQkGgoV
XDlh0OsOmJMwHjAPCSqxksvVC37ZCwLF8Zr95xX+QImYJwqMXCIDzRxFBT0h6w82PMg77MSTXTh3
CRtH/QyoRV6l/hGJInHshULzKnkVUnBLlWEKpMDoK1Ub22+OQwxr1XCINiznCGoSPfQbQ8V9a6yU
geu04dv4XESWlnQ/sPp/xxQuyCHvQ2QI8Ljg1jSFy6meMa1dF3XFZgLmkirVJqKuWpZHTdoYeILQ
YSyXdMo283doFtOBy/sL1FNrR2dyVIDEpsTwWnLrZxyJhBzucnRGNfSDFuEXOJMJSZrlZf/Zu9if
7BBv4OtmseDQ5qLaBIKEhS06I07GuHUvxoEcEstfi6S2E5ycN3GISVP89osrBKLF7sPdjb5OWrbO
agLipjVNpWp8KWFtbiDFMvrNZ0sPVwkU1qBQIR0rTvijnaUzUnXlQDEBbDTqjvroVKP7YUeSTHpN
o0ckaPyODsEA+aYSJLxBZYKt1/VSuyqlDY1el8Ss2KGzAhU3OaLhR51Yv3wyub8Fk6RG5TAJg9DT
r6wsArW1vUIiS5A6OxiXZXZJHzfmQSmC9ldrSpO1Zp8BqkKwNe9REaoGxdR5s5v4XFzgoGNkgbZl
LGP4IB+mShnrNvveCfGVC4yj+sf1JrX6oEaLAEpUO9xN+KIj1eg21L1M9r1aLzQPNRNeXAFssSmy
vVHnUU/nlqT2SqabvBhPYaAFcAW3HeSa7szIaZJUdR/95PLhoCNF01sUMKaZ9D3D2aQEKz6NRYQ7
yMhKh4chAuS54Qm5RzBUT8v3872pkrHAxjLk6NiS0xBmev+1HV/AR0/O5arbwNpYyaGiEo7gtcx6
N+iUgMTJVUv+rba85gi14mWKcSBxC/62Phl+CpFWFgO2xmD9WykIljaqso6u5EJul/b22QsF8vzf
d+5MrKUyEluN+GMlOoLbNvEwcGwNoTIRUMPyzUnvhXcvN6F+nqnW2gVVF52FSDd2ebRyLfteAMzS
ctXlFAqo9TipLqoOz8CZEo/WPIAUCcFheKqcT1gfYVudnJHgkCeATCPABt4q/l2l4X8E6PNNXI1d
xf2CS2rMRBih1Y0R75fLc85qfJQqntmhfBpy3rLPT6RjNbs3Pz5KDFEz/vzn6rpvxzTEuzzbsTh+
gP+s7nevS0Ss/KdzRUA6ugG9WFbMh2PXyi93FToGtiUMeTKnGPOUH1DW+BCvEBbosXO9OTTmgyuJ
4QJfpaZbCT8cOy+4RFG08tceyfisnqt6YtEfzSukpxTkoRJZ9lNtc/urZGXkRP+/RPxTn7jLcwjb
npnuZKQDi6bR1Cj/N23ju5DWVwQL6PH81mWcP1bJ6YPJGmRDDc1p88Nj/STAxR81OyccRE3gXXvj
lEtEwu4U8Tm+eWdrk2wvYJcJSf/eNlS8cM2/xJruEYRW6Yi076F/wEOPaeuJ4JLnBiwsY4RuZ9r7
7xX7cnLCTdFfqetp67diV5A5IemGn4zZjkDzGDmHf7Ns00KycsRZ0RzVxo4Qe4beWMRab51szmr3
sjs+ODmsVlDfWsszXsDFT/7oy6VF+oLqq7MOu5/DNQNXCV0uzZkjq9ddb05gSf0C82OKDIy5y1YX
pR11EXKSqrFzoLUQd8ntqExufLzE+16ybsmaUpK5fp54NiagdBklYf/nyxpXp9hhFxUhBec+QK2D
yCUl77+B8uYm6dYMp1HSmPKbQP9FVFJTconNtRp0hEU1dk9QwpwbV8cGTc5+Zvr+sxckL5t23KZZ
fc2DbQVPFHBjlYlrXEk4oRAsCyiNrDD3x1coHsGGvYwp1LhWBHHJDmkR7lN/KXMXSzSs9hQSHucg
HZTN/V/AxRVkTZ1rJUiTYw+9hc7AsX0ZE4S8d/Iww91Bkd25z+/lswkIJIJsRSFPwNM8tzODMGXj
GJbsxljwrwyY+sv753mYVjcVOifw7tmdDbwb6+nWvOsGecgp8g/CHfkMvI8+FpoRjDzXkS4bS9EV
mbekGRL5hu26nD2ByqDblInxeNaoG/h72Ppwo25GnQNkSjPT17PmWSmNE4vXC7pcavgWjzxX5zxt
/PKhkqt0AMPJhh+Pwuppzgkl53Vkx1/ZN6bbRI/hI3SFfdT3T7pCMvrpTMH6ImRu/BqWW3uJXMaq
dkPvqHcKo8LckEmgNIr5cKNJTYkFZz3XY++rJ4LerQU1aapEoM/C61znJSnB+K7Vv7swm7ubw0/V
wMA9ge9Iuxw2M5sMNOfPmnqEH7UIxag58mYZjvQVxXPF+9sHnC8NFuurb6wj6wcVaJgLLdXsL6vg
mD6NtvBwDc6qDL5ls/1iOEfd4hgMbtK3KutrKX6Af4RQ7Sw5OfFsyoxZrA1zJMvDD785JEEE0A6d
7jDrCJeXXbR6L7f4zsSc1jDYveCNKb25XEViKgZWt0dLBFnRM8kmhbx71d4w01HU/LoZ7bwMC/be
IpQKXwsl4OuPYD8sKmdr/ogrUfRcqujQ32znMKjsAPe6VYw8H+3QCGWzXefqjO3djNVGKIzy8rNT
oNWhuB5536DOnCt6Bu4Vd9fLpDV1xGw5K9VbgemVz/OOSZmU/Ywfr6Gf9o3rdN9mSfy9DCFUKUdb
Xnv14SXK/8aRfLnp2zemV3+LhJ5F2zV59mJ4ZdtOKQfy+aCQruuwXq3n9CJ2XLyDsBeTNzLuK3MU
CgwyhFZa+1C6tVCP6VKWqCSiMZ06Qn6XEYldY3srgUqFLdl0A5pIEzy9v/b4JZBYS01vrs99Edua
6ZuI5yrOkPdxwOkydxnJK6T1v/olbOBCw4ZhB5XPo8UIHfchYD6+7MlmClTHIuEN9YFGIbq93w/u
R9GePjsvoxjf7ySmbnxfIF8Yh8ea+BkUSi86D0PbC3dpLudgSL7it8vAIuZRV52JGaNC2vQuB0ll
HzAxUd2A9ftZmrMJD+UTMc6GxiehCCFZ7YlQdD7W9v8jxrHADMrXpLsiCsfGOOtYSxm0slTX+ka8
XvlBNIbaLVfARtxZfjrxz/g4KwkYk7/wSvikEFGGaFRcl0Wnthapw0NUcBCZaZ4+RsbrUHttucKY
UPC43+4IYgbldm4L4OzcyDvVC74abrZVYMU6z4iy9X8FMqBQdA7Yd+aNDTzgcVuFa/AmqKrepbMo
Por9rxUddqq2HJ7gcn6NRPv1esanUMSVfrlFK5O6BMHYxfG+zPBSqy3FgmXajFdMwvVp+YQQwv/r
bRgG6Ymd0upqL8cCKOCvDmHHDd0R0otgwWPrunTJ/230ntOcef7ufqw+2g2yjB1F7petS+IW4cQQ
rjEUxXsWwYAMg6BaHDFLlo6ebY86oZ7QkFAig2q4UGFtymWtWsJTbhexgLHY6n5f2Itzz/gKAwtk
M8B8hwIwkZhJvYzkTEMjB4rsIfweuAe9IBllPEKEGagqS1lEmpRjBsSfYKwqQTb2AE7vShU8C1Od
bW2+JfpkWldDR4a/7wPan9CLkmk9rI3hGMGIsDTbORxOqA6kNo4EaRvPtyFmOLI0GROMq6S/8n1b
gqsPuuecWQl6LNIHoqF64rSrpwYmyhTSMQI2i/q/UHwkH9IUM2CMiSjRMP2MD/P4gLA9QfFxZ8Ob
rwAe0Ow5UEWiChvWRX7QUY5rLSVxbXBYzbmYKKGdKdjsf5h1cEEcMOajRSQdkPquLlWgf9Y/om5w
XJXS1PDJKFc6MRmUwNfV9ORHBdn/Hvb/v0X0MYt4uigIWWocUbbU5HLiZ13w26/Yof/yFImz2yuV
vKNTOovyIM2t+UUUGHgFhKtA1vyzOzMlUAAxa4mOYYJZ+u0euxyxSIO/RQUcfk+9HOFFyFE+F1Td
tkAtDXPvphmgj38Tza+8vcT3fuLfPhBoaPX7lBcw2UoiozFIVFkqddQ2Zs3lQiLp3iOQISpkDbvO
PmHRcE7Wx6LJJC4SEk1XlIQMRp74efZPRnxa8XRp6FPBB6RK0wfHPhhHbyxb0V9HMSo+b/gRyEk6
juKjoLQYFlTtN3nxnyz7171u+4DhQoMbP4BDlMJYl79fPwwcesxTT3tAIOaq/Dim3mxBO1goB7ND
PS9/Zs5RQKAtP6FCD/iEo6u+XSyoFG6eEccnLPnaOxciG847csLqguaOerDNVqOILJrROFLyBi61
FzhBfmTmLorvZSTgO554wkCLNJu3W012c3w17wz3a5GpNXEotFOn255QKFfWXxM1BfuyWHaGX5i8
WMmvjVjKz3RT4LkNmikawEObzbRHzOLVoa27NXCiJjbQ7/dS+rWEalpoN2reawU5D381Cc1BL8FD
4ED0nS5rM11vHa87OZA5tQhSXyzFkH+Q2OTB+43mnIz6ygEZi8iTTXc1Y/LLKQaT3S2Ks8nwrPgP
hTYgmWYufCpTssGsj3oL4ZmBGEIM3Suf5Vt3rgoqOZqT/zcomM1h4WymRnUMIt+yKUfUrQkqTvQk
2n7x/XzNBrYR84xTVhwLQEf92UXRCp2LlfoytNC390TwmlEaPhYovZy/r4ghiIO7F1t28RTFbdIW
ldN8KtPg94dBHrTNv9gdGCi81u9rut2u0P0NchSCi8peW9daASuRaMn3cq5QTHdzTQloUs5MRXfM
uK6oj08uAo9QFOIkC1Y9mv+kPC80ARrczkHjV7DXIbuu2XRaN2YuGo7KoFmtMTbYKnMyeLs3sU80
MplxgPdCIPyrpdxwXuxuqh1N6qyff8zgyYVkTkb1qt2DGzfvMHfnNNP4w1Zcf7XU9ZGrzw4yJ2s+
TI2lo7sqpiWwFro5/5an/KfXSysHL78LHuFGJq+mnqW49ZnBsS/TrlTPKoOzyQtsXvaor/sbqxH9
CQ//KQPxcAIQcTcfRyj6DnrjVFEIiTt10TGT8QWfiMj67epMap3n8j2GECnyTAgNvjGRpGf9eK1t
Sd+UwrRvi7GNqeICDIWI3FJuUwQvlZCWXxr6k6hodc16BUow8CCbBJOasgqTJqhKMppBK3AY89jn
hkmhIBamn7RYcRaiL+Quf3i0xoylrIGVnaE4wevhjqoKjUGFAndgqh2C77tQSbMbtyC3jV89HcJ1
XPZDGyAsPnOkL+pjH4sEb/9CHkhxWBkdkHlhfpKWmBpzpA6JVrZkir2dGTZ/S+NTa/PxDLbWF8xd
Bni2Ziw0LoXGOdZgqMkGgL+gfk3ikzijWJAwbPPHcj3l96Ty9ukIG2M95sWOvC5zwfj98VThbyqz
SO82nwv6WrGQfQ9wnVH5pAmxmwM1Aqyvnt4P5l7SwKQtRfqFM0hn4gXo0a+ZqxO4LPZl/51NovjD
TqqUq7ujCn/oVzuqHPukuxKoj853TpAc1kbKp85/NI8jmgcmhSwvYmHvPrc8F2TZIs3aBBIh5yNI
6UDDqbc423SRoX5+aOu+bZGxP+/X6Uqa6bwEYX85BgJaGKlJhr/4A8ebmJlJuDG97p7qwc9OEyix
6Laacmfqbuhs5YwKGQk+1OlfhE4p/um8ngyLmKiwixc/Di2APdP9Jg2NcwQbVNdW9S9G8bPO1fnr
Y90e6he//AOGMWnqQ6TnNN6CVQkebgVxld2pHdc7UvR7bVBxlxspczbXJ4k5yB+a27mqFxq/u/sB
pIc+FYAeDEWUacuwvlEK6qau03lXh7KnPoTnzE8c5WksRq6AXwowSPV+rlM+TxzzrM6Z5GXruuLG
9KCFUIpfuCZ76+I9UPRER2TGRdtN3unK8lhF5eqq1kHwjvz8X8TALmbVAN0a/L5aiAm6TnGyw0/v
bIfAJ3dl+3Of3lte1abkxw9jbCP8FNyQehfueWu4SmrDLqGrJYjqjyOKD44qHI2AkLCJcOM+EU1P
45ZOIvzvy0yjMHLjDZnV4lsbLMNzNrPwYbDxoyMsthertTcabEyY48Uav5VFSYua0zoZSypKDPQN
xdfxpVG5vwGg5A4f58gAFO9qos6VWs4LbYzgrJCIkhma8vlnw/d/jzeOWfn7xa+8ViipGtd9kxbu
eqLg+h7WTeh9tx+ZdaVs5+o5VdDX2/LpRNJUrY71BLEdW6xVLILw7WshFjyE9abFinE5/v6Riyby
nOeFb53XTE3Q02Tj2Np8SkvHuba3c0NBDo5fZDmklpjzpzxMppS3XqDMgRtq+m8iwV/D8hcCay0O
k5FXJwDNxcc8BOZrgmjSTGW43acg9UEoPbu6KKFohAO7FNwY8OFMRQArIPg4fFaCuL639ouA/Fwl
JpA30nJWRE7vVccmm94NUHljLbSbzCA6jax9dBxEuBdRTb/UfLe6FJo/wjPg4NlYA7lVusysIV42
o3A/s+iuNbfG1bnXIq+2SEvGYWTHRXawegH+hQieNX9kwUnGdUV8AMJUFe59ewFBhCyErsAwB7Xv
LvbEZjRWsGoSAq33xI632c6HTvOrLqtOomBHr2HQFxNvqMxOPC6P7IdeZVIzxlCO/UIZHvNAKujV
DIHBi3CkkKn/UlAGZW6w1v4e0tFgVQ3/wxlsvVSOMLHvXV2WMjcJGaDhlWTakbqK+z3iX87Tgi4q
DziIpgQCeNacFWwmyugAW66HGiTyBIjKRTQ+x4bAGK220TgLNe4fsXAaaVEsktskRv5Cjrm/+5HM
PR9G0xOvMHBsG8I6WQxWpl6bj48DQVMuc1S1SIsiVqPj1JqXu3XriP5aYhfm7+5+A7fvDJydJOal
4KQsHyUtkOcqRmZ9NvF08pzr+QOcWp/nXfyvdqpqF7+hhf2P1zjB2lfpsgJ5Wbwanvds4fyKpZEf
KPXt1yB5kAHUPdTeSCYG9l2IvaaqY0NCn/6kmsfYmMDEw3QhOf8aVi4Phz9m6oaxjtXwLZG6A6KZ
iqocu9AWlB+iopGyu8g+GhQb4wZH5pOxXg+Qgyb4LRXtcJOJABtl7FBaWuTZJlyrcG2YxlO+kLHJ
KIgkrzDf6j5vCi5PHfL41GkYH+2KvfPK1BAu+979WiEIoo9KxAOQKy04KZX5SuHyiMAomCzsmvsQ
MhL36RSZme2TBZrZ22h9lqxs5cLZA3WD3RQaH9rkw7okwrInykVckJ5ZZNb8QocCBlgjnFjLGpv5
8ZM4L1QkGvKV4ztd+kfAAtU4Oy8E7SzeBfXmQXQ/ZWVUQnVGIfoWROs/JEF5XxOM0w0xqhGopUQt
M8iuSjauScwKOdTFx8RT5tjR9mG91sd0FGUy9IDE5ZgQ3vJu1SuX2WbedkwzloMIBUS6kxdRCmKZ
GLN6V0ardSjpBLBUY3ayUYtYZBqkTF24G7W3qEvIHYFMkiNMcKr2UUaevOQPN1RvndDUlKlavFnv
DMavXE0NXlxsMOwNnUxHnzYwVr0H9+kL/15duNwXe7UBWCBFP0SvyTw40K60IhNwWvjEXDCB3dHT
FJQBy0e57rZNCo9qrd5rpncfIY0aSjxEH0EDrFZ5uPP9GagJb4dHZWK5oqRuU581+W4UfUJcBRTQ
clKSOkDaE9H1w+6RvO5RvcnjIwJXe1NRbDVS92lXGBT4ZC7EJc8QoiZKKKV+ngUCXkct+e2mL7YV
++SlhCH/lfVSIOt4HquPiWS1mtrEPyZu1kgdm2CJlN7Y56t5BkBv93dpZMQRaK7Hp2K7FngevU/m
HyU3DegX+FcWnju50Dgc2niP2ZTbSW63yduWLUAKtWYtPBGH7Erm9AvQeGCOO3kd4MtyjYmxjNzq
TEKzN4KSw/0cbOed19w6d+m2q9mP7sC7qMQovFkSAFnBA+skBbYx94dwUEyUdavTU3QOOJGt/xoq
Yka0nuNyeXQHungQ8IiOnfLl9t6sMTi5HQLL18JYXTIMgyMy6ZNG1wTUfSmIpEBoaVJr+viOiCdA
ifvQOVOcjps0sweh24xJJdGV7jzDq9u0vAYdJryTS6dbh9hJWHiN4aKxmWdzf8+FFMUXa2CmHezc
znTR4LF0eVK+dRIjQYQ179m26qs9igGU8KAwL76WapbOrhX0foCR+v4j97Gmi+xV1jg59+QRJhL+
7I/hfW2E3iCZPC9wsPWcbxZLH4p5WWSR/cybWPseAjUOb8PvDULXn+qNdiD9KtbLGmN0prYhL1qs
huS+xCxv6sze27O/YiX+z6a+hPrF0M6ZH2qpvjD1fCDLIebT+K2nKnWJUfyFvZ5GVfLGJr2/LBFE
wpi6ITfrIxczXCr8DWvElubY1U7hTGV2Bka0t2udhCjg7JJOa1I6xnZFJZ4p8NnPz+RpRh5qswpe
/qVwnPARNEHTj636y1/dmSpKIA63JsIWNXvCTfROZKWqPjtSYBBKj9xvr1DlDqsrgNAFdjPllo5v
yppvsZmpBzfmX4rwTdQe8dfBClXMw36Uo73+Agyyz8+TZPkc0uLsPEu5Rx0J3XsxjilYO8all55s
h5+B8da+w6TqCsYk0MQCZD59sDpNS4gx31G1Js9oJoN58Gx0hRaEDIquw69fYvnDWeTWmXU0mAV3
4lNUqnAWZB2lCC6WUCiBJ65i6p662fZ6m5GM6iPCxZAAW0JSWVkDFftKEnFduzSwsmpw8fBg4Aan
FrQJt1EKkAJPuVJhNWeeDc9h0hbukGNYpsfSgwt3UlzzCQV0UukTX1ytmgoDn53VCkeobe/NaEAz
g5B0V/qgL8BitlPbzjK57s5rS52Nk62VCNYgRUzzzYpBg0VH9qAHaILTz6zY83YEosqC1SLlNOq+
lrNfUZKBX3sB38P39vLdBFBNF3908o3DvHsVrQPLQ5WXobSmYOt11WXc5EXR2BvJfoBB3zkFlj5c
CR4z8+2lPB/jjFMj0hxUpKEXF8feHy1EehzeNjalqQ9gP+cqEEj1MGg7pAKacMdnNoi86mS/aFBr
zmrKf3TrzPgwqibbfCpteS1ihthKxxI6xCSzwC1dqGWm5dTbrBOSg0lms7NNlAIxFYeUbQHdYIJL
PnSpzp76Lca8W7fhtVjMRRljsjJE6sO0746tBAZFRn4U9BXqDvxX1cqKDxeN3lxyQKhYNmATI2z9
bPDU9qKau2G4qPfdnRqRUeMfbcXlEux+K1xTYZy0skq1lgBCK0hT2wLnjH20KEZYRUaXMInB3bpx
d9ckdm3qRUACh32tDYkzGTp9nTwDNva1wbDSBMYJ4EzCHHr3cqyaETAjESkO3EibeH7tuOzK/Art
KB74p2/e9va0uOJaTpDXeJo8ZljUI5Xh7rqrl+o2eUScvxxBzhG3mx+WMzkwU+vP3C2cM5bdqp50
IOL85HI+KpunbXqVzTmx21/W2L9EIhZoNqXoHmsMHozmhFkF076lyDD0kehJeFosuwj/jEIv848B
HP+zXcxGvzlEw9kgJuzztpkga9H/9XB9RvnYQh6vNRSZa8qVfrBYBheoA1MwqVc0Kuc5cyvzuH1r
QpANyhQGuwEnSWPx2Nnq2B0IrcsOEPB9vcF0avnVatXX9foMjj/ORo3XzeOsjOQ0A0EOYb0iTvAj
xir+5bBQK2Ja+uGH/r2UEq4yS1N9jox/KcX9nvdnQhJO2kwLayvdAzejCFPDh3LkGxcIbuNc6lGw
8TvEN0qNPH/72RqXb789KiDR2hmCryFp8yaQuCgcgcxIUMWR0HTm2RkhHX2jmgvVlcMKClL9ZBsh
612Zd9HMTP2T28IPrA97U8Qn0QtKmJSaz8U6QEgnd/oDZEVPgDeVzhBkUQvzl3f7/gThJjZ0wkpH
Nx4KSFh82lutQBiG88c2M8XMXLH9v5Wt0YNNdB6VAO38rDgb/Q9Ba10U8uWWJObbVskqp4T/RAUY
4rJI7RCn89pR3R7pr2ZlEB2xu88mg8fT52O981wyQkkgovaLbxfhvYv5o7PzPSIl/xDuQjnOOu0/
99aP75AofrBdjnt0p3y7sGkW2s443OIUSlRFgpenufj9C1Cw6Wba+4O3zMEf8I6Mqx/9djsegSHL
ccYap0pTJ8sG0UhQ5lw61nnPHZM8S2M2zzYqt2QDZqOxdC0f7ya9VM605bVH+8IWpOSaf4wtqfg0
kwLagJcUytPQM5Ghmy+VywusuzhzhCmU4OC6GGEzBwECGdM+h9jjtUSRZ4P48emZa/b9Y87Yjn67
20ctEKdxBzGxOS3hMrRV447Y37AbP/2401YfS1CYp7ZQPqoTifkwGlmCTxc502HCoq4+qvrXOWNh
3+0YSlG4GHV5NC9T8vgg+CBf/01qjRw5o675b0Ii5QRhqTx02p5LRaynHjGYeLNVQE19a7x27vYw
X8hqg9nJy0AIeX/SIUquZpDhFqaOEK60/tCzGz5EGoWMmM+/WdNYyBNrtluLMwu/HErkhCSbaJzC
S0Aog02wzcoEPRQJdeSYiPwPzSYUaMJl0SHtBCDnNIPjP42Coe9o2Wk3V3GsIQRxgq1DNXn84WxI
gs7mHiG4J6AJ2fMzy+mkqgr6rLoY+aDwWdopRp+dNPSqh9yuo+v6OZ+8kh67nOaLuqHYNDX1Kjt6
TJ2uVSd7TiIMDZVhydevQzjp8Ovwbz13uRqdDmUJF2WYaDO9BYHzAAVeTkqzDgL427grol0zzDRY
sSzb1sD7dYzJR525CDMzBw7DmemBf3WGb3JAa5++lTgjilpMXrOpqkTwSJBaL88VOvisaxGfUFkp
UAMRUKsul08beVMHNDO5wHm8PlktpPfOyOjb6mSMZUqxKk35dA3rQeDdxnzzdZogebuYiM0BnOF1
jWpwBhRRTGO0u31JyFlKEPus16yVBAzqvkBbe8g0yR9nKCK5hACjceVKh/7Aa5iYdH3ebUoA6z/k
putMZoAxcyyOdC4Im4lnh4Uei/De2Eo1z21xx2I7IFrQlovV4sk7uu3RVu7oq7ub4E2LIJzKu4zZ
NwZoUb/XbwLAfbfUQpCwp51Y1ht5g/swF2uzol9s6iqyLNpiTtPCJtBK+0DnZRJmsaxpDcLgb7bs
13OwuT7sZwSJlFzB6U3zVCX23YI8zzaIWUpd9kjN0vD4INiV5fq280IMaZVICDU0Mml/uXS+zAbu
qw5a8UnZ/2PY2NDD1cOcO/kvzqABFnQRQyzrdTS6bFpEU8uXSwuDcGAc3lnqA3NHuLUmL19wlqFg
i0Qj8mSqDOWYuOsF2daRarYeRcgPPBGr/CHsadd4G3305sS8oskhbWxQRBuED9vMZ47BnVe+ugyM
670q7fkZR8LYQ3lADXgvSQRh9+8B21osVvlmIapcbTYaEGYqNfjlT6yNUCCLRMZFpL0cAI5VInee
9//Za2IzYZv9WGPnd8Dmxy2PGvxKLL5uWsDFNxvQkRjM+Rlym84K/wmN6O0R12uSGM07A9QTf2N/
G1ImSSwpMSH4+dSeIlrvHcKApZJkiHQcHLbgIeTLjfG2K9KbANzFa94bxI0l1lbeRVmtyMhVRlhF
nn2YEi1xvR1zSSHeEGkva5jiwu7eYUNbMMIyQnQ8L0dL4+SLPL49l18g17HsQu7S4ggB9LpdENpZ
+tyGmL0eVxcAtgylhVuwFjcitGZ8cMFF2WEOAcAIYx9mh0LxZSzVTVezPdQC0Y7QYsgYtl3iNT4e
6cnKFxoz1qzF6kgwJk5P1HnCNyAsxsvRXKkW3iPacth8RWGKUajgYEF3024IQHkXVugBKH0x7NdM
Mqs8G5XK6IHWjwccZAFCnr5orq2WmMj+uhhOaeHx6v6d+mM4Aluez9pxBenEHFbg4x4ESqDzR5MJ
faVaCAEHgpdJns+9zlnPIeBvsq3Qfmwwve2C3f/LF+EEppyFWOjidlrLuejFOr73WGiLMJFM2XJ0
BOjlIb0FVrzBh/QG6VLE8P0CYhgnRyNV1JKKhhMiT/4u2oncxFrsFxBk+SP2+3V79LL6s99govO7
8c4nA7p4G+/ZKKPHB9FEM6lVaB9/Yg87zflDNBBtgeKK0Lwwih6ZgSqRrP1xKRQmkq2gKh4xiIap
AjnkDJj/EMa2htc/17mrK4CgmOTgNMqS39mltqqYodZBvmjrVFOAIoEocpSTsXpi7h3IktprIaNJ
eOd1G5XdJNdlehNWi+MHk03A1rAS5Bu2crgobdSny+uBz4+QrRJ0N4LGMi27ojTqasj4qqob+2MQ
IatveW1fOiw0g5tkGU2KrJQbwgtREBeTh08Z6P9zvKRmHIfaDH/kj3wiq4IOhij4Kv7hmuD+bHmz
O3cA46oNPWygpqMd29tC/0f+gRuT8dYxAvqCGAixd3KROruvQy+7hd9TxEBdnAPipv840DNi7M4j
ySrIeaCNwQTWzAtI1oVnDf5DuriXzypM3SN0B3Ud1XsdOmvlG9ZkBLReyYrCx/DP4A+IF1h9AF+X
OgWTYmQxofScx/jyzezr9k22DjMgwBTJlMrpBTNbYtq4E2coFF2CqllStarUDytEMo/yyASZ9Yya
hNI5+OZDYqII4T+/YHxEIm2QW3qai2uCK4JZfW6sY6aQVyoR1VpGlIEmbmkjLjQsFsF66qdcX7pC
OrKc5k23hlH84s9Ds6VQJEYvF9y0hqYOkSl0pAnb9WZXaFBzvtcLvogsZtW4OGPq7jc2dMufFnIs
j271upW7dTfukBbr/Om4JZw8AXBHkCpfvJYd2ajVNJtgQZNCSQ4Tqxz0Nyz3jFyeo5MnXrYVoM74
CDKg/fJaaMAhraeqIX6Sa+iOgxink3nJS4Ywl6+hO6NU/+LgVNZQhdlCrU2YTl4hkkRF3b/IsNdJ
vgO3jt9x1OwWSQ5tMn01s2T26mF4KXfosiiL8nLafabxlIkLq+LseFBhv301/KfzQF7fdFQrSVLh
ACCQhq/6Gi3VCmxa562CCi+BDLCDg5Mq75k4wTWOKG1EKacNDBE1nDLDiA69R2R+06AemhNPMCfC
TQzzHtPgEAbEEOl6qBpLoHzqZDeDw26YfF3t7bWxijaBRrDrKJI5J6uv1LeAdk2u/Qj9BRUMPUSk
JKQk3chQr8bNjxhseLlua+QeUShJqtZpZTDwZNVBw5J9IKlEBzYgK5Wwh9CZUcl2PYNyWOeJ/cFQ
uzHJWu/CM5B240mfAVLFo2aF7WbnirjowfHla+F/BEY72ljtEL2XX4Xkioao26oxf7uFrzo4pdiz
fC9QMptPKyMIl3hcZGgYNSwX6WLFz9nlXOXE1OtO7rmf0So2oWFtgH8aOO9/lRjoJo1X1abWaZ8Q
efxaINSUHly2rqNeyBYdf4zXNX6tZGQv3xuuw5REukx0bekBWNykFTA+bnQmmO9MmFjRUVnphNUX
UDB5wbraM3BxEkUyjC/C08oy0UowIZnKFQ1VpzwJD5RHunyjf/fMct+kug0Z2ijOMHh6Gm8o7T0b
pY9LkatiqBmVyQyZu58SL56FkQPW0f7CufqRY7kQB3oyr/qnMABwJli/8C6fgxjgePs+taOPyxRo
JmN20o0uKXGgz5u9mAQQSZYlUN0n0kGFsuYVp4kyr/WcbPjTEfTkHFHWZBml4qfcsRteUvVdz0jk
SF3v7bP4OIs/x7926GoAhNtKkZWtF4S9dn91sRlR/kGfDvi7pWk+VuaQkveQ6+oXhWbobgYTa7g5
28r/STaTBSlyN1z05FsAQl3flHSB8eCrDsK/ZWkNqScAgxCUhwwzJAkz0J8wqRvFIOdyytWxQtBL
0DPYXAG1P7/VDZ+i2xW60nwPO9N7rlcF0zElqqwkrCVqEF9ihVHcxO/jophIOnqHAp04UA6xVc2y
axHvNAev+icq5rtkdUq7ZzJIcIu6K4PeP5krUMZKOBd2FmRCzWPBw1+LYfgx1Qr3uTyh6kj66wtr
dHmuOrcwXLPprQhivdDOK+en6fMdPBYyS00ZHQnZisGS5ORAEGQM41vVVdwLK/RtzaSOiDTe/ctx
Iq0hlwkc7UyqvSdQqqB8uBQjdHA58j+Kc0lv3L6puhEAx6PzZcRAIAuSVNi/TQclYbgHQBKtGvpS
fIxR31uJDOrn6X6MimxhczjRDLMRnxoKMka1hQrK3fcve7Z7WvOVuNhmYAaOzF7Z6gO55ylPLgEY
+3Co80tlSwoUz0xdcgi/9KbZ0vib2i+pHdvPO0luuFRhvxR/Wea+U5q5a6seZb9oFcNlbIqQopRS
R2QA6c0RBnfzkme95l9BZdfQtgnjdIKLsD2DomnXNlzyKCt36YsLWUfb26ukArGsVubX399uLpCX
JoaqZstx46ILanOF0LFoGaPi3OaDP7LVar+jhXVSPK5+yCEfTupqhoJHne24vnKZx7fi6BTTXYup
JXbVvQO+fcfunf04TE3aUGbrGG0KwgxTarXIO5ehGlh0vapiam94fUc4pcWzG5SYOB6ZZfnPy+cA
APcdy/bmrOH/JbqfzR5L+gHsA2az7Xgi0+q0hU3ha+7q6zOOfKDROObIA0st4wDaP7QSOMZ+dS/I
3bepL7doYe9vkU+kW13ghiGFqJ/XdKgIG88BOSOvqCKLkpcB/UabkKPhktmLmPW96LOhDlTq53ex
Bt8Th2vsJysPB8gw6nR/9qG7XSObt5P/jSU84OW/wELmaqdZJ5PkMPfNQstuetkEed3PWR42T+tD
mDyDoliVzMchId7/BuWySciaNGIhp0oxs4/eqYEsnJkvHcjLEFt2NCf+KXy0prN3MUSoqiDiAHZy
L/3fpjwiGc24P6RYsnoLFebwvDbk0ZzEL70wzPSlUNh+WOIF6sPMIfCmHMX7cS+Q1Of8Rq1MWKe1
CIchJBdLJ5YhXbeKoTvdO8b745HGBP3pDewnKEBHuffHq1yKU3N7OS4SK3qQDkEsWRQdeU/hWrqC
U2ZrPkp+6+MoBNRDMEmrmOdHEEVrVVJTCpvAGxAi6Ko3kWZYQdZ8RxpYJbA/6IBcz6IlP1L6Tsw/
qAonNIBRvOs3QAsUnRoU/97R03gPWvQmHTegSKIcFzpX4YAEYdG3bZbWqwIqe3lOG55IytchxmUB
VUBMuvXsGbpOjmhdSyErIOEqlfgYEat9GMbcUD8zvqbIoeGwL6arSeCFfZQrZxiKKsqpjPZSMeqE
1IsKmA7td7FrwomYcjtxidSLagmGg7x0BTEzqpxHAtRu5X6PMK6VHALBHn+YbMsZxchOMqMrXi+r
7eIYffSFqwDZGPHnWM2gXRz2pU6uhfIYS3DxuqT5dnWSdSrAySA2c4l87vsh4c+9Y4bajioH4b+B
IoiMFIpxyuo57NrXiPXpP4M3VoJDDvaCFKnN9I4JJVjkyRBMcg9nD4/T8zWfNWt/MjpJVgQzKooq
Q/4z/+MWbXvaD9JjY2fpbddJ2nAicpYnyIeAjsgR/4NFv75eiRyBNiGIk/ES+8WpLDHV0nNnnZwY
FoEjjmZSlMF0tgyP+Dt2+hA7YkLEHup3JIrOLC/1dwvGCevLjG0j2xkX9s2cLh8lyUK16zxlLkHG
16KPxHxmduKxCRDOBpBqlOQTZnL/JQK9ZJSYeNRndmV2KEoqtvnc5YwJr6EqfSgGrm2x7SLVYNkx
BRnuQJ142s8zLdYzdDxnIrAK/JDhZjQAv/NAcGvADJJfx2YtQhdw6DwX70wB8FhQut9z7JDbyxio
Tfjm1qcY+KsZQvQBnOhEh5RrIr+KpohT+W2/9sWdxjbb4ssLoOUn5Ks16EiiWg/O8Z3w6QaMg2Y2
mmmv/ump9RglUoGq6S843clULZVLUyymD5NJdsFL6XxjVl9NHwXUzhRvtKU0VCSBhwmwKsaIAJf5
+3A6eg8jUUy0Y1dKXrWhikY+EI3JKfjvn7PiZ8f4cFHMzoUrMyMcMGFuvPItS2uWRrBT2dw0CkPw
pa3KSv7luh0UpP0h7esq5JAmdoAEY0HzvLpu595ifQK4M3+fKEodIV6VLChRkSZ0jOciD/iypFSQ
NLRW3IiMDTniDjclg0yMiRf9XF2hhbh0p0wIeBWdgFdJxc3ne00C77tePpKNVK/8KNP2v3Z1ZGba
w2+lhYf3nJiaR9QG/hZEjCMl8Zxxozbki7/aDBZynr1GxgHiN1Sia15BKw7HEmzTY2Sc/YPI4T/S
Gw4BWbbLxUiCDKYPj8oRNjKtgWgMXo6WpiPTPZUYQKjMMTMCTDRJh5Xw5vW4o43m1ueiPSYTiUaN
MkIipm7OuTL3RssR7oxNGt9pw6w/ltT0d/Wjkuw4A4IszZTEL6xxPRJsnknaaIbNzt+BGKV8gewr
POOAvBnM80nJNu+/49i6UHVPx185IU/biB/UWYwJB2KconCpzAGa3Z9POBou4sgqCvrqqzKBCh2o
xKhNCYe8BictMxtrRJGuweRYE9DLKJo0fGhQixBruRkNI2YljC6p/c/rStlQ5H1xqxrJjyN6Ehtb
QOBo0dEq7Esv0bcoIrmn9odn2pSSefyaVuKPZWa5cEt/pnebFhJ9Xc0Xn0WFlQFfIaqJad1551qz
UWcC3c7TkuDgRUm1QCG+nBNUV0kh72UCYV1MphWwutvQ+GJ4h05fuYqv7Z+CdyhRtQtTODt1BG1M
jK3R1bWGP/ca5QeR6O8RBTbq8qxlTz53A4Q5foM62vSLOoYA1z51o1GU9DGzJP1oR7GVfOQjxHTW
UaZLuToyuOxpsgPWSTGXB1i5kStJ7aHI8ivBOfYDz5GH5sIkfYHsMjCqsfv4bQMEGxIcc6+zOqRO
zDga407c0DNa8JFw19QL0i9QRZsP27RQU9nPgCLJ6YARvR01F9PdPsCCqIhdK5BcjamZgq4kvGhP
Ga9p6DUMpuGSbLhLnGGL30PkUdQiFg7lhM1iexu1l7HOv5Jfi3kBcqdUI5q0w57fLt4/jKFhB+jN
W314Z+9bkCLsOgyEjjZOskIltSVHSWQ8VDXkV/TkPM+vIxNmL6/B7MfAWxtKFjUqb7/VSepH8LPM
t2gSoX+28dYMhwj9DuRT2a/gL0iHABwAKcX04fsjrNkos7FGhac44tYoiGpV0ANCS74bOPvCPrtk
nCtayXIIHl8WwsoMglY0n+/DndD/GdhaPwfWrL4/NLI8qTM99Ruvq/VZLM5NR32YFdFLBv9kbwWp
H3mSNBUFApYKKTOZjtTlWiAuOsrlMCyMizEzd4GGnLfWPOuiibGTNTgQoyl2JL57bYU7SUJ/asLP
ndrOHHUqscPeyUXFQ1vhx0+A9XANLuv7vKhjHiaHftuK2GixU/W91+Cx2X4K36sldzoo2AclQvBV
l43zdcKwi+lp1DNdUdwTYjhDy0HvUb+tU0rkii85RLd3rhUQwil1NVI7LpSs57h0DBs/LyfoYMxG
S5rOuxmzTRSME+PKlpElIRkkA7OXqOQ/KOQBqbi+7SReeCZEudCPJm1KMU/Xz9skngiV/noRp9kp
6B3rN2L+rQQqzPiZmnEq3EZzStHKuNQzFcLVAg5n3J/tAdI7IkJhrVsBhGrJFRqK9r7//3JVMIfu
5oVcMnul8AKIVVC1JuwQQmjo3kIJhfokuKt80AKAfaX6AJsB4fmqJ4jOiqlUmeO69SPxkjab1zfN
gjAmfdUGVBl55UcjVrl5KxWyAzuVA0Zm2lHOB2OfS87Ip8MvTGG3v+cgOWPHq8Y+ntly+4SruHcf
H+lkQ8xhJb/qJ5OvlQkKoy8VAahpNBE5J0cPYIE0nxvMYiweXE1Om15pR0/oQ5GQUTrdVH7l1+dx
BYqs4r10pyDVBYFSdzEmDk8iiUa5zABGVz2c6vqLqAXVMW7pUWNzNyYvbxIkY3szJRxulgIszGm2
avaT1HqxcsKJskdyd/IBQsNBgFU352KhO7ouwhDnY8mqCpX8TYnBsVr2+qJ0revzbCpu3EjpAKsg
ZXwRikCBYGvduc2tOUNpn1MuqUUAUopSlWD7wae9Df2XpIZ7v/YxgHLTqfQijyv801SEcddhHtc3
moyN82OkkZG2Lpzg9hkYUq/CWh1M2KBWJh/HQha4X3LYdJomkcHOsrM8p8ijVBslq0GVhwi506ul
QrMDegEt+PFUYcMfcgGnwpigWQrB1A20uKKPrQLBQ0NvR1MeT4tLzqUG1CliC6aVNAEHrreq0z+C
fwNNE798d/rFbAoStnyk5/0Ep8BoaP7XOqBWUzXadqO+962kUli6G8RZDJapoE4gw6PDynWHTN09
oBRzgDIsw0RQlAEqGPory79wpQa5f8F0vNTBM0nyh+i1gCjcWmSpTWZpfFxHJhDmwpdeCmjaV87G
2hzt+wra+jxc+LEljJUP2mSJPy+YvaAphO69i4csn8+crqdKiCtJKJ+ScVC6Np3NqV7ojTeGBsL9
5mPXdJN2dNoTCRaQ8Qg5AaMyv/OkVxez6HMlZps5LwWu3GD0LqbuGrif6BeadryBZLJOX/MwsYuH
D2j5OywlgB4CInx3EkYEpqI8ZqHsNPBqiqln8Dnv+jXH2VHOPU70To3cLF26Br2hK1BXWD0Np4dS
QsyOPs0n8ZTp1w+WUvdgCIRnCe97LGMLvR+Nx51x+j7ZrKE0k2cefIP2f3pWA2L8kpmnliflQKHL
9SpFC6Td8iRpUVEOeXrpwyEIgEkvILK03qfiu0r+MFV/4ZXXrxAO8iIvV8OQMYtQ6doM0MsAO1q/
cLBvFeZ/yeshfrzZlFwl316Onri31QsKMCKVsKHPXzTdpH/v7pPpjKE6p5AswhY/zLlS8RP6EIm0
2NTFXkex8mIqOZBTlrwWHZsAw6Jz3AzgOHx7NLvDqILOmhMBksrjthvAuCDfhRTVeOFGapvrjXnk
+vbHJX55h7YWX1ZS8Qox86KCOBdYCYiEXldHV/0L6A68/DFGepCvp/A1wnX7lSZnwgNW1UihXQgV
ZnoX2emzwnKc4F6o6UH+fmsknEYcSLIEKpDBQXm9CpunXLnKcd4WOS5JD8Tl7p1mdNvWZuEm9Gmq
sXudbGJJq9V4tSauh6DRI+c+2lNxuQZbQ3qOWe7YC7UkMguZJ9GzF8oimKrcsrSzXXI8IYM/s4VM
ZueSGEboC8madXX4R5mSllXA0SWRIMg3Ulw5PBfqhCnOicybC25FBlPqgF9rVBAphu2MYv8TwIh1
2w1wmrhk6Yn1AlRoWN63ouL1QFv2+EGmVSaE8pHDOzwGE/RZXoj+yc2/6+qHHPYZ5cRZ6nCmaa9g
hZGOdAcfoToBodnGJDtjG6KDwI47n4MpuMsap0i8QGTr84HMwFmBYP+LdJL+uSJoAX68JNmwEvB+
X5uyl7Vq+PCF70gUnX3BxHXJ3Sc2PcNHMtf27XTqSaiUzgubMk7JQ89rr/Mjhx8xEIbyQ/JFHINd
aJLDvv4+fj67i0x6gtzBPRfVNYlBop9XfSkwUH5nBsnKZ3GNjDH+tvrzAzNqk/eIbDFyrYCrFPZp
t8PgkKf4zpnyRrGGGMvNEnqYf1bj5AwtXZ3t2GWddET7fC/AZvbilDTmuoP4AG3uwCPT4Isvhh9p
aBxvvazS8328B45UE1YRbCaBJOm0yfCaMhunLb1sIRwGN6PVmqgmJdnNzJHrZtjBTMxR+Hl49qrE
ZQjpOMOlI1kdZ+DKNFODoEzno8DKvtOpxPKvXhL8ntuHz3fBAzD6X2f9BpCbrlqZWEszAXqUuQQu
G3iog7X2QYTy4xzIKmKUB4dGh88fK5XmV0aXWTZO8Lq72/TBwTVUBmwN9ckvMVXFWGRDiSSb4707
thnO1RT4wmJx9wKn2aNSWr8OTKlSPrSSmCuEXL+78eVbOzaruQOJLOlN9ReRAnuSHS+Go3jnExCR
72eYvaMJSY140ubL4lxvjNM4p5Yz7+7Yqb2wkZse8yJuqshqkW/HLx5gnyR3l9jD3SIoJEUmXaXW
MACA7OKkD+xxjVEW9LMARSE+GXFQ8dkQAglsKBmLdG/ZezeVdFfbgmhbOAhMut5jEFX/bAd0ozd6
8sC+oMIszpwjlWHPJS2pORL0SRXgN1VWKLQv6CJmHst+jCZupyfIgy84rPE5cwE5oBmOC9y9t9sK
Qy5ZxK3YZjSL5WNh7WbX4nMtnBE68zVlPCsKnOp06dKOIHBTJlVQ6H5aUxD/+F5zJFVuFW0mn7Ux
3IJgmm9kauXSA+BmhkF12LkP64+akFdIUpwdExHsmkLuc5uZX1lnFRNW3kIJW0tfQdQ41UzKGJdW
/urfYHxWQSAhkGbRCMDZoi3/43mfYtFS8iDztCob8muF6DiAzMFwmyN3X62dCPXaYzeGylCaMOuG
TgKDD8bBRBYNZimsbbNJTcOIldZBIrSmI+yNog4WWAFBjZdBTafarr73t9E0F3FAs0EHT46UNKwC
wjK3Aqi8zNCcl4AMZ/dPmrUyKoEUp84e3loL5yO5sn0HRmk2lcVyKUP4hf/Lrf972UqodrVc+mib
HD8qDxNeRouJtKvVgVY/kYyXr9g7JvoxrjuSg3E2cbsVDHaED/snOEl72tVm5Z/k9me4rFrvK4Uh
9oGYKCK7fe+rj8ba626AqD2LkqcsZ85GiBOHc2eEAInx5rB0AN1z76DzMbNtozqmuuwu3cHxBUJl
x8IiE6lW+VsIyHq5We05o8RTBuIPzEyx4PhEJMoPdKep/8NheicIsBOANe69JDHg7IUW5rjXNICy
Jq/l5uRxeeSyZUprE04EAV/sQoUftI7aR9ZgscUz9Np0oVx2ooa+D30QUZvlBj6+cgTPpHDi7VjK
cF7pO8SASIaEQLVHYis9sxNd9uO6xALxElf/NSN9uUmwYuMN6kuxHPMh2RFChI6v+tsieccvXgy2
/xHDRvuxl87A+zYsBxNiL1gOi/jPI6iryyVPOgMjSjyQuZmWDdnr/GoPrUh7GaEeGGmfy6Z3YSSQ
7db9IiJXDqhIqTRgxWjZu38+japdT4j5rY2E6dM25wMn50xEOzI/JbC4juHLqEprYPcI6Kp4j8s7
g+YKPEiPpp4dle2+BvmFCEBrw5FMiBDD3JzQzxCk1Vd/RQ/ggfAmHpBEHmwaW+uoNZLmqRgltHCF
JJcRmJ12XJLCqOAb+CYK6hV1G4O5MUL6fknkH+/jD00a3KMIes21owtO9cuy8Mv6TCaKA3qHNAcu
wBLKXuV9WEbTXONPHTguEnfPPPaxU5cZmLf9puFLNq3aox3HD1PfX1wo66HqikvXT7HQZEGA6lmA
sHNja0KBz/hVLzv9qSHafbStG2fQKU0zcqw44kFTmMetGjoKippoRScRQyB15JGoZY3y7rXP4fGY
yK+SHw1BrB8MA0fXBoCRn5teIvxnFYnJryoO186+VszmcxZ1Jd5g6xdcKHf40osiLGwBYucuFBEv
Dc/bfBorNm18LmnpNZ4m0bDMlmKp06BJy3NpGokR9wzsXFAErJ6gq+NkPeeu33u5Ws1rgsV0I0zQ
JZsUR3BHLglIkLIhp7VoNxItJEEQOtgKLa0aJ8s8tsZRlSq0/za97MpLSoLfDyCaj4A/6dJv6HFy
0qp8ncL+fGmgLaEiZ3aHB5Uw9RWUVQlTMUdmNZYO3vMtxoseJQYjSbrBe8g+N8FknDcTwwO/YuKr
OWXyynUBLrCQB9JSUcvrIpdzUoUP+eW+feucHLfs00MYlH6ifVtiDiLLW8a6QKPTV3RqxS+p+2t6
1YiFELQ2FrsMt9Whl0qFZzPUbtsd0QDRWRX2zrDEBDKUh+k7/yFLhdxdgB71NLdLSxLOVe3ih559
UMxY9uvjoG5X6VvzqjiPm+0vF0ZFwC5/C3M7RASB8bSgfL9KCXw3HmRu1WNybhTC461McH8jn3Ew
m0gRc9TVYrbPmLTTMddIG5jaxUVrxf2CPA2ftB4ukwb4FVMbqTw0LtNa7ojG8PoBLFlszqPZ4sRU
3eBk90hWBIWnz94woZpvOZnzd/M06nVaI2nPZ3vQV6xxxEbm4eGQ0WYAKtHGzK6ImGpBdl3Hv8Li
p+NaJ6cepeCtc6i/jK+WkeIzcfivqyAZjZ+unZIQTuVuDRyBj693AgPIzPVUUW2p0hIawxezS22W
ZN8SUGhjtq+rAATsmM5fpuVyEGjJFw1kxx4HfRNvrNPPWObBhFZdkfH7NPHe6StcL5f1DlslK5w5
u+uhXORQ270/KLwDT58N4W0tLrCOd7O7R6w9r42zm22CXywkuSg4mL22TuckXut18gW+zp5FtOwB
TEEikCbZFIV/FnnIW0faKHREVWcLjJtJ+PBdgymBU8IdFEolzDORKmrWNQ+zAutcW+GfhuzACTNK
Kptd9Gicrn+j8i05ymGpTdzZuirlx4E2dGOuFnhE17yBr/x/O3U9vaEKLrZLvNRp00xvrqBp1Q/c
NqMEZeF9u8dJp0gmOrfA7nPBAM/tBe4HPJV6aFRfUQ7HDQgji2nW1LthySZGv//tTy9WRRheYdJg
74SUwIK7eczS7AqViw/88WuTUp5ycF1V6pmSBgzgCIN1NCdcYmfRxrGd4QdhqpNaRxQqGOsSxhsV
80IKh7bzsF0+NBipH9HQVng6vszv38fqFfOLEP20e/VCUo1w7d8lUdU+hKs97KLIGnKFD0S2NQfn
56K3iAOofuNLNQnrG+ywovXm9ei7/YyLjYWdbrsE3pkV33nrPd0haMSKEKQ7j7ICIIA1TB2GKgZH
LSoF1QVrjyYjc9t5ivmwJ6MRmm/GeZKy8fQbkGZh8jdC6uErlFAakXDeQOXcs9rTRpndN20td06I
OtwxhlqTaws9/m5moUdWjPDE4pTN/pIq3kmRUzbMKqg4FRZk3SetDrn8otZLx/C0E6vAvNd3goq0
JVLI/AhxFCqG81wOxnvV77HJuhuiHxvVwNNrxUTbZfXuSnTomSYhopyjbdRRXFY7XW267mL09QYn
GU7iORh/UqoCal3YFtXmRHtHGBB9gzLWzGTdvlrd2baFT2Kr8Qfeqza3hjyb4YiRgEeIADpWNoTo
UEQBMMJo984bY25tPMy5iI3qWGXZV5y9vZy/zTH6PNgRUYQ5xPH+S7W2xUC9bWAAzGWeAQ/Q2Z7s
bnW0CTFMsZwLrzuBMAM9Rv0SZhmZrE3fYByYySzwhh5/kSnY/7MEXUfhdBBWCH+DZ/WtF+G409YQ
aEkCFb5QqyhGjoLL0S1pED59/4Diqpi5Sd3j1iqFYd04hC7QfD+18mqN5Z/Pe1aoVi3+eugnFbwo
RBl5I824kgzMjr6Znnu8fHnByrs0xCExMeyI0COtJGOyJnJUj4EJNwvr9YPr8p5yClu1m08vMnxI
jaxmE6SqVan/VZQdf07T0oTajRBBZdPww5QPP/OkrwnaOjElrNYnAsi5lPmS9OuxFAbAL2tNsAtW
VntA3JlV0pQ0O9N71QMN4UxFvvcw3KzUgYpX/WGB50lDtHDGQg+sbxinQqqvM1lOkM8U4SnYVV+m
DO1yFYk0KDaBjHSevdj/J/9OUwvrDYVSqVqgawOzzalxQdyQB3/37/l5It5fDY1ck8g7KgSMFdJ3
L+MtR4yPxM82D7fyDKWJDGR3mC4EV9bpANSTCYbs7ldmjE5z0JDcYW3hPfgr10H22WXtFEShgxZL
GsskhRuHu7KB0pApW/eJyYU1OulidrK6WakYI38Wwj7WnwhmXASYBochMAmQ0oRj3TI4sRMkjRhf
BCH5HSsGKcjQYXpGgQl5dzRBG1hTvW5nq9u1cPMCqLOQRrw8Avw6FFmZMoio8+G/z8mA4frbki06
qpUr6GysswF6LgajT3ZLYqSJ41y6kC962KnuVzZZqqJjY3qEz0WLv5nQdeO2lXuzaP3vlc6YSUhr
7krSc2/GVXUDQWURZormLWXkaV9r4ulYTWHB8FfZ/8wGHMx2GD/Go8BQSDLPiTuS7Y/MIVsgPVAS
yeKTcSYfaWhHvlQ8TqcD6JS0JCGx6L5J2TYbzjm262hnqhHIFwtnbFPb0W8idfCNoiBBEGqA1PGZ
jKKanAxQlSK7nRAcSFG71/3SYUuoSRYJZ2HJjmA8PeQI5jSJwuqgIYoV9cbwrS14zpaEGRVuUg/o
dFNj8X5w5DsirzV7r0sWNdjbB0vsOoZrp7l+c7ySaaWFza0kpPQ2TtSD9cAkl+8LXhwsur45WZoC
pa7FBlslJnjndSjSw5qpX2YPthlbk4LoqOquhhhXgaoiw+VdciHZ6Xg1wmrNc9L3LRcRQ0oAZWtX
YnEnT9da3lwgRXDOU57WtQMPtS5ZnulrHgwSdHuTw1CXwUWuMG9eZRJe/P1mPhm5UwlYmfBPlpNk
PdK9mupTdNdLXIcCc89S1oc2tUYif1onjPA0kNwzVGaNTUK/ImsLfJ6Vb+ABOeS/EhaIdU9OAfgX
V8JgViRaN75NJuLhCZIUG2Kq72DbjMaP7B4tU/FFPAWmvgABnWB4H0LlTddrs0Emcj3482aKM0X7
gN+p6oEy9lUML0+snWLthprvhWfyFtXgIL1DKlelv33h+XSBIF2DAynzE+7vUbGr8JkHbSQbXpK4
Essn6iU8hPmF4+eR1anXv2k9pQiF+/qG3XL9uFaJz0rO3BSEt8dHIXPijMDlBZ485o2HWlrQZAAP
ZGADj23wGtSXwVUGSENyQAJo77Kt0SWSNAa4mTZnHR17IUPmvFSQsjCrdGipY4yNa3gCLi4RMbbT
7iGKnK6rdcqlmavbnH/yEVqafg0+bMD1Q78jrQMOGRBsqq6/ApEs+qEpKydBvdZUA4a8ASSwHqIb
Gv5CQtOu3LJU8aMAc2Yc35pd903uRznLvW2CQ1WQ0j26ErNZfPVnUfDA/CtaDUM8OrRGB2cMtX7L
IfyqtlyzpnkOUTCfy8lrdbtJHPro856gTlZx0gCyfBY1YkTf87lucd+mINshnQSZ+5jtXhCnoLG1
9TcmGIYJETMNwT38gwtPnMfgFqm8jrWDpPa8OHDCT6t91mS6fG/vajzQW+ub+wXpcH2zKkHt18fO
mQg6SSs6PEUpyE4qE4zpakWUy0gTh2Gy0+DOAQpeVOuXXMZ1ZCAbOXZc1lGhuEaSXrue6ark5Px3
JCEbPJvoMrBbnpBMoXt0oZUpQyb12TfLYguG7zgRTQZZe2zMgQ9+4syNYcWQCTPO/jd4XsetS2tW
fdqL08PllSNFqkj7Ds2qr4u3ovAH+QBckl7gXz5877TCqt0aTCA+9/DnCHBxgGtaeaP+0EareDVM
3rbcgzTR98LjTOCDa0Ca1bT1fyUXv2j/7NYqmioRf4b3MgK8MajyrkdYFbq295cKpeXXJvw09mrt
FzUmnhAZbWdGDD52jB4L7ENVZJlXcYMha2XkZc4UXKv+vG8QdS8vlMfYw8cXI7e6cIJ8O2tpj1tC
PSgb9xVNFMPf4F24/P2bigzdIZZLRqI3eoLNJV8XKH9O9QUxa9MpodE33i1Hp0fLUFDMdUgnxwVW
YP8LcGWr+g8wcpReD30+DUjHiJA0McejOaP3qKICIcJykwqiWeR+6ZFAV6RrD4AWSjutjmN+iyEY
TBlDhlJx+nf7CzOZeMlry213BdMP3jzfu0igEX+NyVtIyT1CEEOYHd8wzEmy2yyReP4TlCiPf3xW
2/S3H9D40o2DyaCXjAvRgDIBjhuQO0pD5csmKu0SDxf1GkIVhkzAlBhCsVjQlx3ub8xiqehSJKlE
vuviDfJvtIo+Aw8Pe6uUCt2IWQe3VwDs/NbQA6kOOlyS/W9OfKjeL3xBPyDGEIwFfVQDx9Q7RmCm
Snq88ly+h8FJb6qpAU2PhhGyqTyXwhhj9sm03bI1bqYzZHtIs3ldfrExQlfk+YuE07744xDoKjuf
EqpLvAUypW+5XSDqhONJKoCsuHqVeekJF+toXXDOQ7RJ0I5sA+2EKlvDbj6CLTyQbJaLwen9EVy9
Yj7ZiDlRDgFOis00mX1Gy6mKMskldq97awVsQC1h9IXFaFS56oGyYV6pUKBF+tkvzj+5QgyKnbS7
+iJDslMOTho91Z4dEBzNFf1TUAwbKnKXyBPWz+pqkPPoX8g+aNlFgpCoj+R7jotS/7yYeUIUUbY8
DrlXJZNHjt+2KfBgk+sf+qEpRkTcTPQ47nE4gr+p/OjJmTTgoyDbG5eZybvpECMnGtXBrn1DnxDJ
x3c1xZ+dMS/KoOiMo+jRca3r87GYimwTDALuvx5ADuhNQAFHujdUORXiwhogntOEluoZSe9T2mEM
D6m3q5bfLOEWqnZU9wqpEB3Q0xTiXYaKTyC+UcUKD2/5/k3OakcaNZGPMAB/7rjAhg3dujau4DUz
U+1iuKMfERNhxPYtKLC/6VITEOCuHMEsGb9nMbDEb76ufGyYUNYy51s8Z3ZE3c58pcei1j/ZKaRh
4RkQB98Hxwo+OjiHfcgxanphTseobF0KXvxOjwZr2Y48etjcQYdJ6IVXGa894uaMtxLgaR+j8UZl
BMB/+ZhHfX8hbnpwymYeCTUNtHBX8yeozwWMpewAPM+QebYXo8TNCaJWkpZE+cSPR0Nuba1xVJKc
F1tPzYWvXuZbPd0n7R5s9fccurl+qtG6q89wFWLIiaWGVH2q/eb12iUTC972Oz2c4Q1yE0nsReRP
qJLgBBC+5UONg2MP5OnBa6+nCSxiTAO93CtOWO9NMPPPFAsstXpXtQNcUzrtB+nRpKYBvRULcBPs
nmV1zUQcC8qpF99SLctVoD0rEd5A0oF+RyOmU91G3hrXA3QwC0rnp2MPyjTMSpowo+J5ZsWWgoGw
3Zkjv8Q7J6lbexxR4byCNEz3VfguRzRMtH5j/PO+hPX98gnGBUqGEXTIsSTIDPv8uAajouLP7Ib3
1bWXYlHxPEIaQtCV3E3cSqD5poMCx5uZRwebnsP13bbAEST73+4t6eQ5yhyBDR64tN2195fZxm4N
YtenfI6NqTSATAfkCFnjqEm7INxtgX+X4W1GEVq/PT/Ovx/SfdgNsfOmQIgrwuJyio++y1IjHth+
gnmfoq9i2LP2HLRfPP73OYe7KM6szaxO2y+OxRc8FPAS+Er4E8G/ZxxClKFi2SwSiM/0Cj+GJJBe
yA/kJ4pjNATGkY+2BcUg4US/Nvm673/qW6ZOz7jpdY40aFzKAuUFf9K7MCr4jgqqRiPLoqoloBog
wbtD8ELwmi5YSbuXlFkLjDRWP0S9DFu6lCESwjVwMn5h0OVpZjPm667hcPTK5St5a7SY8tLJ28u/
+sCoHD4oudtLBA3QsTpCgBEnu8tscwS8DqUs7joFp6cUZ/CW64CZU221kG0riytPVoERPrtgltrs
76fyfYBddYn0MMn5HXvGFRNC+UDW6R8ZOT+r1CDtOz4mPtx+XeO1HW5j+DQZcVeKwfXwhebw1kPX
jJbic6pr6fm9f6NrdKpxxlMdtMLTax3C6XcEQlvIDA9VK5kYInGVLG8ZOb3y+mMQCaXN1OEvLkis
sSjbpjtGaKS2szXq5UK4u4LK28ACKP65LIseW17iELHV8YEOMEQA+gEpr+XZ340/oInN/K7ui+Ro
0UujU2WY3l8kpAHkIsZnhZSBk5elHNpr5u6XRtml9zmHfYboQvBEfXS6xfyCdNiR67ccZUibPEDt
kfjGR7zq7bjsxF01XDqo0vIP057hlxbgUYJODycqejmSyesrs+KDVwSZL/N8PGYKq54ELiCmluCm
pY6xUsUrwTmoBICEwbIQvbuV/gcIRljSo7VcAIGG00FhAeZ4dFV18hLRdhFBSZ4jxyhwQ2wa/tar
473CpP0v/UUtnswVUQ48oi5mWzEu9nKdpv9Je1g0GKUWL+VDslJRK0C5NXGlhjOafjkoTm4+GvUy
H3tDg9iDjJhbccQ+yGoInOYlmWRi+XmdgMtuM1XaxuXYYO/T0yYGBvgdKzSYRU5GnubYK7/hUTs8
uYDYssbuyxHm03XJNV+SQeuWu6GsT1bKKw5/UlYOGCSnjTA1uXP1tbsZpQX1FycVIprOoazMejo5
r7KTrTIBmuHL838EQhUu0OqqGL+/9e1pHi0rasAgywbv9zlnklLeW72sdBEKYant9I8R5J7EgxbN
10T3dofiX0aYtNsv7OU0yobMmWeav4XU6cem3U2OaF0QkqzbGd/bH6yt9BtAbmHovs9EBkb4vXDP
DOrOsqeiAuMIv+JfaPnqlbxE5WffvaFc1VvHNp1VYIoazOABP+YyhDyCeGf7x9ZmPCrOCnRNPRn0
FHIhSvmouTO1yH8XDJdJUJwv7rO3nDG2M8N7XLJ6ICtobuODTJt5rfNhKrjIC1raEqTOvWDpmDHo
8XuMfzTFQL/iK4mDCFyIb+pqXSJh8vpm1LV1abt/ehCdlyV/kM8Ah108k2lXLfK8AfLvLn8zoPyq
a7Yub/H06sMRMqMiIQhISI4G0Qwln8dxZr7BSUxgB4PnRQDq7ZxAMv9k6N/h+bWFkYt+B+khm5XG
XUzfCrA0REB7g43d/cqYyhvfWcbPzHvGNvA9u5pt1dKncr2B89iwmY0g1AyeVzFzgCxhpAkYDGOv
7Xm5jSA+VZGCuXzDe1VtyU2vMDJlsgEvJgFxnZsiddEKbAeGG9DnwTN0EeJhBqSYCO4HS730PzMk
0BqLTGAptu7eXRvK8DQYEdWJ/DrEixxvm6r7RSZ3mBciXe+028EBm0VhAcq+UrQWF2yiIaKg1zOP
1pddpXY4+VOqvuCbGcrRZFfoM1wgQNGsnWXH+eQRlZuqLA7IwdOmfGDYpzF8QH8kd2Cl6MEGv+G5
asqw7nuFSCep5ixTdV+QzF1JUOiaH+mmrNKYCV1Y3yBAa5P400sUGcyrIL7N0YUbjpdL7vXMtXF1
k65ES1KKoxKlqP9x7UuwJMO3ES1OFqb+86qwJWBcuQJn8uX6FOX/6HyFEVbSHCDYzCEp53fijDx8
3s1oW1SArEpco7+aQCWcp6nY1ePAALMP1htejjIioXODysVSplvPEmCwf+4A7BEe8oydcXp9K2+W
+aG6E0jDWsJvQF2IQDmIq4HGIKt7ZWiRxedAREKxjsTeP4quuLwOzThuHdp84AK2KTuVidbqS/EV
M0hN7P+zPTWrU1tKbMwGYlzsC7SOnxjIzf401aEOBttDsRsCLCDAeq+xao8LnYuZuA3GJ7ha49VP
j8vlLXCVEvlGD3H6rHd2DlD6LZ/kBK+blmAetalnYZUf6lTp2wfwqiz1qISTNuTUAv/ypDqP3k8L
ORZi2HORxTWngMXkJeNodw31sKA5h/Bl+l12b7BAnK99EfAVa1c0hQly25pLsvF2C+h8WNaB/iDt
zqPGYkUMLkLtNA6buvdd7ObX5ZqJuCPa4zLQe77unsoK7mbKNrGk2Ub9R9uQwcgxwM+6ZEgZceqg
yuFqwqdynEZ47Z2WvM2GS1LP2sxVxbZIP0W70i5uHUUXpRNb0ffEA2Emn7/NiOmYUhYaRdP0WecF
x8KXEDQVBUor5nFgnuExaoFOGdV/n+Ru7Yer5f4NcZ75wcnalOS1Ub83izVlqkN3+FXK8wnnkjpp
Vk5v27wvRT/TBNKhON1zOeMaCdrg9dFP/AuAOQNfjamknbtkMnxP6vZee8r7OBo/y8ZCqX15L4Y+
dmSnSNi1vIkY9swEGvE0CTIrzT3qNanpCFtnoEkrxbkrN1QEZ+cQkiwq6f55vgy+oz88X6at9BjR
X2QIhFdpMVCO7RMahIHuv4jh/GTQ0PtldZQh8V5vJKegEHbGmIi/b/aXMnHCSAeQGcdTUqfO3puD
4ejEluMNq9VnndqVYklkTlgkQ2GNoBUR7t9JLKrlcGCNl1HlVYw0IY3R8W0qd78YRknuouxuraip
NmXQWj0zrF6SJXEkW5uOY6Xce9Ow5I7GjRTFkBuhirivCHvXOXcL5PrC7GTI6Ns0r/TDZzQNgnWG
ZMm4rKLOSHCiIU5vgpCrRAZarJk7YRyPCpR7RFN7sc8a9PLU53v/6YE7EgzsURlt/pHhtpIlDzMH
lMYgIAdNRqRl+tQNqoPv1g41hYkVXwvPOFiIeYmKuTEgBc+IcERDjBFJLebkgahEXVtIpbpUJqFX
8I3VNWxWHNikwjawQRkwmwL+4QFoMOcfxPT4zTqxC4Bo4P3yqPzVY+X5h6MXxSxgGggtYOk48+gB
KymgE3T1FkCCi2lQgor1lGlmYxQvMefJe+9yLbWJkvqeFOLBVF6rgU/vvTkrZEeOsIfywwPlmjs1
7dEYAO8Q21VcUBicAfqDVmG1raA2Dx9EjwRf/ji+dmcoy3uOriF2pTw09ccOuLOMXhl7+VJA0wbU
KLTkk/vPJ+n+FKADTy2v+9ayN/4QF59aRopOpn5JHa0u7y71PnV2CeKQg/6gl1RYyhpRY4ip4q9Q
5gT3nRPCfTXiYMxXMf6XUe55BigaSNrXpxc60HidTxvcu5av8x8DPr5aoQ5pVZO29/e4cfMu5c2G
n5nVvJ18Z9Z38ycfYdpthYajbPLS8YCIl9x8WJDPiJPDYIpYQQ19xXD/ko7ploFFBcbNTmtKBqEz
MO5rnRVKfyUG3NOSUj8BXVAMOdQD06FbgVWmDQOG63jxKF1X+POSQ5Q1zlPxeKjEPtwjTDdYXoZI
ZnfxLisOR0FraD5lGSiGR/Ud3FZ8Nu+jVLCvoau4iJXaKnc2AjwS7TvLFhl6QNzx4g45ScwXVBUs
ndUHKmSJzR30cFMaCAZkJ94g5/lKQdj/s7ckNuKsCm6thiognlzIpgWssWQ3QwWttbxQXQHOOYmG
vXlQSMndJTCeD9tKY5GiPHEXgBsDvg8vjvwe4Dlaom5mdmIRVPdPe8QztLY4I9fQbMzcs0he1oPG
eT+S4Q4Y3IkS3ysBuvRcXQCMUQdw3eycZbZv+IAhXrjicZp6FAMvbrMbmA+Fn2qyzK5+oNr5uhs7
NJQMDl52RPbTxocJHWoe9mIq7d84ObJhvBb//6whapIIWWXw5TgUddO7N7imQzOi8VOmbLlPKCKC
3Xh7OYnnKg8J93V5fBMm1/N7xmnwBHu4omtBg8SbdsOnZeoHl5a1X6/46B6dWbKAwwM3reb97PN8
u2Ml3mlNvqQSNBhyuGPxl95yFw20nwFuu+w01Sa2wMUJ0gZBd6rK0qiDt4DXkvQLrFbwtHgoCdff
iX84+bpJvxNinwmu5hVXxW7kD0Ydv5uSfPG/s+e40QC8DsVyGmFNty33r8mv0G8lxe8C3cm/2hSU
07uvHQtC3sV3dl6S6unLQUJOJF2RSX1f/F83XYhMQtJ0XLljBUlqGx+V7PVr2hNj6wpO0FWwupLf
SLE6RZNMiF0lBheaZP+4iXuH7iV33peQMZSFaUv4zdv2rX41x7BMgTgx22TfKhLiPiPbKogO0F8e
aLFcs6TyCW9Zrl+BbHwX4YehJftdA215wMfd2OpXgJdVtbKxXgVaS4OwKholQZL5i9J7Fpn7NB05
icpAwe3NIJ272UjebaEl+6eH8wAKMIB66RP1jHLbqN9K2P5505hNkLwAfaLsCsYy7qd2oYBYddwl
woiKvY/igY+jv7h8PCETIDZoCk36xY+lj5IhBA7HePSnupYMq7oLhU6hD+AKx+HLsMFCDjxRbm4/
Kt1azCH+rG55kXvdIXh+ghvS4Yvqhedxg/ft5k3gStus1PGMVgdi3QR+R2Wc7cbjxF9eWBbvGlIC
RSOHWT/+RkViCtkcLtSuUaWQHfZGbGWRUv8IMZFODl5ez0HjLbBcWfyrMSXXts2LVhuv/0kpdEM9
kokn/BWcqdGc70SizTXM6oD6XmWfFmEoqOm5O9OeZzlk2vugLqtCYz8DYPLzqTF4JoJ7rWRzrT9M
HU1IzgGiIyMap1RHPYGw5CnL6LTC5jcJdT28HnPw0ufQQZSYc+YtdZw3IFNrq6peAipOu2m0L1SJ
V+Pei3qMk8YdZ1I0Fqb35fVFNuNV2Rh5herl/werFAqM8osPRKQabkBUeZkmNDsHxPOeotQ3KvlE
rJTamBZKOKqyQCnxpq+Tkn4F9CsSoc6XFDVzmr9MG3wrM3x1VSuOVbddHGNdF+SEbbfq/xfqyDaP
AqFJPFZrLn+nP0AuAfvX92Fx0VH7FakplTnI7cdU6xO2/3ZOgiqb90nN8lgBAeNmdI2koz56ad7d
oAi5mxJzkv5XPI2Lu2mhdPjEytQlvIrtOvlOYFGnn7afZ3Xu+BOyUGx6rSmXPlhJa6UwvQdQe2HW
n4lfw6BK8z/j70SfF6BgBjYU8h8Ni4F5hABi0AeWLKRY4dLzod478752Q+x/NXYXo+pSmwaALY9B
vI/xnLc1GkDmK7wNXt7nKeyNYSZvBuJRBvSnh/tygyyqR/ezCQZ1UQEyPNAu+Dv6uRRkX9WCLgiW
dFQAoUCmz1+1LRMG0VkyiYIzEulzWzIxkA0gQ5Iz4juuWEy3WsyjFdG5a9rmF2OiWtvELBVstkFn
pmVknqxLPnMErCvBMViOUdTqPMpkDo40hcX1tLe7evOv6828m/2BXrDpB5KCmurcm6oAf8tRSE9s
YXEqMb/4EmO7CV/5XiHvB0hlLMI2ki3OXrIt5g3ruDks+ibzyTbUFKWypLStLO4Yy31UnoPBzjMv
D0xBJmHW5EsZbSEGlhAXUE131j8hql2BL/98Ovo58ef8VCu8HpQMUTNAw+tZ0sDjEEsgJbZK8R5C
oRCvsfZfSLEx0WdqrmJLzvCS+R4vG+cTQANRrnkzb8zzmemd0d1wuyRpYR63qbY/3VyklNFe5o/H
IEIICovSfkujAMSErrPcCzDDgHmmjXDs/O0Dqnw/JzXBjgNBouT3wCnZz7OkypcwxCn3zPlhU5bl
tmmkI44chz+idquRZJvbf0kxe/9FSDzwtMlD67g/bJ+M3zW9yW6LFZ6yMABtQgTejLb35IFArVrM
b4nmvidLzlqWf1f+eS8l5cdiifQFRM/idPwz0/CVoF/ABK+SKYem2e3ybxSP1Z8cP05Fh38x7vkN
ubO/ObRHY4Bf6i6yZ55P7StRKUOZK9Y5Bu7OKmIZopgczHI0nyxoEdIqShOHzUUbbzIbBYbfUu28
Ry+OJcvpr7ta2kGfH+z3fTi1Ywodtnb1Mv8kxrtQ0MI0wft/UexxP4//a+NuWJOtlYO9Llk0HZob
X9LuiSTvcf/CJbuE8v8cnf1eDQdtkD9obvrhoIp2FEmXPlcSQHC95PEM8uIlBOTaUHYqGPKxBH2R
HGcmV6218Rr/73ZobbZzdCXvBOR3UHte6NMatcuQdNSCOm8Ame+/ozATpzuXpeeLpCe/yz5C0ydd
/fI644HO4RqDiVrALbXQGC/XDfed98sRF49HoNdAsDTH0o5cxqGcLHqj1gyT/R+wkXk4rQd86kgr
8PwG30/l40Y0bEwtOB1BIUbtlQYXOVu/0GqZOVQokFs9y184EZV77vgw4FKPK6X/JSzGjwpQbv/c
qFJ8167WyR5GZqnc+6eRjeQr/zGxsEaIvJlL+6YxmupnDvQekgev5pB2vc8MZ25Y/Zu0NMDFjNU4
vob9yMyZfY7zNp7bb20Ky2mmwDTBsJlYgpUGlOF357JCrEStn4RI8/4OEDWUGbOLTfhaf0VFEW09
tZyhQHfRRM+Knn8qkxAo4q6dgVf+HnrKosRz8B8TE07VjgeK105OGmhBTfXmcvy/Kl3wCdFn/QMA
HfndhvxEGumS6VnMH4v3BsO0SgTwVEjZ7XGAgi2YNEF6Sw+2Z96oUWTBh/CjV+WKQkaSmVIi93Pz
WlRrzkmMtLrpFagQvflJjowxPZ9RwsYqncIds2DkaQmapLAXwDzkiLKjSln0EgKUPlYDSY23uXdg
Nc9MCimDH5+wafmfwsEo/J855jO84gTKf82JqeOyqzk5lRUs35UVhvBHVz7yGM+LDVMyInJTQxjd
G56GEKfhkYcWuKiSqgHe6d8nmXGa4hFIoutQ+9DDVKiupk5U8Fzk4SQHF/tZyKgqXTcHCtLQ3d4p
LzdK7g0LzxW0gtOvZET05rn0uYNOcPNnxs1VNh9uCUzyryDsGrKDIZrtNqhuI3GmFD1c5PRGTIhB
/rsVwjQ4jEmT2jD35hzCBI4E0BgATCXa+a69ZbeV19+JwQYGfhPJ21JAnSN8zYU6SS4zGFrrwkQ5
XwwuKvEr6b4aD8W2n/qjhKpIX4VCNO7Hpj6uwDXnH6CClOPqO6xSjyaRAcNhuHxoaKcCvP8A63FH
WPokIxaeWk6voV0xjtvpEYkMEN6T1ZpvEx3YpjSvdqkEMg7jIa8ssLTcszMf9wmXjICuB6m3YJMQ
hbtx+sDKCcGfVVqaHm3wE84knlyrRlx/eCckq/sErQce+6TYG7DOONCyVuMPKTZ/MO+DNV1Am+B6
tekBPTd9nCxcJxq/QHfKJuTaU6LgtIt5X4jVagNGiL/G4W7I/wL0IOkCGG+eyptycJuhi2qVorWz
/Ecd9vx+qxRa5w97ta8U4VKZ7TM9nqP28JXqnUt18Iq5fGpLdw+gPU2lU/oZIAFq/F6WmScwjchT
UMPsNvxlutCRQrPnApaxFgrrGLQPwaPYsDqKj07TRWtsAhLKllCt27rV5eqxzX02VF3tVCbLDq2W
VF9HW3WFEtAxb5P9aaHZKybvfOye7BSfKs7+X0iJ3I75ZaudGcO4AHkYDEdjRLwYb7esEpkq7yVX
05NRXf07Sqz4iYTTrHOh1NIofZ15raPq/1F0oYGgzmEEiHd6S6KozRSsu13T9iwhWwvbVz/cDRRX
fKddkG415QyIoE4iEetzSs0vy3XnZBBc35eeZSMjJ6U2p8DfP8vFf4p0P7jG1Ge3vChQMaFOwY5o
GRFtO2VDtkU0w5m3cMHWvoyNtRiKTcvqIdOOtcV8ogvofwgq2/TLWiCsCZSlr/xjUUrAgviZjOlf
TSRIkOjvB5Bt9aqh5RxNmnQEz6gFTtfeaFrjk29NQQV1sS7XVwHbrpglFHdudz4kDoUWZ3GOtzJY
Y0yBejrqr14Xly24p4QT+TbfnEVLIBuzZiCXA4Ja87y8jfC/C3IFoEp2jNVTVWzVDtOQp/Kng1hO
hLjc2v49zPUOZLbTYCZ/ib4ggP5H9yM+swtASE2VXM7BOl77QbOOIJdnyQXkFeiYgoa8Vvgvh3Ix
CU+EQBSWLRjsbwAOyUFj1C8O3rzniyPtmdjzwlkriAZur4nlmR4LNPNX0q8sbpHeb5euXQo/UoqM
ceMdub9Bh9HNTcAD8m4gcrDyvEsFzSF4TvGtIJEPoiQgEtNzeS8GH50keP9WEYuiUOgBispoKlgH
78K72ydk7JC0d7cY06rzipUzYZ7rw/J/1OO63Rbpxmpyw9zRcLcKd+A9jXF+m6Z2C1n9jtrmzM8+
NoAiEkIKO2fiTPh8Z6PEg+T3dAH1wtq9rkUwZyXVSigmdKXYa0b26I4PIkZDzVcs1lEq7YL4bDMX
TJ/QKNPN1gTvts5cfqtFpdNFkqZ030OBgQ2F7wyH5/AmDWgigYJEJR88w1n+ljbWNv7sI5qv5xEi
UCFRvuAFZqIhHWYcawYbsH236R4QS/KwYkkzAyZlbPoj+LcUlLpHRTE3TlZGc+dWY94re+4wIcpv
rC74WNpXGQhX9P2HP200wOd6hJOdv5qk2JmJOID6RAjIpCFukoHGEtPWV20YF20fIpAVeKF3ECnD
CRYx6zx+lOfAUVK+X529P+NGmBOKF3lARDtx6cD+lYnyVPIvbUVEx9J3a295C3CqGGpITHz0smgW
FKOkdUpghQcb8dQBe20ozwK7G57hP/IRZ03MdN9Ny4BoucS4mUGQguRws6IvfVcZgGj7HjBWr1sj
NVlqoTXYq4j4/9SJwaiJBgFZTRvsjkN8OxLnRGpU3cxtYFXYY6qSP7Y4xEHQETuqi74oWxbroCfn
6cNTG74pnPA7vJ0FEIxGUljW/CmBp7wRVxsVmYdoOiEpgxyWcaUc5NpkFlMsgILc5Sas6mch9Ipf
BtlwWjKl73483M8Eu29nKqh2aNp4kyAekOPCdBPFlX5A163TEa4YnAVUpDjR5A9YaKzQhofWMb8l
qihV6pdRFOL1bgzq+9se6+P/DCtCGmA1RSmPjn8FZ+zt+7krSj+N341NFRTFvmeUvundXP/S+2tF
+ymjAzuyWvc4EaVy8MaDpkYzgH4+p6FPWXVulVrVeRb+nzVsas3MoY32JxqNauo8ERPuzGk7YDxQ
gK1EWtwRGKvKqD+A/hC2/h9VDMn3jEqPz/Xy10PJAcp36uebDiQmxaIEFn+AYT5C+hhixTP7soa9
giElPyDnY8FXRz+xoU8eGPmyJQ3Y5otsc9RsgkqvEgdld/PH3vii9Sz8eSd1pGNBSNfbyMjh0GC0
9kxoGsDM3CVXO+YNgaDXPtFpj718g4VR0vIfIgUKHmaEFadwoWjHIMeiA0+iFaDni5eKxQ3leJn4
2EL0AlsOca1e5hYOaqHR9WrSzsZQySGXlKCvBaysT6fjac2TcXzajdMzBV0CMv9Xq/8l+Xj5iALa
S5AUZbt9Ls8hvUcisNBoHA0c3r0kUZ1c0f4Ho6tiX8zedRzyAGjnbuKnFYGmVi08lAdJre+kvSgq
nGj3qaGAIPk1uKGZyOyPHiO9Xupzqlb+MsSKnOxNjuMxqp9cYaja1izmRoO5NFaNRP3lVtkfRRhu
ajZl448rNUoy/dcQl4Y3QvpiYQOUH4Zy0tFZ87qk5V/U5kb4EdFJAjjNnNwwQROaeE37jgT+9Viw
gsaGJhdnaVk0CBLw8FiwCf/4Uk2En0Vf23If36/UahB/d1ftjewJ0jP2sXTh98B+kV1QxkRzKs4G
eUBnokgVWy4WxPNVezuPOMd4MHoO6/mKIm0aLJ+KBp/8D5jK5NOXgBKafyFzYfcOT6uMjr9fY2Q0
RnSCSsXCsgXY+L30WCu+MGaJy5vBbCmdL6T4Pbld//fS00589gVI64706lEs6H/DAMdMaVNmS2TA
h4mi3jBTVzYV/Sn9zsX7Cy1XqwP+bTEPMqS4j1RN9fH/bAdtHlBbXhLzw6yCSME4AlYKUtc0f3fv
oIekdBsFNdcO2Fb/VQHgzoWJyy33U6ReAup9mEmxpAKmpxrWIP2Nq1+kT6UdP9MaTqABTZlgYp/y
WHECtvzeZrJ25hIdkdZXlaultTznWFPEaaB1E2ipnilEHdiUWXUIH4Q7/31rCi7P/RbQhLtzh6S0
MEYv+pgqI/MP15L277DxUS/S3Jv43yWvTMJzow7nIYY8epgfcPZQ+otScNXLzG7vEtNj7G2L9OFi
Pzp5qyMY4aNS+d8kzif/FoloQMmY6DQKqAofCEkjLs1LgExn9OTJzhmDoWaZq+2PWKt+SsDFI+54
93/QLfv8rZ56zXSWYO5T6Fhzr0j5WR0Aa5xX7Z1Ba4zsO6xhjQoPTtsoUcPaLufMQBlftJgZrQfV
JQCeA2wZdEXlJR4WYoMvQEm/iUWbew5akkSdNAQ9pJrkR+AWYTgnJbfgRtbuiKL9it4FgjOrUUh4
7gviiVwVEnDS5+H2baUCxkWXKtELCX4ZfIPboExUvZrynWv9so67zVH3/VlHsbIpOLabA6QXVQGC
GQZjj5eaHI17F+AoHmMQJ3cU+NKJ1L03zL84GnFQUjL6gb95O38Kih1uART7/gmUC1n4jZfoILxt
5g6Ng8qMa5KSlUDGbLcgHsTpV3DfTKHoO1ilHmjZMU9tEo20P6YCILDu8EeoNI2QkKcZJefcg/Ln
5DSxm1e3SyrnZ7QFXu8m9FTwuGplsZJxUXnHnypFCIIAstCTtljme8xGvkfXFzbldHRC6wzyRTni
sjp40muXAFTBmU61LYUgRmiT6+HU+Frr73+0CnVzCFcW4fFatxOCvyC1ZzTd2OZs2cue79u4FCfz
KMtxHmoajDuXock1Laji4xesnxwjiBDMpweSu2q1h1NL4IY7DcW2BKUVDIfuQ4t5FBoAKJE4Hqj+
63ogja4GsF9mYHT8miVGGxCTK5Vw5kc5YtaLnz00j1wqHuEKyUpCsFufF9wk70+kFQgmaTw8WwO6
4FFniI2D9wb4CAq77kJoxm0QtsR42EqLDUBaP8FdmvdT509CXNFMefGLlFsKonl93cuo5b27mMXN
kqg0gpFRPzIA+ZV3sW44WomtpCsoiI/NFlYLRkzIn97cDVauGzYoisHZ34tEIRLNaQ08kEDdh0Zw
pkcTIOX2iMdVu7MrCj7taA6oSaQaFJVhAmcOdS5LI5TxOekc1IuYgl4ooghEu94LxwWGxytL9yHU
MQBa/VcIxXVJRlDVE7S6DknSFQMztoxZWmQ6w5ccfLnbw++Uz+xynYBUOyJwDhfmoDrNMioZ1jKf
8qr8EkcsxNEQAqlqt+nJG5yYvMPXk3yzEEbRA3j/7nmFYshtUhEl6v/tCIG75T5gQ/DQNFMfZGKy
ewGsU7Wt4Rtz1C6MAem7Aa5/9Av7L3TyZX0hG0/w42PO5k+ddBsEH9BKe6+gCLYG9+UTzhqOc2TJ
iPcgIf6SqnQ9ukVmQxiTVqOMKUlfCWvsXUZvc/0SokzhujX6XgvACoBZzQdCPFVPMxp34979KQtu
/qmK1lZQmcSZXWEVlvVHSUAwz3aPxED4JVgEn5cOk5V8gXqYAD5IFFS4pp1pyUDhgt4bjDv5oVK2
DRE0/vd/LXnvOIcRAVsK8OobSTAKPww/4yKPyp2Qw1utY+VYlalRScmp8FCDDUdresacOkuy8e11
0JSJCIv7nNG83pey0q00fnspzCfZxtmcsCsEQrknjzpKPNbnyYkxnE74eL3ukkOvpKDlO0nmIdhJ
JdVhYh+uhaTr3S9Cw88XYsbMiZEK39GeYgm8V9j+lKrJfP3UxT1lOvfvh7b38PYo+119niT18JEJ
22YM5gxsVWf1PnQhzmk35OCY48FaOBDL+jQXO8XyDr3FgDW/AQl623OgPQGZClS0LXSDQoFtBHZI
K2okkrKXit0936evD/J0YANng60o59weyg5kmMS6U4ZYBydOKBZlwiWEvul9G3siOPBWtSUgQ21s
q9sUxkvF+0E+7qFjfoI0l6cNaQmOzqar/vvZfm4+BcT3HL3BQ6z7ozDK0mTEvp6x6E/omQwidLoF
P0qznd4f+RVsjlU1+1+xsL2BbLPrJ9o3O5hHkRj/ja+mH7hS9HZL5FqdLJAALhhO6JKQMHgAv+nH
AKq22z9ffwliz3H+42aocJlBWWonMueIKoQH3AFjwZARVQ9RbTkn1WpN3n8O8A+kxDcESPkeKKch
610eUMUCW/cPO1FCYDGMjVaALQdKelNlY7r0Luf2DqvNOr5W3cKv7eaMqZ1BPAqKoUOvggAjiW1z
giqMi9ubY1HJx5+7zXGi5bExNSD5AnyhNmjcNBNwjB2HXj7q0yvmabeilZu2kp3MF19BO0HQ3UJb
on32JseE+kI90BwsliTnng4PRal30cDHaOajUS9gF/5ww/sKp8pvRySETOz3O0x61FecDPvw8Pq7
3afBI8dr0MED0K2sZKlDnCdn3STaWA0FzaA2o5oXsqloehdYCz8BwdtRri8VLP3Y3xXa38U+fQEg
GLwttaA8zXqK6Y7e2TuIvVan3nM5HylDtrKI48SQXoIVAjjVTgv3QjnPUGIY1I2n34xce/7tCNb4
XtFWlq/B5uApBjSbBsSacwhliDUgmGvGIqGQcGvNaSR35C4w0DTI1IB+j2pW0x6UydJocRCMSaRX
zGp5MvVgQG3+KDNWnCYJhrH3ca9Us3jfY0/4El75VlJ5DIbaL+YWZ5J89UxRyv6ObJCzkST7xQIh
GbpYvE8tJA3i1+l04tLmb2QJkIykY0yRma2eWY9eQmJbQLw00e5SBkOisOiK2MzIqOu5MOfR2p8d
dOlpLBywpMquQZJbggyXSvpgHbsTxvTCUWdA4i2RzOTt3lxw0DUmfAaIAhL/7isVo6Zo9nFkYCS2
Hs+V7nSXMur3bn66ILxD8xbA47ASGpHE5VcrrtynLHJDQLrLpv0ftzsN5OpihXJNuCy9YU4VO2ow
zkMbd0rylV82EKryhO6DDEozSCa/B0QmGqshVmc/qPUrUp4eXdsanq+nQ911YRCKn/FGpDEEwhHK
tnYiEZ3es39wRwHwnYhGxh4rRA/hRndBBlcYtPLjovnecLsqH5e+yPnTLFhXSAm1rs6pcRgAQb9U
AxpjRkWqkblLsnyj9VkEP1mX8vSAP+Tk4ZZfEq8DmWSwpEy6u8Sb5fM9RX069mDDZ8fvijlwsq8Y
t0MVPcbs3RBcOypdqu0zpK6JK7rk+nE8+a7p8uT8k4p9HDk8VR5WcRb/gEK2Stc2hoywLB5FfCfw
fm4ZyhfYgQrkYU65ajKR+2Nr+EPIUt0SGeQ5P48WdUXDlC2zkuTxvpCsi60u/pVj8hUP8XdgB9kM
UYTP7T27k01k0rQ00wZ1Dcm0eyNdmGFF0Qd2iR89TV8sZomLx1NUHZx79kSYwQDtxGnuQu7Py2zz
mQNsXjeLoTSgNJuJtEOMQHIdethRSb/dIRsG5SXQlPxZaNJYaeZ567bRtCpdEcQvVxj2m8hDFPGh
MxTQuk4i1MbjEjvezdSwGyrJVJvTqfUN/RFKJxbh0IcKf27nIJzhvG0FDKB4+D0yT/I1VgyK2/d1
CYXaMPplRo7zaPxd56Z8ArWdGqe/352I87oM46fRaueD+oH/YG0fUAURU5Z/dtIK02LcXIx6+o3c
k9zc4fnE8E3bLCFCvCXU9vDTKJQ5FHP1YPZeyFdPCY+LMSAwSgk28so5g6X2rLSAoZDH+hoAxzcz
JFzGnEBP/IFCiZZL1UQRf/Jo4Ois+r5MziTutUv3/jkP2FJhJ8gYSk2HwC9x+W03qDT+2ZmMxQbj
lGwJfU7qa8gK0pQ/2wSUDadLMzM3JBo7JPHaef/6kMxCbBdSf1CIeEcnHf9EEf4K+k+8DgdsAr6/
fNjOKf82Z5AQ0YQTDe/DSwGduMOlS9TSA8uvm/1N/Ps3YMtDrc4j1Ls1Oyoo+wRVRAAIWSHwzcFV
OjUG9u4Ytwy/d0LAZyZuxbqEXSuDMiDoka6R7Z6oWrwo2pbaQwvs4eWUb2T8knOdFLXfnQIZbgWt
S+xz3kT8yH/MiIN4TyAMWMKBVTtyYmVj+40IpupOQtpH+rt4VxiOjeYinconBLsb8KStr/uPr1S5
KRK5/MlwLGtim6djzMDI+5XoBcfBFOiEE0UTAvYu69Ib5B5TPeW6wN4RVeEOmDeNky+CEaB1RD48
SYVOStMhUf1S1V5ofc/h8zMRzJueGEA3MJc2YIrvyPsibXX72dfyMDw1W9VHawC5S93L9tvA1YW3
M83AbvpoPDXTiBvYMksR7v+Ye5KRYey3bz3FUIdNxsCHzkMMzZg4o1lEfOFhCIYJhheCIERbLIGq
9i1JF2qiLEbXdO9R8pXDtF+JHd9QskK1ov3cv6c9Y87DR5SY0TmS8g7C7M4dSVopd1OnEUZKG0f/
RZAWv2KxNeICOBWIntQEodsOMWpnM24Hv9t5za4t9U0EsJIlYLbDhjsfsVlWAOTD042vfzMx8iay
OqYMeUCWdC8fCLMyx8DCIjSkUPIvgG6KurYJzwgfaUXPzUpqeViXT3EsSf6pqo/rOwmPxblWtlLC
36xlgWBUjRWOuvKwjmhH2hSamZr4xgd1XPPS1dFV8viuhwt2SwDUNB6n4j3a3rwIjh04DUtVDX29
GxaioTn79Ng1DmZPR54Vp5PqiYe7wBYZcZWnwPmuob8DkSyqT+UPoT/tvW701dtx4opByE0sOcOc
9px0dQim5sEGsFxisq9NtYXq6MpFS7Z9/GQB1TiTTor9SJIJX8+0SWyQL1pyWIUBCb0XorUmvzuz
rCOtAeW8/Ey7y6wMYBgsEhQjKYnXrnlfgmLzxHG3a8fT2Bxtd9x4lDUUe96UYBWZlcnaEoPZCvza
e2n2VYCkXRmPJoSqYKzLTwjRJPJeo85gh7G6RSnJu96nl88w3svthh+RI4eh9NeiW932JE9FYnUn
1Ve6EDoGQBTTVrgImS23tdhFiiiJ/o6yoo9otMK35gOv0+V9f+xUCV4BY6hK7/+7RcUHNhUPIDyt
qOWj7nHzWZdC8L69na7xMDJ7fU6Dj/ZxnB3tJ7x5QMvfaR7hUdwDSA/+fNmDUA+R7dWHueKyCrFQ
wEVvLVyH7REwGXF3KxUkysks6S/ORR8JwuBuhvfj/ceU1IJ75B4kfMxT+E7f8gV33WfcrOFVsrYL
R54XyTPQ8aIuaX2JVIvcyDBMNKzP9E8Xy0SL6Vc32LsGIQ3ox8pS/7y00kM2cZtBFRUzdiAnakFO
0uUyOA3SiZOWoHmDELJzi7dvidPjHpQ9dqQ2ZInWkJ2ChFAQOsPuSTHAaGlhHJ9Tc0AculqGPN3f
pp0JJE6+hPYjLII+HwbLyani97MRyo/sWAMh6ZAfTvrR1B6IeevNqLdVKeTfSQuKTEVPoQ+RXJ4R
y7a0o/KOcECh7b5B/YvXdkYDAM41mDeY6MzLWIEf+4dW/siYaiWY9bvEnA9cB0ngDUP5fZcY03LQ
uIWwPguSbNqH4tULcFtXk5mHIYjGM6rN2Qm0rSnGlKNeRNDSOMGi1DoFOaKy+19lzXiczGepwNaq
KOi74EAGNXE3xAMzM4j6RLV1NLSzU5JbWJG3X/dhqXIIgFh8a2orzGeDUBWvOdSvlkJ+6HJ+v3Rc
c8Kr6q+kd3cM3uEJzPa8/t24Y/IASaDWXTDGGU4bBmY61K5koyRC9ri/Pfp3ncltree9IqxnIRG5
q/YZwMg/6MO3Im3gWQsG7SReqCSpfzRJdUQeWduJgIdYkAlqFmKDIgKH0chdmebM0i0QRJFavdZT
/6fdpSVrNuR9hsDENRYrxfTQtehV6AR+UD0SVRoLw4XjY66Tgp2kFbQJeD7N0WiQTS4ZsFIBDmtM
MxNJxcZI0FyQrdmD3WXj0P+9N0L0+CwP5IXnc4mxjpCNCU3RZdjaU4G1OC33wngLYE46sXVnl9GN
rfTUbDjsokG0UKN+E8Qsg9W9jqNeBqKC7IkamWYOT03j/XMIvNnPN3hW+dqhh5W1csJ02/EGQY9Y
krLIB+r/rPsLYHpozyyKOeMXGNX8TAJtN78WK5WfTbFbW74f+qwX8wV+UnrtqOgavI2ovigsnKTm
pRTnH484uWqnv8ylEQNVUclKo+by04R/p4wsmg9J02EThwG9txpEUicBACWXuh5qwJqzC1FZUY/D
h4RL2IEqH03/ENrCBEEPNRcTOjd+dwQlLxprNxzqka6bP/fPD8fzf30bWSD+SIrmoZmfqE6+A6dC
AJO9Bpz4XUvaQS7SbgomkFd/TOLgWxQyEtFsdVqTZnKzhimymRNsyXtoYupI8gbIWs/XjV8c5iHT
qa4CKTAeAQjcfHG8hCzEld+kaTNjJJHb8JOZgp+tO7qqbcarQOonlCC8UNTfIoY6vrja5m1JQjY0
/GUUyJ6kihfAhZ1ilUqt0iYU/gwp0hWTqSTP0UvFGr4jOFC+x5GsIm7AM9wSPRUUOaiZ0RO1LO8N
vVhk27lUSPMSVR/xKBE/vxdqLwd6mWgGePrQBK/BCtSRdY/MLlvkKWniymt+Dn+URkBzSg65a3td
ywAiBHegcGfdQ+WjtuzFhojNfzobwR+269ictFh1YUASBWjC/T7SpFbL8k314taT9C53FetG/4ta
tNBI04FUeerb5uU0ojGGmT5+JULlToxMHKQFpKzMhEdWH4Tl1efXaP7+TVpJv/IQnLzhFR0uCCQr
Xn+LeUEPakEL+k/Y8B9/cI/HHSek2tWeuAN9x7ZpvRXIKYKE4NFwZYPyOo2fDRS6CnsR01CqP8OG
HoAHL54txTXf8Xc+ySEI2JqwmP5rkPMMoTdHovtfNw2JzcpCb2Hhyuw4FzZRSVVnKzgFs3NADsmg
yvEkkxQqgg7q0Ufv7kTAwOZVwp6xDaMPTV89eq17srZq4ZcCIkT6bS/kl2aeCRKuL+v8XkWKIppL
TZ/0o+oifL4yYTp/wYukG0GH8zQW3V22DTBDFrS/scrOfRfBbdTo+J33MVvf+PKbGOVZZ0/1YSXe
s3bwl38RCF3GjBhZNpnp2H4XC5BYs3agLUPe5pb/hy/5o9itfiFHm+xsq8mhDELIXgMBO4ntXGw+
cacK/w0fi0G3UgAnKZUXiT1BKQ53C8IB0F/yph0EUMqAMXJ7v+uKTVyJoPV2VS03xhtQWVd2cOoX
o45WATQhmEOUYUM07yrZU1ptii+48xN2PYh+t2nqypegXREVwGRh5exS840jtrUasJKnSh5ZBwbO
8nUDKasTsTSSOMdDtWG+3NZ9NGeajO4JUpPi9QQHC+YwG2evGOaK3QG2PnNiPC8KqGokbdTS1HQb
3g0YLMLQcOTQO/VenUHqc/CCfApkwsHD9RWP2HcNgpdw2/ICBeAA+gyjz8F3Oz8cCpY0wU7nsf+v
k7faw8x108mKRhwjaZsqqsSofLt/LNCsKxF1GIuq34lsKWK1grZskWJjRqioojOxWvAb0CM1GTPN
SrM7SMXbmwfPPgei6LtiV95WYZYPs8LK2ko58ST+iV2rufxEnYg3iRa6oVQ5UUel6PjoRo6s9i+o
WDGAJMjQ4Y5JqaVQEdPag6f4LBbp+/hE3Nzw3pUfg90WkQdDFdQ9OTT3pHZv4tY6BU7kuItOUPE+
fY9BfNrRx8peeSsd3CwUyg986g6Ze2xt7vDBEHdpyC6mIweERtvob5AJon3s6Mm01YRXbh8GEWyP
In8zeS7SJXZFKKemgDS1jYMSghbLcmmx9HgbDhJTXPuSJw+LYQ3aYkVr3E8Yt7KQOI7DIHPEN4gD
EoqL22vM0yFawFIxAc8c3dhWExanRWYJ4q3Uk5CFpmEJa81U6SDGbHWn3hAtFkH4K5WvP/MZ1mr1
Eju/MXDBoX3sLVObBIe4pWxwc206/KoSuGypTf7Dhed4lDYleFtTULMkq7R9xhboLsN6CrQBX1Jr
VgbYWRqcvcC70U/oS4ZyC44puJ2J3mEtpqgcVQwcfuC6PBW+uRRh1cM0qxNyvgTxRToH1pdACjaB
hwDeRLVgcJN3jdOCS9ZmDz0WfjElU/KWzvS4f0VA8+jbce9fsuYx3WB0FzLwNobfCiDiTfZ7SWy1
dnqQ8LQOEmGGr9/cazrTSdA+eO575fZlPBFjFPKJ5lLckZSBOX6DzAQYyLj7zbB3jm2hUU8kqzp+
R/m/q0YRpY/1QM+e3i7LyfDlgPk9KKVR2/bZ2DfDekXQ87s+hB6ubFT3pn04nFEzbF/RQ9sKob8n
CCXpf9zXWXZh7773gAe9rfNKFdjKNYqBsg+yG8b44eB1OVhPilkKNK2QGDXoth5aN4NT4HOU9pRw
Xff7fk9p5StgIDTfSmfB+2tQO7E/zfkp9URSsJbzMnt+sscX4OJoqkmSCauTCItwPABo0tAlKK0k
YwrcSOaaqGsOhmWOrdkKs2IqF3N/l7tcaD2W+OSMvIHCl45nIyOsCH6vGK+LM7O2JS2A8k5La2iN
4pqw9JZcilObXjQ39dPR1jJX9yBWkU05kXv0Enab3lBhbK6kkqaAVsrrq3Ku9J1F19ozelBz6+cp
RUvUe0GAWgXJuMMoFp8+98yyCM9keI101b0KgYc54Zhkr93+MLcfL3NEuJ3FbNlSiSdLBpBYaPhU
dVmaVx4c7+g0DzNK0CF9E1tfHw4EZ4sZuQB+c9kKCN9EwrNwEKFv1HlFcGkcgBMlykmYgo+rlBrp
NfDTixN9jolSsTE9FTwv21/RtSx/kNHC0AqQhNHBslZEE3LdA8gDY3WPsLfLfaedFUyc1ZvcAwE9
dgAiFpPd3OFvORTDMHcM+51rBGDizTiunLvmZm9u0jHP/yW5s/S5li2m6nPb4Czzj4h4jlR2ZUMq
8JGJ4mqBWK1oGbzMt6vCFr2rrIR4+MKDCFFLI0USF26WpJKchX6/b5xKZAyDsq0XqbLu+WUCKpHM
ZuY7WUONLKlGpIgZ+1tTjWK6SvKz2QrZUWCDIyXFZuC3etL+gP1ge9Z7f2XFLnxzHlFRAkXhAXp9
YDrMZRcpQ2jPo48aReK7bVo4e/zmO0jy69HxHrRfDdOvbRve4V4vVYtQ6cGWPrsmgsU3Fwz4onEZ
SbGX1IUGkskU0yPA0dHvrgpKtC/5aL/BSCFQNyvOZ/Se6nMD1hVy+9J/aBZmcmZrgr0w11zNuSFU
2X/PSfLeaFZRRwdyCvwL0l9WiN1yzmQRRRC+xlDGdwDI4ZLew+pTokpPkvi5axQQVqIDNwqp+kYb
s4e/tj8uktDgAZQN8IFbjiN8N0QBQU/ERc8iDCs+rPv2hwSduSFwYNigiE0wiVHJpanJ3fNfzMpp
5RloQtiZGwcPjlfePlXQma+ODSG9C9rKLzarFT7sSpCqLDPLId0Nbhp8lJy2ArvZXsoPEi6o6WLF
SB3EXq6ET0rUGdsLvGK6r8rLyDP1i/bznImUFyqRHuTQ325mYDe3L+CHTHI/AhNwgR+rKpMcvkQT
rsef7OvKkOsRIXWQw2yd1/R0Rgha7xoGnrotBN1XU6CVhuZNnJCNVIYLhTIaU518NJB8R8yEGRSE
d/L2clppAMQ90X6D2L9KWzQf27cwh1GFlmq0YEmb1rr2t/b9kFeXWdRd5OUXTgWydJL3XLVXGPYm
9l/oltK8CHsuO0vI9DiaMu9Z860K00fcBJvqapPEWAEiK7uRQVxhvDazSyf8D71m9GeeO0r/8N1s
W6L4KThoWZzaRQIJUBJmTkBPtQwIbFd3GAICjXx8h8NQpE75RyvT+nAgQeLqsLi6FWHByvpuMMLi
RNY5XDP2TW8lQjle8/qS93fLE2XluYFOE3lC7ct497cmWtuakqrK7kWHweBIyNtI2lbyBIhvP6BS
oGSPCH1u/SNsJvXoaEcCWmWg54orbV62mrmbldNZVMB7qFvqSn5Yg1+M+Atak1nqBMgNqQb7CZ0L
1N9TsQYbr+OfBqzXYmL1KxvILNYyhGm/0v80LLMpwmW239sXEiltU33VksMkC+k7iGfhNxsi8bfV
h+jsZ9902dFxTLr26VCstb7YpXatOIrXFlpdEb1pxG9bg4yki1fGx6MkRUekbDmir97QmZ7A9BP/
E6By9g6GhNeodJmPv8Ox8/30ZjVUqLIVE8HcPtMkiD0OX+J7bfje3qSlykLmJh5DXZZ1VuckOlM7
xinTyE9XNb8W4P13DedyCLkc7QFHUOksPy2/NrLLso+y0NH6GCpYvrxeoEKOfLk5bLKyfjFRIS2p
kk5AifO/5m3eGHHLiuOaoA1Rkdf+lWV3MFSW9Blq3CTgJHjQXS/i61gXUpQfhEvNzbpndmKZa/su
HrUHJBSZ4XSfKlRonAgQJ00nT20102nm/8iVBPytbkf5MvVIjB3KGGyMBofxYzafLWO6YWh7yfIj
TIzAQMr9k/NSI7XGSa2ybSuC+kw6OOxrEgINoG/HSqb3K6kSPJyE8qwVVqybJPlEJjsgG/1lReP9
PvcchfJspAKK+HadqoioyQwJd6DYQk58v9n67isiXsMeTyfzOhsO03HPskiqfkPCgPSBGREmRZAb
bCm+sshupFjW315kjnHnKRm/FV5l3VRbCtB+geaHXM/RB5E9OKyZkDS6rYUTfjmkX4YlKB4unxkg
qfH0biqIuxAoMuLZhYUEllGqepS7iIwYWfDbXyLqvHZ1L3SURwPiyC0dkMVCxQtwukf5mxqwfhrE
MLjW7qdiOY/piNS/gSIwymLUvKuygWpsDk8Df0L8WD2OGPN9Qd98TLI3qWcpY+tmbK66t+tuDWPB
70xwQAaf6bVU8c+R2mKx1ZamjsZkUobQknVIw6QYiHlXHDI4GkArvl0u+J4BfwfP2y30OZpafXEK
cVl6uUBI1Pl0CB9r3Xez/ku+sZHVnFz6cm5SuJFIvqSG/pA1drrm/jrcU6h5o1ozo3Rpfvn2/+av
4lsc5OUp6Z2IL74vSZQpYZ3Mfidb55KsMGRTWsp1lOOzrjC/9wCHY7M1n2KZHo/c5DoHTPW40z+T
Ll1Bp3inwBFh+0itMaXhfnAU4N09GN/bYM6thMShdSow9LIrwNVeEM2+DYED/WMDFqPu5Th1SzDz
ec0v3rRa0y+UIMnjQaS3geYoOvCxhbVf4IHiS8x8/1MP4iEiHn56rjKlyV1rEt6ab9TZI7RKKqsj
GHu+eibpgXxeOeF174XEyCB1L22LAFqZDp7cKWiZ0z0sPzCvdQGgRsUJrWOqjWrorXYX6tpw7obK
nYTGGqncYYnB+mPWg3Ln5wQdoSo0CnnpLTu2IRI/sHi/lh/vBwyJGtFcs3jzGAAdOZeIj+6LcQ+j
/YLRlpRTbdKs7CRHZuZdJWfmz5OyMnBN9SKncbw3K7GEHXwfYSjojgliEBqzN4LgsDI4qRJfwEid
ZeW+XEPAYtl40Pv2CMS/ys/AS5i7v3OrQjCKtffTf6xWWgVGn7zLSa66qjTj2o8ERplPVjAtRB73
CVkFiZEsAUSQvsDLku1bt72sZ2Eka4VbxhqYBlVyYZDPc5ou3Rs9xXjpSY/kX6iocMBSCN1lnMDR
+Zvpkg9c2Rc81UFIHz13G+EnvOyRfCJ6szOsH33OE6y72xEuhOoTWSvxdavQ1Il8t7I/NQ4rZiBL
rH+GMWnukw8TyVs3ozTp4KTvU6s9mPRS3TGCJ0PdFj62nGlIHrocCONVPpSOkEW8Y289YHN+JKao
frBkSW8cLBZtOWfZgkHaOD1U2OjMuQz/iYErGnHNy6rvdBh+FOxQ2IPA0P/830qwoat7x2ySLjU4
FHSYjpEKY9e90Xa7uOd5L3MpFYjKPWqh1nJs/oYdGUHt0vd7ax43gkgk2rTfCUthIaybfVPl8yst
7+YOWjsIVc2fafcVpNVYWXuSvjqb3VB1fPKfbZHDgNrf/chG+T8aGFkuxQT4h6X76LtIJi603kk0
aLlPEu0sdbCRhDtXlM9d7R/h0jXKbACnUudQ1Ry9ynW1UjsVfMhSlsfuCT9X6TncBcrSaUjPA2LT
duyz6QLz/WbBlGKm7WBlBWIdJGg7LkqZsNITM8tVeT4sFyN9mNclMl3NOE9EJVAcQyn49CRsA6zl
qEz/ff4Xo6ymmTLNrSei1M+tOSZCRi2J20S+h8Gq7r8KEX/jsIqiq/IMIwTyEUnZqI/R3qWlm1v+
VcHX1xqdXb7UIk/lb6tsX6RLkwjY3MYjH7mE9asCuFs0WWQ+R6GCjRQ9lU+vsRdlae3Zt/zXoi9g
EN+Pvwjw1No+NlN6rVQtJma71B5am27WAivhzcUPopTkThWS0odkATC9OM7ng55H97XdmeaL3nBZ
2in1g7oAnFn4G3MkBDwrsZPY+3/bRHDHAQBAxy5M7M3K4R+cdsLRTBmR3cDUYqXziNgwBoYhrmaO
NVGOm7W+uZ1VWQ4yY1E455c6g4QU0ZypvTMQMLD1bhOFBYkjrp3tNmHh8inSHhhNF6Q6gVnOxCX0
Lhn0vswnFsBowAVSfv8b2i4U/2mcLKk7omdRmdKeN+UJN+r0H9dvv2QWxjmWc1FED0aGKaYq/hfU
ceUu2E2PxhZ7msiZYIS0914BYtdi/Cp+LSJ7M4bBq6U9ntwACSRhVq3ESNNkn3e4Rz8MJ2eYhaVJ
oPCCc5VFu8c7Pqg5siI08/YPceKn1vfaUDJOLCrgL7W9HRcrvW8aGEKFedRT/oUg3wUj3uzMIAMg
J4+AD6ZMtFNzFcdh6bu17URZ8OEkc4MeQx6ElU1CZrl5ToY1Hqueyisup8bpL3zWcEP99beVu9ET
uDrGbBXl5HQT6HfBlsyPXelP0Om2783w0gEVDRQb5UzPyh04F0v4Om7MHTyKCWuBhJHxE2xOvAiI
0qOepkS4c7kWKAXaAtdrAf2ueftXNRqnfx0soc62yUepoEDo+zDL7M+hCChY+YdVKfbwN4D0FXHI
UTkxgPSgxYEbFizBvik48HgZJ2ivqe/nyD0QYfua1QTQh+LrhzK3Fk4I8DWVMvhaF0xCZaSwWJWK
JTSRPDLEHGmxlifDtdFzl3/DoUbZiL50tKLqRUcMzvtZxWHp2LO1yf1ncUtifjP80kBb27mMKaKz
DDKN4lW8AY8b88AktBS9HHZPnz1Uzo8ug3YwX5RyLBwI0yjsq3jccznryctxS3F/K6zZJKqfkPiC
E4Mz7iSlFVSeEQjV+z7UyuovEGwVoZ9wEq4iGXn8B7Yvpckwenl2D+TC6bRhaxaYDF+GzJXXrJGa
Ti96Vry0+dhuVEn93cm9hQF+nC4TBmr93jXrni+vI9iGWgdN4UEtuYqj9q1geH6kulRKsXUWrOeg
KGCVBv4rN+uXu8qfPnk1JOWcNelu3HJzQAV4Uy/78XvznajTUFu+6DV1LKUQAp3Sn91t6tZcYXxi
lrdAShktdyJJe3VjQ3smL/P0oCxrvD2XYyn5uBfnoz15lna2KvUOL1T4qhq2oSlwBEXr332guK7L
7ZhuyDKGCUjV18ndksA5QTITNNkolPi2JnULGKPMPDOFp7q0K8Ce3VHNEGjXGrWDia88liA9Y+BZ
Pbv62Gw2geF0I4/cfy1zW2+/xcX/V78kE5m32x/Ur/OX7E19PChYLCO/rySZ/RLHY08GPAR1Sq+U
rZICpCnAYnO6PtCd1hMoHA8QDbkEJK5rp11d9A3zfvAx7rgC4+7PWv+Sdx6mPUAb4+X4g1BVksLE
9WWLNwDLbWxNrtoV33sF5Lj2eduP5ApVEDH3SPLDpRY70iZYEcRanUyq3H/1AGCcYkIU3bkt4psA
dEhPT7BWNe8th6Q6gIKddOdHmM19eg0Kyx1PL+7y7pIcHZITajZsBUMULQ2p7qHiLNH6FAR8UxZX
8dbONYsBT9469PezXPIcaOxMS+lw9C3PRYEjLuEv+UaifjdUDmjB2LbxVZ8HQNM3caEYFLob26AV
2ajW3gC24xiJyFwKayR4e5YzfazVOVfdl2+6vpGJxcRo1gm3d2Trf8iPOb2ik5RMa0jjP28ZyOeb
BCCWBt6HRln0JRUJkvhdQBQ2ht+f5YcoDPUUs0ieRoq7xfHaIq6VeQ/HNkyMWwZzbWp9liZvxckL
Mf5RNzdfGmO32egBzb0cie2tkXam1j35y1CaLc0glZscOud1XujINtslVZBOYyisLMoeBNkIefGH
/VvFEkTDLf0ANb+4+zTfCOkbdkOs/dZHaMwQbyMD7MmWPG0Rky7cknktGGKaSs/MlQwSQx1auWxp
pDFbMAnWTXnJwKoiCmfJQLK0KodD9BEbCOceiwVBCnxL9T5BnGVYcp7fcvLpvfSMJYT4cRddVX49
fYM7HYy2codnb+cX3ctyaPpixMaIsywaZcxX+nBVUFIdwkdmvdu9/i8dbLYGakj6semsOsahs8hV
I1zjKCvMGsQDpwSFS8+q7DEB5h02Qa/lU02EqyuS+NQBODHUKGu8UC3cqMjR55qiiL/YZDA5Bl3b
82IQeVdZf9+ocRwcTrLe+/mt7j/jpsL3S6IOWaOMHEnDqhogjpdSKbkA6U9aKfInhWgoBO+tjuQp
RzhNHvMOMUV6B99upUPy8naCpCUBxruo5KoFK7nEI25Gi5asllee318bgR3RHTjWq0GM0VSR1k7D
Uz9rC6xEAEycrzAMpSLA8y46DGyE5v+daEFyWgnQEMCgajWak6GZjvOUZaPSysmRDCnDxH0U1cob
Cb8M3FUqaRplOB8bWi/Za7prFGnLCn4/SxmBk3KbYsi4ShS5Q5+mSzAGIj6aqagUb6uo5jfIViNF
20DDXuD4/jf7Ef29RsIryUdCCmPpK9YeDvBIV9KoLHI7a/QpzsotstlhKInqXMJjr8tB7W35cGKs
6/STTLNHgl0U1ps8E3b4lFjAUri7MujCLBbRUWMm04jnVkQBZvRiHgsGbRimc8l7KXFxaWVUH1EH
TuaINKbSdvIRI30h/UZFFHwNWVRHzmkjJoZTg/L1b+DDUM8wktHMwE6T10BoYz+e2RmU6ba/yCVX
WO+eM03CqSGPx2+LngCeN6oCUEmeCYnuadUy1SpDC6a3Fz/gUNBnHYjU03k43BO3Y33UGKWWAhop
jfu2BovP2yRtRjJT/Bhoivui/dwM9U/onldudauGB29TNaERTcN026CQDXc2PKjXRM3JBC1XBUov
iAYk5XGDZhRTLL2YR4nP5q8HQ3cPYtsiDh2W1Z5XWTUEKrS1bCrycsQ6Qhw8WsN5hyPNasjH3ZDJ
JLkwmpTYZEeqmyoeCiqzME9+3YBuHltpBJDj8/+axvT021qreBhMI1h9XZa7LhS8rWoNCCGeqtSK
k8ObCL6IpxIIoVMJZPgz4fV7j80WsACHd5QAO0rwn+hqXPLm0ckvUoWwGvNcMRhAytpBwf/jWtCL
hcLFyuhCtSoPjEpBO0zlh4VQ/9UF2xykWtrPewLgUNKYARZ8OG6cNwQjp+u9cSIQRpvAGi99NDSM
j639yG/AS7MaBnMemfywJNLV6agNY6VjvjbcY/CP8ACbbkTocbMXCYJ5qIM90ftYzydShmxzMd5s
z16hFoZiwnp5dRRYdulU9ulWsa8+mGbhhRJ9FapaJ5nrdtClE9bH3FiyZH46XnHFN50yhcR+PEGC
F7s9aIqeNE72LCAM7pKglv8+l240O5HbVXb1KhoM+6ePHvZPMLYQIYX3EnNTYi5Z4Lq/OTUkTzay
oiR9Z/5y8F+hJykABysoTxaxydQHjNqDy4g901QD4bKuDhHIwL6mW93VN3azZOokFf61cOhzZdsr
bHO1JGOX9X9KXxQ7HAC3NbJhrDP+9UURyMxR+1iNsZ2OZJRPsKv0k1dqacJz0E8tfy6yZzidWw8P
xTMtG6fLO0Bf5Eiubk9RrJuQyaL8vDQ3HdxMj9YU+Lr4Z5Vgde5l0aZ/JfU1cMp99oGtI0dnrS2s
hwyz0PVZO/6VcKA/SaBxW35YV/LI1Q2g9KcgKWiINnNI2oWPUZ58ShxqJvwldCn+vtT9P445ylEM
ITn1+1nsHixAgpKeZg7aui3vNIp4f+wj3lAryi+A7tKA2k6vZp9ER75GNpP/PwesfZVDvxMp6IyT
4MgnPbX6uEXssGx0E3yEmZf7a5I5pz6wLaolFVqcK2rhQ6ULEAUg3PPfQIoPVbjAmUjAD/wyfZOL
wNrABiidjzy9zZ8Bi5YemIXED5Hoh1vDelqihaI8xP2UmHFahhUNuH8EYHjfzup48yZYUkg1+8Bx
IyTc3XztOwln3dFp5py/BysCQtU1OVdPPANLZg37r+V8eJsrsJnb3/r5lCjf+X1CruKntZ4wvLh6
MNrfGfGIjRgz5T4ctryPh483PePQdP6nWtI+5RygOEb61jAFg4lR6Xo+DLdYcX1TCPVH6E8aNq6x
tJOkusbkca0lItV1MqgJwRgiuppkIcCOcQKhYYua8xwoFY4RVd2nPFaRrPwqHEj8pLUTDyBrAqzW
s0TnX03nuGvEME3Swjql1Ptp0IMMy4QL2NGXBEp9tjdzNMMAHMvdB5lhgHut+j8020f3lJPWv2qt
xWEbPf+PdQRVZtC+S4PPZ3BdtbSH5z03cy8v+FVGH4bwXncXnJ//l73VnucaEmhHui4Oi2NQS1W6
hcKKP5rmSikZaevAE2yDoSo+Asd7EdB4l2OnGFDBfh+cS1kdVOr+cYjc6RUBC2uwS7vfXrx2eSKZ
d1CJvfJTWCcYEmaHCjnymZdC+tPKxqOenfa1ueJvjE5OHjnKTQG/8vkKSR95l93ssqwKhT2Gqa3J
OltMUbIzSTMwD7uJqkuUoxsFMaD7ikyUEMzLjMz4sPyLHmgrn9TeI/QgdDewnPQk89Z11GiRvuKI
NCAy1hyqjg8OdLoNASWO0iBh2+6tzf36STOAVDpN05JhC2FXeVrqnLgNiNnihKiZN4VSBooHFs1W
cYYNUCj3R10UVqNejQE7YbgtNaUDlwVw9gsuQFh+jsp4BYHAT1F259j6lQg+lftKDHewcXMYVZVS
ZlPxSwSYoVRR/RLerU0wZc8/0kOqfYLGcuwx6F0zHO0wP15w46kp4MzWcgKApjgWzsZrd7n+2ZfM
6mMB+ryVI6FajC2DKwY4vibyaVik5KUvL4g8quc46L8GLk3Kf+vV2XJzV9z/tHDUuc2hTY6amw2D
0Z0iw6RZkN7Rbl2IAc1Xsakw5WjSBPAoGa8TZky7a1M3Ydv065GlB2Q3O85O2/KpaN9TVfY8Asyl
arVS7P4e80RAOsQnT5GFAyNWfr5hqQXURJ/mkUgYSgXl8XskGpl8ZFLtSShNxpgu+CHfkveqUb6F
GeekzIuItDDqG3Ifg/zf3BwVMVbLtgOxns6YJp+xvD7b1quBWOuBNzzgVx1eE/oHO09NFlLggasl
o5m68JV7vp1up8gxZhDjGtnZDx5+er05jH3vh4bDV9l/lshiYLU/6cvOt41yMoy1IY1SteoCPy0y
hh0QQjuIzSgs1qRF/R+ZWu0krCuuw0XO18/nU7kuubix20tqUlC125DEgnp/LM+DLdj4+tVkemjt
nMW/4c2AQ1lh5h0T3t7JLkVkr9zJRJtUqjBDdpknzuFzq9PiTvHehoR4H0UGTmEqcaGmykLaDBTY
0GOFBs7fdROUCA8V9iGy1fBn2TYF2BCYplInhV/s+spdIMawWhpRn9dvSp4o1nUlJV7plcOuWQPc
Hcr6T9pGJkQ+hHF+/q8tJbYshm2k2/U+vkPGxeD5Xukksrdoczy+Ns8ipmCtgQ9rn34uDgjBMcD1
Gney8Y+yJz8Ja9MTJO2sh9KrHvC8bxdIjfQQptzr1UW0Jn8b+bxVz2VQCi/W1lmae10c8fdMSL/I
VafmzcZhLMtvFGlSKZ6mc/bkwDPn5d7WFzwIYKE5hZ9F4Nbxn+zI11000ugz3sp46tPCDOEPAZg+
DY4daiMPPh/kDsTwZ+8nD2M9HJKh7XfESQLD+IYo04doJ+6EvF2nk80EJGY5KQL8qkMUj6FmVVBf
cO9n2/fPZtWwHJEgaN1KoPJmCdBJc1awdEP32N9EmjbSpjiU6WKfyZaoEEmzK/1cdsPxmAo2QPtz
3FEerXzYegM2mosDpDrLQ4/qH6n0YXBLVbAwAlvF0CZZzKCSJLgIQDX57ioxA2McHG7Urin4xAKQ
uGKRPPAjoIV0/84sDXYnhmjVd9vAGSApTZcm+qb880AjVzcbVYKgj09xJAMJV0NCDeOfwRj2FJhI
eX+q8GdVpM/1iPgR5Je1BWcN+OKvdH46Qb0/Prq+QDJjr2Q1h1JUzV8nXXW9KB+nd+Hwy5RVydMN
QgxyGVMvhFGeJhKJtpqp7D6BMQtYatXo8o8Q8un2TngmS12iw9hXIlsuuB7OngirSEBn0w8kgXwh
k8P6a+KD18J6bBQDXwrhxwiYRTa/aSESWcl4tXyHIR6Vpnbp43SSuRN5Z5jUnlJARNqk8OBsWO9w
rcQf4uIppDqrUKWR0panjd+SyNy2trtmoZpDwLgaHvVQ4LO4EvpIB5UfT4KL4nkk0Iuy1z1FJIdm
ka22SMnJNkkswF7VMzNXysXeyz2y3tySvfHzZ8WHLyg/6a20vqUcN7l5xlVBkYPyaze4Sw9TXp1L
/6OjxdnGrnQTlXZnLVn+bzr5wC8Cf4PaKyd7t77ksa7S4FaY7JIsmiFfBk6qd9BJ0PnOBMCvj4d8
Ev08DUSwKj6Y+wLMr4/TCJO6OdssuRFlABQ4vuR/1IoP3VkdfCuUKfaPr1x1FjXF7/X+l126Ba38
kiMJWe9A5hYY4i6tvPcSuvEb3eZ6TUzDu5fUNtLHELmO8biLtAZiF5aXFKJ2ftY/oXYZkg6JQBzq
6wYwLVls8nBHfh0PUYTodkF6YbqmVTaiaeu1EwDLHsyUkYJFEw8QCMcplo6LKD1h8YRk+Tpl+b6K
9b8Hzi8fJ8E2QqlHfqy1V1Squ/dr1su0Kbb6gAKFRG21TLXkRPQBDCanfOvDanZF2hvQlDNxKd8N
YF6fRIm8EBSGBDno4NzC35xf7ysPKUQ5royV8enJHK8c+HdpIpYsmNKGbaNfGDZba/ncDUI3FUdT
vxI6wokCtUj9b72By6CBPGhX3tRtGrWYiVDZVkjDxU4DMy7FsSI8fQPxe3+/VmeUnivsI1/fwED7
4pZNkJzIMimr4YkHjdyzu6KaFt+A2RLlaImviWElaijl1x9C4JVB4EkQbZChH0NTegCqmHkJZrkX
CGW6FzKBybG+OLQc93bzDCpYRU2POwTbhqqn9QgRnRyA9u9K2DRl+NYwu9OgT22FemxDmUpjoTE9
4FpcsKT0I4fJKfhar1qmgwY/1PEZs5qOs8AQm6jSmTksScykFPIAnpSdKE0YJMUPztIRrChDFlvO
Hd3bGdJdBOSsGRrRFVcFU7HZCEnwFa5Jc+gdNnsR/lF01vlVd+KhLngO7Kivm34NTDW0yA3FhNfG
uT/gFr9NgLBiDH3T98/35ikeqDezLwqTa2DfiSaNCvgvomYMuPb99LN7eJ5BmXTkj9Q2XeXCG4cw
6u/jHcBbQrb3IWhvZKjUU2EPZgxPPcrRd+JghxqavgAhjoeDP6flqhMmOXZjUOZr/wuIlqN/aKZQ
SlQDw++er9ZFvD6V2TO1qlXKaCM5L7VFzOav/4FNiqrnXjZWRf+NpQvLl3Ky8fwfERO3lPSwUcR5
gMFgn4Y27KXSb1kCRQKyalD7KJsyJC93HlOXX6uZvOTRA8SuoNlejJjLmxa34reacMboX5av6Vxh
Anpyd+TeL+U9O8f9syhDXohCm7H7lxPAMt0zjSWUNDlxbCahrWD/XFf7fKIrOxKErKTInJ/+Q8t2
oBI8mdce/+KLAEBboQkigtq06oQRNeSVPTvPDm55CqxnQ4O9ok4D6b4i5omTRfd+wFcGRfxqW398
EuCIgJmkHARud4mrB3KXuM9er4Z7h/gk64BitNMwuptk2S9hFKqiflkJR+lcwa0hMflXKP23lG5F
GrHP/w5IXsR1MdGqtK+NvkO2CDTVIPATb2d+47uVs1B0+j4IhPAyf0FN6Wyw0/gBqya5oaaRdf7g
G/X0rEfZVUb6P7wTExU78ZC7i0X6hD99Rksua1fU255FSpZ6O9mExuzj4uxOjl05aly9zLY1b1oV
i/9Pm6vKidvKQJlKPdvVz3PwcrhtF6SmNJkrmwlghGsRmRa7U1vZmWH2Mg0EgrJytpsKmnz85m5E
Q/nnZB9IYbtoDfgd36gNpleY05bAmnIg2WJM3wZV0HVi1RUq+mEaz/cTAPuBNI0DQiGPJuPRVsb3
qB98LOn2GMIir4dls0Np/i2KCIx+Foq3M8TI7pl3OXy5IAbh9dV7Q9+MfVD+GmCETRtgZajXps0x
MGlSGjRY/txf8QRv7U3ZCZphCj2zJeQcaKx8uvS0s8kOxDGW/4tZVS7Zs1F3eDgBjSnLXHrBc2wb
aziRDhi/ibtJFoCNsZwwOMdKfWPENAnVbjIvjnX98lpMRrqppU1HT8h+BaIyEK4A/GI5ZYZSGYNx
zqooHBrCOWC0CpOg2XzB3LU5N1ZID3yjsaJSfCEa+JULPQrp7hTBmBgUBdzv55Bhb1uM1/RKAsMo
g3Am9q2flBISPJeT+M1b/wBg7DMbuANOHVPqSLLonksKou8hKsR0A+cOKJSEZ8nbOKhJOslj32MY
CZcDNEmKiq8NdDJ6gDkv2o9M9PoIGequHDCYuPOfzgAZeEL3/AOQcU982HVT6DK8ZpRVJg07zh0b
iYC+zvT5Q3Ow8qJ3Gh2gZ9PI+WZpVYXpp05WAE+NtZFcRpTNU2HZpg2Zu39LAoJXec/8XUJj0jJQ
15M7wbLkFfm4Bez42RmgnsfHU4eo0D3WSRa+hp5dnmnLC+3jumO/KTFW9RfKAN5H3HBkQPBIlRn1
klebETLM2/yrRkGGXxPykrsgWxPW+b4jwdBITI0r80WnncGxbwwjsnsGry2uPSQ4qtcMfD5n9vf+
Xep5QG+qHvrMChbOH/LrlHcKV6pGaIg904o9sbbqMqrv+MN0E4c1zFdmJ+NJkdI2/jjsGlwn8GtD
q4A9/X4eIkkG1xkd2vQQv+evOWv7swIFlIjFWgk8p52v9/OsE8U7W/PQeSH/jBbVYyGK0RIyAEpP
VmgqsEe8FfhX905HjdJfhktZ5ytYAw8rcaNOun94LQf4/PlPnmgL2GOF/zuvgwX6DilwmojjQV4U
SipXSXZv4EmGJ7FzkhWEZ2gEYOVipiWZW0Cn1z7Lw8zf/jFhzwJNIuGzjgoQmiLRhwAcEw8lHCVO
0fBisxzPngKR03Z7QmDw6fqOoMDs7sdXusrBrQSwBsmcuafw/gf7ddikfgHel0Dbxnx84tAKi7Vc
rCIDrux/DDh1TmYOVJjM1kZQXa+nH2XE9iUS7/H+uDdKn888YydG1Utkxn8hEwnta8TSil2u3XCk
EQD/7QZJoAnxn21G7JjKll7eeFzgAs8bNLnPkQ8faaALQZMvfggA9jCrkEXGK1yDH4o1AZhYwmV7
NiAoH0MreeUuJfXx450CliNa/Q6yddYH7InkLgrx+aeEUj1IXCWpFzHSf8KOqBI4yZzVZGVFGhhA
8y9h66t3pnJ9Fc1Ijt1tE+fto0ZOaBG50zgUdnaG/cn8UDRigROZpuFhC5S0wsJUNyxFxpfxqRVy
GNZj6EKNXTSsrCdQiqtxNXUWUb/OtCLP6vko9nGgijScPVM+YIH2sBwaZ/yU6MD5DXIYTVZbkmOQ
gVZi5nezsnmkN3MB9qeeu+xm5nlD182QSlqNxh2Yv+AcHrGpocI1JEHqYx3ExT5LtddEy+/la81D
luM3jg08OuLvlNwit94z5hGcBnwokD9OJ/N98zPEaZ9eN/3eicKd2T8jcDKVW5nFuAknRl+TCqcu
VwNnV32ojaO+GgwLA9IWhxiGC8t9SQjM6zxSv9ZzAsjpqeTroQdbrstE0CHvdOu5ic4QdO36v99v
ZAhYYHXQjWDqqeDwfLwYWqrbEfnr7gxnclVQY2yMJCB+6rg2V2MlGmjwNTimlOTjkAXsY/k4caMD
QxqIDgs/RgEy55kS/1oGZ26FSD9uE8NYy/TDRnss86g3SQFPnqhYd/apWPlRNvduMiLgEZTQuLNZ
G5Z+isxW9T48ATAYKoo2kYHXtk6eqLIyLrup1O1To0IsDXPVux8rJZcErIZ6bsvFhzkwW6qRB0pS
WPOnaWPtolw4DQSBF3fbFZLsGhwgJ6QRb7gTmOONGy1Sn+DmdEkH2DFLcyCaoylEYQ8OcjvcXQTS
PS2N2BpTXlNDCIJZIRI6CzpoY2OXTtWtLFMoOjF86qI9AMrY08NTGa+fXd00h1XU+QmZRgJ+ZbTf
OfxdHMeURcE3nen7snynktEGZNzk8VDMVb3hPryObuY7U+tkhA3lL7jNAxtXGll1lTHLSU13fyAQ
lpLV/+8gyBmqi11KcUPbBckRFtbEwmlFkl5hRkAgbl2gklGtg4gzhrA3Oa71aK7WRayekp3KQJyy
m2YsZ7ro7Vz9B/hzq4cURzBzC2S0pUP2iSpHXX5CpiDDHdY+by1zZk70DFlKlHS0GjpmejK/q4HQ
REet1jpRRbWmgsmoocRvDIn6oZY+Da1Ay7a4cxLJZ6qYINNGRr19bCwHNtvY1DfVoEE7cy2JVPwR
UUWCe/X00uSRgmVzUWR+X43WQVBNrb2KlLO0BRUpMH9X6cWecfdCSKLO/BWK+hqWoCRps+PpE844
wLnTkvAalbQEUL4/Q5otvOpni5JdxSaxUAcqK2bqj5Oh6RWIeKhSrzlCZtRvRYfPzRzgp3qYKGnK
2vOivOWr5hll4NKULSwA43gBex5s4y7i2d/2QnoQwr3S2IgZi7sLp/W/LtnP3NojwMPLI1bPZOf8
p7C7VcDIDWglLyw4ALeMqSvHiLeeCXSaoxKffTzJwJGWXDeZyAUUoQ1lTr5nEWqcKNCmRYj7/Bqv
1siwrr23UjIYJ+aUDDKijFdEX1aoTGKk7Zp0thkQZK565BMCk5h7QgY3Y+/9665Jv+QLx1RNggCp
5yCb+R7F08KtUFqrNHkQbuOES2lrkUCa2dvs23LN8wQTedpJiNSsI0p1ypsR6fYfvpXUOohiEd6L
qq9Rq5oKrAqAanaK42bYfI0Yk8lhHvQxnUuhmUiWjcNOwhI2eQAyyOwX4xS24pOQ7vGz+K6ENb/M
dHrKQckhL4hENAbwUXccvtbZuFE7XyBbXgHKxydkiA55zbTHAdT8ttXio9CWnyRFoGCGVqIkaZWe
HlRkTarR1oucrlrbbzITfneldC2H4YHT5qfaoSFZSlGLO8aa5f4kQ1nY04VTNBt1YTUQM5gLthEd
pU2FeE/GE/SoNx3bZnDd1xJWyQIBzqID8FABDpLshxHMZhWpnTb9geBFSUM+hJ/yLs/DgWwFwwSU
kxyF+/FGwlu56N3gbDDaogtTNRdHJ7tXwCQXMb7PqUDUMrfvZl1scXlOZpzgvr6jXe5eTcyj4WDx
xeUYYZM9GRZPBQgPWzbc/AFneH0NsMTmkIp700JscgzZbVzSu4/QQBb4GKp49LwvnCrHblt16bat
OxcbnkAabpj93dK/UweYQ6vlU0SG1fNv6RE1TxM6yi+DIKU+qXSa0eu7CVi3Hbakr2EcS1/uNCKw
njgP6EyfzPO/wL8qGMC+BxU7d5QZkOq+njd7UHv4TYzdRzKwnuUeNPwGjXBpV2JjnkdyrN83S+Cs
sSY6JwivvuP21mbj46uRiAQPdUlSCO3P968T0kPFxDZxN/+Zg6DiGfoDcLmKjxO7cFPH6ShExFc9
UxqiN4GqXfNIa7/9tXmjDtTQVUm443buQ5LktpKF1zN8tTuqFBPrvlC0RGOKJEUYDPuosR1nAmgU
6QHprRxf3Jgaxb6uWxt6gq41Bq0xv8lTqGTkIQKPqwEOOuwhXwa4vNkdoveFyL+W5lSdq/r3JFDO
neocw5RDYJ9sfuclHA42PCA2SC4UTNOJyQCs+nZM7FghnCPPOFo2Du4y6je2HuTZvN6YLojhDTQl
hZxp32joruZ4vyStmJnN0Grs6v9QAbKdmvpmpbZ8LVa1WvormmVLZFrwRXsMH3wjwOZCv+CeQozD
aW98HFsABqxMDqux6x7aD51g0G9ejsSA7rg3Eb1tbJDZfPM9EmBxaLQHcm+OYoomCkJXh6LzRtCr
htJz4dRcZ0ldPimIqiZfbrx503pxDrQIHjU7S3Xvg35E1QoTYEM+4MM9Ub26HEt+bEJvZvhYzVlt
0ZntPdeGHK3JQYJmOElMviMeoILZzJMhJb9QthSoPCnsr1Iudcgeap+iqE55m2GL2ul2pGBssBj6
IZbWH+hlOxFk+zmLgEMA5keo92N/vLdRg4neA8/w/eddHm+qyNAFY7cDyPGMzGO7A/CSyEvuH5N1
dci0aYppf5Vp019ZjPKLBVmCoXzCobNwQY7wxg3w4jZU/00+q+HZZc7V1gPFys7W9kUk02RkJVh5
Gwd7D+utg84lwrJkxB7J5vi5HGOB6jJPjbI7obLC5YqDpz/jdVB1HeOjlIdMVKtiiYl8+lqaYrWV
nJPNHybwg+s1f7ED8BwosmibfC3EJmnqQppQOB1rYd9Qc0BhYE+0wdPApxFlDWrLXFE7dumHaPiO
qeV5OtWP51tRg4JgOC5tRpK+usjrPvC+NfVo6GQCB7lLbkkTVbPvZ0G8Ue5l9hNMBsA7//8WF4CT
Va5X64nq45QkIod7D1gmIkPH+1KiwIQcMdnL0OeWYk+PnSEP+NkoAPYYDrfOSkxPZ8U1Bhdso+Jy
YZ3yxJ93MWr3+hq1iHjp4CPBAIwdDwZyQZWSH+YDoSbpJ0bA2D/gyz6iVQc53bOzX5ehmqpvlUu4
elWBIpqUnMscYNFCMvk8Pb5cGUA50lrgNsv/KMOSUVpBO1Os6uyAihN8w0rcBiicbyZWdIZas3yV
OqxEC6sRyXpQA7ZXcPmRFGmbnBaOpZBnQqmUfpF8t/4RN6gmAQcWY0i8wRJMqQDK7soHDssNgls4
ra3ILu5Nn4qeDxcidrP1FLtEaSQHWvz4lls80Si4BV0b+rram19ZKiFwC9/rU+ycIG6SSQVrIkkj
sH7WaBQMEVxkpLuKRYC9KFKdw2UJ4N+Ac2+zPvsnC7tjKa2QnptkYOv+jSVXJTSqNG8JNOZrD21n
40rD8CBg9gYRfOdNZrhuXcTyTKYRE5pmuG8DZ8AeNkhlg7NE/PGsYjkhES0vOUKL/6AqyJJzm2aG
Gz3L9JckOoraaUm1dibprSUcBIhYHuXpgnzFWWyXOxz/ioayhdfMJVeTnxY5sT90wgtS4YML2L/B
aoobgbRJaop89czg29PwkuUShLJTj6HY27MC0CHgT4ncUwg0TrTdklbmBXnnwlMttNaTQJWbnwYJ
VoCbSDbOvyrw1bG5uJ4ufzP+09aagWjovamFhO33lp5YJR0Xs84IkenJehE6jrnz3v4PW7eEgStM
0/Trs/poseCadGUkDu42PN0FH3WJn/JlxdQWwCU85ukbdRIVKxPduJz8oNZre0KAW1ShKTE9wOZ2
KXEa0Z61WXjygCYTJdODFpEUBNkATCskPPm5+233F41vl4wo56mpuRYp4AO0LGON/ZX4fjn7p/5i
gOAngbGWxGp71Q/m/HqX1x0hhv6CceXhSv0AG1e6OG8Omo9ayUAavYJziDz1VFJxgbzsF7POSSjt
cOYaGJhvp72lD1h/HYEviX/AWq1DP2yVZ9AHeRwlbVUVftJvlLPD9BDoS/7ZEhVnB7jiNB9V5uJW
0msGLf1qnsDu3a2f1dv8xGnXFGbKjJEOLAjQq0wPUrFyy+zFXrEQ7eKwRODWS9fZF1RygCC6Tcx/
mGHjgj2KIV/osapTFS2BgdqdCEmcWiUT0tc1lw2U3i5SSnVkoC6TIvSzkiUWJ2r3GFR625Ai8rE2
XtEtOnIzklabtdhRiY0nYM7Uy0DBxAVMoKIL19kzh4YehLK2f94Xcs5EpiAhjxf7KMlZIq2Jpzgb
F963rzdXHXPIpfvQu9Ve0KfDcPIl0ayRju6vHISAI1EL7RNFH4a8IAuX6krObAhxN52jMbQIoBLC
JQ9yQPmPnz9WSaqjTIjVVMk6ZN68ds8Pte59+fOXdS2ctsyYBAXh9T07rMUjydci6xgzg9WGMOsx
L/CYD3YTR+pE70XGzaH9czgw4EvTH9qYEU6ETCOJV0BQ600ieZZPAzcBO8y05dBYmGs2FmCsoyfo
rKtMKCOGRIu1nXp0DQMyQHkugH+rF8JxuRe7wpnaEz4wByBtYUE1tb/zzwVuFqENhTLOF7Y5LpL1
oxRYB6V0jJ/5RSTssl3NgiF3OlJHm9Y+pt2nrT3Mc+9BYxSX+efYbpndYIzUU7EqGk/eY438WttD
HM2j/BBUYGSI+klEh2OIdiGXzCX+4wdL8waTo8ltjTaoj+PND8rgzOLbeauNSIyAAOpxErDFC8QP
jwaTofU/LlaA4mNCkrPtgSMLFfbHPAc3Zi16IsKbdEsfCT/vy3GVg6jGxMf6SIqRKUMf4lnLA0Xo
OjZKOd22bm1bX/z29DXUMvy5iaYACs87TKUQgoso9FFXvDVUb4/NV23trLptlXnUFAaCsbdA85ik
lRZDJAgKEwV4TYRcCFi4CleJmGfLis47FypTnqJo9X6IgspJs1WeHEda6F5AYByIOmQvEMBRgRQT
F5Cdn0V+QU1MEWRAT6hxnl68zDWVTa4yLRPePKDdI4dI02yuwhRc+O++l4wr5gHHM0nTMXuTvDXz
tBhmWEfHr6BwatByWnWl6FoigDHb13LsbE81mjZmz9jISGyBqFkPdsQjG5mBCMml8/N5qXsiyqyf
9KxsM5vn64I2H6jr5Ajzk5vZQox8biJ2v+7pAEb0Wibmz8FxZghMeZEDTyMikD1lftctNzzbg5WU
FM36I6FS40WC8cZKvhX3RVb1zwbC3Gt2l2ZnChjS+PqeID/yhMH2FMcro02RnUSe2SglhhSoARUR
ZPxLrEvhbFJgXWrswsKmImvI/xCNXjJExxFzCGkU5AHljBcpdBmjrv+1ZIwS+LnPojqN6rdantWt
DyFwdPM9YN6n7aj+cqB5mQUGr7/8TLnR+R9/ZxP7Ug9p4ky6N7cuylWsyP26mx0SBW2YvBC0H7wM
gV+SAf+EMZVyz8bQZIlbL+EVLGnep5vOzrZP2hIHiYyhgjmeasbQiXYZ5MNzUKYoIXc7TPK9AnHA
PTbbb7NRpUL9GiMAB8b7eAYpFK+FICooeDWTkHzLJKavjUAY8J4x3eh2fsefLFScqZbgl2WEuCgd
BAwYVTSX+M8XcJG5TXESGSwzyPLZggt+HwnnrAeKqQFHrMSfgjVxHXJ5Wpb6HgNJBkiOiBkNJJVB
9NppWlsUT949pI47UGaNIL6SuTvMX1wjFaaI9fKU0pJVhlpXgo8lMIufqrH4HWYa9ANHsDbsq8Y7
RB8qeYWRjXc/kjG+Dzu11odbBIa7ZBf96h1p1Aap83al8b8m4TRJ9cE5rk9L5orStmRY6ySl+ieq
5nb1pb6tGBYdsvUQF8M9AbwDBAIo4BDPwlayaGemsmKhdRUbEdmRDccQbwWOXfgny9+Q2AZN6U3K
kLUDBDBZuWlFZmiHTEScjuD6P6j4qqzqUXwYNjph4M0sAWQJk/+WCJb1dk7JIXSzoiXNCOlaCj+Y
rV0dZpOa0CU50LIfMpY2CuPrGoyzDDX/HsSgUaEFEfGG5MwsK8fD1OyxH2I/iLz3y3gcQYXsvhNm
l8oOn77a6sxTQRvyo8np9+fOme7XD+XFD0iM4OTs2SuhRZnHzwkW+1zZKlt+t+e6lMFnbMZKJtEa
jxdaInh5BtmqfkwzJS+kRtcjYvbJ2USnDmpDMkNwuQ9OrW+dVzsCruexcPsDC+Z2sYiEGvKxUXtU
26jngQ306wPAtzOBmBl12FVzrD0KYzN5a48y3z7WAiZPZpAigffZivZfbRHEEoST7F9qES3dvoau
NV7pdzImA0RQzPJCAXkIrUfpRkMkhb4ftuML5iqnJnpoNPejQLXi4WdRIk7F9vqdtQvkwnzqc61G
7P9zoQw788ydnY3LoJ/FD0Qoqd8yrHLbbl+DZKqVQNz7x2qf3EhG2IszXTUW65xRxNCSFNf2Ck4n
7P+GZfLfSWT2j7IIPvixzt+MssXqhKhSYq9ronK+6cVi9eOGehrLSD9KkNRHbC2cpNWVus1PnJEF
Xxfk2ca27Z43TIh+A38kIUSYHQSmfdK58DDa7dV+yeRxjvM/xtKwKgdHQRYpeDZKefgwXvGe0ajm
7M8WhXMFrslTzj4UeQfV+b/PRoZU7huP+47+3Hb/HrGy7iKGSIp1/rno0nBJC5aYZ/SMDgB+4RC1
CDPCkb0rztqgjl7EJADtJ1l0U6OadmpORgWHOD2K9AnpPD3i2HRtpESzCFewNwrCohfmVCW+bHgL
o8yCPxPE9xiJW9P4aakmmQvBNTSVj6uEJiJehqYxUiRoIjN/0T0Pn0zfb3DS9NBFieuJx0JFEwDB
bcDnFSCmfjhGT5Hvfsb0yV7iE7mmyjNaF+AQNzXVEBe6f1cxdgp0Rlu8sdwCn8wyNWzs/CLJEF53
cIqgwvoIx4/bjTTGMo5P9OfBd2+fVYBOitR5t188egtGFiUNO4m7ePmRstjgMaqRnBz+prgWguRx
MCYDCRNHX4fPIFPdM63C7am7nE2FvsGluH2UB8F9WBna0+2T6xIPrwmQmaCsJ0Lzj9pB6ZdH43wA
WMl9gmeW0EjCa9gAdqjQKrLTnmtxblBw5+Ge0RfD0CgClvyk31n3lm/n8ru7jpDm30sq8lE0pt1K
8DcyAUnBjgMgJCbNUKYOWgstgkxjBczw/4+Q96T4d943PY0leiDrITdtVwkkYWq8wuPkm45r0XpR
ggCco5Q/oFkG4vsXHZimICHexVVNUUaCXA8aUpoIcX6qG7GY8iGzj7y3d3YtY4m6VlAaKS0xv6ih
5XoChypvUVCxhShb6MTBFmoE4uPwIKgXwiy8+nwLk2tOgAXdTSjTJnlvFp2WHzPjUElieazYbcBs
ras7E06Xx1AmP21n1HPzlS2+8gH1vTSjnodB2rg1HmRpLSt2sOW0wjMMgwX+u1u5fGa0Qzlj87FQ
7iPBWPSFKeEovt5N2r0bMcZ5PewYt0GwEy/i6uGb6glHODB2A/jQVwFygBZl9r7vGPyJt4awRU0T
BtBqqYVAhxO10vXmPGhL62sKzwcl4luPNmequA2hjN7EfGNmx0h4pxqWEJh4FgA+xJfIZhfb+MXO
0ELbjf4F/MzPBvHsiR/5OIz2V4vbADk5kqICPQhwxDF5yWTzKJ3Cj+Xddtyr5uW/IUYimy98hXpf
w5sr6OH1UiicEY7vzc0j3bMzb304Vu/oPstE3f2hmK4PNcG14tKr4zk0XwOFacJNCxgNAZ4x+gpm
n91XWIxefLN06gq1b/JcBoPJjW8rudOlstxHza2ziB5nfHKqyM8LIvcmFqUf4MUNnf89Q+AFrJ3W
a56t002gLFSmCc0MWm/lxrMKmi26863L1H299dF2tDdnZr7MO4Vh6u/S6oUvkpVVDDYe+KRvzvOC
m6leF5ybuwcQkf0QlWLqhkROfaewD3KYEgJLZNx439iwmhgAe70q24BPZcfLD+kDfzSCZv+g7L8j
hb8BJu2ordWkQWOHkrPwkC+W/NDUIKpPZQ9Go65jyzuVN9hTfRT8EIWlkqZNL54CBkWe1WIyezTy
mMUUdOubQMeqxWdZ1lMAd1t8pdLknW6BjZfqliMtgt+mlh/aPrRA60B/DiHwokpOSr5YolaMydL+
v/9RqmckNEH8Nwdg7eHElTGlPzuFY2hUbL9dIsirt+bDt1xPfzSQ/zpY28En0gQF6kK+I1EDyvub
AxqVmKYt/hpY85EqAcE3cN1TR32l5wm1Yi+P3aw/RVLC9s4LVf2rFwdKlePZxmG5Uj2i41ltCZw7
X2XlinYm7g2bwuk2rdmhY+asAIpFeE1EzolC+Pmc7DAvDMkisXQzebeTwYVLkNIU5N6I26ghhdj3
g2KIalf5zJKse1tc/j271QLRYuiDrVQ7kAPxHS0ukfLN3kBpwp59b67uhSbzECAPaPIepcBd3/uH
bTCmlw6/g7nxhlbKiyHmAdcCLbgAGMYiCUk7Aoe67cRR88/uKLDCBkiHfZUSCD8bqLdZveZtBPEb
4zfnpREcmNae0eKSH+xE2h7w87Qw+0TqSZnzuqPN4saxZSIY2UchZHf2AlJcitJsz/mwDB69y4ST
7Gwwo5Cb4sKG+isxSdHrEi0JgvsXCeCvmGpYQ76MhX1c1ARPDFXRuVlQg41MRIpFGY2ki3VHp6mZ
blCzdaaXPAUZTfHUoIKqYn35yJtkHovbmY8KnFn9KqVRzHGEAVsZidDyhzlKCkeAiyrYVUblEm28
uT2A3hxeTq2UGOL9pfzyluqMPlV25AtdJOSLl/Mwks2PDo25r7iUS7DiZAR0+jxwmfHdYvWFIirr
tMYxeIqgIKoEfxjInh7YZM91UzJYXfdKw+edfapXoHbzxxzrRfjUCSINwS7ZiuaPs55iKc9hKLSO
GNuqRdvvz7a95T9gm58ZY3xlVd+Smk8uXlJcJXH1S3SRaMr0wkezjzYCdNrQeYzzf5iQ4S0s1ou8
otaj0atsLav07lfoAe4jwGQNc1BobhlrIkM9nF7LZhXgY7kbc0YyLqFzTxR/n0f+ciQI/xF4ecaR
s3S/HsvZ481xPH8whGVwn0A4qsTAs0nC5tGafFMoUnzgIiizCJqNn3dpx208N+5jNVkkBztxP4R9
jU2702FR7vRUJivBd+vCWllJIZxEKj5pb80qvSU1pWtE2DNdLvYw6ztSQFa/C9glppYKNeQj2qKE
/jQLwQgqfcj6tUFtzMxo4Ww7tLQsCBk6tqFn3oZwJSwSUzqgr7EnLXVq+mKME2h67QAK5ukG5sY+
0woW96lQB6l3poukqfus1FGUdNbjBQpdftP4fRQgOzhFLTrgmBo5tqByDGHGrNC93mm6e0JZWSJE
LOeQTpsUmcgF01lcT2+JaWuORYKDwx0x2suiE2jUmCuMD1YGxUlmXDL02AbtZesDwLs+OsdgTR3/
ktTeFgES9VggK48VTrL4msTjwwGj1jcVRQLAzTENdaNC9NiyoISzKknskkLow9J3eMZiFEcwLoxe
xLiFsy0S2tCnGfCNI7ccOhYZ03uvKKAdL+ay+WHxs/EaxztftqrQjSri0XCSvmvkH/bu2RPovKRY
6PwXZ/chVt8USKu7L4auriMJVsltk8f1yNT3arA/s5dclzExtjvFgiIzidejbPNasR4eWzfWuIpj
kwwSDqlrTwGFRSCfDABDdABYDabQ22pknRNR7RaRJEoQ3izCho3P12+IL4eG2CKVJ7vYvYFZ8N9M
A7vMpRVpRkEA9jvVA62/OtJS3x6pFsYLeSpGjFOdh/Ad9Bg+eRC5c/3YN7cbmscbDLfHhqSKyjG+
zQ89FBbZaLF/Lr9u1RF5PhW1fQrc34phTtF9c6CbMRzD+E+ETeJzAvBsOqF8xue4c4I4xNd/7o9a
Mf/ML+GguRTj3SC8QqkrKLbuAznsEEfgVA/BD7B2njXQtJFeLLoj3juWWf/geFAIvG6xhdgQy1EB
nbnxt88bKpFYCQTdAzkktoZv1oXUMgvNBW7VDxTtYNu+JqlurYdCHLouIjj2E9cuw47YBEmBxKcb
XfTswQ80ynlucOLhGOSDkfeTH5GYgdYjZrgn3Owvg8FG86y2dePPTTNnRtiuJpk/vkhBAU12QXz+
XSU6n1TG+3XFR0QUDFdEt8Fo+NBR7rPLGXFg+wGvh3KMTVTBfZHJkIS3bl8Tyq+d2FvWcZiKT/Vt
7SCR5acRtaMnSvDh5LW13i+lsS+R5rzaKMCLgajD1IT2suo2FHuUiyMFFow2fB51T+XTWhIV7wms
yNKhB/cYZSoh4OMFpA1R+D7gVvme5+g6BaVabLzovkJvZqz5di+KUipjYYP0Fh8hzqLYGeFldzmz
m70uFmJewM6s8S4ykmNdkDUD1YfNi9hSpGO5H8I4KAUbDgRpS5IaQsQ1vjJl5oyW56hcfo0a876Y
KPT95n3fCR/EtdhrRA5M6GKwd0Vp3RDsypHdBHRX0Q3e7lGu3E5218D63Au4eBC8Fs1sBKgzQUnw
3PpIDej1MGCTTqS01E+4pm7RG1SvCgFpOUMr2cirPkDkH2NKqQec8lL+ipNYc3KHOmYXLadoDV36
+1r/jLmr1vx4ZiqfgfCe6kOYtTRTwyTy1+/SBkYUp1r/8fy5t+71NRDB4jqbL0nmaoY04YG9foER
thW4h/U1YaRMF55AgLvWKjB5L91LlR44nfjm2IReZpFLovSDlm1FBnUhCdYYqIP4yLChXc2OKf83
JtsCqZ7+R5FMzeZ1P5QXbQzf71Ca+WYTQ2hxkMIZzPhJH+HpQR1otyFqxTvWhRLyr5S7Es1LhpUF
s69v9cGuXEF3uw+InIW0xf289fKXiJNinBlqtrN+OTY0PPouyW/hR4dygCYxa6XC35PAtUNv8vPT
RBJO8o+dX8hnS3KexlHN7Onsv5OrQYY5ndid37PeQIz+dGp6rt5HX2uPCJ63NN70hG3/lDPu6JAN
OlDXOnLWi3m3YzfHVmmKq1syvB+ZO+B2gk8zZuIar00ey5y11VHtEbhto+ZfdU5yUfBb4uVYchjA
tnDql5PhVZhjbghim5I7XJnMSMFcjOeTVYkAHgAHhqXM7xcrlQhSbqb44kSXfUbA4PnAyeP+vZ48
Dgzyq8kEq76YLQX/jN5kaRHnZbpJ33B3qIf63Q6JWvDoYCv4+rZZbfXbqnDqOesJgmPxpPrHz8kW
9IpFsB7HU3KCj0I4WgzxtKkaLTL8AeGOWszfNlxqnbOgpus04pP5K/gFTi2oW3sbbqkYV5tU9TnT
4NTdPk1ftSO6TwJaKFG2e2/xRhcXZUX02lYLe6mQTUxbLiogpF04B2RTFhRvSUoBusA58ClfEIP2
WUZYoh0jV/JmvbwhqtUJdmId8/80BPYQt3dE17TFhMqlPvDKjfPkXs+WcCQOVVndbVvZer4zHAdc
X8fwlVwT5bPbo6yOk7vyY4MM60gOkx6UO19U6pv4H0OeP6gEkqiyWTcExdXnldOraYq82KjFnSeu
nA2xDGD0Xr5aNYgjdvRjGVkSU+7aycKoDHJGd1nTtnHpg8GAGM3OSyM7hAw8rN5nwACRSS8BbKPJ
QFGWXb+GKoeiAzcpmcvSoFT4m649UY3I4szBQl7lha8q2AfZ07H3dRoTMxLVQL2UdnWxEpbspe18
7ZCsglCA/MJA8CIvwGwWUrJSLxvwu8f8MC5PqrG2RjvvnIPGLlljFRUISb4j+XSyaeRBz8cu8RiG
Q2RpAdbOfxhOMX598oQoo9pKDcBIrPvQMoY1MaV36dKxa2Pr9vKqEnKFA0BumPwiQYrqi+dDQP1L
75zI5lNeziICCu4PMpzpM57mY78xU1wNj06ZYbQFzUBBCT/A9ZIjq1RuW9E9o1REONWL5uGLdCOo
UfDDxmH9Ixs4ImCEUz+4dKKn53ovaP9g/yM0s4IACArfged5e258t2Xt/pfqtBUpqYOXVK4ZzOcD
x4yzvDNL1vKvc7ZInqa/qf5ERuZ0gUQdXAdOpPKoJLTA381vh7cS0aMEFo5g2NUs+W3yQbs9ExAW
zQ/7xtv4Ul/K5x7+SZ4koCPq/B1CoNNovnBMv+phVyibbSDRlGG7KoanSamZscQXIgLeqSGFpFf3
sP2oIhji+bJi1rki4W73cZ0/9gJqytY/N/zD8zO1qDWXVZV0U00lVAO0ohlpUqNA71ZnHLDcK46s
45J3F6hLSaIHGkoe6i/fYRRbR7XKd4JJIqm7Dc+EIlIv29t98h1bB0gYeSjXDEJZvZ/jNZozKGw9
WZgOfN8TIevKHHMZdkE94qEmNYifVhV/vXPzuYkR1P23WjiG4oC2wW5/vxAZ13yQPT+w4dd85Okw
I/9PBSV+DoyZUWMNz+FLOk0tvJZrMJNUi1jP0JREJz9jZqozqFHHNNfLC+PAjTUo5VByidtZZpxT
08ehjj+SNj2SrE8DR7N3yOGsfZ9FaTvm5Mk8C+ncVhbTQy7+rNirTALVgz4IZTGUs5VWcZizJ7Of
00xpTMVfNon9NnwYsIisezNh27qZdrwYQXnp2rvNEHNmBjD2fZO1Md5Y8xytjK0+Z6FgL3FkWXQ9
wPOnyQ4sL2Z/LDFCd3cPwrl90fgH34ZRcxdLpNnH9myBMsH65lyLHQ4eG2TshxxOmJNMUUjo1N0B
sOaO0M5UfPfkya8huf6eTe3HZynqodZl46VWltpXE6O4w2WbWs+po+bXJ5L2ZQ/YQ2SELoOcD9py
xP61caLZDDyiuzIJRqgXMf5yvynnf5f98js9Ugm7koaAUHfzH8cUH0f+A+ai3o5WXyMf9LOIZqvz
kzRpBAYCwmKYnsNKnua5YW9tTAc5jodGikBLRqGrXxkEqs0cnRYTwUpe8k0QSoSlXQzJ9fhFCfsr
Xc9KJyvCHI9bkRDPcjMwlmiVXj8nuD5awAYDcBQQ7+03SE73R8ufTPukPKDA8NNVmGmuo+IXIEPh
2zZ5HTTKnUyQOgQ604bS8xv0hDhVs/AYaqWA+QyWBdsAr10dw7uUIHHJcf8wQ6rAs/cc7iNkvLPe
EwVyi+FASgqt+AX7z+EcF0ygVjSe7oO68+3oVfV5VxbIUaB97EvpaCR1OyQhCvKcgayeLBVagEu8
9iTrPiOlmKqNWoNqy4uRt4Z5x9b1ZO9Obz5zYQPJVwudTr1gdT5Ppqd96k5kPl6h9KI17r0VVt2h
kZtUv3NxjDnw3sNvN+CybITFGOLS94fJLmQwLAebPrVsJ6F9J+gP2CvZo9uD/fPWi9jixWiadmd3
KrPv0MpsGSGoZM4cUng9cFYtk0DWwRwQNNcaTW8W05lYu8crPwjo8BOwl/xU3YQS0/7ULfPtG74B
hzujmJ5ZhU1S5XKo4kC0DUIVdUEk5qxZanTbjKq1Q0BWC28cgH6qyB10Lq9ZpUyzTaMd7IQLUM2j
dFToHrtJ9B+nMD8B2Ws9hfd+zWaL3ZRWG1NqkgI0ezCE2c2HsenFiihNG6QC3eYlhAWXtkhjofeV
j7AYtG6nobqfRhpV927LP6qkRd9Vxzn5bFisk8+YubFN5PcD7TgtKr4rHUCIMfQgiGHHEWa4PBjp
QCPnChkkSkJUuBAwOtMS9FuCpV0ejEN7GbbHP/aoUVd+kbUIxSSvsvCvX6w0hJob4enYJrroiQKh
1OjsVZSMaFpFAzFiYdq6CZLxI0UDOPYUNMnlf4KPLs5BhLf7p1AXv3zINGyfJey17QRT2cjqyXrE
es86xwu6O73V9rUt5+FWOCHqsLZqdyoqX515f8n4Kgi0TXdBIBIGO1iDnutkKRl1lsIyCGLsdREf
6qlz/hR2ompQRB0WFOf/urjA/QM93zCvVUtGo2eb/oPn0iNL5yWPtTazNYugAd3YawNNcJyVIG3I
xGfuGDI46noFuWUU6pTEMM7MRJVN8Vn2zHp3sJg+pUbZMmOGcr1F+nG9nZ2NRpDdafZDdhRO+/Zh
DFOuTLcLFPN464wRw97ojrgm48y4cOhSdsjvzmjCF1pqINJRY+LW33eUZF6v9VaEU76UYNIwSGJC
/9bQK76k0qL6kN5kdBeJpDiuwvn4nfBrnY1OUkIWxL2dyvtKGYseyfOQyfEJhc+L2zMDAJVYEQbE
/v7ZyJ13oWDlc3dGX/qR8IWU4X8JQjFHur64hpXWVZQe4PQ0Qjf1BaBajdoV+WmalBggXDGl3kDP
G5wAC5vVREN9VS6V4WdmT9RkKxTqCibVQ6IgjtyTU52lw2GUOYtCSvuQChYemqMdz+CBVErAdsxy
ZjyB2XWAu73ZyI71EuPULhoPFLD9oENiOi/AtQb7rxtbcyLtdY6Jcg3i1gSWg0C7GMB1YpaO+Mv2
uj80ZhwCkHPOxq4IFVuHYEbZsrPiWi8DXTDQLrho6qxa2EUqqtQELZEt56iwAX86fsQmBqoYY8C5
J7idQ0lQWBApNPkq5U5uoitbhK9Tw47g/51bPoe49xqA4rXIgCpySne7kOss0U7EHYK3KiaO9Od2
oPrU8GPxhHeeeFbqYhgQdyp5PxN2osGKT2NM6kIKyZJv27nxIqp474YsLffUMjEUfbddfLcuGqt7
Brw0InNrGhLTDKn49XCh+/XxyLVV54eeWHvoXpQppz8pXQOLG9uvdrH7ME+7Oec6AtDV4iYowNej
/b8c9Dgqliw27C2cdotfkjrQgpuQdQiHBBVrungK9WXx9D0hLgfGPYpzUmZZwRaLJ6pGVd88v4D4
1ck28puwhBkiOXFJme3K8e3FMuKPxKyii5friphwyFLX874y0/HTn1fTiOOuvYYKTxpAskYqFl8D
6wLbVCkontd7aT/Fah5vpDd3R7MM02eUVZLk5ij1klR6Un06cCGz7hlBjow2PFazLFP24fECHdrn
JG/KWMuE8wVS7eiTUDUHME4w2QXnL2jvoVbN4rGmI+PPHejHUlH/tWg4Zw21xfmFI7vnRN54rO0I
zodLjJcNj0+x3mhploGuMgFixlhJyG+mg6a6gXfW8nQvefZOTK4lnW8w/qCfj6ANiWPrFOsX/Y2c
BL8NAsRsXe2foeBgEFhJeSgi2E+UbxNzIeYjMeP6ym7vwYdjQNqCDYb4FzO9TUZ6vNXA09JjM/Yg
h+/5ckrcgV4aAsWt6DT7Kgmwp7aK/r9Qa8wA6drL0U0iuhYJQi7ubJZCvXdAf2XyiLxmW+0vifrf
onmyzAmUW6Bmx5onh+PBBnKJmW4AjtjFiWVeuJ2vGjwpbnW7ZzJCLWsIwS6sht1ehcoucVukXXI8
XGgyILthuDxs2ay4hiZiDsMMTYcdvGlmOmQdDk+oLarHoc507LaC8B+0FhAbLJoQbrtvWCTfZqZx
icRg0gdSAfkRkDgydSvxCJ97uYQ8vwUs+1Zx5uIaF6NeqigOlcTkUwV44e0ApNGvZhrdGsUXo6nK
wD9/Zfj7epN4rFz0JAMDyO6ty8Hktcgy8GosbHJrYGZR9D+MKSTaLNQz/oM0ZUoqB2rzN8Bkd8Uh
KDszAzqRzAJdWctOHPp0cowoMYrjNVSK/nFs8cugI72kr7XOuwrzoFvZ6Utxnx11RkAyuFeTWnAw
kHRuJz1pq6ADGRGbFgfRJY5SJZAuRRdC/O5rusPqarLp/1/teL5TFv/mCblTB5h52B9PMh8PFgiy
dEv7KjhA0r9EvT4BUXmHMUhKsPkgI5cEGNIuAuaLHPQ/cRYsWL6ID1TgEaCMR1uQoZNuuVR6cTrC
xJHwSgnlyESij1sphsnP2NakFUr306w1YeUZ9FVZAE8KuLnMeItSIUB++h8WmuQ/7HTdKF4mFmdE
gQLirUil8/LzrCvIl3qW8s3Ce7iciBAkktMI30Bdmc9rHqTL/yFLciu1+QyiTQyzG4GAQgJT1Qa6
9NQUBJsF5nIIu4t9xeC4wKHsRpFZaoDiUpL8glIWbwdBMXVG+04ZFdUklAPusiszhz8tCFvM60HO
M4y0p3FgV4Nt23t0uAFZj/ncZvDsP269Jwmo/x1MS8QOZs9voToVpupCoLLY3JekUzHt12RnUger
Pyb9TZPzmV8OUhhaVv8pWqvtI94npUqkSbTosWqrpavPNn603eY0Bb0vW670CmW5fuoWvTsy0PfN
i4Mz7oV+xmEd5HIXbpmJ9muuO1ZPqyxNewwn02fptATFd3Cubh7QeXLlzL7c3S3tBDFlk8ThcII9
SHHwHzsQnt9q6FH3Ni0CQ2hHQVaybCuuHXo7mFje56Jggg5QXgQ5M0TA26pWtJIGSStCoENz7pBa
2dugqVSPogwFgDARRAIuQrLiZVvg4/Z+lfSP7wy8oZhkRimPB5Rj1cpiPHgky1MhpS1/aikoXDmd
RFyY0LSiW0XaSakuYgUe/aN9O2tbTFEoYj5PwV+s4b3jzmbwqHqXFPs4utpCsiEoAhsOa367NRHZ
ZQ8X9A4f0Sx+V+TmhQ9uSdD2nLjIOHxQh0vtX+u0b5xuuouLs4Qq9lSgcqBwRyhB3bZZOsLCWZYL
mnin1zfSprPxqwg8mGaZtNpVAkuM1nZg+7tiMVOEfRmEGiJHvnNhaY//W3Z20GBomM1ELV24TY1x
17TG8f5rUVcMPC4qoD/VNyEBx4Oz5IUZD8nmSo0wP0q0yxlW0lguSLIW5PSshDRlmgHwc2Pel33Q
xwD8Fz0WE5xsJFef91aF0sPG09782MhqmsrY3au2SZTUYqi9B9uGHvp3/sUhaHB3BM1A312tdrgd
tmPIHgMhHp67HavzLvb3WpVpsnP5gDvJPR15mWX8WB06YniblQVkyb40y4m4d/+f+dD1gWUSY9OD
RfzroQXZJKfYbEnBVW4eqjfGPCXbl+AmVg53D1XB02F51s8xko+oX0mydz6NIcCrLbpGYEo+uzk5
n3Z1rGNwekpkpog9BvzU0NSA8DhrOnsEbZEzTOV+qHIh+ZWfEylpB9KgePI+j6J+90hKw3cHs0lB
M0noL99ULJP8aXR6VKJIuTQBbibnRravGrl5ohB6tZ8+TkMyeHs9nCuhGRjRE4JIMxu7Z8/JGpLA
vAUJSWwlbxy/P7pJlp0DbjaFbHg5W+2RWww+3gCeKJb2xg2bgCRraFF8IPO0UbW0CppdUH/b+fj8
nHcCd22KBL/ZoGXW9I/4SomQGMoaKcfT9g3X6POzEkY4Iux0CQSLKxb8cK+owQgW6JBceE2HKThV
gMjoYA3wR8D62KAxptJyvxq0D+TqGR8US/WOFv1fWIKahcmcTEPP8z+Tesc0kukUnLk74UaojmNN
LeBC2lrer9mZFyG4k8IuCEUi2XCPNM5G7+gh2udYJnnJcgJcLUfpGTltqImagzbAlPPoXEbC8v4F
Bim84JpbmVp3XB/OI+okgOBgyc50lx9CwJBFeuBAtOr2cMsd2+7Lpj8wYc05k7pMH7x2hYZGC2xY
bderHRmvjw288UPvSz/yLiTL/rBQ4a+k52izDmv/de8RgEo7anvkZZWrTTNDOrkh0ko7XJM0or8b
ev0UhgH0CurEnXddLk936gqblSSqE+q/3Gi8roXvcY8ClH1OBWlKpwd63RWhUQb51iZEzdsq8Itl
7KBwH0OVhjAD1CB9koZuWOfTC9RUd64itC2LbbrgY8eWcLkLgh8WGDryN9QzIu8AoQCnr+zG0MmR
xII8MDXtGFEltZkcdnQI9p3X4oPfALQ1CYVmzdZW6/pXDuPzX1tZVSpvVw0gZlnLFLcl4Rji0VOc
b34pQuWb+AEhFA6/anRR/Zcf9Zh8W4NY265ZU/Kgc7hIPWkdcNNKYd6jMkXXE7JZorgdRV4DwplL
oJXBMxngnqMd91F1hgUB6uOrwcrUvKEBxcvaCBuJrmjkeADn6EQFeWE3oPT59Sn/HI35GLa58Tlz
wWzGfONKsX9NRH86VBPu7lceh9np7OUrJRPlOe2aUZWeQ8c+X3kJiFXlRsGE/ikVOhRHhV7pC76C
U5MGJ9I+9ZaxLwW9kPVtWtvFSEdjmqcBo6VHWIhoK7fQBqEXWGPNLiVACF70itAF6kV7n3/HNvwn
gK+OK/RkBvXzBSMwrzm0DNtoPYzKlMZ5Why5Oa7s6yoA2Zb3X9lzA+LMI5xvb2onP1jD0m4YncGI
QRiCWnE2HOXfK1lRlFX8UAqCJCeaGfAr8v1Y36noL4HJc/F+u7CZs5uUTP971uW2Zs4g7XfF0kcL
UTiROZAtxCa5A90aYDXPGMlP/SD2m4LSED8Nkd2Rq0nh87bXYyiGHw7qE9NIF/VPCtWfJ9EJFBP2
eICj7eKY7ptVUdBLDnNDM0jbLW08T27kmBCnW+2lcW/a7j+kYka+Yy9/kJ51Y5jyJrdruhi+hZLe
6zKCCqXh1oS9CSnsJXxxUv5IIjg+zUeEDVjP2KS+FvfmVDdSoY5+sTq6fYXu6VDNNPEhEshUSyoQ
AzHXwccil0/ih47TBoNl+F6WZOkLPB5dYF/9fvgdxfgsQbOUex2yDDL5RP7jqTHYm+lRctApvJBS
DHu72p7l0usw1YFtIUVIHT39QRFOj6yXaVmd9oX7uqa4csz+NlbTUnsW+pEasGDn0UjdeT/edIBs
mzS8ZCGDYEPJXzN+6hcUFoipMitRR+PqsyOtKjd9GW+N6oC9+hqXrAYg7IUV2EZ334TPk3g1J/Kn
W5fX5L97gcYAAcXFJgiPevfc9STOP9r3COd4nHDqy/mU8F9N15YmE/yBp8EzqmIHa5Sblqyj9Isr
RRuebUBmRngW1cn3NrQEkZEDysS9IiHdUhNI3D/mx7d0JapfMOatnGNlY6KUusS8Vp26PbaKiJ4h
TYCi0L6kdYSIA6jEptK4yMejt55Th1Qzks4vxC88Fv/D1gwPtRaLqRtuTW0Rs8tUE2QhyNNej7zc
aznjaMzRyrO2jd7J0Zl2xXBmQNSVIBiYc1jH+iQb8H+bSUDTFoNWiqxA6t76e0NNBaiqk5OiTten
W92DLgW+HnsdC3eWOtL3+DnxGiNTSNLV1qa6A7rvnvAu6fgG7G9jFmBCh+aHINxle0j9V+SlDZU2
yhl+ZfnOQwotx6x8wMEfBsNPEHiid5cq29PojAO4v6EBcrvPrPuuRLLUbnzEs7WkzPCTgjEoFNUl
g2a7AUnPYPK60a2q5v6oOu0ZRat7/WYfCoqhvrR7VQFs14u4DM35/GRIhztIZv5spKSLN9BkpBlM
QT9Ba4I5kF/s/SFqBSb31INmBCQdH4gAyD6Im9b8LjVcbwrm1FUVC3lktCKVhNjPlwJkVvwoGiQy
7He03BPGlq3u64V7fwLWuRIFzVwoJk1xC5hOaSexgskC4nfxxUQjPNl7gnxtM6Lh0NbSR2N5QUz2
xh5DBzvPBPDfE+ecxtzItbRvc/EdidDIkima6Y8SGFk1MXdcrgpXAcDth9CnXteHeEaDA/g0NfdD
3j7VkG/MK0l/ODSOTql2gNt0qn4DUZPW6gf8kok5Lj3/N6Xw6C0crTSzcFGnwgwdCsClpNYmklxU
lZAhSDvehA0r42k+FFe9vJT6nIuX3t2r/NAlwYMarEjEHjFjFLZniGdKhhwzg8gM3akQCay3Aq6s
xTkPjJu5as2KNqeJbi0HXJSlRGeX0Nglswu+658w1dRY5FtIFctrWGFbELkdhbTAschA0CA5xk/r
CyOBnnhqIFTgY+htkjfzZC3XzRc4V6XOw+I9D371MaaeqwmSSzIMHx0BpgNAIx/MQaD9GHnzi79o
KBzrfdK9QVQT+oTUeyNCOMgQmzRfUnyqDSLxq7vyiwRC3BqQjAKscThpScNr9dqyBn5EOdMYQp5O
ncoklVEa35eBjdLIm76fR8LhudGOONLiBrS1XtilAjNK6IOa7DLxUUF+F2o9Ari0EBk1NEW8FGND
fhvPRVdzP4quaCpmwrqx+0SGnwDvE3GY7kgeW+oqXKQyD08m9TiZ8fyLYiguYqOK8KEL8yLyZNkM
XNWzm61GbKuC3Z7pu0z+uUMpKJ/L4Hrue6e/9x9vz8y2TPRDKeR3VFfkPw1cYYWWnAf6v83IBUpf
b7hXTMz5BGYc5mfYD1cG/RhbMv0HbY/Uf6/piZHmHd57y0AFZFjq0pE0cGYWdcZbn4a4tPSjAbRI
mVpiEbLtV5Gb2c2rMnryKWR2P6DLNZqbhmhq5T105Zj53TGHdKQ9Gf0sta3V6LSe/eBwHdeSX1n+
wd1xy5BCXcZgMyVE9P+xpk0D+ng6P2b0ximhhzVZvi+k5c8iVnLQl2f/4Zhtyj48SXMqVFTUMPjo
77SU0cnD/RxTdaOoWpmmiUqbn6EeZoGUNi/Mew1LELrSiawdNxlQxtCfLqXr+tYwnT11ajL88VNK
FvkWZ9GLqdLcySP9O1/R9omNOm18SeGrDaNh/Xc8aowZvnEHIBAJQNYZI0ws/0GK+a/s5RVPSCa/
1xsuDadXjLx/aJOB00+oDV4kvlYt+8aObUCp5Kt7xE+EYfywpcWZdJzAW8/ZKQX1nZ6CmN/21jqj
fsUdcsEilfwqSvYteog5va1RJtAtt1HwxVue1UOMFX1y8svOSFSRTwPR/O6zBn1DNvgaT2EzqscL
saRGNh8qzsPprcMx9yI69HiN4F0nSp4+AhhtbtlHJ4qoRTt+daL4q3N6BPKOM0YPLtw2c+IYwup3
K2CnsMNGVubWjlaG37xQSaEthBmkndrBYyfqIh9VdwKVMVqLHm1AOZRTKr1wGMraSGhYjHgWJOeN
jiomNTtw+R4v3+QTe06sokurB9zmjaAyeTLUhvmSKG2blayTyZwo29mt2vuoZEkJvXFwe4hbWvqH
zHV1pMhWVsv55szZj6AsfDgEPUZ3fGmNqjPFuq3yoH5550wjtgkLeieHvsnAcwg7Hkr6p4fHb8f8
WmF/VC9xTlCjyUX3hytPnaQw5R0Exy8HrICTdvEYRxp+ZUyHlWdRoCg17pBl2k0MdrBf+tNCpEk9
kbmZ5CF28Oj5aN9SKQTb3vRyzuHUZv2yWhwk2kv85wy9oWe+S2tIFaAQe7DVRVBZmjpREqEeSxRb
feWTLGKal9LqGRUC5Ik17LBiL5tbu2U+PKD1G/pGyT4QlNAEUYnXFhEfow6yCLn0JxAfmoHRBQ9Q
8N9XJliHslcAGouiJKUZNaXLbTRX+WzXLk+d1G1d0JnsUMJkSb/+wzeorXXB5/3aYNrX8N7T6YYf
2wlhUJM/iVDOuTYPIHnY+j2sY6vY/O+tfhtde3gMdwoihtQjG/t6vQWv5W5lVRKDdumYly0T87Og
PqjD5DCbxW+melXmfF58CWoQ609kw0E2vOemjcnZcRo4+hi3ZGih06UsODJpMy8BspQsLrt6AwwH
JTkFVFCVIr7kapkzqau4jhhbItEXMkd1HIpdziKVx3NqbYk73Bf4NwQdeb+YP3Wcm1ZpKV3ZY4HP
VfDsLt79MPVHpZiBhQccispjMqRQvBh5NPI1xlEWbaCULX0MxIoCtkKr4vP2YCKIEMn+00Xr8yLy
/wOXd495r8nG7FR+6m9zS/0+XplR0lmWuV5GGZz88rT2Y3M/KSRnFKRN4Z/zG1JgowKjY2fOII7a
yqFVgcjdxrgEbvUM/xl6NrPmx5e2Vo+/38q1+hIX7f4thXIC3cLFIPydtWiII/Y4Ln3/xBRBbRWQ
XwltO/ilt7FamWPBzWXVLcoj0q76Ar3AZ7tRc+NDoTTlaQ0pN+Xxiz0Q1HtEVP2bMGGUlxZgGU+n
lAUDR/r1ZXrMRnzjpbUhT2ak7QxWYQ7AJDYq1uYLf0JEOdgxgzL5ra3CjuFahxdF1FMrCk4cc1/N
bMro1X3Q16yGupxYHYa0o3ansBeG33/hZqpaUV4NQVY/47xtf1tmYwIvdbzLtkjPhD3llaCjWxlk
mJ0vh6l3z2SRSeMHOnlskpJ1sLok/L1ZQAz7BoxeZNcGZkIJHxB1dGgFs1r4f1YRRdzm6KxpPdDC
PqwwRNUuqB9b0CRS19lDSQeGL+eFj7+IWZrtj4L97cqhIQBG4o7BEtj24ndGF3k9+pQ73mMKrX8x
N0r5t4PIY0fi/gilegJXmBMNyJciLnHdhUnQLZS1MSL+1VMDeEhKXdZHh7A++IfDyA4bQxrtq4H3
zRhTXpZjcPK9cMD8ue1s5m3cDrKcqkVmzofnIfMS0lYlYu3lV7i0YnZx1/kkBnZauO0/81i1dsjh
s3fJTQjFgATxg5cMU0Ugm/Yl35vEd02PNOn2i+LbBkqcZ07cfi+aPOP34jDn6hP8NhAsSuBcYiem
dMvKOFuyGnHRrld45368Rw8HfPrae2g2AIvRDLzPP+uNCMSxG09ihRAlU0A97tE7pmSB8cl2YKw7
q4/t57mre+E1VJ7QvVE5Wt9W6b98vXXbcWv2N4SKgz4ajs8VgpKIryflrmPGw7KoWwFQY9SgqVZj
W9LthNaY9cET6GKS0kFW0IGWCQZyPRacgmg/U4nMWZ9YI2ybkkhRKV3kNiPqNRIPx3W40Jx1CtBi
wOzeUKyLlwLz5QTA5YxJ5Ioe6pHSy5hc03JmntmxMDykH50+EVrDUOR2RpFuvY/TopRb2mhBCMxE
pwu3weTriMsx5BPVmWYC9NdK5U+WjSXoYit33fYd0bYUuhTzSHUKfXuGuOuoy25zzuz7Wv7jq08I
ePalwocl6DkGzdgflbGr/4n2vYSahN2hQIC7IkiwaWJ8+rZ1bSl+g6FlxphstwVrzZ5fGQZdMYZ0
GA99Y3Hui7rMaHyn6imBmcs8HN0Hr3vxYjj3FX+l20eBftWwt8I4eREW4BqJF4rwFqi9TQT3BHkr
EToD3gLx2r21JjHw31uf4De3lNJ2gEKcqP4qD94fq0gjafhSAO1muiKZdK8U/DMmncan+6VfVOIJ
HIuz2eUd9Ra/hAoelyhrLEnsGrQ88Ti0wIKMzhcHiVSM+WN6e6jlzcgOBjN1j3nI4niBnokZHjki
HlYxo2y1CP0QX75//JnaVQfUSFeVT0MDOZfASiHbNS6M8+XY1pAIJb2PrmNZuM3XEJo8MYZUrWBl
t0FGkg46sPexo2Piph7JFmXsDud4WOwXPZBDwsiP6YUMvQ1Ip4/NvTYsoLy6z898fb8e2jQ8V7da
Gn4Nv+8+RBKS2YRJ8NFGeja0EgsJ8evT1WN4jooDdWjfzxfUH9+TyPy11ygJ4AD7B+sHP6w745/X
hJGDtQghl/tb93IXcxWdmqTT1zOMAHnKvvZePKZkVERC3/EUHrduD5PEk4g/ZjA0WcxvsWZcrUTB
janA7VUlYigXaoZu+SqJxir1Jm0ekLjHF9UXXYTf9ATK39oka/HWNmTKiY4enc4ta/wvrE9QbShi
EZUlWnO8E9Cn4RcE/E6BOO3QubBciAEkZQAtAbHQXOjIPo75kwB/zQ07XfIR4Wx3NngqnmdcJNzs
gr1M3X3mph8sGzZNzVYNK9VzhQZZdpeX+RnR4rKFJtZR9pIxczp9y235vd0fLI+fMf0dVZwyudo8
UP+eMW7HUjnv3xMlR+R1321P1MtczOri1wQVE9EMZd20IVCQwqgMtT06bQlfbjbd8WLTTTxAqUZ+
KdIRRE1LGHXAWseRUWACSMZrag5EpI2FK0eIHgq92wj8YD5LyEJGdrgWcuiGIUybxmkfPfADFdOw
NTLvC7sgQzRFofnlbMHP39+0bKemgC7nGJKC+Vj0trlB5g/IiG+nCVEZEffcOg4s7QmV5t3LPAC9
eKFv8q/grx4unamS+THwFR/lf95swiJyV1lvafEqmP3Kd0lGmfrnfcjHkzLrO/p0Tpq2hdE+3bW3
UO3rYb/Ah4fwlf9vhCSGSuVof/tYtgjajDXnZ5cMT4z3krF6di8xjWSbrJ4GNX6HBd65yiTJNB4/
R0pU9yafxImRa5Atji3lKHP3aqUjQh/IQzBsOkzuN4sSgTdcPzS73uZpoT9g/aokd67Sj+lvYo2E
Vr9Owe0svjflSn18ePvnAEMLTHvCokiRvONCg2NROoSoClrdHFflu4tV4ud1g0SyAJV/pWumJFpd
fDAGJDw19TaVTWjbP5lj7qOaMIe4RFssiRnXiFv8coESl+z5qWgAf2tWz3uSGzuh3Uw0RO6uGLzV
Eg50Hm6C6C0dwWCC0cMfJW+yA0+nCQbRpyIQWOaufAR2D4+uUBhZwQeEM36z3lo3SZ9aRnDrMMuw
jeSBg7KytvqbMd/g60CnEvMCbjSncyRIJM7r1g8C5lUttvWn8OFU6Jsv2K5fe/yZE4uYlgzEU1KP
PQs5pJ2C/nWf71ZThTnlKySJ+FQDnGK/KLTstN5s11VMuJFyIotGe0IRRHoVKfy9PklmjA7djeN5
58f+TpTOBmQMI+nM5ozRObsUwPlOoKskM93SiDt3KraUvuh7vjAUhNWLfNli/DJJmxXcX2iO7x7I
GePjpq/m3wTe8Q9MmsyGkXeXAvh1dNFURZOcyfDDdrUwc3J5Gc3dMgbep/f20QnV9b+7ADsd3XwV
rpD5rpIoH+VKE3vsehPIl1cpjCCGLb9jxSvJ4l0nGhYAXUYS0eZO4UB18bC/OUaujJhZxH2JL86T
tregvw0eG13zv7d554nRY3W7XtcnSdgJfU7CetsfXHWcInDshYgTknrb8JS/a9cOJh8pJlbOnib1
OPL5+tilmIJNG7GyBnJVHsSz0dooVVQRLRuU2DoC96PqIhbzOfhLwuegvxFzUIfaTfOwaX6Gr2G0
gzIMc8sUmjiGSQxGuhJJxzMxX6QYC9j/v/M6aBJRW+yq9HS3XOp6XPjEI7Vzw8KEZRYfJuC3fIjO
RqYuXb/WYyWXSjYhmDe4D2AXGxzydtg87zsEcV6Zsqh9OM9hbLUEC8tpQCz4LpVB1i8dxarohfKN
wUanPtfTd4MQYqvN2I1FWMCZdfAoFQMw5unfb9eOEGDmHdl1i2MgGtQT50xfizW66XfChNjbvBCe
Shv5VcAxsrWShwDrI46B9DIKQ7YEot6ROpbg9VR7CyAIi7tkf8JW8lJOQxzMkxustVhUr6aV5k2S
zTIqF4by2Z2SInQrkM3eby9CzSPXKE0pRyevtlRyx0oBRe9Zl260SApVqEDY2L0QEHdx6yLsp9r3
iewys06xB24RU+9toXgAGYBFYP3Zfon/h/xBnI95f8ChN53eDHO0sOwhBTL8a5d5PtcMtz0GvdEo
lMidKmgJ6kasq8PnXW4jPq+UzVycfqnkwz4WlC659OQYAsBu5GgIWlz69PWylbITBuuitD+xrSf9
2upsRxgLpbYIFjWjdNOiMSwaBBY4KgM4sPs8SKGfIfNUEpFQbqGriMIdUZr5POx4JErFtULwbHTF
AzCX5svaKsy7U8mWqdpP1dGnWqSKtg/mGMMDmge7Nt7Jj3yoCW19LJglpX92tYPgzq/Dgqt76yze
ckrThbzriLSbdaHExVSVhY5GKiS1G5R8K7i5VfNBOGrmeBqisZH8hs4wMo3jMIr63vvdW9JFoLqp
CYmGsBwrBQsQcJHI+/z5lQWKZ/LiacN9gv5p50OeDdp3XqzhC92gKH5nsChxF7FP43attw7p5vGA
G4Vhc2HIvv75BOZiuz30agu5LK3JyEX0bSFBws2lSg9ANIAhU72L5vHbkG9PiJ9JSIP3Kymy/wdH
Bya51/O7UnFqTnhJh/2VZ1Vn7e8QkGQwvrJMe5sxQGFxbOO2enwPW6kGdLrKAki8ACG9cfVuLu14
vqvX2UgOAoPqn40I74fbaY5kTpTcJNymf7Zgazfo7fbrxvnq2NCY9TJZ/wI2+2rmxm3wYtgZfwZI
1J8smG1VYoa9JezGBXFrChvW12sf//hvSU2DrpR/pqvNGSvEMr9NJ0QN/umV2IR5fUzYYctzXYpW
WmmDQlzcE600MF1ezoVuz8T6H1Wgf4+NbOkVikStu1M8paj8+yYHt3IFZPUhAonkhRlUOmGYTuNR
Zffx1iu0i8sOIqVtVWArCAv8Vnq2Tu3jAuQE+HbhYwYhWuONWVl/nyA2AtW5fV26J6b6JUiWRs2X
EhZZ0ggCKlHxoyyS9VPONvl3Kt2qEd+sSbxqNnWvpYKWTgq0M+WnABg7ADol/LaUznMwN3MFSSGt
t0sy4ubeQJ/+UbZ7YGPC+wLlBjJXzsoV8gXMJzoBHkH5DBgdwGEZElufNQ/JSPt3Ym0v7O3iBPV0
nH9bhPS+W+A/FoG3R3XFU+bx0K5LH5h3W3l426Gl2APkivGNCMHfDqYphvnJ9Do7QTWIVpaod4Ho
KA7q0r8jbrC7sH9alYBebB+CeWd5/h++z5DTz/TD7HNfOPXYu6ygmg0hl2lwKLYA4h/G9E2H4CKp
+UYrDRbYVe086boWdOX7MAwy8gtgqLJ9BszcGceLgzatTSXdobwB779MzCuqhm/WapgZA93Fw4GS
tQNkWfKT2jafgxk59C+ks/QOgjiXBjByvJ+ol5nmw/4SD+F3zDDaZBllFuCXfMNmxeqR2YA7e+Md
1aEeekRcNAnxmnYPZ6Q5FHt/QGBaCz6SluIxvk58vK7e3PXmBHoobLczE3Zsw8NBNlZ22Teef/i0
eyPP4duwl/T+/zp8yZGQxH8AAP1sDZBDKX3V37o1SyNH8Xn26nLdMdOcWlhEb2ZqgcBnfGYdK5Sv
i7QXON8vyKts1l24utQ0C9p/L0e+SSeAc4JAivlYXoQ9SCumdVsOZhJ3IyGhO40YARfBqz1U+EYT
MKC7k3GdGSlatZUsNtEDkWBYLU+8aDq6owkWwAhnEhjwu07kwhgevYtzo/YVAERyPqGQu03tkCDE
Gj19A0RPFK/hMqCMVJKfvGR87s7TqFk6vZT35frjbrhIezZUrpq9zAshOcv2PnvKwbfVT4MCemv4
P5cKWk1ZTbNFusbL0Q6CXWJ1iY8w7MBicWWjVNai8daRKCaSjssoUcegK3b8XRpiVBc8gr19eJbP
YwON9vP+OLhPbiicu3kjAZ06+EhXg4s4vP8ubweX3mULNogT8zTxcFm2EyY18eXKGMdtKAS1Z3g2
o7+1xLfNt30TaKBAv4Rpae17fGL/11y/Mzd+pddsnTXmVB9WMpDDuavyTXkDB1p8FpMFaQDilGF1
LCbflBP41sHcUUnI03cyzbc24PGwkVx7Ltx4fF3OLwUbZQpz7YFC7zG5WOOWSNnxIVjz5Sq/BbyB
eOe8QSagXUOKQkV+rkB9fiJsvgDmUeNZ0Yc7WAeraivaadusRCufcbhRfCCHoeKp6O0cHGurbHPj
F8QLbhfbX0ALE0rf+UF2C7wTPnXQYCC0BMjpBTdgfj9pu3UEaOV8bnk0hf1lKB7ZYETeMq6MRP88
H7HBJm67QqHYJztbHH8HMqCj95q2DSQnHERIiGJnSPyX5x9kg/7CkPaaQv5FzCG6Sa0jFb7hMcxC
g/JTpd3jlii7uspEQdi8hrhHmv5yaEIRlBdAtmCBrNY+Ghw+RGGKoYY01yvPD6vUT8gOKEKQ/+9X
PnDxptqAZOXBGkSl+8u9nw6QYaWcIJHldirAIJZi4i7W6CrV4a1TBTRS9pfbM2LSB5IxCvKxDfZw
A9MIXPOpS25MZ4140+knpCjZVUOi/mim/2HUMTmibnuoTtgdDBBDc2iSfgXK3fwwmK5a7+DDPp01
QMeCN5q2MNjDEkFZ1ZuVrCbU2NWAqYfial9fYCJImmAmwqyiMqKBOwsixRs747pxzeL+U0vdFjDG
ssyMgpKWDqAfG4MzuIwXL0r4hVgY9y/CpHaU4IhDN5TspMU+grWYjQNsfo6SFPBUTMYuzPm64xA1
mqBP1GkxNPNiMjn9dOPGJWCu82dG+6/b+SFmye+h4Dkq0oUwVgb5TA1xa1forO8oYQIwCa4Mp0qZ
gRuW81JUQwLbmXk6iItmf+OrxwzarHf0PO7EUhkET1SUOdhawW1UlFjC8uSzxU3UdFivSKRJ0KdX
VgHJkfu1joZ4h5kgR2uEBY9oox03Ol2mg1M+ZcJZx+3VI1oMMSP8KQHOC4hWHavGuzb6AFq/80D8
8KR7C1iUpYIUSnKhTzfGKPqzgDny6TcJrvJy5uRbn5L6uB0YBytmYjHxASif8qzHF4ZapEq99xIC
2/uELkX2w3jeRe9LZvW4qIXa7qTvVZnUqU38ZqAYh2dhsIMjHVxgAeHB5tw+qWFckrQ+A5hIGOsD
Ri4xyYwY+IRyTbvoyS4NC+TWVK9bZA2TSSbvgS1NHfc9vCrSzVnRqCdDOaoQNxeNEiXBDtPxBRLA
BxV8swD0rPMVJQhmxe/dJPXIcomrRb3mBpyXluiq+tZUNv6a63V5HZv+9T6VCgyCBePnfcP7DsU0
22XG3cEmefj0r6E6q3Lzybu6FvwOhKzQCX2EkxlM0AC8kkE0Q4cUz94KreeUaoewOAZlydqeFyBd
D8BLPetsy7EfQTwhH8jpY9h9TSJwNKXeG6EkudzVfuDMuPQHGvYNiH0l/YjWpv3PEMN77FwP/Da0
AWJ1pkkEFgJ+vb9LVGY6mtDInm7DhMFQTNrXZ1EcEcd+I4PA7djS7+JIPjpOVzoQwnq0vUF4R4u1
2qzTksp6ncUxde1jPI3wOxBypBHiyk2TLRte6EHRv78NBqnsQBM180Ssbgqt5dp5N3rHUKegnNqK
47Os0Qultbo2XThnbqI9kj4DrxY0CFKdEOZwqt+85XR5Y6Nf+ps1TjTXvBtFlnLnUIkRPYHNn5FW
lgm8OYioWFw1k6T1R+T8MCKZ3P+TSvSjO0vVlyst1q+htX/KT7N27A31sn7xF3z9rNhdxVlKHnAa
CyysGnRFhTOolop7cF6OB0Nx97oDIfGPAfeOcWgEkqLztTvHM8BmR7vOv4itleMnXy2MnyUun+PA
0CCHu3suRpDKTO4UIfbzmc8kQIVt3MEcxbdF5hJF3eG3cVtZ36gMNj+yIEMnaBnDNkUVUEEaYKjk
ymKkVv8J3/MFw7zsBOTNGtJVhZjEga2fNoXDMfetv6BnMen7ccpfYeno4oktiHxn9IidLJwhe6ya
pYXDnU3yM/CAm53U/8DT7TdT8KKPEKSvgSx859QjolCioswptvfS8uD4PidRWwpsmqUvAtp8MgOr
WoDkMHdhIBIKrLfK4xdUeEzLu78SxvVJ4Xb6KENqfu1GwpvQTLYubVLGyGFq1fMlY02l1AyMN7n7
KBgbe9jxpRKYillXPLLj7O1QuKT7btshUHuHKHz+hlmAl7xihKgFs4I/9Irh40Lham3Vb5GYuXsI
7pzHZSLYg2dXHOAYPH2VqExKXZUXMO/VNs7qBXnN/+RbcVxxC3mh+p4iEdjP4E7nA6ikXvFwAxBc
g0/omqrcWjTKyx13qTrHxTPd3yKF7SeksgjM+DwWlm3OPq5Cq3AOs/drqmf4gexo9PrA6uWwME64
qJC0EU+5o3hgdeAfS83T79mmcWDYAp3QHH2M3Tsv1n0Pqt13aTW/Is+dTVWK2KHP3aeTIEGBzX1F
6+HH7AL/wALZ1QN0E6DBGKoqum6VYx8guarK7kq7wa06g+al2Xi7UhOSBTg0wop0WKuk5aApDs5K
aDx/qNGCxfiFqbRSdr6wIO+EGk2j97uEhd2Nz6E2QtocHwr5BBqFK9ENeNn0ZYGYvbecaqL9Qfgm
ss0FLPHV/0bz9AzqVzwoFz0M+99EyNYI1HUJg3jrh4OpYmoA99H6FqJqPplcilVDGOEDvdf5Y3Oo
zaATaHay7NkOa+LDJgI32uuh1HXs7Zo+ZHMqGmxSAPPUbHUVhXMpkIKehoK95jsBsQQQ9GUXDTt/
0LBuxhJB0rWPjv3g60ZAJ3Wob96cchF6mXeD3yi0LSDiH7g5r/UZ7CTiXw0mvZNwEMnVX+gIMEAp
TVOCEXtw8YSIF20ehZb6g5sFcd/jRhTljid9AlbNSsO5708Yk9zprFgsTTCHRB6/rb0HG8yFTYK8
Z4ya2nnnaMswnBnzreXFCOfwT7oT5vnsWVsIKZesQyCc6RV6zdYcwIlieYnjQmo7Jp8yIyIPM3ir
Ml0W6K68fcjauTSl9SCqaZfoNUwXUZxyManHbxe83ub6gbnLVxygB9Dq4Lx6kUEJxk5dntP+sifL
Vqgxt5T0XvMRUj4GyYX9Gz+pXD1Vc3q+WNHdPqwRm9KODSMmqRtzwbgs70kswTRMdJ49OiGJ+bkv
0o6+RzJAfSu1nv19E4wJYtTBwShZkPDvJLjGV3/EAto+hCmps2pwOJ89FGRVWgbfijk4g4FLb1id
z4TERISW09cwFrnyD2R+C88aj6Ca7pOPKx7PBP/XDtjmeUK3q6Iibr++2g18heZv71PJ7GepdBzF
NIm0oQZvwtaFcB5j8y+l4BV6rZZrjHTx3tTK44hZdyoe95CEVHEm4AnojAbrWgBJHqMMwkKrncGG
jmaTl869T9ARcoxenpMdBvdbFeqpZkb5WOZHKDU7GTaChPyl9t4aGzUT0BQi6fDLqJg+rsv7GmwW
Z6nRaUMySQ5OGRSkdF+I11+XaGZsqV/AOUyQs0AjBKnlwil0azXhUakr69o9uv9zyXpwrXWy0d2i
zDSHV2McULsWdv72BNhnpuKrSph9pOeZbpUMD4leqQZSCpw940M9ws0VuEIHaJIGy4PUcEE5efIf
dfO8AuOi3Sm9U3u07+Otb3wgvwvYNsMDBo1L0JNm1Tv8GDbZb7cerzt3C+2W4VgWEpRbQ+PxLeO8
G4EudhBHl8xf16cCBTZ8mpm/EEcoXeMX70OoHfy9vg2L3NC6NRgzKYrotwruvnad6lprg1J2Hw3q
QRRp062npy6WyAKSimA0bVf+YVC0d2v4igWqRNhythHinT2pA1m8PPUn3/nC3N8k3AT47RNXynTf
1i1hqTj1PBcZDh8J6Morl7NS7ZSpxogzfo6QKYpQ+BNSYe3kF3TKf/mTlobTxL0bsf7/tZ7t3JnK
GZthmrzk/NroGcwMGHshVFU0Jtx8silf+pMof0sYLf5VBqgUOGjP7NZYoIzubvNJEc7sxgMFqOXS
tmJktTgs41zvQOk3RztIORYKnDqHBCZM/UgmzMtrzKuDhbkUT6MMdMTqaknz21mDffw09oE8VlUf
UvNymXhZ5ar7iOr2YQSpvZBWSWD3d5xVDPHmRYNWbelw4Hmm7JM9AxcpZzLvdneUtaOl1+BsUnvs
ziOboEsNehvpbDX0QlBLEcQsc3+VTk3ONEt5RKKi8qMCY2z1xCqZY+xbOJ5xUBg7Xz3SKJady1rj
YJ9OSig+GfxMUiDl6Kabc6wSJB1Sl2oZJbV4YiQ2MHBWuHKhNyd0p5rHTW+mcWNYPPg8zQYJxY8N
GOfYmQn28U8ViKOh8fQjofVzBaqNTqX6WPaKk15GU1vwRUlhMmMUc7ASmNvOTMKa4buGzVcgFUIJ
xozccI4UfulWDA2YUV8JRskeHRWNyn/4eicoVOfdE6HMA3oUCFLzXD5oQswAjhHfOO27m1Dd7Bsl
YGMUgdx4SdHEDVADOD9nSiDR5/SkVHxtS7nZ7T2cHYsNQg/Tv7cKOpKInoi/hg6ILw/Z0T3ravmZ
2zmt1ZsA3dLOS/rUfbiRqiSOQH2ThB7Q9E/fHhEwGqNiAeDuKnKhDWzwxsOBunHAktpxpPw+nEKN
GZEY1SXq/1nnAcEf0H/OWhWuMmvt5+QNFxcP/5dLa1vyFiRv5arZTcnhn6JjlsWFeUo0UYcsUG6O
p76aLvGvJ5qks2d/MS/npBDCk51nes/U2LiiBpMvXN9jFdj4XYlkDPK808YDR7Os83iec9sxWZjo
+10qWipO2b7cMKpg1ptdbnkYcw0RAkTOhhz8bc6GPkBakm1vAiSRVrlLCs+hq9HXvB9alxq/IX48
6x+ZC84Dv5lxbRsOErnvJEk1dnJh99KXl8MilbXckthhPR6nP3FD+2F0KqRL89Bd69SGK/S6fAbP
E60+9CULaZka6Rh05rt+v4Mwv7S6VdFwM45drG9GCZS322mSYzq+Dm4m957nAOBHIlv1M41qD1Tl
s9RZC2sTFsJQJS5Zid8wEiwo/4/ix+aPomWJoh7yN2++w7RkNWLv2GdZzHJIg5Uwdq/K1v0K4Fty
gBOsXTQ28pZV7YxUuG+8U0kvt0nR0yrkJGmNr/mXCaL93MndbQN/8DsE5tU4H+i5q2D/ZKUc64Mq
bULac2I1mSjLAGAJIq2VNOhBd8yhe9WJyl/JR191m6OrOIqWIVfvr52hpJOz+mG8ZOoPzJ67lOpB
rtEcZVjfPiCnpRNPCpLeIm0c5gBbPFV+5mK8gUgxDn/NJyWvG4M7gpB/aWXcBFDhdZQg6FnlLKQl
IVyumi2xFaGNZLVF3vPCKXq83j9XgJ+G6+vsk5+dzbXM8lH9YFjDmEXyNiGvNgnTTqwrYCnN8S5a
jt0hlKKeIDAA+SnRaBcsCAV/RvAKa1U0xl3rlnMZYS/nxaxLnndPOkB36fNKZr11kamCZ52XR84k
ySaU04kI4LwgGsRjbiG+sBO8DkA6bi4S7u0+cFxCxNXN73ID6HVa8M7461wNXJCdgoEF6POOxqde
O6mgUc1JJ0Wrni/rWR8vMaa1Kmep+NcRTuRiwJg7/KRCbFv9Ia3vwVu/fTfXufMpt8s7+zZt9qXd
QWXfx9NuV0w2tYVV7Z8271oqVFprsFtYNVOxHUx4v6/qjmUnFFNjxUAFUNPX/1bPirk1U20hGt+q
A+Sm7bY1yfm26HzRJy/yb3w4z/WBp/59qkjNKTun1YpBiKSqi2Fl4L3+2hkBHfTF0mcODO+2ff2o
a+RYA6gLA7XrFOb7+zPsAXfSZ/KvkkJpsG7o3xVHinyGbSeZrMbEMOZj7z82+Ds99Wdxl3YpjLY6
9T5V9fo0b/4JprsvAOxMGPu4v+sVyoOLlTR+VyF6oJoUrsQefGiM8D7h7OHMWeazINVehcYClO3R
9XJBUgve8u6nVa7GfboIP7jFBnmyDmzgU9wcqtXAfetjQU7qCnaZorW/BeFL+sHN+vzKWahQ64is
mQHqAty22Z8vS5WsvypD6PCbGEUqAtkggPd96lx30PeTNmmrbJDG19BZOKYg5bBEMvBp2ohS5LAJ
312YijLzjuIiVB0N4FVJcKWkD1zOuAbR3Gdfjg01uwKeWsWOD8Ny7GohWbaEWPvvy51rNS+UvNOc
vzfyossa5Hw79H5vCGbmRQe94OzrwOrAPmndSLBRIl+OBSgAp69vRI1+zvcDTtNUzbmwxCOyOQuN
Qjjdn7eaNQbv3JbI3VeA0gx7LpHzg98j7W8J79jc/ktlpuJlH9FgTFIamic7ltAMCC5RuNUYd///
MB1HVZQFaFtairSnJYRyi0Wtt+Sflt98GfNe/HVBO1b54YGjyXkJ+P+d4vN+ggM4nQn6N9u6OfZJ
F6LAEz3G253uh4AujNQoS8EzZqBzWlhVU9zj61JRtRh1+rGKWgz+9FqYTs8lGgnDet+raduroKJe
pkqv9Z42o1Hmf6NLqH2+BTZxkhYWf/q6BZgi2bFkktFnv54fbpkk/Ep7wpiTA84z4+KC7wjDGrZD
X1HcBbAHTc96xYxRvFg/BCTE1G9OgMeLu4rqiwMGakYvSKeC/L7yMg2DsPRwtZsl9tIwHKuKTvcu
CVTb/6sAYsvcEx4oQwI0rg5ixgcPze5KhYhyWCVn1pjHBgrKgKmbRyiRAqXB0gt128J3G8ZUF9+H
gNyAfvX+8rKBKWE0FHl+5BY63FbF1UbiWGxj5znjyh6/mZArmPjItve8BdbpyYI7aPxxmmNNr1AW
l9vcP1iBVUi3kDaLJTs0pLVl4uRyKYSpakf3Zldavu6kOFtxTRJt8kBI+A7TezZ92qmAnAc7l259
n/Xy5scKrCXVN3Ra3a93ko2Faz7lZSa0N9JC5ggbEKkx0PT7M8pFL+3WovSwec804pJP2KxRAs2h
2dqrfhwIVBblhaYx/ms+aDjk5/CC4hS6zI14kQmf0kyFJMQRPHAQVzm+NSXOsbA+BkBrzb5iBJJh
+CAIZvWU7sGdDc/e2WkVDi0RKt5hF7colzZLxo6/WJr1OfRON2IuMgFzsS6r6JcD6n0P1/3+KS/s
+SSyOAgDfnBP6bYtsKx+/GRopU1euNZ4xQ9cbeONQr+smGMCsuQISy6s1gmm9Pr5F7PWGT6+SLHA
tq73dQOnxzOcpFTvKkdyitt6ieOL0yrH5FiFhvL5/68KeAxY+eXV8oZiqJPXXzIESEqDySpNvQA3
KxzOdOXVfRbN5uSrJvmmsqXgLDcTiU9p7VycRYHsIU3Z/CUmN3G6Hvz2a0/HNKjkJbxTGtAlLMvN
uPTofoSFqQCHVgRhayq8B2Tw0QrJLCLjCGtbOQ3YYKK23F/meAU53NhVbKTkxQ/Iii1v7KvF9y8h
rRjv0P9Iy7T8CIrN12mmrfO5KJA/mPR2gKaOYPPQX7rRSu8I7xc82MKNvFvxn45ADMmpCbqiwUmm
Qo2a4um96Yh4bRkL0qsuFiuMD+1XQe6CWI0kCx3YsnqC0R506ExefxHVU0IQspdNdahIT96H7GLM
hJmZzDhnejvGPz2bM/okeIiRYtFlEQ31lpMXONnFYBfK8YpfHieHnshpMX/FtB3PtCitE7Uq6+1j
TVOLBFi2OTXFvwX1GNw7vDsmGz764yy1ZHjYaj1Lvx5pSg8mEcAkrCGLLBGbSZ6OI5jF+g2clZUU
YxojuQdaSpG5A+WlsCvTwcKUb2CKVfFNC7kfjk/QauecAcezyUWQ2LNguHd0oN1yoqKwm1VIc/L4
DWhgiAFZ/MwkGmJWg1Y7QSbyBnCRpSlC+/RjyFvyOa/q8Mk7kRXbyffnaRO9sMgOdf01hiUokt7o
oCOMwXvLFM8q3WE3J5GW6OCyu4vTZZsfl/bafXjCE2Vzk6V+ELzZ7HQP6+PsTWxWIU72YW/2n1h3
rYP7yDqDqpMWWftQBPVI+cIbpy8Xrnks0t3T4aV+QK3KZBwqBxzCwcc9mzi5Z230BiEoWfBIloZ+
Gk/dGEaYLF0kqemzba7Pyii8MTqbrnHc5gMcrCc5zZiQVo2/eG56PJFhhqmJJH+tDq2KGN8J+al1
/ASC1rj9Pm5mPiQM9rDGoWL+E8c+M7YgAJdfPUclYmPbIfIftb5eXfBcjuU0LieKo1sDHEUbXkQI
HKowdHwe4B8KbDyhwSSua+h5LNCVasmtqpg0TnZaxkhIepOYSJZChMS/m8EmUB9EbOkKIZ4NOIcY
Rs0oOkAZgJAAx1h5ZkAanrH9hHlNds2xmZvnKR1tut3WaS5pOZnB7cXUS7Do+mH1p/w6i3LZGcpW
vdGG1QZ2fYSErg42OP0PDpcr7oeFxroe3s9X8KRn9CF8mZDa+1JDy1MHJPAtZeebU11AMOCbSRYl
KqZ6vMkaADUcdIQhyEf3kFvMLQ8ertbQL3kmRBmXL/zOBr8GhXnF7JkZYQac/SVdZMSiFE0X/+51
5DB5gG9+91ou+VQtC/JdW/phaL9cz2cyGVMucxMiexjj9dxPnPgEuouwryO/gUXTJJwWQPhs+oI+
MvZK5+X5CDQ/VVgTK3oZ+cFEwqWbBnYnFxyvHAX1/ZMvXoVeLPBRd/J0AEKprVWvMGH7SkLzotVP
z3rThMJat/Hva2aJvR0+u6sp1a6UKYe5Z2MqQPlfkkwhLl21+C7AXLRGt6gg9mCDkDT+T26ugHAz
7ja3pZWoxBeGiB6C7axDiDk5neruygCTS9SqU9+pAZRzG3K0ASXznY9c21ctwrSaLI1oHITRMnvp
ZOgJySm8vuGeCs7b1iDhqecy2hoHGMhBe4XLHIO8MQoDaM7F5nZlHPxAWAGYpqj7YVoKjUACsQ0x
15iM1E33mnqSTPo0DiYqFzdVB/p7ppxXnoL/DH4FZ3pqFb02qi1nAYCkD4FrmEQLqO+FYm0TjKwn
+g5rMjjBb26A9f7LIZSUkAemHr6bo00IHwGSW1uUoOyijUl6vXxN+4bg2B8OSbPd2ZVNS6T2q+hy
MzCRWGA76CuQ9nOKm7VaemwfBKxJOjuYz+tTrYv9GgCiarMq02T/LJUC4rxM3QnGu5CtZps1hQND
aRhEKtHHezHgExAAvhryvpd+oin6KkpB6dPIcQh3p6plsWnnsI/xz9cS2Tes5hEfwoCqXu0rHv4O
GaP/7pnWNM5NZqXIfDMTcPNIe8MsSmsEQrtuHi7+49MSC1SNI1fHgzh6jjzdTILcOJyQn5z8SuOk
Xt/7XQ3pv7h1+ocQGc1iTlKI2vuBC1oc5n7v6GQwTo7frjsgsFR6tefA10pZElE6TwgaocZLqiDA
EAf2JUSOkpMeZYlUTAHDO5N8JoHaDlpsXhtxu3mNzUxs5qNaptWbY/7cS8GFzXkF4OflWzoRed0k
fjQ3MpJQ7QEpqgKs9slvvjWH57fN2UAG0SReA+WuPkZ32koluvnFw71+rhmitli+eyebhQdvSC0l
XFmUM4mNoOG8em/yiaS4XeFyXR46/D1L9G6c6mxrAwCVOnyQZeaLtUQ6ZEqeQFl7ABOz/QBh+iY7
s5pG4vEFZTtlfp1jWPqUM1O0p7UiPuBT9v3FSVm7Wq0IDmUrPR3rk28f2Z1uuXAfeI/X4GzoIUBx
ELz8253ZqxG3jiDsRVJ7ijh+Wq4VQ14delEdpL9J8SZ/R2IxgxeW5R7J4wdseiBazb84l6ITIloO
tuXGnSj8migL8ZqD9Pu1vSgo96twdl9R18T3aDCozZyfGcnue1thQqWsSwl4Hw55zju+eSzkNYVy
DogP8bEbYFlEhlJJDlN9slid/qXlllIn4qHAMdcTseQu7vb7aqeLVzoj0SWqIbDYdQ0kT7SfsyCW
UhZTAvAWBvXKEEPTo2EN52gtBrRU8+XySgUaRWgo4683gFD5knWJG0MqUpSsirEf2VxzLSyoen0Q
E2/uGHut8IfB2cPSxxis4oJZPqjeI4Mc32ILgpK2W2Mhzk4SbnReJyso1rEgN+AlsTlGnO/A+gee
ob+phxrfnME57gysPL3FOLR59nlb/W99i9gcLg0FKjQ5TAheFrVVoXT0baZQzFg4PvOKHUtmv+i2
tyvlcWQNYuoAcCeh8YXYFtObD1nzNoumYGIMDsawajoRdJY8RzfB+fdZbG/HsRhkUNLRzOm0NSIB
Adm1eUGnjPvutnXU2g5I2jHMUw5FnUhVVJkevwQPDAOsj3nwOjEA4/IXwZTcFqSgTfTmKRK8MZ7S
zDfR2mwyhTde4v33dYK+OXEuuNmheeurpryVS01gzqR7FYjTCgoGzLDhzSOdU/JIyd0sDNz9ic92
rFdg3iG0APD5G5p+2MwClATBRNg2QhiOdHv/+IfoLYXgIxFF+Ocz0OmGgc3XFQZy234Tg/l45LfR
esRaaXblaoqD0LUTpwXjKyK63m2S0HoAO+1xJp5BSXhDmY1WwZL8rrvqdu4MTUiwVE9W18I3mzZ1
uU4GpiKYi9gkt+rTfgJk0Xw5SKSKDrYKhfE3ePppXMqg3Hf/LJs7ij+KprhgN99ZsA4K0SpuDJmN
b+fPKQvYG57ctomSJuEoDE6yZt8ZG+Qv2zlb7xwHPLsj2vDCvO6C9FhycLJoo7FpyR1amcAjghIp
2xT0pavWiJ2u7PXONRicZofRtXUDJgOu8ZEaWu1Mue8hm4N/POc7LAmkZVjSViIf1uv44SLHX6OI
VHyZ00rRWvuaOPqM6Zjx+3unb3dYn3/ZLnvdzIIjrdbSm5LufGYtl32KUkql/BLrElV0gS8FOQz1
CzZNndpUcyjlKGFPjiD5HEXXfPwVjHwr9eocLTAGxtExvlcUeU5lb6TMrFGm31+Zcoqvqvl/ay3a
D4RYmqTensxK0afRYf5dMykfHGsOGbEKWX+jngr9R9yv4gYdBetRgC2VCAVQUWJFfJLvDKCnxIXN
czhmwa4FIBgr+1MHZrwBRCtZZ/KJEW+zSmqDq5kxIHEou9ar57vIilB73lnZCUW90OwACxLC5vmW
QRhDksHfYDZ9cxzN4hortg/+GcXxJYogJSSOltIhIphiDjX9OChqzlEyhlxVlF8gBmDBkKsv9ooV
YMM/KxBJ1YX6pePo/PyOr6kaLgSmuQPjgXd/DrnRJRuSZmtwifKAXzMwieuOU2x/xJtvYhs8cQQD
EUcgtMYylL6uGJmzaOs4e8HNN2aPdz+H5D1+z9x3Dg8e4/NXUvOF0isf1fKmw8mCTiCnqFVYySwR
zvT3n3NElmiouKCwWCzjEVBi6dhAJPgd6ZiLwsqMFhyhR1Z/Xi4LgYR6tscR0XRn46EtMRBW53kv
3Yfc3RP1qwkvxMppuoH4jFRjoNcuSW69toyMKMIYaDzXiS1DR2aaeWluPT3EQvQ5RBg412q8G6nK
JxiS8ZGpvXMY/UMHZvdyQjOUB6mzyles+QnrC541o725Q9H9FyHgmSNUjciQk8HyoasdavJrEPf4
1mVNq69d+q6VEGBJqz1IVV/LnpyXNRdwsBbCR081RBS6PD1GvUvLYNgbDVDYTxltRjYuDJQKKD8r
mpYHYMBunGRp09NcnBlQBEehiUSSJIx1oKkSmgV/WVXWHf7vUmyQwqI6Zs88zXTXuAJCUEFbxBI0
vujq1dlSXgWfWCCGWsvFOw1vWKMwE0TCKjwKTSVxjWqmqjw/e1/RrmXxnSr+uIRST8u47tThB1R1
8Gs4Q8Vx6CQwCQ9yvECxZQbtf5vdgolA799a3+G3ceO7vLZIqD6lIOD1Lf9D15FVhuHxz3bjEPAS
IK0KmKEH9oG5XNPZ8EJ9EWZiZCcgel0TVGAb9vK6q4/GYp4UFNozt5/xy4P8KW4+yFzB3BzefuxC
czV0paEb9mNPhuKOxU5BvFWqZOwu1+JJtAJjgm24s99ehPk5tLfdAMuqt1uYxUCgeUC5paJrm43+
Qbqd5+caZABIZWGq/EyHC6dTDDVooiMyS7jc+Lvz/Pwfq/CzLkC2OU8jiX9tFEReqYlpByPJt42F
MO8+y2EUKONMEo7x17Mc7/fU/iiD7HQD7Tq55O1LYzcEqUqJxNZ81hEdVAKZaOVsCSzJjYnFQ4Nd
z/8hTyroqzgmaHhtSJiQ4STMPoHKR7b8uhQrx6Qm14/FAN23+RVl00A4DftWIJHgWzw1nfiQh6X/
sFnUv9bviZRRuEmbz/Uwwf41pqBcbztSXPzlLF3l9u0aU0/R4//amsop4JBihiwSfzSbEdT69/QE
shXWzwxkCPEGU8D7vElALQTMXZ+GGGMRAHURWSQOK0u88WUNu40yjVkxVzIYqCH8IIIeDNNw2xUX
zoidKd89C9Vo31vN7i7l6bZpbr/8s6ojgv4Xikkt3BHTcnugiFyvjRWS0bwU+OjQsBqNKeahi/Yz
UKO8On303XL11aAOy6Xuj+4MsjYJK7Ma463RjDo+ePmJzvkdwUF1NGeju+puDQeBu8lqcisZ+Pcd
YYxX52U35C/VMVOxj6xKl8/MFsV9/YlmQNwVlE0ptSxDw1xWLqdSdonHP+4VpK2BRqs+wH3FneJi
ML/YH3fvvWQ7QNfPG6DgwGLHAAzQApj7xv5I4NtR89NqLE9Fj/bhywLDniFXVdhFWiWl6sjpDPhm
TmQOcpJf77V4ZPAHHapvFRMQTy3UIWTyvSmnJHfiALU//EHJFBgRL8N4KTA8k25K2zhbMwLB+I6S
9A9XmzXi67/3VVwam5uXQry8FVD6lWrGXWsw+4TIbxj7iqXj1KxOwSlnAmF8Pilx+mSj/kYLfsX5
6re2S4E7ok0GEC2Q1xxt9y8LvehnMKfa8lYJoIuXq6eGs18yy8cLn36dzrZZY+CYIVtbj9trObTc
+D37Mk2BbJz4tzueep7byV3eGZlfxkO/pUHX9EFuw0d+qMZSjfmI1KtEfr9Pk/j39BU6K4ovvX8d
XpNGEpV8da5rOVSKGEu3jq2ttjg4mzbHunHsA9kKHX13QGETXVW7foo5dhO3EmG156nWU3r0lQqk
yfej7ZPQFDcmvxxI2EaYMQCzul1Rlv0kduuOnbaQhWq1tOGZG23LPlODupYgXIhFAqfSDIbn4Xyj
RSJPzQmsCSKkHj+SeKT8Y7EKud6M+iZHjp3x77v55BLeJosYMy38VHydP7ysfMFm5bvZQKkeUHet
MPxiJ6WbLQvxf+75xE4E1s28U9L2BZ0WmVUCApI9WjINuJphtlabWC8ykyI7brn4Hmk7PXSwCvAy
3iTaYC60mKUaD6g4umBzF1utv/v1pyGZDFabNPJwpz2d0FEUQhzeeAiAaplezKiVcBJpuuXhhrQ7
YEvHwaLIeMvY9PT1FAf0E2fGm4dR/FxNtHlGeO/UNdn7gtEkxJs2rUmQMwIiPa+AhsiQh1L/MPbu
CbpPefObcqkl0j23fyScvUvaCKLS3ZAwmyB8sDkxgD7w45k2yUGxq16FcVKFedf32aNagh89D4hs
EA9MqLM1rjRYHxSBHyjGUYcRDaYbFVXkmAsY1VYK+IUrl6tq1e4wyqnqjgVALPXyaV7Hie6DIr89
7G+SkQSnD72KgByPIYmZqL8p4iUWcixI2IC8blmelO1LkIllfLhQcXbXr8skgEJIkpROR7VlzLkq
0Ovx4HjUt4tEr4GZASKbIKHAKLUSZwDE0i+VbjUFf+09x1Jw4kJcNtTzZBv5h4q8H6tT6MUbplqA
oECDXQ4siksJBuYS52DxQfahqVNg4YI9xzbxf+Oe9jXSdWlD6f6LoAbPLb+V7NdNBUBXHwA7Z4v5
Dh2uRTPsb6ffbHyXjhysQf+8U0v5zJ4jT0Wjgj8deD9Sex/zNCdn+za8QW6noLK/FvLxU1dE5aGQ
kuVrGEpVQPFtCDDPJ1v1AvIUSdOpNyPAHMLfBYULnsccMmX8BPrQxQs1HZZu4Ey3Mc7PzG9cA8PB
eD1JjJ0W4Ar0SpVwuOuD2Q9OBXO0hfZpyhCQYGWpGZG1apD0FLItm4CTERlJBMn7g5A12kTAXkyZ
lPQ748SNvx0dSqWDekGY5LiinaBNW1l7JAzPSVFFGb+NWNR+WkoBa1ivRWvOicH13OXxZC3qns3p
VTTe86YLuOH9H/FaDU50QSsgepwk+xfYEq5nZwo7n0ORAUxDeBZi8KV9pd7CEN4nxZt5X9WSD7cv
/CiuWhQcQxX/NAe3yVPH9/tbcGgoPRDvNuu8t9JaeBIMgRU3cKL/xXHeaZprGCx7JF2wfr72vNHC
36nxadZX4MJQD8gFzt6QzAy8Rbg3CfaaJYr1TEyrFMBXMhEUGsUgR0MnEU24CBaDpVDoEcr5QfmS
Z+Z+tuT2wDICRj/TKA9M9/+6FqLkx7mucuox3QMtTRAfqbpjOFAb1x4LjA9hJtVZ7+3XyDCB3NRT
WvjMD7D78hGQOA8g5uqgSbvQpzm8e6+s5gwkDWzbUZq2ouEwsitfflLHzHgunP6Jv9G2b8uMHWFe
XlLbH12mN6Gkyl8p5t6UqQ6MOYTZKc0WA+Tk2SomxivM9TH9oqgCSQsuDk5SMd1KtyXQirCR4WWI
tVo5Z4uQFR28P00Y3k/fq8TniAoSyqv5TMi/PYgYDMEXtbQBHK4ebzSSFAu5CjquKAneYlmrfBT5
NH+4LsGU4UY4ZTqf+LsCxAZaBhVxUBiiLbbBn6/a1ZnM0dkSXiBx3eWIQIwIvpHBfLj4QjFryra9
5WsUawPPeUR/d4JH0G3g8AjefWHinqLZGnBA8wzKORvDCJZVDraprVpMlZcCzaUE/3kUhEaALmoh
pLFbfCfj7rgNl4q+xMsW/O+sSGqQzdStgLPVAR9U8XP3FZ/dovAz6Ms/bmVhhWmr4YeusigMX9ZL
7pvyIHZ41v+Pbbp/k4x9ROTZJUHoGCfjF4vnEeJLLE3O+0evwFFYbuAvfUV+eSg6a1C3jvGCuWfq
wO/lGdRyVoCMeWQTPnudT2vyfJpfubqDR4SI+Hb27fZUYNBrb0cTjpBOqyN4AwdeEN3sRXcSvOGM
DocNF+op1pTUOfg5a0Hx35xPDhIVAZochmVlHpWlNFNTgCtbq1e5yRPAnxWklywbYC0iSqHt5nJI
jG78j/bWjRiingfnEYUuEQm9qRCIRcQxeCxXixEbP+XoDCggqX+AHb651nfNmhiikfm2+N3wHYHh
vjbHd+83irGYRvWN2vI6aBBIY97posZL797KNwMUkQjEUctmHJ+d4Up51w3HYSXseYKZnEppxAsX
+Bs+rxmt3nYp8Sl4y4gD8XUbqa0t/Hkc+xXHK6D1oZwNwwyQdLuZEUpFh7nyXSz9Ilb9VowC+Z8t
nmiUu7ZQixK8tYxL72GCcUCB1Ez8wk9nYtO2KRMbm/t8RIvaEZO07Rr0T8s9IkfrrXc3fx0dOZaW
zjnmh3PUSVDchwzOCzX9sg2qzMrOIyWUfCY5fwuCS8M0ZO8zIi0+H6svAe+q2o5+4uHU9hyX0Pie
LkrFj4i1+2fJjunpctPVmX6nM/bfMsEPFeSmG2CUY9dpPIOirStSDOaAl9jx58IOFwdXCpDEHBcr
Eac6I/VrRkjQlAJipdxjDma8QHWwCYHIbvxGI7WzgFjO9hVcZpIIO070nqE9YdOQUqujnSBFtjWq
VtYPvaofW5RDrP1Vr1xjzu0a9HGc6wmaVtJYwx3myevjdgDZopfFdpT4OTc3kkA7bO+pEnkjdgdX
bMzJSxnluJzTfIvdPZm731ZL0mWi1ZGXbtqXmliAsQZiz1ij+L4ZFUVZQvitssRQLjb+pyBzrVuY
0fDCwQeq5cdpQCQHbKVRiIT0q0vE8eNaJSlL64z9cVeZmCL3gKqrzzRq7One7X3ZAWrZJlsAWaLw
tmUPiihAUSRCO1uwf/Nimbk2+cXVMmtHxNmxSvEOym4Or2oNEHGvfYLJQQiJjkobyC6ESphgJsQu
OzyaAb6BIEy1QrxqUCFbhcsxlUmG8BsxqoxCN4MD3gfBD0dDjcd85wREEIfgUEAjr7BFYbygT0iA
7iHpSevM6B8Epc2rt+hARxo9SqEaWMwQBE7VabgmT6zL6TVpUG5WKsx36aGft18I6/eZ2CVkqKKh
SNE25MjfwCXFs6h2D4k8+1eiXXods0BHpT8J/C5sG6ZvU0ggygBNJMzAHWuWSx/DEA9b00EmGvCc
liZS4Pj9QosAjAsMGhttQVkSeU0SJ64xL8TU+JuQSBPQQ9FLHI8Rl93xJ4KQYDw9NJSPq/lYppgm
003yu9p7erxuqnUzcciy9ao/Y5t8GeZpwGmnjFvIRJ1Tkf796CeX/ZzoT1SzR4WPA3pXQpwIteOI
7hlyhcG8xtBANOiCwx5QJY4MsAqa/V4HvyWC4j6qHz6dcCy05X4M6wUhfaFGuKOAHYTPnOr3KFzG
5/I53+bVMo5OtNbI+334Vq8jfAmnFfUB+9mVl5ARGIlzizGvN+jzm9JFYV49F503noRtv/V3Wch4
oRJPMaO8YLskyJsdRrwwdGrJPv+4DBt623g0fT+BbigdlwINM0I04kUMaMj3gbrG8X707/upZRZF
HFx/y9qXlrk6P03kEDDrhKx1dpOYfitYhpbsdbBcGiFvpe6UhRbTPKE2PGaOPmRU5sOQAxLkMHV4
B0BJWCSjAjt/cHgxUjgedrtybnZ6rBHkFVGZpVxn2pw/u/FAgjyXnUDGH6nVhUaC9C1m/hMzu1uT
aX2u9P/Pr1RAtsajes+awy42ik5vHn86Wkt+Gq+9bh6yEbdhXLNraerTieUvpgZXFqH0UD6F3Z6v
+siXbfFKw/v13gT37UXKokZWXWO9gEp5Bacztfnq1c34g3Bwty9xXbC9KBA5Db9TUzX0Z251ch4T
zoJK0xC1KAgBYDlbB4UyAkK9p3GwQfEAKkj0mfyOp8hzV8SiiM0RlN5wn8f3AtyEwDJ1P7L+Q/0y
Rap8ZE7WJUMAcRa2vxOceM/q3prdajg/MJDUypl9uZYO4T+LKxdFYtjLlbE9ILnUHttkfzxFnvei
pQ2HzDEWfSxoFX1xONv8715tI4QtGrIcidfjRbcwX+vHkIa78j+M4PP44Yg0q9pilBAMurO11ddk
kGedEpI1CxKiJrZ3EzToHGb5m6+mRhFu3wgmO143dO3bPBQU6RwXG4jnrA7WNT0fLmEhC8H4qwMu
1fn/2cd6RMqeriQm+duOeTaja14EZapcgzDKqJT7Bm0xK2/6SUbJyJ+SXDo/P/zQhlegP6zhdHr0
uvjL4p+c8+80lJjCX+WV1F1Tvl2laF/cK6Et0ugfLqxWguLubBGYrxZwUvvmhDe5Whfd9xhsFsKz
Qip3kq5NZk5rTmkLe0aD6fMv4A7aEUVOfiLJlYOSyHKND7d542SvO6hbUBmUfwi5ovz4CZOWczvd
un9CidZd58QSeDYT5OcxfyKC19V3wiaeAY0anDcLFk4EBXrZybMKkUkYrQVBskdKjbroBsdSXA38
+Vbdl5VUel4IBqhLHCzPcApyh8+gEU+QEclLtzc/vUx0s2bHmFLePe7ILkdzx0aMkczoDXyyzof+
p079nPU+t7CKspQRdPLHaHTccI7DlHyxiTXxFkHdf3W66n3K5dKENGXXyNYoo383yG3U2+aPJuP9
vzJID1MWp1ItJ8jBXqyaQoNJ+DviPWSi3cb9hLOBP5SYTPB5b4w9+jySwvBcO9UqXQej8xIFmneF
YHYQjotv9kUKIcuchjYJDlkS+WOfFD2goF0vuXWdQ1zzAtfQEXqaSSJ/PjD3wtBb816hpbjynz3w
HmNSOJayyFzY1CszPK1sbb5WpoPIXZiTPPvmIHgzUkCkfT+JL5bwzxCmla66HuFONAQEhTJgkPDr
wlN++36SkGjM/W4IZzIVs097bcwxEZsbgJ3F1z3Sm04mOIdxw/cpbXa83S0pSD5jly9LAkyUVY5e
+Lns+mlHz65eDw9/pgRUfitEFUKLf8iZo6sTE9JtN6GX1/qtq8SMSSohRAI6NleVYOozVfP8jRio
zWhmJZY8D89w7aUu54dOWKcf2sVlIW5IJsMWMeBaHFMGAPuCh8sn92S28SZkmSfmpdqh6LDH3Wmq
AKxmGiUQ3qnjiqu/uR8qSaNyhb2yrMneaisTpasojNdW4XWoyo+YmgfmM9A+D76Q8cjEqNwWdcZC
kzdsMP2G+HGi9R8p+QBcN3uAJKRC3d3aSun1ghBWjOLJN1VU6/347F3IdEw/Sof3L+oZgvL3UqoS
ispxTotjS+IIWPYynKM3qOVk9gF6nUyRnaka8yxvBDq8Cdvz9Fd4xwlmIAzua9MwVV6D4sbOzwVs
q/ar7uPMH1Vc5mqFDLybuKW6KscSL8WX6adtx0AFkeqvLNhS/xlY8n/l03+4CiHo8FC3ErTIcbLk
7RHnuDtGIe/NWZ9u30QcpFhO0DYrPSOBuvJKTveuiIu9ajWJZ6lsxUvJGb1cWePxCqPZFb9i106D
AeNc26uBsUjuOQqND/nzfGhR2gxCzWoJi6IglnejJq3lCSP7gVfdsGsKw+EfecoSNf9bK7+z055d
2EL28F7A1YMT9o8NFp2Tv2ZD8/TISjuyRFcCHpeeYsNx6RqTnq0pAm19LJ1UTxzYNkI3pAzNwRK9
dlkmOCYrzqSFk0UNt2/Uks9hFTlxg8xZpAyI0kZ77Wi+ug750Pw+kwoLSNia9OgzB9oVLESvH84X
5pnFpkhpWsG04+zdU1XDuHgzeoSn+Zia5eH6EhXhEJzR9zDHByecgoKb35IPPZCJ05UBbRe0RJ85
SGBlwEJ/O1RtQIGUIWEKzpk9y/sT60QuvlmBkZcdFw58kKfwgnqMAtKLRpdH8fgXMRZJs7y34m+S
Uqm+P+kVvVvCr7RvQZEf92S6VHBH+5H3KQmob5YQbU9HJlQCHHM169BJ1gEzP8tm6KmZFZkqPxwh
IxqS7/u+tdx95ndUBSXGEqNQQKiA6L2WjjU2AxX3FKM1Ay7ZvTlmlyHIXKb2STPOI/YzT9wqvRf6
JfKIt7GIG1rrD8QGjHyjcLBzmiS1iLW1Fn/Vm7y2BfEImTiqyMEa1b8/6/UpNBANcN1HLn72a0s0
BzE0Q3RHIWQfTMGw5fhHdZ9Zz3GnkhtEIxaeShiXF/lHuhUZbIS+DTdFSusHp1F87XBKrThD4y6L
CD8JA0kgBYridG6kp0FNjnSczmO7mtyvlXDlBHsoN85bvneboXuzN/8eAx7tu/OfcMAt9PIjZe0q
Cl6yjIHcT75M1WVJ+ErPPn5x5aSgWm6l/iV0OoNFTYvdfQVs2soZsizPX7FaTPAJAbpDssSe8h0o
DkeYbuAg6cvXwkM7T2lsVAjcAas4h2y0CUZXAIKIFXd2CPP2NVooyyzvhZoYeQzQs3QQF/pMJhPb
iVIakXHCvun9ZSN2EFcwfVvdfu6X4bAtn0l2oPbU/TiRreE8lXOmAjy+iIZkEPunisGtxKnz+65U
I8aNByGLdWlea7zWqcu0xZsDMhDfmVap9VrdNHqBwZmH7OfvKxQHHsbF2wJhbLwJu440C+criYi0
MK57Tt2DT959oOSacsslKC1+97CWZL+zKxcm1FarUw901142WqJDuMC66rE+ZkDmWsPE33GfAIBq
bAjRS7Bwh0M16T8UWDUe1mbhNrJ0WoNkruLXWiBNQnrJCD6+FHwwMSRe8FQ2BwISwAQ/M/xUSaVZ
kuwVXqOGsmYBmNkmvBgbJSJwM6ch9JBxkqBwbnUjWBcQm1pBlp+Ee6iJhEObxDm3dD7g+/QWgn12
xVFaQnb4WMTt1589uo96+BVNNYpAk/acHX4t5oDgA0VUZv5P7kNDQ4skCUsA0PT4RaOho3pFJZ+r
T9FL3qZgjEDGS1Sn41hsglCwSc+S2ki+ULf8r2IRuGD8pM4RCElxzYPcSzwTtSPDJVjccSJLE2zw
GyHShAn5PSY4dMNvAOdnHJEAeUbDN5HA3uwKbvuuCKAF5ndrkGuDAVI3bQ7TbCQqmIVbpqPbw/BN
NGOt2dlde0ryy45/oRpSvebXyquTeuZhJXY2icUEIiqD5nJWvy/ZVlB8N1U61ZjrvCYDD5s+vHbt
odLKNrN1DWMmv3hVOAW+Br8eFnsA7EbJFeILXZwQ7JmpDrBJoER6W89JAm+ZyzBys0uJiKWK5dnf
be4+lpsDqNxarq+3cHbDUVwNJ4cjv8GH3/5sLtFMSCXagg8LJ+UWpXhUgD9++IglI8eUavtQkPfK
zUeeSkyMLUeKISYVbYBlAInhiowO+PhBb3455a2BqPieuQIMyUrPCGmmHoMZH+ObwqpxeleQS4Pl
Ud7mf3BSItPJ7Gosfw2qVaCy8CuJNRVXryLQuQxJUN7QlaROOhkXi0XdbGx32ggL62kBQ0P+8Dft
8qfDqsZOi+sokrHdzNRX4lfram+h+kVp5pxbnmPxtm8tIgLjaavRRdhU/BkFLriu6BP9QeI7xPZN
OY8AyyzH7GKAiKnQMy6kQPt8IFdhSsA38wrc00mS/fs8AlAYxD9maWp5lo0U0u8uewlyXW/XJ/m7
0SE3ubKsqVlLT94iMCW5gDLyhbqs31odKQsHmv8FJgV9uTu7beKTyVCJRyE5dk9sWdaBODyzrILd
ZCHpuFQMPQiCG4boC+WJgwAX6L7buIK7Gpc87qLYtpOaMXhWOVLt/V5zbdlH0ap4yqItBlLHfJsl
GP2ne5uhi5zqKUK5qWaoJycn9r9ZRIjfMDIjofnBI1xhOTKgTgDESanZYKJQGh123YZVjGc7tO/G
leUogoUzZrCQmb+um6431MXZL2+bhlltjNYI1/hkUZQ2hjqOdFb2kaPmuYA74w0vj5EtHcFMcZJL
rUQLkGHEOkepvVyFk8gzIWBpQ9v7OwwX0DeMbpvMinq3cxniBg/P6060v/t0ldG2qwx370Ujhsua
m86MWMI204lqCgFef0y3LDV6rWIT3liiCxV80xZlIy+8l5K2ehxV/eVcwB/8ftrfuLtD7OBnCrq1
b2KIDdrwhG0cxRghe7aNm5aTQCxknfOeF8rfkJKOzDHWk3OLrY9PQ9Ru7eJbSM1aqiNQ3s1bBgOs
A2QxCBp6HJMaLbZIeFFlWCu1XGxLuKIsAU/C26lft1lrHlIqUqfTInrYA3SHvS+mZxYRpoJR69rx
IEG534Ct2Raldk9RiPFQ9Q2g1fnsbJVMWSefLheArymU7dGdhzoLw1ZBaPGHcxAmM2lB63NHNpE1
ahH+/6+L+7O+7vtJswNSr20k5jQ88gcUReXqknzZDnb4wIUnCloq9NWbSw5PsO3meDhz0whX1v1+
gacEsYq14RRdtAUxgC21jFz3rMBFvLxFps4FfdvnDreggUlW90eGNprkXC9P2U1CpeqjueNVwmsm
UyvZrhvl7QAYsXSXl9rZtlEXKatxgrm133ADvVMbquy22N4NAsdyy0zMCDYaIIICglBXn3LrYYnu
T5/tbRTJ3qfygqN6lz3DYZIED0SXHqJ9AH+5u+ozmjNOeK9KORC7ozIXwjlZgzqTnDaFGCEuU8zW
OvezeXNMcPYeZFHaJghIWpSneync6fXljL9ZQA3d0ONFjlJymhw9uqDkoCPk6TaUCJa1GZK0a27U
W0E2VY6WHEfIVeOkl8e/aBAncpYj49dVq9VcOA8Cp/CzAWxMKltS4tfIgO6BhRPpbo3SZ+LaV6E8
FKtgduCNTskbm365EWKmeljq8uUc6tdNlK/2IybhhHxQ3sgyDld2p5/jugkWcLhun7VdTVpsGTkd
0jsIOdk47bZE88HTdEgnEaX0LoFVjhcVjpnLkws8/xSx5tQG0sdxYOdR9jfGQAgvjGcA7LMPHoBq
mgCertAQkVmOtZaOTalgocXbdLdp1evmdCf1ZRrjPv2CERzyxXUVlsO55W0EwF8JDqRD01vCtrUq
+P0mjGCTeqQ/Jqd0hrrqFclao4eyn/4BZ60+2QlAuxXKyhAbrcxBkEYUwji73c+bkKoXNLkd5V0D
VtGXUc9jz+1Oi6CtVKjYNseZH0zjqCBmpGLiyrCmsVTfdAjwPwF4u0wkQWKfWOAmNEtzPjvsZCvz
ng9JHcAb/KJmgjfRmd2KzhpNmCJx+6XqYKzAh6vxiLZajYikB6Of2hFDWOJ8guIKOQ2S+bVmI8w4
TI8dc/ahJbwUca7UiQ3y5FUjTUuzJ8ir9ijsxQ1cum+031A+kCnBgTx/sXr9JvpWsg0qsWvd+3Oa
OJvZmTNgpHlV4lEeH+G9b1CQc6jjWwkBdf3kxg2Swb6l2WQlW9GuCfvHRhVDdzS478kR0ebQeF41
+VC30gsAPJdGKG9SvMXtJmQFKaizIfD4zXl1QXN+O6QKubnamltt8zUMuC/ma7nlIPQyzs1xtXzu
v5BT2ufZTIFthCcbRWzJ4kvIiGPEOOQSBFbGXbp/x9gMHtLIrwFq2s00D8lWV/KsP408xpV8TldJ
Yh50VVLo+xZ4jnjQtYSMYqiG6JCikASrWKMWPRLee48zNL+l+JYsRqU59aSnkQniawBwEaYq2+VQ
yqJAUBH37k1KdOqTKVaCdnnmwsQF5C1q5qtJi3L1UtgYk6jwOgmfpuUzaNePU3Uwsc3NgRctX0/1
gart0pOwUYWY0b4qWF5s1mAZX9MpXYdaUgxct5QY5sn68HceD9cMrGmjRkdic7rdxRqwznNvQWX/
h09UGM4uHDp9kTCZX0xPGeB+sneUz5nsldLVtjBV0ztMqsalJuCx2kobPnp2y5oTRKSaslyiS+1r
k0u/p6Acuk4RDgDKbvhsr6OrkxMoXa0xHRxOmEJEeLLRQcfynOnBq/qVD71p6I26mcTEhHnxtlk/
EIoLUBsCTWRhdlCMsVkjCnPm1XLlq6gC2cT5+0+cvwYqATCKFsoqzPMxo8DQWNZXyaOjp/lzYJZZ
/0KVwSO/K7QK///SiiyBfq9Juc08WmtrDyfdzu5wam3MhRYN9yHp9ywYYNr1qbZlZTB4Wjjlnn4k
PzVMOtUYGWYGeFDin0xIxoJbvP3kNTBfaUPqkGbZb80zZD9CMclzDDrCKsJ/IBTaNh2Avp8XdQFa
8kn0fHGbNZ8olyPU58JIZp4APcH4g4wpGbd3nXA+U8LgB69hzHruSXnUdufrEh89Fmwby+eNbB/7
sn+LLBxFujv7WAbccmU9PLkGjZYB9A31TkM6L9c0ofAgnks9d8P1vfq2qsPAbCxHl4r2Q25arV53
qMqkMQAsHjXqOgbir5M+iVInoT96Bq4He3Zw0Xif6rkfDI1gCLjnlgygRBmKkGGWHycnjyk6YQJf
r+sENZ4XE/zgU/WqtMsuX2od+FSollHRqPw8tCZr7PUH9le0Z+a40aJHn7DcruoxRYP26BW7NEKv
VdD4s5BJKnnBYfApBQ2BWDtgzI4S7dmwT9Z7fT+KS4jyBOWBBY/+QGENz2F+8d7CR/yb8Qn8mIbI
3vqnVfs4coygAdZxlImUMhrQKN6nrCB000R8OQMO13F1//dU1umzrbyRWaarXDxmTe3LcWBZEDFn
nhN//oU14s0cpRPZwDghm1PmScCaY7fFlO9JclS/nu/lN6z5Uflg5l1NOb9Qddke3w5rgOUXclzl
bdK4UUBjVjUEimTUmlEvZ63MlKyAs2zQhkxOIbj9fTvGrYFMwpP0Iuk+1o1ARKBEFWwHZd4FytJ/
vT95luS5hl+FaS6Pim3fooUlXA8O8xq2ZFycyuQHM7iEe72AIW+bpskziAbXplyHXsZx1Y6M1Syb
8Yh3d1m50ys7H35g5imtTh4fiPGMNI0FRy8FFrh75RYAas02oCh2z+bEFbwX5gxQtxb9EC6ba7Xb
KSVfYnSEudd1jp3h+BPa0HhdRnfFTRqCaOjAw++dVTLDsCzHzVyF/tvrCD/7BQdgqG9l+ZGO2wsT
QSRVf4wKm5AtvUurcS9PAmjmp4VGKEEVvCy8uVma1F5wUUNVDAI/+Bk5yVaCiQfsV3PDMJQFCkle
tB7dosm+xh1qL9Ip1kgYLe4Uc2phq0xQ1ep53VYdBqdfT5XppMGs/jyNKMXNvDi4R3LTV7EU0VBk
k0xGX4hqxw4mKfDYKLvEDFR1/lAdaUaVrQp7UIsZ5fa0kwmpZ7M1gKHOcVnVCoG/J6TUuOueJDKb
soFgzloVYAyIVy2QjqmGJ5ZRUe3z635rg5dy+4ZMmPx2x6ZYqfRA+mG3pu2IrQDVCeKFbdqJb+nc
3FFr7TAEKoO6Jlu51qIkqTWjjRSCoD/61pm09U/oAgdpa19k617yoXXyE975TcyF9t/qtJRIsKxE
Tyup0+p7fnyU7L+PN3Fg9LR6/9R9UMy2dhj3rdBbhZPt/PDV8qtT7FH3QZJhu2SwrI7VluXDRDnL
LfZQ/MJn3UVr3GUzt72j5Yz35uH2bVt4Un9d1fiUz4Yzs8DwZd8kom934HfX0+WcuFgx6FoybVjh
5XXxwPEskh6mzii9BXeSBORfgHXHFZHIq66Ufb47r8OPWx4feiCjiChgF/7f/2Z90qohJaIee7hW
SJZ3yyB8CBjXZl99lyfC7hzOuodaiftDKsv7H7zLCFtdnEnRnJQIe4jBmGywkzkdxBScG14Clazd
dimE8Ujq/YTpPhmKiyJt4N2f0I7aMna/2Z6pTm0xNOvXW7aPLffgOkJ4srPzEOrbaggcNdd68/h+
Mjmn7do8b692+cqa86QBJLwQIe4JRUSZ5VOvPGr0tnitjYIB+XgM3OuVY535T+Fml0HYC02d7TJn
CHCb9b5M608Y4lDllqJLZhcT3WYr8U2ueZXTM7R6MP/VgpkrMvmB9Q3aIOrEy+N85mlgq3TgD7TF
xTewCPxb2lgtAM8r92CrD1X30BmRQzMB/DQt2AWB0HxB7x+eJXe+8mUPQer2NvCcqgDIuzqtX+ci
6QNrYk3OBksDSC2MndEuuQJ66mQByeBsD4s0WPQcDJJ8g13vCzCLXlU/xp/9w28T7FRNYKKV7373
Uu8CpbnTjuikSCe5EYZ8+zFn5JP0SJ6mnjneqtW5DpKpcLC0UKtdkLRhx+13ehZo9mFnPaHORXu+
Y0oR1pAtikeOsVJdmzRO2nCb+m/mFCEvgz/1MWYH2ytyZ8+CjOzAbyOVG8OJb0FAsx54BLRrMhK2
xyvlR5VXENjjd6imMQvs4dmQc9n9mWr3Vdr9N0YX2GUdn5R2edprl5AE0ff1Drqp64CnEYlNCEiq
k+OUDdJc46xM2FYlLUFd7PgAkC7qX97DeaAT15/idAJxFkMu/wyPJDsWkcecsZEB3baS4liEBtw2
u7EOy70xpAp1OfG1DW3OUlbfZTsdIPrgpv91JHPbOx9cFRrAuJx2bYowBMj6iGePUGs5KSTxC5Rh
1wwu47buZPdVYpChBCZVjviag0dYpCQBc5JH8bNOxGWUccrrwFAi5QO9bqP7p6elkNe0kO9q50ZM
CPubE6N56HPEZcqJC5/D5/EU++ZWBFdJatKTy0eGJjPD8z4BygJ1z20iSlNVoK6wKdkOkdSis3Zo
TFoC/fejQRQNqkyxf4p9sz7XrhecUDgsvd+U2jBpik8BnCegqUH/k3Wv9IqL2F5UXGoOVKWC70ON
TPyNsRrlDMpiD1VOH9jxQPu7JtqPiAE01KLcV/nwi/VbnKuK8nJN31fgtcUrietSjxT9DTpdgfZu
WSHrt/1jV9qYXFfWuTZUetCrnNfBwskV58sSufOxAGTXTrvIHktVU4W91J2l/8B3A52aPzDlC8GK
YbHpPPdAJWkrmxiq40elCEvjE2crsB/8+LBSEl62J7iaZyA+SXUtyAwNRTbDNzDUb0Qc4kqDu1tE
SWLCNmVVXcAvT4ssRAyJ/u0iUWt3qLb0cPQPu+RqIgiMj2byf0zdv+vqo0AQLq9Aa4kleus7ord2
uE1iuplljYLx8h1z97jIa4ZRjs/3gQ/j5FIPKu4CH6D4me3zIIx0Gkh6ufgpjnmsA08mHz0ARNpV
poLtzNH3YTXnaAmnb+lAOGWWkyDoGB0HiT7vVdlP/JiCG3Utib4f3g/o7NJe0wxZPQYYSmqdgkrs
XZPwJJC1FKWsA4xnIcCFeYDedlCe3welA4S9dbUMtKyYPKTEzV0vlRzckPl63siqjqIC1U3Luwet
dnVLUdf91wA4cUws71G43Rlvru2IednCkKfd6BGXfny5e4NzHUiG9kHgVMm+qDos3dOLJrHrhEK0
wIwatKnhrajshDWonxtDmBLItfND4d6/OWah5rPxASXvqr+iwFlUzn0ATGXldzJ1BjA4FBOaOol6
guFLtsNXcXg8MFhPfgcvpMofYKGPdNrWxxMrKX+m8PGXbzHuPn0ZOThiCZGwP/5UAj9VpbxGy2Rw
nlNQOMH50DfVMJZq4xC+os8HbpBRcVY/vynB88Oj11rNTbe5NgPHyAU3RnsKrESUyDoTE3BBJQ6u
53iiH5JmoB5Z5neFhjVcAdWaHby+DwYdYMt8n0Uh4jxrX5qoDS9TX7ZpA7VO800Vm+POxeF1wEV6
z64uWuzfnzFqJ8ALUXIM1TFTgbG7cjmLDhKiWeT2pXPGy7gHTCzksHegvDBcRuc677EzqKxUV2g5
+7ML55le3ld+uIU3ovlbzF8GNGddBqWt0WcjKhD4Kw84iq3NdMB0Q6YzuSR8m4PD0tnV1h+NeLGe
+vRNFZLDSfFtr/2qGyYQdoUdcBU1Oc4tU2mM6XhNENCuR/aEKkusy6xmEF0aRc/OCKQa31Em1h/z
tLFRK4m+4lxaHiR1RYfcxyD4CUGftN/IE0krSojljK4IBKJKTIXeVBtSYXj0CWVNu/7ccHPeie92
21fhF6Abk2Bq9Owoh/Z4W4HsmDMGpzP9kWuSoyUAtdI0/aVJKgdaw+f3lgJQzKXbnMSECMCThIio
lfc6aVRCHjdUnrE2tgSNoHl53BGWeXYJkWtDTRTIoA7xIv6KoCbKLp25tAd3dW7wWlWkd/O4NKa0
9aNk0Q3Bk7yBlj+7ogGVmoLE+fVTFHwMjQ4j3EZerObpiW2ALXhCsbw1rxZZUuWNk6rnfHAUeciT
ug+vmkWEak8tIY8nbVSsZTeapcnsruBvBkxwUDghvxMnpDPbP8jpL9TEumnpb4b16bojktusR+f5
a128WeS6mlh3hOK8IrTqGRmy1NUBKJfm9KXHbPDne8ujYoX+DodauVLw7ViRwaUkNRVTW2DznLu5
3BILpCEtpYaqZ62j19UFNhKAlg48ZxUFt42zKNAZJi/VB8lmWAszwr55FubAL/PxFCTUlFyGrX0k
ei7nOawVst+bM9F+YZvZDXZVF883XxlO2eObWvm34c5juBO1fXStpno0ZM7HogepiYve9RWtpdQa
2OsBXkWbogtBikbrJW8pfc01omP04jgeuHFA/bui1pkaw6ZNx83CWoAuS0xC1pjLyAjUi8kr0LP4
wk9Ig6Wvwkp3OdLIp/cANZMPd1rEQTwUKSCTXOVHcKWE7Myz9DhLMrDM3SIV1SixPOCdKtSkQeO7
DrugYa3gPGZr69mLTkaZBB7HvPsEgP+hW8wAYsuPJXvVRs7n9JxApGD8QxuATbPSgwgfWr38IKFM
MKgV1YmoT6zhPGSeXLTKsfjbIW91dEkIQ1b4VeRVIb00hCnmZjGO7UyhZFcmYd3Fht3IhKkzs5au
FxS1JQtO9OzMqBh1UhZh1bAUgRYNC7uPaM5uxkX/IQXdr5XwUJYc8WxYFKg/JpQ9Jk6olONPnP7X
4cqSWoVhUNNjBCJAITPG/sV0BvWf8wAf3F+A6lC2WzS+gHs2TqQjfajCFsSs5ReITxww904W//e0
dvBr6xrInL6Dwt+ZC3f6ZGelWaxnwdP9fVlOiVKSZxZKQSDpCjyzHktpuxaK8lmY1mEgUzLAdsOx
5iUiCqQhxHgU0iru+kCQQy63Wv2XB2N6GyEjXIZzp0OyHH44sSKgZJlLe5WKnLrgtpiWlf5yOcMr
NXnouymrXt/y3ZvRy9EBrTe2bQ6xQ02jdD+MyN/B23koKFf346eLD7PQbpsP4cYHHKwB+4TmgFZu
wA2EQY9LfV9JmnGiANmo3wL0eHT1Nc9hO6/Azg7cNIQR6mC9oxgRZP+pDHUvKGsx6ij4fCc8oHPs
LyDXwucglqOfIByQleeNFbB2HExK8gMCGxzRZIfCfQm3Le4ANL+NqvimVKAMjgEAOEC+SYkqerh3
2yuFG9XQ8PgDj3Bthug/WopfaMsTk7pX6rCLKtPdHKALkC0Le6fltU1kGA2mXkvSvQ+dljKXXk+l
uG1vUsy860ChHYtuvP/kg4j7Kydwe4+btx5eipawn9SN6ofAMXJ/dM2X2HKZGpxwPII+c6S4Ogwy
us6G6TqkgBDPOeMrBNOfNNCZ9iOBGWFLaHtX1KXc6zJOiOwdJ6dFb3QR711BO4BA0o/VQvI1xei6
pajdiZQlbBbNQWpaL6nqbm92ilMAB54BECAMSMY7sSHzKRcCKCdjbRzY4eMvs2bhUcMCRzmpShz7
F4p/WgZV2Hly3cUmXia5lyGRhSrjjSdnl/N92+vzyVqafTOp+k+LwgsrBtL8G05DSV7Y9wd5chFJ
3M05f4MR4hc3L7n8tBWuGWZxddMF4lxiUE/uqvKhH6X99lSc0Ce4Y1+v8vAKyfptM3I+ral5TqKq
hMPm9tXOsf01eTXCC5xbf5ic/+rUUvWEIx9z/i58mSBhMpaitRaWkYJyaSP9r/M987mYb5Qka0Ez
+FpsYLL2JLn3dTVn6wi5OiiG3sg8AHTaWgyz3e4/Ee2FwYRTwZHYVp6GJllSQxEkq0b3Owg3QdBY
glpRtxJDxCySdqe80Y6Y0bEZDfZiUoRnGoz6cG7L9LOF8qHiv9Ib0krblLyjkki8dC8bqZHIe5ck
TdPMvbysd0xME40zdqB+7utBf1IqsOeb0jt+WHlie696v/r3T46yPEnxF57LmWRxzWUqZob1FwFz
wlSZFtOIGLAkFmMiMIN1eq+hu14Lx920LXVRiYZio66EvoL3VVIZsBiRebjtVMxlO471jm83sFcA
B6Mo9qXVTy6jyMUA2+i1X3sCkR4TDJ40HBbhoP7HaqpLEHApO1VYdhlntFX1Q+i2esRqJ5L5g8nr
FnSA9j7iv4rRLh04inKnOTLwX3+pAk1M4yXc7m6siveA6qygddiSEPtRhoKMyAzzuYF9SFDOxR8a
ddFfZylMz5GItOfVaWM1JK3xoSJpOQRR5y2pV/L6VKWebyknPszjVg2YCh5/CRNeagEcxJ8O9jBr
nfZh/v4vXyMmp2JYehlzTdUY5VP38Umq5H0uOe3a/hsezG+KiSotsRKdi9Cr39Ae00iD95tEdLWM
skvKJJZ+jIqDJCgDk55I8TjbXpWGxPm+I6vANP9wbD4AV3zypcgn0QZJjoBghPFU8DlhLr+elO9Q
mbjoVJy7qlSqZOVmLyTHb/OjDr01UK0Je593Dns8Jy2L5PQvquS6AMcvcrYPT2KF1iEu3XkFpQtG
HbuF85VarX0ZW/cnnvqSw7ZU5XZB5mdwFv54F6heaSOiLN7GiPMM4Ag96C8N9wOdU1NYG9JuHlur
dxRXtP/hLWqRcFWLxwgjqVRcuObgMzTzJSt4W7Fo1scGAoP2btfuWbbUAoz2AW15jU5ikvp8aijf
fKGFkeGeZBieGNacPz8mfkoOAa3YkXMFb+qiS3OBT34zfvTKEkH5jYdZyDd7YZ1NTHg7jvZV/RR4
ibtWtoOvMFoCSz+XoXzI6IV7ALGnDH66BwaAeVAIc+JTDx3RTLYljoqPvlsmtiIccFrqF8fEuc35
AzkF4gIzm08QfYVURyDtde7sf2ffpsRuUJFgnOQD+FfWcgCdLOFR1+2SBqtfQlJJRduXciWcj3bQ
X48Oam1bt3CkFgKSB+nESDAG+lzqavLpqw9XLG4GyfHjAtXUoanbd6e1Fwc+Bm7RPpxB4vsVmeCt
PGIhIHl8hRagnnT6VqvgTMJASwZPPwGq/aHeHkI+v5NERcwVnRgOgz0/rjXUcdRw8F/qwpf8PAgY
VzWEbwhuP5VNzND/2VZmyFOx1ipOYf9Zyr0t/PcNlKOHq9lobFaxyCIWT5dNycsviLieoW0Q4mJL
jdy7SIX2Iw9WT6YqTrzkN4MtnpGmuozJZF7ta2XGQC68/0JWnTuKNyp+VNa2w+MDuKbrCo6OfsfX
05JBlilFEDy4L0U1WiiSQiURpVj9Tu4vVjFNZDWcMcaxnbi8sq/B+MaOy3m+2Xx9lUDHZuyIQ7EG
J+F7DCCkJO7KlUdXJaEg2Yq9tDMkY8ahNx/vr/7/xbJHyTBrPDIPPiDPI9kr4vMqD3zRGMb6OddG
1/2nJpQDhvPqPUfHtmNkEgOth+ag+t665tisM1aaCySeqiR4En1k2xTfZO/LyLSEq0dhXMMLImm+
RT9AckFHwie36MC+utybD9E1nOtKG9t1iZ+Iolo5DLtPrn7dSmNvCuw1qgNM2cUaQOchBiJjEV99
w4QqI6bXHNFI1I5ZZCyF/FiwlDHPVTkynpk7sonMy9PaTKJlVL1Qwl2ouGytS6GZG0QPqfw0AKq+
HMiXNnfwb2X7mrCVt8NrYK6DSZR15ZHuzvowW5H7Q+U14FozndGEWqmQj4Hv1JCc+wnAf74In4e8
oG2JwvC28kAutHfHs/NbRyLrXuKiEGVXynyW1bFo/YeMg7hKxx696Mf8R5ZykXDVDI+mSM5y2QC4
y1NIlcprl+KpejDDEL4B9tBT2INutNhBQksJFti6EGP3wkgB+aZMQ7fmSaO/1UegpS4ltQbhTWRp
sSb7GhfaYJPsJ+4XeC2ZMmwTYN/XaPF1S7dBINkUgEtqwYZWFMqKDQmxnKfW4M/0yiuX5r7ZuC1j
/bJry80qK884W2ez4NhfQKUvuAQDWZAd6F11hUgDibROlqZ68PhlLanBj+EIYA0FUk1qbTNnguqS
1Lut2XYynidNRA00pLWQYhsDArRjx8QYtmZ8jDLehfN55qgZja7AD6Ioj1i5WDLu2siCl5ervkfR
4vCx2t02VtlJfJzsAof904byfQwW+dEwMk1EWgyxFwPaYT46x3bNdsymZjMeuc5cYJkyYnvgNXbI
JHvsjkGW3qpnOv7kUG9AfYf626ISl0vleX2GSfXm89grm6BBuNZPt+rzDZmu+reqU0tjiAnd9+Nh
8fOlI8sjL8ROaiYHmQNMeyImhlIoaa8199snLmcefbhv4nGBJclDRuWG9OgefK00h1juCJmAJ7rJ
IgFuxw1+dZkyE6XyD2NlWWlFlZD8n7K2sJlt++YyQI/pg2+i3zrCVb4J2mtiPpUDHb0F29K9ocrL
Px9uVVu1bgXdOf5j8PHtYGr7unIwz+SLHw9nC6NY+xZyOAN2DWOqyo3o9T9Vg/iBgqYIBS32H7ym
oYAtOuFoAXKp9WKAl8MWhoyPGhYkE1z1E5a+ZcqT8bGdoXPE3gnIhoJ8uf3gdbUq+G9XLO1cqpPl
vJk2v54cWwmFO1E1WfmPKaT0P5eKTS8gQ3qtJiFHrTn1AQs6/USzLIDo9gRC0GjOstLyI/esSoai
C29m9NXA6LKnsT5RTDWzVDKBmjfg8Zn0Cweh1iqinUFDcYZUsT7w3ZnqVdlGORicprJSvXRcTrxr
QhTOXNQvj1EM2QAZ9CXr/phc7EJngk6AcVvChs085wvvaqPzSrOeOfNDMyHG8skkudKU7DlWYUzx
YCxlHQm2SEXkoXyD3S+isUwqn94aeCpqVdRlWIeYUaVzwYtRqr08M73EhUjFechgTa7tJStYGxZ5
rXWFpOALdBl/BsRdTVfbvwWf6/77KWGVb271uAXISdCMXRofN6XVjyQQxfWht9bqpORfijBaQ9a5
sS+P1l1qBOaFYxdkIvXRn0L7ydFju/5rGwSGTILJ2bJvYIamy/QEtVYjtOREjfdR85EvfNk7bPLT
/hzfY6PzXIEf1PPIugcL8Kren4mRTM4Bg3/uN0hEwjtIl4LdmkgXH6dvoh82g90tNpndVD6R6h56
jOJd+lho7QDTQzKk7VkwHJBvq9qgzUaltxAlhNOpWbnk1CI4Zv74szrk7r2zEwWN1QDxR9/q536O
FVORJqsJBgofMu6Uz3OowM5bE2ZROLA9yPxgbvPoi6n3IQX+ANvtk9yOkC0ETAQJmmh+xOsxmFlW
oWe3M4ohjWOXGaAGPR8/DJWtmCbZxLF5mQI0VO/MNcfmK+41dExExOwGb2Xl/ItrZ6AP2AHlinqw
ghmoJbyHDQFpTCAU3xAEPgjmDkmZ07VGk+BGGXkKE7ONlSsFDsu8b5g/5cvpZoQA0RPX5kFPAyHP
9bOXn8GCoYCmJ9O0XXlsjvH5usDeQXp8RGYRK1s2n8tCS+Sq7v/+KK+r4AX2lknVW1B+TOoh6c90
UJIbk1H8Za9ytA95TMAwnouPXxHi32sGY9b59NW+uQcTDFlJPsDg9werWnpG2xzUHRheymK6yeet
4vI6ZRdlU1hY2ipQ+/olZlHrKgu3eYoC5ZHJbiyQ0PYI0FxDEcVXgGfVhd+hOI7jcHxtpyWT4z4b
/aHon6VVby9S8yfLOnrvjRVAnqu0PNHYAak4bj/1nKfTYqCBTAi155Jrut9hQeqz+fUuLm7EuTBT
OTOGTQuFh89izIRS5BadBiJzE58nL+L/tNyQmFIrpDKg3wDiJaF0zrk//82Odf4E2AIycF/c9bPN
QuFxsdPyJ+McqyD/TyJ6PN3h35u9QrG2AsK6ZdKwTH4DAUMIefj1lZRPYzM89WS6UtWmVGdGrok8
ukpTZfecwzaeFdXtGKcdT1UctnE701HmwH6+RbEXOlzpGGiwwkArrqczc09QorADo6yRnyF3PllN
haslqsv8GNCcaxzSsQo3wp9tUjNmL5adyPZ+DKEGdQj4R9Yx7cL9LI71cERNk6hDUDFBHHrBCQn5
mkQsugQNFSl/tSvmexj6dn1VbpMB25Y+T/NMXzPIHIdv9QeaB0F9/E0cLyIJzaz5zL2c9urR5RSR
bBclgS0GeOASm6OnsDXf8isb/Z6MdFrc9ZrFgJAEcAaM3jZaB83J9cLxFcVnAP0JI1tBhISLg5p9
qrjijBnR9C139343BxBb+TNFmmsfy6nIefTETrUAlk48ChTjgynuxTbdEQfkLsepz1loC5u35VK+
RkHgnWrTY//a9/vgxvmPTYwFyWPDC8RjlP38Yx+QPlKijqSrNBxCyW9hd9Zp57i6LUqhyPWG78yd
XzGuTOeL79sa8xjsX4aM7xU6D5EWn4u9SZLNfnqFbVSWsWFidF0XVlSOt9Dc5/Q+zIUF0z4vE1GK
fvsPxgIypiM/SS5dBVOg2Rq4UXVAmcBfroBYY7xCY4KCVL1nRiC+CO/1lIDAEwe30GC0O8qqJsYf
UVyxEszehgLbP7cu9833LHsyRRwIkd/p6z9i2DyqUrYCLx5H8vW1xlSkvdglE94WLBx6MBkqArah
QilprXjs7md+6BKAhruICpkI+EbCqvTxflHHRnEVjT1mmb8a1Q28Rh0gWPfvSAmNI31scmzUNhCo
DSyZ7iTGprYixMp+JrmTAVeqLUD9tnqup2Yz2xe+NxUVpIiXAkuwsv21rvd1Ug0DqB1NkrXMYclz
9DOHvPpM9IOGO3WRIvWJ2rxR1ZFg4Kw+Aq9623488dtItV7q5QqpnXIjqZo6nKUrU/KPH/PSueEN
oy5551cIldWlWdjhziF/mHGezpdLkbuEUdH3ML6lCGnOFBKU2emY5S5YC2ji9h9UjpEVAjcLAJ7g
ZtnDwuHLLEbDajPMiJsZ4Ze/AjccMzUa0bDmwSTgsOdd0oTGXKCf2xlnIcdf1K2ND7e9HCAkQZRY
IuAzvsPo9dtVsW0NIm3/fkS2J9TRE7ONsVnW6RzXNVUmJ4kvYIZktfElU5/l+TIehfskwNFOqEDD
I/B4oSug1+yiYRnEQRhJJOQuW1ns4NmBztK7oc9RKyE1iyhDqRhWrxVt2peFEcz1EALpkhzZtmd5
weux4GlWTIqh2aVxzfSc4Lzvr1QMwZqgAoNyeR4Us5g1ypWaMHx6MI1o0/KrBX2wc+sfGvKL/PeF
6dvI17YYl+Bqbjk2dLW+0dw2CSXfq/egWgQqDbNbzrqjKi94+B+pJvVrKEwAdxApJuJj6hx349wY
FJiaM82FCzcPbAABNbke1QbZrMiGOQNWhVPX0SaStVUcJ1a/vsWuO+efsGZGbD7YaFZLNKgHn4L5
QeQARGQXoUG4r+PjW5klzath2cCxd86fuGHJpPe9vDJhOjuvJ0EPCaBEsC2mWcmOyfCWpVITIpIT
AbMdVgxGOX6+3HRafIwZ9Ff91CvkdMdvgG4ccl03O+GzOkNtOJZKW5NvZCFnvQzE3W6rBkC8qWE/
YkhKEzQScS3u7BcowOQbX4KCa5+ZzMPibAatWfByQKKqqPaw427iFOmDRA5AhukFveOPAveIds6x
cg0GaHknuKNO+eZBoxZQYByCynkTD/PDHYQvwoJo+x73AlPIrOaTyz0dO1Jt18E6/o2MXDKtWcea
MoOGPX5alRRDC/NdzUxt+h9/rSBN33YyhP8nacAN5IBsLusNlqmw/NSHou1PTQQb539YnQBECwxp
QcpyHKfVM85eqzvIKdRDtyiw7PKx4rlg1McqYqLGfIHgwYjl6VhgTyDwKFrYZKqf6p5MiHh0E4h5
btpeoVIyNmfId13H0IA5g4KUrtS0Jx0zCIoU3KY+t5v9JeadgYYgvlQD7LZyvLSCsp4HqL4dT6UJ
JYLf+qXBss6Ed0/uO1fffSNzDSNHyIJ5q6+S7SGkn07QoxVXboDzFYcfpUXxDM7BnkHPEJKhIfPe
yba6jwRt8tVy1CDxFqkIDy0L0e8xPIOWvaJeOtHRzcBwHba7iWSfSFVtz6AmPaP1jFbb/rZgzVIc
lmmk/5a+WpKRX3bdfblhEVc2YKntQbPASlk66xewfsy12yBaXv+K4bm+CvthfwbjxJVJdcsjklJb
e3N/rOnAWY58ojAo1YaZn5xsS+m7BYOipAYwq7Rj8kXz46NUJaHSCn/ZpX6cUVEOOL4un2C1Phzm
aIXzEF+CFWqcK/fsPleQiwKXsEAaNuVuKoR3Fh/IvKXvfOvh8Y4le44LAlWngyrznP/nE77ChcJR
Mi+sX+kwzK5SiY0BuSM7vOV5bMPxEx1Lf4yP4ol4FP2nmtT6Pk0od0na/xaDbkzrrg+Qkx8jX6Mx
n/mIfshKjkFQuJm8oud1KksLObjq05f5QMFirwPtF1eokYqnZslTf9RdL8DvjuwofkSgBpWgCerl
bWHVNFOQKbVbaydr5dCiQhM1nspGbQvqK4epNalRSFExOIYfz/dBVBHDnb7mlwkc7Yooh00W4GSJ
S/cQrpXmPLjHqW3wOvK/GumvGBqciulAGp2GYNP6vhwLlDPC0ArXG52qh4T+hnUt8qUHAspkrKqu
MLzuUg6IRuE1gYBWAzbi6MnbKTuqUn724oK7O6uGnC9XEC+tGpJHwWXHzwlO8aCHrOapftjiZrxI
t+JPAL2XgxAytzdNLy9UYfoj3oY/RND7fSokyC4y8zjmokCtZJ+adZrkpmH5kCbqSbhjyy7Q5+Fg
i0iCFrapUuDgtdBCKsongU+pFc5aTA/J6q5u/FB4fBByOwxgRqq0JDSbGPqOm1yRqAyNj7BSRqRO
csdpHvlEeXdHFS8QNT5q3duS2NC1snOfGogpJ8W6jOko/DgvQIBrj05zjl7G+eAqmYH8YypILQ7n
Adc6EAidUKUfsTn1Vkh+YuAfCkHQE0OMK9xXQKI7IvJLk7oHZ87FhBDFOfZ+lYkV3eWgJZiuoZmU
qoCQZ2IZx+XodFJQy1FA/KUSPRCCb5GmiW7qP9UoV0quPgySZ5Z1r8UJZs/J6Pv1nln40Br+ZfDO
NfJhQLmvruTR7QeRLFpNcIsDUhbn/subETxwIt5okDpwJQ8a9HyEqiIQ6AiCRJ7rrMMevc5P0zhA
Fj8OBXbFSF6R2LVZWNZBn6LbiqsUymjR7M+0pi9TfgE1CKcIoGIdRhGqGOaeJevKjZqF3riy6eys
9yOD44pSRnuXH3eKPqZToZLlW8pKxW8Ymp+0Dbgrht9UOe7j1YPY5zte/+3oEfAMtMXuJJsqCV9Y
muSqmcE4k/KfHBEuANYXCUq7d4Mkfm2v4fOpU5AcexS4ldMXeRnkhcW5Pr8j3aCGGKtGBjQvsAIW
CD00XNIfWcrhz5goJYoFOP2pagEJMkEoFuJQDsmmP0cD1uGTSBPhpHygzj/sXa/seGECKdU7ZzaL
Mgq5rwl9ZnXXGTO3b2hnSgiHdDQvYB11uw3nzuvAyzmNjvaz9C6KsIsyXDJg6xxCs6Tw06LQW2lA
98SAuqCJu0PxV4tgs0BrPLQgDapCt1JuR1AMoICqhnbsETv6xfxykmDD067UYB+yGk5zYf9tOZXy
mePtGQwEpqvbDLH6xbcV4iETYt9vn+chovfWCfuafvOM/EwHjLD2/iQRmLB1B2nWDRYRf+nRyrKK
wHy3SdUQyxVoBXGvS6ZWHVWfwSBzv+2BkdoAPK7/K9Am14ZSx833g1CM0U0cGni3IBs0L6oclDGW
tEt2AdXFs01f8LPGBV7+wYavs1nRPkiR5LsSSpCE1oCiUHvxFjzsUyx54bfuzmJTLeUy3QII/VhH
Eilureb5fLfosYk1/Ca0WfY0mKt4OlHWLnyc3N56qMuyUky5jkXzW7tOJHioG6GoU4VTMNW3jRWf
khbtL6ofhM1p1G5sLanZqEQwlEabVj8fXbcZVJcNJVL54raSTKnEEDELgPDYCE4g2bgHNEMG14BA
SzE8gO/l+nJdX3j+sTuInqpF+Tp3gLUyhZkOUHQUEcHCCXpA6IFw2XbIHP9n8vuPER74+ls4ocKp
2nYjenGPP/kliFW6Qyi0l46irF0dLDWpK/h2EJic3nZAGcpaW2HFtlC2VCVYofv6b3ynHg5biEb9
hGKNwdo+E1s4rryJvH5Hk6mIgDRRNIcQ1jtJgaKH50MRz2wurwkWez00jgGYUUr/hj3tH7tce3em
gHk2p2qfVLgEAmHnObAmCd0AYtzGZxWqNx35S8Q6+aphZw+DP3AMfjWTBsiyb6jpBvOGfeRHmvr1
lXdwd1Fdxq2RYZYogfKkWlSB8HadQzXmn9stxfdE04a79/pyF+t6DQ6mEZp7jChdsGCW9E1OwEQl
r5rS87E3VL/iBoPEKeoYw46KSiX/sSJSGnE8YTmWaX6n0MIMi9vEzK1muGI6MFSfxgbloPSnNPK8
l4WXmM5tc0Ys9mQqFkQNlBKgHfxsNwkIW0POo3e1pvRDD9RuTARNo6RNoLuiVBhyzZzLdgg470Nw
80lxQA7g4odd1arXXUaNDg7VAJ2t+ESMfaKid+jNGJPu3J0PBHHKDHow9DGwKcZo7XK3Hd7gkSA5
bT4eCvi1UTyBBD4gqniMQvl5Z0gJ/OHVB9Rnk3cDkGWRtgb/AqXx2FZZ5Rvjb2w34CxvjafdeiDt
2YCzbs8NkihjHYoEwPrU1NxMhVrNkZVm9QijsNq3bSVBeVV/6OrkF6XR9hnBELB/OdKBlP/sTQ7A
OVxsEWkeCN4w9GvSKLBzU+tZm5LamOZOJnqpd7ugJHRtYlc4bDYRPEtSc4T3F9OK8fpVL9vrbXGS
MKNZ3dzodA79mgyrDH91knIpXMkhRJL0L7JZ9tt+RnQn5JmdBrUAQGWhI/O1vXtEv33SJan+aSnV
9xuwW1bPsWd8VC93GXiHjuZwsfsz1qJqeO96tCrhWI6m/Hl5N1sQjorFkJwcnxLZfFoCNWaG1Xrw
qjmwupckrpBRP5WH0D5yRfnhLDT0kQsrxBYp1y1qewSywH/cm8DOPK+Cxf2EdWZKlqrEE/XIoUEe
NkCX3ethN/6nUz6+o6If1xTSMO1ltjs/UYZpGkY9KJjjZDK+pT1m0t+aWiFQOTwb2NKOrEtxhZ0H
2ssJIwoq5i53DQPZyoahVAg75s4bgiHUJD/k5E7IrcW1NuLF1dMX3VQv6hQqWqdIcUsZaniOpXCd
/n2oSfSp5TwRVSOqw2oLqGgyfttkrn1y6GvbKCbJ9NzenA5vi85z39e0X7lMiBMuRQoYDcZnLnzw
svL60Y41Jl8nPwtv8mszSdfoD2iOOhsMMWjIrAYN9o7luWnf3hDQCGCyc8MrfhaRgd4rSJghY9rI
hax12aVqBbYEM0q9mrTNf6N4G2lxkiRNZL2zfZF5LiPP5wbbNO7Uaynd+18tUSXC49AM5durzWzy
vUjt3tcYRrF4CFam84X6yclXfqGLTSFkUgpukzkP4MQzUVP4itNiLTMy0dm04V8uCJrJiUqi//sA
VN+j7CxQUTnjyf0AlPf4GO8zELLObGziO/sTYGqlgcQ1FI0bWHkuhNygKTY/hDcOG2Wox/9R6INE
17TxMPAR+yJNOs0IOmXeHZmTVZGs9WmIaAdJCJhI8dQCZbjQVKsRUe8J4vEp7OFnKM/EfaLbegN/
oTJKnj4MHgJ2RXsBrJlghUQsze7ICGXufdaDfwbxv+YKZlp9O+dZmi3FGuQYNK+4ipsePd76cNTK
rhxlg8W8iyjWXHXtvKl6l8cKoNAKPVybWTu5ZS7q0H5BfXe024SxOQK1/HZUl2JUcsYzH29IoOOz
Rn8HD2KXbGW1ccuLfMGj5hTMSxhRKDQAEB5ntaBd3rueQLPY85vt1semvl2kQRBt0QSTnR5CBr1W
D7wCVG5Lxd7RJ10AOFxKKFEqeOCUrtVQHQoi3rfgphnhcSEWl4L7l6yRO/QgC+WBB5IbOtjybbvB
HG4DcUKCeKIXMUpIiy6BaEnjlUw6ljMc4u+GKAdoonXBgCgoKLSxk8ovUmbR3d3pRg94PB5QTUtQ
zwAQ+FBsTh/w/hrECGaF3HsTFUvbW9ErG8ThnuqSYwg9pyb8sNNhcd8P2gQwDDmd1dxAWIX7veIY
cMXj2E2vRZ4xUpVIZ/9UghUC/y5K9TDNVM+czLcoWKLYvzRGhE2YsJRH1Q8qYnfe8Zwi0NhuUW/e
N/sca/2DABBjPDn+XjNFAatNaQLsZSr25k9I9RB59liWTRNjh+Bdfd8QBvxL5pqpG/Tb33auDNlv
lCLI7QCk/EQVFNscWz2HNT5mYVeXdxXgpy3ogHLdAqiLF9+PLdy+efUYgbT3BnToXs2vEBWKUW+w
A5yj7bqez0W8zYZ/t5UlVh6imOh5Y4f+tkmg4URpzuzjF9Z3wcPpEre1NnIQEksWoFG0jphfaV9f
t/ejNrrv4LKUHuv/KfH2H5hHum6CDLjKQKxZu4dvby+e49Tn1LfeChojf3gS/pyPnDUMC19gtebN
KDawKwZeN0EekyKEg4Se1bc1WlUItqd2f/A7lkEi8+7NmtiwtlPop6cUlZXSCJ1rLl/LeEVyzrmu
oSzzzQ2A1ljqr5Ca+Tf0KLH1mtElK7vSKRlF0BQX1uuDTRfuL+9BBvmpIJRQ78Zc+vEndS6/NtJR
oR2hUZogO6biEvJVwh3betX0OIgs9JUrcVu/eqhUi2s7SwSnDx2sUmBof9lUHtqOWZtEF7AtF82M
wbKYu2oE+i4yNlpRgQgFx2ZDeDkfwD3bOlfgy8dnlWriYBpD8tUvnDCdTOYAm26MCfMRpKmPN5rU
x3rEnvINKFRxhT1y9Fp6jRQ7kpWkmKGQqX6WcsXak07ImQfBzScaBGFJnGnws/GqXyCgnPzZxbTM
RPhOCy6FHJv3mlt73IC5yNLh8yrwM7QJsa8BVf2inVhAfjETrx3phCepKUq4YgQmwoBteqD9w4ld
HZ9bD2omf53e+ZEBglbws/KYMHNN4sgSZxW0sHxndn1Bau7oV8kK9pVJdXwnCWKevMeFhzDqvdOh
9HS99vg534d9NbaRyNkdKBkuv2+eUc2+4BDZOWROfznv2V7eGDJFQ13wE2xoTMTN++f2AX8bmb06
WB1bByC7ZKPyJ0a3jhabmlN64VZVSB1zTo0bX/skDZnJD//qx/up6yFvOeuk2hKIWFOSOgQoCp8m
5h2bkfGMLLh0/5RUUqfcwspsObB/g8c98IJnv8L0l3/aveJUxh91VW5cp8WRrw37JICxjiAe/fTI
h12nnuoWu9GcOCKz/t0n6IvIFTme5Vts0EcQrTW+XiyGh3VRp8Fuyyc4SFiZrbU8luv1d5qbRmQA
ZUHU/Tm1H5O8y7UfzAbGiUs1kmGgL4RzvXOfS2NA32ikPju6lJ/C/Yb5RjNhSkq77mCv1Z99eZf8
UqcYAZtZV2aw4PO8vj38FL0nHE+QlisW3UYRYtOG0qmRwy8CHLPGeWlIxvv8HLG69EIcN6C8thPy
LHJyl+rwC+qWyk2NwJ0Oqt4LeNKeEIJdDF0xJUJzyxLcBbCaF5t1FKWnN6ABTRDUcfbmC9cA5dxj
8L6tN6EXwZtVTsxJ6X2BffqG3PWXyl8mRYVN09Ma3T28roIOqnSrIMqBKc/YJCEdT/Ar/Z1rZDKj
QZC3EPtSj/kr5UuEU5sj1U3VpCeWt4i9orbcPfWJGj6y59Npn2FZWdVv226qi6SgRR5g0o/42eRw
4uXhIp/FnzSrLPxHIL42nPKg1po51olQOeRmRX/Kv0JJM8SvVeIAwO9331CWCDgqVMe6XlwqKbpD
z1aL9stV6GCd5SdUunvFtSO9Mwcrhni8xh/Rywm0eLMqRcJ8n9nBa0Ar45cq1vimuFt73pQc1bvJ
uz3XvSesF6/fG9eGgfl8uvbJ2Utpj6SSDNiYN1zMfH79Vkfs564wvkODteDmy+i2mCnXJD9Kyhrg
eK4XlFsEv9naAXrNhhrIbGH8G/o8oNXtrC+xnhEN3KwTzWuRv13p0EvW0Nq5yPQleq8w98GR2tQ6
ISqMCLzenGpLuvmqmzrepkgwdmhL5OX/m9P6DE08llCr2XcV0gbMEoK0oBfxEW0O/d2l3LV6ZIWM
Of73mIn+wlAag2DFQjXNduiNL2ufLNtU9bQ7dKZzCYl+lMiOXOnavXZgE94wiybWXpF64bx6FCJ1
aMEtNXIvbfGg/kAKYOIUHqfs1fzYZ0yjKsGeiRPCONDl9b2sRDda7hpqidy8y21Rw8iICjtBMjIJ
TX1drlY0iP0D1WW1o16bb7r3fUx7hSN1r1hNeKQoW1LCgTgl4w5bx1EzdgljxOIaA7m2GH99yAd+
9JYCEVGh3iPT4aWmOIM/sBn+iigksM00w9dGY6FKAVwyrEB1HqCuM9Wd1WyuQE4eUgtnREN8LJ0E
WkvBgIy3qwYRFyauQzN8e/yrGk4D0C+ZNl704GbALTJlLt1QFbM85Gn0+hgfPB3dN/z1VOSiZeOW
hbJfIJtg8YMK9IYcd9EWdFRT2wrnRaVDDFlRn/SdMDHxrvsl0HJcxw7gMFEkSAgWvSxrN5Zs5p1h
d1OG3jIqcx9BNTRhd+NRXpCQCe6FLsFUCaef/NqeknT0XwiD7BisM/TA2kWHDakSLF42i9YHAyGX
eQEJzHPzzBNNmp0tOL1PQWhDUHe5j/OLVLvPNIJLY+6K2/osQHkjk/lGGqC88wHqQs3m8+zqH3rM
9+wTxaL7YARZpZJUe1IJfxhUTGT1Nbo+cn2RB/TU7xsZX/hNRwdqRuynoVWJE3rzZ9Ziz1VTmIX2
I51PAiZ28iDtzUmfFhy7hOWj0xk1MFSzXCfwioWI8ZeIyjjASZTF7HEoCM8m/FzOdRMW9moaU8wO
1X2+38P6o912yRo6dVvxpnHgd1MDEw6ix5/dUrIQsUw9DQmNMLqL/MRO8gPPgx4rtmbhvrc+oV/w
vgz/7bf27RGsqzwfDAFg+nQTFQL/cPKOe9N44seUW3WKSFYFAcDllYsdWmy9e0xJRtPkUTo3BiZT
Ekkf+IIpsQPyc9Cvy5jM9/SGyzTPlwi/osJpE0ECc2xtiYXpI55lrMLVDWQPvg2nx2K6SojL6UBu
lYS+5borvlOWwahBJuXXoJsIbuBxTnyR4Hg7l1NlgeWUApnX4dNxuiPsB+9xCtRpBubEvcnZ1TfD
nneUntPaM8aCBudLFFI/ogikA6CBSP2GfmJb/t5+tLFaZlTyzvCK/icviM36jcX5SllAO0k3DKkj
7Ohb6FKpqtspB6Zur1DTiYcSfrD061W1cJzd/Lmmn1nqWtj7AZFC4duqhw25235K1oXgtbFY7lsu
vCpE5vaKTwuIr75fHLidZ93FbWMtg8I+87tvnA5649NbeAXvikMhEJyBhSA7sfXAKf3izpmJbgtd
ocoScJlZBj8w9FhnQA5wnbJu7ptQAx9AmGnPz6cxTzAHdAMkMD7cCjFjsUajX1c4Nk2K7BsEqi/O
61gWR2CyhsK+Kc2hMCHM56eTXqB1lpGjC/FoR5W+XQAEZEelIV3gHQzI9en60vhFKjCkiLIA/aNG
d55Vh5b1gRCWOI0UpHfr8bDuGVeq1Fo+1DkP5Oxn1GZbMuRDYAgXRMBq4V/GdL4bkppbuy1FWJf2
b8SYYbJMkg8qXjh/sYqCVgFwymsDTQVENP0a04m8GsQb9o22Ec3v656CUGEXM+DylhzfDm6J7WwC
jo9wFKXPov3B9OkXi+RBkMCaIHkADFvxq+YyGL0go/U+tO5UrkRt/0u7dMSeFEvJ7M+wbQ/4Kzek
qd0kp/VJ4sIIQ1jrBlUOqS5JVSId9tiq9mqP0P9vTkl3ONUSUr/vkA8DykxBhnnYgtBd0N7jUUbK
qo8yPa995QccSQewyi8eip3w7AVtttr/bRjE68wGS7UpWkMX7KQH2Vavb2np7Ku1B3k/zKXSsTPk
j7XGXC6TCBHRiH6jqfzWGks7k1EklM31/e0PbynEH7Y7Pi+03HC7vndkd5RyPmODW5B8LBGQBjJS
LunRNsnUJl3UNtVqhwjyKjZSDnM0bKumNvK81kimYxB+9d03u/OupRzsOTfoKs+WKyjSSAV4cPHQ
kbLCkJncrAOqiulGxjCLPmzKycvY5FeqhXGbsoelYglXbgtS2wUv08leFOoZZoMJPLfcF905sGnG
qlygDjO5y6NkexdLr7R78/XpC1v6qYVoDLvCSRdSZ8gbhTdaGs/dWRBGB0E3SiWnVFGTdhl+Aj6Y
JMfBA5KN0PVaTELWImX9vanq63ZTFcBn9CRAkWK3bGmLUoRgwp2Vm4M91tFVxygkSRpOLMuVBZ2Z
zOu2JoFA2mKKmYq0RCyCjGkVc7GPUPIMOWS2+P7zSO6vyTwVtOZD3omYiJpsDEp9wBC39pLtXTVJ
/UB18cehkKq7cwC44l2+6ClyaIDfZe/p/JRFEONOHDOLHJDfA1suEAdmFgHMbEd5hgP8PwQxVjiB
C3dKpGff8Q8EImVd9bfPQfJg36UrMzu3GNmLD20kHkjbl1jpgv+ai0MbPQPQHn3G2Bd/pZm1gZN7
X6VKAccgGE4KHLkUw5ljevmYWRQ/RTCtTL2MI3h/enNi7KB84n+YK5tNSakofi4W2vYDxvKfaL1n
FSkUHZHrjLYuAS5SP9RiZBir+M/GKJIcL75opxfcrVq/AMr3gwUdrBxIvz5klHxCPCx3XmM7dXfs
xsIkzoDikaJIpXD3ISdw92n8kYZFQYWvy4jmOhDItRO1/lChQrqQHA940x0UNw0JGlhoUM9lKqpR
JEHRsEDPfdG1UR99OL7Y/J7OVDuGyaNXmJhPjlSLtrdT4pmNVQAkvn9NRNQZNqHl1Fur7fKuhVbi
BBCRSc13F18AGUnGXBPXqCZxYA9fsP1NL3xhDeZuPxWPkM4RhRtII4tC2VjkcVOGcpS50wsJNf2w
rT2/Lp9vHCEMn9zhV04E0Uz5ObHGkkLVLzMjZwkgIKGA/KgvICbSQF9D6N473a2cbm3BvWD69d/8
SNv/a6D8626oPZIxyNr6D0nld4WegFdcC24yDcAg5RRIAHUcZKzg+lordhRzUYLPHMNdFM25sesY
tbNEs93/LupFTWjZ88zBJ5/w8TCziuapq9NwB7112wlsCNTD3WPw485cSmGdkuN74/IS+akB7xN2
Rpbg0F6GRoP/JsuUUoj/ZWjVNpAt8cAU2uAz4wUFdnzbEUaA81pYhmQDauLE9cEaCsJmHNZt77AQ
qicSZQktGMB2IEXfcyt6j2n8y9M/KDqx9S+waRAC/SJ8h2JrDPu8oPkNrO4DImBBs6aRF1kpWzPw
JJTDstHbC+f5GSQaDrXJizLJMbYsO2tmAwPMCDjlGua/Vi9xVDQICCJOZolbtTQX0lEvJGTJLPAn
TaGMf16GyfwqHNLMpO4oA268cU56W9DW6k5nlkL6Orzd0OW5jtT9dHYgHscaOVp/4hX86gEpTig2
4Qn8cLyQ0JoPu0E0VgVhavVZZhiUY8cK38jiIbhs+j3HS+jwfzlkwK+PbeFeeOUF55Rvwn6wHLd8
gyJd2HB0/bvZylNmrCGhTDlXyfiywdfrihRyI5okYanhhhMYXWDKqVJ16eHAJXyZLkaWosQ6w//F
TKka5hGgWo8Bam5Kr+Lea6hQeR8VTbADphkjLp7kO6wmRh+b0AOJs8Ll6Ewct7WRms/MX79MQz1T
yn8eKbft8/VhjZRUIGDciEqKh4LsoW/SuPw2R+n0RjjpennV+XnVsVRgz+ESPd/ptXD/3f5nvdPb
HBk8x6dowXj4l+3XB0Ab4Ra7L4+bVvaBd7sfYVfDxGJMMqfaVJlKLzu6rNGlWDa1kSKzQCqiqH01
14ZONgYtWqbVTopJfb7QrEK0MFKT9uFewOV7swJPz3gXOaCnm7lACHCisDQP2pmDTe2oijQlcA8F
VuEgQoWd6l15q0pEWv+hFeKwO1uB22NIYSdzNwIOFij5EHQsGiW6H4nJHwsqPxVpaxtSYaSJPFXX
cGLiKkI4h9hl86DynDUhg38hfLlJAk2tXPlWArlFOqKvWm+6EPHNRJ4Gy5B9xmd56QCW9K3EaiRw
Zb2P6gJwvTHJCkxOzkPtktbORG6+nleo8QT8suVjKnQzfrm+jME2xGvGp8w3cFn3tW8pPlm6K/rj
M8Qp+Zk3xd7YRooclVeki0/5DtUkM5fxYBgS//w7RQ+mY7XoCziP7H6zhvuo+jFNfmhwn0PBbVjw
E1JXWfqQHjWnmiKYygktxFFrjAA5v1hFdd4tQEB2YZ1SSp+RP54S6EQgE209vFJ6WAUItrPUc89U
c+2wIfLjUXXeW3gcwGakw4UCjN4sLGklkJZ6JY5ntvy2IH6xAe6e1tJcQi5w3xNJE7hAeFzfaVqA
Sne9A+eEg1Zm6i+9BJ5RUnfaTZJSvMY83N/md9bEZcfc5eUXbFke6K8RC2P7bEsMW3Cmhp16Pi9O
s78y0+TBsvidQaXgwee+bNk6Yy1BPonvZeuA7g9l1b4C4ND3+N3AEt8+qh2Y6fsfH/BLjWcMWIOa
fuL2qgNRXrle3Rr3NH/WoEUeMESRPfRINoGtGgEduUSH0xXBpWQTuKcWnM8gSJTv4PXgmH2eUZ0L
mm4FeFyjlYmnBeWG35z5Ol58YqPEkmF1yUAPCOsoyBaZfPlg0S/IXMe3XyXREiUVNw1048hEfZWo
oQbQNClPqGkxJsmJ8pAeSX0cX2+1QPZ5tb9O+xQZLBgKwq5BDM/dNvgSjZEMmb3Xt53wU+ICMTGY
zgBFH6fX4A7e8KmhJFf2epRwOlC+Tr0ixhgNON0CLn36S+szNoQGNhLsiaTETnaCP6Pr/WpKAnX9
rOC15Q08ietTLYqsa9dh7IAG1qqv0pnpWOo+5wijllnpt6Z6svHDWV7Gk5DpTyiCa58LyiTkdIvj
w0jxgHAmpTKEs7ezexvEyAXU8H9ofmThClZOC1HwrkI8rU9wA/XRaICqAThwV+91U0WN2LPudZHb
I4ngyOKJzT0ToYcNlGTHwpm9WU3//S1efAILg/7UUsJw4FoS7Xvu+F3cTVN/qAvSMJamWNbGu7yu
zTjO6LxSK9kbGAbsthDPd3qclFXwJQNXYV7dRpF/gfL4UhZpHjtWrcC6aXWA4eL2Ew6E5W4sv3qs
c9nZnBtjOVbZSQQnKnFLPdIN4TXURCImCbaIVqXpSlv5NsK1d2TpyYJFdGuXdU5UFGCwyWOHOfPq
AGxZMu710CHxBW0wi6laYIzODgRLf/Gr2jUGIX6QQQ34qOtgVIblGyZCcfbUK5HUoO/UPDUBMlnZ
H5uhEgjinS8CfXSNTwSVioV3zuK7KFonoNAPSDanTuaLGyHGhtknClFIQbB18x2Khee5b9WlZLGZ
wvTHBMT0x6oaIe8A/YF1SsLsFqCbcAwx7zPSedv3k77OAYt2AXAMPY8dh2H9tBntQ6cg3ByFphiw
HtWXhtZNtU48Dr+QBXxRdG90Nxy4ma9u8atmfUejtcumodD//b0vwWzKugyEewDDiuPgPkta1Vjw
rTkWudqtp1y7pbWGOF9xHWF5TzgM9K8rh+cXSF8erEgum/n1CiQaGZB1QudKwm1We6kA6uU2PRgc
SGfdwlp12C/GaerybLGAgNAu/rl0FzK2zN0DZJLoO8OdjhOazL5v/fyYWYyOEzSx+YYfYuhQcimc
WufVPejdJPBbpzyFIG4qQHU95K+0YrQiTXXnBO3k8yvTU/GS5zfVloqVZZ+bt4ZTH2W2jC+6DYy8
JAeGUnslDJ+fcHAxE6RhviqD2nMexHl9p7KYeXmXQLm61jj1pOTFwjj7R72UkriyAlSe41BpoAVc
p15rbJbHazrSbTaVcOoLLU/Y5ktpqfofFssqo5TfwN0mpx+l6k17xbe4uJQachZsPe0s5acL0Q7t
9f/zT2wNS86uG9Rc4GAyiZvw0xB4Oelfj0jbl9KWR0ysHy6fUTqdgZ2bW8qVWcRoi9QqmN5UDwmX
tXM3h32qzByMUTLS/E1umq30vzCDSStJMO4gaYgxzjWBKG1p9ObhZAYfW141XQ1QFdPqPHsoZLFZ
jEbeb1WMHVighchOtnMZKLw1m8I+M9XYplmk255msQJsszOmUZdVwnXX76UNmNq6s3UJLOhoTrSO
YKtzw5FLPrV6ao9JTsz97QQUOEPOecbHRKFKFnR9d8HcIFyP2GeluLNBK1s1benj6x71HSid95Dj
yqnABrIqGGNda7J60b2PaIzTXVuDe/DcMIB2BKVFfyORgP/eM0H0lphnNZmfkx4fyPaWkilqlmQB
gcaMrBKGyNf1Za6QRP/glVZ0MPy2fIYorr/DYclEaJ6SS7EymjJJ4aZ71JiV2CHQXsvvm1xFC+zZ
yJT/wkyQAomwuws5skqOPKhdnb/K9J+uqG6HdPVQtIlzohmbUIDfVZz6cG52vPC1pFGHJgPybmci
N+i4Oi+Iq52Bi10jsfqqd1o2zKdbuT8zn6KH0MI39I4XDY+rWRPlsd0dwKHIc5bsD20YW4ziJEoX
1mbDX2EAf0C5TSwoxNf3CXLAr/98aNpD6n6lmTd4GCskchZoBZMvbI/7MpDMGRZrt9YWiu/rfJPm
BJkd9mHP5bHK602QNhK0EYexScyVrd8owy13K1C8NEWTq++96UhKWPP3/IAtjgKZ9n/Ma/n/Drbs
710MgMpworsDuvu5wNznhnvqKPH9V8BE3HuqMkMewj4MNJZmc31HTdyjC9/eObQYitYE6aimGCRY
YJiXAz5Pad/G3BWHb/4o2ERKaoxh31PU8UNl60sUKeCO1ltjxGqxjXSJxZ5KY1rm7oVvFAn0ohiK
iu7uhwygdQzKFEyE7DNmYC6R5nv/8efEZV2zeovnba0WxPAsDr5QuLIA+8FOW5U3QjC9b5gRbPbY
0qyJGeVn2Qe9FaWqyPo6QEtE0SdVpwTG95azeAF3dgY6mZZQ1febJURHTO7LxTILPyqC5Y+asmlO
IDAlxmJjOdx+3OGYcjWUAqQnBJywGdOiUfbZC6QkLY61Ig6tksO1rL0K2hNLDrb29Y4/DNJyHrUW
RbDgZIz3knnqt1zYtiGRqPl0G22eUfVrMcDcipxdqUCFDWjQLe6k7K9wEUlVfXG6Qwq67o6LZ0fF
XqmUWCuFmSEKcm53hzvVofBiGoIPQBGfBdsrSDLDzRf/UK0t68lXRZmmXZFccfX6c9pGnLE02B5X
5KgL27sM9ew9AH7mCABv0y2VNSw2DxxcyqparF57oS48kx4nsMSiyegcJEFRzS/ptj6UKMMt70K+
P5zr8Now3hG8BnO2mTu2Pqt92j4HUFV3Jrh9eX+mCCq0Zbjp9Ya1xQPfseeWBcJJ/6Fs06RK9F3q
mldSLDSk6ZP2Xwb+Jm5EYdK++2JSprGguYKaKgx9+BoDbSKh+2xvDedNddQ4RjmD9lzYSwpm71CM
Cb4A5a3cNcDH/hh2XnH/wkS1b794eVX0UepvMCuDw0Q/XCCLuLyjCBaGBZrVeEA/Hy5Ut6ri9Cs9
pL+fS/Dvs+4EqIvXZ1JdVBlrX9pNrnIuWg8dvTXUMsDxrsmFnRxbPpR/0xZwpjyUC2HTEKbcWBLP
ysbZZNEP85BV6Rt+TvtOiTQ8pUQCHlBaQfLFSLFuXpZ0/jbe4v/9nhF/nesbMzvmKUE3p3f8PswJ
7PD2zsWtYsqNwt1kdxmfGPzdhq0Jctar2yke2zvZnvNLs/uHrpQL3cMt9M7Wa28fKp8cWJcEkpsv
/5+V1Ed29OWS7lJvwfx9ZSQsZXstaQOScQKJG7uVCb7O4fQV1Y90YK+s5o2kEPyw7AjVpEOrGoD3
KMdy4+TAaBQk9NCI2Ia7pkUfLkEUhF99jjmPn3YqgGHQE53E9Fabnwu6pO/A5+AXpSbFJzZzueXB
9xvy+Y/u8JcO72T2PIm/xQr1tsWfgKqPjCWCUEb+Y2C6RMHvjxfD15ld/Njm1M4qeP5eEYZmujJ8
Qap6O1SXqhsEkFpcZTeECwW7Isu3Cw6VDmg7Ngc4xtF1ceeVKqrx/pEQ4x/evKg7XsBGaKjOoGDO
nVRAIYw1QPiNDXZSOPWC0uY61fL6Rb09TrTSSYVbJ2RItpkhFIKYH8zLlgTY96aoZ3wXc5zvC0jt
2zkC/C0lW40haCoxgO2EXKMMG1B2PYRppSiXRCnKjVMGS5p3pBTv3IOM8cJ4qdrtbGKpSzxWVc7H
LeqNIO8nLSxv4385iSIi1r15nllEIRGZEo8n9DrAL3D/y49QRtb8ZR7TJjwHiBKmVxbozy8t5KSA
4fcubdMMuTCQEExj/vdkKx8C8+H6+ZfdIcIP6e+8Siwer0P2OFX86Ec17B9UygGDxjXhxIEUl+vD
fWHxqH/mH16Pv4rqooDf6SsORuySc9kZ6SNwENDBvcZzaRnsZ2f6DOCIPPVkmEqk5jMPRlX0K7YK
LpVbsaioHF91mAm+4LzeOvhVe11EVM9iZKOml1IsktAreoiCYfEJoDL/1TVo3VkyijDeNbRWaxoY
wpns+NUstSkuy7TU2v4v5c8z5az6psxAo5D5dJZ8CzBmHOUhLw9ZLfjjfavUbvk/DaCQU3qSMRZT
3UROqsZVSbYesSJcAXuB+jrY3iU3Rf8wnp7A3wI4C/TL8527PrnrPIV4XSs42L56d79EnLomqpFa
VpZnogpoFiF5X94O2KD5KN7qo6dQAoTzCuV740c1ira5annZFBEKu+GpwTwkLdOrJWsw3uWYYTvP
ak9jXj3SJyAJXCBNVNM7hoDGno1Kzqq0d6Lf11OR5oPBsE6W3gujHS/Epzxf6LaBd2/zrsVsG8G1
7bt4JWEW5LlF7JbfEQv1uOLZ9WTAiJNw7rt0sjWMWgq9G1d1oewwAKD8wQCYkehkjHDhLhjNLIoG
4uoLiqJUZneF/a3IyDFm622oOJUCzkQiUD6kfcd3gmO0oaJCjM31rKXyX4vRxnZFSLyKGWXm+ePR
vCKHf+CL/kW2DxgUfr1IYg3+V79Ur4QBgEwbXP7LC8MxjWGvXusw2nuiXzK4jDMqmkPESi1ZjO/8
iGAqKG881v4TRWahS8tBi17ds9jUKs+zr7qWXoP7zUCUqTX4RCX1JmYvxcDg5rsYfnPztnKJUkn5
PFxGGRYYL2wwJLWgNzAfMr4DCU5ytDeELhnzbgt2GalBfLud5F9wic+cwwu5U2SWc2GThZfCXMoy
Jyn/Kbss0q2kDPP9y+ErCwE+YjQxrykxmc6OPJqQFw5fd07DsyrU2BzcKxC9OKSn9pt8VrtyLzbB
4Jk3J/IAf3O2iuI3y/t+T69OiL/U1JMWD70kxBLwJ4GMQczUrtzmthCjztsKm0UGcyUDjb3zKrQZ
Fal4FzS6HynyYFp2yOWjg/CbKC8yN8MBnd9uR7AtwE3wfqwFnTaERqgd+eI67HsN7sKLrnV+LMzW
CJ9RUL9jwpLsPkj7U4NbZE4Ybl92F4+0vDiYV2ULdzP83d8yOFk1oe8i5rm15I0tSKVRVxMpF/vc
qwSuZjaArHzQk9ekabKaWiR+VUtn9My/72U20He7qZzg308c3GbGQPYpY04D8bLrs9Qg6UuC3m98
gCEAa6LoT0vIitvq3AoAiWKVcg7Q7A0/Rx/YULi4rP1r0C5EnayywMyJy4UX/Eqnr4Xft/I/Nab2
hAuZHWy3kGsfyw1/Mc1Zs79gnbHjogt17G6JKAvSYnReyAww3bTFLHjs+LxDtVrk8THhH0JhSuKm
Bxih+9TnXtwPjZ7TFft4hKMEW4TEOYJULsxewpfwKiroQ46XyDrcO3px0P/tNu3RjlepL0zZXAx+
4xiGXsTloew++zCIC10ehuZpwamofyQU9fHY30LkhxDdNWvEzfnRcAY0UA44n+zHqRI7+LnZQ/bn
MlzcG9kPFo8voQylg+yp4DYdrY0zqeR2sDAK+vBem2PWhOcH1nwhUJtpRbkQjyZ7Wy8BZ2BoHCqD
t7GEEtAWGJyHbppcoSHofTI0pG3mwPLVL+duTdcl6TRhRUFtDOJH9+ozMVuZz3wKufR/qkWJDLuR
3GfklhqA+5X3XNAf/lYt5nF/96xz/DPjyGPPuJndrw79ESeMBpJihm8ie1WmKaIC5DkTYta5mcl9
VCxjcreVX5AS+jZhv/SGWiH9N4qtqDWAPkJD+pLDz5hxdjG/ke2YqqxBU+x86Lce5XHjLRfym1NQ
+bT/BR7zKVvyVCFiBjGgVWzQz1ex/uF18sn+pyLCyKkpanepyCnK8Cxzkf6AQpeG9aDOCgE4pe24
/14tGKUcMUOu2s/oFa2/irzUjyVbZOpe9fk8hmOxwDhpsJjxVuOutn7Jhp4wGbB2c6Mawnjj9tb5
npBuJfXMo29vxtvTAERZfyU0zs7Jn0GYs9LSQTuikA+iwRq4YlpX1V4r5JnEmS/cBvPR59V41ezU
ZCaNFEREnvUdtaIh1D+gFe/OE+oZdAdWvB0qANNx33xY6V5Ko9JccaDUbq4gpkrAlVyP/5Di8/RI
Z48BTMAPI4liGTAaqMZ2OPvLwn0A3QhTW60p5aA/ZGzB9VpNVFa//TWnUcGEl9nwNNWlhFrXXREI
+ciO3KM7BHGz6YjS17aDh28kiW6KB8ws8fkumPjxLAVcpzy02xTbyfl5ZdDUbQbkohkOihx5kWb4
2BSmYNKEvUlrTzAP1zyh3jJXNheagNmKsPOvHZwmNk47HT9C92YQ2Gt+i177tBA+b3Q3EZM1BtRi
NGNn77TRr/rME7/d2P/SKIh070UNMwA7so4WOtDP10/lYn+BH8E6aYSmsToc3RuOB4ogLPSydozO
BUgZTtkO0nLGPUjH7Z+ktJNaWKk0AMaBbRYgOVRQlKpUTyVZAoFVwzbfh4SAEUL5+ZL2IYhACxAO
kGJX6ji7oVwiTVtAQxFhwGprfU+bjtPaLO0V91S+SLGAgK8VRP8aROnVS9u92OITJwcnXYPGfrtU
bQxbEQjJi4sF5GYCmsvz1pRG4gsFme8fubR3NcOEIVC+aPX/VQEmPOW/jEGjWWKA5ntLgDPGgX7u
cnMzIm7WDxCUsls2fhUDVXQDgPXPVi2NjdbSbwNwLV74nbnkbml6dP7W4Rq4f6CybLE5n7GDmy0c
lkNbS3iqj71R+QNNvKnVPTL6clKXoffztFNmRKHvJQJEp9AngI7LJRJkckYK2KtVGSP3+vHrXR2O
CNfklRYpEuo0fcQapAPYSdGY7daZwA7vjqpGbrdbKnGioNE+wuTG9HmkaOzV6zOzYp5JjkBuSPxu
/9oyIgCckVbtxHJke6Dbvwoyf9d/kg5p75DXsq4XtL+7/v/20eSrIq/8fTDF+4Re8wrSWHjkw9IY
Mt3oqC1zLx9lUVqpJ54xcxkU4ZuCOxqSxR3kqrs7vw+myeDFr1ph35T3eWj8dTSKXK8rij72pFZN
N5TW2WKniTqGmBNVrIQjLen9SyJ6LTlRZxyINthEnFHAjj69ZFRymiqsRDbEaZ6b4H21hzauSp7n
glzatxKzVd3IT2RFILeMLMKSwRgBIvd2kJIrYFNcy0jyjqgP2gTB5TuzlFt1XXHGH+6sHSvrbFnI
SDmMcGpbK7ENNxTv+1X+SRQ5kvFbhme1DVVqIlY+zebTs5i8PQO2rfdwtiNgrSlOOaJAJy3jPK0M
wcy1jh4lMY+LFRVWLhVOsmuh7izsXqE8ZimAqBVJ2HBnOKdgTsxLWDZiFLGZO/kqYI9WXl79wftl
hklvjMajtdp3T7zTa20bC0YkkF+u21AfshJHvMtIJRKiNV5hHRK3k7AYeo8Koi6x7muHATGQDCoW
0hS5NPTWP64Dk9xq0tr0k6m6baFmOcieQB3HeC8jDp8bOOnEAUgsv6bwVhkLgvA2FL+ArnvNHpdy
VHrkvPsg0qOBFFjMm4YQxqaW3sFRPjXv/V/82ent79wjw7PYCx9GpFO8NYLTtD/Gt3HZLCa1JqIN
m5xegGXG7jMWqGLe4mBP5pYh3Bl2Eel074RNMSBxrzLsvu4nkcPwfp9XPrPPqwHdE/lbrTRTfzhw
0GhKsnlcDQfMf45to6nDLdaI53MXnQtzENR73nc0VXv6P5iy66MAZNOiCVCc0D57d38IhpBlmxKM
9/bzaEK5210USr/E7JeXylxePouJvvG4xJy3KwbvUz1E1L/DCnH7s+r4amUedAdo+gf2u4yWMKOc
3PBPMjAKEAny+KeO2jNEQW4xG9g3orxV3XO8KLHJVnSgawTu64GWdxJHtCJDz8WtOohBpN2x/jrI
Y9C01ADXNAknID+Kf6DUwxeRr/qXETvdJk3yPJzrbOsXPSKyATmn54S7RcOAiY2CZ+jA0W43ei+7
LnxW5W/GSD67FKVZNRF8A182MiGjvFTawa1ykbPYEuazd1GbRiu6ChdaNJo9V+QIQuRubFb0EuDW
HlG0wV5hCoztHyBs1B4LkvRDFwOlP3G5akfo1gC0N7g4eJy+z4RzBwtsRb4YLzwvQ6i9kvL15MRQ
qkjLaBi1rOb7F8A2v2qPwir+dkA9v8suFrx5c5x6a3hGvx7fcm2H1FnxUHwfkaunrIiUb1oM2O+q
wA2fayGbfzEm2B2ExdA7B6xz9drsd7HP16IUFkPnetg93VgfghOdby0kUBIpwFNcrl5eCRz5alSc
4EQjM89Fc3c3vHuo9UfT9wO/e1fxQlKM7iZVk4DhNpjHHx7MLkFppAa0PD+hH0Dh7ymr7XTFCBJe
M2qE6ftSaXfv3aq8jzuTf6Jb9PetlYngTlr8upccmYWogC1aax73z7TJBk8x6uDLX4NGLxEZaXGY
Hdkdd8NCkXc2fJmvuhTuu3/mGycumgXC8/7rEt4aJWMxLcY/A7dKEeH9s7JQ3ogL04/dLJuPMDGy
NNGVn6hJIldg16QTN9qewb9sZqpqUlYdBNNM2EKlPOcG9gMszLN69HXYbAAQtt0EWSX6KxODlEfY
gARSZGYkpb5Jb3Zp+H1U8VVTmTSqM4mbnyopZUNXDInNBHP9qSKdVq+TIZEC1oQrV27D7d8P0UIx
V8gbnDizqzW9G7xuCnt2KvwKBxDJ2tP5dVpcJj2Gyjag4GyQq0cf3gQNN7QNeMmWOjbqtoHWcsoS
eQCRVL1kZVwlVCWZw6QZecvVRGO6ljlTpoLXXMnJKITHAdQuCuLgA1teFZz6rYcgTlT2M4tAtYdB
1eXmuNDmtWM4c4d08gd6L2NYhQ78Tii6lhG8U0UbnTzlOJqjH3dhQwwyMJCBq/SNF9sfayUYe+f7
eUlIIdh0xWIhTwJVml+ZEcqRmEJqMBe28msfcUZwijGQHze6VUENexryTvXmJoiY84lMpufvURXl
ZyMf6F9f5QLHQ8EIUcy96wxdHkehQiIK8WCKSOGIq/V7tKyGc3didfFmFXfwzGTSpupVf4ZMRE9j
WDELO15ERuRP05RKP2jqegVbIezcurHBxqpCfBtwpcr+agjljW/s2hkPgW/cplvLoPCsg0oDFrWm
u41SjckAavOlY544DxaayxWl0sdeturudBaybjGGOD8vYnf9JGUZQznBWuNWcjkgCOSQ+fgnpOdl
kPPgWQlMWx1Xmb95RrfAHZIPjQmlZG9WEC14Lt4rUTm1Bi4YW4EQ4U6np2gP3kQ9GKIh3Ys7zu6M
fpezI968+Wl4px4RiPTnxPEhnNfPpDKwElILYXwwyJHTj7x1kHZlmTVI/OCuoUskVMgVspD2l8IF
b9NC7kJwY/hmWHgbtq3xRiy4HGGbp8tF7W4fVTrTJjiIJF1KCRS2peumB5RCzY/7NN9b8o9Hdu4v
xRJFiVMHkOITmwJVEvlKoIpSw2W05WayRy/WovDyXGS0k94m0OYlBjiTZonKJN80Kf9RmsCQ7V4V
gdsIYJKLaJD+8fkP0ROuJNgqPZd+epTt1pJhOm6S+d8kCnMDQLrhSPeR6uuSFjPbQ5KX1T5cLa/X
XUHCFfkaSlnF4VNnqOPfPPIHwoXC8s+2pQWmonwOAeseg//HXkSxbuYIhs5f+0CL5k/EEypBxtp6
0LROXhNuRVCQ1Hl6O/SfnrVhQ/I+5wXcmYKWtwSX/lQrf6cFSXzb3JjXS01z+/mQF1xrBY2pZauJ
6dz00RgYmym4p+18+m7h/qqKi60hh8UuO7RLM8CCmHjMI2IOsZRV5OTkcZ3ndfH0FuJH27Nti0CU
gDR8nG2f8EFIbxQ3WDl/UYbgqu0MflPendXbIGraaHoEbtFyO4UlOm+YlwLe9ycIpXu6l0C4Jxda
InGYBBV0YRb92sbDG9hc0Gds7iuOJrJ1dTgJWqvH1TOLRw3cFz2rsNj69PcPRsIRrZOOPOyUL171
shNwEUOyetdVjAMoNfRF6Kvynl8Q8JtYFgbF5kZA90g3E4glHk5IqPuZz/rptrhYfxRIVGYcoeex
M6d+ylqnbFlgSQMDC0Glt75dSLAf2MCEvrTGb/G4bVKGESyVsn2IJir0kQRQe9n00aPoxKWas5gx
uVEcKWYSYhym/YPromWo/wnZvqDMDnCgU+jCOTYJZ7UyvuqIYrXzyv9hDGWDqzr621cn1Lvuoqm2
5lG5AJIhixorAJA6zChrdAEwGGSN7SfQyjNe3EfiUm8wwBZ3iFXhlqeOnxQfAbDXkaiH5B49+iM5
nyjDs6ScxygsfjDHd8Htb6qKfr6rAyaEMMKu6mAU57d1y1KRfoejRzY3qCztavWIGE0JYQLpjwmE
HIm3IIvNzTVvzMq4l8DI+53JZgZmw9kHS53qcd9tmNq+HiyEiuAmjoP1kpwLPnobogyo82veJKCv
9EE7OZAmZlc8H3VoXMGPYeAwwS7pyjquKgqSJ/3CQgoQYyezKWHJ/2Fwf8rbObFlCpUC8GO/oCkn
C6YLcgUl6G7OKhZyS83B6Y2/nRES0YJtz+KLYXUGG/2VGeL72RIzyeBRj+WNvTUvF+W69Xh9IYW4
tNuldNJW+llTUcCM0NDNBLo2m+T1IJetGX8EAGkBIee+q77h+/9CU4THwRfldSblhkCePEc9udzj
L9YyjcfNjy+6oqHJXcVqyy7IW/XAJ/awuKkuwda6iRxoq53V8ikpPIwV4QR7x6gzE5wkl4huMyr2
v4XP+ajGSORXDlx5MoRhPaHqUYdXAmaZ8MQte2pZYYphQaQ4zDg3hEHGLoutC8jlLgdC64vJp65T
sz7rArIo2cpb1NjheYf6UzYz8PXmp7yFi7ENWhtmpehy9j9b9vR9YTvr8vAsP/GdaN7M9F8pkbXU
jy3yB96IkJF9fZRbFarOJ2etupfwt54A789uWGzyfSM+GefD/50XxYrBVJ3qkrAORmIQb2/u4L4L
Bke9sp8UJL3iOZUS96Vh9PAWOgLf6a8fhnTkkxo9Gli+/GPNH+Toyxv6HYEgDTbURvpsdUmY9dHg
vMNQHWbqNwhSA1stuZPUkfF9N93bZD8ps2qNLRdgdY3QzDHKC9wUnV/rqB0XTjI5jCbGA0GkET7+
0vKRN8TRDJ3u2L9Ysc+o8Rv86mK0TEvaLuVqDNSIn9ufGrQN9cG0xjYKL++AyVjWvNrg0Js5v8zD
g10P7pUDV/tvBuRlyWaRB1DL/VTPWVi2JwRSMDH50sO+IU7cELh09k6gThZKy43j1YR2ijiy/NuF
raco8QnG0Q8ovgwprNE2Y/w0Fy+1Ew+pAo6rx2yTxEe10X8ppjzWT3kVhJUyawE6rkDTMW7Uzvvy
AkQ9uuWf27VFzl4ioWLaIcoZFAt7KiO/TCDoU7WzjFJXYvUMDlaW8j3WOpPnQtcPhvFA0qEt+Ifa
cpOeWirFGKrymf6owrXmGGvp1NTyH+YjibtcHiP/vZE1oMQJF/5gxSzROgPWmZcXwUGD5TMJavgY
V6Feo/9nheeEkB4MMbO7+ibEiUEv8t4yPa88PU67g8oCyN0t1JkGos+QJwUOdQriYzOmjzocSeKI
E1hk+1ZBoR6PDjjtHqqVmN62nwOd+sqNc3K4A+rzre0OEYiJ8Gg5nrdBrikypdsj/uZlqypjF2nS
BrJ68Oune99omI+p5M0pLktsepkkj/NCM2DVXVwhpivi4VSX64MULdgTSM9Nv4jjtneykyDbQTc1
P7+7JdC/uXw6BN7HkGyMRnV4ggPBI98/6eDMFqkeiSf/Vb8F9nOGHLlcT1j2KJ58KjGS/4+WzqOC
j7tO5QZfgo9H5Mt2gsLHXxlqPu/Fdldx/TcLtk7ol+MJ3JRITmmQz6pfFSTfKLPWKrxe5p3YYoJv
9ZrmfJ5RKcX8gtVnu5mScUhSqSNaZeZj1XkTASvdTETXSVaEFTqPyZu1IEDHWRHihXn2qgVg+i4t
KLepI4wQk15gy4cBgXAxARfPHgyG0lgbLVPyw5eXmPaZBzhBDzFBdbtRhYuUpO96doYe9nWvBTYI
5ppos5eY/5/149mrD7ekGQiLZBoT2KSAr5vlV4H7f3AeqBrfZmniCeWRgXFbQnDdGzGaRWZX45dL
I+LRH3SA/59cXtgz2+pvdptZ1B7Cdq+ZdKHUVVzT0n8XZAgh42WJnWlR6VLulcTkyEyeefiKnPX6
Zm/c/2uSdkVO+AAoZberA4qKGpInNBXHodQr+2vOT/1WR6edK8dWhy05aVLVYE6UK85em3jscyZO
Knu842XqI8ID2kcNAhD1rF0MAqnfqZXr8bW/fB/ZogW9QyS9ghq5xMbxxxbrVtrPMqL6vHYfuJ+0
FKHCBEE2M91NC1gUxeaUheqkXSqH6Jhsv+CUlPNOkvZV2CucKKjxcL39lhadv0pGAh89PEi4MGsG
G0qcyud/TR8aw4g12gYWko5JaNAs3eN/ubEyxxFSNPfBBPNjYkxde38tyVGZhJaWEzWaPCiR/ds1
2zwwrpiJMOkvk3KD3kl3D6BTYBr+q8KGb6C2MSNchxbj9+kHtrBB3mYosrinnICtKeTJGN9dNMS9
TcY3CyIe7DncmacHinFVp28fSDYNrIz2vSjNdsuU/TI4ccfSPE7ugw/UFG5EWE8BNcYiZ4B2MSJx
XDsAMQ7dPmX7grG/DGyeL5wcZt0St0MDwG/wQ37DzS4dOvN0339IDioYk03gkGCeJEraqSsX/oQA
J3SWfJh1qfiir9Dr3AhW0oIakdwNlf4+/ODQEoV7o+Q0FpnoWzS1Hs3MdjvkVlIr4RkNTc2eCxl8
XynkMzaR9A5E2MI/DygK+zVrDYKYA9jTM+aJCDA6MioCTZgbcN79vwn6yCuWq/qM3bIm/GG12MZC
3hTBN64ESps97mnURvRTGmW7kCNN5vYFkvOqdBl4rQHziqc9RdOVZTVlfS5mhu5RLEwR431x/oKd
47HUEyBORuQ5qwAm9bDpbHKiKCSQkXdn4ptR1cUZSqG8W68rVhAV2SRcyJ1le72mrvHj7MkFs3Bg
RAL4lTgGXAylbEyyq8C0/Zvput1ibU/hJbv4wWNE3ztYOIVEYs7j9jyyZda/ldmZNymGX2e8zPPH
k2k6ZLikh5IWtyfiiBLB25kjxRO9pdViOk1M+Lx0O7iihtE226/reTL9OBgLDWUGg5r2W+1TNJYw
xNFe7ImBpsc6e6rAN1C+8k1yebSWa9meu4iixKuioHJsp0pow7lE/nw69h+4XoJXEFpQo5ZjUZwS
aiPa1DvDoj50bhs0z78e6dfpWTC8EFFyJ16+aJdKJ9n5y5HP0yXbbvZj62YA4O6W0WB3x/sJj5tT
wlcn4FXvT5onxOPkruq6pCY3NLBYmSMHhwNJVbG0GuKPrIQPJ7G5qCH/PAhNFK1suI3bDnE1adKH
EmTbEPVSGwsZjVpQhvH9NYXoUaz2kI7fda/yPCvC5K8lPji02CCnf3EnHik9SVKupzYIDqlb/EIO
XgWBlvRjY9MM/IBW+xTds2cp0bMLNW6BgnwzjkQzJnA+PSXxzVnuH4qe60mTqbK/cxDQZ5VS0UQY
veGWkFEmxnnPp5kez9xXKPVwODOV0vja5m+FkmaHUYhUbxgihAvtcpuQVmBKorNSuvjGG3U6MRkZ
3D+DIHrOcbBG51foGF6NPITU4/PgErT6KTBVz8cU2z5uipVeGCtEGgYsxhVEZEkFAgxcG4hhzvm9
fGNzgJC5L0zSiVtVTdBxieSyFGSX9lLmgidJZ1A0lB+lsN2Rdwcvej303kvuBVpE59q7y3Og6Mff
Cl+9FVLBGYpv7frXP27+W7RX8zzWx4ZX45kl8PBi0MDr2jeMJ5ao7Orzg9pDkllb1fJYZWbQ2MM0
jC5sMgursqreP7+zo20ZT/veigrtVYSe33rL9aKjd3UQOGkapWfJ3YsL4tUMtmKpujxN0Rbo4Mmf
kAE0okrSMJ4wdYCIbFXxkq2+WJcAVVEBdFFj7qHqSprXUd2dgqnk4VI60B8+UBfgWUFHiM5k00dd
FIO5J8FTz4lAFoPb8zAWI/VsjIzZVLsEM4Iv3Dz2e2t13V3j0koxivVINlNjaWDPEhxUssIinYmq
TfBRDlbZ/HVmRPen1ZbdrdXOyVeWa3gS9Ui7XxOCUZvbzo72fAclMlhH6FixJbvZxpiLKXRnlmdm
tydIpEukxU406tMo3mE2qkOyCuIXMVEDkWYfr1iHIGHSyP9CEafw8yVFvJkbK9xBILxpn2ADcZni
z8JEeFxDnhY7ffv0d0RhDojuCyKQyWxH2vMMvf/LBqYxy01+wCYHrc0mCXmSuBE7qqgCBJmmwluk
moj1lVWnymMo5o47rbTrtvhXZrkS79xOszhP1XR4TjMPO0zI+WTuEXIkMZvR6s8Pvo9P7LOFB4Kn
uG1NKS8y7RH1i8xH1Mhi/pkN3ujlw+wBe1E8WWnblDRm0UEhvNyQjIt9d/75irZSRPC7hrKFpjLN
C10Nb8tclGimJZKRNkPF64Ju5G3XTMP+ojVWz0fomxtnpZYzTWUjK49kENroYPVUBPjQ+T8ShQi3
VMduBZ/+04+oa/+fi3ll3RfloTcze61Za9zmPUnc/AV0cERJ4z+KsQLN4FDXniRJpnoIwbVl426K
/fkN+cUlBmOdBeil9YFkDcs24dV1umUqBGyIFlpcrOHT0dVKIYn59G+OKbclWelsEU71fKZA+pjH
W/IY0vuxvtFQ+m3Qw7C8ZCAYYOczmwA2NEkINFi7aFEWXaASuUBjYj/Ua4XKxF09CL6UA1rueDO3
Ru4jiESAm2eeSFsrVTRIpdcQtYBJl+3MK5kQAyMFdMLVrJqIcjs46wSEzrsvJIEOx32jFeFBxE8q
1ge1isUefd1vgYmWDgobgBdrexbGCI+P2R/9HbCqfgVcXVGSfA21HejvUyh2adgrRZ4eKzG10dec
5CZUnhjudK9EtgOTde5/reZHai2GkA7fsWykA9pdgYU5XwnP+v6fJ7qnyURlb1Y9HFI3AncESfdE
Df5erNBZelrxgWqqVFX2puTWf7d6aKt4QuFtbzwXxRje5FDhtXjBNfGVo13XwMk5iEGrW1NejtvV
+S6LWaqVpLxif8krw/bZ7fku2vlBeuc7UNVmjglAykDQDLpdMJ0gfeFylfql4TCmPERyiLIx7imB
d0CzDO/DeCo+KX7o9is/ng+Unk1XRlywofR+emCMCvOzpRCiV0fa1r107XrE9JbWv2wM2KMHg4o9
XR25XlwvAroMfpt3rvZU2c7Mutvv3ABqYuv+cEqZhmvdhe3etGZWcqLDXc8805eAnOSOZkNipp0G
3ak5CE9PIqlXHC9X9KABMqAcAdOJmQ7PbKfGIqWtDgD7p85bYBOvoGuvQotqSHDKawu2kqfVZsoz
O+RfjpZGehxgq0fgbPcOCXY3fEdUoAHB5GuxRkXTZAvwWp1CEitNWL7o2HI9hzM+l4BdHZdusRBA
I/IWCOXIJjEDVsloUFwCHp9hzUodwbgaOem5F8n8CuGzvjPvG8JP6gju89hGYYHQ6F7m/F3+plHy
APCIu34as4HDHAG/ctWesEvJGVUiRguh0X2ewXCGVTJfjZbo1EoR8dwMO41fNcm2QfZO4eYxSzAt
/0k6IAyAn6wi8RhkHtBxonywqctWFNDJS/MHdsRKDzlWOedWSXmFubv98jRfDyHzDCzx2irnf5xv
B3H51CunxZ0PL4D0bxBd9Eyx4KdmHwcHyxTd+7cn82r7KbD2TLPif4mHtXxvsq0BylC+LEOjJhs4
u8hbWN8dJ2ZMXbASvAeA8ejA0yOc2JLjNLeTHOaCyWfAiRs+eR8AkEo1HyWEI+UEroruoor3HpZw
abQ4KYqnNp6ef8VyCTSs97z5n9wI7fE5YnIoKJZ76QPeCq2TeGloLjseDdgOjvpCVemxNi4WLulJ
Gq/At4VU1jmpayapgj1sE1T2qT5uvkqS9miiJB6TLpdvBqEoKqXYiozUDJX7svXNpa6wYIM9PxIN
seE6KBiNIGlbUR7QoS9MCzln24aygoTkvGWUE4jrdybqRJAGx+07nTnLit2XguDHNT7KPu1HXKpG
zW+cKV7jdHq/c4S4jv4kIUlAzDm+CflNTTnyjgWKnBPQfjw0zQbIuxQAfCkR/GBDF4LAECiI5OMI
GiaINDRc6qBNfgoJDRXIQOhPhvqS4Q++JhRIeYIHu5+LWdKMfJzVL9rjybpaLHLlZ2uPYDt5KII9
4YcAzVyYtpUlLjapZ0kMDyuHmpdplcX812EmTAfxY/StrMaAiAS1jMxDdDIY2z0+usg6uXJNaxA6
mup8SNYXgg+nFVyMjkFWFEVx7iudLgIj5Z7TLsr9Rpmszvy4cXUNhEw1BzBkgMbGRKxWvDWqooXQ
iswyY9Ho5hGxAYHC9viGmUEbblaDPcjJov4xE8GfFUC1Id9oxfgbalwBHQHn+vy5/Rp5Ro/mY+sB
JLjKUMYDIj1GGxg8J4Bdw4Ji5LJpSulh7dEmkNobY9J3NEwd0VS4pTyRqoB8ftytR9RQdw1RuPI1
O3hV+QNFeRWZyO31qyWLAmWuRBfaQmXEbFIj8rMi/2KEAAup/P7jEP1Z/CBRUO6OF0Rx3hafhtPa
QyfokmI7tYG1Re+HFH7Y9IYwv7ZN44WGqE7DQ0xvT3MDYtBM7vvmSgX45e1+NRMsPlt1NsbIa5ul
ojauowu1bASd2Pvs7JGvBnwm/qF6K6Jaw7v40U18vuStjwu+NFT6uEOs3Ik/VhsyiMxj60n+deER
4cdHjBuHyxVoM4p/tDUo/ITkP5TmB8BR+TI8nNib6O4ZYcBPSXBcj2c+Jucn4+YKiMcczn0qceFt
0RRCLDHPHgi8LaDjfgN2tyfd2T8PsCoX9MZd/A042BQSRe6EpGOQavdZWYe9O4wJV2JdWUXG1e1E
8Rrz+eXkk9dfEGn/CzaKO658CeJKxeM0CnM8r9S7kaAHPJtFKN9z3TAMRjSabavp4qXWfjJj80Pc
AyA33sD2yzyGOuGCT118gkq87T4iFtwfOs2/nE4Rl59dpePDWNjFlhiBiiH86pnjDyfanZaUWiOP
m90/UZth6SSJyqdOT5b+aUFLOqvUKLnBPDo8ssAsCYjUGaRlt17mNT9u+12BsXtP/rlVBnfGnk8B
0Tz2lp2ruE0fSvMdKz4B3kpdGt5KoXfGn8SFiTtlIbXK2Gukfj6a3Ip56xKxz3BFSzBZ0WcrWGX0
+7iiajtSTCRt70SX+vN9VsTWRqK6QmZs1QqtzrQT+jlyYSCYLRQd8DpGDnSisZ2vve2m0Gzq6/xq
SdFokHqwWyIKMvZKTM3HnIqIoPCUxNA5T9VRUE9yWXO1qyCqHL934s+sATngFUgstGJBM0abw+2t
0bY/nl1uybyKGGUXehkOItObKzdP+Ax0CRtWJPgksVsdvFsdAjuqq9AlVgy32zfENvfVsnL/F5xb
PzmURPucyLipea7xO4SzZDJbBTBrahVkepUJVWLLWpWjBka/y9Nw7lXxwRSM4P+z8i+DdCPYhFkF
NqLZLZSO1LSj+ZPHfD5Sg+pBwIBGhTGAqrczwb5Gp4laELQb1KproydivplB3JCNRNYHsFw6m9vt
Z2T+o/QkK5fLq+OQexL/f7Ei8eWu7AKPHwK6lYXPyJvq5S0GuqMylG5q1rv/3tNw7PAgjkqJE8lq
n19znjFbnk+ucgyVFxEkhWssar67/FnchsbVRTMPiZJsPXTfgF8pI0KwjAx10EMQOgCgKxxSmYwC
Hvr5uWn9t2/fLp7ZegOQEt9rtknctSFz8uM5RWlf+kGk25bncmL9aAvxjAAnJZM1aI7RnM9sIA6n
wPlwQgaQ8s1ryrUYbOl4m3SNqqDfTs0nV6bcpXA4J7Tk80HPs4ARpjS0DnxlWHyTYEJ9dTco2Zc1
tG+LSa7riaROSuwpmFDayHPDzWFR9MN7gH5U+xjHolYLmvc0XebVfAuMw96dFevLCpYOMABHyFMt
pSOMH4Q6xv2cVFfMgfRnMZSqRDhkCfERPr43RFz3jTX/9KHkbM5xpI4mZQC75jhrG5BvXnSf0Tba
LzoGWyS1VNs0bbhtK4XnrIi1uDp2SXouCIjnpCppEAVyE58ILECMR2L53zHiW2c5EIaN4IEiVakH
6r/xMMmcIMii7Al2VdwfOzN9SGDMsS9xLkYHJSd3r6AjaJef4rtzsIstxS1bjJUh3tpJbcYVrfSD
iCZ5z2ZUo8YdVBCPXAHCxnMa6/yu4evA/tJd61HFm80jW3xV+O+riebZ3+eg3DtyztNjN35pib/c
Lw57r6Vg80UEc7qvVY6RJ4gCCGH3ukRSbMRYVjBpPabA1ZH7K7+38f/wmds+/YD7sS5xH3IJ3BqC
3N17TFulWm11gky89HIJpYKBaT9hlbZp2PmNKHDXExB5oW1OeVZRWYA558sUme6fi+Q5/JDndjlO
p9zz8xjwW0vih6kLd9IMtg43wY469SdS7OCYhYri644RSLkMmVLjEy4ySP/Td/y1ZguRWmHw4A58
DeJh32/6KzvQXdIQNXBGLJn7gU+8+h/U8EzaJwGby4lBJkAayubcBBNvjs3MYs5pox0q8d227Isj
ZPZ0cp5L54Cwcae2TnZKkaWkNN10N/EyqjKU/2780WtCcs+SUqlGrlOkM5SC2bvWXPr69v3hTBzu
G82Tb+hEPVJIgwN9vzug4BIk9d0hg2RRUjWyVKIvPT09pedSFZI4rcw4+rQO8XQTSHJ9xeIfHxgN
BROsHpGsIo6O3E5r9uQMkrg+Mbr+P/014eA0cJv81hg37k+5UgfK9P3wlI5Y+JxV97n85KkOeZ/j
2pqVaqyQyhcmQB2rrAnXAD3Nu6QQOfM1UP3CY82ldHDhCqd6UwV9u9bJ4U5n/CCOHHl5n5xdFA2F
zb0N8ZGq5/JcBO5EiBl2Lh+TB2fMgV8hy6U0H482LsWy+oJOl7gUuibyOiyJnKf15byR2IBgKJkN
pGSPIZav3Z9W/mXJtEfVwJ8sEDE6EBueXHmeqIjQZ5cBOGBhoPzC5b6N0XsCy3ghsqtDuuQ7ca49
LEF8iUOwq8bU43Pd/jO4QbrOBp0LGRaoSvEkl+w7zhk6bTR7cx6XP28pRc1qWqtF56c6fdmoaZ0y
Q0ckoIKUEoy82wkTargTxn2mLaMvPiuUMTMTvBTTw0mfdPGXn3qfs3dcrTomrNOn9r6LwjbiRxtm
46M4vY3wHf6Lyj5E93sQnieX70mpy/zCabu9j/ajagcgL87rBF8hrMEFEn1OnjC0TXz4bjGXYZwt
GphjS/i/Y/IZ5kwl6ThgMd9L7Tz5du0u6KYF1WnIJ0e+0bUiD0i3a/RaN0pK7XvSqipCkr9Mj6MB
hYe7J9bQFPCZYs+jLmfam76sW1kuJh+n4oDN1Zn3HJujlGIK5INo9aCKnjR4/wJNHxxRwOAzxZZG
XcT//dFkutXHm9fFINsL2jniSLRavJM6WyVAMTFhrbIqLllM25Hqjfo1PE+gmR5wnrMMwy7V8w3X
D0n7Uz3y0G1eq0N6XzMBG3BB6YtIwvzuvMlW8pmPe6zDGaKlhh+/tfkIKyV9p8kYn4reBSfSqYZX
h4k67WB8rO7ouR7Ia6ReR/pQT5SLFpBm2P6RrOB31ErCOPIWtfK5cN3yRTKZQ+X/UPD3uQ0h9xaV
BZW3XhenZOrQRVXZ50LUt0eqNTnrwZ+eL5rf3/ue1Ph4Zpww3sBuSQr3ycjmk4qKOjcKn+HPP5VL
P3maHXEQtzpAtxQIOqkTGMfSCVw4SxFpImRGCBUikT84slcQmsYBOjvunC2pXrebWTrZZEG8ZfNz
k/MshW+7xdZCviieRwLzN4f0gkRD41wFMJCWNzr1bUtGLXGIe3n7Rgy4SHLOSGWVe7ESuvGkZ0vT
KNg72qP8503Np6A+onHMFCiesLFeWTWtxI1jE9nO9d2pW3QQFjvhUjf7Kf5PSyPDq9Hbt/rMrviM
zUWtjN/AQMqTJcOwU0OGt1CmaNOYhSA80Sz9RBWuhaEERkUTJFGpQVmGrh4P0VIGhOiSn9T0Bk4O
5ibvycb8GW8L9z5hHe/A98KxAGTMspm8+V9+YRHaxANR8bQLinw/uU9MhPZKKzbNjhkTZ4ALucS9
ncNkW0/4F3Z3L2aB5wQMSpUhFYA0lgsxr4lFE9/ZpM4//D75Qhu7gDyG01wSjXwiel1LaWerl22T
xuO33dtxjNVrvSm5b7xNHqcc6fLcsAJovcQXg112TM1KOJApjUQQ5cfGgtZidHvHrpX34JCBGZEA
AP8sP2AsRTfVilPQwKX3T7NO340E2ozXYjtl87a/KIExOCI/ByYwFxT9jgPQWX+oodzEGM7fV3vw
LopC3QSZkwklCLUx1C3AN5x16TBnXhI1KTDZcGe36SciZxVkBjELKXVze5PAv5lMKBXIHZKDJNLk
NF8wCHYWnwWCmcUp3azZtwXt2AY++rNpVVxE7/cxiFtfwZqW9frIqYwFU1BZJfcfcVFOQ3GN+YDC
BDx1HO9VcBdXVewmsDXyGeMqoB3Bh9uPB4sfE/SIw9t7+qgD7Le3EqaCxnt0MowuIDy78TB5pRCL
R1Mq65y4PwOLU7E6uLUKuPuPXplToblBZRwQ5GojObcOtZXpPUc+MyVmDaFTATvwAKWKBFfOPJi+
JAh3i5yMHk232DREE5OtF9548bzNlKt3S+o/t45yMW04eQcaQrdmmFSwO9Qm8UAJGHK8ZTScohjE
tFFdzeFTM6cvNewEAVJJQ/hgUpljibqxGQ4FZpQZkQ/LCHmSrOdth1OKvWBvRfuckUCdtTiQdWBr
3poY9uhPviczk3K8bE6rYK1Bp7ZL1ukXtMoxUGFSLpKF+PHpEcgClpKpL5ccdXM2C8kgYP3O0D85
gxgWiIfTljiqT3cWAtDSt8LTGsafKQYdSxHYvYOdHaACvflbhHEacBte6WHmmyldmDthFfcw2Tl+
y743wwgct1BAkQS6fCzJV9Dku5QKlqpoCwlfmhFHgCnRSFXcatIez7LZxYc2udGX+DLDNWm/iDU1
4i3r+cQY1PqQBR2HWZZ7eF25SY/LcJpnLE/BY8Lu3H1hw5bWvGyzjj15RSs7EF13t+6rf8nbSf83
avRPFkyZjlmq+cGdC4M0pMcI6SxisiRFdxb5Q4aaTvOcrePdxFfdWDH+xZIuZAkk4vAlkF/Odhwn
lR7oF2de9Uwf76de4AJi59JePl/qxlloQTF6hGTh8dXWjHWKe10Zw+G2wm3JP+97NumfYB9htSmf
NmQiUpmfurI+6qabtqgqs3c6a8xDTaNMb0jD4HbiEA6Ag1FbPs88RF4fmMQWuZcxkgDcXsWSR4fd
NOcrVXcvfhmYOXvzrFS5THNeacZxFdcXvLcfGcOZs5MNO4mefKpXPgmUIBPBAnVzyTya7L4Olbdi
jjUnP27+iXHJpt099G1XfVpnKhG+aPm+ue7b/usZmAIM9JNZT6VcutATwshsFsFuHp/EA7srF3y6
Iv4QmITtdD1kjXyYvnO5vjnqe7JBaORiWvOlUCh4Yy43ioo+5bFyFq7gB2blvc7I1xjkIJQIRGLE
1gr4hwFzKgcTXlggouqkVbCjNsy5157SMg4vE2s6rde5RRZxyr7zxjRETqMrq+LpNZtfW7gMlVrN
1Y8t9NCZBF7Ezu+iA6z7BL6n7hNgq9/DS175veMiNjYnUzePQOt+ERGIDL05ELaUiLuuII8wNSHI
YoRUAcHr2oBZjH8a2gaadiLN3yt6W+nYawfSnaYorU377/XOZo7btXDFev62/AGZbf8vEpa5ufmg
LWMTkCZ5Sdt3F4qlsXHlqVpr7gtmrvh7pfRe08WnemQhvP8X1OMY1qShDS+bzs9HYMy+V1itoGZQ
FjGJIk3gE0FKbF27Lu7HtVV4b7tGGXtSzZYw9Y+rE6g+bqBTJJEOpmQKH2/HCtYILminFm/AyFm+
gWDIaj7fS2C1xmXWAEfqeuEEgs2kthL7V4ES1AcZCoUfCPEKDKvn9UzhBeJNK95AZ1NQ+rl08Jc7
eiM+Gojdg+8p3KjlYQ6xHtcvgnHXbaBLZpJZWDmlQswiQly2zTuu0NLM52n8wBAc7nukbvqjeMbB
Gzv/n5XEIDpQFet8NvppNy11YA1fK0/TdjZkXk/+SGFJkg+P9htZY6/f7Z47d9w9Y+1dAOrs0zLP
YVB1VB0U60c+9pr/E41K0hdZsb88t2MHZW8FgLwKMr0kjwZdziG8pwRnmzp+c1rIrt8m1XKLR/sT
4tH5jXkCsWUt0YTKDsHCnYcAsaL0YScDtWsl9nAUkODob+OxM1Aq5+50CRVpNlaDKbVBNHM/37Ch
4SA9h7Wfbjtaep6nsXSwwak3GrWGDmkqQpUuoPxfOiOmEfPVZvlmsF0LBIArFfWYuyYSaI00xdQV
ZZynvtkES/CFN/0/Wj+zKGvpWpAzV3rRtPa3UN1ZjJ1V54aRYXYSaauo6wkWxY2qUm4YWuTVViYN
BLoocOvxxzbw5yX3MPMLh9xkGJCIBDPsilAaD9UZFSRekeZHTVUMNlWwsptcwxHY/V2s6f9PikVX
0AU4YzPHAzq1KiIV0JPEd9XKEnmfrbcZ0uUYNaar4zm9OqbL7czR+M4wS0td7ZyOA7PzPsreYznW
oRU8G0+JOBj+Ou8q60ZY0oDLUzxA82szdj3gOFg5IA6d3mpER8a2OxDq+6x+vr8wQtQqZMSz1bUN
GTs4qINgde86dHsj2ocxRCyyKX7g+q7KrJQwhyhRH9L59jkmK6Ri+bda3QJKRVJpE5BBOrmUc8x1
NpHgWK5VlKowD4i3T9kuvY9/4awJUe2wNDMzljgd9n0r2t17GUgrKv8MH39MZrZ+TiyB7ysc5cxd
Of7o2AIvgv8HyLoKrscu/DwWdxBWIHU6awK+HRH+g4Q1KkLAtG85cEW2QQL/VRTuFtEVICcuEbSc
ErOekeC3ANHJJrz9G9Zshwvziq+8S0oOxf5NZ2M/dwTbZOYJ4XfrwH0A6POQzJK7LFB6+CbqKN/3
yxiQ+5zKb32BeTpPtt5gQTYyg5/FjrA/rD/LTSs6e/uRggXaaQEM/irk1CYZxwnEaNQSM1lWtEV9
OI64R77geqdkWCMocCcTU7VZ4f8UrFOofFOknIRmBGCdsqrEn5GSV7oVaIKmzIlZHDGSGZ/fYKmq
F/A8j6Dw7LbMoKnCtF+U7MxI2OhsRJ84bBB3qNwLK1/vdDE5cRMaRcTnEZUOEwH+KAlnvXf/uvaQ
3R9MOPQGmxjAq3B7QyjeBqpGGW+sqg0lEjT2RH+7TXv94uhQsTECmwXSd88uHnV77PayUFoevuJ4
Ee9fxqpiV1BFU0mo3XrlaJlQo5bo2r/ag4V2U9jSAtWcQHNtOHhxON8K1EukIe9ljDRZeUcjP7vy
g/B5bEdM/lP/n+Vgm0YQvRnL2X6iX60rzJw/cLiQk3mteGmvA9ecr6/U9q5IlSO5j/gGGlnniGVm
aegTvho5cymqx/HvSau852lqy88fdUOgIjfjcoAjIjS8Bc+RT2rlkeRFh3zIc1ibKhGR980WsYOW
A6gS9eI3pa6fBHhdKivYf9xQZTPZbW8gMxcHGKY8soR19RvxNkp1Jn2scF0n/+BFQMCy5z1wavrQ
OkPbdEeEZ+uYYVuCCsrWwaecilRPeRLppaoEiZErZ3M0RtRbEMHH24yAw8e0KcgQKW1M0Ogi9xJc
NQrcM6J3ckxtSzqrklH8RnWKO+LeiOq+aQ8UjvUeWz6wlngAKV9j0Gnw4oMr1Oc13ld8T2D/L3BE
oyEuKKUKe+oLbE9WLvzjw4tfamngyIz/E6N+2t9s9kjNqP+g5szlqze2j3af4VOy/d4Y2jAjFU1A
qqAd9xokJ0gUO/kFaWjEXj1YQpCt/g2fOLc/NLP7SOlOGyysK26E/SFJAiG/2WULlgh1ARmn5aCy
b428we8/4j1eg380721JVRKlcfCLjx6qVQKkUCBQs90kK3zl84+2uSQS23fGmM4U1QTXGiQDQl9y
SI24jZgwahZvi3ebB+fYeeVUmQ6FSldGatLK4fSTWoX4Owyeb9WDiFjGXUZw+SFVjmaKjA7y8PnJ
q6uK1B0/aOX3vwU+GAFyeuJlp8p253FLTfZyusZvEzA3hVSs8yEIJxGNgRAsq3Cba5/Wnar7maX4
KxNJ9J4OIDSfWjktBQ3Zw9DiuR0hF/ui0pX89gumgPQt4uga7E5WnON0Km/ZTCye2GjdEFOgoDPc
7SDOX1AE8Ba/2VlroMsdfcThcVEnIyk3i9vJCDUeyfYFlVq8Ih3pUSogYQTD0Ey+j39pmfEnfvYY
IbjIYrBZ4DZQ8WxVkvryt75G04X443IT8gVtL3BFojCYzyGyF85RMw6LLAw0m/WqTQqJsb4f+FvR
s0sQC0175UYyKIjuGnetmorsJbGZzzc+YMEfTQRjEBDn5x9toFnBWDEdU0ChW6BXNbJPtbLHWKcg
N8EtcTtm6xEjHnKybjdEY7yUAR9KKFIKQYvENW25jOgXgd+4g2wwWRaihKOJhoT8abGvNBdfvO/I
MdkNfrY/qTRn7mJkjJry6gu0zXziNxKGORdWBNIR3BMgSlDb/IyPtc9jfJbcHn4Sk7780NtIjgsU
TgGP13X/0sdIpjHtHBAzjVLqT0CXs0a6C4HPOzylVuU8BxBGLs/vpOItexKiP6wAaqrxkEYC2lpO
RYCLBQ93tZInFya/0S0xU/JOsVaDxy9Q3BxWkqHNBIm3tq/fa9X/ol8RWiLqm23AT2syfQmmaRVQ
zcNCWZzpDsf0rDOo5c4jp+6Z5Ji6AfrUNuO+B1tYuJzCVYgtX+zO9uYnnEr9gqp1dO38mfiwc0nX
b0pRKTKm24O+ZuVX/qoY2ZimItfy4n5qUfNDq2rnusBwuCIg9mzyUuhwImSZyDQb74a66n5Tmv9H
dyFEW75aQ/8PUe6ySVwjEmJjBKO1QmpQBNg/DK3ijx+OywZzyzHH/D29PGFvaHOvQCjC0Wiembi9
QV4D8SDNdB9hFJmG5+yIk9XzUfA8h+vGVYHkRCxqxFWbXLM6WlaU26ATa5DNCCxxz8+xwF0YEJHm
VqN6bVt+7R7FTFkbTddz6C9sOZU3XpnmxflGpnIRiT1tY0wrCduM+WZ2BFACZ77RuEIUO02rUcZp
LM8P+w/6WPFmeOa7Wrf6jBJidmyB18V5lGiB3LLrJSwHeZ87FgAq7dlhNj/c4pPSZF6B1/RPY43W
rFbSjw9g7U7uzW7g/QVAxn8BJqPTEhsn72CFqGPB8DL0QF8kWnLASkcKWNzweIbW8gABkEKTxlCN
GtHTSmrtYWctq3zzRhhFoV0P4zE4a6kUvHfLccMDeLoeARzU9bpn8IqCezl8ocVJZNLDABsEUFWt
Tz2Rlni9eNmbdWQ5Oh9mLNpul/sRJHNbz62liau9cnXTD0YGsnTgFiFl2nIyQQ/d5kmY+6FtYNR8
fdzg5XYPpAXIYoSHcCM5UQsE5HXMys3o7k1vTyuNXZkxdWEcmxGODDPWwsCOn6S7PHJ1YqJvTYFR
n39lQ4j9T0nIpnmXr18yadhdO/FWtYg8Up+8CXeAVHPzeXzBNGHpVCYAtqBzzMbaOJH646MEw3LX
ZBJUJtVGmwpheqN7ivEjNQvcSMnvrPEhXWva22XOPbtbFX/4Tv8qGdHTdRp1bOnv2CaquBpUK9rc
NHmHaHFawR6BlLYGpxEEU3I7HhWlLgMyji81SYaw6syTheZvQEvFLjtv/JNPbeMMKrsdV+VXZoKH
x1/DBc1/X1G8TkfMX3FzlQXNnezjqqFkhp8j+W5L72QlfOSCyHM6xN8PCnHsrA8cgsQERcuN5Mbc
xIVNEB/4oFxKScVohfCK+79ClD/IV8mOyassOYDdyOzWU5TlR922F8yMkHXbDPbAe1wQeXcpoZfA
k5v9atGOVt0KjqQid+1w1mYyHVKbYfnB9hwtOw0TfKbZce8wb/U24SYXoD5tFEE+ejB6b5Pp2Vp6
MMwrWUcXDwoQhV3GFFuhXxVDIXTd6tc37giYox5aoXoLg7JMieJ+ABcVUs7VyDX7Jy5kbqhdIg4M
Kbq+CETg4RjpmWkJePczK1ZrI/WhCx84W8LTh+4bNjimcE1Q2RN2ARiH7kxYxozVi9xOzVLIrcWl
/08crO9aFf5rBE5P1YGcXBXgGiSo13Il3li1oyMoIrJFzDlx9uaN+isRpMLUSgRTm7WbXNZsslC+
2APrYsUqmtgdPu5MDZuRGxZbDQSBKlJnfXw6+M5Me6BowXCTAynU5nWFiErz4le12KrNx4uj5IMe
FuvsQiybJwrSh9j/wXee4lIGTHKK6+96GEO//eMDiKwtxxIWKIwewS61Byqb93U2W2na7ebrOxIa
kmy6gcM6P1mdwSMora800OvPcomjoGn3Avvje8ZsaakNcq0amPfBiVXtWZ0yRDeQJP2HoevzHDSw
86amzatTmq7/g50H0f5F5zRyxOAepwW/Cj1M63FDt0+3U6BPNVt+ofD3chHk0wbdOI+YOkGDzcy/
tU9P8FXv4d1VDUZiJo4m4X3cO62MJBh9GsH3ahh++YY7pUDG+keDxo/dWRfiK2tEQxIdb9tB6OYA
8gDgT7NVT3Alrk2HpX5B0HbxRjStrBRAjshuWSi1Tn7E8FrSfszT8aYfBO0+3RBMPjU7iJaWb/k0
z0PlVks4X3jC7wnS2iK/nThzofguz0wCp/N5sUEfEhE+HrpuSe4pxSnYtog/KvJZEWVBz02dSedQ
cP6xNu4NtSNHCITR2VV8wL3yevqh/l1fHGBp0Sv8cpypuQChDDaagDPmNIVxwx8UKQuX94GZMo5Y
IXRfUyUMsu4e/QA1iDsBfLwylvt4R4QogkmlO0gAeHuLWeChk0/mBfpOIUedJYpebqYvkQVaZAOe
91t02zblNseXn4G6gWAifEXfsJKdfgeacaSorcdFG8Ww2HuCRHZowdG4Mr2I4t5H2sBQmMNZrKov
04bRYScweXSYEihUiD8bwlx1UHI3VjXVd0MXBoAu0vcNJ9hp3nV8Zr4hjO1k1X4vSxU0aZPjI8Gp
CRAmsWiWloTQQDsSGZ91UO8/hIOlc+0Jq/G9ISZL1mhpl5xpfeIggU67JLdBvPiW+vynZognYtUq
ugA804AKmq056q4li7ozvlfT10varrL+mhu6jXnPtLvhxpTNzzLET9kXwHof+4XaauVdAQLfDPXS
RqdMy3asc3RaA72+Xy99XyMKAd9LZUKOD4heIEX/+s3+qh+VBusUxnLnhqB/2UsYSE7117rEENDg
eDV7XoDKMiwnXtloxlvdC3LZrahMUWgQP7EcSYDPhChlg4evK80Mgnk+L70U+SaD3FmnQyqnT3yD
OJSLCSaK+rqcV7OMbM6+TN7D3mEdcNl0r/LKXgzNVSCbXgxXMLCZF3SgW83owbnWPTTNQfPlj5Lq
tUn90au2DbCStp8RGTzsgFNumYvr2Qefd27owffEbRdhN7xn0f0ev+XA6SHerXFOihMayZEDkzvE
6j/HusZsI1dWDzIBnqVHOb1av+BFeJjZd6RXAgK7xBDGyLcjpZEg/gYn788UnzMEtOEb5szUGyVh
P3DyzVVM7YV87l5AXs5/joGCzy4FUSZvE7F9oB5xRBdbyZggL2aomBH4PnE5iIqYCHUGlPlYmBbj
h31bmLhHEssy54FHu3wviWak7cDfOrTqzLkjdP66h+WAsLTMeKftjr0hMS8NCYqfNECAOxnYzMp2
+iPrxR5eKL6etRyeSJWSMU1ABWV2mbsoFTelK7a7JILetVe7Op09xT3bRFPsPH/MP7vCxpEXMwJ9
qG8s+Xba3XaOVDjRu5aai487HgIW2iqPNRvk6i3SuU/C/AN3ibx55HchB4MdnbZpIVFiUTQ8HW6O
EMnOb8Lex68wx2+bOSZR9yfl2V/nbgSuW8QUvvpwuuKV9UqJWV1v9/BUHI1aNoKp0TyZpCh7T5sh
xkbyvQe6nX1FnuVOUCKHPJLucytJf8Gbt3JOGm9JCzkdgnqC67mdD8DdtR00Ty/VdHuarY1JRTWZ
yL4kxcuQ9rM6Trs+jA/Z5baXebAoF9SOUHJQmKpNkZLMk1DH3Is+d0tIAsxJ0hP8V7PPRG/s7TRb
O2DKKYBSnRqka+F3YjZtKK8HMvgo4o0yBDkipF2/NRrScomI/164yxxjSjeBJkH9uEAlnXyCMSXy
U03SYLhyTadSMKDvQqCX7Y7R4DP0p5OSon1qIUHZNqk9KXDrjToES60wjoke1PggJYDXK8DdtmgY
kFX4e8OraQESzfOPQaBrxYRmzVihFlo3iir5FUaJy6yPTO4M7lLByiEvfs+vSpYfF1nnZZJ/ezea
hDZU52Y3xBqZ55hMhvgIVn2drSnUd4S5Jj2YHNQPhhlr+UtsmsyFP5R7Hf7Unk46GLv3AQLc0DvT
+yCkCTND7Olt9EG2zxodmBN7CvC4Z6kF+RQYjv+TAqo6bNec7mDQFhitaUFsq6hKq+EifwHecJ7I
nsKbd9VAy/ljuqTlGtNxBRYPOniSgE6FyeHAxC8CERusmgf0IVN7QjMAv0ZeJCjdyxYOkLqcFFCk
EHHp3tTr91Tr+jl4K2WFwh8C/nYbTNtrctfeqk2+lT3QE2anvPp3dTu19SZeM1SclIgnOzVPBQxL
7oXuGFhKlqH4XTLjfRQJ9BA6iL+3BB2dolnJt4VlFxyVkJd7/upPADKcE/O0/ASDgE6Et2ivDmNt
nshIy0IcbKkEV19KR9mEYkEI7IMHkvLelJnPBfLmhDKUNjmXpYL8gRCxxtsw4DkaAiPdKR2u8x3m
utIWuMExIBS5NvQLUAtG192d+EB2IB2w8S2bxWIpy42FK0E6IKISlPkmteGzz/Jd0XvV28O3VI7x
Xbnmyq5/HQ0a2+iL7nCrdYYUcVuJXFsrytjFqOd66pqUc06YgLITh9p3ndu0RUpILgWpBiBr1gQJ
mXlJmHgV/7CYLVOPmoDu7pU/yeMRWIVH3k42u8EqLOHq85XQeGIf2GN4pM0m8Tz3F2mYYSRKQD9O
HGxG8lqWtSH7sLRdrofGvyr3f/mpNNfhb9mRpdFHKBflxfEYm68kFgL9hWjWdTcgwMe/1CXZVhV1
n1rme7sJbxNQI+AgheItVHtBIATZO/pBXGIqVnmkqPvrbl6Pr87JWf5KjHAyIuysCjd2q/rQiWnc
iYiCVJsIbq4B9YBmdCLqnZ7ZAgB7YStgY9DYAeF3L05pCrn8sFQ0XL4XGy5UJPVV6t754N6ZwnEI
hBNQ4SE2aomtFMCYn4eVeX/JUBU+VCrPHBR+22d3soKJuVVJDCiN2EEata7fpGcLv8cJlrgA9HoZ
QKs6mdct5UCKDeM2rRSa50uioF8LmLqal1JkSGTohED82TJrnkLNO0FdewqFmUTF1qfeX73/PgkF
DaISA7QCmOkDuRcCsiMBYJ1KQ7hapYoleZXrhszgtR78ti7a0lgQ/t5nuX3H3YHqHRPGmrhbXsN9
kTGl31gIczWXlfiklualJBSx29zoVQhaypLqYmaXOMjAq4TzmgLLGsvqOj6R+F0ZDWO9iaB/LmGG
gQdB7e9x7mG/7Emkzb+PbGmhyLVb9sQQmU6vOg++7V/ui2VYP2ZVzpvCkyQxcLBC1OUbOvIEQdcQ
Xoa++DHelnLlWtqLqqI3c8c9G1rQYH/mV3du/w1zKNW6nh9dQ9FXo9x0ca2zzpm6xUXsVfHXTeGA
+iFMUGNrnRj4ByrF1vU6n/FIknWKQdUF6OKhxLPyuauHnz3iErILvgwWqP1GNaoY+nVxwd4W3Py+
KzkoJeQYwg3w77CGi3WPJhEjXPC4uJc+oBGcFHz1L49gXccWZzkOgO4jUHxqMM7np6wQsFKDcYUt
4ST8wT9JepiJhuuZdDdNSo7MLeVRkaIEKR1qxaoZR+vYneUpYKoNHso/1BTxjXuhIJq7G5ZK/D48
DyhghdbkYsYg43N4uPci2cLPUEy+/cr0iCbxoJXLTPi3Au4aCClIco/tepQzGUk170WC+iBx4EHF
5s+eV3qeZ5Eb+wGp1ZQG68zQzC0Tyz0zseRzzuQhmVOqVtpyefrtCb8Qg3PM386W2unsE9AYM+Lm
h01XNtrbMfWR9FzNgP6ekonMKPwrkq4KDMDm3YynpsHV38iXt00DYGc9en0VfuIGpFpXawBdNfYn
gZZhxK0/t5PyGpe8lOkEOeYRhgMeB0gp5enzco0Bq8ffx7UUYNJ7BSdkQ7HzA9quEuwn3yVCXhxU
vmDNZwXXL6NVDcQXwLV2E9PduXtAkrvBe27Y6cwdMuY+RtLh9xT37wE7UEN7pyBNIDMZrGTc9QeD
xujqgrbXOwahjrbysK9v2mm6zS2s1yry2flRq4YBXScg9FnYoJEQTYP7otyuX6qZgWgh2XBptB+D
D/hGNgIBHvS5rtJJ3Iy5+tscwOaB9lbb0ir9PgNKPzLiBNVJySM0fqrVeudeY9gCoCF7eI5Qt+s6
beH+WDpIQXqYu7S/9/9XVFHAoIE8nrKWmwU3DF/iKTiQBokT6c36BL1QNBDz2Zsj2F2ZBxVuS2Zw
B5a9D0KRrcDKMSwGkd7tKxzMLIvGW6a4uRteWPPZC5ME+c3n5u1apqX9hAA/z0I9EStB6SC06qvk
YGRn3Sh3lb8l6qv9FqjiG5xe8J7OM9Sel+qRwPEgiFdwiGO5kqf2WnLGQnMzBXINnl/QB2tBUnCn
fopnn4A0d84opV1ba1tr+EFzLUUwhRo6AlF6z9MMjieNWYMxlLxPwcMD5aFtzAEYZuCUibR97WFe
TrCyNc4IaX1SRwrzsydQza4NP6TT8iqAQhTsJb941y3RCD9+2pGDr4vnOOqS43WC/RLTa3hRfnIR
j8FvAmxIoWgv7TCC9AzkLEn6VkrGos3JsLCbLtVirBn35xkGFayevvpFoX0HXNWZiy2GWVQOMkhi
KF8yBAkfshIyUwLxjkzFoluZEqEeURYIDQZ03Un7CiKle4NxbHyQwV1lDxLRsHsSCJzDmcASg7zj
G6w5Nndbla5VmXk93cvUzYzMtCinDV6FQXZfe3Gx7540oFBFHT/NJmu7tHr4VTYpEATw9r9WZG3Y
r5yTFtAhEuNS/iM1tZ5+siX4F5RDuAl1g4BLzUAGimpaRV9ew0FSETKDLlj4D1szHn6yznaiyLNq
osbk40hXAE91V7kOOjGapyDB6sria9tX+gYfZ+EXf05Y7QYPg0lGRiS/2JnrBtExtzs8AU9Ov+si
TGGyzAqjAUiXXnAvYfVs12l2fFGxHH8KiSEdpxCdr9/HHmolX+pjEX1kLJe+zNnKRUBYGgIIgsAP
fwxI+ItvAWrLd85TdYcwZpBfemYbhG8XBhYVFcpdGH9BqXUvF7z2L/1pyUY0mjsbPufsQ6r8CNim
y0/pxgbKmkTf3Yte/jL/eDZ1J/7O5So+LY6sIFLc451cmwr6pBCB5vmF/N+M8FKdytrjvbIphmx/
cvmuh/2yIKrw2cBLcygbjojNn7HnxshMgD3eo20lhKFvZbrPqGKaFo6R6mkDYgDbIcYCfJf8MF9a
ITp/Usc0pjdoYXbPvN11I9XUh5o2d/DK8Re3KOci2GT5jlB9dlxuG4mbPP9/1I5ibEF9KSiPey3h
qNRCBz2YN0z4E7vCsVmQ0ecnudmDEveuecubzuavgaFubp7jGkxSplwGj0oMTK76hyyPd5PBYW7P
QRV53iiRJBKl5VF1qJb5Ui7ClboiTC9lE+/4NuujaXJuNhlwSg0EqbU4nNp/hBpc2aN9HKmOYiNL
6TjYqM1C/foPZWX/6Fj+ROc4IbBv5/EBtMYyyRwZ7S+JYHp+pvpBs9R6WvO1O9vBZT2ed5yX3A4F
B5elh+G+FS1x7ncT2EzpnYlx1fmok2wr9Z4Qxp1sLFoYzo3bZYRPIUDK1yHXfBZ30GgODJ8GFu+h
ljXBE17f8qnV/3g1+aRFMJjailkT6678ytnFFqhB3J5d0aKAX8S5KGOwDSZKknATTO04xa8xGLfc
5TO0HsgtpVSS4LaaT26mHDM7OihMpR9dzXSoL4NyIZVHKQZ7vUIt4ZrsqOHQH7asGUCDomnrtCTh
4n53w2DOUwitM3WXW9Zba+OsuCXJeuAji7SJawWgjrQmfj7pbAelAegkuRxMRfgA9v2yBGIrYF33
XWWlPcjCgGv7vXmweel93RhDmAqQxUV8g65kHAirpBIFC20XtbgDkoqpnxvM7oVRLzp1HkW/RU4f
4ZC4nSF2rENrItBuXGFu5P8qKtL2cRYUoSJr44qSNTM0Phlc720yrc8zKKwcJjDo2hNkJHvl/ROt
o0XEc8wAEi+8Q564xlMxorjBJtljE6wY8U4NrYU/JicuaLQuHr8miznYLlB4WBX0wWHtbyXdeJZt
2ssesW0gpYl2keKGzCcc7Oi5aRfaUvlAWnPr/i2KKTgH+y62YmWmuLDRy7Cm8UVt2nCFN5zlH5jK
Z1HIz5E1lCqfFG1ap6zC6D91DrAlb9RSqa6jM/NHSm4swWnkrLFOQSZ5cqvpapHhVyUHAB/bQCCe
I7Eu3N+5UNVBvNzBhJI/fMuKuZCHk+6bIo6ah6VX75S2iay32v7ctW5gTuKB7SXbhGHqI402FcDW
IubG5sc20zQyrHU5FFVq2yFd0DSatI/U0R6HTqh/Aj4DwNR4wiKwievk9OxDCLmg24eX3js2D29/
SbG4Djl5c5mTnyE1qh6ylgtrHzddLogxrQmyzekIsWK6ousmw+uZbbRp+CV2yTsmAVyMpatl01Q4
6gGRK+wXYLltAeKCbnZpPH0g/2vB2yCTTbOcDST4o2LYmyfo482IrX/kSzi+Xobtn5JrP8xpFx+h
2Sn/GJIR+vDljeKc905ObUJk2Qf/lZeOlA6a4tyQxNFSJY32bxEuQAxqgd2lrvhz5iZaJVVQMrK+
SwzAkl31dnIWPK9pNevmKPLtuNOw3gzGD4ncTnsOp6MiNPmrqyRDeCTr57mt6ysLAxVlP4J/rhIh
hcuMUfJuKbTs01kjEzAnCPfAwxK/mPqlKreKPKxbCA84cRL6g/lwn+SVWrhogZur6OtZSreLQzp5
qnFavvUvPeNdc2OlsVNndi1GCej9Oa8MrDhjFXb5eprWFQD/YSJ2rFpZXkw1vqiUogphyEEot+0U
G8jvvW/yNPwBsbGvz6nCYDnuLbC6+4QrJPye9t+hQuWcOlULSE/2fs5DS+odCrwronobiua6ffGc
VRdKoErudHPXMUpbW/VAtx5QmkrAdEbLjPRK+IC84JRU8qDx8kmevidL0XQM32WRmoMIDvLq29UF
sjXIzD83jCto/2sdcNqouRVp6OZZdjAVIq8+f+c+3lwAEgcgfxaR5QAWD5zE5d4DPg8WY5aYgDNM
s0G7pNXdRuko14JVMW08+pGW7uTrUfjHGWnNgh3oYgKJoUwJ2iXFr7QJmyMAn1i1U8ASe5FYC+OQ
h0bbmDLLSKBakPjds87eLXI0D/DkrwGL3/zEmh6oWwWyd8SYwTIq5y6DoALZuYRRHYAsZaCc17NI
mrvK+ln38bMVzSENuelA6WNxhd/Y3YYsoH5BGImNoeIlBbeA6ItZpm9L2dWKmXqL6WObMujVyo2e
dBHGXOTTPjBwuMPOQ0dEr1hYknsIM8ZVSv8twyUUsObeOHOmjk/qNC0FzdSFw4sDwjlfG15tzsZp
lAnaUM7xrNg80BAHTQ76VE6cWpWPP8YlDyCuZgaA3s8PUUX4SkgHVTDoqY5ofSJ8RIQ4v3oq8MbK
blAK2R7dHoGSJd6lY81ehn3Li70/01zYc/kdceIjp+7I+K5VGb/hf5pSLwyCUgdyyk1YTd3Z1IPF
m7KUFbzSQVcD+VHH4HVReyXI8UHFaRKSGPkkkRaiED80pqq05YpQ8H03DdDAyLWnu6YYNePAdv1A
28n/KX1cCYJyDY0Xwcq1LyyEEaezT+PWrVHA6pdJKAty/9/EANN1i0z2C37KthBrG3+veJRUUX4i
NN3GwuKVe+3ut3e4IJvVfsVgIfdMIaI9BFDFXnZc448uHlnWMvsBH+rTT70xyUnVhgxDceJ/mjYb
2FcQSnrAkLsNR2SyDJsvgZJjeFsWnOnTpLVjmXfft/nYgS+cUjLB+8jCBJSMWdHE9mnLbDKyvGNl
APyci8taDG8HmvYvydnE6oEmiasbg/9K+q6gjupS06SbBg4kUepf1wSCHfbh21GEqchaVLUg68H3
1kU/Wf1sERHYeIikM6d1vw9P7KfyfDr+2c2l2yeB0BG36tVvO++KbzoCoO5zMcYrRZIJFGTuzi/F
ZcwivdMMxzqiAMt5FiJIgfZsEzhcFlh6GqR3OjT+yWFXe1OwcEOPvVAFeHKc/t7f1P2GAnaWP7Dn
oXaQfHZxgMuCthDLmk4LWQNg+CcJ5wPWDyEuvbbBJnBLzSy4Ial59JPSA1oS04QCOzGcPTFRYVP1
ptpNC17AJGRzJoPiN8jo52/IE109n6qSha9HlfpWrDTTfSAM3pM9zGzOfoAbovkYflryVw0Cp7wL
IRiOjjpXcFbfJj5EprZI/KqkYYB1HbgovroAXswVCZMAQt7fZ645avFYcLKoMi6Owe+zImhstdpk
5vPyDEAp+olDWny0sQbGPpYZc9RdE1wwNiTPMGftfOhfGseATUzhqjJwmGYJG+ywsnGDdZksWGea
L68Adp94dRVtapHT9QY99SvvZ2SYEGYjkWqNc5FMT1oLgzQRbXrvWS6WcwlqzJuJt/Q2AZUK0GrV
5Q9k5KkpeFlnXbqsKC+sPMR2Cj2bcdWyCbHrqGyfrkUPQCQMLRiXH564KCZYqi2VOP2opzHpjMm1
OGus7yZl1zWLNFC00rsu4tV9O9myIiVvt4WIn+U9ILQU6cJPQwlqb1bxWJaieyAIX0quBpjmEN81
g2V17O6uP7CQxC6EfTbc6hFwquJXOHJxU4Uq2aY4VvIAleNmcQ5de+prz0Dc3BPbKmJj/OjhMyPk
s8q7ccnnlE5+wJDkRV1diwXlh4exNPvmRNwsmXnF7I4vvcAsDYqOiwtgUTEVoU6Qyib6+baB0Ka1
LpfeEurhv4oeIoc3977eJpZf3HIykBYNhCsFumAjodUQOpLLDIeh5aPms9ZusCjwKGX45d0SW9rC
QZ+ecIIDG6n9w8yBVwK6Fsp73BJkWLLAfuCxk1gsS6gFv/8XsbsxpkfyppxxdjDpJkhZqoKbmr3m
ZqUG1/PcMolWjXalrRwGjo/3DBbpAizNP1OzxXcHid1x8HxQo8O/iYVAdEhY2XWW7HTCSMeX+5K2
vlJxcMfvkyqlYdOhTDflihNJjlUDL0/3NdFLZN+eSgW0xBAaoTKH1F3dQR/e2ur9HSAYZb17i+x8
PJuUdTOfyJ0ODdpKMMHayHpE0hcywVT9TIDGspHT3J6quPEYFnnZFjoNEwBYw+rNkjau7LK4lx+W
FflHkfeqc2VTHd42cykgMVG7R30lLnBv/y99KIemC3fu9jmDS/Qzj+booIl/1ukRo2wtDqdWtcUL
w2SGEgA3ZaMgEjKnAbKXC66bFzVYC4f4uLvbVyCq9m/hpc/eHzu45j+KBXLbwjGQ1h1GFCQdS4Pe
OC/RXNsz9b85pGLKqXHVIQYnAMf8Wfxzs41AXyHWFkaO8inCZp2TcqPgcmkCEVkkC/SDVL7qq2xh
7fe8KD1CjXr81Wvq1UyhGz73uL+QCVrbAAtE/qm8ZTYMcADzNi7xGldY/j+s9fOj8BJkgvNiW1C1
vKyKCJS/07L/Ou4o+QPtjoxwpo2G4FZo7KvY8Q+6XhWTpUxHQNPpRzTlZ7gNV048rHDmv4Ii/btH
nGm0Kv2oulc0bgslhMjNjMfEGwF3vqX/3Vf2M7cLP5/xZL5/xBT5P7l4gSISblOpaRm75FyJAa9X
Z3bGy811i4ZHcyaUUTlLSbcM2GIU0Q724bY5lS441kh2qZYD0oqe22p8UEpxHaICqMsAv5ia9pzG
usoq0+gRPtoo+9Dudk7pmEFMOZlDHh04mZpiNKAQlUXGJZWeC4Dkrjtitsw5j2OplL2+UVAdv9MC
sLODTYnQhEJAZqmFBAyHPTpYmqokcSVqvfMNefnqSXnUdsgkDlNRG3YEG/KScJBxCeH/PFeUucjh
UPIS2OB+6aDOD9E+DeQpWCoznNq/JqgbbT1ChBO/KEca4loh83tcsQymgSbd2NmyhR/x6uxm77oc
wPcqmbBr/FTfsDBdfbBFu1S5Rq9Zmr2SRZh1jKQmgnUn+MkAJftyzwVC/n+MGSP1/nfhG3xrXEXp
uINgIjnSyGQ+XUgv3HKs300YF0EQz4Fy5dz5Amy+m2WpRbJtctKpqIGIpz/ssxvjeFJCwxx7XubU
rhOXZhyIm0T8ZIy1PPSdL3TRxl2h1gX3E5IxjsdNRGn6nFwoBW3UKz+ReXIzUxAQ8Tha0S1+rrAC
63kLoxCQO7JKfMiIh2g/RopH+OI9AopPvIg6EejWIKgvKjtOrsxh2yKa6QGNbTzSgpvP52itTtxh
7ZMjDTAIUP/Ds12PJYofzD3sjXY5cC571Lah1AuCfOvbVD8t5XyW7avxruNn/oHOcyTxyewUT24E
9wyPCp5Nncbam8e8+OBwfUCm4H5UOt6RRHMcJGM8y9XB/A03ygHWlsdIzPKmdCpXPO/PqV/khp4B
snwqKq/+kuuocRRlAYFck3wk8XQ6iC4YlOYdtbYnpB3b/A5K8dq5uNj/3E9rN6+Z6s/IBJlBf36D
p5G2grHB1b01myyQjj0hoXZx0AZIXsfEYRncIenBiB5xgi26Yp7sALbLRa/lw7qwRlhs+cll4QAt
j9Nlew/v8WU/hhNm6diJfaI1H617Vbd87fmgf1yLB6kotXrmhdkvbvPnlb06qmhKND/PS+ZpXwTA
m9Qyy8ZrDFjdrmwxlUtEp2A4LH4WjipPV1vEgyroB4GkHXHFHPcQV+U8Hr6Dm4PtBj5eTkREiiTQ
TmqjO82i2Fw9FIG0PTl6JYy40Xn+3gDz7r5rj5vABTaI9iIKC/7LXIWOQ8VfcBCINFgovp/3r3g2
kye1Pdjr4hx3E4f52kNLpafNhmfj6bidqYNJ9KibUNi0j+SleZ3xJ//xcGM58H6i1AUTbBGFmKA8
SoEx1wJkJvir7nUzNDmM4PMRBrOehKdBVVwvwlRUajyVw0/d+ofQF3E5rK7R0tBAo64JJfqnvlPN
alRVVLsgdfeFjIvN6L/2nTLUspGzS6894eTKUXMfI5LXHbahos87p6nWaAzcanKY/iUXRCJGSeC7
BRhjrbfYQkY1Htj5EmUhX/he+vHv3uHr7fKk4vNZDANk4Z9Pi2e3KZ9KvVmMrq4E7z9II/Z/lZcL
aJl6TRLyVUSCrInG99OVpa+2cBcmpOLmDovI5ZOIT67Mdp+QzseIp7kKq2euOf3yw3/JVk/KIWpb
qMnbpN7sJF3fhI9bu0f6jlFC+VuhT/PM5rA+bh0ek92QivAnaSAnSnjLxsx+stzPkDE4RU3cq+WS
4SlTsQLsrgS0qOFXHprolj/tVOs7A87N1fwjeIvHOpw+ZrewPIeWlikeHBonRzVC8G1xWEvYBIO4
z4Q7jDKT8gnikToecFoJNVIK9juDYLYR6cT+tFn67+IZxKhFzxd/5qk81QhR0pT2iLTxd/RHTee7
GTxd1qUh7kM0gz+p8yJXKmzv0D8/FhLjU6u2pDYK6K9/4i9SjJ6Mdh7ZVVcXHneCcHNZgdEhg3jd
PUjqOD3a4AXLJc7IEO6bNzPa6o0jwP+u0AhGKo4D+gf2tZw/W8GdnM1qb7kSPwU5e8C1t8hoXGdL
z45eakd3BcHwVwrHnO5Rpu4iZLyjh8B/7G2IgQURGwK9b6074vBMnxK5Ay3Ajx1jmHsC+RsOTSPR
dt5IeEBCSGl09CuXvSvzcW3m6qmHnGMxTox1mf6ujFCYCJLY9l+PKdP+jIPaURGD81gnQg9/1nmO
/yXUXd+6J+LBt7QXXSldExqDRY2nGvF9kz8P6xuGdGSMyVVZ/Kl0pXOgUkkvDLmXhzg6aeE2MRIr
ydA2BCJIptBZ+xF4jtdsvd+12vAaQbNJ218UGZ0Rq7g3cnSuxgF+8FMYVaFokcdYsxG0za1eZl4B
6GRU4BqBBR25NDy0QNi10wLvlImmE+9n+vGM+PxsEJ9Px9E2d3Z4jCaKhZsvfjmkCitORglo2M/n
m8lfzqnh/L0jQSK1S0lBWqaPVVWs66bP5IvwxxeWHYz+OYPBjW4RGDSe2r9oKr1W553NmIjrdBGt
GwiN33KaDx+wcHGW+evYrvvzidXHp0iGdof2fLu0DjIfmtrhgTwrrGd8dIkYcS9Oo3aaYwi9d3uw
1kMPn5w18CI5oJPumVjO9RFo389rPSNXbnQLXE43u1AB19uzklm/TF3GNR0jPjqbdenuVFF9BfhT
XI81DzJ3SFP9nZ/PVEhSaJ9uuCz7ujvQERQi4npHStW1I/bJm1Qyyv79HGdDzZE35LA9ImdVfqmV
dIQyINQiB92B3U2w/inCDf4dqugL3+KloLN+Q/XAtXSbt5wKPryACFt2KFKeANRb7EfBbkecFLfM
P7wVm+39vobJwf+2xtunkCr4jNqZoMFm2UMzauItFD8WQdp8Cj2xbRoAe4XobqOvnikTmrnN9PLL
WO+YO6RDP9iemkk2W1ahAHg2WllwWlqBSflrHU7mxpxa0ci9WQuAztqWEmqXlQtdF0oViYqQo1sk
bnBXTOXxdgvFdu8exniNWd2Qom9p5vJwPPKeY8IgqM0plDEA649LP0KhjKh0XWPHxUqW1PGU/1bo
fB9cpSjbWdW+HNZiTpDRUnrAntGUPgW/ZxwMS7zWhqRPERgA8G2nppYXYye0QKEMZja6MAHh6qTb
YuQdUPJkpaczRU3zh6UeADA0wYgVlHKI8vGl2ql1V+WpIiwKEjajmk7MFzjm7l1xIFpke3xnrawZ
C6XoNptGU69c92/LY4cShA6QNjfSU2BxUBwvvaBqp+sk5q3WKVWKRVLC+nJKmkPw1BqeT7H5Bp/5
eNWYTRPbRuPeZ/OG3vU8GYnYdLiYXxo3iDNm8+3CiHBZFh8mfi15emEzgGSrGQE+zucb7bwNhhLO
42RWxg89ERq8bhM+Enss3+FZV8ZedG3wN/qAMx1yEMO7xDFzAd8XpQoqsVbD8boNexC+IKWvUeL1
wKKrrnihZ+kl/VE5brADRDuDVZZrtcSAv1o26h2lZmoCd+bacWvxe2ZnwC48CmTB350FipdeOHHS
nLMQmYdFBLLa+I54zjkDQFRldB3+kOchQlIUHYADgrYKLTLiJ99x980KDvKomGW1D81Sxo1zzJ43
S1gZp3nq0xSZiA4MwevqHn/49/z7UX6jrVDVwjN6V6PJAJuwDj9b1LixR/mocZmCie2Q3Atsbe3Y
xDG3znIo9cNYdyRhpwYQ0dvYGNfvo8dhKBVLPzH+UESgljqpWKMQlY0V4GP4Ulbvkgh4t/MMJO78
efFIo1P18pZVRPretnuYVP6f4eTbQMJdc9AcGZ+5BS0Wnq2w+GrKnwhK02qghPgBnR8toYpdMql9
ZZ47tGkcQDLpM54Df9a/6wX0QJNz0o0suqohX5ASxiEgLtLzwmgUI9fKzacHOOcELy+DOilIEe1Y
2yX8190CKWvRUrzEZI4TaB0jOhuRHxL0rEzE9F7b9xMNOVXyMcphG/0BK+zWMr+qW+J99PraYBml
DS2vLToBjG1moGrO4lt0bVc63TYIvBi5Fg04NgstFFd8JtpC0tcCMRyuAEHeUtj7kLCMX70D5fTv
1ao/AccpjXPbhMilC2CNkH38KTOcSVx1nNenYzazRiKk1Tg3uCAIQXcOCfHRqxN6hvOYJFBFl5jz
keCd5LAuQng/7eDNdY2Zl+KG7mED6hZWRdLItbW4EoGQhMPAG9mDpQNXRUeH44WYXGE5gJIHtcP/
0JPdZqBWABxsLsAUZ/1r/OK7e37SkAISFqwrWL73iG8wFDvr3nEfs4nJ+mXl+CJGEsn9J9ksqRTB
CqnRAW4M6mxmLfd59NtXKH9lU0vxXk/ih8Q3ARK09xSqX51ru8+eSVcz/+CXlvC/hWMapkulqwgj
GnCY7+1A4Sjog6BrGTCBzAwyyemal0W6+ys+vmLrNkGXt74pZnoMhxU8wLWaE3ZEmsjcBnhkZPmV
WZbEjWgy4uXY+8iEWC/ju+0REcotMMyiNW/lxWoURm11/+gNvsLtMIdizo46Iqx3z6vuu5OkmyhT
qZTymON4rP9o6ybnewDWJZHQN3poqy3D4yrv1OuRKf4M0qwGTJMpANE9Vzbkpxvi32FA4qxpp972
qxY/Fm73C4jZ6RfHiyh6CT4ftUNsSJWMYp8wiczFjHj2RcRezY7HPqW0ioXbsEqb2DTM1U6ZYzvX
8AIi3LrHDvWrdme2FAYUcDkK0G2DKcIfHPahBCJpsw4yb7BtSqhc1MvsM13but/6cnwhZ0mGyS4R
ee/koTnkzDVg5Zx4a5L4wX8awGgUjYPCNvDKJItyW85tniDLYNBxE++0HJeknkYRDm7VLGV+azRJ
HwVqanXoj0OicK+UGLEeGiaDqvEQTr4ZvjVWYc73KJx8i1NxWRNJdvB80PZdO9nRf9Iu0JCBrnu+
K315GnqN3p8VrQuEUWQxFWy3fp0xHpNPgIlqeUfSZPlpCI8swqaRzC3+3YaPwV0IUswk76jc5x5o
TKRrUjZyuXA5qbnp75Hxq31greszXTRnra3qJyDvIpA+EFDZ+uursgbcuHt6IqSc+/Rz/A7sEXK2
ClH2H8ajna6wNu+0aLRzivGBVLVvUDtv9el86i16RpVx7rfAfGggOWOt2G5WltzeWgrDk6eDIVos
Bq84LAGwLsFlnVYytmEjbcasI8cfdBbIJplNzTFjcHYC9oNXfTwhIInK98jl0BBxKHNLMl8hcEX3
YcVyJ/+KIk6a+6UGHt5sZnNhQGIMs0P+0Smd9VzUWrZaF5Q1oqY19g51vwt7nEOhsMSoBGbKY3Or
7OGQr8nic2qKsmqXMCvLpnJo0466y8ecFOkngrunZLWjHFkqsWyoPyTVr6D8SR7RFoxVu0gRr/lF
uUKF12N0KhsRl1aS83VSyl7G+k4o16vkSZdUPiOxyVrrtsfava4V/p5mcGXrXTiBw9//HpNAXU4D
vxzBaMvp9NQbboiGljVTLCOuDfdCqxSt57m15T4/s3d4wYjsIjQKJK8+P0LUTKIokfxcBbUV0TKG
y8ONT7jelqWarw8xvsNR/3wbaWqb9d+wd4jIl5B+llqiemdgEiHjtO1w4Wm6k2ptEImWnvlmKNXd
mev1/DxUMMJFMZwD6w3MjHIJftgU7HeDojVoSrO8vHoZ79hB01Qd52uwooZRNqLHYaCo2u3RMbVx
2wFArgEVTdvz4kPaucM4mcFHgEuUPrlNbRR/xEsyKqpQmkSivAKu3k39+zu3RkGOVU+XZNKMfTcJ
Dl9G7zlCNdiiNvy5Uaz6e3dQUfT8x+9PgHXtaXoH8At/zeXTg9DY8Sr/Hx5n4XzpvmFdEqfnTcbp
Q5IWsoYQlNGZ/Ujat2en3ccKY4fdWk0zpBHwwkSkx2mdEWhBzs6z7/MXeLdDfeAjlUw4YLKlNb03
T/zODUJM6wusgdD10ryjzPw2fygCiYIo9r2aITb4xb6pzmgfqBZFfC2U4t+tiy8vRZUTrEc/Srdq
yBzzFB9y8u8Sreumr3kVIj70BxtBMBnJkX5IhOoeU4akhd/uqWJxmxjwevNdK2lcYqGdIsT+ITyV
DilUGCrpxXt9VOHT7z+79BfXrsDXilMOnz6a2+xW0I/d0C4eyZzcTuT3xRtL0ftgEQ9kvpPRY0pa
7fGIO8JrH341czpONidGCTnjvw/u/t+TxsxcYaoSOdam9Mt4moRJWM0xxIb/IXgGQ4Awy6v2y9hP
Cj+GrwDpS1aanKLwoD2+Zjk8tVMGDn7KIpLUgfQSSqgTBYh9HoZQ3RnIC6zSrbGfQINDDVpJTs7H
BHnqCOIgA+r/hPdtMoQsrMIr6K9j/DSsShQt5q1Vxd0hca7gAvramGZLsIQrJ91sIK4uvXiC6OB/
rGZUI87bYOGXTA5OKe+94C2d6lWEQ/6Qh+hFkpTGKADDNALdHi5AqPUJaY9JiFT52G5yTg06kZEF
2GCwApokWBnvO7z/2HRAU2AFC1pIislblOl9n5SyCGaLDYrOpQZ0Z7OvjHjocE9sW5y0xRcHwWjk
BGb7KNFyhpVbKFXesdMy9QXWvXnY7KWVBwocOfw9xQSiRMl3mF3EPHd7b/SQOzzNLWThwgysZuNP
mSomF0G//C2XxkHZEcIB62iZ4zhoTRn/7rsiUvoDrFcoRPSsa+UCaYlfzWCA1eKJfknlEFs0Qc5K
E3cf7/VlN2A3on4CIaU96BjVw4WzaM5X860B9Zuiqap1myMZjixag5BWQAmqUBxJyjPc7U4uMRBY
Ki3rIdMmJCE/jN+e8YTWs0U7bBcjRHvd7cdrrPGE94zTVAFKC0Ljvr1lGRGoSbLyniGbO2VT8KJE
MYqBXTka6o8ZbU2+tmV2PBvLqXixaQnLkrybpTdk/YzGOCtHkuy8lluQeVJrOeJNGzfOFF26PTeJ
3nf6y4DwlKfhSVoRH432yAtZS+XpPsT2y+SqLHpbbmLAlkvjcXSIH4+Qwh3rhj0mwIER0TQF4na6
9xQ7lacG5k0PsMdsZvHRm8u8Ge+hxyiFSsiuXyDDO87dJylQTeahZCSJss3jDw2LPUmAOfJrGOJa
AXHPersEaIKC1Q8yCaYFbZCae8V/tyIMO1J6A39PITYpspbTTpK1y4qDOWrLofZATI8hxfGkWd2W
EkswQIurKZ64oo/UzVYtQ64xeg9Zk3GZopYnlMOj06XLki6t4JkSdCpQtZ3SzTZ4mDhUvxzNcYje
UT1fnEJadrJ0IqP22PWa2KIbFmKFVTLW0VOjvoevNod++L0RK/Gtq5R8s3S1cXrZQxaaUuqBJAJW
+V7z0+QfGx+sDyXqoElU1tenxEZNV3gNeRgq97VAS0lyHLbTKRY2MU7P77d1rCcvz2Z9tvOdn7Pj
X4y0XYTrvXh+VIjXoyrlvYQpkRhrL3AfvuNRUJqc3BdclmNRN/mwiSUlAevOK8t+RcU6fiLvRqSJ
fdRjbTbp+X6Tlf/HYUfi3tz3k7H7+IQ7RyKQZrbseYLSJ4pMX0tWcg0GOIvlvF93XPTicaLI0fuO
EaHR2gYg4Z3EV969vp7VSEL24XK9LASZCQXBsYbKI+GHqieWxGQbsYd+sj9J5egE8HzF8gzij7db
3KDRDNzKIg/mPG3zktXimQfZc5Z+JUROFah7XMWTHs+dCIHU9JArnhbHWgXeTk8LAnlJpLTh/RAJ
bkx4IqoBMEtgtFhw19hkG43PmxjiOBrPa7y96RYfGH6mUv7fNkTlTtNdBkxSddiUuS1UviODG8Y8
F5QzBvZ/7ZilPHbH/x4j48nzrsgYjFUtISTqP6Afc2I3YA95IcQPF9VetXj3iLctI7a/yjDvn9Xf
cXRJLmQPS7Azt0YuP3IOWYi5byvtMZdkBJKt+5ovXM7jvSjTWfnWJSLtE/qRbj+YG8MUSgIbFJ61
EUHgZEO8E0NguwvsucQAf/oUF21M+aCDKo9ybILybwd6p81+u6S4IPkWpfRpTWiw9qLk2nXCwGzb
kwb50rrs+h+68NevlU39rK9nfCvuUWI1EpSuvpLnYDOOm+YZN7NO5s3A79pCah7A130JloScvN+E
VtfXCs3+XETG59BFCZGTzPtMZlGRR9o0GepnDMvJmzAeRV4UGDNZ6N2ULVolvPFK8JycC6+o2zeT
0NGurIiNCKpb8AwZeNZBTmUxrPRv6l7f25es2XmEQZ0PIdRhv+UtbLB4aLIx156gclqOShDOU6nR
lHEVY3Pe0BIkYGQh0EttsJdw3gX46IaiBv5wd0XBzdfoxsTHSRsOxp5A9n8lgMXhJIeSXgPCbuU7
ed89GnIk1Exyx4Py8Jl0nuCQ6S4tyWvrHHmoFyo4A2vYQ8eDJxKkY9OKOZRyjmzlThvGRJ+cAF3x
hmtqeDONpMIoocwerkUPrb1xu7rBnmsF04/t2sIVqRXXrA6mqMjfhIEJgJ4cPwUS6hujCD9Y9Dgq
WiJ+aENqJwziVZypqjXQCyKQOQy13GTJRP5i4qTOIj7hMgjsqnjQIYJp/a4dniP6Ogs3Zvm6iXwj
EiewHn0RCzNFX1FciLAULP1LnTXROIYbvmY0kkFHbJ3j/7YBJnuaYbsNrmH1PWcuiQCihmuhd9ka
NrrO+OKxfWu02j11uXq1KrPKRystpu7YNwsH67p8VIQyA9M+yrEHzJJNFT9MDV2GOz6kIq7cal/E
cdkL6Bs6tXqEzZjgWepn1cl2/3jyGP+Ja/0XPK9neeiSI3RlyBFSTC4RfTT17MjetwKM4Siv1JQF
Jc4PUQYtoWqSX8uCwthPruBxXunHNB7eVHiVniv02eQPTTF2y4d/2Ad3v/4C/4FfyB8ykXLQxIKq
nPUuh+JqddHkdnodp4NeCx5astZ6E4uM+K9DUc7aXoLjqM2V+FN3oT2wp9z3bC+EcRc6IeE372k6
tgy+MpI+zOFibIPoPzRwo6yxketD1vIpfpxdWmbaH6zZARZtmK5R5HChrGRWRA3P83sJpp13Rxv1
4hjqYnM+1az8FDmP2P+lY+TcTgW2hct1taxiDIW9l2jt3aM7cGf9qR/Bl/LLTWCpo0lJIDoFxDj+
aetoccQGrkOVp9z3opFCYeJku89DKmL1eXkZS+HOjSR3/raNodNKL6bxGvX/CIB5t0FIfmrub7OH
UA61tGmYxSJ5LPTLUdqDS515Xa2x7y44nuN6CM9w4SXDpjGMjCL2+1/Tcyk54bCFzDZoYJeu+kql
KO2Z0jlXtEyXH3m80A1mHHkkXi/eOxJ+bB1Gtxp+L+M3LAESJ/gMz4rUFv7QG67l6BDzEaATCs5y
ZXiEL5OBgiapsgXwHyVP3BDiLj0Bzh6i7DfADmtZnb7gW0Vwkj7+pO7zn9+6Y5TsPVLE+brtUNXT
J4i4zqbrNoWTRuVgNSbp78t11QvMB4li3/RcVPMEv1wMNjgw0bM6h/zsNYynIeEussc9psQQhy5L
KtpTE/LBuCeGujQucR3jcDFSNdaB3bQTPzPKSasIQ911DRQrDqBc+Z6z0G11unL0u34toyaofQ7y
drZ5luKmG6+vzAsgU1cfOzztVLw6J1RsjY3/L2SzelUwtU/apw844REAr5NZhZYQGhGOqetdOBy4
5rlnRM8JL1NBxLjdj6Kk0/2GykCjK8M2GCYeNBs4GvahHOUpMvCPaZmxa6JPkwQEs/6pfDEzOcRM
EW6ZtDwfqzORrM/FP/IcW5roLk08sQWgynq9AF2ij2fdNVFCPW52XvGliZklL9ktdJvCKXx/+7KS
rzwGZvhgHlnH5GR6cGvN4fk38DaPAgAMGgXmn7TWOeb4+k/TGRtR407qJps0+qqUpEBigS7VtYQU
xSfRdosppVxxk7WTi6b5Pnt92YjT8Xj+eAYlpts0KDXqeZa3b7Nr2sCVaw4P11LYL20Q638vCNKZ
grKRR37W5MTDlD1aOlWbDKPABat+4PN2eC89XhnCh4ptCJG3GOnJ1dgsZVI+EomM1jqSy6wrXbEf
uDT362m2cdIZ4F7VJn3fTxudK333rs/5lK8iz0I6x1OIBLfIGUjTGpdrBOvPz10v5jFXhAwdDiRt
SXQqiIoxlPUjF0KUeS/RMb7/iNQxGdLM1vPHRTV3dUfhZGSrYQdG+uQg0fAomhsEI7SUvMJhawsG
WwnzeUF2OlZl9wcwr3QwWsN84YOd7T7ywL9z5nAcSggi7t4DP2v1HLLddym5v8DvwFE27zqDZe1a
RnRqG0WqC1yE9lAo6eH6+oWHJyx7lWdcEhCEnBWXPTrHWLSq1uXO+M7xAw4I9bRP3bIut6QDBUFU
vqhoJdsXPesPPjJClMnVodXu2uhEQkMC6jjXqOqFuPCqAvRyrCLgbB/1csSn14L7eyS21a6VLbSd
z5h/OP7o6DgN8xEcoSj/W8LOsCZIDWHColfyVaKkcJlBxwUO1k3xG4mar4RQXZddI3OXif22Ne/7
98mWV2goDKLa1cnSM+idSaIzEbt7IIxzBG/gThArs7oc1qLBERhde62weDBkYPgvmvjoWyvysDaG
uUZ6JA8NgVbpkgcWumSvfkPMPh1txTvLdpyBXKEoRoSjdUA5tGj6PpyzAKfS5YvBi0kWMJQ31cVM
CCpdhlq0BXwBa1n6LqjE7ytM4z/+7UHxtOCFlf3Um9aiZkh1qXG4jnHEiUulOb3W33prMKYG77pG
SdEwaZ5yZ+tXAmax/44yksfN5m72LGdeN+zD2NIpUbQQDWYuvE0jEM82z8MiiHVwaSWOZsT62UZI
F0RNEXlYeK0xd5bZEThGVRC7ZfCl0zkFWpe+JE93qLL7xVLWWIypYwO6a5SzGyN8mTkELUzfqets
bJEHfZhBwuq3/dMRlpafXyZI/SQY201Wagu8hqDsrmzAjDrdkeDhmeR8uDptbf3h9n7nGv/8e5Pw
mu0/PYuQtSA4Qaj28G4XnbU+txeT2jHZMPCE9qhbTwkFueOji2hn4Lub22FTkHm3wlhdQkUBe2Bt
kMHccDx491HKZEGpBOaGh0E2oi4QyvcqqlXL8l9ML0wlYPRfOn9Pgx5hGo7QM565IRshup/6zckU
mNBaShiWDzzeA+lVX6nbEry0OIE1EeY9ZqNrGDUorhjs5xEWC7P0zjnW9aNFZ58xM/Fx85x/F+F6
ZHsaNcK89jO5vE/Nnoa+YvEM9M0iHR6bPT5ilJWkIIjTX2p0QDTAIXEYCnlMMxDKU1iuXp+xNbV8
gYfeDZx++YYzb4VLA90uwTSkG5n2JbHomRcxfzku6fXUEuWqUPKsLrp8eV6S1qHprzhEaYcWCnew
3/z0H+Q38KLr6/vsaScp0hEBXRDWHlvtFNao9LiSe7c4WLiuSrgX7LHAoYjFO7ynaMhHJnsuH2Tf
WnIfYk3EYoMprR+ypT3q99tZf6qmoJa5Q4yXJsvkLOtZQJYV4uIyz+qoecx4bl9gumMpyGE0G3T1
w0Str9FDbzSiKWRmGYJwcWxD1zeztxrnHHUhKn1rdimJnN+2nZSKR0+B4SulA7AdehGug3BB8o1+
uADWD+cH3OD5eKrR+yHot2harGvTupj7Yiu1Ss4X9ur6Zx90yRDEfL1bLYGbb7fA2k22XiaYyR6r
OVNSlkXwZOx4ASqIworDKb/XaMKAvrFLo+y5ppnsD31t/eep4W9uwEG+zSIoLMgrGt5+rD9Rg12H
c3EdB07tKOmKkDQUe+6WwO1hCXlGmpik1Whasxrz82ZF90ffJEgZIHLqdnc4Zi9LciTg4Dr5JfBa
NHfJbAIeyp4QSQFGpcYx5tM+EdkyXZ9O1eOncwR7aYg/ik6u4uP2ScbDjKpRGO0GMrKPpxMqJxi8
WqI0l6PIeaP/VbHQfkwSrKJTqutLvxs2ZZGBtFSj/BfrZv7ThY87H2vi+CSadphvQLeJlFzIptTG
OKASbmDBBCn6qwe/hRsqvjPquyCCbneC9l6KVHkD0BZ2DLIk3EtI7w1w+gP8nGElQw1fu9BSmEYg
griRx6srFUZHzmC3Ftmm0qt21K8XFVdxoLn8BttrDcYemDBf36ELYoth/FUtZgQVI72Clx5a0xoQ
3FdePXaPJ7+Y7L8ZbgHFwfTe2hwH+6+oWAwvpj2UBqTFa+dbtOAZ/fp341p5YRbJ+ufxB6bTuPEY
8JKdpO9biSd4mhXwXbBS8ebEqweN/prdkE12ZoRitFfVLg4T5FhLt84gBwemqjQEOwBDZAj+wvXv
ZSaAmmv3dl5MEqL0EyacrIpnkFVIId+kNZt+/3xrOwIsAuA/TXN0mAY3sjezBxMz8wV50RfJWjxk
Kkf0xlwHXURRrrnUWhjYixrHjHC8BibksyRZEm37ajwdDGh5Fj24YPdrMqhAw/Stmh07VW9Rt1Fk
2NlaxbcgbHVVFQU66JsMu0xSObuLq+Q6E5tSPZqeLM6jfBYTiHOA2KtZP1OCeMz/RQ5mg2HgwheF
7EDJI7x/r3SENGatXwc6h9dV/CnMWY6dNcoQGnUnz8MA4UinOAzPTyA+cozTzR8a6Mj9SsHKtBOz
KufZ39Rf59hVnnCyw3NdufrmFajYqKf53ZzXbqp9MoheCrDcXfZMUzsPynoxqKJY3o2UFL1L/mTv
Jccvdm2p0VS65I9uCoUgEyfjPQ4s7xgOZr1fZUg4xEiTex2PynyoeGOWj3v5zF3/Dy279js0XWIA
YRXsyOfIOvMoLObNXKQVa3NGhAmYckW5gM0/NtuLOLK1ko6NLo4BJoQpgB46U2QfdN28Tos0pW5K
IPOmNtNNdrIKV7SPG0JbfS2TLrj9TvGZWGkPYRxC4AlazYEn2Yal5zJ9fsNRGLv3rHPk6ryGAvAz
r/nrs+v670vZqBJaavCrUffIzW57jhozq1oe9kXd47ua3+Bs1p6WlmP1dxf3VDsUNOoCJ62laGWg
PiNbt+xwcZmLNKO5P9z2suJnTnoJE4PKfW/nTtYxw7nDtBj6r8Qi57qT5bgGcwuQmmgMO0nGoaVv
yNbev5mJQShamJaz2Cz0uHs5G2jwJswsCjt5pQYPTJts9wOCfTgv+W5bVxSAnGRb1IVYzcn2wIvf
586L2qmducGaYA1DJodtQbVzj6wT3lA4m1aCNMHEW3N9WiP0yzMQIguDwYCl+cunAMwELmk9q06V
WTIP6yul6rZDmHSMb1sJHsDLPSWoGn1+gWQurvN0Rc3IR1g3jiW4IhcB2TiOZSdE2verKLLuMTJY
O/hW5prvvjvk0T2uCWVP5NofLBRbBUuzlmsjzjUB/i+n6VtlU+wA0pfUqYkQv8W1fxu7mKldMf80
GbW3fOc33zrcou+eS7cbzzIXy3pY+1kNq0C7beep/eiJa9onJ7TNdWPg0IGHpZWX0TbMAXtz2X/N
60gi/uAPHKLpkHuOm5G/aOTw/no/XiLgGRJgapobmat+UrqrsPKjxZWWJ3AEE5cv+b0C7Bt8csAw
9yTIsTJRbJJenR04Gk4u81xWACZMCBXLM29jwK86yMXrLXBtUYE6Tx003U5AyRo9N8rxJzoCBL5o
7ssV5Yaq5q8I5wtRyoB94K+Q5ucHqvSX0QlpVZGgyVPGkt4OkDlxX86H5llAxchfzd2SoZY38F9h
glyF4u0ZSv+UqRPkQxW4D0PUOtpLdUq0+w3dzsuOT+9B14SUzJix/v+F8uvonZG9qVbEIkF4DRSd
hDocfWLUSBAmHNr6X2W2EY/CqFiww7W2iHxTVhdUVD8OdMAvmFNY9bJ/nEmmOrYphneQKjPhw3xE
Mt8tQtO/6fE1dP71PlN4zdnRhMcxOgXlZ/w0irkeenlN8x4OlzE7MI6rF+pXD/6ZxBDYedfFb1H9
7oOixmH2FBxqv5WgxYj3lsuC3iCxR36ydAAkj3gyKthahGfA5VVuy6ALR5T78qe3RZCdveONcpNv
GqKHVyTUkE7BEVpfKOTKmTIEXM06NxBlcmlDQjn+JtBQFiu52m4Hb8iDrS6oQUosadzvEYDGKerH
ExwTMPClpTCE5lr14743E7AoD/paPysJKkacv97SLLYEeqi5OP+x1r2fMXpyWI9QgbJ3oOFRI+Aj
vjGUj2R6oqzrFWmylX3CSA0YTLPbygItn/974cG/MU6p7fL8W2bskS7V42UGzCHrABPmtW/wBg1Q
aHTekOojmYcB1oM3ZxAalzY5kbcrecvh9M91pYVmzv+k1w+GNbpg5OcGnhVuzbxFIt4G0YQFIa7C
ThnBukxLWGpcIOlzTwCHKO3oe6nPJybdS3YO03QhmHupUCd5vEztADUftF4ot47mTOrMTkXYKs8T
4GBXZBLc+Xb30aurQov8S0tkJxtINpt8uqJw52rVeL4YfSxpiYOCynv1QNrY/qj1vhHBVK6xLm4H
Q7Xv61YSSMe0mas6qNP25skq83DtcVYDXUsockjtixepV3FqnpiEgEej6lg58ZAFofHQgEIogt0B
JhsH/4Tl+WPwHV1lIPJDM8qsZ9XuBRE3kvmRqDDhdKOv/cK5t7Ajpo73gje1640Qx7NfZsd/rmdv
kxqDrLw+lcx98JBeSMjAg30ZAHPQT9mBxoyw2WpKwckfUkLaQUEwgMc1VryF1Ur6/sD5y+45p5LU
ThTy025m1GtDnqKmyONYyU5l1wFeRQWwxwzZq18utlUNlVHYelPI87A1IFft8xWV3Z5ghNGKU++f
iiFmZ+Kp+mrZmLWrNOaUB8vDo8sI9q1Tsg6AQCbo2fyY5bXOm+tFbIJnQ8XCNEuxOg516BDkwSEm
T5sdu4YC6R70GXQsOG2M7HrF34DEKSGnmsfluWQL/hslbu3YaLRElsiCyhivZwHWAVF5xi3XPY3g
wa++fQsWPSAgk5059tfrJcjKNax71SbWYeMhRJL7NbsrbfRiq2+RdyPTwlhoDiLALDcmFarORjQa
2jxYu0ZqU7gR15m6fVYiIVmgM88lICjpdnjXN+apVufiUS/ponalD7pOeUmEYtrCHPGbys5xGzhC
/YyX+Q0DW7JVQ56n9PU3vGJLBCxN64fDVpqP9yW1gj1a6JEbRrcPhOah8TiEyzuQOuvIQ7CfvObC
bPcB4iI2Zi8PvMupr0PUabnzCsqXU09o3sSLiLJTpR7lL7bBJ37CqBDUG0Ffukww2/70LCu2CkFX
HkGv8R/I33HyRY6ngaie6DLgHdMxZ7TkOWKEKSFzbgnj5AGetYIrKj5tXn4Hn3CNRWTLqYpwZHhT
SloBH+BWq0U2OdSCBYetETQX+rHu0cmHvLjx7IU9/cttUQk6gUP/7DKnzL+mWSoWsyEiMBIJEroH
vHhrUaRMiG/QUxZjYreyVsQDC6K2XqmP9KMlTJl15/3SNED/XJFjEJPVEAFWK0ndt4vVHrDqoYE1
WHU/03ALAWtKfcPQlMyVe/DMqPS3isrcnIjC0a1oel2hjWCGMtsoRbj78cbRdtutZmA82hVML42Y
QDe88/mNM5eaX7FngJ50di2DFN1Bnm1gG0Jp6RZWh9nS46X8pm4EZ2mArx9oMcI8zlDl5xMTBlgh
pFtK/hi8w1QDz7pfIpkjUMJLb2jQg67TAjgAbXP5BRH0h2pVCYHzHh90XQArnHr75TKz5zXdEdTu
j3JZKS1Y4Sntsyy5g6xvUVqZpkeayctQGLKu/Op9t9N5WDdq9ihjGwBS6V0JbMuZScmPg3viDWPk
x3QBcW8v4mvXDXANCA5uVr5cpjm8sOmEsKVGV8xYORJ+WKC0DyQA5nDvFy1LZ0kVu80qCPL9djDF
bbkZanSxcMWEBLzdMBv8vDFpKh2oYSOStgM8+D52QOQAC+/cXvFe3yFWtrPgjRjt3g/nsdyegYLd
d/ApMllbAv/CHorXtiTX+7TNjDYIMcPRCh2QPUR5gxVZ6MX7MjiNVbcDhpPFYfaW0sO7PtE1JHks
A/EhsvZFu/kOPFFXVFa12G6wSK2tbBYh0pWlB2WNI3INu/zz24c84ScvPi6HLxP42jC2bhS6B10d
Pi3xweX6EvJsCven8ewqdZaJmhPMvuUZpKEXldYTSKsE4Y8fxn+aNBV3d04UNHKFXFvYuuGpTFQZ
w6KL1dLRZ7n6ddWoV1opkp+JD1McKWzL+fH+2tRDrGflmyPYTOxGBjqgfDLxnjamsJCXVQEAUiIl
TQW9bS7i9H0Bilr6Ky63D7C4ppuBYywxDRKv76hZVyyQd0WIU+LjKbl6bb6UsFxwoC7kdNOi1j90
Y3BYfsCzcyxFx1pZUlOVv1rj7DFK3v5kuX2HiNEzyAwki2X5YQqB8K5WTDYGSGSYKVO+ffIxQs9q
+dAW5WlbGCyEtzhnJ6wZ4IkXaGmxHqA4dYmqcqOWmlgWbHmbrMfEnxoifL5lzyU9N3/KndX6peMm
F0wXVb+kjKLsyGyER6K/hpJPQSLIiBe8JA7TwJQ6ZWknkog6fl7c8nNYd6T9yQyxIN61+c+VbF2k
7uewKofc+ApnRPFF80Iub3zpGo3NZPSbTCAEl1Cp1xEXqWUkjQ47rfthyxZE3rWzlqfE4IzoZVGZ
Ezb8e9p1xA3cbvrVEp8RCkMhXduwipouiClGKd5sPMbHHSpslSl0Fyxo2O63J39ADJo2valieqiS
CUtYhNBSnDrOT4U4+fRQ/IHGxRAl5kvd8DCSGoSvHE0jl/Y0rYLeXEgQVTBBgrZMo8A/pKZtc7FP
ZcgKepGQYrp3fiXtmUvcmvJqQwNuPHpgp7+nNh2MRHf/uPLO0XFq9Mg30QyWLQMCATAR5C4XXSs2
nTlGP5tQ6+cjM/tQyCpsHJFu/MxWomABVfR+bXSqfxWXuuAtyqsBHuVnEXIiBc2mYbMLyFcsP0Oe
/vordOiXiTAjae6BcUE1pYCdkOCm6jILUFECoym03/N4FTaA+yar5ItSFdQpZcbEay4Rlsz28Dcz
RnG8UQqVf4v0WeEKla9bgWcXmQ78bLipgfBQpcSwyLcyT+6j81UlCEM5Sm/wBUl0x/uoQo4waEzm
YaiVwGNLMLylmu1AL9ImqujxT6RPlpy05r2O0wKbq+cwchEccw+ucxic6++XkGLI3sdDLzmnmdcU
Aknl9fYZZqE5D9WLroC33bPcRGULZfKB8M3P7NG0HmxiMJ3sQvTGNL9bYpltEl975SeSglU/ys2E
s9crZhjFHvy20nfW0sYTmuv13RpuOiWkbgsaVmGsuttFmzxruVGO0hNBCnGmoQI6QQHa/A/Mch8Z
DPKdFRoIuIt29lCn0ju2MQgWulD+DN9Lw7LI9Ue7jFxrrnGRWu/Xb7u8E6Fq6SWevO9RdOuuM+CA
OlRrBYTRoI5by4I1fS/HCspyqYqmPDvKxdJgWOXWaaaOQNNYtiDkUfV1UO7RVhSYrPuu4CXJ09GX
R0Z8Jr1JxKT9YYY3w2osvObiNTWt6a4KWRS/nfU/2qWyR1Hj2mCGvm7INFqk7jcMGIhG5FrJH41Q
KoUIYqr1gxBP2uAbYmei5VCGN2u3A3PBtFy94ogfqkShslpHdTFAw/7bk2jtrQ9xWzgXFUdhkZHC
Ym90yL8/33QwJPSVzeywBafnX2wceki67/mDQ+0S2sSEuu6t60boKDzi6k2f4P9Obf5hXDhxWnl+
Kv6SecE/lktnkaiMOTry6VhOsuwDSpxGG3bIgFjUk44YMkSY4tBC4JxAwUqTrOqT6fe9lcpoZ3vN
0Jmf6fY24E7b3rEfuDg9p2/cUHVNulRvP1j1pVZGFxM6EGkEicgoUwe7CXMq0TH6xa6Q3KfkUqrB
yxkzNWsZjUyw+anYDlay2idXwT96uQCGISFltyKltG2ug2H7XbIh3H232gzp4NUqAmbiRGhG/OCb
udQYM8EpxfjK4Mt6aDaQUp9V8W+RiEnPro24Ogo56Ljc5UZ6V1jt5DLnQbMKMrsANsYS96oFbte7
pWxPmVxkTIlcagfoItmrYi4Bb0Rw7h6GxkfjImsU6xUTs/vR6768K5d92y83ttuMpjdqTwM6o/FV
qHKUOPFXS8u3SphnfKyMdlhZBOm9C+wOKB1L/rIaE30viDYpAt91f24Q26QNsr7IqpaRF87H8ta/
OY4fOKmzg2iQGTD0CCuZl9hg+AOO1/f4Di8rX7Tgego0HaSVftIbaijqhI6WVjXkPgyejNwCDNhg
Ru/gboFOP+purN1b5MeOopnf/7FKwhLURMN8jxjCOUEv+nnjay7A/icdhjOb1E7pIEEBhr3yv5qs
u9CL4xKQFPf++4i5/G8QcGUf3fH7jFSjMLDCLnJ6+2v5w5E0cAqU0jqb2X4vqQfJ7o1Gq4OasTer
XrKDk7yLRE0o/C4NVT+be9QTd6eT5O6qkdV2qfzTes+VpOnttlVi2pL+g4W2fSx8HwllAnWFnVrP
pIXo6SAFFSsB501ybJS+U7bItjx8DjARmnAgLKLkdGfux+4IOYo4AnxEOC680oex7PYqz53tlf+o
/LqFH5WHtjmf1M8aCmnUaDM6xNADw6E/kjOlzVicupC8BSCmMdJ9l148L9f7mmGPbXaIcCTx1Mxl
VRzoglFoa8Ni1QCKomGqST65taXUxOYo4gnZ39NqGKfDb1Xz0DD/hMoQ0wxalWzH+hMh1jwD8zlp
CbZd3Z82BDJy5nIr+QgieTVk8aUH9POGICChxN/N486G2m0uSC3jK/me8MZBoxyF1GPTbYl8Cc9r
+6lkpMX91E44Tpnflmm18Oo1TFW8Wjd0yPtfJUqsfCdnhDqRIK9mjWpVAyATmDZaMpbTsgp3Osyi
qzWb0x+Lj9fvsPDCGYXE5DbyuawvsuQoaS/3tSyHEDmHRDVqpHM9cJjI8i324d3BKpIe9iiCX8i1
LNlPK8D+Dab3ECgCr3mPsot3RASKJ0msT9JWYImQ5IonU4PYdccRKiAANXp1pkLowM24U3CM47OD
N4TobRkKg9Z6uIgfcbbjjdjuQlHADF31EzeuwDswCBenI+eikVcdbvq4e0BDJl501DhFvhBJxoCV
k+1oaLGxCiahsC3Jo7mDH0Wf87YyEIY9xwRso63zdEqRda9fnN2577a3Z7Ci/1GRAnVo5XslR80M
y2mwIOytZHXQNaE49UZc1vovLSSRdmIslIhC0qwn7GeUxJ68M5vC9WCfY/hA5HOwqY3woln9GRLh
t6oc9AX/sJJ+X2/22xYlXXDE7GbTz3460VhUy1aZ9wL/0lPJ4uV5XkoHYeQpa94aucWX5jrbGD5d
/CcQ3sK1K4qCno1Dotd0R0na7ifFlB9RMHYykmQELNnQ6EwgIsteHcqqN2DMGkST/HxJBvtxuN/H
RCZ67pJdue3tTCyN6ykOiokXFDiQRl1LFSMX5uvVw7S3gOYGomMQWABM5r0zdE3J0B2n8Cop6vj0
uY0Pzq6it18O0S5rLVhzhRge8lfXsfCZGuXKETRZ+5UccpcZ3T7PsWPSKAbcxwR9bTQ9KCHFFFXR
2a/G+KJAU+N3h6hSiSo6dOBwbKmBDOuw2EnuCCXelTOJ9prZ7j4PtTzyeDEQuviz6Smb0DeFi2cU
g+NGN8++/lHtkC4XgWJSZtkp0yNVU+Zrn8kYwcq5GtNwymFqTsOGzkTlRbzb5qW1QjhfAe8DrweK
AVTIOEEu0v77MAOvJGQKFJxVncOFu4FZ0NlcaaQ50IKDC59MzWqw3QoV0h+YhF4ao1OOETrtAdK/
LqprRkZmlbj3Nd3Jlv5lr54GNmquQIBB41W8hxucy3mywH2t9y9EINBFU5KP12O/NS60jKJv0K3S
YA0d6f4HDLQbUPHiXqVhRy3YE3uvrcShxLS/3oNXohSOn53aeDoqEaq52ozl3ryvn0SyWBccm4+v
IWmE0PWixEBjjscEqzqFt0vFBxZEn6IKqbic3D7Ar3wY+Ox6usZhUGXLtruyzU5WdcaSCTye+87h
ZgwXS1EhLyvtX76gacw92KmzqqKJ/q7gJf0zi/rAGclWkI3F0I6Uc+NGrpmMi8dnBb7TIV28L3vE
aVNKpnGPYcSIiUfp0KGHKBfZBboTKmHQfCKS86HersMmjv+hN3AYQZWCM6w/nXce86hVsMIiY39M
mVLbtOZaKpRDz6zBJdXDMxeCunSliKDadtP1sSv2Z+DMnNZpnBydcVIHm55HCJXpFQmm62hyB3r5
mOWT9ecMx9VEUqJuTsboNtSuUFyjl1k4nWWPT4RtDVcupHmK4+nxgCZndbTRFCQDFX6aUFzqeRk4
wqJ7MAu18ru7tuCmty9vj6/HrFabjCu44Mc1yyvRhG26WtT/luSFRjmongt/1KwpU2qKpjNMUy5C
3/AAhKiKKaIuc8XWiqpuetNdfx6AwvilOeGQbVJYldedHkTdmWk9GEPssuOFtbCpOACZj8pifwxr
0qqTATovKYxZPVA4j7gpNq7pfHiGhapICAq58bkPX8M/em1HID3PBgsqz//mTTjSRIL3lRHeTpRe
gLfSzR1PTz6OWzgHyRnJ+g0OlyqBgLI5hw0H7p3k0v23gJHp2Tf+DYCDBIZJ/ThabTJQRI9xjLfu
BuWi4ejQLro3BQr5PyCwxUlOHkji29TV1w+F/U85g1/T9Qnq1IvaDB1bxZ7AUB/IDqVtXvz4qmBw
LO7ysA2MAebyaMTKjY3luBASvICrj0ptYMJzMlXmkWh/G4uPuxu4z5q0JzidWh/uYpC8deUXAr+d
nCQFJObkWsvsVJANNo2wlngy4YNdFMgp/9GH6D278oGj4qPps6msf2VEn1ZwbAMw/66YHwoqQgyb
mdiDPFIIzkk1Koe6HxOMwx08OKbwFwARjxJQJMYp2nv7cOI7VwDGT5x+8LeZ0pbSLNk3QxBxeX4q
tzWa2+9YxmFH2tnhX//bLhHwJfVGLJma/fUx1PCb4qNSCjmgRK9PSwwpJFHB4EXdAnvAnVtBqlE2
QuLWcQQhLCKkzVZhoJGRxzPXXN/HFN3gKkiSvgXcJGbRqSTnz8H6LHkysfKmrJjnjUECUTunlGqk
nj/lRFgwpnfjZZfJ6/Wf/8EGoapZlKSly/kLaer+0QaPq2Eenvu0XZjUlY+Ov6J03ONeSqu71Oxm
3nEkMCmMsXxQGcDpHnLzX6EQ3SbWMrBky0xVYuGFh17H9qojDZjCsxGuPdkg/vMHrp98X0nWrNN+
5eWA64MSIkLSRD0oAVxCOQP8rmDhZYgsF3iFlKoKDgtZok2hZh2GG9g3L3LDIu8zW9xPQ/3KHzMY
0jDp24ebvW/THXdiam/I1IVCM8m/L98F8lVXfMJQguQXVEUnRdSwAcAEBMuNUY0Qh2WCjbIs39y+
9Of2IBbFNmdaOb1XAGyEIwKuK+usXGpr/Qodw2XZaYvyS92VCneJPOLW/+rcJA7PwpipXVlXBy96
VpbARVVaK59W64v58GJjqWdw34Ry+OY2WyMP0hEOs1ObuPTM5Tn/5HRdM+SZfukcFM3C87PZ+mpV
4DazoSuYahlFodBRc0DTyVsutIZjOJ0VBS5ld0tlVTYu9PDEUL5psV8IPYDrTPYDE71llTgP11d9
aLN9Pg6oHiM83yqs7p7pEbxzWEyWC4sOxCFZ+wPXDNw+4CR0wXwvnEGSSvHVCAvjImxIgPSFbDhS
FRB3InQgeJEp5yv7/a52+p9bY9dJUvz7CBcLyWGJIOSY7vFLrNbZVVRrOZRL4bckkNv7xdcw26jo
DbbfeXQRozRU6tcPRZZ/G4IP3r7dko6GpldGQEH4F3g3pvOKdLqBCfE4mpTpGdhQQhdGY5uLkAJt
WUBC1QuyjERtEDrgkSqSBzyj7AiI4mJN4+ONGk6tcO1tImFlcrTnLH69H0/+KHF3SFDd3VIJkU94
6uP+s5s6UDVW7u7T2TqRkhhnyDxPzEcNZdi1wvj1dEQQ91RP1AoPTdOfgY/tCAspO1DkImdk7Usa
CF+zub0SuogoDwlG+fG7S2gQ2MF7MMV+wuMUdLgBoEl6726mGk9zGAFbyNFymy9olQdnIwbTSded
Z9T2Nx2hIUXAODW2V6uQRf7D3EqkGROQ5LbmOEZW3K0T3yh8P/VS47lMZrx97j0h4NnipCWzD0yN
M7DO+OtyWA9gETzJ/iPjSSglFvlP4BOinrzrPhqrOiyvOYfYE7EKMJ9WZLVvxha2e4l1oxsA+FBE
KoCOl+ofNTc6CfSv0cCaXrE+Do6Yit3VE8fkaxsO00Smi0akLd8wMkLHF6QCgOk57Lg/EfSMMqVr
nvwe9STHy5i7zZNHvFCE1fUnXRifJnpzAJDnBEzbHlryO4OZ0x4f9qXT7P2LjIPnFptKyoux7lxu
JGcOmeYnwTAlsd9/3WTvlmeNh3Z41fIRxh3XK9WHMhj5+Yr95ZkkBw3uQCdSJL4iXOt4izv8Odcg
rngrZmwPZS/wst3l3HJBaB5YbrxNP+MaHKQL5jmfzeaPbrEio4/vY+ot0ucK3DR44Q6QrUa/c4v1
afYNj+96UhrFnFNjNrXWWL5xQxdjH8gSgDffqAwtAwbBIrldcxGVOHQQW0Lu6uz99xZ+n8cEJQSw
qtwyIvl0Tx6SOGzOZ9tA6MgohdH7mjkWYFAODa2YhRm0NZ5H0wd6kGTkMNShve7OyA5hcLEClVCQ
2pJSiY5WtpXy5ivpijFu+u3WY8nD0M3NAOE+mTsw2SZGSCfsbgSra1CEHhFSvq5r67FR7kHYdgp7
qxafLpDiIuokF3xuihf74VadUuh8qGIFuy/Z1HjzvPlgT5hO+mSo+yX8CQZgq+xNGxcDqUUJPMES
0PoowD2tF3Xdx7yg319QnKom4UBe7/OucnWMgQThlJHMFek1ejAg0h2UF3a8gZN3x5QMv9FRYySc
3zQNFIh/yVQDyJGkAySuyNbhFDrWk+s75dJXECf0ZjIKPZNdv1CVs/9nEf7aXySPzH2k3lkQHQ+P
GX8KChcWa3SZ3avTeXSl++ekDU3N9ACIxTh6AkRUFwMf8me2naQhorHFBXPiZj3GwfNMJjA4Opi5
GFiTpPUPdMuQzFRN7MYdlWxAUfNb1VGFDABBLQ+Lviyl9g3MB46ARE3NNzRqIFKdZMq5T8uxgOO0
rjGKsaaWTAWIQlZInO70a+ntRnzEao9uVc+O3T6V5tp70xnOmY+QVieFdvJ3UDeHYFI64HR+O5m9
dkXxf7FPVScOUEIEXOppCEJALGf1i1pCU7UXKyWrdxesOwV3+2MPwvMmsLXQXPsY9nYyj9+Q6lh+
ScEAI0syx/ogPKU6hVYpRkeff9nTRJ6RRCeqy7Duzt+PtJRT/BvRii1C25nwSzOqsKlD8gU5ngUK
TDaNfjel8YxuzlzCn+CxwueKliNiFdLIZJRLG0TZNZyhVaT5W1MfaPMoA9X5USdtfb2tO3G0fSJv
R/4/g6kRz6GPVrKCri3DCq0fIA9h4ak1u+UCF3x8XMhy3Z9rNnt3JtUBA1AXIAXdf4FJUAhG5fXZ
9d6oDL2k8rIvF2c2MV3iV4Rn5NEj7hQf1cg5FkrI2kzx1g++BQkWBIvrD7uvswNrbAqO1MiNZkdY
c13cf7uHLmvYS0wkMDAu6H/vx7CrBvJXy7EGDRVD4Vv8tn/IDKT/b2oT+JVVRsEq35STIYm6lzRF
15wZlIshdWL7sDym5e8T7Tt0ooN53ASLmUY43L3JC8nCh5lvHEvIjaB9RapxB/g1G9p8Qw+hfCTj
NrCT4FfknEIujLV7OFw7BRZSh6UEnNRfcEPmgQjO784pskDOOlHQ8O+0V5u7n3jIpzXIIqLkmpEW
hm8KmbOW++DvH6YQ4lgNReewEUc7okmDGjriH8vJpfDl94eFjUDHGNVSGPjbQg9tnQwjMOL4MgOl
ptJuFp/qxuj4SD0KkdJugdpySRz9pThbU910uv6VXWyhBvpQ6cvIu2SsHd8eGMzLC1xbRdgTAoHe
mxdKYc44zwxiB5xAkkJMdxDNqhNTadECaGWl4LjA3lbNlN/u0XX8FSFHb1eRpy1J75kdLqg0Ya8+
ONoTxZWlUee7dqPkCwiMb63KFa4c5rsk7sb9S4UMfqb1mR5R1eo4kKDH4s47AihRegR6ByWhUyle
ZGMjdesFyCiQH34I3KNV45PNC/YROFC7JwXWc13EuHl00nbtmBr1tAoapnyVimDamtezm2kF0w3N
gOhY5gl+91gd+X4OUCxfSdPM7p+p/O5xFbRm2MT7Jd8QJ/qzLP39CgsfpJt2qnA87kkakMwpw3NA
rC258JdnZX3fWn6CS2dA15i0T71iY2j/teNFQ/3BmwQprvxm4rpn6vY0bWIn2RQf9Es8nmzBIV0l
RvYzrzrGka6sUY+8Qy10veWNC4cwaCWrbckiE5LYPyjoWK31r+tixJDsnc3VJ7xz5MdZhWFyvgpu
7HWYM+KaXVkfZrVt3CPv8rbJgwyb04pyBZYMYu/5TjYvVpa5vDx7eswzBONWKtREXmAByi7CeXYF
KQx8y1ebLB/qT0BMplQy/wBcSRN6eiY/PCuOTBCV4sEe0uZ+PtNHGoC8BoGMcyX8dBmHlRjOxxVA
pkdiTYGNpdL/AcjrovfjgbBduqBvbpHRzzqHdrLNrLFuAHL9jI0JJ7kBm1j5quGD/1kPZf8Vqzpt
K8kj02Vi6gEEv2MK3LY6l5uNhDzfuGflZNAQb+YcUwwmpxRiN2NdmkWuQ/gHywcjLbI4REA3u9J4
G43jut8X+svRSFuuU54vuKWO8t7C9UrKz1HZm/KxUEujMO0ny1vPO9qLTrwv9KA5rDkousiNvYMg
EmkRiwkzTASFzBnEPERq1A3Ylf8rTekZYTqPkLDKCKa7M9jZyIlHWKgjAO3k9dlgOk6o6yvRG1Dj
8CinOZnlww9I/WF9HNoLuuTWn+4XgXvO6cdJWooUWBerldmHCaUCnB/3aSGHyo81QyBEmaIzR4Nt
R3x5/dtzFuvLa/syeKLAWhXGgWwv4fC3vhITL/+MvmH4Mhg50A3fg7Btn/sAIxUyVZdVRpAFP3i4
uh80ObirBFSkWui6zMH+pLqh5AfbwmRYXGffEnQf6qwbhwcb9aMds4PsxJHICDfoXhU9nWw4rLcV
EYRWN4+dVS+EAPWPk+TErpyLxptBtdFjRFGPrOYObuQDRrgDqyYAlf3EB6GO6wmuCaqqDCh/zZqk
ri3YEZz3tjT5sS02QTZvlCrH7p98fT3VNloOJ0JRf51Sz6SdVsl13fSxnZVPuw0785A5nM0cB3fY
HJnnn6wU0xXL3N15n1uFWMBVTEbTTXmdOuQ1rdRW7FHqi31YWbEgiJkZiJWwjRLdkop6Nzv9xx+l
zCoKZT2oXHP9y/FKTr70M3tPI9KEyANi1PB0tKnKg2A31VT8DpjLj52N9wTKcWGr/5EYKLI3WLc5
qEfvGBxrEM91CLuZgP/JHU4wjBGgpYMQSa9pk7PQXinkEZwT7jQbo9xt+cgH1TftbL7xFw6jNlMu
noPBLL5gCBUXw1s3TGiVsvfxtBvK13IAzDE6WkTBSE9y7EU1EdLy4wjuFb8d2cd3GM+rPBPPm1un
sk3imUw7tHyiEC8czohbrLXFYRRfwG5lqX01JX/Z1i4Ds8AbeCOnuAbiIBHBAqDZxEwr7xXmmDxH
fP2n/cWbIWZuUvruT+LWzF/Ek37NB8h+r68MqYIX/FqfK+7fRDUUkmoUlwZUuqh8nYecuRtfkQiz
U9stDXvC68I1BmKGR1Z7rvPlgLc4a1w1t/4aFytiSl5sqk9EbOSX27zy4o2OVgAhlim+qkSFN+SX
RUL6nbKC9OAr9Ts1g/Lj7E0vz23izmfeN4g4dt25ZeI13Lr/QjP/hkBBkR6ovkxsKBvCG1HTwrMD
UvkJ976qJSwBVsmcGq25+X/CQSdqEJJLMykgqDWP2te24MtSGDbboQBunGyAGgABRZCwHI3+boaJ
UFj7FXL15AVSOOq/6w0Tk16gEG7GjcE47CBb3ncfAXNgzwW+EgElEuMMXyy/l49DWjXR4xy2zhkw
1QGpg1eWkdKwh9XrHMgyylULISWUuso2/+T/F8R7/0K7zEzlRSgimzZzOrX+GE8j3QbVL4k1XNNV
nM84mma0zN1QmYpmJpbYrawnk15Yj/kycT5+WBHirbgzIhlCfnWO9iM/9EH2NS4S/OUYtQOkfucW
J2C8igA+chUvPUEcnfjbZEX1TsZ/4MBTkg6SPQUtaM2G3SHiRrKwc5j2gCoMfRW7ocJQbDvJfWNm
8yueeApcNU1MtEqAGlmnuP8TfSbYTaZhNcxIRCo+1ew0w0opJISZU+HkgB/y7a8kDgxHfY7LgAjJ
7pmwkFfzyz8/zfmEodx3dq5i8VgW1KW8cbcNE6Ae62tyRHpmaKP6dpVAR5VSiXQZNwk/IQ1nYItT
clmd90Jiz9m9wYXqbnR4DZLkmwyckh4TkISMovidW46w1HhCoLPAgI9BEX8Fs6+68UJiXzQmP/Yy
TnI687aWBwt7gKk5kn5La36fqXAOKv6WGuDj5ZdQzg5bVAj5ZFleqlG0SU28437iANImcJuVB4KR
KiEOdya5x9dVAvcNwRvnnP9lsBquf/v+OHnvdf4jx1hZXzT4vQxAV8yP3My5QsBY0Hd7rYYcZQHW
XT1ixPcV6JutjO8rYfe5aohIOVU9C+B90rBCC+ixSZHhN6R5uM9UGOmcjyrahLAiRu6Yokd4+nRI
mSQpB2miChrOYL74pxB0EcY3acng06NfMVh300I9P5Te+cg7QnOk9lQUx2R+7LJcTht49I3asLNh
ZHgM3CgiciT4RQFiq1RUY9DVLUG+OaIxjOXaQmfIrjPWM1fWcOpRJT4YdjkSesIm3aVEK4aFiN0D
c6VJdL5jeSxhBzr+g15jny3dMpJG6TKvAoCym83b8cMguMjGFoyrLC6n7d2IiKwvbq2sk5TCWW8N
zkKmUWdFKTVibOaOs2rwM647SRdAQcmYTcQA8OA39ouIlbKmyaUgJAJ4eyqs0gKXwxezdyBrVKkR
kUFHOSPvvHqZxLYOgYt7HE2InxqAKKpELqDkN7N1OuYuFpFyQi2clWQk0eHG/twUqB7aaot5qwpi
Lh5Sb04dKfI7Q0HoAErjtSv4+NkI/XfcYI/TEkGrUOLNYi8MLhxh5fLiw3/FtriWUHQOLIjsARPs
1ejSmDukTPt2iH7CuqoVuqBeTFAjqGBIqEGEqZa9mU6e98hw3EdpROl4ExMF6fhOc2JW0mT31+kG
aSstX23VHrFhOPqew4PUwvs6viMEh7CiF8tuRRAn5hXemMH4eiz5odPoTHjhjKNiiY1KkK8qnT2R
btA5hQD4hzRmxApNsq/TKe2zeqgAl+htiHo6O8r031jAf+wfa+wHKhafj5ETCiomSR54YYtrHaPD
nKGzJDQhgBd9gfg+gxB+9y/OlU/+4Q20SX0AawHgshtwDblwV/EEqzU2ASI5WLdJIZBiWldrrpcE
Fjyl8yEkQofkDX2Kz8l7TATDX39bTs69n3BunYtvBGTt3Vq5vh3c2CLXPn2x9zrpRs4lG5vSqSDh
EXmGIElQrKj57JHO+Zd4llnEpLQf/p1+qwY9K3HcjAF2Ms/EwCkMC5k42Lv5qJ0MjJDFzc4NNICs
Koh+19GtMeHjjzKgUBHFlPisAG1IcoBBAKlOy4mrrRgFvMMu3axOIBN9RDfUsMafzzrSg51pR7UE
HxOe6/9bZ57xx0NT8OR2ESZo8BxSnBLR6b43R2CpD3/79VXhpTeT+99lIgYQ4RlYk0hxgU34LHQv
W21sXgmw3yzGowIR73yyMF/IZ5Dx7TiE+9xakih8zHyyHYJYW7AT26riODg1VhlqkUJPg7pL6uNy
Cue+mMN4tlIAgQv89qhsGMrVI52usaG3J3ONqlm63fqcNP5mpUKYk0Bfe5tQkD7L9nGm250uKUXO
G83ESweL18pp+0X/AHME0IjgAZl2t4qiSlraJMqEB4VXswuAZcz54LJUY1MNKez3Vj80SXnTEx6u
BknDcNDGJm+7t0OrqMl+DJt/746BIkNDLUq0CB1LPZXWI8+vJMEO7D5dzGke7a7H64tTUt71jkv0
ua0w4VWfFAaH9/FjchPFETH8MJqnaslQVO1xdVJOx3Y0sC9MfuvKKv7Cao0qzXAPIH7OjqkaZNyt
7ymgpGj0+n6RYaDc7j4qmk9tnXHbxR/XIupOnq9xE4hqohO/POfLF8IT9+j5sU7r3qXtbJOyKcKz
MMjTY67fh2ZPYYErfhq0/bsC07+qXV0+/hpjoVYfnQkkrjqhjAlu1Q/PGQVU06wD5HC30u7H12sy
g+9CswLDSKF+Lfgb0lKqPC4TWqPQP7izIALGQkbWdH7+3h3zKcNmqUaP/SuyNzl5ExbDA53CokNB
3WD2K7+or7LIOMMyUpFwrM1mmeHmwCH1mFUKwRgcbIXfv5KqtfK0obLmMi2/ir/hR/kLLMXPnWOO
SS0zmlxniSdIAMC384ttiq/z3gvygvTtdGTHBmM15DbfkcG1WV/fShHMrbdaoTfDcLgksw9cX1CV
yDl8APbETDGK0pEG3C88bwG5lmZBo7uXNHuEiW/Yec8taGz++fU/TuuxjD2j4nuRh3StmDlVOKrJ
yQ8zXMMYl9DIu3aY/1E+9OomL2vU3J66AxiUYv/pq2ePdhz3fWVABm1mdBjtOnlw9WFgwsqXl8l8
M8VZ3QO+denDJvqGayLmkj8eIoxL982uD49DXMn/A521r27Fz12TDuZc+6Hr9zZGLLq68o8sh97s
UnbFnE9nr5z1jFxEafkNpV7cMMJ5u8LBUi37Ae7sb8HJwJbUWNxHVoy9Se40lRjXid+1ZZnvju+A
yKAIeFPgIgJ+Buc4fOlh/zXe+MzpF4kro58R3gnE2JeyDXE2vNkxv7Qwq2nY7gwtMiqBtEGjte/p
sFjsOpVLA0MQsCPLOCC7u5+KgP0oVYZ5PcJ5yMKDolmyYjtA8vUra1YTS7pij2yv4B4PAP1AP+JN
Xx3m0k4s5HpXrYmJXt/xTZsQvMUfAeHoqkQT+wgs5f1dZKaw7VOM49uMAlstWTpFxcQ9yR5XXnb0
PjxfTi2ToW+M+ubwb+q7Ko66WeMckHrP0Qif8smbQx0dxARUjmhPUCvWAW2FsIRbYKMlMyQd8g8M
gfXL+2kmF+5iJPByh38x4w4NVcQGTrLxC7F3CfdnQryxR5mSXYjBsFPg8DQ+CC4VgEzKJbeTRLOx
Uk0fDzqVt2VIsyb8xpKh2tS3aSGpr20nAmPBsUPzz3Q/aPwbqvdxZ+tsHW1rL3yqVc2D5m8NJWrD
uDz9qjJjIIVAB5ipS0rTLClVISraCmIHq3P2whD5Xv1i+e7pn8SfFkfvwL7rIvWw84PikU400U8d
tFyNFqtFiyOqzoB5SFI0Id6wXA20jtVgb9lfmc0JQNLy/1dDfHMUHRQTi8/6P6ypUNw+rCzroqVT
n/KZk4tTED4hvIX/mN+F8SqQ0MA5/EuA20je6GbL8wBzJl6NkHaAx1ynMY3zIgBKBNxTUYQ3/VHw
LDG9cFnZ4wtGTxK9wNt4i8JC+c0Vd96Aw0aJb5OWNQp4VJRiPggahoKUXvXe5ArNaD2rKXpIeoZ9
IJe76eSNRqYjajL1QMb7NTcM6KpLc9qTtQUElgR0FinHMCq/02+DrLNnBDkl3+Hp9gtPC2XAF0ak
bMkfNTyqFkn4aPlETzVcdgeaKgK21Uaglb5RSZsPAvObua6hNkLjoWlIFDSZc01sboSTmfkSDe8S
AU+tRm/wuofJaMEIf7KQ/HHNwevhaJRUP148vWB+o4R9UiW8WFJA+w7/thTno62agzv4itka/h1y
bhNpWhl0W++2KlHRbhzUV8YJep0n+pzQ0H4j23k6DmUcnHbSC3Bdsez7iW0X5VDfpSPYcz4NGLX7
EZXuSnp+1SPCWyGEFt4vPbdzXZ5j3hJvPGSzaJHAnHttjxh2ZjXSepWJCPNPxR+2xOR8YHRVHYC3
mdIArj1buBraJITzMa/wPQYaqZ8ZRGitBcHdUtCiGY3yapRf+xXbHHWCiMofP6UzkRUjixBJFdbq
2v3eazdXW7F6o0MR/FRLshLrOPEm0xOU0hTRzEBJRdiGQDC3jsbW8NMgCWxCEEERiWyrtK1w5wDk
8G0zPY1lzA97xsCIrb2v1xO/Ki8XB603hx5mksC0Ia+9vXBd10/F96RfN22PIQerRcPndL8k2TMr
ZsyGxAk06GDPNp5Ct6Lk7Y7tfZo9ZeJjzI8OuSoB/kawMfXB/kSzBoA89dcnK3nnmIlx0Qg1ZwPN
nAC5WgW1VJYAZQsXdUnQOoYNXIKDuBX6+LcqDzekNWEatA3j547dtlNJ8PfkHqScjo1+MMpES89p
BeKAXGTdtMLiwC0VBbVCfJS4aEkyilanV1y0NUuhY7PajPjDNB01viJjk1+KarkSDJfHez883N35
yn4MidPHrG23JNre1kWZf7KtR41hh0ZtY3PmjWrsg1vHF1o92Xql0fofzmjF9iHjLu8mgriKPEbL
2Qq0zsm3awqmERWUY7ozpFLMU9s30MLOLyPc9FOllnq4BE/ONxIRn39bZUomSw+csH6c/GE0dpN+
w/9fNhVuPXSeS84nGERx8gACKUeyxNMlhu4ujg8sBJrTnnfUp54TvI00xoWsXQm4kd9Kn+MednJl
a+n9/aixRdF74edeCBz8ISPGjYzglR/kMeuNqSW+kBEI83p3Kz7z8EazjDjJf9HUGBId6lKDqKVL
mHYyQUSRT1dJXN54fQubFK6sJKynnSOgIBct+k+IKd9G51iK5I8Jj0NITtO/NJZpnAxCBaZfKG/I
HT0dPZ4p07uHzQd4HLgOS46o3IgjgxoS1j5/K2MB7BrAI83W3+YDLyfyxyOYBOEcZQEC3V2N23KX
1afOJjQ42aMtaw9cZmAKd3x/SycJG1VwvwEbsUvyCPCC51av0ZFPkEeImyruY11FRyH8S0JX8zQ1
RCfNK8nj7NX8+TdPbC3HAv5HeQBaPw+uPVRASkTTh4vBfsjNf3SAJXqNGh1O/PFZrYywzgCTVzdj
Zj0xR4pM2d4Vwwt1fPUtBIGY9RILHIjRDo4eD7hz7AmP6pfCJxsu/0g8KYchy/ZDUKXMKG0hf6Nn
LyhHIN5Pqp/IONhs26VbkFOZ5SwelOJKNj8PYXYT4ETiqfULVwvKk4WyTdQScqxmPOKUcTD8+z1g
sBp0hzwFGenDEi8z+WvfSIUhUkdzt59Jmi2t7TAgsfgzne3PQs7ZdBFq62+mA/9PvrrsuNolktsQ
JSm/w2K1geuRpEmHy6xifVcp6izLnigQRdu5amNtKxpU0TZILra82L4HVKw+JFljXGVjjxC4kUMY
mWauhvC4CZu2AvoWyOAzTFMoGS+bmQOcrY54hL08RsYjQUR6mUsCd74/7CfwHTzk59yCEhKRsbP0
ukP6mINXhHQx/ez6IWCkwdyfYxMxl4dvSDnTYEO8hz8c6tNJU3Yi8rP31se6awLek97g/qZSEJcu
e1+hwKgxBJHIWhvyPr13LAZ6R5xtNUlGLNRaXJ6BlT6sXT+ZAiIrK4ZV+QK5j7yjgr51ZyagjcYk
8Y+HVQxe9sDt/pbFSljnyslYIxCxYm2S+miEOq2jPZn4dc8Vn7l3LUBBtK7j1O8X6xsZNdtsSJkz
VP2jRO5uF2K/Kag56r2CSlkbPbiHGXKCni9ySFR3m7mjQ7RzBi9FjrVWPHI4j6+elRRUUKkAh6Fw
he/YfF9CCqPy10SbCAHa0RpQWrvfH45lWiy9b2ekOB/q+vdxZb49uKVWLeCMHnYMVQLreJFF+m5H
JnvAS6qvBeGm5hygZ9HO8djZBMqh30CRVQHj/2nT0KLO4NrjlOl3X6tW2B/4mHR2aw0zG6aMBJzW
YFno6EX5gIx2Db9i8xSIQ6e8iKFP+h/lXi1ztUHv7UAQNvReonC6jm2MIsTDFsT5hdevHWthA1pf
C+xlBqeEKPBKfMsJ+8FkVuAiHUX2SlEv3Chg0zDuWZN3ZYHYiqSDgtgzoPNkShbh4KaFssAD/81a
AOrJTN1K/OuYNK4znR8R+/JtGIaxpguUoS9TNGB6jCApvmTmtrjbz1ZrMD+I90gm8zyHx3JujAde
QQd55ZVPZCteeRRIEbbIWkF0OV5VKbcUM3zEG9Kto0ZYupb/NUXMBCyGiVfkXyuas7VU2yEH3udn
csVw+4sErdHubhCMoldldB/dyMIgRPzOgreHs6WNvUE3FZNF/jzTiYDhn5+jjNDFgg91HEM7Mrmu
WkpNNKN/Israhg0KLm04kt3IVnER75ImvBQxajbUejD2GA68WHia/4lGUFPfaX8k4JM/mhIB0fnZ
s4WrhwTSVjgHFhz89KjcglDoC3x6IfLgH9R4C1cEvk7kpHCD73RIadvUjg30l/0vXpc5RwPFCQbZ
WxGIloVPNcotpxKTTSWkKozM2e1TW5s6ksc42GeT1hQpLDC07ezGzuOk2nmQsW92d1OXz4FbM4YJ
Cbe+TDAJYoLKj/vvLdrrT7rglC7enftrat7EWcRfH9K/JDVjxNQQySrFkPT0I7ioeMLprTb1i/Yh
xpV39saNXnzsblk5iZcAPKslPdquPaFBuLM+sXQyNTo9ecHwn9E0J9LrhEHGD8YpvQPPgp38jbnT
MWHxD4TKdanXcPCtfO8und2vidWuGwmd9GW15lDqQTCiKuy+gz2hnPRiy27YMSD4F3tCSfszIT7L
B9320eVtW92MfJ0NbkeM2BjevuMwlVQQE39bxt0ZW8PdGsvjJIbpyPBUoodCKg+VxR931DdqYiPY
BEd6LjWXbKvapKNy68XHbJM+Eph1ZqXI9cm8li2UBLsoq2SKyyxNOdMap1hrGWQ7+4fFPQ7JQZMQ
v3aNqLjvFhaQNWNuc1Y/kM9iHmD4cwJMIaQ1AJYE0hQuYzVWw71p5mQPKPgGutb0E8/fxFr/f+YS
OOxHZQoVY4CwEgBaw36SRRPBmtJlrOYLx3RqgIK4BP6io+O3ma3Jn/GRzeRMbdgQncjafN/nBEu4
DQvMrXstex5BaMo5Q6WYCRMA0+wYR1ZeHaQXYIjhJ/CdTAHYMCw/tNB/x3C/iAl3g2JszJdbliDh
f1CXiAIj+7YJ9uSBwnQSXNaiLGnnW7Rm9fVXMt4361rfUEBTzNsrHp4HaTzLdMRwfJLwkH6dqq+P
6c2IcGDwy0nKvKOPM7scnNmWxo7XsYjAc3AaZaRW0quYo+CP+inmzxQ5aPT3M5ise+PyH4DJeHkS
1jJQHk2D10O3H5zR8u/0Dk8FnLkW6hkEI9wL6c4zO+0DDAsQouljL0ObyXTbp5+QYOvpcTpphg2J
Y+ug+nEZ5lOLB/chzWECh3nwg09lz6PNOe+OSX01RmbokFssf9lSCtX6jDmMs8DzF4hrU1i9IyND
sDZwH+IupRx8373pgf6HggVPtPPs4uTMNX9+5odCYhtmvglAAXbSWN9T6vNlenvegFsEqWDTjmGL
oIPmMLzKi55+V2Jaktc7PIMFRegU3BaMcweN12jrDzxyhFDJufMrVaSE5SZ/ocXhAc9fjlDGvRA/
MuaMD4Gx4HDBDxBOiIrpHv9XjSKyxnWluoHewVFRWyIBkRMF0Uu7Y0ZLlUvWjroh7+cIGp5so+HL
Ep3BLB1o4nIsydYuA1VtIdmtTskFR2fKvGCwN+zRgab89KKTC6qhiVoct0P0oX+NT77/KFontLxd
qBmWRt141U0y9NRCOhUps7RWFEjMcyN+Kt4N2Tv0xBHUIvS18YGyqD5WMq9CJ4ON2MobypOe0GKc
SItlhF7MFEvM/VyOl/RZ0hE6kV1Ie/1ibzOM/PNXkf4vZa1oCc/DsyRyqJECji+5IkKDyG34F4CC
1WT4vqK3RTaWFp4QRoZLKMJhALibI8uPzFLBz5TtEsCQHWZIe90BQWYR4u+Yr31xPBNmwaHfEpUT
hCIGncfIc1MBmr+9OCxx4QUaycjhyxWxOcuaFfunmxzzbh6KsWAa08fvueqVID7Dr+EXts9ls/Vm
SKvDYwrmDtwLWS8xA/Re6f0rvjx0qY9JWTprv3ig5BQVURa2Ivigrp9b4bb2eO7Xt3Jy3pcKXwAr
BuAUTydoS1tub8rhSXqf52AfmKEKdnabUqGcfOlVrfVB+GXKMsqSnBQ1UjtRp63LNwi362WRMjGY
VZq2yyedHdf4Mou4jlG3odr7JMb+BtWB8YE3TQhE1aaPs8+rPgFUmB8z8jMcA84stZpgCAQtYl1X
t3zxWNhPKwg3ci50eoscjAUPP4GH2L7H67iz24eW2VePQB0pZDuOaX6oxVYziO6lEyYQ7fc3353q
2FDci43yUj83Xssdel8YB2germ1i0hOuHM7AwyRybNO53tBOCIuMd4OxzujaQKdAMCYfp+6shk4u
n8rnzSMDx5FnrXFhm/dTac/txgD+I4qYm7X9QE0azGaJXG1ROsVscm4cv2ipDRe0smfdp4Pjliq6
Hm1Ps5Yu8Z+PoNOAZV0t9nVk9LY9bFlmJXLgnswuNEGL+iFyVBXR5qEMbyc7QSw+BABx7egylvLI
dIPvR3cPbLqBeXMLhhRpqlCh10Jw0HqODh20/jyCWkl3/eXlrNHKTOd7p9cDD0DmC4OiednHbqgr
2GY/dEOSIR2F1xaQrcN8a3yoo7VWRKie+5m6thFdhzIFWGNTE6xcEma7wUWm+OlUyGrwd9XO5bK0
XF+4htA/LCwNLHNv1+iyve6o7y/Qi+cMI8dQZ8NYBzt34JLXnON50ELyN7rRGZ2ZsdtrLNw6MYYS
VaS1ZetT4KzNyhJfk/VHv6CKDd28T05onoIXLhsl0iK1FCt1WJ1Y2s7ygyHFRE1AH1VK03uyE9jk
F2902xoteKaO5owriFp1+rllKBP86pAqGPLQE4Zowqv4lAC0nBAF4WWL1TNYEkLT85Vo/JgJ49Aw
NW0IV/WA/QGKLzaDK0FM9XKanAOzU1VXVu+ASlbPmaker0LD0P4vQ2dYVmZEqDjkOe9mFHPki6fK
3/+xEKrp7wZXIiTjh6uxRbIUj9P3TcSHKzrDy8ibmwNnmmVXD6wWFhbQz7jt8pGfqMaw7cYYAji2
xPC72/qKQ/6y0TPLaeUtCfF4fOwrKqsmLdW0Ywfv8jrOyJrF7P/PSBPRuhpAv5e7s6dFjIXPtwqM
OWEkHSFpa7zzZiodQ05zBjvD/XtEAMeXz2F4FJNBZNl+d/OTX+Rm4HQqKEgpKwr3+KU+gc5nT+M/
i/TpKKj5hK2dRUSF+TD36E4l/r3Tz3umLbKZWaTOhwT4zHxMGHdJnKJoH+HckO+tVS9DEeIl6Zzc
qLbP1gUdlnTAUm/p3dzMp++VeWrgh568i+iVjjlb7KU8KTQl3DHI/bKr9rtAh6i6Mn2t1raLqule
brKdaCH0gIrNFqatZSZyZDHxZy8RYfK6EuOtTUgGswPeiIevtTJK4apjjjkRCLLRPya+PPfSab2V
v9dDmcMD+Me7jW1+EPNzSTl8WaKISeQqYktc+r8LITORizebgdm5AWfav5SVVEMEjHrysIswnsqR
3i4iGjSOrGQ/ewJCVz/UJ71NhwMsitzGx5Y10q9gLz0UZYDOD14R4mH9WY6M02VahNBsRUsTdEbP
rQi0RAF+V92wkJ7EI6FmWd17eVX65T67SAAhw2FPyMWDEiwGn+9rxluSLC5ETKjHldrHzq6yaiWn
8QblWY/DTwfbx7jKvSE2/YnPd8CdZtNNGCXHa3FjY8DbFE0HunRnJ2m96Bzk58CXq1YybinS3HwZ
xVaMKUSBD/PDhj3r1/TWTu1NMzCRZiXOl4GdmeZ1d5pC5yxQdu4bZAz2sYSkrOwNnLjopjSpfJy9
o8xWjnB4NyWgGECsyCiQTtQxcd6jVuulAlSBh06WB823GLil1M816Ec5zhRoXSITJJcKYm5VYZfb
OyufczaTd7qajfkmXM2KEfSla0DfCkmo1vwXvhmGRlhILTwrtO3t63mKH/cAUiKbx4LNDe9K8r2J
iJj89r5S8aixpfggqlEsYC8KEkNuF/cnTpc6iubOPY2QpXLSAblIzjbmE6w4gnb1YEy/y4DvDBA8
bpP0eQw7Zt9rbi29Mbjl1K8DltsBwXAOSfbOwCf8IxTlnuI99VSRyKCBwVB8VlNgNhlMzvJwncoo
8Nj72rONlVOFh0Pkld4RxGhmnLrX2aR48xUbVh5oqfTVhiSYugNgZkDxLk9cue+w/gRfWBAgBIue
5mrk6luszJp/Rai40c0hhOvdhq90qVKNGPsR6v4Et+Lah+K2cjongNRsjG7O73xZXqNaNlHSH5gw
75R4MDYPeqYcQyLRgI7iww3g3C7qoOSTL4qiI2VPnL+HR7XZtdcgKp6L7tKH90n9kbv9v3nD/LH2
FQ7SMR/HiLGeANRLh1lP98qaRqV9G6mAKvUaXm9vOwiorcWKDBWi+LBEqg9dr7FsV1GoqEk7FdbV
wxO+QdML3Qw5wYdwzVA0GpUmzE46uRQLvxPwb3bK8Bhqzhl18L22nNTAVLCkLo5dxuftWxyupcWC
0JrYFcL+dUfde0MG39Hfiw/g4zNOYlP4iyARfdL7lmTSAn8qWhC+IvVdgUmkaEfqCxq6wSU2QVyy
0gmIa8sR2iesyrtqgQiTO+5pcA4yfGXA8OVLDdu5ny4BtlZBfdUUVqJ/LeaTR+PMdS87/lKhG+Kv
4De/QWRXkQTEO0loCTS0lZE2FWaxsUE/Hj515VsyzVyOzVYqm8iDrHUtVgfX50S85eB2r9Ba5faH
aX/YmnChFj+K+C42jf9U0FZqQqcOU36pMfYax+cCQBGHiYoVS89Fy2VTKjveIKjgGx/d4MIe8IoC
qV6EgeXR0h63+sjpoaNBsniAMogOw5mojvkMffbKhU5yo22dNpBs/CUI9qD2BoC8BWTi18eCklwI
HPaqb8gzSEof/PxjmmTT6pIkgwQFTRIr3TTEjnfFHzn0Z2CFy+qTxA7V1yKfhqxRC/cMlph7XqrT
37FLxc59LF9+YN3ys1rSR9L5zWl1v9D17U91st8NS7KE2pIWlFBqCK6vyOWmY+Mhw8pZTxtd5qEu
/xpGpYg42fBrb6A/DJamSGbWGBaIRrUQK7dosel6eJstM5ylzPJ9C0nbuJIiocFDbrhhJ774mNKB
KXIIZwOCyNdoTDBOtrbnqRDgCFK5owLRUED2PxXglgqz8RNlRQVq3IdJDfNmWJRA7cw9SF5rHxt6
vT74DVzMF+9d0FCOGj1gTmgUr+XiY0mQSC057JFgY1BoKIOzHVlv6WDXM47xIsirZeJOcsKf6A8Z
RG43hDCnjbqdNG0kzqemIAWkm/aKtqLGOl93JJS9Lwp5v65vGcOKPGn2trsbtTYazPQfPIiY6z6K
Ceu+bxaVNLSzvKMV7ioTEJEAHtdbzyzTXq5Imkmc6QyoMpUdktG/KrhqzQlGiEaqb/M0PynlvEYZ
Ks3/M2FZCZO7zAeyenfAK2/t3zOLF83sX9JJyHnmHy/K+/j3Rbi6CJeq3whKYmaTY4RXGi73F2Lp
Ko13XGyQxFa0eiGg0LRVa54D+xZblUnSjUZcQNPOo0nghVCr18b9GONg2EYcsOnFnYMaqIqflizs
TjpRUtq5r8ZbL2wPLiFTj9R7GraG69gGglIlAkXT5M4+VWKUL38rcPY7kz/l8ClpXWLW5yNsw04D
B7iKnuJBmXHaVjbAxv29Pokwi/DYOwQLVOLlnOr3DMPnq1oO2J1wk+doAi8sV1qWM0CzZAQYRr3j
Bn4YSGLMI8+Khp2gNh71BDCdI9X/0o/hhclNw9iaRGatZz/lynBpk0jEihcxyCImS2ZAzJ/QabKE
t7XPZ1mQnNYOKzDCn3Y9rLfUK5w1zEUpOdDthQq9c1qZQyeQEBtLYt7qsZszLLCAWEdPGYuqNeVr
Nt7dtQM413gTeGIt+ZT53/ifNX50w5ytPDMuiA3EaSr3goX8jvZKmPOeCEsZzqID/sCiWrkSQLt3
D9034fzWyyxLBC2GoYXuqvY3wK28K/XSmtiNNIQ3ssep6TpWyzV4F2JgqDjgRg3JCabtf8rGnJno
FNOXFhrw7UeACxQ0KEiIszZSSAVoVmlzCe2R4AKKFG03ynKAGHffX0Y7Xc701Ni79dP0js7qOjDp
JFNcxEDSsusO6l4eohFMZmFbjT9+Mg9Aq5nkNNUOYpK0D/yLdw3duQr8X70v9EHUWuwRjNilrbLt
A0vAhbLr2ss5BuZlZ0U1pwkMheUVFlwtpn8EUljBUUNzi4ErhiJRNSMV0ZyZ7YzLnpxEGRqtG4b5
fSVVQAy8UxLFQGk5kJJ7kLqAiOAn52FZmGC8yO640FwBx/mOaTD7DOMik3Ea/e9McOey6VKH/604
aRc2HTYaTocJg4i3AY5HMGw8ETQP1hlYzqhiZIREWVzkzOqsbEp64otf/4hJV38OFcfrU+KPRDGU
BQaWdITBGWITY5x68hOz7J2sY4+DXPwove3jmvpZWL44/umgihWW4gAYlzYuCQSWYd40Pjc11ZOd
cRtuCynkH+5wr+xQf670+AhxUwCIlt9C2Usq9HPlmvuD2qyZpMeufMO1ixA0vj/djpWI9Zx30ZSA
SMtpCCkfwWqirltUbMGzEgyOvN/EGiYmbGcKHNbC4izavbFWp1pPz0pbEuuBiVWMrz9dRZMmtAZ/
Yq64jdDlQU2NEKdFJx/HeHA8QCeDnpRaJ9Nom62hPWfbWZj11UbVJSzLmiMIi1TW2VWYNNt+VwOw
JASMMAWtUOHPfNv3MKrD3WY4PB+E+lYTCe2Yf4TaqKgTjmu9kzbWLM1/S6Mcy2YSk3JubyjuPMcz
tAv9SAKr3y4y/HTJIcxnyhKE+qqcftpbWLfvTyVhpQpkU+JXkpDsGPdL72CFYZsOhcnh4/UYWAG5
wzi0tbuFPAF83ePFrBIfoL+XwchaLwF/AFUJ7/t1gAC5EgjeO3cs9DE6r9P/Jdu3gS/9v/FuCnXn
hNmXKkdaO844pA+9b24D4a9jNQ+hPRoCqv5yoyW/pg1PEWmEFdPWQGvyrCmJ5eGvcClPqmkZ9WwQ
C5H6Cfn17BpFF5VnnhurgRCi/4DcmhElP+ck1HLNSOi8wuK+xSPYoLpUmsdersKW0Iq1bQxzNByF
Y93VzJOscC7WkpWJDJs8hJpSnqSjRghLRaiGWHiEvJd+Fky8SBJwyKkd3pDT5QIF15YL0kSl4L4z
fQpnV9gO2n2OKbeFKTm9IPySOfyUPzUbRSHWfHKY6/ajsrFGQpTjihQdTVd3E23ROUVmVdCBVuaV
ezlkog6OxzJjWY3vREZxocCOSae7NNbgzoYWnP48pOOxSv8dus3PHszXyT5BUPJtvjE6huC5Qmc/
dGMIlzgPCuHmUQjei6QR+uIXEIfIfyS5ochGLLmbSBFUI7m9plNMuVFvS2GNXiHBwyNE8lhTAj2I
7dVKnQMr6vfIWyqGzXcMcVsPrvRx6M4utDjqrK7nwwXBSBhYz63Cwq4BnJj22lYgENtTkVZ/+hXa
DSO8BjTgGcG6QXFOUVAeYSgiMr0mCGt+vu4Jri9IGQA0E6dUFDaqRbHSsvPaTrOLHwvaMfRsQYcr
VUqpwKGmh5WSZq1Y4/dKl1ibTjCWjPmrpx3iQzaNm46WXXldmm1VpcuWFKeqEFuS+r4CZD624mVv
1tLMLx5o64aRfDGS9Lvmz6AuWkcqCVlo9t/NBEBHVkiPF04ZYz51VEi7ptaEQNRsvleSoTRPWv0J
rBApUfGYrWN6BZaOF/ZbH+txksz+/vyjmHGk8jx1nAo8mg7Cgwh43ydTl4Yy+/nu6KaEjCABYsfX
EYO2jocJZmhYXk7pIuTq9e5S6pxVuqV+bHA3Q28nU2MI3keBdcz0XTPJBvDbiC/wNwe4x2uYgMC2
hc1XbQiWZLhziKmagBoGxH1L2bNX79heoT9iP3BTkT7OwgJRv2NGq1hDORkMrIgney7NRYcdtMvG
KBheqn22z7ab8GoUt1yy8klBH/UfT7GwNPXUOwxf06I8dDczh7Sr0ZL3VI0ZH7qF/07Z92AMYRGY
U0pafb89HG+5N5HJIpoBW3z9kuNGToYBiVo846Hdhspltts+R+FFh6dpKWtgw2uEGWotW/0nim3Z
9mGPVpicqbAnevZSsLNJL+VwWNzD9UugIP1CiNgU5FTQ1ChEWAuoIozjuohWNJTZnUMERu491B6s
xeVRzZYUefoXN5y+9Z8oHsePQPmjfgGt+Z59HGkJ6Lca179pmtkfz0NuGveokxoamXZJRgzNxx+5
iW2djFLlPCPWOTLKSWPDdv9YhrpTMiVbzHeZCLHvs42l7A0jYJ3hg1uwo1KnQvrNyvHci2bERQDL
woL8bzzTUbiRafZkX9FAjUtGFmjHmpnkC/CZHAra4NhiDgR7fxMWxuAbRFYrlj8uZ7yO1nRHkoWh
x6UqOecpUwkHW0F7Fy+xOqkLZDUxvRq+SxWleWQe9IjnDSUzQB9B6mt/ERPbZ4LR1Jl5r55CtgPk
zThSeJH4BQ/Is2bcilONHjxipIXkHIpNOWppsdQYYZGMU+dKsDmbtXNVG4dHPT+x4boVhQL5seqv
IKH7SexxmRVRIht55L5JxMepdoHuD21LlWQtM3mZ/x8w1kSEgtlZewqLAjHPvfJwue4NttELuOte
X/nCABYuDrlD9d/JGAUL9RFU3xSOmByERmcu1EBK82yNsF9L+8s8dG9pr7EIpy0AzsppU4cBC2Ra
DWooGWSSItzbTh+lcKWGETxEBc5hdQMCxV/nR731xKjRJ2x83IW/4kCGjk6dD9bT6PfkV3Bov/9+
DGimOS/ZAIWKmo1OmY1XetZ1nz4AUJBXG4wPEQTwyNsJAu0Qu/gjOj3rWJRTFeDC2NQ//8qyzTIb
Nu7ardW0QJ7vFvP67YU/+B5J1LQHHlFqjxkXmA9dq6Z6tzxq+12errGfr1aHu/uoDjVZ5wRpOMDo
zIoxGxF7NNAWA4IQRWFokNS09JeGgc8AGRUHNhacO6vE8qow1iWUjtLY3luJ2VqySWk57QtMvngl
fnPOln1JRjL48mNwoeAJkDL7Qrta/vBbaPrxdmDqAYSCon4ikZDkiqaL+NSYcLYEp7MkkGb/0bDS
fHpDiAeNAq/omciHt7spEE8pbnvdgy8fBLAEVtyVcPbddfqYAQRt4YziF+7BwCZ69IP71F7mk3ZT
Lik3Xpg7rmp18FeY/uCsoXEKoM0Hd0pHZDsYXn8oGXUCV+rOim2TkoH32d4VB2T8oJ3yeIz3QHiy
3Gy+esKGOakrfFkpWBFpSv8ZZBUDH1SkDvaBry7InThBJWs6mLt5WiL86cus4+cufRxYQR0d4n3A
K8GBbz3niy9eF6/3daP6EgnyRPpV1kvcQHXCS/tIDL7a0i0EoI8rKjo+kc2mIDs8gpS2d/N3jHZU
O67cdNzcm6UBBOnXY/GsQI8mLjaHI9kCPIz2fnn3FZau+zpUXzTPIJaJ/onMrF8h0EwCtkwOf1Zs
AG1RMjtN94x3MujB3TBziVCYC6r6O6/sW9UfU0xiXsY6M1/urgyJ5mcg3CCtqEoeUl+zh8mEemtV
lFDeR35s+HzIaB9AI2mXrs42adAoCCFMVY4JwLnKgjabj5LVjFqf3/Mqc6xat8Jk0FwUDGA/IJ/7
vsSQKOZJG2dpEHWb1aGDCRKjmpajpK6OwGTRSpUF6xDVY8d7+lHj3DZycIPWbsv7JXkGLE/QApUT
eXen7wYG2b61SH59VoICwP+FPGw1MTF7lsyNkOG2VDrnxwVMEZUey0tjKV5LSPt/e7/kkL4NfQo8
3dmfXKUokA6QDqRiMFMdL+X/VDo+bXYWCj1qFf4Pk0bVPxZ5ZvMR7kMjcQ/QSjDxPjQOteZEhZ97
U/x+M+h5JrZbd+AWYFYgzCRkjeLXT2CkbWFI4s+Yu3ty2CqJCO9eMyiaG5WkGxM7TO7BuwJqZwka
fIFcuXoyviP4cKVrysV8TtJYeNnq1bSjzbYav/OB05xMzh8mYOm8niz/T7sN/yjgDY3ACM3zbS8N
DJK3PUY2gnzse1TSFl94poKmCsaWDlhy6SALnq3q17hsrroOTVML+qu4NtA7/WjOT7jYw7lLwIoy
Y59kyNCT0Loh3j33vDW0n/9mH9NChVdJRKUTt11KE0sQWdghqTx/imVky83BDmH3gOIvHNs4wlzh
Be95mYbVD88BqgjxtR7oF0uxQvvsSWBQCgmZl9aZV6uYCVz1EHsQdzUCqxdATsb374Pg1wdF2oXb
OVvEru81Wi7V2czzUsPPBvdaDchjU1RlTJRnzIqKIU7S8i+bm5uvl6On3eiQnVZrg6DT03d0VjDY
v9OF2G0Fq2XiAB5IfOudGFlBpzgLUpW3JVBPZDFuFKNUFTGFg4pI+jZF+hbBnMz6uQM5e/gYKaZ+
t6qz+rtTI9mDCJM4rDd/0ozc50mO5TdzLk95qRLhnun1KyLSrJx/4g+DLfHi67GfEAszJiPLu03Z
LCqXCD71LG2RZV53Dr13GaqjxEmx09YlVJO3jsV6jVF4kE7dBiLy9X+YtaJcfNREoNfSzSlti3o8
N39aLYXYcfhTRhmCp8vdpaR/6VZSiVEqkbch0tddW85U6Zg5LeHCA+qi9iW+qU/u2Z3zsnF1lxG4
q1FKzsDgKFa6WtP2xQ+Zf4voEBF/aytwBYr73cbv1d7Cuy66FuJ2U0qqIY+b65RNfL5KWNZYyOmB
VNcG1aPfTh3U6Dc/KzslxJNx4qP0hbLaz6ByfWtDqj0y9gccXWJI+NUcMTgl40VuZ6HBS/Q1k4Cj
QViuRCo+l8dOfgIjx2B9Nug5ZFQeKqQfp++Z171Gj2L/V2kgTLwHy5aVkO14Kr81IHowqJ5kiBtG
PeCVf3CgtgZ82EzSkRAMZfJECY0zhy4uLOSXun7i4LEViT/obeoYVPkatubAFqT+fH2PsXP8eE0E
jvHvpy+EPNQIr+BUqriKS8NULS25AJcw/2JdN9WQdNehVVTG6kmu0ebus8zs/M/TZmsY4tuk6an9
0INTeSa54RHwyfjWHYh21SSEhJwOHDv1SrJyhx+9GL7I8pnJnhNADsZ6ebNWx2yKJr6kLzrobaYX
hWGVSpu9ccEwNNzT5byYtBjlWJ8Gip/WYnLpT+O+JbdqCizZIKbUDH2EUVAgrRG9kjtXe7lOWrKs
x1Dc5CF41+nIBq4kQdoimYm38mApOMplyDu6nMxM6GY5QIM2VbwYCdYYzUn/rP/O0hzsr4LuABvd
MBxts6cXm4UXnAy6NHAiBj9Cj3/eANjsnzHwxnIivTiWDobGDK6xNzkOiQZpz11IzOcfkkG0o6vY
kgg7kw+MWWtLF8JI1z20gAmSLkRLYCFBnNO1A0vWdDlLGFkZkW1sseqlJIx6QHz0HrHsR/2pI4Oc
L7ZXRjGRtzweHJ+PcWa2TizeZ+FAQinmhLfNuckVizBy03MDv9w01wVCGi1J5e+bJwyAo9T9IIPK
9nqp9WK7y1QMtMPW8R7GwZBtL+pG947mGN68tE+0aqyQ6AFpV203UaajEMHKD8z74cxWrzDq/Iaa
1KwNTGh3jdKbf+3NPExmxljQ817yChNhphsFQ1rrGWQmumoLaPJQl93cl3fTjmtO98yfN8iZbq9U
Ps+PES7sJOVLyOR8/R3IC2D5UPi0TXvhAKsd3k+SKX2TvSJ3kveiG0afLMSBOb5NhcZv8ULmKQ2j
cuhUl7LVJAypyft3zbnORnWkNkA6O4o3xOYOjClcLfil3YYq54Nqcujhw2/4CszFSEhGw9nPqfb7
2a9AqW5mrZXyiGm4LGONtlbY63ocqpq1/ihamW2rmT6wHq1xeUVfZYdWOnvuS/0NY99gbsrWESo+
2gLFtDyHRNjQ/fA7njj4O5J+4okxKWLuQ0rkObHwTd9zHUfyE5Aou9ipMOMYzyO0piGnbkCnSqJF
2GydB5Mo6npVJZp8vXfoa8xStyuSMrmw+aMQQ8+2cbI5bH0tKZnOKy4jTw14ATFbGop7jQZjQRU5
/Mu2MLz25QznKVhIlTzlULt+WYotZqV/qWCocJKJQqT7JHvkYk+Re8jAgeaOfQfGjcw3wD+KVSNU
7BRsK7GcT8LgreF54GqW6orFk+gApZ/bNRb/3H+cmdhQ60hI8wbxBEhWssT6sscQx4N26GgtuNlp
nYPXgAaMVxx34SwAddFXi4Yx2pCm6hZqb18d+pIEmBa47Eu4ZCPPeWLQYh5wxSBcB/UTVFQhiNbT
Qci7HJj7X4zqacptBC+yD4gNuDpY5yMfia1JY3O+LvF4cH/FoKTqzrWu+/8QWFZ+aBZKiIAbqOeY
v3WDRBafHP3vNIJChheTnbwtom5krB7j3KFWslpVKzscgQMAFG/oGfoMnZ9qGk8kqeSOBdJgK8ER
fr/kxYEHGXha+njqpkN92PU3+SC0VoboSyvNqp5W4BCjub0etCz53BMJrBm2SBv7mvlGODSefzMc
omsJOmaUc+vFZ9U0otgU7LqrgtjMmFXEnEMl7nV2KHj1iXGiaTTTJx2sBq59iNUGRVE/HZfd4VO3
PLWkwvl1Tg8/5PiOopBJkBC7v6U6juiVcbnTyaxsnNejmXHWywtDRZPZsr8vabOQXOoPV8V8CW7g
E6PelNZ1weo02m8RKUR1aamubzAv74egFqlgOOWBRPREOChIVrKp8DpUegVpAaMVhNVK4LVPMJQh
Ox3vllCaiOx6IUBBE6RzJ8q2v+fm3+f4aYTUUwMX04yJhvBV3dMavnqwayJ0sRYA1ErG/59IK8Ie
//Ipk6dkYGgz+aL5A88z8Q+JRoLXR4Y/Yt/hPMu1Sb4klyuw/ez9wByGrnt7SQEuRje7B4IY+Y4B
QDQxjv3waRJMaCBCtYtfpY7eoM8zp8CmzgqZrJBPnxt5SRSwSVqhrGIcNI2pKkiMGY+dKDnl69dz
K/TNgPuj6ybFaX0Bn46EFfolFltuTWLteSjfoNnYkdFPg/bqOPNmqimBLSMJmpXs0DAcSHJh9fvz
BnzShshBWXcHsLF5iz2lY43DcLlL5hSQOReflQR8zVvBTWVgrVCm2cZ/eMdCJC8vm22ytAR984Lc
84Ud6HdJjUDNx6RPpJ/sB/SRHuJ37xkP8hTTFK4QW2Vkvf5Jtfn9vfdgr2mdeGRI51HOkdRlyNcQ
u6sKGTqQ/gZYYGQwqs9eZzddfgQdoZ7LHAUCOr4rBbZ2xn0jljPzrYIkhkG4KtUfXzviAk3zK7Y2
3OajNGC44Ll9aqCSXivD9Oo0gv+Q6EKOdEKaYz30xujmmEbgP2WzdRn/CbpugHdjqrwI+vXAvm0k
UAEkgoRLxTEnMpU3TgPFvSJsv02YaPNLCDG7YZSqdZQZWToeEZ5EMyGbu1lyTr5uqomdDV2gT0jq
JPThmGcdHQHKwTQ9BYy26N+qjTUpK6uNftGpMUjdWaW9R1tup0jOnm0KEnLduDsETTxJV6rBHijM
5ts8rEYWHd7B6eUF67Ayo0iWEUI0lgp6IEPCzbdsxFNWeNGgXq6FTP71hVb/jX0F/MKiOxkMH1BH
RuOWqq88CWCAE7gLqxvVQvpaDLVzKuqZuY1t1twryjOUdG6pwt3Fv4DiH8vITOLPCjYe7fDtTpWT
8bgFG5SdCDY3Ia80parBXVryZaegGEgozQYT5InDSENRKtScXNiulhX1Yer7HzSHY2Nrp6uLrJsT
maeqN18ViAKdAiLg95nT5Uj5jmgurcIi4iBniFH3QHVb9X9k0h73Rle1LzYHIaIaDcuxdVMt/nWw
yojrqt2BS28uuW1cx+2aNYZDdb1i4lf4e1dvlUxRCW6/iQnnA93NUp80eQWL5PvFjdXnmhxKmnbc
5ahvL2ODO25ftDQv9eZPuCDstHDmbrOYaruMEjaip0zIFBobEoQNdu/vnhSmvOlPxTs1E4QcwGJL
WpsS5/+svteF+JzCa1N2UpZn7mxuYUtjGANG47rOx/IVd8ti86ErkQDURAONV73OMubbHKXktZBU
a3mkDNIsCOGPwtxtU8sFM3X2BCe5Ae9t7hgD7Q+GcFbZEdIoSX/POd/U1YZeGvnyVqJlk3wVNlHN
UG/0ntJ+9xPN/cscp+IuD0JM5k/GBinPRWZvZJFVhqPVtuBBj+/Jc5YLlGsNs816QxiDVRedm6tr
7udjIIYZ/h+w6/YHuLXm0VCkLW8bP/s2rmoS+OqATcXbd0rLLEXbuWYuPFwrQVq2Lm+SuRn5HFQj
SERYfP+EEzXLUiPiPaLe4LFUzSeGycT1USaAK4pB2W7Np2o3V4j3OWroBk9iXvw5jd9Hg2Hybhus
KJ2CedfqUujB4mgu9jb3yd55/27pupIRIviVQ9Na53SUouiAxkkutkG73DspJUJJMPC1rb4KzeQx
FGk3MIUqeBBiqApiWgWtOOpq1Jns12RWS9nmI//zTjhbtfk4SUO1bkTgMu80zbMrW/Wslx5bBF7+
Whe7WFJ8T8OlJjMHvSC9lUqeltpCAvxgWroPdKyjhO2WpVAFavF8mFAt0L8BeiufMg6D6q4Dutn0
zNGcR5b2szQxyCEdfaZsrSy3kuyM6Qe3dioChQcfWOsZ4bqwiLbcBOLTYLwxqbpk/x1dnisVYOvz
QYwgtc3S4x803RpON+Np83gM4Y+0d4fu1mwg3pc9XmFYoDzqRwShBeRMbtxpAD/63Dh88+Y5+2K/
mAUxE6Np8er651VpcxuDhkE7cNjymiLqcEKZFAuQkPwELW7F2la3sSIn7CCyr6R00CsvSZ2HwndL
KtjqLmyFESzhHJz9o4yz99V78vIVxtbJftGAhjhK+2bNMOWYLsyDohyqXgMG1USu+U+oD+HlmyZ7
619r2KjDYivHprufWGhCJZGRSqmZxzvKDFhx/Vjwj/wbx1J2ukGWNf5a4B6ELgyxyWd9sCT4avjY
tx8ASu16p/mCl9WtHwjXd5ZG8BJ7lKjSwzG1EaL19Bp9/h/mka3BB7TaG2zDIWVp0B78HjN9ovln
ue1zw2x1+bqHN03svYOXiDoooPF/ldN30FlxCJp0+SmE7SBYEajur2+/yLD8ZimcsblZf772STx9
eK9QFgU7Tkoii+gn0+krt6Ix4BJf92FEkpto9ZSosSXxp/F5W0ONdBHNV1hLOF3rhhIfgcNZTdXW
CGxVWVO8fqCc3ieoryZ9vSxHoSMlRjeUiwzdAFAaInkN7rRLv8VAOiFs4CYvG6waFg0p+w2HFWnn
xRxPL4btB4eUP/yexQWbmOGh9bQDVk3av+565s0y3HpJUkpa07xEVFUCG5V0+7zHnfa/aJzHxEa2
hafHhZFfpAen91wc3kl6AFZb1a15CDFXjlV/ncIuc07G3hW7X0dmZQqpveFl70nnwTJgloo+OH7/
J/uCRUUAidkyDKxXpzJJGwCHDolQmEWvv/AcHIqUTfCpUlwGRYQ0bSi0BYu0IOlIPdVvSLG7YVO2
a7/GX46NrEKCwQymBL+7oRsClHHJlwmha6VEwHNY86+kE8nyauwCR/qN7/Aends9z6lMxrc5V/CE
lWpL3YvMfdehQtJS7xjY13z0C2iXt5NRUxnqi5Af+7Tume+sLgKfDv3ErxNFBhergg0U01Altdzo
s6Zdr5XORX+jXcWmJdiNKcXiUQ/kSKYyE6wwP6/M+fzlKSNCiwe03itY73JBykBLQfP8RjYozgKz
jyLrHOvfaGeVd3TvBw2R1oOlhxU5XSDkS4vltAjM+gNF568eUtR5EIZScNleBwCGGPhmasQixfXr
lobmKyW4/PJSjshvHP9GjiZZuzk1IN3aAsIGjJ9+DK3Ub748HQXAaSqhU/G7BFOEXNeeiPyhs61j
OrPOYjsdViQG+kGmLGkVcw0beOs/9H3qIuK0usjxq0PSjLCh+ITdvZ4iHMc6/nE7yScd6khuJsXu
uU1S/EN53zx0bzUVtVhLO53ZpIbSepth7hA2SkFZb6PI4ZHGt6bMBY24/2KIAJaFl54Szo/SYZb5
NjejvryN1tNyp1FhhVK2H09sd0oa2q/2btiiuqnbzN4ww8Y05MPqI8LWvWzqP7swnMnHB8x7d6gL
4n7cuyWypbNVaNJZqByr7cpUEX4B4zsWoljO3lwnB4KO4OxP1cQ+aeZsjB9hXSmjw5PZ6H7mVU6F
6p8bocNZf89sNM0cJsMJ/QjqMuqqLX2a3RTpC43h/xXQrSJxqZ+pL6lNzaQItAvv/bhXwPhJx9sQ
igIDLjMyJlS9tC95D7MrZ7PRjM32DZKCxStt/bZMbS5MQctQ0tp6sA8FuLNP+WNVVFHndE77Zkxo
yWDdpfkpgcvK9+O4kip9D40I38bjNUofl5RxzIFprlqZzxTnt0GVO6tPQVBeWEbxU4w4uFlVZ9hW
EPSSKew2sLurX20DouJ1qG2qG+LkUByudHW9VDRKWiyDZiY172uCkBZJa2hPhk6FC/VosvpTFCyv
Z4c1Kflmv0sQj4GK4GoKm0hY1q8UsGncx3AB1mp/MPJ+ju95nA6dylZu5L0YGoZ+1Nz45sDd9CEh
1J0WDXJVh2XsJQrE7Ia5M+Su3wIvFsNp5Sbi7ftaaRt+OUCFM/aLepqnrFtsTZaxXGycjpldQtNE
JC0Ztc0RduXK2NVE+7IDsfXMb7eR4LXUNOoGu+YbzJd3oIpPDeMGeoXrMlMcSfhhOIxAFpVbSSsz
eoV225BbtFrPzUAv3ewcS0iUOw+q1Lz7zlLj+gY5bkrAMwcxYL+Q3rwh+/owkhLE2nm0iebtO89w
sPJ/qrE4eM5mhFtNMwZphDnw/jbSB9ML9iUK6Mn/z0FHbXQoC004CixhrvN36wVEAV0ZceQemebP
i+MVXl5hUJch3yy85K0RqqJDtKaDbmUbZ/LnfwzG9vol5j5i24N2sxshUuAdmoW15G+tKrmObNN6
od+yZtEkKHC5sQXCrPrNDbdocYSVtrlq+DrSf3i/ozfvxjI8ivRz6Ig0Sp30dJtAS5HY+YAmS3/2
rfCGu5ApDChUtWVp+IJbOVNsOwd562ZUtaFOiVNq/N1mTGqzXMvtMBpAeXAfTgpl9TJMzG59TXVW
Y+MADRoShzQiH/mpS5uMMij/P9X8Dy8IVcm7zje4AIFMpQ1ki9a3WLURo5AvYHl3PTIfYMkQDyOp
QzHqOOQNlKrm709kTyPSOcqXB+Bz9+Rm2vzbKeIjH7UAqvRuGS0C6kXxxsiL1bQpuoGut9Arb0JY
AeknKCGtH7xZ9AAZYhr356ePRSOXg4ueh/DmfTsOv8E89B0wO3yM4qGPsfkGxpw4FcNPwo0b47T6
9H040HpbWgxRT9o/w3f/z1O1s4YoYADfJMCFkjsV6rH7huacGTe2ZL8w6MavHA+1p53SAfXAZfnP
N+zEqjovyAixhm/yKZO1tynnZXj5enrRbqUsNdPOuyHg/rxJHXcVV9WC2VrFIipfVROi95iDWY3v
D7hyO2ziLXAYK2sUZrkb66NcOu/Yd5EKTz5sEomNY/qyuKG53WJ1gqw+AaLKaTxENGBhL9jRw+c/
/pcNNOYUYdTbGzy2PcJH6/jT0XLA+wooVRQxiheE70+Z1oDwvgy1MGG5qzBT4pa/pArDMadU1Q25
LSJ5uqnvQQVuDqvdXOUPnsbYe9XzNK5Pq4+uuoPLOZXP13KVFaEOXsukZ9YtXOCWK0T8Ao1zkwhl
+YDMK9Hm/6cosSOYffILdqx8UmnyZRauE/vhFjaDdUDWi/YXCPB9+rA2bKjJVfE7DlWXldd31mZG
r9TaN5uy9snhkd9G2CLbEMryNv2VLDkyptqPvTIsqLq4A6mn45dvNLFBCXZTYrrPwUUOGON3kXbc
xEbLjWQ55kG7nw+C7ICgo7bqSH4pCqN1OQEuUYB5RSGj+RgD6vcZG59r8N4UW7QnGX5kh8Z43UvU
Sa1WvPyPkhtt8YjvFaqEx6sSmys/XuLhUqEGNddsTn7gYLi/kj6ymcG9M6OQWNCx4EFBFIdJaBOb
5FbwdJ1YAfciwZNnvgEn67tYWu19y1GwrorB5yr4ae2Capk/R76IW/ITVJm5xoUjjs4DL7zmBiwq
d/Y6Qq9qXj8tqrrIlpQUXT/CwSn1SURp4gurj4UG6Rg3Qg4HuaoxYsyJwP+quLVBatthbbHig+bw
h2SMWfgYtb3V/SFOqh23QbvSVfaWzRayQ88MPyl9pCkD9jY5J5+7SP+n+JwrEo594HPqqTvizJWb
toZIuKEw+HidkNyReE5v4Uv+2Awsb0F9tumt/oY7N9XjxePIiNieyGsppPLLgYYFhM2YKM0NWtsV
AseUpkd9q9gajDCytqADvDZyLocs9LWB0F2e7YkP+HthtUBAeYz2ibe2JUNe0arba5u1Js7hCQCv
tKv2jlQXA9P0kjBhH9cnGuzoDP6N36275h0EkIsOntr70oimKO9hXPfGdrpe9oomwoio9CWaWNyv
1v3sNq5C7vIhqR71gpEigXmhQ27m5ETSA1Ebj4FO/I7RP8ml07V+7NBNrdirzjUTcXEDRUQ70jlo
h2yVkxKQuUbyHHLqP/tePPfPb9/deB1A0HoY0Vv6fSTgVl9B9RjJHoSv5OernbFgEtXYNwU1zkiP
1OicA4kOaEkeClNqBmiSpgr0wKByEcwNsqpeMd1+BBBHdPbDW7sX3He5IMQpGbHBVadVNJg/nc2G
Of/G5B2AMD/C7KSBzTcKh6gZhcP0I8oviv+Z3NnfWqVANZGaQYNrNgBcUh5The5WLBMR2E6d2QoA
qq2iAu72GRkSzN3u0fM7CVvUHUgBUpjyMT8CTR5o2bP9ve/8H9Pco1jo+kx/sr3Gz5s0lzp3xPlp
O5zN/na8K0Aak8U+YSKKDOpL1oeZFkZ06j0egAatZc+5+6LZt9v5/WjK9RtLr+3kQfCwMXJxI6Qo
1Q0s7XM+ds6QPdrhwUozh8FhtBeTV8uY81r5S6Izvp/RDI8E83LR9REqx4yZr2LkcgGsVwOrWbUO
4ahZjanogjrgSK0l6MT9IyVLRTScfuHpX/Dm8NAIeZVEdCHh9vNg8gt33CIFHOEoPonL4Rdp+CBy
/lAanmv25UtR5REhGeZCFRJt30fEuv4YbGGQY673ucXfIktUNZNJG9lVyxzUh4gBggiMW4+m3kEi
tUeUE1FfakiAGmy0dX79qXP45WCGOQDg0lyM1ebdeI5WoXRX0fBIKrXiLsCKaDNDz7F1RePuoOvY
1e5BucNQ7uRCrpDNztgKz7LpgiddarBqBiWQ7KxkamizwBRmjpfFy1S1EUquDKFvSsx6gcB/xSjw
2kN4xu0AIOooJ8mPnwKjGywfHbZm2X4Rr7uKPoQAPaTVatPrpGbjxFjlgRTj5kNeXdfXUQwJRcJr
W8C9bMc32zPzXu3qbFU56t8aVXE571cNJilEZZVs1StgOLXHSgIKkBVgDY1SAAzNy5zF6+WcD3gX
HP18Q6uoziVh4ilglrhHooc4RHw0BDo/NRUgzJJkqUI8ZDfi/q+n1ORsdHInwkzmp4llnXX/Y1sM
rfiBNSmIKQKHO/I1l0cNzITSirgecfRRYi96fTR6j8z6xkG2cykK55yWjCu786ufSUwSZGqP+pLS
+dfSqc6URO2mDXGeE7elfL9IkEpDb5lEIZSv3crD6Ze8oQaXhc2gQ4bBv7SO1vgIEtsBxEfA5xMi
7cUaORmK0w9Zr3jXcMG0uL0QYR+CQqYHMwRwzM7CCH4UOMfGcOdzrBHBFrfwsxZXqJSEv9i8/jvm
K91RSS8ROXPBl2nhbpQTlctPgE6RFCrPgE9uRD8wjkiyOVcc+Jx8Qwz3t1+BGBOhTarDOYS8ZAcX
JWuxaIBohhzeM5rnQP8k0GGNVUQhw9XVoWwXo6z/D5aLDLz/VMR4uc5BW4GDtJI1NxMCYx/M9DZH
bA17eSSfys2HSpElRrx/wV0QuG9VKKKQlr6YsfZZYu5CHuwYY3PMRvFlLfjBmrVgtTlJBxp1p2KL
xy+p7oXyMp+X0xKQmz2IEpuhZBZ/UAcasBTD0DwdOwDj9IL34jaNi5uU65FqP6iZIWGZkJjLioqy
KTtUrzDtSO5FMngOCOORt8vNsayHcpxfc7f/D31s+uSXlh1vW5UrlayjPz7KtPUq1hsR8rc+0P29
qwTRFl5vsd4dW9BSbCGKPEB6on7afpWVRrqBVjIsmLHDQPCfOINTMsfWWB4YyknCBns9iGddl0mO
gW6ssd4kjYaAK/RoZRNFBKOxI4nkz8cSj4sZnufGn8MTpjAxcq6GwKYimiCZLKVqFrleKx8zLMm1
DNDtc5mOZNmKbFtj1lrmilvQx0GFN3QWSv3cKJ7OHzqGyVCc/RqbCv8em6cBZbsLsEjDZn3GZ4ML
5LT+wpGRxY5Agny8rbEsW7BbQXWfnCADH9KC805FnliTY5A0hFxgt9noBjJLjqEaLgOkjycDRJJC
UVqq4R84gKnAILymkojEvAxDOGzorc4K+fsDkCePk9X41dSRo850aEm9E6lDGEkEKumaXG6J/jgi
7ZSHFcRlR9Ty4pc74HutO1Va8W8+L981jcQI343kU6HulT0yWRJVoZwvsqnT7hLZ3spaRfaXvZWo
Twf7KBX4LY36pbXQr0Ea16IE85raIl36knenaixqoNAZTmhyLfIIK2o1n/yynNEGXy4o0dZv0rbl
vSjG72mbniv4HcIsrDsnPZxZh+64lvq/MngHTGuRDaibvDucNdAOZe1wxD8fkBwGueatOssmbvzG
9o6bUQP0nLmVJ9A5RYRa4zr3oTDJ8oAiGE2gG5vE7V0BNt7G5djpcygN+RDAtK8pCtCFsTuYucRz
6Wb6yA8sClKpaNcrh3NIItG9x9KndxH3WA50QYtspAonY+Uz4MmA7BnOdIuPCB+rVqalXi/hfJQ3
8ejaEtqOMpWWQPpJbLcdHQnDM4Xe2tiDVheJan3CjyZiwSlXQKLWtxsbLXYMXdMKDcBc+meaIaQv
ldiBxa5GZ5tS+ZBEG3bKYqfUEiYtPxjFZLCstPemAgOfQfOnu4vs4UToPM1XZns8QkhEaj8j0RMl
JxOgG/cycAK6KeOYhd3lu9lOAI3NiLzVSHa0z45Qv7X4FXtMp1fXkCL1eQ3xfS/cNuszIlITKXAq
DzDsbT9NQav7ghT9SU4eqwPdFF6uLAQD8WY2YYg5zpFurMR4SJjK6UeXlpHQGgItcoO8BbbjbMph
WK3mPtvSMWY3yVrUabGnlZkkiu/v2shW0grglYsacWH/2a68X7tZUI2hVh9GTp3rijrgbQ0dG6CA
+DRRJZ5q6RkUCBy3dfACeQ9JiBU2uiGDRar0d1tWGXTKqPNezwNdpf3/IquQXPoQvCdwIYm4nn+0
F5Nu5aB/ktMilliidEigVEIwTC0TaRfJ8mQAUvQxyPxPJ5Nbv25fRIAuZLjVTfHmbnD93jGUszdu
Mj1EhboUroa/CZ8PQHyNg8oPOzDxNx3WrSc/T73LlkkDAEYIl6NOhspp5zL8UkyD7KnCmzvPyPMD
cHHHdieGQmy/jUZ/cVde4ngMpm5poXGr+nJKvPePpuVT1mNT7eGsMcKyoh4YNjs4X63ipHETk3oV
2TEGnEpTtF15iU4KKXaeQiaXx05aW/7XHScru5QEGyuTrF8ZgDBmvqj93wr+xRlAzcUzG5NAFsp9
7vQn4tBamXq2V3fGHbpDAOzuUbHiFSLFga7V88zym8Sifbk/3QRR643544S2YBfl48qWBwp4A/Ny
dn4UcPY148mgjOTJiOirezjn4NklWXLoE0bGmMSimXMIntl1ZvXA0BXfguYjYrRJNcpL0wYdPgXZ
3YWXMTv/jcAvDqECddPMF+tCbRLHE1Pe9ooUN0jE3pY5SqUEJ9wfSmRvMfiSXHeiX/lwEV9wFweA
wNRx6sFz24ZL6qbbWrEn5iZCKse7IqyA+Dy5fdgY/6R6SNn61jHHnzH+TNwkZ5gc612MBlmYDYkB
nP7TKFOE5oZqXGPPGv5eXurDbKG3sm9t7hC053rHu4TpsPMsZQ7JNWTmmn5p3sNINmn+sy86IbpQ
w+sLE+ui11NBFTluGDCZ7r0UQpfTQKo1f3VuQqsRuLVuU5fCvjDBH/jKJUbKfY2xLZTHWJ3niH8f
lHmnrJRVhl6InCSq4oTgR+nW78eX5wU0Ih9g09f06Ju5Dug6XI+CEnnZyQv9SfEXb9KXVumklX8X
akp0H1C83fn33PqVxnUwdUBRd7h9cD/Fe8E/WJ49sPnp3/IsxGkkjWQXpIRPd80OCVWofVDhGqcr
I+C1Tm/+GRec00r3L1oYKZBa89+8CpnrzEz0MHS9IbpshVOVvvQSKr0OL4uOrah396t4UDpHyJ/4
gJ4MduFgahq+aatuPwU5+HqqKSEKjWB/blmKPXDxyNS/Aiak7Jk5Kxv8JHM/C1HOP3Ke1eXjomaX
MYzel/VGsMcFHssx5TSmbGqUxB1hKRcH9lJ3G6NfL37iy85qrI3IFoeNihsAeYNhNGXQYQ06/54f
sGcds0rjDRoSX6amz88/4Sxg9yXBZP67juK13ns+DHUoLXDvT9JxvESSbM3/EedVSGYM9mB4aSID
QajWlaaXV/2ACFCEXafCKzag0JxVhX8rv3SvpfDUCR+LHQR8p14igbPmpmwS/K4lUFWSli7P7duu
CRs+IGLXjudHTF+OaxOyuieXMzD0hm1zIU4yG4n+J/0bGuCDE7RCNTFUwW6ZPamn7Z/vL9T8+lqN
pgUBslISpoEZSBzn/1822zziE73PfxJOod0wHyE22PqmYFHZoQjyK7arskxGnrE9V05ZISQ5hl1g
XNZztd+mpthCNxe5iyocGIqqM/YaSJ433JV4cAXGh5+z+pfyc44YrkZQ1w52puaMCYPYNqXdJq+g
1UijY9ecuGw6RuwvFMRO2HOMHYWPMG2FgOBBmVX2S7nULz33raz1N2WjbivKubEp5H8XfWwIlyHc
NwLWTZ14s42pY5ZyzCzMwpv+t7tcZvJWcfDFM2mXn5sS3Z4HqLf6jaYUYUt4LfKtK+CGDqFLFsNd
Vb5giituUH8D2qsY15dyJ3H/fLVCtplyYLhbDXjNk64VHTcvTres6G8XAokki+7B830+5v7cMkXA
gmAgnB7Lndc/efEoo4gELdrMjui376lVdMASKKKrSvLP5SGjqN5zp4wFCswLDcXJ8IY0QqORCFed
sWnB2TqFlqJGdOHYkwFHYjWZTF2kp57gwvnmJzRVPU4d1wvERdL6pG90lsjyVGNNZ95ljnKPZ+y/
nwdpGhIss3OGsDfF1aizS66ABDlXxn2u/2cWzoXSGSnMjEJtaEl2y819vM7ico02v95y1hWoC273
lq/JBUuRa18F2C9OsQmufJLv0Zu6XDsMfB5lYUXa2KXl5uAVMhnhwAN8k7ShTyMpCE5xkHtNwMTZ
CbGMOWfWoiLr9XqZ5+dfItkGPPlyfuRmfCsDm245OXP4mal0sJS0wedrnP/9OH6J8UgknTa/wuQk
mSGn6dTZmMbRGuSgu66KnuFeK5avQLbtusjGq0QflExY26FC0TSmiBOMwDWfdwO0/HyQPAQLVmYn
zJs/gRrm+FMJzeNVQ7dPFUdIwFeq7jnMmpXsW+nV+AdB2b+S+Uwgvp//taFqd8fdyXS0rgB4AMsI
8L6RLmWPrcL7vSAmBxj2Xnqte4gefHL04ZPJFeBLsxgd27qd1c4cMdLTNd6sOghVW/XxUX83g4k0
mJ9pg/kGEnmP+SuEUDEA9e5na7Qm4wS/TuS/YtnVECaxq8C2DdRHXRs2yASHJ4Ozcquka1lmrqAs
klXwKADj65XHOaRkVbncKNb6NigQcJLkwe+l9yphOM49OESgDriKllH62FOBw4jrGzNgMEGH0c/6
49AQihrWz4pCHMgWoxQbtNCA1uyh+BvkKkw8svllOnM9rkBmNbVdzplsCA9xCR1+TAAQT1bHfTFU
uOZMDnyvFd0pkTmgVWYVrqY/XfMPuRgBaOslQC+ia5vhQpNFGPeU/oCCU2SlAvOjJBVgcHHfuKIv
lLWLDHFbt0VEi7zAJrYI8vEd1lxRQnc101oW+43I5uJBylOt47O8/0xSfORUs1KrdTAY/ye1C3Hs
q8uVhR8s/m7elMLpqMIZ6vAYkzbygxCugzneG1+MsVMvFgTenRLtEHJe7G4YEBS0jf0GorzJp5iW
KESWsbVZeGj93t5hPN0d2HAQyDwWQoAm4h/qZESTAHkd0ZGX2Lx5IJTt95PyVp6AwsbEXK+IpvWs
+OrJrv9MUiVnpBG7HCCvz4Ri4NdLfxtQto1lv+2rJ5FZ9kDYuzunZ3iwqkMtGoJKI/z/fECYaPOo
dRBxyQSYPiyKcv9nrHauEB/GzsKQcsVJKAcml1k83gLCwYbjliraweYklHkeqV5Jzsy9WrDyObI2
Qd8zFKC336fJ/wwC4APYpiWBkJjVJb5ItQDod6KuPErEEDXEr9DieDMInvYywdepGPmsWtbUQmB4
yV2Pxjg5AUFOQWKU7xe0kKFFSpUJLm+wYw8EK4yMtg1bAumyCrQrb3oOF5KFxdClbXTCNFpfvOyL
BTP1s5XckaP4N9dsma8wxgvqDhPed+wZHiz/PklPrfYhMLOjmzyPduiNDq7X6YDv366fgRm1GrOh
BewymjjVFgaIgMGJRWCZp+3jPLqNCjYVqrzRD6tvYho2W6g1JY5nEuon9PlQtJzCeUbqrF4UD++l
FxiB4MTTnZa/9QZpP53+SZiRMmeFq5b6iHU8jCLjhpbXNfvohYo22Z7Q6kOHxtzxfVLjmG5fT1SR
tHGWh96vuPsjUki6uKzQczBAjtOAUCrmlAoDskkJDBi8IGcZrotI4Zi+ZahpQYM9rnDDFkaFvhMN
htsGjVhF1ilowxRr9FFGyKILv4j7SfspLKdfZW6uZi5CiW8bzkYC1nUV5egsuLwRfLB5ntu8k6C4
9CUsiSOAUky72SeZ3WRZ2eEd4A5npsIWxfWqaeqRjrlS8NoB+NoUx5Gd/f8DoFjVt9C9yQw64V1z
3dZaJjt+isUhrOQeoB9ueymcHJ6jXATB3B299v0mimMHbtUSCBxTVL6ap4/3wThT5HOK09FTIg+x
xefi+tuNKma3PYMSZXmjpMLk+pywlRWer6eGQ+R/ytIe6d5sDh3jDEcIkwkgZvG8j/BpKuGI1vSV
R84ttHQ+YOKNazRwRqDS9xVsyg3CjXaNM1cPx40AV0TbOl+kMmFR91O7jumRa9HCuRY7LAePtWNN
mneA6RnlCoEEcYrICLYeQP7sSQR1oC1JJt5lH0eysvndxvTghojHPAVil0VVxoAhrBjLLa91T76e
E9LNT4Gir9W6anbLCENSJoWVIO0JJtFTxKaog87/uvqIiljkb1zSOY2f8Wx/3tTFdUTPlUlqaYYM
4NePTjW2iUkXqptC+OVob9HbULxQW+bq+8Eec97F4rE0VoPXXDq97zXWAxhUOLr9On+MtGbAr73b
38PZ7A8xG3jHhn4a8Oiw6eWKmFx6Wgy+Nj2kD3LyYon9MWSnhtxheL7aFVt4B1OxZb9HtlzcmHtd
oHVGnitCD7j3CHyIgXmmxmD/1UAB4xiJwe6tHdc4TEkcrA8UoDsXPVv9kB+J3FS3+fH97ji77X4i
aWwY0RQbtU79lxF50w2i93kcIrx9dnGZ03hC+cIuKcX8gkCZOcIgCfgnhUzR8ZZAXtKTWxpLGP3D
NIpzTtM0lQ1wuMCpyZPAdDjFUFAzDOJKwPqWNXc+yEBkg8AOlmKUs+NeXARU7fHsiZdLFZjUnJOA
KKkGHO2Rmim/xo9b6+8Jqhsmn5LkK+DdNE5y/LYTNw1HKi+D7sz7D0D3j0ulwENPp+AiPcIreFxU
mqQsv5qKHp5O+oF19AikwWzRE8PEL+bQpjm2hRNGLsV+VUI/XeRv4VDH8oGHVHDFxLBRUEMHW+k3
wnjwHfBZHsCuxdoSvZEoD1CrwEW7sPYixD1b12idwh6lokpyJ6eshy3XQP1YpZaTOk/a4nFcX8lA
PTNlbPij/Yri+TZBuH8gBqQVyJG/equqzj/Fz7eGVbfc5+keL8aNWSp4zlbQFBhFu7MxLUivFoRj
Arodpd6Kd2jpemvnY1xd/zwNl7NfU7QHzp5wCkiQqEy5a6FVhhQ/YVzf2Ou3enJWtOWG0S+szAn/
XMPbZ5T4qv64jTyV2Blz8PSK+samhAAyqqwRG0CBvOBVeC2SaRbh2fT/czDCAXylvzS0FdhOf46c
WZl1hiDnGjCqo16aF5h55DGMmxSguDrO1iJgnDm2L6lPo11/oJ/3d8dNFAPotTVMqWyiZH3mLObl
IjAEHr8rRDmi0w0ngBrZWBPMKihMgqa5IWpBxsY2OODq/Z+esT0Qm/5XJCVj7HCsI7Lt93UsNes7
mZMN1CDnNyz0w3vAYy846gGDcPVUrFUi2zX+98WL+Y9kzK6QRHEf6wYkiHYn8VzCsolTLWxYcc+O
5xj3n982PpKkA7TwsVOrq2KnJ7F6/m+nB2m9o6o622gysoqncGFYqGC9aby5YI2Stg5QGNruo6SE
BrovVaidaJmRzOWr3sq7bpfPkwZatvAedQWOOgW97VWfOd7F3KhBiFvxh6SN0KY5Yub5HMQKpR8N
nGJmviBiMCNohAQZDqY55GL3q/cAoEFrZ47qwBxylbXYnyjK0KpkzoD3KZ9SfbAvOS3RTAt9AuKq
/yDSQadSpQlSv8sDgLWON80BJrC734cMz/lSSM7gw5prfZyrEnSyQfxsJnE4M6FSj5xinC2kZJhJ
qRsoUa6Nk6Db0oYHYPbY2qzgyVE471OUVXJ0Xcgeqe3X5kbqzFGcxeYSVO4SDk7LzfobnuFnEh5T
Oy5QUwHsbKXcMuKU1zmJABdGUJpOmHC9EwaJ/924r6X+1dk3tx7dNuD6o1/q8l86RYJ9fWxkQcOU
LpV96SbDyLxOFCkcJNbG2I2pRLHy+V8QXrfpU/ABYyFnVjggU0TvJ1U4kjUKXUHz6pFr0vrFzBiN
c8CrRNwTjnKmAi/FLNiwMD7ogSL7egmFQdP0VPdBEOcblJzThjn0aDPTKotaJjJMqRpDGwH3MF47
Z2KNDgd+JZIDTYzG+kniczQWiDDCm6yjToWsnfvWDxcmhWWKUOJX9GO5YJFS0/KZJwFp9lcdylmg
TsytFjv5i/JAEzM/R8WiLNqnHm8SIrZ+r8nDboVSy3uptjXzkVq37aDdBalx6UFZXuuqtd6E8mZp
DkBykq07N4jrahMwmVvecNA1oDJJr3Hpr/gVfDNWYMDwmzg6mHKbUvg6ZBo7YvW20EB+ucAY2ECQ
12fg2Dq8u6MFXIoAT32FvCbiGOYvFbFWk+KQQD1khOkO/ouXnsh+9m/W2rNOY3nS+o2/Vpcck9DT
KEVsVkwmAIyNzHAe090u/3OCbaCs7gtrqiZNJ8enRgqj8qgmFfks94EWappVS6p/3f4ClxJcIfNa
Uk/X5mViDYs6lCnaN/N4iDMA3DRqp08yNka7wVn9vFBxVxkg4R+Iewdug4M/htSRkuxMzVcq2Sel
pZinmOns3+SmaPrLXN8I9SPay+HpxtMABLE9seEqxeq8VLfJT9/d3JXsa/LvKN+n0eXTijXZjZbY
/MAPQwBdRZZTSAO5o82k6wfyomimMm6E2zlzeHi2pE32TWUCMPw+2sX0oOMMYxCC3rPr384qS/OQ
N3CqiC5p2AFMaCc5+NVG441/Q7XQROydIEmP8o8BbrR0wXdC4sr6M7RrtgS17RwdmBSYr/a0Uzfd
qmvgP3/rOp5RjsYaXRcgPeKXlESuh1xYQ4hqpUWbV0+1uQXya0Hr6ug42vcP1tl/AmM6pqsu9rBW
PeeXCBBtZatXMwXgB6dAkHRTVc6sz6cMeq9Mygyw4JHjTf2Si9Wo/EqXB6AFmfkXFns6g5SXiAdV
Loc7OdAQxdewmus5gAG72ngVLQfdKhsgWPuQLyJn4+Ajgqd+TP0r2nj9/rxBxbfLT7OYzvSo/8db
5D0XDHFmK7qdXADc0Fqo1d8QatETtiPNiLQtL+2fmtv+KP3FqH8nxubUOAQZqBuIo1OMs8qBHV1R
eR3rxiVRde/FUI8Ik8GGIXZP0wNnfsH+x5eypYpkIYueEPBL0cJHhgqrQotf45uHd52fFWgAdpAm
KyoQa2b+yp+FWxsiTaHlrNVtKQ8njhdNDYVrMQfBf/bmEZNn6qnb9u8h9GsfpOo5G8VbDRjIZCUc
5DTrqIqEXDlEu8VO4nrRC9y4GRJAcE8+fYk8PR6+/E0F+jUx9e+686OcIehFObznpObXtz0h9S10
xkS2yFJTNggFZzxWuvpkSWwXURzZr5FkwEAPK1xRmHUBOBKTOPxBbMpY0m+ZekFWjQhtfL+m0iNA
TtovDbP43HgSaqjdL6nrr9xr3oX9J/6j3KTzebMAS50wL1S8w8gsZ4S4zxgKo4vwndU6FT+Tj0jg
8yLqh+T3D2lo5ibHfoi02MoaKsXDIz2vQRxs2leLumw4hju5Ws+ad15Lb2f2Ktz5h2IVkqsmIm+C
2q5aHn5MulGRDqLxAxgpMeYTN0MHo0MN5PGI5tQQ0NuNzEzmu42EyWb3pD+45sjIlZJaH0j+7Qr1
0xqo44mFpxjb1Br/Q4+5Vxj9ZiILp0lG153gXnvOyBd7jinEcPr7xhgLYUY6tNaCI6x+fFXSutmt
tFIa9uSo3SHm68lTGQpr3aNoGi0D0XsHGzfFY9WDDNJrW0qc1al2T4xxh0GIXVAntEsTrbtHC+2L
u1/Kqa9jESWW684Z04mLbAZ5+Xdwaps2+JwX0TDEdlK9YS9XlseNMI6DK809/uhJaL5fuA8ep3g+
G9EYZr1vfGrouFqmfLS3zU9OREeq+F90sTWyETEztRV0Pf/gdeRWfvLAG0XmEG+d3ZHBx+dUzQlp
QDjmpiXkhQzpX9YN7rqGAcy9VXO5Yw33aSnc6Jsea2C5AnA9+fpSjqgZfW+SVzHnT7vkaRLStkAP
KqONN4HYFu/IDKaO+Idvyg/MPtcQjw7bDQ1H+rW4pUWPn7xd2LYxuvk/aqwz0twOYQYq12gqV6o0
h/4CE+JABJ0MlxHwbzF0ZhlmTEiVwelpsfVEPdc11emDIUUQcybylXV8ISFA/B1iraQS7J3gY5uB
q20dSoaHafkuS5jsMBjkpwEF3SsLt4DABEuis4ZMLQjdh+3QbAb1OmxJbF293NHxj128Mh7JZq0B
kE8fGqdANKO50gci36rW+lLmcTie//YlWI9I7dlM/r2rom0QtmBS6v0DTsHqInRObmcj7RBi57Yw
HWDNPJgquPhDBtq1uhbZXkgLOO6ucQWZkN2hXEvMGiKt4KIR2c6tgb2s46cPgnNgfAIZoc+5JtDW
IfBxPXrkCOKvAJI9d3B5c4/BSjDUHAVh/MSV6Rl1MgmNl8NBzuSg8qPWzA98qJl78hN0jHDzic+0
LH2C5sWZsHRzNaUe52ytCXk+vp3vilVTjrqkwJdWEP01hyu2KVHAJTtYTO329PKrgQGcKhHmVmYm
nZ2OaXi/5krfpr24st+G0vvKLWf4zvsCTkCUOv/w0f+5L06et1IcIJw0+Xm5LX8LnAOXh/cx9Al+
pJMFUjTL+Tgld2yiE+KDID3+3iX8xQju6k6zcHrZ/0m7Ed1rQzbrEphX/OjZVb1l//Ph8wdaCjVW
dLpBGul01xQOeOqrvAriRyoer4UQzz/ZSdxD6k2G3uyvv5Ya+8dwL2G2FbWqY8dkoB+4qgVYwmnK
BquZMaopCwWgA4X4n7Sw1cQfUfTt8cF75N08bsiVoLKMMYCl5kZsNtUL/y2HXJcTlgDigAiWy5PK
wJxMxEh58BI2ZBsNQYjkALx7E8/QhHHwU520RwHs7uVsOOWDIbLi4QlhG1VoXcDq9Qed2LoBWeuo
W1t5r8Gkjl33meuqh6C15K2esyvwT8mGN5mWoyeoi66Q9EcPD0MJsB9VYLvkd17j2fJgrxtnvA2o
K8sPrpbSLDX65VHGJyBQCyDsUa+WCcx0PYOqC2WiqxaJkOOh0m6uqaosRHj12KE63TwlcbTSL4oz
MtDpdjCJhrAxW1uYVY42GRhklf6qkcbbkUiBcAspNYlr/5Ng8a0TizyX71r5Fb4UQ3VlIkWIWND9
RUqhBXkEffCMrB/csH7mEVxi4MXqLK87LNYBIPledkJWNxQUqITnWe3GPMUnDa7BYq72BogFofdh
WVG4ULu4/tYpmzZF0n6VQ0b1GiHCSmSQZuOIq7oFxqGZwtUze1nF9uxkZ+oyJmsmcRjvOsyGuC2C
A3CQukPKx7fkG1x7ddsVH704U6bG1cgGTehWcTIysyVfJLy2DPNERl94kLcIlNqruOVbw5cMZ76O
+LHcD4u+E7d3vp/N6LuV00SkFqMviEjj9EKnKkSO25fInNQDgvUwELAdFFvwZQZNbGj85k9toCtF
YYf5kqCzMGJnHref6W6AZQCLiR8cjZzmbzm0V19GGk3Ea0en4soziTgmnioX5/UmQOV7MyU7iMYc
r8CwtfkCIGwWLa1SvYHRhrI6B7bF51IddjyWODgipSqXk7u1kjNQCSLjzCkGyF11E4jraSZLvgla
MJ8nl6Xq+OQsgO/j02Huuw4wiwfAH8WD0RM/9eC2TyiBsXAp8HhT1CyCBiujfP//XkKDvnOh/wmn
uEgc2cMQupFko76qLrnUw1XqkKYSWTwaj5MdoBAmxuYo74WAfo/rzBSJzqp5NrlsKVw/AyiZd5sY
AfCwISL7TuHiT6CnZr/yh9Y2NfKCHVVHgi1bc7Qq19rXTxogo4isQ318qFy/qON2a+eXTDJktL7d
Tfu9F9ZxdsouJT6FiiNcr6KvUlQ/qYLwjSIzCd94VuyHRzD8togDwIfxcwfklh9urYZCIyz553HQ
Qk3lH9fk+UKb6r20P8Ixu+WB8Umf8aSFKISuwHs7jlNLG8d8z6d25Ee21T/dR7QFvUaldspUlAwR
fGGXVmAENL/RTWGwHSQtdNES3+i/pHlbAeLXFLzFM0mDfTzdjuWzzxW4k1PNeu6MITGXqIwgj4ID
UmDC/3JfrgT8C3yyFIax2H5QTTNNantuipqQAmzdjOCvccMOtxA1GBCZ3/BmpVQvsNglW40QvILO
DUdWDM0Mm1H/ryFJ8qvnH4pBo6xES3OQuVjYa0gDS9M2MMLqjlf/VzlPmNOUs7iGZD+DWZrlIuBy
BNFJyao8GE+6u4Gds8t9DkDI97VdkPQb3WpSkLoaqb39hoonpHZlgBnUgaCDcun+NsjJQcM+75r4
TVmLLm4nsVSixVM8cBWoPBiXY8QduuwP7+MghBoDlxJqNq2B00kV02Ehyp8TlfIA35Z3xcxnv/eT
Z41Fbezi6vJQltLUakQoWaXeqbS+qy4CKO72ne3+P8OwobhdO0XY8DKE6bMk0g+JxUhsCcl83Qot
gA+QFGNRV54agAuKw1QrVbT8bqFc6JLo/DBduBS8Vpq3Ymifva8sBhQJeCa9nU+5CUddxLUInf7h
Wi2I2KhRAKWf5s/Y+XI+RUalgsTr+lfNScpn9b41kim7P7JkMzCMVKTl2pSfKmqYiQwI424X3iXo
wmxDcpfjBKcpGQZy/O5hUErelhuKHFp7hf/DNm/J3/GSH4oBI1c7DhjOHxo9IorX2knX2I9KN4ie
mrpNKRaNxceijDlbY9FINSgKHtYyVy065QllRYzJ+WXw7lT0HeQXrAoIj+H3QxiWpW2WFtkYX2CO
6LFMyTZXhjEETUIginyI1ZsooJ1caKq+IJaH6SzKdLIYfNFGFUvLvh7cDjKlr58/LHiUO+D/awns
VQyBmDLLd0+pKa6/SWSwSmwQSpLXjoaKCCtG/gd9lpiyVTFmmKztxEFIIL0FWNQlOIsjL+RdUHvc
9x+ULlzp1rCSjc/LNCZOESGfEY64Fj8jKXFYcq7FWcIB1C5JFSgz8oqklvQlAwluXS1EcoqKg7mw
yDhhnmhYXwEVCxZpoIpnXWUyiLdmDWCutNOmds73aptOxhcuPLOqSJxkLj34A0MOI+V1nFldmolj
7Cbo3jbex8wYgJG51la7wFbawC1+VqYTk68DqbcuDQ+5l6B4rUQvXWKfaNYAfTcZr3pOBbmRV88H
Nxzp98TOvedBx9J5KmaNoXsfDRNkB8beJT8e79jNfPj3UpB/K15s9jfiCAhzYGY3zs0ua27+cOfE
+DHs4rRpDRqJ8E1IWKzTJTF4icUc9+e10aU7NdliyQ23XbVTvThTE/nbLyVU2HOLmHTdMDe5jDAV
tcxZOFFHh9ZyNppRLJA835fQK16N7qn8cr9cEySf0YhZkZfaquF846ZmEPdnJPK8TgWzRENsMy+s
OTVPAppK18PbEo9ycGzwiLGpGbNyPC4J502cDMsUqNxFBBoz8ICEj5GuWAyIOx+BWH3a6wz+a7mr
huMJsYhRc6vrijP3xv+JWm/3hH0SRJ/7qvLKxmEaA7rvyNGPhT104SDwu/dBk4iEQ6NHYJreFMRd
9i63iRxioUJmHP2yX1mQTlozzAj8SKNVRMhVJ1J5i1HyTR50OxOea3pHKQ470BUnwJ55YT7hAvTG
K9Z6es5ZKR0U9G2sGaQK1SKyGSl9TegjfMIiKOz20YUnAMtVY5u+JwOLu+NFrjNbeF7Z0ueYLf7m
oiQWhIlhionS/apFF8hULL1gzliLcp2x+z+OwQOcvRHesEPgeiTIUxab7kriczqYGnsUm5thUlrF
lqQ4vRVWQCdAT9qX3q0VpAO4IPS06I+F4bMmiR6Nis/mvR+09EsgHdcFUdE4/No9DNOo4HjD2skn
5zWu8WPdXVQrXSHEkEz1nke6X8QlUiLWeXsi60F0FGiU/4SrbQFtvJYQGIRpDI5LwcogWwZnOXtX
SaItqKWgQk6+smOmAjvdSeWbPc5gYyleCI+grsjkGzK3TGax7DlEMv54KDcYb19QxoIdkLm1A+Z4
et01mVJAZFJgCIG15xa8bXJ5Li3P8Hszi5Mt/tz12ghEjjlRVxQ3qobfY2cUXn/smd4ef5omCxiD
pTwoD+7xKh5TEC/KdSo1sGfOMIllmVHzrBH0LUCyzm53Ssowx4N4z4PYInLL91deqr/DgRGII3qo
ZHJkA+wqFHnn50AbEgEYeSN4egjR2Hl8L22BrLj7A9jusZQH9oF28Vx5lRmG+YhBl03n7PUR+WXJ
vMh5m2sHyi2XI1kjCk/56IFxQYQquWaDOdYvHpN/Fb4onmlF2YoLXC6pLi5E1H9vWDNqHWWmGi9f
dsURdXdk+Tz63TGs9GvUxcVMdeW5QJSRRN6KoBA7qKkR+LeaxRGv8hfdPVLIf2RK/mbm0+06W06e
6UfQmzz+toDm6BBdX2yOYMzFPSASB62r2BB7U7cAFkaGv8ke9W4fGabI9fe/H9jnLLdQYbSe9sQJ
isffZRpGbNP4PaIThDsl2CwIaiJAEZZm550m9VNe6iA4fIp1uE0VTzvBHSsY174muwmK9mPjEbec
aN3UdbaC90lSU1SrSvu70GndwDFgy+KGfDLtuwb3ArS49aLyIQMpeVFqi5Uj1zOg+KUUgdIEmj3z
aVnOWYBt7JNIvnxq4VDzOlUH2/A3d8RW1C/cQVDtpEgBN6GRX08+iYYXyRz4r017QdvzNdAsMovo
1oOtzUb9P4soNnwMew2WA3Vddn3mYXZpoedj1gHQyuS3HwgJSKXacsavSf9lYFnnJFlfPGGpTGAV
Ogy3JT4Vcpwpl74ikXHxvTvr+mNCTc6NskFxsIfSTElQsduocC43CWQXhuc4WwJBvl7kd3HOJFvq
qFcWIGRQAzefUl9wI3qxrvThY8YKFSmYZYwwYCk8c3jMd45W+FVxSnT6MrrX/v2NDYwu9oM5+qZL
gJrrsYHwpdTwHv6iXVb0HvhbP66tZx7pf7DobF7FcSeG1NtZ8BCjGdlhgQXMirsxN86/utWpwoZx
JjO0qPwlosQLVyArQS/iIkQI6c/nwKRakDanQdpCMcgnWEfv0UH9vBW9SHCVagQXLciNCeKGLy9o
DBA+DZ08BQp+gA9iGNrE9VR/hUb0F7Z0lSdqwGsxxPBHoS5mQxtNt1+nEPONJ8mbuRp5Kw4m9siW
aJfMZHgI2wT58RYv4jITX8slvOo6ebLjM0WaujhOrbntAv1k7HakxNq/C0PczLIny2s1sCj+XXeO
/muBGZpNBvH/U3qTTbsic4WOfrFpCjfmMOfxGdYHNdoiCHsSnQRBsYPmIy/PJI1UYwN48XIHTFHD
3OmRMT7hyzNxWgzdqHNKJSnLbWv+eFslxfvwRtQgK8VSbffSi+2KFIQPl6DL7u3RuImTmjKD9BVY
dkUJXfVrJskQMzJDySQNjw8Av6P+qmn3YDZSQpCtrVIhL4QOzQefWz8SIiUx5BNjyPD3uiWrWd92
a2nQ5TXOpt2o++vZVllv62XvkG63TgVhju9I7cXy/mF0BlSFPwGI8EUD7Oa9fWhDHdpw/mzHr7x3
C9Hcfi1/OdsaXDpqjj5RbP3JJxagH8PABIBY0I8lVwIBxmipkEOWMHmqLeMdETyCzaiA2Zw3FXKB
93ArIc4yQnYqLbg8JhF8x/9bBeKyzscK+XiCePYqyUWVVY5bJAYVJjoytUGrbN4lIOYkWaE6LMys
nlX75A/BGDOJfHbZq2sxc4rUZ8bak2vUlkjFfHIdfJDApbnYvFYoU8cFRsCybT5OLd1gK84iD/Pp
EQpQFZ9wqiPoF9z1tgH4t1sMlVUSNxMaasZYy8FpgLQDLAH2Zq4Qug1FyhavY87TY408UmF6bVKd
/btf1AkbLt3mE60djSx6hiELdlixrgvegqL/wScf8ILzmsL0XyG+J6vb0Taacd6Mh3Cs/agtC3xD
yKVK6Bq+OggdI4zHDRFFBhT1dZTb45KeQz/xR3Axq7TG5AXWktq2DKOBgL31ogol12mhnhApuYvd
wtu+jgQZKeujNDenZjRroDPQPggIkkN/EDsymBzOM6xlOtf5747KPh3bMq3cOCPiRiLjMYJ3nDtL
dUuVkevXw86tNROLACEkJ70f2wqTn3MtUADUNivdVL/3VwBzftxqZC984G9Lg/ptZGto8nxgU9cv
GUVYog+ppshg9YsOMDzOuoJQLKPRYKhB9t2m0MKz8FEtq255iWIEV4/gTeWS/M9JsiuTe1wm8NP0
blW1+fmSu1yROKVNkOVJ8rFk3bwTPLdbUbUELVMhBc92auwQAS+WSgVsQkPKTI/3LU+ZuhFBeu6o
T4KBG+OsWQjDIVDkhD5td5LWmJIe44EQyWQs+gOvGMoyuudyueWYA9ND17AXZrU1Ihzta/7s9GVC
O9vPP3CmzYsZxrU9qnEjG2uHEA+EIhynZTIfXg262bAahqAZKLaoiz6kAhAUWE2oPbH4uk8T0vec
k+BH5+8cAq4JgH2JpCeOjW5N55SN9P8o1KvhDr356BG3JlornJlz92jv8sLWFvw1dwH6mGC7T02f
0pAQhHKlS7di9DGDKwgxfa4TYlpT7ZjQe2YyaipRinXthzHUADxdsNOgZbuLHMx4d+cJwYcZQfZA
M/OSEGOYlKhgNz4R/r9Mpn91s2+HYQi62ibXU55InfG+MZqBlq0ILZOjqj06TnupiuY8E3TAM9XM
o0jGVawJPaCgRbcg/drNtuNp2xyLRaFyNJgv5A1gLjvuBr/Oq7hOzjb3px0BP6wjuI5/cAmiN7eg
FiUeKI/NGj9QyLNfZhZX2Hd69553kCY/5MQnAchfu7OPGaWn6E8ES2Mr0/R+TFC8FfePx+CNqHCG
hw0Iedlm2xyKOGEg9O008qlE50WJloYaDV2Nsx103nrUzpSGl32WB/mT2nv4KSiJrD8GxHx9wmDK
pZ0eSdmsf9nS4AwHQhPp0hA0ptL103C2Mpwyi/RcPUtgdGImGMKnRmOptlCqiTXFxssoCMBF9sH5
TvJ+gZ61lfkYWvEWvAucUWAYKok6gT4fhmV7FrYaSN9x9OYZwNY2VPJwyhpZrGENN+FsRlqdafAv
iaNQQJWtYEZVtlttKnN7wWLaS79QGhrPNQsl0Dc+ODsu2bhto0JXF5KHlT//YCd+4MV9NBWYGG0y
va3swLM2X+o8CiknV+CVBBGGcn4TKUJ8THdbLorPWjP4VU95C+S1jmygmlilESeG9rirm39nXeoC
Ba6u2qy39/nQ+QGACM9p1gi9KUVDp78cfjuzsQGvTj467X/I58a84hT39GeHPeNT7Sg1T59lbkNj
BSEFouxzSvugJzxfWVE2E/WRQVwcLqVvbpSBg5k4f7Bi1UU5NM625XDe4buFYBeihCAZo4ZEwG9f
usPRdluDYDZqh7g0wqcgLCoOw4O/HDKuLmBF1Tx9bmo2B1e1O3dofuNUO+C5zE85udxRmAb9N6DG
4zIPHI2X3B9m+qvGS0T/RH7K5MPQp2c+9D+9rLqO46XllS0QQk9J7vc27sE9uMl21iM22sG49M3P
O9xFtFtoJPgj8+JguxN6Klt3qq6ubkeV7cwFbnEky1i/RMS4FXItLfft0CUUjHJYLtF4SeNugm5G
1ct0YHb8cc702Cwh5lDrAHHUtHXyN9rBmO4oLQOnnBb78dpFv4tKhgCJdRlFBWtGD5G6/m9yMAOK
FrvnwY++WM7JTRDm+tfpbNiyXBzG+pc4m/gacy4rW/2NKOP02fe/wQLbpim04kDPAFIvLlGey+8b
oNzOaZ+LqZ87TifBIDsPajyxM9pOPG8EjlZOBc+oVQgMbgxHOzhLjCDmOqfkgQPhxAbWBAvOXT/v
YdAzgI3iroufJAWMNxx8PGD3BQjKnocpoodorSczHmu0Nb3/lEsdjCFIRU/8nao/UKxXpCC4X/r1
zqcSlav9scYwglVaPEqF518IdFr6qoefglUHvGj2+EG3CwlqPcYNs1J5JW4ImlZcZZEITwQZBwFx
m9wuKuhIV4Dd+6fqq3HsOzTXpn1kSoLVzWOdpgcGzXBpmcA7LvyWmrWRqBmaiyxfSfBJWFtApEPy
uKiElAkJrYEJGnuF6vseA58m26pKhTuWiasS85VHiitkJVZhYLezEc8TLMmYnNqg4goxYUr3cPB2
4wLIGrwGxwmFVM7Vw4NPo8O7ZILSB1w24cC18lu7no1Ioj67wbgub9Rnbh295jbPyJL3RIj7BqZA
8F0gJnKX22P+c/3WZXC5+FysG/o2r5rn+yFVlGB+6pCM7bU8lILYfJ4LxGdoMJAhre1Ss5fDGSEN
Fv26zVju058X9xWdkivsp3ycVZWLv/YnAtXsibjYgm6PefpcYhYA3UI08e5f1yKJo+SbbaJfwaXv
HjWOLzRKpVlJzDKOL/Zh4M9vsOvQNVtaqVMkbyuTlJR92I60JXWNUEc+UBaOsHunsOc2tVXw6tMI
vWOtmZVNh/IgJrudM1bHCpEhG8ZWFMH7O8CyKtAqnyRIdC88AmKqyBfBInZBsGSNJEMOioeye5H5
oVgKi1d74vbJR1KgcHOUvUX+aaGagfbecS5JFLa/85JvgiYgpXJMkDpPvoa/8QT5jZAerLnjZVuq
UjCN4ex9BpWz8zGQjaLoLc5AlmZEJT+zcPzBH9IFEvCSTydWuY/YUuBp06bD9XIin53vZlLGuHWX
y5CNAN6xpLDRePrYd4au4O2DMVFAHXLHVYC1F8YloK5EoHts0XcDaK7betRJUJnEGDRkcUnXC9V3
pk1dEMIImXwhhgb3ZeMA2Qnczcc9+hJEXhq+bTsfelI8hxuQnnCBqrIRGVaGZcB8SyR04IwqFgRb
BKraZPowkfO1UhOuzPdnMelSrrhzjCBCXKYCC12diUp6jStcbnJF2HtrIGvluB/t3Z4RbSoBNmHW
HOZIQEDh2ZCjKWPTYsozkuJCuqwvU51KrGOSFF5Ozf0gsGkUTFVkoMA20WXZYe4QiL/kRIX77roG
kofvQEtXFStae30thBIcbmlgw17M3KeKK5pVP0ynhYc60u5wuENatzBHfvkJuDuYIZ2HxgIeCX8U
4C1HodS7+v9zM+bkVGhdjIYxXLBPAdRp9KEpAZHhHv6tqtMl0mVfcfQ94puealfAuKfHH8Yq1vZC
+/SCsHmZOX3DXhndON0nUVL7ECGif6h2ejOl3tp3Kcqa5bcvsHQOJzM7XyQUht2XLjFBSxW8CHpC
LaZQbgfFQIinmt5Q7d80s3MwCmpJ6bDXutFNOjQAm2IHwb+7sDpoGgvzi6cv+l/9CWuL6sBVH8SR
Xaizyqil7sDMxbFuG+lnITiaAJ/387HNhroRO5vLGDftVxIo5XXENosQEIss2COQVa9PeV4Erf90
RHJ9zO8FIyPM9ar4b5rMCJiqEqFw8a8EJTJc+0gskusiv3pVRj1JEw7AnjZ+EapB6aw/kk48cB1c
YMRG7wHPV5QykTeX4r5Ikp5WtFkyNb+49Hk1VebzHuKYUJp8xkSLvVEQ7rdNyoNpGgjA/emkibck
JXjD5aHjwmelA5+s9BCyhQasasfeBsKhaFQl9mHa1aK/GOhAV3UgHS51QzmRcdND85Vxq6WeUWVo
0mlOboN66PXNHLMNGyfrDdEgiU33QABFwiemJlHuuMt1+cWM7xsDedvhBN9uYF51EB8aOa3oAZgu
02+YLx6AG+3lQCYIx06PuFz/+cgjPBt6fvaikkH50iWAtX6+h7GohG85wrJbuj30r/en8BxQBlkN
w49/7whQH8/OnsM1+dNE2xhk6JYYTCQ2L3jwVE1HbKK384Aq6OkGhEW758PisZJNL6ogTS7O/rL0
qPeyyRU5JkZRTm3H6dBo83OXRjSVWuIfEOjRSu3LQOcg+UD2CGJtPLwAJUeiXCCaZ0qgB+DwgKI1
vjLUwUgWTIk62Uvha/zv5Hch0su2nIrFHJyBrlpBj9zXRV6hetL1qQxQKLvZ5Eh10cklI9xGoXUz
X3pmTw097ninANZIz8yNhY0v+/mIzOBW+lh26aE6Y7VnPC3lBsCN0xdJi4GUJGBEdHRw1hArwUr1
lHvgsE6FVM8w75Az3S0S14696+jVmK6/2J1PxdT0UKS8J7SFzaUTv4OsBlDaT3TvViBtlSmc7gUK
X/l5CNow84/esucj8/fT3hWLhkXGqstIvxFs9aGWbMYYt6VGaQamDbTjDP6039onfanj3BHyjgl8
X+ewPUWI7heat8BnUlX9s65wq4CUf5u+mwfRN9xgHG31Gp5T3+RcUCEfJhewyUlzSgnW8198L6ok
EHAR5kez9p4Bx6tDv55deV16uREpUPmWiDOOtvSxXeW2oo5fnvfRmL2Q3DsNhq09PJYPmSkJIM0j
dlL5mXgoCt8LBMTMmTgSubBIncFFhuEitbpAuDOwKKN2GNM4ugaWRAcyHbPnQChvleJlRtuuaHOI
JkssuZrLSRk1K7ykczOJtEVTVzrWrw16jtQRL1hiUKY3JEPt9dXxk1w5JB46AcP7edqggmKmVH0C
TKPnsEDjHvkNhu3XpIMSBt+sMt9R+YeReLyrmXSkYG0b9Gv8cycWKxP9lI9yg/3V97pBzWEJ8iG3
IrVVhstfCYbTbZG4yq8c/E/hoRkIz8fqmyVOTXL/2590dU6Ycw6PCDdpj6bjECgdxVmsNAA44EvJ
mWbZIEh7P0LhZgXstcLVhdAA12qu0KnwIOaMn+K8wMEestS9tQbRH4rt1Vt+aQedntNYEAJ/Gl1p
pdzgH4TGCjKyQmSbknl+mDdyLPQr8NcVOmjkB4dgUW7YKNIh6y/oH3DEWw7pidqymjie/ODv7NXq
9bGXLnWBGwlW70oZJnKvhco+q7slIqQOrzjL0e8mqAHvQGj2o4/vu6qM8kENJNylj2tlDinlNPUj
E1tnox+fYQKr9Fl6rN45Xb73JeI9eIPFQLTP1ZfpZYwuUf60D/PTI2lbCLAy/FN5/+jhk8bZqcZ3
aHVnjELgguO9CCuMJaQEL124lUa8k4Se4xFNiYwW4rS9sXGAYCfZqtuBRtnMuZzRFhckbjh+smev
0lp14vlEHMCa7Rzrc6Yl0mOr8ktlzjIXxuxbXJQHlE3YULYbyBnxTGOPEnww5I8cjRU4bPusd9+r
3JesYUaqWKRPD/+6QOT/34O89nxMASrAeJtVvSMOYY8G5oyysVUXlzfnBtT4tiNkXhrAvvVWicmT
On/86sLJEIevq0HsE90DDbUfyCPmsHZXvDY/jm2DD6I4NTnr8xm/a1IAlhWilF7bE3zMIhSe/NfA
LTWvCmT5AH5sukiIfUAfvfINqn45RmUoL0mXr7LUCEBVkte+KKtCBD0AKLSFsNTmo4Blk4ZbqtHC
72ZqSa+lI5iZSAJN3Mhk4ruRbtZ4x2F1DA7bLMc4DmehKAlhGcpNvCbd6wdueNOCS7dp8Cq1Rji9
M3Ps5wubRiaJAzCcVEI+NNWN1YRsvjQ7ZI3iC4Jfl5eTzdWP5a5pZgIdrxmElOBAHX3zbwM/WBZF
VmWm5mV6McTeb6d1Ow6Dtl3IK+ugZrQFLr2iDjSkCXkDphH7mHDCHcaYgSrVI548XUxZFuNaNK3W
kuniJ5Wm89zexU1XeOabYgTqu60tshem7sS6rw5cZ7EXaV6hVm2mArdMAZXtnDW8VoYvoixl7qta
uy5XgYfkEHieQI1culaNJCZaJ+Ai8qFPmA3VRRbq8JHcKYUXp2IKMvYIlO00vMWwaRFc0jbccAab
1nw/4FMKfoAGFMSdazP515iNMSC1Pekt5tQtIN8GPVwWsK3F2y4ko5cqrDHTlxlWyVIn3taDdyWq
fLGM5mQMtWGZKD6cBwRetZ/ypZK5Am/ytvifgg6JdPzh3pJKJVyJejSQAK4wgG/nqCVENo17rBNb
sKlNK37mu5lwh0RXjkLUj+uBFkl1dQH9cZ1pU/1/46u2SnjtCj0Vc0q8Y6cqtp46NWpO3nSa4GM4
ZsUdFdkwzuqiepBIRQqTY4mjt0oR9pvdEKQa9UlotgnOOY81lgQ8xNN3+q1SMu6SZCNQBA7UbyGp
wSLIbzoU4bc8l+MBwG7D60sU1fRzCXcS5VCe2d/WBhM8vA84HHWjF5h4y9Rljb54ljh5fo95EbNq
KFo8eOJDOJoUUYfoiFjFRAhvEkn8CKcfZDeipeJ9ldcq4wspyAdoCuwaA6odOvKfyHyGKrd4mW/U
5mcY72uDYCzLra0l86gtgby40Js/qeb9Nti/Nt6VM+AkJJHosOd1/Z44NpCqMuusmI1Sm3V4wABU
FxwiObUmfuXBTLCrExE77rT5YacqI1k2su126azO4/si7u/CiR2XcOvDUK3hMPPxXQRLJZ4roUKk
eXU+n6OSpMwkDiP4h2ieXjMyk9HYKuZ4hoV2M5038SnD6zkOPVtzqoCEwwXdXl2nASQYT3YbJ6nL
VKkVNwBVH2YPIN1AjoWkZ6ZclzrC48Oz5zdVIMwgMEvFagkWKvmEcVcIW0cRQXl3b2bFM2YIdQlX
pr5Q6DVVjRtnHUOny6F0Yak/s+DgE1Bu/GnTddeUq000ekrTyJYUBU7G4e6W6fSpE+H9r/BKQMh0
KqGR5JnqncwCMLeH2pjM73z6nLEc7+jxHOf4sGYtE7nvvtT3ZTO6FqUMFkIwdimZuiKwRnTy8XxO
08lNzbzHUNPE5NhMrSgmOlJKDnj0XmkL6RaUNSf0QDnwNfAPx52haqCtq6Fsy8Ky8XRaax14FQ0/
zaZ4AABvdSCRIRvjNhYRMykMHZxguIlddGRJ3ooMJydn/FfXrxHhReuE2mcCcNIoBwpvn5eVu5d/
VTFDQU7Z2HE+KAYEkXimYOZlce1gTqH78b7EuymUTD/Xfi0wJr0TS076ZTV/xSOdjHi4SKjt7Elp
AIJOVKWCl9uk88brKHdBm8D7MSzOhJo20NntsBeOPfee4GItSplFtrgSSERl8MK8LMfbzL5hWc8w
+kvq0s3s1QbVwj0c47Y9RRiEKQBmh0edfWev+1KupybPrFiQC+JOSeCiHlBgulG0jrgw6Ibu85QC
rm2v4BQR5ObYV6abzNgKXa60ZybbeBlehhyySz7mu5lJaaFao2dHW4/ntnT2rR0CJ5cbZhuK7xTI
fYRUJYrcMta086Lc1ki2ylqPGlY+kRgXVLT/qfPNNGqWNj+bfmwSflhIEOMrozz10GFSWQJKLLpF
Q2L2jbQPnnLSrdI1eBPVh6mO0XDlF484ZkjdNVkELs2JFhAdBWte08TKDBprApFp4WUvjsar+ZAX
gKvHYVUUVyF8x4qBu7eNPq4ipW01D6Ebeg5u2Lhjl6BIhz1UJkrhvYuskQU0MnGpi1seTO4kOOUl
qz/7EnvvjIJaJTeNsu13bFgWWM4Erw0xUzk3n8FY5rG7Bq7YqefGOCv21c/UbVNJjwDleR5ZyvTm
74beMhgvsGds1sEjlCCaFtskLWBfQdKHtvhCTNW5DBlO+hoW5zvWBOeN5muTgMrBTTqHDhIyupct
N+Nfg6eUUALfCT/wPzWflJbL1KVMZbg7d41JTi7VaJXmBo8TvIITGdnGnI8KSu21pDjJ6iGkaCcF
W02H9pfJBgy9dIxGRZPu9RisYrbaQ1XRm06RpX/YQYZF5leGM0L2xt5wcszrPPDZ1XBv1ajM1Zkv
sVnrGBOELlCtuFQTL/abaazOrwdPE70Wd5Wlnx0h2+x/N8UFMY93geWmOtcHhkVt5px+D46mLAXA
A2tOeLLjKwTj5l8cOrGge/F4JPoDWvD/AvzfuTzpREA+cDz45RdbSrBEnfJU2z6cs/h+XC+BJQVV
xtzMO2igLNQz6qdNlclK8kraRJmzF7y7+9kz+NV9sNqH88x+uC14/wRnuXB3G4xvpAuBRdIDjpbB
Xnr7kfCvq6enXyR0A78rCjrrHnwKsYFZ3VzPlcCGB4klvPJwkV6opKrOum0T1EvinSk3fE0t5164
JENqyty+RE0teivhb++9WmS8ONeWY2KAbbzOSb4V30gWklX2XIsBrs78M2yj70GATeyMv/hFAnQm
oZDVv/KId5M98jtmkliL2dw/YvpwRP6tnQfDvAUA6cDeFy6gWDqO7PrRaXvWsJjcE+Nf8zTryrIO
COBgF/8eMgwENsjFtPZ12o4JUFUXjIcw5J3RFQFuEKmNAiey8EFuDoucaadS56hn477TGpmrHZJu
+XBnQMjL2wCmZhEGkjW4AKszdqIlY0zfC3TKqF5CHQgrd5+4C+2whqHyG5qa7se5tZwNcufGtpcu
NK2W1qLHLYXiyLKS/k9Cvvd6yEGzkvE5QhR4lBx985jJuvh7jrJSgr6V45sx7cSI7G6y7g6/QkMA
9TGQlRyqKNiWsh04sjGUSIhUuS5kKGQpkWRsB5spsmp3ikPo1FahGkcWwuCPad/8z9GZXJ4HXuiW
K+ItMggNRfiXyk6rTqIJ19skZLktHsYTJZNrDa225oeHIqfT+gm1S0b1FZqnMxHEbM6MCmg5EVT/
Oc/0vOxHHJCA04FgxZY6dqsXvDToPzV/tGjeXwubJ6Qr/nbu0Dqz0hM+HwczZHa3qNsZYREccZTB
0kbAVdy+54wL4dhSgDcyqh+om9U0i41/Iq+fWzdZKDYejgS4HQKUiwIwYSht0SiR3NiSIijTp0rC
lYLn+Isx/0Vpd3Hngbd6dfUL6I3Sfj1X3fxslOJWGTr2O8qmyPnnD89IknU0hmsbfg0OMMa+7u5e
hsSGZci80bzTm1B1RHFKfThjxRE1BG/40DChzAqpj5excs3Ar3Ljq/vJ74mj/YMpaVKk9hHzwlY4
OHmNLs/Rx5jtV5b7WIsbXR8Q2VGOUE1yJZoHpsu4rjMQrNczTjFwCuLeYZJMsrsYS1L0zRLqntBZ
58U5m3LFog75AVD3c4lRSpvGcZ1GWcEtvVpYUvEBmNeJPM9m/eDH541Rrfl/2CPWAOFE9Ap6cUWJ
33eLKhGAuiAml+ZZ+ofhvruyzH3k6PYBOZOx1UjKmMgIH4HHLDQ6ViaFRGXcNSEPQ1/ZOgYG6ccw
WMkBJFjhvEegECOWdxhV/1EXEop0v7gNdYzQ4ulG8FxKVH8kdq71WB2XNR+UCzkVmsPVbOOYYIpH
apkUPEcRmFLv+N5U9hUmMU8CexFYxfpNauACmxWb/xWZBNLcMc12Mx6JGGd+SNT3tNN7lvYkbwAe
4tErqEbBnB5J97x6Gmn5OAapCgtCe2ap++Khw7QDKD/tApixWxy5tkcvKd3oQymeC9SYXdV/fCWh
SGloG/5nWBAaK6aYDktyM5i3orc0Ueohx20tbmt8hh+6+JFrSKAv6riPIFbBUPlVXNmHRnMxupsr
oNDcJmiAKYneUMCsIKqW0/3GbITZgEFGEuf5+62l6XdUPFrzJIPznbeKenoLgUWJ7qQxyqiyKa2X
k/VbF1j3LLjWbL/ixs0T2wZJVrkneiBWCzNe8v1Yq/lz5fakM36SFywTisiWU2l6J8ZdqBD3aExk
vbfrS5628Tr4speYKSE7fYrNOIl7Ta9P8fLhLSy6p0QWLydPmYJElCeI7ihN3oJXWtF2lpm2nlQI
Qs98EuWYgV8D2dINbk+B7if/W+Vlo5dv+RqGbQ5Mx6HzioprXhOeUvlZMQ2huZx8GYGLEchua6H7
YeEL/loIJ+Y0Y8qf98Y8qR4/GGzPySoyaG839VGWQeJhefbhn9GN4J9BolfrBYDAm6daMnxPelZx
1oPOqikoL4UlC9hggbcOPB07/4r/xvilfTuj4R/0UOyuMRYvM1UJb07XzX9JIqokD9zxs/Eu1YTL
bxRcx9vjnrOVcp2Nr8APIZt10KT9iwU+RHU2wLISOQ0iGZ0XBjAD0Y86xBzXQIqdIgjwXMFnkJ0C
A+a1zM24aRxo68ozW8nE+bpzj6WP3Zvz/Ot84X6UbUBdM0jl0B0uTOvRXFy7fPnhUUWza2nwpeZN
rBTRXB037fucJKUsewwIbbdH8gOQg7GbrLaAbeAFolMxb1LirHXCbT/C0uXtJEixog7G1YiydJiG
TiAJA48pMd0JvIJYjhXtzxuRSRogX42DD+w8CzM9XgXZ5l3kHVWjOJxQI5TjJqKUW3VSp5OGqm/y
/f4Xj3Zv8Y/8Ap9YKzpw+hnPKGnYpeSBZeqTb1uq6q3uFZeIRo8L7uoD2uJs2DiSAng7C/YTVaTN
5yVISfKKBU46K88YGVW8gDVL9Vcm7KY/wnq3FaFLOLtI+sBNYGk45xnnTsDCYIQIrQXfWYYaVGUj
A+IHp0Z/7xbC/OecOzxNIEmLqZmSDd6MN00zu8KjhvHdhW2zgeVQ1W3fsIAec710B85KCNg5yAJf
q5f7te8MwuociA5VxHzYutMZO0mGT4c/kQX4Bz6FkiqUQH6hZK0RhYcQ+Y0NdDS2UXl5+PximUyZ
kxH3JMsDjNv0FAWZVBYQuROsWWkyKNVzdO4XVuEAtZLEYr+uKoWpIeF9E6Tmcskqq8Wc9yY+Nzco
FeQmNaoIHyYCsLRG/YKjjZeV2K2gX6o87cXVUurjZPMqzZj87dEh0ArAWB+bSSOcVlRgrzRvrBF9
dMVtvmMnnKRfiEbifmyZHG24AbvMzoStk6tGSBhm5jHCznqfRYXIHaxNGcUp0vkTzbE4UwN6iAtg
RZ0SuFtJELsTd7Mjk7ne1NFRY+EyRjzKo2lVIaYWW7RgIaKSOyCs3zLMSXOkxWVIIGSkOaZ17Rnk
HE/t9prLtlX4zAOdNXP8saTJDTBp/VHGvYfzLn8nbuCURXoNORtYJrF8aF85/4FRH7Ndws+XKtjA
C5/CJUHRU5fMyCCiahRMF7N2yJcu+4IEF596fqhCkLqmDGbMnBhrpncXCYcm3n+uPzhtlUegT1d8
WTcz9HAiYHgNGb/4/OuG21I55ftun2nOXDV0mW9L2kw7RhHluqu5dhu6brUen2RfFuNtDZ20oseM
w+ow6XWMfT9nHpLipzaFvx6bBCPlaDXWHBiEdR7OlQwmriawU8C5fXF9uGwDM+0uvPlgWnMA9UBp
XOGCP35hF0C4F5fyu2Vgchh+mw7xvX7XCb+WvsgMRoOcGQ4YW+lWZeZUi/LxoA12jhvdbtowIUst
3p121a1h1ZgU0dft5mLehnemLWbWpPfkm6oP4ZW5zbIiqz5hghR4mp/T5NMIS6iabR04nODy9Dll
8ya2/4JoHVd4gj3TvDSUapSk2AzWZYRm/7QNuv+QhTwidyjRcoID4AzmD8ZKzez4Q1oyuva4bauO
Em01fa908GkUYRZsQSWWCuOHdwuV2x4i/KEsPyP25j3KMixWPUE2yenXY4dWth30qeltaGPVgLIK
1ub/fRa8A9UB42uUUAXXGVOg0q7QfKLh+eI4vAMd5/b/vRHwV9BMo6YzY3920e8VZyCkLV+q5lDK
KZiyPNNNbKK/1IYCv6rWUIgh2e3fD+ktSGsLbavtV9g7i8cC4TivnmqTgtBenu0EzhdI71B+6F9J
P60GAwhLE0sYt+AOSmAH51pdok94KuVMEtYqZeebyY8uT5InmsRFJOU97tmOWFe9EJ2HgFGq5E4j
kItihDTFPV1Yp6tsgG5RwmE8l4/sy+UapuTLkuyY8C0QLRpAEqOysrDkeF4o9QfUF9V3QTe/dcFW
5fnmS6kobEDdtdZqmAuOnOln38i61zmVK7z4V6fOc9WeGx45evwjtgUNn/UlULy7ppKje9W7UW4u
QuaE+L4Cg1tGtn81E/OT4vPd7DVkuMGSxuHNyLumg1jhg/5ekaf/pcPBESTI4S8iq5QNW+5cFOfK
igguYvqMoYZYLN58dKs8Ih+ipfpF0nrpTU7VKmOUziWwUEVoWjfUA1lcbOLl4AQeGfGw3aF7TwRn
F/BjdlHTfSJwLR+wb8rtwE1FdebX91ErcIOAh4gCR6d1Aml0RPAIj8DQVRfRUC8ZyPKR4hcgq27U
Ucc99xUm2CGdms02vcgJ54XQ76Cb/niTOLlapXAw5Vsr1hjDKo7P/xktkwgbtGzscZCHhUJucA4h
h572o0r8ycfypRcRp5YAe7nDMY+OT82Zhs8G8ZNWZr1OHnSQUWw4T1TOsxyI5U3nP1dH/Yjwy+5p
3JaTGWvZZ5QWyx2+cGTErrn2jZoGKnsimXsZVC7ykn7cmLCIGm37Tr24Mc2/H+/rHhTtAThMJUg1
YpVVXXgfnzglBsLdTgxMyUgujaL1TfN3KVe1qND2vEJUcuWWxnGzZgf41wOcT5kcV/WzU7+KyDaJ
wK4zhSMOGf3k+Up+aLeAMb5dFd2c6IsJv5NCVG9AX2QA0snIvtBNBFONNCYk/6KH2MQi4RLSw1fP
R7DNLa2e9F36/OuP4CO9aMdchPDAE/TLJmhCRiOWjqWUTVWQQ9JaHzVdN9nhQDuxS6IKl6XnlvuB
Vt3CfqWWBUA7UCz+qLpEmOHKklKqaq/kU4+qJ+lQlQg9sGCpMXrtJqD1bbh+f6O43X+2Qr3iGW0B
WGy10QCmihfA03ITBmAREWT+rUtWtRtcZd2Htt82QWqAWr5I4+8+YZpkk+lqptYL2uQ7dopvcI4s
1574nOsVxe0lkxK9DJE3GiqwBXdw2N0yYKkMe61rCb4SjbBK3eGxUU2hysvdz+xdPooka8K8RbJm
K0VGhtDvvuM1HIgvIjySzxxA6WXi+nYYlw8ILMYINdhkGq7hwZteu08RE7l+mwzzPFQtWm+xk8mo
gdVC/eSaMdIE4Nw4QMDZxFcPF5lLfASkEMIbh0G9qFc+4sBMXIZozKRCqmlnnuxUJGcoCz6dlKyx
CjZxvrtozOgppXrdFSZD6TPxlbZ1mFnc0m1nnUJzb57z8DHjsfi+zhE3ltEAMjdSyvDpXzedqOZ0
yZIrS7JKud/e0l8p9FtRxbnGSOiqU5QF2thF8h9cMof0UKUMxgJ2Fl5JwUG2JP/y4so7CspZf6dX
F02p5k/AsxKKK1ZZvU1ohm62uyeJ8f1k3KE1abEf/kPUKvHUFCz9H9otrD21tzGrlGMRiFpGiV4t
YqUad4zi4eRAN2BScme4TaxoQ/YytWT0upmQPZ8OKBsKdN8PtL77vXMRC/F6vnqoh2O4kDZKkv4+
4scdDmLkTu9IAyclrV3Z50Ace0Ek7CBBcW5WiOzN86KO1Jg7kn43Q+jiv8fIiBzrpbvFvBLg9tA+
ozc6JUB2tIW8BfPKuvWEDe1vRAUtR6HNT7g1eTkMrCeJywFY/HaYUJwBCg2Lts+nX5AvkrdO8Tqj
UAQGCeYnaVTiL9pWFbXnXGxQABTs6f04OxowJJHC35JY170furFNXI7TSAKcu6p/g/h7RCZldNm8
AH6jYzNxHu8Qofj2ix5QubIJkW+NHIXbcEHuQxmzVXsP7ws2NxpRTf4NUgNCXoIobxLWXalr7HDV
pO8oSXU8VuWiqB9ekHGus2joqAMFKWhh4NmWDalublbQE1zT2EGYcYxIv3XRgvu3dMyRo5tGm0CH
CfwhcVZxtg6wZc+1ClxQQBT+/xyEKDBZS7QbkHQBJhEetybhOEA81K41o9Bi7nEk94iBj6CTCCyu
qBVyn+MBV9OM+RrXxzpuRkcyvnlrVe11d2S10QC8gZpUA2u96p5w5sF+XglSNv67yXNCKSNBNunf
OrG/NL/a8qLOIMB6yOO8Xsh32eeVvuGuuUYvvcVzz+n7oE2FCWCLceggu2qmfh+iUOesvXsFWkgc
aV7Q3v+4WcEt5o9rZI9dPXcImjjz+UNzC5It/oC9kczyFye/DVCXfBJ2g210dViLxMGHiXweGuCc
IxCDbLXD0JbPmE3ndmwkhsfSdBzpkrFh+vbD93GmynLj331x/RkPDp2q/9+GTtVr1oSxCar+06tF
t7/aEHwbMR1j3puUVgjAA+W0jFIY0dBTBs6cf2jA3nG8bvSjLN6ch/3tKEfz3iaJxCjpI943wnj+
P7W6F7qf1zVt2i1IUf59qzPlrKSyinRDSMh+f1IcrrDkDZGJoSleWY2hAwdIp12UIw4YNrXTYywi
4ipZCgO3AfydsAdoPZYdWz4vLYiSKd5QViHowqnfo1RYRVi2PJPAdm6qs+rYGVm7oloIz/L0GmDy
WPE4ra1yOGXqqaENcXquEhWd3q+65XJHWN3aYzdiamZuv0XgqTA4O6AwD6mLUwmXlIj4VIS0Unzz
Sbf9uoguVdY4DKrXNUe8nNamrrd6UO7JjAdpZKIp8oaMjzxtddaAADvpKbzQ/yjYr4NuxY8qPQjm
eRlgrwAGA1V3entnsx9kJkTGLzuDs7JbqtHG3BHG+fkoLr8NTCatHChNpanYPYDDQBzcHN5v8wDs
/Xbkp37uXsW2XC4I8E0rI8v5vYPvB+pH13t3kkX6G6+QCGx9F2N2yYLn96rqXyKxD5zrRJVX1H71
N0k6M3vwNycHzDhWAHuh6AQ+6HV0Ypal+5+wmVjK/iT/03P9D/bSBCHRNXTmPsAYi+nxd+rJR5ws
A9cpxtItc0qawihhUDmbeaWMTkNLYeFJpnWY554odlRzB0ZI+MyVD21na19UnlHQUys9l1mNKBcP
SoQem+ydhu43gN20Mk3nOdkt70129H/c6DS/8sv4uPiTXgK8RqyGj/MvTXG4LSGN7nXDuD7Dnm49
KCqBheDIzQFZ9Wzpksb89fx7e60cf0cCFrUQlgGzF8CItVWS3KcL6Lbve78zHzP599SLnxNNGKKh
joVTFKOGK+i9uNxwh1qTbsBki0UFWb85mhLM+SVJ6Kxc4JD3rMX99iYbzGkvjyYeVapQXpcAy3NV
U/yGtkPtkyukzgxBkCmPmkDz7WYw6yvTj8Zh0Qx7wastHy2NUwmXSh2j9U6TandH4Mz0fY1oTjrG
V4wZt4JkwzMQrwjIvqGpWkVBkqKQ3pt+VefNaCqFg2uQ95FsgdbS76LudvyuVk73OZ5daAbpN+o0
yCVR9xDbsy34X0c4HCJlg9KanFxBeXJ/+LUPiTlICAMpHFXO7yTo596IK8aCqSzY13fhWq2nXDSK
xj5HfNE94EaBvepnJJSAism2meOypC+OtQRoNhXYyzWHcoE8okBwjKPetJJXgoTbmyCOdg6S395F
UDkkUZVXUWx/rAwtOJ1o++MnwHDlAkEbt24BtMAoiblWxM7ktpzABLXDVtlBeQJt/fe/DoGfVg/P
N53SMBkW2yc1Sk+mUMM4ayhDpCr6ELaQAqGkMmFTGVIcwKSAx7EYBXngp7zP59V0+p6TTD8SJQMw
TaVPZ48A2iIWNOib43eUqy9Tarn4Eh22fk+iVVp0rvpeJ6gTIoA/O1de1ZmXHlKmsMCDbVfR/Vc/
OJugMXbtfEFzSncuY3WNuKq8S08FKAZPjM23NnnYQqUqHorSCnrTiLbDlMBxg8P1396ilbJC9p2C
/WYUTIEW6q0lXAUFx1aZCK/wO2gbVRCIiVWGFLAIF8IAjQQOzQYM0nytqLBPnrH34ZNI+ztLmuk1
k64kiDDSG9I53ZPbEH1dHER5t++83GeDGdrbGqa3YclhbyUphsq/Y5XAnfGVLxtigSx/uqEBFYlL
c06vk1BBa9bM1LtXHaLBPDhwjKjN5wBRgO1cuZ+YFT1RkmEoTp5+8XETaIbDVDjMlG+c5hltknp1
zfSMN7Fkh1b9QTzoEcaTBX+ACjkL2H8ZpIQbNq8q1A/DXGVgHvakVWqf73ZmWf5Srl24YSAN6tHz
aodbQTNlZdwEk0whCp9pdMTXXb3kGZM3e7AjjXfzG1KdUuqxdWmv6Nikx66hixuPuGfLCQ85LcVH
SijxUd+5XylxBza+tEKeo7DpoYXLf8TQv6k42XeAVSQHeWMK6DQj4r+j4aE7OVBmFeRCEkkPtwcY
q1bKG6UCvejse6QRtk0yxfMG2kTmTic+YszkZGpwHMvsj1V1g1a0W9Ak3H3UQ5BopatICeD5mYcj
l69wa7qE46oetY+IQqbpmHBuhXYsUxhQTGOotpbqFpCRrB6DXeW15cz3ZYGmk23bXelHwJ4PeQaI
uihKXtk53y+NrEmBxvIbmrCRMwIuhdVXBHznDbrP7kYWZUZQ1kiJuYgEU3ANqGWfEu9BmJ0sAGDp
9GT9MnsxewWenAgIA43xHu3Xh5D0yckIaFQr/0yHSqCtiWJ6M9JrLeiTmzjwUL83Y+JOHKnz038o
Z30KpYLaIeQMeLeMnLklM141TEXakmTgHk1B57dTeSykYV53+8KZH2xk49WlWqgHUB+cBS86t94F
H8t3/YAlCLg3UckzBD9ILsTx18nPDdrG0slhu/XbrwM7/85IEHmo01KQnB0Q7QmeAXViNX4AjQxF
myjx3Mh1u4s+BvieasSYkXvc3KnmSQNPzvECt2KYr9c9wFNA1EO7/I43d2P/MCoXUudnLNitefuS
pyiHN64StGY9AA8d2W4KX54mg/lZ5BVoVB2WlsCH3IZdAUavylUyDSn25o1tHA7G5M4Q1v/txX6R
tQNIpIb39EOemq+Sgjc8FI/VaWoWkT07hnp68WNPuu67Qj4dFcpuk8Y6josb76o0l38gl6ez6qLU
6L/o41WCzvhLo2qHD9QO/NqKqsYuVK8/BOhYVO7zk0Y1Y36EbngWf5RY4Iir0tTWdOJioR1pwpXn
BV0Zqqt+XbxaXRA1p4QyFUahkww1tkoLIpw95RAScla+5+uLJqQbPDM3tU1/hvu+sPnCEIZJ+wnu
Tu8UKd8yJiV9u6X/lVC4frsA39wGLqrydBAd5thZ6avXST3dBdBfxwN1B67InCRrVwCJGTkevq1D
dDrCbjjAfsjpLVzz4Q7UDsyX98EyxnoSRAOWkRiCKf2dB647pUP3O4dOQwEBQ9ziGZFGE4i2P80P
kQVY7ZE+tosFbSyyr90InT7BrbbCa0o0+/5bMzBYYQ7IjZpWB4PkMpBNOfoomDau+RucBfQ36YqL
hwX3IuQM2lYNwxQ7SUiEqeNEALBfgqaqudbh9D7HDnTZWmE+4enFUuRV2eRRn72BBe0cegVEtJaC
r1hFMYf63Ky15zrSboEMIo/a6ufhN9LsQS07xRKotLONv7XrdGWUN3EBpth3yZRBb4z5v3a0I+jq
v3V3NxF9cUho1MeS/dnT948VtY20K18hehRQjuMw287EgrnLpxVWgou6VtYFpVu+L5Zb2gdHXQ8q
/lQ2Tbyg73IjX0xJG0g6gJ6IGOrvZGYvlDEi9AN1shiLXuvP4rTEQ8r2crKOyPF6iLNn3mjmMb7H
jj/3gCRYfMbB7DAAhkBGjp216IZOGdV1OT7rA6XKYLZJ/7qvyBPRy6iMUfX5IeIsA+RijLDwgaSZ
nuUKoT/mjEQCBMObu7qIDh0cGdAUrsq7Wa9BB1Vana4YgjicdqfJQn8HAv/ieQG9hgw0ckTwLgp/
0FBTrFVFJ2ZRKmFLk/Y/kdptqxALS8fayKfDntPXs1/wACXl6vABOCmT3CRRxOq/fPNNvIZEgXsH
bUT78eD552tE0nBGeUeV4zA5KYa8lQy2Z7YiorhLtaXms/vvnLzmKl3r4bNyoN3NsfwsFLlxiNNO
KtLvwKbRIZsP/ihoHiLLKP6hMR8MH1Gg+cbUyuQkabFYbiZD5ha4hW/itI4A2KNYsymRLTaAZgK2
amRkhWsCJI31ux07RoaRt8lPdVM7jNDIA4D5ezLaN0Y0X1G/BxybS7bbTBypLRxQ6fIwRu8ixWaw
qcJ/PNKaVbawi4ry6XN3niI/N2s4KvMjGY82TLHU7U656mGS1sgTEBKH3IkBP19kcpV0AUsq6vJf
AKFfOR0P0pI9HGynj0JSMjz82Q0st2no9PnriswDIk/yVvox30VQqohYxjtmMd6w5ff3q5eEnpgY
2EJSvGYYw09AMANHUgv3MdcIhfjhNoQ8RlddEhwqRcgpkF2EOyScQGDmtL3Dq79e63ls0koaFY/v
/LxcZQGI8o/IrPjRCC+C4vokuYWSw0VpJ4Cwl7NqzDAHCqnmpO1Ug8nhqV+XQ9XPop7r3jvAwEnw
R6Y9S++kjJCUInIP0rR6DA/0EYfvEcmufG6TwwzZkIad3LDCOJee0YczKIxjbmLewYuICn4uBy0C
2PTBf5AGDX3mORX2cy5CMb+MleOMfyx/pXmACfMSOZBh4FD3wxtYxkLhZGdvCu6WLCLfS+yauLa8
wqSeUW1OpvQutoNyxgmMnv9lgg233pc69D+nayJd99CGoWKZ8BpDRRO4F5O0nmdj5k6FZn70hXqj
J9884SemBAUigmcjtNICGT0iv1+owOSUlXa/f50Y8lELpNDtb/JfPerwFWIs471CI7mAJz5L74XG
onmmJWfE814WKwyxAjF9qWCZDSDjtuA+oU1i4CxOMZPZ5KRu7+ASISAds82lboGlzyZO05Ditg2x
baYUlUCOIxnaGcTNyJxYN4VVV0jKMJMage8SwelmEI29oBcSnuwUBEuxiK+EeAKwxYINyOgbYXE4
1vFGlaAcaJSdYWDD7ysWWjtDNJyMm8YstTd77uDl49RENX5TO0neoDWUVMRMv4R03qHXHZxpFRaN
4CnhcmP0lKW8Tq1hDT8M+ZHxRemYyB3Ke6vkeS9FLxXtYgI/RSXOYdHV93FOAjm846pLuZhVvWme
aWQJGkY/l2eHE3cSlGQNlRjf82Qid3uj8YSnpYcbJGVTrPbxbcvrqoFsd02NCRhMib8yRH4OgCIv
m0L/nVTeSeYhATGtTTeZeNTgLBJ41Prheip4fvF5DlICJhWqRfhCOeV6dLlWa2R8A9bx3boU/NoP
ZlmgCrDNbws9SAxCAAJquE0/etoD7ByRmTe+LlMMXsxjMSxaRYkDsE8wzgGuV6Z+H66yY8XwH3pX
6ksyEkaTT5meAVcrktI60L8N3yxxjc7AndoEEKz1OOztBPDJthhpDs9XiEY3ObA16sgi0wygm5jn
JsSFXL0AFln7/cVua3Tc8beFDagc6S1AqkeD40dalxNECaHysr7xPl4lHC8Z1Bk50EnKz+e2XR6P
bY6xdsqScxvB7cmrt0oUOR6l1f5FNbzQFeiVM+Rbx4dLGi3pqzZA+tClECJkPMU4UAL1NFgSZtuj
pKdreTP6kTAqLuMvPuaXaNID1+3a5omFn28pkqp1qmvQCXNBkkZq4D85YqwLLx9wAOSvjtE8YK+S
lVgqm8toaQBl0nbYWFM/rEdUWRZqW2jkAxqTYpoyfzm7knTEbz0Jh+418gNAwD2/gOtD/i9Qagzx
xilrXFEts3PxBD53bF4dfidFFHTFGy38wafkj7q9CXRRSt5CLr/wD07uRoOFnenIbN6yKUc+chne
dNk9BpTx0CaxdfBnAWM5/kBEw72C1AyRKACa8CGTcwe5sEGbKNiL/nNL5p9l6JZoDd+VCJPtcIi7
jRmBH++wcCOo8Feocw+OH/+/wYEd7zGMs/f0hPwKMo0WLiOwOuUs+56kQSuR29ErGkhYjQCKzF3X
CrVm1P9FiINqotftoa5+5JksNgTM7DFWaJWv8Fku4ot5KyHLx6Kprt7B4LlwgT+TP3OId9lR0aKU
iQn7c0Koz2T+/Bc/Sk4t+jPLRVtYyNMUUQlMEkxzP4kf8XFc9dFsd/kEgbzAiBqlvoIWLKXI2En4
5syRklmxZ6CKR7AGN12N0RrDLfkikNxL1cFgOHGWMwxu75nepMC7mDZflD1KP4pRuN5u+B/GDVCU
yFQeToyt3VFQ9B66En7Cwg+uP8/WmB4O+cGPjPaaD7v3wQvIaNP2gs5Icn6xgwQLrl7zX7HUHznI
PGTw57DiUQv8qpm6v1IHM1DK+M0Jgm+pGBvVHxOFuJH69X9PHfzevNISfkZ0htxE+YsixAJJW3Tf
tFZyZi0lPptKFAGabrF2GmAcGwwC1DNvRcP1BUIvQPpbpUMHHwtZMb+19jbE8FnhrBwZahJLK0Lr
Em8wR3cpTpDx1/9N9A6fRxtJixN5a6uPTu/Tiots9WykYdMC2g+ElLHZMVV61q3OjwZKfuwV1uDH
tjRxbbzsexp9/FTrzhzeE+K6AbtCc44Eysem0Ak8tp4pdnhA2jrpJVsJ6yLZTi/uFCTOh+mNR8xD
eEe0x0cWTm10Tg0SqKz4ulZCImadpKHrq2wjcCDxFUzExZ/5wZXk7ZTydDr2L9Awo6sC7V+jW0qU
T64F50JgWoFCyYSzB7yFsEG6Ic1UBAGRk2FAU6DwhZmhkUjuFcbAP6hwkTsH+78xEwqECAgeSk+0
9wWB/tTwT8hV+ZQPeMFABE80VukGyVV7A37WvZlv2fWSr9F8CkwLuUDkSEvja9lU3W21JiBi46PH
6UvSTCi8kz1p9kGwcneBxQ5PK7vdXQIv6SrZ3NBOtn+i5OynyLqz4wREiDoZSZLnSjDEGY8ESdJa
tWRsK1rTpNfj+LDM2byEy7aiwkiAqWUtXSt8NtOmuccpdC/522PuFg/iqwe7gaQO4EoGoXIVrtr3
VItRMzrvRq28DobTJl/YI0qewUvdLfs6jiL0RIuf4FUc8JAElXdzoUQvEyvwH9z1YvcyxH/6Rt8J
vQvAkyZImh6540mimkmHXpcfBqeLAELHdF/DURyoUmASg5QKNi8uSjtkihIrIVDAtnIsUuaYzBum
tCdRrSz4faoC/a9jPw6S98WVMpB15aNfG0d4qHOpvlso+DfPFg0GqrBS7bjwm1Tk/LW7scnhfj7L
xZoMI90dYyxnjYzRX1miEtmvp6ZFd16oBhZXnqALMYq1Mppp8gXIg9uo7mM2VdUe1/Cb+V9wrVhj
UJ72o2UAhufNk2Ofdk5yxxyBlN+KsU9B0D+AhjjThnSdtIWcUPTEox97aLHtS0Xu4j6/FAYWZAZv
SUAanVf83seqah8dcq3pNqTIBCO0C+PTDJUqyDqetyU+wUabaJIxfa4bzIkR6EGUDZbY4nxOXkIR
IWz+/rppsRhvDKZIYHrezYXWkbrBAdtl/JtBfUq5Lu2xFMdwxwNK6EFr9mjMp1/9jSqRcKwwU+7q
Ov2XFa7qnCNPfQ5rJmEsB61vHniIAt6h50oH1dq6JCgORA/CEDORNkNw5OdCbNtrL7tPf9dtkzrQ
ugxgnCG0qrV+30Tz/nDR6N92SwzZ3IQuY1TzSDd0RX+qlCH00j48TPQIuIZ1hwisaONonxevV09E
LFcmoRx4oUW2hL4rgy4IzUopZWsQsM+zCEAx/5MyZva3DwZ+B6KNkSC+cdLEErOBEbrRmi8YgJyr
JkEX86fIq3xgxz4SKUpN4A9niN+J0apL7OwO9kGj6vEpGn1NqGblxjpEVT/vklv65uIh9/8PC0Rk
Z/QC5XJzBKE84uTbpJf+GRpsbRjq+KCjs1SVpkZGywlCW9oDLBmRNyOT/kMuLnzjeIeRQpzL6486
knVBXNpNEQ5jDobhN+kO5OyuntyMyhil5Kzv+KQIcNduhMrW0aaMAoP4iQ0fwzto1ggqS9H9nmMq
AI3hybS5BMuOzCk7e7/NhcK6lPzB22cBGCRIaO9WcXBgKe6tnSg1aW26tbbiq4pKGHMgEmC7klbl
R25p8t8JfCytE/PIOnsZmh6YEBYB/r70n8s0ZTrbN39YOQBMDOdfxvVRiEOxQO3I0I23d/z7QLPl
j275mmu+gDYO258cvME6vZJlB0KTccT3nsi/CXlHTRHsyZTDeZjqxPsY5v8EzHIpPPjbZZwIQJlg
zhUGr9KZnux3PWK67rbztv/x/cYVXJkces7YzpJvUzmA56EsYPjzndhxqlC58k3LYV58RhpKM+gA
kQDb1AKY57bcVXqANfH0aDZKcExZ+Sk29P6b/NtmT7jPMrFkk4fabg8qWs02+jyNM467TshbUsWo
1n4Z44STI/Os3EpMVRvkz+Rkm8Bx3JbLhELn05sHPpU6mGbEAD4OgnIRLM/CA+1pQOdzjOD8KQJP
f7Td6Jnzv/g24mIGRGARn4WSlb/Ewyns8dNrYqf7QSuZd+SMJLvRgJgDMG/27MNOVfeAFuVXBR6P
Hm5HyUwCf3dfOkM4DdnfIewPYmAhb7O93f3Eu6XMXQ6J9Q7P3XrbOcjD5j2RDD1QoVhej9PRPWuK
EGlBvZBl8e7ySKXLfbKkcDjaTPFN/1vMrV1QybBStzmCR1fvHQNBIaSiqBrsl1PCwYXjjTKEPasx
ea4DpGLPD8dkUW8GLbhHamZIiqMDYWeOWXCZN1gIR2wAciAhCF7CkQe/3/U9bm+Yp0vTpf5hwTG3
bS9aSF/rIU+AikUXI/g84TAk69HoIDWm0nArEOL55R1/r417a3VhldDuzi1ztL/VFsGAtG8dZ3gO
fE/dathkPw1nPcYGI441Gbh6J8GM5dQ1L7SywXPy+kul/O8G1rWvh2k3opbKCAG8NrrPyUZKYcNU
oltJb9WVW/fSOV0eFXnLRKutxJD0KuebZi/8g+S78THRZpyeAKmkBUbG7KOrBqNGFJeub0DJK22g
Mj7Osik198VVmXLczfevdm3xHgH0FjoWQW1F1ZJiy/nwxGJXrandA8T78tyQRHat3kaQIEuy7c5R
9notdlQ2W78pzA0zRZSFbybhUBFQIuU56WrR1OxOA8gn5U9c917i6Xn0qOHJe5vM1Zfp9A4gqyaH
0yJAlqQSrjzzWgRra8z7PAJE8YjxpY1abhzGd/SsY5y0rGZNXkN6DPS1vi82tq00YjJH/EHTobJh
BQwFoPBiUBMBUXjkU08D6/6Nw5jNHDRbJXttH1nIWYTycqI0hA4Ylqcl1RUuuaPqBl4OBnivRGU/
Qbf1I0kbzjIMRGffHYiGAZ1qYGyDk+QNFeGDlgkXcw3uHEA1C2KoKqiCaJCF3bxUcHEHC6HmoYHK
j93zowOJANqC0yrHA/6EEe4BlsK40uuMFdoXnJ5ldpLXXjSnmQf3lpQTwzhBNCLdDJd2dHeQQaAc
chTn6kAJNzpsG/47/N0JUIwyxITHME7gyjrpuseXE2WtmDmsKEX50RQCqt1JHARmrlfgFgcuAY4q
GUOI7BJ4LNtPxE/9K5Ehh4eqgOfrfH66SfMYdXbFu8ItPQVc1AymxdS7NHPMdDqazaV2yMr8GwFs
hVXjbUeTdJFdZ/3Pu6e84Xaz67cMyewdqpDxuufyvx662Sr4RrFPLdnhOo9w05XfDM4N5AV0Xskp
9s3LgqeV18HyqW0q226T6XykxbUeS/SwCni8MeFHtgG/b2dDqiwy2AqTmEAcR853H3ohPB3eakhv
5VzGzTk/T1ndEq2w2U7X/a7QoVD0vyBhOpw6KTxYPBYb4aoQjWX/4eqNpWYwqsnrqyn+nBvfAuoh
cTG6tjwHy51YYGtYEfp45WfgLZftkIKlCRy7r5TvJvyMsNrHsWB9lgPnIX1TBk6GR+Yxw3Be3wSL
IxyLlRc9JB0FagURIoJVkEkkuWuiQqhg8qFfonSydmnXZDjiRERgTggu691r2NRzbtxinXqZ9z3x
ly6rRMXXKII+lMgQ6nVQK1DBqYlI4ojL7Qvb/CHnOb4Q2dAbTTrOl2ILYKvBpvV6MkIAZAslEHvA
MCjuzHrOx+jAaNMrlKz3h6Q8mFFIObvrg3CcmcfEuEssB11VWdJU6rvwyVQ98cdY/8eHs1nyQgo4
MYvJZGr8Ui8AnYdwSe6IPJjF/saDsaCNp9Lxqc+wrkIA+UjvBI6dDBZxJavVeWixxuAY3i+Sw0FA
aw5bWL1hhBExbAyuuvumGLY6y6FCsBX6tHBa2QVeLA47/vpP4TVkXtYUZ1SGPukgtNTkSzQPXkH4
CNAD5OBDomtdxM338sobJlCOcOySj021Ohg6zIUBpK+VbDy23qKGKNUXx6AB5xZFVSrZZ5oEFFqq
cpX1AqRUjMPJFfRcSJovp77AHCaW1wyIv7rgNw3WSkf5Cf1f6CasrW/kTBIcZ/knhlZ+ezn4Vrvx
8tTE6XNS640cf5TrqaoHJQG+QAEP9ZVGGtM/OamFozZ7yCEmcKLmf6PfjWeZBycAoFSp6xh8YV49
AhU9PGX3fr8giSeo70OQQutMPdavhVue5Thjdvh7BVj5/B+s7KcKuScvO0xRffvT0dY9K1OO7Uoc
WI6GzsSWd3GFMXjxZEam8OzatoZ1ArpuAmZiFgHs49hBicjJE+ro2qgGzlS2z6liwMDShhFfWnUF
zph1FH89FuXFBJLd0SV6xoDWfPXQOo8K1nSVF+tfQyAK9XCtFoAMgqPsRdW/i2oW7/wNtPj3SUS8
0tJ6J6CAZNo111Arscrug7/d8si4G8g//T1WbkzYtbCSQYVE9aYXMeqHFXFB6V5pmthJrR1fmy6s
7duDAd5cuXKK7fskc5obmE+djmiugZM7rlF4L33rsntAaZ19X7/42ELuVbSgKmHahgrRxcEd5buF
/Lr8QfJKxv3e0Am733gFuYfKJSB7pd+kN1aPE2KAUfSvI8fl4aHKyzr8VQcIPr+TtvHAQ0CII7xi
AlvgMF8YR7Lkl0UwRhKU5BfOHrKEx7IQolZy4sMp8uTXZezypu4SsPXPa4B3PbHupIeam4jNPcMz
X55TpmFx1R9pq6sjGEX4FbgAwMZr7CuX5i/d2ddFd8X9WltOF1teZudXZ9dalw8HESw49L40pYRI
Y0rQzxNX7Xn1gQuxtOWhvutVDuJySs2VczICC4GZwD3wTYIo64x2z5H/my+LX2Q6Ff+alliA+Ec+
aYtuMSn9g/H0HyblIZqJurWXvPDAhLNqT3aZeGh93ELi3xjlzW9kZrN8gmUNergHj0sl/uJEhQGP
AyVmHZ5qS5V8CAlsSUecQdACDvifXvJH9iUgOCY0WIEyFhAyZB9UO254jnZVbETbMgH+zkHM7M9j
EsA5YtCvfqt5/h4Xt2qZhUEwOFjcPQ4EpbKNBrWPJRx4nLbsuv7/uuvaZh71cctdwsJKaB3dlMtr
gODIg9I2NdFDVBLJ+BvpSKg+mMJYHLo4ZBXszgmr98o2iXawrwp7vn7tJOlkJTH5CpO5MLauEfwD
OPmEQOWxA3mhWxGrXBODIQ9w2V/Hls3dsEGouuQWkurUGE+FSlU3oj85N5kyMF/V6hlKqvtIrNEU
G0z6RkWu0WJqlrUBsPydBVHx0DsKp3d+4OWbWseXEngy5ukdbKjXkDJzsuGr7ZRFEJK4zhJZkA8P
eV2La/uZHSxFf06mtfalysQYY6QdY07JFeQgoJjSbHNaVJj2zB1x63pQGTdlB5OAArhHcAkag3GE
3HEQZPiARfgpJ/WnTXcy70e7KMlYvNiCn9sVf24AZ0ZcEv78lyb2C+mD/dxYSWAmsJ8FCRKRRB/d
M+Y4y6Gy2Yo6pU/bYEVaVO8H3iRwi6Lmeaj8EN+xMSnv6NCZ9LKZNs1KI5TiDcG18J242QT3gRu7
9VmBbz9HxTUx0N4J2rZwQubRBmIXNpl197aJY03etdEYQ3hxYeGVfsa1g9Bvjaq9u67J26lRnH+W
98GvQenoitB/c9vk2T6qbMexpC0VmCJQmhG2G0863Z1Mwf0CLPXw+dVDr+KQSXs2HCY7dWjBEDRz
+6+HAHbBx9U/OZCGrWJYAMeZMaNZHzWyr/pDyaXXOxuFt4hCEeGVHfK+srUoeDg5gMPEDVaNyFKL
a9Gp7Rg8IZr0bIC+yB5a5HWVpJS/VUFBfOGB8cwBS5CcX0y361vBD5q2r7nQa35kiDJfegi8SPvr
ARokIhdsoZahFekyQ3COPqwsHdZ/fnUGnUTykcVV9uvgu1hz+xxBTAUUz8RmFUSA0S0OnTKf5rO/
W7EsClOfE4a8aspzJgh5LH+bt4clsZpBI5erLFrnhY54WJnvgFzsqGSsfkWZAlu08Sjm269ij3sX
TPBmNXglJSsglmAm4KmGOSuExZtak/tjeWAW4B825N5NoeGd+2m1+OhjFZc1tkFZhfS4y7M+9Gt2
a6SsPFbXG39wAuCN+4dakIoEd2ub+A80aZR8Q4tbD31qG4iAEHXQAFOjhEI8nDY+YswFibu3xOOl
bbs6/CN1ed3h1eInh5Z/ginh29NgLpCfsK6PDY3c8tiYZLrN3WvChDLTWUOLSpHO//SLrDiToX9s
66UaxbIilhHHPm+z6s6IY5JFOmbYWyP/eP/QarBZSXq5JR0txkW8S18vHUXuYwS4dM3TyLpRwU+u
kwugC6l3hCxjmBslK93F1C2LMckwlnQ+SQQ0bOdwbTxzOn5m3arvlHMzpj220rvEFZTENl7Rspb7
2PHLRTzlGeGNF2ht1bHvZCu4/2cNcYbZ05zKKWGdv9GkaZb+gheCChWirY0JWLydOvf2k1UBcx5F
zWiRzGyaFA/UHrZnYPtTyD9Ymgpd1983L4HB7tzSD0ASCSQeAgQlN8tlkASbEe5b78xvom2uxg+x
P+g/VlOCjUOIECVKtGUqAS6nxK4wQBA0H9yW/yb68KoUnyskE6BEkFINIwgNH2R5R7dEZiu8WSkE
Gq0XOeQzrlsz+llIXcCkApygi03nvUbvi0lbv+D/MEQMu9OJkbPP0GYWWP4tiofwEYPz+PQYgTbu
giRyFmQ1oJ0GlxEt+32y8B42rkQrunbjw0g2E7JG1/A+0xNJH2X+Afb1jrDKl+e6GqxIDLwjfuzI
if1bDSSjtFvXMxV7dBRogp2EwODbzHGeCGzOuiKwKAmhUC4R+OAeBZwVS4QyIa4ykeEX1tIZSACy
scUbAxU5p2J8aLmDsnaEr0xrO0FGqxnMAp1iyUQJ1NQLAUvVAeMBNz8Y8XQn/wDELYmDKm/ObmoR
ubs35vYWHH79BlFLnVlFDtzigQ6XijeOenk8tQ8yVRgA70mAAG5NRwuZYHNlNIPja170/G3OwkbC
jJlxQBUHxyUNaJdB6Q/N9DDJne+qBU9cvUpgItKpGc3BNCQ2NpvsaoBdF2KCcrPP4CdJcv2+4wuq
UQqtYkQVhLEdRMKmjyVQG2yVqlyRZrMIFrwh1YttVJi1KHmrRQYAVwbhqNuHYPwDVV19KNeQyxvS
CCUhJt0jqkKBckpL8r6UMPUiUKFnI+4W3WBkbMRkjEVaGUNkF9ZwHC+jOY4DHuGFi9XLIAXaHD9b
mYn0VaUHV+azNOb60yabol/rRzKLLebB9bEntqtSkxcI5S7xwDXQEeuUzVvjUxjYqOMUXSbBElka
aXd9cJOgr/6xL04JjZ74AGeIrbZ8pJ1eigknHxq5/nWueTxymnY0EqjNVKFi16iQuyECc/UsFaOb
Ff4NZPvZ/f6jzM4OyJMe453/1oGa+2MUlGd5xwoRmqTe9Jt6FJ8O6pvlMj13yO2BbZWRBIOEx3To
yXYAOEZS6yepvRmWY/BW0emnXussmZi72ENpurJ3mTultxfEKl7cbM5/TR8La8siYGk9MlrM1ZhZ
Ln9OVqrW0TLaJjwiRt5pmaq2ki7cUDdW+FG8+EfsMAU2lPQW8/GJJYKtuJ7vuSovkBK3X3N4K0KQ
O3RwHQuBX9eOky0WgUElDwhI2BOiz/7QKLZ4xAKr+DqjlYEI1IoFfMr5gKKCmZ79lDNQMUSIM17Y
tZQaqYcr5ibWURNZdq1d6rCjnkBY55CziAEW+f9QSfHshYcLWfYZ4d6aKPC/EFGCetKl7Z5JueEg
CrzyeItzBPSt9V+EN5AcG8BC4l9afvMwXO57LLMKnuUdV3foyVGKJ74kfxLx0/9+5imPzVR4k9W0
vTkBftUuCUHSARJL9Z8eBHg33o6zXtwlcENAf+haOVBorqh2Uath05bYhaj0+xH5dr+fVHJ3bdu3
XZhKvuFgY5TfV0Vz/t/gyJ7/BtBQpxrsjRHuNRW58Z5dQOqn0OqgPRwr+PJ+nwIwjWzx9IFar18f
FrwuVG2F/Rv658sGAY6ntVBwvBI1PxZIb7QzxsG/fevyewR86aaHT5xfDw+gM3bj+8+b5cCJAiyC
fPPYZJUkAq0RUL7fzFIERFjCD0W9sgYOygYtiHm/awdSfXNvacGuPrwgh2JIU/12aPw8S84L7I4v
QllYi5uFXCkYEoUPoh+lOnmj7z15S6GUQ4VPDbOoakyh2+A15TH0nsOqa4jdO0b2W/qs0RRk7Bx8
6QK6FpM/2NwVkNdrJ2k876PE+v5C6CaLhuDmgh6YDtLo1+BpGfCNBrhVcJoLSiwfgD/Q5nnuPp5g
SXKlK0EA29QP+R+dSwhaCgtU75TBFX/D/kwklo5f0KRXLJFPycR69ESrDDVPgtSX7K4NsdPS6A+o
7AL5zomwW21hQKhHtrvyIMvzs7MVmgsON9MpJXmDBRKv0hBWJYUs0bEE+hcrU9p+AWz/BVuoQGeH
A/EWKp2/9AdOalHpXv/29+UIEJ5MRMXOzuH+9Wfnhp4QbKtYoyLIIqZs31vXxAG0gEI1kYj9esjT
qrbmb/cdtZlWz63EXpPpHeKiyshHIO9/yRiKVDpL3eAY6vC2OKbm/tsWwzTH1b1eYOGjkK1X5p5E
h4AY5AXNPeurX2GxdyaM2/90V1KdpJaVh/xywAfK1Q2S2BWO8Jf/KlFviBd3oUWUX8QR2cI+JIy7
DlyCQr1hgVCvk11IX02yFgFUzRh2dJ7zTMI9G16TSJF8axzcaC6bOx5gzgTFeH5bFOZfyZoT5nxA
dY557+fbrzzBhc82+VSIhX7Zyd6QCbpRcweUzjB/M/qcTxrQfuEJ2lIbKIvD535LiSrmYyS/bE4g
B+XjRXQpmzs7zQNqbCSaMnBxmOYe8Kc5UqiucX6hrzsqmYCdRw/qai68aV5n0F6ak5jQa77LtKZU
dBfcqUOF+DN7kJonm9C24m+TBHyrpjiCd70Er0SbiZD6SvaG3UeHgR6fyA2zfpX7cYQ+UfEWqs9D
k8268kEudJqAfbU0tZMoYsMb0CffKAd/+XkbeV7UgS35Ds4J3pHZWAt1aodL9U7SpNsmzPwAMmSY
kaIxWV5i77ceGwFpnmzqaahqaagf2H/1T0rSZ9ult5oUpKkdoYn6CXaqutZueDOOhjw/B0OsvK9O
vmWQCOp7vObA3sXhRX6Y7NinBDKqoFqZyF34uueSJglAOl0JUFMnLorHUfVCV/EJalBMJRHWICDR
rUGxDfFOhZOzu5ogRIQ/Y719X5jx4GngFitmDIQMdean49J9t2pLrJiec23MftlYG7gqVvE5/h5e
y5VKbaeRuwzjVwyuIsOa6xYoHghfO3EVt2y9UhSewN33w8o081oZ1fnY0/w11y8yUuN9tyh/cKcz
/C7E/1K2sflwnAFK6ZXOYfUFm2/GsiIJLk4UrQWt8Mv/+QchApn+FQ4rI1jF7C1rdp7Kb8uwS3qt
evoLWt8eZeDoFV0+ZmEu0k8gNyfvPrjeYDB2IEOCOjB7WvqzzloDRftR1WTA3ohg1k1YSSmjghdw
247Us7dO1asCGfSFyt7E56LyBWKjT/sfe51mDQ9ZNd7Q3vebKT4C6QJv+9a0m7+OiTHgJq0BRMu6
utwWHPIAQPgIwOwI8P1i2+LPghexw4qB8YFDYgrTFKO89jkiDQTaziZYnmAMDrnea7yeEc/9li05
UtUjHfTbVjPGiBMwHO/euGiDPgojJfEc6jvRMY4HefY3e7wAjQNWqAbaNPPBvhyIdEdSdcG+cvcO
TNxJCHkBmIS0m7Xe/ZCkwqBnHzV0Vf0u82ouTqU3/oke0f1B4EnnoKNp6hidCZdlpxRq5s0QK2uS
ZyB8LYYkzkbQ+EwoAXPOA+puVG+RB0mP/W5ZoF/0X3YdlxmpuYqoxgQgUz3ajwbiKmZrYImV7rDk
3FJBx55FCKEVZPEy5n2GXGKxQhgdK7ZlXAwaMnI+wGRCtqRHLt7So+jXy1ffSZ+qpFx7/pHDeykD
1C1KR7tBaUU3DkB+N6HQO9vfAStTPMGn7SbcZNoFJe+uUdxhlOHGG4aSMUzRx3vzpeNd5D9Sm6n4
3Cp8Ea1ymd1TTM7bYlts4znlKIzEDZC1IqO/sQCOrTW4a9qlcwNcjssZlJEXXwq6u1VZi647oy3X
OZoDFg0uBZp1uviCZcObtd1f6Fg6DitXtyUxJFummUtFbibwpTmzvrKVhL2NlUo1YqzcSj3qFlAH
J4tHcnqiRYq3ocACmQPzt0FKfoDoT25CvFRiVt4+Td9y8ZnfWkQ0kPnPkzgZ+aMInL3ySSobCMEB
G4pflHq2tPC9h6tAASeOp9X6SoiRGCtIezMXSy4r5DG7XDsStrjCuEg7s3egLtg/kyOCXBUFk/2F
hP7RNnM3b4o5cW1S52B6J+qDzlWwMsrEwfioageYCzLnHuNRRvqe7/iX12SO9+OE4Yi2vEkV4e6F
ma9GFv0GtAKoPhDyd6Kb5KadkHRt5syaqKIe/t+IINrJ2HI5DGqSIN/4UlW1D/vjbbaScFAmc6eL
FyntVU1Rstag/EDYac8kJkK+IqADYdJZM9B4MMkvlpKSW9/jNGKfyUv0WPBtTeZf/jalVKP+MeHl
H2DBbfiFhDyUlAx8/AW7rFBT2Jl2x9AZZ8W2TWgsAXrvpMLAykuK5UqljF/kAQU5tCdyQEOAoZ2t
LGy2eBnCo5+imaA68wDy32JgwA/8mQnRpP/2lVzSrNHqMCVI6o8SfTP8wjQxzXMU7xLD6RpU2Ri2
GHhN6sDqT4s7E+6ba1NA2HjAaiUp9biISIlWQznP7T548c+jTrmHiaVxWYRl0Jy7f85mMFt8wuZx
xi7bG3Ab/29v2oVYuQLGPo5dWQbxPFwYlBUws+l4fjxLWRvX3+/UlxxVSe8Af5IcPHqgEZr7hXc9
siosY9SLGtbOtqQWI1OQSCL1YnwojczLTLkmpLKSpXShbrzVMMzQS3TTmddK/4TZPviY/I5B6Elg
/G3s3ARil0TYMRADXt2FQ8hB7hw0Bd7wHwPkG7QPh4ZgLKPUJrMlUOH2cFNajXd7F0QBpsOIT6jw
ZiJtYG9ubWldvVcqSECx1hPD+0YSsBEZNGZWgsc0U51VH9Xfz61PAZTo0iinazYnKXXoQg1q6X1c
c7jrmhjgklngpM4KSoir85jil6lAG6AtJaOf4jfsoQrIQIPyRG05iy3bx6lr6vnG9wh1JUDNtDDY
TsBNM0/HvIrHGSacWh8vK4foE/JIN4or0V+ALv3xzjq71uB08+qUWAFr0Ci31Gr+uUNMai4yilja
bjtb4dfIpLDEWszsQjfveisYkcf6iq10wOozgI1n1a98Fzu3DRw6uuH/2J895feYPKIS1HCYMjk1
7JpZb1wltaw1dAdDRnqsVCEjzxPOpcjjM8AYoDh2ov8mtSjTzxRbqXwbkD3JH7KRUJBt50UQVbWW
j9ZhEh/OYTpY/yZmaQFmmw4gMV80Y6gRQ2gI/1SsY3bvCohOL0qm7Hpbpvow9u4MwQLTc9sqtah0
gwV0KRxKfbq3PAMNSvRJx0BmlYeYfzYK/GG+fS8BGpzS+LvRajZFPDaoytGRFSsGXcC0Yp2vtRy5
z6zfXs5qzsazL6rsIwWaoWWCawEFmM2W79SUfiWYN2qroNsw05Jy590VfAc3yzi6KJW8eFia04o0
ZtssXBSdLLhAYzfnPXa4d9YyHoMdqEmMv5WMlec5K8N1Li9EcuYsvfYC+Cp9QflfFTeN8GeUYZE3
DXEDHAaDgjOz5xzPz9cXvjwJDGU7X6HpTYx0AglaxzhbYSNuSbrn1pk9gVAuiUNK6oaLGilUagYA
OgnuVoiuUfwExw3w03f6TSciqjG270+0/yToXg9MPFEJvphKMAmfPKC6G7OhrTGHvQaBuHQSCHKp
ZL3y/UCNz19bo6PM3q+xUEXlskQ9swJhC50VwQOdEY8v5eHfqXk5Wn/oW21+xnNu2egruAGHiO3y
RNRmNTGEk2EuT9aMQal1oJtgy6aIl2MmN0GXM6Povn2Jp11nAehI2IzQER6FDGyu5v5dcUGSCXva
pYTM5uSZVOlZDL4Nq/yK9Y88kBc6u3ExmDQGxZICUpzXUtkgN8z7RGHKcY4fmpCr6ezq39zmrwTS
qImNwGiYcb9TwL1A7Z7HPHXkYlK2BBqla2MEUvxhG9VyM6SFaDfTpL1s/IZFzzPfroTv0FANfUMO
6CZOKH7EFZFeLlBX2zGQrOxAvfTeXuFJsDAL14uXtZGHPzGuMaJReec/yG2NJf2ys5iM7N57hLvL
M6RMAE3+iQc8W/BmU6WL3m8MTedJecqSBIl84cS4pM5h1PGPRu/QBL+fK96/cnnRhvLiy7PlTtdk
Z+zKuXrzuBYAtD97HuUouWctj6Q17uSAeHMlYqmfbY1RMS0Jq8jNS3+Q3067kXnVjGiL/f2RA9uB
aDH6mNYQEukOfCS7q1giUXbs0iycRlV2xsrbrZtAvl3uVm8eWCYHVHt8HzQlC9BwmilxiEqlGRsE
GFAbCtFL3ejeHaku2anU/jko9EUAK79uTqU07KEUtdxqMKrg/NJ5y15UpwVzGbo8YWLwRNs+8W3j
59u81ntxrIh8DZPT4hItYPCDA+7EOB0RzBsDS4GALRFoVXStNvSLoazTttq1Q+GzjxxZor+nxL2j
DHrWdMBLmBrGwzZhr46J3NJ/Tf/cm2O+AoXwZZCtyjNaixztLJEU1WrtKnsNMga+ohDRD2aDslmz
G2jFae0IDIDsCvzjjeY2DXQHBHDEO0EjfRT/8Ya70XE0PBWxcBtnMPgEbm9mOL5E/XRvlag7PE/T
JlGB7HJAFor4Hd5nSxEEW3XpugHSL/rpOBO8GJeZXy7wR2nuLGlFFA73BYwQoTbnDnBzPWfTBvUD
HH73oB/lmtiTKoQz8HLQXKPnBqks3QVBxKEItSQbjrR7sqLVndI1u43SWD99o1hR27hzgYuZ8xcE
PnAbBhH6xpkmLqgify/EgpnY3ECNM9RmViY0sOh3kyrlV74GKgQEUhiTBUoDV+M3h2gETnkrOHW8
3hv9IGID7vcJPPlrhGAdhMa1o0uIpR8bUGqNDrReMQD1xtDPoFSToUZChGU+dQGgLdxL7OXj1VWe
Rz4a5BqimJY+W3fyNQng2beGFvo46cACtwdRxzsCNlLU1PKyQgYVIMIjT14Ec0aDMAZvjFqYdYgP
4o7UJ7fC7DiictN/UM4SVcvW9dKPc8Cv0z5JvgZbdztY0xF3sdq3uPkajPZDX6VKq1BDAZkDML3r
OB6t7AQVtA9kPenbsi5NA2Z1OXd+seyQ7l5kjt+h/zWIfeboYb5z828M/50v7tkOXlTEvh+K0bca
2GO/lDPWttY3cvv8MUIIbb46+pC5zHjCpyQqa4n2lVJx01mWd5JzONXufyxfRelmnZRb1l78tO01
x1dCF0zLXpJNRonZt/kDJ+UhEs8u1I96/kyulI9ShFgjzLR7pepVm4xSFQRbp5clmX3ah7uUB0++
qkrMk+oWcI5X7vI30LKct9kyGHUwCLBsCmaclyOutGztS64I78O9pqiwq17DzZiYHHLUobYIq7IF
Yje0unA+W9Rlqe79sQ2rC5ibISYyoFZ5UE2J+AYLeuBnJ6Zj/nzwvC02iSpnDXGBCRY/IwT/038V
WnlllncLU6RXRrDj2dKrhaRsxV40+CiWDNVheORKq5LLxt3OcPKolSQkNCWnACfG2SdhVtCMMAGD
CoznfmtLwF0I4ZAqrHShqDkjVd3GcadY6i6pbceyzRhdGGn1nUbrRqNmhRtlpC1/pv7kFxn1JiHO
bhwl0pgAkIfedfgq4Zh50uI12f/3JuyhlVqXLsiNC697/na9QH7fjhHCnK0YvkS/ZNao+5Em2Tg0
YNH2ah1ksCRg+sIUGgC9KKJQER+zC4buMFe+WzmJCy1VIFqf2Q/HLLBY7HBNt3rldoali/j5GuFh
87lyBeZQabil3PLwDCl/u9qLLREeOiBOcDhupeBhC6yoJddWXcWffgvmm5C2Es4YDfyHRO1P2wLQ
G2+O5hLmy2GBrexEPUFuESjQEzsQd9YZUdZIYbI0OlxGBuyMYM5Epb/BxRds7zPu1j8/Fj3rqKLB
nEH7xWOpUE69Fl78FOyW5HZbZHz/rt0yRYMrUZBxTBkSs+yRHwpl/a24S3N/1ptO7Ic9Q6t4bgAZ
0PPvuIR/YHp316OYbfLlRT9lJ/KvHl20XdC7oKn2yPI06UFuOdTkRseRjLyLYC/mysmai1xHXPzO
p/fK3ACPN7oB71V84MFDdr1ZImFTIRCN6w7M3gLp54ZpI1Pn2aHUGDq/H3NhvynDa+dYTSFP1PUj
tfNw0p/4qhSIcFQvb5/d9L/zLiXBWCuudslccGfxtJKAndb2qjKborrywJ1XJUOx7MnywLJYmZdx
yDlINN7CnyDt5YE3QWYnsxK8LUEbEqEsrYEQvpD5DkmtWIPWha793Wozi2/GiLoOybv/I7I28Z33
1oxoVk/SUYbBu4AGB+6ZS6O9z0fHRG5IpVQxOh7NKsFZ6CENjjX3ksExahQmSsWKoUaf+nfnUGKF
56+5DAsYXdp252Xa7jdyzVTgwCp0yOignegiCF9C3bS/QvmvlKsI75bNmN+mcIphgt5pSJkXNnxt
3buLNSGJFreB4/3McN+LyOdQHbvwgzxB+WZnfx8MkylyhydodEGFPyjGl+QtrwrMGo2PpgM9hBHH
rR9N0puQ4z6eZPYERR6793LZJAnJx6EkwnXvGT933COp36qIubfQzi6Z2qqP4WacNjM4hrYdy/eF
L9uulV9ZocTpj0nNNgoNzejWgsyFwobtymLTeSgCGU2V7TQz3cnDwro0w0xGRbY3iOkRE4hB6+JV
UA/MCXO665j/8Fzr4/rn5mo976hk5ZaZJrXCfB4vbuAKJ9t3bjPg4bQk7WaptYl9pSa2llU3ON17
iZMXC8Xtn7MtGgWEIi2KOeMQ164UX+Wv3gfYCze6Z2uBVR+FzkMr/61QC0RkPiCoEqdCLMQUGmsV
wetECVNdPffo/vlhohH1GMfltlK9QL+v4yt9A4OmJAers/tc/DPpIQQLhVKQ9wl62WAzw2p4JfHJ
cUPPGdHF73AEGH6cOi7Qsiftng71u26QWYR/SfdxL5PCb5ij6C/91Jla4mZcetehJnMTFMz3RN7D
Exn3GTGwmIlgNPCnfKfUr1tJ/IveeHUawtYoYd98ytRAkA/a7JCgiwGh+UBYB8VuYfIYEJWqvHar
vCIHQDQSo5A1K3fZHnvesM1d8TqAS6LUElxPxRWVv3Se8jP+bXVF+xqT1Y0rBsFKAPLsebfBdkBF
vtUWqGd0x8B0k+LcZbLALPcgetMIIrARP5QSmL+/EI04SbNkpscklZCKa+CH+h5X+PQ6DNeTcEev
KonLL/gP4Sf2WtObl3RZM6jkHHMjQ3ayr3knKXhTl+RpZyiD6uH4tsPIPj+C17+QaxsqmNO2X+9t
uyu1emZinLEgbgBSVNCnYeWh6fd3aj1tvhKoW/k5k11mCFHI/u1cKxoTxBAw+2YLNibV95vpc0lV
BIbsPK6m3HTsfBcR3JlJuqHubu+c3N+p9W0Gnfr0eMspBi54ZWSj8ZXz/8bepO5Psf1yd99v9MaL
BCVjI4qS3qBqC+LmWAot48SxoTI58pmVQ38P1uVxh/fQyQDdPgpmkmHjgbaYemWO1ql8D0XTFRlV
BtaFuQlOED+VfpH73Y9C8ydoVr1rikHfJT3l9MzfBN/HwrAc1XtYDyyEOcPmCLPdlNA8x3ehIv7U
heb6MPA+25Cq2C3kIVAvouR3ATBvLE56qsdBD4IDx7/EAKsM8PdG3LnR5AGmmio65x98ixgZcaHv
XfR7T3Wvk0DezJ/8SusRyHiuFPIO8DsKBJxZ+7SKWvWwh+IyX3Rys8CCs3Yf/Km7t9e7mgokt0RO
uZHOENhw44dE2Gb/GgSrTq5iOgejUe8reyzNHqiNUOrLOWghgZ5Me0jEttF+qoepg8eP+yG2+b82
jDSDIeucJ1RrSu4PzLHvuK5CsoV/DmZrLHYa/BMyvvmS5vKjtP9R61LiPjeiAo/gkKmUfk1G+CRb
IvALxLSGhQ/p4TZcmPOFlf/cJ6bueHk/sdy/TPcI4vQm20n8mO+GXubu9KKpB6DGyIidCt30+bWr
zTnDgmoJkCz0E2oNPX4+o29WgsMGwmofTvMxIiDciEpSAAFGbhLCjCSYNbX366Hutoh4/8HlTc0h
cmV0x2Sz6yEFZtOOgeGQ6JlAoFBpnPuwC5ItZ9xuPqkMYfHFgw3qbf7g9FkU7rlMM8jHcM1HhkE4
lq+6RwY7zz/6NwSUYCPgdT489bkhuGaDaDnMRSyMiPVnoYbEskVJZh5BdlWfr74kcJYAhnOo7jsi
NiilnZdpBlh5B9qKhL1CF/KksWm+c5PMV3Tyqkl+0SGOlH3S1/qeJIq6v33lSttAljlql5uKxE0i
Ghr/k5WpeDD8irtZfLwlIQJyH2AM3M8YWWwU7FRmKUuhh+xkdmK0/DNt5ZbZkWESlOA0voxXLShf
UEX1i4p9zkEXf2rmbbe4h9sg9vlwR/w5huCZwhm0JFIniGUXUBjg+TuDdjl2BcVMFNEnJXaGeoT9
STCGPe0Sja8z7ziM667/NpBIQDN2na8BHkHEtl1W0P06j0yv4XecHD5Gku2Za3UzhbGalwxivqIH
stH69hkOtLMOkHXPJaT32uObP5TWT7H49XnqiGpFH4DK1VhdFCUD6zPY9F14jevjV3EiK8+yrZBD
lK7EM6McBP5GAAKwmRntYwaXSdlWMjTLI4PVJVVhFlDxOUJdWzpIzFgeG6G1frR7X9EafnjywtWU
oTorkdAKPCTUQ9daHARhBKkmiOiS2OUE+frSs8aH/oxHqpucqPtn3P737MbVSmfFdwbK8ueu4Tym
3OuHpx9YQVxvFmKzq0rteAaZp9tTCD2I6AUGH6b4f2+FOycDQ4N8YG9J1+ecc9untT7N9othKtyg
+JcOJOUncJ4ae+gZcVvnR2t1ubNiVBpEs2v4d5giK2xHBl/5nQMNr75vOir7SEllnsS4r45B1ubx
ezqeBXmil/P5h4gxLcaPzBWhycLTzAFd/R0rcKEnGs6ZxdjJBpbXp/DNaFZap9I6QUu+4Urf0QdX
KEanhSogmpNO2eDZbXx9usESUYvCZwk3hNVETnMycTdkPQOazwHVHZx2KAMsW2GMXo2xNHb1N8im
S9l0JF/2Lqokc6mVvNfjMS0olHTcyoLM2p2DA2AJ46z+vkluOvDZhlzbsMc9Wx5wQUWms5Oh5yYQ
3+KbDZwcUhYEX3J8Yqc7/gCWRPkzCxw1ij28/BXLzXPSyceAStivMIOdLW31bmpXyryozb2SEV1M
DUX+wqBi2vvYhbdOs7WsZfEMhPf2GIcuW9rTt13Dp7EZ9Rh5CMh1TwoIuMnJx+l7FTlo/a4FoyaN
MYxnPo1eNrd18EacsVEQwLB6011Ok1NqDbxm+1//p2xuVMoS9aoV9yM7dsVXUV8n5zdUcDeg/mlQ
dRXNVif9znDgPjGvyWWSrao9DM0JzecKtErYNFri/REsVVuCD5ahdl/8YQu/82ku/XW7ubuQEc/4
94gU7Sw9GtA3HZdJzw/E5w/JCZ5s1VMczzOmbILU+FUcqWEAwKirlBz52FscDRNhZrOk4dXoneoU
p5bhZWFtGdiihKuNoOtBLjrM6uO/CsaVhKq0EdKt4srrmxsp3miTa1VSlb4iNSKwCAIgsFA6ckAY
F2Qh10jVS3ABCQGgIetUeLyRlTngvtGHRLe8SrZo+WXvb1rysOY1Sfh+8JlUrhBg4kVwMYlzCEkZ
Wesu8RInevlnel76U3HNA40xvF0j00l8SDvqU6dfiUphHbiqUfY9qhu2awT9XCjuCy8JWBCNN1fg
a0dB6iq67eALGbvWXSik4wIWKzPY5N51oWcnBfGssRy/Au/AKO09cgcQ5YtMpcK7bS31WH4mMqGU
z/FYcUUNSXIJa8Al1RGOEM5XcFoPX+QSWE4ERu/c0NQNeo+LIJzQWolg8LHXt4VLiVzmK+QL84iv
xru1AfRIra47YZ9tQ3Xc244Z22Yn0m76rDxfFw+91z9OAE2NWc7xdFsVop9Bg4dU+qn4QiD/sSZD
8tviDQrt7qWIUFi48U3alzP217DqlIAU6ws6fTzGPlXmnkOoSbfvtZ8Sx7P1pFiHN++QUnb38lRS
2veiLxGAEOAbJtB9fAKAXzSBVf8Hj/vpDRyydbYk2RVAP9xcZM1fLqFpBIu5W5+QQGfjlSoXKlvU
6ihO1ATiQ9q65DjdeS6pCRtjrl1LAhV7/SESz5Lnn5AszJ0zIf9Q3C8jsjlJopZqpPnPDFhqKqho
GzWNOV6LskbpQTVyjWAKweVKYa9Q4E++uAzw9UrLDfBDeaEhpPrgRxhjf/iMTtmI7PGbBzwu3Ej9
2HPYfll1AYM962mdFs2wx0ezez85id4hrb6XsrIEleoVLyTAvwwtXKfVg+ykmVeEypptQIsNwjt5
wC6H4UZp68C9arf1+k7HAkmZgw5NJg5insD6MjImBjr6Iwcm6oRQB5EyQ9SONmtj1+CkMDLrd2EK
IosJ/Lo3aHXnnWKrLgMVZ/zjTNNvrGmFsKADe58iLCGcbiLSB8xXZNs24MIJn7EDyNpfBr9aIXxC
b9dz0fbM81ksHC41n1UT0+pKQxgRw70q3t7ICvNY+2jW5odflsyVfQsmJWFDvtwsuFovmthOy3V1
y1OsA9qmg3ByiBeBJTAeeTNtsNUT/jN2yt6jTFca2JIPsuW7CUXy7ICUsxMrX0DZQXQye9zoM3x4
qpkJ/I0PJ7iTy90mOO0pphv8NtXUn84kVfXeX9ne3tNfuQHUEenpBA/+n8a2nK3C7Kj//9omkIpW
Hr67wHiQ9+34o360AuDzIdxFGExhviB91Yl3NFPvKHXn0FF9Elj36ZBFnxKEL2wrgh8mC7CcJeUm
Saor3r7LlIA5IA98Y+yP1jpi9PAtfjlElI+3BGK+SSOuimbI19/nW8tI/O5RHAmDW/yLmTJVEb3Y
09+RXAniJN19txF1tdSqPbAk2BtrvqiXxhZXq1wgI8X5AbkOI+7VezsSjfP+09O2vRsJ8AcOpYUL
iBtH/zVxCMjxZEq2R7z5x9VXyofDXVuXr9emN2/l+T5dhblh7VJzll0A22SXT8B3NA9L9lgu9UVG
Qr2CDcc0aGeuFrpckVvIU7pZkJBnhciqkHCVOqnBwZy6K4AC2Nmokso/tGDaEk7kRHjRGEc8jskU
zmIDutBulpJTGiUmvFZMpaEH7z2Ppa/vawCSUzdAjLxjYpPM0LaXGYJCNh/j0JoPqJfLfRVnN+hU
giw7qRFjAQJEXUgn8024NcilKJfImhPEv1L0+qbNEfEbRvXYh/plIm59gZ6BNXN/10JrmGPUEvoK
BLgqgsesUzcrGMXVUm1xZkEreXNozbgMYigiiuWLk6XSqHJTaTIjbtguRJj+GPgAl6djXRIfSyrh
JoCvR07AKzShB1YxWUtdTdKLoABKp39uvUcZICFsj8dmrES/+hwYCGkonxum3FiBgav7L88favTn
oELE9mMpfDfBSVB38MWRIRUMSntOOzg0spcKeMRiu8aH+hYdhQ9QOHCZn9sWFoaoGaDMa4SEpoif
0Uxds6ogYQUG7rzQfHRAe54UEO4Xm2pME+y1cE7vBNC4mi9UzYS2obNY6DbgOsXnw7oCHQpuDeN9
x9I5u0ZBoDt08iwKfxby6I51vTcKFYewWnmpulC3DL8R90jrUkrmvNDrYSX6IbuB54ZbdE9iF7DE
8oGTpM0vsZf6lL1eyVLls26CjyJfRmJXjN25UNqCkEsjK+jVKkqOWefHiGOAEPuO2dC+97oh/GJD
VPNQKxTVXxllS23k/SSdOjllbSzyuHSeC8UiEMax0lruQ77g7M1KeueZUA2AwLFAsALDarrAKOwv
t6qUTl+qKQ1wSSCId9JYVIVUsfqc01wvUMLYqysKk6ItChZiU12F+Voyfd13jW9raTNXCMiCpa+S
CwfQW5DwzX3rNwYj7DAdU0ECe+1nMfnd7S6OufGVBR9Anb9kLrTHs4wofvs1NRereIuJAFDA512o
B3K/K2GYT/OldeFAQmlehqf6CbW1Hg9gmf01P9jYgkE6VSKI1HDhpwAGmbBcD5gaFt51ckrOkeqp
bY5iKX70387LfirUjMzC+WRs9LQxX+2Xi5uIZdVgWlB6z1N3MrMg788zIImzRBy71YdPTMQVMY1/
H8AWA94Qmdib7j2dKhB6Bxa2uQFSi895J98Zg7wTmaIj79JDm+qx56vA3TvaPp8635r43lVC9yzf
wn/nSFiZam5BsS1N6+MMXrro256fxjOP/zQJ3VYY6CdZ0Ri07pnd3iXnS0Dnf0Wpsaq47ANy9/b3
oBiysXcfPkmgdXfHQOTKKABtnXKSDk4QypaWx+iEluSWAmbzBqZBHpfrv6RwL4JcMcRqOkqNGqal
tWz6nhGZ+FO/OEkLUHUPLfHl9OFj/rHwphOTIl16rpeOxMN9bmmMI/UqV8s7Pc07+wDAx7fuTHMU
zpHSSbGXR4I9iMEPo2LyHdiJC9w0E8ApiXHlSYaUKIuxBvEVbFH/5iciWmvx84qd6Jqbvi5Y2K4W
CQl9KIp+mqNBlb2I/h+CulPVriu95YYAv2k3Hzk0QlkW08vuMo0bMV+IftOXgn5wDd3vlOKo3kta
2OHWV9IbY1CgYvN2NzZRr92XG6zwrhwmmfwgSgx+ZrcEspSFXdEv6FtDo7iD7cRuBpinGq8ZpTPi
ejLwCdzF5RwUgQX/TYADNcBNxDdLReA1l/IoRdO/ogvFFouLikuDtaZAyaebKbuyIHkYFZiVWefC
Dr/8r4Fg7JZa5ATv6qK7GtdrwCC7V+Rc2gWrn0/YUoC57M2IrXY0AHHnhLqcdfMy8vG135qsBIPc
IlZJx4RbkLAycnRoMilzOpAOUMKHy9dwUQurUrwfJRyUoNu9V+6BD//kB26sYtgBey6Xr3o507Gj
rNOEodmmYhIFJ9KHKE9HK6lnKF2OKHNMqM1TZ1yHaSxN1Exk9NfeZDFlUqhfU9jHd65MTEEoutxU
KpO2p/rNOK5R2PvBrw7mjhkOBZrM8dOmy9Opxx2vpAO+jS/ApufUpcSa3Zm2jNP8BrMEKQaO7mkv
T0n9CR4MVYjcARlQoAneNs+RepyUc8myG1x/eWUxKsJ1DoGHg9kVP5D+XDtBfVcGAEKinLCdE/vN
3xB9xEyNgow7iaNLMoOOD+yx8jJwAZLl/6iwFRSqS6AfHY7EUx9QoAYx+Hcs2iB/XOWrsY59PxWo
SGsPnxx9YE1QHnMOBPCe/ugY9QNAuMm3bZ/zNLtBdPx1vbU08KjTnJIKA3dR5vwBLOet9oHSL4N3
+u1Hv+rp0fPEpWMxqneT8FhRd5FSm3jx4xoVU/2LEKWqbSB0AhuSGkXgHmWzYMtkd9WF7ZEuNQHr
5pm4en/a7s92qtg99Qfd64c6HWVYCMbyfaUGV5rsaAbaBAWWdmoTehcalTXEjgZeX7qGgehrRUr2
NXyEXr8aiY+Y0y8tiI2bzhS5Nuo3uVuwKctItaBsQ/xMWk2Gvea2GCGlaLiGOlr1KxftL1L2h4G+
QkwExmcRd2Kv+rB2UoBrkvCVqkWB2LngB225F0KMk1DXkJBxQ2kKhriP0nuAFTGPQDkvDLg2zVUC
215hBHEXF32+/5nQQGgbTyZ8GPpyJBpZ+R2BLfkbMoCiSM0aEaawzNN0bEd0GazTEjmpQ/4WuG3/
R78xeOf6+nkk+YlggKgEPOh9hSuO5cUbxwHnrG/d6na8Sx4YtZvA7bZhueiwZQ7Q5WsiuRJHhAd/
GqKj1bfOoLYQnNBj2nCtZRng3jEdFOp//6ePm5gjNtNJrYTiusnMFdSP8Htqw/mvtdgRmvyxe0FK
j96Uvm6Lzu60QnfP3JS+msDgks4Xsg8XbrbRWPsuYthk+azCAv0PcBgHpEYoUiFEXs8LQLLat00u
Fv+b4MMaKFz8TAOn8Rq48+yZr5hc5j3VzgJUscFhM1hhgwqWhEcm6BSYpRfSuqrVlChB5NJ7pu5e
p+ypqc75VB7nnoX5rJidzLPWxXV5hdbtEmzp2m9dEjaSo8iEd/T8K/qbA106pMfvkdZNS4z+dsKi
7RqnWllykY4fQR4yYA+96Fr/7RSGn7PFORxbqENTy6cYs/CXHOc5S7jzrPN2Ivy0VSzROfV64pPZ
JQm3oNgGhMVCjnFX9PW13V0c/ngCDTWS1csR7aGIiVVs77pWREAxeX17oEWWN1/YvdP+6WUtSH43
NEoRvnwgrG7679cB5m/NyKtTgZfysDZ4+ddNqsYeJ4avfyOPzMNbvimAfPr/Ea6KiDRG296UZU4U
0rnl3nTOdtaFg5eJ7Pd8N1XoW0ibOpcFjcFuUNHHMUzqU54vU2tDIZDzhF96F4pvzfmlYqYPUMBh
+NTOjjYP/UKCDozXP0Kb3IOI6KW5YMo6Z1d4DC3JmVEiGezLJNdoOHdZ1qjKPLeR53k1XVDUZ8Xn
g3fpM3ZY+lN/NbYiFxKk6LzXpmgThCBwrUNluNtV78JtFdKuHJVCZFiBLKEQZ8komNQrzxw6dOvk
lw8utdlu086NzEjBH/oMvpqSbLCAoSFYIXL5Pa5azCGXchfHCurMozvzH2tzhplW/B1hnJmveyTy
8RJ9ZIIjYpnBlEFrseKxGzw9sCX9f4UmhwJlXsuywT0ON94D053/jo63xsdBy1/snPwuaIDKnDkL
QxzidujgmU+eYuSSFHwr3LaWQbCYJiixCz35d8ySJPN+ksLCBKc8XrOwbXcjX2g7dT388LvbPOGF
TfQ+DXOxHH2WVCdI8+Y7M6ISAVC4KnuH6/6jI+1uSYJBocazme68+M/L7ONR4CAJ4t5Mm19E/3vq
9E7O3Pt5pS8lerMIZ4c3rC/vmBExCNskcfP06QHK8TG3YU8hdXY5Tcj+1xX+C3aGoHSRvvhXGTni
ZCNWUxvkEiSYAd2DfWUbE3h0k+BIvp44GfZeXjbR2deprcUDCFc6ol24uMdqJSi88P2FfUOnh6ux
rtOA15feYok4jMWkq+XwhZnNuwUCTWsG4W3xJjRxOPZt0vU2A68HQECgUNwFfLIDmYLNF6pAw5VI
lw1ntMqh73zNhrwiupIlznBXpwxTqEdUb2MqgkHnavghTbh23tQS5yPiB0OeQZCrP8CpmBdHQHQS
86+nVnLN3t4vAKO1PFVyddyLSNj48/KjPR4wBV7AMFNOzsH2lcSuduIwaJwx4NfmsEjLRRAzTOEr
D09TmQEU6yxCQzV8lUEYnLxAOdbLLHEYYJAUR212QAf5q0+cb6P8iPup6vzQs8IgYBFIzUrKy8N5
IojazoYjtqt2AyZ00lZ3RYZ7N5dx5jtxSyvUwLz5rx4UCf4svZrtw7Zs2+JalDAI/rx5+zS3jLaK
y2m0BqgWy2Dnz23A5ppp72WLubeao7SLcebm7HmuVypsyp+jA9LEFcgf1jD5Aa7m4OQTB08U2Hwn
czbGcbIlu4f3ubmib+tQsKRsNu1UEQ9zjqb9vdsWR79yDNISmqcDQMVUdZkRmqyKwhSWmy40fsgR
y8PRWw4bXXZ6dtnClzASy1f8usEXQiK1F/tp1WXG2CZgn8OSBxoWvQxdXhWx8F38kILnVZ7ZqHIH
x7PHBfTkklvCqhEdne2m42eEbdi9PpUoJwNkpbncE0MC92lNj3q9aDu4S+VbS8s9CmyfhaI2a5qZ
QR8DolSqX4lZh0jt759AS4yvP3gkVHoEjDhWeheAShJoYqps06DAmcpoYKSorA+MOQqpXWuaKsJc
IcJJd6oz063BwTfrrUyWfgfJQOiILRHXtzpFN4blG88Ryf1UsYMCvHcfZcb226TcW8dS1MkZTe2U
fLgquU8KLei11gm9lEawEQykwuplqbyrwSUmt5Zgko8spaWELDCmUc6ltsboRI7hH/06SgaWIOfN
1lb1ToMB79Y8qGlJMqyYCI6E18kc+RvaOj0I/sWKHr6J66VfqXrWOQCxMwqKNd2vfMcRWUTm3UIu
AzPEunaa0JkDpeST29AG+GNFnfzEJYLZkLH1bpa3i8Gc1+ulA/Cwp6aMiJVJrUaHV5IWN/C9O4Ka
cNjot4wSgg82vclhP2uIKeUNYzg2bXYMaPwm748s12TW1nvPVt0F4DmYTdqpTMj4Nw71hAPmvbpV
rmtZuPNYkXnUg2VjZGpgMSP8GP8S+XCimH7aujCFsXGEy8VvnC6qWAphumU2E0aJYclTrut77mXP
KYYUGgngGjTuTwqv3pG7ExXO7BEMFFk9x2mhdrSXerp1fw0cCKitFAzQzA4TuSHg7AERwL4r78Cq
1HZBnnXgBR2U6Ba/z7w7hhUzWeFQ7gR+aZdFu2oz27pfeWFQJrwYYjR0vNOyhTNgT+oF72VU/J0r
JiMg/jlnOwKFhLPTeTAMhWGKpxLLFxLuu5G4vUN+L39ZdQ65XM+2NrFwutJBeZCk97UoCImXR1hc
QV5t8RC61jRsvZPUVbQ53PzrIEYpeH0uvSaYe/meYHqkpAf8VWH/Vuwl+BcjNRhLkSZOM2C3i4j5
ONpkcJDnx/gmQdQv2O+6OUuJoxGH3tAG9i5XIBsEczCFImYvy8dnkLCl7c+96hV6G88J7KmhRm4j
FnojNwWMOSmRJ/16sVBJBfOUNJf1ZXmfjpUY/SxIPfI3HHrUQGcg7peLaUuqnXg+UOP6JKO3vbQk
GjpwuTmkxcVMbpqfV32/0T3ejmenMVZO+XtKHTCJwmscFzmbLaGiNFfNacTJjV93N6XAsyxr8e/w
E+nT1yMzrAo1BK6MzoVXmw1x7S8po1Vjl4J/7OUEmVhuIF4twZMBiEX6LInbQ3353ert9LiIbr6v
u2abIE813ulkWnf/M2ZvvOwh4GJfnZFLAB44nfndRk3Mf8qfoOliSxow7wRyZc7b6txxJTz8hO+L
xMvFXC51eSVDK7aBYPuRbBziw2hj9a4jS49PPkcCVJmIoQguUqbju33npUV945RbMGQkvTHzl3/1
9nK1b0oIRGNBWau9pbrlzs3GrHW7hFYuvqy+dCWTQ8LDDRPOrl3yPLTWdOfSpgClVCKXhtL05K5X
sQhKLxeG2ly2cKlyl1NOA6VgSEu/68IlPXu5HMf4EIMASv6YsqMy7YLv3H9j7djr3Un2MWj3NzXv
70WqdC7cP1QlHV167KSps/ACXyfEcoHA4FJ/STqbbr1Q0YHv4ZsPjKvOatwiDAYFelKuT9hpb4of
8cL1yRShjaHOm6nfngIoDU/7/Wy3sHtQNRIepUO+vqdBVeUTlm22cIoRpxMLkKzRreyDCAYYCJyO
5LfB23+FDP78ygrwHdqfvp80JQqzBKFShpQCZu5v0ASFerTmVdPnZf3OGZHtYqbm5Sjt7l8W23BL
D2tnuFVtuUGZRbLjHYYEwEI4twvM7jCrxVR+M1C8DfM9TRinfZu2ZEKv4oonomQYfap77WVGO6wE
VoKYI9utj3NAdHDr1c8Q7S2cWB3QD0LYtZaUXYUYnyC6qopEvEnC9RqNzE8qqPhVVJCP5EOyT9fT
hlPaX9aFX1qLc0wdlMpVhSAoPdIxDNTFAzEaq65kVzd0MqjGh1BUoNzPId0qc1rj48JQqmYibAP6
1PA/2Ydb/8n6sWm3+f7PT6xGZVCgX9aidlVQNGl4r83ewl78K/5gJSRWUswkPTe4za94Jk4OUm5U
fQkq1X1euV9SdPzeQ3D0voL81bf6qQEeDxiakiJnHA+6tOYvFW77q9OFrGPbXUnhA/pTvrQyF9iq
MXbcnM/nG5fhkW2kikZrGCGxhNcpJ0GprpJxd9qamheZrPRgrBuDSWBxJtcrAFO2iYz5yok/QeM8
/ABLSWykQrywI1E9BVI0ardtTXqOxpcR1Ub7JSyfI3FtXihqDKvmY3Kxcbyt0hpbBQRQpmrs+3RY
rCo1xJAZk3EN3XzPukuXq5l89fHISYY/pDxFVik6kuI+DprGnp2S8UL7v521Tkb/TEAmISxpfoMl
7oQ7OYp0nl9NxVRhnp3uVyOXfLcqy5JQwyPl/oPEwGt3h0XH5CV0EiIL4Jmw9zYrIvMq92Z0qGj8
nnwDkZ++Dv+LEOcwL41MaoQupIzKXMDqzeZ0KO6vXR1K3S4jNQGd4ot0zIs27AdSSrloFDq6XpLW
kI+OsFHUVJ1ljRSsFO4bvXZjDlDfOCn71G5jZpAhAnA4/SJCMEr+klby4N6qBRFbnq5qPJt7Bvgr
BfyrGBMCA2jwnivEDhRVdWYnaKS73JUHgBmcvxG+IQV3islWsVpudnN5eLHtCWU8pAZB7kDlJr+5
KaYXZD4eGXgvxCk2Sw9JKZMnaO+Nbr+ggM0VhKPTIoUfUw7jrJvDTLXp7fQfJNU/jHxZ57/C2yhr
R4O8S/hrt4TfNID7mwwezfQQRTpnJ7cdFzQAao6iXlGjOYW/MfT1hn1ffhWIyOKAlmZecEzy+Z/M
fjexRmqGZwujgigs1w44cJINQyJUZpyopXPYaMzwfABlzziA8ICqYg5ojGoIvWB6WGWuCWim1IlM
jNRnvPs0kFhZRbLPuY0l9hGa7oRndHzM99K69hGW8wVRFuXBx2duva5APQa1VNVjtfboaXtKYhFH
jeFe8WtpaFWJD4Z1B72VYGdayYZyf+/MlQ+zVXb2Kk8AZGWaf47B907IybppQvpNAxdtiO1Pw8Zr
XPGKbvfVsL2znJxy8Upub+v+9L4eQjvOimDosInYMvl+YhyMeaUtrQyFgHpxPEr4oQ0z3uEmSyef
5vq4knaNOo8/A6vUdTOk+3GYaRlVTccKbU5EGwYU5IP9wJOkcw+AEDKFflqGOrjexmjftDVfTJ0P
Pm1muOs8AlQbcDu8hlXkNPr6X8VsblHFh3agOubYKCY0wLYDM1mGr45FuKuiO6kzoQCqsGVEVH1n
VZo+m3WeLLcnCqZkBRVszf/eSnqtR22UbgBj1D9SnvrfcAtvrXR8RtOa41qLlJkz2BYPIxuoztPs
0H2k6RNtSOAD7oX++74V9jWbDmr60hQp6M9WVghN00NQZPGGCHclnVXuUrG2aYXSvN3HszxOyXzm
2Df5ZKwG23jBcrI77BllQUVHk/lvMZM/zT1YnShF7fOA8Qd5UNvHB2bOR6pehUhKx0/+pSFg0GxM
RyH4ixB3Vr3oZyFmaIA8ab/+mMAQ3AFzUJzlxC+Sfb+xpWxOUQs5l3WFY94qNFtiAi0+CE4cJUNy
DenYhjeJKbdrQcCJj86mlkQ/4ErwQ9QDPTPPPdsicsJvZJ79BJCKpWTPs153IGSo4515YohY96e4
VrjlQ7lPaxItePCd4mQRhN4BzNYPJBQv4FUwAEMjq/CVH36I+i/eXtp1Xkm5IV4/+e0zffWGrvcP
jfAxz+pp7JCtLh3f01gXx3EnGx0HwwDkZ8gZ/dIdF3xSliMvmcQdA/GKLBJLMeIO9lX/0mf0kp+Z
G5E3kWO9nVtkcWYDlBJ0/7/nsH2sb9RBiMeiU4NLLr1bhz6bOyxlgbuf7buz5C5kdUxU2WrqqDuA
MGBg8lKjxxjt2ruvRvjxVFPCWyOfFzuWOWCJLPn6YYJZEyH+YHY7IjChU5bwRRnWdTngNu/rKe0+
MwBZ1TE0/DIXDdEAhfpHuOXGRb4gbPLX76RLcNqr8K1nIAyHuIWyVXyBBByygjd9bWB0yUsOQAnk
OVNQsab+7oOYrwu0S5Q4DXn65tqoZuIbpjeDKinf5sDtTZhd0EPWFVHtZQ00xiqUKIRVOXVzCL14
dkHeaPWC/Uv6eegTvbDT9h67hIYmVERHCwncA9pSKES8Tbrndep6/mGNGUI+DUQa50QuG6+DY3Nq
7qIZYq4sJKj0fBWXcC2Ar94fOTX3vOqsvzw8PEhLdjkk9M3VTGcEBVzMQDS4aa8+GMsfS4kliFVz
iVZIUa0/7hUt4sd9gTvsRzCrz/904Gz+npTz61CqKaGUeRByriLIX8EOUYkEfwx+yyO3UWbn982c
IGrdPh6GuUt+O69YIhp9phUwd9/8JKYU9HjfKcG+/eYfYTIeMGlCecbTcnbnr+7IkSf0wb/rXD66
sRoPBy4eW4v6REe/q7/ylAVzXtBde8OGGs+bqjrwUFLPuC6s4IwUAGBV4V+OLG6Qz17nDmB9rSCY
qYBTd2aBRJ74GqTpPe0ZcNxxZGpbVdkDDHL7XSLtxNGSoji7myd7FOvXiJR69SRqtF9FHtohVzo7
Y0N+9kSpbWr2ufILPZEn0XZK0FqxWF37EaGtYvCYZVxYEvq8+jxuYhpAlx8yjmrgIujIi/EiIiNQ
KgCkN8yzLUYF4PeUqPnW75p9GOaC57Oel4vFUmTVlA7qgNOdYgITVeNMOsgc62349KZltV//rxrs
DE0VFBSQvYIe60bsCM9/u8j1+SUZmQaqguyiUVcXc6PFf5EpMm88ixQCtXn2LUuOYtyzfomzVr6F
JqwtLyfYSW1nESbe2tNbPXU8X33zj4Ao5HzouvAhToaN/tblJODCXI7DMCrNEtS/Jmx/ew3+IZxi
I5Z05UxYIb+Tsewa79CGCgePYmdJv2Pdv1Il1g9i95NHF3ucZn/oi7EDtxaxxEqMZmvBl7BVE1lL
OVkkAVYKbK418cnxzMOQ3tljH+JQYd3mm7oJHG5GQU6y2YTeQ4ps7TBKzYGejK2uqxDqQs2AN2BW
rFIuV2vInK6Ev5mEnLaleBIkCpjm1e0y7t0KqeAO4Ceo5ZUtGMJbrK5MRLARX3pzws5eY9VhIrNr
K2nLjPJRH0rOneTi8JwLRIJwiCamy8ySqNQMAlctoFWAJ+2JxjF8AuGMsHP1ydtP2iaX1OI4JvXe
J2KS8k842yUmZSDi6dr86eRQimSZ57uHvGLdjaMthsxhGFsdOgFMHZ2pBT51cPr9Iy3UPrtAcTBL
vW5vUNNi/LBicMi6OCmIFw7M+DQLhUyjkq1yH+P309lanlJ3jmyTu6mPZJcMPj3lQcxGCBK/M6hN
BqhtU+U8blSbEyS6qY9ax9bZ0+wnfaT21P9b8YZZQ5eFm1qCdcjkM+7iGUxDl0QAi+RqvTHL7K+N
0bWID7sUx2W2wNQ5h0I/Xn9z9vx8fz4d2CkKAL8ydPVzXNmjue7NaYsZICa/KKD2x7H1YeYh7dvc
G3Zg9SjSkaGOt/5bm6bLp8hi45VLjmVlcYqcjmwuwOY3ah64Pd2sR0eU5BcXm88ekvm+yatMRflu
Aa86og2QZ7DZbX0uOB9JQBOiy+udnutf3IT722qTGJaczuniBAcFlCZVqsUpHV9Eyj7DBVg+rjN5
T9L5G9Ooxs8te8Em8l8+0NDkR6S7Yv7fPAfCd00mAfSXE57EqoVyApkpEJrbZOyfuA9iULMeKc0t
Q/XMN1xa367aJ5pcUDBvtHXzeBHeHclzIJKotyUoCFyC1NLqsGtSle9K6tJAcoYNkFMmfsCmvb89
yKrnEvSg/at5esReNqDmOZVpMTouBMBek7n+2ormSnfRPodsBF/ayKHh2L3TzOKklS2MzS5JRnvG
BbJEIClqA2M/B1AcNEolDrdxjszjpG5nbHlk34+mqbZ/+k7LncaIWbaNcETOhJck1R8hGImxFpCp
iF4l/4oLqUzmLvawGdtS1yDBoUyN/rz65L1csmeotWE/n9eIyAchOzyCjhNqXXc4Y/1n/mHgRT1T
ul2JK5OARBqENbwwU0D9BlZUBdND2yZhz2useBSuBkkR2uug8c+dd6IFrgih0p9M8uAqz0iBPJ93
F1H0/kdHyeyk+Q8BsswjbyfjTp2I+mBdaP6EF0rUmDn/k4Ibt6Uhxzl02qu8ibS+fdbnPvZnR+tc
xIhGxZH3N+Gcd+OdfO3MS3EjFytzyYI2Yd3TKYWLIuiFdPj+VVqE1eTNskxYOJh6OhZavbbq49ea
2GQI6OJrhZsJ3qb6g1up3PFJGS5bZv/CjCAdKqWtUM3BUh6s0uu+1AMs9Z5ZbXCI1kWzbJw4bEbh
g9qG3Ue0hI10hbVgbFJBrWi/GM5uMtUIijsWRN8UegmtWFrzCc2F+4mvQ4xtdUndQZ9+Y1UGL3WN
lxWc7MfnB7C74zsXhp0nYCZEYmcUxqoi6qe16rj9mNkk1tU6o5BxIMQ1XJC6CN+W5MUSmauTd801
swikmv5aXFUHzIuHDl5sNnetkGn0EJrboFEohqh8V8/BpZ8+WUfwBCMdK88gBOnVSx4V7dv2fxBJ
koXLBYO1BON+5UOYT03sa8xU5Ur+WH2rmTuWkSyhngZ7IhOhTvOv/ZT3PI1P5rJoka3/VO3JYDDE
VnDj8E1Umc5PHzzgforYFgP15Z+06luCW1/AsN2n4gvP7NmUoDDDTj9yvvLNiPovKhXOV4L7Sw3u
i+mUi42WP/KslTKstJnH/BDOXUljnUfeWF3OJWl9O7cnG/25aOnsv58lr75zL1kX+W/QxnB6D+SZ
IKJEcdm45qETPZkFHEIBK5Q3cxYmBw/UA4OZkPDecH0cGTapJZTXovFIG/B3ka3ya4C3othDNyeT
H/p/lhi5Y11rGHBdkc8E5Ar39KYfPOBBDRo8A/vWCcQ5NiNl6zvPUaDcrxeYpeCT4iRyoIIMBccw
rDedP/pv7jGNSsUmDwlwz3RJoq0Td/Ati4n37UpQMcm/CbutJ+wSRLgLoi6mJM/2UZGhFhKdTWWh
S+DetCPqs063ryxFgtyAuFvDMykJbbf/56gQ2L+Cd08Wv3xstVcUyr/J3edmoSETOKlajcfPuJ39
0QzY87/3JbfC9csvZNmzQdcvIUN0YPjATMHLIJpWRA3c8Ns+zFhjQYWcZYexQh4nNBOaMMWJLwXX
NwlbtzlCosLYITEpGgVEsBPvsumOcu2YX1SM56h2Q+cuQzKNqrdccyQd3eudESyL4XtYjcAAx3ya
izK/IShMQReoUy+PgIgNofE/oir4cDZ2h3BQrKcyb1+IVmQzOgIgjLFwse35vUfIp0p3cQIp4rry
sPRVwdeLKf/Y6w68pefrw8bz8BMF+9EEtqW8PzcJu5qV+ro2hz/CAAUnApZyup/MVPQI8QZ4yHmA
ftoozTYl+Aur/cCK3XDCPa7h9SPo5cbOfBo9gh8OBGa7BGANoQtOdUibofH1N8UJ9PeWR/n81BjU
wZyyltoMmIOdtq/j4If5+vRAioYWF8n/qehWUjAvxdCIR8tLRl/38DwbMA+VPzOq8NdMdwyrNk3X
M9FU7OlkrXC8ZZ6D2tRp+sE8aGb2Xp2HShLIseROKaBJkIZ3lx4tsbHJZ6UBe4LfLoZACWn0p7oM
ZVxyqIFP+Kyso0u4yr8/RS3EWFYRl/1OL0PO3ov9SS86awhUJtP57nDtVSGJyGHOKVO3YIaecvEK
03KgDnQ9HQt2lJdz8yaF5W4jEZ0+7Aq1VLSy4kEbz6kEevImV5c+8DmJsI6irSf9/gxBfzCUAyn8
QJyPqvD0CvuLI4bmVl4jGS7Pjg43hfi9SqXyPWgyvyfRFNt11u2Ptq8iZSrIPzcBgpJ+l5cBmIga
i4CZIdRJVPC2kbNSYrCwJBLPmLxS6W8Fkc9wWHXTMfLsLbIHMuWss+QyIgnQh+DcqP6PK3nA42rM
WDzaAbSOFuL65X9i6B3mBxvWqKOExRsa4S4JPv8jpDy33/8cgrwYQn8/frR76AJnVahP7jwobuyM
PrpE8xTOdYrR6h037ockUSyniyAXElFIDjNRhqfx2o5wxdwatbLIF9OVc+32dyGHP2zyAKNP46rz
xfk8HVQ8AeMhdTkcm5shrQ+Vvo+yXnd7DXkCPeR5fbY5xxq1IKfmyfSWsrI0g+xwnuphWhjgRGJe
5JPSc+/c/SEEvfQJ/uqODytbzxE+dqmN9H9eEyh8A6s022sfX/KjDXs11XxsNPWI+NMHO8RcfZA9
iZ3F1fiRH/VWs9xie2DyAZ/ROaugiXkhskna1MyN5jvbHdwvhed0Q9VTdtZZ5m5MlKFS+IcR46ca
7LcfRc+trn4BqCLthoW4N1YzanHc2vPs8CEmCcbgsYWqoBws7F5o+Fi1jOCDXa6rzpWGmgVXKgsX
m4x2Gux3cE6sR6BXgI0CDNUoRUJAeZdPgRxsG5dwSw+Eru6q1n+IYs8RRNIrpsw8gZHctZh//1Dl
Ncptq+9s/9v9Degl0ovReyr6/rdI3vPRg2tSJ1/ySZ94qS9b5OQfFD1RXIM+mvQATykZAje17VBa
Gm/3A8QK/gxky079T7w76+K5oHjuHHPhNmvnwm23hMagafyvs25OXmRw0qmetsBcQkQj+zk7Oiz+
CN9NQ6CMr7XlE8b0v4vnFlEMHqpcGuRen395/tzuAz+DsZJMaMn8AaN7Vkbavmor2+eT1kt2fTjm
Hac5LofNSevzlhQjgMBmKVWNYjBMCWkPz6pwvTr+m35T7UoLizRSSvmk5BEnyd3PR8Ikq11Loxj3
7irtw951dozWGY6J4d0g2uuDa0WK6O4fF3laKdoFq3InOPC8enF7EDM8mYo6AOWb3rQ94B4KQ7Cn
F9SiTSahM9Dunja0hp5JFD7t+ylRNl6RiNGeNLWbnq310QcO7LvarA2DgkSYHvq6Y9MVLeT/WBWX
/w1oYRdFVdGbYH3M33heKOpMRr/05BrR2/kQd98ATgYpXE8bIb6IWZyEX50TSgeurHT9ZFvM48Ux
r9g4HZ95PGIevVvaM/9Lr7yboZCOueBkQY28koS8bRGAIkDhzwecpeh/xmisa/CSKsmyOsGyW7xc
kH7OrtmgQPGDsorC+kwm1kDXLOefjXSAZ5EGO9QpL5pqL2ZGNr9qHe01XfMowpQZBz31pTeiMiYU
zSfZXNqZQkIiWoml1sBY9in+gbjHDNQcLwV1v1d7Cvl9/Lg9+lKbH7O2uJMawgviDjddq0sUi/hw
UwwnoPL/DIgbhqJEBI39S+Gg84RpBftkK1DRxkBgTVAgM0hO+QsCmu1DP/io4egNos5Sc7ygA6/n
ajlTiP0UDGbrwT9+c7FHK1qZBSnmPupOZXL/nj2QAZ+VA/mPut/qfl/VTI1B7muckFKqKOpYgA6p
ZJGtiMSUsmKlaStWzwbVoP2PLRQ1tHiVpNyJ8WMjTawm8paWU/HMfBtFE7ow84ng4IKF5+SVAowf
ezMHjFVd+6LxcluXDLqqDR9owHml2oKlavo7y2+e7ebCuv5LDJ2BJwq8P1TTl1zyj+PZM6GGtWr4
UvLTE3O6A/h/02fzXJ54yCX7wEE6gk16s/VDfozepaGarWCVF7/tRo34cetf+6ECgOPdWMe9YgTL
+cGEHuLrFAzckBnp0Z2L15YQRX6q0mmS4MdWhFhTKs6ZVPMrXYiQ9pzxxn3uPOFqHzletpqexrka
7YRPjAQlWX6AO9F0YIHtF6dTQ5y15qyejm90F2FwRDfUfmbfylLwgqQz+d5gLfCBPMIJEVQ89S5H
G30dxpj4iUOKracJlxKApLWjv+Tg94sxKBWxmiJdvSbhZ/SmvCwIH+8rR5ewIuILxT5mNtEL6x1q
cD88bLOifC/ZJYSrH8LK1sQmORCI6KXEVH02J0rKPyEGMNk9CkSq8XoYeAAaDnmypEuvf/5VKWwT
V7SG+F4qXJxlb7Memb/NC7DFQ9cSPgD1cJOIug62e+D/QEiFOhkFyfb5ZeXaIn3m/cFc82ICIXnA
A8X5bBYwjKW9Zepgw4nxkc9ZhTQUu1M2Eu85kMMQiBzpU9aiH4VW6zKjpDhtceLmQm9+sAJ0g7Aq
OuiI7D2UBIRU1zB6s6iAVByfW4KCXrDQgdUTGyKNA0o4SXVXvxGJcnANLJaTrybFEXh1mL94BTWj
Ux56KEI69z7E7l6AvbsZ0eps1jGC9Oger0CmyZzw2qMINE45Wpd6Zvh9xWJjBFvMLodVbSts10Si
jt06+oespExN5kEV5NIUrhlaBLtH8zHstWy3KHdcIiduQHcOMFkI3W7YtOSSyv09IlhtDEY7pzSI
nWB/242icuHnJiC+FikRr2ymaPa8f2Uhyue+QNgBGq9n2Ialc1ZEGwY1ZDIdORrjC80dWyzPR1aY
vfbUY0Q1WcDl1PBZWxNcJOIHIPKGB/fXIMGZTBS/prQ0Tsz2vJLDNEVr2zNQBLhseFH/pOh6/Mtj
nwfKrRWPpT3Oshn3bMS64xR+1nm5vPh32YJ+6fhDQyZtav7tBXvQ2daGeVB62aH9JjvXD8GLLtbf
b31lXaa6lgM058bwiw7FASzLrVSL/yBEH7ajQFeeAOYpp6wV2btaYG56kY6mioTRAwPqeMgehRZR
0w61N+Gri4tBfaGTGUVs3DM53TUfuom+SWKC4Xe0ZlcEfmxg3Evmf4U+bCOx9FH98VTH1S1s60En
irVsPeMPrD/YBR3Wbk9YMR1apfLttyVbTR275Wpe2sV4P9MPXS0435yoDvbAwFPtOYFwy/c2obhQ
y1cp0g6ps1vcFbctHYE38xiu7FCy1YeixSkfTZee5S6m7X0UEOUSbkTXdAMdsG3GIfx1wyqT+aLY
JvFgcp4K33pegAev96eTXLdFT1nfTkK5iVxQbTDgrMzi0ZJMF1bLB4+w1vATTGx1Yj4Zj7F9Df3Z
q24gch4iVX5NTfAK88P92zL3naxM9liai8kOEEkVpJ2AK2vYWNwtzXGZIuPX36rw05nLYtOoxvX1
vktgkzBmrkprH6m8+IeXb3Yo1UWKALfB4BJls7FY//GhwP39Megwuayjupju04Btwl/rTvHTJiKc
EZfU9f02wqmkLBPd7wcOBcy3eqBVn2U/0feAgkji2WjhZwCpc3xLojhAHwiVCXDYy8vSBHlq/CPh
MCLoJ1lKBCAjmvlq6J7HOJ5DsBQG+UyqJrS218HP3wG73S4efdgtXPqqkXoWKG3ff0RYcc/Dqr50
KuJvoAYFJqwWbDh3+EM3RpkNK+wofjqd7m4TAUAifGnQ/mZP0IABFOAHJQnR4JEhGPSvf0D/9MZ5
OkrGanSx4V7GIEBvexehUij4ZnR0kLaidLRbsp08+AidSZyeIB+xBmnsVf2ubgqurtLSy5WinOIL
JcohK71XzmqEMKA6C/xcIbCmPqeDrvmjo3fmVS4ma/Q8Op8a1OS9++pAsjOdBvNOLmbukTpIdcKQ
6+2CpBox19pOr/J2q8H9XBna1FgUHyn/DBiQeuPK1ruRB8671pTGhXafK3nUKXRInZXBAQykOyUP
1VWd0RUUjJbCuFu3mGWHRyBY7k2WJXN9tvKGqlGrJqk1UJjPaQ9hGrYlz6Mle7agBJKg3eRsHDTX
lHZQ6pZ4uMQAhcvpjWTYVOJYkmPc47bGGrfLxPHE8oQcpmoAKemi9FFrT/fkfcnTxDmLr8aGgoKU
45VM9vm/f805ySNljnpMc7IyhrfGFM/5aY+amQhK1XxsV+uzUCzzVAgTqLXW/CJLg0qaA/Vv7XUK
ipbscvlCAeB4Y9cLT7Hu2O8lfa8qChtwydkxpHZtYH5YWkgsdxbZEMyFHXjaR/3yMUr93a8mxgja
rH9UjRybr9kAFmrn9x8OYAYIX/xRWTAXndhm3Ok7u1ibECRukrdgioeUpGph5dHPSfXlZ0XPJDxy
Z0V+vmWj8OKeZ7SsXR2cUIeDviR4iHP8bMd0r5lb9S65gkzFYCAi3/UdjEi9ViA0lOF3aphJVlJC
0JgziKKs2qs4Y1vzMLw/xV0yeujdBJ0oeMNe0aXC76ydk0iL8rwA8+JvNG+kVdoZBzw6eQXBcV3X
s9OnvjJtUbXhbkJ8MAcsAqpUOESfhCEDzjNEdpJ5lAOlT53GtEKeafH6QflK4+nDl56EnXzJnqa9
PfJpOJwiTZkk+l1CPmUmKex5umfgmgxrXyaKSOrh0Cr2ZoDDGBF0usBcC/Y7zs2QpyBi6PQVXyOY
xvs2Ept3J67RyXGkKPNUUIg9X3nGorfFdAOLqWgVO0vq7OkRK4CsBl9B/r2ZuTtygJbnYzIxKNaM
qTn4E2wNibGFnZWt2a6+VQVXCGVTFybZMPjEBczJTg/4C6HDgMeGF4LGIsD8dtLnnET8MUvlJ3tw
LhBXEAJ3ulnmZ5xdJcFXB+00kWifTIo3JN5kCx+yBRqMuoqs3lk2vWHc8LlSNv423ocSJv61oFzB
haB/SqQBz37AdaYr2U8v1N2N7WVpisTVlqtpKP7e4qg78oowU3d15KObqQwwN5FBaf+7dV0L+TAA
wG9JaZhObcP1r7MfX+A8n6eQtTl6gjdA5zcW2FYEqyi2O8Onu3IFMLtjlKvY39m35w7x7yCaNFu6
EYUxV2mdvo6t8XKVhPstjpqKVIJHx+6dty12Yyz1DtGojV5Gb+m9Vg7T+vFwg6Gxx2i4GxwW6YXu
7hva/D3BYev3JsL0W1JcYIDwqXqVFJ/0NepWgrI8MGalQES54XnK/ShZ8eqpARLRuKiaL8/EdyeE
H3l3GW9Vob4uLwxOTAWZ+WX7luKNVe0JCNBSVuHU0dNs9m/SyPVX9Dcfg3Yk3TlIOLNw0/h/IgK/
2Ytz6TRGzeBjgXEudYAHl9aNda1wQ/7XeOYTmSIYlzC/ry3WSmLJ4Fm3pchWN6spK+1aaS2HSRXw
eXN4ud7xco1HY5sETC60jkojYu0ZjPG4PfKnSb5yUY94/jPcdqVHNvmKBT7d+owXLgj49XDrya/F
Xusi5tWmASTIk4ZsmsSAuqNcvxw8HWpCLELOF459HxNzZnPQ/p3SXh9vqcroCCcHYJUxNKZzu3LM
mdioPUw2Wd7C7uShzLG48aA+a9KbxLbNNB9w4ENqjonKP5nm9MOtoDYBC3lWfFFY4k0mmFoQfZcG
q8oK/1g4wEjVpVvYSRftON82x8IYdPe7PJCFqavqI+ndIuC0lGRQR95OU8se01vo+krZbThzy2EM
IxZA518HXdbLdRdnIp0rkH3ldRVIbkv1VmqNfLBqp+NFJlciQ/2wnVOcAxVXN91A/HGpVz/NmpLC
+8XeTnxfwZxUPVwc57IgsxHbmcJt/j2o7wYSnZY3lhGdx9/vcUCM8Vfb68nuyl6KpDWMug3N7Aap
MVshWTM5Jf2h+oxYK9q6K1ADAolaPwm1UF7nnfHtIfp34EIOO36I8sBl6vFMNwf8Le7agGB+UDlo
6UcS4+ZZ3JtD7KHwls5An9q+QZFrE1qikqvH3cVPqtTMB5i4TclVWl/igt9dibRr4MJeMlnPJePu
pCMggNzEVfgJqu0oDL2YxoELZxR5/zxc22e73rXOESn+RFjMttJPlgHpl9Es+PwGh3eqDqbobTIQ
YORME3bLtyNQ0/3TpstXc5Uzq5O/h6cVMRn4UwZJXEtvUN+l6giXwGrKiJQKMLdQIv6XBKmxOi4v
rz2DiEfoYm5keTIeeWTXqIZx+d29NnecCSd10U0BZwSshIWmjc/pzuP/IeVv7wqtqWp8WZUXgRDs
cm8/0ZAEL1Pta7JyHqaND8B4ESr/zwob2rFEUfeOr8ML1umKChdr7pscE+N13aA0xo2G+RugkKBg
dRiVtGcB8RPZXda86O8R+yogrfg3JExMNIMsBfKY33zsEnih7v1dxNz50GwrjGWZhCi9aJ3Pa4iC
sDMBfRL0hK09XFijwNpIIXY6gAMY2Xi2UCNAQWDPJYO+EceaZdsogMcdoSCMRFljG+cNsMbABfhm
DSAQjl2qzqSCngINpslX0oyIaFCKbpOACOsMsbj9Hy0T1SNzS0zaQBRA1ekfs599l+535EsrTl7w
XusRsvhWAJBl8XAfboCeZ5DPIKmv/dfgtmJWB+p/BNZtNG/froR/1PM8cICkm8KcRRsrd9F14goG
Krq8++x00Yin5bWRoFuqC3RXYOkh66U6njTl5y2jM//sj0n+nv9N6sQtvIhBmV3f4b2joiJdygzP
jVA5XOKxtAo5jWox6YE1B/grgoiBg0s3LWG0k7uUj5j21IMCxV8qd8oxlF+85eFnW1rluC5yXy+m
p6OFDmA/WEbP6/3pTDBp/x+Sk222euy+ind/fBU9p2Fc1lbfN3Jygpc78CT1wPKM+youML0at+P3
1wtOBFe+BH0vL8V2L8tisNCmwRnbQ8L7qVtt0a6f2ij3oe77bigjAPz/j755lpt9TKwGobVIZygE
m/IoWZOwoGGy82CUN1n0NzuJooXBfRSZw858sZGoLbh0tmC0hobXomO+M+6qsMyqp19Z/xRlZWHC
et0yAU2njgTyXFuL/zSnyq1NXsZ1S3qdrPK+xZTiXrFQ8Ka9aQHLr5+yre3whGZoPvVDPXXXuZsX
Hf0EkXIX6NtGcxQooOdBqel27wyw2Aer/wnwl/5Bz1VmjCXsPN8uEDJCoKFA46J54zryneZhS4+1
Pz+AQ6vW6kpGG88g+epwJKWv8q4xEzn2nXKTOBhfZdXWifnIm2MVPL+u7aNKdtn9Ka5Jzz4N+cpe
dPIbpsdMLkpQdregwRF3baXlv0kobPYMK6CyoGCrpDGVb5tlGIZFGzkyfzpBf5IYjaSE+WMBDiJM
zHLkQ2aE13BuGkGattzVin0ucBFfpWhYwZSHJbscGNwReF5N1opjfplp2Ng2GdBMv4iz4EMjTY32
9Nbd6EPlkZpWVsR9aaOQqtGbVb9Xafa89e2l1sMp8m+uXcNnRb7FON3UPryl39uUGTsDFlqq5zv7
LYzT6icZsOGOqBKrRzxnJBS6IrbUfQzVvXAZM1me3MB6aBfc9P+JZgTe+WcJuHNp3vjUIKmNuVjJ
EVTnMny/xpD83Nwz2eLU27YsSdwUx0pjBxDzFCknvby+9noyHm4CBuoSjG5+anNWaAbcxHSY7Wf6
L+bL6OR1lX8Y+EqOfWsjljbPYGs/iQCcJAnZll0vMcjan2/Uzig3zvgrA4S4tKwnHF3QgVzLBPxe
Ta2qAxM2HjNHERnPevqgRxgt2UcWUZdgY/sEd7AtlOM5VCe/alKL7ferAWkRZiDXlLzgq3Fj2NMb
nmntunFQtc21VlZAiwZoojtpMfJSRnu+O1x7o/pM7JILgo5Sbj/8cbHvleArZpv4ypbUp85DPj9N
abFrvc2I5sz8JmOtOvVOEbkPbobtsP6M5n2C2wCy7E+zXS+xdNMI0uumCWtf6J1w5U5KlolNwX6N
f2cxIr4utTN3MnG3TaehIgFaPAm0yKZ92X4ok7DDOXql5/2v3u1Gls+hCBMPARv6wU7QMVg4j1jY
1heQdv47cPJYy1lyypNDUF/9vykb25cH1o04Bz4G2RheG2hr7d86yjdiR723B1R67NWhfEEkIH28
Bf6vldyFVLEfaRgH1dEzj50yKk+T932LUWVv83DWMtkaB6gFQ6G1MB4DXVeh3QAa+CsnbSATSbAQ
UYqGsE4i/1pWk5lgrXeukeygTruBLmfEBGTc5DKE2JR2b7dJNq3c8N870O8RpscNlZZwoWk2Nn0z
chnWRf8ravCkD8IcJ2cmTqadVZK2otTBVIw7LQunELyI/Oq/dLB+3/yP33CkLQ/6dPFq6rGMKWyR
JyaFq39FAKvWpPJDqzUxXVrguo0mVMKgs6wVeYJ2yuXOD9KEkPthS00Q3KcDIYeAXTJyfkb4xH1o
1qGctxCmlL6nFgL4HCysERnQOCBUQpza8WeuPv/cF6VeENs5fBJ4mdipHzbk1muUc6h699RkyegN
ENgOnLadG8Tb8PWahLaBers0NCPZHcfT+ZV6q9thQSo+3DReg4j/+EBHlEw2tmTsxDSA2XXqxYki
jFo2IQOfksPLf84VFg9CNYdtTRovkghGdmTZ+NdBJfgiZq+2x8IXozuLUQVj1wU7Gp9BpZopeT6y
RnHYf+VDgf2wdnNKLG6lstJzlPTlZ2pq3rPAR0ttAep9+gOnbx/lCEe/vJvTbKR678hMZ515G0IV
FKT4o+qZjktHVcHyyqtvNgysqPZRxS/LMAMgR1j5Gz93M03Q0x0MN6OmvCr4Khmc6Cu91IjLGX25
i7QF4gzW6Qs/4gwLoUUjx5r4KnzTxV/F2Jt+IlwEOXE0uzxJwOHQns25zPLlu+Bj8y9geLmizcmS
EdDc6DguHT4eRqTWOvcP2cm1tXfiuCCd0/S9mRO/UMors0KkLt4nplbt2qxuoDd10Hn/GF/vHnA3
QguPYBEXVRSSaKk4wRTR5gJrUgbbt+VQnAk9td2381CUOUO7BPZmrJgTKT5PAdEkczZZBljckL1I
9McB68qDzjM5mZXPTmbX/FW6jj7KPLiWhkvdbpz31lNc3TqdRzTq1+nCLcxRIbfkmf//ejYpf7Tj
viLn3dmydK9nKAXM5fUC+pH36kPnTeoc6dpTrUR9rvnXR1PYu02O1w2gOWWzRUGk+s3NOuQ4wPNW
QPRAG1jvROClASH9hOLquoiLrPSwfDmSxl3hbR80hm5f8NfhhhaH+aoP43MfC1jHlquN2FbMOR96
/BctPKkp6nzkf+zQkeuN34o3YgtYEdkANM5ptUTcuRFxf5caZlFAVW1XT71LtBh41kXGC4WqMDR8
hbuRU7XlCDgZUiJezi9xGYuMV4KKY6TUWBxKLYnw2yx62i0pTCmiLEoI3ER2Anu/fdkhUQWwJn56
kRNhOLzuGTd5Qcuw1Akj57TqMbn4aQ2A10TwTYVy6ujxZGGR7V5oaw1t6Tj4pP4ghSROI5wR+VkT
0+k9MvW2puWRMF1FA5l4zd/WhqRbGIxzy600cM3EXWds6Hg9cV5Tg8/PEQhmWjeToaUOBukqrIwh
i0roQPJDN50daAMjhN1ADoFmnEqNpsCZ9fo6usp+CtKKcdME7ATKhKhaG2Z3Ik1FY3Q2xJdDpeID
acVwO9wTqKA9qCperqXBVHQ9D5H4CdLh9sI8lWQIEiy7N4Lc8AyV46/1IG3cQQGaTcBN4pYUsavM
sZil3avNhIdabeavPJWMvWlspdLA9qwHOJuoYWWks3nAqYqwcGLYk6vioxby1IUTc109KqMo+GQJ
K0VOAjGzvwDFPZlF3HGVzGNaFzS36G2PnqYH0sK6zczZWazmyu0mlw1mY6alp8wG2jIYQiy7xcyo
RKfyyhIv6cvzDNkC8HBkqRpY6RqveYx/OyBT03yWB5LLzEChcOupdQUvf88gT4P6gMPOmoXmsXP2
GNAXr+nROYNYkGdP4iW4oJgCq0KjrgkwyOogTQctqOXi0U2XnzG8pMgjNhdS7ciW2AVCsvSRAHVA
FQruWq4dC8phjLS5i/gvPMQfxz9PWJnD3fZV8CqNhnhaCpHKYZVGg5jH0CUqMeIM9v6F7FuTEafT
8M4qsqLItee2Oj6dCY+dD+KsfHwtswajZifVPPQBQ2mOnWocgxbsugL227OBSC5507tZPisNJaqY
rf3bl9bimGaHgUFoH7NPsUFHITqO5s6CNV9KdgFSeIpmfJtMGNOh9dJlEfR0ToQQ0Gvv5jZc+0r1
RPG7N6H52TfJ7OVS6AXGg2qq1RS9okohVc6DVi5sse0apZ3cidep23jmaQUJtJTpM1pEld6WygBP
PJ55kRm9SObFmbxOzmBjmb4OHE0ejzKkaUngF0bd8FISFZ+DxDipY3Fy1xdM5w246dEEl+EUvEKH
JKtt/gNuYjycgKA74J0CpnKkGfuE21UJ50D7WLYcsUMMejugqQFyKjeJoINO5MTMv4Xgb7s52uyq
tFHnmH6WJhn20gryQ9eiFERRyoSM1oBsC7ens6LwYOkSKV3GfY/Z1iU6eWlHR8tCBZ7/EmMQ5rCU
R3QSgG4CfwCbbWmKwSb1SDxdj/5nXqtiBDop9bgVluJLN5iBQl2hDDKd8ocyzZXl8cQFu/ydEABA
VVWgt5GpkClnqsiITO5IOMByKomVRuENMK7kMH6Aaz4ZslTWuWlIDXifJYrcEB/sMt7tlh8ejlzh
4IeVveNDKG0xoFHfr7Sqhn6qay1FMhCVBbSukt74WhfmqMD1zBPpN2t3Dg3EliCPkXEosFdl8b+h
f0njPsa4ME94fiFnUmRfmQQOmhN6hVPINpmqjywG+7NKveXZqM3acDcNL68VvCc+li+NfhKJRmvC
dOv75gVXrOygBGil8dybEBBxRlEvSxOsogsZ3uh1d1ZWf+XBpjk9DtXfJfAJqktRF8DVO5nkl6D7
6JcOZDYhf2kAzHPYf76u4LTsaKPjagauRYyAQuCkb6zTms4VrsFL3PSHcWzwY9k+biHbahK+tA03
QQV+CRbZLSYKxIBNyvNi/1liuVT9yWFCFkzRpvx/i0EgUS3i73dbv+orjbwDZoaeRgY/th7YckFd
V1q4fa3cLaejHeAybCvtQfAyb0DjFRUmEGFBbf2rdyCw+a5LIJk3b+chGYdl89f3hiG6hS/vAIyr
jEACcMN83sNuO93biKjbsN2lhZXc0SoPT5eep7Gn+t8nBuCPH4H4/OuprQTPwNliv44hDr6QOlLF
rMh7IxaS2NBOOm2bxtDw37FThmgCgenWohVUXGX8RSITuinmCR8b4CmNrZk/3jkOmFNMP4kfVuqM
AplyiFKGpImXLlzd70THm5igy4Acz2hub7cU2N1qgA+OVzHjqKq/4dN35EcyAoFuV2sZ9gib0NhV
VKxCUVvuDrwxU2Yphp3tM3M3fKTYv/TeXGQNnYssIXlpTtkwhdwq6yR4sjVKbKgypo+vQ2jlIWo5
R7czWSxxHDOx6t46stthvrIkSTZeYiLfvEnDnJJ3cVb3baqJZB6UVLXgXBoi9K55HGp0aqLx/Ufb
0DxuGCC6VRRjsis5+UTplorw2kbAHBzxvELXfFtTEnhQwTuYeEAqnO2KWK432hj5+VrE0NyA8bfv
ZZBTUDjlz8UpfiegzmniQxEuxFTtBGkQ3E7Gg4/jNtXsmITRT5NZbWwGvsQCP2EnnwkZy0B/H8pd
797APDmLJ1XtGUibdUQhGiAr3VIEv3K6Wc00ieRX0Hl8VIiz9i5Sv8Rrpvy0B55ec5cgc65bY1bn
KLpf7MiH5fRyiwObJ2lZPgZBkhmwa2g20tqmYBHl72/7V1t6gfCSk/jPjR/6ncsVuOU9zC2HNv6E
qBLQDnOLGAAbBu6fzwcHc3coYLNmDTbWsI1DjJJNbDQFKOw8Q9RtSxDGWkjdQ7I9tWKcnOSewBhd
WQYfshj0pErq/dmam20AzuiTeN+TgmSwC2aGeZI+/U/PYsWBLX/Rft73q9rKFjBX71T0cCIBT+S3
Yb33IlLOXWluyeuC9hq0e9a1GJoyY0pB2GyJXYt1cDbrmB1kXv9peFOCII2YdmLlYwd14d/w/Nut
6o+/b+TmflNTCL1eSimjOGp0w2W+Qnw01Q1lxg9DUxK0CQ+UhI+9vgmkMkXP+foGyEeQ/rCQqV73
M150j3qVj0VUZ0I3EP2BQT263gA2bSBgIaQjI1dDAhnbr4A4yLFCT1GZZti0dbZtd/ovzYxekWpv
3KE+jF3rB1S9BXErl4srgoeTP6Xvh18+gDFnzbpUv1VtpuCuTedKW4yHdQbEuoxeGThlhDh4eyUW
pfkrjR91ALhgm1p8IDmrp4AFXRcp4AWe2DjdqE4M/aV8mHZZotyq4Nsdb9UTTto98/tE3gWmrTI5
NqGiUbudTDeq7aCoF2IgthYglRluMAcNX0S7gpYSj3ZNDG1bhVJWeZGgjofOcA7mJQDV10+GqzeR
8WKWxi714+PKW0VAS5uUTLgKpxitFjB4I8C92SydQopGN6kycd9f1KNHOUrN5wU87LwBmkgvmu1h
TZW78ady73SNXdLNNUA6lspPdCTC83TDFPJuT5iJWWnL/iRmiT+p+D/glQTSqy1h32OLp2mA4wOa
JXwH6DZnrj0AhFi4+b+K/s7WKIEfR0EM4zM+5Mymn9pEreSWnMzYHc6KlVQ3xYNj8ouWDpdK5Zdd
pMRB2ozrQsxthtyubNFUOQu9R0UMDs2jysOTMMt6IZ18GA3i6vSpJw+diDTq8EDGMayuqf0AMfnI
+LVyJiC/8QhIOvbpx5QkUojFGsYzghw18UfEfe3dsswi54FLpKy7/PjnHF+rmLYyLz16S6DDK+0R
0/ARSngcXNU8pM0lDUnxzHM5T0ghxyP4/mSE5Vog1TsxYjRmy+o/0MfNsLT46BGHaZgDb0OeYBzy
07lnDlde0+wbdTiTUhuVzOTsqMLVOJNEmFEH0OjfhJ+3rHq7ymlBTyNRUotsFMZ4/6jURHjbOoDv
JNgXEqgTbx3r6lKEPOCKcnOLpi2z58ODgsYFs+PL+c5y/gl9ZXaTExMeVqs7XD8rcpTFOmCnCqqP
uUrrfuHcuEuJmRfFzhsdx/Fbct1Rv4cITdlhhljgzXo8CTRLGlcCmLvrYq1P/AoVB6FLSCEG5iXK
NDHlCkeP99pZuLv2pgiCefEcwDwkOr6IrYyQpfl7AptcDBnAvsGPN5iZj1OSc3xMcR1S9bBYgQGY
PU6qS3oUbjdXh9xggkwgQVLBZs4D6+T8gpzPKGTx8v1p7sDhrbl4AUJrlz/oV3JdkZ2r/szF5Xzw
97YYwgPmLFP+Mxkf6+6p/hh21RTLOX7td01ZE5UX2b5ZR1zpWzNe4KzBcSqL6bOppr5k+EJrULtB
oXKZnirX1xFpCwvcFbOq6qZj3j9m3f1IpJHAqfYSuON8Q36RlV3P0CGX/MML0y2i0Fvm3Nqjt8+Y
F7qtN21T3T3TyOUyZHsZMG0gHN6YEYunNsmrV4rhTWoyBcvpOCvQ6dS2csLVGJ3sRgWp+U3i4Pa5
46EPS7JQyc3u+UXq3P5lFcCBY6bsGUyo13r3ROdfvrVFY96DPQGut4Yzn7cpA1nSyKNP25dL1HxP
Og4JWZm0QL/EERpaK7UQ/yOtihwomOkDPxlaLEiUEYRpimlhFJQ7y1BYb6k9dE0a6eIEbNjX6gd2
xD9ujX40pXCqOC7EBi2g8jHkqnowaYmEB2fsI4y/m3NaJLJ8yIGJ0fM6NCGIef9YIIR2wN9xiLqN
ySxIsGBhnUAOQhmyfdIR4776Xj+tYxqthw4aQxZVsOcy2wWjpDnj6OVJT6dIYaSyaAl+MS1yUJ//
UcS8b5fbo0vg13/7nsFXuNnsuD1egNjBTO+YNJk+wW2RNG2aoRwQ2mwbx8FUZumpC982RaqPyWse
cg8dKo9bE10gaQ1bO0AUTnILg2oZgnOWywn8gcpnLqzICtv1hO7ZIHlHJqIraUNzCBR9XYqdpHId
BAw5R8GYRzJGz5jTa0XgjFEePLaPzLLsJsrNJOYI8t4zZKRksR4/Zuddd3+DX+0NSDl5QaBDxzfN
JU+vXQmjAp9iXyedauQ6UOGyMlh/54zYBoMSnsdSXG0p4hJmflraX/RGHuBOEPvvpN1zx1jnKzbx
cpqN3EmJky1nHxoMGhu/TQLCZnqwxRKzlUbGmfFT9gZAfcnS57D1ayu4Mc3WSuiO7l9teBpWWchE
IbKWm/ICA6HcohItVY9G/zeJzsAQnDdZLpKSv5NNN24VSWYaL4TuThUg138AkXU2kF+5GTmIdNJ0
ccyQn3gF/mHbiwlM7TPbD7DctHsbtvwIvyFnq2nR1jVa0X5pJcPnhTEmGhdQM8oO/5O80D6++ZDg
2tINE6czwjsnOwVTlFm5CD5DJ1NQ8ouZOv1gPYLY5eaKWNxvayg6rYtZfpuGrTi+brNhrkieWTL9
fFfRIlAheevru5je8RDTFM+QTMGsf9O3JGwoY9TBPqdeIOu28QSi5ILJ80GhBjR6vmLrSfpefmdM
PNEL5hzfp79K6MeLjYDBq5xqwhuj3GAp3uECG0PRiqzLkeJbtYNJFnRjgoWcCyjznp0MEkzjSSDD
2egDr32pRgA/qdIHowKhPtfbqILUEURh4VmtuB098P/HsscDX6yXRg+GafxhnZRlWVfRutZwMOY9
A4Xk2GLBXkbuBFTG6V8xmDV11HkQbaQfo1JlnzTjLEm0Kiyem9bKbCFL3NsDBoDSKZEqoGbObB4+
zsy6Pyta4BckVItiIGIaW5nYDR0zYuBYQ+9aWOby1LK0i2K1EO0jOu6wQpTAG4g7jlDChqNUzRcS
fH+/9zfuT9/LedyFHhOnm9FPtCwc5Grxk2YqcsvJ4+FvdoNJn5wmRU+rSavxRaC/q92WYdPKt25A
FzEbKMnt6lPxVUyYyOLRFEqpkYK/W0QkrbzWcfN4gWpRnjrjMAdps4hjs6q+SFRnPnVDZYoa5vng
z/IYlnq7xNsoYyxRs7ah2lwEOC6fQTg5EUB9LNSQ7M0HHYnL82Ry9WwjzVg2ElXUGw0AAC54D8Bd
0q+R6D5Snned0xrDuoUY6kNkP7Kxbtm+eBBwIAjDkWGb5f03mdj9Z+NeSkoWwdWhlE0QNJjAsV9t
OQv8hNWHB+mEGoEsZLufIrZs7xdfcpiyp/sUoTp1DoXH6fZsz9ddBxPWiy3qTPz5hG6fzLVaDtvs
XC0YVMEPbZjepDlEfmsECdAVQs4xMYuchRchPj/awkLq0fVNH/1jyG1qvFqacHxxud3MPdSCL1Uo
B9OBZPYf8huELLghDvnQSsQq+7LYIa1ZM/sQjic8BjULqf4ebRU/ZBCbcQirkId/gNgfmsvYFot4
oMx6xpkoY5wlrpRaNoL1uMVHWHSUHyR5u3sjQWIbCoGsmGo/Ju3OoI4IpEwscD+UTKeXMuqt6eOG
y8NVS1DqzZeiDPiGPRZ+XPVHUriJAqbYXb88X7D7I+ixCgzsn9tkpPQRjvGxUKtTQhnnggoJcF6/
WLwLzFXkd8piLzVTy6fllAUWSxaLaqQNGK34AzTEmUW9C1OJB22gdJ9AVI3oOjw6JSFBStOSaPlI
esvq5A8HylQ2cG3RsRN/4oeDK5SE2sHGlGugvh2f/OQlAz8XXQioxc+p0h7rhFzXfM//VXBHIJ7j
AyN2ISx1uoMDKc7sGO51hmQoD6KBDBQK4KmlGTf6fH5ojHqiHzTa6LT/4Le0E/2zVzataiKF13ag
NPKrDfAiz7gpNNTYSGK7MX2ojm2eJTBTyf2KMny+RZVb6zWafYmbakLcEMpQp9pvFrKfU76c+p1U
2vPkVNK7EnsnltUkmAHJJ36DiwURVDzZnimimRRdFX4lR8x0oh+qCwOcfzezsm5qdfKAtDBj+9eL
jDp5WmnRfCAacJFv1UomClOgrG12KsJVT+cjCBcKSQJdv2PXh9+xeBDNBcKwqrMMEijICePlbaK5
AHAEoYrV6vP3ee1HYC4OKa544lQoTxGBt1hoPdB8zNFHCpEeIUqoX18f2xW/pecI8wqTInKEM8+5
3aAtktTnL0o+MqUzK9wRUIZTNLe1tBhQwN1l73dAnvagwCVcLP1ceuXXQEEVnVzu9YzG1+SBXz7E
TQ18MLLJV/wTuIOEztzMHZ5LXLq4aNRiZPlFWWHVcPt3utTxmlv6pK4+YxPchM8xEv02Q1WJrqEI
o/bX3bKItoPxUc++YLyQW+f9lvLBBdFf/GZkr3GtlClbkqnJpvQRgTchS7Q3RomlD8SO3RSVDDsZ
VYUjdO5jFsMVOKXfTtl13AP52AEHwJbeclFfa8h67oxPIBMY7XqYBAxm0F8qajHgjU308dlItWnA
/5Q2aHPe0Zo5YtHUbvzAlyiIOTx0FrVAAHk9ruBiX+44YFzSFE/3Gx3t59KZ/7PbfDUXd1A74jLz
zhAQAtugwFJ6mQoo1ain5d3hVS2yMlz8LJkhu6JmwhhjI7zjzlT34NqpNWR/1w3k4Xmf2HNhP5VP
6tsfAjHXdotTekBrDbVVVW8mfOc8e8j40ttmxLOf1R7puUCbBEv7Z0ZHtPxBZdVdUUaUM68h/1Us
UYHkwB9/pgLBwjdakPFEDv3StxkeKIEUeAZFUHd34WYF51/R4+LXJ30fcHQ8/jluufDiQM5njgu8
hJuER8SHadrIh0JCz4iHkyV0H7CYjyZMR1tnHa/Aqz+EWjKhN8n400d2k1zaeo9pEM3YRi6pXq+o
vFegk6+mo/n1zLrkNEtq7NvMK10nY8f8L3H3lZte0Dc74MjJffS9Zd1f8Eepo3teloorwk++5Ar8
Y4sMiyhpjKxYDR/A6IOMtXuVFQf2K7UFwQgZzFVMKx97BB2oeRHv7+BWzypHw4e5zb+sPIuUz0Yg
oT/Ak0Yr1X0Tm+FX9N+RvqOnSji4uGDj0PP9s2Dbl/bIAlMmXWv5uGJtaMeuOxMZJzaGtDtegGSQ
b4BJxXxjPOLzB3EX4fsTZNvQGsOMgHZlM5aebzgs90uftv0W/bcOzj14v5ait1rbRAkpgc0/2C2n
KhiXiZiHDIURcNTGK45LRwWfj2WhiP9Ei7shDOaLIxfSyC7sfcXwJd4JKHH5GME0r06pCvwiI7LT
xKEbq0/W3dHnGs8Fga792LULdb8vG1pfGKzeFSMQ8PyLyGb4RfH5RLpEFFrFp2Vsu1CdslsbvX4L
ypUNI34+03hLrBZY/pfmnzajAK7wWYdL+WGh7Bz4gkjSHCWpRCpHKL3s+HrFZ+jrIjxs6FyYe1gY
YRGkQz5FJ0qKyXIQbXEPi6l4AIeFwxXQIuVVRYt8Kd8EbngA692LcLGADzMM+b3/Ro/KPxvv8y5X
o8yMQpcMGNVtopp7DrEjHhHW0MaH66whnGr3YHkX4fJma0OpcBSBUppktHav+30AEw8ES8JgGMZH
x4PytfRNvimri5zvpsk1cMrL59346D5rxLJ47N5zUBydI3ano5fuF/wG3pg2kddVz0wI32oFvL2S
y/TxW1EM0UEJ3fJpTuX6zdDXgZWlQ1pn9ZzTBbR5I6d+lY6o/z1SMtv0Up3xEJDEp/gstgZbrOqA
gp/z5XtazLV/+9pyLWE+rkYCSg6ZdAv6wpZfkhCSDhC71a+w746ZoUsNTJzw3/sH6A4YnapcptsL
RY6gAmJVVP0eExxolvu640LADvYCjMkQ/lNBgmRkNKI+gZWKzRU0w8Osm21F5SbnPSVn8GdlzhLp
G6MNkKqi+ZJnorA9YKxYUzyZjFS628pAMso2AzhjZvdT2kqOJXEFDd/14DONzVBbo7ptSrRQlpzF
BFT38o3PAcaRNn1yjz8qmZLmdqIpUdveyMsvBPt1Z9/KUmLIwFqP0wuxlKKOmrSmxZgM80ZjXF2u
rcs3ItOmA+6OMosizIjnYZ/+O7LQfBQrni+e5JJTMURZS6winiSu3GbfPbshz2WsQZJf83NtBDpB
Rrdh6o+IBkZjBh2vQ/2u28G+4ham1676zQXrg2B1ZKdYIQFvOCcJUFxzqxaOZi6CCDOuWPYLzrZ7
tZHcHZt52IFZz7AWYwu+BYri7RVPlUid6VokYemOMxki6Lleb3Mux5iZwLmIbjvVN9gYniqYqpIq
7Fry0XpYJCScRp7Z20mqIXN7m0ZDSJ9c7VHNIN8sLEBc2bqpuFEGX4/0bbKe7bQj0g+9nvbY4Zsf
pOhAD11JcEsUsXiIVAhG24HmGI0e3eIMuOkTU8DnM8eGzbKPK+olwgv4VqULw0mYEGUP6dR2keov
PnRAru3SQgxnW4eiM0RxRoCXEpZHGRn0JizugNjynKqY4parhoyLl291sW/9HJL2CtwxWuxeQEMN
oth3SiMnD32Rgq6spzbsSJM54lO7oerzgvUNkKvicn+dgkEX2D8Yp5nIh8n45N3F8R5facxlHISs
ghHqBaGW/Cs/xz/QcgneynWgayjXxmJMYkDP4aA8svfadoMg8H2ofUUQ090k5LFecDCHxL+aYaxB
QBlQbtx7tCusgoONI4jneXdY0xqAawhVLsY5duLMhA/y1ca3pYMIR7gYoVRi/gbuVMwzqek0VCKG
iFPrRIYzhjiS1DYh3R8uxMIXx1L4LYuhhBLR9k98RNVTGmmFgJ2vxJxcKff8zekNWkLHDNENoo/D
sUuDoCWDmLYvXmlsVmyGZLgCuGaxIyJ+BFo1IyzoegQYYIAkgNvQ/h9qnsqi9+GvV2WlfcflTIlJ
VTN/0HQuliUHlSTXCBkVnjmB76RRUuFO7Y0WuW75EnHZb5p2lvtOKwL6nwfoFiVSBrNUSsttoSuV
afTnBAu+wK9Id+bU/13rLaDpLTh+CJABbmQpLDU2y1nUgkzzD5u4LQf2lhxC48sB+i7BqMdhJ6Nw
JkQiMScsWHKeFE1F7nzYlae4YsflVzt1dRThQr4y6wUK/sBEFAxR8edOi0sJCuTukWntzdS+0EWe
8EbRVIAoh/1G1sf7UXJW1p6EGNnlGl+rqu5Mkqmmf722L69IjrwgJycPzIZGDhsESK7AbeKEKMQm
LhaNHWkV1JiW5YE4fyUDohUZHL0n2ZSO2Z9c27GmzTkYWFGFwGRxieAAdTdA4lxblzes8sbjsHoA
t4WP13SauIavmETMrZmxbXYjM9VtV1PyQFNG6mXw/EILu493pVj6/tQjloFgIfbhw/fZU4lkt/T6
JAf5rMqTB7SyctOZkU6X/8x59ro+6JB99udJgvja1wV7zWQ7oEqkDtVndEIu6ZaPVWN0Lkyd2EU7
/Z/4XYP25yqKeDTI9XMXp+X1Ufh5q1nUHy1TGMJgymdqccP1l2tGhIc6MUqy/LKqZLW9N11MiT8b
yRSvCkbKd9pxEEz3l6TySMHFXJdkwaw8mKZjqmVYuAg13S9qvESiz682L9zBhqO1JkFVY61RxkY1
qtPsVcVaZ7467W9ssTcX9mZgzYgIOGF4ypM8ZfSu6XH31QDmaZcSUtvR2UBf+FxFfMPcTOETYzIg
OUGr0HFIh64fLMMbBuYGVfO5bEK7UkDeraXkewbmTIchzs6j8/24oTz4N083d+D0Pxky0fUwMVY7
gv04wsuiWkfyOhbuIl1pdzgAO+LfACgWAuBTJLXkWcoVa1HsDMMXjn4BjPj9MGQ6UKmMhETy5Qm0
0TEt26VxM7GtMftDLLNlkZZ2rn1G/cPjL33opXkn5GT3HJGk1s9FJp7BeLCYGgRdu9/kr+ZXOywR
kyYbVBaoNvOpG1g/XIB7KnzD0vouJ7UTnV0yi6lpVUNshGVA0t5gP6crVkeyPFt2KQb4L1ej2sh7
gkVX/E78QBwuCmv3YZSC4XMWMjLoNSvvVTAsCZs3EHiH0+IRO0V6+CXTP0aiWHr1r94HPH3D26kk
+qLpA62/lwQa7cDLubnGZ/45OjNSFcrqxChrFY+1kitmR/8y2Q/Aw9C4tu2EUppPqaxnV4LmVaQC
OY3HdO2AXnY9sbgmd6rkw7IttOF+7/MN24CF2vesXCHVUUkO+txfQWyMoAi5EY8qoTo1O5gWpw1g
D/3EuRLf8UC49hRQkBNhSBe/Zg5lX5k2iwEri5/L/U+HY7kCnDlyX8x3HOLVbZ+jve+OB4v2Nu8a
S0l3Uj+oDzCpCuH7GVdIITMc1Q9FvQk7RjuUmNwftZqLi2H9+CD15iVMC541KqhtEnGUzL25oLOT
m241UZvC4fOmVkua62Hq7oyU0Itcqj0+jUKatSR0FT1q82S5tsWlPP/LHzsMsSXbKR0Vv177hBhH
F9xWHjh4Z+uYvkhXyvyaXshE01l/Zs9EGw+9Ykg4toAjLqIz+aKIrUl0kXTCh8eMd416Y2WJjeBN
pIMWTPlcyXg42vffQu7+5OXiJBtbjbp/sQ3MdF/Vstxcre9RML19FYeXgIoFxlrhDG1tLDHC0Z6k
8oNLfv/2HD58DpZhdAtjqnqVjOhU91YvLoPj3eisLQVB/wzUGg6BiV7RoEZD4c4fzQQXdwcud6HR
O51ukjgpQHSwSUsTZOpObHSjoAQSUrn+BfekeA+nI1Y+lxf6w3ACMvD0hZxwfLXRHfLI6OADT985
L+BakjbPNg91UMIGaqevWj8iOLhdtq/u4BXzXiutJaxaM48NW/7H2uRzb2EHdCFJMzQRSBGymJya
kPHtZpgZNzAsjHp5WDQkj0AMqRqypUnY/ID8YGyB/u3Hqh9hTjsRlJ6YCdZLzunl9snmqmQwEH88
+qiETA/2SgSLhXu2rwIv6Z2tNBGLRXRkVlSJmRr9/y4LyC2x3cD9UyXKhp6QHFLSne9jQPHKacIK
YIkId4erSLw9vdXo+rSBvkZRkrcKGsfM4SEoirshzrGfWvkS/UkQSZw7Nw1N2x4w/Cmd39HwirRE
ArMnCfDLeCxei5sTjGV/7Rl5RMs+ejx4UlCsY3tYFb4qmpzJcQJJAE3jVMIpzFtd+6wT77gIwPks
s+fWrPGinnsDssJdS6YF5zELXSj7xrndWEFB+6jC98bdr4eSvM3RU4xwiWs+VBYaIQgAE4xYxTj9
iojp7PRQmhrg1uOLZGcaOiTjqNw9HtYDbpTRXTjqc7d0zpwu/Eou3thjEi6wAliQ1bK3xUwAykGE
11tyYWMe+LxM3bdjIWv2jkWd2M53ZjBYkB8QZs6QYH4UruPOOQr0yvtRqxR2uR5luAC6Em+CLlmN
fA4yg8Ej+VfKacL94mtHvwOdGumRstxCiYPqTCwZxIZiq8hGpDg1am9quLU9v8mp/dpsO3+5ZtZb
7hSZc43EEqny4fjWO1NwxSjiAD3wIFB+sWVeW7CvpWrGn8gmdr1MHj260yhynLtq0EgxYAKfRnet
D5beVWSOCgBWeq0xaHmI7sIbFBmyTeHQgUguE/ivEBPzisKXDt331MxBFDGi/0KVwLEjV3p0N+lO
Lib5qWM4kGE+pOrQsWrZklHlFOmXxSmLFP3C06/2I2q2rLgxHCh0Cu4xtfygYcVLUeWJtB3CH5y+
j+UA8AKOYhy4S3khVf4hHoo1IW9aq9EXy/ZOdF8IwjMVOsN1TxwOCf5Q9zDzOC4pSfWzxz7xJWIp
7xtuPW1WSAb4wLvvFA2UQxut4DIkQDotp30XrS79Xy6jACVowMklmE4+nJ6prjgti3ggrUurPHzu
ufe3kzU4PkDTmKsEdJWfMD+0JQRmr/N73GvsPEZlJ89JOo1+lttbGmlY/bLgp4U3pVQ6kcNSxiiY
0IbsjACiSnZGKCiwyONPueUwDgTe+o+wuBVCrAmjKyxlX/+04VRw8u74YPjZGsutaNQ49qW4xLOY
q8EnPCP+KotNdIpKAGAslQJkYin9Nzc5/HmdJGR8wLg1iJlsQPUYx7ngaXj3hPOyldWVX0/H6v9Q
h5vQFIp4DLnLbLvbl9P5S3CG5jF6kZQNriCy54z5ogPP0OE4dTBEsVRXaPHjFdOHJBVCZU4RF+VG
VFo0VmII+KeXn0cGSOvGsvzMQa/vPCci8z+4kuQVudm0xO26YOrBrVCAjcyGO17MLaITCPLIcKKP
3Y4VdZ0sReRMFmmiYV+S+wsBChVuL0dZLXlJ6V2qSWajBWA/d7zb26PKnCbx0+aPVUf5DLjwRlLh
JVF87yjKf+JlRn7uz/eSWnbCTrJnYzNWznXAx4mTkhYkgz9YUxbN3tMyvtXiHgKZYq/+qAaZeuJ2
oU6tiWBsk+xkpUjS/DkJ21zrhvKya44cbdmMrDnexPlmUz00MOHie8c8a/d1zzmfe6nRXWEr/WqX
1ToWGsarud3hp9ILOsPsJLrQXwMGa0dfZ8Wz5cKeR5ySMK7pILWBfTspQwlUPx44dKvXR35LSOU/
hsP08FbNx+q2277o6K+Of+h3rLC4DbT1k8pNQk5FKmtygeBfSaptq2nyMq72NbyA+23Dj1EmUDCZ
vF5E2m6k6XN/kW7+HLoBIepebsN8cbX8J98YtzhwhTeSIWqlCcfKr9HWtpKmjw4+9IlRd70vGR0A
VIpUDllbnQEvsCUJUUIdn/cO8ZwAvKP811EpLN8inQBJFF0JSsaELc9conIPmyTKKrdhHau71qLb
6gpdUICq5saZSd8vp40zxRuXf6VxYFBiDcAwBqca4V8gTfaktJ9+GOsZynN0IE1jl5YIwtVSne3m
XpSZ5lCRPXqzKWjze/OV9tiMMH6PoaGZhi8mPC94hInKy7krBN6lt/qmx86z9arIT3+mU1BlYi+G
5e4V3D86UmD5CeUXkOPhAxRyT/kHWqOn1Jvn9jgl291uL8ZyyIIsaPZyiUuby/7jr+9Qb/1Ib/G/
FnYUx1eT5DiFftJsOfHdfsNx89C8M2PD2UmuuFdA5HZRJKuyeLP6oCFJjkLQ9Tj0sis8M1WJhiwK
noRmTw/WhW0cv9aasxudhA/InqWU427zwqmvyc6y/kDGwUdxJ5kQr29fTKPJ6SFuaw5lrI/5gvye
83nyCsiAQQSTQlRjX3J7ZblHcu3CwMDqEiy5cre07lj/n+cCVe+qBga4lvm4vSRPyKpCUxIG++qM
ZrkhvF3iBPRT1fTcTGjron081TZUFDwZtZ6qtl3FgyRh2bejZcpyRUTmgrmO+vIKrzdEavWStokz
9YlRa0OkFGlpMQh/+rWn6RhDRyhDD10ayVUozfY0a5EVLmIwkSSIu3mv8r4vGErS18zI2cPnZxVr
/r4HdMwbho6ZaPYoJxxBRsXRsCB/tUkk9NAGB692mUiDbprBU5EEIQPUwR9y/9TFf5/PRFacdn+m
wBx618R1a6EO3PXJNCCUygFcINjwntTnaiz0DsP3rPySBVSGo+0bePNSTIuHcEW0ktrt/E1q53Ln
4z+hz+nbT8VRdB7KhezVAuHGXnnX1rtlp0aYxOb43OwlHUWvVVnsFM8DGMJ6vFSHQCFLFKkBh20G
R0R1mDkQodMEA+aXQYgfTT0hs44Adsk2iC07Obcuxe3hl8WTHPf/wDVgVM2nDVrUE5n9NewVENe5
MZubR4i5iKW3IJZsy/tfDqcF53Wxs4RdIRdqMroiieBnhVDuD/hCrUtcaf6ijOpl50Xb9RUlIsdq
rn5zT6w3UiHwUZaS3+FZ3vvcBIIV9+nW1cysKaf1wG50jSMnwlE5SS7r0b4IWwXVsigAYl1eokxS
opXG8Vn6lRAck1vSlOqlzIaPF3v0e43DWGt3IMQXA2qbpU5pYwR8GtbmNV5sVIbvxGjrspI8xYAT
bn3Lltg7ydQQEf3IT2gj0U3QHtMJyKAicDAZZyew+W+oR02fMqxbpZdfaXOr+yXUlRYd0cm5Q6d2
sFhjfJR/HCrZxTl6uxLeiz6ViIhsotrTQWP1VtfOYYLV2PGYd9tptqC9WZ0DfYE7XokQzisOLGmU
exlAN6gAjh2cmVJ7Ymj/01GKcJXeAw1u0X1uFoKqNdp8h2badd2OD5svYW3FTqzw30G/OBC0MDEk
lcJ+KznMkosvTITlcKOWiVik5QyEpZ6tZ2oNGAO7RThCeWa6YZoxm5OCc/35y52EUaupJ+9BuDMd
JAxKdhQx3cO9WHa4lDMRGRkdy1xIqIgmydi5rIZSiJI6hTdV7HjfP3w+T4d2VqZYGDIHPtgXugiT
XydkXKAdpuiQon9fOKxXTa4SEVCVFxxeWbz2+/RBTPTSKCYuZFmHkZQN2nihlJFDrI4679G70Gpe
osGjNgiebsSs0rNuUY2XG0mqexTc8byHf9aUtpjI8HoNATG68TsDHSeIj/P5kTRQKFAl+TKlUyhi
6PMLHUDjWd0NwR7Ikc3i1ainuSSKLoEdWFB5aBWPwcCGL/y2doZZWt0AVmhg7ZAoG6+9ehDuLbI1
Qb7LyudZRxniMKiaVLCsm3FT48ac/zDeZSLXoVcgHAEzpxq9x+hsDt3MoZScxq5yFuzxPOwn0p6/
alZkZqLO7gdcX9T8ippQA5DRtuGzzW30uePzbAD6ETbNMuHKUsnAF4pTw95XBP4WQwtmriUMLHK8
jiq+KWFcJWgwQnCY3ND8ry8WEaJdB8m9oHD9LYXnJOj5AXrs7Tt5TJgKwzAkh77ynw1+byhaCqAb
81APo9ezQm3m+PLchd1kPU+2LCMduKo5bPCwXPINM3zhNaf9uUs7hmFiinO3X+5/Vtv/TF2aB8Ct
cRB5HFyiLrX7ezvbAYNEVITaewvJZrFAHRi415xdp2D6JYiVh32Yfw3/dmlv0DmbIgDNXWzTo620
NzGRCA47p/FJ3dTN41LshIfICxKgZufLilZ87vpJSrC0D9QZlmSwDYeOT2N62Qq59OxgER8zVLXq
7tWlx7b6oqzhHFBAUt+uIiqSyCeu53lAStyLVWzNupGncV7hG0KvytmdAOMCDeIv4dpnCft6/f7O
HZrVFK03nO2P7Ib/v+hYAetOOjeW2/rC8dZJ2ujYC6UtHnDc5XsAU7gI+YYHItvs4x8ZF6vyLrOq
pFal2/sf+4hJhKE2VbKUrALTjXqUVe/a8XwhrBz1z9nzaRzKKbqRdv/3UXtPI9dPdPmE8+DWxMWq
NAsbOUKrbEpo2Dpf/DPoRMo2tu/KCJR/I8k9V41jYW2/PblGdVCGVlgZJhI+nqIUCHA7zgG5K1lo
wHiVmrqU+IpAKcvtiY5/fYi+t6V895HFbZR6FBcjC0mMus/BJFNrj+gW37hTRUk9pyFtGig4RUzs
SzGpq5O4fV8QFME0Bd5xVq/ZMAFOwWU6Azhc8Xid4kDG3b0AUsyDwF/vJRvoOCAD+/w0jvVcMfTy
OrFgiYwvE+CZ3WV1nUthfkl/dGlL/X0kEktfnWcyIaeSF+WUL6VJJv5mkixMQ34DfJgELFiu2g9W
dULyu65cNyIhlISo8AULMBG0vLDNe/JonVHxdIBPHB7F4iLbA8pgK6IZYjFG6iVc1FScEVJEF3L0
DyexkIGii1sAKhS23z3nCvAjtRKPzeMBo/Z36KTNeLttWLB8dq6gI/FZJt/0K7/neHKTYMRVdP9V
jQugWC7BWa0iYIMkJ9T/OigKkqEmPl2zhG2BtKcoJyOyQcXWl+aXcrkpdz3PKBnfKFAKjElx/ZEj
pV2ULssTh2Gq/HF5F65to99A7A7ETdCmNNx4Klv4uNRzun3bbTmPMJlB+lL72Gi4NSanQMvN1IO6
BrHEYwRICIZ1H+nHC4AfBG4F2CoDSLG0sSQ9b9u7vElP/4Qj+0zzjm0e+9mh0V6NJQNdtENfALTg
QT4FRJ43Vf2L3hFzM4dCnmrQ4dHJcfAAOXT7J2U7bauf8DLT7soWjl/Q31muzxGo/E9SvepYqcbw
RS7u2LOVQX0DQf/XxxAWdsp0ThkdSlyP6b9k8+TA3hiWPtQMSkdtyiEYn9cjSJGYDFdXA8RVGHjw
UWFucUcB8giAXZVj429sln3RRBjSYUwebzb6H6d5PBVSp5YPhlRjg6sAcMUkKaHd5QFa51k5zut3
KkAEwvlSuMnJPUpsCwU5+ugOMwDsJXzhqw19aBgGajnXeo3sH8xNonQYuTaDRIKy2zGWepLZ56Gm
gqq1ABj0m5N4puU/uf+bqxLOkHnltSDb6fRArIagOEKzJ98QI8BEZ9CMloCUJ+A+u2wMKDLvkB5H
DFY5qEYd3eVbS+bt4AJs1kRqRgCUCUzkqjXhZDA1BE5av/IwsTnMjTIziP4d8L4DiCuAHUwxLrGg
/3wPVOXZTRw+WYnPeVwycwq8YZnBINRYhFAArOmV85A/Koc/5fuWYzKG8uxLVmgkpCS/Myl9N4hh
pemzK5ZGPA5ZhUqkKiA9Tsq54+ebpj2oSWDjLh6EXPurw7DL8JvKQ9lGR2pqFRgPoBPrshQE7km+
Oz9AVx2P2rp+ydoZoAEcg4PAjU4cNVSxBfcctHHJfjEEeyYKStqNtqHm1/Qh6BOhGdAfRUy2sBRK
zyUI/SfxL9ZiQHADjiK4hUOEZ/qMY5O7oT17OyQ+xPI5YzFnvl4g7O3tpAl2YmGqmo3IR3ZgE9fg
YzSHp4oI6Fg699Stf8lDx1tNBmwsu+Z6vK2ePD+qN6B50DTKgtRCmAxjLFGZnCzFq/23caBjxRx3
cPIliaLeFxnEK76hheuTWfRGejDmXSDZE7kGYsWd+EdkdEXi6cZHChyfB3j7I/LRAE9wUtB5VrpR
9SUkoxKcjdIEwzS5+iNST0MRDMpUruehBWvPi/QI2CIHcNpMO10GnT2JQUNoBPArlFk3cYbca5os
TPw2K1lJKSjTlpkz05RMoHaECikOPApQYBx889VNEzah0j29Gw0WMDbJ0z5tTfTLoSa5u9Off3Dx
eFJmogYUe3Wj+AvRK6de3od2LWwJhTgBCXFRcABsNVtM/4YRInP4VBMPt76W6yIbVos6Psa64otp
9cKRKZboNv/vmtBe3q9xlq2WShZm3Exc227ElfnVmu00Jwu+TgQrhinQBVlOjUcIclDOjg+e4hsN
pZ02AKdhaX1aoGfAijFsWtUybGE78HgXCOPGmVoObMPc6CPBxJmeIKl3rCoZK+23/NBy5cgzAWGe
z2/nMvxtbcLRs6aZLkElRJ9ln90vm27W/5lbiuRMu6hzM7UnMNLrFmSMqUxYMnXKvOItuFckRxWg
Xhh3I2E9jIpbF+eTNx3WiHd87e2GTwug0aB1NxNImlXcuomUVPEz6ND0dDTMFDvP+iHqrSZHJkTB
rCiM7anAJ6JHAyY3HtCAFb5fSDgT+1mqn7mgS6QCMjWXvWzyTdOKIRbeiThBRxdQeEGkVRbZMdEI
HfCjEygO3/YvQbqkXb0xPDAw86LcKgYFEjwAkIVjdUlYwFe1cKQwal8gXRXBIAdTqmd/Vq0ro0A0
dBgJYVB61FXnNd7qcb/NzNXeKWfb2ZEYZI8ENjjOAmuaJPD+0rlLq4d3SVEtob8BWppU6lTnAl1o
04lBcFJEH+nGXxCjZ3+FLOm38BBLsBkxNbXOskDyK0rp01BUNx6V1MioXcigMZKWFfOBgcDwbrLM
akKI61oWYrO8gHwra7PPCRZW3w1Fqb5T4jk8neEKmDKzMy3h9qZ2i7C3gz6sEmjEz/kQe1ZbSHvj
GPQ3OK+ba8uwIOPaq2VUpudRBMJVYts7SoAN46kkfZBObLeNnZxZV6DtWtX0ihvH6HaLS5RVGuCA
PCXnalBbsQBnWUVeHOYTwHII7bi6CKV0U7pOC1NszVcqeoHa52iJKRtB/PNYsfzac7aFkHaRe29F
Rn6+jVMM2W/ibrQo1iHBGlpXsF+fHSB/bFo0a63eUmjT6qrkHcbcF6JMvTdLod10oK+q+Gf7YE7U
G4iHhi1k07eePbVU1Gcre0yNo+f/ZgNqFrR5Mxp4RlD50QYc4KI1qfySwI4wpCWHIQfOi0D0pisy
SZ2ACCI9MEgV3nRa2Xmi0HXcdk3iAvHwFauc9/FUo+bGPXUL1wb0ipi7DzcW8x0BJsWj9fKiZgoE
voc/TpeoDmDQ1QdTlA+LuI8Us8raESj8dY8LHtnAcL0lpkEIY5vNrXng7P+kk/AAxYVQtGLDj4Lc
7yp3LknwAFa1X+XgiRnaUtPLBJTDdL7cGTAD6FTVkCRnj/t0BQuY6SYEz+fZ1wZgcuAXakuzyESd
H2AE6eHWhucW4LzFdRE/dc5HG4DlRvryQxnrR17qffVQgC5HPBuNQB8CgYw/jsvOkGQ0hVNOrrc+
PoUNLsZdi+zn/7P4rD0O5yq1xda+rPdFtdRrZhkaAy7isjO4Qs9cZU6sHY2EcPuWKYuL+36eKlWt
fI0av7gAHB1fTU0wixaTDRkjCwJMNm6mn/fUAnrP7ZI6a70WE2PmUpSrf0qelc8pftdOsGNONEJf
zpZ7CNpeIPo8gALbHzYMVELW+WmURcWc2L8RlykxeymBrQT8yM/x2UPF7lYtkeDG5TbpHf3uIYmY
LoUruom2tuJrXequTBJXWpPLS/bUDRfYR5DxyXpRP2gs6OIVPL64GcPmKPKiQrSZKleSPJZPe+eK
UIziybvmTDaExYOEcZ1D2no/1B/Jhxsi9Xgl3d4akmtT4Eyu/1dCi6gOpW1xU+SyNp4mWaecI0BS
vWiJucRUf4l9wfjroTMs6h6stKa0jO+WqKmCAt+zYJAdtZ9I5mO4XYbQmrEeei6sK2uy9WSLqySn
UFWtZPjEOPbqUyvEthtW1nwO+U3YYkkyohzArz9qEsY49cW2Sa5KUW7XWWsxJX0u3Kt1N6NX9pTh
dQ+bL9AwoVDHSnBxGHNyQOg3rRRTKofgy56TIoSDXJta7r73NqszOujqg8NMSj/wmM6NzW/jmgBE
0KQnqNtbInylzVm6f9cH8WyQY3qfM49Ueo+HZOHKDU7IqPs3Dt1KBWijtXO8FYKyQLg0DOVtPfh9
vHVjbdSETG/D5HuPknETFha/sWXGWmb+rh/lXqSS3bM+WnB4WEMLL33pZzBJAo8aMAEme1GD8kGQ
wfN19OUoEIfKpUBmjVKBQ7VeZfum3qTA5x5tz/lTD5GIFh7PolJDbn8XUpnPVezxkFqwVIeK8Dvr
N3WSMSuKG9230RRMiexhjz+5Ns9evtnaAGaokzvm1ix7nnC564bxuPAsyC9qx7+4NtgrUL0SG91O
raroTg9rO1XMxm1J9JFXf9VqCaUU4S3q8Wwf5lMTZUbiQt1f4W2qutqzEoiSWIVApE9j342iyF9k
xOzumo+DmaCFW6QRCH4YNfKnbELKFjhI1J8PfYHHXozys8erIPRGoZipyxjwWDhfnA7JdzGfEnDM
cb/6QdbBphEUVsjSY/KJcHD1LqNvkOObUPFOt5lymDDtUZ63hLkqvs3DVbn7VU+k0Aj0/GPy02yR
fZOweNa21iwLzoCQMil6gKjQ6HFbwvoIQPL3tQdYOElb+S+jCyun9HLQbn0M4agKydWR3ZaEfxVE
gL4mMm0jBMKIcjWZsN/7c/MnuxSMtjeQ1WmVPAx7+ANOMLL0SgxD1gHMsM17HlHzSQ9OyYlhUY2x
OYCtKwEEs9YxNrH5hgTrgVw2TOQ3F1eSSxHFj93fSf+CRJqjREkZyH5/IULNQ492cw6jiWgTSsjw
BRgB2Vg7c1/im3h0Kjq1h/WtGSCMUcQ35rOublXodwq1+R+1Z9hvqoh3nnxHHXu/qPLCEadP68wo
MqvmHiIlTuLTmbTDyith7hu3SpJsKo5GkjwMhBMvHqmHpnMcfi0wsPv+kk8LxKUOM92jwWJOm1x/
BTjuhgKmSgUt7mDZNNCYYaiZy9uW+6siXevdwjVy1jhG/2KvDdsRcMofCuH4ErMko8GQ+x1SN2ry
5cqJzdTxv5Yyh1YGZlFNr2FFXh1qCKkqtBKejrbBPQVUOHq5NX1CxlkmUkXF+KIWDQiYLWpe9XX5
mAv+ItkD9RJ7DXSl6ax7a5rETGMzztfSuIFCOUGro0edlX39R3Pf5gbk5P+/bQjQfVCIz4U5Uao3
KjOc6UC+9d7p5wojwS+WHhvAYAvTROxjb0Wd43cHqjXv5j9PmCRmgfdL0ILVavMgkqXjbwxZgn2Y
Vt+S5U3LaEszgQUNpWG0AWCabHZEIV/is/Uc8UeJ7cl5ZMCboaiJiTvC99m0juQXrHVnRcCue7kp
S5C161TrX8Ia89keqt2iJrYiGTBgw2+BVc0yRDTV0Jeb5PrCdiWvc/pwqIA+9O30Pag00KvarufP
sHosqYgfzR6sAnQyBfgZwFo6mz0sg0YBeWTdTpFkl5BxAD1nu1SLC+uBPFYVEaIUNTX2aJdWTI6N
KQyxKEvu6OYGpPDItiEJazBVS5L+9gZgPPZSIvylCYmhXePM4TGu/y3NIyQt9Na4c+ubVC+THcls
zPaA+mx+mTLZWexDUjt38JbLOaj7o443hh/ny1XBzERPw9IhhNWK82zYQcYc9q4thUsPrIOVQzp4
FtMdB/+WzJ87CbFPk+JCJ/j/8uk8nKuOU1VOL+VEIY/8HycxoWsRckTOVkt6DhmEfmd0OXnheX6+
NAH3RdzADLh+faUME8DE37bpLOMOuXKxoA6O00Bk0CvD8KD9OiQ9q97S0V1oSfzQQbBDuvd7MM+i
D4KJFqva5T7XAhtsx9LpMsugCifqVXpNLMoIJRI7ZVe2kZRjvU8usjK1LZdOr5ArqbPPHltPsEBM
ihpz0r9zdBZqMR7Bikm8yFB4FomwQwgwbyZ/7xjNMswkIK932PWcEdUd5+WORHYogLmdCN0N1uPK
cNdbXf8xDiK2MfqT+FmtTVbbpgd6Lv8PVxEoJeDKpHwc4po7VXFEfl9Yics/EZOfuU7Qya3tJFmi
zhZ+vrmymMhpAPVMNXeRNhjDHC/xK+a3+VrBGywyD3P5qV1NcP+rFn5yTM/7+Yw1G8ArT1lM7Y0x
cVLqzg5n5fmnrFE9XopYtAk38lnRwC0fKgbwLy8F/GgZXE6YFWkukPhHeH32Y+6p3TV9Y6Xc0H4s
Um6ZqGceDdDlhHyobCRG3p2vqq9/D33QJjNsKWLvCCn2kLjVG/oCAMi9Q+l8nHXOFr/pU2TRMtX2
jO1gM1dDSz3jLoEmmDYZTabb5Az5CIVNHXhUMqc8gWgSZt7shWBBI0fzs7NBpM0xwtYtmiqUszjb
Pp3zYjfCnfE+Lk1qMCLBuga4hlvzahAvMewbtWndDX05Ps/C+4ouFsXlXAUptzRMWa10W0wpq1jp
sO0P/k+CeGBvQP1ut0Ej/Uq7H75F+rIgreYT19NApgWEWGnRSbPRqsjp+4YViB3Mu5GD67cqiSEP
KxqO+F18UWYa7YrqllylCijad1FrGOaJkYAahTFX+BTyH26fP4NFihLCXGn22XcKsmPrLOdg4GV6
kdcsAA+jJl7TYD2ZpGyUOjDvL6QOAL3PS8BQi3qXHslL59kNSg2cuseQ5Ha7vN/xLg8fufX2DpoJ
65KbJuDKoWt9s4XThHwry35/yaSKmbLAJF+HuKdVRYwCn+3iH+SBAZkQCvIPD1PvoX7P6cYkc1wI
YX2v448yB9f981qNtTaQIwrnjKvUEX6MtiEkExX1T6CoPM3XQKlbTSluFNhfan6vqhhLrYYnNhOY
Ut7jGi4Ruh6HNgFGK7iM/XfWCboeam3W7tWrv1kmReRC9AuMHFnyaObtSWSTCLI2kmHNo23zWZfN
qI0XEIz6kuOqYP9fQ9H+vMXgbog1H0u3nyl9ZMmLCZFe3arHO2RFva0TJg9Wasex66BSfE7Dhtd9
aZD5HUMkRfPHSSOCJIQi0jU+Gf4gJwMF85NJuOp3pAFo4x6RwdLuenU+ZfRv+tAgJG+Krpm+reVS
j+J+GV09jRRi19KNuzMtRU4pD6KVxAZy2+qwW0DCMj0Qll3W/MHZujFIJIRqDKktpB5Kf2IYlDZW
lPAOoJ8LOY8smiI0mYbqBiwUyU7yRgS2CQAC0vL0aB6WQfWANlCwlC5CURUChxYZEV9xzws4YjmO
OP3qWSQPgTI6MEZOeXuazp2wCIPgAQFbO4Evec3w8BrPpVMncCko8w8U/cBn48evIafSCGBcq/we
M+GC6Op+wHqvO3tX26lJUIRVgUcnESU7HgMqV5LPJHADcuIsP5zgY39CF/AiMpwIiYIEKAu9PavV
0nT7Nnj8mHDwcBmcW58huKpLl7cDHRyUd925aFd3G0zRoXfGNviD9Bi4Wa76F2weeukxZ12Jt0uL
cXLK0XVwtOeZ0VOtnoNf7brEduRs/z5I7QAL2nlRLyatOqkUVUIZSYuVBjqUU9F0d/LH6tUjDW4O
0ji5cmpCWQOapRHbjCveyDLTqoZp1AOBj4ngJOjYnCo79JrmbMLcoWnVywKbXarZmtLV2qMLX3ae
b2HmqTJPEAtDR3CFV2y80jG4iJIT99BgjJ+EXSqlZUDrTAEG0JqIEq0bQYdum2IlMpecd9k6KaRu
Tlhsn1H1aE3R7UAeVWZsnyBKagXRL4q+s5RyMyWypD8xtr/LsNdivz0BsbKslzAeNx7Pt2HL2rJP
8HhtPEHcc0V6XHTQklTEgczMbZKAV/Q0h9JqQqdb5rz8V3MmoP4rJW9KBgPyN+RhZvxMlzlHgLe/
c4anYWBgb+JVDBvS8i63DE2wSG5fGAUmZybhFKB8r+mwUuyIP+S2LwQIrcD3yquZFh6tIUua2oky
vKY0MUqV/hlP/go3lsjiu8UTu7x/bysdE0pDaTe2yJzCDSGUNEA8r7KOHaNiyg/YnlwVFyCASAMD
Wp3OS7sr27AzAgoyOnhykbdXerz2i49jpIUWh538PCVk34f8iA52hTPQDvcH+niDc5TzERCYKulZ
4DDCzbZVNDnMuhlqyn0W+IQEEHf96f3baAC4DP2wlKeXasf8eknpttjpU73Fk6PDFsKMpFKB7GJ3
y6vSsuITIaCU3eUZq+Wx0ZQjizQs0VLS3bww0etXL3EMxPl4iakYk3LcvgzmtEbh1EdPfYudpbwU
SAf/88Uu5zzRY+4erncVPawQ6GTQbLjGfklDJiSJHrXB4diRxTY/sUWjzq+Lesc2YikyHB1bfJqj
cGDPmxHDFgAZMrvRrrTAo/EGdTCEO7tOyiDh45rM+GhlX+y0rEtddTTJzgX8uy9sTp17G/LVNSYX
ZYzJ9NHndMiGyDNJhBQVaXHkpsi/9HxB7dWFpUWopOaNk4t38i8c3ggn46PocjxBnmF6wBXrimca
ZhGprQl2yTOQv8FS2r/K/by/Cp5PH9AHN8LXJ2uNG0LxjrrLwgh0HTynEGckZwEaQ9KWbhlciSYt
gDu681WBLuVy4DcjjfMb4AY5yKccqP6s+7ZhEgX/vvKsEGA4S92G0i8eZohpf/54yV1HCorAw9km
FOplHkliq2+dSktU7yLp9loDkEM4aC/sLIqOfP97/F8IU6pExwCMktqgH46Qo1XC0eHWKldPRzMt
FKWeH738g/w3KkDOR/zLwQFJsuqsk97lIxHjZvBcAAhs8E2o+g1RqzAnhtj0dyFBr29T/+Cl9J0M
dUl8x3/cNeqPkp3HQqPrSAViYWs6byyZ4x5O5git9lJwj3eGB3u01X+UuNHTd040t9pSqd/pmfsm
Q/dJNsZ/3oZ3J9FX4F6zQ6k/nMlsS9/bhqstM3HuQ73J9hQDlWvQRZuGtMUkPbiiZKi3cJzL1hx3
O+qSXmiMKQNL272SJWvqy0UEWf9NDeNNUfZd5KICcYJo1yAK3HCejuukvOKSsAHbaI/GT7EGqm1g
q1SPBXNJvAXDFr8boTgD8M5X+kI4eukTiisDR7EGmr5DBQ58i2cYRQC8KSq9P01mpJx+rA7xjJWa
eR1ffBFgViIhjO3P7uxE2EXTAomA6nDDSTq1iJHjyjdxMKMrdG/C6g7IWmoKaHC+2lLF85gC9nKV
/PV7TYy121NY4zwniydQeRaLoMSmnNm1zGAiHPZnYuKV2mPlwAe2H7BXj1BE2NsVikwIuEc81Dfy
8W4D90MH0tND+B+c1QSUQxg4LkguW6qZd6x6WQ+etp3S+mEL/aCkovjklt5hooHssX3AV0D0L+Iz
ugflB7We95g6SK8XL+xaZmYetEXSY8/ie6jnK8rcjxu0bXTByhjAFDlmuT8C3//zvrq8VcA4jUsI
H9j7lnS0l1luRYrsdNwBHmCkv1Zrcza0n8hrjgWFqTBB/dgGwX6j/E8ooP+hWdfV0emvf6ctrGXy
aNgppuRb8jylW1bVg1I9WT0y3uLuN+X1GiIadgNV0GCR9l+Yn/4A1LsbSfubmh7qvfFK6Qggowdf
CaXyuuSiN2Edl/k8/7e7wvhW/FYuCPDvKRZVX2R3otyTlHSfD+OzIJeS6FadZsSRSJrFmfffzOV2
hv26U0bzE1IWMfqSQKERNFcmPXNhwE8ghlhB8qpjhlFEGBHj/Y2zaErPbB0dRwiPs9ALDhC9u/p4
jg0Vd2T9w+w1/3H8C8RAXzWGiNkdu186e9qyiYS1WlVV2MXD+mz2VRjvFnJqcjDgK/L6W8yaq6W4
NGe9MFp6Ko23E/GKKbv2o/hB/a1Nac0KnAdz/OSH2t31/rCXoUCDzS0INptnzDVJsAZdG6u88iVk
RvEdf/Qe+L6iMmDtjMXn7bCa+tEf8N9p1PTJyI5X7Zl7ru1DWH8vIzHd2pXf/YeWWi7hlYLfc8Jp
+7f7QmwUygs14R4PwhR7BXbzU7AQiRAAkGMA3EHkUxL1/VzL/UVl+vcAEFHX8KSvehouSRDzzDhH
wMoUGyNYlrFC3J2sdRnqa63rWRD48y9QpwftIM1FtdkueORSh4VDo5a3P22Wb1w/5D2VrJcNdACs
5Z4em3zCYNcbSN0u4r+AHB+NNWj5331O2ARpz4gUEQm69EHvzS7egKlXOlQ1FmVaHl3XG5c68SSZ
pCiiMbkV7MScpckq22Cm8cEtU27/ZBSsdQ3n4aUp+Eah26hE/EPvN4P55DsmbWwg+LF/SkpM1zyq
fSXNi5rC55pMkdlFHd51wdhwe0kUK4wRl31KWhkD2b8mqJXCS3PjEO8Du3U2R1KzpZQ9PFReTDr+
/vFsQHVNUXavdBiUTrJDMeB2cjd/zWwlplspvKGHAKD9ZFwVcWuF/ZU6QpnxQ5h09yMAyV9bk6mz
Pe1nLVf8r1ohk/rOYnhDex+b6VJ02Dd6OxZ1sHyOL4XBVaqpwpi1LK3m5ulH8eJT+y2ZzBQiH5Qf
RhTlkRKgIANc49nW/85f3xzOkw0M4vVhu96rU4bInTYRbZS6mb6t5zvafSQTHftLmNEnE4XLb+Ve
Dn9+RscdOhrwiWHnfl/OuopY0SplQ5imTF+HK21CFC1gmfya3hYX7olrOyNXywenCtQmBC2tlL60
LSsknvptjQ6Wbtfkxr2MiPhibUrYSuIOrXu1+pYzNKPP23rWhXmMseKYxjjGO+ZAIMBDcsDogAPV
K4DhXDX82J3sb8oyHwQ85DSMixle1+gJ0ooAvT7y4YYwyPiREbO2cNvTtIhrk2f1JBV6AAaVoSSW
PL0WXhtWLQqLP9jxtFkWoUspuG6cQpPKqhsNdKdEpC8ySjAhHtLtSZ6PqdiC+JDiDSk0L4JXnVb2
0P8ObMfeDzhtM/LooKfMuupJ4fngbGIfZwk7/O6o1GEgdemfouVvgjFjr5/fgLK0qYD9aNs2t3cI
JoVf069n+KVDWzZ/W5yeqAhCsF68UOj72mu1Spp03eHCs8QM9uR1Bgsv7O/UBjBOgkjxSh4pf2t8
3LdPEWmCyom1Ane5yYdIVs2QOddxCPPZlL2DkS7vtgjx/cgrz5ugkFaJMFzIncmemd89h+7+4U2J
TEWH8jx+eMUf+zxiKWSf8dkVonn1LUuYsd99q5iz1hWPnyZRUZa+wkEY+vqxJvbEpFDG8c7icy/k
WZhtD7xbN2iksOn3hhGzpbYUxnIQzclDBPtr47GlvyV1FWF7q4SjsnaV5hgB803HgaaWY9FbfgGa
w4KmTk5Kklj7SC8uq9uWwfnjRGEToUjzZGwLLj19LDoGfOV14yoNNgIs3myMvRYjqyYmddu0tl61
HMn8XVcAmVZYNJmnhLxymCEuin+E4iLRg8V+784TKCglh+qmARst3LZic5hve9rc0AChJmwkzR6T
poSKmH9JSSDBEtOMkcdWByS9gqMFeHlg5HK21BkvJCleUetDXtnMq14wPmEdNScfPFpKk/koY4f2
jXK8+htrzH3IYzHFQP/zfYx9P+dql2VDvHTBTyhu8arrNOUj5Qo5TR8sb/sXRrdc+YcrlcN8eAeK
+55AuTFlxNOXpslm8Z4ENnTX0w3sFbAODevldY7jYzArQrxfLmf3G3/M1poMPXbdrBJSFjFvngQA
u77ck15Ykpg74kofz1W8T0b/RC2gFOhAUUHef3bwMZaUlSqHNyRD0woRHHpTR+d7bgr2BcqgL5Mt
Ly5Vbjt0TQj2WdqaLadvTPbezaDsi9jFvgI6rZRnEej6PJqLOIlGGPXuCDZfJsKAYU09GSZdo3Fl
i6dyNWGdCTtQmOcNbzCDM/eVbiD9NFdAQxGeXsV1TKBSe27TnuYz6CvadsjEcID38UzLI96SgK2n
1T3qavb7ie2jyzDHeoYskX0h7ltLVb2HyslnGTmfghK2iuEWUg0cEoSgBj8fjUoZqUbiZOsU6hSK
ai6wyukL3TjKjyGC+PXHqhQETikY/EJyeq2xMksw8+BbFg+QXSdRdHuv0MS0Oaxjjta7gRCJ1KNs
2IOm34Ad7M5fY7Vq/4a3IVvpUTEoXCOyjm+eP8oSiNsgsghf4z1Ht/RFW6LBOyiU6dK0isCU2pL/
CYmY/MQWak6FcFZPURnCglnFZ4ciVU5DVeTUQKNG2K075zDCQgHJ/JUQAF/OL9YUGpIlnmzL3cNN
alNxIxvfSOT8rqQT23k2siHsZ3fsLFlophHxsiwKGCwEk4I1M0lYy+mbUottW1jGH9hUPjNXOO+m
EUzfkBVa4otiL+PlZTEl3JzRrbwL4hO18OJoQstG5OoUMluwCcWagpJMncL7Rm4+B3lBqzK29+tN
u+F0Jp9pgO1X3TmIAnQTcP0HOrhIxVlRooPU9/ZR0gqAd5xBJ91VVPvtRUJ9ukhCqQDVBb0cTvn1
72WPBNBG+Je2zv1eDSY9qtNR3+lHFXydBnW34kFfACTClK8UOTChc7EucLSFoCdTwwgv4LD1XCd+
YN5E/HA7BILcIk3Tdk2NF9cq8w3D+twj11FtzTAxmF/Dm5RN/GCIOxZktogL0oDEja9CrE69E8te
8M0nEUBmaT8Ufun6Jbksr44GN5+zDNsj0DSG/NpN8aOkDHIsw/pDT2A6T4BxopdxxLcielWGWLPh
Gfc/gxO0INPITMamQhd8GlhzcI2BN9lxI3wPO0u+0DxhnCdA/taNwzd44AaTtW4Iqg7Lc8XOKLYw
RcY0g+vx6W2i9BQq4BkiWzCgTM3+lv2TRpkAUimVq5LwSyh83ENQQjsb9Whlk33wAAzhL1/6iffR
ysCuE+U3PE+PooTktDNd/JKGmiT/BzG3Vrx2tOXu3UjzKdKkc7jG5TzVedpRC45zBTF27C11uc35
jHfhavEuZpI/busWDpG3YvqzCEGNoa3HTJQEbAIBC3xkMz9p5QsZsq6bmhvEEQieiBeXjGztKTuD
99gHs6ZJzALg+DgZ7bcuKOd25m+kw00hUT+PXErm6OsIZ8v/unJ4MzQZeK/1TX6lgLRgLjYZQGzu
63s3BGpFozeEnsffvFF/dy2FAEKPYd/TzxNVXyGKknYsatwJ7LkGFsyiKJSig5//YfTfyrULTDLl
SKVAxF85mZ+qYyccFx6zN07EkSTydyRVUO9Ohr2ZEy3WPfoW/n1ycMn1gwV2PFlExxWUC2+0UPhT
E+dwwoi1v8yyN2OnEEc3lv6pDWjyxNeSyFIvVJIK3csQdxgTgmXrG2GLP/8ob/IQ2ka4LwFVfdLM
CSKTluF1M9eNzg/NKC66AR/3RKO9Ov4GxdK7wtoEJmAf1WiZW6Wjv/Q9+wtUGyyoPrEaY9XVfe8N
Kc2PwJDy0P1EEFLVQjZqZG4QL23l9Ai7HgW+9+FoyVNi8eNy1oq3A+snhf/jPh6j9J59Z44CF2XA
QFgGrTY8ecCN4FrrrAtN03Ij7bAtJIYrqZOw2LDvzB5WQqFPfh9bI/bK+SvNL1l8AJHN73tD80zY
w3K+teXkv38wm7srbl9qIgxcPumhhot+B7SCIEviwhzdRaUC3BQEcuZNmx3pQbLzpV5kH19PdkUU
aBTtKuwKgpievRz0O4pxRDa5GSixorU8vOkQ6HZxdLi9f8lbmTKlRX1qrrFdIJZ5NkBdN6GeYBdC
NnVhF0e3fmP6mKRvkxd0GRHeBu7rZErjcvQpEz/DvmEhCFMiyi1udP4XTcfvVLqY3qR0mi14Zhch
6bDz5UEubLEsJGNsb+p3NC3lVxzTjDBu4UB4nfRGSNshYXIH6+A3K48NClGWtGcdOnFadA7n4m46
kWDIzV+DsNt+II0p7OgTdK7NWgcdpb0vkU2npymyIuIMHsjVVD3JpmnNqOfB7lP0ey3kUJGC9/ox
P0TccrLIpieYDPhPzIvXIxx4U+/rldwzicydKVLNd6VHZsmMk2HO1263KFuSVp/+QuBLb9QjSYrU
QBTs7zRN8fxAGGUVDoj4XWsSSFKJ+ZfeBAphJvKjpGeFa5TyyVYfncUfiQFUn08Lie2AxnDSQ2Hn
jOGHoDH+C4249nO9SrtOov8hp3CXPW0hp8LhtXCnNCxGK6UxxmgcrmyLseKo46I1jglLGeFpofaf
rU76yBQdJUwAi/Melh6SpssDA95AeNtujlSx7QNU4Gm/RDzkmflfabVpGKNNdVyWMfp13Q2Bl7d/
+502KceOZ4kNWSgP77DWslX3/m6UxOvy404R1jZu/HE8pmN6QhXnKL7Mc+Ffp3CBRB0B6pHMt5mK
0fuFjts61nIoTABEuKwDzTPAH+9WKZWdFNvpS3rHHlKXZzJFbEcM4gizjG96awmogrXzQZnWwjSJ
QUaY4G7A3hY5r7KYReHcCZ4BV/J6nkSJCDMij8xZtdS9ptNt1fSr48KPsp/iHpvUBRMHIt/DHouC
OApf7kAzz0LRWAi6Fe4YMACU4zOqY6s5vSEhIl5PBPJjQ8SmVOjU2EtqHSfujpiAWYj1DQWGEVzO
EqB+2z212IwKAg2EMXmLyqCQ547kriaDTRfL9bzUhKrF3TMRgXgRzpSWD8U+k1Gn4EJqXuLcEsST
h3XgvpqrFSNrwqkqVCW/NvVAsxAzR6Q43BuUhHT9v5+ppCRU4IyizOi3NNrIhtdL5mKvn6hlLaFz
r8LWdHSZt9V1BCN/LXbNUKqPbt5WMWUyOwsPk/aMlM2XaxFo3noN0bDekIx2l6ZuDw8Rv6OnLH2D
EC9T22D/Qmpo+V/a6+xqXVXySAuaCjsTOwlijhkpkc8v+unwnP/ekghRytFnxpnzebCbiP4h9SVt
jM9tAgws6JWJojMMMEz8sZwN6j2E82y/R4lkUfWdVC6BvMYAi2h36y+SFfL0PbsT1Ey3T21PZxoA
O4Pf5WTrfYgZwVsBo4miuCRDTsFWkbJVUwQFVqHZKZNGCXCQ+/UkfFGMmdTmbbbdzlY8EexIjerF
P/a8EP/QYDq8UEei3ZqHk2sZ+wMUfkTvT30BoyrlpTLGi1S0cGT4dvb3vB/NNE3aC5LR9V/fHzjd
jlw1qkmr/7QlOKTdFKf0c+dh+pAomaYSrwCPLH3CAqd6qaIBVnFc/SyoYDgjzasEptU0lDNp0O59
HbQRWt9OmKsQmkavBrrZw6I1PeaxtLCcPXfi9HWiujUcJyUzcJIjGNayhmMiJycfg0HQtQUSRV8l
RxlJsiUz5uA71uAmTIApGrJS8O1J5zJKxUMUO8QHpyZu0XEJW0S5P4F3ckvr+dOCNIDi72/D7KH3
F49SPxtH6FyPe/RRwMoVwLyddoHk/gmHi0vwkd6z+BWG/elwCFMYBC99H8LvouFUK7Tb2GIqQWmJ
6NrlhTMg9gtUaUkS/0n6G6JQDeM8goBhkh2UrElMDGtbDiBLo2gfw4vFckh67f2ssUjcq+nOHpiX
mAMwhRnzTwS+pg6pTzNxra+ZhuG0lbo1wTSXqxpaPFXs9h6qJZV+u+PrLKZUUe3K/9auKrh4jxey
p0o7Lbcm53x23HkZR8/FxcADLE6awv6v0HXXHrYdhmSab5q+484Bz27H41nQ1CY63LXdgOWtvsnJ
e5XBkUS290lYpx2N1CJw7zq+gcfLouea6MpJCJe2TYQpb/H+6ZZ2KXVb9C2rGuvWXDlcQyVhPdQj
y7iL66mqyg0y6IP3SEL9ysBxpaDI2rXaqFP82gBnjDFuRmalZFS9ggP+eaxea7MOakELN5WflBG5
eL1GdXsi7qyzzpwOTCKuKr1K1tOqBzGZv2vVZVwP2g7AGE+UaGOZDE9BEgDRS/g05XBg6FiltGVT
Igm04/GmV02yZH8DLZhlhssB2MIdjsiYtWXIEyJI9hddyiGFgupNvfyMtIuRAnEYPIBf7Hrwqhh4
q9NSmYAIbWlCnVv3bdInHPeTFbjTLlxT7uOXBT3bIAEtjp2W0jMSULVOfpkdBWCp2Be0Ti7g1VOF
6WGSm7gwYAkbQHPN/UXXiQ9s7ThJ5tEJ6nf7bqp/FpSVhG0ukOw7+sBtZrNnZ+SAy3VygcPfhHyi
fKGZ6DF92yCgrMTPKXkreHYweSzYzUCWAnkpulaqaA+VPIr6Xlpq+ZNapnD+zmccelep8I/5cyvv
1HTsNsTtupplLwz+tSIPMAcsuFrhe43iMh+JrIBDZPwBKmoCdi5P2057Xv7teUaPzN0HIF4hiEiO
syyxVwbg2CcE4kktMG8D+ZN9Jty+Uy5Zs7aAhRVnqj/RzYYmc/E+roVqZjprAyhJrE9dkPm4SXVX
RnPKCrxOwXC4eHb8Kb0yBTboVyxXrJspCR8QAV2WLo5Zs1CLXFWTjIalFSYcUTBXpRHpGdZ8eZP0
movOl0aNxiAVFkki0gBPBQYy7eeLbfHfK1nSeIODOEJGQ4x/jYDOkkCMkgxbB6TgI8r2xwj91MWV
e/kVEZGwQeVJq9I4K9/03JcSO4Mk1+9f/qE/X3/12blmaAcdeZx24mcdNXCgzxIOQjtSwokCkVo1
wrd/WPYwIExLQ/myp+9dK0cqn5BaH65ZVv0YZQpGCjBtQjmlCVGjiLPzPiIJdr800HVtRxjIZ1c9
0pdFe+bPIbh/RzldwIZ9+lbneItu0IyPJtrRapS+vcZPtqTXrpbZPuvWd/PoSZT8Qk+lNgRO+s0/
NBlePGuQdqV0teTGIs95YQmpGHOjXG36r8LqsMTyN4plIXG+hCuge0ZA3sl2SSsrBOkFQ4t6p0Ye
VPJYVvLa4upcSUxS3IOenmIZpMTGFKjLlSa2tY8CgdQAycvTU37ILaFDKs/MZseQ2nIGhlYqEjuc
1OY2rSkhjPcQtt1Djsr1CjLp3hNE0Yy1TSndY6UBBle9IAM7LXtLtIBgYNeZfox5W4NgueKE9rcw
Sme/Efekf8pqUb1ocTUs//uh44DWhqxwuO7n3Q2bV8qNLlfYV/gAQY0vw8GljuiGlffUTLp2/w5D
ArWBhVsqO5qAcvzTFNEZzTIr8YCxAd0Omr/WRp2KTsPYdF+f6xFvvUsLW0RmFMwOhox0PX592HyZ
bENLKWCRnQaOtwYr1w3TWFc9Oz/IWePVYH/+a8nrX6oYHxVzNFogcbXmAq+ZVu2Ri1qWBUeFvZ9i
jiFX0MJx14kQY6mu2mOjM0jgReIoKxsJB8BSm6AdBd/N3+dTFVXnxGTIvdegm9CcSjpSLGNvReew
1q+GywxR7n2YFRBnK3rMI2SC7ZxSOu188mNVxoCPjvmCQL48/zv+uI2lLjUN81BX3Khyc/W0+TqI
BbqKzDbkb4hp9H2UCgO7/43O6ZR59TJSGfW1kMgo3LQ3tAlKimL3kV5bpd4ayphNXk/7K26VaKBy
o5EbmHDp6RoYxrwbnun0ig3d3UFiYr9ekUUpqwUBgWTS3Zx8nUQGGDBw8XXESo0EPaoigQjMKId5
YmYjAjO6WpCPEBXYhnhTPHZzclpy7PC1I1iCutqA+fq6z1uInuXMyc+aslhvhLxno9t9qirZkXwu
w/nRe4g6RW5ualER2wHvuABzIEdmR0MxOrJ57yJr6faWTKk8vG2al4njpTuoAgUtxEFI622qJTcx
HFK03YzMJD1mZg60dqQ2WOuxshLuSlfbrM3Ftok3nbppCt7bLtFX2Rw7r1FrAY76cwvB+gJgnHvC
hY6F4/aL0aJaE8vyGU2pUYmU1o8coGv3x26C4TNXmgos2OiOvMMueFSnD2d65PJejZfygUH4j+Zx
ZmyUz/wQjptU9DGIk5DLktd3Q7BZYxNFyUZqBFnfTdSLSI7gmCjHByO3lW24PFXdSS23uhxPT0G3
PD9PHv43ZDJc7H2kv3J8eTJfLKNuaQDjoOYCqd5KhPa89JIjXJyMf1a+huNt5lvEPNSDul4Qfdp1
J2x20ocBJ06iLWxiiUnI74L3pf+zNhQ2Wb3+5PjWI5XOc+NEP7VcQ7/JKkZZqWV/oeA9nO6sKMts
nFsC3UJoxGHJm7Rep/lS6MoOtz1nouPm4sFZrEeB4n/cozo//FuvzbU1U360nrf3RJZ7E4AAdDdn
DAMmsi8P/MKqNFmrTu/RG+hiaDlXSTlZTJFfClfne0M3QcB2yqOLzltxoF2fNSraSblsE0GmWXyR
XWJ8635zQQevi83W4Fr/wqYsj8J4uzvLg3uTNSgpqBGR/TeIF9bA+OnloQSDFKVtHZRN8C/Ync7T
SmejDNmuLDxISrNWvnGEoD7cBjEBGBd2ZiwKibqIiywhf4onpMFCCXvSafz/fdySOHUGftiy/QW7
RsF30k9LOhOjKP99q4lBJQ8V0RAzrSXkETqQ3i34jvXsiRJ/X+qicRtWSGjhjtujUqta24pY/6q5
FaTPUpjl2/XPXtxoYSvzyC5bfzigbGIeul3sUtw6Ku4hRK+r6y/7NItzp8xAFBn94vX5WxqGzwZg
gda12j2eU3koDZOqn+F+j58+6pzlI27LrEkgxvtYltCZmMFRg8NyBquZIAylGPzzdzcYgtVAu4vV
OR/UnSdycoVbinV7Jbayyw/mTIa2vVUxWJjnwEeMmrP+dPTkDypiDxGSVMj9qKJh1dPjYjyzwrzb
kA+5IIEajcmnDHXJC6+s/pznYTdfSsx1Mg2F7AWPX2Pjn9AUVSf7YyoBCODsQM7ckxi+aCDWtGev
CcYFbuqtHSQnfDs/WUuIIE4vhAqqdBVUzUVqIeXKDuKpOSwyth+/D2RCRT7Ok6Gf0fi7WI5G8zMX
UrP0SU9+7rqsHZzrPQYOc/9wrO8n/ufPrz18FvlyqUp2ronCCTDyum4TSFgZmSeKIzonfnG9zTlv
fsvJ14alGvfA8SQXjiAjGDzG5QXMdszg7CzcoAa7zDeJ0mXv39okXeSfV7whM/z1o79Hu3OPYdTO
Hik/ibEZzSu5dmMXk1VTze5x08bhRVsZU95sdNCqo73urDd/zouDiHwDnqoedIIxdMqWwIsvl2Ba
eRyC97ML6uvvXHH0rNlQ/IVoulzAWoXaeYPo68VHVKTV0mJ5e4Spsr1R1Gq1LXbeAUlNqu0aoWHS
sRiJNZnMUerhwqBIHqRSjWkiGbMiXKouApnBtjAb8RT/FF4THGEp2+AB1vKy+Od/SgalHPQAZtNv
0QwEfk77FFbUHYj0Np+zDAEkBzW06ERQ4xvQ95e49dOKZaBDOesPOYYR4x2/ELRjO8TEI06htP21
kYljjq2cyeumOKVLicI+3CluYQ34BsWKtbhAXTXxV1QBDsPd8jtV4siHtrpHHzEBgWIWiXYa4slV
0/D11veVxkEAeRrYZZUcFnP/h+2S6ipaOMAt9ozZvWZ2SYVudkvvNKWgTWTIc2xxmkV8vthqTfVK
r6xjIVdczd3EaFzw9L8B1+xWepQobU5xLxppox8FDIrmwhoyT+LqVpMKRvBiP3liIeZ3BpXtj1Eg
ApZNT4jpviYZqXLpJjUAm+NZS60rcoH7hhKUSGJbQQGNT7Bk8GaP1I1EoZWpdOKNxQKicq3nX/VW
G7Sh5kc8AdVOCg8rtv4FHQtMVn6DbXT5SupQs0WQYK2YcBAXly8p9uGyEUIn8pCRdJp8j5vciLDz
vXCXcTDbb6ouAfu7s6hqn1YKODCSXqTIBkpLac1ex6kC/49yJ/ppFdMDnphqimeYg7Rjo+0LtrJX
RH7QPGql3TRzwnwiNWQ47e39DD7cF8EzdJLBKFc4ibRMuAoNn4klvjoTJanf8u2VrpHg1IffGN/i
7NXoqgp5NEREXjAdbfL+tyi1cBb+JWJTzbTBrzS5qr1YPazcc4vJrxQtScB02GNBUURKpCaJfqqK
kbD3VOTgOIPvOiPO6haE2phdfq22Pnzy44HeOGPzVRCe7kW0zmMZJu1IJACg/D2T5HxlS4yuESDx
p1Q0GPrM2RdB2vc4shDskbKw7dSiUtoEa+QJcaB2Um+3cV4TB8xwyW1DWSSWWveQG28BD0NGlAkG
Lo5oDGy44TYoeoQs/uF0ERlghEQzgyhGVuST7e7mpelRECFeRqXDmZRb+IU2EfOizxSXnOQnjTvz
tpqgNRDBqX64nfFWFZ7wNACH82qLwansP+7qRZlSur2FNEG+u3M6AZBB4LaZa/MPdAU4yXZ5N4HG
G0xKIfofRzErJHAQFplgILSxt0HAXcevClDAUX2f+kP2MvR9MAAQ/x+2EZXvCv26bgbQuLSO0qwx
S1w5GyVYKvFztNQj8/522Qs+U0prPNsnXX2rPCBA1TElK5hgacofKM7jzVpH9e5WuD55sU3/kQpg
JbiJGF1u9b3IIQd3qTZz9D02UUJ4Bs0/IZG04V8WWP/vM4wVX0oQ0AelT2idGtyg6umFYrLUPH8n
CIY1UO2KBzGQoZLSmPkN/sbAPu9QBmk5sLpVowcHmJpBxyvzP3LOGkGYJ81Wx/0d/2y0mawlMlrV
OZF98AcGFq2vq4QmIfTMPSaJuRzndl+ZIrKGEGjt4vY6Vck1jyQQt87N6PPgDOXobm2lWzdwcMX0
m4w4IhoB6RQKrNGBgc7FyC5QGZrIW6nqZ8bP4kRE7SNx44CXsryQb0ewgLmd9B71CTWpYxHIhoUm
CMEIs5eQubbmKhZ8+TMYhNk0c8JWfMoWPjlgH4v4XybDhn3dnRJSt1Y6dxs2R3PQHRlwukvgCuu6
EWmRIBT5DzFlR33lIwUKC4/zjA73xTqSkp27PidCPK2IrhDlNwvj/a0qsWb2PLBbLmG8Fio4Hcm6
glfupQhIMWQB37d7cnzOT3NcLIkdywuOQj6jMICsa5xxYv6/a2wH1Mn5ZfZzS8sU1OsENJPd94Q+
gva15j49TG18GqKwYBsRBhLYKLeOmtaw2fI8jY2hJP605Bb0LJVjkfc0ujDQg4BsL6+2o+YTvqYM
3d06fGDlJLPNOTc0/Bg831UWahjyNZboRVTeEwZwhK002Rl0F0J5pt8yFSCsyugAxSF6r1Wm1ydh
4qM/Cl0BIfPXwwNXetjJTsVWBYoxGxtkRDYC1xz2HAzFnpSb1oIQgnErsfeKGRkUwIRPhRZsbyln
mL1S7jd/tBwdAnWmALOkA/Apute0ZktFrsJMVV3i1rIFI90usvrCWmQGngCGQj9VZTwRCzZzc2Dg
CPffn7bQkzwloVzGxrUA1Fuohv04qrVCcih162wYk0drWrIHpdDMP/fY2V97C/yNIYNxmMWRzy+j
Me5/RoEU7IdvIri7dmONKcjb8iFgYry5WZpoO/9MP6mYzmpu49zc6WKA7bA4nQHnIEcpeQyyvl82
Dgs5KaEKUie5xIxXNV4gFN8uVLoXPCDUob5ZVQer6yz5oryzYZ/7eEUPccR2qvvc73WQWlbpXXdb
gGvemRKUPWXggZ+QCHfuVl0K8jF0ZxzY2ns4DWh4VvkEg3JOVkFsflC7fGrSsAbE1Mqemi597KEa
wpKncoPwy9sTEM1FGR8b8Y+jY21mGRIMRHIaeR7Qt4TtUtdZrFZn0HjSeNzCukICOZuX/PphNFCr
gJjmDqA4jxweStWaTQl2duLozsyG2aw83OHfkuac2dVfpVZ0h4LdnV3UkGBp1nRaK/3PXG2Q2ISZ
ODpUIVBJe3v8DKwFOqsI4XzppbL0E9OoZZe+Otoo0vYh/PcqFDuRTvXAZo3+VxlpPM6hk7F/ShAH
9XhG2/TgPyiPYlZAV2XDx/1X+1d5CNutVV/VTq3R+pF9w3Q+buVuYIeQa0QGVvpY/cXeoA+A72o8
C00Fr3tTtvPJEz4wcoxfv41bym6/+DpHUzEShKTYoAHwvl3fXIe8HMh+VomuGkNUBZbvl6gZECZG
j+PUzg9odWajAyu2xj+J4tFqhRzxsnP9/XVpIQYRCu2BMtnohmt/k0HC+f8gDF0BFW8VmNiuHcIh
hY9WFNH+EqkVn0Wf31ThfQvYwJDr18oTDwaO93RFMm27XpAsy9S1byuUr2hWQXTKGiTXsyNhVzAJ
Nlr2mxY86OwggAExZyeJI5DGQDINAq3qv+LB55UXrmeQnf4trZbzmdRPRQj2yEB4bug38ovcfiST
Lj/1TpK8/83sQ+z5Gqx+HupEnrCgpHggqD3BJuivCcK2CNqtiXpRCY8MfOf+QGhqXfviBBx/ETDD
CiK31uJUrVT22fKsRf60KsYSNxMJbG5YhnrK/g688tHo3SbQKd87jQrncn1JCs635rkz8dCE1L/h
vzBg8s6C2V1IIQ8n7kWPWKG39oWKblUSMWTHPquXB6cGdcWKWuKg5B46FVrGVsqGZVcLtwwpIG8u
DL2YRqQonus0RrSNHjp0uZcDb/bvEop+j03HFun/VnA39/gvL5l6qyUsMQcJJLe98q3jTlinUu6d
hchTMj0GuL4i8EZeUHc48HvSJJCbTuuzZWrawssgWd1XCjYB9gzUGxlsFQfjighELUQM1sy6TE9p
e1vnt3Vgg4FObOcwUiqW93hZEe4UKvgeztJKpXanXcH53RkIlQlyxRKyzIQCv2E4FQF+MALHJr/N
4nCWRVaGrSNNx+OCTbnLlC3mkpjzR812biYG4x+0OvJfEZSNRRuSNFLa/+AXPtlUd9457s9ZtV1d
OnyBs7CWP/5mXT4t3rrz2NgR7U97lpKW2ymfuyBiX9enzm97UzYOZZGzQtboCP8JJ23l8N765C/C
AdAR3vywniKko1T0Igi8qPYMyBGEG8T3hh/ncLD1owoaZE6wu1Hv4TOmlY/kAW8Rhxjq2vyW2LGu
o3JsB+RNWk96wFBCVY3hMsoaQkmW9MSEHUxxvJlZCKNvihCTeksN7v5WqFLlnvqLlaBejCRKztcu
JE+MktISaRcKxbuDEyt08BiHRl6fMohkTHwJlP2SYFqIT2uudFWBhCVtdGfAmi/jY5MVvkXYajkX
C8+5I+msQtIS/mDvrlMAFYk15GdoO3BNHZAIKPeKoYFkJZPS20qIXZg0gcefvYIIJdsGJPQCdL7K
XlZDJ7gPrJ3/Y/9Qvd0ci257XdjP4tQUYaui7VHmn/4A6yUO5l7ElsHUd9M8a/pk1iBdpFLEZgr/
hpc5S5C4PlgsOwTVNqa68eoAPgY/xGxXzNvlqbPmnNdlidE0ErXasIvs6lLaBuGbIDaiG5Fo+LBO
v6fmj65hTOTDtQ2TlutupriOy8KS1z913N+PNKAqICdwJueqE0/7d6rCJ1AiLqsjHFkuM63Tu6mi
sFQuvhjz/4GnxXu2jxdIroYXsZTDpgA9MQErF0QNsLs6Mj1ynrqBYoPkRTijAYaJWjowRZGEiDwl
FCTXwXD2kBJ5BjZZXykHcETF8VD3e4sHC/0qA81PMq4lcHZgeKXE8BH43sEQlOoszceYL5iZxjy0
MpTBlLifEb9jyHV5ioMJNNPl1nIYEhSUe6cHzW5FuGiI9j4b//TFZsviC5MXx9OI/fOsnAhesvPE
I90YU6WrJl8G1hiAc8446OxooKt47+DxmB5CNqLLuooOlJH/jIoTky0QD6IJmLNcrwIkZkIvctwh
x9ZaFUXCoP2pnphYke82zIsdNhuPEiOaI9asQGFyhzyb+tY6+FcP6RzC/PFWmH0mjmAiZoamjXgV
k5MYQ1UWbQKPcYMlhCqczusz2dsQMMdzHKH/lsBfO+TfDJhWMLpUbezruRg9WMbWbyufOVpXRpVP
TbHJiPzcfYfFT1uVw8At7NovOY0Ril06DL2Eyl2ttuQyOGke0jwQza6MKYSoNW4NdtrPLZI7XaLm
ILhmWxAtUyuSBLOP4tBjtC0FE2dWLk3uqP1kHM6Sxw9Yo8aXyAzEFDmPUaX9fNRhkabBPHmKutYx
3W9Iqt+oegEJYDnB3ocUwGZARE58x4PDBglYt+QDig5u944akOfQUNnstQ5tlhpbsbzBanQIHZlm
TyifCrb0AMIldV6QsdUVUmaDXn02FAWQYm3jBsoE5lrA35vhFfLuLQ1ztxjDCM40AEYcgStYQPOu
cWQ74bvi6prqOJEwVQJiX41KaSSEFcf85RCVF70ugCDL8Snidh+shmiJqu/rS/ym11ulZ+d87sHo
FktODCWJtCWys1jrtDoVpixrLXCE8Z3C7bh4ZTtDRI5KJ/Qafv2tLzNzxsEYEpdJALwHzrTgJA8O
nZj/4tDvn++2bc3TG9RDSMBgSU+x3oW973qlVdK2iPWSIyKpOUqDF8PdFQtr70+JrbS63QrxEMGR
1Om4WBnAiqPL83aT/hVw2jn9yzhTq9Hs5ouMCuOwTcbOOV0E3kzTGfsuyXknTJwvYNW63I+Oj0Qu
WK/LcUWYE6/uAA1lpKquBPqzLbcIlcl/7buvKQqnqdgrnQw1EYP+9C+IGzgPLulakhDf4LHUKiVt
9OcvNiOxCvC1GfUQAEt1HjR9I6KJVmL+LPESiopwnAq7PDinboWIN5qJLEkhNhbQiFR0dXzx3d0X
Eki0Y62Kn/eX1GE0YzqmMVfFGnZHlVdntZ3Vo2DEd6RGtCkAsEmU3spD/vQJpJ7PqAT1izpqYvge
NnnjKdcP+lgsibGqy6SSrhNm8ZVG6oRKLGFTAJm4Zhcj+wKfZTvrOc4lx1b/G3qhaGDs0z/6JKPN
MM4Fm/ktktp8BbeOClyzoBwnJ4L1rR+K0BHBw+mQ7TUwdtJ+8akEIOc4EBSgjDBovb+W1XSsecPD
hbHGhqMkrZrUyZB2asyLNI+h1NueElvP0mzBtQjPd91vOlHlfVTgatPZaEGNNCT/RgJknUuecBpE
g7YZ82unSeHxfas9/MYtmzWd5lopvClCIX7Hf6dN2Rp6OA6py2XJfIkqXHKuCK64wGqYou8kHcAW
ovrTeYQ4khCyXT+0NyqRD0IXD5ptTZ4Baa1U5PBv2N+byIkreJ7FhV7C8A3RPGilKqV6hnwCxuw0
hBM9FwF1ZNpeFeLGes2WsmgKv+Yr5A+GPpXgpUdC/D0BAnG5c0iJAtLNDRTTpsR7usWXgCjZ5ZI7
UhZ5GHVl3XNepSQkW6fiQQZLPM+8Y9EzQZlQeSbfUtmddhRjE0obNdRLlm7Ye7iGm92hEbe6+2XF
GFJYWfeo0q6GfZGrqWbVW7W1WFe5e1SBs6dK2/esi8iZilbzppSyE1xp2n0IDFGV3ewBZRf0sGbL
7XATpnmrfWXNCS/KjkR/lLNS1eV++dvXD514cDxVHVv1Qv3s0//ze23pwChU4NymHLwhCHcIhvqp
KqeXEqv7Z5Di+YAZJvQlKjeSbud+yWnG0DjfnGNGOKNtekAV2kVTS2UcQO1OaP7ZdgVrZ9M5sujW
86uckq3ehQ76W3GPxiOimUiIop/XSUhO9k3ufe+TCNUOZ/QxkYIy6eO6fJFve4quA+8J1csO/mR/
dxS3KRmpADlBbD8a8fFwqRmlwr0/eaPZ2znR2lH9MrFPVoOSuGTcICxwrth05i2PDhBbg1mdR3sm
FgC+iRLJFGWJtUtb4HMTva1QyUGb8Vhhzu7jff69F7rD/sbH85Ts4d4doKNtGZUFOYs0XBCW6ONn
p/1t8YI3CASU9vl5vUa1l4CeEBR68jpKloCHgDwxwZyQexkQC/VNvhHRPpi6Mn9k9a2FlhDFEM5a
10N0znMFzNicsVBMa/Lj70CPH2cjUY19AhykZbkQHcTvcvlxVBqRGVTWf/w80gCaUVof/zWqsjt9
wpmSuM5CJK3ZF1XfSe/isKt9O0jBbAHW3N3T6YHeRC+YCIr6hrpjX7iD+Riog85TQj5UGbOAkJMF
yxktKgSsicY5IuwJIQv0glhm2aWCG3U0AzyiyO+dukvX8OJuTAReDQYOrtYxdDzKOEwGvu99DLZw
5ykXS4UTTNA9oe8HMIRGpsFX+mQPz3pFPMUcY2vHXeR27rdqx5La8gg2ptyHL1D3qtNXoFvp443/
f+K3xne9rQDGlA+gkSWD1MvfrRumL/A7q6/+jz4Yr4R28jzu+iWgGjS0rPzNBNskWO3DhGlQWRKA
YI3jagsrGatQeF3gjmI/dFYJw8y6u2upIAiRoGGwg4yedYM+KiOkGyjT2TWhF6W/OJYIA2MVhMrm
FOZYjfauBMINY+GGH1SQpOP6jKWwE2c38XGiIrmjXmYvYb5xlV5d9uWGRYM+VfdPujh1XLBzMwgG
miS3ylbvUW2T+HCeSKZ8XexFiE3mh7wPU7Hg6LimQ/jD97dSP9hEjqBKPehqM183TLUN5j1G3gTd
7RpPx63SZwsOwbgE55vjr6qlfLOzNOIgi8ulX3xzc1r0bl0GVHutTUFcbxf6XwCXBr+bU1crJCFb
clJQAUa9X3yf54cCJY+eIA/dHglhYBuo1W9hvNnpiWXv3eo5pa/aoW6zBu98GlbBL2Dz8VJR6fQz
qfIhdG+Z2QH76MduKjwVt99imKecpCoonoOzeJa+9UIf89MsMIztONqj2vJb6AHRp9/WhKez0QH/
H8+GaGmA+Q2XBJ0vx8iJLAs6o4C0ctd6K9QgsJHWpPIQc3W236SA77nf5v973twvUDHvvMec49F2
6o4PHRfO+hrfW5v/9AuQMGx4JRtK3L0mnJdTv1Yc44S8ITPFJJ+5humoEBNFWcBgxTP9Gzt4UJjD
lH8ZdPFrcmVPIcWs+Vpy1hfSjjp9FJe8ykarP3TDSva47O14wt6SiVPZSSyob2zdhkiJYyiRDNIE
32cqy0sRQyzQxu72sMdmWKfeJW1ohgfshuPMG6KRoLftAdh+BAi6/VK0SJNyzWR/r3sZCam7YOVC
zw1qJsTvoFf3d3vb1zpC/KlHv2f422/x+t6tAWbqORv4fFYGULuBI3W2kK7QcPD5+Epnw2n8u7bH
582Psv9boswOOvjZqntnJlSImYhpV4clarwUJvPJW7OoDSlV/c1gH6pXBce1ZPEy2I2tNmCby9af
JIQIBwSt/B7ETvvTlWLlfu/SX7D+qO1diJ2U3KnV/RXzwpWEbA2+o6FrprR9PXuiJWyRQ2Vfgee2
6rYU4Izbg8QCJSgmY77I6eWVHLuRP5py14d3eMKO2PVO9jOjAxm6nZkXVU6b3WWoPSZ09SOY4OVI
Gef/0XUHM1jVw/3zCZYeVGo/9S4Hx1cpx4J4WDTJg44JrhLMIpFTZ+kfk54sLm/nFA6dcbQsuPjh
l19GdEqb8+dxSv3HpTPD+hTRR1SGwHgWdtNgRfK6oH762j9IGeke9Tsymc5xl70qT/QK9UrIYanI
jPjbNKnEOs8LkSkb4vZ0kt4YARGkcUwvDh/2vrkMs1CIb7tETA/0UH59u72SunjiFQbI1RN7KVWt
jIf2pshlHwNARZ5sPs0YhmNYMXvFg23VCiJn/Aq2kI06VQgYwo0VHSSqBZqXgWizxxB4S98mHpJy
RboG6r47Tg+E5UunImcReUmIexWwA977S6deLwD2N8gfyTrlXL/AUxKdcklfTAiYpvmvWN8WDOKj
ZQRVOCmuaFS2dShzkdb1CK6nlXPmsYygPP/Pdqa14AkrPgwwk1JMZMD2anMCfoINRzIhWD02eCfD
Cc9vxCloldWCQPLNBkVHjMGd4MLUE62w8NF81IhkoXWkjJse/yDekZZUQBnNurJlWWQpdVkY5ubP
8bpVvmM6JyYRV8H3vUii0cEvTO89Mvj89yzMU6d57+L37TkVod9LexWvdxq0t0v9pMnhVilWiWqV
VCzpZVsDpj59GhsPd0TuEtubNNPjRS/xjQHhZ7N4BiuLyuQWK/oJpK4PV8Xf9ajjViKs5v+st1IY
UgUVarCZI4nIJWiNleeAuBZaxi9er5qdKLqtv2zyj/rHLeMaLQVC8m80KwKBnemG053dv75gAINe
0doofoN16n1t4pqJIwYomMpCoN86xzs7A+ycks20EralTsgwXSpAXKL6wyWJEg4SSk7k3iZ5BM2C
qGEnO375A8UG4Vh79mj+PRkRgu2ON5K83B0JWz5jn/KaLRru0o6bOIM5axK6vORqO9oY1YhrEaVb
FSDxCOW1F1q66Yi4U/GdVuFBkKlXwpRp/atD/oBE7m1XRzLv92GHJBoTE9IT4TYIDnHjgSAqsRLZ
KCtoP+Cuvfxy9RIYmZyXoBupkbgYMSGLAZg70kMM3lpkabsbgG1n57oaMIWfxiehSMO6Ac6hxpTj
zpKFEgFLZupBJppWrNn2So4vMCuu6VW0Qnm+G7n1TGHmwfKo2sGCp7Nj3Jvfd+AuRLuoffL2/eT9
Kh4n1s8WAtS3skOeaM+NuSOvwRR9Yld/NkJttzc5P4K6KKKZuzrKr4CxIuANTcMXWyHuf3GUmkGA
Y2/Fahv53rk/wTt6gzg1ep3PpsuwqFNWFo2ZMAl8g8JdlXjv5xQfZIb9DG2aSZP+YBZtFM+i9lvr
VRCryztK8CqFr9hmSC9mZJ+7t8aY3DwL30xTE9sYdpNgNkD2eL98WdSE/S5lNJ+dNy2z0+VK7zZa
bmaZIkOqy+qVQ0F9utdp0HWnXpIgI80N6ZA89PkF/U5sxy7WMvYblPh6ljLZ4WXJ/WQa8DnBhuO5
psOm6eNaBIvYrQcgtPNvyRWgtuqludo86ASD1pFLQIz33H0Y4BZPiGBlqxpiFkIc8bsjduBeaxfL
oTxmhs60M7pgIdovy+udvMF9bAUJbbsATW1nbm+WCWeAQ1d87lpjZvNSkWOO7f87ESfEi3o7JRL1
/o6EKMdOtMiz51KFprUeeiCsE2YduZjS2Xv9KbkZ8DwJ/JrnZstnbtVuOErRuAWJdO/UbDg0L14a
CegBVbxAx9xWZMTfZmWb9Fiju8pjCGqt4THUvmgRCINRyiH9JbCw/UuSkGRPVonFHIVMxSgXnXFf
VEXpttugO6x8VG2CXBPrJzTLBtMdzle22VKCQCS1jawSyxPTE/gYidF5tZAZdCqT8JtvMESnz+IN
rElRPkCrfAUfr5AtKVQ8wB9nBPn/ZOczKtyXqL+2FZjm2zMPBBfjfPww3Ffsz9U1qn+CDCAx6lUW
M2X2KR4C08Mc3SqTjptELeNcWcGEbXoUZK5yXSAlolILDFMg6hcKn7fsSJk5CUOQamd9tv2/H4u5
0x0ejdWZV60g/Vl/HDrT+mA73Y7sSiNK+NMbDebOnZRBHdLDFJFHhUKCnXAks/GgsOhui+D8Yy8/
P7OD180zY/L6vboyaYcrNes9Lx3ABa5KlYTL6lqNXa0gTFyP3OXZNsButiuyi4XyzhDzsg0+pKdg
TdCNKFyQyxP5r1lwab9rxkmjDGrbKQ0R1iPbibXAiQmTtNSrPMkdrYvwykBGN8AR6k8mDdDCOq1I
pO38or8fHzzcYIZ+vM249Hfs68uoZ2RlofHcmQtrJMog88d6/mMtKvgMaMIEJf4tLzQnZTeJsR21
gQ8ED/4GLwXUo8bDscHph5sIzqzZPMFNXMmWGTNqhvBvIeR3dvg6IRvB64jDHzkUx2SCS4KT257A
C0pLoH2imvJbN5yPDw0zgFqhVB4tv34CI5bZ9V35m7osiTJyrZT36toCLJrkggWikRqb1wWdHB6X
prg7JT+7QKj+0yhSAWgw6xLpSh3stenxq7/uOrJXKnBGZLUO/srRbkc0gfUppQrNBzs73G+byDdu
q31L88UYJtU/6t60nONaMLV5spQhyn9DvnlCIYp+xTiwfVpQ9GIBHuuBCEZp/81eOqdFRV20i4On
YgzG0g6B0+ryFV28A/+J44naNkoLAB/ZWAFWkRE5w3nL9Fwwjnbj++4kaB9ye2pGygGKfW13eOa4
2wcUWzj0zsdzVKZxsxTCNr+VmYq86/rCHcUC7Z/HsFK1JHcxhaaDOzGF1NPTUipOzQdDzvHf++D/
y9S5vZPoUV2rCwgPm9kcQiPgyiBEcviFwnivPNlxhmHoi6r4WIWHoIyBtqqBc5jONB1u/WwQ6TcA
jRP6llsQrO5ldH2qekKASYcDbh7LgSP6jo6baXcGfrmDCgOoYfxsznh9qCywssqRkFHQZWXN0Lah
+tB6FzhnYFWbewGBkc8TW1dKdF9MnzOhOox8vRydFNuxlGiQPeYcgeXwDLg7UpUxk33My3D0qVUA
toV5jypKrT9xi6jPNpCRLGD16T26M6nAdAqKRALpWHELFujxzC50Gyo6Bg/b3HKuSCa0/QHoMFlF
R3vindhnB85JFTyV+BMdE+LSRDw33jtkRckQZIQP9R+FBOiZKtb8YtL1Vtc1WuYWSLhuDKCOn/Tg
kh8XcjY/MkHNNINyLnibMREKxgv6JWc6ZUmlTU261wraV0TuJ6riKEmCLo+2Uswa0Sg++6myQefD
uPTHK0uTMSybTHfFtYTX89VA4R3HDwb6dnve5vpmwdOW/OAbUn0gYL0HWzKVlgOaco9b0nIMGHns
eLBCebOOCX397Omu9TCu5D+5WiTNe4tbYN+J05Z0qwS4eDsKYUc0z5v049Fm730ChOn9lXz0+SOF
SFwYpfFY5Cnhb0qS00CN4F7ELpgBG3AYcMbkUGUxdLHdNOXzm5Bary8ckaeYghpR1+FyggGpqJYR
jPIPAlm6Lib+W3YqTdxlq31EkG4ATD3L2yLzX7QUbQQtQAxirViDTqT1tLxz4qeC2nz89ufBPXNt
WlaTcmHdZ9oQ4SI02pT3oLksp2DEX+e8Sukx2gP03mCKtNcIngCXrmmvF74DHqw7P0iBRDhtGunP
ede91+mU+lva7hp0JDuy+oqZVCLgXJY+WsdpC/5zRWlERfqgSEHkuLBfR62Fvz3WjHNnsQUGzfa0
w4/p/PtXNsmZD7LcmMGHyZBXBVrtOsLSgYF9+qeU3B39sQJLsGdSwZQ5Z2IFtddjs9hzn5dgKgzK
uvS/nhZaJwSn8b9wlUFvD0qVdHnh7CIK++VIlhfShHXuukG93GldI6iW1GSCudYyVWskhXludmKC
AyIL9pbJwz0hG7gEkVY+VfF5GpDOwvHSMxHLJN7n8W6lh0A7jxDc0GexOwY3npftsVAoV3kHcWu9
DK84jthp4vIV7DzI8uXgw6vxUuz3POP02t/seK4haUQV3bEKPYHjpgIyKPFW171zsgTWLTeDh/+9
K5fKVhcS1k2xBsr/LcSeF9J3MysCwvaHA1bNr6fplwMX6FSzMhiU/fxFz7u/na12jS21IZETOpHm
4+Ica7jmSvPVf/LGFJ9GYEg+msE6VvfvvUGNeY27EfbLz69vd4jC2clO5yGbVNI787b3y8Pfpkv0
XG0K5RfPXdsDoZRMzbpugc1/3j26xHLrLskrWD1ga0i9tJEbz/tP9CS+LC47SBkwv2LvnE5puwuh
deHDAM14y6DbL008/Ulpq1Sbt3b7t9pSjOD0ydhHQ3c+7WKFfFsyEIoH3HWz/4rKBbc3rOrTLlHx
LH4NM3WrSxcfGuZJmmTiNv33X4uL4MX8+WGOU6/8H8yYPHIXIbtgfU4Kvvos7ZYEBhkdcQXJgDdt
iyqomK4G79wSNWCZDzNh9jRp8gJDqykQA9A8Ljwqov+TMJWj4IEQd6VFz/I1dfc/F3hAwao6kKJZ
yE3+SF/3VJRjBtc9AGg1fcUPwIFa27TBmyBEecfCAaUBq5hvsI58pbJQYDUzHb2eXV35+m/Zd5do
1tWkveHpX1kW3uuwYWd0dSt5TGOsyNYgtWdYv+c5tPEuNC9P7oCzM2GhVXsfPl+UhwlYpXCnbwyp
wgRRgR1h62St8E339Pz7nJo/kSuaheCHra8gUOhiLK7Ey7irOF66egJVzWpsekq4vWwU/Kz+Gn8K
ihGkbJ91GUzdzxCqPzSvDwLeU5VWjnNABKobwpRsL7YgKmCulY+xwteZVDtKXctWzi22asBc8Gry
49AUl0ywHUYWFYNWJs7TE3MBSMSn9NYspBSymsdD9qbxVZjBtYS1a0AGPt6y0lYbPuTSeyZusnfs
JOM8+/if0/zyb+tAeWgID7o7HEgwPs5MT9sAsEES/IW4o+/dd7yeta8ifZ76m61JqulZc/fgG+Gs
E4+bFJ3ZtXGDej4wPLuSCbHafb2Qk2nia87C6opg9OxnVFwcyj1Rh4YpqZzk56Uzwa7C4TXjPi0P
27he37hOmxYUTM0RLAvboVlF+LwvpKligJACpIcUYKOV4E95gUUdwtfgND8dPQG0S6G2VMtTwhwp
GfkUuEZzAP+NsNj57NZIxq1TXOcmHL76YO5fqd+xkxTYvmx1GdJOmnAbWbgyylyUjk5y6owAjQeb
nnbNgcldOrgV9gqqC//z0iNQLNCd36akFxLrkONDpuKOmmdHaelv2oxXY3Vn0Px1u4mwcRlF+G6V
St+iKtGcs213F+4i3goP5+Pex2amPcjEw6pP7eAGNN0au4JTyw9xo9iDNobc7gp7YJCJI9KNsCIi
dVTIDdlNrqMKW0bVhJCwV2GVEkIUFrelBqPu0iJMKaLOE5rgnzzjdnmzUGsc/7isTL5F2Wk4RiNl
AJeBPDnF8lQIPlP1+ZRe+bvMTWffz+oxdqhO8F1ZaFifScqB0AexYQYOGuCXadrW6Z7M6rnCwfEM
XbsEpodEQwsou9RpNtnG+pajLmiZO90/a1YJmCbNXuRXYQHhG1mzfR6joRt4WtVs67vklE4Ud38i
P+061JAPyRovlIEU/4Fk1y0DXk8YUpkX1/r2HvCE4U/PP12K1Ac3JUPojHMTLMCiF3t4s2UfEl5c
DTtyvMoUKAakuLQbRTWVsISujbhf0WPt/zfU8K0QoxIKep4i40CjoQnQgXsIJuhAfncyVaO7wdMO
4K4rYku36WsI3EF0I2PZjOpP4hwo1VuWdkzPzX0vIJEFuhcew66YR4h1S89vgRr5Gx3syPzbAy/1
N++4v2qVdFYhavx20PqnxC2bg+KwGHDXcbuAoP8u0ttcx0QABNXu3ZyQT5E3IW4UtvpWIazEyqhS
7yfhnGX08cXs7Ghms8UofW/R65jomVnninuSLFoSvHm4DEMN+B3i2xAbqp8BIaqIuJhWFgNWMsgm
/8G09KH7xb5rjJKSRov7X6giHKIF+00XtmJwRAC7VBmT3Eun54AIp1KLOTCh+RandnrGoYD9sKaO
UWzCkPUF6VgpvtozpI23C0wvF40y7n7uLZLUE96PSe82CTPf+lHkNmcqQvHfHgU83pjtVemqiCJT
Tb33BhHMBmGjQBgkeyOAFoZZadFHgk3jSeGal047JHIju7LN9297ra+0/hPgqZIux05QRC7G0vMd
AWTG9vuUloccA4ebMUgAGLDZnnbq6xP0uCQPhheha1JZNaCruepjI4IL+zglTYitR2rbR1F6yz5p
5IgLvmkgrmIJIxckVH/jY6j+1N5GhdxrT059wa7NA87wRId5F8M5dEJK2gLIwMc3LW4KHyJ8SEOb
2qbxF5KtpjUvCGv5owhjmAitnDQtiYJoanwudgwwcKzgaJl0BgT4fLEvI1qMXzoGJxyhZAPLn3Aa
HBJgeQBg5C09pQ+51pwXK2O/F8ietQXhcNmeovuj9PQGKED4Ziluh+Dxl+1k7zaV6grpIH5DZbjf
NOaA8aveHYzCxIofyYUQPsfZhX9ZkCKeY/yMAQ6nQKq7YSmYr8VBD21ObTx6t8QcBTNyEBNkUzkm
ERgpbyWxUFS/AU0XO8BdxQsEJ/7ps9pu1R+ilvD11Viyn9Uu0cXDOkREq35TWErmaoUZ2WT6JL9N
eqCvAP+6QkAYFhcYkrgJXrkXRQ64az98KwY1uC05uv8y3MW5ZNO47Nc837wOsitvtMlO+00FOjdK
k0L5gkH7kKteMAvmEzT9BD75E1+bnpEcTp6gAKrC+vMsVP74eH7Cp0h8PtYFLP1VZna37cmNjNUQ
FHa/otANB9Vgyt7ltayFVD6K0LoXY3Wn2Ej3F2KGXM00KU/LthRATztXUaPJ6XlVAt9FWDZ3lwue
BUoVUiOIqGJlnrRxq8nc2RgRrkN6qHo09IPsEZy03JGhqQ1m8OzJmR0Y9aozP2QYyNN2hhoQ19bm
2l7or3fYMeRF8pGkwTLwJdVeaLZCC+wHW8iyb6UO4jhRTxKPyjIx/g1UnIMFcIN/vWIdCyhDjoIS
CKvrTnxlslS40n6VPtUAsxyT7ckVs4MYXno77Pg5h2eQMTCxaFbrjJ3H3kfRb1G0pDOhvF/xvTRY
vKeXEtnq/N8FP3Ys72l0bdW0grSL/NDTFVY5V9g5yILj/hzHHJ7s6tnW7WVj/rxxnEZZGLGsfv2Q
ZnJdl02KK87/gfn7sSZC77QTdFPAKK7hWgIQ2conGO/oObqtDDliSCM4RL5TVqWS3g7WsWd7Lksx
rngVqxB9lvMc5xFnqG9Psv83OHrlWO9nM5bbnKLGperVYrrBmriK0PyBNE32P33PxbyJBPc3RN61
w5UoYKBLDSKltzSGjnBNKhMc/9ySdJ7eW86Q0lBjoWJ18DBpeMCz/JaDeM2mE4cDPQ5attlejI6+
TKg2IKjpMUqK45VYxR4t8Gomy7MpI3BOvyBXWg5TF19Pxj2AYuV4M3IDDVOxq5n3r3TtDjpcnL8Q
J+FyeHpdN9SlzA1YIH0OBNAoH1K890KGIZ4EtM21JvYrd4A1I7FY+1lLk1dB7QpYyQxw6VHLbQxk
YLcKjbv8YwEKPUHoLqiGtSFMm7chmV/c5otw/CjmX+sMZW070Z5hcVPilgdo8LvFYkiBDKZMsAGR
qOfbkuo9mg2ZI1nOa2rq9ZirpLtBJykQobvC1uMA4FsWPLvrlrZsTXn+HmJUmDcipnzRVXURg+gp
n044cYRlN9JNQYbKkYO4cuFPMI+04CYdKXlFsS44p0a4GGQAnbGBulWt/w3vbwzTnaKVnyvSUpdP
+NFt5SFK74KgGy3mIPdyzom42ljnmgkSDjuqdl+aiS2aDDSj05oS6KIoN3X7gZimkcauAPXMC8f/
zXMiird4PztjfJbyr6ZkqDx+M8h/OuI+G8zlad2CIWYhamw1fzYSpfeDSgmJ7oW22pevr8wysVDZ
UX5sPznDhzD98OCXJ9npFCyl0Y7+SJGnl3Ib+dI5Y4egNZz2eYGrIgtohmZGPaPqxgd1wmyUuJ0D
RLQEWeei8AiB0vdKURxbOyyJ21xF9BFk4n1RtikJitYaRmzkFG9ZXGCt/6t5hdPwgxCTILU0AQjj
bwf16Nwldn8kfq7r60VuTtx1DYbx8F5GYj5onBJzY44qkYNmHVAaHsgF5ugQ1H66ZVsXRrMv6J+Q
MVOIwNTL0RSisv/a0gj6I8h1QKNR0jOX2MYwaKCL83dBidubJAWm/B16zbMKOAJSRIpF6J1Kdvuy
pdSKS8/p5rYV2nxE4CCKTT+AiuxRxtbxVj+7FFX/S3kFeQm1G5vgyyAtpzBtkDvZjfhYD70ScM31
NANUPfuPn235xhBXZUDt466xi0kVtnbyqN8r+87kA/Zper2qXbN/VQMBRZ0b/SCTHZNzZ+ng42kt
ddoqp+2lfSQ4GWE6lStMOAWmIUo33gms+lGsX3mPKWqVCSnA4SWVeEKVNlh7VWk8A64E7dgYxc5H
xDBuAnUp+WCQ6O83Wz8iiajoJGGhtSlo/7L7meEkpl5prjdWEvL5PLxguxBUVWHmHapC79o3bERs
/pCea2j3g1yNMMBzsHrVvrKdJYgrX+aUxIyfTA9YoPlBA9aAp11rJrAEXDe9OKjPJCwADdsYTJm4
1hl50OxsjyLNpxfgiSuigeGVc661jR2HAFUigauMyVL8tYSeQQ0AmoAzHDoPaSeCSFm+doI5GovL
4iYeGDkQ/BYiI9HUKBHsyXsZgmU8Z20rlN86OyaKDg3WFvisQeCsFOmcisjEuFomNFIH387kAJLC
w/1T5fgUDFxOi09B+cb/YFoSi1HaFSY7YvZ8RB/y2jlfFeevUQ3gLd0LjMlYOuuskOhNRGmwskog
MaR+LwNzUZGhty8BQ3nn/rsg0u1XWnYHwSKecd4Y1Iq69SzGatohsQaLcN/b1gRB+hqDYbCxb9ju
+7A7MUFFS41Y+UYe0fBzPDLtd4tu4rDeAGzaKNvbZeoKiyPVXjN+Dt/neWc7b3/0NMY1fciaNtqI
aTPhzAxrGCeGTSEAYaivsidW5/jtOThFfYuySnUhnyCA5JwDTbf1b9pgCbLSYrLJfVny8+hjvQ05
NP3fNYUaR/9r5/1FtpQt7Ci8ets4MoH6d9DtOs6XrHlgiNHGQe7N+jSM3j4Tf1UoVDi52GXB1iJj
SdyD03qgiCmTZFi1lElSac1vF0WhE49c0/zE6jQrq2IWc/VeE00E5ZrB1ClOZNPVaRHju5ZvbASC
QtBcOzwrXcftL9Ao5HPfnEjmacppDMRnAaTnmbKdZVWjbu6XwTapeoiM4HILFQeKoiH7fIWYzs/t
0X56ONfLsVn4/vYpwXJUilt55LKlu+0XNa6iNHeEJzj3A+3tRMC9rUWCVNkWzR50TIZcRqExHkdR
nC2/au3JJF4s20Gh3zU8JrsUxusII0X+5WJnQqlbHJTCdIO4bq9oSi0jHs6zagbp8gper7bZWHU2
3eJbl4lk4iBbolbfda+dm4ySmRPdT7rXIvvGq+EeU+1s8xIRc8tyTh26dx2rmHkdPpKGAeYDNS/5
MKwSQBmc8EyzJUUpvkBAn9cJTZdkc5J517OG7AwreHPVT4/lsPULfOoBHskW/iq5LVqCaRCryUC5
GmUSgqTYKl5C0/tYJZd2MqYUJkGmIwjNon1uzEKCoKCjV6ISw4y6tKhAjuGK69N0Jd1vYRlSo3ZA
WhrdcV1PgKCXiOKaaODGlWfoS5mF5ujVVgvARXLZHyr3PqExFx+Ch8Mft82Kio5pi0MlTDp6TEe6
AYYd+Yh1xTFQiAIOFxISkiq1Ryix5s2akP8RqvfADjoxteORDq9XzvZ3LQMrOetBwFf+F6qhcpyK
yMjeDCoZmWIuoqxtsVdAEqCo46XTUOglgppJKuSxPscRZvUcgRAb5oQnNcIy/rcor3kA5D10/q9M
+fKs0PgizawRcgEuGtaYByh6LxfWvMeHNicfaEaOKUzFiBLg7j+94BS/cR2r/X4YLi5fizjmCDY2
s+K/j2m5Zu/zR9XHD+RSCvy5IrI/zDdld7+y3lRlVskZqC4LX7ZwnyYNtw0o9IM6iuYX9GAnQ84p
mL8axE2Sd6ySoi2ZLFCjOTk3c5RnW9UEihBd9sErC7XO1jvb/y/LgV1xgFhXQI9vrWH1vqrUfaPm
oCg+A8juZkOS4tweuyQqZAeQZ3rXw2avbLkn+zwucTcR76tEF72S0GcgZrU2tB9Lz3gzO/KFkZf5
Lf7v3SU/1uy+qUq1pV4qOTS+W2xhli+nVqNFEIpVruL13ai+/+r8tsVobelfRFDOg4f/yPb+kIPc
1+utsr9M1S3wDrIkYGR/iWG8oTYl4CDHwoLpuPy0sDNLvA5ek3Vo4JnAyqnrE+4Uln81oCkZ8RiB
M9ATmh+8I7J0Vu1fixzP1kJrz+4bLpOya2rILRBH35f7ZcGBck2AaBkW0RppJIXwaGEKswnY5lV6
kd6fTfPz3QcYacMAseO5Tee5FH8nY6FbeWQmOVyij7IzgmDUa9AiSVfJji/BWHYvh6/N9Wv7B6iL
GxAkQY/Hnpdk7+wLknEKYwP8gKJ43C+p/Ra8nzTGQxyYXzqbUF368DZH5wjdui/HcSm64NCBFpK7
8EEtgfRnqoc9Ch117hyhFROCOylcSEuQl63fHXpEMDVOvIbxF9g9AQput28ZmeyniHDcJBqWF3gq
JAseCWmy3VxHCGJ3NnLwcCx38q+maFO/2ljQRg69yFHP5zjLyvT09sSSSD/PfkmWx8TzUmDROOok
hx2u06Z+1yPmFSHMAd+jS6hcFcuHGIWj5nc2g/InXhpFgW2ScT8uvChICdkgRXXQgalpocZByYCa
xtO6XPjPjfn3V2Ine99/zuaJiFZpq6VyJmRroemIUIZh9/403IRufxY/Zce7BcE/Z3pPhBk7UgOu
PICeXT0qIhLcrmyOoPQfSfDpbOYe3lFM+had2c7WsLkQK/qSwPwW3jzCI0i8NsMur0UsqPIr+qsJ
Xhi/Sa4DkCWGT6gVwrLtH7aczSjUN3zl2oykn94+EPcVRXSLevg5fequhLkGtDbZG1Pkh9EBwUNU
lzPlFQ5M2Ko7R4wk7FndNgSL8dBWt1yeD/CoWcFAoFjpAyAAw3Bqdk3+V36v35LLjKqoaJ+SBZaW
yhOCp47IV4VfswoJIL/IAka0JezTKzKki73Y27qbuj90wj0weqQ+NYiV/3yNrWOQP1xYuxWT/rg7
zKcdd8gtZaFtruXzAPfwG8yUbhETouXpbDvc/2bmOsWE6jhAXZWJCq/bhQCszjsybVAXKsjYD51r
BWZLsoeh9ump8CYI4/QXwnRnHuaT2FtMRYaWaB4fbIwBZ1XN6do4pUzzhYNcJvRkiWqvVs4eww53
+bmkEOw89wbGkuZ6salYWRqaDS89bVMD0DCFe6T+5/hn7C5lgrNjAPIPeauTbZy1M2c95M+f07OO
7jNYPrnQS7MoR624XyInF1x4e2i7A93Gilsoxmm+TpC+wCwvTk4dSY+DLGKc7z5yh61gl9KD785Q
QfFJO1udvukZyEC5GW6D/gp0azMrMPRMqhCokYWM0tBAF/H3s8H8voYyn5yo0tEI+6u5clFCDVJ7
c77PatdJGbMHHohMTLnfHUrTf+rvtTysmvl5XVpurF1YnJlhVhRJ22DAiwwqDa+Htns4WNWsmSQv
X1e+I4DO+A1JQlInCBoLEt49lPDA7xwSZ9gImmPvQAQbXqWce6jIo3BQXlcfTcyfgWkn3Vxu+d1c
NuZwx7XF/3W3jXlC4UocqFuFPiC8HJWR+asnMHGMnocOBhaUZeXnUYfsDucNAeDPq/s/11nz22w4
51X+NujdN05FqcUSPo6+nOnRmtbIPqMkajoG8Wyi791J9+ggYyvX+yGY4MHcFqluZTQY2S7f7A0R
rI8Sb1fVtjXCAwBjYMKTdECN/ptuD2tlpKvsInyoD7Hz7XBFURUmgWncBMUnTMO4cNw8BznBHGHr
QkdyCl3w6Luz4fA88uvqK8uGKO3jXgw4Xp8mtRA5VF2WWWmHIo7fbtAVPhcAVWXio9nAFpfKqWYD
K+DHW6Az1XaQBbQavGoMzKaqNZhBj95wEa+JI+OnRxybByKEQY95ZgzoL9E5rqgjupQbnea7dEmq
2CnvK1HpGXDYPMSln12q1Xxu80NKu80RpooSdT8OP/dYG/DgE78S6VclqDe93iq8UwZ4EEjs2SKq
h/BRvYO2d8rgc2WlVYwsGYtGjvR4pDRrlnCPlPUYKO7DOa092XksKjNtrnZ5bv4MeqSzETBpGUBA
nf+2CzsoYR2gT2IQmUPWv0v6QHBAj0mxn2fLSPqgnuHyK+c/XUgt6NE/ksXtjXbl6SBivW8qHhFZ
2qKzXGwJREvZtM/lnQQOxP2KVs0Sc5goH07jlLde7TCeJZagfOF8qruKz7ttrs1SUKqXm6ivCIhD
xj28ZMe3KlkNPfDKFQURQ6wb4b/GtF29OFQgkHAq+wSKtUqxLYKwW926Lxk/CLoX0jNcn7pVcqDu
n1iCQSA8hQ1egO1TBzanm+diuKs1nikujjA6NJjOpBY9jrM1LgLmdDxbIoIl90rTXhJTEKZoqrBE
xovuc84F4bC0s7+Bk8sKc9VwyGs07HSOW88XXwUhZ7PH6Xl/hH1CfnkDE2NLsAZEQAQqIMbL90QN
URf40ZSwYPZPyr/CHgv3yiqcLfnfqqsbnbsNrOn9B/zkDVDn4MqgJm3dGMrw2iQVhSNDKHzZKUUJ
aZeh9jz3SAT8xkjGou8KzM92IfkDoxNWnCJC1vR20Kl2vL/Ca6x/yAC4/j0F32/2sJ21kLYBR4d1
Q6uGWZesu3jsFFsDabdUtVc3r0ShgNJJSlgnw+MJlDhTOS10rGi+xSq+L366yc7ImTjzhroNVGeV
nrq3neFB2UOEvXstHeUWlUbYchiWC8rNLwb046Mi+r1UcfmUXnZwuIijdoCgSSkXmJt6klW2Z8Mq
ZR/6tAsjJiimJwsDvHRGPJ6t5JKkT6MamFMa184M7cntI9cuCX9K7x7LpkBZGqAEFQs3bc2iC5xl
AcSB3DwhwHsR/8MpPmzlFa7qTFx9x9sX5V8PxwOHP5f1uc/9ESJ1Zvjc+Qbna6hpVXZEPjaSMVOV
kA46TVdG/h0TPzW34rfrTMYTFL73XEIHXzwbb8GrIIbIKu+GuuLu0MtVuv2WhvlRVBTKzhuw++Px
hauClZC0rOpeLhaejtJMcacVRvlunZMbFGnkEoxxcyuUJpmbv/Klwq39PLR9UTfjFNBztqaIZAAO
RLsY3mTPgisCVIkqsZ623gaXQezuk5wEZITWhGKrAG++IuKOaLXbml4WgFOzOr7NanmXMs+RMaM7
2ooytVVaWgSgFH8RWU/1IN1ozuXmQCk2AhIoDOYZG23TytQsbvX6pgQ82+kJdz30ue99ujVZIhi1
6r5a/4G+U41Ij+X1/e4BsdcAiosWdhEfjYWFPPPLBGdcH2WWiD2x9kDTp9xBxjLdgcX927Pd3V9r
1W5f6ltXZYN25Z+63qY6pMJkrZTwLtgenRwrWU9eQmnhKaG9kRcDLUr7ezbITVenQmWDAk2e7Hzc
hH61R1BuOU80Zj43lK0XqhqkrL5SbUaRBmyCPIYVvMgrSFhCANpiLM4nc2v5bOwI+yqrn3YhdpBV
tlfCX6R9UVeUEDB25Xx+/ubW3TaFbjokCjOX65bChcL30JjPwNhbNSgpO1VMld4FnpkxmpYhZOSU
wpX8eWXmwZQfyn5lJRpJk+R33x2MiYzb3j77d2GIXge1kIO7RjH7iqvSw6ccaLsAZnca0R8WlwQM
5L56RGtuhlHfeOJqlxWbn/I70XrkVFYLw21w2MJA24kePUbR+UhWYav/kPZAcUouk0KJ056GRcNj
msCqZW0/ih6XDHPiSSrPA590Ds8K2MzDh7xeWRKvp3FznpbhNlZk8nKsTcwjdFtzgnc81ay7H7tJ
x3KJwUgH/VqrHMz3/jqzEWQP1hP7GU3Kc2s+Dt2ZVlRacQaQV5Whzu1euAY24wIpH8jTwPdIF+vC
kFuac9opgmrPODrPrJv18UOsahHz7tf4HeFW6sqnDYG4qtub34irU0dNMtWnZrlc34Lxgq7+StJ6
5NXZyEgi0RauESHTBGDzxQMLcUtXCVHLwgKclLvCTJ250Uq7488vyX/TpIhDCtyY+SoWd3QaHONy
P/EJItrbpi/X5H+sx6JwF7uOogsqmXTdy2SrWii7M1ZwjxHkIgVXVJqBH68i5LbfFsKQK//imC+r
sBFBpw/ftUc+B5c+7JIdbt3SSj41BfXooEOdBTyQVrhz2cwy/uWLBzAEhqhQzSmhnBEgONKNbF+2
A4K9MGH7vUXYL3VTXM30K3ca24ysPo6UinlIOxgiY9D8Yl4L71UxKS2Bs7taSkpgwqyzcTJ9c1n0
1j5Oa0F1B3/f+RVFPI6RbowM+xfsG3GzzfjK5M3dTZTaS4oVTHtRTtdpMMiY1I5oUhlR7HDSc+GK
hhmhXv1IiZxwKlCMYtz44G7yBtR1mKzljSSUzKJrYA1dLirfB5AK/N19uzDeZVaOmH0efddSFu6U
m3ZElW0Dr/H8QglZCg91zchGOhGC2co4oWCS7u4r7dtZT2ulC1YKQhyvkCX7rrUEJMx1b/o9Z7/1
yEin6XgE+3p8sZSuevwc49pc34q9waPcXCdqkAwYM9j93R9JXMPrWJDYlqSDUiqkAG+4pbe/eQM1
RIenFlJrNpxfOAtJfTOMlCr2qMv9VijoW1vZjX1g8S4y+c7LqxPGMNSaGC73sLD3Zm1s/hN37rnO
JAaMn41CKFnjGDZcoc15wRydE67ohQN0UaDQZCDUcfb8pyOIHSAdnDH1iEUhSdGwS53tVvNPxGKS
o6IrouZOhCuhy5EVRqpVxYCDlMid2n1vJZ9Vmrr9NPpckyJ1+QLZqLuh6Pbq28oSxei9nTzZXu7Q
lRGcZ9mlDCAXHjVlaIA+C3YFxA33BZct095v81j69xbcRIGS68b3Nx9slOz0syQd1XviDhy5fRv0
F47rar1ysbhoh5tsNr6fA9MBth2WrMv+lsN2t78dve5B4K9fCu6lvnJecMp0dijDdNzpQKOLs45a
oIt5rfbVRBoFiINa7nICyHHeQbqNRSWvWzSwr1/hdjT/Ql2ckfelLz3cCJR1xC5Z9orVM8IHAjXs
lj1AoACrS1LVK2Jze9iEPVp0IQ6e6XyWFxShWuYOhd3w9BzqP+WjG0BvlClzMNUe0IgJ7LzEiGeI
6UyBsDouSEyK0XT0uNetpmW69R+mUhVce07UfUBvvAt9oORxeHxnr0RjuYQezM+QeYu93PSKmJUL
f8lBoq8QttBSmMO5VjGXKjQ/PrrNws98HTHcqEk1DL8n1HD5gHp2tMv49aksaWEATBoistPuW4eq
0nohs90xGXAayOHXaRhOSCYEcIn/GqxWdu2bjMmwRIljsTaPkYx8TFB5t7pDNeXfpOF3+YafWKgY
vRJF7VGHLcDQbzG1WUZNzZfbMc7OQ12iadaisnt+/rl3+F6IQ2+MkjizmVeMeGLYMbI4cLdCjnyC
SwHX5loC8reytebe+Q/Gw80dpV2ITw7JGSI204EiS7XEU0TnPyyBRw8ptxwhxwFFSZN+14yrVvJj
2CbdbL9lSRTXhf60ZvZRKZ7i+hWcl2IzGvrjibqUZCDzlQbs+AtxnU3dVgBiZDLeE5nplmXkxoZp
+JRgClS1t8uw8Owr80ZcNt06tKjWfo4s7sHkjRfVw3JVRI8FnBQp88rpPlHVZVMYI5FUxHaJV89S
ZWF2YP5Jq7z5L/i/UsykZOA6QZL0C+2q9uzybpx/w9uPSbh2Y0FoGZZcSrT3tbJHUMDmcktjKtO/
JMMsM75F6xrsIvJ/AO94U9tKJlOv3vFCMfAfG6j/HDUnAhvp5W2Iy4izGULVf3HwZOxXviz5jBt0
QxDeUAkHuoukWJXvKlJc8KZX3qhiYRz+5YACxNNSPMvQkaUjnVjTeU2VBiGcdYog9UzyHFLiU72j
gP0yH2WfFlWpB1XWvgIw4pcNQMdWssq2Pbop7a1Ws6xrTD32OH5GpqfJ1xgH+bj9tlR3iouDmEDS
0QZjC38TUF+Ggf1zl12QNKo/ZMVQiH0cVNjaz9xwIcx4i/Hd0kjVAc2r4nrOTj2IB3P2pOL1dhnu
8HCpLrliQzAQi6/f/vmriL6uxzyDOSZTsdix1MTzGumtI5Tvj9MkqIzF2ebXdYw1y2C9TnjZMhFZ
D3uzNMoj+iJt1pg/9+NL0Kv+5cm5YPY7hAygPsmDSMPJbzXY9lzLN4JAMXTNgp5pmol6qjhI+vzA
ya086IqhlgpbatTGR2DNrMrisPglm/hkunSJCSAqQX64dHJOqNet4xR3YaDtz+W7Ti6tob7kuP1S
98A9iTZrCpIIL+LZb7QwNJPp05Yc99xQTkcFWv0SOBWntKfQDST8qkOP1h+RwRFgt5le9CNSspFK
nxfCBY4qj469bbg12+3oo3rlT1z15PHii9uQGQkiu9e484jAViyhmxkEFHeJj/fhIWmI8JlD4PAZ
olH0y4eeFItNFev0s0XrfFcVtMtIwxPPBnMOkM0+Ne1S1rUJFbXK0YqixVQ4CusyqzwZZ2TnMITw
lC6AXDvCCAhqmh8kv+FPho2diWkxhurUqWYm7x6Anb88DXlT5imuM7BhqyILKBKoRyyLRgP31cXG
94B2s+JZECiD4GiXmlMsrmp24FTpcexn+CHg5EbxeE7yz/+pK9SaPc7oY0eJkMWHLd3zwVa+qEtA
lgyD1MbbKoHr4FWqeYThWjO9mKrr3yETfPRIP3lPcOvv0EKa7f3M4pL+YoO4s15y/s4hH6N5xBkX
F4NvlT4/iZ/CW0an4ys01oVqcsVMRrwPzVRrZgHVMV9KG552RzD0ApTWPWV19LADxCoMc9UlWn9T
QypD4nUIf/EbM6LdAYikJpiCfpBMic/cSgHThAoZA4sKlHXg4Dy28mbnbbxqq4+MWV02PFneCRmO
DGRmFWAaHeDc5Qqa8fqul3mi9h2bIXxmi+seWcX3x01XovO9INFnTwCEqtNA9T2NJN+igzZcQTv8
I2NK2pX/2gw2gsT0i6Iqn3hEQ3xikYsjzCwnfkeOvPFn3feEIMKGXRr82otF/DtF4kvygv/o/VOo
E/7kFG9pHIMAIU2KaccS56ndr38hKx1eUQqvV2RYKK+GRk5Z4CyVArPbzKxcGub+Io8O+JAls0he
PoxRmzqDcls1c3yRiGBx2foWF3pHXsf/Ra8OZKVEp726MxT6y5BYskKd2GKRUgj2NBlkD9Pw+Aw5
00Y3a1N3y0yXAime5Hg+INnVTUlXZ3ys1Tsd+aR3v6nLW14/tRGnxDYmSz+LoS4kQ+YZ27P+DVqb
KIET+OV0dVpURLna2lYS7lWZZnk5wnZNEzyBoBNcEwUhz/53n5xzoRezto5gQjySAfrGZ5I3eocI
xHXQXsATqDsYgqjNLpw6kwwggo/dkhDWhz4nNq9RIMuOH1lfmuGmxLJJDYb1yUmlgD7T9WP+mli9
2yZ2Qz270wMPTFn+qKrtNoUPTZbz+ovIZinQ6xs+ugG/ZVLR+yzn9S9NDQ3/V07LGzGt4s/CcRml
D6PWLXGnAUaaN79NgeJqyT++lsBJ849GWGsjdQxxtI9axzp0vsKUBmzXtV2bjRDaFQmBAu1wixpc
kNsPKq0q4+V+MSVcQBcmLdwUXKBZp52M9DpTmIyfcqL3ByivI/R3TzuEFRZ72/36yVeUTGCSrL4d
vf+hJ8/7o8KDT5YHl2LOpWsiLmx+I8Ld7U1IlMB4DE9lSRv6dUcRu1iN0D3M1FBrK9Ah00Xhideq
UY8bGacx2Rj70bS92hIoRDLHdnd7gblbpNxPebSVpHoDJ7ZvOH+34VrApE62uf/AExcspzJ4VVt8
gA19BMmYcWW75XRS461kLwa2aO7MliuI/eN2C13ZgBu2i2/G3m3aFYvXcSoAwpiLxFRUGjMMkxRa
GcQCCrR0DXPxkHUyAjR7DOsQHdUyz/PnEziEm7xhoAXQRbWEQLLkqucrYsYO74nWsyaM/TZRwU76
MixAcy7AiHREeoRIjubL/WhwrOlOT6cISAa7sGi0Xjyn0bUwk6SPDpPZEVKBqS+XlXrKcBt56dIB
7h9iqy6rKTLC7dnSvaoYReYLnuzsry4sRVfjbS49IJDNaAgfpvB5pZfZx+ZEnjq+DIQo0Zor5551
n+9tqgF5TStwCRjJp9KWfHKrZ+Q8rRS9v4weUA6v2nQ9A3YQ2cW14Nujx0LfiKLGN7drxpyyhXyE
U8N01xVQ0fyeGme1EWQ9AorVZqmL4j1M+zK+bauqAAbRZLGHy5RLW9AJyh7FVyzFHu4leJuiV5Sd
t/zvC7QiSvz10WdJvgPzEDzZWkqym/T3pc+GEpFT+uQaakVc3H/uxrHdEQ1YUtUz5ZFzXSZBUjP/
LjQaNZuI0NLodkrv5AAMEREBiGn0GDjlG3NgooJouPSzM2GfAie58k3jRmdDb+vIBsJw5GrOeXqY
/pKg8jWEUtK5JjzIfrP9BBOCgsgavAWUPHJvP1S3OL1EpLNAk8Axu+ehV2GL7b9PtXGQmNSkEAqf
pvYHpfDQvFRle7OCmHUiQDrgZ+P6IAWgfrZ512aw6UrpBBBBkaAWVh/GTuzGC7wEaIDdFq+7LNPM
tzRo5pJzQy+sYI+py7oV8bio7oUzN8gSIVwbxuhrOFx1i88V91UQjJe6HtLm6hjdLxQZ+Sw+Y9OO
rafJYqI1Gi5iv/TY7E17J3MpLSOcuiqss4NB6M7JlQWwQjelHW84CokDAEmv+7oAptx+WjvPe8+D
oNFiprC1yCXuS/EMeQJAlvvgB7S7nku+W1EuUXro45tIE0PgvlDhvtoqKfdm+8DdQZv0+DT09oIj
v8bdi8kHKa+FekVMF8UqOutCg8gIdyicRaN8UDqlxOrCLEGRLUbefpUrdxlcNBnH1/D8I7HjYUJO
wVQYFLXTL4nYl9hRvK8PS0v/tzshIg4/YjaebpZGELLJv7FENQDVN2l2iPwImS/cx0WsqA0hJiTx
V/yMyI/eY7yLTNUMa2HLzhoeASisPKdpmapLYZaXcXpwxX7S1sLIaX6ckaUlY2Ud5Xt+3IW6gMeC
SNPoxKHRHvhvzscg/77AXTzyCVgvVRYSnii/u3SenN67WvEopp/KPcNNznR+DF3XNnEPW1Pr+T7z
XJuCIZtylPTXvERdPLZrbUzx7nulLpUtU6wwmVqCT5A3g4wmJNkVd3AzLQG/pajZXzFwBj2C2Mwl
cDYgHQN37VCg0jkbz+S/CaB3o9e07NpERNY7yhUypskgnHa3DzUoKLaSQNCW+ksqKMSU8XBvA73T
fmOzpcKL3dca7F6Rij5Ed8tXQ/P+aFvvbVitzFp8LnSlyvOeww0YKJWzL26Aqb7xcNeILvXcKzfo
T2DH2kXBndmrKoiEXDEUWToWtpCePStgHiWWeBgaTq3V1379a98OXkzp2FHFrypQG0C07ZoJXhyq
TVaQhvOVSn2aRckM/aQ9sjrPklyHIFw72pDpAuRMifz4jvvhe3k39rNWP50xXuPk5bRJ+CrIoGvy
s2jIioGX9wuiJR1+lwcVkJk2bSbQFkqPdbnV0TduwzipLtpBW84/HZcp4ohvcU8JZKe1H9r8esmo
i21RWqyzS3v04a8dyP7uwz+e9P2SKcfSGiWBxaJtSkdrNiHZwphsJ2+ThnsIqYHpICHbcJGxYV7B
1VMGRq9eXlj9Yo8vdrSJBi4b2VYVnwk3paX/h5MygSXE3tWMSRhYa2U+HAYM+09KxVwBadGWWof+
GHmx4krebINS5ixIC6TB18F0XHRDL1dPYAtoN4kVZrVywlKw76gIarMDwfrKxjrhrdfDMC+hCFI6
PhSQLkqkaW8Olnti1AoD6LY94feiq05Ew3pr/8Jd8QKcxGH2/60X1FkKr7LmbTr6R0ZeuYj7jbtZ
wHDSVMGy0eKiYZve2cG/p5ZT4vAZi92nbQD348RDCX6eqs6oI/lTqKNyNxXtKS3EvBU/sDkkQR96
A2rDC2nuBJG8GUMV/K8GnqZOh+O+ukGI/xCFiMns3Xcap/+u10dmz42FqmBsVjHvaU8BKlRrP5jl
sx+VyRDVpxA2n42br5XpfcQckF1zB5nQq23neMmQP431UF2ZMzGLsaK3GrKkXEEx/cSuA1+fEKRx
Hg+NBJQq3yMq3cxlYNUAObnMO5U+RVEvzk6643anHyMoXa1a/2TlUa4AJ2Sfa02+vp0LziZ80IrR
OhCmT8UMy5XUCMK2b6hF/jU0IOXQgFzuE7mMrR5SQAViKDPi+4AhcqWY0sOD6rC0SoEMpUJ6ZEVP
6KCMKHjWmTkHIqiMJC7v899jJgrIqNJ6650Q+wtoY/UD4DdcmG6zN6o7Mg05BN1fMl7AVlgTtlB5
nsVxBRWnhebRA0wwAgw3mWai0NYXCqTSEUmrJPZYZSHkBPtTxWpciCVqOEjoZXE1U+TUJ8S+t6/Y
jHb3VrPTPGLgxuSOJXmkxKuShpr3uHzS66Gf1T5a3GKfF4Hj4IaluEyC0SZn59HyyM7VVT5/0+LS
toV4oZ7NKjDeYEHpQ5x84w/CjRVtsrP4SNax2S2CKDQwOLQBRUByyvOpZ/8rYi9I67OJCEDnjkf8
eaNLWqUgmfPBWctcbIaSsd4KzMCrE1E2Pl0bBFUcV76Ui8WPWXQJNRNgOXmorJGxjyRk4ipuwgX0
wk1bRBnaB+El5PuB2/4J34b800WGoS8TyPk+xKDgYgTG+SElIgcHU70DNihwvjavZOcfYYms3HJ8
fcGWki5mn1YYEtPPXk/7ATXK4MjSamUtPHmlZYVvXcQMo60OMl0HeSXwh443AxEerwOm687TKlne
MY8SZVVoYIo76ILHvXOw/BRGiBY2G4z/lSowvwti8VrXLgQ9obymutvjTVkrcCl+rRao4IB3sPxh
Hn+urseQNWE8MEvrBkyGuXjiIjscOq9W9uE38QQ7f2+H9n7KGqfHURhlz1EUKPKDNETWIw/CovzM
41Nhxps/7FLAnDqNeBEiHk3rm7cogxiXATVoVSJOupE5HaA+Hjtjgeots+SQXoslXyG9K+IGHMnq
W7XIOQOvXf0KhJwo1eqA+MfsrBp8yVs8wrtij49mntSWPCQc0oFHa2F8r5nK30IDdyak7gMSNxB+
ORJJSzDjeJSiEGP8XQkz/Dwj5nTmJzc0uFWOjsiBF/gRS5gGvWQ6gXqtH9OWzuOcNfg1mhykpjqC
LHROiVj2owFomqc+epNQmuZ8GrkxFvf2YrMZ3sV1QzCV7UXfuVdgw+jCjJfkbng9MRXEm4P0FU91
GDaJCo5mPBrXAkwhMzVoA8GJdJr+bTkkNqxeQEAj/N6v5oQHdnB84DYWib9cr51dID2T3jQ0NHyn
ckmPHOEG/tTnAhQawtU8MX81zdY3wbN7rZ9/949oaOUrRDs/F4im4HSuEvrOIDNJO8+gr0qN2tsi
jCEC3xuVj1jPjk1kyhoHnOnfOxQ/SrCJXZtsoqphjRNKqwGvT6Ia+Vjg7kcg8KhjFYiluy4DWMlu
GkraAhTDNx7Fc0PojicwA/CUeig82OP9PfwEpk0y4JNzYPu2PPnkYkfygcHjNMdBoB4YLQgqjO+i
x659XMiSxmxGoHofQ3HI9zg9JoTIrq+rMWuC/vnpPxgdORRXmmQOkrNaQDCgocKdoiwOb4fz/abY
lIIcytyHE3xvNFQRPTcJYd1F+h4/Vdc0aZzmn05Y7X/VY0arlDCRUtBFSPYyAZQTrBd0Rog9jpFR
CTHbUMgtYwoLZWi7S2gVaqpHha5NDtWHcmaIACWHhMYqC2gOmRWnJnaooIL50xOW8HofqQlgl1a9
TxNuBxjzDplfuxPR9ZoPYMMouSW/eyQbNbEj5+gX3oCbhIDaNayUR9akj85VswlcbhHpEiHFL8X9
Hl3niMT+lTgt7AJoUW99DI9TqvwrWqdS2OP1fafSbOUlAC7nE95Z3rw91Cn8Vrlzxeq94Fh/ks5H
Dzk0dfZBbaAxrjZ+zbNdwxyRJVj/QxtA3jyb39nQbvwRxBu82ExkEWH3sODiwfbbjSyi5fYOd+ls
zGM+PWmEMHJT7V4c6uN6W+Wp3ZI3pdBhuQljh7wiuaD7mLsodZCChmqO9I+GGS71xTG3NQpTgatI
PkhUhs22e0X/H3D7UY7emzgj5BH5ciWKwj4G2PeVi2ULIlvbAIiBkyeDLgGC34x/mcCH2ch3UDj7
rmvzLrQt6dPg8lX5qLePksqGL6ZhJRZp7UnjN8eBVy8iwPLIvNUE9LLcvDh73XkfEixOmfbVLTdY
BmG0h8U3gFOTX0biuhb0E5fZQf3mRv7BCCBHuHdpn6GHb+uyCZDc1zZSz46kPQdBtPDQC72s38R+
Tlt/bdzsZbm5nMhuCl0ue/LTdAmAOHOc5cspe2cX3BNHAeCEMx0MDRVEQiNax/3E6qCkVGfHghGH
/TaNg074Se3TDPqAVO9UkHei+xwmfgBZ3MDeiVBwWU637kjh41u5DpdTwPoF72fYqjZes6oe7Lgm
YaEEnzB3mJL+3wMy+bHmDkieLShOEupcc7slM05hwv5gbFNaqaFUUxUc2oVaf+ZwFbrlsd6ldxPn
XKLdX0Km1zRfoqEp2f+H6JddTS4LWJ5gxjSWGFx/AJhst1YVE/cD5gr0tTfqMUvsaT0aYedluQoT
2DbKkySDFppetUvnzWQXLpQ4GgqLWzFKuIlCi4pCugIr0VFwQ8C7xqH39sUc1FNRTeJh1wIT748q
xNeeHtsjiucpOfc9EAxxqBihwDpfDSjMqvn5Rpc04RNvoQzPpn3Q4QyYFOAdE1sgQLzOPp1FvxI/
K7ffcVpYEzjnGmMx3lyDfOjr2Gncu6UjaeymdnjfNzTTPN+J8edbeZL3Jh/BXTNncOYVARyHsxFo
kMQKSokPNZL0X/MQv5uVbSN/i6O2bnjYifjdxmFiuSe6juGEBhEiLpOcBCF/KnsG8y1YNBxn0dtu
CcUNI7cEs/Mwgb+pKXK5TF/XvFaxgFuL3f9PqJfvtlMNXyAb79lLwIPjjCH8pmvJDb0m/4RVH2Y3
I3IbNgqDCKhwYUwWKucwSGmY/oPk381warSCeBZTtfjdl12K5obIOEbc/JI+19W8GPkOVIXDIL9m
Tev4Phd3Cm7GIOTIgZisT6iX1uRvPyT7yVYFkxu5Ig0XlEi5eoD/bM6kXTpD988161ldNuWTnFFh
2qfC6HLqxkcGIGttPoQyCZmhzCGbERNTm04HJWPBAam2Cui0YU0YzyyAx5aBkJLM2HCoj9M92l4c
G/XLIi84jNGEtiFASNLojBFd4JOqZrJFi+BJ39sPSa3K3oa5jv9JyUdK8A9lF+1/tBdCfiJXLfuO
EhUuyL1HzMq3QRNjKfiYQd7BkNoKvAjEWT4uQ61w8cX29xCntvHRvuHTHftulr8dwUnq7yG1hmf5
lVVJDgbvWfvaZAQwdcVlj2/bmwth3j4XTlgOyxkkNZjoo3U5pIoO42fMRiKqEBAwMR6w191nJtfh
6M5TqzUOxdG0q/2Cs7Z9iex9NnLv1gE+EWs6t0opo8HypLeSqGcUTQvt8YdMRMjTyBSjGbJ8OEcC
Who3GVn9poluNhCjdwOmDOCuxgBnRxKR7NVVGv6CX7i15Wf42JKRnp9ULNPQfK++3E+4XX6wrwVJ
E05yzxYIN1NNLm+xMEBM4My6K9mQCCCZCkEi+tRVkU8XSm7RkmlmcphPSaBr0jJDrg1pQBIBbVsS
9jhccK2QQj+xySST51euOI69d1Ja/afIxX71puSGFAdU6qncniZ+zwMasDihbJqf/GYXJJmX6kYs
MaYIyXegusctrJq4ZEQzCCyxj+F5nDrudoVPqamCdwNx9pcuey2WdGsL2fCWa24TX7UQUJUCnaMB
eluIrEzwFZSDta++u76S+4DudO55z4E7qTHgMd66lD3ebtWVEC7B6rUHIK2X3RU/S804UBdXXcSZ
lXoaxg+VzD73JZJoc5u4d7ab0COj5OdJ3Xb0Ng2K4+F5r4fyKrnp6ZW7huygx7B7P4acpKqtdu6n
B+37jhGPWoGfkSbqkY8iqCoRbvjOfoaRpDGvI+iJ5lNdN18p+WXUYLHygdBYBxfpSFg9bDAqdjMM
z/x3YzD1q7VNi1g6jeaSxm9RCsOy4nwASzSzMUCx9lJj1oddxl110Jy8qF5gRUyaB8tXq/AUk0IK
S8dj7mlVsCCDc75B64oq3LC7DLeqxCOKhhoHfkTv7hT+8/3F1RNGufhOHvxc9xGBlZs/DzBcvV2G
4G/c/vtCuHlRjp7koqoifb81b8rD6LDt/zS3txz3mJcn6Jv5NxTet6s3hZti5/XHgoDbi/0+xD3f
jiwL7Yb9JhFEYLQlFQ0UkOtYxGvql+udLJQ7MR/UP+arXf/R6B2tFa+MZGy5BN4rRXGiUqNNzkzk
0HW5Azo8MuxrLhsjc3RnqUrr8lpCPSAkb2r7m9Aj0pEjL09BJbPvHPfWIO+1JSSDIfLpJDWySvtA
ynwEyT/DZ03dMYPRtapGCHRFPgaDfah+/scyBUNVC0C7lNf/y3Tmb6L2yn9GDhIRkA7ovNbvRc1G
ZlUa3Qpb4JNd9RIuDdBJulOIxS9aXK4+Fh/PhSrZmbl5KU0SvkB7i2okS2sn0so9x9zLXR84LwHD
79hvt5D/RCx/MughpEVVP4zIKBPVJKQmuQ2C0w0tcCwapBsflJbaFm9W17CyDnNk5vy1h4rrLOea
fpJuGva+NVl19DwT9weu5l9rtkMhyOgeiZ9isQ1ITGJM2qqRIcSsflpc5igSK57MLFVmmI4rKzLA
qriV99Ei5NyyWpmp5s81t1UxH3+3YQmgnj1IZRzDbo+MBvWl1Lex/ea4DMpQpIW8R0iWRCu1Elj/
J5btfBvO1Brt4nQaK7uMexUP3tpXhuMSTWofxL3tgg/9Z0IalROMMCn02WFGRGvFD1XRosYF4Lx4
ElDGNhmdeiL5gsuyepCfXZRrqt2cnxkPrTzooXzaMmUJfeqQh3co6K6Ue3lh0HODgBTBF4rpb4Cb
4CyXSh190/hs9UZXA3BitxfVYmk4SmEaIYW2i3Alr7I0BE4ekd6JUEuspRl/0DPteuVykckHE8Sd
lg6Ay8F1Ui79cS6M6oCS27m76zzkNJUhqNYuJ/ydaOH3P/onSpipdBPCJqevUIQ9xNEAYIxiDJQf
IhcOXFQOUwH42wbsUED9aBrC8CvL++iWp2SZ3viyHBHa+57Ir9Uw7gyYdrgoT+UWfgk1+FlQ0vvE
Vc7jkc8QFoY/UFpIrfLMGi+uzVwk3U6GUEmb90qb3GKoCtinK4B5dqWUXMfCwL53p3/UKNdrShd/
9MF7wblNS+3GYM8YvrxoTz5MrDsHILv9WIGMWDJJ3nK9pVsl+JzHmi8Bvsa9q+HVlvKRVp0fJ73Q
S7ij0NPxP/+gvoh901nwpUqF/AL9tdMgFltbGlGxfA7kAhuNQhV1O+qqFMJLfX3NG32a+tfrX90+
nhZ7NS4TDCuViYFEs52uKzdOxCPBCCxjV/fJlseAj9TXrSwbfpVkzeLLRTTZ2eQU3I15bs5+6LUO
zY5h8QytdM+uzEwMwSMNI2tY4iTQzGRoTI1bpIJfselVL1S0k8Ace8Ha25hu5tSYIKweY1JedOyc
ijW/fF3TzPmgJ0YrVFOth3oNBrtbeFW2nqp/JyX20TjA+LOKZu/WJCdK+hlZ3SipaOCgLi72rjrz
O7+SJR6P0wswtwvklN03i1xGbHfiSi0N7wIghcXs0LPiKjsOSXeNxN97WoXjlWOwHyLb0a96r6Kz
jMu0fO3QRbkrMMNi16ZHoEn+9rr5pcePXgAoqRDoo1UTEsOpKXlFL3fz0rA5zQ0Eq17/TQkeJux+
5/y5IAUrtZSl7JuD+Piy/yLOHbnJMpNVz+h9ZzuRHNYNoNVapCOYjC5zldjlQkYEdiiWNGVsMfl3
SJD4ll/6586UUJ6wVVeATaV3vJETABeqmMe1BGCiIjkM5f5LdEQPmR23Q6Zwgje1yC7TbZywPgJ6
w6jfkLlS6FjKv3Rg7Aotg5A/px5MtKGzs2aXNHmetKFExtosGn5b9W9f5nqJpHBANjMwB+ZA2DI0
G5Y0fo7Yeh65q6j2V1N0+3PVXoanxOPjR0tvm4q27hQYGNjJ6j5cd7LTxGPpZxS7JhWty+uVQcKM
OKfRlV4l04fA9QSK02R3d+KbWmN2Skw5i5+iE0hhOLXBa23DnAgsqOkDBWusYnizgmMestO//v6G
utVxz43cqBCtc5GhwoHmwoG8Hsx/f+W1MQuIvOBYyp3+MkT1QFzxpNxpvmgOQ05nwL4KzeTQ3I5R
0HJl3KE1jC7JyAuIDJ45A4bUFQ1W5xGvn8bRFXSnTdjJgWsh+PWMxb8zhovpB968Yic6RUuTTpuD
hS9sCAvdJeABA+OwxjDqdwJCJiT6JvQwz5RJ4oVt70Dsjjf1xg+NBGvaX1UWfZjmczo7+rKE1xr/
onp6lvtrSQgDUpFWTIyF+BePGSH6Gz3UzmldE7J7i/ysV66FdwkUYhBSSiA/mblju/BLGk/OQoU4
yu2NAaPfgrqXGjfQeS3Yu7qy7/QyuyL3EVaiVAdZIT8w0YxKl/ZKmKRhl2xgC5TjS08sQ44fL0vM
1pqzZqrj2Xh4k9mwAbLiUhquQoO3MC+8O3OAtqude4G54tG+pCmLSyuMfR0kpEiCFqu/LfLoKYoi
QmMRZ/ByBRYhYtLZAnCu7CoEz23t6YrWVkackZEziY9D0DoIfAQ+OHgQ7/jOvTWzNGRI+c/el4Gp
yv4T9TekBCkfN1i1xAOTqKMJJVfSpEZiCsRZ3kOmIlwwD91l6D5Wv/S53x7eQyuvqrfl91wpSo4E
lx05M3IOWsApj6RQ1vzFeJqq60lUXsvBZ0f7IFyehwgo4iUJoiGaJkEZt5yvtHWmETyCEnZN/bYk
JkHwd1Ee53wBrn77+xTqPcRXYQizQfG7mZejytd35aUoNNQxF1a+V2VBCCMZmtTaPTeTKrqksbAz
ynjZTXrWKI7NxZQvywOXOboZQapEY4ufK6fS2pDVm/xhKBtCId9nSpqu+tBsGLmFU/0FQnsgaKOF
Q/Rf0DtiS8KrVo32zA5iX5OxwD8S0/CUmGfRWW8JIie7afyArDFxgRezCkUAPGVVWqT7mZyQUwvV
zZcf9ELBZ+phMqL52USP+mVNsLxElkLUc3Z4JvPVQjA97SQyzU4xxC33S+WG4eWZwicTQXPJj9YI
Vm8jJbqw16jYB317hRSCNUxlGMAowzRtrc7D8kJLv88R5Ip6O1xlJIbsHFNxdkp6cZg2v7+/iiD8
BNeRaVENAXv2BEINKaAZ3CuA2XQLjWZFq9lBmrrnltk7L9jcwnfH+OX0H+BjR4WrP8BTmVuZJal7
Nvhtviz1IG8FGrnWJHppf9+Gk6NVvL9Uf8Kz+L5T7+aZsdek/lH3S4U1P9wV4i9h6ALnWCGY2oVn
7iXM2s6pphwb4qGmpuGecsy5oojBnQd2epIHYrBZrBcWqdoNN9mvJpJb1xWo8vXI1e0Jwf8vmJIv
oxdLsc3e2iRChaFS4mkIcrHABYDwvVrvimSwELS6dAGrjsW/lkTIHmptTrQjxgWpQQRV9QyKVN93
ukUXytmCTeTfW36vAFdcqs/okev2Qp3UaiqP8OnRIU4gfi2OuQcdZsdQLrOYs655mkdJHHvEbwiN
oy/a+oNp3oAt2MygYYUA59FrsvDP5Udv+Di0MK1QqBHjQIbwx9iOacCiJOgyOdOE4FDj5OepQFKY
lFyx/mMr/u8Gw9PGGhsBSrXw5x8vRMwbhvUP6eq4qTgLc6K3q4kY01FMSiNdComam3EaPBgqWvzA
X/Hryg6xo1xOYozAoZfXxnM70ze41Lkd/eq7yBtFn4X/89co0uBKNp1og/AAVPHj/ZUDPhKhbeP7
xzY37sNKeYjbG01XmeEs53sVB1IcKrcX2wL4jO2tiJq8s7CKt3bCI/S8SSIAbmAoKIFU3pa/Y5J+
4Kkpx0puGr0S/TxzKVSxd41nw092umrncRvS5fJBkG4l7sCBHrOQY0m7rOTV3aq6yf9uDTC1/nZk
aXhJkMnbDvMiHB5A4W3ZIEb+72EQmQxbSGaJ0xpGOr6Uh6vq7+tKxh66DqXJNZ5ytGX8MQFCYTHd
Ine5FodVCW1XOSiXQFWIe5oUs2S1cyqFjDfIFIi1zrSG9sNC166/wBQF+66/ljX7Cim4nfQR8WPR
XkOKQbyXdtDkydp8rb4xjL6RpJ2vONv9aDs2IBioN8hCsvjjNvp4H/SR5pcbukbeyq0Xoi8dBij/
iT7/5v6ffq7SlZ/u9WTGiVvXXpvuDFT95lxnrAqModQrKW9AeT/vNnwKA7oH2jjcjWM3kum4sqRy
gPtmq+EvNohtWb9zfxJc2QgrrkWqSSjRqtUrG5Vjlsvw+xvQUCBr8YHZplijz+WY1rgSRhie5q7/
ntQ4NZq6BLf5JMgRZZQVka6XDUf5jmtFJdpbpWsbc1ExYGtxoh+062nISajtoC5FHSNsl2Rxf96K
Tv8kYqqlLUxu4zcZFmchjaM3Tv2EDLAwlMY0/Dj3tpOZy3ZIZcWQkih6INuFo+M3TNxrwBe2mLWg
YoiKVt6NC5KEKGZUTllg+Ky6+vog+GnRdA+M8jHc9OjJ/fFTBTNq4fu+r4JndWCyuFqvUsCVF/EC
2QsALXbTV2wO/FQhHqgZ29Xe6lGJmjGo7hLu0UPzcECniG6TIHpoNP9mXlVmEpuKhlAuei8863zf
ClSkTYY9Ypo37NmXnq2dp9+eU4kuhgP1GFmkAc3lY87lD+PUHJ/b8F4M2c3zzdJYxyDjJf3vXCih
2xxYuCQJCpoR72pMghOOGkI4scUK1L1ULCoUIqcGNQhpahKvaDnlnLDzHHLMdKa3moXQaT+PyJZx
3le5D8Ki07MO7UjAum5HtSVCR2WjlhvkMz4YNZ3DBkOPBu63iVN4/CGYSyud7v6BvExergIel8v9
zK9IB6cmJe8/BOsHNgwCwVYB8tjy3m8BkZhezb4Sa3ZLjde5nkGgkVudniOSnyS+cepwp/IABTSX
5Gzh3q/Gc7TYoH/C+Pw72DbJBc6ElqP1ZK68ugclaTpruwVRRdGDgB/APgRU+4XSztUUd7M88zOf
/DsRv1Js3uxP2CR852+nCrr3KSZa4kCW4nr6RyG9av1k7wSZ19PxbfeS+T30jNTCdlvtK1QM565I
o11wcVAGwIUryo4LN+uKMvCncI0Sjntv+LaDUFHBk8rPV9KF0JEDuzhPQTlYgGZL0OJdPZoUp/rr
pOvTw5PbNWbT8ePQi1tK525VrX/jBcYcHVokrOQaLPrT+tl5ZtO1n1J9iLnEDiwZiVyCq3OijPzD
189yoyyeAK2zuua0fR6YkJKEaXaRM+qFYUphqumpxjI9fSCA0rqVg//UH2MHotIUWhscllLDax4G
bbpA2UaRt9DYgu8o+J+AWDkhGc3WfiwAh/RrT/oM/Flmp+tMq0YVHExA04IwiBE0w+UNKA+7flG0
L/K3/7cLHlaiECup2ftKEjNe++F4u+mCpkgg9qonkuNtIK56UGG10eQg9TuPID2LzXfl8ss0dop5
s05uYDHwq4I//O6LerSoVc9+I8ltHNzs4ri1/mZHX8oRSK5nm8eqmVQehvQn1Nkuub7RPXpBeZex
ustcTKR8rGSvNXn4jwVvdUeh0z/0TUQGougypJkQ10RxxquPqkT/BG+p/VvJhzCa9S50CgDv0QnN
UtLPhEyJdiIS8uhEoHBgVMHK1ybiJOOVCjZ3D8lwvmQY/Io0DIWsKLRC66OcKzG896UQTqwunmuM
YEZfc43QliUJJTumZa7aaHvBkTtaFPi/vA/C8pQLkEArGFndGrNsQhpEXnrzUefwgDwY229SJZHB
XLLLXSVcGYez4zlWQebfoVygliPz6dqMftvxzc68GPCAhxl1w7DSroOm9+AAGFIg0begLhFBtVly
UNPtHeYwFxByrCrzOOBSNTG2SZ1FbzFrM8TpTjOB+Mc57q3TKMBJsqoF5HzfWEaiIvIdefARVbQK
3NIQO2+KADerdfDrgb/GacdZICPiHN7n1O26sXWb7LY+49d8AhSk2Z+53S0okCpBGOKzl1LkBXAl
jC4bfU5qUsYwgOEUPKT3Q7Dqt9tsbkYn8BQOq+UqX7IU4jl1k06vucA9NUeBEqJLqIlErOtNnpzk
S+HHviMJUAuiEd1PmYu1THC7LvORdSNxb7tZ5skHeoIdLv9IJURhUSZMcW3en+D3/Q9c5zZkjsUr
jgzWDom1W9zGJNI+QNkuC20KdJutGgfO4kI55vGqsJ3hRZCmGyeiZtiVKc1+TKhlHsvHiUop+j4J
33dH6MF8irs4U6W4CsaP9o6s79dvAcbUvDqWd23IVDQzqEwemhstDVjjHoe3so0Ja2zxbixgJ57X
RZJLZrqpSrjUKrwIgQ7lBd4VcY8P9RwZ9O4+6df+FBwqGs+qWb6Gssc028XF63CBkLM4sO5bkugS
QTD/LATBBgrYZ1PPwMFOX+Lk+2sjLXL/V/UDYBxuP+WQWktXpsjkheMNQS/dNoUo/Pev7pmHO5cI
1swCt7Rc31ihz83ZZ9XlCJdC/LQ44+Qt438SEKl0vOzvcUOaaYQuzi30LDSqtU/fmLC5O1yFGCc9
bxLkwDCoIPleiGK4OESCB3G1oNIgEXtnnJSbaee3Rv8kWy4WEMMxQ0hb/l7eCBqqeQ38C9JZ8sFU
Uw6K5cbiYghu529nCzvhW/CxpStfVjRICc/clVJF3MitsFiTXyWHnI5Zf0fK+3a0SvsTjAJI/Pge
T3fMrUZXowCouriSjB6jTSWHEDLe7DlbMhwezMsbYwZBi8y+oVed/gdFXvm7zkex0t7FnPv+gLP7
9E6LbKRBZemlIOQQuVWtpyniChdFasrq7Palyp8hJXQ7O/xttFOoHAIPl9zATS6e9YYiCQHKf3S9
y7AmoeYSel9jlmUuY14zs5HXdZH6rcCQuVFyi6+MkibxIO1Jk2zZAh5BZdyXiYMq2SHydhVMtoTF
i14w1+Zpwe4YL7IqnLAEuN5uOloxrOfm0lQgoMB11n8QblPDtZI5lHuVzuAufH/2/cqrQoqjrSpV
FoQ9oKvyuM9WDnsX3GFlI6Blexmu0+Q0+Zq6KMExkVmfCfPWJWBa2WGm+6fLQGCz8yS/VzLDz/PK
qKMABnP8pcBnfHqbH+J+MilwfrIjr905v1sGp8FG/ONR2WoRNXBbShxuHaNLCyLeDJiHLCBlqm2u
Q+t/LuSC4XtEdGf33O3EWWBotk+No3VQg2g3PP30obgsMovFv+PRmyDpFVS4e7SBU6Qqhdqr3oz4
1hMLL8dflA9UvSiwAXTVFVmPZWvlCFc1yVqaXQC/nDfy1wiGhF/QDpH7En4CHsO5TRu4EECvPcwh
iJDsvqRkQwEvBKWS7YKHJfInJ7j9O7Htu8CzUSQOv43U9AEqaK/Fx9OARkJX68dF99uM9tSMPC2R
EWwUmiWARvL1MDnM5RHJ1B2UEBU0rDidV8835eou1s+A2C5Fd+yrH2t+F1jctBMn1425bsIsfdYP
zx+0MLm4KeYQswuYCBJl5we1t4AwCXVsDix/Q/GlhS4Di0qOdFdtppUPIpmzBHW8Qpzq1ZmQkKqm
aoJcc/QaLAgQcICQTfbE8KH0gv1Rw6624pEAwcZavagYg55OHVlGPlG9HPiV+uu2mLJyYnE9Ow7Z
9o6xik/Pl/JxGHFcPFpIcC9nF+o8D+7ldIjwk6qtDB9Mx75dohnUqGAa9ITjXONEHLiPUyKDMGvc
tFhZMX86Azwo+BJn8rDH+rsnMEeefD0fArxpv2SzXHzBSY4VM9UwAfGmvnCUvFrTiM5P+M4jBKyd
MWkRZP+3JlVQ3tEogFQTDylhcvs7V8GahjqfIvg7wwzjBoxvQK+9obsFfg6WHIucdhLqCq70fZej
8CPB1sji0zgaUgiIeE5T6PfcWz1r+PYgGkTGmZmhjhthNcsldRLqamqffRXJSvlZqxFg/e9qE00u
2sjQ5QonrYQVBr/FkmArCDNrniiuK4Oox2rL5Yw0nWlUMuvyridqX3Q/43EYPsMRDgLw7qUvPAc2
lM+33GQcwAKcNA7VGpMaqIHbtDweYZtbtkzrH0lDOJaYIz+shFx12t6N8gRBczlRS6V0LvnEkkJ6
DFUrGOc909L9S3MpjXgUyoVHI8nNu2DVvjGA1A0Jn102L2AKZNdTPhjgNprC3YmCX28ucprY/ssH
boQXsyfiTXn/8AU5jSsXsH+MWqIvk54lGPUd2E8mV9V4i5tynaLjfQwywOLkjrnj/w9sf6TBbkK5
ccCVZnYb1j7vrnsmH6VtCjS1AEIYnxDLDETYbOIExenjnwIprYUmGS92FKOpOWd7Y7oW4um0b6Nz
3fz9H+LL48yD3FU6KYA+dO9B7oIi4K7VeCRcLZgZEQssQu9uWCJW71C61j2Qz/JPB3FnYIHw9zcc
zKXgCVTI3kdGGQw+bhdtmJ9evzdLL4f+20N1hY94jyq5F2UvrGDcQeaJn9h+6gwfH1OCcQyk3eZn
oBSLSTLTcae5guTc+9s5bzZdQ/M5vKQ9Mo+Vv2Xz3BGwvCvMlrFoUy87F0z8l2LNEkw6tAaUfiUf
1gPlY43EBM48nJpVMImwyfq9wwT+2+fZ+MFoNlcmlffWvLZAmsXYKqGgD3rNV9I/fZvTWQluiOad
vwmUqQPO5WOAKqnScqCXDCXMLFBJjsI2ennqdzqN+Kj9BCyu7aCrKe8PPfAJAx+Ybn4Z8cUoS/+R
eAYrrQcf6HL0je2Prk7Bh8zm7Mm+3QazPZW+spXf4kRm0ONDLhdQYQDKdCNdIIQ4v5oaG5kWjm6E
bPO22lymwlwdGVos37U1rFGesKg8SJbi4Z9VHPw616n3ByauBv46qllEM74JbxM2L6pk1YmreaA3
lHmZ7joLlyMs1z/NUfgZRCe+6eIjHlo2hf5n8TeDLEwEnAZpzFgZUxvqa9P/DSFWJ6ODaJQNEvSG
G7zcLupk8ZHphZqhbk/C8ZaW1qpotcz9rbOSexIzXLk7fmSZbZppXZl/YOUbSrdHtzPQl2VkMPoS
3EUUgnObNU0doFkZztprcz9/ZBSzI07qrxuzx84C7CaMPw7sU2WaV+isNUeCeSB5cK7JOdLEmMO/
xnBmowf9kfNTe6BKNlXd6enJU0L5V4WMxW5jQ6WRAitp8WUgiPeoy4bVDW/ChAcGs2pmJTZzO0xT
BRzrOcxCFae/+fHvhyY9DlsiG2Fww1JD2Z5UkboBstS4iRrPIGr7Tp1DCpjYX4uRsXiEdqTu7ez9
pDZOYHzXAgRkBk7HG/MgWJhjAkYmPKM1vjZ6nY5dp3YXt2ooyfjtfVj4wLcDUeLszkelI46Nvao+
rm1YAh/Ls0arPSJ3i334onEgIrFL+9pfQxoTVRz+tCYTPXYW5pTRO5U7Qitpl2ZM3c0ib61UpoBI
jt5B9nJpdrah4rEFZXgs4WQOktbVd4wRDqG7oqMms94ze5lacsfFnnOzSRGGzmQGcF3Ha2s4slch
A4l0sxcPUkfEH6Zi9eGYUsKeEKr/2xLt0MeZJOVh04z95Gfd0s6iGURcZDcTtLMrpbyuhavT/4G+
yRsmFEwCm9jmmw1OKniILS/ALwqAWxUXPuA61UFjj1EguXvYQ79Okg3EbnmSH92n0SLfO215IyZg
mxUrKuqoUcQYH3O1sVh32W6ApZQpAVuC9Y/c7oglInSjM5bEp8vQOxexnGJfsqV7dNjHWdKmVbkh
6FEGDKmU7XQV83QWpp99snHTrFxy3evaGlhWtqY/gBc2He/p+4SHjT0Id22vz8kFd4mUz6frz4wB
wn1hcKIWmf6E2CFYcX+MUyB2Jd3Gn3cAc/cS6PsWA4ha6FxYWxkS9Qour+iwFHmMG5lNljlbWrxw
UPAMtIVotNS1fPBN28iyDWIgmrw6QQ7ECN6Pz+4/+ZwMdXddcXQBZOnC4UbDFz2JgLr2QIuiIFXO
Kzzhpc/9R244xfgVFpBPtzPrpFhUxSTYTuWRqxPvBtc9ULGRdimZsuRc23HcPaZsFwgkxGEelF3b
Td3ZMbBJt5P0LgP2OLJxOow4clYTXGan/u4IQ9nnQMCtgDFB9/e719RchJ6GeTuJH841h+mpC4vs
Y3uOgp3sOxFjA32UHJCnGQSAJhAj6llWY1y4Gnm3aPp2rcZnXBtQejkHlPAePj8CZlEAQ6M/1gn5
XsX8wAzWfor5YaXEXk5J5IGs5ST22NWsdar/aJ9j2Num2S7TumGQCjjH8/pjSYO6EIC0CfvbX5i8
4kmaQh/ySs78qnZLIcebWA12GkQuLb/y5U59Z3/3hhWF+DFE3XsgSMv1FeDDwW671Q+hm+n2bLDz
4f1JXnfMUhzk5ix0Yy41Sptki20cvDSkxOfUYuQh7SEukWyKITar55DwcQEq0x6OdXMcaGzwZ4cG
V05jO/IGwrr+KGanHu+be/LCCpwPX5Kp9Rl0PhIDZqFcHYSz6LzH4CL99ix18fHL+2MhuH1gLFvI
f0pXwtQrSWApb7AFIbEylt09Qna4C5/2DlFUa8c2rsLwzwyaNnfwQSxoE8Hpgst8Rkr+5N3nKngE
nINxbPKhnYycSRXnzkiHpN4jek5evgYVFHBMjSmGH9byYWAl7tU6kdDI1by9i5tCZk4qVPI00TPO
vBH5UneHsUA/YoKO2XtoI0UnYX08pd/sxpH6ErvY0fTWCyKJ5Zj3i6my3181iT6pd6WZ0tmhT/sA
wThJEGpNe1TUXdg7R36YToAIRCRNfpy2TJi+g2refvMAPXUPRUxwd3eeb35ySTzXG3TpnHiDu2HF
scY7WS4vW0xLtcUJdGTLrMRriG6VUXzPTSEfWRtu9tXBBasSBkRCngEp8uHC9kdJ025IaKXyZSTU
HhFELwVRazpXR0GqAojKuPLujf7iwnsfSQ+IEEr0q3DDPB5zpFgG1aFGzVzjg3CvznHyh8HYn0Rj
oolWkZAXm629w+r2RZTrvIiSIvAqqFZPSD2usBGDAZiiqxM+sf+ZdfWkc4kdrpRSPEw8Zw92hN4K
31a0+9NZGPmpUm/S2TaEA8ynbcngihNcG0BMY536pBm/n603wqVeF3x3NjaSi8HcWlZJWCf+A+EP
6Gtjl6k962BWNzFyEv52QSsZpSe0k3Zn4J00Q5boe0UQZGAOTp9UxzFiinbXuWUAJ/Amwq6Vi/w/
8igMCnSV0qjvdupHPiKPWKXaWdVFyN1j9qBxy2Lgn/hQTocbXTUmpAIvMj3wxTl0ffqmbcAExpJ+
FkudAJZ2VlG1gZWpEaG6Rgsdp1De2JaozfjFijTIC3r2Qm9K24svPWDcgynTwN8s9kohfHb8TPSd
H3vZ0oTyzupOZdCIxx4jSYlx5es3HulV5vRUtio4gA/oDw8I6nHmMQTNr01j1PC7aP33Wka4DaJt
VEynZHabxkHn+nedhgZNLp3rFYbBY4q+XXc9/X/R8pOmw9X1Y9BP+7rgRBXgnjYT0rGeNeLS+UQR
/cRMr84ST9GiZT9/dXjpEgFd3++EnaySkACs83qxYBmWPRZr2khhS66xdAeI05x6n7G7peE+hds/
hA0piqj+wzJdUo5CxLnZdS0Op7Kq4RG4V/YmHotFmvvnuT18/Yu0LwY1ievX2ru7pBZ9wSzRLron
Q23x5cdYsid8+jcxjqDGK6EjYUX30TSYs3Oh+zxkIyiowHK73UsJVhU0hn+hxJzlegXI6yhMM0Gy
o6Nu/dK7HriLKCQYBKHmx9ZSTibz/aqQ04l9TC8+Qa6HHXvlBGMd4zbYyao6APBKpCw/wDkgcec4
Ye3sXLU7BUd99KPPTaAb5l9cMGRAE9mdnSLh1EEsrvd/s8xibDmX9GC4Whh/N4e3dOhO95djjjF2
02HJmctz+qgUS1WyDhK7xYizKDIT8zMyBeU0MKRMtf7XcrXI/hZnubTQ4ks9xnScCbm6mjmxUnDF
O7UM/99UCr8jRUvzSFWOAgAsQrdlvzbuUXXoDGiBuXfTZ6tY9Gr3U0pcXG4gbmeaOj/0PEtOlYxH
fPk948e6MVYxSk4AZPWZ7zdkbjmd/CbvCFMLmhMRd+8JUqc2RmS0SiuE82Fsq/IkVekhbE419Hbq
JxkgFHPXgNvk9VN870NKXZHWc+32ShG8cqIYn9r1oljXOq2kDGcnOKlA47LNgC1wqkcLRnwCVs3x
UPkBhSW85M5uRzz5WEPwginaOARRTBELiUC6a0IRPkpK1ofQVWw4HUhtqtPNiTZIiF3KtPfj2W1o
yjz2Nz4jbPXy1K/yid++H1+W3OAP5RytXZq81pYtYimn0ErM7ZLAQaS0G6NSl1FXC1d5zaOzqXkW
lANsD+oG3N3KlZhwcZ9zTtf/7n686UKN9AuY36RAq4UZdJ5GHH7eclWbYufOJ1v5J6+8dxJi4R7Q
dgsDU6ub4EmVAaVE38ZR9ivzZ1o6LkooXoPtMZAOelRGrouN3ZMeYRQPbu+akfvedNLIuhNRipm1
j9axdmlPdUMLBMBjsMXdboZZdjVPdB6w+axbEK4XsyMVne5SmYFRX87BK9FcR5kFTvMb4kq4AJ2G
hFSuxnwLYci8YsLkdU8D6yeWTGLUILsTdDLacGoXFsIFrNZ3CPvioGzLqYgOZVI4yRT8OF6QqAa+
/fnTzWgLkMgG8fRjNMUUQuZfr8ZLsGXOIcaQJVPVvZHx7KfaHpgR4g3659CJfesw4wiR1L2fyVSl
rdi/lgH0Z4pvZ8HMSaAehjb2QtPcnhEAHcegiETez3w5Xd0c1lYSUvGG3zZPgsgy6tHOnIsh4/By
ef4y9xcRIjKP3P86V4IxE2qPs0ZxDxh1Xc024vaw97pimGYy/jPhkgO7fYoPhoq2LfNW7JivxL5W
bJScqfRdIuOwRCfhf0o7IKDd+xXYRqcViC+y/lU0p+2y3aFUkHUwuy5Hs5Dzg6ThPYKt4GCYm+3A
sJmqnWZSmvSDwj2s8O+h7q5l8cvfYD22PhwdOIql0/jgkkl0EL/wFzkFBjJG6OgM6d/ura3DtOh8
Ev7gkfjeJHRVA74WGTC7kWN18ic0U/Pmau2G6AJcgoAE9qZY/17Ur5gBeglH6KocdoVJ8hlD//wn
ISC85kjV+t7T0li/bAkQevf0TAm5OWAY0xNM4nNlUzpuWVQR4JYA49+oqAy+FTjrkePmMNTn1JmS
2T8bi3vv2THMAYymPO+yTP5IeqxklKsYWWQ+K104rW7cKET54msk9L0djt7yCNcVkG7/9oCuLiQo
wER/s6/B8JCmsVmuu3zg/i41RukdrA2+ZjDu41VRolNpIMcBqGN7yWv9hmppWL1efKmv0qekZWJl
DemB7cm/RSurga3VDm6iu+ro/S495ydI5BMcMGuL/dYRoAA2nf57oRnYwKn8R917fnIJPL9f8tXK
V1VI+/8GsW3OE9Y2icqNJTwmjfpaV6WmAvHY6bUuXpnjKsJidNnZHaAtGLl1WszYc9zZToFIabs7
mYK30Xd32do2caB7XM0Jq6oJYTG15imAN5Asii7t+JxszlgBK3egifLZ5g4gS1n7zNoTQ0uv5dJO
t+83UhJNHjx+tKTTjOBeSNOj1szz2SNry4eBy4I/2Pmu4rASCS3sRrivOBHdqxR9Dxf1xgnYfr3w
/2fCPnesOwuFM+T8k5lCvA4Hd5bFUhlAdRvR6a7EgkdPUNn9jhpmLptqRtl1wAuPTOuz+URSIHO+
a0Z+1vvUXWKmGKILB2DS0qpcLiNCu+L1+dHYMy080yyFcWRH62HZvfskhHH9+auISUVnavJLk/iP
3lLRCn+2HWnrumGnqWSB4QVR++CqDqFqUNpzmxUeBHqqhBvgSPvTJ9oQSUaFBzt2xoG11iDGnaLY
E43FT4358RAFBA2dG49KFf2Nneu7LOvtJrQwdUbuaKcwYZHZnbwDpF9qx0/jel0NDAhcxRlIn0Vv
fbQUaPBSWPg7JNxj88UCb96gGUH30F+InFqMoxjW2ECllc2/WVQZrtMPMMQNCJ+qI/KzbeQyuI4L
RVINAQn7hnuUwVNXidc2D0LQuT90qj4xga5d4Gu4usgrPDBRN1nQ6+cbv721UV5eKu3/iTetuksI
Uwj2y11g0Wl6irp+M1jMQ+hWWIEam4G6JtTh+j1upyHX8dGB5Qxq2MrzGF3dXaMshbCOW3GYPgZQ
kwq9Ww03SwiPlOWg9LYWguv0AYNkG9+skmmmSWX4ZuwI+A5Kj+wrvPr/xKLHYvAKJf26WJ6BV0Tg
YCHzWucPbCpKCkasrZ9zbPSX9DxGK/hj67ANWenz0kPuCOOiSGwrvflIaqfvxqnt8EdMEZJ6rUvw
RvdmlyzVorqvYkXihT0+QYE8s29t3KMXS57JoOUZUydTJnkbCZ3r3hfev8l5FcdZ02Kcp+EAOzra
79/gBBRoB6qsTaEMaBrCj1vlmwdAuxHHJgpd+upm5a+S5Rdo7JZfJ5FQ3EX/s/+Jcc+6i2Z2I2NP
Sl2SsRXzXZvG8lpk8dJ7UBH0dQPuK1ROMCuDIS2VzPK9WyNuWkvokeIrJ8QGBa5nMeOcU2t783p5
c+OUer+Vjg9YOI0Z2J9vN7tnK7i/kZzkB04iF1I/9vwJoLLPG4ONB0FwRKAZHYi9KMbGT7kUe4uC
4R7ubse9s3Yyk1bBUYHKdOf0Senn7o2HvKuOULUfeec+H/nCcC4t0Tzef7TnE6unzcn0TbgPvnGt
ZoqzhlyPK807YAXuhnqNgSbSfI6M9rHXn18EFfKwWuV2kB4hTw+Fv2BfWkCLyFXmu8HN3HgOFR2d
kZMIDojbUnAbHaRieJsQh+O7NTr7JsUE3J5a/4cfKVC7S6b666thnGxx6RZBH2wFSTE9uY8sGs14
IYrggV8qyrVcm41ZVMg7eF7R+mQPoGA+gpv7JgyPMjGAJ4GrZXlM2CC00k9Dccp46r+0OV83Xy5j
nMW9dyjoh4islxsg98d/4mIzjJGU6pRNNQyOyvHxLbdEPk2WsExpRh7Z0oGXptI8z+9lZAEZqlH4
uOi0jM1+An8wkaEZ6M7dxdYBtQQAKXokJW+nj9v+xTdsqQXh4+JUf/KZ6kN1o9xfdIi0MkGP14b+
POiVX954/VPgFkMKsYD30Ja4gXAUx/5KlillRTb8aYZZ3zkLR40im0eKW0O5H2L7ppr8dJlMcVxs
kQM2+O7519sSoKV2CyxexlGqjdlpLfF8u0gIL+4QtmwasCus1L4wtOHAdIHFez4nLOKCeyNngX2k
voUTweTfcWCvj1EjDstu3+OwCVeovIzx/NEWDEjYQMl0H5RV9+ubLvyuh/aqneIdK0o6etSrMD8/
J95l00DQWvPvYyTXBPCP5zbpHy2naQd5mkRbj44WHmH2Z/AFRs3WYjEPSAiY8Gm75jW6dO/j6ghn
0fKca6B5W0gXqMTSVCqOpwKB3ss2qYExbIdAUFEegl1aKMRCOqAoCshpz4C8xsQ+E+Jx//reJbjF
BqipLmH7zbwfEDASMzPluR0abQSAA7N+2SvQ8++hokYD7DYpYogPAFnVrfR2E7AtskDI0ljTZ+8D
FyfRPihIPglTeVwDbL2J/yt3yaRq5IEVbEq/JriJ8WvqZzkgXs35hJrujens77RLcoyA0p/mIlWk
Qv+rlgJkOOZZ95tyH5zH9cAjxUVqu84n7+admmDq1t4ItRv9blQIZ/2gquheVgStDHaAChKaryL/
teCE4emsAkAZD1hq4a+CB+YDK/tZiBB4n2/snzMKVkDt7danxyhZ+v0qqOWLb/gVWYIXJgSx3sw8
6m0/Gak0lB15QI/fOjDhxl3JxensTulWbgDmak3xeODWhtGksvCs5Az8BBBAtuqihi4wBsvRiT7u
DWdfdsxYS5WSDNMFGVzbbGiW32976Ttka0EHEHX3snJVIwT2M3Q7g3wSqK/ftMYsxuM+AOQL61uh
GkBHn4VQPkuV56tkVcPk4ykK8sigOTw/AZIlbEZ8Art6Dvpm4rewbPaaIw/H97edXofPYqyC6/GX
58JD4tgIRo2K5JD+NtBla2xtzZ2VixJJGm4d3g9WAaoQDoaaVO06bxeNJREVTAdycfhu+jgVdoJX
qbaV5GjWpaJEs4vMpVoO0F76BFwhFJDVdh2UpbrtU1zOKkX3VnpjDfGmUL3KY2BMG4b8P7bzuOpb
bXiDbchzu4ArShNiXuHO2tZxFrGzLSpMX3Hv5BsiiGUurBOpA7zwTH5BmDkO3eAcCH95By1jq8MG
BEuxK7//YozXZYUJ9wgIKRwTIl4/8Xx2VtkohN4mGuTmO9qjvfl2eivB79uT3/wndUlXts1uVc/7
VGzr32T3lV12LEQNSVANyidMYbSjkBK/rfgKaSKlYC1WIirPNGwODBdOv6VuLO2KvWIyVJQgppxd
jsLxQiDJkth/Hc4Jt6GczJviEkzLwzNJBOChWuMV8ttGAN9+9VHcjlh3TCm8hdvZeoWT8c/Cm9vq
8NK/ZvQ4Qadf1JARCxPGeFb8I8Ch9+lT4pt69VAhjr1HWb++xiSaNmWHihg/p/3A9DWTW/kzlFEM
LrncsdaiuPWRjHvAxiB4zUTa2WrWA1qKXL6Br+4iORVanEbAT4+btEm4vmMtLjC1n6u5NcGuOsUw
jtcCj3xhan4JLnj2EGfwHslAK9XtNavcJDcNnKheL5Kw+n1ZH5FztuzTSZnBFNRNUrrfirNj5aNQ
MO8G8glkdxozoqwLvs+nQEbvtfKDHExVK8bICYlTtFqDbaJsOL+pP4+5wYHy9UgT6UIzb8wUFjLP
H3Z4ut+SL5vWr7O5j8ZHipEbC/calMyKoXbLHHFaJknSD2nbR3rjdRlCKOonIuXJaNSdYEMYfpMR
SjqSPNLYCxWRyEA8VwednBjuM9dswkUGs4D/di//IPRt4Fsmm/+GNtBhsHJpFT6/3yq1KC++HBSr
7GfPYZ0GwSHhvEOZdPBqfONAlU28jl0LhPAJFxSq4xqtNNLzCdzF3JJLDTiVGgTLoGPV/ahsIEae
G3DNGgoevOtQDnoTQnm6Tzai7j0lbqXgW0o+nSTMC2mcUdVZ4SNbRAx/M9vlw+6q/7DV2Tz1/FTL
3BNfVinimbWs/xHatMo3aUVfpaSvqI4gZgsVzWhbInsPCf9tdAFkiU2ePq/bt7T4CeTDYSEeFaUs
qGoK+Acv4FCCeDVOsHno7rw+K+cXkR/tpvDHwRTtZx/nT4B0tmfuOKQCxU2wHaE5wUmT/oPVQX5A
I2RsGlah+EBw3ZPWMtnSJ0Rk+iITLn1UGEF1kPJkOeMUG6ke2iRKZFInFizooZJp8CzgnyPlsPfE
X4WpLLlerKjL4O7ei8HRePxP96qcX7dYRneJnaTI/+tRGX5pD+gma4zgsGF0emdkZo3CxJIMJVg0
7DDcfuP/l5YoG2/Rr5dtt2AxvwPbUdAKv1ngStlaCfM0z2oDreLBSOTfGVFLu+KPuuAVjafbKbmR
y/KkkHNZYJIdelPXA9J7fW5NJU23VbFzpP4ap5q0H9UVGDOEB5j4VPozIMfuUKRMCGyXC91ySpgp
qU0UNvyygno6Gh6GxdVdh1GZ8kwkd48ap/LJpF2LOc96R+gP3RA+VRyJx+VN9EIsSLocRQgejscB
DyxrHBDWZH4I5JI22IVTrtjdpJBHfl11DP/JbfUyJePoIer3wDdL5DOjten45F9TOtEtHBs0mz3r
DwYlFOPgLFeLrPUT2X0u+nqDveiVxuFsnYvdyfkGE0oKE9ZgmRdF4a+ugi4ycq19vYnrLuMCuzE9
C4tpn2J/1zzdjIs0gb1UoMJ8dHrwAH4OTtj+1g//YrM0AN8dWDm0mee308QaySOTlXafwvsb2+M/
Vox7NbL/GJtqlg/+bbHu11HYVuVjpyqvmr5mRN3EpBhKm3ueFuvEDUE/K5jRxjYSR9IVK7utls/u
5pyVMSfH4vxkDm246fQVOBMDHASQ1OT6NyY6iOGabJ+ULfo4tvbDJ+miGbqerFh6mmmCsjayV/MW
labXXiOPvdv15SYtIXxc2LlAS1pSgS/jq5xjlt/5I1+qF4wrUrO5PX3FgzfbL2dDiFlDMM8M/RsM
7K4b7VxyR922tlfLDhq6cJ0HOJZnA6F7csIGoytR6SYERYUiJd2JsF7Islv9wnU4DuIzu8slm6BD
lEjXWchuBt+HIiomPaTjtgx2/0MB+mWZQ2scSJXVFMbtADnjIJqwSfCDsvGldkLkvuXrWH1vqJgn
+e9xLQ0QO2GBoeiMxbHkUxn2BB7hIUbMpJAwrjVO2ep8RzvI6IT+kocfA7PNPb6DZTIy5Zz5qm7t
K/R2iO1W899CrOdIF4bg3w9Y4pdTt0ICE9pSLoyoC+8/Kri9eEiAFYlq4NtbvXVWk5rMGGXD1+1b
4dHyY0TxtI04f/TDjoGza+dPVF+amTNmLXtlCFAEbDUzW/+afA+arN2SdgpsvHzfnH2VMLu97KdK
5V/5kWfI5SjA8KvRfkvlakmlmokX/jUm5XkK7wTQMYdrUDDWQocsHK4K3nlHnLqhInCroOcgJ+YI
7pRlvIZJBogm3Q4cncxbyTTALbDT5tkDSqW1XGfbuISa8CZBqXbmcZpzQYBQqc+rUxAwDwbMjIOT
ODMSP5Qo1Ky85YmVhotKxiHwzxj6C8eOVh0SVqeUimMPyXEkEyIIcIYqXH1IFHf0EPvUebt/0ZLj
PPsfpl01LuJe3Uz6hRXbttXsw0PikFzROq1rDtX5dCo/SHOPSrIqaZ3BuhURdEnAaq8NIgiVrWuI
bcPFYCubaZUwE8JRt0RohMnR2A/Q6fOn0/OBi0FEsdPBO3uZIbOudKIUexQjrmLR2V0PYl0ECe9B
+j9hiCUi5IGHT9DJ5+ydnqVYigY116Urn42cvg6+NbKvnrUbNZME7x4Hwi8uvlLDu8WvPkAirsD6
z+JAV91euN0KXSe5F214GIIBQ8YlulxGIdjxNsIRc0zK2/GGrYQ6jpbDin0UJgljKVo/OsGAwS/O
k54Ma86xaGI7QvPyfnXHglmJZXJ09hKXvt0vZ9Vc+gLpYe4Ra6kAX5TL+njngqGp8Ol6bpzV3lHa
c4oxSJjnCjhn80fwx4w9RPsdVTFnlu7Jikxl6SzjiQwAlYFRVOnyz6EOaaa7p1YAluBa0Oa1fuJP
Jsw/8PAAkI7NbkwAPf79Dmoq042FGyW1x6X0P2jWD1GXldc5D9ocPOSouCzt25PDq/j38FXVdbpZ
cZX4/+UfP+1Q0SE9xlyKCgEFqUocOyKQbjiTdG1ET85Wl+r4QjBfY7k0WH2Myt6lyQ0Au7nePR5G
WpalNXydJlXWgIHJjjylV94oe9gZpw9V4+eUUkt9zSHZxFzWS3dn5lA98DgxdPaAwlnitxw07whB
nQfyGfQQvOgOGasB/sLJM8NuIGn+McQKasClkirzXQOd0SVvXoCfXBQowzMwJnroB5lPUpBntIA1
3qGFW2noxZMCzZRSTFfZhuOajfmIpkwZXATfHeHYpCL3MEVYwI/hRF2Mp9SvovO5L4YnosP9a7ht
VHBQak4n3b3EnMXk124bBhTNc0VCggUSel/qmUzKLklSn86F2/ceIH2X55LDsCQlWJQ7FXADyG0r
b1WqKzX2zt94LOaUF9cmuS4hUHAarHyqlM0j9EMN4ST4i6CMhUhn+SZPLasJ9o+9xb+tTDSHkMQM
hqE6v4rOI3LnJ2pVtt9RDMpIe/Z281VPAjkgG1sdidWDBzc8Vfi9HeZtcACGKFQsaR82nL1EBnxX
NHKQcw7Slsus8hYDo2nforG8a0e0D8k96kvZRJ5PaCLoi+rlIIh3b3H/rhseA2bG+VHi6Gs3/Pom
hijtUPc1BOxXfIxvqPbQoZDpMEjYISxxoyF4n1RJbvMwRZTAgonA+vpjdy0b2NauFGpdTQWXX4yO
i2FT4dZB7ll3QQ7NetFRfgazTAO6E5GD5vhBhxAUJu8IVxHIM3aIekmY2CWeaaewPtf9wtTM73a4
g1u1JiA3p88QQEezCnvdJntD34uZh3sWzsUTjeI+5iBPsHENMoAXkH9CTS1IffnSNAaDHL3Mi3nE
nhT6KAj90HdZxpaBKgi0mM1HCqvTwKUiCklG5z8uetH+9qrhpVZef7NGfR//xkdYBIGT9UXdpvM+
HM8MjWvCgXdaflNopUd4A721O6NJG6Bx65VafG6tMgx5sa8485D/GBg+xBkMiNHb8Ri2/UPcKlb2
WoMSH2hZjfObml3fOBf4zFBoMB3YZVirERsUDL+ofWqtC2bRD7FH3TS7OfhDfqTodWnlegeTa+1O
a4i1vj1RwDDDQmRNtnf3QJ5cq1Q/1BoXaY1NPH0+/OFEtQd9L7v3Nb9ocNn1PZ04VpaeWx02/qmF
Gbaa7lYsTj0Z0hlZm4qPsdNRBVNHx5Ys5PNdoflYHtisfDkTFh2nrXSIoF57UUqLo0vYMV+Pi+Zq
ZAvvXiND4ZxZQAqC6QvfwW+nWM0HSQbqJ5jhYxI54sxU/W5W4WLh8DzY4ET+i79w5pSYdiaSDjj+
2IvxnAdEbhxSPDP80ndvuh/Za8GxmR8V+qcruAwaAEErLFWXN8uT5aPhi4rq6AD51S97lhLQaOC+
o+BzSILM7IuFWbrhmUfMd4zgFMuW1hDGNRdaA3p6O9tqr2WjljdPk97dDOWsgtXsqYqdPjDAUADA
kyXZEdNaRYW10vSYLn1t+AZv54ERkRtQ/QcFGSdJv6gvMfm6Zr86qBJuQKKFtjx8c6z4hxQPj782
nul86gnAdReOVNbuciQP/7N0ABY+FBbJZ+BR/M/v0bX0FTqZPmhRqPAQuu5tPZcdLGfnb2CINmEH
vgPWgrdyeEJbrHgFYMUJGQt5TOp6CUh1ygSxuD2UJ0b9fIk13EFxFZXcAvCK+voQRisnMDxp5A1l
brrh9uOpfb8K846zy+h6pdaXzY1w7JMPyEXZ7xB+sViq5beMATjG1FqnWvHJE2X4i/w9hV0xHCqc
s+NmWfSBtcaGSfKZoIEjhIOLDmYyemBmNRY+h0PDVZWMfaOcJOCgo75U/UXXvroZvazLh/WXQvWw
IZhh5e1Hi1QpkHqWg2L+gdMnWPUd4OHqcJg4QqTx7BWTVO+BrzE2CsT3q3S+jyxqcLwvQzpo7pC/
seTWNzdYHUI7tRZ0NXZlb4Bbmq8U7URH6hPplckUYno5/TpKZgmzLaJuO+463Bo/j3SMMVB8e1DZ
hPyMVndFAhgKNJYWiRxOcIFo5NVE5txNN0MCefjDf8KsaVl1djRx4ToFj/r2qhdN6Z9IZvltXiFD
y90pnWJYJiej/R00GFsKXQ+S3MNCp6VPU4yO+z94e3bCzNWqlb/kLaPDQMwQe1j0GGiHhKxaCRh9
m8Ab/2aLH3tmgdT92Msbl7j8/Kshcu71ESuRV1RSDL48V08Snvqv4dandJ32qiQVbmt7AF8mp5q1
gX7Kegs7hAV3chro7Z2rQXvBoL62AbdR1cGsUf9uoaHkjkqL8+Vv9pYDC6hzl9FYUh+SUhXCinWm
969p457htrwtpXaTNTZb4IFTX2TBdAxGUkF7aNSp/wQo4Xn2G6U60+SrImSEAesIgbtKCYafUeHs
tTyk/P5uSGyoE2GHODKhDVrlYtTeiCXdj48h/vzN1Kopi5pgPx3+i4h0ukKFCdZRF6xn9Ew2qQCg
GZXfk7V5+NJf+ddQNPTwhjo6iej35FZbDWilg3FX2bF3y7av0XdkPJAf95goExBhxfkqR8y0e9MI
770adTxc60AQ7OCFqefF59z2T4IFyQq8srzZ6myuk6P1XvWpNPyTWbPnI0BEMIwueF8z50FEfSxn
5QUNTmqvrfUtAL1xBnNK4JyF73NPY4OeW4T3YT+94SrCO9P9WXm5WV0AxMo2pO2mnkBiJRRt6Ctz
3pyrZybYEGVjyU+RHRJKn3PrPsMLAJxuK3Q2KNEx9afcIBA7MlEe8R0K9Ysuf2WOxNTdETZ/uXNr
rOiRL1w4C2gVGTrr/tQojuGVJqIb9HIhUphoY5+HflJvyJ1wmZX7VCtWbm/5scvREFOyFDvZATOk
bef2aHuhxGZpQBCaD6cGXVzd+gT3Gaza4BQYLxr12CI4Pw46XP0atgYfDCaoh+ZNO5leLIoQpGZA
oVx8nfI9VoqS5GF5OtXlmGvUyzBOGUC8pNq0bTFmo+OfAwa6Wfnw5OEywSfzB6DTWsYodfcXCLZj
vVQX5SRVJMdjIcIq5ryBoiRwiM9f582bLmTR5gPo6vAQ3INgDqrZ7db/SfmcYVApxZIdcCyiGhfB
GgSikcFV5VM7rP+639Oyl4Dtq+djwNGwPS6877MWu70sPxIYAZVYDTipZ5NSyboOkl1r2dKvc2YG
s/7xLQdW5nvXcxnLwuPDTcGLzxVKjDj9mFnbQaHveL5tpQZJjD44oJhiJ1ufr1CfW9zxM8bRwDxr
7uIg11F0U+p95ziiTTsTxx/WbGDC6E7xXiirJbAmT8G0MUKJDeN9RqHdQMAnOiWn1IOLRhkQCcQy
/H8j76IMmYUKonvuMfIKktVzpFzn3KsSUANQvACgrOklvst5Z+a2ERd5peo4qLYGrsxq8FYfnwOq
mpCe5clJD7Qv7qN23vnXysQ4A71WMBr4Al0hfWnkdsazY/64vvnh9Z3nh0gvyOrADNqRhTnOo0ZC
cbF00tGiQkIAB/eW5S0yLDCOyLb4C1s+cS8Ls181xiogOR9TV00/aq3nM7gZmlnNQxuWxezE8sMm
4IlnT5LXY9HmISnJ27cAqderYBg69XnUs+ob1SKD3XRSe2zznTdHnTXtNqqytfgN3Fyq5mP3Yt/P
PO2FmkI41qa6xd7BY6EdbLEyyVp8ey+A3RpCMgchI5GxHHFo5JNocTmIpC1RpSadeBdA4YrP2nyU
6zQgGagsLEhk3PWrPhcsfGsYwz37BYwXPfOsXDOTRd4FHWaZfV/4hSCf+vC7Y/qDM6Osm8nGqFbe
gQDI2kOdQHmrK24zyhWIVCMo/gbLv3s6mUVNj0u5zkM6ssC/QY7Crt/YQjcVsjga7ipIcpkxEvk4
RRmK1ibpn4PFD4HJe4btj3kpjg1IvMxJ+0MVvss8/wioT+GklS3mTJAHxuTQuXbawTQTmIsUUz5N
8EvWmAMDyjagUFTL0ugOW3K5458BApG8kFOaK62Dfh4sT/I1uaWE+XV7SRCCGqz+jzjgEyvpEEAx
cw7o8jRMZNGdB4dqOuS8/vP1zI5tnQvPTW0RTbbuFd9B9USFKRd8NrM0k1jmMXNA/0Ml0rPelFg0
LxMjd7Y9A1Yfl/5dVkGKMsBtcxRL0jaXXUjHW36tu19Lb9H2xLwcFkxHx6cXnJb1WXfkhYRXFgjV
KytDBuzKTPBD740E/1A7x0oWMe+iITisgXAOB8dLSDu1uZrTKjw4c7tmXNrAPx7a1UtlIjhavyna
l3hlyr7A8xKM2aA3yOyNJwkrIi9xdonxbEDvjums1kvK1lRAUiJrB9ngNvM7kllMknRQ8F9OM6nq
RnPrgnrDAjAJ+cyTiMVHl2bQQ37HzvgGRqYxMBS6nSkAFELAsSJEACzjJjg839VY1bVkrfmULvkH
s0bAqT/w011TxKXMY8e+rtYiDDWFdqTuYtnjiVg1g0WYLcke5xkYjp0epRi0TSNPHkmbRaptxKb8
6Sax3oZSyZ8rYG9gxrVJ6sITpxxhc+zDWgjjhQ1/4c7OkjCXJlBTFv6rTJKQp5FokhMVfKsbXYzb
kyYbpohlnk3qBoKL5RoYRBWfgOsEmY9SfUxR3OvV3vYuIv4c6K92mlqDSaum6hLx8PFyxbG0CkLY
ybhxt4AYH6CnH7qhvxkEdksdpEgC7bs+qnLsMjWXyjsCiW+SozSGFsXDFQM3/d7qJycWpzxmGfDL
rIcG1zzEpCRnWAkvDyQcYc4CqJplfM0UW/+a2+Oi9pzS2vrFkMl+NEUvXhKSQxoeo6Qkf+1k2tB/
ZHAU3tMz4B3mwgIIqNbzEV0Dg8RkrwcjFU+jqc5QIsz9RqL/BHzmzPLKAWs0YYnWCUOU91gVbx8A
Qycd7HwT5S964EYH/X1ObApGKtZjrRZ+NTQ2iq+7JH+jMjERltcEwGGsRWIT3VNUfcEIp+KS4roX
Dri2b6tQCdif+UAgZAk732t0Hdt7ZBYES3hAFF/wumm1m3iNFphu0AfOiLHnCsqPORk7Rw0wka81
94PWiBYHP6HsgGip5rbhO5teBTlhHn0XJKYM0thW2EMwVDg/4LjkvKRYP/3SLcXf2IuQlnoGbg0b
02TEVbUsrmf9pfSnlKbF4p3Sit2Mq4PDQUje/MMeNYbltblW/bJBDyi5evsiVcbOOZ89m9tjIn5r
0XsNvv4DoROLEJeRiHztlFGMbz3QGubJMv+0bk7X83jr85cJ48axjRrzqwWK4NjtdI6RNhgElmex
HlymREiu3WzIoL37PBWswUxoFXiPKBxLYBw/UaUf/myle0WwHMhstw51T4ZWIBo09mdhKrVckA0E
TORR/VxyBAEzFh371uuAeJ7bR5bPvUwcxSCelImRXt4X/zwGRXLGtFpP0iR+pHStS3BCcOcYsW3L
+fCvCr2g2SGEOWcsbIFI15rCc4RDyuGb86ZxUxpolazk8v0RepmyQO3YcJsIV0BSTRjsNTZcHScr
AybHIbLr1Y5GkqN8bATaplz6ySH//Qtu6OP/HBdpfyBUjBNwY0pVPKgPSOVM8Xw4CY3I4rsorysM
cIEsKIg53os8mluoLW5dIpvO3/Wv4ojzGoHLV7dUVHFtd30LWlJol73E/4GW9vp2V+5ShEQkLUH2
m7zvSh/X8m10a6SvEzvWLlmIR/S9QEqvbftWAVtWZvobBta+C7ZkCvMN1MyFILMHrOWclqHNKqp1
Yrar5LhBIOoBG/7j/STuCmGyBVWP1DhPKIbzjehT6p6VYsl9lir5XTbCzzo581SbvEMEUtv6YVtJ
XXsCK8YoIySj0LS1Ih2Jao2vkOIOsFjfBDMf3kcKLL+yrqN5UezM1tiWexYO4ipchL9lVJc/PWXv
+GeCYWxmnJWLHaTu7v68APXzHYD6SEkT+F4+ThkQ0NIIUZwFvU+iL8ef/BSLCFYbuDW4spZoZynr
2T3FxfXuqPihmRfiAHa2FQUmQYJYyUt8H0GjY++TWcC2jwUW1DkyuMxflsEXat/YW+AW+OU+R/lO
6Wreewj+KJtbc9NygIui78FKaXVSJXCEjq+I4B25om3EZ5XGqjMsAjTHw/qZtJiRJPW3i2DmBF4Q
tjBmpPcf5BMGPyx+Da5f1Iiyrvl1gXClqmGVp2A2a7PyoIbO42U1arOmtpC8APzQWnfNA2hMKhHD
ZVG1uOHNpdE4ZbKxEn3kHtQTRrv0nahk+xtB96KWH31RnwvDQ2gYy08k7xFtwscmdRc6etY/zqsP
NmedQeA0Toxub35N5O4fnufQOQqgiFbiG2TW+10EpwU0GfQpAsnu5o4Wesj+YU+KM6JiR8FuQdLe
RBLDqqgha/9S+P+FXyZh4qSQEktkgEUD+QtzpHH/TNwELD5M9rZou4DLuGc0WI9B3DjfAwKl9Qel
n7KPb5l7F9PnGLRwoWlU+x8/nZmBOvMNlQDtCySauxdXHDTvIHqMO0xjQz/4szr6SAVIAwZOOZQx
TcKY8NrNxG4bX6mnmxg8qMXvMADD3uujpCP5Mhqfjf4vKOLmGu+2sYNLOAj4a4uMW9UCCKJDw/Hi
nI24H0/jOZbkml+XzxeT8Ud70gPb80txR4FnW1U+XjE2rN3q13NvlHpn8Q4zVW0LjdoiwlP14BEO
WPlw9ON827HjYig4np3bvabIleHeqi8ClIeVYRIzD3PuQWCqI0UrOIPu1EQsM+nW7qBqRWPtJEqs
UirB8B0IgaytMJO88JbaBaJMUCr61UBxg2i4pJxgIMiHHo//mwDo2yvGNSUp8/BOr7CDCs0acSOK
aWGreHH9Xz4j3ge9VT6d9XpWxxn85TLJyXZhaCGndzEA8/lBK/r8liDnfCoE+bBDALFgVBUSBP6O
BZLF5djBDrxqAlnPTrmQ0P3Mwd/rRuPvwR8h59YCZH4BK67F7ra59ChSvjq3cZwiksg+IGfpEp3s
arhPRFPW+60+ORo0zbnwrvRYuni5MXT4Kaij24XTB0NMm5gZlLuI8XV6haL80NynG8qFONUPtARY
yeQH0m5TBrdXS/YgNyqVIc+CeHo7zz1eD3IBFCyqNXyUtnUa1/FA6Ot0UMAb3NKZhM+lgkfztqc9
0nQ+ThE1m6DooClpXIem1YRjaAZnxNIsLfzMPh+Ag/buw86R/w9IenBCOuglzadF9nJJe5zewnsj
7gkRWjqi+gv6zJCtfclRhsTMojqhllDrYwzKuGhuTTS7SOrZC+r2RC1ZoZAQZkYfJystdf0JN8bx
2P/GkiFzPQX121guDgUdmUEmU5Fl1J8VJmXexdXip0VYkr/XYz6BFtaJ/HyKilQ+3AzT7Snta1H3
kKZo2iYkNrNzD42Op9xipMT7my5qGaXAV4sZmOfo/bH7z+KtbfVPt6z3XlYciCiMeMKsBvXfDNvR
sbjKLKdL72lZlZBejfkeWdt/2rOnIaaJMb3/608LJ2lpsw88bR959stQoC7SgpCk7CoB+jGqDhyu
5LtoVtHGNhKAlCYyWFv8a5B0WSuYpaD9dQfZa9KnzhqXgWjtNi5W35h47AqzvH6vpeaElF4AYpvJ
Bt5dJUgRavioNYSmMIiZUr51acqRri1pcEPgI6uhndwf5yCMkNLgoUpbxigUv0ZlOzIT6LeFQFen
QpuhJq0UfBnyU6+dSxS+KoP3FePrJHc4FtSLcGbKYZ7cHU4CBad8E53wZtupNbr4lvIS05jHHF04
Xwgc3S4iCrqeWdFDqcvjCCEcXc0mwf8UlwK5QNZmJOPPgiy9Q2yWyjMNJx/rR+Xiye4GHE7oE1lq
BokEXyO42l6RWmLOnE5LUmMOzHUXp5axtaKksW3tN7R+ZojjuE9BB1by/Vbuns7sMGqU5bPuIz5m
LYUz1r7gs66BP28eEQCLaE+oJbiP9I1h35GmozmYEhirxY9Wlfws1l4NKkl+PQkqlI08Yd00/5nz
c15PthGoUMLfEmgELInwToGno/rASnC7fc8U5lrqzyCE2kP+4IjrPasX32tlt1s3Wypnfnn61bFp
6fjvxIoNHovbv19fE00d5PFxurWcKN9Ix2gH2rMEXBeE4BjQUul8+aVHnanFxPfnNtvXVJ5fK+Za
NcGSJMkVDLr+JdEz2soaztK0DOHQPuSmyyPEEUZtYgU751kx9/G7C+YqvoNUi7ZJmjKJ/o8B+hK2
yLLC2cFhUd/YQXuYYmJfFfx8e9t7gwYX3GJM/2KiYIiFwTAEMcDXQqg8OIz+YKu9ev289C/cNct7
QEWojxrv+DURGsnt5+gC/4OL1oDQWQA3bZJZsMtHWMTU69RtA94JDVXdZVerkSK0AVsqMTbuBfP6
1jT4uOTRWNq7K1k6W9VRpHqu3fVTx2MaayFzuRsm8qZEnrzVFH6PgtC2aX8UgTNr8sackX5d3I2w
nmUTP2nCT+rwpbxx4u5oUvu4ji0thZcwNdCCTZkZv+VnfhhLs1hfFQwlmkZly/Jg4e1LQ7gJm410
i1XYHzPnYOls5MXqVi99BxBWBWt6S+oUf4q63n52qriX9wc07l1Trw/XEviA4H1sJZDA9MMNUpSQ
ydSA2X4Ix5MqKUshhEFih7xXjUGvyPvrKxZ9MN7KLD5zk8OmB275JhMrKhFkJ/KC5qhNZqbRCNlo
ihPTEeD2fCDkkNlCkLRfOzmnK1XIGr1T6koXgw5gGXJnCFQPHlzC1fUtF7bkhvfBwJeW7b9ikpXw
cV1paNuKyUq/xqiI1h3F3muhm599UgWaROu2ciNRwHozXvEWw6xdLf7e+bWqm3LdmYH/g86m5i9/
+USnPwO0rGtX2fRzDm5KjlhHeyzOl4aY4zlPzXfWo3RvVN7R4Cvs99rs3l5MZ/Cit2w410Tch+AS
MWz3tUPYJjRW5RV84RxQbErSEtF++ppQis66BuiE3C1fVX19gMfr4+LZTne4YhWkuZU9hCkBgycL
umIaa0gSLX4Icae8hxlNOIpwZOp69lhzIRm6UFodYql50ueab9tGEHl1SThyzvbHPAk4UQHrQmIC
ozYSsA4Cm+3Wz06GaDudlL4SwTBK8xdSYOJPnncIMlJ8VgncFmafqKbmHYlEGbIlEHNBw3iJyH2N
xR/suanyxS2cFjgokfDAViyvBq+FvLHcN/mDuAdmyg1d9pyQnp45MpKCMRh8Pcob2tF5QScos9Ou
5nBnMXhe9/ngqPveXIQlLKiTh9wLCv/wqQE7LxTcAEcPVnBB6/1TzMwGvziQocPNZwTmPD1KXWIS
oDjDYRoENlgphsPwVdS1tjGeAQF4E/fUM3+3mcJzR9pbIWCBvaQO+qCeSJSeS3HbAkukFlktsjj7
SvBE4/wpB55mUpG8/af3a1CwVlEIaa4KYjHiCgWusXC8coaSBKguo0BqC+SY9mGhDdphpESqHJn5
SUaO1eBBh11O6BRw9pQytLNuoaaBFAHuX4uKFMZW0vwnD7i6WlL2JeaLRk5Re2zZGcEf2Oe9JEYC
qb9u7N6cNDRtEQJj/yRl4z+BWLc6ZHFWwgVYVGGV/Lx5rlNtupCdXwUTGpcbtQP+Cpy/8UsR2EFG
yEd0G4m5NZydb3XlJJD6fcDUwOKq9P37juPMJc5NOC4cI7CCzUsOQkhaUTPdJKnhXuP3sRu8HiON
EGSGE97N1ZN33IeDItJQABT8VFFiE+KHe5kS3JTmlFfdgHxuT9zTfOChEo9Z/udESWLJw2YFj/js
UusJwjpvDbH+Z+nSPE+ArgLw0NvBORD3ooGjL5PZw6m0NQCW1ablT1MVRwjLZdN0lHaaC1uHx0SA
SEXkEI6QqzzfMkwOazL7rM+0ALAJzq6yCO3rejwE2SYwtewTRCb79kFKGZhKMeyjaMowDmxZsh/j
csruoaFdoGIMgCsvBbjN2Hl1TyhTZ54rHZZKSFjaZONglVUg4QKgAbGq3TTnWuT00tzse6hZ69hp
7uIPatT66qamtThBI3ZO3ODKNfJbwcIiaaEo8/K6d/uqPHNa+aTSnRfFT71Q+wwFONlbmT6c0ooT
kTI8jfdYhFjYbVodV9eLLv7I5BzkOybzUot4ewpzH44kB/7qby/wDHn69zUKebkf3lKkx1pEOdtR
5XiCMu6sA6Rf7me+W+PajA89vkAMsFw5odEh1JtwhY0PvxA7qT7umhFLjeHbi55V/+QIIwqQYVh1
xec3AvfsIHWQ6gobRA/UK9DVTtlUUCDbNuy6Y+i6BXUrHD2Z+U57baqVUjViHEhTpHPVNhbIfn4Z
0lzy9lDevangWVgWLQKgnNA8Cp11bFyhfRbLbj4TaflOdpOTwa5vUrb7p7Sk4P6rKFAtVtdPkHe2
svLM5HY1tDswfAjuAC9LmQky9MpI+GkoZj8H2UIMvnSPVa3N7QNELJJpiMwcpQcS9FrmMcwdAHj4
/FL2g2UJj3oXGJoGDhlQmLtHyidLyVEhdPjIXm0siolgjEOsi8EHzyzLD8FJG+53xs0CvdbC/98S
NnGSLg+RRKG2ResweXy60L9mrkIPPb0A8b92YgiuNMD0plESvBV7sgeUiDCGFNOw9x0BSWQGoR7m
ZIg+KiiR7S29lQwej0XQyz6yGEB5Ed7DiWOgdyzQznuqdTx32/fVYPkqFPJ2Lt6H4SGWC+rb3fkv
gPUmNWOMbZ2iLuWh11OArOwolzIXsILsHwF+12WNymmcCBLknOmLzSMgF2zC7v4HhacVxsYrk8D2
Uldvs3agHBZKWzR7hJ3yjEyw69U8iNhSLDtud7OJubGzHaMZrh77uNDuNKCPfQUXk9pP4XgFMpkN
z/bIXsDL8ipDn68G+6vByMFYkBGzC4/3IJhLcIafVfCtoGIl4t/cEgr08R6ETI28T5ozJvP5+Ju1
9M8iVzq6D281Q13KxyXlHtiZyyjmm4X5+B53XIM1Tt0+xaFXK20+p6Vk/ER6KTdWld8TlUg1Q9E9
rrM1rkbaiYCcH5CZlCs8Ryp9QamjwrTKhJHWdKh8NDRTfdiINycXIICOo5AkjYaw4/KI/14OJ+iP
kRMZQiTJu7YRqGjFr2C+eDit/KiAkrhh+e/QR4gPVJchDQA33t1T8hqAztc6zLrLx4iJ1ACcx8WS
5d1W0/h7DArx8JgUkEOpMgLuiWm3x4LY/zTPhrmapXspCXcmx/GPB7qMofMfE6FXeREZo05G1Kgs
Bv/9rktt/P72N2DPgmrPoT59xxHt+a1nxdmdjFuOLJ/71uK4JPSACLegBxyzIfqfaodxsP6TDwpT
9LwNWwYzquWrj8GzD3nvnwo3DMJ4Q2tmmXaNKRmiayWynSbqugEtLTyoqOdtrC3Pz4oVrDbYEU3+
cIgMVO2cigP0AhSpTsC4TIwTmdMmpXrG1j7qfJozr9pZ2Pn1KRkFClWfcwclKXOsjvG3D6WKRJod
ktazfz5BXzFKwE/HoHjE+DLcsICTEziUBgPHF1fz4N0yZe4IRYml/D7KtcXpD8gp6xfq2aSu+3nv
SBLK8lGz9Ew0dCq37aEKcGg7zrUryF5txN7gsfv9DbhN7txhhUa5w3MDbBCArAFklu6bLFv2MVBm
ePrlodp+BhhjISHVJ0Clsja6PR576vlaVMVjJhKhr3+37XYXLoeIk+aUj1zNpRlXFfW5iYF0g0C+
pORK60ObLn1Crzl1YHv3MEYCew9V5IitPYCPQRa5Bj2IZit1AyjIHJvmM/vbk9zrkc4tL1RZ1Ycr
vYDG35lSCieLmS37S0Ic8R6UwDXf/dfxIu6BfsIG7Gi+rUO3DtxMXW6JcUA0iNkGSzVFvyjZEzRn
MJi49YTHpMl7VooplRtPcJ/F0MgTY16NFUZp48scnaMt7l0V91yGfqN7DmnSokash4LmzvBu9Uze
zTyKTyJ1ciW8BEGFjE78WFqoKruFNztLFcu8XYDN4PDGTP43cT80zBmiF3VKiy4vBTh+pOQxRY4B
FnTmHdvsadHWKwmxcIi5i+zVlJ6KXKjmtfj83KohbrONiWTKF5hW+y0jzf7tFEYlHFyjdWBgijnl
7gCzWiVrP8sh9yiaor0xJKYUO3UqZYbs8H0yRDsEV6IiGRPsqL7u5xZnlSUVMgxQxC+S+/CgEqTK
nJ5l20cItcocB0+2MuCiyRE40SAd37YHvPrLnPHivR/MFbi6momqqjA5ZSjrg0rzUdH6ciapUxrv
QYceK3ItGgAU/RDMzNjHmi2cgV3HMPxkvbtMzskexmFvIbOVwbyBMlVt15tRxgk+vrr9yBykXcIo
A96wvMLVFU00l6NkG/jEVMwT6xdziXcroNPOrymIfTIicTkYAJgpDN8eWtAVn02WRzYgPhBh7Tay
Y4GWD2vD8IcmM5sLEGOA4Q7dtEwuRtt6UackilRSlU4L5d1d2Uqpy7s/pKe8Cg+hlAl+c7xW12N6
wroAk8HF0fmKmvcI9irdFRt4c4EwIHxodvpm45w5LrrJf0ta2DHj6GmXv8WVLTQjeeMp2ytvCo99
37ydbJ/eTtxkpzQr+vENhdG5rUcCvF8VY8CL0eRmy/vf+6Dw7yT4RC6fllKOeMXZNdeg0KhpccbQ
CJt3D+CJ1KFdh8JcBIHct+crQsXIE+yMaY5mFxzyqE707xPohyCVkDqPWf+shvChcYVsKyujFDmP
F/qeKKbQi+0oIbJKb/chUQe4Jns22VlKUvhDm7espLHsYR1phn8X6zfaCIqxLElUBcZKJwcEgIN7
MpBZYsOxkKzraVs1PmhvYbQok3ToMlkxg/DLtpVExZuhpPcd1Nl7LebDx1vWxvzY2SFE7sTBRfeb
SHxdYKPRdo1o8yiGq+bzt68RILSQmBng3QpdkCHWP2Jy49KytNe8SHKwTwaheVsfjYYOtx51XWFn
CD1Ou4T+SSLiLKwlU+foYUHFcrbhzfhIDKdu9sTJyCfF7BxYy2Q1xvl4egbcnnv/KR/pMzRNid+S
Pcj6Wv59MppqwFdr2sjM+pP935GGaBv/AY5Gxlic+3Bw7ycQUNEaw6aPEucm+ZHuD3YzrF/JsHKq
txVATL2c9xtcXknZs9gA/gJ9z6cmLiHlOAsxDLsoIlhbI/jiWOwB29RLxcx2QBMyFv4pzDRl7w1L
jneLRvxByV73O2dsNjisfmvaRKP396otCPC/TikghT7goXzlrSWMzwUnj96RHp11Vvgo+yaqq9E9
VUOU1HSZp3tt0Rwy6Jxan2rN/frCmtVwghEsAFbI5KXjmG2iPuQ3+t4kA+moqGnN2MwooEUf32Vl
qu4KxzxajnWt1N0k3W8cyiSMXag/6eYd82q3mvmWduxy7YLiZwJWMSnZGqSozIEeo9HhiskNb/qP
kHp2MIlVcY9KUIPdQW2r0vTiFUTSV3bPsZBI2qwWnF9n+Vq4RDdVRCo2fNlF0+4p+HmCOjnQlGn0
4tkpAEtnkarvYeFFk1ToDCTCG4rOr5qjdRQ9YV4kOgx35gpHkjP4BVvukjer7nmz3vHEEKRrheSA
avcCgW4sl1fb/l9qFstfYUzX9PQwYYvZDnuCPLlRcQXK/Xm7Z4gU4hZ5GzB0//8zH0EcUBWP14G5
phuzHgKN3aHsRmi9oIL657zp/MIa7VCtmZ+w8Dh0mBbNG0iKP7z2UGuOmVsWYcDPXSmW54/+dE3S
xbU2dH4aWqWokdZ00VNJUJVSlk5KiGwBS64Vh+GW6P2pO0EU3HmwVP6snEjB4svHnZoEeQO735YA
UNYUHWUo2hsE5tKnXQUGBSbzSpBuU5WJeVnraOqdj+HhvKKqiqy7Booz5Q1/kOnfmkXaf+Owz14z
sSDh3wKPMp92iXSywCjxQJqUoJjy6hpgqyM5HKs0ztIjBEG1Q9TKC2iEq0q85WT5tkYthkKoNYfg
HUboLWYdY5FyoqyIUIfQLq19C2qVSKTuGNB9brACDGaA6fL9K9byWL4+gQEW0Oo0JFTObw5mnbr1
ug8cMs1rCsoAeS5Ej2MaoQ4z8aao2GIUqc1uTDfWIw1SY/AmhUXqNPWY3l4UhnGAYfw3lAcKnGzy
1ANUlwXpCeaWhH9IT7k1d0pRgOJ93W7HwMghpjn1mYvbd8/lpd+CBr3lz5a/hYGQClYwIZFmuaqF
nWqa3nTkoG3/khj0Q5/SQ2NSUz2Na3kL6AyOSjt2FwjzmOZZy/8NADD8Hdm/mcFuvLVc6+wgc7ot
nGg3ny+1PYbxUsTBtZJGzpKTID8IE1zR95CZ1V7OcazvGu/R7ptcODUgtQX4R8fw6/U0d6CkEw0A
InoDQ/C+TqaM1g9mNvWTW4Nyl7CJR2wYE3Q9nfe2rTphmivkM3xze1dk19dpuHtF3aVkpz0ipEiu
Ur2hmfRTgH+7/I+76CrkKUjQJxJkrTFRomAr/VLn1/m+RKDJ8rfSjajVGJqpy6hNU0CPhAU8tOpY
dOjDWOtaFUByoX2yDGZsX5JwD5EB9JtgGN4jK7phtUn5hTxmV+dAP47iwIkZcOH2BIcoQoyPq2a/
8iDOemBCGguUoK3BBDBCs+lRuki20CCIKrcq3q+x0tLAn6LyeypjsLjJWeO+aDgqUHI6+epVYmdW
8bXQZ+0gh1BcKAVBk1g7MrPk/1mXigbavATLembITPTrkyasR7QbPuaGjxnax7CeaD5TiGIyaoj6
ulW2imgIZex5IEqeHQfmmzqOUZTr5c2kAYMaVK5z2XBB0qnoEUQ9iKjEj4UMOfm5Pkh4DFxDu0lh
Lb2l92kRxKK4X00mXhRTT0qMxqpvVzo7azUqvcuhsiNMT/0zN/eRdrdgoUKlvBIMFY0pJY6fKoOs
v1wEGEFtbj4T1E7nPrFINL0hnxPOUJpvKSYkNFjYCzUiuOgrsHTwnI9Z0B9W7vnlxb7Lfu4F3qGt
LLKcU/UixRMN4DCd/19KsBa0PEWF40QsiF9Gzu6JsjlyUHjj4o37ekN53SRYtNqR7UlSGOEciG0/
xhuY3EJqrSn2RA7EViPmjIL87L5EyAzaWCbRwceptagEUhTQ0UTkRnatSWnlPpls+y81GIQ0TXvj
W+5XAKuqlybHUbHlCWxxdx54/OEYwJH3tuneSy/eh6OkCTcyOXu+/HSuRhM8cr/9z1r3EtXAuuTn
F9FJ3NDWDbscsGhLYRfCssUQTtt0BKXM13bTkmEaTQivaN98D09NkTz/4K79XxZNoNTSc4qoXrGi
Mxfi0pek538QOIF2qGCvlUUnbubOcw18iuXZABSASIdkHEBBvuPtCttpN/f9wA2xJuasZgJYbYHB
wVKeSuJiLM970/tU8jZRznzqo4Rki4xFa5kJJ55zQ8/HhXr9/CcfOFRIJS0tun5s6zbEwRRoBHV7
YmQldTfd2gO1LLUZnZe+eB5C3+xPtDTMQlqEXdD4tkTH2s8+vxZQhPWO829oWTkC52hzcIz7v37N
s3XX1/g/7rgm3SzyjAcNPRZEsNFp7ubB1Buy3A2stSv57OQJmmh/PvGQfDVeZF/vnAO3AU6ljXvB
Og9R+pQNl1YB+RoH/4OlyjUmfuNK3itnF7ANTRXZoiB2zpac9a9/PUn4QoSfRsftbQXJBLmr6mhM
W06HMf0HjG5KwIGwHoSgxQijFEKNCB6OcBC0GovjeatD+IGvpzpDZYV4sYeA0RY3mn9xYfqbYabc
C2E7qhuiim5qwpYyxolnCH3utP3TzuWFN5tuURLUeZeQsMWszOxBxK6o+Lxyefm4/TDaaLRY36rG
bcW+c+MJj2jOt7C/jfeQwFz5hIvaJtRsyhroLAKqG4Br1RsHjdlb1M35wVdw6Qm2m41d5wkaG70P
5n4pEFpPk4TwvdYA80Gb5cGJxEgM2qfFDsbkSgxHFTS4GA36MDtN38gcb5lFWlIf+n45FQq+/tQN
ZJuJJASvhhCwI6zPn0kxOu8vaPhMyyY7/FwIZvAV0KLN1pyXoNCVVTvOcbDx8cFm3+DG2ok61x2M
PjofrqlCPPJbOBKyfehGfsk9uYdD/gWqKvs/qum7K5Ne/0/JjMJuRrZUSWbkVdEoDEqZmRkgG4M7
N9NJLp8cFypVNd9ahYJG01ZI1P+Y++1K+XKAXmRamPcwaJXFvZs93PkJGTge7Vb/EJM5QXw8mQEe
ovEXRqgjE97eQhrIonXGDtMmu2h9kbRWY2m3tuRcOI8rycmLIro/a4ubhfa4YgUOvDG1lJRoK6it
Tcs5qJyoPPeY0lAGx320DWzmCBH2rj/wIF8vXOv3BWgdWtWsHjre+WJrkZI2OVYs2RmCIjyTlaFo
m71q8P+SxBQHhxwyx/Vd7yO05/WDFvSj21qyJXEEmQV9k4W9mBDiDpZpSbxp9kluNnz2pVS1AwLN
/J+Pbtx5XzgBKf6vYuBblFMS1FKn/zOimUBvu8tXq0P5U9gaPuyXo532IT80Ui+ue4OPayWyIAIk
gy9QD5+Sgso0fiFGcjydLwdRvYM71W3PVcyPBMqJJFjOnSNUkVXWaw+RljZkSQjzG2feRK4Kn2ne
z2a0rPgs1LnnHzn5baPdpGS/EqEfEKeiOIh6yxCUusT3gTOB8eXuvu45GF3hJ3mazhF2hDHLwZtE
A/LQpa5/i0xMZCgWEgCEjwiM0oxjZ3xUE1oExZczYhnikyPXBdiZaw0yaMhLSvtjGMNSIBLvI1ht
W5a1MHaZSKYjfcYaugHOWUuWuYjroHTCIERSkOJvNN8h2wZNLCkM47g1k3I2etjNwkvFp2TH8Bn6
HSw+ThtoE4IctCeEE6ZDymHw2FrnvkJtZKFvo2t29b+g7pgwpxK095I2pj5RIFagRfqFPcKu2uuL
SOUmxI2uAETY5tSY6Y9bo5vTGBJ9vxRA5OVSPbe5+X8FvONC9kGmoedNRYuKq7xYcacDRXyCqFMw
lTiJo+9331zCjgdAqJZ9Miv555R7qNingwU7H3GYj5uqyHK9ygH1BG483FC2lSFkuRxCBNXhqAlb
cjM+OIGBLeIE1P2BQ4aVSsv9vx2hF5dIO5wz+yR5GScOlDAG8Gt4htlKNzT+IJQqXMu9Xp6i477E
X9meJOyUjFJvF7zsc+Wl1lt3sXt9c6BSlsBSGXVQZbmlLlXRo9kaENzk2hCymefmo9THvqCyQOIb
tpHYDVs6mVvl+RWqlScp7KYZtTAwEE2LrbSUEgUm58NRH3S/3Eu7BhvsvKLioz4JLed1GNg2t3mP
7wNfCSMKMEuaMq4bcaNLKRz8dpvMddN/dB7IVTOwZspu50el2mHChD/6JlVUPC5Tv4DXefnEKxjO
yLQS61q1HYbnrEwm2anMKK0BQoQWK1DOTsBMVx8ygj9WYFpi4SMEHXfkXGwp/ltMBWDP79jkDR0P
xb6eFHJD1y9a57764NA+6jGmQ4QaVizdCFA3pjaCHGVMqpaPhC68XHmmr1CuBwNIXF83jWcrc22X
zcA7CaavJGS4Srk+3d/1dls+Lp9ZthGOn03eTFErxC+cdCz7h/Efz+9GdtNqHVBZyFFMFy5OuWXl
9tR3GVfZeEwHCfJP4DKreEfR18f+mo7MK5I8lk2rs4LXOtsYhWiBoVgfqPtQwr8339xEEBMy9gNH
irkxhSMu77yr1y4oC9UHdjABTf5soBJaVxF1dzee9gtuIs3yifhMXqvP4U7hkGBi1IGScO1MIwIk
FavDnfUbs5OAdc7oF/jtQHafiTfTurOiGg2A0cVUmOm1nTYkFrS3L52q8MpZOB/6/4o97cHHUY1m
Qsdxi6FrYX1AXQSaJOw4PqR+g0vgLKx8L0WUE/2up1WAFHoLv1AyqmOXRCWxupLN28BOu7DwHaDj
+QWIvgctkgR8G/cqKPIO+W6vJBIClr/Naaex9Cwkm0Hf4ZIy3tXYPcX+vG/GBrl0LW/KjMmQH6Rz
jkh8uF4/k949kkwTg82jHbcV9stJVM8/sUoY+sBFxJKK78o7BlOUFDvsyELdHDqSo4fnrYpwjBal
RevTzavzk48WmW4VIDaLO5W91dbqzgVlTenKwNv4mEGdvIxXxryo/wV5z7FfSeIy0YYhaGIjxT06
jq7+zIYqld4r6kBsK53QXvbnSI+19j/9Gli3LhNclFTmYfF8GVs15v8ymAU6fLiu5KQuXl63vJuT
j+4tF332odLDfp/WFVBnPCA0KDa5mHGFMjBCmbnHWOlVKNjDYuWOeZjQk77VpIrc+RkGuPfv5WBY
co3Wzf0fuChdQCAy3S4FcZklQ1n3v/M5/LAXlMqLL6QfXm51H9RwhBQbDJEklCswIJWTV3SfazEk
CeOhF/6pT0nnsYsuodbGV7zywQcsy8gK5m2MiJhGP4+oBOGjMqDJFRKVs1fPq7sUAxGCqONsdxTL
BICpPXTisjHIdKfbcIq0i9mM/0cBN4kcuyDKEH5Ha0Nlq9nWLwS6dWVYSk4OFqDgy5QJvPCeh0MP
l28Irv+hH9A1CqtcTba+Ooz7YVmLjxCbhCiVQN0PBG8OSdvD2QXCcISoxIuPPOqQCh3BFyV6ZQdw
V5STx5/RV6rbAfY+TnvRL2ixiUqCfod+sxHJMaGkF063v5tD+ujjkeoCrbVBBRPHqXi3d9gVGvn+
+RZD3PSZu6r4Mhf59BvtIa9HJCnXAuo1x2k1j7biYc5I3b1JDRKlpWO6pw7U60LRNIe5XwEHJ7Xa
nkcfuQgBsa755FuhTPWQHpHkyuvchcg8ayrdmm/cR4k73TLg92SbcQFt0XsvLEoKtklbIgNLX4rF
Fg31zkusY9+3OiAukKRa6puIdwlOOsMuND+p93fFVc+AjvqZDy3ws8uXQb1pt4m+WkgWBfNup8ak
6spw3tuOLlxsJunn1o+tqwwO9EJ6auNJXh2iXshkM4CpIvFJkmJs1Wgf7ykyCYWNyP0TvXepnHaj
R+BTlirZHzcxFBrJuIG7uJOgV5bczjuF26tfgOdai1zhaN+dQwC4M2BzChU6Nh5nlbvGxovvX4wP
4sVSHD/t7a2XADr1XH0TflLmd9Bv08+YF6aQ7CP2Wz++z9M8/35RDlDPd9JzKbAMu4v1pmAJyGgp
G3G8pdBTjErr+uKtuJzPtA+I5toRXN3YyZTSUwuDBmuyCatCqqabf36F+HOSVBV1mHoYNGgeyTaz
DfwGtacAh55XBrvQAnwBMVd2dNVNaephvaN+pSvWpjdxSUTMvsIVFSNuNmVYlSTqwopdNtSkFyUG
GOYEzOrZM1DQt90jaVJ/awAylB0XCcKYSlCFLLqZAAr4Bf6h1qm8Nvh4xp88bg2+dtR3NrV+qhIW
copisG3EcOyP5zfAJgdA8GJvuVuw2e9g3nwrcgNPHmHsLoL/c9WBY2Q1s32hQVZDK6r6St+xcjyW
YEgUeZIKwSN3bXqdALQdEfKybq85HFCHD3indWe43Pcn9uD/kLaRi+13fkaCvCI5y2nfLF2x64dc
pRSD0yjsSeJVrqw6d+LqgcaHiV5bxLnryWaqLNAAnC7/JzG3vMKn2dRTzq8H4l92taEbKhsHIpW5
ywM5SpqXvhUeL1Hmq3yu1MYe5JQGHl56+A+PORpiVtm4X7C8wQwoPwysgkcCo6bFFR7WvSNk8cGk
T9KTcrXyLxHd131JXzeWXaH0zgCWgkCLqDwjiBcnJlhoa5/H8gwa5ohkSAC3cbisF4Ba11XVLpzb
8ZOVw6fADKyaB6lIOcsW86I2FNn57ufBS8QtZgUQ+G3B8+p8/VmK/h0YjFaciwVxm8zVW3vM04Ez
mctNwhPrPDHc+a5eppDWg4h68HAk1XXcHJ+RbITeUzcVtieZhuPRZX5WuIcwo+7YkW+KrIKf/kkO
5S8UPL5n56Ue9d2uF8EYM+RDzJhmlu3aDhPzLPvBefUqg53aTCpypZ+TGReWuq8LrId6KcRAIDbw
yCw+4kQ+fkiKwUnLP9vPtND4eM+2zcgldFkDehOD5cvQppTqA0yYFXhaq2TAnZNo0R4JIbX3v3WS
TghjJWwnPApTk9c+fls3J02b5Icm5SiBMjKHw65kq4MZyG80KECPGgCnDKYNv8YYPUtUQfJxDpB+
5dkZTd1xSnd9Wz/SflueSh6xpMV6gEPTwVOHxDsFKXIKgXzj7ANZYa5rkNNO3XfOW7eDTM6awXL+
UoZkvt4/dJavG5tN0umNnDlJrsX1a0iZENyi7HO/6mmK3vmQ3977U/kUYUiA77Qk6HuYVkQ62VPt
9qYZtrYeEBmjYKbp+StvZ327s1PG87Fwjq8N0iBxX8fDZC5l9cSd35oC39NDInI7+MWnv3FXR8e+
r28X7dZQg0FNZQvG9yombY98orXmRw8ccUA4DnFZoInbaw8+FmQnKJ+qegflYH08hKmrxa6Z5rd8
nMe8ztoQ3LF/IW5v9suLGkPGTYJ6Q+g5MgGkY8C0DAhWd+GVSRTs/QsXclYTZut4x2cbQ8bL1CVf
gBssVnPM4weJp2wi0owKe3z3y0JHgOjjMZAHWhSaquTAenh/FnCdwpBKH7AwZU2siQgFcZIlRBJG
3jG/PNgys6wtFs0YKQV3rJRbal35RtF27fmTzQ3fJHzuL0FhTZsfmFzIm+ZXRcq/PevkfdoYjN9k
63+tVVye9S2nnlQVktHCWv6aPpvDA3iqzCiDWV/ncZfzh02sRyYOvqLc/yGSKa1iCGU+S1RayhUV
kBgRoU3sgcFaN8PcLfmsBe0xgnmblb4EzhIv48x7INLGkIJ0XdablPZe5oBd0v5crpUzP3t8rGgC
InLKdcqnM0soWcIKltk+kBLRF4YsYublPj3sYvNPvW9gp8xIsL4Gfp/kRrtsEhT7jUUBi+/pfJHu
Kcxs8ZQYPFB1ycAj9O54ngiWEwXNlfV39QzN3V+hHtKVSllyweg0guANA7G/Uoxt3EmWS8nLGJgM
JF538X5/Xlc5u9TJJBx882fTwfB026vxKKgpEoVBZa9/z9iwVTnBHstq+B5l8P3XjHBYVzqxtJt0
r8WQS8BcoxQOVvmwUn+PeiYx5czoq/sGZGYGyHpgvpRdc0zQSb84wkPKVgRXrrap/MO2VNs3sxCo
nF2jvv7/9RYbT6YeCAdFSB9OWMywhY6JwyQkY7ww1K+Azg/OepyPromddVBT9bQGw/R20pHTSlar
/V1xx+MeyVMbp+XbsNcqxd81KWVYyQFAwVnA1Wzzu0a7horJCkqzEdPNapf+hMxqcWPNbj+DNZlI
xsaFh6168gjwBL9IErgZtzIHPIkrN2Zp+LuRgWYRJmsSPbwBfrCr0wk/Nu91++rqm/TuyJA8E3IL
QgQ0Lp/e4zih3VCraF6NmgPTZOZaGS+cpBAyUTDxMCy0QSrcI0bnVtjFFCM4YOpXRhoMW+ZypSsm
ajE5QJ7fCgTWFSipgTzUt7inm7Bxv60wwdnT4IrjFUoGAeb6QhG/v+ES2f9BHkAjwr/I1ybK2hZK
MyATRt38RxcRRwn1GXAwlxxLOFBE2LiK1p9pKPPBtAsjhPaw060optoJGmPszAOJM429k2kj/Iko
PGdRdEYA8iYSADOvwuLkpiwhSIBykOCjbb9S+qOa3h7ljSlsDI0ZD95gRjhutoOk32aQ55iSZbJK
nj7S/5WB5n5Xl/BSLVAXcrxPKFDzGgAZLs2s2uofTv2gb4OhzmFuTKZyVmPsiBt9jT94BZKpig+h
gav/lPsmSUXOLAdlUjl38VcIEmnfnYOas4P9HfMtdEElQlEU0+OfdSeJT/OvDVTl0mHk1bYYjd3+
rqtLBlwwtv+vF1ukZK6tjZY/mUM4kXk3roO7tvo6AA79glv+RpoM05eFJsucv/spsXzQcYGNkoTI
hywhmIKJhzeEEVcqSTtHuGMtGgLhmgVo2ZHVHxC865KHk6z5HKPDN2FUK/9SdHorhF2Xi88XLvcU
u9VrzPOxAdCUTfieKYGJVmXCBrmPws8McxfIQQwBqAN+NS0SVaVbrlCbhX9tdwTtyRuK8yd7kyLL
zkiPPoeQrNDOH9ZN60JjDN9/QuShaMq7G9nSfJjkIYm8ANcc+dupzvTyCp0rQxKMtSPrphGzAgDh
ShWeau6gEFWyi0WAuWlFJul1ShGGav9mTwZJrDX+dSdJ4n1Y15GCq/FLWkwIQRAy4WtLlW1ym3x/
1PdOrDpzaNMmPqLltHT/QVR3OgCrZkk6DpxPgMk6IipgbFSRCCRTWrqeFUWz2fBOsCIN35pARDVl
8p45fUyhq3MPv01TxKDVpbtN70C8llLkRsAaDpU8gFhbbvI4Kpa2Glhc0nIjGzGP4M6iHaNZ9L7z
2hTt1INlS/XScuhI6c57HkHfovR+k45G6zudxrZ1YpAoqp3fX+ee8643UT1a9gsvgYT66qiIPtnu
cGK7tHNOG8sskjY4XGotPx0Yy0722H2KZOXscSacrukQdXxpy/GASrC9fFSpbRqqrmMzN9Co5UX+
U80bud3RXV+dbZ0oEvGytgJlHhcQq6hlW3HPGA+0d6yBiRbOKQmL9DwW1sXvSpohXXQ2mun9Rx9H
gzPqsHEaoyf8+yw7oImkikvUYO1Nw5oE5IU1ueqr0mI516QkMXuKenN499qyLouoMkJxqyi+aZxQ
FT+tI5xHpNGpZXqQd7GySpeUrolFYsnlq2VBcyxY+2nj0OhQPC0wH16zxAfcKx6DDf7Sc0DWS5EY
huvCNQIsMGZMgSy0Ra8x3yqhXFcyRglel9IEcXcnC2cCW/QDZ1SlSi17fxhcCbfAcuMtffrpjjr1
P6pH4WdnGymma1zkILfIEhyNe6BhdVz9X962nad5Vhu2vI0426/ePsR9/NuxEhn9LUrqQerDCJkf
lByP70+2As0mxZ6XwE1cypaUzcY4NxRC9decMWVuthZsqAaSJTXhEw2eBZZ0MMA+BSXK7G7hi8ik
VEMN8YtTW1C4tyBPUfLGxGgY6mW8lZm3602a/bAWsJIYQJCiIk0rTULX+hMWmzS0D+ymB/jsvOct
iLUeDG+/gjat7xjZuHYl6SAokh1Sw5yKyrqqYQWdLSW9gXSJZMhD5M1LcIyKAErYbi8qM0F95WX7
8UWih3JgCuDJl6o0JjQzCAecQNKQ95JeXTsDzbQLUXiAxw1P0971DiyQxCsDdpvvvx8/80lz633p
q7zb8XRr+KCA3D5XOsCpknvUDfeGih1vJnpb69J7e8eI6SBw/UmEo64/lZhYJDcib3VGdJGHM0oM
ryf0eBq10HLnzlMT6wDbAtg7z8CpwFylbwMLDV5kMWtr8eZeOHFMWYFaAOm1GT0twiDE8XXLWbYL
cs0JFKpyF2u86bnY72mGII8z2e5r0quGo6bWZCAasHiuvsjtP89hq0l7rmSk7RqlebX/kOHYrL8Z
SH/qLfZIPaX+efLuoz22o5MUjGD90j7trgxo82wUfcX6YM2BCsiYZHnohWokoY/zbe4uOY+XexAp
djtxJ4+7g8Rh/chshhfgpGqktwXcPm7/bdObpPHOI64eknRwYaonyrz3Z4z+5goN7qyH37YBJOhw
WzjAIm+bRz/SrrWB4A/eCg/FIEDDi9m0HQY+G79jGXAqYGxwgIYXI+htjXid8Cm4LPzrjpRSwoyj
E6Y0cf0ep+KR45gOr5XVE35ShC8qeigX570OQYJiFSEf+Ey48e4xSkFyl0QKlGzqXr2CYNazcjQY
dws4ZC/E9zPLd7Qa8Il6i/GaW4hjFuKxZ5tpq84rej+5or3mRZ1856b/sPmxOYxy2RLDNz/6m+8H
/tfhLxsnsNvLZVF7PTqJN5OV8AaavZr+xFvW2zG3M7vX8UCEcNaMv2jIv3X8JT2EYdGBpdobBLRL
9hKdEI+5xtumuHEs+7vSGd3/5NohSEMmJ7Sa2c5jiLW604mJxZjXE5le8wP3nyPEZdx14xyTFirM
lXHuaaRIaaMorcXi4pC+pKvpicxJRQGoShInifU9A9268wGWGMDNRPGjunnYUe35E9WWSxeHL1K4
VL+N0+8UXob73DkA4Ymm+G5EVsxrmbJyKu23gOkKEQ8eNX+E29mZvE+NCg6UdnrqVqEAJk8F5z0B
kgWfRhkhEyLKMcc/YsALF0ldEfAnOEkXvyEIEHhSrjF+Gs+69aZRphaQIQYRM5CkdQFjtm5rtdKG
rxaOgarbbv0/Dk08A+KG9M/WKEsgYak1gHlQmTuy8+tSKMK/3UW44APpUq6hj1GC5YejBitK2ast
poFNkUSYaJIpH905bwAC8DVWdO9P3t3N8GTjFNyEJn7t+zuwDUXo/mG9OT70Fduteg5RaHv9vfs/
UbHnQenM+nrVn+eLkekB1c71OR/JhN8y616wkNXrpySccGvHO0C4ttnn8AxrcdVxXf8YXt6dwguR
YLbVuZx1Y6hHdoqFTLbXQMNNxo5vm5gkKbyQI7gArELFLEPJhSNycf+DetkwXBfVOYor1w8tUBAC
DhEWfDxeSAdrHMm1YDoCPkqjcBvyDLROEu6SpBeQ1YDJqXq98jFnYmN+3EOp1mQ0J3nDO5i87bTZ
RTvnZFrFdzWslgzHAsB/+wrDzFiB2eXQd7vBowYhkhJ7eEFpfrKrwMq2hOYuSzR7hgd0Gu/B+Kzn
yrHnKlsRML11H/tqfPNd7WYz27LX1IuuMtaDaaQ9g3isfPcZx3RCr3RIwqq0s4LdfdjqGFQticv7
qLo41YrGnOmfVpr09GFKZdGAvgdhfGA1x68uOMsEOujBJgiLHtXEnY1LLG7ivcLoj8ue6ZueHzkz
zccJpD89CHlAkwNP5g32urLYl7YdOxFRi4Fbzz586jF8nFw5xJ13OFJE4hjddZ+rovvlHHoo5NKm
7llbXItADjtFulaV5xX8TWmNTRxZHagbOM2fG+go7rVxgGgW9YJAWuH/ixzI1VLl0FZBHE3LaApK
0mTsGaB8FfYGUBzCoqdaDmi/COdU2iuVK5d/XXY3bTx5iR/fw9KcIzL+UnZr/77RDSXhKpUh/OsY
ni6eWW7YM8M+lIXGiAN+ge5S1RTO728H3nYkZ9lGY4Kf2vMEV71e5InXZl8puqxQyHtXkFSxEVi3
HPqQEM3vkeEBtNPwA7MaAJvg+KkESffRGBNv+OzHEQxNFe7mbQWh7uSNhQ17nZKiWdjQNli2572n
PHm5JVE2qQ1nuwp3K7HWARuVq/VZG6wo0s4vVYSnWSnodUhCiK037GmSI4D43L/hU+s9vW5EybjN
GW4JShBOOeDouLkJNA9IbrjyJVm/YBq2Dv0NpuCYNsYimnNcHVUqCIyt98HhaDWrjAKyfMte7kRN
f9Xwr46c7zzmtv4qGq/RDbcVmqCTBtHhGDFH6JZWj3fuQqiSxQLNeWT2J06oXjUjBLWikBtECpYs
4oIhtvsKRDcALvfZ6OT6iE3cUGZTPVsN2MaLF1yLVpkyavPPsWfDI1lWwyjJLUnnDH+BIaYur00v
k5E0UphX18niLQpC3r3I3wMsJMiX2FsCKzz1nO2rizveJBxy3KkYjldrdTscrJrr87z8Aix+BAc2
8l4VOvKQHEwFDDbe+zol+dxTREC1MIgeCVnPcWedGITom5fi5HOvMB8j1ioLnHrZCTq793wsIltC
rkRdpRcQLFmeavJvs86+1Mzb6upVWKAUU2ZxHzLU7LdWor8lockJ6vFoCml+5r5Zvjzhn6S7dXW2
RdXdhP8NF+myvm/cZ5YiIqVVj2Xt4h6XfYi9RWHTfSb8dgHAESuiD2AKNVVTfpID0FpmIex2UzWj
gIMairPaSJXWZjINvsHMXXfKGCCQEyRt9vOchoy4r5tMQzfzlSjsbW2u9uLXD+8+kAzsPGoCIvJB
0Bn2PIaMb/lY1ypQDrDDcwL0MwAeZUHBHss5z/GsT2WXkbow+jloYUWdKRWSTvusP/ZjtEQoAuki
VDIlRG1fWElc/cTo26MgpeejacQ5f1xKlF8fdxKLID/5z5yQBrL7Oh/pnGjDkNZ0ux4aTeZ3lPZs
x/twkaMu63oq4eXXbVwlapiYRifPohIDpZBwV4VswUm4wlBKriEMGZrepQiivSE3TMGbyXn0YXy4
cj0yDjwTCSP/HhiX5MN6YI3pz7n22YIc6/h4l7g/+vqVkAT7EtDacH3O9qqLA4LZHJT9HoXhdsDo
aC04So0QK3QKM8b/EOeXgFNAWaCbtFzLWfBl8/1x0yJvdnOIYRRTPKJXB4V3xers/BrlRBqQUR3h
FxowdKXmYyJ6Ts42sXe/x93Vrkwi9ZtySqHlDe/PlNi4mkKPnmcD/kfRk3ARM9ka5YUXwAVkU0QF
sxvi/6yhHHhl2ERnkTA8HWBApM7CFiLnYwpca4cr0kVbTqlfVNOwQVQNvujSxLMiGRdR8mnsXVQk
mB7JKEnivpY28zatUcTbPRVzDLH6R080xpTKc0Qxz4PRBKqBg/D/WdeXtMKpevBs2a874fyoFinq
9qyTC3TdMn/jPev+Vzs+82L2A82By+m1w1VD2tos60qqixscDaCrL1/R81KQ/Tm7OWumao4a+lRs
3OGQ6EWrKg3XxOdSxAPWc/8ntZZoM+/P13NMWfUXUAjjjWYYdATXqU9SQ1z/uEku874b48bpGgpk
ke6USfrdH+6iNbhbTLL3fwgTbOsbsTf9GzfMxmUSMX8ERz3jJp/CLo1LGCg1jG26alEWQH/MZ7aq
Z+wOhBX+VsCMR2VnuhG4ro54lQ0A/0Ro4lg+mDctqnFDfjy6SqNSABLQRaFq1YI34aBoU478IVP7
Rxke/wYxQCM6GnYE2DMiuPro3wX7GzV0K0wSvvIUbPYMgaI8aIFYgVWQN8bx55AOp5EsThnWNcXW
UAMeF2O9EfiBicvNnhvmoj3dKLrjTr8B9347v0/EEpp+EgWPaqbMtTpxXEm8gMU/KG9sK8PxbiRa
BNDvODpJbgD5wZJBymonm1774Zcj9oMnnVxjKCb9ZqGN4E4HCjBJRmPskNVerVLXnxT5AjT4b7PP
EUAYmcoM3KeFlfQXwI9Urvt7ffg2hewWGTLaFe8nw/GNj/kMKnXy6EZL8BG6K747SH5i1HXaegEG
tFglU6uu31Stq7cDAz2V6SrycbosTU4lMWl2ymPb9NeCpNTqbshkjF7eMkJPjQr3i79Siceob/nU
O5lYNw4X/zW56QVnuhGGu0Mt4jaGsib4EfEwGb36dChxCDpQNBcjF46sgSyFTMK5F1ABgZzcr0bo
H/Ekv3Nx9mzQLMkfh7QZ85AMcJmn0kF7/uSMgeLAbylFEyymtwau2MFNeqVgosvk1/tdcxwaVPxI
knw7cHKQHdAHrYydaDus9aZLZYVBUXeZ+MHzlmgb9sLeqiVEkl8oSkS5IYy5Vhl7I1o7jwzb6h+E
g4Sx/2jqeYoISnz2B1m812Q5AtBWK82+8V/PT+4RduFEmwcBvWWWq4FrQ4mi2uWmWM8pbxZC2Mps
dJQ2pByTfY2EeY4rxD7uN5Y9pQFjY5BVepuuWaS4H6Jazl+URLeYF1eYy7KiHnUvZikFDb4MoSJy
DRlI5job4anjXdNFkI6KSrPLGuE7XziUKELPKmshfBPLTSbR02az9goscKIRL9FXarnjwKuJUbgH
pA/G3ksH+n+HZfeZ83cVUt7uTb//AHSzefF9EsCxJAp7D8O8NSImLOb8k5VYap8dSSRB3l3f56T9
pXGWEmMxsFYJYvx8f92l0mW3Co/hnnPJS9Drmel31/SJ9m6CUTbw1ft7zzK/FOnvFwVWPWUZp6q4
tHNad9v1t/yTvgYBw3IVQm4tIP04Zp3578RK8axg5PCax2lnudaWnZfocy0EWUOPWGi0P/AlwrRN
haHjOknA8dBPPH1nWhWTNUuJb6NjDodNq9qbF/7xaBoBhV3FitauXuTb6PJY/M+knkRrPHQYNm6y
xGGfm9iMnHg1r9MN/Dqbrt+t+gpPFHW7kuqqSnGv2x1OUHOkZgxdp7EsR9dVBfdDC/v5t54Eq9af
9h2senpot4nv/CxFU2+2VV4ffn5i/f8Cy14dOCa+GeWX1irUwF08cMVaj6dSVDDrXK3sGuf3ALmd
ipx+wASws5uk9pLQN5+0l9oVDjBA6RJh4HzBqY/WXdOdZWwERlK3UkaKChONArjSbx8veMQaTw+0
+dbo+GkXC4Uvy5vERcHfVhe9FawnizMN/7X8ZLvlzt7e44QafhnlKp4IjD052i1iKt8yXoY07ls/
Xvb11q2hFTA4oYmZ6k+JiAIoZRtX4V1z0eVxMKCU4GYyvOjSMNENxHd1o3VLSH0cmpJGLLukXy1K
QFnjMDu/XLCrDB2M+xX6+087MLoKY4FK7vJm7z3h4EhjsBNyBrlbk62tFRBYl91abaZLVasvfUtF
uB1u0YZ0MiBzKF9XC36G+udk1ALHhL1Bs68gu0YzZGaSrxWZD8+nUgaWE+TRiTE7o0kDIK4jMxC4
XIdRc3NVH1atbI5wB6kGfOgDuFJwGg2vjbz0wqasBPv5Fabsku9LFZ6YcP29zBgL0DyjU2EdFP4f
GvEY/3LzftCYpXX7Nei6eUzHtpb/JrCxDtBfhDopQ3fKWp6JkGXLtS9t5bblDKiE90FSj1+3XQop
xoOCLkC+ax5bl+fyOm3jYQY7C8hiEzL2eOCF7dCCgGnvYwqcCCVCD2SnJuHhHold4RHAlDLXQqdb
aRXiDy+dDTpPTjzbnZ2OmAktWGY/dyA6Lh93w1bg3iwhXRy8ti9XJZIM17Ry16m65GyhEtxcUi1G
gmjwGTkybHxOEvdWBzcn/iULlMxhI+BHqnL2pC/OWRsqHNITH3sjITOruyjctIU8ohvRwAATITJQ
/ivPY543sSvtkVRqiw3aIbo++dCdBCRETSwCXAzkxIk+0wCQOC0OeOjHn9JutnRTDXR4rG/G43yu
z3QutP+n2oJ4uwXOviHntaSfK+vD036U0nWVMFXPuZ3vGwof+E0Ih9pMgAIHfKBJ4TJBfA1/F0ak
Y/Bc/BEzB2ck/GBPaXnWAGtbHZce0MNjdUHnLRz/5MJBotHommnEQDcYM5AfM52oI/u32uJ2D5Y1
G/aLO83iWi5Hh695kKZpHLRWDGpYUh2Vb8E/U7IjnJRNWqNM1GTN8U47DmyCy76kWtqqnra7RlcA
9dm5zSRRD6Gv2cYM2JUYOSfCXssdW//cW9k/rO1mbYjnbt+WUk87c9obbXt7IWxB+D50wzohhQ3S
pPy4B3eDK+pHa7cNz2Xdtk8UQXOLujX6VjcBf94dYrEBaJNmQwL6Y3v+F+JY/2g7VsagXLSxTtKY
lNKiCuPYECOP/0DWyNG9r8Nf3cqRZl/M4EgoOIq3GITKW4Lms3FbcZf67ORk6xbpm8PcS+j9tgG+
u1gcHHDWfVxGz3r13WEiNXcwgORfyL7gHZTB6B/Ww4AqUW4Kh5iGcrm5dfm8tmmy1qJWD28V9wSA
1hOFK4qR+lnxe9Tg6Q7XM/3w8sKen3pU7WbsiKIHvtgVslZv65JTtGzRGdZ+kPQdr8MqwF/KQbC5
W4pqB6r/PnTxtnTgkAlLG3HRlaq/uwS5O39YgkWofrrk9JNcvctqpWu+3VkgZ590TcqLSWE43GAO
vjQBJnawQI7L1Hf/CvXtsz4oD6pEe7CpK7TqxLSyR1r8oFTyWbgsh+jHyeIHPOhhw2U47WEQ9Xts
xukja3idkBGtLFJ3vn8U2lkbOu398FJMcix/5Ec8QiOtXmW454pZsSZvBc0noM2dGPT4HxTyrr2T
6FOZRWadHpJgMrgFN+YbOgo1ZnUwbF+ykwPSu+Na5Z9SeAX/39p9/rXmUiQ3bN2n9QVQlSee59DP
Zj0yavIcJs7eRHC9HH/kN4I54MHZZb19Vmge9uDethvEhilTKiYmON36zhYJjd4c9y8mtJcRgqwu
G2cOJkVHuqlo4Ezvx9MdDZra2YhF7u5AIfhlnuWTV16Lb8xBtZw0l70m86DYmxIRQ/e5qi7a9qVL
qpepkI+d94xYyCfZflpF8Iia96dhM88lZycpdXJ+iApAF/d7Ky6AOuFZZWSXc5VowiilN85Ank0W
CXlHttlv7+H1XgYJyO99mco99UID3t1tNy+5q8CHfTBVXBTA1Oud7V3+AYYXAb0Or2F4EM9N4uNq
1OUf5HgsP1L5U1v6nABY2OY4mXYaYI5lVZsbhh85DkWIcR3A+1XPw1GiNeE3F4CbDvgxmiyTdCgg
VV50AHOegRYI7cqZ9UWtIjdZfiPUq2rRERyHRo/iQ3iPT3ixlGdrABXKnq/dt3duqongimGssi7D
bsuJWmvcN4iXC5xKewG3yS0IHkBjbVePjo2oE+UvXWR4J/+/kmeTdkysJ0zSM8u9xM0+fA/3Y7uN
sqfVFmYJlZEp9PESp3cpp1f6Mm3P0WHmeScNUFLblupOTCy37Ax20zp10N6i3R9WUaWZhSHvn3mJ
iD1G03uhdqNTpAHs8c02nb83ubyAJkDTviJahHx9MdV1BtD+SJh+O2rsN+w6fLX+9GGOuOzuhid2
YYnoceDWC2ekRfgeTEZXTBUnNUIGxuZszr4QKqm8qRB8vkUvmKFxAFAHr6xe11/WvZdQGwxokmA9
5l81xUBGzyEdpf0vc3aOGCw5EY//3Bmx0BXDf+3ouCqin9LFZO9UwljoKYjgSAL2e5Rx7JMngF7F
NpnyYab6zKlBzEgMVjTb5o8bnXf3/pSo71NYMLfFzw1hy2J1ktBWwltNvbBh5UgXeexDV5060lVR
45GfA1x31w25XMvGaIffw7kOqXlzLB7VHMPF/pCu3f9Eaydj4w4PqEeBa7bCcBP/YCObiYWMKss9
74QGQVfDHsw+571MPGQP2LhiwzTplfmgrX/oK0pwcOStP/Qkffpx/yhhLnxfcpLv076jGeGLAy2G
E+xw2BS9Y23dwgGyMTNuWd3rY5yvlj+fpA3g4vq3VBWDt2oc9sItMgAU1YcA3/QIG/FehyN5SWt1
q4VP0AKRiMxrpKjrCMYT+1qernBA6U4eDbL/ErURKmmm8ag9AgiNhcwZKTQImedAwpcOiY0mIIeX
4EOwrd8CMnzMk4l1drp/CBelx6sZc04fqt/qaKMagl7P/Wpy5JzLOCCys6afwhxLmmAjCgN/B0xN
3am3ehxNn9jOm/tddPLliQt767v0qFF1yEzTi6F38/NLER5k0z7QbydYLxfHkUc9wFHx0utGg9rh
Fu1Tl0MxOgMs3rsD+kFtVqgndaOmmNje0AIEvLQ8SC0vKb22k6duRk0a2cIWuMFVNayDsg4pW6hY
/hyBJeH0FKYepC3BZAPsyb3zVNK7+5ryvO8TyG4mCZ+2g4dsgGjJ8ffrtqsNoIdpOUT030wXqHX+
A8GGbVD/nJhmJNmdi0gg30ym4rpBkmvk4kMUKtoEEOdBmED/cbEPPWnEauyHPlYZTIBbx5m4QQca
onHxZXxrQdYTxBwOdu4EvqIOgbRAl7oGMaZTYGKrHC4LWzkLfgGx+uO/EB1cnpn90CWcHIBySOF6
lqPF+WeZ/zjbd7b71ofU1W961mDbXmLm3tRJS/m47C5UWhnVoMKxggsnY2M+ETHdxA3xKUuLYgAS
h86r6cO7Sohpoqd6fR+SrMKGlU3TMKwBx01Kym4c7ZhpHvDItrtIA0yvctZ+0l/wC+HHLmsvPnQR
ObS5FH6ecwCiMJvnEUirm168Vmim1vRXLp+0UOoZ8tETtG/9wSG4LOLWoCHPSml6eK7OgcMSMWYN
bRpgXOOMZMS0ayhkZ/wPo812HjL8Pd9TD0y3Iy8O/T206mbTFWCWQFEnmNj16JWn97L5BBMWBm73
0/V6/p18+aTjUs4KnI+QahvfQdcbzUAXE1fnJH+1feptWxUZO7TpEz7x4hCUWml9CK6Y3H6FGfYB
sORKpcvgC+2bEsfhlq29ShcMoT9g0pwkNRLQAPpgO8Baxn0jHyF7/BxBHOtcC0gNr/n1Xl6gSjys
AmogIH9jwKEoeR9AsYbFxDPpH5vmCDfAyQCqc+GAT+/DAGo2Yi9U4UJVT2lSMvE+APPJbo2auukF
HOt6TNOLCXY1bOJburKdSMWELJlklQTuP3O6yij6YPfjhJkN2hsLFQV7Ae3I64Ak5MtnDNr8IVni
GeyOGSQwf9tSK4p76ndkmaW4q9VFUi2GgGsGTQbx2HdYnveHGw3vTvBvPKDKmB9KjOBUxDuWMTRv
CPwB45D1zeG/weClLdmft5ZOUjXj1RBvwgkR/0LwIq8BUPe4RMb9DKdgeE7Fx0kQdLMawkJ+nmKk
Gucr2d7eZyK2rczhkCbUpC6kmYQygUtcdacfqZpzbE4KEpPHBbCoWw+Vixh/KITti3gCAFGFuigE
oQbwBNq8rePC2Ifzsm0c3znVXdIzCTywalUd3UT2kfXQr4tBGNolWsyk3kO1cRRA0xDjATnCPee8
J1Osmb+mpkfazIeaJzCWwSN+28vZ+vsXWObYA+D+1nWQpNP4ApUIJ2scMjjTuF00SI/PBY1nC7FA
TFhe+bptxfWknjUP/OFxeJPRndneiy+QJxHMJiG6uDvMGngjj8jK2i6b3mVV4GacuG4hNC74hrTz
hqxXYGgzspeGrHcqjHTSlkiAGSwazg1R+XP57U+aSOycx0mM6UThDQS7d8U17lHW4sNEvyAS1/Qo
CQ2n+qS1yT006uRXx9p9SAr3EJ1W8wp902DHzMBVOXYKCnJN75MSDp3cQzF9liwrtYmzJaH9x62z
c5hkdUu2QFrXrl2Dq+EZwVXpWuW1uRXTGjDb55M92M0pOs99tnoDkTf5u3riJQGSHFWtgAoPIQZe
R3O+PhiS+RxMJ+I5gCu3pS00STc4ljLMlZvNa4nOpIZN3Z+64iFS6kmLrh9n54jdJshgb56Yk45v
Z1hNJZ5it/kifJwKwWjgEFdBEBL46afSmyUyqOM53jhVKzrq11f8eZTcY8Fl63zbdOJnz5BvIMRP
1mJ6meeE0B2imfup1OH4/A1bRndPlbCoEgyWKAqOkifrnxg2vZJMz3neEhRjT3C3Nm9QgFLrtK/z
5sqyJEPnRO5n+ha65p4Nn5rjVfWs0NmhXHPjXzri6C5yIiGpHFNj0U1xD/c5whwLmQWkILiihOni
uBsp0TzFZmQ2eYbSmZhB40SWHFSTAepzaNmhxejlofPz0AMon101tSBg6NUCy5w+uToSzbsGZ04y
nbkCrZTe0XGYoQLOqcLFPK8zlDXUhtnb2H3+R6NDeMVBLqHKluV9YuLjDNITBIrO/thUCG19bvTm
Zmnf/+TX3SBkJQGiMInIZOZ6157SP0ec/NMO/TJzbwOwFBfyA6Fc04AF+fbNOfW+9qRn700bf+1G
XLBMYc/kX3EL4MaVT4GDoFrBMmil22IEvbLbGJN1Rwj9H3xhuE5V7vqKwPtU5zmLj2zr+5ah2D+2
u02j31mqskVr6YOnBF0tH4Mu0ECAlZaScpuXgt2Ye/7tZiq6pMmFYEEu2iqCp7/l4roAdbS0aD0V
tz/4Ih3T/Nrm47t6qMA8xmkxNeoVZY1zZfYNgXExIDTx8tviz4BFfhZpl2M/+yAK/7VNhfBMyNwU
/lBbG7CwLen9NAac+GMOPKDvfhxZGRBhzqgGGG7+fOMsgAluvklzPj0e6Rv8Xe/NdtFG9sE8tRu/
MZ9C8GZy5VEUelNPY2ady5oAs0NVzhxlbRklnLFrseRj0yQHxKc/q1c9BdeZ9kGkzmH4Hq2f6AMs
n0jaGs35Fv4nQC+LFaOIZuhmI8K4hImEd/kfFIurKHFbbw3ExkQbd1ASAfRYWQHvfIBe8OODs8B5
CzNkr5+Ca6WarwFHYBe9TkBG/kOYKeed7gFOZoeGtbjvA3miCascufQGtJiG6FdzjiaLjTxCnmpV
Gz+YF9HMUWHvAzmwvhezqiqpvZa1hM25aDsYYC3Ei2izrGneHXKQenf3/ja7oFouA9zW8xv0kRy5
jItOZKUpBIvVnHUIh6l6qNObr+KmaSJlsPiIOAFZBAkVOA4K0p6BxwNYjn/fJrdDPgln5od6Zgs4
NirZZB8R7oU6aHpDEtooSpTSS+IAuwiXbnABW0f4ro9KJqELuaX8x6H2TERpp2jZ9E5y+5ssnEkF
6XTqT2I+3AyHnak6ojGqWITLkwvPtQnYM60qBQ3iFMYk81uKZJmFarIe0ekA3CvEgRXTqJFX4PVB
MEz5nisUtWqonPTnRtLXbW4+j4knhwsrostUauLVYLmJBxPkBALlvCcxphbmbtA1KN4SqlsgYuVe
cIPixqPE0sH70v5hXnGRE72RecnO9wjkq76oVzrK1DG2HU1qeXGfMdgFaZYG94+YgMZNzfTpJz/Y
zAMEsbpsUkyrCxC/HGgR2pkFk+sUamuSjMcX4zO6XZIKhFZy1Q9EpUyHPhomGQ9ab0stVJzu0FUN
SjOtm3ajVDvik4rXDjrSxSRqUdNvY7EVJgkRcpNqxRgud+Bf9DIu1nFkbzHxiRVnlPJlR3ZNqeXQ
jS+QntSU0tx2wd0XHoWs+uuumKf97ig8T8T7GOOXGL5uQP+Ht2Mvkd4y+AgJMOfKOWLmGA6Ii6uT
LyKuXAshuKapOCOYYPqr6VgNiqp3P8LZvsythnynOiQNeFT76/TtaW1GEZnrzzb0yQn9sc39W1ZL
dzwCR9t1ksgkXxpEthgvBLZXX0JYLVd/zfa+Pv+uDKllVe4j5v41DTYReXTiIytzIUWC69O0i6z7
yLCHgU2GX2lE2NVo1d2Q9LuuTe4xqHIX2e8lwBd/6XwZs94vlUbLN4f4D5eMa0cZz2AQXrvNE64c
JivsuS802DEQwF3FCjORukGdNuvitTDOi2LKLs8Jy7lGtc8h5Fi3eDcb29o7t6HjjAEeRT2Lgzvu
MxAMHp+7rgMmgi4OsnnT8Jg66ElhNX40TJVcT7bmz4EWDra9uJZTGUb6uhk7dzn7jtNifsQU45ZT
hnujONwZv6lywiS2TIBndZK6dpzGB3TGEdwwVjehnvsnOPx0C0W4iXwzcWaTQnelg3M0ORxLENPi
iWbWsH97Xs1ANM0nhs0qVG6w76W5Sm5ReO2DpxREX47OncBnCu4Ml27epUmDzDbvfKXoVuOnxxDf
h/atlz6o6am6pqxZIcSUB8BDQiF94MmbOvgck393cxwfJsdHmuyBU9yK3hXC2LzSBTEPSQ0tNAya
9w9SKCScZUkiIJTtirrmDQ7f+xvDF8j+ko6OgMbL7wYJo9f1ZeQSMP4EJrOG1dF14Kt23OUJSyMu
dLfjEbpr2pJxILMCzIuX5B3/s4vcrScQHa1hKB8BUkD2PQqBW5Bsyb2VzQJxQ3tudK40fxste8Hs
2Sez534ONRtiGPKnB3rzkyFpw5ETGeDAk2YMd7neYkGN/VbjEBPfqRrrSQgUpu8v7jap1lwFiFse
/ZRhHd4q0DvOV5qVataVqI3YAKqvWKU/YmuYWxpSjoG+OCbOYCN03jvjtXngWwrExt5UlCAUBaVu
4EIrV3tgqH52ZDNEUpf/xZ/AFEz5gyUaRObexxRXONOrTmmrLIGYWVzZzEhyF9ZucwgQUSy0VKou
UtJ4Y1AYbcWcUrEoLV8GIRAzDPUKZ8/V6q+C1jL4GCudFM6Dv3sW4iwg/WyyFj02qUlseir5UsYF
rS7kK5dgcy9Pzbh63VjzZ6pKvP3q9Zlu1kIh+CPV5K3D8UrM8YHF9q4sip5mCm6JXtY1qVD6iZYE
TAweeVZ+T/+VhuWEf9cxa6SvOm1EPXHXplhEJjFqH4UlbUS8N4y+aFumZszl1WIKv5kXGW9L0Knj
YWJ2Bt52OmavsBCjKTEJGabIc7WgbAZPutK0Y42k75MA0ZAOT9Lipq8u7BIxRbnxdFRfyr/y4G2s
gDRiS99rflvDQOv4OD0SwIRDWtE0IOAfWtTyQ/XwSNEqkU70tyc9+fMBCwIjviGEouYOWUm6WlFB
8B2zDc9JhFIrB+b7PR2Adq85ICMGcOcys/KbhwnRWx2hyNNM6oyZTx9rX9XHTrZ8VfY1FyEoHlBL
gjifjdO9Zu+nN7nC4Nq0gXSF+l5tjGtooOHS9fpzhPzVTwulgHEjf1lixQz83Fg4F5T/UZ+gLBOJ
e25CyFl2Aqi/bzfyCiVs0iVWJWGI4dZk6bFB996yNn7XS9NYWOjWITneD0j1LbNb8BJrpUjR3pz6
5WqzIbrkNVRmhPZnqU1KtxdABAwTCzk1z1Fm0Wzes25LS/FGi+TgxTHQmvDe+I/ewwYM6IC6rceu
F25H8MJSjJYksPBQwPBcKC28Chapq2tAsmp+mYdZg8l2B2QE24o7u/ZyDI9qdUrZtOr7Z+DW34fE
ZzLDni5zCRjXcxfZsayZmQLhoqJU3bljxVRPS1tzFekzy2yBcL5NTUPegJbfhOkeqEt96BkvZZWv
+ugyi67vXwt+sTBd/XirL6WrvntA7kzFZuYXbmqeLTTGTgZkTpKVnzmXXdTJ5LcTeSb9nMuxssq2
QzD6MeQ5T3zvZkPjrmog45QRfbvtsrma46g9YuCQ0DigUjyyQvfWJNEbJweMIquTrQu7cLLPLR9H
px5cQO6kZwFiOXMKA0N1Df6yIJ/d73J8caGPtp7ukZN0qugnQQ1OkHxE9891I3jF9o4wJf6IAcRL
PdK/13/u9tNoqxITHgvU01cqR16Mf/8aD4PE2fhOZQAsAkhD1AUmRhfDeZqfqLxvpgQ+W/+BDZII
jE34CxWq7QpemJa6g9I9C5ZDuX32E4hoM10WKDcOxbbGdAmQHedJvjfrJdgNfZWivyT6yBv5UXNG
zHBKYtavLRigz04SiGJRhIx1OMytZ8g45Esgkly6rpbKZQjnzSaX4Ds5RA0uXfOHGaMgtzgGTz5m
coABij4fKSWtaJwRsDlLDYvamPIlOuGl4cpVfp3PPamNxKZij/FJGEeb4U1NrR22ovHoIbDScqUA
V3G4TfA+4GraYlEb+5zbwezyObLK/ePC+rrM5MKDFRNikAufhQOzEswH5LuK3Cgq7JZ4O7lzmv8E
pMWQSIcRHLqrcY0hE36C16uiR3XCH/c2KHpmz8lPren2dkdxe8tKJe9ao2GRGcPz0VZcsQQ7zMTS
hC0m8//WAMhpSSHMtoMIF57P4VRc97L707imwVryv9he/QUDwkm4CtnGK+T0IuQvQIVBkT9JA1h1
gySDrKcL9XiK47Rm5ST/+UQKtNQCpxcDB8S1vHh3ZKZq0v/JRIH1GeCCtoqqR1g+DbZLuWuv7VBH
EJKvUPaKvm7Xmebztihru24l4GaF+UpEaNC9YeE/0M4lLW+rRwH5DIKG8fUHsYmgyfrlZFSZE2s0
B4EiXk/alDnUHD3XF5p5U52rslHkE64W7ipdmF6Cxh31N7Tmuw2TwDJyU889gfb/0i3IuG1Kg3j/
ZX6fqTF6e3Lsvqjq/uO7GZQzbr5HRx0uz2QWLF+fR08NDLoID8o+cdL9GX+XSDnE5DAO0hPjcyHd
9r0lN992PcTn7tAuoFNR3vhskl+mTZ9SVxw2ruDHEoJhWPXNFeY3/n3bRdo5IpfLRT/VdD6v2z0m
NCwsev/4vnNOVn5EgAdpAX4blATHxZxpTyKWiIfP8gt5YsK0AIuf+R7XEEVq60LhXw7bSvPy7F0y
uRTkT01LAudPHO9R/3hn46I2qvvOgaZVXiHZF5LMPdBD41xbOm1xHVuwHXBCdEDn0OkjPLR0jhFC
OFQfJTT76A8Paa+uIZ0MwXdf6G0ECEgu67dM5oXW/nYaoYfkWp7kIXaCGLaEfIFBbtx0z1YILyW7
GRAmuyPAyBsS3VBfGJ2SF9Jh/dDfUfMMKXZpPMW6+SoXc+ZnQRG6JXNfZG01epAH9SnUGh+agR2T
WxTQLHT9nOtRVy6gvC1sMam5wo0As3dRHYKSHb4XQ2Z0vnbh/W4wTwPL435mrJhzhNlLWLt7N8k6
YwhB/Mv4iC8OzhjtDCrcBiRdpdOheRgq7FSbY5dRmg9/8cZtvSuOPBEURrCjUV3ZtjPVTobEPCTi
Vu/e1PkuOPrwr2yhU62F+X5zU2lP+DebivM4DKdqnXX1AOw3MESSpIYGPhxusbOPc0ydEw71Op3I
9GlP+Lu/eqhPSQX17XtD0NMbGJ2ATCOPXQBWY3SGt3j8V74L41JommLYp6YCTwtL9OqVrV4MdqX+
czy3jt2pXTgpqrrCKFNxuVN5pipZT4bY2RftrqrI8Z5+9osAtnC2x+grbTNffYsYN/rzfQ6T4Oa7
Qrnb5Nq3dToe2i07WvThaZ8l8Sc7rpdFb3B21ElSw5k4aWqdbmzzJRAa+TGI8Ydl1LTtLLo4LKdI
U8w33giNbrzgjBFK4OihCO7BV99v9Ve98Xy/XysgtWIzBvZC4VwAU8orc/bNVP5XftqqWvaBvYrJ
L+uHWVNWlj+Wj5G9Zx0XLx3eaoKa2cHHPDMSvkRk98Uqb0izjeAF0fqQwG7NBHt2STSMoy296aey
0GhhuBOR2cTrtHkjVSC0HWMRMfqTKM/O8clo5mkhCk7dLo/wsU1IThHh3RIHaWKun4/uIzmmdltj
U8G2UWlGhYwiKi5uFbL8mx+DOy54xbE+G9tpbvu4NSO+vCPr7UkpF9JNM1bn+Koqb+kvZBOZzhVx
OYw4Cb3++G6ixKAxkrc8wfGz0ec4y/vrGSn+1tYq+pmfjqkzEnj0fFQT9XnIiLIecF/DPkZ1hNB7
3lDxyGdCTEd1Wc99nIRHup6LFHSE3F5HKJgysAZaTteUI9djhXeFHha9FGh+OUOoNgAuV+BomKaL
oiTVnqpTVKeOK2p2gANBU5j/blVvy5SiVoo2O9wtlpKZ7HC/bVEEcAmIaTq2BRo9rBdnjG5w+Dor
dwT1yExho9OJpjsbFGg5AP6LevZisvJVr4eHe2UeR8crrB3BDGwdZ8IE3Y82XqoFWCmvryqhfuit
25ujh96OwZHI7jPbsuF1cn1dxqodxfeZBgtzFBC/CXLWI+n+1V6VpvASH8p6wQgMhX/MZjUUSgzN
cyQqBUSLhmUNXz8u2C2Y8z1v16C+8yojULsewwqbgtboK+YHtXANAKAF4iqbNMwBd3hnaCjvEv8V
/YClLz4Q/rUqknc1Ve6OPXI+hXmsjvoZsBfSsYuce1SaiRA4HQkFenTMR5hjfliqzTdasLMzl7px
eeDq+gryauKLWX6SR6ue8VoxODqyG3kjfPlv4S6xLFV6DAb9H6jkbL9igojSBlSFy/8LVNeZbU79
r4/FGqhvU7dthlLyowZUgO643IoR+Ljr94F/e+d/nldoq520dQ0hVIyGy4jXnyyGZKiytl0rrBK3
CxPGfxmFdHK8u4XBYoSnXWG8jRZn1XbYgaBT5ODn7+d8f4Bt1uK8tEmkq24sFP/heAxH0jKcssTS
GWzGIDYCbjXkHIl0YA8NodgJshPciockmsrNh8X4fiWVZLOEMIHdyUlXVivp+QlNw9gJK38ZhBzs
FMFvX0S9hUV4QdcxSuzp4P//tJ4pIlfcwyDvpQvg+LRj8KFCISWLxTOxIWFMyYRWAZYSqGaX+hKW
hR7GoVhDIkhqfgjoh+BgsmwgtxiyuPFZahx9n2R9qnO5bg/kRDvnQBctoIna1KkP3tud7CfYPmmN
x1UugIPxXfc6IKoIckypwl11CXG6GaZjXCqjD7ep3AK7uLXvKZLTPuBlRvQl2pBcZ3LHOvPsdd1C
qr2Oss0nl4Hqj2RdVuti2TzVAluhiZF5PpZB4zVFMMRYEhG41Kzsp502Xlz6GYwRyfzKTNaLJWZf
wxEMIJy9uoJclclnCNSAtFqiHhiFUIBqce6d6uKaeNbYEwAoB+h9PVMO0r4TYFvIfLDfmxfoPs5H
aCkACzLrJay313OVBKv7sZ5w59SInN0ry/rihXtugKEQY+wDLPJ8JS/jLTXKhJByLP9p1tQGj83m
H+2kb9VG8qcqADJmM4IW2TxoEF8DZzigkm9kSYFpicmZNdk7DscQ7GxdFCl98ehs8gbivtVGqkt2
tnTvkxzanNiW70MrDknmTWWISQp++FspOisSkTl5ZDFsKvZKHsfjfGLXxgtUPNjtWoprmsz9YY8i
QQkRKPIyFk4tDZo3wVcsC0GgtkorPbPyz14XEN1hYVQZxwWv8nyo+BgR+2dSmnh/6KdHAJGpCKqc
UPRyXlfQE5hdGMjFkhyoYoyD/GcZoIHU67gMlcccnvC9pvQuNlH0SxaaP3+sbQAWqFVXQ6BciNMu
aW/LtRCL8cVyafwdsbWx9q+QnL9nA84JeA5vJTwpi/yRJyWt4rk4RQwCJgen6I3dEpfB/xCikd6G
LvDO7RuqSO58M13WHMCMSbPJgaKAbkcda5YNOffwAgCDi5Afc8c71id7+lspBpBlXR1PXxU1+Hcn
pdE0dLYv/2dKsaDc3OBkz23rW9Trm5TN02B+wy621TW0ScJG/DfGIvgxEScoUhWHPJeQjtqym3fx
GJ7KVt+UqsqSdYG7uwAHT6L1N2lztL4tr4X7ciAlbfwbZWveim4wTasgwQdWyVlB0NSTACwG0Wqb
H4PeYJxy5JN5JPiScCGX4urvB6FUikOpmGUtR8OKAyFi7qMTeggYuHts5c8dTaYHMNv7tanN4ifO
gBoTg/7q+kyCVoRYJnZVez2YfnxLq0rIn5AYgNOqxxfOx9Wq2dmwhxPnWYTDYiViDUhqRbDqC8C3
KiT0itNX17CCcYbFsigH45CrOAaX2Ij8ieTCilO8EXm+8lW1J6mtxYIB/M/tbI0uromV22O1laKW
9X1p/JLYTHO64Ve9CrMCvJv2yD73Lj+NTX34aIWZVuSYg4FsbsGqMxb9vEc40W2gAka5s6XzNE0w
AzZoK1MEvmgFsSpbQ2rLEbTiv4rwoo/5sNAM+hXUCVmisoTpctsKCCQOxK1r9lMhRDgZSIGCqSwI
cazuZjvgL+QDiN9+KElNllBLohBRdiD+Pd8tZVSST2Gv3sjxALJS9FP+dvouwnTkRaisN25CQrV2
8D0ltxr6jew9yI0Rm6DmJZ9aWsyLVI7jpKX3wv2bwwmYkgJrGjIoSPdcSWrz9d9nMQGUU8hu1KRa
VBwZyN1jeG7N6tTW3jYMrG+cKqtdcfAghq6xozlGo22aqLfRdLA2MLlGWm9xXEPgmZgET6FH16fb
G/bbGunJMc5JS2wiBF9mKG5yEOTvztTOfxQzkFLtDmli2yZ5NRptv1Ld792aOw2oWSogmgKGn/T5
eg6A1fqYXNDKJ+w17Mld8jGbmDRnNldWLPKBCLY9XzZg7v7Q49NRqJ43B8SsBSZzOkM+oOgaaQXK
+5LBZEuWdPzj5WTFpF2No+ZoWoIHBPvfykoGT6qnCKeYSaEFmx+NBM7Y0GBTpdcs5X8TZCpOnASL
cHsvmNbWnA9yBSeX25fu5zcAiB3mxLaji0urh3DR0V8nL0R9cKgttAMtVo4AGezJDYQxSlnWfCng
rz/slKMy7efm0/Jx7C9nL1EJX7c1zR0vxGCAubcHm2WErbYrnSTdpBB9sqZS+1AFqa7IxxZ/Be0H
3hrOqu3kNKPjTr5PvSvXY/eH31tcKcZO5OgfWcq+QFK2WfM5SudR6YCoDudjWp5DMRKA11Caya3p
D1E2QFCnbU5AkLKIqT+3VquQmmmDnw4G2rvxqeZYSjgAEAYAQjyo+xSUhw2KXqIOoBR/gySyBpg/
TBu/Fe2FF7a/9qU0rYHyroSAazFlSMnrilbSywC0vqlKgizpTt/WUp4iKsWtI8Dp/bRQOy2zNr78
iBuF9PfRoAzAUtXje5LM3UFUDndqh7E+tNVmvVmeRCU3YquFIhrWdH7YIbNEJ2AOMdXc3nlDQP5t
WDxaRoHcLiBbIaGqfQTi8UyEDnSPFEPGAxJi2nWQnpgdpacoP4tctbLhqnNxmLp1n5F/bpMwMzTp
oeUg/D5EH0xQsi1UGLQCSXW3iGIK2LIX/Vn5UhtKproATVdShd/qBjX8GzGDAQbbk/kEYfWdunBv
FRG4Srwx9SSOIARck0uvcPeKU0ehQZIWwadZIcxprxjR3nJJhb9wEjoiI4gwaZO7Dey5zV1wTOnH
r63RRbf9BBMiWQBT3apEyPfNvfb53CkP8N3Rzp7jrgT6lu0Pt50IolXQpN7+f5m/7NU1bSl3mhd7
0ULWzll1QJ4NdrnUljsIIFgPGimkDaZX1wqRuAcFUsLRxbgUCmZ2XtburcDKDFvWaE5ypyAiD2HJ
yAQCthCf0WGe4omZ0ZRZdmCosyYPwHjxKXUdCsCaFeLhKYyB3xIZvS1mL2n0Ibfo/2b5s/jYDpV9
zoghmpV+B9RAQoA7QfHHVRtHt3tw/ft6Z0vQcOk5sayZCEv68SyYdxEVaF9ZuZsTQM4hiO93Z8u8
WBa6/99kQbyVDR6kyEH65WcmeQnxBN3mYIrgipfPbs0Yo1qUhVHHR+F+m6i8ohCD7Cmi63pG8xA3
nf1a/9epGfXXvmGVccI7HJ0iTGgepJg7HgdnhASbyhivhvKM6WzNIwzWta0oANSNSMSMLMnyBq4+
MVwmbaD/XloG/krKp8YBYGUtqck9zzYnupDbSRi15IHYHaeNyX0xWHPK1VnOswErIaD7TxFB360W
jrpq2wyZfCBjruI0b5TogySwO3PwAIufHN5gjV8jBJhglbBZRgI1vDoVDH+17UiQOsVzzsGp6pFp
R6caza61904eiBnHMxQ68FBEtaJ6zQM4lTPQCudy78mRPxkOt/kYtFMjigYp+nLM7AVaINmcufxy
Z6Wbpl1n7h1tHmKbTjyfwekxYECbUsu5W0+2XecE8WRQFc5i/m16EiytzRQQIh4XW7JZACCNBAAG
TzHW3zj3WMzJylD/2VRn1WT6mqMkYMqN98qGcPJGs2Ag89pIf5HtTszFYYXF9ln44CO7rSWof1Gb
HLtc7blg8ENcyL/s8UIq8Y2HmCjekWsO6dzrbSoRUIrNpeGRUsraGT95eJadWkPQuYeAnDGQiYPS
iuGMJl47gohymzVhNXAjKIDGHuQ8twLiXkIy5xAdRkYiBKeOpP53J5+lfwWxvYulqh4tB3KB2wpZ
meQsmPfjwNQ4oUjxVoHOgR+8rMQ4R9WvNW16YPiGXmNRb4mD+PcAwf1+WFM9HWx68N4eqP1L0np0
ozTysupqV4BGe8icQWhGAfCjvjBgfaiBsAE7wm9vznx5Jv9Cv45msHPAlLSVWT5EIbiXjHQJq3J0
W0IRMghqD8MqFAxowgJuFe0/9zh3MPtSeq/wKIT0u3/M86R0FSZhZ0B04eg0k3cJHr6L2sWsdqTR
uAU5Al0e4yXN4fr2Vl17TQpm9NJoEwNEP16PQQIIOIeKKNNYq6Z3EeAYGN43wsOloyf/sWHHoAEa
MOCcUoX/a57ANCxpk9RzXnoOaNPIFGAEdQZ3iXU2t0FY3gtI514Ak90diL628biHSneDceQIJ8Di
yoDI7b237seQUB79FIjFgOhwC/UrvT6xmsmCV8+ee/ktGueGIYMAsxTozBqI+qNCwcUWi3xl3zyH
nWMqnEU3P11fFpaEG8X6L1unaxpsTcsZLe+ZyI8i3Xxp5Ul1t1ru2G5otvuCf+JvOZVOs7KW6EaA
cqkhhzpLGGUo9rM1giRHrZ0+nUxBJNqBdRLtwIeJxd5d4hDvQxV6BYbV8lM51gCcjh+NaCGQY7mq
nDHSdyPM/5AnWZkeOA4rqbaVQITgS2TanD4fwVFNjDJEe2VEi8LVf39t1ocRXe19z0L7XR0ySd9V
ol1fLczzAVXi3EyCQqCjg7KUqRO48iMLSHcFbOGIMieQ4yc7z0LUTRtXxk/PMwCctRBLpJCiTJGP
22rBBSI9ZJFCa5n9WgDO7lSCgIZA9HediHRQwoH9Xf1GSvR17jjZbUYGIAPsvwaS/UISdoja8ekv
QZzU+bUVoW/H7YUNvhgE5gNwemp3Wabdpcz+wBcUdlexYGbGcEELvi0zBTiuDcXMD6GZmMW49uWf
UjfnA0DECICz2fM4CNYmbFCMvX8OKEgH5DA1hQ9vJ6wqKnL6gSiz9cL3wmWdBKPTJjpt8QbuHLmw
4BQyMqK7cfjmZvvbC/y7KokYV5ohUC2QrvqkQapcNUgpVVa3AGDFI1O/fyQZQXELE0baeic05Aor
Xm7IlQi68SaPKktIIPm9Hu26sAl/wgduFfNhobFtzZKKCNtZDp02Bu+RTE9Ek1bofjJmKBPkpUPO
YukLG/L4ThYaKnHLBEqb5assyhinWEDgPQSUaFViOwHewqV4ue6ElmL4MEOtsvGw7Tj+WyMUiKiR
efd8W81o+FHupr4WL/YI2elo0jOIxx5LjIDb0VEYVeJgBDKFD1b0zZBrFiZji87m2JONg3TFhAXy
tHVCkEKI4QhY7DNwdCOS7hJNjavKN5waHAmzKj/qAJzyZHnpC1R9LPcgBdl2FWW59aKXDxgOOg3V
gcEtHGt4GBQtOfRrfIizxmAYDT3vUwKMStwhcb/srdtwdUT3ZPXUfrNysKfbItHQyMXJSm3eQxQ9
S/AHtHAhrVfpbxgw04/yS0OEIn+eOJ0NSXuKypGA9svoWennL12W8dlFdGw/L1WOnhD3cu2w/hjQ
mECX0TrbwG3788HkqiBnBtCttRop6c20H1KY7343Pjy3YFygGnlxfwa2YHyDvHCb+rL2JoNSO2IF
R3jzN98WhWQnnHIPUp/jGA96CeFEWRjM13pT9eKJFVhqtrnBfSUMINNj4ySnskASnVBxHdNYuLPa
mBy8Zq4m7sXvOqdRB4OvjwVC+74O7tcXl8AtLrCb14k8hHxM7f8WVk+0BPV56Lwnypr39WYOo2sd
adQxmNVKZubmX3Ut7mg+gm59pRqXnBAY6GWlE4sIGZxt1Ty/jtOEAulyqRcrij1vRUthj4QrU0bX
zZRiZSeFufQJAXkjlTiu0MtmyPl8MyS0f2AkeIkls6vA1sHDUcvlhEDAexkVV4+KG5//MpcY3M+P
IOdP3wnLsXmyo2QnaEwpp6NCDLfPC3aQMod2EykqJuJABt0SLAl/SOJsm9zjU0PQrqoxQEdEaLlp
+lyUwy3+GQAMhGJPbaYnkkGufYh7L2R+C9iE+rldKAEA/E8T7UToI0sMI+fgInAD/BtfIqYyqUMc
G+uiCdXmAi3pGeW0N6GfaBY4kmcs2ifiaJfwhvamgDSnGiPbIrirMl4VXp1j8Qjk0ouTzfEe41wJ
RfwD2Gh8rqnZEtSqll4rDEDrvyYnOeGl+iXlt90jYCgdlO6uhbIP3sXH/gVpnNPGLZG0Yb5qyM5F
bLpGUCPZFcy1KPCXuuJpn81HS8Xhx2qHO/uPmjq2gf/0OqU9VaMDXdT7iCouwUHDtdw6gmWDk6jJ
DGJA2Q4jKwLTKU0KMgWKpWczeFu+c79lKXtmiFfmdE8o0tTdWX7QiuUn5MkHgy/GWSckBiiX2uC6
WlAZn3FTm3Fp30dJqSRYSGegXdrM1cEo9mYCC5CpKri7OuRbohwOnNEK2qKTUfkE1l7YHYzpZE0A
pK7le+vF+a8zd8qT4dInXOEKFlDlnJQEsEcKV+4P1DJYLbayKhp+Aq1LWvlyC1YmIItSW8RILW1X
l6e9wW3Lsu3mAC73XvIpIrgvOffo2QWu92PJwjDe3qOYUjH0WhlmU0W4eenz/48TaEh2l3gYR6tM
t0WzKU/kjcncUNK4fP8nu3gH9gS/ougwqPq2FZeb5KWTGPa6X0qPWV6d1XeIJYNj+7gRu6t2qnSR
nEcK2nKFMyV3GWm0lBh8SvA43Gxdn3ah0lFzppUEx3YkAPfEenyayVqjpsqpXBdBl7jubhUiGOCL
xetlQx0mlBTvLKPwyIQhYDIXnMekdqzGRA4/+9e7NaDrNxqu5zyShbeAbE4jVuDsQTxEk6/g3ALl
RW7l+lF01pOh65UiVLCSwLUHObcwmUFk2XhI2jaFsS8t6m/QsEYzHarGUTLzaX09Mzp7KbSSJFXm
4WYlsofviiOEClr6rt0/wysm2lb7QxMXjHIvVEcC75c4tjLxM6hvcQ5owRmRRtZcfo9oAxhRovPk
HU8ryo8l3OISeJOB4zJhowa+u8TXSv1KtujIgEreXeTKu5UNXdFG83PCgtmDdU0t2Tgemwl3AJEr
W03r6GPD7/1XNsBVUwQ1QuzROUkODr+ZiR657gU00rFM50WuQmwbbJRkdU3kl0QhS6zcdip+r3Yn
DnO/ZjVQ909n0AqFdkA6NOd1/P0ZDfAOuybqml9Byju9LI+zmuW98rujt1Zy4VQr23mS2LlaWfy8
8vjyi/tC5ZA3HjIC8V/ly5s7FgKQ2UcrQPAi59jk3DMIb46nkoCI5PoRZ3xdCraFTNTEihcBYFRn
shp6qBBAh4DfeuNsVx4xYqjNI78hwCEgDYlBh9j6Hdrovc9sZrRf1Fj/hemEY480UFd6+2EV0mg3
7spg3Z34rkRuOjTCgiLYXayrLF8EVCHWmmgdnbOfZ3jpauRI++kGP40adMj4jwieHmO034319TiN
Kwu7Q49flINA+cPylJj0rWaszcYYBTz2JPDZ5V8bK0tkS7BCx2VRzY9FsQoByseyOFo7AjemzUaR
ARaOFCanF/+NkoOC6UGq8+hXyp2jIz/nHTDBPH6zRXuytK4qi69L2ZKD8ksmi0xYEUW+M87S9dy+
dGK/yr04b8WsOQYdpuz4apyu8RlEekaEGBNUmZVBSTm7BDCu65RgXH0b0qtnVny+dpaRH5mNJdxL
hRMF/5obX++HdFrjivl6IAnnAqWOQoRjbtUrF0ap3ElhFm9mfM9vST6RprGAz8S7eOMUWW/uFEgN
YyCz50A5iIUPJFrgUedWEU7IqSJyYW0zH0DRJxDDMwr6dfTscz954771rN50u3jxXLJwM5WtZWXs
jo+L7enzJCrnxMNRTsISQ1zzu0RZTlBD/niwSaN96q7WMQ3pZYI2jDup84aeM1U1easNYeiQGR0X
bibk0xI3WWeq9+HnNcPm43wpSbBmKo83Bk6JUxfIole4ijvhq7mLDXM6zuYg1dAohZjNodnvp/ex
29sor2JsuArf4k0JEuA9jPlvjkUZO5xzreXK8t0JxtzhEF7Dkc5ZwsPlf6sAfVT7CEMfSRdQt764
Ep9ITUGcX2gR6lg4v59JyCMrjbIlg1WSuVNlwUUOcaO+nhwTeMyckIpZRa/PxOr0u0FOvB1OiKw6
ABATUetO658aGKlTjMHSZYSh3I1pLCerLXOlyEWyKw1jhmW8DPB+c21ybp+QDfWVQ/MR9HuXPdTT
Wv5sJYR5ZEOxaicgn8mZvuu94BgsnloYadGTrn4BLL3g6lHiSbHP/dfN/oJcmBOignF5ACH+eFQp
bWVxGvvXWVONGTxsPYbylIACy7ZJ1Go7C7oB16I3PKqZ1bLyfnwNjQ0lPXGQ1PrmBPXUwwOBWCoG
8wi9GapvyZIs6bKSmk814YkSQXZQd2MwZqqftSY2aG8qMPxqe7tPWdkc8YGNqinpROpMx6xqCCrN
DhsOizHaCdcM9vllg2sexZdGq4kGCnrIbbWZkuKlDQ1pcMTm4u7+4zTzX0HU0l2XEPod7ENaYK38
+Iliiv9Uw99mZ8tRf2lih5rzDRWSaVaP/cWfeoa6zUM6vwvNpUOwiKXwl1s6AB+sXj0WxNN7Db6g
G60mcclioSnmSc1IIzSQsLtT5sZ+mU5mnscbRds50g7N5AHneoXbbPRBtQ8qj/CdZYlvoBNK62Ed
JcSqzbfzOgCJjxzZBNebkse67ot0z3nf+KLOz6T/nAyF8hJc5HjIG+EzI/oXQ4Yg7hgObwLcxJbV
mzuJaiqi83YIFCbhgH0qtXpu+c0Ko6btaS1MICjw7vA0DoYLvcGDnYSBEofiK7K62p5w6HSk2S3O
c+hvY2Vhvi2niN7xkDOL8ev4oojZ6sVYH8WzJO4B4jepfv3v/tQi6YeZJXzYpM87I/tNXGD2DF0V
0AzVsa25cdklNAHiCqpGx6mY+5U9GzTvHWv+H/N7icokAPawqMBksBPfhbfdU7E9pDNrSKGLcdae
MxtT8amX6yyN7mGhX53RITOgZQ7wxqYukKy1oPMhtWvttShHV4nFw1LN7M32JNB2nypfbGevjXec
APqwANjVGv2xRfRl3x0SVDOKDY7rCxRDz/Sq10dommlQ7exRS70jUev8wivAh1x4Azu5NpYSJRG8
rLS2wBnRHrr+Xm9621R0HZbc6ATlW5sr0W+MABAkMeXSD7OSZQD3ioKEXYBkTDIMHYow8c/LivBX
hqcQPWswLpo8UFH6xeWlheVk02laJGsWNv7CdwjoOGEvqhpykAXJM5PmKujWdAtAGgCqewO7E06w
L+n+ImSDRNApC7lsID94WlGaZFtCjg99KD+W57poq+v6x/STa7YdA0YYJkI7YadY8TfS83m4WvNH
eLMI1scv/0Y7+q1fO+ChnY0qE5zAIZBTpJZyWUVqdwCcLiNX8+m9ZGm00oih7qghCOK2h3VFEcey
2Hivygg/p78UpUGpIDf3bJzqQojSk+LQ5DyaVRTPseJ1m631PNmZem2WX5PJVVo2l3tEcJkeP1ky
IqSCsWQqXw9sYimA73sSW6OT5ymX/dCN10LpTN8es+WUVZTwsfmxSKgYfJQx7vCqTEXxaG/6jAQ/
Kj7FGNxN/qCSCovwF09D4w05Kr0gUZwCp4SaMTpcU/PXQbjdEzBh1j8Orlh6ADQWYbiMu8jGcsHZ
2ka2GDSnI+FBqBXXbjdkiozqPUS9TQJTG/8ui+HVJfFy4x3GN1RKBACfMqt2rLOfqYkjX30SFqV0
8T2fuLgKvyItZx4+Adnjrj9h/lCtQT+L7JxxRyPEX53n+k2Jrd9N8fE14UWSRr3owN9JfHOIozR5
5bqMsmWsaPCEh0Kr2x2xj5wHtcGwY1X1Vsbw8loz7k2yTNmvo4g0qDIoaNOkeRrwZWFbX8C0GfsM
iXKGY2mQyb82P6gkF+dsZGeDTAQiBl0AhjIzORPBdHoDPLbD8v9wEZqgA3zI8PVFHyuK5iYTP9oh
FmXC9LWA3TdtN0pPeJsjt8RXO9sEX7jreNakepMkhaAOtsJ43N6dNOpXeGIds8UEis80930GI5Om
xaxWo3H0og9mhCe1bQGmWIkELO+kmqLYQEKprDt/PdEO9qFtwHzoUFBAXqMxQSPfNcOhd9jIB0jb
ygU+efpDImcMCSEbt5Mn6SEQBbYj4auFoocGa4PlHFSUlKVrhcyQLKsEnm8bbwxY6QY+1CnvOGmD
5Mu1Sj0DpOHjmrm1zSpS+p7f+5Iii4dmm9E7dPlGLLSSrqoBVu+hs8aWzxUL7TeyszqLzbMMFtPe
TV7BVDrzsxugv2GUb6hX66bWNjYE7D7I6P5pn0hEqDzsdIx7rVS68qzmFkSc+xN0k8hP7i3CPOZH
H/HdzOorK7g2yU4WPPP9j1v+V0W4fq/Gf1o/Ldq9N34/7ffMalNsqOFwIZuy+/ilbNAgD8pIA5sI
+xDA5C94ZyB1jA7n13fPusbxxMZwt7kC4uqj7qJmdcmaQkhJ5fPrBwnsLWgrqzxAEvSm7GwT5c+C
XSzqWbIaacO1hAfTkW33g3BOTjMFBuG521LjGqs0HpObr7ND2lBqXi5EfIz8TN6M9s40fPtI3CUv
qWwc/du0pZY/rz1Tu1PN+4Fzl27Ytjx2yBbbwPnHifPPIFRjFasvA9LfDmyam9s6n2Btd+y/9XHL
I4J7dw+X5F5tH1ZD0GUAF/4McIwFTTG17ngRcqaCu3F8CNuHaTm30CkTK3blCyZtYtzrVdiRgOMu
hBqtnDyqllGJM5t2kQjQrWxZEnM9tBXbZEgMDDcpQTZpV0Bh0IEJARvSbNuozkVilL7BSNQjFg+/
YBsEugSxrAHaPhaH4XK4o9I7Mt+q9sG4bfgm/aUnYo3aOdr8yJLVHeIQJirAR8tVelqlaJQHH+HT
WRdrEulWB6rfZ6WJ1JQgU/24OxnxCz5LtZitDHKeE0SzqqMF/7BcK3/vhHAaJR3HUZkq4B9glKCT
R7oDBquplg6/O5MSrlXygxqjdlU8CqbDJUKd1plrWhp5HsCa4uivvuPS/fuyPQAgTq+iZCLuNktc
sHCZ8dTj1UreijVJawuXqdR3oeb7kawHf63IaHhumHfc+GPcFkKjVvlrgrVcggKZPwNsvm1eKra4
PxUpiNz/0foya5azTLUbf4pWiDzRN58Lu4QRaP43w3eoyrZ31mwvYa9zNvoeotYEvQ39B/C/i5U4
s6QxWyXJo8WZMmXhDeNHoKhmIT2E3xW0KhGBC2hnqKxPcKV9QVTIhbu60jkFPqyvpG3rfgKdGOHZ
z0q6zsZcIAZWhlSMdkeOd1WFlQJwtdUwR/k1ZR83ngV3iroxTa2MR/L9lufybRLbOuV92IYcmji4
45inaHzIs3wvVr6bmBApx2Ir33rdqallWKepjCjb3GPTxMGBnzYlEV7gMGqUEJ3XhjgbuZTIInH+
+9/F/Kdpg3uayYNBN/2PHCqTWfC0s8LJsRrePwkHwjfqqOjOEJrNnlRPsUD2EiEMZ/1L8Ri99yU7
QovuF1fK47Or9rBgUYq0yZrNErRSsXp84vQ98d8Bip6xkt+unEjXF6yY77daMAGtw2PdAdx8dVuT
3ST+gdsXmk7surnwp9hTIPXl9pCZBxQvoZfyeF0v6aZ6cTvOl5aws9OCj0g+AaivnikH1F4kitRx
guNxHTvh7vliciRtv1r2iwPc67V5mTkWx9ygvQ7y0jmTNewLJdUc78WBn47j7uebl1wEpcL0YdKa
dG506HVk99OlQ6caeFuufyeMXd+kKixggeGpdLbZ/spC5ND5xAs1Pzmc3YuggAmrXOqmMZcDyfMu
wQIQb6SfBiLRh2/HzuIy7fsLDzCbgAq0GyrzJaYqh5ld8iaheyQmk6pPut6ZFRXrbbuBzhVwQ2MV
xGqbuevS6qkLcFNKnAex9VnlIr/unv2OWBeMsXbrs/lRY2Vw8/8qZ3G8RXtFXb2otxMZcbjJt8Vj
DHw7jGs+ViqIpJ06YPIxHjOdMotumxx4HUerq+VMax4p7PVCK99tEUHsl8izV0NnTztUIqTjZ1dh
e6id70luHimK44EDflomZfXilNxy3UXN5gMvjQll4TkfK4Sj14XnQx1JLybkPMrVtw2JBVdhCadt
+J9SQz2gTtvQivWTG0ha3q4aI2rU5jlJ5++NivXMHGKDsg17fGqfRoRbPWX1Ng7JKScpddnuQg/f
UCPDX3IHi33cvkpnBk9cPTMnTx3kyPuC82U4ES42Nn2sMDMkxWx5HQdyf+0ncL6a3WjenYZDd4/r
+816flStdaNlKBuweLkvFilS164XTr7CWe095wFgWI2ItwHCXWD2plw3TJ+lUK9NGHd118m1xwfp
W7svMnc1rakT4NmBw2nf9f2dqRZA18J3fNGYkaKQASJGToQMRtfIOzsecLDGuO0/YRDpG7sh+113
DwL8Bdx260GADiqUbjRwtiEYh/aF3vOP3bjMbIS/zCuRGId4cVJlhh2ZiZg8DlSScUruQFc2wJD0
eF0oNlkbX2puNNzWuXKh8jO7tV58fBTm6d3vEzuw4ssq3OR6x/xhEgEZ8ttPcArP4c5KDdnUhSeJ
c8aeYka4cu9AWHv/RvYJCxEmGJCfpROZp+GDxhGz42RdtdH8r8DVQDsd5qo9Z5P5XmzRoVzF6mdl
5G6uuHAA+NfmZru5x/dT2mpOWauevRYkHhnNx0CgmqymQyI9h12oGWvWEXYZGSiInZu0qV/FbKxo
8h07rAAaXPFLbirIOh+/uQj+RAqBfjfnFtxcY1/leSyP7+dN6k4yTukE8f5YH8jqDtDRwqW5+qZB
tHjWut5Uhhenm90jZ8uq5SPFygvJgRGCWArB7ad+ko8m+FM3nIvDLpEvvTTgHcw6oD7fOnx3Jh2a
EDt12NcCXBjHE6RL8JrawvoWmZZg32x7EN0VIlrYBauN4uJ6HUuWaFNwOFkgoIlQslCG5aw3ylsN
CB7bsB9Yef+f2m7PYiCzafXmdwpnCShg77R2ObnEbDcbeERwcO1VlE6zAjsT5fmPYFXlbXwD7SOF
mJvpHxdLDH3tvcA4eKy+s9Tib00v4pmpeJqzwqSInx9HihiqouydEPKVFzlYqUOcWlL9t9SMZWrf
FJ4D7ZP5ixSWiN/+Ess4qwkjNAzcdtWCb7mnFAATiE9H7tlwidcAGLc2xeYAqPYQvb2EgcSkkf8V
MN4nBGPxcSm1Lt97pKvHzJhPr8jHloFcYx6cvCdHCKuUCfsK2HG7609Mw8HgihCc0tuYHdki8XdF
WILQbS3jGmYbRebh5oJpCuaGVhDRbj4XEn11A5+qezDs9VBp+hOQgIV/du5+zScYkiBTE9mWtetT
5ZA1cYVpfXIzdfK3Ge+q50aJPoUVFxVujzfdIo6lcuFuoqWQNzLBUu2a9QLFcUxnS/hvwN7x07xB
rKcRQV6nwx9Z21OXJltAvoYqkDsBorW2HkLSG/YHaNG1SpxKRp+6eI9AZ6brVDPMO22oJJ4aL0RP
tfeFXlRLK7J2vfA2hp4coOAn++LO9BZvMMFogsvh2Z1/oiuzcuRNlGdEt87LIQYxew8OlhAHgXZ1
spDNYZf8WFJs62keTEEtkFSfOBUxpOKsSYfoHI67GgItg8iM8IVfyh/31c4bRBiOT5kbR9Cx47+o
IjL3Q7x+VK92UlijR8U7eTY3tvzdYJLu2jVDbW0FPKdbxZ18ubxNSgSjS3q3qDZz09Zq9z3FCJBJ
jYUBdSRtFfADZUbIh3idT2pNI/yVfqZmh9K3vEF6ltv7haG0wOhgnwXOgG39/GwkaxoxnTODjK8Z
qXJ+Xkv2eRdr7Ge77WE3sL+bFl0x1H3VKcjC1Sv9nRM0QMlFYc1LtcgciNv9Xp9Jh2/3eXHVYoHr
fyiLF7/GHoZ/kCPnpHOyul1rB6UzGsn2/qkPBhm1n0rfFyvRm0IwLmacVHUNjm3p79nDjPROUIbs
16AJ7IynpgMZyhs9TEczM9pZc6TStmhZg/jtayZzguNH1bl0I1Z3PXv0z+UlGyGLmG/MKr9ttGmn
7bDGJq88doWc3wOgg8eWMz921aOknlw+n0hltG4eteoO/RIcKloIsgBzq7ueynzSj8Pt9MtnLTwn
/eg6zpi07Zy+NDfJ0burWawVQyE2H6cJ1i9FfTw1d7hYb7XEjH6UXjbLLgpuZrU7H2sxzYYdENeh
C0lBDmNMUNrQ9y/+7vWya954iXekop3X3OIHgrkBUBmpm5uhaU0S6MN4SUoTFpgMYl5LZHM++fkE
tnsp4q9pA/onSm63KCk6NR8iTsXyoOErIlEU2t4vJDNjzMZYqDSrNXxF/DssF2yBtUfipO7dR2HH
sKltjqoRdirJwFp9wuGzJw0ycHRUpz0M8WvLaHFqSrCGaCXhSyzQJ4yA7GaWORAjdazj63jVbgsj
izUzvbO35EnltWf78/BfQWS9d8Wpjbfqo+FmMq8viB88PJPpSLwtxpoFE1joNsV5kf5fOMCimsiq
VCV62ajwUyH4K9DdSW60ZdMGLxPGWGlQ5XToF1TLItBgxZ7VnitsTXoZfm/er2aC/pnEZA94SaiD
21CHB1/cUbZbhKY58aVTYjS+ILYD9F7/gYA1PICuOflhPiGDCkcrRxTNL5+g/rguiWg4LC9B45mj
l3giYsPj2/nJEPhXu64stc/iXZXSqoKHOHbbfQgaD7vPjg3y8ZWHVIu0Oevn8FhbyDb0QnDT5LCU
as6iIhWXpnxhAhoijMbQJZzZhujjV4RXjt+Tkgdy81rVqoIcfGPSKrjVjAJn/jH4ctfG44AduVGg
btGeYmklFxhB5Ij7pG7pnfJ3rZUdYbUxDX5hNpNxafKddp4qCGcRUcH44lpvwaAcTcF6BbTNmm8T
01DwWAs/61hZ4Jv8LXL5na8v5TYwOjhjgFSmV6npF3WRysQt9aYO50flxAxzWOZIJpjScTYO+DIf
omP6t7JkrI2i6q7yDCEfDydH5eaEJjfTKVGITAHyaHFiqcPGCfvuAOvgeICFPm8x97sLOzfFOGl4
q2GGkyF8NDGLn4qYS9wCTJe175bMFXp0mQnmLk8GIXHdJcm4tP+2PzL2tTfOEZUB7JLlMX3HPEBO
45C1VTxJBSMgrd7Ak/b6focl1bqbeQxT2x5helJ4AdR62Q16cOH8sCI4K/qj5ZCahQPCswmhAKgk
/QID2HbNY83Bl1cmr6nz6nBYSU4RdvXKIPUzbL+dkqstERUksP2t+sZlqY6Nh0mamZ6GzyZGA82R
8MAQ3K9czOrKL+QX+1EbwbbxDFj4qFgsfEfmWZxyijUKRokTh7Co9UEMdHOJhhPqhfroIXnQ0mv5
RiRQZPb99w7SSLF8hGxi7CoRNdAI7eWWq3m/gSQV+cr6GKu1WemzXHIslR2kpB0Vp8ieyqMEspR0
HVRkF8sknD3yFhj9WFGGNTUcRlA+fG/Vxc6H5ccJeDxgcSDZUj4JIM1Oa6B4Lw6uQKAJITlZ/R/n
2VHPA8AjcLtRm9Soj+9S2EcOHTQcFIB4zkorrQfR08hBtyYYEHXSMqY4a9aD6nYilzgOuc/boQea
ibrvfkQ1uuLWlcMj3YW8bYLejjtmYYSZJhBXrtc6Xv6av1/9lGR+VOLS/qNAk+qVQAYzoHc5erwe
B1BHPqd5toBPHbr1LpK1CXIrKKESVeORY8z/LhoRuIPKWkPiIc0rbTf4SCGXZtPtaoMXHYHovL44
kCg0qwe5v1pT/u5M0SWB4Djq6SkHbvMniwIDFUqGwWsIlAwPQI+HCkYEeRlHZuvSD59Gqu3Gcgyj
sTlRFhpZHC62luUO0TBAqnIF62+Zg7IXlJRK+XX77HMzIYXBSDuDCYu3X5Rmf0nJUpSXUxlO1uRW
56Er4/ULAyldKxpo+NSX/z2SWp9fbHuqhBXQAqb6aPTyIa5TKwJ9R6GQcQd8Y5M2VGGphXSmIRzK
waQoV0iCPRxZYA85K7lq+cj9a6KF4izOemQcYlEsq0SPj+uzcQExrTpAXcAQT5ti/mlOGGwvsxQ7
zCpouXFmV6bWjtchQaBbDElWZUaaYaRpHctOQCpNjREtO3L9K0uvY3X9fOjebrh+6DwTYQOHF1a4
drJsPRvb+Yeo5RFqb8DLkjXKXILZS8NUZUQirIVirLmhU1iU8B1jJbYJ/nb+7w4XZq+jjvJzRJcJ
OFCAgCD4Ld0e0IdBtFPf1KoTn53HqG7KtCXFbcwdTBNJ5fl2M8C9GmfO8vXIKQLDvlj9zjpUWZLe
7Q+JfE4sW7pKqO+/vR9DH1e7q8YER0FZQao20x5kn9qT5nXbSnuQNSY4o00dBjDL6ZFn8kmgWNKb
qSCsX16xNuGQ7SB4wTCMeo3zHyoCq9o+8GKvxWWtFrNiil8nIORiJWT3Oe/RLjnJaTTbXHjfIYGQ
j6p1JZzAaOlZGMnXo1+0kgvblnTIKzIOy11Mv7c6UwmiRqbXhQXcHP2f2YNxfQB3Ly+i4rcJojvD
fvXTtnaBVD7uYbmlptZubMJ1vw8B68lFDy1R89snR8BbJaOYCZ+vYggaulnfOmTt8VfnF2/SBy46
bGy+IXjA+yofX7JqeApb3yXojyDtsvK4IuBlyqn+4rOZpZ9Wzss4H7H1p9a9vZD6e34alfkkJg3L
Yh70AN9q19jc+lnoeU63Ifg1FIZNckMjy7AqPgw98aHnq1GxziOuwH23TR4SDryM7Ft1BXVzF7jK
NebznC7Di0GxZAXzv0ZTE9d6y8PMDC5ed2AwwkC+0tI8gv5r7q7YSjMcQUSxuOac2OUBAOX7j9AA
NP22I3ANidBaViyboaPL4Y5PoLI5RaxHdp2/vCXFwrPYj3GigqrMDny9qvkinZSCIPwCc0UB/A0P
1y02NXsjBQL63zClHwHt03rwaGvpQZ2V81v6IUDu1EG8wwk1SuVyy0kUjprzJ9vp+anAI6JGVwwm
3uZP5ruZ4AXqwVvDVPwCKALsZ8dDOUWjAayCV1CFKOMoGSVYB9b/xcgAPDmn5LrjEECFoV2eiUZk
bZfpKp336/i+k+8rKPknzl0F9BmoZLVgbUOxE8aMvSFXAFQF6ZomuQ+jzYIpWNpeFMr1AOLBxcIY
+S5AbvXnvlXAP+oIDKDta/0PpgGUnrGpok1vjsH0S2M2kk2mvypuCm/Xs/QVD17CasH7+BxIwy1j
vAbgkOhbIAE+eZnX/v4EoHZz4n+ru8D9mqo1xpN9gnH4g3OH89uzPlGXfXz7nsXgsnunI3aGNAd/
H7x01+yH3i6hBk/nc7ZcA1G5aTqxm6BOIU5zxzvuGcb8W3ZIGm1Lq44teLv5Ea9gZSDkGmEetwvl
fTcfwOkF0ia4H92UbjOtE8CtX3ipBlYyTFExwmy7+SZp2KoLxFWx/J93+SkMrorp1sEsaFJeGAGs
02E7htXBT9phlj4qzu+vlnSDA9BB5n+kTv/pWX4ForbMpzk2ULLIRCJCRWCp5Zh57BypVTFFUzZQ
C4rSFQVxPvWdq/OPHm5HVMFiCs6KWq2FYJ/GPj0a7VWP9lRkV4XwTQE7NZW4eniDbpZB50Uf0Z8E
DQOnw1VS+kSEb58kmzJ6WGt5xwigoWc8HZS9ttM1UVwg5PPO76hspVm+8asKn2dDto97Nqu6COv9
6vddys7vvCiOXe9/J/zLdB1Cl6s2gQUQ9Zmd9hu7O5NE2qYcZiZ0kGGmz8m5kPsPHHLD4ngt41YQ
38rx9YoNPdfn8+guJ1xqB/kb0EkcQ/9Lcmd+fduC3Czlyt8k/On2JoiXXdQRQBooKWJ7rabA7wrh
MTxDf0y+cJkv9j/lM4xzy2HvKHorvXUjTHoaHDEVLNm6xvoF6DS5G6cBgGW+Lm/cwIZwk3vZeQHH
MV15EpbhdVyjq2yoS3AWulU2uCSeldnMNEnzNKTWM2cJt/kEvbKGupUR2Tm4UforzIoETMazPgF9
gY47i+JrtVlydjfiHqJVUIJz7Vhd81w0hEpcnelRqMdZxioMX+AqPlm56Uuyo/izq50IsegrH7vg
Bl5/MR9/T6flZivb7AsCiAX17H3PUZbA4H8CeHO26gvCy+CzCv/DlBOiZSHqFX+YLXqVomYca0fe
ErXJtfzQPGJ2WkR+Llt8rGoZbWCGAqEGc2Y/FOegQE4bX7aYUAF6hWZyC9B3t2qE5/HXzl255JaE
CpEP9AqJFp+oac34cM63y7r4vV9pB/mG9MbHK46GQRvW3aeZ53OmyBX4Iffl+u/rktEP8XbA69ok
CY9SMIW6sOe6D6atlzJztYEDuOPGdQYjUbmVyevJR74wspSZdPx+5OnQwuLSLWF0TcxxUKDPvpUE
K3dQ7DQc6KS2b/D77hGZLV2XR/1ZM/cgU5moAkkefvwV09pr9l3YrrWtW3R2n+Jkx5q3Zlp+HUUz
7p0QL6O0uP6idyox4v0FB8zvVT/lH1rZNSsWGqGU3qVB2siTg6J3X5EmQSxJ/LW7zdHafcVd5Pgl
FXPPxAL5eY1RON2hXZ7gQJeVWbpQtFpJeuVfUCorywmCpo0fKAPWlFkmaHblJByBqUZjAqPdAEqg
YG75R2yCXTL5JeFGgiaBLlOyE1Drz7kPUUBInbOWYp2anT6IDBXnfGiuOtSvnEPAMV4EHpNvLaTP
fTr9Cys7kXa/y9SVbhf96MV0DCkbZfVHk2Z5hj8em+ca290rBSkULnbOC3tHaIK2GMVBc7gNxME9
xJTc/eX4bfQfBD8qcrdhNinVFjnsTn0ZOH+SL2nYiZuZonB1QBMhXI+8nOeoo92kpeGFkq28Yuv3
BTmRE9uzJBGjzHvKD3/p2GNvbLDDHjtb8mbFivYanwYV90Xog0glku8MrRozdTLRwudRMWb3z//p
qyiNNPjk3j5OA1h5WLLuz/S/rpN4zIIwpKbUwn9QLZ/fbtLt8Qd99AExAQPySoqZ3ufbrJwh3D63
VNSl13LwfBNcld33z1Vlw2+tCxLvKFV4gNhVdOwoduzWjJL4jNhGYtW7woC/WGVqibc/B27zmnOr
0tgBeoIUvNwS5HKKwlMi1FcL7V36lleQh9nmIfbS4I3/gCRTZUJ1FYL4VbeHu2Y93Lj96NB4fqBc
+yatr3x39JqVXJe2t+M21EiY4EohxaubkQzIaCP1MqaLmKPvSPFt9qmeP6QHmu272Im7TZpPaqpI
FCJs2WwHf1YJOwzm5r5zT5p5dY4N2YLS24OpJFKadpM9px8WBt/sm8jNsln7/j4tJxabdG/eRVF6
0gPzaUmpLzR3E8F+VhjVafUQVSu3DNjtaBl3DERxIBs0wBNLsCU5fbR0sDzAzym5BKJAwVpGa+5F
1rzEx4dRxDC3u1QSJA0g5Jof92+jYWcTFiPaLqAVcskbR8fYt6QTbwnEO0jn6cRJIOuxcOTJq3NR
lOwgGR+elSlkhUbEqLzyEiKy9stGaox+6zNXyK+KUBRGcJVXSz4bqeYDbS1fax6/oVCNnteQMKSw
4K8shUD0ybZBz1DIdHbR0cGjKxapcFHyniSblpsuy22utDXRtq8w+LxxlJCv2cE0PzLbaWV73Xg7
7u09O4Y4H17FIswg0az8V1ezp44x++Ie2x89tLibqdZVFJYBdI8y9ax86ZHvObbTFs9cM4t2G7Sy
IrqWQZjChAmPzwcn/ecX6X84TLirC5LkYnmMZjB+TVthqHYQ1oH5nGauCWlwyoFAkJEK19HFv96H
Vt4sml5sbnPl9f9o/+KO+PjfBwpOW+GHiXzqY+lcG3vWx15vfxE2PfvSedYAHaFDB9gazbOSBGje
gg2pdRbGXWEXO5QtNUaoJ51NVe6IX4sdlJwN0TbfTPViuLsJIVMOhossaVzuOXBjRKUMGyuGXUEk
BEy2YybBf+m+TEHmcp8zULWXyDWj8CqwA5L6PBCoZapN+O0NgrIaTxSgIEGaIK+eoqPT1KDB/aEH
RI+/3C0f9Ay4MN+yZB4uDfpkmq5m+GJxvvHYK//SzgyUvRBhcaO2wz/oifyabfEB63sbJxlzW1kU
K4QI4yw27JKM+tFv2S3IEz602VNL0a1+wWF3s6HdbDmmwmqd7CFS/NUrGLiZ1l9PMWNcXmSbAb4g
gHMF3hPPz5HbIeXpUYd8j0ERFTxw35BUSUhULdItWQ09sDHGYQ21SNv+t2uiOmdDcZi9oNe8qNv+
JJiQaSqgofmZWOqhz+vgWfeKT11Ezdk/o5M2fnkGdBSLdhK/IMEkkbCJdq4vnfVHFXVInKx6EboH
ZUvL17k8QcldfFZGWRhmtvglj/iy5Xtns5/3kn0UT+TCP+vmHKlJPmlOBkwNWz5Z8Qnw3BIqhniH
jGSYyLnVrA2iri2QVKLuQA5tbuC4NoJHKNEfN7DCYsUV/eRc35iaKh15dUItkoTYy06y2sfxioJ8
YaX6heNzQTsgq88WQRb6pbST8yBIBoQRWwWiTZXQdRQ8eD6CaPPLKjNaFASVSFcs4pzjqGB7f7nS
N3mzduNWWm1gq26XI6sTvE0loHIz8SLho4RcsJm6QnNm+88/KNGpqjJZ3yJgyaJ8AgDhaf7viE+2
m53AwU6h51I5OKElFa6TI9/fEyQXj9GYEOdiNmWQJtObNKVg5p3wTnBg+itOQBF5Dkqd4l/21gIm
OHSGe5s+33MsLpnWr0phrGKLULqAWJ7gZgibfMpE9aaws5bZdOvkRuayO7Lmg9QGe2dpsXM3Q60L
MRAqDQX9vIjvzx5jWzcdKOycZVbvOxmgLrkQdhztGUuMQIEb01WZiSSO4Yi8Ikj8t5CYVBsVLzW5
FoQXIrr/jzfBKNxSW3y4jOdbqn/MmhHRWe24Xea1YThDJkkUDUPwZqVKc9wHZvBV8TZj4NxUBhI+
JDbdGMXV9O+cIdXNzg9AoB93J1Lwwbd1qM3/PCHCRBMQ/mKoscbIDbaAWikZdlJjUNn3aSj5a7y4
aeTIgKl3ddVWmhCOzgmXbEOzoXG+Dgydg9gYV8z1eCQKSa8XYZYL7pdzdNn8UZYX7ZcyqpnALSef
x2MKKkfFAkpC31OkELkCDBFkEGKf0rbn6ERLqL5YBqesnJlVko6Zcfh/kU5rFnDf9xnAfPWNz2mw
PzTYV9D7ZyL+HtslFO4oHHxpqXpSxUehhlpfeDzN4ER9fJEhSvNKMdeBeGYfAc4+YuLm8cn+cBAf
gPrCEVRJgsW+62arEYUHT3MUMgj1JRATTo7rvOS8y8Y6UjOcSRJwE/9G6TGdVn3VWYmnaW4T0nK+
w16tn/SmytaBpqXfl72sko/s6y4Bwl2sNFHjp0y0lnURDsXxGUBUrI0r+57JNOpN0mFqKkFtDW79
mK3lPUOEKUn9vybimghcNm48CWa/9OYYjxvvqDl2zRdeyLQpvK3+D6ybknJ0f4kWNqhqOcFJUrJF
piIRu5QzDWfVBDljV6iH7MNobTlIeKCGcGmFHbVKLzOwbr8aDu68V8Xj4LIkN/PqCbip4VjAGn0A
HDehN+PT7PYwpjY1FZWZqrECkkLv1UOHi8RbAqOCwbK0e5ZKnGwuFcnRzom7Aj/4fUOBZa5bViRZ
M7BimIS6Rtxrt6cf41heJHbj99gYI/Pm29qaiIJpeLhg0acNShiTDyNmPXizx/xTEkXf5OBQ3yJc
n+GaqWDxF0WIv8WUilKZS3VU6u47zZn3oIfzBUuaxDSo59OUdFRsXm+H7SCOZV9dGHcvtq+NDbcH
sVBtBdzFAGZSg4/mvefjG5LySI0shUGKS1EbNpAfA+zr+piHt+RcDocVEfqhN7XGyrkFwP1JKv3k
YD2J9rrtXZujI+zfymIFv4M0+KxZ6MJoabn5CB40kuGLYBIvqIZ8YsPOSb3c5AK/Nhg29Gf5qVf7
swX5/6JZ33En1abUA8ZR1pux5tjcb1z/cSgqZx8yc10Wm0Dke9RFT7yd5ncO3IvaQdIlHew5bHF1
ZW3MDQEF/DDgHAipGG8b4j1uVi80zygEFCZI/cj+a6VM3PsD55wiwdVo0VbZIOXWWc+Hqv9c2hj9
zRf0KaTtoI7BnnTtDt5TaWbUYSAeNEYLA7F9lgImMGaE7I22ufYh+1wH3W8PAgWMPw5xjWHDm+6K
8HV6zrnE/wYjeUqmmSl1+pCQsOqsLzIvtymo/hqKSa1r8cwYdCQITrlc/Tzbigo75ufhzLeHIngm
qkhZe5xKEVedDuUOtOfRz++bAeIhVEDrJvEKYw6jmvuQdz/Bj7z87WGTFR0aGRtHfahASCmPHwTP
FKEdLAJpeJc+HW9NtH8+hTj2kOnLbc/590BZR9X0bhyPQsA6OCay1uTmmivahVRzNcZ/KeYPF9o5
TncnbI1+5ShokAwyFcPNQ+hDi+MnAjz3iS128Uc1YVPBZ9v4fL0Dd6wE5z31voIbzMGg7CCuQjt2
pgTXAWVvzW4vYOOD9daSZE1ReKq6EzVpYxOL748wPa02b5KKExqQI3xkGXNRDzybhJOorXTGV8zl
/BzSet3846ENnbHu6NO5kXu5df4FhCxspLGyVItWWGHFnKA3MJUgQ1MhF78ms1PIoCNYMN3U/vdl
Ws2BVY4m6C4I77zqnNKBjHOeZWMvKCslmGXOJlKYkKk9q5apUbBzt+WZBBGDJYmNnxHeSCVkz94h
oEdzFT9Q06p0zyUmP7CNMt0itEDU4Jqtcf6DjoC39fqNQTXQ8TwEL/3YpMoyubeqhyT882/gWoFl
vVdCdC1J8oa4pVSdCj4HEHjw7LeNHnS0KwSD3c2FTkm2NuEjNWwqCxXqbHWy3x39QJiyTa5fT8BC
4KR1cxT5suL33fidy3OT0COXqKNi6+rgbZ58QiQG0uHNpIMCGCLokMfclYJMx0Cpc7KMHwkBQWC5
OxWkAssxw02bs3Hb6NFEnW8r2i5Zs883eZRhsLXAyZStGvYeYl167/LL5N3McTm5XaLrPaBifblw
KvxOOne6ab7nUEOiwNOipjrl1ypdW03P1y/TjTx0zvvIyj9z8Tn3sT5MtB3Vmd2gRjF06YKsOGfI
HpRpnYEAwT2ytwRH+4q6+SIxQrWfl5XLRTtQKFu+UGkXtfM/ld/D0v3xkmjyX38oB5Elq09y3TN+
3AkU/RSC+B7J+yh/nrOJPEOVqbyx/z5KEEqX4oPHSAuWm62sL9BCFC8VLJww4CiXBhKCXppgzPDh
4TgM+mnbY1+H423JFT1kFQp65DzKPk8+YJ9VBiLPHM7Nt2YjlsxWmtAe6ZcOe4PITNORqVO9u6/z
XZC9J5pVincm+2qUouC5HGOPGu8OfSVEeD4JHXrl1lrU3Tw0jlMSMhdNLu65sdzRvSIYtYnbGiE+
3kL2mkgMf7YJFthyCiIilDGtXbym7yhYQWRE/uttLRpMdOBtHrNhOLUJ9lhMPjMbsmtuHvdXvZUY
hxDyslqoXkyc29/m1id3DwczhUs3r3ma1Nplbl5v835R2aHsaDo0S8c39pdgkba2lO4uYagrzpu3
ACR55CozkxedX5cn/eiM5QS0u9+1ymc+MfleOqRInoSxH/uYLxYd2L1+rMrO+POSHcBK9yex5dGv
8uaiOCYtUJrRB8leVs/w+oUFgnuuGjJgxXqEy4F6CSp+0LbH7xBfZur3+mz76MdrECgcbXR8VDGl
cL2UW0X6CpVbjfAOY2pFEAS5fSG42zf0Z/0uWDgFPYv3DaAYerDa92Z3TEPe1DikJcjuhpb3jojq
GJ4asym+Lu6YBqzy0GNTmvTuCN5eW917OyNqaW0wKCNRMGxMWwAyV7UtXp5J2i+YSxOPzOW27QGa
hfA8ThlHn3Tmg1ALdj1ADM6x1qEGR9+GgDPhmhOR194Uv7Ypobg8RockuXG6MrxeTuz+uuaL6Wbd
WncTeqyJrghBU8vFCoXV2vAFrofiF+qGyYX18RUhYGsRp2s6/SVUoq5CWBkudosiMOfGbEejUFze
ZZbigPz/szncUXWNBXDRyjlh43p8IYbj7N2LDvyYjRo7xGDiY13E/Xxs1wY9vfA01lfAL06g7mL7
Rxj2Acdbas4UMAx631QfT+g22cLyiaWR8H9lLFhXfA8Sip8w72ZVQP+xyk9CV8MwiLsYY0jnO5Ot
RLx6Hbrv0GzHE1fHIexvYpadLsGKwHkkjJsNnk9SROKc1Er8EMI0J4I/NFuAiTQkJAGUBotaQCwn
Te9lB3Z4OXu3+lMB12codpBQlH6GOAOHX9OqqjT5FNrLGQkOWyUa3JaWiwuynbQ3BbfiIRFAhy5T
4hc0J8EUoqf1zjDriPBumd4yHHw4uE+mzTx/Q6Nyy/ge872czRpxXIEG5Rv9THEd5M8bdDVtzQ7g
iR/deLltq2ZprtG9Sh+/iLlWnNFJd2DkNNVF1DLZPomBVDYftR1yS9dcsYWrgIdahacyuACBVCOH
GGwq04oKgbEoeYeLdD+uJW9WSZUWFEl4cPhNW/nerlx/819YAvm6/kNI+Jp0YXi3Hf9uX90vgLTD
eB/j/Qy9UJKuvauPoVWZLbZTBYQnxc7lhCAQtwBZsuZBBIlWh+MzrtVBxxl3CFF+vDqeVhavla4C
ab0eMTNt08RGHUwAT2FaaPZPk8G8MtykovOS2devLc4uLC07SZhhTqwFpwpjn6L5drTxj0bwO0yM
qFWAwkkHMwqiosRWzYZNoRpf1d6kBXdK8pxT/Kg4Hrzp1+i+yeUnbulPPJKidDZSz2KvKnLuVXHv
udEJfPWbT8O7gqonjpSeXv6Xtwc5goRGi00r9XnWrgEWqIvA/8Udo3mGFonjXlNFtrvxGc9RLhMA
LmTdqjfgCWsWYa/Vfo+ebvZRrgtHTIsnpVmFIr5JOI8LAka8x9wHMQzg2AgrwR63I3a54tct184G
ZgCM/XrCpjiTvDoTDwBY3LEn211Ouyh7+/ylEBoagFJLveM4shE4XesuUJG7ucNaSo6N8P4h8YSg
Yf+OPn30VU4JJgbwijh4xlgdpVOOlBd1+FrZEHP/6RgAwaFXICRpJGFp2dSI2NbFaCoGta9gFncc
JcxEI0GEkZQopFPpYmN3uwx75PP8Nt2CD1ayGRlrF/FJKUzcL530VirKwLxMLxBGb+R1JWoqsUbP
phfkecvygCuJBvmGwvs27509289/LoVoYvJoMH9zEbCYsiwDHxlAqBsJJn/voPC0XfXrBcNyHHJP
wQOX6ar/qGUJ4G56b15TpJyYcOuaRFg3TDOD8dpGgSKzlHLS9TT1y1VVvogEzEc5w68490rfmeDq
St/MXVSUWNIUNtc5iEfshMI/WyRJs4wbgz0v2W51vWxMxwcpE8UksP56YH4IQKCYkuhO67BvHMto
1x2vfHGlQd8V3Gpn+w3pCQSn5klKTXzCtbjmkjRwyHT1gAO/Nii5AY1ZZFvCEXG/z8YGS7HFWMFk
xG4JtGZUUBmF8kqr+pzmWFL9hQijq63DLrD0oqjSAndB9xYPbLYGxszxyZ6hilS4vQxxUn3QCsNe
kVnuSQ0Qx6WS/6EiLp7toKgaTOFEayu8HVzjGeNAK1JvTMByVZ0jBq4JcBlrOLPx+iCxoGHNCCBL
eCOMjPB8W5iODfe0NkYLv4JL8L4/JeXFnX/h8v6qOzdQ+iu7EefAt4h073/HoXmom7uDrEIWGMaR
NIoI4EyIFWxmeU1e3ceJGSGoOHmTnRwpGE5Zoq00wUrKP07mkhaZcjHxSfFyHvLwaNoF2y8K0gH3
GQy0VQVwnZ2K3FVGgmm3N7LEl271cjwergXRq/+d+m526VGnSZVUvNfRvL4dsORH8dOCKYMDab2Q
AGyL8NiZFKM7l8RvvuskXfxlxanOnd51RIxp74Rz8C4Qb/3b1rUM+PCeTPhzcIj43pHOJL39FVTV
diRqIPstLQolOjZdSjpB6hg9WeUQQ8NaxBB/DiibM5yP/FgOWkWhk4zwv2bUrRmAlev1DZAJUwiV
/HGHQPdd0xXPYOyFP/wi3cD+UP1tj2FiPv9xO1jHcBLWRy1gvGwwrn3cbBzHRuDaTyTNtbOzP+hf
wBf0R5BuzWB/NpKSGJNpEEKHZovuf0ixTkmVw7mtWvZ+6JbJ9fObNzVkfThFtew/FROY91r/qRtm
Khpo/qJa7XCqQPyIkhEWdCN+4PJOd9RLvoaAKPn309XTISSgI2uSECHl0/o/uF9DMoNM0ofGViwW
lR+eoWF5ow1yWPyj+mGSe0MOXtI0SW7HJklc4ZqOjU0KhZuhNzOSSDkokCTDdXa2Ypb02nynKimG
eV7A3TVblGuQ8sB+FtPMwvjTZMub41vH8Si/5x5NrJuO0Q7vxoAoo4SSN8uGmGIumOsRSJr7Osbv
mhH9CQsXVOsNhZI3IZQ6UHAGO+dozAEuGZJS4qlv+HBS8+XAd5lq3LCapEx2Z4PHrAp8zBr9NY9x
upuLRjwNJlAqwnYB7Mvw0BU+pJoV/p8eYg3m5FX5dWR19QozZwe2cxcZcFDsmyF6gXX5dN9OT7U4
EF9LDn9EL05C8gMGk3AhUWd6lWjo9Sc+32VzVXZWXGscZ5podhNYsOXufY0P/p1YEy0Jul/+EGSO
EEABi1090Dr+fsjTYX4JF9Y9yqbpTcWPMsASM+ds09TbdfyI9OpBbnEPN/Ke7e/u0VAbb+mbNX5Y
1uw/EFCvTbODZ4uGoFpo7JgA+PHcPM46YGE1eXuyUNmcHH3Sb2Ix7X9l5TGDRaQBWBBQAih0iogq
q3BRKNu/wCzEHjbsCXVFvuGLLzVxi8Uhp8lQyODggxLYDc6XdyGN1+ATL9VXWxInCbPjWkMmO9vg
36MaNOxiNCnUBdkxhjvlrEOfsJCkry5owXbGxIFfIjgF08Wyxvd5ABMxHtwjdIjHfTswrJ6XczTp
Ghr1ZTjz+qiUV7blGCvqYNNbBNWt3bxheU/bMKTVONkXYP/kFveBoirrPBAy5a2qZGjlY2oeoeKC
o213shUv+ZpGjt5aiQoX8+yYRZ7OKNyjncaWS8wfDUQmLmfSvPH8xfc4rvz02r+fS56RS6IjL3fk
q4VWAhLSElbUAiBBPxfU6Fggh1WA2m+It9NIdHk6qoo77t0EA8E5HmMbOKMC8M0yRiP6pZXLF0lH
dXGMRiXpro9mL3PLJLnG3VsSpmk4sRSSsL8h9ADYgNzOLq8r/bJ1CG31FRma82cynbA5hJeHNKHF
5dJwYHTpVSD72lB4gLCZsuw8xGySbhWh8LA202cwMHE8gFQUehEirzseaSaMB5955EagUaKk6KLB
O+lYfcnbFh81qm51DY1jlfG4lMJvoj/S6MELb224+JK49lknpJr9PX+M+nTdZTGIPWfE7tSi3Z2w
WcfNTkldwdMn+s+YYAqUZhWRzusLqe6nq/qUmkalcnDl2jv3M7YHdiCVtotWkdyoPrXxr5FA5BzH
pN+6VPUwIXBNeA2Q5cRnmIphEDN835hUOdgTPYADedYk7albJgDs/bhCF18MfjOg/9M1hDqw3Ect
RrVyZqL6gJoaYEWdARKUpeql8r/TvEcLRex9n8izAF8OebcMBqBip7RSgf7uUZpWpCaQYE/dd0Xd
NIZttIm8JhGs5Uf2c/N8f0I2LeGPoEZUUTF4WjtItnKZ7XIRDBrAeNKOLKQ5ennl4O8z/ypf67kX
+wr6EdjKmKc2pa/wW0Dum+ZhLXX4oQN/FEyyD0LeBjiQFCrSTTiTWmq90RuURf66OjnvaxmwudqQ
+1rLfPI5Nw4ahVqQYjk+NNPN42KWra5FPxNQK892yKb2tplXx2UjyA083qLpZ14JOr9MjeIifm5E
4Js5OTJBecmvzfxZS/WCBKQkIKyywtHA88HjAsdjqKUbvUus1KN1CqUQpxDKfDOjOX5y/vHg1fzi
ClQRvOxeG/tZNlqPHB1iCExUt1e2febdoGzueFTgrUPVcRQrTDzvGHucgP5m5udXF0VOgG7hoohh
qwUAmj6OXNAvk0WJyCdmwxzFtfjkkOv6EHc6egCcZgLRXMaEe4+WQ7QLKvwM8ZtOPnwTw9jC+J9m
p+RVq9RlbI91MrRbQ3QD9uHlmVBeVqb2v7T1TsW+eSKpoG5Tv9FsAQcdy/GQyz+pAO10s2FSdnVO
sKGpcyATJG5ODN+V4DhGlh5NSp9FzmJKuw2BYO+OENb+iLBfCXIk0PqmWmoybciFBR3tOxAzfs1O
8vZ+4FfvYRxSD5ouSgGfrszTkIKa4L9o2/hlOLZOmjvofSMrFBYAHkcGrt/p3bndMCPZY8gYdo96
hiYfRIirE8QDukysBRmmbdHIOW+5QRPy1rznbHofpwWIzrodxmYraRqoY193NC4OtXhJQhdTsnSu
S9ekzC/7DgIyR6SPrXPSwCV5wt7CIFZtxKttFt0Hen4S1y8VMfWYd6gWv0sazpjbF/95h/BCXvb0
NKv/Py+Ycc+15OK6nBs7tp2QsqyHUpdO8zJkIqniqClreIm9yOFA+qsP2TLNM8j7LNMD12NenwlZ
87yXzXIY2WBmcsZMUkdQIeWbTu9wRsi0z0e0fsrOsrZ1dASGPImM9JjXQgCTNeVvDITNZx45921t
sEilSZdw9j16HTueoaKCEwCe+EJz/re7ZxsjlW/acqunBiFeMfyvZpzxCkqEMK5ukF0OQw1gRJMo
xkLX94lzd/duc37pIC8QRHgy9vTajLqkgUbkd0LR3EC0PV5X6oZSzGd6xZ/Cqe7jQKFhXr+4vuu4
FDWAwVe44kp1wtxJTHZbEqhwwtdDMGvgpUjiFzKAsOZjRBZtz7FbPYIUg9EIo6bAb6GCroXb53Bn
XcGJW6Tkfc1YjQMTvrbd5J4jzAGnbHTJF14drrvUf4qp+fPvn+b+Z2i68LfrJl/KDtmB2iIXoVK8
4M/B3jsUi59e0vEcnJkPU5aF6uF9VKbG75ZrUbqr3EdeZ/cY9UEfny9mldNSyJ1GOtWA/ZAzQrxX
cTa7Jawb60umba9PVTif1vwFZss3at6KHFvHrUgxxG7jjTsQYkJ0nO37W5siDD0nK5esHdAmUeXK
QtJWxqdzYIuLSKAG4IRCdu6olRzhuVo7J5NqjlRWK8ePpoluOOf5VmBVnJxTroC3yHS8w195YxQd
h6XfHnl97xiqCyzUbX9mkLbjrQRo+CoVwI8aS2wyDLyj6hrY9CznsaJ6vCNW5oEWL9j6WIfxxdGQ
Do1bLJ/rnDSEkLPtb1vhmPx6Tk50Jx0sLLBDNnEguqdd1QR3IQNj3p+6F4VbnOV+VhZAjpvMjJev
1YE/NZbWv7Q9Cl79xBKaLVVssP1jNKOsnVd28ldQkMyUGOg1pJma/nsvJoLgrn+Eh6N4p/Y0PU4c
8Mam4cAKuvkOYGfNGymyC+29Bbx75FuDu57T1q6jlI+e4sO4+nQ3Paz7FOtEC0Bpg2B1AdKBz8Vp
FeFK4hcU2jX95mnRAfJ8drz+oP7B29ldNtVIKjEBwfsDXBAigYnsBUIluwI/OaxBVX35hR0jBrBa
g64ICLrNkDNdY1NWJ8zZMdrQ+wK6UOoR5W1GY7kYRYkRp9s9m5O2iTXgUgA/+PZ9MKFwbBfTxrpF
ybI4cdUa//HFv0fCy0GuSAXnZUT44H1ahyrx1NBjziHgPWpoxL2V1R3NpwuzPKYS02XpdhbaFGST
8uQvc0iuAtHeMvAniqDwQrkBvzC2xxXyLwMOlFJRlLODk+1u3zGNAnK3wQ/4mGGnAxf9aOp8rDJ9
PgSxa0nJ8W8ystESPEW7lwZecNFUgkJgE7kK8AWmI0y+ofueo1qPpBOSBun2Ph1R3aaO+zmdy4+t
vMav7qLD+ALea2qlNJeO2o0tscLbEPJZR+9cKSxvhbqwtN9PQ5M3w9T9Ot2YreQkD1+4EIix4pJ7
D+pJ7A+iZcelE+ukAs57599E9TXb8dTlSEMG91oDLB4apURVbsSbFS+STmbcI7qtnrV0xNcmJyvD
Nu1cGl+FgwpzSdGHI6IAzFySuzlLSJk+HoZn4/v2Jbr/IMBT7l5gTT3Zh0QqUX2RjnkYczJZki9l
mOKH///3nnY4FZOtKEsbCY/5wtxA7uxj8UN43tnektDiciE+yxerOQNszrmQowOGN5W3V1zOXUkj
EXl1QXLbrnOmiv1V3r8w1OxDWoTLqRy4CnFanOTvppobpvvGfBE3FmfdvDIYq5OsCAhBdF3knRYi
UCuEQeLTc5OtJ32Qs4dsDOYoHmiZf+wbbULX3l8+zy1NeoDZ4uQpVRXhJxoFQKkaUr02Bh6vsD/Q
9Nryrlp0enTxAN/5AIsu6z31DcMYEB/C4BjWYfEmHLDaQwHF3lzhlK/ZV5z0NsIUrQhYscSUHn9w
kE2dWQ4s2QpuvQkTaOXt+lugg7c7WMVBuOW2iBciHi6JWUjm9fWGHs3ogXmFvDoj1GH5a+0SrV5F
K7WK39b3aG2aw+ZfzDS3NpDyNRbCFlV/LXMF9LSEnhRRMHG+KrcYr8yBhmhnW0rEjPocAeJgzKbo
CpK0cu2TQS2+I4Nv+lvA6mJNkJMj6mHuk4xlhTeGmenTmErTn6AWc1pKOK2mGeSgMZQzSVXNondJ
N12WcTIjTC+SkmVxhbo+XbVlNtTdjKsZYcDVfmDNgyptJmpasyo2dUM2PixbOPl0G1pR5cU8RZar
4MMAC0oexAFTl6GaABvPOk3H3nkwMINNXIFg0uNIA4w+AZqL5u+BY0U9jPVpstlZlkKPdAql0wf2
KL/j6gTSoczD2KwSt6/gtORB6NtxKku6C19zWm1jRytWxA0oyHN48LGg49WI9eYHU3QTTOedg+C+
cpau1Z8KTpbyPnVq/blCMw5qtJlDu9vXrml0AAfNhJxQJIpTGVAC0fMP+4AfpSuOwKDh+THHwaby
MTab0zCEtN5tieJgJsWlbFPhSZf5vFtuYaO4DZmCPcgH87HFQX2iXZxaVAvtOuQ8AkTPVD7tsroe
eMMEK9x0Rd+rqPt6LGWP95MfQ3mNv+UI+6BF/ba79f4QEDrCyfGjHs0JmFpdKU5QSog8MEI9gie3
qqzx/ZISneyi1oQlOnINQCY2HTrw9yknRRiGG7zCkjHqjBIOkwN/FCqmxkIND2qPKx3ydmdHSWAO
RfGLcW5+t0+G7QGG2Wc5gPhG1mYmJrWuAcOf+P3mjd4M91qaw+0pNRLOc9VQ599taytwGIu3R1oE
bln0famdC08LZ++4XWBqZMBjZDAklKFKOrXF0Luza1/xY3TZcwTlbykjyfxMKOEXBE9T4DXlH0yX
cXQt5oNIEjrBYvNwsretYnXYVckapZweN6aM2EXFHZs408rA54SSgTIB63sb2+GTvtgcDVBgvoGf
Sn/pnOFHVzLeWoIWQL93NNHB2+bGkeUNLJGaLjAAKZ4eG59bcG1mUyclUR1NqcbwmrekdGfs72t3
7W9NrHJ4tdhW1WoCm407vl4W0LxLKYiqFiSmcXlKIcmcvg/BY8aljjhoi7Y6Sc4WkEo/M+qmhYLW
OUwZzBNTZzFUWmkLYFNIy9RhkUi5EgXuhEXljF8vDU8i2xcmQOsMM7K64uqXqsnBfu8PVgghSC70
OIo/6Qbe3QsD78fo/FZ1Tyx78Xgw71t7DTe98d1K+8qeDIgLwNEc5w9aWe3OgtaFtGwX6a0wk/CR
viGBYfkSOKIV+AuMyJvl1UY8M+tmJsh7s1FPJwEvxxZENk3G5xpM4+1WQQ/Nw8i13sbOJjLoW6gU
6rF862TLXnX4y9HKXqlMDRotgIpwiaVNLc3YhJnRYLhWF0Q4GrKty3IAn1VUF+oAleEWkfFT1W+Y
OzXRIKI8RVwORVaOGX58vfht68e32X18ElqAGKnvFDFBRotdF+yYlKyAsipHJ4mo84lrM6722sR4
/SAYR/IKZMUing3m5npkvYNLDVms9nohcPWdWGKsJJ8Q8aesAC7RZER0UZiODK1RS6b7fB3bYPB7
GxVkQxfqGvLDg46iB42GIeqgsmP6prDSgM9bRrBlE2QG7qSqXbO8YdZ+K8WyRQyF4TMli/LH7yQp
YwgUzMDYUoYBhV+cMcGm+Ln6XMpHk2I005+LbAU6Que8ywiiOOm6OQV9IeOa8ualDxkubA1NAFga
ea0XHJtNxEqUXSBYFkAnKk28ZmxBYgAGvI3h8uA9KallhuVySiIp2bNxnW0FSwtea3pneSorT6k7
n55qLOBFYGZemvrmf27rMcAW/j0HXzOnTpr7yfUIGpwkNT99uFPVCT2h/6kFM88d6GrrtiVF9ztS
iTgdG5mpJR0sgdADuK955sM5uWEKZb4p8VUmnUiJb+DF+k8gDTCBnoSbqahnmJYzs6GNqTlQ8Hmu
8iJJPQwOhyU2fWJdg+IOY4PkHRihX/ze7bMmQ8gP/xyuhOgOFRZF4ov8oYfhGqeEmNVLP7Y0DLuc
/oG0zmYPLb/uaPVM8BO4/6MrtVIoyyj39EdtwG0CKdko7CEDyC9TUfImFdt/z80DEHZSMAwV5GV1
F9JcRGUiH/2QmygE8neZriGpEKjCWfFn1HCGMYeN5HpjuTFr4nXaLJAJj5FxenZRyVSIPz2CEKN4
Wt9znx14E6dAy0eV5ft3Cr3n8fIgCsybLSnEjPbQCBAqS55VbQyIBLDqkHe44dPQeamALc/KrH/H
AUEymb3FtxZc/Y14r3F72GEOqbJJGkouFzqZWQJE7ZrRlTZuAuqc5ds9x/eFbCfg1EhbSI79DKTo
khX9mW5vPvTH7CPeFgTWaxl5fPDGa4wT+nlI72A6BS8xUR1udikxqPJEm/ISM68k7qvyrHdDQ8Qz
Dq720WT1hkv6fN6Q8crHcNYsJd6ijet31kJOyxfHf1/gw3CLgzN48PhCPZI9Rivlze+34YbSfLUq
bI0KHkTRnVW2U2Z4mmpu0pSiOGKiD1hNu76hOlnELhJ83cBQWRd6kHcUnVPkBkrU/q/9jj8oa3h4
JqsxDtVTF1BZcZcw6raWb6dPWxFdP372YVoAG0nQp0j36xA55AeNPF3ODM2MWm7DVQJ7WqF71veC
rMEVFh+115ZuRFjHBKndthc4foi78vJYTiuqdTDqSz3I5W1rmVRk491Vk+WKVB7BwogFnM35bLIJ
J/SEvCuSlaMRR7eI1fs3F16s4h/Jlh7cs5QIK6v4bmdNpNNWUiHEWJZl/KlKqvTIva65gvXpCvBy
jt3BVORt2PKo9KH7wZ9Vk2TrxSJMnsWuLJ8A5GONemkm0nrFghA5/bRc/gUKuxi4ua1Y97n9gNHr
hIVRnZVPbZMD/fg3Z2InQ1buUmjTLUW3UyFctrXswFOjtPQvj7EOYYIO3pJtJbByYGLMPVszzTgw
YJomCyYBJL4PdAsrtFg4gHV5SFe+hJPpqQZvF7Ev+oeQGGtKroWtiKfpRJoPtLJg/rW87QGCvqCl
USQBxhy+gweG5XNTtsNWJ/Ub90kvnKoY9ujUhx3i7gZu/YOQWq+Fl1zYKvURw4uRYZaAmP0bjSE2
2ysidTwKOk3+VftbqMxJdhk4XrEhuWoYu+isq+VWNpNx/DRaQ6oEAl62VuSQpZbTnYbd4zQqZATA
iR5Ny2k4STJjAhbIt9i+oBL7LYuji8qe4T+2wJo9RzHaXlRl435+RHhBU0kBagMfiu+9M6RHyNCq
h7c6RmeMhsmpA2r+unr8ovc8bB4YHBC4aaNFB8ROXTRi1HZuraJ8P7PY0f7lITpD734YOFfj5oeW
KnwikIZ0r0xNzZ4gRn4K2/BIpDaVuAEKPB9AiuPGEjF3hsB0BGfQPbEgwIEl/hs9PBSBGjoTRJsw
XBj9cltJaY3lXt196BrEb4krf+BaxuXqp+BtEQFOpDwUUP/9e4f2AfbGf8PYypCZMAiFKHIPhs+s
FHlBQZQMPVBhqap9BjTnToSiPsK9Kb/7sRc8hwEigBZdtC/GIMw5hYP3yA04CVpVnakekdjlOWY5
EtE+cBiidqbKNAsSOQjFQVsUCoMfhXKvKatS4ENXoY3CwciaDmfUQNQfauF6TGrlW5qS4Gus2FAv
5xxNwJ6SzDMV7XEUq17xTTpeCJWC4RL6ZT3uJ4z1DvtKAqAxdoPaIAMeNkIEzhHdGMKPhUEdAFx+
yLshdfJnPdZTLzMEIg+JIpHqvxQ/27ChAiKM+HG+RpfaBTCd9kfQ9WBoQyEWwAnmOpGTINURQIOl
CcYfmrYsSbsy4rCqFipCd6DQLyALkNTpOHyDJEFCHggt0PL/uDoaN8UU+UJb6+Ffu3T1TRjqTlC0
eBqCPIHts/WQnLWF1pQnckdWUk6y0HU+pn/4VYlDWK/1osKmnNG5CTNVdzb5WgskOPSzbgQnRRLs
gu0fPoWPAj7vheuLiQ2hKhP1cvJP9Evi04omoTnjgDKmIY1pjy+koYlhJ5lTnv9QMx7ogUp1SguN
05ul1qMAB0PKnlz7BRTURvw4yul1dXu0IJVbfP/3BnvCHBk81MEvv7brxBScaWfXbGPKq5InS0qT
4sClBPpP3NMSoT0u6CvVs9RgWlPKS7F2I1eNxpmgjwLPmdr8ZFu8tdaMiS0uwb4SUfuHhs0iM6to
m20VhlBfI0gy5OkFcsfMKO7HDdWU2vHbJOm83oe3424qYlEs8Czzq+gGZ57gsbHR6STrgkzKStCH
rwLItw+9h14/2Ylh6jSKVdWJ7QcShsHQAhf2I3GCfSt1zf4xOHbIuKMAIkiEEkMODd2Oa81lCIfe
q8aS7zpiTKIgJSZduNRnsPy5UvGSDcgXPPKQle0MPONKjXbASAKe/G4ygbYiBCl1q1urAUAfpGKZ
ZBg+zimkLOJTJZ+P411pARnNXJUneYZL3fs+oSZaV+D3qZjS72tpYxwQuirXApIkFzuxPxkiknqN
Q/JjKdiTCjxiam86IN2/Lws5k/OcpJUEmf8Th0dVrc0BKfHJkfeglSqOrYwPlwkNiCSHwpSVyNOa
WucSDKhw6I0PVH+2KjR+BKBazSDvSiT+tkGZ1G+4a+0rTvdY6/BcHwHBqj8HGo5hhjY8uuETZtR7
ByScDJ4Q+6DmnQ7yD16zt+YkCN+ZbOls8I1qwmAJUj6WlFdCMreZsrTLmRkHRvi8PJCNKdf1SrZX
v8TWso+fk8Sy37ngnyxjP065uwOJRmkoKBLrsf4zaOkA45dScKEiTyQTbzy+PoYCUqw+A6ZB0b2V
uVRnWUw3o9aTgNfBTW+j0wWUQ1riiVdbDAY3zz9+Paxn2jtrDJhQcYYIYqc8eUJD1dLgBYW8UB2j
WwwoD8WVZjpTcPFrRKE22r9bA173272Q+NCBEctab3NAbaVtmkNxs0sw6MD2Ug6mxvav05uLFJRb
xq0kIZgLCnzLTINrrCQNR9PREu2kEeMNm+oMCGrJ4jvlHgAFAwCHCz+DibUp6Hzigxh7AdADYai2
Xk2QQseZJ2WoPmPrJOi0OPbha2QsZIQctMdoXiQJ2IdttkgL4cp90HW9sS/FiZMoIMPnR/WOCOyL
B/+bcfX/A9oFQy/k5+ZHkFfZ7tqj3iv46/tCmsi8EuftTZ1kmwSs5yiNhCUj4HoXk1tjvMhC7b9/
63uhQYrEau6FJ0myQgqJpddmSXoIi3cT+9uO/D3l8iBTFwiTvZdyOrO1wYllSr4jaBKMackHgiIB
lk9ktkVFVvCD2QFCwcvqOFyiec2r7YIUCJlHHgjlmqMK31ys28XWewhtlYeG+57GLUt4JhdSTqIx
503RcsXTGHCdw9Pu+GpKe6DwIo94Cz35oGuDifMhSV4pePrndmC8ISoc/rJHZisD3eXQZTy0QgSA
ow+HFN/BBq2v3FIqMkukbT9hBW/6FaG9QbgYc1nAIGys9hhu8P6iOpdfFqOltiV09jilkQan+0fN
f/SmXoeSHPWobKpkoC9Ji/Y4ERfSj/D5UsAhT5qg5ZMCmTJwOxXmZKh69qFS/bCVjuvMEib4ywS0
O0v+ZuHO/igzJYi3/VY/eiI2oa4fPu6GljY4lahw3vgZPqyiA6FqskWHB8ZiUNrZddGkliT0iUiR
Wc21IFVhuyZiqCriJ8JFCllO40dPqoCa0P84yoFc7azoVbjyzA4tBna0oqZP8uMy9NFgE9Ae3ucU
j3wqoWNBjOXMxzLTXwhE6xZATiFLpBYuS1hdUmS7g6XkCpFQ8Vg+X0KhBpFCFwZnAwKJABKozn0M
0BaUSNie/KbBHO6qCi363kMIX0h4KJ09r/nRROh0M87H5hID5u0NW0mRY8h+IFju+Dzd10cHNK/V
/N+N/hZDzYJ8HXcKDihV+hliD5PAVl51A8NPmZziW8JXbtyApKEigSqaeIWnWgY4RGq0mCh1FmN5
lylTx5HzMLZ5Lxlj3v/zejZh10C/gW+p3vCRSPwppYnMe9y1XBhZ6WSfOnUnOIcDZ+y7T2l73Ish
Bv34anikBsT2dQsy0du8HrTKvibwsf55avg2Kjw4VaBZhpl2iIM59t6JfIkwqKRL3KR/40F89T6o
hC6w4jBCeK1ibEb9mpw6+UXX8gD6EZHE683ccLi3eYVKBfGPCetax6hPnWAzSZTzWwpiG3yBfROj
MN5dR0lfekOmYHXGNkIWNV3iHQa4obv69wNJb99uFRu1E8sFmCkBhntBZeWoiPvcjMaDUsVqoQhf
Nohts+VPlq1bx85w6ZajZYXuKvaxqBDI1b+1zRXgT9jCZp5PcERoFM0cum4Q0k6IsujqmF8I0bA9
M1Xxn1Pb81bC6BdTURW8HGKG01gCcwMLaa7dMJZVmEZXlHR8ZliceaUgSToV2zwSD6wRaoTkW7DY
Tp3gbvpav28dyDmxfssXAexldDQLU7AaoRiK0iutBJn1EyVYnQWgMGBQoewUWSXo5qfw6irNp7xa
APxZsC1X9zl52rhbuxPAjrULZ2PTNIkeBD7BCgLx0fV3e5cJjwcULajiuVxmy8WptF0EyGVDW7w4
rVor+UAXbWJeYodrb5JycfoBrjFwB8etnwMdDNAmWSFytJt1Ka14ZfnzucSfONMvZNVquEEtX6zF
1ipEfL3YT0XXwwGr3Neat3TwADUI4o8t4pFglH8ZzlV2FZKjVHWteLmJh6zSUhlvtddHDGIpzxpJ
/o8ksbbsZrZwO+xi8+xNhVDbl7c9Gu47hZiC5xToKDGB+lP0AIUAOF6gTc9lzFxGan76iVojLaNn
BW7rKWpi+gRMvHGOwQWiTDejHsan0GtKZ5DswiDP/eBVRr3h0KSCwUz6AXNMjpeI5juslIydHWmv
KbehWr36rINcURrY/oBYU1TrMI8ZNxjKZdavKBZRqvnjMvkCJlOZvq+kIkF8b9SIBmBaPqDGJ79/
4ZeuuWnTqdI+Ux2CTvGWFt+0iVYx5tM9JTUR8XSYq4TaH4BI2jM3roZc7tCs43TFnHYvpSS90UFY
QBpf+edWtLhvxG3tzGnba0O9lb/ROjskbEUmrZIgfn6B6f1oLMj2l1RVHpzGkiBPmN8QBwtFxsCc
GGcL/v6BaeamVm9uMDB401VixsI4qOF9b2ixpU0+dB33lSONtcyyP9QQgtIew0884dFxotqfkyhS
yGb3rHhTAPMTguO5dGwFAtFaDm206q0sb5JrIAj9D5NvpM4VBaIBCowfk6X9b/BmP1AEogs5U8RZ
9WY5aA+ffX9d2Cdb4ZnYUdmpcOLOnGiCxhPXaId+8e17S7fdSvmKGHB42r6pYmyC4n9NiJ8O056b
d0lpuIAUoa0ECvbyAAM1x17GXzqGW1go3ogBogztgnoP3unI8P3KO3BEH8dmtbrVcImo1fZ1R5t7
PfZwrocH9Q2WHpn/arrIWk2+sfRqnkJMkZrRClLRBRqeW848Uz3/DEg6f+H0MVbASUegzmO461MA
Lr48R4yUCg4dOFdGvPdbhJPxJ9zq1jEkcYi9Yxy/E3pt+gkJw4reke6zQkUNwK+TmC6qL4D+aXGn
yPmyqtSgUjyQrAP9yRrnfdd6fTr47x7mI/VC3j8LpS4udBEUZD8VHEJN+AsV4LqdP5g5UvV2Yz6U
CKSSGSs7FZoYb0eWjmx9p/PEalsR19ij/pMRVmjfxgk0re7gKnNyxqfA2/UAhBrTTC3gT+lG6RRC
faOq+ar/kewCjDqDmqNyGhGgyk7zwLtCYc7C44fOX6y4GnUcBXa2CvP53pfIQOSrH9X75ZzC6usi
Ao7zARkHq6h8LJqBf4Ad6ysJIrDWT5c5yEZ9CNWJy2ZsWEBwY9bu4jK3YgH0OwrZbmWe0szjYkjX
pd1GOYeGe/lpRAMG8NHd4hZhpIvcNvnrvioSO9nwmKU1d0W1j8Lz0yXBlb+Rj3RLHbbDauWsXBh2
QAj1EoS1/zzk2wRLS0pPvn0XUKV913yXmKf/NplNTNNScYO+2orHynbyYUCbxVa7Nsv4lFv/9//7
/s6Gt36mIFUQrClKFv595/9naHjsoRc1KTH1LImv/Rtksv7hR5oPTQxtIyO9DflZoeTH+Td6P6V+
C+tm5GzkxiLG67J036ZwocuUQUFvy3VHBolRuxabudIxYL2rdJXOtxL0Nqu7eWKZ6DjA7NjYVft5
5ZFlj48B6jsLHon+h0ehzuB4klvRbywIBzH7jitfnIaU/zc6tv9GTRmQAcoOZy8H0fpQsatuNyk4
q+35QId8Jya0Gx+CFO1P/NDx737y90mjHrZ1FSHRrwZpSE92NFRPaKKUXqJkaj40SXNeCj6yPhrU
1uibD6cU4DRXbZiYEnlZvoGxWmhdyaTULr+LKAFXGGz+ONIzEsPsKm77xejcywYbDXwTUGXWTe6/
eBIe2ibOr31vMh5ujy/LnWQ14fLqcmNeHehGqbH8yc+fygTxG0ZQmNyB7YhjAPn60Zh9uMlox/Si
E5eRCl1+ex8p063wYW24dg4MsWQw5a9nVXZeftxV3Dn2K5RqLmVtnU5kATPfoAp9sHX9gObsYoX2
rEVj/NKCPXC+F4mF7UyLwsLYwC+6mAbAqUFemU5uCDFK5RnvuBsMS6qUcGCUEngO6QqiU511o20D
irnlLV3LbxPiyAbVGomJHTAdTn5VJlh/e/D1gUAgaLZw9e6+4ditzhjMpfyV/Ed2Hg656Mnr0SQZ
0uJWNK+KBen3wgSdvS+OM4pCUdJJfMFTH/RU8Dcyj3LuCnJMWo8ZMpc0VnKUCwqR7xc6G1TZRZru
j3Nbb2bDjJPBqX1ZVUVACPpn60atjaIv6ZmZPhwcmHdFOrGoA+3bCq9x3MNE+L1TeUACQWs5GYuE
MpUq+Utm0GsHCeuHo3NRmezTcBO8zLQYVzald00ZaCEg46t1fgslfkGWO5LJsr8xhK9z/Uc43osS
lsqzjQQyDTF18JWT7P97TACVtqzPHMKamWzBkdOfnVBJ07FO4lu9ui3KoWbFIt6/l6QYTwgCvNah
1nNSrK5Q3zNocAqHua1xj0ZV2MaCRER9/CEGcMB04F05RiXoQEH2AU+4nydMO+baILIWj4DxYwip
ontD+MWmsad39Us05Pw+Akiw4xnhOUJYBcXvRIJnTn788WDdRJDjBhxl9pQSfs6LjwdBqaDgEz7m
hO4hSCuX+sSdNxzNGTdHZfEcK+9BmL5q7y7kw2Rokx8FVd9sgSx4flculocI79nlPVp7fSuOGf+Z
O989eo+kSW1J4717nfJpACLcOlNTKoH3VL52Bv/br3tmzzesFCivPTEo/EYCOBdABLjdIOEVZXLF
kdIYbhc1cU/ebQ3Zo24ByPjBwsES5AG9afkHl72PPQEkgkZfSy7FtIn+wF2f6sXVC9yVVPFSMPiC
eUIzYn7lHyxYZsJ4iX5XuNcUd056ifLQGJQEskcFDGomGArd6h6Hw1J73GmPdAlSr7abWGgJiMqG
j7g/HWmUgdYr0Pgh6Bdk0mFzm1HLeKL6uAiPu4+Z7jI+3XFq5q35ECJv1GYA6LuNjOu5hU42uAc5
ZdK0WG7GihKERCOY4dj1eC9e9300/PHR6t2W2vegY8kk9hOI4ndPDtfXQlZyWFI/oOVmOG2o9AH9
5XpScNiN7GVH+BOtjMCofHBYC1pN2kEtYq4dIpS9R3jFgXemU3VfOcbEnZi5AZ50d2LcCuZz6Yzz
qYtn3pHBNUfzRtLgrHFfe4K3oCB0aAMhR9qKSFMSq5WkFOXiWj0FswVelI/t+qSTUa/OcSYVnBi7
J05mPp+fjdS2Ajo+FkqkurQyBuybXi1enW8st0KXylQFwLRmpVYdI/TDohHoYNM4w/InF9KAk4Mf
6GmRX8tsQMx7iuTDWmvt+/6QCfs8lKyQ9lr8CxhYzypuPDzq8KXuiopUXtexjsmvxap35vabubAy
5vuwV0527jkLiGAyudexAC/KdqJM0t5yVQEngXsUZkTrAmxvY6qrbpuC3ugaOh5pRiziD3TcRLtd
KaMQw0H7L8qCb8mwHWYfZJ082EPTVqmBJ15nxeZjUrys/LdrFpVOispybk8CBkXYsQJpySgd4y/S
SYn5cdPZLR1aijK14FoTm4bQL7HMbXzfDLYxyv0BiwHEsqJXXiPZu3pLHP0zg8qJs3Icvvxvj7NL
Z5RoWM5y5wnAv3OP4Ywc+AuUloK+aEfkUPe1rqOWz+5xhB30Qc8UZTgzoZZ+1sFeS8ACnseQw2O8
ZGR7aPZeU6Wgs90ZbrYdQog1iUPQ1k8e7r0uMt2UZS88EgdqIZp+hbCYdAFvG1GneGC7ZnfZ8U2G
WaoWYr7rChuES9CQ3IK40VxYWhBc2GO/hT9paoMo+M1+bTXBH5To27CLGkBBhdZ2yzzJWTRWbYA+
3yHAJOCJF9qt4DKabChwHP+mMO22WPq6lyIH3XwG4rehA7bTKRDL0w+XniOIxaSiTrbh2qcA3rQu
byuNuIPU+cog8t7zPzfpcy6/QAPjTT0z/yzqgl2cRoJirvSWakNwsgZhRQs17EYL5x8D9F8yZpNw
0f7wJZ7zfByilro8/ozXvTc7wgALsPAOZODJKPntNRXCh+52DIB3psCaiRTRmAaeBJEQ5CeJ7flA
LBPPTDgcD374zj0n+tpR9mDY69dIHpm22AGzElKkf4tOruZYf0taJDYhf9rAoJY9vKz3tbHh/Nf+
EwpAMwQ4a5JThSB01jhhpqbHnj4ddDHjMtOaElpWdPkPTLQYDhvrG9sxlfCOL+b/YGot5aRddzJb
DxHriN9BuTKRyp/jorSC26qojYxJdRSEA6Jt5bvenQ09cGY+TJlwXs19TQlUa0tTHsa0l1uPJcaP
T3rDWfxHcQN137v8FBaBxxu9HmByYU0vEw3BNwP3tWvFmi9IJJ38krZcWIGG6s1CsBz83f7Fg25+
a1xErLSrzJyuUuptZu8MSyjjAgd4/4TqxkPyA0L+1uk2y0DzkER3lGYqU4myqKLyDKNifjR9CQod
VvUKFqVJW+fu5hxNfgEB4Cmgo5kc1OJPqt82cp/rWX3F2SK5vMFHZGQqIDpeC1MPj+iUbZj66FtM
3eqvh3nfRAzMGBWs3LBnh93GuGNaM0sxhKYuJKKDt856LuBhedUmUvMKXN/L8Mx/cjO3YIAzkdem
UU057YtkeAwN/Ifro3hXMnnxsIZaDAoAfe0Mb4AWDdfBAuAvADSmEwVz58B3iibg81kx5ccJ71XT
qet8ryN1KvSNDtHmZPmSOHnN+ZzLyZun8ch+jPUWQi/lUIhCWtMXCCpONc6HkkpXVHwjYXvEDChJ
Q8S8SfNMTgMvNZdlC2zLgvOqkB1l3RKhdtM+rr56RPLexD0Wp1EIdXS96J9uTOJJ+MHr0b65aPEH
xqgifm+5gYuk/y3pFgbth49hCy/EJB/AfZvqY2qLdOTqoBcIybKFy4Md0psP9VXIf7+g65MOGnjc
wALJv5jZlkN1YKWSJKfUJ9UoY6jt1Y2OdlsP64oBHGcEoKYzNROO6YJSf1VMEFfLhtlsHZsI2Kiq
i7VHPM5X9l67UYvH2k6ThsTFXTSo0D2g91KqEVYl3WG/Ipe/0cMfqVP44IsafHke+IIHBX+NysxP
YUvHcFYX1mT9edF1IKx/CFOyoJcBidoOHgjsizH1ma+jW3hrKZZ/T8XMdFwPIz8Ej5KzBfQENirY
B+iaofo/PLI3zUoAQSHl5lS4sCJiJzc+YQfSB9my4S5J/PKlb7EO6r5YBghqi/QIbfmbDqJuY+9e
w/H7MbpSzATGy1i++Zf/SK6GNYdsQQATcdZusiNSPQSom/E3BIxDG152RRWmzuqrTv7YVZkNdhRA
2Kgjf0nnj4763XlAZ+EE82VKpZpJa4hUTnVB1/Xtb9xaj3TsBU6z1GdsUNv+kCHOrW5roK1E2xXm
DGNJba/j9tq/e2E3lxcfHJqCk5C8dHN4wepwDcLYDhNJE8aXNyK15oMYvT6RWdyA+ItigbqspR2l
0FNHbCfN9t7DZzF4gYSQWO0ZDX/PM9gmLslVv+SqSqnql4HXyUeCNEnd4BOGo5QtL86iad+km0Uq
dFHRwfO9ITYC9RQPdyBTihIwjX1wmAU5F4VpM+ue9LZZoF9wS+8FdLnw5lCS49IKuy2si0+J3gtL
R0hiN5W8Llx1dMN4MYtnuAg3hhY57FTAuqJRxcyOgYwhEoijDKIdATS5bXFCwT25HPGSFEFVtk42
+3hrJVzhe8CgTlANMc9FHOTcIjjk9UzQoOnQrW3QwMIauf458RThHofGAAabXGyIg/emfp7PTL4C
CbZv4E4pdlpQdz6rUuxMuBf8Y9STNtJZX0l29O5rPli1zCAv5heYXhPKiaBQMAM/SAgL0UpvzcTx
DFIkIpLKkpfgB8mvj+ot1Kf1Ry+gnrrYAbdFkqirkViIoFsTsOjUaujhucLMXZasuKdoB6tFDkYS
E4votaUAUvvNfMgW1L7FFcALGHjXmVPiDmcBEuGypP4y930T9+t2khQ8qM5q3X+IG1mb98EWcFpH
IH+KG/Vjezi9gvHivcVIEfRJZQSe7J4/1Vi2hfU8+rRaahbrMePDqqmHFx6uKnKUOzdjpzeuQODP
qXbWLxY+IZaBK5t+jJSvtxKBs8T9CJ9oiT5+swDN2SgHMPNnpCRzblzP2luepYTdPIgtncMxFdci
30XjHqA1CSDFYn3NuVZ6g/lpOlgcRh3NgBqE2+fBVZVSWYWv/T+dyGBYr45thNSgb+R39qWFSmML
+7Oz/YZ74O2uJGOev0B27QrMTHY+LbURMUR9gOj9ubU5gt5CWVLlPSTLl6AciMFl/cmho73d3cqC
t0ZLpasicC2XgFivyc6sN3YHy53/Z/+330kXRQpKgdXnDMKwVQHVYyVUhK4g/FKekg+snRuosfpQ
8pMKf1mAuQR3/mMMyBTh0NXCS04Sf36V1BQ6KzXPnPPKW4Teh+jgeEpoTqmP4W1S/cCNZ7oeJIRi
2V8tc/DGrMdBuaI4NhJOx1Q6VwWBsGRjYwaG2BUSZwhF1jWIMtLfKsqBe/Ns1obOHVDXL2gGHer/
Uco9FET2t6d4jxaEdJFbI2g1Jno9ux13jKEpl/JMDZnTGdejwbP1i1DyMwehGhI83Ilfp3KdlfVF
ZfxyU7YxhAWdA2f1cUrU4ZFmtdEdb1QXGRoXVtdJTCe/bODkmBwpy9F/33Kh7f+XQQO4RgboaC2y
+cbpDLtdXLUx1mym+EAJ+lokz1G7YWlblvSewfNz3BfAVIEdtZmYviXbRzW+VVHgCeqyInn84kus
uXdC7+6yJX5YcEN0I9JqDiK4w+kKflCLACEVmITI3PKAAubuqjPpDHsZd8329W4Uz7lPF0BT3tuS
2xunN4Shm3+WViRCqAwyjiwkitmaU/lTVj3NHhcckOMQFDwixnhWW66HnGpwJRzPmQvW+0MU/eWe
bg76UVShQiLLLKEU60lhIabCqG5B0gueNpxB9D/jF4zMPIpWlLLeTgbomJyQCf52N8VzPhvCYBoM
8VpwSO2K504WhiZmEKgQvOB/jpNG8df7BbO8vFRs8gQ7mDkVy6oXKol9/9WT47VHP+4j4QJ+vGzN
HyOIomAIF+VGefg6g7SOE3NIfcn3gUFXfc458AE4t9q0j3Pw4Z9w68pVJYT+lZS74sbiEyiQ4W6C
fLGP7wg10ATYN7NUuSNU8U6fI2wLidKPdh7RYIh825yUnx2jWPg+c4e1wQOYHKzDMv66j8FjcU7G
Z8ppgba25DwSsz7W8/O0YnSzbDw72AdyPoYMXSOaz5DsjedDq/D+CGdyeRofnzpaPzkzqrPhN8AO
Rv2aQ4d5qjGcn1VUCxGTGLmXlgS3MG+HSXHIhqQpJdkSShAfdo5QK8U0uZw5qLIQWEWlnjtbmqMV
ySyDqA4wtyeXvnVLwF5nCZH35v0/ttsOPcFW8Y9W9OCzrVA3+eNikbUlaL6jdiJ9UYSXQKFGj9dB
NUdnDNWDqdkiAhDKRjDA+QEbCWW4vx1ceGjR9yVCJ8FgfBqL2Bvq9BRODZSSd7EuTbebMP9jqqBe
2i3ao81CwmzGH8sdOT2JviiaqyXFfrcb4qdz3c8uJuU4fAmHgMeLEHRfjJIYQPrJCnP6Dxhc+hLw
gqf7PRhAEdLwf1ZzRCI2Lg2r/15KPy8eKUHSH6Sn443Btz5l/9E1ZpiiQa6BMpJzeoFpcouBGxtr
2HL7AlLVkUOoBSS3/owzOtEEDKCZMv9XHgbCc3uHhBDyN6aGnLgxo8RWQdy2EWupVkrgCj1l/2el
VGsCVZmm/66AyqWFxTjAybLdOG4+wAO7UQ2wi2bUJ2zRwnHPTNUdDmce6TrgU9zg9azRIWHuAzkS
+spLBBg0P+kLdgntoUxxPvAwSOfK/3cnyeBzBVLozWpY3qrfXPzDelxKIxlcOoWp3SseDm4+wybe
uQ4iwyLVxj5riPUfRsEfzcZef7RK66c/MzDrk0vN8GEhmLFmwgbnE9ghSgDQ43HTqQSrwim+geAU
NHef/ze03VtQCvmeHlmf1cjrylQYXS3/pXMHq3sfatT4xDy1hRAK2Jx8hKSlBXciCyOvXr1d/WVd
VXLoMwlSxEu2pcOHF5WNlVXBtcbtLcj083Oh/n8aIwX2atg5mCQjQzxmWQoxUiYNkZg3PHPIUgd4
3ymPWGIlgPayP3Wb3X1NetPlEmsSJ2YmtJXME2G5mEBGXZX67eZX3/V2fXa5HXlIioOQVb2SlR/j
sl6rgFjP2wN6OdkjlX8qX3eoF4yXpFaZ4OZl4x6jVs01NKN87QAGxL0lhLhynraaBhRSUe8N6Uho
vvnd2cQD1Inbjy0n7bfRZFaXpS/Y0YA7dbEipHWUaOOKBuT5f1kEmAxldQqYeZm4bN9uneHBlrNx
NTg1rCQblgdj/R95dKa4za4HVxF0aM7YesDVr70JR5GGU1MPU7V2r2XapVrFaf93GHYPK+MUASxK
ia7oPRHYvkhZGzjp1HD1DrG1ZPJmPAyGkZrvY6QnMo53NS9yzEZEPTaLylVVmki9lmHuENPZEJ5M
20wW1E4U78TGz3eoM/lSmXtsUT3aR3HOv07EZYolIrt6YePz/lh3d53ZVjstICd7CKi1/2Vh/9zV
OAZ/No66dJMXSdFFKET2d3/CEZZl8TnI+l9MWDM5WrgS3lihh+v3Cd6JUpS+nisn+hQrBGDe252H
xjWUqzdr4k1fDvmxEVlALHkxUOahP1qhaHGampPxLNtvwraxY1Qv70X/QEXx6RqTnFa4pnRyL9Od
OQMUSP8qokX30sFKl+V6ZURCRlXF0rxT2DHvfv9VOgH4wuoxF8n4xNsd2zT29M+cxJnMNLlrebU/
GMwynX6d91KvE+WxnVnWh+Mhdx1wijhGdL85TF04QQ4qnCUoad9lgkPohr9j6ejg9OrSi0ts1zX/
5KCJXkXCGwbL6vzelN3NqZFLxvhwqhnfQxTIjtz2bdYEVsSVk3d2JlggR4jKDlqnKF2lP9FGtPqi
T3spq6kewX/AQoQwXpetgh7LiSu9mly5WFxfV89+iijQSxll1sE7DVQ1dEIS19hGoDQ/cIQ7mHoe
tQWQ9r6XBxdQnX720QmSu4TEkKJRWi/o+KJkjCrVEp/h+64TJ/MwJ1skwOusQbzcyXuc4i5tGT+C
XOo9fdtzftIiuMepN6XVPvkRR/YWFCznTDOTxUbHlbvSzKqzelPxwokCxvS0Ipmle5uv8zyXz4iJ
yRbUiZCnxFY5/jr5SPEDeQDnSFBd329a4+FHjThE4BJOcNmympLefPhys1ZYwyNL0gzbecAvwYv3
JZI1+fLGdkF1e75eQMtSyaitCFkBZhPQJhhM1YdbAlf6cvctnyNCFFbiX2k7sDaDjwbTda0OLWFN
zXhdHcOWoL14jZ423X4HhiRfS458m+qHAMZtxdI1gTR+MM8ZyeVmVnLfTjQnVpIP6vohHEum6k3l
dRqxPV/LQeHv+FjoPbcOTG4oY9+blQHWSjUhcHBIm+CPVPR9+PaKyDbIcDkHapSEN5sawhrNhcGr
UB1TrIFIms/ocQ9sxUBue8uD3tyXjkDiJPKkH68SUNefSLyyzkjPflH/vBHxzWWX+t0l9+4WkDQA
jAw5jixwfvTmwCGnBt1MwYwKdUnkLyEo4RLcbj7C2uGMOkSk9C0CbhZnHpN/y7TymgV5GVIlx5AY
CHD7FbcUcTm8T0HnGk5haAXm+n5uEXF2AAFOSkFqdaJd2IH/js2nPiW71UJynrNorblCx6030Au0
cGmf0q2iGptXrvAxjt0e9Ru/8LLsBpOT78XcA24ZrfcN8SVT+RotVKwL38uQmjo4KNa6Q4pDAH7p
7NlcKOQN78BbYgfYk50Wthgb0ErNVkyrsbf33SHRj0cFj213/kpSaL0Nfrc04x7n0JtOWgcEmNOc
qIhI6gyHxfkEwB37gpgjP9ARr0uze4bQ3JdTCpgyB5dKuC3NZaXd65LPolWfW9e2j54WdvS0diio
uCnU1Snw7lTkY25iPgxWrChoV1MJEkKCdcyiOELDIM33FQh2Dmtk/lAvm4z3XewwjOQ96oPDRhaQ
OVAFBQlz1M8R6LVZsljkyxe8JA8+9Bg1Yx1pGqhIMY4NmGVSG9ba4b5yAWJueq01fQrclS5/hmx2
AcjOEnzHqAxUXwuPDJwVkWRpE/89zmWgeyxERxStI+sHIynLxjiAAnjoMrpclN8YJmAAYyxMy3R7
HTJHzA5D7lyN1QZJ/oUXP6thmCgv1tyEdT8gbDCArRp4pCGZro/4cjVdqrd8ZWKcXP2Ef0K+D5fy
Pj7M9C8VYgi1rwf7NYRLfrVwCUqCMGH+IcCHgi9cK/UoCZOE3o6IIvJIvkYBHy6vblFBoAsKKamx
94JtF5+QC61DsUWQH1HB9abrYBL11kHceHUhCeorb+Swf5jP0+0MxgUyNStG5pdGEvo6wK1eYKrl
gCqvJwTS33xel86nsILkpW4nPb9hPEG9JV9f34z/P5Q9cO5VgqhBIPqf3Iq3F0U7HzToG/qyu8W0
VpEDnWIDDbFzIF6qjpx67JFAW0y0LkdrHo7akjp3ssSIGqNV6rieXbVruT5yc8x2omYFg7mCJMPs
kPpyU79KgCTV4O1xj0iORK99aPsB3teyZCZA1nc+2xvNqppARBAEhqOcmkeEuq6lhu6sGPCS/izV
TVLXcyhu7qu2zigRjqlWB/W1JHUZkk9UFZzsIGDsVctHd5k0TC8Y1wSM0sTUYqOzGohLuhQVH4kz
gQPn/MPlbaPFUSMqDMpqxFWHBNtZUyujnuk826vdSJMhYM/aYvqEppuD8i3regICschqOAg4snz0
UHO2AFEu89vzm8NxBejWLsyS9Y79VYtlR6Y8yQoTyUT4C6gPMouQEkikS9INtLJsOr5TwOkQlNGo
JxsqrcBbSK4bnTBtC6Wsb6u3U5HYI0TZQTND/60bS1YnWZFKN7bFVWXvfNkhTopa2FyFOZhBiJpr
fSK3ruc2323yvZxutNQZrUHxIj/O3A8c2VnsZbS2h+WjCq3elg0e/StK1ayF0VLNo4L/hYgTLB2g
gyi9wk29o/8LSdDlWHcIWeVnnlqPJgEkHRfL72wDeQTiucgGLAkDaRM834Yu5inJkT9ungZ1b+tK
Quzzb70cnGZstwH4fli1jhjFyyL1i7aXC6mbYkyQUn4fmHGQyDRRvaFBgLnlO2c2DLu+RpIfPvq4
CMIILwV/DutfNLS3dhRUqSLTP+rsQJPPmKuHLD9Q7xMOQq7ZJtsoZTn8R8h4cRr9UoRsDghl6QtR
iwhdLgi+MqZrNCWgEB8oOp1BzEYvBn4NduSsTWBIl6exr5Dm22sgqeG03Pyo+fOkMoJAQBfzcifQ
oHlr2eMBzKatilErDMvTQI3PCk2t+UCBtz9jwX+lv6JmVHGyslogvVimJbORo5LmbsIhAJCY/HKo
T+GecHEyuDgU7Sc/Vx0WRU0kpgcviQ8Wb1SbKFUIaXSIfZKl/uf7l+5qUSJ/gOHG/Zi1/SCNjYtf
rl7j+1jhbJKlS4OWGypL9DYmjdqFw8/+5m4ojy8SlhNyWLt+DJQpkAytUz3ApCKj+6XD4VG+0HAr
k1TG0IwdfI5zw6/+tD16ugG9Qcfx6tfYVEqeQ9QXHpVJMlYx0bM16A+m/Tyt9Ye0QjpUM1WFOcoQ
ulnDg07MwmlH/hXohWntVXyCYLbYOwlO5Y/HT8NpAdVmT2OtH02BtwXCOULVdTju7ov+wMm/hgPC
Zd9eFOE16Kc2vXkOuaqjSnvMXnMX0hwdfhOYa3L84VbqcIMk3Voj0uAbz8xcTrtIibVIHuZu6S82
8vTMS+r8xJNOdGy9Std+4/9mhzYbVYGDA/cayKT+fIbUQ1B+bLAMTKCgOi6dP4UXVBTuHGbtpyVE
vu/OeQ/eo7hFCP0JOTUbPQyPrjLC9lKlV73sR1SZ5pnc6iZO2Ts2/10S++5RkZIFwrQ9mUpR+87I
zbMSIg91GUr7p3Ql4vu+1Tx+xlP0y2Y8xA9TzZ7VaEy8zeV4ng6xANni5k7dwkF3RA0HwmxWcOdj
VPpBILDFCxU3qZDJq7MlSq75TorACks3POMFL+WDQ/M1EfDiaAljv4a6t9uX1sRS8JaQ9/kPpR4z
cwSgBXXnke7lx25NG4/CO6MjjE2S3Mdc0+lKXtiL5zbgaOvVHyJuMzO3qUQPizfhF5QpXC4TogT+
FUX3Rzw+jIpOty+Z3DkaoTzOIfzX6ze10Vb+10Ew6i+/1tww9qBN8/eD7Zv8VJHMQV1+2mXg53da
bjWEoTxlFCxjNOMs2qVr1PjWymC8OC7PZzyYIwwNmWgzGu0CeLvi0aUl+pMq09bjgGgoYaTnhTBZ
9XdHy0K12wtw+RPPom86E1tNdHIWX3kuHeLO5OFMc0yBwIbSCTNwZsm0EGABzWmAyLCksJjFkDpW
OAwTPqQMzWNAEudgA71hDRCqa/t9VYFV4O6wWKbEwmIymxz5pAfTROvB2ttViu1dM2vHeoxq/XkP
iaZ4ALdek8Dei/xt6p/FsGuOapwlPv4m+9AmmD5SF3NuIkuI2YQGQtRdRDhJAHdr1aWKisUBGGTD
LyEG0cT4zoUGLMysm/nkyUpFV6QIbw2cGaYJFy0MfwTRtXRPevcMaW5SOewfuD/dxh7wjq3o6mNs
86/mWU68cdZzfCoSbb+BZ4BnBSJb/SwHxKxBuJOkZdokjg/Q9Hvi8amn2pnbsxYHNUBUGhDI0CZW
o+sgJ2CiFKrrLeo/sx8TGKw+31jA3eC0mxXXjTOABHRzLVNRVwQZbLOou2WW2VmtH9HqqGjban2O
5jO0pGFUhn7at+W7PJ5Ohledo9MNNrmXjv7nFSfmmiA7ehmwHBNCJayhgDSPPHJsh7b0ub7wX105
e9/WXb59otXBn5oDHDFZpuW6+L0IBbrjqiXNJRSPO3POHLnQ4p58orSXT9mJSOWv+0q4GsmwijDM
xtYO0pYrtsL8YQ4jYK9eCLVbNOFRaCWrp6XqtH+phVq2RXl3ktRkp6GMrYLq+QdvWKfZJ3C6Oi4g
AGXqZBq8zbyDPl0G8Lw5NpDkhcgPgRJ4SL68sJGHyARRQmtfYgbJ/d+YPC5GcajlN1TOW/MIfubQ
eOvjn9zrGs46BxhjgcFed32JMebLHzyynWb7ynY0popkAgIEiLy8b1IDYvTDcfGaRqVVcDhvEL9I
F1GrcXiljR4K27wZ2B8fKE2kbESA9E+oyHlQcJyinrY3d9dZAygUW41CRLTRE/orkIiplObfDjwy
+Q1dSMaXB2juPZ8INu8Qyc838KPGWag9SkEttGLoUC7DL3W7M/8XIMhEo6L0qPATa+WjK9ZBICGu
ILIzKNP0SXBsHge60PCm+/h7my3IKy4R5OxEAJc4jTl5El+v4Th4WYPD86H9kYlSIIc083W+iJ52
bTSVC0gojJBBvN0iIaHEKGbKt9xbPdgJxaGAExqmwHc8ltq24XnM4Kp/Sqk30LEGDGcs4Ii3ddcs
hrRs12ii8WeajMa1X+HEkh9t/WF16vIKYwr475JRZel07CuHSmgyS/13Ky69v3d6edJuxB8hVkhZ
A+S+GFqDeexmvb54fdxQ9w3QMwNn3C7pfDwin6tIK1atScTn11QQm/GhhfXWIyuyZmSHEFo8mb7T
lyMPm0gPcwd3XqjQH6l1tZQnJrWrCyk0DDrriJpRqeX+mkuzn79dWf/OzKfaPxCToqAQ0fkz43ws
PzXMLD3qrfBT0Njt4x6WSzw3hp/sFT9eHn+yx02gzvvnRGXydrvSODuF2YFOL+ZzAmxv06ANbcI9
a69xUHWl3YeGHDPemMpjd30BVSULLM9v+Z/T0IUpZABO/Mnc9yzNbvQD/ngTascl0skp0PcrnLyO
1WX0PybYxInvxdsKWYnTBSMW1aUNqeibF85nyua5jkqAWWIm6jtVLqo8VtX1lhE7pMBh/AYJec10
um6ftDyf9ru90FaVm08OOcurOukbcGtPcDtku/Yw3RecVeLY2lQEle4sGURWxztSkxSnmjibFXzf
GApgDZEMO0KD6stQKxUlCUelLxho+SNBYrAqWqc5HfZOWO/BJXt3bcuIWJf3V7XVdr6mBA0j9sCe
6TwwVEfSj5SgcJRXiZ+zIBdv9C8yFWfa1n63dUoRLENtXWpOreiq6MaTSn2pvf8B8hu3PEFJcVDx
TQ68qe9QYeaHZLMm/zj/S7wo/G7hrTyBg/NZ6rQfndyxr7wznGYbl3KJK4McZA7vlYuqJjVaVKD+
DzkaPiojEKL2v4of0ul1gGyVa4wxEaul+jxpILqbbDsG84UF4mm/153YU5J04/BCcWYS8oQQFd5T
7BMr+/7vud4CQVLFBI9dftvplyPxWpccFE4ufmHhreFy21YQ6eZVVT1og3jYBB4pFKxACtQc5ec3
gsCPvJiBqbbN2B1p4lHMv95E2vm/1Tvb3RJO1FQix2qHovC3YUv1h9OflVsONPHSDks6YyPe3yp2
sqXP8TgqJDjyL+Oxw2nMNt5fUQRHP5xYd+kMOAmKaY0ad7NNOq5oPufujONP42x0xoacdaZ/jE5+
UTbsyNsnl+hqEUOhK4hlrTjh/63rlqzAkQBlkOdawLxcYrWQWiAQR94EBu94k92lD/i7vBU1qvp1
rE3rpNjOO/PEd4BC4vPqFSjnp0AB4Be0nRV5Kx3LAM3P/7D59NyGX+2SJ7Coji3Yu+nyzduqILxo
vH/u9oqtgz9F15AUtOE5twdOr1qZ9x7qy8G7LG8s+hD0PXWub+aBC+Eok+HHnHZ48qVyH+EVJCEo
QY4Sb/VSJxVoScaL+7MP8A4KVMXcOS2NY0k9FtdUVIp5xD26/JUbaMPv1bx8zgz7vabqSSZ4nvrZ
64U51iEh6QOi02AnDlkfhbB5m7LUWZUu47HejdUc5wBzNnlwi1cX/q1xLDlJJqOUN+7jnmOszHjq
y3n+v2yYqwIUS5bfv0A3hWLLuwC/G1zBo02tEo3/kVmqhYFBM+GEbRba67Rfhfe5rIAMt1z+b2h0
jZqQrtJabY4WznBPhII+qqbpLzk9A0b8bVhfuNPBWDcSAbPrc3FEgFnSQ984ceWFVdEmR5rqj/1i
EhaG+qHMBoGrrrM5VGoICe5tgievYiQVuEcSOPTe/rv/uwdqohD0/2+uIZr2Lg/KE4xMqCjRoCHb
ZmPDu1DuUc8veofWGYRwB3aSyiNKz2RdfuFlUbwG4+lBj64eUBJYRCBd8QTkeZBDahSoq2emOPvU
CI59g+c+hqJCvgIiEapq1WnBqy7bAUbrSBTosPqxx0TfItl+B6xFLGldg5RnZw4r4kyOby/fnetm
H88gu5TeYgi1kW4U6zOpoNNtefd/l6VhcBumbVyxS0MZMzrbGTMFRR68g1jyk/qbHkVmq2hfK5HJ
zTbTtL2HFpuOHmtYg9AMWLGMMEjTmlSPhviqmaCYg28TCeRsUku3UNrJ6Ygd3WiHOVQD4rO7Zc+k
4fF22qa+3h0IjRBKFC/iDnawgRxAU9p1HuUCpMLBy3hPtuZNZ4SxGizNm/MhlwlDYPPkS7kNB4mU
YCVo1KQsVHAlWMkN1XwAgvhbBOVPUolf3xfOYC9PCqL/XL3ml0PYkHytQfIkOJ8nRMwivLeWBftB
+hZ6Beed+oZvpx6c0b4dvt44IQmHnST9mzyKY4s7iZb7smj7pIfJ9ZT/z7Ql4mkt17y91cxev4Iz
9QmoLLcvT+Fr5DCwd9MYmIp0SKZZxYJhVLyFin3gQEA3dy/XZ95tcQgGpE9hCDH4kTKjegHP9nR2
RsCezy/lDTwNtZgQ6BHn3Xeu+tclPg4VOiy7cp8RyAYjYAbT0HziHDjAy/He3uzL1l4mo8x2x52x
/wRHT1Xik05MOUsW7XspCUpkfNeWFr5lvclXU8229ijkE7zUIYCkJ1GRFN/uEnqpZDaOMHTktEO+
NQmZD1m0j+PycLjAowgpcs6fSDijzKQWiIHn0pRvL5D0CmlAxpjMK6cAD0TK+5Bu1lcH2oytoQyN
LgP+qyn6O9tmEmzx0L+xz2xzMmGujyGCgx8uYDKnyK3AQhRpr9MEAN8RegEn0IwuFjSFXIo8JD4p
W8vy3LtG2zWHtyx1c7OmjQ3omc6spKiE/wTPJYoeEJIHlzxMW4bz0/+KygMQBkX9hfU/P1xdUuAm
IFza9ZfeXZgQJLGYe4bsDojP+kKElJ3NATCYMlaAjd2vZ2AeeNYwWk40bumSzV671dJzpEVctw6n
8M9VuUyHbC9TxZSvOLd3E432CdMZ4modCSLsXREBGTTA5h0SQMp+nMgZLVWVGkvoDa0SqtGPgPoj
s7/R+khXsOaATg4wY1fm5XWkXFEusa03yGFD/ppZy6zef8/gMeSyoleDkjuqs/Gd3C2bWXr0Cm75
dnhSkVxJdI/yxCcPMdpPWNVu9/u41wnE3fV/6IFGzOqU7zHldKRx7D9KYaX7g9ZU1OsrdB664KPR
GVUzpLWfmm1HWbGzDJkbdERrFYCfPgg6X9RnCW5IGD4TUO0qcm5NLg+8WinzIJMg/TKoRPemCP0q
b1j8+MxgWzvhPWE1AQKGdDw7CKisJAGXSGWazJpafLE8HmugCwzE/2mimW9tMxLtNr3Il2USWcA4
p338OPmgg5Vwvomrdo/BkWtkqiisEZo5Vwet8rgIq//9Pu2Z2NDLugWSSE3soe53VzJXhnKoNXGU
3pe6VCWnKBbyTh1VhgCEMrgTnVjQTvBjYIXvpblXAncOws78v+qnCH4FUojGtmzuWGMfuqiLTzDe
4AUb95vRKeRj3WBxEDNbbd8jaXqpd8y88g20bHFXOsKKc7gbfCI44iBH9bFlrCBwfgXIiIj05CF0
P9jweOOmLAjlTSzWYzpoihO0NIgQD9BDfkZJwM4G0dSpWNM5Y9hvVfAXAYZkBjcYmFY2QNz0eOok
Uzd4S88RvHmWQovmf00uXruIZSQDivxbRwUjGUf241BMCiTuR6dYQ2L8CNKabot5RggzBX2iBONh
nlafaRAYU1pd/D5hPzA18P+9OckEWQ8wHmexeVdvnpSD+WnhJe42kyAM1V6AkLkvDiachY5oLoux
b389JjA8qVaTErjtTpF7ln1vTO0wQVkO5vNKvZ49h0K4iXqNdM+8hP4TjYhRIycv/ctY00XN7NR4
mdkG1NHGdfPHQm5H404dzM/idHxIlbkK4JZ+Tpq9EVyf1qO1ab/yeCixflZlLpAk69A8oby+ud7L
2+YCt85ooCnOFDHi+Hx2gD4LqpFQBaxDWfyar+d/zvWtVPI/+FDaOB8xeDRPMDoyysv5uxFbM4cd
KzWhv5tQoy072BJ0bANUvT7zFKKf5b2LRxwIdSwdqdXi2nfyOrR7vuL+4FtDIbzoF3knSLLjSXp7
Q87xobt7GKAJUONf9pD4jEkCliAKOALKv85mpn0NsvssZ1rk/q+QkZ2wS5tbuVNWFaw40TsZrURo
wzh0jr6dk5dp8Pd/5schH/onweJIUfrUJgyNRMJXwDlq4TQCgxvNmccxC9gpUrxY0GoV4jIgSv0O
xwZHf4aoNqdTvnQzI+ozHfGav5l8TNwaypwp07gAmxzLYTAPrSQh4QXuSKMLUzmg5IIpVcK+YPkE
+en1/+yp58G17QFtAjVQ0jZPk4sihmg/wiqoUGMJB/3MbZ2fJO6fwgKZdhuXfaEoGAthcilH0oJP
Ehs9I3VGkXEtZcBYKmUixdFwLgzzhh/hwNBWWR4MVNQPpmoyDnbeGOgzPMLgfZOj5cv9syyOw26N
sFMYyvqna2FJ0EpLxVn7XFgpBR6zyYlksEv/wuW1ynoosvPeYhVcVVPGuz/GNKNSo5DMeTR1dMdr
v9xCtTWXiSZ8fI6cWTixcu+PCuDcWm2O/2ebSP4LvKZBQmsKM6HQXloPllR+kPedmacmAxuueyBA
L+rA6xN7F4cueiJRSMQSP8NXcsL8I8aC42CuQLQ8Ryhfn6960oPpDzA8AkCaUDHcyuNV55pFrEXU
pv7jGZ32Lz7V8IIe2yt7ijLP7LTPmzoy29oiaXVF48EVugodf2XrmyB5hmYdoZSsdfYzgxsPQH8G
rNa4kPIi6Xd+luH+0JQGH3sQmxChYOAsbUJw7cBsUosMnhSnfaURJrs1ScgEd12jsONQaVPtXzyl
xWE6ai2lldZP7Zc5GWoX8Q+B1uAzTRmjZKRS3zbMvVTI7GLh7nuHx5TBfxFgk/cBdkvHMqz5d9BD
8FiTA3tqQT9l0vsFT3o+cS2deXgdaDL/1f2c2csJ/AEbPggPi+euFAWjWEtTgrkiLlA05CzjvtmX
2URDtFfujK6cTkt0E3Ma0qvkQIZ9jNtGCaF+rPFZ7s1QTJh4+8ZnbGaHmi9Do4wva9+VJGH98MlQ
NIJK0kOViAND6/+dvO42bx7sFzZmK5NfIswVLaLnydeYbALoOET2aom1XRXwjXDEmjTcvvzLOA8d
SED2z1EtUVxYZGSrfdTnkT3pZeNqDySMsDXkncdojv9S7+TfDBhRGxbOW+DrTVmUVrYxW2Fgjk/R
8WdsAQ3A3R8nkWufVhy2uh6EEA2WAmmY5dmdTu/9Bf60EoqZcKRADGaTDJ3aKl8KmPWx1FNBGFTV
EgliEiIn6UMRd48PVmHJXh27FwZIdNqHTM/++ysXfBUyDpjk9dPrY23TxmaOTj1pP50dI1z3Gz94
Ny/aKM+BlK7dv/gUFvNTZ9JXFW4kmo+xG12Y8RrL8LQPxfEPHOnngF7VqA7QtSIKhpTVnq+3fSJu
/oVQcZPjaimaKDi78Zj1SM9p4S9gUGJ6DgBYYVh+qdiBR6ud7aqrUaggqKG6LZOVgRU/sdjTASR9
0tgVylqH2fQELfE9FgnuG8Zr8qeL9Zd8j+Qwzebz4WXZ+KUNzgRjRC5hmawO00phe5DFE3B1d1eP
1uGfNIezbKY5WemqVF0hkjGhnNxC9JPpdc7T6z1c5Bozyk/MDHYXg+K3XoGqtyJR4yR2w+DrIIs9
TJlIcqpclgswSnK4VBbKmMFBFT54sWqgGRb5G06inW2kJu641zxQ89cd6MNKIna/dyB8mTHZ1HR1
tttkgvX/be2Iz2QWMgME86IarVq2Gzv0o392zO1u/7GXItuXtbelehXm+jDBDMB/fKYQl/lqvdAO
nNju2gAZVllxEmuxGhUdHq3ndA6DM+wauV041E4EViM1B4fFfix6CL6r4ErMhmeMydZpJDLWpHGP
1mPOP+Fr1A65BMnJh9UqQdd91OY39x4cT5BDWoiUMbPatb6pIdT7/5NmPcS3ot59CGIcXvFV4BmA
aksmfmD3lwDJByjOTlP58gtkYzNiwn1PBw8yCMXUhoC6pDWHrFLSn730tS7Rcp5/yprg1htz0zmr
MHf8hRzkt/jHZ25KM0vAn30CEZD+F1q7Wn7odRbr+O7Z/zR3sPhfyI2pRZJMk31OznkcYBGRPX8o
e5IGWCJ1mMB92Hl+V4vIkv8ftBW/Xc5E9YuNaQGThfnYYmPmtQXoEtnKe4cOcDuwpwGTgI122nHA
7p5wz7F89O/cyeNm0vzxmQ7Go2aMtML5B0QqyCDpNTNrKGIkAhLRhi0/wteFV+mZl1HkReeTPjLH
DLmdbo3xQU+6yPYOb1LWwzHzbC1XTtw4ROdwck4lly8aiP0pAQWIkly7sTJazXRinu0oI/qofCWS
dXleqNe5mm1It3V6/v4qk+peDHoYDxGSu9Lz4MfpsQ/aQkHiCkP/K3Lzlz4NBItqEAIAU9S7Bm01
fib/Vyw+KaOa4lD6/6WTyjyRrZJu7HoftqGJnM4RCxC/PTN5y7FvTzzDm24+/JnwI0puFLL25nPh
TVCIdgXY+aATWLrtMHGAcQyXlKEiFMi/+ORw4H22foAaY1Ug5vlYlNowpCL4vxtYMdUaxEHcntdP
DJ5TUweq1PHp9JEv27nIf1D8Lr/QHs4F2/XKsJRIsDD8yHzG72CcKcJlrn8genLB6s9gjPI8/mLr
EYsOsLzqlC4ccs1P1b2oWAj7mBzD4hQnxVMgQZ6M89LOvWCuHMCDrjUH64AF933sEFTaIuyW0xZT
LhW7mFOtxb3wi/Ri0hW/UqRZEaB6/TDOGAJd8AWXBfmPEEIys2VyARTRrlHi2cu0N6DJVG3vqkE3
C1HkDj+etvBPleclaaUvpeF6uzD2xmnLU3VmyLKhE5k0QBDhRq7kC35PQz4gLnhD5/WBAnZaZ09a
ABxr0jnjTgw9Hqt8bXsEwpX58Z05LBGk/0232e6CUoe6KbsDOGJqx+cS2+CLASFNfEkn1ssFyqZs
dkjJ9GHIBYODBAgE0573wFSYqHQdaMNSWyiwV445DazyJ0hkeYYeZ2s3wSFMDqWJEV3wPqIiiuwQ
H9ZfBX28uDrTEN5EA1fzPq15YO9VywHBckApU9bj8yHQ31FxrOBPji6f+e7GSdNPK39KN4/Yn0K5
/IzCbPDC12EBhqmUAZTQbKXt+yxUUQ8UgTElyAmulRGmqmIwSvPTxNFOa7773iBJPp29ZKmaZQv5
ijcZAq1icMEf7y9QXVuev+n4iAMI8ixfuc2e2l99iQT/Epa0HDexFpA0fICVTVTI2wo6h7pADEXs
l1Mc6T6i5+x6sYxwERTbpO1CygVsSatQ/WDWe2qlCK09j5cRiYW88i7hzVVGoG8jxIEhLsEYk1jf
A/ymvsJ21QspzlZYgRPVMz2Sf0KCxxEDAmz/C6HOgV0P4aCUaWanr/jRQbzcnnnKD9afHcoBos2S
OvD974N0SDC0rAMWhhiH5V9iYcnMWr5GPDSFXfVwiQnuTKFwyvFL8fmuXu+Ctl6RBpqYtYq6GJfm
XVBuN+NU+/JGKGX/SOqs5MalObVRGPpYCwr3YMqDpt78eQ+aaPM43EGQWzloCgnnfVFEtdVSgKTk
Nq3ZxwAb+KlFLaSfw4ITxRrqo1606p30bDPiHUSzsQMg7LGT5aTEjyDlCBuMBDSK4MoTlA87ESK0
tc6bCDBZ/KvOdqPJ8pjVhlkJaw0pYjfgIbvQ/v3MoXHohuK7QyUQ0mpyp0Nir8KNEm5GPmeaGmvK
lTN5GIZvTTm/AWcfmrhEUpZp14cv/hNnMgOxIhZHeMeiSuAk6wklNqFn2lPDxUEbRJEh81092a81
qExA7QAPxjKXqpcjz5UhKr3p/ak+zwcazE0Fq5vZA0B+ZEhFs3dMYUfAK8SZElSUieK5TDnrJvwV
60H/POSxsgvpcD5gnRDOM29fTJ1F2RJ+raSWDcj1AI3Xb176whWHdcwfY17StGU8Av9r0MNqhDy6
r5l0/CskTqD8WgPFDbEczT3FQDsllsJP5ll9YEE9swuI22y63dJzRU5PN45JQJZdFFaRMkdJ1LM5
pNRK97GBRmWeB+1i4J4YSiCs15RIErH3e6DjYsUVFoTcFGxpcGxXekvN5hKSa2ZpBR9UEy0RX2an
BVKFqY6GkrYEwJSBFEIswqLoPfzhB+5ckkmpMMa+4VQ6I1+tm4mF1kEW6rhW/+2wnsNaDGw7a2U6
h03CWjG4rV84SZAqSXwQgNS3vqdBOgjDRMsHk9BBNP2h5e4PW3OwK+bjaqoUaeJwnFYk4lxiEx1d
gl5bGHNzMevQmO3rpR2Lbo9xG9i4yKjr2FcN92ZdVGQuGpKWcenY4t4Np2Xn7TpQypEeuAPqpLL5
2cYpMEX/z2SGTcSxQID/fG/artJrJEk+nOGYNweqehIRWGcT6GSg5/TyyGskKZKKdv2mSqEjICMd
IakpusP2VxG38ntgzJZFFdVp+B2FE52PFk2ttHv7nRlYYexQtlM65ISBSbUHo2Prd4j5RLOnMDat
h+p3VOjdp/qbvUl/D7tFeIxENGl4yNcLOV0jRq5cqNuxskP5E6NRRfcIf++SF+9SIdd8ybOudcPM
u5SJMx7EgQooAfeS1862fAYv1b0H5uwwfUzRuiVbcOQbp5GHP8B0U6ih1HA4RAx02oPyApVDQ/sQ
1+WiFMnTqPR1hO6ASsAxpEys5rJgEtgeQZaj2w8Fg8LPrKvAtrigNNZbvNf71UpXts8ywfSI6wZx
XZDi4fJ5HfX9rG/Ob7NiV3jJX4SA+my0BJJ1wHlr/BXwKKh5iVAachrCLsHMiNDaZ5QnSbSWHA/A
vAEP1LuMgi9drTtz7kmlyCZLO5HEcSVvaMmsalk+k4pVzSpoDWbcCtgMxTgR/tzgfj0yKiRZVmNE
vw59v5yd1hmPkeRY1QnvYcg/tJPHTl49Y3cjiKyr4pqU8uwses3yMuVtu5a+Sy58kwJMvVqkSgeb
vnPSmcjUNNaBXzLWCLLtEXjyqHVGmf9cwJV1iVKHjlVrmttSL7g+V+meiMGWRUiDajo3KoWhWMIA
YwTntX+w9Vy30AVXmt1cZ9umVA45YLfkraEWt4km7DLwb7+0K0/eXeUpEQg/4Iyhjj4gg5a8JfgP
OuCR/6SObfe6LDLYPu6pbcQoF4+hDmkR51isOmmUHxSbNzVMTvajF13WppVvdfQJ+47151kQCNhk
rYardwcCd6P/STs4QiKbidyMvk88PR7yLI6t3lf+rqAiZRKDasQ2afCb5kmW2bZ0tj3eNWmuPKXJ
echoV/XHKMKN5JdpTgntUG7FsBwrOqlMRM70XBIWnE5mS061Hn3EjyLm2K0U3kZNeNzy40bwJVai
fMQuyEgvAPCFgRC3xgdCIlaeGR1HT7T0EKGip+MmOpWtbIiTv/8jkxNCLl9ML6PzDLqDXUwiLgVi
RTQPCncDBQnSLNnxOVwCHhdkjRK+7KZpyd+ZfTIjbc2vxFiYqoYEj5ExXPYERHw1e/C3G7Wg06Gb
IkfP/osW/QlGv0GRwBFhWXXYl328vzkMF+xa0N9A/9oR787T39indlhEJuwkvNeD3PV1AuoEkogM
37Ul1kOnKbBzZjxHpB9G0T0LMAfEZZtly0kTM/xiVBg/dofS8ip+d2BiS9qg7oWF2gX7m5G9UDHF
dwm7CWSoALws18x2l6khFUCrbrd7FcNhuSWcz+u7A4piOb1qgYje7fIHsAxHc8zn8vLx3Z8re/kl
pVUKvkafhUL+bcyHUb+gwW1wG+BDfJilGY5Iob6G8SrIdSMJ8ugwXPEEcJPoaa9UkLvGY4QZQs1W
IlGYV2c1wHeDhDdbFCDQXnBfCSKoVp4i3RYptdXyXTkd9cGu5KFhTtWu37vVkM/xtVY0HT/PMt6b
DSS20neCuXqAulnaE+psMzNZWfssK0WsGUn9FJGj8KnyYbjwe96PNvhKFcP3wMYmVUwmuoH1CJsQ
VFpqWlJTeZe+gPQjR40+LZxNJRqxSYtlxZ+9yKITMfI30/z6jhpggCZN8Zldm17VkG2+HzjI0V8I
MKDvEnTyAR5jp+/9J5RlZrhvQUQfVgVCca1gpP1oQCxDZ/rSAX0mk6ZdD6jTaWAhVQGRpVARwgb/
r91w0wONDBD96ORTMGebt9EfvJIlH6RXiiT5PtV1zNhILxvmcJvTLhCUOVxDZcVZk1aezQjoPvSH
r5UbIAzJIACDDU0GXLoDLxKhlM6S1v94p+HpLmJskI8KYflX27NjWKUBYEQillIQ5SbSpqfkJWl/
gO9aWEO+HD/R2H4bijkZU2tZPItRFI1SS3Vt2NXhx3jKxIQgLA5QUrLAZIBybTf6+42q+jaVImnK
d1Np91mD5sRg9oCaAF7JbdjYQ+zTwmSZWpplCa3HsGeiKPB3dSCW/3KqNDp+nsqKsQoX1QMPPAto
cMHOD5z2kPiNIlcKat90kxlzVr//hkE809KDXRqToQEqEOUEMajq1qEw3gLgEFE4iihqJ/BRqwPy
crUIYzdsRe19zugl+SIst0pZ5VoiIz3Drryb/yp+Lul2HyGu5WXoSsUge0u0lVKIaGOaK1tYIqbq
CnPfhXZJZgdinTPZjOJIR+m15mJSS6GD+nJueciG7fLhfMaMMOYBjVtuJRpGfCq8MExOlNO+1+NU
C9GScGB7evYsHpiKnyaUanzi87VaEbkrBtRxXsJuC4QIR9mHjn1cWF7/qaZFWqJUFtXCk2prG95I
M8NIXY/Mtkp1jL9s0XDheGhdGBCKU9+twl0OYo/CcYVWtZjUnuJwI2cfqQcKm/0A5oeks9nNhyJ0
cWdrgeJaXMUWVmvF4U4B3oovCoZs66TDsxS6VgeyCvNWOs6D18T/zZ/zjjSbV7qCxG1KLKLaX1ms
tGuICutbI0wZm32WPWdcWlx5jOK40rpJGYSxhew+W2OUK20R0vRzYZuU7xadpAc7R1DreLDJi79r
xj7ODvknpZqoCjLyra1fz0BabQq/lTKOHbDDOGtTLzf61uKvIER4dfXiUdFrBp8SKZZcEzS2x9Nq
Ti416I2mC90rsVCGpa39taqztRvwPppA2PRxDF9SB+14gSOofo1YsMAJkknAAhEifFDyKePNRGIx
Tj9zqsZ1ic5RE/SVK/vPOqhc1I68m0XKjIouvqhnNcXIRIkyWPBPaCcg3FGBAfOouAoJY0Fm3usw
Ry/pY0vunF085z+yrLiXuWxSrlDomk6IQVsTbWir+bc91yz0GEOPq3+jzi32o3PoWEYVLfxB94on
75NRq3Xz/Dzju79cOcGnTaIXIJ1Lq6BQw93p3vt3VYs6jaSlrHa4nCSF57jbD7jjqSxHCFdggIX9
KUKMPCU+JPbZWDfhGFthmmo6T0PG+tRCVdIabcru4I0t+MsnLTuJITKgyJB+3sR3bRjUizNmLbsJ
2XoNW5+BT5PzkQ0LyhaKo/kE1Lt7HPJJOzut01/uplqpuK1+y5udiTz60B4PPQhUReW66ZTTqJr+
L7I8YrW50g2gvomcX6xtIZbgxt6ypLEhoaqzc/BbNvR7cWnZE0+I2gWzBygGLqTdcGCnUMUAb+HU
CSCshzKVgbcxxK0tsiK3nlZpsaVwN2ybIoHXEvYujC8PiFZaWW9G09REh3iVhWT2uzU8WZS41dTh
YUXY97nP79nK0jSfq69K6zqVvAVxnyJutYeDTZXI4LU8QPQXhYqyL+GmDbDOG+28IfwtxKo7JaZF
QreYw1CKXd26Ci0+oZtKvAp+ghPYPtR97mfB+6MB4JW+Dn1EEf+gAbwIIg9/3ktlpjCCTfriUt3q
/RpJo582pr52In3FU2Fe8pcnpZgFa4ZS+0PVEcWd3/q5mypifOrvStKpqY8b8MAqbhfstAK/HLqG
Smo+XMtncD6okmqYA+6wwAlUtBXFBak7uuV6F7iguXcpE3gGESF2UYF+svk4siu/EiCZUlnmAoBI
07tLfmYi2OGiqVorxuZs87c4PVN+H0yps7/KgxY3Czh0jE+YKRXLnq32mpjG/vPK3fe1igBS1P1D
6Wibus7PFRUhXjnNm8KMdP2wqJIDYf/jXjFoul+k1IJmU8Gn3JCfzVmu6ox+/yjuKx1auD/Rk5jQ
kHCVBu0vbK/gO2brhxHYIb5Rpkyr1e/hwLnrRP9oa9SOB2ZzXggP7tu2Cf6QfvQ16erDl0XAHOni
tqgCCeYNrv+N4L9Sr1/6cp5sqOKXWz1LbgXEu2o7Eg9CzK06T2vtgySuglRqhMsRS8ZqKXl3/gYM
/NCmv+adDC6y201lBlXERL1eF9v/wWEuydTqni+OB+MOG1ZphFNEAAtGui9a5gSY2b4eghB1u71E
oMhxSPJsMFyVJjcjUzn9n3z9+Adjbnwdg+C6INS/On5zif4ZzvOuyQIvvL1q+9+C7Z9CEJI3SFH0
ZYTALLcaoQu+MyhniKuYE813kwxopJOyunTZ4QcJce8kANlPt5HOD/xASs5FT4VjXOHrgLyvAdix
db2alcsM/04Io1eV9dNT8fHO2HcftRUtLQU8/mrJVHLaWj9VUtU2P1u2uJRF8MRL2lqH8Z/kJqsI
KMeA/quirCaK68FfxekaXeaj3mrDsBLbDYOEYAD6b0W882RtAH5unmLMJe/fDvAkesXYVFdx44Y9
Tk0myTwqqeZJ002QQi6uqplPnYve/9H9tVQWtahWp/zzRD+Wv7+R+1u0rePAYfM/wAJcw31hVd4d
hnWQyz/IqLb4BGs07EVxWIvnJsuSgpfTFw7Zd8rl+hzRXJFZjA+XBQDBJL7voSDjFN+SKWW+sc/e
oQIeoqgmMbEksFOvtGlrtkNcx7nQCKdAlMuFZ8pmnn71IbPyqQuMl6f+hcHDcy95dtmgxcRhdH97
nJgdy+P0xLgjQ2kIQjB/q+eDzQaFtfndZnT5iBAiJIAybQt61DsEwFpsS9/rLRmC6TIm7GGsOvYi
KKEfJ8fV7USvxgVm00tD7wcl43hGVfzy7Zs6DuxUmzYts9uSSHvhQwjYSwlNDj6C7VEaivcQsB0/
UkqpwY6MwY4YTMq+EU5RMo71C9P7tICWqz3thpYYu776H1/6GZESPynB/5BTPX84RlEsG81jGiqK
7oleeKgvrKif3La9W8u/NAGpUhyVh4wW/j6R6agMYhquAS9Ev7cpWOkbiG5BsPI9ONukMXAlW2TT
GC4F7QKp+iGbAmP0qPFy68oUmeStF9CMAtNBqmWjWg7wV2e7QUXqBnygnrSKadyrvlRXQPVPB2Xk
YHiiQ9+ycHldiATgFenzM8Ei1Q1b8kIOItF2mo4pAXlbNDtpVxZ7f5zJEaOwyREX75w/Vxg2KeTY
LVgPVKdRSlRXh/iYK2H6N1dUXQMGRimf/Hkx19mwatsP389JbYgdW1iK9O/4TAvNT1EsHJWSUftM
Z//okt7dcw74SBF1OkWBb+uC95k+DLTPvhkZ9UlguYfm0KWtlrb07j5+05wPb1xj+2EVjcbbNxPI
h9u2gzR08HiWBI4QsRQ9KaWrygo0jmt6fYcSVpNIfg0p7vhd5KkggBMpwCtKLKNK5N7dkWdCPlKN
IXv+chS6D2Ft4aTvCgfpVoz4vAxi8Xr6mMCw/EpN+diVHW8Cflz5Va2DPEfiB01+oYXwlMCiQ7bc
cYusf8YT/K32JsqeZ8BYVLAuORn6ZXDqok8b7QdXaqo/Ebg9MLy8jc179xUMcADn3t6HRApX0frf
ca90iEV+IrNN/oJ7HxRq1z51vQnK8aZrAImgpyFknwMwXXNjJP6nyGRGEj/scv5bpAxbmYbjwNM8
srN5QuuPhgsoUvkJeS7f/AgkbXWqDcIa4x64QWbAFHbw33jlqaaQP0BqpuxCiUZfM9hHGeKXwqtB
6fGbNA+T4H/sRpwGePnWnQ9ik3wAcHcVvP/idwSLJU+bjmI9Z7a8yt45TyjF1t7sgtlhDFbqnfv8
912fQZEAytdRHP/96PXL+eXZVMm3nH7oa9x+PVuhf8Nc+zEtQAVv8oebO6r2ntpFV20I5OisFUvX
3QpNE+bGGO1S5WCawk8C2ow7IyxsvjT3U60Zu74XQ+aMudrIrIBUb+zZD04bE7C82V56qbSh/JXU
/Om6WD+tr4/anorI0kx4ckv32uhMRUAPNPR1DerK80aZAHMe6tQ/jKz9WZlsMsi9r71bSvu32r14
+6WTdavpt1eijctgZ1dQvqvokAydY3YFu7UI4YMnV1DqOtnFkGMzvXcoBE3JdwCzdsnrNRoMfJBT
KJBrYEL50Mcm/WryPaKY48tGXzPuUSGC8QSLl59Rc/8cHJS9lDv8CDKfgvmWhL4d7OvGBYK/CDKV
OkpLVnxOvsmJnUzqrg9kZutv9xjEjy3BqTAkYXCs9gfkbxkTal3pw07Z3sEX/6OjWSRQl7DjNm6b
dr0ZiC0Zku3JNzxkJ0ofVBT4cl2OHR7m03i2SzIHnEgtbiLgHRJwmor/DqEj3D3OHyOJm9eTLFLO
AsNjTFX7QLTfHs4k0SijUvL+bRH5iwqlmAeI+2v5Z7TC/yuqZK1/SOTpfwmnDRL47viXSVJrMUli
MxQm86hs1wSnZ5o/Arh7ZiBhuVzfayX7jDMZR0pkP+jiaaY9lDknQoWrCmaaVp2SvcKCaBpVD/iI
E1/hfamAmg7nOLye1DG8OMNLi5cZTP1+NWGkRfcNfr7o7SJuASxpqq99xrS45dFi5AHmO4xFpsWQ
yEl1mW5WJOBM81lxZ2hleve6S2ZIldP2Sfs17zorlHTEMab4fkGMVbll/NuV7iwfBLlbt9eMYVFp
tX+E6hZvvHgU6Suneby8B//AxEMugqz99yXyD/kyILtWlEJmkLaJKU0fqSt9yfTt4r81D/gU1Hne
x9n2ICM5DuSrdzwcuF6nvYJ5tkPfe66mVwQRsgDx37aFyfSpRhe8qhnUBaAHS92GnLwKU283p5pC
BcdGtvB2IFMbvXgG2xHkgtB6dX13hdlEXmCQivg4odmLf6Dp6Vmm+vsdUM4afzgXwmsn3qMfSsf9
Ne0nTjzkJ93osrVC4ryAWEvgJVl1RCnTgajlslIl/c8iEX6UaXBgQttpgJWjD7XRbXUM11n30C+R
P67oCcI6+w/gUZz4YmnhFBbJMyrjN9H+XWQNhETJslfOcmgfoHNjD1s4Z0b3Ypa5iOPW3ISIbA8F
Yc8SPXAmIhGUj23tLrs8HrF5mY00RNgDslntbJQqByWxFfvfUpHqS5/cdv5rl14dMTurNZdhQ64H
uWVQbF3yUQyTE7Lo8oD4zYwYSRe0pCvKc6kKI1vB4kgPRZpQcdUDwI5PFev2SZutubIGbzs2zomy
O40FcF0HcKxuM8jpphrNh5Jdd50eFtSi3W6tXXxX/9K0d6hyRECOjJtfx8fTqwjSKoAZdRf/8NvG
FGKg3D1e3l1ATCOezC/BpWiUMY3NTzO0Nubdtsx/CS/KAqlf5q3TcXxV32p98EAzlt/ZvzEHDQZW
nr4iIX6XnaHhjfkOUFA4ri2A6KZ/x4Nw6u1DxkvkYj8pontVcV/90rJ6KBocqWnCPa5v3seg+zQC
6TfuaPvp0qL5KNxWteYpmjXI+b3SEineR4yQXKIRY8teyJFpsgPmlKrAHQ6+9p/0+fQCBkI8hSzm
nODvheY2LK/vI/LlhZc0R53At27wAnre79zxRFt0oLyqewpYelC2HhbbZsj9RdqX7Hq3/c0JcLZo
Oc+BBfLI29dlChS1aObkXa+2mRSsDEl2MT+bJyT3P2xaRiQkQ+eN3R+lIsLxReqa0TqJgJDwMJf7
uNa254ZeMEWqz7kyyuXddhRuOPBgkP7DaPYwJBpRoMS96E04hn58YGDlWA5cSFgZ7+T8WP9qNUaM
tkdUdWOgpfuJOhzWqTxcm6rrnY+VgJypQCCSa2faoRmBRmtmga2flY9fotbXDYCwwCJOiwxeGZjX
JwD/Ni1pt68XqaZuDJjnCpK58Tr5sE4csYXbOE2nVeQXe9hu2iWufYR3/Ajw2pn5yq5Gv/RcAw9R
uR2BgE5Hz/NfDT43YouBdbZDMhZGC0Oltw4BlCTzbm7PekqNZbLxbFzUZm0/Oq+KM5q/XAICOvus
xwHXph1zn+lLRMR9YQ3c31J2mFneNJG080reOJmPuviyluIHOab7VEL8xwQ2NNhUiL0u1aJadHQB
/Ti8Sp6nLJ2z27blzaOgnO7wXq9Q2cE5GvF9VXUn+pmRdjtyJ/b+tOJlg2XTBwUiBNmMwT0gb+oe
6ZqfxcLq1lO7v13PjCJLvLkCsczJtuKQ8tn/d9x2FynNRTxwA2jv9+usJ9tdfmVWRxsrs2Aa0+y6
+HWTaU/oImJJ3z5oZQQgKcbbi1iavHmc5kRlYw1aBQ8HulnEkU7UT4GpsYl/E64zmbwSsxd4a+LP
umtImJKmTeOK3bJjd6LiffClEd62MbxnRr7OgrRowPzgjBwIeWykD/Zlo/ZRho7FGNqdbJA4OzhH
TiAtMCdRADnEOkjZzv4zbxgOfhJA7GX/CBYH4++NeGjAds45vNsS5CAafirWUYHnkj+Amgd3AzNa
D80ij1j4GLbROKfPLnWcBGgzpxc+KcxH/lTz8A+V+hOjhxCpqso1hFiL+i804g/II2rMqIcAz/1/
LMxRNfqD4MmLAqr5qwFb1EdroRvQv2kOXkNPpqpvT5CwRMQ1Y+xQdOahkOaoCAMhIjoQXuJjFDkl
SJmVZ8UGb5HuHOk4wd7HimnlC48M8e7bJMeiGbCYM5olR6C37xG1JbZGyAIqcle1Nx7HIXX3z1TL
ulljSbLxfxNowFvaqJZ/YUV/+AoqnL3cva+fEKPWqHLUPaFbx+BB+zORaIzQJXdKVVRVOdtHtuN9
8UOPurZwMxJZvhnMgNpznCSAW4TZGk5NWgMFzOkLS8akFRC3b58wrM0eT9MyQ7GFz3CqM7Pd/OTX
+bAafGm85ccNUjZBj5kyf9e/yFPMEPvqENi7o2+esRHwQF823+pBL02whfIjLOKk8weFRz1143+W
yWYYwfxU/ynD9GeE94YwGc7YJqu67V+jBl9ji8+KWUQDDfajMxJjPrqCyrkkn/4aVz8uBuWfs9Vi
RIbaFeUYBJWYJMeFJ2/XiE0pXer4O3q6zu4bctKKi39EfaQ/0ZhWjcwy8a42SVWi5fXE54OXVt6D
pfXpqIKUKSWKk7I+8EdWzEG5YVcQKMzm81URJ+8FxF/F6iQg4JvXamYwwN5FZ5Q4Y1/K+TA7J+5F
Mnbz3Ougch4dQb8GbO/U8tkW+KkIybk0LEH2s9Ils8koaRt9010q2rJ4/2kaLGoraBmLNOK4rb5d
n5ffG6rZRSyjC88fye1BLL9ie4bb5cD3Nm+W+zPGwiX5NWp3XGBaVx3XMXSHBxN2nSBfNVyIn/9F
gcxYtsaVtESkztqBniiXhw3xyl5vraDLclMxMou8mt7LtHTmeTkp2mVd6QQw1mJqaoC2fKPoyHkB
BVOF9QuA10uqcSK9ow8Cufpp5HUs0XaQMqQKHRE9NlJTuEL/mB59xJ7Fkih0tMf7IMbfCRNCRWtB
UbncblCo3eO07aDJMTLAyx7p3/ciRzhtoX3VDL/U7wwJtf0QaO9ao928effSJq69i0GJPp6EkIYQ
fKeyWAdM/59uYnZSQQIqlYnQTThrRoAMxMIfpd/xJjUrCKLV7mQsOlCpS16etNTusmpghfYrucQH
aH6BPE7pKvDnZQz10bibvPuLdn0EDyEvDBvAnQdPYRPajAS/hhY1yZAawCDcypTMf2oQpt7Ytv9t
RPOaZp8+iDWBTfuoaZM3n378yP8cxE8+Q4aBmYtspOBccy1RyClyNOcGiFBBGpMOgSgiAGOZogu2
ocxO57eTvTNXC0fsGQcd7D47Y/KFK3Z+J0SmwhI2qE9bB5ymQuZdb7BRzodiikdizC9Za3Z1R5B6
NfIcJWfEdjhsKK5Fhaq+j9s1GMXG7bY3Xz2NeAicB/rxkCUsYB07Ia16oX9F0s8PvCMQ9Sy5Ii22
lCsEwn7VenDTjQUM43tFJ0IhjfbrmjqBEmpFm7zsRr1176dT2lP4Yh2YNfon7BwXmB3i+2dGZ8am
6w293KH/E2zVZKjwKeWL8j2LzTC9izup+z1k12vghaCRtrUr+G1Q5DkFD8JhPFZLMus0KyhnvQTX
uLvrt+zQ/mW+MbxUo7ZgqLHZG5spL78PyAo1uHG+R8EB9ksfO+7zI9SDIf+woeFtuSNxwn8KHgLR
OU4+4Au3abBYTCOvYOPksQ8A0ydJZdSzSNs/SJ9p4l5YALHTRO74bTLQm3lm5ss2JxslD2w67y/q
dONAClAHJzOVfviBNM+FS3VrbGlzafmGoLKJcae3KUGl2ySS9JXdRWVw6SxWoSSAvNLhwc4L9Vip
dy3c/HbnF7lJF1dHd87wVHt9zSgCK755ATWJ7Xcat+GlkJ7L+/LeAiBqt24J8G18UhZNqgkcPQjm
8E3AWVe5Wt/dLe85+sR3Uh6SiVVsCgIkT5MHBDfOdGYlzEHLwkW/xTbrh7xl3aVaET3mun6vTuGY
zwkEOIoxhMDAeoY2rKxQSz3NMPeGOYVbKPItH9FSXQb6tPJngwX53eaLQTH8SChyC1bbmgaIT/cV
aN4yNCwgqHguNjmzjsN4co5zltaoMA+dkIxQaxoVf0KvuUkDJFQ/BEK927hempFG+D10WefXW1ZU
srGVFN5O7bp+iJT6CiPwXmXkwmv7edZBaqgADkVhPRDTXdKpLj7rP8ZNW/s6/0JvD8wq03UiPmAc
RWQaOHisOnkPiwAmPAttJcnVtWteLldSm4FBzDz/Wy0nNdL8LlyRuUEO1JwdYz5S6jKY/6e9nLcb
21GvVqt8770cteMXK0NDOBHW0lKeWDe3jJYVZ+/OzAh7U61I5Hta3RzXXZQluP584DUW5B2WTFCu
E/kielaj2HUcJcT0OolScb+njxxDKdsEf9A007xaWpgz3OH8XLK5WL8RWeD3avo+Xk5sYCQibZHI
mIMv0oy3wz/jmyMEtgDjbgGJGWVU7Qf7/6NUFDtbdjZH9YoJ+U20skh21K4CZ1keYprpBqnfUEDU
fE5c1ThWnI+whd3sTap84RUPmKU0Pm0SqdTFm+1OEy5V16BJxy45Y6VgKNTdsd+QSB88/7IPd4+x
dSiZ5b3g6kwFpFoPWfWUGZPYITiRhRJ/Lf804ew1ozwLHuXWCvuFBomkvhQaFvSyebH4tWKC4/uY
abAdgyBriTlR8u2qRBp/f7auV+BK4WFZ1yuGpJgzZO3zum8w/Ioa5TnfgC3sWy3pHX+etBl7A4aY
OhEVwX8Jk/upXkA86E7iIUg49pK9l5oa+QkTcm/PlYGcYGqpb0lYBQjOTfSzCNVQCXz2gY1a2Qof
tzhqy8FIalSPrQd7aF9wd28VnyEE/H2n5LdU4Dgby1eXhcgV8lEL+Fcsb30zLtPqU0DZ91FKXdCw
+jX4SgvHFk54FSSt97VeaPlJ0Q9CxYGTZXsbLr3r0FncCiGMl8kRxfs1jrj8kFL4od2SboMI6/Lc
5G91ELxVX87YO6EoOxrGkNFwzkvNa1L4tQJijHjYnj+KCm5VckjIJxngP2io1f1v7k0BXDm9hJyO
E+FjcmyVpAPvo2sCvmGsuo3dKUHb0h58zmJx1J8blPHIv0Rfq0aYuTZvSqVf6w80SUeIz4qOEE/q
5+6ZYB0P8GzxDCnZhowaDL/b4EUPhOKBw5DBeYJSwsgmsiQgUQL7JkwFKTPEpvHlD+dXZPiLV+Wf
QWeUIVyfb1ZNwpkkrst7iO+w8Ztz4UQjAuRn9RK0PdXiiD3nztAJ5yv7AYEFCEETrSAQp1e90RGn
QfidxWZrcDGgqyA+05R6xFTuMtGxEoh+tJqimpsT6D1WjX7Pl9hLP/1JsfReoZEXcQD8JrAUQq69
2/nnzxIjDfN0LNir5WlqpoNI4EZv0x5TEL/jqF+v7HyauO+kOIpiuOMBfTzvasTF+qgcossueKXV
T+cXgf96QWl4fG5hw26KyVIjRXjsUQPo86LJljhB87WaELVEQUuNlsqG7w0xgMyLATBaOSPF9hVf
PZw0ZY/k6ef/UEtMYAcseSdraya0uC9BgJbLogc178x9dbEdk2TncE3lMcAS4j2WrevjuulFMYW7
0vSsvwEXTuui88FkdWaxDZE5nWDGdCNrdahIxcwgzBCFv2QsCbVgNXIslIhTYiL21Kz+qhLRNLdK
ihCXYk0U9z65kE29qnVZ1WvTWmydnzzCOHE7gZUN71B+6DY9P54o9QA0xyVbibID+SGuadWe2mEU
TPzFUceWmfSDliUT7AyASChY18UC+ulJvvZjgueR9Hd/nx08YP2x+0B9bRuk4GtkUD8bfuz/LkHs
GarTgewElF1vAsrq8CP8zKiz/i8li+U3cCsKkgPHZ7hjpo9pqHAagOn9YhaBAkI+x55jAB/+P7XA
edHmWSw3F2xNyr98lDgEOL8iZrSezpYRFocHLkL3GgAolQrAgTgW5CB/sI9eDBnh05mPeuBBTgvn
hEQySMyn65UVyg8c8fvP9PJaRHTUGz5DYjm2WX5MDXk6fDHgzxni6AGrWRLbtaD6ezhxPKXjtQDp
iSbgUQ8Y2B8M6KxKkiVmfOOXDfsm99YYPgJtC8HzpkPB6AHxB3j+XGvfmE9NHG/qUQ+mO5AVV8gc
Z/VLDbJ9ebhOoOFGpAfbg7HH0QjJJ9FOIMi6ZsFXNxFGRtd9w8EWf54cEkps4KVlfZkO3lq6JnrL
Fdvw+utGLtl/6KJnn8yX7HET4k6PU3TqfgiOQ02YuBmy1IJkh/fusWQtCO2ij9JYE26vjajeN8iO
d1EvfIybrY1Sev9TXg0kDgLaJQ+ndt+4FypUOrA4GFV0HBBe501GOndT3dKOM4fA8k9hRLF3mIX0
9TcQW9zRiSCCQh3RlsWwN9i6k7cDAYRoWwYOYrxMbEzoGPle/A6joy4Q8POGWTA7jhlRl/mhusoO
UP6xK3tLLjdUVO/AgbJtFM5+u9DwLFGxwJGHSGzngV4FJpQwM7XVoWD2IfIeeZxL9I9Qb2sYHPU1
DuhG13rmz32kWoRrQGbTw3wdxkR9U4iNGqMlSbeaG/ywSRzXEngiNhZ32gqIpSUUHv2SUGQ/Utti
VW2Ih87wGzvVfGfplzVf4lez8t070yLmL9c8bqOGQEroXz0rL7aC8JrQBuXmbTUntXMM9Y2yg3wk
fEg2gm4Y8RiztdO16KGWD59gu0yw3sYado4U2U121GILf7LsCp1n+0qmZHRyIp4AIMaL6jvGoWjX
GEgpvFK0YYkIydg+rr44HZUa8+0x1JKZrnUkh9Z95uBr0o3zhUrJbDeBnM9pzrR8XzkFJBzX+to/
eNUQbhHBl4fU9z4VA5bZY7VNjfau4Gvt19P9CwpGDAsdlvZ+40m82tHhw7sqtYikfliFsMMjj3xO
fMXBkd4sc0KPZMTPKDznzwwUbVK1oIG2QY6ci/h7YMPENnv5QrdwdNSKw5nXFEG11gm8eVBXJtHW
cAn3S2PB0oxRqUEToSrYNdinK1Ina3FDvejEUxTSwksrlmasJIGBXEQx1Q7OuhPaSbJWbe0n5sO1
9K0+JH7eZq3IzqgC2u52YQ5sHvTwTRj2bkEI7hOsA5RopVU4vj8W6uOZMtj7oftiTs7+MEfgMPaI
49zXqMCUqfWrD/gopaM9k9cm+v1dBcwo6ehofNEpv7bRGz3dXEItLETsM7KsHKnB5GK58TUSpiE8
KQHSgXAIw+XYsXElN/kieLzWjSQNQZBBGEi/NYZ8vxNjZBEPeoG0Fpg5uxOPuzJxJ2h+Dq7JhwTN
5svXsQMzLMSjurTVST9wiLRDd5PufqbNaV63dlwN8N2+q10XCzqbSQ7UhsWFC04zT7pozz8nkrLV
sPnFRwodVnPfH45y96JpLpUH62OpoKxGUwV3gugU/bSweY2NuTRTdtYsufLS/jEIWSonp40cGNKT
0j/CfEf0V+m6b1gKgC8h9JpVk1zVikYfTcfOW4W3d8aU2UvVYdOBO7qUr2o4Ftp+lVYzBzlvmUCT
IsFGaw7tC+itLgnk40urt6W7rH82vhK/JUBUbfE6SkedB3QsZzwkLdQshQvZrTqJr4Y4XYQWh3pN
l2+RBgg2sZktSyqzRQ75CLiiB5Ug+RgGH1w94rIzFiYnp0tLKbIU3ywOecvsKQDenfdGjD72oPHk
WszmkOKKrASS0aYcixVyS0zbdE6TcLN3eZClb56RGnE62jIBdxevxnYzr6892waJhHKnlk7IKSe0
6ZaHqZu7IeDOxKDkdZAc9GGNLsUhUEPVop6IBMgTz4/wi1BLIjaP1ubtn5LwgmQ15uP1Sk+wITXL
555KK0ZWSwvT36LshDAK04rqBxHpQwx5Z2ksQ8xQKjzI4Ho/USGo+Y4JtIdykdRsLHE5+ykpiUfQ
z/OHlpStPIb0W1a8qiL9UAl+Yaw6AGpZUXJ2m1MYxIZU/u8Vq9H34kg9oLrEQ376v6bQdJmG8XNE
e7DmeS6O2gfo+XlR5hSacYqB3mqWk5Mh2K6hM/bFpG7nSwPUMsIEN16ZUDIddkvNlbj5achKiU35
5YzUzlDjgHjoWMItBvY6GLIju/01P9Gw5eww6Un9G5Qdbu/83EYZhrjjneUO6KAkvD4KJ6UpFVgy
COB5RgFAyJlZZSzZlB4XvFFYR+gloz5jG+eU8UGw4RZg/B+HSavIgtchnfMytRvqy5WRP6kOQme0
CC5xy8gRZ9qg65YI+OteXgfDljB9uxIfyim1aj9SMmaowhHrCY/WmgwOPA8oCtX/fmrecPj2GYi1
azWZJBcTF+0zMfR4pDYr55DPQmWNvH6jPHFSMhwuYeIwcGuojknCxUGRYXpzFlv/evouPbl1yqr4
EUjNwK7Zwsr8ANwnKdDDNvwHCWT5c+E6S6QH8UMZHkX4p6vx7szs/8Yqu3voZQjl3LRWMhApgll+
7vVAHvKo595EWQzFP2lc4qdCyaDwN3VaVNrK+c3oBB83nXlXorjdvR1jE6ld/H+HPyHPdtDTwV6L
gqQBjg8fC9vYjSCZX9guD01Kio+sx7oJ5Wp/+untvq2ZOS2AZCKvjA04sFMi7h2EbcbK66qkNKJz
vXxIjd45gz+cdBa+Iv5q45JB7d5y7b3gySySOFdW42AIFFbtLEuXJGvLvqhmNPrnQGrPPo2zuoJp
NmuaIHw38Q5zFe1UMcn/Vuiq4Wm5y5M9d/qk2P5fS0WT6foQcchiXxbNRFqy0e6uriLdRz93EZEH
19IhqF7ZysviK1WtIw7BhUi7Fttr0o0VcTF2GMx/FJWMhGeb5gtEXBt3hfcT2ITPQaeWOxP8vCH+
FGOSK8GyL7JyU9npTxzHoODxfIMY2EMvVM7mZut5A98Ccg7fpHDYoK2HskPuAPVy+FWxAh/ubxM2
6qEXulN4CLZceUmLjeqszvE2GvptwiyoLfDOlSvA3S2erihdO62y6+a3qAEj9U01trgTcY0fQ/b7
krq6eeEk39AFwW8wfOqtqDFurAzXo8X72SK1y7hgkRypp/4qPQdmBks+0CM4bfr1hSz39UTOo2k9
OXLISL94rnCDTXqbKC5Pv0O5QhRybtTUJaXbfNbtwTXm53nmgh1fjBwZabjIAQ4a9lg21Jkte+WP
Xs5ATejbkO73q2QhYlJ3Zj1NRAUeq47LhmrUkbU/P8fKAIpA+6eKTCAt75KLGqP8lbpFrdEhG+v1
DSwK4QdQHZVVNiFy98SO/jTIVOGDHDRFFKtmfov4c41gxIoW2vUwpJfrYiexobfI03lM0ij1HTfn
Uz++IcT2Nca+xRCg47F8pFtf51mHXsYvk35wtQULysPtatljRVR7iWpP8C5x+pRU5uNXU7p4Wuob
4lGMot0nfQB5Kz7lvgVGeg253xSV4AIsAtLh/ychkycgi4riZUx9pfjqhdycCzplYk65YBeFxB7d
4dJ3nM3mKmvcDVL0E1MWRKzi/J2yb4Ih42SoBxhkQeGiAp0376GNpB5mP9DXyXcUgH83gdBWjtIg
NXXNuWqiVfWyEO/3ls4NxUMBqvbBwOv3oCIAjrZehvXrc0Jjuqc0gwvsEHfpYHyxIOggFbfy6XxP
VNB242bc7yGMDa8St+9enTYxDGxTpNCJ+TTgt8c6gHSiXaKHCxxUj6T//I/xggGOggcZtdSOOkKI
fq9B8fiUN/NS2qYc29IDafV4zOcbWxHFW43U0NdR170z+9dMawYe1M2TcHXzHE7EPBVtaIuPIIP8
geFNpKibYyQqk/UI+SlhfbTPCDDEKmHMtYdWiX9C0XV7YFgEw7KIqavnh2Tz9GhnOTvDG8kLG4M2
YkBIZLgzVaVO0hkk7S1URzTM2ktr1bZcnXqzZtHsTnzxQ692grtF0w3X9Fk7U24pz4a6ktyrPY7K
82IIreRu6a/qgGkTtaXPQDr1DqwW1+ZfyIf+XDjFVjpwc2aH9p+lDaN6N0unvHLAKW2dEsrMFMX3
+Thfv5FD6hdLTvFCdaLArXcaOEAJvfmTkmLrUrzWCVfCsPoz90I1MSjVZ7TIYVJtLLK/qytszd/V
IxSSwl7RUOTXRfprZTdS0ODkf2XR/ZHqP8HiNTJJwIVJC5bGD/X2KVO9JcmiWxSRGTS/Bt7T0+wP
l82wXupitZetGps/TWOv/9Ma2BJl5Tu27NVauoYPWj8oNh7NHyorYRmowHf7imV/UF/O6V7daswA
1ptP0YVOzex3BOTpwSc0T/R6DavzBVcSgImQw6g890DwcP5CYP0kq7BnZfZMhPvctDzpt5HYMSGQ
4K/o+BlFkAxJ1y2GlbaxtTXKC1GaVHAtoT2oOnqBZltSEM5hXSlW6nY9WCCFBK2Qt+QLDH602yH3
FfAvH62Z7P3IbnlnlvgeU6y/a9CQanftvZ1c4AG+uoYOWhn2fDxXEUAXK+4wf8+PudKwPvmokTsQ
xuQ528dK/Fd9RmkNDT6+8wsJ7TLHNxo5yDZQ1J3NPQAVPlxGHkrqAZCc73JwgrNPyKgntMcrwxSa
/DOzm6gKV8V02aKlQ3q1dTF0n1neZxGYHg7BZ0Zg6AA+9Ra9Qmob+gcawME9RtPO2Q7wSUuFQ/F6
rUwzqvbfU4MwWcLvDdF8qZSx/oscDynXIZZ4KZNCthTRXXYfX43RWnUQ/emrQBQo7bMeeJzzjhjg
o2+NOuZ3sfVOOKcP/M6OCdB8k9BoxG/1/jp98VQSOK3KPt7ym2XNVW1bmojZxMubB28cno9V18JL
6OpZ4Onvok75dXODwkAQbiPbzlPonNlDp/FR+1KMH2pPYlpneQDyThQIxaOvhZr0x/kApaWGm2Hz
TzpquveboPz4K9qilwHJl00q+yRywXW5JNeResnyPJuUF8f2jh2TC/lFis9n7OZcTB0pF5/dbu4z
62BS86qMCTVk+H78uf+x4OAOdgrCoOxAjFIwFbJH9nyVQq8tSGLfwEOWtzBZwkPRLyY+AAT84aaX
BHOAXU69iorEqph+tNtj1s/waMRLL3ouLPwlac0eftWctSWBY4axycDKpUifYWIuXUJH55byMNcF
ejER3OrxdjE42Hum3BBaPkjysdRh1/Gf3zPjr9GcWl96039c+AImRg+nytfRaOCFKD0nKXHu26yB
CPXrXL37JwVOnxdQTELHjWO5oMhEV5GS2EdEgrRfdJ24IuCNjv+eEUfdOSDwY+1gk5qfCRfYQHp1
LiutT9gHVLuLQ7BkWx66FtbssyGABbUvZNuoIXqZcZz1CF+74g9wrxEw2MmU4uojqm8a4qX4ySZO
gJhRhwwknrXxUcvmrH0eUI4cjiA/rWDdLpjRBPdXHdAqorlnwXiejX6kbd+loCqH1gOOPqg0Ubhu
hO9/d6UJgZufaLFE/sLhqbn7KpheBvuMMuZM7PW6A5bslPB5HEEj+epeP1lSk/wM6UrS7Hm7FErl
86S2dRXx0hJ34Bjh+l7wA5wFRQhnF+ZSfONVWPsmQ0hud9BuURsIxDZiE0vktgB8vLP3X6lWXwWR
s8zuDzfuky+XwZC37aYQsifYYYMPHwSLDvj6vjYIPYV/xVWC7WFn5DSl1ChJ4sbQLyLdVB/U57O3
2yJ//rdKf5U2lryqaib6MiUGB2pWQIbaiyC9jZtlTkmbHebDOjZJu99MSofrVftt75jQ86G+TrwS
nW1KoVgY2eVUod4joufNyM1VIapE+vllqzyY7MzyEdEbUlpZS7xLC8Z/nBtv+8vQjjhdXoZiKcTE
Cp5JurB3ykb/jKsGIULN/Lx2TY4RdC6ALI2djYeOoAb5DRBvpw2rB+snsQBwPaDZYPGGfQ1F3QWo
2exWKLaF0wZXFzZh+sFxEoeMttiIaFQ8gXpYFT3bY0WOVFfWU51euCmuWsPkcHFCq+iwZJ2j/8PM
fSrYT/d41Laazd2/nefeSWh8MC6x/jkv3Zi7pA25GZl5ts+ylSmH8Uv7wZK8Ug+yqyAkLwdfsLoO
YXILPGP2HvfNobqpq/xS5DF6FzIBDkx0QxdwWpzesdFUwTUQ0YlJpxLIrGBXIc1YHQhSv3V1189W
WdfdqbMOQ3o1x0dwSG6ZCgeNjeOeT8AkIwUoKf4uZvdPuBTi0L1voGuHhxg9yv4X09G69YWrQp5u
u08GvnMQmjY8SExu5BJxFfGWG1Q0udL8MFKGvux58TgdjkNrEW0kZRWMY8jb80EGTCi6bpLFqOMz
h6u1+aIXOYN0QOEBoSRo51aZOnaUTRpHjDzvQ0mCqFiZPw8fAGeitWWWO1Efqop6BLyMEq5l/H8/
t8hyc5WTSmc+1lsiDL6LWCojYwF67ip9DXGMYWDZn1u5LI5SOXolk2/AsdzTBasrm39qPjgFpM9w
0CW4FQv/hLEjyj9cF/XMA1tqY7ETa23q0xDp77uZEvd4YpHYV6N3THvvEU2+8F+fd4AhDWW8zKeB
U1sE0B3NmHnq/HGRE6UMgdcs8SzJapo7OfhToi1hNZuiRvrl6Fu2DMkREbQGr/iHqyT+7/Gjk5ai
uEecAB3GKRLFJWYmOF8w5tufDNl4VBSMaXuekBgEa2dqnLVj/OKAb6y0kNI16fJlSrtgdS8/Nbjy
L3YDfhs+m0NIuQggKzvPtRWooWcIEav1F4Gu/fZi7U0Y8KtEWe0jM9BMmtsPS+IOP5Hm7YH0Q6Wp
ceNWvqooJ9A1iAcLRtHPOPJtabtpRlHRuKJpYgLfCUegxDjlf/R+VtayU9aTCV16CPwKuH/E62Kj
a+WPinaVJ/QlYp8frflU49spMPIuW47wAHCRKAjhesCLhhPy+VO4/Pd8URpqua2jXQKX0gApOwXb
Ts0uQKnOO0n/kIe+j3hiKqvw8V/mhVq0KRMwA8YZp+LAA/A3kpeeyVRx4cfODCq4wVPmzRODjfut
AxmNvwWPsJse3AOd82Vcow9Ci7fTQUXEEoH0WeyYMGOa4TlnK0d6D6HlOYuN8jGxZSvJWv2fqcKP
Y1Gcfn5Ef70qUQmCVd3T1YiNNMEpMdGouJJXg0jd5WbBgncdSLupTtUpOTlnQCmxo6t2hdDWS7FZ
z63XjzvzJLQ/V/m37uprDP4scIQwNirHl+7DvOOlFsiZxL8hEZZvQagaeKMVsH1ais8GHFZiTGrO
QP1yWyycdb+iLV5rURYsHSVWvBfnGWPuhXO5TQ7UI12xC+DJevLy1todBhn56YLQRLReeFG2wdzT
mJe+WnvuhyjMzX84lntdU2BtDH/JwhmK0B5J41hazi3n7m6r82lMlv0Bz76SsshogQ/6Rk7aVYWW
oJ3wCCR6Tv9PZGZ0DFIWzKPlfmYmxKUG3QA1ZITNSAV9NcoY2n1CmL3Kc1adpWmcg+qD+GbNIo9L
WlQAAHWNb7cdW9vuoaDyCy2QvA1CXfm3RUN+13Px4sHWv5Adumuk9UCE2jeTqNDV1guveRttbjhS
a3ZK8wAVAmhdoxwfMGlXydBQdWLe61icJ4Iu1rbfEcakcfHxK+W0DupoLbzQ7txvIEuoU58N1qaQ
ZNbyvSXYtLrC8syJf3ZmTJ4s5g33VgRYxKMh9Hmki/g2WgI+S/n+8yT72O+puFJAWYCBkXXMydb8
RT1SmZHL7RS4qEMklFmMQV/gxkCofKdmNIa8eDKQeFwJbQrJLIT6Knzyz0VQgrd69TlE4ov9iveF
mCB5vk6hh8GNoFVKBvuMZfCQwG90iN19mqaOGEi2hG7WUPez0tNOkECBEHDBJ3uj7OfsPBx7DoNL
hrVs6FL7nWpm7vpt2/bRcS/XLCstyIzNmBpreFNhm14wOkx9386kA3p3ztkbesSjSm1efK+IgubK
aAc1En+q47iJpIwmqHR1VnPMxDlMxWdvRNpBGtnxk5I4Dj+Ur1ORkLTyQF6+GkxK1JBIXufsA8Ap
Tv03vN9J9pBBJfJqT7s3SVIjqFND7IiCHDRvbbBLiWEWD5EJkyz+Z8xESCBaTKzw43w2h0hz5Z5P
3EGQTAXKBn4noNzkhV93h1ywQgj2uecsgdeCddn6TvrK5h+MX83gkQ0T/LxGZHzh+jLhA2gglGmx
lJcbap9xvfU1cjO0HzH5WJGctRspGhZP7CjKSK+1FkI1BRZIZU01fnM21aUoBEftdEw7lJTYYVsz
Rgvkerpu8AD4WBla5rwcStaowOYliufsw0xEOJ4HVo1sgpEx5fRkKHDYzEklh16p4n7yxdZxPhEz
Dcp/NQM/g5ppSHvpgJWzrqRH/MNDCilnvoN0X8aDY9Q7Y2sZ1t9w7974329Bqn3F8PnK7EVIwrue
YIstBz36inffu/XlcNzgOSVb/bMIh9HTCUDn+8/wq51I7zq1SeYieTQ2L2yJWZiFgWKFzKXOpCZc
ShJEgWK9CRCvyhdVY+aOYI8MEZIiCxKVXq4RIQuoEo3v7Zu4nfaMtRfkBeW9OIia06qOAVRoU29J
5FtkFaeg5RtHv9usLggZtCHA9ix2zNzkU5jaqIOwZkjBeZzaT7q2gcEyk2YyMJ8vxPl32tG9WGad
6Mhh6TCS7rMLb/nkimLOeMy3zMDZ0eJNZmW6T44waefKOuyQbiSb4C7kBW17U3wAZGC9Z5F2HiqA
xjnBB5WA9qQYjSlQ2FmLCD/pCMzN26L3fGEpFThXSjRNqkVOuTkJuKwdOZiGvoQ+7rozKXpg7LaM
xVP8X3UjV2kxWCA5KdDrjY8BsOyyoPb3bNPng7jeEgobEI1nXsVQw/QwKHf3VSs8SqJYZ1Pb8joE
/s03kiuhQBBLYmdMH145MLsbNB1hbTScSN6fqRmry7jnVr3bWm4goUeFGBl5j7dT1t5zcfwOdzrs
jJuFxyqqo6tumdRSmbr8Tm5lNQe22/NuE7It4zyFMyauUL661YxgcVcOtM8jJNyvYDr7QIcl9a8D
+NIKPU8qGabS9nX1gUAhR5wlvIHtOLHJ559jKrXt4kz3nIfFM+/h/9/KXQsUFyspd+rQIFlCBcuJ
+6nw5tbRbSPVrMhu4Qr176lsQW4YVjUlx36kcNT4X4ZiOtv1taUi0l467Dy8guMV/iZMIESuT6mP
BecEO/ZEcO5XkvLsKdfgRrj6ws57zUVD5OXdLOHt6ewh8wcSeyXmHmYw7taH8mYKtRi7G79fDSgN
J0e9OJNND4rQsmp4K71nuGwlRGR3jkbc6WbigMJI/lM/fUZoH6AebTa60vZGQTdUFetR83RhyhB5
mZiU/a+RBeCDfl1C3nsty2/cw3ZALA4Oz/G2LxwYksdigWUwhjivkIbmuufoCc96lI1Wbs6CX+FN
BoYNB4+kmZb+0n2lBOwcg0fkJjlQH+jpy/m5JVRRxJAYZL+1Q8xKOrOc3vhQKGuASg65WPpvW8qx
LqrlJXfR643SmrxxKewBwupWOOvLTIHYsi9B6kYllbNGRUbU/fu0uBBlEMR6Xx1TB+tFCnq7t5gG
Nt87J3s9MOIRsJFxo0+Jf3aaVlzbTQFjJ4KVgApRyVNZKSVATlseQNFSM8NbWvNgp5szTpQWCo7m
/KL4PpqM2Ejg2wJs8F8g2NfrMeLfm9aX8JJ/O+ZuK8Q51Zuo5lihjuzCmun+BJX0P6enlTw7eZPV
ajbYkaT0fnpjhLMs1KqZ2F8iQjII/Ix+NN15+5/mkmY8wQyveMibs4796nmjQ3jNYKtSifecka7t
fvj90TFsiCHipNH0fS4r/GTUFmMAvhilhu0/O+364zaTLkMbFTnKmWks+8bU6BXxpUfPqz60F6kI
u4kVNgR54KgJR3if/ySLyVL5PVZvYiP/ePkXSosDzmu2UYOcyfntygkKDzHkr0OORlFxMjEjM6h5
UgOBsdEXSMP1JNcC4un4fm2wonTKPilWjxQ/m+f+1RhJPP271d9eSki4SJrNRDZbMKpt7sJdmSQt
c13YPfL4PO1GPqUIkMZ2gpACuwIDEfvVHzAkal4me8BO1Rv72Fkzf5WbArdSzd/lmZlbe7z7dQ6F
1OvWwqNXD/gmX5cm7MTP8AVMOmDzYjfhJ8JJzn5YDxtjHkwm+1vWv/FZvMXUc5+vI3/nrH1un0tI
qPxu0DvEN6dnPTBy+DodXQPnCz2WcCYDXi3Jc2oTrZcY7F6sh2EaAk1h9IrDhuesxINaTmGycTiM
pIEL7aGoDu856mPAsBoii/XpEUQwh3JngESwXXG9L/2LjMFaeAWfW/+lnGPnJ6+d3RTlgLQWwnJp
1HvLhz6VqFuyjKpxo2Dw43TVLRb6nzFan/MRdy9GwRAjZeF92zr6N6Xp8onu2VwSoWSg60Xzniht
kkMi+vNBlPT145JQCfwZrd0qir6Vpa2rF/sFdDSjS5YYUkbOe2+25EuTAgNNYZUtw0ldNZmSiUVw
sR2x/Daxt28HixKhZr/rA+82zAcqSVMVn6c4wOmL0dOphQYyXrCK8TapmKrikvgzV1ofmaH2heCk
Ft0g9QkeEErzbFy/zEgkCkVUWLr1xuFl0BI2CZgBPo0jvrstLE0Y+0WG/+U19yvLg17V05cYsOa5
K3uX6HyHsuTnTCWolE++nQ0b0YGUnPNGkJ0wRIZwoSsgIiWHJ/eOlmJz10/S36fnPJKaAHQHt7KT
YGth8NfOERT44P4o3As2SMY9hjs53Z27lquKRzF0CBpFENI9K2yAmUqTPrIc7BX7qBgeHNR7ppwb
ENv8JZkhLfNGtZ+ymuDUB3n3Fpv3ntRt6D5rG8ROjFPApx1aFOICMDc8ZphotOqKv1BKCeMWN3BL
4W3OQMh+4Ui3OsQjTd27cRdzwZ38WdV0DYCkeTvkGEACGCHQn9orEbFfexcPN8HOvpYP/GbWXsUp
HrX5ICHisllPgrVxVTx4EaYyzzSVAwOIXsg2j9a9GoCnCmMf7enX09qguo/59y/iENvB2wGOtYaU
emhUCzWa0+nliCtyt5ya0kD+QPrcKSPzVFXxHnEXiNQf/WBZq5Pi2O0npIwRR9BRokJXM/an9iTs
Wevh7l/rNg3yxA5xltymNA1s0Vuua5S9mJ3FIOfbnTbAVKuDrsjHzZUc7sP2EHDhRCHMcs3SDjTn
AfvJ27IJA2p7w2NVDWdswuZ/MmaOGPM+/m7G/5+MWAfNVyzbdiU0ymuMvYoVVT1qDiK5dUpUPAm7
qGshXRwFkD2pJ/EUa26mboQ0Smds9WY849Nyhi6LDAmO3kWgPxgZX2q51gx/mK9NKWrZrSQi0neC
LT1Dn3A33o1RW1qeya86VZWU2XImccWOKzI+itA6WrdVrHSv50UdH/bxa5pwyScqq9nrkxNfwg+a
uak+nt6+XeayxcM10wQPKbBAYXipSDEFVU0Ih656FcfpevdloukYZXUFL6JhX5obgMjGzqFt7xRz
6IIRzn0rOX3cQTPsHQYdy+e00YJhT9Pmp+88B9s7VyplKgPHrbI7tS3rKz+sOFe8Gzv2iItXm7/c
FjzeNcYXD+bJIO6C01Tv1FCeYxVsS+lpgzBlytLLdhsUd5EcQr3Qgd/D0dFc9UObaUI0G6zKjDY9
29lzojzFwVbkQ6e+LDboIoay8rnm5GGkI4ZM30G5vjGXTXWuWyOIwFk1mj2XDqiwGwxcxCx8PM4+
Bl+31Xz1xLg2rO41EhvnZoLNMfQs4y9CJjpJGWb9Yk6j8QL+Mrb+sTtKkm6+A8/Bx9wMgoDtvfXD
pmOACInsgwjxsoDhQf3P6jsu6XHet/YX5JyE7BmDmIa4EgIB8NMo9gHOyX/PDBjkwp3JZ8s7Xzrr
xi6z99+H0TETV3fJdRlHvw1l96gSCFTQpXlPRz2pw/8dZnhES6JwyiqPLJuz11ltcr2oMVdDKoIY
PGV4SWF92mx45Wp253agScu69mGnnuYIn1aFwSE78Nsr16Gs2d0GtEPblvQhOec4mrYGBePw8Jmc
U7U9khL+/nDhNgvRAPG/ZQ2aFEQ51BQ/jwuY5jIgmRTQ/bz3YvvXC4KSS8VJ652bI4B0PHoe6WO4
EqdF5H38UHRGl6B+vjsDArum26wPN7MXENlBekU9dC4gsIDx+fl9hgDCXwc6q75Gvb7u6UNOVNS/
HVbffL20T6KQkM93+MNUd0rWxEOY/eufW/iDnhwoV7/VXy4oFUEd5XaCIX1nXlLQzICiCQExm+NA
iTTkNUO5u2EG5IjZoSSllAfvKFRLruyr9T0fjuvE/4RHCJG+zuOqmK4qBCGM5xMLlbn4CuGnTJ3C
chb40O1MYJ5qf24HOIr74MnaIIA85HV7yVBiGni9jWR4hJ2yaAG2211TBjkl95wVwnrDEr94riEC
OsHVmkQCUmIubLzLXywJIV0+KkECRILcw1P2flQb9ZttBhzTNLtyijT4s/0rs750ltjH0yxRh1At
wCrYn3DJ6ajfu/v1br+bLtIK3ZmpcOiK9UvCD2EC56ZKNTAPvfphemT6E9w/gSOmVX1M70mprckJ
/DcaM/h2mZdSHt6ffC2XWZ/kyDI+SrrAkjBag5/My1wY/6rx0bKh8w9N4Ygptc6XTKfVt5TAlDMh
7KZMf2P6d1DUayLsVAUKCT5yDJ4qbrZE4V5w6vIlQQfcpK6zjf8SFR+nsRFoQKGOWTP+o5+NCKOs
i/E7CCS7ukV3vmFKaKpbxN8pFFUFFziMzevjmzXMNRIVizhikXGjaSTYdM5CE1X9VAXsirBZgxio
szezgClvwK10tkgOUqDUblHQu9nIPIkW7Aj9EyLsMb6YM1TdHrUMD6DGRrW6YiUchm9PpY2M3zeE
hPZUcIu/5ka5bpy/IjX00juyLLf4FiYeU7mAVKX0tVDM0OEKVXMIxf2uSbkqz2MnMBe1bkT2HeIk
RLkjd0+tAS1WArZyiuzo1NPZwxgEGqMZr/Dv2y97LO88Fqq9TdGJlytVbnk6i8JDz3h3Nd1zxpVA
gqpyPq+EkcQOpdPjfB7EGfCHn5pg95JINB26IUEOunU/k28jErs81jf1GRtUEWMbfF0s0VRyi80C
JE6qOA8Io1dc0XdwZfZYJ6ReGrd128gtmWHUITeZmEFcqci60677OoX9aB7+5T+IL0WHN1shkxE9
L/BxMBg4/DeeymqFE1UQlHx3r+k6Rw253lHUPSGLvf0NW99Eg4EfqagpoAS/27SAn+inEk8Sovm7
DAlHeKyLEtx4U3Yn17OmFU7pYi+lco0hPCC0XEutkFThB1m2R9x9tp8QoBLQJymgWNtnvLms3Q0C
2JBtmNAWo5vhbI7QWhcpMIGI2Tt7qx011FWlse4P8xTqxenzt7tZCipmHjST1Pmj0RDVf0PQAj+P
njiQnmY63tP8EsNP285NFE1yyw/29vFJ3F1k//htN/2X2r/yfiUkv7f7EG+CNKLVVe+w0HH7QiQy
bmEiI1TLDJnc5Cw+aTIGZwQkMsEZ1aEhRKUkSCjAxh721odBES5dNS/ZCT5FNM4ldLyC1kFuD/Ne
Qh0K5JBe5cmCmldXT/nSYuf134PCxnbQxnPFG6vtQ3W9AAdDo0HHI3s/csoC6c8mNohsXiAKXcjQ
T5K3xexDL7l/04PiruB8y9nZB5i/wNkHjZVICY0JBQgRUiQJtx3PPuBHdoDB39xveFAcgquJSiaI
SOAurWF6pnm+9O3KjJc02auRRyJK5hKft/GmHYFw/SHdJuIf2X1OkxSNHsc1rmmFePVzXh77cOlT
yHzbUfm/uxBBXgvdkg3+oL/pLqTGNDr2c+PnAicerZ1UJHSbMC7V6/VEwSBevjlQqTTkSWjPPAQE
HcMLxa+lr5HnvDxQNz9IpQVusFIkjm1cnYamOZc0O00I2/4Ta0uPnZzohcEm7w1tkXVkXZMB2afJ
hbALFePvnqqL8QBdGWqm0NHmuFpQxOa23sNkZ7AuCrbFCPTGtZFqq677NV7YP0K2VytRhACoRZW7
2qYkqXZD2qB6Uq03g/h3aIAFbJqlbH9Dl+ryNvfbjgOT/YYR0JCfhdjzg+K8a0SILZkJ0iPPte8U
y8xfeb7M9dtQyzjhYf05Nvd585AuDCVa48hUFKFv1LnNci2NQ0YCtsPcF66pq0rzELryWCffkdYa
pmlCgW7sqp264FnmwdLcWXH2NgLbR4EwGb+SWyfAIKkhNF2U9Zf/W3iNaRDmwyejM+FO0bY6p4Vg
9ZwQ7nJ96sdukXUb1MGObC6GJ/TWhSBRolrzmQB1T/vDoOtk0iZQ3lavJ6Hi+ua0AkCDTaCVOGne
TAgbth1/avnMsAhWAIiNn/wB4sOUwEr3TfnyvXscJFwdBOxlsFzoOYYRpUiozccYfoIRbRJ2f3s5
smvBQSz7MQMz1m7Y5OTnZpbdzVt5NTBjMx+dV9K1MCQWoo6Y55CMWr15HBliNdNtNZtGMYu5d0zq
44lp6sUGtb8JrvSuIQyQ43ushkquWxBoDyCbi4XgmA1sfI+mBkhnIXGfBcNXyzwGIRUse4ovW1DZ
xmGReN42eHaajBZXK9T/V6AeUjfB/vmnksDa305QXogc2HliRy+WBShzylRsbYtdPlyZ8oxeZDfx
EA/GaQDWFHDNtoKGwTAzL5togI9IDofThuT65zOjCQKAbAWJE40Z1PhGb7WRLMVaf+XBEIKohRz/
ejgU52eMTu7WcyQzP+cxC7DMhDbu3SXZF7tG4uxZkCprwpPTrDvZaPvmrP9ZLklIE5jyNpT9IBsp
G8MuQgOi+EubE7GAb4GVZqXJvdWENCF9sINNtDKs2y3dxfIuhT1Ttfo/SNJR5fBUW/SXr9T4Jrkp
2GqKK5ZABzjGJNFHhXCxa1UVwW6IeCJzkf6/zthkLBiDvYsM9ZnDnZifQ2KJsc/+f3NiBQcCVZZi
2eld30L+5w76a6kU4QQq0mvcY4EiO/rVMl+XoYizyngF77kJAxAv/cAj03+WJbOtOblxZlWS4ZsP
H6qqO+R+lYYKMD5TpK8QQeBicBQpxG/lJqNnOiP8FmPCe/14hyWpEg6ezYFtoFVCJNxjf8FmRJgG
dn16Ljx0ivoMV0veJbecck3vGqcqj7EsvPqUk0DmtRNP4CJn3xEDeF4RO/zv/y47/C2e9Y86LmRZ
2kM+luTroEmRLONbCbn9DVPdajBFenLMSJdfBTJqQUSNzi+R2r7KwZklFNNGRHI4NiwcGA2T5gdP
pAq4v+gtHOnCV2Ia9YlPDZ7rIoTXr/PyfvTCGaNGQAkgqpiewtmUyxgSjhGisGIEK7QcBY2oSEj8
P7qGx15HpzzZHkYTZ3llzux2OL+WP4HeMas9MjVPh8wk1cgH7pOcXXCPdOfB+us7CYqKf8xUnbpM
8QScsmP8AY2AhNKy9SVFaODinG1tATBQ0S+3dhSHWGU5dP6m1o8RMGRZA6U9g1RSE49I6wG0vmcS
29FcyZ20rN53RsUZRgVXZM+xHVjpsPrGStrXiuFHKL5LzWc1d8wJkNEgbgJ6iBrb43brRIDRrzut
nrOUVYX8ITxY1KD+BO8St9u2Nx7GWOceHie+snGZvAIvMenbAVG55JYujfreXYLKA2q5iV1saWR2
mosrf6qO22bSKcxwvW/V6tXixXHF2uov8lTREQzbU7LcFMblGQAjZER0Yo+tHCnMVG6WB/CSYjaL
YVeWF9eBacFddpYWKdvg/Bp3HOualNY3Njk61uAeWzVAE5ltzhEr9sUBzgWvkEi68d69sWlGi9j4
/TLNzJwDq/jafoIh5rdDBXDHj98miKzgqmrW+/GBKdxPA22UgiYvMT15olYWRGeFBPBATgPbeU/G
dryk+02B2mLANZ0mUthE/q0E0I1ODvkkJDSiqIzGfPo1SdsRASm9mUt+G2i9nRTWjvuNlvFSpAVl
g8OqgJ/QR9tnyeEA3g9ZOy1CnQlmC5VtH/5tp9W2pUvATaHEQNK3IQPnQf1FS9JsC0vIEHwMTdeh
cw/3g0r2oJBdOOYTZh7lV7Cggu4w/51LmwlZCRaC6tFxTVrbl90q1/E3K6JMttzNLDpELjiGpYtb
OGMtr1SFIA6fO813QZKSAv+vWfjKt5ZMLxY/V8B0odl9IkiyMh4X6yq5svaROV45f/uTPlNKklMQ
vVPnD0sRwXXHH6O/aleJDxMQvZOqsXU+JVwb/mLD8LRIjOM/7/JgNJSdUVS00cYou2i1uIyWO5F3
I+w0s70xNMpFeI47v3OEpVD0cESeYmRNA/eHPipplIHCC5RYPMcTrfCuViJCYkWmDwjfLY3PDlSq
vYfWLmrmZ0iLYYOxcoPVTAszfGWRwsonLrxq/U3lIwxb5MFL/nQ2Zafn2xvP0mJVGAUjXpb+KDHx
C6P6j8hUsgEtSvgr3eVGxAsPk71wmd4pK1msUO8iNdk6jRB9PTLuHGttY64LuKB4yG90On1TsMA5
Ec0DVm8dWADSKfS2lCN5hYTuxS/NUCcP5zC8gglb4vUaBb8oBoCzi3OeTUY5EkbQHNFpbFI+1u6s
EC7lbKH04d8yf+WLNd3CBFAlXohzMLuER06krA+rVOzLMGueQS683NXwwtFQuTuAuyoBB4pobGt3
S2LSteOCFC/1rtQzGxRe+tNbDIQLe3lWOyhk78gq7gjGdmz5hEf6PvwC7XxfANl5L1hyogWwe1/3
yCnKHHYyNwwp75kJC0gFNSAfzN4qKdBiIsuWX99yXTZFJ0aDmCn08tbWK73wXknQUIZAyfDZcmbi
14dByKwkvtaRryCYK5LbUjA8wEmvXum5tIyFe98iqctiI/ISh2p6Id66uyGTPeqk2v49aVGNdpRx
ztAnP56E0fqcvHPPMWxrUyC0K9zMI3fp+DViZ/Va869xtLnAObryMNR9tL/DzRJD4PP/BIwZqk87
EL2EciWKjAmJRXYTvcCjtFjzcMo4MsRDau8pCttScC2RltaZ788TtltRAkOBUvoyDMoIPRUAiWh+
CwptiRigQ0+uIKKLaHdrj69EH4ZxCYSGjF6dk1oJrO63ASjfVYVuS07FhOjpsSnGn7vcRJMQWWPv
uVflRRVumUzVFyCd+k+u0YhycmIjCXYDyIrPq4c2am86RhXpsEyuofelBpxMEwl4LSGkwsaMePoA
4M7F+Gvw3uQdJBUwcmMhMmZWhVRVij+PIHfeZ0Se2pnGiCx9ii011MT8c0vAM3dUdFpA5lj2O6Mq
qXW1SXc+Q4siCz7Zya5cjpCMfriyezHSFNQ7XZlfx9fTizu2Bo/KZzpU5nu0duGTITdCss1p79bS
jBNWqHnS+7yqbvqtKafaYEvIEPOxeltPn/UvxBIQq6mAqsZ59/o5eckDTeLwZGb0NtyVrOFtDH/0
aIRtXOYadEIgQVHi8nKdjHShqViLKwdlSQbtHntCOb14Jdydd+8Z92iMYgh42uX/wzT+QP7VnDGo
PEysVNykrIVsI3H7BBA52/3RaKAPjE/VoCod0fJXb5i9K61o+H1UbOTKhIbcyIdBUqvCaZaXisAh
QY8h5+ZNwQA1f3z8GE8bVgK7MI2+2IBL7+oOKMmxWF3fkfzihbc2Pi240GBfXsPU0W9vBhORFG5+
PHwn47+HRkKfvw70DUFPD+VT3zd3qFoWpyoJJemLsOcA2Dd+uA+5lr4qe82T+glF7H77IHT4S0zJ
Ha0dQlDgmfrYoeGRD9kugHB8lF4SGnbnkqB0quSHiv5kUjTsx5yT2Yyw4zEED29qbtT6fN585KjH
N6uYuta6t1ozv3Jl0b+NHsakuyEppYca5+ZOGZXEnyiSxPvd+MT8FaYjLjHrfCV44zro+C+H0VF+
o/jnxnAwQA/x6F77tpB+Vd0p+eLSDVv4Lrb0v9yFxnjp8KsqYN2MKP+GsCyjJpRX5fZ8UPKWGZmZ
Fik23J9A8ccrvY1sraEdL8VlkZTVc7ijnjtgF6Q00joxKBzVTA6QzO+nFUxi/M2RuI3pYbMTE7Nn
K0JvzKTWHWk73HH4dE4GroW/6LlSILomw2IyOELky5b53oab2PfiWm9rh+MOP1Zt8hZpNT0sa5wY
Mkl6FKEJTKg/W+N54zqePfhTkSa0MKlnTgaxqIuYfCy967EJUVwb9nwBxZTsZjWFS02Alj1mCCjk
4MRxZFtbGW7ugUUoGvx5H+9T0YP8EtwG94DrUEgNnKy6T+g+HQzzsGmU/V0iN7CEnt3DfrE+YFEZ
SzKx3G31kj3fUUkF5vE7Q+P9Q8q20BeGre10ufuNAJzo1lHgEmkEWpoUBlF9Z7LerkrTMYwPPVE+
bb+h0IXD+LVxPWQm89VCiTzYUOpwpV17f21C5EGgOTRtPnFxP/0uXXVKJg9UDvNy0IZulmw4U9AV
gtoMbka1BE/6gvp1vCW7ncIEPmg8+NzfpCEpPkBlK2P/BScX3n+Ong3u5yzFqRHkH65qIFYCCwQy
Ac20hbpCu4D7DKmq3l9wrR0d+4/M/cprGtHOVKoNDRgcfLSa0FddzeJGOgZstCaZ/+DPXXuMsTJ8
/NHSf1zXYk3UjMC9u1prRpOmIxm7yGzSGQThVoqrfhqIdt7t3Kt19hwAp1pFdt/MuXjipOKa7aXb
uUmijFzEnktwwZnZl5gk8PZmK4dtXLA2v5UG356MU9A4vhvXeXmuN1LmukL2OzOlwQ/HZC3++AUO
gxToz5FyRYIyTTcbuUheVq6LGmVs94As/1/PknkffmVFAVStcA77SjHSjNZBZRtpBbGy7L8io93K
GroxuymdhYnSS/hkZYE5j/kJhUvkzqshr3mNmA84YhPFOLxC4fsORHeFLER1uoj9d8sSA1Tft7MM
6IWrQS7viCFHgdUrXC8ooyWZx4qeXYoKfPnmErt8Lv4Pvb1JSXPZaeeKyYCs7227a4LewdeJrgTH
bHuSENz62+ugkjH40UXDIFJQ+WLOe6yjgGnERwrP2ogKotenOVKzH4AuIcnFiQIIJEmfGEXrINpr
RZ9zO8bhkQo7lvvtnCqtlRLLo1E9A/w+0aO/AwV0gYNIwqJpkojSAth6y4XnGCCoZXikqkcYuJHT
JyLMY7188RqGjT3GbvUWveHHw0cjbVcH4jVR2wTlfhInu+cMtgfZLdlqyNoABRrbVk/AldA6w5gr
rnOPZvkwRe2fxrKzCv04bVHt/C2SDExIT2W9zoe19lH7ITDxHcMClXOELiaHjZXk3IV0+fnPby3t
AkBwvabt6z2Dd6bc2Ci33Xp7lKsIqpNnQuNofMQxo41tvnHOczvrwsBiL5SOSOT4lu636JVX1v/e
bL2YBAd+xCQNbu81LmjWCNEMPnIwSLjoLG1vF9ye90x5oxwXt9sm12PrML3Mla5mK3omf7a+QswR
LkgV/dr1FoJclwh1sLRPRJDAw4mYlezK8mnuEZ9/BoI0WUiqjWz2deyiv50irQLc7GuCFi25UGf6
lawkWNglay2OmBItbykqxHARXWItluz4LoY/pcd+sAPLVBxLG1iklBSjaeMnPCO1u2z6RDt43krn
UiZzvy5Wy0/KKB0fPvXnO9ITM7IhbBENiUC/C3Z8/XyO8Xg4lnoc2Fbh08voXl9MQqT8WuY+s6Qq
YE6DhsfJi7wFcGP4nRqpCKIR1ObzoRutI8Lo/8wlVG1l1PENXz6hOmUc8nTIQkfjen/z6b5NWJwc
6zMsXznWUA4DPZ20dtNzCnfhDE9yErZaH82MnAAiViOQK9Us5HyGahyBt/Wc2TnSa+t4fH4E9EkI
AycygXZ5KCoYREHwfpNudhX/w3thAR7liQpVY0XOA2YGx+CFMtgkj/Iev2Wr+TIMfc+Go7xtCmS3
Qv4gzjYv4KE2ekP/yTFt4u5O2qnHFab672Ic3toAhZq9NBiuCSx4jHm0uvG31F7ldr1PXmQlAoBX
LdGt+fu7Vos9R5F4l7l7yiaNunC6ybwAN1w5KIJ+ek21Ce3xdg8fYmWmkx2HC9V1GQZNnBl0qs+/
kaTM5fEK5v4YZIdSER9/jsLVPUqU3wP9OgLXUWrCHo8OQjluP+Y02RxqwWBkPvs6vg5Xku/kJWOj
hV0wKUK0wG3WQEIDh6ILBy00KsfQtlAWzxiRGnILnG0JLUeRFrxXX7uibamOoJ7clXWkUrklvTiT
rj7IEfWk1HYS5CMwJI96+YqdHKfwHhb5RvMtkH9cNJUypNYZLVRWcyGgF6DEuigM5ROGhSGe2Iis
rgAJ+J2rnVwdOfYHOo08PE84tpRO2UQR/e+ni2F5bzrTt2RJ0rTDVyFhkbc/SHGJh1DKfl6mYj0U
wNpyMtEt73lV2HCUu6o1+hkzJXY8Ix+tBbZcCag0v19milklh4guf0k2odscwpu88VhWSFTWBobe
rdpuR7TH0XvxWn+ipht+xbPPSKCp/5Em6NyBBZbETmz3mfHSHNxlsL7Yb/2g0AY7/O71WJEhCjtw
TkG8cj2Mo1kiz8VqpAlUbBkt62OriEd/rbg4XnWxmz1MJ/yPCG9gl/yaofHexDwHY1gY3OSunpQ/
BFaPtveOT9p7TGR0e/S7JIn6aKzmyWJ/BlH8MNor+jzUJFZYqGDRHz72Q19Y6Dk0EXNCdXotdJgI
mB2zqtgyowhIQhrl7gsoFj8c2Vxq9j3FzlZ5IMJOjCfsVDh9FgvH70mZ539t6aAej3tehhezhFGl
sSvlBvdyo2LmYlDXkcUXwr1CJaRj5CyVqfx97BqIMZZyITZbsJHGJK8HUKv+yTOjrJBypFCL4DF7
j0980oH5BQlwa+urjsRN8wwYBqT4JRqZrHHQT8T/prLBOwTYoBPgqf7hygMcshGiPqRW6ai0iHLB
tiq0+W5+3+Mqdve5eyo8mvj4ZfSxAmtTm3qYayu5jBFgXXqDjKBRXqdl03CYGZX4iK3IeAhRcZV+
1Piqx89TciirxDSpV0kZJOXH3gsJy5OmmI50b2RPiAlY15MS8FS7b6LRvqbVTMFOtF19I2snTovp
llyieoID3ae1eFHt9YkR6fb5MLnkNQDvj11/vd0STVTy7Ev+CEGwZHkRpMWjtVkE9f+etN2lNR0o
3KKHL6WLw/BD+LXkIYXnlmNEZ6TL+ObmpPL6W9DjgnmjhhvpNs9T0LJOitb9F7n9R6kcj1xCwgqh
YlmjhuQMlT47NnIzksmXN3O4zSp/53zQK7TGGVVLhKmJ7eE0G2miDMd/CQJL12qoJPYwV8Xdd+2o
3xeZkvwh8BthLMaErnmEqTf5VmIwKqhCj9mnUmnpdvnb8d3pSSXgBVWbXNsi8rJkkatalPC9GZRg
iagvtP64GksEZE1rosnPArwvM+5PVfeWDzXf0daKvJIzdqRpTEJYYaiZoiiGchGaZbc8+CtE4kEC
tCcaEp231hNsMN83T2XvW3I40+AIUHkrR2VmP94PAKP3yLDELPwXNyGznN12EfJnLzull10p0sdV
12NWOoQG+kyCxoolsyBjBu8eJNuqhCIgk0zHNjH3J8kC2pS/w5Gh8/ryAubE/xqdRMw4Rq4dONxN
zt7DeEx7xT3y9B4AjXhuEg88yD1shy7x34TyjUrE7iDjLsbX5S8IYFEsH6opAS+VgadGr0XqqZ0a
dWnKQnokbMRtbjc80bFq+nRI8MtcgPWuegUUlyAD9OsJtpjWw5tD7Kj4KopBxslnrxg9fSopMTSv
dxGar9eLkAjbciJ4sgjBAmAYDl9aZLVIQOKMhMTZWxtAP6F0xQ1ln6c7lZgkVSkJuKS8YkJJUZTX
FO8M69Xiv2CWJDQkpONxjXhVPzNVKsIswFhJM+r7iiuf6kiL1rrhISTMqEFd7XdYAxKqWzbhD/+x
CMiduHOj93NPqXuNAbd43Grld+0lK4TOAp0mEZ8buzlNWX+76avxCF1E0dohbKZhl3WFXRRUlbF/
o2WXDiRY8atkmAG2f0byFcU/IZuBFDKskP78AM5882FrLlu2U9U9mUnGgtmHuQV41CAx/6lL+vnv
PCVLV2MxdrVjmwe4ZBxBOAxsMBSTjnRk/4A8LaupamaSGX5MdgYCYTGJzclj/SvnZ0ewfgYZ5Glr
rzOvTR4LC78RD2HxANWqhSMSDTAeb3p+/77DaPsfLuDwEGoTML6Ca+5L62Ma7vmPbb/wuZS3zjgH
HNme2jjgGiqMEFx9Vg2WJOAhQp05rAf5P8Ha33QD+yuqiz4Ac8KrU9EeOl+ra5013rvRyE6tYFvx
pIJysPUDDDZm0cl318mRQdjiRwa9C/jd9Cs0l9PutKcrtfhVRGd06l2KPBidOdgwLTNWTt7oXxip
4XRU4VqM70y72wrtfzIfxKPsqIYtsDNBurMsYqrd7uIL1JkOwCqv70YjGDFS8XXCTBVVW9nz9Jk7
0EU8qCpS2P8xTjdH5QBmn98TGKd5LaSwYebeneNIRh0m3Qzm0uOi38Wn6n8Fd+tYrkQrqJsPFb4h
hR55hIAJro6r/DryBIVwOPrjFTzG5kg2utsEvL16VQ42g2rexYXdS/uuipUpb+KUZ8wuEorrCrC7
TGEPkQxqwT8NT1BvJta8Mc/1PqOvXlTsSesVRE4AiZY4S4K/ATAwpxDL0L46gQqMTvJFg8ciWlY/
1a29I0zA6P6VSXztvaLZCjReQvz9T46iBXBqbiv76c0Rec8Y2Sdk3eZjG9dO86K20FgxCLvA5Xxo
GqA0d8RBrPqvPrM9qdITtS/y2My70oFl0b5WVNcPMwUXQfu79JEk0aGdRtkqDBUy1/jq5pgG84RH
rpIv1PVa8BJ3zTWjAp13AiwzJQ5lLK8twlHiS0yNULQ9+Bz+nHBoMGp/cB+388UIu3BTMMVYbdc+
71pZdxwoqG1vxA0fjOTKE3NIB9E+Pdq7C+N4Wy603lQSKa4ZvTVhEux6K0KCT2ePrn4jpe9mEa9N
oAht57rBX+3LCV7DxcVmYwzrZk4Wk9oZg9TY0rVdcncVPyBIRwXFPokt34MQeLh8XuIYOkA+L4Yi
LdqxTuJr8cLgH3LfT9M1+t4KBHWwLaLuvP1vkZaYQIa9hA2rXjqSte1KPW3W+JRRkT0DjWD16hXt
2y7/GtQC0f15inlC4PmF9OaaAQuPjG+4Ox9OUWeTprzMRwvVNf7hUBazluLNKFm/+mRKRpWH74yV
2PgEybhHGAAyGP54lPRuJz7WhS3jrrsBJp/1y3Y5oKKy9e2TNikXx7Piyw7Iiovi8PgTWxdP5rnO
BOn5/yQH6FJ6o7VtbGF4mX69HmYDLpJaULvPckR1L0v0PYifVry4jla94BEQEfnN2JTT0udfRtJu
HrPtgucH4MJ3ZJi+6ustLG7RwzFn9vW80k9jEAfBYE788tdZsd4xUAQVtoWAtgDEPRhZwt5Rajst
whMbZaxNHigZZNWvNUTyJTabZzPaJyMEnAtFR5qBuCUbc7UL0rxTW/ZOSdYZu7qAUuR+T0mrxpxs
Pp76YgmjLUNYeMI5BWhzZTfBiD7mX7maox6oL5d6b+ZGdvUb5EFFW6IGA0LOXDvdS2atvEuhfYwu
G7fzDRjOEoARaiBIYuQa9ToPI8EBI5z8pYQrOCW6uaDexhCGG0rh16dBZRbSp7WD/CcdDKWBBJqv
6yIqajQCE/7w6soZjz0NzDc6/ZdWwZsg0iBjfei0TR0kvtamcvJWg3Itoj0Ch7jpzDB4G3Tp3OeK
s48dINuGfqJF5imCTdCz90xNdk0+zdqaGge3iiLxGhbdKaUqvxBeAcIgM39JisJwrZ8lYccQTDnc
1VQ/8a8dBadbdpUxjzfMGz4YZOdiHHT+hgm2pwLimvWqfdrWl2fLTZaV7TaVLt3xhv2hjkJ93Qrq
F+eo6z8rWUDSJ4c/05f0FenVPfxw7S9LmfCt0JHvrWxWgTJAe9WGUVrfqL7Esp6qY979V5jB3Vjw
ZM2K6I97kSM3JWEbpluk0ultRY1PqOwX+Jj34DdGh1Bj+QUWgn3i7SlOLpSMM60bEUQwQFCaYq1S
4Ukt4HIDfGVRz5OvGKvbn+UyEsuXQ009PjlKTvNZxutUfaOiUdQfWMKkUInXZ1thcWt5gAY2BQ8M
YnCO7goBUYdU4JUXbsRbTfh0M9254zeumXslKmFPwPcvJwdofd9Cak/Heboo42hju9HG1io+3grT
dinvz8EPYAOpWHKsE7SZXpbEIoy+Z216IWAHGcU80MB7eCLe1JBtRquSiAJ2X6THU7k3CfclX28a
ofEclAnKWlzBWAQasJy8NCZiAFq6pLl7m32tqayWuGi5qBzKAQedkczioI+5Gdgvcto6YHRCrzp9
KwK7ryhUaffcs7VwzQ8kbBRiAGV7GK2j5nco5CX4eg1Esdr1PUFi32e92BEU7ZF61c7g8LPYlUJH
m5/Z3IlsBiHeHy9sitO9XY/qPelHcMsTtVtYByBrca+mM/zEuyopwQ5Qe/4vn5sMHpntdaumtNH/
n9u4GI3DVSTEN6t6zQCZyJzkKfjxb0MHaWlDNO/sEJhleLQPNQjM1ZjCOhpcu/b4PO1GjvP2IXuK
lwE3TB0ShrYFP+avZ8EDZ1qLkAEsw+bl79errM3a+pvBSBnKkExItAGj3SByjg9AHRhEuUBPq+LT
wBOiqZuraOG1aw81jkkErFZdUc6fT9AVP6uuVdrCpficp/deew5ueMsDJHk2aOCEL/dhzb3uB6U/
o+i41HKQH9z+ES+7l3FbDutEazHlCJNT5PbTM8bfGIF7XkbKj1ptJEKTppP7wEUNTMAgYsi+KDqM
xkgI8cx3xGRVEcyV0qokHKkRzrn692SgKyU6JaO4rV2xTnPsaKNDZwFTEYSi0RfckM5G2v7n65JU
Z7hGn+EOUoTvUQh35ey8nCY1TmzeU3/e3i7Y10Qht8mVZQBo96ombgQxQ4TsCMSzl3o/qWxM1wq7
AVaTQyKx67D1QXzCjG3AJqaj4avAXuv+MOLobX0KMwMkQPxpBTCyTdrvrNktaSI+Q02NxGsoHcCy
70Egk6I1EpTn4bmW2xydbSlKjBRbihLVAhYyP4VjI9wb5hE2uRMCjPhREU0YYki4fdD9NbSewU9o
u/tJJdgtShQDXFheyxpQ9QYj1+5EmUuLRuoYyACi3Qb2bWcV2T+46zZNHCH8Ntyd3yE9XGOfUwxM
Ol7CBU14eI9sMXvIxack14X5TBdWnPRn9p7nPiRyff6UW8Gwz5A/unXJyzqrslVyDADl4MC4QWKH
kPTa4+8T5G2iW8D1uaOXyiWFMy/AbPW9RT9Uy5aFl2b8f66emQ06+2/2IZPhvwrjCcYOXY5Z2QlV
XDSHPPrz4ESgR6NQgb/PGwfaS9pu0hYma6FPdy9UsNu3zoLea/uhyeJcMbsyLVM4Iq0m8bqgaNwQ
tvq548Rf2rG5Yba3dTs7R99nLPhvakVOV3RKDOkL42gHPntovCWSShR9runtSHCVdXS8K4zIzHMT
tCDcljkMdbKAZm3PCD2JJ6YqM34VZOHGHY39TOeSOJ1YrCaMxumJGkn8Q4YgsmzRaKaW31Zp2kHN
/MCBu4o1kovQ7q5PGsvC65ryKqbwYo1F4jeGiq03TTW4uuqrW4Vr2sTPUDhtTex0BkVmqZRXshsR
GYmnzEf6j9ezV3o8zi84gCDla0erMHT+VSEpFQOZE/Cci3Cfk+vlmxxVDGNnlG57RFYOBeGn6F+d
RRjoR9rq2bcAQsGOv7e9MhHzFmxa03qxH1Bhk4yxxewiZXGSgED1oqzQVoRkMufnyPUKUUo9wO9N
+WGjxdQaAFa+UX8LLDcJzMlRZ0P1Jizt2ln7XONErNN9FGf4c2cBZYLMT/LecfS2qngZ+Ay6MWS6
4ZyDKV2vjHpMhHX6DmDd8ekn+K0ecGZQ7RduVTOmXcbNadspffA2xkk8dOxMORNfU8HVkjgm6kgd
IFaYrgXCO8Ru9tXIrYwsSgpQf+TQapoUflfqdGplCkG1JUljt6VjhBmMUc+jgWfmuxzYMhSA8XVT
pcGNxZsS16xy2qkkYDYWFCyZlzgZErZC44+2bOFaONtcAplBN4YKV7onbgZSnVXGcfgINHTWAhN8
Dnjs+amk7UVKfSpseJuKL+5HywP8f/nJZwh3XTUfyi8rAdWVpAJ442HgSZyqmFiKjawa4ZYZI+ir
zA9MDSCnHHW0n9UnQGUYu+et07+EZnWzhmcckHelJgQ8Z4/b9Bb0sFS8KVtNe2/5cNiTqK9911tM
r3lM15CAFKOkexvi5gB/9mqPCtKFSNukiagUAbeH8jjxhBMdrcLFK9mnN1ukJNVEwAaooaMPvLCQ
9SSSp24LQNL8gLtkSkWsIXa8oSgukUV99p6FVHLhFbP2DNLMJtFR8KtLT/59UNPGctZtUVLyS/Ca
E3IVsNygB0KecFYTSPYXZUcspCor4UQ/rlx4XKkJXN2hPEGnuCK3mZiqRXgkp1li5O6kRw1639Fi
YRzWX+ILy/Bgr/yin3Y7/XwJuLHgksVpaY9O/tx7jW9l1i5LGm7m0IQSNpCM2wzCyzgZS/m4Vctf
4t/cQt5SjVOGzj424bXA0GeFriT6x6r8uW0nYpUXmht2ePy7Kj9laiyOqZMtAlYOKqiHnZotlUB7
76Re6dt+bg4zXOEpPQbieWqTLk3kVdzVkzMN1ijn7j8DItHLXOZszOLBKPOOD/Z2CNe5EdJfEO+O
M5gczk2dMAq0DwoJXp1rNSfZHEG1qhWxHxx+sl0F1ZIOPyaWgpMTkRPz7lGaQslXHrRKwRFdazCR
w09GC0ZAqHCTBjgM7CfSyJ8cN77VayiTbTy/z9QDEQFy76gsCYX9ZAK2dhKkDWzhh/xxVUHfLfF5
ECIyiStgxrd6yPZKji8S9g63HUiXwf4ogx4M8vUpIUo8L29aV+aCsfrB6mFS2Z23d3q3vmYstQlG
I2rSKHxmVhD2JExzUZW+fApKSU7fuTF+io9zMWFGrXDM/riScOwiNSDSaNpdRhIKATW8EBbDB7z1
0WbSAUMHmNu6KvIvjVcQtjmp7enX2CoLzEEw9oWVOG7g+cK84H9bK3q2TwFatt1Qw8BqVP99o4eL
3Wyw6bASB2WDLObq5K6U2NI4r1Wr/aOndF9eHxx5n7fNXwRnivRNYhlN83ASBCHGna45nW7bDNKH
Yr1ytTTdhMWTJas0rlMbSBKvyrtNcjoGe8ORTnLHMkjBIb1ZleWuaWlr49TfOxXXUgAq5u8kMPNN
DS/RhlJFSiedyURrCAh2ikr413R4eanUdTLsT5A8X/glBamlBRo5mMS2QKX7Qye/olCuCSvcI+2P
KrdWo91Ry419L/ZxRfHo1afliZQZ2BBi/wtZIxItdKZRFjRt+PKeKzW+1i7J5KHRFEeaT1lUzmSI
a/+rhCAuZeDN+4BFLu/1Ki7+rBBRXx+tu2Ba4HuCNRLnl95GOhkNXmA066sX3EiNFcsrSvH/21mk
gBfEJ+R+qG1JFnvLPbXJgnCUik/8fnjabgQKPiucCfsc6aByrdaIs2N84ExWOgdJJGjHwFioNeth
KdmTv48IpC5/EbtfA9Ks0jY0VFYBok0ikpsCnZv+cpobWN9UUoiWH2LBPYelM/QtkRjUxA1Pkyir
Jv4iQHSoMvOJ/GliPWHADBzwt9CGHf+NTRU8kX4iyqksfd3CGcs84WWSyoWyXJjpkc5oJy9BLdsd
AZRVBnRIdW74BGA7hVOAgIETmoRN7yP356bL06oRAcGp2gI+0crIxlyD2bYK4agmXjMMTluhoNtP
jougHWJq9IVso/jlYhNUUY7+PSOm+XuReB3lkCrGiEPCShUfMzyjhcQW7C/TK1Bqogy2u8LwzRf6
M4syb/Hfo/K4Qljujl6j+vh57QpGsHYMwStOZ3LzTfPusyaheCAXVtZDxvt71EL/iQ2CljPz2vpD
WZbk0we/5mH29zSsvw2lF03pzXGyMekqWI7X3Mtln/v1rFcyqZ5Q9cKQJ0DglS0ZExNRxfwxGgaU
W1vppwny8hSBWayTHwtONmdeBHcplO88n6G2X9hekTdR6x8Sr8FByejb+2l3MyS7lLuoBVHiYkTV
uKoKGcW2HJxQQoNdBz8uHJJMzZB+SuGoH/1whl01pb6fgrTTmo8Uo+oe7KqB04T8CkouTLRoNc6j
qd1T2aMJirpMi6z8kak9bBXB8GRhS7TEAAQwKsEVFWb7IURhENr9vwlvmXG+sgDfe3/6d5gme+7L
5kx0al+iNEG06RVceGczyHMjMqJBHC5MnG15S5RzXXFGp5p6R+BGXthv4eMMwfAeDL0k+SK0SSG7
Dk5orz+d5MygGn/h5lujR8sHA00ko3y1i9DypbkNM8K1s+EWwp6MHtn/7JhC1ytHmSlglSt27bX3
y2D5v6DGbqazXn7GDDKj5cI+v3wdJHJ0MPeDOnBg5hMilCavfp4m6s9UG+Y/DRyaL5blDZjOsE2b
CkVNxOv1LnvjrVo2SwU4v7Ku08y8v0hFXJwCV4b3vN84kD6rteMqhryYqr4UbMXoljLqeLDcfO23
I/dRDci0BrfhRghtLrI7UW3+Fo6DWcAdPfT137pXm9VfeJwqmwHrEobYn398WmWHHDwEfy3r4EUM
GJ/kJsbYB/ovB02KNw1t1b3PzTrTPBGlTwyx5804ckrJdq8fJnS7NZDlQxpETVS6+HONhrzyYyeV
/54mdGD5i8HKdtuEKh3+ylHwvaw989PezQXIsFaCQVJP6xamJ5Zlop25RZc+2mEIyK3n0BT4YbXP
atbqbMuJSACanGGBXpcguu4ZRFxOwgoAVNbxCLO3bB6lUOhFusitYyEqIfz9KkNlpdjDzRPL5/6y
lM2bpERarlmp92Xke9OSA+RAcdYmKGkpTKpuiX/EOYfT/uZ8tRejMZA0ZIF42yNM9Xq+IFdJ0+Df
Cob0UR4X6u0VuGL+2pxtl2xGQamqj25ExM+eEDFzL05mb4EgQoXwuZf+0rpg4ZDN/nFRPVMsqxvo
uWueFeOIXznBBzF3WY+yhFzNG1pVMEAplKH57UAELVeraUHxzCf9qN8IaMypUA/W4XxUtGcEcjWY
rRSjDt2ydUfuM6XeTMy9LvQ/Kq/FULD2Kyjfy0LXn1eiAtCuqtRxSihbCBh+QWyvhCkLWWS11UcT
dU7VF3fjgtP0bxXkrYUSpriKwvycIpNka/vyAcF73zLV48bxRRzv/GTXX8dHyNRH9NlBHMsJmbAN
E9sjZ4le8GLGgEwH/L1Xj0hQHFI0/I1ljT+dy/Rg02xdRoWv8T8DGYYamKV0Rm8Bmn7RkS6NRQeO
DIzg+Y1tOwA0J/PX1mhzzTsv9DykZppw47izlI0wK26j1qraNn/RXn8dOnxBc+OFLr6WEeMljUmd
9QhwP8A70zsRLGB24ecCzPUlBOOl4TXsFVIzy7KR3C29sXdsVkcH6xqAfAMw3yju0AuAW6i5dpD2
lNDcRrtborBcCfobJvCB99Y8UvCtZt+9ZgZ/ArtEcEwaDtGLLRX0w525m+nRsLjXxJbB8u1xDUk9
HHw7ZV7pVY/LHkNS3V2d1VRkfpMPrKBxqptC25DIOU9eyT4EwPsqjsVD0/+cxlvBtwOU7yVkm37M
qsui18QaHznT8EqB7IuzKPQsnIu1vlcsvVB8gAjuTecp0jo/BH6oIecG8VdwJjIkvW1IntKcrx4A
cDM5pUdF/UTk26NX/VImwfKwtLXj9Bx8SN6CApfOhNA+UtIhlx9APtIUUYz2EeO9yGNJQ2M/GMeq
yyLUJ0MT/v8NIsMpYKaPcP0ZGS1xosXof5tPoJb2PItMijf1Bwtx28lh7FLdVlUGPLKs088zYD0q
xjJjZW6Q4ll2Ai4bbLEJbbNgNV83cRYclwzhNHdbHe3Sw5IC3xn3jJlgrpSKL85Ht06Twtj8UIbB
wcs2oACTVHJzh5QbENVZ4gtyTby4EtPd5CXKup2qtDQwSqssClmdgSKHebDzCPTzDXDaZCaJQE9i
/bwQxrg+/FfnWagGVKofSlEBIC3D11ZNrV0/19WBx4JfALDwBd2jmeMmGgv1slk+g99V49ZD8GOD
bmO35wESlCGr5iEWRnJeKByMMTO3Vc3ykPSIS6LNZf16RKwelGfiyLBmkdx8FMWWNtdBWhZTqLih
QzIbRTcvunMbP35tKwdScBHVBLsf5AGNBXyKmFrp27kywxDqg+UVyyNvEmU/buBt7voEocBT/6m4
USauFe0nWtKGoIRC4h/oe8q63U1TIQrQrFnZ3oKH1wm5CkAuEKFNvoc2OmyK36AaogqjXeAfT1JQ
Day1XKcMC93EglimxnrcQ4dOudK6PR4X9FKbuUzYnfl6gcpX1hDSSN03efgmov1Wf8+Gjl1l6R6R
vCrVMXjgmtBoqfxQ34zk8N0coLP26pv7F/gT66yKui9uVCxvsMHZJefMt1947fa3cfAEl6OdPLVq
H07TFljhSsLNox0dd6VVSmkXkRl9PNGE8t8B33YI20sT2LdDdzlUQbVXyzRDw9rDhrW8VSnl8I8r
sx65VydprkbknHQ7EumF0/hO9XIGui1eGQ+TxvV1xscL/ghKb6qnOTbsXzrg5fsKsj0xtTJ8eAEw
eq0Jg62S8bkFxJG6572XSUGND4NefFrO6mYdMuaeGxDJid0nlM0y9VXZ90AqGANu/GW6v+DKJbd1
ChwgJ643qljlnjdaVXGoSjR9Wy0QeCMurC6UjdEdSeekg39WLohHoaimaWZU0gxfje85thkK+HTy
rXzIDC3qKQLDWPUAeTs6OCBiatOKhMExFv+b/beSEM0tM+ESuqgzMss6j3gNCYqh2nWszlyGw1Rw
oMtYAF1IQd3uzD/qeN9UMlTuY9kFyfkJDB5YS5mMyA+DqQaGfPsMZqtFX6dK74iJ1M/5SkzK7rE9
3KZ/vrnZ4VzUdfK3MIuux95eePvgNFs7mbKovKeahqP75gSEgh8UBKC4L04MSxvhovWDwkmlTnwO
LSXmKDzRiP2GZ3+J55EkmoY0ktm4bFnxw11jnMep5mNqJFUhWJejSmCs1lQLoeYdFp9kM5Mx98HV
kyKl6qVgsYLe7CqCnb9XkivaTwvaliU5xNEwhGqql0/cvQwGAAPVVCVAD3Te/4w10XU2HK0SzHHP
fQmB3h8DLcdLnRliRQY5M0/GMfbv8vdgGIfi1VF9VqrJYpOtZYjnsc5MkCQB3tgDpPfroo3M5EQr
LeSsnej68WoXH6AIOQKaVvHHBiCHs+D1U33p/Kyemj4LWFQmYSLhkC332XRU7xQVXqcPsfqRfpg2
bsVw7WE1AXJl/Lm2iDzHC6l/O/j8ZNt8hpri9LVzVVvvFF8c6z8ceDFQFw5nHos+K4X0Qbr/XJaj
PmSKS2jgHoHark8hMzTtTNs7UUjqQQbtvsJLYKAoOacCDbKX5QihjCFSwzSkC5n7QQzL3zzK6eQO
AeiQg3ObF2jlcLQ6bsiL2guJ8uGUWW8DsWfYlo8yX4cxc10T5iZckfM6ng3jKrshRieNC864UVFO
WxSoXUgISsU+X8jyCmo5H29flaOg7YA/gvLJuU8TePQvW6MXw05srUSKT21P5P+pNxDiCqZpR/kX
PstWFjLg6WRBtH+8jxl91mDYB1pQI857tbUtqfRTumujeWo1tQQoKzibQHf3a30nXDG/iis1J/dp
bFEHtvvvylY++aUzkTC4GjYZp75l2NHJe+Jn4WoLpE5U08CBlUdSfWBQcatwI67yTm4VtrsLXWJu
714TxwOGX4qe4fH1c12UJjQUVFqH2VO3AwF+H5nu58Y0HhqrU+mxTQgAIDYGw9gOr1JVv3MNHC1x
eP1OxBhR3dVMBYG5EqDinu82/ejy03EQbciHFHj/xAQ0mWcKsfM83As/adFu1FqxkYrDPpWJSkeo
nkqK71gEmRDMecrDhIv2z8z4vFTQ7zAsfCloJaDCkk//8STE8txPJx7Cij43H7OMYca1bP2+kyyD
cEncREaKNarV+A402x6P3AjspAm0WfP+G3HlyV4BGyMsGX2BOz6JFEHkH69H0fFwe25eppOmrrbS
CTdkvTDQkJLtVcIOkb0AeIp8w1waIAVOCDhcKnSvADPQY4gojWhy6HKp6Nx5YNglhJQTo/Uj3cwM
jeZdomZjSV2H/0hnEZ4JWY7t2A56ltMmqycj/qmNHKsgez/3ZvXa5lKGlmMvxF5V5WJpKWdTt5ab
2TXkQBw6x4yVt06lzNtNZ6hc9zfxkcvR62rmMcHws4dcbPxlzBFgy4k7PnH/oe0i6J05/b438i9D
YjlyzUhVr4HDuKjS+H++BSVMRRuAs0HCa1RCOEvB5cjNBhxYcWkFkWVR4C1cscZWR2CfQ8TiC2Xb
ynzgDd7rjQbiy1bBTjYoGg1yRukwQMZ6gpo3qUNRoQEDmPATTd6kqa8rDvuvdvnNpY+vb8Rf5iYy
8jf4R4G8BLFcfS/pdYM8k8ucWZ/AgwC9KsLHuvUk22DTEDBUrZqmlWt2meImzHVSVdnOc7pgqrfy
E0icpLlH9YCYhmSaDu5bbp9i6kQoW5zyExhw5XboW5aZpn7h/Q00wGQmVBO0Gm8E9QvXvjnI1y9C
uCAhY1XUHPck97Xmy6aElVGBkyhQzsylZwEnycOGrA1pHKdMF3QB0i9o9SKfZZGTV/rO2EjGEIt0
DbsH6zCBsJCfHWvErzpSvsByS5cBo36wC9ACwCCVdihsKrNQwhkuAwWRXDe0koXpwT0OECJ4AKnF
Q3BwZx2uLjF4kGqxXR7+I8uaiw2WXkKQUVPxBMqMFsRtqH8pEl5FzfUbvQYVMfI33JYXSohyov69
RKADEg5Ws1dzTCZcjoa7Y6G3Z7S5VtJ78w/g9C8dhb1pVHzgfmUF4Ui9bYIMeguvmn8lLMdZenEV
vch+oaE6rJxoF+R/gqUCvR57tKyzOvXxCTMM9g+/rNhRcvsJPyOYHDUp3lH8deGRHgFtmAvDjw0Y
UDAzlsRsRvvc9ErkZ4Y+WxlkDKEJsNF2Hmxbwce8D3jTElLKAzohOPw4JB78ap7wGY795ivLxUyx
Rhocg4zuvkvHxJNzBpNDj1dkSbOTwH6dzDN247giz6s9e+xNC5lM7nGQH50lIDzq4XONLEcx/nXl
jkKMAmRjIhcOmD5lFnYYyzae7HPovdqZLzJA/Ti1xIpnVaN9NfAhuYF/cK3cqj94BKIRtXH6NdWw
uVl+tUMupuUFKrSeQ35eOzy8QsALZzhecyb0pRr5qZXkhwxEt5a7bkmGsQx97fJSj5HrOOaYiMN5
f/m+/HZLgJOMrh5g/SuxS1IlGyqeIT1fdMs+UT0Wcnt58dZVFS6Om6YTCYQ5TrOmqGbK6iE7cWRU
KYyHOxl/ByedxV+aYz0s5hK9BJd5E8qy6PIYdm3+tTO5we03cxDK3Wt1x4wu0C7jkHjzEf4ADKSj
oDPP2L/NoSndtpbsJ6O2xXICnDieVv9rWgLztruD5So+xSsWBYBdtiLJdVqAJ+FiNxZghRT3pvJ5
aO8AXmAGOHEC3no8r507fi7wueQQ3bfQp/lOc5kfN0XMx8Q7wloyE9lTij2PMkpdEZkkvBiRKp7c
m8MR7MCG6qAhYl3ThMNjtP1w6ekCJdIO63J5i2wUutxHkzr+AEddiDgEuP8XJdqogeHW14LdyrUI
edVI0oAQWJUB6260O2svEcw99ccEEPQ2jPqHjqMP7L2S29pYHO1/T99SSPoSlbmHX/zxddJIMjUC
E/RTnxIrZNXy938uUATQujFSXM+bJORQ8Ppmx5R+rM4+V+BCVY2IItA+rIrGnnRAtUUtiyR15SFX
apPfa8Lf0Rx2ivWtj7BP+EuREiCezFRnmZWxgPRDkL543GJkBNhzms+hb+szgqKt4VkLnN9Qo/3u
0eVeeF1rfit9iSpiUuj8afG/Avz6mBpfvtqxXHzHmZyXr5LKZHItkBkni3vcQ0y0QDSYwrb4dx2g
f+Ha72sNRWK7zA4HNDfBYrBXvK0S6GD0d5/+PrtKIGyXAEzcfTdUbi+isevlnfQXbzJ7vCezzYpg
0iQOua4NqP3iFCj0KC1r3BoyhS50voUBt5hsjfPZ9W4DSqoZwt+AKuYpcRw+ppzE7X6m5rifdD23
xc4fUYCMqWQM0ICWK1prV5HmuOVhuXFosRIzpdjbgH+prhQl5tcS/HLJLo27yS8+pdrZ65NUXvLL
Fuq6DJ4Smn0WCK2QzuV+311Rf1v/XahE7dO6Py/jBIXyZVZcD31sY3HG+NvyklRgxM+u6voux+yj
XXmZhuyeRMUejQK7iddXHpMAdA9+zTh/8yEzrcjTt6YfL0yjHDMKs1D4VR0jlIcA/esbgWlx5jLl
+VxqdHsm3TVvG3zIUF+toXxiQXTWMQJ+NrZUvjSThr4+VfGNJCqX6WpMF6+/jwCaAelssRLZpZC8
NOgCt/3tz9TIPUx+d0mEkimXC2A/ybNHpTp1YHLnT2ttNBTeaZf1yFe8jjf3T5wAbFg0e4rd1hvk
VY6tYh0D96pNW0jeJJn3EdBwAWTmjbmuKjitvUn6C01/iFpYuRku8R60V3OrnkIdJHMT5TWheUDv
fabRKrUkEx69PBnmphiOiTZYtcf3EswZuvZmWoRvrrjYLa2wvxzw2D7jmT5kCaG3HS33IYQPPiAK
5MrFqjgTrQ2gDz4zwmiAhptGGoFiyLMAtdpnp1kAtLjK80hwLnP3uo62goHhsJlDazsrkRfhjg9s
glc8X2pseyrjsVAsIdk1LrDxssIBfBz0grBc+eco5QhNCCbu3fX0WCZl0keoBFJCLzX/3BAOMS6H
kvDL7hXepBMub0DYLrRo42/oeFzGkju5hvf2UsY8yC+Xds3VrRFLylZ1srQ6EpObJ310QyZfu8tJ
R+5Kyb6y4r4B6+fipuNCMQsbT/ATRnWVkk6osx5Iz0/GMPYW+pExU9V4cZuHJS2AFBSLitlpRLMs
BIOxQ9QGs4akNUVCxuNqWP+6YWEq6e/PhQCaridgXmBqvZrymH31yfemCL6qrxNjqyjvx0hfuilz
a87VNEnv8iRQbpUj0RQ4bI3Bayf6x1znw49fkcjp6gUuDTedMp51XFpsInIDze3qLOYRqa6JnEP5
FuzCmMElsE14uG5hYYpgTH3Lk1YORo7V2opgOHV4SeuBWWdGrqgIlCnFKwkgqEP1zbI+N57Fx6OH
xNpaSJfEmqAiaoefV9AsZ+QPsOgQfX9pjhEA2XUu8wbsmbAb29atmu8YvaTawCn+8fvuYP5ocmuu
7x3UN0RuMVwUXmFbKVpoRnaAw27z6/ALfYa35VBqMIDR34bKMSRw3uz+4RynEtYQi79Vc0J2UHAQ
5N7vfQazQo5hiCm63FmgTItR7pB7k+fdbAeziBGe1FJSxPKV9UtjL49eoU8DRS7rzjWy1BTFu95j
mac9zr1pbe3AYt5YNKmIomi5UHv2J0bwCoy0YrsQ9pM4ljZJzArqMvSqKOMudGb2aLdfH+q4NYB2
pO2zE6TM+khY+iFEKZGQ6ehnSfuEPbHc9juv81CWUMm13W8PNzk9iA/u34QZBllOfsco0UcpL3cp
PnpW4mrSUjAi9mDKnNqZZyCD8MlSRG4VDS6Sua/3/uhCupR0XrcFQWNLQb3NpwaGj1VjeEImGAAC
eHa6Y/UyvtomYirvaum6/NLo6dqThv/bBenTGGwcjMkTRCVOA7MDVveJfVuRzyntu/XAgzPCufDF
2fVhCDHmJET4RnwdbhZ2otUiumOSUnYiRxYCYpp3FJnNXkl3+mJLtMW7J/GkCxK1Q5WkiEosqkoz
WF3M1qpeMnShdhaFq7y92Co5K0bO9d7TengNQEBqPBf8JIFAempklD0EMjIZLYP6eY62vZWQWN4c
jnI5SXKq37n6gCDhYMc04EKRNHHu3HOuF/CcbW7x7emS6LQefFkoaRCKb/kn81QGPW89LLncGMQa
RCYLRianl8McwFSp0u7TBfklXpXKuZV2RaZ3S9G92Vzbz8CRSGJeeLuSa6riCQUdUSiDeZoqoKmX
0LLwRu4/qcl8qrxVAJIohB3tb5sbo2jDEFQqrfBfTjM3df4p963nEd/ERZVSQ5JHXB5nxbqYEbzz
k6x3HJSrUd++qrGvzo8QLD7nWOi7HSPLnRbw9B3hew7I3gmAK3hOAYcyVs1IimD0gcJyA+KHxjkv
ySNqrc3khC9820PwrjQ3zIU4fs2ECInfZlx7cVirHhH6qz+yXmMWYdjF9YSxloHytGfWcDt3sQmQ
ljbq8chAtKPduPRNPFCA2qHfajZLWRdKQCGMZAZP/v0I7npVFkCsnRa9F4qkaw++lRYVXmao/jjX
jGteqt3AkVPFPKmNVHPFFl9ZMYtuGKNsJNTW1MyRE+gSAia4iMDkjAsXwLoYCOMLwnUjF/NNftCR
FoUs+wHP5byKztmTC5xHSnv7QSp7SmAYsTFHI26q2wSompJo2O+CIQLIbga8+u9SgojoMRvjZdyx
LvflsKY1bWKBgL1Gn3EHJvZVV1zAHhZVugqnEk9whfNjnE+xk/11FAkK7lqfB9w0SlBIXtXAondi
4mTRAJHUzeozTtZ5pKcbzZASoWtABrm0I9qqcIuxjyKJanuyLMgzxv0F/FEX/o1A1v+s2pDBJOk9
Lx7oBp7bF4nkwqyBU/dF763XS7aOWZ8JcwvSyfTYzLg989rmRhOdFv4gAv0OFIDGmyX2LTAi9Zse
BR1X3/648snU4EM1UVBS9RMbGn38EZRCfZAYElZAvHAXlA0DQ3FVG3NK4mndj4EYB2V6DjVjUqqD
dkqoObeHoWnsvsJUx6fTXSBuooCws5q0P8HSeHk7eBGKAJj+gsc/FqEVEg+K75Q6P6HEMfB//K0j
UjRx0k+RowaAIDxzld+A6XkCBQ+YG6LLrDoUJsZCkryKaOz+4hRhmiel9WzIfHTdthP1Ms4BARib
ZS/QXgIUtyBHYe3Xvm6sRpa6z+DP0pU9RVwAvPCtJUYtD9uMkoFs+HLN0LBg/Om3UBklarHyIHze
p4Sr7L1MNeZcugD7Cnj0HW/ibyr0nEAbUgecA9SeT7FXz7Prwbp1ItKQ7f3mC7iC+Nn5J1g60fUa
T99mo9SkdAsMCLTWq7oBnuAoz5t5p7c8D1UaG2zIwvpk78SYcw3v9pqNiU9AEyv/mekAmzADyuCY
KA/lVemni/6niCEweLTq1+EI3x0YN60ghv80461dBmUWD424/1cred7RcKblLoLn79LUX8zr/+8z
VL+nhfUwi8xMLFF6Ufb3iOHXzYX4hmLZnyEGLRs1d2TW9AIJ61a7jqRIFINDJQxM9JogfsgS2w0w
CpSqKsGc7puIBtqnwIWGYKqbB4kbDVu/3FW5ud1/8rA2h1/tHzP88UccdRSiC2lIAamJ5r8oAVJD
7+b46flgUOf6W91mx0wRFG5/Qc3RzFHVfhocDkUt6Yg1bOAQ/uv0rdl1xVdJMdcygVgzTzA8SSgf
ShTGjQDadGAHYrtKXqH3nyeNfbMYl7Z07DfrybpcvTsM8U6Lgs5gxUUswu2rB1i+oazauqRwXq2c
Q6pr5hzXf25PW6C5btCKosVdn64mMSqwR3GqwmuccfDGJ9Hbk3QpzKmBonJdXmWxu888LPj0Rbjt
UNnmXamVOQWPZQQwiD6Ovc2i6mQlrc7h7FWxskP1vnpr87ysd3MrxFGkqBv1hBIjOLIEtkR/yVzZ
VtdDQd2ofghStnKd1Z+gxwGHnr4cQxLl+448V7CFKifuhYlnt3IwYWGxA2flwRZZ1Vcnkvz6dyZA
pNLwihKv+r9yx+tnjzgscIyBIbuLmBAphuXiYiqCr6X87Rn38HeJuSkIa5rWg17SdYkfMV13EsB2
KP9qKYsQV8XYG8URGHEA2XUdcfTpwDuE8kdir0htVtm0IHX24E3fx6Uzz9jkSdubu7o9teoixQ4K
R1MbOipnDo6lBTqQ+WTDrlvEGI1MeMNq9fUuEHhw5QFRp9q0KAVdxWFaSTCERWJxGIVSERqGJfTg
eyc0VnXznww5K9BM96x7RfEjdSxFGaoA+tV6paW6a+Funpm2nX0Frouod7tpva0J5rH1HVq6kJOx
UX2j5928ae4RKc8rPxme+QbV0G75tRpsCroC7VMVClC+amcTYBs+7PGiVhPt2oiuI3bwjLAe6+et
nL5p0YCFjzASwUJEZp2DMEwanzsvn3DC9na3Uz3IBa0vSHs6pM/0ygy1lhzeuIsqaLpnrJ+edeUR
LpeY/L6Kj/hbcCbBW7zZ2XibBUukBz2OmccT8LeJZRHrWLn85DpQsdiZVBxZXx8DgmH7ygRNem9i
+cSTykx50josz+3VUSYRdM09OmF+bn/L8DAIDVDzavLcDm5gQEzIdoed4WGrIHWTfLzqzzXbhpPl
9vlxngLDj+PSaWLA48o4DJXjwhcg2O7gyNI6nvY/s7q0xYsE379RHgyI1trYRfPDbmFXtssOGb5H
aT0eNxYrW+1aRq+KrvgDVYwniim3KlnbfP4mAStKirqKMpIJyDn5JPOQBdJ+kME+GX6rm1Br4SQ+
ZVMGP0ddFHl9WDo01Z6mjVgTs63IoleKg2eJm4vRMX/dkuft8u7FuFIpDwhHdt0fOSV9J/HhOgr/
QrttgCgNEVUIwdPzuLsANILjtK1GpAVVtRZnYm+YnutXyE5eEj1wyikqITHbUSAnq6UfB/AfWemT
qvsjgjpFY5e6bbCPawD0idziBECFJDC8Y66dkrPfFLZhbAKavy6Y/XIdqW9HVnifuwGjcko/LHj+
DpXrhe9TakCiSB6Mrv90Fv/Uy2d1MMxqjn48l6CbSYptLCmhteH7rE0QjabwKGjDY3Oke2jA0snn
2nvvbTpdY0iNsBj48+yyWDgMXas3d7EkqG7cYtN3q3ng4m8Y10L5f46aAwIfkKvV3btREMHRQw8e
fdNt8b1eVbdknTd+fwcilxsXc658aJCfkM/nERH586ZocqVTS7nDMZ4Id5+OAkGbZwEa79k2v/u/
uRHPBAVNfIpKS64UTRcEpiqFU6DmyQP+Sp2uHU/NDMbYZ/Z0JzaWQSRx7iTWWNvOiMSLFOC1Q5t1
9KrwaPSMop+Si/lCbjZpTq6EmrwewKPsXp/0e4Xm8xVXLszFVV/y6ujng9gL6MftN0CHaRqTePjk
d9npdb4mIao9HvmKecl+oeXp5OT1uxHboKN9b0lyYz6bPiyEZ0jVGga3SLZjVN4XKQehSlHtWMs0
/k4mErQ6ydq5nIdxTtc4jA+GIGRQ+MNw6NLg+hBOuvsFPq8VjJ5CYMN+9xIkaqV4Uv57adD4CPbU
gb0YVX8NB0bfzrIP2Vp6Rb/88oJQRMIWOShs8rrtNh8uTOnSQLSflOk4KOgVuaBgMi8dZxr4NYi1
GhKJsJgZJIJbDwsdBKiE18omu8uJBO2ZZPy+NJX0Z+em4+arbym3k4hS50yJG4bDZ4CjWvE1g7HY
sntsPQFEBm2nEHajY2Q7fWopJ1jgKJwZVfSIiKzxE1ozZ7Q7JO7Rrgdny9PurYF12+Nijij2Irv8
/pOGHFgiduriu271BlUey9kNm1xB0GTu7nCaDdsi1h/j0Ek9g67YRFATTV9ogPjoGAb7KzJHWQvr
8gWBhNPwu5qJBCfJL3VPA1pOcuEyI++vHbF129iQ4VxfFjM+I4bU0iTVgBdgZYFmA/irwxbN5R0C
XmnQXA2pDL+vZPY68xkdxesDkauNUZJWDa/qOM3Op12OLZhH5twmRzm7BapQhwPv21mV/xgd0Fap
InzbmQ8fUAqYIvCAZAY6ulviVsN/UF4EmOQgXy0zrG/vh9TRgUFBzVJJKSeIyDXC15s0Vi68TSv7
X4QLOdfo6aScdQQ8OPL957c6NK56rUtpZL2hOBGIIAd8sOpuUoCT5H2lTFQzCrBDu0EfiahHImil
6KDRAMiiZr2ucdmK7mqU9Fmem7RkDB1nbiuLWZ3UqmPz8yMxQHzKNf6i5+m4/zNWx/oPK9scBBsy
Ewq1WiXILXHI5ihORxrn+TX4OGSFQQu33M2EqztHuhW0vyAv0I+9vTWzI6/a6Z0VLQCJ3TYYKp6h
CJ3mHL4rBdpIg+JXLj7AxdtiTmgsVINPYzELHDiyhJM6zBnqRSXy0t91xKznEHAnwrjE3NqEg/eg
UD5rVBxvSA4wf3pboKQvWlBkUsaYfWvRztpST5j3ORJ36rO8dpf+gMc+xQWlJNPtBDwQMt7XlrsY
msxSOB3VACnfECkKLCV5Usi4VbCtVBKPMyA/9Oz/OrmByK9dGuVJ1Tsh/N8EFPFPOIed4GXD+DSW
DBXk18X841svVh0Fm9Xlc7qOfHmI/SJv2c+U1CBa6LeZ5HxHHKt4HjisUnEw45IRVjeEMdyhHunM
TK5I+Xju0FaEQt9l23Tsan1x/0Q6mlqi9ul6GMhtAIpZXDmZNuhw3U+DDVxQHCq+BNFDrJyXeBlc
wx1rlafCfyyr47IbgNrplThDgHqDQOHllj51jGvIFz2SK71XfBdxkZRLYYiH06PHYBlTyurSCB/N
9f3j61qkfnlSS1wjR9fOGe8LG02tUp10DqTP5hbi46v+GyIiPYLQbjMkbxHjFquMhVBzV9ktW/fA
xPma0CN1Wa1uad93RJX8mzKTj0GYKT8p2v72uR2jc3kCUTGuaC8UQn0y5D4tgt/nnwa11s5M+u1T
m9XSkVlD7tJMDVKT10Xs9S5su7CIdZdSJGXBEf3mMKvh3j/PHAW/bLLU+zbNRITmL46+OqrIp9io
ZEuHlWGDIBU+8EwBAgdMyslykJNOYD74860ubGVAcKU9k6HQMXGqT7lMBEDXoSqhByqiFMSzX22e
lmK/6fs7pu7+qYLBW8qRCxhOI/8T615vLx24XPPfpvinYARhpmkwBE53Ja7GxbvzUyaiRC5XASBn
j3OFhXyl2uLX9zKWFjkM8FBgjB//nXn4gyIOXMTkO/KVkDSuXb0oBL/71gdIS05Mkejxj7XQ8hVO
1Ek4v31BE4uNcmjZG64Zkj8YQs8G9qCy1Q+elsrF5Z6QEX8eKm+GebXvburxgOS//8V1oN3Z9cHA
DcfMWw7SSg9o8K5vdsd/WjZbRkYe1sJCBdDsgHVkXoCustTiWvfJVZFpHPJ742d6nHa3bViFa/UF
aybUnWxMbGA19WpFXFl18Z6R4AG7ImnY+wlEKnSPM2tXvVq9KWfd6dk1gNTONBKq4WryCIZvVQx0
UXeZxP+qVXZgvmCpkJozXkvZpIKb5JAjtZVg/LKTaUZpvnK8zyUyNa6ldbgt783d9mzSYHvrSUxk
9MPyv9iEKAYVA0BZwfAJPxNkTwpfaEZ3kq9zrXnlI95HbQl7RJ8GEBMT73Yzti5ueDXQgoaDxvZS
x87LnpgKs+MjMDY+rEwMo/2bAVMDBu2nHtK5M1Lg7fDsRk+jSxeZEAzTE3LNiA6m8DrDspyzaiq+
EkwdDBRcfu4v1FjRcODxHiANb8hFyS4ILF9lG3t/R1GE8RjYkSVVSdx0sTWnVS121q5S3sAydjuu
lTX6nlX2gIhMYysD2543XEE8mC8dpWJFWNyFQjM8tTOHt8ND/Bc45r8hJNwRh4YtEm7H4SiYSKI6
/GBK5nqHRPZvOu6AJp3g86K1IIJoHhArcTUiQmxC609n1kBo4WLU1dO+6qOO1aC+kGr9PVr2tV4M
vpt/DzY4qPjof6d39cK+/HqtqbtmjRiMl8qzunjDhQ5a4MNGqUqh4oHsiWbgYGlzQulH38KNuFSN
ctOVaMaksBsPj7eVsBoxLRZ24cl1Uask+desIb3+MDD6tcMpJK6sEWF9cWWxxu47MaYDiQCFlAvX
29kkdI5PaEOy3JKX5KfOlrBgjCHJ8PXkJDpz3Z1+SqZZdgC7sRZpjDelmRI9z+APAa92DgqkIXNo
1/X7ps0sTieqcEaTKrn/g4SRIzMxnWsaKOJR/6YIJo+USeGG+af2iQl3rrWkudSQ2f2UthlAqML1
v6W47unNt2QYKzvQ/cvLYlJqjL0e9r1yd7x0pMPOpTx87nPElC+aO5nArvopzneV/1KRkq4NHs99
FuKpOM+rAxNhAsoGk/LVFUpBJrBDOrDNqo/2j+9wFonZ6Hbm7nd9vd1PbD4K/NibyOyExL6cOSn1
oNcDE8HirmtXqZZrWAsaRLb4So8l2IccBWmQhD5HQe5ypSrrGmz249LvDJoJOmg4g8hWTlT6oORm
Ha2EIiofujNf86hGReied2Cj7+c+VisomTGu4R9QudbDe9/Uae3x1a+NXKBEH3tG/ox+fUUtmlQR
/ALfw+fRXlYEU6b/uWCSJ7miM4z3qMR2V7MfS435vDTqiKgjg7cRoPf6iWfj6h107twEmdJ2hBLg
2uPvr3/ksj3WPLzs7qLyUOKPUZHCNqKficbUTVeGMi+VgsfxvSspyoUH64FhLHa4qVZr+mVuA1Y0
+PVtvtadkUxtITPRgOGaxqS3GHtMSbGsSgG8i8wPoz9L5dUu4MtRZFQKan76navEkUo6BKlp1S22
xxdUYj3p+NRcrsDyGvtjFFnTU03rNimBjMT/9ZqPdSaBznFDQWasPcTODKZTDjXZZM8pIC85r762
egaOa8djNIhKPXl8gSmScsam8iZvoZSGzVNyX8wemNLgdTsarmsdkZRA99y7127y0jjEQDFiOJjy
/LogIyVFbY7hCqSTs4zXnpJRg1deq3e4NouaNF46mto05CACy58WwgLT48XjQxR6lokMwcaSfeF4
NG8YVbEFcHBF3YWH6T9W7dd7OK65TWtHxZd+uRQyK50Ou21CtnMQWy9Y9hTm2GtHc9cu7MXO0i2l
87brE7YUswQZOGg7hedsdEfdkstfQQ9AATZ0iPbPFTakESV2oyiK/yj4UpYyxfFadyNJs3zUbqsh
XnZSksbsziMSJ/oT8uarYYFmc/ssick18GbyaKuG2w6RyiqgsNf7dQ277R6P/8UTSnM/1KEoB5w5
idL4BWpVTb9S3kxwMntvmvHaii0+tZVZX0tRRTMunvr1lt10EY39+2bBsZexkut7m3t/bYdAtJPs
/CZZRyQOr/6U5e6FPEu2lvVt4yc9OSAFwGIkFvZLofzmtDC07FKFF/Zv6pf3IPSVngtJcX6ezKiC
HLpZYV3oiU5fGvY4Im/s8wXu3AhDs4UxmWKgtaZcpBvQy+1IxfLhylWVBJl4XrL9hW+5eXEogIax
btqmQ2r60YiC9xU2D1d/XhFbfudDJASkxrobpzO6V7l82GGEHvS0CrZ8U/xy/WHi3B5oECmdE1hl
47GsC73BusEPKq972FSmQUzuWopRPCVi4C/8EOZpLcTtyBFCdUUzn5GVP4+ZR/CctQZbwkTmlY6E
cwtJ8ARbAdUFbkrY+QMoCHz2cFo5F5eRlXT4pS5bv/88m5302Q4be3Xr50yFHToVaga2UUYVzqSC
HCgD+wDZwiBq5DHX2iqDA/uS/NcLs9VsFvDyVMDAJ261GUE/r4g0uo6qSm9mi9fdsjSx6vmcX3/W
EoLOskI8dx+2AjUpKWREqAAVdyu5y8GIWgKq2TYizxgJ9pdtthLfEeRPScouGYxgiJ2aaFagXTdZ
EUi1qnDOh8R3ZiptBGqXi1h2LmH0bnETdbh+m7T/EQq2gm56eAlNiz6nLRON3jnl1Ur2hmrpVrqS
iDrbdWuWkam/FY8g2bgKOXMb7se8Wg/Utj7jc8bUhFSWAi5YVZAHulWwuYYvb6lmgT01kSHA6HnU
ZDK86eb05ywiDW0PteE7ezKTkMesyzFb3s3j18w3blDIhtwgE6fbh1uQHbhBF+LqVmif2vReG12o
PpBsUm71UxizlXtZpZeY9gzQA5YpX6TPB77HytJnTscBUm5OSJtIM15t/yM0/pNctnFtDAdVn24n
n2vDbCj0YAbfSkj4nH6SxPbxCTjZ0W28IM9c4vptDG8dPjg7kqkYzbhqmIfAj05xG79oWxx+/yKO
VK5epDV/ZPUoDgVzZ5U+bEP708e2NTtyHMKcBs3pbSB1q+jq9UkCBfin1/McS+BjyJMUypiQKjHV
sCYcNH/K1BJMt7skxZOtOhblFxJ0wWyBDWHP096yzI3EJoiFkZutL2dWrD0hscwQdxH/zf9njEeG
nVbUr/1+7K/Gz9bVyyiFSqvD+Sjb0y7uQBSHv/yO3tYnJksw/RJb2UlGLrhDLICh7kCF4btoQJlb
yBU6fLv3Qq2w8zOAGejb+MlNNqI7OxjLxrbVcf293umhMSkjcIWIEH4AtApyVjLq0TYF4QlH7tjj
VKiOKHwuGus7sOYBS+JUM1xSIPZakQ/9iumhiIiqV2sgG41SX2SbGcLMJKT/3i8bAl1koc1HyUEH
p/GAZR/y8rPJvYTN0yB/W36EvxEfgxlPRuJzVIxJ0AoI7OAB0WFSJK3SWPpyOZWcJuzk9IhYF/Zr
teNQd06cAe/JtYfBCmBMfLohYqCh/UJOnhmpLJgCgEHdVvCqxb9sZXIjIuj0UPvHmbtzyPbQA6az
AuRwIWqSmMXHCfmSl2xdqLGVnVfYr3gi7hVoHYnuR+9wOBxHQSIEJBHE9FUMdr2XuyNhqfLvHYEv
C3K8bMhzTRIatO32uFFKXCKYFXNLycABG7360qE4qtPBjbAon8om3k/HmKIxC21hMBjUkc6tOot2
UMtOA7NNKkCowypQ96pUH9egDFaU/0289NJEBQ91JSxi/RSn3gd1l2NBsu/BzaAyMfsQr76nQSSM
cF4YmC7ynlfz267veT9MQUOmI7yeUtUEAi1nSxcBEuj4sjvx1bc1g+KAWxn7t9RGF/kiirXtLlfi
qqI+az95t8gLDLCZNsnFhudy4Ro/7TA9oKclM3ElogG781E3Wqk772hs4eFVjONgKXXAau/lv28k
BQTVcX1qZn8xgP42l+TvCKpNfOy9Yp1X1EzbDko9zlDvDE1NJJHKJn722xq6h3HaOAmnXp0Lwvka
quuiB5IMLRJdFTVBRwoE//rwNrmbG3FtvpueXv0cTrq724Gjullyvhhj0cOW4ZRBcB1HBk/wf74d
0+EGpXdsBVSXLrom6lXnyKw8Oz81fUAEhEccZOO0fJUa0i8MUYN69d4J9YKINpXPXLZJ9Az13s5b
5AlM5XWtmG1SlP4t3RXzE+Vw/48k489Yce1BE2DBSqd/1PQ4LKb75Ave2iPhKx8TIHSvH0biIo2s
denHzdIR06hckWVXbsRcXxP50KLlPAqlIQkO+/wE9kKZFnwEU0hWLsRRfvd2GTjZ6enHnJo63nV6
M6/M+TqLLLiixxFSzxi9bW+T9fDLzVvvv0KWExrk1TnK+u4N28pZgZfCMCsFGj5wxutIY4Qr3+GW
cXU1bx5GDcEK1slFfIWPhXCYygVBVMkNbqUD+ll0ANgkAnp8bbPdVXsV/ATRQf7swn42BVa7htu1
hqtEGMjgNrBU6j3TjkmTnOWnDeHGzG8ucBIDoW8N89rS5FRWe9FdAqUljYPaKSuKJlw57kL6jMKT
m7iiUi6svFs+IwXZg0/ntGI3ar12eX6ClmhcJkTzQ9WBsfhup+aAH+ZX5/m9a41Fbqhs1Q85z40/
RT/sapqWj0mWs/FwCOtu+7EdeBTp4SARLQhE2c1TwbO1lj0MrnnAdL/4njBODomqTvXZFo+EeHk9
GfZ1zEZmQ3XUr8h078uyGkbZefWxXc2gw8QJrmhuFzJvYUYomW98Mmv0YZYB/G5SKN960bWr2GpD
ED24ahWez6o3rydMMLHL2/WIllk4qLHbU6RZ+/9ePXTT3vTadWPDPrz4Bh8/WJfn2afVXJBjd7DI
wmtdKpPzy045iHrEzLoB3HyFXDuK13hIVRZD2eTp1blMSZKOFHjhN/c9nJVr3U4gYcsETspwLsrp
4iBEc5dvF69mBpdkCSmHwD6fxkXrsBvxuczAzMPl/X37FzA1uvrNz+1U5zvA+F+h55/cugm1OKKu
IGvR6TaGWRh8w3lcaoqNdJg8mZbNX08vAhv5yhc+dNAag+0c1ZQn03Q3v//nOfDE84fg7/0VD4Ex
eYwj3t7dVm4XPxrwEjGYwYEHm+Ja50JbOeyHFUqaMN21p9Emh7RXOP65AgziXmOWhUjakwnv08Oy
krAFOuyH5dB9yrIfVyMcC3qznqULGMk8K97WheAbY/XrhMfsnyhsvhv5Ly+bTqDHDfc4lxdCEKHd
f/nDoU9gOhESHvi2bx2rEE1hm14Nmf76ty+3KSzl3STENcn5j5h5nIpzdveRL+vQIRhsc5O++SZj
9Ke3pVhyKtFA8EnH94Yms93yKNkHkfeGiLUXtCSE8IGbNF1YzzTmCjHm4zn70hyN0VdPy9shmuvo
2kZSr7zMUVmClwO61rqehOJWbDtYC+lwrKURvGWHtu0EJgRwunL6xwM+stdhUpWwJKGOxWGha2SL
5/WyEbuzTWw/t9557W2MVE/413dvPpCsyelj+wQOdR8AafaX6vTozxJV5VLZAuKtbcVmRziCCU0m
0g8XvEgHyrRkgN9oWR21tvYdOEyh19zndvM2tpJeUumeFeJkNJQhKziW9Uf6GoOjLS8J38SV+Rkz
MgaUu87k5zDcNqNJZbL/FuZG612SEgOhPL1Uv6DV6Puye7+KhXmXv3Ou0l3JdTAPA0SxZpuwxquX
wAgeM/D6QU/hvJB6KA4BVucGXxHJuDbVegJ85rMSr56SsUR3qS08udQXjkYmBd9iaw9xMK6YBbpM
76676q8vyquM/FFuyJsjFUhDF2N/2P+MPsnJcW2zu1zFgabsau+7mUiXWCr2CFD8+0hzXz9mBGJU
oaDbriD6o04eN+eYvItFreRlV+AJxim6VhbpyWD9x7AGoxi2Kq/r4WIfaxxAKuH6YJuj22xuimlY
f0Y7dmbfAO6gHBW1F5zRwM4O55Qd93PMVQsd5muE1D19erCZsqLFuFWO2RGNPYSmF/Cw1kH3fqaX
JYtuxk/Dun02a3STpl5Cn46Mz6jhoGHDBKUHifCdJZPZ2mTkZUBGPLWk2QCZGUu/xiYSR9jkhENX
j9902GxypWE3gZfxRfcnEuMMrpMdT41pQjPVhixiNi3Lyyib6XWJEwyT/H+AgkGpLLkkl298+YlV
fkKXRx/dHdVFHq25SlpqpIwso/GNvvAUlzOmuzIMpueaC7D2dlpfpXJ8+lPXe4gNZfOp9Q80G3KM
Z4FuTrb7OinptQaCb3CEoiuefVK17O3Cavk8Ahjqq2MQd//Dk+pEqVX5KxFLGjX5C3qbuWGLovhA
ru19umJmPOkD1YvhbzYrGr7lCq9z4xc9hhH1mYlIWXQFEeIpWC6NdX0YnGZuQMCbGjuykeW1Xu4P
Vvogch2LMQyc7rYBX9cCPhqX/TLwM9m17ifu44sPRmI64hgXY7v4pjHJ/avuWD6K/Q36AK++RI5a
uCOAoNCi+I/VYqtS0ClnRhXWUj/P2CSOTbA39lEbf6gmEogpLxuiT520z8nZ188x9ZIKlyR627NO
wcT9E0ouLLXm1KXJtZ/k5fefNinxBPR4wpLMzauXYfDhbE8fet7fd8mBX/4aH1vmqyT6HhzMbnYQ
uzh+sc1nDCTiEYLRP1mKseS5+9eLX9DmdriO1k3Djo0tHaGJF4AVwO9hHp/mowJ4mTNTG7KYSqYR
WfV/KRj7UJGYGXUWflMHann9E1EIjCdYhNbBujI1GdAomc04tEGB1wBP9zrx28G8jPvF4HliOMVy
hEeC5JmTlGKt3PE3ogy2r0qxwQqeqyPB/zLsggyB5nlX6J9eSB1bvBJj3Yb51OhQDJdPycnox0Lz
540FHWFOGJdBqJNRau/MzrG5ZVOk4/7mSSwvVOqfyTWim/nT81NNRDL9l+yX9dAu5ny7LSFkYrn1
1ZFAdr621fx4zBOpqC1FsLYQF9TKjz2Br7085kFM0v7Lk8gpq5SLUHPBnB1n2kxBck8C+iov4usl
g9oE+OPCIgdnBBabkbj8GEMrCMP2bzc6i7wu70lhLZphM3v526hC6oL0RJ5zjcUV0cIC5UhQY/E2
xaJQP1htEyGXTy9lA5u7R2d1rkYmH/ycGk0JFhWmuIWeuHbA2dXZubnoT3W0X2VnwYBgm2MfxHY1
rbJPNya2Ut+gtv1ex2xn8AV69ag8tqH/iEFBMV4rjaWfERUzvju+OzXXQTMRI6KGFV6P0DyGa3bZ
BVTa1EHDVcpc0lg5kttxogdgEvRXaL5UEXs95OPubdzEH/bABTbUjcgxs41Env5XpkB41viohxtE
QdUaUItuqGnQCsAWqML4GuvYuaJm9xtUcdVLB0z2zLwGVBi/pQKFv7IBbpGXlS4tFashGWRL6BCu
WRoN32eA6S1k12FFlnYlXmap9L4GZHnXbyi7oZANap1ouiku3FvXEZuREDLGw2J6NQ0EE+LjAIC9
iHPYiVPDig+htobjubUCGTgidUxulEexfyJh1psB+wxrjBTeW/7ymMjXwoOThmsodL8hqGcU1j6o
YER2d+W0INOWH9aAPxfHwnc+0pv5nHD2w7I99bmIa8tovKVc6J3Yas8b6deEV7ral6fiDwpKqBbv
sSusBPdoZiSXKLKaGQMQS54qt81KHr1vDLOiJzMSBkJ6d+in3MYmdGajrh3nB4EVK2B5jusvg6QT
1k+E/y+MRnjdoM661e9LMFj4VFumiYdjcUkbgvKiYnWNZVxUGgaK8zqBsyuIE9spwsn57jwFGF2H
uUW1FPNZ3rWL1bZ3j4JcecQhDLujKQC+iTslsXlCitOH1zuh5W5VHaHANKNrsQVHZTJa0ZR6oseQ
t8mCkDUmL5kuwnlr3h9fdblvgA3j36e17X9uWknCGrZwA4E2b+hFpHEKayZyaGYdVcxiLN0S6Ftr
iEbuYOuZaQddq9sY+gVOoMXuIP56DfbFEbb5spFrxRCEDP/AJPnwqB8YCZ2YzNFiD9gop7RO3vxB
RJW7HPhoU0UrPhLUPEqFg5NGF1Hsc4AwyN3n0FW4TB7pjsVQdLNXHATFq+hN9FcbojW1Zn/Dg4zR
vBgg9LiHHGja2icsO4RQ6dDpEwZlGVGGFfEaWmHOt3SuSkIiIjmlDrQ2xbYIFXJxQ7XSOdsq55aK
XS4e51dhVCbm8+Rz2nAsU+tU/0HyCN24BC+iZGS6rCUeurTWh21F9CiDyxU8bevJnyc1uTS6ol5K
u8DsTOJoZ6QRBWcCn0B+E7c224Rg9C89d1s7RuCp3vYPJ69rFkCwvil04O2tVHgeaGW5HdWAazkY
uPyZQ7SKUaXb7njYErcop31wE37uAJbT7od7X35MP6skKlLu9UFc74/f9ITncoj45T4JJJkOD3Ol
nKBqM0rJ9bndKfLND5qAT4V1dLVZNl8nWtydEo8XS2/KcnboS0ORVsfLPJ5zOIcCrSWWZ2iAgBpn
e8M9FRDlmpcfchP/BpBE+uyQFSh1LH2XldGa/SWF9+ORYxYVLx0CRYy/o/4RDPKLbdFAX9P/DVOW
sUDklGnCi51lSZGsI2d53vKMRkclvQxqe7j6ljwncSz9cYfaM7CAudRmi3Ceei0craD9GCCvV3VY
tPnPE+zQELgiG0X7UN8ZLp9PaqU8Bkj0gAJPWe7r89YvdKWd7GCTo6i0kmK3SlOwSRWcfZKvvUDR
QoH/vCIrZpYpjnusx7Z0SivneXCFeA/zYpWam1/cBVhYOFKGQQlAIl49SnO9dJTCw3Q93v6podwI
uQh8vOtgWK+uVUzn6fw7V31yGUC58Z1JK8z2wmRIyqgbI+AY5HSpPXCNOvWd50rFlrKH0sE1K9WT
F5lpbCN0GftVgK0RmW+T7J725eA/I818hqlMIY2HDdoCy5o7OGwQ49GQYjdxPtKEh2K8dDWFtqGM
PpJdocpiJtG5C5MO2LHfDpNSEI0G59NegihBp+nY352J9KytjPVH498dv6kWuByqBSILO5aokGYu
o7+vixiLCGFuPToxh13ppGpIAEfDdykcoUxrsS6Fpo4vfYXp7redwvzLbgilT6TiTF3OulyIJOhd
CciRip8Hz25m182cdCPy6uhmAtzSFoe7jaIxiypC2oPDu2hFikF9KsJaSHrluTk8HiRPuVavShTI
bwAYjKpCshuR5SEpC/X+ieETS6VOb6bSqqaasG51BktScysqQyvAVOjXT9LT1qWwS2GuvAIKqqKm
YXYVjJaGMiGMBL8XgEw0U83dYsgPlVFqWX+3g5+izKJqoOfFhhGlsZd+/teuss33oc1txYtKoZFk
JIOv2OyMp+6egNTGLnbd7sn/+cVS1Nv6anwLRz0tvj8Vtpoisf2RVXgPbKnURBgJpTfgRQaHrDSH
LlCoivhWTT9C5Cn7heUZcvE6SxWWiZvo+DSVPGXi+alsk/Yy/M/RdmqxCtp+7chOdPyn790vYzZY
uDkyyBk87Usk8M8jOc2iD2pZZ3Bb+w3oL1qeHFW0v9X6QTNyyfiRMD5D3YhxEJ7zXAQZpvdxdRqZ
iLbFJ2zG4J+3u4ZCg7Q2ll2R/6cPBlB/nON6kd+TH1DzmSstrFoqOP9l3+a1zfI5VY8lOfSdrjbt
ZUN4tWedDB9/bkfu4q305bTHth06GJT6hKXnY8pN9KrLRvwQKvhDO802O+9QON8p4kzxQCuvDn8E
vkwXVzGqMUOT+fTSTexzqtiZt951+5uChGPGMT2GgpKAVJlpnS9bxMRYTe7tUSHD17N7Nj9br5Bv
/8EG5MnXQA9341+QOGLRX4RzrPZFTjXsQVMGNGhlAj3eis9nv9wQbIvmiT7KtyjZ/9QWearQWBSy
62jR3oU/n2l39qgGG0HENlzRx9LCDj76O6RF49a+ZX8jQGNSMNMzmWJkOvx2+Exop9sVDd0816lI
AApalDRy2NpEuCF5Rl5HqBneVDkDKL8Ga9GFyzF9f+adtzmRm4BcF2sr0sbqWF6tNElhkH6x6tAC
q1mFYeI45l2Rvp7wjTdb9aMMgPdhfr3OJmvc5m1U8HyrhoUB0MhlZfC3eYAK4SwEGGCswGifeB1q
QtxKqoxMeVmu/reACB/5wYHmuQ3YOQAk6+sTMBf/7+BY1nKK1RV8Mu0qtR8VwXBOuxqajtSa5KEU
F11ig6M3p3U4il7gmE3sds98rfnBir0pfR9ollB6wMZJe2LsBpmSNMlLJPTMY4cojU8bcyoUT1aJ
elQaotpHkozg42OzjOIl6uAAqGMPQeQVxN6Lk20aTCZxSHxry10tFtPGHwlWT1w6eR5vuUFfeyIG
HfdV7lYiTXm8idcT+sovFoLVxU5EP++FJ06fn0adcS9t9pM7ov3PHm9H8i3Y26L936yWs6GlMLvt
Mvx1KrgNoMAZmAnJCEEmzKuCBzqv2ZwP9z7VvXntdg4IXvgTDk/HMsehe/MmzCtJud9/Fm7pS4GI
3I4fbyRqsKkMlls0286z2mAnnXnHRJ4s4fNJ6LlJJXZkHBzA6AMKo7UE8t7WEIHnLLedTQGfhgB3
bb6VVNXLuJh6qaQCRgSfvvckzWs1/Ln4OJxB1msUIJMZ80FHEth8CnQJF7zrbJpmN5IKdmkKBkUE
4yx7u8Ukji2IpvXe3CQlLlnBVQWJjsuGPB4+797/21FZfIiluMdgQNKpQsTa+/YjNGfBkX/GKTT5
w+lLyS4RSvrbr1sEhz4WbZHkhcxK9wuATGfsyoeuQTM5yQScnI+1cgkH9qhsbczxT63Cq2EuOMc2
nprtaQnlmd39atEfmTikM0+SIP9YKoZ3lYicTD1fWOzsQiHk4NaKiX7VdkIYiegA8aYbe5M7WgNh
n+JJn57tTIrgmO4NiTvsWf/aoYXtNY6jGUL99oSb+QkY8NlUHeLiWX7FCOjeYwm72VWomvsz06NY
dLjlRtxt9wVMUBzOOzrLsmGEUbLIh24o4suPUahnwPlYv3VNG4/ZB+xcsAzmfflxhg7Vr6YxPq2b
LtVKATx11PyvkLlaDmcLbwMp2eByZj66+8aOeFuCAC4PtI8iHy20bTN/3Vzok8bllv3QW9sMt4K8
EerT6vOJy6cM5My3oYzTvD6CQU2JpZUeKvu/GlMrYNE4l3pwc2T0sQma4moS3yJj4DVYX2a0BdiC
sBR+xCWjfVZuKbYcRujZrJDdT6K4ySIGTG4pv6py4PQhtZ2xY8q/KWX47XlVpjXozTxFQ7X9JTXG
8N2MhVfKs5FaDg/RR6GVOS0yag8N71byNWi3thoTlW9gnu6kkrDtDBQiL6upwBVy8gLaptsnf/jy
mNu+zjqVMneuGgg5qYs0xgqUA2ry+3acLK4bmturHs1bSB/h+DIY+UJVxchB3IT3FIThw3tN73h0
cShsEPXsXfqSH0/lcUMJhN3GTvYXOmT5mUWyT5L1gLgB3EGUofCdkxucON+UnStRUq5hXJtCp5ct
LEm49CfbPj9SnnTrkg8+ABV7TUPtaZErY+Q4E6C3RcMbrbnyEe50atHB3trx5TTuCIdlRTqeTbXJ
2bSAAGtZxF+7TWGELV3PmroQMbRIV+LA+KYJE6DbCQlMAhDif+7yt2OruwSTL1K+g/wAyN/xK/Mn
UpbSVhje5e4olFKNH2Z3UlkkCoufk1wDOI1NMk6Fe7ERQ4VPZgnVAPjTg70L8A133n2KicpJqOZ4
x54fnNDoI1uW6DpyISI4/Fxx1jfZD5SiyCzDstdZhiRlOEER5y/TKLqV1pkQ9qrUBK53mJeKHNF5
DDrpoYnFzT887JqPTkcZpZzB4axE03XU7TqtsP2Q1IKtYDTGTkgiWMQ4cl2deHk87Sx3H5DBUAM6
qdRQamZzkB0CB9C7oyh2ShGPTWnZUN5CY6v2WRYS5C/hwllXM3ZBJ8V0MgmkTS3dJbU6YK6qexJ5
Dw0xysdqz48gYYi9xgNlEhgR8JCSjySrYfwAdL82Ryr4SZo81l/2GnSlxjpZ71yJE6q9c5QcoGRb
cfr1j2hi9QGaWY07eiAfcPXQwdHJZCT4hvykUBLBp6l5ADXrnaWr1LdbwdUMxQ6xreJAG33ACKyG
0wQPog9Df1wi0nWX5sqzL7YqE4ue0jL+mGPP2DwrEudREF11Nd69ivkVKCkbjIwSUJGhbh5SsbjI
rK6aNbDim+9HOQ6KqesCTOWXKRtQxS+MtNM2fZnJWhMWUN4ZTMvjnGFTBh49XP2RGZn/tJzZgrOH
+XbfObWM9NCBIhxb3gsXXiu0j/D5CkZl0I72AqHvBwgRNT7GUhB63Sh6NIzL3cdgsNjVNKy0uF8t
PAy6Af++8Drxtseyacf5xkB6ThMt16mYTpBXhGii2fbg9UQodY2n4uJ0PhHC0Bf7frEQMtNDm49P
TS/PD32CWQjns3cUDhVYDXPj4N1WLVpXY8B3pk7qOCVBSWLK9IT+1OV3N/z67LSmpjVrwRAL7Gr4
D9fMmCGUq4C7rHljAXytMa3OYZTJnjWUK8hGxKdv4Zxdy3vV+68nBDFNAo3P246BWFtVBDNEX9ab
NTdJYSGxhgnQl1PFah33MrlrzaxgouTIXSx4tYz7pNQIjSZxvb+tzoG06q3nSZC6qAOTtVnkAZ7g
njMTUb+hAqQJsCXY5u1C5tir5RJS169XVtPuKgggeNvaOiTwR1eiYDwuVSoovtcYNdx7AfkHJqSJ
nwkI2aizgxmMqpkWlsrwCNUTEpMCuI5HTyHzOfBtgCXD7rsgirXqZW6hgyz5QnM+/N+vPjbW2yE8
QkUeAYhRSuiTSuuKkrnSEjtEkSvOfzCT1i6LiU9f9SbJXfYzyZuIEQCuXFHqfzEmktfQNNlDZ1S1
TMGc73m1lelTBG3KOCtM+OdJiW3tM4tB+UO+s5LBr7PPHfCPIQ1N8rd/7cAGC+ndUo8whVSle1kI
hcaEhKbm3SpWqbAQiqcSkG4r1drPqaiUGqX46BtZqiS3wKgQtHf64wykgWovdEBkI7ClydIfR4dE
OIl5l3C/QhL6L2bmwc2vM1TxTNQIb5LtHOSUjptbNImeC8uKnaeRLThwmA1xJQr5DnvWGjsAtAJv
VoT2tk8QFpLsYWzbCLE3rOeA1JfCzzCzkXKvqGia6Jk4Y3mpygo5tePAhvxsTrVQL2RW78bdmF7U
BRa7IPTp66flU4H33WeIS1T0zmh/Td6ir0LvRX7yierHHvPrWmfz4/YP+JsbcpXoaPx5Sd5Zx4r/
8puLOLOWY1YJg6Xmbx/81YLJAbmgWKkIWKUhiah0uYlUkemrZZgR6k5WKtk5oRgiu74fJiR5hUnK
p9w6JmudaE3UfxZ9CLLSw1HwSyGS0wRG4ep4+DHwxz1ibz7mBxkepfnaMGDiIW49FX72r6uPVwCy
YvEcEJaWMV3mmbbXsA/OJRT0Ok9ev9JtxwgUzSIg0aMF4/98xmm+GH6ZmV4sdIicbLgPDqHzEYjI
uzcUeQnb6eYUwZpvyrsGnGC6MbfX/Gmpi0sgPnIwfa7TG4xh1GE0MVI+85jnEn45CERQKpow27Ds
K3M7nRPm9nX4VhIac5Vww4O49mxcVa0LyrsPwzKGlZIsZRrQYGlxMIRqI5l2ZZetBEyn9O4G7KO8
+jZwvzoCMz5W5nZOHuzoPE+i2G7/6iM/0pwfBZpLG4a9mrUGfdtrdxHCsiYjgWluuweH7Cm5Po11
SCLSawWqwgRJDRQO4QQmLwn9E8vnpDIDrhZXLzV725gvkZxuiMHOlqknOz7COR9GFgrkeEsljm6l
S3+M2y6wRrNKVDCkvu4c0uPpGa3jNOyR/zx5epGVSoOwQyJwkokkyi/+GLEj38Grxv2k5I7KHxwm
5XEzbIaY3q/gDvV4xUQpM37BvsZwuZjwAyjxc+nTaEZRxfHLVbMqtT8bowPI3FPplv8m9fongsDE
+NDMA9YvuRHBnD7dQIQIxR4H0M+tEf+Qxd3fEklYjHuIUwqgNJB9aP59qyPvmOMr7sH84kEnKwQH
3DJ0K+pAubtfl6w2EH8Didra3Mta9JDTV0uTnfvbrS81WL9aJJY+qfYDMnTDUN0yZL18kNLQIPnr
L9LR+Dbg8psOOhyPjn0Eg6Ts+3Pj8/x0EhKB10+t+JaQcRLR0Nkg9gbr2O4y00mEiPe63Z2IK/G4
VcABmVMpiQxML/Wq5MGX5gOmI7R91c+8lHXO4OMlQja0THlj2dUoQcwV6oiKIMix4EqYUOFdcho2
MGN5Cu0QB4P+nTq4I3b9lJIsvAF+m8PeYwCiXAymwYRgBhtPSFc1zFFwtXdno1IqE4ejJQC9bBm4
nraq7QkRo6NZ37kS6AKLtLSvviIbQgfg8q/lEJH97YudU+Qfzv02Qg/xXQ6ROjZ0pqfmW/rrbwE2
ZqetoObkrV4F7f4FMB6g09/vyzu5PA0AYQzxsnuIUFBVppseetGHXyOQfba2XjbOE9kJo4OtIqMs
siWMuCWlMXfGURaymq5cvoVVgui5ehPfxqs9AeL2eIoQ2YEHqKwOcsrBOzygXGZV4Io+5h7ldu8m
FNz1YRdXepc57Nok3NrgzSG20jzUlJrrvcEysbNwUyviT1DmukaTbNlyg5HR3KDexhQg6pFvLSk2
ujC6/yino4hyM+rsCSMFNpJNCv/tZsKM/wgeBntqCUy4c0Qqzplc1VxdSr4cSA9e+CCAhVRNPRXZ
rMJ7IkVVzfhaYupqbHBsctTT9PYOyyesst25b+fKtcAmXjcr97UFnXgZWSvE4VoyZW6KkSvER3x8
iT91OTx3gQosxaNQ0ddohoGMvvChUNa43ZQUM1qXegP97ftI48bx7WPSnBp+Biq34CHDEvS6RxSM
fEUjcDkkZ77xym3x3wIoiqZOQMkFDOjtkrMfIATIN9H2tmx398iscKWenQdII/HsUqf3uO1auq7A
6G03u2yW6ijitChE3SObVG3l/ojyTBkCiVEnFXBf62e+c03P+Q2x/bjwhnnX8kZItUxEL001+ag9
Qc0mYXbfeBufNXqKftkYAjeKE1gEhqVSLKNhiAzR4EhrGwylhB5zP24uN0XGHZudFhTOsAQ7rJx7
mVzn869c0L697t0pNnJRtdaTMtrrAEG+N3O6dSI4ARMSSCsT2RTsWMcBbRg81a+m2n2Af7oQTku+
GPDLR9Mm4gP9vnCohBrpIfJ15m78owVCIJUmSRT53u2Tza+0zEOs9rdsZdaN5cdeDfau3f1eiFvo
U2qNDt0wrkLnU87eB5Wd5QNlTYMfAACwIDgDrnrAqvq90AhND5pWs53qkdcJM16qmz9fpQgyQMys
D8MkBhjZ7DvkJXXB2JU01WaogmTfiuDqFFn6AdxjRtGKB/FVDi5nYW+M4174NyeiDkKq+xMXRXAE
2Q/WhR5Bdbn5JrZsOU40Xh5qDQjdSNJ36AG/gO8TVw+pNHRVTJKaiKAafiDyMEBAND79E//MEJs/
dnQJeiBdKx9PDI3U+hlahgQZqAKQ3d3s9p7YyBrsN8A4AKxfew+7oentND3zdnIOqi9sg46RWiwx
rh0+1DY6S/XxXQCP7iJZk3N5XUDXhk9OH+SoCgjZ1ijAyXjem4okkeew/Iv8D+I8pKlbfm8za4Ly
YcRUEmateHNVU9j2n14/jRJ3RalIuYfltH7/iMD6rczN63h7Ysl2JUWjyCxClzwLW/xYHTpeJEwp
YPRSWCqxCUHQASj8P7KzlHWRTXIf9D2UShgUX5GrxhAT9VcYuz2NTaGUP4egX9zeBbNaSXeEKqBV
hiGNkpnxCkF/tiiKd2cNRoMlkW1bAjJKwx5fn0UjZGL84sfbTejdT0ZQaIdIvYlcVWClH75AGyXN
jd67Gkg7mUgTI+Y/8O7bosyF5fh1jjFvihRAFqOkrqhegdotzYrTuL7v5EoFwKyjt00AVD6K7z3O
dK32z7wH2dzzUX5Boib+HxBg9U+rnuKkYVXEVsbDG6cMOoULj6qWn/lwBZGbPjA4zPLRoodzlhVM
fDopX6/C4g4j6APDx/JBrR8GfSe8hT4Bo138ksDtINTQgdjBJann1ILI0h1gewFYuWCEDjj9fH69
kEDGl/FMmNylLDmvTq2iiFasiXZMSOwH8LVC0nRzjPT1bPeY5W5JnHE5ug7PhfvEM9FUWs+UAcKM
QnqLp9xATcFv180l9DTjC1gPU6CJUPhwAe7k9movQSPLlHDWtdyVirTxHFIPkx4f+vZqA/xEfyIR
skrx0txRf/dCfDsbZ32sT4Q0eqxi5dkDI/ily21PPD4gVXL/H4gxghj3iN5Gwj3euKa0ussIdTnw
4brDjmXvZrms5Rr4Hdt5JuIgyd5InAOrBRCpDz5zCEgBGOgcgYEar1aTEvQmNrRDHx5Ktzw4njTY
fS4Rcpj8CWDkMvp/Ur17AEUBNysAJqeXbuoZ6rBz1fEXED5vvsoVd5Y4S8Aux09mttYo6Ep+x0A1
SefM8fBSZysphJk70nQXrS5qvOK4z6Drw8U8CPW/Oi0UCb+oCt+y8Oye01vKbtAemAi6IJs+GkPy
IptY6Nx3nwVLEndAOyNgMf8kVS3+qJ6j8kwZa5rFbWRlXBZWFFAB1/7n2yeOMSEkmecSkmVCpbva
+vHiqUb7qQv/XYcpdOje2LY3LJrwsm2GM+dxrI0AxUgCpexC2xkvX0KDm/817X2abiVoyt4Gzbms
8k0NsrbUYHgRRD4cwjSXOxtk4Hz/fpckrav2RlFX7gtRWYNhwOn9SzyJmkT2woBQDqhMzseCP1Hi
obsnKcvD+RttFTe0ontJTIvoduRVZ0gjRSPXrh2c4zXa3cLOtXLZC2x4aPwK5VblQ9d2bjApN+2N
OEDpXaNt7HbXQQVmCXSVHDoMgiCokIrgKw2YglRp9+iGfkC8ckeCtbXBTtOb05odGIc9/eNK5u20
x+2O2Vd04KDePuaMNgE5+klBP6uFtvR1Qg7xZLEkIMs6+t064MIZMdpKWS1Ef5JtvWm5mXW0X148
53Y2SozeSvDPoMCFF3+erA90ok2cxPLlm39ESvNDz4o4Av1V9dR0pdwS9A4D2E9x9hEIL0KHinpb
gGpnn+AOEtIe6CzoOLKNeNhiUO2oG0lHnW6l0gCPBEb+52wHgQm5qNpwr0ixbW/BglMWg3ODgtTv
wR60pZPOELKTjvilZY6PPcg5gQ3E7Q8+IBZlYCW77zQQKFKmSVYvZcptUWLVACacYcR6pYIWFQwR
5Wm1xp2NN6pnnXrA6JOLDytWDAE3en7LP/iYw1oZaODPFNK0EL983iumdQu4muLAXubZVlISqYrY
Mq8Hkrf411Nrmm03C7qkk2ZWLMAcKiE51HYVSwSagYyrx9bE3Ppe2W5QRrKHo914HIHz04AzIJxx
q/l2vAKLdf/0IIj0831TcprJuPPf7LQ67WTv2IoOte9C2ou1Nc1k3uYYVib4X0DjucZ2SXb9mC9s
58FqwAJnOLQ+XOflEWwqtAxkfVWrmi6nbRgIsuBJiBrbjEn3t+gdOVzp3mcGrKsIPcW/ST/DnxTF
8ZH6gzKjTOV4+f8m96+FK2hra16dmx1+supqCRn4aIWCTjI1Rvem7FJyFSIIahVL2BZrcdR8XA0l
B7aOIgnB4t7aFOFaEeIE/DuCf3hoS4pDYbfQbCiyE93zy7v5lTtBZKt4Qsh6/2jTI2gUWm9R0jWb
CGaPbns4eBhF3mDLTOAs7rTN/H/r5qRMDaf/hpUZ9fLWjUNcYYcMQFZQW0JlNPeVH4IqaQ00XVYC
9Zc5cCOJZ2UJ5qR1M/zise+x/b+4pu8mlaWVizkxvh8NNJyL6CXWX/mwjhnIjodB5oQE0z0yU2Yh
WlfK1fh98tj9WdsXEXyIzr5+x4nthzHryGphLn/Io6EnQnYoyOEnYVSiTAWHApJxzBtEJz53PzK+
eng0hXG0SNF7WFbxLbLkiL4ro7CX3ptDWZhesh8sA4V2Q6RCyJ/fUoUP6+IrfaKdTVuK4RNPOq52
HRKfE3GF4aCHHgTwP00XKy9fyM/SVo5tr72t3RfHCo5iivCbRkC/qmEDu5Qu8EmjIuxZQYXcsAfr
Og0W091HuWx171bgMvlDqr3ZSCeKS4iXCIOEm7P2Laun/DxOraMFOqYF/txvXmHl4+C3lg9WD+iE
0FrEQ9ggmzdMj/sgD1SlyU2WpSlM737AINwZNWe6D931ciG/kkRl0y8TgKDpzwgR7Mkg7x4nfUG3
zMFpCfN655I6fCskeIzIfcJxPSauBbK8RYZeBLLZGdRUL3DKf2wl/0ircwa9raFMCS8yxPRZ648w
L+5OlOgT5oxJQOxe6Rc0wjlVhyYqCZq3CFwwbFs40i01y6c72++Xb12jyo3NVTutuSBUJYJNn2hF
zkc90XH4lKQt9M0sKqOscdmdP9wnJZOBxKVBTgSA/D+cYbR6dzJDPuRw4Mk3MVnTM6cfzPG+mopR
sdmXd2R/vEwxgIhUJxKutJoTXZSnXHla0ybHl3WULbNUkVyp0r5fRQ1wcoXSp+2x86kcZBZDbswE
v0rLyRX9Knt3O30W++wGhjAYdMy7FsnD2Z6XddkxtMX7Z+R44ZJs5RaZ1/AxzmszB6W7POf7vXOV
51fJqusciWOlelA0TbK/iD7KMac+0p3fBU1KW2Nysq1v5YzVuOTbFRM27xS0+nNrrkbprTSRfXqO
0yI5eIMwtKLA691dUgPkUoLzfWAYHGvTO20MuNF5+mncX3C5gJ9vN9+yRqBMZa5tqr9a1rrzcPEf
iNEMetwNl3J3NF8D5F0faZGGhaREAgek6HccVnZJNVd8bGCGcYfYv0engjucujT97Um8Z3a/Y9w5
j5VSi5zhk8FuieGXukuPNx3mUKW1cf1wFddBp8rLiSb1FPVUunhRvR7Wc0hrKLFJadMmBQ626lhJ
cz66+96CuH8ysWkczZkZFL0LnH1mC8wGfCICGlYJBujH6nc/cH7FvdqhUprD0rIxxGcLgmPq08ja
NhQicfH7yUL5NoQt039PKb2fTm9PZjxk43Y+vcva+cGNpL0cLCHaoWXeG35liaQU7GaMJNGzEepd
GGoNgy21nJ2NvRHvaMNfSaVp8dmM3kBz5ulTV66d/4SMFbhPGWCvMuuWt3UDopPzyBsA7Ut6kdZ8
cftWD6QkkT/hEhBAdMXxavM3phcbVNxdEva+PzSNt3h35mv7+HqjLVDKSDd92luBIh1JCgttrVEt
8Y6valqOtLNgdOk21CGhsQqeWxwhUXeVR1AaJ1zMfxYYARS7Cvqxco3UsxTA8DiobxxyEuT1MHs5
iDfJuOOtet07ATfVM6yWPXPoOrQ2hpokU88A0N2zw2P9OSSJpgKmCxfxASeGUWeiJAJWYTvHmu+J
1weOtXKVO0nzopTjHWrKXtMs9iLD55/a0yGj/4JJWFkSLozsxAWTpAvsDaBCQV7yzSkY0SmUTi7N
UNwbEn/3HHUj89zL0aep6zf3pFMLdpNW24GiOu6h5dS3DFDweXt3N7iZv5TOcXKRcJBb5Fc208e8
ClKaKHTzeLRnUSXfaQJeIEs+z72NE8sHqxxA6mR9wihPd9mcIYTJUbaVoIwy8n6qjDqDvxz8vrxB
dBuJ0ZlyVDG9kgpC5uC8t/RzecNtK3JsUxlf1DuIQxDaLGBmNPf3hXDoHaC9wXrUeqeXB3UifzpI
ayMwb7XQrsr9WAIerQrmfDV7rcCCTu0bjnRUSAryZFFrmja6MT4sLEEJHbtuTfQiJd5ILI8qAyEw
Ic6PXsmmxDpFXitrGDRQDEur9pknLyW4Edn0Q7QwgU8iePfYhj90vcWG02ABzxLEPxxkHdJM/JMw
y8WTe9rnGfVfo2EPecCfCbOxpAX/2cv2ivJZeECfpRA4MetIzcDbcLiXt904dTLWoMSb4soXL0yH
BsZXXeH2XuhAxAW79UNAQgiD58aEC7CEf+jUY6/GrBB4JY76qScMXIjHhoPTXJFH/WoeVhlNw+Dn
dByKiQop60Cdbh8ecQ3RASCXov3DRkQS4i5IfIafp6iYQlOWuyR2xgWx/ygJdBmRtbWXwWBMy456
bhnKt/gIBsPoCCvoLMWR8PWnVgj2yQK1ozukP3aHyMCuVlHPlPArOLQ34riqpUy2oJ8DFWsddZFn
ROJa09yWjb6q2eTh35OQCOfObt2hHrVIH5FZRWYsBbsJIEl1+J3TcUtHyigKmD7t9jCDohI4BpnD
2nMqdfZ+4lX3o+S+BtlxsBCwZ2ArO/9m0hIGhFm3eZ0V48kvQTTr8F/PafFjtSha2V82pgCqQnjK
Vva4c+1kwg7lSyOqhA/JKI+t+fYaTvQzy7qiqA+GcFrqcdd8JFXjmNwI9oZfJ1I7rhlDodOfkquT
RrtBmyfgpEQg8PhjPujXT4/50IONFGTd/Wr4Pt0CYfaQLlOemPVZ9nZA+Tvl8DHuk91YaY+OFF3j
u/rDvM2xtL7u6qyLlEhhZGOw1xPobwPMWSo4Pxn2BkezsNve157r7TNMTUjuMN3aE0WqdzBq06ag
MQ586x3zjd1NpjdY3ShXgFfH69b++dx71EDb+6//gdVrxi/rHU76eDH84uMy7uBseVhOofLVVw0U
Dj3CLyrl7aZmNKg6RZLN0O2trg6Ghdv389ZKuh6rp61eILtRwqaBAd5AKsWI8oAp0iF6Gf0uLGsE
o6XFLczsC5EKktghrirVhhUkvgfnjID8l13c1Zw3t0N9prYfI1CL/pKJsAXLpNfcW1Tgd3Qe/6KX
UIziNuoI8KaphAkN6rO06nOAeCqXm7GUgwbiXjqOqOeJzfdYspRcdXdDvxz5mUaR6dKP2S2gcRTF
VPfu71LqjZukFNXm8koFl2aJksaRSSbouO3Nabzvcj+u37BdCioxo7xOq072bCRziYTUumF6RYb8
FD9wU1MSgQJHefnXdVu20RWseABqhcDOlXZATvm01D/UkxVuUjfT40Z2CoaTDLLK6PuiwZKq2t/2
WL4k//s+kgpNyuz07VgSUp3HtY6tl7f+nfQRyTYiRrr6D+kmUMpdT9CX2n6r20WqdR1XXISY/kG3
zyAzoilhUMNlAnX8rU+rTNYGwH5L+YPmPvZzV3boAC629ZTkL9cUsntYTpwH7/48nCab0bYCIH6c
3pD6x/n9Xa7iJWVilCes5vpiCtNsqcvHCf/ku+qZ7J1NeQS+r8rE0Yz3m3DGz0V1ZgjL1rycKSTK
cepnsB9I4VZKGTOd6C7QL8ux+mOrX7iDHQkXI5oeZ+/Npw9+/O4Fyb8iZTnE19t/l1EnxBAh4OhS
Rvrt6Y4ug3PTgBlYOATYiBIi0yv92c30iWd6HLvCA/M9X+qBIsVX1tTRlYoRzDK546gmxOfJS8lu
ggHWsJl7dQrpL6nrLZfRrd/3T7YDgyhBc58MKOhmNMp0TTAw0lFTZrpgS21lBk3Rwvb4P/6lAZcc
Z+tb9aNcPsM4KbB2SqaFW7Tk6gn1wnv/olFgd+/kmt3f9eG9NvJJFdxcX+ClCp892WBNJ/kRUcar
XHvridCVYSptmNyoetKxTG3CrzTJcW8at/wILXR4ApXAxBDsJZ1B61KIL8bB9dUkXg7h7VSYspzA
ZFZ4+mdemro9PbK8iyGG+LHs3cxwDbTcVxWMIXOWA4LKxjMpjQzoRPGv4F0wmADpRg1cYwg4fJyl
aNgh6C3Ix9WX7PswwGK/jK5qJ/VpDomqEs6eDRSV++ecZS0QTSQ2qnRAJuk0TjP1Xj5Ifp0Ud/qH
QiXWRr0NmsD5xjnOlE+SM9S0Zgj1vgc9MTnwpvELGtbLCiLxyrP7L4jwpt/0fFJPdqscwKnN7Bfc
zy2coHz2iVfNHELq7YzJ1aK/DmLP22sGyFiLUTeAksFoDE3di2BmBFM4rYqmxkg1MzKI3kHrBXkj
Q2foiut62RvqWB3PBd84nWbNFTEZxe/HNgvWOVfSPojRUhEAxSJlcJ6PFJbDnrnBXZHxcG6er+6O
Bws6tP++esH1O2njx/DUEmfk24TsG1d9AMBxkgg0hi6sn3IEdw0YgfrjaA9MQJ1jZBWnTy6DEHVc
fLd/Hrt+QU0zNtjie9YEyuLRKIbolkWNAwgJi7donOLaaDrddYVxZjaeyLHvSf4sF/WMvIZIGL6X
uWsTBS0vwbGZ/m6seuy5bYcgyrpZiU2+r7ld78yBqP9g5NYaMtj9oQObEM8QjrDX7q4GgwLIyAdg
dUEKJPJrf00UYVKJqE/NHrixMogOGbnM2IFQh6rwvDrB6xOvDHLH+8+xO1my2fzouW6zu5BkppBb
8d8CDqRtma3GQyFOJK8NlSdAHaaPlhgaoPDc4PqXSItoOY+lAle/Zb1k3h+lcZEMaOyUSRB5w1Zl
3ysrLR19nMq9J9CF/EUKoIcV8I+sOFPnEQ/uqJjph+2Ipc4X38qJ/bVv+ihS1IXxb6gpV/F6gQcA
9f7l4u2qxt/US2mbe/ZGLVQX+zJLarr9NL7yfU1k3+wptXT4VXq2szXM9UftkPARcU1KsU3qO6J+
9AWg1CzJpdP2kS7zEa6RrTdOoKtsFgDxNLHMYOmnfgjjZ+MFaN6PkXC4LUWqf28yenLWPvKZ1Vwn
S8V75l616dWgEa/GY1YCy44pkQpgk33gY1NukEhzz640GhjnYXXiVBaIi8Pq0t3qk3UoSdqr7KH4
otUmILVCNMmOVd+HO8+KPymlm50CHELe/ueR3i47aakeek3Lq2XWH727Qioh+8eGTPfOnJc8nNe2
4OcXtdNP3wwZoz9UKX3Os3B7Dhhx/pJdT9rPf5xbn5SYjWHCW1MXouhKFFmghqmZyDU2QkD4vFir
mQm1FqjsXg2P+9dgyK2Gnq3qKrtZRVPsIe41FAQ/l4d5eR11+qhkF8Pv+lPv68cFQrxuc8l2iuej
7VAcgBTPF3e1Bskc7GkiICL/x/+HnUIF++rm4ThfvA5s1/EI+A3JHLBiatgw9/t6ySnTTQSfzz19
FfN2NfN0fd71KIAVGaBHaRHKu6cSvjfZMErFVfBdjTKazBhNYblYlziLB93pRGrreIt6E9fJintx
fp9k9ssHnzXOljGgQHoLIKtiStZ7DvG8YiNy/5ne7Uz0MKFCioMuI2EfO/dhhVu3GfntV/YyekWQ
1hCVsprVdQbawJHDpfon7A6Yq2q2gNHKb+kaeN/bUtgJ1Vn6yK/tFm1PeichV9vkyvzKDwm28SK/
sEVJtTK/y42ZdCyKDgsaRx/ddRMoKUbY6/SHDs1ev9PifuDUe0HI6dGiHfAi98g93jktfHZ6ItVG
9+PPf4FtgwAq1asggWxn49FocBfnt5yKl2ecVciqk7R2ZovD/JCr+7fhfJiU19fM0rySFFSWJsTs
3On5I9WsLDLhTwnpqlF8nqbTloKGmr0Vr0Iwj8Zaj17F1wygNaWZD291Zjr92tug/FH6mzjPgNkd
Vttcqf/6RkG3m9FFBPop0OwxA75OsYn+VsujoiwCPdFu1OnJaT45eUW9mFVX47FgPla9wDW0Q3xM
KGSlUMFBCZ4D08odWJRRl0l1yqaoW52uwVP1DvtYgTfSw/vsSNQTM63cYyTEITDDeQGEyeW34hKH
f6YT4zt/Yo44R4iKdpk1SqEqiIlaslsqQXQNqKYdS97uF/dskVMLoxzOJWVlhSGFX99wE/3DcIKj
jCcFuLCdaTvRQls5p0CRpeRA77kyuezE5wYGIsOdmuh+R8QpphnHft3/g6UP0QHMpz2dZkaAfQWm
3/7ETdmAqcYQzYNmGPzkorLUyGWveSd9zFTsMGGh2gknE3sXngURop9IGUvE3nYcwt6/kWapNTU/
ijGaDoZP4FTK0HvImudETY6cvk2YHTn9W11Va2/BxrSOKq1Jys+n/IBcoKqWaitzPOYroXrAL8iQ
EYUwVLrEvm33+Gnlmf0SPUi/fUeCtDcxCk0BFE8ZQvHh3CH+ToltwdKjd2GJRelJnFy/tHNj0bvr
AhOFvbWoPLv78kTPZEk1VJC753UpU5av4T0EZYiH4fOFv2yyHmOkq4digG2bFWTBH87oV0zkakZP
z289394wVhqQwWHIY/udoywDin3jBlzOPV6dJkTl4jhgpCCOoJ5SFPJpaAlCVQHJ3SCSL6Jyuq/T
k3S/ZL046Epnh8Wjtzz/1tqXLR0OjoEuxbfpa3wpg0AF2/79fNmCj3nPHO+rl9EcIVRgYXdiaZ33
qIEddiWZyI9LV0UPdUBz8HF06Av5wBOJllnnsNH8WHVHQZyKox2VFbEPB3z0o/+P0G2/ouAfIlI+
8r6fCgjqB3XkXrLMPzEp24QNxU1tSCGX6deiWS8Xq7N83pImbHRh6+/uNQ2nthd8i29oGmTZ3Ddj
oO2lWtGtB0FWd7E8G74Myti7WZn0ciCHDUuF/CQp0ccC+JO4aiE3y5A221SzEAWJ4s1gpmvTsGXf
j8j0ZKQ+OPFSD8IWxW5P5KwlWU0BIFronnVcjnkK9EMOCTvSk+kqOiWArmbhc8XYaLGxP18tHEJq
4KiraaV+SVsGkbzeZBwwYffU8NEWVQjZk0wfMN2GIOLGz35wU82FHZufZAa7rJ+uacL5q26H42j3
MjxaDCOY06KedZtToUGZ/B1BMOSjKWZRS0qEje0BJxmU3wu5lzh0LQ/I+go2eNSr3jlAu1YHG5ex
MxQwy8/LsOJnBfOs/Q7TsRSUV6T91pAfNwU7GNWC6D4jvpEjw5rm4MZVKz+mwziVSCTxEFmIBXqA
feJWJ31oXxmkMjkRk7+QJizS6FbLTJr4q4tKQCRWw/J9h8+wzUW4KEiDg75oMza9v6WeG7qwuT4O
9MLDpurEj6mxIUepN26pEge8BgBP576O4S+EinfGcs+aCSe0s5Gewo1O++3Lwtu3mtd+Xk+KDNGo
aoVpuHNBBYUBzV7oCVRMi3xWFyS4gbGaDWyocek0uvFdwzvk54vNEWWUASR+PIa8z+9SSLrS26Av
W0KNw99i4oE8LUTbTRDI82/FrqyPxmS01z8704kQC+fVkMA7nm8armyqbr+4UQ1MHN9667Rs6A3m
ncJNLjxqdyRAKfxdR83FhAij+GNUKZvloeWB5fM5nu+XfQkDAp4I0uY4QyUDjWBoYIi6Myjn5Fw+
1Bx6T+e/2w6qknX7mIoekfAy1RGaa2ji2+AkT90DDVfKBggl2liyi2JEwURjjsz44wU2gIs/PvsC
2DyEBpB5eOOJAfAkht3XHJeBNb4UsEv1qI2Cc6uAvHvOl0EFRRUJ/ROaaNXPYjrzkzTjx6Q6iOGN
2nyXR2rrgWFEALu5XzRR2MlxgwMioS8MGaDtkc/ZVNAz02ctl0vxZaq9n5prlPLssHmFXqJHD0ks
K0YVAnnHVFKdP02Uzmp/jbFGHe3Zr5aNtWMhsYHNNqfbxT3KYRITbeLVMhF64aW8NNzxMpKaqkJY
AHfB2XWe3zzmchaVWvuC1D7anqdL0jTAC7vGtwJynvSLzVlvBg720RqMY6OzGHRYmg5XbfDHbd7r
icWO4Si3SXbSwLtrfWb/5HfrIHljFc8Fs8Z1poxz5AJyU66Tv/W2gAybc3M2j+vmR1ZrDCGCQkrz
GDUyUeCeaB2sWJBEyWX6VIO2b6rEXV+CMIHZHH6K8DFi0gS5t+9ZBAp80xPHuAC/+z73maytLS+X
Bzy3pjK32qOlB04lvv9sYl7HuGSDb0CWcxFHgtcTCsVDlrgW1hqyYH/wxRQOL46voXXuiLmYeKmN
OmqymWLsi5SEG9M6i920QOqg4BzYdD1qtYMbRQJhc6PvAqXgLlaayhLKVZ8Ps/QXAQUO0br1KFkd
mqGb+XpssMamAXQYVW9u3BkFFI5PcqU8yAZH59klQMRCTO7Pir+L8kKHWE8hdH/JFM8TcS4bTYGf
G9pyWRvfSa/aInjRmS1IZMFsUgPDsjVgDxScIkBoTrg5AVFXBreuXq8+UCFugv5xikaoO3MOHirP
WnzDJFCnPMR8AN910nV+8+fEJqnNh/eIoWO0fxAqmGflhlym3M599309WIvPThQu74lLRV7FWG1b
RaIlz5Tcohu/FsOJ2VqLknQ9FIl4FqKfFfw3udvRNgfFLGyB3/8gsdB/YED405mRm7D2GspSPy6y
Pgj7LbO7EJTBMAPFmZBpjItaHI/o+UDmAm+1bKGYsZ5nATdxBhNtAWmdqRbr3JiFNlUS1qAPFtXZ
dG10P5CVAVfCJTYHUvAi8PKvdh38kqRUJ4v18nRvsH76FbcQ99outqzkBpAdoSYetS9OypvO2PDR
3+9PNMwPRRNT+gWC6KHrWrSQCIX5LDRwH5UK4rJpfeGwLWfbyLT3Ts+d8c9/PHIJjoPAAxf3n8+U
m7KTnZcb/EaEuXeghuWMae78rSR5u8XsX3rbG086sM1fbLH9+UjkBjDmbHtNdmHsr4G5rLx4myjS
S6L+frlJKJ1zkubev44WZdwWmbCk/crzKEdRfN0LNUNvuK7NH7VpzZVLro0nFn3YoAwNzFcfILVw
aUz3f1ftx+yWeXBaeDOp/S/PgzoIHhwR+GOc9wKoxDLfxUHqiFJ+asrWqxSFwuTs+I+8jBalF0Mz
HDckIlB/JhePUS+/EUm242Q00nxL/sURPq4woTK/3+JzrYINlrstaM+Mh0DB647nfDHp+dYYVcaJ
q6ui0u4yibIECXyV4vqHdOTcCU2k4zMcVV0oLWwD5Px78Ze62nsRWgeAewp31Ctq9J/3nBlf7EHF
Tvabad0bTCJc7oUh4Bl+/Bvn85fZzdnyQD/1EEUa3JNRx6+6WYiwmvbk21wLfZtxB2GgbngZtZya
Q1EC1OYNf0zwiOCTly/U7DA3Ol7OKIbUsXJaWqr1DPp+ABXdpKEds+Lji0Ods9ElXN0K1m4J3ZBh
YDLTvwSY3rjVmpd/RxSnYxcIXe7HeywvQT5TLKoBGPhYkEQDO0euJ2RfQmdUO4oMQ3j44Kn8EWdU
7lkLujI5hU72t2JhGCFNBkK6uOlBA+9aMLWmXjx8L+tUHPih6fEn9IY1dhIoDPJZPWg84NrnRuBp
en5dkLzoXh20IMaiVg/jRcOP/JKkJXPMTQnXfP6koHVoKJYeG6D73dfsnofCVZoXn6saWAWwdYUY
uZV7zS3xtqPZ29ZjR7BnL91rmUkpJLxwqjGdgJc5DoGWKKn9UJLQEkLLqpQiO30OePipEGyOU1gv
LqI2/2BVVZJnfoaupW84x04oz33dD/tYLjClZqyaxCGV5RIbQgcb+cSpQwiIiGzJtKhNoCM45x4Y
7mm/KMlDQbGyep+gNCGKEa5aghlW1QPF85DmMIQch2u/qBd38pL3uolgi4BqFulfZKyYNjMgm7ZA
vyOFWIy8BRAUHUMUbvXxxkku9DH+HNSVmULgrZxniUqH7rT93OUruEcG5DWeZztXqfZ5BkC3/2+k
VCoicFfXnE4fB0uEr6O4ZoGntCK7/E3fmxhDID1qQL1gFa+wnai10SaqR4vM6Vf4yLPS8STYJ3bH
kNtmNjHCxp/wuKadEB3RIGCyUeYtkYT2qPMxtQse2Cs9JPcixrlLSKSzuG1Q5i+JaGmKLXrAlo8j
aTlfmBtZSR2Ks+R1lCxADUp1QMHliZd6xT4rqENsfAvFKHjUsW2bMtLHZ3YYPLKCeti4xx/MHQfU
/ByYIJPa5IMPsA6j4jSDq+YEzatwv0VhpgkLeCnC3cECrTENeGwQWmpeTVaI79s2XE+yofWHg7LU
hPBkg2RW1OTruKndnr8pYWeUXV2YxRa8QaSY8dyPvm39RSnEOCXJfDCYWK9NNRaa21IRT1dvUsZ7
PC3LN8gVO9gZn/ls8Dd91PMxy6KxHvv9Kms6hglFuplc8L1a0eyCkSoj6IEiOnQdK3/w6XuEpjfX
edH9mz4c3OZ5+gSt8yVatAv4QlazgnrW1I7TLHBshGlR5s+PHHovYl4xhZS8zDepkniIEMlixZrX
8K0Ea3GuHa3keSRHUY8SOj4OF3u07ynn+nQY8B6JDPr9CrBw/NWq4Lp7fNx30uAfHy8ZN607Vayw
wJtCwePpHhbs+qR+WYOZ9mB3uMjbYvTGFpY6vPlZHnG0R2mjVIfTU7rPwPorXoMvVp0jBL16DFJP
ukmKnfoHhZYTayUYakkkLpJWm5o3h5w01OnAjeNJVzpccBR+JXL5A0RAQ9D9A0ExvW5DICKdjWQ2
v/yXFRSIIZ91Ix9jC5PkL+wmNTSdqq55PxnAatupXSyIsPI+mbpy3Pw0SnMnCTZsdVdEAQngf9i0
Dr5ozFhdObGFx/zOuxRXTCPn4iCKn7YTn2hFYWyIJsikXbSVLP9Ropa8cQS9+IJEmMkIo4GJhQzC
sXw+lensSxFGl1tUuOI9XKT1oenlVZavgytCebg4repjfrWAi1d3qPSaXWABczqLguEvybFFnapF
0nHJ9jyqBfMKebuaSZJLTV5XQE0nfdDsxygCmG7Ee8lXZLw96jy5pqL7yLjo0uJzlUWtKjVshceQ
WjcKX8TPCoC96t0LOpNTDJ2q85izjPhgXSRlHoJa9kWNcmimr5Jb1TqqS3Rw0yDbTAA0wKs8hCsV
O3CWF0Pt6hSYMfMsW9ri6gOCWG3Zws2pEKCcNsPWOCNXmpatlX99MHeWgFGugDoeJaUgMqY8m6rF
sA6Qs20XuGSVlC7lkjJekX61D92762j6QKut9UHskV3WUxcDB/YJ+a95aK1vPF+ks3M56EUpfA2F
sp9jG/wDDIpw8H6JuRmxgmsAhJOAdT9KQFmw0SWiHkURDuE7mt5pxeARsS6+eB2GnGLC0bs40oe2
NNQol7rltxvFpNdpnzvnptOuhmYOsbkixxGiw1GzsXTca2xYqxv8cJ7EKLzlWq0dDftJqAxAWuFa
rZ+pPtYJpkWkDkEEVoHamh8Q7H4VmI1Gqano6Ykl3wDlkRqHG8Mg1Ww6EqKqek7IxLkw0wFCbdiH
5eY8eUyPQUr6E0TeFZrmQs6tFNwFkoY+AQvNDpKIxQKuun+YQPej+eulA+hgPQnwPjV6k2oDWN9Q
RlwdXi6cB49oFdoLYvi7n8ohVCNoMziz0kZ13cWL2J6FUDZ7hWmxNJ2zMIsOY0cOCSkFolq/3+fw
UzhPepXn2gJuH5h49Wa3uwCHcoQFiJihvkf6Eu4TH0E+6S2PfU1dP5Yi6aytR5ePL4Slk8xunqHk
kgt77hAg4kROYtkJvthpUvmlPyGwsZ+WBem/htkKHGwHLHdG4Kr/cRYjLSOhxce/sBY8nAsdEn5R
jO/zavNuSeGd3sQWFu0QRfgPRwSykmmFgq+lO3RjoWJks9Kl+fMKR0JiAkhYd8E/Koes+Dm7Ea1Y
Znm0YhBo/jzUo/nUslo9TvomfAsQakCtkNYC3DwUWUlxFERjerflXt4PQDJt+pmGWCt4b6ZOQYor
Z93Bzl5QLCjpKGUj/cBYLnxACHryMoLnc24YFEXW/4eM/nY1vriFLi400HWpk9KSBhzBHlC/VTAk
tIQAIxjexvhiGwFk0zTfGlk6+UUyzfx56rK41PlyqTRuZNEo7dP80TScw3Vd13NrG4tDppDMYMTc
c60C1TkCsJfaX9McSfdkFfRgkQO9EzAcBW9VjiPzTtmVg8kpAz1WUY/Ykz43CsKoYStGgGaYts9F
LsmKUjIgpbwvN2pHNJyqvaNhUPRsQCtecpKLoD65xLyKc9Dnh8EhrrwMbGuvYtzfUuRSlxOenGEg
xZqdPFgC4D1021yYRiXbyh1nFoDLsIft/bY48d8Z3sshuRzUNDb6bcGESLeZwOIbsBZNMhxHotN9
YvG3r3nJ0E75hG3/K9MAlQ1QADKpjCOm+gl10dCEjPyZUAvThX0FzA7AIMjkyWikOrz8P+hOG7wO
toRMBIW8WnLqDGqE6JiCTOiNo6EgC9B/9UKXJ0paIzlaC8jpkr4hKhPv+p8i4WGqBlHswYaXTnLR
e0y3WrlsBrNJHTuABfRvwSOmNJDKi+WkOLbYjn5uCJ8OS+nec9Q2nwV0GjHanVEWHhZAR5AgJ3Gi
7EkUQleXDt2GDkv02aUPSYwUCTBWOVO3ACDT82ntU0yX2OB7by8LW69TcyFn6H8ofMW7E/wYYWdA
tJ5EFnWchhv2S2mH3C3ukJma+iZQgEs4MgPGnxTBiE2eIIoN5XfC9v5d1y4UNhDCrrmUgrsT29iS
piNwshk9XY9LtiGMVWDTQpngI+ePtRXlSifGb5kdOPlpXlJvcYbQOFE80Pzuv+60xg/GJN+mWERq
Cg+IThY0h5/xdDfZw00fs8V3fbWDQsM+tE6AFVE6kPAYJGxiTDEoEMRsr4KgEqsBLDxVhKTjzNr3
5/iKCK4eWO0TTdZ9vXKWiP+om6+exOEO7l1kgEE0aMS0h+kB6C5v2VsXU70+DJ23zmezPcQCXd+a
7FQ7xtrKrpkaen1pMXsIqNxq5ci3RL08NuYVqCiT5xX1b6hrS3cf7b/Ng1NON/VwSBDuilvVDVSe
L7jBJWxltHv6/ZY+rIKGCHbv/5xJ0P7kYhK+Mjmj3li2igRohAOHpHhyqLMNlDxPuLR0StS0fO4A
HhwHgDIFXMjoHuX0K+FVZmrI9uIfYM/UeFWO6bbnP+ZkbuCc9EQB/tOeHlAAnWDQkt4lQkbnfmGT
5KJpdCO/Mm7gMf+riBhqP1E7NPjLQY614TpLiB+ghsp87Ar/QK/EI0FTBvAAtrIDEp1OwXBzTPH/
LNWXsyLNDQ8oY/80yR9go00QUhLnqrBGsajxGocniJ+wPrVIfR7FM+Zi31HjiXqwGH9QIJRvt6Pr
v78h7MxWbQdzde7lEtfg2zJpe/K6d6NuDK06r5/p9RtzDG25C1ohPhujvl7xvYc1creTQygfbiYY
k53sZgEd94YthzXBAzL1t5xFYRl9jScTcPg7kiqaVt5e0vGerfSfV/Iac388vjMeDFBL9vxahZdv
rxzmsUtNGgCeEPi0LiF7JblDZqO2waWC3xuhr4gqtTTA5OAHbBYRjn5t0cYh7tqYzLALp1ymBhIg
bjSzn5gSnxfYoftiRt3SM4jJN2fpbviYTVmRWcbqJRGTF88+edA58vntk3sn44BVNv2XPrrJWqgx
50FJH06acpFUgs3KNTC6EptAlgziMnqsm3S6ovy5Nw29mE2ycegQefS+qaFAeGqlMX2DLRnqjDnw
hWHN3awfgDFKEEZFfTK49Kot1n/GJTc+Yt/NClXeocrNtMZCRNU2VSCg9zOqx5iEjEzCcjVGpGU6
5su1/UsGE4ic5flt6JJ3mfW6MQ86zLMfhr2nrVKTamueHVXSA76YUAyRJ6iM/HINqdIxQOXH6pdy
UQLMIrcfugyw4FDCsP+ZosjcUVz7Q5KuxLLEMrqELWT9rNpXRLe53FFvKM+dzbbo/Nq5E5cM/2d6
khLmjWSqO7C6/MCHSiSkb3Ek+w6rZN5e/JchXaOftJ8IPqm7vSRFxCIxqh0+w+l0pj2Vgplwdn/k
j+q8lIMn0ZmCc1yjCHTkhQSgizLtyAgiDvBeUlG5nJKout+BwfU3xXBxCNPrdS5KCvairXIY0nju
ixES25F8essRZiUZ+yR9hqsQAI8PlE9txKwLiqzxtCCYC0SMMm+LRxiAj46dJnRyhun/PiPE/nXL
w2uKtLqVTgV7VfpzIqlHJ7NPwye2/en311tDQbKfAJ44lCapSA1foddSm3p5pyS6c/JCcPYSS4hj
u3YtoIUUAXbgUj8L8i5y/D7bRu7+u9oC6Oo2dssPKLoEnh3Ec9TRXxLvlkgq45/C9agfBnjVMSCe
atfO0ENA1nvx0yKT+GXlaxyz/ebvWDp46YMS0BrNzF3DsQASHkkFBBxixbfXqKbbG5kIwouU25XK
8lKOZpCOZoExeKtcvXlF+6u8I6OHZcwgN8eQf54JCgEt9jN2ek41dMYO+Z0w690iimSyd8sha5yv
ozfZrxJ32Xw1/vCtmDOCv9qrpwc35h765Sr0CtPSaekfeHGg7GIZl8iDzgpYJcU0AghtkGaw5kgE
JHogPCpfUSmMdMTnwI2s6BrroGfWD+RpFQfxHQ9isosanmTksb2YNQfB/0jWtJT6ByIoDuwTzRSw
henrluRNu4J3hNbHsT0LgzaIgXkwelHiPa3OpexBFeuHatPh4rEuNp/2QmyDSVn53tMvHH479imS
E8Lzh+M29uddtIciJN5b0X9lrgQuM6THYpKv7WhFF1z5TViaZRp+sMTyqfNrWq5vf7kMq3AckegT
TPHsBKD4wXtibeOdwOwIvZanq/JZ3tPxbrDnewnzEWNP9gz2+uyzVexKlZzshdC0nP26790z4GwK
hXHyhzZUzgkxoiisw4LcNlOPs+GY6go4y6339fa2eso8HBK4HohSknrHwhKOG3RpDzl2lWgKzfAk
bK3IFXNPElFUBtmvjFmzJOStjsStiwTFW7f/DS57cq4l53D9MBhGyDGUYrRo2pZ+B7Rv/q7BU0Ue
YweJRFAoi0yBcYso+DOpQAk0P2KsP4X75rii2W+Fo3hdmLcC2gqe2w9SZLL316jJ1bNAMGZA7UIW
T19ux3Sl6MFUNb9SU/xEWjmWMgAcQhVZ8MssiWPl0pUon1+5Rj4RV+Lom6nMZthosCd5QhczRUZH
JsZxsPNv4MVOx9dbOFXN1VNmDOpzCLZQd/38LtkYU/IPy5uRmkfJoDXiapaUeNiveSyjlukd52qW
a6T0Tu0xXoEtQ1f/R39rvLxlhQ6NjrFEceYLaAAQDhqd+hP0HbZGULPs3pBdPFmfYs8KcCfQkP/Q
GePTES7mKz0PyUajd1WipYd60sFPAlTuzVdyHyyXc8nePx4KH4ANi9XgT4iCqJqTucGzjd6sROjU
J74bsTbxEDB2NRVt7L4L21Lcaxmh7I8a0VYP5eeeJroKYAfFXc7A5+cS63+a1iDJmLluWMLKg2Ch
IF0dD+gxIt5b2rkOyinquYm6NKluNPdQ1xjH/40oT45qHojxfj3luqfJD7n95BXfeQBIn2BJLFJS
Uykpywp/1yMCojEyRy1MK9sIl/S+s3gKc7eFxhtyYm67WD/lhTPkdvJzHD4HVEhoPVzIRtDUJ2/N
ml4si17MZEp9psYtZ2x7qu5XaNpBfBLF5Vucn6/g3UF2DUdrAhHUr8GVjMhyqpH36DkD4oI4kmvY
U+USiLp8MeWcT9hw7crtNnInMCIy1lWpvtoa/dUKh6tgL8jEzsrWONJIS/JdoByW3f0yL6tfowXt
hRlpYaRQLhTROjvOED+B7OdrPz3seZUWH3dr0Iic6DealFIdhqcjLpimDrVdpoRjcHUuYz/pHQFj
PFWI8/mQT59HjUGc2BSiBjnvtNMXexFhQs4Il/nz/z2j/7lkTIn2X8yiIAEe6XzuBw7TR0VQbr+X
Y7H34Gpzuf7VmBsfH2Bk/WaVpA5UxCGcSfWZB4MLlK3Yfw6ncB4Hgiz9Suo2g/miLN/qDXNjAvl7
Q341a12uRl00+RO1xS6YO89o0Zpat9WQTBcimXU+08s2SDnU9UVRcHFuhc41QGkN2BxuwmGl31JY
BOvRYODwYAV5w316YNUJqCjsJ0OzdcpD/3dOWVr80LNlEbrrseUuN58c2AMrQq9FJoyMn9VBjaXR
VXenUBjGGlQMvqayfZ7vX5tvMLx3nGkX836VXgyXqrx8kqmqqOJ6pMlNiNR4+0qNUljD9oqt0ZY5
tOCNR/05ysZ+Lha6bjomeKJOFEA7KIbyTSka3yY1xUVCmjhIz03YWaUVJAnoUZbbIaV3DpB5v8uZ
nyZtdOruUziUq4cUnXGnuavEsAp0KrKHsmPHNYtTWkXzAv5OdI7ebG76a1kj79f8FTAerH/222Q/
K39plm0vrUhUrSwSNBN85nY0HO3fCoYg1cBWVzG6GlQTdsQHmMwFkUGV5i+oTyKnYdf4KLbzY+KV
spCPvDChqkck6kzIsGBCF003a8gythQ2oh1CfxpAkjiRZMBE4oRx1aElTunKZOnfaRPcDAuoRGm/
1JX81m3yJSuD7aQs01BjP0A5dLvGrsg1P5I3rSA3LdyTrSpsob3ecx122Wmr4ffw4SiVSpa02LiE
4fT5Uu2yiApVFvHXPbI0SJ1iuJY4mZPM/1qPcq/aIl1f98IV1Q/W4NE6Wm4Mofr6UVlF8h25RCEs
l2jR7xEeHUQOT97+O7iUKRWMy/9WVPkNzIn46fQ+oeGBzUYhZI2IgPgZMXymSNrjeJKbYNh80ANC
XXLuGmqytTgbnX9AkHVyAtspSEICmOFtxBlOVmmw7oNZH62vrcXLLuKyGLM0W96fKoAA7S+8h5yf
Oll9s4/SIITClxvLUuOkujkJVEXU1cKP8lMTpSYTiwh4RhJfDJcPWSKPyRYMeWtN848WO0cTA+XV
RXHcroSE246qP3i6yFnjn5H8XmOHjw9MYpoJFr08vnv1LwH9CEe4iF81ahbtjpNd/7RVGycBRWI5
bcYpHE83ZMRCL1V2QE3lcBvD1eXexeHWJ7lzPgr3CwluMdjbl0wvNYKhJnvpXLRR9kKUq2PRZMp5
nS1tXWV71e5pmpKMOspEdKX+XEfRvD8JitiDwodYKxfikjUZzWimUCS1FLZcrUNrNrj4EolMN43F
cUADwmOQH82LvvYoORcU3y5W1XOB8cgE5MHqqjpy5VFL7WcLN12GzvrRb0Fg1LJXSVFx8XYAEz+q
DXob6MEGvJQqNt7HTgpORo25eYTlRb7RKbSa4AcDJf/stIwPpbeqwFzMLw66IxCanqPQGPe180E5
gE+4Hye/jKjhwKAJCWUp5dI5MU+N+Q7MADr7KTh95TyJgPb4mn6LzrICNOugjsbW2umNILXlk1fK
DyjCDxF4t4f81f8TSp2SRyuIoVgkbuBUXvjj8EhaVSn97Kzqsp4uAT3QD2ti9cHYlC0bXr7eI0CT
tRplg+o8FHRo9LegiD+LDTavuQfX9Rj/f/Dtu0bnuMqJbsPpKf7LYx33LEn/6xUd3Vo1fX53yyex
xxF23/2daSd3y+XGGGYUL5XWqG0QR4P2p7IYHbDrVfrbKl8PJ2MhpBiHtty3vOlqgx+JNDSCIP2/
b9Yza3qv/iJgGbDFoSlMESdN2YoAcNzPR1AP4Cg5gr+4gHvxJ7iVh9WctwyBd9IgKHsuIqzTAFs4
N4Yv0ygNZ1T24M1RiN0gOXksiwhAHCc4uROCrR+3onJiyyfjUIO4uuD8mDylopHNTL6DpX5JWLv5
JmrhqWPNHHtURJol9yiNYRAYzVHqI8VhGAmHKPN92W5hIZtLrCl+f/aaBss3gt/FhefIndlJYszH
zWe5KWSFd7IZHmggLsYpqUJZyvRsM+WY3WZYVFncgO8SlA59sqYT+QIYyWU4bS7R7nY1F4ClARmS
xwHIYEjLKafuSvqLAlJtGKyaLGxB/9L2o9PM2zBqyHqa71C1rL6O4VEFseE/8x0USr3nnjNUEMhe
Br3cympsEjy0NHwEXTKjEDF5rsuDNZP43hSygngy+VN3zQyeUKhiY8pgtqPPA9+D6229ss0gzVfW
z/VN8rYOsLH8Xu+hJ0tw8VmIRsDjbDsZAgZ1o47NgnEocVeeQ0mrjpg5c28UOzrgghIitXAQee5x
3fscs01/wRyZJCfD0wSZVVGELt6Wb9EHd0MrMiQ0xrAu/obcg3QtpP/nW4ydHZgTEnQnVPPWIZM0
41w3S8AZy9U6uIaQH2kt3z5ZZvoPo2UuRJWEkua3R8zPTDwDCSwIdYuZxvFaA4w+dU8B1s9ahMSq
+KlEDknSDdvuLAk/S995874BrbYbtXXOSkTmz7vjnBCLsOVypyCVDJf0wzx+9Q8Lfpyd3/fww6vb
F0wWnjV3+KghHQCuuLDxAYNEG+B/vBgYVKCi3j+j16PsIfc841Tpky/SuZGOUH1AEX+Y7lkMU5o/
bR4kU46ZX5wyBVFBxs2J3kLKm3bcZDVI3pYtAiLYhT3f9BiwoSieMSQErBsdQ7frzCp7Gfw0+vFM
OHr8zcwqaVQPhGYXMmUHnCRsLyKFmo75fBddwVTmZ3iClBk7+rymvngNv7mNMchpi/bPRdhaZew9
vZLWb679c+tVASbUyk+S98W3/5l6RQa2HgMdVUU52nE7UwjGrE/Z0J5y0Dg/amx1bHqm4+gg1+nI
gHkuKzj+Pxnx2bq2xHpfQLZFIflTB88mEyKT+MhTZwtqoP/JJzH6NuyXgBHO5LHvY6mSZTAhWyQn
/eHAN3NM/c5GzHFSyqZPXivV7pYImLpx2kuVla1CZp2Nva5NjuQ722FzQ3tMnfCIvj9hImkANXd/
yOnpa8w5hSTBOk0cw/Vjnd/NWBhH8Sq3c+HsdVR+JvPAto+64aveJ9ZNKOA+/kABvpMD11/osNJg
qJouA7UkkCGstgO0lt47PzvaEZIuhdrtsEiX2pJ1BChRc6rm+2+s54qSKXln34ES6nRTQnP/iSjp
gTaCp3c6I6aKSChnMbR/vb1TQ/JsrKQpfhSA8LuEromqbRE4aX+qfvwLZwFPVv7cr2ad9v2gDyM5
k/Vdj6qu8KnPYnaHykfpepHUQEvKmif9WEY+kx+9eebfofSTNoFn4AAMzZZip4/3cNKUbXj7jZXE
KpLHiHrGi48hTGeWdtcSnxqxqJFdMVDzb4N6XSTZnwvi/kMpxOCGqWuqjSAD5aGUuTVRObKoZweK
7mBLBWUhHigytumECmVIyukqbjOZDJv5pz0e1Xhf/gtyrCqpO6GdfrptAoiVHpk3GNEMnPlEwZGf
lcnCZsaiVq/UzZU9N4ex++JrizfShbOQwopGJBHmMQbWSmF9Oa61QvDoLjYpQkN5miE/ecgQ5jDI
XU8y+JwP29fTXTFhDkO32k2uhqt0F/FEm5CRNWtZqYg8+IrQD/Ut6P9VJoNa3JCTlmIwrXKxo6GQ
/6I071wW5ledO9aarzJpZj0Kna3zwvJ88L415zEJ3932wTHC/XeuLS6/gg5PxuXn9kewWW1zU5wa
4kOnWmbBU9hB3KwoXw6Ya+1FvRvBaCv84ncKOoPNxOvnjAcKe6iFB3pEZ9baqJaapz+/49j/9Td1
E3ZDopEMbcFzhkLxK/jhMJAxGKOM0OE49ZodHmaW15HK28MkPC1Oaj7pwUihmHhNw12hY7TWmJv7
hWAg4dtI0HwEs5wgqNnndeF6HYxNcX9Vf3SKr8ynAg4PJX/SOhqXkGWhPs0LfloAulysDclz2c7l
xy8HbL9EGUe9unzdpWgysqxxDtvkkSvKT1NnRLLtG4j1ko2+gEsv6iesBZQqkfzdr0m3JN8OtXIO
/ymAEStWxo2AHwHGSpM0feryPgoHxN+KRUMO4Z+zyc2pqnqd0mQCol4BrpCPjBA6d+vSjf17gvh1
/2lLaU6ZYnZFl7+e/79/AafnJvFTd0SAGPClUqpi+5vbvB5vLEq1m7SM4B0SjXVpiLq0609mqT+K
nyFA+1DpROAAcwtra51NKcYlAgQ4IK0GHHw2Oc7BOFCLuLnHatiY1mgB4N7yxmGmWvXKPh6utul/
eUgi87KpbZOgn3EyxXRGh1xhjH7aQ65slGXY0hKlXd75zYwNGaxeQwXhlIvAQ/ZvLDy6vRgiXDGc
IoPsYr/lZxUeR7hll83PWVD7Icq0kAWbsP1VMGqIwEOviHNsIAIEN6y6j4Y+75Gv0UfZrvin53WY
HAHYAyDrT4ggscnb2ffOFLxRvjLbskuXm4JjPAKKDSjEkJ7GnDX7XYkiE7+Wx1sNe5tSInoYo1Nr
kYy18rcW8ljk2urBeWRF+5OkdC3cjeo6DzSdxpxLIzLLlow04mt5GTaOjtKOupemGx+HN25fhYpZ
hPEIU58PJ2+WNkGhGGIvmsUu/TeO9OIT9t1nP9SZkFP6RroNv94kKjQf56FQX36mApRnQflsQQmx
m1Zt9q9RBrDAjm+f9/On8rvutCQ30VN9W7s/wcQeEw170dD/H4EClcN9U6FLBetxBAES//1QeZIP
qVZnR1YLcnX7bp+R4J2vR7vf3SMVjAlFEh/xXG+g5oSPnGd4zZNVrEvC8IpiIpsMqY/87dXU9l1R
frSZjtZIJuaLcnEQxB62eUs1QV2U/pI6+U+i8ZBFOL3IrTsmHzC5O5f1mdIJxykExFl4uxY7ZzTF
jGUkZigOQxmMttXQKrptgHdIKITlomifztbUpJUNt1egI0RZ+IbnUbmNYKTXD95T+8P1LWX2T/rR
IOIXMejb1Is/b0PSBL53C732R53KvNNSZ/4IK3uWTMkh+ebfBv/PSoEuSNpEX+gm8rzxEoTYHrrY
fC5rHg1VuS7pmiuIO1l7ps5IIVk3H21VAzpNC/9mZTeNhc3VNyqb2KbA5YHUyvi3VVrKfGKN8rPE
oqBgCRp2oLd7hqWH9mGbkpfvpl2ywZgpgn2c9ObWMeX3/f2PqCoot6ij8UV07ga/RnxS5FfR3TKc
snOA1PK5CnGgbJyIYLGZTyMTEwbLLJy9NNR1vXe1Fdpq6akl5Kw3JgtsRGjM0FtQjYZ8bNmDVRx2
okg2xPqbi/B0tAaJ4Yft6/gvdJL8mSalvFDmyyQuoa+BWeCplMbqm2SJ+fPTkUvrcV8NqCdiE21A
sVi1tY6MnySRSRJEIrUMFZK3Ev6eNL8DsipNTxE9x7TAcqXg4VHV6d1fcYC6vmAl6hAcvYNEL9Wr
VlVJ7ZsmKSNHBvR7rJmuMGkLwqjkownKEtv4C0IQWvf9XM9jRXg1HfMwyzB/7JzJHi2UC/FKxBR0
yksnlmTTS2wKV3/8Bssjfwae/mQPtH6Tq2BFZDF4+N0/+xU13DziFPbd6QAOYtFNY2WRsG8TWVWu
Kft/DHLL8DWYV+oot2gSyUS/1zdrDCGS47p5pRf6TRHrqusBhnEzRGXR+VARNZ0WixqNcOYNcKSh
Xuj8xSRid+oG5tr2IE+IPBFl7mgSYyghfMzkkpNqjDtLtWAW5JIY24HAjSn4gy8fJ+raxztfRJip
TWCFrqm8hmu+55xz0alMSHCB5kLMavbyBzyqVI35q7nU8mrSRX8S/WG7ylUKJS0rY0seWHw3glmG
bJToUV8cbLUX/2VFHTkR8RZJ0+D5sHqW/j/IKKsWfLNkBubRBByIGqiw43oMeACEM5Qyazs3HTwt
tALjyLQ1sZYCdRsv0SPfHoaC8+deAiz/B4qB7NZDsrndZ+7EurQbxhHABqVK+oBfZv1oa4dxuRty
TRzm13QHHhrQAo20RYorA30xOloJCY8wjAvlPXa03yd2lXsoIYOwwMnP/3DpfcF/4R4jGcyYS3Gy
8NWIOAYab3uV7E0pix/Lyp0cioEiaM0jTBdKSNEVOtcnxGVtKO02VZ4Nw7ILbGkLJNDoDuGQTpL6
a6bO9BxFxK16bFOervc56yH1ZNEwyhE+XKRfGIVuROfALPfhWxI2sTX2IA2N069bvqthsBFtH8HO
4uYBAXxRYl0c4FmozTldo9zpkp8RTOiOkjFB53YnNgYifI7zkzDpIuZvxW7SwtX2qSSEQsSFUR6u
ZUDsJ9+TUukppAiPCf44Rggrt61SDgsHe8eEVAUvnZ2PBeleEiBLUaEKAzVYVxrP/v+lw4jaTQza
11Iiy/tpS48lGOPC1A91c8JdCrB4LF2iFD9epcpCg/cCgIsT5KuviWeMYUp+0BTCN2zoFrC2LaXM
mZyqzmG6oveonMELXvqV/la/M8wVnjjgNpOij/bX69a8n0tmJS4r3YLb7q8Pt502fhfWrGsY+sKQ
h4kDi4g3J5w+IgxLSNWavfnnWV/JOpGK+SjgAS/jSrJFObaSbSzLoafPfmplZC5YSRekRQX13si+
2cxcjmpB0wC6Z6bynT8MedSS2/xBaS8WtVuzlouvkq+pq0dg9LXBodh1HuILSXiVQyyZfTnIzXnO
gVQjX9jv7IBLwdt7jsE6jDFXZPukRBKPwdY1QWArmhbgWAQRcYuxaedoMH0wQJOHNz1yAzvli/bd
318Z1IzFNQKNE2+9moz+ENZF5nFF4c4VS2Q/xWJfFvCMDgZtDtkIh/OzJtMErPfzz7h25dmAAn8d
3M5rzPd3aWRXAZkzhei6u19Q8TMv8GNhWqVRo9ZMjaKOCaSyAj2B+Snt8JlBjwKXmu9noMs3eODd
wl8C4Q83CarzGp26paP2ipHLgdziNT3YJrx4Aq/cTjiNe7HssPraC17ZJHW+Qzs7eOQJbvadycur
/fdCCoNgb8yOZOJx03hCPGtDEpHJ6l2KXtvWhmq/DCXzHFgmhjQWbNel6hon09EbJaTk+O7eWbLP
qMamXP+JseAGAJrsNY7e4IO6K6tVesews02O9VU+z8DkOa/GV3eF1zW5io7eaSF2ZuwRiuXZIeQj
7IS1cAr49zej2AiWuam6WooAv9w1PkLAkw7x+7hXmGN339S8WAK6oqvRv/4W/TsaHx9v8DAgvK3r
cTA+aWOo0mVlGuHWqrdU2e6fzfGNZ8POJlMcEPiAi3TYsDZnN2KdfS+DITcvP6+sW+g6AfJiY5fT
HU1o+tN11neSOQFcESAvPsNtETP94xcGp7wZud4+x0JI7pgCVprQmvMBYDLwkmWtmzIYE3VfD5YS
AD8l2ABtPGZz2SfPB7cJm5yfo5uTBmcyFSzsdUSfWWB0X6MitKMxDhqbVgnW6eYEv/IgvmhGsXPy
VMVKI8b1qXSzpC2+o/VQRXksI+I043rxP2G1ERm+ZvVm452IwvW/Ormpt+99ckW32o/AqZpoCoQV
xHB8tecuRlHt/6ahYmU7gNGFsJpycO6cugGDDetmTlmNPx3UynDjH+GFQ1CzWsZdcRB+6AtZksbf
HDubLf30vacRX4S15N//EbsdFpcQ2Xd7kuUhZIc20CvWrPp819gOMtfASURlsSaIR0sl3O+mP73k
8jRta9HGHWsoPxNhEvE6hLuxee20zfBHi+Os+++F0yvH2nCPfLbkW2CVyynlLunR7f93Ta8H0PxC
Vp6bBp7yYbvy6mL7Dm68ou93wESJdISmJI2XLcpWbtfLZDUm0N2gLVPEtdM/ThVv+W8+bByk9OcR
of5S4FCQ55TrDIWxqPm1fcCeoB56XiTtbC0pvY0QA1+XXtHCKOjOxkc2yCbKF186ZooitGLzAiz8
6H/77jiOYQUCOG0OtpiCOnYOb+V/QP3nc+XRHvoo6nt3Y4T076ZU4rLkgC2PwdW9H+7RMZC/Jd9w
HNi8vEdpN8KY7vqbUROwHRkSCGr7olvx2w2VHyPp2UQtI26KKU/ZYH1o161gA/aG+gAR10k/mOWv
uKrmHW07a96xhRDYbFw3oU1791k+O0+nzHid1djNy3oFYKcVM9EBqMZ2IonDxxJSKcuwDVYeKRgX
zGiDJwts/ViFL5YFcxLuXHLTTuULVlQV9xqLpxjBJ24YU2iceRt8HYmPLELmCkrrgiROVwwZGXm6
JmjaYX7+/vLjFA/fUpCnrlB+8pySCouwpzVPgQ1djEqCCE0FyXGpwJVf3ZQ2jVbjq3nadt253tq3
+j5mVAS2tHQZ0H3w0/LAFGVpTUhGyThghanrqt5ustmUptdoGQAqeuKLCpGZnM1qAuK0kRMj4Gjx
x4lAPVGqeH0lye60fvVWwZYyLFaq0r5Zr+zRfCpppPiX/370q4b0RJZ+/WkMCymUt0AteEvPKctf
VmY8Dw1FiZBpdHv3iI4hqRv7AVKisAEjLo6id9myeYeZnD5Wjn9vYHBaD2nlmnVNXHVOfcFvO9Aa
fOefXiTXjJXaCGNxHEJMqwktAla8gT4ijGOfOihEJDCpm/ZvuH3AxRB0jTMilhzlpa0rxBrC0DFL
x9STbkNLVwM3vn6+GENtur5GYzDElaQNDQCuHvigQ4aIgEGziB6eZQagcr1bjsp68KlV5Ioyo8O5
Qay6AoNKmtm99YNfoequy+j9dFq0m8NKY+ejVsbPWJpTZVfCt3Qeyv6ZXvTJuGlxKBTjY20QzVNV
UhzRDYtJ/yDOyKcN60f7DDcRypsYQhMbjapcUbwz7KbVa2NaL5F6Qt73Cuvk
`protect end_protected
