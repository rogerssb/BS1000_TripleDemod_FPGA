

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KHi/M3BTJSmSi8eKDRu6qrIgjp2MN+sO8ExfqFjNoz4nifEO6ThamG/rkDMbSXxMz2F++qwB3LwE
ObyOGYRh6w==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lPvtggTP1o1s0S/BMx9LZQu6i232RIiewKIRL5Opwd4xfKcIB55RnLQh/DfI5un2YDiG5ODrqzBs
53YFw5+qwZkrayznP702MyF0ttPzpcDmL2vac/nTlzjqfFC4j0wySLMr4znjW6VPvs2ZvzlemdKD
3tIxcCeVqWKrCOUSps8=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
aYRS+BKRB5/m4zN6hTZ/AfBWYEU7SU1ObGDxbJxfBxyjGukFkOyFS9IcQxw1Ea7B1mtsWSAuoOkx
j8Ke59/te0OKZnvbsDG0LLD5S7ZuDBHdQKp9j7GuTpWZNWZO49nhj6tRqhlriEp5XZSISNajWrR2
hc8jpvNVTPnbX5s9FnE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
tQGDmfcroz39gXkUVe1PRT2McDBBNCtvLFHrQY9WjwJubYMMcjFTag5Yw7re4rvepYO+r/OJ/9DK
ePsOw5kBOR+8SZP2gVutLV3OAYo1bC3KXcbAB34omDEXujSTdqlJHuS2RLXgyEzkTOWtWb2ex8ta
0Z7IckG6OMpV/2MiQnXPVdCs3Rtzj+p32Jn0Y9MGUqQPtydqC48CssuoTAiDcQNANk10HG5tZT2o
cVLgSC9kaM0j+yKYWK2iNANyk3KqQ8k88WFuzJeBfjkXwUtpIATjQlwJvRawCmaKfIdjqv+PDAP2
u3jtPfaC/UTLWDRMUYBGUokcDsteHHV8HTBgog==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gbPSrvcpZbGRr+8x+sKTlnUUuh+SGrJMWhpyMd6nPLQn7eIDUiAz0N71XlB3mrD8Zo3p/VKWFWY5
WnDov6UMLVGUDRCMkS3BXIChJ0ra4iu1uO5Wc+cWlJty6FIZuCcz2IkBvBejfngcGJUldH3YInks
mh04/8GnG6PVkc5wWeFnqWxk8Yas6e5LvOwCUEgdVS+6/smRqGo1pnNQAMQnR7wJSwtzPTswLZgQ
YzMo3pGFaONzkQFe/WG9+Ptnuktihh/FHDP/6HLw+SpMzK/BwpeBPj4TI39Bl3riyYmwrZt/XGI2
g8RsVCxUTOhu5EEp8NfCRsKCqMyGNfwagr4M9w==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
aff1iZjY/l1xrqAWU30UAh3ovbDS5gl/X39DQ0k7RDR2SWkjQ218HJ2chBMt3lidQZ3OQRI192OF
5kc6to3ojCnXUh7TjVerzpKk22OA2U0nK+KedW4iyi/FTpx3IViMTNftTm/NT7tN7OXYOD0dl+3Y
zsb+a+RgQNOBHrgYgK6YEBKO/iMrZCdjv7bBZ+Mq/VQH7O2iau8gmkj2AvaQBBA3iKWwLf9Vxsap
sLsC/+KiLry3ofDpiQ9psV2WD+N5YjkylQHZEzlnOJ1h8jQw5+NLFRGVKAKNot33U+7pNNtLzelO
YMN+OFM9r1j8f+eRjyGHgataI1ETTztqsGtXtw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74064)
`protect data_block
IRztpW93Noi1cL1MZFuG0f1ElkwLvf2V0i3H7lpzj3yd9BAyPW4Lvd7QSReBMzN6BIelseNo/KWq
2nAXCKx1Adkxv5mDwULHmddxC4MpDqsIcSQrASMv8vypRooZbeB5157+oTjV0EZy3mgPWouj6jKF
/WMW5rDKvbW94/sV9UcHHlFL2duFRhTr8i3FBcm3j8QsqxV5yIVhCRoKxyYtV05AmN84YJjCkwxV
gw+51w7yE94/Q9VRaTWr1ncYYmjSiD93ysNHFc1vcBIrzmiSOnkfLwGjCA3zHD2ES0dZzqmCPImF
CfSGQumXpqBtLLa0ntNlSQY9jSoCbl8rVX9F4aGeQ8jDIH/fm+yw0x/+BR1/rbcCk++MHcmwqfGy
BKj70tX9L9Z4DYj4qzEgHmfkkC6fBFGm8aP/lSf+UlMaqkqKMOKhSiMjfiOTCOvMUshJ8eG6h1Wr
PxjQTS58mk0jhQ1J+1/3HBqzM4zptt6375n458m2N/cGb5s6SzYhklQwodbwu+bFDDletD6gkDGp
GJOsI3QMMapjqpkBzBKFItiOU9s+CJaqqaRgkjQHqw1rqPY+ELn7braAqvJp0dcUge6CNlhVGq54
Dosq3yJ8E2gVER/TR1Y9By7N/9OGbvqHp9blsJ6pwb0b3DbxFfcKbgxmPzCMCo2G6Po0rXf0kQR7
VuwdJL1n7jBb7TzESomG8dt3Pzjz4RIospMXPRSmLd+4snpTWv2JsQS8DY6oK9T5//NJG5STusHK
dkqGuLHAHLlt4ppiLjV11ayzr/328CntxiRgYu4OV4C0h+kyA4u3RCQaDclzpAv1IIOEw/yXU4Hq
3LAQtt4kwz+VkCZHZE+XpfeM5gL3MMZzY0YP8WO24OWuq+gr9Hk4WyXk7z/O/TLn6opf3FsorKjJ
Ak1tBa+uD3269ZGva9SKnzm+8UHCBCTW576zZ41T4OerjWhdudQZZBtEempDD2Ne3JbL1XYkxDs2
MLlShh8URD0APStQ2fsMMmjR9K2dtutE7eeIKad1nDQEqf+V0DuJr8d09T3xkw2kU8yJILdr/AvC
gRr5YEYKN7/tLJHK+7yTcGjqsjEQDJ0cfGMqlM20Ei1H7ZKr0+m9YNIma9+qloswsoSAuCZokPm9
0pUpNMz4oRinnx1++ec6QKqm9uXJhM+rFlXNc/qJFq3S+g86iHSsjFYJpQJTw/op0swkwuxJNlzW
JXAL4Za3egZMs2xStjFFY0+RMlWnbzMooX5uvDBONFkoGVePGFBEKW0JyKwb7NNI4YH+A3x0E39Z
+4RPTLOJ4Pj4beawx5tK34nZwWRTs8PBWxU24gqAsl9u7Mjf+x8w25sxLps91lFBXPQDMEXcoTVD
oF9DKt7v2ggDrZPUsPO3QBKDNBCn+h+Ru69i6awSaqRK4jBsUPmqDhlqc25BrKRWaUAGPNy+zj4u
L1+jzIcLXMZyUZMiPozfZRnV509Sb46hdKZ0Qi/lRwJioZDqG5DPVkX2Ky1WqEptj9IFGqJcPctB
ypMX1oJh5L/WEnh5raQTWyxDNX7FHMubJ9DtVcy9mG2rmjo3MsbwOMSAT49JLKx3C5XgAhjvChxB
QdiqOb8X+Qyr2iNFbiY51uP6//ZlnoOhRMZL+kMRC7cIb993nDf7If/0SVD5o0KYxePT00Uw5T4C
zhOSSbk2g9nZvzdN8wNk6H5oGCkxxAZtTghHFxwr5i4CN1PNMz6gqGSr8zLBvI2BZKr4mgu5G252
Zq9RoY3sMcqjE70F0HLfObjwrj3qP/tIUJr13W3RJt06bck3E224GsiOGdtqiZMLXq7TBWnRNZN9
WMzFuQjm0VwKbtkccN+ohCILyhxPwd7eyK+DluEj96R+okavloC7o2mVNyk+zWgfobATrfxHfnUV
NN1IwpGFUibOuuoFVpN2SIFxHcXAsSgD8xvQ0Gg742aoEdnQegEN+bapb3YZn+EpM56DWaf1Uw2o
eCwdVE26mbsEnmtK5OoaNKWxxp+yNKHh8+4OqYk/kcLWkzfMkh5HqAWGlOVA8qTN+9tt5KV8+HJY
+95wILCUWoePKB0KFK0LbUezL7p6MM8TVjA4m68HxKHUapyh6yxAapHDtSO7LDgZBtxRl3ooHLaQ
LooTqMDZYNvj7lpOTmXZTaisTCgu5QugOYXRkzEsBOLllBtCAQusILh52i483R9funDS1wIf3k6Q
H6os8b8Z6qsxiSfuv8yE66h2sQfpr2oPcYbfIWDH8JpO1fG4MdDCtpfZzVMFk3cxki587+S0+wdA
6NYIt9whus/OY0BXIDeOUfmN+0ONMe41wuawiuLsK1tF07FW5BZ2MYDyYvNQrccqn8oE44FLp2Ki
mUvNnuKQGFaHaz1ScBnII4Ce3ANhAOmnQ5MnxOxr80Y6c+KvptfSVJfRShcobsJzrbWxRrmr8NS/
PfjDnU0XnopKme0x1Aiatv/UbDizsVg/T72TZuZ6Qr0HmTChkGp7ikPtZsvIFJclJ6mYGKzUV8BK
xHukMHYWgerSORjUGp1Voh8quzY3R/CkVxTxrx1Tliuzsw1vxsRgwSXAgteLKf5O1lONWw8wFPtN
RVhuQYq07Y+ZeFdOEHh/+KdWhbrxjCMtiOsj1ZE2zyh/qmo88K3gDmAVKdlamEauBAj1ErycHoyI
8UmtRa8gs1W4AIKbdmmUhHQqFQncobbELcJuFmjB5Zpp5yXtkKEusmd3a1zAhyOmU6LbrlEp04Nt
D1WNTlhyMS7OpS3U+31KuRt88raXpaT0nSkHdJLbIo49nezCjqc2SMvPoeCLhejgdbMVYXqzrhXw
K1tkogMccP6IIQaIFQPKyVXcy7DqukB7sgP9Fgq4HVZhyGOEVhikxLXyyt/1xYSooQRjRPWZDgjY
I+Rv+aGiGWOGYukb/iE11MgMUsj5Wtb7Ff26GssouBCf6mWS6py0X1tXX1TJRScNUBoexzumMy62
NYCGLV2Bw2cQQMa8UEHUTWHG1/Kg+QMDIhD1fJ12tweFu5bubbma8lPw3XFrgBV0oGJDr2ILisZ3
tKsnS/5+LsPcHCoOU22oRabASIH5yNDHpkWC2lJu5lMzpc0vRiudANNNTwMiLt5G/EjU46nCot7m
Fy+IsM4HWu5nqrBbV6zd6xTR9HXqvCCVCr4Va/E863pyFzEZwijqqBf8jom7I4dvuXVAyINSFf83
g8WaaejlL4wEQhuhjNXgm6JH/dplJ6VM3e4fbmSH0xCfGxG5u8OI5Q04rpImJA4Eohy0qROdGbec
9W93JT/KylAmAJT9dMJ4jMDJk8qR1J+nt9xtcRDNXz8B8ZLNU70GrC3TdXrUUm4GyGuFlpEPLW8N
qTDW0/0Iy6Df2ejK/WtEvTv6PspHcHaqHO2m2HUbXpnonRD2VDK0znDZDfcHn/DvFsa61oJKO6e3
drQYOwkjK3Cbfi7izVSm/HW9NtFZQA1GKwUSgFRv1EpWH76PRpXzLTdIcuvfBUUvRsoaoLpl9mOC
XyIAxpEbGNOrJNi+TzB1JPtZGLqlILJFQCf3nSHc00WrkTgofIErykyuOwJHVQ8tR34GklyM6lr7
b6iFSDdZKrVTr1MN6ivVpHEoOVJ8KuHZKasYZZCX3z5UbLcu3IZRHdlWCQG6Sb3XGyZMC6/Qg2NI
DTPr4btgy3txCePV97k4Hhov6TvlxxrDvZh3t3iFHtc4YM+lch05DtVKQwUJfNNoT04ddSJ8dHiL
SdZ4r/hNPmW4YtJ6PxIETO0EVk7YxWpHRqybLgxHYQrnaUcUSO7FApyt7AuOZZCrY7jtSo/Dv9gu
z3ZHwT9yFD6+kebM+TrXByGvu46Og4YOwz6iblD8J9VXIGXhqx+i2UYxjRo4TmveWwQ9kgnPkgnr
It+a7Hy+Bugq/+z9QmBpSHwITW7r1hx7SkTfOhbzZj9M31v+qniNCfcVM4X6KpHtW/9qCZbQacGi
/1kM9fTa1/4Rs0BsqbY/blf+Gc0CQh4JTa7N5Mq0E+dnQGRnzHEHEJp3mWGgfcoK4fbudJZ3jT7J
YESvpsiUu89ljExry2fh5j6jWfNCelLTPLDdVFQi21d8v6lAs9qbgxqDhrLeoeHNT0OoKUqki/MI
VG+6LYVyA2nRwedjwZxhgk4InXTVpsQxDovt9EZ0sLuHG1TU3xLjM9uzpSKh/pp+mm0IO2DWCu7X
Xg9yxbQghJx9CuXRh6R28y9GXfCYcFPgOwQ4u7cFeQ7Oji1j+jyVzdo+jGJ/WCJ3DJvuLS0YFwjz
S5yN9H5KjaiYu5rCAFPG40JRYWobWt6gi1RF7ESN14QJUuYE0/z6VY5DsqsPxe7NCNBZ0HKXiLAG
SUqumHKYzon0F5F2fdYqj+nU/vhRusfNKQwovwdSOX9RMwThnaQqiF1aMMyGaIgwQI9MbF0iiNh9
6oVt0o1Y7pzKVQt60lB6j87jHzAEhjHNFAsezqTcnUcP0z2DLOCu8f8SUiDRvft3SBo3b0DCNyYm
lSRb5G4i1KwIuRi+dycUdx0EKR6atAxFBIRoUPliCnZPN8g6xEyXaDRXafUAyjnwm7SW3yH8w07e
Z4S9CzkE0KAgnLMSmRKrpc05CY1TmAOFCgzKNS5a5pFusoD7NREsaummW3CxCVWKI/PWqnqe6IjE
zNpeH846OqRmOazMpci6DgvGWsiWoHwO+TZ4tutWjJ5n0sdcqmns+mhOjQEwuEs/O/+aVRVbr43X
Vnl87ewlgs9aLMRNBimEgpJGoFplOEqYwGrglXmUYIJgPlS8FJTA1AlzSo7sy7QGfPXq3URP3kUc
XWleljvU9BNCmU8y+ZWoXnu7BX9DnascHRB4/+4gX+NaW6kGgthqaIzvmWJBWg0FcF1mXswq6rDe
Hs+0hJnrbAjP2ZkD7X6qH4e6/5OMtX2c31WovPWYMbLcR+Hy0VW5OITEaFtbrx8B+uUcVVZWM8QV
ImBiUV+xMk08ntRqSmWW06VjV8nForYzK4WCqj7DKgPR1yjVON/JthCpXSlgTWf+29E0SuKLI9/I
28FJX8qruMSkOsFDAPlkpxAwJhPCY+7WUGwy4z1MWYuRNynKLTGmzTeBA/9y5mO88M6sGbzbCsty
k++HxYanwnZv1u99LgtvrqHSXbxpVIys74wc0Pu2HtDNrx6UKowBTzVwMoscOFZu+DLhoPCLZ+E1
8QkaemMsSC5zAlhuIIcfXJPJCfav6+TNUWKFnKtNW6bgQLPBlrlW/yDN8RWNj1v5qRlLRdgs8dIQ
q8QmYizCOVRkhu6NIQufQ4JGegK9lgDGq392uzg1kmrVdx2bvHW5fPAqWIZbJf6DdqOWV4t+glWf
mpU8wcrc6ltmvQByOALS4iFNpUcNztp3un78x0jNqNZJrn+mAN/alUnG7msbPxcKaA8KexBtCA6n
h1gGBxeh1g4DOE0fxoxZPGJhvkaZ5mWEWnqwzfip5f7lZtOnpMxSk8LVMjwefVIUoh2EZrUpEaB8
KEZ02rn2fZTa/r9ggEEIpcoLeB4kS5I9qkyhIe6iwmMOlgncxSHbvqHeQ2vbaJjhhawo5LMfNP79
6M546C//YC/fZIwmm0T925e/iYI12J4OJSzT6ulJteQT3bdkA4UrX2oKHkqZ/wKpNhGj4Gm2VIbj
EcUghUdxHPj6XHQQT1mSmI7KRSB5QIScFwQNKvKETs/Ok+dXNRz5en3eiQJKnNgWeZ0BToOm39yg
k2Pk/w4BBHmmv54rEOxR1/IqvPzWhgnCkWI7TAbGb0/GKtmq4sC4Y+9TCOpc0GQjX9zrz1bW7hZV
y8/45iyR/oh1lhAA522XKHiiTZfM42neq01fHkNu7k5VmrwY9jbGZzdcxCai2e4SYgeciNHi3oFd
rsl1wxCOCA2/6qYXSF9mqb3PwNOl8hBsNNCIjdw6yflCnPzqcMmwJ0Dzc7BIxBeA+XUFhdCmfOzL
g+XnJ0FGj8rJm2+SflnxUtamx7F8BsusOP4vowBkMnzU7J9soJoYFruotYfgEh+eSmLzLfW6FQwm
gdiNqJ8bIpK3qBXYzelW1Qe0C1DxUnXJUXYbs7MsMfxTzsEIJPcVbwfJaglbcBm5l3WbPSI1MMx9
iX4HwCmRD9o555Ppu1Os4DJC8Jo5xXnv4zxkot49GywfQc/1K522TvOusXX3FkT/c8//uqWBwTgf
Cd6mK5A/3C9glAlqpmnC4+9qX3SJTw2OWBVzh7ayWZ8P+0rhCxfR2ZWncCbUEd2IGoEsUTzZ0ljS
K9+Hrl1kkUKrzMQCujATjk5vTeAzqZZBMAVWC11eAPw8DbQ84zaY29va9kwnHU/rkndSxXh2ZLB5
lcHYAMYvmOt2TRAzVnXdeRtdXq2zbSIZeZYtmgfdNmC9chKVrIhNyRtr7uopDLCxSbCQT/DltndD
03N80E3ZZJjRaxnd+q4e0TdRZvJ0XhqMKSG+p+meLCsFEnTanHQoSE81n8AllY2L3xyweDet6Bex
RaObk+HmKxx+UdX3u3fJVPvPo6N1G2GIEEDNihjq2drJsBuJsAtvw0yWZXOU4Ux+gr/woMHi1oAn
YDBhg3lIHgAsBUUXp4DQSXLrR+wVBaC4rWx/0fgXjfWqPInjY8XgoMeuR/iDB8vTJjZOW9XLxnbH
N5MsNIsg6D2CPd6dRL/gljhC0gFeUeds+WYrSuPi3mzbSfOe338GoFY1AGySClzu+mPCZXZuQ/3y
Ob1TSGgdoDhQ2Kudt1s+7YNS3fK2arLCWSQcsVP5rzgsjvkg40z3okx+Fp7Seb1TpOXfyhS2yLV6
0gRjJYs6IeaQ54DfqCE8GQE7pryhImjY53SWax2ppXnPAC0vYAMgCKBO+Gdr9KSxWyimnr0sfhhB
pJiAfs0QbcPN8nqGWsXwEA7O17JlMTvbENX/bXSPg3Uc0/qpj7X5V6CacqHMQ0swbqIFffDVvRZy
NkErg45wi6akeUG0qWQcGYWvDjCSRpFNmvO2m1zjIaQ8kDitwFzwQJLtGwN+OXBHzcLsitX5U2RA
RLyW2jYr7S9pPUt5H2+UpMdY6kAXp/O6+7AyjGpCN7Of8G7puq9dupJfBnTiK0AUhzfnhXEDrjoD
Ia4fatpj/qpylP2rEZ9g7tnLsi9GkemFRJw+tSAfl5sKriTe37O4H5QkXYPSZBkZ43oGLdR9dKx1
C4P0ZQQ/upAQfDl0KiM7PR9kc7RJhmv3yA9gTANyWPqbGwt1UW9X2MfrhzNa4n/Gx8DF4g6J7vFK
KUVjYU8Vf7er9jVjsJDbgBJH7C2PeZ6kNjZHQojuPzK9zHtaJLtxoCcN7yikMtTBrQhO9GlbvvCl
nLKucv1FGRp8wc0zFflhRng2482klh7saBvjIoR0apTc8ALj2mbHO6jcYjoFVZzf+GVRndSXg1aU
nfgL7hNxN0JorxzRQZi2JGCNRGxgjMSFVLtOV+h+XfqPTnzRH6006B0/jXm2pXlN5ya+opTyquFf
sfxi3vm2ef3T+tUOhYqwEzSB+qh/RNOBSGCAl9A1IPA4gxlmiD3tcRWJ7zjUfObTwnJH+ULFnpu9
pl/VeACSs0Bk+w3Ndo4MstLdhw5bIUzYFNWRgn62D15jNmPj2f7COm6LXjX9dXzyaMHp2ujMY7cJ
aPQFL1K0tLn7GVTQDLsuFrytugNy5Uo6WTwYUqq6UU30u1ROkO4QEKaFrNbW9p5NCjLlTN/VWBE+
ZEoV/UTNDAMNU4brnuoor3BU7cdMvX0tf53QRHy0gk+2dCStHnUPfjIlfm0+jrwq0ot8zwD/BzEG
GT9K8tYaGhnRNMkiT2/P2DLrsDBqH/CA3YLsEAIjbNnCGLr2Osih5ueq+XxZkcudYsDnMLT+DDU7
mH4g0JfGyLZvI3K98entDSkrFho/DbEsurVGydkeh6RpuULwSaRMtiQnbSh43I4u6IjRgvEDUfzN
ordaqOV4opO1UMmw9Kx4gSlT17TJDjGvQkFpimCHFOsrh6f6Wtq7pqX+A0ATmp1IGFcNrSDQr0Uk
jWMA44LIKIB0PsgAfms3ajzBeV7YT01E0vjhAIp8HPVhMqEKQoi+VIrFG7CaM7sdBFW8+EuuMa52
vjlwmTj6n5vr/SHdz3F2v41iZyc0OoJap1apEmXVqrmusflDVz4Y9UVerMFOVjAePZ9SSSGpZdbb
aCa1vxPnHU77M7gHHqvnVV3x78a2OjGu8n6sB5DaHsg51YdT/nG926U2XiKS45M9/LO4jwafyiJ5
FmPG5EmqIKmGxN9ZXV76xBNfOMimgqlCy3emftbf5l/IyhMo12CwoGwhlXosqeelAUZwjwUOqZR8
CEXnZUN2tnUn7cZoF/judkfKG/Zpfv6oVpk/BAXNsm/qYacTPh6X+lCT0Za0lHGjnWIMIA9xxsE1
+wM6sdnhOgF5kjWtHJMPdVOW7NoNTCHL2R6zqNoetMOQDhc1F+Zcbq9PSDQn+PvHGD6uEfx3+jk+
meEjht2Cs8vMYw/7AryodHE87696+inpi8V5Ol6wOi7RdGMDxfz7LaqeQYf/ctiG6OPXGxShzJ2W
dJQcx39zu9Ptc0Em7p7ZKU5baMAa4BjPUoaEEBnAjs1Z43mLUOlvc8+zE6PbXHCV3PopReZI3oS2
O+ntre4t2X5oa4RvxG3kb7JZ57YPaMdtvRPb61vowEmypSP7+Ptsnmaoi8uqtmv5/s8mLJCqrLwt
FmTQRpER6vKf8YnyPCf/lMGWdkGOvS+yf8cAr7PfcJJv2UC97FMFubnp91ope9tdDXE1ZuYHhJy9
CA+6xpUUrcWDD64CVGLR60hjohccQQ7R89CvWdMyAmwrwEsBnsaE/3MOEEZUojD5kuqbo18shTg9
4ziyXDmFit/MZ27XRvZVxTlMpLzZZXkcUsGJBQch6mSE8ZyzNTsbKbVVVMOxa/V1tZrGnH4R1nCj
aqgGx7JcuEHYYyLFNsh8D0sa+KKJ/jZKKBX44uIknSEnIJZRCUhUwgBUxqqBOotcVrWin1pzg2uL
mYEd9ql/A4ta+K86Pp/4a3aNSmlSq/Qrur6vafJgZh0g8xCt/x2KbsuXVfoPIL9FJLQ3Q8YhtypD
KALPFXCa5leAEwfiby2jq2lHTZkBGKHacJ1Nt8RryZWF8wh/qdH8B0c4Fm6VYk5aGPanBoHHqE36
qAL00t3Cll1DkDVy2U6cWKct5lS6xGD7Hv1zS6rrkD8bVuHz0VV+U28EwxJGzGKW1Yg/QvFToxlk
C7hpieBEyH6kLP8sCXv9HojnqgQAd5DaGg8sN+MOE8ywMJtAliSFbflWF17rRv9Mp5H/RTbRkQ/q
+DiI/Sx+DFjQNl+YeJf2NpdRRnV8aRExZsP1oLI681uw+nQb7D1dC9hHfdZI7ksW+ATfhc/QgMu4
i2rjFJ5RDgFYDn8G5w5EfUDTegk+mzLZW2Wilo2WQ+VKeA7jnXPvF3orq6fRQg9Zs7+HAodZ5hkf
UPjZi48t1o/fM71kAPFBYE0V4UfKBseBHiC960gZ/PIQoIA6Ojc3pquSqKyKAAZDKB6pNzLZDaWz
p36xLNya+q9vGy0+lfkJSeZbfw2GypyABjRnJ3KUM8dwq51qEXws2ZXfkxK9A/eEagKeaRIMq/wn
E2CwNYtZoEDgSefi/U5FRmOsvXf6ZjYbcpmHq1S5Y+Z00UHKTAWPMWW/TaPE6EuMyJSyK6D3gnHb
gBn2UADNHQ4hgwIjYNaCZ0aDmQRWMXplSpyhcfwXSiJTAOHa6kutpxloyk7DCptA1LAxPLr5FsTP
DYIXa8iu17bEis5zzTM9PdsOR1l1c43x0SBewWhYZBPLLveEipCMVqDt8uNB3ay+sv2G++rGZTm7
4gDk+HyRchjR3eoYx8Boarh3v1tH6CUPMlElipmndb7UQuDon4H6BWzgsO4yhJCLP2VBrVdsLzv7
BsyfSOA+YT0fjCbndAIOKYOydk4hE0ftbGfh0fn0nX6/iLGZs4lMd/9uIA+3FR5ioDASucOFOQE9
/SYWr/1DE+DVw2coWRp9mCuH4csFH8kIKhL0+4yeKlc8WxxW6u8DrdjBZ8JAazmK6MN9gfsScVCD
wyMCBPEKcQvXato4D4p49wUzbz3fOCvnuIJ/9fScv9QKwQjRT+lLCgV1/7wHEcHQR9W1F/SOhFOl
VWoAILH63CLcleMuvSS90NA3Y5d+eZlQrhI9XU9yjo/slQwJnLvVHTEJ96Y4zjx7LbSDfL6c36xj
tXcBEnTnOafv7jQCWRZE1/xa47xp7/vH4XWKdRx3cqIcrQM+bshwvGpP/IkxHmlJam6V5LbadFNm
dM2yTpJxeb6FbnT+v8zxev4wBJTMRODmpi/8T5rcI9YWWEr5UAL2DUw2DowJ50aTKFW91gBGLhAs
OwndWJiDRJOZ4O8cw3fII3xrC4/w+0MCBonCMMmxcjfYf0oo2gz/5LF3rCd39IiYS0/VLg9ETceT
PrP63ka9aKbYilKbBUth/9USsir2aEdHxvMdo99Q4tKlJoEZ6ZzaIDjwWoVbO/TvS5reG96mpryA
WMQLcdN0mFvVEDqWphjLKOhc8Ste+MReH935crP8SnaW+dAWC16axuoIZ9dbtl3KKo6ap037jhkR
5o52BVubavtZQ0TL6vE1c0gXurXSQlniCGyh9iB9XTWZPp2NU/OJs6QWi1iHjwC791o4JwxykqaF
I8w1JJ0GBJbFKmLFyCMMRvwW6x4Y/IEslddI6oCdlY6brnw8A8R+fvuO37uOqkE/pDCUHD+BDYnq
tMb42N8wa5BHmbzefAc/aRsyttv9vFSN7xs+E/SIYMuJbYOZKxHg3qB01XqkJtdEPfxUAeJz0DQb
vxpwnhperF+Bs0rjYI0rWeVYITbFikdj4eJL9M+eqvTgaf2DJcqFOzJc9PldzgudHc6K39GHpg9Y
fRcTFDG86pJf6BDPI6kkyIqISTRxARIKBFcMloDLZB1qHI3FJ2TXjwK85JByuPCebL66map+I6IS
nxWxSWxJx1X2XxESuvGqZZh/lqLrbW/3LbC6XeFU8RWJNck9r/AePe5yRpGkFQWtF0e7ThcAx8Zh
GyA6Aib+JfOMWkbiiCfUuDneqDBSgbDutGEYsIYCKuwN8Mqec0bzs0Jebbzoi8PcyUWnW8NTG+DE
Uxxbal/yvXp29JNOd5WmLFtnpe86w69tJ4PHzB2NlLyTy5myeqHERPO8Cvag+SDaA5tVQCM4JEfc
UspKfifFMRv8Qy9vgEpeRX4ywdcgtqq9cyMKD/hrT/z2lIXl0EEaz9oXorJjYfiL6AO40sjZkBQy
2DRqL53QZBHs0WEmpPuBiwhdcPzi6i707f9TIeNZ5fPh1SdB6v3cpQ7igtYprY2UcXEXxOf41eYu
O5hw4HBNjdViTkdRYkiBACYT8sI02u61wMl2vUDSgtEwxAmXjXn/XFvFL3RdIwBdQpD8ZK1FS6SS
XAky44zzIrFn2Gbp/CmK9fqO2e+6DYl+urv4e7GQt2PSLXadGkc2Cl6wZ1MjUGTBM8Qrg2qqb4Pd
O5DAfAr5pqZaJVB4qu9sYf5AXzOQQOL7KTbJbBEldQZYdlL72PWApHQiDUthogwe7se+NkGrojgY
bag82iQVPlIojSK3TAQSzkRRbh3yZ8wB3fmXxyYNU9HBjQX01qgbjFTpPEXEYQd+Ye6DM4CpY3IH
Wo7hcSuux+sGR4HJpGjPgDhh3HRf2TXLeB06yAJgh1rL2ueLYX8Ewet3LV+hBXCK948GmOUrKyKM
85sK6ln+3HNLcDoDYUWHNuCUU4j2ZGtZPvzLTz9J6g05q4Mpf+Oe3802x3cMnZx61yGnKqOmddaZ
dAxnZ0xPCJOHpC9REcMewJssMYfMCEJFye2wu4lrcJ7Cq2m76yP/aDnx4g8jUU2AtqLfEgjDdQPF
YGa4m7KRBFO+kMYZeCnK+L61ubBiE+8+NOhdnL5H6YZS145nivzndX5EswRuf4gdRyJnXnXVcYXL
s5mNRSdhOEIG1CeGQTmv/KpFhtgd5/t7Zq+8FeofU5fTYQWTWGF8XGy4F8q4y4m83LAmGAYkhjeV
iDmH2cm34jJ74MC0eOMG08Hmw8q5ZfrRfob+112WA+O267x8I0PJxLNHYQ9+x00JoYyYyKggd3R2
rCQXpetlUFfqD+nhNEemXB1C8eCnsJHNBzy/rsOWpfGIBZqamYAmbBB8RCFw5Wsac5L+VoKsl8LO
DtoaeAu0vxNNLuB1QcArpODTVUUEAZOdrJZ27a+n39DxJoxGC4PygF9BKK0dXkHl7lO7/8SkEFy7
drtG1v6ZbFDZKUT3c50/wmeFaatKLRD5KIPquXeJHWbhNLZGTA6KubwMu+T/yuxpZUf6DuGTT4CL
R9pfbWPdz4HkhwKogBXvBPX0qiLe5IKsibGqnuRAzjtYKS4ahtgR2nejl4c+JGwWdeCGxkBWGGGI
uV9Gyd305dxAVykJ9gbH79rRLyiwHD/ealGmJREArerBeRiWZb57Xu1YPu3+iMXgyuEUVwsXPkk1
tjssyCW6qfypZzErt+mRMbHFcf/PV6IXkfirKQbDuTlquseAql5rDQrliNSLm+ddiI3x86pHL810
z5CINtVGALgV3B+WFC20Z+kkYZqLqIpP8D+k48rmk3qBsuDO0uJuh0q+a+apdfmG+u2zUIPhMODM
9ZZM0z0bNfyaFp4liICnPbIiXe2EMPBFuyzVIC4Mm7HCY+VCWFXqri69zMG71zqODdyrWUmqPXQJ
rqSdFmsr50uDSVZlylxoqQm+m00/qJGfAEjLhopw0SMW2MdQLjGgZx1m29yOKmCORD1cBOYe+eaU
46EiT0naQxKJXA84PCkm+D1mnpRsuPLevmTZQYGtPkt7JRdUwLWXJWww0ioU9g4bRriRISkix9ZJ
WjpKjrfaD6LGg70uoisigHtKGTmL2q+2eKPW0E4kHgg7q5IPOlFsCOi+IQLHlsyDGoUVP2iho8/p
1tP6hgFouoV+DQ6xZ3urjcBp9IfklZ2okMRV6smaIg7k7QZPTaE5rrRQyQNj54BCy2i6ioRk1zMn
/GrfM+3ZsFFtRrTMyLVtFS1CWDi13gHHTsk+pQaASpsJZnojvuJ+Facxq1Qx4E1haDtnEoY3e1sy
95Q5rN5WBS2l7C5MClEmWlAoNngwG9QEg4UDkYFb8lomAiU1HDZFg8J/5HaswrZyUsrMshAJ8IJR
wy56TsiuWuJtSaONz041uhJfsKWcYskEwsbb8QgzB1UEqKwmlQkTwzVxzIsM4VX9KxjEvAk2UFkP
gv8UD5YmXuFA4SHRJX4WNvXcqI1h/jfhjnEP5Anqb/Gl/O95RZRHmTHbTJhE9l3yIw968QQiYorn
Tp6eptcMSaihIYF8XJDUBZgUY+wk/F8vKTMr7R1avEgZM0avU4qn2S1R7f3ubs1EzzQw4gOhldWX
jtHvEOvGEDX1maw6Wh81wmTyr96Ic55bmPivzSQD+IjcyQ0bzuqEJtcQlaUvZM5k3QZuZEoMDFEs
x1IJCYEynaUgNcbhHBJNoSmodblOHIVHHvd1Hn+3A8YbZEf+SudOdUmDU328+BlOlz0nZmMyssp9
IRBfJv9IhOL4YcA5VxHHgu5Mc0ja9dQK0EbFQz+zM9fII32mFfF+V7Q/A3RX/elMrbCV01zfnYbv
OQw17K79KaPx+MEPiJqGsWZMR9alpZ+U2bEnimOHpV2gZwqrJWyNMXPWIEfX/iRknM+F31Vc44Bw
ZP83WPwGRorRfLdWjHS8l+ostomexunAd8aDuRVEa/lyVjoUqNZACi3icsb2tBclV4ZP5GQ2n0wk
PUO4hi0tcPrq/0AKnOcBd5037o3ryxUAOZ7WZur3RjBYPaIZ7QN4cu2Auvk0+IQZQhSgfldtztkR
3PhvWFHA9AXURYGhkit1SSkl9YWGVbrCVMSHvcBDel36RoaqzNF0FrQ38/jYhuYfemz9SpIe0pAJ
UWEMMLTc2pYMxkGB+ylfQaHBuXgERE+kAlP25XqQwuiMz5cheOxZ5TPHcF9uzq75e1uVpr4VpGJe
T0YFUsHn+kubA9ilQTHXfnhybqTYiRDofog2lLWjO9wkiab3RTSdsduZhnshv99/JrE9OtTNMdPi
FftaINIakHP2n9A6OjW+kQafr0YCy3cN3QJWS+lIgIgeKYxiLjrSctHQeAB2TPZFeRq9LZmy7vdb
q4nYBIoPYC5n4xMQcn1hRXZBMScUPViouWoaO+I7E98HO2/P9SO01+uXHFhRAntkdykQ34p6qv2D
nWxiCJ6HltsbfJyUkVdqMfr1rl7gMOvU3Htdv19wtXeTg+uNoIiwJwi6E5sSj1C3W6vSivFSMZrX
t3jStFIcL3SbLXzmAJtwBKd9BVmpIZ0JHWceUY+6yJ+mMluS8YG81EHFQp0Vo/JCf8egEMhZ9KG8
jaOlTiQ8g/U6v6y6Lj1TcHbx2814uS1mI2szJc2Q9Lp5r2adiJ78FiZXMui2rCIY8U5xrbqG30WT
cT2hjYKOOrybukzKAFW2n3R93oeRrwyKVT3WqMeMP/QTFKKaK7w2cVlZ84Ck+B3RQdei3vnl9wVy
bfZNM7H8cMxZFngmRhK34JBXGmyYY0k/AMsh7hE15O+Ag2553szgRQdfJo5yN04lwIjZwIuJCF16
RDhkXyeJ5TObdNahkwyZDE8GVdi8aef1U0C/xnSGKkgW79615RGIQuROTJYiocvz3PcBpyuedb2Q
CCRdCiY6mNYDsYYt6ucJ3PDS0likOWrx9UFMCHHU2l3Rq8BTokdnK9e6CtKdv2ixIvAYd0nmhC02
c26Siu9z3jX+C0l4TdrDxv/YnR3YQOj69+vhNsDER6EbOAuvpe6TOd0VGaDjX3LKvAzWYjCqEDer
FCjz+Dkuru5BFNM4dYii3aChieCo39nSDwsNoGbRopGiiTZy+MM5viZafpOw69wyOBrD+oHq4Zvp
NUoHqpgD/mDmRPlptnurKxhbagLC5Fnchg6UGqw69Uq637LG9IefzBVFB9K/kZFGDxGQfWRx0yPb
54rqCxGerOuFD9P/Lk32m+ac8LxDL1fvAyBGKp80RhZfzL/hA3C6pqc6LP86KlwLX82Od71mT9cf
SN8bKNC+zndlrOGr4Ittkd8pjHWGCkXKRaCyA2XE2YK2o8aPQ2uHRYmS85KFYtxAuMmMrtAYA+XF
sPKWcIe+n7RHO1anwWTJByA5r0WO0QRisrI1ZRLs2vJO2cS9rdcbnsxC3FLdbBjYbuPEgqRh+k+U
tAVFyiFktn+Fw+n7X5KX8tawoqe8QRJsA6MheQEwbC61+UnqjWCnzFwNioxrZemH+1JT1YOUsqb+
8zBR3iMkrtvgcKxQoJ2pCGEgym4a9eYLbsqsphk+WdkZmBRtPzEtSgVZ/fu3zjanLAWbNBwM/amU
ojt86Aocs09fdff1v8Bi3txgTS3cA/nNJ9yelIJ66B31kT4RilVBjnHDUYdNkpzrcyippIyXnezo
Z6z28JNfDVv6PAewLzz7U80T8+VAcEf7xJB+svYts7IqZnIz5bw7bWTOOG0S4UyrnVK8IIYB2/tB
iuQDWuEnYpa6H7UszeFWtb5gVK+u66BS9TBr4FKDotLqO8CJVnoX4DPeLUn3K4T3t3HRuXvzi6PS
OtJcgA/bLPAjoriIrVcmswJjGhSMn9rwY5z6kot32iQEYxb02nPiS6b+x2FFxPeVS2WmKsv4sFxs
+PF/9nSe1xipW64aQ++U2/wGU7pa54dQ67dgYSexmUIhtnpp4FOIzGgLwOUvUfmr5Y+a0palfLXT
a10pWSLrnsyfLRKT+8GE4FcAZ/5UcFKxaqc8W7wiwUrdyK3vaxtB3HLZr2+3i6aZLTJ6qJCp8YTz
MdrkoeFgZShaVxYHDjj2pxkykS04zvqjsNmpR+Q6ya1JoziRc8zr7U3Z08oOxUXRuNO1s6aF/t/q
E5gT7EOMnR/NioJxEwvJPznTrTnrt/VXCErbvn6KaVeYvQg5iJ8ihr4SBD4KzfBQNLzmUf7/BiX7
LAAXSdcnyq7GDhLmuxypPFv3SoeCJXqvqogwd208+HVXQgbCh7tTSg2NAqe8P5egxPm6eqBGrnKG
dOCZcwm1EAJNv+xzUr0NsaQj4hJnqOYjOfW0P88KDUK2eYyzHgV2HGjk0yq7H8UeJvyPsiVr2EF8
afDnk9DYdMy7r9f6pJzLBsLvtmitbAWxIXec5zGdsdiPoOvS3PJvSIR1ziOpt90z2ctRYmqIeqAY
kT6nLTUg+eyO57EyccI1nSjoAyVLXx0PohoM54XVAL43MC5xeWxJpJqICSOa545Uq6F5CsteTEeS
/oTNxz8oK0cKLQig/JF4aWaMsKhzlIDS0NALIiLVlmuOiJaIqF1vV7waf0/dtgX1Y9XuMlPqQCig
WHZY1z9S4iF9RMspc0i7gxaBQVHkQNhFdaMVwIdlXFO97Mior1K9FjCPfWNS4tafWHIzm5tUXXfo
DfhErqz1jA7oY9rmr9d3SDT7Z5BZnwoLhDPaTf0y2zwVN1NJNtr/nIVnaGdzUvOhc6+DzDJgmSXz
gMH94HqhN3FGOVXFEM5zBPeOn8xPqm93uSLnVZRQ08yi/tVHzeo0miAKx90t+7ZUxW3ZhzwjFWcl
0EdY91ekB+1IK1eRhU9NXI79DzTiPhuGbTrIB31Ky4gmq8jdLFuJbsB7d1Q+7eLvx3qw+7xbQRTd
eztKnp9JsBb6/1Hc0aim7VOXRt/pBKG/BHKtyJoKbZA2sPvh6Z9pow7FF2qWcZUiUeVa151IT1An
/4m2qbLtTRHhe0MMSDxKPZmrsnd3zO0AOm8vcnYI9BngdP5d4dwiRUWW6ayDMZorGxxHYx1S7Px9
5HwIxNRai8EZPnI4wCudtCOmEN6xTgkMOVt68BoNkyjUc6vCACXjn4QvvFvUQVtxkOXs+hXsN6QP
hId/8s8XzNHMp853mdMprzderx5bCzlOTofUeCQiKiiz4xKN0dRyV3PSN+uWiX6YGu3PGNQpu0IS
Zghek8wZwCG27SOX9ArfRINr6Ur4p/2mQyosstfB/Sr4a5P5/YcP/viWcVLn0EAmy3dT8kx02l61
NlBBdrtVogzr4bzqEmTOWI4lgfdnqzmcTahxtBI6b7OB8C8bJ+R4eUteA1c9ZHsNPFwbNojfsJo6
8JUc7pQRxULA3o1SlpaAAHO77pAZxTy4ydoudATBJYoyNNOZ4uJjB7xvWCBrxdjSRPWcbCexIYA3
KweTKlFh1ROrP2eq2FtUokTANaSmhY5VJgTmXmJTMs7C7cJFyzNUf0k93VsNTlJVhAbfP7zhzZil
QZqF6QMECMoylDpjothl6TAPYx44ASNY4/lupXXpU7hqwDlCT8l7Ed/EpvxGY4b6qtM1Vcig40yf
VXx8Jd48LkDzQ3iRbAtM4thFmTm9Ov5yhcBTNaub7UyaseDaOHFuKaXhWxbSFDMC4gp0/UvvJCiP
ysBEkkmji+q3KG8PIn7cDTA2U4Z4TNc5/rmWPKSy3My4nICSugea9rABrIB+DAtWKflIXLia8Ikd
J/CeHKZ3X6eyCqO1225im4dDt/UQvPf5dqoZUAEC35in5T4yNK9rBMpWPWUXd4WZxDCzaguzt+t/
pk/dKlLKYzXcXe0PwzwQJwB6/7qRWmnHylB32rKY9CxXZXQqzKEwVafbdNlfbGf2sxw+MZ0GWXiy
RfVfweRNtmlbM4WhQuyFKx1rrn9KiTGFSNZHemAuCTYAKAQz2824Sm3JjVa0uaB+rSbBRv4fDnJX
UHgmErpG1k0neHl7YEOtKxfRud5TBuGi/Ldxa+v9SV8tAX3O0whisXanZkdpgCXoXqYIauJZS+xM
OEYEikccDJgUlHWTcVNtnv4wdXi0ph7hirsf70m6bE+HnXQTIa+bNAeGsMzqKQWR74o3a6Ql8MbR
w82NLg6jNC6if0IAuCd29XR4wWzldZRh49A5md3/Rda38ViBrqIt1ZFY0v4y2zkEC4+pafQpjJCA
f9huGco/1WCjmPZJDvsfMaS4P4tI2fp2dEW3qvgcyU4gfn+Kdv+/L6nqI5fQaY7VSenOHiID0t4q
Daeur+gC9Yi2CH2JBwQDj0slWJtK51oOiRvVXYcMxSpUpwJztMzYLKjtlaj8qS4EB4jk0m0p1Gp9
WATO2BNo8QfDdSKYMWj6UrFKt2irVD0SEfgpQAA4tleUpWLfL8VHeLxSKbtJ8XjxvA2Zuk3T+toY
XMCUHTa4+SUeK1pSOH0Omji4cyZyh5m/DS3BjVRo+rfnnPAzslnT/tes73kVfY14u9iAVYnJwsoB
CKdBLyIKe51UdvjWhezn6/UidIHv7wsJH0HoBNshp6iJx4Qdb4ZYERTi+n+eV7JbbRXYUSVsO0d1
YSQWmrMkM8ye4Snp9giCf6GDDBNSmuW2/NrZtfi5/HW+xtnWWXgm3hEX72vxgVgkpCG7Yd3m3Pbe
4rompkmNuqXiy+wJjz/OZ9VhaeQRuSe0mqY45v3TW8D3CxFz6ExSYJ2iDHxok66SaKK/KhKhM0Tf
fVjkvt9nsU6SLtmDWCF0tQCubDJPMfKiH2sXgvJufT2LADdDSkhdp46885HUZAzVFL/DitEHGdaW
LUdl0MHfI5idvnqofqetnuwRGyoiirzlSt09dZizS16Bzgm5K1wKjZ5/TTZZUd+2A+DQz9KiimmS
K+ykCj5DlqKWL4W2O3+0sLlNUeyfdJv0/ws3AHpHPtokP/H8Exr3TfojF+5yPDlVWNuEWrOQxkXD
sDeWqrOw0o0Ckdcy9BjDNzycbxQM5hfHZYpaABFEdtXgihmMFL/UBanONCEubA4oLVqBhL1J7gW7
1puuTptW3Ad8uFnKdVdRbEln2j6i4VHchfO2GwTl34/nDgF2eaVVrjP5e8q8A1ee1++gUyP050Is
ZD/p02lHnBh79PlH4YmzbGO4Wvqs53YqevykF4/kCzG/xsnBPBPuFatG1848FCQVO2ya15b05eLT
m+9baSIqsfV47T3IVsJ97UYfyAinWnssef9O74xbDkGsQ0N1r8yrUYpl70uQyqrgFo6/ZmNLZQvM
OsOCEsHhQu/UYYX6IIbc6DG75ZmAAoPY96lqpSPTI1n/bd93qWbw29OT3iXFWPeU1IDtoLcS1v0P
eMlT+3FRSQQE87YMdXKsioY8l4pPnL4COnLTNaIyLgMglfSu/zesDDdo0C69iClQ/v0KCeU6i79T
0LZnswLcoWIpilBlGlCpg/qg3ZXQtdMTkC+cwFhUaV4VOIdQ0On4JzfQdCr91qTdajtCb2Cp4NxQ
8EFcnss/D9v3h6d2fdoz/sENCg4LfgYF+Sfo6VcsgeZI/CaOgr4AaETWrpF/rL648NNO93kSju2j
wh5blHVGE7q0nbNjo91jtcMZ6Li8WNQWrx+L8+cUpZfVwo4VaERKxDtNi9CZcUBFql2DnSCTHswQ
bBcBwTxQ5ghZob9OwKrMLF0dG/dys4T+l1bKFXpbtX7aJpHsgX0gZSfiSqou7p1Oxc+lP6UEQVyj
SDe9ppAKllu8eJmS5ERW1z5AXwmtIeYVvee97t2EYCu1ZAoQBLidseUPcKG6NTbFf12Y+7vmHt2h
3ECpiEADnGv0J+yXw47O57ghd1xs8qTS3p9LGU/l49ov9T01mllI6lZbG3OJDkd355FtMGIurS6d
LFFYPcU1I4sJ8LkvD4oc0QekONTIxEW5n6SClkfHAbMqBs7r4wAvuvbeC8ykgL8o8u6eSrJJwary
3U/j+baylZ5Kzr7C/WrgTlFJaKm7p7CEOMqYrlGCZYnCr0dhgbPZ2CN6vYfdeihj+CeVKGCdE9Y6
3LR0Zu0CJSCM5WheoNXrIUBetQ0C2F2nLNxUKQHhO2by0voQN6ihasPR6Kwx4ZtCmj7gT+PyHT6O
h+6jYiKUamISg45cTHocZ1rGA4/jJjcint+93bTMX/YN7WGXkrvd7VvHNYwCe2G3zhXt8mKan5O6
6Rl7O8YyDvzGZycLqaNnI4e21FVgI/UwM6ERmiTRvPwf3ghSgruTSY+SNE681AJXoKKjUwiZhqkb
QCsqblukhvZBScaOfBscC4w7bjmGDi06jGswUN9kWYzGJeo/LF2dVQM+xdGoeQq3ZX4pCh2NWvoX
0rpNlFA7p9KLylXB9T1DMze/jtbmpZat+XZI7LGGbInAMZ9lczapqPqE7WwLr5eHejfaiYdmlyD8
zBtc1EvJBF3PADnLH4DSoLO1rSuLRNxlQ4ZRaQSgd/7eiXe4ijLQDv8+aZZwnwdKsNUKUPvnvQIh
wuTrpCsTSAka0nOWRypWp/JyluR686VblTDgOHAkPwvcybKbDXIU4zf2TTU463nrDUqwu5tHSlqI
pyfjnbb/1lpbRTE9QHbCqmuxaV1WAMnmMJtXWTYsPgK+ZjoU/X7L2h9Yq/pfNNOaxtSxP0Y4LqfY
KOhyFV3+jw1eCUOS4w8aUxXe+AFXpwgBR4+Ws/dlHcYgnsCrjIO1+nGx/p15MFGcDHcoaiZeMzpr
fkpwWs6U81+Ivan5ELbv4RkKX85FFzoXUjKSuseiHuyhos5CxHdtF5KDrmsQySQz3/dZ+9qssdZu
ZD1isy+s/5Cl0BPZjKxf8TlKM4Hm6YRUptEcd7wOGVSWRD/pk8dmwD7P6w2fcMtBdVkyJk1qZuyR
wiV+KXHWIKcjcrrQGLibZyKIXyy3399C2ZGFNjbAvyL9nCkSIMK3sxlIJhPvZbnvRd/WaIVoMAaj
f9lW9bmQczSM9ojuxWbMTeYyl0pjz09CSRDNyagEy40Zvpkl5GEeHgLi6mgf4DIMSzyNBqbopw7G
vKQvGdFK9wFA+n2ES6/WFCmuCNZa5gSnh8HqtLbx+pV7vA4nSTh/XDj96BiVDfB3Zf4DP8023qf4
Jn69cceOgXZPkJ9qrvNzxDiKIpLD8eASGmcftY/sMHdsEOtPY5z+sOKGNyBP6rL3xUKjljs0XkHD
IaRgE0mLsH/cEJjr6FUQk4guFA5Va1doWL1kOOPQuGfFRZPwdYgp4z3hcaf7NK1ALwxejlzSwdg0
NGDD2fTT5muQw+DJ+1AQTzoSOoIDojb9skh39eEFfVvKRDfkXtIBFlOfMRtkMuonCIHzgrcw1QIZ
dQ8oYLYOR4IcR88oNbp6t/ZBwySCWqBd5YGlylCzC+TA3TH4+CW3UaLuz0MJmCIYPsWjngafuIIP
x4zRSOTEKmfkkl5ZvmvhyFaVpr0Ay04+iSBrkQ+BsYyEAtpfnqZPybA2onHyOZwv2+4wiFgV92hX
EMIUnfM7Y8r+o4RSxU/5gVD/9idTPFApqwIPhF1hx11JeXnizj+9qWOOJofrYxBLScIInlZy2EdU
4/Y5e89oMk1Z30Dp1/FLpfIDSxMdRoQ3wGyu+aqFT6ZzfGqFtddAxOdS7OPzUaXXjmwk5hesgZkj
pdz3v51Wd01bWnlKKqQeS5z8GfpV5Ag6I3NvqH3+ujs1sERYOkKJYuAt0MwpIn0JEaSssJqlvDwL
aAiK0M8lKG0FB0ZxRbxI+eIjhIDtDeeMjyUg5Huei3bi9k5fRsR2G8PT4nvxZoiWoOnq0e8/CfCc
uH8EGsiCEBhkr5dbMp8HPz5Tidm76DElrrDrAArTZBK8ggkYAebSdvLQ6dVpyjbEooH6Xgv/9rmu
zvs9QN33upJpIzeBypteciXLaYKaMofAXLskNPH3tpK8d2xQpp5A0ArkkV/O8CxXsGJOKswOLJwS
aHKho33WIZKje48m35Rj/JrXTiv/QAJEIkRX7rAZofHuVCconFngyyZdZZfBqidLMjraTWIwkvb1
Y5J4SZeKiPZFjeRonVyDFLpAuN/7bcvXK013LoORopoXttgxeXhEjeJB3+uny8Sl49YWk/BU6K2A
xFkenjWZB4/zl2o9R6Wmv6359/HJSNZx+IEQMbloyhCUxJEIYaBbUUAlu+fYHz7EmL5BGYXGxr/+
+31LCzb+HT3AyQOJ1RFO+jEp9U+sTcRdtmBJXe4MS9YPEM6kYEDk8dPU/2Rfvkm6qpsuODnWVqFJ
3djXlewhVrcDk75PBdjbmiWyy2TMisjo8c9LFJP9gJsz/D6hThBvugc22+3jSHd4TnCA0RLJU4di
C5BjlmE5fbUBrqFBvrjv0FqBvF3+xNACRYcGsCJ9MNHaBBpZ27xOC2dRsGjYc98YZjocK3Kw7u91
jgx4fcwgBxpWAXGmtbNx3lH2aR1pdyP+etU3hFg9hQ0MPM3C9GXMkHGhwC7WTd++npRMHW29Hj1r
o7B+QGEJmulKLA8ed/FmYuggN1svFHZNdv3d3KcS4K0t9KkXqqs7Fimi2qrXXukT7bLCQihne4ye
GHAZapVZZcv/JHwzRXyo+FnPzS+jEQcLD9XOjBxMjtL4vMllL92XMhMR+ZB+y7Au6a7WiFTHY5ya
KS6CoUbQEBUYg39T/1SDithEDGnRamCfim3nokPrqaHE6s5gprH/h9uPEdSZdQTTyvIVg3WYwnRs
m3gwfYbvhQh1Cqmc911gefUKtnlBOQBzmbF4Gs+hZTGM1BLZTX/ldLPvkBz3g8yW25Z3uZONGOh5
6ljSA5X5LN8GSEkvDzQuWwMjTGjfbdyL/q87sE+ejrzoFDu/DVyyHodcNY7jf2duKW8QkiYBlJfM
ckPYvcH6EvSMGWHwXON3icVKX3+j4Fc6NxSCMsAyjuWx3fhzeVWP7CHOMjmFtyXPjhlDUivvFN8p
zJ+mbp8VAg4GLZ4VW8y2T4uxUENkkyz20WDwKothKBKfT/hfnscpAa/CubpCZgjdEKn3OuBJzVQQ
5Zs+ADS4UUm4hv6NImwuod79O/DWpgq6Rzy6Fzq8yduIqvvsW/6TWEse9SXXcjbYneXknYaAcXS0
HpiSLuG4zz9RinAZT4ZCUR2YPfQa24TYxrcEupTT1jaRBe0bDvi56gTENH/x7iFR6ptuJy6mp6kf
Ue2hDBn28jI/mrurLTdfber6zql8s4XPt8RrqH2Eo8I5fmH2I0pzd40C7QOCeCy2VLkcF7/mprPk
3VSh34OO7sw9HnyWJENLzeqOG2PwB8gJdZVWhS9X25bL0UVm/wGqQAaRKYK2ULDj6ImRlMq0V3mj
rIGICyCAFJZF/K6zvqZvH+Xm676+IrUfnUrVY/F6TlRXTLbDIOsCxZA2IagvKtJHNi/+mO8pR8A5
4ig/lMbPBL36J3V9W0CDLaxPfJavnKq/0/7c8AmJIqVcjT5BT+aIeFxTktseuO0l/5rfpwu1uoFA
ISE63Lg+VJMnYxqBdtGjdRom+2+kk9dlV13RTdDyUWwjIgAjW6smeFKE6vEBjSjAn+Z24wKfvZiE
ax9YUGw0KSYMgi7usaOD0EejtcQPtIFzTv1GF+coXpx9BY/Q1sx2y/etooiMmT8tBCAfGSaw4zF+
+5lzLuI9XbyUZ0X3arAKBKN0z6Nj5XhZJMSdSuiu7i1JojuTNPHHD9PCHHUhYXZJhChYeJ0vSuQF
s0m0j4L6exYLaX49S4umUnk1q/l0Xvvg7kCds6uX4EtwxFBqrasIfX+aKzrb2VfdCZeXnkLfKDlJ
1YqqsFhcBmUjSg7v0UxvNiBoZn7plguSuWAn89mYLCBPrTsd6Z+QLIEPVzfTE8Pg5dz6Rrdvi/mf
rqthD4btaEOH+x8s2+GJbCgunwsBKseu0rJwSOg4lwI92UUuo7ISjW5gW0+Ud3SsFKf/lI6tKZpf
9iNca5nBfqnLQ2Gdk3TpVcRDGp212IPWvqxGL740g8NAEYez85q8bDF2Y4hrVIs8bcoAj/RMy/zu
V3stkn1kPy8NN/Jy8j2LK8YEVVvUgV7MItpc0aKf4AoONSsSp7rqHAh/y+C2iTp0+P0GJpktqPi5
BvZ51g4WN8uOGJM1NfciS/n1hnQfkrRbvilfO78Z5atmwy1Rcd0CWCbWQQbIm29ESkDKdLlHKjGH
d3pJ1f6wz3vajRvADC7cbSeXo4A4UporAgLpqYvqGKBXXXvG5kivkZD1aqb+/fjWRyJYMiWueV1A
vyHCA6cLnZ+R2vozHLvLQrYNsIlzfmALbkDCBKjGmuuhlbA6nCTkaO25f5r48KZWt8E7FZLtB+cC
NGw6p018XiZnUV4EwhIKxvJQ448wSGf66Eu/rTY5WFXVEVu7PNEuAg7hNmCUlJDYgCzjjclptBQk
mfVLA4mGxQ/8joWtYyKTWMZIx2mDAXEJvbM6QdhIhq197Omc/hUeJPeorAa/ZKHg7oQ/0RyBPYea
VwO2VMbKja1XyQ0qDyWWTjD8Qz5/WZJqb11Nu9hVd4CLLkGjUnkHaCg2mGLL9B9BraXW2j5fzSmC
Em2qw1pw9WS7YErF5IKG0dWhZBwwRxS57jUDLRzksQqeioD8hWJGgYtWnnKFh55NMxUIgm2fqHXA
GVEJ8I6w6A1KvzUQ6Tq/puAMEldWb/rM8c1vBfgtf0N2MNAjRlj8UJ7TpfydVV1uTbrBJArqIQEp
R6XEbE5I4dyJn8k21MeBro1+8U3cLaux9aQYSGZcI484EI3uS4rWuozafxF/15ki1yaAVhw1j/YU
QjDAGu+11OcpkSQ6e3EMRG3VDi199jzknAPSJoZuB5Tme+vt/oKJDXDf0F3brEHd/O485m6fux8r
83XXgQ9sTj9eKsSLHmJerzJR0VJBBUCYUNV5uVg+drWIiyURzDbgq3hmQVRa6xhYCoU2dgBNYdHZ
vcJAbwtYLTxL78UuXjZdgwut3VszXrnJMbpXvAteqJoGCjy1EbqtaLP5qtrgN88sW3ak5b5P9Mdz
Pe0+3GaI10FXpc1+QUdWIQ0PMKH1FU9KWnobcBhWx0EZpeJJ4Y38P0T+GMX8iIT7vkxKOnEqKrkA
0TUeaLVzksiebQwlz2+kjK/K/XkttnOyFk11m9NVkN2cXEm4ylczi+ZEb9qB7eplUC0Xndet0NIG
JMlHP2wUgRFg/wDAJOTbV76oadj/VL5srWCw2RrbjjuV+1VvN5LBJAHY+BWglew9vaEF4QRiayYZ
CFCYHiM4dOKil0HpI4gZRZCupoVu4MFW0GtFhdK+KZThpQ7Y5v4dMIFieDFjy4q9aVExxUUPttB9
rvlwhhgUesIqpnTSgS6TcCm2VxiwDI/ipikhL5GReFfBZcMMeofBbsZVNJBice4qS+4U6BuduLdM
lhE8cgjP2M7H8X3M7LPpQSM07JsYqIkjTR0UAS0pkGggUzcrwQR0o6YhuQAg9TmDJWr+k4nhEwCp
ueB6n8wNwCWGb7oYAigvTwt2EEX7aay5H1Hxfn8GFYzYmYdgEInOnv4ickrh8SgDOcBI9gW7ztDm
IuinPQrFAoJ+wC119WxS5PGvXj54zixO3sE/g4NV4tXhQwvG492opfAiMlF7btMOO0exOQKDuhTN
TjJUkm+IQrgSG7krmskhc0Ou0LaNQoJ+5/bzxnccS2ryQZciySbxSfqW81FQ7Qyye55g7W9O8cKH
7tMuMEyE3TXF8gNhceheDXHXs15bRO49QgLNeNmRHAfG0HQ2g1LfNt54Dx4qJ9jVwLxtGDl0Rkyp
zh6zwfsVNO70K9L5OU+LwakA9ai+fP6FVzLs3eSo4/PEFf/3yDhhu6EQmaQSZ28aLoOoHD86LYUJ
9zrHg6f3osk12yRYyYwDNibeYxhU2djrjA1wwjYvqgqyLNS3ebUJrjpZOdfBmaUvFrXY44wsk4jw
1DN0MieE6gSxCJ3C/A382coje2fiRjh5v2yw/HJcG9Azjl5iokXEebIRap7WAMt7aCwlGVf8crwi
gvIb7gWZoWM4LDaQIclnGypiTn60YUqmVCIl4SCM2PitlWJjPK5Qzm63opzZ9hf10aN4imKkVkGx
ef+8445ionCTmvyHHT0JhgiDbtANithQsZfhZsv8JCJ7R3EIZNxnKf04FGbLkOtY2BdkPtp8TS47
6He3+IsVEX/bBgbCJB1tUWOTpZBavyJVGVJS9Iez/Kds2g62JVlGomILfx6coLACI+0632I8jmUf
IJ0pPNy6tNi879YrLTPSKCLAYziFj423jsT9mmQKUKSnt9hG723nRigW+wGlMHEJTmblk3Dobjio
BsdtXjWlPEq1uxi0P22X/DVEqgnv8zsoF4efqUl3kxfkO1TWIO9kRBB3da10oe/C6Oq0a87iAHpt
KCatoVQmSU7Sz8K+phwmK7ftK1WYX58LdVnzuap3KnguafUtSYVpYIBMWPSmUII3UA6GcGKzIRAH
XX6lrcT5yMBtSiTguiAs/S3wUBi4tVdqcZAzp+ZtxPlfWV6dS3nz/LsDk4GleokTTCPEq11ZpO6l
z33FzCMyeMXpLJv1u70Fcf9noUIogWmw7K1+fe1mlwNuKP1G+Cct7tIUyg/CFu2erZ6Euj1kN6/y
oMf1zrTNROlGXNvskOM62Lb9SOWkx3zMs17wPlw7oV+ZNCicYJQDDrYcRgl2AqMjl9TvWKD/Efnk
vbLA9x4PEsn9GXdGd6bNlLs41/TsdU/ThjiuoKuPYhAL/eTWaeada7+xDwjAu5FQe+zDgxaPURa/
1QaD6cciuyWCuhR4dRxfDdAdElQpe6Fr3urezUbMDk61iK35hEMo8T2881+Oiez9OVeySZKkJ3N2
49DaMyg9rt0q0/I0OnYuujtLUFQgTkMDpmvveqxfraLEfBHgUy+PV0mAyJzZkEH+it/0qWXHFHG1
qB8KWdBp49eZlLiGxSE4f1fcmrRygifN+Pxz9rEVTHWhBvkngBCrOM1vM8E4BfVXghVv8STGcPQ7
lgzziVA5or3OKE+VTEEvaXIUHySQ2x+6+vLMTk6eDo4qcDi3Ui0V/nWsjjdZ2TF/foELA6hePaCg
94OiWjBEVShNih0mpr+XcbLyrBT8bPvw/lh+6oaovIDM5lPYZ4IjfdePdRz9//g1QBb7Hu3zfC0j
M0bt1CObz12p4uFd37ioQ5UH0CvVseu1JPsOUCA4SCB2bTS3dfSIyrHNnDRI8U4tPYdZ5a89hfdj
7+OGuccLkU74L2TgETEzCgs8z+4qrcE3p6InQqZtMCohYqCxu4y0SEo2l4z1iASkISopsh0gw/qd
NKpPyYyfxzpXj8lvJun1Uc0M8FiPNYJv6yI2gZejGFcswjqQZ9qGle6a/VGjV86bJx1rXFqGpmyF
4cCKi4gazjiL7eVfSktfdOXnClLbqJ55tY8d52wKEn2IrP6ZUHPqPaIwfGBx6fI8qDUHTGtHYw/9
RHlH12O2oaR1OSFlYtwZ8V60lEO2HB0t1mF1JgDsgdXSTrhVYPsRKiqVMlyNLDgnHyTSzrctXXYr
IPRlZ+aZS0ce5qQsfIvbnvQ5z8sIEf0u3u4coYPsAOs8SJPLzU/a5+4v3kUwPR98ggmAj8bPx9vs
4QCTqsanMiFOqtao0bmDej7ueU/iQh9CZTu8ESBQ2+QJBdz4GsylFGPCdOcbgYcMA4cQn9XvSUFi
29SBav1E5YGeQDCcwzkK3RaHXnh/FtlHn2oDcP8MiK/l0bPA0hvz8DbvknSlo3febBqSdkQ9EzUr
BL8CRyW7StuygYg1n55+dFHVykKmIT83TCQEht2pc50ZCmqi3NdmwzENoZUWxs50PLGmoNVnPrYp
UlqGZzREOdgiAyUPNAm5gowc12H8obmixny0ekVkZNFe07Z4zthmsPAQGrG5roI/vJ3oMtn2LW1u
0j+QShpoJs45F5+924mLQQYXTimIl3Zvbr1Mc1TE0aUKgVC9AMSvZpgcTfP9Aue+XgJD9aTNXsDc
N1h3j5LfxW2hQZo6LWp74XLEJjgiNPnblp6EeAO5kIjfs1EWqyeXK9XaBal8yUU4Vv/W5n7PhOzU
G9Ez639iD3/bNhWY34KEig0A6937xiB8E44sVlv65HnDMoAcjmSRXMhyiiaxUCl6crZ2hSSgwuXe
qi5hmXDKhbDv5tjQS9PErsl6llECL6ppXvB/inanVA4TtHeuc7eRaSPFCOYGRTeLSQeDbkCqlVcy
Rj+QaIL9PDCR6q7cdi84z9XQwmU/7dTmEF7THQDKmAhtdARIoTxLIT1d2gYoXAf+t2kzhqJFMMb0
G55a44bKrPTqW/OA4AhUOK9KLOMVZi8qK9yc1C4F/nRYaZGc+8J0MNQTcPCOUxn+rUWSe+o1zB+n
udSchlijHqohPNw4sojXHc/nRPC+s7iIxaZXlYVB2gjgd7/UiyQXQFz8tllVyS+Qlw+H0yiX5ocq
Azhx8kjp7kkgBSzkOllxwbyUCjuo85Pi7YdXQjyFK3+eJheJstm1HWZjcpoc1ak0xmc3D6CyokFa
2g1SIdo2omia/ifmeqDuXOsNIj9qmleBvwfs5Ajr0Vwao/dXL/hO2WD+ESGCfP5HTo1k4XzyyuxO
HWmR6V7pcdJeuFOmZrhl9cxtKPm5eH+AUl1P60eayFT4g6fim7ZV9w3ODhUJ1loPrBmKxFg3xO/1
rQKcmanzvmOSDKnud4YdNC2AZ4pRDqcwm+aeTJpXxAcJhdYbcgIpDJaBevX5Ub2QHohgRVhRt4Ec
yxQBs+n8nVEaOLQPBTiQekkm7FkdCJcf8/jiY17hrXOSPhRavN784YMJ4u5OSNFClseLLXSxj7Ab
nadcQpuVpYJ8StGpIOcEp3X7KS0twJb8FVO/raDnfBgTJZB5qaLmYnb59vNoUOBhNuXkg8LPz0QV
hCj+isPxhXeVmhf0RQsWbe+o+n9sh4QJBY0XT2zoFlHXuazHob3xdYSxOPSHfaLpQydgHwFAbvPp
5LFUhEC5JicTnTA6awBEI30utmWcbBOcB+3v6styw7HoIXSxPO60Z4a2H71/17hZeqqSZZGFy6Pu
CfyMoNKqTjq/w6p3ColprTOcFHOzyaO10KF+XfWP3UScztAxsC9zX1S17WHaHNLMKhqqJCULfGkC
V6+/MaeD97AYDnBbqw6A6TzY8yLsmnYpEbM2/wV0peFA6yves3if1lFDpbDGPeYl2B7p8e+xaZ40
vCXUTxwrnEmv0TK5ZT4jvNYVwMUQtvvUN5VodcwWJnr306fsw5uBkH+K/pQjFl9t/syt+ek/6rFW
uU328+QcY5Vpa+6Jc37gTqLBb7ZQskjNgr9qPqF+Zxs1CtN9MSGuaomwFtHSbrpQSKFR6uunADhy
/3+90Pww2yTnpn0zid+gvVN6Yi9Eawsk3k0T1sX/Vxb/nmrkYsp8eQgA47rdSKKz4CcsbhRlLPYC
vfvUOAnVAwO3D0STHuVZRcqdVSCUzYSxkEV4pXeLWt6a1kbb158WpeSJTZ/f9j08sWlljXQ0Vh5Q
p02hd8wfc5nHkohdQM/x6PlysXFBDqL8KQcVVY65HKdw361K7soCkNz3LCbNShSoRMhG6Q1YKPxu
Ur8dIW8LOATCgpGHRvZZquDeZVXa8t+ro63e6bs8fYkWw4DBcCEj3ZDr8kVP4EPBwkduDS9I2cnQ
wCQOQR2cCxvR+wi10tYCw0/l3k8keicJIi+pIRNtZhWS7aEQLspsig6oLJAcqQc58PnR67pAkheW
vW1w9JDKhWG2w3lFjDPOoc0KCy6EhK4IAXMmzh1A5e20M58hmW/zv+K2ILgOcNbOKO6qNqUpexvI
Xjn2v3dyVL1pMdpgYhi9KQvgRzmylN7f+aABayhT2mioPsiHi9vABKFRTrEAmoJ3EoeGoPloG4m7
4OPWEeOWkh7c91BXsp90bwWlcAwZ8Z6tDhkJQv1RVmTUo7VeJu4FXUMKUGiExYezHPKT5QZ+f+Vt
D1K/70GInFUxa3qNLdVwy0jCnokVq88Jd7u+ukGRDsKXHLYokC9ROjCXpz/2XS8E2XJNJWuiVKaO
6Alty382Jbo3S30mkjkb2mAwyw4R2xDhjT8BhTHM2hFxH4hfMvdhg1cbky+QMwNJ/PLkpWW595qY
eUCHSSRiO8dXIciNG9J1l/4gfqFGRaGyUnpZDrlEsV+PBmBY5ZehqnMVBP6rXpqbl5YUTz5F62vS
DQ4LTyN0UOnXE78YVyeliXtTQ0+0nPcM/vP5OAfJ+HJtHqR9KHYlHkHoJ8r5QXspx5MM6qQoXljL
2qbcr/EOwB4mUgYWvpu18VMJK6MF94Gc8rCqwA9HZWMI82FHfq5N8lmXS/qKqEyt1YUMMizhymJH
9VnpEsXC4V6MFwWQ6c2GkNFgeyxsCrB9JYe3z1kyP0F6nfKtWQRYs5R2zhenbG2zSn4tYwpN76V8
l+cVdMaUMOhiZEllbMDkEGTePgUrrpMr9OSnVXdFBSNpVtXAB0Y6x31mmjbSM5LCgYj9FWl44Sdq
17VhrTOzf3AHX8QGDgQ5tpwkFoHADOML1ed7Clpbfk2w5up/UPaBTowFrI+2dvtblWQ01x/CYtB9
WMeUfEAF00EFsCqcJZXefhEGmtfpTnj8mFbtxndYGmQjVTvWqJfO1tlS0KHY6wGi+cHowyNL/fkn
y1XozKUNkgfqZinyoQ6LgmkUXFqmY7P2HshsRidjKVlXGFmjkAXRRel+vG0VzCdCyyaiOngwulBY
4QhBXBX1a1k5qLkLL6T6U17HgouQoTzlNhKsMkkStRPPpCnE23VhCrCJOmbBqKwAk8VhVXF+HWgT
iUQaAl7pfw7G3+aBffvyEBi9ZEPxaiLW7uHIJubeUEZsNIjdsvTxB6apWSauscKOMdBnMmCXPAV6
HPPjOxLL7xlkhNx6gfcE9HwZnF7N+fnXyj2e8QkgejCAmsfC6MIJVifpR72Q26vroGWH80E5oX8r
TlxR3H21E+Nz+MJkBjDNt9RhfLX9PSJc02RXKGL7ihWEoXUDw0szuWisKwClqGb8ZKwV5ZBiRlfx
ceSXh/wF1ZyKdusbngMsEMFjpraBfAg4koPO1EnnubMOZOyQmBFJGipVU2KhuSTFUuw42jQ75iRo
aWoMn9KanzjDSDSSTac7JSaW16I8CT3C3ljugGqBkp6Luw1Sm1NkdgEsR2y/8N0mB/SlI93ubA5N
YGsUgxaTEjiLs2JgPD7ccgzLJ+VidyCQyTx+/xLbZGSErBipTGbEUFkOvIFVfz7Ftyvw9vGmqx9H
nsyhFp+Q0bjbQe5NvuvJT2ykLQZ/et6EckCUOnAGb1nTu7EG7KWzrUKn794Awu3lllRL5lbT7Ukh
HcxfSrfGsiA/SG/9w7Ht9SDfLm9B34hnzgpFZWtt5x+5IGzR+xCZNgZCkSvBc+PO5Gk/5c/7y4D9
YQtgMeftIBYYR6qhg0NtT5BCh4rNo8qDJ73iFsp88gm4xGj+c7JKxIn+SflC60jASJzSmKb4k01n
Z5DxtPc87VzEWQdip0aiYAsnwZkUegw0JuoB+Rvywo1xPRvRas2Eb2nyKALTG7z4EaJmp31Glv5o
D3lEkjnKPzo82n97Hr5HiLb+1yxA2nZ/QWqKT8LPW4QymFLinOVFFOgasgYIA40a+9N7MSl0O+Q2
ZCEyYAYBzMTH9U6lANjf99vLv8+bAKbzbzN/Kap/+Q6LsrHTQVoGgs2Hey+fe6495GuxeANBT3oX
ESLRk6wOOmZ18kWzRQFzMJGZxjCyyeYCp0iK1x6DVcoqAKAGzE0K/3RJPHpJwmrL6uiSB4zuzBEo
OALmI9fkmQDmixfhGbVGpn1zLcwxmXcQrBhi8D5/W1i5e4UQqgahMNaEB63eb4t9Js4rO+C2jilD
0s1QQAAqw81NQrwuV7ZaUTl4GCxM1B5JhaghlsOpDXJn2gbM0T7R+V3U5R1wdg5/rliCDabc+0Kg
mXHauw63TE6ovugfOnJAgalp5/HznJFZp15dECHclEpaNDavNLnUzGV6Ea4SYtS6BbtGT8dQ1xNC
BqdJa1R+9M5o+S+iYMVyZmg8mSIi4rDiwm8Fr6KALpv/JYdbkQ2Maeqmuc8nb08xeasaE2af2qUL
jHcOpswWcL+LJ+v7uSjJ1hBJLRUtgKdjzrLlbLxLaVA2Wqaabx5O5oFMt9C/jaWBeshJV4bV//zR
iBhmWEJLNm2Ir/vsr2nAgX35ru1SNI9W6ipYbfoBttBo9YSG/YL5LmuoYHChIptjkNm/OfnnDWMo
E6S0PtoQnJKKFp6RVH97HvqCb76KBIuRsYUgnUEFTJ9gie6ML/tT+wgyLWRpAdYQ1oRUw3oaAAeo
uEI6klwxGOm2DJSG6hVZB85NQjd3s4O96nh9AJUXmqWHtkTljUK/t+72QvvgnFtJ1ol5vK7D2I3q
2kT6qJLOkA2iqKmF+BHC+toB/E3j0Yba8A4Wd30E2iOGx9hCZPxDqkVyl6nbF6L5jXL4B8bnyayJ
dR+SWFUq4Do3FFao3NOfwQNjBC75k8rG3cPt6Eo1T8TOxBTTdPIY2+TrFSF2mx9O/PFtMLg6zIg1
pVmgcNS3LZISRDOMaKQjkPOKn2euTsLYag0UG8ljKn7ZJz/KQA7hihG2QQmCvn2F+kXnwsL+fEow
IEIc+g+p8CAEsa+21Rr/l48Q0HXvEkq1hJX+veUwOfZvgIE/jrZPn7Q3mrQ5r4UEGcHubzdZIuqy
hoGI90KNU+iQ3MV5X4mWcbCuNcUBYDVpO0Oj6aTWRQnDmHg0kFrL509BgUeU0k10iiuaiJsvlH6M
IiNwC6x/ht9Pu58X+eWQFRqILisb6Y7Z6nDMVnoEfHgF3aaCLCexIVQivaHfGM70EibDLBUSGFPD
MDPW3jJcJMVO/3eOZ10h07Ic8BqkB2+LV/MyE/4MGpfWNx5HgAYJwN6sbldU36YmdtvtL7D9YxGQ
+1nSyWDCIfmFUMzbxjRGMdwO27iS8rCe7pXyP0c8itzwv54noCrPAoUTbQOZdRHqdcipPTviuWc+
dKv067nPxt6xZM6hNUYHtwWNIpkSWR3xYiOFQVQQiOB2mJJYqp9NJqNXMxIXAnw3acB33po2q6Ha
4TkLkEbD3kXUF4M896X+yipqk49LA8pZAokHaKVX1z3JMw+yIbw6qmU4K3w1egIo+vPd6kTlkist
nPZberDRFzXhQ+hHdvy5og3qhVz2vgh4BMHP6+Ns3vBGPVFMBdXqFYwKy73zpzUlmG3W+Vmhvymf
3aAC8jAIoHbVp5FBgm4TZhGcZBLYqZK0d0dukdrtWAlYRf3w7Kc27rA+J0TpmCL6G5FQjwyFz4p+
EWKEc6lhsAzdFRLb2VLLqONBy/H2rnuM5iCcQcdpBl2amHGkwthYyj50SP19fb1Dx247O3TIOqNj
p3X48j2+AFZCeIA7O69GVliGN+Kw3Ucc6ReF6Q+LHEOf0KYSpMiHsuI5Oyj7tb3LeoqzAmFeT9WA
4oc4/HdbMyzYzgtjcRplrok/QEZJzdyoOxq+yuWuQ3KAHkviprjdUXjsJuZDMDU59+vzzc6OycTk
2ZgpxJKJbtC/WWE9aMx9H4QgM+13DDkes02MwzYKNa2wFKcNfvsSm0I8D2YAioC7zwqCTTp65s+J
hEEcEbaLskhXLRpyCkRAV6myUQSbS1RtyzQG30H7faWoXUVukKmtjS4Cc5kCIWMuB3jzVi3v6wr6
g3W4RiwMJpVW1c276qq8UlPLaZo2o/VsTpcC+lUVcEBOEhjyEvQrMYgdyxiiuzKnd2I3sBrZDWAo
9VQC3eiLiacCpvJCJC+nTvPDiMnshJiwEcZvepc4+ElI9/VBiSw7STO148tB1cY9i5DgOEt0uQNA
RwOZHZWILm5V2JQtsWyyIzpY0TH4ot/5dUHrYoY1C80F3EXRN3jEVASQYSe0VudFzt+i5u6DfJca
wydeOw4JW/En11X4VaHVHUQMe6VwepfRXtylZgUGIiRJk7DdrGq0cACc9nCdZBl+QNp5aBX/fp6L
T9lVM3TGpVpUIKjRZJcCRxS2PeAuX086SLep5JUW4M7StEV61lt48ofdf06Xylos372Ju4bxNXuF
tXpKChSMe5ffXWnRpKKbguKMCKR+2ZDWhjSCbGwkRgQUVIOuzaoiZKR8PPsxxMIg3F24IeVGtcJy
lgnsm2ruri6D1hwM4VdB9xDIUyQBsziWVH/Pe5OsfI7h/03ehWHZGT11RTifY9Ml3vZnJbuTExcC
AP4V2G20xiMFEg1KXlyPcgguRlkm1aIWU79nNQvV7YenEh3AO/9/auLWSZsZd/YtdKBTNyUcbkm4
6PL+rNct055b69gI96JNJgQu9mcT9Qb+cL6IQP63KCpgSiG+niJM2/gJiucpDZf4h1Py6z03Np5u
lGq/6kITpEsdJZI2cycuG1kmgxNrGeHHT/ThU4j9b+OVOfg8TJOHL7dHsWjIYxYcaOwkIZSb3D5X
ycnLKVnjdJ3WynKSQRFpsw0zp32zj+yuYrDSwTNYJ8BTQPvq8gBBEvUEV9E5FqR45rQFIVsw5M6B
KbGsL5P9K9d1i8JmLHFZp+IMMf6XLBqR0jo/FBefvvRxOULqlD3sKqoRs3Garm+jLXOyfg8OxIdd
IsjyYi/yahDC49BWfIc8qq5AarAZNlIgsAQ/AtUV3695T3nWcFNPn6ms+zE5SGXnoJVwRWMZc4a1
cN/w+uB2u/c/ZSPc1Omt2waql5Lxq3hQ2zmLlA0UUQaJz2ZTM4lSKMNyuWxUnvsWckIvf6CLnwEi
hkptPSQuQwTm0FY2BgFfOJ41PexzXn9ZHmGWb9F01Ec1+MZWCOU59qRFAEM3d8WoQLjs+1JPQVPp
Xa4g7hUF+Rd1N5crs1449HlcHnjHLJdJSDaoRTvFTn8s1PegvytHwEpyofEoHgkxXFO6iwP85Pom
v0gkZOnxTf9nsgrPmYcoQjSlojeY3u2MjxhJDqPVhuTNOSnQokC/gEg6sxzvyOTWT1Rx9QlTXpnk
2oa8gcREDqqzGzLPDZEaC5y1dxW++9koZD8+C+QxiHCsaTU4bHFCT9w45w/8fYmOB++DEAs2dKtX
kTdefoArLQios+ULQFPOXi5ZMuXdnGtZdgCfp7ywD6Dv7/cZ/u9hXMtuh7TCS3tnvM9gVKmZo2P2
ULlrbdu5cal2blr6EG59x1ku7hSIleJZcjMoUQxu3/r8lDK6gphcP1JuZkYW0gXs0ps4OtI/paUW
hdOAnZ00uULqPhKsPrprzoezbXk6UsvmoRTwrbS9W+m/wzlesbK6Q60pw9KL5NHMn7Qi9PdRauwQ
seY6AOfwebOxvHpJ+V0D9iM3Zt7Ivxr09ywIXwZFPy/r4yTOivCrY8ptl30U0zE5KBV+E91sgRX0
+lHh+52jR0kAC9AT+25aTbq1j8DUhvSf+2AOtlhobQEkSUBdCyvsBFfPnfqpqsZXGN+jHkWruYZR
fmdGuieVnLz01obJOCXHYLHA2rs2DLuhbwvFI+wVWBBhaHUzU6+xZ2E9JpVXFAfzDNM4zECRslDo
iZ37CPBVbcSCr2JSnS/CUmr0PDDheEz6K3UmfrqXgtba/m6SE0O8jgoyWw2Ur1+I+u6o6RCWYG/E
ZTiilTF0iq34OB1gW9XULETXHnQms2EHUokEMpuIb/WOr7a8VJsRB1uf4CdEVC1VridSiAMKlU2y
3/ue0ArI4x+4lNZ29SBGvHGtr/VsgvoohXf9aVjAE01wgiSVevL/3FkJ7G2o5IioPkA0oxBVx/vo
/eUjY1HwMq5uu6xe9MeZwM6ovBxRbtkA4D4qeedlZ4UpEy2ZTbywugRHrwZbA01rHwLTK+3Lzvo1
AdhWzHNUOoA7fo75i5zdOQm90I2SrMNuCJYWtdmjr+sb9YBpDZxqMHxXjw9WYV7393r18fjzg2QJ
oD5nnER5wM1zIAWI8sIlYC+1cMVrqbYbZgJ4SV9PVvIzS7CEe1wdQjDgKI5GZu//jp0Ufq0xlz4w
581vuvY4tiUK5WfOxVSa5V9qdVC/BpW01uSMB9yp+Y7JZo6bcFAYQnn8tQFPbO19HiScPFtz7lNW
MQNM2vzLPFQlHhce9JNQYQFdwtQDiSr8xX297LDa6dIeTF/wTX91TYHicjg3fEDo1/KRfC3MR+cK
yn7Nk21+SjH5My0S6h+RqjN8VJJKwyr52ceOpxoc0US37WjzIOht7971jodNFaqwh+4lLAmlZGpl
n/x9hGjzr0TmPGwA+PdUT0CK7+UYztX5pLuiZnfj8K3WtVHoKhioDa7iukqqXAWAL1xYao0WLxUN
gsDnfpbTmLxGC5vUjCKBEzKVnyQESL2XzKE/dcZOnGbdpL0a21kXMZzkuQPYT2sWHsq1Iyv1rhtP
iN3zz+kdCY5ghSyGN5aMaeFZCSvPfyMv/Ci3o+usiuD8Lb+E4faHHgkrPcdy473NQFXvN9Nkq/xb
L7KxeBW6a2ajbsMNJIbACScmyeaA5QttEsIjXZpUDSmVjbaQyhGABzlkdNGoRHXRTJ8QcIDsJXAP
j74E22ijmPRIPqAwbJKwiKv+Oz7WWVAWzkf4NXnq5HDNSFnnedh2OUEaA7yq7fw0bJr4UrTwaLpY
pL31u16sxJC8CtGDP03+w3XKRhk99JKxE1KmP+iY57Ct4sGrJ1c/ZBuN/SIKp9N/xxfT4gWS1zoO
2Ea+HA6Yq0Ex2GLvdY1LztrfamXscDiajvb6YSw4OfP5Gt/Rr6+ewGMBchRROKihtcXFSLA+ewf1
e/cmXtplvNJlA18uNz7mk0n9+ShsqBxYoH4BlQXHgWb3/30PqrQd3C5AbYciWtCmqLUMc3yORkU/
Rcuf9Tn0J2XRfR7oO2vEN0G1Zyd+DEgWpfTpOMu+6sA51JhmWpW0XhTvFyx5js440DSQgH7fFV9n
P176dm9WCwlrOFvM9DseZ8Os5USf34qJUeQTGG/eIP+NE2pgDeO/vLPhxnuXTBhaQScHnEq6EZya
TGYPFI/N/ORgGAdEjhogUjc0sa6PTOGJL0fgTaWW+4HB8e0jXIYmhZ5GOw6JlRytSadQp4UxYeLK
jC0Xe7oBxa/bBdZmU56IgeSKCOsLjgkHLtkjuYIeF47XJX9I8bckP3AZKsx7VYBcbkjVpD4rJjbI
TZFMoBHih8CxOtTEtq4uD3TSPUqhWlYS2TeFTRIL4L5zjY4q0bScEintOVNt8AvYW2R79Q7ab93G
qyEa2r82iqF9zD/RkLI4fm74IJbTs5SbffmNe3UW3S2dTuXT14rvAOnEDQ9mTfG9IH9nb64oVgCm
Sy42Hkp5di0DLJ+pIMXKZ6B/3w1HjgHcdCEEs7fmCsmVKWb3ZVd7UOFM0iHlo83DfIuJScV05Df6
HxYQkqluD1mbN0ZBFhPCgXJqyDdyvBVLlN/HICevcBBXufkgIAc14YRhQwifmQa3KWbBAUzXsY/l
B04z39uUKODSM80+WEsmIoPwyGnjgcZQgkrFLhysAVFXECJcLT7Mjl92TuTNaC3Xo902QkB2AX+l
KsBnRktQR5L8upICvI+BRSnw/ZC79d+IMCuV4wIKkFNIcUI9EteqzKafyNylPbcHMaGn7mVXDJjH
d6MMcbA9dzOm/gzNRd2raLdQRVKKxpCmqrJ3Pk5427LmFhEwOTsz9zaQScEGck8qxCRUcdcB+mkU
7OZ0NJRk1/Dk7LZrzjQeaxhjpqDNmBNtsKDGfw16RzNjg9R3S8TSSOYvM1O+9IbnukrF7ngEXBkT
YVyvPB1tK6RmnNz6GgNtDxHSMVaAiW9CoIG06WB/WNtPSDM/YQgVYpIIZXhL2xwi/zxEAqaRcM0P
AbNAF5Pmv3vQQ1FLo1flHqX6mVscW9vpO5a5ewCXsXQY7xUW4wJclLLXq+SP+kt0WFcbzh+9J1eB
IPpy93Lm8Hiu6vaMk32Zlrva3PQOMoMUG4ry/jHjBLHyudzUdHByWA2oM2zjfuol/Em1q7LedyQz
SXgKkh63C9LolH+qmiSzbB/AMoLfhd3nYFJcGRCu/RWSV79Icy0iPktyqKhsqsAryLI/Eac148a0
knvLWnjBnDXlorHIWpUkQx1Wrk/RKpEQFxGI6FqKxlOL27jzqG7WkVZP0G87wLYM7AFUbhKScs25
/Hpkz8AP0Z+S7L9TGSUg1VHqaVgGD0fEFT2Smesz9svmy+pUhUiLPk2VZemOJjn3PjM9Sm352QkU
tv5GJ6i8JssCJPHFgo66voVAOgsyKxD3VMCY+BrEuJT6ApVnyfBRq1QyoGSdoPHRS4QkzYwNc3Gw
tgTAXuiRnMFdak77D0+B2aUGGS4UuwNlpgFBV/XowsTlJ9rywc9VoWFmkrAL3nDZHJ3QA+zZAjHV
Fiy0N+5OQyZIiXt9w7O1t7dFcEta3X98r/qe1YCzBrS3XKHSSzND9Ha3ayHtNxMXWIjxwdaq9MBf
fffLtuolPaOC4q6RloWp6JcSaL9b1zOtjlif/c3wqx2XA/aGMjsmLOu+n9+4C1uYbt42GnulQot2
6jVWIaf43FOMVY5SPSUFMvN7G9p0R480+SLEMC3Y9JOu5rPDHTDwqiUrPalZdud1QLQIFrJYlE1/
XwETJdIezQFuLze5PQjR/gP88AfEXU6+Kb3ObFUVv6oES2HBUeFEUQqkFsJWi6dcZv5TYa+IdF9g
AorAED38EmrZpG2XupdeZqCmhNa7CSEN3qb+82RBFJ/YPxdQByT3F6nYJNmSwG4jOE75Jr9cxM35
vJueRxZPYIyZv7ngU5yeBq20DhCNFcHLZA0GTEX5f4J0rXfebbv/05yh62Jt/ZHQ7EOQpgY5moKX
yGlTSXoYpKiaQSIP+vFTW7zDS7NEdbnYOvHl/KKW/s0I/UFMrhVEGWXK9Iem1T4qwhzvF6xEOhfB
k+xYMMFiOvxpN5RvqrLqnhZrrm+Q39Nejq3ngnYCAZ/ddrALS9YG6KjqNumSzvSdWxyb8wQaLS+b
PieAyRi6GCWioljjxVaYfEklvCJpOtHXrnknzNT2PwjwRW05egXOWFgx1vbzsZd1P8xXlULfQtSo
olM47p8KiXzShjARSoX8Ul64UxIGbfZTxh8gu5iCN+uAhburgpI4L1FZzzOQEs8y6s8W8tboibXb
Vdwcd96qVE63lXLhF8QfV7VOVOiFfg4UHaqeaFpy11dsv1+P5iMIa9Q5s0T/RGj2IKtTcM/5tphM
l6L3BO4qNajCFkDIUNGy5h0cD5ljIDEQ0z5ouzIIhGwXnufUEcn2ou+Phm2eXiXGlGKjbeyi8Tc9
5ceBVn3WFj59qJKep7zPCLvvmexYv9mBIu7NymjpIr8OmzrXmDHWfPaf+AQ/G1WApLAXHR3yRGjE
bBZ4RL91DYbO7/bhIhX7iSJs1YVwsDYcdR96T/OnYwK8hfNje/G9MRoZ1e8xY7cUTvxEevOlppAQ
HxqxeDsdQqM+mZsQNv3hXFhpwB35E3jwnhXd+RPUoQmhw30f6J3YD4ulyiYhuknHixEkiQLVb42W
eKGGWpp0sMVw62pUtthOeOP2Z1HUDsFEzFfcoKDIt3bLH3WyzPttI9aY572Hz15wxEXafFgFHMyo
6ZO7SioGRakc3kFRjquSuXwbG+xkyzSI58dBKxXrg5j68iL8E90A1I8vw27Ir5NFoqrGcZW35KyQ
ehDGrRw/WYACZzyNYCb0Zr7HHe96GNv/WUdZxKbqbfj4Vh0q6MsTjl7CsMdtmnerDWZK64ATYrUq
hajxSEZqbn7lJf9LK3NVocBpAs+Ky85qjdybV/V/rISfJKTbJyMSBxUlnaaC3/vypX6QGq4hQkKD
rb8eLtN4A6J6G6pOXa7Fy3GHRwOurU4Og1ciwwTQCAUsqp2cNVW4onqxTUdzRfU+g3sqXV6FENLV
QXaqAShjMh0yxIJxsv4phOxXQwaAdVua/x0LLHSe0nO63yWxyMfSCGHMEfg810DXEI0o2h5v8ev4
TUemmcyJmI6ksuFAimJFMCaswLFRi/4wdvjTGawQqYqqYVxfoK5QREcK5/OBb08+fyqrEhqV1QSx
Mc3GN6LdIwV0gEOqv/qioOGYxLaGIQ1KuBFwrHTK+F3AiHlJ9lJAcxEQ76ZRfelWWH6NLh7+z/JF
7PZZ8I6x+sxHg24w5TKXJ7HpSJTL1gRBIf0oLyX5Zk3DMG9o+K3bvwo4P/ZN9hsqJHS0vfSwvs1r
ImrQXT1gMYTEtI82ZMsss2ppWKIfmabxbUdhyKzykrKIUfYQUms1RUTLCrwqsXqe9q/O+C4kXqiB
wi4Q4srsXcKJzWF2h3VX5SkBqiTL0ltr0TzHS7hc+EGwwlDz8Em6w7Ooe5C9cRaaqwMVHFVAqBIb
HEY//QBV6j+Uj2DZooz1H5zAq4DQGmmTJ3/zu3eq82cJsN9jVOoqVN88ttP52tTMjogWskJ1eusu
tMJWVKcUKKqIJ7l2iTvRumKMsiIkDJl/e/oh0Bltau63Itx+fTk0YJ5QbDG8m4OdN7rAv2TehMtS
V5SwgLgFzyT8lVEUZQxft+Z+T0vMSJyZS1nA+tm28UAukJ8pELNKoimeEYNGDk7pZu4+r1HWURRd
YBc0QUiw+3vtxKJjxpM/pbmeRdvGAvA/MPWQfsvLtg8VT82w/warzCW9u3zN7DQxPEbElGiRnI6P
imRV+vrWE73RKoLWEkQsEGV5BMZFYPhpmVGr17m+pSDetNVBfZpxK0Ks6s/Xa/6j5Foo+HPswuj7
JAvEt2UPE0DkeVWomHC+vmQ8e3G+uxcLnnpdMODCa4lCmDpsX+3M1y6+JElCaG6CW3JAOfdPxiqF
YmBbDEdWuCWSRG0GunmHSePCUa5eMtoBuT9162FxBTf3xd7oQ2i8jQMKVB6QBp/Cks0C8X6N0DF3
q9VY9gtO4VmvsnaWBFjUkn5+JBFdEN0tSYA0Ll2ow3C2i9FxUCx/MDFf8yT0GhnRvEWrihKUYXKm
XgUFLQIbEv8k6S/vWbGdUGhTpS1zzxznmTaB4XUis1mzZkU3CJHIW13Jep8D/7suU8jp9NUs0Mt/
nV5SWnzTogRUQ0u68sE/59zMIBPYWbAO+NQcKoqY7xKwNnx0AP5PVzEPsIYLVvHOsk3l9An3M1Jv
H3RIpnJZdXma2VG9LJOPaQRuiGALCEFXFwHuyV2prOQ7s23Nqjn2xNMuttgwWZnoAhOlp1xaKrqf
JqkDp0dCpTKu5hFPfZk1kGYugvkEZORkg4Ppdz6DbSYm/cE6M+QqCZFbH+j7AFrMoxqZ3S4eR/9X
PRPbB4X81CfwNgoEmeT31esPdY4/1bcALIuNMyISEKogJmDOYLp3FqQGjjnySSSHroUxMx/kWULo
UB2MoPHeXUwsYrJIHXg4lDcLf2ttyUYtMkQXgqhPqBKgEDBr4HW0UaXb0fMwfUZEYYphfrr8xQ+l
0bhkip285XNsowUqrVjWDAf4mmUloonPMBI34bVYCgAf7hD1E4nqTMnD0+iacnk9nd9BL36AaaHH
T6NFJtlpCI3YG/xMIz1O5/gqkzHrga26onuzOZUhVH1x9t4Cg9CXTAMD6lkfFFBojwIJKLhuAHnD
28aEAbMxC9jYuC1A6BIRCXDe2rOYwfEBK7MybtZUmTZfZ/DQq/WVdmk40fmOjbWyughnMQfWkKP2
HuBD+bV9JKzPg2eOaPrgeykCNchV8UnqnSFaPCfGLrOADV8emoSpBe610Eu/bec0vy/7RnabOupa
xMkPjeR5/X7wUpX35hM7Ux9LV6RB4PfHimgAqQDmKrbxTJml5V1CshlVKhtCstkfeTeIYwpIyHCy
DLZa/I+E4DSTABrG4PgEYjRRP8gHq4KBtO5U87RsEuoTo6gX+6wuNnLsFne7vvDAtchluvD84meO
qEN+QFYBu2hccfxLdy3IOQrekisvRMTCYj5GT1ntMPQMx/YTDmJy5JSgVC+SReMPMkjvI6Z4qaxm
Byn4HtUAFKEN2C8xO/sEhX+9EOEed0RYKsUqXztKu6helhW3DwXYwLBlgEDe5oLgAxeQ0JsDHW+f
ixtUCFPe38/O35sS6DC3bk5qvZ0n9Id4QLNk5HUlI2+ziFhH+Zige8w7fNSq0o2wqkbQC33Ho73K
3NQcfxw0rXxYvWqrv5iz6hspbnkLGbhvfivieCduvYR9WzBSLuhv7ZUTD0yYQ+jGuX3YJW41jv0h
HpeyVHQLM09keFZ7EytDhOAnza5XPW1MkT02Jwg39VMXXf+/Dg5enlC/yOGG1ySa5pSZuq+4ngmF
JNBjabY0s4DneqVpsPxZDiNGio/cx6M/cVVczyy1XDoihri27ysYP/8lVCszr361Kg7+BhPm0zV9
yUgyVJy1YHQFJaLUSVOt7zzLg6CDbHdFn7cLW45KjyZG0zr/MunKVIEwWfcGUwS+03EpQBpxqWdC
6STLUUwJwudiW11UYRXFliDTW2F0W+izXwf1MmVIfn/G1K4h8CuIQRKUv7TLDlgwbj8baJXl2/XW
Lw/ahTv/KfmZM+55Qso0J5kOrcBXTNdDRxEuSv+49IctQe5bYVCxe4SDABNRa+0u0YP62DMEkoMs
urPPCIwfMBFGzdYcdvNrb8KczgWEXmfpkAg7CaX3qrhQvH0OnGQcHAmStHP+BmnZJ1BVQm4L5GNp
dodtCafJPbhABlvS90NyvSVgPKKaUbLvtDQU0QYgQOT7jPG35XcnreYDhFHjwetMdlU+5Gg/ElMn
1fUKFa/kIimfiO/9/ld6zBFkiU9X4NkWF/831dG9xtxSgNCz+kY1q//GxZfeTv6pfYV6OJkOAb4K
ner7nAPAadr758FC1E34Qu6bhgNyz9Es9EOM3CuUmiIkyToe4Zpa+qFaXMxJXACz6nmZx72Xo1iY
CwoSeaQau3PVK3lHmyItYsxR51JEA6wxR3qagiRHf2Aw8FQApbJJ8joREnrq7n8lsjgpHAkHJYwx
nATjfu3J+S3W+nRPFpbwE+B/1tUCnrJu60csAbhDf6Klq/o8vEph70E9B/Azvskcxapslid6XFeI
LQJe2E4AGT6U4OqiUztCyUg1dhSuw/9RYhjBa4+CspHDOdsQGKmM+xUmYhHq6mmPGX7637Wc+FXM
gnp+BdS/nHROzgiQspfW2ERq6aRPh6sj2MBW4Vp6zYnetXtpeUbRRdICvWmvc1+0e2OMA7PHv0ud
47UPkdMdyAtHkFoqTgAVselNA/DFjJmSA987RlF8mzGjvMsOIM1FO6ozj4CDR83uJu7hhvfpWh/B
6QBcHIXGN470mmWT8JVhF22iN8xM4MD0XshNj6dbcCI8OCluGClv3dfFJQOqYFIJqXhDcXhhphhQ
FmOKAEeKZfeBkPdf2JPEWS2vH5I5ebZRMX8V6VNWE9zDShxSgiHM831lI1uVTXAobSivy5Bw5blc
IZ9ca0nx8yJXWwKbQ8Wpn2E7FEth0OywK3RWYV0bZ4ercrI5raSPyog55K+FBn1NOuGlUWTpijWL
y4dAyR6gFW73xhB4vwC30dYQWOJLASS/epLnHDEzW28eQ7FVu0sDcd40dCppuuqC5Q7DqNXrJFqY
vPG6WrWO90aVaB48EFaJZdoHxvteeQ84tpI/ni8pabNKmNu8Rh75dpLRNtXrMNj0FhwavQ6Sq779
jyfbx6To9t28i7ovX5SoCtFJF+2t+kqP2hJAW2SrDCQZLmAzH6SxZhk2iVcfOyv1gBAH5gViTo7O
F+2fzuL2VpON2cHAi8sYgC2BWUmLeQ2jSmYsslaJetHGepTBz31qvioyfB8bywx9qPLoZ3hip/MV
g47cDn46K0F5z44ysAUdn86FvThEhMLhyLwGpFyLsA/7cOzqBvzD91f8R1y42bA/O5LzsF/QX915
yY50XnP64AVuPcRUXxsne9VrL0IzvatoTJROYbPFqSAhP2WJF/WrF+/w+IFuIkw1YoQsp9qWNSu6
/p++lLzUxtloMdgbzvCSWKJNzAIJJqeX1EGsOnAiXlq16mOIXpDSwjyjPzyvEe/GXv/2ZlN15Qzx
qcLhtRj108z1CiwvvXT7eWjv997CQ7+WHsPqWzxwGa5fHlkIs03gryjnTAUy5J3zJJdVd7FxGXN0
9asKhR9ndlmoV4wdbxz7UNKBh8Vlw5iqLz8QhqJXZPI4Vc7f3telSCJatnJyisJxeI/eo90bffYT
efdM21W7qxlhDkwP1ajBSu7Lr4dGZ1zk45sitY0wvFe3ECpt3Q4KNGI3QNLG52NWHD5gs+7tNwBp
AFTG3BgDaAcuxFmDx9JziKApsg1Bsu2h9ATdOurZpSbOPrSpQLDnpOgxaDXNol6FNO9+NWIoeljk
6X/KfKz5ndHhUrYiTOy+fs8YW+rbeIVNYNjNmFHoSOHLNBMHsaiqeqIdWLE5aAeU5Wv3ffozLSeX
a5fBALoFLyIHMSUnkhrJQM4bg4bEuI/xtoNShZYGcsB0edd/IRqfjSTwnTnVnmeLBQ+v9y9bhAew
E8EF749FZSM8vkg1/9JZcSYB1d7cZXiBVG8R0dVSUYg/PcdwpeMACDR5DsO9lGJZ/0m1DPMpqHtS
AoDGifVZrktG9evPORHQg68ox9sk+xRRyq9i7tgdWxsG9bqvMwm0petc+l1hZmZtvo/eogsuUcGD
+DM9qPnYtxyoKmgdrXLBq+uryf6tiOBqHXaGw4bM/NNezCSGnyLcuFFjiMBhpo6xM3q1eQ7nfqIc
kdLKWT1wg02++vNWWJ2jQtupCzFYYE/g0ks10tw6gz1ej0uAZvjARF7GVu5wB4q/bBFMcDdqTXIT
byDT3FOtuQWe7c2r/czL0boH3Mta873IJqnXaQ7Z2hbmGB4hAg9VvNG+Qj225N27WxPoD3F586aL
ITDQMoqREMRyGyZZxTXjMzkFlMdaFinKvv1fm4FkgDi+VVi1MTOa4KGO3wXu5uZxSg49VPaH7Byb
AYUQRZlU+tozfPz9WbF339xuK6Hw1Qd0KLnhaY6rWoQVxm+wpq1ycikt8wL/px1XWmmRXjTVKDIJ
toNlAhSlbWSI+0/8h0w5Q+ryfgcYirWv5KX2n2nJJnwFFeHgy9lSddwulbKfmHtQWe6QmxBoQpe3
c5wdWXzshoKE4pi+PMuKsQINj7EoO4AeYByZ1ZZNjtZCt2yX0cXgm/jJOpkE/bQ5UyKrqC+gdp2r
355NIzqxrR67XuP55yhhFOwziihkTsV86hDap0QnhTrPkXCwGk/qUgCdnbOU7tSZfMTl6E+FcRB0
338c+RHX15d4tuBPaSqq+yEiJ1uf/cYcA3iC9Wz3G+UXa8XKdHm61Eq8xLg6tf5VY8MD7L8xLfsv
2YhMgU1IXJ9PTtPMff04/N2U2tWftljwrnAnYZrbRvxw0JJegKz0LVitLcdgcJGO9B0N8GsvXc0X
X/7oHSAm6Zmghw4UIckIv4NzOyrWnmrOT3qAMxDJggLMFp8i8Z3D6v/xBdIFVSMre+PmLM2WulSI
h4R4ZvJxThje9JkcCY5grDHbe5T/y4b/Ewi/+J1vN10xJES2kNBi6UovEf/WYoyNnRPK7sg+Gm1C
L9cY1gtgWDfMaWwGsF9Dra7ztw6Ax9Byg/K4BBOdsDSbkPCu3OKnlcmd4IJ1lFtXlRQk/OEFqcAV
eyZ5BfxQG0m6ls9vbypTbxHae9IsaeZdCanda15+xUqBLInyGohY/u1QptcU8rSrh48HWverN5GM
zV3nkgAvXc9umSIExPg28pzmE6reaj4zOMqXos3xjzJROPZPhNE1CmMgwFrzOws8zlyLI7PF0wuz
+Ozs7begucB1wx1gEudeHSvO1HDEX1ECjj74C7rqD6Th7mL+fypaZu5kySKXUf08MtDCSV+Oegri
9FmWULVfm52sPtgLNeiIY+6VuhA23Ckpai0yIAyNI9RLIY9RIPxCyiOsBMBPVfnsb+Z1nqJfhBbW
SZH8MWsjvDGmHG+RtB3y25LsE4R5Q4NA1U7V0MjJRbqKPJvUInpthpeJ06O6P6924wfeBdj43jDf
Nn3nSa3n3IxTvQwX2hhYRXIErNswpFUtlZzS2LBBPoxNeJgloxYiQmf5mjdDJxjGcDXkscgwojqB
NAxH6V03gs6WVebTCpfW2pvC9l4oe0Le4f42OKtiKiUyue7aq/lCcYRYpwxP8uum3Q/z2fCM/yBp
GaM9I0fek5iAEeLTNT/pb7ZYQm9HZGju187Z73/O9Aq6igFTXhcazmSJmHh/+qMB3a4u7GYOZA5N
iQfyTFOq5VSzd0yGFeWWPXRGk0c5ofvJS8Bdl7rhg1FOBT50uA9ryoVFTvMHBEtz3lYhOzpyihJS
58Dl3u8GSBBampuEHStpSPVhdtQzlocgCnEcwnMt/YdEeaI7qCONmyAA1VxuPUDXmusFLykhfEyN
HBaQPL7SI4GeEGh8/hFDan8r77up52ZnymGr4YQZCbHUNiR3mzvhkvwzgBsi+a2aFKcJkfirh8UB
sR+AiVGXny0IRHNgm86Zc5SX985A8CH29QI25IBsUdjwR5SkC0lQlF1e+2C9a+RIaMr4D4YVfyZg
eGcryjvNrkjmDueZPRcrKUiK834nai4dYVMxEhCtHRuQC5EnKO5tuUICaBBM1IrSoVw7F2Wz+6v1
dRYljdmp27sEB6iNVXXYRr/6zN21EE1hWbQJLpaz6lsQbO1jh8qIXerbcU0lV/NYiSLtF2FYuxWN
jLitne5K7N74kVwPrNkg+i36kOFjeSZMGzZVvhoV3txu6Uey+50WI444p1PkW6tLq543Jj8Jh5rJ
LvKJER2u526MiTT/YK1Dulu/UCBkjkQx7amx//LedxP4sYRwXTC/3YMS1mrrG4OVNsf1pHF8KhYm
FUT3kFvf38LI7D1dAJ59SrpACDhjf/MvuUryca3Ew9lf/Fr9VfwJFBo4cfqhQ45KC485LO9odoVx
KNlMsOQXjmP3bq8xJscZFCq3CJolk4NSwC25bCN84LUZGKOHvNF4JYuetzvOYLts1H/cSG4u8/8t
zviETLGtjgIXRvkHx0lTG6AjKMwHtHRexnnL2No40Ox1WzXbvCBLHjmf3MNo6+miS2HrHZGmsuUB
t4vumEjcTUMkjLSKX6mk6DcPORVI3sC1a/01sEmXuP1Hw2fiBqfSKWQmV9Ef3MwzjYAWdVFtbnvV
J0kRdbmaRIvaBEsm4wZFMlGfkfv2ZW0+gVs9UFEDhdJ8Tt/E8FGT0MYPhdFlSZGasTfPX62TbMld
t0ebQ5zSatwemIuYhpXxPMadBWGu1UaKUzNOBov6XHgXWWjEihX59EtgYvLmtjqo2CntylNNSbKV
HkZdYybAWJHGiC4woFy6AdkxdCZa3gdf2svpoLfQ/0WarIagReJ6YZjKZ2m/xdQaVQFKO1+d+REZ
81VxcAKxYZ1PYIB91Jk8tL324PXwCiIZOWwuoccTNKNgwPFQs+Yfdlt4DW9c9LgAif1ZR0gxHkmC
YvjbHA07IcWbfI+ihKIldRzD6ROfx3ad+xeMHRPv24GwnP8Sv6SB+K/pOLeN2FZdLQAxMWxhwJal
bg3GSane+qJHjzZWwB57QPdNq8qNZFeWPBb/cRD/wAUlTwpjuZwI42wSaJA6uK3MuAQ50o5zF8s6
BhriG5NWU0kkrFcTO4kssxKgKpzTMVyWteuHe1M+3KuzZs/mB93zJH2EpthWKW5TLewURKwlG/2M
tUQR8tewhgbB1pLKsGc2uMoOELOhcMkCHidBXgew/0Mb+dw8Dm0AfA1aJ1Jlkqbwq3JWb2Fx7JVv
RAiFa7A3I5zDe5ytfQfHfexaHfQ1uXMC5EmW7lgqDr4Th3KSMUpuwzGTAAidwrjBzFG+KadltCxd
vTqrXgHKMY3qtBLF9J8n24pIagtMmFb11uCe2Oynu6Pne8vIXXl2xRivnD0AfojSmgchF87bgbAu
LsXET0/DuHw6Dr5c0WmEC5/fgnIAPBk+xHzQTau57OkG7rbJhC9nK2LJe+J816R8uBQ+tD4JJ2ot
jENLaY+Km+uCQkss2+7xyThYXdu8aRgbQdW8sH/x7Nd3oSbhm4djpbXBJXR2GQcwFkEu0KMCg2Jh
0FQwTuNHWj72mzLgZ6eyWwyh5oz+jjY6/ZvhGFnd8E9NTPXHjRs7YFcJf72BH252OMw6Y83n7KH1
fxcSB7d49ymD5tCfigmP/pjG5Xo18CzExL+lOQOqmBEV/wt8EersXsI+yEyBqObsz50Qd3/Uj4oQ
+YiIJVYjFkPR6dkLzVc+vk6c/zwaRmtNydnoMoanVQGb8KHYhTKQHO6oaosVGPPOSXTyBvuBm96X
LQIFakoh3w6I3r4aPW/nfxLbC2t7LJUOkZm0nQ6CRB9J1MSG7odE04wFVrByGTbc/z85b9mqGIZa
Rv6d0eLdutwgeGAlu/WEc+E5Nkozw8KiBQnoENunvvoDTcA1+UOKxNSQKzPcTF4r7htIV0bPCLKP
o2M92fouzuzCWjBv/oPThXqHrjNmXQicDQT/1VgWdCMfhHPWAE/beBbJZ0IuITe8TT0k6avgOe3L
l8pokBnRzxgcTRMkBsb5XXvEoDRM/JO6ef0pMFfAXntk+icP0DBaLgEdkn68dn78jNlQsT3mvxBg
4DtPtPlrPWSRWgfL5svUz//DiHTcCXsPB68HSCegjfVLa/w8Zl0PoBNuJ3m73Aa/xDYAC0WliENQ
rAoMCFE4Nz+nSvFkwaeiKYjmIE/fTjwmRytXI8c3SNf6SO2PC9rzQPwWh6OovenGymBfF8i2vZoR
kabnrO8lcED2Fm/B6jTdfERfQcGk3aPOSTvABjvEgRFb/7q3K6+9AaPURp+walE6k8B4ccCQPvYO
7TOUP+P0NrIaN01Dumpfwpz9KHnvqTNphnywTcFOLfrH6B+5wzMoe8YwDSB4BWFVHxp5nKwx2Fzv
x/wEV68yBxQa6Zsw2rPWeebMDCy4uJeb2PHEYGBWouSKeULHbytZOiIU4d88d4z+JSJnyfbYm7DW
RE6W9xmeqX44JRm8t7nLf+Tybc7o9ox0wQlWCwjIn3GLvlFmAiDIeoQzX/nUGm0nZYn2ulz/EdUk
oohJOGSB+1oxF2m4nkfSSDfe0c4wY0yPH9AaIb3iocCs5AjmYnd3GvGdsOSH8NLsepuLN2J6uBrd
slCzPFphydAvz/mgyUe+hy+cDryW9kZshllfLyb7p1GLKboihKkhT0XnHLJZzscsH7eZgxgve5Qj
0dlXMCP90aKjg5eRJcGi82L7mMaavGu68OQl1pShCPq5RZsKDkiBWiSDrWmbsj0WrynejfY474kY
yPocxcAqawJ8WeF8lGUxpELFFIRGkewiQc3J1YzYYYDXmm8up32cI/d1HFi9O8XGKucQVDURMrLP
64mt9rsCW7qX86TsAXBqWGNWmn7K/9J68C/I+ixStzHElO262J2iMtBcW8b9Ucib9yoI3NF9oi19
+CYM6MNQfbnA3ICcXNcCSCMZ91jYYO18wRHe6J8G9GbusS2WYr+fSWbdK4bwEoP1Nhh+gSSrBeiI
0DyHxBzWt4bNGwigmC/TRRUzCYymX3FvY30KSBFcUf1uhQLcWVW/REI8AXPo97Ey8R5kRzWrTzlR
Oj3dQoVtrDsWDXJ7lPXHGuPLSoNOos0tWOwvryuB5qoEKd0Gtl3oqTJhsRHcJb8XkRTSCmJjF9wh
HhxD58SuIVVugul/2WRNxHU5lmtJy6sLgxs3EWs3JiqcnORbqtTI8Cq+xCHOLXyYNd7GkjqAubYQ
Y2ezayQWByd5RFI0noslD6ycx6Vai6983J4jgIT2sWCfkQgVdkK+L1EmwyB8uaDkJyT6Xlo3Vbiw
dTmgmu3eokaibEVQTAPiRalX98VxSF4WsQ8ahgCSdCXBe+zXmW0qC+78EX2V57utRlrOkDzqTL5C
Nazw5L+luIdTECdPc9mvbazyyarv4RU1GzXe4D+2Soivim9r1Kl2lACYQs/ycj9wTwq9/6bImLOQ
cQhDeaQ1ZlKaSalY7noyJpFvy9B3cDF4qI+hL9RSxZjKTWaW0in/BOmKGt9QKLK432AAmFp1Bcyu
Vh3HYyzFNCpdz5FF7OkWjdCTUJqP+3ARhe9o33PRwV08eetsPRQZaTzG27vb5XS6zjEgazko+4+Q
nyJ7MKSaU3dHIZi63mWzVNS6T1GXKSi2RjqKu75qV+xGtDjNYsfzCO2ZHwVvXRYtTNhXakEdbC8U
N9yorynuaRueFgy/emI+TQyFgf2NNQJGausFOeA45sJDOsQXTJqN7MF/z2amypZ37USATDbBGyeq
DIGSqe/w2Uaw8/dzQWFeIjmqq8TqyIFqoGRgrOBBhp44BdElBmtBgw8uxOD8AW2qJe/SAa3K/rc/
dpiksRdjgs3rN/IRcmC2zQqe6AmC5K76lDNxeyz7tf4OB0fnYltUm8m2PxB6akHQljLI6ykY1SSL
3rOREe/dwUSto7+XUGuYO5blCMxvl+7GPDgPFGUv3sA4sYEM4kkNygJ0snfsZw66DnB/wVrR62GX
K1NdAZTLNiOct991M4ZD+Bp8hXGRjCw2UGnR/S7g6T2mP+AjjETlnaZluDtUKAKr5WMuQBnhho+u
cZgyfMa3k8cJKw7hVjp+qmVdK23Nz2BSAkVHPekSSIpTaRWLlC3hQCVmuntHlj1QsnzNjyccnMfZ
R1I1cHCa7kcbp7q+SGxiEkBFRDRU6QbqCN/ByqXqWGaH3SECro9FSmanxdCGyj44n8MGHpBp1uKj
Y7dWenOGmSGm9PHCFyzxS+avfqm7twMy33P7RCdBaBKlumHF5u8mKyuBbd1NXL261DuXzb42qytE
Nw29dCRuKnSTjofT34hJcGfEjiaslIOfbLbfSTUCOIKFJLsqK0NS6cEZAj8WQiq8YOy7hnZeItgw
YrcYxG/hIoc8kN3wSkblNaotNWOFESZ4hIAHRrETwXECaRT7OQOoi6t2HhRBzUPgPnEUuPKuXcPQ
urhJFrMnvdHpe4VJZj0Jn7B8RXWSbYCDKabOh2ex8OJQM7ldLjDks98ATpmporfTkjRM64+B2NKs
cVbAqMDxneiWXFoiY+M4PNizQawv9qrMz1rC5uDcGge/oIuTDim/fSZPqeXCYwog/kh8ln1BmTCC
R8mSnQk/SoRMavxZKVIoZKLHO+bHkA2QP7Jxpy4OF8efPJLX4qt9YCzGzMd22B66iszSksiubREs
WLBsgTIEFoxL15wLcRgMzFfyzSL59WayQHUW98arg0hUvwhP/1Der2q+srLSzvDEWhp4BNlKAgBO
zidPioTHaFrxeNFr4sWNNgXlUtrF99VtvzujbWqh9WYIJ6XbX19aUAB590KeH7+qRp8K5z9pKjkM
+IUAJpfOG/WWKEBzLIBidKnL30wQU+bGkhwFj19lmJJhukB8K0P5YeaqixxERLHahwwJpY1TqSsE
3ETBE6yO5/1mQxp4+E/jDX1JInp0Camr+oAxB0jXBBwCnnn1vuYH6R+6V4WTrpCMDoRBAESy614H
l9odMv06z9DIzGt7u+iedBMmtWnxWzQNt5JEDYjLNa6djeEtlR80zN2PoAf5tXVjUZayaKKUQQKE
bR1jYEEWsk+tf+P5W4JIy72TXDAd3Lxy0BYvpJbeyWAqYITk7EsNozbPxymmMsvaeOaxIMBwU+wq
dCp3/e/tMjGmEnVFhX0c++blUVSF0kZD0mGvM5vVeoHLCo3MLA5ISebDUjGwFURd4WpmVr28hnRL
5WoI6s1U9l+3XPVMA1e7OZ3pYuW4E+NIzlX6+aYef46vUJ89NXli6kNe0zDmgblhCOf7DyePu0gv
1/TwuZ0P6OeZxV3mY9ZZEwcWlHoUlNACgVX7m/UUdQyclpItVHK/bPg+IeR/VaQCnBjfMWn0bY/b
PYEou0uvar52C6pWoQ3mRnB5X3zBOb6o161QxfISYfeG6P0yQu+sqlTjNFOAOcQGalDMQheWqJHL
DiApI5KJRvDEhUFJNTTcw0jZQHwUNKXLJArSf+5Vj1GMDjMKYW5L1zHGioM1uRVptO4CLnK7VzOp
S0kKFImw6yaxwWh8fO4zg8fr2fxCIhw2NtYYyYVJaGSttrNqTUerIvhE8x9LZErgiYcSLn41JCYJ
wH3Nuia0ipMLB44Pznbj3GD1bdZQjhfTeb+WQE6M3GstutUQGklgghKSu9IWwSa0+vrSguIwEwMY
DwVrGrsGV9MfLkIzLZEat4N9wPB1hrgEfvoZSqn6v6/RQErJkaRX8d7ONmVr6FQSL5s+33jwwWcO
YBXi2edl+NHH+D/cgDY0fuyXxBjn/aHMKjwbK1N4mmKhIi4gnKIaZRrIgWT+NJdO5lCAIrSFaSKi
gVZDtPuMEoQJI+FGs1L75RD6dXQ6ee7wJ7D5yg/DKAR5ij0KB3pSfPTFHHSe53TYPQO0CSDC9A8S
mIxv2OT1fDYEjkbzzJNJjMg7csmStwLTvlo4DHe57mASwTKGXnHiuG4NKq2OyugCItHS4kWPoGN2
4nSFfGuxTDry+viBuw3g8XYgkFLMbhdghlyq6yGA9AijzrsGfCwDY9T4i8Wfw1iOk2b7+dq3ct5P
oDFRD6vPYn3d6AI0xSnMVCd4lmDilhwJduKIX9M5APs7lnRj0y2dsereWQJpoiFIdar4I/xW223i
DVlW0BmaDLdRbZ8UglfzZTVEWmNZp1cb+1okVsvF5B+35oI7D0ufQeiuv6UJEqkzdiFmJQNs4vrn
w8lDyph/Bv9IhUInnyRkyGAqDC9BZ0OBssBFte/+OwheWT4rOoFKGQFpEX3oAxH7YCUZaroSF5I9
RB/hlgkcdSEnBHtw2mdH/VCwdc6jIJ1akaSV9m6ja9YA/A0WQ3rf2NYB6P5gx3EGhrXW0b3pgRQw
uazLsxhPhyA+m0BzBJSj4+ZX6TjcvbCXNKOxJ47yPnI9LInx0gsKGQJ36iZLc6KFilg/SIAmS3M4
hX/rEhgeFTCglO0NH9ZyBdQO77kEZ2ZAwH6gF2rqcYUTevM0yZKpF3pOu+oxRH7cDttfm5Ehrjem
UPdKYGUe51lEWTaILJM6c95YMogwDHcJHzjDb3QNhFhQVV2jkedXdHYJSEwne4ruZAZedl1weY5M
w8oNr8BZ7G/G/OMdw7GGHKZ1EL7UKw9i9ZfkOw5sYAQz+YKjcaMHuVQsEYgXejs/FcPyuDHgnqr6
CGitlKyFVGGvHfXwZVx6U/k6ZF/hkMuZfWCoVKEXvCRbEt9EwRe4UuHkm3rwxUE0FmHCjZNo/Pt/
8ip/s1nZea73dvYOE9ioVh+k/VPx5vMCuvRcAPxqFijRXkDoN8FJmD99isas1dojrBFxlC7dpxVI
neNhay1emZKyMQILVC1zlFH0yZ6oL5/0Y0zNocEjiKOGDXavM5qs7yO5M2YqiuVZPRGgybnoKSUd
N85En57HeUza4ER+stQ0qj72pzpWbf/UTIwj5pxaLnj3WoRjZoL6b6gk5XMt5OHirkvUC8IlmGW4
dqiInGQbIjLhZdA2rug2dEblG52Ddb7NWr/fKu5wavj0Jdj10p+f7FnVJQkdB2Gx4GSLJlDA9QEC
+ohq149IU/EYQxLR9J2i2O9kgwRyNjUnWRkM8/+Cn8jZV3GSjGfAiPHQ2vfHWPItveN6y/Eakk3i
F1UIspOP6L1LDniDBzndQwDFb1lukDVQM4I3B7vI89ehLATbDAXk4Og3CopKy4S98BmuLWFQbvQi
qNXFZNHddbH059s8vPnVqpBwpIIfRdDb/pV0zhx4nEIXl2Z/+DYySgoUeuzV5YWD0/Z90RImyyXf
7njsCxaqlezczByYqbxvcs9+DDyqq9QjafT1gvoSn4BSPIVWcxZvdsyoSOMqJ7vLuilho902HWVT
8OSPZJJDv1jX6SL29CfSJySHYDbWx+LaNxNoqho6v9pcOfLMZCDxsewOIb2PfdMEjd2SZwYwIAAk
fUWlTflw3h2KYiYVJO01PPLn+Ub5/U8a2pBbANQKw0AtJ5gdXcz++QI3jaYThmUYEWswfI1T+HPs
9GwS52/wjq7lmsl5JoJ4l2ILsdTDA99OAvi1yILsBbglY6nUmE7kVP4HvG781cxlRX9yciDLIJRN
H/d8CgdAV+Iv6zYM/zGpnZYusAdOOciy05nBS0AcWSasqrNTCPoVVba08Vb5loVT67XuN4rnhr86
FnUYgkSJHF4p/X9UGHOwk571xh/EA5jWSJ7jPfoLyAD9uBzmgYhbVEbJrwwNCKUOB0adP+GZGyG5
Y28g2fONWPlJqUxKMeIN/oy+LjlAhVZMPmnYEuzyOXEBk1+5SPB/gnH9lC5pilh39XE/8lpWtUfD
oZkSHURiOM2uPrgvvE3+XOjP6wIX2/iz1dkll3zyddQYFnLiyGqcz8Cl2yJVZwC1ssP3G2RZfwYA
vQDalnCr43hEcdsJuGbOKuiUQUJCOff+pMi3DWmuzSTZ01mieQXfoILa3V8X4sDm+1dK/NYS7QHN
O9yUxucVTrrxf6bkV38UrzWJ+2m4HYNccCiwT9Fgm3aCR1ehtt4P63RMN1CI/Q3BMcP+NGUM2VMz
4lm9oJhm6mZFHBlYQmuNiO6b1ck85EWYAcHh3qUAvBFoR7Jr2PoOs4dK+t+91CzfZrQYI9yUhEj1
3V1h1k/ZlS7xDPekZAgjx/V1SkX4KkLhdRu3E55lU5IAiVATx4/+Gv372iHVjZ1j8CM55H8rTitm
4bKI9bsB/a7c+XBc8kapgk98IE+ky8tzgySpiMzU3MakEI6qkLYrhYyXV2XNmvHGV79LEnDDunTg
fROKbj1t6WIm2iXg1k4kEzdXP+OZ1Yf7ANYegOb49hepSd2uSxfaqCRpT0IG2HnP6CBCBtqs5981
f5zmJWBzMsPDnzo0XacXgiDpZD0YLxkvWF2ErYfCrPMhPex6rs2HVvrpPHgzOPb/4URAWYNgFlIX
ATWM5FdgPvukZmpzGacG3rcRddmDvvt0gb3JxjKCW5rdGIVVIlps6QNg0O8p6JbEETfxiZgIg7w+
/dbug3C5FjAXqlS/1HUFtTReZWFFx5bWj3OhW22ybzywFs9h2oV6IRNrpWe4pjtM3pVJ2pB6W1H0
1qBeXb9CJPfBYvg+KWrJH0TEYr5KmISDX2BA+yISqqbr5UbmWCh5tSV1kx7W/keC9wc3niaReqIt
1/6ClBsU8LAPHLGFIossuqNYJLfc0SKARL5rl5bSNGuwf8YtEGjNv3rl7vAjQvoXp9J34J3HET2U
fZedBSR7upcQAqZrIRYO65S6I2NwvEibqbd9owVY5VhFDO8s0N0VHFpLaajQ9HJ0cmIEYGF3p7GO
OXUWLBbIpfSD9pjRkHzYMRJfvKF183bz/hg931l+URfvV8L2DL7aeXnBnOrnxo8EAqMJISyPX8My
DoOrIz4qCOxfSHVa4fRJDM1xMK6hAUUX84ZhX0+aB7R5nMOwf0m5yKPUrUsMXOnCeXrYjARQMX5m
qWsA/soFwDPnvctsuK4H4i5KL5EoMbWEdn+ATuSCLg4z+wZTCLo/XZsahnsZFnKFZXTU1LcDYbP/
J9jXp0L+KwpGJOHHW51mmDyPzic5lyuL8GYL/Hr2v9ivmGhBrUCdSplqtUU/iLV8jtIToLNvnWk9
I2lUhxPQ/+BRS2OLnlgEtuwqLObD9exKwKQbGPNNKAYxyL4jwiWOxerKZy5cDWvPeqYC+UdxHNX8
BoBuwUwR3U4/yuaplDzhEmR2SmaU+YqpaVAH5Gp9kKGdGa43b85zxRiMxx8YikvHWIwV6fTq6emg
zvC8GMfuUucGGQeD+Twj4hOnUNv+CS/cK5LWj/C+qic7IwdSvoBkBU00QQDUrs1wAPH2FKyhFY5t
7UDRRRxqQ84nZYyr6oOlMdxI1hNg+pusF+NkrUUJYCKuweqW92ecGkW0qsJ2MyTx2XNlfa2UgdzC
F6ovnE6cRcb4n4YuYBeiwfBs1+H6ihO0ZwTa5STmjWSfjg3ttvSayeBDLdFod3rKXJJKYw6B5QkB
FKG5EY1RAK+dGG2Qp2xTMh6K11TMx66KTmSr+1f/DyXc8IOgn9+NetFouhfiEtBQbfJ9DB7O8Rk6
hlzSwGTHyB1v0e/BFF2NZz+zXssvxBhDcWqND2yd469aifPbQi69KLM4vfcxlz3l8tQFYIh772A3
/cMMkwvqN+K543S6WwKTL9M/Nf4sRT8TGAchiNRcTIQD/PcUDWp1H7p5wKCXIZZ8T842dql2fPTl
T9mXI2gYIxH2YiGmCRh/DRDoNdi+/sftS7uGJXl62xbiYvkvXWoUTriaBxwn/gxZ1N0kBuJaSLl9
dGrfrXYxamMb2e3rLQSNGaNtzXiHQm9T2VtJKBmoU7k8y0ocDM6jxYjpqshYSy/2h8Ne3YSKxsQY
PR5WrYN6lhECzslmnUIGvlJszPddZd5AR3OtzGyTol2cWxIfEB2wKsU58rYUqTy0X4bOnyLi+PlJ
2yRiLRD3vFX2+Uf5kQBOQ8s3cfxCErTCq5RiWIjQjmnXyscL1u9+XuX+sioGHyg7h7VyCNT6nHSa
x/w+Xc8m+AWKKTU4p+PE6QKJytav+MtKrgknP0NTQorXooeE9qtAKrD+pob9pt3b+oNNEClTCYzc
SbEqtXSNd671EkJlGhZcrE4bVpEJFDg4NwQbMqIFF+XuMHg6u8mxXS+W5nrYgr2piGkZAERDQH08
EB2Kg0s2nEV9JVm5S58PepCTReJjvZKhkK2ltk00h2c/uOTbcYBgiSG0aHQEKxGpbm3LWUVk7WRU
UmrobxDz7KqJiBEVJt1Q1za5pmYyr+tpWMxUKZ5v2xtlyuOLPiMThogzZhM0dkB1pzbPx/GH5W62
j1hq46mqvLel/55DCF6TEtfI19IR6WJseUxjy3zHt/3f2Z6rogmJw/p2V+/yNqXlSBv3HWz+ijX5
zHtWCmnz7/FJW+Jz/BXfwJ3xHWHB5mngK/XyMH7D6zwnCtD67O+a3Mey20LpTNyGed6bojiFe5wZ
4qtniuHSrG504DAef812WQmXJKpyRBfJI1NENcehwVRajHL3YxP9568gOl4wjp/JyoH280AT2D6W
nbepKf8hFrxV3lBSHUdwH5efwVJ+zvLO4DfjQzmg2vQSapzHntKTE71W94V/hqcfLmP9/g1qGHrg
SdKr8w9HeYXcAFYPu5gxFdNrpuwaB/d6LgQWR4DMeQS5kTXWrSswAQtyRTY8ui/I/Xcrcr/g+zqs
372G2lRVfzZ5Q4H6UovZf+IiiqFvMKKMyktaoAOXFgOc1XUx95WanUvWLNEAMdbD0bfKKCOLX0xl
IhkmQBvVH3UQuQIf1cahQ0AFG2KpVWj92q24Yw4pZlvcplWuJUy9zOr3A1q0y84sLtykZLyul89N
5y39rbmsWSya3q9rhq7Fhqi6EtLe8lNhwoz7QuyCiXwra2Wrl3YavNtCNfD6E5iehmB8mGCiTzVr
keusOxcE2Du4LGkNOiMMYAWkh2CvGmz1m5qifnVJ5AQ804iZFZu1hvaQsPbyLQm6R+9sxw/ItLRE
R3ux5Ija23nhtHfWEoxIzEdev2dHCox5vAlo8Fm/Gx5N8D8YcvdZcaLftSDyqzg/ov9JZOsfEBKz
O7+uelLA2VgTf0Uv3qz5YiLr5b9vnTbeEKDUQuwcTK6zrjybPFS4qJhc/S9i1iayLbgsxccEbp2q
eLzU2ASsztkDabjP5yZPupZzIgkkwyUL/KZrW4nVoW+I3No3F9Neew96Ui52psM+xVP2fLQQHH8l
hCQsu11pEVyF60rlVEKyqiOnaUcoibGyd1TcVZZ2HThubiW+tlIpx62rnZpOQEIyrYCsQDqPme2x
iezf8al9mlMs2dSqk98w7EWiMEi1Ndo2WjwuW4KZpi0ES2aNVDlfCY/AoDkfLrIpsAmNsO8P5YBG
+bmjBcJQBHq65+JXyI2MQYpGfG/4IL9OAVMu6qfAY/fF5esmKEyJBZjCeaUKUDgpNHMG3by1TgpD
X0G+qGAVCpEmpgZPL5gmYyJVx5T62PQbufUWxX6kwh+0yt9AKYTHmfoYeVCz6+J11x6F3fZYiA4Q
Nmui/hQ1zf0E323OEDVo0e6QET+3cvI6xaAt+5SQ6tPK817G7AXo+Gck3RIzCKe7+te7kRLouRU0
o1S3AsCJDtAUZnXOnPrSB5E4LiTM+2dYcn14c0xdtGWH08tKqd0xS65mpPHCBo6BvBNNwyMH6IVk
g6Xz6OaxVXP6gZt2SwhqI0pMVHY9nrbUFgwudO2XlBfVVls1RZQyHG8rTgEY0ZORBDrNTHCqaohO
LD0RWSbycmk5McCEeD6lj7Rtz01DPlFjrOC9/rlQDTYLO6YMikXRm7LQhWnE6ExSw8sSA/wroOmM
WK2MVwPhFZbpzyyl2Crek+dW0cjeyaTVl5tYjx9JbDX7Tmi/4YFdLDFRT4aw5hB4GCStRQgYxg2f
aosoE4qb2g84p1eWbsbuH0uL8KHzl21ugs96VvNPceGoS85em3hXG5Dol+n/wfScBAZh8qKfgaqJ
/Cmk8kCcPiHBVihRuvxTLrTPncrHDH5T8EZbD/mi3o6K/hLbPWCANPs9f6jBlvW30/dtJlhqKOHC
xpQ/o186rR2GZZZbujZMTB24e/69ohvVSUMISOZuv6Xj8rSELyfsgfyOBQ/osfTXfnfug3/9zyp4
eapm6Svp5wa/TiA/2/qtKrwbg3NTJd5mIWYFU1oB13rV/2eBTnZ6tcLp3zRV0F6qX4rR+OvyGXRO
SRWCxGjLDyFb2noF5vhKZmDXu3bHNFuyfzhOIxqgaeSglBZcMv4nduEv467saQR6cEznM0dLNRhc
00FL+Yvn/f2wrEU9mMQR57nIu7YkMQkdm2yTJE9Osrq6vRyk/m2UDSlzvrTkBUiERwJp2U6XdjjH
kId7C2mE4uP5/jnNhEhvNQeCEdQoQ8yHZ8ouhVrCG+Vs9ZjQ863++WgMeRYFQgSW8qOkc4H6/Aef
gV4hgT9fk+DvHrtro82sHdsn1aiFr8dhlLyQAZuiKYOsmlEtOFmlfIeJdOzSMKKF7O18OcisFkEb
qVZ1gV6UALLsy70XnoW+dXXJNRhclizLf+d9SOiqIUiJprdoU2hqUkkwLKMt/71zN86u3JGNjlrs
DtwQPpQGLKkn4C6YtlsRTPqBtD9KRXNdvugQtSL1sqo+Xq4ADRMGdV9omVq0+L1dYKaKp2cB+48R
6vO6YmlBmUUNT+ImO6H78fccxmiTVgihvQ5kTXu4uOZRS7kiqtUZ24e+j8l03YMatgQ7YyNp9NWD
0eB/Xj7lIFob1fMW60ATksR+Ub5LcjAVP6y4YiaNzcPgNfFtvEbrvf7Z8BRt41T1UN1Jwnikhf6X
U6JwxwnuuDbW5SHJoEnyAvsjGFPW4TZAob0h0CnpLN5YeWupjrxRrc7oq7fh9yyAS0xt/WdlBacx
q7FnXPAOalQxFpQt/cvYtDHYZ2SE0NRUk6rZEMdiURhKwmRi4XbY15yv9uAWDWlLKX2N8d1ZhNqW
o/vbDM2qwMmgGIhcQ6OAqlBGp/8DBGdE48kINjs0p4mkOHty7Iw7mi7Jf8GV3j5AqCwKCj5q7EB+
MFUrFneWR3a92bif3NMWS+kqN3MAqqijiSJRhPjm0455aBF2hUcRZfx13TsZn4IpKa82K8Zi7yvz
f1nCKub9FH5yd+KihDVMfo+CGy4SLEHoTHHw1a8oEROc/X/bhg+UPkpmLR1mZqPLgdI21eZuQszH
Dh/qhxiiwW1WhcUU8vl3NRPoG7NO/aEWfRn1sR5lCMGzrW39OJJdLVRtWVpWrEzf9659m7+bG2Mc
wEK5m5NFSQpgP/dgXsPhu07nQ9wZcYosSpYHTZK1d1Q0TjlsdYIThUMo1+aj+0F1+nUdcipGBfjO
dpTOMhgJ0n8eqoyyQaf1mIxJcrI/fJd1PFfYfxw0UngZ1UGeulByjyOV7NcAUN+6iN9R0ATkH/CM
MdLdzYUykVErYXWrZgX832IceIVME8SKZ0IZggD/8dx3carg6AhTSNA8HGSUWE4E5L35hJO6FZ/J
pSYf10s3bzvogrBqY9DnVPzjgrLHw7WJ9Tt3k5JP5XLT+hrhywLfi1aGwnayuDvHKFQvYcGbXq3X
sBZvZsLtV3STxJiCmpg5u2j0ahL7Uhox/4Ew6oqIMELPso+1oNi0JgOuVbo8quXKeh0KHegb0Hc7
+kvVR8vesAnnKlgnPuE7AFbG8rQG8EZEGCvwVVdNLl8oUPa+vvBgeGuH7Of93/FIPNG1uEWvOtr0
4lb8XIiT9Dmr+kSatlLTw+dlsuAmXaWNnip1Qks1jgSFgg2lK3E7xCXI2DHTYwAiRTVBAenSxMI+
67CcxpgfYzwrijF9gBiHsovS3YnLtY5vCnfdeE2F2I3QcqkOzCnAeQE7SK3UgLcyJMuOXCkt6K6O
Yz2VTpSDCE10vE9ViGwHBV9RN8ybxv7jKzms4F3Q4Arqe1XYmmavY7G7RihlLTFMtL2Yfx6pxfD4
j9p3ZyLxdqPHxq9gUl4G6y8v4nJAUW8S2qa66TjOZSWTqAPMCE3o8XLQzC/kLS2NRrHKHQ31icd2
qKPvZsx/b6fS8/mhLf+i1sT93bgr7afFXUcfroZtuA22m9yJFfA+AmdNiMKZhLDYkGtT6ZFj9mOf
GJUIN3/ajN9/+BI7Ts7tXzhOkM1qyAsOYMwz9VrFJmUIaqcU/G1mx9Z1k0vi8Yx9RyHbBefaHrE7
KqRRigFHbOzoRg6+6bPUyNRNA4v5gjGpeR74+/ZtYA8MfSZBtrCEkWFhmCy5Zgs23jVjpE3GHgud
lN+0s/t2mXMcaS5pJb4+f1BGAIHhKFkB59DCaDwsGlv9OY4CA8rgB7yDl3ERzmLY1j7p9T2iML00
xw9kT1m2FMKkgcRNkNs2GOBBtpq3ywxyBP/Jdc7hBO15FUsqpWqS/IiKiqTvc1R3gxerMLlcIAgH
MmlBUvfNFaq7agbDbKdqLm4UgEmOjoxAh+f63dZlLXeEpkJDVPoRL4LwCsIU2/ue/NlponP31EbH
wIveC/D4HQWHJ6PQQJX1bN/Q2HfC/FOGjPus+YwjkJgtCdOoGjxORJXu4O9eVWIo25uiykZY7tOb
hNeqybk4rAj8KhAxOQUkcDlFyf8Sl4nT+cdp1BNzibpQXDFdMea3R7o3y5uhDqwX7EGjYz89SDbm
ORmOo6Mpvs9ojmi5uqrSXL48H5CnhzGFuAbmYBUT+fHAsR7AM7fskjlb0Wm+eVIuaZwVag2BPTMb
W9slObd+SO6QJlLIbxRNiPJSNYr/daTVAoJ5ihRYesJ6p2+o/iqPrsAO9FYXh54XgbfQBpuqkpVe
B7EwpidBkeb1HLDiG3JJq9QRi2akgUjJ6J5AfHKc8SwG4P/d1PDlmhoIGt43gx4cIqzi89F7YLjp
hpjJJc2+5LbuCNsH/nGv+g9Vxus66lDe02FMIuD666O0GAJzJmdR08/QdKLC+y27k1W1UqLNS43i
ip2FF613AcbzMDB3TiE+bEBIMEvQ7uuoknfuIVAI3BZXWiE5Iw0MY8hjxAYGJaFvnpwNJvrGQXIO
EwVyFBVyhW8Q6qU59rvBC08SCG2EGNJHgXkVkziMz7qGiKrioxxkeAi/aFkFilnvN3/qAPRiwO9+
x9xYPmUgZH2UiSRri0YdNRclv6ze1n/vUAJYTJGeReaUkhTuSSsN8J3YStM78RS6u+AyNk49Rk78
qDcHrbgg9jwyIQEbwRVOnItnZ5Z20VX4qv8lpBRiPsB3Q+yQrJ7hKLXIU7t++PmFGtZqSl0M8g6G
vH8x5+r0uYBA42yyG/zmihkLv6VggaYhHuEsBJYKUmBf566g0x0bYJqPyX/i+coa+muxQJ3dsdEC
yGSdeCvBqDKbSfSNMS8ccdj6fzV2iyysadB9kpXYFIPVApwLgjC6rEiloGXEKm9yMru/zZ2L6AjZ
e0GdeUfqiQliNk5xHwKznlL1mR99BtPUrW1/S+vtKjKonRERIYgQ99tqaGXKMrDBQCx/5H5nMI1c
QN4oK07aQegeFOBA8us+lS8eFhFHPdvhNEAE2kD6Qp8yWO1dbzGqDfAVIp1LULb7sb7mmb81pPqX
Gk6BpoCrU8jx9SSCfCrMbU4i17BBOKDR+tOzgo2RgUHtp992UeOAalgoYGkG5jF0sClR1vaMWs7G
H2sLflLCXo1HtNJfwhFVr5PXscoLqjlAEXZgA89PH1hjEvMdx4EwGQgXQr6Lp3Zc8iH/pcEBbhTy
iTvbtv5eb6Gfv+84/QwzY4mijGaI//961fDOti+YssN+KDApMZj36HsiLvOc4xNoosNQzb0zp4QF
HcmlQKO6/JlBYZjI29/HRJL/woDLsc/8RXK0hI3XDEaAv6T97m2xqVp8+FnpIt/BROcHI88Uc+/O
i/mqBLhhc5/QB+tA/doVc881a67HZLgUPlEaWfCFrnrZrf+ulHO97I2LuqP7Of/WUaLlg20geRbG
adnI4ObTiidjfaBsH003RSrPOTE+HIPQ3gLK4mg4d86wf9tK4idQ4YaMnEAIMhZh4hJiSIwZIsOo
zacD+gueo/BJKkKvChKopD+m6XM8Bo0/sQ+LAWFWXKDj4nR1pWwGtFn+HLoL6/q8BC+Aycxo2y27
nDb0CXd/3WtBAXVBjr3iKU70PhplI5gBhikrzUVNgaHjZejtmBGgTnBB86Rp47u6F8M+O/RBDmWP
7USzO6shEPZeJyDoHs6IxGJE+JKTtGN3IAcBUjU/ZxG5is0x3Z1OvygC98RbhV9jZiUovUcaTzl9
R6O7kLc0Dm+IpQwQ57xVzMb8yizK6txqbcwgNz+uNC80R5g1XLZbyXlHH727JiNLtQzFWEY5Hwn0
EM2XMoKS48Y3Xi8Rim8NVo7uSAUq+/DQidN8e9Lwrymtj7LzcQwp0bPK6mnxjQ5CYYup5rT4SYWM
JaXT+Ap1FdygglI5+VDEobUN5Edw8SxfyuJ92E0ioLuVWvWtIM0QrgewzXFfCzuv9O2ygvVHNRUc
SZbighFrkD6JhWgvGi9iu5zY8Xc+ZSVzWxjiLtDpbP92IDuk7OsiRDUsUJL2KntpLOisuIRYRXnO
I/ajDJJhYa0xH1jFO6EkGCSgVp4O+Y09OjV+krThfeQgdyBPKz4aotQ34VFuOeakvzHBYMOI+kbu
Zy2cCbW+oM2ymfdvSYWRz1surQbdF0A74olj+3Lab9ptlyRfHCeliptwwhbJiVXpHx9JizO+r8Ty
cSl73xSWWwdqEpLHoyVkoNNsJy4a4iauEQwVMqRmgWZ+9KIca3BhB/Kd7BvOiG5MTkFFkg3Mum64
RfLpDsLV6+qTLj3Ib/2kib4DQrq03Iya8Nta21+jAB0QWj75/y3BKFdHlbg5J2Kq2nOlndzujzQY
J8jP7x7qp/EqJQ+6JP05Pw1ldSktL7VenWbYsrbcmUZAm/XaTyQDMNosc4PwkoTEpxKegGB0pRv6
QGmCBZ3awy7PgI1lxn3bEptJbpq4owqdSMBe+nompsB6omHemeRARlr/FDzB2UjywhcYbW/c1mBl
abEVCmcqDy7fW+vdh+nbhjKJiPzgRDE+CcM1Z1FqZmROR6zqSblOPWPWMFu3M5rgsf99AvQJ91cf
0y1+Ia0d9zx3E6g843OoOa/tpCUbwoYAajP3Q5QK5p/1dEKYhmjQrRkrHmez/v9enHwVv6uc294R
xmmYKNWsnMJOgh3OqvaB6h13Ne4q0IxScVj4Kjy5LLvhrzxY7qlyiN7XBbM/8kk1sDkuwMJAZMRh
yQ60PhqR/KnV3sBqNXQkuPuSh6YaWqlzdiMx6+eQreouWkAsivjL3EqnpoACl0yxkA7X4V92Mpv5
M+Us29JKFTET2ptog7Qhe8QWLXarAfAOSp7V0amCU6j+OFthT2B2CUdaVzWv3jM33tAgmPDdm5tH
MuA18oKjtTUctuN8KyTVSDfXHS137J/ZNrstYpV6TYhKOXugGLa6Cg52GTReegW58wIJMtxHdyqS
z8U/4+F8je2KL17pk0H7w6Xw+82jAZM4Sz6SqZ9zyzwXx59KM1Cunfcu3nzVZ12TphNP+1M8hqPY
0zCkg/tPMJl09/BIGFYIA6wPfwMOC/Z/EuXLHSc3dIohqWPJre4TytVHkuNQDEBAvAwoektmU1Av
78Y5sx5h32CGbmhKJ05ZNIQt0vS8sDqSkO9xFiSb9osnMmE72IzBIP4ITidr+fkT1UG+eMXMrUz7
whpP0C2XoSqCpckSg5c1RHe7pqc2gnhmCRf7XLiwiAdfWVaA9phCCB06VX/nwf3I6BsiOLUB2G6i
UCDaM5T2OZB0IRJ3KTVu4VCKGl74Oc+yrslrxI68yI10Dp2nKCRajT/7uSGGK/4w4N9TusWroNPS
ZKGqM6T3e8rMc9MZ3oVJ+YWHwzn16EeKdPiMxVcrCbKXCw8QYLKMgq0WOH/qt//nDKbiHPm+0mYK
haarkbezHc11x/Uw1VuKgpJyys0pHxxRBnwZ2YNkGQVAhP4l4N/b61tLjY8zLgdvTMexZO7ztJ+Q
REvWYQxo6AdN4tcDolpB91uYrqNzapey3RyrD1zPzd57H8WlDZhntVbFMfwEJt0GU4j3PeZfhREp
Kx7j3sMZXUfFn6O7f11jmRGtFZhAHXCC4BoRHHV3DsmN69O5u+x+eCJBRAbqDRPoDy9Oira1938O
HdBHsI0Nxd9TAmkBFQDlkFpASgeizMX+VWRtaJ3S4dl1/XtfvCcf6A7/CzUBjZwxW3kdDkLP06U3
/XVDzPoVWZ+gtWFf3UHxRg7/dm4wSHs2LXcrP1kFkkYoG9BV17K3uhSKxMQj//WWQv3VqTqcS1Or
zqMeRvp0SZnJiqFc85ZDhuYUF9TMCRKCyi4SKlA2kzdQJZuAVPmr6q1SkCvZjywXqAiwwDtgpSbk
xcPxqXZ8orrHuxtA/NvwBjsEwNtcbcGwKIBc75s77NWjRjDK3Y+SCNeYvKuOcmYqStyuzPcQDAHK
bbXfqoMqX+COldD7yNrAFFzL5dqv4nJG33zujOZ58oGeu+3h130ZTtfj9BrnNMlN0VSW+adLrewA
Fr5Sdfhk3G/+oEGKJ8A71OXQEOwGADcJAQD9QWUecurfNTacULn9WXhKgeGq/i6comSPYuLEFu+v
U60kV99PEUoPjBzIclSUMITQXUYtqxm53Cb0IDJnHSBQiyWJYwVBMFVDNEpQElfXfjCy6RL417KN
ecKBy2JQcAgWfb4xSACYF9eMY6lpB66JXXEQq/hkn2MdqkA/h9FYHh1xCWHPu7zyXwoWL0xRuHpw
qPASM1cpNBTk43gVKe5tfXnO12uON1NQox5m57TEzE27yD+h8L6bCXBrtXnLFVDYZSXsi6H6do5z
yV/R7eiFIxMTHhWZ6xSNyLf9Cr2h4VhZVitvfYpweDEllI/CcBwYtoDO25sB03nk2TpEkMusKpy/
hto/7lTKbSnEmJ7cBhpBQnseVf1va9e/JqLT16eB1aRXInSBBCdgEhYmZWA71M8pO97nawlj+tHY
5T/msIc3Ov9cdHqR7hOz/HvehQ5hTZcwLT8LVL+YtrCJa688lt+uKcmGe71jfpfj3vd1Af7bZAHI
i6dwqhqmruGI/lyuoXtEuck3PyWjhbBtwUQ4gTv/H6y+bQKdi6g6H7cZNtrGcMKMLHfpg6EHwGzx
4s7oChX4cj8ppArxSmmxB7VndrqWPYoduvCDOe6FPoumpl+Ru/NhQIQo74u80pznfnTqMyx64t3u
FPHyrgioJMgre/mLPEalomkHvkb7B31dYSaujd4XWcLpRnapkWaKx3lExBiht3kjx8O6Y+mmoaFx
5D5XZ1UFhCRrtrGgOZvfmO0jEXcOrowsz/3j92lJ1D3J2/+IpoBQXJ8QwtN2LZOZIY6DoH0rHjSJ
RPZC6aqzTxLju3oTFfchFnR95d4VtoWXb5fVoGQF/yomQpyU2ZzD6ugL3wCjCddcitWlK4j3+0+t
8v/CgRmfTapKLKBxnvqJjp+dWFiXbG2YcPT0WcvC9Ts/cB0rEb5XWWPayhgLONQIdY7WIf+RcjP8
bLz+8k50lMzVYLg+it4/4cPiguFloftslldi6iTZ73dEaAkbRa3ZkYkFsECeDbJo8yBz9O081YRM
I403z+TezL9y+qSlhdFaWB0xIw8DFg+f8q6/aKSyT+r2R1WW9JiceBUGfwU3K6nWUS5DCdfhbyDj
OIVQjXudFbrOGO301QYjC+nQmmg8TtcwCKWmce0BQU5ioEP76lAz9ole5qUdEX4zzxqd4R6QQNfU
jDyumSKyaMa7mTE380rQ//WIKXEx7fJ60f9V6Qyna4814sepFst2Zo9rnqEFKuW7Xr6IPj0dsC27
NJ1kmLdPK1vHv71SZTWKUM9lj99yB1KcYR6WbZAOAqC1XrAh6lhpykIo46wdMCFWDeuOSx5MdFBH
wXviNzu5LmNMEsUU5gwrscY9lLZgGVbQTlHdmNcPaBq2UDv2lzp8Nm0i5FgxEo1RNtY5u0LOMhWW
Dhg7xbJQn2GxWyHobZxa+vWJYxzM4yOokgPBnfxjIG8k3s0rYXgLKJrQk0gJeIMFIpHK5+iDS8v3
Rr2s2N1x0EIYhCW0afJL/6341grMIJGH8GtcZ9L4BpTUSopnH8qFS6gnwoGPTofwv715RmiiwdC2
RDDj6CfecADwojv4CV07iEMPx34hLTdxgLrJKJTLTa6GlEmAkNqTzl1D0sO+7Qmuoo1f761/011B
61kLsZ2KF3IKlzB63tepSbkJ1Q4k8P6WHm3p6qv4XA1ehcQ3GKjNmFxwzbcNAe3dfiDwIXmCIVj3
c9aLlHy76bbWzRJ0mc2sRylcfygTjIQdUAvgD8/ViA1jwEL8pQvP/Xv1Wi+3FeiE1UNph2oV69Dk
oODETSr5F38ZdHOWVQVE/+scLE5vHv3fJSM9yBPIQxOAwiBe871Y2lvp1pYoGshBBvySG2oqVj4K
rN+SVOl5R7YiiDH6hraC2XfK+zijj6y9FJMejC10Kd0Hr5C4g8oQc2Rx2gK5scoD/242JMnWkjJc
JFJ+pRd8z1BOKX8d6UihKCbjR/m5Dpe3PBZsDrsdnvN2f4W+vjPwbKZnEqo6zeGGvCVZD7La7D4H
l/DkRm30dfSIYq6s2RPKMptTpSdoJmi1N45jo3mdATHIG3vyo3rV12UO5qAWdbmqInicqaqI2fKV
72K52LF7roDiHBjFU4Mmiaj+nIqzW4UwGvY7LIn+vlw2LjmPq9obEFi2OSb5hdqFc1wdpjfXiTOT
hVFU25Vq7CT9Bri3yQWvxVlNCscneQHaN3Hao4SU7MJUTKP2Dq2iPJZteUokiQbwpP6gbYlgpiRt
tZJ7hW22ZVy7CM8oQMkGTDdth6UavNqXf6PW/Go7KlKNHoY4NBMSVb4MAVQRGe86Z6LSXUVmzCCG
o7qaWPCw6etjy+FHxeRosT84InwgxCZy8FCm0p7O+xsdffHzdZBLyaSbiKa9M12PN1q8vG14FhKA
I5hPtQoQ2f9hIhpqCaBuTRYJAI59ecW8/vJxOg31Fe9MP+jaqpfhcuLXiwX9EfvbLa6jc4kJXxs5
OPkfV5bJjDwI2AG3mWpCtrFZR7JuchXc4ln5F2LNjTOf0BYW5YWUm4ZSGDJwWaLZkj/ku+EVTOgz
bPVyFI6w62z/hJXucM6vrjrHvhRRpaufolBDeh1Rt8Ua7wAr9NkOdQmlQeXd6twYABHZfSHYwBSC
kTmFquLtToE0RgyFJP9nIAwkdpl9YJdzHS2ITOL/APbLZF9EaE3IMarxF4+YaoSrlQgOyFlN7mpX
IIu8g16xuUq+hiMkURrFQagp6fbn9/Tvd60wbLLOfzPbstvbqRz1Q7wtgEWWqXOzqOFM1ah1oOA2
LQvXoTs9vMsNpoXJmeohl+gZA8XRRS/AVLrxy04MdoaqbfLtwcbc+tJj2JXW4XbH4ZI53Hu2B4zL
ZJ09Hh62SBNPeogLKuyim168KPqATLmf1/jV6Gzz4lt44aCBEuwY64vJ4Vxlet+1HXTEWSXQAFpV
Lyl6z4ISYTlY+JSBznBIHtAvd17RbGfxbwCIRJSuwBmOh7Qkqkba/RXcttuj2olWQLb8C/m11QxF
tCR7xZzh+10FF6GKmF+FXDmsOq64SOf7O3suY4yeWX3CQjQBvKYA1qxCdl3hnLtHcZLJr95yZkMN
BDd0FRfUDlegOBKlxDPojJITsAigjn8AtxOQKop4cMIRos2Y5XSdGzqXGQ6VxfqkITn/Y7kjSipd
y3P7BnUc8eF5/N7pKRgjT85XV2JeMn07Yds12m7sNKUEA/Ds/SOh2kPSuEuTIwumv1m2oPQgvJ/j
qb9PVG84CQjspK9Ly+3mCuJP8/6ksOIAY8ZxxJKWFFMagbel9SLM+1eTEyOv8QZHNju+GLWaGbJY
CkGPu+ADLJVIamkCHyt2YYec3rSJTLT/pCg7ncXBvAka6MInA0dkFhEyz4ckjChDakzuRMrJro3K
+UtUi4V+BG3PwUERi1AX3lHkS41Oea9cbMK0CBQdQgyScvaACOAlnCFlmdn4/9fS79dmB1TbZERf
hBlg3CaDRUrVGzq1Q1KKSTPdO+D3kWt3USt+3blV1kODvaIm4MdpqruWLJkGQ1helkKvGhnLnElT
IZCtXOFyeAPnLtyn72vlCKZUqCZJ2+t/YcVqwE+pHfXHTbA4vR461kem2ByEcJDeU5lF59Uqiz54
J1kB5rfYHAd64zaylUfkskIzG8GeUTW9zWqN3umc+raGsou80d33WQ9b5RO5/mGL246OEgjaTEuL
cejrv5lQm9v//TLaeku56zHl6pWpyXF1dA82h6OZUnHzNFobOlNDcRMMXLFWfyYu8vC+x752Hblp
KuhFBkcIZNRBKCLMwXDfd8/ZHg3Tr72k8BsULy4zwQbzCaCLUUlnL8NsE7YYs3Irex7fNV7736se
fxgqMgazFpLziPSBgdBa1JoKC2IOrn+2UWYLbowQ2FEp3PkjX8EmA+NH8E/+4/vdYhgKKyBini7K
6V2V2z9h48IJEsWWss4uHjSViLJBpL4OSwP6Fl7UfcrQE7/SD4gpfHN7aLY9pFmAOFUM3NGrsk20
kE36QWlh5lwwzrtD+V/uK8joLjujZ2HaUQQZJSBrYe+mqb5CpcVWU8fIlq2t+ZVj0jLsSdiVpwRX
DcdGloCHERxsrLT3DX/Azi+vz1VEZstD/WsmSRBAhLrm0FSV242DqCWYrQDvtcZ/Tg2tjni/g73y
I6C82aA8eF8jb54D3jrHj/TDQr5DVgi77eTZBZTGpvMDFfJGaLQPKgffAPT5eaH/AJZR+RT5QBbk
NBYq1t5R3rkpujCmKCjLhKB++hDlbO5duF/dkj6mb611qAW54zdv3hM0HaS4ajcx8XCH35BPYN+z
JvWeb4pDJn/ErRYWyxS+XLc4S3PAY4BXYbZHCw1rRYLiLf7oSPs3g02d2mUldZpVRyTqavYcv98N
Mc67njiXQYuStZRQhl36YFPz/RMywGPz8g95/DJa2KWASLLTpqlaWaKo8W/8Qe921OwhmhP+3XIw
b+7wAGsG6DQd3ZPszM0nuBxTDmNE928ryJaMogQeuZyuAywU9u5WCDyLoM+j4qyRPRJj4gcfUQ+s
N601kskERXgjBaxSDGfKRGmq31nez12AEJ+xPsO6mn37IhsvAM8ORV2wuTtGl9exeVbB7NgDX8Kw
+ky4UipN8kKgskh37Ph7JwBRwu5OVAQqCknB5PTJ5H4Qa5AZZz9ZsYOd8keaEME2Pxlbc4R1AmPy
8/Q0MW6tP0kNSwTveFKjG3pZuqVwxcX9GnXIMs6bQwUo7BlySgqChlx9CxdhA2oMaZsYHsTuJhP4
ZX+KQ6AJnUPEYJvx5rl5ZAiyvZy0BfrK18urWgtr1M70nqthNfcCc2DzgavjIqB5Va0Jfc5x75yT
Orp2SeV0bLTJCwYeF3ELMTKXDWuR8/YicBd/DiIWixKtmPDj7qErzkBETwpua3vcsj9VkPpzIf7v
/eRXJncDXkT4BnZ7YViZ1t7GhbvsiJm0qg6zSftzLeWwr9eP0JeTJF4ioe0L+nNFOGzWHIqkaEUn
xT2bj/UX04lYDIb7W9TtpHjiOX3KsNMdLru1zZJ8LbkEEMiRLYdLg9HbASXXhsnech3PWVW/UtfH
OeSO4puuE59y1z/oRdrn6PfAglPwwPESxMyMPlVqMpmuD5cE/e7fqDDpl/uhgrdxzrNefClofYp0
u5/EKRZUqVRUYfdv6IQkH02bZfgDDZw/ETvHEQhcbkTqbPUbEXs19lWBjTC7S7GyreQypCxHbv7O
ivWz2SLAW+ufqtwg10Ms9E0y2fQmCbVg02bg4DyJ47qAg/bMDJqkbmiAuzH7ytoB7BrQG8uDy+nS
crJKK6nQeiyqccKyN8d2Dz4AzMLc6bHYt9NnbcQ+jT8CCDtTYPwrg5yuWdOEtlUM/H2J8TEEsaij
288GiwiIEDxXk6YaokqcB3leB22uzKD59wnB1eK1XQ6dZL00Y2GmBMfJmbSi3plsQVpSOgMZIiYn
YkXaKqB9CWbnL5rSUKCoO8HrBFDjLeGleZ2G+Hb4a6rIsc+avkNp5BR6fRgE/leywenWhXcXNx7G
FxLLIa47SvSFVWe5h6gn+WPqy6xO5P0egIV1uHd7wQGJAWpJdGTfEr+hgaqmxCtzJxXWHKBfKIUG
4+cARKxBAwTp4nPieEq4mYBKJhn9D1dBTMu+CTgzHKfTMEzAeKi++VxpNXHKn7PbUlli24jufH9W
2fzjemD8dGoLegslL1sVsO2/j6NrLQ941aQXd9M9xhz7fSLFxiBqqQ7I9Y+ufrjt6VzaavtTrmyF
kKwBA31/J3vEhD/onZO4k9EmGrEbqsIHiAKEeMQwn/91/5k9+CJS5eX+Js2AT/lJwWy/l/dD08Ty
BpMjzPTj2d2gEGhOg54sw0F20fDioxGb5BpJDJMTUO2XwC2vM/HF0GB5tarKFqi4r1wqoEVNj0pB
CSv+FJP29Vvz4/MTtF6bgU8lbgwu4LkKI86rKR5rdUyNNB9UyDKcysMpqP1v0tZB/R2FqHXIOPM/
yqZ9s1wE21T5gLUXbVvCnR7cIF37cGWYHxJ3+Uci6hSV/N4Loiw1xfCG7yAengTFK/1LXrjCFUe+
M2y5ZlPKtWagmGh4mku0QHn5LVLy3eAyViok/D3dlLgORwNMO5jYmLPBD8zPmLys0oZdKk/zS6Et
MLlB8fiyHrGCYxxN8WZoNLc8FdkxHFXPIfsLqjEbEeeDdEXJXnK1s0wk756AEB32MbjqzngqNBjc
lSS/2fLM9qmf0fm9h4tProy+S3yLsEqr78HZz/gNGXvJIb9ugqrn1Tsl93fisx3MZFZ5rzsbTKgy
ScGJiI68fHROECJm1Qp4xZwASVkLGVU2eCLn0o902vzzOQDG3cE0bQN/fbhjDYWFd4Q8R1t6P2bt
uto+Je42Zen+ptnupY/NvCsgNLrvJa4lNsomGw9OtzJ+jZQQEHplC430rIgYD6P08K/LJWnUGXnA
3SCofg2aTNEUP2IIfZtVKsIH32A5ZDOArjlMYJIQPzmR0qbvaLGdJr5K05tCyP73D3/0SCw6l2bh
MtncODibLe5MHYvf+IzyuB85Jkbz3kDY9vU47dvI4hi7zXoD9IMAgI+hx0MXoHhgOsah396w5I5c
8pcug4gEnLevYFadwb8ovdnYK7AaN8PVmSYrPUp2f/OUynP5cDZJRM5yuD9P5OZR0wemVIzWS8pr
XO89tORqMHe3uNmDNsxtKrciMDyKGyRZ3xcnbGRUqqOdTWZjwWluSpFAFgscsrVQXwBtCjFxmqav
tUn5BTNnGuZIUsC8Vn6zS0Vt+PS+aEZ7cRMDDSx2Mhl8if75OPesWv3MDAmX3sWY5b5e6qZ+tE46
kLq3cf2lrJhcPDOQAGBNjbWLpoaS8njHG/MJTUJ1UsfAJBsIjFXCwwsjb8DrVpLHkSgR2ZQu06In
Vjc6TeakiJvzX/D5gdrIF4gK+dqAZPn58Oy32BpjMY7yFfFG3x4PhZ3K0VVjk3VpVnUjH1YbWeZQ
vD0+wmtFb/dKx4ww/T59ogrS0Qnhhx7pOf41WjQj8MofXTG0Qawj1R/4g5vM95416O0w+UJYaQO0
lK7ARRpRxaKF+bTxCY6julEnp4oi8UHrGEk4AaElHxWvFaZBthx2NgMCRi8/sTorizT2o9q9BzJM
LhnYRRSVOfDCk1wF3PebaKbDsCsYI8AVjqjaNUZfpeREdaKRPtoEPpi3IGdwRH+6N6hGANWGMJCv
sqkx5Nz1tuqqmTnx0rZBcQex8ey0aVOrW7Ol/5qdK1BTMtBgcGBCa1L4+why6WZvD5+//ikgm86/
z/8plMboEMtWqCHiQMmhHLNz6HRjJiCucfShe4zQx+zlwSiG1GAaoNSwiYgL1Id5fqGH5tRmXU80
tyH9yUSolKuHjak+/UPAmz1JKtcv/pbZ4ZlkKBW58/GUiyJ+RkTXmBAGE9nj2SJhayyQbxQigNFo
re/iL31JXzIPc1YueOpVaPT+u6BHrJHeIvEAK85L/PD5NIBuYziM8zOZKG5yK4UgZ2rncDfJw6xz
a6HCgv4DdtyXnJMyvz4WfBMBLaDubzueMYat02jd0evNmiYvgmxjtVHFNtnmrigdIOyBGSmtKjfJ
vv81g5fYozk0ccnljhAnlHjjf6TEMCrKLab33gZgP2rx4S278xxJ7i/lELzi5KacaGlgynVEpaYo
DIPLZSMubxcGwpqLXkIpJNCJton53v8K8obKQOHZFGpfBJUruinC/Iqa1nqkEml9EQC8Kz/5WJCz
9VimsfknKwd1JWhsTw0brgtm5RYuXn6Lsi6r1Bx3MxF5ABzgNoUDLqv8IaTU4QGuuV3+bAJ/vkdn
1By6IELdyQflFiGNoPJ0Nunr2HwLmmoRz4PPwuxJqL4vEY1TqSIpGHEzIuNWKQDvSiZMWlPez4km
xPYhTUWjLVhXyY3bWZNEyVU0ReJ3H6+cXOAzRkx1HcT9LyJJslL0SotY1YF4Uz9Weqtvq8iJU4eK
GjpK56qBeMvANdZ423/trunSFH3TvyZ7qVqW1UnZL0Ge0O4uEorWa/o2y8fQkouvBDWIPgVOZ4Al
F/9mmAWFlbY15/nIt74KR4/tCxkxKTaDY2LUtxhJ1ySqf1Dcf1NOG6tEyxqZ068HfEB26b3MqyVU
IK31rgx0XPiwfTfW65byDH/EMQSB8IDFpApe0VwCUP3Mu9tKmY56T0J/OpjcBhgQ3m4qwRIuapIz
LSQ+3eF/+YWzCVWQoCe8dCPF/SQ+y/sbhNXQe56C/dtQKgWdq+rsvDvXtSU9UsrSa6vJKc4/y8tZ
mm/S2KEzrY6gXISfhDrrGhLFU7nIBFK9U/UmoZ18conaafj5cMhZ2TogFU/OqJU8gGfFhvnyMuTC
pw5At9M95Jjerd4IwqSaN5EAyQVZmYfctvJu7K9lxIQ3WzXm2YUgCjb18xgHEJ+8ftFdmD+4JtyH
r7YZfzHfGMH4zswu9LmbN7gLi6WEJoe9f/ZW3x+mHi2qFmE3XFwjtJMPNnoyngbgFGzkxuyQUK+1
bqTxAkddhJJ+tY9oO9sILLqmf86xTqtu1nMRCf6nluAT0ExJBmp4PkHbd6gsnzAEUcZoW6iHhaDz
SNqdaVCpylzuMJR66hUJY9Pli6zVyYuq8IrROiFuYfO/ORa8/LUsPW+Y1G+DDEAqt0+YK9iYvmXr
RPvWQTN3OmjU6u6qmrafCeK56lZo/15GwjsuMZj/97Mnuj7LVNRcGHZEBqwFyrNCS1VmHeN6bIu7
8PiYOXcgOG31TlTyh/c4YXPiIWr0+pACIgkNuw+MMKRUtwt76U7o7Jiuz4r6LoAR9dNREcUi+f2T
fOYruyI/gqYh9TCyASqwzzbUg+cfFPT7mVye3zN01wsf7roZ5TC9OTebhwJpMMC/2rEuWUqTMaMh
n/3ENVganlT+Go7tJQz1nhgbg+0aWPlVeWig5t4hrf28EEe9XjzM/NfFhW4yuzfKwN2d3+iuNnPI
LgRwZgOyGUYmgrhVLpz/6JvN8mO2JSWHUqjv0cSatPFOZiKUbS6WsCS40+HmtJigdWtdTBb69MIX
nWFuwO50ZqLPFIF97ONNyhik5i9VW0ygtrFlQz/ZKqzh6Aj1buWib8OOJgeDrlV7YhwRFDq2aNMe
6xASCQCf181/vqidPV6/HbKFW6TuuGcirrMazPTb1zfVmQfLlyw5D5zsvzm9GGEtrkpLntvhu/wN
9uE7r0k8NbFgRmCMmGuH1p3ZKpOdH0hNE/XjaC5BZQw0Q+ED9EKbdtj5f3zidBxvqerADaxKwLY7
3ztveV3rROFCbaqEGhuV93M4GevYUHnEyhkqc4+vG9hOkFo355rexnlHgsMXJbGUfzQL4AhXfaed
V5AmhkKDRXH9eVPy8+bR+gtHLwXC4cFUwc6jCu15hK2TVw3t92jnJpt9jpo7HVBY7bxBvwpp3hnC
Sbzt+L2DAv5HVnmeM8dxzDLoCtyAT+As5bATBLTRDJyyHJKb1kwOF1fhwwBxJ/Q+yO9Y0A2yFhPJ
xbFWfJHmTC9n2r8ut47uBtx8d5cSxvHQLJcMF5y8ZyVtGuUbacgETrE4JlQIGSJm/MNfi/FEOCYA
QoztPhjwRzRaO1gLCNedklFLuDkDuJlDTaoPt/3eKNGDCf4rg2Bukfnl14kWyQYQhyjmcP+LXqYK
5SDBwX0VRgFIQmGOcaV2kk51CB0YTwU7iSujrFLdgLgN4BKIL9k5+ZVR7XQnCRrpeA9LYVm1fNlh
LlBY4ccd61AM2VueSYqZj3GQ/bACTrZMlSsujYdR7pCfTNvhQSCJOzcP5OlJFpp4ofsFfykIZiSO
bzXzAG1d387V5N6947x5skGKiJy6GTp1stMeZalDV9ZroP88hT8HdH3KqcG5mFY5rmqZGh/dBnk7
jSDBS+NTGwCNp/KkkkBVjYIyeAdpJmpcireLSdKOKPgJg+nkmWbPRdAjxuh9u360lRvN22M4AWsb
YUNmrXWYG4OarOP3h01btkbamwbHChNFb1W2APtp0HA7/GrDUI3HNwLJpgYb1qduQvkChRUjvgyy
KQwStxGBknHBhr18mM925fmXZtk3LpmZ/diHva5CGQ3c27kVxJeCzeFroaMUX05c2FZCfWI+D8Vu
YCAe2CcyPOJeRW9V/tf3/ZczQNTrkYh9hTPEa8+pxMAfJ+rMorQmqakDFIF4x0BEkJeGc2OED8Sh
4wfhPvp+Zg/TosIAtwEsCGqAEzOa9gRv3tZUlE2HJYWfCDMH9kMNGKQy3DQPliRFp4FyM/FdAAtq
KNGEa0dJ6c9y05UAOT1pfIKdzSgKlSjGkjVf4MAqWqDWXEwtM87WgtWasaW2bTT6tJSYLK5zj9WE
3jEUdwDWk2+EBsVmZ4cN7xW7+ie0GgfLV4vhvmBKL3rexyndlrHFalItQ+cMIsbIekse8MWERPrm
UvjCanNtWa1rgLRVXn7nrbImv/Ga7wND/bBbhCA28u5gVsSs6NTV1Bd6UM8M/8OfoVC0oh/EcBrS
1dzKefZERVzE0brI94kLQrUD4sq1xCe/ndWXEhdMj8yvCvXMp9APhfbHh9P3fatkZvGyRKubwTGF
asmCYai1yiymBBbVxLRhzee7MgJXYTJDfpFt7NRcQR1hP8JCiFbAn4PyxLNPK4WtKG6u41t78EeM
tQKJI6YFuPsQxPXkp4cbRxPDZ6+PT7mCBJNgfIqWHGLXxCkLJPNswsKj0KR7HTqCWnZ5TEEOOXT2
CjzUFRlSY1mezPkiQBD/MysT4Rv81MmfpoX97xuxBOA2l7VbsvTBW9nLFbE1fsphn2x/owQ8124q
Z9aWH8YcOYT8ThtLBnd98QW6wX+TbJbOJU5lssgyuLr1ZdbAWrJXZRGOGD8Ysc9KA3mk/X9hgP26
GABuU8dBlfePTbj2H/Z7N3GQOROvRszEg7ujgIwV2Xq7cApjqt0OA2i+0FAZ6b5EwODIT7/z56+Z
nds0/HHz0y+fnsE3739NjX1N1CKnqiZcijLGDJ64fb7mKgw9XcagwbDMioHsdFAake5OJr7mw8Ze
5qFFgv5WTi2+MbLvrxWXOpvp8LZ6OQ/jcK7ckSQ+Z0L2eonXygpg2ACntTJly7w68d+1YIGcL+IQ
OMxonoBjAr1hoAuSfC/Q0cf8gF9KaCQLc2QhvhcHnm/Zav2gFnWQkpSp/pA3jOQw7QCqVjQoWMZ6
skTzaFD045dcMjlyQfu7M5UDXD8IEKrTLRiemhpH0i8LR3WL8yM6A5qIJ9QpRZUunbdjJUKr9939
mTZq7wD3mMXkz6YhfmNUQDi93eFysOvmwtFOmFXt7kOqXMZixXnvyPSp2vxfyXdRifY6Pw9cqr2u
UOt6Kgq/Wlkpxglcw0uY6VzyRxYXSuj6Pq8EDlgrRligYCv+o5/l/imvUiVMXuTXoTY/5KNMCm3I
uhwtzDh4qkTiS/XOrr7yt3L5G/s1X/3+gbXUifizbMUZYxA0s8Z0ZyEO9QWLx0CchT9ohErC9ziB
Vzxxq8cmqng7pxknUOwi6e0GTU39ZW6oKw7+XKq1XUHP8jwth2ghkpq8n6LOC5huljO9nb5prW+i
C/YAD/JaZ9TF6KE+GVa/pFVoxx30+javGEuezu46PgUedhYtmOOxxPdUMohSSLM8MaKeL6z+lD9Q
V/ln+EJy1wGpYqBoLiNC6MxzEyIYpqwVd53XGXhY8+ninQulRi7NryN+UKewWLjkQ+teyn6B7gLl
SjM3saa84fCPviRfR5K6HGk3+2LIQCr/5kUAa8qPFxX5yLVs7sJsXOv5Q9RLgVL+mR0CqhDlJC1W
GsHzjQNFpY9WrdUmqvN5m0Db1rFJZVJM6S+DQG1GAOT2RFXM09MZtpPNJKrmwsrwkd8EdBtPq/FL
5sOSto6Cb3Jum96vzRxKvtaPty/G4eGDj78Y7YomE6AdoJuvODkgjOkLw0WwenNWqkEK5/X2sJWN
1s2DWMBt0ibD/tISM2o0vBsAAmlXth0ircvGoWtLWEd5+oph78NaQ9MUYyBtA6dwEyAFxBa2VNt2
7E6JlL8HCwH1/u2TiWD0k+3cIFydy0YRhV6hniXyq13/zEZO4H+VMw6B3sb1QCEK6pbaD1ugd3Ak
mDIqQmnryVVqQjKB5SfTICR18wV/cFFeJ5z/nnTqEYIx5JMtfjVuUpery59rZcw7nEjgwg7TiNxa
XM/duzoSTwd/+K8SQwPovO+pyIX5dIvWdH/j/tHj5Fwpw4zE0bde5JzsgZRZUcQXDPwTL4x47MTM
/W9sEFfWEuVw158t5H+iT8K5KwhFZ2LZQKRrSAUAKGNLI7T0fC0UcRGlGobStvL/Ng64sWC7o6nv
gEzFyiqHOL+N4xGk0Qu4+kmJrNaPwfSW+gVQOd6sMw8iqntE8ZKjxbEzezGcK1RJfE89jyi/ht11
lMV/r/8OzPi/sqgBt+DMPijlzXQxGgCsrTj5fMzruI9I4hC2wBVkJSh0W1J3ulJQpYeMxQIPDrER
+CbS4qhw9K2H5OPElEJMKwHPrt9rpoXEXtwxrtC5KpyRMG0XRwwtmq78ZlP8iM/4k2gJBgtWh2v/
KNBDBpKuj3RtnoB+nXDPqYcVVezgEuL8bope0h3LnJrWSWEe/tmqWAlG/rGzuYdvaoC3NL5lvCXP
6zq9E1dqpdoparwvPoMR7pmMBEOLoYltl+CsJCkoNp6PTq6dGV5Ljr3fe7nlCLFma3NMf5/+lXEV
UYt0F3mk/B1NgNk4fjoY9fVv028zjXujhwf1AuEU+AEHTRBxB3uAZsoWHo7EsoDfOLLlXaUdMIPh
9h+hl7tuZytP1NAonfPWbaRYMHjyLuYus21zmFCARn9vdKKQ/LN0u0P6RaK5nNWThjyjIei2Dnro
57YH0+6vCt/HsTpKxKnDpV3PbK65r1GrLfHgM7Ywr7GLo3nefQG2OLiwAE2q4P+JhhtWZbhOSmdY
wC33w5+4kuEZ8UpgK8XS04LgVM/JKJK1LT+nWkRuX5xalNYQRwLI6lkCZi52ZsDAj1VgcaQujS7G
b7JN92jC3wNdzodOt7B37e9TaEH2DBngj3FcBXYoQ+kFKlD6OtkFlrAZSsz/XIXOyA3D33o+wv55
lpD38/PaXSC3O4ts07VVU4mpl5IMiXYFJSKJ6Iq/5hHEVrS0tHor+xpVY7WTt8q/bD2QOiuc0Had
LOSnE6gbt10MIwl409gSE3BY9ueXNT/RZKLsEPpHBXkYRRrsSzCurdhH8A1G3z+7LvdNg4gzKTrx
MMdJGbilkuGkfqY4j6AEwHPNpZ4NWh3V5UBwo0Jfsh1AWKMaE2mcUHYJk1odL1Z+iPyUiZNgfEkm
uRJROAEpW8uny5i1yunKqkx7gPfB74dMD55xdCSv5vd2+P1gUUrGYrHCW53IrQifWgOd1uDnhcvk
5rAjl98mlh2ZSSMMKhA5kE6tz9Pu/FAt/8yTudjw/NX5VHb0L9UZBygOPEZYWmyhRPm8S0/qRaLp
l9ZTQuNfUs6hEU6/s/WJwkzQUR9zTwmdUYiEOTAiStuA8dVr7hpBUhUVPRDqAENMMjpPBcb8wBGZ
hpgjjGmkZs+oVxnh6XUxZzSbB4vl5dNSI92jAfPg6wB0Ym8jc8hP63pNvzUqph5ZsYbDk7BbmlRo
2PhRcwSH+VDwyLCI+EDrF+NlEH1CNE7wlGdq4tujqzehVwm6PNlPx7O811jwT6Lir9U1YISpCKfb
r/aNZoQnsck/TpEYx/eK8dD/nBVel4eI2/gZ50MyjN572xzlYXh54T5PdqDw4f0wNTVM6FYGKtyK
MaJsXT5O2CXIdnqHkHMywymoxRaxA9iINrrWPHFJqNHz9HpHkdbU4HnT9PkfxtiPsmYol9uI6zAM
njUz8gJYfXhKzBNezyTUyDV9N4KMMt29zZHQgJXowDtMY+1oSzgcdtgqEiDXISQ7q26IuZlMuVvt
8fO9ZB+b0BXb9K+BczNspsX6rwEQ0o7PPLQ33yWhOriz9KDrXGphG8Rpq9HKiU/baBYPzrEfjHdl
29QbIq52pKXZLhi6SA7d0Vq+oBpKJJhUIad6HHuJAeiElT8A+x3TmRR1GjpMQg2HBwrqEFjbqgjg
wOVgvd4mFBaNhOpcEDu34eOrif8VcVlaaH7BuFVfmSRWhJQaFtX0KKrVnyxKoNunoQcfzxWL0pNp
wIe6zF/iHkl/uBl0XBN+La+qlVb2JedaIRUXNdqrUCMkUXMKtbkJlwvS90k215gwHza9Hp+FZchO
O39Lj/nZz7MIvmIcr6yogSUM42GRsV2M+e28XkZdaekLxXgPdjzYhw8dFR66jRkUmnHMHnNoAlXf
x9HassrrMgVIE+nbebPygyC2U25BxULMwydIk9YhePQz6mG816vM+rTnp/aq1zQjIVa20jsaRXA3
cKhoVFI/2m9KwGNky02qZO0R6MAzKazw4kNbWFQqVzeWPSomXZCbDOXyyglxGAWtPK3Leh7vMI63
V6jPTBfpRrNe2Hup1V0U4BoCFelAfIhePQqpZYhxjGVBUV8fZ6rcGHDOuezgnxrRtT6AZeK/J2HG
qZ7D/7lxvIJgpnl7EeUny2uN6y3sRu8gmq+8mS7vydYecOff0lOn65ubhS7urzdOB/4rKkvzf/jN
exsIZjb4yYCOAu0EHmV6fmxwnkE4LHf1oz3cSxLitGYKT75WjKre02FYvADPucogC7n6aJVHX63q
AGAJFucACfLBgInhGXDsTgL3H3qBC5O2fsvL+wEeKuevZadKF70iqj2uYhO8G+OdCZ7uGXOoaQDI
RTh3oygkMkrzLwxsJcIjrV+QXH6Q85thMlO2eR5ULbsYqvFVZP9Rq8xkw1CF1jAQoaKDWncBPktB
g0Ler3hyNDaQYYmp6A25IhqR656cpf/M+IL0yxtDSDSsaUEkzq/PHAy6HTKchRW2G0iPDAgFSeq4
TPn9DlUDpmgVMRvoxhsEkVgNGOr3t8lvvI/GgZrZTdt9Lqhs2d9xNFQqbsC27y/YdeswyV+2RmzI
ZfFw9sinZSwkJ3cyoEg/mspXsM7TQ2qFNuq2lWwAUoBTCCDcitxd3ppvlB9yZZcZWzkKhxtic8Mz
L45HFKzadVnyaImX55TODigfvDQ/XIMeDRUQnnGY6fSojCZTXofm3dGZ7eqNO4ChB+PqnMyZR/2Q
Iop36ywPpAVc2lGm+X2HT/nCFvABjhSvdJUdp6rwzU4mtpqCfuuVpZJLJ+fFPjbf3rgzniC7DzvT
Ql/LlFP//9pqrnBQMXC6s6RinUoLUCDj3t2xZH6YF0LGPCe2TEwSbCXMwwJwvyPwY5lhvwIIEn1Q
SAOCVVsCao3zDK59a3T7WQo5AvB6MwdZ7Yh3lv62O1vzNgN1X4w33kof88yvB4eKU2psQX9p6W09
9GNbjeLi19cVQj4lEVoZvFOfoiWzWRO76hzUa4/56aI0Xrq+uhGQZAFhRNlHjT1DZNI9g0eqgSuN
df+tkorjBxa76lEZsOznztmnkv6uIHYAGKzvqt0hxTDO+FglTIrVz/xRbBdJwMkFsMrG4SzHW+vz
cMaILPem6eqLZ3eL2Er73OjEAUPNA/fV4zrtVqiayButCZDq2myuaRwUe9dCetef6mrmcbwuFhO3
KlBG1/FhLDgYL0gwALUYAH5VKrMRpait1a8N3HIsxPzWLq0/5VLOnhmwgD/uYL49lGgbaUx6VwfP
IAbOpYZaou/b7awIKvDWq0KNjgo5IMCrlBspl/wP2rSkN395UYM164msDd3MnirqA52GzmXoTuGQ
e3Hn41lMzIZdNvSNkEtBgLnBMA3D2gG6XJEK6SbHxiQKcZYgPJrtqp//FZImr5/KTe2GtC+XclUN
hI0y/pj2Dvv/850+liWkJDcUtQwBGgpjX1AjNBxp1zFc088nwol0++7N9B3UIA5mS13ywaUIN6yx
wjOLxAOca3zRbcYHDjlpJvIFlfGZRTbFeXlrGIc2ExOT4nZYpnI39sdK5UZ+D+SwxOfZ145kcDHM
Zcshcr58n0O3ZYi6idffMKkHgxGlt59rnpdZhVl2LETw3w9wrfeAjpJ5gnQH6UBk2e0WNa6UtrvG
QETcEwjp6zCTWMPLGWlst0h2J6k0wIa0hh5btduceS3oYSDNvBIvxb5paU5gaBe/xryzKfCXnfjh
PtsjgB6ZPNlKdWEV7LrSYPjzOJ10Vz9d3R3hri8dNQvTurioVYH40ATM67Ky4C2ypKtPohw2m1vS
CGPyIf2iMJLS6rlf5mrPRsmxHfr7gX1/EwtoKYp7DbtNFZ+P2t6SUDxFyjSbXoVbxpwqmV1b1SX2
d/bE6mRnYWczsE/Ec7fCLHkum/tWzyV8bEr4Q54eeFxfr3+ktfPcnqYzCrqoZUIx93w5Hj3vIz3b
cF2R/P1iAqNpdubZLK0tGJcyWIHWsxBu7mFiDLYDkFQy8DpcGAm6Mt7WYf13oxDICGy+Gl+GxVaq
WJUoArVakiKXECg2kA/KWLpg2iiUbGfg/n5X6EqYeUW6d3Q41Lr4g7MpTdvQ3G3in8bFq/w4qt/Q
X2xxTNcif+4reBRDW0A46c+Ng+tjMX7pLSiG0SUrJQrpLOKu5fozfZKM3LAXW+h4XuQsb8cepkA6
gs0D5G7Ibo2s4e71dqqAJ7izXQ9OuI0gp0zgU4RBJxhW3VAxNxjg/woPraxYNivN3y27Vf6DpAF8
DDCKv0OqM/s+u3jmCn2tk2KC6j9RFyaIlXEOTrhaVespinZvPNFemiqRVJbrELeeBgqFyWpcYyYU
NMlXj+w2eKzRCMa0BAg1IFjowHcsVx2Ij0b0t4R8vTJKmTJITIG5OCXVsPjALbH6Ugpzap2ERvQn
LK10P6EQ3EFDgNKgbD/W8TolIbxDqqrqL8pfU4tDrvmJs2faRp89mTMOrwlLZ24rhbRh/kvNqTks
BR3YsjepVKQ/hQcd23USIui3ciX320IR28MFmm+CnALa0ONIUTBjDNEP/3Fg23MS0y2+UhzfOC/X
UpJnndawyWE25y2SZBEEvDQO4HFBnB753J8sObs2K09QXSCkqoZYQkTJ7a0MzRB4fVSrAKOF0yLJ
J7TFXXUftTm9L6leE91x+c9zfmQm+XiT3YWcYz5hCeyp9M8GLtWnxw+2WjEi/quLJcwUfVGgY+tc
5wuyOPX6QEvOlrfbR8kvP0+daM+RPlf425IFsKWpbUnpMe2B0Vl3x2TYX3Nq5jk7+O3hs5otN5LC
Cm2WKdH4+uShSRBv52BIIxxOnzY3WXGhig3I3GRAgHjLLSbrT2ldBxeCOdzzvuZPvmgl0s1legzM
sU7uoRfK8yiFVnhPprGQbfiRo9BMjetHboxJHYlWh6h4PM6l5HCoBCX832qfwKohYnLFDO/lU8+j
zOxwO2C/8ZQg3dRXJ2nhCss+IPLdZFOja0erhL+gaV+ubPcylCQjJsJ6HvPRdTkwl9ZDvQ7Q1C76
B8EIpuYhdmJlYtJpz6iotXurhz9OOghNTCLx1zPg5Ntt74BY95INGpCkXOKUT1bNaaHbiyxv/zMm
ylyV8W1OavWUcJuUZnmUPIm9Vkut9H9XJGwwNJHvpDUF6aYeyMFsg4Ybk1sORYklhgyuHS/I7DMP
nBntc9r6I9+ZcYAhaYdvK11/EnYuP2scs9X5/cE8on76+AGudsg30vICXoma1lRj62DQ3paHBWU6
rDD4fXNER8HdZYlUIPqT3tz94lBctbnzPkQmSKQBaHc95htl8QGM9itKssZMVQsbBkUgcWjdE9Dn
gfAPDjAWmbRYDHJhaW+TIs2Q61ZjOmtv7AgWdH0Soo26NFXU5dYWeB+6dCkwcol3LkaOdtKWQLQl
1iBvbcEIzYuUfLaNHky9whz9It2xv/dMsuFUB/45be9udojSzajVMyHopauBm8XrQg0mjNTSWz4E
omOmXp2A2HFiO6XRiq5dOvuoDs51DNM7WtEm6JEU3lBpDgVrtMBhgmg7UXqTvYVPkYgQn5c09H2n
tOaP1jiK2+xkLx1dkEYsaeS5gjljgAA0TEXBtrIwwQXFhcr7XpvIJFuEcJSY20R8xTxs4tiI1Q6L
5+uT8aufcIVVe4F5gm3Rp4xlDznPRKTug1Mk3g1figjvORAHyNxE1bILl2TfuN7RcMC0NpamnsAB
lsXCjB2U/8OpX7SqTJcgrVHlSJbyJc/174r2n1xI0H6hy0tTH6tGJW1fdAQulFNp5K6d77LisMF/
wKmjxH/WSee+7Qd4kZUBlKuwxNBHEAw+QdE+ixK5H6vw2gC2NcrHXsvoCqM7NEuzYIdPmYsO2L7R
a1zIxSIRERw1qD/UwYy3ajjzodpFbJl5yoTpPlYDNzYOQ0j7zI00duO/IndbExwEW/pvST2BZ/X+
7zG9xDbkj4nK3DsR7R7+N3hI5BEoXboSnCU6Z8KC6hlCHyLHEy4KvZr7qnBL6GxsQuj1hHDAK5MF
+vQW2uaiqdTOrofUmPeWAhWyQFfIY7tBx/kqzDPM3PRt83XXdWvisdaJC0vC+x7yrp/5vXfnFn7z
qXQ3dgaIulay3wAvQaLLMye68W5wmLcIkvvc2Sj2HyxkqKX8ejlxsAvDWl+Z4ilH0RbT/Mmfgtuo
UIOrTdmkQonIfN0/sAZNsunqeuzfUZIjrYlhlJgwTUxVyoUtVJCP6zHHPBRO1DvR7dpC7sru9eeJ
FkegH+/pDY4GuUPGFg3+lbKjRQORV3pGwDSjC4xWxwYn4alm8XDSlqzz6nGu1juq3fm3miBW2RhL
0it5r/17YMJb8XsefgmlaTb79TanZ794nI5iB6SsBRfGi4fkTzNQLVswlEfsUynstOEBjvjQ2OiB
+4OyTU1mxrpGUSn2s9uaTf55dlsxRUh4315oG9zOu/cFjnbqw/qgLu3Et2HPSWhmgNkvtAQyAIuA
EajrvFeBKRAtzwmZSmkM8zXsUS4UkHmRMHxm0/K8gs8P7wDimpWehaCjhu3N57WO7puVTJhpzysS
1wdzUryB3KDbOTaxYJKFKDOnf4apG51I5GafFAwvBImHvtOCqO1FIvrKTzjtDN1sN+Y8VkSCXGur
AELspA3CDGIHkFd9QZZOfbVqr0soutBSf5HNXOefbzSRI4yHnb3sKZQ2Z+sAgLnn2nhvl0Itz7kI
+Vl6/tvkpvUrq/bMf7ZxmV91UwYHDCbvFrxfwNwMNAxp5L4QlCaa6/JX7dtb96YyMSl4ks+EbXPG
tAuDGHKslKkBSZqz2XdNSGYaFOAKTVQgxm3p/qfiXsRDqVrWRslaWXko7l0sAx9AljLyrlRmeicE
ZYc3sxAms93uYkZWf9sUZu4metzxIvOhWJZrmtLoaAHimbbRqsqfX9GYUlvKQIctUBkYeCjQiIA/
VVGZPtlgBby/MLyX+3LNwqjTBbbgS+pDVVzIO1Xohwjwa+zrYjIaDATmh6qVGuAfQO6qjLX150iA
66Ard2xf8Z4hZKS69F9ckuoepG5y5HWzcFATWIUvOnLfsAJJlYEI0b9sST07l05Hgts2DY208XU0
sYZuM8A/g10eu/Bo9m76OCK0sPXenQzBzS4VnSEEL5VpwONWEqIWR1eW0joBSV79FKmDyBGn1i/Q
lI0Pt7L7hpEWtxgmSK/KtQZwoc6CgEx3xoSgYmATystev6f+fDH7bhxY+heNLSLdYr+ZHKcgeRim
qTYdWuY2Ad4XvcPET1U/t4Em2zm/p4dm9IHpUT5KS+l21gIaDwtBJqoKzhzEasdYxntJ3zCD1B4i
KQWXc5jMOo2VrtEUX1RYVxBEYruuBqDNyEA7XbIVEFqdAlnDj/+Qbi6Ly532eSnO50OV3fe6xlNo
ONihMidORQlfbnQZwWHJQQKtdkG2TR3ED8CHyK2DeMaEirK0KHgk9j0lvpXRbk5RK7Zqtw+347fW
alkX5dN8lKdiCXYjNu4A+8rwRoxkxTP4EL6+EVGJKNwzK8b8nRN43mxdjFAu47VvzUceKydICV3u
wVeaoc4bPi2j17M+QZmudGXucM5+/5Z/W+HcbA4yXW+wgBLG4jVuI2IMVZt47oVSo2PuXTe2zb7I
LI37TUGWpgLdKEzVeYWeEVyMkJpbUYZdy7kCi+psumqChH15DO+HMmAVTXkTtPUIPAeRPgscWDxR
ltTulIvRGE09hwH1OAMExTQ1Y8OqSoINoMfG6Z6IQkHhr2/cv+By50fbfXyc4tiTLb4z6XQ97ZjJ
r9rWRP1gbEfvZmYBroIZlBqjaWGQ9hP/UEx7t8L2YZMbckLsUpMHzV8D95B9dGX/nmUBN0slOnmf
uMcaBO5ad8/6Pi53E9N+FSZavpWHbJ7Ur0N+KLgnlwk5m3dFSSuLWyGmRfjqZjIkD4FRaCZcCxed
whXKt8yMPPii3D5FPYNgv2WWEa/V4KvtlKe3XLbo+HxNAYTJYDebWHL+SUXQ2542EUbY+7Ri/HM7
TnZ2ccPt/iH5YW/D//cZQ17U7C07dcK8fzo68/nKXeXsLxcZZ0iGFtT7TKzNGAOJKnWrdXohNYbK
+ML2BvqxvU3WdBGXf6aJWr7ZzLCtXslOLwSWPWVb9R8lmfx+CfHZvSSOPVLl9D4mhLBsWkRtrFX8
HPGkfvOaqWvRIhAMBylHMsOiGDzdnsg/bUnBwLTbhHRLHI/PZzV9kzxDrM39jWDz4ukn2XKyZ8LE
LX7Q3CxfYt31KvDM5TiPZlNdjLrXu79eDiWiGZLUxK+xKV2AbLm7WTzbkYoASB9e+K7KJIeUln9L
j8VSafi4Z+ovFGKJVNtEJb+pcn6bffB6SM2J9HPjOoGC9J0S5Ac+OxJOcScfrGQYsZn1wqVuHpul
ETNpnvTky2vxjUTYWPPcF6eDMeN5v9wQZVoEX+0RkaBTW5nzUMWtrt54bdJSFpKGoNKM4fszvhyI
eAO8Mlo7P2ioO7DIal9lGBZ4/aqXfQ8JObV18+C4mgYEwLCwKPc5sFVcZh5Y5NfH6xjybAtgPYwE
HrTWjvz6Q6PDWG6GIXwfI/+5lye3w04ZMudvo2sOYk6R+ijyfJ7AiDfHxuGKHZWlUH2KnZIzV9EW
Tmutw+A8p5HYGJOxdhsQD9Qsj+NaH946fS/S1bQt4y9UDiFoq9i2vEi6J61MEDfYp0UoJ4jCgRRw
hjjKKxR58pFLTm7D5fgLAzT3Yfq25GNVVMQS+FR4B6Yzys0sjaRzYMttiAHXrlmCLDrxPCpyJinr
hPueChjSmJ0cakT8yr8PN7bT+HckeGxwnXTuNBnSShabeVhcJnrmIBTDL/Khlx+zmgFYwBHJEafp
YFK5ifjum53ieFON4s6WgB1wsbOVp9d1jsK/dQjnf5iwmbXhUkS77BN8s/hrSw4HP+hIDmwSH6kk
Zm3wYq9NJUTp28++XdwVl+kdw/gkE6C9CVGcwS2KTYCA/zPYSZ2KHuShQMoBAyZU+0gwBPnYrtW/
STuWyzboWwVb89xrLHgyh6X7k5Z9h/wAyS4hlAfWm/CxsIwHMvQjbS4e/rxb/GPvLOR2R+lfRKry
r0D3c31pXY9o2Prg0Yt0qkZSOpLF6RoX5q66KKeql6Jm/bFWmPHLSXKE+PXIh/2UM9x0r7d4Gn/9
uHjlM2kTFqnx3bZSOW8q85QJI2mJtcwM2J1tnbINeis6SOGZ0gRRxKS6xgMe9XSC4r+Tw+6a+qrr
TEllQzugFu8UKbi4spXB/zUrw1YqED+a6O48MTjTbNEoUiEW1hwNEGgTKqI3T7Nwh5TjjD3LlAtA
e4jh2P1KPEOw57tB9M8K9TxHLGyuUOykDJvKiESHhxOJAkVYRjx0Ve/YZp2HXaU0+6T9esdi/hV6
8QuUr4pmydsbpBlstpLlEsndvzY4kY+rkryoxd+AdXIDABzbJNmiPcwDs2wsXEQMgigoYwpJ3Vwg
ih6+eSN8ftZRXEizlRhSi3OE25HFd+QbI6caABcs04e6hNENxlUyCbfUDfBsYzTaQm2X6agI4qCm
bj4oRsezB5VqWAQAXSdu+fn422ejsYJodAgxb3l05pEdYtHv4IXhXEYc9j9sR//omde/Jnt69s+H
dz1hrPzamjdhd7uuM/GY0AOQcF2jNqH4CmWOtldaj1F+8XxfOQB1NKgDWDgmiXpvzRbqBgWpu1xY
YQDo49ytpPqVVkD7BvKy1x+AJKhZcVq7oDDZ0UNe8kO/maWYAu8L7T2OHE8MVeKTzcjtfwYl2WPh
MvWZTBtUzgj95LthtlRyT3xuIwjfdLqSQABoyN5uu48PhaEoazz9HmSgrcwQlvTtKa+2MvBdxAjv
P3gvPZ9YjNJGPnK7gIyzTb2W49uUwLjFsRM2MMk9wL/LAvrwG6/oVXf40TtSs+rc5kXUJzV6KGDD
Ee6nEydzxhgAhXQjaFXJrl9YlnyXB57p8kr9nxEKjGbsXPR5AAvXUhg8XiKarRyqXP66q5pxZ/a1
0KTZBq9qcUkDzYdVEhtpqkmAw7MLkwm8F2SuGqJIno8IWMNY1FV+7FjanF4yNUSfWsvEvdXX4OM+
AGLPvcabGkBXLs3F07BsKt3yxskxlgyBk4Shf1DAHaJ5SETbyGNg73dF4rTpm5j/1Y07X8VI0klY
Oq/glRO08Tjx78X4PSftn+b35Rds+0ok7pQdF7fvnq12uhwuhT2aqhBGd0UJSz2cs6WuXA34fWE2
gNgH1IgT2H4iZcdjHgy6kIW2s9a55f4fzbe25zPZ17uvNgWpnU+9MZuTDmptJWNBmWXH6JQxFS2f
knRtxg/V7g+aUbFxPrxZdbepMg3xEung5tsgJsSoaD0mmt8kblMojy9eu/KJ2ZmbXq8EVGyEg/r2
NIA8rlOgiFvaU6nqG7PeDkOMd5UQ3pH7sGfT3y4XU2eEWCAWNZxkaQpbk3D5lNVGF4B4vpisGQiK
uVwzlC1LmG3sJ8Pdvx0TfybjkufTzL5hxW5k9NRU0wZbuwQ2QnFZTyUePlL5nRsRWe1MNRJaY3TY
bsMjLe5ZJ29PBtzF2Z3WvexrKregwFnm1ioQ69kQqT7WJd5iXCX3inhNjdeZzY3McveDZ8ug0anQ
QYomT1sXZFReJm1ONvG8GMN6tIZCmCHMHNXiS6DN3ggDQqwHz5ZXA9J6ZIKQFFk6HcPyk1VYfGXj
qGw2XvUCloLzpeS0ZSbi4dEsmeNTJO+P8Hoq6qviW1v4qA4ZGnfm8+sCxkpp06UkXIkG+2Q7/a/C
AsUIUcb2oUEyKV4tTDgFqHjhQdgIjcK8axJhLLJtohmQs8oareONnKrmXLs3PLh8jqYCKwC8yOzu
3+zzLsG/Xuv+A44CgsG04bykB6OgD2vbYc8BPX7Q1WuyN6h6cWi3pWY0KjwHZ80qsxXSoNhce4ej
7U8JnnuVfKAXZTuKL3HtTKnOs7PksfjDbl5Mgo6O/vwmFOD6lcfig8A+MUqURbLxj2don+hQTGPD
4Vn9WxhWMpci496Hfj5UyONa99X1LkyX2+3XwSVuZRdT9HXUIkL973bvMNFCrQTDoPuWRuk3U0uV
5gmV61fjN/8un12XzUG6dAWjscwhrzk3J2Vi+9K20u8cSelqBchGLkBzCs3003aRB3/OGa39hKqM
2xo2uicINfLmQZSC9EKPXHMw1ZuiSFhcotwEs6pc2TjdFoSJAUNdevpxsvQVAjjarKfBPEAhL2eR
o/8Dq+SSCmgbd1d0dmFjndg++2F8KhCb+2CSThChEcbzJ+os3znk4NPv4+p+s1O4LhdLNkmZO4sp
2TlPzHu4oAyyvUC/F/U2j02+jV7NpH8IagsBlY3RNQtL1cSyjVWqirQEdNABpOUbQFFqoaGEX7GG
/BjoOpBkvzw7Z9YwVlLGQvJC5czVazUvDyy94LUQRE+pD0Cfddm8sLxYE9Z1Im1oOpI/GrHTfBcZ
jIH7tqCP4SkQUh2knsMNUDYUwXt2llsC8vobo2eushjV9BGDLXPcNpqfIBSqiTSzs1SonTr6LBmr
uy345ogV/TzSkhFotHNfpNQNhoxeab9NRStHsSm4XbrcWz/rKgU6yDp8cuIsk7UtyaxAEH8Puna7
zyNuOLIl0NO13ccOIjjYGB//3E/Dem1C401frClyxWjbhkHm9p79TadzJc0gPb9EHzvSxaY7f/x+
+HvN6fdgLLFrcka9pUHmLKpfR4gXkGo4i58u3GaMl/N8GaY5BmjlVUtFCy0pF1eDunZ3u6DNwgdE
MgNVF42muzwZlQ6RsEDOlB2YttB+hzjaPFqMJ9eFgXM99/Wiu8e8nuQ9MuPpSOVwaLRaDHbnTBWg
vHU9xGuw6DzsPlePfl4+MeMj1qJ3RoBSKlBJgp7TkgKl6oKuyIM4BsJMHhhVaeiuFObroVvVu7fI
4d84SXV3OxYd3/peXMM9u9jJiBs1RGVSaxKRTtRq6ja8H3aBeo0s1QaCRTdAL6NHzf1YZbyXvNI8
PPRT2ASKVAYM6bGbsjcXpW7+wN7QWw/Qot4lQicZ9Rz/0tNaBk3DK7OHm8xn8/g/I0YUilr2S745
O8PW7S8XKqb3aplw6mBdOr4UuNFWOgcTBkYZEmxj+xOdv221CRTLha2NNq1eE0ggSKRcGzOZ9WGo
x1niPUQQxrY4v454px6NuHNbBBtLnRxUgq24RdXfHokac/ofsUxlyD5dwYO9t9uqmSD314f+kl5T
o3Gbp8vVrsnEDuazMmd6z7E3EINfMBgDv82LVe7AuKoGn0v7Z5gc9aKwzunDvbuygCRjMT4xfldY
tDCtjSMOwL1TDeXKPCw4NZE5Wf4jOkl3vtkHVaE1ftzE/ait6oTPA+d5m28EOR63uoIMD0Hdfb5x
RHrilGnXG0ha9M1gv2K+b2b8ri+agmkdqlvfoEipmJkcCczuXXcpUZZXELaxMKuf9V3mmK1aRtqo
kjQSHg3gQXph4eeL5GXI0OEVuS0b5vxwOoMzGhFetqCorxfPYA9+PtZchxWQQjpDhNK61MNf1S5h
3cKV1cSO4kh/1xe+z9+HeYQGmoFRZyK01wm02+a6a2qG21Bra6nT9DkTO6wgAB4YM6DNLKz43tsC
Tc5PlSLxVTGpxv+Bt7xbTbvyfqeCHg65tS/wgo7otwksLOHWt3tylmpaMZco8zHPwgWx5cX0pyAF
XQlJ5wtw6ws35vzfNi9/+JaMQE2rBBUmanWfiphmjE9fNsI3+X7vVsUO0j+tSFlYUiw7mbzfc6w6
Qh/4b+HGMx+2JOjE44ePg5jGWkl1FuQlqQKI7Ro24PcijFvxJMvVROxAAMpJN6GzjKPmcgvxOAdc
dnir1Ylt0rT7lfq5CPzC9EUShZJjmTggrQkCqNneoSANL14sNtksXZ6yu0x9UN6jD6Nn3mR31O8P
MoiyMemBCBpydyGImKtiXp1r/7oSGQ7nU1DTllbuibYyP0zTJWdppijgBKDbMlf0rxJRgEav3/0n
cDBBe+083Cg/EIRt3C0eeD8I3IvzXpJYUh8HmO1XZgPZ4gpm1cfsN/ym+gfqADoA4z58bUJyWAXo
AhTGQViAC/BkdbzYWV2/EH95mKEbrcyQK/fHrk+2p8Cw5pf4Js3jWDTWk7uFrDZCdz/UcOmc9AzX
EaNUpBo4EhuwYcSjIF85cZiwUSWjgSvmmG3O3BZcEtgO+YsstTMoSuClA1sFcu9pS8zB7xO83fTj
8+oMuo+f/Ewqbi1gYGtbUuFigzPvw4SfLo9/8zQDTJHG5e9pCVyiYTKd9jOltyxue4TEPbu2f3sD
EZmmzmzoQTgh8YaAbYKkrI6P8SZCzRvt1m2J7raR1CD2ZGZjXPW4U/gtY58dNM8S5+rMebHkDXu9
Yoc9k6LBSmQ0q2rpLQEs1X160gh1B0Hkiotpp5HQoq+2WkgFRPCjR6V/WsiA4WElEEnq8PUo/eaO
iqiv9yMJOTEnXftgW4x7WBZ6Le74aYKqqp2Rvx/THOh3HMaYOsspTkifi7CLNBcqYJm4FOhc47qv
5+zGBrXLO01C4crAMI36GUFOsSSTG8xO3v2cDlmJaiEu1rQ0bBVMecCeCsfi0lbbGmELdsMypYjO
pvQsdS4pzwz9jvoPwphGtL9/Ht0lLq9h6frAgR3Yc0Wy4mq7p000HVJw49wN9n2aPLHv7PRB50Bc
wNbAKh3g//Y68X4fLX/dFBKuJiXLw0Hi6XU+cc7tEgXXlXmQod7jKOk7Ys4/8DsI5t9HBYUxMt8Z
IBRynmrrlDupGlcRJX8yDFxMt1L6zfG5R1xigw4HrFAJAgG8Vsfh/G016qR31hzbK21HDBPxDShy
ycYL9ATA3AGfZDcJRdfvzr5rCs4RvplMHoDsDQQCLaEspfwRB6muiDDuHq2uXaTlJTSy9WwGEs1s
j6GEasegGEl/EUofVSDtEd7IPsw2KVqYYbpft+9B+i2aZTeKeZKgc0Inf32mGwk4LNF4KCPnYnq6
VqPnLJRFEDrsFwtjvIFe9GAefl58e342hEWR8DXsEPtTLMf5h5XFvx3ECwqzAM28uI6LStBK8qrB
NEBr76eVF0aHSAQGF4QfNRlV/8+N0qY/1AQfWSZ/kI9+Tktxy+/+qPpky/W1+wBIc52mOfOXitTr
QlxJmgELFF+kmCg5yg7knZwXOFEtZSYbiWZem7Bzd6uLWo7+h1Onf/KuOTTz8Erzeyg2N1PBRERo
BAeh3QGBM2jhhJzPj98PKV3xnZcxJxyAmgMoSBajuwVHa2Hk046H+3MVk4PYWUTWf2QyVBz7hr+d
gVIoPh7Ni5T328JPLxbtJs34/jo/1VHohvGA/zwtKrP5Tm/HHY4gwX8Cq42RW1kCNqrF/Dyuzdwt
lNj4ZxqiCjdYOM8MsVGzsZYBE2cFjZDRwfnHYzkyqZDSHd0Uhb/7WHmbOT+aVmLYNipDRSJIt79U
YVrW3J18sAiUOsoBmH2f/4lpo1wNBr9sF7QUX04KNcsCoJ0NFucmSw7+10vNgPhdwghL5USa8jtq
3znaSRHj00xcoPDIBa4Ast0bNz9fF+/a0zd5Cq92uEB+6RoHHIjMHZa8sszXK3ei0RnPSEexjUei
Vtv54uiyvGtxEIA6cFveNF99pgAmSzm0L7zecinSXhlMStK/s4+9Do5Tygtv08hSBOdgwleP/BIP
+D0UkwI6Bp2viJjQTHFRK+lRlwzwLi9DijiuwzD0smC66tTuCYh58A9v0HGkYHXezrJkneWFKQoV
/ZAce+PcIFgdULgexw65VZ5rvVILGMfmhbmqqW0y++7m6yvpcmT+E2fTOPjFsrOLKt1LvTsRlsmU
FkI/VhOui2ENYsK0RLHdSVdtdoJCoQgBYMGclJzjrCokLvh2QXv3wPffQvlfIZPyU66+eW6tu2BR
fTmaDXAbK/5ygit5PdZJqfhOiFnVHgoqVo//y/KS7L3VXW4BhJVzRoe3/A3J9E5+ZA3RJKjw7xeO
D8l9rp2AqQBfRK03iMfZR+jn2veve3EZ9ScgknYwKdg28gw2tIRGF89/TqkuXTziUYeb2FWsYyrD
xHHTAVmU/YBL8HZIDMCdhY9IcWP9toZdht+MYkB1LVnxDH8Mz/4j7Tn3A+z6/No8Pe50oyMa5CRy
hELO/WtkWBoYAu3etlWOWBszRhviXSz5NcTWEDwR9U1nCJRwv4JnXTi4VNFG5VNoEcrkFI6SA5aF
5xUOIoszPTEbq81+0RB446cCKNc6pPbcx9GPN9m253niRzStjqHWsyB3+RZZOPDWDdXTpnLE3mwp
VJ7OQbeTbozYLdN4y3LnbzVTHDB2YELyqBIlC65ej7jX9pmTUBspeRYtLY1+2UYYHkvxR2F0w5Ew
eaoS+Oc5/M9psy4QfOn6oUpyZ3l/jObdkfohJLpHu5vP6N1QlJg6F+iEXN/Mpaow0sJeZQgIRDaU
EV2tR8nb7GFSof4EW1iPGp8lXFbVaqiTutKkzU4jK+W2qsAuNieEu5jA0YHPhuw/xaG3KWsYwck4
GYSQEuA8F66OrPNrfn/hiaWb2jla+k1u0Cm5hdwYSu9+RouhHDmjUbFwzEZClbgP5WOnC7mYOS/s
woe5U8ZqhHgACDlD1N3i5JzIEFSOhge+th3HsGKOc927M2SNKVVF0WvBBFMgpVfzeqUUMMUFYKl7
hMClQfywoPDzz0ImKRJ6jj5eTaMgHS+V1uSN90YSX/djLtQPqDuTc7x5szsUn57EJLxLcfql7qDT
qZZExxi/bsbM8+NrCyZmF3i7z/EYMViljjf+Kvx/CXqrU3kDfnIJEr2EE4wWoFUqVdfa061/V754
1W1Fdg9GUZuQOScWO6N53a6sTaVUUIJBeIzcQ18GLh0pIZpgCpFL6qC1ehCRPzjdzffD6Pkgy6fJ
NMj5fIMKXr2jrxFyzPaScPdGlrzLmqYFtQTit3Zois8eg1rjGb6v/779w+Or5rZoztObnmPw3TAv
tEMbo3KV7BhOi3hPmaceTKCHhCif4PfY/2fPLeUQeSZ5r3L3A3xckRMFa7MSltPbi3stCPXvAzIh
j17t+eLXAjb5eyNPT/apxOxCMUBznwZFPUU/MeFrSJY9NUHxp843QvBTr4dtfYW6055PWu1Vjg0g
z7nt3yLEKruvcDgaVldk0St9fB1Mh/II7XiH2iWUR2FA7azE1Q2oY5BNZ99ZYfsKAXjQ8RT3y1bc
98bck7Umk1coryC6/Tv0uKyiiZ/ILPX7S+p4b5XM9ongVhGkcAbdvCZKWmWD0SPYqyPwFZ/QIj5Q
Tlk1F3QisXgGNdB2/5zcaWOZJvk4pcbzXdGxwhjvTLm/bo7/IR0xeBnIScuRVK6p6YLpIM1iAbOk
YlxxHZv3ODxtPPpwh/kVzyGxMM6m2O+cFQB0H9nR0QTHogKKMcu8e2ELM7u24lhwW8uD1OfETBXK
SnPLHYJE2M51gQjl94fJdB1ufWx0oLzAuVTjVbYrWfQDDygpG7S6he4dkiMAZbATOeBu6049aQ0a
SK5Itmat/fAJF79jRxLIupFp7qQS7sW3SWMotrhnQympBs01t4InjncUxYheOFoyFjCkzTqklM3Z
2avDfwXAha+L582YlPg71iz8KI0ZwWMVTfVeBrVYz4wJouW99t/ekwth7E772nTpd+4pd5oC95uv
RR56YroNQg3FHYme4iXPvcQqj639LIrvy2HVp5ZcUN8GBevo/I4Yw4Lj+9hqiCsQjI7vb7OcKl1i
b0s9tzUTXGGBd13lYcY4tzBEh/3xkAC8ofdrE3w9BBdbyzO9R9RAQjOnm68IQAJLjQ8+10yvaSO+
yJzNTBVO0HE99lUaM8yjpqpaPU9Qr2CjJnD5hdCXZMwhxBaKHfdjOXIUrE0DhlL3izWe1xxibRfE
zAP5OmItwH1taI957cE3DFiAmPp9pmUNCGjRcGR3nS19u8NhJooUK6gpV1DaO/hxKYdf9RSVWMkT
Jr7lhT9l4cMdwa87VxZdNBb/hlpnhOkXdCKMXhVKhsqh980y4nB+XpHh6jK6Advb0dTDlctwT2qc
kic51lExVIStOPcSRa/BBgmx7THnjT/H6hkrRMnnheHba4UkxzyDOTpGl7Dh9HC+poyrJyxCEkZ4
fMG6sOnubwz6SGeFovNtaLldYtwHtqKf2QvjBsktnJ1YIxzeDeykyAjpH8xYOI0+0BdmaETlNV/x
hwNbL4HAUp6tw3vxV/I/LbFP5RTJSePmOtrJt2/XMnUlx3Etl0RM0SEB3GcaBSItbg7TISDAV5m0
67rRBhGT1EdMePUkryYDBJH7axx2kWs0hUEMqOkOrSOSs3Bzmrk648ZtPIQjD8Xbkq7W+e7C+P69
Y/4mvNIVC4Xzgjdr6lOI/Xem4UB0YS2AFjV6Ox0wjuWvsPRxydMcpY9IpmT8jlX1464j7ZpGz91+
tJolHqbPHdY12bAGrnZkOoecLAAjWPmCgcLv6+nBMWfZyhTrIgfJQliabNPrlg+VRvzJyS0svd+B
3gCtFH2DYIyu3mrxxCDvT5i+IR49RVzIyBe44jIfb52EFFKKCwH+22r5Kryv8DObRjvg+AMim4kV
IMTlBVxLwT9sHy8RVPq4qFs2OiV2XIva0M+FCXhuVRMGytv8vWLp0/DFNh0J9xSeLWPrKIk6/0m+
+R41qNVfLPKwuz07Fan9dtkz3ovnB3Z1hc86qeJPtdJvBLIW3vX4iJAOlxDjmvk42GWMQpCBgYMg
FBiugRj3QZoVBhUbDLq3ewTSmChW5FzwPLiO6RI4hU/4sIO77yvCkGzDJVae6+GgwDELBcePgn9e
SI8ameW5C5bt7UNf+B2AFolSEgb5W+gVaSjStmlZPhxYePdekqZFOUc2RBPSEDOeIevuh1bH0nZk
vBJbLqy0P/hJ8klCU7/QFxXFKE50vdoFe/jRu8VV0IXsZUEbJ6FHhJxrbcIw3JZ7tdhx4TRR6b1c
yBFT3R+fwZATxaF8kCAZ7KAJtDOTTrUATVHqeopYg3MVSwEwSDRV77S5tbNCpzXhUQbF7PuWe68T
2MqcqASMl82D1v+T9Gj+gpxOAGlS7BVR2ejUE4sC99nsc2bT++p7j0gbpciB4V5p5h+jhG1Qidup
WnQswtGn+SfstqZ/sqe0YmSHiCAp3BJeDo0htEYjlv8IRcJFDlMIgCZ0taIUipuq1TP83j5UtZYx
WiTLY65U/KAGTCPpNgpnA8w9fzE05LYV8ZXWW5Kp7oS3CXXkjs5ZJTDhbduDVdYkcClrvbKcD42F
Y5ulA6pHBNfMa6j98h4f/clpho/DNlw4eeZcQYe4VmUZ6B5FhYKIzpClc92nLriUwWCsRS9icU2r
tF6h93FqIfHaQIowCq3M/Xs91ZNbXJOPkD9/6c7MDOgweYtTsRnTtFM1XnRtQh0mVbjnLazKMAjT
PApoHzeKgmkNTp0JlV8hmO6kDYwHhC6ymfJHFqjGeHaMa8hnPigDgaPh1qQtFccPL1UwEud7CcWq
xqXqW+HuU2icggSS+3bswsp1U/LmnVrpFIVeBIM1UWRcoTKWt+05QVUnL6j+6TCZgwYnxfI1AAXV
vIy7I4oErzwqlIGU0KXyrqozPWhvSeSXXtYopvt7sSA0fCshYGHQQjXwKdYRgzS5NcE1EyNA7X4c
XOz3ecWu9TFG4iG20ESQOhOGTaM+4kkt3SVCAraJAZHW7NVEoct0O5JtOpdL2pHu5bwQ9vtdogj+
xQtQY9UnBJscVJP8bFyEj/5akoTWVK7DKvu3QGGW09ujPSU3Bjj51H8QpRc88oEtw5tuqbBvK871
a0S+7UMPSDyNDp4L6zStYoOlj1jgQEi2GhIIkumx7OTmu2nwcQXaXN91uU16sC2TvQ+PXyeFg+FI
YsdgYgHMb3J/ZQw+MYXQxVvoIVMCk12OC4kLu0qgxbPyn6I0agxzC8P1qozLxsKvpdqf/e0s5lNH
ZmPxl3Ipxv/33PskO8KUNU5x1LiqrnwWSLjctXuX1jZXnyejnvcXIaw+ozRpzYJ9gGzw/S2MGPQr
P/OaEyrV+VcySsUEqcTaDO4Hg+U5KM9gOb5ISX6YlAQX7zWOvH3vnftzeoUICLRZuSVzcrBFpKxG
RsI7V5BjjINKBBMAgzd4sGLdvLdPgf2ZhDNhYMJVqAortPLg6uqZbNB44mil36EsgUxrj+V4AmfH
Z0oFoyC4RACu6V3ehxx1scg9etDC/qXJIj1HbfZT9PcdkASMA5J79QdbpDkvY+0P4YYzDyh9Yuws
xGax6TsGrEXb8VX6bRiNeWeQv3vrzryw6UnPzVvHc6OiPN6kyINGgV+iEhpLxovSrZ7GQQrrLxIl
+QUVl9m2Pc4GkBApNsFT0Fe7gqARgj/zx5vJDnAzva9aYYQvdpM6yT/pDEswDDCOnT3kPOgdtC72
+tzqVisTiZV0HKLKy6/3y0dkN4w0xFbenqQgCd7uO0q5VDMgcj/eyPG8LkdILDcNwf2LnAZUG+K7
0xc5rCLqbwsMuMAEWiZe6MBCVkoSsa8BOciZv8G+LJpD8Ceq0Em3o2fYAok/gCoBFRTEsx+XEWwk
65m/HYtLBlLbuGAkH2ixbrnwauZMd2E+Ui+Hq+LfDq1G1fyQNbnU6DIQvTM8Kafi7MDcC7uCGuqX
CWn2zlx4jgw9/MGawKlIqxpKPyD9fyckg3GSfXFqV+UzWvEmRlZi/zgnqdvJO2dFxCh5jcPcQC1p
1ycDhmp+Z7xDtU73x/M7y5yKK5LgT2TtmW6iclgjO3yNNbwT1DWMVnj+QECSLlOv/6tUptHXhgVw
4NCrwsli4uWXamQCpQH7WqYOc7F+OvjzCjEC2p0icGYVTeB9SrZvoQldFnxJCa7Vl1Sr5FDchMKO
Z7BXwep58VA1F8G32tvZ8DKuHfR6aOwML3i7tN1Jc8lwDwnjMmDsA/pds0INbXkX/b+M2Ct3goVe
053+kNfrvjrGmBdKTshoGG1VQSPp6sHF7NPuie7g4KmQzMb0VVF7xzhOLIGLGIl5GzuWN49COLex
uiUbyLDTYkaXGw+jm50JZxurnPR5UaNLIRlM+Nmj4on9E6VqhfxhaZOCgK3cZNm7KbkLxv5GkePK
R/T+YekCAagh/5QMcc8tOxhxaACDNPwnrQV2C307nEJWjetFd9zs1NpqdBDKt8S+WTvlPlWWfVBw
MlrU927dSOEXhGz+NgXmOLzpzi3M7bpI82nEn9rVveZuS3zuCSmH9I4jT/vjgslNPZuXEapNLQak
z1Am4kU4a76JngbZj1fyPtxKtlbr8cbsiOl9VL/G3r7OQCoC7CBJl0wseKUmP36qQ6NnvRwCj6cx
FazTzJHByYETJN0wXCB8H571Xgt5g8c6hApj8hIHQVABn9rtD1xv+++uQZFFDbDF+tJFw5ChPl5n
o/uklVAOhinCBsKyo+xvLPejwVent2spOOAdMVJJ1eISoDBgIYSsUC0PVpukqSlhSyo0b94tfN7d
rVQqbzk1lJCalXVl0QBmjJU1J0NosvL4/p6edVJEwAM482OMsv2xYJwnLOJUQ0zb7M4zQ5FwrwYI
Iz43Lricf3OAVCQjUCQvEyfgbyKhg9l2Aex5hlVPsDqarRckliGxcQ6Deb1/+ygKY2W9RDXXuukc
540znbtvAOItmvBjyJzFaC09OSiJsYKdWmCwPf07rrFS4W7+avtJ9UjdIE0gI9Yjgwy0P/f/FBoP
FvpPIOMVRnCH/QI4ElzyQ0N03NoNdTWZey6mwnxEqtYkng+7V+/AhvhAzGm5oY+6XPqU1Iq33sbM
ySZZwMjKEP+wfoOhPDlo7mxb7BEAUrxr6Z9w8XMTzjA+4pRiQ6D3AVLxG+KwMMYA+Y8eqY+hcl+5
tyaGgVpFV0I6lFgRChkLppi+TzihX4l2O3SCM6tn3MxnZTE7RRNGnzYiitZM3cLLNuxgkeusDNaF
emFbg1KyX/j2xnRxdL+qg/V9K6R3xgX79etqzUH82i7wNwghTyv2PjzQ4waIphBNZZGVA+hSCBhd
9dqtUGAWFnUqPmtKi7qcs5pi1vEh7R89EA01sH3bT+C1a3QW0k1kwMB7isBCvZ3mfoc+OqDTKWW0
GKsAdjgDoBapuJUdsbv8b850U5GOOZrqftT+rIyROIoMQTHkDcDgK/CS4u0lQxvYPfg7sP74fuqa
n0+Xkq5TFbVK42O4kx7yFgjh4+cfFT2wuqwdJAWJdNoIdGrbe1PIAjvBJwOVCdYVIBzR8QEVb/NR
QQiUZpnXrKmcoD2PHJmA0BnJlPdC134uYoqjLO8e6Jx8pHL6FM7Qt27f1lGwQ9bAukv9WuRMtFPp
4o/8t3w/803FuhsQsytjjqa/Ut/DTdPua3E3jFBUAXky7LmDC+2ZoR0aVPtMo0UMYhOpONDx2NVN
d60/LbI99ErWkl+rj4idvXrhSjB/rLHjtLcgvZGbZQPOULn9DhPDr5414aE4r0LtTaIrvWx6uyNC
IeA9XfFZcxXfQse0PbWeZAI2Q5Sm7wczloSsR9iX67ycwRN+MkIMk7xyxGVY016k0xr9vGGvz7ep
XeiWyHieowYNXgA3bNUWsSTEnAjBO5n+6X8T9YJghHclkey5Kj/bv787Izl67np2FFBU3lUL6SSE
s2EI5ssvfZzkCPwuWNEhaEalxU/aQuMvqG2l5sjyRRrkCdHGdZ5vBEpPXW8uz+0OsrpOPRxMIvbP
0rnNy7fJj1FhLNiOIgXSWgyV+x+kpkeuk2J7U105ny2Xx1iCTq5QjLcg9X1sWpwFLSjZbzILje5L
BQhhJ2Z+5nV1L2Yfc2vEQ8l2GwMmeaPFk9NxvKHxq8OV4bB2luJThdBV3SLiM3zh1GEuuL1YQSuN
GQRZiOb4k4Q0m8x1x9nVC1QZybhi
`protect end_protected

