

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
c7xxggHXTVqTLOqNp9SGE10nZyxQ+KnXNaIB29bib8W3qBD3E5wqL7p0a44guEKX9DID7QRgJHUE
DDZDL3rhyw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nq2lZPKYocqsOWqzQIKkMfDY1mRu5M5W28mD/gsl0IsEv20UFZPbkGMvAOPzPMKFCfZE/w/tojuJ
lhzHqYYkkLr4Kq8flbR7GJd1pRVcLbgB3/wOm+TmwkgJW7rX9tcmcD2JVbdG4cQdJOK0+64Cxylr
tE/5LALuXxrjIWoEawk=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pmatcigqBUUC49I5eR/BSIBbJwg1ggOOuVwmghOlqg6b8ps0Y2ETJsI4hCcIRjxBzXvOXeVRPa30
P/UQjviF9LgD8weqVeUChds/h8BYkoFogiR9tXAtVRxkbS0SsGfmxC0y5ibJNjJvQithMhWRAZC+
Dwr9mrrtKYYsQm5CcTo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wE+0Gfid0yGB4I3Snko6lAD1/lVbjYM0/KXoK6U+K97kM0ZPMubIIe5j963HoWOouUvolyk8DUCn
+wopeTz3sbZhFw0jKZaUxuU0EZY8LC6Zxqe1M0rkHN/z99cdGrW135/VFy2wdmKEm46TJWZQTFog
zBkithdQNCpkyade743mA0BiZh3GfcYXW975VHcp3dl93e/TPvi5T0M/16u4zYWM9rFHx2jksA+4
WyDHs/zsuw6VF/wp0o7N8lh7HkqlCuJxCLzLlbqjUTIXkigWjDCqaTuhEeNtnyz68gUi44M7hvJN
4n1MKmEREvbdBzZlINBREu4D+PtMbEc8FYDT0A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vS4gb2gRnOSxthJ2WQfsj9If7xTAT++28bS+0XEFknK0ihZ3bFqByxS0n/ooPW7ht1+YRqkP0Bwv
DHGrTFLq0vsWcHefMIyZ+UJHSveyxlI3gqFbCQc2PmHI3Hk1ptQx0iag7wj3U8OCAxM6QEK8ljjG
jwuJynfI3U/QuygIY/+Goe/gwxxauw3UkIqpJIgK7v8NOZio/x0yv8vRcdgzmF6U+StKLCRJyoLQ
PkDJwoGm7d40BPdVSj2RT4NyhPrb7UCkyeSPk+x7GIvXKW2z11dAWd7PDXxWlI0CUGXNpD2sgLv4
5UJi/ugUxzl/Uc4eCoHpsIlrWzZF9aJZ1hY2eA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f/1eMZvZi6ZShQtYgxBNnqftfBNeTaHK0Vx9SbbwUYYuWxhS4cCZ3XYMj7WMeYAmz1xzCHvXD7Hz
b3pcNKlusUVQrCW3BsAGvjIpvDQ74z/9o4pHir7N9rnRK5Esxy0d3rZVu1wPPBR19t5Cgyshydr9
Vwm6f+mXGH79J3qPnHB0131Tn1wd4+yC9PUqELEH4RxLYspNCwtJR0Kt2MLV7oU3qmX7/KPzSXaY
3CP1zTsIkbdt4HvmuZMF6FIhi6B27/hrchU2oO2YzFmLaa46cuFM+cb0bFn1l/57EVF4CGgUf2Jb
8BTWEBELQQYeQ4FSMEsMugLMgP0DmmXZ+W8Mzw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99632)
`protect data_block
WHJu26Sn6nVV2w1xRfZukGtgNTD35H5llzrFJrTyGRt7lrrS0EznNZKS5S/8/Da0BmChwvlP9Dse
UFvsQwc1EuhWBa63i0f+fiKc07G53yrIxZZl5fbK1M4m54KEuXljNQdNMveH6mWRNbSuV7NPCpjR
aorjV+pdLr9BvkjfFpUrajPz2WDNfz6U3SrQUk3iQedo/Wolkac6iYqztdFNNbLb77PJWgyB/jxo
IPiMPvhOh6JadOGZDtlHVfo++wQkMkoSG83SGZnFysbZomX9FZb9AkkLT91sLz6nrDBihQxQHDJw
tU8Hee8/QHR29ZY2vAT7ELBbw4poYqgNm+FZTcr7ZWy16GxSdw4gl9GH1XO8ITX7VBxHY6WU7EFY
wuOzpIeQ3G9VJdqZHebxnSTl7Yn7nMEPAl9mw2VWuBFtTBvrOYMwweVLMZad7k4JO7jNC4qXqmLi
YxPmyGmFHe4opcHzPxmsJyr6nNSd0JTsOo/d5DYDepPC/n6Yid8Hqq43LqVdM5/9vsLMaSwdPiLR
xSUHaOHYpdW+2IYfIBpdxBRA9NAdVw3MSJYHwL5+xocDNCIiMLtXovzOpwEAxBSiesddXCOsX7Dj
EU0YK74ny78XV59zz3oZFQ1qePa9T8qMcTFnzUhLBnsnlDhMkpucUALF9CsO9kFmoSg6DNszgOuN
8AFYlenePnVlQl9TCn+wI3t7KU5kAk/lRAq17WTwgx2r85J8EeeYtISkXJej3/AoXojj0YhdQ7qc
EF6i+gXogpZgjaB/lTY+/Q6+o+am+iyRPoSJFKiuUwG4L5ywrGLr+UMXOStFDzzQwakvjS4lmro5
Ieq0tDK6Q7ut5D0dgkDabeEUy2FFbZuVv25wePyKKqLj69jeOO3jMNzwrqIurbI7Gzjg+nocolQ1
3zPsu5lsrQd+pHNvTCblNcs0XNWPfbLUscda3GoaXtx3YzHMRThteAWAbJH+jokiD5Fk324d1ecA
m/mVSJ2hWHSb3aYZimtvzw1fIjQa0mgBGqZx4rxlaao4uWd/7VFbMdteKwDYRtJp2skVQZg1U9EC
Hn1qeuYDXsIpHArcuGUm2tByg66pULiQS/FaVneSZ42UGRpaSrgiXMy8Lru9t1tDN0q5NO353fe3
FeeAU0HRiR7WoZXiTON/LlD7su6ju+PTrXTMbvmm81TevWMym5fUnSWllzCrJHX98gHdMxtOwXYD
4umGhRar56v+63CthT/OB5IkF3sJZwBc4YglHtYxOV3pkUzWpWLhAHbcqOe2LzMAo2rcDT2hvutc
CqD8su3+j0fd56oKVwySjUNCC2DRBw2PleQO8WU9LzmATyOlx/hUhoJJm7s0WrKZmm8yh4DpXfXk
xgTkQTvd0P9pxnpwXyskiLYVp/ULugmaxiSvpN3S1lNtk60w2TY/igIlvk0Wl902i5+Ca/GJxIVf
3daDQtzFNFQVwF4w9GPG/YpSY/xluOmGZuJG+FIMc/HYBiJOzHGTvBx/Mjgdbniah1P9+s/nwUdc
tiwT+rGZtuCeIjqxG8eEYgZvqy6JMuQidxaCJim7Tapj4yJSQ7wDRh79WvuuTNJZsmWo+UVO8t9l
PrwMqZ/cjnkGpSL67GkPaz/hAMqtGSHjVNDwOLWDu/FJAIotDlljfEgXBpgzPgx6X+B4XvTMbyB4
4oQbWIH0JCY9GYVfp0i4whRUxIUlp0SbkzMRBUJx55xeg1BqWWCmV1SYmzS9Pu4nN1uDKY4f2FMV
8dfCn9vM5B8dKARfE35pkliCjcaZ2RHZV0fJbxsRK5h/j08bD7vEaxW52sEtSKJrV7nzDIY5L57Q
GNWML8dnNa17Sz4D78PXy4GaraKpnQmanlJdRS6k1uaac4885LL4jKe1+TBgHrDBlZj6eUtwuALX
sfb1sOp50Kp8/4CrzchmNu69mjP85jF7HzvWGP8dnYms/3kvtQI654FpAhCOX6rkVYCUpa3DLhNe
B1nMwbS06bSlMuE12rIAMgWcNzA2ZYv1a2kVAyzAGLMYvtOgWmWkhZaMbNepoLF1fh8RiEgZaRoR
iayDAtGUD/TVpy+IE4TdO+IjMITQHKh1UHUONEVotoD3Pa4kyYDmxQNWtR+QvPuDJRgyqlecP7A1
UhFyqG/Gdsy8ZU4UhnAl4swVjbDbWpQSMJX3RqiGAcNINUGcmJOf1GJA6UfH0A0j0xwunGSKyp0g
+S7UUE+3IglBlN9KdpE/0qhvAKHYbTmKlOypQpaaWB9x13JjnIW6zp7czWqaPc8ZY1FW5EPFsCzl
aaC8l4+hdTJbftTsRA3JOCvbY2lqQTwApt5nFRCuXfHnz/NfhgAS1rdXlEF+vkYaigwDY0FwBRQo
lYi6kmxfAkHgU8rzTnU5x8N9+fKImIzRMXFootjGF3ajbuQyMFR5bKH9dE0iDJ0ZtZT0DmrkY4mc
STpYxTQtik9Kj5/SCc8m+VxvhIwQ/kVdXgeJyZUUk9NxbNbm+F3QItnkuSVmXm7nXgZVIASD8qpK
mGS9QK6aXFQcoaDfvpWvzsvo5+oQsGi5fpRVQK6hCOsf4vysWJxiCeoQCwgvzrC3Vw/CLpaxnM2s
57/KxVqJBNetQictt4zvDFAzaNBFVTRsCZme0v+omQOlBwuwV0JqN0iq1prttDpXYdV5Sb6BYJsa
4l2+bWE8lC1mDaFCfW/XYgBoWTZCtaaWO1VnfXnfLSlvMtSarWOPdruNYyV4M4spASEBrYiPkpLS
wDn+LjYV8GoydGlzdkktbJzmmFo7JMvSYwl2DuLQc62Nf7kusrctFm4pLzchHe0isRbxEP9muLGe
dD6HlaA0ZQj2uSA5TYKXomxHXZU5Pzy2zr/kihs7WehduVbAexT6/nwRjUBIDQKfuRLDu075UYnk
OBqiqg/mB/O8so7BZOhByz/2T2PLsvxmdJMnvRDNfEI8z1Wb+zmv6xolEGNXYfOL9qeqwYQZ8ud6
h5zsmr3IH63gXMPw00ul2xakIrqQO2cMN9aCuU3GDX6p79L/fvsZnR65cr1iMA2dCNjob2ExwUP+
sNN0VfuN7MKzVTr/LKapGeyfPbFL0MKD9RePE1L42CgDw0/PQLYaRl/nSUO03OxAdZkp0XHF3M6w
j22cpEyups+5zU7X/nVgjK0EznH7s0KLYFrswOJjJEC5GM9MLL8YWxeleAuztKtmHOnq45i+xEpq
YmVD/zwXwkkWVEGp4WTt6sSJSTiVnGKVGzXaEin695zGLNYKn/MoIetIF1owdMwKAz4jKfd1niD2
sw4YKAyWgOOMpau7udEemkEP91U4DxwZnDYCU30K9aygQOBXcbWiiOqJB7LuRpzzdyskEoxIboJP
Z4m37KXikAfN4mdARpxVcYTXSG35PcliHehgB+Xp0SGYX2i5nE8yEK3irgfNqFa519IOAgmADbUO
GllIp4YTHX0/yOmb+z7OA5io8wz6txL6oYkFj08LK7x3Gn8uQRqSZbzXaiIvVjLGL6DpkOc8SPQc
Ol1LD17muY+lfcic7SsILCXY6FTIhd+sTkcrfeKNC/wZJNOCXzns6aDSBG+CDO3Bmqt2aDv57bWq
/RFy1vO/5YEdGkKYQv2qiCfzO6g+1x3UhtDK1iTR6ez0h6QtOd1WOJM7KRbn8pPbgMOYP/EXAjPk
JmpfmHEeEVM7VL/RAsF1b0nlgmVcFzGpl8+eFY2q2pA2fXo4BsWRpaUF9co+ydwC0x3lthWbAttt
FqycJxsiNZ+7/5IUyuusTjwPqD5Tm9mGRmT0dA2KyKJ+Aq/ASgCZ2bCgn3qrj5QK7G04AmHEnp5h
2+vrAIp7stpbRLvUwCjFWla1rhYDI3mYpgyH/jNQQIRf+vRMIsyFhkWqcreR7F5PQhQ/uZGOSLmq
SsuvO3zcWMj/Myi6UN1hPygHBzKuZ3JWpsiXFL26xaqLi71SRjmwEd0SArKt7S0aHvEpeE8bDUTl
4m0Eo+K8HGbRRFwfq2EwrKI23xpINWzcwi/WZldjbMtaNiBS+DsSECl4AHEGWZHU9RIYQaDguESQ
F1ByNGH/TDTrGZOgfo1NBFNXn1I7nbzNY60N7/71f201a93m7W5pQ8K9NdHBUs0/dXqmVprZM13Q
+q6yjcDgb2S8o9XLjfkLI3WgMKXCqrE0YTL23HKZlPlePz/bDVMgjI6CLco/yJL/b3h6aDnnaCj+
CtNVKbKsKwgG/FMtoPQ49yuqFSqUY0kGnk0qHpGVQFMhFut51aSNmRd53flKVSVFNbAhjxRFVgsA
GHdg/k19dP0Tzwb0MA9YB4OyR/bV5M6VXqmBcC3LPNx5jU3TZBH4k3WdgjM0L805nKO+5gh9GFLb
tGKC9UYYvwEr9JytNu/4o5mVnxZzn6qIs4J3NhiuktcovhmFC1ZSyyXLP9Qn/9evJAMcsbgGlyVy
YGQJ3CNyxAIPTlX+ToFLh5kdCH7ypBxj30RR9VoweNRiFB70q61Gn8dXnaM/Xl+ZkocP7aqZvyWi
BuQ36pIhELrPZje/1NGyb5bQvOhF5IGa19nVwRRxlTTkF1Qu1K9i1J7fuxPkfbttHvqUTSDvUeb2
6OEde0SL8ilIkv3DI83jzFw9GxM800UL9U5D+GTBoSZ+vU3WMCsfhi0F3yEHQaUazmSamJ+K6sq1
hJq9wpsxW9rWRJ2VI1LHbVRm8Z3O5jz0B/GvEUiAaEyPiMXkcmdyyF6VSetFWvxBwZXUvlf1PKkq
C21Nmmj7DDvNtxAjEWR5gKK1IgG3egpahAy1JD5Iw5OQ7UAWp0Rn21ezAI42y7zW0yogOZ9cEvuX
NbpQg2jtKTHinz93x4YX3up7iawk3ulxCcsrt4rkSiBivjh2vUVHRIQ0cT1A2M14twOz9KB4fb6p
/Wb5QbGTTB3SIifQ2NWQzl2/VSeRk0H3GPGIcvh8xAJEyNJAfprSSCbZJ1FGsIOSlwkaaY+4zzv6
Zf1A/TZnOTrDwl/fEjC+aV+QYU72LrJJK5jNOo8tm42CjnXNls5w8XWhbkUteBgSRt66GSJoLfXn
xNdjyKccN92dHhgpthDUxl8zp5jlZM4twZYpE0GS2+OCeVxDeFWS93rYyUfQnScLrPjtdTmCvCIl
HxvY/4F7pp2myYd01kdL8aiGm9ISjhneMCC0JusPOPDNIj6bTl63bYJzJmnizOEGK1hg4b195SUx
ifczirExISqBxlJXlSpOdaUBqW+de2kVOmtAw7aUyb3UvcTgETHo60WeN4eBahSrIUO6qA7ThFmh
kZ/P5onO+HFPyT3A4eTWZLOoHPHftx6/GC33dz7jiry4mWjTPtKZ+q6xk+rtuGyBRuPrFe0rE9TL
QhhfISmULfdlZrSxk5i3/WEK75pRfniPPcCYA/38tTRofpl/EH9ZUcpvBisASEzF9Fhc8EA1r9EJ
MLUG8V8SmyygCA9GVmUG+JrrzLaw8NUgnmBWbbFCWxh+uI+z9496T4v/ywh0bj8+peKYOXmNx3ay
jBF0vz4s9DaKY6jjNF/WJgeIWL5bPNtfbPx9CHMGCs3oIjxMEyp0TdSe4ti9wcQDIqMX+8E5nqWT
IpmOb9VuBEjwqVKkkapiQR4Z5/lUSvue3BYf2f7FksxLYgXoy/3WiCELTTRqpM5J2OyJiFtaFomJ
uSEdyfA/vPuoZCD6gpCAPnYLtY8b3Dmpze49MJjMqoHraHJPZgVMbflC/iqIrDGtShBP//0uSKA0
+zgsfJfRNdXNdI+Mw7UXgArm5TLrC7MeEnCwIB9xcWhuc4IQ/BFnVXA4rXRKzqJqm4cBjNb182u8
NE6dnV0nd/AE/5Pk4bS+WfPg6DdP8sFnwBBfkOl7O4n0vP70AW58xz0MDFC1UtZpaP/NxNbL6iPW
Tj81ks3vHfbeps+cTbydq7KlbHLqsjqODdNKC7u25pr8xuimF0z0lvcfIVgo2Dqm2uFHQQJrpnr5
evvMOoV3s1FGrFDEL5ImvHdih0hYP/O+jSF3+1yqUh6pZLYvx8/bM6pQX5lkCGykVZml6jqwj0Sw
rZuWH601KM49U1Ic9Uvu3SSsIo9Zk2QfkodC5vSWOFkRFwP4JFk16y5lumw+2fz7DsLzUNddXMMw
5+w4PG5RG7fQahCSwy2xmpbWVmfLLiFEpYawUI3k+SaeORXOFZfFzbzEE5kx6paIw8GslgNiLebc
gpms4irlV0nVqPLdLt12fDW3f+bJTkwOEhtCa8Hf57xS5GA9jEs9dPTjDAGwoqFuUMlNu1aDboje
m2dyH2KbsAHX8rVQVLlE+psTgHbtj87Pn6EuyGZUy/ixOj14Kb4KJ0Sd7rh5cOVg99M4f/h8HSzh
DV4KjPegeO2M91o88bia+YTeZpryfQHGwuL0NcB6pqP/nAURf7sTLPAL+mM/ZR4zCdcWK+ppEldX
iGKPNoMtXxHXH5GFo21Uln01H3gbRUMLHLStul2w01o3gycn2NE2b45hAGFdDQNCBjttzMzIuwWH
WPD+MX6Cox4AtWrNesyO5J+wX2it3WxTT+iGYsBpCEHRTHIlQDmaDftf3z2eCf1xk36di6Q8P7R5
BDcOL0w6ykc0JXklYsfgci4GWMJUT8hFrSslATKtXiL7FbdZVMqH/oGVE5iOUjpYr+wuT1Nbfk9d
08JhCxLe3vkoCpy0kl0Ld35AJjhHh7nqY4dvJmKHboSUgWUvLiXdn/Hl5bI34TkQNR/vuXnz7dOn
hIwrCc1wHy3qFvrKC0fTc+YxVKBM4bkmJVzOMuWkkcAPgZ9MEoNIcqwzA/gF93wVNphH2e3PzPwK
HWfGIJrn0f9d03RQggauNnh0/X3o4t1Yh5STvcX7OrlZBFCVek+CyXaBkExt95xvYY0RAPn6oO5o
NPaggtDlr/ZVu5q1Jk+f9awwBtJbDv6xg1js0c6sqOSJHdS5LfKYaLM6szbcSBd280QnB42Sqo0h
Xr8wgjPcdIjAc2x7nFeGG1X/P38C98M+qQmm4FsEmF6F/J6OHr8gl5DOFA+No9I1jVxZKRmbRIkd
YgpzKQ7cyDvW4ly1ltDWvL46nhjcJCyDN6DYoXZAX5s5hkvAQTB4J2QiD9o4ymXHAfEJtHViuSwh
wkfJS3uq5Df/zcTwz4hJYqtpaoFiZXm2/m7Po3jVRnPV47iOFHuEL82ZvVDIPNuiR33QVIYb2R4E
OUfHGHiMahSc/fNPgx0qhhtYobJl+zxbgOthfHbd9ArOTqonAHnE59zERIqmdVnD8XsTVah95KXK
AFf3j/IKNUdO2Q4hjTScTYoxirjCYi9VovJGVRlh3YKHyXfsVRp3DnZFc3pVs+sTI0LpSy1VL0AY
1NqXf+VSvA6sb6Dc0YTaLHlERD8shezCISU8+LrQKVv/0tQGEwHqOiSKzkc5XsQ9I7FePsuRvbKM
eLy1S3+ewHXAk0rGW/mdJUOvvlvhGHTlWJtC35L8mk/vWATcJWFKdsHyA4iBvjuqs/H/4hXiHi8U
DnGYRpMghKUFPHSwb6lJ1mvr/acBhfILzgoNAY7+ztqWfzy8pz935T8Ua7w6rlnvm/bl7bEh4hjj
65fnjzt3FBJgvdd27OdeUc46Y7yaJcsrINNk/8c/8wZycy5cXBabBSqrQVaDsrPIWYIeWBxcI3bz
+81fhv/K7zFJCA6dIB/odoxhPVPqfMp9pAe7tPKJGWgkLtSltx2UbjRdQAszyPtnwWDSU+IB9E8G
GNshFLoL00KiGA81NqAFIojaSQAI2wFmEV0V63GmeBCzWwODMU2B3Z6u8g2BmHbCHAYvjV/7kqdQ
glvS019YJRXs0qucksJ4IWYDIioQkBPd3oAfNsVXNqiKp6Ris+GjcglVeHAUI9FP54fPNE7zTidu
P7MrM6t4OcUhD4PFmYp6QDnA8ko7Yn4mvj6eHvvrhDRPCT7yLG7uXKBQHb8qsEoQXCgkVfaI5NiQ
VqgrpXtrYT8evrSvs0ywqNWBYO0WmvZYp5KkSKvhSzZ4/51cp4BfTJzgFEPSitzI31k7PJ4xYW8b
Y6D6HHvSkuY4LTHRmS4pTUn9DFT/ppYdKlpV/SZ/ESVx6gvUWR0FSUzJVHlLXcKqHrCqqLsQ59sF
Ib4oDiEmy4PCcmOmPqt3DQpLdXtGnG8Pdi1dP4tYZRuJ2RgWi93VDvQAYwTx+o8LORaw1ykISEIY
gJOhwSkEI4pJuSGxn78j5ItSJ7WenGtu0spYh6sKgTgX7t13fXSalZTellXrLn85QjGEMk6S+7TM
Otji+BOwqQdIwNGVURk2cEojrwqF4Drcq8CQAEf5x17P2y1nmniEVbQJpozn1OrlRKKd8gLjYxwy
Wzy//JxVA01bN+y4zEsTptXZ0xLjMirEHwpSZ1piR3N2V+PkQevYYHex3f1AbeSJMooK6XQ/trQx
8/2vvPq+DdfuftyeCluzUiNDH67f1VY7cOYlyYvf0eOoOTVkZymnVN3f55tXLShVGt3HFAJm/raz
evgYSj3C6opxnSUQ98t5UtaN/O2XAah1X+J73g7wDxrLmh6y4CQWBnvNapCMxupLYB2pDzN9Nw84
e947UyMNvispWaTfdj67AshXx12t4grrlOpcEoj6njWGo4uWyxSm+R93pPs5YWQo+C20hLyieK9W
j6+ym+1i8laadHKJohoNhkQZpl7iM8z2vByHiqy0Dw6TO6OcS63y+NKsRXc9uI+kxXdC5Xx8WMu8
VhRbON6VJ1oNZvtaI7RAYvwXQDpGU0Ww1sGZVqvhC0vpqEvLFUvFhoQOnvzQMtU9PXw+ant9dhaf
T61ERuThnI1se96EI8vqhGbaHv8M5ic0x/qSZdl9FSLesbokWhcj6H018lvc4xUW4SP2Sgoy/uhN
ah75mpqNK6VVTekD7T7MdeszxBogvYRP9fVlCGGE4qfoMNroAiZML1Xy6R3cPyYJ/cwY6o+oDguV
OgOqJEJiVTs73hTV331MQ5Iz839RrasFfWptgcD3OxHhlIHZxkq3wxVPCstrEaxv8n/E2Xftxkn7
sNzZYMtza8ZQIIhukJEPX7aQbt6yOxZTYsMy75NexIHtF6KTQ6hWSeBQWtCN8KjfMF3HmLGk0aOH
DnklMUWywPgMadpOl9/Ui82Yz4Q6DYXTnDMoQPKzvaYED7HdRw4rHKpS65NfuRAfjKRuuTzyp9lZ
KpGHCvT97CVL6y8hiioiTKsgCJyF4IqYnAKAGxaQNy/DgEPfvfd1EJbYmU9ANgu/Y/2xt1Sf0n7x
FxTprtpQxIOfBlRwP1/A+xBmYQRTp4mjrdh4L8+NZsam3tu4lv/2KUvhK8zuE+lc+xjMB1ZCmyCj
h3mvG+vXTsZ7IrEG1Xt0h31YDj4YjNiBIMIpCtPbioPfNeMyR2F/hssg6+xivC0rM5DfYxdcgCSB
RVW7bjbiG/WZSOvGfCbW7d+Lu+hD6m8mZ7GbHtid0d3P7yc7ZSMICAdpotB9R4YzqtZE0e/hjsDK
9qFaksEHgFIcGeK5Y9FdL2FZIx8Fj/YUXSw53LspNcKa4lQ/DmKEOlzHbJSFUX2lDOjcsFjTkqEG
Px0RSz5SCYdWUtz+8YvEuGsQMV/rihfzGxWCNXt4gjTHr1Np66LfHhBYh+0DX7PaJmUxsN3QZ+R/
IASsHsjZ8Ubr1F3o0SfI81PPmgJmqaY4IJWnGi6wszM+45Vu90240Q/mL2PqFphWRlxz4eCWD51L
y6Vld3VzrKmM0ig4a7goAf749PNyEMXW+1aEk5wK1tL1gtzS2UETPkaeEAVPsHWzwyUmrxp/Iz/4
qLcwPgia+oGh4k8cAPrMTuUp8Dl99tRC/eF/gBc9fsF3jZ5lNKoNK6NVEJKrf9yhT5vrnzCpTTdT
+7ztgcHJdHlJnf2rsmVCO61mGnn7v/TMx4x5P+riOL1mkFaGzCF6gGToIQFmUgZc7t5LHJ6zJeLh
JnTuF0iKvrw6nA24ByW1DQddAhT1Cyd+GQgkfXxbIK+uDOFb1Rr/L3gEDKkhIXpatPxt4DQVybs4
iNP7LFWootrB29CLglO1hyp5CMeTXjiCXa8/Z4J0ky9/jm1Uf8wZsWFTyE+HAaZE7ykNknOiCHWK
1aWVSfyPzcOFbBVXukzoX+s9uuBd0xfdKXPfWhzGKnEchLtb8caoiM8kkuOUgdEzSHraGs55/F4C
bVN1O80YGdBltvCbbHc7L/xZ46O/6SOohd4lI6ge/fOc9nxnPLE5cONPnRGTgVSpid6inyx+dUP3
9Hsk5Tqeuq5Z1rO5Xti+oRwVU7RMF7fUsh9S6CYEMzMQ6+Tr3apZ7sRKGtrxyozcuoBN5bFzAjGU
erdQALQSq/11XQTE+F9qAn10COJZz8m9jjZhuXk1Kq7NsM0HN4JSUfSWci5PZddHqCMO1hzA7rDp
IG56oyjyRwMHVGqQFSldsclsFYwoxKDOJd2+L40W1O/lGmIb34oTLmtxXLPt1OjSmIg3g8ADHsxc
QV1rLh11pnkvzRjhSUlW9njzjnsMFjLJnOrkmgrL0OCC6CEQ7o2FbvoWGjs0zEgKT+QfeiyV+idx
bAm9czr/YwXQPluXVUNcSDtPDk2PPf7APHxC52w22mgx1BmBgZ3LhGUKgwVMsZSISGdFWTs9IWrl
uEZ9/jiM2ssg3rQ3tqODgMnWKy0NraiO0awhv62F+xjzGf4q0trTFUuYu9Kq2vst5SWY1AfSAiZF
Vc3o07KE3KbOxTj5lkYTANSv518oDaPq7ZAEdVKCrHdtU6Kue5mfXwbLnAC/5+jBjdUUaLzhfjXP
D33/ulNL4u0ZfEtC61OwTMIKt3OGtsn8tMylR3j/O0+yLu2INMHX8SonSDfuOmetsykTMtHw4g72
KDtsV7hPfESlglehmvdjHXfhEzpUckh63oVWoxQxgx2iU0YARZ5i78ab7PJbZ+WzkGOZ4XELVUe/
rwzFcOF+5uBRZ8b0igNII6LxLiu2vdzqZyk5pB8W+t7PtGWZgcDaI7ckOGfpd9pCyWA/uv3bWL/g
obsB4TzJlYcjdqY3QJ9BnLCDpvirE3BsaoSlntSMx3Sw2pcyQf3GbaLbGopeX8VANTWWAPnQW1z7
elShWBUXht444NWieNveFxA+Vr2O9bSpqCKWv5jxSVL6OJcWjHHGk7d+nDVO07PTaKSri6HtIF0j
0v7hKM+IFB8hiRS8DvuHkNmJeR4XfJ1oAEDk1R5oaIAW1ZUxuUsilwbce6vR0SokugXn05OFlKSr
cOmFK0gd9FPcijRP8/R8Iw92gNqIE4OU8EWUpERW0BS5+G+WTMtML/MJP1XB6f1URLAk5DUOdVnL
riZZUsBvKG3ZAroSC/Ea8bHLYuFsjFiT1etYaTyHw2HnlZgrJ3BwE/6cgi1XDAfBtQcFRlIx3Jw/
Zna6yGhZHEu2DZ9JXAc2uXXnoYHeCW9c6K+iSu+o7+zOJQq26Pq6Scc3Ovsux0NBlYxAXaOwX/qB
pHOtFgiTx/MDPASvxPbX2fqReIthI7LEGezKUdwdFGwa58S+lkxKEx7ZFF9K1zD/xmemGnVnyWQV
pmtSnVoAechxUezrxwJFmHBW1N2/LQdE8RubbjxTsmjPhAIjtT3Tk8lkNNHoAYJdzg6yeVStpA/9
7ifG5Y5y0+IBKm5hYmDR1olNfemIJe2G3RgDytXAF8wFqPUG6UhI9wGHuHa9/Vr/H7cqbDB6+bw5
dFIaDiYSozTAUwweFznvFduryV7c7Sr3Rhy0BccmzYnOBVSp91sljLkfvmFM4A4DrbdtB4lYegef
Hk6TlYt7fE/6ZGHdotuR0CoUGOhBAhOnu0wcxJfHdRXRYhxA58NVCNdug2k2JC8ORnJGAeInYWyK
pVhIcuOPnG19zWLyxE5AgprxQSpouDoob4cJdHFTqLh7BLSya6pSugOLVzlLVCCpz4UT0Rt+iSpW
qBjJZx6WnFgQypWZID0nE53kQBavYpnYfRfTC1TUb1xtCMJNsvZHyL+q5Wnk+D89vwuUC3Rt4k8O
rT0X0nRMhILpuvrQB0IoD7fus97Aofp9+rb3QuTMMzLlW8L0CFz3z8N/wZeOg1q7HW7pkD4oUf09
XKjhnYbCR9A54n3Awb42SjRBlM/4Te8nnPV2t0kBy9dPvoROsyFiIsB+gaxni5kke5n0RX/7q2Xm
wKTAuVqlwxYIlSO40JiPUTUgQ1u9/c4zaltgLqV9XjROHuv6m0HZwjNviIy6srms3Dws3UP/GHzO
5JOOyEe9rGN8quFRGJLTunYjPiaLFrdxrwdEmsuCEKhJqH3X73zmzJj6kL72yvichu8oHDbKBWZf
iU7ORwFbzVkv5YPz5Wf692RWuVL9HahUBm7lHyW/Hcel/XAon2McfRYS5KLx4Fm66oVQru7Xw8mS
EuqRwurtN2XtIMFSZdEIWN+7Mwk0qwVs+ieWNIvdbYd6nufTFCA8rOyQQXsAOutH+UkT9jMlO6sH
hc0D3+l2lHX8Ic5vkJv6rAr8SwazxX7QckI9KDH/lUXXvnQPfnxAdH+F/Aw0w3c/zWmdmhvI4kex
ML/b+VW6fcc9tMeN8xOqMzBLIMcZdLygUQz8/sONF/t0BdMXvWf//aYOUKqU7s2L43stHfQIi3X0
PwIirN8uPcP6adNX1nMEZpPB34MQmEhoyUVJPv+fPWnUoOboSK3UPpMwchuIG7vaS+Oz0rDJ7YrB
6ElhJnkqPLmV/Ou+FXMEkIb4M7DJ95dTBW9RSbRct5QwooXA4m6saSgjQTD5AJX3P0i8i0EaW3TW
TxRIbrCeT0153P+XZJLfwJXj6OAKYORxcfxc+LSLSK0QsPbtqyrXKuvB6VzyPaJFXpWLPuHPLrUN
dek4XlQIL8j9LZIUDEZ7yAODwHO6DJsg4VUaBuJrrYc89ZfmBvc7bDmLMMrB4PZrKEW2FQqlZaM+
gZVkf755nMYhXIDeEU06W0je6CvTMCR0D2uC7lkTcehxMJ6okMJet43NIw/R7IUjtSLl/32xKj40
ezDuc65rEZzrxeXx4rirv7vL4iKr1n9CsVY9a1cl34lmpsswyJM/VqkwniRdTlz/ZbOj+165K/xb
MZUT59BdmEpEw0T1Rl+R2TNO4J2D+/AhT3HJOluhuC82S3g5N0yzWFmRcNXhqayzK6veHGYHse3t
+9qbecxB6Tb58ozt1vQoXQzd2LHyB7ZwU4vDMzSfjtibbnd0oULQxHMQchEAruQqgygL0RSKZuEn
8GyHSZkhAeUXLrCFd58TDVdfRUK3vC0D8irVd1N8zr1J5BJIyDE06cZIJ4WtMLumqJMrWU8WhSqA
8Ij6ehvY6P9dL3vwZfSQBwxcMWSj/IkeG2Jx212LEkbT840FXDzZjwWTRl+CPNisG9uT0dlFz6tG
+Fvk0iY86F0+gHNfTepFgnUCnYQVRDC/PU+U/xZS2DRThyUQuU9WdRM3uEN2icp/SXJDKD76Un6M
4D84BrdMXGxT10d1CwLklDO0E+Pqez2gtCszN1tzUYRkYBe9kVeKCkKmlR6d981cdXcjJF03DFzJ
qCTTgvPlofjLu3lKbfx4aFCJYVKZ2WjdEycq/W71LrZNfpFT+ek51sGZC4cvJYy73KCKe6nAAdvg
zMBNSZ6bsD6NmsqXbvwzR9wq9oquN1nJJizF+jEq5HsBtjYC4h+jk6TE42bCwX9BygOqNjtt83YE
BSikNVrmbhsEwMXVNqp49mLrAuoMiGee5sYcw6F48jVzyydupydSXQGrEJvk4bpxS+KXCWCfgFW3
6c1Nr2dej7T6Ks02mX6U3z647ocie79Lhvq9MgVZQ6SF3WH3Dfm1R2Uy3aPKmWNa39MGKmdd4EM3
+WbxGaTQN0hix3hlqxSO+wGAH19Mwqrfb5QRoWw1TOrtGg9sBg81t2P8uUJIzoklk++HJdTd7hdi
dfsaiF6/sthBVS1tVwxxqSEp5gRfXqw+4f7lhei7rxb2F/Pq+EMNJSVBTUv9Q4KFfeQyWju/nk0R
mh+IUlXRkdcxamnH9vw/Y2ac32JM89AcQwbTYP+837st7ZRJ5xonWV6Mu4gRnwPk06cVP0MyCOAP
ayTtEzLj2P2brXzXhBOocr4ifXRTGdlI2LKG/xDU0xGo6IGd8QhlADy+CKkRSI1LoNEAxUpl8Nrl
1c07ID4NZEySDVKUil549NXfuca4nzAV2TCwWH2/N3c0Lq1VvEXCKSA6vNW9Lz6uTDrGBkmjERlS
foEQ6gw1H0Js6NtmZaPH5O67tTNCclyR+sC3vkc07kv4YHNtUQUF/zfmUr+g1qbMyilK8UiZZnhx
boCxSY5SS1TZQuiC+Zkq/CShKJ8ZKlc4seEhOV82gfUIyv+eKkoaL3I+0ImROSL1OFdZHiqUB+ey
Nzw9vdiV1TX/k4a1NT+KRcqeP/r2HKYaDDeQr9aGRcuNtax81hfiYObOQHp1CsHrmPRwrIiYHUcs
bv/yMWHv+NCwHuE7LKL0DXR/3xXMgQ43Wd312reOO1aALHjKUxqJulgYK/Lo+ojogce4PoeOvidD
y+Bhrf4zudigdIcxHHsqPqeuM/OgNQZTiA5hKWAkkff3JNqK3RWeAzpyNgKlw1BPhCAqqkhRQW2F
1aAX8eEvUioREAh8cMn6sTgoPlLr0Geia7jQQFzf9SKJz5XuoX09LAL6fE2TUow2q60DCi9pfeLK
nVwAQsF1/9Q+pNsoI6pMLtZ04HEMEHnbyKHbJCcgeOydgeNZmhUyAaIJQ30dzJvekmPYfBFRu0K7
6GB2DPwIZk1cw28vT8klfZkSfpho6XDtciKhVnaZL2nv6N3y3WqjtuTGPoqGhTOD6BeCj4x7L0NT
Zxjx8t10sSnS6XqPQho1JVwKc4Ox4Ju8xy05GGLVSIIwmw+oicF5Y4t1SrK9SaNwgDEhBGVZ/4p2
/RsEhtBiuB0KF+INwJ4ypwwW9/mpkHroaVU/NARjuKvK+FZWA33vzwyMx0pODWvQ2+bwEN9PFV/x
OIhyPOrPf8Tn63UHdQFaO317IdLcbkNzCIppJxaSAYzp3fYlx+C8rXNszGyho0vVC4cxmtslsUQD
3Fn6BEzxMcG8oHZqAbDLI9panczgYJKF2491rc8SzrWTnVwMf3+tdblfQgemMC0OAEjTkISIKxa0
vkIt0a0Atw+1426xsqtqnWdP3b7AGdsB1FzQmkomsKjp/1uAo3t2auqHHs2UNDOLsvV2XLhEZdRZ
i+rWklxTM1SE9eHnfLfEKsmluWPSqmUYQd8zb1LfCzafdgS1yrddWV95zDOGaEbEYtJAtsICKkLD
nFB6mMUm+F/Eiw/4R4v9DwnLiIOihkWAl5fqO71dWqxZ3uv203pcKbDexvIRm29kkCSL3smxqcrJ
42dm8YE81Lla87nYQmCxk8ewzrMeNRMaYPLkjYaZkuGj3YS+W+1As7uo3aA2AcVqzVgYgpsqaCkI
KyVvepL8h2ZoztLAqGDnltXZL71ZXAHNEVnCkDBt2sTQCLkWg51RxTYM2FJFzfjkIs5mbunbnD4K
aqGlD6bZejjDDKuAS8p4MduXe4oFbwyLqCYMLhA1C/hk+uIhw4ICpds7AAMBIRzuBPexPtVJl20O
lnc80ujCEiLe6v/fIBqhxroW994O5RnIN4kljvMYZoGODmUljVuWYy18PiPVwBzVVMMbnToJ4Jfb
dNE55nL0WSVJdk4dR+v2GyqKTAizPOgrpu+cqz3ZUtS/21ToulnHmJ9pVhB/O/J36SxDClTHw8Ws
29nxcXDZGM1ZK8+1K63I0sh/OFZnrM1pNjsz5sG21VDV7axpu/ATx9CyjeGKeMVXLeoPVk9mB1xF
AMHznzg7mEBTthqPvVQAW1UgCMnZPGSna64HaYaGRnyZudcTTY6vbcnRwP56nNTBMPX8QbNdbRHb
TJby6Xb8mCC/2+MgAnM9h7o7uXULzu+ANSbx0HkEbA1a8KrnaHK6N1S4RTDLbJkxDyPoGUAxZktj
1ZGHoCpCB5KDXMBGQqUDOPFAKKMIuDeHVzFhxsRYH6BWyK+uRbHxh4NZTclb5cpqb5uOn5G4vjJL
wJABP355qAOARusWGerhcvXjzMYQZBYAK5lRa+6Q26qTkEU6nrOBQ+gMrAXSu+i1upBWbJZLuyb/
qOjK0fNsuKFUEXjH8tJda9kMnmlKRD1Syn2itYIPNTG+Sk0QmJyPHgVDA2xP/Mf0WFGYjYpp4AW1
BLPQa2n/CZi1ylsq0Xg4JsWtJUk0LTBVRR0qZfKQE0dYu/JzWmB4cgiQY1vH+NzegawTL8TyEHRQ
Z/jYTFsi7dZVub+aM9D+MXOsfSTgpf6FgvQVm+hHIpIWltXrkK8YdeSJfmKUniDTX7KnDFNkB+ks
7QubrSMaBWzVTgpT3FK0wlrge3Idn2YgkWGq0Jq8DnQMkmJlnGXU20zFCMyDVyqzJvAix1snEFeG
BlHr5VVJGQDBHb7cA8PWPl+Ozt2SHIPozHTrXjWweExV2BXhFRAoM0yY3QUbpqLme5Rjbm1qKDgZ
UBn7gqQE0IZtvxDZm9IG9VdjI7x/vB0l3PyNaWsP0TK1us9/ix93O5HYaFlT7wtn9dcRGbsZXJC3
L9uzSqGgCC1+xpfyOQmyWHF+8sYDRPphcoVauWVTAiCVUAblf1XRaSZ3UGP5SQUEzW59PMe+8QpQ
x41VmrMb69ay5xClZY8ZyksLsaHbmXca9XS4yevoSEnAgZy6fIQudDujDrTmbrSdS/cDOJVLs1qe
kVB+1OQlY0QGwSP7C9NoFiAZpRU1lT8pC8RK5BbygNo2z4qddo/iFLEtceMrtazb1sWx76XXeGJM
/thuMuPc7jO1HCkTYxrKOAaCIqyN2bgRk5s/h7v803KXAVAyuOCEJGt6RdLVDSw7DCm3yvYkZi4N
f1sCfW1coy2Q122HfIPjwwWwnM+wOvohXkrFNnpqgaCu4Ihz0C2/MbwcODKasP43isuq7FzIC8zE
ZW89PMZ1KAbjLN7y5q13W4RSqXGw0/UhgJeUsdT2Rnm7u6p9qM662u6W/Rw4W61A92cSZf2730lm
FgAlVHTpEqXrhikdUhXEmP1vh3Z5wNR5G53dW1wPVr6fb9vQQ2U3ZcxO+MqaH0khN5s4ps5FFM0D
gmxgaYPOnrYp1MXuQCM1qCrdGt3OcurRd3MqFoLoy3ukdYejoOrxdlT+qsTZyN9WzCxYGCujJVyh
/T6LCr/rxPRseaoi5E0wp9xnRsx0Z7u9epPEtHBCOcS6tEfDXgmMGHZegZWlnwuI99Ba9RSCUCJx
Im1VwKuzXmu7nN8uKDV2LB4i8sJ0uT71OJklqpk4CXewYWmuwXqahw63YLAS5FlYGl8i+/VvdrwS
5Nw27du+CKwL0LfQ8FwUpT71kofYLWPLI7bPZ+dTlHP1h/9+H6A0h0q9jpi2R4gJo21Oh81jrTdV
+V5VkUaaaTNFbzpc2Dvjo180RPueXxGpL31xkXvIciFORpxGYoY+hHEC4cNNFmlZGcRAMP371sKl
c/8m2+WOA1hse1haEwv9jjpy1DSowPVsV/fbkk8eEhkZKj+n0N1jrBxFdk1LKMyG6iNad/WDGXRd
qo+2RMcPyXM5igbEihU4/j9psvaO8ziujnb35vIuZXNojjI9DMKE86NdWIdEwYcL/7UqmCDaDGqc
uiBAZHWlpGXpOxHk22j4t+xhebkKUkH8f4gz6SWeqhY3gQdCu2eYWgft8pCx6+Lg0uHvTQyiXTgF
FFkyEDIGxAm6HqpryzjPzPV+19jWXNSE+EWkPUF2+wW1EbLNTIzPqCBp81/qc9al2uOfJ3F3Mo1y
blBqDSudKqTqbNSFmsghMPqpwCtGgKRTvDiQ7zsywDtoONM8/SMYMV/5s880UEaS2AVAkSp/RnfE
QYWPYvjDALmOxSRBEs/RS8VYPF5/RLqG2YyG1wxjqDrgojYXDDKQZ1cJvc/BbSeWStW0dJ8oOfNy
Fh6Lt2uXED3RgdHfj4VwrcywBCmHRnBCC77btTJOvFL0N8VD//B2JsIL5ibER6dvazH1DaN1MNk/
eBdAMJnPatuuZUUH5+roiDCx6WM6LZKLUnRnctkogsvs29/kYvSZtXDlQDGxA11jZfJGTqmW9mXo
CTiunRGYyCGa4HmGJfb5mNOETNi4AsEZ1Z+FMOx4hIrRCOxYXLqG9VoodXBjGyEW/kXnt6N0zqIV
xQMP4LyOIu/gKeSqeuJe0o2QqPIT5KIzRjeKG5lnzQTI4+mvgmjEvHtpQz9yVzZW3b4tF0A+opzn
5CivhdZu9fi91u+7YBMjGTPplaNF9RDyG4Bn2J0jPYgVIIaEl59JRUU2Hgip4xvzwOzcVjvLbz9o
TLbDl6jezXOppot1OvagLwpz3vEpqP5sFeP/BMNzjJj+n0JNZfi1+r7INoavQ6SCz+3ivFRa+BXb
9j8Mr17Y2cIRvGwAx9gMhs7NWo2gH+jwqWd5jmWDnm3XnTUcphZQo3mmjhnNhURX1+fHERZ0yYeK
gaBWAO9m0ZYC4toRx6wcfVsStb/+aso1Sd30mlLfs8d7S88o3ptrZ8ZWiwwX7PO5KuCg8XAoDkrl
JbHGG0HToxj45GzJ3J2KZEUYFnhJAcLGEREtX9uVCdQ4F3zLTSzLLRcQtNmIb/BedzMRRcp/DwLt
rqV72OqXOQO7AMI6kf7+/QBqRKnl7UfnyVuXaEfUYqZ5djs8rm4PsxLEelijxUahPo8thdaVTVNp
bpHCcBozfnY5gSe1s1LhqTVEZbZP83Q7B/cQ6UFQQZzWvN+CN3rtYCtAVyjtbz4N0z0IB26oF22k
JgH/I74a6xnQXNR72Y5CzEg0pUEm/lnLc2ehUtVkytEfjWbu8dcAL3TmeGt2gWdFgw1znxv5SbkT
DacnH8S03qMk5BT3FH36xlKMr4MFExMKWjghlLY55wjsC84MoWYIQGjunz6ssp1E8X7W1QNDdJC2
jjsEhnT4USYM2Q6AwOodHUVcU3vA/ZherzURmWwGQfdfoHUei7Xc/26M+Gzi1eLtEXKIgnqqt9ju
xJIF5LwYY9hdCMn8vYbs6C4yONFjG1ix+Q0LVHMWVszJcNpfu4tbgNH7wTCRkhM6W/OJBa5VONhN
LG6SdTXr3bj8/Q+169l3NJGGvxQiYqbJNWG2JUqfkRncBsueJRazBlYxh30fjSGR9eXTzGgihhta
kS3+/kdcZyQHHYD8x7yaUzfYMAOzX6VccqDGvt7yivIhuxBJj4O7PQm8PTS/vrtMXiyHjzObTdf3
8bAivOMvlexjZW5Lc7snI4wo0wLynLGhW09OO0CQXGN5xYyqxzOBWzafqsgoWv29fSgbE4Z9jvwz
63YARARLEXU5D2mEX5sJOZ7hp5pfZDvxMa/ndjA8JubdM6142OOBVoy+RBbb4bnRxjn1YoB/yt/t
0lIklOlAc6D/ZOiA3PhVJNI5tjzu7uOE8J8QHjVY0++3Zvkj0u9RtmROO16EaqbJiySCY+Op4KTX
cuaQLVWvLg4pguPNp4955qgYKlD2sBNX4NBWvl4NIkY53y1juVmUf9jlIbziLznuEhgXnFZu1Iaz
nsNul+mq+5B9hf3u+WYetSLauZ/KjysaxAyDiKVNtpo/ydisKq6Cyrj0zAzC0BUY28ddrG4RCttc
xx2pmavGiU1EDs8uD4u2XIeKSwXDPylkhAf347W/Nkrzu5INUZwv7WSTKeSLTlCkw3X2SZjmHuhl
L9gk5IgncylnSLLpIz6OSI8fotJ7FNoa4tPoW+7LBJ1CVWUtfMhmrq7vFgVo28rm8130keZsih6D
Zjz4hcsLEndhbT3MCQNJpjZzVPuosFfhs6QBMXGmjXNPYtcI6kUVDf5WZO0Nho+D794Ikl1uQjbj
E4y5Qdnt7B0vfvJsWRSwGi1rB1qIZd/Ss2vnG58prAqk0bAfmsRsDM+e5fOUGyxLSfavTmRMIuYy
kkLqd0mLwmYiciY0gTEJ0vReGWzDBsvoYEXZy0wEnmhJb9Wn9PIFZ78aRFdOJcqYyimQjqaxDPIn
4JzTVbmw2hpZXeSYq2StHKLaruWbzsPLfdMKDGEYrQDqQdRPPURdUumCl8AGgYlN3/g72bp81QnF
534SnVnKshzph/fI8LClBE8oJQwfmTiji7uYzQpJ5t1itLD94YEqDo+5SOKZ/io4B+ngrrJqIl47
65Bnd+L18N4ojWcc9QmzQjFZlg5Kqgge3uM2YI501gjV++rcgLY1Le2Nl2uyUu9TZnYfSmNttjTC
n6cLYXb/HKQjUCIPq4VlkeHcNjxRVg9KKF7k2F2DHvZZ+86mRGqGo2qnwI76SPaJFuVuEZNU9WgL
UmFuiiVkpj8Q4jEa3CS0rbCe8t10RrYCkAv0NB0Ul8rYhzKwAakotOWKdpby4XJMKBSxzvQezrtK
9I6SF3g8/4ksBglDUNX2NYISa/TGlLxUdwBrN9j2zUqyO9ckbtoIw8duzF0NNSEKORfdgEhpzkpa
AM8Lby+EvMnnMnVZH94KkfQLx6kru1B5rWyHFuY7/6nNenrJ4PnB4EN2aruexiPNOXDvoc8YbFSV
nQ2bxNxYE70lvnaLfuKbMbXfP9wzmRftvK5dd/ruJb5PhtwK5aka19orQZZz6+8y3YXzxwwqPfPW
s1LwTY77s52ehwxLwUETTAZgHevTD9EV2Es8SBWu1/BpqhjMHeGyqZVQhR5eT48SdbYVJTgrB86o
Ka+QIYY/SBj6hz8okMowhEx3+GaVBfzzEPSK2Ew+X/92uLWLyZTVQRTf1RI7+A3Z3JEeQzQobt7p
a0pLZSjt7b6LKkFvVIAebnYJYo+1VWYjmGnrCVDkxrfJjyB0M+USoim4T5W58EU6RZV4LQBGa1ap
uVM+Lv0eH2uoFj3qlplSlg64OxC/lpvLjmNqQbC4TjRlTh1+3zcfttGC7hGPiI28QCAPSPyBKCc3
NhwNLVv9mx8jeVru/YIyVGo+dIikGZjzVsOSY+JOs2i7A62mXVLF34E6AcmgpDma+YnOhky/jTDT
XdGUytKZhMr/NgRAY/T5PlDXIE9H2Wq6KzsBsGnXW6ly35eCQDJV8cZXJ7v7pw/UEiGiUtHSYuRJ
seNqlaR6fDElouyBl0GxIYoUtX/rrn7V0v9HmeyNxsjVoX47dzzI6hvgaVfHvmzpHFWvUd7+UG3v
IZ+0TeZfRfxFLO+t+Nneagy+IRsYVO3bBYG/sai7LgRra1OckI//nr7VUhrqVyVSMq/E4BXz9m+7
P7rRbJPgsRYN/ujo8rlSuqpVAniruQK7+QxLwroialkQWG3qSDymS6CgH474Jof8pQP5Q346oiwY
1c5n0ei8ai/ga8EXvQSFU3csJhSgDwSiEgIAAkvKDJDLRsZtpsALkDpnz/8aZ3nTjd8Se4HALo3X
NjH+tDSqy0XHea7BlUtduSmC7OEpVMEbktGH/1ZljbTG0qyBtEnZ/uJJLPnMSLvc9FOK+6KxQk5i
ohuimo+ozEl6gQKVMk4d9ABgS+U1Ccql3wXeXuPbOVgXvk14sd1TOWMo7MOa9RBSlnJyEEFeDg6D
qSWtHeV2BC34DmZ2bbMsR8rhdaMM2wUpRLw2HZcz1/AVt4SoQEpxu5kxhN4MlMy1qCiIzgbTSFTE
AcA61xaY6D0tF6Dat6xcDyjj5i5X9dOTDrN79ydnemsQUIOxls65Hs9ypfe42tR6wPn/xATzxHki
AelcgHkOEKB6m9cccUickfhe2q14gV8BwtLXPXhqD4KwTktrgzVB9QkVFXeIbJMBYWmeSxIj9SZ/
Eek7KK01RiuMN2H+c6Fhek9oXwXHscar4g/VwaFFRifIe3U9I0zhSuasjvSYUsNcUhwPqjJzDzVL
HrGgzgi51Oz8G/7sxwXtIMNJjT4lnA7gQe13283ixtHumQTd/k9CY9pN/jE+jlhhgBa6cPUegmQX
WHzMLSUocTQ0PCNBPhHlIE1UFN7Jp2glitrs9v4hkxi3ROwGgPy1DTRFYfL2DcU4Ml+uWIhJoXoq
8ZviX2e3hjt4hG/m8cJlvGWaZti1Q5jDUusprci5pgc1ppPItPv0TBB8FNlCg1/VIfS5cCffBkp7
6w1Fl29YnkLoWoMs/Oj4s1NjjWJMEJYJlRgbKqRwRNre1eVPGgnMFGlPHnNTAxFaF3pMTg5oI2b4
2qqdLwQsJcrrCPjHXuPYJzqpSnDhSspp2QiXLTIxbIjywsBFD79ENIjYBS9nkWkFST+lBq0Xma81
RRboVOUfapKxbR6TFbZh67lAAk9Or6tGFlg8XVVT+jJkJsy0VtCRx8irSbpCp4Vm1CosIEKqAKw0
fh5cOssdgFbQ1v73HfahVKPhhhbaJclUmFR4Y8/JUg77LaiNlkCcBC2eTszx7FDERn6fU4UdnSAc
bgu/rDNEnXZmTJge7xULGWZ6Nc76ft1KK25gTqor9UQgGHo9rW5NMjFrsv21gxgFZ5uRlLPHqQN6
W+Zz+iov2vHJLqNv9+bVli3UdSDf9BCxw2V9z735/2lM3YgNAME6KpOaTkMDFUYuoWVd3ROTQ/SH
W3R3etz7Zg4AIc/3GLv7dRFRshZk8I8zPedMctkoUkn/CLP6zjWTmAbk4EuCMfDijkzBZqxT7hMi
0WcXRj8wTW3k3S8/puLZ42ucNsNa10wuj3VP1X0p2dGV/tM1PqBhqfdpLCRVqlPiT35yhQatRY4f
dkZbENaNsCidfcfbmPrO8VMJtZIVMpq62Gsu0Ob+nGb8j02kJQNzUKV3GZtPE9owhuwHHwIHFkMN
zVcckXB+jN2jckUpMG586464y1U3kk8QUMSHPVZFmxnZfLVCXqodQe8dwFLPErOsrKRV/GmC26rW
hQ0Zvsf+r6RmdT74BxPZ3JavmacSD+YLtiL8+aWbAv4ZSEtlifwkY6M9Q2TalHJwu0IKqnp/k/f6
zrBowSvG0TwgWjSsZjsfVDaYvSAqPvfJTN1FYC2J6DywUZR+9BzRKs6RFmLsNm1lObc8iwAybaPH
P+ZBxZQ5vHQ1vYweneVcnAi7mFZSpgPd8JdHaEwJFWa7mGBznpo2ALZP/eWWZRIeJCae2zXPL7eC
QJiaz2ZupitcHmmfqCfJ5xKDu4wdI4f53VLn5Zp7ThMPb+8L7gOfJ1MGmw7VpBtwYcJ5n+kcaLpJ
1B/5U3yXyaEOe3TUo4/7s+ZBbMUkinPXK6GhB/JdI0eDV7mUr3OFztF0tzvc4xnSjEnAZM4kwCQo
zo8tUSIXHsZ7h3PXtSGkExW6animaah1oQtYylmxx1LRFKrymDwCuWcKQcIUQqF1Jt4tFPonbfrx
ef5VPqirBX/dn1ySFk8P+yJzo9u/V6GhEaz9SetmEDrIvqVk6v4zmTrynKp0tVvmrPvnooPnbrme
sAzarvDHk9kw/RAUoS4ysg5fIdilptwUFsfqKz9NjNQRuDnL0Sict0OY8DNDOU3J9nFAijCQ4Cdx
r8EvKRitz4K368OtX4Ya5786GKfsXGQfLS5CGnIcRbzN9tIOiny2nWUqFM47MivHQf9SErNLnPAm
/cHmlDDM/f8jKDh4IPMiNnJmBpURoVZAXSkTVQlDZXtCfKiUfxIUwodWzTVO3772fOua2HcHVNf7
9zS9nEgNiiTiRTk6ABD11R9ScB/7kDO4GFDhl2RlOujhnxL/RbjApSBsSojJnMjgX5NJpsdiYu4f
rSkb42jkKE85egxSm/K+RJOvWCO0a3LdurpnBjB7mrCDFF0sEDwoE23zUA5WrmbMDYLtfMkLCbMy
NHxk+waXO0U5JZz57d9LJiUcXsq+TDJqngSZuoMmoPWTxKruvzeUoyihfD5L5sM2SS5nlJtQhIVs
yF8jFjXwsFrTEFLdUuRDSMbH5sGcSelDmg3nKj2otFWx7Q6Nqnl8gaCyAxTiV3K4OLz97DYHt6QK
uPDgFr5AizCeUeOZhgES8ZXok7Q/y5cipRTSK8pTeCU08C3B8qGGGV/oSo3q4U51LNnFw2YCop8d
qehUqY27vbaDj9fpRCmMOOc+QVJeYDF67ZvyOsdgbOsKs2dOr7nl0Caq1I1nWJbzqw5JDjiXycBQ
zNfCNOcsUpNVAizk8ED6ICPYI0dYgSkihIKgm1ryNXu/V2N89JWdLmgmXTNB+iSZvqphoRtfSGQM
HhkzKLB+M9Wwn3ocLy8ieQsFxKmW0xWGSbsda/EvLkRLLcteX2frrmurfEHktpCrp5NZkOEHhKz+
My6vt0kptrhAVwOgBIesh0loa4JRHhTW1xI0WUG78dloFV3pdgpzaLyeXJm4MQKXFSdJtkcj7ZlQ
Kf7wyrzDe2nkrm8VN3R9eakcKq+1/OXFCVG506BQf0V1O0UavWEqSVuquyRxE4n8YuG9XYfzCrOW
SJc/eicWXrns5m1WWrBqmovhkC/AVW1Rle8EqHQ/RJBjn6Sn731c9nmWmQ4ofvYcV/wMRkhooupf
dFhIek/H4RewDrKfedfhBIZZnrJOeSOUYsJXtsNOjvyGWIJBfrhrZuCnVbvNvTlfamAs6rymmgh7
ZjpEz6z+0EVGalQEAtYyhmXsV1hYID66aAebZBPJOT479XEeXRS0ooWmgg39Jj7OU9kJCybH9nc0
GHb+5nEdlrlSAY4Ev2pNg+br3b8zUtsh5UVC6r37bj4imjL3J97f1L7zfhWFUMA1qgLmXvv+1baE
eWSz7wOfoxV7fiUlfjrsVb/VZtYqZkZmz2A8Y4VH32XQvNlmMhXD0FZRV/sLFhmD0IkEwnCpQAPY
E7kXjw/OMERABxUoysaPzaxEeCy9/KAJCN75aZirtomxu5cBDdK5UhDbNMHVYgcaXY6+H0WHokS/
hSyy7ulx6cjJF+cZHrbtevMZNcoDua9jr4CXKy2jDMFC4EGkEaQXyixBS8k+bCeXNAePLwsUx5au
yCGn5BvugDFcUvktpG7eTxsa5KvzpHIZq3S1dikMgqwmMja9u+jc139aaNNYCKKTnDDPvmjaRtCu
MtO9a0S1m2kK9cVyvLNPdvyIHYhyUlxM515lK1yTxdYveCDB7vkC4aAcgNLRNvDDWJD6WZZ0qsix
lZOy4+NFzYRJnAB1iHubjbbmN5pdyefNF1wVPmpjI/BNhlsA1LWbrfIRTcHAiOyhx1fmQjb2aTwc
ioaYeX9W5uivJBbnmUez6dl+eZS3njcW41UyyiMS3QhG+HqrMucsANd5WyIRhJtB9O5d30lbIacK
gpckdqjQYxYjTQpJvaSmHpDFQ3Y+FmYN51tRQJ2ozGys74SDY7h0EeD3KC+zmXj7WzMptnRRl8WM
z4MzmIf5ubEiP2KfNF2QsCkn/KJrhTx91poPj2Vtc4rPbqqB2u31Ll2PXpnea+sMkuGJTnteObor
AIpOgVIyxd5KeX5PR7Z6MTThM4OODIdexINDXudHkbPfhuG01XtiNDbo0TqM3/zb51KEshQ1ceLd
+K379h7DpACnluMz3wdbS7/a0pIs3aUfH64IxalUYbtJC6b/4SyQoHksFLu6EpHpo//N7ENxTjOQ
aOXdXVRiBMHecfJ7EkCmZnCmWckEyGG6dDJZByOQpO4pIJbVmbtHtUNxifdkUO8T3zkjeq9mI4qe
mTLLur5Fj5pWDRk20bMsw3EV0AxWT4sdbAFEUr3RVCoTrVaFtf+6RMaBfF0aw3pIsD7vd76Si999
kjKGFzZKNJjmtqtC4MWq+MQQwPTjqeecUqaN6sZ0LQpTPLkAI95jy/+LDW+QM2Dar3cBtgFOKlhv
j0ajLPAvnsRj4RSJJsapos+wbORtlfGQMvprpGqNc8sg+l80NF3hx3vs6TMfj6DEQbNIfZD6XOTg
j6mOsEcFVn8VDKNQ5IMhKKShHgyHDnmP26MP2HEub5yz8u4tzG+qnQsa70lge2DSNHArB9i0TZ+T
vNeFruAUU1HCXxEIDrxbRfepqJr8eykxrHrpkgJfpCzwMKaDwXyOCP/GZw63zTrhowce1dxYnEmk
1dImllWilJvd3x/v4oxiRZu5LEGw6udRDMXPOZC9ExJxPBtrtSwL14+9Z9sJDAWC6h6EDHvYq4Cj
pYHN9124cVsw5PWftseA+YtNDAhsLCHfo6QAe2c+jGVkESjLWHa4D/gTlS2ziq4MVVPE6k27Nmnx
I1GJHJwCFdHgo9aZhWQ4S0HhPfm+vsDIcBRHWuJSxQqmNHOlU2hAyVEvUNp0be+Sh/djhmEcf5aj
E3aEgnuYGy9y7v3QHmKvYrlLYW8RS3rHoxAdYW6/mmHr3KXDz9hfaBUyBUqwEJLnNVOt344tE9ke
IHqyb9Hli6hF1uXC+gbN0/nq1AIdddqBl0gwReAkAycE2Uvy4fXg2Ge7jlxv7fTw15YlGGsYkJJ/
0Hv1Spk3CpXBeVm/quoGdgRUX9VJXyBL12Hxn8zDVG6Z3QtJbxjJOQGk/biTkWGBpPfOySjLzXcp
gLaFDvcVs7n8l99Du6L5nh0mFiayS/mQL34VSewwr/SqgUVLWiTyNv/Mmm+kcK3j0bS4uww4RwnU
DgJ0hdKN7qiXAX4LS+jHaVvhJUD6OfznWAMqbiQYNusu+cVaV/VW5I60fgjTtf8+oO8P6aKFhRqN
j4jI/2jad5v/jv1s/6ylpa4v/7ajv0amx7ydWtNu5Vyqjh7XxZk+BHS2hTf2aH/mIQFe5xlzyo8M
druOAtAjr6ya11flZMFZK08PhUXtEeoNyzMe0XIDp2JdRM/4x4n2G/XKUXbiRX03T7QjDGrOfcKm
/tVChplberQPtu1my9SmA5SvtLlkV8I3t0p3x6gOnvCtEQBua9lSFHrv8/gZO82yT8oYuyNf6ysF
IzorlI3BxANrUhvewlXR1T7++b0Bux7XAwlsBUPc7eJv033aB9kPSBjoDbbXjAINzDYQJHR0pthR
PZbFMs6bPw1yQ4dIg+XhnYMMouTVezJ+1ExWDre1urb15o78C+iOU+ZECLWh34weIJ1hqHKF24Z7
je+bt4Y4Val7cgYpMxiejNJPPofhs3ezbGz8Marc4dKplzwQcqeXcvZUjPI20lOEIrJF5d56SjMT
W7XQRjACWsb4FAeVHF+ZH2/ePivlA1M3J/mNzPs1SJlhswu3R62rZ3u+MD+Ru8SS9XDZp4CKCcvb
+118eMKM/RpSw09RypnRyAyJ4yMl/QNWUezAG2/qNaWx8541IA+K+fjtV0kGrFrwCLTX2X7HexEp
Bf2bJ2lKK4cz9qOcJryiGa1vLZidEUTv/te6q8k+u1WWINaBIzJeXsbO07+lkPEZZdRU/uO3SRaj
4/yT37y61XtCbVKxBzwSXtepJjAHKrGSrf5uJ8oUwulROG0zY26i8ECyAASai0Q33nROonPgKbkm
WmTC+tnBZQ08RDbb3BIcOAMnk8iWyCics0vu2kRYcyu9cUUxyEeU2ExsqC6e6+Oe2U6nn8fvyzya
fpoPWmD6Bw6+CtKjRL3tJ6CFjvE5Qy7Pk6M1Xx4xvbJ3rXUBQYNTqw/QFb25iKrMH8Ih/fdimpHi
bqYWZJda60sQISzNNzzvx8ZPLRXl7WtBO/O+IHr0C366XqshObz4nY+ZL3GyE+fsSAVHFJCVzsaR
LLgTSRr5l8ea4BIVc3YKej62K+C1oNrT1i0rFsaCOE6D8iHRi/z5935H/1Klg0qEOl/pC+ty5FrD
od2cUM/B8bBZ2hZgM42MvpWGlxxZHFcNPGDc61vCajzslPeUmBjjumzhf1GNvge8xbndKXoYCItK
Z8nvrUG0Z5r9DlBWcWyh7PVMMW4ZqPpS0I0L9xG+n6bNKe/q1FjgQ8oj8PqfJinpT+ngUqdVowbV
qdJM+l/sskfHx5M/Kfu/v1nxsFpKogN3u3MCJib/WTgTnDJYIxS9ITlMx92NYO78avPgq8CRC4d3
GBGdC2DrZjDTN76itFRWyry9VsOCxQFDT1AbF259NtoxMwDr9hGkA1UAnKlH/q7FifJsvWa/FLXl
6lFMLlXqCIklToK5M7SwPVkgyJ09NpJyUFXkle6b456GLKOu+h0ITJHM9+w1oxemVSJchij9fZfO
7jW+HzmCigX9XZy5k4vBQrEy+CVi4lLKSeJW2UuNKuLswVPBdSK7tbtxCC12wH3Kb+tjfG0p+5Qt
9/suZQEr3qGinegN/fX408MnWb9pLD5Qs2Juyu/9DgzVdjB318HBO7uLgNag0+mNlI5aWU2M6Jwa
hymZtzd4tgSRRVk8lGgT61T9Q0QqfpBZdUrmvCQHPonygWQIYEpDJwHhRCzszvZsRbguzKa1AZHm
AgU3udf+zbMRTNB9VivgfSRn7MHP2anlMqpJ8ZjlplikHeM3aqyz6WxmjoG6CRc+NEwl8j/mzX0i
5BgUF5kTK11fb0cOm1cazoEA4/S3ft/AFBV6fndF6WAzzGHok4POmNZRGRyd12DiaIhzH4Kwxm3n
T/v8O4FLc0NXouYGlyPB3BXNj9LQGk37WCmfTZHHROJYmHoye6VOwnyWrUnjRhDrHQQfLalNotrH
RNef/tbSeF0gU0+IGcvEBqtO1VdAPou4BWsVEMUmp4aNobhVZQvnRjMkTk+QU1z2VCxzVjcHWAAR
jyUbTvNkr4osHtab5J9U4e4kjnVw/HEADPC+36wVAKU+TTbnuSLILLL4nKKMcSp7ZLcfcGAFMTLT
gaX15dZpPYbpbN7B+JVSnG8Un7BUs7+zDmScyF+ZalBWFp7po3YPSlhgCrEB6orzQCVGTGwjUWAS
a1sZTeZDgMl6Q+wT+kehZ25ZDFmieGZuRad9CPZhPEcBmP5PGa75a6Y7+WSMZxugQdnPrpLCLLPM
pbv8pKBrOFkEtesgnVKPyK7RpD3g6tm9QBkxZ3fd4SB9frtSTWvqFF0/MuqM8E0p7D3P+5eXlYwr
g9rkwp8LqVG0A4iVQnd/lbjR4kZvjHBkBMzsulSoytCId0Fso+TVJiWGd8ug+89m+k//SrAXdNHL
ADdK8OHSpKZbMtdV/I0PZoCw/zork/kMFsuySkUdGXdCRANGUDABZR/MYJ4LaXxgVyoznU+F4Ay8
gm9NGvZ9PHWrkwgI32kE9jYPM5bNirrsyQSgSsvY/K1IueHAPC1EFYqWUMxNW6j6QIEl065wgqN2
HuZcTRXf88j0AgKzNaJ0o92jYNfLvVKkfOuefDrJxHv0TSpDReN24GKasrL7YWa1UzSwEZFC0gPW
0w2+trTC1Uafvg+rnLpJXjre7vQLaYCyFAmYymXA/sZXq3LMfjhzlG0LrsQ+JA4NBKFXfzyXlNh0
1Prfdngs/PIJ4xW2O/7DLkBGtyftEny+ZadHqtfoVtC5wb9d0WmvqCeLzNp4IDNDMEZup6qrZkkE
/TeQGQVVmgnJwGaBRLR+qWvIgqsSPBXh6/GOYFHqF4ePFdHfo0ccv0gw2QIKrtQgHaqZpHqAMFQH
5jqg1kaPYrmE0pnsVqDhjUOgzyYJutCNR6NoUweS9/VBJZhrZmVeeMk5uSDzbk+8z/3WdeqZeyeW
NYbt2KgUAa3fJtAOOhL4Nb0A3YMAPSdD6diHplLRyakSCMUORrusN6fq4xrasxftBPuN5yv+EkDq
JkRmoOij4I5Mvn7jIKa9jAasylJOqeqt6f501/L7kOVlc3aSKXjr1lq89YZltKbPvQQHjHMGFM4e
xWlI1FMKtMR/h7t+JfQKFFGVQ53OBDPGsZwNszBWuIh6NmWTKYb/RozJsAQZtv1v1erOQ/V3zPlR
c92zfVfkfPjIDBhYJK92xvI5xOgZOtpvBJ7R8rzkREccDl4mOcG6rAs9fHwsM2Lh9ZiAzP/ROZZ7
s4vAvnK47p2GTf1nMmGuMT7elH/hFrGaSsn+Pbtnr9YAwHMT6mwoaZ3ZTZanUfeilesldAQHo3/0
5L3TdUS3RMCp+K5xJ1RRlTHy+tCnbCk+rbraRAoN9bJO31OLlAnB8V+77xjiQpq2QXAjUjNl/71N
UaX3iwvg/1BPdPoc1qqo3kFJBrENZR1TIZZdvUTXLa0MGxLTc2DgOsJVDfqdVlL/6lnhXlNC0Vnp
V+p9VR4hLEDe1NBMgMs/LJd+iYnlalSmHVwMjsx5Ti8+THrGL0LCh1joHjbLFhwVGBz9IrJ9Acm7
51c+UxzoWn55iclnKr5Fs58hFt/GU55ijdGF6w+3K7scFAqJec67tkvIGSavl3FUk90OcORy8Dmu
lUH8t1sXPi+7RazOtnu9Jci4o4O+XESOZOwC8Wj4hZNTHc4pG6S/z+JNPayT1Apa26LdbR+sOWpo
ukZiE1At8OQ+KBP6Nl4m85Is6o8P/mbdSRZk2ggjQUwawBekhD5WzLffW7aWiSAspb62OnnHXBgP
B8/IVzzTCsJcU5JAEwkjN7yUC4X5wKA9V+tfDh5XWcW9VSmZHk2Qjs4gsSXdstGHBrh5nUtjZjHn
unr1/wLDV//5vVCgS5auu4qFPt5W2VcjZCPX9K8bDljxTRSTKjJlCbk0bmrVPFwRPJfE+fXTONt3
MEOTVxn9m6n+/cNDXXzeth/7rSNWd6gJRLTxeiOpYQfmb/jebIXVix/jnVXUqU3OeJKL1zRYh8UM
UVCvpnjbt38HO7Uc0aYZCvHQBZa+xk8kQ7fjEn8KiO3/RwsGfusBAeZ2C74dPNy9BU60zOFDzx4I
Al3ZbJXG6nZaFyqxqw0/vPHtQWjbUfaZ4x5gRvTPTZEoqHoiGte4yRrV9XMmuSdF4uoOZYgqmUY9
ZHtCo5rZsV/On7kyag95rsib7saES2OallCzCG1fubCzWewlvhylAqg2BFCx3TxCrWSmOmZ4puQ8
uVsJsZHsjbmkyvtcI2W2lVaxObQ6eeVdYa6IAxFtixJbLU0rbczcGeRtnFVHHs8GvZ7+MJXuCr6l
FfGX10e9pzPEJAV0gnzWNNIMHaUM0Fq5rD4DCRl94vdnADEWCp2nbFbyn7BcGpGUiE9VG9G9nCcd
bLr6JMsmfAQACRRo8q50A7Vx3l1o0B1rjMxOk8O56CPAhGi7yeENe3dzodHp7vIhJRjZIimuPIIx
aKOqtY8ot6YOOzEuShlL7R/utblSt0lJW38nK0S4M039gzQ5Z13l1fmOKGFAl4fa9tgBwJIQ/qoC
hLvUD+UqQfymXM99upNejYnVqQCAlf9zH1LkiczszHaI+2pXMDyF9Gg3/H/sg7N4ky9eLTX3qBuA
HhzMV9KlfzMvttJR8Xn8BsJjDh5w1tcZnY+9/w1fVUK+PFjRIM2N88i/BX03Xyv7R5dR55lv/4U0
QCyntLXWkRC5pFf0u8FtT0tA0W6j+OwcyhtKG1zXEtJ6Mzwfck1CsB4nZtz4u3g/KoZ0vGOa657L
a9M5gwtX/IWAzesn2kdarUVKokiZgWXyzuYrFBoxPSzf5zBoYU7cG3RD9JGf3sOYdMaTTmdZDy6b
JiRWMgj6eBqd+xQL6Sx33t9h34KAMyP9HPRULtFMQRhAhLp1YnsmBaodw35D/f/AQqDZrPKVlAB4
RFdtuliwCm/FE0jRI/TmYy0Y7lke+7hd3Coyqa9BhDEM6v5ekiVaJGEanIsnniYfqearz2r7ndok
tsvObX9mxmsgYOXWC9QDb1+/niLJQzJOoIJv06T4OeXQ77+GvMtwIX7cyUQsEcMTr5U3Z6KPxu8o
/XDx9Vw3W+iUJZspCPVxCPhxRDgvsfQ+fnuBu4+hDCl/H13mggZsRSBdy76bFinZS6UFeD+VYJia
0IGueAuOQOc76diMwYUhJvBPCCMo04EI6aK5bCsNrW/iJW2wBe7BaVTKkXgpiTOCFYXSbOx8+Zxi
oTmls9FTrm63kVZKKFiMfTlEpNa65MjC+9zeF5sfroWZ6a4/Tk62YgcH2CJeIk6coUtbl6sHnhfp
I/35d3OR2CbA30+VUpHp0hDbk/xtYKOwML4tERJgWg5Rni0ocCsRB/dgt9DaUFtohjEfbYJt/Fq3
uxIcFZHDWaIY5rD/NC3CLv0uKlNWm3R2XZ2FjW8kuRl2vsJRWIvqI5IyFmPX3jP9thop3toNPYEk
7bhUCpE5+4O6AnahhH50IR4l+e/n1r+lKaP9Z2wicAr1qXOhHRgFfwZSholDNgMVLNdlQCt+lWEK
R77Y4XYMqnx1lpSkL55WhhvZeRTspwCK0ALYVH8s0g/5tjnb21YDPxHQF3Vh6OiuyMq+qRAVAA0O
oVKKbOD/t6u3/R7+NOUf4kLBmyt0Plwk0dtkF2P2Z3hOdctR9piQYHFYxGe21SknNr5ZwwJPkPXB
0dceVDM2LMcdKbyqWsJ5FVYluMPmFC3D89+DXoRbSkAw0BeqvRlfMe5/ilP5x1LieHtVeTyA67Lw
L+IB6AuPsdUZSbwGVq34qBDJlZfLqIZUiT1V8dgBZiMagGmqlPrHA0kw0bJit19jIF5RTxWfAyEK
wtPdOZstJ92ODGLdTQHKxKP9pfYUwNzlWnR/oyqFpICOIHXe57YXufiGdeVvDYvH+fFy25zXQ/Hk
/boKthdFPtqAd5PWo9zDBMxWDPCdtnj+Q0THB9wdXWn4IUsw3O0R8ZYBJ7ROliMhmmXi/VeLEVZg
sUtdsyHF7Jhy/cUMn4LaIKbV7kbQYEqDJfOD9uH5+tC0rl2LlbZYQ9rFtdi1a1l3zXYU7eRT9t3i
d2UVKZLkQdx2Bbfj6HLKvkRrpv89IEjhWJNkgTYTAlqB/3WkEY6stOMRWSzTC0CzGipmFSsHWrJq
JwN/b2UX5wmjC9NJNsUvu5jFKIyH+bw4Q6wbsMfwC5qDEkADOhMUzPX0yjHHtmUQ+u9189RH6EOW
m0Y6dp6eFJj2G4aeu8z02ZT0PaVt9STyPe+olJwTCuvni91VygPXW7pl1MFFofBmoygpoATZETKj
892586ZY4sQvuHChNAnlZomGodET6S031AV/6hd3vxM3vxKXoSnOs/ed09sRl50anAoFLbKqygqe
tW+pfMLFPce9Hb1OzmwwxjtnSab2CA+tPAPUx3jbdsFc0vh3hOuknARXrOrW6v3mFEnz4oryc8Rn
lKBaExCkJrz0Oec91/7/b5ynrjG2vxbAV65/UNssWi/rR8KxFNA2GTjS9O48aOZFm/16H5UCdWKJ
Cx2UvJPLnDhzodkhPN7x6Y0rUcJte0fWRZulbhlL8R7xidgB+j4Qsl5CvE7b5qVGqVevFbUGjb+x
vhJA7X0CDgHqeQiH9/sAgoXWda7AJM3xxcWA+P+VhrjSDNDalUvGy3vYrSGGqxty0KXJDZqHarEy
Lsp/xSwRJD8br0UsuORbmUaZ6RC8ZWLlDZ5cqduAc4CAUAN9LH5yrKfQRwf8iehUOUJkC9qV0K3F
zXNOo6QMcKOGCNZwz7KlidaZVw52ZVr3jjpHoUcKTIauHK9SS6bB4tqC2bSkxusq6OZmK025+GRs
6zo/Uhcugko8NtA2qzhE1lieHfGE3bujjg+4uz9x7gtMYhTGMG9896OEiakALXuw/5SD5TvVQA7l
9U2hPthmOkhze1TIoX1MVVHGPt722JP6ElCTbnqAc6m2FMOMVj6eVsLstlbSb7k4kZmlA4kChZgD
0kZfxMcgmYey9usOYu41gaQS7bxeld+zfkXDaGHKJ44wQe4QXiORF2V7YRHU98cgXTYELwIMnDQe
ikTRR22EhynnyjyKUa4SpYoRcX4zRa6MA7weqQzm++6xIhs4XxybDSOJM4ohHz89qAVp3DSwLhqg
hL/sy/5A3GMIrg+oWyM78cb7dAItXQT4Vg3OtcglI+7Rw07FaIFzkESzdFzGAgjqi/r6aq2yG625
Y9sx/+PPUfI1BPOx2AZ18PMQa+1JfUQ9KZOL2SrBkun+DSnysj0JSfYM5EhnXuQPbpx3VQJfzRrN
mNN9yAxLngOADWgqXd7sA/l4nbQgjqK1O1P2pThGL7Sq+h99pQIeK0kQ2YbnwFOMji78V37JaBeH
FezqrBrnZiI3QGx1LxMqPlp9CSee7qyf/dGJ/xoDys7ZKfQ31NFREBV0OfWP2fEg2lEUmCCXQYeJ
f4oxZIx1LpC9KBsLR7rhb1zs0a/m9j6FpFIZ/iym3LrHnBV/3tQSP9npAUyuuZV2r55uV0ItjAXE
fhAYNRKH7t7KWXBYx17Hk9dFAjQzYhCfg5O5v/NDMy2E3I/nmuqkHR1lCHZJkQ1rCUuvLnq92SC7
TvmbXxrq+W6bcOaNC9T43XE8lpUliHMmxbROOAnP6Ejps0T685w8WK3QCfswwthAFyi2NV7oQrGR
Ai33ZXa0D1WJ+x8HelY0emrgyDs9yCrBt8+5MYWXzjmCpllx9fdJzsHS+NlCuw6fWwv1I26AE3sM
036LNq6AdB+jKesBJ7L/BE8wy8M3M1WQIDRyY4ADWec1+VnON5IpyrXxA9tGkLM/IVHCIPP6v7uP
grNhfDzp4BYy4M4P3mABktoEC9nhb2ASq3ITnG5uaYCe7lHtZAHBgzQ/GsTgWMWBcchYl0OYJ3CK
Ch2n17LcRdI8txTqkPvrKabd98Lb1rxd/OWiL69WleFyyMIMT0BDa/6E8BLw/67u/PbTYdoXN6Q5
V6Xhtf/yHi+zS+9Sjffa7f2wclyHxBx75sbf9TaW19/hwSZ59EuC9mMczMWVQdaJx20dYxi2c2Pn
rzPCU1O31LTvLwfWfPzHh0U/KR9LQ9QvqPeJ/v8/talHIb4wSvGB/PwGJ9TsrU3s+wUy5r6tqk9f
7ucmm2Vz+m879/MEQMXaEsTkZqvZ8hgvOWpss9wosdIzL1aO94BueOLg1xeKAbD3X4DHg+tkmJlO
3GhNrrP1hxCOL5aM5vE90Frl4NdzNawpacwmLGC714XiiMZsAj8FyjhcoFKLS07tTxj2/jwvjKom
j2kjiYN57waLAsHb61BoliAF4FtAyXe+Uf/0AIh0YW7f7O6LsZgzmsOjVRFFZa0eupyauh8zEELV
08eRrOkcNWab2hO4yXg5Wai0rOyP3NuMk2d2d4jQT1OnvCdDKVUoeXWGRsrT34VnJtwKVN0XSeEr
HSHa1B4tg94d3sgiUWJsN8HKXXRs69bKc/AtIKfxPN/1KojsaTNn41KkZqTYMC9BSQvcJJTbSn0S
fd4BOxSVZ6Hd/XU8lDzVn4vTReuLYv82WzcSiOLWrQndhxiGFsjBcyleYCd/ypkBb/T35yjod/8f
3V0CDqt+BmLh+FOd7h2ao1BPN46QU93zTxpPpyZpmxaIGoTph0v27DtJ65PtembksZVnr7FHCSt+
I77EDtu3c1wo92u9u9Rx1Hsy2hK43gGy9cHAiukl4h+XDpWoIEXzePl4/FIHdByHSC34xmz38PDD
KBQKGj+IS1GY8nGA//921jwL2SAVW2YSCePPBWSigFKFTjiB8jBoYiPxtMprPBUmjMhfK6YYsKYT
EFRPs/rpamxT3AWt5uJ3l4tZ+ilG1hA7CXjbJtdxRosceRaauLuBmj7AiNmsaYm4hffZQnYvgTbH
n8vwftAvFcVzfPtr3PeI07t86lzWgokrwm53WkD6IH3TSSbH6NUT0CjZrXYiZwg+fxCHFa2gGBSq
0LGhaKXeu9VpQTW7XWTVKCfEfqH3GtZIsILjGKpr+1kL7+aAvyZrW0RB6r74xbulUJWY7hSEt9td
gIScjt+tqx7g3fPWGE5B6vzJO+ZPHn+DUehcSRVfaLoMwhNbzarDoPfl66l7hsdjFk03PSEHZURO
10ITWh53MSOGV5vQvKVVpIT5JMA0esux/WaV5ASB/gW8LudTItTANOzWF/RiSNIZkOjEFkVIed16
+YJpz1rGjfBa71RcaR4Rmei1YNwZYdv2qdE03v0YAIFc8p721R+t4+anOFocm6CgySqtq20M4Znm
8vE1gYzaB2tApobl0qyJ09/f1eYdCeijUwlLKAxi/yqIZQuSuCMWz/Hv38SIMLjdF+OCWYvkJMjx
Cw5e0F3EooM3V9MaHtVDRmHKj3HP+c6UOX31rM/jNKNaZuXPhJcc+1J67tATkO8Puqe9fq3YhKbu
yOefRCHxgRJ/ryrIhLcgv2/ntj/gM4MRd5ZMvbfDZkwwM8NeVnk8cyB7ptmrMtbm+V7fxWGi1Q7b
Nmii6oydmtFEllbVOGs3vy8Je4TLm/crI7z+u/o+8FnI8uvx3/Qbs9x2DBbClnMr9kEG82t7jDQc
bkOO99fWQx+up4om+C+m+86i5FugQwq4GObkV4p2A9fvJtQmYS5diRVNq0tUMovN4erM8AUuuAYn
aHh0helbt40EN4XYbHz7tfNB9/g+dq9scO4r265j3rfYXgyKOfgemXvBQKwewZjgTA76ipNgO3rW
ZhBZOrFWxr+8MaYOALEjMCwcacNkpmWEgJLfWXM70HZ+DsaTJcGQWQtTGJEOnxrwUr5IjJnS9bcB
+fRKlhExlcRV9UhIswI6PUElKE4uKmqIyz6nb/niG5UOr7OMzEz3s2WpPwqk5wJq9pWZQ7KfwB3o
E5Wqvmt15+Ctqfevo/LjDs2eD87Oz19OPdeIPBXjobQKU1PpMWKD8TSRyF9JZ07rsK3WPw7OPICS
J2XsW/GCyuIE7LmIWgDQMcGRYL8VdKub5XOIUZ9pLlZN8RwKJ9CGh82v5gIuQsmBrCShMXI9P1tO
2j7mmS5sFfgsW8VrOlqHkceh1wFviJ/fnQS/Pl1kJNISu1nv52m9PYsbU7ysWB3Pqcx8iXj7aSEi
tJ9v2EQrxAwNzkc/MGAd94SGrRZzp9zfN4Ke0LNeyPNUhz2DhKRm1BzuSVf8P6opYa+XpjKl4Ftr
WdXdpsOlSKUWHD1o2N96iOGjy8RfvFAES716fnTnPvq3o2Qp5OQlE4wwdCpYFq1q0ozMz1vMnzlF
Ma6dPubP/6KDt+hXfoaOmQF2q4L13VH6E8Hi5LqOrhpYuQoavt8PhpFXEclZrVpD5uXWNSnPMBWP
1lLeKHtGwIZwgW7PfpyEaX5xol18dds5DKLr607gSkEhjg9IwzY1sTZsRltG+6hdVBG4a17OhLI5
mOnGdEt6iIvQGKzQcqP3nER9blwPuSf0dv6EdpPR6sEMr9WPgjLruWlkxF4mwMlaHOaOSkyhmLHJ
pI4pIJgmJYXtz07ORk5J9zBeJWfxr6b6jFNBQRDL5CwmL48VvXcEUEI/3AIgYQ9l2oiIyBIKGXlS
lEEQjGVGRLPV7U/DPg16YLCzZDqE5q7mgkqrkjtjFu8X0Rg+7qnnN3XofBnJUHGNlD7F9etEJuFj
9fhE146uAAFsPq4QqsuC38YXWxlBaXd9Wr5JmWtSHiMpwp1C2KobRGQyTjcxqi9C3DgsiNNxtf1m
cznWzfJqhMSIQas9uNmEfV98vBPhZIuL+HTuBhyJaHfY1BldSPb9tKrcYj15y1IvFQT3Xw1kJyMy
xFW7umFK6+nUCdDiH/AK8mp8bv0U6z8R0xrXRqukJdzkxYcV92RoncHxhZdqwwIwT1HZVZu/YUa5
VgXh1uGo4oUst7Nag7/X0buwvUdFYXo7dd1s7ldK9C+LRZnGvEevWJfk3ljrO6d4H6E0k/aGHsIs
QoI1wCkos1GXahI0c5jhUu2un3J9bbiGnQlygNJzzr4uoIe3/kQstuZZnwqi0hQ4Ubw32p/w4M4R
6A84wji+7DU6lRnJEdVDL+7jg6QNFdjk6fX2t2Tvl+Ap4S8EOu/nFNuKL4RZWLpGMD0xmc0WX5ro
Gb7wNlC8nbb4CQixMx8or8QgdPRBMCyMlLz3ToQZ54NdViYSCgYjCFcbX3SS+hpesuSjejPBW8je
c+kI3LzYObsb32BNW5OiiNAMY6Bt2574E049RDjhxaxY+XnXH/kYWTQXPMG9dV6MyLlTmoUPwgTI
GRwGA+KdF5Wj+25mn8N/ACApF2HL5weDpvsqd5q1tICWIIPcsh7xnc52xZKNsEUY+YyaePNKbU+f
xDkY2tlMy5No3fPXNJgD4Ka/gBTjrJHrz9/Vs0Y/D4GN5o1arPIbDELzuuuBEDspezRS/JApvANl
JfcjQfiOd774RxjOVP8w2FFEsljSpUAJGqMmT12WbPw6Vz/kqfRdMwnL+C7JmK5HT42HVHYuSRYz
dybzdJ8d8S8q93ik8ze5A5vVOCoPaIoYgZW+Uo93eHwHiKze0Ij/UXkmoT0ylEXLzW4IpbiURUj1
ywcQlekA73iA0gnSxvBols5b0DUPZWI7cOD7EzfvFbS7+hGDb64EI+aEciSpkE0B64312SJzKj+i
n0Bw/FnV2E9oThjgF+1aBZ1ph4eumgNFuj5SvMsd+ksj2VA5faNzKg2n/uGp6LcJZsxMYFv4GaXw
g09d1Az5MfClX6VjJA/aQxs3a+lsnEFb/NfbnZMwLUf7PQD0CiXnNf7fId4Ivgk31dMncrUnKgJb
ReZ4bE6tnnlVW6EPJWC1praZRHVrpWQCGHrQlFwOxUbvdCOmboMXJLYYhLcP077NXFXz29ACltw4
44wfoz5tjGjef3VI5kkMc2gibAfU3QfHxhC3QPNvcOT+sG7sv8TLYbz4UIagRGSK54LtngTd3/9c
ZktfXb4K/qOOeLAnTbdFSv5eYcKB+/CdJ3q4eNbo999iCVqNwUM//BIuQZg5QUoitBFWebbTL+mq
R/03wpfxJy1mQJXMvawcC54SBzD0UQEgBwcl7E17cn508A85yYYB/sVGIbDFZ8D2qBf+Fyd44Fb7
mmwYGri83LZPDHeqmJ4XRpWvwXZ9/N063StfyqEYQMbFfPVJorKDb9K5ZIttIH604MwhgBrqptdf
muf8mS1KNZoV8ghFOkHd31JSsJMYVZcoSo93JnbIPeLgP6/6FAmragppTrwk5JQA8+FbxMl5kOj1
dUBmI45bdC3+Q+PzuZ+3BTXbVdG7T8r/5AGzKeqQC7+7q3RB/0aqakFwxzMvhruGO1kD2Aj0FL+o
d0t0KyIXLVWgw9Q+RHwcHo9rSpe9632U3YFl47CvmK8pC6Ay+85JK3GV6cLnZN/9SmiruIoIbZDy
Pyuc7AAxKSNZaJQSj7t1BxSNxiYweMbB6BbkqqeJ5BGQTP8OyA5+qt/mVlWYBQslr+sMurc0LljR
tb65v4jLzQjcwaKs43uXnzO546dIjufycGj4q35Ks2/cB9GioazSmfMD5rkpI1SWrC5nyAge4O8W
e2tD1zQHpgIjRrSNu06Z+Dpg2PLI/UQ0w5MnOc0KOeaOHWa6HjRDygw+MXezFqzkNi4Xgg+s1H8X
rx9MnUreRTpQ2p9iQciwi30cxCwwhDoj5jBWz+/YVCBfnwjnwR0TxBILzdAe+9WdDpa2/ALrykpm
8xYSHwDul/pNcjn8rZJDqbiL03GyUGhh7C8Vi8aoKHlIuFTrpB9yYgqUtu7rVILEllk+OgyQhzaZ
bOxTWvSzBHVioac3+aKAiiPgUbZEtqTsJTt62btkpFp0wKuY5iBECWVpB2LteHuyxjIBaT7EaAMb
XTiYrBtKLC7q69sQBn47e/E9TBy1UfnRlHW2jdz234R+V0MRFHaGNJLRNB2BqM+RxmO3W4jXeEng
2i7MTi5tGadKCDXoTg8GvXGaRtxNHR0J6oaY6RQWmNl31Mh+LbG4roGW58x9kZKMZr8WM5Tmhnjb
9BEpYGxwvh7HzruBQKzzzrmUk7HreC+eGgj6JdOlpbGHml/tANKY/CEr3wwCIFICAPvp5lUgotoA
UklAnBzdQkEnMtmQRydUXV6RHq0vsVakg816ASN4uMxT3kUZVs7QwJgbbHuh2ZDS9n27fbA6HvB4
5FEhfDCCfZusyuRVpGLj3SLQL6oqIQogvdd44749w1MNIQfwViZw6ErJeJIk0IIzgG8S3SrY6PUA
roZtjDGPBiozQmSNsJsxn46kDUPlpv1Tmjs8jsN7XBHc3IJbETxkkArMVhIiy5oY021HQWqnOR2I
08M8+QUb4QJIPCZBsZys5PygGCR+SBTIpsGDbypXHzvaXhQ7m+JWezDLVtpf+mmWKRCYmLM2cPuZ
39tc3e+Io3tYk3105yG5/SVE22uX5nqdyQqQftSDKfrciITYsZJIPz/oxGwVbozwfGhtGlzhCCNp
7fsgH8nhx6Uah7ydk/zS3w7QPBQTuCLP5lYDcQPGCl1rDTuZGnEJzETk5k3J0GqrtRFplPiA85vB
onRY8UfOdpY4nQs4dvdc5s39Rsshvd/oTfMUG4y2880sLY9VLirUK+K48BzYdTJ9g55D2Mf5uuQP
EzHOQq+cIoKGFJLwCPh4YpAgIv/1bb8VKrA8WMzEuy10sjyZDDxvYg8mrywLFnRf7oUEwGfoy4ev
/ANCHzo3b1i+4d5fwU/hDYVnF5tpWQF+YaOOtagojqbx8DeO7KLC4yuKO/o7qo8cV6bFgbiPZOZn
84bEup1P+X/Sc/hEDZvnIx7zNajqWC2lVi3HKoC5qt8JQVRXPbvPAOr0RAkDXJnWthj4U+CJRh9F
Gvj5Gmi2Xidh5JrjNAFmNcnSbdUPt6UQBuMIuSmiqz77DfVx231Oiy95nBsPrJZ5dzpRaNbRJY/Z
t8dc9TNPxT08dJBlmbdc2pX33EzJai3vng36uiAc8pswa7M6eZ7N1NwoBNGdhIlr6g7s4Fmkzkhp
w0IXc7eoHp7kPZvyrK4Xg/z1X5QzqtRFX/zZn7MPd7R+ImriC30dxIkd6Af+jizPQWZTEOUEi5Wl
pC0P8xJjKxVHfgtx4xEZPOAiSuL6dVGLLwq9EuSVzCVm9sEX/AvY/2CSw3BwcziuSFcgf5+ny1hC
/MbRDUv50I7rYJbnbmOrHXjGhzDXaLXCs3On80/evSdkgtiqCe4H2NuqoYM18D7sKa0SDt4cQZuc
IpPZViwIPDYTIqwZdokc3Q1ULylr73YMimFe7tdfb+2afCPe29jhj35oOZinRZq9IVkaviqGSAOc
dnD1lzzl7WdHTBex2A0YNKcteKYgawjN4ZnjnH24GRdPRoX7Qsq1qYWubfZWqUbsPqjXBW/zEh8F
I3RdpKmq7+4cXSUvaN0GYRdNzBMAKWWW0ZwoNXF0wr3r6lniB+lNEdI2HVhTg2lUREKbETaQsAbZ
Rmi63MIgEg8vSVPIXUydH00b59cfSNoxDBA13ZUePfCUkIpxjRdetltUc0iJ2RfdPQ04WIpv9P5E
u6OburT+QZuHxqF+kCv2lVGjaPygQyO90e9+sUUw/Vzk2az71J0HIMrNg82OX2Q1sPsUH8IXhPyX
BNlNs73+elIOEhUwHFjTM95ZsXEbvPgaeh67WLC/dDFO0KaiYrBZK+0GnvsRcwxyj6dIOFToKknK
nQiy6xdA6Amy3MceWUALS5bRyh+wvYLhB0Iu0YqLNaeAJ2px9ohVx2NKleOOoWdj0TaOUprPBVsJ
W4CcXJVHK8ZiWVMlFWdLZHJ/KdQUyCZVhYShk2Vt5NMvq/USpdxBI3RjGHiN7nWhqQxrUOcJLird
UItmW8NwMlrug+lBxT8ar4A+uoiiNc8FZ/wjDqssLHsej1Nh3FuzwS5INk74OWqclZP1iPROO+Po
V3w7SBdbfABGBMbBUJDJRMR+eIa9HMX7ZobAmt/Jr6kt3TibkgtNniTQRHWmNdaa75rRV3LQ8QcF
5O5lU0qVngEjYnuw0s0fiutEQq3D6sgplYP0ELXG+e6PJM5JZvXjbIo5/nY0pyIjCgfnh1a/VCiC
0/4ubJaCXJJGRBqhLEYLx6VmkOXoRn9zDMWgaNPNRgzi3lfX2JiGKXZ9flcDVfJB0el1LrCZVjwa
vTwu9BTWsEwvxnZlLWc+YuhxKhDJJKQI818s1kQS5BdFE7hJfhQ6+/vBJgtCruS8ggt/SHKBxtxk
4KRX5SLV1kPlpGG1vdslTDOmWxBTvP1iIh4nBAwxAnQDmGP39xytV9ujBgBLCN5l1+eKIOYWokzH
Ifb4Mn6kWjDJyrJ0XfpTb9H9hOChPIKCRdJOGMKJZyUQKp5L4xtfxt5hHxBhIqStZ5x0hUBIVavx
n5bf0wFSRjhhBNbA+qUivyYRmclHSHJ+gN9ANnqpqNACn0GmATo3Uk5U7+1Tp1uvkGdPChy7uX1i
8pspVAg1w9Z7S/xn/BkyBhvaqu1/2YPuLurXwT3OB3MswL+/8Z8EOOm4D4gTCSg6kfokH5+rPb0l
9W6BJY1iW7cgciOX+OoSCVnjV8GuGTX7vNN2BYDUpGkzjxGWNZbTKEwn+lzcbzZln3AUJrQHN1hj
1f2UsUdo/XkaXL3R+wd2e2I1K27H8H06hEL067j9u7prDorla4B9YuRtmJdbRac851Yz2KgWrmB+
NdAQmuEowWuglRQvFS9mHxRJPeSojCGQBd1qCAlomY+Ubk/o4wtwF2+Bgw4pAg0mKX1nNCE5JULk
X2Q20xGG+2u352mAXwejrHCnJTn4u5kLQIFklzJ4X/qaoarBbCoCo6FQQt55PnoHddesvnCyxp3p
xdl7LAsFeNjS0GEvW5XpFXjlqKQzeQWjpqz3ZAZh6xL4MqOgc1Rct1C3swh9fQc54Bt1Kz3yos5N
w1VLi19UJQCEr0qfN9rutuV9owr252kKjQGCgTKP8YqYwPfMDQrt23Fqf7MyIazUNx098ujGs1Mp
gj90Qe1hkZqmbjT3RmyiRhPOp00F4kma9dgSWBvHQwrParn/lcXPSd1U0RMLWYh4ERaO+EStOh5X
eB8jHrACFNDY+wiwZjIn7sCMpnEbGScHJNnxVw9Qo0TvoJaI4ukL+YnJzYv+foaZSSohzYoLMXml
7JlUEI7bVWCsR+/5G7fWmCMwyaWsw/jUQHFTxLcFvF0eyPjxEJ2rgWg63lxMoHq9dZfbfpuCfZ5A
//BdQU0RymnEz9BWX4/du5msjIp1pB2pqEKRpmyUApe/e7Sy36z+bESvFn9Wcncfn0nX+wv1o+YG
M4oqrkG04fzpy6BQhRDtf5IUKO15M2xBnyaPiRkAQVVI+v8q7+NkDbZKrjf0EnIcJdPgGpcd7jBf
NkzQIoTbEexaMvyhNx82E2I1gG6x7BnPyRHhoB47D6RROmZnes4GepW8D7v3iuCqzptBHPmsOFHh
gKO00Aeb0G4DXKP0PJZesrRffGRxpJtyGLbslSaKoE4jirNukhFSIMMssFjIUU8qRDrUVSInUpgb
tMinYzYrCSQ5XPR4HpzzvWGl0OkT9WI9PLnkChgnjXxIOM8ywY3uVuHERXE+xqrjFBFB17nfMMf4
xtXz2ICdoOgmU708/qMfEjMikncaxHlMwX0aWpawfzvqb9BMIaVrJKp05qaAuSWUOcwy7+j6U5A+
2Ei+6c+m6QnOIKwSGlGS9f5SSXYLc7un1xFOgrMIowutP4jy4KeybuNqBHvQvPA1Td1aMwrNDRTB
tD3cGpmhFsnDlSFbJWlhbm4fdCPqTo8iplGFgKDHE0H7cqi5f4GgeHwH8OMh/7Dzmv0v+P8CHnCO
8WAem6G4n7SXFZc6K7YtwhE9cK0njuNN2h7UptgjIgd5nGtg5UNubIG9Nm9f3/l6RARHUIXTezJU
posOsBq4suJxku67nr420car1uBpf2uCS84yt8kEHqEIZdoZlmHjvxh/Un4X8GR/+wNo6BdsZLxO
nLb8PEoHsjrA62kAIX+LtUGpUSOXGMehUNrFITuc+9zkd6+NzHPC+uKWNjA5pH14tBT61PDhjjC0
nFERjuHp9eMHZelKOx1zFPubA3OVCfWoEXuLShGXysHtmd0f8VteFEvwW2t6lBHxAMbX1U+eC/It
3jAzdHHWu4TJPPVb29L600U8idPaKkCWo996LCQy9aqckkT01LR1yJ86n38Grpu6/Zc+Vxef8DEo
al14RHdB6kHDTEn4Gf7LsneyrLDemWzGSPv0TtNi7TJ4RLnOumBi9bEVOs0HJdQLtf1Vl0+oUBE8
0HXTK6xMexicwtGinx1NMwz1gwTYfPzcVPSXhlt9M2OOFW0xIdRlSB3rijNvsg6JFff7jwbwAGDG
I1Ghtn2Zf2ZOe5Fr3Zm08NkGopbcf2FzTYL/aSiJjajt3SyQlBKKYVpPFRPWWvMZBEa5ogbfLpNT
Z+rCEkbearK+Zq0WAfX86t84lGJWAE+MzgQga+9NxIQo6aGbVWKKYRtjaWlzvjTtjTqPMXF0gqUj
biCVgf39eIOcdNKnO2NizKKJ0S42AM7J6CUIZ8AL+Cmp9vKqB/vRMvSDAUmVKbgUF5dcRseiD3I3
12yFCOKfzXAN8tO3gQHUKRkhycf3Z4CCCOGFZH//LTbPL4I4fkSUJiAogjkzPF5IrmVDSXZ8fflA
S/S31oI9k7YoieRW2YJ9UL50pn/psalYpmjXXSA5NRtpnpsUK5gdLIAKiIk357tpd6sGFxkfjiUV
yG2soCU8xq+rIULtQDC68A1Sds4WEsZuGs3shHPLKy29M2W0zhZ82FJPwFvceNfNAg48itoO0MSk
IvMExLj4ZbpAWhq4Nvffsuf3S+XGI/KLe1DI3gKFBqH/hksltcDZRmnWN3yKIUL2aVN0CumPRIRu
q5whUnPvq9J/F0fsTKWJIZ6d/vkBmoelbtFKSWURZuD6ARtUiW7nzZNQ5oROBXeOHu5Kxy9DF4ls
/cn9qFsTGv8cFJsDERuHMgVyfttOAvGii/i6mw3fnuaArp8C7QHBwiip7EJknR408KM1H2P6couK
Bu4x33alS634CxuscVJghswx7CCDiBhOmL3Jy+bHaCIXuQJYXTGp5QeKchNma9DIewcOyXoj2TkP
AbP2vmQhYXjcE0rdFa5F7M4n4Mc+kW82EZSwe+Z3L6Uzlg+lzeRZaCU2BGkBcBJDjoG/2zgAywqj
Git9VlEBXLGY86XHZCyDAiiPvFlTn5KObzmaoPdRrD3pnVdRuWictxhN1JWRVuSSksT+keGRcxY2
dyqpyL/7mXPK2d9DDSRPPxslbHzyODJbEKSCQD0ckpbErY1G373q9vTZIq42woAm2GKgi8u81UW6
g+2r8gs0VS43enpn9JlAfxNXs2sLfDS2FP1Z6DI3AeGoIN94SwdtgTKgKEJ5QolUdHKgUgtx+rMc
9dQTCq31TdrkNT6tGryMrWWmVpHT3eDraH1LybQr5cb2Ggl6AmUcWMjkSGRli8YaKDEy03gLuzIs
Ho1II8phRyT+uxKv0UHpsy8b7RVyb2Qxv5PDyl323fGkpe8Yqsv1oWpRNTTLvnVoZPbUb+4ILWRE
lydYu5Vb50c4v3jZ4Yq9IJs6Ala3eV2xS1RzkXeIF+JBCApO1M85E0kk1vG/sNVrBbIlq7thPE/j
M5iPKUnqT2lDt4W9otTNYU9oht1T9AM/GsCowTah5dSOAC0Fpu0Zr9b34U++AUB+OX2JBSsRBr8V
g4SU4mIDduATD946DMSj1eBd0TrKFJlWwZ5Ks0DsE24u4JIPe9bw8lYZK0LTJc1WNv8WBd9G4oHK
uX+LJtOa8etbnPpptpusbZnEvIl4KzCU1UXmk7ZrAXMuAZCZ+oQo3Rt2V84Uf1BsaGGVmvr2MlKF
Bgs12aJ1bceyDbr+IRGyKpuDMKMiqbCJVXGqHTHEsQEe1dymRz8ENbx41oBHfGOmyLC2w0Aju6HN
FIa3qb/sislFMFBdEnIuETXgf8WfM6SsjVlqES1i+/Fx1pgdEKd09pcZXCX5tQeHzxPmL5Ky7Kmk
Zj5D4AJ0mlYbfd6kQvho1ioGbPECgWIfjEttQzxKaL6hwMGJIPAAMdfxjYStFXOC23Qb7/lrKx4X
VM0M8I0Z3z8L8I5hSyoQpogorhtyZevBx6xrbtgq3gxvRNQ+4OhuR1uhWkbYLQW1lyBuJOTsxkSh
f+vH6uN2E/bhNSvRHKIvzFlNv8UtEt6q60vZseWPmjkUMd8f2M4Wo1qvLQDIBywoL7X+Gq/KtMtw
5SQ7j7Z04seLBbtsTbZGeWC2fHiIskXAlvp9kX+yuQOkAOgAYT33FzCeLT8teHQYiSUgtAqfEauf
oYZrWF/ho/0S3g1NQHSY4yWmDxI1HmZD055xjbOWqmVVmHy9JJGXIW25f6ONH/IzjMW0IOWIvlMM
DJl6UHgUcZl+awPw0Q2bf+EypthO9KWoWDc2dDBN9ojWBPVWVGUKTfbpXytQtxzM0RZEzPXIZmJO
M4hkkJ9iyz4U1JgP5dj6fRyVTYSASx3vRXy5lhLOehowEtJT+QRWE+/TnFjPpDeBBt4bq/s27p6N
WS3GvQiPeAztaVuQFub7TIwRlHZceLt+aTPb2CvMR89iq8cwFdw88virgniejN+aj8D2fxUTrscK
PONUb7tlKUu9Q9OC7GMmVwMizrUVBqRQLJgrGEptMwC8DwtszSp8Bwou/FWtkJHFoViy4H24eA4C
J00UoTZgNeE1QPc9ZWgZC+lrRYiZ2AhL3+HrV0J45vrJmUYP35UZUFu/zT09HFsDjxDkeZaghuug
tLU6rKMRouWcThKeKOGaTiFF8m01gxQfMA436sa/crEaCh3oWDdJ8KqVy3Dav8vizDFKPDxqYCkH
aYJcT/DXREXwzwm8VokaBa4Hl2CsyXO4quIBHEhF2GR4dqqNZe9Ug5jSOgVUsz4GHF5vb0TDOOdR
FJZHLvBe9JN/rG0pvI6tb4Xgsq8cBxnogeRUy73dQAyEBmmnZpyUyb648SwcrD09rZOWMqgNGeXI
l4jVyvTX7bB81hDo5uFwSJGLWdFnaxQyXFI/EwvoICV505AwcaYYy2u1mB0VR42Jm/A/RVJUeIBQ
HcMyPyrKLV8IUXYZTFpXpDC1B2AE4KphwqclAH+55apR0sgqqX1rPSxsnvv4otiW6wzsgfD2eHKq
CEMs44t6FQNkwfOSblUuL/hwuAGL/1llx0jC0g/fgIY3uroYB03xRG1mMn3x1W2VGy87xFjtRg5K
DfxjxL3R4VuMH9Nl2wjJrbA6nquPouu855CzmVf2PajSTX3cSclXyBT9/chUXl/AyUrJHnlbeifZ
SNp8lSBWHGCy7iksb5f4ltZvIAnEOjLQdf1zhkUidR2HYaaWjYUcIrYXd3PjrFtcM4wEPzWHhNyA
tcx+6l4wH5TPXJyYJ9aK321nGe7rUFvo+fCrcELcHLaRc6NQmn9dtr2NtDcAsfnwIn4kY/GreuPT
JebYo+6k2WIPMcaEsxANKdDnYy1IRdifpTgGGDh783uEgaRmUyvHTaJH2Q+N+9LbjjnAYqb7r4uo
gHRu64gsfm7qVieTcHpMMiMuppRAuaIQm9nMhovMRqTzBa++Lw3101RXQpfVQAltgPLuUV+pRaQb
6vSGm4FhcH0rtkkI7wiOHaD+WxIQfdn+bjnr24Kq8eQgxdOgZMsYfHpLNze6sS8UmxjZ1a+fhYVU
NFRQrW79chmRVeOVqV6Juxd7hZ8pHkjx3+zhKyr+Z3PfDs07CcNECJKTpW4YD+4lasAj6iijbn+K
2jayo+7CFUHoPh3D1p8UG5zDPRb8Q7zWsojYviXbfwVRmLD6ISgWNzz3uFhy3yTSEJV28LuBp8Yp
e0nwQgILsI6lvn3mH5nXI8AoxtXXtujFd9lXJVkm0A6Hr/0cHM4mt80Mo4v3xuV/i35zuE48jhaK
hiWUEoNVidCWm7h/sctHkJ2CGybCPBve6/iSc2pQmHU7TSkJUqrzcdByKBJ6XVRzgvZ/TZ18Mcrw
c7frsoEAB+pJgH/ErnzJ8EkHL0mb9gs7RA0kNXO/iO6ZBJWRZUEkTknQudd6GmhtXku/9B0JDjDX
RIQO9Qs5lMhF5m+p19gXeeLno3zn5WxED4/LocuYZ7ksbB5X3lXTjWY11tFvQJOO29GHXUuof/+V
oh8eudxouU0fHKuaBmQ1tvi8DlP0041nIB6X5OAes+czul5kBPKwrNZNiolezVaoyme5jLreKio1
djhVuyjU2EJZtuBqwxT2iRddi0DPFqu8Lmq+3K1eNDNrW2fHLsAAHLQ6unx3DHaZRDlkl/+suRi0
SrbMGJw/ChYMONQHuZKdilN+yhyYjy40ZHVPcHPNi5LEizE7+lE5sTFimBF4Y380BwRwTjRI+E8w
OYGnzF7o0dLrNqOHiRLTwYu9qzvzv5U1ouCy3HA02hYD7ECehXuvC+Cb2/aG+YLZGjcXPSsiaxax
M8R0l01RltHJanTMCy0iLKebV0n9b2D/PwQjKi9wbuYjiF/+rQSTE7ou040GPauvm2uR5ezbuCey
wlSHM6lIvvY+lSX9gZWglelK3XGdyAT+d0wFsVUB/RT6CqYU0KYBy7jjybNTu569z1tzIApHcayc
uVnQ/bhyAhjKaS3i/vZSCeiLhj/MpYhz9jXWmJcg3ZvIdoF8ndF31XJXb0Xwh9rxOnnxs3519EMj
6G7xN7UEI+Y3XPesuj1y3OsP0BvFjKYtm+Ypg7LS9+nt6AJMKlcZnDADJUHcNUnMdxRb8ymRltf3
Sxu+nrnETezI8bqIxkFzEGXMtScEm1+cyER5YdavGYzhkXa08/5EhmQo8pq+XUn01Pqi9ORPa2tf
7aXVsUkfyOnq2Ny50ouDwGf5AF0usHt0S4n6mh3VvKFDoDOmsvpIisIcUlyq7tPCb5+jkY4pb1qh
Hfrurzdl6VfteRjk5FnwR9a48GgHdYrhK03yebEtK8B64XxpIC2TX8Z61AIjD+IfTxPLydNRtXVS
U8XtB5BGg19wNFtPgB/6IPVB5BV6WnPYw4VpYTBf7bNL0DLq05DMeSQfXl97XBwQwDGzj4o0vK9v
J3u248iyHxaS+uiiaCupULK7/Hbr6pN/xuxCMxtZ/8gnP4bvG5h77s6nNE/ldZPxY8QowdqiupGT
ABuzjBEZobSZ29KrKBgxHlol4pBTmUdiT8om3E2U3cRZBR3BYZE+3vrUv5TQiXktqDXh05Q0jiJp
zo1GZerbcVyxfHbURUf8dVLgGFZu0iDA6J6mOgSH+JrrlpgpXh6IFvsmNu6HC0miGvgYCSs+Glta
kfW5fPWS6ihM0RCIWqp9VHLyiOQnX/4onjV38fqNTsaQQMdh3nuYCTlwW+Cno0nMXyeySo1nA3Xq
pclKnyqgsHQK28k3xM6f+IGUWbY7cStYhJvOMQe2EovyVkJsaS5UZ7smZeT6eK46xORxrfwLH90s
M3sDP2dAYvSRExpY/Z4RwghjbLTzLCnXJBzdgzQref/zMZRZRY74EI+8dpSwuapIDQDgjfcU6L1D
UN+F8fx2cLeblxKsrJJE9YPi0SdPxSAt0w9c7aVvRvE2fOziBsO4nGcDK/BDGf0/S4o9GBl7/gxf
btyfvhpgjzm2yHvcKH5AUMg1ji7eZhrw2NNsPNcRgxReNeqvqll9unC3cmUV3fNtZuoAFwSmXT4h
q3tCb4s3juUEUtw5XeTJm3tJbtsecJPMRps5Og7zpShah6Ynyw4zcCqnwF5V8oWLoTDZd8j7HKwW
+imf0UWEVIK2/zWJNFJl39inUZxPKzMJApoPz7A1sTnjNq1Zc9Ky3IpBCQS6WU+dShbyi9eMtw+h
0akgUI5l4MAqMrBfd8YrNCesm+AYGR6fVn5Ej9ox1cV6REiZv8HYWjysxZy54SFvXZoQsxKnR342
CIp+w8mkMpublz4RjOA/orNpAaSSw0lr13gyiZOohj73bYvGfKYB1VUmLeGRnOUfnTQo58KlJ1ec
sbFhJRMt7k77tOgSczrjj06NCcshc3waIWDXOOSoHRaSe0kDuTp2zb+MCedOnpQMWrITjPI9HcoD
m+pw5LTY8qBNuqyHGzPA4Bl5GSGoAmU5N3J/VcF9bX0h1RH76dZ/RHuILlwbQay/igPOsLDzzSUP
avywIhRuV4mqc42Um8tjd/8Olh9XXCwTR83zRWNWmQHGUx0h/dGKLH0nOaTI0rS8noQb+weGT4xy
76BREuEzDsCuQVcEFBOosm1lFVBy34cCCc6sYA2aiVBdCj/IaYJ6CsZEkpic5fQeewR+8/Te4f3r
06CTAgaVpSEpejtg5svK9u9lNtO3nksDlrKtXkPeX3UDicf5aijkfOmk2ThmfpZfZy1KJso9ahck
Xl9BAxR4iJVk1dZOO02NyZvvsJpgE7ogNvnkYQWL31baM9yltj2/3jXRxRsteWyLsHQ6oEJjFvkN
h0Sh3G/UmihJY+/e5AphDYPavVoCvjxU9fhw4pUQGiEafXsTT6rxdsRyCO0Es7Fme22LpLjPjQor
l6/rpufF4kH3JFrVraG6cQ7vX8K9y3nEi6M+QC0Y3oGGxNogwuWAYHtSo8PNIDt/YoFNgVLUJvSg
OECqi6rQMt6/CmW7vwuQ7RlFtFcblHnUWHuxCSzlVKR54OvAZ7TcDBGn2nBKgKBZG4P3O1epHPF4
+ATkemCfN//D6lOCyr6hPIm27WSqWThW3qmBuARA/feGuU1EO+cfke0ghWAB15JWh23F+F5yQNza
ipGHn0WyTlxiYRLHcreqqu4JeSPhT88swBri+Lo4ibbxWqwPyPI51THIfo2FA0v++77IjA86xYmk
BX4WWSCAJ/Qx9suGBrWsmoWfVTiEeLtd9s1TvGigTIFYdSiXF8QJ+1DqZCGHO805cJS+Lutkyavh
dkvsbeTRAjmmg2Q3k4IuLKlkTU5lDuRV32nY9VqfzXY/S8MHn8o5/kOC81N8xyL8GKRfUg7v9Pld
V/kSF+YLp+cHDAnZpwQ9waWwbbd+OuBMyipsKA0NjCi3K8752tWbOvmIQ3u6r13nMK0WCGCbpDhD
dEII04Sd7liZM48vuym6oL3q4F3sdGoiwxcYH9Fs8nXeqQ+KEC2OFqVaR8NZ7aSgzIKsHuthAY33
7hG/GocUhOWXE7GcCXDknbeTMAb9YLlAc7KA1gQgW4bdoiHXUHSQzpceJet4mIFadHDmvU7VzTue
c/npatUf/Ri+IVxYMHuxED5wkSxmrogXOYChX+fZcwN/Pv/x7hf6VcFEqdrieJ9a0s0CAM8FUYun
dlrqnhh2TOONK/5qku2MBByvIe+DO43+pYkTnHVUAaEJjEfZ1s7EDyCyaQDeSvN5dJolD6lKBsEj
Xy7bGfBjyIvv2LzBUewkT/4gP67NtBGSykYPXLO/EpqEBZ+YRIOZv8SEj2V5ISjdMAzl34dWR3iZ
H4sb4M6qtTLL0MMvCvyO2HjBT7hBsgFuTqWcFycy2utbNeJb1+Ys2QQj1WOr8OwQ2fiICLcCWaB6
QXWOSOPrAx1YrzTqJU3RnOtVJkYNOmPOIoZd312j/wlHOC9DbRAdOmmFL8c+YuLJ3rS9V5R2jM5B
nYGLJfh3wHyFl6t55GVvtv0jYhWVWyxljkbsLQ100YBkrR+NcZKFS9kE4GeIkbABvLrbW0Q08mlq
H9CXmH/WV7/ecfQj0RXYa22VryQJPsqm+vXDyRzgG915DJVPJbPwyN3TVYsVchC17ywHboa4lyhe
R8F5Sl9DoiEXIC36kGL69qDBe9Ah3Z2KjTq6fXEwsizO+VhhsINBNB1qesMeagh6L7n90MVlymGk
+L/dTLzvfdyhucF6D7jgqLteXqWzCbMADkeExka+l338Ts7Jy1f3D7ps0GGIiJoOqp86jf43qCGq
ttYPeUBs+HlzRxxj2g5jV1oqFLwdgdEWjeadtips6DZu95iR/weUNTlK+AlbUSaVoKpWN4jRsf5/
76g6b8AJ4Dm47EHD33Ck+huj2UEmIdGeuli7T/9WrERFRdl03814guA0eIP5i8ZwWaaSE33D8OSf
cyZIiozAPN7xHcb/+E3ywVYXw6vSPRi3D1CfOoGQNA3sC0/nNslXTA1JNb03n4PvtmB+pYWko3Uz
NW+I4eBk/+QMsudjOO83XOy+C0fsbe/YRZ+jSkC5gxJ9hM9j26kKg4kcdgm6nBiyfqSOcxVFy8PZ
pyiFfsI9Zijz33WPBXsk9XBsTM2WKk4HviDz0lz9ciXek6OnaBq6i5Q4eVtdjArIwIrTTcynvwB0
hxWpCZ3M24PFSsWn+S41ZesnyDB2iTVPY4Aahq66k6EedCjiey59d9I6SMrk9Ckff0PAIbANXgdn
c3S2OJyQwftmS2DzqpWznV4YNnr8isf9i1NpFkR9uwZc5WYWmDwWWkH4RhzvkLMb9CIScdKVW5pW
gEvjBpYiDc4eZVnmBS9Jx9edo9vq1HVuB2oUIduAbt75kdq8JXWmC7bjKpqT0ePtZzcCybJbVOzF
kYTghBSidsci9OtPJdHaOZBbcWU9kvUOrTeEBe5Oc+Qh/g8puqsTbJT9hEbjjjQyYpFS+MrruZPb
JWkoXSGzOS+Nr9H9dprac0q/qnDTQZNFrT7GygCGZ8L0HHfnF632uTl35Tkr9gBtOyqrdcl9TzGQ
tBXxQpjjXBf9wW6MYMntVJRABuOlJBZt6OHkEB5ZG0E5BYDNotW4gTnl9gvYHzZDKlOM/om98DBF
6VfhQ7dS9LfAKan2dTE+E4g/sIiuqoaWXEC6cd7JRpYlIfwDgihqtUyova7V3L3SdmBL77wunkYs
GLjAmtJYZROoWXe9uT9uZdx9PQd9lT8SnQb4Ds2qqAm2YWXU6Kpmzze6RlN6/dPPc0JB/LOQsE+V
PYKZocqheOt+i4tVBDygwDjaH4z/BFCDB7BxCUJ0x7gbSVTBaj6fCIgitPuiIlCYX/ZSerSJk/Fg
+3aiaLldEmbruGdFuZ40RZoC78ZqUmqkNaoUe/prLOaYdpp6P2a/3iSQ87t2DzaBkNMSCg3/m130
JQQJthppH/bgwJmHsx6y/1hcTQHuNnQcFQXAQww4R2OK3yx8wswwgjDAYqBSM4hW8ohNMGwvA4HN
tQgotzJuf3z42AXEvcogoCrp91zxpUOGxAIC4Gh5KTxTgMAwoZLUCOioAcuq9RJHvBGy60QmJ4wM
fGswT+5H0v6c6DXmE35Nq13RSnTokA6texvqrR9gbBS8vGY6l2t0GKjKoZsQsMfTYvII+uf4WVp9
YQ+GDkoqL+eoDXIP+Z/P8VVB+axLuEezGVRL7uWdCh/leCu+RohMzZU8u0JwclvBfV/VFh+zg3nY
aYekEUKnjWf9RTjvEshmCXZOH6y5r206pduqJrXREK9CvmMSVQwCL/uk/KtR8dazKX2VUiGKTRxC
eejkhFZKxYo3Df/4gP6Bp+nh4SFe76OvWijLKWFIV37u1xoSEnLIJGDg3RCxiKKO+rKuKdZ9/5Wp
JkMDLd4Aw45kjf8Jxs32rt/2nC11nMuVDj0sBp0+9XXFhBICsZfUUsXErUOTlUV3uVmDZHSkfRMC
zS/hrwmmevG/3ojQ+FcAVf2UsjEhd/YwnK9PiwPNPVnyt3be1GOvyCvEuqvA8Z3c1ZyHgAyG/c36
PESwrv1hGtAVcNY6W/fz14Os5VDQvFgNUk6oEMv+wQwEIYjVszoQK/pXDXHl3bhLxvRxVPnTMuop
8m6efyQ3oZTiL7QDUGjX90fdye6LDF6U42jfsJpSSxzKSmfRpiFrWMTaUqQWJCEb/1rsVhuAF6jO
1BXsmm5o0DBltApGlfom0YPv9wlYQ0b9mowfyDO62cnkIYretF+A6gnBoKdVJhyF5KMm0Ewzsqqv
P0cwDd3xbTAxjTsIGAoMlyE2BXaYT0KfHnXuGNZc58Oq6vUU+CQc2YdEDEUGYoXHXYIucp83K/A2
MfPuSqP9iaFgMsHzeLKwY6ACXtEw6cliNMvMDYGU3XoJJz669KdlnNfNp7dPAWm71zrPpCnNOPCN
rwe4UGc4INkNg+HLmOGGKShh82DnU3N5TFuZ3TpMRtuUxUFP5FKKUZ3gLvjGkAmqUrbvsiMUzfSj
Olc1tWS+XqBaQXKZ1YIeADRlIMpwK9Ihf6P10NnuUC4ckmwthhTUiUnWRD+vxuSAjy1PJcpg68a0
b1EM1LMX5Mmamd6Qxt7nrNnsr6Dund2leX33LEWklw53yTEU6/LQkmeSTx+3EAUD2YcuZiMNwPps
SQln67S5eOiSeWVQS94MMQ/QhFp4ytG/iz+ukvH/KjmAi6r0nF6e9/HFfmxsqxb2OuDGbICwwfYN
zluLFw8darwzcj7nWdB7abbXzblz9LG7s5HzQ7F66EZbrAk4QISk89QeWaRyMH/mtejgvVJZ1h1q
tiPXzPRjJLUOGsWjsj7uK9Fuslt1noovy8RPt0MM+/UbNQ6X0nlrJkxIt+cR34FkaNUByJCHPR6H
ArXSPmuAKv29jfC5zlXhgaWfyXJMKQO8NC5jLg5QdlDdKUCrzJ/6lgpCo8fnfq6ZEPXP2mA5XgnA
olZCmpawyE2cu9bIgnaAdwkaDxJLr0vimLwgdcifQZHINlDCX+W+H715xQ8Tu8g7lmCSeXikbxQ7
B9Ts8lBLqEeqE7ptcFxvxZ69tBV27ayL/WS4XKjLkBpdgM92XrrE+smGwy6+r3VcEXLL9q5FrYnY
QcxLn5mcWsCGRYOE8G5VVv9pgqkq67uyD4X8InTX359DSWpbIyEUC1rzfceX3fYyfEnCE0uDl0eK
G1Ip/sOlWFLHS3EJO+le562g7HH+gXZJC8T9WwqeDYfY1sfCrYHXeQqKoM4c0OnggCxNUc6yVMvp
dU+GWj7B67Q86P8MFjkSFDB9cCT55sCKlZmJOiw/I2+F75nGtqQHANwSwdCwqwPt8Pc3qq2BDupT
A8Fg1CjjWTUlTD6VYuhKL+R2r1ya4MJ7DKftwHoQNfFTqyoLtZ5WuY2tpn7kLz6s1pYDJPGh8G2p
OhJvCIMgO3gxk8fhiAK5XB+k6WWTwXhSqosHBN/MuWf1yi7olL+3eLiJhLfg6qn8WFC4raBJlz8l
2tLMw5EnxTgpN4U2LYENnou6LTkR5gOx2CIzoitO0hFyQqYEjHRZkMPjWlUwZ/DcVmCza4h53cxg
llxq7YtVqXNwK/THJV6CZrhq9qRqLCTb74tA70C6mVh5lMc3dZ0tFP+ZAT5NLntjHg/ZtuzdzjGC
DiU8E8ZfgblzkAbqqjjpHFaZIh9TBhrZJzT8YGQ6gnJgTZnZmmNq8zGScfqWmt/6EmANLxedIgeE
N8x8NQIx+mRvnjF6iN0gWUUPxLoLzAjSti+l2HCcvTInHRH5CD7BoQc4OHqFkPjmCUueASa62uzj
si0ggJVm41iBL9XQzC7wZUO2gsVxUYxy0Zu9ClslKkpgO42sHRh1ouKY03RjNbD/0mUa0PJ3jP2L
ZTFyGxN8kHHuDoivyejAF5E/PXvLOUso60pnkA0gCWhaSlT5Imn2S679MDHFAL6IUvobwYwacfwZ
nEuoBVc+5r0x0Zwp1QrK/jYK461Panx5dzesut7Ulow5BiCSYy0mQlmuSmTLXgw7pPyAqSv5f0Pk
5/uJgSpweEvbAplnQ4EYuvzDJ7kDMGHkBPz2Z5kgD7hYpvZxUPKxJQDM0P7UIlCtldhpUTwaQJB3
XelCZfXFvSIl2BYBi1XRnVX5vx9jCSmjy3h7YN7pK4FSJOYHboPEpWE509HZ++p1mILJ5jQAWK4I
1UQ91YoJIgPEcvRGrk9ZNH5wRrLo8Fq0ywdMnhoaX6ng5uvAxGBVPKYrkNug2xxoP33gm2x10LDt
7QtMxVdMX7RA/9T4wstO6hmJszMGD9ff3y/vstr4mqeyslXJd0cazVDJFgsMzTjXjQVARnkR1M++
usKq7NyZu5hCHb8rKSGqMKk6/HOge7x+gdDS0bGsvAmuHbhx069GuX3FI2XliiLlnWfvTNTxbdzv
jZly05F36MX1hYOmXtnDMEvEFQ7MQACjM5tbBgOoAZtlKWX3qH7R373Oa7J10dgxDXdKSj+JC8a0
+g+ojmMyuGNVAsvdS8ZvNuuG3JJ4KuV7D2y+yZbQrlvbJ/adDMrk5ZSzVbIJU1FXFGAWK3KpgBkJ
XC7tmy+2XBDnbLxQQeC48+rpDOYj5gb16BTQGvlUcFhPau580pHGf/7VSmTJUPNGFWJhssISGEOo
N0ahB9NhaUghSW3Jk9QOiaFe1eusInbp+F/QveGuBUvtWjaTtv42hNOAfoXaNgZig1+KHMGb2Y7R
rW9b2QzUjNcqE0dQpO4mhWQRJ9NL2m25zLhE/4BmMe7hwCpkAycdo74WGEKE/fPA2jlRsOektufK
f6xH7p41Kt/Ffs8Iu6Bdh8lRnjaCduOYgkwLOMbE8WXrNg/p6upzXP7yqvkm2sXwRIZLmxwGT8Re
WN+moS7tkBCZfikFAsWqQLPFHRX/jfT4iO+fQa0LmbSREYMGt3x01XP3QpxFDP0lMNltx5WmKWoI
q0D7BbxSdxFLeyS8yhT4I76oDznRvdqc61AuOekpA8nImrvzOFtifo8l5n45yGfATsT3cS9ZlnVP
KgwDIH6u637dc8VHXE++XoczuhDSEeX+4zkaS+bRPVW8LXXV7OjcT2tMxEPKhUWtMj6yWplWrD0P
0KfAZh0Xyr29d7Pdld1wuEP9DXIOoRaDhnUtfDpsWg+NDrUfqnJh7dU80JIIoJSdUB4vKfG3U+F+
p/HNzPW/j+uX/b6O3p+rH4HJwDBl/fpfOkBseCOAbY/e1K6cfDSNmu0vXS4FLZR2YiX0xk0FcFtp
YN1CNuwADVqLtgGQmndWMXNzRPEMUUAmQ9yXxFSFGwALehiG2Nd37YeOrdrjvlQ6kejPUFJkeSRb
yjB7A3U7lKXt43aDh0c1ktTVIMR8TeONXNo1+8+5IK5FySLyYMFgdn5Z8rgERiO/f9lKLCbynTu8
nOH4ehv+3WQoZ3yuQk4dBWIW18EycNQdRgLTiaqy49pM5Tgh+jtbbuvqTF/L6a1fnvg+teIIttU2
VDzAViUTaiZKdLikHo/43ktmpoMdfVsZrgQm6q9kp3/Nw6QUU23n11RhfSqmAX4oSi7piOnHp6Ya
/Qx++KuMBPpYDLNgHLKmx5sRCx2w1MbGbcU/ofuuNWTEGCjJ59Ycoozm7F9lfllyvaPYEUVvN/ru
zjt/bIWGrYn0LGl9DZ7O0nb6DM0WN68s62czTkOY0lAm9nxewcYUKyHiCBxdfUCPaeLnt3xFremp
sLbxGsvhbkOUsPZUcNIUAVqJrQvmZRtuvYGo55wkdqfw36gN7yXcVUaNPNcIfWnFdld366bpJO+D
vzQRNywzjDpNiwnZPwj2YkqO62KfWLgKphOVAgUtxZYkU2Jg52MnCOvMrF+GTMsX3EDi1kNePGL6
gyx8zWakzZ+Ee1TmaRU2ZZIuHlzZrXT2OC0ESY+AQE12GJgtAzyXi3bissah6lTyZGM8S0o6hBmr
vIoTgpgEE3AljJk9fUog/ffp/3Famw2FdXVhhPLlcVTYV0UQ3a4lBDibET8aRDWWU1CtvXczeQ77
TVjw+R1TW4j5AnCGzC7IDG6nD2ykoILlz3cXJ/CzHXsW9lOhMzJLv6xYBaAkLxPhneq4YK5wWoJt
IQ9hp1xnnRDqW/KeP7OL4nJCNcaTeEqNg6e8pyV4nj91D27/KzXuwA6ha8+GxaD4DKZytYhb8rWu
kAU2VBiAV9gXmcUP0ekYjCaWCQ07C6Lce44KpCLnjOKnS5f5B1j1WKKRU0x4o/g/U1nt/muSkSid
7zwpUy0ZkU71Zh31qZYsuHc/INcC/5z+AqdPfft43buhSEiRKOW+pKBlO+32ISCJ8IN+YuaTJqZe
NTfY7BPOsRQlf8G/OP4DcnowXiU25MF0e6epfDt4RATsiPmqdSGmKedcWokS7gl/M52/r+agE00v
ksGc0M6VKnELvaDU15ZB2H2kHGX/hafjCk0VBPBl5fWIl6VwWQHwomKaAWZWFFcrQk+RjXYVkoj3
MYl7rh9gfs4v3Qi03PBztp0R8mwGmFk9b2qzSne7qmLdiyyFbDtQdtsCNsfOV7QkTWfc95kDow6k
TGZyu7sobqJh9O4+sI2rPDiH6fBQQvs2P5F1DjUETiwe+rno4uOwcqNUi8TziR6jlcaFywqXohLG
vF7r/x/STpiEkiU2if9/hTA/Fr6BQL2Pt2JH/n4mFWIWgeBHXYlJKzr2jbQkFqJe6D+xjnee9qhf
yQHiNyP/AC6Y6Lv1nm5cycuTNWR8zrtyEKUWp75yEUJExaC/jCHgey1a1tFsGRTTB0ozlCvSKxvi
nMUrRrE4SjyUKGPfitjkxduG3foZgyMj/mdmLOsLi5kBd5Jdk7EiAPOpdkzDEQSVJLeLQ5G9PI/G
l3iPdloXy2Qo0M2pRtCgx4Lk8QdX+V63UHU0R1DnV05xKjjTYk2NrJBZYsd5YOqXs71BTz71p1vl
d83M5WDkgRvxs4EJAfjOdyOfahSYeLXKvFZ4UJAcSuGhqR2fMm+vjNChUPNeIUpguUsAyVfJCMZX
tHv996B77+6sziPDk2qITKAVg9Kz24bFsiWLFJTHRJG05xanbHpQaut4l0rVnBez3dSJW7FRRfva
QmFlEzZb8hFL7FaZ2vU/eUfRFT4lHP4VTCk5FYak2U1J90l7+AQN2Lumj+P28ZI/csziuKN42mcY
lbr9X2Or4zJ4l105cxyBzODAuAFbC5yOZnwqdPfcEwVxF6f34TRKlStJQ2OM5O7aPSe2J5dn4kA9
L1cwU8nWWUqSruIbK0qQ5syUUZYKIxJenEDSkQUnVYz7P4lKPzaqOtiI3Q+DFWDQuj4465JKvLOR
P7Am8pdWyZNM5pA6ICA/+AoiKaJEqd2luBUCJa+N8+iDtMyBCXqUR4oCYy5sqtNWmZIsANGDuEkt
aD79OCN2jDpaz04XbGKKs2BuCbMP0BBco5R2hqmLULZYr1yL6PyzQi6NoYNaAr2soaAmQbz9jdGT
8dG9YWJEDNoE2j0xaO9GQxBNG3Yug0LXxlT2MKczuxJqv2uuQQWnpFFRynSyJiNqh5sZ0/9XyaUF
PYeroX6ZjJqhDMavnJ5GOcKoEC2MYd6gOuTXFTrFdkBNAo57O7wXbjsskisnKJcTJLyG3Jk9QkvE
/TulEoMyKOgAWuEWKx0M+zsU1MaHXK1/ERqi14QD2Liu5J14PUlihOT7poSjQb2jqeKls0EWjOd1
HQVcLDK3nyM2OwXL/DLgNsj5q6wpOLGI9xexiUa/ND98BwypmZDA1VZG/s/XgHBA5dHmbUGqF/fq
WoIDx8Wp9cDa7TRGQmErJy+Vc38r+C0A5jryYyXTRoXOVhHCITpjpLDiT2LLguuETnmjRwDzPpgp
pPkO9tnH1mCFGbI6uav3fmMXV4d/I52u15NOhOjQP+Nxw4EiCu0vJhzGZ66ECQgmSKaf9wj1zqod
v5UxyPw+IR1ymFA8Nw1RV2ZEbSbY1nD7u5yyElZike/xK/AgxFkrxp6RGwVx9aUKbm/14BLdCY+0
YUiY3HKo+YHc+qIi+EjM0i5dO8lNgdQXkGJwTZHuDFUCsWaGHJu17LD8tL61rSI7mVin7XyZyXMn
JxIHnSgQmFdyS0jXcjKZe078BTF6Q7B/c4FrkL2VNKY3uk0cOr7hDzfb6is0HgwgUVQkJ549aWVW
9OpXVBhHzjvBzz/N5TuKBYRn3Kg97+nPX5IF70PvPnya6/OYpf+RK8hbMcDi7JzQ+8e3f6odfHHg
SSNjPVukPIP7D9qjEw771nlmtmzpO1QXReWlM3DyCRrCPSq82DjSlCGmNbWQnI5UXPQrzSCI5S4R
cmen5owEYMffagzRxiitM4sfTc+ZMxPA8t9RduQNgQOkWvQaCZOSc18u6NDGs6KEKKZv0lB5Om3y
grxpYuAmMAGI9dco8gsimEFkmGgELfQMpzvw0uj5SbUjTDo1zON7EuDFHX1NZdLAyxJ3BHKun3Re
c3+vqNdE9MT+psgJhYWeQplfkv+ZQU6gHQ7HYlxVK5vuNIoakPNyLJdCjMGCzK/XOOfPYIOqL1Wp
Jrqu7yTIs3D+EUlx1K5tsQumCwfSvax0nchQSaVKTJzPU6DkivWqx93Z1m/rRvw23bS7BMq6icsa
1tQQkY+xxCKWFgSD4PfHOAAgtolccdGUWGPjnWfDW/eslRILOxRhg5TOV8OoJGO32auJ7wczxmG2
yID75pw8QIOEjc2IOnq+pbfNnzfQRW8qXdYcX27nqKquAYEK7noLYEW54lp+4dFOoLkzwxFk2rHb
8uobg7XTa/R2DS1zjZwur7NqnwRSqjLiHKfGMZ1zY1TUpR7bEoAW7S6dj0JWs7WlLFr8ui2O+hin
8dKcQH8D9tB9+H04zHDF/FiGQI6Tfd4RWEuVYUeBXLanS2VMyTtH0HEPo5nxu8n4EXs70sa3OILv
Mt0HQX3VPV/KGdp32dyUxHh7F1zwSNWSErhQt/EyJhaVBAR6JM9EQG50ntFbMQXAXllswETe+CMz
B9cp6Fz23okBWD9dDz10LZ4IjIR1JZKGBWLFzJM1hqP0Kv0sI7AOphH31Cfid/Ss/v3qMFbyvOoH
+10xe2dHnAq0JdWWldvfv2yS1zTf0g6r5QShfrQZELBIg27T3Nci+tfhtpfETbMyHvS1+/wDptOv
c0XoLg1t+tzt1uVSe5fl0568mboG85lxVEdrHdX3wMzEpNHzGjhDn9IoR35Wre4CapNlxAEWlOhP
KPkLiB7IfpGFqpHahCfU+YoR6MAgSQU6EJhKT80DWXJhVEOTCjwC7aj2KeNjoTtx5igGL2OkWyT6
yjcmgxbOFoBtynbFNc9QN8qGQV+K5zU4bAFPgyPh6F3JeIH2Ot63qlfCTjvsz/rOsmDG1bJJuCs7
pcHmM6X4ZeZP3JXs+lqwcmwm3lK0/YgG5PMdErlLBjghw0h1hP/mpq1DJZVuOZdCR8SDyhXtjx2C
xe6hedBjxZsEmzDXiZlI3vUg5pi+fBVGhXZZGXfyZ3URRHV/LFmJvZAM+pH0fzOseDUoWMQ6aQMM
Lts8QDwXlq3SlD5I7BL0b2hm2vqBgbOaf3xqbf82uzc0jt3GwSm7ebZLl9VBk9hgdaxyjKczpjdu
mh+zqk3aCPu1oJNJcwBOPAJQbMAlMgtCbHo0XVg7h2hBTUjmMgfbAVoncm4orwbMZ0kBvgdlgP5T
XgBBX0Ud5Jut64zin4jfVv0DTMTnM8lSwIGuRO/U7zXziF7NSEIDkpJz47ViRvIkJEzlCyoz/FIz
6yjUOw+oL7twudGu+mPWibijfbgn3rSiD1Yh95Eqd0oMK4zpXP3ssOkvayMX/O1qQ4MvK/laL59/
lurzsduenliQjzNSvHqvMTfy6vVrZA4abovnxcHnHmD6ao2IezU6D+jUgVsrz3RJj8mlyY4VQam6
Yt0s3OEvnXoN9hb0xHPBaTcWNc4NbuiiJxNHEyGkcTSrZzZVx/NCXahAA2ps5s/asv6nPtF13m8B
iQcBHVa5CnORyX+0xeQ0oEjwvsRWo/IPwFgIWrduM3UPtu4sHwtoiC8J2B6VzamYh27bvHQSomlQ
3CYnkGHSHvrV4P+QCT2EDqkIcsr2YMrKQV82nZz4xkkz6bHj4lg+FauDJNp1efMzK4xZZyMe6G/B
5uybAJzRZSF9nVKYPK/5tXw5XuPb6utVdGwSzJxoiRx87iJxf8Z3/rza2qpXlTzH5Vo7ztDw6j3+
l/lhvxqJnGTG+6SXT9Mp7bc7+doxWP4qlL/i1bgyQDUHJ3KbtLBFKTEvIbU2Conb5iI1xSEliAl7
+UYNnUQnNDGm3azXUQK8O0NX1YaQwNQHm9rSi6kq5a5Zbb0S5WmhUoYPIY1H3h/s8o/YLQeg4Z/w
20LRiFfjteVZIDt6A9VIawigdsPW9wsUtFV0TNOI41QvgFyyObPbco0c0tbZJmh+SRoPYpFYy45I
F5I9t8lr4Q30V/9+9akdDCTrRavPqYhr9cpTNWr0hslBXyDdoGrKpYX+nQnuvYMaLww65o3/cYTD
R40Zk7z4EcgcI2bNTEOKkqXs9yLhaKB/2BAO17g0Qq4HWRvi/HgiLV/DRtnLabW531/MNsJ+LXNf
g0nxrmrVjaSFQdcjMjrqjlYrEZPUAXvfEPOoALwrFskFkqASpW8pRjLM5oJMunffVkbr7vhzJhaE
zO5rxeDGLkWdj8H2386d2oqrj097Pb89+1yfri5Xis6v5yPa/utxcSzSinA0r6nA2slQuhIk4rHZ
bb5Z6jtB5Vo63q0DduP8IXIrkKwCnZGR/thkq2PDbRG1FZXQotx6V0BKWsanejT5uWajkdtcNMER
ARb9bj7RYDinPy2RmSI44ENJjizBbhHBQZQyfXZOaS6G9A8jDXb8yQ9hRMZePxNNVSDwckuhG0R9
vkkCcP7eB6Q18Pwuc/PEpjS8qndSPBqtVxloFdU36k0sOwB3av6vdnmvug3T/0ZfUN3b9N5mZgIy
+5ztYRP/coC4nfTFl1g6JU10R94npnn2x7N5N7U/k3fARiY8mHaHH1SEs31Mn0eaaobdEPUwTVSl
DrRpZg/1m/5VHWiYWawK3fycrGjonIzh/T7wviATeA5mzi/+4xzRdzpTVdVn/jXF/98+y8Ka2z0F
skInK95MApFaPeLKagKUtss3PN83t8XLkSUDaRGFZyZTsMQoQzowIaJIvSTySh+Rthy0nXQyYaB+
lgyx956Vb8SW36TRUvOyvy624UX3l4cCcuoKhkhx2pvXjoJK3c4eI7g1mAUwyJnt1TmJFEozPGzT
ibgfx0Svg/q2WTB33xk5NtsLZRFbMOFBrf3nbGMd6tVgQG9JiP8i+r/vr4GbLrFIzHmj67rKnUaE
yxUuFha42UjNIERucNw1YsN4XDJO91xW+rZt6b+HZVrsFh3drrhcNDQDCYXDANAAKMQcklnrqkGa
TUHVXPnrwD0Sx2x07wAS5H50xDD1+QCYEgZbqUG1I2FyCdqnah1+vfKVKPWxVl+9jjLEG8+B4NBf
M7vi+/PY+qexiYUCh3UE6ynjEWnOsMcf6RPWG08TOaSmn5y4uj9SAFLuZAjs36uOMZl72tTBgy9o
ZYW91QEbqAp9KqQUg3dw0DLHu/WIyYcSi/xulgCcwv8jpPBWTxiE++zXvIE+syoRPWec7txCQfvB
gn9S8mPSHkGwH1rdroaX9BumqqyAZBJkBmqpoalTpY/1g/wbB20zYtQ5pN/y18N6ZyJLHgeeAi7Z
smAiTqH8sx5Ax4xP1i7nCZJM9poJVtkj4ssw2QRH9eCggK7us9EHEgAkO2XbiqfEs3YIHSEYYLzY
e1awgA0ekVcXsHWbiFoWXhrQMKOtaDa+5PvyQwATpNgDLFnuYGT+SB7JrPCKnNnIb0GXVYtIDRZT
CSaGGTxHGRK9K/foYZIk4CWGAkmw+v9nzjDZQJwcXyBS00dhlQ7a5RiQA8PmhBk5uq8We2Hv8G7a
Fs9iSCONqfJwLWBqGqNRgg2xI5Eo4iKcQ9Sfq+sLdBHsF8AEzg+Nx5urpAR7SupOAjGq7OZnQs6W
vtQRxcSVpAcJH4FHmbShvS0qM8nqH5zXeIckg+CqVAOi5f68BC1WrndXdMjBErZWJHR6h9Nqkldj
MwxV2xqOh+NCiatbhPAfD+Na9wODGd67KKxYKFwspo+4BNQ0DmM3vHQVM51v4D68U4yxCIuFXH9/
VdHF8lDUBmz95g+Zb7L36vah6VI0dPNl0UkYfcUuS8oravOOc19JTrzJJvrajqiWCVhLzw+VMf0g
1bdPGFwC+bcQL8SqXulNZJ9SgoeRzdw+lohgz7pvMqIQCKFkGfDgJvuA1A8x76QH3SJDwoCM5+5A
HUhDfQiNYphvIXoW1lZY1D0wn5pGMtyw/ZcYuUZHNB0nQ/UO7RPVwFCu4G0qGuEOsfk1Xj7BUMzJ
udtDna94ql6YYQa16Z9z3c3A9ZljDWhc6A42892cBiTPOUos48VFANdKsFuk+UZvxAuafX6WgtB/
yyIr6j28LYMSjSESrX652umo19IUPyGv8FLVlAKxpyz32C1GzwFBQ5ZrXnnrUWdsIjpmFvetQEtr
FhfsOMa7eKfJflLrMkqTr3LsOuJxIhArw+Fh2xa29clk8Ei9NR6rRNQVcD7TNX7wEWgRE6vQ1MyY
DIQQ6gh6R6fNoGyFO9lB2Y12850P+dnEgehKwmEg0xGPg2FOZMZofXJk1o8UcYBJY5vu43QnUj93
/BIWPTy2jSDJCUM8YakbMLLXwi3RkjXUMtDYsyCMLh2Odomrn4rVP+lA7T8ysdxreiWCdX+F3mo3
LCbMEaIIUK3IC1WqsyPkopzjTmOnDrHoslBu1LellJCQ9UcABAe8Gh1Ngfum2nO8leEvS4TlV1qY
E07KvsdfQJZnQGCpQP9nhJXTbzncEexYsQUWCoaX6kZJdMjFxnuM+81YSwwEZ4icovmDUuCmIqoH
yP53AbGoBTm8UQv035+tVVGsqRB7Res68X0d86SU737laKdtR9PreKXmZr1s1guc4m9Ude/pKI1h
tgk7qKSngRnJC7QywOsOAc3stXgqZ9lGc363sETLwxQfmHULabM9uwrRRiqyMtkBFp0XvU5pVcMT
7OBDQuuqc01J49zjBEPxIXulB0o5s5D8vTqXWfZOAqktKAwS+KPynoin1pUOan87Zn55ra52S0pB
H66QaF3nUdU0h3pHrdRL2qHhBtip/1/d35yUYryY5hn0jmfrAWn1aUWgWHD+CDgI/oOFNQL/kFl1
nQymXV+gdA4++qt/aQhbEcK3vgYiByeRbeUycOSmr8DVQ78NDgkDOf//BYiSFbgkBwYd8HEGIM9z
qGD3aOitv0EXeUcxaVNXJB5MlktLKSb6IgERoEbafVtqa+tMTddHFhxNHUKWWup8QxOzxxaFTGFd
GmmsWQU7eefWTkz+P5G7iCN5yd7PC2D+tAUhTw/pLhMzT+GaXj4QKkxtjFjGQBBkAu34PLY/1NHn
z9zkLlfAZOYxdXEXB2pTL2aGOi1lbids3WWZYEHeAcYIEBaNCeCr+IxIgtPh1NuOiQl+MRbw6pB/
qyOheTFd047vlD++U02A68MmZ42AGybh33sn4Kq+D95s5fWAYWsD6GXlHWrv5REr/ZAV4g1LUSsH
W0kfyQrvsJsRp7+uauCxN1Kn+fqnGLGA6uHmZUuE2MQR3fl550M62uWWTI42WWvjTig98RZqPovq
BCKEGIK9We8wQinJubmZ9+UiHs+Xl/YJCBNobp3kgdNVgSOC2BSltN5DsakBg25XbjWszZoWXoER
jyu4NhtUtJUaHgGLMHv8cLsWWcX9u3R8CIitOchDubyX6Cuv7KWiOWuBuR19OATsJqqNlWZkIFnT
8WbMewb8Ck0gNnxrBhH3oOV0/ziV0EubC0NIHv2+dguu1Yw9SKA2ZPnjY/6r0CZkmZh3zPHHSC9Z
giU0gt3gSB2IfSGyU8KnJLiO9Rev0yHOkywlihTl63tRehTQIehpyL7ghzyY4S6WBURjx6p48YJv
AexAtsqZtVe9cUk6yVyvk8k12weWIshvz3xBJlvBCB5hfooRPOovrVqvo/yn31E4l/JZrARF/EcP
UdPldXUVFaxQOoeLlOLdw3y9uhYGekYE9Z3gVRiN9ydvGWCex4c+GlZvc0yQvzFdQKJzFBscgJ74
vDAjFdcO4dwEZry8ZqEv6z7W+FjRXdH1faw+Bl24PYCGu2fFs9bbwsTJwXRyboGHybp8WoyDvNrc
/Pex5ueE6Xc/cerIpSb43ZRlHvVigirTDfpj1i9qRkS0L4ydospGocWX5mOiEZs3Db0u5TXkfXYI
vnjncXIg1DJRdxFY9tmVTEdN3kIvF0hUQXeVWTxvw/Owy0Av5TF1Hp42ovKTZ94GQeFovVwmhkii
hc+Nr1NFxGdKlFTI3v5jsDHDyPMbQtZmkeoHSRhVg3lsLdol6A4n4XTeuGv6pEk6Qp51ot5xZAlf
duhSAlnBgciiJCzB81y2i7ntWnOFikutd57UGwhcCp0KieRnUjeyvawODKV9+8uynhCAWW2Hcgf5
Y6mQqXrUkeLkFKrAGBSPTvyBdgOw+J5pKcolP7Qb3+O0CPBCrxriIVNOd6HE0auz2F2JIQNIgFvc
ilprkXlem3YCDw9mKz/X9O0NlBYr4rPmiQvsoS467rU61n1xN10lMRQ53N7svOZWNcjRXj5VFOO7
C70M1S7VXHisg0ulBQvyMK/Y3F0wfpyQ34fB9gM5Z8DRdhw14Sn1OJ7mL2MTB1AnO9cnLBl50Gd7
6WNAUR57YRO3NG5iYf/fkWP/NSA9E68FIG33pmB8GVWSIuLRC6hQZIy8K9S/dnfjaTF/N2A7qjc1
IMTUX/q6nENoxKW/RVpTLL9GNAl9XcR5iljrGuscFqgW4U/KjlNacU+qAdAkat8lUkvb6upN1r76
hrf+stn1epDkJZTdez3w5US/sop2XBlZTD5Rf0NGe5HgYLzdnv+SVyx29LAPTykWUUF73sSOfARz
rD0nz051ziipgH0XVwTca9UCCtNEDcUoa+GTw7Jk7Mbyc5zwx95KiNyhHafjtMPwvdL8Rjk2Ldme
JBYeOO+XeYqVVk1ztW632HXaOa5gVps0KOm+k9OJTdVw2LB8Rpy/rruzZSapMRqia312tCNNEgiq
PcIewf9LAv8MTE4R9prmIGSzer9M30lucsIwEq1e4Mz7oIAaPwOOF6dwz3fVLc6Uknc5uDvoEqrm
ReJrWwy0J8eZtSZVivBKnKQkpKYgk6LUrmwluUJhH22w+S7MQTnbDJV6tlYn8CZJ3Wtnwm+vu6Im
NpBCtWyI+PzWf8v65LKukrf9iUdpIjhitafqUH90E9LiZ/SAMbQsUx52HcS9xNpbqS2H9ucwHKAe
WM0jJS7hIrAXTaAU0L29/9CsG353dkEb/ZqiQd47nbmngJWtKBFlh8bKs2bmIuQoQB/H3aGJNl8j
7eWUHN6mxWnLvoQyNwHIBS2Y1GO1Zch3jlqBOe7X/l4To1cCZ/VV1Tvj3Xtuv/FYA/dxjgjRS78z
L1ewJrLbn5hjx3CoBJvkKfnBEnWCQh1ehPhIbgQKPLYdFpPXGtHriJRNg3Ih8GdopPR97s4pUm9O
XMAqsHV3PyMqksyqfQRAN6dVut5ykwnpGLnKHaTheL4XrzHVJWLRGCY836HXhrzTA95N3jGBJR4k
DvMCtJTy0jDcReYi9UC6XTo74FOh6pqZqvf2Ogd0Nafkp06o+qLcYkfwrmprBZ1Vt7u/Thmrsspz
6vIPuiRK4ljOXkd9vsTGvBwBk+SflMP6r0xzg04wSUg4l04zcoy1bLxY1KH/oEzmzMsiF0U8HQtO
m5FTT92dbKQCu1i1YAhlFTKctvBfaYUPdxGNXQq1nb91twYnGbyEXTyGMpL4//+YBm7hyNVTh+8b
IcHdHXFjjB3xkPaJZfGp+ejkWUU2fyF43qzyAGaStfES2iH2YAR/6y0BATGx8NT0ZQHb2iGz6af9
D6BcTADRiVX9xPvodU3qhwyB0CtBVX6gRaMptuLz/cUzO3HtyCKYNm1H2I4FIVu8uYuS8v268v2X
tn12mx3ztGnXR6juokJGgm+kWLLecnUNrj/qFt2BHz6t/zvdjq9DhNY52xz1q9YedD3I0C0QZg5S
mJvcUkjmE4twi8Xbu4FN1NoyUxW0AvHHYru+57ZRoJQA2xcpD38MqZiyfu/2M0CHzBNWCX0cy2/s
Dvzraw8NnRxqBBojEn2xwE/ta9cEbNxHZ0F601+rgZSf4PshddYb9mM1vqvEszfVELZIP1XwWOxp
S8wzU6Wufa7fTh/O1scbCd5PVWn0hI+FLMAhy/EkCGvazl7I40isvpsnR3NccNFyOzvf8R4zh2RU
LpC7Qp9adna7SV2d+In5a9YhhxoORNRS99PWhEGvCXRrmJiHaRiZiMYZCKNK5DlgZuY0U7QnfXR2
ep+v3J1GkIWyf7jE7RIQcrgW+BAosDm8x0Qvj6QrhNABJ1HZq6dNlsZeL9Gb1PLJlyC2N+9Spvvw
xN35zjL093be/I5Fv32dEOSPvUEfrAaQU6tJ5slvdjf0cVYwz358WJagxl8tIfOcwO0/7oMwG2+6
ZxX2/hkL9k4vCinQZUB9yoy+1aoQ/wpZPchclCQbqxMjeJ/sA6p1LGPqc2yfrdE7ICccW4BJkqoH
ycInb48yQ/bJRx26yi4WNEYAlF/U6gwwWSVjnWle5B+scYwShL7bLOQCR11luBxaSRu7AQKZ5lFj
/XlE0EaWx46oAPCnxLtiMo1+Jthj4M0mAHYZdet1qxdjB93URuKc4cp4kGG+R89ALKSKeImvGrWn
9oN+xX2SA2aw8lz4wL9AKHyeVmMFqxIVChYcqVI/V2LjRPzebgQ9oD3Xo2JWe5B+Uh/pQ6RtwYzF
WMPsu+byHmMEeeFSfMXc3+OskE50AuNj52/G9esZwKp7q9pLVXcrFEkbf2DuQk5yiavFruL4HSSX
VBzOU3ju3dMBGLa/gmssRR3o00Nm2rEsv0E4PuGGiS4aWSzF2qW8ArlRgdwH0Sl0LPWmpLI2Xoh6
mzFOqkTgxdS/VNumIgPywFF7cylpkA9jI57fFFATfswQskjselt9nKQ2msU+60Zre9LzgZ2oRgUQ
UkS3JdEkSnnGyAdkgc17783BzeZ33DiGuu7eRIPc7AgSmP5b8Zn+fcsYNnAmMgzONzrk/I700r2o
ffneNRXz5dVSjUkB9pEnLNrJ437mYKotg3Zssy88CXWHuZJzYoRt/SQibHmKV4FBUFbB8zs5S2N0
QEjgdhJZ82cGUu2n4QVxYbC4SFKx8fiOtuQDnBSLeDu80Rinw/tw4mk97PMNY32ADrcWCKOza2KF
VqiDU+A5Ly1UISZHUUkTotB9I7oJ9SoomV08+WD/OmIKTLZzf5XXCCkw3e+CoF3hww9lzsiV/Y3Y
P3ObthruFPJ4ESyMOlci9z9ToQp9Fym5De/8rrnscgPCnHsYyfIg6kBPkfcUMbPedvvNAQURjTK9
HMll5gmvRiii36VC+dl0qCfoOBfX3VU98TutTMK6rFxCR/DXA4mK5RhX47QRFTiUkmEE0Fz8yh8j
FsElrdW2SSc+cULUH/Q1lobh24Qugi8MLjJihfR1V48Eirn6DfLLF7P8cw0ZKZxWs5ON0H1gilkK
maHF2EmbczI4QyXR+z9b67zQsJX/NCAZcmazoN5IdQQGRBWl475KwtSeUo8Ivz+La12D1lXT2wDN
vISgT3/XwH9W/5r3NxzqSjocidkEeueiGzMX/o/G4Ng1k9MWq7+Dt3PxUZR60IXUk/VWIb7kRiWt
jArs1H4sDEwLaPR9xunh3NdytlZPEj10nmGCeD3zlCR0L/kLDr1jlF3N92LRvE7QVLbWQcn+L/KF
nvDLYnJjmhm/7o7y4qS74NCDaIFCwDOuPjleMXJr13J6a7JzVJykEKGXWKZJs6Gb5tQQnino14uI
jkp89012io60VPEcErZfebU4DRhrB5BG9gPyfwCciDL7KODl0QEwBFOU14Sf3o7BK6IEYGzcV/9c
CrAvaniTraGiW8MYZwDCpWq/Isg7qple7eBUdJwgVfbbOd9mvXCOy1zlSqfg2IPtEKCyG6C7Gh6d
9Z8luAIR9cRJSOfKXA0UbG3M6nzHHHiQPEdspZJtwtaJ88I6AGu2ehf9YOjd8lYBtXo7PmGbMiVk
2w575CC0Zhel4diQeU8HHJi7Y8ej4GPBbIB1d6lif7GToiEucD+HjkTWn/E5zVl9HmQYkybGFuNa
rkGnDfZGdRmOVuXit+cl3ac5UChcqpIy17PMImhHgPhade4wbDJSGi4yqiDgDB5eXwE6jOoJMlrN
PTQDE1Jh6FVZ2XMfooLiARygNoPwR+6MNt38xVHeEwHXiT+/dU5vlmgjap2DFeqVC9v9hqWINIRT
+tTWylITCLTAp4/ubdwM7uaiogkxSb0aghdKNptEF3kPsgAHODxn+TGlbRf1e7mz6i0Tu1mKEjQ4
AxqUSO+Lh87QOJ4KrIpCs16cBYaYmNA7WxCJ56HO2mr06Oa04oFEQtTjOJud5wdShqss26lLngcn
HprW/z54OKXRgaPZO2O482Qf/AGymfmg9CywG37WIY3HqLtMFwmcO8oJwhuOIpAAAO4+m7wRPdAE
3zpoIlLcwMPG6zqDW5Qjq2+Johx2GfZy6NqyHBxGcozQYT385WF+BmfNR7bwVQClcr+w3qafB80u
hOsaOHkHuDLAfSMQggsW6lehiv/NIHGOdC8yd2DYVQBOzO5KH3KkptzW7X0PnRFh/+pM4N0V/VWS
c/PE9ySvS3+N/SSsKZCTCheHUqjexHR4KTaMzyDgq9XK1HzcXS6epBM+MQy+2ctmhUh7cD7dLDhV
eOeQ6q19m4tSQ/oH7nX96SDXPrwHMJtE0TZKNWANfQ66K+PdydXvVWgm9plEr/AR1dF7fBHFHg/G
EaXamxvf4UxpybENk2zQ6ElbwwpZMWMr4EDgFt/tjmJ3B6MmmBJBybDrgBfgMWCHgCTc/XNAAa5Q
RCrRdx9GHTd8lgoje7x1WGXNXMKeB9apLKcFlFwTUeluYj56Q+pG8TzG5AFdfx2QNT6ff4VKsTfv
Tp9H64uUfiD8oRdS1y9uZwUZKLLnDncz4IJ7Pof07XyE22Td6u0b5945ToYqsfseqhHMMgqwKIeq
3ub/vn+v6vq8nPup8XQLRhtHMdoIRMkmRVrr8G9GtBblQgEWGFd2ksEzSfLL2pdzyBTLLFuodz36
FZZb0TTVhNPnmOtTIdQyF380+PZKwR5Mk7eF1HALa6tJC6YjFVcxiRKgMP4BiPF6Aq0q/yk5VVlf
tB02YjRMW1MaiVAjbWNtxKo9zE7RscBfyKzwX82/APfgn5yOUkPIzSD5pdDdXNK51fa26O7WByXr
8WYgbJKMgaml9s4yjRIHAB6PwQxT4Eg5wbhk3GUff8jyXEzrvBy29/0vJqzDeFztJtSUlyFttpWE
6NQDiGJhegBt3TYi+CzDGQRyqcGCRTmNp+Csump//BKxcvDma05BaGbbOXL4qGU4ftliU+b0+o/p
1LQEoO48Jxi0pvLBAJCSs+WbftIgwb4gxkBsdbFGbRXZRGUabWB/CxIk1biCfsn7L6g8xz0rN/NY
hMwp86L+pYNTXmHBWvMq5s7dnj7HdAIjd69k82Cw0KluZ2Q2y61q2+qGRpLaC4zSu2RN1lyMwq1u
XUH6kyzFVMJLsSLncfWEC+av2oGMRCm4NC8o5wmdXKQONUcS7KYIVdqsDzZUVtPbRXIG6IuuuKPu
4+5Ou3PdsaK7ER9kqYO8zwlhz7aZ80OplwtgS9/w8qEHGz8LeefxL2n6nIAVCiDjOZY1HoXdNq5Y
IA1Z3dxyKqgDK8UBN4QCYTLCXcuaPjUkNDT1MVraOGVcwSXIe0S6SUr5ijIAVsZNk+47DOdnHyKR
/P6yna3BAn9g+YOzTRxM/p5tsk88R6Sx3CciS6EF73mAxhquL4CFiRqW1FyseuTQflSH63c/81hn
4qtOjCbTeFS4XJPQBI8Ml7aZq1zD0KeqvQGnBGJSUASZRq+en0dGEQATWf4yS4Wye3vsYq8uO8Rn
LINPsn2c2lW8AFt2bxBQOiEwIYdt49kcaW7EsFSKN4Y+ddW6wo/h9IatLSnErUBynXU+kO1tsg0J
xlWGXpw3M9+RKtN/hcd9t0bSb5jIQX3D4kXIxebXBZuv+Q2D9WZLnamZ6cF1oNgQ0DmZcxp+858A
niaBPgl9nC5l75y+PgvVlpbNkW/8FA+PTOxQpB5OgFXMXZbus9lYX8OPgBdJ3vNn9QBn2JCmIlr9
xx6vs9FiP273B8ULG76m9ZkHsVuGnASZYNtYmIxI3e+vA5wsinae7UGKia6xPS4DsGBkM/fYsn01
P7lzZDK1ROq+yhkEA/w821uVMEypO/UkV2ijYPPVJK1gfJy+C8bq8c04LHNozJzzkrpcTpchrsas
oIlNSYXcZPWUNSrjvc5TaDtrJh3ltXroV8xkwl6luHL86PiwoXJl3QuVRsrlpJ+SNSUEBlJ0DCby
5vp1f3+BS+57D3XhlvWU2un0ZwyKb5JfrHp4enr4HaRjqXA7OxlPPckdIFFkCOkxyK71QXEGYMZq
yVc9tX4c84jrJqgl85XZumEJPh/pAkOrgDEo/rIgyaiWQXFzVBPtqse/q2W70psFsBIuP81JOrdR
igi7/PIAi+nZARErICXPR4IqAJDpExCVOlAcyra5QB6l2wzjKiLbFHCTvAcWGAo2zOtHvpniwWBy
MpGD32aknxaFgLbVjHIu/1rIGPwdR/A1Z0XLiqDlyzCfIIRve9laNPeZxtg7/VyM+mtPNEd3uZrK
ZW8/vFs6N0O4jvE/Wc++umuvsTcsxunVkcdIsCSoLn0pi2jnjw5yOCh237MZFDZBD7OAHaV8qpxR
f4MxVWcwuTXgIirY0wst9INi2jv74Km2Odj4htVtR20Xu4UDy8MdHKRURWfOJ+N681YBZl6g64R4
ynUupD3Qxt0VemKefSCHK/BYvPpc8NnymH0zRM4wHoczCnBL0nYuM2Czo8d8hK6SbnL0ijInHGr0
5pQHb9mNvqEQUTmxvmaq+ItbsFjKnfekUCXC3x520dh2QszDO4VtWjc67+VBE3LjsfEuNiHfEOBC
fG+K4ymR2xA9Jep64NxyppWGjB+JQYP2E1t1znuUMZ8x1gxYdG3FA5W86MYwA0u/sWC470XgdW5R
I/bVMbemln02NJdseNg+1uI3YPneZNZuCzWveeEd+IL5V5AQajURbIVB0G/Ep8MBjpm1s+yCWa++
HGDVeQEHtgnYpoyhXAHWgjnJ4i/vdYP2jZAblYJPWm6yOh2Y7r5G1xjaHCWwJQtHgKEW8cZyZNGD
QQkX0TrUzR5yJEBV2C/CGH5zewm+R0jUS6Ae0QUs1FH1ozH9uMXEma1Enc4/uS4sI+ccNTSevFyR
EtNBDs3CZ7bI1kRBQt/s/wHAqE2xv6OwVzOXLR1sorOWD+DK2UBwfkMtDXd9bVWaVDaYbwuFDf7F
B6fJlZE7i5JKIhN+X2yB4rV6zwB6jUboQzrB41bQkBdCslTmfe0FlotaWbEqxfzLgjEctK/OATJf
w+QJDQMu6hEZjlE+23IN4icvrg285eo0T9S91fVB9S+Em+ARAfMlBo39Cq74YtxPlUwX4jEEIQMp
KvHqDVX4Ou/e13Rl4ihvz71rmR53Ggq7mphGqO68acmJ03iO04y4GLXcH2uhGAG9QZEWXH7aSOKs
2I7aJiYFgelnTSYWJB5k2eq2qkdHjX3MP13M7M0MPK3Meo+7qu+jguV+Yp8kSkAZkbfywnZsPU4s
hd5BgXwNndIcfdLRni/R9/4x5AOIIoMOhYz31YfpvVGy0mRSjgvwVyj2pM/VSt8Y+S1kB3DXajV7
khaslsQ311eFMSAWPKk+r9bWX+S9suZ911xsCvAEHJLv6Z+sH1dULDM89ni9x3yTqXvuU7K1sU04
z0gmp8LRhmdScFc7HTjJK/HTvTTHgW+lHTdGOQJdo0JahosMzRFXUA5EdNbxDmoWfH/pgDwxvcd4
tzHHkpfF4os38eZuE/mM5lMP9BmQPv7+f1pa71pfM8F4MibC9GM9bM7IW8C4B1etExB8KimtYr30
D1JAFrMMlWjFVoSSTlA4LRj5pdpYd0NFExJ15Ow+QxYVphRPL0SE5H/V+zJYTqAZ5NjUedmX0afm
HeAVtZXu8dK3GoxazQrh6AJeEQo+J0eRfEuoVXfiKQFuYOVuzwv0+Qr+guqEZYJgo/A/+4UgGaHz
93gE3TvpD58iyatuq9y/qDV1xBfZ2FNlqv54SEfqTUMWKYRxmsIfPRfsvR7PhWfFqoxLGt9cmPUR
XslW20vk8acNUeXkvJ7sjyPAR0aerrm9maa8A5UHzhs/7Igr9w0Dds6E1k6e/kGZsjdNWKK2krij
affaRO66P/n+nyoN7K3mWhgdeXolYgmOyOOSmd/Bm10LotfKCQ/sIupT3hsEr1uDpQK99CD9n98Q
Q4pt4eLn5sOHnQGbLUr1LS5cjAuaNDtK6tpmcfVbiGOtgHoP7+KlexSiO27X5omIChTYUD8Gu++l
0XBSNp376oHMXTnTLyQoWMZM0h3mzjFd9qWGqJfeIxQhHG636rDaJD2wcWm0tQ+lC/IY27zp/Ntu
3TFsM4s+66AbN+O0MTE2s7w2tklQWakTfDv2KAEYPFN0qlNc+y6iQU7Zpg5U7+X1qd0fMwighK2y
VRmQE8Yua3mdrv+1wyq0VpuPFK5esijC1KhPl538gQAT9OYwNOVuy15kRAqutUawMmr9m9WNr8GX
LLk8itYFL2Ak8d/JaMA+0OnxmTE12txurc3I4zwbO3mbV+H3ZCpdS+9LCTLu+AWFmedWyTHcQSus
bMKTFxExFc7IHpEodSfk7JkgXUDgr8xEIt5pe4Qz3PCPPIGFV2cFKBZtuKR6ujeexYKtjA5jEEJp
MRj54Z7b+doChsFegT4fGTTuUNhCd0xMwQHq3jm6QQoIUiELyXHMvPOv06+/JmEeqcpbOAXGQMLv
ckFXsKduJAEyP9f/TVTEJELvf9z3IcEwub4qZ/chiykMYUeAETbBawKnhWb3I0pCeTvsgzxEwZMt
bPD6J/2mTj1Bo1YWsRTrK6MnVXmcVw0u4OQzSkBahJc5YFbGHRdoJAMBzjp+XkYfipiGB/9oaZd/
+Ly5aBh58UNSesEnBnMAThIiFx9ZRQYi9z35zVdaTP4N0Jqhb+lKfjycx7VRkGC/9hDLD+4UF2ul
NVmRL89kX+SB5q/p+GQlDREUbzOCw5820RDyP8VFqlzoYX7T9vCfnvIPI8rt28T2wh/tHOLpwjAk
IPeWfR1+2ES6KfuU4vDtOYiRQRy0hZjS26HpKEjiOZQ8k2uh893yEjbRFG/tt2nbd5aZjijLnoCf
12BV0KQInzpwNCEO0VVSLmdSkvBYFUnPzY1+RJ9sCEJn14PRNy0Xr1MKyJFCwbcUJ/HPz+FhqS6S
eCgBgDmJ/p9xU7qHZZ2ORZX+xgL1drg51vewt7eZWzmvAmPrSpa6Pgv48msKKmttSM1w4+Ur7ZSf
uhATLkg9LILT3kNUA0B+/m0UNYeRlJJilU1vblfps/KQf1A+watCsz/Ut46/8bSXkYDCXMi2km9d
eK+94HgiWt0/qXXfIqwgSdfg5xUjBB4XqvCVvDYcGTQJHK4vgg2D0Pg4cIb/dCqbGVIbpa/0E3w0
bCvqSCad06RokOU684zhBg9kABL2ThZ+BnWCtYsZgRKzwmhhAtWvy8186sd7AexdCuRoTlGAmODv
t2aNJMWgjipjHkCVrbaxYSqdeEpjEjJuTXMIZW4rnBcZByEDss8+TFT/Wr8ZPtuWROuzRXeDtVyZ
Sx30nAv5vl13l7BH1tNhd/E02JPs9Mi+wCQVqvBNgGOjcu8dXpVmL65PFng0qn6aNm3BSjHstULY
f7eUHO3j/fW9Shs1QiaxGm5tlibCLrKtwMxglXuQuEdEkFfnKs0OEFpKA5FHVUUx41ooOD/CMAw9
7Av3nNUPpIXvxPoCQUzjE7dCx4CSubpsbjm3Z8PZPIGujr6go+XzqQMbcNxkYj7g9Etnd31Fv80J
vafs+qriCeR1ucnfmKyPcJoY+4PR7CjYSholgNHbushA4mneJTC07ntd8bsoE7Ld/4DFgDlxPjNf
mTSR/qNAKyVhUHakWFbnhUTNdhdR6WZwArOZvu0uS/lfsuX/nNgypFnmV1vAIvdCOK4tIf6aL9E/
NebX5eGyLc74VuBFGNPqaXhminoaoq/UXSJwDZDhiIrkexxpVerXmautMFkzIEHneIN/SMcMGJ7I
wFqDYD84WTqIiX4YYSEGu5IHk/jde7fXZ5bJp158eRrOU33ghElX6xm6+Z9DoCAioiquFpQbuf2S
MvSKc7RdaTp56ErWfIjQaLXuytFgQsRKZVIu62JVsllLc6fA2SDciw1dNlkcntt7EJOb2aB+ru7n
cdju5Lo1YVVRhh2r8iFUglXdD6906j9bLfQGgZo2XCGkrhwDpLAHWTOnlQ4GLFGAVq3uxHLwva57
yD00rP4eifPdkxnZk4CZ3/M4YtW2eEH/e7rec3N+NfsUWnVokAquEwRP1a2AQ5PsIbdUgzskJeVz
B4cBvVt7apcg9hWP+B/Npku8V7ExT66BKDAs8MAXXqP8iT5Iqctzf3CKU4zXCoQv2Z4z50hQs9NT
6p8A6cnkAjR4BTYYE2fc6xHdzRl8HYrJz/20FJc+9vwROnhsL8XkV50ziUiamjv5NfOEvBjSE8uT
CRrbM7KScBH8piFg8dbuzhzzPoA3/Ki0FwTYlc/c0wOykUWHe9B+LBBE22SJQiQWC9879nuIGGyW
XOpM6UX7T1g0ENMXNiZQ2TZqHLvEvd4VWlVcCmtE99wazS+FIvjAM7SMZ+g5SkMI5N/pnA7Uata/
GPuJy56g2zNUcBEqgSjTdFWoVFTcfnMOqtQafl4yq8J3QVQgC2ox/41J57VOKlFoWCBJp7C1rugd
a58hXeW/pdmsgkE1XDU5a90uH5MF35TPp7grATWJFLx0HDt0/PwSd0jvwDki24dB7D6c/YUklMAG
XERhzoC9k8c+t60VIbophI/7pSkiwRC6WTdZqwQCtZAPCBTIXYSxejNt1PDiwDuy+BCBuEHCfy32
eHKn0FIcn2vI/eOMHPKMS9hGQpUce/KFtmIPq/XB0hv7wmTUIPi3B/S76i0NiBYGqfdz9j09t/SK
0uBA/1s4llbbP2szRCqTophZ8d+YUF2A6G47Mgh3LDVrINJgmqCUZOri86aJWNMN1eG8OgJupAQ1
nZakS6c53E1QYH/kZPPNwEcKV9x7nv7M3Hj9NmpFeY6E84ooMs/4fW9dDvRFdD467oGp3h226O5R
2iNaBA1r5kDW0FM7Qv9zgDjq1JFp+cE9zl3K9jwaWnpD/MdA6mvyqmz1ZoFWHxPKX5Nq5GfDGAGC
Gm3ylWlSWmgWC67On2SHcrfhRwA1TTx+73uKoggy1598fMwnYDKUYC9ck5bifdTjaytyEzYJKP0L
kdPjyg9h/L50y/eQlrLVtyCV6BFyqpEQ1KDywRoDTk7wBzYHnb3LJuzWrT+NnCZdNve6GQYSBxJP
tcqL9ufuCKROWWywTJ8OcXHd5QGDvFYNDWp2l2N1IFDGOVYWMclHr8PhbnEhm6m/0xaoBNEBuZYl
ZoIM8Jpq0Hyvv4QrdaEfJjFrK4/y+axOg7gf+7LjXp85vvoxIPdOxqPH4NU1L+9hoezA6074zIzV
HKy/uogNWjSYviRrz+C9BmMjIRbTZnRAwm2dMRsZhjQZ9gN4CiD5j5+7k5zKIs5jE1oKiwZy9k91
rIyJxt5JtRC32qe+LX0adoCwHtSKEPwRxnH0wosBrc6vznjXONCChBoymvxBOJnNRQsdSzeg7XID
wX6uXh1ZcuYbi33ihViBOQoBVmzZH3fMOsunwi8j6F7JfecR5/SYdwzVLdl7LbBMMEu00TNEbX/9
FfKeRyPoSBNHhJZ8AsCc+bN9AZEc0iKIDEV3V2AlG5KTfrVS81pYsshcRajBa48LEHoswsUCQ+9y
rkU0MpXTbEl3zq/FPZGJPoxsNUWYGhnEkno41tUHRhQ0EG5qvpvFSi6tpBmswnVjnmn/1uG12Twx
ygtPTsD9Zh98dnQaJh8Zz3lUqyLe/Nfqofn2h07gtLTLM2czGWBoYwO5aq+QuQ6OXFZLjmYcr+kL
/YiOzXTMRTRZzm3+V5L6qHOqOH4ROVUVHqPnULkKBV/rGVKbaAaspB3Vq0qsPrzP0Q3f9yZXrzmk
wfDR35GsVRW75cGKGebX2lFMLk2qh9ZobhIy+jX8xS+3J+XU40UXXHB3R+z6IWc/Yjd3+SWvlg6t
udah2xBYHyCnvl6Z+yy9VkUemXWaMHonwf1drFypPO8oWPHGppj0YTOmTCsaIUvdwEk27iHaFCx7
gjefRDfczhtM+ce/zO+YUm+pJwY9tEBBCBJnNKkZ7wQB2fZ3RYzxJkCTlf2HWg46O1kjYnd5vCxU
d5E8g3DKC4ZSrhmc5FGUx5/ehozbLaAosu/H0UYnZRW4DP0dyOx6uLOHU+8T/VwxeVVtOzMgrztD
anl91C6HuCRGM/Hu73xkmg9scY+H3lCWeD6emVZ3LaN9T3nmzeWOybEOUE9zRGXGwVktGCnWIMI3
1OP40bPOLs89vs5CfArKFTkwJcAlsNq+jG8SFMcxZeS1QGsXyPvxhkMJhJHcu6+IG+uQUSBSOtf5
blHTAl97tNRT+o5lCjWwjCn5iwRbzG0qoEevfmagmg0wbwxh+2qsuwwcqVwHPp+8tFGcgK7QWMWT
x+E2jpR/Opd12afQjDv9gF+7fvKWIDxZmbNtQ7++UYnmEZ/zC34mjrqeALeRpjInIOJohfaCiwDc
zvo8v7ZgX3sUOG/6kqQLxocTbtmwXZi2Q1Dwvj1h3I961S0+cqIyh91amPkidMgTR4Z6XUkgGB/L
KRuVD6RVohblydlhxlY+hDiMaNn/VnJr0AkmtJGtNULZ+S36z1diUxiZ1JrEbP4bgEQaHQotj0kW
aO5hk5xp/zWw/PTNwA2l8/hJRe4GmT1X/bP71P4PSV6G5o3xtzAxioGnY/SS8W/gZBt22KP3oEFW
Bq1AM1u6yJyiFn56bHOXjw/eHdL8D/Ni5iqOh/U0Xb4hRCrCS/HSqYQUfCVxCHhLoZ58/Mshg8aR
kasqQMM1lLpsb7wX1hf6j+X5MI2wFyB9cJoIgL0vyuoFxRvbIL8y1DYZa8NxoF/mroE796iupsSh
Zgfz4OK7wMTEQIM/b9rYkMeO35Oyl40sszRN4X9WDRynDqJOxoSiyDyjw4iHG4ACen9G85NYjA7q
pegFHAtKEQB5MtpJN58x/QLT6KX9bVUsS13Thj/AYQWIvfTIWo3F+ExEaMKNMs9NBxl3I8ZPWwHB
rIUP0LbHHAhqyQQvTnzQVN52l6WVZQ4RMdws2IwoGk6yFg8Q4/dblVgsrP1T7Ab4+Lqh/VreQMlj
e9QEZGnKb+qDZJFpAvqZDkl38AO1VBufR+DmhuhsSQSxGAnwutLgnFTem7nhFZq4QQ0moQEK/OjI
31t5SsYuLymrr6PUvehqaGJs8Dt2SNl+54Z/5Zqw5K/4DLYwKMPtu7cmFn1arZHxeNWbxeaQCqXE
ay20hH2xShgGC1J98/UVISgGiaIDR2gf/Fx1iENAo8jNf0zyawCfsWXRryFh+lGFy9Y7j94UUAGC
wzTWdk2kWTmSOPnp475c2t3G8z1iAdbZ36OTw+pd6YVm+oMkNBmHdJu+bEkleKBlfawAt4sY53Xx
oZXPx1NkZbcMB418B6W/xM/DLAX1mUfzPBopSbgK4EFgPWpYeoOZakh329W4snmYwZaUoxb9v0fD
SsVcrltz6lRtSpmu8Lmxto2T57o7H9DfkfDRf85StzxZKjAXWK/M3wQG1PnBYqNEDNMC/0/1YgG6
dbqqK05NapId2qFlumm1+hA5RwDA1G0KBLkHnLuetFgr3RGcJNxxxptad8prxmwq+4Y449pXREqd
25FW0u/JPcZ5NKGzMnl3nZSvXcUfEJkjIr4ccSNunPOeEmQYUIyI3jWG2ewORroHg6/V/nErdIWR
jz0gj2Xtuw4zVur0J0ifv53Z1MRD8kwH+QFlfECQWqI4kF+fupp9PCqen2NDCnTfwPI1rEZI9qWR
4l0t/KKT3nbI7Uaw6dgTC2zeIknmVelmC7VL4bveoEibMwv71GmBCvbrd3bHXqHV8R4m4+GoVS2G
QWOLIeI28zNq60xX5j9iCi4PVSmFx9ql8Tlv9JXLUrwJ5E41APmtcYeh6OESLkYH8I8KQKsClqxW
LaWW4jCepjggMsKh6kuDDSRGEfqcUUhEZBHqBXtro5z++gZqATa7XJBYb7f1LQipFLFm8r2aBhTl
UCIfTCcA2kdrVYtn4Dn8ZVjFfIXbtLxTB9CB6VWd38fD6nVe41/UQpPpJYcK1q0Lhzj/zSs8YpHD
R9iFalrZKm8jLW50akUD/Bg/3I/An0EgyLR5XkS9KTp//YLVikfIzkooLBhRgFhJbGYfDZKQzACb
/cTFT99Qyzs7K/XHlN53nEqOipoE1wcyg71iF5emndq3BjA11LyDEELhl05SpiX7Xy//j9rd+Yer
HanBL4GZsj9f49Otdf2neY1AVOavfSiRroBxpwZJcRNDgBa/2dzr1i9Q8HrJxfsBeFwiFZsWw0Me
p3D6d5kssepKfMYMdlW8ftE+kXQs/CfiUMgU4/XCqxEtUdL8LvGVl3see5O+nhM7rL+3ikdUSVso
6aF8PyT8s62hvXe8ys2Mfrrhnlf6ekc/ueIXCPATjWhYf5z6PznXL7ZYZ4jVdwS1I4xRibJUCprB
ryV5QMwVLvDTb6X6ferm0rI2JptmF/lM92mFjtMbykUtaeA+08MhmglutfQKh/W2hCHZ63Sc0cz5
zF6l/ODn96yPdC0vvYvU/0ZzZfn+vNb//7VSa3Ib6kifcExQpO4Btzi+CrK/PgehiHGbTAXv2kgO
jVBmiW+MuAuO2QDXYplI+cqDsQVrDn+xlZApZfVUKf0wYbNxL1qyqKjan5sUcqyRLhNJiBpuDgDP
yAsZsz9jBqnM70xRQ8pnGLGoXzxSFhNHBNrX+AvjosONKfu4avANzppsQsKBFFvnk+Q9WLrzuupw
/z6ASCrHj9DXSf45QOGuDkIfsd01mklPbzP1RFGt4LrAAimxuLUEZwYa0bK5ovpnFQq/BycGRpjb
b4Tsa8CUPpP40u5Z2+rF7oSxtjP/szfM013/hNcweI9dfR1uBd0vJUvNPswwghDBSrPmwrqLUqXw
RKpezmLgxtKsPKfnfv5540FiDxVo0sXNwCi4UJ+bz/JoSEX+S+v8DEZTbT6/32rqwreG/5fq1acG
7kCCBcKs0qks0VBs/5Hwaa5XtCiXOT0ck3DO32p2YQL4WGp9GOaoZzxoitZc7IHgarbg3scs8S3M
aa8+3P4dgc6HYcHtYfwhVf0a4eqgT+CPFhXF5WCoQ2IHN19owj65FNkeiMCyMfJQ3W6n4448xoFI
HJ/5AklDENiZaA3/rOo0rDr7d/jkoVFv2I5Da8oTmvoOwj/CfzdM7xbYV2t/xwYG5t+vxKOKBQ4G
WHHjSpRwBCd04AkaRH/Gd7+qLCD7xULiPtf7WxrXbQxoNFnXB+LNigb1Z2mgfG+27eu2zHa6Muh7
tzZ6CI1BnQ5FRmo5sxtDK0yWgcIjN4wzHINn+67FeR1AaOjtebN5/seFpJUvIavuQOIUFWXVwecb
rwD7WLq9CidfbtnJKKHwFoFq4bPG5IQvrHCm4EOV61iGEG0VM97MNgV3UbCQolXNq6bIJ4su4L+p
Hqy4TkVWcfn8z0/Z548ZMJdUC65Rd0w8FOWLGRcVJIhuZsXaB5bVa+K28JjYF6aKMSn8qB+OwTAW
GfIzILS3uI2niUAMLpR81fhZJ6yx68UgbHl0gk5PEqPVT1gRpytyZDh0Y/UNkVmiSB+14EFTRwTi
Cr/h8KtZHwUmC6xUvss8vu6AyIbY7vCmGO+qOQqXu6rcJOCKP4fB0S/58xUBhqimfIAv2ED+BX2c
55puir4757V/WYi2QbGkTvsxmiJo81z33dGo19fZU6W+B78ijsUZQVap41EhX76BmSBDJ4ZAk3vN
5tDPwyxeTdf0cbHGfxXNZUnGxWCmQyl14m2jtYvHtEe0gOP64g/6apZyzZ9bZFZRGo8D43WfYiTg
mjDyQSJ+5nbhy1SUVHRKIVYiPBSzgL/HwW3QkAIQ8dfNqsHu4epJe0hc6Ap5s4D7G8kH7P9Jnjir
eERjZDlLn+svxzk3FYt+OvZg0e3GkK230E5JLss52NiSaE79Udg3bT+FgQDXG9vs8NcN/vNj3v0M
3wkC9AC5B1GytYPId6v0IW9stHzZiCqJRyEtk6jIpjociXp1c9tZAkciuruaEUM9hS+5xaV+UJ3F
M2RQeMBb+vIaZY/WbasW4IdqAYutNI5MOuiabAboYai4P4zs63Vr0vl5Oa03Z1sHgqZxWYDh8pwE
iKreYra8iv128K4CvhHgH1aL1edRwFhSmlPdSBaZv9jvynxGOhTo8RMcUJ18LbFLluERC7a5ZVMd
3uff9/KUVs9ftY/RIE65iq0bS6Mng9njaYVhubiC9eayW5Kc2TAGW3dw4WyeXU6TFptsHy0LxBSQ
1c0WtoviXANVX0satyrbXOvBQCY0608Scjsh7suzzgjxX/V70lhEG8MCIPG/lDIUcSi5mFY8SuWd
zj1ud9UJ5gnC2yQfEHFc/H/CKjTtor0rbELlU4BUjiLx2yNsjXxvfWyIOmO0z/Nf9ISxlM4tDOnG
1LZ+gwBmGC1j9voLUzrwlXHHQf/soeGSx47TjPDW0BsQQ5k6xN7eFUvbxzGV8kZxovrdTEKEvrtq
Slc7VDrEUzZcWz+eGQSG1evJZntZVecZmJqPGOTk3LqBefo4QgSRjmJT4w7QEa1TYXh2+KhXZOoJ
CT1fBCptui2rMd8V1SU5sN2dlQ1SmmHRB1HMurUbHulS1/TBhJGUygp6AjDptGpWyKQZlWCmf+ip
sE8j89iQDuyf08wC68Gb5dQoqs0xx4TGX28z9Ytea5JeTo/qBYMxA1KwyY2oVqzjDL/XzDXUCmPf
wjbaZJJaSO7LPQVZ3SsKzU87UZDXoPc73alFk9hAF9ClNAoHMCKIuls3gQNoPhDlbWv/G/uP3FJc
0JK/319A+DBXdfP+tyNBJr7gTvDYuTfFVv3rGxscAWp/mGdA1D3Y9sANlS34Q02PXoy9EBy9x5FU
S+OIBYSU4BhiXlCouWn8YCwyJjm6UfT11R6qLSOCfmzMBaNNQ8fxORBmd5GzE5ALkLkQF4Fac14k
tTsISRofCux5DwhfASjvafkz8f7MLKBCOspqJ4y6WkSLLcjvFdBeNg/mbaA9KegNeJJy8+/60OZu
eU7m7OUCatl6iu5oQXjlcawL1+0XSst5KciJVHP+VxH6SfcOa1PC6W8blIwF5wU9VW9lJOjTXkCS
0mJXeThqR3VFAmIwcUIwI9E0rsH9OX7Q00DVaMMXi0+Oa5ocrFCTG+6NsDJn/XaSO+inDNLrxh+B
KUUxinnmMy2A6JdM3UIrgYy+2sMqxnSDbQ4ZLfpALgxhoMSgutcTmb1/6UdT6D8znUKWp+/InS5P
43zmIFh0zawwnQdOYYnXMXZVxSW1Dj0RQ6o29RCakvZHMskK6l0StUEzbhZqtn4AU+aNkotvGcim
m70QcOwEfSsxATihNlVlS0QMh8iJDerjEE3H/qYevJHNxCbph0jSJl0XHIzzF+hfRxHHcEABfEQQ
S7q8vQqzEsdQC+C3PtpLrdIHENfwPWEgcEr0/nYmEcdva+lvoh/Sy0HMHlpUGeTuA26NaMwXqNZ0
XTbjE+WLQYdI5p67rHC5fT9copSQjq/C2Qh0Z0U8f3MnCSkK2n97K8mEo2rMZEE7NkPHTpLV5Im7
FcoNgCOuSz/au1NZJ48E/Xe9JNwyJjiKzstqEpTk0dMTK9lvFQyZ3SL5FLFFMuCDpCvBr2hOxvAm
tlFMN+5NRXIghjxpkrA6Girx4FSb17nDEd+dOlQ+nTWNJo98BKZzf6LOjRnWnD330gK2g6q55Imv
KBsSoT6yR6E8UGDnqfNcgzUjTNBstKP+LdNN8kk299O/9PrFHUq6m91y5YMnSOBuVhXBu14Woa31
Fy+yrqtGxsmonkgsYv2J0/giyuNI5JGBrHE2BCJjTUutzRXO/6CXEazTJRmXXgiF/QhJWwbbJj48
8e5EdEa0Pow9jK82yVk7l/Hb9on+YuHaikZWPecpEMP3+7hNuvxez5SojB9lyEW9c23IlOMIQBOT
uu5kCRv9Rs7SINZejzMQ3kl89U+aZjogCP0KQ2bLFNMCYtSn4V5emMECQWfI3CvN3aKYqQcuyyKi
SRFPSMz4g8oOV3w8lOhvREKFLar9V88y2Sjo9PNwSEYEHN8H4Ta2lidqX38kIiu5IQD1FcvRXk/7
JPKRA5hRdNFRlOOu1jYM4nmikvnhr5qv4PSZfFHvYjh32prb9X0nBbeIml7QwGCxsueo6Y10XLep
mMzXfTJ+a+vvyM9299m5MW8RuZpIQKaqlnxfN0cAdL/LLwHNKRMYU0nuiZGt7fxLxbQEmJgNXq0p
X/8L5JGH20FtyeIFdUbgN+ydwjOPIDdDir6JlnvfW+JZPqZAKGUtFa4ONO0pXiKBKEwXtK4vmMO2
EOx5iUwoXem2e/0wKUBpcL7CFxdJVrDTAiVN7PKRJT1W4SZjTd3SxcFz09Hvk9CXJup4FWMUMNU0
s+5dkFCL9zdsuYplRbS3iUN8PGZwoCnIKWjw2rTBRWJrdxIGm7MQojkubTfRkhwGprDLYDP52ozM
uzMM/5Yu1ataFjlzEYBydOla8vFhBFMwMFeLUgRlbRcjFjAqq/hUWMZ7x7/h95FLD6yd8xYH9QBH
hDv2jdQyJqxypiDubqpEyjwXzwXr/MNlFm9klgNijcTd+hi7pNThU27Hej+JVaXQgPyq6U4bf67s
q5rqj9YzcNEu1pLkX9CZ6/UgM9SL01JC1/JZDONJcqYipIgTTu0Dzfy/xpHsIMzNMNrk96C3rqoR
IYJNiQbUIwltiKz08x4CKa6DTfFzLlPFIQM3S5pkDe14o+nwYIG2/qXLOI+8tqoxTNN5+mTn/Cpm
DBy+avbFytVz6ZFDwUBP0vrkvfRxQmL1H0tIvfCgC9mY3DlvUkdUkTlQNwi3LyF/1bi0RLnMqV9N
iP2OggkARxLC/Bn50056UDAIR22iWF2OPSClBlF8Vbzw1dVsX0PyJQsnWaEbLJRyYLYt4z7LDHQI
crXWcbo0kqicemZZNoAupMOD9ykmG1ieu+swjur+gtMEF4KkUuPA6lYA2Jm4yuK71tk3qq9jmeoq
5pygSEa9K1587FcZBIh2Em8aQJO86PAFU2Sw53WY42Vfea6+yPUploR3k+yUr6VD3orf5Mgb06+6
TDTHoggRbKPQnqfM6a0dECyGfN9uAodX5EBo5LPDXB7dkXAPDP+u7AXVd7hKcWH+VvfxonnS6RHI
/YttZEqHNwL2bMmlJgJl4BRk56JWu9ydT/HtAmmzlwKU7Ne9QiOi4kdwJmZcqOY+Bi138CoqpHKU
A+2Pf4DBtk1GT9OGirItg50QHS5KHeFyOKgtX0Z9EzPjF/RrGwlgYZSuvmq+x7QlOg3FQ774eTRY
eGUvqS4ynPUlnEV2j16kxnFU+Vaj2Q+rr9RWNzpigrO9XEs1z7Z0vqUsMmw1XikfCAUwKHvee9vo
ts1szem1VH8M1fjh7375ZV6UvnkwjLCdCuxVwJHu5daWTzTmBnHx1u8U51+reQOF/Thdnxx3ZFF4
aalaOO7Wy2ndIc+9o8bnPwbwxOYyXf6PxzukFGGnfqKxpITBkVugZrI4Deg/+TAK2/WsNQ/dUCdj
Q9OG0a8Q64/R0bU+K7c7lq6H/AHyq9R/yHqKmsTjLe/kPlG2v6Cmx3VQVfFBPOZguLLhh6pgnaiO
aXhRgUWVdyD2lQX/b4tjEg8ss7v56uC7HqVLTw9odcE/2OtQ/tmczdij0+OPivB0HK0DQRzQsxbn
RJJoOj+kejTPE9YFt0H9boBDmY8NnH4Akv4WzT0b5jy9Frn8cDdD/f0/K5dyb066CfwJBaI1IUnl
UkijRhKxy6Sa1mQWxf/e7q6OWFpDIEnNUOFiI+sQ5RGlBwWKHj8dS4daDhM36PA161XZp7iw77Tc
mX/DpFrDryV+aPVyGTYf77VvF/HJEOYQnQ+u4YeUMUJiBqTURc7KKUYGZXcu/4MHMcwz05MfU9pV
FZBLeDIvFDHVpAhwPv4qJau84b8QpDxkFW/QAngiTiZYdTaWucb/M8tY+CLLKmhNhhj8iSXPswEf
jiHypp0EHbyZKgXX9GIzWGbPQwo9PWqGio6yMJ7eVep8p56+71uOEvMWMO5cu1ZiBAoxtF5+pPvS
+uhBj7rReZMm90JTGosg1Um61sYXG88sxNbJUaFgMxst4l0EFr6rlO2PU4cJ2FsFrRZMk9VHTY52
50mvnW1c5CMGXKf1fEBpQwaw59J7umSSxhTMXwLe/o26ZQ29T3Asdd5e7a5/7TPDcRR7vwvTbt4c
eAK+4+ZdA606k7HLqAbeE8zXQMkPd3EQ6/E2Zo2bmH77Xw4PLjS3gGMJqb8+xK09O4kRCdr4zpqa
H3tSuWSqty4GcZuIDK8AKTKPyS5LHXWEkuS0FkUm4vvpwZhNlnA4UXfyEVGpH4uEeEGbnsOGdA6T
dUx/cj27LdA2iH7RfGejAjnjDYmX8Yje63ZhtgfXa9fNS9Dz8xDqqx8Eo9IE4NEeJ7jd6BaERTqE
yJBu5W4UaGlt0/juohvi3vwVGms4tPQIEYgfEmVzSp6sjDmq1EIBSIobFVnGBQdn5n/gDsrPVnCY
VsaZW316ESlhKIdrUufgMDnafyQS6+0DGVLiemhyCxV+EYA9dSVxVkd3NYSxpRkX2qmg3wYSO7ks
T1LHSBUnfrXLmvPQwa9h9vfstPRHu4yEhr4fwUi1DkJlHrnoXV73U3iXL/aX9+5MQf6032obhHb8
7Ae53b+2oP6n4jiQ1npJHvKeSyGSV+Aza5U5P5pcfrWBQO0h+gCmVa87ZVrcQpPFbXPp52W/js9N
zOk5jtCIoBDdM05d7i1xtM+8Rgwg1SSKmgwgINNKAPGX+mHku3U4pGPsbyw42JfauddsNlpEnWA9
Vjj7/lJz2N0kgil7FtYfeR1rjl3WwViG5dI3CV/znysieTJFcKGQ76Mmwn7DJMx644zziR3FPWnG
N/WjkKuoCaupIl8Dvwg5+Olsd4oYmIPFLI/kSEbylWYQygfjVtxpCtA/wbgzLGTD06/fIUg3HkpU
mJjiS3L8tWfeR2lPJs1waEKAIRdWbFvhuKyW6CRaeHsfPVM1sz8jifcCHf2fDl4eCnOsP3CV3VDn
SUEHpZmJT0DDrlRlB/9DlvNUk32tPncZ7PYByBop783ql6REUYpmfl6dchy7e611fyT+1dMgAI3u
fVUS12nhmnTaqyuSBmCCwC8hZe0j0JZJQjfQQ0KLL4OnqUR8WJjweQ5AOPCUeKpse0/tVmskvM8r
XR30n3kwRJyQVMzSXABTchHIhKEmtka2rwFyeEUwFWuybhUHRHuj5aZ61umYSR84h1w3cz+9Kmf2
QYcwlJhAPoBxf/QJUjW1v0HeEJ448LTn/gmvuaLmDQhfMhPa/1BgIorBTeOuPlxPKRnJwbtTLssI
4Faf0toD6G3AWtLaKtnGELtQ8mat5PbQJpN2mRYcm4D/X8SbU5ySyexUcJiqSRR5aBfozSEGz39h
PRlEZigumOk5o4g718VFYVzUichIII1/qBMTOpXQFWBoP4k3GoGXQE+IaXQZJezp1IsO+qQPb3pN
1BulUqw1u+cX2vc27cORekdEwPySR3WJ90djybm4pQuOT8yLe2YoDLBAKj9IKaFmsY7d6x8sGBA9
YV32GWXTj5FJ2K6V/gndDd7lPDDPDMF2j7b7pam2RcPLkre0uCXD+kj2j+cusNLIkreZOgQbooXi
9ZAJ8icPLF51HmjOsWubpsuIQ7Ja4bXfgSQ42ljVHrrfM/UzkwtbJvxciNYG1FLAS/u9RBU0M3/V
+h5C7+zS0ELBjqNjf4ZVdqQPmWYAY9fTbBTHl6Szstva0MIL8pwXWTXCmLZ5nHJdNnQG/RwkxjRW
4xjc2WmHM5e6zMecvrCavKLBgSpFoVt02JHiLbGNyV9US+JGqBfdeBlcdnzBXfq2U6jXmHZeNkZ1
pN3ZsSBYnkT5X7XEJV+3clbsZBi1f884yx5NaJx6sszu9m6cxfHwv2rro9g6UOAp1zPIaQgm8/08
4XHT6E2VAZIH/RIVeFs3nELUV3eU2DqEoKlApvNqgqKpwt3Xjnqf28bSqWJV0ZkFXqfRy/LzIFNw
4PXkbPHhkR8eMgQuD/CP1g6Wq9tlqDFNXSyuoMurSRokmeCJh3sskyO9e+VcF+cokUZNLV/pEWBN
qosFchAr/CZAtdApYWgq8a0S0QArzKWdVAjxaKLZAICQhLKNK2X6O/I/w27XwUS7DXIqHxBduLHW
cKJrYwmD96U7uCUWqwyq6zN5uAi+U/4/GX0wWI+mHxrIsLRBVdbuUblH3/A2EJ2pYKjjNFnZTsxP
o2M1KpXz7RGmoCZf2YZ39baozEpBlC6FRL1/UqLTD6rL7Co2g66yx/iI34IsCg9w+wQI3z5ZSWvG
Em9a+JxiVAvrIBEvoTxdbfclTPLSl+5gkSJUL/4e9XJ4NJzWilCxONXbTuuWWjnweQ+wtNpZswxq
grYB3GkPFOiLdDafE8Tq5c1HkAQX9PtdIiIwDpD6FeY8qE+x9qqS6tPPYU1Ts4hYfmsJzZETiwlX
hykZgSe3i5uGYbkmUh0VuvZXwd8GwuAWbXOfttvR37vT85k5TN5+qy5GdsOm5slpaCTOD4RKyufi
4tTZsAsSbMqWqe3PwGskSBrrsCBdwSk2XNgCNxPQH6DklSEQXWZujdY2/lsVGXmPYa7q7Un4OYwB
UedsbISh4yfjRlo66LUP0yw10PWFKWJtyuMvm/eSFKIeKAHZrIcTXVSEVRNQ0jxPDPRpnONYZS5A
SlRI58jQ5y5/rWQob7g775ASI5ErDvLMGuvccL4PAfF3czA1Mg3c2zC76NxkyhCujIZyR4AB+DpD
/pQqCBeeB8nphjIBgyh7UJWI7byN/vufjpoZ7yCtPOHjev6YdZszdLgV2Ia1bVvODPFOM5uEFglO
6uODColWBARrFh/sOdqOyF1nal2O3TjHA+1ssP+hqVay4lpC/SmasX5F+MqmrDq8im7egppjP4P9
G85/hHZ3i3tMfUQ3nu/QznUIzVXxG0g1SxOW2sSOxoAKSbwSmfuwWiRYtcftW+6Gu5PASFyDXplj
3/Eb4d7QSRNyesQHmowpQK/8zzIvFp1RA8kDrQg39vhXz7232vfyx3APmgZwYu7kpBbC1wlsfQDI
frZ3x5kpu+APXTwgBmSW/QKWLrAHbtBn2UPNgdIvY/e/yRRjXeVx+iBEYtnyqGxXj8r635XzZOjt
KTHQ8drHQdC3kPNzwogq/Kx/vCE53/arczNT5FW7hhcyQz2EBAlRUEZjX4Bf/ylA6nFTqCw5enom
JYFVIWKXSVc/OhIhSw+QQyFWAFgUOZ9iFMytaMLfRV9BXPmPkZElCuXDTsZ/puXmGJRbWcVhAzCm
XOfQ/YIkWZIFMJ9Be/xzOiG+EBzEr7N0poZc9n5XN3lphUnflwyjXYQ39Ncv7llY9+3GdTTfEC1K
zzTiqR6XdFef3AocfQl0a3J2+q/tYUVyvHfeOBqko578DwydPp+zE/hc4aUoSjIT8KCn/r8mZuVL
DG6aRVTDE24dtGxgWgcL3A/xldVf60KxKNVwuJyWD/VAflhxuvU28WCL49VHzx5l0loGlQ+LIeGL
t8bAEZ+AYW2rIuPBlJ6+y1SDKV8T3+AMlLkp2YvwC9HjXA6PuIxlFBvy6sLYvmHFWGOwBqkpm1ip
wurZGuBvJhJi9V8IXjYhivfeO5v8xxsDisrC+e8e1WV1OMWH39O/owG4Ev6j48as968qUSOJnkVb
3+8vw9CKcyAY1t0JbgPe72sonENSDVFaDqLbZBFJp41rnSBIH14wZcmb2PXVZzY22blzXQ6l98kR
o4egdXtHIXYZ6cy8BL8FetZUGVhQZ9UnGTQqFb/m1oVzP0hxCLfmQc6UGK9oW7N3N/58CjrmxmaP
QXE9kD3URSf8vjnIFHFvBhh9sqAMckmpJ6/xfWNXdkBGiDxLxwa4O2OLWbF4v5BDAf9nDAWsRZHQ
qfCPa1UNwrI5a27phMZooZ4pCE0AquTnpYLCfje4jBniy1uDg2ehkezZwtEZQcuRSlmKGIV+JTzA
OfDSoRJN4biS/qFHVDoJO8k9CO4zMOBjT5n9lTNiqKpk/F6o52XKAw/vXkN6QZxJMz5tyBuPV7hH
8d9+6jnp+i6/TPXOTWIq4a9A6UeehoUwBDnMlAm3rmtVlbQrSrdcTxiChkotpd6mCCEIZoAHz9uU
jiHyQ7a+QbI4N61blcOpEAi5aa4dnKX6Iwy/qIHp/MrzPC0YlsFHlbJfGIMcqDWQvxPvMRAoDUQP
/pUbHV27nXfVGkif+OoiyPuERpzjHL5VREvK9kvNaHvEwstD/otjsnoRWCctpIFQDyCOas7hcJMl
Xlf9AJgqa1hM7qnqLmsp64UPTstTh/kxUjQS7lrKlqzk26mfmj1nKj7Ttl2ZFeXybwj5HG+kzl5B
3jIMQ7UFrbT9dXjsFeOdRQPC2nvWFkagDN3Qp2gzEu4d3IyfQX4g7ACGzx3zu1BVaEgeOnO6V5dN
PqejkcNU+PGgLRjw0x5RRdHlfB0+43VZljZAWxwDJcVhmEtbEMxBUD/5KKvsU/Xuvfb2WtHVGNhT
lBkcCudiNjqqzDWkYvIBdkulpGpKnlTf6SCIHKijIMHuOcgtRMuY7TQE2oEXIvhHJJ4LKZKL2Jwx
asltNwoexGAjQkhnUXF1rjXR7m/yjNnNBU2DmB3CSnldv6VZVxzipSrAezrpmxzfqBB0AP7NKbjo
bx04Ngljorr2zpX0VnNL1MfzjS/wypwGl37YXPcyJSFrziYf5PbOcUC4sasswnmKnQC3Up8mrvKH
4RyRQae/i6UEfnv2qTdipBzwZl3DfSPlA3wr1DE9BzJxiQh5k4Ux00AsvO/VOCQk8WqeDme5mpdK
Rh2fNqCmHYBjza24p2LtfAz6sX4r+AbDVuTgJ52HL4EqYPED5+jrGJBlBrkStoKKSxwEUhMBGsIA
14nk8UFrqrRcklMzcxt+riY2pcccRTINRwkLqG3FpcX1bcH5zx/p641a6YlFKcYk/RZaTz+hNp/Q
RwyiD3zDF7jRc/unV6HjuCcW5y8pI7c3vvY6jY//lGwIB5wOYqfwGs6FoNOsaoRKxs+wEO94yWzZ
Are87kGBy98bvp+zS2BRm/FCpYaf+gqJrzPssdXoCCz6w8fxjpS2UwwdJpL1PRpt3cVC3s8dSKZZ
WjEYXLpZydLRJO3FrTcaTGAjYqncw32+8fjJrhXo7TLysWJVTZ7YEl/90fvAcdcknk3P8ivmPY5e
IWzrwjEpK2LqRTSVH52zirPEwdphPZumTt2RiH1SoUGdgQeH2brZtoE7o8GjtlJ/1W5XBSg/NCb9
jXngvxYYqUeFatojrekO9CmF3j4etfzksLgxg9lKOLy1VV3ClgfC+nPDfQorxPc6BFjbjaUoZl38
K9lXZ1Bm8cs0w0whlHnF7F0f4sMfYDUQSzSaZtJ551/n5nEGtYf+Xw8uPtMhQZUuXXqKVosKSAn1
a0WrYiPTRuUAMtavY2Z+D/FAqdl/4lcrRWgHiLzrS9pOUEl/We8dh7RRpc6Xnz93DfvIEhLaB8UB
5iAGcQp9k67ITPzxXNEnammCDrEUXAm7XwoyT4XA5Rb2M9pv6StzmSPO/9IWdGOd4v6Ae8/35Auj
UIimim1lYiRrZKt7NQWtqCauF7pdXQN5BrgmphSPlMj4RQQZn602dKsjYaNhsIQ04e6p9q/zPjjo
iuEAWoTj56Lf4wL292zry6eXFuKtNTZpDriE1HLw+Aicl5j6Jbb8ftBchZYgLA1+Hoya5+u0gaDi
4HQvqPKlfmVl4ymj+DeGecoxe9plgah19S2DNPT/pnQ6hjGVOUqwyc8veoC6stP1LK/Xs2yMPWa/
g9oSYe54PLerGGo+wfwzcBNs+7t5CbDehbqDxzjK81ULSf+L6KL01ZzCzOLth5JRnU93+WdV/bLo
3hU9J5g7GrN1XWFIIOytH1Xt72dcaJIQMsXFrFOIqLKvBD750JtKRs+SVBJ5hRlgc5lyLMIPSdoK
TUMlDQarikPMRVLw2FmHZIPwzt583cjJFyhYBG49yGrmBP4CrBp5SR6rvd9d9F2z2mRk9ar/AqTY
aiH6etD9ATdDTvtCRB+pLae9Kpfvnja6JRpb8+6BO0UGXCdNFgc/4qgKXdnubdLeQTublzeLN6Hj
JyJ8C6jC7VyTc/wwRFa6LnsMyFIDe5SAPjfKAcN5m+QILG49Bij4KFwRCloX/TCacCH5JcneAf4y
0O9p85imfoZnbxQy5mWsdUaRdCTU7O1+6dClPW6Sx1Jy+TI4S0Sznpokd3mwEmBes6E1YFXfehnt
3mDm8GKevXK0B44fpA0ZD8XPpq4/a7Tkttc3CC2Nc5I89yfIDQNkEQvy5mDIDxuk0ol2FdHyUgl2
uEX7wd54mk6iLdBL+VBDFXz78p3kKcu62c7hFPU5x72UXvJIhz+3FNicmZngQbJ4Zbrpr09ICf1i
hLvNID3gA3PuZkodDRt+gArkwvJyTQYRvbAbBlQgRLQKvi8epQJ5neW0ICRy2eK3QWUET7lkulEC
PSEX1AYSHEdKD5NEInPgGnGPt9NUOAvSo2k3RjTHz3F6ZiKqLVs9dtc5TtIsR6bBM3JjV6Cw80mr
yp1bEOQhmu+BSpBttGb60KGR2nIScb09PfZMXyA7SIigr37eufXQFm+gZ/McW/1Jyg9uHFukLbua
zWrUe/qc72KxtPEHvVyPwws1O5YVaKrOkqUS6tlMFQP+451UXHA0LE1sbhFbd7OFxhKG173XfVf7
dOlaJfPhkx+mysD7vfaPFrk6deMGAwI4yv3s91F46fFHNSPEukdB8Yj/0yC7nlO2oeB0ks4m7+2F
GaqfZU19OIab1iDOUZ66a1ln2ATrHN6HrGQPpZ9hZMaCrLNcYMrsZ/Ww0TLsXrDvoxT1H9r1beJK
d+psRO48V5uee2S5xYki3Ff0EZEBWB4lx0wqWkU0XtgB9kM3pVqr2JfQ4i62gzK2aPBRcmItPo7i
gOPefxNeTr+a3yO29mYr13mW6IAPzM8GkgAe0odTBg+vEz52m6N/OXtxD1xCDQJEdEHKpavN/1gg
p47YK2hpdPRsNg2lhpJI9pOaeMoa0/dSi5pm2ljCYerdmqoHq7O9oYTUeiHxTcpuKzgJFAiKOpCx
YVgf9vnG7r093a7hHHr92j2GWQiu51cGkbo252zv0F4SgZJ9B2tdp/5xuvycnGbIK1/+TjQGuOUo
60JaS1phmfPKN1c7rJpUMFIHPYWuZx01denS2Y8jA03qqkAQly2BlGK7/ICGjxQcNf+d096+jpS6
p3A5z+wUGXn/sLYiPXOxAOPuiL8n6QQfGM42HbbBg6GdRBV0K0rClKC/HwNli9i5DWa+4Wcgp4dZ
TW2XbfavPTg4GuSZ+OmD3QqSf0IAEHp2KxPcvraWEPHExRLR24umN2M5QPxXZDH+50UJqcsKDEtn
NSFw7v+Zst5hH8CgKe3RM0A2OBdahv6n+fRTUtI3HdxHxTeBCgnBeEigpDn+Z2oybRS9Hf17CQQV
OkuXaBP1+VjqxH5zvZZatj9fyXN6tkawNXc0CR1YWEQPtd3j114WCtM+8KGgAzP3IkAOviUvNIBz
sNHCQ6V6Wi3KK/kfX3W65t3TLIZx80a5xHcAOkPNnc0CccakYRPT2LRhufQQBVqIgJzLBTzUHXV7
U/eARVSj0pPWPw+fXadFCwuCHbc3ujHnZ2G6slIj/dQQp8vhkyf/nd846UbvpSK20FcTagTxVMBw
co2IZe33ikVyfzmnMXR+oUBhick3IAAsowQ1gXUk6hmUe1+Np5B5+EY+wLB4Nutq29cmRJU//zZ2
tHF+A2jmge9qeN0tBuOKWv38jh5otIUcwAgeysAvwkPCqjoay9+QX/zENsbBLJehM6CZhe6qqno6
ngxiLc9ClW1oiBtiRD/S5C6I6fj++9NrlH7o6tiOLCRxYQM//6XAeo5yfaXsjbZ6BiSgAwfC7r9V
AzcecXXXi7+FkkW3ZhuVKbhz/UBcse2ate1arrg5xKDx1hvF1/6q6ptD93lzl5+pl11X1ER5pWdF
dt/vA2QBjRdvEf7JC9hbcjgcDOui/J7eqqeCY3WrTXIEDug8ehuAiy/LIy2JscyfIi+7LsMuUiRw
2hBDJY/p8zS7LcFeuveY4zctNGerGSZlxbCUIj73FRnfwv3e/n9SShnqhrep7K4lSfqwsVn/kiWG
uzTTDWM+NHo23OAstKePAM8jrB9JF9YvC7k9sL3iIGa+KUTtBuboLpQ8xREenVIkdp5MI23rus4y
u1Yc2QQZ4p09bY5KWUhL34N5bUQcpmKkpokR4k62FCBqo18qU6xr8YmwPjnqzvcWc4B4pAgXWkJ0
dhwj8HB23WCQhTOyKIjC7yV8wkcj6E8UlVXHFpjPPg36awEUWMEudN6S4IUOgH9wGkiz2jy/N4tZ
pt1u8r1hHS1t/+DAK/Bp7D0h4TBYBSx8kn/3TMc+5/pB9ctRtgtb1TC+T4gi3d2/ayd5depT2Evj
tFjbq0N5XU8Zzku5wWhYYmngH0WOjGhWjMig7oLA60+InkSN04Q6kdYgmYV/ZXLOiL2I+J7xx0ne
KyngoTLjGy9Xs8OUtVAHLrIO7s3gt9KhNfcLBNNXZEsfwlp+RRb0IuDZlHzDknhG2m3UJC1w8pfu
aFpAlp7ZX5yb/J9++IbFKvJtDhepZR9JNGYxtUSJEYYE6vycxday2XI1HGg6RU4HuxS9eOOaBhv4
4L22rOVAPa5i5hbuOT4zTLyQj0H/w7In/r67bJx0KdIWIKLoI7X+1GNa/yabtEkxQ9go65i/04Sf
6aG9WZQZDpeGMq2Vtk8It7cIK4drxGq2Tnh6BxhWI/sZXJz2CU9C9/CeAHCn7o0lBKh3AhZTcXDX
IjANzqWH9aE4Lo0iw5hOHQfzKBGmcpAgwAvJb5qDgCHGXv7F5WqTXu9pRVulGh+YzCiTkziYWXNX
TmSO0LHAgg3i8eAve3mO6MFWzG5EMRuKhZbzUQoWbDDKnVxGssPv5+c/4oxWj7DwsjdB0N9Yvmvv
TNvpyecbARsP7bI3hPHSfrVQv+CX1bqBQsekULeDRbvpEsxFKAiRFdP6aW70vbFrspy0xHeUZSZZ
Bdsnb5udhiNq1Ix+1fD4t5/xqfVxN7CdzViTEWt70gHbJKq5iO7HXyq/Nx17yXrz8rWnZHxilGTp
tf1zR+WYQrul/e4nTsy4lYV/dETIXOLa2sHA/CAimgZFRiK8JK4Y19/Tuvv0PAqVAmhWSBw4g9Li
oUl8JJ3lpusg/Y+W5biKV1d5iuc0M1nw53or86cIMpwH1OhrPUo+tmpbsoKEA9iFCA/G/1wR5ToB
RyYnhPZReAalzxNwW8fvr7igeHYQQfSssiMGlwG3nhE0k3oEI8VM0lxrZFCCRgM/aYzxwdjjrusw
aaK3e2XxVbO7vPfyNA4FBt35ot9j6Yh8NkxQnJtsPT13+JBNCJsPiwLgm5WmNOPned9IL1XN7HeV
oKLMUF9oZydPsDk7FMqI7vgePp6sc2JuPZ5W/BK2WaXAcc25q72oeEGVXFR8g1sEj7m2EFyqPv/h
mhuxhnmPuAdvVd0AZYO3ZM7D5geo1x/GVDLBUn6OfClywY0tPFOdI3FBwYaDAd847FEiG0NVBR4v
4OlvOCJ04YVyjYfvBFj0a62piOVjXyfj/HhPtZLRAAZXK0rcjHsCPfXghapIjEKWNXuVEJzchV0e
T84z0ZwdhvR1u6sKkXnKpgUWNYu694axB8wduKv724dUYWxTqgITnAVctPyUzKnj6nH3JIKm2zcn
eVedLCNHdOBnGtQDGf4ejIBDC9R4IuVA+YX3gduLrRcr7fj7n9LAtjoR+Pa62pOQbHSPHsyYVKJ/
j+dsIwJDAaFjwI5xX8nU/3BdknTKybYLYjIUwdq97QLBGdC/xKUIXD2uTNc417MljQTBp3qlgvfo
GYj6IGDoBeXNUEuENQm+jW4520HUHigcJsQMiETI8XcV3xUPjV24Qd0egxenY5QoSIYdUMvPQ+4r
WFVkTQeGJfz/34cqcOeVsB6tEUADsi2mQhQxQCag8URwE+GbqQmIiMb8SwUeFMLf+oD5jbRfIjaQ
DfrvtCcaUkTpfyO83u/I+w8RvkYObgd98vTTYgrn6bX70hlXMozSL78dXV7bPEOXZ+WIM/EAhIKU
kU/d4bUWIXdSmJl9NdB+kGPATmSfCYZUshcX6CGjPtJlZfglFuPpNH2jG8J6SiVZ0Ng3aIGqgC0m
jZG5q+9gdbErHcRVY2TQe+DvDk7VOs2coZ/JhdMNmqFOUG4aC92caJeWJcX24oRxGxZqKR1M/AYl
6fVbGus87h4HzT1RkvvU/nlIKV17cIR3KCEsLbEYZSGX8w4F5xbuevq7Jm75kU5GqB7wCgMZyY7B
guXGGdXsEprA4Ok/hH2HtS9GgQoQGiOcihdH7yU7a6efNx4Omk2AzT2O5tq3dFb3pk41CpXMzFFp
YEA0pbCq7a7pTDAUAnEnrRqwEsAX5l5GwTWy0ruFA9HZQorZ3wCO/53nMQhV/Ac05M+QWwP2+3FB
wF2NpURAaS7FlsgagvIDaO0ed/m25SoHpZAiBvwvEXPCtTjs1iUoAb/a++6KtK1JvyFLDWj31AgB
/x+n8Fp/mNDbSRrzkmVjj9X/LHhIrVfJzw5RriR8AgEcRG26KIxWYt04qKEWSc7JCeGQsu3rMlK4
SeCqD+KM1EZuZstwbGEa91/74kg+WLWZKt/9aO0cpl6e2FaAtRDAxrUgpQkY0S00JIPxYH1XDeuz
CZldCwBMPK9/Mi8GEbfDCL/HBmxY9RzMkMc0bYxKtpISI/Q7vFf4/BLSdb/utgHu4XhlyTfTEii+
ffRTvqQ11E7o16iSW/ApXyrKnhl1uCYjK3pd94CNGsj5DwjVbqqV2bcTZpF9OHViCXzQhjinxvlX
57mpTkx5OsHFNRO/zwVVXWWET3jf+T9rqpmUln2OenV2sjBc/IoQ0g67YgFNI5scrRQm7Ss1VRpe
jVdTKBsK63ep/psSORhETXnemD6y6ogHpEOf9b1PV77Anym1tiRVqtjeUv1rVYrHEBss4IcObgYY
7jDsTsI7dD40awQdul/NGIUdsa9NMQMp5w94QiPcs4HrXGObBSZyIjZb/H5aCO2sblYBQjb4PAvv
pDrhomBPeXJJBCJNvtkIpL9fYaMksByMVyCiQbpzUFVXdIe11BFzuqY/DQLFwy+Sc4mKYwrp9ZMP
uytEaRARf4bga+QsaCcYwlO9vx/QLtF77Dx5odJF5kTyZKJtl+Q5mgffx4nL5BScP5KcrViGNc65
8QIkyTxkQhRGorDnKw5VFPZF9/VRmvS0rmkk0kaKO1bHG9C3whuNe/Rpus6lmxw0Fir3Ng4OshAG
cxx/yuL5dOxTs49Xz1UQtd5bimGk8U2WWdcnpuHCI4Dcl6fd1+Oe4DmrQoJzipvOLTTd/f3CU776
FZ/HIAHPRQiKqJLS4b2qbRArNdAnDL7bRPjLtXXNyx2dy2LeoCoU0Ld9nwTtK4zlDimYqM7LMy/b
HwsOw7DvJaiCB7bh2VTjBkbvtJRGle9SGTEsx50LoSrdALkx710kRCf77L/mgv03pc0ahoPWXZNt
pz7n6B69qlcQ7zZIGH5UANvQQc6SDpdHhCTKM6ZS1vTznDSwiWdtDUTDnnq3Qqqa/lUfPCaV+mp2
hjn7oVQ+qjQGmYjW2DGP9PI+xNlfoj96NHez/pRv4i4zSEaf50nEVOmI4+IFh29dpQ7H7qUtQXQp
Jq9SWOYnEYUt2/i4Cibk4Um8bUw8FXpOYtpV9pazv8eu1nDLbf2pANU9ehIClxW9LaXfzUXEheV5
UuCzBsfsN1iHZHSJlcGfue+iOet3bwaJNYXkYHjlzdGsxGJCbnN/noU/4Fi2P5mGlkO7m37EDtCt
W5lIzZDiRIdwwMJRzzpTwMDBWcNKROWAXf3Y0dhTNXmpsn0hx6CrRc4QBRu2QgithqMNbTfRPdTg
CI+q5W2jdK2Qpzy+W6N5YAVGX4VsV0gTIlhM3dn6HwaY4wHCroPaEj4JaVadRiLo62vlPPGZRjz4
mzPa3aCDj4CTBfww6DnB7XeSfi7Ek+4GRoD0UpoT6o4iQEIvVycDVJEiqYppZBA2YAHVe7ql/qVl
Qf99PekQ3yWKNOX/ttJ4aAxq0+nO13KL/Q5bpuT7JzOd+1pzKibn8vb/iMW2q8FRVThWkuoLDmWf
bf0F2L7W9bZQJpG/4Yh+gT/U6zv8RJA4mqeXr/5O7Cm6HLrmXc/+jAX8mTWVgdfeYAkg1JxNYEsM
bxHwc6T5DNJw3mROaeOZsFmye1A4MPyixgK6ug5rfc4UbVeRnn7Cb9fKb3tksjinLwN8JPwg/Y5P
KTRVCxp8ABZFjyN/BoNdxhI84aZJwqQbL/YXMlap92vnX0HYyWUEFOEZSGppPuWJo6z1OrcxZc5v
W3R/gZ+4ET260pARWkFSTunCvhAIJ0ZYrqX/m0ulzbB+cl6cVFfdCEpTnr8rkBIPnDVSG0wm+x8Q
zrg7XQp0dL4IJw6kZPYiAxrg57Oc7Gy/ewiBmWoVlqlNT9iIPbQm2vCTVdAQldL7LFtzKWjXAel0
U9ok5QYSHEV7jOIwXBP4r0FSeaXI9M8lKNFDQl8Ukg6GpuZ+DRyPRdp8uCw367g5gBxI5oE/HEv9
VT/nVBBgIbXkAjFEUF2xELNt1Yo6Y2XkFElWf6HK3sYy5Oqu7feWNRHsMDo+mA8ksMg/7RmZ1G5c
GMEpVa0Awf0P5Em52as5ma+zcQ7vxdNDbva7FBIwRLRRUabQas91ZKFQZb06cGmdx5P76qW7jdxP
TU8RQ9/kFFK9mOX2jpvZ7CSVYPxJSmrOkQDNt8pj3Esm+MVNnlKihvHIMY6bhWYyFXqbFF9i2UHg
vVuN4C92o8Y7iATNljkieJ+bjbNVs8fWR07ODrXdf2SO2brsTb7F3WG+QIulCEZF1+z7Sf/DhiEQ
Ghlp0mle+/aoeC1KwaGetSDUaoUxtKvPuDhY4zc4jYUPualEXb7uiU9/LbZuKITpc3W7+81gOVpc
Un7a3tnaIQZIZTm2RSbb31ouc3Zhr0Fo+EUm+04jA8KY/1QUp9nIipR/x2Z57wM3AoxywHdzPK2F
PMjp/mQlOTZd1NDXf8grGkrKMZAgCJQ3ibNJ+Bbcxam/aJBkKjEeexhsNkZfEpG4H7JYIyBFMliV
dgC2IDm54XTSVRG1WOWxYrfvalOk/PGh/eTc0ZiqoQEnNmWZHsPQ7rJavPLnLkVyuIuvoodVT7rZ
aQZ3CZx9RMKE7aUTNQHyfuZ7Lvxw/5S1MXTd5zgpeykx+c6ysl6DKfxbiPUoy5cfqu/4y0kerE0I
l2hvJqaSqS4QBpzl4Sjpjx2cNCT10u99tmZeHQafYbznynVmzb6Yll5x/YHC6lm9oUHVEDDMwIP3
CsItFu4L8jl2QwvXrBJZ9dwBz5fCO6kXtCW3dq2PGJhomjMMkCLaCSqGW/kg7c3VMQkDpjWzd5Fw
3uaQE7Z1wGJwCm+1+XkzVShGUtVy9tZue32w5PQFtRShIF4Wg80Rc4Ukt9YaR3P2nW5YuT+fBWtt
n04gHkSARN3XwH1YTUwVROmJ5lh3mcQz9wEX5QJh/PGvPPe76aMLizvHXoReKxhF39bb4I8l5NPZ
iFQlhUsCrjGu6E3mD7Z3lOyUETrgj0Ivh+47oHY3KqL4sEuhKuPyq/JdZ1fdE2xqOz2/s3k5H8ys
LkxgqL6QiVyNYGS7cBWsb7g/R64JAGwBZM2yxF6qhjk8qJGDgj0uDN93ygg8s6jKdX2CdTDWYWP8
8DixWQkRVdXkLU1U0TaJEt5Z85bkIwqF7emgsOVKeoa/edMUFiL+H3901MEuhFmCVy6GZ4coHu4i
zyXVhy1jEMv1jesjt6sAlEtgC8Wv37Z8RosMgh58Vf+s/IpHvNoili3diEYe+maCyEb1hNO6zRj+
BVvnKvJPYEHxq09BUHGEfmosfJIhdGa0Wym8Hq03Nj+sPrFHVCLNwWNwOttUAZ03w3GoxUt2zCRZ
Vm3DLVGxcGczBhrJudIYz0e25pcBDiOVfAv6InHqVW8F+Dp9LLHMevYikhYWnSBDSvEOMcR1vc0h
yD1YrWVTtc3VWKgXBt/0VPLnN/K1RR5w49UZPEkaR7pa1sGz0yytF3U+W7oBTiZz7kfFKDzqxehD
rTgc62W7QjfrOpuEmgbHzuU51AlThxuNKdWpxf75RAxFXKhF+i8GYIDz8rksmAXnS4lMJJyfMJnD
jBSgISN+U/kj2/3I+r4FJs2ajeRC8q4fa40VUfM0p+Tobcb4f+0mlNNGpIdI55PM+XQIc176pMxa
p4++nDsXgWaJnCkQ69PqZtk0l7O1A1uKK9Ps/TX/uqOgfr66p6it8SB/aR+7hP6wxd8vsFjTVME9
7f8LoOtsl3td3nAYGXbTB73KJIQJYvsWjQ1X8ekQeSjdnYeEFn8z36fue5zeIIqdNaKJE8YMAQSz
Haxkc/WVnTICPrMVKmLl+HNNMLasP3qEtOVvhy1wWq11OXmIcnKxpzybPSib4T6ssTl818cLvpxE
qswzSXVBsPh3qaCor0UZphN1v3sNXtbo5BItzysmNO4NfKxq9/x85ZX+QptBvUxjqKXrw9VLsdpb
Be3Yw//7uftaq5sBbsrLaAXNKUHp/qbNaKJgv0u2b6YXU1kqQoY7YN4WgdeOBcMxFEwP7AACYfdO
vG72eJo2r5SYM5GGohFAkT8YM1X42q/do5BYFRfnUKKC7NtebWU3jDUmj8tWrWWRKggqMSA2t5Df
oVYZv122+1Zh7V3C4Gxhw3F0FA5pxBMlFkLEIiGdlyx6g0zIfoyCSylQ13PwRTLfkyTC09eFaVIJ
kbXXA5HQbcNjNFa3UBCY5bOdkRXFrrpbMjCIcxz5ZarNvpY4NBqlpSwTG7fWUrZWW295JVdNct3n
6KQSbtA3603bhalbfqXo+XpOhHk5mU1WT6AtOLBSuF8Auzq0tHOspEt2iOdvZfNE3aBLFPMcSJDX
EZ5mN4d2NuhRbmKPl7N1ZFpMZkV0ExGqkWXOKJMLkd0DpecClABG+i/YM13vzWM/Y10GsnmLYjHi
RB1Ftn/t4p3M7iQqEW8l1zjNOKAjLCCREu8SQeTWmYIseXKtMfGKPtotIwo0/ayZQYueMvK6Xi3z
5c9CWX239IIR7CArcUH95/PQepPOQaS9q1ZiUbiA/fExtEgY5iW2IYGsxI1PIhPYyud6qM+nxxtg
om0nyz72mZpRUy5TZieFGptxcC7t22lk8nS0o5kPLEiD9/ZqdNu+JwvgU4V0lPT5EP9sG6q6zbp8
lTwuIsqV93dQ/XHjSENVRWHOQqljZMQFQaFx655qFXWPTZt04YpxZv4E0ev8/U1r8ywaCijmpvKP
s10d/Z9YZkUlC0oE1E66/6WAGxvd/u3Al2W7PZVwuGSM/pYJQpMBsCLhOByErzaimKTaej2doRbz
CIvCLMoFC6/QtowHRy0AI3gpr9K/rCaDnT4OkShW0km4o5LnAZ2D/WlqO9f0Q7ctZk1fnVH2HZfH
nfq9pmDAtNZ/ObgywT7Zqh5cYMkVqrO1QVvp7wQ8ghCcSDR1BBNoS+bgHkebjWN1/93Krs0z5VAR
W5TMzGTNuo3uv8PsuyWNIKIMxptMgj/NS5ePh4klNxcaRItPIypzYtmtxpEa13q0vZkRCRTINlsD
LczXsupjhU2vMMrkINAuIkJi0sHJ/P14oZneJiAanR9I1weUz8q5FaVcYEpdLTQZgUvX5+OzjTCw
hqaVWRGi4ymGnAAWE9Jt4Sv5tsOU0EGhfNwPF9kAlILx3a2yqM1I/W9ApI/ypdV37RS5rUZil7DF
BWxPQPWDW2kGOjaU5hGYrZYhLQ1pEUWygQd9Lc2A+VaX4wKu8ZJyuJs3UzFqpds7UQs7PsVhu18A
l8OGYhdzn4g5F6kZk+pk1ksHdo9MG9H526JCL/ogHqMIJ1JOjvis8W8Mg6WwrQrLohxQQ9sGIMXU
oqV/Mahl66wpjOgO7JMuReJB4XP/t0VcbtyclgCcMjdGw+aau5qWwqs6qIMYT5IM0LsfoxaAlCdc
4y5+8PiEAgwZFGRDKOk3y+E/WPk/Q+PHvLj0y0DyKW9SYckcnsaziZSNXk/3i7Gn0KJ3ipzacNRo
zXcpLV9z9nc/o8UN3YrUkCVp24isd8psCSOowzeGsc+OKDV6R9KiJycpWTvibV2peN+eOMvw6zbj
yjfENmf7UoIoE1RWoJqakPk65KajBHSF/G6lz2b7Wmpq0UWZXAv9Suyt0b0a01Kc7kdeot96XQSW
KwMVDC/5PeURqsk9yhhhNJHejaXbrp8EtiTdAqbejwbKTb3zyHRG+mBfePS0fXsm7bBfzOKqh0zD
dbKzxP4tqn0OPposFd5jANC+ngSfWszY7RsM57O3o7QCH+KNFMYeczjeAfQi9WXPCaoRCMBPCdFD
tdf4+ABifgj5k3E0FUxpZlviaeTb24f0Qg5ORPDq3vyIX5uvihkpMKBIuC5RNujS+7DZJaADdfyL
XwH0esT25Gch81+VLPk8gc3CvnC+06IBigvS79lkmVLIfNzqk6Di72k61JfQJyAOVx5KakONJE2T
/zC/cMDbjj7sGznJ967hX9UpTFJw6RBONz+f4qPLzJM7+5DJHKRxbCw2d+NXztRVa5qKIz0OzOUh
t7oMZmSWmgnc6mLUBDdfa/AoQbniKB1mKLirC4V5gfSehoDsGICVfA2YNODRJBR8RSjtj8fxKqc/
EbnQ+kdytJB2G6HvSrzTGkmBEjRLK67Q8olPPVLc3osSsjO9zIF4TDC8l1yY4d5RchWImixb28dj
a3tVN0r1zwn9xtEpQkuDSXmiJbmKfhL5c01mpM0IlX9I2u4IdrQjz0Rni8ThVwW8eVpxQhNC5jJT
z9iPTyGGD8EtT25IrMkUDZD4Gv4G/sB7tqLBtIKV/GkJ7jHxG2W6lx8dBulwaGk/oY6yTXj+ulxr
PvuOiG7B2muC/F59dPq1+vugwtp7rUupyZVV/r1W8C+aTJPEVrJLLNiZWD1f6FvPzuN92RL/cJoc
aZo6GdvVMNu0N6nDTUgFUh3qtW0jxWUP07t7zgkm2tS08KniXtZGvS1khYc38Jo6IpICvwa13dUi
C8sus9IBCMT+rBm25g4ej5+rsLclA/BAA8SXlgy/0jgYoEUfd8KiJFg13iktu/AqFWddTnrEVskU
SUG94sxLh5C/znjP7ua4JscUIjp5gGYHb786LTablMgeQqp1OYX7m2OE+xWc790G5qXjrFkvQjb/
XG2TGPYHKmD6p7mWLtQhZh/dg8Ywt2BYWv6gglRo9GUhFYEwjZRcvC9nsr2cxqh6Qybt5fpoJPYG
Q6XOYgsAcZneE+lLRo2IWiM60ZlRmtypwFwpbQD+KNFZHXpHzPIJhtqG1Qhw4YDvqjtQ2lmeRabi
sZoVqezqM9DlVKvofKyoGWRXAV89hcFXhn3CH8+IsLjXeIPaaeDODcfiWGSphShmqsOquf5OIPeo
y0qTUXp07CtFNLItSxeVMGd7lDBlhKHnnRu/h8KMceAMyjsfZHnpryKy/uyBmnBTy4yYih7k9M1H
RUOQUFg4fxMDkPuuRSGK3EjKalTfBQFlEqwoGracbhg1s9JlyMagzsHExiUiHh19seke5SuQQMoe
fEMnQ6xZYze/ERbT/BqcVhAXtzBeDcm/RGKynldyOQvy5N3R9LfiysxxkmhGgpLq6PEDPRAhyU4M
7M1wDyJrMJJipIV1KvgPawJCoSdZN/jp9RTyjj67I9++umxrpbAoR3sKQ+M/3S/3rQ1pHBTxW/QG
Jbo4tmx8ikux0SR3Q96RNK0mc3Pf+FIYifD/pB3uWPbkDXkw2Y4F1hLPddGPgARjYkKwDfPMU5Ir
oyGQ4Z2u7hl/P9Z5V5b+2zIzFp7q+vQD4jLnQJA9Fblma2jhzuk3z0o6Cz3PiW++i3q9QUocfRPm
1VumIMZndZspdLEoViA3+kAMrr9u4PWg+VKbUt9AtRmoVh1lCY5tYcRhKiISQwg4Js2llOJyWrjj
wbKhgkX2iqAgIpG5iDIye+WjAcHtIBTBuNxAzq3AG6cejn20SaPD1L1MstN9G1T3ftpwHW0rwr6f
BRVIsU1pZ09gKbI6J5hVLGzWw66vpKIgub1Sq99iAYWgj8sn8uhxeYuuCIXnCDJZQvhoYC2zb7Tw
2hgZnuS/3npLFxGxoDRq+s+rQRHPBmYjQ3qmre7ys8j6h4ufhtcIKQ4waXSTrIORYqcQrxZotnZo
cRYZeG/cM1u9xYFZC372r0Ph4cfrTI+Je/iCa3cv7HsOsRmk/0KgXgL9+3k1Y4/vO25pxE1M7voB
E5e4idbAAEQWQaR0bZN+TNxYuMEL6r+sa3gY5j379ZgZpxqjkSVD4yxCCJaTGQl0Imd9/0PKWOJM
gB0Al+GoHFXg5x+DzB3SwFQzt6uQ+criof5y0CntAx1YupVl3ctqkzWq7eOZ1WtfQCw28eDhcEGp
tNEuE+6h1Wx3XFGxpjeanHoGZJzbFLJVBzk+BfFpAr4iDs2GmJpTYGCDJ9rmRu/Z47aR2g3nyJ2x
BipJACL1ae05Ax32PPDwxV4D6dcugcygM6i5zyC+vRp49m9tifnutRrBo6rGxll7oyTzgFT10Cpq
sUl6ysS4HGRb4oFiFW9kEedp/KHQP78GfioucYcHkNsLNYimA5D7nmgAqqad5Xjc7SatayqOmqlA
MjFwZdZ/r/xeEtLghJuPxYqWudDHshR7KGR0d2xB/+giJ2WNudeFDCJW06rsE8h+UtVFf7H/C23/
YSI0TlOHych+VLuS4az+OUDiW5jmYLHTUm6bvMpQLiSOJ07VtmoXIWeC+Il3U2YeO19JUarc990s
pjdYnTBNfQMDAESa3GaBCADJMk+mCSF3Krsaj2Bh+CLG/7Zd7OGXXY+u/yRPg4DZ3YD/vc/wb0M8
snM1De4zhSW448WMJu9kjJ0a1FMhAUY0Y2Jq63dyHQWOPPI/2Qtx6Tww6R6/Evt8/jumzf8+FFxv
HUnWwSvylHxKCSKj+RQvGNFeTQ++bCkD16Zy5EyI+xEj50TTOWKNxZmssJBOnpuckZHNxJGZo0FJ
XNY8L76Of/3CW+lRsxnjs+M9HPmllY3okiHxvhFbCh2vwQQepf7Krm1W7PdwD5QRVJ18fFPLQMAF
3o7d6nLZSfj3TndJzTfnlzOHQKgwqSrGYj7JVLmJtQqiGhEvcs1xQxhxthAliglnHUhItEzfRjEY
yJ39zlpJ9LS2gpC7+kAm4Z+4Kp/Le0ydOw3YDwpGsTgdrRnp9Ub0/WVqUWk7v6bEpebrtU3RcoDI
BP8ROxdcOwUl9Q5t5btrFhSVhPKQjIpOMf0TF7Mvm2TgQdLKjhfiqrVIkvsqPfsyYnMEAprYN6JN
afBPVsXMCQ+4eScl8pokVNWNGd89jX1P5pvwGEfKVM+VdXzAagAI/O4khWdL5Eg11B9JgUm88Fwz
40yBlm+IriLoRg14SFbOBJEwvu3Ax9LOElutCfOCWfijvffQV4PGDfAyRgk1XnOC+PpN011E7pfD
Ftj2GYhWwlNYlAc408kZg9z/0u+O5zjGUcir4w02xC01+zTZ0q1KlqgB5A/c7QmBR50dbzW+FoOm
A+EO11l6n5BCQpdmK8Duqxzxttr4trWNMAbBZdQK1WDUJJ4MWdPRpBuI9hySPhgMv5qEy+Zd4NGT
dYwj36CzW9UtAdEwLUbrI7U28MEYdavC1tjm/ON4fs1i4DOmGkYVanhBknSvR7zRobpd4uA8FnfV
M/UgfupN0WiUW6LpoOLatbVT0n9853BJeSECCFRgnzwlQNjThe+mwVfPbpDW+pzgfMmhrmR5T/2O
sR5N1xzpJMvS7tjkgJX+bEjgRWueV9hMGIg3TMn/9XMU1mfGOTISzH5d5+3H1O0aMDRn18iEW6MO
hueb/uiji1CPkXl6pLvknHslbIDdNjh8Iy7rqYBgZpfkcIktkuZiRFD7/rsmaZkBRyiPXvA3dmZM
uEp/kWD4+wtChyvIOHDZc/JbTZsn6afl7vSe+3bIxiOsmZ32SprqzLL3oD6VKDE1WVlZ8IX4l9UA
3t29Yn2TBL90CDZQrhDN1Mt409ScKGn0cIot/CkRtOz2hP+3NUKc1NBQYISc6mxjBUqcrWf2/6YB
CcOWcGJLd98kn7udOLJ9EFMV4J80c6LXxLRXCnjVpCiBbN37UScErZnweGT1Gz6jEeXSrAIHrqDQ
ijO0poncLZZg9yTADt4usBwgje4bjGiM6a7ZN3tGHEzNzsRuLHs44eZ3P7Jrr6+kmhAoE5d7mNER
wLwyxTAcMEYOawirpJDs3zxquwmJqhaZViccNGqUCUnjyslBhbaTNtdv2L/w0JsPVdmJkPyNpHtQ
jKx8bM1q41Ngk++qjfXlbjqXe8XvEtqVAg67z0po2dhv+jE8rv/ji18cCuIPfdWm5zUN7PX/A6IL
mhI3504I0VZ2Hn5mTaYMm0ev8CeQUp+hiDGqI2BDmjn3iu+epmOT2zeZxKtTLyF4mrtMko6Ba7my
E0u5+R6avQdJ8zk7TrI1YWOJ3eib+Sgoxwh+1RiURv7N+7s2arbDF6p5hnGg4rpgTVe1eQvwXDz3
Mg1jKGXFII1MK6eEcbch88RSI54wZ12YH93ZvJ6utaj8qYKEQcztDfSIlOew4hoiN3lX32jkBjKf
VQy/Nbs84QZU0hbDg3eRAjWW2UTUpZHvaWXMOBG45vFG5IbTfR58AGY6vBqJzh3GlbBTfAm3Vv2R
g7bPBsad4IBi7M2hBrXePqQOKGgdrIqyW9R9QyMTTWfSf5hPa344PNS5t25Y2fPoe89nDp1BUHmC
TKd49VYb8ogvuB6uWEq/ZV5+ERnF8yH1ugEORHKqzuCaA+rSfQV0mZiDZASBiQ0xQXEKb/aRjoUh
KaLnz1o9toZocIa8TG6YpjoRzluN9rkos15C7VVCsbyhEvmjFQ/Zh8BpwDa/WjR8ZdM0tlr07aI8
/sXVK9xOfxxRU4+56ol2mVsIOsoar2YBXimGaAu8ZVExcFliGVDwk76v0NVcjnG9OaqaWnlFEXHK
YiO1RnlPpp4BWehphJNaSVN3FBeYKh2o8xBAwNw7FkyC3WDQtqfqGkn5rHHUtpu9w1cAJDJAeDpt
F5Ij9CDDs6LQwD7rn5elbpBKeJ4rxWjktl4KaK9KCpY1ghPNu3B/T67zRLFG52HtDshaQ4BLkLpA
gl3YO3ztX8RqDt25z72RmStTQdFpFTkFmxs3UjlBooT+4GLD/aUdzsvZIXcF1pRoR9VMJkZZ15zi
m2aKpaiUhuW4kQuCdIDiXs2WaSYdn+7uqfZWiCHKjK+48O1dkEe6IYnz6vwyS7Rn5IMj8ctXvfXo
EtcLP6SjAhujxqACW8yJoKhaqdwN0iKJwh+1NSgisfk5V7g7dICAy793bzsUY0IxnfTDFuPb2qU+
HdYCVK9r1Q4pAFqbBZ+gCVFAcJo9gWN3gJwhq2Zz7kH08Tn7+WJ9IBJ2UcFLyK0lQkYTFo8BA7fF
7qq7GwttIZWjADGxusqcs8qVRHoVx+3gifEADiwAPMXYIXFsV+9DsR+ZVoT8W05RmJgBoCHd0G16
e1DJ7nHr5lK/oe51fmnEYvYzr5+8CaS0pcEdguNcl6yepPHdXEB/9PJcPkagCROoJP3+5Wxd+I+z
EGFmGtuH/xplOWW9MzjM4onlIcVbxt/03SJ0sqHQlp4Ihz1EfZkXO2oiuP1pPlfQFBsLVlViFD3A
VriFY1IKszJ+uAQW46/hp+ULudv2FCcdb2dazepVK6lSfLZyL7r6t5GpDmnZS5TSXJYwX2H9mApo
CjJ+c9c+/uzyvzCUYAPagc0V+uLpqz2+Nbpm/QV01ol72KMtirmIZHdWC3wLegneKBapuI1ieZOd
W4DVXr/6Rz9G2xpTvvf9lBOqhIlISTstRPj2QJCYq+hL2jKrMoiWp/yXkqZTRLsQBKd20sh4dh+q
ZGpud/4fRHRHD2b6xKlMmo5G/0g8pYnK0JWwhLDq5w580zkR3o7T/HEe6CLw2Xvs6ndi+o8X5UcS
t2BcbzbKvJL8hnV5snM0vxbbu+5ivWC8oreAaBkMIienWrCA3TyWgksOnPdD62/35gvg5iortDjN
fPmTHVtEZqN8rtXSmTgRZrl4hqwE9nzwOQeC+QCDXohX4W6n7Cq1TCTHA3BTrEotT8xXFgHZO2gj
51DKysk+awRYPb4531qVmeC67Ze42G1zsKqtxc2eurZEeWFeDvgZu4ANlfNs9TT+PXhSw96HxR51
ZXpN5BEJZqJzAORz1NE4Zs6eipo05HlMUnY/O45xNTMYZ2DQNJDyFKrSIYfhIekKKOz1T8YMoq4L
d2T8g32fgaXxmKd/gNbZg8+HAbYNXnU9UfjdF/euzbkFLQzorhq7o1Fnj+tVHtsNN+Qn+PUk6dRF
MtQK4H8u+3ZUHOWR6CXgY0/52uKIRBwDlT7rFwUTVJs8JDvOSp04/HwxGXd7C3ZqU2607mx1N8E9
HXujbfQEajd/SiY9ILzZkr/IdBfOU3I+XEXLaWhVUhuxyVG0ILUVwyHmbR8WJUYfiuC69fY6rkT1
bzm0KC59EuiTiIBc1zmPjc7XgkoClPKbTRPZo5bQSsTUIu+n+u+lcTjfOp8gpFIZi0xEYmy7wFL8
eZ4HkEndqGAkxmeuSrK1fqCKGtc+RSF+lLlQfnpI4w5/D64U6gir4npmVmr7/DTxOScK5hscqWn0
jYevlWyHo2Q40Nbe4+17caBDv/pGc2W5xuHSclqvKIdm+PJTFobDyWpmPIh3cQ9JEt9hNmNM6bzm
OZmIJ6srn+l7Nlj9HXecHUZ9BO4eAkiVY7DMv5135obGWgRwmLVsG5l/tk3Gwk8q9rsQ9mgVnIJg
nKg/i9UJuvUX/OWDCJl1uZ6m03z1XpnNQ4M3kRMuNAnwRpFJjczJUjd3WM/KK0c/8x0ktYOf55m+
vuKfjO9OAoUL3tz5731ZqCroaVSK1pje5kgNz09K+xRjdD6iS9LKx607T+/YQgTJ6CyOU7roMbXY
/KjVombAmw70E182aD9KD+bjMs88CqMnlTLknCGWpnGA2e64BJ7Thb38HCxKO29zOLBd/8Cq2P3E
fL6By7DoPm9k40X/UtTzKi/hbP1cllumAGkIHfNPbzyUFhizERXegObHDSb3st7NwxZcATWOgLqW
LJxNXcnpDIOWpE2KiSiFzT39G9SWFwXscmiYN0J3XENSrBtSTfAooPWYX//ZGLRr2fbceb6OwWgX
ZbcbnqXdNyi12Gyyx0/D5p4l5gpW7X3ZoGosrf1rIZSWWgBbabXHotoKunektKZFHNd/C+DXSiZY
CTzKnwNfyfR7ppu+HRaeep0UpGZHipJkc0c5IRpM9VnK4ZFaZFJkqY4PVkiqfj4pwCdl01hpQmyE
5Sws6CJ4hb5xeQ28tOKtTMGqsUFtEsAtNou6H/Jjip2KEzNv7Tf10Xgeu9UbB1dm70EyRaCan2CR
XhIviYnvnK4voYOTEziz0G+2WMOU/Vaed7DPjuPpGnfwehC0TElZNsP0TC2q0a93ccvsdKtf2gF4
RDsetqYGZlE2x/PrzDVR3PdV8TRoytfSDmGhAARyglveUOMTEwUQ3uK0nGJQRA8iSrNpMYkzi83z
0Emezjk2ndnSpkbzIofLLfHKZWxlrI2mlPi/qCC5IpYM0L/ne4NiGcCe9oOQBdVV7wNlFgAbB+5a
Sos0qKRmfEa1iHgHSHh8nPBZPYxEcnjjHPlr4C2nATG7+hpi1/w4SByI+RbVk4qSSsbB0gsJD+co
Rh4tSnrZ/qwtRG/cmAw9EQLm6pAobV5gFoIY4+04T/e2XLw19T0hn4hZczpSd7xVBcMXB7KBUTmL
JLbEmO8u+lsMP7n7yJp/y6dk4iDUJeXioO6bz2WMP+POkkXIT56By+erlPBxJ7/sGD2iqqcc9ATg
JHOeKL+Z9KekcdHw2eSZu8CNpDjzQjaGdNA/Ew/tDPmN1XC14gfKbB71g5H5ODSFdsm24p3ED5Ul
ZdMa3DBdUNYOM8BE6/czXPC1xFXcnsX50GZPj8xG8xiNcViXe/bQSAmMJd5+nRpwWu3Ef17EhmAW
Z9rxJrwkKSoiyqNYQmPdQdr5uWLf6p0QQaA+xlHAIHHtPbgucoULkCoT52Grmoni0R447ql3G16N
MZlFupLk2TkXT+5fAMqEtFJ7vDqC4ItIm7ZOQW0GXaZfJVIwgIMD1WB1+XveRAXSWYwT5I9YkWCU
kpj0i1Mvtx0qgPpz7YWbto1IQiWohmmcwUbSne5X7R3/WaF8mRY73Q29jymOtPtetN0nWdf9r3uy
soE/j1MhABSRSKkVema/TPNE8ctpuYXMon0cnCXqLY+e20Lyx0EnlepKdXVkYaGJ6fNKsMKr+XyK
T2ADdUHuhJDQQaxdpk2pBe2tW48tL0C871jV/0A+7JAOvKFavPJ2QxrPUtl9aUeTNc41QiIN/zgG
IKKj52HhCvSr1ndcztIuQ3I4csi4BUzG+tTOj595W7Vxsi3s2o9gziuV0FAd2Pu2YeIHhznCnKBK
EHSSgeF2cVpiRnSigGUcerPX13u28pap9XBmtgwiB2NfGJJUCzdGzTkGb75QQfZ6CVMBTZEIgl+o
heOzpQcy91RFBSFjlw+kMsUS634pvjUFcIo+p+RjRYfa4Z2A5n35fyhnoaQ7LqmpmdpLNtoZRwpA
BERUHsAlPiuSjwoUGWdp9EvKLPCnOwgnMUb/9R2Kts+XLcsZN327MDCmyWuXJEMTNHbmdLM7+DGq
VwFTTHivKwYEr4kk45+dCYFZ7ko0MknWFrKdwaHcjTw0F3Ujci5xvVGwFap+nTq6iQWEABJXLJrw
vL5ZzbsXxbPpwtcPXvyJGKnGffrtQ41jfE6tidNxmMcs4EH6C8bnjYR7L8P/cVh53vov4O6CMhji
WFuC4h5vQWqDS22uMPe+sd//n2p7ISdC0MhjvJhHlIA3RL2hI2C1DR0Y+vWdzT8/JdkjSKdHfEUI
5wVHGN7zvhT6hXPpzGxg6lcZ2x1DNKkXVe/wV/1GmWS+NdUr4/XnoSnKbTX1RqKeGyrAmE84cX5n
O0dz0Zo0uqOdVB2MEtXtPNyqe/XoOZr9fZG0F47KRuRP9sZT0o3x8i8X2dcOZvjBZVZ47FijQ5+Q
ZRd7UuKU3pdMlITJVb8j9yzjLwvukuvUwDxZCtYeeXVfmZt6ENGzDGODiKLPgIS5JuTzdOY1gvak
+mbvUXZc4saGxVNlzUiKu4eko80OR2fEJG2tXPvw1ihBCAq3Nl4HqVqwjnF0XQalVL4EJ0SM30PI
pFDrHbenLZtEKIcH+Aux/hDJDzsvYMHIYTRjAdSlGjl45A0IyDIwIPfpTlyOWpZonL93auWFLrYd
WPygoD9i9uzaYkjgH6LvZ8EytFOtfkeeKNDeUNC5x8LtiJXcViA6NzoFZnZFcqCk7nYg569O06x4
wNbpxVIkAo0wu12R33Mz2DDepQnK28PIhzGI6zksz9JQQ3fw8O6rpF8k1/NvGJd4Feaaw+Jnw3zp
y2r4aAbuIgpFRixmHmYNTny8IZAFwofA+USyuEJqbm9l83ZjGCyNZD68an08TlobNnzCF0ObX62s
9Lq/3mBG3m4TWwhT9KZ1TDYNH/wC6MOvP0HDwGD++irafQ1XoINxFXn4B2aN8Lg3fTrhK+hjjqzc
1J0Cp1pYwXw7nUYfGoeQfA0+eOP4cLl7PRLPStDnTtqG44rBBOwR3IDrHRySM6Dx9qSAUL1WTnil
dgv7OnRuqI5ur/FZQLY33fSK2ptYc3S1TWfllge9EtKM47jiZ1ogDYI58OAPJ4wVNdjGsJjK2fXy
R7B4uRgmoeAImEl3y823oZIBZwQ6E1TKeDsfY9TzBziB0LCo1ulZO+VethPG0OOqbOPK64FiW/q1
2pzRktgwPMbqRpEpmObErT3qCmfOxPPLKmay2k4Y01Sz8L4Le0b9NhPuobnA5KaMckVN7Dca2rbz
WZDuDp+AVolKWzBWhpOMqt8oTq/qjNdV1zAICl/Lo0mP7pvG/LM8G0WO/uyhhy8U2H8qqAHA9O0S
sPtbQogDC8gwlbGHqP4OgmEre73qR8YBEhWYKvJvQ9/8o110SDzd6IlbSkLjMCWJI50ZnUpYgmwA
wxJZm+iUxUh3JSKn/v/7YKBQKf5Kr/zczKXMs6apsRXrsY/nGKxv4LDyAvJ26P7/1mi3W3BvNqTq
BsDXMgZr4BuOQhO/KFfXvs3MJEyCCH9NzX4l3Ty/YBKTQ/po8QBj+DlOQzNvgj216REz3CJ63oaw
pY4Huzk+Xn2/5/PhG1m5z3mRWOkEI2tVZwapL1Df/+n5kaDryeFlLpYrhWC9qccotPbB8fsZe54M
kACR4GMjFK79+r/D08wxmz3puZ3dAEuMmnACSG24qR8tTmdZpAsl2rchDJe4QGY63BPGoXRzRYT4
lw7XXjmUsDbFFOWcOQybkhnBqM1T0dkiM5yd+H7qNGk8k4wK7bDUq7avoVVi161yRxluRsVM5sUM
2ALcpqv1NksqYDPHcgvRxQsPtkrk3Ep1JAXxwRR4a+crxSuLRlFtrXiyP9fv6Ix82ALK8w9e2LVi
fgu+hVXR8oGU/1pIYqQu0XiVw3+Ff0RGs4sccN+P8tAcp/rLiO+PVl2/Aixm4YVjMBh7YoLdRuSU
rzn939DoJuzkPsU/wftNrxlCPNp2tDZQyLGnNrgR3yBDuJ8aGR48a3abx8c60RXN9gfoJ1x1wxu2
X5CY13HQCKZuqPsVCcYQEay30BhpRy00I8rWvmtaikMQmcNVFRR7UiLWHsZ9KX6GKeQm7WB5cz0Z
8yJn2mHpd5qRDwSpaE5QIpp80zHSmXWdFdxlWccjW+YD1RvTpAAj+dM5ui51Vkv3PF1a27Dk/RUs
630PZ4OOsIxLIuRif3L94+c3cwWM0lLlzmK3nCnrTMXv8wYiwYFjatDbnQHpmgWycLeLY7dRT6tC
6v5UH79Z5JyGqJ263dDRJVQ9qxPaWe6x6ONXT43zd4s9a42xaEUsGZQ7jwE7YkXzCOG9m6RD5Vfu
HTzTlgtmHaTb7OXgze2Lde39dpfXLQc1uy6hquDSrYkaNKFAP3kElVaPJUAxlukSfX/qfARw9ZSA
PLiDuT4IAEVic3J9uqwsh3QS/2mHjKFUEQdsO/4waau6y4y98AEVEe2N+y1TJRvQjxz4WGFUN+oj
/V2EPIpmWSukc8zApLT3EpsG7N1sMHZ+/wbt2zHWiD+DBmXukSsIsbWPE6R1f9Vd4exNQaefvbEw
X4ktFtH11gzqZ1NSTfbZ1m+SY2YYEujKE6E/AmSPmt0RmUIce+44kf4830Vcjs0UjEqF87ObzQLe
Z42sB1Iy1EGY+P0QN1stZY7lvXsZdhmaM03FrXGegk0VRQfY2HZwWRsJ/zQUh8cY5veE6qVxKV3G
9lOAf6qrcxWvifuRJLzO+hTDuzpCLM0qOdfwEtAsG97bTHLBmn8AaxViLK7ED+dt7BHaYcl9eW7h
cPSG9Ib5zRtE+0lSGit7ga6acuHqlWJNCiw6uf6DxQb4wElYTRWoX8QLU3u8ByqdEDcl805O+paT
vAMAHdsD/J2LF5BkT0ixAaQr7fziR/9mfX/GRpiMqMd3WSwtqhB+63MSkVoZXTU/1h6BN9gk5QsC
9mclK51zjW8aX+oh11GMLcpIpu/ug8ORK0zmz6bdQ6TP4b6+yI15uNRE1wP7lem72HOXe71vWtIb
wS13tvPtQ18+40B5BQMaDVPH/R5FwHH/mMu+wDuifJmQf10Jgkk1n/5DBcDsvwNyUgbAlUwGc4g2
D5g8l8iMzSwWZ/Ho368mQGyH11sdXjXGtcrZf7hT56XpMMv+iVylwmckg6MN+2GB0+dAJ9AtJq/a
UznLC3DRYaMO9F6coOlhV1SpkoteIeDflAtliE/9k1PCr65HcQMCzAs+hH2dDc9nohdSJT6OefvA
ohxGOmk4GcxK/lS9O+b1E6fyVz9bz1BDR7Y1ISpd28G6VpaJR/porsWaQdJs0qPbFj1dhlGKlySj
DV0xZxMsYR6QvoH8lSg5OfBPy/BOs7oEjpM31+8wKoJy/mevWOAWcRyofP59we9pYbk6k4pzrwdP
3Oo1fZr+py6C2Dsln+bleOwJTYuL7SCXsYwsrI2DPnjRGHmktXTQlwd6enyJl3Uq+GkC4S0swdZg
SXjAxjSUPwmunTvdKAIEafB79oeP1JLKqy9eT5fusMFY3JrkOuYXsQ+8vDZQR3KNT4o+xpb8iO0S
MviXrrhvbPEKu3iScr54KbBDDCoyxmgzivP6Fe9ia+r1eLWhak6j1+hQfuJmtwaIUQGSDy23Cw/c
u1swPi5Ki2ELwup1rjRsYyRX3R5MKsyociu88Jc7IREvXqagSqTbf3dYMnSkPC+dF+JN+AjEOFBu
A4+PuAHvlX1cyB6ZU4JO4LA1uARzr6jwzXyiSA87SwKXKl5BjwJ2oCqvXuYY3QukqmjUt0gXwigs
cQsesn87Ijja7Kpo9taDAxE3ukpofG7yoZCSXv2slFZCw8M1/DwwBuZ7rKwmnLfqxgyup+aS1lY+
7SrCtKzw020rgFI1LwnYUxUqs6oDuAyzaDO/FSjS7xufk8UsyoznTOBmzPjCMS9mvkCZQ5vzoNds
iziHGMj8T8mjjgzRQjByx6pBfD/HX0BPAXrrFJLwpL2VwZFfAVfd+2miSg5fVyN/wU9Gx7Nak53k
5MQ0dlkfeqoMdf5igsOGFTD3GRMDzdFdSyHFJbfsX6DgTO9b9KHKFIMjPxFrP14e4+n0Kfox7hnk
hbrPCdAp5Fqk/z2XJxJqAFKEIUBCXvINQf1be5pLX6viIvrPQigPxA1jjN1csmuDF8RA48MZXQEY
r9M3K9iyGAh8EbbQzT2P/TX4NPqiy8dQ47gfwBqmYcjz3uMXfhol3QBNsocDH8vR4qyeN6luRm2L
r+ZfswSSNlcsRLho0ghb8H9JM5YbBf0D+lTe5ph40s1UkkEOMYkWsvstSoonVlXMnhfl8tooFE7p
d6hlSsmE06hXEbXnfEG0XjXzjBQ593Ern9HXMUM168tqftxqKbK71sAif9BC/WyNUVJbPaLL3oq2
x+QLd2gWpMcFgn5wIcsBCTTqYgz5UqJJ9Bth64lKZBwxRn/ALVl3omKeyLApMvNlo/FToiAk8wkT
9fS1YmNGPqI9p9YdBHzUZWJFX9Jh3bQL702KqdedMznLil9hYt6Hth+82GexnykLR8VqHwPbY+eE
0+kunVzzIDz/DcEnOLDDWwELbqBUDhzvR/D37DmtQvHQkuP+QVl1hEnSVDYZ//eoZ17bo9UmP7W/
OJPWomPddABJmmDP6I289LHGMxklu40akwSUMp1jkY3KgLblaWPvVhFA85VDBm4ZAI+JV2M7HwJ/
XXKNyp/jE1tPN0pbkV6cES3ZuNx3mDwZ7O+BvvLCAX3ORACqqoQUzE5Wa+neFebXEcyKImRkq+eF
WYMaovxEf9tgpiWy+Cd7PFwJWye2iYwYF+S/tIvnuG0gvYb3YbX98F1H3nFr8xEe5JT4bfvgxV3v
yPyLLF+4MDcHXOy8l1nNiy9yYZDzFopt1ILjGKHOVv7G0jDZllC4g9N//Sn+TfmLftotCbpNjYe5
BOgjK/jnAFMjf3gepTx0V0eRmsSATAjTcIHsLQbiYYz6ZLLoCROrDITmY3pZ5AXCbb0Tzd8xEI+m
hCc72kppP2cNGm00U5RSWU1BVtwQ0oSeoLqcAxPfsvkbTn7qx4Z/DreGP2teiuWtz5kZnggCNsCT
apT1gKYBzZZqdyCezRfFJPSjRnw+PcgzKUf9ZxcEy/ulJ9U5oWBV6/hLB/dHKz1jzm/8mNTSbsEO
gtagKx4+NTkKmLukk64i7mV1LcNbHixTttljctPlfhbV8AQ+S3f72/h6fVtq55srVOYOyNLKf0TC
k/I8psdQn3GOvZL8OMLzeOo3NGROPzbSKTp45WA4C6Ed6DZOipCRp1qX1v0OtRyhw/iTNeMwJOp9
LQ1HYyHd4H5YuJ/Zw+0EZ2fMw6wcbVYH6IDCSYzDYkQqxuONLaD6K1QTdSMoUm5sjjoCrmHtuepo
oBhVI9VDxFNOQc5DUwhuuwDMGLeUeBA/+sD5+D3KPNOPuFtZD3ad+jcQupfK3HatP1n80p/n4pKB
yj6nKC81e/n5uZJDHG1qZBdjyuMnKxQN0+Z93JCaBuhMKa7cyo25wooLHXW4uvLCfaTVK+rRRFly
x6NztfryFMhcR3wFq4stThK0WLYU/cQHo1csbGF5iocfJnwXNsx/4YGnoVSLCmlkrKrNy6mh2vJ+
rs13vLDgPTFMcUMQd1rId1fdSoc4QSLrYf3l3SSo+ncsIp3QyS0MkfiNPR42oUH4kIpFPFgLre6g
JlHivhWBemTgvAKvJuQ8nnULu/3NALTLw4E0RintQvQEtLzeS7dR4omWQQlPenGkJYiLgrEFPmAF
ZlKfWHSyf5HLwc6VK2WsQKtrTye0tlnXPEbKbrcFOhbqiY6it+fd/o6h7me8VpCWYrLmajZF66yh
Ecxr3Cr6QNgq+qZ771KDkg93gMqgkV+oW/DKNv+9ZTuwovAN8RJAhZvM6jJotkdADTKN1vNF6lQf
0fYDSaZiLnkDazG7Nrkqt4pI3oU35md3X05LpG7xW4BfXiKQ0Y+RhN0USdtbp1b/n0+mRswhm6C9
zfTFxPtpyYPLo1GLnzu8iEAu9IrMb1GEDFAk5+unijgUkRGJwb4Wc/zkQiFIxux5fagIWjLtOBWl
yCIyWLh+9cPKq+9JpCx88baLPAKlAM9jTfl2or3Tm4E8maFITAH6EGPO+gh8C8+Jc9greeZlZGhd
CnnegP+as3PeucRXBj6IKOvv+OhHgj3z5NTNYndAT9aGOgyQj4V++GnofalxyHfoO25/1E8E6Nag
HQnvroefa/s0pCJmgHYUKbnhk8gKTTZgbbkMntBPu4LzlEszbJIYnZns59gkR0tDwqgIGfUoF52Z
bl/bjlaMN4VZEPed4mt4FboL3JfWOMyl5WfMPtJb0YAfm5dC1EovPS2TEhojMx021dAB5rZAWqts
7zc/O+C9vTF3jwQdOmgOmicMaY81JRfDmtTqQVS4baV+y6RRXWiCzL4LcUHqKfLI+DAmS1uLuA26
+XTYQ7CgoOWBMPLtiq9+ROsbMg+ZxDk9T64uqm+04JWtiBGUqd0k+2eAAO2zEHGzNGKRSG0V1q/V
e1A6vSBBl/6L8uszZEsV8lcOKvm95NYEmXcp43U8/PX7VO/wXEUNy+vp46D7FatcQihPyxVZTM5T
QS0G2zBfBNgBQvaqUW+pVKqs04rajI+2akj0PNUoAjYhT6kXQIJxVcyll5a/GX8xEyEkYZfeCRy5
51EVmZ/hv89tFQn9zmLX/2LDy0BpyXj14nbWvvA7M5m/e8H5jTMT/loiYHqE4fuzXSgJnR4k7Acg
2P78kf8XGkaunKrCFGcrx0hFTr2d7YtgzRI4ycTzgvgpSUQotT9Gnp+qa4MY5D/OVduy/9ZjXNau
ix3iOHmpK06whvydGj3O1uQ4iQ7iasxdq9lVBGDMDA+yE3ud68+sr4erkl+GcnCkMBxFQqX4QSYT
tBVobaERtJ2dQNX+BQebTOKbZT3LLtIHfCpR/OZT91Uhwz/f3r7dDXaEQPKfRenczCsuu1jHaesj
d+ISIX7PHsBMYbSPiMpWONPPmMY8tyvwQ+Pp7+VyaDB180Ig41jeY/Jn0IrdH/+N/JJcOhbW9TWg
9fwzaw2sekBSZ+AjEr2HzRq4nqBo4FnRWzf7QJl8LEv7Q3LlaAd8TnixXP9dZNjOGrixcknNYKWR
ulXpQKx9J4YV6UHKdzyWGYVqgDtsH/CqT7mLFDAQI6heYX402FZQRQ41NM1ghOF5owmRYOzpR8I3
81lDYrnioURYQaxNJ2OXS60OKD841eVVBosU+GNwR50Y85qvL2NsAPy4GgXnVZ+CEl/s2btWFfKs
P3lgYtagsyFnevdHV+e+xWANjcpxkV4KgUjS6QooZCdcBPTvEAQoBJo3Tiw0pm/hMMoymoLN1Jbr
2ABFuqVc/0lgnRI3tIBe8Atr9Iwp7XoNfBddBPKyjry+cvahJuH92WBCyh0GiEmrnR1nlAMkdWsG
QPd9GK73dmAUMSuSUGTM2bv8OuvBD0AYJF1YZAeePb5qfsqZT4Z8ABfiymB+HV6NOoLjNazsu1Bx
pDYeuR+q8C5lYMUDgdYepm3Uta3b/amm05+/RedfK/htHNa8jARyY6oQRoCLXavyky4Dnln9lbJn
RYht6lYVdCDhA5Wj2dka25Eu5Lcrv6ZlRiy5mCG5Az3hx19cbG4l+v5skTGEDctW2jWd3hte3RUR
YFVRH74OY7zax2yUQ4U5SktuvGBEliTm6yavR1sZjoMEaMhcSkc7KMJHzZS48V6SoNsrpxEiZhbc
1GRjt2vXnk0HJC+Xpy/RStp2S+qlDiaAGziTx+kaFt6HyDEts9gt8kf7KftWjAbqmeCnbSXQyZA6
qwGNZkIbD4xskvdUAWcJ2mjKXOoGoV+If+gZFIUF3iICBHk+ItiQdT2FRmDMYXuDRFEl/MSsYLzw
EOG9V76ujVWCFRng7p9Qre4QBRCuLjPC+tkptaJH1p8EjxIBziCrV36DjhqCJq1d23AQmRfV0yy9
/rXN8CWRc5oqTdutgBqacbFYgA6bsYDc86Sm/I6gUSIOvmisR4EjEKtKE8tCRVX8mtHgXS1BY8p+
3usOAsEWcBk8tJEfRdLsqYPspJn/uCiOrjfCZsaUmDGtb8ZslKLne4QDT6M6+PytrQuYrDjG2Rt4
4RgtYK+/9QJ755cg8xPchQpAAWXaVNk4mbtMNQ73pFUv35so95zkQjiTFEKo5kwJk1NgFFkUydLr
ALi+wYBukDWHpZ47KBispK4F77DYUv3AieWE7Vx0gOlw9cLZz6rmxDTcs0cWiAQD0CtkXL/QspoR
tvImzXFnx5Zl6xteWNCjofhnwoSXckxPI5yhGQ2sKrl9vLmFQhWOKrfSJQHiIgOYDVHvCHKqwIhn
zIx7VOXBJ89MHY3G3JpeL9gYsMQDJn+V6ouf3N89HucleacgS4wp3CWlR59sFcbkAawmBAB5Fyx7
rgADB3ZaZR31YfviVgCmaKsiPplQCGYKtlslFyxJxYvg+7QgwgQWCGsLDT/rDgLrCmy2tnp/uhuS
a8HWijZhF6CERo4sZrRE3ciJ14OYGOE50JFcF/qdXrvcTnW7Udng+MkI1LbW3FBqGWB7gJqyYuWU
f6AwAGnhNIHgxJhd6ucEAE6agDXDWylsARgwFqIIdTWFxW47Bo2mTsZ9MV6MrPOvxPidCbi7Sa8q
Oob20OWSyc+QPWBkz4dOeOWfbzu2s/3SRLbpwneHq6j1Ed9F2c4wEYOl7rFVPiOnae5O+NBYDVb2
09U2q5QUNUQNU9yij+RWnxuufV7GkqwvtcLlLR9a8nOtjAAnDimAn291QPJzjm3X6JV4nNqL+ifB
MzkMbSjvgOyUx+2K7ykhel87rtoQpgtPo25Vz2HOR4oUjgMRr+IomodgmFXuQLac4kWM0MjB4iBg
PGEOKhdc1Fi0SHhXp9l/jDZ7OztTuDFIxpd8txKgCbHTv+XdnfZNsNE+3C+kc9IAmumzl5zJybtZ
nJvTbqNHkwZXx9Shd2XRSvvKB3uZ+N/h+xwasJaE9QVI4Ysimt6pX/JVWFCw5qu4nfBwGZoRmjoB
e+YmqYK0Vb0xgE7bB6vMp5DxNrjEeEh6FAjZObjg3nROVq+XXyQk0Ymi2QbgEAdL1X1hvSPdct8s
XDlKNC74f/ia6o8wgjSXnSapTmr8L1ohTwkCd0AAFiBdEAnAwmfhfqsnvz47t62kySlRr87m1v1R
P9XKyOIYWckxS/IJm/wPrtPZE1LoVcut8WkUEOeazcJ0gVBFuVkbYfgIhodZfEaGsS2dXoKN702x
s2AniSiWAqW2PE8PVuRCbONZk+kNtlecFfHqxJE1qBhZVacANJo7OU8Y9xebKRdZhgiJnbFZe+OU
7ylbVgV4ww2SJHgRscgDbJZK3LtZHtVPfwEaxLnyj8FiBcbtNqUYfaK83pFQsUFdB9dlaVX/RC6x
xVeOlGIcB4o63EZzK+xfZwB2Oxmv/xQrR+GVDJipTF2CsU6WqCiA1Sdk/teJmTTHiJ5mJDt1CnVw
T+7YAen8Nq3L6rS9F/lPOat9F3GZole2SVyD9vUPNmJ94SNYIqFHMrV3lAqAHyyB1RBKw8us0c1Q
lzFsykl/hG5f42IvDFYqxUETxvuBk6gDEo7Ouft1+t+ef/ur3CJpg9zh5+UM/G/giwvo3i8U3Ycb
FiTeR+DdTw1wDZPbRA/6A8HIT4fHFTAkclBFgFzSEY/TwaJAc1g8LY78d/DwxZ39zOIv5EHCPeGq
ELThS1dCB+w0xQ05T91tsQHL6OdceDi2omdOrrZMiiRXOcQGHtcJDLpryZaAUGohqOLL42oPV97l
8pKjKgIzqY4vOYZZgmH/s9tb1ofPFv3xl7eVYCYvXi60Q21ATPo+VKQbRMZQQ3TQ39uXuFwCQxKP
erGNPCGADUQdrl6ZcLIThDDAsXgz0tSnsE4lwY5wRpyh9O4xjlb3IQkMEzPgoaD2X9/eZkNHFX3b
xv5nPA9G2E1gEV1fu8WjHFu5eCCQberG8KHGbCca/urshq5twYtMx2VppiCnva5iy0ERaQ/b3Tk/
NtD6o4KJhcoTg2ODAA9oPUQnpLQMGvFCQfpERqaopN9+V4VtofT99cRBoFlo6kcRp0VjxY5c14zb
L/6fTFyaA9Nw1RlHENXhK1LiwrMdVO1I2USN7CDRJfzNOPvh+K254V16tB3kQJhAsmByVENFHWa1
TF+HHcXa+mEKZriD2cLDroPrNdncQDXdgUsgzd1kKq6rGOmNLpjYD1yjfhbu+tEShWQqBRhEDvSr
a0BT3+ggyp21zjb9QbXiqKzJqq0594SRqChYQUupZbPBf6NcbGobdaefbaY/u9/ZDFH6esn0JSiL
QWgZxZ6SMox/atdE/9YzvXirz6hj0gj7p1I879E0DsXzj7VBTU7DcK6dTPC3S0ZBM8f9IfHZ/tWZ
SqeR9yiyTeUuICNLidS5Kdmf6Y4f0CsCgEKxAS9v6xR0YUKG8xho9tfmeHm/Foz5kSOYiqnv1zff
OCUKW1iYhojoU929LnfPMdWfB3VEdQ2xQRve+X3XiKY5QA6y5eI3qAViNzKsPE32ouRmrivNWuPF
OhUydxWNfRYNVqCSCA+6eBfSDE6PrOQI82Rss9QvPPwA+S5hGQCCVmtuO0urXGhghnz1jteRYIWU
YqDgSsPlkAIVjEELTzhlx4o99h1Yx1+9bgBq1bfp09enuRLAlN+kSHDVCkKdvCiVPWRF7h97NEMZ
iHC9Yr7pIf8zk+slVB+pyYV7VgO0be6TqBuDhnU2ivcKh1wHQKykmG6G+YLrDGMoXiEP6MBQAQM/
87TmnoPgqEvgxh4I8UTchAv/NW2ei4t05/0c2m3fOXapL7xv6qWmj7QFlPI+MKeeqCU/YedYn4zO
drcamI6Pn+tssoJuyUO+9x6p8kmaOtBwDVNTnE2B8SHiIsSLrWFsWAgaSd/MZLiiyPNph5zpDWE2
hh5sbr8kfJciRzQBpmOpfIArc/KvZCvi3c+j/qSjy4pMkAo34uFU27zr3zIXd+h18BeSoPsTw22a
wRCqIWZJnDjDDjFelqDtaVmx7iBYI18cucRRxXoIQ1uoyo7lYwBhn21W2rffz+LN+IU3O3rbYu29
HON+GWhu4QHDGhKCfd/wcq2FXr5JZ2kxlX3hReEz82u8XUnzGrLTKKcvOuyYJjhAhn7Rg3W/x4ab
KoIQIyVQ69aC8kDlzM+XzYVQd+TBchylRXAeaRMicEJcaQjn9SBewBsXoEvyYX7PbUFV0XT1udgh
FSG1sCSdQBtcPUd8H+RlEScBLJcRomNbpRkX1nF7vOx5jD4R+JgGWQaPFZFWnpZ2/Gya0KxUssZC
ks9+IBhWkWn6I7D5j/Hl+QUm+17zNJWw1xJTEquV1Fhxdkwt4KVieeo0tYXq0uDmM1gFLQMg5GWR
rdXH0dGtqQucicRJxIDN60SbX4vahdRJO04zLBpQ1Zcm3LZQyFuxEokHGHpkGyYvbeAC0/BQkOCc
iatunXULCcV7DKepyPNUYuiWa5oMEMCrozdPxgBXdYYDY/xpSuTcOO6l0g4ERbcuDGYZwF+CWGbO
GB9ncwn5MpMjQ63nyCJiHajLO+As7OYpxET2RTsSRssjtpQWcdvZ/74jhM4eq2JCMtua71VsLC1E
qjQdrk5z0xX2SXwoRpPzWmH5XXyo1GypMxDY9gsmVuqqJosh5hppDqmISb8Zvj7f3klb6UyE72+1
35gDP/Ezuyw5tbGKzf20hXH0bJcqkpqBssLtidv8nEFZIflZyH6fEX6PoRQQXbMgyJ7Yz4db/4yp
0D0rQbbtUoztJ/UxGTqzCo2IQMIp3l3zxUnDUmaTlkUlG+5QZ9gDvXhwDa2crQmuhsPKV3KdVYzk
gdxD+pV9rjHJ4aVFb974GHh0kyd6Yj2h0ySTBgX2ih+hTJR2af427CnmLOQXEwn13xGIhf0U4Hog
zHR7gi8GluZ+0LPSSUmNM3vHd0YP1I8Y8yjhgLAYLwlS76ddC3cSLRxq87lgrgyj0AG3vDh5irz3
6EpZR815k0YiKqitAkYfR8wv1hh06km/jPKNHIcFcw/K+lQzSeX8gQswbKzpqeviOwb4XYYHYCWP
jkRXVHqJBnn7OHH8gvz5QbCpnNRyjedbGgR82985VCNx9KsRNQib/ILkefzNUVg1j8rHQcjkl/Wy
VREKJU/q3WmYyOeQ0kCltctP3Quyvx6GT/SQfAl6ODxW5SdfnmekvxDzXfQJKpw2UNg4ZRd5yYrl
PCBgNiw/Mwy5mbMW+PvFdJE3d5QusWjmSIJMs2mIMx+te+5OosNUu+AC1LuGzozBciHDG+uSnj5a
wSKUYIGzg0eNzVLEYt2TSZs9UFSQIXJ2zV8ETCTuLhBeqRDCljq09r/4xsJ7Fz5IeOvigsonjtRR
yYNzOc312btJG4G57lieXJftNYomnF9yPupdBTAuuhEK5jpkaVX0hRE9GLv/M/PiMOv73DRGUeIS
LwNA0lk8wxwW0+BNuoqSAnsomiW3d5hiJLgDFP/V6WcMT7RmYYUpyitaL7JFofdK3YAieS+Kq9gn
bdkJBSZj05HfNR+HgMIIgWR5KzsFw/YreqW59QnUpqKFikGIoK6T4GoIozxAES3YCDbM3VA6nRqt
IgIZIQRzdKMgJtvf8Q/ngA06d6AzM9U4UkcfL5/OwrJBLQGRD2SAkZTF71eTrYBCMxHq2RvWOeG1
OoiUDJD7EjGqCUKYM22iUW3aXdWOj1N2/nxnDIwrOYCoxvyjncwJoH51XZ/D46S6M8dNtmcgrmfd
NTocT+8NpKSUz9UgcYeBZFLKjWQ+riy3g6P/lquQx7W2VqsMMSo+P9i73/0PQlVnPLznCAI4oDiP
FhRjb1jpEYhspiuHvM6ziAU44aK+JLL56Q+NIRKcIjYXNiMTQOE5JdLa7SHAPpDIXyCqMOXDLa3a
n/NMpbkTuRwl8sBBshbkuhCtpby9ixl7HMonDDBS6y4EUif0syK4LN2p+7wlbgbHBBiVYD8x2Cjr
kk+vFMFr00BLGQzy5pyl4Ovwmi/EjZllU4TBD3pmklT2bnq3Xz8rPnNQqRwksDsdOqIv1NhhxKXF
t71ExSfAaceSN2L+6vxPB7Ly/1qQRklL0eQrLyP1Ma7YLhgmPh8XhD+Hrp+osTU66SXObk2wh80M
x59leEtpZqk0Yk4dVzFjFs1auxJ4cotq+biDEHd34E5z1dXub/kY8rRpEOoxB3k2BoEDmxuETJMV
0CMYGP5lQuXnajtCXOZsohZLFJI7lEtWleGrXDMyK24l7aDCm200M/WkQKm+jPk7RVHfcIXnLWSO
wGAnTEd7i0Bb8oVgxYy5NpPm4YzM9V/YlKyctFIE15EHLz5LasON+lfXnIQPligaF4W8pSk7ZhUQ
6zzoZ5Zylte3Boo+gxEgeqfvppN2CwmhNav6AAOB986U60bR0nLcKWd382uXJ2Z1O/41mQyCg/lN
WvmeTymaUmNwH9h4aaiCvgKtIKNjHR0s6oogExZx+KzyCBEqHeqlD51DAPCgJnDLsG6d2Pue7pjl
HkmvU6VRVmzmLnd36MTIHHpQak3furxqPmz2twuRQsC7BYdcOEY6T67f2G0teSBjRv7k0YLqyQzP
bESfY1NxkrqXa8rv4uXzXFupLB/L4yDTVsLyhM4zGfo/gGfKge/PZEpjfe16LvF1dPkFpV595dSP
nkA0oJH3+ujGtLlzrbOTwstlsq+opojnw9iu3J3NMIHUZjA+lok9QSyIKCtr+0LXXyKXDZagFll9
439YeH9m39vZLczatZreJVkG+Qh+7sYJRv4JBKFU3+/ZnOXK66/Qz24ULFptJ9T4KKfn1+9dqXT3
885rVZNJs/GCpOU8gyb3iXXm9wLpQ6h7IBTo4tItDalDbH2DWJHgyz6+zrdgSrS+GmsbolhKqhKZ
YnU5CNrNEomOpHcC2s10czy3eKT8CDdZhJ7xaBfR/TlY+McpkQy0YJJ3PRkDnln7Ivj4hgOiQjig
R9Ugk9TyT0yCcwtnLgE017yMF/QE/SbIuN7z+pKEk2VaXJTxoKjCvv/FGP+s2ZsP+egMJ1cACBEB
GMHSxKB6VWVQFtqCPfGDLH6lXRlSHAZlmy1MBe4pn/7tkZwCnvR/ELA+vLBlAazEk2+M4PY2dE8f
TGt7Yx+hiA4FZox1Eg4rEs6qK8wnAtG1hW/KUVBTxdPuiU2SpfsWzZmsihCGEg3ZCRL+/oXfE8yS
6Ij4cnXX0nikbEDj3uyEJI80bEEr+rBymk9b1EmmqStMYsf/E3ATMrZckIqAoYmD/q3rf29hTaYf
trw7zY63Pwg9XL7f/52uq8wIxCm0eU39OcCqFtL41RfweNhCXg/fIrVRwMBPVnWT8wrPx1q7cfdr
fbxR3e1D4xNxer9zXKnisSG6GZTTwtdpaUmFAS9INAt3wZCnD0KN0YmnJ3lv8DryfHGV1sDcGZfG
dYj035B9m39R7BtsELjfHl7CV88Y7slnJ0A3pHpgpDZkKq1RMRigCY2FQ40hs/QHe/Qr/giArsvA
KeDWXxmrruKNCUf6Eoeqr+hI3o0abJ9tEZ9DQPE5xcTLxEvzrcIbBD2T6FZdC2hcJiL0hyxIe0Cp
d9QBQCiRzTNqFAOUQiYV00U4rZ34Nq+KzLQpqSyDp5JpNjbZkX5bDBkGnVuShW39dlkOHIvHdj60
WGmDl09KUoCpqMzftbDuCRVdClfcgqAzyyuplMrQnnIeG3+3UcpJkMFEDz7dZldX6O8a6Da48Smr
CzGnX+c5Jv/wuxRmcA0dZWVl1aSSH6m2lTsIgT6rrnQorTIWZ3WzzvFjFYJfLoOMGp+TeW7kZN0b
gehsMnES+4Ttc8tH3CsrdZIhvM7u+JMahPkYM/HD+Voh4AYeEe7qoKSBuMwGILGMVCq9PnhVicsp
W19avlb1K6DDL70/70YgwNyPlqWvfekdPXD/q3ZwYts2EdLtkD52D7aMP17U/q8pSUf3Ro9AnRdy
hy4hSGPn2bZIAjHnmnADToYSTGB1VdGZJ30SqNJ7KPcG0LXrRydLngIPgJZtNOEQh3AB3CfAtUvw
vLzidnBfwSKfz5W0OgiQhH/sfkYQ2DfcBOBj7mEec3FP6ZmdhLKfy2FvoWiBouo3KdXj3Hx730aD
yH1Xc/L3qhasFSYKYdNHLXMN15G1YVLP4e9jAESOwLQEOzn1fQn523rm545Su8laESXdrQdIAEMn
a/9jAd1EGJxx2/k1dRCS6rwAKhlWDnJKNEAQRt1RMTHStNlNYmmYhcu3mgnBZCYn2bZA+ByAeLpZ
fHfRWkOPb7tirqzwW8fbAWR6YKunIsRTnu8Gse/HLxS1gvvpWYIXENdooaESO7OIwxSBm6jtX9u6
lZKGtPrmY17/HO8/ZKcl7Fc0LHmz/MiZP4FqzLGEnYmErT8VhpGfGGQc/opcQhSKGAhzdvcDiMIn
xX9GS3tMDtLINChLT6fuBTJD1nVdEO8p78/1yhpEo2m2f50ToEOA2X9pw9vjpAPXfuErzR58SUlm
Dw9XYVUm8sfTRcKOOZkuFm7KtxiKKA9pNTPit2FPf+uJoI4Kjt6Fz3B/Jfq1P0pTGZ1QYYyIQZT6
+7KHo0mw9Y++0FZEM48K/ZCNhPAbr2P/tZH0h2C0sg7mCthyXjVpo+BSLJzZmJwDz43D92+nZ4w6
sKj1r2UdxspQLie7g08kvAjbUwFOZMtABb+8vatW6dFdI3Fc2vGLHXocRRwywh1xGlez3sB0dQxm
5z/um0uTOTbMbaYmQA9dRVDTGxg4ecD1XYbIIPWZVjYUbAsspavmwNHexhkgERxq8fILbOHie5T5
bTytPeNdzm73Rs9mehw5OJVXMe4nLx094+LguceluSzfnjOzse6Szvcb3DL6Q0+9VudYaXRc1CvX
0e+9nydFdUbhfqJV+b1IthzmN7wotr/Y2LNiCRCbEOHrbXbqO1fvmshOtJc9V+HJJqpMfyHvmG2U
QSmcm/vd2p182gPcsj9EIOtxw5tdtr+cD++ayMZgtW6TC8OQSAgPIAg8ZX1NPF6fXNtAvgbwIXv+
8DoP3Th9OSca6ldH2R5d8UoZ/TGsGEA4iptcB3jq8twC5nAMQP4F8JrWHhUDVMOsyghiOV0bbJ5L
3QRcTH5bvHaR+ZXUgDe2cZ8SJ3mlnjpsebfpww1ljphe99MD+mkc5d8+JuvsXJcsDZPvwD7zVFOu
RPFW+/jXfz8/qwx9ZWNbOROS1YJrbIfjHSR2QqopkPaGULxbcB28woKv+q5Vfh8o2vZ3B2Py/8wU
GyduVIwSIoBlqWnouGBj3P27vGmqcB5uVBuDHTxEvGV3btaLkiFx3jl/b+/qzMmrGhV0P/WJiabG
RnL3uOhcPYU6KOtJWj2gl4Pam5uEQNZxkAt/QkSyBX9U8xfnGuC+NC7qqALQ/aYga3Xk9f3XwYUG
Doh0vfRM3UHLBnAFBgXJbDyncVEFOFBN/K17kkRwEWVCyIgSQ1kdbl8zDBgO04JCoqHzxv9sfewQ
FS491LJja7FORJtzgkIDxinVBayEplN4gsoKQuW/Q4id02xeLf3kVAYloIlucaOBoqwNzJ8G4sQA
UIDqc+kk8La6KUe1YongJCUKOTOoCFROLChK4rNFnafhVChsMHp5Y5/mbEomo/7XV20Yroyb6jXs
igQeaLvKLtZtl2N61zg8dOnxITFL1nlfH98zm5+H2Ah/V7s0H5JGRvlKJxKtH1orMVlLqU0UsB3W
/6tRf0HoREwF7lAzPluDjobEEr5tjOV4lLh5ykFlB67XiLHgng6lEyeqS8/hG7OEe4lE10x4YBlc
hb8k4J5Qd/bkPV8RGzTj3VnqaJXEJXXy2XihqW75bs1ff88JX+qV6a4J3nVyegM7r87DmYQMNbfD
n5smzV9PCmri8DILGjMRnp/sU0c2Q+XidEbNginej4iwisMOf5n2rC1DMIaWXGbk179wWk61lENB
4mVTXh27S6E9QhoGkSSASzgXIHaviDz4b1OdNGu5P5HqK9XDm07dPprPoz4d1VhBVFlYlGdsY14G
blZDxsGy0kZmb2XRe+vXBtZD4Bzh2uwLmGeR3RzyGZuOI/Nx0CHvUmM3fG5mUufWLoxmWc+Pv3Fe
mZofGJBWbkku+usBBYvLUc1ayYTrpT8xhPhhIePRu+RRICiHeaIqfeymeTDdl24oUd4zkP++b6Ym
lzAH495vUY609YoCYD30RCWztVQsnCcxp/n52kzuSydtY6H3b0pU+cJGdE9atLkTnC2AmMAC3iZt
uyCjLgGhSrHqyD2TkY2715eIGl8bc1ISWoADzBtCZEbjprz2OJitvsJRer8DCm5iyZ4bucx8Z5MA
vmginl4dKuHfDpsNVrS5OgznciRFrwFi4nZZexoSzYcogzPGLgH7aeBQEJXQHHQnrN7YxrSZVCJW
BacUojnrPgS8jggC9Ajhuwb9F2ygnMLBO6O7rgHOTOQePguiSoYkB2yVMKBOJiFC/OSR+KwpAD6c
nqtYa0ZaR4Ekb5Pmbj40mdmcZT3oeDOGdzYkdzbiVEjdxR5IsPuICYYcIxYAuKWtNc/WMUwdZZSf
NlF4nC+nNc2ebyCXnYszkzfRiT2jsMB9RWLeHID7O2n9kfed0K34u7RfRWc+kW1sqzQIdsB1Ovfj
OXJwtU/9TTl5AFoXg0CZS1DGoWUq32tclMIOJkc/oUhHuG6yBiZmThMyRAfQSecaSsK0GyeLsBJW
Nmg+0B/QNpFLFddReKit06L6wJFDqm34UFgVIhUCuhhDS7ReReVXv2E5VHvyWgK4JaMKWuBkPi0w
ihwb1IhzCU8NC6sgvegiPvgGkRD96s5xokS2Dfhq2VYtv+Cvi0EPrq7f01xYyF+r4it+EYD9g1rj
/e+FPffeLWRaIxg7fDpBL33ml8fI+ZvVjSDBELiB/sLSc9mKxc4pMJhJymeAP3U1FFMBwcjV9cXy
lvIGvb2sOCRAciBo3ee7WUAc71zt9E1RVMryLSGzyHkUhR6XeTgfLIogTc3cl2+IWCAddVl2xQqq
ZIIKwGD+V6pe68HAwndbl2NidDWy0+DpdRYamcF0UMep48g7y8spr37bOUXy6BZ6u3wTazzCmHq1
y0l3nFy0092P7Et1ZtCPo3PxNWy+AzG5Sux622XkBXccygmsgOzz9yomrllmDl5VcQtAXIWiy1Kw
5s9AMpSOJacyyY576Y+1tcbR5Ac/F2cwZitGio4WR0O1fWn5T/rIsA+xnU/voHHh7v4B1vdoZmNX
aC6f+kLTSm8z1dm4R2YUfQ2EDLe/jjgeC2JhbdMQ9kRQR4UpWjgBUqSM9PPSmAgt4ipgCU06qNw8
oLHgZ8uAu4LV4V2AIQ8P7dg3FXzp+mGVX0opJSLe8Qd/bHgUfOuWISFUFwRxpLSGxeTPLrAKJubb
pbS5jsmm+EYsuccWGrHOLxgfSw/Ry0SxBQqjD71bDBhcNqcwkeO4dr9dL9n27ckTMOKOp1sym7Gm
YubOsvGQN6cU7mq88d03QSkniz+Gn88Sq9+e/M/833kTa6+uWe+awKWZ+S65trx3Wt2frkBunFzO
kRlWRq0B5jGzj52FnV5xrwXqiZ8gA8yaOdvTdF2OdVtE6FNwVR1gjSsQ/DWJXLeEzmba7IsInYS8
wO9U7VfJQmqM/paxAWG8o05z2Mb1f2Zmt2Wi1RRdtDQFXwpcGcVxt2RPQfX/yIANINyJxyHQdNWk
xyf+b6AmnFLZ83W8FjBr0RIAmaZZh11GuyXBdSVN+U3yTS09UujLZ0GRaY0mtCM/h76+YgiLftgt
FiKXqpYf1nsFHfc6tP3opDvef23CQ3v6xfwJheaVDCQh/Vixsbgwap+/xBhGNZQ4cN1WcEVnIOuP
ch2mu8/cfygFomHB2GSHF4abg4KJn6Z3HDGOa5xo4N9sqhUeNyi1Im07KiX5mn3E6+/GGRYuR5gR
FJvDM+iVRrPKdT8Xx3NuthpQDMVW69wmlyPuuDvWVkzxzXUJKLrwhUE/L3nVWCEnzTYl4ePXdC+Z
tuTksxBAdSlijxKCZTwXkOSPVDCLW6lPXeZ9EtSMOl9sgNlEAau6HsHwvvZC/QewMADbtZvVX1ld
TJ5WmJOf8dDPGRb7l9rjaiWRJ21fn3yR8JWPYqdXeW+iUHHDweEBmhO3af089xpnEpVcGn2eXMkE
8pbWgsIIY39dda0S1kVOA9MC2nmcJ3q403AArYIAkUMMvMvGk3X0RHtTf9RG63hUDA+nFOb0oYBk
bfazc01glug5gGga1995qMPNHnjqgGdsh1GZxEIgmrx4zqaAlzBMgunqrmDaW0Hvqx+EOjR30nR1
53D0n2iY5YH1Po0hfIKV8EJJGgrFz2/WoRRv9H9wnH2xG8VIIH89s2Kfhwzr8vtHEbVvW9/RThcu
ztvrvyNecgE6TQy203YZimNcMn3x5U0loVGTi95srpsYPD8C7dsKWdg2nDsgNYo4qCwjp7RkcYb5
MVtY6k9vKYThjyLTmMGJLEucObNfnEstKx83TcqFxiJ+Q7QTqzYJxNc6NDQieHMPlLXcxuk+w91R
KYInmfsYM0XY66/iBnEF67SYmY+PoGNGXe2enN3HR57qf8Bv3vInr7P1F2vpXMr/DXLOKxMy4cns
4tyHpe/CZ6WkbH2c74VWCIOzX9egABU3opwGikiv4SdpoO1QqgVrhlTYsl1mKmYc+ncqwrSUg/Qf
qXWrusY5UgNDPp0h5E+dsW8TlRcfYewoimvdfOjoL7SsEG69AwP40olYSTFJZBuXo9qpBLTfvAPH
0g+xmOek6zCXSG3to4yW2O2grRrl166UJ1jYMeAWYbx9e/CQpi/ubFereZYop23ZP3BoZoWIfbzS
axdU8HkYzG8T3FHyKSpw89L9Nc7PSIreSyXYUpijjG3SFv9DxYQ1kpo1yMkRz+sMhQbqH1bLIb0S
iQhEmJoaD7zhCIo7Rv4O6DQGldBoB0cAwUs/jFQAp8aGu7J1HceLy3d4pXJc74D9Zy2uJryRZUx/
O4zDj+CyC6m00z4Htzv7BYYyP2IGrBWgmVeL34OU+TDiLMqxQ7XSKsbu3UnVd32mfmthXWreBGqX
lTFV8GphpROciSyUd1MkdTu4zm+W1jMP7hon6JZTBkOUh+KmGXsbrlNyXaL5qaeIUHOVIAoxftDq
re6HIsshuwRpOYIZ7uhtiRZl6K6o3ezope8fZKIa4AGxm/QyaVfWQbkEDFR19d78quUH/0MK/sTm
Ll9aRqNiXgXW2/sxciu3ce9fc2BW1lC1q6V0TJrFbJ4jj++Kb3tGK3ptgFwppFSDjwdoJ3znz7fz
X0nGh5LCfjZNts3bjcNp5bKT29e8LYQdol6shoRDlWOYof6epZmqWaj9EpIZUP3Ej84IuC011QVW
BRz4mKn9Ok1KJvUIUXXIanFzVU/IXVnvDwg3BAaoJsBxP5Qy+c4rOOOHip4k3bJmv5oIt+QzXXLu
wd0H6HS11fOo1UE8AIRXYcwnZpRAuqzpNxM1RABBjeCb/olwiSeUfOcrlP+CnDqT4kiZz5GdJlU4
AF54eXVZevY6m2+3TcsPu6lbmHmRdgJ1OvH0GvO5I5GHgPfNTkRu8uzS+GGsLxP+HTJs+XECRO/G
1vynL1bjcyKRIjt2Xgy/JfDianoW8hBAlweNXqW0FlzSwTuyCALrGyM7U5RH+ATqKdEj5XyBbC7K
1pWe2TEuyvcgiL1oDXfm5EskS3VGFFXhd5kAHBGLF4vscYg/ljBDpUP/Mj0Fua5j74kyHBzhPxbc
j72rcTxWU87V3/N085PjADfdIVRyw0MdNBEGL68Ak5P8qH0lI7dtt61d25jqqhCkVzeQTXxDBw3+
bc3CymFSRst7FZUxBzpQmKeY8kSpnIQRK3K7ZyM1aIhE05zVyrzHX1mL1OLxfmngmYPrHuerDqFP
RUUDL9dhv2XWTKxY8PJYyWUG1pMz3mM1DPadAaS2W9XXnqSXEfeubf3weJseairx93qLHUFs8awv
NoKiM7onZKecc+LLToGeTzF7V8Jy/NYDnMmepP24v6sJ21UcffNgUrDVKErrMq9iLb/suelNqn/H
bYDQ/23TaReIPMF8s7mcFbS86P13ipHIzkz4417PTXQMQcpTbdkVjx36fogChgD6fhfeoovDphTs
MjCrtOf9ZEuaRxTcGY600OavSJFPzVkcJLNaTLEzOiHqXVAgEROD37mUvnhk58XWCxkQ1Z4czatM
wdDajOmniTLudQh10Go+tCmp9XioKaq7mZ1HlEhP8lkyoMW/FlyJB1flM3wRmvW3KCgYsvBLLlDb
BPIyEqUOPYDz6pBBk2YbGxZW9vjp4u7xJBA4JU9tZVA9y6Fwhk39MI1MoN+xisTSEzn7Ze+gl2dE
etalmUKRZzclcnCjA7UZ1DMkvkw+NrWhUXEPV1rS8sFQ6Gaxm6J3sjkACYc5Na1kkQ715+e2VOFO
9Jr3QAtUOCQecP3Nsd5dDjepQdTFaZH8efICpqP817f7gfvsRMMlRkSOQCchEUtlapRby7PYnlXH
GIs+ScVOR4It10WzpDRSBj5l6I0dEjzVqLJPGFsBbhl283VPvXc/aW1j9QEa1+iCunYPpSzdD52x
KIzySBe9LwtRMNMf75ZlmHCDRZNoUtu7ozvwfpkkX6AgmtogpKAIzeaJc15se3XE/3KKX/CYon6/
Vu8Zm3p8QJseho+eZBBN6LFjSVjVoEtvrdwCWt0hiPzYZ302zJ2sk8RKq5Z+49Bt3MJZvmlHGoCE
EZpB/hUpyYLbLNPHPylvaY8nXdoqz3NSINh4BLtNwjcnnfsa0U90EwZupvdGOUc1flVUu9JePOIq
UVKEb/vUDMj3p+m05TvwbnUzoWChkWRU4m5FP8bkNoHfhLrhse06015bxtCpgCLDjCvZJmjf9QFz
QoHnauN91AsFC5rTgdM2ATBEzsyRk3P6bLHhjUsIVraZ9wGXJNBjiHdfTSieh57Stna0KuCu0BhI
FuMs/k2/uN2Pch2vd73/nsWHl/1r6NiXAnq9oY2H76/+LkDt9O3EErkTSHZN/03I8/jMgtnysLdg
IIPMWPspLd6K3AibCuPWxlbxQIRHmgsXa+PmEaw9CLlfkeVpROaI+bbr2GXySNX0wKrxvANRup4D
/DUz/k+hgvtrbWM4VOohuJOF17URcY30bqNJvQ6Yts72qYKvveAIE2ehsa/F+AsYUr2bW17KkUYz
FdGoKJXeq9BBTF1VLimTXLusef+3GZa5z//pmJljbtt2x6ZyiiHWpG96ppl10KwIT+WXWHloONhY
/qYjZ01PYtLkjNvVMPeGOl4G+I7RC9XssnF5P6qFpfc6s70TINX0zo2b2wP580ORrbA6+oAUgP2j
2ekuaJO4x8Ta9Drb4Rgy+eKMJ5kYhjWSet3I/gdmF58jnKQ74LZ0ZeJUUp4NjZ1p7ZimVODd5DtS
Re/6c3Y/bA420yGm12UhOjxCSnAXtd0HvwLKZ8rBxGMKySFLvyQASg3JKQBl2OYLK20M7EzkQRCU
F/oLhUDCmKK1P+IIugjNZgTFFVGbURvj7yxzrGvMO30OyVPaHjrOSuXE4ilK9rxTPA1l5i4KygQg
en/trgWx0sw8E660+5Q0jV0cPKnIr6mJWhLtm3wP3ACsyt8Vm7/MZ4XOi3Kg4fkASJA5BNLic4UZ
SmEWU2jXJV/cXJm/gEByjxg2Jc+Uy9KLeGX7JZgL1rtkBazDCpW1cpBudTiPk8FfaUWBdLA=
`protect end_protected

