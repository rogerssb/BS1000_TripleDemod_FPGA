`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
k/BYGcITVzkj19j2HCuCh1wA+/VTFblj2MFzTMZNbTSHTj4w+cHpukw11MhMCn+1VpaV4XPk+KCT
F60iuGPAiw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E46yTwoXeRY46I4q0sknAG1i6oVD9Fby9HJTDGmhPLYly5mCC8LOLeoAWOb2MChDrPQjbs0lo0pV
f+CFyY+5CIt4nvyaK6ks4bOkktm8k4x8SdlR0YtaVdd64mBwZuzP2CDguB2f6VrE7ugyB9Pv/D+y
PzNO42OY0KKracv7T9s=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yaX0EGpfIrjKDq88PFxDkQ1Ih5gVPzjdX7cjvCAtwWOJixqSt4eknB4pThz4Sb76SURO4/kG72IJ
X4MEkZS7pR18pfDUs0oncDNZ/lhY8qySVVP5KvSvSGJvuEd4y4JWUPlS4pg+mBSQkD3ynhwRO+7t
/q5f+vhDl8ABSWnlKqs=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lea0NTFYyEg+GckCXsxSFBANfLYogm0qN5YvRb8u3w8ZQu4vVwMbl4/WN0QXKfZy2k3ZxNQKz7Dh
oFdjoeGsDLzMnKSnrBT1pHIi9PGOiLLrg6Lvgcg2TM5HrK3jIayh/Y5AnjoZLBttQ1q5cMiS8QeY
cX1MV+cTx4ovtKU+NIUTJbPutsdS59oWDtjR8DpN2LnfIJ6nXUntisb48CVYqNKGn3QZ5Q9SeW3b
xwlvAgIsUXzx0rXauLfH/BSPN91Ja9JgI+cb4+D8D9y/xpsjpMIE8qGKkKZT9w3gDP0xfprRY/mz
eayiSfKIPy4P1XQfBdDuTHG6udNxb3Gn/xvQ7w==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BRgljJEeP6z6vVvDwBuXh9cKW6awpue+BLUABGrJ/7mchmbRYCpvdol/LFGVHX7yiQwqBDAClMv5
xJ8KbMro6CvlKPYH3A6NBuEbPnBfCSjWwn6p89wdQeA3stqsOw19i2oiIX9DAX1HNpBtiJCNKdOK
0nLwya3/SE2z1/VR2GIcR+tak40u+wRkQbZKx6m0GiWFvcZRKPbiTLTFnTT+MDqgRgoAjaUHaAVw
tP3miNiSXswdta959DVvVuH/uQeXipnpEKpytKyq9/QSzS8wsRDdWG0SzDLLITnXMD7C3/ZfGirJ
+MwqxM9f/pD0A3k7376qqv6kz6YBPfyVcNMy9A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t96cw5VHs31F0QSbsQRgm/N4gTp03rujgsz0kvvkpIXlRIuQQZQ2TMZI+9F0Kqm9UYCsHzsucT1R
e9dnnzUZ1azv6XAhIozJmAJx9JNqEKctF0ycLby0+bxLRoIts8dWX+wrK8RjAivYtKbYVfImpn6A
04qoiobCCJh9Yq2eE1Mw5yELVbAtnkGGTfEezmcsny4L1DIRf4A1ISPYemouvYdZ0B5OrtXZDX4/
+6fMrKMr0hHxqHGqmi6lHskRbI7/T78PFj6oG5Hoaw1F78As5mttBqvaoC5ux5GCrNuIkguMTWNE
sRdfJrMxL0sNJdDNsC2po3KppjTuemj+5sPkTg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
ILJdftLFavjgyYP1mskNQsIEXBtHOewS5a7Eqq/o9Jdky3Uytm74PysUtD3A2jsCmGhfJq7B35mi
pGCKTjCgd9a2pPDdxmRou6ZP6zRgOeBNbHx+CbcDzq7/oQsOcpW12VfcAMH6EBaLcrhk3Kv335Sq
BJ5iW3GBmCHFJ9ioDv0eIoJqLZ0YYW8F9LIX6fpgbOPgZkwzi50R5p0X6XjPFRFH40Nsc35TGJal
4Xg30O+oqCh5RQwdi83mOoH0zhAIJNFhTvnzCNTkDxvdFkWJLwg1aFP7K89cr3wKP2V83hwTFDDP
vANow49fbn70OA+He+CKoe13jLvcBFW89KmelL43cmmNOa8I9gvi3c7tzQLGccrqvw7HNhRjqZIg
/NH6MH3xQDh3Cj/CP5VbsdS0DKGXpFdjvfP3JEi6hnckoo9/NxDio7yM+/yLDRgFYLnvjYPf+pIb
BMU2VFZsnidd6rbBzoVGJS+SEXqQO2pnrrKo/ocjX1dtFEUmsP0y0YmXtKeyh1I05g6ds0yHh3Sp
pUpT+AvkXGE1G/tC1+P+ygNPbKc5AKRsmoxscZxeOml0xB0e7ZpwGnsi3aKvQ1Ma8q2SGajhTywq
ulK4KbCLqY0pxnUUIKn9vJRjVnnGz0aCv+WPQydVKOvlcff4eyf+yjNkRrc8Un2DBWrBv6A0moon
ypry8baWVBTC9II6qvbz+kw8XeVa/rD/dhR4p2rbOJ/cK1UYJZ3Ymy1UnUW6+GUuBeCJ9hGCeW/h
pxj6dJx3ODuiVRBpK761PSx04rKOniR22PgYWciGXlNx5FZJuki+z7PSc5hvmBvIqEjnV7BX1a1i
CnNEQxDnizqyDwC61x8oiNs60fozQvJZrRjG47Kec+iea9bd0vrDpnJIoJSt7vOdZgN+VSjlRpTT
4uT5g7rzPSOiPFKpZjhML/GtMJRBVDm91erAesgzflE9MvjFWLaVWGv08qQK3jIbYaAhHx58TysY
hs7OddP4Txoq9L0EU3o8vZrbVTtd4pWHbTcguAb1oj8IaShEmNyIjQqYGUBoxZ2akY7b3Vg2Dto2
qzuzOnwLbWgbZ31fAvETe9BW1xQmtuj3rPZTI1dpfny4agcoSaL4GKosNhTa46n3CHUl73xcGTUT
4OlXHTFqbSuwMEUzLjeojK2r+5DqFTQXm65nMcksgB5unNfkJqyxGut9sz/XDlJ/9YpgUD1xOmRS
Bgd9Vwhb2WWGTRlUEzU35mk22E9g9GEkwwP2a8arX+f4cJmCggOuNYX4oqTfw7NBNExMur7/6kDO
tt7c/LlBaf2N+UjUwItYkRw/+KooWI1M6VKOD1bF29yAmYuM7Zj8lXdNSSFAalJQqH5D1vXsIMJQ
bp/bZI+TkJSMlLLPublRjiRt42zshGUdx9rdFi7OemhE1X99giOEzWzZDC8xkKTYKeYBASL5uLr3
irh0hukhs84ekcxMEjbbOLRQvsXkSfkHp9UkeNpenSnGPoPtK+80ZemyZRarPi5xisGQKyDXdla5
SjgLzUWIRSjwB+S2dYq6vLXb3LL2iINuA2EiNk+WdSaRlX6ByFpZNvuu2mIlsd7Duwd150+gtUy6
5Kkv1l9fCbUl/I4qG0jIpG+flWUBAGBuuq7W6F3cFo13G1nGQBG9EKiM7B+J42C+zy7g1YQ92Z6/
e233q4J1sPly1YPCCTR7R1Sokk/GnyZ3qnYOhGC9YmDkVr5j2zl0kn93PTvbvYuKJuvwpUh71pZn
Cdr/NrdZlTU/CnuWHLA8hV3UhW4kEFc/rQlE3M26JQL6Pn0fDUA84NyBTuHqFWLQM/HUfyw/+p+g
iINL5XwHaXytCH8SCuE5czCoL3xcC68ST56RlbMaKdH5gpIdmAS2gpyIJ7tXFHXqP/AQukhrgTVN
mELl6G+g1PfFboWJV/WZm3FoZlJej/ONXcmnBsWp6FnVbz9vSBPtwBjuaFKQTpkCpVhoi3zNI0VK
Zu4OWQ2zZiF5bAlh14c1Th7mRaLHdanGiKvoo+FRIszOkDzPxg0y9cJ/JKuGbZpfBcsytrvox+Nz
K+z0FLPNDFH92sSVPB9QxTp+NQu8NKVX2Ez1zdenOtYxOPe4cbqSL/sRF7QG+xxhmk4jOeO0qjpP
E6BiqVIpBpwTj2Pyqi4uS1SG7Ht4TC9MHDe4krTTH8mA6rFFaFP3hNHipaTgPZLMLliavtdui+yK
EGBjoQqc1lfJKeHJTsGgCd47teHiiPemEPLMZDzKIwEpJNxHcoiMiMP9BqK5iuK1/wjqxjHi4vRv
K46RVSp2EbSbC0EwyAifz9F++kIuUIpdLjNb/86prSStmJkDiBSbinoAv//nwqZCt9c32Knnhers
oSWr3zul+nT9UfrVp2G8p34sMZOmte8SBHRhVRWsuv+aiGLxaVVxM1eu9WL375l4pxZOJuhYr3fI
YBMVf2ljtcipkOQXkBmoscahSu4/AWe+B79e339z67MEeAqvAhUid0rNQtbtPzRDe3/vLv95gj2p
b27hmvcMPn6jyHfaRa3Cb8NE8HSPtdpFStKMa9wd9zgTgtPxJVqHdokEdXkRgscxeD+OzKenJEMV
gRBoKNxWB7+RnYOnbV7hf93ngK23S4CSw5JX2sE3FwS0UM4MVXqEdeJG0/7LGu9BOa8lyGwJiNDZ
1MVDV/RuWnL6F/V2M62E6z99cW+acCgu5LN4yRDCaYCWKY2lnVSnQCWAPfxWahhGpvAdeR0pNgtz
PlqW9U5yRrSEmTkSLqN9Sj2crfkb+LgUGSEH6v6LW3MwTxj4aUUCXE95aig17iES6XV1bKVmLAtG
/Br2ECMgw7goYS5/90xmV6Dom2NUCSOWKrMkBpYsuFw/x/HIsl2gC4pDvkv45nyfwdS2YKoOpUAp
twa6Cbpc6UH23xYI4nZZ7OSfPGPB7G5+u1ODe+TYJJrUFgGSo4CW5NjpBS0VBF4etZG5bekKBkfC
Z2jNKAv6RkefaS0alciMB0gcbiRJyvWDE5+I7z2+eJ9+kVyoFhjN0J8p5pQwdNLYI8oDm44E0pF9
7awLwkPKfxxPtpJ+HQNnVVXyziUPj8Jyn4aW8wpeMnXtMS9j7KgWvf6MKRTnwvuWqzPP6kzn1plf
o5RMyzqMjuZImXb+N4f9v+3XXo1U5uyYtn11oZ8Jy0HZE18Ge7/sA/5mjcj+TOzWF7tjbx45nVj4
+AlqPQFVkf/Vwd2N+Bzba8nOncqPwJEe80yBzsBATiYntagUIZIsYf+0hKIXWx1oSyUC4rAeFDJb
kwfM9Y8W5kynHqqwrOOnuFPiEoyDGIGRkgM4ykfTR8UxTcEztXanOX8/Bs+TP12it8LA8a7RSvWl
Ap8yfuL3Vbc0dCAGDUe0SjCbtrRBr3sjbVm/3sG2IePJ8tEXYk5HipsjyyAFz+3nhSp6TMGyHwct
FdZ9WWuaVdmcNA0G3HlGCJHu9YEeYrBIpEUt4QiTyz0/JcOZCNTg8N2+mSU3HrPpQJH23OZd4t+B
dJAv4qiFqoQoEnnen5Pfud1eXsY4ZLYIrcV/EiV22DGdBOCjbW/8/aKepG3g7ILqZ/ulwj02o++j
hGvAJ4pNS3YEixVSXFb2/1HW8oHLxtjxd2andVBSxAIBAQLE/1csAApHqWU0RqANnzlnYv8rV26g
7/q2G6W2SJOqYwzHCidIlbappqMx+TQH1Q+JD+G/aoUuPLtifReZzZwCX5UjjVFhCOtiXtLadjwE
L0Lf4tIYqgx2xECB01YejZZfT1lj1j9JipAclf0qTnGgGZmiHKqpLpWkSAQ1566ISzlaM/ChGXxr
kqw4XUT6QwKnmYIYUeTvTvrzNVlllRSPbNlYg/CY3CvyQQciE0beJ2Ahu2lMpbihTuVVPL5mThQK
sQj/zbHRrf57GZlyUICc+XsNkwYxvZFXO/hChIar+/c4uxkh/OJqirr44yPDyu1dUG3fboxKgsT7
KhGf8JU68HFp3cU4073DAAkBz5x2rHeYKM1/XugC+u8rufsp9fb696LwEqsKsxF46Fz88vBEDfRs
I8X+zvwe0MtyFXiyYrzixUibo33ggmmMalZkn4iUKt4QoYS+5GKSDeJNjNqbjGXYVhbcHsw57jk6
D2AomBlRJhFFxooO+QB2KSBbtR3V3ya58tXZowegvdZMCbO+8ExI3FF1PBReB3qa8+r8A6DewFSP
HvYYgYQfLynRi2UGPdlf6i6C3GMeHPet4mfKTxRLye/Mevv2ODlotg5YDJhRgeBc6sJFnOUbWuvS
icb/cvWt1GDLsxN5XaHM9oEdxaogRHlmtkwhLLv3HX+zb0Q5p2NSfDJKv6AywQ3joUJ2usDu1Krl
SDTigllPajixb+lYhfmSubJJfOv6c5vZeO4hIQWZDRFy6m6JWt7ibG63k7tHvgzxNFkhQLd0YReq
00Pz8m/8YyQ6VTqBV+VAsCdbL7lJIR7NFNhxl6FHF+BF9JS2YYCWrVXmT/tAQim87r/soEy+rCc3
m6ASqASWeL0V4lP6fP1vXFgAhHduwJkmViQyG7UMnjEhsa8mUhYq1cbKvWuCjMe4ZbFu/TeoBcUd
vAg26GATWUkHLk1Kc2hSZ/rXJ/0WbekcJaiMOYdLA6puIxr4JR4ww8l9LEiOj6d+BEEplYGJKqyj
MV6nPbm+JSQqYN5U1woyNsVSSECeHhb+HOCLTNSACGy1wXnoX2lmSNw+KLvWSKMtsrzLoHVBf2ow
9Za05gT91CIXVXI3vJIw+pAttNeAgW4TfFCMc1R4mI+A9hQBhg1aRxqx23qtP9RWB28iA8dOgn8p
CpccMgHBkPRs99hYJ/s6YKXh/kWZIL721aD5ovNh/Z27fkT4q8w/3acS4AHCoGw7RURVF3G0plie
EFCCqMxVdk7Cn7IeLSO0NWeQV30sNUOybSiZAjNJkg1+/qp061KtOLuG8UNKlW/2EkfWz9pkdhCg
a6Wy8E8L3M2Ur+l+ESeXD6fII9l96mmFeEwq0gEaSoNHK6OxZ3VFp/kA3fdL1mTm/en7ouoKeow0
SGF1+gnrMxPKjKDc5s101aexNaUCVDoJsQ+nRmFy8cQXiukIBuXl2e+a5GNb0v+fkCiUFAB5fCTI
tHwIgZ/d0ctOZI8oz56v9PtQ76F83ZTHwwUqCNZT7s33o0UNJGMkmM7HqXBxC7F4IWw1Br54FI0e
zGOaj7AMJxjYuveMWlYiHUj54s84bRXOGxEgkuFKKdGwFW3uU+hyjN8RglmE0ACVTWgORhXiFAXz
W3bolLgKSMZ8INKAnV/5rspuPzDxeJVNTx50I/h5tTS9e2KAxgEJ1BV6HLUDMxjuWJovn/lXfNt0
PMqXjIc644e8E8Gu3M158UahP+RESEqpSwbj7NtAENiwa9brCt6PSAefO5Ofe5/CusxAtvUxzbP9
01gUp4vkhAfYlf8ZIprbvtrugO7ADTLAEMA5zub8/AGbmJ3Ok0AYY6gc5xtozrG7uon9K36tJZ4U
h0zUnjyLcyqHxL/+DRzTkd8XWZ6xVDiXPLsHT/NEECukdjtfjQfr2QFc0DAtV2FGaSb2OEPdfLaa
ZIEFtoCAPwruX+yAxbkMcLfUllJtY9t8eqt7Zzh6EMlIWLL2QTVbwGu4hXRADBSJvHWKkNOPZfpB
+2L29l6if+/UlFTJBFo00gyq/d+9x5YDGmD2WsaSb/r5uxQP2wEzqAp/VIdxZlhYbkoj3tBZ1sc7
TLZ2v8W+s3LXkDhvR/APm5ZzeYDWiHTkBAfWM0hrkPYkuSgdAldhDmNLcXjet1vkzaU0kxy32rvW
EVm2LDTPfg4bg9q6pPxCxSW0BZtypmmDbsI6WBfTjgs4Bl2G7e9T3n3KjY7uxsERnEsMTSe2u0Ls
YprabxefLCRX+Oq0Tk/nz7cRL3F8nsajO2NHzTZem4kb28MK0bIaNdE4tihludzNrRYmoWDg7GWg
jdBSY+VmOSzGqZHfro/8yzKLzpJSdT0YV75ZPJzvnwlFipmf+PLD5JEwXdTKQipuEvkhg/S9t/zP
u2Nw2h3p4EyDm4kf9yqYihky3BzwoMtvapsKTNdEOXW8+9P4ad4kQh2970bWAfmbp6bRJbayW4uS
IQ9tPiy7p6eW5tNt6mKtG2nejdqq/YR3gFj11cm3IGunQKTt1hhwUI9R17oDMFEbvxQ+Yf+22f/2
fHcq5YI+1flz6aRdgUjaCAw1K76rjUQw7rCMIO2mb4oK8UTUhzuvj/yKIk6lb6k2qU/OSn9523PF
bcfIos5tJQ9Te/UrZ6j/AGV3IPZga60adcXjyzF9BADulnwEgBZMZoy2vtfNcLwyNrjQ9KPLx8bj
ERLP0wUf4bvaapzr3GxroaIHMCV6sNnSZ1/SzSUD5fdVTQEdg9KbKwUEUxi5gTB4L3MCVp6JaUXP
ZhMrJnu4lPsoLM0aPMjDbApREZzdSfPSmaj3+olp0rxjbhNol7C5hQnQJCWJCHhKRUgtqIvQ1NqY
32bDbz9aZaQR2zZGtUYSsFQXHkIMKfUDe94q/tV6YGoZdsFVaHEjNXzBVExZExWGoccgaRcODBDW
VHQ9VSuvNE5ZEzdUtPtyGj+Cx1KbSYBdHOF2QFInAW4Q88qSlwYBbLsEvJAGiIQMInjmQpyzV4tK
tQZdGhsoMmQAWUBE3t/lwI2NsrGMdSehryVATqeBq4YwT0KyG+iYlH4ABsTs2nCbsTXUDeZKnqBp
Yqz0tGHUNzWFZTnRwXyRzSz5LdAeCBdrqYSOZRNMkeli6ACFQkSHl1mB/aZGSF25rd9EIwxvnajK
3NrhEk8eQEVLfBN4Ip4kiy4mlk6kePmG50wgSj/g/w5hP+L64n8gn/BKZqsfgSlb13EsDDJlr9wP
Y8l9Ijap8GM6Z8/p080TWTVzVMXMd9AxW8ZIvSgK5GPnqKooz9UVaB1c1bL4/2nha+aCE++C0mz/
6oLa4hCCqlxZqTIuzQuxOPPyDvBPeSqWiduFiMUHQuOHKQYJbIpRE4ew6A1ZUAjBBf3dIuubn35E
aNdh/p2RTYSTCkAch5sN38RPWknAUmWX89azttBOxkTfmRF7baW+iFSqvx/Cn9uIxe2SC8WPI4s5
xLWrSaE1cxzXU6Lo+DpX0FV3xyIykrB3g7Gx8FAZAIqwcfqrl3oIOkBQtfvYkaY+G2l6i4PNh48W
8Co5oDr5ps4IQqFatc4oR0aDLSiwSgoGZges8MO97cFIXZA0CVHyOo72CYVdZHRfG8w/9PNhTsgH
n1vCmfabCHsaBMl2xdN7T3eUljkMI9/BIpEY3Cl3d2mFz8H2Fhp1JNON4y3g/Nei1C/KE/2e/mvQ
FjXwr8kYiZhQ3EWZqExYJYabcCFpbYOpLCrxKnKYL09Xcuzmf1JLepyWuj8Zr4cQzANjATyJgBW0
2XDSa0lphd9c/q2ceu/r7/otcRXVX8MMt3ANNPDcUIrDw72GMccUlbm1oPK2H5QRDumP+vXR/O1i
k8AtSCwijP5HUYIOKEDRhmW3+dmZucksrkBR2QhFRIfgAEHRlKm6Ic9Ahstkca9eQm5bv3Mx/fUM
A/YLj9P2z5YnHBfmRZkCo4OiMDCoMdaEIdquugkVDt/Os5AQB0eHxUaW181xTMlNMFodPLrsuqn1
J1igXE3Wv9c4INnG93HGncX30Vud1zw9Dcxl2vGjiW8hHQwH/nUw5pGJQAQydhFqZZN6/Ifpcq9v
jhyUZNPL7g9XISxAry0Y+rxtI63BwmrR9O3nw0fhvBt6pDKU0k3jW9vDrT96XpVYwzlQ48TAt7AU
Ko9AeOM9Tgy6ytW+00Fbhjl50yx393QOMlNEiCACAMEq7JpheacgdFkcURoeEVCAipVVEiiQcEyk
LOTSbqdjeJgzZ5s028SXwRHo3NFeKAuTbpKZGoZpVbS0q+p82iVlJMS9W4rkpYRv1AGYJDXhfTiF
5Rz6ap8NpLhxCQ6ZiBBZjVyfwhd+OvakarBGEjB1fdte1aVeCef5ChA5jZwkL9NQiMjqoAaLnszu
3PMALlBpAY5y7aIKyCKbRAK80jM2FWkccBWJkMDm+ZaKFZz0qOche6KZkUnZRBssI4guK81siCfL
CdfHO75TXJUpqr2s2vedKCCC37FqSepR6/aqdwRpvQ8N+xiuEUhUvB50A695sQ7psbT6sWtLsMU6
J6xqA4lmb5AKmjDUCilU+pK20CGp7coIOvMbTICXmwBKt5WQmJ6lPrG6PLDAcH8rpi4fr2nHoUCG
Sq7Epe3Pl9pUOGKB1iytSxoFpHre9D0x/Q3WQMh8sJJ1g9b6r2UtDU6i/l0g63nFJ1Y2PJ9QrQSK
JDGTPV8i7ZHgzGVz7TxD93qKORFKw2GBCdFHWdOaGAG2WgpXoCTv9+eYVnmU8AK0HIZbE4P99mtO
Q+4WBs0Vt+Ry3Thf0KVmTzpdn4Y1JvHU1/yCFljTiyMDHhUhrjZe/cS02Dng+KUM0Nv2Xqh8QlsX
kRzj7dkrJnXVMUGinvRYIZjmNetHCrN/XHPAdX5zpZcO1Juu1W6LXrsZ3jAERBKErT/cSKMyIcDC
TDZN0fqm3CSW2a7sh8BYcLqOa4D2odT1utn2OgRwMoeY5Cev3xWqaZUVZ1lJ1iTR5h2zDAAkQGx5
lCMWyTXxqMiPaOl3Kp2de3xyNPtbBd3CTdD5OE7xaUiWpZNiBdhfVqLcuXFb1jRpML/W0SGkGL5z
ISrd1orDJWW5nBm7osqSwW7w2DP+smrdBcZB9CgoRJhekvFHpZzzC9X5NVOJz/NoKWWW1bzggNH7
SOPua+NetB+SFaPqkP3taU9yyquPWEiBRVhEIO1zPPC+6OaLgW7MmqRbJL+KZbGUoGUYjREdX/oE
44FwZqejURXzoy5EiAmsUi+it4S7Q9cscLI/+gt67Q34V8wXqpbdu8zr2PYkJNpC7zTE4XEEYgRR
yw3kg0aQYuAJGxJtpoQC722BqBLUsmb7CU3RPOjRzPrEIGqxc3grzreVkYpR8Z10H7BFjQEQnrui
eYRw+l/8YgHyj94p+LjJCPv5gfKQelWK78R7WTgSfioq5ez08LV6Hi4eoa60rJcK/hg8ESOJZVWe
cXsHVJ4RPt/9ybconM9opOFlXm0e+OPrRYRoZ/qbqDRPPPCHp4/F94A9uUNAa/RN1/dYDWja3gLm
vnT5/jC2ENy6pa1+Y3O/7LyFkOiyOkZgalEmpbn17klC1Pk3DAtIaXJw08hyeNK9D+HgSdt1O/fH
JG/LZK5mT1TCFYBCz48lliL1PCyy+M2kd3bL+u6K4FGRLD13IrZwSOwslGwSTBFN7aTfBiKn3/8e
AlLtMLd9haTZF9FnvsCw4xd4rnpa5chby/v4IGvwCjvIzUkSyVPGOptXKp759c6JdVN9GRzVFcP3
8odkCOYOQ8WGL2IMNYwumwDP+orejSoZzoz1ZvjES7bB/HoXC8dqW7H/h0+TGLq5E+40AjvRGvdT
2PUd6fAtYSPTfdyJpdpV2TvS/A03TX38onvqsIqeeLk27+KgGHPg0PXjyJ4KGMq5FPSdlDZCYvzB
n4DBlRBzYhShT/nraX//JwgWXR4JyaMcmjvGCoAoJ82KOgemHCs13wu45lJUfdeWx5mJx7Mj8ruR
VYcpi4ZMcjEvcq2lJuxOiQkzIiU4rZUlpCEnvB0u8nieaEk1C4W1PLQGPalyf90nQhSlg3fzoSql
U2+IJPQv2afQ8RYJsoYFOYiqk6TJCZ8eQXq9K7ecoEGtZS4YJr9iIedEyZwC25qMCgTvQ+/990Bi
CUdeX7vcj2LZqG+uPQsK9PX4os4Cy7OFTleoBn+PhcZ6H7yPBIQsj8n95D8tAAZT7tKBFApCVMQh
+MOvZfdryWR6I/pfrOrTPrUK5uUeXITRzftR6vsAKrd+1n/TcFJnyx74tOX+Wz0EPAo8j0S2XL3N
rzSHhFSdDCF3eCRNaJUCaTolJWXNWkALc20RvPJGB3rYaJYYQac2bbDheCYp6gTWXqUzeaDx5MxP
2+D5FmiVFf11oDAszZ2j8o5nkQUh+jRucCw6BO7uwFJH2hCXvaRsrDw3/WQ/zDO6u3Ra8Edukwqn
Q6WK7ynjeWTgJykC04y5t7B+t2EJG0/LAzyXdyBK0oaIZrdUVcz7eSjilVWbnrI57YWOefQObYFF
Ior5zOMcr2dAeZ+K4AeHZyNgHchcq8Px8umcAZZYzDy7mRtE1AieW0OnN8b93PwidJ9OzyLOHybx
/wCiPQUiYPRH7D0vCAvQ3Eya6z+WxKSEU85dne49XbzBl2QjK0tB08NoLxBbkKUMsUNKA6fTRnQS
GDMQrZNSZbeQ/BbGJxlUDn57fWwlTTwjdvm2hIF+WO30C+kK8BpvQxK2XP+8+m8G71ZgTtG52uGv
WnmB9+ZkQeDjTLEMcjTbBpjeb8E/rprFZvCZ0hiOX1tOPDg2MATUmyfBn3XcLk0p3gEmy7jREUzK
m/QRl25tWgmQZS1kDq/HJaWJT37DesZiM9GmA7kU7TUS1bQUiIkyOLJu8tvIOAe6X+uf6h2hZ6ak
QqzHxLnDBM9WZ3L2cgnxzVgmyXEaLIp4RcJXvCyE3Vc8ynlLamx4AAlbGf8tBs6yw889W9e9bEEy
NNAXVfSa7HxrY5HBdPGaOSmlVmR6sD58Egz2ONKnVnxoE3DF78oeXUyWGeFCP5h1JC1pQAe0uGs3
JYcCoiPA8g44mK87eRzg6Bvg1SnAnD84zrZdIoQbhzVELAa9uLg+r+Pmg/H95U9uzIvzj9K7Ycxf
uNggpFJLKlVdG/KKUMBmsXS2I2gFfliKeBIxDQxvD46Yni7rBzrbXZfCbhN9MP1jrQAIqQgTfS3G
gzB4wwGCiYG6r7e/Bg9pS8jGYfOr4yGYKUTbRGD9CqLLECYQCh0W9pYSDepbbv/cI9BSWjpZaQdg
J37v21EX5PNBc+Ekx2JTZ6u58irXmmE2TU/cidZyEbiAhjZEeqzuA26xsFvcOAOvOnp079mrwmVI
wGwc20BYqSfetCoI8AR2rStpAM6XaT5QRXL9J7MqlGp/IK4CopvSjmriShCigiHuJc2IV5L6J5At
pYH2Xs/GdqNjU8GH70nVjtvI8t3KmvYEcSgdQhIp4bscFYCHDGoMEnk0QmvQMRfZlaDNWzJqLFAG
oK/mXedUeKnQLJm2JW3CTi6jwOYc8zr52ngyQHCgrMwtqbaePmGoGg5l/SBgFvxUEHR26Vh0OVpK
Qt+FSXXXrUPlAuAmYtLfdVYQIxyYLIRzJR3PPsEhuCL7zrGsL94E8QD1JAJVp97kfGvlicRg6uqy
BNhwJjPJaRUlJCrU/XzX03DHMSv9Onz+jBnq3qbuRDEFZqrEBvz/hcF7x4LVuvrYIvyQmq2Yl02f
nRfP8rZl2YEpqNqDP8Z7Dnmyj4i0+zcrbYE57Zff7WqdKow/3jWxk82qXWCNc8fZIE3NOFNk5G8R
XWGnz6QCwZD8KpxWAmqbw0RsPz9TD+9BKJ4LatH/J2N5aoIQKnlk+h4TgFFZfolvB2ZdImxQVL+N
/eR4xMgH0Ff7078+NVeCZntupYXkbk6U2iToCKPMu3YsFIod7oC5LbtBMm8Ha6P1LO1DfXDud3/p
1jtHzakh1LmRPEBfJ90PEUTCNBNq8Qp5CqBW+eea3vsspOP0MK5dnVdtHYFS/Ie9gykIENi3UZDM
xRCmX2mSYJ9fV9y/HP08D0eNHCNuEYqQNTl4GSlsr9ccDpPxyYuODXvKo13lvKFJ86SqYhdYCDLh
WCg976q1DObY7Vjz55RFfdKbuqyE2Si8eWgDa7egJ/VTretMuTJUF2vwf5BKsI6/8YJBUzGf7wqX
ssrGabbXFW7nDFw0GlNn8ejU/s44+lXVP34vTIUdQ2T41eNMLUSoXbfDAqF10u765cyUQ50yqvYs
0F2QOQ7lmbx+0D4pp/eDzH06DT5Y1kH3fSI68vZaUVokVhGGiDd6Pk8JWe1w73dHH7dK4BFDXDFr
cPsEfIE1n+e1dbBTJVFMkYKlIKtwbd+16QX34FtEbv5bip/jctaxUQElWwNVpY9Z5+VrJz7SOEKg
DzLYgqTO6IKWMN4VCd7EmdU2Kd+L5avjkeSBrAmp6PAi7wYcPjnj3FFP0kHQ7GaqOHtul2tbjDmZ
uhff2OPy6T2Jz/xPZexMi1u82wv8oD6ilasQ5b6fC8A3oEbmuIP4F6nk6piEMtdg30tNOXZYefnY
/ycB9Jx43C+U/YqSkF0DtFUsXeydhcua/sAgT6hxDjEAk0kzm1sv7e87A8J1E2GaYNtVU1xxMyTN
YKEQzKA61XnT9JWGGz9i2iXk6gEe4dUc3r67txXqwv3dh8axyN4p1D6z6KIbXI1xe77JPKPk2DrN
P7OVjUI3COGR5FGUMYpzI28kQS0/pW9F0xW9OG1g8jrpDGckV5qrqYyuMYlE/zp+cHZgYN1xZHuS
C3WNPPGzOtR4Pz5lrb4zvUgMY9o1TMScCJpcqS82NKBdLGU1thXPvaFpKx5IyP0GxDW3Ne8mnSdL
W9mWQSJdMKm1DCebRhiKrkiAgGON3pVx6A4Qi842mekJb4sEEtHmZDTPrjO8Fa6KeWyuKcdVH1JN
I5mvF7iV6iAC4xQPQSLSgKIciKKfHyfd1z3GnB27qovg6CIGZ/1WTO5a7P7s5xfRTQACuIXKqO5Y
kTiDZ3byR8o3JWYoESH+EPHc+FaRklY4NLNqF7MMBdu0Yxupx/CO8009T+9gWGHtcRPlisxm7XRv
AROxcj3SY/I4kVZwNLYSsSlt625AKJJFeKJ4TLfTMLHoLqIo/ygfREwdNYiDde+GsgLz3711Fpyk
eVLiiSoLYregnm/9ILinDcBR6tNEIOs1k5JXFKY0FDZxuSQarLSxOqM8Fd1wehzhbNzM7KdTLHhR
kjrhUfFT8irKOXaO0lk0B/pkounydEK+2CoPcBke4tF5fbVqH01f1jbKZq8JcAbdbeB/ylBkqJmm
J+/aVmiqOIN+f9rs7xZDKaZ+hcKC/Vpnx7n2fufMV35Jg00z5bDUTbS9gKWuxKsjNXkG3rld7k7e
ztnBf0lNECfu7vLecs1HU6Gq6GRI5fvEM9f4QvlHBLFGhRLfofYAQPZfcoFBN2D434GBxSw7JlRu
XyMjcpGQRf78OSb+joMxKQCLI6Xb5Ha4sikHF/Fwyp6xIYTW+uf6cKMQNAP1494+cVhaKzPjjx6t
RQU0FLoT91XEbDUmnPbomJ5YiIQoOuYRPxskxcNxQNmyQmM8UP08QtkDgIR0+GjWqjRc1/KAtamb
IOsa0TguweACZLelOSfqv8AvENQyY3OicPj9vVZFfobYaciAyceXaHk4JoYfT6fDTgnFbvdJDMAa
RMeGoit16XRLWaKvZNAVQeDKLnrz9ZxqO/zBPCdNeoeIszfv7vWMcsnYAtxKAKQImWOBta/+DuLx
TD6vtMEV3jH2Iu1rf+3s7qx6B5S4toqgXwKqj7sTkbMnozhpJshi7mfYSnNNPo0MR/r9J/t77Lfw
rVPLIJnv0ME8Y22pFODCtpj7+5fcaungrXfAzwU1vccUVCIGhH364f9USvehuMiKyPK8oEpqqUx7
ob4t9pgffljkp4bWrd1zXBSHBHvEfuLA+gI8yFRTISvxw7l0In1/COXD2wFIt0ec3edrZ323ggcd
bDqdEgc+SyQLxuZr8ins+MyQpu1PCPVXHXinUBUomvG0ppG3oO7US+ZA0fa0gk3N2l2VclHMvirx
BgOfoJ88HgCaLI9zP3MHt+K4eyToAYNunC8bemJwakJX0vJd47iWPGoME2G0gh/Xv55tpwvxlOG8
AQGspq7mXb9zeuW/InuQcJGVbSmNFEURskQ3wAYJ0CtuVopNdsnXBp9958DzVehNEZ9ZJDBkSnbQ
L98ipftJPxcvAJknlN7sE7/sbxVIOfq17+5VFR6w+lMBIBDIsGO613r7PdQcGZ0QaCQphxjunoi+
WgoMyxKgNLNnv7zL9Mml4zNZRdwWmbBsAlmw5hJi4lt9hhe3FTImm3zr3aPDyMQJvHo8CMdSIh9M
EJyw5VK86XDXHhLOaaHgXPCm+ldbx7IDyw9lCvrWgNYQoC6174JWW+TRQvzkKY9A+1zK/B2PId1U
BErf9y5piMeBfnfcYenMfU/ofkeOIcZlHc5eoMiOHsItjxQI45Dy4FDLT5cuJK+6txB/U1F3ekd4
r9M3VBZN2dZoCoixdB0ivTIR4xyuKhHevBU6vGUpQtaYtBCPaQrGhjXwDwTCJKxmJdN3XQPA1LHQ
uIXqv2Jv3Gj6Ko9PPrOq/J7L2BxlV3A5GZM9JCBXpkVmzLePNggXjm7IsaDWKNO5Jczz26Of0R9w
4AIM/3qAmUTTGi/XFdSU3Ny1EoVfAcvrrua3QylmNakjWATARiltBR6E9QsaGEuXdpToXMT4OB0m
0Zm/+9FL0S473hceGhP5ETAmrFsmPL1Mgk5yMI6FGsZLiTM87KEK881d3dYtyOgnc73QVhrgpeWg
9/v3zkMsJ99ULlaFmaxLoG8tJQVZEz4z86EUYoTV+xoHpRicYx5Cd4FWmW7QmckgHRqH2MXaultB
VVd+8KbkyvtgW7IDuGALJsUETwiGa7t2B0Z9UuTcehqcSkRQN61tkj0I3Vk45nExIOW5GPepZpnN
Z+PLTiSXadBdc6fNm0uKfP8WGKYZtajy9RsS6mfxBdvTTEgzDgJutHMFJRP/cTO0Ro8cyVPPW2NY
/34r+DAp0H6zBsK5MseOQSZlHrNyVGhTRErPtVitOz9Jcspci/+48IncFe/e/MThaXY8CbOUCTM2
8ggpFy60WZaH9oGh/FgNO7V2z80Z3Nf5uukpv+2+M6Oodwt7KX4vjZLXRIJowXPbu5kEQB0gk5C6
GTkBsk5yk+CpAuLc1XZpxsDVot53UTpGnAoGMx/MJfOmMyKv5QPYjFA8FAzBNfQJzgVj8jDjhGf/
kCz+tlV3ogsOkiFqORFH6BGlCXk0Qa52nKavkLOpAdjF9ov+j4i0N283JvZio9X5HlkVsFWb/KyM
cC80rvzA0J1GKBkQuj6J4udSmRW9OBrt007UKVG47ZSupjPyNFw0QdyCfTvwrqzbJ8mH5nQk1a92
NcIGhN/0Jgrbh/qs6DBNLjAUAVFormNf9G7DL3xNGYswoSeR6kaighyWH0zakXApSbQuNDlNBSUa
TRa+hb9XdcLE1mM4mi5D4uSLiOiQ3lmBJ1sxo5f31zaNGNGJEMqK4n1WM0hafe2km7tati2NcJlp
HUx8nNWtgHUaT2+3vojeBa9R/9KdH+kFJGGbv3+7eYa1/Dw8JoDgSjZtKe3Hd3QrU9yQ3kPJ9nS/
n5pcWiq8ZQOImZd+78Rm7Xzx7Svg0tufYYhLlJh3A0v55BwxCGELNVN0b5xu/YIk+0auPbrqzqq1
gaAQZFMpCMdypKkVirJZ2vZr09gbAoZtxE3oDkQCKfxiaNLaHblZ2Di1KH6HI+kcG+rob7t/F2VU
P/rHcqw0uIVM8ibrU9VD8a/9yV1aHjKirRHQFgHb/wWf9WqtdVCss94RGOVC08HMRTYPvLUNkU+g
trnQe4bcp60zFda342FpgZ5rv7nu2liH4NE3bi59PY1Q4myzcY7OyEZFeVk8aM5prJ7V+aTITE1s
skZDqvzO0FN04GbLGYj2i9pB80vwUoRlqd/z6Jay04GsMzwayaCr7FTz46ao8ls/PFWl4J2NS/R4
LaKYF3v0PWCAh4KBlmBH+xJRDEE424Uic4/IoXh5otVCJ49AjAOJSTcRVqEiQMsSFujnLQkpXRI+
c/R7X8XYTwAX1dqCC165B3oJQqenf98MRHuGkv++2ORZU7osKSSeNSofrDtyhXvVnLhawbZe8l1D
I8aCAaVCVEvFM5IVhYot5VKZm1JNmnZeMU9RRmhR6k+oP9QJI4ergpF3fW7bLyx/KO+RRxpsqKLy
oT2229txMXG0qc9jGWk9jALGcVD8ZbOzHV2dQLbFNL6K1R5/DM9hOnuQiMykFSVHedMkvP9AXugN
OAmIUzlpUEMG8NS3pi5PaxNSad5/Mzj906T2/OgMrZtwwiF5Jednnn+0LAd2pwDkKen16qGoWmz2
iDw3CqlEt/rwxHdVYcB2ic/jx3rok9i2jmgeNeC4ODBe6Vxx3nVWvLbfggtzTlHjwM9uqj2Q9bFC
mbKHsYDJml+cIp/H5tbbrRuqPJVg1B6Tn7BecKjtHD4hs1y5QGudkNrsQ6mBs52UNHb8O4BAR/GS
XodxigEjH5x+xp69lzwuuujLJyH4EmLV0YvQt+Xs35C5n4lRzn8xTpOREKIpOe0jb6mrpUdfrIsI
K90ZQstwpsJ1YW6JIIWYpiAZELSrIx4790anUQqbNy6G1d/u1ycP9vYeFN2fRKRMH391+jQzeFP6
K1TNZij6NJjBNSCKnHVr7g4GotY19A4mn7N+t3Tl4jTd413uaGemIJov3MZnmtadQd730EUbcvYG
PkC4PA6inghcYH6v7awHv0YfTee0zWCtUTfKT8LEYsKbRrJFgOv+w15zGxN1jjkajKo7rlbWiubO
VCp/LbLecREi5bES2y/GhC6KkUbnJ/h18dYtcdd/dBFJsrXTnXjRJBQVESl0J9G+Sa91EFkr2dCe
AZqlXv1Ul8mRA3+GS1EPpu04pXMEndu+YpnW2CkFvAiUQ3ugmerLsf3iMEtsVfz/chj4OGrn+Adr
LpjaOXdPo9Z9898NNAJw33Q1k6YIMZZTrh3DCXiS5gWoxLxNDKXO8er645jLPN0cy2uFPhH2jisi
CsxEH/rtuEIr4C1ecCRRAm5uNDnoPLsVP/SG+cxhg3gTt0DYVB96A1gisuMqWwdt+WZWwHUQunUI
sa5bUHlUXXKoA3IMo//BkKItjOiIjXFkpurtA+knzVOI0l1iy4ZqW5Aa56xtH4BLOMwWfEXSvStV
75wL8ogd+j5NTGwGzfz5KQfcjsjAl88rkng98ZjACrE9Sq6CMtLjdAvdOXWFKlLTRLGsagjOJr9U
LjttASo3YjDg25SWC4gZL1VnBev1Dv+hFmCQCqGYSWCiEdpa/9PyMuu+NdAlVQwoZR4n2IljTDpj
bbJKFTl5fce39hnNA4e2Afn6zj3+Nck9OjrOaPUWUbDGQcAgmYp5Icekv6X0JZnzydZF5cy+8QWA
i3A8ggzLBT64pSPfMJXlWpXPUR6so047KhQ6wPWK99UFH4kEx/lsPYo5acYKTdnHdALtRiBL+Jow
kEHfILQ7xKnzDdaJmiMdPcHZPgUuW4KFninmz/mp+xqA3eYQvd4yfRarBVXuvckKsmHxj47P2sy5
YAsNmdN7q6fPN9T8QcD8Un3eALJuF98uNn3UvPej8VIFKtLKo5jr5cvy8CLnNSlhiIBLDFJ/l3BJ
emaKivasompk6TAf22YHyazXiwkOSZrV6W+JwI2rJGxbHaHqFpe/ZSvHKNvyh1qeqN75jGaIeR50
3M9bjMnpDu3rcXRWsfeDh15jjciJK3b7k5cBK3wWaeVRz5f5Uf1dL0oe/vnm/rPIyl7W/UYLiP5Q
e3DOlXoxnIliam9wwkDiYRgR4nlGjn8XaXbHwm2pjjIgO7mbntSm3hNBt7abyMtiPHOEpknKRaTp
pCHH45yekAAh0n/BTcR3+NC5QfR8KWdHkivik5+vJnu9Q+db0R8k8pwxKWvZcjAWQn+ZIzeJQ0vE
fHkUHcInyDF2gVupSPKXFSsmr+z+y9w6jiQj1QeryVHbhxCldyoZIG7ELxTdyiIBpLQ5KL49p0cP
Z4sclFXFr5ewzhwaokD4FZO4UflXP5xqxkfjBNO7v+WLJ1q4T5fNwUqi9AQJ4q+zAywo51s2+QYL
vGCtqN3RhfLaAhxgjSPCSXQjtPlLZZVnsk2iY9AjHv3PiQn0N+r434tYYtCp4XjGKJfmdhg0POg6
tKQmsfXacgRUSCQx9sK5o5DJtQZH8wc6w4VQ77hJ36Af++N1rDgAabTb4lkHE5qri+GjOOxYreNH
8aY3SjW9aLvfF7grr9q1DgypWKK9mybvWg/jHIDISDtD7u7qrnVcfLobJKWZmjkd22XpzNltaKdB
Aij8KdVyDBaOQIcuOWwVublroJ8To+/KQnNwEmf4vu63DPh52GF7jWWTKLlvSbSFVoCWw9355xht
BAk4myoQ5/IEMgvKyiyvht/48T0++7t1okHycIOzwr9ZaqFxiYDqEKYkWpVvrWf9v2XIBriCA+AP
K5Yi3/YbyREeOhWzonSrOm+qqDAOgtM1D70tes0dRNCZ2gKFziRrDe2Fi324TG3L3Y5SKq6e0ivu
wNylQhVUsKTC7M8doWtPs/Ur+3bqFWzcwVl6Pua5kHwo4frgUzcxQWiluGSQyE3NSRaMupT61gX5
cwTWhTc2mUODrB7uQZ3wiNlbXmuUzm6jwh4fORLge9jWdAHPnU9Opf2uNSFCRIgJOGKb4wdTIsFI
7H7JzZJnej1WSAuKpd1I7TOxPxB86uVxW7v1po/xEwg/3sFiI9zppy0sCRr79XC98S6iPb7EhTuO
rogtv/kv5T9Z1Cono1poiY/+YcNCiCeu6hBU5KbYM8Bo14G4VGinjAdhNO0ggLoojQg4jgWSuBaC
YY8DBTkNTXO8R2zTRkMRGUurA9l0oNgojQgAlRmptFUOARGUZxUSSbGfo0Wp6ZYNv0FVlBS07tvI
CGoB8aNArIao2QaV+i8cQNG7sPX15mbduVXGQROxPVhMA9kgDXJXnK1YGF/i7jDewmJ96d9F1j5R
pzEcA3z8ruRdWQrm8WFasTyQJgqpBA6BmtoxNE5/y6xAL5Xrd4X+ZkDot5DCafCCBohfZpNP2zva
D4zuMD0YuTnaSDmgmclqBmiSabugAPP/ss5uRhAZm/7gWRfHjYPEtj9nWujG55jP4oP/QehFVEn7
bhmazkmObasQhNxr3JscPdIqcy5YdNlOwGGwvjCuRaUQDywIGcRIR+M8fd1xEo3Sy/FWyqrT0r1+
rRLKKo3bFg+QenL2GzpGlMtq0INq0AEYvg7IVe2kd82v1RapScyYw9mXSKuocL79UnMxSKQV6ZB4
/rTEB04sg8zt4Ewg/Klc+XlXhbnZ2fw1JrhCsbmsfog/JO1gN8NxdMfWq1qYER2B6Cb0cfkM9XP0
9TBM5K0WzOW7wEFR7Hy5NKUc51GOxHB0uBfY9eGJl9ybEz88AY0HViYOqGZBCM4qKGU17w02vnaT
YT0AfOdLqRYVu/lkT2l8qOv/1i+CghBzOs+3mTeP1J+VfrXlL/O406D/WO1muokfPKCDmObn0uUd
1v07gCpbqix4vTVBs1w5IU9VWXTLXDSaMoBWv+jkielgVEdsVWm4nqnPsgDIqVxGiqm1Atax71yM
PX8snl9iQG2Ou7S6zoUfJ/yNoyEd3mxI1sTe4pZa0raZ94M+kpzMtqxcXRGrR/IIRjmIxyDQMYzm
bwkYsMZjVsUQ6Tch4BCD66GfqgJYYmeLOKIdYSo56UjOYBJi/lZ6vT5n7AWMGudughp5oD5FDAFi
pO0UXDNP3g4d7m0zqp+Yg6wAj53GOfoxPqbkj8NraJacbVbb49p3vyIZAldEs/J6ZZKBhM7NT7rI
fWmFThDBHGHL+JPpX+x67F0uSdE5dPXSxkK7T4djYD1yPaN0B2M7FJ3jDdrwRYCcuiFmbNqMTnoi
1ggzXREWB+DEV5+h2M1TmlPZbmh6jCPPgPfv+P+BLxrIPwvRJTXz4hlTg6NeiO4Usqlpddyxx9Z7
6/kHiQq50zArDRp0wHuXp2dOsgl+ON77r05J17gL3WD+kRmvtU0KHTmvghqThqTz/fqZpsh6308y
3/VpGKWSRioyxqvM62jmjbgFY+S1NrpDJskVbQvyJvKd9rSxA+kw7UqfNPrApN0B0Q0bJ77UNpz5
o81+9e/+dtB/G3Ec1y8WWUe3tQ0e/dyNCVcrZ4dbkEez7KXz6lrq40vrkIDxNn9wl39BltRucoqx
wyjEZ3N3mjsKFeRnmSdeKywSgvxyXwS29/4dXvK5NLAtQT1QMzGouaY6f6efivTuIg3f1AqxNa3P
F/gvfv8xEG53tuCQahXixCt7YfNp3aEpLLmJ0svWYVRXmwAxhpyBapntP8OyB9b29VxJu6Y99ilj
mxwzECEqz2/xXwGUZFTpVtLDY+zy8gq+GHjlpyfl5z7Sc+7nWJblNle+PVEV3hXCl8NMI6KWbBMa
XPslkAN8c8unJ5brkEN1eZqPqr0DRr2rclducC0UlySEZuZZdhWcd7GllfcaRH9r0zIsmKeN+qsy
gpVDg2anIdb1io3gRdcqaDtAoZIW8d+G4a9zH48ep4LYoUPJrccT3m+Zg+jt5qxs3udr/bYddIOY
OeRmMhLYO0h3A4YZsahl+GQKcsCGrMlw1Yil1rWSni/qDItetOIWtYqj4nNxzxrN7FNl4LZtSTT6
AY3gFn2zQHyIvVK7rsMPUAbS6Vug8pcXgrMs5/WOvM9PvrahAVIsuRarUvCQX0eelTbz9ylRmCI8
rN8jUHTyNlIb0MZrDFklRSHEKOO61aCg690cqt3RP1VVJhQJm5LeaW4nQVdWPBrivjyhmrCCrjqN
odxAjGCtNikTd28pw935XFQBHfjzWfncmU/OlwCTnuPsLFbE8nlknZkPxc/a7EsohxoJR043JnS0
OEFmj3Dj/zpYi8asOJyaxG6a+6bMEL9c4Td6vJqNolblzb1Vt2nC7cgJN0MEqWX4Mq7L0e+TYrFt
p6I1Q1vJaeY44+s40GqZTiz7Y2ui9dLjCyN6vnXRegboEiBnTR3VriR7l821JMr4f6CbIIweVm81
7gSEWMyEADedXrlH2CyBw+5ynfchdxnKsxXalUs0fd/H8UBuA+SYFVeMV1LcZZFKJhOY7MrPEQH/
wYVFgmJbBH33D9jk/YOGUHCMC0KPFuJLUr/2YI49IxKWewLw01Hm7XoIHOaP7K3E+NrcgIXj/INV
kAYHAEIjGt8EE/XH3xQ7Kt5Iun6nWHa+CJ2+i3UtNKac+RHByvkQJBSVBWWe49MD0cYK78yADrle
cBJRWhVEPvct78doCVQjB5+Cb/eFyTB43C6bIBmEJHyvcsWmWR2Lpp2NInY5QFYGbwfWPvZqWnOi
EQSGV3UGpla2RzQN2zSD7j8z3DDEMXFC8PpfZ86hYTmjqHY7gZjazNpkbrF0H7YXKkUBKZ/gM6ZM
rvu6EiMQFAI1S2Xa/Xw74XJf4qv1SCcL4ILJjdncROOLQ9ta7AwPN46BO1VzCLU6ILCmE7IG5SuW
2ZrHtA12UegD6rbiMcUDkX/2Ba2++mGUFZxRL02F3sDSuB8BQZi+Nl9xbfyGHUFWFvfQIpW78KdL
+oT7Y6LZMZJTyTWRqcX/r+905MFhWRN1VvCcizMkTQxEWeQJMQyMpu/aHaQJMsObuuX5ycpkdLD9
NcBORQ5LczFi3EJCxTRUR/dtf6+ptvgqY3YHBOdm/oZSSi/y5SAKTKT1sAaprV/xmjtH1OZc6WqC
q/aeDvAB3Mic5vqGFNguK38Y4FHPty0c3JV0jB4D+gyN3R+uK0tRhlpn8CGK/1VXTkhA1a+BmGNv
7stO1GmGZlYk627AbmR5QaKAF0COYEarreyCeC4bATFejlwZ6/u+M924gosAL8gO8UFfPq1m6pAM
OVw6r4NzYfoQ9ODftc6ZgnqbCWYQ3eM0NIXu4EHmVIbhcAqOxLecB+LnE+MyFNkaAwHMXuqeKxjN
7XLGQTFas56faX2nL3iidk4hw1I/SHULs36PCdBHWEex+buqx8tW0IBY5yGaBMluFnrIpFqV29ps
srHDIDCl+zHZ0Br79obUJFaoFfTi1dJKToRLkXXS9trNqFfOuqb7i3jSnueRFZ2OUom5lnWZmBjc
3xlFglqdfuhRpS0tahsni+T4mpGbg/cvxUewUv3xYWkMlFxOqK3JtpB99hiDmc6U5Tnv7UclxrW7
qXeQ3CR+Gaizn7DcNReCeDLoZUerong+axm0wT+Evhycu10HEQ7ZdVV247C4P/e4+OGC973sdMW5
fCN+d3JdHxaF5k0P1HqOlrooqPIOnZLtCGyq96CqFoUcrno45DX0Jgg2qVnMMyvyH1oA7vBMcPtU
otf1zhMMDGU3K4GvYJxf7lKfh6n/Cyt6BjRBQWqCJQj3hI/XYKDiTB8BAK8YxE35l+KKWh/yVNtI
TeVKG/NG8ExJ5vqgsCdb8LnNpLnfirPtwrrjMAKQmMpRDhnRi6iKfgEyho0XRs+fCQAFQ+N+Xr+Q
5CDyJ1sflwvR4h7H5EPyzuepMph6gqPi5ZObxMTkwL3jzgms80oNUArg8WQvg70Um2HqSOh7JUW3
c1GZC+maF4EqFMogE9npUMAowPrH9C70Kv8VEDH46P9e54ilhhTNpX8A31lU8AR8tLE7fG4QsYsN
0jV+n1yR8PN4u3LxBOYJ76oEaxBZRBuuaAvcj6H9eD1Ajn9yYKwlZMTxFYyv+zv3UeXkVCD+5Dl/
DNMQhHEi714KXKVnaHofAMPF4eE3WNGfl4dKppz6KKTAI+UTfp+PzasjwqCzv95UMgjnqwuRrDH3
lYQ6DCfbEdrsSj+tm7WjwVQ2C9OEggmxIuIG67qubckBaADgmBjIbDwfc9V44UB84vzKIJv7lHKh
2y2zT9w8Et0TG4s9oCXdy+bWd99BACDwR6O+Mhm4pRcqV5hKgSce8Bnibs5ODM3SIE0B9mfL10HY
hOWM04Zijti2Uk5l4aBqRLRo515jNQjgNjhrUMSmFpQ30ws8WMkY5LhLBHPBBmqvcDszCFm4OHb9
Rz0jbiReC2+5vvGsXi1fjyUfHQOx4ELsPqr7SVp4Vk/fVF02PEDDhzfViozhG2XzD4MquVyHrGUi
JbezPaXScvEZg+MNVpH0I5qg+nQe+upMKBLM1icxpKvoV6px1MeHxi1r6mekRnpwPypijnOXmSY0
zd8IfgbgErPezODnXsWkNTv+9B5T7U9LIYiTXVKJnj91aMPDYqQPu8RYJj+EH9bHhdos2dGxheSQ
nHdwcbaqpehc4w4k8tk1w9RgMpuycd9WLg77oMV78jQh3kiENHHKhtVaAp2lvmAvhixkXXAaKIVL
Igz7kPWu1J/cTMnuwqslnFHR7pV9UUaGiIsibP0bgBe4bBFL/gm5hRzAhNbOBfzDDVsl4kxiBPQE
gLaB8yFKPpKIf2IxnkOOaAdTJPHEBgRVxE4/2tjA33h7JSizvVVv6H2wMA8Rx+5s6L5cN8UkLVy8
kQRL9TrHHusNyKZMn2t1g2nujrqBq/0kPXWnxEPvL22JqDOZhjGpE45RyKWcj3LOHRS5prdqBBQU
LVbzXVdy6S6qlkCwAPwPSVhb6DqzokJ3Ty2yeYtQyeSZpLSj6rMAqJirbWDBeZklA/31WaP+hUXZ
0nV/j8MGksGpQieIlSZJ0RWFtH1i4O+2KgZwqlkry1XdSLbICnVYAP5aL0InnJwLeetP425xobSw
v8eXPUUUX78iivMfUK4SCcV4nhnYFb74YAPhQxM/iQl+mEpxU8CU+I/vhSJUiwQF2Ol0uCRnB7FN
owSvcQX0wgHB3GXOk2F3VbqMTYV4XIsrmrLarxsgFn4Y555jkWj+kOXoK+GgzwD/oYw/V3VG1I5i
Dj2jW7avcY5fMjqc0lp3v2LkAVIY8USWLmiMKoUtk/uuE28ebVJOpe7bICU6gGfK0gFdG5V6pwVG
lZXd4QXXlizqy1In6nYkWt2y+NEEOUwdFo/7VL8y21yLo3L8DAQdH7CTkTAwraAp4mhY0T7QQE6u
kwdqIwLoUqaVa5Ce7IpHqAyTsVpss/g5NftLDdeKqJJaGcDI/lILWQK6OPFH0q7392sBbMQZyO9W
aQLlU74BzwlyQSh9JKw2Zbmpx6GTH9lEnRfDhw0LKddWsYip/c78+QNrhu+I96jxlL61kKV169Cd
6T/DuObdYQ7zMpnWnj4AhsMTRddlFpesfb1t8bqdZmO/bqnymLcKZq5eBO4BepkxZ40h4NugucTs
AHyUaHS/nQ4lq52qlfiXmfXMdpoKEDpLdrqHxwlnhQ1YOI5SxPLAXVeUGvs7I+gmbQmIwGm+17Fo
eco1hQV7IyBVGx3OyjI/xAkuj98lDShwGxT2NcnBPdskpdBOZNJmknTm3mtBOZ+z4sFaoljPuVJx
IZrvDIN/0v57/HHUY3HbrV7Q4apmWkyRMLPr2wEYj8ie6ZTf7J9v4auRxlGFoYZGStrP1c2KGOhB
4yCUer2ybJUckDy3piJ2jidsaWdBpjULduEw/hFhuB80NXqxcVnokMmqNHslrcVisacFclijFqoJ
wLn+eaoXWuuR9msKkxo/3GJ1NvPr4y6rrIxJ7CEJC+yNjBRO2eZBL/vnC9wCW56D/JU189yFNrYx
HPY9nPFvaM/np1Ms9NWp+h0dAzaFU0Slx0ACN7CwFzLhS3ILOOdG/38leSu4ohG4RrxJmqGTR0WL
wXFpvTx2oGDoXMPGgNGsRk79QY96DIeP/xHjsE7LgAIRXnfzFcHJuRsa19Lsu2Jlw1NnxshIs+4q
B3LUxNHHzf1lBI32l3fBe+dYahso+sv1XId4/1uue9TMWQ/4o3MofoymZezHFStl1VZ4WtrXCNit
axF3zyjOxXMnwSx10xcTmXTfW8fgS+vrEF+1siFOMf8LfeHOP7QaDnkTNjbhdog8MyYx0oyTlJOQ
J7yYTdCU6zJCyzQ7Qu/6XkmPiuhy8mAMFWC3iYNsu+JTrc+3IveFWmBFlnqTHFggV+YF41mdlZwG
kB1ZOkjSwo8DzfN/qtGec2xau/5D1DnqgiUTduvkKTvXBNQNo+xxZbaNx3S605+OTGKXewzVFZ/B
/GAo0/k7h+05cNyLk9WjZioY78LtKzjzzwG785xOwWYX4l9XUL7cqYGc247gWSfvpVu1++2UoiNI
WYRJRiiSobmvKAUfiKWmtoLb1R/qcLTsqoHoXgwZgr2aEiQE5+QrvQ93EzVxAPuk0LwDeImZvlX7
qY5Y095+3OFi9WLVJ8/rrgW0h4aUsNTO/eDdVhUumSSHfBp90s7b9JGaYiYxyhtswOvRas/2F1oQ
BZ6wg0Z6TpUYmI6Kc/D+65sGLrTTgJvcL7kgZ3qjDX8Hqysn+hV9gcSR0YlkZKzaHOpBDVeYUDjS
cPvAaD/17X2vd5LItlXE19J11wJ0GQa11qPYPvpax2RlTj9iqZnmRrcw2TE8ary5HfBsVP/Ww3bh
wHEdrLdhDl7vlrn++lFqzsKNdGAvkyjdLwPqzoPxQy8bZS4MEbv03dvzg4F+Vja0DnGjhxxMINjx
oIZuEMvRyMANCaTJtHOZI1w8qSW6ABETOOkYB5Y3J7NleNeNDqsOXHB2dWOUVMzqbrJx/bNcAK37
q5pFoWXEVJmaYbTvwqpVv86Zfc4XjZ8R9y9t72NqVY/tbSRprYmoAgLqnfwM6azczbhXtuDJDa2L
8JkQJePMzZPvkBUR92I0tfKyECm5OU0ZPy7LlqEtZI7FPFotWGE6T0AO/zlD1FtYntSkNAwfgn/J
LjibNAiPsinhsL86pVhWOxGtMI/u4kkgq6LcnNYdRfIlvE21lRrSeBdq+zTF/pC4jqLQ/y1x0nVk
HMXaSSaQtdd2Bxwjhmwr5N8JnqsrBd/6o2/rIjtQhvHOae4bcuZst+8mWWU6oeLYXI67V5uD0PDC
8YKReRdeuhpqTpV5QrPtaSQP3h8r9uU7r/I1qSEc41B9gkEppPx4dwFZcFNVXD19GKhzwFP3by8z
NJ+HPGRW+elOBpvuuklYrdhk9k2DdEzL/DQcnUFjWfKCHyY5CuyP4TDTxFlNiFpJ13mDzO9yfqq2
3mt5IzpRaHXG8AvJoKxtt26XqQOZbQQhDVMyauXCE1n2jEPw8KQ6u2Pyqhv5NbuRRDSl2ZejvMs+
gBqqEjQ62cBYgx+mfLUO5xjrXzrgoSu6JqUNYNg4Ut3RwwYIM/NCaw6XtSrhQnDiaAvvXq/Yts9W
/uSmKBDOy4BA1RTpTU7OxN6IxDniQ7ldyVQ3dOZBX6+eQtKJ47rHHiafvegC5eshyfabEhJGxQa/
VP7btyqH6x9nAXZ7QvmTKtefQb/CFk3volGpS5ghBBAsCdeOMQi2uz+lEPp54JT2ktQPylX0/D0x
78ryI1K+WaXKI4bWFKCV9y10yMz6oFitBGqq7h5Rw3Ezdt2NXcCYdqS7VzDZ6NI6ey/vqTkzhi1B
azb4PmIT7ImtALjC33rKcpd93hoynX1eJQV9KAo9ftj/dIx9YMOuUyMHKjn1KEr68VsuGj2gwHNw
SOf2cUfu7d3BLknILhe+E/DlYXjn3q6fQ4Fp2wxaadjcB2nVULAX4Pvfn0VvuAS01nT9kjXDRgkl
GwFRU6gxl2QhBnNtl4SbKy67rVM2L7txi4s8/nqFzcDvaQHMR3dEzzDBK8XebAns9sJldE8gpWEB
LxXKTgM3lLzVPD9rp6C4TloEXM2pKcQMoEYDOjXcVVZLHfoaF16kXmVxT/Gpl/l+9UXdLz4Az+xN
TcKgYa/fycSxhYjw4OPMblxnRQwPlBv4Gblg1wSWsIeE+FmK+382bhvkUkgLmaNyDNkwtHcuGGtD
jA2JLuFdtML1mDbs+OUI5yEU53rLLk0u/FmFF2WjPZgtpTsY74ScHcXGcC5mwNaEyVtOeOyxH1CX
Rn7bjlXVRbthShhn4uk1/qyAzzCUJ0D42RThnbwK2n/pw2amtmWZLTUlIjt6eC3M/twVV5Qsu5Q+
gj5NCAB0fuDECkQra67S8DZCKNBNPcL02HOXb9FQ/b1AEvkYjaVKnWB08wz9yD9r6K38jUkoN3sc
sBG7YX9UzTsS6XKxaul6RULLPqCud9yGdk4l/um4ETUoQaa7GSwrmtoOFRreEzBtj83s5Joh5U4Y
bTGFXobnJ0XrKeabFPma25jDUb05Fx/p9EtwjAAKYJBzoXM3EzqMVzzBJSJvBOxXx6hWujpjEBD0
MsJddWohZbq6pdbVaWy0d6wS/iPDwi6fJKGi9tUlhvMqpWxWRicNXZGr3Nxr++yO6rbHSsWMlkvS
OTdgFSXBYJTgFCuFj8lB+HPnHuqSd47AuHwfRMHjhHsz/O9UevotJCRBBwH+AWOCiw7vE9CJHmPu
6dtaxJzN5ENOE9TQZOllGGu9BvMCAdlFTdZw85vfNYF9+I6UWS+5ZbMu6pOd+Z9tMDwVkXCY5UO0
Zhc/4bppORUTx2FpMsCJZjhPByaoB1z9m3m/UffuM9l/ySP0UWdCU57QPJD8Un3atH4Tyh1ZFHog
C/estermniRqxlOhX3Nl4DfZsR/vbR5hPFSWKIPhqItdU2/OBwXmm9uD8hBR6aKlqYCvRyOrnkRg
2A7lqUsME6nSuoU+SNBTYl9lthZvweFUvSDnLLdNCnNpSZ3t+3ixbiCbP9vRNSLfwNkroYQb/K8g
KZOySIeazn4MsLaa/8uczUu+RpyGfvvT17SuYDyteQCE1eSOb+yfRY6KqAcPrmaCBOsJzL+bznjJ
7W2LpLXHEdexiYD6z4fdX3lEYT8O4V8k4uzu68z4qDqvs6041d0awpNSFrJSAE9cskcAcwqmJ9la
BSqEFl2WrlwWLj0KpRXyE9yZQ6pXeV9JLdrlwLtMlYVGymt9tElRcTyyjo2FPc+JQt57uhVWAjJy
Qfie+/DiU+dA/8SZRZkSLhB/16TI8SaPWFNR41/Xvi3/IhJegtdRpnKCQfsgwCYmd0ewY8j6HwSr
ecitdezvUl4upET9XV6Xyo+YgZzOQXzkRJpXwaTwyvNCd9tszNkqL8YuBMDHrqliwc0rcpESe/n7
B2ssk3LJkWrz5RAdEXvAVuN6RS1f/DMNlYJE0G6mJtc64eRarpTr4fREypGro/8JkVlrpWA2j9jZ
E4Bo+mEzpupj60Vu7VWUKHbwZIRlruXxKm69V4DHJLET0ohgNHmtLJWMO9x10PqKxT84G/CYI7+3
vmATkvJRBkHwrQgCnbmIa/Za34pFmqnQGn0spKtaimeI1ajLbJc9au1WMuYCa+hwQysYx+ss2g0B
BIQOOz1D/3w+aeT7X6kfGQdb0Bw44o9od9vfcCrHDA8GxF6lFa3bm5nS1/1ctHeB4+Z10og8C0zd
dmFr2pWeZQqv9vyrl548a0gPhuy7B5kCdXoIMN5q7B87RwDXKSnTClE2wPuBb1TeCf8788DFkZIb
geoVmB1i6IvSa5NbfW+sf9Pin1rMifOecq326ziwzFCa5p5n9aEohjc1gyx95b1tMEGF5Ljuqn5+
U1377Sm7BeoD244unyEzVjidcTXMfoGCUpjjkzV6V4bnOvI79+KoTgBXzd3+sqY4KGh5TcsuIzVA
hkn4U/jIPft7Ma42lZJWaztBvsk3z9YaSNbKeFF8wfjdu8LgddGX0J5HvgHHxOwAo2DUjSkt+wVx
vWj0GXhxAKBBOW+Y2rvNU0yrpkwjTYU2bjuv5f8l4G34D69KEZXoOtueSudwrsm2qIGlJVPidAOw
1HBmf/a9q5EciatSjTiCjPwqJuIQEkWvHjJ8pSuiE4B3a7V8HsB9UyylF5I46/9BTNDVRFSp97tC
me4rl5mDiTFZtrHHOIjS3LmJeZtAz2tiq5osvxMdWqIexjq0GtlPhCFGdCA734hL2CGWisrI0Kvs
h6RBXEfAfYWeBJ8U8TIunA+j/U9YPt2p2QD5JaRJB4053rAxNxJS9ZpC7YJo9BnXvX0ZzVOQfuMO
AP85mm2gRWC1K5eSPSMIdC/MHeEWVHlek4tKco/LIp8SDwElXuxY7lomBmUhbRyr8pYzp+vsJ5nl
dKlLFicZnKOEkZUFZ7ohiAL5drJVdEmEBAIZQ10OEs+hGeUZPVjec26qlACtitTdL1L695l7PGpM
/EMkijrnh4SJYdUCgNKeVsjLBlM2RtXbltVQwQZUuYYnikuC41HCNQ+LBnhHiC9mt00yLsnPw3zA
6V0OKo6TycbGTRRnRdXNm3XRTcgtJEfsIWv5R+6908FQmmlT7LIGh24hrTemD1A3f8Sw3bxdknif
QEnwLA5263JSpY+xTdK1Fm6HhA/n2CVcm2L+pzdplUoN99Rhtf/BSyOOHeFZ3J27g0sqmgJvYq7l
CFpdL7PiLW8XRcr3AVnZuE+tMy5dGQj+RZy0jYrKLqWblcDhTmcGiU/Lk1ppUmx/a8KYlFjoBy6r
BkcUvApptgYc7ehUhYWbkKI8UHe8Lyvoq33P1J3xVMPgA8OqzlMejao8vD0BDKAtHStBVCdvgGn2
Ipi7XjzJiQ43DKiJzKCBjpIEYEAtiPp8YD5y3oMPFTGJUSRhwkdpJHNaxIzNGhdCO1VJJ1FsGzhj
biVwsXnLpSfck2byrKV+D8hrn/o68bd2LTECgRfSwgk4YW0AO2/JMhpfTnC6ZBHWGZMF9GeQh9e/
1cICxfHeZOnSzeE0ulZuxLf9PlYS6rQ3fOnpIWVtQ+rIe089878/lCHMODiYXmRlMFIGVBJcFqRp
fbN45IZtOxcITaSBfhwSLpMFtcaR6j5j8R/ZK1yKYpVeQkG3OeSXs5lIAyx55n+lOcG3l6uSZgnr
fG+UnixnTlftzykZLA+frasIFy2vxfxHu5tPa3xMIaiQ0ibvWKjB3YhoFXa10Wz5un4UJI3Ir62p
w7xtdYnj+ZJ+tUJeaK9GoFzxb+R7FbAHyH2rQrA93C4jbRNGjrEmuVu4wucFSi2GY525+8Pyb/SX
Rq2UVaVs1U+X7z77+/7swNcpRltS0Qq7Hoxfa9mRh9YslVrYAw7vDJgWNukCRQPEQDtCDho07Lg8
zabRnckk2d/x2fAeoQOwvlFJAbKL1DZqbGYc7G+7mJtL9VoyE6I37VgXG2tqrb2m1yxxg4OBVGjZ
fGLt2SFYD4KNaBbrztpwAJ3rcQvLsobMPNLZYIa0I1uG3rAnUEGmbEy+Ng2n5EfuRZEgRptUxtKX
vD6EYLrThj1uuEco9mY9O33QAKPb89b8vTHYzrvzxUslIPlu7lW6qsBjbYCsEbWN7g0LdFyyCuzh
48VDZewUXSuqSofPWqVRDjLhAc7I5cCmigIGGYFSK50Nk/xurznUcUXS1NTgHLiuhEVAxcZgZGVO
/XSgu8zb41Ojz1DLvz7+IC3d4YRgvubxQOouSnFsRD7RFnGA19fvvaudcziof8gC8FeBqYYAiLbk
QLbn1GlsCk40wkTxo3GnkIZja1tgjhBhMG5X+CTnXkw3kYyXpKqGR/9RmNoq8PEleXQgBGLDJoOE
OQW9HhkKY0e5xgxGmlwJv+WzTHzotDcRzR1PvThGoaa2i+3HE6/iC0fM0Ba/Amzi2e44ISx3b7n6
I85DfmKungDYJwnyZV6Log1XgaeaAwJuWkQgcPCyd6eg1JwHLEckxurXhTKGCajffBQGx36ff13+
TgjXFdr2mwc0vf+KAZ0AmcY3X7Fy3bQ/ayu+rJ0SxoTDm0g1ssg115iCMQJ2dMBp+w+VsYc8gCby
YqOV7UMI2J5bi5M2O4TrybnuBmOZ5umksQjfC6YjvWnU08eh47s2a0jakdPXP5m4Rpbc227VnifY
wMCDFR+9M/K2oKI8lWAtKfyYTxHicuOb4sVYLLvMBL7/KLV82ZCgTA7dGxT83CgsshSmHRiSbffF
l7XBNSjb76bnltFcFISuYVgfxOCQfMoRMmqanRMI+Kb6o0oobO7HZmomhAzFe4AbhGYBzp+DeD4G
4WVJucmtcqeRFXmajYnA3/1URCdpiOe/TKWMNZLhtzi1d/jlOScuv2cWbcoow/3OaJ54Kd0EfeXz
ncaQA9Izq9efRZgIVJM5uHhIW0fTM4o6Tx0ktWmuwvWY53wANEHGyOEz77FuuKRGfZCS3Y4neZ97
d0nGxWpqWHj78kRYPKHb1+ysNahCj2Xw+4iyz3xQ54DX0AJ2lZEQQ9fOKvskyPX0N+m3z+Xxec87
Vo1bxI5a9NTSYavUxrRJgzXNzwsWYh0hwQygF2g2h9pXlktkyRs7tJJ8T6FPHu4WaBZs9k+3hS3M
p3wh+WvX/VVkoREuaOGKhqsG2fTgtCnusb9vmG8MWLJG6F7nEwW8k22GRvF1qbjwMH6ybmqhznMs
B5EWAm/HzwAgJBgL+QPyLZqjH2CjxhwCselX3KERlY5EQ2cA1xs8nEVaXAAOQaozi2/jCDwcV5kz
YTw9uUPJPo8lIqaDnbG8UPToh68m8KP8izYdoQpCEK8MEqYk1Hb/64jd1ov4sCw0T/XM5Cq6NB29
s1c7PS8/nMWA9lF0JsJhAWVNJJL8KrjruHrb551pZ6fBFFPTYhUSTAEMxHKvYedLzJuGXp1fIHNr
1uEPl4MaDkWDVLX/pj9K0YMM6a+OpCwj15e7IlTrA2SiQJSyIMxApIHGnPfx8o94GIy3jixiQfLj
/blc2zibWiYcf/dyh0aKg7ywXVB0gABO2DIl8bNwXRvb7c/QiGm9P5kO6J3P5YGIewVDx5JSvkbV
9+sJe7JqA+Uf2bsCo/5puOB3m2pwLpl+oHu2STWV0/j8v5vgyuJbjUaJQwXb7aLw9cj03doAvAFz
aYxBmidMKnMQ1Hl36fkmCzv0VF3AWySvvtJ1jQmi6nwVohT08ym0V275WLnLEmHazJY7pHupXNQf
6quFAKlbGDEmkS2zdWqlmRLLF9OkSxEo0KFoHAIxD6yRQlDtVZTYULJSQ7n4kOU1Spc9v9ISe9Km
gXhJLH3ZcTr6zjvcDMKbTvXgQYEmZL2y47yxlwcO1TeAD/oqWhz18SKQFbDvehMjku23BdBewFJP
L/lYfqH0kZvR4J2lc+1snymijbdu42gnDTK7XbswHNVuU7tXNc+epcjJSzhh+8DL6crw0ZT2rn+7
3c0X/p9e8vBOXq90u6NURFTQJzHOldOSJWNNDDGSxGcPTHN8QH5ip0S/Bn5VQe8Sop3l2LNhvnL5
imvfzVAJk/gFXTLMrrl9+C6aDrCv3sGa84TzzeosVV1sH24w37GL6gmnOQ0OP+wNvFPQW0ViRTRN
bHxzhTiweMlawqJxqgLRy1VCPP6C+Yg4/FdagCRADhJBQqG9cVVJ4xf2F8IF+DOzUyS/Ll6Z39or
wZ65FML4JRHsVg+SXBmFQhobuCp6pZwwo8rMdq9qD5WsI+FxNdhQHI/sxQIWatSdt59/NIUxE8VP
Z9UTWWuz//hfZ1pzsHZGMAF3cH3zht/vC6uC8t+fYu7sIX9boJmacpMYWx0WhHnVHTkZkWwbkRGQ
Sw2uNDRMhkkOcDCHR6CqdYSh3tkFou/jKgur2KT7b7CxbmNrGgoaBN7zbJkOv1qxiRNZu/NnQ9Ng
0Q4B3dQ83J6RQoVth4khqTtRv5QhzMMzXYV0Ph/jc5LM3uNorCENn7n15d9AfIlyKI2/ayI9D5kd
djavgf11FSvRcN7Kz+o7+IZVIU+IH2H7hpyJ1tvoq84Yqg2V2Zw1H6Ht7XtxaVVXkrfN6zrxQtZB
paxRFORbwzATVGYz6iRBpxAR/aHH/vRBvVkfBEQg9FvQBPLo+V2YQOzyuJTgHV2y3WytBGcksvXS
MX87QLFsbmp3HirWEQ5bQVnaEppC+SBj+y8hZq63qcQSWWrLtTS+VAJzNQznW0WoCL7nRjFWQtZa
S/TpwmhNblQnW9Okdx5CkHWuU6g9gjfcxFd8J0ZKLffjGYhOQrKk3f0bTghISLqFT9KggBsKzv67
RWH+VLYSx8MgCs7s0lCZJUhy1KhF6D7sOvGVcSw8Qod0NmkwOpXU+CElIqJS6CW4pnMyeMseRE01
wdfCcClmtzZL/hMGxevo8/3SEbpeeXNtzfBfZSXzQv4sFT+6eAVbIiVxbfV7lqr3yCL0tIiOZKtV
uXu0GCFKr4BHQjECCb7+pJzIh51DM3mTDXRWYdZK6xP0R0UVkhY1z01IPrY1ak6vEbcx8kwKpz+x
3pyMeB3M4OEiUBPNOxU0OvGbFSGmM0z6L+UzVuHTT9gb4wU27O82hI3AFd7LiwaHmeSvDzMCCduz
JEw5XXq4CxIE5KcNewc0CCfOqvFwbPQrtq4bru+31pekLeBH/KFFzD27sHq3+8R2R7ZX6f2nWhCU
Vifi5f/mXWmWZytex557NT0GE1RMcZ2E/4uhQJHQLP+hgyqzXTQ39w9hR092ONED8sJJfP24rgVl
IiMPITsdzghbeWR93uNwz/W1k9LceFc2ZCSBx3Zkg5Xxia4DukbzbLPJ7Or+iy1Axo0qA0fd4qad
8gEPwJoEyGy+5/ENpAQixyzp4wAf/VnpueXEfma1xmsRFG4/4j7NTa1GpI8AcvnFv5FAr104JGo0
QIYBu2rsxqGh1pMqSGKEej4lKUvBY0+DYtRiYfOO6Mjncwwf6nh7tnzylOwQTmHJ/MKBG2uMRvKd
8UxoKyzDx6cYAfDQM4r/fMxAX/KDFMNbWO+E6SIPL112ywcoxaFheaqyxSxPjmTY95QtS+U5Z3+n
BySXWoxslkW75meUh42Kwm6R3O4TEkRhAbvJIBC2mvkWItGGVOaY9c/wjdbPq8iTYhk1wMXHq0lD
lT9K0MBvMce7tv4FsR0A0MyUnbqSdD6NOM2OQACmFLb4WmKa0n11/YJxi9qRiseJkX3banSyE8W5
QhLfk/Wrhh2Rjrf7r5+I8MjYgOKyObWtm1gPrkUmMvPUl00c5jlnuajoOLUGNXIzeDAAu4ZIHU7r
2/qXKOQZ5PJuCuYaM9U4ytFKAV29KRrbQLBDhbFMKVyJ7ugMjgSWYxZ48xXHyF4JpsbExwLOSsxz
8EYgZEDTcBg5nXctjjVeOqikM4dsGqqKO/HyGpt1afn2aOApTnoWpMF8z7PKcjv4RHdzNT2PjVp7
CYVTBu5Itqnu/8sGNMB5E7/mN9ygQaF3hHC2gdouZAvLQsVZWkHDtaLagvBjTs+ccw7jncb2tmB6
x1/gE8kBid8ludMz1Q/jsz1BNsy0T4D4iHl79fMKWAA3xGDNAXgrrbTlaj8DUDzMZFfXYUNU1Wog
eT65+KBYpw48fB+l6n1Fw5kL1Y98UIDlbuKYNkrs3VxlzrH3LW+Y1DdN3b5urqBB9lWi3lJ7mPRD
NZ9XM50VY7pi0i7Xbm6UUBWW4h/eqmCMlSRZy2Agi6/FBOR7TsloGPxqbeybHqc34Sa0X9ZkjcUY
7OiDQq8v5JFZXsOyIHLyitZgpnt2xY65mXFX0ZTXpxvaXifosGNdej88VxbUCuQoSrdE6CibX6xm
xImgO1j7xu4yCGIONF06N8OkhEj7FCu7Kcz95PGQxSF5aUV+6zZL43CLQDlCqM2FGGGMIdV1kfSI
XrWMFgD11pUmlrlqazhD6C+fOufTHNBRN6IBgJyc+ivIytsqPvn4C/S8wBqlYH/KY4IXBUkOb7dc
RAHQbhJwF828oph79W6Nr6F+DF8rWVHaoBopswo6/kn2Neix+Cfq+fOiGKfp4EfgtXeHR34bD72Z
VZZZzwOnT0kbn2TXnjfn0ugnM16BPOfZOF26YrQ+yzVgcBXt16PX+TpooirYINFy9/U2nLV8HL+i
ZWxYD61UcXLtEKoOKlhfYky2jUZ4zS3GU1xj+OM52yC68tK5wB87iefO5lI47bIJI/YR82q2laZ/
L8ocAJqtgiOjBFtpNXEL1axwIC2fofvkELN1kA8nDfYIE1oFyXWn31UHgjHKrwFUdfe8s7gghxgE
PrmU5V7eFAQXQJBn7G0NvWTLJ3uqfWC/B12v/fFG+2Ju3DXNn0+dj+Y8tNrUszav61y1F029pKJW
VZeGdhc8ElGwF0ioCzj87egkIKfTHgUcKtGyM5wJ4TIfMTSbrxI+bhOT5eb8n+T15bOR7dDTbSNj
6NnUztkaNrzyObCnS9Mn1XnsYUSlfj18IfZf6qF2fChgKbVEg1T70dybn1waI8Tm+YL6YOO5tfPb
9Cal5p3jrFRAcFIbLy8mgnD3qjuenkyC3fVnGFfpNB91WRZmK3tOKwVoVJXpuHDQAFTnABIoSvfM
qhULT/WygCG7MVuoKa43TfriaRiIgrqHRXIyXofrOFR4WN9UpbJV3FVzp/XWCYO1EGoX8nOSCVja
5tS8sCOp7LF9EWXTCfi047y3bs0P6zbTcyM7AdGzliLSCz8ioI6ZmgI9X+dTA8+8EoXQ/+QfzJof
B49B8lv63rMv8NwLfWJLW7xZiE6SXHY3XWFbGZqlojmJT54z5tp6QMJCBqvnSpiT0y28bAZjpVeE
5jmlCOe/7pWZMhHN1u5sMUUbh12biu9HXoMQ6JrjH5igmAnJlzPWn8cCjve2fcF4eXFfkbwOXAaC
vfUfH49qwuoKiXu3KB/h+uz1T0AtRajfR2/XlVMk3SJ6U24iBpH8pFrqRvKyC9nV6bpru7ALMY8R
Au5ny9GGeHaoK0n4MfI/qejmGBU94ua8eoRchLfA1+m42/thxtAsA1Gzg17juVnwnG/H6c5JcYiN
3VBxPVSuLbOURqOzpFSmKW7KE8DBn9HDB5iGJwgThxu6gqmX2k5JuX0LpX3FMA4HWKAVdGLOjuO2
LT36PeC7+zmAqMwKBfWjnT8BQWfsf0jMdmaDhxv/MZb5Szt05gtnCnI4bBjNWc3XCggFHvcspsiQ
ugMeyu2qtbx4/9Ju5H8xBVnrZS9m4AynB4uIW/5IoKsLD7SvVzEtI74lU4G6qe7lulFVCuJpTs8B
AI8/KIbTrw+6h6I6dAF58Qjb3HFa4fogZJGn0Sk4ex7/V7kToJQAOH6XdGCc/c7VVZWcn0Yb8LPq
nba5aq8hfAyVE/ZfLSlmox+8vFXzqyGTpQC2NFLnN3ohTwlXYqwvqyAEbHjHWZ1IT4V6ajzUxnXG
88YkI4na36h/b2BMXW33Ubw5SYQDyxoYlyDJ9GaoCeJlrLmgZVQ66dbg98A+Dc/Q0p/o+FAusPLI
lcVojAV7GLMVZCjhXtHi/HioGIIs2GvYLP8XtCuRwrId/cOcXzNySCYw8Wv4StIRyy4l7YXss9ue
6seG9nL4Lb72ooS/3yPLVYNN+HsI0cXlCzgtgHHXRbnhdqCuzU51W8siFbPVrNQ/paLIq74HSPYZ
yxvE9LcrbV9MAAyaURqPfkGaXL2Jsn4RtfkDXhFMDZabsMiU2DsvqnC2M653qhMlnXnwkayzEzSz
lJC3isDnqRHVMllxk28P2N2XcrmQFaTpw5Ka38+FNnb3unNzFYMkUEO0snUd9d93ufzwrso82i2f
Qhk79Y4oroJ5I+tSb/HqEBHdyE+uAXHfoeB891UNlcBpcYkdskunJw1TdFv7Q77+yNlflurdIAks
Ri9JZWN1haVZolasgokcuq58gYjAHQ7Cxr2HCKIZUiBeG24/No5HNrecFSS5YGSfi+SFK3bSSBKy
YIY8PxiIGwZn0AIauuQ7UkRJCZdOEQXtwa9Q+w4SgxIkxB4s+U2lb1UWhh+eC+Vr8xXEKxBkZV1p
N2huaidC/afe9ug7ywxsdIHbX3mPE4M1iW8tzvk7LmKF6OBckvxp2T1uXZdzKCCAWnco72mVEpOL
DK2iY5YVWoBeWFshNbgVzjfIA3xYyHdX1M43lTFyfAAYjAa+HenXg7OxRPwuPwRlKHc5ASZL1TUL
xIjDd+GCtGnJYTPXXCMWEiiN5LjJZyDxbxArTixLHgRPfGhC73NOF5ponXAsBcl3yWmDMyoOMHY5
ors9MHhxXgE91zPPLgOHwrkzJB98bIr8YX/lKQwj7CVnG39FkEkuREyTQv9dxO1MznQzkZlrh85L
vg5C0sjIZZ6UoHzNWuonmEH7QAevkcASrj08f2CXShCIUmw6/ruNNJriwGY+smKUlg6tzyBxbj9X
v9JmN0QgVbI5rT1mi5asb2QPTEOjsKfBsVBTDRlHQb88FgB3a7/Y0a5TsimSJjSJPfYb3saT4hWH
DWjN+ggQI2tpIOV/iE27AtMfncj8roqleMgrVpwgifdJq2fQ1FEv4vFFkqFBh5B4yFqqRJG4pS+D
k1qcCu74EtPx5p+BQqOwzLrwb5ZAsUhEIP3A6x8jvTsIxvgUuF2ZzIlKunvkzURF/ltGmSWLPz6S
iYKgorf4IBZ15a4xVnVcDb8SlgG7fzbxOOwINDbFB5bEwzaklWzxdDqrXOm8//tliIpRv87lvrZk
pOr3pWRRWbiqM8xufB9IskvaTwgi4fRG+0N6RBAlMMImbwQyHgbHoVHv1Mtn98sKWX5jtQYJYD/0
LeGAdodxv+qVO6uhaDeQ6brDRq8XhUMwg9ilWb/0WdBuOHcc6Kcwmz1l8aa429RlXEqKmlhKy6OD
m7p8wb3yKU/ndlb4GsjEzUBOhTcKdOIjJSrTNMr/K5v7fP3BMbnueGpZrjTyI+/ytl/289FFtM1w
Mg6dO6j8xU5TaQPV9CKt6ZG0LJIe9yaRFfIX9ysZgFqeOQmIaRfCFIOMzCWNeOK0iskAJZxo7+H5
5r3Eiu86Qlr8BMdwVsQPeEnaJkFHuhkEf6zqMOnH/ZqsgD/4pVoCca/peeEyBF5N4kVQV8RTlYAC
nyWb6wBIVz5ljiWcMi00Qa+dbVwuGabncU2yFQNI2Wild/lNOKqba6r4SVck816ITGxUdZ6RiJUn
LEKbRZq+XKv6Yn6cFmT+JmYxqtc/qWC1uiX+ILCNLiPhKGUunlQwRd2/s/z45hzEgsiuKMq4IAbT
rs+UD7FsLpK9DpmGf1afRa84qaVP03NC0frYS8pXt0Zo9aZ4qY8/wnRbuiwsbTAam4rulMNNUXqa
cBOk0y43yn8asPecsu/sKhOVSw8GONfJgbwPPczQ7oeceEbs4RF0cRaIavNSqAUZ55XgCjMTij2b
iuPvtGokuh0wCWSxvEapLGSTcFPeV03k9zqaYhFmB1DQTOjS9ioxWDIdY8CU3BBIycda/xRNxwhi
PbEYv3c+vuFJrTj2PM4xwvaE+wXJFRLrHjgUTQfH7U7bwsXwIBSgI1vx1U5nzryt6ZSlspEJeW5Y
SA4Q0mAJQhD35jXwS8iYOOS/jgva61ZKSXl02jBNIz7/JiiEt1k0ME6bkm2AcI/pZ2daviTP5wjh
F0CUA6d+r4Yz2B9rytrv3tfnyr6fOsEccg/h/PD2CcCoJ9c46vUqsZY4eVBytTwXjoJQTY+DB2QP
sEWQRX0PfmJ5SeWyHlv4ZPlvVHIdDsN6LVXD/PpCfgzA1198Snh3XXKVwS6tpzTbrsf3u1ZtJrU6
fjE8v6xgCzBKDO2wZFuGFYJ8GCHN1/8DhG9iTrs16N10Zs2JEPNNTWkzRyNYRZi13o2J8vA6XpAc
E6EMyHgZ+FqSE3oDtbLyRPx/NWQbZKzp7mczQxkjCWm1qD7a6qH/JT9FjC9zWd74/Tw4WDqc34AE
Yy439my7LtTkExJk2d3VJ2GFgX6DK9p4M4B/N+alxOcYKFMznzRTmI4v6n3mh7tnZy5QyULaz5Eg
q5D2S0DuIRGQvPkStKnNZgK1j3LZdrWN+IUwAdufrI/lFM55H7ntES7QzbSt00C0KgWtnmq2WqFd
OpdF7JBVcs+iBENW7hWmTu41oUFdKJvkMt9LrqUwig33wvC6DPEVNdMftOzAVkHn9bdZAMrYsOM9
ekN8cBD1Onkp8AYA/V8RyAIvjrYp95O3z2yTrhm0zjEdc5GTS4Eh5eMlAXdG4Tfuz0A1teR7vrdb
ZjCHoRCB/zZLKROxoDcXDOjV+g3JisaV0Sx7gCwEk2ZTsYiNbzU6QjE2RiuHOKioNu+2nRt+0Pet
DANdfvRo0/Xrxzg8w+ckTjgwSL7NsoPBuEuw4sogGG3rv6TEgy+099WF/igrtbgJSFhybt71O87u
/42+5teolR+HqE8WKnxsdA6wZm/dx3ZV9dQuocLDvAPRVfvuTIRnQtU14spw89z0q7XFukH7VIZr
LSqerv1DXSZwdzhW8Xxz9T93XI9feAiKtIoCG8KBVhe0nZ5eZzCklbYpomq1IkljvQ4ykIq5Qgqg
c9FFvjK/ix8lG/Q/6gOOib3/MQR4y5zj0q8zvxIk+0ILyCNkH0MUUA9UFKDRyUnlOU8UVVeR3XLN
FMSpP/MOkclyJl5QajWGkBpBKE7lFWRmKhgVBs7oIXHktk+sJnJW2T4Yrq7U3+K1S5ES/YaCaTNT
L3oJi15ZbAXPPzGhblUoS3h9hSKXI+xj+kzkOJxL7cpDNYVgqfto8LgTstbsLk2Nz5TvC4ObFEm3
2nUID/M9O5OmTFkP3/4h4knrfn49YGPWpY1RWKZBPFdLoczv1kfM/9OVT7+u+5CJ44ALGxtXKCG0
KZRirQI90Xrjf8PTB1fjeMvruMtWX4QQERdCiDE9d6ROgAhyfcigvf+pZPbisNbifLm9e59doclW
Xurz11ignhMIsiAyEJuC0yJR7+6A+mD6JMXej6IWxe4nTqP3Uz6sEF5GQ9DEK2AFt8Fqc4bYvrYA
whsTxfBEU+4xYTbZuyjYRf9ON0Ta8RedsDFDvLnaIJEYXAkDUu15ZGXigamMavzoNvDxblsB5LPb
+gZhKJFzV71gp6pVAj3ribgsgBx2ZRmvqHcEijoWrq6Qs+jVePLkf8wAJiFaQKDnQdSthi9WSQjj
1eMDCy7DRwtWm0D1pvGl7KTxtnz9DpnvlxAQ6DMx1MZrQgaP8uwVXTDZHanavvm1Fp+xIMOkrzEP
IRhT8nGwhwpqzjbAM6rzjy2aQXNK6qNe+wJl/K01c7mxWG3JHup/46ZUHEqQ7g1lRaP24/6QSAJH
4/lYo6aDF8l93M5DElcG543B02/K9DDa1pOgaZPnW/URNar2EFiVkKyzDQs+msifc9zev8hi3Qkw
ii7aR3ssmnYnEAOOUc7wqFcACE+urRCY/+1euxHA6nHAX/yQXFGiuLJH/bdzj2O/Qb8EYqv8mma+
/9Ys4gjObN948Q41n72liWyNzpTSO14kNH1Wd7X7oeL4+bbV/Uwi43aXUhBn3d1rYIrZqpsqfpMW
pU+J2P6vTbCCqb6aPVnaxk4kQgI/bFL2uUZkrSReUbhkbmkZoZ5tL8A4bY7qNe2an+T9PAwuB3lH
GpZrSaQh0edLmxohh43SLuj124Migi7ljdku/ezTxthZT0wzju7W0pQ6kFWExfG5sAp4sPUk6a24
cm/utZSrv2UhZvNcLJLvljV4skdWUTeJ9+RATneuR7D7VYXtJTmWxPswnAm7lQ9izVNeJGq87JZ8
+kUNn0Ef5h8a1wYvjeOvw/sF0szQwmTgPsLi3xz4mrn0ud4Oay7WXG/G5WYCfgjxtomkAw80aU9W
EIJrkaNvHAEHKvUHaQyNxAu2iBZvRJBaE/Mh8MIP4DR5DLpzVF5Fpw2ApMi1M/CJVCyS+49P8oC/
b4YniL1281p+p9VCXa890ohjgj2agu3wol09H3u2C/o23zPoLWk7dJYBU62fIGuHPDJnKxCoqJMH
I5sQdrT5QdEezl/7B4W6MZq25lVm8nLD42iK5V0WyiT/DCG6tmSpBzsicFmpiATqP5hefTsNAO23
378FALtombGYvSozrkbwBrtANdobIhdFaSh6aveVJSIomg0jrV631GIQo4vmmZtuHW630BlrCHbB
D8GU980kR2tmn8mAvJZk40mRWT+DLeweBG5n18MiJ7MLHFR9hBkZApa1fnKU6XYTQXdNggvxJBAT
QE16OfFAsUe2T1KqYW8tqrlS3Nu8ZLtacEBtgLJtlvXOcXdSQeV42Wo1hCQG1KcKt5KF3zGjzWTb
3cgqyVLX5+S+ej2/s9gQSIS9UBN9JrkOscikwn65en+RJyOTgfKm0/zflD3hmHyuOyHFAeDOXXYv
CRaq++9SNK7IXJk2kULsM5JiFDyoqsw7rnkIexrJJAo9ZAUrLs55cborvDhX0+3cSjwfU5BIc5QT
Bva5p2d785Aq2Ns20uewiBbiqPge3YSa1gvRjokUFzxHWxNk10xgEWYBK4C+MXgjTa6MaokOppPG
4DU+xOO3Bi3l3z1y2loLrAHPdPdVGw/38mRnjEU0k0qDZ14js+rTpkAQBDghf2BlmNFRN9BX77LU
1UuHFQtvKvOgvV2kYdptVCbb5nGznegEpuejlpng314e+rxHK+crY/c0s3Vk8TAGLVCTmNhYqAnN
C5XdbKf7dpeIevL1HhoovIXOetP/MB4eqRghDSmTg3KOJDCm/eTz8Hr1Uiz4kuYPgOOfmGkcsO4p
I57YZJHckQvWQ7DjDP31Eu/JdZjpo/sN7OVKMf9ms86HPJd/0j/sTWMD2TOBNH1gcLbHora4pzqE
zs4iBdOKeFYBbglIYf3tbfWlYkUdXWFUWvY7znl2ZQ93Lu+0aJhXtTNbnidpkWXkUCngYqiKFbpo
PszVXoVvALjKjxpWJhhTLcgzj0+AoBbfghdUPi4nGavNPiR+dinMHbaFdkePaDRFkMQW1wAkAalX
d8OyHr8KcxwRzcP3R+NcvWjFTUJbLdSL7x89Qq9Mio92hhJVb2ypDGrvXtoC8gNGVtKo024Ak3Ah
POE7YiGsSCQQdigrkgCwyGycRz3CnjG2y6n+aCVp7Z78q1inx2EybAu05PgcSDXnK9iRC9AfnU+n
jDoSfOKWHChVWypIvaq1jSNiedUeRMemeKw7AYNAKUayWc3EjoPbjh61zOWb/xv2/zk9gIwFVLYR
QZASzYD0XYMp2spMk1ovymNtEj/a0rlZDQYrAoZpHw82gP1oDU8arKLw+Mo8zCaAzr0fNUDfa/lL
JKcv8tRLkFatiBbN2JdkUsn5qGZnfOF7Nj+w0Pa+9yHUwitfEXvFAmFzH1hPJlb4Dxw+xYnbqAiS
4CRN0XeqGHOaorItucSk2QxldavzZ6l1vPUYoEo8ReOLh3vcJDw5M2aRhZTm7GuOS9ZOHMjFXbmd
XVUFow+WQRuikQUpkgSYjzcDrMd3qNUGaKqoC0GJ00rY8oy2U0kGid2BZBA+cb6/uxwutcD36nrX
EyckW1hWeLq0S25cLVLpRTc+RWqA3E/bsd672qMdJUGlWDjUubT941N0ukhkEf5zHmdxQwLkWAXu
3KDLXZO3ycugFooP86YcSIRzTWADGuA7OJy/XcccRX/HoE1w6yPqCasBzToPpRLaQGXSw9aYBc7D
5/VTqBCT0Lb9woM5iYhDdDFc3FjaxiuUf3lbJ9hAleZuKlG4CUQuOqSkr1XIZoOS+0p518zLmRp0
CPAJmk0nJ5okBOWTc2ALapziRGNuQbUDRuILY2cmGv3fueGOy8ykrvPtTicjbdGqUe6ON8KLKNyA
KUzluz2dUPJ2AeUinJeYzb5ZHT5+n3FuA5DEBxTlj1bL8TKsN68Z1+gXE/zEvd3y0Bn567XTa5hy
szYSuqflCJiM/EoaJDqluDoP0v8hU1lyzvWniBYih45NXGeH/oowhAo76s9HxxcoiurcYzgXYOZz
7tjLC5mxFpWW3tSAkelxfWCUCXpygd/08oEZGeSdjC13W9KpEg9rs+4JDcmKb32O1QUcXjRgeekJ
XTEDFZy1e8bqQKsCdYXnmn71RHQWfD3g44q1959nhQa0C5ma6ZqhvnUtudzSkTxDNdBIY1toKafk
O2laih9/oPqFUyH7tSaXYtl4Lrl1g86aQSxWTi4K2N3CcUgs6uMI+7AGu2UxBBCOnngvEX2sx+xY
iUl+BRCFdLPOHdsDHd5nMrHLyUixvdHW8KeTJZZ3fZrXGaIHQPDfkXA4wHVW1OH8wnj+SkJ8mHi9
OGM02FJpkFHK85igVW325XuM5SPpwCryms0IO1NvhBZuQaqmtwk3RQlsNZjMP/L9BBrpXlytCq9j
jrMhFHfItSBB5PhOIs+uRe6c/DrcygEzN4qTNrV1loze6j6GsqYZej686OukFqIc7qq8OcC8zMAF
oyb2e2xOq6zEj1mKFButZiDU5ZPTzdnVMLVWVA2EFD0xIP8vjO+Qmv/cCfko34EJ5sVjSX2x694R
JoGnvEghtFDhrMDjw2z6Cce9uoC3lIJEj7drOwQlDp2E7y1ifvgZmwz+iaRbAgwybL3SLGcP7RPM
lgI2gjyX6nPgP4kcLYSNsCCJ1IQjV1GGWoTq5lOgu0n4JmELloJUopBgNHMH2Tn1QgbV5x0OA3tF
aylRL6zt4dqNtBQNTeYMzEh1faDfIiKAHz/P3yMCgAdjhU7mSc7GLKqJD/4QkrKcnOb749WTgdVc
m31LQhQQf316uXS5064QOb0VyPcpmD77/PxwNEQk5Ix5Kz4pf8c/t1ISQ725DLBjS8bpg27egIei
rvDW7QrKjX8J4cDOjiqnUVgFzQoMxq/DXD8cWGOSmGSexx2k8Nc70hqeacDRbSTo8aMFWbPabi++
6v1XoF0TXyMYsCSE1AWApGfT3QweR5jBU3lk7PksteLoUMWS0YNOSpH9EkPv/4Qu8DXY/aXqvVL4
AN6K7DBeKYDgwW45qYmeQ62Ea1RhOEXp75QCo9HdN/0wusw8X6qg5NtuwZn53u5byMk0iml+DDAK
UPT1Ax5KH81FCkJ94rz/bZgStDDB+MNo4Z7Ye0V4zZqGxBBY0rQ6RhXqOWeT8h1zM7zHvnetWtXK
WYyXDG2+BL7gLPI5rPXWceK4QQJVQyIV9rXGX7In2eUsWhNFJ5KjLeOEzY0bcNArfIyGDILdJPuO
BrcZ3kE3aTZVmEfYnErD3f9HWSztf8W0+ejGUVHP/C3bB6ubqxKmf0bnD+Ju1ZD6jTRiM3ejQ2qq
bsDAP4t3WWTYQ4cKQ0+Qrzeu7tIbzdMa+rQLzsnD6Ny6zQV9G/Gav2B4F7vXrG8454Zd2atBoY/W
YwDceMckoe5jgE1lalBNsUb8Pw1vKpmI7v01b4W8ifkSMwxNCgf9+BZP6WqM0feODvCaOM10+r2K
jrKf/gm7PlsKmdL8JWU9ywUCHre5RNhPeS7QZojaTfibmOr0sGxNOyhYRLO2yDZTXlyoIX/FYk7w
7YKmYLXswo3bHzZUc/4cIFHIe7O8D5ZJwHfB5+cmEz0rxNVR+zeQm4Iu5c7OjJmXtj5KXoCZ4mz4
4+V9NdW1vJEuGr1lczfxEFPLZ9ZRiSKJ+XM60HfhAXXqgMdkz1he+gvSXuHdcc6WIEDVFPqaLqjS
iPmybDUvDeEShc06ymmKY6tT67pRWcGcSXRI8yWqgYhMXOCH15Zs0wqOd+nIh6XE+SbBruML9iIR
PX2jCpPAWFxd1YLURtGWYigzM/28+5+sGHgW/AUx3fts55G2STf4w/ydEQOI1DxAROhRU5uZP5cT
P09gWVE1rm8sqjImN7Mqap84wx2tVo7jSCqYoe/gojHXxCOgvKc2Vx3SRQuNhNtNHdYomQNcgFeR
xpCbDCszTLoBHw9/CM/qkV276DCXsVb8nGAZslzueMl7hykvYRQDsplx8ZBhTghGXKY2c6ePJ29+
QrwVJqPG0eQjjWLI0CUolG9hJMPIROLPQBSb8R6Hy9AT8SNgbre2vsmmHuUknHmpZuJcYti2vkl4
XF3EeS48s0sQVn7h6H9rJDxdPzv8juiKAnNQLQHJG7VMGm9S8c1UPUCVkug5+6yMG7Hwc9OungJ7
RpN1Zt2kT8knhL1n3qSNkxSYuao7dpQPJe/HgRB9avtLggkKgzmmFdVgnvu38hEHAxgfzxvFAIGB
oVHSZnkWG0j+yl8JE+/FzChG6N4Zjxghdp6dnM9vB4LmAGWOR3ZNfGTXn385NlFnnLq8+54uvIHU
iaF2v8IEA5CNIEej5j1jY7hKLfV7HiWFMdvlMjtnmIJpFk7DGkjJW1ipD2HsNIQWb832iOfgwVol
YuDRXHXJkIN5BuPf6gVITtS24slRtaKkFpT5gODs5rjm42arSexOJ503dO1oUxkgHS+0isu/NTVi
USMNryZpCiWTR38nj5XB4bqN4/QG89rpZORDaxw1/8JLbuu6pSww9d9WCTj8DZOKfW4Sbiw82BR8
mLCzctRBTms7Kb0JAEM9pWWQitPme4VJZnkNj/qJmOzs3O0OL8bL6ggUVJv3quhYbn2Hk3EzqfiT
CHt7Nt7HlMuRhzPFHp2PZM+lLkLvHaAgscmo66npv4xcqWN9v/RcsaVrcTIGDALdyxz49eBr6su7
ZwRwVgt5sPYTxyNLM+7ADJ/QLoyQX2WT/YF0XyzF8ViCi0vmV52RWc1RAPtRPuesFbWspZtpmSgo
lLWNHWU6wEY+BodDCvVvuhj2m1qsiWVmmw5quJC3wTklG9mXkSngKwZFLuZfAq7H5ep0PYFggHtz
txKVuaYRMc4KJgqXOSUZ4nEqoTc5JIxcqjCSwoQRn5SfByB+v5Ht9iFDEBo34lqwxnWVa47rvluu
7Ln1YDWDiatoKMbndn/UFOa6ynxGTVsomMRLdddPGvs+whYBfKq1Y5GT8/+9+TVBOojLEdolpfMZ
+3YD00nU3ZMZiD/Y60y/qFw8Tg7261OcM8CxLwh+gckW9VPOG8hFPTztSA3UOfs0xAAC/aTLrxA2
V9kCn1GinpSyeL5JZjem6sUCy96LlKSI9oBtz8Y51HEKWpRnMGM3PZYyxeIU7RB0MBcbQ36glIzI
pMvSTb/e37qwfXyQ+F/GqMmRyj0PpylDDCYaVtQAkyyBwEPRWvxkJDHGgFiwGWtplkDOaYgzGVKZ
Pa3a2rTjfhNonI0y0eog5YtOPP/zR+gMpgKUVAziNFggq58Xw4uOoRmSchfB/cGbyuXdgLwLKqXf
WTtnp2Kv1InxLNhI5V2YkalPGjP9lcT6nyS8ZOPTBTJcaN2YCA5d+s9/WRgkMQsHF/dxtGeUBV5I
fl9u9qualLjAoj3y3y3Ktb950LtSSIMx/R+bhMXpxx4tIOs5pkE0ogohgTEgD5lTouCE1u90u0IM
1BE0z3jVKBT+4gVwJpyJkoxdQFKvQKc76GlI+m5tCAYuuqfmmm8yS46Sk1i/nc0JfohNUqEGNq4s
gH6F/pymCGEzKPgVzCZdBBdwkkNk/wtOKUAPX4lAp1xBeQG3OIlqpF+p8yTfbEPFOdkUTPTH9VMN
bKcHj1S8NnUvYdYHwSejH9z5i6ElrrBhrhVf/Zs+Mkc12HTY2JthZP0cr+qzAfe7+DNz34bOOLRh
9D3XHoH3FVq68pytEXaIib9apgc74VqFGSfwWxZzyeCHa7FwIfHoN6ap04erb0X/f7jjolM3AZbK
2jGbagbr1t+pJFB/ZiC5JiF/H5umlpgsvjFzUihUGoNoOw2M6f1G8atG6OyD+F8lRokP01Nn4tgy
JnZC5FEO85BvpinjdcSZbE1vOpVHX0nt7QhcT206Ih/slGT/I6yxZ1ZZcwiEGcnb84Fj5ElXqdHy
wHsnCQ+fSO9rbullj4M8RKjJZwx/d2Mm23Vj2gzPM8mn3KHupTZIXT/ok4d8CnIJDRWw9mMbm6tO
3nuYhJOYGEIOgTCgj1I8h1PPql/JWEG0u6qW4GULEz4x2fneituAnwJGcS1xv7aEhT2JoX24bMj3
Vy/Ndenbs3eMslVmdrKPiaoxsfQ2+h++chX0vPoGxn51gYtEX2dq+1Ei4i3GXy7P2mXvTssAR4R4
EfXyDNLcXKF9qF1NW/kY04JHiqNMM5ytQMdCU1Ip1aeA7Q7mm6HBG+hClgvftyTB+CcVIlyuMTmt
y9GQPLcQSZiFYaXWOYUYtRb9nyVJgpBTkKiZU+ExoVcadk9jMPo1TaH/KIRuhOxFWW1ub5DQ+Pc9
Utz7oawQxLZUCHUmP8DygcMmvKqQOyLCwRrYZ9A0swYxbOwr/4yqurFrl5oGXVfO5UVtgNqK+6eu
RvYabmM60onH1QiwcLjTnBpFAGQx213To6exwdUT7iyPzcpFuxU+55ESAOXFFrjFRhgqn9tnFnv/
3W/YxJQqWoD4UX3lF94ocFKmJeBreY+CzB8+naKayZ6M4LNVriBCHtfpAcKiiZ5uZwKWeGndSoFZ
dA+dSnJkFXE6+0sP7+xG7CxLaQ6dVX4MwcqNHU/3xjl2nKQwpt95slQ1Uj5XK8yD+G6C3vxgyJto
pLPOnZAwaF2yPl14Gk5YFQvYBHLd9gSh+jVFKf/dWk7a6PW3VwUjnj9LoLvOkxa7JHpPsI5i2+aw
jdPYQ2tKTNtwrLQC2xKC83JCyRInIVCZvGyRQ05eHhka+KUk2MDoQzcUEW7BbV2jCx9C7dpKN54Z
X+Z+u+A9LkEDc60Jmp1Q33fzT/qZ3Ty2kdJtlUQ3hhBwXBYrpJYdy9E8L4TTJi8M9wyilXnAzgMb
jle8wz+7b9U1xaeSkV8q65S9iYZcki4pFJ4gFXRmCpCHzvX6A4cWUl8Di5QSrdIE1UnJ7jlOSatA
MJUtTL4LbGQQiy+GKeJAEd4YN6r2346jJTdqkcau2PbQbjeNBwlJ8rlVkYjzPF2Sw14qIWpOHuu1
hxIqQbuqLyxu2dl4T0h8smpD9GK7gz2i97FMQ2qv/85XE+A2VgAQ1x4TnsszaKaeE5bs4dOuXGu5
eTqXN0jyXcQOTSSDPvgJE6xu/04ekQocgJEImVPe0nvsRoAjjzi2E5JQTxRkITV26h6Zbp3zM+Eq
SVo+Pmc1RldtxYpwkztH+K3WSbKntQU2mxJfVzkqnAZ7jjYjubcLMoiUQh0TpCiGz2Xt8Zo91QUy
Oi3mdrsdAy5RiLN9R2OWjUMy9sVLw3iiGRhzfBcsWn/L0mKtz8Qzqt0mwPkwjERQ7RI3Sf8iS440
NHlOS9rS+vO8NVmoSMoEg88rT/fpDD3T3fz3eftqF7aToClniIfc7SBOjwXI+kVT4OjbKzrb71GC
LkKNN0kBTfqql72KcENsaVcwBpShuW/XaLjB8Uz77mlMkzfq7oSRoXwkbLuKmSZPM5nhw9YalsSA
P54U8W4Nd0FQSgXB1e8a5G7JeJVTWoSAw0UC2UpiMpgpSa2vxSH9FIVsMd8uMnqlOk/EGtR0NTrG
fo5XfSvEjwiAZGUARHQI5nSoeXeryMCQn0hnVaTfk1Lm2b7P+tSfjQPG1FaD4muvXBVrcjNmacnn
qLO8U4J3nDfrAmtzy/TD7+Y1lNhzVtTnBjmRrQ44FwN52vOjSiuJ4gS1HxMf97k6GQFT7Ma0Eqw3
QUkk4DSaivCwoN3bq4117QNbPgtV8PK7QTT40d+ozfKcDwmg1J9qKdyJ7yjTXrvp1wsHFcvOw3Zv
tO1Y2ArnpXBO++DygoHTXiVTeDMsvkcmuwPMDKlfeHiWGPbbXCtulZbhfueSdqKs3z7HqXg4jaP9
9OyGU8QM4JkbYH5D6lz+o2Pxdl1/1n/XRM+i5hIIM3ZEb4REjAX5COkS6Werr4Ffq5NQKVgeNBAn
/MxENxmDxaCTDaAdIr1RjkbOvBGzGVfm7MkUAxT53Ot4vVWg3BqxD3ZBFUfvVsLxKuEbht2L1/dY
W6s4MunSsM32dy/V/4y3x/5rHvlVki3uE0dTLL3SQ48pYpDk6IIK7c611nC9hyqxTBfWsIv2pmRN
JFQVxuRrtVecpO8psXQsjZcTQrrZuyo5lKNG20TqZAa9NcpgOUEKMgFPR+cUoYYLpDU9hs6qObza
M3QKfyMbetSpd8SJmYAZ+B0i3AsUgX9klKeDYNMWyj9P1O5EqsR76MYHBF7iEfuyy8c7CjolNx7P
kpYThil4ZLjAB/A4Cm/CUhuhp40/pVJFFzvmU12oRxlT0sMP8lN0VBkchSLm7/OC9Zoe1mUVq3/j
Pw4QubDgd5D2TH4iL7IziuReIJIMvjpnQ6d8E/xRPPJ3UFFiU5sIQRmlE7zuQtwBORPVpMWflxAw
Hwco89WffLUogOFdb4FbQYZv61yGoQPIVtjo5+XkpYh6ZjqGWyuf5HMy9jSEhk97mGCLFTj6Cd9P
vzC2hIL4NI2eT7VLaGd1wZDvzmMI5hikmSykdrEdYQnHFY59UyI/hz80sOgI8UnAW0DoKz927xgS
5kJmGbFZOr3NazrNFH9rSB+632UTURTKQAiGHRKsaduxErfv2IqeKDXPXLpqvIb4//U5HPuCZVSc
TtgMmRoDoS95iRKFN5iDobEWDGNUePHTBIO13OmFYajAWlvOh/4ubceH/yiMqRb05nzfoEAsiHwU
8OdIZect4+sRGfCpa/KRRme7MYIeA1xih71UlHoB9CxuKMWstW/6yVE5FMpAAJF39CCt5rjZ3Gwp
xtrwvNGVu0NBwjhuVYtxGE4pAfF+WIHLnANKLLGf739V5JkkuRS2CAHoLDUn4mCvL2JTUtosKAaT
KtUKk4MhUFvK5ivrqquW7Bmgqm8cNd51inBcXhJnSMJ/Olw4SBgGMTm+SBAe/e2jfBm8d5iwD9e/
YQSz6ATkJC3NzxNZbWrPjmQU+bH/Hk3zsOS+hrI8k3Vqon9PNkQ3OfXQyMesB1vEQ8CaSBHvHKMQ
tJvkPy3J0/lG73IdzQFkJ/7XVyRoHOnXb9IM/w6mQ1PmLHwWlZnXbgr3me8XyZUp4wA5jZWy5aut
0y+QgQCsIlnJDQ9DGpBPVAxZfr/SxgvvPU/PvDci03SOYhQmm/whU4sE0oB/z30RpdcafJnuvxsW
7mnqhO8f9XbQ0zbUqsQp3m/VSwZnBUgoHkf0qqp81m6TQ8+GrOSXcxCsRqZQSL+VbIl0HcP7t1/e
LQOJIhqGmdGWVcIXuhPJI5cEiBen1k19tjLmmPBB2faeU2W34x0Ga7KdMcZv3v0srYPKKGmZPsbi
HuFoQk8dnGS7oTg8k+yVOcMiyLxUjjmP/TzzOFX+bWO5bkzrP8nkiEeN0TvMQtaSfTmx4R7h/g7x
6sxHqzjkkZfBZV3dX33y7OVeV9JrS5KsGu0LigRJc7Pvcusf86VYQPYtO3C6CvzId8BdXMc9NTr3
O7QYppMyBYTGjzBMtDYvWE2N9aWzUssA+f4q3mgyWyooZw7OYjMeNT+3ntdUUCkPTKyc8yxTVTiE
x8MkrTZaspxp+ybc3VNLSRbuYOWlhYSk1VqjnuHUGPg+nr++NvRGzsdzFgnPLuyNq1X8rplCS6mk
mkfQdPXlTrvaPIpPjajwXhCo3bQidy74mHCP75KpB+z1KueLO8dHTCrzlkxdTj1f9VLcsgdI7GlI
ggnkTcbNgV6+6Yb8w/27RmH+7XT2EJKT5mimHgd6Ifiow3IYmeVYp4/U+0rhERYzMEG/mj4IA6Ab
Zwmdt8kbCmDkqBHy4FMBVxAZxuITk2YAkm3VIwObietlr0yyOx04mqJay+YJTEwgTDfVlgbSMZvT
5cJ91/P+MpKwDoarJ0Un77LK4xKjiW1W03o28/ntNiTA1vxKqs+wZRgO8Mab34ZEbyrPkMbUGJOU
J+AyDx15fj5k61ncIC/fl2ryXWTqGWt/mHgLNosto4QHD/l4NVcBFRBf2disgwUFQlSPi858Qze2
3sGf3cu0/PpLClOGaQZZJIiAtWydzv7OsgRIV0mW9KXeHGwjpWl1zX1G8AN4DOYTDi0oAUP4qOo0
AlYKgY7XLmzIVpgRBhHvf+2qCGKlLZoQcT+J7H+2Bj0SICMzmQyT0vZ42/sBqNOeEI6greIiuUiR
fOj+xvl/9k0GNL8ObS95cFdfU5Hl/ypn0Oi957m8xg/IWz0UDDFMFlLdGuWgIavjRpN8I2rU9Txm
HzoGEotQG15RBpQU1elpwO2BqgseTD3lCajIN9lyti/wzJcmgWcKdbo64j3K8QtVERJRZMMCXWAy
Pb3341kaYt/GtzTZsbSFaKM3jgEw1Z8FXoHabK/nMecMKjpk3zEgbV2Bl9bAJIqlbhZB98igYxy/
Xwv9PxX5UocAL2sjRR+pu15ZkD5ViowfjphIasV7L6jUgLhmMkQcyVjLGu8tDLN3KvDer+6SZZDi
I7lZhh0X63mYV5tWIMwSE39AEEt+euDcaiK2nxOP8K48rMFos0mm0CLpEXRUVFcH1N2P1OEZWann
K8t5mv7kWOYWJUEwdzuCbM2JZNOW5Z0+01cphGLV0t1eb57u03h8TWpG/iSDHFTYAa1YdIFPPBz5
z/cPqB/QmuZXKQ3s4fVZTTB9egoF2pVJA07GWYNwQanHIt4NyfSvbPgTUW/axPaSyDFst222cdf5
Yd49wbVMcqlEVl9/faTAzMTH7zS29kvkhSWwZV8DPamBmpnHiQTOILCwuQ8J6RbhOEiwBccZ5oAy
Nu4FN54IpbVT18FklqbB4FWD421C9an5CrAQmDBa7jhSrEAdL/AHMIAVNC80HxfcjVzKaPuu/mN7
k7SfQuBVj9sX4qRzR+Oc0JlIoz/qUVWnabXTa9wKTAZ9ymMOfE1QRDA1x2CKkcRMWzZMjzgEIvbu
fHF57lckHIEBuF4pd8kCvE317/PM/Mavs2hrZjoZaPVuolAGrMInJnvNQDl2el1En05vu9vPREkZ
ZBm48A691+Egx4PyTmdsGDs/n3UHtgAm/gTvE56Zg6Rn5HkQHH8c6yomCmblnJlNtw1G+2Ue1hpc
a+W+LFp/J7EyUy+G7P2i0gi0cCZ/X+NEJeTlDtE3qEoq7f+X44KGQ0du3nz2nmgZaMv+ikaENTCY
GKsdKzn0aNJ3Cq1FsttJ5aLjTL/m0g3cTNFhPwckvT6ddQ7N9A4lEtyNpzHpOYd/L+h73UYDacVf
bfncET0+QLUd6w4XUWZPVVHDr173s3iFo7Y7ilXdALVWV/cT95PsJeogXetPD++tpF3u8azitusG
+GXZEZeY5ZI6uqKOXEvGJnNg2zSJ8MhAIEdrqGzfa9nYuYIcByQyhRSy9LNAHfUUE1aj5t8r5+k6
spvXQOeLSEyOR2TxDHccpBI8j809lwXQ7xFopBOMsdiT4kU2wJ1Z1souB2BP6XPJoTyxaz5BHu+1
X6y3fhJRq6KJIlWAfX/NyJHooesSTIzqjFsazeWNWO0NbNIsOqTiD+f07jlLF8hM0gvPSJ99TwKj
klaUgtBPBftZe5laMvMD3rVoRS9MBD8c6dPOoDpUt+ZdxE/zbNypyVIRBSUG6SAcUq6BlmAuEcMD
+KJvtp8PilJO/wfpPgyV2u6+nLDMRKHlN/pBdeK33F0AS96K4Fl5exEDaG8E/Px1zNqsHhW+XWw1
/1yWd8EyCst9ZXNt9bcbVe1fblS51p/RED1zu1cC13c1CVBkbGl/ZOZBx/Jh+IAGw5r1rMSFU2Ka
gaQ5L2HnoJoNYSj35oLQUB+WgIa8xVsCdG/ikXJybpX9dlKSm9JTUVoE1L0uK4HHhrNcuzPrNeQz
5E+9ExIoaf/6kHg0EYEuuqwsHtWAlcBg25/DW7iQ1sZouAcxEwhpXRiVq9Vidck+WzDDsszTCh/C
FPrp306cKoPnOOCrzYMwvQqPjeSZIkEEDhW5q+01HKG5nQCWqCBjv0ODnqNAxaONnQqVvS6jI6dJ
vl4bVh7FhH5vbmJGyrTouKGjx4ebOO4/B8ofjM8NNQGCodA+1ZfaLwwTSU7U1kEyTkUL0L1UMdna
9hIsDC+JUFhWgdYCWQWIjfN8xPh3TOGMgWWRVLJKnrnE6rk6AGwobPcKHCYYzn8ryLZkdfZJnXA9
vy5aycRqTx2zJXZ14iKPud3jBa2L3ugfswA8GSAm1JD9d1zWhvcm0ISk9MARbjMFi6jsSh47gGoM
jS2Q7x+2FdT1pb2JJmUJWKaLvmQhp4ctI9ysTTK2F85VzsQraChc6hWsZqjL0bDjLmCJCXVAagK2
GWXWaIRjZFpiWMmkRGM01O5gOKocMZymh1z8PGPlg1j76YiLTVGDXoG9WCnoeU7Fyb5d2lvbV4Y2
QJtP3e3p7HmeZBTybTS03cFnfOfwg7RpCmV+xVZ5LEoC/MSynuRlB1PgAWuvJYzYr6btG+Kg7Ntd
QPgiu+xphYPbXLelVgI7QvV4f06zdmn2oBp/72PXU0ls21mBuvWVlULoZnEw4fFqOnD1Y9q3Ag9P
dOwPn32CnNlo4kUqcSg95zQAZHxwI+xafSP7lVaYwvBYZjKeWsUfI2fjAxCKmUYODtj2WlhO915q
zRs0G9f/3TSCk6EHIims/H9b25cW/Zsi2hRlSV6AW/IrEgv1CFT1boI4JCayoEw0ljEa36313qvq
9pKW/iCaWlnHqPJUoqQjtKGCwr16SBnFoizI/hNZGZ+NPzoSP4+gqJhtGDUB44cNZ0VbKEUnIIgp
shzPg820DkP6F9hST0heOCa4hj7PJW+Px+5Xu0vxUCiwHiCZvACDaTZ6bJDu9B7zRyWNqi+cy9Hz
fKDsyrWTf0/F7fURD83iLctQ/HyB2eaOh9K+RJ9cxEdVH2nBoIRTCrh1FGwb3uGA8DAhoqniRZ3P
LOCcTZzxYHBPpDSviRSwsmsXos9jDOw693KUbojCYpBIJxZXYEbAUMyw2XAU3UMLRtxfmrdPaAQp
M3cbdGwzF8UFfsMHcV6fLSBMEBRmoid2BQ76eA2TbWKZcknnbJw/5m22oqeVgluvhE7d7rINMO1F
0GV5vjnKsYyDulp7nEPCbyvr9vgbqic8tKVClJ9opKvOvkmg4PFabsrWUHrygR2MA9P4K0M2Vpxn
/7VcF3qkGnBCVuAHi3Z8wMC3M/yB1Vu7p6OzFngzU+mZSzG/Vhku+GC7RWrXuFdLbHh5C0Xm/o5/
BVQLq9CLjqy2UrbXUGyoUO1hllkZnd1FVK6Bwu4uKm3JrpUgVf4O/FRkIzFrc7UzpnSeGjFM6H8F
zASKQmjmgOoQGXtghrzmiwJcrZlMypj/2Fhutc8byqyMNTrwBrTmLVZW9U2HueQ6XXKxAgXrbrwd
efMsKFzEUnrasUnsSGfFu5o48vRhz5L9qAzkPge+i816U6ijGfT0BPmHwGchgvS2m5l5t0qVJQrL
mMROAQ+ngb2mh7536DTcGCe1qjrPcYKJAzQVzdLaNll6S2NNLcJqT/LLcnE/+VMXBK4WPaLGXhiW
/xnBvUEEONYc5JdJjFcyNS5ZNqQrvTMzp6BxV/8mR4+rXy5fouQEoZ23PPHrWw8HYxUwAWUfJErt
2JgH/uuwR6znTtV1rKdw07xhZKIkzx2dy0vuIIy1PeXV/iV0kheWDriZ1ogt+HvadWx9axhXQn+J
46LaZxc5YId9KTjr00qVsVUxVJYaucROcBHb8O7rDgWOyxtNXWZUsGWS2Z69yjMbQc+DS076WuyI
6dX36VZsvnBF52s1mFiSY1GSO2iHSOqrG+RW9x6xXS9gPDMl1jSrVVvT5NmQvcgQr7Ay763PbGVS
/fQx+YHr6WA2eIX70vPZm/sK4VtYEnzRhoFi9fQXP1hS5EUWahKaazhhcTcpGT0V8VhRiwaDW269
KBN4oDxVNWWEW0wAvWvyW54mw7M/gxjqo1cCQpCa6hLC5O3+h4BFnwp0sM1/7GSuVAj7vyIDl9vZ
K1nUGOl0/LIJeElRFOg+7P8uNUweKxOWWdxqLlM1+HZt3xpydEA8raFOwveRPIau0sQY89iqLUGI
GnNP7/mIM4Ep68SRTMKOkfLY4bQsciLTrRMkA+RJgGIRLETII5tj8M2qpY/LGUGSwHALQ7tXHTnB
AfrJlkl/2XWnW4WPJhfYlQL1zPI6mtDZrvYdjjbOJPi8vhqProtu5I0eJLnx6kShPml/d/lR9i6b
Eai/ZmhHKfrFirM4s7h8f49EJOyeUURB7yu6XMD7oWIHXpLRb6h1U8/zjqo7SOfeJn8RLIQMBpaY
ygaGPF1zptyYn1souqmgHa+i8ixEHzRmuGVD6sA6PbZK4oDLH+TzAfHs4uePZWWe+RhxU9IT+C61
B57sE1OagSYmg/+eRju/m18KYhmfkXKOCC8VFQn0t99+73gHB3R+xSFcFG1DYBJBkvdc7pED2wAb
4KnW9QE+Z4kk2Sdh4py5N1xAUS8UMnBztUhu1II70J3WulXTp45hTT5m1RQubcXIXvBL99q88cYp
pkMSNOZ21Pk6s8yq4IgcM/02jSW3QL0E9OYgxGaBeiLctUiKbmHDLQofiRBCxS80ru4vk5sWclfG
WKaD+UePJyWioqjzq3CWpWjGf2Kik/sm79+ZB7X7u7tY62yceHDtQYptubBCzmm3ANn0Ruzn8Vya
fcg1IScaZIVUeN4Lxbq4TthHDktBiiiIU3F5nPNaTYv0HsmHeW1evur0mMLDBYv+q9nlBnmPlU+E
ZryAu/6iDKAJWjrlYdtLs5YSAWt506/uCVQZMd8e9ugmfGHUiKKgAkfPka7SAQDSOVgbiF5QpC2E
Kf2gK+g7lQ2RPTT7dTEoSvrZweKUI0qTlwN3M+/ismeOVI6cTmBtXS6boC3t78xRRkiwEB2d6a+3
c0BvyfbC9yQsdh+FldOKzth7Xs93aX600MA4MM+sA2u9pABzV/OscPWPG4onZl4RY17eX0esTDyT
GczKGGMuDKA5Dqwgd82dPiDHva4DcXc6xk/TV4ggush6Hv1L4hTitLku9+AonuZx16YxTgQGVQKc
Nu6dQFqxs8bhcdEnalmCmmrS/PIV3mQViELQTeoc97JEXl3qk8CwUKR6o1DqGFoVpAjxzscSMVtI
MYcv7F0V8yySMla6CquEEQJtJyN2aFh/wC6DuFIb+i01mXSTEQZXFtARkD/0Q0t3KTdgGDsdI4A3
6YFwU2E/kGI4Zb38uRkSqm8ugdP74gk5WUhjZvpCmpYDWptS59FgE7+J14PNfokn5XlvioMSR4JX
yiRBF2kH2oEi4AYnf0IN70Y+heKio3MOqJrip1pUbh+Ruel2U0BOyhpdyqqrF/PDKBijlscEJsIv
iiOtOYIvV5657cc2TuqB+A0UgjcV5L6/sYPu4bQFrt8S/P3kp2nqtMZ/qD1JT2IOoJ5l47a91kbw
Mp1QONyErrzLoeR+ie6mP2tPW10MhWcF3DdlM+hlythKYQFER9WQ1JjCWCcyr+gMes+57fshhc7t
jlgzwkCsKzqCMw/gWQ+uc/Hid+s7SFq6gFxxKPrmZy4jBCMeYRdtUNMU9LCppUdqRRq2CtyK1AR0
YmDGaL48I0DIevGrvOclAlLSjuRApukFaPBlPXIfKuPC7Br+P0eZllES/ZfBF9y20ljYnN9S5WBs
iVnqDy7cG/QTd6rQckDJiVCq32TioB9U1yDT5zgbUJaKfn3LeyTozwKqjBTtgGHbJ1Qviu+NtJQN
Wx6h+WIyOHBX1H3UhdDjA/UTekSB+J1B6u5mcneZbuoW0cfeDn+mdVu1NpbzjmVRVy3qCGL7HHVF
kReEBAz5hlqlIu7qPpCkwdA5Ot+zEkXaityWcKTZXcNqMIZ1Xp73FZ4f2XWDCTYQYv5TotgWvt7U
dI+h6+cVecxSi8t5VFW7WXlqaxuPML19hFRoHz2cUQBwwat1cFS0fTP5XTyQDLh4Jmp4TLa9VtyA
Vhisk1zNhhKKkr7V4KTORiHCnQfak20WawwWmrKzy4JKc4SQsJ0MuiQOGhnY05xqxfq+zUCgav+b
z3xhCnRMxzA5W03zHmLLpwjawJ0F9zVuE9thPKdlseXr/PDcgabuduuHPKSGFAZD5QyQn2wxasii
Wpz0cDfUIOvfxu6konzRbI7iOYKs3dtKjSn3yNxYB4jcoF9T/KmST9y+WCVop/QeZCcVA6pmLwCq
LbvYVFvlTpTpJ5YgNALFvfsh1QCWrOdznNIz/+3xf0vbFbiuVEyovYPpPfB+y0pk6d5DjoaW6UuE
G4WLMUTB1HwVsIsV/1G928aQUb4kjxIODuGQt3gweliGjFccNh8WdLJRop7mCFumlzTNLwOK/GQw
P3ZmntxLvOOS0YnsOK7XCX3KF9OoeKGqq1NYb4LrbEXbmeWyuZYXfZermchnH11+EcdPdnWGiyyH
WtfFwlWgJL8Airy4wmzLCT76mzyh8SlFKzYNYYsQ6pN9u1j+alEW4I/xAcudbvIWf/mzQ8Qz76mQ
5XLe0dJ9IzYK6fEDLb1YsjpLt6XLadTJOueUq6jtFWYQ2MXhzgIHSl+tea2gfyieFrheRUjVFQ6O
+7k5uNvoOiTHFwjQF1LEOYuktdWu3WWnChxylkEwZWSpGNRG54PIIZD6D4gFDsCTVqgxNCZjJWvp
Dw8wTliwCOvWotgIuSesgCETKqGRL5zwp1bc//VO+B3bg+umd0xjrwtJwpAli5lmfGW+1GQugkKX
kHz6kIt6kP7uCWXTEwczMGpfrGt1hEX1+Q+Ij/gMY0/O2Pnhhvz37o5YEESpA1Fmj3Wo3XJ6hxJ1
SmctHnQSNXYtTL6X22PDgE8v+YiAvQUhpchdYQ4i3K+cr/D+R51qUdRlCTaUl7zsU+oiFa8f4oiy
2gN3RWnz2+xD12X2FSdfEwziaJJNdUIVZKsDZwk6KHodzjA//QXgIuDOf/i2CmyCJ7Jc0m8EWtc7
C21nEViflh2EVQ7i1jaFckxNEQjCfqrK8sKpUBa6KP3QeOQMAzLdD43s71JgqUZC59usQfyT80LY
1OcI0H5wXSjkYmGpJkAGSorVGtXCV87xJwg5UznEbYVAL3JaSVyE7SRzBVnC/Y8oI9ujyESKq9jV
n4KK2r5yebZ9++gCRZg+AcOeXgsnbYyupaXkszQp5xv15V17MczzUoHkcjiyLC/Jyqwps770rqSU
WojFsncCU/iZT1pOIfxuJ0kp+x0WKPAUHIyaaj0J03sSA643LRbQX+z9EVggEl5zakFW1mK23zKA
YB+yT+Ij7WKZOusuzbeox+thFvf4fV4XFGSh6grFkBcXwtmtKtkmj3mGCCT4Eb5Oz6L6A0jA9x5I
F/DXCvVBG0kg8ca5+z6bFbW6f8Ldgryeu9d4hk42TRCQftCBGvGGu0RpDY2TBAGvJdUA/n8j3kgu
bIn/d4kKkTYvIe0C9ZbBWZwzXfu+T30tDBHEd+XHt3t8uuStVKT9ZR3PISOAgorP+LPHx9ywL1Ew
F88I3fnQy04bCsEm+hFYQy+nKqnhCov54Q8XGCyOIHaXz08Us5Vq1+6uwxtp+/TJsXHD+0jxkKBP
bUKdIoeRSF2CenDvY4Vz+xJJX/5b4QtlHwMbakfx+qEhWbare5wHC0vE6+A80VOdptpqNUoZc5lD
KITjSQOWCRuJenPeM7qXCqG9mu0kEtzIGFG1eO4CkorOex22L5KYmYrctKvoV14lAVpo8WXi3Qf8
BnXt4QNr/BkMxwiw0CLl2q/pK0VyRtZ5OyiMB7PwcFuRoByO03fmHCzCQpMXb4Z7usOnIdE39r5Z
GReDlNycGyoiKH3TmiyQ4vORFxJ0UzqABXfIjHDFBiXdfOdDxLpMg/xSJg8EL5iDqAjl63mNl1aR
f1XyPah+PWvRPPDeJ+u/7nsnrnRNw1mr7xB6oFG/z+CCAjMVxMcUL53NvTh6eLCTG94IxxJz82Av
faTJ/lee6lgJYFpaq2DI11vCDbSxh2YC/UpQQY6sqdC/8Seh6Cluz+G6dOssOruSWVUt4PPrL1Yy
1k8/3rdqBgcO2Hv97AgcKMAgZr9lwzgG5f/KgQjb01BPpeThI184CyVGRYqqfMMKaZ6XBLPD08IW
zOt7bSckAUONa+69qr7dgymLmkiycqJd6AsKvBquO7EqnN7CCTf0GEy6mxhdMX3iy+qsu1qZrCEi
9DWfma95ykscWBQ3KgIJH99nIb6GqfRpC/ziiMacY6lmbfJgLeIzYIVu6MpoB7p8p9/zmLvc2Ovy
5kRQmb2tP9YnQ4nwV3/jYrBeXK4SBa3jHrNzkJ1cfbDJI10Gq/d7ncBr5nSBre1AkkdVeE6RyFN1
1cX5XND5LQHvsnPVfSUNZ5zlX9v9uURIaYp+yAug75g+LPQ6pDLNXEgWUltWC2esemEbk2EpVLM1
fJtMlSZJCNtUVNAX2AwcqzNzEkPSeBsrSlG8L4+T9ahYmdhUZzs7XRDbq0dXRQgsWE1zZ7wKLvuq
Ef9eeLoQHLp07HjhoUQnSvPH90KbiTPFmDjJS7RGaHTwr7s+b0TbHvBsP9Ggp46oGE2aqKQa1gMM
aDThvKh2phGWRrMnm/xWhCBO5pCWiCJM8AwlhbAcYZQ35cAj8d+PA5kw71GpX0KmmEKHyXZs/iDL
d5hLg/BezLnKoeBkvIO9u2QbhKIlFac9laq9suYUMKLlA6g3onMwOBynpj7QebzbpnlWlNjb160j
c3Wxyh25+wsC5gEXGX7emcFDiWxAu3xjtbmmJUQux+TnjDoXwIuKp5UsklHs0LKHo8Yc9DQ/nboV
2V7r4iuHnLQ2TTDmFTuacuO0Jmw1MXIS9HYtluykP89s3+bSBLfTd0rKH5yOOhZEkTmN5Jx+sTBy
N80or9yptwQ4a8+aMSgIthn4GxHf0QR5Xf+uDLX1rGe8vEVMQvq4rUhWR2v1farpeassD9hknUXI
KFwb3MJFj1kIP5LEjTrmkQ1NjvYE5v+BHvmiSs0cnqJ/V0mxK3NiLGZQ0I7XJjr822SYx36STagE
LANe6Y6T+aHnCZWs1aHOP5P6dDHNtTK3Jjo+NoOebrlUQM9puZTeena56PYhJtNaistQJR5dHKR4
XdA9ZUSFQe0shOoWQZPkp2JlHvJXOJZ8J6DVba/7cx4O4gOQPPlay2rpUOnf6w4XnPuNoBqrqwoi
hJOXi3qiN0Xomg1qGB3IricYbVL1NeheIjSTBPRNdtoXBvpNZ0gjyUYcMEeNIS/1PvOI1GdhB2h5
n2+PwqIRc5CefW1q+4RiekdNYmTMGLl4BoJ5B7KlnWG/a8gqbi3H6qldg58srs9I7XiZ0dW5NCFr
IF9tShc5wy54si0ERZs9ruGUpbCNrZSN5AFN74IwGhH2AwU8T4gN53g3k0gBbVhTGB2Ri3CRijnt
HWrqJpRO3Myb/OqNrlHl4KEStkvaoXNELy4zSvh1eoOpCme9AQIJa1MVuzHA20bwk7lDZ3Q5ErRb
fo4QkKDC9f8YOikKX58DVlnWpefFEy7PAz3+RUNfx2VZIRd9Xww3zafLzXWKcoOLc+rijGVLUYWl
aMbS/wz0uXSy1kx6aNu0o7CDHysmlZ2zGP3CQCeTW6r+BnJnG/DXXCFVrcuxW/E0pwqKcSqVA19g
0xM/Ho7ksIyTftS4x9HpW4qOPsxzr9RnMN3pjQIcPqpjn42BBIaiaC2XNCc7LbIoZFg972/yqOHU
kXkIEExrKUVkRmbRw9uxvITFqj/DdGBHWvpa8ajTbUWOqcl5nwpgFvHGZBlnA2gQW0dAXgFEbarT
IG5mr1tCif9tOQfvJrSNXmRBgtvSXb+WY4I9OvXfOY9WT8cI4paBhQxLfjZ9urcYr+U7X8n5Jc4V
wcMzSu0NPm1g43qV9oKRjPKbjh9UkCCqtQf7iK/7dSnMfBBZzGtqMv4cR7RbHgNFkK5V+VKhcyBo
sqnxnhsLKMyKBv8tkBby/5yF3C5FUELjTMNkQjGo/mFUQItzJ2ub7giThfVpfdq6tnwGgwqA+0bW
1yX2D4MtHhcCa8mIfF0J0kn0WugskSgVUNXgrWP8+7q6If+0nVs9z9W/zINLoBSRjhj4rXOlEzlH
Qf/E/9N7/0JK4F9YWyI2E1+NRu+4012HlCuAvReBhVvoRRczX3NfFNWZv6dzGKRJMoufbtQvR/LR
UY8jGXKNj29zxwRTG8KbGx+LcIRih+uRHEigF6NHe+d66IYD72JjdEnQTHAPBXTH3t/3Y6KiS6jD
Ux51m4UgawAXu519uZy1gLp65wloR844srSaR0T5wz9pjeQJlXHVsKMXWj8JeZYrkPzqoeNhK5+9
4obscSN/+IL/WMUF0EAf/76gNk9M64dyWjruhTsZTwKcgYeI0kxbcptCLX0GA/4/nQ+8RxvWrta4
8wFGWDKng3xYRVmYwEyTTaYDxcpKyXfaAeRI/nTz0UNcn4/p1d6F/P/7jn2Sd/Va9re9vBwCTrge
RfvDdDrrl9H9+5xv1qTK6kM5Ml+lScsafFv2pbV0sUgvPnfKE5ekNf+ufSa4jUnCOCyJuJ89oDcs
VJHTir+8LLkEiI/+ka+JTK5MDokwGBv/dGiKSeDxQ26ysd3Df0/LJ4rXV+gzcr5Xo5LORGe54NJu
x6ewYtdPsw9uRfXzUPUHUBOXb2jzEthXMzbWoDU+a6OS6scG+REFszhCj3m7lWCAhNI549/vXaFU
1fhzx8kik47m05Y2uI7DqoZiz01QjEckGPvqgIWaHrXfW/CSbgzaDmTyqZZgHt4vW7Hlh/Tqy/ZQ
zV+5ipSIy/HlXZ/N3VLQE5hTEDusTf0bQZmoY84juKAP9XVj8pExO0hr4DTuvq/PCiWMPdusBZ/5
6EWhUX32UYzDMmsFTueZaDWNrMxbThLhb3yakHmgwqH79iyrmT0UKVmwGB5A+FcvMBvnVhhD9AzJ
8JmUpNpm15AZsTkl60JqKNBXkYXhiN9JP2sDKyz63gDsJwJmCNcshZ2hnhqkooGUudH79A3w2ctN
Po2pQV421jS6269/mgxEvKF3KDIZRU7ZCJ5xOXxYhD/RwlC8YnLFf/jeZcBhkBtc3glUH7TTNvU+
Vs+z6s70D7PFZ1QWBa2T6hlSKkKSaLDbR65+UQ0gHCnTjsVjfr/CJBUctspmKtFJRSCp6OD4ZbO6
ZSvR6lrVq7V+cxj8ooEodDmGO7HTCp3Zbfyg9Skf+AvpzXMs8xSU3G4iNu6uyNFNabhFs5Ub0ltf
EM84XH3Z/EfvuGw0hov38UKLwxhJ0Cmz12VZrijVO7PjqtMnAP9Df4zlbUX+DmbS3ZQQ0e7vmV/m
jrLImWZeClmypA0DLNVBoBWGfktEHzyisUmnzp107sl21/zeqlKpnSlJnh6qHiGsBb5VERRXVHnI
OXr4FlapsAV/+wCOFX6FSMSNf0lnlCFKSWjMKnYRGF+RxB/Y9hBeM+lK6yjV3GjLGqpvXFBNs9ID
/rDfHMZqJRPf85bh4PsJPefiyt8HbHrIs5j2jRjps3iBKwUkbGjRryAbVduVYsV3WNE9EC/bqVwk
JkklXVgpz77fhMgVsxX6wUoPj47+3LHqZW2EadvUQbCiweCnObHAyRetAeXDeoWfLdid3e991aBe
1aQYl401Fo75m0cojMkbsSzQ9709aRmwEIWQlt48GnFQ3orKXBba9nBsMRj4YewbnPixYh80mp0o
uiqieTYsPx6MCxkgM5J5fVUka8YZsft5cd8X2XfQZaxcmZo2ZP9IbzGuqkk3ZxOW6pLkEMDsCif/
bOgALFZR22bjRsrdw+5SH0d8kIuWylWXIRj7CiOWDCrNCXVG6vQiebje/mdQgYzUbSix9Up0Ctz7
BmWIQ3uCeMeLvg4bb6uHeizxuqfXgbJ+GrkaHkdtUpaVq6DbwZYU9cWmudSI+JSwUnXS4n1av/kY
F5O/q13FrlGP66MPjx42qnN5lRGmXEBY/FDghK/mIqrLbLW37mdJO7rqg552sgwQ1FbRE1Tvoofy
MLft3cHOfTXRgVNsDaOiwBeaGmP/Ly31beD5PY0AYEkSOyY0c0NKVlpQya83MWUvS49y/bIuh1+m
QryRdnjFPQQYeE2hrIvEhEHCiax3gFSU1q4DC2OUchuRox6/pT0VfkJK9+VyQ4vcgzC9WMAEL4eG
8GQwx93DYvumcEIZfLeKIhP9cKljDUcHQJ910v2amXWRB34HU/2wHMxfem+4keLMUy5gFZL15JNo
cMDf4KfJLrOyI62Chb2JuuT7zrkPP4NSfPLlbwnbzfN86DNtn11f+peCeSPJVIRldfxHz15IsfLz
c1k6x5LJCWF7P/yumklPb+iJcVyyphMSkjIyA2x8A3RJJKQCShopW5pnUTZ9O69MK3ugl1uqbu9l
7GZ158p8REGmmNvWVTkb5BIHzEo3m9wdIOTt4InxAYJMI5AZ9BfcJKPOGj4pZXIlxWX04kXKI/Mi
pwlBqxJ1bNwANYTUAZ5i2eHACmzwcpXI6l2Zh1J1g44b1FmFDgy91hkWdHOR6XcMbj/A3kdinnNF
pBSmYtz5fOtwRBElKz0OzU/V4RyH9mzd5+nN0FXANIy/kkD8m/IaTMEClwdieN37BPV2poLrjSK6
DybkRVp31mt8l98jyl1g+crQqpsg2NE0p4fBLkxZ5XhZnpBXnRF4gMIXMtg4ggGH0O5muK9J9fbL
KA755XV3vblFz0wuW28jP+ljoGIzzhBrjvdPxbB9oMd0JwUp81SoRGIzU6JM+3qCi/1l5u+yNyRh
xTOfnEN/F4HAdaVLoCDY7irj3DXBUE4ZmG1Ap1AgR4/JNCwRKTW+JRl32Zu3Z3HQgzE7INvWQVaa
iclC6+CEW4gBScvhPfT0FJupfWDnQGyOEPl+EmcD98eM89cKNwfVLGTlCG0B8Fl1lH8PepHZg5no
aKcHkXv3GV2XoDvZCk5GL5nC4yBEwEj7KI02CRr3mCtuQRgtIQo3yQe9bMYKXzcL6hoacABLNGwL
yyWFj7sre+M39o56qXTnja3nuZGiR4e2hhj5vsdFyga7+i7s7wTVQrmXfhXUNtmxB7+Kk2/OiMh2
rM3eNfCU89wqtgf7TJBAfwk34Ezg+fmK2C94HQvlftZjElLRERwGy79eunOk5DvAndR2CCQw+HKl
lSutWWkmvE9lciNVLA7b6HclNtJbRW1CjZgT6zfu4LMnb4ZQ+K6lr9T2hQxBKHBSRtI+iBIuE1MZ
vHY/iYd19wQuPocaOSXB5fbphflOIX2cHnp1cM99l2pI0/II2guTdNqnJSlqDg5qzlIWKhko2324
Tl+XI5nU1it76znhvh/SH1V4ahkaemosLd7MI3a1TIPh1v/mjswc8kaCw8/QvVk5lht1dylwVGZU
SyrrC49/DnL686t1UVrs7tSJFY9vll6a1fW8tVKcHQjs1ZBwzYUB5SC6iDIQgdPkZL+iTNdIH/mM
SAr+P0oklcrRycq/KYovKwoh6089bfh4fEZEEzHs7CVu+j7mYZUk6w4R0ghz3GgfdE45qi8OK0AB
XF+CBVQ6d4R0SkNLTu9h9QgSYw0XSPJ2c7Z73UoLGPGwms/pQ7nPW1ReL/hbVIa0V6bSaNO4YjZz
7sqFkvXXQCHEsn593Jk6GM4pSpvXLSd4U5OypYs9GzUGLqVcANPjdeLtKMllrgOdZqonlE5Gq4DT
C4Q1kLR6yd6eBGNcyQUraI/hp6W+5YyyqjuPAPd7I+EBXfsXNk7sERSdEglaF9SIwRz4hnxg6Udb
fA8T1kOjgZaejiktjvsKgJHX1w3bgpjVdqAS3LESzSNFaz70P05gM45CvPLVMFAbjAkuy9kJp4gC
vfrhKwxkab70L6JGDXNO6zoOm84e3/pjpY5dM4CQMaodlzgjksng2aYU1pAj/s75ZVtSV+jM3vwh
t5caczbmL5U5MU92s+e/sgaL4WvHTbDn6w7P3Zslk1zOX0S0DbdlhsgfTg6tIIaWKB2YClBKJ7zU
abcH1gT08+YJd0GG2BFIBt1ykksb75+VFfkSn2QIQizm6kkrX8kJ5HDEW2RZjhvUqch3jrevNv91
42ttz2oTyio+dkBAVqx9DKvNujeR01DUx9cPyLMTvumOGlzCuZwQsG8sszWiCnlMUBUhj6hJ5gpi
LpgENQK8sLUtWO43fvwv79rSQw7SKJvT5777GCFZ9VQqZFFl9d7a9ZRlqKviYbRgb5SW/XoRkZ9Z
pSwMSubq04oPF34Zc0iglqLImV/773s+ONpFkRAtTkL89JDLjWdF0KpSIBkFxQiXzCf04QD5Aa8G
fthWdydt494ib4w2NKSzaBsUpe6Y6e49oOAaWd2NRlJqiGZW9YII75wsMQ8n1h1QnOtpw5QhJV1a
zR1IQs/9q7MqiRLsRZSAjLtY0g0bjA1J/MyfMyV2q/RMv0AyZ/OKVi/W71/4RTMIkyO7Yg9B5QXM
ECABeUNafn/x5QTAiyYhq3JVxPmHOD3EW/iplF44UgEFDT2Emo2AxyhBNM47K60y7u60NB2Mq2EG
UBJTlMnstzLgWxlZCUo3xV4w7HZyyUL3kBMks00zqTcG/MJI4+qwjTMdbCfXdqbHMxFQcxHH5/dP
As6w7+Ewe7LEBahlCv2JC3evdXHylKWExkAh2/E5wUSsCKZnvEXOxq74BitObz4BB1FP94vsWs6s
iBVddgXl4vvrfvM+/MPJvKlx3RUbXPqyeCA2XyZZgDZTtVObQhXUzCKPhr3rJZOLiA3IXfdSpgNN
Db0LWH+5iDzYPbMZkKr3j5yH1eGRadAR2WDUfJAgq71EG564n54Wqeu3a0P+0yOwtk5lrZqz4Kp+
KKU5rGu0uWdnh4HNe1qfM5wer0GSNRPW+2YmGw0sXvC6F0G/f7fP8u+gTG8fYV/U3KbJSnXyas7h
XAdJX3D/jSKAYsEhmNOZaW+vQQkkUkSeZpRs5XpQsLSIOIntk5A2lsjnNycMMb9b86QzAkqSLGDO
BeM0xH4PrQ4Rnq7dP83fLu3C3Ga413MqVIF+rp7K5ePg1rodgHgadWY20B16UctogTJ/UMeRn40v
CcgP/Uy9hV+GWJVu52AeVFepVg2mg110LiaXsuj6FKNf2Rgp3RF65+8imn/TCTFsFKVxKkzxrKrQ
0vXAzugjPzE1G3OZhckrlThyk91slfghb3kypjiX8iUum8XVNUF+qqAf1Nh6z+d5bVyJBK/oLXg+
Z/Dw0omDOz9nzdV2ebnM25RlePcY97nD0VvDNuwpjGMQ4agzVeIg+D3l7m3Rmc4P+/IKi51vF1yv
QbH1kFMdZuElnEJ8nLOJ5U2gnb4gHomffLhU067oemSd7o5fOXxVH8Mk0ty97VQEdTLwNA63j8q7
mecTA4npR7C+bQpBhm+D+fNIhhNk41Z2HhAMLabKpnzlFIRXi//SF/mYtA3d06wOq7Tf8ZuWhp1e
Hk1l4HCJ2Ok0yJRYuinCpK4MCWA2zdaa98w7T1Tr7Bjrp8Y9XI2hTSlGQUCsCKAdTy8pFkZWTEwv
Sp5dc4y4WcwtH06U0VbncX3A59mj18y6vmEl0aLyI8/K9971k8sdH+CAMX4fGoNI5FojKqEhMCuf
qqw5FDqEw0W2EIVU0T3kNEHIJY/ZwsRNup1w4tszUh7TeotlMx6ThtF2vm9zImMU7Bm9PikIStxp
4C5iR8AO+cYtst0aVmWrxHV9uzb02MtEdAkAHUOTOEYAwazIRRiZ2V7HIZNR76VWQxZRmCOGuJ3Q
TSb3ANznC51tUKMvi96uQIOOhOKqJsxpXoRcoVenNnBOPbdgp9INxGSRRiG4R8TYvqNTAr4tPT0Y
ZvMJ7AvNj3mAjfceTQB1yPVchFnTLPXv/r/5z9svvYLWjcMn32905+q1ym0v5s+0AwOB1wFvIDzj
vWXztmuY1fmoQBTExF2+40TI5zMpY7naagL9ph65Gxx46kdknAN8R/Y3UZ9jv8DQIkW926eEHisl
5tWbUdM6g33VA8japAxmGcBgMubqmJcu5wAUrjSeXHTbp9FuepJZuKCr/1gMirFVkPtnmLh4wGo1
4M+s011jkUcrvFuTx40aGZx5OJrRUbMkbNlc/LaIf0Fy9pP+qE2fUivW9MARzkpcWpLmwb6Su8GA
G5GrBunGX5pP0xZLhxaKEsyh8Jq/GCVirPqO7Zeid+Z599E9mWBCSLbdh/a0aWMmli3mr3fXN2wI
1WtzELVNqwD83t8n+iJHOOWzYhBKnOoWjIVmE/hcVeyIxCZ7d23OiGMakTMe0xsD5IIfObRtz97r
OYBaU5aLHDo8SInJY4i7aylcHVqNv5YOZEYAf1lo9+OQrfHLQcdC0QQ0UfJh5hLyMIy/+Bc+gWWi
ZRskAlKtpnnXRfddgiazJ8y0q3GsDGEol/Pdtt+ymZz9lZGhfG10nag56Mdj5L+ljsabjbWbxftY
pXyZtm4Wp/IpJBav1WzIQHQQ0ELgIHxazJMDFjNwG6Wq0VmK+UN0JVxLomRxBLUseN4S5U5/lZK5
GWpPO/oLVrdlhjGfwv3G1gDYn/3taxFCrX6vC6wXVw0e3o6YZ3pw9844TdcLvYe+yepLLANZA1CA
FR57qJ3CsllAUgw7//Ex79OF8fTJ0r04RxFGG/iHnErD9o0c6Dapk/FVpi9QHkIbAVFUhTNq9hMf
Hx9mFR9qRb65puA3c0t7mW0F/Ur0UwaOF3lTx4EQXpJmcGT5rs4t221DhQHcIBTxO/BH1K8TVYub
IKK+EwlmXR5gTSf1drzUGBCVkoBrZKR8miqcs2QKrnRtHtdz2n5sUdWqr6BVU5abdzAeZAeBCEcU
92wDTp1ZutYIIiOrKbM6eamRlDoBDVg7YLevahB2m3tf6UGqU7KDYf2WTIALADGAkQkk0GKyY34A
0KIWhL2DBg6UUqzLBHbzqT0DXNFlQWvWDBGBSjFC6wqQ/HqInQvn+su0ibCnsNUCi4xVeOOah9st
KyadeDOpGwkl82QODpp7SSdPlM4hQiCaIerpKwpY4BKr0NMJEul4OL98xCrp4AZfu6HB4zm0MO3E
2KUH2gEDlLkL5rg2dvhif2wx2B19IjyKyOx8x9vnzzpfbHjpEEN+FO3xNY66G9shOhd+LpMO6765
0lIq0P+jjc+Bvz7U0oTwKeJMSBy1nP5YK/ruA59zmnjzG30kNtLBrMxUVLvcOvMBwP+ZBzIqC6av
2OBrhAkP9I3Cf3zz+Gc+e1m6mIo7HoodcVFAO0PIM6qeca3Gbn9421HVlETpOZ/F1WpJ7wwVUc7R
xTIyfWFVPp5UaBU9RNEaacMiueJGmL8vXT4akY4rww0YfBiA6b+ecy4gPU6c1jc9ZkaCxbrG6Hr4
3JPLR7/a1fdYwn0po0oOB0siOzqjzvf6vGB9CFjxKPuuNgmgxtIqKGUXbhSYQSmqEihpCwvC9zCr
62suO/q9OfVSjD53hLMtO4vpUXuplYSJ3esCzkT+wPojqdYEmy4Ggb8x9AQ1U4NbU3olOzl5NBjt
t6WgvPhAcHrza4XU5YbwPVGcR5G9RHoSe5LDJCUJ0rBllXaez2Yn4VlUm9TNr+QHoloAeVE2XNJG
NaDKPTpMZ6qOQkLNwBoePUAUrYImUpWNqxSf5kYXj7SQVcnR3oxfuScQsm1fdqyUVdK13rO+q8if
3QctbGYk2iGWorhCtXtPOUCRq0Yay5CJsGjn4czZLks2sJfchsCk/EMgu/713MIc7QpWClK2jgZk
W8iP8iI5NR5nNRAQ6uoHKEclg5WUPAEXXVo8hQeR1qi1hWCx9fONBGOsrIe/y8t1ZJslxxbJXBsj
/O52Jy++C9rmUpS3od+sWJ9i9UWEZsXF/jfq4/hmVojU6lOl5jgdq6Yz+KI8Dl0TBvqPTax4Gewq
k9cCQvA6xUWvCCj3IHwGZZLC47jHTuHjctTpezIHZXi42HI4iA1cUDLM+NJR7Zmq4yJQym6MDSE2
RCocDjdGUoEcQUmqVgSnYR850P5eMILxwUrAGBhmKcWehvaWBwNZQSqe8J0hgqIjNjj2Jl94Tttd
V4lugMJ65gBQS32YbnR4PwLC2knjVwm+R+tpBy1bmVJHtVcMMtBeHC1U7/ux7w5xxxxMW90KBZAG
CMbO3lHCnjyLYGtVx/v5IhylluOUYdgRqKR7yB5NeE6wZF83OeyB1Ehkgs4gZ2SLbolobuMvI0EW
LaYdAKU9Sx+VoxVbXYLGBqAE4SGbdHrVY6W2H/bSZdnDuU9O5UEy9Ze5eAvLEOWwRtV9EasHsOGi
p80vmtNWiWEA2295YKoxe9CmBfw7zy/VXJjRXrW4YkLHDMCcukZgap3ku9RF0mWvgCbFLLUC1pnh
5LEVzRg7b+C5G7VWDfiJJc+olIFT6vRjK6Dy1BCGlcyWFiD8yt9mTmmCzGhCO9wO/UGTF7IorDPw
h2trSGvMHCiIXGeNAqgpuMhtr0c+CUQCT3oPQP0s6qlhH8rbp1ELNgYR0SBaGBMZ7suE15Z03tII
jmEPpxbowknrYPAwL4LVe8hts1+NzHUhhUtUd0eZrx0+xjvKgAh4HuDAVEDN5WwPg/K1CUF3Vi1i
Hi42XrTIQP/LtfYhzh9gbER7tvFurJvJQVyQ5PrHR+MmGmrJG0tFjj/zk0POEXuUS2tTKJjITLGf
CKKNN2jvCjTN7iRsAH4ZXtRoiDh6xEtvESVZRe3pz6zhmIdAWQ2yLgB80UU69IhMJ8suUUHHqYtj
K3CxckS/ZcjsZYkuJJpcB3g70Y0q7o+DqKJzdsiiKxNltY2vVCTfLhlYfUUK0uiIHqZHLHLtDjFC
hjmyXXQTaBPr37+aWGLe+etzW2A6Vwt7J4LTSdQ5jjugLBqWarluhsScvyvKYjWNayvTlsnjq2QT
2srplcFWFTAohykj3tAeRCVYScAz91lXqdtvPNIVtplr1xq1BbMmtqD/pPXBkpPawGtdf+cc906C
kpOULqSWD3SsbtdK/GxpQZXl2IFWGBDEM48p5mVvCFHAuXGIZi23f2RHscQWlbYF7WvqmRKIDuUv
EYwn+eQJT5GRrw4OK9jD6oIPi3aAEB1UnGkW1KyxO5uVmWuwQiSuLgT/cz+/P1TTw4RemqvgYjPU
fYOHSrduG6nTi8K01rQ14guhxbIQ5T39yaQWMxMdu0Jqjdlw6yIiXz4pVhMkIoqgAQH7wQfWWRWs
wiJCokYUzb4J5fLegj2/xy2NMofMG8CxpSm4UHE3Yn9uy16gSLVy95gkvW1o4Ck9g9z/GVC8vFkd
Hr8UWMrl6B4xRrbACI5KGIIXe4I/PnFh6QMfDaF8dWYzoQ/wMINmfqRXPGYX1R4FU9c3ijieQXN3
ly/iT67bJaMATaPT1RC1SU80rVTL8fehuYyvDeWH21psXC5aqGiCktcmRYc1qYfOjcFXN/FwEE6w
pNdLF7m3o7RBIHmUn4WFFfY+sU97aH097scLRCfaZVqzJc0hSCTTEwcmij58/zZIBR3Mg2j28uFI
sGnuUIQwZRzRcEy7vIqgGyPvS0AZVX5kpcVeIVFMKZI9PsA8zIiPtd7XCajqWKgFVdoII3oonHsW
jf5kcYtJzgNwR65KJSZKuV3dBzQMpITlzk/nrBSs6jIXvHH1tiR6wjhXRiQJdjH3SQA9z8+2oh+r
9zxVQ90ZB0mBZpc1zrq5QM+awGjLgnc6fcQAkerJShYir+sn4Dl++FjBkrWtOKWe6K7JRcUiKK87
7cukj1WvXCzRIdAh7kqTceCev7I/I/Zd2eRbhhKHLnTsn1287N7meYRRx6LAkm7oMqzXBzyKOVRV
PrgiXCd9UtMB8T/M4CTAvjdDC86aLO+27J+Rc6K8LGlZhraHAK9TPW4atr7clxc0gZfiX5u728hf
x4AyauxDaOyo/uRN974vYYOXNBUdz2+2FumELOHIrym7g5OruyvVEslOFSfxBqLwoRzh1OWlRej+
OqNATWkXVzSLNLBvGK3kSkGYigQD7YgbAZLxKQvucIjSP9h3lthRX6l1TudBITIL3s+KUNtNdm4W
7ZXPqW/ri8zPtI6+IEvOYEIt4mtIYlVdNv1HAkPUosMcaxBefNcoUPfYCLOoUHGEbRts5QkztePO
9/Ee16P8ibAA+LTImiu9A3Pf/VpfgugBLga8ClgVXAABFeTPWPN3hIWCH63WPm/6lPQoIOQobr6P
v0n5hEw1N36TUTExNMmJ4VdUEjrHnCGZD/DITRHKmZqZVpOwb/kylvU+oXoRwlPy8EMnm1H6PulO
F5kwu7dqH6wQOZZI0Ht0vD3LmMa2V/8Dx2NXjxPj17dHXe5tSAOjGzDaNzJ8d39siiI+SoffF7Wl
zjf9XTsxgM2f3t9yNck7sucs1mOZJbF4uIOSrzdkP874tXNeC98lKqmQS9HdbhE//rf5WicnMiU3
DCnvWmUqkcOoqsRTJgcpqx78dbt3T/JoTPsSQe1f5dEho/1DfiKzhbYY856uKrCPNsf26iyzmgxW
RrsXb1PYV4yDntFAKKVsPNWe+gYuo6p3msxl/uh8DoUxm0SWFfzM8wJ7nCpKE1sDHnSz8+QzWwS4
JRJkQpOZmHUangIs8ZaXN+IpIB3PrUJqEllZ4RjaYuX4Atc23sGTWWTZlYyei7f/24iQLHgX9g5K
A4iuqSDJfnva4aWaQ5wGP8y0UMkkavu1pcYlRZ/rWa3P//zYJdfRTZhobZjy56fFMDIrYWyHy8A0
ILZ0c4+zZQzhjWLoN1LsnJbdARI57V8ebaCCE6bDBL6fQKzkkfKdGrEBEzj1HWqdcb9A7lNfay6A
0rZUzi7PjKCLX8u7Yk4KEwwZvx30+4l4VDkkWOfsaBAh/0PkyGuqImu5RDRapjpXQFxQOUCS8acM
IwfCk/sMQ6HhAOuGI8prIp0QZB3uUSaB3SWLuq9gVzzLq6o1RYk8Q0Jf/YUcuYROW+ppkcDg+Oig
XquYsGqFsrAtQHGijsJGftfGpad7XwT6/DPIJIRtQ/YaXw7BmzxwTGDLkzRBYWbaYjBVPwP9e2Fe
hiZ4SSIArY+V177dtT6yoW6zFaLmsV+64oS5wo3tthhOhAkz6iTMVoEjzOL5E7kQYvxZXzwAZ1bW
6GGwm08fMZK3MDZ591ZHBVmig4oiAtSXWiSl9KHx8toPqWZluVCfPqwWrGKf4Ktv8X1kyyTBbkCY
IgoT2UNZSsQ4WGK+pk3C/Z2LEo5q0P+2yt6kSWiA2q8J8kNGAFH86IdW0Hxg4J6VHY3owOpf//KY
uUlyhCdPfBmZjZtZmyI6sF6MTfc3LVHlj9aPSma/WWmbGZOXeAwkNSE/Ddd3Hi+M/PbtROlRVQw4
eBz/7P24Rh0JILwn3i9S0fw3k7Vq0b4O/Vu0A5mTC0nNd4AoAYjZ3Ty20uGoYKdCAHCtu5EWJ6Fi
/5QML8W0eHfitNIrFVfvEUHE+gVt/FjqiPHsB9R5P+QeOclrndxHhEJwJhCBixX8y+oxrnpGclDq
ig1BC83pCc461QtVdsmCmolg/0wGU8/HVAgVabA4yAC3eeNwONb36QVBcicyRu3k50xFIrCPiJCS
mJUR6iEbrNc2QU70Vx9xeMw1cwbBkZ/0W+SezcL7oEQazVZ/Cvi5IDqU+wuMaV6FJXkLBnj6hJ61
hkTxydKk2kCSZ67KALCNDXyr7RX3AyFfFVTUwu9YTOM8q+0hTghxlvn1/BH4WeWnvmYQnTrDm7j9
dB2sMEreCZS/eoo8I2AaTzJO1en9tFFU5L3cahBEeJfSfp7iefkAsHUn+oBUlvPeBYYboJX2h4Jf
erGrUZJE/f6F1rJJ3qjQCm6kNj8lM+lZhNiF3QpmdLHrMKdh6j+d8Mu4cSw4npArmaC89Qhs12WO
ABFm82+LdHFNzsMOYfBC9UJi23bG6Yt5hncsGXHAu3xsocNRyVfh0JehK1MP7kcDZVykWNiyAsJ5
Non45HrweayyxhDrk2pl5x3Sais/QNKxHWSLogJO2QZBgsxfs5mYgFO8sKvUnU+Wf1fAclx9lyHC
rrUt442DP15Aa/GzN4q6kylF/NaTWGD6bqWMVLDENuXysVdsyqO0kzPj2HYevZYOOZ5PmfuiAuce
SxLyrIS4hbBIGeI8DBA7xgh8GoueUD7dkYFeMkCBNJBJf1lJpUhE1FxA7UCLTGb4psrZ0CrAlYyx
pfipfOxkbtQbFag5rdXI3Su8fQHllsWmNK2Z6zLzZchLOH5EVhjNmXridkypYNHw9FaupWrv5+Nz
pwVR9+bJ6ynKGzrAtXARtdxXb393EAtMTaMKeoe9Rh4wXiZqqvL2RNI/kUmJHLQVDbl9ekY0hNXO
PRroibCtUnF/Ky5Bz9yBtv5lbaE7wDorJgqH2vvjJOSGcfTDPxsJT766CprUEF4nElivEtCQ/aYb
cAAjL6dkw4JHgTB0tVki3kAx/qpc+zCCoZh+DxhJcbYEu6/HUHm1IVdHp7QVh77ME1ruPAUfipsM
HZQyKyeVLGqAu8pTrEXRQNyTeS/xhojajXFwl6ErnOJ0Ut5PCtFwd5vb73mgPtiRs5JbyBRC6//y
K82gf/0Ug9QoejBjkDH0AG1C/4E6d7hhQnm1Trg9kgvpxnzlQfhFgvZ7QqbItqYYUS/XSB9l+8fZ
GY0G8r6S7wER/3XdZf8ZatM/2J7EJPV68Pxcg2VoVxC9/oz90VivFDt2akT7YrEG88WamhE4rxYP
voIrGO8z1qoxO+qrK+qq36soCLxfemSEh89lCJE/KgIaOyd548eIMASeQGUanpVHoUlwGKIB0jog
nqxVaRUGXQ80Rf4dXZtrERruiYNzv5fVlcvtRjsOzbusOZE9UvHQnEj/GFMZJ8vIZRbvwJXeUClm
CWmESMWVUEPHI/YtnjhRiwIW976cC/ggt6RhKZ+8e6BA60J6lSN57DxmBHIxlIWjpk7SBeBqPtNZ
ZnVPtpZ2NZO2U+1D9VgzM7qmcytZ6mm/IcWPaD5I5u/I/3PNb9u34FMwmYbFne56iCuEDXcTfTxl
Z3Id4Um/ZMFEV07Sebm7Dis36Hj5Wmo1kAu7WEoGTahOM0t/QA1I+YwICV42ImbH9Dhz1UhzzGaZ
wnesUSpYsGPoip5TFKsYF0h2SJC4n65NyRtT/51v0J9N1/I8SM99fZ6TEgHIMtwtOhS9t7tnCIs6
Nr9HqLQammsE8e8KNesxV6Uji7XRBd224oZkvZWJNjG5LouAnJtiERvBu8+a8/zt5ri9dvHfNsc5
AvBX7W3oKpFHlD69e0UeAoh13wM65nEp0JKiU7Af61Sk8lSoLChihsireZCG7SMOReZMUpzV2ZMO
O9g4vZkGuEF0Mno59ZUkmFMLsWyJOfgtVsh3sumrpxpVdsxWn57DEyXaK+PZ2PmzTAf3YumwFnem
6kFd5tMB6UIgkYmnV57UNnHqd4ykME2TVVXGcnGuoWiiErVAzuqQxBsLFcUsfHYF5YA4/lNgV26N
Hyzo+VgYns3ek2H3hG4BHmB682eu92JDWtfm4LRqJMG9KB9bjOCAlpL3Cr2fmQ2BeRFC85vWE06q
TviyoFg7C85VsZGPUz/TBHXBZ3v3pib72OEuFsRZAoppv/QVyLZCproD1eKgXnH7D+/vbeEfQREY
PBtEzXM1fvhvORNAe9x+7U/rglXrnC6ifsnio49BUr0pGvjpzycqh4W9LWBRSOn+TxXF94itG78y
+pgQthZAlvIl/7jmXICGiCrMTsDlDrpHINLhzgjvuestGrWJDjUOvg+d+nvWJKYeU+MLkcIRqLJB
qxnatGcpm0WHX1UuJzE8pJKnaObHedyi6Bi1mhF2EyCQ+UzSTeTLwxwsmwyv4tG1HfLMAzRpnuht
9sBnsh0k6rzN7IegrOfNR5PMTmYdVsnRAmmuHJtUslf3q6nxRHemlZpEQCN0+YIl6G0TJGlXkqLw
J79YnPCUSWDFIe82jS20mzl+A9vK/gZ6dgevXkvQcGIgqKrFypWQFVINjPFelb8cHLMxzdiR+3ah
XPzfK0snFY3cfiNAa78WN3DBKxpMkm8m1MDcxUwoqZfzxeCXAsXTZXptmuX5g4/cng+clFsTf3M2
j+T/qPqJbG/1d6V/trfArrqgOV0d+/M/Uaq1KMsnKDbQPuNapQzWjEeTPts3GJS8ZuQcrcFRldrI
cbm+XDl3mLld4etRXwoQaH6QvZiJwp7QbA9dlW41/DPAgf6/ILafBL9d49lV97yUzXiTb3+hryy0
zKu9LZRNGf3+zoKJ9o63e3HM1uLlA15oscL+3dDFMN/++O/7N5QBMkMvhyri4aKoGL63itzwsuhS
5TYkQABKJUCo4l0p6dCJZWZV4SUYJ8aI7XCwZ/CCN16T46l7dKA0m4r+5OjprU3xUyUUwaZNNVaJ
09ae7Wky57bx6exlHpJTI5XZj1sOIgwzEPqgnzYWICarMIsyA7g6FEX+Xg97/zk/r+FnYH3KEL6z
FOJSDwCJFeLCiMNdJDHrrmy9ndCuZrHSzGkzNOGMoIn1AF7MLl8i/XHn0hnXGUAPzVuV3ngm7jTc
J9KNMjeaQLGGeW8hXjddbio1HN/TolquokTePtZamlX+r0kUesHLFSkLAUlvV7CzzGsgPI5SkfA0
xE6k6C6Ueq1mwZQLi7caAbulk4+5Id1UlO7bRnfzAwCtHtjGoxTwz613zCA78o7k/wiQ+jLkgDNG
4rG7/Our+NRgcjJfoJ8/Q5s79HcRjHPm9Kum7+M/cbuQ/Af149vEnGzmUTro5N2R1jSDu9oZ/C3c
bd1DRYxqhqQAW1schcol1XcuSiZlDKmi19XW7d79PnbsXZlT0dj7ShRCovxEbalpaFqch91P6kzm
8+2FgoOtdZ3u7OVfxZpYwS5kkEGxRNDbgSIoGSQk6WN+jXVNAFae8TZJZ5gTA3fdYAopfwBrGaDm
XocS08GmvOdDdQDv1vzL0UMARaNH1CkuZEm2pEnW95f7UZKu1c15lt6lsE4/tvOrgqlCvMYzE0la
DoKhVH4dGvbojyJsu5xekX0mhVxDjt9hqSlUIx8lq3o2bN0fn/iWi8yODS7dBxR22DknuTEy27iB
IbEBF7TiPj/JTHJL5IFmmgGtw8e1xTpGF6C7DcpiuvXj0TA3Vvmsp27jYtKsYGUDuOACPBw0mDNG
azUZ4lGZUJGN6I1sHE2f6Lu/OZPYkrT4aJxTVSTOP9/iTj7J5RTa1unCRInRku3WtM5R7FTj2byf
hdi17vR4vqr1B8N3PHgY/VYCAGAN8/aAxYFt218fJnNEB36kGjCXq+viRd648IfMxANpNqHXoTrN
mjm1HdRHxiJvV8y/W/pmCNTXtNUFdm9YHxGkp9CKf2kVjSem6RKHVZjpv2uxlXt+ak7n7+LS0tvU
I/vns0YZxCcW021xUNmfMLFs+QMbsmfoBQeB5HrGLuNrIxi6UrwAxj6Cj48+Sq0rtfYhs2i7ZP+w
rUCg8rbfzJue4qYY2mMvwJf7Xkdjri6F5ldYf864mPfhat6OYqnfwQ6dgZ11CLrHX5iUzJ/iA5A/
TQfQ6TV8pGnZajDXiYlHm26F9AdP2yfJvif0US+npnbMuybrfXkUDhJX+gDDY9nYd43MxDkPjCtY
jFVo7Wl1LEWFmM6hh65yjrnuqpdS/HfG62/w0Rf4/ACo6t6nTfYKnUBLu16ViEHJ1AS6ohxJc0uG
JuCWotySVp2MfhmGROGRM6KgOTOL64ryNO1eS2lafJfUTKIt1EXdbyw6ENSbOsIlc43XTEzurrsC
88KXnB7/2o4nnOc1CY0MI84cuQ2JpG+7/FbAJkfY4An3M6GCIy6bqP6OA79IPt0Y+NsltwhLjfwn
kc0BqGoIOVHzLrcsyhGcLqSkuSUUyNbdXDr08M906keELMUonJkqq++p5+XjPRzNLmmNkpdg1Dxs
ouGlh+QCh+QMIs6DbOLDANj3mIzsWLADtV+mr8gUWs5ibWd/GGQUrBqEQHVw+OyMOkUaeNZJesPc
uL2qMKxEetHwE4spBeH/bbC+R4SkQhmq+wBGjk1wSg1KabOXzN6IyHc3jYXPu3UUed9jA9Q6tzBt
GAYZvYrw0+2/UucGpjafjES5/xAHqfzJX2hoy8LkVGNLL3h8KlRvyvCML3qyqXb1uf728HEJfbDx
DjH1YO+DqwQulRLEjLb202rlPmg8bNbf+g0fVrnpbtHx0ZuBX0QQCmGcIajVryrzSpaYSQjGqYPi
sTXMSqo6MWDtAVsLv/fFUYhlaYwhDK+L+Nyt5KUlIo3lxWwvob/ueoAu8zkCuQgogRaIqrA2wEaV
Oc4OH8Vl4RMOGRb7fex4XA5lHikTZGLprmurMUq09ZehOLAA7y47CkqGcvpOnexp3DYm5MR++QwL
vaRAAs89RoMAnlCxdz6j8GLY77xqugLoC2Gd8RDTUY2fb8YDpQB7bEd8QFz+9flj4I1DcJS6H91E
NZi8YT4SJ0FKeMpygf9HYKJ7khZd//a/Ciyy+EVt6MF62GZUQsLCBnRf6IQL5dgm2xVGquqG4oDT
QwMzR9ebsGRZXKG1P4R9FCQ7RUB+3FkffoilkJbEqS2tZamFpqWu08XjUCYUsnI0PVTkYqSRMJC6
D0+7o/0J0M84KVsACTTvjWFQn2OrLa7ZItsG/NhEUYQJqJkrtieG+t+4lXOsFIwY4P7pCG7Yz8N8
zXhsuZK6PlBNh8bkEgSsHpOmmDcqSABThmR3xVvEUqRrriFdTRt5fSp6OLhdh5CdQCbspeCkEdXo
ru01nVBiZN7MhngS1sPY8oBdG+YupZBkoPJyNfbE/Q4lxY68w+rAKLXO3ZSuSedPM81gJobRj17i
Vvz97NSykqu8F6yc7/o85bBjZjGeazjJBvthYAiiZXvFu1Mq+b5X+epu07+RsyTPrBYxoJGAEiHX
vQSN6avyVlbH3uAgkgEVfU/rHyCqPyhDvShdzgqrXSioY8GmvCh6wB6tVecyAREoeXvQnCnZ3TxE
nbe9KxJqQ9/JzQk9UBlnNIoKCftluoTno9T7voGeQMa2whkwBrWRF2bEhfQcq+s7V2gT/PZ6yWub
rTKcRUcmnsl/ZcTRdHS7xJCfgsTxTQuw5NUaJeLik/cwyhXhuxzouuB0IZ2ZXK7tWPaLYyljXfo3
xMv5zTdyNVrVMajCkLgQ9IVKZCq6GED12bIFYOZTXKa5UXPxVsdCU61PHwHWBV8hhIn4N0CULv0e
VDAS0CREKomtHmZhcX2xhDlP9A6JziDQ8pucAgHqpCzoj9tpQn5iWVQQm1YFHK1/xpkJK5wxDG7w
YdSUEr9TTL6oQ6dc1mYlcTZrk6/FaWa+bO1DZ4BDOX/YefkU5acaEWkrA4UBHuEEL2KvCu84DNx1
wa+WvCgXxvL3AFTacPzZiFCXL1qA1BT9ymY9bLlNDnhnCbSArUkxqDB+VhR0Al0gA1YVh8CsHZMp
6vzisO6WOEfk5RW+w8HFHjXwKAtb0+EwI2xYKgK2m4fW4w1yXzHUrfbMW7flpj60IGXJ9LazLiAz
xbZ4IHNGHxDT3YQ1un1c1+7zG1Fx4jJ0YzRYBzgcrD56bW0fYrLhucwINAA3M9JqLk0yyWi+4WZF
ZLzvvFYAxoFDSBKaY809r9UEHIDFO4bZJSmDJgCbhXQb+3NZj/fcf/l3R9HZMYOHTXi3PwNZcd3t
R0c26Jl3Nv80cCNPR8T+XFAM0rO6G4ivFBlQbG5snux6x2ukOdUoIbDj10H0uMtJSPkPJ0nsU3Ng
Aqnbc3yT7Cub18BaG0MvwOiU1YcSZJcwaKf/tRizUQVM5rY4uPnAfQ2EMtjux7G09x7kBnRHQWE9
HUZByQBpNWUHoZpLzdyFqYj2A9XQCVB2W9v3o2RVOKqn+2/xdmuwXf4gyV2s3laq73XT0BdlGVtc
RJt73Q+lej4tkv1L+h7B6G4/+XqX3AgAKuEWaeaCgao5toIeWhQzIyvYQM19A8PwkP0BJ8j+nm7w
V2sj9RT3OO5u3UvLGY+KdemFkPMqz76cGXH4D+LMFTpV+tNdBo9e5sGZoTRNRoGBen0VvNfZSj3y
UID/t7inCoSS8mh9IAWconk1OlWKX705q25f22Eww92JfVDaA10srfSftVzqW7oWgGTJBlGVI0Gz
oOC6W6E5yYKSN3GxutKtymVumIHghgBCdO6JcMJIP9nn2Kdjll88MtifpgKh1u/XLiDGooms2aot
TGU4NIvxYQFVWcP2crWiW9cXzzqaJ1NvuluZy3SQKWaqByheiiIVTKh/q8lFXD9AUGZhacOPkLdp
VRt68ETlwmoFbU2k/xHOCzpbC33qVnpYMAvr5mhy4yBkhfwffcye/y/4+5uFtuCl7k2ymBQdtt9m
B8X3v6xSWHUjfw4SllAkE36JkrufB5WFmIPzhwnj6/zmR1G+WOgWxiY8ajAKRTfsMv3VjaGo+IuC
shxjAH9oImRqU6g6EckSnOyoZpL0mcgbL8FXlphiDwKyowH55Sh023MdPpG3ubtYjuPidn4AUOC7
sHDKh0/9kKVheyA2ycWrkK1ftcMT5y/+MyCJw9v0YZqYObGWII0PEsI1uGd935Rt+jhsYzYQK8ju
T0sgCxdxOACqB0aLD8vrSjZG0IDVunB8hJj485kI1PwtxVE8nZvrPm5/3hWB1eRpTiLeK1QGtIu2
72ojwkvxcC8MBVq08fzySyG+rnyLjdfymtSCoFW10fFr3tg90OeEkjM0cjy5+pgpZwhdu1hQPpsC
ye9t5by9ca1uu+Vcnse/6C+AgdZ7XNOBhumkbTMQRDbnBUxK0MhPWkJSiECnxmn68b1miRTd0/re
H1Jevt6UOfRk30yhZIRIiLqJQbM9Hqz7bvjTTL0aaQ62/rMWvM8qUwnS/z0xcqJTZOYH2hv6d4f1
RK9hUNWsekuSiymygUAzQ40ielUPVXgcfiaZdPQRzGlkavC0YbYQr2BBHtx7BylYDfJxb544Phm1
jLyiqwRug4G/7HdURZOatJDm2+BiQk/Na5rC5h1jStMXHWdg/Wm4w4Pz+7UGT4BglLDYEaawRL7W
7bazo9cWADp4c+ghavZc0K79TP+AiTm9OdqQNYYbuuAWUyCDDYEQobBOwo6jEPtjpi65zTxna16d
ko7NVGmB9RjYiNP/8e9hr27qH/nKha7vmwZfFPODUclENn2mI2SWGeWmPNn7JrSmWE/7jomnr4F6
M8MJA+SRSUK0Ofm702OXyPF8YXzWS3BVuN8dCulD5xMo2djd2S9f2uu2h2CKTBuhrhsKHG5jZqgd
J1UuN1A28zqCEoc9rne9Emy53GE6YHQX+MaJY6l5Pa/g+AZMXY+inryrabY33ik9NDGVJV03+yIs
ExyQ5s85QBFimIONHRCylccARrcXF3wFwwU6aZaGcxiEM7LjZ/iD1GwC6gn3LL+Z7VHj8swU56fC
KLHWEHutpgefk579nkGBGaeeC+ig5LjGceA0T83dbFteqP0vTilcs6kjYRY3kavAu61vvc2LQnpJ
PvC8wbt5JJHlVPyelOSqXjmov0SP20G9gWyWzyvVQ/0xll0XM+OgKIZcjSuBErE6NhyUp0DkmBKo
W7an6RaZGYc9bo5OW/90s8oxYvMCm/yYwv6g1Lqh3iK7+cOY4sDlVrBdVyr5Bz5zzbqOxZdLYd9f
7Kw8cqbbQbB4ofq8598pWqNWbmERTTihh4W0g7JXIMlyZDoKW2NfFrmAimV6FPpTw7N+WCpIPQu0
0dgFir2ZcXPt1hemjubFdyHkaJfPiDMUxVOoVI/Qh7lYhL6nlX365pjA3kCXjxEF4lWPWS8C95t0
0aCvJFYvLraGGFRD+VlRaGdyJxqv4+jlmqLy2EDjkzsK181susv6Mt1WmuENtSLwzZcGFX+RkT0q
RD90+mL6fY7UfRRDxJl8RlZCbHN1c1Ld3t4aLKGfM6sVSmjevKo2C/0xq2sy6KhMkbqAj+QvFlaB
gd41xZSMI6n6hSx88q0xkkSpsuQM98jNJD0A9/oN1cSLDoiEp7jQMv68/OZPYJzaZy5kbhKEGmHT
Ab0+C4bUHZH6k7FntQsA2hRBhmB5GvFV0XpbplZXHE5FaPsgm2hT0wFA74Ondgnyuy9sOaPGqojk
uYgyNAM/rYFo0tj1cVjTNkv0H8s7I8NvuiGAlx/EqDC1Rpip3Ub3eAdcwdg6S+wojfN+OOAdz1B+
5ys/47DItyIWImSZQg/dfMrL+71o3/3D7PqC4+QHPKl5t1cGVGmZ/NDPdo477+BQKbs42LVaLOhn
E2nJLSOQknUcvlBt7AIi1vn8d9HdEss8QZI/njOFmPYWKGqGWatFDjP3KHxA7V7o98dhiib41y6e
jKhmGg6LARS0qXSqw0AvJC5LN8QpSNy14bjI7P/u0vlAMJVJR2/57S444QJ+zUx0O+18pyW9duxD
PgdTpIRnwh1aw6ify3cWX8yMZg/k4BpnssgjRBNYChIV1ffq8mH1Xa/eT2UVDLxRB8L5JNXbM2Dj
pJgCovy5jtM+URz0YI/Y62bwO1JSSNp9JwWSxWef4mBAUA75TYDkZokoRxD4hw7/Pi/uvo4fUcLk
442TfCkkKN7KudgUA/3ISWerxS+tMYITPw2g9CUsbd6jz3kbAzTgzBWEWl2QWhWLh73+p39cSzG5
l9r6w90ZqH/ALdNiM/JNZsDy5kL4mzFtDKhGaVkMxOh2NL23/rVz5DK6Pm8ayyzr4fL5igH3I1E/
qwvFOo1THB1nyXfvRlFsut4fgrdscxwhEiBmP5aYZ7QEY/qmSKo6HgRHHQWtVuhj3QaSvPX3Ek7o
KbeDqZH+3QLIf/UJPMXx+fFQqiovgwQ8kS//h/JgTd/qCfkoS7tm39RLfaCz1PsyFIulwzPo1f2U
uJIwaVSbwPqq6ZtK49s5QkfHA8+SxhHB+GGAP9pDXVYc6WJDkBPOGbJiZDUfsPJd0/hjoPwGowCl
8lSJ3K5tPfpl3LEFEaGfaXL7HOGqXW9nd529ILwCV2IB/5SsthHXkq4go3G8uoBKP+RxCvN18qzD
EL8LNTXZU7NgfCi86oZoGYFULZGzQMBtWr2jqUu5VbsCbQlxyNIpoLTufueDBMp9tyU4CngMINZd
a/Z8uAVYihLbAJvM2B34aMlON1kZN6l7i7vTUku3kBhoB2DRkLrFi9jwvmMXavVGIdbW7FEsXjLR
KVvd4WqgWE47ZvkY07TWGmij6X19jB+2EU11bLK0AQVRUBNeaKp5I/OrJB9+dbKDT0lOXjedJ3NU
ZqVQsDmkjBHj6YXHmleDZQegWnm4vmodlFS3pHdbmpRTDOi1WVxXghaxVWcBziPtim+Z0nWUmztw
S2A2j/h1qwvN5e6b7f/PrM//mGA2eKZk7Js5YVzkh9z/KiabnmBGkc3ktmNcU+n4eblri37cYikv
q9iutk0mz2Nd/kU1y+xNd9iBJ5v52mu0Y8COOgfSWlJHQ2KqiBXnYQAesZ0m4sZz90L5ioSVLh+I
JK1qa2jSqnkM9A4ylR6kCJBXLzLpQ8zxQcvoHnDcLLx0yFnZE6LKKWmG9dP1f0j9vP5Q+eew00Qg
Dr0lkcUrP/GkN/M1sNABA3VvKD96uIxI2oMn6HADe8fDYgonm3XuVmvziQegksAPpRgxhirYwBBs
5I5wjW145dG37qLm34Ykbf/D1CL4xz5RdDA6ktfBv/xegvnRhYl6xR/ldQqkny33TPJDu6h+hxy3
cQeGCFkO7uPiRr59j114oBIDTVa/Bm9eZfhkYz7SFS81jlloWba/tbN8QOHteBq2Xa1uwptLTyov
PCmDvCOi4YUs3TMHe4Qun1rbYlCRDBvGkk5aK1JdQEoOD7yJ7bH2PoSkD7ZtaLn7IeG6BX82EGmv
1/Yl1a+Vi4r90iO3YtOmh7utYfGXJSQiD/TXvhoITFLSAN6oH6lnrVnhRjfYt0QrQqmfQg9ML9Af
5XjXUGly/omKLoW44IBFoZVPuXhCqRFu8kWpWQRPRvDrUVz+HQuf2UE5aynRztBXN5wQqMV7sE8z
3A2nsLdJYRh+zOuVPRmETetfVTsQnQFg7jwhcVKrZ2KyKK/GNHSUO2FujHrvnX/YPP6dkC6EKaBm
L0BL3zeAJzDqpJsx/adLyIYZyARXhuu28kbUmlWKO5lpeTGjyLYzUklNhEN1xjFcpejb8peMTBTB
Ks5IjassdGxEOzE3b1McjL0ov6b4P0quPfQ0auWQKztnRzMfPKb+mgXTJ+vAg8zWh+d+Yd9jhmhn
e6IHKVp5ER6Ug5xpezMYmLTvLHfkwUc/R2h0gc7+7ffdHX2moTvLX3skpNsLL4MmjsGYlfowKYlV
EK09VRZMH+hDlcQO8ZlZ9kQWm1s3y3LHRQ6bKigQYdNKSrG/ehMio5XsPKFvQ9jH2azmno7mwT2U
zUVekslCm7Lnrn56NIccAiJ3D94p+nfhhGPKDhueXqr9wPSl7vLxJnbV4uLABa4mkK/kPxspzuMD
SD0zKna/fs0zFckOEH9lrY6A9i1zs2QAY/z6x9trvjZBFwCEtjk6eril446XZXUE+wAqsC4/kGNt
LwksjHvjPOJVGphawXqLxHFrW3/aPbldsaIE3liqP+zOxYpoVq8HXSxI6b1sUFKA0vH8tRuXXO37
d3h70vn1UpAJaQY5Rzkbj6kmYN3nH0NJBW9IxmyaorsGyMaCA08fb8tLhlNf5cExg1DPcb9ShJkA
u7Y+NQlyXdL8ikchhVzIr8E+pLW0GQYllpPfWmscvWo2tyVLxxvStpnbrdCq5dOQVhPtOuyCxqGw
qLukdBcYyKb7Brp2Zd+Zr47Gy2y0+ZyIZHl2hkQnuvzjDC6b3Fq/o7v+BzkuH+SBvGHrOfixMrhu
XGzNWkT3EJ5giZTINo3Enn0CFndDZ4L4Ht1fBLbAFimbYp/kKOT+Rpv2Z/PIPcYk7TnoJ9YYCL+r
Dx4M1P93nEg3tDSyVy4MPiFbfgBOrB8pG5zMBI433R3Hdj6s0snC8YKhJ4ss/hzNj6LUuXOOcJZ+
YQpSEKtgkozYx+8P8y69IuQwxw24NSaFWG14flU1iGymgr/1dndIiAZHTfPL+eUi3I3wHRQQfKmk
5Eby+W4DeqVRFIz7sORRhsz/vEB+Po2RJpiaZ0zTZdovO3nKzoZqaMfqKzJvixZPsLb1HlAPyJ/5
rcP4JcUcX28p4XRH59sdKyFymITvBMiz5POz8DXjjEBcLI+uRRieRSJRZq51ICiTuApC9IfIPl/t
nIFrEWhkaMC8sCkIZaM+yWq/Kz8C4gQwpFsNHxtnOa3XOpfR8z6+peOpcj5QT0U8C1IWYxlATeMg
eMbA/AGVNIvey83rhP+ZdMjVfaKDpJAv/20TIbdU39GF4Qc/f9QcPvwm40Z8IHDkoOXib5+c00ds
k5JM+/HkDn7qRCmEfqSrfO+7wnGcW720RShpC2tDj6kv136uNnxlonQcYv2JX7mHX8vr3aJxwnqi
AyfK8NQRxgwp8v8fQKxWcSrwPuvks3NStaH3Lyt6uEcnsxF9/U9gPkIm6ludqwgL3zdfDGbGJqYq
yMPQV2Fb+4xI40XCQLnDkxBtUb/vbT71MOKTuFou4t+S6zFWlrGNFk+zGCMtZcTB44vcLUjyrXN7
KZJIQV85L9QHGwm9cQcXAmKD7BALqjK8JO681bu174J1w2X+n+YpLpaS6LRas4BB8ygOPAzwQvmG
HvkzDFqNdM1hrqyH5a6tP3pyR6jKuO6Kw0ROjNFot5MFl+p1AmcuevLvI+2NO2L5RkZgxVrllkJr
zft/JT4IGwvqfeQZ6zbzpynzIg+eMR/EyhsUEUJ0DCRHNAQH0/KHO7xxk3Wz2Sfuxcx699g8KkE+
CEcFei1oLJa3ZubTNIS3zOvZmD7vW/C9OohuNUV9GAOF+FXg9V4kBqTfni5LskEe+cTRcF3z62y9
b27nNpgbQjguVjoZz1yxJFTxf3wl9o9oFahat8NBCTt76WZ4AzjNBKnvAKDKV+bjk4zzLJ2lcZHu
h0DghDjvcxRO0fe2OCnObHnVrtHLlU8YOi/0eG9V4kUFUM2I9K46ZX52ZnXaELCczElJAUGqtUqL
j5TF+e9+Kq1CI6E7rzPi46+nIBX0n/aUKdHHpTmzOjcBWvr6GZ5L/qU23hZRIDx+R8n+PA1aShr2
F27TY+veLRKZjg+/oxUyr3PCH5gnB+qOwSaNezCddSlLQNhVgPw//cQp7NtXhz42AEzyJpocWNkN
/lsrblTHWkrRi5sY2to/SW55EO2y8P2ScMJNMs6OT8qs3cRgQLqYgDX7n7DEnX0UuBECOmma+8Hj
aB25EAgPz6ENvqSCFIph2KLS4UZ4QIVdKvP8i0Tj67NLHcQ4Tgzm6+r3wI49UrfJjOidGoSWNyAw
QR3mMfVBvD5NV/sjJHY01Q5svPE+ZwuAeoVhWWE+AIwxaU+j9jte8x63QPhvEQYXBYBm/r+45A26
h/v1ttsRBM+oNDD90mm8EoFIQta/eZZW+YIrhcNbdx3eg6Km0ATVBVenQ3jbNRbD0+IvktVjvsxH
TnNx6ML+rOrchmG4Sd/jECm+J0Z91oGh08qV8wV2WZHGLu71BxbPx/d3m35PfPpqi4qwLPcsgqXS
073FU22Pdaec1PIDnYwRHgraookuUrXJ1xT4bv606XRTirAw6teV5UMHiqWdUVhC+YLN03mzOw4Z
oIlfoaBiCwyczaMP1fnQr6IoZ3abzGEQKJB9luNNNIEmL1ogTvNVe2qLRC5vIbrCA8CUuJIxrwb6
g9nzxMAozEJAt7isbmf4xYVdEzCqmSH87jy7BVtJKLZkLrqQWz0m59qF25e1uAMxl/5Rr/fVC93N
Q+Xby74Nz/RqZKRupy4KH5CVwpLSedSdjH8bMsnJtzB6SKDcMlBSB4OEit3IMTvX8fRShEb9uPkc
Oqo/MeVKtMFjzEy8p9yEWYqLx/zPo9Tq8sUBoRmruwPVhJLwRl/eKYF68PRJuSqVWxHj7+472eJs
dN/HuLndPyYOHAzVy7iDIRYHghfZl57ialzalMFJFRXJ69iPSbwJNEdfbmQs2oWPdoiy4kWr/RT9
IB2vEui6FKHi4miJer+/RcLF7pboOrs8qBf+qUjGVwPjjp2nfg3d3h9w4HfZN55fE7RdXt1miI6G
kEsRiZRZZI6ZZQpHEQPJ7GgJ5yQio1PbLNgHQK+oXb8xgDoDNI76OGaBD/NRso23rJxO1V2AozB3
B+wcVAZXShL5l8fbUwWxJAOGHta367azB7Y+CEbRraU2zJG0nEKQTb5kOMKPs3QlPhPA9GFDfB3W
Y1Ndr92Y6Xt5FTgqwr/BJsE5pqwTsHO7935FuxjgjdYFrbc1VqE6BgjfgyxuCqtpv9s4/I1HqBQV
P0ceBsC747XohVlz5uLFeOlq2U+SspdPPJ0lo5KPsCyCZNel9aW2VIPAT2+95vg0wZ5Rgn/03t+m
udNV+WdHOTi0vrVf50uJDvEwpeFDPvnza7qyO5fzbxfQGE3LX+3EWJLbB66p7Yo4GYjiq2VRPhD5
jmsLu8p3WOi4tO6/AkHr6mnh9MqnkIJufHMi5WxahaGBRmCsHZ17H6hB2UCe6gRrGYmWnB8FAmdR
aa+IVTEi9U0WOYrZPJ7hbwQ/JeY+hxytGaA9Tbl8TapRIFFuFG69lc6BtoBFpAWsJJQ4zPTgmEiT
Nzj/K1kZ8JuauO31HDmXDAiWaaJXBVaKeR1bV4rOr6eUaIMlDDoMvOLSLYHynmgaELSZAk80DWPb
nsUgqGl1sIDrPJIj9KP7vl9KpCr1BHqQ9Evyl1WT+OdP9UQC4twnkUUmFWWrdIxD0wKmw45QxeHO
DdRbIa2Y9tA867nolaRXW8bRSeiAKmxAFQnqUXvomLBKw465GcaDi3Co5MnMqEbJv+gGJY42+P2Q
e7Z1BqLp5Tkb5jGCgtrmw41swDMO6002w0QgfoMPnF68cKat+dhQs+9Hp5o3fkgBGwKg8b3Gb2g5
dRZvh85O7X6MlmJ/6ZHoEYsXfEExTM7LooIJMIIwbOlCE2fJKWw6WlEgDSOaAaH79p2SIsRHjsxQ
Rw7YynzHodZMgqptWQsGPNbBTwMavmhxnGL37F0odskpoDbMAFuccLFvlgiAW573T/6tQedPmfYk
ijr4k+UwOmYZC6RvKFASpjjgmZgjba4pDBhlYFclFwdT6O7eHqUxwxFIKhOm8SNhbMQVNNEpCQZa
7bjRalrfFoS/+Q363Ml6jlx1sip8KBUDf3Ldbq3eX5/j9oDReTC95v6gat8fvSk79AgdADjcMavl
f4i+ol86NGZmu8wM6ILC/hnDDK1oPj8rVcFhmCQbFFTk4BYjTOXuUOIxbT9MpdDY0qYY+gvSDBAG
sRZw+nzB9aWxG1bKON+i2xG+/wdy/3MNSwJyOPhiBmk+9krWo1UbNjr3c+DUTnb0y0i07XJvSK5+
W/Lc3D11BulW9a2nKIAHGOyeBaWut0GpkaqSLY6ngRCO+4B1A+bsjPEfZvNh6+hJAwBlasPJt2Jv
BNICGyt5UxOm9wXruhO+dK4+7ULgyw6Q40sX5nTJi+tW2mo+gkfTfJxJTUbNDfFl1nL+hAhpGU/K
JgyVe4X6fdqSeqj9O9NJ1D0N7BF75UwFjYaZLd3quF+l4hlQfYywiYkaEEoYULJcwOhwC/LH8U3g
naRhizcutISFnm2lkEH9jalDjgt7C594fm/T/B86SCubgQC3Ug6f+PJuH6nNOIBmJXFELYSCHi0L
h26V1xBTvfJSEcXcyDKhGUDdTTu1C6XkoSamLxS5qEhwRSHHzIx0huKe6LMQrL9ORxAkGVkshPXM
agjAKEwGoh+masTssFyiX1S7YAswzLXXVL5vjuEIO1LgKKAgB1WR9RMsgsyz/rJP8Chj8QMbi0JN
0EJy2TWAXsjdjk+DQhkkmgzq2WN6Ov8GwnTK+u3AFddCL3J8DH0wjKLv68y64MGvsW9cqoaZqyXV
/SmeG438u6AismgwyjEgPkms07UiuLsTIt5MLJmOIDa18xOSNy6mSFj3wBqwn9XxYizjGcPrl4X8
EDrsZnsVcs1RuIpY/Z/NgIxCl7oHtiJKC/9Yu1la4JM0aoz7CP7p/n5AqL1D+Z65SU68u/jt/8C4
8srhXdZBA3eX7s37kGq9vFiRNqK8K9BC9CO7cJJ6hXtKnkcqJtZsVX6DDgadK/9NrOKrakE1mR2N
fWbB+xUEiR96tRb9nYU20wR894Vl0Ijpq8x+nzFop0S1pSAH7iFayZwmsR7bAHjsVYHSs9pzSa1T
9ENRwHXnHQ/ShAgq5NZh6pufBYvr4i2uRaufK4tyxcMTTkA6PNQpLLHV+5GQoZsDH7utMC1mB4nz
kp5bITGcgJpCmlr9YD/tDy220nZccoRPUK26fELj1XcVRctMka9PuRs++bIQ9woyt3N9PpvmXz7L
M8WAbl4KyMx1dzcyToR86tMLZpIn82s3iUjAkezVZmZYr6QCNtLoQuLnMEw7dTQj1RaWQckaKpdh
5v/xnNwBkOkmOTE4LJng5l+qLH377+5tWQqzHpRoIkp9vcjkq8SPbOyzUy6cNxrS4AgIPzolgD24
RkkUp3K2nmPyvw0yE3HRnTeQxdJCdQlGijX7wBSRuNd6zR+Uc0leWFkKChSU+TTaPfk282hGtmqR
MNcyBurgTWrc3GGH+LOOKg7Vbe4z14F10MNdbkd6s+NFQJ2R6Ae3bvi6hziLWc3thVrPb70yqY4b
Yyi4n+F1CtrLD9V+4aXfsr0yFvXqPUXfIJqashGigr35uSQgeqWoHNDFCdyBr5Mp8VZb54x8GiAd
eaLV/KDb1FUi/69W3Xjg2tTeqf9DD8jxeOlJNY/Z6l6kg2pAkPMGGhLwnlSEHfHjjCatKkT8bRyZ
N5r383NKfgomOxRnrqgAj7tEyzbL6CK1MmSQo+JQH2LFB3rHtAPBE+yQJYRR/Jewj3N0t0LY0kd4
bFXFQIEoaM4P33iy+H568kpfEba98DvoUtBCjsTqFmfRd77LUA+m0SULIxhupOhiuhEO2HJmgHZR
yhARpYdomj/Wwc2dZn7VGHpQo5UkwMSOtDPdXTtqAbDxJMujc+wT/2LpMmZhF6r8Qzcnm2BD9T7Z
9U8j4/BoILWIA5+ggzKDhiNqZtJoHCpTpNh3QdMJTQZlVkzc3q4ZGH2uUCWmvsmcIn2Yf12zpAqw
NT+lXf9aSqyCrlcsmNILL+xRWgnmVEh42cc3YGFH7JwFg4BLd1L3uewP79R0N5f7JFWYYIlqs6Eb
sM1x1MZt4LjauTXasU1h6xac4HtIKfQXcwuKty7l7VZtkcqeMIQ+GWkM5bLlymbD2YSrRXh4p6+p
5Kw6iBHDMVaLdkD8aVOEI35mZiqe7e5IPoAr+mw7vfKeoRJ7gHEUOlFdDBlEPFzvaVWtXQi5euj5
yO3RtHpKxcaN7ZwnvHtqNUPPpbLvVJn/q3SvCPq5zNSDa7zPR3+ZwXht0gkvk+TbT3EGgeTy9xGk
/Ao3+qLlJ0bPVxWQtLg09Kv7nCni8tl8akDQhiYV5C0YMPFDeE5fmDSjFLUHqxa/Q1lKuhujbT7k
QFpTRtm3z2K6DIxN3BzXdz2YK9nI/WnotsjVnYIoxiHjpW5Y9ol6U3AhOdy2zUr+C2Xpc8MypGgj
1/lmoYewCWyPGfFVkN0Oh73zPn2JJQFCml8/YsmRgM5i+JBssk0+DEeyPvuiP0nPvmPgpBYnC583
YNuk7R6AO8tExDOB38lbFTahT/HAm+vqEo7CuV5sGuRxv84Rw5Q77Xy+acfQ+EziQCFMtvNEZbLZ
i/apA6ogbhO4WXJSM2J3v9CaoJZJiwrSzk3jq+mKlYWVaGlwpA7qi6OfhAAPBq3VjAzWYer4goAu
6BUzyjXEKe/DgBcQOZTRscuz5+yt0EkQckYvY9IpHYOA44RUXs2E702voQnop8dhqlfCJTnBJLuU
JOFsGfhfvJQd22vMUw84Vreo+Nm/TjcadhS2h0RQSmGX5MeUhe/PRnOI6fblQZ0T28+CDWf5ZYET
xg4tWyye4iGacVl/42q9WLMAUZQtRiP19zaTys/O5vn32ESa2+SJ3/dLOl9TL/tSWWK++aeO9UuZ
wwsWiWqqkgDFBW1LGw9+I8iHoFF6aHDxdQfh3JjdKIwjoV+212ZBgjwfvjZ8A3ODIdspWD3jYLjF
AtuDqUS9btIUME28jKTGrcR0F2EeK0FJb4llPvjmcPWHreinCnYi6OU5VI6GQYq37UMEz/RB3S9I
GF5z8BwGSg0q6c9t30fBjJNwaIgWaZQqc8hHtktXGRNbE4JWYpZwKKc8c9p7txC7IrmJXtLXTN4R
C1sIY9swpnskXRs1rmKkl0qXpg2Em0FmrbOpzq4X2dWsIyY+yHYlCxVOuzrTa/Yu7MYR5SM5nt7E
+N7TeIKr12IBipglmztex3VwLGaX9MLiX/UXW5T6sRKrFrvLIiDS/Zfhwn0bSQgv/t7uL1jq96HB
1Ws958FHJOkXaupjgtE1Jgn4LUF7RwFTw9z/3usOPsJzIRimpkpPHbW09lV/8IJ6mm+r43lLmMqI
PlOQtJhaU37D3LNvKYeAn7yW/QNMwOdhU2g+PxV2vvP1hkDggcgoQY/SY4FpEZgUL2uS8Oq9UtDN
ZENmlN5p0j0QEX7IjlWophXYfNPEHnU4iECOjDuJF2I6SFMuT7QGlLYCGCr4h3TpvBxXiJuwhgTd
hlcpcoGd7oIESH8kRF5LGHK1P18A9KOLW3BVVtfg0KVbLqnbJn2VmakG6cdWliyZP4El5BF4Uz7g
eKyDhU4lfKvem3PFoU1HSvFM77nbIoKacRSLXuNlpp31qsusZlDShOmyJ7JBDJ2NpMqZSZS21IDI
y8q8PvJBoUKewpWZBgCjMfq8FpAk432JIGwD5Dtu5icTZYUKvmv48IxDRt9IcSR+MPZeH90hG+7I
uYyBKk6YylPnuvQOTgPIwRR/WqTtibhn7DqFwiKyh9+2yJn8HoJZ5kyOiAbmxWHAnVGfmZGFPXJ4
noE4aVDsqBIJ/tWazfyw2ev5BIWp+wEguOvej+3K6RPtV2taEOMQuZghXJ2isbihTgQwI90yoN80
xuTXV7suvZsc55jBRgpvNHlecE3jL1VVhuQ1vT7ciBlJzixlFFwvlf2Sv48OlRfEV1LQI1nVVqlO
OwmjSXKGzOpVRDY089yqRslsw5j/zlOvL/qwPZ1BF1gY1TOv8ivCQUlQwXxo9bfX6P2iiBa8X66k
oxoOX0wjRHpskXYd2rzBz6vZfIWMPZZqT2z7l21LEuM02IAMBxBU5P4QD3U2aFGT7QC3ZCWlFfgo
RF8qxrqXg/iUJDQ1tc7yRGW18wX7k7uCy6XlH3QyEn9oCj2mHsWhFHsbB6QFXSofW9QJZqzqf1Iz
h+EiUj0dS1no2HwMkVfUYao/ZuKrGOYOlVasfmMsJXim0/s32eN7Mx/fmISX72EwQh6FelzzdvC4
2y7+nmJgE+REdYckqo4+8tdSxccUDe4le9TiNu2yTGSbokQVcDVY800ACd4kG4e05OmHZ1nWDz8/
ugNGM4SKPcyu4EW+CmIp0MZ+qFuAJuPyv6wI22MWnqhJR1qPzG9laIZ5dXdzC328JOsvGK07mBRb
MmTa4GpI20r588p+tvweisOtIYi2Z2dZJKDyqUGYIa7QiY0zg4JvsKoYfySw9QL1LBhkisKOaQOD
RZnJrt+XRYuC+oZxXoFPk5V07/ThZ3PYhWV2y/cFVCqHzAVAmlUTOdJHc2eVwt0WUmz84pMSZHaJ
F9UU2VlXZekZeqcXsVbQBirNzP1cVE4pgTDoMC5PbN9VGN3+1Mg9IPBWXxcKAnTwY3yhHS0XDNmM
OS5g8NeaJcqm3aJsWM7EoW9zQ+mxwwPgb5n/4HP+JNFUp+10nLxkLjRbLhDGZvmod2KIZW+5fcv2
pb4mefmWX1epR4oEzEF1YmnMNEEy4fBf2DAaklAFIvPLuMKEtlxTPfqh1g65SjxZHUtqrC7oEqL2
C9uWO+5GTcNYTfi0uFiAv0LTJu7d1sQqKCJCGpAzSiCEq0Vbn5P2FZkSCPXYmMextagrirjMG0Oz
DOYyDGvFBEgP4abeqIIiwUZGbZouxSsTHhtEGY4hOGOpkkVHclm1Eml7dqxV65xaRMmP/HGvGLOZ
+EWpOMXpvf4WFyVr3Wgcv3P4NUl1jpPkmLvWzL9F05PJUlB5/fHVCQos+lnv5y4t54W0LQEFmzKB
hZ/tuLzK8X099L9+DSX8uJP9uvqO0XPeR8/rf729xCRRLcr12Xby7P4RbmagCDplQ6bDIAFZYTOO
UoA9y8Vbq7LYaMYws3l0ra1lD2tk/MTscGiMKciiXZakxtgeaFJ/tBpdb4rAIZwvwubi5eZPBuUc
JgCPAwrM404cjpZ+3gXhUqbnuADcTkW1e0k+BHKKY1//U4rbRfxREopwGXhnPfZM7s52hmP8Q98L
lOqvZUfADtQQZ+YOl/RzogJNotIh+6hCfgIzrXgPzchv5qtjm/2ifOYjilH93f9ASkJZl6VRMo5D
bNB9xGdgQWM33j+L9VBnurynMyCbmY0RiNrnL23XxohZzbXTi0lPQTRKmDg+bKLH/W/EvUGEoVro
1JQM1Hi0/Yo14ABYITUmziACTKNF74k+wjNAIPc31opxnk+uZcgFjliT7EIXniuLikT+tYj5RZL2
BATu0GzzPrtU7LTwh/5IH540n7Et0zVk0LgMp2QwjOmn3cskaeTech9zsOQAAGmRASGC5lE2Vekq
ww7ygtJ2NEQ5jo/bpLpUtxg/Q8mcKVgWYSD+2bBIc31rtp3JFF8+VfPzTIaxsMYnFqL67HXIhSPG
MxSTORy37mkNINIS9smrkIeXrYB1abhvtVu0ttwOxui7Apr/jJcyT5llaF3DNpTNGKrJu8oG6hiD
DgVEJqH3UkuTSXt14im3hFzI5Wi2j8MLEKbF5ID7HIWoZf0B2JnY7SYCxVSEHr9tQaWPHRhin7TZ
PexYiwBoeQsD08h6NsMCBEBODvajJmMQP2y4CrJkaJrjTJ6jHpf1S/d+otgXkcIm2og+/43g1/h3
igvD+d0CGEirMUsKQocuW7+KnLhnJZqB4YWWJw69xmde14zcRjmwB9tPFkLzv8a6aDdMOKUG22P9
9Uv7S0Y8TlatEqFz4/rK2Wc+aSVZgNxnOusyUKF9UjZVnicvDqchrABL8Gj3JV0a89vWEzVnPAuc
nooxL3gFtx3/u5Rbf2a6A/fIpJQd97YCjL4+Qc25SQbbdEgwLarl7SiGmuKU5VniOnglsXw2x+xa
30u3z8K1a8oUrUYIzVnx8487zs95nzWGBpdMBb0QG98OQRabeNt2KsoXuavC+QhXboT5NSrspFni
NshL8Kt+vYgQF6N/bTFRedJ4HVRmjNTbGtuDIBI9v5jkJGMb4NUBLqWCYg4R2gBHUx9aq8+Rb1iT
8TOqEc36kbM300JpU3TGCE53fm6Bq7OtJzNarSFSQat6X6mmKsuqK301m5ZOEJUvUWdqVHKJVa/f
YEIxFHqk/rLKbaGatjzeRdF0RLzBjkSmXWyWJexo9VASm0aRt14e+deHgOndNmN/3q0run+bm/fM
MH++2aHmDUWsBP0WEjdR5oXlApDP84yM2EOAw7EvHkVpFti1G50DBrswhM1x+qN5FpUS373SMSek
0n5evTBXZVe66+LtoiH8JvH64r4rd6DmOWqsj/f8YskC0/3f2kS6A7EB0viZN5JrfhEF1TGBMpMD
rOImZBFDrq9vGeox5c6TEWnlPtywKLyt1sBj3tfdFpHpHKkLlQd0iGs+DEDqWjopJRRVWRIVACTM
AsmOroV8uAuJDqruol3l4zmOASoVSX5aEDDEY7srb6m2fFzYsAWAcf5reUjedtW7awRbs7LVZhFX
Dg5t4vNlOU5OVgWUmwPp5IgszWzbGTlor8DwWIfPOMCrIpzVwKzQfC9ONxFFPE2XEW0YKxzH6+I0
pYT+jAdPQOjFsbxEXfCsIF6Ly1YXJUqGE7PRm7bo0YExfp5vWVitx2VdJrxckmjaRp9+wh2L1Zr8
maMHo5IWubj6l8p/QDQA6cRv82xJyEKieLo12WveUw1Aypjf5lN7QDe5A6keyqxzGj3vBhynEnhy
EwxRaV0WlIUChi5OoiS2D8XPelGjLMcV1wXGkCM0XAimjq3EmDVKDPHxAi5IOGenBkzC0V+I2CIx
Un/lWEcp5XgnPStYK70EfZv1v4V++OihWUSdzfUpqf6S3WGt/I+n/ZXx4F79ML7gvVPcHNdHHVDW
QpTosHVMi9rVmT2Tq0DclXLLDXnDtF89z4jaUvQ1tQGZXijSI1r0VLuWghkMCdMW2YYejlZ6xNKG
Z+z1HzftXxFbqqLH4FYKQzW95Z6tMm1I5LfiBEjV0baj2oPRYe9lROKzsMy2/zw1bxGoLD0Zo3vC
Q8o1Be5XDr19BIkwcG/yM3CkelN2T1vtUiTebBeCfahPn9KoWK6hacD469LpHmc75tU7969pxrbR
cHNXYMmazDrZHYNgnfRWdBok5j1SHo3lrKGSpzVTi9dWIE4mxbGiG/rEpeCLNUV1A7Fy/P51jBNt
K49Xhw7JfVQ9FIdIj+po9wBZyC2XkNYBoiWBYll0c4Ruy3A4qLIDoWALHrC1YvMy98+GaQOXlYLR
thuisqRXAuevmPkdR9rtgm2JZa+1xHtcFUChtLE703ELQbnKDHdc8HgIFjtNmzy3LVNbw02ofYpR
Vhu52AO/5J03fE0RZZmxD3D0Y4p/+sTZkNJN4lr0+T2dFGAX1pVeKKrZSrHs7qF+yofM/H6sCZhq
dwf8lZFbXc1HzHVqzjkGr9G5x6HQF2mKqCrLfOQ0kBDLUbgrwiRKKpadodoKMH1hzenDZVMfJiXI
5jLF5QQ+MXu15bJsIOABcUinvDShVX8xgqRICES4v1VkL5FsU+vc9qXVRUxPQ1Jht9SRMsATXS4I
SLQyh1CXgXnsavcii6Oyarvtf1FnC8HeO6n83yuPdIO2FzOdlE3YGUcvPnznqagAch0DsiH0OGWd
QYsyRV1nTuqL8Y7yTfF3moK3z8N48qJ7ZkAGNunGiSzb231Ie5mckgBz1ZUIyTNdOwchOPx7T6xY
+EYa4WbGnUraGXExYYj07NQbLbEXDOFky355NG+NOjftvz2+L2dnMNeH5DpYur8/b0djTS8WOXFZ
Kv94DzyJ5basvAWeyT3qdlYgA7hCBqyMfoIt+Es8VfwKjFtBreU5L62jeaSHK2MC9y8WrVOR37GK
Q4lCaEvncgiU1zypnJZJdCO/EMNy2iZP2aT7iii/4Ek1jx3o7HhNdS/6lD0faCKzyKyp66ZfzxzD
xPJssUpgVt76wdwsww92+P4pbj0MfodKEdrLsTStkSedFJc8GX4myVjHxrq+6L8eXX917vxOsBlB
++0rygtpxo1GH+T9ap+zd2hJ285FtyV9pvRFddDzMxkmaQmPkVp02E6SXP6BYIcgpXCFZvtc3zHa
lpRuU/kbV4e+Yar3GIkiI4ObEamDg5+JqXLki1vzI+SrStW94wWvoPyC2iF6EOoWNV3fyxGMi6/h
8JmXW1xzOpKJa68b+dTdinSlGxt/+r4pchAl0QtrKiWLd6Q88wM1/9qVFM/+kjw3HqSH6gsqCcfg
g1+Uujwh9rpaV4zjdJg7M7TSoFh42whPF0aboRNRD4IScpLg4cZmQs/gNfn6Xmkgpa5Emc4tb5PJ
kGDT88+rKdp5xTc8a2Y7DFMC46PFFWrpJZgXv9bL42mvMpx9GEWkYb6/FrQhj7tIE4wy+GnPYqsC
HVaz8yvKvzo82W374DkB7/z/jI+hev4IpIWGHko6jbiIVIDRonAooiXX6kcDxkOn2uhvuvfCo7ce
jvmB7mllNn+enJPyLCAzbAkMH0Am7VVzD1U/PEiqTK1jbkZ8J2OjYZJNae24dtu0KnJ2eAWSHIty
Tm032EArU7FlkKaFA6hkPxB8yPoPo/eg5BSdjh0/I0xqnnJW1p/KP/tWiFD07BMXaX3r8Wd5Kmze
1ARAMJTUgsEUKZfas76fHHwTBUFOEkqD8RVJnmknt5gDS1hyiNQE+2s28yODMMqhpg+o5EPPhuky
ooU5Ca/416P7hbhJUrFxyeYNgNuVe7jZcGbsCo0GGVMWvwSqliCh6QIxKlnbQKnysbUI6i2B/qnR
XofG9NfCW7w95wL9Vp4GxJ4ahTQD82YL6TpwuLQ9VOu+UR+EoqVGAuGNiAG7UpUGczXkca13jLqZ
CcRFOvfmDJtbWsXLbjT3TViD1/nhDHcWJUlGCt6gV8y7iE955Dvdc7OvYuyI5Jx12sfXY8HsPuOj
Nq+UvaqOl/9ioJ3ddnSXNELzp0jRvht1nffi/54UR4ON4Hm1DGlHxJ3uLJ636wbiGTSLhP153N1S
nv5PUjenZoWdAzh0Wqo6TnlJK75FeMmeMFfTE7NhAFs3Z6Z71vW2UXXj3cSS7u9BkteSpcjiFGAB
e/K3/g7qiVtsDtbKOu0f/HSB12HBbyskcds2dp6RwdlokdE+/CTZFPZusx2OQYCU3Wi8XPVMUytb
sLIt5l036482JEpbHfTuidbZioOyE7fLRrBTobqVOV97qnDoYDojB2DhRLOW3+HtMoO7YP1M3WNc
iaTPN+yuqqZOCXupete5UCwUutXcu5Xd2f4mWq4k8sJcfPnMKQQtqVNSyoBrA6uAs2sVm+rd6QJa
feVecxZrixZTVLxeAYQQjeYNs/UU79Tn+h13omCeYbfrTgto3rgymKZCCxFn+nlYQBi5kjryf5o0
5xpMrdURpaDj/s5y+WnLNx/sAgXHVbfVn0qw10aecMSE8BwPw5V7Jz7iOZDvmAZdG6W+1yjOezQS
SgLyt/lIir1JpabrMWOE4vOBbupVUxn7tv6O0SAlxsVaviWWX0BMbtxHbVhn58nigf7BGureUPRf
rhYun2ek+zSXKN1WN2pcr5D1G5btHGvsO122cndvqYtvo0GMpsXU7xpgPFP5XTlUBqyIDITeBb8f
mSqYm8jT5cASRO2AdXPLmE5T/dQ+2cPJ3UviMSz/TIKK9RHCsHL0AO8U+ioG8+ukNram3K0FxS6L
Wc8RcP855F5W8TXS0vEUCexkEiA1KZP4M9Gy5H3N+OdM2MKvHB5v7pD01iDeuyvqNHCN8au3HRIQ
zJVhpEEJHQZ7/oLc4TcLhiS1JiLYvJMs5N0Nc6zB5SI9wCMuOA3R7zzhcYT9a1aJ5F9lxmnWsYlF
IIdjs4s4slBxJkSVBhKTFswv3ngaXyEteiN7rRktstYA7We2B2GQTjs82hW0vcISMcX66TzkIPNw
3J3snyRWhJhiKUx0SZf1OHlxjs+T+cehmSoekzBMMtcF+SGno69pTMYQjKm8kXYkpOQeiisO4W1g
ZTU8QVjEUWEQcx+fzKADgsE6P7EKgzXqx6AglRAixZZk0i0uwbMgN4mfArewMowt6ymsZFX15811
wNhSrR8b3virAWNtkXKSkmPsCYtG1WFnNmgdqy2b/KwfnSAmuvfD+rYMALEY2VrwDNcdISViEPjP
SfAg676NgsSfk4II0Lt9JoGwwORFl5aH44e6ybttzXlMeTDhKIfNorKCrJOyrA+mDDWu5yla/9M4
PeBqXI2AQd6X9v6m38V+DnUIH7/pFfOKEkJJPIHXQOJZB/LdFi2B6H1caOZ8Q81aWemIy6XCMW3K
sVpy0GGAOKBXdIlKvFRJ4JLjptuPhLOaqn7BQJVQAeqdHkfbceb8gmO2NmCLiEbf/0CqoJLlVtE1
3mknuYTu3pcAiuSU400eSPvFNOmE9fI0baA+h98yJnwkTIag7MK6gcicayzOS6yMrK0G0+Pe7z2y
FA1b1moykwPT20yOnQ4CwQEvMtlqji/Sz8GRDh4u0vqm/0tkdPOywhb0qe8sEAvHDaENYiZbV9a0
qMic7q0KOJGxcBaqF2yO60v1t/XKDXFKPRbb48DrynvRKUIOLCnLsAyeAYG88lKU62MLCKueBXgJ
NCb1Rz62DrzpEIfJMVSegnMZmPGVQUMjdM5AUEzcRpSo+K2ZDpRu1638pDXp+il60q3kGGnFubIp
Qh0XPsJjZNodDbGL6TqxZ9UwT6UuPlNzcxj6LIJ5N0APBTbp/dnEVyq18F5PhROHEYMwA9suBihB
UGbm2vIG120hEFmcJ5XCt28Ft8eIfgbfmfaq4wAVtmIkfKH5BpjtyqmSdQYfpk2qeHOwRQ8Mrs53
4s00bM0NNagSEZSUgV9wbIhjXgv0GIz06+kbMRfEh0gzmW389eq8y13MZpHyvmy6s0KQrZXomtmJ
Y1L41jcH3ZPSM+AJr0ZrmFYQ7MOdPI/AYVpecImDM5FkEgPoGv997R/IQlhra7v03bvOH3YyrBvF
F9wgMe51mpikeqY9yCvNodV4VmQftJ6oYljqIhiHgXmMply7+GTIRp7JZZaKgrDvt+Durtr8AC5g
uSgzYycY/d/16Um/rDIYK9NpEB2yawMBMmBHX/hbNst5fjz5b7uy8fyW64qF0tvwT484L58Sv8Lh
OyPNdJ4oCcLR6E14Fczyqwa53sP16vMTbf+ONLXLNqQGSJ15vspm4p4qwxYAshmtzii7xIKXgFXW
kMr+dLicmHsnJXED7zfToXw6sQL2sZQEP1txIiderEzsnuIzqMntERPFJ/7tsbSDKBY0i4G7B0qj
cEQ54WMs16yHe2ZvJN6zhQ9a4DjdHzu5KvX+lQL4/IyOdAgA+9ITSnkKsY5M7GpIVnS2f7Hdnkh3
aIvP7IrCEn87GTAA9I7thRBw8h+Dzq0bhP89ySfg8M7oYq+brahAoUjc+jvvqvPPtLbejOZxXdGk
q+4AqRFH/mBR84Zumz4lzl4Il/G4W5FHRZ05KHtUY7aQEwB3w0IPrunt0/5S5nmOIbehQMDhzWsH
bmobLtsEe9zpq5cZjm2eHcSjBcy5mCdvAVvRHKs56jXu0Jwwq0pOry6ZxG1Bt5bfjteTiJome8p5
gB7uex1HJFNVdQr4X5g920wkQhA4iE7zT0K0a2s0KEkilOw/GsPq7FIbafErg5fnK2We5Qc+ytOt
zDJf2O52SLK5HpwTDETSpXJoqsBD2NOINoLFItML63KBO9VgE3mb5f3Y7+yczq0euW7CGw95zR1J
5jbx0e3XhvZgupadzprupsbcjSlsr1b9Burkph3gD1bscGRvYUjwWlFT96KZXveLV7gRRX9gTT2B
BfjzHjjGXCONfla5mwg/yQSJ3KaWGvLctINjxszkcqfoA2ozkaAbHswL6NjvFQdMR6bOGyPHVNy5
OUiQWC6FhW5cZXRq7w9IjsUrfpLwEEodOTvNWTx5Xz1BdURdSy17L3sX+oNgdp8TNgc9J1J+5Xz9
fz6P9t7Hdg23yxtZkOA7861dC/sTIfgZk+/qHVrFO48ffgQBCNB4em3dWcuVjqSL0JRxOUe2XszK
aRFOJARfRV3Cb7eJMerNCmgitcPdZzVfuGa5yyiydPyAyDxu84UxWv26ulkrZM19Nm5150ePG76w
wy8Ncs0/ztd1nTjrSyzM4gwR/uE2VCzfIZpVjWbsBLxYRZe+pZo0jwLpElWMj/Dz8yJUyXht/0tp
lb1ovg01ONCJw/XGcNvQJjgZe3RuidzTEOsnyDrCfuZOTAYsgzonxOPgfAcFLuP3AdVMTrf5PKcK
6SgxgBUKaToib1yVLGOVp8wdQj/OpBcdZReMpiTdppJWpn/TXrHJ9EAd+FV++7klfwYoHYhVozrq
RHzKlzUvBqiOojGOwN1ouNQSdPVGgkDPrw9FyWz2oIeiZBoLFRiB87l8MQ6AgjO8FJ33ufMPe73A
9V3NvKvg/TJKQxIceAlrkFrMpYQiYqtfi1UwzWQ0luvh8F9os3pxupUj3q/qcUF9xce+BxvDi7vh
EPRtizz5Hjb2yFafaEKPYfrcr/oKvuKTgnVNFxWWNkuWdFWapA2oTY9C8QshXddVHkTJNJRB9IRu
opf7m7wHKixwkmEcg/QHDtGCf2csOJZOco7h2fJ8UkQFXiOIOTaVyoBgpe7xdrZIQAwz+Ld9fxCW
+/7sh4rixiCXa4n6IZvjMn4oKgvsIRhHxwWDiRVY0AZz5JlHnNvLx6idDz+Ggf9EHBUzQ8Sg+qgQ
WrCBYNMiQjJSJ9IOwGjY65c4n/I/WWzQ+4gIDf2jcc+Ei2+4WwXBmgRWiJ+vC4r9OouTPkaIP8+0
d+u2OCoeGDuC5rdaa/mRm8hpsJs7sSUcKsT5nehTokASYMhI2xYkE4RG6nYG1V5HSJTcts6SlOPe
0kSkGTTwHZqvFXpjkQCAUqJDMET++w9rv9i7y09gov7CKZAVNi66eV6uuJYaF3yP5kgzvG4Y7eF8
o0+s/3FqSsVPD/oSHLbp/9vip2lLtv3uQZSb16144KWoOfSnV9oWqQlilwDIpRk2brejzOZ+fO8V
wnaEiCjn2eev3cavRKyUncW8PuP03yjdc7s0nwGBbwZJwVqnDRnbq2FBBlqGRNMGzEpkkayqr3JS
jExUq5oEUTj9hjHbzVtQaUMvt/g90e4RHMIqxM9qawYcmAX5uNWpV6OIn22oFjY85M7VuY43l2ev
xruNSaVLTjrabk8FTVT85Px6/2lZunFF4c/la/dqEVvNiFgGcQfkjsSB08LfzKNYLKpp9Qlujl+t
9+tGLUaaSCsY3zafYAKz5ssEMIN8T96NExqkVsgXR+KKFmqfNGo2d0cyc3YH5Ho7T3SjrVJ0vZ0P
r+hT7B50aSEGfgQezprfNfCvliGlrmwKuSMfA+1nFn2/08WKwxviHRK/F5lOeAmrm+1UnHOdJ5gA
oUAlCRKKjtPjJsnLOBeR8gsoqOY72s6nDaTCKAJplBBdJnyAbgFQVhMhOk3XloCLvK2m/GJELW3I
4hFgPTiqQQh04ZP6GJvlcSgJDwKEi1uybRqQLatBCHUR/zAB+k21Esl9rfL31+1kbzy/c1/sZjFJ
GP7Y8dsbIVgoEtJV3F1ccLpOOxpEeCVptvZEiZ8IIzQJ6FryH1rY/3h0axTXKjFO8SHzQ2i+dozN
8PHxhdEqRCd19lWq1tlvWC/aEN+38LoP/BK5k/o4mZDNlhhk8MqyNS11nFGBmC3Nj0RKcF32+Adz
GEF3Ky9UQI4mqq4dNupjqhW8fhykp39qOuuSxutR7x+E3cI5wsFMBfKHNTwyFQDDM4MN10bC8Dgx
oOSXf5+reAC5eEhxjLKwwhJ2m61+WBRoFVhAdCyhsIQXRNI9JDqWX5pKCNAIDgY7sTq+koYTLpfu
1K+mFStz6pdJZDOiQ671N9d8XcwgwgBsbT52lnNEwKQ60ocwIiDT0sCTKh9FbXTTWOZqYa+wwl3b
TOACC3dXC84lF/Oy9XmwIzxraxJhQYD8iMlBMWZmzhTSj8dCQk2tSjszshVu2BlN9xZ3xYWMLMi6
esEldp6E7mUvKiKct2zcqTNC4x9U52oog3A4984+GqPmcwDQ4P3wTjp3k0sRwDUoItYau1CX4o9d
MIuAPZPN/ErZoy/S88liI2eK5+zzlwGJCZf+lI+vfjoQuPlZi2mKjPMJLYu3rgIhk3y/3KNg/8Qn
nYtxphWY5A2mKiKfLIfU0vL6RHZ+mTzvnTZvbtZv253Ur//DxhNyDqE6Tte9vtp4WSZJjaw9hskE
BgASgQO5riFnjJrtAvCkT/ZEkuEYAyNo+hSJU8g0vmu1bOpx8zqIltr9aPGFGTFh6UXaUsleP8sQ
/tEBKNblOtutuashM1lhYVdB7Y7fHBO2zgwoFsf05JkNOIZxaI8W9cGMuheWZ2DzP7SJ8fHgUSLj
eAMMWI2jlYQnNu5tMnEtVCzMpqF+mvUx60KGXlqM5EUdTkFvw4R4cP1r4jQA01O1OkzPZXVToa2m
n4tXC71LPWg5oULYmXdXcOsQNbUWd1MEXU85HpJsQNmBqMhcNGUVmK92Md/HxvZ/q3ahMLR55ipK
pp0d8W4evkUg+toXjPo3N0Wd9kpM+gIDm1BinUxS7GFZzISOUlpOnKJg//L5G8wXfFWQCttfkhnI
fojZrrMJDee/Lwi0FOzX/blMp45W0WqieUA/UjefOp6Gjqke3qGHkpRuekKDvsKREJGJ/euP3bF5
w+1GaVaMwFh4tdZsNWsjc3BJPPmtnWBvCklEL1N26qTaP1pwIXv5x0VGvhDVFaJb5F9QPKLHkjND
chJvCOjAfQfeFFSKggSKLlB5U4k29AOjtWpgtGTQ0bDi8oQggsyWFqeQItwrfu5CmblIsCCu+tI5
/ozT7aN2qS8tqa48bDg9gTZqOogZyVm+mcKDGz8lquRQ11mFgkHHkWxvKI3vCUH0laAPt2FNr6Xp
W43AZ2YtFhNslAjl/vCL/MoaMHsTC8Rac53qv/NTc+9k3lC12HPLUoMYWeaMKjJqqFMcMX+d1ak2
lhTqvCqNg+T+GfC3QInqGywWOC2pvYCx68/kdx8Py1Gb16hhW+8tZ+6OZBWsPLOAXgzH+JXuFmS/
ZLl5MtW/cRFENi5W/b1cAdSqSZLcZ1WKsbqT8dazTflUPm+edDwJIuc/EU2Bx4qvNrvVcoNlY/YO
2phtJ6OGF5YSq2u5bgH6o+CIBxWa0mCmporXt0Rvkah2BdmAWe9r25QWwUlX6b+XLKdeUkPoX5FH
/VrGJ39Ezdiz4utC3Gg4J+dTlaHSxnd1n3DCUz8VMWeURszz+erbW0hcIM7kgo1G0BhDv6o1UMOP
kC3s6uv6pUCRG5XHvoyByRdbD6IawPhZSnPy6h2hSutqHppwX3VpzxEBOcUgUVgQSfJp7bdFIkDu
IbA6gZA5qrCJ1GfIYREbVVMf/5meFBSkBQXrB+3XY8TH05UFhL+tMxeLqf+HY6QZPuuzzX0fNq68
SmAB2n2FxSCPl5nGRfdhv4CtcIZDxvtekYLRcWoV6XdM/eX6nVk+A0yySBA1G396KM9mWPJa+yQc
L+7cUbNnBOP72ylmNbQoRJkGEgZbZSXkVQuQxJjUmJw4kGs4hj3UAfvF2AXmMrvzDEFNBvZgzB6A
1jPP155Yy8PdJhGS45UdGc8ty7n+voSXQcnD4xb1CEvuyZHOpko+PnNw1x/v1bBz2850r9T36dpj
55F8AGxIxb9EOsqIl7cgz/rYSvfTK0HDai1KnYxFZENVGZxKQONKSyaKyQNyNwj+jaZhwZ5wBcP2
+IQbsQDlLL/Tqg5tfLVfYg6BaFCfEpDhs9ya1rfHn0RiLxrTLfMIpsaqa/DMc9oYPMGunDEyKVOz
3GgNbZ6+7dPBCWOG2GKyhPCQ+FS0wEm8AUiSD/yzeLZYGq5cQXHcJR4U3cJeEQLLwzgjOtOHldJv
4c5y+/PtVIQiotEq+xyipm1XbekAoLn2hnP+aitHXTOHl9ffa4WhDVhGxSawgnBL07CvqDB2lObU
6r+EcMk0D2jJbQEbICQF19M5P4KImSi/GAgyTmQZYif9bn2hqftoMZ51b/HTvCKZxj1fLn2sBT+C
hNzCJi+7RkamoFoqacwikBGIfFjXvNS9485RZ6nYrSVCrGJqE4I9rC3ye5myn8gnk9ImpLB9RBDu
pdKYuxBIR7+MkbxOg1fJ1ZxHK87nEVbSAu+I9f9PUzs/VUsNVlWjQPcc04H8N6ThEjWtywk2BtlJ
Qtz07VrzGFRK7uN5nGoxHZrPQZKf2HPwJxr0uappodt+wkMGE1t/SUUrkl06ALVv/mfzAAOf96xB
vdUYImB1Jx8pcU0Zt9vtLoDrsf7FCUmCKpOiZicWq0hJc/3efYghyGpxVUV9nDp2n+Aama57T5j9
wixaN0kHX6SvAM/mjnniMVapuZIodVyCNXLNBgO3sqwwbhxrZEpGZjMA2wwt4VREHKr4skUYCvS5
wvdLlKguQS5CAscDA83m/qN6PRXT8IOurT5QY9ODL3Sw2aeqYVrly2Y4NFYyNgWcmdOES3YzGh9z
c1D6O/FY/ECg00aSeyGZDsfbhGxbZv3GC3SmoBMibi4Gq3or90lTT6a0GSLb9fPG6uR/fHFDuxHb
XmSIumgeys2T0yCr4LA64zwTn+O6CI3OUFKto26i/bY8G3NBjF0doE2qSDMySODJM4dzpxEEjq31
+//1CcNK1kUOnvxTXhTB6/F+ZMLVNCxVed0jwxBsATt/hevp2qIsce8yewd0zyi3QPMOh+SdQTrr
waug9dcypS+wmPiC9/PQiQ9bzHAEhU8sse+fTEuqCDYZibQPvdAngOw22thxo5ITrumTTCR4A0BH
SRT4H4BheiAjJ6ZyTStX2mqBLQ2WlJqWAODNTytjQNnyWPkyjCUo5HG6jS3YKKMMqq5YS1Q5Lop6
sN1Q9c4gWu4ADa3RGkKQtZR0fb2gtSoJ8LXIGTriIgad8zQsJ7xbv8Moy9NwBRczRmdy2FmokL8l
JUqOixZvgn4/mdEp5fha7MyZAs95r/r/ONBNMPP9awkiL3pSxLsgHqiLJmJBo0BCXTjdplX/zyBS
kr7mrD0p140++e/l4W2QJxLiAuzpyS8NQyVZL1uPdURQM+dy9YYa10lhNpSuBHbWPZGOJUhkw/O0
z5lOoCkUtjDKOzjTDV+suVi03jjdNIvDeuXw4Kuzevt2WqOyXYREUlLl0HLx3rxx+Y7eW66wEUW5
qjhoxWgrvbx1yYKJED2667lxhRAVQE0FFp1fyVpqL7QVxbQPndF8BLPqtUrKtQOHVODP88QN6c+p
nERKrcuoqDMuv0R73hdPqrKgPAVwygFFZQzW8VD/bW71ytu5Fft4PF6roqBehsS4jHNm9tJAxBWm
Ep+xL9Z65PfkIQPPHvtMcBVBLkCKck7aLmFVir7auk389gP179NJmUKsuUG8cVgU+TC528MNZEet
0YtlqSBFCodv2baTBISb3L+zcqB8EBFWvgi/YVOcI5XXPvqpe2Rz5ADU8Jq1/ZBoXHPP96eimFKC
fOe9z6deZfm6HIquSFQT10uA4cH0VGXwcuCAO4BkjdDGuKmfbAC+fAKmUwdpTQFH2bXZzbpCA4Ue
jyc/VOWjIxpitHaU560OO11hIWlOBPRdQzXbr7XO3UO593FJQC2m0k1PLdIE+D/UN2VQxZ7EUpB8
mYYEOm/2JJewiR2sWFlZOqwXzUFyJ1Qv9nE/1TTIoolkErf9if6Q9PbWP9thdlMuS+hHZK2NvKJV
qr1wGlAuLfeOBnAwsQ+nFlJ1uPT0mOP1ROtRpah1ZvlbwvR/RPt2HHTHS/LxpiRYSkrFR4Ja9KYT
EVKoYbzREW8El2QLuhS8WAxTCtF5pMsEVOcz38gjUPN9t+KMou6E5aKTMGkPbE9IjBva1Zx0d6Bi
TIbyfVsjb33XQwOBhe8zmvL+iu7N6aWVZYZOtcNb+uRS44sA1POyv/Q3eDgQ4VEy/HwESbMVY3Zf
143l8HQom6zqKpSQH/sODZnbHWxhTfcdp1Gmi4lxb2HgYg8jKgLE+Bde1IZ4/P/2m1Lxex1HC5RH
jH6s61zWKj8Awe0HkM2d13YoVHDOZEEz0eN96eMf0RFqE1yLDs/ibiIKiABN9eQcQFX5sHcjR+ed
8R3jxzUmbM1uFwxlg3oKY9YsUh17Xp47m07TIch3kNHTV0r13q7xaMQ516oDQ9rMvUmDRH64kZUi
o+QvtnAmaHB261i2WaZ97CAoyk3dCRuJEnt0hJlTBpI47magIk3RQv696s9ub4ofIp+fyl5K0QuG
ronrtqzAbNrhRw9xzLaOUzYl9vPW5S3/rSwXQaoVUg3YxNCxEC4IGCerflQoMtytrojG62GG7PUy
5JjwuL6LfF9FGu8PTTKFyTicz1Ed8XiHGs9Y6ZHusNsAtvN6kZzbrhaMURvF/vGlvYovylF3ChJ1
lGslI3ExemLNDvrTKsPwBoGG4LQBrm7Rah1P+d86pm1RR8F/npcKdY1T6pH60/bmlfzZcnwHJyFr
QrdspMYa00p9vYI6rIHN8ELuDZxjSG7vHR+TMVYajwA23+YqRKSKx0vJu5vhBJbhhlKup1S6aXzI
5P/AxNfNYuSEcwxyA3MItDFXeSBuOQITNfBfdW/2Z1ZkeQHSeSe+yjI7tTzDL9t+cU+z/80mJaYa
MoZ+GMoWYi1mjCunLdrjOc4Ni6Tv+YdPCi/W1RrD5gaET5n9D8WUyv+xitagCUtEnOYoERamWdIU
5b3YbnE53I/OGVr16iRrQGcTVQVuPIBzicgGjcoNf8JLTGYKAkQ4g79WaOditoeLWJRVhxyIPuwW
JD3rB1eEH/sCeAYNs5TfHToMMKGy9dC4Tr+m2n2dA5Y8hin3z18AhHlCQuwtLGUYDyPF3oO9EWES
66nTMXCwa//OpiyJs6hEB8Dbp4qTk1K5O6kmGDUGjDslfeS8uEcaJLVxKgYdq/XGliSmusFhvTMf
RpZnOzlNYn/OPng6Vadgmruw/RXFLdAcZRTB3j6Bx1B3HnQtTDb+3zxuMW0G17yATg6zEQlM/Zdu
M2TldZ4yoGK/ONQCM8sNRckLeqD49ebN/LsSXkC5JBRFzX3ovJjZTkZhkrYMDwxP9RSM6w8fd67d
K78rALycs+Av+edeubeJ8xBF5+13tDLL/fwrKuNU+sENvx/5QX3BRJjVh+uR2ACdOEIMEsmhWKY5
W0H5k/ykPjF0hAwSKjJZ8l1clAF/ar9D4cRojMfmIsKVG3kElOow1eB1Fi/LQ9QDEH+YEtT1ft0N
dt+rTCYlbPTeKpsr2MEWIWjreFSJxoulcuff01ualzgx7V9eFJc3i8m5YxRJwqgCgd583cWrL0im
DyTU26SfKK6f1O77RObE84RfX7V3Vbi+95PvYhaK9fAH7ZJksLCDfBB7PXapYytGTuHrIH93QzyY
Lb03Qev0jMxnjvjHrQGZm5lrzw7HHfvb2eTop6/Uq9w6Mub44aOst2aWZOD3DKu1DKsLUbhgMCqW
5qO8j0PocYnEniLTaVmoLlbadtYIs3VueT/2GpUSQZw2BrXxPt4DgT7a8HBpMdIT0wuVBd46lsFb
kDiJTshgTd/jSxdkVbhUnNxlc7aglQpBv4EFOKIkPlHShCcxgokU6u1OWA1HPux4u/5v2A8KtoYC
xogkE4y/B2+anPCUxkqYo54uGem09Ds2QTkN2+skESTp5fRs5Qy7t/ARxXPe+aov/iYuue996wO4
/qQ9XOaRQETpNk/YkoCyM2uq+X+nWe5pbN0DVBlt3bmSLqmv+TfhNzWjGAG0pFUxMzyHKjU8t5aY
dPRFpm0kizXyMwBXqZfgzFdwqww/DBFp/EgbqU3dwpDo+OwEEFbzEOjqPTNPOOtxxUQVwNDQlvyX
XXUJbkB69x64ptZTL4JZABJCcEm9rFSPWG35pqXdeh2HlAqpDwRw67DojTi+AKG4xDBc2w76g7HA
ep99dMG0qogCwZBYMB4wZEj0li3WwrsGWr1aXSI5H9/dYaqxgPhEbtoiUyV7DP/h68ELWemm6/07
q3p952XdFW0TruBxoIe0rer5/q8HGQ7JQhJKwIx3F0mpAEkGsGHw7mqC5VueIqirfAuAoVGSO/AC
940Cw0DONS4OrQowOEnCVJ2h26QMPbgjof2J/3fB9QYvF7aexGybw5AXqjMA3pUY18VrDEZPCiHO
ecbioZ07XA0ZQP+dxK0U/VhvucdVZf8BdfqUeVZfN1SBwlEWerJKM5VAqrgGYH88WDQe5spSOIIE
a+tcniLipbTQyTX+ixoBqWQRs+2C3jcvRn7sGmkAsA1SnOHq5wVJbSxCROM+bXcOMW9o5JYvj7+i
yZ8SeE7TPh9Not0toGyk61ZYlbHP7TIkzpVP8r+8IG/TuRjREryf862BZlsMvl2AK2HrvscMvFMn
UU68uIu9Ce7GiyBdsZsASJ2wq8vYE00FOZpv0HkaQ/27UwWK5p3LG1Z7ZHv1HtKRvq/ViozFVlmF
1r77gwPW+MhXkzQ5fbjba31N93in5hiFgZEe3Z817d7Y8p5af1wHByN1UbVbtpv1xcDVwD4BNRnR
7UZ7ZMRs8ym1GX7DV/iFe5M/D5pS/2SeWF6NnbQKb3IrTnhd856mlriQ8Zc0ftEuOAej3XyThe6p
5Nx6HqiduES/MVNfPxkK77MLsSRFw6ADI00zAUXe5L7z17ZyeGgHxiY6Vmx10wkA6r/scdU1nN+X
4F/1LQ8cTx2Okdkch1nKW6KU9y2qaJidejpUF+RqX/xVO7vOyjvEqPD/csTtDtVqoHMOEo/NqAIw
H7xTwTxFrCjXv5e25nuuZcUu5fNi/EL4Ua6HVLjZMUDscPGb/TmZCcLJz6CF3eUbZH3RNO7KQ6a4
RS9/HEkpxEW/wFdaJpQzy62USEngsySerXcjVX1jhZURmO6pNrWENKDE2w+dJtHrqXdW9qdFmx5i
2e2MqJzM3RwApe/UulJTnFDsjn/sCBgDtUTeDFrAMhUPryQ8+sGf+ybJqLo4sfhShWN1GbnWRAbF
2eStNwkEa5peSsQy6nb6BoJgwB576hvwYek+UdpfLS4f4q8cQcbQ/ysUdd+GuTFfU9x2rlr2jxXR
/N/1kIOcHv8RfAx34cm3/Fwluwm2F8nmm54JllEAgMnEpYil+kBIU6PFX95VvmGWG7nPSRXPe8AY
MU13XTNgbnRRqZXIuOAAPL0dM4vXvMQXZLLwOEpPGwUio2xLZEW4uFHYEom4iFwbKQJn0W5Qcgsw
xIwAx2eFkUzYrLF4osuBJqXbfoZL6pD2War0h+JBSkGjRLir/kwC579fHv1AV9C/Vjzuz3tRc31e
DGPwwoug1Zrh+9tMuJTdF7hK91oLcD+FcQn0Wc1LFILkK/wZMZhynli47WpHwy8szfyIVEbV33H1
NpwOXBhcqcwf/dRmksGNaUFcW+72WRrS2pbDn5GvVtIwHZtV9JA7VWpI2OeVk99gsfVuY1TtJdOX
BHMqRpMoZI97uisvV0l9zppOq5eMkfDeUdajhr1LfRj01DbPZQm1Ax+TCBXhLFWLr0PNqcMA8zcd
D38jss79xRseUm048HyWvBblP2qeMFYzGkEP1T3JqcplzBdHTWmYDEKPN67JvnTpvpvSsFt677pa
GkORvQWh7uoWprv1DxjAeR4WBSMVvd19SEWUv4Jip8C0iIXTkDcZzJFgXM0d5L7h6sGu7+oksgbz
8bDw5YtKIIZU5AliWiI+wUpCMjmCm1n8V7rXwk2VYrO1DQ8JtlCzTVWpG5us9YBXFH2rZm74pBbk
3IbWu7lTHiH2taMMyewIfu26MtYXnYzmthbZJufJlTxvNiCnxAGI/s+QiSiWW++/GqjaVsf3hkTb
eQZb+6ituANp0U5rME9R60o5XmwZ1vIvPa+KSits4/nWhkgGdPPhELV8rnrQg8NaSW7wwShMmv0K
/JgdCKG+GODBXb+/4/PWSKzb2Z/IoVUHfMRIg5aDWUKndshOFpUlRUSAsnfqDg40yP2KKPWt8TUS
WfH5N5LIHb+fqUDKZj9azzutxhLF6apgKoQkygaXIjtfo3qhtCvAWMCJC6FIo6mFZJV6l1mmWbUv
RNGGJyQEdrsrLOfd3xaC8IQ4/XzosuGcBW1WJkXqecHdwroYRzZO3otBHa4o6Wirg9D7OZRosh9h
AgArq8WWwT4UMBBUiYSvLt1vp1EgTVpdqFrDOIWpJDi6Mho2nq48YV9mxG6xfFbYhuvxqeLBNZTc
bsyrwSHad1A9vRAcGAW9cvU8jpupQjeHKq1JDTbuwRqRR1rVonTdelt46PfCj2YigXmdOBG3G7NE
KBq9nJe4AkMY4OVKBGzNz8Ma6F+oHF8Pukqu1fl35T9MWPSDk0I0a/PfuI/sTao1eLFJucr/o1f0
hYA6jD97ykRv+rwf0/oz2P/CKzSM0cMeDgMu6fFcSVhTSnugdd+S9JCu8kUbqrsboZ2dlvlyq/z+
6l/1Dd1tIH0wH+QwWzL4q01BoMET9NFZHBO7ZGOXF8PRIiDTQMMkGd7DJ0sH7Q2RDScfr8qh3Jeb
iCRI/9+4fzkVgtBbKKlqONiQUw+FbBTmc746MA6MTt4WAIVQK+gmyMmHhJzjgmdc/M4X6qu8SvRe
IOqDDyLaTYhGG4wmlkQMMsgU11uqvJPoqqAUfES6ZOaGr5FY1iRftocQdcr6U4XlysHQHvj4abqN
VzDxWQkyqDS++OsqGMvO0HYszWHYquwSdAz/LzIdg7vLKUF4ks7Zy1FUu0HFaRnX2M9Sz+uCuLzM
nzDjpGQzRaW6GprupBP43aLKT3LNmGO08sQAsx4JAwzcytZuOJnt+nbmMG8TaAid+Xq4EOGA9nUa
bvTWLJjbLgC3BAbZ77kvTsvn+6Lvkj4kH+Cbds4QCO/0UhORBi8ixSZMfDHBqRx6N4wILeIsjAHC
FthT8+l3sR9qB1b4JKeel1++SZwAPxzT1Bet3dSsbJGaFHgE74qvZr77DNZhlPMKhilXl2VDKGoB
uiMjujFWNaIq4nSjX8kgRoTZkuVZOldHcwAmjgzo9Gr4pO4HDt1y8Gyg1eO78NG0zMijjaiNZDJL
u2yN4qqYdbGTl1xWMh2X/G3Cv+XILS2g9EYjdcVfYkDH9xZUIFc1OklMPZD7haBetwLTJ+yz8ZZJ
6Rb8Ypfja+XFP/32uSSJ29yhQoM1Kd4uJnpZE4n8NXr0w9HEcN295D4WYc6qVQnk+0YT21MJVPxx
4eFuAZ10oQuLYVDXvdSocYfq21hHVML0Mna8K95J5Div08QzlF50aU4WxvqmeiyLEFM/izP3D3iI
VEdjB0ABZPJdE41fD3nfjm6+lIr1ahqjAZdO9jHkBg8kMobcTcn414Dq2H4dxhRUUn+a2eQpQ46E
NrYr1EeRNTKqAsD27uLKQ/49J+KzukGFOHRAtob8ZfB/yQLTC+PMmGAcLYcOgTnzqVbe75oWtgHT
TfaFFnPdFI1bOu8UlqrHRVz0PH1TFo1NbV8FUAMDYQvl2Mpj0yRoZaVtuyE2nymxX7aGenkoDjmB
fb/RDWUoJXcufyrG8wBTtbh2X26Lqb04lhWUspJWOip7wuJ0KvGxDtJ/AUeMTEJvmHFz85NhQ4Xo
aDkU4CU2lEcrM0rjBUWJ9oIvliPW2Jsv51cEOjzENfdOQ6b1HSdBm6qdbzB9zIG+04frWssiJEdI
ZO7/KQgtWLF3jj4twovnBPlpAzQdQstoadiHWoDlFGK2sNBMpARAA3Fbj2ChbeOWJ34xFe20f4Sj
EmkX6yRwrF1woxknKwlvPpcDm+09ScVP2cVgirt7dppq8GjgVaKFaOWs1drmAPP2ekqajmZOqvAp
IRfzIwhCpb0VlgMBRf31qUk1W34FhPJ9yQ2O08oPiA1XazMYLTe9bVeHe1FQNLiuC/+KF/wzbIjl
7mAAOqQeFySQIM4aVFvl45f5tvSeKk8Gf4lZF1deteHbuoXNbTAXBn2UdfBmCfHGAVo/nxNyPi0p
yhoNWmBHtubYaAbjq7SSUhtiCYXWZXpFk8sUmpfxvjOWCApqE9Z/FvUkF5z1DGGJmklMEGX86Dh5
vzw1lMD9fUXojJiR+NYONNcWmoT6+ahoMB2RywEjWAYzwIqF+Q0f6lLrU/rVl1sMZZnxEMrQfB5i
qahSeKevNi3tXK5UP+vGQ6Isy1bNlAGC8tApvv9eznOX+popWnGP1bMu+6wuqxMzrjxdZoUN8wc/
/Wls5LOWmnPlTMugm9AMv0k1FayDRUJEZmNTiiCDIPbWcXavFrGVKnyuXH+7azNk9/Dtk7g058gy
l7NZlzAPxY/j0Y6NGUA4Flm9tQUZuaParIBKoRUpxDrdgdxp642ooisCbUeIkG/w6JyveYNV/XLi
qI4Py/hsdLKIJXgkV2uwd+El5lfbwGu1vZu78KpnwMxX7duxY1oEkvoi7x7J3GEPpUdxrJsu/2c/
ZVFCDTHEvsbbZmuCEbCDfSIzsbrhuj9Zi9N0rCHLkVBi95VFcgulYgwK8NnM9kRa6QAt5kQXG4Ne
GKItcQfjWlaVGDgomuN6hJ0CEXVQHtYbtohotuXcW78sHc7LjsBZWzgRjCUOhZuYZXTaRJ46pArJ
h613I9qmahdE4lGAy4AiSfwBj+tdTMq3faGPzsDJLy+vPWUrqvoY5jJsV5uxtOxg6Qe+4RunaZch
HDyN4kJY56v5Scbexa7wtQniEiTnLvKDihuFwxvId//5/LdbtgAOjkGuDR8h+DdjhToH7D/1/uu5
KPbx5Pw2pkMQ3NyI8OfufvXQk+aY8stz6PrV7cnkdirCloS5jNG+ATAiHc6D48o13vv29nz92GeX
m5wcUhPFQgfHkgPXH0NbmQlvC5HtoCtHRxyB+mzaMS5CsSJeValHII+K5xhv5QlQULeyTTjr0t2H
uneTmJa3aJzzTqHYM23ahh59g5QvLAQ5InwRY7OQybtpi3UgpFr5YuhbViT6f04Ah+h+8IcTn5vz
VXiNlSch4utbSokhR35xbqd85Z9ZxEKy393CDzPn6V0C/MquRw7pUbCtFbmOjz/ND7yC3uZLsXuI
tS7NdlnomRk8HFCMXFVnBJEcc1QW6wiq7OngpVv2EccV/88YfpMM+oRy8na9KOhrVlkcam9IbGtU
IO3SAKMDzRtlgk5Lr6xEkvu4joD10Sifn7QgvdAZRRGwOs+MPi/lDFLSy7wI46Dt5UGkoebsBDWf
24rR1vkE4C3JFJ5gzNkkMV68JIb6sZhYtifYh8dI8I2P/G706/Pme20kOnFzBK/8IhQP8sVHpXsE
tszwX5jQuSwD43qWUhc16VSDwybrEbw8r4cTnxKpv4jbxEf9YKfOJUm3iqGu++6E8/Tv1c/s2MQ8
bpbdRB8WaAX+vYhL4pK9DoJD2R4qecJynF/nj4eWQVFTQcHOUVLSoBn+h/wbp9vGPzzeE3ptEoUQ
kq2Ha9YD4V35+wbvyh5LFd8ALaGR1DpckbrkNBqfqHK4vFq/l+FbOzGsCsm+mdM+5Za+gPWtUySc
Z7n2WfEF01Qxsy9AHR7rkWNipgD5VD/RXX2tZwY/P8lilPPSAXMVGyF+0AW9gQX4bQg/MxVRdrGN
qUIy+8Gxj0igVL6nMNZepylIVzOd5VAcTjL8ZvGuR56x9lFr9jDDa4j8z0OW7ruro0qarBD+YgNn
qB+/uSWLF7qtDLHJSlusMiNkNuu9FojNbT85lT+JLopwsZOENJUC/7MHwwr4EQR29b7hVpWxP7I/
sLcwNscs3n/z4gBQa2FQZGJbSisPXnOXplnvY8CqvzuFBFBvI4btU9FfF6BylhRSz4NUlwuz7/jh
lOYYeLUCikeAp6bhti07AtdfngSCv5N6lRQudToop94ZnvW0TQkzdb0sQgTdso6DqLhdfcc/L5bi
sMx0EubQU4jSLoxEJP0RkaJVqi7EqMy/6gdp0fMr1ERzA7irMRH73QIddwOiJoWWQhncVzDKO91u
GxGtBU61ZP1QvXVrsGnvj+YMohDXgkrUdXgswG7dyOAQRxM4UzgMv2owmg06+M92ce/9rwfU6mF+
TygByiWqfqRGnV2ELn9N9r8AnLQ02r7pBsZgFnvxtgmyNuAHux1KSmPuPwJD4jGuKC+pfN1eIlEU
We2ogZQ5gYXDOEprC/2dC79eEHVRPiEgdxyKIqj2vw8Tk69MvzGrvhxE/ZjMTPYGAXYSiMNNLjWo
pi6hqk4XyNGHNQwlJEBLezN+a8zzFvvyrXp1Jbpo/5jjda1aAMnybmNMB2Qi5JVCk1jVUwkQJdHG
rI55268/AwvVDWG2fYYfyQ1WpE62wV9FlrUWOD4214J6dqxt3bVR/9VbAelKmOncnEjqxcTgbvgk
ZHYlp6AhFepU5AmqobSImUBSgVaPfk5oTU1KhbONPaQDypXSDq2iQvRNg/sh6PCoAV4px1BHKS54
z/Irr1tT4ymzBiOwdwOQg3yGamAZQvyWbF5zrZBuno0tuAx0PBw9IRcBvAF1rHsdmJERDtaHxn56
79bqZl4RmbsT1ZLBmG9QhdQjS+6jZSZ6jXqz7hByISi53+BRtxS6gKs2J7MtE2gj0yMmiQQMmrhD
06G0xq3k3t0ILYbdnGjFgdGo4G4yJAzHoLWWugGoJWp85ingzHpAgKg9T7m/bHD9aAZ4dnEQ4sBg
Ize3mMIuUqXr96V0Qp0bb6vMF0aDH96HBnm/3t3NJutvqIfTzFxhl/nv3ouvWdXPrqAP+voVYIBO
WQ7P26uak/WP9GoxgJklYqvHKD0t2o82fqAMfvnjQPVfeK1KZjilutA/zvbA2yklv5sdNnr0WK8D
DDkI4YKqLDhCaFWebSVT8NS84OmP5UeGd7rEGNcAQ1PeaxSiUavbX5hlfL/pVgrmSekf8qx4Ievf
14gcOz0NyShRBL9oL2sr/87CKT1/Qq2Hr1q5/Ld0p9SMm0u+getG3/DW8Psf8wIuqvGZxyaKHzNA
r+uQPWD4yaqVVlvfPQ4SQ94/2HuF8S4sjhiq70VERPj1C/p4RrE+Pl5deWiSrmyT0d5PPUGZd2WN
oCP1R74UXVK0KbXuJYyFqoi5Lzst9CvCBSXgErFOIzAwO0xx2JvMrsdyps07q3IoHtIj6pVX3Ye8
RITDW+JFbRUIiWJV5fSZjdZ9OO9WyrHzOghBUFhvMopScBYm7ZPhau1LnGyTtbGy7PIIzJ3ceTkD
sLW6T2udRDmMefEqWV3B6m5o2lEBZNrQSsI8ciLewQGM1NZyE8dI3C03sRJYCFe59nua9db7BoDR
UQy6w7QTcnmqy6h5UALGoPA5hu5pzEuN5al8GljMyxdBnDBApNTyooImC9AkXSuBaHjiw5LlvMDJ
G4THJ8/0rte5fVlR/qeeGP/+en220pTBb5ObV13hCqxtKN0+paOR9+AAyQvOqkPBbJBeT1ozicIg
5/I6aDz5rkFX6o3FMu1hxWOTzV+bHk0mbMYZVglj8ie29fo7AiTbsAuxhx5tE810bDl9meLFxPwk
dAZ/t5xF8kcwkfBWErUyPNhhJvZZfKRlENZxyG6cRBRJFCHC1m90UMxi/p6lKe19dpm6F8pylkod
KP7cDOggoi+wjxUIzkVHRHk9eGW444/qF2YPy2b8CF9z0ct0psIvLCzC91w1RzXmLVOhBCGML/xx
WzrLIkDnpX5N0gDH6HXF3i4hnFXh+eFnHCwM6grk7q3xUcB8gKOxu0CnaBudzuwLLxAJuZvgigtv
fr4+IS/PJHiXOUDexGvhHh3yHalpnZni+1im5E5vF6QbjFKbTSjjixMNsuvjzmw1cYDv0Zw9UB0g
MWT1/IRXQlgasyWTK2feNxzmSilJRbMFfAyHkqfhWu6vcCBpu6cx15tauu6yCGw1Nto1aKnRfGcw
hXaSQNCGAwzZLWuVEvReWeQ9GRlYMd89AWRn7uYSHGdvJ4qcGoMlt1eo0o8Fr0XvufPQ1VxRKH5s
kKhU/OLR1OVnT5bt4qUh9WaCdYyveXFScqbuopTTPLd1wfhAjLrlVoHqFe002O6zzFvR/lIk1Ur+
0SQRTbLV13OFrP7LV7EadZ72gfcyVCeml0/n2J5sY0Ligiv5Lzsh91sGIeuPFGiBVO+dTkzb8LZQ
wx/jiJiYYGK9odQ+5yz6PxhFJ7cU7fVWdETYSwFbVKj1afNaEl+G6pBhwotauA2HYkUdG0bzD/by
7jIg57viMp4P9iqQzfSHzJIJoHCR11V188sC1uG/zj/hJF1UwfLdtYBTTZYiBSh0rHtFeRWHHE/h
Mb2VkROEV8SU33DPcjzOC1QBTRxZwbHBZQqQF0olxz5bfoMsVYtGrWFKQDn8USK6g1L4XcqlSYUK
p5Sk9zNhDUMGaGyskgrMDYNHllVOPZlq3LBBQ74Bt2xydlFGwD4JhN4HVfdkrqzZ50/25NLGLE7P
Q0k16IU6iAuvB92i+jt/35wSunaNoKwO46h8xGrrmB0gruX18I+V7tKsl0ZrarD7OEhQojvo9YcA
UEYTYiWsFmANb/TV+1yy9+UgYuffifmBUSOhtu9VJoX/KY78Tc++PYNdwSxI6H9FxyEHy9FWI/qb
GLAsxrWkTsXgvO+2QrLkBJY9w4qoJ5F+IFktzJFkFOGWsNb66LOya5Al11JRS4PkOR/24pIpG0Zi
FhKUKseagHB25LdhQygyNcVF6iDuYnAc5xfcLPo1R4/S03KhvRvyuP3JuJsL82DxNf4fxl6F8zc7
YHbgHd7003ucWRi4eWviWG3p3MbciCNb3xpqcUqEq2d2fT9APmCBbq1eWy77kZcYP451gE2cfWjm
r1boC4k581dz3yxIUOAlK/GtfEZ0Qn3IF1pjvxc1QLd3HTQjouaxw/4wi+X4e6ChH8lCm0wSNNdK
TMrQUldvILyTjTOvGOYzCN/qKslEVHHGJ/t02xDE8Qdq5EJ2OP78dQr0jT56nMIADyVwrT/ZFFiL
hnbTIL2L/4boSZyvf5M1M7cZDnCtKvp79cG+kwZc6V+DWhIJ/hfCRvJcRonDgwFyZHkHMIMofr/f
aWjkkJgLQJ50LOlUhurP3vWH+Retd3PYaTSQKLHNEXtAWLRxtvWRah37HfR1Oi0W41Bqgnf34Wkg
2nrXpbThnHlcrgFtXE2bwZVGTyNftN7S9zJGP4F9hduXs5P86lQtkQIHaCEKkUFFSAnnF/OFtX1Y
HM84fq305guUpRN3Ocb84jo702MVXzUDM1RzB2tl3hf8BZUg1zSsaTxQShWmqnsAx7nxr5Ydca7O
4SfBYwCMlxCPOwUaynVisYvnqBBQ2amdIJr/sKEz6MShh05LZ2whA/tp1S5HbOjXey9Tr3YEs9AJ
5O7Wj7zySBG3BB1eyq9r5hB3etr75CbPM1Bd4pb20YdkYJvAl/J1ZA61I40SVD7k5O+BYZfq/yfx
uewUjaJtyMbfb7LRfYhLiH8/dDsslsooBJofTBkOPthQdDY/KQm8rNd/LznDa1TAAKKqt1pecKlC
/yK3geWR5b18BqlaLr+JaHVEG/5QH4HP6YcbmMGJ7faxUmGjdzjGGmsW1idgU8YkAndzbLeyKL+f
Y9r/IfKYZn6AzCmn+Am1Y6l+fYTlUb6WFAmYnAhRL+NMw1+Wh5D/6NiwM34ALTRMMZInstBMCtuo
U+GnQtUTG2yZOvZ3jJZlFJPThWCBBrXyVX4yZlmqAdG7rKu/7Pk3fZGWtYTy8KcSrT09vuc9fo5D
M4kUN3GC7l0KVKYzy4Gei23QUw37/TEdfQjepAYnfqoxGw8hjqmxspbP/EQIsDHR1jUChUilt9uT
tRkPem9EAoWN9efguBTI1V6k8CQ4oF9od/U5ApnqIewhj0qPQvoDYZfFB+p5zjUH2zKkmT3pXqM1
ewIvRWMUqXauHUgyziJJAYlLaac0ekjVOWuTmFm40CRT8IBdNAhx+03KFTJxrtDeLq1UD5k8e32l
LKeyk28xlJncHIzRbUe276jqtu3jmZBs7Z1coomph4Hkqz5mc9FqPb3v/Cv2r+mcm6/2m/yXO1+I
aN5FpGbKNC+VOxJ1/ohzE4Bt0X+VqzxvGzQfOB9Szov5+tYchRsisoZn0YPokxKjQ11oPgIN22Y1
nn6PbhilLusY14N4LNq1/s/cwD4D6UwyFCzfiAznS1YbSYdkN+vFzAAIIA3M9ENmqScEV3JOqsJy
h1EZJZw1uuvTco3CV24aYAGaoifwgFF5fr154JVI2hE5jxBCoxAfr0dBmx70qUtydxgoBz1MF4mo
XawQeil2AG+H9d68gw7wKvr7xZkcjUIT7V/q7UboJ86vRZ20cbN9HDgwZyJefg/Mn+MHTSpo18Ri
sl7ciEWQx00DSYl+2dq6XgqwqXGemvgQSouckeYM2tbEHMVZRJH45sxOu9chNhv6VunwEVRxZfa8
oiYrVpM1QbxlH7Z/GVA/ISi0hySu71NzCTfWSKTxYWGC2Q6NfoVuMspeKJqVC3RGtcjUdmi5q/B3
dRwZoJVRuAzWukOl6ElSToF1qlRm7GBVIa7CPfEE0CI3YhrXvbGphFlE2sGJoZpP23v9pwrNS6Gb
KnoBoosM3GF92uwAai8iZgbfO9QzwxJYGjdOeD6TSrdX7cebUdpc4aadzIYkmK+JWmllaW5czj9T
Q3A1aLUeCOuqSQu0HZtAaqPkCGUcaq2wnMHEd/e7FJvq8IZDU/qvK4lZRon8Lnff7jFS8bXnEM9C
5E58Zb/bCet6jbujmB2YTpLjapa1Vu/1tKGIJT7+AnF+Vrrnq2q5gCy6OjKWSykY/V0PJSUcZR9J
waR40NufVRPmINbQnmvJL4hkNezb3oQGjjTDPtLmcrOCgW+fgs7Kgnfj/Vsy+eXL1UXSMg+OQm6y
NGKnJe8vBvBDtGYBE8raZj3P/B80jpRDQN5OPLIsStQi5flM/zHBArynkNEQbk/N8hwV2dWI8fiB
GP7XiyRjZ2eVSTqent/xBm19SwVi2WMHu5a4yPgD6TifKRSMzok/b8H4yQ+euDS1990bkTIbewlg
4rlhTkzZqzUepE6kydbIVsH5ibMkD2CrnUZJ96+TIuE8U1qu1xxqjzcUhWzumvYPfsF8BnGWNEaH
SPtJpfxJMfAAOUK3zIg2uUo2DocAywpxgCuzyTBx4pMZZ/bBCLb0tAPnLmiToaCaXtEKe8/kLjk1
Cu5XBZHQGsPlEldZBnaUvYx0uqWnZpymlEziUktIwRGyKFPQ8Z7FuE9naVsFcoliLrAkUSQ5w9KZ
CVcNE+HCJCUSwJaZnHQur5+y+VmSEvaC77EEqdFR5XcCgOD3RSGvqi+LyVE9CxehmXdM/w9CaFdi
t9PR54Tv+wwMLmI3+Ya+GfzfRdPz4kCmvROq6hx8UeQrkkKsbwni5qsgITuEXUjXEOI2sxG6IVAC
uAaeXjAhid+mmhOGJW5p0UcJg07m0K/Ydj3/swx2BWDKWnNbG3LN/S6aghua18X6XrAUWv4AIKpB
MSNQpo81nbfXxBiyOOL/lD8bjhE89uNJEZSU1gr5ZRQaNm3jTJFLQCIVtXOEnkkY9QWkt+TKHWMq
S4xYyxR5YvIWXmMFmD9V7+EosPlsiqRJ1L8ryQPCe36yp9WuFM40Xn+QavZMINxmnr6m8o1zjhyg
UkhJ9EXC5me8t/LV4iXhseUVAvUYH4zyZ4Mked1WFKbk8w1ya/KlPxummoO8i3JvevNjP/71Iz30
lcTQr4U29Ht0B7s/gmt7mFzuHWxqUukH+pRryv28pY2FqUUZWI/jqyrTLcpksqVB84rX1v97PhIr
7Zc5KpGxVzVaBIxGul96i23RrlVQ0MVj9z1wezzbNp33IPXPU8Wn68vonE35EO8B+AObrZp7MVvf
WiCZ37ODZnrpanwUr+d8qzScAIj4NcwQ68AYJn0/Nk7P/Gws99+tyA2+Rd4sMIQYx03O8/kI1ieU
dbwo8B1c6SyGxv6IVA9Ponw4ct0DXfl2sk0SKZ3YdW6ncQg91uX5tK4IXnxGO/dmjdItK5G6ZT9Q
39NOGszBNeVPCwe1A64zAtyfaNG6F9j/G6OE2a5wgVq8yTIiPvoG2P0uLnsSKUKuCN5yqb42IcIk
v5ML50tasPtfUME1PTGqafTFSOYBRwMP3UkCvY0Y796pWJdGdtIIWl2t2bwc3jt1mb386QHKqp39
9tCc1Bxe/XZ+a/HB2Z5lf/ndoNTbnjUSYWn6L/SOIkTwAPukVTbQhnMpwceHe7W/PLpjwINp9K5W
Sv5zfauP3nHZeELoxCWBWr28ycMVhvlLWRZFQK3EiF0BoP0Do6PzfOihnnPktdGMOPHBCHeRYDpb
iLU+V8B1gBJHOTFKqkt+6gDreEMbMBiJthq8209d+pXzza3bS3GP0Y2aJvU+aE2hE724t5dlLRBy
+ChWo47dvrGJBlSbnTqGcWh3bEnCqfWYwNCdjDd/RKHE8AkjTiA1qCenTghkr/DuffoSkebf5Eh8
FKo3HrQNEWXUKeOZ8COiQzYEXqWsI9oUsBdETx+0HA2A94hkJ5vsjFjRg+NzpCLl+wTKR6JU/Ngv
LDI8TU7BnUsJRL8196uGiIfyt34YpPXsQU92+PfUs9qGFA10yvPDY1J6fg+gSrnAk0qrzitJEVmf
mCN65QFaf1gRm/Dmu0zsiRhB9XWSTk1cflfTfSLR9BjFEWABalXtGIvahikEwdF4urcEmFtkdVmK
JcB2GvbU0bWbCGWR4aZPZBd7CbuH030BhJfz/9KKiEQm1LCOmohwq+P4Bzrdic3tTphIr5SazvF/
fqJhiDwXRwvcWB9cXkdGWTlyPRQGJG1auIPYW9WA4x80+kXIlkzGYRYLqHtIs2fbSf6/UjUm5E5I
JAXha/SkhrHzVhz/j/zuEZiDqWaqKaT6RpKP+ti028m/v7gqdr0f0JRaitoREADEOkU4g7XBDbSB
1M+iVYtf61liAg/5oueFF7avh+/2DCscpPgetcNqDbDv5JxnZlCYfuq3voQi6ADIXVBE6C+artZX
BNZpRNBmwRY00LGWebA/nXmn3Y2EXREbRtyEFgfsoLZVq2CQfEvf+fYAp8X0XaYuLGzscxemk7ZD
cNAav3mYhpGXq+qM1Z+L5Yq3uKo+tojc8Dpgeq5v5YVDyBoEsSegH2lxoMkM/QHOjISFQyNeuJYe
MQnMUztu3CLdQFd/Bh/3f0xxuZqHFTBGE0/eCqnR3Cc+I0Hj017aYaW66ex+9Xgl8DT/9Pa1TrwR
WWTV5twsEP8enZHSWsj7QOZP/vga0UhGr3ez8sH8yNxcdjO86ReBT63xQJB8wT/xu4ofLedlKwau
4HoNMvTzysnk6V2z2zwEFXcST7ouOUrLLOs9XK2snCpvHtWRaPblFiL+G+YwYLa4ppkl+mwJ52wC
Hd2NoEciIkC2AAI4k+vfol54g0KEVglcEsJcRlr6zwsWPssJC1468mYGbyno1DqylZCl1d71oAuT
HjdQKxELrZ8RG0e/fgQkLwy+ZPwkq3JhDzMtC/JX52YvR19NbckfNtAwGPnmjKkp27qQMpX4kjnk
nObjg3VBeX6oLR9s6hMef+MkPx/cBaaj8rWBjtPfCfISVvWQFSrogmWucGe/q/v1Zmdi+BzkAmzy
hQ9iMWzxg6g+1EbJSWbFuyN8mgUGopLrQ1Pd7WhrNlChWzDJHWXTN8eC5+sJRmbRb5zw3tsuufEr
gUu6mr57ho/tFZ4Mb3j9fHHKuiHXBPP3mq9pX32WXBmCKr/QE1WK43zleQ6fKg8+ozL3lyBkFHK9
yOVwg0VlZTHeI6XWPI/yfen3RVeCFaH4BQy8+2xuaDtoa8keXEZzAMh+PN2pwJsw3BO792f5MfPR
3GQrZltxsCEbRVNE/7Ok0pVCLNJzShlVBnUfrXeLxTjKJXWdRZzURdyAjFVxpzJ65svsCewzneeL
xWkXbMiVLlDkzEGxp/XbzhHWXU2k/jSyoGmgHIHsJkLDhEaSEZelPVdjdLWuExaoDouvTOxUQ70u
6Nl47yx9CTGLDvvWxT8yMPAzeKujeMgBzC7ueGpKPGObCEZyC+ExcAjfsYFvZd42ZhCQsgFrgNmH
ODGhXPDdGDhDe5KUOzZAcOJnDSr2UumzzTh2IJzZugHvxr5M5ltK1C6sPFMiBJleJ+EM6mDAazRe
rTrU42uANvCoX96a16EyoriwluDCUiiFEMlu4SUfzw3m619AqTP65zMFtHAZ9+oMJwrpuzmbF+oO
ACpXSiUl+XC141U7e63BsR7h4gUT+x2yVb/ssrbbPTPvRYO9f8msIev+/02RrSeUwKjGeDCyEWl3
tG+3Qdwdco3wrD5MU4M7zGhBS/jAqNuPXX2TLuY4J0LaD6NWdjPrfOdm3sLXMFIqvF41wBXnrl4B
X9aWpV1x/pd4fHJxKaWv6+YJzLri3Xx7UAuwrxtkUON2cKblvthXcylywLXu6/3b5qVFzYZGh57s
kaYnU933zrlRWwTFwvm15cLzKu8HqJDltBUCFdslN7fcsH5rVb9/7GHp2cHPaovl2+cxXkigJzXO
OSHjp8Vl4DrXdE/IkcL755mjjZFo10u8SkWzsGJacHNEV12bmbxQYUXGWjkPllaKsFiv7sYvYJGG
vRSckESPj5yeOUOrhRlxWhB3e8HwnvGLx60GFyTVVMD7I+GR9EUt8ac0zpAYna62uLXQj0uB+pzs
ycYYUKKFld8hwhbenX33d4X4uniyk8qbJjMXtvNWtGkXDEN74BXrZOAhky0zuBRyLOPKBr7m3HsX
R3lPdwcP8IqhbMEC5Rb0hs4aFWXWKxglW9n3iR/jybIPQQRGPNxrJho7PBEYysPq/4yYPdcN84yG
9h74hsqjQtS02w9/7bYnGRBp/E0SJ1+N1WxhKnq4NoE49oyB0UGkXmfejnUTsGNOFLx+wF+e1W86
J0wCoLt3ApOD4V4Gymdvo36odk+rR4g9Ar4Pvlfu4vU2Ouci05VH95x34t9+vRq4c7zipV/geOTb
sO1Tif8Sci8pl9U1LutUJBmTh2dZrLy1+QRmnu1QvadYM/8l8QyPRa9Ly5TSaVzu2ebICiG1lFAe
yOcjVMaiGym736lTz5VdyuINklFiB9hPW74EQzkhOak/mFheEIbC7Y+sbt71axltS7INvV1o0y+0
MzR7BWcj2WcbHiVnktNqryVpWnP/jC0Nc6ViUgdLJZNmslAaJsm4pGAwvL4PY4DxOqLdEbzw7402
NQi9lwu1Ae9wiZS2t09Ib0wsxGYygBForTbl/TVPvqV3EO1O2vM194a2KbtPawQyCbD68ZM1HAH6
hmE2V17uaNsJL0qd/zA5JVh5368u+PRK8RpC0EUAK4x7IDuoPrfz2dRIGlpo3Gkf34IS+00TZF0x
L1kBdfl49hyzVoUjc9xBmFKL/AF8fp7VeVhvAKELg1JtCs1Ffw/l39GL8peigr4SbxumPQJ4uXQm
GHn4tgRiydUvJRmAzQ1tWSnboJaOv26jCft9HfTMgPokshVvMTpK7VtLrEbV/CM4M+Ocs49eYHvn
2K9gj/8+FObEjxAghAbl7s/8NACU1klUPov5KNiBZvLtqwIwPQBV3VZaYLMOdFD+RZN8mRTs9PKp
E0fOxUR75OOngVwQzzlWA7jWuTBj4kdPZ/Mi20Gfbql4vYU2e9zq8MAUpXsYNwkWdegLWm2Ha6mC
FRQ1XXmEziCJfNXsqkotm24jBzIgY/TurE4xoEx/wbIH8KoNMTeCPZyjDJwlLEFdMHF+kXx39L+M
xG2QPiB45dhBQN0Dt7hku+BaTewOkZubTYqa98LPwTyoJ94hgk6oY7xejrgIUX2/SXcyARdrgOKr
5jbGgF1x6QsZq2x5qHuz01VRUyaDu5Jo890W1HNW418J8zp9a+h09thjq1oAfGF563JxDKxh/k9N
hS0c1cwYPwOqbWYUwSgluct2Ketv+mxhoDI5BwDClTu5OfJ+ewTJhqevAsVAdqcnNfnTsZEzfRDk
PHm4DRSNNbLjh0q2EzCqPk2vhlu+K5K2KM54P9G09NCKQl8/aDyeh4tfe1XTbmAkUIQAg4Jqoahx
lVgDe4Jf+ilQdwPZEUJeErisYS1YNUibv/XsDjFTm7KROYeyx22c5yq/+qXyr2+yShuURCZfii8k
LY51srhB9AWCEn+UWH89HCfenJEpBeTrZrXvRzDfw/Cxa5JSP8jmO0yDTfRv2Fk5cLSoEXiBD3cF
yJaUb8XFhKCKMaPZfpj/IvUPna33X6MM/raXWXzW8Jn//QuJvsxAV2VIHiVNzUNBlpoFtktencN5
KJ+NBz0JZpG7xjOKj8309wpaNcXTxGY3XGf/A05tiqMTgb4QVYTYpyywQtfN0bxBYxF2ghcx8Uw+
ZfZ+SJmrFAkCbmhNR+kWaBHidmFXo9Tg719pINMOc1FFc8PAhR0ucQL6t95z0GQ9leup6OFptmZT
k2yXPbqTFLUKGswHyugnc7Y85SMFIVW+KDyFTzzQIMZXWsAJMXvGA8PVbgmVRAjk+8dEFpQH7cHE
jp+/5hyw9OCifuO8zJ4btrttrU06ZnI/VRfb/h59Sn6/GuIReoRQt+x2SieZkcxWlBoX/X9TZkip
YUR/Ugp3XfwV3qIzFcA5lL5u90/0d2JAfMuy7QaVMpR9nJoInobsjU779ee7fK8G9oV7sRu995u4
dxKP28KuKMGAZvHBsczrPgnjxOxXNA0vpr8TS2UGBXAOTG6wXC/ACP7MzvZCNo193BCPJzcGhm3i
9MyZhhJozbZ+rTPfus15EbDlFQu2+WAGlXWWw+JWdv3Ewjm3lNbuo9rksQdf4wYf3p5JHjYatXT9
Mn1rvMdJLkc/g6tVVsG1UJvzPL1Zauv1FORDA3WnAchGlHkITCpjW3PM7eWjnNYLHWi9Fme39Ogs
KUK1R/fBbVEbIhQJOf6eqJxiHNCVh/3+d5QQwvfxTYvDSatSKn6byMvFcS6ql0AjCBaEyAItbhXs
Joad3c9PE+16dH3Rzoz5SPNX9DVT6U+L7s9ufUmlD6RGx6TLljSmn/E4k9AGIGMP1zg/eT4G+QE1
BWFvZ/moJ1LIRtUjRH4rEW5qbJUg0HP6Rx0yttHwSc/2vGPKdHdgS34OVBwpjueFqIkIjhcou5Ha
wI3K0p3ImWbU3c6TIIuLg4XlDcxEj1icSQL+TpmiO+NhN6xEFYOodARJoS0udGHVoc+RFGMkeIu2
JyAOf9reAkhK+ZAl+mZwwR9C9BkVBa3sO2T+l37dr8h2Tii2fFHI3HsfqIIzdTY82cBSLDQ6dVPF
u+vHaJGh0MjaSkbul5Q3Ctr0IlsAHAz33M/mVNYnUrwsjMu4vCJKS01+tychuNcjjYq3/H/vy0L+
umu22FKJs9xpPpNOVlDvXg9wwx+T41oq+GcuchTEDY2xkhPulANtQOHJIwUur3mJ/8ju+g/tN7P6
mPxcSEqUTNI3BJ9n86MTLTNeUFzogZ+IX7PqoS7J2cxkAGhPmjhl+eWPBPJObHz9J8UWavjlKWlQ
XwHyfDdEmlNeT/bGC6FdEfjjMOiwpXgrYRupDhJROYkPek5yZxs7nJHskQs4pnT+5DVUf1Hoxrjv
wTlPXqIkCJfwU6oobZKRin6f3vAppi1qConFLaieZ6RaC04+LoalAaoE1MoEv9hqOfnzfwcSfHGD
AoOzdJkqlnVx08CwmRh6pBIRN8Qg4tiEcV0Y7E7NzyuUwaARd8xP9G1sPNssfr+Y31zJCdX3y48v
Hnresb5fceFBwHxeD5rbAUB2Lzg4aXhrYBg2uRLw/E1Uz4CvIa30ivhDRddi5/d54ZGBWeygpZ1U
iAFA8kV5naWJRDeI6IaqoZJic38l8EgbXSFQbshi3qpWaFqjZTehEHa+T7bWuHbrvJeV2N2ynXda
KABSKJcU9JptzzrDuEZzu4mYBidqglViQL/E4UROLvg80KwadfE5pIOtW6NP+xZ0VZNN5cR6v5oh
9cZc35bTQj49cjVqYNp0gEehZ801P6mPjvNFT9umpSHwb2fFinsZtrMLPWHGo29IeIWwDRIJ/lHR
Hq7GDOAGO+/siSvevnnZcu2rWzRfH4CczvgD5jTtrjESRx8fwawvZkGy4Zug/bD1TKY/SBYA1adP
w2hoDZmeLVrQQCoMBIgu4PCCaj+7aiaxp9CQpqXKmBIGIw6waHoISfQWpqv1LmmXMH2TsRFXRez/
lZon347NLHY8bHEW3z+TpEn31IBHaZxu5yIE1NiKCsDSj1hIBrWjXylIRxT4HpLVFu0O8fqDrSgX
15Dxxqfxs8fQRwc63CBpOHNIEkHjRwOvIkX70MekbVSoIBWdAsCbvEWj23liIFlcTOFrE/g9c38U
L6qiiIxTDV1Ru6S3/n+4qLdzoTomuEtJBMhS9032UKJa8WKN5NiSvjg91WXLDKhVRe3IX129Wcib
rgimWrpNZ3IcOOs94hxD6UNYvMco9DpkOEEbyQbGQSdqHl1QBzXOOx7DxTMNNQ+oD3LMZ3PacFi8
9gle4Gsao2WUYzO8Vpy6xjg/W/I7C9J/JkyNFW0GN0Uz1jmDxLuR4aVD/RCO2bJA45o63UZXYOh/
s4IydpJ40dVj+5+vKeUhlXivvii8nAvTAuid1eufLnQa/NVstnKpSJCLN3xDip2zNiuXdr2V32Rm
gq14HlWLSQYdDR5DZoOid6X9ObvrIH60bQdzSqz9i7bE0Et3jjit16/vz1XhMHM75ikS5k3PW+B5
GTDX24CwzkIFgdj4CU7Qg2GnQmuoDRUIhthEHa60mCD6Ujb8MILeHAgTjPXEnH7k2lPTpx5w6J8n
GzpUZ1QoSufyBOpIzONtVnHI0mlSGPWnPXcdx5EMKP9hKEA7I2lxa+jr3Tcr51GHb9FPQaQ0Devd
hnR2zrys+k/NBiEz4EftlwH5++9Ea+B36uexyWPO1dHwbCXJ3Jxb681imbAAameLFixPecxFhiad
Q1zdKthjcuI9RLewRIRvxULyhMrhgBMdgWJmAUEudivSfT8YWJTM+5vp/+CTznYMrCyfFeO8v+lp
ap5POK9IGcNUY0dT6sEiJEdbt3CmnMDXpJDdrXJNhvkfpMQ+og02drNncDk43abC3HjHls/ao4WC
2Xppy5fanFjHSPPvfJ3DED+/+WQ5ytw/8emndfdRdOHxxX1ybtPwcEb2/I8M/RKuCE/cND7ySY58
MJHcwNiju8sFDEQ18p3z06GirFeFjilRlFNrXf8W4TU4bU5y60QBjOye8qoqj+jlkA+Jh9Nivq84
ow097CViOYaIg2TO29KeLbrvh44bRPeUMyDdBJGKUvNcjBExxkcpEAi2w1jPPb7zM9n1nx5WWusd
ODM7UeYq6jQaPaNSGCBOUGm2TKbmAWNoJlJKzeKcu/+b1x5chCKLiqtm1kdDE1sLhAxjRzNKObnH
maP/AxGlJ10yCWfwzz6+YmzKpniozQCX5uoWl1XGWD/EjNcYYqCOTlWqitbibVwFP1P99FNDl/3n
5OGmjG6SAyF9jM7sg8uGk6zAcpDcpNK4G9fr1+v0S7o/8+TkclJS6oqhJAHn2fu7/KpB8iBM80cA
KJOX+pCOTAp6xMh3f83y5zA+ERpPE9/hknTQvvKIq6LO9xbKHZ7fy+yUvugpIv1NKv5ZgVeTt0z9
VfMdc/GmkvlNVK/29yDY42a0cI3GTPODE3DPTKmM468NVnI3etCznFCUwcX6bjL2NooI8YfAw6H7
nGwQv7obGubF3OmmsuK2m1FOODnxInG48lWQscSkl+QkUGKnUfwWE8e9gSfKX/IldXvjJ0deX7VT
kE44RjZiYl7TMZQAZ81imngIsfL04YIY/a8o4QAjPcJyGw+uknfTBjZWMJ/paEA96vWmNcv3GFt1
e2/5dYVa9skFCbcVOMo6uz5g/VW4OVi3dMtaX7lnFMeY2bzt3NUC3qpqYKldb8OYtyjekMbaRv9L
R2IFB/5a2lkLLJu9cGLFFOtbQFqDadjZUZB77/v0EM3EsILaj7JdeUiLnwCPyurHHgdAVmfwTowR
2+6JUGFzijI0FSDEtwfS/DejF6C20JJqn0+mprbs7cBP7gi9Q3ara/+a0fwfS90HWlIOiUQEmdEL
ZXIiPEGknzkbMjTNTuEUUcSdVUB1OalMXNjFR52OdBIssUF4H2nSo8rSgeELcsG9XNdnDe2iihMc
w51WTW1w+CxH0U2Aus9BX5JVocVP6HZeGluxbuabEMAorDxejJM7LkIXV4QyfobfKu1Maa8XMfx/
Ltm2k6IEfCRL2qg64faa1hq/tqr5u/0XyKAEaxzExL5rgqe7FY6WQZzrwpQ9weF0AwU9MR5j1CUS
aQJY1oX9dGe1ksYBxeGVdbIA2bpGvnlMJZ0wD0+OdrLFzfz+/yuPyV06m1wqFnnMU0607MJlthfq
AmYGauoj5qIPbi1UW/WxFLWZbiDgm9bmesaLCwDwgWb0GQHsqEEPZU0me5gB0VZYSJ5d3frPqhSb
pExTFKRGg4P4I3EtU068r1sUAH5pVVVN7lBW6zq5DwLwJ5YAhtYqTwIj6zzmgUZmWKY8843DHW/6
RAX5q+tKaq6UOTdojP6fiCot3r65ax3Z7BWQ5OYCF7/+ITlWNitLNXGKw2kqMuc4fGYtUP96csfU
vR1PVDyotTupBW99AGVdTOv68Hbciw5O7P9n4l30gYHkX9742gExO2wC16Sy7gnIkp+ajA3Jjre3
MfLmftVCHduADcE1rBnZM5CeY7yUkxcZJcS/wN9dUHTAe8EXqqheD5x0q28H/MudpVnckwlnYKOM
Iey620B5SzvfIgv94m5SPcLZzS6/yHVyTA0uwRKQ3wXwqXVkCqeyP9ZpafnAwaLfjQgM6DvZuv39
wDU0FNoQyd2AFCi6CDN4EHghf26gmgc+wirc2tNNsHDrThchDgR74MIf31TB2rr9I3oPlM8+vlFD
Rh5La+hHxexJlefH7uCHIpvbKL9f4YkYbLa9t9VUQ4Uz5k72P++Bc7ZaJEwFhReGsWRh+El4tFY6
E47Dpw8iUF1OTnfIG1oTW2tNtLhU90RAQNWsVaiwY9UCJdFtI4Bt7E8C2/qPNsHyw0uxaIOfDr4z
Uod9QMWL9tEinqKB2JFhNGRaIapw8lv8ZBQ9OXXfj8d0TEuytGzhB5CUH8fBlHw4/sVlAtseGcco
uTUKaMkVxituJ4+aO4oTWllsc6iYFipnzdV6jpCCZnxEBoWatVM88oV+m19eNR1Cptxiz5dHRJWc
S/fOOcWFxMdecijs5nF09vMirDcKZ29Bi5aPhBoMXdPIzp4y+oEVGvlri+15cfs0zljF3UQtUI5l
hWmuAlg/UA0b4VzChLSM8wf/GhMbXm9gVJW8FpEwz1GZPzs+bGakApRMBu6WnnOR9DA335KSRSeX
jug+XC/wWmtE+7F/tDt7Vn+AuNn7uSoIgJWaBCHHWEu1wjTp2pPe/wuAA7BIOJam5V4MW7tYSbNp
TH8mb5Nz0NEr6/x8yOaZi7c8zP5FrSioV6cuRMqdk5xjFfxscEhfU/WC8wvqRG/AI95uqRvuGpvP
PV2lMUYGQt1QdcUNsFltUCKM8nnEAfjMMr6hrQpgJO9DqHGAAT08IfV4MnEehi8rEa659/KfT3/K
vEVo64Sz3zXXtDZL3Y27PcVtPMIzBjsNxwwWhDZUx5hlp8ceMubRxrmzga4f17/ypaDD6HTCAz+N
N6K+jiiDQPttwzkSCPiGwBXbCoWJw89GIANp3f2jQ701Qczfe8Ho6K6/+c/ajGYFULMYoaSEs0Yy
asXlh5SlHvBKY6i5XVlNojhxSa+8/Yx7YWtjrZPjU47jqR42y9PBmVZpAFNQ7I4VmSg9KcxiQDrK
R1pGAI1wPZAPcK25ubVGPQkupkn2tm2+lr7NQDsATjfYr7WOvXxY1MQ4xQhmkkOSyAqOZ9AAj5PF
qLsUKGyn4R+5iqpZILR85x/Na/wj1y5/A8/t6Zs6pf005V/UqxsNJnGydlKytcgoAeQkQBZVQiO3
l89UBAO1SkcX7bzFyA6e3evN+kJTAGrZFhuNtSFUYTeoDXuJC+9oQk5HDh9yeVONE7WJPggZdCf8
wiHseXV4qxnbURpdLvhQ834HccaLlmKQZxAOHOO80YoB746DHQq5lQvS2kBohYgcfyxCiWNzcNr/
LxP8nyh075m6nOkA+BkB9wDKUMqckApMur6v8PC7Z5Zj71ezrdnMKrn3vmhrExAXSp8qZbdOC6Rq
N3wY1NonLK0U+uGXBkXOxK5xYrk+swZWJUtW1+j1C1rcqbBlD3uiWTCQL16Kd2snYqmUs19APG7Q
kDXxzx3r6pByOS5BVwUHCBXVrZlcbm5dg0Wr7YBFCpFjllp6h2TQ/vrB24G/y9OptBDlzTbfy/Ba
b2ir3b6Xn1YeV8fT+5nPy4Ql/vM0JetBe0to/fb2HgUExB1HWuSqI7lUbSoKC3OlAIquz6vg5KGR
kgedukg+sWk2rPB5uXkFwaetaKEWO1jvqKqCoe7teIqtYKbAZIJqElH7YK18vM+SxCIHvJU3idkF
T18JTyGh0iClW1FRoRx4BV/LiXjm7Zmc7vRhEImMzOD9lzO6BN9dE68Q8wbL2huTn423iVk1J1rW
QQm4SHJiXJX/TD2LQomZTnnJURg0LAgQxmmnOYvAz+ZqvVMBLEPnWRO20aNd5qlfgSUW7LKnAIBK
V9Fz8wfFemZqsLDG64uSFTy1MDDW6q5PMCOR4c4HniBLsfBioYBtQ5xfJ0AIQ/Y9TKSBv2sG2Daq
yANW/ro9U4twBg+KCKHZ4iSlUZA4S8ZLQVN+KG7uZzhXPB0w0jwetxDziarW9kgPaUSBf2U5j73d
FhhxZu2rD2Yu1/RxxXYM9kQmWJyVU8XNHdLlshWY9McMHFalQQtdlBAgHlrH/ck0YeFv0ZxEyR34
gezeWnfkIW2kTAKsYNsrDH7ZjL0dPcKioguD+7quWKGUZ0l5ZYR0VJkM/jp8f+817t398F68NLfm
ka4eRJk00oR6Hz/iTU4VCcUeltd0YXIMMcWFbHt4ZFGwKkYdKSqHmtEBny2a3ZkLkwoEMOI0Z9hI
zaostPsJokkAaCOkO3YP/bbh/4VagFhyyNnKme0YwofYtHxfpT8bFZFJAUbvmXBE8zpnP118s6XR
GbLIRbew48RftPPli638A6EJnFFjA4y+acCWSkN/r/tD+dqbgnxVKSC6exF9kzjXWqKiYd8f5kBQ
OwCvFJhsjw9iyYlRg/1/fhtAFL+a9ues/AnblEufGZSjZJJcgtQlVBUSgTyQigOwXpAVMwKEVUCZ
DqY5HUbmExAxNg0cwbP+rRIrMn+QVQK3HmqpZNxDuJeIuB/8ngW7eJJrh9VFEjn7bzekS85Gh5nC
Z5tO6tQleOWCFTXFvSd1eZWliMWOdKiFLNzuAJLlkfqpvK7kOwMVVuzJJJkGKzJ6x5CG96A0H4Y3
M3ZFmkcIjmVja4k/7gzFtWAnq1Z2vGgoWVHK29ym6YzTstm153U2omnRGzfGeFwCQuL1TLd6Gp/z
HNf8LyvEtHgrizvni8SQjQnErLjBLM6a6g43vepfEJAyfobG/V0Ivx3RPqKxGaX6vhSsDo9pJLzv
oFnzrF0rHPJvim71aXZYFJQohi5d5/pASSMNqbUdEhfbh4E/bZ28P3WgDsgkBiTNUDc3QY9r7bGu
cLhRda25ydlzpr32cUfDIJv95GYdFtTMjSktuPIffVa1UupuKUWePRqYzPKFFWs+kQKEGXZ+ksXv
BzzFM0HxfTzFxp48D0+YrEOSpgZPQ+c+YC6Yb2jZ01yAi1SW4KTWxAbxL7xd27ShwaWukDf6/JKZ
1U2cLUn4WNgoppJrSeKgweAK3Wxyx1D8gg/WRIFfWgniOfkXROkIpzuGbFMMgX3SfvlfXhybHwWv
M067PtRgCSUqhwryF6ffhzzw0Kp3m/JFD1cxohh3Ut+qIofBHDnka+bNzpxV2XZzVg9AYQwxTRYY
Gj8BNFpV0wdjhLxWJIQmti67M5Ox0OblchAnWkEhNlpNByImFOtreHXX4RAaEYy5wGQYJJNTXgbj
MuMyfgv7O/KhufQIBo2hdf8I4ke+kMG+0wsH/QG/rTSmd+Ivfh6ABlYwWqBhn+J8ditbiYA7tlLP
BScJGT92yXcifPTbGjzKT2AyAHAKcvpL8h0lIQI++JmWzZpNPSVGea+H0X2M0jBY6a2WMRYrM4lz
2K3qy06kiRSqEfDZAYKR0RRvskp/OGNaIrh0shwoANqFwGlM4qp3NReE3NqcD0YuvqafRNUCKwi5
tZ5jeuru8O9sttKmh/oPhk42Un/PJ22ZVAsFTmt3RhndHhTOojQf1HYb6ar70RJHy2R+HN2pEsv/
zWsbQIVXKA1C/s33HPpGf4475MPFvzJcy3QqtnD20iLwHGC8q7uLBhD75/enIK1gg3QXsES5HLrU
qJVQ6TZHK1ntCVM507M7y49sGs6Sv0Zx596FsawLHHYYyaZQIDtb0Vltw2zNXjW+tHYo8hwHwO/F
EPef49jfFS2yfQ+R6qsWjVdgNMgeTpAm1Bh6zwueqkR7LlzmGGkaqHPODyQErQmPITKpU8HCfacX
45za6XQP5uZ1CNqEaQtilGWzx0my/oZ+HoAzaRALiBKf0l6BGRa+j9e0gNKZaR7XWo5ZB3pOmsiw
fCAPCKzK38ffQjopbYy9O2hMKrhGZmhdgRTmvZvExEF2YQljhu4bBmYWJCInGCtqVKPDHK4wRzlB
dBqb/ogWHVmjbpT0Dv7WGgAkPYnSCKze4VWVlNOu2ZWJzRRQiLmwUV6S2xnnHlpJH7531r71uDHD
OG13kn1/+7ry6u9sfQTnu5FaWhIb3BA0wUr6lgcMIg0DpCRXPVPYUVv3Mvp4eayY5ttWJfuBDhdV
rgt5fsFIc77giqRZ3KsP/CUYGzG3eY8DBF54EZznp/y6FvnID79tBNHlPwESZkr5rXCosm4ObnoY
UVUwNj+yF7jbcIqY7eYNdZrRjK1tKfAXyLXtl/ngQ0/itb/L8z1XImeu4u4drIwMl6K8uZbYa5bz
LAZD8jdQYTqI7oNAZ4x6MmDG119u8Jws1Bvwhi19+cc1E0h1Kdba1ZVRAnSI+nCNbWJDrMRmykyZ
cptNySNoWTHPQhJmpwCAbFpvG7i3DAGUgKY1dAsaRIimuf2OXOta7uNjst3LqNI41Wt1VY/QzB3d
h5fP/Gz8tcNnz8Wgk6CrfaJM1p5RzgjMv6M3Gbd5LxKwjgViXQ/9IKuHSEd3ciAlNPX61a64CB3k
dmkGrcUcGd1nYjWxljm23PdXZjyyU5mc3HE4pKMbO/EzKJZUh1BL65oeZUjloqfO96o0hSKD37Qh
vDn+i4ec+ysZTP0uTfo1o6K06e5o3os1WTsl4qGciPbgUKILFWsT898UrqGqozh/eo9XmxqLplbz
xXYT05n1YsPGfdbqb61PA+yL3g2D+mW0xjJmyA5Xt8iLFfudboiGfgrvrRD/zL1UAdojPiX8omE6
QchZNrTKCsyBv5IXDuRa85anMPYavC9q9LYZhlUtunbFB8IwAQIdKQGCekq+Eg+I8bw/0VGZt3k7
bA39+ncaI2xZtJqX8B1mdiJb/p6yZ+Ex8gluaSzl/GFHqdNpDaeHq0UKvam/awd3ithBB3Pv2Z95
eo92/RGqDfvMZgUsXsuGvzQuV/yzSM4cYLtMlBQjDdTFhnm91YHsGYy+mv0WSG9cg49FuIpJfz97
ABLO81cPQJ7hTauk49MUS3gGeAzYclpbOTN9yV11M+jxAJawEPhzcb3Iab9eNErwlUtM1JnnvQME
3ged4EX8sCE+BKESCs1nXT1Od873BHR3nm6C4p8Q1D1QQyDHZ9i64AhlwggqZSCp5Ye2Q8CU0b0h
Qx7U4TYujWnN5ck25hsyHdcgVzZEDYP2cXzm3UpBwtO1HwrA4AW2sCZBdrP5oLWxYl/5sWN3xCK9
+Jtn0R/qvX4Gtl1famO2/d33dyoBdq0msOvH+T3woyQbr75wo94SFLLlZ6wVy3wEBNzBsKlypsxS
6R0Z8UkVRozD0iczDsz2gN/ZGsmCDWvOe9W/4ACAN7fBcXvFnB/mr75plEQZR5EDdEmgGUltWfjI
4yx0ce6l6l94DSeV1U4akk8/gZVjC2BFxSIgs4z+lEgmfIWopzw5/T0cmW66vRW2LjlZiTOjVrTn
kP7ECWuMG2mTktfffA3ApJxL2XwFT0lG5gnmGlQH8scFZNux5UUpRZFiGzTcG0BnWxFMBagGy9on
yHr8OOWulZgnLDjZyKtlI/maJaq92aiddHb5aJcJPgZhqSc7oxP/tu5JSv42H+AwqKa7r1JnYlm6
mR+beUyNV/OwUe15r4IcoTH5WCfwbejF8jGNerODZGN6sr0H1+bDHtQFKK4A6169q7bIXa5Vmvxj
8FQl1AlcXr7kUISkId6+zlVHdjUDbx7J+MetRq+bju2qG7pMOj9CEOywo/pQU4rj3+PK8P/PtPph
NgCHbo/Ww6s7bQEFC44fuEpzxBb8bBOzzPrr9ZTMTde/L37UubRArsWHG2TL30TKCQ22920dNeFQ
Ks3BgWR8zMyuwr3bRGLwnGhzR8r/rSI9Dh5erornI37nN4FzVVZGGjK3UYs09aTtKww2XwWQ7oid
zcYsyURqa/6xT7i4VONIoafAcH5gEcbBtPfmAlokQgUVIraWlg5BVoEU5ahJxH2Ztg0+Lo+ENOdX
50d0YAhsE7hHmhS5k8bmL1Z+/8lfaa+joUqszH5ScMYF5zlDHUnG0Xup4QlNKt2mToSiYfkC84rL
re9MP0M2xUcPGMZNevPkKiQiKQrsTKslzPmxRH0/BMBqhl6AytWCnKHOw1WcPeMTZYdF/uFEcq1v
oe7AFG4ccEIWsjj7q2rDXm69tPZKVl6fag78FrAD0mdVPFndwuAzDPzDh70uakqxJoVVaHasNyVW
Jl0qYPgXiFhFG6Yt+LztCgCrpgF515qZSe6VaXuZPKJOQD1xnxhSckSYTxl/s6BrTpOBCl6HvMDD
qNdKuv848SxxlxBWc2Bf233tQA4RoVaXrnzm/NPGl8NzYhtZLe/jsNs4uPbtfWV4qS5/wX9mXweg
wc+ah8Gv880gOJcVsDzJWTPT+z/3Qb2vHrMwS8MkgowcshhwqDgiNSAgSK6C/WZ2mTKaRZoFCFLi
opvLq9l/yuQlotKx/6YT5M/kVGf8soWkHjGBKDPYRxT3B7EmMGE4VaC/wvEbvk0q6ZdiwlEuRHVo
UcO5Xq9/x0gRYn1PvCvqUamb8GHVFDP78s8J5tW8rjulskQzAckmbI1UmuHbRdkL92RlzCPsI1JF
EK+YMrGniu4nw97SH4i0/j3O3i527u9h+rpv/yg25YpEAhXHVGVzcaoDarTzKLSs9zs/Vl+eSX/Y
S1qjU+9gbKL4P9C5fULolOr6Qu3G3HJVDJ/SBUT7OAIpTA2bRJeH3UsTAZsMZ9eKHcCgsqSFimTZ
CW7gqmpwgKedHgdS/7P1pdzTi73CULcmPaZXpO90t5kKYWAQUbZSPrL0TSbOiZBFR93ycM0E5X/X
LYXiT5tRV4v96l233zOpy+v9zyXmMEY1yTfVg40mpb/k9i7Nm6lR/TbTY77TyaiLTcfKkhL1pOgX
pbmHOVNSm9ubADmqsPuBmV/CFTQECgBcTUQ/koI3GB2lIewLD57YOrq+PhCigfZhvUZyy3wzvkvy
gc04mhBggdk06DMbz/P4Lbt0QQkb4MbrodWI/UcecNCQ/Ncfstc4zut/ChK5iaFhAGswkWKx5xk6
5JMacpwIZboAbNbmrJP22DP9TRYGke2X9Z77VXzB+GLs6L81b3ZIm/wKK/4l0S3ven41QIEtcPlF
Q5VLLSeojv2C+/CSf9+M5hDg6s+PoZqW1QanzMFJFW87iOa+yEqWygRWFoVKVJyCpYEerzmBNiQ1
Bx60yeYT+pfWzFc5KTDyAw972+Rgbe3svCMQy94OzTMyDddUClmUeu5UEluVRlbk3I24rP3Kfe3q
DZJMnQhSobJnq4mh4f5JehdH2F13tLNjifDvy2RBd/rXseVfqXJWPycgCCZnd5+OEKY0ihQ0MB1F
wJ3DUxbxMBF8yRK1e25rnph44zpF3DDSoALwdQYBh50TTVUcgtP7dXahN6e6H1g0lSYvuK11nGV1
NtBbmc+GlUFfVdxupd4cmplq4cC9g1R7JBXbWqaTr5F064iYHlnvqcyMAy/R+b6aL+RpjyYQoQI7
E93DCxkhcejAKs7Bnaxx0Agt2ur9Jn9J/WSxK6F2Il0Dh9hIOMkUTLNcYOdYkymRSS/7Q6jmXsLu
8hzWS5n7rNsIYVjLzcpGeh/5rzzcATr1L2CgoV3H4vbR8OHjp9oGKbD2B4ui8ZaWWLugDyFCEyil
joA3Ho4xIz2mKxPT8g+GnEW1tifw2EbZRXhchAEDGl52apUrcB3UINaFNkyPbCHE0D98mwaBIXEc
UX/8MPuRyqRpO+rHei/1iDt2qL5rV0QT3u0m5X5T/BDMqAtw2xd9Vc0E9KcgREL1Lt7ZV4yBHXrp
R7pqKxinjsgRgNoIOC9VdnYMURrYr0zIfj8ZGd4g2e7ML9mVrnSNzPDtm6SxUcZQERsX4DIRiZNW
U0qXs663mAx5wNvId7ezCSTjv7e65qTomWc9YcUmBSPqbwvpZ3ZSrNxI10n6ipyZGpoFETDrOp4k
3cjyOxwcgOk0ktz8+V7Y+s5L5VOYaTxLKmjWz0Z9Ex8j/UBDiENkWN1X391NLkfi7UMC/lHKukVg
KHyKj84ILBwOBQX/KmoI5QE6aBbLvWEw0TL/5AAC+BsjkrMkvg7TsqtR5u/7AVYnxiJ/0OsVbx93
nOu68/FOC1lAwsFQ5k9MyvK2aZrtBK5lNiYsGqhb5XWLiRLzN52jchAHv638go7spLUMPjSkVION
+OTpMi5qyBcY1OKbgYhW3O410qhuIilZX2seT5nr2A+TqWA6fA335ghTIvx4JvtF5TklimoNKLU3
OrbioF/BBw2seTDWboOFuS4l4xTEkteAb43spn4EUyjBBERygQc2cVRt3YtzLNRd1JsZ/+xzLsen
XlAcwybnF0CsrqiaJJ5SE1R342OPwvaojKocLTw7TmT7uAMqkfq/sjxbnAPOynP31Y3yBTnXYmmw
2aN5l2K7fB+xZKQivRRnsYVWeb7C29RagLqZ1K/IV+CC/uVPSKYK5ILdDCXSVUh6PtFRmXcSBu/+
hqnDzEXBEvpFycSu1Ic+Jh8rV1X5OBuHnbIvS6lQQCaOn5ZMJYt+wCjQ44KJZta+50BKhTx7vjdR
gV7BNJN5afMY00Vqpxy/uSynFL0MnmR9BS4nO8V5fUa6/Mvmvr79RWoH76+8ONnjFKcyzCz9sMtP
1Wuvns1NT9ycQBRNhDXtYtDWmwNjruu6KIrlOnQM/9Z2npe+4vXhy1HBQpuZqTsoT8WoLfcSG0vd
LfCZHer9dkScA+to2CtPTCOzdtVbLhLU8md/KFaO1iPyXcVcFN4XN683XRqJWn7XuBjxb6Eb3qkR
eAvPJrettouOg6nPNLJiPdZIEOSy9nXo9XPF2ZPdpsOISI6WFjCoFtA4vWPuVcU8wCH9QDKGTnW0
ONNJ1pxepkPkq01dv3OeXttB8mVuVeT3FXHhpYmmUTxn09PCRXNAX+3CqigRHooFogOZ4BGXGvyl
YhJwM1WXTmf9a5y2q7ah6ysO2v3CGFwGQgSZrewSvTsY9IoRzYXZJia2UzLRMVe+4Fku7rgso6SL
IKQOxBDstlOYo4fXB1QclYbmYxEwHWHCVBElUkDnmmV4q5ylPYUTaAEVxb5yGwsBVzpkoE3D+TPa
Xk3QRoxYrVN0wQ3E36iH4rBY+5NTeeYmd5sDtvyPcs2UWK7RZRzValyhBv6vaECHZN70u/B3vN2M
aTV+8cDVsnh0+PFsOZDfrgXguByWwsIWYq7oeMdvoEGV6tnmPEBtwoBq23ZmuaXFCwZE0rdY0M3H
hPOtWm/VwqVJDaBdnPhXS8NuqBZp2gw4ATgto8Xi6250+EPLmzXQ51eG2n2H+YkI2T1a1Pp0YZvR
h0Q7DZRSoR99/j2yrmmFc9VepZU51vnnDi4uBuzW8iAGQNOUVQoCA1R6C7Gp9Uo9d4PEldRRnNyd
RkX3Kpy+R67teW4BRj+ELraJjKzPwFgb0KNNT7B0SfLYWaUVCAc1oNoMDhkk9CDe3c5m6PRBXTy0
GgAyJoZh5/2A48lpDH9sdC2SzhdzuNjDDPFJOSUwbWHw0hhmIWn4tGF3juSufG4cQQQaURKWMBqD
NSK6exvQSs0kvYDcufMHFr0+XriGALgXkF6yDW1IRjtvjnY/U/Xj6aJg19Jq8/tNyQwD5Eg/yl/6
p8EIOxfgmEOo949jqkinN+p4DG4Q3d5P51TmcvxmO6huBLjGWWg3ldJ4yuZgeTetl26eFPS3ICJZ
rSw6vZbnmHc62aLM0qCnry896j8dJajtk62GV4+ARvI2HyNNGmkl+pJPnu9/VsNIe9hK3QcZL81E
A44Sm6GMWLrP/mzKRbQxR1vBOnnlRTa5BK9EZNks284XqkFqS4SE4kqMUwYIfQUQgP8eOGAyXLbe
3nDfISLRLS3NH7HWV5lBQNv/8ATz3JpDgTGWCFNlQvWCn9zYeXdxNyBqmC0lXvXVR6a0HOAT/BAT
4DJGysIh3iumBKwpSGJbJ3Im2mBenRDQO1kAkHOtEfmzKtOSBSq74+J1POkVLe7/rrbDdu3QhNYt
b/fm1lkKig5vq4/kyJOy4oJq0B1tjuYpBsUmgpRnN9g7dlRV6pItCc7bl5N2kBfy+7JOzuUpsMhv
i846xTIYdGcyg0fKVf7gMyLC3GFmrVb5M1cH3SOW+R5gzqUWo0nTLnwAiDPjxEzc8CV0fgm4/stX
wuodEPkK6Q45v82wj3VH+Fwngkdw/pfW0SBsz9DAYKNoW/VTCa9nr3IKJuedQxf9KMwaXrehtJLU
C3RIiJBO2t37Uz/ivxAN4aIz4zUG8y59GCefJCUcia43yblQC6n59F+Kyq96RCMa/GTpRO+jKoWz
fgzHdPB0ndFaRe2RhD0w+aeDFyFz1V9DjcxSktYxDkisYj4INqs1+j5W4fJA1KYXjWbm/OVoTdFW
PLLGbekUa0BaMlg75+Mz1p0wvVH78+qFsaghgC1ciMjc2LAcLZi3ZcEwAC3icBio39FvvUSI12H2
GzhuIRonH2DStMorGolJEm27s8vcz+EtAXskKe/W667u26oapoPd93hQO87VFgsPSVNTG4kZ13NO
69v94px9b8Gw6BwdWoYPiqXN5HbsNy9NJW8F7/8NanPAaenXLFyR/PAjsQf7MF1p9ztmX6huIobG
ueRlZX8Iuj/KJEzFDPeGXmhXXURM6sJ6MzRRAtw9Ps1zH00B+YCgYi6BxVkhsaZy0Ijpf3HTMI1o
IrAkmC/inV+R9zrLGfQDECK3Hb6cW8MVYQ/ZIe0ZAQ8HTp0qlHqVmZnmR9xpqHV7nwpG97Ulrrix
esfnax0usdo7F0uTLtLPgj7BqH+Yrp+qZgWFWZRIWc3FlE+R46JMJzodkwXvK/xzUBp/xv1ryfVn
E52s16y0DTD9jFAY4sQOCgzHZb+RPDHYEtu056V2MQpmI1cK71Nx+K7rochr1QwDA5ypJdAfpFeY
tB1PbttdGIzDIk3M609c2B/VPT5f0amrai00s6y2nrHWdHLP4dwuow6toPpy4x9IZPPLha4NP8O2
EyPlxXMfveQ3WP8Mqw7+7mMckWI+dk+gYBa/Bi/hAS4gFMM7CHZv260M+Br0loROGldyK+uET6dV
iLpSMRCxnnB2BK4eXwiuL4slda7fXkVyAPuKUaQW47pwkgr+B7ZMmbq447FqcfvLju049oO9F0S/
t9Rd5077ee4yqhEHDeeTYv04bKfQ/L/buF81Kd1PKBFEnnPFbSmnFd9prWDcfK6Vemvm8Py0wnHT
IS5FS4EYdC7fzYFsWerkrMVaVJjPXOw/oQahKd+jQZ0mL0p/DSHGPkmnMr5luD2/PcrWJVuwN4xV
0U0q7Zb6Yo9gkPG1qvZVw+/YMRnAyN87DEJuIiULluEPnkHScLRvfNcMdwds01S0V6Ngxm3FYKq5
v0kgXi9gxe54yrHqZkoBmxmaC8USO6yybJnI0JJnmLOjOTdVdIi3NKbHgpdEtjGlDaG7H/G2EH2e
XSoemNFzl0LaQuswpRofx+SL8A3f5mCJYdPSqFWLcoYbUP3Mgt+c4dcMSoI/bkE8mM/WBNlMtqFb
YJmXwLlkJi7CgMfKwVyCrjDtowNmo/i9vu2puCzKeGdeclG4D+Nx6Qv0vCPL7WvmFKwjARorkf4o
Lmf7twyINrzRbrYmxQ/hHYy6pgca6SUUA6FqWl2Y/VT5ZAx/gfaQIazKNYwICm9rX7L0kueiKiRJ
s4JvN1yUVnIhkDJx4Cfz/1q5eBMumuk7DISPKemaFe4jlbOnmO1cR1d6fnDR7RF4joutxNJRE+Xi
H4x4c+79kBDZxt75DxS6O/KOL9L5nc3OqL9bAP98KbieDaJeg6yS9icFDTUSvYVcOVf7Jb4oQUDC
l+cljJlD/K199oouAJZorXD5VZypwVTjd7LLfcBoBsTvlzvsb1fCN5xEQl1CRO8sRtrXfbUj4QEg
oP9A4kC3FEKabYP207/9E2JTSw0BMBplHMk0GxnbS1u3G2V2MJ4rANp6xS3JsK0v7CdLs4HKB4ky
6Wc81g3pXAL/KwG8zfyN418fXltzjNohV7UvFHXcvDHiAeSUbmi+RqD63atqkOEEb8/knIxfsk2F
D77IA/pF2TGjtZ0f0wRo8HDPEM5dUpDzcKMHQsClQhMY3V6jeiEdIjySRGZI0nV/20QlgrxDcH+O
/vgyxqYIbYwtsrzedQ8j+MoD2z+vyOfrfVxy2qIKHTUe88Qas86KCIvTpauMV+HY4kwvWDOjU0QH
OwAZdYSWLkIffKUBnrd/Eitp8YZn/7da9sraXN5+5XCUgFJiCfipZWlIOrQPzUn852x3yIJCNai7
w+rJmJntannWr6cooBTK+hsMXH9bo7+Mk0INegTfYevj++CH0odAsqrXDu5x1r1zmOMW6xEYW93L
6jhV6x6HSY+/KPfAieBmbPWfjCazoOp9hUm/wE7Zt30NyKEyJsqbkTagPt6egCQYEptk2SWb8xE3
SGVPkuYIVjQ3SQP14kLXOkMbXnARfVxX26cDwj4NJKU8z20V9Y/W3ATYqHCBfWssnko+dW0ydYEX
1D0HgJAv9o9yXl2fLi4OKrY8rooswwofprazrvL+uhM0hPPW/TPtuYy8HxckSs5rey+MdXRi2Upg
YlmAN4yx5XVY9dIUH7GgC8lf+j4jM5GlBWxE3GnyQbrVDAIxfsl4yxf6cViFyzp4PHEhC2qvlEtm
zKeC7QedvXP9rD+qGX4EkwLMvU4jeJeQRGEX1SefQnHEAksnco1LHY53VgIPTjLvCDPG1EDdpQfh
uSo24RBc+9H8+E1NyhzKu13amvJmO+cMZ4jLxo2YZVqAuX2ssduEOsMzcJc9GKHsKF72kn9wVI0G
gS3WyoIeR/esWMtLbIAvy0syD2IrLiSzw+VC7EPvDoZI+9Kp6nNVlhKO/aOJb+au7MWh1js3IPH4
zCiWaKAy4OnR+wfPRZuJhRXv5OVyhNbaltOSFt3OcaaEypc2MDVKLn9225dthffbAHFTzP6lgke9
mmOLBuR0aHZMmyzhLsjMQNk3HshXaAbr4wi2+g3Z/GRo48QppSzLHfvdD2nL+GXOcQ0dCKPFG1Gj
FQQ1jrbVkGogL6sv5JS9Lvz/icaVGrkM7JxyEdWam8MXd35nDADLABabsIi3S8JatKx/tRF1wDhd
twO1GCmqufmeRZ0Gx/NkaVZmoe5Bazd316EOpAGH7p3idCFfSp6LQLMmjumIhzaonMijshJE0ZE1
gN4Z9fjGLho4yeNgD55OaKYTiToeWvBMv7TtY9cS3N9H3w6F9S4mdI6ZmEtgBplIscW3Upq3Kehe
Yl2KlABdxBs7blgweoAx5tK/0y60HiH7Qo5E7gwq2nEQKeyHmAc047SJvVZDx/YfEmYR9l1jEQGZ
RYKboA51WyVrSfSkdmPVZMkxJBM99ihb97s4gSfXjIcf4lebJy4ei51K+I8dAOguG8HEISY/XxGu
Rwlh6PJUdjAJFs6VfXkls73GNC/acnsjbWvK7RA8qo6dslOJNNkbJfyGvWxNGiZQlD10rZB8wJp6
/SL1CZy9soisN6oX7vN5zgKDj5T6DBlGaEeq01jJhA31KtWMpl8R+fP6Gqbn8iB3KhrP6l78LWA9
87g4sF/4tmqT5Vhmkm2iCPyjxqDIPsHdrmVkPOQfwNHf+czLQt0PSYrxcbYombYS4ZmUSEw/a0Rk
3i/AWKyjZkvloGCQSCetP7n9JGjGVMmMFAB0dzKlQXui6ALrbnxLS57UnFyCzMcL/ZNGHrROldFi
DaY3t4KnLdms45nNzsF2dAABDUqrkP2NC0Sfywtbj38KdsWFFNQqM6LOifgUx5gcaxtiWl+vfSPW
00H6KiBsMP7s3d0LXudQAlS3Hkv6h3+gXok6+7FWD688ZeXAYB7jKdlfMH7CSbrNiUnlw+wryRwh
Wnqrzt/kp2TMNPNtfXhoAOLNeAFtpaeBiqLujKKiOQRmvuV+UNEDR5q9TSOU8tXydzQPTH8Ytrf9
YLvlubfgV5v9L1nDHVNHuUEpbjxTzNj0dSCnevyeq5DFM9upGOItA6wwfViHtFBGfaEFJnwthJeg
Nqwy1YNZiOFqh04bjX9MynP+PKfux8Gxg2YqgTh0ZD+lawMD29vXEh7bimxOb8mByEPLfq7YD5QC
bK4OStuMwKhxez2F3m4/e33KZ0W2/nRagVZjU6yX9wM0REtkm4oJdSYi9Ieueq68qB7NdpBXamkb
58aCfKiSYiwEDAgYdB/cyZlzolWGSAmH1cf2mfhcl531zcSnPnzWe0xC1iefN9quwaCecDc4MUiH
GQQXmhMTR2/GevmV4ma9VaxaZIX7wmOV6O7CapnpeRHcA/vws6XkOnKGCMMYcs1lDKR0YrgQ14Ad
esAXXhf5/9GhXUT+XBiFWS1KdW1jTP8AM9fs1D2QUpg+nHY71LvC4CQhtQVSfG43NM94JnygNzR+
o2cwEPaTpLySrmFzR+LJKyCNo1QPQodHqHpaSPKVD6LO2yviPg0vnS+7xkaLfRPQDn/7szMWlr/i
SizUrdznPqhrIH8t7aiH2/BSdW9JjGCLz1SDGbjbyXmWzzYU8Np4yZm96GF8KFgxSmqqvJCGYlgl
LIc/zqcSxsaH1cwu0Z+UjFr1dq2696QIP3w7zlWt+evl/maodW6esqT4mhvy2aJiYYXxYsVSaQHL
w0aU2FFYs0DHtpU1odSv/G1noLHtPc2PVs8zJCoFmKcxl9g7bt/usaMRMofo6eKUPMUvEgZQMrt6
S3PP8VJ9vBVHIoYE0G7W3zPTUcTowUBt9f04qG95yUEcBsBuwG6tSfLFNZJ4UF8poe53VCiSTCvw
vODmrY/kcRZiW7Pp1ToDSK35OYsq9bXio1RPz/P9zyp0bU0IGWkHmTyakL56fRrDRP5wAHpLZ/GF
Mg444IqqdX3qoTvB4KZ45AWEQB1tZvuMp/dSMvK1TRQljQso0aYaF96y8RzgNuqnEG0ugeWuxj98
mlM/6oZ/xjSmYeqxPMd0ivhNUtYI1uPeP7tVIYhjPQdv5FZy7QlrpCfoC3F8lE4HwDdbPxZ61mPw
LZo7PwIOU4eGeWnx8xmMwIwiUx7nKWEwxp/hmfo2F0sMcVstCOHqfPJrFBBGGCQhWcNGI5jHubtT
64jBL5jDFxpl+BEGzUMfv3xMtYNbDJUPWd42tsGl4mznQ95luSEa8DXR8G6SGGV+Ye1ECK9QVbeO
Rn6M48jKQrD/Ly862OwmuZisPFZ2mKni4cqrALnrAYh6wo6fn1sPrBh6pZgU4Zbt4+NJPNt33UcX
JrKoBqSnBCxsKilfXgAMAZEoEbDqcxz7gW5QdrWpPHlNUkalBFhdoxshO8Cg5tm2J9C3j8K0oXco
DF29uQwGXEIyVD6gZeh16cPD8R9zYSH23wJJ1AMv07wtcZRpO7oBPbkKFcSlaNJXQrkjQH7Sv6w/
XaPwnq8MBjkMFTrtG85IE/biGizS9X6JamO18Kjes+hsztlhQ5baEUlfboF1+VwM8LuAHahjIl4h
GOWUzLIdrf9MVXt1+PidHOv5APnUVJu9urTEZndhj31MEKiMvu4C3j+FNyIRRa5uzImP99Uymung
ayNq17ToskSroqXCH1T0e9exEgyt9rRwG2v278WjVT8cPRrGKh6h+houFfHu/uvZe7nZk8d0JLDG
+I6Up+ENV26NWEKxdsFyponP2CS6DPwCStzoeIYISrXJziEmwFQXj4DNlwYUHiiH91ojS7b6p0Ko
F7wDEtRnuk6A5wP5VVhcUcMh94IvbBiqcg19+2IARrKxXhvf/r9HNuoisFLjyRvbmhXXeaSYg2Sw
nGyJqVuzwwu4ail5ugfStAj3C1mCbYX+fX0E4+NEbe9Ivo8OgMm7pa/ZJryLjBlHQz6k869vNm7s
+gLmUQZPn4iO1jkdu4sEJ4H42tsrYh9yoKdvd8+SimUdnlVvLUt2CmO1QDkwl/JkYKYFavZPjI9V
TTvRfvXMP5qma9d9jmqi2eviy7oBxakfskvfVvq/y0j4XtQg75vQbNY4x1ibndq6DKwJofY6NQ7r
1A5jO8z5h8hPJ3lKK1pKXIv0s7iTjfOgvqInA19P0HcQFQ5ypmANnamYPd+9SuC/X6ybc0s7h+ND
4No8skBjU1Hq4Bvf2SQcy8R230ToI8ptaf4Ot9IZtKSs0gW6p/9JTlzyBjr4ynz3BjMh90cgldTd
yNLzI0fwcE5qVV/wJgx0DIh1Zh96ZQCaXa4dVrQLxipL1Zd4lmoReCIIQojOxImD2ccXjEWBt0UU
KvZt8s7DRxyPCDeovXNDI9ErH/q/GManIWK5DwDUiYxgJx6oAn3lIsG3dnhwKlASP+WptbasJEJl
CqvKCgBn2aQJ/rynjM/WHzSupdNKlFA8HVNoCOaAUQJfkPdHCoy9TUTc2RqxEy5JN4JZvmkh8mdK
UGlXDgjzHGsQ91k2rjxN52bQHoObyUlHg4O3M8VcH7NgiGUiqrNbASBvcxOJtNijmqOdVHowV3zt
vo4ymaPnJKIHbJ4NFEtkGn94cxuONI2XAit+YatuyJRV4vrpcDAN7Nx3Ld7X9m5msYyxcW3xw0xX
d10qHKWUTQ99edUnqtDUljctH5PTm2IrdMPTEnXDgZOcXa3XONXJG9oe0yXcVAJLwML9Hxr7HJk+
xyRZ31wuHIHjPj2Khd4xb3xyoxlO0KZMO/BDZFTKiBaEb92vODgT+1klbOCFPnCS2HAUdE0+8hG+
ldDb8tnvBW4J4G4eCmrdvswwxAzhaFeiPmr+2302CehajjFcveLf8+Nf2tTawWDCxP9qP4Uqmb9B
UK7IHCGzjO94NseU5NQVFqLGZaEP24BGSWcOOKbjIiZktBj06jZHBpeGAMiPneqozCv/FMED8NRV
986HZQjsDgCGlvuGGHPB8WrvMlHiPEyoGK/8q9GhXhyCXEGde+89ih3exWK19nwKs6bYc40yq5qC
RPekPuR7NLk6QRpVl8a2mUjiraKTE193Bkv+HKiB7QpvbrRCzfAtvGQ8qBx4mGw9xZT4NDhx83ap
HW5YBwX4iNLCmdTQtO50l2RHbwDM4V3gZxrunxpV+r2FUJEdNmRBFuVPXR0YfETExKXrH5+JlLfJ
nvIbMu8Trf7hi++E+hEKdWWM3ivQmgMYBm9fyMPai7dNuqqKb46wNL8txyvH3BBSjNISJdlsOW+m
bL8gFPVIR7OBxRjmZmwYvjrvjKCU4+35pl+V/ZHuVjz+odh//7IokcgyS7Ittl8Is1bVecBWkCei
7sIHK1B5fA2q4b979nMUALxj1mUixHnkZ4xJouZPGuki9Rt+ERt8Ea7MYTd39YvgVwSimnd7JmDG
P3lc9xh6ZgGjnNg+Rr/1qIBwmmiOQEaWuSW8xJoogtIsGIaaS89etlrE/FmsafbDJBuSDJDVnII7
7ayXq/ad6xqD/mowDfoL4q9HLiEGTj56+dFbWazTaobVDIO6eFk8iGrLuymzuCKpakYIY8q/j3uG
PGwHEtjoH22yg76moRCUXL37BvpP9CSo7ZEPS+lmqIYJ5XUpnrDawg7IZMMkY/xowFwO0eknj+3K
37W9Zv5RlN9QDcozI2WdUHl2Eul4rpkLFIEZxisU062jNZjv6qSQhgDG+uLCEr3QzH9w45m0OLuW
f8HGLYcZAx8LmXlMN9sg2veX94aKd7Mq8/wdfBZpbotkT2JTfJcKW2DtH27ugyKuoKUvPEd8HCt5
KcLrcYOHhIj5HQwesZg0pvXnvPRWjJhZt1Nk8vq9uOplc4iBq+I526uEfLnvCb77tYwVN3eYo+h2
E2TCaxc/duGyGHOM9g3QAY1wR3XjV2EH65iD1dOy37jUSqhZy7TTq5pgcdBgarqpNXtFGeFAjBWy
KW61ITQWVmYLQ9+MLV8EEReWeP/kv2Kke6BNtLLFeomiDyEhTX5br3vx6mtAC5LC3K9SXEG0Jb1c
zl+UcF9egqcFjs04LzWf0ICHwCWIwpTVEt3ks3JJ45STjs6khI7ENrYLgzc8gACi5kCtBcYiPzon
TRw4mNNWDgOnfwsV7t2xtcJQDCzNM3g7W8z6joqjnCBOYWDYU4X6QqBMKZ6pf1xn8ta7T5CTmbiv
871xp/VoHb9OXNhyxd1VE3b2oxRxb1ou9itld5YFis/lyKYQrqY9gzAtpyxC+iKy2sI6AM6wN/V5
zkH2PUH7PhynOZ7mmsWzt9qpjWFq2BfAUfPLr/e/f6MT9XQpTzcmAXeYskJwrjuIphnz3W2BzsY5
cGouakcRQvNxsw1E2goSWb0a/6mNvggreoHu+OVR5fl6NVtg2KH4UET/Bxi1P/M/5oJv7BSQSuzC
4buCzd2HZ2heUdJlfuYJmQMdskrFEwCTZhf4wi/Qc7OOjqOgyr31r9wMrFyrIIsyJq9cfc0EnLkq
ekXY4QwOYLrAKXdeq4+xg9HMS8ez0dLiWh+sIbzlKj0p+LF3k2dHeEMGd6QCF4yWkkN+KGfasCDN
h+DUQuaEKm0zNeXAAMu65aZlCll70crztSOKgqbrHGLDam7RUzf+3BxWeElOSlI5BBgf/k0i1alR
ayEowMuvUg4oryZ2az9nexHkplgj7jzZ+HsmvJf04juO+Es5K170zQNEoZzR4Fnxa39gXAqY+O/J
OM5TkXIuZgDmCVaplUFdbmkMapnA7umzpaGQ0x2Jf+vFcuYdfhz7SNDV0Zr8adxw21/kGWHMcr2W
rhb6x8X00frlgFxVowfe56LKUqsuk/x8NbeCNqHA0Hx82sJ+aR9WrvrkvDmGRd/c3wzwEqAdpXjj
72WadzlzWPQUO79PlRjktLN194ujA3/vMJjANunp4cdckWoOYRbi0cmhBDNMA4HGXwdt5XYqUMuH
Al72Xed7CIyc7IbTC7J1OyG8gVIzkYuhev+1BBZbwUrTH9yjn7b0xKoZs/lkebQUzFuubjvrNesy
6G/ckBXls775HB/KWagC3dfg6zA3opKXaWEwU4QmnlcO67UAxwaixNv3A6YKe2QCkcjatEyNu4eH
i2IpqhnrUAf+r0qAUtqQPuVJQQtHGIhf4Kx9y7XU1xpBo/msr8cgAAMWZYSnvli3Uo1CD6yHbE4l
nxpgKg2N7HKw4UuKmFuXrtwl/gsAFLeX3AYCvTFfIZ2SvqKQIqYxAQQim+DJHpNbiWvlcgMT0M34
lqkyKyiAEVUs/a3sqXiLj2mzPKhgw/3a+06cwMJPEAj+orrPMszj5b9NhgAsyWwWvknABdmEPZZ4
7A+u+of5ckhI+Yurf+UWt2QdYB11O5qlsWXruBshmELVMkLYe/JHSZ9BUzShgjRwcTJ98oS6AxTZ
7ba4vZ/nla52yAvGcVEhy5UcO0JboWi+Nqzhf8IYN76nC1wJyVrTebPCJHSYBvLzp/jKGuCdyP8g
cKZxbN39iez8he9Mm4mn4tEsjjpblucCfsshyRu+ucQ8xA540nXQZQiu7byGCFRqduUvscZcMmLx
9JbmKrNQwKJZ8Yp8GU5+e372qOAYBYeoEoRAwGL4DGf1Yyo8DMTPa1wQTgVw/wRtAR2HHC7nBUPx
R3MHFX8zUmifNqAmrNs9A36iy5dg6wqrjKgfezgIitEznMYyAYxnh0YEqReiNuAdUN6nl+KLjv3o
PisUapZCgFdpxcKxADun3gjJyhJ5xVIS3/ld4jTdtX9cxhNlcjCX5ENRxzbsgvAGcLcsPOBx7od8
mP+a4mstzYGBC4srzob3NTKRSNQlpc2E5e2z/aPEh7HpaDLFRpPQTy2FQn8kf9wGXFqIeyw/llPc
XPO2LOxNzJKMS5uUPvAXUVx4tnP16EHFVrpkmuqYgA9V7MM5I91XBLoebZ5jf7T8zlgtqlvgvjuO
tOyCtqUlkI45QuoKKpBZWDXzeuzhVULiIaTelHxKODO2vApuw95zqa1mQPibHgWKALx9CkXAHMCY
Lj6wc4YErI6mBmBE9QY1QNiytgcloHJVsKpG/u6KnDUOwkfv3IMv/LocpDl2tA2PXCEkfpdNucrs
W6E+G9bxBERnBrM5ooZUyWb5gnLw258cm8dJSEakCoBpIwyO+A7DRRotB1e5PuXDXtay3vse2G1Q
Wi44zVka3PYAcEghVV9btpdXBLxqUNzgEfMUExY468zWKwlJmO3p+px7SFJHTkje97dld6ULukcQ
4qSX4iCJKlSoYbSvpqffdCU3SlhznHcM1FSUA/jWFhT+jLxeeZ8yP4/LZAsuAdEvdEMGm+0GOM2I
W8Au2m8P4jyoqQ2I6B4AdX4NXPKQm7SlBtVv1tkZzWvjJ5L/eG1hvI1tklXOY82gkz52jHFFEF9f
mRN6g5MSokP26phnXNEhCcve4Xq4iS33+C2sMoMCVPWPKK+IYgz9v2vwp/neNZi7BEhrQls4Cmmz
8pwnj7iN4sC0CYDP8HXEWRmHx5k/ic4cJz8nMn4HrcUTPagUVQUpL0jNHLbSZkqVFaayxjjbbiFB
pBGheq7CdyBQLHQ6KrMq8MdFkBSftKJepy8hpUoBaZmhfEGt44bddqFBAU2viyXMoOgwL4kxgHTu
aTMkd/c63VzDL42rfvK4K0b7qk94cUe4phoVSc0umU1Sjp9Zx0sl8eeoUF2gmH1eEcmWLBrO6Jn+
Hc/vZQaSttj5JDZOPVyswmzzM/7eiA5q2ZjKtbzd5AcOpfmkWME+ORrJCYHnfVVa3nxjCZydy2eH
zxllaspAnrdaTQlMI1zCa/bCjYhIBXThjSlm3luDX1zagy4pKBtYiNTVl3w4d0Enxht8HeCez/55
XdslvPs+WAIf3PqG3r+P47gET+oT/wL/Q/Thle1iwIHvP7DeGb+Vcz89WLAFqc4JoGIGJDk2b30f
3XgFEPygxiBZ6cPEiUp97Jnfu0ioIv9lijc7IiQQsPQcVcFJGNRKcJf4nlW9M7sqDNlwqD8um7AT
+4BtSBVb/WypyvuJ/Wv2DPh2q7gvuGMsjykbVTPZXqLwS03THB+1VBCrOYT3uJFX1uytD2vmmaac
o97RP7CEOGA58EcZoxl4GgNlFenfkMd+4uv0JsgHq+CuwkOjLGqrrQ1FLuytiYTp3fKBGo+vk9ru
gfr3fLMXevVJU1hbgqq1RtePAaBns4D1HmSHgZXg2RfhqUXhUTcSkNCDCTptFzm1x9I/GHXylyiC
VCyrZn1bp+nFD1hdRKu+jwibASuJXibFqPB7rmbz80MlZq2n/AM/Lh/bdaQXOStG8t4ZXizKfKie
bSqLcBG+6no+fdL2jXA8vAyGylNOl4q0IzVW4FExpg6OODPThz8lO3YIk6IKvmViZpu+IFM+WtAd
jwf2mItoHQ3b1opawobQoADWZyWU3m5ILQfNlyl2M3MRa7yV7jZHjRQnInoWLMNEx3Xnys7qDnJx
MhjsI2wT7+3q7yMCkLj6inIjo+ywqtJvDtvF4CXIkfbhqVu9DwoxKyXQSdKVFQVCUSOWO18T/R37
qiifgHGx/gSgyB6jnJhm74F5rpjFkqfMg944ibflA7j1zafxfFhE6gztbJi4uLPITeh5no5o6pC6
33h0Seu3g4WzRO9Cn+miJN9/j7glUtCE3BV0oCDdw/55GG5Fd6EqzNlqSffmsK6ceGsxMj3PA3yq
4vRNh8sHLks3mdc5aIgPqyagQPsaW6Jy9Uyd7+tjWKu9W3I4x79GkA14yPffGgiA35qavLW1Xm3y
cLGoKi7iegqR6xxFElHNzUKYgaIs8H7mX3c4RUT+jLi3QN2Ys6eWhlQGLHdbYOILd2P8Vy3GuIi0
xlQBx0W+fEzj+ebdOFSTut+wIt5z+/LiOtNmmK1Ms9TiCrDRCtTS/8mAhMOL0ZJKgcGXOouh3fpm
2wQ8UkK91uOLU6apY4PJDL/3LrfGXyg4t0kNPWr2ED6MCwYxvo4gr7HuIiY6M9R9BtaJ7wxVqpT8
xAc0cx3Eh9gI/1/yfRys1DNm435L104Wr9NC1B6UJW2FeXhHrKEES7DkcsWHp7/Nj5XkubTIJfpE
s4xU13Ykt/inmpmHQG34Xj6Uxlk32CzBY2BAVyWBlzKAxn1m0x5EP5V3Ttr6gXS5w6vDsskwaqt5
MZe4ngoNEMHJ5kA72N+uz21x/j1wYWjDXDhIcZ/thXDmhDJZwXGOZvxE0WwKFuSODs69oOWqK0UN
nxc2iS/OfNP+X+AWJRVSMswp5bLQDMQl4CFW+Hktpu/MF3G/qipq8sNU2c4vhoRbBMW5rYJe2ajY
R9zKOJVe+1FP/iyFxbeQW6+tWBEuHLLFH4scJJSrsVEX941Sz8S6wFpkt5zfuJUgXld3KYiKEcpR
GqkfSKjvuxaYwiWK4WRfPC/WqL/KTH5v2eqW+XxTiR4TPcE3EhOu9KaX/5HMq0eZ7WOLthlIzZyA
Dkt/GERBe2HqmnbC2B8of85nmDgAbVwZM/8akRnNqt2esbN343uY1oDEqybwU5HGtzkbMQdr3sxp
r+8Td96ita2ltgbrxvtlvRHmNvTogUnWtdtYEFbwT+asAUUhvwzEx8CYBIubPXDulgyBNEEofI3N
IjR3H1iSodBqTNLScBGymWedcjqiu1Qd8n/LGG4qta8dPh6eQSAEKA/Mh18seaxvZ5ZRu6gZ9cA5
A3aP9oqukRsGyRNvxpotlOeSPvHd7rUNvYr0g8ZaDj5w0ISJDVxUF5DX+gefRLfnX1IIBVPSCs7J
TUwPdiR/Kql4F3QvoLfpQTAROla7NlTee4/shB6lAYyKgwrqY4i0JlONKl3qVG2sDMWLOnKXoQei
iOo4YvCErlrWPnfdni8gIAc3LsB11i/rnall8s2k79fC+AIaiBdTlfGeLv8zJAynG4wA+h02sX0S
e0zKq2plbDqPwSE2L/bClqYlWcjPMsHbKvK0dueSNcACL+ZG10zdspf1/wNaeVmaZNZQN1ifUBHm
U0Bq8QqOgNjhh1K1On2wzuQGWZNs5qJZ26JzX2jszvGJvQVGdRbqMMvYrd+C12i57CxPRgCl+E6b
hbKOyHiSmh9C7ZFDVtS83H8Hs68Q74JOh8xPtFOVPY9d3lB2Xj5S8iwagpaSpst54LuiXqARRHqQ
GQVAFUYWkV1idMBbwcS0VG6bH2fx8zjtfSFnBFb1rcQIPE9IAz3YYlY1ZY0VQaNTruRPSsMNOfF8
AZEhHQU/dnhSjI9FG4Uz8TcVUHxQZUwMmwW0CUsqJbJWs/QvO5VvpSZjq+J13SxrecNuGN4AxBII
y7EHoGjrn1vd1HeKbU+XId0lRJTlYICtHt3Ouf8lumPGg2AeOpEzAj9at26P5mwsmcNAKgbDAA30
kFSphb5VoXRmxMwmETju7nbzLZkZsZ02mGfl9EE2WeNLqnofWA6tfXBD5I9wwWjwFzeMW/aGPRg8
6c1dRKL8DLDmNNLRVF+Hx2jrnn+hsNsSajkd4jJPEBqgtgxFXeoSADMzg2G/8IlsWjbZtUuNvA2y
SE/DH4j4i7s6w+smDCwsOnOWfokooStepppctEHTcba8xApkRYyM/tHAo0s0PDoj0Qk9ru9M6DTd
5wKg9u76OqVkenntzUXx1lsU2Y2MU5JkGiE+W5FZOuApHeByxB1QyGrWCWTEWgYXwOvndTF4iZmz
g+eBAw6fm6YI0Yacy5P7QnH6oUTTNxl0K2R8gdQO2xqP/hc7A2eOEZ2zDs004bq3/hM6I5i06sRN
A7op7UrdDPXe4uR0oX6Ydh6ke+WBx8j/LF7Z2A+DSXrkQoTtPyk5O2YLoqh1QdsNBlmocAjPW8/n
7SHyaoQ08mgfQoWImMiFs24wQ4FHbbIckI03YrAU1KjPfWMtMhkW+4w99TXyWf85tiNXk2aBhdov
Vnj7J6ikd+3ggk+pIoviCmv/TdsJcKUVxqM2JdZt8gYxstcFnoRN09y7RVCReYG5gVMN2mj0HNzQ
Kmgb6/czEum5nBmQv//57YUmokhjGnVaku7wFa9camn1DD3y3ogwlTZAz1yR8MsRlCFvGDpx/f8H
fXv7GCwWsDFV6qEUyWMRlitG7v5VzqK8wldSKXWDvPlPeZbebes2HSdUedRK6g2vNqhRoXGnHFir
RobquaYj4AP3TiqgupfJ4BJNtwyyDLkZPfmC2DinvW5Sv8L5wrjxBbPB3lofWoqVnQWD0wknZrnU
dx2We9I7Ccgs8rKka33xatf1f7OxPJH6o7MHJMLi7yvf0HVHx8MQsVlQNLupa2oJiKTdZQy0SrWA
elqw7vBCYcaE97DY8KUm+GMpO7OOEuy5qYz/fPQsDe/sgo+J2GGl2AU1L2KwrDn+bTWaIshB6cJS
8krf0K1FJI8EjhKvZVS6hc92CSKEx5qU2ohqWKxA2x9lzcT/DuR3MOpgmK5YQCh/Q/iLKZVfsGXt
hKzXVoffBxUV/2SMVgj8YW/I/oEuonO8O9LNGUVCZC3aR6TrKFKPbzLrJiCbXcmLv+nRyO2vp3Nr
8+fX/Py2d1DmFybIE3AE35Ext6UaZnSI4ZNZ/3G0n8yDqSyq0Zt1PZtKzNlhx1r4DzNHCozm99AY
bbOTzcImdyYOZXwLaoTB0k8fknx50H21wwGmQ0iwqEsTdmdXMS0AFSnF10gMxJKWJ1GRxWn6zbG5
sNXyTgxDUhRtft1IMWtBwyDcjEyivyQia9/Kjyebz9E4AB1vGSERQDdIClJYyanvXRdTv9XJx/rg
9bRy9IluHRZN9u5Bl1z+u1L310FTBYo3IvDTOL665K4wpmKcrWZbEC9zXnePGS1uP82OCVNglNxs
8WFDLKi1XHqDZoNGnNvaFYTYMpVOLeOEwXZah1lcPiGQg53F3L7hElJrvW1X8wtIInhZLz5i7wAr
fWwewEHNGXMUvyZ37f7dTsK9Y1Di1SFbOI1yupvh5P+S6MnX214TFcvNrZvJqwb5XpRmsvJWoGau
337ZNn/sZ6ZUI3T2FjxyhFs821xq2bJAcIdW7kangzkmi0uCxNdL3zgxYkKVHYTdjsnrLMHcXUz3
aAM2JJHJu1t1N92/ZNBuAqHKPaAjE1v4VJjvhiKJxoNfv7ngyNdR7HWrJL4ZjCCj/L0rRv+plyqA
05UruuF6suYjwZLHxQDXFfcgUhlG143tsNvkdfO21exCU0R544wNklwrxP6DB43eck7rHaUZ9M14
ym30J+1B1s4RuQhGOnOFB8JxiDsFPCV68rUvhf/JQ4ERo9oxcRX5Wvt7Aff7G9hXDNxb6xsb8hQf
oCj2CFsTwkltUTXzZJj/J8cl7Vjubj41ci9Vb+UIS0vv6+grJJL7T6gZeBtJF/oD0JeSDx7MdDNf
BxIpcEw+uHVlx3eYOfuCAJua1dLQEflWAsaXWhYPbznfDjVmIdjfixQCUKnu7Q31R5fDJEhE6Qdj
YmvChkiQRiivrAQrVWQ+G3E6BEfDpqQqTH9r+JDx/vrm7PwRdfE7sAMP+I7FZyMMt8fnv556mx7Q
bklqxw1l21QIdDh6xylenIL9xY4c7opUVMhAVfSDQ+mqOwbUqSX4A1L5+ETg7Fpu3aXBSsFlB1d5
HIOPX3B4Hn6DkOPTm1hmUK1ebfJ72+h7gBqGVcASZlbM79ebmpgI12jgOSq449MZJ5NRvc5nzAjm
FSJJrllKDGL97zf84wS5G3jXpIesYVOywvfPPcG3ZYada4lrM01f/rsMXgkW5D+3GII9uwwgWiUj
pyL8Dloxdgb1IqzPz3h20tXp1+7iCoq1+ofGzqLKfXuEvqMeLaYutRbyvX0N1OL0MQPs6+Kxemmt
Vg7SkeBJVL16+Ri1LN5LpDWHD8uyyk7hKqjUPhU0O6R9wLwkqqd0jlbtPeDPrWKxUP9AcwEoekaE
pSccFbJKYe9Xc5wdoPUubICmbX/VA3FAl1Go4fYk+VSSqvAIWixzsgS4QAcjdbOTftQF3BXCCz9O
wjZhHUmNYccy0i/JhobUZEOtJUJ3AwxSOU0QnxtHYyXHp9ViypuAkhAiw4g78pRo8pCIby9y/EP5
O0iNTBbjdP+UmeFZ6CXkYJjNbc9CSOu024dDBflvCYp58IBERsIrwfmU2AkWqpsoWaaHAp2hDYCG
uFGFdP9an7Oni+/KIj0IqQXYSCWKGStVxw7xk1wKFOCGDyT4t3QHIRcwGawYMZSxjzYby93LzL8p
+j3KWbNof9I4azb0cuFbSFDTFrY+HN4QdWhTWuEnA19KqnUi0VH27k/WT9dxhQ1h+aAe4mWYp22R
tM7ZHtz/WTXN5tcCi2kB3paa58Nw6JoL7V1ayvwVdeU3nt/02ZI5q9rIXYZlTJjdkXPcO6NbzQyc
/uDhqvHBJZQbLDoalqiKc/s+VCbybQ2Wh1eUXyQsxq+8T0y7wivYauEcm4oTb8tNXQBP4BskBZ5v
0JR6kZ0n8J8cbihZckboyFhY2/x1bLyllgfkXEVTCq2/Pxy/hra1EClORijW2cXH4dK+cYnq5CJc
RY22KqCLrNaMqM+lzCkutuQO41jsithmD4IzSv9KZ/FZ9VL9wJuNXtXN3nJiCnluJoUeTOwsJofN
rmMRwGFiGVtyBfrfpmJh0BeXn5mqRUZUVCYynWTX4qPgAH2Lb+xW40mAnf92TcmeD7rA+yESgKwS
vMKNrPqyUcR/uW6r3Sh5lHp2uo9rDZ7NxFu8hAQZ95i3KZq51BgaHcuEdr6h/yYtKHUa/EYBwnw0
du603x4HEuzgEzwSqPNsOE42ROH4LYd1KnlpeE0Rrp+fqHoZ2f0tVZ8sjqrJYVgMP9d90wmrEYFg
VSJpomzuZu4foLyr8lk3aC444PddwOK2eCZQKUXj0h3/2sfgOmHzaxXdaxTASCM0yIgIPZHS0Fh8
zPx8EMdTvhosbO30KOx74iCAJOaIAM7oySzUyTxr7cZ/HHZstxNr6EBKbbU6/M1YnykzwEDewlal
QYRQYu+RxFTFAso9yoxW0gx9/I8q7xJr5a3bTHEVBJLOWyXwysYHow9+dW6jJL4emxIuFRvV+vYc
JBcwwGKFaGnIXwnN61I67u8zpJ8OW07No4v3hzZHCn7BD8hYg23ayrtERnXudP1Jm7M5t0TgVlIN
+Qt3GBBnTGUMvsXR4t95YWIvhyw2gwAntxH6TbCNp9MyW9rEVV0PZbazu8ifyqHf0qMS8v9JvJ2T
7el+LLxgejc6jXmOtfwT8LnntDEkIO9WEC+h/YSJb3R000XQM7eM9Su8u7EjfzxiF3iNqBvWtkyy
/VEg51X8mhyYlq8OvvhgNKuTfcIbhEwGD+Z4717btDyYiF7Ri1hwZlPp0dOQb22D99GY2WPrPato
L4Dm9QERT4IjZMMEYZRlzgxZX1RLhbXGSUNno5evTsLdyg+Ooym6/lBm8RDftz1QFqVKxGojtc4W
5Wou8aduyqWy2/AT7LDkJh1yWde+xh9C4YsZC2EfrQO3vHOUtlKeO3MIVQXDzrXVsimy1s3mFiva
IxfhvH82Ob4Fx3byj37z3m4gCoq6sU13dAdmNVdPC8l9hGjANpUb7if9Zh2T8l4QHTmyJDZo70xQ
tUBy4BfqniQ0J5+7KlYnLHefcJWhttmjNqjP6Hll5BkDm/yoj8shOOgk3yNAtt2wTJ1h4PzmRETV
aF0dJTykxrQA/DeWfewiprA4zr0+sboUrJ4xm7z2izffODQNIm305yHiSmhr40S811tNnUIygQMP
gUNRNkQX1ZUxtLdRV9UA/bfOZ39b/bQ5fG0VSG5pQRvyaR5v7SrUMBt8DmnVu/x5ZUyRi7YQ6kOx
fzeAGoMBf6B+kGoVeBWlZ1cPMLw50S5oTWpdLFoOzlb23nkPotT4mOrB34xEY4BptVubpwj3zTmY
O9dK1UgAUFk6TNHK3TyZNU/U8pmP4D1AD45mF7Vr4vAL/6AmF1XGEhUT2FJ8EMVnwdHW96Pd+KXW
S2U8gFdSijVoZEpeQF2r3haOW5KljDm4jCD+aCc7bzA1Yc1b5QMgN2HHDqvP54jKFqqwigkMdTuu
pcl1ZWR2o/oadlAxguEPsyDxl7LFLMtpcw7YiDqYdwi7s56DyFmVwiB/iqFtplgcCwm2asY89eVT
czQHrWl/WuRgj9CMROTa0SQACUxb58xopM/xnoc10T/Q3jYH8VkemEf2QTYqw5QLekGShfS1OU+Z
R4Fp+Or4ifNW+6BQuUi+95j/91d/dqGx8wTiMJk9GMEs3I+mYNa/KGn4MUvKTDm8GHO12KtK6dpt
AzyztNkBnmU6fyUJiFg5sIABDA1WekljUCw22r40cUI7nLQITeHUtswxdnaLapwsYVer0elP1OwF
OSH21qohlRl4SHUkxHfzrvP5BM69xVhBDRx9dVIts0k9ioHNvqMWZ+4M3YdTDFsEvoskXjnB9bcI
yOZCmFclrOngH2PjZZtB+MddLYgVxnHJt5DRhxepxlrkPFYD/szKFUDuBY1SiVZn5ICapvzLXD5T
aqfWTgFWJTj/8rEFLBsekxwuss0V05d/et8mTaOQfrzxq+jMG48SV3zVDDirjKf0MFGSFTHZild0
sHD2AW2uBJmAJetJPm1ziWTyXCjNn/3TxwhLRY5Lp7Edab/iQsx8rOsdXsf8nnl21f8ZSsih9Cc/
3dNl+OY0ZLRGCOwQJ9O7y3D67wP8ibZ/hJShpVKXXgND+vk580kkunwi04oCiCMv2+rYUr98Ypie
dTPbGPa8OtTah6LtP3P6bO4WJwz9WLpNASpQlZILrYzjgQKED3t8SCRSm9ja9DFE+MFYYuCJba0E
ntQX3Rt88uh+8pL4KGpQGmZ6AnjXEzQxVNEPmRU2SGUm4n44HUA8hfebEK9pUsYpqXi0cZRCDayt
7yJosUOQfPPYZsrvRMEW+W1t6Ss25KbcBxQHRxLhINQkeFvvlMZUHmsZbR2K6Y2nRS5Z5AdgpHlh
JI+mXXldXOYOT8mAzHNpIthBVX71De0yIG22VB8EE3nVMX6xjOMwDX/7aavti+l4oUcoJvJFsuo8
RVcVWM6jXYKrXO1ZEYe0ZoQyeVjxHAl7idOtVXA3nH6F/8sQp8XnwB/rSp8vS3FEOtFRPaQ/fRcl
ztma9BpQXVCHcLlHu0b39Mvpbug1LufmkPt99qbrg+JA2DX3Smv9BXvf3FsIVr+g9ect/CK/IZDE
WNoheb93B0Tpg3mmi3hGm3VXFljx2CAroVP+rjrGF668yLqRkmipoCwmWe9yz/ZqLxUFmvTwOPDS
UYmgb3XLIlqTkO5kQ2BBpHqjojbgTKiVtbM439QazSFmIo8SWwoMzWoBOCR8/qM1Lk88g3lMh6wB
54QXSg75a0ILdJkG0dIbKMVdb356wsa/UmQarlwaPJXUKiVM/fDnE7mhZo4H9KsWOmjN/sQVgvRY
vkeGAwfH5jbapbpcG/h+FUNy1qIyti/BiJqwKOgrnRHTxej90XjUQUMpS2CH/JrzQ3dK6h1vdMf9
DJCIJa3gzwXp11AFCRfen+YU7LMc1coaz/SKangLGroW2ahInFTm6v9AdYO4Ri8fj5201WdQh4F1
oBHIpRSpUV6JJglkThC9ulTZkIs55sc8NUzhrdw/5FqHK5LKMya1I/CKdYpku0da9lKt+FDkwMN8
r/LLxwzUfp+Ye7zNTsfbzWoR9ywdOw2VvyAzl8IPuwms0Rks39kdUG1Z3sAPVEw2Tplexz5UDrS5
bCbPNRl0Nvn1J9yV/cM3HGcHg9mnpbJ0IoAYAr3XO++NZFnD2LcSzXpZEBmaPZMRBl3SXweGtGYR
M+AlbGytfUM/U31cdx8kZ9TruXw//A2k+mYVlLXL8eh5B9Y7SVATF5VU5ooi7mr88XhYWAW0O7v4
8sc2P4/yTXICthynAi5/uYq9fVBqfvWj5XdRwvLSZ/CFPd1EPANfdDIQtqOXkwMbE4f2N4Q7yz2I
S3cTRHb5JJbYejB+9S2BChYzuHY/uBAyFgbWZIgiP5n7pTQ3/gW+n6fgGeysmoC9odXerG3utMnH
Fne+pWoOLUFSMqoY0DHCPmZSM9+sg0AQ/ohPUgH4TXTXKUT3fY3JvdBjnWIrF0aFwvOVW6bdgDEr
cyr2687R+8WC1lUhZ8UVoyKCZrFuBqty/pb8bfzvypLL7SpiQ2KP1S+FBPKzuINbU8XIYtz+pjI6
1Nn1z3Z/3OtWMUkWQZa7yUxX9HaXISZaUu4vftOFSAB5LSFsEgYyZjpBYdMHP98HE0upHvvPnqjv
u29vgqjAvPd6MN1qZqB0yT+6u/NjMxXJwQZoy0dU3F+WTGLMC5pKTs8jQJ7TAmcpFAOZ6/pgsP6V
QsdydaiNAUdJZGiUCtGRmplPbI/oZU2KhwWCIEZK8oIQDad0XiHCYuW5ByEQfF1jv4KrgYQSrOaV
AowstSM8p0RKqOS/IGhOtoRBfDjegHA6KG1f4WG0lg132YFKXZ0dtFGg/IXNcREKXxi88v0c7Kqu
EpXgjG9gLJObJOqnydecGN7E2bTmlyE72OEYcyLTa2pJtb1YjyBclAMyF1x+smnI9kWekyKrJEcd
mg9kvMRfyG2lOtLB6a8/U1U5jB8gHNwXb5ElOaLrk/qk/th8pgNqtKZVf9TOVdy3EqiBmUck8dJZ
TEx+SxCjRWWPS19n0Rcr2JvORAFbPunCZ380QNXN4Vi/exS1EHgBAjSYYL4LBispawqjlZkdmkpc
LB16M4HXdO79z3IannHjYsKPS4hxfmOYDiQgD9MM8bNHaZqBIeiPnW13EMiodsTgVY4LoYelzws1
71YV8Ag9qlmYFMOKTz8r/Egy2ldYDI5OIb1gZeINsMByCSigVeVc94q9J/RmcjJCsHecoOyg8bgh
Laf7Hq5yzrmXTlilhZfdwHndKWTTYL5yPKWH1qvZkUNyFkjdFL+pWp46s9Dy3ADVQiN4nw41PytR
C34uhgI7nutTqj+0w3jPSuId10R2emmc3M/vbt5AWy+mQooJBuXx3jof9WgpSobTPtw1cPzgWThC
vmtndJB2llCNeNSF1VsSjq0PELHR9ijkLcCtRiAQSncoF8FTjV4EfN0I7vU3gMeeWYXLpfKa5TIZ
aOk81U3WmvoV8mEsEaE6X7dq+5HwyxmrvzgR8Q/f8azYFlLbU2Cqp2aOvbSGXngl10NWAob3x0WR
6PXNXda7GE3lww7/szwxl6TeO7jJ3p7Jv7rSh9Hg4OawJEbOfeAAAkrep2mIQDv/PH1T5GLSJ0d7
xS/fndJlbEERgf3lwMLNPfmVIcWDET7J1svGCT000hYpJDQD2hiHNLmw6Hvx9tgdKP6LvFFGZ8al
7p4FBfpWwG5fpKBBrk3uqQjy489wuuFab+vU94P09Ip0pnT1Bt3Uw/DwGuYg3Qg2V9jzFsbG28le
Rr1dmvxzaCoDDcTwOdkuDWoiQPXBsTLlNJ7CHsSlH36s6TnS+IgErdRnm8sd/YW23/fqBg5PIfEP
WBRWoXqOHpiLMw7xaHmWhuzpZpXkjJkA+/hpQFVnLz7SbQ3gbwQVS4ndxVeieh7x7nb4sW/dyN6w
btLQPxyL3O7RxVo89jyBuzaxZ6+PlGWraAMpPQglT5ly8l8CDIo6bJT/MnbcFspVfSIpI6GtFKOo
+KLv+BZFQqZWgiS8YfeeV5elPQ3dQ1OnZr4IIcxEKxWh/7A3fJ7sTq4LUGWNhRkY2agv6hE7OQB3
zj8YRTaoeq3LuQG71hKJ0AvlRebt2wXfH3Cr4ZLBEIMSkqmnCwHHKv9znGGJZFjYKAfx8jXGc5yN
HZ0+dMiho9cP6BH+ntXJYKelXnyCaDPZ3f0KnmVlTaQ0orr2nCKaXp43c0HaLam1VJJ+L7LN8DbM
F5wHFWN9QOUabzoogDxMTLjzrPpt0F7JDoN3sW3ISw8rKeQSYO3pENhl8+mWXnk0UKACo2QkGLs7
hmo7WqObRWQoIeHS2p5aVQPritUu1tZasIgPImZN/zRO1fRfDAl4rPH8/x4pMy3sPQP49pqrcv8M
E8yHPWr7UTSTvE7mQau+njfVLrn7befP2SGCKWMFBUa03LY68iuksZz4eOQfZeDkhw+GEDcIU3s2
xt+j4D61vKFVJ0nRK3F60gWSMqAmeq7U1dbS19ZvjrdlXpmJ+LSFq8Ha5nMLxfGuwHHsi8ou6maw
Ki5rok9XRii+Vf5neHdiR0FV8+eqkpzraKD/aX6rqzEERQVGFGFGQbe7q1su+zWP0hl0tcAkllCk
RYeU7+Ew0+3HWAxwAwOyCsuO/nQ0wPqlBMfpkIOsB9rs/uY9kdUnZzsTOiRJldCm7++5imBLm2/w
2EFBSm1V7QY1XxmeiL5aqe42RSjcuEGRZUZcLD0U3h0YiEKK121tfBa9Touh4zBa/JDANRol3Hb0
afmjUNwH0PDHQvHfZelqKl/Udvw/0WkwHVqw77wkZmw5xlW9+y8eoIbiJn1Mm9NuYqE+j64uljO1
r2frhO8FXqVoXdYnWkD5jyOtJ+ALNdN//G339Sx/9xdquOfRWZ7b46gO6jz5w+SnRloJpLRFJFtm
dgstRQNL7y+r5rB9RabzVqeHl3Et4vYOx+Ih0LBgGvDXBTe1WaRV0/buTONGA10y309oTtMOZlls
xzaSMaFyHRhjuGYHS3rhI6N5ANsn+Y/Xpt/h4KujaIWE/ldWjR2KioYAqiyFKBpFXbCyNvdkI7/s
VPWAs8MAQh55Ld+0SGiaFg7baPXDeotSWUl9qFTurd9rhWiLmgAL5c3A5ew4/9q0DaqC7W6L00AX
OOjmRmDkaxWcpGRKo+HJ8a8WHS3u4+LpS/qU1Sczu+7zFw9+/OrU6pUSgU3rCe0pvuwedhwBafyL
p//KiCYmNY6nAbpN9c2/ETtgmWoU3o3xDowMOvAYCWk4gXMhhqBJBv4Md5wP8plcWnMX/1DmSK3v
BOEYo3DBZLrwn/RNlBPiZswD+sfyvdgFdNI16luWD8ZrQ3w/yn+499zlrHTCYukvpEz/ErwKtm12
uLvgiMvRTKFTPXveA/qT4I1TkbYRW5Il6pvhwBuRADcrEU89/7k3UcgK/MuxL+f6L/haPYZlHJJ+
7gRX89umMITVIDzy9Me2tCrXMxSztE6qxfd3J4KuAIAUgiD5bQoEN2Lx87/rVhCWFeGA1jckU4uS
FdHckWowLKYJetsewvPpPB8zYzcRc9lfjTzuddun0ae901AMreW7GrgDylYCJ1bpV8blV6Q++gSW
3cyPbFj2OoSzkIU7qwXg18ZTg6T+mcJ2xwqYOG3Mz4tSlvulLo5IB8rBTmOkhYwSjiS3toSIdK5x
JaYFPuHB4CHrm5d8pN1xqZkwNENwbIw1R2Q67RNKfZQJSvXdHI/HqfOg7u2x/9WqIgtUeIWYgdtM
6NS5osnmhW4vZJSOIzbxqPE6bhpivdH12c9+lfX2VHuqzOT9rOn32KrIP2hc6a4jTT1lyvYvpmMH
oLcX5SMy/PffJcJw+FjYIrYwC6M/qR7El4vj9qxYS+DTCXsJGH6Et1Ff588CUx2Scw7fzkPKVlMf
nfSjCfahIGXq5wNgtKgf1zhch6POhL4sUYU/PLsc+KNPBYjEDNj+RqCDgvsD5ULkpor5AYFoXsv4
hYb2DQe7MOlu5KINDwd+SejNerpoxfOHO/UQBMbxgaeBRDE6/Hk7W9L713rP2UqHimy61TOHJBhU
EkHz2TIxRFeAeCBNNcqNuT4nFIOvEpqBgokMnH51O0EImTI0amcqi/WxY9A3H8wNuSFig0Pdkf9D
fM8YTS/HXPsHQbHheMeLP3A/LrWklWfVNwpbcMaM1XZGto2wz2NweMR/Bi+vhY9DFL+C1Xyi8iDr
hf9YUeQMiMlTEMtHlOwNkBtpwokFgADAF+sn/sBF1e8z255/fAwY1WbknU1IbUdGb6PQxvpIymRH
ghbZXeIk0xRfyQf+62FVX19Re7JzHFgx0FE8kvdBhTuw4wE0gQLIOpOD2q64DgPRWHkmfvZWBaXK
E0y//nLdWHNrsu22DY15OBf+YEZZL5yV/Y8H0ewyWHVAXk6qMqjnh0XXyqLJW+ycnW/yRbCW48Ga
iAXJm1wNTzUw1vD3pomFkp9kcm+KxL6b8FaDvYX3lc7p+q/809ninNicmY2Ltm97tTcTtDJNRBjS
5V7UxN7L/ZzI11tzIaOQ89x4rfbM0x4KGPrUk/kUa9dPrhS+1SF34R9FkPWV9WSKC+sj9SVpQez7
UUsISL62chu/MNQd0gri2pi9epxaw7Uz8sE0ZB224Q2E5USQm8ic6ptnspVavGQcRdfZC+1UHdqP
/zSpqbGJjTxVfppnukEmUkSikcdjlnM2NDwdin8DmmqV+tryQH3tB2Us04j+EgwXRe5RlWptbXwl
VKyt6kKfXCpI/coiDvMQUtkmXOQqjcxq7FhEEVi9i+W4c6M8PU2JhtEr5FmNfIKA6Ijm2Ypj0YCD
+xEkE7QkxDvj+bvWs2KWIvk1HWMZmCYH3qyWdCDN557X0uIJleuNuxlTOiD54lPSjfkoF48AUOMR
3wuifsw8cw+8Ig20V9gAN1/Y9S8xPDJuJ6VQy/iRNKQpeHqXeiD4ynSN6T9SO/NoPqSlOwaWXBLq
m1rtcCdxuAI3LVs2ZNWbPyY/bRD91/MHeJvZ+yrlTJYUHzKCrWxox8WK10K3zeCs9IR+gViXzaAz
1B8aqr1Ul7NyRlsCaV+2+vjs+OAGc+bNfLDIPYhA36xJSd40oi4gCiHiNF2GsAByI4eh8p2T/mgn
JalsdNPohi22d+Kcay0sjIABH+mniW1y8mbLBtN6Uofh6iSdYrdMEae1vz5frvEi5NxjBBcS+bqR
BvXUZVt+cZVVcgUaauwbnoOAPxds1R7nfo+FRhFwBbNZQYniQpSPzA6c0tooEjVwY7tIUWMf2bpT
yBaHB4xu3pDvnrwto1QKDH735GpD/si5I9tEbT7/5swrat71vwdYVTfhBMYiMgK16GXUvp4/qxLJ
TM6Jmdm3GbfE7oqH1PnSmZeuu11v6z2xLHm0FrvnG0j1wBiBxjCy+GCwjNOlT26Uix6i+usWc1+G
DjM4cqCZ/GRxXe1XM0XjL8ho/CrUUfsXziwM4pvmi1vKIMox0E1ARklMsBoGo7LpDObzRdY1ZBEK
eZM9XZi4BsWBd7y3WRSILnNuF7WMd6b1MKoMmK7lEnF9IZ+ekizzvEnBXs/b+tJuhjX5KfBCFBqk
vVdaP7KhiJFO5sd6SNaNi3oiWa1GrsnbOeCgLCOJDLYGhUcDXbE7O99uaelYfC/u266HSP6A0VVj
nU7EKwbU+K5algSnrfqq8930TrWpVxt6SgTp7fbvY9w5+X4pUxFXue/xd1IbRoneLhMm+h3YA4on
Q405BPUF82vQtNHpgIcM1Qo0Klyr2+YnixpR/J1dheFET1LFD60squSZ+HH6/pR0QZRYZK2759xU
3RZQPtZYg0AiOIheTt/a4pli1gz8uSPfJx+mJdlECuNiW49/0CK7Rbio6A8hj9H3Awmud/YfJg63
S2QUNByA3ldxmW7p5eZum97emDcXGgtAyJMtovmf5Og2P1+5T9gftO66YqM7ntQ/pNbo1VzhpsPD
fXBQ48FJdvGX3VtZN92Jvse+C6GbuqrfqG0/+SJDjSH26dbRK3XHIGtG/USou8W6oTpzk6yGMH88
1ZFRGp08N9LrrfbyRur+sAOwpZIoWiWjBrcqIF1RaSJc1+DuenR7JAfYf6Q+Pr4/EFjRnBVGTybt
8ZM+0j0koofh42NM9ByoLTgr3EjR/GtxIlKXuq9Fs2fJVxqkjWGb6jFlspQwGVhGtox4Y13wPnY2
hoU+ZiwFnRL6d3cQ3g1Lts32SKuIZQ5Hf9Tc/8NACP3nI0JPy+J/QG9S1qZenkC0deqXzNJKHfm4
wSXrRvK7jiDBJ6xrhrbB7oYvPKIZqlr/MxzgTNsiDfcqLHSMOdiYILX2gzOQa39gv2hD6rZGgENE
2c3gHhd1OlFThJvOjSQx6idJi683N460S4Le+Vk0OApI+MHKuhoi92jPAXKM01DRj0oqg+aA/FEw
XODfQ099MNw1VEdb7FH0WeW6GgBZyC8nz5Ros/fKGy2NsF8NypDBtPcf/5f1Fhmcv6QFN9yUjrU2
j0jfVAqh2N0TNt3FgKx+0m/mX0Z+QyFL0bFTXjgIcAVaLwMNKZJ+sSDDqgTzx4isNv0qG23wEoZj
gJ1WR1w5wVg7tDfB/mvBoSCUaKG3vH1FAnzaWSM5ExYZ4xtqMMrmJwYNriC02jTduizAx3ZZaJkT
18sAaNsNOE6xT1iwMS+bxWzcJ/8DswMR24NhGNn37c8xNnRBSaxLdQjJwgErHDCEauHS0wxnF8M0
9r3KoKKw3JjQ8Eg1QNTrEaBZZ6DnhLgThDlXMtQy0g/pCmXn9xaN8b8t3hXWwXdS0pWUZbCpWIE8
CXhy4JhYcNYbwgHDdIvlgGVz+14ZCL4rHt2nHDIO3l380N7UriEm1u0xASA80JToeIKOTYu3+VM5
Et2H2SNBThgpLvNcRxAGwg1vK+8BIs9wufXEPQBsIIQFQMyvvs+WpimeDtxTTNMYRWO6TXkv1g80
87nWigQoqWNdOtMh2AnStqffC4HJsgFDeZrAstKNWKcVpaIPFybXdhN3S/Z4jwtkhU8s0kKPhIc/
hbwa/UUolEgXU590W+cqQDKHujmKQz/yp/JBYDaTBxFd8E6Gtl9INeP7bGvHQmvuk4P4Rc4RsRix
p904poNavCgcAiAl7xEXgOxLsEeH4LxU2s4pZEwLmJc/vlGuHEwhaBpOIabQUdPZdPVSJ6SF0NVc
NmVBAsAfk2v1yxkCiCkxnAQPbtyI/jeM6EPX6czIqdH9HdhjAN7Bupzm7kWzkSi9sHgn/rSVeJ0S
uOnVo+kaQanVexH2WvhHqZiGfGj7w86M4jCdICapK8M/BZZ4SKl2Q5Tgr8XtRi+ttvpTIJkw3/oQ
mE5y439cUAMcK4bXI59BvOC2uA1ubgmPz7NxJukLWwjNKCcmtEemcAhy+UUywIMyk82dJEYCWUyC
YTxRafTqU0G2DGUo5mBg+ayykpnFCgrMM6G5rHJJew1cb8TXvZEBiiGefCX+PcFp6CCMnBbjcUTh
S+r8QTvxlGBYYrIrAvtAyLkSobwqXFRdlKSuj4cCj9uzY8ZFdXRAq5ON43zR1NRt8soequORKqxY
0tZp6kzrg+NbIuZn9wIXFf0DORkfJDwiEjYp+1wWX/db+ujbRvbx6FLZ4nrsrHsJCwob9sXYrxgb
ZWiDmDcxrcXwlh+HNI1aYQ7au/4y61Bw2Efws/0su4g9770ZF3Cg7EmKDQF99F6gnwDI14XQBahJ
EKSdMjZOWU3Lt7oHthUrE4oiyJ6GfU3JrnHttTpLlgToS7VLrGEvaSbOTUZ231xJ5wumRQ1Sr69Z
CgyOgEE7fCFURsYkWjbD6HrCRujVS57gRMppbaoab4TGhOxzqB2sK+v8b0PKUAxJQ1sQw72iRO7T
AT4jMXV5esKaAYEaZFEVuLilS0KTFIOxSuMQOP05vdlGjDuoUWjUpdL9F3n7aY2jOW3lQcDNH8lv
ia65srNjRAmvMPpUDwdEtagQJ1WOp3IcJf4i7mtXW3dvBtdl45EGvBA5UP7TpkKvNh7gIF0TBSzN
jaK/dV7z4kdWLmOy8dq5IINZp9sUBO1KTmQCZiztbwzUSumrw8n8WSQGRBdwy5aKgvOpD/O4Bksa
PaiivT0TtPChulLhm0LCWmdGsIuyTNZ3Zbj79RpmMDDl2rSieiSMxK+g873LDEeqygHHkx2fZ+eY
2QrH/LBOnyW+qBncZP/JrumHgwUJ9T/97SnWM/BQ1MjXXeSbCwg9z17o+5Y6upFQ6ihv71L3FT1w
FJFbj9cav00efoJl5GBOqqsuv1N2F+czEyDNFhm1tDAFIaK8sFsvDEqZo6Iuc/dUKIfC/JkXKzs8
i05+GC9osudNqjvQA+ERgoxev6MsKsNueBQ6xgpWy/iqqPMMfLkXlkwSQ9PaqtA/LwPEX0toodhC
rxsuDxG3T3hX+ikfnbUq252mpyrxYWEudIcjUBhlpDJ39i+bwY5xe4TT4QsmV3VT33y+6p6D5YKo
8GNdC+hGhJdo41LDjlIK4eeAXCXHQWP3cLJ/hTjMShnDRKHYCismrf6A8RIJ/u3eiE2SK+qGV1SK
dNTiU6PSHk40qyegWfjasx40CZ7uvkW3dzfhZJmsd2ydyw6BbOH7gIf2r4qCNs4rO6wkeqEmddp3
fuv5SLfFJupcAlszqDwAPkb9M+pAgmMGcWBaWCi5cwKZAFwUg0zpYl2JI+vBc68mpkEF6k+78qmA
XvWY/FK0ML6EaE+TUOAhkK66yQUeB5jW6ypxd6YF2djbnCgSkUuV3K5HM9nATyOWleHS9eZIeOqW
fbUYotz2zqPIW31zNEqsbqAK0MIFDUNga38ccxMAp065NO4Tmgg/AQq60exAt4/Cemop2S4rM0Ci
POHhS6GzG6jEo9wl6LLZX9SQG8s+DVC9KHRTJCRCyDk9o5//YWBkBTmuL5X+QsQ9//klPPEmtdwZ
8iuTA/d1+uEFNPLsXN1pK0SO6oQWd9sDl8RJAM1RUnrpMP8792a31XLi58Ee4d8eY9c1dgN42zY+
3E7YRgXdWRYvu6Pa8foMt0y4Q9bOCuu3capXUC5J9l2Ga1r+NsSZfV/yhMC41O2Zh7s3HnUuHFqD
hL2U/WhbDjKx+AAvoUldSBI/0/eteSkgzsWi0jWZF+o8sAV0QlFr4d8ZYQ22syrMphtobK158dfQ
zlelVkbIYiAMgkgzTgSt7PJ5x25ixFYkrr0CkbaeNqfD7SmHKk7Do1VTvs2pOLKntN/aQlHJegbP
r88axuAKShy2BM0A2L44gc+I48FMTxNOak1YvCVSgnoxFdyFZHI3hTb9Tg6pSy03qybhLIunsIsi
aTIUo7fN7ovvOmJ+Ice3mshzHqGxVUXym2xuyg17dN66IiXFFOLPvCFuQf6uziV+GzwAswBlVxBE
PODf2n/BXYZtf/Bfio/MNW/Ys8+SddiSvpF8kknFYXyjBSjIqT/yTUpRKw0eXS2HuYEWdX3DQeiH
YNd1ZAgoHX5HMBlZsVyCpbZyrttxZWIWAX6ePbs6q3Mer7NZWPw/pxxMOfdvGrQnAy26PHqvZho+
GOEc9O3db9M0nv76nDs7PHHec9xndn4ukaY5XAYL/MnGII+32tnVXnTxK/OxNtxVq4+959YWabg4
qzzdwX1zSLnzk/y65b1OowPT4G/G16Nd/RlqevBILNu5z6DLgUioSBMWtWTnRHIDkrZoakIFyJjo
o2sc9gQZqPjL4vbAnSYe6tXCH6XzUZDyAY4K/FtBS/uDRLVKv8+/LzrDxG0968A/8c2eXK/YfMyH
PW3ETZV76R9jBIblkZWNMEoJO7OwObTJCcnyLriWalKUDFF76HR2UUFFhRUt7L7OpFeCoS1EkH7f
QZ7OLWpFSZMSPSl7OHPvNLnlZgs4frUe30EpQkLrkBdAuHRgRODbhr9xrIzgyD0nugy25zzGpIkZ
2JNjyVTqX7K2iiw0A3ohMz4EYr8pxwKT8/ny5qqkjrN0kx/a0UZ1DfT7tMzVouHhsd4pbML3XtFq
r7ujkvWdewXPAs7KSx73ABfrs8BOrommyr5LUPR61IUHzvE8+jabgrAzAgzbTRp2uDgXQfG2tgHc
JBvDK/q7s4XY9UFI898lC7X+Iy0MQTT+AWbS7jEduOTL690pIbsNXPmCM1IjIfIafre/ldpFTZiO
97rzQUPC6NLexOTzJXPL485ErsrW7sEekpflJUW/oHpGGbmdmYvDz+6GeZAJxUARzT+RKqJZmoUB
/JrUMyei/MnkJ+fImIoaonYCo2+VWjJD/yVt0wwbLSWL0piUFXIWalf5GabAnqjUvprtutkquZjZ
qccfwRR3N8opBFno/MDelJ798GutqZyXnRf5bkkacwyW0+XISimTjtdVHggYSEOSQ8iTT6y4ELzk
Yz21ZZ1V+dvIHqtzn7IwBw09QMMkV/wFDQcamKzZEfCGFAeYblA76FARSL9cbMlicIf0uhpAXqAc
+4r3s4rUkNLhox6Kl7buqOEaw3SfjF6fIxgjQzrHhJ1NV3RVmxBE1gTo5LqNqggcrcRsYwrZwZYm
TIGlYVu0PMADc5cZmXoWmcVZoMMm90M2fosMiYyjn1fR1Ra8y3MvN+90D02PVBvbs5JlWQQPyVIi
v4XTANWom2Dn/gkH/YpdKYVjYgWLSAgY2LbQWKXht389HRqQPFYHSuc9unJy4EaS7e0iv5a7I0cI
THdWd4aLkHiyKn5pgzSMNtWHms1Xq1lTD1ojPXAuBFxVoThNGVkiXjD2MKTHdgI5d7S/eko+peAZ
9LMG226nYuAjo8Jr1sgDh/5NW4yToROR/5M5mNzEjbE9d3Ekjufkn7QI14hSUst85AxbKgV3IOxK
uyxDQ0lcDjjwj8FSQX02AV87IRvAytDsMjCO4IdKk1ee/Oi4C04V5sgo81INIybjZKGqBRRZYejB
cI1AxLSpnn3dZAzePCeI6T6Bl6h29HBxAaifZSAkhJSm4W1geR52bJLHgdzTUHewvXS1pDgLo0J8
2pzSIShxbxQ+RhuflMFxeyNIBD5CR9yHnWoI1uGsdYa3PmVbugITWQO1syrsfU8Nnu1o3nN12++c
hlFwO+nPXARRKyD2v0kuCA8r6COZWSMgxP2WMRdrsvaI5XFFnmy+Jl2x7VMbrjvEul5DVyBDBSKu
HR6VBuJTYJDb6whZ//RX5XjsblqflrvEA9OOmmTCtQsM3+yRLQQ+bPrgPkJLh3zCmiavEAY0iHTQ
UUquJo37dZegomZCltMT4PpVNHaQpT5BzcKcrCaWHr/P84opbtlchTEdowA5+WQrWM3lOmOka5zC
qwTAhLmpSbOappWN6j8Ikf3yvDNRVj0eKQ==
`protect end_protected
