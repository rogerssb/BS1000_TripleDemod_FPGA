

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
MYxa82wIOdtVBYlwy4/Q+gWfpDcqU9LOv+vAXX+POwJQnILHf9GLqGb1MA87bCBrfiBBU0yv/Mz2
PWB4gnNCsA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YvhMY3cw0yDTC9muVdcpXe5SBvg+YkCe6neHQJW8HFbhamEt1ykdxfBkyDfp0v90qgpAUJVj2fOf
33TJkf20IvUs5i4GLE67n4KKhhDy14jYn5WAeEt5uSZ7GTjlSXhuadWiIoe2q1lkKGe1AoWfh/1N
Sr55/KEs5RVvnIvsU+8=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
h+VE5xEgbKgFFO5KK52GY4FXHBtgVMC1GWByYpGZCxXDXUBFb1MHRqDH9ibaUxAO1zWAyx12Us6u
kmi0ukFDXYm4TwCPCrJyJv1lmp8BBgAs1lDSAl4KhOMz8ZI6F8t19IFQWy6EjvVRxXPDYqwxROl9
8Iw9mbHYMTgkVXI28t8=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rPan+OyqpJHTIRYXpbG7IXln5NiJicGHWWeeRCSCHPw29b8ZqhJR5J46cihj7eGwAV12gP6KZ4lY
HF2VwPW5KAWxoY7FBD7ObVBGyQJHGxarb+v2u1K+LsF0hTaG9WOXR4BSSW1hPgpKuF+Eb7mj5OUG
4K4q/DE/TKs2YS2fZwBNbznVvaD7cnQXU4LKI+rFIlKjUJrws2fuJhXFAKZQpyIrV4gQI3urA8+p
R8SYPQneWTSlc2SRP4ppuewpaTJ7jDyYmcHzJgrzA5iFGRKTKlFQbbiRfzClNA2Pr3zVPSPEDu3m
CQ0qg6qrFk1/cEB0RluL03jNEU/ewROjWktLzg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FTESDNXPsNu3Yk7E1rUlJEUkxqgHW1yYULoZLP64VVuoX0gE7Ro2qqRUDwauaVpPTH6G5tBeWbeO
lcLOW9TpcGCf46C82wqaLPuM0D3OMS4E7Q8DFyEa7QlqsYK+ccCQXi/Z+lPV2IiCeGHbn1Wsezr1
npz0I/tjCfeQM19xJjcg9D+xeZOvbgRLSvNjqdASD/UdDcXDKm38HP1Yxgba3BFGSue8AgThpmQZ
QVeQJCq8ZO5bEKqK52J5B754+dYVcfeOPIQirUzNNYXt0yewztRfbEdUmH4TqIbw9lfyJCxsEK/w
sfCLEY9QmULGJ9wWjHw97jBnuFWfiB4g6+X0Jg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
w5B/y73SVX1HnEfEDAJggjbtIJ/M37U8f5iD8eH3ipYIrJ8Iih1ssqi8aRUBvbljYmWDOWDO0UJF
PnQ646O3Pv7t4X4LLMMN76Kap4WM7hlajcJIM8CVzVeoXIGkcoqtsaKSGBAcR8gH6vQPCJDL3zXV
wj15rwPvS3VnpnoCoaRwo+MpNEI3OY3x/BEMg1n5sbr60yCqK65qXSNZqG5hNO71gEPnreERpPsj
0+fpKsW3eDFt/QjcfLTFy/WxoIBbGh9kwOZn8Pr+3U2v/elDSvJ3sBmgvxrZFLYoR0d5CsKDKA3x
zOMm8RzBf42d9hOv7qsY6X+mf6PaPoEPVGtn3w==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 99168)
`protect data_block
vlUy5cIU7tONmZhhbKyDMZhEFbI/XDPOK+miMXbjLxGSmcVk8EHYpMutCwsJyeJ4VrCUFCS2UkO2
C8gi3DispHGKn0XQFpwMec2PxeA9lYNEtwL51SuK2xo2fBqHoak7e4uzybgEJB5sN32mygnm2VHC
5PY1+hfQeBScBaQdHGWbEv6jXCoQK3EXMJZdsNApyIieJF9Ae3bJXBVM0MKnr5Kej+WJkOtdxpLk
TnTmnSMUgu6nfLVo+JU1b0qtWhjtuWTFzdlRa3OBZ4qFrkDzTkDQJLWxHd1S3ul1kX+K80YIGOCw
5M2ghYdED4hWdPb7aQjVZ0QCU81rQgu8nuiGR0OwK7ybvHIVPe2SbLapYCiQ9Yg0SVZe7SGJ7N/I
ZX5QP77TXf36nvQaocAU4qBpBR8ONi8Qw5HuCIeu/E82F08u+auiVpUc1YsEPpswmyG5IhZDi3U/
VIFaOI9/eSY7vjki1bg14sJTFA7rEdpKagUd4m9vwc0ZR445OB5BZmvO25IiBUHDDslM6RjdEeND
b6I/QigROfr3NuKp0OPSkKTWI+QtfCbSaVGYy/D15cRQB0DhYZ8Mii5lMMAGS70icxho+FALg+I3
iu2Aa9Zy7kWERS7cVgidseJL9wMUn8NrJR3s5GtUQzLDLzzaf1aznfZ4JeKCXyuFUqmT20A0Aocx
4a1FyfAiVR9ZvjcVC2G6wlFYzrYQ79Fry8lO9boRIiu5THG5jKvgf6ayyXD1wZN2LcNncXxzpuh6
MshH7N6etTXYec6S6VeNshu7g752sWlPSgZImNR0So0GS1q5fEaPFJNawwMMVHWanVJyGF+vpcm8
nkn0KDEC4IM4w7VPtF8FZAEhKxM7aQx8EmGfJ1lSrvol+uBV9PUwHARC0mJutwIuAoLHlPWvg0uG
hqUkYzQ7WBIZCCaRsYUriDwrlyc+PoJmVGuc6NMmFG+PSNSrHhgfn92wfs7GubRSN74viob2ZWGq
qJMsQSQ7HiIhOEGHsxARf/LhtdO2EUu3d0AKKgA5ODc9fFS/SQ2ZBBU7INOjWZ1AeyO6G5zhmr+e
f/I6DeTuvFeELuHu7ce1hNbXXR0iBx8kKQJmELo+2+Tel0pPzhCt02bOwZiNFn2Ppq0qj23CsyL7
VpFI7XNXDd6VWFp8RVBic/ivvVG23Nv95aaX7YD1EkpEasf+fioqA3j3Ia4kttCc8oUkwQk1P8ha
/m59zBJg4vdTXiP3XlRiZr6vL3/WgltVJrb8Ew/LqqA/g/FNwntl5upJWCbcf6UbP+73CI6kiH+5
Uo9MeKh7xWV/mF3JUtPEk1saYTTjCuSkyes+DDtnA+rwP9kPPmun+9Hi9y117dpkG/6RxYnw2GDP
09gUDjlZM7NfMaibPk0lXM79cLJB4kaQRj+lESByNDJv5xmEralPlamAkGgBX8rsHs9eusg2TTuc
JHPTE4izeo7FjMKZ8pqSC8CYdCbs6+yhMnPAxIL/2f/pidsSHGHCqGnnVkNYiaqPkPPbCqOrenQZ
ZWeNB3B21yjZzAa8M6LZCfgx9tS8dt5OeADfotlfKJpLWeBXSgEZe0Rn1gH08Ico6rcMmzRIQjF/
l+z/CQ9o+OciwiVz08wrQRD1t47C++E+b9z3r7aJbts74EwAJ82OzChlIQJxD99vKr5QfgqavHup
/4E0a0hDF6YMsTfyRhD2+dbngJIwGkKPbJ5iVVLG29+nsin6BzHS3g7CphqRufWJL8TZWRH8o55S
czdrxc4x0qUqq03sRAnZ4KMscPBHma8jip8BbmbI38K3xEs180EInFCyH4br5gtJj/8CrP+9b503
edX5oJkhVQU3puzFyEl1IuGhvzeMAojVcEbH/6CUskFJPT2IL7oOuzwFdO/U2tddWbMrrzGwQT+4
U+X2qZ4Rg3GtoUOorzAVwZ1BYmKaFZTQ3Q/X5oNR0JFivhTkL/p+bVQGwjtk3QlALf9MvdWpzTGO
S8SUWZMP4N8StqhWr71zac8StkBNt4m1XF3BQcOztIPrWkDphUpiqGojqJUTQY4J9c6tTcK0vD3q
lhBN/wCo/rBZFScxaRx7AMAWAFLo5184RRDrSsncby+cTTjHCNit9myHlNxwdetPHd3evdEOCFau
5KlrNyiL0FVNXathmIcPl7Wl7Z6P8KUGjVHOfSdj3sLNFXqK73ki8YgvechBmwtkMbeQpAqjG4Iv
lzo6wZUpiPAs67aRgoobT8ZTulbT63bMZmyV86W0GbeJoGbGGft7iIqflic9BAy8Q92UyOLSva3W
RFzO1pkdFcH+2ngEXaOPobxZt8clLI7QWN3BWSZGG9ghbt4rTtCGOpkv68moz9zgUTDWxFnOgSev
VJGV/AEs5AZPoxXMZtAs3FEAEW5w6CCGzO9TgS/YpYV419/VCf22QosdBH91kODEEeZC0RlvoapZ
/PDon7PbjWi4HO/M/1/5xkqzW2E7eJxhx3BO7ccMg2keesVSmTH7FPMng/+bCi4nCW8dXwqo7Qow
goz41KDBhUygvNkg2vLqBuywVxOFLXDJWtn3g8L20FA94TAdqUZkp6eDeZsVGU1ZquDsbRO+uvVx
zWJwheHt1mxB74CUEhCOVVvHwdqbnE5/AGYwMKFmqjVsCrcWMHq4GmaUuC5oCqHam6MWp8Ez6/mj
S2yYfTj0iDeKXsHNaOc+ybicNciy3Cxjf7CQu1WTPwqeLUgcvE0WCn7MQoGggn5zvhXkmFMFAxTw
P58Qbpk5RjIg8eYJPmbk0urT+TVETY3JREh63OCZGyJpZcMqFgiGY0ZFTH+xvAH3MoAPhGOGY25U
1sEJWzDUco1z5sy5gDOL+FXSU730kAvCv8M4aaJNpyDIzk6MQec1Z1DRycRGbF59SjQZ0bkXkGFt
Aqo4NiPyHqf6LDkJE/sUJzSpcbx5QLvLci703VwdShisNMBg6p9/wHXdtJTWqFCRGfg9CZf0FhPP
mmVLI6Q9c1xVIaNUiwpv1U6A49FQFrkhe47slZg64lC8zZDX6/zoKES7M4cqPEgpmTE7v76gg1bg
aJyWcy+e6i9g0qH6JAhnjzKhu4kuwlr6fkz8s+cqV/aLrZRtU6X9nN1pr3IXpL8ENPgTHll+cJHG
ID+lQSY82Z4lvlOdmsGzTFul4U6W2aINz4ppEZKDrHJDAGZhHGhQnc7m3CU67N5+sPgvA8zWyVLT
X0HfisiFPdEcyJ7iqZqmZtWgJf3upEXmxEQFXY1A8hgZnGwVpO+XkdiKAOXRiabYwZPrEHZwt5wh
9zS5LL/Et8Jj+7dLCsbuu/kQRUAZb/nuk0RSw14HogqUzio4y4nq4Y2g8FHYLeHacnR424sbfG97
bsEt5GA2UopGx8LCKgIPuGdNW9ZI0cWAQAN7R94Gs1pRg6tDpYz9pkNAurePNatKwvq5U3tWU12I
c3njsLggKz3FVQxGJUUv8YzCQ/LhfULxoIqbgFSDmWor+9xFYTznCUc0p3HDjLL1AKlPyvFjtmGL
00pJEZnYgigflkOZSwbsmz4QGZweALB8ESRYeR7IhxznJ4WJWNmOXSRb8T7GvNfQIUsC8eZ3vw0m
usORSLAjb01H3/MlG5pBVewBNYU/uEAR0bXzV5yM9j/LBAMV1s5hqfNZtAqlWzOlvPFzyvkn9ywA
SdQ3eVfO+2xw9zF5RzMNVspMPDQjAKS2JFp3rHEeQCfczOVJMSIoYoRI1lIf2fA46/U9rvF7pHcn
7OAlO/taKHGL1hH2MfxIm5qvKYpT5TlVOyUnGFRPz3GXL1HMvUZVe/WyJ61xXmIwYO5fAHgNTO6G
3lPVOtTHaqZIaQNYz623ORvUi5evrTJUxOfx8fPJuCbM0NNACeNsMKXElu7E3Q9gjWSHO9zTd8BL
4vUZou6WLyMm4JGm/Q/fiVHzXQl/A1Y3qOXCEHoe1jodDBwcxkbsWTS1QDQUX/RtV8LHZSjWHneZ
EvR5PyD5zjCGJOk2+ORtAds+FkDR04i/ydZfpt5NuXE8TgPQGp/gt0UIkDdIqiZFO2lW4Ivbqtzd
1GAppXqRYxCfkhFW7UaWjsnyVTCD0zHS9f9ukxCe62VH4p8ksJH4fqVeJ892+ET+u8ZJi5h+utd1
ic2Y8N7LQ88irgtlyD8ox5j5YQK+jMstk9a1HAk5Z/G4GM1q4eUW1DFGtBWUY6zooX69E0y/Nmew
5NW4QWXXue2+pqWDrXPqGcCXuh3eiUQoF3/IJ0ncMJOwi3UKgJnw3hosq/A9cL9Qg6EMPVYOX3ww
Z3hqZ0vNPVMPC37psipyJpS+lAZmB8+RDXPr3I8qhUTmCrSvhA6lw0AtfKKYL3y5bEmym2/G+Tlc
9smY6AEYMvY290fGdWg3RgVxa1LIf9KxWZ81dJXOhVHJ1WkmhJ4OS4gtVYT80vL3ljPbNLiy9m/Z
pmX1DGIwxctF2qF/H7m+9bDckLbE9XT7MH1Gqgx/DiAz1X8WCnK3KPaWm7WZtucnd1alXE4MoF3p
ACO9PsTrSO4Bo1haMoCoXoQ4TRZu2AJIuSej9E/WUNVm7tO/S8odxjzpb6T/gNVH61cHSYyg1bi3
LyyT7WMSEbNJm3fvdfYURqncDBLTKmBoyR31TGEG9IKCY669ZrLsv+barKOZlI2Lhg1ozakPfFrd
Zqn+wLekIwgZUieQNo4v1rno891ar2wUnzanLcRrmTtsmHWdEz9z3dINNDtL6RkuJaAr1ZzK1D6I
rWjdL1cae5BAe9dALxLwAB0CyIqJnF4SWRS1w++JCHKdBzHsUWnov2wh35oZ1lFyvL3ZpX5YqKdB
GPKN1MSdbwuvXzFfkXS8LbnsdA+CmKfyUGj18PapSDPLvVEhTXM5iT2DGbo4HTwVNMbuxX0J/Ojk
FDf8R8cVkALCj3UD2LLN5BJL9m2Lke7fnddPN/qhmFPwTbm3D20pTngy5gXxEZK+1bBEwXi/VVsB
U6MQ9rEiM6d74GKIgFWDwRfdGMxLZ2n/StwxVt2/9DcoeuXarLl8zimADskZUSAtvWRp44BCekdo
BqDTLjyaiZZtcZaDQBR9B6DfD8mm1w9oJSF2tMaxsNAapYoGFSCyeh0zq/Rk/KCX3PGKm9ZnlIht
6/RpO715BqK3QpFkvOyQIMAScyyISfEJuFiWpTjdO37IspcgsPDRiG6z26ZtIIwpUMAcvuLigZuR
/iT+fon0XkXBkjQn1ECQbC9149DoPTB8knR/EeetYtlcz5Y6E3aF7o2y+r6Lf6RXP4BURjZZwkaJ
jRUK3NFKRdkxOlP7NIbnN4D/gQbuUNU+5aFOjcRdthjO093e8AtmD1WH3LWMn4o1xMuxp2GUUJdd
gYoT0Q1fRJXMPMDCje3UJ1vpV/sehyzd/rBdIsYsAnerAgm7ILAK2Uh3EDjMuei4ZWANOmEQKVTF
yMrfpN7zUS05w1i0Hl7OE9Ur2HmM+KhcZnqkNQG+yi/HNBZmwF0IMwagv0pfJZA/kFcJWcUCcfcC
bzerW1Pa7i9MkG5mw6F3sxVaR0V6YDCzAMKPjHmu0KHL6aF+rD8H0Fcrdh7PNzb1RxGtV9d8Ok73
E4TYpXDIgZg+rhubRdk8zGnAQOs5HFzEtqOG6CYXTLMR7tz6WrBECiLa/OT1mSKWWdwfwP9zWTn9
lT6ytqUhvKTng/DwThJySOgtUnagW/391YDunxm+Z4qkrD2CfUtJsHAN7bFx82qFbERgXnYo+fdI
oZqnFal66+3J+Vl3TJ5Q6T+tZ8Ox8sHLa8j7Jg6TNEE2efiPab0K6VY8GXBKxl/XtJcGCTfpdreo
Cczztyjm6x9ZtWw9XDSAozcjVBLlh33bAuQ82CmNkV24dcu0b6NbNozP/GS53gKdz1dB3+Th1f1I
IYAqvULEj8k94rAImJEaKbb5Efr4yUUU3mDjecZlMpXV0Jx+ck4QXSqXBkdmo5GfwLboU4cZFxel
5/PCzakTcYxC5DmQf7ihKlNkzZY9oVp+03ow6U1fDYuvvuPZM/nOiTbvp3BlLMLDHJArzjK68pjq
Tp1xCipwGhTjKEQFw8OTuM3/lqJ2MsJNM4sQOel5U/ht847TXmbjf4kwBsIAyE83cHp1JPsrtW3e
8+4PnNhgkUq1pXmeXot/7T+JO9aMIVTDnHjM2QraobgGUD4n+zRxtaa4adj2nIq8nkg20XQqMljJ
tcQxj/EUdmcj+eRlviQFPS7Co6XXPH8Yds4UiNcpoCLVtE3E+IqgOnU0JKdCnoC4w7KYXPcuLaFu
nuyCk3k0q8GTLAWHdKl2g1YsqZdOr6kKQcGLjoMf2QK2fgQq/CjJ4LV4vgx8VGG2kBuo5eltQpq6
TsB8Qvs4qPv2HJjRb5BhIj2MEmMiPSZoWfvQ3i/4/DZIOiIKJMSy4AY+azDBE1hgwYyo+Cwr1iJP
+4kyoANOJLOjnFAUV4bXRwy/VLBM3buleh+BWKdT9Rj8LqORLh2djFVDD/g4yz/bEkLXnsag9k63
AHR8zNz/DcesLL0vqTIk2TKmf0dWeo5aQIpcRK/SBIhUSNWNMpiNFgcDLHMKBnZP0ACHBfzyBUv7
we97E6nruRGwxJKm6rfMhIEWItRtc3kqkOuFkD2N6IogJcelOfLAh1gCN0yFzLtorMTjC274cNZK
z2X31Ph3MIpXmmcVw6ghvxedIwCIbD3aM2Zxa9ZSIqCvxywWNPNwPvyZAmV5SIEI/gIygbBQOhcg
2MQhFLVKiiy2tkS18eI+W9fL0Adh8FJtg8PmcamHnUSRN8xRejoXhGXPvItRoLBaVNGE8p+mJbpH
81lnKCU1Tj2EI2PI5aLXef4jgF5ni2lkaIOBEPBsu6Nx4nhpKfHvpej2znKcLqdurEj586J47F/w
nCx79mM8jLkrrBErSjLClbRepY/yuOkNTZjWvECle9QBelhweWxqIm+8emLUxaqzV6R2vlntCHJX
PYfnc33SGx9DFdTWh5mQaD63RxGo+wVBaScvPhriaaQwowasSckpbVgAnLzdX5mGMQgO/CP0OdY4
OZeM1bgveCByWsfd9lOg6PSJ3ZmW3658hscNTpl8+nZnut/JS5AAtoxm+Nwgh6mx4IoOWrRLNSb5
cFa0KNTLyNHlSn2MNNkRHrML9OG9ANBagIJz9lueFV0fsjeUibv81b89Ua7BAgzJnIfe0Y6MNpqy
eHNZG0ystqPDnpqJRcy2tWjLJswQ41Iu92cG+OPafGJAk4WvFNC4Qc40AEEMcnj1t+tkKVv5BE4n
LSaRJg7EeNsI8VNPaej/EOdnczQF0UMKmu08WNPB351qolwvT6mbxTV5PLmVF8lKPZV+7Lc05nZ/
mTGFX1x2cV6sYOVOYIvZ0ByOndSDOj2uxaatLorMBWECWDb+ji3eKvem5amVrHDx7sTqURtZZpZ8
b7CAcNO+F6cUfsDbd3rkzDPzUfIWaMcgo4mLiBCn9heOE48bA7s0wFtLRS57l0NofYCf0ld5mxla
o1kKWiGvIIKrwu3AMnSX+EPJ/zyEyF8QM+7v7PcYEaI8f/lQPln+9wZNGMjYlQULX1yaxEdFr2qT
pN2XW11jJu1l7btdM37UNKexsElq6aguLM7+4F5p4ZtTSIHBCA2NJCKZJFLUljEjEv3fEpbyG9uy
0opJuHIdH1OXQjJfGAdDWgpek6QjtPAWZu5puTNIlp4iK8F81FZgx1/UK3cw4lq8XtSa/v2yMwRy
wupudIcc1EzUMZTYwHP9xlXTSclldTJDsf2dlQcRUDNzhyJQoBgmQLadb33FbnNGsBI3Xq/Vo0w7
c1E1AbbQXFCgXbrpGQXzaPc2bI9229XGCjbJYHAgOK4qkuwFzxC20iDc7DP1B5+hed7iaoTZU8Fy
GNMj7N35dWi2O7c+2xJTuz8HQtyvMvS1sr5UxTmzldaOm7HU3peL9qKvphRLQ/sm07WNUDdbid7X
f9/LoVXO508u0j0IwALsrb41N5mGt/s6QSzPjn+WwohSw/PizBj58NTX/q9/2Z4fg2QJvSl56hyH
32YdNy0roXKzFRLrMUXIm+/1CMmDDdMDs6Ykn96CbG/pGin0zrILX3Yn8hP+oAsKO8Exz5w74Bcp
rCpxLxufYNl6Z802iJqoHKt6xXZxg2NzzGm+knRzuFaF3wl+D9org1eX0kx51SySrYP/UN0JKgj2
4aNAXaaXKZIscfepVllyqpkggMDYH5HrktA9djRXkd96Auukj3fQHKDOpSf/LzS7nZnETJoCKHpZ
5RauIlJwzgj1MAuIa/DrNc5++QdhVDLqxacMK925LBEmjygh/i7LF9Rv/gmo9KilqIq6Sd0y2vbT
vsmGtqk/52OLjazZuxde4FUXfKAwKvW9jrPbEfznBiIIgPu1psMZNbB4kasacPbABBWEqPuKibhK
qYd/AGOJ9ZDlVTUZUeYlv6ZPJM7//KHZqpfML47uUi02A/Fx7J6vyq3CpPx9+A2BFnhdB7hbztiN
wCYM5sWQhxZdIyWgLXCZ3b5VyKBb6ic/BqdglHj38za8n0wqructPNHRkTu04R/fo/2LKICLSULd
sGSmF8E3Nom9jY8qB9zIOvaFtwQktHeO2YoxF/b76Y12bklwr70vpuqORQHvVsil2GKAlSoJu2kt
7nBzWhFkGQo4NYae5rr/XIDLPMeYLIXSEfLoIrvLlmCJ7wXL+IOZr09y/u/vUlegoThz4PwLE1bD
SPk0O6ZMY3osebtcleyuxef7BZHRx7GJ4+HHmnBUYp4FN25DQrIplPku6NeVZop5l4PSwO/p+0x8
zZhUhMgtTLt8bsPoIqDr8Hf6AmVf4cHnC+DLIzeL0xEqyHSv4XZT/1M/g/ko+NZ/8mYXneAfnGvj
EcZU3UWD/6wjI6kdeG4Cv6SxWwB9T0C7xd1YUi0slKF31raDI3C3CR9LVYc5IIJ/I324VrMXiTvb
+t2VbnyjYtgiNhTk5yubZnSMyxvpqK9tC9+sk+rCgE0ueeSEt0Vm68Nna078HWlM3bZ4BoOUBDUV
zfSKSNEh7iUHKr7B7rEmXptkvHTPBBbLG3WJFXY4jcPRdbo+LLsmaqSgaWfWARv9nFSSsDFe/Cbf
LdZT8RFegc9Y/fNQCQLooqh5xMNNKVnSHxW4SDK7RPjTYxpoyyQzRhEFs7otxIH54EwyYacvDTYj
uvrKaNJm0arw5HkKh8+RaQ7nAw7FIiqfKX4IskFeiWtByeftzSvqHkVZ0Q6wZIs32+mllxpjsYsI
DvBuWbHqese7ocFGYjncaBkJIXbnCa8ptKm0fSOAtZhJbSSaGsyjt+lYpCSIdGNdooOofeXKUEWL
i/rSxQpGxjhNtQ772tPEIRA4MwGXZq82yjgxAjW6JLv6IHbTAGsfSjOPDAGLKmB41NgBUeyFGjXN
fXrHjQC7D/c0nc1t7XY6hrMnCBO4CA++aMIYHkVpF7ob/UgPlnZj3o8iA6z/JvXfVzGFKs+2J1L9
4y3J/jYaF+nZVOKUJ2taSw2I4Gc9ulTFaN3GEpv1UmaCQFppAKZX9qjBRgyKIB+n17v5zpC6+iv/
Dvc5pZfrp8KqCj+U6cwVNEOABU4Lewqnp4mmieoqfXpXbkDSJ/ow4IaReBp0W8Y+o/elQkZj5FZU
1VQA7/OWQQkHlgTOP071erXIM3bM48cpQNIho9C18TeJNGur+knWWqWmxh9my/NcMEuqWMTbVS7/
oDjxx5jX9iAbBUcQQhMkeOnajkqO8Ft9MVYgA0OUv1pKxh7fQ9ySoG1feiW3aoQzm0O8PATsazx8
fwbq7ryVD4GRo9PxYg/vujNZf8rfa0ZDWdMW3BCjP5q4GZuI0rLPc36/6CgVbwB/iRM/A5vnF92y
23hu1DaDU4pH3QJ8ZaWRA8TkADBy3jEpQ994k6KoAVliIggrY3RdGFxOZ6ZogiLGWMFD5o5hU3ai
6W1mU4MeY5RpkaC5AvmBm5qbfCJ0Ky6T6WW/C0QzeapwZEdgdU/twMJ2ajTLyjgErlD/+Ny1frB4
NYkfpZRq9dROlHHRwQWCvaRWbxAxlB16gbHt9LykW4ADn6hKGmgvGYaMHff4vAlmX/3UaY3sle1f
gKAmq6uJyFiKSU5mBUGSKlPjq0njQJ1llHDymlwk7yzSPmPn/cjYzCNnTU9+yfr0xQf8Xpk2BiTk
yxI62mC2zQ5D0m7V0nMAb+yzpYS5JGgbdh1PQYT0XfMj0ypPRjCQ/5JbBUvLpGPlRGVYK8Ilmjsc
K75pRVUr8suF5uih5QH5s0x/2EIHKSusgnQoyPw3plOxI0M8oo72YC2HvHQsKB561Bivl4yW4l/X
dwqz9HzWldNh1KA4VE3mZGLD+fgUArzlSsXjP0H0orDrsUJ8poqBF7+cT5LUPd+rLKNxQBYSdDwQ
XKt7Kdajj20si/gw0y9eyUi/J6mHMLR6bNfB8zL9XmwbNtv7Ym4UYIl4g79lFD0yhj11SerFOftb
7sgoeCrM20JmSYrXz0S/dnbXHjaIweptGfnc+vSVGT2/keF7SLmdj7NJJ5Y1zapqDJ2Bg1JcgexE
5raLvXWZfu8jcPAdOmFWbWoNOrEg9rc0RGiYNGPmj/7Ba2fKsiNiYhP9JLvrQ4X2PvvdRHOEbvQd
oglXWhS/WcLCQVZ8uIKzklBxRmB9VjGHDYbOtIpbTdiQkmn/sDfQ6ql5nwYFFct4xP1XtW1y5DJb
Z6MLNKRHzNjPu/CoSZwUwxaDrWTwfhkC/RKdfH4beh+E1sfc3n7aJijBiKhpW74YXGyxnBnxczXj
AWzQ89wk7ZvTAR6MbxLp03FsIuDhmlo7mwfB6py/4lEZYoQPMOUcb5DI/EttE7Vg5CeHssjDiiv4
OPYjPS93QCcZ1h2GQdDzMBQjHxN3ZUBdZZvC8E0/AZ5ZWwSnta8vzHs2d6qrrVh4cCEbIo8DUUGY
mKQdk1W9eEd1ujgYUXXMsvy1MQK5ssHVDfOttlBr6jesF1HyuqXex4AaIFqItC2oiougWO9KJ42x
AljBse1JLR++wM8BCQ5gWpA3xPUz2pq7pjN9cU9G6zUS8ltzXuuEKQXZ17ZQj/IjD9n/qEdgsCSl
Wq78NYb7pLjj16BU21SLNjH1vd8xEIwpSZShLUgT+MNaRYY5H+uH8sgvdyHasCQBNvCsBjKj75IF
x8+cs2iDxSdvvJrykOEdJa98omfolQqNOEMAZtTh1jhlLdk4kLRbFyWvjrqEZi297Pb1z1yspxS9
xYzbdItd4zb0iOWwSthmJ9ZB5bc38V5TsqNjkKWeTEpT7rzctVTZftyn61oBvqx+vtBOSAPGcLsI
CcnJ4zV8eNkNiw/RIDWszDpKxsoSgw3kmKZQF8uxA3QLbbZzSLQzCBflzvkB9U41yPth4uWeEiKm
qjkKvSJajrf9bmAQGWDL7I7AckdNU5AHKqK/Ytv9gbXGucBDTKE6fyoXcIaThlkgmRbr+6/9SPgY
773qg1a+qY3Tm5usPKow2jWK4hVI+UWzx0i8swGtSAl70SM63RRPrPjzMgU26zU9b/FpIEusuQ6R
nqdkagNjN1FJ86UrLRIvMZIrqKDM7MZ3+9H0CZARPHqo82JAXxG2qGfqlBEnp8uNGSwCJfCLEgtS
TEAw2CSRi8MILr3qJkBPASXOcGthLDZzKrGnSJVYqbptRFfT4szYl0apM2axHPvztC61DLMzyXwM
npURJtxwuK9J8TYIIf5y9dnmqZzuUqkI1kpCUkezawpj55y4spcUU0dw7qC4hwpjgIWDS5HFYJoR
FE2lyu3fhx67ZkJxChiu4leBeNjNJhLlh62REC7kzjNECTOeqABnns1SjdFiY4WNK4R+SYMZxuj7
0bzIHKqBSGeKxHBDdK/SoQg6oYzgmKdHjNnxGKHOWpC+NuwpB6yWqBlwQh9WKMLbOQi6hQnEbEM/
qegis0Zszy+p8tEME0WKO3mBWNjTTQtoHYvlV/Zqqm0dI5xFMiVthn3/V7WKXYFJcBggpJIae8V2
4aaHxj+97PJDJCT5zPSs49BzfFivhLtJtORq5JBn5OHMCnMb9zreW24m0DYZTiwDksLvhB2wiZPb
4EI8V5gDAXExbpsjJnkrH9tUBm8yrc0gIM0kk0Ydqa+WW0f8r7w+S6JisW+DUK9hUI55uDRMfZw8
bl2KfhtrbMxbqkJOLbMs4Yy6nWZ+v4+CVH8OV22zUnW8aG0C2VRTxo5PftBUeSTBb6NmZiyVEKaU
1FN5UvAE6MnZNanmKrjev4WaRCEjfxN7SAOld2m01yczi/FAtZe8eahwcB53E/A3dRGlmIPhSfsV
/0vsJ0n1+p+8wYAe6rWFemSH699ZOwWq8ieWkSx3N2fJJ/Mt5WTZQPfQ86jGqIim5eVEYEmkPTi5
SnfC2a+lfdIX1AlgB1RRo781ZG4JlkvNM5LfKsR+XQR8tD02/Fv/VioZuVAkaE5XeGnmXBiB5x3/
z67zdoe5gAkI7cNn7MwzfYAv+V5PZVpFszPM4pGL8PB2YAploBa7/wuL5lVhO4nMRLVorG47AlGB
L3xD/vCwTfyRWbBkFYWkYfYBk9jJ+uj57bMuKmGF6xaUS1xFUTcba3km7kTbbKKdvgdalzomnZC+
ani9iaIxshIp2YrixXHzSnzg/Le8/1kijBkdKUPCF1D3/cQ2wSids8btlVMyjpE3vENGg2yCIBh+
pnJ5t3cLBvxU3NaTgufBsLvF8p5l5LbwnYUZac4CSK7dTrYcDvmrpWORvD+y415yL+e3dbdHXjXb
uLXOMl+DmW03bl6zzkoa/83GJKrEQWkmwgBOiR6Eoje/0Ygc7LR2I1k+tzhAJUgVJXYkhsBZCGI+
zzV3G8yXoVtmr+Z3XNzcixYb8C2m5MHTs+p1zma/Ke5Fj9nmKoyxVF+itRuSXIIRdBV4CfSUAL0R
HobgmuPVtbsgdyfLkg4UdzM2TgkHQGWUHogbf2Vsqn7xnaZGpE6v1yvpYPzlS4wbY6w0SSJYVPHz
NIQRHp+EEOAStMS4oJKAcrq9+mcrvtJLJDJ2ra5W5XaqL12Yv7oII8pTFcsLH/c9j1w6GHsp7ZpD
DWDRKkJJSIkhfhzn3Fy0BXGP8HYTeF6At8HlViklt/Thez3a5KYcUXlMaqOgR/yB4JuyWt2TuqCW
8zg7gh7TgSlBIdwhX7tDFaDbCuYb52s3gtHLYOlNLOyFMuGaxedOoPUdczUcdTO3gReGY5HfyKA5
0+ljVuFz2dKc5E1oW0BlaOAfoMPhXUPQ5SoJoLvF6bC5Qdcv2AO7TcrEn3IIkszQ6+C9ce51kG/x
Rvv8Ktsb0DMVmIEQCRTPPpgClsgF5O0W38zIM7Es/LOv1Zpfkoh6mWNeojnw96yXKNVIsPphJFuo
X2Sl7C+CO6tMjr5bbMKSxy+rmIyssyWhnFmfLTqe+D4Vq/l9dfZCAiiYOnIBgL6C/xb/8lH5c48f
hwYz3YJSF4Dcyy/KDF1qNQ0sMj0wT51iBehN96+51ZIybhcss9RMtgRgFgs1Ov4pm+1jNROBkM5J
6GReKC+3wC6OI8M2QjS0fQRKMOg/sdealbbaJocBknlceAw6le7CePjr0eDmWWVdsG+DClpFU8sT
hqXJINuH8IP/auYyUzPBAqNkUH4K1Z6iwVTS2KkIdwssBwp91zyJ2Xijc9Zq31MYyDxXiglQgA/F
Do45THHqXKzv8JSPtoCb89dzSGLCIBvToj8x4nCjFXpkZVED12KxQp3ppe1UU60s2UamqqUjuz/8
WIMxBMqdNY8FOxni2ldsZCLgVxwDLj2iNUV0suG/8tC4xFdDtRTaxF/lTFV2XtH98j0dtbb31Wuw
R15WfzcCNXz0C0mTI1c7Jy8mxy5Mdc6d8JpUW/uGuV9uZ85g/pC/WaWRRfaQHx5l2org8MxLOu3Y
NCW+T3DWesW4sAjSzvGJ4dwHu5JOtlJ4JI9jimo6NaU4BhrkHhDzZNj42Rv2AKrBrU/a76Mozz6V
gptKwLKHJNDMw4lkMuuBZ9OXLs3mimwepSkuz6zZE9G0uX7jlJvxDnw/7fdRNmT3qG6BkElLs/ao
/0ZTOOLhoMGUfveagfH0V83HW7VTQNobuhnAGoaG8HnRC8AzS3E6Qj29pHBwRLVBOcGGhd8SzD4k
w2s2T2c9Iqy+NarFSWyD0eqhS03X2q4gJTBuaLkmXhkb8UOlm8jyKHVTWAtvmJF4H6t/wlCSxo5w
a77MkCbyyhhYXMIq1MBkY6Olk5Ue1FaMn7VCko+0iDW2SU6BR4V0whTieSQMrbdS/VG451FPFCBW
ORWBg1MxPGh2Q7poq3NWuKGrF6NvQkTZNI6HWLciW1HkNmxTOkxPDxkQXrWHU+hV3Kv+Qxsp0guU
/bYEJVUrZ1k6zt3BODBH9ZMQb2pjneufzVrRW/Br1j1eG/zy1UF/2zM510vvEbtjkxcUgiDnlUP/
o+WmSVQE85uvNzNKyzyUkqDG/mg531Qr9UHAQc51huietT+15pbUb98BbQxdKFI5iKjByyuoCdfE
GYDKvihIaXppuun/ATu829G2/qfZoVg4gU/E2NifimvonuuXhvt+QlBQOel6XvFyHeEkeSfr/36x
/txmX9k8Fi/ioqkokyPRWo2SqCMZWGH9f/F8k9mdefDfnZh/m4ATnLlIl0Syu/0Tg86P/inoR8kU
8c+AHhefyBlU2TmTuiz115Iq2Z/1r+Y5qjAxBkb0aVkKz1lGBJOG48xNJZOYe1CIsYsx4e5q5XFW
KraaE+R6IG4liyIITmvjFiQcJaWHpIhctbXcoCIrMV1HqzbqK31vt/97mcCyfed6/uvZW9yVzmm1
AXIPeRz02E1aoGnq7OCicBE28KSAReJ7htZFQHdVSgW+R/C8rcZ7spBJep/L9FVYkS8jgHuqYkxM
UHvA5dmGOB10cg+fcrzPrr2Mx7oxyhzHdPLRqUjqx/Gx8JJgd+0C8aWqNres7533uMUZxPGZzKqf
9bwf6E4NhCpfFgzsqCUjDlrOzgpa7NuJ3rsfYrHO8DckfoFX/tIcd8pPIHENS++1lD//6IWM9yFV
zYnjPivpBA1LxFkM3PrLAyvM3FxHAYb7s4aic9OUpuvNhzTSugB8h+o05v0SF2FWYCqf4rAZsBlv
9vnea3iQEaQGsGH1ThHFGex0cS8i3RvSpcEQVXStu774XCOGf6opf4QJogU/6u278fl9Kb0AHPPi
qBcV6/g/rgB4zGIDHyOONVorvyykiCgK8+D1dIr6Rwg4a3QK7WRzVnznayGGF2cjg0Xri5hPSJeq
sgaNvIyQrOiOiVu4Oc103zKmXk0+sjCLnyYQAkl6ycjnS3zI6i+AHny8tT6WSXKm16NZA/BuWXYo
WshxGrtsQqAh4f6/fISt38y7/FFRnIJVcUZ9/04mHk6Jx/DP5Zp8zx/WAm4senE7GY1R4zvUJOx9
OlYwP5X8giP7OfAjGN7+jGIAztl+YbF97Enm6DRp+fKlTs4fyuWp7/nywfB6chWhMhV6SUGwyiTF
cJ0LqBM7wYe+94/tx5vwGjbwlvKOPY6/AWcmvg4cviu/L1yMbxLA4LHqtkdtdP6CKcusvakIl7xA
0HnanE1iIu9/vEljlZNFbx+sr4cjZWI0WSnCPKI6dkg1yh+IMXDDTxFbU7ujig6oCizd5DiJuw6Y
hUqFYY6rvQaUFy1+zotDiHWqzP4j2JuWRCgWUQlSVqmvvgMjpqTyw91l/qfQwDHl+plt3O96RlPH
HA6cd5z5ZA/hxE5fqPakrJ0j5LSK/t1qN62X1OIA4N4dIX6UqghhBKtywvRf6HpkKxCepLTRNYM0
f0mH1b41HK8rKF+pYuP0vGAZ0WJXkJwS/DuKGhT+QZyvHlnaMsukC4fpJ46fwtNqemIjZgpByLO+
ueOCl5tCyBpCO67mnAac6V/egn1bx2zlqN25XuQwEIAguW/b/EfbXY71uCmo5+ARlCEfUysIiV0y
/SO83Y+zwDBbExolfhJuL1yJ9JRDbJeU08nl/irbGpq/T86Dq110RwbNItWr/Y+NqD2j4kenjE/A
0/dRc4R4NlP3Xjpytxv7Tfq9YaxsmzfZcOf2VpaGxy5ycfKhi3xHB8uDnUUoXBIq95dUlGLuawra
7KZZ+f6jeQ8onTpk5SwhIXUMhTdYHM9lOoY/xRHiwmdYIG9LFS87jTidPtVBJRuwNJnjYUTzmiPO
v4qBmpbj2l44Ehdy/SP3MAdhINnb7HNYdYYgm1ZBsS3w3DBKobcw7+oLaIohojod9TyI8xOIEp6X
3IL0OCbKFVRuTW6NC6m+/udCrRT6osK0jd42zwRN5SsTpGohUkq/bluBQBfJjgqqOyNoXy/WC7t4
uZotUEhnSwkqXXpQwkKW/QABKd2cjnaZtA4dycq/npbKngpANu2YJMxc3Ie9nY430Yi90GYG6pqp
LRrgugGaH19wU8g3/fXzybFvxVilMe2P669EEQdLn1eVWOd0gvqlSHn4LIagI/vxXiyrqyxCM/Om
MqvB5RhnmYpJ1i0CWEocEbFJjds0FEjSz1112eeLg1pMofchVFHj/mx7Ndm0ZHlbA7u9wH3R0s4t
68F+2zjmksmQus+2dysUS6h/6KtQU8bXF8EV1dA2KTv2aU46oO2CgXRQrkJygYBYR/TN+sGRkUEQ
DL1AGE9K0rl6iFHmSIhlhHFWLXo4LSmvX3UC2O5oAk/mcCT5Cr/M2Pmb1D55crYTm6oaRYCUQ4b7
D4Hx6LKq/4pK5kuEg5vEcP1f18saQC3jdZKSdTaK1Y96O4nQSBl1JusaosGOSFHrGpztauF+3Qy3
CFglU8oqKQ/SAHr0NB07P1la607qvmD6CHkyhW0ofSpzi02xepTZ6jHgpxq/c/UjnswjHkL8EsP+
BgV+U7ub6MYbs9cdZD3skmXUxpyzn/CNpR3Ggzti3waspa7JomYvh0sKdD2/wMAtY1eoA7OeW4jR
MXyLP5l3//cec12UppoqyDkaAl+dc+mFPypu6LBslAFihaMIly4y3ViO4Bz9MT/r8mGTUOVHpRFW
LsHM0GGY8vtG9BkjjF44GvS4rPVOH45o+wsAuD8LN0zbW3wfO4zbUTF/bVf2ZEgFH9EBgZxd8p5s
1EbrV5cWsF9UYHMchQ3EGa6q79O+cHapArnULDB8waTqq4l3jzSb2cLddO+4vuMrh/S4vALA4qYz
o1AlmZpeTf0v506duEKvdQA9nt5SrqC4SAN6OvwhNmF8UGZeg2WCIgst18rp7B/BgP6F8VzHTOn/
UfLIrNLCVyDbcCgLUNnW8TRg0p22++0IuH43VZkF1gnIneA1Gtree2OsMxdJkWHMHFMhhAxWIAWv
dqKboCc7/B2Z+yxm883eMlO75lb3ByyeVX+eJlm6x3gFvjjtnzeftA3Hr4grY/3tVv1zTPlLgHgd
j5yahjuYurJJdFLS1nkM08jpd7gWWtBCPiRqzcAhnxCMyN7JDG/nYuaMzolugNi6NIzg6jeixpsl
UdhGAyeFsqyEWxSM3cxydA87N+h6a9K8kpvuGu+jma87n6QxrAfDkaU7Mo3mmYuO4Z6l6kLyRcbz
je6Tgnzli8NHTv0XMC9Wn6aWRhPwyLE2EcMSKSDy3dYQ4quih9rxolf+IfLnBzZ+wRit9wDJThgA
K2B0da9MMyhw6H0SySVqpPl+LwlqT3yeMYfhL2Y1dRkuGZVLmxlCDn7wSeOy+ntJKrJ5lQxYn5Id
+j7EeHUfjUjMHXqrqRb5UN7vByyREP10Cbyo1rWQtDKJsQlLiZ3spWqxk78JHhHLKwR/lj3wQVTS
u8QcPSn8vX/MWJP6RRuDPTd4QGrsRQlv2uv+LmBPUc6RiJmCfavyBK5jEU+ZX8eeIZUyZVFPpdom
Mmclck2pm16jtCjrZtOkq/1VHH/reOASq51y3CujcScnstGQoEykhUO2gdiWG4kglN40Fkhhuky/
B2JrarBHU08tftLfJ36vxp6Y1kIvclk7GXsx2Ap+qkEAInTWJd102rZxmrj8Fc1GeF5343Dge5AB
sp1zsn2wUC+QBxCWfaPs9vPMuxi+N5Grfi/ETq36+ulpbbL5bOtiQLl7vPu2AuNAfsX+qWthY20+
KpaX9YTs4tWZ0ymEpgVhwSqLPefyzoWEFr0d4o5qtc2hSAu6ukoQPKysoShmzIbV+x4Ie2KcwnO6
Mu1QKrFd097r9sNPITB/7NjJnEASwOdcIILcJTKfn5AuM29d72id0CYcZEbPxjcmK6kNu6LM/oNt
cZPbViMtnnVAqbBZTx+zzZMRukMa5iAuLzKmt4e6gx5wilhrfFbxMlxdUYcPiMjntDOXt6N5HBLA
rvqBNddXaDOhO1cRkSLTsR0C4B2PGVyYoQyHvVGAOYek0LqOIl59VKhzZUalW0ICA4o/nOsStVZt
o9Dgo2vx5fBI2xXMQjNeX2+HnFE8aHRhvs6Eeefh1Mvu1JQsJesObv9vgTprkZ6ezYsqBzlDzV6z
afUvTniEcYSo/RpNA7Ujjq/1rXUFxVO6otbKFeiQAa496O0/0r8VFkFIb9bKGlvkkYa4koPuQq7T
/jl/HYW+hbZH7WKF3/33W6O7xbLtBgzKZCKZK64HixLvuzRYnXUliidosGpNQGy/h5T4HCxkIcBe
Cb/kIjPzxBncxOytCM6MrM7ZByYNLbW1Pz5BnBqEHoWpd81HOAFNI+n9uMt7biOoraZ5RPgIqNxf
vWKOPVr+JEsCx2CjnvC4tgbrzhI8hBVlKRgbi4Q2RTcKdc0NS9WW7xn/v2euUFLStCAdhRa8V+oz
XzH9s50WX6yZc23LA7db7gXYi7kSzMrnWqAAMJk1GNMjYSHxf7GEDky91mD1xvKnzChlMQsvcpto
39P52oOMBTPqyVtyxLr4ZG14IgGxLfl86urO45YgKuzBTROgNzpayPWJKLCyQxVlNCqlRteYCRBO
MRY9M0z2VvQbXbC7FiJq7ILa35hW9VpfDYqrTU9Dvhm3q3/+8kvEhKKmcpp5RTjiyTqwikx7heTo
OWy/SuezE7fduAhyOHgH72R1/61f4vn/Qa0A+guOTnHrhT7UvLzA1/kGIH/QgTBWg+Sk7T0Jv1ZU
apnBe6dsJU4Rf3Hg/Za0KTSF48KpAULA9iqvjmO9OmICcBwK6l/ljIV7dqMAWprl+6UBVXdzp4UP
zNoQTJY/KngUzrJevruuFgrELjabOlwfZfSGKZfjfbaHZOZZsI+X76qvuFVAipXcOYrMbVBoxmv1
gchFwqezQjr61+d5M7hwOUfetBrZRnQZ5Pn0Ry77znq9LambXQPYtsGxXlA6gkwrPVJ1hZ6SzQkL
7jVQslmdUpfI0WUviVhKXHiLA7ENRaZs3OBeWgcRHGomyCekZ+jpaw/sZgnhP3SXjV4rbIq9ZXfa
fRjbmfkoBLPKXd18JR4OqAtWfn0vCF2y0BKowN6yhDXudIrRNbj9Q1NVk1TZwraek/XOMirujS8+
yjMXyJFMi4Jt/qj4Mdh2dBWTfatz0c4NXABNMAFAx7UcbtDlYNj529GzemK+3Pt84uyN6IN9Ixcq
FKeKxQsiMqLXT/DoVCcaZbRw4hsWKarEFNG+uTS7VEeX3EepYP3gGZI3K9m9CuteMSUMS8lBomGM
W3e64DFlStSGItjN5Hl/JhMAvbhTQAvJGevRU6DXkhWtcFJiWb9WJb9AiXT9pStCx0fnnCV9EAi4
Mhdx+08WlejWUYZOKZ6W/sAefJUMn3FK6zpKPc9jvymBB7dL5jCG32hSf1dl3MFxVmc0peKSc6nA
o69xRjLT7K7wyQwkGVXOphBdT8/zUIdr+4N9oN7HjaeFbqXRGGoMWAeFIFKrsO/vuy+zgjSI9aVT
9KSqDyQX6Y+rNouFM0U29+aX9VCrZOXOX3+hLF8lwEtHI93Q2/vftJEnBncxJj0Q+eudeuoXeX39
qLGc/tBzohRGbnuJFZrQJzDnHLmDjROJIJO9n+C7RJ/bR9keATV8CeNYRrRhgrLi1HacUdJ6Oti2
duT1N+4gDsgpB5w+D0+eCUFi8hfiL9QapCO5503KUsDd5dmExuhwfvPUFnn/oiob4Uz3soQ3YkII
gVgJ2kUgvbH/YrFGyyT4S/jZDF9BuRg1xbADnm15T2G5w0wGCZW+s6CjdXIVaq1E+7rZECu3I9s/
XnVuMIrUPOn+SfTjkFX9q3VIlH7sqdRzKsjbnSqghk8y1GahH61JIItmOxJjsxnAEtc5DS6PwRdo
6K0JLRFDQJs77CfV3nSMDPYYuYow5mHvVfJ2AV5xhjAWweyqIXuRGzUv1tw04J4pHw8juoOKgpfA
59pYe3UdryRqjenqiYOMzWvcgI92ZA4w7R9k2okHBqTYbyZmy2qsxduDuy2vHQ021RE9ZjyHqzhj
4TZ6g/a1PhSWD0671Tm726l6sUJ9femdIfT+mJxW3sKCWEOZKmPdUiYIv8v52+o8ZGlFSMDSUNlr
USIGLzRaVNqrcwnNZM90VEiHbuDCxrAP7dAdDIClx7KUyIocO+Uy2OGa4fK0Tm3d6PPj2ufnwsE0
KhtaRRLWXO9998bTOVss5ei/U5lC9H34bJaeY8O9S0IgxSA8m3Ew3vlrcv/XqYvWOen8P6juXGIi
Cyf4z5wzLf6PcSzkFVsCqcdMfQ8KqemRXbd0V/RQdyvRDbrMiAe9DFz9+YFnwtH4XkU6FBjPknAU
J7cgs62zeLQdceFKC6G+xSCLwphsUwzbr0gkxxnh+ipiQzwNzYJQEUALum9xo2fvVNu4h7x8YheS
Xz6atvCdHaq7YBioBpx6PLhyV1PKXcDxnEMFtPGe1MXirrJFnBRhLayFcHedLj1x8PIPPfqusbDN
v6pKViaGUCcORZiOoU/RAAryEQnXjVnrGdLEHPomLH/sANWTaV8XcUf8IBqgrCccMi7RBf3KJudq
+lB+Og/8a21faBJ/fF7i7r6Cf38krg3oq8vekNw09GORy6dekS4jSYd2jceied5sgYdWWzvznJuQ
9yHM8X7F9x5IAG+CcIiIG/7VX9Zcju28ArOatya4sE7mC+lkeOO5lKdg/klqTnxYrr3O31SrtpE8
YYIpuOwR6UBiQX0sBSHjCtgpYogFds9PJiLoX48odS/7IhcXRUUtY9jYa3WGtuGVa5TFWdX112fS
kLjBgiwTrW/Dcw2K85EZ4HyJiTjZOdpMM428Wv4XNv5Cq4N1yd9zRmDi9ZAAuOTrUGkTYas8r0Hy
Oz8O5NfjxmBo1AHFoOiy/7zcVn/hr2uu0wmOACkIEP2GAZJXmXfFxgCgvACim8dJK5U+R+JFw+8K
KYVy8rrC0YtuxAxNs1C+/0gxsmxCIU82YARzKZL6naJHeCGKT9plnDoTWrMDTeIVDA+T1Q+78B2S
ZIK0YLzI+F+KAVKPRQPl6du1sYNZBLX8e9AV+2Dkb73lYGmZdj+8fPL7BkFDLnvHLl5+AOo+HGtt
kKZbQAXpyBko9TBIt9LwtDWRlPZTg63YzQJ3PYCm7yLfiTjBydRwjxcHi6cVyrOQTyTE8HMI0DVV
FlIiphPq5AgPzvp9ipj4d9RY9jXiTnirJa5pS/N9c3rKDPeoH3hsrPZoMtnsrg+/3xMblIuS5qHT
cjMsq4UGYxh7HWU/wrzLXfJONEQTQipMoT0buAM8zAm1KSx5QHanQgGHa87L8KleLYU6+qJg1ZWP
rViXc8enOKIzfET0sVOyF4pNgmQa+XuZ01DvO+kAwzbeza6kwwAsMKQl+mzBx4+zZ/HmGEW3D6Bq
+LekUGxTuf1YC1lJH+3Cpvym0f746+KV9qY+ealj4tNwowyt+mYnVwECdLE/b8Y1OB2GW3iXJs+E
fOiCkItj42eWumxieUgcCCrsHh+HQebY6iXKvCA8DdU0BZudMW888vPuMMBTcjxG7WguHnqkQczO
n7/Fuk/mi4TK7LAZ51h+TuGQl1sdYl4z8TNehiYT5Woqr35SrSn0KZ97sFstK/8TiVX/4lJ6Yb2/
HM0VMaxa4aDIYNK9Bk1Pt2HAkCAG3w7XUaVUpc4abBDq9Q3LTcOhrUDgLRTKYCSY54sJ4j2U1u9N
yxFT7Zp0aBMh/CVvr5Q8bVZBstJJoOdCdSLQgkPOoB/NUXy/HlAnMJTis6h0NzlWXaDxPoDIdfhP
2EhS/DX/Y2DlvJOD3W7oHYzhETgHsd/g3+FMXQCjfnShdPEq37qpt3s9Po12ZQjz7u0L3d/2Rjlw
cgbTYzIJdNQXSZHp2PYWCb0xhSCaJ+97TwZ90E9CuIQ7c8RBVYVd1RXEkoNluXx626+gV7msyoKH
8RNJhwUbQqQjTDfNP9ceySArCQmGN8C1nuznJGliB9OePrSqouRoXKn6W9eVSHKLZoIjsj6FvOAi
/Ael4+EbdiDIeZnSH73/igYNGRf/Bu+HmF/00E1u9hPLnXpCntJO8bacCAwGh+GNEc+iDvZfX2w1
8d82M+Cxbbgw/hKGjsPy0vczuL38iMBa3nRm233jfhBLClNqRRnpetUDSoI77dlJFPO738SzU6fV
+zoChcudedwYJSXJhnizOVo0Jyjjekwud3FmrTE1l7cJDDDzuuFE7gPdt62/qO2N9U0+wIkbAmyu
1/4gAdZR/kVsLF4afTEUpuqI0hz70odud12R51RR9I3AEhnD5dacA336umxQ0dnLi8matWyalbyl
kaybWrDvCuNb2cWBq1TZQwmr3k9ptQLFZtWTyVJ5nHwmL5EJC2oIwYkK9O1wMigJgiUb4uH3hHKY
PiMAPShngRymBkhTl8DdTLdUUB6niK6J/CM9DSrc1C5YU5UAhHv9s0wD1vK5A/NxZ8asjm64vcLh
REg1paSfzAwTqD8Yfs1TCEGs1WjCqgbLlWKBV/2k/SlmknECrpXnWa40Imx2u4uEo7x1rT4v8ndO
r0JtvU2A2kR6w3mSuF8tcRsFLPTZq3FOYvc+1hrFT27bip/0/ouMS12J3q/fzc9DRPGi//W98tOU
VzOa/FMC2W2793W8rOkcjpQUu+Uv/iNYTZkVoVKJdEZ2NSXZno5wbAAG6wNW2GgnGoweSMIxmeyp
ne0K2OBxv1TsBKreu7RQgD8bPG9V7OI3UeyLbXhO3nrVd0c+1+TcaGmMfD92M6dSnssdd7zMdWjs
lN4w6+JsjyGSjnT6LqcAfXdoO40GoaJy2FDfhszvrn7sdpNphpZUWzUZgo3c3y9ZW7Y2eXnZZcoq
8RuqynxHbeSyuKoeYHAhJKH7jCZ3Q8lbzGy8XI9LQtK5wphVDfPV3GIBKULgyTX3+nr/VIwKi5sq
eIj/+idXyZ10AMgj6a0vyM+hBnD8LJibWNFgSGIbn3264uIVAamLGDLhfKB8W4LnwGYESHdwaajP
N+Z0UO+a8Zdce5soFnpSq68B4kx5d3QFHCcTDkeqTku7y2rFpQ3KnLvx5rh0WpayayQlX0AkfeH9
BAADLYS9o1c6JVPM/JMGgniPX+olMKB1cm5eLe+yDMDXHy5axN500nx99ISkZxTCKtaeiiBaLLKS
noG4/8u3vLR2IjrhmXFJ4YMhMHB/pI1t3CThp/+eO4WHgx+cadS0Y87S+Q39gazrAVKO0iVjvujL
aj9EnJzGMrKDggJjxMse8WkbFJnzuktZdaO0yNol06yzoEPkwuugBOs3GD9jL4eoLb2jpRmuHjtx
t/noKwkr7+keT6vD2jsIC1Q/vFGIiu/t0pLWldNtu0MnoUIIVOYSo6cGqTTUux/QPumPvH6zMMRJ
4tTQNOVcruKdY9FEcF3xP1DRo1tmnJkPk6bfEpWTI20Em1r+QiYE3OXLmNTZ+Fxg945AX6rrZbep
wnh/XXcT4YZaCmjYHiOLnGfNvr2cK1DB+KsbnX/mafDdRlAt+9nHSQBUZLijPyz2KevCtUQsTBiY
rN4NCzzWtMjBNQGwICtqRrm4H9zQc9kfWae9Qx2WcF8hW/rmBGXgU7fBB3LPiAiIG50dIO5nG0vb
/QygFIT0fr0E28kPOQQAHEVWK7QRx2HfJDICJxBs1h+y/Zjcb5o89p9NllTPgvx0E2Se5B7WIvU8
lQV5kgtaGs9ONDuJk3ZFtQ4+SZl4GYanPOf1ZnRzUbeDTPY1TKZxPUE+BOKzdlt5NZ3sqmjvtLSl
/VMC4kxTzhZFqwvhGtHTtYDzqNo0TKkFWYfuGPXLBQRFwjXWBqoGEXklks0CudrOGAqkxqDOsZTC
IU0E4P92zaW3gfkzy/wqD6Ww2OCiu/TWxQ8r2LildhHaCgKzTNkyxnZLH+IcvTAwF6B2coRLVJaH
TZsPZw8ko7xtAEiQfgPo5pclprrQfxDMbJ0ROGf3OpVu3ThSKB74wlCHutMAG5QrgEIW/FHjfUSg
2/kCjdZ78sDJi4RHpQvw9/ZTYacrqZjjTDOEXCoKZ6cd1MnXtJ41DfKqga/TLtSBpWRdlfffCa4H
zribgyZlOxxCzMVO1/iQ8jpmb9KTGCa80ThZnx80X5yDVuVXMDLvUdVTNFdfgkdoExJYSdhywBv6
3bia9SvXfYhKCrB6Yg5obG28RUupE1pPGGXNiWP8F4kriPcLBmmIYtRcKPVnLjJIHa4dEckTkjZI
3ubbVIv+UtQlcdFsXyWfv26u3ULNMkerSLC390/C9MxtdB5hR6IHaeskgCBJafv+6aL9rMVCOGX8
s70xyHrVHZ5QYMRe1e/3XiyHtZcq9s5e8Jy2oKjOdd3MaSuLaqbHCn3T2nWmiNjQm6RCVGEY1Tlt
JGdWUo6W1SlRGbAVwumSJUEl+kuRgSJC3+pQbpyu/jd1QMO6aBTyDhkEDfMrT+HGgXvn2aDlBd4m
MRBz8svczK4KPhrt9wuUC+P7PO8IQQO8Lizco0mUHXrTI17YKVtVxI4FXhKXBGbfJmlP0HEJJbiE
vbGDmu0YWSJIP6nY/Hu6LlB4UqAXbZaAIzikPksWuzbXaEAhFp6d+Sy1RTBNQYe8/TQDsp/Eriig
3Aa+DOQF1lhevQM+vPrqsOjVJ2QYh6if6M/KOWSVyBJahvj0UOCVb0SRMc/tY36cupIB/6aAjiBm
W5vtrl4wJreQlgfWQdqJ7acxAcLG6s7tNZE6srQWFUZcjExwPBu0q06p4n3Yf6+KBR+9HGTCe2tR
i6K29AApYWlv+4aLAIgu/MFEfeBzhVfrBN5/BqG8jYAB8uJAbWpg6vApPx8XSC3cCv/fVHMThXcQ
I1/+GdVoaus58LWNUi2DRZf+aUfEV42FU4EKrBNCi/MmvI8BXEWhG8fGOh+IWe/j9GH4Uck9JlmE
q9y8FHG2p5BtLG2l6GcGyJiT8m/QwBfkzI279L+74RqAlwKQoSV+2rBOEpMpBGGXdZ26Y69Nbzol
WGhfw20RnORCTymbJEcZIYaCujwuX0yvu9QK7SuSaRZnHkZcYRpT9udTNzqDCT9XlgDhK9UxZhFA
JcBEUJR4wvV21VKh7Irn8zqEzUDrJe+3jrwKzXoEuVjwt/jbxnh6X3fVAo4RhxLG46QfUDzt2ZR9
UL82yrv8D9YdMpAoMvQ7WxxvFlBCDJEWS3nBQdFnt/ugoQsjg68Mo5gYOq8f8Gbkvio2+mHOHH0Z
o3hKq0/3pFTmnSqb1tRqiGMBhNjL4FOXktre34BQS//v3eyf4xJFwPZa/fWd9w3TG/4JL1FXt5kM
g0gkdO6NNGMVLNkXft5zgEaPq51trX4yeIcxixJl/IKPVugLuy4VLLMbEyYM56pcSm937W+CxGZx
vpHzTYzW2pD7tY9zTeoLq8W4bb9NjgBvWHa+NKnlmxp8a6O15Ble72NvXYbZ5DPuCXGcWWBG5tl6
ZRgMdAxnBaCl0xv5p6fF07QwZhyynLKCkZxBJ/E5qAWcc4HXM1s00Mg7AIK7kZNtsXn530xuJUXG
3yujO9FcoXJrQKjeUz/hgVaP+ukkDGWauvu5hkjMyWtjZC9IDJ2V4qBKk/G4b9/JKgIMHiJW0as1
OW6XjdcHoUHL6TlkUcAPZdvNJsIi0/MjGll0eM2Pa0USzajG09VhMYjsu7CnxGW6BVdLNqo1zUMl
NnXmbPYCpKq9UeBC3o1Oq/fhwTkA6rcZRzejE5JxY360tUs4kt8lTzmYr6rUV9IsKgDSr7QOMB0U
XYbzBe0NblM81pYTtV2m6HR3co0UhIybY7qI3s6JaGtbJBzzdyd+Nwmbdo4/HmLeaEb13XrpEIWb
C27lU0g39h5ys9RB4qawYMQ987hvmvRa+IyU4PfyYD5Mia6TqZNv4yM+cudIN2IMEkDSOLMgD9NQ
fICU0PfQwKeG9pcbsJm1QRs/Q99tHM2gqx66bLsD7NNeRqmPYtBOv86zRD/OBJi7VrG1o4/Lc38J
8YQhkJ5AZOoi4T4PTvwoOfJLMNlQJrFCQGVcmwZcx1TSary1PgxliLnC6zCjNpnPITqp7fAdsf8y
hsep9nJrFy6JTDNWSZYtxM32I5K3GtCMRaH03/S8CzlndnsupChKrG2YRChu2/RsL07glblGeVKk
ld31LBCRGYz5yuURczoZA0tuKtnE/EjVKku7qbkCWjea1JN3FhURTwe4/uSNngeIrf9T3Gi/x+OL
O4wkM3Fr8u680cXr0FutumB2TEsUTMYs7Rb6ggsOVB4/bS5g0kN1TIuCK7LmdfFGxE8jdzT29rk8
sPlpKPkMU8LsgIdO8+CmCPuDptmLxPczdFyvkshEjY+ug5pIT7augvPyA0/oJCvJme+Xg77Kns4A
4dZp+vWXpc+g3dhlEUqt65zbtMXBwKxr1zdg3DcUVsYjaKIdRXwzS7rtV9DX9AX9fvtclk6703nk
RnSBv+pnC/WVEXpo67Evd43/bBFN9A91KpYwN/1o/oWb9sbggMw+Tx8NzwG1jaEafqSP0RtIsB0V
c8GJlZH5ZGBBKJ4faYpY3LYUKdjGSb+a6Ne08uQh9B7Id+9jOhILImbyMLy58a/UDdm+3t+mwhNH
XXRsTR37eKd6AXVv4BQuzPGETEUZPnli9xXVma4AUcW4mCLUJXUrn4l3p93YeoYoHtDwKrM/kH5P
MxNPtySyvAB506HZ6BZPfgttGNaXepa5MPAgjZieEhrYhYhUaHnUbco1iE/XsdxRcY9ObT7i9pFb
VCSl+yPfslK/WNsZM/2Aa5k4Snw8NN8Cos6KCBnv4w6IF3ymoUWe8KlzyPcYSlcv1IlXupDeV4cE
8/fFlhmdXgx/agfXg7/J4Wgl8weG/PLIohCy7JgeONg+M7BTTphWVaeWgiIozW3MRpbzKxXzWic0
Hbk6nkF6DQvGubOduH+yu9+/BY35jYIZHKDK5pTHnw31oPalCh9w5OoX1jo0RBM3hewVPiTjGzAE
/XmrdythGwk2FVOoNjEGihFEfALQjhrWfyMAf9p4HWkyfo/a+tEz7awha4H9+MMOSOKBa1oD8Pq9
C/Jax+brlrqvmOVSiw8Kj6t4tINQlbQ/EJaupFp83cznjuECATr8SQluqEc9cIO21QZecySmEVyD
L+4x/o6M5P3bDX3EfbAVfgIlp3bThPzlB/bfOirRFja1rDrvw2e+WhYu17fSZX/kDZpdoo6hWDxi
ticrC/YPKjhjeDMpXoXtwLGlfR1yu/bfTTr9co73AzG0BnYXB6fHCY1rVLuJPxFQxx6dYZtxMlZG
LmyqPnXkJTCIVRzXZwyfng36ce+o8hcTGtXLk7O1gC8dO/LSc+dZR+XFe0xzMgHMiklIgRImNzVs
8D0JEqa1zOmXclIybT1yZwWIN9CNvpBxyzqK0pevGPmvQIL+1N95qRmTOMlctNWzN+/29ZfSmbJk
p+nk4rb26/iGnhRXjorMheupAlUDJ4GnUwizpMT5I9wO/v+R/DxttvYLke5WjthsqzfHw2hTBWpS
ytV5eJbam3Ho0IMSgplgLlYslFXvlVcVlpz1+XGCh9w7hZXrVfuqhm5GSgDxUVQbp7UXDrOPv11q
j3oqlcWsJ6wgFjbnpYoFZN/w+jveZ3zBmN6rkbHsUOjAfa2HUe6Yb21w0531LooHrfbUCMW8x+58
AdI09sRpXlrLyKiPgqc2XeNq1xhwwp6fh7Bmco+iOhRkIqMXn2PP+MQMgB1AzkCi2Wz6MhdRjKvm
v/floYD3g8Nd7I5B7BRuSIEO1fOUspyFNxB3L4b1up14WzqVVlDbV4eeHPZyD5WARKbgIVHZcW43
uUCOhYsO+srY/VhlwZ8CwqZ12roNwUKjESxzYcbbdO3xaIbn/OBsrcytMBpVgpIcmt8xyoHg2Dmw
LBEQ1AgzO4dsODckJerJogsi40z6Cp7bNmig+BqXSP5TQ26PBKjlOX0O56aRik9/j3bjcfQWM7Rv
MLHODv+9ljp7lenZbcnh+REKmCNUwx4Hv4VvYI3WPXIZ6k1M8bzIIfsRSI6Iub4p7L7OiMH000s9
FOAp9g+bCdxgOK3UDZUxbRZVpZZmpiNul72OodrBUqhtz9p2OEUxlyhEp/6ROZugYM8/O0G9S4Hg
cpNHFnIOLQpjTdIkH7BKiiXNI0OipXZxdfO9ogGzEIkAVmzkMAaouoZgFsPc1+fyz9izMGHPvWHX
u8J9svvlUgxfyJYPUS7cIbVZDvzAcc5J3sv2jpciSWttLY5QSI/H7I0VvWIG5jCEPQajs9vm/NgW
DP/aEeOtJcyuv0vMC8VhebiYmwO22EL9Qun6xaK+MJ4jBk1pOCeb4CrVk9lCuLC5VWjE7DE6eSMy
i4lca3cAMeZ0aNjBz1G6WXQvulFahld9uDwCCISNOQ85FOuq/i5uWcbbnrqzTEHZgPHcidmU4PtL
24oT/AKMLmq/1Dgr6ZIAmHWVfT+Bh3KSfVVk9p9iFnEpslj6tJhRQCmldwUER+PUe4X5BiRHOqZj
90DHk6I7vSyYuzShULN6sMv79oGaAoWEIXiDieP8k0pSGp2qC6mUl+dmkA0jH6Gqd8gP01GlVGWc
wa+D14mY+dF+bzkcrK7vrUzi0bEgFYujvnOpwcXfMMHhQKKx3vr9D2vWA4m1MzwFxOd1qfDfaddD
Ksv88mRByd8TYJbmDv0INyyfws8p6r+jv/g3kg7zuuGRiDBb835OHFKNfoGJWOo+9wcSjjbMRlvQ
vwQNLfnsZUYj4N1P/CxtI/QO/xi1LvHAPdjdqF2BEGQYETI1fb9FpCU0pwu7fcq5Nz5xO/W6ZNwX
pHcUpBsndfJ2f65Izhrkj9Zd6NaYw6GjKd9VdxQwkiTkjGQ7+eCdA67i19c9k0og1hCiyxX5hCi1
AgEMjCSyG/zusNYX9oD95elfc4O00DYmaE88w7g/MTGJjtpoQ2PWjVrWoDwbYCW9JS91/OXvfzmD
Wtg3+H2sr8uArJi2yZ6yx7jnbXVW9CUcaYvXErK0z6wcoGpleWnqfOarDskUdM8w5tbyWYu1thu1
IdqK5oYEWLHf2ZIYu65JPRAy3+mbDyvsU18o+GAWpNxqzULCCIM+51B7lQQ00RUmYOrZtB1Jj0Sc
xoXXFtzm0jvjJib86SH7o4YoQrtshpOjSfJJQADG1bjiKkcwTWq6nfM0ghLi2KSAjDz0HynOhKx2
ftx9pYbj39go6FMO7Yi738lgGAZMWE9iB4No5nw6GspjOaIky6zkRfvWiimY1EbifZ43dPV5dlwK
exQoBSg6EXJfUHrTsF4H7mHNr96o3yu2lMj3GvNURQA2kOPkCIURBp3btRLikETIwhBbPvbOOucE
WEtP2xOPZvueF6Xb+k5CkQVJ3N5jHbI/R1M2joYauggArBXaMAedfU68tOx3IgrHGGhqjdjIcmNz
IFnZH9VBlXPLwlDdvaWLmI1iZrRPqAQq0jy0BFpigiMFF/edvwP2rq8Z62y9F9zcq/+y/grJIcgG
Is0a7UMfDKXRAuZEugUskGKu3X845/RygxBjx0ipPO+ZHs6IorXqRKZ8ceeIMJmm0ITy7sWfjQqD
N8jWhTxwsyxSrTK8XZYdaZTVZ7vuCSwBN5UXuKK/g/+LWTFFrxDEdXj0QbYv00X7gyZz8tjR2iMv
04cTiH9M81lh6MnqxPnehOE8u4CCrt/kK+C0VQ0sRoG+1D5jyM7UnFlr1vf4h8gLErCoFoafIjrM
+lbWBY98+mOrDRs/tUnanI03gAJrxZONmV7603pU/L88swMUvtBv/qsI8ybRxjml0HC1Idel8C11
cfcz39uk9TRilt4QhiTAm6ioa8I26JpX8lrS9w78seXcTzLjtmBxYlD5jeVDVULvwlXfthLhAr7h
Kj5DTL2lPz0/6nQ2rQl+kUsOgwS9+ZPIGJXqOVyiR5Pee+PmZQyZkkw/LTiQgfXQvf3NEvaE3Q0o
X264wKbsk6okMVCYeyvTu/hOxeDkZRxbnw8uiq/ffemkuFIq0i3FEkgptlfd1B7xFh9H4W8QihSM
3Cs/+hTFSM1sRHmV1RQEWv75ZJnm2qQVdudYF3p9rvVAjoA2vzYax5CfiXguZ4kxc4ImCwzJGEsT
10gcNSkhc/9LJoslQj/oTDvl9eIrqTKyJpie8yYj20wFDNHiLglFr3Jjc10mx2N0vQK5jjc/P+B6
gCYNw6uklDXGJvy3mbz846AEfKgcvCUtXKdX9CeBu5zaJe9P2AwpMhdGrLISqvje9W+EjO/lf6YZ
XV4XSorxGjYgvxAJv1b/gzdFiMmaJtu15Gt/osHBu4bOoyu1kY+E53NLazYy4Zv1SCm95iZTKvIw
OfsqBLZQoINrkRQv+7BBr+C/2xLPi/TL0iVMEWvKoAoymn5iu19KQyMQpKumyeM3u3VBIebVI6qV
mpKT+Rnt9IV75ayrvDX5zv82Xd7wqB79q8IanZI+fVUt0L+FuCUS4tDZaGAVKf1aCk3plIdVWHLN
4akY2b0hRpqfBOAkZ5oyR29CkaLhzLrhPk9+CKp1ltDulIKkyKb/7ohNsEmYs3KDTpkioxQUBNnR
SCs54IcRsPT1UsafQCGOzujkfjef2PM6ItTJQZs45yWa22DSPPaJHg19h2FJ+9eRFwEHwgN7auIS
rQRmQ7bKevq/pVRcycHekFQpNdjIclWVYUZcwaFjpTXaxEOre2CaDzWitYuRwM0aUc42763Jc8wv
yrp6GZYBzbVetA63PeFUaz2PwQz/8f2dM/jaHjJi948CvhMC0snoneNpVhj50w0MWDTUP50ZLysY
VRtqSP+TMV854W9cgoSxfdeZd8lRIA9BoNVs3dRiQGD4XKGVBjgJLwyO/Jx0qVZK271iw4bhmkMK
VNZEUEzqwUq01vP60VpwcXQS4OD8D5gWjX1xBJSHgQS5WjQGLgC/5HkTBWjlOTu+Yf8CzYUhn3fV
WpCVxpqroYHmokzZ2SUlPa6Bp6qKtVnc4UozL9yQTj1BwuFQQOt6GGuQtMX1ItGB/mgB/wj7ZK+K
Xs1Wnn6LQWpkVBIbrn6ELo4wp0bTl+EJON2h9e4QCl1ETf+JW06gztVv491AbD/2hEQDDJMP73NN
llKwUeiBAPGUlGb3OPZvvmra+v9xB7lWYfAYePXHUyUdMGeC6tP5U3APdRPotIp8MK5g/e5DC1IB
qkXgz5Pw9Qc0x4BqDGgO74heUCsDxY6uHRYq/o19oHWagSIOP1QVg+860JQG9cCarsYHYw8olUhj
Xc/rowW+qCkF1qQNJPMOCm9GUvHvYEaKr7YsnObvDqBc+Rco/CBnHRLW69hf1IYh0A8W1W81D5n+
9jqgzUTZjnbnR8QP1e77AFdhRXMNA6WjUBJDN6t2AHPDMJZ8bNhuN96M6UhOjQWqAX4tlxc2A7pT
HQXXbJZUuGv7xQPVgEd0e2wUG4xbqgTFk1SvZYSVeowca7AMJDjwsUkdcn2yQ0JLfT1lV+HIgGCe
gsA2aAQH8Eyj5WvcKnppShBCZTxTUbB2nBwhg5ERIUzx5vwLSzQhtPol+Rf4hrrwktQe9y8rxPbe
J4y8EfT2yuXeSqy1IGrxkjMc0NRhAjW9FJhQXbQhH4cvNFZIc1hSE9g6Ds58NJJ6VRErVe89cNvg
6409FaP9dp93Zxwej6+47pIFAQiPSv+XNJASGpX9lghFANVm48T2PnOaL7d2criLD2ksyh/AX+r0
/4VBJX04wdiHnO9tqlLDb6oh8N5YXeAcAPZAkkaxvOnyO4pV15iccVPwIMdzSZ/u9IXS+T9gCOIT
E9LFUoUrtZRcyCOcymT9rbq5+2SXY/59DpJxxGKJenP34tNewM27Fo8/+d1+r4V2xLUcX3WE1Muz
p+0bKiiguIzJD3ERAvPWTXxVmTGshDwqZ15qj0ziRzPUFpLSzZ60DzqAUXmUg6+i0RZC6eRFaf1O
vYtDeLvFlovVxSNpQzPQ7Lg6cY/DUarlF5Ows4bH2nLTLtmKkGMisg8HZGIP8flLdPSVmwv08jhU
m7UTA+5iw1bJB0oT5wOLXPbxQKJTCGCrIvgMCUtCyWrytlmffDNmeWcdrpnfnkpTtyyvMjmv4jXU
KzQetHpHHwnP6mwq8a3XX4ZswUxM6tYy9oDylPWup5LDjNJRZNGzcQVvqOTTKHktFLtQDDh0SCJS
FKeMIsTLHlae3R/5dtuZ5soB2rd0eWKh+W9vfMGnVrYjid1G6X7333ZdXNsUobabqFp35DxAKFZM
oC9a3Q+uQ6e/mjE5Y9Ac9QavcvtrH9SVrvZ/AMvE7s6oBVKVikJgn6Uzr0D4xUeRjMNUn3YfRoa9
jGFjrENvx2m4HMqT6pq9MCdByoRt0+dzLHRWTgpcQ8qq/i+hLTjKSwBmcZkUSW6PKa8A7mhEe781
SD7fFUJKr7HnXcKpvxddXxXCJs5p32N5aHecQ8o2hAQW8sOEilYOaQE3zbVkVrHNSEM/S8qX1r5B
GriK4JCmPqdIPK8xIPoWc8rheAJifB2F927vrf2GDpaGrC6/p4nwwnd3opMP7PHgO3lTSLYUX23H
3qIxGMEpFvbd93v66uyrG9VNJRtPsv7N/8vi9tQFmL/8Sr4NjNNwETF4seaNOczTY7lxzgdXiR7l
JaJ6uFHhzw0yRDszOMX8hYOZfQ5T37pATKP9x5P9CfiEO9pT0h30+OQRPYbGurMJhkm5uHYZJC31
oR0fgZmRPnItIcVAtHx/27Eowhloo81oye0SoMwLrzu0hL+4+uneD9q/BE3xRHv1ubK3hFk2C40T
0F6mKA9tzgGVWM4U5cW6TudF9Hd9Z29xqY56N2PM+4gAX8sKcp+Sx+s7usR5o9/XcdZXFGNW3pB0
ieI/ydhEJ7HbvuPw5y/SN8FlGia2lZY2+h29ZYDf5qDYR98rIHGzwNUKqvSIz7TIQO9NI256tJ3q
MX1oWDdo/E/HCsPCkIeCcc2OuAk0qPE5OaiEey/dRIbXztY87UCSNnMLoRjr9qfexlRcHO8Mvy4f
kmVjcHpGaWA8RTP8eeqDFDAhZIZcBJA4yszbh3StwKJYWNJiqLm9Rl/mx2z57F0MJH6CnpuHSaPF
VbmBN6tY+fmRUQXERkl1CYK5CLKaNydVNPCRb2w4G5e9d6ZuN7xu44TUpoiOQ39EkEgJwidrdDtR
8aMlbbchI1iaOGZOYmrNcv+g6m79tGlWcZ4cyBc+oVVByHhJBzQDb5zSw0MVJrXEeyC2Rm39ujyh
vkXioSsDhc2sOMh53hpETpoPuOqbaglLQ4tEwj7EqxBB1VIfiV3hv8IkhzHzQz1+GwcTz0RPullW
1t7nuE7IDUnZzEcdR4t0AIDMQbvJrimXLLO48/nChPCJLgQPxb+gYdNA/K4z9IfMH/WJtng1vxPH
xAMq/iZH9lAnAA3rclqzuRXZnVGGGuPdQAYZp62zh8qS2pxKzY2nV5mU6zjT/0tXlwhhVNSjxp1Z
H8u25ijzb198QDqXD7yPSFCyK/PR0qngW/C0QNz3xLrgfnYLHsbpHmgo5Q7+9otxQdPPjIsy/94D
dZHFKg/DZERfQFdQ4fPGa2EoaIQKazPNTnWsS81HL/clcbtY40zNEsqXLmPbsMQWnITy6hVLVVdN
XiQ7YPno8PRliFUWXrmYGt8uMvzqAX/2qIzyrhv0awBeghvkVyoZOi6eVZWqcA5LeKkCN63WmoUy
dix+VkH0amB9arQHBRd7z7tPo2M5tVH0ObtheDt7ZmMds9a8qqItySAuvTz+fAEXGHNeI4KFWlVV
5ZDh2gz6iy4MIBft7jA2tKP9RpRV+qATZgX5eas9LUdhA4+3YYgd4aRRRJ9isj8H6iUXNrKx8u1Z
aGI8XefMz5QpMJuS6ptQ4c6azJ8ImhWRNGwNUe6hkHjgRfUhkEQsy6/3Vu8KQl2UppSb3Phoy+em
HTz39spEfL7tKXfQdP6TNYzZO0tHpCsuntVhzObApCsedAnJgsp1dWc7Xe9+i4AnoGf2G7+mqEdT
m+jEyV1G21/6iA8OQkbuV8cfMNbzhaKIr0CL9UMR8tm1AFdp89Wu6lHEmO2YbwKmHiSpzDiA6zyF
tI1v502lYvQj++dbHFc7IWJSLXEl3L/cNSYWidCsUAQN7tA1UZYo2p+0wcPp945iG9JW8hpfERrD
MsCr0iXUVqiMpyPsFr+/oXQGLWCVgeBQMvGQx26zQt1htG2FaKxvRZLJg6vT+OeiDDXkG8DacGaH
C62HACdUJO5aTKe93G5FDtfd4WMVteYxl+jCk0skS1M62hvVKVh2qN7XWvpQivC/5jCcAuv5aJLh
eP8J5dptJrwfwXv64Dgw1DDRHoGZ2pOVY/YhteFkIRrNAuY1pqlTGScEPTi5b9d+DE3nYwcBS8dJ
wUxxmdB29FpmDU6EGkNXbT8kvJsr8vw5yUa+T5EFRLe+gg6Ur05DxmDJ46tZunabUKwUYrDFkMAk
x61/B2vvxSwWmsSmvx2yRyx7CVRCyBVW/zkdPijKdW1rb0UYIILxMIdl7fWaGy+06+Zy8T+59jfj
Lw4Mf1G5TqZlLxawI2s5msHBIxlU5e9fTO+ovqdeStForBViyto9wsk2cfNtdNfh+D/fAbiRdsCl
TO8Xqa697MuEj/O3lWE08pRLDFK62/QQTmuqvJa1vUncDhB8LW4RTo0di7S7cGzgnUAzLQck2YEy
KmuIADjZe7KBhUifftTUpHXGer2amd0pByGnbrsELcm+CsaB0gr/FIGRRvkmcwE/nlJZEcYc9Eyr
YVxxSLIvtJX2p5D82uGJnFHU5xjASAY5qvSV+L3bcQB4qkTmX5Ya60ghUQVRsolrpnZB/YfQLUMU
p6/H/rcwM1wruSQSZqJ4xcFaDH8MWhnXVstL2j04EwfCM2NIH2fHrSeTF/WeOizLZMKre4YGtFqr
X2yPwFfEOPr95tsOYUIVUjKg6DswFnZgOZrVE6/c1gL5Ogc+cDIt6qb8CxEn0Va6Jb4hkgkDHM+U
UPLCIOfgZm0mpBnOPq1OyTaDFo2khRcX/q0XEY6FXH4rMLIvi+Oqyo4wRtbvhfLZ8Tmd4PJ6LST+
BiOmcBOE0M6imPdX0LRjPa8mFDRWqmuExHfXaco4UAPczESC6TFaJnH4I+zDQ4YSHPYgv4gm6PMm
BGMZ7XIrC47CqLQOmkCcpIcnrqgmjAebv7eecPDYwid0JJBSj7gOrIT7E7NWNmKP95GVpOa3oGUL
dwGO1joeg7n7CEIzi9ixfFisVYqe8EtRZC+ASFh90bde2en/ZoXm905CDQON/WqlFROf2wHwwz78
2V6gyosrRzgJQ5VQmySbqAUmbo7ge95eebUEJQl8Nln8l7QIsDGet/r1wzH46+Qd+NmaAYlLlMoN
S3sNLi/L9N0s3dj5CzGTQw4N/+EQMWHywCYjJyUDknyMAKdVdTKW2PiD4PY905+zBmVdB6M7G64h
+62vSM+o006RAXPFaRxK2xTi8Hfet+QTrLs+E7aPrrhi4SmhP3Dv0s16jO6PlKKuao9OwmM1kpyw
YIJiaXbf/vHMphHc6gOOBuFAlVs5CfaHnSd2FPBlr9JcZUUaT+hgsjUaFvtwxNInwC62C9poYV82
94HiKYog8rDMewQst5C/IH8LVmKd/J4gy3kjj+E7DM+kkC55CkLaFRpTc/Q4+OI65S8LVafaojRI
5TTppjD/3LvZqgHx3igLr+JHSXTCCZcXjDmebqClHaMPxsCqbJmzrR8cKXHuplpdeRDf3kCMwwiM
SMzpu8pAL7Eu343vpzUqCJn7MWZAQgL2lF2bI4p/XhuN6kA7+Ibe8BhPcCGTAs0eDWQi3KEtdoF6
XQNp+4orWhQDO5iurrMxAzaRq/AZE6uMQLg6gUyU/IyHPZZ5DgBzu7EvhTOhk577yz1pbfTH4T9S
7yVw5yfzuLdkY9g6XEUoLVqhIW3HjDyZh0uMIZssbJcxP3n6xalpV5AFp5c9D9yFYpA4o4SjHeJM
ofmHuGUQlgZ0n9cA2WyRDbM17c561mP4YN9FHweHfQIMevq3Duck+Msaum4Ip5rN6o/EqxWiSuEy
lfHQbQ/Tjijs9Y0y2scNQ4Mh874+ormLU/muwmqN9CdcPxTyA8V6bL0hxsmktbvFeJkCtx5P1e5j
G/AyiyKBB5CpdnEHoNawrdWxnj4f/vWWspoTxHRUnzGyrSjbGlVv4TxwW184gWbh+xxGRoAIMiok
vvqkI7mJJp57txGVSreYhEU2gRHwtZ1Z7r860BMsl2XONexIicfcyPkjJUt0ytH0IJbJMCjregAM
NEDBiP1A5Mv7qiF1kPLeumhTxsRwotSGRaJN4riX6Lbz7FbBs+XfVpnEHfkKfUh0yBsl0oA0Fnv8
xW/JJf+y5nkwnmt62xq9eYkr8N04rcrNK0zFNQmaQdy/SS6wry5RPvREvJFmp+r+hOKtTzg1bEft
Ro4V84M8Q1iSQcJOJeBVbHpD6S8ooqh/1qkx9xd7w4K13BrQ2HJQi9zUuW1YfeH2cMmYjsRbeAMh
wi76daAMECKIvA6pQq/0fvKfMoT8ge5f5aqI3g4+RU+Ukj/tfaQgp7xvjrUIX/heFRQyhMwQBTg2
9MQA0WIfkcpu6j6Zn74eJf2b5zhiIMpa2oixk58EbLq0LW1gvZGsWeQAlmywFzPXpEBOxvunMjqj
7cP+AEPXkvUa+iR9HKJIC7FSE0IKG+Z//HgZ8w6azFBKQEy2FR2J1VEcSxQu/NRMSVn5l+5wt2Q/
j/okP3/ZT73ri4vAtz2IxVtRY1ChhFWirzJSfLWGDUxSdbbW6fyC+cXunTi6KsESblrg/U0/WFOt
BnBtMMEeKFVk6ScSNGo0hd1L5MX5ktG5XA/7FE7kWLcSZgdDGg9HCaROLOEucfmEmFqx4b7KRPdj
Tt5VVlxxJh2qYoQP8YxA28PttukmW36Ap5zJChbKdVA3SYprH+yna83Rcg6Gs/kTTbE6Kl/rQckO
7jhgsKfL/q0ft1IRn88lD5YJLwrtPXRNsNcqfu/6oG5tFhMonENqd1bARVn83peWu3z/yYYQpbfL
/nfr9IgVyr1QR4msphjQ6tVEomoOnrWpKKTxPlmNShxpLnMPAYbMgu+6LqMoOPvhHmMeUUI2dvlL
37E2E9ZYk7BrTrNsH5wfZt1kpsxKXJtiRhU8GrrUFGhF/rCQG2OLEfRh7HXwbvgbL9phRhIsFQMo
eZqFkxYENgjBcM6e7LJCbS4Q2Dl1Oh7uyVyocwnQHHw0xi7ylR/suVfrlyecSmSfFmAMyPktbnEC
RCzao3aijx+i0xzVnWrEISiU3uUJX5NkzaVSwadLsx8iWlwWZQcrrb2sIVaoTAg0y7u4jHxhA+5V
AJTT1VJlULWelCuhJwyT0YdgoCTmLAS/++5/5Ovr4twxB6eWFG67QlHsg1t74B+WYXF7FrJF4zfr
6Tjpnr5OJkNe875NI/Qae6dsZypoiy6yXN4S7moFvm1b+r19/GWnjSkfoJ6L2UJPdqY/ZGngVbg3
aXZ5Z7kyPwjwnODdNseJJszjtJPEO83RFQOGb8PyC39zM6/KSzgAXSfBWCYn5puworGV0dDSjnjR
Emn2nJtF7GZh6ju+//MItoJqgi/3yNxTVg3LdNB59prhZF3Q83qMMriAE9vqgvJBMQTxaGYSODCz
LjQ5hrxh2Z0z/ECFsobQDnZwydp4MIpvjUpT97y4hNKExoHvf/6iTQxPk+OTkJWRcQXamn9pLe3s
vqtaVK1xlaiXZJPsukyn7MmEIODCoR9FAS2+dbJU7b1jZ41YZTHnC851vzSVNtnxMZ9GtH5KHMQZ
9ZnbzG6mtouVO/lZbVg3TvBxeTzcZ1kTVB5c9OOVredcDo77oX/NJZWWy5ZPmj9D/S65AzABBdsS
rOCddpZP8P82c3NUD+J65JqLlXCRGmsUFsCQS9581MqGZqyzkALyGTWwrdm+YNBdTAuUqfNRrm4Z
2TKvH5E04TRRoMiNO8ppTqxAgzBgT5JNwTGg2OoXjkZ9NS6fAHKys/vJnOUtGezAHM7tnh7Sfuq5
0V5bfwbFEWapUtUSvFTcGM3BTawVxdORBf7g+0MsUHKx0WpYZFCqjwYjYbwcmcwIDoKjQZOFs5mT
pZMFp97V56RanimBlULjx7EQe5h6WkHELdfDcz3VUdephVPIhssmsP+dxRLtDTU3j8nkYAav7gsv
C7fgWjXOdveFMw4MsTgHcb1XMDlWuV0+lp50dD0Ynl0Q5d8RV4uOcTvPs2XLTQJlo/uIb7iqBPRP
DIJUfXd6Uz1RfV6OitbS9ZIrasEjWAdgYjrUcuBrLc85jjm2IYQWFb4blvskT/Ih0jCFzSTkVOxR
FgXotwCElrRbYpn8SvYn4Qkn7i35KibJ9XwpKMatnvFD5xhQAwAqXULEUi6fG5cP65IztVtIPNs7
XYCwQKMTCINlmd6MW55Q25Di/U/o7iV41iz3jsR27SPi0l7zxLXSoWk5ijs4QHxmVBtVLCNSS2Be
FqI0Tx/iHFpLIXgsrMuN6HWvgnwID5ziIllC+06XGyi4QEsDQfz5Wi/hahui3YDI8DjJ4iwMbGKJ
vrdgVbEHh17qUtqaX5SqmmR97EN8UKerBhicmtSbDDStrAVbMMQYDVo3bNjSEDsSXa8B6y+xveOK
vxzMiTxlYjopm+uuOaFo5zkVlZft/MZjbZetz8jK8a63/RhUkXN1tsdX73cz3MIRu55nfPfrMOl5
lmdy3cX8jIYREh0Eagm2ecIMqFO2SnjVYt6mGeYL6y/AOHwa+bqZpwMwGRdHi21yuv9RRye2l5vY
5CjWd5MLVFFYRtsEv5z2KP34VLgXDnhqHsEabfTs4rs8IMAhtn71RQDw1Jj5h5ECxHVujGVtmr3C
xN9aQKxbbxoMXzoloeMYvASXGxu9HBt50EcPY0rbSxN/HB7nX7JJA0Mkn4jIX543Z6rVXY/jRVvY
QctCiVi1SNfcVY5FAz+i+D+GZwPVsdIsPNiZUePGCc0HwT+4Gfi1v/180ui5Ag3VjHnRsrlHTH/Z
UvSO2yI1/djZd/AX4EXkAB1QgOsO2wdGjbb/5a23CL+5RKs0Vae/jv5jp8+34w2BY75l71hSeF4k
mStMtU8HFUsoQhaY4IiJ7oTGHBUY39EBOcq65cLH2f9XpNToKmcWJmKNlrHZ/hTu49KtMH4kVUX8
9GqBw1boEUi/Au+ss827VC8jcBDGD1gbK3Jyf4H4+r7bL8o1x9ZajRN4pk+qU7qWYOWRWAGa5/mY
JAFab5JajBibdX6kap3qOvYmb7FmrdYj4XFKy7aKNBO+h1GxVXSH3EZm/CoM8z34cibnj3okAsMd
rjlAYHOLx2szLUqPqVRk7bIDIE3djD2SQZj7cg6xGIwIxd/ducEvOCQdWPvUWAp4AZv53EOYgeM2
PmiZFi+eLtmGMqrjCmqYKty0qmDxQ14dQvPP7xmX8VDmVjTjcE8OaXP4+4PR9JgeX4WFCSGJqsbq
FZz0smXYU4IdC3QO0j/sYUSQ4FUkmK9XXZbv5vSDdyX4TFXh++1GcsV26H1jxDOg2hvN6JA0qTLa
eXEscpnRNJMJf2Zy8GMQs7EoF+FxfrpVMZQh1LhBVn79Gkh4Rqubc9QH3vTNcGVcXTaNdax+aSBj
jdSWc0Mkjr+p632UmCvUt3Gtcw2itsjK2jfJdTkBk7OFsKnqsdpj+q3kXFjqkjRIGCHiU0YUQiV1
iP8UU/cieiOHQbM5TXKbbB9sJrMpvfTuotVt7+mfpUxltFrFHTWPBHDe+KHcf09N3ziKtJkGqXkK
Yhu7GuVlP581SqnXuistiyv2bLeuaEtGBuOP3q3a9oTOTbPWtjPOswo9XdoDq5vNMC8e+/UKiLg9
gvqezhdlw+GCu7js2Lpnyhz76bFwx1wv9/zI3CDdyNJw1dMXSOVfCuIeQDhl6RRoQLk9rJtpwV7J
C12LxGVt8Iz+mBrTSRNMHquzu8GgXzOkUTLWQMISdLFMMWjEa/+/MEzWvD8tXo7a09B8SZhRaIri
KhXwIdYLlzYmAqlwFAuCDW+kbexYqAe+Tg5d1bBIxIa9/JJdO/rIY2kA3fobP5cZfQUTNHfW+7Tb
e7UBdGgWmvlj3yPco4Gzm2vuF4wNmboY+BepUDtmZMu8pMvzswsUF9eyg+gG26bcGGKIzojnItIS
KRIEZ2WKDOx0C9HbEmQMU4CYC84PPv4zl2auvU+JN7HAZFgAKet/K/DO/oHvhgiufIevelUIsc//
06CHt5dRF403go7HmKJhS4vZjO1pPus0j+ffXPR+9uqEXo0pKMKmM4GyXOJNpBFa0I3dHV91JT26
Mww3aeNJYVXqIlDEzQDPyddYqTl3aGRG62uZnzAr45ZNJmK1CtdAiAZca42GBkpkTlH/hf7DquhS
7FsN5UVqFtkEwmGe13PrrG7Et816L+cBb/eCe0v+6zgLHctNAh+0pNzfCWo8Vv8GUcgYBatSgB8/
z/alqM2aD2Hkti343OvoIZ29tZdVlTTmYxPr3L4OBJ/xVSrodmSkNqe3jKmF2/S8Z7fkF9zxAjRS
thWYiqYPJyRWK/uSaGZKZ6z9jjhjyepSptHa4tmKWHsGodjtrjGj9QOv6jGzbpdTaZauPSGy18ck
ogw56kFdwUXpc2WLShavoK/7ymfKecCyccRQTgPytpt6I97LBKeEZdcKz17yRAqFE+cVPFFGCk6Y
nE3b79RwsMMKtVkfpMi0sBKm6vcd7i6Nz8X9ByepFqXieneG44QR1zPz4ebXmaNJ6TBoCsMUukbT
PwjegUYp0UV6KenzBMf6iOyzMO60/oAMlgI+i69EZSv6iKU2gOJ+0iwQ0S4n02EtrIW7pndI3eTq
hl1uqr1HweTLvnk+GlZpLdhiTK7iZblm8ZwmPSLtLHSkPTy9A/8L0DKgx8zMvFewqrekcAnRtYg6
k91FYLoJb+C1zaQ40rkQJLaHfZgQ3sZ65oByfqi/R08X8LgLpIQ29W36qmahV3A188Za66TnUryJ
86vBqWI07x8yuzFUDS+W/8hqm5IFjtEZu/0+JplzHDxG6Hk1/bBY1VFEOMQOoRdd550EACPuSRht
QpLXrVZc3rH2tLDG1dSbtnKDuOwtoNWB4vZ+P1v5wjnKX3uNDY7vYnAnEDUD+StjRfGtbHcgylod
X9BGV5YEKZykru9/QkWROREUjZ67I4qM/GdDUvEQhDVbkCwHRiX4dE26auTDqCIliYma9k0bvJn4
PhSR2Kbd7oGa1j6PWlXYPALy8KKFcp9S6Ua50LZn/qw36vwywznxkvjxQJMfGmCRl70fsVGMjrD/
NyxbMvRwEuLMFL0EcgZB2W1LFkdXoXJU4QXs7N0H7w5AQs6TsuKvJKSDzTc0tS2Tl7eqjTZR5RQI
UOIooDBArwsDT6SOoquAS9C+c0SbqEL3L22jNGKn/8hoDtTZnRo5yvBfLrklUY+hPHnYckRoNbt9
Igu2gUbJFEkesLZG6IVFp4GEXBZU0NhpsZkuuPbk7RZtyXyYarMuFvF0NYirEb9p445I2WYAqXJk
zr8n7KP6cwC4m46LPY5Ayh1Y8/co9OlxjOBQb/zfHrCbAxYS4KVTuOnMXZm/J/Pb6ktY0dHNnG0o
y6f3Bxi16T4E7D41qk65jOeKFlHkQM2nfjwIWnUVkwVgOxNqOl2w9kqX8v5pD7OSb1pvFWqdyUaV
f+EbV89I+8ep9yrmPLVaeNKiuoqOm6RIYNW2s55MLSx2e2/zrmAzctKOWh0ER5dCpYFqFzkKpIxM
Xicimg57O0CtkkMZmV9xMse1nIspCLgBVVU6KYPDkaqtaHnXzNiF7Q3C2l+mahy/Bb4bhLwcrpNr
faBoe7sdI6pVHcLKtzaitBDGmPBkAIR/j+VSxc5QeNTfv829zlgSbx5sKlh30KyVWCumA7i0tiJ8
clwQBL+UK2J6qIR2o+iTqGo5qLq109dyvHyS6cUh9hH0AuYYjz1ImJoSSPj/NhGvxoACUt+0Xvmu
DEfupWMnijXjW/4GcwsHn58zKREy9KbNUKsE/2kITNXyLCIpmnm9v37qjjNM0rDLjPrWwGffeZCr
lILMRW6oDXNZFetvzOhDsipmFTb95qhtnqRt7eLsalWkr7OFIc9J8/gePD62vtjCEzMWCu2hpvGh
iv4uKYasPqicA1BkCi8YP4JMNTRE6o0ieq+2BVhhrCszHfRDJ4ptMeoIt13mLSx2CZ+dwsySel7W
zmkHKO9XOeoapvuvoeJWmL5EpeKfdlWroRyuYF4czPmYzykx8PJ01Qpr5ppCrl7k3Do6n7GxKWO0
YrYVTATBZJmfBiPWmgbdQmqm0Qng5m387OUjdOkBN13aQsxS/5SHi0gxLS8ncsBaolVHRDMkAma3
1UQ1z408pjfGtzWfE0Bne5nhNRMCBLBIlWmV3YKIRuve25dYL8eNiP9BfI4S/gdoSftO1FKVma5I
ffRjEhHMan7SO6G8dzNdC3Ia0bcX+xdkt2Hr0OuVFlsaR5xKm4I9H4669qg9CL2LZHFB2xYFAMb/
dNA5V1aIRCDc+x/FpdNeF++aWcTwnxOO/7P2RR/wt0lRaOpG/QIq/P1Nr1/YGclaWRm9+WJPEi0Z
QZV/nV+bffe/+d1fm44oTfBAJe3htlU7oAafZKKgSGI6jsoZ+85y4t9ABQWoHBDIHKLf9k80SkkS
ocPgKCrBSbT/wBSPrcS1D3nW2+71Rr21bkTiAsLhpRo8L2E/CQFz5py+oLn3ag+I8VXL+6pSzNzx
GCgmarhFUd1Y9rIyNtuEOLfUbBM59S6GUmUZNDcsCP03Vb1Adu80mCq5sV9FmwDJjHuYkgoaSNJ3
1GunNAWz+f0f4/ee94CzxrGvUNKTttlXMtj3jWlS32KOC1LeDKvVmEWdwhZGME3HpMguc7W4hq0i
o6Xv8pmEv4dQPigtz52/c6CPoKIcQbrZTxk6sxb7XYWGoTOx3Q8Em9IQ3MDCEe/mxjlX5j37tAjn
Gdsw76UjKTLeEVbTzWT/Z4Y/Im1QkrDiOTUfQhZsXqUDihK/LcisezTB4Bb3SN3wyNJaMBx6fswF
YxGxNDdrzZFDY7knVSD5DsPP8zYBp4IU4adA4IANj2I9dvJNCzzYiiZFM+Wpr+NDWFe6MoAKtSq4
grnPaJL5uY/MG0fnfzBPR1zVswiUFkAlRXneFIuS/zUSX5uMxtfd39wNxDxulRyh35hMAGMoV2w/
q6msx74DlyRNqPOQxGXvv1a5mBIYZIuOdcbYet/l3FL7wkTpcUgNVa9at9ZLLHSbwO9KmwI5rwhM
MizZ3xjdlPYbuhV/5j9KoNnn7oSitINQ4TXzsQc71xGFvVztcNltZZrdpT1O44L75OFsYCtdYyxI
jE+ZkFy8Q3Y6sHzkuf0rmWIKJdHoMP1khhZEMyZCll2XzuQruoosMCHP/gkok0ssfXf/sSsvf38B
8sbTYzCcMP2ROEVu7BI9rKue95HRgraaO6f87zaORO6idZCn27Psr+plA+LmIFI45shHAGKBTf3f
z4oTlpcy8Q0LFcm+75ljMgnlLvCKjucf6U1Vo4VgpTCtERncfdQzxffzmZslVWMyhJRjP9pdwGNP
z3M2GOC+/th2JPt9DfmLvoOL+l1Xnepf6faCsFyxavZqs7HFijyI8aJDpBQYfESRFlcFIaHVbDnq
XBKdPX35Dv3gpfex7UN132rKvm+k0PPtqupO+HWAVVmosEm72+5cyg9UrsYuSo2I6K+X9HPeubIy
Y5OE02Ja17Eu+30o9nrgbqHh9aHhbsakreEQHGz6OqqX6YwEq/t/xhSqQ7MSC7uhey/F3eyg1pkI
xuO6vxpkkpj3UlP2P1r4Xu37OSVoiVeL+FbpBET8nbSRinWr1+/Z/ByyWdRxRPjHMkzX+AqDni1D
4WArnbKSPs9i74xdkFoF3leU0RK6bVzGLcpVeq9m5x/VRqE/xZgCm8rF3WHut9VealAPeMD89r/x
NcJiOzHgIV75XjaVhjVrTZNyyYEPLh2aNszy7ZpPMhwMbmjuwDuKTR5y72FkRszx0wCqTXca93y7
PSsFPogZNx2FaJiBV7xdYDAgj5farNEBcyh1Tufjz5wqluZ0i/i55hf8qcvsFH2j765jX2edyrRa
s1BM/2pjr1kbeQVOZF/ZpVri62aYCR7R3IT46W7mcMbJM5lbtui2JjCpestiMiLSoIJJFgcpN5D3
0zN0p2mBkX7ECiRAOvQRAlE0LIClA3aKK34MYy/DjzpgaJVm7IoHB1FqtO1MzCC+dMRmqwyBBoTW
a2rdiR78ZJZKdToPCGt3Q7QrcUM7+6xJXZS37BfI2TQCi34kky8Gq/QoV2dREnZv+b0YZ2Fp0FtC
HTHh56KyTvf79OvlQlScFWBtQFBI27I8OYQ3QF78wa3dRw38XoHVxYvT4LWMrpsiEfh9ftNmlmYF
CDemrGXOrf8mpSg0ybNVXQPnzH9zMouImdgEwudpuBLVfNVr0U88p/iE1ofTKdumzV2Nzs83UjSx
AWG7b0eN69D62DQcI7iRfp9GVZaJPsasmNynL7iVDIDMcIXPjJHyl/TmO2Ju18BBkpOdoNUsaeYU
bwGRyvPSQ3iU1AdQMngUiOICSR9S0zNd1FDtdHpAHCnatJZxZt+UYCWHbnOSqYfe5BacVhZezwtL
Ie34MwgNw8sHAnTxCrzbFET4hh2qFBhkI5WLlQ4InCLjb3LAhp1fDJLWOIo8S86FjvQlg5P4ujWT
Oi4AwwJ/Hn3KCDBRKGPR8uBj9JuS70kJWXN07+CNQJe39+v03g+0dQFOcDs8mLLFmfXQhOVnuaNq
H+Fat7lNYR9XXIT3kJr5CHI4JuS9EEupP0pKSyhpmvwwA4AoYCcSG7JuZa9tIVTyVu5PHy7dcsut
UDtaMVVV+QPWJtcwAGXRlYz918yLvZFb2NVb7tKOJ8JvAqEfGCHkJ19ktc5lulo2SI8sDK7aVB7U
jM5tbrjRIqXXtUboC7vLRzyY513AwmabnpdAl4XISboZH7rPXcr8ubLFefMkpi1pi0G3+tyTakdJ
wk00xlkHh4RZfe5nQxvD4T7VmeoFKCK1sFLMRZScBWrD6YSbyTogQ8ofG9/bedKasZaXW9MVL4vt
fU2fx0i1H2/ZqTqbmgDNFV6QeetPtlBCfgVkCh2gLRZnR1FBJGneYaj7Znnc2X0r93jdIiHP3LAY
AdZoZwAf7s+xncVJD5yO+YA5WHcET0HagO2wPiL3kn+3XMqodTsnUZSDkXKlK5/u5TNbBE0+XgYc
jfN7p6YDAWu9e3h5n1vfdsK+KoJVj+xG1uu9oOTBme2nuJdnP/hRf/tuS5SWJaE7fR8y6KvMczCt
mnxGFRle1Y7QoiQhLwzvRNEuJAXPpPnhvkPiamTkJf1i3qpQhUFecIgMNo1OZ4yc7yZHScmfPE/r
FQvBfl5afGl45JkmKroii+bAk/iDbpIo25u/6PM1kBiF0TlOGHJfvRG68yrvigOqlP7++kNT61Hg
czNnBpP2GthWigf6RvCgRD+zrCuZKRD/LkQVf1i05z8lj3/ufhAMYMMI+7n7clnYbJZ1NCKtlySe
KpwKTHIcFsRGEsRblpcL3f5wBMmY1+XkECKMFkDoQErWdNadnNs+Jc7wV0iHmT7R9Xvi6Ve+P3wI
4wEXnR7DATih1wdNZoCJfixp+tqNuP2RVwLZmKHBYd6FNuBRwlDd2D6e+WZ9UiNXi8TA4gyu1Ey9
CE6BcjI3WWsXTAYvDvZmgZZOaoANW4pHYKDcijm97Ii6PkVy7e2gCLN2Ba6iBfS42VNjJONVQSR2
dN/qNVMdrk0GOwR0PYBUpfj+3spw1XzDiMfb/gBrS5ngwjCAiZFzZ5VcTJjD/wcNCqO7TcOpqKuT
MEp79x0YP+drlcDMpDsMXcPl0nP0Wqgj9EA6rwC7XxwVBQ29W9mxTBBpiESNQ6mNYDoOeUEi507J
JaaefMoJqEMAMvk2Tpnyy6YaeaoA2Zcg3B9SB3rTQptpPR7Tm9uA4cRsMvhltz6DqH5TSWRJOU5q
TimbpJxfnRvLpyvop3ILPK4s3/UjaefxPWnGRa97DnK3Ts9+g0hjvMFRSy+56b9xDOB99yAxPrSt
XKbkaMBwZi25L614h7RehaSnFqMlVqZMo8mL72aQdCmJBUYJe9tKxWWJNxsazwUrqeTWhV71XK5P
TNyc96IJ/iOkNHfqukpYVvzqr5CyL8KJD9vUpollbqzXom7yMG+ktN5WKI/X5GBN3Yzn7wcozAcb
WWBY28PHqWElA7tYSO0HfIV6apYNT7y+/CZOF1aPbIpsNf48PFYxytRJk/Af+Mlx7pjBV2WlQYLU
r3iOHBoVgcj+vyfTgTZER5+NFOwjlqTbDW8x0xiegc8ZjU9gNHrEfyVUEBa7bi42Q8B5fNex9MRf
PvirGzJv8Y2l8bs1HTKrsZ6v8MMxqEVVpdZnQNu83zmfP/E9iYNrqgRKKC08jRciFHWWAokoRg0x
0PNQ4V7mbiPCbYcuxH8NEpqTG7T3oT1yWSxDPB5uOGdeDUZAZsQtQr46+gEsSl3DKiXCc8pZOepm
35t7qNRr+ykLmiu+eHLopNoUhBAyI7AV+p0t6rkfHbIRfnrQsqulE1jQmOnDlMcOW6nCHLkkgafi
XaASo2NyUM+CE4ORz/lyXlqUaR6sas8YMmsnYQ7oDCECY2dsqTLZDqVOYhYDPpF68d5zcToA/G77
UPPplKAYQrtD/w+F3PPgH3gFQ3CB7HTDOFGuqEnHku59BFEW+tfVxRG5c69C5034+/ayjMLkibuk
eOlgD2Xa+W5f1m8i+zJtoq18rPMRgTEVdL3fUYYHiRwsJzpvTpmWbj9P61KuUMIRlwNmQTwYfofx
JJgsFFGwDutuVWhrNykWO2/Hxe+aEDeg51gUPtKmr+UEzjj/k56L7mPsWEn797+LP6iQc0rui9bt
3ldC2t1ssZQhukOfYdzzfT3wt2rsh6FusXs2Z8ihtYZe+37lQ3BSCyZax+oCYwpRkmRa6NNAzWAv
PnkfVzUzyI018IyFmFFvk5CN+irfTqOOaol41PPRfDoTpGv5tuIwAjLCKbqc95e5PEuqA9sm1MSN
6fZBBwOiFjiz5fwTNeoYBhmsh7RpBdXHiKL3gM074CxmoF/md1quUrKwHIe7BUWB1TKarP+G1Dy7
fBVJK3sPLVmYq60bkejQbVNNyyP57DcCuMtgkIKLTAzJQj1a791ioCLkinJFui8cjO9dK0hcVudj
44bRePVkXVBD/o0FJphGQ3/5+kmU7iMjAJerElOLH43ehcJAXt5wutb2bkqDCFCuwUYjkrYnigVW
SmStClYoPAW/3mBOWKleaRKFB6I7TUdrzjg/1yyICzxHYoJ2BrnNHzovlfZhKKYD/ZLpsvNG3UkH
9bFkjSWVC+cr6goSCWV+Y2HhqXhw2lqGPXgow7qN8NmAkZB8ypxy+0dE6Ox+x8MMxL3r3/mJcKg/
bj616Zp2RgmZuqpgbb/mMZktnmER3cFgaGMFBr4UgF321Kxi2TBSmTMF2H08sVnizRhyGlvZQVlG
Oxfx3U9Gbgt7SWUaodCXE3HJFyyHG2Y97oN3nN1kdOIyFqNKVczqykV0dN8zdbiBnjazFgtnNFLC
s0yI6BfS812eUu+dTCIANvDzuB267t9OBPX588o/kMChBKpNx4h9igfcYCVsv5dx6EgzYsJ1l7uZ
aJX8SxjT2IC1ZWS1zkS1r0qYT8bMsc6RQrQCzRVOzjwHPOObPJoJLOOutsM+XM+WfsRvZcMx4Mas
3C7IsqN4kpMbTuCFTCoyDy/MPMssO6RrUXoovOv22NvHyelOgl+nm68ebSclJ4TOtdtWzkg5ag1w
/Gkyr7wiELrEC4TiWbjPOy9jriH32XCKU1fWhoNSt1pdcprBUhHyOIzbVp5lvTVFAeavm73AMoKc
ZjFl86SaksP/92twxhVKl63RLq75KMIQPbUBS/AbIOGOlQIZZU+1XFhkZhBFg4+knmJIqvs1YOvT
uZGuW8QKxR5YuwLGMVd/K3eBu9COi/j5i6BBRuomwDkObW6pjDMf45mUngWni6cfbjEjWJoTZjGU
P1LgA3b3Cc4HWI+YZ6iEVojUsQ3YNRBV6JUPem1rB3tpbpSfsLsRPt39agi5Gfj5PA44QrLcbMmF
VBkefCimqO7+KIxqAO5pfi6MPePLAl6XK6Rnk2CnjqGJHGwO/RUNxSQElyjaMeDocym+ggILCRAg
W2kYElHt5wj+JqDS4yKDTYbfmV3fliXJFB6rz2e/Guxd/vj1I4BRmgKJfBAPYp0QYgMpMN599FIy
e4fLMh7qAzs1kZGwnJCWxzhIZk2ie48iiPCaPsKdqkk8h/W+KOSa1YLkIQmWopUHl66GiUBaqJSu
0uL5k6rkIdtWJJkB1LB5lq1QTHQoviW5B0JD/VDX1LVD/EKkg2uBQrN+CS+rQeQw0BDV+G4r34TT
7nF5RSHCVS0Nc90ylZbfHa+H/wVT0SKMGZzJVofIM2FZq/Con1Jwkyq9UiimRBnvMkeUkoZ0gjfN
kDoUX3ronA5xvAn91mG6nCBw2AxNSa0huQncTbMuCY9N7N/64+3AhIZdAGDlUuQDInnL8Bzsn5I0
8XoZnmXruQ68DGMc1UTuHBrj99zc7Ynce0KFl+0cd873sQXYNb7JZrAbiHs/Ms6vC9fgjZ9y2vgu
TLoFZ7d1nxQ+7pYI/N74FLhKbWhVmVHEoBjdJDQdhaujJWF5lX+vWqB5CyleeYdY6aO1hl3S7T/F
AJkEEl+QnI7vCDt/dSQs8xNGFNuXV5QGz2o1yQjuhAfhNvvBcPMJDnURKXNQAiB5HBqWdUsL8Ljl
EQ5ZExd7rge9zMouuUAfFYEgreblvBhI/K6eDdI31b3vCKDjA+kOfQpkiuuiq4RRVormS7E+8sqy
UTgeBMWRKoVg+GeigjiuJCsdhLba5yH5dkDlmtrJHlGgau7XolhBWYMqGx/w+6MZ/O9nucl1oNn+
KJTwATvZYFM39ckLLMPIbU/whVq1138kaYxiy0DDBCB/FGyPzMnQ2YuFDMtBkNGIdRyZ1oIYs9Hc
kOQDwpSonaRhXA4PQO0UHsZsdb8JJBahM2dIMd+AJrCqSjGCKJIikIeMcFCD9SYku0q0lVu9aMDb
a5u00C74ybQSnSPiuHToSMWOXW0iRlAuL87iZkGEVUqCodxnKlqIOXGLFrUshrEJtehOmBisWuPc
8MlGpAITnGE7Gw92BAmB+hQ9OWUcFUa20r3WnHl/uNL3+zPgObmWIQ2T592gMVvUaVT/utqu05Bg
51vn/SnTo/Irh6+TayTiJvUin8GaAKsPTlWdZux2aaVcsON74Tta3ZOoxnjeVqe627k+Zq/5vRBV
Lqus/l0NimrOh5VAf1RQf7yjjoHKaFpP744BdeMfQEavejSa7wMis8hZCFm5HicDjxq9OKSIuC5j
sdMpsoowgfeabP6X0EA1rY7/W4ygtml3KHG+oqMHiscJY3yf/4Hc2pG8aob3APGK8ctCu4uURlDc
/XSybriYDdSvhBEaa+9TGTD3H2Q5YfOpbAvC5zJZT9RlhXed8AXtKfHrsbWyNG6ckWHLzrSLrUIH
Cwp0EKEM2HLccgumsdq85LeK3+6SYfzQRA41HQCgfrwL9zxM3gAubFbuf3cilHqZEpcEg6BVn8Yp
G8bnh9e9zCEQuuTNzgWvJP6xyKwBJWU9gvHG7Jj7NNfjcWcdedzgY1sMwcxW2Va0+YfAsnlKPM54
9ELMqhBmPhvnwrUq3OIvhbVDhgKEnbOGiZQHzs/NbF08xdcL3bkWOVivgPQ1v2IWgFiqCRqHTZRp
Gy5TDA+3Oj8guDMKdbCQ0Oy+ULYab5YV9NkQKTLmYfJpF7BR5qAjX+G3amS3r95xt45VJVOwpSoi
WnprHXHSzyzmB5/3z4q2iKaTAtxUfr3FGSBD+7ZUnWdeQ93zW5KrEbMfNdx3A8fpLwzkyOQDpsA3
jGpbXJ/P+trlYhSebR4Zd2EKOeqsthZrGIxt/u4emi4FW1GTb9iF/ZeI6xLfgbiAn4KGRKIdrVJV
1WoLTcZcK5uO6J8bZ+8hR2m66vxx4vJN7Zkd1VZgkYc8p0H1oXFqQd2nMB/uuaX9vmjmalVSHdsZ
EiziYjtEtXmJzUAltJMri8YQYPnZJqFSZ0pNJqFnPHO54lgmIIyg3fATMcouHnfG37cAV8jq7Qtn
iiHioxcRq2eVBkvDEfguXZAxDWFsQEtQXnQDXSbJz4IOmi38Th4XZ3cfz9Pnv6R7vNlY2hpKizt2
gKATbWeePN0SngiZon1IOfbEpMK1Sgp8pzjNzY2uaOCS4Xoe1I0fO5+GUR68jrTrhrLCPqnZ2L+H
g/ET8u/1y135d3jn+lo2AOAJ5l/hl7yDY4kZ6XL+aY5fFZLDZSwoinSiTtxPhEFo7vgtfW2Mc6BA
uNR8aFWlJPLHjL3Tglshai24oi4M/crVirZDIyb5M7jIhJY0aljRN1vE/7yIueLCXvPpqUO/p4R7
ISm7FO5k11uK5MG9seLMbXoNzxBi9T7D9HFdyLh/uoRrI+ywzRg/Lou4LyPaBvXKtGRlBGCanUjC
/Bc7SN+rZVm2OEFc+WnOHfV2B3v3T2WCqnthKZm3VufLLeFbV8zivAGhENv24OAtTODTLn8v5YPE
Ga3QPRxmV1txZrA5arVeEO23SDjGsRfCW2iYkOuqrb2C424zySFF7hkVK7/fdiGFGsIr1kZ69Sk6
B0D1+hAYyfF2Il5TmE+6s3+IulQeGkMy1/dKD1N8kHTT+AOYYB1/c3DnQPfqg/0pLybONTmQApEj
pqfIauwRru1TI/A0UmSExgK4xSVjkzxNX01MkwYk3UqVzrLPz4Y2JVmsJThtDCoya+9nbwmTharm
JhNFUbWQ0iIfF9mLLCN1UZzMf525XpGdj9q144FK6qQJHtdwvw5DsFmzyVkeQV/9Rr2wLdHB+dB6
z4e//ncoJmE9bR8DRDBYcF35J/HLb6SCUnNmFlb2peUUA1B/ENatwcHsKWABiKrU9yIc5Pq820LE
yFZbS0GnIZsBbISlaPetI2shS9elDwXu1XL/kn/KwBeJSXVyNF35ktRcTreabNs7EPvtWFDjamKc
lfipBasIFzJJy54g9HGHGbrJItzdvxf4BMPnjM2qSz3G1r22167E03bmd4CLXryUxqhoBoUYllVU
+4fH2NcuitdGtme8JvBCfVap6ccpRtYbwkzr4s7Rss2GpJZ74GWYzNWrRCrTelEDr7lnDOfizDYa
X0qJkwS/VV4G787LDies0lIdkAH/tEg8/pfgk+yo+8/lBVofQyeiNIqeq4D3TRudhTU1Ig4Sq23D
1ZVN/X8R40dxcWtyDp6TvLNURIrYG2D27bJ+I2OMC5TuNlMWOPyuoE07XjiDAXXhQnNg/gZ6y1Mf
kk14LS5X4AIePftymlqX1iF3oJ0Nxl+U1tYc+yDU5yOHBuN1/yO8h1YOsekRpbQth3azVo9/7xVY
/+KniKdsWEdgqkd44JKmUhlcnrs4fiwo1V+HBW1OH/1RuVYiq7kgFC1vxaXcQ6whYeIJKUHaOrbZ
VjFKAE3gAUfHELICkIkXVIThOIeID6rX8IHBkktZnDzdPUq4X+ptSAvyCgoHg4AV93C8+BDBgn6H
QgvbbBDiyCOSC+QNYIrHdspk59C6BAkwQ8Swk7gKzsRClXXe6Vhc9qnXyO9EIk+torPqZewIP9eN
3rWpt9NbxQCwiZSHEUsLaiq+JzWm32ZmUe1Bo6+dnw7gQja2+5P66Wgx7P/yQg04G5Z58xMVjtJf
nIowiOW7aJK7EYUtcpvj/DziBFrOWn0AptI7wpHaiOymfzCVXE+S7g5LHmsRWxvMzMxnyxI8L2aO
hHYXtwxP6/KWkE9rx/kp51X2ODQnYGtMth1NFMvz0JLc/WsHRpYuoKBNw1LaPdb6PPvoryabLOhM
AH/5Cfm9Zs5/NNRdYspxVFX3fWB+c5IgxK3TVCRrVmig/B0QrkSwy3MpoPH6d81sYZ8MSf4P7b4U
phtb+A+Y0JDY5PEbmA5tZ8OTUYVEm/ZxMpSxobPEdkuDw+iRY/UV/sSgQ3pFoO3r27iYQpAU4OVr
m7hdaS0kHGoemdqRm4R0H4OdVzWJ0WEbW+CNPaQGLANsyvgve1Hzv57AtsoQ7A+QkeDBzEVsSaRM
A69Dm0Tu1wGMd6WAv2dmFbm+f1w49oVH0djeVUCEHG0adzgzRLCDaI8GxVX7KQiHJN6FklqU7Bph
LAotdwBdfYXfVlZJnie78rHVltosEZMaJNqAGkpWfp7iXfnSnEecsjDzpqR+CTWSA6mMtbx77DPb
ApatHo1OCg7tBddAYol3sQ75G5MmWzJPpVKDt2qNX6ETJzyQos1t+cPraqB9YCw5Y8J8+jCVjq3n
DzqzlnrdWEKZZPKL/6WJPcMGS5HnRKarROwp6ZDfSx5Cxb/eUPWQ2G0tHFYd/XSdQkm602wZrHMv
IfyLaSg+wXILA+dACB4U/YF21IbhQ08xVpaaw7mTbP5pCrNQRohs05q8iF2oOLvjC+P0fBmRa+A2
8na/fIPqKizGwO2+8reneCYQvC3fR3Q/qxO+tu6SgmQBJgVCtZMd68i8Ocasi4mVUIHm/XqEwDEK
zwUN/dJo8WVFVmnaj3nfa1BCCyzdbf0KKd0ZbJDj+DB5uyKWsM/qVBX/JZgiipzUq5CzStT8hhXA
0KVWMLXdQ+BU5WbNNziaSJHYJZIKCFK6eLnO6Glbk8JCdqO0+4ipX3rwUu1cSmwEjpmFyklIln87
xSBROdqKmnOyWFr7L22r7QJxjj8Yv1QSj23V7nAGC39B23h5W0ijA6QvWcya3AlJyaItYIarLgfN
RA9mxpU0oLglmFWoxuaeMx+UXAt/e/58sKtW3XA/2oNSEJ5rCKfSrqlC3WI21rZ1eBtAufEqRaVc
RjJUiftQlwiXkMKLGDUCvksMQcmlA+SlByI0L7u0/mBFPa4Up/J9U2F00ByTNjYEpP3g7dIci6MJ
AdMuSTUwkhptdr02LjCLBId2CPsiHuvirgGCf7hF/rKKjbXgkf38+gAmZBwTbF7Ou9LiupYFI9C1
KTwKl8lavyCxOfKbmLnZFnf3OyYMCDf6A3/xQwmw5yFNgu/23M0YJe8yWc3TqBd6uh+GEOle4McA
2Z2+SChs8XDBiSI0xf24B/1zRW/EtyEds9F5JJFiiYlSmWsW1m4tC5hMEYq1KLET4Am4nU/Vymmr
wK5zdOu+d2NXmVjuzy1wnLItcMOyreFkN2IbFTqqNfjupNexiBva7BfIVUokE6091yflLvGWMWdI
8yvLvcg0pRCfOHa0PDJMvZwC5pdSm+mXfeYPQa1juvD/YJhDp48B/7hGqjdYn58XK3yJKq7Tf9mw
8YAHnKovlsKKcjor3VdKI5OcsCP2BH7g6aCNd037xv+ii+9rr1i+wOqu21w0HYINHlWXkw3fhGXx
uaczDo0HSs9rYJ5JfwYlchASOUEWsmBbmAeyLeuWiylGUtWFp9fsyddTzhrTWF2Ty3PM10ZyH3Wg
G5+XGwhTdApybKW9mocdRdD9sSsYYAKRyF2LtHf64XsNsjy0pzKhWeiLn+nlV8LfFyJK7ztWSISb
Shu6+ZnJ1iLASHsZXRBLIy6F1RyJOw3czwr+YeeGyD4l/b6EWSvyN4M7Z3PV96ZKBIx/DER8ePpB
trUBpP1HRH1/H6+t6gx4hG+rKjNemY/8p0eqgEfFM2CMAeEtIAII3w0rWlhXVZaVSpGPflhcyHPP
tYSN58pz+TsOSqDKQYaj7MBGoKTLY15A17zaoF/mSKfawLDNU4stag56Vn+oYDuFyfFypy1vS0Ws
+mE/nMAaOfryK/hwhMdPRLN/jH1c05lY++qDnO6n9IAON14+yLZ3tzOI678iwnxhhZywGQP9HS54
kaYsFCIrFdAbombkFBMCE97tT6DyfrAiiKFiyapNIiOa3i7xpL+XIu3DEI7L4D5mKLBkAuEygfoA
GCnqcQm0V30GRslWcAXjz47OVfSSWa71AX7hi8NEgfxVBIeaUFLBwwuhPFBO9ZeZTmwXOo5H85lU
Pfc4ypSL9m7KKNWpHrL29MFjOp2EICPAm+CCLrbuec4EfNHha+lsPHrFs/exkDJp8eLTH3Vs/c0T
oRzxPndaZubYSzgXymq0EZ9egQgrvf4JUVNZMuiChTOGSpCfiCyxe0CNhDwjwIRGsnncEMIhi498
rQmgOyLz5VQvphp6l/qAfLyrVTDz+tKsCx3sCxP84s99iUHXiBxDW2d3/70VXAbSm/lkvrYYE52i
3Jc57RgNCrM4A5/DisCzd5XkGO4SN5d/Xs5z+sxF9AO18KhxS/4XY60IVJLwv4KNoZ/THFFeo2C2
W4b1Cgt7Uss2aMgSm3fYia8lS1X0H2UoYWRmnyBE0L3suRmaSMr//EQoSpWh8sh7vEQdEn7Fb2gK
Dt6ssglpYM19tdKBkSKSUP0h9+hxXGC66Xv1iIMGZ6iW40JOMnWZ/vXRv4x/xJnSgadmlYa6BgSX
V1lO9PZIfxIhCN6AAwF4zrGVvqknGpTvAVJr0/tLCQ8PNHBvJaSYujj2ea5Pg1yl3BWZqYtG4xxm
kzLvG8cSi3eSpMurMh/nW1qTyS3JLqSZECttD48EskCrNB5jK324IXkyhmWRqCAkz4i9/RvYuaBD
+Ii0sDcx3QbZuoMojbQmL99YgcvqVXxnqJp1YUsyWqzClAKYIDDEL+aha4BwfZ1exfUfJW5gE+ui
UA6Q94fH3CzqumstjpAai8bLgbR2FalFJWPRbFNh5nH0Li2Pqr1FOrMx1/MvoXb/7T2Byxt1mYWp
UjBh+O0CNJBUYpsSp/g/PRItbT3O7s5qco5I+hPJvb7X6x4vSKb1sFv0xqFYg6i1tDzAS3AtSll0
Y0A7RnpAZZQ7XskhBIjAGE0LFhuZR5DF70yvCvSMfASYfhYFOToMZQcdTNyHGgxvScuEezeTs1pg
KeuEepvT3xVTeosOAiaSw9xz9zbm+1SRUKUytUQwRmym7YLwwyxZjodhhucUlVzeb5aLfPoZ8HEg
Tt2qbOYeF5VUE9Exica89hSQf8CLK8UMEhiUVwlv1UtGdCmhs29E4o21RfDbJtI+jZVNOJu0+6xU
fcXbwSbo2HLvHC4UzMZ1GxRjV1ALLqQCDpNJs785YYVnMFKUPo2EOcaG4FwVlamBEIa2PWHT1Ho1
U0EZB9VmICFAh7ENQWxGo5Os8vp4jlgidEQ42dfAISx4TdnD4jxxQxw1PHBCqKi1yiLAWqdZkQuj
XpLNOvwmZo5PMb4KyIekNNhNjeV8hMSKEzXto+63Tf41qJq2u3BTf/dvRu6lJ0LowOUY6BcsPzZF
JCuUD5zh3Fja7rY56UwnC4thbMUEtob+pVsaEPqVrWulTuoHYhrIdD5ZUW+qdND9WsG1la8BP8rO
0A3nANvs0EOjw+2q3ryUlNJHDXiRBKHK5I5+ejSEmbNitMXZvEIdBhl2LUH94rNljH+hvWbqFslR
+n15pT1MxcOVLJRpJFs2pEC8b1zwbb1zTxTZjd1Ny5wAh/0X7wA21b2zN/ojJuaeGrHmu4EKC7/6
WJJ0x/rx/AGHmXgrWdBfISqF4sRa/x1U4vb7+Xl4yx3u+EFGQdmKRSVGcOTR2hBoMnMi1SCkhj06
d3TiXsXGjbp7U2d4T68hFynXjUmQ7/AQZUXyNLUDLTsSYiOr+Hiu+sZrO9CS/d8QrCftlkd5xR5Q
AzI7tET8GDwemGpyg6EnR240OTRUCnKOcws05Tdvh2kIqtjeQtdamwXeopHERV7PRSMtkZkOYfBC
K+O/PZdVDl/H3Io025sLqDEgbZStZmSquSRrtujtIEfBrI1bQEcE4wYq/gXfxlDryoC9tYB93h2h
mx2MyeFQD7tkbHNakvMmrJstlp4FfVEv9Cb54PRv4RCqxq9aMqiLIpei96o0CdDV+BR4iN3W9eM6
IQDsVCd6In/OuzZx6P3SY5YEGYqD3iTpdzbzKE1o1tO8hcZ1zq8eRv3XUYSQ1T0H3eyWEvei19ik
8pb9alv2bPS2xQ+W9vtM3gG05ByjI7GfQ+rpb7jQgePWhqBGRdWDw200k+tTt8ApoY9OHDjjfUQs
9MdOrwcqkuyObJ9mrVFv9qAX993X4OaArz71X3JNCKqbEoci5oaZgGPhO40dg8mQc/hP3BV7ApSk
UeWuNALjekZkHd6M0oKv2amg51sRJCzhlkFdFW5u/cutLpk2M33eQMl8YCQ2USx+9j21s3fCoM93
ZvvX5fGZRkZGKKEy3kkVr8ecLsE/yYBbiKz0JjI7XhDPXy3geohNK6/sWJyEeStO/5k4qbzu89Ly
vQfuZyrCS0cXV6ud/SCQd9JAzKjxHa22ZPrROolQVcsF3sjYVeDCG8MeJsWzA2SEcH2vAgKpzGxc
jXp+S5MlXr9CW724uDJhJcfXCJmpJxl3NHG8khPbGCTv0wpUIrMMkWAUvDg1+bsEe421JjZcJsP7
YUi/t8jhmwo6bQi5KTKREYtc0rSwtkphWmTjvA+GvHyw7NlECpeMbWXCRJP9euL3z8ZBZzNw7kIJ
a5mluixxQ7wKDwGfV55byuNFUOemtDgPimnsLTBV59EWEjzfb7Ckcy0tHjDZ1wipjwvPNwjwsBfr
41LMrFUyZIglvXc7LTV9xi0h3m9zpTVXWpTzCGcVQVDgXKEBepingFvddEaBMZrJb59DUYD6AWe1
Ikr5GwOPwitRafzCB8HW9kLIvkWq8Hje6QEhq7mFmq+ZBGK360a/vmB1il8IEp0ovN4lzB42iK0z
QT6DnsBs+Dd448Cde0BIkpM5msMjFMYsAPSWbkwlGkD6TvGUK2AezlO8E553UxdUX0enRmSgMwYv
sJaoT/hm8TLmxod3Wi7EZ5DAJpzK6iEHAzvdn24PjAspM0ARZC7fJB0ChubHxGW7IhJIHaTVKwQs
FVuzG9MRAcHhV0IYACI7DE7MMpRpYINHcSNbV3/Zm2wXSSYknhgo7UAjYbNqyk7PYjJzEccRv2PD
xan/VVtwXIm1uKycM9o3tuS3Ji0E16H0f8sx6aJkklFWBJiNhykfJQLkt81+N4qquKxYz0NMb8lw
iunhva6o1iNVZDJ5YOYa2XHyZ+Y1VbTrDk5A93j3UBdhO35KC8vWdnqkOlseT91w2bemcA87fhd4
j4dOprf5YQrfb1tRMFxaTqJzWAKkHEWbyJIqgfLZC/9hRBev6KTnO8lmeZTiZTAsIo2t5JoWuBW7
KJMwPpBnY6zD5FTHsxRWTLaUQNfhYL9n0sFIIm7ssNo9qNEdeIwHWj9R9UZQCsI0QyE4nCQK4lrQ
GUzsiwzVXeS5IHZux/vNtr1XjhuDTy9zz4x6f4+UUyl9R3arGAPxK3SCqQROKqMMeTGvOs4Q4kS0
/PjXjEpq0A4LL4OA6slpJdcYSWj8iGSwOirqTmuLslqOaHhSNzVve3aFsyYOXl0z16imt2l53nd8
/5ee31Tu1VbVrD1DirCzKhEx1pAVWyQNiJ4lvcjKPgXNFOj34iZhM330JzR13qNLhMOybecVw6id
oQNXvmuBxjlkzXSKYp8nIZvdf0VHodSrxs/k6Y/swjGDaTztGJc7DptLsURCr7uLDyCLEsYnx5BV
RvJBK83SP+1S3mCJh1xeMNxJjJikewur3VsukpeLGihXooqDPjHsTudDL2XiYUiexkBtzwf/B6ny
StL7Yjjpcq1kTEFXOenwvMTvstS4WhC0dMHNoDeSFbdkT1fdTLyVQB61dnYm0qawAYeau5gB4FnF
6Cqd5wlbgkffC/54JvdtP227iRLJG56qsioqbOPHhyxVd9DWWcadSd7Xidrbf14dGFEC5j49nSGq
wPpy3BnK3KgLy+GNnxTB3RQbw8F6g/XPs3ZcVu037shpK67xw3xj/zweUlJk0duc1aSZPNv0Al9s
B/2Rf2AAvrgp6k8iyFticv3bMvPakehtP8cTbufRG1iqy3d4/VXRZ1B6TkR6rGRfZpjd6vwFrhCW
u5dTqrszloAhtJnOSFP+WwqMIsGqUw0Me6+6AVMN6jea8CbleVU/FZzgJgr7XA3Vgne5SKmAr7W6
P4OUww522BQXhfYBD+iwL7ceISgdoOkEjLZPfXbhLAGSRS2BghSxa4XDCgFYDOyBp1CGwVnHeSO8
C0bQ0jQc4v0K7Cpx4IZ3XZH+2dl9GBJrtCrr/EtmLrDKAGIKOWsV3Nofht5X0MeTLXoea4/37AHi
HBzUrSXAv0ph9MOo0a36nXkNozUK3OLJfAQnSq/4v3MVEwok7PBg5zgeugwPJBia5oucvzTa1C0x
rI5phNMZ56ZDGNptFq+x0DXOl3es+ypOhoEUeKgG5hGwogZassjEwGc7JN4feRDhjuZhVo0S3Ttn
FoENsw8U8cRF5WVxLLh2oBGBMOt82D4enBiEFA78DmpbiM83WVht+Z2bOlzyQpSz8YkVcspRTb34
7eUyJ9MxhpS3Xs+BzFGtkCI/7dgV+VK5YfnblkEYiJLUW9t+Yl8yVnCCXe9JVtH+MJczHhTyAsXl
DRdNFAR0TH913pK9UH7olfGIvglxSH7fGmFbmobXKzExUFOrJM+3w3ej8bFpJVVCc9sxEWkf9Aq8
mIAai/fvpDFbmzoVlnZWWLmHJrybqcg+PGeoisf921+aIx4Mxdt5jxi2SlY9Yx5TMvF3qEMNYvUp
2xx+CXrMQ1YZYjws9ReSJCeMP6/3E6RnLvG4cnYzMX9R5O+E+GpRnCoOD/cwHS3YkGmTlx70Wi+y
kn6UySg1St5iGywShpZiUN84GKcOILrEUdRvc5JNiPsXJtFS6g8+7RfniygxSFjZoB1WLPIV6Xnw
pM608lU9NsZeIPfL9T6YxuipymwAP5v8XltQUDA3lBV7IvT29rMb8Qobfwf4AtTjlEb9sJ3e9rOt
djY9HKzf/AnEx8HJyaAk1cTqZRYIMEIuims+y1AFbJL6GrmCa7IUAVNNOdkGHjx2R/o4N3jJUmIO
cWZsKEaGj3L8Ie8CaNGCDwatEmBjgdflLFK3FEY2mTXrGO+7HUoaCVvEk4fp3uDPgbv0YJ2yJKQA
UC15RUkH7o1YcvdldwOLPGj2zVe0ZnJGIGeOPS5vr9tc5ZxdyICMIxf1KGxbLgaNNoB4Hf3WEikh
ISzMpcjGCrR9+e0GwPWQzW8HBJy1pH3iyMH5WUCcq1tqDErc5z+tPHxZoOK1IObrmpK/ExqFegEC
3h0iOZ1tYclkLP3I55mQYdukVdd3ymNC9mcrJMGAxqUu8FoBzUH1tpc0ogjE2CkFfg2Km4WpB1bE
PcyU4AsQGwKEbySUIdNaY72CazRWAtjBRnhDKk33BytIPPe+G1aDfTUhsQS6HEbcNvphZ9nfA8bx
JQNkIvucva3QFiDSjkTnrYIlXOU0he9/X7DSqw6ZIpWvVrj//E1NnyAlRncFRVBhYDq0zr/X4spC
Te0Jy+eNxM0xB3hY6gTLPSAMfBsIVXhxx63hmNb6MRDfMnSZ99Is1YKoJAfW0LlNBOtG2Vndc5HT
1sk9kDb5/XIIy3p7t1Rv6xOwFVr4v1IBcshS0fYSOxK/TgwSbQALtjVUo7R3FRUiGEZT60i7BkJH
VoXtl7lzH1ON2jJl0njxjt9eswjS8nLEbACO7JEALe4VvUVBSX2JvxooL3fDgvq4WtO02LFSxrP3
7o5GfivH3FZ8ylhcxq34cHDcwNZujTVVfFc+rGlzkQJcy1s5cBz+Tu39NM3hNj8MwMGDI+P6QhW1
mdeyoaJMWEtyo++7NKLQK1M4MMysVuwjcdgsnpUj1qBr78bCTt+bpQIeWaxHKFlxbSrHPwwlATtU
iEI3166J/V5fqtLEFCiE7ap5R9rUTR5xC/ulafJNe8yWvq+ptkSD3tNk+iJHsddYDfSXmpAAdLVG
ZHmqJa997HyHeUYPKttnW+wie7Ma5TRBIengmBk/aGoHHEgmq5JYQkl2CwXZOC3JQo37GocNw34A
LIVaxpGfZLYDGb9gONQdcJMy98gCKSrB+2bqlHCIRC1dvgdD1942Xi5v1lyQYBgGEk+Y/lWlGKs3
PiI9VqQOyADFNCjDD2DAertay1wOoCI3AZcbeIF4Yx4V+VY6MfIQCKFOewykGemRDOD6Q0ulK5rt
xLGM/tOoISA1vbw0iCASRyhOsxAvbQgtmPVr4fTWO16e2lJDUS6DykqLMzEGDoo0FY7YOjHQgTrE
HW8SotPNGDVkCWPCrXESSN/IEqgQax5O0PfP4qXWS6uG2LVkfmpy2VcHUQq89Im+b72M2G25o6Zj
XpiX/lxIPj13fgUmiH8oLXAyz0M7JzgRjrPcc7VF14IXns9tV83y2USsRtW3lMbBUGd/4KviwLmE
bhu/CGTIvq01i1rm4izmMVVt4PfVsxJcmWNc14+vlO0D2jOfYGI03Fegul/4YL7K5rHSlW8qhZ/b
6/PE0LwhkLPZigKEShytH0PmXRyTtReKXmIN7k3IQm9qaM2TvOxeE7F1rk1F+nWD4KykrcH9qunD
jc1D+g9EpEwHP2j38px5KHnKavzomRi9IgbvbNFseDyi8fCxG8JsBOXuzhpFtAGLrZ9IXYfugh2V
EfsuGy8FsBBiJwoUhKNNmceB+f9S3eFnl3AY2raoFwoIoH+9I5V5AfJhU4md2U/eQ0dW7zNyaGf2
xykWdAOaFjkMK+5tWsrf/rapPNpzvZ0DIXFVOe5bsug3tp6CCA5UpfzBuikbXhuyv2wufIL39kqr
TvucxbCdV/4Ojcc3gUXseA2N7cOsZArXfX0b4Ep3lZt+VFwi0GpXiZqOQB/cF+KGbDekvJ9lwAIY
KGb6HSZe1Qf0EPTzMjMTucI+9NZJReJjb3yU7urukXXX+4z9bF84I0XNlQqarmutmPenOHWJAc/p
tLzylBiCtKe07UeLNWE0sZLo2zqTSmno+uvgfvLSVb0KFQ2v3acwneSY9r4Q5UqVQKVljljpuv6M
FiIvltzDrbWlJyMqNMZNUf4yE9XEhNV5hBD+tSdHpOInA4Ngntx8SK07nZOIMnvqpDRXALw8acUt
4TtDq/lyOzlINX5TtqGj/Xa46MpdUKKB+xXuDyoe5WOiPHS+wdETbkzz7KFFBEohMxWDTy5YDKAa
71QctdHfDeasQVaqY6+0WTv91iUPnYYfbKHbEI3vn9LSe+/QzUQiayj/ddNnXXW1sVg79w+OHea8
aZJeZG0JwPOhbKUXpzW68Op33LCLSYb7SEsvC5jPaJLS/in9jpMKVjN1a+6UsdCTCIhqV4pgIEBH
XHzULwHKKKN0Jj9UgEL0mggLYMJlZZgry7vNhz2oonITnMHTZO6QmVbxqQOJMHuPyqVPtQDEhniQ
isTGy4wqH8v7QYE5mdFYJAEtGEDwkQEl9KrT70Zn3L1GpT39DvObdEEEy2FLsrm/nOm90fCNqVHe
g1Wzscrq9u2fLaQHXu4azeK/8Fcs0nGcG5tTBLXy4gQPSKS0w0hL4Fm5dMAmhX6gRJhbGjqGwfnC
ANFk9+vAqDzfpPCzLb07NNGNb0Iy9gt4/p2h+malcixyl9N6jog0b0eGrCRrI3CRFzh9ekbuF9uK
9w/74U5BOdglV5OqIkEiafzBre0hUf+WqyJGJqZI+ZYoOmyRwgfVlofSo1rJZVq5Hva2pHEYx5B2
G9CI/OwRbIdkL/80ZSfQafDzPKg0rmnUCXUUhy9se9FXKw62Y/DjCPNPaUlUTXi3lzENsEgaxWaZ
EXh422q8975N0kzOMtkujqiC52n1jB74al7vXzjzGwobXNIt6P3Rs9eyCenNGuIlfX6kTUOpAiQn
2rZw+/RrIpN/PhcPrmaocq/l42RPxmHKQ9gQ5QMgaj8wWJ0/QUPSqabeqALApW05EJzo/ks0Y7ZH
G3C5ui1IcdwKLqVUy+CqRQ/xcVIfQml7gpyRejqytYxgDcL2H2C7MFgsvDecE3yi/v9Cq180PKsr
rNriMpsho5K8tJRKQNcNar+ExLWelgKaCHhzvp8JCllejVvD6BOmPPEnz/fZzFJQNDEF+d+ZQhOB
GwCjCs5KWeBjMxe7iChzHWGyzxM7moBL0hd7k+gitAnenohpCxlGgTitX8MlvdSnmjiKKDhPu16q
8Ap+kipbKQCcw9+5tnz99mPw/6gmzuQ5t0M37SMy40RrGQ/SASaOFEZqwQv/IZvfTTfYkvRcQZgG
hYqT9PxMooUfP11XvxZW65xvLMT4J59vaorbEczQ6aHLqS8tF9EKsu2J9O0PGidqYKCFU2H9/neL
HEtmndWq4Ge5euEHfIdZbv5qSPlTMLEorif9uwtnu6sX4RFEar2Cpr7TTWLBBByD7MrMvAoCSu9P
y40fkYPLSPfR15DYItaKSxWKcMXdfW/RX4RqzCb9qEbGCWRCvWp7qYAuAEotZRTpU3JVs1n/rt6k
3zW8kzeMHea57UdRTXJy+iuFshELKX3XPAoGNs+XbpoBp3ZL/VDB0mqdjeIj9zp2M37/3K6gDLV8
bZz+ytJGoVgXl5aH5q19EOaLl+tnxxSRImtBXr99gFH+1gfx+8vfmiYoKce5xVL+Ngg2SaE0qzCm
7s/YLP2GYIwcY3a7/Rx8srVPK+E+3xfrik/HB9asqx8T4ErtVjWmd5ELemMS4W6kgqG5zynxnTz0
6VyyGZl1PysjidME4dEkaEjWEDy21xMh4W+OFPkUJqytEMFluH+wmL8Ydvo+D/GjfJ80pfCqcmV7
GnJGAscg8BcSkadbH4KqAwKJCAtz9ZcSIDX2BhT78JAmKhqmU3MW5a9mOZ4BtZiDWrswn4ME36Nf
qCem0p1PlFqlGp926/DTz03TvlFAx2mweCm6i2VukCM8Tmp/PoYPltM9TcvkvG20xKN0ZEQ4oUa5
N/8NKh+ilm1xic0jvGusMaQwnWV5FhB4rKJbhpNd8wp2X8NXDvBPaGiihrndkS571qNMqVWc4j73
TKm15ansxifVzfSal88qjVoUt5ytHSmbghi3JQosX+E73/GxnQ4tQScb8zYdXIoHJ6vGNPzuD8bL
m/hdHjmhVL34+biKAYvq/Quugd3PtkZtk6VzLpZzQaliOkc/AV1bdpOnfyDiW1kOdn0MONZp4Bcl
Ns6n5+3gRhhUjpT391r2/vRe220XKLY+uS/hLZPG+s0m1B0CK5pEnoi6b2I1Gt3AxwDa1yCZX6gg
RZEprprdR2qusoMZPtmRDl9+Xhqrro26U0bqWqlFiSmwfspbX8lyRPsnefvnbb04gqWMtJ5Ylqpk
QwfUg6azSeQ2UDljAExCw1845Po8CEK5B/dP13cXUU8ORg8YQ8osc2V2JkcRuUUPX25iOuVwTyOR
zGS3XqHsqpxLDoQSE98Bul/+ynusF7AefZkcmifNQEB4nIzg9eGuH3zE5s126/Bpo6qVBSw+7lR7
yUf7iPZf4slADnbmEYN5YCH0OuOfejmkwHbRtWEmlO7EXkIDQLLxH1JCQcafJO8KaFTtQOo/NF11
IuRw6HVTO6bbuHa/VwwwpksILboHLNWcUGygQ/Prs6JmowFvt0c45Q3xlhKGUS8HonlsiNGlQgUu
YHGDOLss/7rWT4kmrMfP8SW+CweXMmP+qSU7fy2agVXb1PHdmoc38ayLGx001foMvVcIqqk25W9j
UfMvrQUbX8fHZm104lS6JaWTz3S6VUFJtalFa1rwH8GZc14kVIJKfFdXnK0x46F39x/0tosvOhFH
TeopaiXEnwVJXFlGWEsCIED8cK+2RFF2UI8xQwldlwdVQgMRM7LSDECiOr5Nx44ETLVL9+0pA3rZ
t2WdXn7iK4ID1kd5jEtvrqmpUZCXITScEOsCUDPJy/wr/VkiE5kojCksIc3pojEJQS0TDOikFJ6e
/32jetYk3mUQ+66USBa9Q8mntkQoBkQdpVDoLt2D14MmHbduQrFexnKkYj2bvuRlmp0FheeTu0AS
4g+4OkTNiQiosDsx6t/N5t+xvkXR6PanHT+ehqSKqKhjYbhtNazG9elv/jpTU0PtOnLdpwRVeanT
CYgJ5kA50sKCpe4oe9CZzyuLs9BTk/Kg1tHuOQbr2p4z4nkXEYx0VafFg6ZJTs/6mlfC62ZQxRtZ
XgHqlHQ7KO/VW9VjrxVctFs6vBhmCtmP6OQML85DFFX3i8cNtTPLTqHYO8HF+6z/ma/q/mdtfjDx
kJm2gqubjq4njL4aBDTRJ8v4IQWe3Da7GSocAgz32o4lKupdEmogRRW/kyJl2Ok4vo0Xy8hRugtn
OzDO6sClfxXEex34gALRm9Oz9uMsQbJWHeKMZ7GFZ2nyjuWTa3HDZ8AqfiJyDMbcROGRUwCfIekB
IMzxH71Ht5lQj265+2bKbQTZv6rF9PbNPMRIEeFjGhDxyr17ZL+ZUlLz7RV1jQubkH1am0haSg10
s5OwpLpnRABBdk0gmbcEzoNRpjMUbDzRRdDi/NXB0XlEwavFW8lrRZ4Itcock2meoGlBLWWgsI4E
x2Emstz4YbvI31ME5H/ONSWRXaZYpAcbJ4aHpBtFxFQbHe9rRNtirGo90iJxmPoVk2pnqPbVLKoA
GIvM4MT7RN9sT5Td6vfyeHYzYzgn/QlLPNXGVDV+4TbkHqdpAyr9qTkQrOr1ARQSJ5op3EwMYAHL
9mhDlCxlIlICxgrdNlft+ANcESjijB1Uo/Zlqo4Cut22xF5277MV8D3g7Bs/MdnPKpa7sHOZTLll
odnurbQumuevehI+z33HmZF2418b9BUx10Q5mqfvscGBd6DC98ooXXEFtfvG416dWygU64fEMFtW
Lx7tHvz+He4U01qloJqx3qLnZKX6btVdZrYFnZ8d/dFl7e2rxXLRrudKLmHjzE2XMXkPGoa1+pKO
enkqz4fZD0ncFOWYwK33dWXq+BiQJcdzwdouzSNK+zBHQ/IFQakZ2pKTlX9l7RwTLMXi7FDqwD8U
H6+DZyG2F4Tl+8IC/zPOGAplPZ03Quc1Z9hbf0ih3g6T/7nNnbVyhoUw0t2nvEdd9sxHKxldLwzW
kiBtRTxi8lKexgvl1ryqUHHL1bNLVVYhEUtdk66kOlChdkPqIa6TfQ792EuzGkq5QFB1BztBVNp+
I4HjJkb7QPjecArxWcRiFthOpMBzHiEdZBMMz6cSpq9ljLSn7KfKDAAiZSTA2yEjQNyFi/z7QMrc
8VxyIwgblFtu6/QVTiqAyQK1CNyirFaVN4Wf1pukLLmXaBnvcvMJsBHtBG9xPAiT9XaQce8kr/F0
XD15btqUUNc2qw0ZS1UsTrr/qfRiVs2eKqzBxcJmTS56ZFnBH4CqzC1GRh1mw54ISL1d5LtJ+pJ8
f6BfRT2kqG2SCJlMFWTcLUqTqSGKvbmatuiRvnYQ5cgcjcODuZJG/w6cURRtD0CjpPZuPpZI3D+F
/Ne6eM6KM6L/C2TLH8Ck0v0f4+3UPECAsXcLFURM6qgDUbfNAQN4mB6n8GbaVDGBN/ixn0+tDPcw
wPb503JV2jNrHc2XBFlGRGWgxD9LeBnZ2hTU3T0O+H7+qYEyA68aUBGrTxZqXxs0dDCfC/3K+zNj
ZfInhgjOtIvhshEJcDmRMVnpn9wr/nlZTcL+YEz5fbJIf6XeTiEe9dOoaciAoAtqldZ++hzFwDrx
o0VKS8MYd6kLrDRSxVMjXgMQ9lrs8rmeq+hhyMRykpN0Wbb/CtE85w3GWq/QnislaiuAdFWDHHLM
5DKjg+xjHG57DlfduplKR2SPSn72A0F6c6ymfIB0Fh4ISVH2nRLy3yh3wwR/ddCNZUxAlzhXpFR7
LQyPDoJiaSyYSWqWEF4w4JyblnbK7CMeLz3nU2/j4LChycYhgmkWt4yUnbi24retVytcLJP8uuSm
PAtdAKFqggShk4xW0Q5kTyEP46kJ6SHJz3LZhTF5gOSqHicabSsDR06I8oymCi2HwMv00BXGZWS1
toYMTQ22hDIOmEBdDPJ9qOcgO4yfjLYC5PHhYWbjtdXYtK5r8H9KIJDhVyUJn15W+bYRDyF31iwz
jHViILBkBRHnM45ouQgR2k9gzDt7iozPGnSO5adalHVE/bLi3So8ow7WjlkCQTq8SBX8OyMTgx5d
xdRDTehiwgwogP8gJC6SoytKU0vuivbNZWsAY5Fuemkkvev+SCuexqAmnG3p7+cxWTN/++106EZc
RuxNyEVRd7frp1hR3Ee7+2O2BbZz6RsfMhcST9D7DY+y+t7Cx/7Zy5azROhGPIuiuDbYkj2IJPIg
sk/2dbn+xSMv8QDxlnVN8rWDiYeL01GO+nakaBr/2FinI7yAtYTcZCe9EelKWa5GTJsO/SCi2M/N
VUEbaKtB01HST8TdOURaSaLtMy+YYrmEr/uK/xy6C9tIoqu39DrkoeGkmn3y9zKU5bjB6ytX+n8m
wx6NzuvsPhMumxcs8UP54fIfoNxZlwbZuAvm+V7/J9xPLGXcm2MbrkdJbiEBhdvuA5k9id52fzH5
pGnxGYIYXDwGLoCQZwZQKgYFkfUjxzkCcBEuZ/j/b7UUqII44SaktDoKJgw2TB7+NrXqrrm0vTNO
J7afZgdQMmAKApwBIGmMF1nNLLGO4HYYpuCzXOEIe9UeQq9YsOW+R/vYuWB6s8zYakBjgZ6/M60A
nfya6RLqylzRaDZtfe5kq+eEy+cyKPGRVdOhDlQ3tch7JoAhFsH7hw8fn8geQtCRTT4F5njF6yh/
+l087gegVbwzMG2XHOztK+g2rkVH5mXTf+45r3/mDEw8uGFwA8PjmyrHuywsSRERVnPnCvE1Y7pg
zLODBxVdLD6tV682dcAt4Gaxh9GNk/OrOVlShrYjcab+1ekEYTG9t2QnoXX0XpmrTWRkf4k/w5bW
bNaDrzpietxOHktiBHWuc9QpmkvAw0iu1chOcxJSaIeXvKM28V6lof+ND64lMcTqYqBKpW/a+8Ip
w3IMb4QtUJorApiR8Vww2vMVVoNZSBPxzoSQF4HTyt8K9uFO452KY64JQ18CRipDAyGbdUKm0zfe
dfaoFH/K0CWeDMZZdM1+fQVtOVe/C+R9xH356OPx65tT36kQu9pr59NYfQee+9jOnSdGModUw1x7
mqNT/1YMJvo4QIznvlSYKzKcf5aO0k+BO1TJYQBxKg1MPIJ6gHB7GYl5OhL3MN8+IMIXGeY5peyo
q3UAdvyb8Jh8OCdlDXv9mj1kooXu5StgXCFp/C1zLKM5pfVSlPWTNQDyR60nBkcSwiiWCeBGGAx8
6q4y0YCQkXXihTyinNNNRiUVUyo00sDnq46hg+twQzOCZUvLoKje24ScXufufT8U5z2qheWRQsct
NzwFi2lP7uQ1WBk6wX9pnPNLwci9JGebsz/RMeTSkTF9vtMMlyOAtIXGic9oZJr/iR+ouCaXIF00
18vjxipy/kmspOAYhVZdj5sQhAHaF7FCWyHaKy/al6u8u8CdO0V/2Hh8zjbK8zpS15t/HUGCwb8G
lEQmBgRH4qwbJ20EiP7xctTAo2cTOhlqr7yzF/JDZLhwx+vFHdsirL7pXaRt0cReelMgIH5jrBAk
DwD09Nmei5e4mz8XFNqaqk6Tr/IDzyXlT/6SCdVoYchDaGflfeuD/nnh9wRJMuhD1QSekiYuFITO
bUXzQbTil/JG+yPL5Pz+acl0GcIPSlVtsa7UqNziH8Wr9gem/Avu5AiRBzB5EP4HIu3lXm8CTv6s
8BqklphwOX+4MfhLLtRhwP/q73LDsU1zjmjdnRlmQ5fDIGGPz0bZ40fNhVXF0D3V3QRMtrOljkdD
4987e7iSIgnD30oO9bivDJaXOtBzsmpAu7bXxanS1URDyq6zDyLkbmUPsy4weM33nQjx0FZ5e3N5
XwdysgC/aIQaT4W9QfrzfHJVlaf3wtqdPZ02VtRDF05jEI53eTvg5FNvsIayqIXpf0L9yxv2Rio7
F3TsmToQRjYV7h17gwtzYUq6eRGqKKDDRxqh1lxoUURmoEAwfw2zkCEB3NiogP7di/wTVDdA2Cpb
JTiNBu5IzzwlDlQOOR8DbRtY7xrlQ1IVeBFBpsbQXj9kJewMM8WcOtmd95ytpV9ce6VruJSyo8Az
01ls1HCtbopebiOYyHxEFM6Dxtb0V46jnP8gT3IW9CoJfwT0ctKJkdy4/cgcd1FJU6e/xF1CO592
YUv5dwpjkF9TyeM7PKvEwmu40vlBq2uQ/5HwHobgGh84yVZ7fD69QBGrto9PK/Se07wPoRYLi6Ol
fHMKLNP4TGMsPoC5A/hgbC9N+JcADTHHfcHMFs0FLrZXp6I4vpEIBF7mR42/9GZfW1SBBAYA4Hqz
CuByEyv7D2GanOnDF8HBzWpoWiWfDgG3N955MhZTsCnaLbGZIZSU8egn9dGhlHetbGGKpFDOguU4
Z/W2wJAdpZ/K1jmWydhpNcq3reJAVxSb8819zQM8p9vs+XjswBQZcitTPxfY/nUXCwEEUmDXRiQs
S9xNwNi6bt1G+GybN9KIwPCz26t5t5xJ9Nd8AeIGgZKBpOhkwi38WBQ1Wdpdpq1O6/lZVYxv0Zpl
rjO/mQ7DEaWlJ7fbln+zP4RoTZso9vEOE6K4QOzXV3DDxJ1IQSfaV4W7noF21AQvfFYlXYXi00ul
+RMILr4qECACdEo1QGigyELBywUxnksTqVrUQnQTh/n3W9vzG4KDGsJbF8p+IoahvdAw+j6UvqQu
rwrg3U2RJb6lTFhATUSJl8IGuU/aofCvDEJ30Fxri1+qQ84b7No0aUliWdq/FWZCmPr9GHKPZ+Fi
Sxk7V4YgtArhRVXro+exghHyHQcwd2yHPBMbbFFvN7PMPmdkGKNmNx3tMESZvahcbCazJXCFXY+X
ifjnyf5hj19z6pvmLZG7A7TeqP/V1FGk5uzpjHJHPGWpkzb7rbPEPVgzze4hx6jFqM2auzharHYt
FeBy4Xm2JQyQ/ksfkhkVTMId9K2xeqG0SuiLoTAFj8w9PCArcWP+R3ErCU3sY1j58N1rTO/fTqro
v6W4ot6SSkrVIBN8Bm+Prx0VnX/DJpWVUIJ9UKSj1sdnD2QWCRBrcde5hRUQNM8WG88zSdySvBSb
u/7F+DCqAdQL97z8IISlnMDmmyVYPG4AN/CgI6OcZqUXHZHJQhVHwkmZTQp+LcDWJe8HCgWNz8Kg
HRa6bcAxxiyjPXADvncUCJ7yigWsDCBBwzSQmK9p6IfpzL0ctgVXwGS0ctb4kiR6hfL0OavBARX4
h+fHrHkrd9aX+P+BW8Z9HEwdBVBKBMPfpnwdQM3vup7jJnGy3yQSP9kyHY4LMalCZSq7AXbxxDHz
/qhLRr6kwSFW7RuxkZOFkbYpVczHwaXhos6qelMVHL0P+ZmbTiLXRKCHWtNGgnQ8d1foJpBUCVZw
YtV8EqJtjXBUffQoMlYk0gsp4/Z8VHNyVjDzBxrz4esLw51+17NIGBVDRlPeubEG8pN7yNr9wusZ
OTlqCgEKXjYY7mrGoWBoNt+1p/tb2W+bACl354RTw/xnRfe29A3KjthY2uqPq4sZzRsFQBZIJhPT
W3nSD5mJBK4szFrIuZP1XoeHTfz0Ms5Bz23dwv84YwP4rojQAna89ODvAjOuHoth8PwZRMkcBKzF
2uw/jdPmQ8AasJmTG7IUrutXvZHc06Ho2PHkyxzdsf3PNuYeMkPisLxTd3gWVLZz3rk2jHUVvYYs
HbdVToRmeip6TYx0ykQR6AWGKk8NWsfSsG6AiPrhJXzdwsiReg2WjletJrr548KPFSkvtsNWSk5T
Cf99U06FcW1hjUi5cSdYK1LwCHbZopVP6PEpS9Bi67s8TUjkUBHJa9FlznWVV7cGv2eRUANysrsC
zQYueYFyYYufLuFOqoPzK/IyLCzJSyh+gVruYQUd6cTwVkfdixOq6aMtWmLnkF/eYDeQTUqw/bk9
J8cvpqbaHqXyliXsPiAYS4ro4CdaCSlYdV0+8EsinJonNCxUbz71b5Foo+jK/TCmnGr8VzocO3sZ
2nbEX7qsH2AAMsvaCcse5DO8lzluhkOu6nezC9tt1jGZXMkkiNuTcVNUA8qdm/UE5EFcWt+K5kxK
d05anwaOCkqrGS7iBN3VlF27AwGSJim4AoWgXWjFnqoh5Im3Kc9SkStVONbniCorkvsgN8UI1jKB
oqMkH9HJNViE+gtQhLFv4zHL+ESeeayNqdhijZM+4ow20VVscJ8q0BdgTrOpm8VxejZrU2kmOis/
Mr5T5Sfj2uuZrbJyJUWKIiCcbVssTusi1EaXWkL7R7tDFm82R13V6ZTh4KrarwVyj6LH/eABKDgM
fUKf9lronz/CuyZOk1Bd70jmtuibBSK2+CNrWBG8Iy15rnmQUt22XiDzL6o9pmbUySXi0UsjYtQD
sDQNcyaTsBqUOIlh98T7YookhnsCbQrXW4fz4njaGzAutvzthlvqu3luXpcRA1yo1kiOw6sbtk1H
/pdNS8E4EMSLhS3Ezd3ttfLnuMOxyfFp2X6U/2DeocCWlALDtRAmVXySo61+JUlbp86XRI9vXyaT
V3d4kvAbrcNKQOW8CPkt+HJFfJxPuoit9H6ZAy7sXdAMD2hUQp/NiLeYbQTa34xtuu4mvU8CuxO6
JitwklLnFAl3OiW8OombcLXycxSUNtyYW3Y5vGmwMyWCwUx5ygCibCNT7w906gV8IjPUhWcWJExg
8DeKWw8DjFfVoM8ldAJ/IaV4SuDGRbAdCt0f0r6mTxA7VI0Mh1OFtimjDptVjoP51/kH7JeWGL3D
G1J6pjUkKXSFCflmDOghJARbxhtkqt9v5txP4+TE5dB+e2lyPa+4fz7CFBYaHR01/IMXjuvDAXBZ
hkzkfA+9jZbvJPLm08+LNPrm2SvSkhH58FNkvhiQ3ZB929yS7oOsgemqQDf4L4AnjWnM3MAa0qXE
yuq1l9+UKfN58hiNWNpFQWZzImhGZSDA0JaPJOM3Ixi6rXc/JXT7HiiMF+g7Ps21EfiBKDPcBYfD
BMvuYLB0uysnKj8HMp+Hy46F2TRutMipYn0RzL6+zw9mTFmlxVIm2lexfWrN98y/F4MtyulanCvE
yseVniKLhRwgUmRPQF0xSjFyA2+dqQVhbeIId2INu8TK9ebnH2sPq7RN0aXlgTsEn8qiUJwBwvMa
cvosVoTglvrAdB3FC9mQtjhYBUwJutjFihCxYs0KQiM5xtY86+srdXcONwk350259sdxXdyss+F3
YKSL+fq2u7nmxUrMUtOVqfzVwH3ElSgxgjw10ejVr8XOgALZ+AVazdzcXVf8X7Rl5AxMnsdGaPVA
VeeN6mmLfBKe51f2ucVcVlHAz8nz0j238bQpfign9oDemTJO8Y1qC/TnKnLQWQpxT5TmqizTRQGd
qfTzBlEAJsbinr2ZZ0ObtvTVSZK4p8lgZaTm3eRu7o0nn8DhZy5gbk91zJErxJ1h/80tUbceI12g
6fDAGIuPYJ4Knd1JOdj0WBpO3N8qnlkg9x84TTC2LSWvVTsfOO2RycFkoNhlSOzOENrNfYahrV7w
jSRwUxtc63Wis32LNfSsrWp02bOKewWqXFybA/XjN468c5xGhNGyKZW6zbZvYHyzXoYMgokM7ll7
d6pjFf1Si8510HQPL0npe/D+Yka1QMMehuQ+n1n23G3ZaNNkLpYmbgn1QbnUJFIdY5sALRBnKq55
mLoBPiiD7HCMP/i3UjxVe9nNRfhBg/wKXg832aSsYqtk7Zd9bszbSZkEbkr+vRzLYxZSw8oXWNcq
jjxL/7i6g6OnNAcnABV2amjYFZtJ+8nrsa+clXs1VJym6w8LD+0hNtimgxRV3+AGO5ZvO+YexwQR
reMMT1YH0xsd9yqiPoafjVknO9104RjxUQOizoCixGEoieMCqZS/GQiUbkVTJnS8qOmpP2lBTDIe
6cMV8FiyKoVKb6w5JPvhl45SorezZRJHNYFMHN8lhwswBL9lU+I6Tm/pM27AmJ0I4zI+BcaQ8UdI
H7xnc1Z0GRYvPGSFrzWU0zOQcih4iWPKbe7daD5+Vw0UxrClyr5r7J1mmik2ynhpldfHJGCsdGzA
F2FKGbv4DZOnOIT/MXLElS71eAn7PDrTyvVFfOVYAxUwJrX1X+Yh+Mo816KmzYNPuFAhvyf33fjz
5Fp7d7DBP+/UM9peDz0dmsj+KG69wbjEp65fwmCFggosoyN/6DGjydz48qd5MCoQiiOV/SHpmz7u
inNSO8qhmFRJH3lT37j0ZqWUBxYQqYTK6MRaUcFEZ11EqUD7izIOD3orTwz/0CYPrxPXARRtYHzA
/k8+lDlsSHX7ZWRac9y1ZmrnMU0SVm7vb6w2crHEdU1Frq4iOccxaf3W4iQ7zJKrOfNJ7CaMq5dg
63auvJoX4C0Oeq1kVTzSVBPPgeRAC6RLgoDP4mjkXhO+svPQkfdjGvRW50pOBySLCEgGjX5l6KsG
Z+albiVwSTDAPhevHeVHPJbNdHKC2e/aw+6K2e0hLSlnejlcnLm+C449OsHWtSCp8PfwpHwiHzLR
U8yj1bnlmEXPd1Ts+W7HLNZ5TXj13nFzGEKc8RSch7DQhXx6k7kDfU1ZiMwMuB3LEXqG7504SLEc
/dSvqlWXuTiH+AZL9QArvczkX/y+OimGP65X7zAJmiOZG3CdTZxNbrQ4NpNNLM9yFZAPKRcbDatO
dXSTKMBlemKzTxoyKAtVoyPBdEUjh+XNWQH7hKHC1ra8oQKxsdquLajsup0kZs3GdFgKbF7qA1UH
prNmlnhYl0rhzvfmmKLZgawXWLE9q05iI6FjEu4TtdKlRGHU/0V0ROPzhQPTrzpsx7fZLeTv+2vb
maJR6sp9FHdrMwr9YdpD6TuSfnlHlan1hqOzKUkof8wMNykcpJK6IChJ9/1EgDPLq8kSmWc8B4uy
hKQdKuS6UbkX/EFn9EVQGVXacQy6N13DH1B0Vi2BB8DKtqKnaIT2LfnRg4orEW1JUe7ccDpzusow
2W7R6UVAaObRLai5iLav/LfJggrZVacKrFHaBCWQTPTX6+/wWdRQrycP7DgVxIsPKVyIJyuoo1p/
CwS/7Gj4ki2EjwXdwZ3BUwev7UjI6JurkGCFKX4J8XsCMAsPRst2UYR0xDQVPxl3JTucgmRQUc//
CfUAf9ZgochuzChRVkj7d3pLxJN4fBBZ/V7PjUjb6UAZ1MC2vie9FJPx3EjbIlygQqd5WDAOTobs
ZslpfvBMHbqanLf7cpCFkwmhzUQjRXZd+8UbiMA30T1dyHtts3lK3tsiqJ5PBLfLrkYicCPuEtGd
kudtWrW6V1Hr5ankPJpGS72vMj91nZ+eY0owvbAa1EYqqJfEKQMORpCTYXM61ABr/5Aq03EUScdl
nmArGxYptYh+6TNtJEWWU+d6DzhDYPPKgssFfQDzEb/ejZPn/Wqs6I7QQA1qmE2kFxRgnwfh9mNX
BTM5Xb0PHQ+eyjU0TtsK8qnBncl4YsB7ZU4NhodUHBgrABVNtd4m9ry7/9L6oZPYiyTve7ibmfrW
uDGmyonCqYERyuYWPfS5/faTa3mpXqM3rgJBd0O1+rm8+7MzMSMHwITfdsZvz9SO3QxYP2+m4Arr
vlxP9ch6LvoWVVT2Z12bUnImmT65dtgh3onb5ona8+5kWhkKaobZdL5plCJPIro4dsL86EzUtVne
PDWV6OutjR0mIe0zm4CFizUttutaQo5hxmo0djPbCjmDsdU+/93JtxH2sK06ub65FtNMK4Zmc1vu
4/jWxh+LXfbHoT3IMGDA9Rv278nns4xxpnMNKf8bQ7YALUFDLDIpihmpe0ygmDyfJ9XTEmg/EoI5
A4FsHc3FOsrcwtPL1qX5OsQieMwT7ESBoaZEXsv7xmc+zkm6uCCxaj9OumnQo4Cz3/kSDOeB1Sav
fBPETo2FWC3MYzi0G1R9JQFSBrJHKLoHlEhb3NVQp9xSEKyDOjO05Osf078zTJzK3HPbompiXvXD
V7WJGItFdxLGcjcJ4FgL2YQ/hWs7flnZiEvTVSugzdTc+6+G6d7/dmZCjoU0727HNlHXdNgMS6P+
p8d/vOVpo/2V1RXIM0qSfnUoCziJnaJjHYlzyjjauSCXuarPCgyHm77bc+U9xFHDzqH3HXsuAT4Z
G9R5vrHV+NXE9DAArvaub/e4wawDBPsS4xXpxIHY5agIA32oCKBO6fv33lvxQshu3olYKb5o0rX3
FxpykZlWttMK/ERk/HN/2QUR9L0+Qorx9e9VHtMBvNc8gPthANAUw59DZGdY8HoPbNWt3RiES6VN
B+hgGE1479YZS1xjbguss8W5CEAn2P4nLSyVRBTi3Goz4kZX/R79H9t6Qs9uju9drxfqqHTQbB+i
VeiFWGaQYNCJz9MYsfiJCdh+91Ggpa+Id6Iel1TOoQbr+iWi2rfahX05TKL+g11K57P+UsUkTfFX
1BdE1sgcezpmi9yl0okVtFYV5DT351aeihE8hPknSAC5p7xC8N28xXKxhhYgF+BVxxMAGR1mBh+Q
ICOXooXGxXMyw2nehQZ2yrVRw6GUUuSVKGDxl78PoGvtRBJ80MB5BWW66JNx/blSb9wg8ayXvS4U
QZCi6nFC2D2JqZJXhSe/V6GIRrHBH2AQoPdSVOCDgbUm9WBtZBShT5FoDCfhc6VnQsldnTkOmYsv
+mFxxpcaNURn4mw8fKeib9vY+Mwrqim39LWoVdfG/EMSnFVnqEx1eujwdvhfuQ1ibDkJ2O8YJwO8
L7uOD+AlkDBXykY7eHo9On+0G8Fp5YXTtEqc3dOcrs5RDO7AOne2RKYk4fMJq2G8ncKMMwC/4Kak
HTJ0IWoZ+ahPsGvgAoI9qNjPH9er+hm8qLD9doyYQpjhxpAf9cWw/UVez84bEU9iC79YVlfOnfiT
zS1dJ0XWeolF3fjk2LMaO4w4IdhPE+G92LVDNT1Q9QCvnnFpGMY0Nr46uc1+s4hPn8MaN0EJU4Xe
eP2idwr2FoFjOlvBVSLB4gRo6Laf9PzHbpFMH0gry9CegaxppHHXXdv2YSIilAHmzdOg3W7MMB/D
WeZ6ddygNRoOkKZdELUWGccAK6mvhYLja/By2J/UFL1InriKBqnCXaRETb7n2qZMFduwHuLBFEBa
yk2H58ZAjVPOc6a7EACQbDuM76fwBIDUwiJYs631lzqHAJveoZe54LheReyR1eri3BtUAqJnzkXu
OpbLq+1xokYZKqwifLRfvpKFA5njgHWadasV9wgELjDdcy0Y3MfNKxoP9/m0pmEPS1kgC129G618
fGocQhRNqkxrdgsTh9G7x7Wub08yAcm3F+r1TmOdSY3iM1hzQIOKom95NRydikq3clewyNndLLf0
NW0nbPDCzu6eEPbbA++hiSQ8vBkIjlnHFTmDGXGDIKvOOvSaTLRhTie2MGkRz6i2jB1cYs28iT8Y
2Abdx3zP/Yio1VdKNk2BRZgskd2vpYkIUd/i91M3IRgwPKaYUkksfagEaDI2Ucml64wXigIdKB4+
xEa+tcai8nnYXrshDAhZb8YFun0riUMu2nblSMHfIJJiSdOmNvHA2frfmF0hex663S6Pm39GIqm9
u+lIm3O5cHXioB7XU22iP6OPmF0PocH5LZe+imgyAv92GkFUCHYm+Ku6U3qsiuI0KDTA1Jbg3qIK
xJi5JKInJI17oYfSqEXnN9gSfprhfmwccGA16ONgWvQumMEE0IroRpgy0dyo3RC4OxPM4dIBGRWm
GF5DRLxyPcS8LRY1qnBnPonCRJskF+Srd9oySqnFRzYN6cEGcE56RZWWryezF/bYP9HDxwSwXTqM
vfITuZB9B0FcEyY5YVDK204mTf2/qubQj7eyn2r3/tmJ2oMykAiOikg+3UdV+f463dbWjW7Q/haj
nUsULPFDF9Z7ZcPAv+iERBERD7p43BUDB2ih53L8fHn0PwJ2nGnO4pvHrqvnv1Y8WJcnrYWVVWv2
5DqXdPrhaYuctYuMwTKV1pvudU+B+hNh8BGzrv2S0ZnRq2t9rBbxGgOL+sAMgyq6Hlcq+6+uVXS2
t2lcoLHexGbryrJoP/A8XZrhkJJbIgErzpCrt3ZpshzIff0/yYF6Ntahy7r2R7rv81lL/e2BDu9P
FaDYywbCJ6Fw+m11QKFAHyDFmrvQpD9Q+utO8cFZ9Tht4m7jMaiRfX9fOtdal/heFYV9oMkiVDPR
Qy79dv4j2ZkHBkqvi5q86SgcKDQfGh3XEy8OiRNgYqCyoqN1bm3rWNArhw2HX8sC4OkeFjJRH+bw
0mvg1LczoBWyaUNi0f0qE15GPNop4ERF30a3C44Sb1Gr6pwstyZsmCebTuU0QugnET6mWC4ivVkH
lea72HmrO/X4mVNjyczwdNNcDt0xM42f4EynHQD8YpNt+YXxDWbutEP/L0qJ3ztcNinnxrkKWZQo
r8FXciLWJeQBl6o6Q9RlwcgRDi/Hbq6v61MFNhrASoLKUtEeXnYMnPR+HX+7V6Cn++2nSEKMjynv
b724WwrvY6z8EDIy03bHPTHEc+1bz2X6pHw3/HToq1nEmKISzESTF1H6QzKa6WgIi9kV8PfOWNZS
Rod0XTxO7IgN4vu9BO2J4s3786NTNBatzr9DFOiJ818RFnqnhO1MXabVzlbI8+6By6UacApk7XrF
Uvt3gxj+YtDxziVONF+jf6zDGmngYVkSXcF0/CKYYmk8Ci+qz6z+d5r0z+7rFjJB+uk2y7duCEL8
vY3kefM9Fhil//ZTpW6ZtzSC+EeFR39d2q1kY9UteuMhXFcW/UYrlik/AkaBb3Y2NBzM2nEWfWqa
VTLNx+yV8q5ZIBNHqA1omC2e7tMFi7/J8jKZzpw5o3JTmcrb5AW1hsrzobmV/8p2rPY3EehC3eVu
Qzb7zHI7R6GHIkktDg4yxrwoCQ7TC8Vv2dHWf7EJLhpBXq664Dl4Ih/QSM/qCdrxF0jx2QKStGrj
Qym07hOAkiQ9EQd2q1RwiiWLKQ3DHzya1Z8n4lvQtBR478hGSQupXfdI9sWlA8+T3wM6E454hA2q
yX+cUeOg04/EhrQanV/SFrEL6STcGzJF/YgpGEVBHQ9cC+AnV4y5tSMELfX3ZzfHhT4z7iUK6qYY
UaTAfedh7wTHc/WaDlrWr0qM2Lese0dHCbUy7005DcQI7K245wZw6HhRc+rQ+UmSrB8k/XOnghYE
wtX+l844jDIh1Io9En6bGPnoQmIsSQFzK73EiChpIILx4+Ime3DMXqnQNfSZDt75LYqh/Uxp5dV9
u33tmJ13imrHvwpF7Xc1x6Wdapr7x1+7bnMHWUl8mf6su/HSXLK3b6ydgCxjwGnZCQ6sOzMHGV05
J5XznFqG8ZTo3GadpOSwV5ez2RyYNOZTElzd9WSZAH55x1EWvoZugz33dntNaAJ0ebBcaKzKO7rH
rPi/dVFFFug7yQWSSnRqwoHGddXlcMUJAhzRYR4b452GxUqbZTZ/dVaLxvAWperY/3pDwwACLSVP
snWnGpjHHKp3i3l5f8IXj52Tq+9kdtc2Qg8Do+y3j/Nj7Z/cxmA25t+1Fisp11ldJn2Gl9OKxQRv
LDtdf8K7Jsq12shRZujPAbzD9VfbC8JCdZSXiVUjGxdshDOV3hEANw/u2n8VekJuWDVpCIwOb4+L
VqIxB1LJNfcqL3aLD3N+Soanf/b0onJCTsdQov2AZgg4HoU0fBf+nUaDQEYmxoD6OHeKBxvDe1bQ
4Zngf8VKxgOglAFCZF07AGp9KPzSUIryrTgwwDcCtyk6jIrMeXIfLSAoDS7KCCkkpkL38t+jxPKg
X+0yWHiNuq9YobEAb4vFmi1R24rrW4E4tz4HRImZx9KBp80SGWqG+P7RsdpAZquiRxkul8P5GP+W
lvbKl9324PqqI5VNq9tXoa+CN5Pqjo4sUH8tIzkAUr7227TtXz6Zn2W6eYSuuuzfsyEl/5twVLna
PSIUNjXL33Ds0LW+yV4/uQY9p4RnhVlen13hiF4Qh7sBndo82XRybF7lUmPWlBi1yfgeZ6uDo6kx
W4B3uMBCt00HnQcCiXINgm9GdyvruIi5AnppxiQ1zNbES3/dGY7WVW1r9pcOAr95SW0Om431A441
d9amht9AKT+R4Y7h3ebcElucHU4tgg1NqZeVCidr5uiiWAZJYoXaLXu7Q/5BEA/prRte/jpuCgdY
XuMcQ/gCC5mY1oUg43NdofgMpZhTZj2LHMl84sTXPhB7wicKDnExWcQUys3HsmJ+Xq1JBYHfH4og
Bf/XeWddsScpK4f/sL/yVM0K38Yq0JstS1Vj1NP4hdxmUm6ENcI8bQ9gXs72tT/mm+hhiwx5DGZg
HigvwSnCbXqFRfaSPIRixfAANNsYtmfbtS1FfIpQfXXANme7yAFQAznXKF7KgxdqcUloIu3Qcukv
z9O2g54a05sbh65oUPr+1IdWh0MT86OWVXGi/LV/DXDEvAGG/g12qC69Onh5E2s1XJDLNwcvcIrw
B8yPnXta0RRoAANZleCs/AWVgk58UhwAKoUz2z+cJs0GSeL/v/GmqK+pt5+Am2UaIbpy3eJ7x9Ya
dk0AMwECN3VgifCbqZyZmw24x9mS6W5yQOGJcIZB/mRLm/XrKPDCVNr6YetWRFcu6amaq0cxpfOw
wU0nbZBvtaK6rQvJP14v25eY0BtLXrbg55F8WVgbUU+5wqtdXjtCJLyghVHij1g/fUvR9uBPPAue
6iBh5zSUTnSbqDmMoRIsY0ytn8ytCq/m/5p1SzTRtrvI2CDb5llcUVBX3xvXOhPhGsuiUCwNunVk
qnLxeAhwGmafcKLrwiA5gZY5TNJiztfzz4tEexrtaR8cEH6DYJKlj7cR7qH0kaNS67qrEYxPZXJQ
uVes3dr094VLsintSo06nexTnmVidYZsR2XLku9I4F4l8OgDsZJlzah5dss+Gr6JC8Ntd/GE7xR1
/mFmIsjqN64DBCkxQkzWHNXyLiQ2DQjF9nDf8YiWpOqEO7/JsD2qYdqADUwiaIdX+vFUnI4bQY6K
6xeq050mr6cBv+laMKw3cy1fbe3W9TH0SFurdXL8tX1M4jKJ/9BwJQFlFLdh8eofD44cjZA7WID1
NZEbq7jUv49mEq7NFxds/OXlsjszadPOrVXQF8jcNn/oxlx1BSslFjdaWMVH/Z3ILygXsHslWAX8
agNbzCDzD+O+lSLLeYnyCxSkV34Edwry5+MLSVzDSaep+2mcpFkpL00xvhKPm3f5rCW/FZ7/sEBV
ZDMD8CbxmK46VuITd655yV9eKioOavmV65zgVxtetVtzoUTH1p+MoSpgQPyLMtSN1nFq9qsI3MSr
2SNI2LQYASyWVOphnLyEv2S4cPRyqt72tgwpFaiNhPxONnseQtlr4jancK/VA2STqIrH81iw2tto
R58Qg0YqrIHniCw7VJ7+FDiUQsZDXtjlD5B/tvTcWR1vBoYVWTCKLwgcVXhsYKKq0qqe4gmbiwFz
+Hqo9Eiec29RbkZvDJxcUPsvteD5Au3py5myUGWVzf0zE1icusIJ5SAOd6K5zPFlgK0nCs+TkJEh
mwQL8v12bXnAoz9lDDXk1EUDpM12wP4t2O/yvmA3HlR4LTkYTjxh8senkP0nrfxMaNxvkOKkRbXA
kJcHicVR92gKEiw2Koz90Yim31al/34aVFSMlLXXVyZ/sR0KVQYXuylmqrbzRRbG5MqQc9T5guf5
0zD8HfV9OjhZyRgq+KsdvYaxhBfOskEkh34hfAqqZTN/JG590E91V5h9jDi72f3su4IqcYw3qkYl
DJ7r1s6DGHuYSv7HEa+Rze5eIooX0f4BmyR7y/Q2nIaLcaZfV6XruTTEcfg605c1N5+2u3CxfCnp
ppp1xVoOxNafVoWdaNUk/1z1FZzOtDOWVqmWyoWE2mA2uauRC3mJa8jV7o95DTJZLBI+sVo5Po6y
hnSD4PcfuD3zOW7hRu11gq4WzAu/LspaQBcPuGQJZwp5f4NhhWOUlJhpidlDmmzl9NN0TOLPLB1T
BhPCQglHf/MWL2aSWM+Anz9yvPt0f05ss/qCk/BpakTMVl9eWw3vjCThCgDU1Bcoijq1KvvTf+Xp
EJF5HW+UdTlxmFIvX2pSgNE+Rto0LHs0df+0kbWJs942GYi0u6lNPKDrDKc1nPCwvDr/xUlWmLLB
XbatXGSnM3KEzA3HJxwq+a/r+8Ukgt5FQJXZUVZXWx3/eyH4q+dtIwMM1lytrAP2IcWeeg6XeRSj
GX0zE8yPt8FN5NhE52fUVqmaXCBdO/M2r/gUs+Muup8BEqQCVCYy1PhY7S54+rA1JrcWEUdGwYmX
Hs9u6QHyXb1VTB8AaR5+ZB3Tn6E3ZbXKI6/4CbgIEIwPoZAo6IS1B7B2OmTrWCxncs8ceMVWhSMC
yxf0U5nLvFntUKOvLL9DMoBtaIHTcEEk6Jv7m222V4NHCKdT6N4L4HTlyX9zDjwOldeTT0R8OYJ0
CqWKtWhNONxQ18uSMrtWwcZTZLbWszCjqy0o7H8zs2UASBs2NeCbnMY4FS4q++q66SklEuJi7bgk
us5hLdDiMSu/o3gLfLA/TfjEqIUSkXF4mpcUHeDPn2LkCZmNSociSZZzseoa7Dlu11x9PqGznsq3
oVHpZRmkl6ANBUo7OfadOg5+SSspgox+HZ98kZNHA+KYb0Ab+hYeSfst02HSciF/AHERAAa+kvqM
K13yVGMFdtysw9DjK0e5cCMbUAc1XfzUdYPAM4kxN5jck2KSxJD59LKxt4SnLCGY+9sIfGGR5AXY
FJ4nF2UoO+7DRezyhFUuCQL+3hS8oVKd6SwZH2NVRvotlLZDxt0KIJOe06Eb7vORXGRkJfzg7+YP
Y9kvGKyY1oVE98CP+Ps7RYdCBZek91r9cKhwjz6IEp2+tZwHdPkivbWhvXhGsir/uxp/V/7nqQfK
hHkyYny5t+UxCOToEZJc7TooBjEwZ44u9YN2fwhKGqq0BfQjvELZkg4nUtjZCGrMqAKa+piFiZBC
mUaTrPFWd31pYmbvoY4olUUS6ykc9fbJjn731zWFJORIrn3jzgcMcjmgmEGPkMaWllzuPjmCqUat
ApDicFbXWSLNfyF2vVnCUCJrZYgTgwlAnRwlYNAYF2nTVDgqha0yvknG0fdmTqEdhYQ5VS8BI0iH
pSH1EWnbhp/8H6wIynuq5mV3IJN5UiXc8r3ZpQVr4HCMEBxb6aPU5D1DhZXw+c1wz73JVzVBrH7v
/o6puqjSfZUsIGzfqNkZBlC1RFj4bxgS8Ey45xm1ULoQcMTW6oAi1ati1EfIi8q+7VDTNNYIN7RX
vRaK2HSpym9L2qNEVYFPNG7RBhUeMsDah/Iu2/Iz8dtSnrwi0WzISU4bTAUc5hmJLJcsE7gzFBuz
oTAI1k2kZ1SZtUA1Q0plUdOp4QPbfUeOaGZg8SN/CHXNRf1FOrC5Bsdnt6BAR3Rt1NlmdI5iCROg
AOOQ8hEg3U/0t2a0sE1n3MHqybaVhk3tkE4gfLKNylVQuE2Sbn+uxSXpuYpJkm5Ws491WFFpvS5R
zs3w1N8IjMxZBk8vo9EhqdCalI7Sp/UB1OpN6tLJq6jc+IE9hMfd7Gvbi9S3R+DRFg7MeN+w9kw/
a2Mufb38U2HqNQtTFGugDSJcFGetmZOu3Ao5hhxZsVGB4RhQNrUQ3LHXoWyc8H3DzdPYfQUmmUPX
KlvJMAaXKdK3ehnG/j2kvWqg3slvvEj/RFOeoQSBsayyHuf39Sx3DBJw3xh3EXZN7Qr5VBsZhrnu
I4ysraRt+1uexGXaDYm7Lfd+8y1I+EU4MCJo7Z8K0nbUUOXpdnjW2Vha++1LnhDkr+Ox3BNjWczY
2DMr0ClQBb3iEk81xfFleqWarrnvKsFqWBXgItUXXX5AcT2j9NnP3TImevOtSR+wC4yOqvqDGaQ/
J2MFAWlLTk1z/CWc4jMjG02UVLhi55iuZr3HDD5tUEJBtWX9WeiTRMGa0Op28JY3km9ZvCObzqN0
7puVmpwytxUW7xLujBd6ZbT8jjoiV5gyl2LFfi8vYRhpNhJdCWG+WDWb5EhZm3BBa4+wWEqIWLha
nqkeU9PTnAh2Q6rWQWmQ8thabV4gRbbcwZxNRxUHJzchn3G1ta+5AA/XEzXtwUHeLXs4/O4G4XFP
MC7wItRC5QX6HVPRKeunWoCQf5pMHwHtxOQqzKXbexFa+dIxURv2gycQm6FK4i6842LPJcjjcTak
33rfOzPTRxbnwLiZGWRJwMwSPxr2los+4KxCXc4GG8UbdBGxMZxXlIgqkPdaLTuHic2hVCJMi3bz
16c4ZlAUDUhRfdFHSs5esDTKRhWQqYWgkEEbDWBTul1kN3D4pDfSWiXMkhb6O9KXYSRvMAL3kXnZ
+SUcovaKSyonCnor10vddMRqJ8015x3UYZQTMPMz9JMN1tCILz/RxDGNFnNXt5G4hA1N0+4q2aG9
7Rxi4QA1Ys3ULdHAjbIaf+t50uw07hlIB9X1+b7rOtfKj7A8QhkSo5x8PiJ1lgzutnKJ6VkzH4CR
1saNsYVL6AqQ/JFiT7n1pMgTs+34UYwzYzEy1LtyXTLT/rmWcUDxqaiD5bDUgwc1N5n/MB1kTzJb
Uxt6rJj4+yCzGqS7JL1Kr4CcRxJ4SPdX3xEeJBdsL1v7r2N2WtncD9n+cTbXbLtaxK1dedk5lobe
TIGz2MwTmQVRYDQvudIq4FDNweGFocAD9vayvmWfrQevBB1mvrhlJk7l92/7vgitAhOWBJvSpYSP
TEYqD2zVVZY9fO0Z2gcHoOASQYEQjjvWG55u70S5en/G6wmDSS5ypcZ93qoMGiaAeBssI57KcVSq
lhoXkhbeyxr8BsSBF2jPuRB4Wl2htuGssKa6OmjaDBFoPMVCpIVXiwPa0O1qWwQ9RDBWTVUdTv7T
dVS+iYs/vJoK6rseA1p4NQMRmXWyWGxwhD9NufQSvWTnb06yymljy6yIIiJX2d75veRxTwV9kKuZ
CaT351OE9ojJ/0j08kTS6lwgeKFi53w3Frvmr/7Ck/z6//0YTGhgqM3ibjXFAh0tqO9FrWdGh7/b
ZiT+kJ6NxwbzT1fEYNErk/QCyYLV8LRVnrkXyYXFVa09TJePIm7VWM0wxahCjaY+d1wheaMTi5U8
Yf6RsY62HVlm81oJd3KKWE8iYEoAJroS8kH5o1vb3IWMvw2HIe1KO4PTNJCsxHPGPSzNJzuqgCEZ
SXqwAGEib3VVPwgx3RXXSETyhSOEkjszt2cvnc7xnjQo8croF24up9AbqnIZrZx42n9+nrIZ+Mkz
NS0Kh2tjmmlfpItwQ+/NqFIPudg4hrzpMpbBZYy0B75oQCpvYAbfG2jh2WKqLvmbg9Q+4zPB5dYa
2wBv9uTG1AjIkC7YEPkW0srhyvmFeYiqI7jdTg7cpZlI7BP0Xq+uYGeVPt2l/YNbntd8iPcYtf2s
Pk1zaV3POpgeC2fo2zBiQp6w9HZ185znADpkywAv8tZLl8QRtV5bBe3xcoWOKpzW8pNNzGDQNrNW
/p6jaTlHfpvel1+8K/1WqYWyDcYJRsGrjspiQa9u5CDHPE+0lyaWQ0WLLYDXNbmOqrbD37hUEJ/9
WDRHmPAiwLVwF1oos//DT8Bs34M20jt/wDN5UUmAhXHOaBYmwbve6f8lK5/2lgxk/gbKNbDdPGI5
U7zs88jAEUlu9091SdrO1lLykeJGih8zuXapkWum/Rk5PPPOJDA+mt4kCZlak+Kn4ydZqaITytmw
RCRRF2lal96u9MUq7wmxbAtrXMSycd+pak0NUUaUOthV1FetE7d8KXl4CtQlQblUrCfPe+oRwsLG
ZNlWlPkOJvWPxeF4dOwyY/70t5C20JFmMQbJKh8K3GsOKCIY9pbzrFLKYH3ld+7YycK3nJO5A4x1
92gJjNC1Mfi1toZ5iPazhEg+kGdto+etP9D47UsqGQkQ7RDHKMlD2BMbtlpSkb/Qo9azSmZ7aAHR
P5J3iqQt5iNc1brQ0+5QjxqublYONp6nzsWUUF8uRCjV6om+/wCw54RgAPvqnG4TB/IjGt1yhTyC
3SwfBF8SNG6/0/SOp3oQy0N1whMdZhnoCZtlTs8wRtg03x502tICVsfsy2jF17EFeAeek+KIVPPR
eZ7J+vHXoBK9y0bcxLdzLmYNxE79OuuDYujqywIqmU7mXz0jeu/PCs5qj0wLLaOiXTVzwUNpChBM
D+Zr5ACq/IpiDAVXm7v51rLT7ERUsyojtUDnxarPrQfW+JRUKROrviwCHQWPKi8Pe3ayfDu7vvaN
RBKE3yljq627PtPRS/7VjN9BrujmMNU5w3DkGtIVvA0CHwBwP4BArkGBaLVhfaapvSVa36DqcsXp
yTOpRt5uuHlr+8JMi2WeQQtRsJgNjCKOL91iJ2HhGcUmnIvScpW2h6eotMw9GcX5dNWy62k8YHsP
a87FjKm5llNI9sgxHauL68XbOWL+GXlAgxiEfUu8Il0xVIfKajXILc7CTH6yMEfNG4ofZo5mPViF
Mt5FZcswTgGC0knCyMfJbIbXAA74mAJxeti9P0OVq4a4xjM2ME0xoJhi13hR3ldZRjzj5HGXY/Ol
g7REG6z+dD/u4l9D6pVLNTf3qkWRs3h57gbL0Ww5GguCMyaUhp1Rgeh2RnZDZY9JuFwT0cXkxNYX
KL/SHM7rmwPCSto25sqKxwsC3B7FtTcGGO+eDePZE4Ye/+SzxLsVJXphWR3TPZMyhaY1AU/k1EWG
M5bRH5JUpisSqd5Bie0DhBhbknu5adiHBH9HQhcUqeShnh2q2ONMkeBhzNED9WjZG+/TQ4ZzxI6P
XXyb79QPSHvhZbAqIwK9uRRvhoP/2aW6EuulfgDGqstVgxMUZMaRZEZkiT5tbdj+uy7Z6wpBWwNG
LQ7m/VKR2ghreFb3zyo5JPZMLmrH27DlGqq6Og1kZGqXTc3X32R7BEZbGTkSqBEse0Izkys7Ejg8
Zu9E4jSH+d64LRG8Z0ymOUux9XSeEFJh5pi6xpqSIPOlclkQUw/APhCbTd7yxaRtOE/JPb2eU4ct
93AJoHv9lxRpvJ+80SgSVPSnRSSkyIVKonObXyJS2hXN2UALd5PqELTwZh7/yYhbTjtDljThEogc
fGJiKEpcnbkjNvVAWWN/7fUo//fOW41CYjYTJ3iKRiPillSvEZV+XbSFhud9i5OTAJVnumMF6wlE
YqtqzsXYuOabIWr1Ot/EgpxuuwdMegiTBLys66SmyVM/bZ3SuRimWC3nRkTu72RenAT/nGT8RhzP
aDj8sY45usXHu1YDUEDbe6c8bQhfyLJK9M76TQSG3RORhKYssXWi2lQuhhIzjBZGlTK7OWHolcQj
PmpSn2Ksh3w1gBrEv9T8SJU7fJBEDiYWAieXBuV6Bt4S3asfFmNUXzKuBxFQKIaLNVPjeRqb+Aw6
F1b4Hmg5tim6KUtQaaDw03Tm7lwjkf1H9yM6Zs5nP52OMVqdm9unHTKPKaZFwcYEwaKnbQlZ1pli
G0b6Y662BCudzmTa07w8eOrQ0/DcTcyif08owfNAcT+4JmRx6vOw+EBt57J4MmrwA4PFRztyMWB/
IjXYbr8VSkd3rCXtpeuQvdaAI1C6/yWMfS5E4DZ37Ee8u72sym61GFQ8uaDl/9QRRr00jnW5nneY
vsBXQWBQGggM7i/lMvNLbIIfnGQCN/TWT/AcuJuGRfzGeUDDr4CPsEnMx9kJa0ILQAJvrZx/Jyhp
V7/blu5cXv/HwQO/g9RhlZkn9NvOeXqOSme7QeSkn2yvDEXkA1yq1KKHeSeREzuOSDC9GsmerB8+
+6hHBHoi9H8dgtvCx12uMliSK/TYX3AuQGrNPfbdqt2nbmdqmdmY0qpVtt3qPm7hnTQk+bdlsrRO
I80oMC4nVPA7tpfGUdeIGtuSAcpFxt5IeWiPJsUedXMuD65oAvucLgh0eSceV3mZ7sBwmOh2uGOc
zwkTLZtq13jWpE1pKZOnKf7ewWeirQ6zKhW7PZC/VM0QLQKic+5inQBEOUYYI+ZM7pYlL5w/IviB
3SKCmiFSy6jUfp35b1lf4YL+R3+4/fM/W4nIOmUjaEKqpOsw1J2edf2k8pynEfXgmy0Syvyr6nTP
qY0f2DnE0YuW4j9pUk5nLhn+8VO479uZ1HonwM8ln8tHdOkVTjt4QHoDEHV4E/2oIPbbqjqbZhLL
3LvAK99xqklATKeaAQg2qLqPZZ6jI7EuhhSdvuJyGM75Ew7aBLrI34FQo5Y9xoQ0NgJVhriQhZ7x
EImXrehoAeoUpASyE2ur5Cg4KEuJ+kkKp/OOxn60W0ylbqdHdnWdp4V5IPin7j/We3bYTOP2MZtP
qQPth8YAj6X9I0vtpeIiGwWGtSI+nS23dz9a/KsujVgruAOXvlzH0BnkOROS8ffEqMb4USbTHjuB
3nP3WtSVRuJEM/6QKbey1dioqCkr0prenewanSN53WRHtjpnoNV3RB6xk1zycIE22tLRzP7O9paM
hWxHeNDejXrYYU+wSlklHaX09+5m1gg6kgRGyPTEF3+MF5hMlLp5wFnWvv3uyKEBSrP5qpXwyLuk
4+KmlEfxjgpmrrWKvNCFMeyigOJZAAQFwkIHL3YFktHvDUvnthBPa/K4biYXFgaGljtXmBkDMgBT
VF1bRbCsxQgtQ/V03HEZ8YkuAYTUEzMHQRrYJpaS6asdydk/fihaM9X00cHMER4XeHL8HoMq7eUG
yrUQZTGUl1dFTEMBxUxDIDdixspuGaNeqwdMla+JftUYlq5og6MoEIh24CneiCZTzK+/Gvll0jBT
WR8kE8Fr2T+hCHtD6ota5pikWL55nsvmXUjG0iOEB9f7fHgum/NOZgMchfTtlVTaJY6Ut4Y+a+UM
S+lIX890enscj5/FcNSI3GQlDdjvuJJEOsKLGJ9ClyIzsZ5aVZAk2KQ7qGBM9Emztq1WmtWpmoMX
pJS3ahB9Nm1QTL6nqSvlrwUm2ayueQWAsQATCgjNhfwY42HG9IdFMYUOXfcSYNGlzawQXLi9DKqq
cpdHVv656Tr818e5CN858qXCxSuZSlJU7p+GP+ZX2H3DMIaRnbmHVfq8V9l6KFp1N8D8N5ZKlAgh
zi5lTROosCQJQ/XG5e6keIoBTbUNrukHbgBUX6I1d7u6MO97WwShJgORtxxMz/aJle9H3YH49lHC
5jssO5Zg7aZP1AueDCTzjslhan9RL4OIZh0a3WuyLyn5YlFNjEEPKPKXo1vedm4BIqpVOiNdq/H6
DXphI7RD5YcwkynDDDDAQ5yxhznHWsrqg5GAwt3eUQu/via0IsoECF+O7CfWPtxubD6AEEeAL9ow
0zDc/HkMDXcPSYZj7gOoEx50dJxVLuf7gvZc2FfOM6TT4nONI2bfNC/gGQSyg6F/XhLUCjW+woBy
q4ctuT/kX8nOw6/h82PCzam5hAczRCzUWb4sO4DWJL36EyrKGturihGI81ndw3Ip3hUSJhPoT59G
Ko8z8y1HGrnv5bt4rjkgtxrn+Ux4CoioZdCkl62/F9OmkQlePZqKICuzeNcvHD0d+zDQ5zabVq5K
Pk/nGqyeOiTQhSIojvuM7ez3aAGC/+NL3tiRyHr8Aw/W+ur8lw5ELJCAgMJ1+n0hdgsiR9ifgEIe
VAdWY/TItr9BMbaJu9Fv1WobrnytomURfPRZxBgjjKlq6aLkm3E1gbEZ+TikmMym0fhzILGEBfea
nQmWS203x+PaAG7E/AkXCweVt04sDQyL15funCIgYnyYHW9eREZ/B4DDRjfPK/LN2OzIpf/rqqEW
Lymv3o0X1eRb+LFhso4hjKJfH5pbUy3YQq/htgNXvpqXsD7KfIgLkxJpThQLEvodY4zs+qPGH/9+
G4yXz5h3nVy88jRFriCm7PcX+ezd0vKXii+DCRK1qzwI7+mgOziweCIr3fb65L/s3/VELXO6KAze
qrvKmvyGGg1NU6mK7WgiUwWz55fFKLjOjuE1c0qlRJMw3xRAxdSU6Kj41jS3/2EIqJNp59hW60yI
GUe6AKYda1br1lyBHzs87+npbt9HAsjb/Lw4/vXTrTO5Kc0WITLf+aVjQx8Riq5IOg1UMFZZBY8R
4sr6usnCyinTA7kgT9czHM+sYtcqdbEs5a8ofHPIisoH7/STW5DVG+AqU7dPJ5eBfoi5+2N7zKCi
X25NuewjMMHreh+MEHyM6MXlAEublXmZ5j3iALKbu3xDpIde5Qw2qTKiALoOgKFeAoJSqevYrsNJ
sULOe9rzH0a9PGsrhpESi/9RuWtkA/YyawJdilzv99az1dN/x5Hq747jVBK1YcAhekn28N7sHVBL
VSU0Faz4KSn9qtaZWRYSppDprmE292AjsgzCF0GK0Mm/y45J+OvKZtPKzWRfyZ1G7t5E/1gQUFO/
EwLDMk6tTLNsnZrcfH7eNhkAPLyHnocTCXTkpC0ZJHaavYSsCBDi+/5jmxdhNrl5JUmYx+0nB4Az
HtVFkrBDxS5shd+bnBD2cGnVwcXdlbXuRO4iPvUxlumvVPgYVBkNk71l1GLFuBAE7xaLwg07JqZE
L+d4OAPwwg0oaM5tO9sJrksJRmEossF6pVGubgUypKZG+7RyTw121MpAxrZVkuOygKxwWWbVL/b1
ZHt93C0exjQPwY7+8VydAyLtO9CRDi21g13qT8ycSWDA5fr8Hks+ABEmCr1CDtLoW8IfWdxcKmWj
1P/+hOl5vzG7demiZPrjxJ9OCHnCpM39B2srJqHoA9sYF9kwMlaYbu5QDOMwOSWZ+6eBffYXidl7
cQKpBwC5JzRlPm/1vBJgXOz+3UfawySeSU8BOmdeo+STkedFFKrRV2uu6OaJZxyz02mJhgYE3kcM
fANQROzENaxwL4oZ1mbdJjVEEOieoHdMXmAn140Z1vbkquRhJ+YMTgPonN63TsoH49kkSCYx957X
cz9n4PiyQj7kbL/ZhdJP3atebVqkvSUygSy0ajkoUacD9HHBh/Gjz/LsI/5Xw+xR89gaJnvWr/a0
7RPP2wO4LoVf8bZoDfkfrAUFJMD+s2JNajDMjfWhYaHgVkEJ2yu/epm+QJ6fS6kHmYcOshZoVEIU
M/VK+hJ0M+P8Gk8ybfH8hzQiMik/EglQxAD9XtKEcAQ5Fq89JeOxjxPtZgK7iPYivGdQ3tZjgLVI
pyIs0n+/bWnyX76jIZoxlJYNqPRUjfgix/8BlFKxd3o9Az+HzficQHf4ngOnKHf7f19o/xRUms+z
INY6252bueX5x/Gl7iBKl4H8a/G+mS9Z0Es6zZCnSIxfjt9UB0YWkPSvGrsA8D4iTjW61D9voi6/
Mu53tyBrBntkixDfPKcvglZKSQTyhZ0BwWy5snpfzh2FZ9wkF7vzLPYNzfAGgLyMKh/S7Bm8r/4v
EJMBm4oYVKXS5ghP2ZVl95WTIhgceA0ughwAGRLTuZu5ZaHwCe7eJwPKTDFVcmVdfCQ8nw7cgQew
+SLRATnCq/5GONJ0DGX4LlQm242FmL7Zbf+Pb/XYK3wNQWzo3h41Pm+uMhO1/4Nk01b3nsZTG3HU
2s5RJNOPpBmpS0x94E117wSDt3EcwsBI424OUy5Q/Nz15shnj+6gGBvLJGfostyNwz89xeCGSeCV
BWtioWnT4u7Q8rbyahTW+uOZ+HB+pEeXf46u+zm5hAAZ4YFKKfBzGIIc1XaUz2Qktataq2DWGSGT
8OKXeO8WYkd7GxKGRFMCQHxtoh+Zi+rMjisBSBpD7f1BN/OQCQkZRbSK7Irul8aeWOT8sW+Mf6fn
Za6JNA971lkPgSHYiuUFn3IiodyaeS1/q+aSUAbACfvTWCi6NaoeO561kfzcQFmCfvsg2nTJorMF
zngYJtcT8azUv12ZaU7nIe489f61GjFbhu38rkHGYsxyal3XxqprqpHmtkbh16hAphIbsdYlnL/B
k457azS8iRTbotwfPW+T+wnumg/CY0wr1qKoFWSGNoHK3JRc76BeUHaSnf6kn9tmRN6P/4mNoZRt
J3QS+rhTLu5ZidPjomZd9pnK9RG+mCLcHgJY7QZnuI+U0vcbjPe6CdcN5L63NV0xioC/aYnqkGhX
mSs24GnpTmrCICgAGhQa2x+884jCx1uKZWdB7D2wWqJvLbyctHIn70jis2ewsSUzd4ORUS9qeUxe
EuGOXNV/eXVLx3iD/UWmTtBrHIdL2bUxBw5vxKjtEI+wrmR/drkemQ4eT7/S/b3Epp0tZemBOYnT
ph2Sr3gsrtOk72zZgmi4X6iYBC2jKt4SXDubLWv6ZKI37MlI/72oPkw4muyy8PHstNkVtX/fAAMA
kTueKVydl9tVaRUuUbnaeOtrVA9ed2VSaughJouGQJq0QnSsRZB441PkeIvSSsIMHRkL1CvJMFih
DDwUqQUQe9abvG41LNuQcwIWJecYzX2tJZzQJm2RliQc7EQ9DPWkuUbAqT1xPnF0TYg5KUIGuEX9
9x/JWXkmpimXqyL15y0t9FYqho7IU5eG8Ez6sMCHyEuNnSOzIJ+qRuX0nwuvDQRFbK2JCE1in9ZW
qWXSLUhe8tq/rvl6lwu9FCam5r8+NR9zls6GZ5ObE6Aqw1fYrUh8SS7I/jHtlakagxqQ9LoIzXEB
Fakla2ZEDBShnPeBygxBzFoFXW4hYV+CaRInQTXWrkoKd/9vfD8W/wZF7kVxsgMgMp8DpBb9g0Yv
vYqKP9i0AwVoWhYIy9hsXqW1TUPmIra4kNUKZ6jQUdJjE5BqhETxFZg3BQ0JLoV+jVE9fkYsWAbZ
IiLhmwXQxxfhFV6B0vnqx1NuKPVEn6EDNd9xo1f/ET6E9bkrbehDnkwSI2gp+s5Ujr62jfDq2tqh
7Ku2EVN8QCg3o5PB8hLcior/jI5prAxjyNCQiyCTsxYHRffy0GHEkLCbG4eVun4YSnXcnarRPFzI
B1jSxj/c8P/y24aiWeXYp+PBtmuxUPcBiBv4w4aaK7xii1S1TZGQWuLMaYZZKoO1bza8jDk9BD+A
VLSveFU4BvEGvnAEOlcpdU0BHOd7aDCGnlLOPwAfMZOkZgxRBzUTN6Mrckp4AhWwnPeBuU/teyaa
mBOd0zYS8vlMR3T1JWQopmc0crMB6hiVnGb0xeFge8gZ6aHc0vS7DgY/yyB9Iw3+0kmyfvFy2m0E
K+g6IBSqImbEaK02M/rQ02ennN+vOkOtYeJTitzJ2VPeoHvdoQjr9gZQ47hjjviRQcjOtY72QsAG
ECQ01f4c+6LDmoKUObe/ekkEI745D9MyCy66uCZCQNiy64u0wM9KXVlip8XhyYwfksyGLb3Nz2+a
eozA2j81nbUDaIMCMyF/HgmY8yS/7mRekc/T/oKEGonG9XiWFNgSWBz4DvpztpTDiq5ou1ndJoND
4FYoy4BXog5nW3h0LbTN48mtC20oi3YbsvvZF+gTrBNlEA+u84Rzk6/6bceZtCvCfgEgdtSDgucC
d+jQcfSmfrfUnHntwwqdhlPUHtPivQVjdigLTZbUFQduvIjpRzti+AVtbXkbk0dP5GDNmZ3QDGNq
N2N/LbRlFebwvZoP6QsV8LeOJ4se/lqb8DFz+R1M2+asbjhTr4R9saPdSzQzZJsLO9Og7QQHLqAx
It8D7TCY8x6X8tZvX7a1XxXaHmKwdTnAWZ88ia5T1uTknqdFauEqTm3h1rshzOzQAejMhfUiFOF5
NguXwb4P2ofQZWPh1QjW85YSlMNm9ipaNPegkHLNitPH14sFn+o5b/pqfe1VB8j/1wKjNPV/tHY3
w8IELDIRNkfbQ9TfSEK8Hdg+L5ErWeFqbCn+LJjQuIQGCPVsd/UJmi47zRSTg1vPxxcDWw0mJIc9
UkM0eDSwI6oKl80I/8KWAxV7dD4zd7BIUJZKb56xhM7Ukp6KXsQGidcz4XgZZ370SfZsQZ426/92
sfkp0vUbV2ezQSp9xVL5chtRv9kcqOT1cxsbtw5pcNNIUJrb6jWDDFqulwQtxwAsaAqZJiGxP783
rf03L+R5wbGl2ESDLBgaYh+QJcCDm+ly64aUUkDHa2ti6o9tnSUO4arbbDWCfeSJQTERF/yfD+Yu
xoFPtIMQ9VFQnUnw8Ho+oOaOKviDPSYyRipitdocp+nP5GEwPQZ4tQT98G5AZmfpXPKPvHaNlWao
52uSo+kHeqCnzs6TWXnXPKBu+Am6KWXU9gySQCgKJMcd64upi8JGbBvVcrmcymH8ST9sI2u8hOcb
Dnxyqqg5I2Jf41HrHl6m0QTt6On9H+fw2pRqdzznj3OV8ZWHkxisj5YPxb21sqHaYhwX/e01Zqph
z0F2CzxF+FeICM8Ou9lCIDwo4gC1SCiBV7k/K/kodSW1YMLV0fr53WqtaxfRt6eI2XWaDdpLrIoC
jr5PPWqieZtRb+d1ihn6ebfRhr9fs40pBEEx+w5CeFXetpxjx8/rcoG+8b90JpWM+7nWkMYLDTGe
dKP4EvsBfHrlJlhqNNwgferIT4aWhLvmZnTMUuRG2L2xbFLB/Eil5PZjWvkJpjHL6dtvJzymN6Ot
ePDjhanAGuagSbfxsmR7F/wlFwFL7pqymcyZhkTgNoZ7Jf71UCAELcSbIyvlG1FEPJTllgQHTj4/
jsPgNy4dVb07jNbYT3Yw2mpzS6TenVGRX6Efngyj7TxZCcrGgnC1WJv4Afi9T5f5ukWaqFgMZFWx
aYy3wOVgkvKgLG4QFIk+9B8lTEKT8F8s9E11eNdHEzY36+Cf+4EUsk7lN26iSSO7IUvXJoQRzzHG
EFytf6mGleJRpKRSOQVRr6fTmeoShiar4why4CZ88Q299dVTe+01id9PX1WFZ3XYRUkGqwfKqGPL
OJNIzBB8m1gL8dDKd/liDUAal0JsJwGcVMVjwCIYFay11LOOkOY+8n1zlYqQHneYI6GtSG3YXHuB
gKk0tKI9A3Rbaswc6bjzH2vaXSPfJCViNK/ZtDgh8tqyOukOSXwM17TN+atLnlajoypshvQ0mvlT
dX4p3C3cFkrZ7azkSCldSU2rh8UoClxmnqf0GmpPANa85LbFLkOtXBFeiX5x8bEAqSoKcU0geMWv
gx2lTzRLB81B6xmiO1lSPSksCRG8Lli4HJ065JjuhIjlElayoYiIc17F8q3rGjuEgFN/twLYkQR5
6tf2k7j4Kx6cvlzbO675w4Ga0di2HehkIwJEMaK0aUe/MjnjNHwigWqLVEdVWOqnQI7o2lfgjYAt
IYFe3zyNb0ibRYoV6vwFBz3zX4S/cEjw1g89hONBkJtpZOiZHtJLpOCrFNCBkPOZzkEhb0g/kPPW
lHGEnQF/oGWKF2ITKmFa5zz2unFeb+azKZLubD+PdG+Tf2BzsXblur4V4JpLxgaKdCj7pJ58dhyv
C5zV6dzxnUgBcQyTmEeAi3eLnUGsAasCbsXTY/8/0RZJnZWAOB8eR2elcja5zwg01uUvDRe+4yys
M1l/XNPS6mbwL1cql1UzXeEBO2dkTAAN51Gi2Ygnz1UGnI9EfEHn8DqxchqzoO9Jia2Yc+q0FuFU
go53yiIgPtY7gpHux0bliT9FM2zJTwJP1aI8iz0AHa9FKOBKv3qRJ0C08T8VnZr7ANmzqLy2LS4x
CDV0DPlLMNbmOMrv1n27rV1WMST1UkWMVuwgD9fUKTg8STiee5EfsAoUL/H7VhdvXr7CDsfiVEl7
lcaDh+9qh59A7mEBX+a08S6Imxycg4wyvlbQ/Vqt1R5+BJC4KIYGx908YM7zdwRhJ7ROrWgUAjAp
jkd5sC6WBtYASN3h22Y4fk31nuyDfkuUHwh7iPKKRAxZjUOHCUn39Rw5OMEBG/DAMk5WBNuzr40r
OAnMvdO68RIZdVVQEFtgLbN1+SFAmxpkFVRY228Ud6uYPsHOZIq/lPAgXVdxdk0NXLiV5bDb6htV
LbEKa5kAyENXJurY+S32OJjjuNoyFeDE8lA/DA4heCltXx6axWbDuyGH8jiqS6zsBaba55Ljzg9s
XJ6+c/HRlfpsPNsh9zPKNHWvqC4hj+vnfPspJGAfspuuWwUdMf0YKRpuZ+UaS8aEJHoE66dL49ZB
Yl9DXC/HXE5D2sSB0POwzvup7RVgO4cAuX8WdoylKAhEGyd/O/bfqOavNimVYdNVK9zS+Wa/7W0N
urdFXC+g/k92o7LJzUCg0JlEyuCMTAFLZIta2h5Sk6Z1RkRZayCtwvCmkB3OSuqOgdI+Sv4aesWk
8Fc64/cQyAMLH02OYkx7R5rblRX0Wa6xr991530iRtOrchD1NP9pbXcgqv4dq1FoF3Us2dFIAz/2
A/4MNAbPlgWiuXNN98jg72aH4iZjncsBHoTDUetWsglurWXeBA2N9B91gbUr4xPNH5idSUgWwzsK
5u4YNMVdERPc/Dhn61+vL3xx7WOVHDPYJ51COYRww7lxVVVWoKQ2GTZfFvRBjUQiq9N1woFcpQxu
/co286F8wEFVEJXjp0LVXr2Za1Az9EST5hk8UPA7DIQ2AxwitwBQu1Q/qHsZ6mEx5qVw6xK3mjVe
662CzXkaq+XZ94npA/hL0KZ+vlFJ82J6HdZu0GmorNTZHZQGd9DHMYSHeY6dLGLeehQDzEkMdRwx
LpT9S5ZaFJanlkBogaZNB6StmLQAu4V+xLqJOye2ZoRda/n0Y3rg3vzfMtbyAM9AwxAeGpD8DKJt
CStKBGD9Ugf0JK037Py0VvxUoz+3GEy40HjTx0JwJm+z9p2GV9omgqxO7s1ujvc4O8tRnNkFUjV1
rIdndN32H30lds6Jlv4nCeFGdBmxLNKxsAzDVlwlJg9kgWvDz121q6wAgG6t6L6bYg16sTstszq0
pN1MoJcIbNcEu/Eo9hATECz8sDKDkcdFOwlFxhJ37jvwT6ggrUxbFkKmf8c4+Q5Rkx1fXyEkIOn2
IE6zCfce9KhS6StWuRpzsdN5KChPYdwekgOyFuxZW+pkWWg9YcfT0r4BxLXelPmBr18NIRsIJy6/
K7XNXaw04inj9mwimafwKzczvjcQW+siE1JSEHJPyLy769itfD+zc1T9drvhwFGSzm1ekmUJbjqU
3ZPz5jydMyinL+hf1GlwMaUYC/ZOi8PQ0idxQAVUH5/rDaMu+jZtNVznaUEYd/CTRVnn56tTzI3E
pl4znW2un8MzFdvhn1lDWQ6ZKiEH0qvvTuYEAGXYUsnW+tBByTmMy6VfM8Tz9t48JEVcVHIQhDJp
pYO8JHVv3yePOQ5dPH1WPGaJ+cd7X8aKoW50ZsQkk/81HZMraRVJT9//dmveBX+WhOfqN18GDdWi
baCEtrmhACuk3Iwfeh/6SfjYJh3HpopESJwhszAFmPX3fh34Y9o1Ncf2TjOyO/WtjycpQubyehcc
p2Y1Y0m73Tc7ds1+1d9yrdT7mQY46ql4L8mQnJi0DoAMFECax+DfI033bTJAMkXUbju4MefKLuEa
QQwHL6oS5ApalFUD5qY6pc5sbFDd+B0WUD7ny172eaDzhHIcAz/PnsA1LTfflaxorbp8vUJ+4iOW
fjIVebPdkA83kvQUs7UdlWp4U/rEc/J3sA/+sSOANe6efinzB06IiOHuLm9mvh+CqHDvA7XrHsRC
2079jCHiLEQpfUPhR9Z/v5rej+H77OZJXHZnlC41ph+HnmsewGHXaAgCTy4q7Dxqv/EMkTJg/O2J
K8AbRT/98aPCHsE2y413Rv6YCzJfWhZ2vQieakeQjj9M9m1pWVwC1jNPd8gsc0Hx+JrYYFKnd1Kt
Vq+Nxnm0dGwJ3YWXqQj7SViAvMozZgxzl/LKsYCibS7gBlJIi+MlRh+SOtBPNL++QmcmuZqqhwXO
6v2FjG8T0636tmx2vDgjydYdFBjuaz6hKXidRutAAKqyn/P2XzXLEhQEnRhqyXgigoNMFNqo8MN5
4MJN+WCIfg/DxnNGlLhDxGJh6+7+6hm5a336u1tnYHneiQ2MEWd3h9dlF+YbeourVTjN4RbpRcII
s3q9aEOlgNt4XSwsVZV9FQY+yuwkSpP/IaONmV7Bk+eOipiWGhwcIQzwTEvwwvxkmDSeqC7lgv3x
izlYzQ2bxk0DXXu802K0554jP2ZV03hPXaRaD4PkUjwo261GdgbDNW2e+alGch2Zh11MYDLdzTPy
/1avo0b00e4zQVTcr4veAFfT3NqAbSwFnQjR4jYB9nAbRmcS0aPacNQ9+HnSYbMpHmz3WsCPPPbp
c7FemCI7yAT9pmRZrOiJEmMr8bCZUWRc/HcZ2DGSFPif5nx5AOLxxvoQs7S9yLiJxN03HYiCbTDc
QG+s7uicfUW0m/LvM3MpIglV7I1jpzXist2NYTE2vH6M8pwpu111VwDwDLGAtptIATpTk2MUW4eR
Qmu8p5n97uGBj0GKYIwpgrxDQ0KIEZ1Wp5vl37FcI1wKd/2OvcmME9bli97onw7Tet9LQxzavd/P
8C55F8z326yC9wXSSCC1ZgS1qZCDFOe0++sM3nS4HqLYpwEmXZ2E6ZrqILX8B8jk9P9kYv4jnBAE
ftgP9fkzR1VYw9IT56giZgJv8eABxgvA+7s7oSw3ez5MGIERscsbJ9bfRmolNHRoyWIWFoXL56ys
urHxvaN5/2nYrnHYzPEtopIT07fLJnAcsBMYL3emrJanFOLgj7qXux11hRaY7vmW5tGo9LzRIYrR
tH3OKFTMDwH1VzDLx8bRfappPEdtjf+gEdH2XUDc2W5yrlcgCw6GO4XdgCoKSNWaHonrkK0U7Axi
tXh3wWrQm2KyjnCc83cW3/aF1Mbhmia9ONcO23h/w/q7Sgr3psNzwnU0VtUeaEOgVTf0h67VlvP7
Jyc+QKDq2cndxSCB4odU+v+5+cVLBI4gYn0obWYyfUw7FAPDlO8RJOHzubnZNYAVTfZhw8qdze2c
cBaFwGT4LYBQUb/D/MEO1KbiieKgtaKmsP3r6vzNv1lkKTerBCE+lpfEuJXv4nYzuMgGwHBmx+ID
ogjset+QSvVG++gTGtJzQXi7A+RhS8TY7rkD9d+SEOCltPN0d2ZmgjDzbtCL4thCX4jh2wkuMCNZ
CchfWtogiaZf7275pDiqFsc1A3d8W8/TfvX+oiAQtG3Y3e9gitk7AXflK8EiqLD+tiuljYWaXhYu
VZ1p0CfBYtPNZw51LHQelk9e+9JHAiAz6XROv4p/bB/hYcAXixgcYw/YDooZDm5pmnKOnz6zQwKV
ZbSekDYYKQX4WxsXPsqniAOYtrMBsASOX9KJuT5hOzR29aFCyiRlFrMyAkeZQQOMT1Pk8cHDZS0R
35vtdVtPj+TludS28f1rNAMAOMExvAEFYOq0RAVs707Pi8NIXnbpGAcJK8BYcq7kAIbdnJ/3AEkV
W8AoJV8IMk41K7Z3907Cf9p2rU3fkNF1KhSEWXe52a1SVGflzA6cf1envoyFRcpAQ6StlwTTmCqu
PI4aitVlfsWdcZJGGD5+sDa5cTu/cwusn9uaAEe42iCB8AC35U/hl0Xg9DsESplaxo01GHnj8T0S
vGnKaTyBdU2TOE1FRFcN5Y75BGzL1pZGWC+o9fODQVki80gsCYLekIzFF2dlCYoNZYByZPVkCfQc
72Ge0QTnwXJcNmMsDtQsCLXKGIMOVKcpYyE6mE8n62wy8qOpXZuB7jMRD57l7Dyw1DiOa0plXgbT
Pv7vilmv0FEW6QHxE1qKgDTSGSaJX52/79vJ0+LNZsmAfzyUcVWlGyI7JBts63LRPlQCtY1pgYcJ
wT9d04bXv1hTrM7weHCQNmtY5Ki5z5UvpMPj3c01flyQo6nfOQEUkd64UzKhjREfqkmtJtAoNskc
cow1U+j4PL/00a4hl7OWNFcFUAmZAHpikx6hkDc9WYCi/ep1OP7mORZNcS4oYU9yrJHROB8PN97D
2c92c8b5mflmj6RMnIn37/kRHdr61b/yrn0a+SQeDe38GJIgaOV1T6P5l+jdH+dFNhLAz8ehbmGv
v3Qi7T0OnBw1T5WAy2BFAUJNVXLkVXfN2DU6VeNjITBWzJ+0wHqSOO8nwD3BdSx1IzNVij2DQDI8
yYDFR/flP3GMcd+B1piAse3tvWKTggFQi4813omthRqwWMxhSBdeF0hvcIm+7ag+2V3aHFY6Z0Sf
21vVGNa6xt8u5Ys6yt+5PPYKMulpe4zVh8050yu2XRMndws7eos24UQ1VdU/jHrAfz9u/HTNoJ6T
+MSkDgNdiR7denZ8QSvYlax3DFmljT2JfZaxAlFfivv2yIF9MhPzUEey/GDIstvtvxbxotfkeF6y
BjDz5XTTHbY2VCO1q71xtqXeWcm+Vq8RQszdDU7ZVKGtPofNv+uUKQEdGk9QwaG5lH5PDmqJ3Axc
opcy5wibCqefOCmhL0XUQNEeFMGh84yNGp5YlVb/RMth3/fax8uRFV1e4gHjeGh2YgQDHAe0EtOU
aanr49999aUfHYgKJeTtPdg5998elxxbAea+YHa1zpFqAvv5AyPscS3ko0UdT3oSN9Q1HjaJOCsZ
JV7dKo59JXeY6Zlw/EiGpmSIReE6CXKmtNTcZ3PdIVrJgzvsl9HC5rzOcXSLg/I8C1GFWOI601SE
TMtFk0ir67WWFAkVQjwhT9/bzxrZBMIHw9DOnEPdfZvgUTXDf/iK7NXSqtmjztqq/cu0EviqJF9r
1fsrjxI0Q7BpwRFqX69Z4VcAvNN7BdVTCMzFvFefVAyrvz+xoX8P9n47RLQ0WUcSM5GgpKKz8aHw
UCj5GoWMy0LjY326alcMyGL1moOA6bLYD5mOj1hZDz9FaVSuf0hsk66Hd5Qacna5377FuxfPdP31
HqPUUEEOQ76MXcJ9Sj6ujk/3McgbfZKMxvZodzC/nkPY0oCscpwXwAOF37zeAKeSbCe4hhpaKui8
lmGL0JPwkX17InJ9J73uaBN+vKQx/stm/qQ6JTvSlrLFy/0+dALXQvAGdyAp+yftTOJdDRqmPpGq
jpZ3u/1l0sddj1M/mxC4XbSyA5IKlHK1RDkWDUMoTpMPPGrJxrVgb+mNnGv5idXYZHqi96qU8RcX
mQXBajjRsHr7BIUWZrB8dtuOxFXN3W++Cg1KIDlomDjqKed3+LXVU1dOYgSkoEBSQrm1SHQrl3CC
m31dfNUHaysXPTU3McNZTttwRIxQdTgMe/K7aGV/ctaHm9KHNSiiO/2/+i25VZYP5b9L98L9bjio
W1g/WojUBPffG8V1zUmW5zeha2j6u4OHJRA9f238nzFnzhzl8U7hlBhHugsJWI62yDfAsCK2KjZT
L1TESw25PCXtk5kbCkqXCAQwA4kon2hfDJGkIjxsbel+VicUWpa8056uNF0ojKHroMsJAg7ZfvFG
/CRgJmmSBHFakTbzM4UbtnNhtiYYs1D8MfjD9Z8d0zR37F3qLlWn9IIzQY6OuF/QfW5tVzWoLkoN
BUYSjzqyS0MwunNFsZfbalSktwiwqU+zzGztxA+oiXCz8TuNdfvmETWIpRFQZUedJloLJAgEg/1h
gsT/Ku+Vxf5f+Cqo0DOdc0c3YJ/CAZGnaV0or4A3QS448CmJ4Za71B+xACHzS9i32zgwlvaXt+yu
y4iQFd5/aeCx6DL5Teteo2/zkpe/xcD2F8SVEt5Sci+fqFoo0SWCqjj9wmc7v/THvFKYFqndcz4H
e2ytqJPHrMUXbiN09yKkMbctK8j1M1HhREQeO+sHL0ihc5facFyDfr0n8ff+jSbFo0Db+92lduCw
iEQYRYQQxKIp+LnnMYRPZ0rknkhhnx7hORLJ9ZEj4ARFMZ5qwUwmnScii/S/9aXUEZb0WYMXyhX4
YQ1FNz23/XdNvsTI7rAmc5TrrWLE6c5hfh4mZU07oW/RHryYb67viLcI3xj2gfhd0/JdBTMsyBW2
JjWidADxZhlMxb9qwgeXTYbY2xTNSUG7UjGm5KX8Xtv1GJmPCkK2OuayVui8maL9YHc0UJfWwPYe
DtwotzGa0vh+hN31v0M620424tRB9J9PwY9TrtKFUuoo7GSmB2ob2HziaI/WAViTSF0jIypawNbQ
vdlC94mWjWeJYPIQ82pG2g32vAXQef2tf0JMfHBms9DXtAw52LKce7N/1HqOCGzXNdWuh4/QEKDd
BAH6P++AeoCYeHtLQfvdN6MctYBeipMbKs4t1FTuNlm8X+FJPVIBzrq3Z6ct6Zp0WndlxRJSklkx
KHCiWBa1BPiVGHL8Q1Dwsppx+fvnixbH+fg5A+oKXJr8mleSdfPLFgXn10OahAumc6/MA6lNC1J/
Q4Nd19pHFU6Ng7GZzGiGMYZjjjU0CVTjGHXTqLIJrXnNHyKLkaDNX2a5/73lTJKmyBChbfNOrNwJ
ZxevgT4Dy53bocNZn6LJWuK4Xq+Vlrt2e/QjR7rMIVCKkH7/0VprYx2B1xlBZ1trtowFieva/3eg
hZ/sqt0ElSsJBJMU/KSs6h9ALv0p6MBncRGdCNVltLirWfl9gngDO4gl9w+ajEK3tVEv1UjJr3Qe
pU+R+OuUHhjrFtZ3bqbsW5ySS1/7AsWAd7Ploal8V3i85LxnjMHTbfx+QH+F8Iz0+V+cSrNoG8XD
4vuLn7JezRPUpma5gG7j4VpLd2fZ1ObhwFENkSrf9sh3+chUhKrI//LJa3vL+p088UIPvBL43F8O
O1qv7dVwEPTXxlf4nLMqDtfh9cLTKtvlcLW7VAjxsjl75oPrkwCg+NtDrcFIVaDaoJJHAYHkYGWr
MtYRxhyT/ufFulxRgvENjdTzKevPjtFCCKXEzomy9MrtmQ5jpoV0phHnq80qE2nMTeXafnVe9a92
0l0mFgzyixCyHqpudDPCK44NBwqa45rfMxs+E6NbrfPh1pbyGKfGrIKZie9j4UDLmS30o+Swgi8U
aGkDKMpDCv7NP4/j9aFSFH5C/KAATR6Dtwda+YU/1M/NhwBCzbULywKUjZdQqVN/ghwr9F7f2r34
sWjoNFjIXUmbtPTQ+aUNTSM4VYitgW1/eLmWOGKMIk9I/q1R3Pc6Aw2OSnkZn3JFWAu0n61Lu/RV
0DtYiYFpLOTqOWDcAh+ep7ZGQrYzMfjpLuxSEG/oJ44D0+gMc8g4yipCX1usxJfnXj97AlK778bZ
uj/zbLyNzZ8Vb56Efw3UMqWgvf6WW7aiWNz7TswCt4tbYuzLuqkruzQWa6/ypFmLZXYpe+Dg3mp3
lD8+mn7eIj6CFF+dq6LV8jfjaWiNSFIUwEcNE4iuN9gF4xFKyDn5ipT33l1W84aau5q2BWn7MvV4
Bo+JhlRsGktZ8fegEXrWF5OXhj7mKE2BH7VB1LGqB44OSEhPr2BgnUesipp8j8gt5/05ZmS304VX
9LeNk7OOYzKm6ztMCifGzwNn5uy4++X7iVnzlcn7bMxaI3hsMqjV1wDY/awAprF00pqSsK+Wsc9R
anCcY0ScuNLccEFp+MwkgkY34AB4jqD5aWMG75m/SL53McdOpW1jcMKd0p814vMNoMxMViLlA3yE
GogTWpb9Wf6EaqT3Xrh/1na1hA/tvIBQkZuip9wzEgxEWgMHlRJYwRmmBobQqeOUnlQbXqCZfu0K
ySQHTUo4w2D1HfzbMPwO/N6eKI3tW55Q/nZYfuGDHcQyoDeU0Qon14HCIIUYu9l0rYi6Ezzwjsgi
QZnapMxJ0ob2TWxCG4vLKMSbxy8nvbZQnecs71OziCygMvbeMKW80J55/l3RlxG+sqFsQv7R4Mfk
J/oY+N0h4bwlkJS3lF2M7VbpTrGqzYh4WP3b1a2oUShCEnch0ZBuyloNg6Njwuc0saFKiBSA31fn
KBWNfTzF4Vz5+PGhJWkp4/8+gynt8fhR9oReafEg8pMdWRNQl9P1nj5RPpDVx/icmzSXbJHliD4p
SdtFStU1JoYxWW/F23AxRjwzyKDAY4cQRquhIMVxSUvAYGgrpODac5cjYq/a36lYnIBxkGSrs3h/
ubri/BY9eBuUVJKUQeWBWGn4crZpIBUv6/pgxpaCLlgfSJOfiQQo6OUTFyNThv8fuAcqV/1U+7Ka
InR2crQKlOUJ1iY6ejDGCvttnrCcCSym9ncLswJnoo19p9bzbcDB1OkYFoM9SEo/5oNuFOIIt5dW
r15mImcuh/bDCpkxoYf3hlqGoqLJfrJMsTcSth7h3+i8Oq1IqBB5OQdmZCpHuoc+qmtUZjp7u+uu
ZV3H5GPXlq5xvAQto6wlw51quhm8Nk+vH+XSHK22qxVU/dGbKPZzcbNL1B+zxSrdjsCFhn2+6RTV
jCIzQvbyX+onMI8Im2cF69DWXRNZXqWBemS+l0SjeQvktUHP6Olp3pNvonR3XZHGreJsZ7VgdC7t
I/MeEIIU7vm6qkueE/ubsxB53uSzyIESJhhcVMBzxMucrJ0b4Rb/UxwjAYQJqKrJkIaKfMCV2mRT
1w3ABWSJ4TPxSMg7pWtzpzWUUFeXrelmnhV0x4KOwTsJoWwikEiiFWvINYOIzo/1nEdVBSrRHhub
o2ZM7Cqyd5JMgaSyRpTF2YCDlTGmVngWDVL+pPw/uz8R+gU5IjNdAsYsPOIPhi7ZwDAqmqXlc69O
vLpyC0loUOvE3LOJxS++Ii4gXxvvgjlmPbas4iwFIWIg0TAoKT9YxY1DsJtqXm1BkmZZ+QgKWgpk
51Jzjl+LpD/b7YHnDzORYBDBwrXP56bVoZfQTpG/UqdQL6FuMQ9zOXV5zbnyUA/2AmPcxvgExao/
UC0e8N9UaHIZnzsFwc79Clgj/tEpUIN3wH+Vf3LljNcxKXzuwrhotwWJatZtEFIW31j56wmfqIKx
AkHN4USxq0J3lpksgdR+q2CZ2bC0gVI67qgATagFZMKFkP12rGSZXTRfrRzGW3jjDKP3tH/JV8Wl
KdtxBuLYyWOu5UdNqGXlnzCKPjjnIRGcPhQBaaiXx3yJvScF8wMnT59UDO+z41YW9pj5UHG3nXam
4WMf1Wbv3w5KPIaNOIGF1Pq4Dtuu5X72sxFxSNv6J5smyPtp+UxfYGnzREKWLWESp1FOr9RfEGtA
hcnj+2QvqwGuJapPOKgtnp+QzFBcd599Uk4hv68mhs0cwlZSKkVeMZnissTXKbjF9qCI2XKv5e4i
JiTDHUu7IrfksBnMARSqaedPg7zXNvvtso46cd0rV7Er8r6KqVyUXCgbC1+NOG7ujptJM2s8+4M6
Gpc/efE990beOmU+Josi52LfVY1NoU5/QnfFmpuHuohWTlBoDU3uLA0CYqveeNavE4kNeqNEwR4v
clW0sESGg8GajZGTdL0XsDS9LEkNxRe8ovDLIBQ1hQl2sxWzWVvS+qdZsWVSJ6yB79CjTazhrjg6
2o8E0F1v0q/EWt+asu87OCdtX1CY9OWcU87wKhRZRfaszF2/2QY7yNJMXwSuPD699hHDNM//4P4K
jlwuNQiqr/0uZC+Hh6tKR29tXU9g0Tx2lpyAptsGcAAJGKats/RjjX2BOn7y5FyXIqob8lcDHBay
RFiRyr6HMLrFmwBqVhltWXaC+f/Yz3FxsfgLPWDiFLW0DWgAJvjr8uEeQQp1lo6KWCQIeK/z4mIj
46p5Rn2c/y6KlIw8d0syeURhC8ZmfbrUwQDRKF/36iAso3qxfCpBkU8gGTsK6//xH0EWq4wZVzgX
qXUZH+dcgzRx8Sxw9u/kjKnWHJNkJ78+z+ZvVYY6sMbk9CcUpVCmC7aWKAnF+1lO5bCddWZT678M
vnQp3bQQOhIKrs168vN/ZEoFAQJVAsSQBT2VJCcOZuZXgA8n704VNQ4FlRCaY3h67FtKlpye1e0M
ofLJC+O2xWaLcGv5Rc1MNZafbZlwuucCh+00AbMnad5RxdWQjMbzVfcKAapQcuLJJUvdY1HodaA4
rHE3GvRIbA9hOOCyxywXEoxEHTdzj57zNcWH06XiSfJoEsx1Buv60tnXVa9R5n8Qv2aEDXitF6AB
SVP87zvu/dtbF0T//17XrKMLOu4G2vDiYU9ovFuAwYjvvP9wrzhQXEI96/r9LQZRodR6MFwiT/qW
hGiirpIWR5WgZy4Uk2u0NqX4wcvcDXSl+FWIwFS6Or51ciZ79N2Hhd1PIRDh9jZ1gMPYzByek8nj
+ttQsgwN4yZiUXHZMJlsaJAlOieOrOoPNNp7B0Dg4ssiQgyCamwhegQkLBH8yXw+BfNTe/erjKqZ
roxsiIWO8VrYH80pDMdrLcjeolKZywJWfgE5BeFRpTMb0EgEex5KAtLRqHgNmHcW2Nt61pEENGn4
FXrocBVHSE3yuoK7hG5/8K0DVHFM3S3IDA63fRNK3gNETM/MxxUsBlDKqL9ZA2A3fCJvxiHmaWXE
TQeHzRDN7e/jOCOvw9aNmkFa9mhPGAkBaW6IFgJkc634THcAtqYrUgDEe/tJY3bODfQ3a8gcN28h
1nrnVPNQyZzAnbx8wG5+wzzsRv7KWRxbfkYFksFhJ89YaaPEpQ96M7De05b5f2toIld4LqfLDCck
G96cWvwU4qszURKLEV36hZkbGqMNJ6wB5GB5vY2Z5JajNd/9mo90EYUTx6kUxequIrOHAS94jydD
QLUi+dTTbHtOAVeKKj0fJ5xJSI8Fk7XAKVKphKJyQ9FcePMNM0S42F1jPRbrcmHYaB/xcEPHlH89
jZmKJ6FqlRG88y7YhRx+6LgRfqRrhXcVVvgMZTq6MZf27oFQT+f0tl5XSb6QutKiWHa0WemVgZaC
SUi71erke/37Xc+3jx11R3luhD0u6dO3IWHFevs1KEbGU0ZSdx7aZVX5pbHFo0PK8KaJqWcnCCe3
chgXS3EPR0QYCug3O3zWpKTkyiYpHf3CFkFIX6lw4tk/rxmexD2CxrQi626vTDGWTaFqRXaPY58i
bE155rBfhqU9CIKwagNVNYdEPLFhj52y+c94g+cayFvtYG+VzIechHkDbBwqOx6XljLVTuLSGFiF
r4cO2tYp3eIzZyykTXBgx+8CIuWqPLNM4QVkurNXGlrm4E//KXZVYeR3Y+sTEWVXtFfQOFMAlyL8
6j2MZR8rS7zSrPJoaD+w/084TTVv+DP8FJ2WJVTUB4uAun3FB3D5yn4FpN9jE4UlYKuyvWAwdhnS
kKhKTlWC+8vL4RVznjUAIcyRceKFY1p3jbk8ifpNzFtu3No8k4HHggjBm02WVDm+rL0nMX1FpVxD
ypTKO3SKaP5JxCdQSHs+1sbpkyahv9+pV9CI3VP5mHZoSXSQDzggm3Q1euP6U8XjcldmDbJSadNz
QNFPVJZQg+FWXj2Yq6LeGX+iKRJ8QxHo9L6vbPm3MmtaphqgV7yGaLsNakTkzFKKpn8c2HWgLEpx
heWwtMjef59tyWrgl0UYfBYMKxPa1AnqMxUvAf+/NXlthW2I3QWPNxg11PQBTjPJj2yeO/WSI5u5
7zLtFbpNoCo9ksAXbkbaf87I2hTksCVGq5L9D5Dc41vWF3XW+DyAjNUlvBOqRybhnKTBd0Twm1iT
2rhlbx4FrheWsv7YxjSeOWwo7IYeAypL/PN1W1DfTglf6/DvFThk5WYJMMjV+J8DquV4SJbLkdsL
gdBIkFbIPGdjzO0LpVTGus3fe+ti4Gymo7no6AjQe8hm9N2dR5MUAISG/F4y3m0pSMvQru2tmlU/
M4U4+c8m4aUtymxJhbsJZFYsswv6OoUvTbi/hVRzgtmgI1zED2jpkWgslQa6o0qbnRtTQDj4pOM7
YPI/qECgZXEIrabICDr+sOG1OB2V7SPp9NBcx8Nzi36AsMCVE8PpWGMpp43hEXW4q+Ozn26vOPUH
04pIbLfc9N2MfHe+922Rrj/SNFCqudiBXdqVONQMLu2sCeCPLPKOMm/a7UP276lzujQer3A+fYXP
4VWGjXWz9+XLwOsPRHtSmXWyxg7f7WC9hkYUIW+VXrgPk/4YhpI0AB9S/AYw3o85+UdWpd4HFIB8
xrvNia4zIvUf4pyR6Gm+sB4S/420bsYYAyzjwVw5W2If5ztLfdiL3N/gWgyQiFQe4hFiUy6H572w
8WXiGOSETlRSjcgEWxkwtbikvbUxwjbFRKK3tOIdFF6N3tvF7iFM0/2IEKZHHB51hf0sx51jT9rW
hiLTiHLseNPqPz/t9DWBkfdr6RgZYX3uuMpscvT0c2UKDJdZePA+h7qBXf6pMnWsTsHbM8PfS21W
Fct49yG4r+8gaD7LUYlJ0/S6W2YQi95YLf9fVTl0ROekLT+jCQUCZGGV1rYWoCmebiffn6rk8r15
Ni7KaeoDBn0JXZVoISqV5chnkMOUjVXChRMT59u5OydPFeuEEtYZPp1Y8UlvJQHBDd4o8rGkhQwV
Z/cvjVR52ZG93Stjdm0FaJnfNuB7GB4t+2jyg3vww12UKcXEPUxj1mZyzIChz64EHnN8KXWP8Jgc
nHFYtztceWPEanyYm2TmgJWnLU9LWxFfuuzBOJW0Se87290EKB7gV4n0xaOeVknMBMbwEPUFpdSE
PsnzHVAqKiPUaGC1aZGvxPwbVaWG5egZ5oYfouJJHJf/2d5m933VNQpOlGiWVEaMiUp1tpEeX9GQ
18u/DNg1TOLkJ4H2600n2Mkg85i9Jd6pMNMZqXpgciXLzfm36VCPBPzRG3OXVN80yKJcjJfX7ZO/
jM3oaQsWOHyaLomECYyPc/uFekCfm7nT5xx6+FBKJzjtVQBZjJX1/6FMQ4OW4kqt3BmQmTUwY2rv
HrSqF4EGxS8Hc6QeJLpZ5O+0qgUhUDfnE01I1rnD++fvcm9Ey1F09YVDz43TXtrVokKGboA9OkSP
G70BbZ3ocWSHcebL51PfagMmqzHm9Npc95I0HDxfUhWdq8mB/Z5sPVvrckZJW6gUXY2LB0B24ocL
73r3YQsXpcXxeOEEPYmkWOS95cZstVVpARqWg28HM9PsRK/3bG/hpflXN1H+pcGWRYVcTVD8JIu1
4mYTvMKA33R7U4CSNL9FRHaP5ZVEaqPbGVOwugmvTGU98JA/4gIyjYgLMJqcYZiGWr1A8sPVUW2x
jPb36f+tefQqht4CgnCUWUJll+0CB5ntNTllrnVufyM6tkG6/HnNv0el+9vzmOcsGuU86w096NTp
Dtvxrs0G5Qbg+9SnEUUZpr0J/16lYl7bPlVO1ikiTIO7DTAhC5qsYH0cmI1aP5yc6E6X/VwMpn/l
lM28DClyYhsmIchrVaXet6Ok5p7xkh+D4TcskKFOxzWeRq+QWNXvHfx5QT9ufNje69UezXoMItJ8
PJZTL1ohdg6mhPDgaUVZPsWjG7GU+63/pEYbIbD0G6zjjGUkI2Ul6KpPM0rEriUomwHUrSEnw8++
NLaKQCq6dUYRbhBH/mXNFH5nC5dfdSqg2KlVH+SXzcNtzZ5+/3uANATlMA+3dXvzCH2JPd2uGpvb
i2fkeP5RuVX3dht0oTPB2kXORSOfhR+VRAALtBK13w2jHgVtRw1zVMZJRCtvBxKhe4FbSlZvumg+
4HOnPktJdhM4TVp8GYMQRhkC1728as7VGhiRK1Qv5up9yf6fSNTdcvdwMITGN77KDbJ22mlpcM67
zte0pB6wJs5X/mGqi5E0BQ44skBmY/JFOETQc2jkZjkk9Ql+uNxaaAmbsNZfmHpbP599H/SHXFIs
vBXlWPoUJ+q86RnbUYC70+tTuNDg8MvG1rlAAzsSX95qH51ED0hWE8f83N4EnxIx2BCC4x4FMllj
Zxp9ILZDO1gGRjBpqllPn/LJqYQaM5hIP6xZ27K/Lg3Xh+qlO1d+3Ct9xEONf1pRFnJnpiOLAlAX
KSU/68/4QrRrQWw0TYjm4EzjSLVmeZYH3Pue8osOW2OUP0Nvag+4R+1VzHLiZqJ1QMUkxq/FHmPj
OaaXvfD4eT4Wp53lXA8XQwYp1r3ug8RN5InSYRWvSvcXFyP71p0nHtyI/YjjhFV4eMeTukvpq5B5
YofnetpoWFvXGASyiEEdZ+EmE5wQ5n3ZtSX32W4TSYO13aQvKXDbkpFvSjxijZ/Zz0hKJimJTSpl
8qJJ1vI7tuNul+JCcuavnmt4vI4ruHkpT9UWGgMnFsO5iGOcExnNeUW2NeGbpJTOfi8rxHXDQ1EH
ZjqfMP3C41CCeZDSLGH7G0bpclE9SZDA8SnLN1BFddscLyJKhecN5PMUIZ4ZuNvpgO8k8IwbVMau
L8Vym3i+90p2Qai2pI/+7ZO/PqPRfIzrZSYtCDNWJRB7zZzCvKYdRXk/C4pK/B5RkS/DE6dWiHKy
GSMzC3N8svwZK+WIpmVJq/tQ1IkKoDfPMbyLExJhWxy+AhOD39Wm/NN/1ldtUkrCffs3tG8uLIFU
0N1YO4iJsUwAzTN+wzZL60I0guSoHbWdz0+gWvua8LjW5xLejQZb7HkEo0zPeTVWZWkmiFxPorWU
zj0a5jPcmUFVEhp9zQydDmy8+u9bnGTzqh2JPyHlvcEbKG9KSVz57r1BBVTjN9pUZRSqU9QFJmFq
E/1vjwiAwk6yqaGdt8B005HfZymnfIA5+m2P2qmYyPnKZtk//pWfKIHmshXyyf0nE7/CSr4y60Oj
VlC6nyIcOov3Bmi5l/nAp7EkMUl9hCKtk3pmPaMgPDnQFyNXmUJ11QYP+VD4sAr82ImMMugR0E9p
u+eBY0ZmwJhAMB116yvmHOVYo+lJ2wijuE25feeBbEwsF5ZscvBVcJ2guz3V33YGJxBEca6O/NpB
7sO852oVR9COqDAllYDyAOzVKt5DlR2WN6E130wjPtaPiYEHVKEMa2Fbl8VbZJjLkMFYDZlpb6MX
MxSmpeZY43rWeh38hIrx+pfa9DOghH2qhnyRNlyuqG1/dcFidBIDw/QCf3Fv9LY8ZehKqtF/4L9v
kk+iXVPv531KUcmHSdds6cGbtRKp1zD/cEAZlQP/wdn21HdnadaGzmSpE++6QHBrdLvzE8bpSX8L
H13DQYDQCz7YUfjxc5tvAKpBW4u+0do0lECHmTl/7uDjAcRh/sH3frMrRFDkdwuwZFvtt029m6bw
srr8nsMHyRXVs6mkqhpukY1x2c9KtHRsqEQvKiFUVGYcbYgpLwFVTpp8QPojDnZW8aUKtJ8CaJqw
CZxgfC5TndehU8UZrd636L+a9C1Cf1jE1XK41KPHn4MciIIWYoY52ZvjykUkzinSSZYmHXe4etCc
M4SteyxlyNMuwEIqLpVrcYJrmnKdMGC2BpRDDCCoCLMCggWjam1AD0VohZSkzrbv6idWFw55cEeF
vun5WVHpgmis2s0QTnhaJPJE71ciixrmTo5dVNNfiJPmtLycYplRxQw5wnskFiEgRuh6nO9HTJXE
k1U8RH/iBGD51HGuE8pJ0PjSIWpA9m4RExsxbM2BuWCnsqScoOGoef5i7LurQ+wh02kctlpGO6kk
k7RvpWpPiCOi9H87KAjMIisdBmKTkBwmNm/nIDue2y24naYCxZvGn9aS4VPkSJl6HeYtWCAY9SF2
YSnPNpd0GI/FQOJ8nK2B0wA611wSO5fFwObrzmrHYxW16zlPf3KR3vul1ghcAle/mBCbETQ4ZaH7
MW6WEODoODOaKfWMBtBMORtEdFZmpcjd/zJ8lEOcZRkhgBdBAjV8IR4vzIGyN8mjKv7NYzxP66MF
HOd+62ueRTXjUK09WosEAvymZpiix3cWlrkXIDNpScDyaySZM884Hub0+CXhTGsB/Xlqg6No3ird
xATVekFRxvOoYZEvtM/YmSOOUHjiwZo2SEnaCPahQZEVezW0OfBL+pMdwqQ0blbbf0eay0A+iWdX
ObgCakp5yeAS6Pd4QrxJf/a6B0yYz6OBpOaqE6pjVDBGJxaTywjwBFvI/7pk5+NTx/NrrWSsMCUY
35ND/2SJi+JJOAwmQqEImGHg8YVeGJp642lvgoDuvo5KhnPhXoDvDBlFA6boiLy2yLB5wLc4h/G6
fLQoaAbboAPe6ax/fxuF/Xe7CWJM+E4l5JuG3lk4dEqZstV+wJ7pAOrSQcCw2RnpNRpC9i7MQ984
V5jDZNcUmQm8DQ62SHm95p/ocd2/Lc9tYjXGlpgjbLN3EtFJV0x1Uv7bhxwE2+ntMvLYsdmn7j8X
irmBgMGZc6n1VOPjaITzulOKGsqVYrTpsSg53hhz+k5qNC5hv9o1WcK3+63SfXkZm2Z075ALO6jS
HQvOxadH0eNq2JpkdnSCI/bmYpvKwWvxl7dHllNU5J9wcnRx1XGlz8yfe+A1b8kRdmrlArCrOeVg
BjroD/G5QFq69igQG/4eYRVBDLkTfoAYN0lj6wcSppUkIVTgS11ap5LbX9EtkrKJ1lxL0a6Dfy+P
JvM1GbjyelNUhkIxExJ6/JbcyTvG//Ru9TV/Hm38VTnrcH6rxT3EQEmijYQBKxiOJm/to9u3FUPR
od9ZL/LOjjhZYsDb8HaGbbn33w3J4FC+RZG7G6kiXnMavftbxCNn2BBgvX9/nRDURUubQO9kvWL1
BlXxbdrTQM46PRoNtZsZm/1fgbpIn6qXVpdnx40aE0cVm1GrXa5LWP9Ed75RxlD9cEAAY+GgLkrG
+RW+siPEbHZO0KDm0x43nFw5qmUAeiP+4xHnEanSNwCOIB4sYrnndMLOzT8TTkq19hWSDz8NKegJ
+VY1hiMr2ezP/TBXpSiNm4jC8GnhA+xWtdBKnsb0vg9XlCBE0IIfwAp957BGIbPCymlSOOM2+IXg
cCcCbNJLpq14r0eZKQ4CI1b8JHhbgplKlp+6UGLysR6drVWwpD8Yi9hRsddlzRi1w2qeBQ57dYkN
vTdReDUgP9TVjLI5oOXADTSA1ufRl5MLaH8LarBg4K48O+8jpIymoZT5n0g7i+1Ip7Ac86QNDY9l
BlYNd+c+rE1waT19RrptXaiX9KqsJQXqOcmgXKLVnLGIYgdf3NM3KAf375gllMHhnkw3tY5PoRpq
T41jv/jTg1HPzfZzCsHhMPo+bhFOGsnxRK+Uvy/j43E9vrQhIur7ymjyKqyxTIEbv3I7hSxsgwdZ
x1xs7BKUSOrXkLI0/eaL864dMlIxZBSf1agM/hZhAwfp9tOdw1Ec0h6Lp54tm10m8vzICO77z8v4
AAMxeX1wFy5yPJhKwj9WcyOBHfSUdI2EWjGsRaSEyVZP7fefwcKZmYyTitrN99Xy68gAR0tkd3G0
1marXfqTp9V713k0XyAjrm+Sr6vdX64ZiONCT0BozhBOvnSN8o/uRAlnX341nBWMeOs3vP7AGtNT
Pfaa5z0S5M7RKiFn8J6gjugFP0evLoldj6ovtANqpvzjW9jl0XL8O7libyz6K16rglONqH6Obr6o
EUjidZR/gcgbKSDev6zgyqk1iZ0Vo6Y8fDB4kMFy+BACDdo3EnPMTUCqSoUvRpzyaZldYA29f9KL
DDM8mQXjbDx3JroCt7PtwSZeEKWb79TjyrjJINRo8k2ApF9C2UWggts+8PP10AbYsArTjCK0q+qM
kQIiFjrLncd0bIF11yillh0aYbVYk13NXRveQGWUEbRrxvIDQCj8Mo7+9V/9bP6vyzn8VWupbL2P
bRQRF0fZNBri1fPJN1ETUF1jwy2gF2J98ojqu3ZEATji03BarC2B6eYPeLXrd7gn0Z7aaL+Di/Pw
8ItzLBkWJtDaT2iF0WyksCIG7R3LFS404Ih5NUQj8lCsDWNpUi92qznWrV+R8MxZf9S2xOnDmvmD
xJjvwSBjzAWm+GIPzxLp7ITg6PS7vTIufat8T7AijfcZmhvlUAuwz+CHdNEW1ZloIc2X48HO0fck
OHLe0R92xsxnAWX7Khvg9u4wO1tMQNh2ZH11PfLGjMIFalshplJZcxWCJ+kw7Hi6fzm6MFgbFVWU
HlD5ewdsDb6ZMd7y9W+CREDNAqDo3taOigiBtrPZSzjkoPyz1KWKK/QrNvX8IydIRYcHlHNZSanD
LmqtE0j10hpIHg44vhKY+3Sf5AqkokaJLjqdUNtRh6YbUkLVdHERWoowzbmjZOPJgS89tD02lg4u
80jJPzcFT1Qgig21GCLMA0sVYZJO4nPU5sK+glfwhoNxk+eRO9u3fdVRRTRROB0/lj7ciIOkLKnG
xBIzAVUaVKpozggLnhzPIrMweRT9gpnC17k3MXbhjF0NXo7T2Op1EX2WmbxZytp9RxLEe5JWt95N
kKMHaqm90xtFe9m9XlDFSeiHvqoW8MBuauMACWnMvNdlSWoRvAwirw/DXJwAZDQgCO5/gDpRsVAJ
8KXXN9sFPB52/dIDZ9W56kPdumpWmYT+ZJqbSDCmUkgnfm88XimCgNk2fQbD2BBwnfnqUVT+60l0
065PosZf7PCLten6eyMol5G7xbMaVcM5allDPEdUb3J80ylqfDYsAUlcZEKB1RY1dgUkEZ8rTNKm
7HBe5psFdfW4keKMT+Kqj+8ww4XKo0XPTQPLk0yooZ5MNVSe8j9I1N2Li8dmFVHPlVwh1Nal4pjn
T8mhGyqfgKe07aujmVrY3PKnGGI5WDUDHNhN1f9+ljyuVPCgL+mcbozIKChVxxsIwzs8+kyIfs3j
v4N45Msmxdk202FwMpdje29VT+P5jPBbHtiyEHZutGNIvsGGNg+T1NuZtKZ/7awk61hYH2kpaifg
X+K9aqkUk4wu7y7xtY2S4x2YjjwOlRVeNSG9HK4dcmc5ruqen6ubY9q4YCbzeUFXc5c6nwiy/kZ+
jwow2zK2w9fuB+GRpGUlNxb72bdPGFdO2fVI18MywkLRyL58Kf/UakrnmdcglVnOtXEDqVqpJ/fS
FgAHbbCoVnYCcO9nh4eUVYf7mbjBMBIq/iOn00BcWwK1mrPKrVH2Rrl/wUlKdK44MbSxJ4sNzLEM
d0CGZlvBa6raAc8c4MGeTTRwBfqcQ/cY6CMhEKLNsneQjBqzUxeBcAV8CaszM/d/m4mQMK4R2ozz
BRFHdA46aTmdO9hXGod8tNN0Fp/Q4LYyt0GW1OBT8bgtSo6ipnInS9aZolRq78F115TPq57jP5el
DZJEW4d/5dbCeDJXoAyqGDf4mhAZ+i8XGlyKhjJem14H+lN5jeyfMX2jAWPt6TCvucYcIpnWNFbz
J2X8gvAw4n9mnltu6MUGKMsnU33UQV3wndKCCRkiOF2auT9FQ6MMMyAd6LTOS/dcHxlZVGOhKvUt
5bNNOIt3Ug6CDEcIA0uaHidlS22H/an0+ue5WA8+0Yv99jR4aAUtvrD0fg/UC3TOEdqm8tjhLliG
ZOu7nrasXUG9ln9hnOGrsN8XR8iJTJjIc1Gntf/Gf6tdGdUk/XiPXRbWMWgpB9/tO897Ug8dWv7/
frlyKOXPvIMKFz2TF+wyAnVBk7ndHMBsF1GZGX9VyHideosoopJ+U3d4PRk6DG3TuZuBG5wQL0FU
vVL+pOzAbF/7uWgGw6MXxA1mjJIyqdNWar+iOeN3U+mVD45d6M2YhvpuGhtOEZl22MNLTxoaOgBp
2G8jCQmHEwPPs2IGolJGBvmu2bVr9J62JLwOT0O+4CNyG3N4OeM7y5uxLifhKy4yZCUcjkxUzAKh
sZyAvHHggsBbYbd4JMTNmzaMa3j5tJv6RgJs8jeKgabULp9G5e4nnDbbLeXMPHaDNM1E3Wn5VSJq
/9sm2cNpwwJp0zqFVBE4FrDbJ3cu67XrRISbCHEEudBHTM4nEHJzDXA0awPOjiaYn7AsIdjjKSCv
SAd1RwHkeUjbFnCNBqSdPjdZJigV/AGvKovnGvV4/X14lcPL6mw4D3MgeS1K52BvDBC91FgNrjhN
bXMbRI/oBqBbNTyNU4K2At/4elOnSR7VVYbrfDJzlfQAOWNHrEaBpgfAFZUKJttpDCQKT3iva/sO
fNf4i/za6rP23kvJnwm1+1rtctcUN9eO6u6a3+8ucsmPDMYtFSEhEhNdFumGCxxsBy0eDodHdhaJ
7r5eRCc3GpOepRd0tpqnGRmCtv0y9QbHSrPd/8Nilz4JXGxR5nWzrUfR+nLcMIER8GmaNh49hLZy
484jvFIl3StnJ4x0wUJVRLgxTYnIhPQueh4TdRQ3O8txYFGKA8HmM/AMzHYfulntxeceFJGIqaC1
4YdryCthJn67YdV/1Vc+vBKxFyIt7dfPhbJvw/ly3daZQ6SFUWriFcNQLRDBOo+9ku1c8lEALT78
uUR+cXlg32JaPPfk8HqUs0Wgmsjr8dnVvXnx71i5Ph+zpCZVOR7e3MP2w6H1PPdjIIN7ixl3pZ5h
LIquBDAElUsWQG41asxbQ7e2bWsNZH9VKv2jGyhH3I/PlDseVfEC2+TItZt8jED8Yz1G5NAPtTrc
ZUBdngHxHu8AVyD/mASJHzGNk9xoDE+EfsTVozOM28ZALY1zTcNJs/fNWqwS52607XjSkzf7v1Ev
2NWiNx654KiVbz6kQPXWgUyJkw/9YlyeAXWqI67ao3fMEW8AsIwJmGvyq5zE4P6zWjDLeFT3mDfQ
bvAYL625xQ/4o7aDUwSfM+Vmv1mEatVBjG9rc8nNV/n3BOw2yK6+DDNuWSO7l/Z2Vm29AtSqBBZv
4d7wavjQHxNI/XA4e2/98FAmAr+iVBCzDLa0Iqjbe61ENdDidBHT+P8R/vfN6caIVkIYx49RMkWp
SufMEPrgGw/euDkLGPO8rZB+4HK9gHgEbu2jN3x9YM92L4jn9cj7WtwPVMQFAR5sg2Q/ZzduYsNL
wPDwR6QcYYrXWo07uMmsdpKskh9QOtnQlb/EW19jbRswqksHAxyo/e9GtrwhSPKdGBAvXunmXUaV
BoK8EhNTz1K1Ri9zfe0ODYdqzYwTb9etkAGkbll3TQJhMc7Jz5qmh3o5+XElYKhZyEb2qe1rFFka
WnO7iiEuO7NSf9AYQWFsqUL5hy1mAH434FNQgN5qxdg0stk58RKvmz8aFDuzd5Yi2Z5auvI0fGWk
zDcM6eqvqMqrnx3OtMcxFwPCgmVgC71ImFgwO1zP4BbimyHDy0SAs9gOywqqAMCZIHDoF+8Kglcb
WGp6bBIupNRGvnF9Unpwzltdr89xdbinc5XLerUKjGP9iLyJ6H15SChYWtct3r/19bUDiwZUozX+
RV1KnNth5wgaUxbiijI5eY1MwIiOfYkwyV7XhuccUeeIYjlLU54JMnmjGpG08WxhcV8H7GtzFsEd
d3/pPkhKHU5vVaMzsT52R6tmO/FXL3Bj7oPZKZTGAs18q47+GhZg447der4GcvLTSsf1KDpwjBAg
Gw5cr7ihzCWRxlKrOofnnQitzP+ou+Ca9gmZXnTcZdny68ZEN+IhaVDEG5jnwhEXEe8cShFeRF5b
5Gz4c39PaddhvYLZR84AmOGDzIYIE1nukaucBCM6Q6Psxbtx5TJTFq18d9v3iTDnPkchNjY2rxUT
fxTMbsFQC4whN7vQZVKG422iVHVo9rlAIMdS4SVPrxSVmeML3oLZ5BCEaVAaRToPQZwFZdQLJcmH
wZJxqlXPutDlcLwiRBPJeBqKNPczIWQAVqyKUr72VP8cN8cwdUDQxQlv0rTWPSZTcCm31H2la166
wDaVt3yFJryYCFternEqDxe8S4JLTJABOoimvaMWjFm2Yco0BgEtLA2TTzi1qgTvBKrf7hhlGCWD
Dnf4qNZd4DisB5HM4X9JklgBawwghVotTQqKAU8AVlKHgbtUyi9lcKxU6i0H/neliLw9dl/mjwBl
CPw+BfKZeF3286tiMkMOTvMN0hB06GwPcBAepba9ZTJfwxoDz9SQY6wYA5c3qromebI2SqYDqMMo
0Y3WBHKMEEhkPTHJL/wYhxzSGRcGgHxGlID4Egm0ZZyy5Y6c5ZI6tMZlXX2XVTpaaSFo3VndvBBv
w6KoxF1n2uOGI1W4MQf8prZ69bROXY0hC2bsUXiko5mtiJJia/CgldQzesOlNm9HBY7IcwwZqV8N
fFnl1GzHJxAfompU9wLTuq10rQ9YigiImrH3kk4hcuB8p8t+TjL41/em4SO+vxb+oQPS4qBiD1O/
0nerTUDh7UQ3n9JE2ZDOWWf+P32hIaKGZ+CEkNz62V/XmkilUFgjaydOmc/S4Fl9wpFcoZs8E8Q4
JKqiBQ09Vae57f+6mw5OkjHlSWwB2/6IXUkY7qdR7LppnW9hmmSwhdEwSpVPp85r6a/Ko/nkDKAD
/yF2a++OmQ0I/1NxNQgBt/iVBDYp9pPrNskP/3zYIBz8EKMkpBfXjae11QbLbDJXxcWxrWa/8gzn
nNUaQ+S/yCplAyZdCiZB2EnonoPQNSIlARlefkrg9L7Blfiw/EWI8CasXQDAegykBnMck+M+pR5u
ZNEYTWcEJCU7sRFAX7AEhauDdvnRGt4yfYPFJXiihwT/BIEWYPpFGpVItApKhWR51WwcblgTtX6Z
nHKDLzxLEpASnODNe6Se1hxnh6kH5pTLiOWANIzZCEmUTlv3rYlNr31+L9qLrLlx+7VSq7sBkK7J
BKgnLDyqaS2N+vTnS+iZDZNg6ZX+vQH+5+gSpJ6RyTlJkegBL/mTIZndfccvjBfztiAQIv7S6Khj
r7x35Z5FFH7VMkoeSISYk9kH5xy5si8Og/6FF8NyGD8MlfgpoC2zxn3jB3gjQG5Fdlaux5NohVN8
Oz6cScDu8nOS4akwUDyBGySEo1OAzId8npmzOveE0ePndGhoglBNVz7aJH6dj1VJ3qdUF9d/9tsn
on292HwtxnP155SiFDB3pPeELldTgO2Iiyl2oWQhqfNE7sIQjzqJBdngpAXz6I0YTaJx82y1j7mI
hFkyuVg4X4EpTZA4BdW72pACaKdbCQvunxDZgP17JgzznEZBpVP8ue+eW2J3Ca3N2whvY8OZkJ6X
tL6fehtPrRrfuZPvbJCRvUrJvqgLzPIFKjbgFDKe39Ndiqgtvm7eENEhzs31PxiAISVFa4bCR5lD
RaYtgkkAXlN9YzZikDpgKRlBPJZcSBhkK2caTENmXjui0O0nd/9o1giFtaoFrfkqFxe5JZE90B+Z
3eGDr8gSANAFjbl7cNHvLkmPkj2ZL6jHRpsls4waCbVPzsnzYt0tKUPd1ybmjQvetNbCQMmojAhy
acu2opaVWPwSaxXQ75OaRQL+tiuXqrOk34e0SKPygGiybg1iRRJGLWg5Vwbq91Wx/VMkDr4LY2df
CwQmG1KuR9AEjzR+MG9UQqFNx5819Lno1m051tQQ+xC8beLrwf1AOcfy18l/icpVonEWCY2GgIjU
WjzFd25wgx0E8KgVxaiESaio6wyPFE4IfqlGivmfE1c0TJYSVzB+nVg1BZB1hXOU7LDOkNdtwh1k
pkm+GIsDXruI8XPFaKCByF8qddeSlUnqN+91sA8eYOioTOKNJnP5uGovJnkHSvlfJt7RVBuXK0yR
oRFlKR7p7jK3OwUEvsQwuzGtKPjTRohwg/JRa5dJBcuMAbfImNGhNRhwzQvjJHLdirfJ70LSJHDV
62isadK7/e3diT7Jhpjsiuu/W9JZKW106zZy5KJH+at7SG744CClamH1rv6DuXVYhBProQAwOlP7
pJ85cXnzXl8+MyQt6BTj4jhcHVLDc4tNkFkvrfb8pfJWPcoN8i0E5wh2Qg1MBkNbkDw6I5plUZIZ
zk0NQ+VeHLQeefLdQGY8D3pw+SZVxj2LxU//MEXo04sOcAkbzlToAakYwMFSWnP7RmlNIKlxZ4JB
zc+6TGKCm2poyw0g2x0VZKmRoA9JDo2O723hK90Li8A61wEHganULeFJTi/VtyfK0IlpQCL9HjF+
xFzTwyO1Eva8yFDHhHu+/ADvjt4kS5JX+5PU5q3YhXVFGdNkUuk7ewnDs4FxxIAj6J/YxY4PfA7Q
GLf+9sC3jwiqoNJJ9Pw7C/5BDXlJ9oEPdEVdpjsWgIdRt8MssqvhyHFDaPebvalYf5J+a6xHVerx
bOyelN1ynRrJHjV3KkAXMLxs/FnQwBq0zOI0F+RLXhvFQHm/mDpfmPnvNyf6LUYa1RwMELFQxXeB
6Kudv1qt4yYpcscJqWKO3yj3R6pG8/UnJiVxSdDGRyiQU5Sr3hvJfIsYxVDgItSxiIJ4G2L3j8Ms
DeR4zCZ9bTDcuOKIckEQFmo2Ml02TH3LYDodTVADbwCPGClAPAvcnrKgy32BZrgRKW9JywdMrnPP
m9hUUxJk8KM2LZ05gvjW+BGIisG7UF4SnY3ifh2bdaE7dR7Cc47Q+UvUT5VoKNZOjE4mKui3GZje
IofZibplihmGsrBLWCH+gUiRFsUg3jxReVdnJnh3zrMej5AmL8erpzPJdmVtMFNQSsqX4kDUF9+d
/3/Y2kaSUcEdokAIW2qZkTseDV4qh2tsvNlMhe5ZB08SIQklSP1cVswf7gZgBq3WMsEWyBBZuN0h
mp0VuD41vloTSikKLf5GYGaaEbnY2kTvqCDYAWsZMwbCsBnHIQ6pgZMUKJOEstwKfR+CFM4BBqUe
8wfl+X6OFFH1/85AVUNgEqjuJAAZbUjz95bNnPBU/oVInIAIdgHiSzUq65iN36vzWH41NQ6kr4UH
51w8idWAe0JY0QGmN1cFmSm6DbQFcPXPnkzaIQJt1DeH/ppRt9RSFF8tTqEXVD34X7Z7po79K0db
I7swff9BU/tv7pcVupZd69Lt08XaCKfnsq5x565XM/MMzlCVy08RzU6rJAfWNGGtrjWoq7sCC9t8
fWOv8818AxED45VP2JbANz8albUW95M+YNsD6BKrLqEnhhCcqHlhGF+k8s651iZkAbOXBEvHJmku
UOdz27LJcdd/G3PNssgPv0RDjbSYZu6zafioPaaDmNdoRfF10DaiR6yM6n+Tze5CSJKS77aGvlSk
HWRNMadC93kSfc3223FgL7C++f0LW9YJJctu29fdHAUnxvGsVBU/JM8ETStU0A5xcqwdGTSPAYdc
xgnrbydN8P5cNscAtCJj9W54nj1ZrUNWzSBuxCpp3DJ/dg2fbuhgKJuRvQm3q49E1jgD1mTJOQw7
wjIGf+Oxl3r/SfzpTLpg13Xaw40Z/h3L77KiBPou+PKJEqaYO0ACYYC32sKajGcv48IrSi99Kkey
HI8mq8VW94fTbzJZ64TH7UNDfD226rR0kRo8oR19pHpUT4O0Xeb18KUGVQgsvY4O0YWZOF9F6Mc5
tyiikHhPi70nkU6ILKx3qRVPDbPD5j6py31fU7ui3Qzi0O7F94iboxoAUchWxIrZBKW0eX+AFMGG
GJccB/hVDNDEwqemrPZikxQ40sUhiuZ1RO2+Bv4dklVxHQOS4YpTQYJIXK+cOIiKxXXu5KTZnjBE
il47fQfO87cZkPO4hSUKUs2YvXgNyFlpZsgAxILNMfue/SbPdAKZkZ8kWpnBILY6SMUvWEK0rEYm
5rDPik+c35j9YVjesS+xkBLHjkiv4fPOUtz4WsHM9KGTAIVnPWBUtgV1Hekr3eiq+raI14iUsvJU
Pzv+gDOcgLBO4JuFLXK3HwLfMWEOeqogKIRjHTVnChgCxxIXcMHGpm9Sl68nWNDocYjSgAMtiLnJ
02BwjtBQJ5tGGr4/CX32GFB8W0K+urk7WtPGpFNBwJY+0ekoFSeJcCMOezmn6RTnAjp8gcKnJC07
8mAWBhl8lJckxguQYV35RfQZul3riB8NYpe0+DKvJtMpH3MrWXWxZHpGLeIfs9x8kl4j1pna3JvV
cq0dIUQNdS0joGofsHNHECtk+n0KZ9CPylFxqKMIZWCTcE2g3QIVCyThkvDQEdPukIhN66gAI4gO
i4eq6w2jnKKtPDXx/JNfW3nBr+2Pt5Tn7pE7MKVIjI0lVejlbwn51wDr0TincW3y8JKNV+BxAs6H
Z1kMouEkON7qwNwvCjfu69mJpB3WQKsJ5LWDZdSdyYZg6UEp4ATUUBWhXOGwzo1b0iDRg5pAZs/a
AjoljsXFZdjosDS1RPwsVpOEiBLaR58Ez72YRuRo9RdfyAw3yE46zGWyDlFOGDEkTG44IaK8j9ZK
TtEgIxOQA2SvO+oTVWGxUuiTSGQgIouw9nGgj35c1xCXgWiaHBmwcZCpVZXBQV2obHg/JVx8BkPA
vi+9LRDBWlCTgkLAMZrjH3CW0J1cL/P2HANmPZxLVG1TpOWjH756uWyo9lofcGwTXJNJTwjq90fT
P768GGoCC67YRLjIFXt0FE3LZvnvMBeiontXnMPh7e5NjTK40mH2Z4AK7zRkdEwr+F2Sq7H2CeJ6
yqgdzZ3hE0hc29OZIm2HDTSHpcTFRK1Quq6CrRJFHivVtXTXygw3E3BxH2IbvsqGTmbWrDsVntG0
ge5Toas2hfIRo7C3Xq/t2udv05PWj7TrYj9PERgSH9oTKbhLcA5Aalf5JEFvrdqMYvQnUhAHxtY8
7X2A9iyBDrxWbQ+dguaZrEJwD0i84T3ZHnZXz4SphxjB04GYDRiqi+5DVnn5e4k6vXdnkVm8KGzH
nM6gnvgsVQZJt50xWWPL43IIEXPSkHhGJWxDy1ZwV5gpMZpfRBn3ioHVc948fkb/rSMWyEZUmRYu
t0/X4ulUx7lEl9boO+jkXJADpxEDcVchvQ6RyCVY3riPk8s2i9fOWWxAGkQdCzZtBcfAa0feLXF9
Yn6fO741qHMQ5sUrngTKcJXF+Sz712bogElCVe808uQYeS5bhya+OPt0H3ybBgqV6jJx44Vnl79P
IISgktYfhGQ7tbzX2uRDHJtdq+CaUHH1BdeoSM33S3wQG8fma8w6z9Gq+TEfmVVD6s7Qvmd7jAi/
0Wq5eR/0L43pthLDUd9FSvBugiNuvO5DMVxzRAIizOwu0mw0E0FSrKFKT3PB/Y0820lgNWPhH2t9
UOHxi862eiG4LPl6vSO6mxSrA3FnJ+sZEpUBmetKtaMbCu8N6RW+FasdLapoKiQDKIZ9TxIHdr89
Skl15VcvMKnTVbbENvTiagP8GUjyJ/nt2PSF7BE0Yg0HalHAUVqSAvN9bpD9nv7kBH9yskp3sKLq
M3ERJ7xcP4jOQR9ZKY/y0LvfzbG4BV6WIFNNcU3Bknv8yzFQtBjYiBRD7qBgM8ArndzV8brZrkAy
NVvlnKa/PLb68pPI6PL6vdXvP+PFnU5DLneCGn0q08HkW/wzymqf3y+z7au0fdSfggx3BrnXB3Zu
tHrIc0yD1VrQZtDf0D8oauDu9fkBryV+NgiRwg7nHageTUmtAZ0q7ozFZMwuk+9BdZvozShDBNrZ
FateSUqFbK7vMtP3/gXOlCnjggGVo1oWKMIN/DyXU67kDiHjESGDZ6wdbPYmBzLHudbRj8PKhZqY
WuBsdK9iwD/TDCZb64NcmQqTpOCAgkbBwQsiFV/Bz/N342WJ9qixqZiAotgqoa8ecMswMZ+sE42q
s6dTKMdTChr2nKAa7hAVeefqQSQ4SIMi2oT3S7yzKB1h3RI2qZX0R/XtCpk6ZTlbV1r0qTFjYQyw
kIE8T6uTVWwhcPrBImzZo06bhV3NFwrKwcz0remwoHKt7yTt40zk8HJEmYywLvol+bGM/dLVTMuw
DDR68Yi5BfV9KZgS0ORic56Kzll81pS3eCE5Mx+EN0wlY1P1FT+tDVpZSoLK2bYqKHL8TPfPihnr
vsLFlNUIKI2uTQG+QYsqaGppKJg63RdeemDZKeO2LnvXseeNdHRUxC0mS5/bH1W3QCC0G39ccCqD
gxQdxdDp/rYoIcZZaKLp78hw89bx0mCiws4cJy63GcQnBz1FAHMTxfsroK+vcl9FZGL04l2OxnbI
+r+UZ3GYrJIoqMeMi4epq16JxdxiNL4i5bFyMPSEOk6w6h60buC3/0szJInByWSkbfBzysE2XugA
6gNHCN+lzmEgr+zGrvTd5nRQtXKYGxliHdWH2P9CzRlb+2nkQJ8lFDVjD3csAwiro/DniDRDW/yG
VVphPXv8wYiiOHsnA3UB1sDlknTPQICHMImosTsTnvVXl09Yr+9J6Oirt2ev8E99woO2kEnFGcvN
NpFBkMrkJmm1/VUhdhTaePDNv/1o/K1pCreJ8IqUAFOyVIsag7Oc105BsWjomZzAIUP1xvCWTMk8
NMU8iJCkmT+BRavvpZ+K4G1BJs3oRWZXvaISFrHk52kpRrlLPmEATAX4v4KE6to7Nup2pHpSZXen
FH4fxSljiOXxMUieAzyPo2r4RLO/vp38zWwlvKLXohwvHNsr+NnS2EEuIX7Yq8rwlM6OQJvaedtY
XppYC53rI7CnPeTUqbbQyCoycKvKw6rw/WEPYNHMs3sxL95tbc1VAlgX0zzxkzIfM5XlapruP0SQ
iUQfaG0OtMYQoNz6Ai3THuVrgUH066FUaJa/W5jmHEUKnDqfpt8vqc0cC+fGiv7tU1xW9+prd1so
3bF+1fGJenQPtVLsRZGRj+9GBX6sOzdgtmar/l08FkKDslwrldrFJ9w14YwiCAsRWIWqKZNZRw15
QU9JcagQp2iwQNWblwoVfrUfD1mwVcGx4CyanMWJkYTFi5lPhpkSIyhM0x1VnMmZpkOGQJkUXPoB
llQjqCCzWaoQ1wP0cOpSuDB4CtfRHNJ6sdaWtfribqj84TsrnSRcBTrHGbE4ugN0okKE9YFY8IBn
wayoXLr90PeDDzZhaEtoxIzH2cdXN2bnvWG2Rkiq675+owosqOZyqLvoqIaUMn6pow7b7RgDBgZm
LJoTLjZS5exgquOwIXwkk19Jq8RPT7+Xt2RW+hfACT7mCQhYp018zFNYZF4K7hteH6/MJcE8uGfe
WUS5UH3g5lLg2QLORMPryoTquM4T2ykEjUgSMqIvTuYki2b3U796DgNBme7pikvMgAFELLuPu/z1
GtWKPGwIv2ZHqV/kJaJdTzyPzUBAUZf8j1XL3LYBJCrAEX7ZTcuVyuQDz4wK/S4ty/sQIdqcrb3P
1mlmQkWu/54Ivopr/QKuGsQPcIbFbOeFh2onK+YejvccWn+8FIVDaab6Qn5JAIGqpgtjuyzMpT/g
BJIbiWytgePqumPfZ0+dn3RoY+0Hp74a4rzSEkZttUtxXzSyJaXPrQXa2aIA8BwYJwP6InXajKcA
vaccLg1GIgaSdytUcRbFcZ8mQKPLHoZ0Ld8fft5UUEYkeyvOzlE2nlx+IZpuaiXVdR3FeT/uF7Cb
HhYi89Sokk9OrpIPNnUqWVEZp6zJGpzUhkbl5JLiEV3RhudwXxzfmXKFaOWehq4ohOoVM6TfC7sU
vDGdvOHY6rIL3WhqVm0x/A38dTo4Pohw7Q+52JX67u9a3k+2WWvQ2K8uqJCuPTd6XBBUC+/v/lJl
oEY+dB+p6u+GxAWDaAQlkgazIQXdJtWVG+00sJlwL0k3UvdIQoRn8IaR2twAu7HKWZ1GCK6MOGuY
8CDp+F/MA0oDqj7A7HnjYoixDDwAPWXnoy0dUovV1WwOT9ZZcxWff53EzpiRbC8LDw9RjRLu7uHn
A4nNwikIGEHfPg79r1ckKRM/3vfPOS0Rkd6d4uviw4HPlJfXlYKfA7fvj+22Ar0GUKMnGnFWzpXl
EfZVe5Hl/EYrSLonugfNqZOUKf43ruOKwcoamuuBiuvTXsftsVwiok120fzkLoSK1iZl+5jpsgst
EoE1VLaZKdq3A0bYRRWXFlLDeOQvSK6XYYarYsnLY4lufR8j8eNWfecLXm17lIJky1SN+o7UH1Vx
Ltb7o0qN65chqXFWPFO6zOKjJrshDrdfNQeeAlcZ7UY2Kz2ull+vW593KxCJoMiA71AwmYwrKIxg
HVk7Ki2Qtqpm/n1Xi5X8P3i7d50p8d858DtcLKByMEXvbJfltTAPuLL9poqxpD3t7cXgXxTRPfZP
EZEeFgTmQIg02QUnMojxm17bwtCBfCGfZA7sTPOlxWkVC9X7IKnCrgnIzzq8JKMQRQbpgpEeFD9t
oNqHRCgqMpCKKzNwR5zwQ0y0KTwxlvQsjzxx6RVwpScrsjFLMBHH2tVPPuWDsj24dDMlg1sh4Hmm
umb4ZEquC8SnmDZ0Cr7sWLObrviCFqpMi5YL6SS997ItQgf0xexzEDSKdfFZEcc36tYt8MbaXJmF
W9zQwMW6rb8kbeO5b9odtL+xNvWosByY0FOAw6hCGJefaRqI2L6dSvmT/zQAdtmlc42J4qLP7Sm/
RhHh60DtZwiGyjDIDUR7uMHd8tytMwUvnrmeZW8BvNMBYCaTUHe2l0IjQo815ZZA2fkv5iEokwmU
2g9NHXAF72rHF6dzwxJ3kI0nfqJ/0dn1CaSNPRqzTHh5Jwt/tgoAWGVbqCivuDnzHQh14S1V75xw
M7jIvJB2xqxPNqW02aDFfzzDw3uUAmgYphLL+CnlRTdZupN1O5AHtQio2ho6Nvo42YUsLTe8YEyO
laLdtn8nQOOZUr0ZWj8iGxL9bzgcZbbPnCchlf/nkuMmXSvFNar3feTQbZfY/tCV+8H1qq78Oc61
SpnswUy+uAVoSx+hiHtNsfQfi7lkh7Z0kZE3I8/esU2crmzGYn/8vKpdpmKggOxkhwrUafmw2/ti
pPdozL1MvB36a/z9ujqZpghIOz8TvvIaUEc4LxuQpGAYf1HyIdkLqidEgv3iITdeXV1Zv2X7ArUh
HtNmfKyKZEA5LT+93uLBYI/omAsBUmcU6BcCCUUkTnES3vB4cgb4mZh/OTx2YKJrrcWtpTrEkTYt
q5ZeC+QQHrWDRhY/PAb+KYRucYP8/DpHdEmDQ4AtzU/DhkLzwU4aXBWUHV4RKPfOBeDrIAYcGcmq
ItykpCsXZTzB1pyctnWmpB/kFGy6XBj0/r1san76y9v3VpfTlA8/aG6lmzEl1mW0+okfjJ3HFlAJ
q98ouNseTlIKeGmnTiOwzLoHk5MqQgvrxGzXaLZI5IMWJi3GghlKBcAymIJyUYgECjrFNjBiLt00
xTvfmnQD8hiczNx0LHui1fRGi10rQ643N1Ws4VrZ4QMP/43PsMKaN1TJYZtMXc6jRPhx5A2mkBQ6
jiFymnK3gXtzCGoo+b99Du8WTm8rLMgv3oShetG+4xdw6DeM+rHLcsWiMaSuDTbDsIda7NOxWK2U
o/Ghu1gVhZtFUwUQCjORnQJp6V3G7eu501KA+6Bp/P6TToghUPjUrsEoIIiGhU2lHdnbPfUiYCeo
ylYrnoTm6opC0leWNHR6p3W2ldUkv5Lc5uE0Ixwu9yKiK/Eg8si83bvyMck+fmBYfr+/fc/H6nhO
pC+dkJQjK0gwoGBezNTpKu0j75HL75pm906YKvepB9Tn8RL8W9e+DFggOqDg7LBSqNzGUgIpD8Ge
/Iub32BFnstOQqOJc8kwxFYgc7Ns5JSogP9PThgram4iqjx7D/Wzf5aiPoS004MibJewQ1S6VmmL
yLrqD/lXng0+ZBYfo8JLiz0Gf24uCbeYEKoMusCAL7NdwEqDIW0TMZbcD8orM/IzZj5K5KvjfWqa
wymjqfBPZ8Jq7DOxuTe1XqHs9ZFaJwyNiLxCRjomM4iwlJeUGTkXefRvsRmIPfUH+qSMA0SHqDKl
4MbvoewzS23Utd+wnk+1vGUyNNro2SA4oSqFayuTDDfmlAVfX7lxDxWibjt4cJWb8dBwNwzTIb8r
Ymp35I40CgAvofYp17h4rqGKHBWdd3Y7YPKIYqRfwxfA3Q66oyX/Rzuo5Ze1Jukf924owZoL+3MY
nlpQ0VVivmYl3jPrRPlT/yNeQxroav6bGAPFmtkf3BBUTh++XhfrU5MsriDI+tYLBfgfxKm1dwEN
aHxcYFlM7vpj3DUGqABE3Mej+ZIg5/S0LD695Bs5ijn/+HkYqA/ld4/oHiieScoERiI1kxAdbeoX
wiJDyCicj9nolKxJMPzu8pFxHnqG3Ouytx3RDbhgz6Lcn6S/K4MX3IslGVUrxbo5DMWp4aef7ujb
B+R9iUNz8aHfp5bFH5QksnIySt7jAIfl09kNNgsu5yqneXFnMUfsm2LoH9iiYwZ8QYTcu7gX9eqj
qPomdkhE+fdjftaBBVXK0hy5NnDCSCDtASIAio4rr5ZHnwmQ1nm6C5kC9lYEXfuNwUjmaGjKzl77
JW29ScNuFcyZ9tX9URjU/WBdHJPaFA88pOW5rZov7TpeA2jILWDPnuiq9xGG+aEXp4hZYw2t0jvn
16/W5oeIyvSYnN5YONn6sNfEoSej9+AICRNKiNB904Pv3CMwULY5eaGg+BkaZhJT7ppZ/RwUSwkb
BzDRVaUeX6sJGLzidlvLF9gqG3+WHnqKiqLSxQdNovsLSo0VGjVQQBfGp2raOHf+HlQ8014FWsWy
G2JEql+W6k5lZcFHbYaA84aZUnnktfY8z8UnHfSSkYRS9FhCzNtcisWiylH/NkLmIQtXdWrA4MpY
aeDhtpkAPcONu4LrGbIOHW1p7Z9QuHiaL+lkN2kGyiIwyteLECmZQMQx387NJnnXd7DFMchaq0Oa
nsVQBU73iiE0QXelCJz5ra21qsohQnBbeoKOQO5XA5nRwxChTaaS2jp5Bj7desbOXs9+2Q+mwApD
UkokepwuIyxPOFvDh2FfkPa767J35eiPH/IpBIletrL/WrOSUJ5FwMRyvQUyfMWjCsVif/nsFI0R
18WEi4cHgIrQNskCpmuwCqOwIQ/6D9RlPLPa+Jfa6FT9na5ND834hHu4C0zdfSkWrFbVwRS7+dk5
cYrTmAWmH1sliM+D3q9EIIlqcGyCznE74yLH4s2Op7aCsduCEc5HEMFxW85izeIdZiAasPVF7MYq
MxfIwiF23A6ZbNDAtDezu+Q2pj4oh/iyhE08QVQLKmVBfjczovHqe3q7p8zwUNtzxQYSmTGMmQY+
RnCz4aLbvfmm1SYMfU5B577IRu805sG/8kJjUWJR82L6liYn2c6IbvGjsn4jKVhurOSOK4nthZNN
0e5WXu9r6x5DaXnRxXNFMjVmqvNgG2Qur6viiHGvROlFtg1sTofFW8OvBTvpbKrKC6FZnGU4Rxwa
78H5xQHYHXt6RxcrLlMh4SI6MXHlFkq75nqxN5dpeA665Gm4QZttQXQGVXpSZBgrjYTXPc2AN/x4
mI3Bbe/cOZ2I/vAwA1bL87Ff1BhjoImUr4J6eCnRxrtC1cGqXSL/E4eAYmKofhoIoujKgn3/URQ8
2AeT03rF2KOQWElBCJzGvm6G/AHb5LFE1tmlVwpktQu+Mjfuc1Y5IubS7Oz5eTETt4zwL8brqhmG
6DbgVUpzPoaBKyoXUOknRb6fCF6shippZnbCdyHa4x5SH7rLtch8792ngvlrVJzQvcV5dSNenekg
vKWzjWFWhukfIf/XGn6MqZWfLV2OcIEnmcNykL1syVvM6oh2YMjRYKO3ffq7z69jliQZN/nRakxN
W33ALZKFa6hO0QFpTTmRwoRSGGc0hmuyXwF6HpJfLETpPKSAkfZ3HyW7xs5dnwKEB0AYN3m0Wcff
GrWifFv9XlP9XXD/cYKny01IgAeaI2mbnbXLqjiWXZJBPwx9qNJz2nZRxwgutb4nqNuzNn8WePBN
JRt11N+elSCKjNx6Yl5ycij83pK4xPX/wysnIdYYffqkckWQedSoB+/6qXepiAJZDPJpE3ZcOXJx
Y0tpWkDtOXtxPKwMwM4tNl3RUMHHfN0TcP8qEmdqTPlkQ6nE0maLrQfG5z61DeHHe9fhx89QVQta
dFlnjeP8S7YO42GJsh3mpDAfkyV5fRzvueG0w+bEE+vjbb58YqsjOj6GMcXqvn+WLR6OQpNU30/H
P02fd1TcYdPKQofebB2yrDQKa42EkknvW1I0rLqu0dTksSIFHcHlRSWbVg+zGJaCeA0fx3TipcZ6
zLUZKiPr1sdCZnRIXz8rN1Q2SBoNFK7l6EZ4l5IvU5/iF0f+8hXISlsdEkvGrKLJF6RyrrgFcZfR
n6dvF001fgefeEVF/52kjYJMv8/Z7IJL4TgoZhhzra3ksQL/m8q8cm1/lfZfn8ZSprBI3JA7eh9J
Qy7cMUsdPhGzMkZOvzTPhmzW+6T2bUf9xV4aI4ShFf2YWvLYlGWPedBLT012e5SVd1LDINQSxDnD
nUE3PAu5oyrc7ltQUoLAYLeDJzUyRPxRgUewmUV8bsoHNkv5fps11mVY8iackNKQfyloUccXD+Lk
69R5cZqACeZP5LxwXSGmRuZ5QsXU5Jp4XoPlBL5+vFNWiwJf7B8sDCdgbmuVrtOmNuEpE4I8JgKW
tkp7l3tLQnz/PcPQy84p5901D4haZD4yg2HiDOoGKGF7qryURaddWoOl9g2E/ZenkDpTt4VWNhn0
Qhn/AHBeR+seadL2FzfEwziuBOBlcFk30KpQT67fSwiCqDNy+WHbSBUm4OIl20TU/dy6EFBqoC6I
fHJvMnU6BVHrZfuxtlwZo0dgeObNSl9UUbenBgnOrpNzZxE4+C3q1vlUeUaLrR2kISFOS15rZbAf
4pBQI7kTXEEM1pMR86JUM2MOR5jINZFmVMt0/Po1dv0nK8886G/wFCUgkhQ9OYuq6P6Gb2O7ufyx
1mVikRfdLS0meD3zwI6ZxVIvRGmocDXkNWwv5IY4zSFdmQc8qSXpUwmryF9/B6wcrNTNwOJzneZZ
B3QcDGdWNzuMtw5SUmtyeoZNuO2iNL7aStM/MRyjwB+kSPtB7+pT3LWJrAyyv8QCtYrOS1runtUZ
sizmfFHlcRpv5ZlGdVHjZhUfneaGt1QKBV2+yED7cDFwKu8f+5CN7pIs46LFMvhlr2eJJP3WcU+z
mzxjfQsRmrQ0pgKzHESG5xUGGDu69FfjVOckDpXmP6qd9EqOze1tpT27ELw/U//4u+pvPgd4FRmz
869l43dwqtt6BNQ/stvDTioSOD/Z51ZzIGRIbT/79TwnCZsNn0cZPk5tEFeuzjve4DYa9PCaPaUE
xxiQGFMURRKPWyO7l9YvxbSzITDqYbpVVCIlj1lLEh0yIpifJNz5OqvQUyKxPSEsSTgJv2620L8B
xaWa7Om9MpkpjBWm1SuaztJmGsLU62Y1Gi07O1Yl2hyx6OAZgh6vAJ6qWF/3ArP2wy+KRfEgpw/0
pBk0XpjjaZB1iz0gDRI7e3y8gdma1R078xgLumiunavxKnCTGZdRu6gm5fqcaiAVnFqBSDliXHTv
EsiUtUi1yWeWR7uuyUeOMIFnOAC04bjtXa4bXz85w16HjVVPqddwcv1my+CRHLw3aXX/UC5VoiGY
xr7F+iDKlf5aA3a1gDprbtEjjKE/4lJDowZRSMBY43UNCQSYLpqUOAnc9lpzgqyYS0OLvF9d/S+H
RiBr9CUkU5nfeUtt+/tVY84rR1BXs8RRtLw6mOI54peGGyrUbHGMsQ0xUoiq+VTdHL248NeCcY3h
JQcJKE8NE6GWkzth9kkKHO4NiRYrmWsbrQNQE5z2/CHuO8bdWp5ZBLxttbje1162CUo2b4Zs/oVz
kDOj0qv+z5tFTjHu2y4bQIfZFkjeZE0XoKfJrphURpsITc+ZaVl+jvBKtodivjKMtBuYF/0TyuuK
JZFE7SMsd3hrQQA/BbKsDVx87t0STjamQqnvH3qiQmitB6FRmP3WHRBElTc8fwN3VwOer/BjDfXA
3syIK4I88RSnb+WDgEFhAjNrmMDD5+5VtRVqEFcE+mHdUfw+NI304mVYtXVkedAT786IJxNQTo4u
lKApIpWufstE16ls87Z0kn51wPzf0k6P589SZbCJb9nzurDE7VyEqGedreVhubOm0PxPfQvdg1HS
eXVz9g0Bj9tAJCB7czu85uL5RADExEj2ZAQwPBzFFu5rStic8i1E3BFYSrpPJ72c08MmGCg+SGyu
4kWAToj5ydp9swmkhXAFhfi7l+p/G4WoKJCLa25NFU2ISzmpfQdIFlyoMwv3VLXZfWRttZMGyn58
kOmDYf4y1K4WbV5HzTmagMQ8hW4ePJRBHl2qnR25GAKWDkbrTSpfL83gSlLQf7fbPAIeh/jkdGc8
JDlBQ3P1vdnKBDNBZHFqG8UP8Lz3/qcIq7ld8MM+9kCRd4GUedkJCSq8RQ/Su3UrVeeIMSPUSLuZ
L4P0gexkUebB8YCM/Ninp+N+vizr9YKTtyKQKoYuA6uoVdcqddtffhw6z+4O4gDNcYlvY1IbfouV
3A7hyQ2RF3bYVzgOCUQIcFkacLxkj3gnhctXA+S0Uqwv7OflqM6Apw1CIO8ko72bx8ChrE/S0KZk
rJzvtxu3IUc+CjdEewxmoQe/wB/nxoZ4oRwnGIEewN9bugI/KDcl+Yj+D0E3w45iFRx9mO3vBhNs
W+cVfr/bLH6l7bc41jGYBmyb8/drJSu08J9eQP+67sTp/H5UMKOqYLkE77jZIjHK+2/YRsoQ0o4M
JYNrt3h5JrMeZIIvJAewIGmdpb06HpBBJH6QmLh1gJvLcbU4WTwwwuGU53OMm6gDk9TCZVOkCdX5
8ZFsjcELtVoLeg4/VJRhB9jnO6Ui65Yk4QIkpQY0C9/ZWfsQw5Xm3LRxxyG7fEy6TBFmW7ys0y36
NyZNYNX1XnB4+EytkCAxHUc6mLhL0ZSBoosvWJIIUsBKesRj5ZDS0Ay9+zqpK8HFKxFcQCpkv5UU
O8X+EEZiBacj718jiuuJg9OHUm3XjgcG51A6djtosZ9yLPha5fxgGDRRWGusHET/fgYhdvYrlwCj
fat3n2x1yDFuB7qXFHq4//O2yMs6C8miSXO2YEjkphUbsIQNmDVvpUcS8Sa0F4ig+y5DhHcTakrK
1PgVPzLPo1yVt4xwd1DiYBDaHEY4sPsiB+5U75wp8RPbDer4s9aEwqtJNrJMqRiWPYRK1RrellQl
0SEYbBhvpHy8Dj2C2Cn1ALF271RCukeAD5dD71MnDv8RQcXOx3A1PuD3an0uD+6XMYwhSdtrHTSJ
m/o8G3azjtIOaDIBC1QdGsMsUWJLQRy7k39wzmY6Eyk6p/p5s3YwuQl2LDjif0Ivp35UTFxDno9L
hiePIJhYo/vozUynmXk1G55lsuWa6gNV67iekEapjNRLWVI4+bek00+MmW9gIBCW51b+5/Lh7jzY
oJfvwv0C/v4QHc8Z6/8zv3xROvtKyyyPj8Mp08f1DlUCQMbk/tU8lL0eHRu0Y7YQSpHX4t7I2IY1
ea3EzhlLTFS6ky+u9CVwPoEW6lpn7nkbm+51VHCym49cxVZCuEU+ppd2xk1OGEAZ6I3WyG3AONrO
U9x1hnO1LzrNge0vHlm7Fu+/tYJH0tNNcc6HiM/3SJhmYzBwQpzT/e9QszilY9raR8x5JBTzx87+
ng5iIi3+pEMDUESx2RQp4HJt/E9v4e5ea0WMvGzqwaU3t3wNlXgIP0VYylfujqK89XTGckZ6Bnyo
hKmx3TEqUAlwI5Z9I4FX1LT4v0SiJWAm8tFz1epUyHoT3uAUzQODafmxcio850CS3RxgWCYL5CK9
6AInEncpadXEMFEfUaXOJ9nNgEN3Yk264sJ/QpmTfewjbJDbVKdAPz0cNICrDj7uhxATQMJ54mvg
4Nrg9qslrhw7aoTfxQZGOoUx6dATCsyPyhzzd/2d748yjfBdENjR4IJ5tWE3u9HXGWIJMbZ6VZbA
GU6s3NVPJ306ps1qu8Bcn2Uu70LN8CwtbGPzmFgAOmGBJxX5+eGlnjNbRDjlk06lomOLDzDvFU1Q
WBz3MCUFjy8uq9bTOiPZ5qjZINBrHOoWMrRrhIYBiP+5ine6xZWUgfIhfJjAHNvNEx9ZNl0m43sE
RjDKZrBrWy5OsxSaFApHOvCvdqRepUedA6XeO07SW8Fvvkm6MSQkPUjDMGgsjEOtfSFHn92P+eVe
AC4jTMYUlngeUb2uDG2VX9c0VDqzXmbsZFatIM8JVMB68liUToze1jZkmtCVarvVdl79AfM/t00s
zC0ICcLOWtFno8ZLl7l1dOJHjaqtgUk02IySECjKedtsKmcTk5rXo0po2WtIPNqkMURX9NQX66Of
OXyeMkwCX1/r3gFDk5lO86BfrMad3h+vmWAhAEiHclTZdE6mHnNVbgqHDdjUFpWkHHuXjU/1Hw0/
l5OeZ9OmMLgcf5397E5rdr0elcKxA1/SQYNhIiJaQ4moLilDSjvDyLJoUvGMl1ONDQtjmA3bish0
WoUfplZ1H5UYO+ZA45Bbc9Dh4DpUJHprQusaTLrMjbhalZk74XRjdMqzHcN/w5IBlTTJqDJj0WdS
oU0MqZ6padmM2uXiYnSzYgdkQpw78xzFxRSxICtBKZ9UCjDqjszEZH+SVbzNkb1uKvCgqf+Z6my7
4wzkQGNXwKgvDMJ9VV3PihHsavOkbEjjD5Xm8wzOyEmPIXGpfXM1mgjcIngN95wrkqVNUetE9vKK
xzEL1ss2lPmiw5g0K27jDaGC42tGoe56WuMOXwjii0QwvMZGA2ZIpIwtfr0+IEHGyLnrLQoHzZxm
VvkX9zhiGKBqdk69SVqnibYWyloTk+f3EJGKZKUjZq4cfiPYJcgwhzbzPpET8BXABQhXv29xeSZ9
ZPYPEFn6X6oM8h762tGf3veuhvFyAXYobSDP7spcENaSWFcpQN37836LYQbR
`protect end_protected

