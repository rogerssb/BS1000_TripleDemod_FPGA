

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ms/kGAvt+G3oDCnERO1eycJ2b90ZudbNptdHH38L+Y4GQelWq/dBA5+w8lehdDT6+wilefUiETrd
yzOT1V0X6g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ma50tP+5k6PHGNbYhVzuZHTHAlUzrRrURKkQAn10mVQ+0FA+BJrnWXMKGgYaN5PW5jLKRkqwH6f4
+OPU50BZRC9O/gxpvVVAFHL58/d2/vu5JIbeAxandLPAFA00Gkku2vG3jj5JLesjKHuD6dx6X7kt
ltc1Xgv5gMIosw2XoI8=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
V/moDxOKcJZbPbLpE3UFgrzhtYX6V25CwXFIfGfgEujL4kSJhdHeqUaG+J680LW90EXDUJN4mV2Z
+5/J6wwTqHzq82YXHEiFHyVn+UKfS4SgLyuITAeVkbGJ7gYIetF30b5cEhtrK947V6NfEdKEiDzv
+finYCL7sk04MMrJamE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZeR2RtoxAcS+eEvdoEOH6KignhKIkusNMpfM3K8fkH+CyRP8yJGwkrYREoL7pglF8bT4NyO/nnN7
e94uwKTGyQV4b75DhIrvlVZdzQb64e9V7E0Hkp58aVMVrlHLaDoDEzLv2NcufFLAROTHeG70dTuA
psS/MdUEKT4EIWY4kNfxRbIrPwe1NVBMyZm9ANTNsqFv8RztSt8Y9DmcsjQgPXvdjXH7RgOe4UCH
EyqxbXFWetb4BHORSIwRDO/rHW5zc5FMALVjZ5Pb3ST9gzQpNKfcg1d2CmubDXPFLQVhqQllXR4c
DtZJQRQxunJoURUONXMIbEV4nVEEVddf4EkOEA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ta6p2ELMVjppL7BP1tvafGWa96MSBCL/Efwc0X2wpgefM9qftoAke5Hr9CQjRrujaAeRDnx389Xq
ZCNCqwMVw+BU+QtNG7TcRy6KVED2eSkQogAl48DeT4eRRkdOT4/PKwFOYOf26ioPpeJX0KCHBA28
MrYyWDTrtKSlglqzB5lGEQh7MTfAMHZtKzsIZ3dH5/XmiHxWuKotsFMIW7+4vyUqG8iiz1QgQZKa
rKhkzZh66Tw4SaWTtmiFhOWUmAVGaA2ycli9svcdoW4uoRHZmubacxWVrupNeIdSUUZNUKhIUymz
OYtEXLYMKXFPFuJSg6Lf7HSKNTzWZ6gkp8Zgmg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ftAN96inAf8l6/mVEBs0oGDx+TLuDZe/J9VNNs9WygRsayoieIiCpDcxcofMYgCYPhQjxmAueFDa
tr7WJHxy1AtHMXRriEVgahexvtSLFeUKVltgt3NwoM5v9xZdgz9vtzruyMokKiLwg/J7x3DVEPxx
zZGnmoyRfDY+Jz2HpbpFFKridenliFuNkbwh2gGNv82CNMIIVMDFt5la3+s+RmGMgAMPBHhciUp2
iR7N3Uy6PAo0WHs0CynuNPk213K9X0hgntcRbDiFysBjCKRspfRUIa8vLasutwFQ7KbuiaeV7qrG
6GU4yaAXmnAqkTUo49a7KmR7cx1OMdkAGRLlNw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
GRRZxPfhF0jHiQlooY+xh2TIhb0Ih7hmFcDrQIP/vyP1drWBlVrhSdG8gPXU2XzWL1IZJZpOJSCw
P9wobBCS5nEPSI5Crvc4hm5HNT6X+5iVQSsJSnpqvEnBr+uw4YgJ+5hQJ7BhRH/QqfKzGXXGxmy7
RvcPMyMvj/z1fsf78QN4Zf9XOrsK2Y0hQvNh2Rg80mrr7VXXYBCKdEsy6Z/oBTqcLxaxcl6BFz46
0iD1fMJLnr0KppKdka8uM2X8x5FStudJ8nAyTfhuwF5GGCVL2KHi8vsEUqZt2MNzs3DEP5pbCW6v
v546Zu8FNNRIv9tFU8iHUWoqvHSmsTsZ1h5MDC56Mr5pgv9/Xwu5EXDQF7Y4ZfHLMVDE39fdGNZa
rssWWY1jwBL/O0XImTQnIk+mqDnED771ExNFzhsjPCl504oCejOZ1ujgY2KdMApYjRsaeCfG3KmH
ARvF7zMsrdkfl7H5ig/ErNgE/k54vnPzE3ekMnPeld03cSRwuOLj51cC6gGWpj9/VQMjkQChoa/2
rFakhsbo6dkSVedFui9obrNNav0ctNMAQWALmUmvxsBfTXdkzKmHR7rn6l3CCEJ5GFzoFUfIVPKK
kuS5nVOwh3m6Yk4a/WET4Autnojtw4tMiQL6t1lWcmWxsKBNpDGNl6W4UhHWNvg7+1gp/98OZpPV
OuWGzFMpZHaaAx64J3AWdjtryS+izFwOQS9k64Zi4QYKbGhNVgvkyBGotQ+QNxgj+ojBsGAkYXeQ
Xnkgae0ROvf3VOk+XfV9+Jq0bh5L1iYlcsSXpscyfpiNz8cMISpxK6nHP/nKkKIg08OOqYCZPZ9D
UirRhUK74FiDxiSB73sZmYRr4Nm5UtUodWYHatnP7l8tOKIDWNQ5sPQhLDPHlxeEnQCV8yVkqNPZ
kwrlPduHJeO+c3V8L+DELpyHXB26744LUlgjlQCCbZggc6LUp5R2ayy1envwj4O+jNjMFh36Kiub
Id8TDSxTLUK8odAAnxpqMw364jxiy5JNfXTuHQ9rWzptZah/1lk1JDbT2HBqsfUnkH2XCVtx4Wl1
sJlf0J8al7XY5qStt9nkxHFDh/ijcVg4iP0/H7zjZQSFrpz5P/EDj6zfVMUeU6WsRXVqrhyywuoP
xQAAC5c/ZaDpb3n0hFjDLUpb21OQC393WPesBIdLHPuc+rPN1p5XZ5NY3QkPEgD6jLJ8vOkcdTS8
AYL9ZKJTvRQ2RQ+QgewF3unQV4NiF6qNhSNFqWeGyduNMmcDBeuf0BgAFpM49JwCApWKCI0MHtHL
LWM/xxbgqW/V4pJ9bx8D7LR5+Ic0cU9yj8hOIck2PYFF3RxPhcmZ5M9b47knWJrESgUulftN969z
6+/6IyHR7zB1SKLM+ezgxoAidhWa3BYA4MTiCq2guI7WU4VYmjlAblytZsMu4EBqaQ+GRTd3neVh
IHB/wz8Iy8WbQGNMforaRh/SDZxiAa+694b/3ZM/UJqUaP+FkM+b4xOD/OiV98p4z0JrKIO9ygyK
o/JGLKhOO+eMKXVx+jjgjK1f8LR+SwY8iInvbzMbLbeVNZUAnmOB7KqzDyajtA2+zP7CRN9O7juJ
90YnymCuEnWrPesU2i3CUuxWeh6R79DDY3J59BXgcLrgpWHbNhUdC9a5U6/GtjVX/Qz631cP2e78
rp/VuJpCO3CilHn13uoWUDcEe6amFHS29WhzHy6EszKNYgB56GZOqdNbGkGx1aXHC01wGOzB4Ubr
6gGgdVI5+vnkpCHYc4Vzu3GneKfwLxtkyIdiK2I4ezsUrkxM0Yy52d4bsYRWU0PGHplhHbjdfrc1
DRcN30L7F+NNgzV16eSlqcXc49qgJjCrLq622hROvlHfSsli1nKyIVHV80J+nNj7QOVpA5JoSi6l
2jZBULPyfYoUDuMSxq9qfIrgmeSHBnaxsxb7l2vpoYQr53/25sfmKerYBJAQJ3EKT0raHALqaU+s
Tftegp38ntsbHjogd+dLtIMTmlP0QqMC352TlTrXCpoBmBS09nkKfbSETCP4SWpLjg/cS/lYmgp1
fYm+HrtoNiMouSpLSCGn5CU5f4CmWkXtVHrZYCvpKXrIlMn6BuFpm7sUGmg8mGloe0DUc+m7Yy9S
bFJDXvEd3kFidyKU1cWEQJZUBHoFEb2kWC4mPjpQs/Xo4alTHejICV7OdGtN8iIoP0ZzS0krUjdh
jH14g7+aFtUjCCZV1Y3smseWbGOjxkujYntLDHZ0wJ2xjxDi9V3w0lFlmLbnj6pkLrJKy682tzNd
8JmTEvVftaRJ+0oMaDGVwJ0k3zPu1lMnTcxM/XqaYWkV6fG+KdBiAlRD326d5uGewJ7mNQXctpvV
3SyKhaUEJAGmk7N/WC2190t6CoYA/ggjEKoJ/XCl5jXsQiH1sze7Itrmd34KdMLWrgFZVA9GaziU
80x0RLCa61znWOB96bkveltENq78/CMkrCfzGAjmgroplkONf3ixqgUpfSWuXqaD+fSusmG2nBSK
XbgKWE5OAEpxnRrPf687aycilMdXouFk+QLaDe7WvaMDJegHsDFkafgCJIzDtkLA4BsH1I7jaHhq
W5WRdXD3jbuR1NOiYSWgoAEbqo9JB6kQksSyRkRHCEHzAGopKSt/2aluuPhBOohDkp+ajEiv2TpV
yMjUSw87+1K5jN1pOeQV9Ekn3e2hhUu15en/VLRNOW8n1ElOZDRCFHYnEBVyx1AWEk631f3bKQJq
70vU9UbHz+sNMMS9l1Dh1yNEVj4eX2nNrnd6lg0gWuWXk65BncPfFOLjY20qCn0j/DdC+o5LDJLS
s8SsTgT3wbwqhY+EFN5KLGB2+ofOjvpqOO1OASTeVyJZ1ssgmtfwT6O7IKBYmAWD14DSlxz9uiGW
H5rh44OUbmNF3vSr6NvU1Yj0DFa7seVwQCsU8+opZAOe1CspfJ/TV+rJViL8gTPVBLBkVyoSOsiC
Ijte1pFoJhya0aCb1P5GJdBBCJtM53+3t+V8c/Cd9fwPz0J6oCpg3YbKpjdtPw+w+dZ4wqjAsvgS
CcUEv3dhkyfLDnuGZEuXmng39KeRFJ/rJvMgEae1zFttd5P6A0lYIv360VfNc/dcykNFmGEBaUzR
iaCTvtAPFvjDFq+m9OP7Y5F1e9TH1n7oOjTLZbS83+h8pIRWv7UcWNyDA+VlM0Vvu2mV591Z+DYJ
/UJajBgPCgb1vvHv2rC4dI3B9m6b6jH/I8FIlIGpkO2vjgX/HhQKjuGSvNViRqtu8zKYi+1LKTtt
BT9eKT44jMoth4vlaISjNUayimN1xONXhEuCtQZgGynspMHjLJtLaXRK0GIXKbOEGLPRehtyq7i0
0I9B8v8l2CyR+YWuoGKhx9FFdat9e6jn0YVozw3jxsJOW5FLVn0rdVW/Xbk3bk7CuLsTgBtst6N8
4w0Q1wFTuR4t40qbH36zKoqWfn6sROEWPvinaLt7ELgrNlf3kQMc8eKDxq5m1fi0/DsS93JfFxof
mr58nBF6RIKz2k80PnMUMzHfHCSGXSTh8b5TG5yCgEVNGfkF3k3I3+1P/dxDELG9pfbKqEQFCNHu
pT7cPdNpCOquK1QT5V/1N2/syY2dzWcERqwFpqbPzmfbQV3HejTyYcMyU3owaq+qfnWn4545kmrk
pUWh5ajg8WKVoUAbOKy9N+3/EdY8vH/Gjf5ua2xGVP5/jMfbJv1WSqijFk7Gjho1NouNsFznMQ7g
wAOy4GWiOXbU104nG3PctzAQOtl2hCABPcroumPK0ds6B0sBuYiXXFknA6WFmRUX1S5jAH7eQFmS
3kCe/mnBf1f4teLdWVq/8oiIjupapFSeMNvCC0Vnj75Lj/n5LZpIFVG7vHieLScEMi/zvrny11Bx
GuZc4j5rTwYwEGdMSQFQSf7k8VD492zGmTaGm14YDph+OHmBCtbG+zz7NnD27tBrPkBpf0cfRL4h
jciUPsxoHzK7W2ufRBSERptnew8Qnh3OwdLnOjcdeanNP4OzWG1u3LN/db6lc4Gx7QbZujCYU0Rs
cjpdLRe/Z0gJH4/KBZG8CGIdsy40abJcm1v8Xk6mrb/94/pNAJPimPdrdTnyZTgfIXmMp5qK4AlA
wmG3Itfv8mLfzIS84Yb81n7PKPNxQDoP1ggUWZZq/RFltputavBs00hWjbndsze3dkLrfmYwm9V1
vhriMOv1o2HmRhU9ozJhDQHd1BANoo3ARmOWHyB/5nT/bGu8zH8P2u7frL/3ARDzJsklEXcvY6+r
EoiplKVpMsaQuhfYobuEf7CeKjNjHhPtQVNnKzJWMqWjkchD23BlAI5vylH9Pz4/zSBw5y3xCd8p
WQtvXSklAVqpMDPkcR4A3YgLJWuhq4V7LN/DTFBCV1wjg8dboMT1lekgIsQa88mICyM/2SrjiVv+
VF/zCAFdaCHgpPyAZvpUY6f72bQn1Nnpqwwg0FGmI7/jg56EkaqT4CmSW0HPIKX0bOb/Weaa6l+c
05m8/XujlvRIOsNJRnQB3v8f7oOoFnttgJklpNUBwBZcYT2Ak993MDfi7WBJepkSGqHf1WUCP/3K
M7c5pQdghUwtEst2m4ylSlX6KkHWmKe4wDguzyLjGu6DGttviaBmHk7sxfpCYDTDXTsxDBYIW+V8
mqKEpuzGwvfJytEUk2vxhAOMX61+IL/CZ8rKMobmBzx2calrNcVVzYnvO/LTaCoP7DQ8HxvVqPwO
ihaSJloevZl4791oyGMUYqxHTEWlegqdMMFJ6Nf78Wcf+2vgK4kqBEMt0KSpDNCPBrZbMFipFmo2
mUJYLFpSCQpSZGsYucI1naStO/ZOECU+pFY3jyNgTynt+KrqAJKifVne9rJs0w4a8zkp6uYMYphd
M0IRq1C7e2rPOWsYl/JcKEJG71i00mjFWdhIzfC4GbF8A6nI5MICDoWSEamtJur3N46tqGl90FuC
vHyBO6IHGCSDkpLpifH6BDhWeu591rSH5ApGuZUzrkkXRsmkmBhZ8cskIgwP/cDFqKnWUQ5wkYts
/GLCdPwTuoLSmBmuKhx9bdTUHGhAjt997MY147sDEDrXusw2nHpuAAgagsBDgEA8lkskUZ95npG6
5MYNzzxVTrOEW7wssRxOZ7pDBR2nZLt0B3mdaY8rhwOtq0Hbugzx+4r3Y3U5Luofxe4hHvAWgIU1
55/n1qdDobhFmHYtBSrFMNjCVVGaLRmnDOrZjmQZLfFx5qKs7bJ+HFOAKlVTwg3IhD9rofcusLss
VDkoYfsXPqq6Vx9dSI954Z7GovUr4EONMaLwbH/cmcIayRw5wbX54ZeF7lKy363Znah3RNOZvplR
yp7SF6tmCAUbgWInTOGmVlBrFbcGduDIX6Hgs0r8+RVdUhpzk/kjS/Mtj3d0f+SLO1izZkOeQHpf
NFIoZnLwpoqdW8dzY79ChVPurknlUEcQMgWX2CyptMtOtw4UVFGHoDyk8aT2bKWQOO+07TUgWbZx
8w5V3QYCRm6jk6Zmp7A/SkG7642C6Or5wQT+jss/maT9hktU/hQza/jqNpXEWCt96B0h/FDeFblX
q6CTea4ZHMMx0f+p1W1CV6v1M5BubJsDtG+BDBnpc8HB1ZlAlv3gVvjhvBxeLTvrGsYKICHC//7Q
ZdqiGRSYeFd7YdB7KNLq+3gAKi46q5REHcOlPio+lfJQpXySaq+H4mnE3n0Tow4iE3W6R3y/GSIC
hq3cQFxdBnthsES2G/e2qAqTinaOrALvcTDDcZmk//h5DQps0ohkfdhYuu4yDJ6ff6nqRJ7qu6iW
4G1cWMI5WwvywGu1NnU1FmYHTlIcdFoxiBjdLMzzKyWtEi6mHbvybqRCBfyXeLacjQPff+W3n96B
cItAWk/eHxUeuHCoB/OsrJF2ah1hXMzSkjvjkYjZqF6kUDdypyEyOVdPJnjGarjz5xMJGbCSzfpG
IJphxnu2iOGxptljHB/Aru/8gHEP0xUuS1Vab/pZxawYn8STOJpWLBOtRIgp5gQtansixe1TnL9x
6U3p7dlgLo3WK/PY/ZauOVllPo8syLYsJxq3ImbfU/4wk2CP3s0VL9TqR92afLrGyN5ABtM3bIrH
k3/HdkywrXO2LNePwy25N3nwyxpFbOF4Yjy0y5seLFevyC6v3e7ic+3KICLwTRh3RAK1Qa809XRt
o2sv6aKnTtqSkgkvd6hfhvx1ZVlG4+D8MMyhOOC3Fhb3rD/PvSKbLvETrDAysmHZICNsf5NF2SpH
TOp6frghJerH861+jKyZ8A3gEHo3ZXZ2XXxQ865b8ZGZWJ0ZgNpGVi+zzsGqU2e2WYpMjdJUo/vt
tv1JBzMf/fDzGanh8ouwqJioe790WjJSkJO4zbV9+4E0yZMrDhm80iOMLhcXqqLHVi0QpcyIYV27
6v0vLZ7IKTKMjjW1kO9mvOPecreN0d2QDEEySuk1gGS3LQr2AjvoL1sa8PuM9h8mLI2RmtI7Ml3Q
9PtjFEWt3AwIbC13nl+apMeXSDdhQ4XuuzeFlc4ybWuQ3gEfyJjmTaNN7T9tOPgvUUTQ4zu4t/JS
w5GBZs5RB1RdaKtgRzmlvAo14KDehErJTEgWo7Xh9bi8qKNGt7ida3rWpJm44gYkjOcxW7xS7CFM
d2SoIi3rxmfmL4FtfqGHsYnAc4eLFjz+gbAvQXumJwvkR8BC6eIQv/2/d0b/tLvGDiqSwviPaL20
xkTJiL8vEpAgWVuSBGyWUMz4sjd5L/RsLS4qml9OHr/KiMpgH8W/A4RjTT/hNWsO7HgppRCg3paD
kOR5oyo1vFG5ClgtvFmEee1nmtZbJMy6ZkgjRg4CRvHvo6Fa4G9dpoMq086yaNHWURXhaozAjbDZ
RqCIHSHWgveWkBuHrZNVVPju1KbUhtCeNVT2BLTjNuvGBNObf7RIhsa/uzU+txbkqxueG7dCrJjz
TJHWVYUwy0r+Uh9zBMg0+G4O9buon22daDQuIxlso/sBK/pVJINhn3Kxds6Woo80fwEXlK5ZD4v0
H634FsSdBd6wbwM44YTipZRLHZh+/YqSPH3UctRPsrtbOWPu8oqE7fYQQZOTKYPaXDPay0WxunlW
5yjtdTVtyPNCHXATcMgBo0Mvrk+3z9lndS8euFevYShbGpwXbnrZ560MYgIOYHFqMSsPJcsw0K6m
OxJgUmKV+9U6gHtcu2J8P+GMnGmohPdgk5ISV2PwGvE0rmewpmFY/qZyeH9jjeZ3wbEMtOU+76yJ
ujK20f6VMrn5VM6rVJe8Yi9LI/DGVjXdDcj/50yIYVCX3elL0n8ZOd5IdzS/kOwJeIz/NEZLoiK8
Hx4BPW+j9vYOuvktMbu1WmMJBXxJAXgJ8sbDeDXOeFjNVq0042DQt+IEWZ5DlIKTghS3qbZdjsby
ZWtC0aceOQirHRcq1rWuErLd/a70tKqXLv/b3rWxDep2If7CvUob6jOA/Aglf2/CI8XN1DX1gRaw
ZVgnSUQQ7RYXjwfQ2BJkGT37bPh/ojhtUbtvmGwuJdPPlIbVzECP3kZ1x5Tz6U1dAGnHxmRzeDf1
SDoApfoSxxTMY+mA+5TBJqwCubK6SQcBJRFAWklNgq9rWtiY8pKKkUPxGYs9VoHIUz6EQd5I3nM0
hLn14CSzwwMYKqbZhEeJgQ45TqyZy8wNnKA9F/1TtQk2pvyQQOlzmJWQaSiGYddU7HcCkNQ6qOTL
oKXJTgCtZ/qjofF3OkF/BlY19DtZfjBgT0fmVJYhgdnq2z4T0eKnIo4XO3pOCDrAabvxS0Udpxpp
cdsr8UZfx8kxtZpPkrsCNdwmfLRuLsH8Hb6CEIR9JExQZDZ1f4CoI1HB2Wr158BCDEUXH/iz6gsT
N6I3Uq42Q9F5hOq0lhEjM4Vrb9FjKXPXWn/ft2Mcpc3Fj+ZmDMI5j2W6zC8oFaxFdWdyh9bEwhCx
ZbmVtt5EpEiBAkS9nXewYBM/iraAZQwItB2JlJl0HvFx3zKPjh6x7vOV/7q9GdcMvJbzBSfGYX7U
qNUYbdP7ne7mlckR+cB72AQwQ5mATqQ0hsGgr896PfXZBi6dp4mgHIBSIfLXYomwYkJD7we9F0Tg
nsxleuW2sd1881fsM7Hl+K2bzD2iREZSc7VLUuLC0n6r6zS6qR4IjDNY5RJrkJNbxV+SfryqHadU
QJjvuCoUJcgWv+1Gp8Vi1BvSVXNpNmQsUJ4d8wiqJeBXVSO44nolRANHFnYNJsvyx6ni6rtnGt0Q
GSOhgZwTlMIHKb6GHwA2xZNcXlJI9whzHQ546B3wCWVyw2VAqCs2vtyLFR+qfctHOtM4x3cQiTwk
wRu7QCAgzdPFrf73g+6QPtSYaNR8+gB9SvS5eaa91PrRamavKoLXxWvJ8l/dWjyazyFrPTmPpmJQ
gyVyOZVNUUdMT4BBA85MKqpvZWhMmGPBfR5yqBR8dY5YjKYZtjqMj+41aGBZ3kmcCIbon4vai0NW
Til81Bc0CCehClb71X1nfrDQ2VfBPz26WUX9yLChg/mFK/qW9L2xr7w4uE7RuVTPzvG05/vCFVLp
10ptD/dUprtZJWp/KOJ+qK4qVOcTxUxADO6Sya+3OylXNPsWDipEV9sF6fnuMwELoicbB5ET5ewN
Mrd0Zh9aUjLt3W7VeJDihxoxD8xS1lyFamt/YNEVBZ7B99dbtv/4An78jQs0z7IIH8ENySDGbcHG
PuSb09Wg3OgR3p3rl6NYSJX3Z1wwtFPfabnzLfkDLQxrpk4P+iRE2h1ouh/RfRMwC+cnONY1z6Q+
lMMlV1iYtOu7yNNobs1HWiv6Y525LcFahTLuVgPJLzERIv/qas+ZFvL1JjhKZ+ipPGrSCnT1Rz3q
v+jowjF0AEzVrq9ujkortQTA+t45ts6PW0/tCrFYf9QqtYyPFWC4hqW/zO3iSBfbfPFIHb6WtXBo
yfjZYtuHuDGr+Rok2De/kDiklJwWxRd84baf0yy9IjDmARg1rItVKqqSfNHVlkCwCXU6xy38vniE
DnAbNkKCbUJa9wbW0dDBisOfu8h77nie1XYHkX9IvzOS+6qh7aFV2Mh9Uti0hxxdCdQof1UqTtx5
XfbZeuhkFTq82Dq7jbLyfa1Jx8E48NTIWYst2TBSRIwhr1G1hIOnGyIXIwDZDHOQFJn6GAGjrOzi
vTkOMh+jjonJk0am6KGbxfRGCLekoIy6l1EFMaWNpGaO1jJLJzgtphRkLzMMfTnA7bumufHCYQSs
QyoSxtT+ks9y560SX/SVHvzvykpGOAnGPwJXB9KUGo4mWaE3ybuETYGxoWhQ1BKhbIbXeyOlGkW9
4iJPg66CO5VBebHw/i2BhxofpTdNiDql3JAdzF7eIuDIGzn8+2kaEbHmLXn9feylC6Ay5n7wXa+2
3AZaOXxDJXsqUVfJFpT1xEsl1Zl/Sh222/zbPZ6yLJX6yWAAGlRDwbJuSL3sldlZLE/DTy+NB2yD
GrQnsTd24YULRJZk7b5jPs2On+CYB6bEqJp1apXs2wj6joQrdeyjQ5tiXPKwjOKAeCeX5gbEuJSb
BkPckad5XvaJ3+B7+simEyKSSK6DJT6vnhC1O8n8KkZUWHLmqs2vNlTOQi7he3qiIsO40N+12Jzq
vDER6LIi2yHUSX5hAdkEPxtRWnhWHVMhyTp3VI8ozHl2sbg/m5sVQUTNaBiBrdAM/6Smn/Ffn52G
xhTC7zf/ZdAJQv49JzwF9+9Y2rClxzHUHaZpsoGomK9Zw97W/4Zo7CzoHmAxSyh5L9L0t0InnDa8
T6l/BzBk9ObbzdI2PyhnAqgDqdbmblWAtj3mMbwBuxKdwWIs9lLhJuBIVzymxGzklicd6+ZWcQJY
SeReV9kz+FtuZk6JguC9tT0633YJFX0mZr+cfIm71mBw6xZAHGuGabiy6kh3IQ5vSn8bCPEr4cy/
+sFdXGVPo2/OxdnUV3ri048UskdmPwylknTtgn9TPqRUd4bHgLdro13HQWqO9rbXuBDURaRc3yR/
ZcYDcnrKYNfDzMccqn8wS/nvbxP3pNUtSghG/Bgq0iNwAZssm4mKPxeSR/fsE+xoDab48LeNyGrY
kPLI0Xd8iMm0vKjo+tiuJatVQjr72Jh3j5k0xx6tZQCVfBQmZFy/fhLJyIQetGlBi5vJrEDSdwQG
m0AKp0aaBIY7aR3lbMx/wWxvcmquqEoOOu1ldY6tOmkdOZR1lpFQrK9SR3AUczZUvBZ0BOE28V3P
wt4WV8izZDBGd10bZlu6Ea7SNJ9Z++VUSAQ0HLVY4nAGeRusDLJ/7yTAW903jkZh85VqAhygSPyN
GDD48LXVrZ3w5eNqhWD7a+BZ9LB0Aks+9e3XZvvzqOnhRBWzcayDtQZihe0qI8mGbEzT5sF4i2qv
tt28Mxb9M51ntzoeoi9vqSH0E8s1o7Zt81+xMqeXOeNiJaQWJUnexi2BPTweyC7bdBOhdERM1EQp
6s4YO8DHMd+IkkZvheX0UiNPObtB6giZKAWZmZHPCkGi/fVuRK4oervclkzzQmOk603pihVNa7op
9ce76ttjSuCGcvRmxElv5yPAv2aig1m2NKFNprT/C6/6DuR6A9hlDma23cPKlWUFyfyS4C8GGLrP
MWTQR52XyipLQ1L9tPlBNBkNsSMXeh2HkN5l3/XyfGt3YW0V40DP0CyY0fnWlYO6Q92JLSKajLZE
UtncCN+XKoUaHOwJcW/QK3DofssC3Xsdbg/FLjVKfvWlZaLJyLyhIq/pw5uQAPpyMY/P3tvfitAm
5YAOilL9nIEi9utlveU0DzzwcSdz+yWjJnzawzjfD0MipFU019fRurQv/CVTrg0tiBAQ2UdelDWn
zN/awUr3AM1w3sy7hJ6LSo8c9T833tN6jbguqgu59RSMkntv/t0NJlEG5s/U5rzB7ALR1uRJKpJ9
56csExrTAWqqkvB1XxqS8pA5vM1cWd/x0n5xmhUYNhqrAGl6YOTfBVCCP3wx2c/jlUbE0irsr3L5
x8obdY0JP5J/FbUp4obTB6aRRh9C4io8TeUn5Asdb8J3EwYNLHFSodJLEnqiRvVTE3A0lUHELfnn
FoWOB6b0HQ+YeDRBGHa4EQQbF7+wo0UQWPzdoT84d1K7komlXf6Q37x0Z1NAyyJw5Y7N7pL00GuD
ShHmSKsV0vVA0M1+M1cSnLjHaFdpIdaF1/XBrTh62ENBz9gbzDO5YJB/TTYn5L+lViR9edT25XVj
3xJBPs+mbnSD34qoaSew4PprktoX18oYTSjzm4C5ZrSLRUjqA1yf85F/2+ZoVsvdt85pWh74Zv3P
G9qoytX13yV5niOPfCv/QGl4R9aBRpTMTlPUIrVMNSxpM9P6MdKKthOxAfi5WwEqyO7K2kkwh3ak
m98rW3z51h4uxIFG9nzxCVpmTb1LwvtHs2CBhiSLZHCXgQ2Mdyf74v/rvNa61Olv3Ou0izBdb1Oh
grkWKGATxOL08KRvCT9FCxXrlo1ee7uQt30EycPi9xHjn6okqc4j3XgvBRRRUO5bmDzgTqgKLg01
Wz5uBFGPV16mW2tDsGvmgEl441fXqmNTbZBPsC+LOk79VuaM88+BTdYnwxyEpvQxU6RQBqVjx4/y
ynSIQoGd1ZzzvLQxEt15kguarcKX2UA0Oo0weqG8DOTZbl5e4bo8oZ0/18ev/ZZaytkUhox/Ukco
UCpN3kh/avcJoAcnz3smlRWOFATcHZ1SDP4QMCLrjW2lKAvIx5XhuqCUWLgbsZP/riMwxIYPwB+Q
yYHOgUDdc1+JT7fMMw4iVp2/eN7CsrO0iOXziZz/a6Gx0RKqxyBayXlReZ4rgFFTUNfQ/ncnwNb3
MnUcshUdhW25FViEEm7tTnOm4/L1dQMbHtxAaVb4wPZFH8xXbCXzCQ5CfmaSLjq0JcUJpJQTzWCc
ROWyrOSZfEoatgxYugydY3aKQKRMYb0SzXz7ZFQQXAHJ5Tckd48zNN6wCwf7W0+VoDp+34xge41N
vGX1I3FzfKXKxhjccazM0OhBcJ35TSjqJgRlhqMG7Nt7woQs69bOQPhlv3Csqoe0qzdHyUCTJWU9
iiiwKxd4r3sovhpMo/nOYh6FsqNKfoHyYVqPwYP72ZKinkz1bnVPRtofZafTr/Uriz4nvon/CpUa
4D00H3lsnBf/ykbAmFCxV12ZYkr26RQJ0OQc9OotefTDH8IIstD9Wt0f2f285L8LFt5Y9j1ud8+z
s/oAxJ10LzBNGwshmsLKAfjVJSjvKhpHxwtVC8PPQ+QJ2ITOR5PRfGh1B4rlQH4vfeF/4X2vpfn5
nA2ccxR9Rbi4SJLzn0Bl99TMZjbq0jAcr9Hgzi1wY+T8SPGwNCKCIcCZDtrn2cMj6vgVdop+F4Id
QX3VdTUt066YlA2sSlwYfDptjZ+nMqliAizINhLrRXBhlm1L31OkKrIxlQn0dmCvkDrF4xzX3YkF
DjPFB8Cmqg0s0PvAdWkyBeYfkcHBsPn13+75wlbXX+Ebtt/hWfulPw+9Ig30r7dcdUdd9AjuC2GH
HtBtDVeXXLlX1L71DThxhM52p8gyj2spZwfu8eCnmmO7QQqQkUSmyIYgHlXHmpQuuKjedFNQPYZ+
Rw4QQE47J6+AGyp09gNf+w24BFhndciiBt8RzdsiJfA3PgcQCor6D+bQty/IECRKul8upQMRghGW
1oMPSTDDSP59+D4KeteeRF4ehOkjSuzbH/0ThmwMrzZ4212vmhuT9kBkmF4zG330XMNLpdUBaEcB
g5RQGJugomIvU7Lnneow8bkyADfu9fbx6n9JelVRCpBGtbh+Y8p7hXqylrrs8srfJSIuiVviKUxm
GDo/axNtw3G2pCOWE7q22X0/U59DDXmLP1LMc7aVbclJVIHkyLmYpwgCK6/VsA57UwTAxmgUVNsO
DbUAtRRpJylcie/W+d47ur8F0YCz3jFO/VD0aG8DYZnorwd9FgHPTetn+rjXlJyLM2ZaGnQUzLu5
9N0SoJQVNe29RPKOx2lielItF/P3JmyblYBvZMAjCrBlSYEiQosKsqmY17sM4CO3Omr35wciL96i
JYVw4k2k98Z9vn25CR2tFwJ209DG9aokCsNvcun2Ru7Jgx0G1lgO7OT6GG1M7hF07ANpo0Vpk5cA
bO47bRs/wYUyPs5z370By/hLnZzbcFxa29OMsivc0OjcijRqaWRqMUSYrgEdxUET30gXBF2LnBV2
5qMWBwn3nrkss+Opi7mFiYWaWwFXgKDls+Jrp0Vf3g9+CZwoOnF7rIgixqH+583yMmFLX85nXWy7
UNFGUDUybRqQEOxo7LpYFxTTfVFp/6OzWSNZ/CB+RVUQRjY1U35toZBEFdWmAK/WHOSX81U+wZ3v
1sjdawC/kAoxFiyCUm2wRVw3PkIQTN51Xm07/RftQASxtEBjpBzwD5Jm61TrgXWK2NUp/nqs42lY
Vsy+b4BE99/ZjGlpG7tpp9MfwSa/KOQApYmhNMa3+UETm7dzV5nPt7RuqmcG0cJd4k5PsvIyrr6E
ESyKx8NAsMhV4TM+U9UIE3/XgDojTvB6nUvbU12dBlgms9kmetzyK5cIkS/vzc9RxHAocdswbV0U
8khWf2+SEllywSxZVpx1a4z9CplL0Jw3YaXxjOMHYnVCtw935SdlzI94B3qH1vWNOxmbzKSkN4+O
LeFM8KoYqz0wJKQmov5iI5x8Cs7JgFuNqTI19M3AFUZAldaZZ6DMoGlJ9ROKl0k9wb1U8OHkgk5Q
juFmLtvbbQq3/Xl62IWF4SAW/3An2WTXbFJiC9+3/xaph6vpBCl9eL+zBB43fraxwPglxXwxZ8JY
EffTX3NCyhPdm8o+LxiNT2nUhCAJqMnD2wx2+KjhmdirDP3MOAHdjMnDY/hMu2xViLbpvKBLwqDs
/0zSP8f43yFKZrWAwnCtja4Q00r4TSZrfoWHZAROgdp4x+ei3kZe8XC3EK8Hf6zlm2NmZX0p8nPM
FoLLYMgiL6JDxhOn6NGs2IrJUVoWEXuxRlBffxeFY9tz0tk1rkYPI2pgJ1VU4fD1DSWqFgp8wFCX
NUWIvVqTuLUnx29XuWVyyaRhdIwsriTGOLld7xXmCrgoxAY+zY/Z2b7zDU9rZdqjIPI/QlZqYjdt
x0p7gmjHclXBegAsaDgQ9e1DUNbHgARxzWortF0J9sKLMp9RQW1K/wNxyjebTL3xE6vFhDMVf1Au
yQCvgenGOykByiDT9pXZ2doNGhUf662yU8dgl/0w3nouTplCuuiEOngXQmx8ioSSltc3I/9eASQw
Txe4eut+DrdlqwTLTDKNKQcReniEf+iEEHWTw8amg9GN9JDZN+k5zHV7erHuASX1s00tzq4VZYDH
JwXJ0awYaDMa1NB4XsW32tdYP5zoB1pBKOml5ThBN2oaBtPIyF8VRorWluGfzMXORITeRvPm6qnw
FNM2eMGoFIN0qb0OZ2UjTeoThJjyxfwYsjK3od5/5kuCWDq1VYYaT65SI2qmWVSVfWfvCaQGQaT/
EncEmdRV8GELEwybgUmzMIOzCYRt4ozHMuL3hE0bPxI8Oi5zf5yxLx7Jmd5n22a+UM5+6/VhJx3R
3DuSM9nJYhsacwaxTSLi9y6odp7DiyGUqwObyktc2haRJVSSZbOl3ke9nYUntc1pIWFgEoDnDyoR
g5bC+kD6QHxX/QxYZyPWt14cCwT0ShnttBVhJBNT6xoZOiGJPvFwjVkpto9ls1YkzIBUT4bU8pRr
eW4SNVA7i94Efmj4figrzJE31rH4G+zuQaE0UWzmTyMNR/z9BrjU1H5CBhs36fI9z2AXzeSO9PBC
noBqLNyJS+89EEWLlSVLvb1m2BcqCETPDSSbOH3mIBouCwePvH2ggFxXiLMw7e5o51BwmSnyod9B
bOw4etRh4kjh0cNesLcnE86QXUuxM87oX8k5iYF3iz1c+ZXtdoYgnVnu/70Uw3+kz4o8tb4EcDyr
y5NzVr5UNz5lU1BQqEN9EJLy18y1W2v7mhkWPqN4TGKsJc4izm6PQ+Y3PA8QX1L3CuEVUKTU3MQq
96NzCVp0VYrB0DTmoglNYac20L7j+VkFnTdnEE2caJPkx4zvi0Nk8hLSeBbY/gDeMq98x0nmYJua
M/i8yL+Ee59LMUwl6vrUcmBE41oG5H+VcqGjhi/uQ7mC53u4isEhfNVkZdaYIfjk5Ask0qFuDMvy
O+Nc2k7tSj4AhwUh9mxEhHRBSo6C7BVUlOB+dmYDb4ekAy8ENfxhRqkpk0ancgivfZrzeG9bZkn1
LufxEpRNOhdrZDECSSe6YPdAfSOuGGfTjRr1Qyl8wfIxgAQbhpzXG2/PaATWz4MtG7zM+9ip+OVb
pvWeQcJFiGKtPEakHEXwGjVDoFhWyaxtdKQesqACry9JJFD5lmFPvN5llbAGvi44QMuhzj2M4/pN
EYpuxG+PWdwil24Phy95IsIfaRqiP5PSrxToZrwZs7Ny64ghXL2JkQHA7vXko9fqD9bAGdxL2Usy
FqH5lt4a42lcls5RxN8aK0CUb28u1x/ZBdZ5mP5UxGc88mulbosYxqx81teTSA6SL2am9upDOf2J
ash5nU/75lOLJSaX9E0rAu4oTkUjUV84b47/kI+mPHpoYLvr2SgqzEpejA3G37djeGtM55z5AX/R
QOqENbc7zcVuw70pzoUx7SqVBHZS7LZwaIWP5hdzYH1JeFInH7U/CNzIZo4xlOCSrDfrxDP6ScJf
ZMBoAotv+DVmEm3NO0KY4P9XxHWzCamhMQCI2UGdlXpKyI4mujYf3JqsxNaUT5LtB2zuOLCpmpLZ
qTMpA9JT9jmPmiE2NsD7QUdgBtRc4WJ3ZNA7aE24D+NQUaD4V4WLb1mJUF0dHckuyPBZmPoo4ykA
wCbXe0OxAJruVOKuzrg0tYP0uuPrzHGtetuvI4882mo2aBlNPfGYOrEzavYJyj3zf0dZ6kqhe848
UQPwbkZC0eNJvdenuJ85QYhS5J1864tD0aP9k8DjhQVf5dqaLOdbwbMlKHxV2P3qMlX8ZiHglAxV
Bli5y6/OLRj7AAaRxdKz7IphDp2kbNikmXPE7J2Y56j2pZeen93ZTPi26JcfWmPNk+kS15GNy9Yq
ZZ6q0YIIfc9v71VC4Q9YrK1XE2kKUKm2gaQROvG7w+D93Myh+MEAc46AJMlhQW8oePzVCAYMsNww
A2WUZVedr5HIcqMkm5utDskETt5k29d83KS4eG2D/Zr4jAYSpbiDlcSJTCpYM2+v+6UmCSjA+Dnx
EApcmqyxDG400+UUjFbQVZH3ET6Fq4YTYgdRZTJIdK1XMYHkxLNN4wo4SH0kO2RedIg7+Wg2nF70
KnO19/PdFrW6Q0qyIKMqqAGk2RW0lBumoahA8pEnBnRnZsaEYREHNjn9Xs73YfpFA2o6jO3/4hJ/
q8OHyIamuVSvUsa+zwlxll47PU91Sp4YfOSX2xl0nX8S8IiehUhqdkYjgffjjSlwL/4OXYVh4qLP
w2EJKiyW0gmV59m6ps2oFU/XFq9l32ZhecIZE/740CMLfsQcXZoU/rE7UYM6XktFEKWG3/iNQ8JS
FxR0/+7mgtW+IXr9IT+GVpMVUEkQO3XUNn7/YOTScJJRcb65T/x569UKPkQmWftU+inT4hbWFKDT
4ERNfqRlhiUH90C0hyU+pueAwEAqtc6/l/nYh1fDncQ4FrcYv7OChyz3iIVhANsdBnRnqg8zhRak
yrHYBGq6dLPp9thxvatP6vqplKbQqJQgJJVyFesRoh9w67bUUouVd9IalvVe5F7SOmmfzCvOZL+X
wmK9x4OWaCrszxDPV69LSITN2NQZVgPlQdi1wJKcJFna5SHNAeipco2L7oQOQoBcmLqsUgcQORrp
IN7lblmCMn9aETy1HjRddpBfqS+iqACM9nCEPz2JLCzPPltqL8+nHLYYUqGEDY/XaN3h6MaWRSmO
RNkDbWzFQpfr8k0n+0lT4Z7cJ9omB4cZyVW8ocJGpNCI75xXTwhNmP/VbAJs89eoONz/ORh4HfcB
CChwkw8dwK95OyZN4vfozvw8LpqHjeI4HNRTanJCQ+4Qzf5DiuWKrasKrtlfz2cEjc1Teq8uVZw4
60cg7l1FpOnyErFOk9+kSkjLui577gXA6QhI6E6LVXwn4yzCjL7r642mwhum/qsCWg8oX8JYxpVO
DxAFFgCAiEPY4TGqRILeeHe6l+NpxAOZtSx+xzZYkQy17Sp+r42PqCw2IWtlqcysGfxRhmkhw+P+
VqHoq825ofDEIEjGJIwN4fbdTvhCgx8/GLwX3X/JYFamz45tHqEFGWw4fEV6UHuKc+QnU/CDl1W+
/XXN6TZtPghWDMt7fr7PP0ErxHzcZz/qwKsaMeQVBuOlxVxVxe7sDWro44jNh+ysr+3j9uju0Rjy
5APvpVC8qg/OXw6Uj2fIGjbe6FNeZmzydtWFWZSteR+QXrWLmUmafPzE2ncyamb8GHpctA2J3rte
LSd3t2aKZyMM6/inxNo3hEBp5dlH2VFYSWGFO+jKPmRYV5xv5Eg73lmuTIQOsFTPLEPvZ0WEp2be
MNXj0fT199fF2aRnB4L8ZC1mVrlMlxGZVTK6K7ncSh1yzNMFhnPZPAe4XckZAH/qEbkto7zHeEyw
hm/30rQ006uLnrZM1lK8isbDclhl8mDvrkTR8N0Emd0QyJ2DP/jX7XiKigLaZzrk+SQkNe89TMjV
qrIgZbbJbzW/IMIr+lQrIv2trRd3eilFTGJOe60SyqXhoxdo3id6AcErdcrWsrGCbY8A0bs1+U79
qVa8nuZXNFdwpzurKUQut28h4+K49Si7CDvz6zjl9O3WpN73RB/PCHn/rJcqKzUdzzTl4obGNX4v
NeYeErIDZnxYWdDBadaJTtVzeOLzFRMme2pOvaFCmkWgDkVKRGXwL1eVYMWmpvEAdROarSRaBQKY
jpNxNSvNrnuPgGgvZm3JT1xwnfHl9gxbN24zhRHQ4zIVmuscHXsB9OM2RZuUZNQiqrX39IN9x9Kj
AElO4ZOIxeQY5zQtPxTcI19ChAL+wQXDWx+PTWo8+eRllOo52neuuw9Z3bORQfHOG6PYN4cO1JRR
zOeKKax0nLnrzmaq2fEapbzLhVmp7JA0ayE+uhzeeUXVkZxcWurmnclRat1cssZzOSigOVuhUS5i
vM/OWUpup9FSr5JQqGJXfKbXZM5xPaGy7ee9bG+hEAURDSLa3JM83EvOimWxzV0gE5meWcFMowmZ
mYtfNx/yXxXQ2T8q29KC55+1x2eze+8Ho+xTPI4Xwbe7phSFpRl4lPcr1JhTyLSjY1eE0+mAF/ay
dfy/FW9T2PBXNELsu6Ddt3zdhc4+sFyVia1oczuBTFzd6Nom3jAprEdDdJG7N7+tmUXYXuPa4Qmp
7SZqw1A+HDUnPM6MN7bp96Si1bidSa2EHhs0gTtv21OLERxlX96ZR7ddMnJ3jaXqlQxZ6KhK/Geq
fCQh/qT8I9P3tbcp4lRGEkp4Awm/VgoFlVcSGI3cJf4VkRy0pRw+OAKm83Oz6wH4iwI48lxbTSn1
5BajUtCtHR+ooobYla0xtDI8PuDHYVxfkJSD4qo3mpPUlRuaKSwfKzn8OXXvdrLP9o6Wi1JjVRbf
O9aCTIPDVIypi3iRuhOoO6okPCDKDs1TCUb6OAixwhMKAoBLEtEAw3NzfOm8MPuL+SSkuHozKcXk
ArdshnCG6nOtxa3JznRS1Ce7iQyT5nC/sWCn0R+Iajdum5eI600sYKP0lgODmT8AgBvJhZUnqTIv
byJjXBE7f2aowNvdQY9cpyMoFhuq69AhuZ3c5F4lA7C7qdqnkRmmeFMVqpW1W/wWIcoZf/IOh7KM
sxAEaVkiQ4Rrp6+HQlrQ7KQG81KiIAm3EV/VYndUPyeZd+amHpF7uVxdibwAzTazP32VLfeOo1+y
EZGNkXm88d2p4BfxUdULav5VcrOI7kDuuW0q/rJm0Thvy9Z4BjltVCuCF26l/RyHKLz9JpMFs5cM
B+DIcxzSivyzO7N15iWhBeMRP/AP8/rC7mUmVA36ywXcqb+kZuUYDvuQzej8JS9uuWu6l4AFQ9Em
w6M0JONJbsM0kZikqg+28G2Dde9YdoXvLUnN9MQzYQZeYoU7Y8Ue70OZhyRUsxon2uequ2nTFsj4
tOV8r6s7Xv8xcEYIL6nxDVZKSAEZ7krAe1lQ/uPvCX7eyuto22kKqv1Kun8q7JOvUOccrPAgyW4s
zSyUvo2XDI5nRbAEkJw6Lg1xir0tyrjMq3E+XpL+x4IQCw65NRZBI7XCr2ijBTGPX6E0orU9+Egi
0Mb0oJM3+BlKzHtZ/L36g10W99YaHCcijXCwLLSb2ehlqwsWGexE8fhRimOCq7YIxy7uMQXnKFdb
8/3kcEnG7cVs4kaFDNRnbiaFwgkSTBqI8eaXXh6KfwZ1Fn4/HzoS9OoBjs0J1k/TUxiS53iAcUkv
qH1w8KY8hK+t7WBJI19Rzgmxx5p2q1e7aR4YfmMZYxSP2skPJizyPP3+8emk1xpU5YSQWSwqbmra
gYP4fL0grhv6k76O3lOkXZ2XMJCGXVDi5hNW6JL8FUqwHZlg6/uPd5aZvd2eJwis0sFGiFOYnPZX
oWNAc+sd7tKe0NWv3Tr9n0DEgarwhKiiUGbuyYdavpfULByzb7UvAco4p1W3hmhpoxY8g1+8Oml0
+L8HiQpKrf8xVFkFlF8cYs+eS6z52KvigS0TLjAJgzmeyZfao3sW66F/IvCVVa240dE1Ea64T4Ci
yOnrlsCa7QcMtMSHXcHOdKjJw2EyCwtvpXTsGbYvmAUmCeYqgYqpWorIwkzNiw3/ln5c/FxwybbW
KNBeP+p6TmCRSxaK+OS1Ze48KqBLwLeLKiwF/bHFj1zWbyRNpTAnWDwZuyaxwv8lo1dH5zVmE7ao
fvhZ4RvtqZ5tOCZ7enwutpqCUYXjFMQH/N5Nmtmsg3rE+orADcTlFwBfGjWBboyncbJ9ssP8rNHm
xKH68fdkEG28Z3rpK/A54Ptzq6i1QyYTKdiktf09hJWsPwR2zp3X6BSzvCEChBCOrLmWOEyO5iRI
7KRyov4PU9PBS2PQgHhd0b5jezMAwD26Y34VxOf3yE/IN+xzTpR5k5tUJ1ZnDk0RIcXLOcWs20PA
H600+mJ8TcVmhNfrcK78K8egEZZkSSs8Ft+WwbdPDGWtEHVTeo45z8fD73m0L1vLHQTvI6kMEaeX
0f1D5CMDbQWwLVHS20cwIGn2RTALUkggFSxAROBZkRm0+jNQ+cGZhYJWa/rfuazl9v0UL73DK0ii
RLGeCSfNTfjgjqm7XSnjaKiJj/LrN73j7/Pbfzhs+sbnQRDq0zU8ebGWQWqaCIyGuskAtwT/19rW
ujOz2zoS8dI+MfmzGoObc9V1Wj7cNL4Ij3XY8RgH2sxQ4yKu/ya1dVH0jm6b+yA8OaOHwRkxgF1z
jwiR0FW1tJ9mdZDSmAYREmOKJVUnlxHLwLkLmSwyP36/OKs/2USsE/IvZklF6X/NKvMo4JspBent
dPmVV3ryG9UQLTrNeAoA+yxSmhPww5JZSXeGtPAVCdGagTSKQ6WqSF5nRy2lG7/34fLKkush/Gqs
0rEJkP0AeK9kydWJHhghzAC9eXkKhcPCgAcCLjc68KCY5T7aezzq9AT9rPfel1O9+xhxU9Hiy7VH
WJSsilJuTVQlm69cBQRq0WliJirVI4EA6o8f31+s6U3O63BZDqAmRp4N31U1nOryZiljAt4aEQXk
Y9vrkl8utx6wQ/xKGadzfMWzSJjCCAq3TD6Xk8NR6ZmbmaBSGvF/DIL+ismqUZZla8/Dz7+XR7AB
5hfXg4pkRFp4vIRLnluNWbV541LxvrtErWFfP99R+/qLVkTnZ0xaL1FclwJw92gxfCtNIPpWPFMM
sTT6oakl6VfgZUnKr2KEjGx2SNwrSFpUUjxHYC/PvnTT3/s9tY20fPz2POc6c6+kQ2r0hqPi4TUm
IOKA7EQ7ubyzl8YFLoayTCGKdSWVEBCSytLnSYP+DHAni3jN/Dk/7HFe0BmsRBkgs/3RB1arwrLJ
8WN4pFHNrXvlCUIYYX//qFxw1gDReKdmgALjllIaOutkBLv6VQunHt7Y9RIWqyju4UljUpg2YEAK
UzuS6q7kv+sfsH+LVShyePWWie0fG7M8FKo5WgBYh4BWh2v0L4lZx7AJPt2BlVzKUj2vjII4u7/5
PeT4yPV7/e6tZPKSCwcrPXYD5JAag3wlJjXE9LOxya+Dg+fp0w8ZwfF0l02uoculmAf0Vd1nYMkb
DjO9M6WVLf1OCW+MLKUKx57QPiwJgFysbRgbk+VW3FlZXzGkUEMFCTkb2Y4ypkF2OsElPtPzVGcd
2hpb5eN5xJ0IDu6GLiQj69kRz2eD9+MLl8P6JMQyK+TPI/gLcsAzbVe8DEo+zGliPIW1tXg/ii/Z
q2OJ62im56Q2X7xfZ027gImsvXG6xfYMnFxizXcCpXyaF+cL0/ifW/9s45KnEqnPLaND93SbISRF
57afEZBykrahwqFI10kvpfq4YaPWc6cmHLxHcnDkZBbYx3863Kv79aFffvzqEA/YY77tikeO6+nM
a4ghly5yXIg1SCWd2jtfMKz0L7vARl/ifqfIg8YNb8jK4K40zt+c3BgYvYEup7/ftJM5uQaeq1gM
7IjuzAGkXbl3CBpjb0+gP5xQZFOgjvzmQJYqzCCuBRkk5xkEIfFotPSdRALVX6V8kydDrQf0yL5v
84+9FEBj79jX0uE5eA9RW19cSERYOtZKp5Zma6Ggdka9NKiC9yNylXtoIudRcs48VdJmE6cSjuWF
c2sriT8OFILHcUfKCkCTrgk2RKbOm7T1if2gQiNsQTpGSUjBRY394S11sPjjOYuLhNSVQc1xsgyM
5XRE9kOaICQklKZ9iul2CxfPd97ZvbGvA29lEvnlIWnuK5Ej9Ed5eJXjRG3YlozDBp8TfjAaL+mw
F5RcE66ETXzcaEfcmz+SbSb1xB3DiMJuP4CLHOzXb1zmfljjHg+Z0OnBg+3qBz7WWiII0UaWUwFY
aLhe8a9cZpQPn470jC9HYGsDGpWalLEjziT6yMk53D06v5yU/WAt9hzMPlDW0SEXY9EEQeDvj+RN
MgNep726I1w1rqpVv/gjv+3e8p6iynN2ous02sGd5toQxzQlyYR3Ny93ZvA3bj7odRlGgeExOuQs
6y+hx1sY/tj9a+bVA3jGv/DhdA0l7aKU5iKB1uzWUALnwRd+XnPePVbIFvRDfdBp/ifWDAeb19b5
mkmh5TWVaSIJTWpAI6JEkqXClXzHxMvuOE2cXDA2Ofh6UisIDT4bNv1NDXItNb2SvRPzZBy5TiuX
NM2O5wVAZAXCRypbHjyuDYiaFdlfKWlLjh9ZQNH3gtotQUbNqS7PuQAdQt5MrgyUhrVl6Y1iejKr
1brC1yQgDNHQ09v1EjlaqImcZ9BRUXpYtD0gAoLgC+5uX51EOwalBAoGqf2ZihD7QPvi/JkomiUR
P4HmFOVzCNeN3dcD/opCCJuBM1fHKToOp55pf74YHWPAwcHmRBj2vlxXdCkYBeRfqpCdpUSVyoYA
OVWITTvDDMS+KuX/U5RYZCsTnOZeXxW96RLNj/5UXeIn0nor43AdYbXcH0D4uBTyfI3Yiyu2Za5e
iB9Yc24ZC7hObs0pEbx9QWJA73N6R5FKu15BcTW2H4zD3YBfu7NbpAc3WBDnDsZzwBtfq6P9+LMQ
r5E3fbwAozAbnigQi6yCebzda54qtX5XHs7R3kY55Km2ntUgx//R4DL8UNno8HD6NVU02Xs5LtrU
jUpCnUtVxKkSkeVN/mKSQsOc4kX2iTXM7UHw+4Tk2l7CZXCYfcc/7vnoobJ08SPSWONUHh4I3Wjy
D/qJpoX1CrcHJ1QsDzgrURN1P705D4TSRG6Pt93O62jtikrI4iynFIy/gJrCt11pxGbP7An6eI84
5klIsLxtbLcn3r4hrXpoDih2PIdtZ3/GXyI8virlSSuaZOLsudMDtHbUGZSkg0qKS4u9DtE2dpV3
SC3eM9zTvOQUEt+V+IC+pbrRjsnH266VHpv+qhJvrN4FwdEBqKEHmDT90TFTzIR9ww2DBcLI2daZ
nBjtyefhEzE78R8M5ZyTTFqEStY/uLYPgQduBBuLtsd/AEhGt73ye/YqtH/6zLi5GyyM4O/9uHQ5
K5OQYq1Sw0vyoIU4axgxZBVkk4s5DMgmOJf24NDbf80uLcKkhfaEggJWwrI2NvAUxqYZ3mbMqman
KM0+h/YsX+fDsMHBFKbPllOI4LhpGzEnTxDy+48/ao3rOqZrStHzGmi0ReO9BIzHVuDK4WT1+KvY
mor0TpJbWYWuxh3m4cJVMhu8s2w0hesQ+rrCZhCh/Y2SuUtFP7R/K3+CMhXOrBYB7hVYkeP8lMSz
rjIk37bHcWNzy+MkerJ/LsnUuSZ0mNdwcBQR6fXxbT4frK8Ve4FuIT7pNxxbI4Orqd3f/YoOgj8J
01/KEhthgZdVbw69n0FThAhFSZDkYvi+HAoXHh8oRTH8eWGI+ktuskhcLAVSOpE7ZHOBHLsvyphA
D9cGS9hNjV7MIVGYiD+ZWzFjyCWjA1irVNCJN3ufALjAsiFbziiXCUpba8ni6UptydYYRPshqTvE
8QoTa+Qeb1+45fwaxFT3TOArodIr14BaJVbeCMNwnSLRdDz+66m75T9ZsRVwD8CsNR5ljHUKoOJJ
7KYGjzpB90hZHKPatRjyyDnidIbyWOynOI5OSOJqI+/SMJtSdKp2CtfMfdZ79KJXSTHH7EUyGUuq
3NNOfczB3VZM8dNI6vAcugfobOc+KHKegpJR13zxekujq8vOQcer+KhFouJuEIg9BLauDm+f+x05
9KWElPyWopya22ZBr52hkZl8s8qTYEmLx9QMojG7WvLohqj+Sa4e9rk07vyxnoRMMxtbWgVTqVLn
s0cis+SoxcbsIMsViFklggMzbHi4bJ4Ny77BGAg9lWcDBUJN9GDI2ACxhJE5A/dutoNYua2myBgW
EYJo5lj6YCZOn3nuU9lAFhlAjrZIa5qP4UaUgTHnL27Ro+EegLTn3ix6t6MxE5QYAbCggY+iO3co
8BU+GxXSpbuat//dbhdCjN7FiyxetUByxbpn3gXdU5Lu6i99z5+V+87Ye1YKgJoWbDhiqxrg+aHA
R0e6H/DEkZt6HB3AdKwEf7RSLFqbof3rgO/iuFAFP1a/38GW4VDssL0SEkANEqfyAN8LwbG+diBd
UWW/l6/yUtfVvXWfvqtlnLr08G9EIMA7HIx+/Xr0SEN7wGTRNFb9eke6njXSe3T9izxJMh18/fMR
b63Eck9lFqD9OnFzn6IJ7XpB65ueQBQ3p9t1Oup/3tpHvbJqP96tdkT5RBfGi1Vl8N3tXmRZ1av4
I08WG3OIQTSatX7dHwZ9C6rOXmK1u1Sf3LmTIjTWE2Z0Bg+MABOSnZTJCL2zBiKOijgBhZm8x1lf
VkG459nZOJhujxePnWrwuvUkEIq0QhvrbX82qdMbavgU7Q8TMiXlzEQIKh4HNbtVRQ4JNHWBr1In
6W0JTCeBbtrehjRI6eNv1+M5QUxF2Z5CF3dKrPKdFwp/NWh90sWhgiMig57f1R6bK5Pd5ogspp2i
EXjBIxFRH3ZvbHAp44UPZ/JTiwYlPwkd8vKJe00cNZnSKLMWFKWdvsvFBJtxtWS3iHRkcxCK6mDH
LCrbr5eL7nuzxGJycAvUJpSNYoQ2z21ZyqNLp5Ex2BIB4uJBDvPVNvBGhSjTb9h/YW2mNnArN3O2
NFt+2MkXimQxCxEQVVUOvh/9JlQI4QRKesk7iDPrBzOsSq4N0UqVGdUyZyi21Wyr8ELP5KwJcXJ1
CVvLoWMgVFwgMmwzOxgKuiCDyh7EcTfRdiwl6nAmwcwmW++BKyH7priD6YtxFnP0PHNj6Vw7FuIW
iMGVQ4RcYfatfsNyLACw7CaR2e8uDUMesytTz16RkM2GjltMAS/wKGW62XYBbfJSJI20GzewVKqC
ZC5TmCjxBGozNwAXcK1775XNMH0sD4YZZk+95o9orId7otR5kij33Pfx0YOI8K6eLBIMTkowIS80
vRNB0J8KbP7lO8sZeCNLCCjrpltCjeOT6ngMXwxlyFHVNp8V43kjz6ObCXGi+FnrOsa0CuEDr0yb
JaNM35sdqz4sOjUSFMc6ihYjXc4uS+I3nrOMGQiABJgcnN8BFYZ2KiXwmAsEo/TtRRMHT+J7EudB
6OB5FKVQCOLct6YoCd3MybRAPuzXWnHMoXI1sDdQQIM5vMk8RZ6lvM40S4MdpKyPH554bGtLkhOR
TQ3S2qCH/rJgze6NfUuJh9JxnNRxDHiJWrNxjWOhqFadEEAaDATm8Jtj08B/GBLnEDdUZn2dlJXH
Cz2zSxZuBLcztpdoGbS18TWL63+JniD/Y9n44addltg1WywYx3yqyPVbJ89Yz9Kz97fknaMSW/P9
jSWXMqVbIPiE28Ac2j+LBqtg/sOj/tKiG6yGhrWclXamnJTOW+xXDTFRHsISaLmRawN0Qo0Z6HtN
CmrYo0nQfUP50WK6Q1dJP/7Kf6jJh+aTkTJLo/6xwlobk5uIXLmwk9uAbWGwI9dMcNwDCb3dSlag
f3J5k/o2PhylsHxvR6OKjLj6Echi7uDMqqi6Ybv1bPA9dE5Vv4o2S7W97cBPl7dHmj7czyQ+lw1d
ZLqb5KNXYfLdjR4w7nkupU/+NtDpIs+oCrMjz5g4ubRlk1+U3O8Rw3ygkCRrvy2Qr8SL68T9JvWd
qu2m5ZV144/I+ZsO0xA58NJGSO311qXKllrGcEEMzaayEv7UgxriAhgwF5A9pc43JQcoT+F5Yiz8
9EP4IMFYaKAYFItFOEwtacw3DFsi6w0/gOnEx/9swVUwyZ4/dsfXNe1vKFFLeL5famlbhOhBKZXv
wmSkp/cjp55hdLoItNOzXIZ7e7gZfmPRCXIjki7e+eZk9p2wLFGeHI7rbBmCO7QhYRYc3ntXyMat
k7MUy97Jjfl4MqSayhj6RwlKeeVe4mXASZ06pWuh2p19k1K4VIduChTcCXRrO13PGwyDYXUfIifi
4a9mONjb3hCkg8mkD+t47IICsN3bK/2EiRNExOUAkew/dco5FbcJTQX5+PaQiqEiv8q9sXjL+tzX
WW1oGRStMRRqIxr/9+wXiIBxsKFy/8x02edkxdmgbLLGwH9sY3g14hxG5XvRijKdPs0cgsg3v/du
VzzkNgHiNutUzY0A36lyzSGRC/FhmbvsBILcwEHNwlEmDUwLVKwLWIzjYz41SINNiGDSBW19VYPQ
VyGSodvvIXfLOBtTdWbRydckkZ6A6BhjT8AL27pNz33g+jVq5uX2i3WjL5PK92urTlB+EG/B1fFi
bgoyNjtvUH+NJzN1UNCcnfQkF/Yc009tOq/3nXAGM7oe4qOW6VP2fxFJ/MGEhRpjHFUAFQCoiclT
Bsx8ZXoG/nuxjQ199g1o/VHht7A0bxOtwhJnT/eYWRF7Y3Ydirnv+AVTARcxUlh9R8zSJ48Rs/jj
RzJoxiPGdeVC4FSsm1y0MTd8xei3DnEkqsJjogr86fxAw/dkkqOAXzK0zmrQK5zum2jZAasO7DIO
dlLjzY0tmfyvtHiri6+Q8+8fHIqSo2QWgxOutRMyDFUw6JR64AwbLMdag4asB884+wduHNYVGVvY
KOQvDCnLOIoAQ6KD3mSNM68N+lUE0UI4HwJmit3J0XXLLZWMwp1fCHl29E0k3pJSbl7AwN50Aa9B
ma/nJCkqSu5xbS8e0TdRL7Axgtyjz9JlMeqtyGaxPVVDYWVuTRapLSojC4XcMOQp5Hq02/6pb2pT
KunQCSSdL7vUWvn8l5Clv6MH4NYHXCA4M3cp/BCRELW59kIM5486JNY9DNkQqbG5lkAFx4yS0tvf
XxUB9ovKQ6i5l6zdMrXFPEhQ/7T7WFBVqE3+PzONNRYJvVR/TFBaLmx6oSXWOnoxbrqFUPn6n5j1
+Mz/2l3DOSswbiNUAIWdNgF4c0MhUVOuK6FxqQLixLaCkNP5Jib71WAHmspOwuI0kJyaJHeBEoTh
8ZGEiaz30M8183d3SLTo8x15kOYzGLnkOEqfTHxxtKeipoiuHN0wF52wtAFYu6LNBE3sIXxsR5/O
eo3s53livxnaJbcfsyKkgMQHQvVtUhk2T+zhdYyQXRbVGBrB+5ECzbEi+ckpLAvHLMM9iVqd/KGe
4JhjO/5QgmNdrIBgaBPgAwA9PufTxtATazg0f2w41SKDP1YFa7mCFpYs8Ki1SFr4riu9Kod0yrfw
wPaYngEOTze0G88GcnOShvH5sseNKoz6w9oDeG6gfrWLMYzBuu7hbu25byX85V3ZiqqvVhY4c6eC
DIYvot+6u0niwoExTKTATyNgyNPTz4bCJIJVRAn3+kWZCXXgX3GoIlQZsaYYGMYoNQ3PZefEcAYu
Fuao1EEhEUA0Gj/w7M/A4qnk1C+YjEa8vedyf4yWF9V4V3Dpk5HwswOJe+R/+if+zzLVR4wFu4Me
ExIJsA1y7ORGQu4Kk17K1LCp6ERefLpg1gELbi6MBjn4tNRCMZjixfM/ynzdxFmKIoufTiswp4SR
vLgSpEY9Yp1c49akiW1coUGAtHllVUcHjHcWpJD4hlp6kNYK9+ndvePdtt49U9L9RzzKjFMBjOWZ
5rwShIucEcwBODh8jO4hUt21Dratr8fGgFhf4MgGpR4wGYZqH/x5HzbauMS9LfMqg7bp80miQuSa
GnOxDFTnoU8qOu8mgPE0OfYlbg2Ejj3brcHuibm2NcFrrjLwVkDSm6yikSr6znqRSr+puTjuVgE2
epCLr9GbZj04+IGpqNZhsBZBKAiHyIMnx34cn4uyTvRZXkL9/e/HFanSOG2LunA3G3w3ARMWDh40
Y2IWyX3BO3gEHbR56Xmc2jQKSwdWxvNXfAlaqhRuoViPtZJ3oY6qV86C3lzCPSsw2AHgzQybI/bg
aX9tOp2vGDcUneY5zI35zhyIlZLB2aQPuASCVKyu9L/nMMErfqS7iC2rvgIXOaJwCOERlzw/zVSh
K3oEenOpc7htUftlBnAWOwLPH4/1gaGyjGf/+c7cKV2EPIcosnehVNynHH/9XLlGQ5FdHH5xOhun
bfF0zMrIA7GjfqKQvy22cF7OJosXygVowCJL3/T17QFGAQ8glEpvSUHsUbb75GeyHpKOZyKauwQr
BWv8idnTwkJZb+9+jSN90pQ/O7x9GoJpHUOv3thPf1Z1y6WMRbJaOahOZRc7bV774puNli2dJbSk
Ynp5hQJbTZfFo8sGQqVFCYNWalw7Toxa/z4EGmE72PcBWCQNLvOUL6/DwCGWilmzuulTyJ7HxzI4
UCPN8pMG1D7qIXAB7bUwXkjKveuSMflW0vcREhk4kc5ypWr/uLefBK21LGT8ZQXEphtKj6Hl79rY
50PYq4FI3Ez/eMlfIvewXFLfY6xdm0Y5WbRGeTN/0qPq9abe8hU45VQp3QUh3uZDuuYnAsUjSqu+
oXmgia5oUT5zYclxpsU+8an4xd3mAwzotpSdYOb44J0tZ9oWtMMIV8OSyYY/wY+PaJp6+mt02V8G
uc0TbMflElxlsaS03nIKJ4c3PIA/YgSk51h2b5aCEA7wtCHpIZwYWWbnFgLoeeoXbeeJzLu541l/
4JcLbV+5qSlsp01hsesvJy/dD3q7IDdQsELAx3Y4voVUAlAkoaMAnySMwyw3Gk4irMg4AwfaFViB
KU2YUqz1jv2aaKwr9K3yd0lIsOhssmQbOTXwsGmaF28eSotq/SdJ5uGi/NrHQlgCosxd/Jq/gI1P
K9pNT5/tKTa1b5P6QaQH9hf3hi462i27nheCdFggjZp/LUmNRYwu5yT5VdbSyV669lF/vBFdKbny
vqikADXor7HVibMF/8tJcbgDWE01pW6ePQU6GyNKoOKlSwxkeAxTJfuC3h80BlTb6X5WzeOwcnwG
7OX6FJemArlvaCltIEj5yUwMGuVSWYYEMv4w2/VGQM29lvUBKaDq8snaz4d65qXFzMXqEq372lWv
o4DpFLdMWmRkeAmsbJsQwxM8rZWadtKA8yASWW9bky77Md/ag/MM75mi83G+/AhIEOXT8k503gAF
TU+wk+krjmpixbjEg+BSeBpQnf93tRih5OtxghJXNKr2kHVn74GwU4cNfE9u0CTi6lEXD97QFnjt
z7pQExDVAYlUmTdb0Q3Ii5mx0ftnKBEy2MDnKIbwCEDhNb6GBrIzPycv+i7hija/lA87iISjk/V4
kL/YBaHisjLDwTNFLFYWDeZEp5y4ln0ZW+5hNQ2U1KcTcYKdkUlxGiVK8Jhyru85hocxop7QGQ5H
X1uJpmETfUfePVHWxMSWcRC0cRxrxGQLFrEEsirGIAbv2+AFsU6XhA0fpM862yiAgbrZXxnxqjYP
cOloeZSK8rCDiA8hNAmTRBLCqaTftg0pgDaqF6zO3nqGWj//Phn9GeFfTc8lOjM+pMfXuDf7Gv/b
p2Yg0pkXsyr40MCv18fobjkx1fbJqzrcZKbvQEEEgKmSNsyDF3t+J3c11ufYzu5aTVh8jJq4U0G7
zbf6HLufAn0b8+6O/bDS7iB/aGufAo7mGeB7rOau0ZncwZqQz4kPPZD10l7jtOhv+l+EwdpBaf6m
bmc9G0ZUZAJqMsmrAb93Jy9ibUONVmnajo2/+Q0994Il8zsHoiPYs8cjBHo7GYaerKdkF2tZa8SI
nmELcQ9YtE/jqWMCdOBM0IbeFGbljigVNoo9WDK9ACYqN9lHIJJMRx5SwSKl+fUmGyRZ1e7CzvIc
ZKp6g8U7vg49NPZYUevWa0l2F6KfEjQLIZcUg25aZZBWANTmZ0nty3RzgaE320xMMjwNzl/Y4izg
ri0NyVOJRmsgb0pGFmFIkWb4UnmmbZRBvAiLUkkE3Zf/iF913xoHwGJXP2AqZz+YGEx5oSY/ZIED
ptzSdlDTnMfb5N3oOpjYn+5g6TV6JsYLV4eqbCNvfPggQP/DCJPfQL6jqH3HGo0WXJ8o2gRrcban
nIlzxvRjw4i2GJQv6ulP33osXR281NVl287QqOXH3CQEk4IaSfXOEk8ol+Fe4vxwciwdHKMiMTbt
r4O906Ws5a+PCFf99F5uV5nTSu3ZboqNxMqVmYpUXe1OZCZCOk7Jh7jcYQM9oO5N/6salT9VXa/q
lu7siSk4Oii+QWTOSSAqjG2FLGhPYYUiMYrN2g/nt+EsbS6tmmq4y+Xh/Vh4+9ZDjTDWwBLLgj+V
Mybo21TtsA78hYgpQUatgi50IlcfdfQnKL1nvT3EWKaIuKv63fGo58Ik3kOqVs0ZXxR7u909qKye
ek8rXrXc4spp31bZ7KMdh4BTgdorRJgZGIZ0N8K7OoZBw7JrFgv0g1pbQ3+QsWNZTmUgmhiij472
5xUgHW4w1Ysg+44cnzNmFX9/rFQid0S2zOpMM5E8l6PlsteEUihV1PuWypE/Su5gGEINW3IWDsw1
Az29TOpR/t8mBb9L0+XVDZFSTzi2oIHVga8cfj5oDMo+i9M+wsOIpR6wu6xOKSMBB1s8QdG+EBNc
zTIv9Zib/xl0mydsDhgIsWADi25EB5NgE1Wu5QyFcg/azF4faMEegnfhpJLwiOE3t+Ju7u1A5C29
oDy3ucVwIeliBstuE+vsDRgA7+ibk+rw6YmujZVw
`protect end_protected

