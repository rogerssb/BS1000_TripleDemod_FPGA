

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BJpxc8xtM6CZ5534uckhgVnYBZlZvHtFtmTqHp9IntW0n7yfmmrOhIdnXBGq/t13v7Oqq30lrKfs
NHgdu2tIgQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HmUA8u7PF8GvQZrYK5NY0c4PacPkMESC+n/jKG25bwLAKKAZ5KD9gxH/YekmQdCpqxR1vwPvH02e
RL/FzlX7yzSQzybQxU0bnKnlYmprOuxv6i1DyxuOZ85ATpyQnXzkMCgBMXnxAFU0j3d5SdEuzUeI
HsYvPtqAWEqY9XPHZPQ=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
xlH+oEl0ZT1s87bGIICjv8VDuvpHIRqnhydZhCcaSPCDop2dAVtf/47zP8Ir6N9oth3Z3JZ69FAT
BFnUShsYzXQ7O/61eNw5h5VWsXjyOxugZjgmd7NPZFRtq5SdMfW0CXINZ3I3wYkEqBsBKTZW1ajU
cJLPHxaTFHDKsZPOI5c=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
j4y4YtOMJzmNVfQC+SpXQ+HrNa9I9R+v1PKEa/3k3DPr3wDFcvw8YNexH7RC7LhhHX4HY+aNW/2H
Zv291yoRESMc7eeZkyt7DzWYWWqiV3aTj15PN3w2G+5TY+ql1CwE2141XijKMXCi1rr62hzPWsTL
H/Yb+iyGBth9b9zYJv5KQVWG0F0fzO13plv4aIXe2iUWcPsxukh/XJe5kBJd0Sxzk8ZMSC6+gd+K
Sap5osMNamJKVcBc+zOSe5PtNa9Wbhl9Sm1NV8pDrBoqYdg4dM6Gkq8a3tdV9d7V9uhuExNbpIrj
4MvkL8aYhk8Mb5cb9FxXphEGqq9stA5x46i+tA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZzkyHFgJay58tUlWxXVl0YwBkuy4/z+IN+39/cq+t+DRbIsPGbCsivT+mLyFd/J/00810d2lx4A9
qhPM/pUEkFh6IJ2wg1lzqTaKcPF2gNgdx23/8dVTROakthDCU88jHXWOz8oJRg4DfVB0B0icIwyb
McAW8OjA2o4UmfNqAlEhYa9rvuUdBxMnblcfE7OLOi7hKEcLzxGklcunyRu0ai0JM0XePUrG2KRh
b4Id9AzjyBFH0YS5xPC44zRfGf0Ytm7AVGWkr8ETFG0IiWyYQvsCpRdK5rr5mxUpxoTGlxx2B56W
XnQFT7WDTMJ1CsWZwqtmcfwlpfCiIin1Y9ZN6g==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Mo+vR9a/HCXXBZ2bVK4rFGoC1ibJgF+bwhtRGr9PnhDXoSSplIOcR02HUBdqOABn3idUw/P7Lygr
OOb8XgyuHvnF7HljDCdJeidfov4bo/TJwy9LRAIu8xMDN3y0D2QVqXdBC7ysWPh4eM/PhbWoROpb
ksXg1+uxMyRXW8AoLLjhgauxXYQbtk0emtnNldgU0wwqWlo1YYrzPx7Yk5VFVdv8wM6OLXOfVDfX
wjMzrdO03trTWHe/ScHfRbAUtKMAY8FFzftZfDPaBU0WI1tjD7AsNKJPtgL6DTSY9/XefXLUcRc2
Wv38UFxgxJ7TImni5gW9jrE6vtskmZ8LT5EBKw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 920768)
`protect data_block
+Y8OHwp2oORQs/kjDQk05guUrdrafEPsk1Je5OC9KQ06qxAuOLUHtwvbz3B9RiS60V+87Fo4/e3i
BmQyTEZlDKjzKJZc4P+7cOK17G7aRuCH/XL5v4CdQmCJXgb8sUkunK7drK9qtlevDCCeXxpkzcTx
Y9ksNDZj5AY07rSpn1FMAhPFqzbfzkr82+xQCobEbYqtKmkTbn1FkbWMCRar2bmTTGTz61x1YAe3
YyRMNf19Pt73FlJOtlJFU8Rft28D5i1bMNjWEZXgnukR4a1KMTnY5/nJ4yYHee/iMjFFWCsRnQIv
LTwEdcbXDWj+rvrg+D/D0NgIuf7BgfmneIK6FtanM5vkIXk3g4nLeMm22e5/xIVgQyIF3jxFqEIG
5wRIjtP8LCgkIKfpx+aAhErI2dOmp+zL2A/fcpIuz812Czw1H4w/P6qlg3UG61ROWLbN3/vSTvHF
IrBksS7YqSPvFWQSa9k/vYWcxY156bPXwYvJF4boSC35IJc+OIB8P2iF8IGCGnotQ2a5tfW1uNiZ
VLVeN3Z76Ieb+1QmIn03+QHPUYZI3OlQ6bLoa89Fd3h1DQDbwi/zv9OEqSaGJYgx020o7t9kJswV
ilen2KZOeYdACVY7qNhXOMX1JUv/IDyuTgRt/ddpO4QRQnkOlar8Z6zeHJDgEMagNJ2Zoma8JeZS
+2YYRxvQqd3HqHshrvotOzJ5ToE7x4quWRH8pBUfgE6vXbQ2bhWouD9/mUprT/VUBGeCO0F4+Ls6
anku03aHWpBRs+z/mlXWRuGK9K+oho25HJM/Ka9X9JBPKZzh5LWWyWfdEhe99QLmCQTiAnVV+jB9
+5vhqr3PITU8rAyeWRYsPx6Nmd+JnTJWekGkQAaAZriBAS/BHvT6lrnxTD490XQzivPbAuCL2VL9
b0sH7+x8dXa/XhTfsNY0gzU7kxHEO2LQANpuuYA7V8EMNtT+ViUuu08ttapFadvRg/2h2QK/oG+0
+1Y2fQ8w4pnLwxN6MIfeGPwZXZe36A2vli3RLqocxacDBFf3wU+03q3pwGYfQDpzibLTohhIYsbX
vOfqmkrhqga22AsfGrSUxUmeRKG6wRWiZy4j2Kha3PMdIW2XksgnBWeDRPywa3Jfgx6HUcKFQmVf
jTX1sxQFd35gk21ctHE/fsDmpH7DDyxkeFXPKUApxdIxE/mxZ88GYU9exvTa0Lv4N7n+DvMT5X6u
fudKRGJI+MBAyfflkKgaq6sjYFgit3CuO25u1ehSG/qtetgfVPWnPAfE/4Dyz2XBGRT3ci0AaETQ
yVstBczhZ7gOjKq+KsdWvKRbk46DB0amPIfbzgQiNUXv1L1S4vX661TuT+wz8JgACxF75yi1BqER
0VzE/TDmXfnVX5VFxIWB/hBvgBTAtM1zArwFCmUV0EJDC+PH9s4N+KEAuHbQIitRQiGI8glbLWhL
hcPvvUiqPRaYljiqxt2NC1wxJKlXOKOsvR9Cf3xigU1gnf4Vj4doWpaV4eSdbZ6DkdBCb8112itq
6cdv4snVLYLKkGsvYEkx0tzykvX36f4mUuj5RcPE924J6ZfvSpPTBl1UKOKxbCF4649ruNGiWyxH
jfA0wngaSa+ZnHKSR2JjYcTHwjTUC1nlUhZ5AEabY6Vt9ZbjwnZ99MdJS6kM3G6RuRSXbg91dOI6
x3yoEGYnnqroWPQF2moxKe0OUY2RA+IECX1Js2R2Pk0p1Zaowlc0zbHknl7CkXt3MthKmC0YcBsE
uG7Wm0hfcE5zUGFnJt3f/q+lTlloe+GZ4OzGiTSCN4ZPM6VBibNOKWAMU+AzeCZWN3U49twOkmGP
bTojF/2bEkQj8fsJ0sKvWNk7mHoRkRi/DPVO968tiFIMMEhRvDid4JRAaUlJQKKTz1Z6o9p0qP2v
nSBDanwnEoYafKAJ/f18n80lXJ78n9TXYHAD5llRXW6+vxtEhylFV0PpUQzjIDM99LueNtccdB+o
OB0RnIW3itXdMb/+IoCA/nX6qeseoeir8GzgXzXFG/PPA03nrDstSPKH6hoKGkHfGKAFRJOzrE36
bP+VII8pZKXwoLYqIpG9/W91m/NfLjpUL3sjbT1JeIfDdNDgtUKSphhONKO6qMvmUgs6DJXGfp3F
C5w8oz9UA3DkCTIW41QCFc8OUFU2mkXzFqiMKaMrqriqhOBs+sqqihTxgHwXQ4BRVDVCqMxhChhW
/tv1rq177I87yHdJ+t/3l/8cYH1An4O1Iu05AvdW08hoLNshG48AZa40e7L7m5IFdmTNKF7+Dakk
t9TmQkO0FzaLKL+iyoZk4RRr4J8cHR1XW+ZpwhsEe4GU8MmZcustHnw4vMNtIFHq2eMp1d0I1t8Z
A1znabnQdZdjwW5Nz0JGgrfpkDcW6Z4aKlpIGCIocaS5AUFluRV2xwAnhgUc4RxHFPEIgzS96dfi
Erh1EWm7G4aMUZzsb6td9fl5R4Xr11LxIGqyvjCM+q7aorYLP11p0cc+9XfvWCEpw+R+80KMCiiG
b1BZ9og514G5oH5dkMj75nCiSECpm5fG+Dpiw09QL6ihNsXtLkhEnftJV3RlDCSDNIRML9w7BSv9
k2vUgCelrqylII3H24RC4zy9Xw2lyaohOVhDpvKfHbBGeLZxwYRsPGa5nKPlVndCvC5F0mAYvxIl
7sTo/1nBZsdtmumqF+VQAYSvHlriAgdGoZ9obJdfzBKEgk3ZH9M/KlOK2upfFNrAJw9eeCXzlwqP
QOc954uQ175ZA/nW174Uavlc5PpVv4XcJR9qfdN3ooxqOCT5N39kd9ZckWgGbc4fbCofZS04tLZ1
nHeOGfgediSGYAghcZiQxtgn7/gSfXQYq6y+cOif342SeWBaC3bO2wFqZJDGyOte2RcgjvEkvwUO
idhrmoLTC8MvIam76+HROh2OyPrYp8aQvKF6Dq+tHF2nDKL3XJ6Yngkzo/wLq2FelqQVdA9m5azu
yiRp1yN6GUlZZzO7X5c5ve4x49BcbAEsgOVzKadte09OadjikWjE6KK17IVZFzC9k+JgPcBnPS+i
6i2qxAJPChRbcvhjEC6gZxc/xKWh+1NefrpKD6tbQ5jlXzQ/FIuKuZKKuxShZpM4XuxlKnndAEcb
K0nRQeoMUfJJ1wKYNfeC2tWq7Xj+cxgsdKEnJIGaTTSMgIi1yy8/TOTbxBTTuYfHSDpEn3+2V4MZ
Y/kuG6uyk0cvjf+jOoEnKyC9e2w8gR8HTdDEPPXXERO1XKwsXOh0Sdf/j73KdQfVPa86r97Hty10
NGGLq7PQNgvNCAHmfxymTIZIFOG3hb6Kn0ko2zbZo2OEputCLEtKj+Mf5mwkjR2cTXMOkqoDAeZW
KlYVEhP8UB72hgcW1p06L50+GfzxV//IXkJtv6w5grOQlInqKur/eB7qRcnk8okhuFScR6YzU3L8
2G3qJFwZH3DgkAx/R7i2eM5XN5FrAVcihtv0o2GmTz2l52zdbxhG7RTLB052gUSnDzB0vSQxxAj6
8CB0i4hZMPz2P5tyzm2/uXe1JvS4DkmbodO46upz5piXQgQQN+U08JxGVBj8v9uy2k0z5KaswUTv
IiWy8BNTRY/pSuknXU+3NVBaOWLn/6q719EUepKyWSBp2YOZ9i55ZVvx4qQVbiF75FnIUiJeR+HB
u6YLub3lcA6/mLvYnvaJ+a6Bk4BxB4y3Wq+MCUjs3IgW6rSqdhQ7EdDTC5MIU9sKCYBKgrtspAUq
OeU82dBsm/4VJqglydvNw568k578xu97SlRDz0Vxs49yoXmAmjFzm0S4rIdIomJN589crFCaie4Z
o9lI0u6BJD1+34DgTz1VESsrUNPvGeU9oMk/zlUkOrkzgFAb1/vKL579QKyOjUlMCegkUAkDFFej
nIpyrT9pMAI5KNXNS6yJRyANMsC9a+UF26+eqIYerKLGJfw7Rpm8iFmQsDcEb/CQ/SnFIQeJaE59
9qtqUx4JFS6TR4s0EqINPq5c3e6PpIinvyAtfScv6avIgbLqIx/B40QKuBfnSpeCXEiTGO5hCOCW
tSoZIQ1KDXVe1zX8ukrR5B2/DMg06EYOsvUVeQVms3+2rHxDhDeHkyDhvP1poglw4Wn2r6oHqC+q
i+A5M2UMVqXIm53D2K9yAU6gdudp72xFHZwHw7KIxs3E18+SWwjKRA9/aYvNn/pbAdwoHgZ+sjB/
D3C3q7ZVqU8YnDF/RoscSZhAlGIb0cbvqtsbyjRXrlFuDOFFWdULO0zoKIaGLqXsQyIQ6b8y5PVy
MNZG10hKNQrwO0fJYS893DNd+VCj7U2iEA9QqRHulMniASmeOEidDFGj9UtyuHuwy5PXtVoZfFGu
XG41dACH7HURzKDp6xbQ0GGsmSYgtrAE2Ct43nWZcMxmtY/XIefZbGHFix4ddYJ8gANNuQ2Er6qp
+JjAm/Tq7nIOwKRo+aNyu7w0cFFk/jlBQ3P7umRJakxoAH4QyA6/55ov9Be+BkLGfsYgnU3Cxt/t
8rB8mVxfYKUKrLej5nKaVpPtArATndUEugO1ueSqG5gHBgan7ZOjqXeY9XyEEysXIKY8nFlIm8ui
2ZKKy96LW/6I9ZO8BMQOpQ3vLHxHqcTG7oMZvOpxCeZuEuoV8D1eIHThZac7YFOhN2zVNspdh87q
3qCirlsjQGumkKWnrGGJIblgFP39Y6l6N9USGh9D8pe4CkaGQgmM5mmEkLFH/CVuimtJE4sg5EiL
g0YTs2gz1N1qYfevTspMDcknNkxzvwtdnjaaCEkXmgnoaWipyZVz8DquV8polIkpgPyvNstIm3kD
crcA4E2xZcp9YXhppFMZdSd8N0s8NRA/O8GHkyEhsxeVEF5OPBgIxGdZg9aFx2uo14czFBW6ScLV
W9yK64JJg0iam/yfoqEQu111/UvaR7SpiQNRv0JqrbfcqjWMzuBOk5NIoffvWcTtjkT0ABD6N1cG
TBSpLeqpEj81GtXDi1iVa8Z2vrUbTBNhLSfsP/FJYGcrXfGXnMptnB3p8813uxcZkpv6I4lIdJau
htDHTwyfxlDMPBDJPqWLaxVqAbYgs8bXz0vDS2qhuIzttkCvrwRXXomT8+m9ybcYxuFJJ9hWh4Vb
TVBg84tdLU1OJ+7XM9C7G+Jtg1F6n81iw0k4btRH8SNnhFKc+qbdknfQga3VdpNpCKWkB+jMxWdh
1QCDqiNwI1nPZo+9VWiD3ZyZ5vVCpNqVscuqnNyLOaZN44Cqg94b0ALlrgOfPiQBLVOxeW+wyO0q
UJj8c/1wcBe/KbXAHuDSfbO3A0U2/eqF3PfTcWH4w/MOVAuacKEA6edSflau0S+HAqTrzk39aYxY
RtutvsLpFOEoVn0/Xxb36fpBZde3Cxz6K1pL0Z/SMpVdffnRpnOkYDluHr/u5tQWvlw/iffgLdy6
K9h+sD/sPa01rNx2EC8UN9jVdouRYo08dnYpCMdKB51oMQktU1ZyqRLCUiiKW866kFIhSPgDWg7u
/KQGWE2kydIlDUMb/k4sHtb1lf/WP7RIbm3A5c0bF/3vczzC3wbCgwhiWfi/YPmZiL23p7EfcpTF
hoFNxiO62qo+ScYKz1SDySN0dRXoeujZ8JGDYjZnKHCXacz+lkP5NzMx7fQ6EXZIywxHxvDcJ/x+
lc0jyofXkgcNA1VpCZqLdXuwOQTJSvyOmVzBWNHhVRWPArw76bbOGdqQhKFsoSLwzMJXiw6VDbAn
nCE5VRWaYyEdTLkWUnXdlY6Ai6VDAJ9RJL1HlPrMLnlWRqO8Zux0g9eB6jdwLlN+0Kmw/LHxtVno
7331+eXNymWiPnWBt1cIj+AnDUuhxpyDnNDIRE+mlZ/v7geNHWIOjFQ8qxdtf4lIYptThQhCLOpY
caUcJipjOhG1gtIZ0JhG1tLxJHUSM5uQRqOolCyP3tCRof2EwrKiz8sX+AvSTpOAkD11rIBDG+2M
dBOKiSnFpP9UgQllVvm45+LYKmKNuFKFk7y+dGpbcJAc17OafKkIUqP+OspPvnV0/ZCqQZCjKqIE
jUif70wGN92CoHRlSJM24o//6XxbV+7AAUc1DRtpx9oAkgKJjEeMp++0yuYzg3BiHPEmLFzUnmxX
dFtkRBxzcp4o3uJBNLeVzoBAOSUVJD4lSH6pZZhOIgTmhIvogs/JvpxOUROysDgF9y5VJkHl0QTV
J8y7gl//+C9HrBW9YAi3FHK8bi0d38AvtjJqsCectBWWOkp7usIIRczrRpoFhOSgR+fzoFKq10mI
8Wk59p4QlyUSPb2vGqdB2lG1Dc1t3LonwIp4JPz1mzDIkyk369YwDsSEzHRrF87qaMW5TdTDXo+E
UD1R/2V9580dJtjHoaPtcwvBqdXtKbzgEojsHOyxwPebaMo0BQ6HlkNYDhvMAZduT23I7xTV3EjN
HTCVpV2OXYA5zA/bv2BoyyLqqoSQswnr5gJZqd3Ax8beL+yYdEA8cS84bO66HVjAdmKNPyXvYEHg
IC0m4trSxmXTsGcNPMahcfPk2U0cR66Fl6uwiL06sHxdo/ql6PxlRH689T1iHM6+VNfmohZ3kwyN
BZgEaPTsDRPihEWdtTgrlr3IeuIDHiFC5lB3CMoK7UNRf0iTnCPoKJ7YKSxbVbAPu7un375u6yae
szJni4WMWk8i7RuQ4O93FnSGMsXZWJreDOigUXFBmcd1Qzu50cVxaP8/hATe16GOvr5w0y43FAWo
SWBcGQwXYMBtYZmSmMuIwrLA+Th3HbIvxknpDhYwyUFyClTXkIqj7Kh91l14IDd981UKpsFNHR6D
eHwAdLWe2vulFYf/brYm9/ELoeYUBXAgaShrrFtYWxNBeUZ6Vn5H0dJvK1+iF1+Rh/BTAqnV/Mru
I0ud/ywoDNRIsOjoo8w9Vq+A43jZOcO2GYfv+PbeYUg7VTrNpiBV5iXwULWHHJbwuX861tvegzKG
DNxIXNGWkiYOoUz454gaCY70oMcke17NMC1TFCXZxwfJcVZP+0uKlrszKFnr1huSUjH44XwHCUjr
YBqvPJp8hTbkSY5t9BMtU61p/yTjOuGaCkg7q8raxNEN7Mv+WPgcNH5RxGfDOgek4tlV+eozapxR
nWXBC2lK3sWM9blrHoyI7rR6lnY/wTp0PmJpuSKjXM/jP2H9/ivxSYl/MDjlHF2ju5wvuqXEBocw
TqR4Q6OzWXBX3vFEUn0nj+ym85XH7GQRlKXL/E863zKrhI4Vl+AmUIFWXgW8WbovzKXH7UDz1Nrn
HfQXOjp9kQuOsfTOMWG4VTfwJ6ICHlndsuwOXFwLrTNv4QRdu0qVG7OqVSvBZMsH1FvtysEQak5q
aTYaS4rUiXjrl12cJhhM/Y/QvQ+1oWkQVde2cJXy4QZcaP9TUQyW6idZX23JgUMu4HoicJhik/zO
AtcWneWkY5j4gWNXIXyi01SCtdpUv+AjsVflOUc8AUQwGbdhyOpKU3OxkAs7rStKK503Yj+nflEj
gd0HqrTfX3JSyJCEcPozwJSAkNSTrXEwP+f21kpDwG4bWHQO7ZqZEU3vhB8vN8EEBW/6q11XCGCd
Ws7qpwJB74buVnRfDSjeOZD18s598r3qxLQwwegSH2qMti1XkIWCKb8VmFzSUKFoS/Rkx58K/eTT
ekEhB61D+7yfO8ucc5ApSqC/bLKkhx0cp+TntlF40pRIvrp0WaflQ263RG/gOdEoPa/i4PkrxtJq
x/edRA2zgPBvBE+SC/dIUhLUcuPwjTfq130ndTI7Vwu+Dao+pPNsGfmSlW0khexA/ljcsaE8B8kr
QMOQ9IDSPQcrdxzAn5FeVjTjL2+SCW7E+U9iO4Qrxf31ETOdUmrLEAXtzjtHwNQrkWjeNA//Epfo
IIjYpsztnJlxjZXqr0HSSFhSUZdfw60g7VCZ2OGkXgpgRteYhs6rmzsGO2x0W3X2zCKSyUwyEC3h
OBniripbYh3vk9bksVJ9O3IuXitdVwM5d5B7MO7MPOpvupIQhMa7LqG9RG2DT4Gx8lh3MWsxMRDt
WVwUaaVbFgDo+66TRQWWJRdk7IpVNXhr44JXh0NMk+vvmzmMie2UHo8SBJxQFHkqu2l5fGKKDMXx
NLxLuwYWxbpMO0R7RAU+hshu5YRHVQ9sH1XdGRDT0lWcPC++595xk+4ekA42YISevKr+0ou7K8KB
hI+vGptTYxtEOiHozcB+7uekL+X9GADzsJKmdzhJH0XoV162yJsr6nHXFkkkZ8NmhwC7rOHYv+zx
3Qwczt8Frlg3rLgpTc2qZBsBdGGIjFnps+o5/y50R9LFM11nzbQqj8rvaJiLQImqrAA8cWxhvNs3
Xa1hD6TJCyq3xUdIPWdTMf7OHx1uK0xHQZ0LJ7wyaQs8eblxPkhmIl73MYC0Y4n8el3c2MmSTu2V
VllcR7FFGQ81irU2TOhIqq/96IYjDnm8biuRfrGHozB7OCD/PPIB9t0cOGRa2p6phMHfNpS4iwUp
yekO5NvFs2q9xk5nRrWwQbi1LTCB0ReHb1ZDdiucLDiHUhTYTDrKsht8JvKecT/j+ndhGE/YaoGa
V4pkXi1QTwKwpDBYqDxY+6AIKgqZWrdHPph+4TWiktGFYwskpV43DDtSXFfuH4C8l8xoJVpsFLbx
AeOvNVeo0ByKhRDNF9IS2SrWiT+NUNpAwib9Xxtww/u3vWSXn389+9yvTu9gqPaGN5ek9imSqJA7
v88EOnHfE7svGoDDoEg66GVoJaQ90BX5xvjwmV13l9YjVQhoJRq1J8co7oqUPOzd9p8J/omx0sGB
zX7Lni32IfAMJiY6hg/mNRzlRFPdTuq1J5xPeYNUXpNZBOpetWBtDb4+TorJt2YteeBGRH8NP5Mb
7YOZGdf/9drPG3OD6I8ds8VVBfNMZqIlWNitj+GWOxebLRaTzK+pikhYOD8Iu5ik2I9OPO2RKzp6
d9tlRRdYPXyy//Ts/YjyFFvWhY7hoqwwoDON9NgG/NJarGxPpPqK/DpyNDAKhb6gO/9+ORWTQqzJ
4AnRujnFX7L0nL1PGN9zSSjFjq3ja8kQehu4uQ4iGcGAHyetI0FoksMJU0eCvl40wQea6HQnf2NS
wO/jQJ/xemLwxTEyGyBJdlecY66DovCySil1ODJWIxZFznnwo4/w/cM9ebL5CEqUpuW9p3nEUfTA
t5ZjFDBb3Ia4xhTPr6w+kOCDkDVNEPTD1ZGycx7ooRZnuMv9nZuQoFmKqAPb6oyp5VKUJu0yBUM8
Rx78b/3SeJxhW5KlHeJhMMc8KlZb1eJs6dDQ+0e8zqsYAbaSiWSDcVKTpjJ9BpsK5TgEnrDD7GIk
fj0geQ8i9gDVoniBF2Z9abA59kXojB/esBXCuLDcSn5fcxMPvC5s0pmGyjfBQ8AGU9lApxa8lnJi
DWggvFxVeKLG6tuhqQnfOTw1YtRAwRllKludFgQhk5MFhk9mX/igeUJ9qOyCXmlX14eRJMq8Bgqs
uEZjmD+N3xRiq4qREnMnmBO40mbIswqh48I460KlC0DO2cMP6OdI/El1h852mO+pZOyDd42F6dCc
X0R1pvOItMDONFiP1/k7QpKl7zaoPp2ePuUNT34attx67IA23WoiXdrYWltGwIJNKchFIMrNR8+O
1/twfW1Prs6PntDb1cQf0GKVk+iS9YR6molrrA7AI4m+PQSph8R/281XJ0Yg4yI/rEoarwUGiEFq
6wm6InjhklCdqZh5u+UJ/h8yvxcFPdnIHltBIAn2doyfzl0LEzj2e3y8UlShdwn/g/oG4nkCXj4w
G8uY29JyEfkenCn9VE0dkHPyOypNDgPLPS5aRZvpPT+ytmEsyoYSoLy9X1m7QfoGy4qZwhVoaDFx
4p+aQWoYmP+bS0SaCPmtP39np3ivFy1IJ11gIQSQoC5hWe/RzOc2boHH4/0gubi5Cb0LUI5XXQ9Z
DnePzQo/iZJKcQDKp3X/H1n/WywMlcpS4psDcorXGpHxBmYqUFWHh9hrQbEboSg6Mraify0f/SvV
E/4iHqkUEXp3yp4ctvcEWCkqzXV2p+zB2jI5wmbpANR2YniVenB/3KocuZmmIDQoTig0mE03VCyL
3u04mxW3S9k2EINcmqfrsByw0YQKllGQUY+3xTlPkBOmf0upbq+Z689Dqul9quZZYrL1m9gs+uVK
5wr3db+KhjAfEPt8X2b7XSado7PIOthbc0rztgDCRMGFZJ6zdOhoWOlOT6H1f2OAgf2MSrDjk+7m
m2tdSAzZvPMQeKZyamTGpDJ6N6jim/HeJ3K5g0KHa8cVPLfmYhSBgNZV4iTrE44sFfdH+CZcC4PR
RNQD4qZeqGrIWNs0/roDjAzp6gZYBHaLOcQbU/ddilZiS69ZD+ry6PdAkKpMDBN7WXtoajULLWly
j7kFdmV45/ZPDPgwHvejjtLnMipUpdseYXH1DBSFRb4sfdU+tIDMz+OkR2Lt1//c6ipdXWNTsB+f
x3ODSFKl0KpL96id0PZRfb8VojST+kDdPFnRGzoKcBSpF0HZt/IHcSKAGIlOLYZv6zn38trNr6VE
BnU9xWb8EiCpMm2nvW/xF+p5iDkkaAAU1mCxbydzfpfNLnif066EX5Vi2qS3Wi0KzQmXNcE5V7vh
vehepFDqfo7GrRl0VhYpJ8j3ntsO4IDQ0NEqlqfEQEbwKxggJ+Sdba8CBEzo22VtEksa2qOSqBHr
Rlq1UEzddZCbeI2Biwi+7DkkdP6HpKr3gxv+uaugEsIUmghaHjHtoQfi4QB/y0D8MfxR7NvxpGZL
byejugzrQMmYnskn6GurMvXyNWe6pxG0rCHcNtMGYWyTZhC4glKdbOFu0sQdtf3PS//LPkeZV4r0
FJyh/ENY6YSAMOj0UmaO5Fo7PWVF8krGBFt9JDrKYGEQez93HxweBVOUMEfnWEXvQXBxkDCRzxHe
oxdSn2yb0oJq9hQw/w68cy0hZfRH6IKmesXQyV4G568jexiXqpcPkZllpSz3i1LdzhXpSg+/pMEq
UTqli/AasrSXOQuIY8W7di2Afg2Fg8D3A8zeFjacKPgqxntCfJL/0gw2G3Ie9Q5Xi8jNIs9hUYqC
X9THF/PejbozBqgphKnMofLuO8111Gp0oPFp1gfhVC4T0Bvw+OYN240qhmXf3QVNspXyXH+UyPRN
ve61EeWC8PU2rqDq1STtiKjB6vq9zP1Kebpsy+RWhxAE8e/SJeRMqlhMHR94jpsoBAHexV8ac38V
hGVV1rlsEivyCJh+8IpylRHWkJk6GLtl1ua0UG9sRrpgIO0qTRdlTgjmKUpsMsHESWQ85Q+t+gpN
j1S6cOqQWstTaLOz1yDRrJTv1c8GMGGH8tkcjzs1rPuuha1eswqnlO8F8jkBIN+dhPsJ5QArHrlk
Ymgcobc7OBdROooR7LQNW6aICrJpKKP3MXk0wZ7SD3QXzV1JrJ8hO354IU83cXaHyMaJyTvIqnaV
0NA39QmerNVfYjjhCgUaVHVTd0hVw7Sx3gSVLKIPeAAFDlcPCOMNsUsFE68pO3gMfmTxRhcdrzZz
x5LmocQZ5eS6NNnAx8FgOusMvLOefuL+Ul3oQev2WPZc8QlkhPOdM3QRT0Zy6dM+JmTU+Hh2j3Fp
Ota34ugX26QbvGPhcQUFjxa1Et2+Mrvwm1ESdbv2/D7cSZV2dfBd6nQVa2IqUfpuA/xCzYdEwQ+s
auBhuBBT2cldEgJcc4phmf0NlfhnGPAE9BqC1bJrqY0amXCL8uKcV6vjqKd4yct3TAZgWKnhbKP4
3AnUJxvvBwIlrED+aa4OjOglXps1sq34LN1a/3F3JeIbu0VJWMzacs2kkrRoFJV6FBoE22XoHJda
+kbo7pcfr1NNE5og6dDQ7sMCCHZp0V3fntjoPpeOR77OjfgJsatwvIhI7Vb5QWk/5yGCtIaEjhqN
ci2+1vDVVg5tY1FqS/m3CaGG+BPppATxRL/gu6Oht+u0fGdjyKrMWiiWKjhsjOh5s0KNwSFrPM+/
S/9SUNy2DyiaOD4l3Kgn02KWcnNT0G6fJF2gQ+GCTaAMyNzQwC+7lxlMm3FpxPVmzYdoaRETDCxU
3lXj3877D02PS345qGAOHLPaBGHfgnIR5pis3lZ3if51hNpf5Kua8vtvzEiY/lbyoKCXWrpFDbA8
NhEpIYBvKEdEHmXluloeHS2qDBy/WigyaxvK2zqErw/ficktTQXhp4cyXaV/WetHBiUNnB48KxZb
Dbev17H9RhxxIn1CTbjUqV3mcSJ/mIhWIFOppte4RX2Jks/Sc2OimMsCCiZjsh60WmhC1fxF9Vp0
rvKpZNy+SWz/wZPTDHiPMXqaGdi6/lyWSVVjFQLKhrQ5y5pxcdQzZ1wA52sZg2NITF3O3eKZ8G4d
MFxyZe5+6gyMbAkyK2Pp4PHYxc/ADjiLICKS6RGlE1VkyFSAqdMHpp8cFJ247mmEu/QmMaVcKB38
GjEoGoeeBUDuhrMTHg/OIc+7ubFRItGxcbKn4KjzfP8usMa7GJXlNlvr/UWmKWRghOxgrp9UNzcK
NQLLngSX6yUGbyIPEx3y+SSZLKjk0/Q8LmesAGS/2CHCF5sUl4GWTBpCd8RCFoPPLal0POx+pfFy
dAH/00pV2B90pRUp7pdz4OISyOaIeBIvJ6JSLGr7QGgtUiHbegB0cK08CQ07FuYYCLBFAxm2Yz8w
fxWKqGPsu5u09S8sD2JCaAak3xe73hcYWVDJ7W4JafdtT80B3z7NO4sHA6cfiN52hLApkfXZbcbD
//5kpvVpUXh7nICAn2pzCzTk6FAswGt6MUfX1I6LIg1i8QH725ho7twJLj1UD6tzhAXlRsxvbsrl
lPKGhkzC+d1I8aq7FYQOBA+U0M3YoeaIHmN42ymiPO7hdSXe09XeFp1ef/OreRMeu5ncutdnrCyV
1mlyU6PRHyE2pD3ZJKGOnuMJlXT9NjFNDtD98aZunmJtJW+lP3fVgB42QUnIocEyp+IIZSyQpMFC
a82q7f3k/kn1SaqhB7/+Vp5QVRGZWSl08Pdb4J5/l16O0OzAh/XxXfmBzYMHC1JhUnmN4UiO1hfc
9AmTutXCoHE3xX6jBSe+iku//axmNUuVv/DsWk5ue1gAx9Av/bWJtF2CXmkl4tUkz+wvSeGHMwk2
S7EgfFlTP6dzfSTWVD1abiNonflAvl60Mb04e2mP4gE8mgoXrOBMlWGUdLM07vW1wtte6uSehzqd
g2SxeNWxZ9Hy527fvJc1+UF53mfv8h6f7axEHpkRfyVShfYZmUPqprWPkYZo6sayMFqtLwfcRd9Q
WSaE/O44OzZVb+ArIG5pd9CfWMTLmzm5sotp5zwro+kbq8VFpuTgq3rQqsRcI7x6iSXrIXZk5I9m
BZarCYhvuZZIBWd30BAmMkw+/8i7iH3OFyP21XhmOL2k9u6cFXNWuNIWe0QdL/FL+LJz4Bpu7/Hd
7EmMK12eDOADjzd4dCwfeAY3YyvPl43Q+cyDEM3Sme9f3fhT79xnFivMZf5wCU/xDSdA1RODizri
tcWc1hIxNljxb4C0h2NzGSY94TzUsM+/FwMJcjci8Pv3mW9zTd29LoPQjf7N947jwBz4q6LTIl07
rXtHT11YcgmnU1ofmEvysX6+BmgAQTg3fYKVekbPjQYPKKy2Z1tFk0dsMdINL16d/IZxiMGKWAf9
vi0VHisEIc00GQfVeN1ihCvKkcMGen7f3ie1o4VQ60is0tjP2YdXJgp2ZTH6Tq7Aly3mIa55/03G
KCKp+1Mnz7yThvI+bDTToyr9AT0sVyB5Zbe3IdDqCKXxC821SzMkXcY/JOfDEsajp7K0qvJwp1Op
OX1yQPtlC67g39qQi3rd1KTPihD346z1FQglmqfWrZkIzMJ3FGb9x2TssrzLAiS0WvHZnegepEBF
eJJch9MK7eU3m9udpGZoUMpZcoBOqMDYRONRK0px78SuH5/YtqkSGc9wuZ1/7IECpGSRAB43VQpL
AZm8QicqikK82PpCJoOJsAilWEReuN5Nf+fDSTo0vJiHWEUBHV9b11zJatgP6AB98ZAnCLdpr+cK
i070ubq46qYH8YDpa98x4x8zGqsCpebKTCofCOJ6K03SlnF1/WexOtDw4l7fAVIrHIl0s2jzUaqg
lov5l2zaFQ5odpU6HkKb6VAqcoKGwhK0M3TRt6/wp9+eYnSMOGO3ldZZ92Cpk3T4MrEv2xE+cNGU
vWKqeQ6fQkAqFYGvnpR3aHbmutaJNB7uLAaodrfxW+Hkvy0t4xCSxoHs2o9CqHntLcdyq4UEDmLW
y+aW0m3TMCcMiobJmVim+LHbfU5dx94NeHD7B6Fbwab8v8PSiOfnkj74Oo3eKmrCBOW9e4jRWwdW
RwLDhx4L9QISFMXx0UwpRQiNjnaU5Mao6SOZtB5HUfsRG9nEs90X8p2L3i3VwFAz69e5Fcu+mt2p
Ae+wkGjCxCZQCn1UiygJ9XTOYEm+lK1189kIKQRfwKCnfDZbVbuVftjBlYkmtvto81b6He5G78y7
UCmdwv+4hvPVGyJJXySPl3HBuFyDynOeFIoLf6xuQgduEvMRBqejbFcC+/m1nij+NdGB/0RXNluY
0fzS+vL7WhJKcXJ9qc2NepK+N6AfMSH9c6+LjmqIdRs/o+zYrRylRUySbLohZ+/eCjfsZM06qYYO
r//Pq1qnKSqYqv+wGbYx6eMVHmaYNoCeyjO947Y6nw/Khfx40M5p958XXrbiASVfj7Rti8lQGcgY
dpNG+8ox89HXxbZaFfDQAqX1Fe4eBn+Dld5Wli2p/1/9Gkj8eaP/4nw9eu4yERHMCRUP6iZK7iGT
1xrK2oA25LyDiz8fH8i+crMiH9IKW//8gC609gL/t7yNMc2s4XjSK9++qRLfrCfjUIjbWNrSjKFM
7QRIPWGNZ9a2BzzpXOZDJCVKt6t7IXp9CDLww5gX5TZ7aUThPwV7OchMqmwUcfBci/VHaehqcs+e
tIgFw14XBsR7RY6WSDK701jQok7MwLsjYHzzJlLNtxwq6ILLrYKSzoTttthEdv3vaXmxh8cIWZu2
WB3hu0AUUzDBWaBkj7H3aAwxam/Gz/Of55Ua1RCriTp0yydBOfKe135iZ1BYhkMbZCwXM5BKqdS9
Pydrrx1W3ClqqnlaVW/vfXWqaWmpTUCpGQc+CcY42NZxn5BcRrzNC6IkYbSZ7h/0kvGdZxlNWB/+
m8FQUbogMBHQRpEerXUBlYzbcSGYrrtX7abpoJ99B0TQeb5/L5L/RQZEpe2Zk+yF34cFDNO+G138
TamPIW1MrvGggIhQHvndxkFtU7NumvxiYFsViI9EahJDseFgflnqZyjDcpPPzIDwPVE7Hf6hfngY
awkkBPgIqIll8b5UqD6GfR2++GewSZxPqQbn8NfT6jh2EwgkBhmUFwRuh2aNbsnZPBIbVkQr8mTe
xbsvHesBU/RL3QjbPgU+gJVaqmqP9fB6beGP81gasmylHA6zrNuUS1PSNtDoqiVAgG5fjWeZL6gM
149ca6R0i8+mSXyyuQ+isSLvKYDrBS6j+HGvE1Qf+QKqTI4aB2WQSKVDTvj6+zeL0njG0Rdouxiu
DpPi+4B6WdV9Rw0aITG8RAPmazEOuOsWx6VqBVAMsa9uJE3WNuIwC/yI5NqnAf2Ys9cwcRlL50wn
5v/9grbJBzCIjT3PHvIkwvW4/lTaeAHDYb/letN6wVBR4uoxoj/QT6o0daTGhn6DDS9JrY9QTqPK
zklok+k42hMGjyPKMQ3+H+t1MW8PuD5C/LC2vG35T9n/jt4GxthkOqcdAmNuOpfUIR2jlGn2GD/a
eo2gQAsP/1ppm0PViEZN0gQw2gTcYjyU1BArmAs6t9CiqedBReOShRw98vy7VLVLD9LonYs7q2CL
z+Ej/Z3revzFPSXD4de+QoQwGVLWpOHDWOcSlUr7AgSxpfbbX1bkzFrbgm5RIzhdkiCi5g9pBwwS
gb6siAeMCMDjQQGLdIGFgK+v9Shb6ac+JQLEkmeGsRWil52yIE4sms///vHg11TEXnJnu0m+g7vV
EBp8ZcDjIsJRYiQA5l2TKyxraR9n0U87KwcJaCT1M8KJKNYbYX4SzlzCHi3F6/fT7AXnGRJHS0xd
0lSGNSYuk0RK0cyqywXh5p3fbhBDRk9pUTIY1ZPQhs1tQa7JCZEBlr6xvWyioURGz01tcpN9V24t
83eTUuiijb7Njrig9/1UhfSet3UN/HixmNw8Lwfw4ux2aRfMr3SmEZQJCLLgyL1cbKXDSiKzmRbd
dAXR1uS+Af7edh2U3OVjS+S3vD+RJKb4qWhDtY2X5qUkF5p4V3DRFZdXRsricRA5upiLcHjRghmP
3VcJXRaCM43GfV5MRpCBZBiHFw9T8aMeIDfZan5694jAoPg65OS8cyPsmebETem/CUSSzv8qtfZK
1+h5eWYU8P3BHqYZjlVbUBzaDyuGUM7gt3Nze1M/KhF21zoRCr+EKpgn2jdq23nPyHS2ATieEuWQ
meHj7CVPwvRZ/1fXBLrCNfYTuFgMfEKaFsHbVcOgkeBHKwlIhbixS9dMHMH30lMoRTG/DDgPTKHu
PTerwwEYoMB/GpbnW3eQvWI8yp+Haf4pUe74jZIDJbY8vujNYqZONJ+whctDtuYn3rFLRTXzeBGB
1x/wMjQZ27CjHprfMxFRTMy92MmI3EaDJOn1L2FxsMkjj2JBSouOLxA7TyhSHO8/nXjRU6T2D14R
MvwLEA0bDccZ03NnLrmLxy8O4sExLNnmtlUxR6E2ONmhQYMbx9l/czIkKeYVJ1FUnCA1fhVeOayt
DxiOgz9kKyues4b9uh2VKy6IVH51NtEXYpXNmHQvy3IG/7BmhaFNlyu1FLiCPV5qQMksQ3HJJPAF
3d0hcNo6GSVfGWwUF+gv/8cM+QRfnNFXJA6skLUS+ffqVGzQ9VlU6Br6wN51oznzR2yDF9Im+nvX
zHWqyHrP4sGVBDfqzut29BHK7lkPzgcZxZMa2VqZXRtxGsFyZ8zo0rKRNBUw2a0qy+O+ioItSOU1
oQAVlk19TiLsF0Mthpx/VFGKkXwALsS9rU+zdb8nSLfAopQalD9NFo9sjy37xM5XBMd+moCMgByP
B/W6nqueWVnRGKGn1wdnDH/2peGakUbE4XWQxGBodsvGuAA5mR5sarP2T1do1jwv7U45plj1hg6s
WE4nK+DsWFJ+vE15l7+CWZ+iW34h9PWGjMM70KFamL9KGQV2PshLw4DYL5c+upiP4i2im4DdKWHl
2MkmblGtgdLl33k2PGL9qZXXrpz6qGtMGrBHVQCO2qj29Whs+14m5OedMMC2+BT4nbr8rCfFXMHk
vq2N4kKJAoUY3XhtMigNYORjngBYD5fbwtTBObGCFfeMPReaLI1YM0pZ0xLfA1apavza3CKIapyF
ByGualbrugElbBUaCiP3eCSsvfx7RQiJcBPoAMEUJkxt8/ntAzoGhEIN55gHfk3tQJHXbHfAGULo
CSNtyiLHIV0voyNEHI+ELZYiEPQzVWu1JNP+EilaWKydhHSO9b/SzXjSRgQJpecyJPUvlqHuqFcs
09KHouT5jP0I25Vzwj5HOKVePzytClZ6A8jSimJ0a6xzolBGhdueKRxWXx41m9dM2NQuMiPIFnT2
umwsXorwQLJQ2nqIAL+QumR0+2tRQW/vykyGr+hMcb1cViai4qZfP+AFLjdZeR9GM3vF53Q7Z+WY
J4A4dHX4q/p8I1ozna80j5AGO4VD1opFwspq8zA9qGGvjeWfuiRovfWXyFyfCFu0N3iOmvoscvLd
3aNr9lywcOUcOTbhzGxM1PZe9uiGWI1Ssm5WostjnBR62lvnysebaBacL4EXHD08dyhEqNUPprir
IAKXhJODyKY7eKbRtjNZf6AoxH2r38/KwOIZ/bnfTDDflsvzXXoZNXCwmWA2XtXzEzwrPotwySoZ
+SwboZz2DzdIpEqamJcXg5XJpZW3mBuEbTzjeQ2E9Q07FiVWWxmcMZZbmExW/vYYgHIS/gW67nHA
UlAUgbQOl141F992ldzIySf4drsNtx7lEHmtNUF00c8N1F5Z3LB02qwn9UDMqFR/LJR6qiki+Ddh
iYVXRJX0wwGUCtpRdWc4i9sudEj1zlmqO0tW3gPaxvp9aS1eUXfWvM9P8Ik7uj/yBQoUNOOvZp8S
I+tiP5lZfKgarVEEMO2+nqAl0DMzdzhuMXYctPKy/e+vCg8RsQ9SyFjgllt03a1e2k7AMYjVvfEE
7NcVmKIA+Gbev59nJtTfxHHJCOGSyu0H6Wy0gwEbnoRNl0/38QV85AdflNHiTrigf9k2ThAYzrPz
wgkjXWEHQnbJzKPS5uCQLUFbtHtszetYMg5hMZWMgWsRbry7CreQyEmbJGhATvJjvz0zPIIuZxeq
wsHJiaNCPOfIQqYKKzgPmRWa7AcSw9CvbG98G1UOs0tv/1Y20VSrymGCCEygSVBoxkx8msObU+TJ
qlCtj4UlGksEU7w6Q78wW85+XoCiJ5jkcGhjJ4qxXKtn0NPZK/QnGJgSMxk3uXcYfNdhJi6hsSZn
VCSnjVEqm0yups8yXxW5HzKxd6Sf3kaLFzd0EgRfHj0KoaQeFouj0Jsh+oJSkDkcd282yUOaC66j
1g/uF9XOswLWRPPFy1De9N57wwtkP31fj4MbYtRrhi7IamK+1dPffpbXF6HeLFjPLybwiJpidFB9
WPrJEL5DWk+xBLA2QBFb7+nsMmi24Lw3s2INn39eNz27b8KG+FAxEpwyEM7sLwTkeibcVv59agaz
RZ0hbjgGG2F2A4b8CcvMBIKikFLsCPuXo336O/+/SbgPTwDut0ppc0lXKawKbGP67hLEQpNyy1gS
6MTcIVWHWM6861uJ9Xj3i/zQr44P66NTZ/5vDtg6KcjDtw3vtFEZ1mc7vFkX7FIJjL+Av0qmsZg+
iNyH661bwiXNu44Dqwsn1x9zInwJII1gHSepFWX8oHKlwmJswqm1hwGyZx3gctoMpQ69G0th4k0H
Wc3QQBNBujCv4LcuaerESXom+ts71hB7L9/YnDGCOjSDQ+tQvRWi9TjFTNqQ5nmn+OK/niK62vBq
VaJkKqW9vZp1Xg+CzOj+nz8fTkvIlKpllGqybHk9xpinhwVhYfrtQ3HPnpXDTHZfd8SoD3qXDhBb
JsMeabR5SleLXSAimYaKRYba0Bq+AYp3wQsMxkHAFlGB11GC9SHJ937TieKaUpkF+frLRX39WpXY
RY6C1OBOQa+xISp2KV185hQq4D6dnBeYTJESD7dS766RyoP+4tapXwASPVXxUVL1helnmxqQZBHX
JaKRIlgqYSE4NKPpRMFeGlGOnySm40/GFzn6DvzHgFPskV04FmDwLkQGxGOwl/Ewzv7CydL8ZXQ0
5+Dq5DyjCeiwbQrEhcQ5KLDMQ0hiFzSHchYxi5u/2sl9xH946agqV0Khngl+JdAwz2IQXCoBPcdg
beCwyED5HNjhjxo+T4M3QqpErohDB74L2oQrgM+78IH3FMrfTaRuPzz1P4zFDCcM4l7pxcsR3a+e
gpP1zODZiZA3dk+apN+j0pt1HjBVNRnRgILicJDJIG93/fCpr7sz0acFpuBip3kt8kMiqep5qAra
pWaMKFKCl6MzIbU6QGsUyC8Qk36AkhNAnCMsvuePwdHVICGXFwzJV2YEmirVNFd5pd5zRXHw7VzR
n+lGIBxUJjgJI37EA7pOTdC9MfM8Bu4n3tyPf/mk4x/AsZoVKk5v1Nd5gqHSAQrt0os1ku9XPEjh
nQKUVBq1j6EtaEOst8RZERNShz2SFWY88g011FRKL4O3lBYr0ffbcOwQdZarxhIfIMOnW3SpiGzj
VjgP1a9DfhcMYE5tYVeT8liZ9wz5FJwW6wgGAXeedKLmwGIKaryMXHxbW+TsD5M5Eo2frmMyjKUy
w9RdsJ+yfO+yIUeZIXRC02F+txloNaWc3iW06wJOZbyeviNqKXpaqaYFtCaE4hrD4YWxuj7/hk8E
wxkFWGVj1PTdLxi/2PZcYpisITh3Hfqy/rtxazszRsuWTAgGbfxiqKSiBARIqisd/s8Xw+95jJlj
KYHR/leSMNiXMIdvT6LnKKO2PJRbHgNODE38vbCkYTWxlzSecS+vCuWMFKOtOv+VsBLUSd1XYHnL
TSdvFDHBq9eRJ8bkrwFC67kW89IDRfumDqEbr6m842lpmvl+AJsA1pq0+54sISDprX34q/X4SBYz
zsjjBcah/c9vnIdbvp7I7wUn6PtXqKzDcF+5X5uk+25UVejOBm5YdxOFYg11xPFmylpUg4Mw4+i7
enL20jIO7ir/KIZ5JiJqgSuUOX0dEUPAmJ07xSEWANFbNwRcRuuep7TM23+5WWvn4hiT8eoffShk
4ZNvIEKIpNL0NQCthHrCDNwThdyzcV5ZbCry8oHLBFDsDwP1BelggwHKnow/acBYQtsUPksQC+7Y
H3ZN0VajsuU85CPmkV1YYZm19eeGEQ77F97300Zl47bjn8tW8C7BMutHGXOH9ZBbZDNwUj9GTvma
AK1DH6lySQva95oqgGuSauJvyW+4kd406oObGD+U9rrYTgqC6Kj6G3Klrz8oODwdBTZfEFieDT64
oCVWCXoMsEQDEi44MWFlbTTQNF2a3+7slRxhvO23j1xII6tGuFw1CZxAM0TLg8P1eUj19gxgeABe
CnVcyUOHRDJiD7FBdm6VQRraIO6ZR47mA/P+l6rl9OrGO7g+uSx7GlKBfxrzc22Prl6mzvJaDT4n
KP8eupUvrVZ2E3vdwExiJvvz7tyJ5J5j13Ygp5TfL1Ws9UWDdpBc47nZUGJH5PHIFs+Cv2lRIPKb
8yrAH+HsjhgcdQ2SytnjDf8joaBgd84GNNupl/KoiyDJsirq2lFsMl4fUJVTKJXcyole9LaZaxP3
+psYaoiSGeuXWLHOF9eYVLG2ePWiC5sPQNqil2AmP2/A8Og4fJEVMMLUO63HE8/JEWAhwmlqe30G
XYULZOEbESZF0bQi6fH5ijZXcDCS7CTME0IBgYyJEu7f5qGqRAdJUH5Ni/OUwUa9kQI8sAM+2Z0U
Zyi4S0RC96nzBNcNMJITI/M9tWCSV1TxUuJDvGA8Dowvx8ITPsz9KvxfU7HUj6Dzsw0sxmMqneZg
v94XzWs5rFr5lQOqoao+i/I3QqykqkqpGFiulpC3wVtoEtrhi9P1F5GI6I5HZc0AdYKwelehWVUf
psMPIEfAiojqsXCLfB0LfAFm2wOLGer2P7VolL/GwoMKWnPgSsOM3jp4mQIBDR+tiGlstOuR1uJJ
iBvwx173rjmSGwkWSmC2rZXP67wG+s4G1fcpXisrT4duZe5VszfZ6k/dqJm3ZO77mwS3vKrGRQop
5OP4y5+9obhkN65ebL+WLZBcx+1m2DHjHOGNTfufjQefnsQ3lIpBLqSPlb/5uAgcIv7V1KZHb94R
CWYf0Zl0kj/7K1WEsn4CQ8R3iSaXyrCSyBc4/66Xb0zpRmYFFuKsySxrKbx498bfui5dvaIW26xN
dFBQS/oZ0Res972/fG6li8sPItlvXpkrOcvDp0wJeJn+5DU3HHN+ucfLhD8ryNGj4j9aDst05n29
ILDdTycw0GK2XLfMBwVNU7iDWC2R5h/7GqqsKH7+gLD/Y5L2/J/ZqwyY6UJyqFHnIASZLPXpP77s
EPGxgF6YnCfyMf4yej8sa/3RCSgwRAsfGYyRt9CAPGUQDsGhRdjaN1Rcc+A57WEeFCkx8e9zD609
PaN+c8wuoVNHU91Pf9IbEEYLf0f802MnbTJyA4rqJe0kZkYTd1GlGxZUQhMMSstYfhlS8uf06rFP
6vYKPYwuPfY/3wk3KNoG13urz/CCgnhbjrShxn5FLnTOq2S6HHtSYUPoMCokwDxvIXP+3UtZfdHv
pfQZFvhlXdVegJfrn2B8oShq86jIXg1BtrqHs56PHfl2WQQksYTrKmj25xG07T52HrOQ9LQQx++B
arTw6LnMr3rOeD1lCLIwaGP662yaZxDj7OgASNji9j+mE2f7CuQEum027oPScOhflSrKoZRVz2Lc
r029a0fRaJh3Bb2lhtTM1r7MGLd3iJVxMuluy97OFBLE8WLMyW86yU87Rti4bfSlaIhvnPuaYM7l
qY4fqh4r2MKyINGuzGBCNZPC2n3sxiRPEluWzKZ/PVIaQhHRRK22HpYCEZoUZT49XYH7rVAIGyKw
YDvYy4pV0hds8kQkM4++578JKdsA3HA8zCCX4Hm7mGE9a+9a7WOH8WIdhx/7OEmlgg4ZXZjbjqrZ
FzB7UAebdgc1SJQNtHMWL9LhieyAaC2fsLj9rWaPVlyJ23XgEHzVv0p/yjVTLSaSjGAL41HKOxSl
+An4BpO7qaIKVoOWkkLZ9Q1SzHy3t130Aoop10O5+LdYkSjepJNixS8HxEe+P/5UCOjEPDmBRpmz
aa6EU6+lmuzHXngP145LNb57a1/g5k+zlj+MDv1+TelXnPWii5RBipfEpI9npWvjweGocV9h+uew
MEBt9hDk/Dd3ebEIZ6P/W59knupgzLeqDEaaIphEcTTjf0dLhVtVJQi8xMnoqd0LCrnnT58ru5Fc
YasKMiLd5Qg/bcoeRSF/9/pnXYlRGmDvcdpdj6oBs1XCvJy2i6heWED9F544cGR6EnsjIHzN6Ij8
S0EtbuAibS74Xw6VP8S3vk8pbB66VxUOSPTm/CdBcDvRwDOKlQDQiK6EaQN/sVWsVuY7c3X2/YWS
6mx2LjPmDDOl3lLy5H5qyaeJHcbvP7cXN0GhK3N9reGhyUcG0B7RXjnzOfIyfO5/MyGBQK6cz7zt
Z3keylgl4oPktfLdflWjfrrQEwP8h8Kc2aSqGZGgOmmcFIOeU2gos+47hjC1KyxIyGfnOZLgOZgp
Ty4xuNSYXVeYCWVXYQBjMXh8PmHSwT3YUOU/zyi8+viAICNNLIYGoi52bSl+/lyr8kZaFxP2Vzz/
jm/5d3hesbwkXsPQwxQiBYFOiJnfsggA0N/tR8ZBhBiZY4DioRn/YfgP/8gcC2htp899SbbFJjXV
jm95P0eKdGjtOow0aJJGySJEikMuUEAc0WMUoi2kUJCy1gMdEt4+5CX8zxKYEs27uKAHhqKaoz4Y
+H+9zCG3eayyqjy2jFgDF6VL/Lc7sMfsgC+I78D7IO9iQCJrwzeLvHMl9cFYc/01Td68Hbjj/Crl
aW2nljEYhvtAPfvhk81okf/Ui6hWOFapWjRYwf4Lp3pDsQmh2UumCZWKq52xE4VafusppKxB26Dh
fwSdh7Xyp05Aqr0zw9zVIc2fiAhd0VvRwgThYicPfp1xALCHtTd4mSHJr6n3XgOYeBYsMnSmj9Uw
YJ6j9ydNL44nOrXCOjCzf1A1LFaBoyVGo2XpnEVfnwmnXySqUmP5DoeUz5SDbYvUwOzxb8RCHj/W
ShRxUkdWsASAFwiJWg3HVBjF/I4/YRNi+OkzhsksGe/mFHttvs3DR4lYNtCvir2xCLJqd8PHpYVJ
VdqMz7EgjvhFFjKaxvLoEyxwY+R5oKHcbGqrBFQj0ye8DuDRUKd+l5dys7tp/5Zor6pwpBNpfRhZ
YB8fx1H0SGy15w3FXPhOcuAASG6YeTDmOENB6RcLaijt2nqfkF5ZFIaroH1ysAtRxZDpLHWU1Jxv
rGnZ5HUlDCtZ+ZYkAFmHLiD7DmA6rhEQqtK734KjwzpIYA6K43GR0U7J7uEo1Pfi38wWm24ZZgqp
8YmgpyL9XFqAM8SLdWy5kNPRORLDiyvoK/hS/V4AyivU77S92JIvS+W6tBtip29UleSUFbxhfDZf
TgFpDTx4grGggq1DA9LadZP860UesatWjs/FG2hKFpkl2Mlhj9hBhTALw/Gh+0/1xq2EoFW5U4G8
Ck/PH49y/1If5clceXwj4K0D+YX4jHnbF1+99or1PS1tAz0VkLAVeTmDMJntXM0PZiV1WqtUWssN
L9lTj711YCWcOYXXOFinAshGdH31mcSbPe0DbYA00Ys0GxlvM8BMVdNqI8v0U2oqDqtZZcv0ypeS
m89nT7v356MQxZn/dAnCFxdtlLAYHkdduyLNZvgeJpb3QO5avSfpsa9vyN205QiH/GeUJrhy7mlB
y2jBlvkyIbCU+Z050BkdPyo9RBKFq+ul0aQLv3WVfWMGcTrXEaz7GW0fbO1V1G1HBrkZJ8ohMYVK
bg9LpuvFLU4TQsYSRNBh2wIDwWyPWs0+ZmN3ibvUYda+hgpV99gQfAb7GCDRAYqggrwmYobq2uv3
2EE0A1vE25YTHKyd5LI0xJZdnykmc+ZEXXIFP11L3uPZ8Mk1zWpy92WBq8tJbUiC0OTmWwxrhLe3
8cwwvmrHMt74kH4ByKR8EuAPg02Qqks/56gtij+iiYngh2zZTCmvXSQ2OSIl5v3BEHwgdQkFqQma
uVJ8ZhgkCSLSvVwvk7MgR2xC03kKYfwat93CIE1dwE9ENyooR7Mt0XFGFkJ8W2YHCzaxJQT5Y+SZ
REiteEK93D7GT6SceU+gTqjCEvccmV7rpOgL7+94pKx4H6ebDb5QKKoTgFDp8dPgeHq42IyQ60gR
SpQhMwK9Nzi5k/bisifV8pxKKJFEgdI6EUWa80EvEy9tsRVOpzVJLLI6NU/Lyh58VDSvdQrH7GHZ
n5URjDrqaBVVmm9v0vHTBkD37lZ7vxZqcnja7bFSmjGS7t2DLjEgLj2u5a7p+LObZ8q+PYBWq+bw
P9bE9Nm9EpczTKode7p+lw9T0NHYMwHhhmPqOVABpq8LUvTxn2qcKNRDxKhUNhbBN4NmmBJxYJ2r
LXvgt2SajJMdSvUSpfj5cwfsoGyzkrW61uSUXJtz66zDy08b9HwsXCN7OwyAzQFW08rO8qucXa7l
V/UGmXfnveI/4sUZpHSBJQDWWnGc9u/lxfKoZfqr7ODAx36C7/c7xuvny9kUX/wGhiGWsVEKAiU2
dNQwDZh6wKY2k9Sl5RCSAv57/27E3xwhrogV9lDDufVYzUqxljHazHD6G7tkl2vRK+qmPN4HuqnW
yG2PKr8Y8ji2vmIKB+tMp/Sx1YJv50Z/SC/zha/GMco8iDV1EbUZo+GnDPqkri0ILbs179sZiyHv
w5cMhk4ywL2imLOHKWIdmFOZpqF8/0VfE64uD6YV7UOVho5xw2fB66I+oks1d2K3byNRD45tV9DD
QIXu+L6tQQJ2oaqxbnuq96AlBZIaFlHJNnde5w81KY3soaxAYG1T+rKX6QtB48VL/zYcf9u1ttAr
m6t+3SjrlVS+RAEuDP+TYrIlKYratUdk3rK4V+h6sDzEJDjaUCu9Pq784SoV3DTNP3JiOqG2tMwR
q7leqtFDOQPNGvKLAh5VTKJctFMRz5gbjOB/2UCHuriRLmB6iLuvvpH9Nw6eMPilOBhq/eRCu56y
dx3LcUVq6SDTbTZv7PdSxL81Ce1cS8AluflPFB+JwRp4yWp6QjKClbdvLfJueIbLbw7SnuJsHLHq
6Ll8lXYvVP5IbQR8w68yuC+WzE0Es/EF2MD17uGNYrx+8oRWu/srxrXYZaTGoHM1ZrHf1Ld0LdOE
Sl3L/kpDcpFK5pzB9gX87qc9JRyplELtjTtaKLiHOsqS4OpL5VrVP4xIZFo5hQpBLnhysHvhkA58
AIIq1wYB+7xbYxh9BktyZGaNrqKkYhMbBYVGYlf8f9XvnoX/I8ZX/mb87plJirqCOHI3ZOd6GbjH
8f/ojE3oUrFcUjEUXkT9MV3XISECQyhvwZt002QLNuiLGpV93Wat+R1hSgVkY9nzankGKqIV34/8
FHpu7ZYcU9zEV6S+8zcFz8xb8V9N94ny2o5NM90m2iPUdVi4jRh8GRFjyAExLGHdsdFhqRzO5wzQ
D3bq+h6oxat0+NgQcBOgN1BJQXLvipa6fj/2c41VN2FnsFVjrsGZbFFfR/LdrlZsomKFTD2nbjBu
uqWMrgkmSSZFyvbKta7NMfM7du78Jxcde+C1aJwTLwErRRN4MvsFw448tm8yR2JEjulksK1Rf24n
kZXeHwT7hzk5OirPWQfaFB+grwyeHGmtwFEi+wMAFMUCFWnaEtFSwq4+xBLYJLVYpkY5dhaHKwVG
6zGDnjf9iEt+7gi/xrfrwY4MZvvlJB/z8iUWE10vYhGcX/56rdMTxb9NIGsN8Fc3Ik9IWuR/0bXw
rYDhFq1CGTjI5CLSAgFCIcU00ProfSUmToC0t+QKx44kq0KTgXVP/y6mh6J1EfW41V9JZ+tNpRb5
iWHFnZCRhBTSYE0ThcWPFYikkLo+VsjEiwC99JEK7JVltiQeSe7UmpDsg+e/MJ80snZD+8CSMHH0
eK0Qc/HNv5FdWRBDUvnfkDr4XBOgwERfyzS81Xt9/T4vmch/VwmbcJDGo0zG+WhLy1QdXpiMjwAZ
vD8XFCEuLB5vSIkfYwWGqHaz0yH4KMA7awUR/rI6xp0gC1fho5gLZWck9iFApIVP+qweDCSugXbk
eJLrnVPF6xcIF3x4Kfp3zh4StqVwEgbhI+M7zGfgTFhaKg5iRzIYZGJ1yKOuZBxL5uDSLZ9Wx50M
/JK8fHkDRqHobMmJecWu2shy8nJWQITv2aqHX4tDxl0r1slUUmZvQKVuO53Fqcwvn89ueEBD6jMn
Dy+MbtY/n667zeUakB8u9Jq2NxXiGf0rBdodU9Ok9QRxnOLmoZbvbjMY5qSoqixxwcIfQAc39Bob
bAXVnS1+76N5jwYPXbR3Fi9ocThFtJEw1xETjIpEm7aVILGd6LSM6P85/XYD4HFIEuPSaVJ9s2AD
duxbZtXkItpEKcls6yOSmUsXZXXSNuFi7IFr7/TrBE26e6mVVht6jEyEs7AMLvpu9NSdrVvOYqMt
Cl9/7z0NfGF1O9w9RqMwxWTSrkq1PlTcuLObGqJUGNNOeIXXL2yMC1Aj+Q/144ZL6XNUIt3pMc2/
tly+VvxHzZHulcnTmK22YXOs3qW6/OHYcz8zi9BqPfCQ/e4poFiWuu3ReWPM5QBQ0jzye8M2PQiQ
imXiLOyyyhLkFIL5II+JxSwoXR2zNK5idx9IiKOiJpIrxD0ZTEde5vzNJbmFM4TObAyXx56ZKhjO
Ol5jePy08BDOFfssfLb0W+OyVUDb75qopFTQK5WPbLxvfG9RIWs1YQ49BHuGr4ejmJq3TFGkRtQ/
byTF0c81q7CUI8ZaCrkuYyK2lBJ7kbPnkj6yfkCoBBiEfu167JOMN0tOr/8bRqRk2M9c7BaCzMrU
ie1SBSTWlUARQ2HYUJ2v6GhUKYqFdhqt4lGGXofBwuQUM6Xo+nRdTr9uXMq2Fgcnde+K0L8Pm00E
n6IAtHHfgAN7CZ5IYefBN99j2ohlOfe3K5J9ze3EJasfnrJI0ypiu8GZYacbtkuupj4QI5eiNOtv
raN5lfSdWoc+BhAm7qK9PTdozWlFEDV/wi4gDnOZ05eORDd0S9YciGfhKtMzcRKAINekoLQODHF2
UMzDjv0MeY1fl3oRiHw9zwQKAfbz0trCgdRBld0/T3uZNIonsLSeLusrDSWCGE2K6BW+A/HBcmqL
iNJ8CQfEEnP5ioMBcOX6asgyjqaKnDjpwgLHOxgGfT22yjla/Xmal3dMbyUwsim/mAjjy/JzRdL3
yG7Hoco4VIsdZkCDBJY/y3Eid4Oqnx87RcZBDXLJ9sngLJLpErer0jNc4FXB0CSVrbuEKVc5i+i3
PfMbRt5ntHkBO/xqAutcZlm3G4iAokS9nL9m4Jzvags/0Bua5jxD/8/jfW2NjI1eqEZy9WztyjAO
vU1Xkp03SfiOM+Dk6Toos6u5B4iGVxGi0tucqbh5vZM0nzJA77zGB3jASKEJcp8X5evuSBBN802N
LKE7Dn3Vyp9p4sZIOpUUsErZeImN8Dnp/7Od/VMdM/5nBe7u935djPY6uiWNjxGTCSKsT3ofQ0kl
axJUZWEVS1SScq2HTXd0oV5Pw41r7/bZYpxK0GMkwCYBQLs/DsYQRhtqcME1AV1+k8230ADE/O4w
7zUrd+NoePanjsh62Gjd/hyjBSS82nvXISoRZt/vkh2/Q7CmCSvKJhMTfuvE8dWtXQ/tnIg3il0m
wmtn/ocAOkWEcF1VfloIrRKSo3U86xPI6kyvIMKzSISubgfqo3cS9xlka84Wubp0flZJBYZHEdD1
1rBQ7l6q9Y5pZNJb6EldpLF1FFbNwcCkh/4INuchibTymqHTXkiuP+4DayB9QeD0IyfO/6ckJtMt
z28/FV/853kGUUwxWDI3yxx7+LCSzWtzbfNDVwT+ZOkuMuh04ER3H7NwL3rTi/Zw87ilfS+l9x0F
rGRLnnX8dhfJwKsAk0ZxHwYqLt92fRZ/mRuM+3SsaegYL6zyEjQhdsylVpW58jP6fHTGBj0CwM+x
ktwfS4Q2QGxCVzr3lhYj0O0sNXkBqEcQzXUSFjliVk7wS/C4GhkfyBku4UOs6NIakF1LvsIsUdgg
iQ6Lr7jrqxf5/ktx6uZZc2tAujY3YtSF6iwFg64ZieRKK6NdqaTFzavNNibbNdhqkMvrkUbQjx0A
+4Y76zOPnJ3GiOnZvDKmqhE15Niqr/06l6/ehN4gwLS8HdjeUw1eYAQ0O8FzQDK6qIDKa8iviJd5
g/5xbSs/mV3BRi7R0ZWdmdm+Kp0o6oxG6A9uyAYHYM0cTlTBq2c/uwm5whtIVn7eUfW8VlW8vWC5
FMN5b8Adi3dZm9y2msihv0x2SKIHxXMmyFEuxnBb+OyvMx7J29OkCQyIzjm9jZw5XPQUeBGhzAHM
InQpEqkfKbkwyIM7Eowfcxp4kDaGt6BthlD3UFpr5bdxZHmYA1ISdUwwWBzHXH8mq5R5rdJ8fvNg
X7twZPRENvBjcwwPCdi2G4wI20rKsmibWBc3tHfOMYhtuHBkqZiA5awRb59XpZ0+PGJRjEQeo4iC
5dsZWg/Z/cqGLleWBmG41nugO3ufZDVdUwQduv0iyj1rOusf624L18mI4zUVEzwQ3D3cXDbYaFQL
WbjZwtD+eraWVQ9NaLj5zmrLr0F7ARdxJmF0poZGRYUQdANqan/QfE0rvKgFLCj8uB3/E07VUEVh
PHqBjVjIbNIKG1WIKGjhfbtdROoZFUpZnlY065t/+jgfZX8p5iT6k55ddlref5+CNR1KGFNuHKg7
DqlzjsSR4944e1pKnMM7sgQl6Q/g8zYf97YdG1TkullN/+FFGIela6zggPBfxWF0Grt2uXcdQKR1
o3Zkzr0MSf1Dea2Z6wKCueW2scssPAeKkzxvzhxV3iNTQPV6ltvq4nZpOOy6XXmv3kSUvmBBHKhS
t3ZUP2Ezn2NdoMqRO+0ru1XrmpZk3f1O6PKI5fDbJEN6Ecqo4u/bOvxGStembhvadEf4/8BqApeE
8ue9BgpuNpGSbfLn4UXtrzjvBA+1wHgetoVC43bUgahA2ZoySCDHmn6DA3VlxZpEQILzxYrjvbFa
RbwqjpTvrYGrb3sVCE6BGtYllvZ1osWwrY+21mrNRfoY9aPflsoj8IZiO7/CFFTPZePTWPUlo0xD
osYiAsrHdjGFVS+WiqYQ8CMDG225VLV/AUOLk8VUAqUmwB4/vZErnUogOVT+4eie+DPrIIvtDMwA
bmvbIt8vEbmD7UQcUZhXgm+2wKQG72XQQ/KP1jzZRf3OWpLQNageWSnh4qS2oNMKAYaS2qUQwor+
Yen1sNFzli574zvf+MjcScRwelYuhwS8+JueBpojbNG77Xh5YB6n54Jgtvq55vpm2Zj9XDAeFzxk
EhFz8T9sng+B8Uv4FCwX3s2B/Z5Yq3K6UyxwnnOXRYVknKD4nHUSp7BmvNRJB0KoSyCb+dc7w6B6
kP5gdV+5weba285MqLSYkqhJyXKCZfiD5i8bauJ/5Yz5VgCbhMcEDIPpQLYKtmO9LAQLn1Lb8xMf
rnujtgTlYmdkJ0xuEJKnfEQphac/afs+sh88XZj3zN4nuqrN4DSk+SvrjwbbKDLTUB1zBsy0zDzG
IzDXfINGHszNr7urDlNz375GTEY9KujzQy5ffWkWEMC1pCCPt1fTXy6+u1dcPxzQ12YsEAlhCN6j
etINbeXMLLg0yvfbQLQmLDBXip6/PRtDZx+Ct6iVQD0uvFgFMMTVMOTJDhiUpy97TguA0G75mxIz
zbxzQ2ZYpJcdgUWgoriKuuwy0StY0253BWtOO2IKAqaiuw6CoiVZZlnLkmzPCwUm+CPCuus22iCe
85TWbkbX1XiC/BKiPRGocjNyllBgbfHlQOskMc+gVgLTXtxohM+75voUk4FO7tuj7oCs55hY31ks
qj0JT1oyv+C2vRmQvwwRH5nmlArJSh27GZwF/z037LtjIKn58Lze8iM28xGrhVENCRq2jSCcYuan
83bP9BtLE0a34H2NgiZyMwQvwCcRvSXX7PSj3NTFO3WxfVIDyjITQamhcKQMeVKa3ATOw86UtSD0
hU8BRdgzesY57KtgpksKCWgLxbcIcihAwR9q8G68XjIQe1jtKBQejj+2gyCevFXtM9Vf5SDfylVg
eeaNp+JkiCjIFUT2cDYuGWXdbOv24ru+ihCetaY+KLI+wEQrMfJ51VZaDudtrr/6yMubTf0kU1ZU
NlSKZwKA5NLOC/vE69yHhrQhojVIDpXV3DyeDA9J+loGxQX8bD5rYmP06eY1t/5yPsNfOrFyxHHh
qLnWR7j7ll/J212X0fbna6M7M/IvPdx4zjq+bE63uTAsHW/nHk+mHTFzWwTHb2r7zmlnJgsbkIL5
eaZMemnt5DoHdOfbV+ptFF1Exg/2JN63WXcQJzYZpQzaF6zoWOnyNn8dxX+lmFrjddBTnb0TV+Y4
m2p0GyxJinIaU06bUkfFcsqcQiR/sh5lA9HDK40L60F/EENSpkMQG9QG20O5GnTBMmRxiU6Q4RmQ
PZZksPzB4DuciTD95O6uo9GjYPRyMYR7NexVvBwAiyDjDe8V7VahAj7zRJrNs+spejBaZXHp+dCf
h29gDHRzY6MUuG+/ADJTSg6niHOT9B1nJ36VkCEo2jeRdrDxdf2TyaITlaebUoRg9t80zgxiq/Q8
H29oP0c9ed5titzS98c07Z1Tyx7DyqYKt77F77G0POhFw40uLEVHIE4rZPKj4ckXwSg2ox0OyaM9
SucDTYWFuh8Gb0R7wkmmsh63Txe7o0rZX2WVgmMuVTxrlcg4LGptncg4HImYdDAXx4n8RUsbTng+
LHfpFsCE7vXETViDVfobbnlDYJ1XHoeuUS+L1Kmwne2/nDqi8B8uI5IY6JX6k5B2LyVfdyw7q/SM
bvTy9HYjLBf04Usdye+PBnwXa2qFCkhXmDHfO20b6xP2+EhpZwz4eUnFHXi9RigRgxwU1ieJa7H9
zwfUfTdvfdnWGrjMfAFwNN2hFLZOPp5AvcJkz0YqN+eqDgWzlrlIex4xy225Gw/o2smRSK/bEv6v
G+EhSFYD5G6Gvg2VyRXASkR+Zfrj5mVoLOqtIbTLz7k9uiJ8ci9Yy4aqz6t+wKfXtUSYnS2GgaS1
Ri4Qh5+x/pk+XM9Gvsh2MStSSWBzodfx6ZgxHVVSzdh9/y6eOuyy4pt/iFigvgIh/EAF0UFkxnpN
pRDQyLdfdZD24sfB08MX5j7cT9vkQ7gie3l/6JZ21uQFmcRErm8ceKdPBCxrTp5GiM9i0oyVySW5
F7c7KSMbc5jMfpa7Mh/pE6XceuTty7FbIh4ufaJM35D1GcKZyx0BeiemgMCkZYi0/scqapFdOGSb
KbY8XnzyOumzLnSkFYnODjzH7yXQuE48vjeVlI9CD0iF1IGolqd1e9fBzKSk6ZCmNZuUQf2W+PM4
5qWmsujIqzrnLHla0KViK2j1YvEnkQGuV4/GrFGatpsFiP/gP7BrYSU1+P6gzTksdvSOpEpOa9U5
1/CaG7Oh96DbPrVMQIIjXpJ4+pUKI04bQWrz5pTBii1+dr5yrNG7X8WGrwoH7TT6XavYLMF/YHo7
Eh5hrAR3h+FWkl7WOrzNVSgC8x4yyXQu0vlgr8MJhHn8/dc93QQf5D+Hlgq2WNPUmQ3twkJqN58S
/v5Ww9rCAssT3S/k+bX9Nlxgz/VZmv+eeE4252fHcojGsZ8Hs4R3nMR6MYfNDLstJWn+KVkwX55A
rJWMjyUIUqdJNuhFjCkV+7YfLhHsLBgZ5/Xy6+mqluQeJjkQ5YNdRbBBMVNLhRFqa4LbwlWLW7na
8rDbcvQX0oYHvD/bYqCZ3QULtjbwIuzbM0H4jRWV8NqVNFhqKPkvWG4pRek7L0uRmZk0iwTlNCw/
3wZyP3tVCIv+7JoqMAEGqeA6Z16Oj4pQz0ieue1+RoOWIPrqHvC9BmzazNN5zpRcfIrnATglptcE
AQzY+qvGMVCATHn300q/B8hJtjecSXmYY+8Ve9JEWfcPpciTr93nJcxub132tE15GyQKzsjbAYi/
Bjs4Ozm1GdNFyHFnMGhaM6QAAtrSUxU9xdIJEEzSRbiM3542LdrDh+GgKGKXxstplbyGawiKidHd
QtYssSPzfTip+q8f1mrL/nTaBEJc7ztn04vLhejoB3xEw5eJ8JLt3BlpnwH0B47A8Irhm01BtGTB
xqzahHMF74jV77cVwthNI1QEsZaYUcxhOiRnFauYN7H2KVg9NbnRWGDZ7Mk3ED/2WYA/ZZ0K1LLU
8sooL/GiI97ISri3Wh9g3b0vudCc/o0Pz0eL8u855DosKmIFhZpWYQzLb/jlE10ZP5k5jiT1BhWg
Zt0vG+Fstvi/Brizblg+exwWTITZRQQ7tF1EbO8HKEiyqzeijXuqgySJjvDYg+YlRoTD20UPFTd9
iHtVzFoQVg0dpvLOsnZAC0kVrSajyvvPjnQ+keXZB+zM6MAJhx19EJNWHWf3r5It3y39AcZncMw5
zX/DYiiCVqyKb05kxAlUEKaKa5TuD1+9KqdldWlXfwgEmKF6VL+0JW5HZFrv+Uj9CWvwMvjGatqA
a4ruyVVZDEiQEd/3jgX76U0LLOuqxaaS9g/oFSPwyavjdeEPbFv0RypCqCJX6rem8eGADCeEnWpk
uYtr1behoFaLUtYHS6mKU9oOKrncRaycTX9NNZS/i8FUNnmTlLMJh+i3R/DoCCo81BGI0OA27SCU
aCRroIiIMS7cXFG2EEPjY7kFfMQ+LzKA3YWj8RBZcjWjiPiR+HphzCj7tvPRy5hi8D3rs+hahApV
MWqGytXiG/IlDsqEFPHGgLnixm3LC4ibKvGSygTAMfm8XCM/Keqj2ev2xO6LPg05+x1rocoTLskm
KGz7Wx9m64VhBlydd3DBOl4uArpXCHFdaDvIV83T9OYUAlU3HTyOvAmyE2cs+twaH+/akSvqTj2K
54+Q5b87d7GN6zvQK3uvDRQO+BNEBXRxXiySeV+RbP87HGTRhYcqjYEEDjwVOBTGN3iwAINdXf/L
DlRDljqloxxk8s++2bdqZnB+ROSaTiHVh06InNgAOEVXOLOrDmu0qnmRlM809dTe86AbBSM+D1j4
LRWb0Ze3eQoBtJg9YPyq2nl7eG76MxWO03TQyqiq5AB4fpmm58h+kl/vvqYInl8dYmuD7dgIXsch
jYrIVll0R7wWNeFYSSV8JT/QWVDKsi0sUp0LJltDXRFLZtf6/Ova1WOxE1b9ZJjGWa1rN9rR++AE
GFeq0sdEGaC2tj6CXdEnQOvj1LZETRRsQqAhvegpFuK7Qp1B/9wcMK8+0MrxiEkMKklXuiUxSHoz
aEIuCLh3rkE5/poww0Y8wwNZbaAwB9IJsLrjkgszY/495GUsE3baQxWfwy6dd3JbpeR0OfaUQKcR
V5L8xczRt9qlfiHTqmrVSzlDLOsV6phzCVzYaN6cn0yMNT1+u5VGjSl2xU1tInR3h4b8o3BxFEyc
+aHrB1PEUp0l/SRh0F76zXqUUqj2Lo/LsWt0jodD2dB1qa0ugNdW/srcxmmMR8LQ+5XshwwC5uJy
T6YBfaH5KX3/jhz1gSSBfoOSaxFr4hkPmH3s4ltuh/Ahxgja+CDRzxwzEIIPMKuv2oHq866onITN
nzWq787l2zAXWR1ECwXgnHxX0po1fvl7DjxcO+e44PJ/UWkCI+rvaiL2/U09byYE3Jzulb+ov7Gu
m5jEphEZId9VYuUP0xxdF+gfrHrbmK73Fps4bmI0Ymqs3szfoPbZaqTAL8XGs8h3D6hoVxC4ETyg
0kcII0FPx7uldcJtNhoEAuLJSUovftqKmNr5ZpZNqEsyLTShkDaiY1uz3JrGsIyBxaYNdSuOkDSj
BGXOzM5qvEve2g/vPMxgQcYhMpeLJlyNZub2bAH6gW9nGffbyvvOg7/YuyLqp6FoyWq/rxPyhBrn
Aw0JiT/NaG1N6RgnqyhysyjJkP6VWP7NtJYBNfDnaZLdHUnOgV1fQNLs4DT3VRmzSOYKi6nUCUsq
DBa3ZUJ9VNRjOTKpWwiuDbKk0bvymSlpLaREIa3qTMTMzCdV69vFCyrCpEQIEhRR0MvbLOvPGsR/
Y5xeA+Yd2ZvgpRnkNsCrwlI8I2y5K7g05jcyGsV1B8EHe9a/6kCqeShVlCe6jA91pQ8AztW2YJxo
HKT6fooJb18UGJCv+sE0KaEh8XoGql4Z5cL+60XjszNVoS+Ogu0iEO4Ch5/su02lPr2glFNwl59d
YIdeqIlzVU1W6eK6olSQW67BrpNyXOONTXH7TGUnvtaq9KNtwIigHBhEPnyPZKBqTWwRccrsy6HG
llqBYEDn7yTxfVniwgBgaCstvVSKHhPp5bgiM9kU9PzBZuIDQjgxStMaAyKU9jeYImZBJGvY08Li
I9Q6Q+C3ZcifIws5R3o3moWVh9CN9iwJ05uDK7VEI9AZgyLk/m8B+bYm9SZPZ+n+y1OVXVjdlmTG
JGwTPk31eLOggFcsr68muH5B0i0DwDJVpsCVGERtlRFejj1tsNoewc5AuQKfZjxl9YTFi1g3F58L
SP65X9tSEPjBfeKMHVHXBf4DFXOkIAongVQRF2VW4njYj6Ti1nJfPh1J8UNoNYZp18lcn9vfMJxf
J7SbyUE/O88O8bhZ3S7zkFgTcS7Qc45VkhJvzCxDVg1iOSbaRqIz9nZHA6oPAXJXk2IjcgKLw8dd
tfouKVY32t/BQpR/oZfVGIJz7NS3Q6e7UghBLz6xj/QyVkwjHovUgjsD4Jwfx5/KYpiLhGcUdeOq
273YfuCZifwxAuPeCkF4GhVU+jtWb9uZYC3cpn8Ip1TrMq9C6Tc/2rARskgLJuPDGtQJpxRjpzmS
ntBxwAYRcZMtCzvQxGzKq2u1bXmfHr9qpnJ1CsBkn9l3s6hHSzR10zNX+cMFTHWco7Pr3r4fA3l5
cwFS9RYbYmxMf6ljTAY5pKq5VB2Jl7WGBHl0ZrtRWhEW6IQdAPkFgjQpMqHOy7zABbFVgiFu7jBB
ZDE1iv0wF8zDV5WapeILoKSR4v+SNAhvhLvnwANW/C6x/EwkeiVLDNE4l5RX4rihDP9dkY/mmjDu
c9uFIogl5MFINJetr1vhOkZiUFDolhyBjxkZPsPlm8GNHgBjDdakc3kJljP6GGiRbE4PKhO9xPSL
YmEgcS20v6CBWl4x4s6UACpJjxnuV3YJnYpgNtOyIQhl/NHk9DI+6cSTt4WYet+s1dhGL502cVhd
Dc3+Ihi1B5EZR//nqzIZfL1LsNAEMTDyP0l2M/gtAdTu7/1CsKMsjh3HOevNh8TbgBN9cN6MOpZH
F+hReS1S7gmUgKVvFMeOswbJ2JZkwgMhoPyOT5cnOAAn7qyqWKaF1HAlikRcFsnJ5ZrLXOmkEuT8
t4cfLPl26TXeSMfU4WELmy2PCH3NpFszRkaknxF5kw3h92sJXx56bEaPhZNMPrMXxzzjwUpd85S6
bTEj9erZlDVLLDXEMC6J9yws5xvaitNKp0unTpi4fsiJDTpe6C7lt7FdAlw15jfcf0mJ757i1z//
KS4M0IsHLNHgE5p7Rjp/mQxxukx/EVqnu+x9mYcouoRiCE7H5E3Q5LBudC5nQ3MmlELGlfKc7Hgc
rAfIt8/RrugIvqgnRp5d94GQwYbs+U92V11Htf5UjpSnsPVMNni9VcX84V4vKlCJYKORFdZDUZOX
Gxno+xG20Ofm9hlm/QDeDOxO0XTE2Tev/FfjC26/D064yXj6V86g7rPScB8GaQufUZh/Pmt6ZSRo
oKiLpDf2nVkkT+ZXMNnh1rStctfE0+JNsUaghB4wmgvey6JkXj+5r1aFOEDzYih3L2Za4t6qkmqL
nWhZFQAf+wsEeCRo++biIEOCJWX/8VCa1DlYBaF84DmN43fnUnBi7VMSUOcBaiRPRzPm89tI6mnZ
u1/kunV2UmCWeCxK7h/YenMlpSj+rIKEFb0o/hIzxhawgLLw2KdGXi61Vt8KpnkJ1TUe7QMgY78q
KXbn06Qocgpac+s90xslvTZFy7aTUBxvswEURq7P0R1UvcPhE5Fgx3NEX0AHP4gUQmrAn1bFEk+p
pfAkLxXBJUkrQiCpYY0EAevhp5f8RFNsgrRsLw+47RteKrG0CMf+d2KZV1fsQ/sqPtK/xCBHPh4I
C42454tXLsAjeiQfVvveDtJDxd44Yx739miO+yXWpm0rQGGP+WCgcwOizbj5LRUpV05uEAiprlX6
fqcs0OCiWAbF886hCJjkg5JYaMmW5D9QJ9V+L0R+zfGWCnqPLuXNyEquxe0ulttgJOcCk7JvKCSP
Kc4Wt/3/7JDca94tHDiFYrLZbYW8jkK9blIkqNXxDRFY4v1JW0d0KdX0N+lhy+OIdYXxbxyZPWwU
KntSHeGZ2kXIs/d6pJQOyK/WsJgzV7C25UJ+KdOpKdKMTBSsaaQfoWGsKD8ItazeQqSufmlZUB8D
u7o6rh6cfCu9RSVxTjxZv15qtoT0CuGBuQOvvX4YlR7dXdEaih349hoE2Gjpn18s7rwYR0MEjbOT
xAtM4gA0Kf8uNWfqJKELFusY4DP3zzFKpbl2XKWrLQfEHfuOUmHQ8bmf/SosBYySgDaBlb9Udp1z
CdBszCCVzI0aEa/aCaYHBDj/x5Np5yhHJXYDK1l7kWjVgzTvCQGBQq+bvVHNlWRdAAEF4WuOQyiM
+y+FD+zMaIMQxUDuLhil33EB3wOF1X9LAGHsqP2kXLsCa2LdBDwlKUTso+GY/pR6NDy5bQxIYq/n
EYnXFFJvwvvuTjiWIA0DGb0FjeRYr4Yiewpl7yuBCDcxWal5nFY5lcKu5UVNSR7VehZ88/2Npvko
sR9tGmVAA/NoTRldlwvkpVIx1eW3NgAreln2i8ELWvgQ7Q7lgOP0TEak/QayQ42DulNeM92nnSzv
VaVAPlwITPSeDvIk2xUKrZJzO3uispU/uIkNSOpuRSdCBRxDO+SjJsUA7bJl2pTSHVilZxjMrcHg
7KEPVGLcAgTGC+TspaEUM/1aqVm8BiP8YSVJ+gU4yxDvCXf3wGcmXO1vbCaCfwmIIDqeSXDCwd13
twAzNm4ayIGJoXdguDQAXUDWF0RNjycJp3am+DiPjbx3+5A7dsPv++aQYWnB8P+e+aSvBVOXEKyj
TXgPBgAXcxjm73qtaerbS1c+6X3gk45VW9GdTEjzYwhZue3FFegxgvAgahmPVLIutpu9WNRwDCmq
ttPbiQQgzn0MPdVzI06EtwF16Mwh9nqc3x0Y0ZxfKDlg8VDTonL1qAqhj1vR4wx3H5lWjm/z9ond
yeyTpewSujoUxdFQy0gpZVD+CxnhG7qZrcKemtRrqzbMumANMr8N+gHI1+LcschI0ZLDw5DHc8X7
Y/E8EuZd/dWU/BT3TB4uUbi7XrglY0LlE01jqwyArvPyqnZ7aNcGfzJ9F77+0bxLCq19mMsQVjAx
Eie0wgl14eWQYFlJ2L10DZoMN+k64Db6DLr250J9SmVKj0w14l+u3zH+6GgUS9uQ1+23CEuLfU+/
t+rzX88HAXhXxDhSGMFZenMetSqLsj3EULlIVc/8WmUFLd0s33MN6LXU25OY/8DGHqFQzCpGwuI7
Dfqn5SmdW396cilJp11RYDpTaaL6WtRhjJZYZuZw6pnMqNclgUHkDXNlxrhXNQleMqW+F4l6dlRz
ONUuwzq7HbDzG9/J1rSBN9VPUsvX8go7Z1oo0fYza4jvM8lLk5hNN5ugDt3cHBmHpshpZ8SwNfJa
Xy0IySmCbA4E8mI9A8PiIHH++54PUB7i64CK/8U2RDUpy/s6rvUlLh+WsYoiGv9uMgotjWSA6Kq4
yhPmkDjkv9caXGcKTKT9DM0WUNWzMv2J+t4zFNJGWPK7Yxmd4MowVNfCC+kXeySnuS5O4tIPved0
WiidFQZgtCYf4hjaEMWvOWXAuKcLmGC6mpoTkUDw/2FNuFUPeUfUehGBU0gWEA/d7uiGp86fTcp4
nqufALqvmr641t/hGs3kod/Ls4iLiJniVtRz8cVPUNfn3oUwn9GUhdURJJoKZfDy/u18nrP7yqMs
t9WCJv0O+7D4OujI82NzoaWPoQ22fqFAkFdAgq+yzqlKbDvPQyUwBrtCjssMxyX+cN7yneoaf+fB
7JTUf66TCq3JspI1NKoBYIKo0sNNacfTfaye2fuQqhFXzeaV96Lyu9Kh29AlYonThVcNPG1zT62Y
HU/G5OliLi/W0Ax9u7yf4YUNu/c9wOnRygZJa5ap/vIdCHkNdEg2B/rDX0f6ihZXu3xJjgWCAxkq
4ZmoqL6Ru6Uesral5rEj+io4xCCvaWYlIwE2C9nb3XAVjsPWz0e9Jr9nCxgAmtwOm+mB2yO/3WpA
4pdm4v1qKK3PWz5kTZ6aTR9t9yH0SpvukrIgS7pkAQuzPFW1YUX+hry3n6VRgLt41Ly0vYRhJNmI
VSnr/WEeKqyH5z/7gK+YF39jnC42/JoiYyxyh10tt+8+UdhbVKEZ+sJHDmn/DyxXQfCCHpnMpglP
FM8ZCEBKWUTOGGG7Eq5h+f+xIOtuEx8uLORHwy3wlaBaDu5ADqSmN7C0eijTuc5E0a8i2KDtiRnr
SDU+DrOe3umfoeWhP8pNr5PsPxcYSOSjfPjlF32q9hGbnnMSW7qrzogQm+FwUghcEEc3+h6L+qxz
9+eRlKEInwrRd3Vg6F7sLix/Jrm5YUr3M8myTZMFRcD9GgkwtKWzIGHeOusjPhHejLZR76Gd+/p+
Od5GBhLFMP/LoTjHRfizLLviZ9A5/irHrUjZnGfzNDqquVWVAtOr+wl1uwMYj/fKjyAh6+er69uY
vQe7PQN8zbL2VHx0wX5U6ejc5idmZUuaYOLN0NGLZ5fKsddxZlS9oFcXVr6vrBm5wC92aCvy3OpC
KUwgWEhw1sUYBhyYBHnGgUcuS0r++ysoxZe+BCnceR+NIrkV8hf/odFjjVu8CH5zdzU1tMyiK0tM
1/YDHeHIKjZ752kINhrgyx6WNetz8UhHlPxVkgqLbABqfFG6Ycvsyy52RA/L4aA2JB5WlV2V8tTR
R/yvQ9Ts1VGYdc0UvsnR0nfFul0Hwq4raLqKr4oWJiWWlHiqFQ1Kg7aUNGJLkxHhfI87lEVTfGK3
wdjTYPbaYuOD7HbYpIG2R+M8GlO8Y+SBenmyY6O2XJeIW0/xFI5OTonYptcZUmMhXP4BTrVAg1nv
6NxmrUSh9gSMZHdNPk6KU/qnDPUwAEUvxYbfiC5+qM3B+t8lL5gCKbd2Nif2BmN105i0l8m/mcib
1aMUJCIOakk/noUicmIWHzeCuDRnHdLOk0oDIjEwflULMv6JKkYcBWQuMovsfZRa3LCk4lliWCPF
6npFXafl4KmhvEhhxjZbYK0reRPParMxt1WAOiY11a3T8M7PQlY1tXR9SQJd85C6Yw/VVzf33lTb
onNfLa77tZB4rRKnLgPEL2IQkK+UI25fLW+k69AkmPW4Zk+s9OnoQzW0SYp4U235uLY+xWo6PRqq
PZe6AYtXHYUdKm1QATOrHFI3hRh2lmSK5qBwvC6dF8dy1V0n2Kk1XafC0Is+o1l9XB4KiUFY1Xpm
BvHuLQEfVy83sByZirqiEbpDkBWemgIOKABFSvf1EnHJfgaFcBkb9EF/CLddPacMrLWHGzqo9aS6
PXeieVb7dRnYQ2cLBrblTOFLK7QJa4Z97s1/SrEgJoloxgEZlbZsosoqkZPJLZo4tyDaqHKU+uTu
XlfRzbt3KO2JTO96nReqwd8/uTJi9lphrnh7h2InlUbwj7gf+Lg7t0CqhkuzGfCh1pDvqTzzCVgx
63OhGZ+SOA9wCyab/fceUbjm5vta7PHNWca3Ch87ZcIS/zewiL2R9+IjVDHChLrlxzi3ImXG9Lcb
gUIyq2J356hpMzPzjLlzbg0rfrNcmyWfrXRnNxxa0bnbaMaQILeCQoEDkzN/G9xTZAPQCi/k2k6+
/K+x2q4/T3IUb3pfN5CsH0dC27X0ZdPWrwGYk+nweMvBiZ3LikAuTofZA3KLcERNC35/tj7Yb0h1
ESzcinSCAhjNtaUzA/RUfRI+0kQMmQB4gyhzIV5ewphKFyBJ2Z+iPwJLYClNrDYpAYUer63B77j3
jDc7HNddU5tcxtmJJmNRniOGU2HpEohLLII8ZGRpEDfqOkCA/I0byVMFj1tIWsuHlGBswxSxt6aL
tPazcC7wud6kg5SBPwZiR/8DeMFZ49sk5ubNC7PPS+n+AhYax/rxMu6fGcf+rVwPBXZu6EJqrevR
MkLJgUeOt/yxd3PE/MPbUHRx5KhfiheW72LQhrIQ1ncZOC8KlUeGhyEjwIHaEXnA1HDIZmVJdsfB
0nhiO9Lg2aUvgzQK6r3wKMv1by4jJtUhhMuW5SIHLP/UnESmRxrkPc8x0qULCvNa0xxeqsW3oYJU
s7QVJDI9UA75IlcUSaBN25otRB22Nm049ePdUzPwl4CpvrOv7lbr8QcxawLdv54yNdOEDj1FNof0
SAXdfM1vyvwFKlG6tGMw0IOvmMnvalKtYaXWUyRJJkjlQCrrkThOx/jHRzWTeMVMPBijs4Q4hUbe
wrlR/i/a1g3SNuhtUAwmEg2ND0aNXNKwzKfUJovOE1CzUC9aDMjshptLlDxvM7OgFtbGteIyyKmm
IV8tsJ0JG/CzFfmuT0yzqr5fWbZh8GUGFi04wpjdHLfaagFWtMTG0Phj/LLAbGvtlr07pZ7DXKKr
4ypEHCcXgV3QLfZ5GxTqtxftLtopRAGtUG84+YCBttALJTFK8wKBrELt5tscxy4JqKjERtUUW3b4
f9gvQDtJ7xX5IpZs54KoWhDula1D6wDIB5tOx0UqBely6M2/CSeBSHJjcuB90lpGTo3fP7KD9YPR
OGP2lBC4mo2G8gLi9Z4dy36MWHwBqUPpwnXiQhIRtJ3927s/o6WGXvAyEV2d2m31n9gTVD0ITd8W
8dy4yWk45v1hkixwmRbjKsUwtWHVTFU7kwiM9Tvs/mJ1nM7OmoJ6jYU8jh/7YOCNMfq6FRHUiQSV
n4zW3RLYpbiGqW6SitzsqPuHXVBq8O21Vk1kGb7ibsNr3rrEE1KPD//gwTqGqweTfg2UbLwCIaow
TYeHsTv9ZYRUIZgqrlmSIAJO+ixFbaZVFe5nYRggBD7Aogmobs/64k/dwp+TXtTmi+IuE9ZxkNNs
Br2qp/33UPB0IhuFcgyA1Ka9WGwCl3o+9/qB7+s/dOk/4RV+oGsZY7kvu7uSShzfZkoyRIqBU8f4
xNKcyCiAyc6CepAtfPOxJWpUCUMQmOUv5Y7fgJazeYfk2humIu/AuhImmspjkRGmyPC4a/ByLrgd
GpNpOqKvfL1lX6hmFMO/S8bqlwPzy2WPs+niWC/e/Qfje/eg6VOiTnNQHCbBTOI4PKn3LVuZAPM5
15Y5un2pXnRVRrM5MPN6i6JY2KnRdILtIZEHN3NUcw10sqD81PyA7lGEGxtqpCB7q80et4nKNuPG
B9H1ERY5It9C6FrJNLDflgmYF1rE6GTidGG/7tWRBh0+TXjiHru35g7tYlxzrARijk4Woo12C8Y1
PCSJUjFtQy5Q7eP3mcl8HFoe+L+43ZoMwKwoqoRFThfnxp//tSgtFh6uARrQL8rwRn3qCLGA96sg
dkEjjq+jDRDRHnRtblBJEuTKKDBZ+9Wf2w09uUKUUq7wHXqbjKFM6WvgRc0TfsYH1Kq8NCYe0cx1
VRUgf9ZQxuD52ccX3Fd3uscahje0lSuQ/LcJUPEba7czlhtsD6P6BbZrazFOehC8FA6BEt36R84Q
B9RjqeHyW60/rN8UPY6Di+ot4vXzKYBpVNSFKtZfI7b1WIoESICMyFrqH8QXVlay5QdkZOCNT14I
iUeBIPwlme9cBOJDi6tuXTA7hWl6ZfJuaHMScUyJ4XtvPazUHyilumKJGVh0AF9jRhKjLR+Nuolq
AgYlT2WoZibqASLItCP/uOVz/11ZZgEZk3kkUOm1g5SG+sf4KAsBOU6MtCP08LhCsxXytRxawRPi
niUPPpp56K2nAqoE429dNgJkCxLsKZarZebt9Q5pDH3iiRoeSZYXLb6H4a5Qq8EseIpR30SABNCk
5kaF9pL3K7pdUwrMo0dSwREebMelSp9UBD7GDwdVUpTB0Bj8bZEMz35XhpSpfF4JIR3Vw09sj4RS
17GIbHCLii4dKFDcQCnhnH8gLXILUQj8yRQ3z9yiSpcqSUDFnYYVrw/EeOLtbeAa6vABQpc5xH3L
IaAYWu+HzY4DeZcD9JcLjQoE0EYwP39f19Z8fXk2lKjHi6gLvmkTRGgpVFQ6JqPrRjGEn8J7tfPi
sh4MFIgvXkbv150ky8tRLPUEH1ESQr/PkBFtbw7xxcivKd0cRGP5dMwX2OXqwty8Psf55VKvTkur
GTuyxWQKk7SuQfB1nci5crxdhPa447UE66S5TNrYen74uzfeMJikdnIIrrumKQcEDtvFMgZy6g1C
5IHljmYehtERF6QSy87Yy+S304v1TNq5ck77UTXunFRXEzMvyDJBFDPHFG+MteGT1tZRCr2f4316
Mkb3JLOt9JVDb+hXX01WNhkaBgS23wCXydWceV0MAdityZmLuqVM1qSGuK9+XmDCuSE5wkI87o5O
GlphaHXO9Dz3gCNh1B7cpoin/en4lfRPEQTgVS2ynunUfy1TcVzu+VdTNRjLolinnQUYeP8Bro89
QwR5yrEUkcx3hjjIU77Es+en1+aQNGsFZ67+FthEAT83OjYanmpC8IzVSGkXV3Lp7cwVZAOAzu4C
YXwqm+l0TebF67fP4+4T7Kpsn3c4ymt5kF1BlDQhOaVdGj+W8UgqIkEP4rlCcK4qW2kfPxFgdVsT
zl+EH7NeVTpQp18zBFv2f87dtb0O0smCNFUxIZv2qeY9EgFlzJ7tFjh1UfZVw2Z5s89FwE1NH7sR
ZIXyRciVmP7jgQ80k5bWGkVVqt+zlX510bmaC20fUchsXPH3yEHGGJCdTdD4ILFMCUfvNbr40Rqv
sfDRaPz2Rnd0aaJ1sbQ/c76v8dqg+LDWWJr1XD3j7sJh8orDnHSqu93HBuRUJ1IWeCQdxuLWl9j9
QGmMyBizI7jZvPi32l36CFeqh2lc5vNe0OIaXoLiv3+iEiNRdTLWlHxXaKmxYy56Co5HZQ9He1+A
PikS6UunOl5kbf31/cD0D7S1cu++le/ik/MZnk1QZSOjO7mG9xtq1c5OsmCGal7Rfo8h+DUYdD+R
HJqOlHnOObVBmpkrQjMa3lo1EIsIW1UT1OeCP1AY9+CEqigHpHqIHsbf/OWaE48Y7mnIzqOTR37D
G3n/uSxp4Uu+9zr0UDsQKgcl+Bn8XynWsdQFqHXtVbLId11CxEe3e63L1sVuad2Wjawq/ALm7ay1
rhxcpz/Sk+LytanqUsNIcctHZO53NifPHtJa+LSOzJZA8YwOvSQydFqa4OQfcoAQzas/7EB/9UH6
2D9uQNZKASTBNEpVt49tm/ANchtUbuUSGXt4QYA2XHjuo1iEDrfQPwaHRC55JsnGMkxTmiecdUq9
PSatWbmAQCQ1IsAmfzfs7IVGvh3a/QwqGqR/5PcrbUG9gXGNk/pP51e5Cie50AFglsNLQbUE7UR0
7TeF2/Ml8msUGv3vyOvcPpt5SbGHOnNgpZExkBZX5ylTqWfrYlxrCwPGcxfc+IcN4UdnWcDFxvBB
RCvvRDBea94dPWTiWr4FbvmhCKhU+FxIyl9xAmAlBznVmLJipuUUlAs6c89J8XxX5tyS7GSLWkHe
PbYXNhrSN+Tgddz08w26CXTNzcVm7Qlht9rXCji6+N1AhvUM5O010JW64Q7G3esAoZrkJSbSD3n2
Vmg403EeKacPSTiBTCxICxHXmlRLLneQxRZ6poQELVPftpLu0Rqd/FFwWTE0FfJX/NVFTYzS7LK7
9cJP+FNL5aqMoLaDGUkl0l6nw60yTKxdUHevQ5QI9nh+Ojx40v6EUIh44Qgu1sDXcYgc7w2CGwhG
PT2UFil+swyAXEfCZehC+xP5pY3vLjn7XR5C2WtijSZL0w6mIuJ5XeKZ40tJAQ8zByHkEr24Qauw
CWZcqtpsez9Tse1z2sS84HoQ8P1MP3Kob6VfEJkCnZ95yAk5zzElGr/RF+wu15rFg35q/yH/Bu3b
iKVisTGh5xUqJVMswYCjzGDUuOgevOtheFe1K0l/Ltk6JETpMSQQHddgWbEUROtUwu4EsngEVVkQ
Nbpn0Gi+11qiMu68TQnYU7xXe7rORrf/aeA/9sziofLOcfjaLiUvV3xnVCj6nUeHcYqx3Cnscf3c
LOHXsg1Q7hs/fCKt4oV6JTa+abTdoXfJ7X0338dUA+HVC9YvNcRVN4+IrA/8ThPNrh0WttSa+1q9
Ye0bPs2N53pmoStxgBSOAEyscQlh8yVqMKSSqhGOfX8lkTSbtwRpRuyNDWfLiZB5yTfwzksMx8NB
NJ8mp13d/uOagK5UzKF5JS8pPDBfLBW6gjK0tnJn47232GJSjSPwkTkJkRj8RwmHOZXTN4dPJ15J
T8zLZs254lD4zUGx5HAW2AiJHhbCacU5C0Fbh7p7X5cTlKmGdJ/7ugdA8h6+pVsbfQyxGjLVlYay
YMYDhwKBnUoTgV6U8gSq4m+gKO7Y+bwgk2dxProyjeApynFxi3GJjZKgW5LRgvUqDgS4lmkFZOt/
xAj1WThZ5ZCXz244MsgLwRnz400qzCuD7c+2mAkGKnW5m8CAz2Krkvz1jwjoVOk2xS5zwkCzPBIm
72KWYaPyg5AJYnYhkr2aX1JsRIkronqw3eOITWcwr+bKQHlXFRnBohcU6yNrMQvRmzsrvNgFKObs
Afxrcg140hV7ygr22YPC13aDEgDpp7pzP/lyVCT66otfEqiwMqfIl210yE9H8tmGvQhFq9NxRKUm
xAo7OpC/OfO8hD8GztVtnx4CIoENObgOPNsuHSBKkyk/MbvqfkbxNhQOs0VG7m7q7Yr32g+2qHtp
QDm0Pn2/HG+DXJP7VS9haSMDE2xwzZ//Eo5TapgzhYQseq5M5iG3U7iinnsROUo5ULppcv8Vfzwy
n+0MncRS46HZrfYav2o+QwlmvLapXGTnQwZvT/QOvFU7yHtMhYDxO4YVqsT1GAKfRWy0M1lW2x88
bxDRuFRxSjvHPggZJDGqNyQ9DNDLUhTy1YPcN4YVQaBbeu4nBGd4lWBlaRszRUmIwaU39iMF/nX9
OYqet72iPYvMZyzyFAgc/vb5CBjL/iOjBNikgD79CY2oCZd80cPMwGHsLWA/2e3VSF7UG8D6hsoI
sIyB609Mc4CeboXMgWVM4WQE2/k1nu9cAHwoRwcMsZsc9iL4DdmeFnEmWvxHbLzA1stssKjTHMML
WPBuhzT/CoWrGrBbN3BNDId6yHGPETiTqbPuTpc0OrF0nT47MG9zg3MogoT34UxV6qKPXy9QAUY+
Vxzt/HQNecANo55h5eW7VxRDjhrf5GC30w9W/AcAi6wyOowUPpqy+NGYBKyJ2qtnpfg0P1n/cGeh
g2PXZIMLSyCU3eXMUH/S+KbsOOqsDBU6y8SfS/pg/EfVLnyUOS/5X3LIqT3KtJIb1SqudxG7d150
2RE/yka6VZ0QMGI8eTgf77kR7isuHkUBe36bAHekWxq+pbhnRNVKKTDMp+ILCPdNYYxdCdPpHIWQ
G5HEzUYlojZWTzRhVTyGu9R9pc2HD7SDKp242Dy2mJkIE0fvnnM3Eqjv6YPuZQQD4CoEOgs/IOl4
AjTU0PCOt+al+0VgHuTGWX+jXeI2DNhKy+lWVP5rI9mPAvpBEtG0p6yuiGmXupMicOTjONaOb5+U
S09Yjzng+flrULNvAvoweQyWbm+JKM9its6O22Ho6aipbeBnzkMQ67E+5Q0M7JkhFY/hxej0a6oP
RIEZJo7SbnRqLlrbnDpq1/Jz7Ytaf+fLiFBRjmwE2JsYQTLGeaEVO1qJfIdg/TrB6ie0YSzdK+8O
avmhtLG9gvwP/tBQGPxrOB8OdgqkUOGvvyCpracvnxWIx5x/I1JeXylvJxOo/NCDE8G93AR7SOOp
7v7yM7QEEAO7WoFdYEj0HE7mnxLfhDptgahV3Q/64MIUk59zrsj6RvBbJlo/eSjUgzhxwvIKjj18
XfI9IFQSBHalIsKM5GMdbPPxEokZWF2EC0yuzADqt8phKxMbRrSTk2A0s9J9hspZgzGwZOovhy5X
KpKtYC3dy9SzWJIj3wL4L9+0XvxQNtvj2PQfxjErwi6t6NRm0hcdH7/OZRkq+D38kclItTB7YlRt
DT/7hhWpr+yHy9/bF3Sq2cEiFD2B/GuhLXMgnjCkpVTOVpNus6/iH75LmNimZmeapr3vy+NGkIGf
M7es1PaYgx2Aon3mLBsUzih+LssnrKBm68DXzfFtO3FTGvTHZVRfiVawY8lZaZl/pzy5AgNQ+YGa
0esazOeGkf2lyD+pWt2oyB9ZHiQ6TQKva/dVhBEpLE7CI1pC5ZtjmT4qeHtlf1KQNHxJ9QVVqnXR
OXMYsoLPfY7NwPyWKWCcQx0YrRC65OK6NYoIZ/tL0LclRkASo3csc6CD2GV5dPf8q20OrogOLfkx
G9CVQbGdSHA9DyMSBVX8WhmdVoWw8CPaEyIlWRMdbw00h3hFn9nk/jFNkqgsZ/xqWfvbYmwH7OiA
aP1teVt+UBUTntxAHeTEvksn/GuSxcBu1BTV5qrgFasY0nPtQgLLgDqRbckafHiFsPlB++97A1pO
GC+vlc701CEov6yjxk1R6RWOGMgsSQGLhQn5jYsDuSCuyAKliXuaW4aIvsiWyyPlb3Oj3UdaTExs
yBzxVCcFE1ONhnH7JsVX0soMq260BH9AcGW6MEa7syztvNoiFlNE6PnHlMbey52GwgMNK8SSxKQY
eA8oqZtn9FZTxMEpr9ZMKC90QIub6/1F+TchzwPymGtNlSirV65C2dJxxso2g+r/gIIL2gzPo1yu
+0iOvnaqhsrhRbF8Fb2UDga0jZ3Der2zdP8GNC4pauo/o0cw17nFibxDg+gonkM48TKk2W9//Tzm
sgULvPp2zFV1ejxrXgDfE8MvRa6jbjGooM0p5ZTVwNAW6Amr8LS+z0m8IUQ3zVWjTfgjG7SoC+9m
0dUwZu6ojmw2kkb+743CQ2X0IfBaM9mhXZ5PRLRr1SWNkav7ld6KbyDHemt0WvlTTIH9ELXnPcZN
w6p9eAIo+Jsb1YPeinjbmq1eKYlMdDXFNKjpGlU+/MQe+0Dx7m8nQERlGcZtWs2VjT1pSVy250Yd
oNSHTdjAaF60U+pwa/ttgce04dOuUo+7OpRzYQ5wPkPEGCxZ+R1zUBzxSyanXh/iofmw7DkJl7iS
sHRXQYSqLlNVvGroWcXdZE7/whyVpg+2ebUeIEv/8YTGXhxKPql1A9Cfu9YncFRGCNDYhTz+NzZx
b4uKZZAl1K+3cAh0lW6AoefOG0XoUnZaE5cAtCHrp+oLglUdoxxWuQxrLsy99GHabbN92h9qidSD
s43neDlKd9EyKEYsuFAD+pcbpAsq/Cfl+WbIiCInrEK1X6Gx4rEby/ogPcuVU3Bqjn/XLjBfZdtv
4z0hfxI4IMZAX3yKTpdf6KPphYIp7zpJr0klF80v6juZvJkgTeMupb8wJ0cWM0Jiwu7Kl8nI9/M3
JmzHk79YiQeW+V4kemTqs0/t6+fJUcJxZdTPiDXi4clR7K1nPQxrd+TvOPffZkzg5UOShXS8WfI6
abTISjPHTSW8FnvROh8mRHhv+lZGR4p4+/OCH6U7IdSzqWig2ftyXXdSkBrRoeUEJaB788Qnz3H5
CLd9emj0Sz+mDeQJ6PSDO1748EKun2flNHt+9QD1jioYQGO4LDU+g9+UsCti5ECovtSHAaVTZDnG
xEC6DlIRJFnKozGcjMrEo+UL53IU5oX6d+uVRCZMRZcSVRsxToXoHOJjIQcmXtzMM861Mo72or95
n2x7CWT+TXJsUhfIUMgnsYcPQVwZRQivVtmb7BJUJvlqTOAHxBUTjoN1kWIfYqKdeK4KPhvMlHFB
vgvC4ytaTNBQwVRcHgJ05oUYd7YShg+Ib4T47ZKkJJyz3k+WA1OQHvJwiw17J14Qvs5rJVaeXpRC
NhACTKQwpg9Lr+AzJZC+Btg4dLfPLSfMiYLjwHTNjBWZakAJRh3g+5AEMOA66jAIeh7oufvI93/u
2MTVV7h1SuecWzeQPqpbQuje2PUCuq8EYnwgHgAVLg7A44WpjD2jWKnibeac0x0iUfrqClVmUVgE
KZjdhwEluk2opN2B/9HIlxNXEnnf6/nDm6LWdwzHy1DR5FaoKfIc4jHXjS89/tKuBXFphANwNN+R
ist1FSvOz/ekb0L/N5KaHMTgLU5wfgoOPwNTMNUiLI+1+Ny5szGh8ogdARk6rWOlfCMdSPG6EQr8
/El0S3h8FDbt9q+6+IzSHG7Ao8Bg/uXmkBh0dnWdBMwS0ta1m9jTwxJGiQ8xhZqDns+bkQcbkGEN
JocAMSlmQg96WYAXk3RKEZZPiv/9kJomYJFHnUbiOTWZajUJjPpUvLI5gRTLFf7dRHj4ey1mio7F
QBu/NdwSE/q0GOv8550NMUzjnPXGIYSqgT7RM+lh62E+mppU3YnRe/b5pqc+4vcEspnPgZFuwYvn
qmII1RHGPIW6DwngzjsG/MJqlCdcV9qWd9wskbZcrDIU/rPAT+kMcwrFKXa7R2HrRNK12YMvuCoA
3Vby78S60iOhZCQwUO6z1+MTYVlCtrjWVWmDQS3OcJIfP+l9FdsenTvcJ8Wiy6JSD1Jv0PNeJ3nP
J0SkAlpUUL/fyEh0cT/jXRdYZg9Nu2nsYlQS6MQXK1uplCnJpvRplufGu40eqphQyBS2lmbI05g1
spABjoExdeo02MRsimyF5UKViq7mKQLgZGRwIyn3R+Zf5FD2rmcpxQVtWYs4rEetE+LvHvdGo9in
9liqcm0z3z1FjTdVBhX117EwQqmj2W8aFv0un/0hkHREWRh1L0fKExVigkA5AeMOkUlmnm2FoXpC
2j0QJgzjTm6H4HiNxjvi13/lpKm3Tttf27DJgXeeedhzjrYSOMLxF6gWKNR30Gslt+mlpMYNhPiw
21PwgQGElePaeVnYy3Mey5LftL7HLnUNJOb6BZXluLjz4yKUtufs0hgNcsqPIjBeArHu5NrmuL1v
qPFBdftOKIWZ8C9Ka0vkC4HvRR+7njNu6ovODrijopwOBoO3dImXK2pWGuTRVipydOSfI0ETzZry
snIKezmNzClqy338/vxcZa5uzDn8Ilt0/185LJf+2FH4qQCBXAd/QSaC16gVGvIYXGX5wOx/Wy+g
XNTYJ8PrmHYxPq9pEgX8e3cvEXYPV+kOO8HVM/A5Mb6KJIoG7qtyN8efzHT2tUQAMBpQdwmcuG2e
7k4dao2ghjGosrQ8Qfx93G2NeocRtE9NMJvYTY7KGYRX6KMI4pDUFE2Yu05Tr/GtLKBaO9uX9H1u
/Ae0kMHQEfOeYy9fmEHR6Mgvd4iY2lQYOf3g2YVIEU+g8tXxJ03oTlJ7nGJpnMgZR+VWm0j8/CO4
60YdvIcezJBv3/2JGj/MdkxfbOA6pzpKYh41zLI7O7bcoXr3byNS9Ev0eh30jUGozDwRAuxN5nWe
b/W83K2GyTdI8Q4Xy2g+XQrriyPUGgjG0P0P7tBe20yiMWaq8RhuVtqn+oK+jG2jFL/iGugPJDwV
DiSUz6eTKUHjBMxzxADnKiuKdiKStVpFhN2CsPlghIx86Gz27U9cje2mpJwKqEsYCjehFtkDuQkC
LxVcSbCleZJgG6LJRxbajOf56+6kjQpMN3ogl6L6QxFqMtSVOqOK3ayD8jPOoB3vfVvYtbvso6/W
T0Dju68//1sf7Z+yNS6lyB0GzIoQcCKQZYpj/Cjvw+yoP71u3SThsDtufN1qDByguZ8dVDHzVRrd
UjtU6WQA9fIuVA7tqLBpfz4SR4RjpZaTweR6HzcY+gIzHCGEOuYUXlUPG/nCH7I0nKouZ7RIRbcJ
jMO/gbymU45Qa/0N67pRUocwnRPYWOcbqI+jlfWFXDt6N9WR2Xff8s6AnzRoXN74mrZuQEdqS/bS
6VRKenRb+ZAso1ajtgWDh4f4gfJ3lsoX8ko5nBe3BU09aKEBBfk+Aru1CM4+Z8MNHCMMJEY4RoCi
cQZM2Xox9fEvXmfjXEMu+t2mCFW3KOyljrP42e/+M4Eqxaw4JnnAPKnFOQfHQaGeLTo3OG3Q5zUR
DpvthHjT9Gk1qfpIwGLclH0pHuj5XJkhg4fO80aQF7wINCmCuw+FQaXHYbYyQcVv5xjIXmVw6s5N
Z6GtvDTpX5OEEaln6/RJ1V/q7AYXvs9wniflPFSnSnZ/RwGs4Zsm8IqOBRdXfTBMxTw4IusegPJZ
5++LjiFXLS7Er/7I8lGSo4ZAYYA9EUVd2ttsNQpyPoSJgkk2tHBSKYReJqixJ+R3/mm+PHAO49Vw
KZys1/T6eKMvHqv36EEQpVd6kG+aQLIqEWerdxkqon9XJm27wwblegx2pdrnOwCLMVk9UKX9yNye
K3n3nP+GFM4Q6Q92XJlvz6gQ+KWhmT1LIStj/0Zeapqrf7LoHwDInTr3O78us2VhRTVzAt/0Ifw3
UOFZuN8710WTC5mrcydKSHt0kR0XYTrNalsOLfY4fZWaK85p7ofVwHb5l6vPyWirBs0vLZWbjyQU
FmThqAAmdvJHGGAyghKWR2eQFP82KbZhd6nM2vkQVRvdvV91K825wo5KN0f6ElQI1/t1PPFSSWwg
Tv9Xyy785FukHFabk+GviqLU0JizrpTfxghOQYUdVX4ZbdumY+0q8usaQzaGz7svtfEFT69qyZLg
s8K36dmm6fWM4uPn7CO5BM7MtdJ5kgKJAnWzjpAw5c/EpGpP6gHcKKce7pUpkCZqJXOYLMx6vIbc
x/Cfoq8Z9OsDnaOubf3peEtxUAAG/mNysdsVk2FdWwf7eeBGEJmbYefIz2jgsNluaYEdGPD4OMYx
umhS8Y0+YEuZeX7Od9TfWLp9L9XNXnF5p1+98S/0j7EV7/egfb6FFk2mRfHZHWkSpRcA/1Bxkmgy
/N3jdmRZGZUgaIx9M8e6vIxaLmNwtcZBUpmpQYKyt/zXM8cUUm8/9YFeMk0DNSqOcrtsPL3wr2bU
kyj8kZw5Vm0v5ET/Uk6V3/NoNz0t2O1v1U2ySMUoZZPWr7v6PYvs9r68rxjvy2FeXsEGebAJhZo4
Q8N8u6+qJbftoyk5v7MDu1et5BlTPid+unV+ZdAPkZnDy66GwFoXYH6TFx6pqoUP80lAdg50lRmD
t9avMy8wzEEJ9vrPAhXxvIRuEvcrw4wg1Cp0Py+JWpt4FxMr2bPiACZM+vGXPiHjdvjo1HqCmwBE
L7l8zkKIdiOVvObWDTQzvxlDDNDSKS9ZGZXGPWBcU+lhQoq9/DOyVabRv1iyeYWI4wz3NqzjkUj2
p2BiUEtzKtaD17hjfrYNGMt+0v86MmPWiTGpg0et+NYTQiKgDiCXXpC8VL6b4+lK1oL8PF+PmOZT
VhzbYwx54VTCdzJauQE/VOGhwzX2/3gVDB6rctjdXXaL9jWybO7eYCVpWyUlahRUzF3wUVbvg0Xd
RNE7h6HVezDsu3F34gn+Oq4AfeUJmcmDnQ7zKzlkxv3oL2vEIwQ+/cBYPONfiOVsItf+zljTAYuV
lPn3OgNQKyU2fiYEH0bjfcs5aR2lxqRV5zwWuvQ1MrwOfIrC0Jpf+sK8oM4QuJCItnzYRxGa1H34
Y9XDwvLINP3XTkSmC1w3Wa1eJ/yGIgoqXQpvroolFpyDZMDvLxT0Q9fvCSwf/h62XvQ1d43TWQFi
D3N9co2j6fChisHdVwlHAnTtbjtf/+JN0p40sfAnUzJKP3xpSHMmMogdT+0aAoTje6EsAy/pmOtE
TeRprh7Lway0q/NgsS/I1Y/GerKxecKYFlDBgRcWqbTKP8ezktSqsQbowYTSBUL+cmey0Zzzll6k
qS9rf593/ZeP5BZ+7tWUi/MIIDaPMJf4Db1OCv2fyRS8SNU+XTrEKOR0KGDbL2SFOSEJAgN4CFIo
0KK89CScDDgY9viOwXcwEZtuJz8exR3HoCddw53AEI7IQHX64l5njouHgMYaDXS8z8OOFJLNbLuK
0TRqEDCzZy2hYNet3XQnJyo7BwHufGlFRJSSdFjNotKwdkZm8cvFPB4LdSvid+NytSWHV5QBUiaj
45dKXSaY9d6WUBVybrv50wOcloMpPyrdZvCjHTJkS5kh86bW3f7d5/Sccm+taosSzYPhf5H7l2tX
7KM35Yem4Faaab8vMyAxJVayr2VZafQBqEPzGuDdwgQwlZSGNT9fFtp5DJWPO+yB2wNbHn7H3fj0
SARLaPi3uXlXq0LWDpT9AB3AS0i2UgC8i+XqSr/1KljL68qUI3wdoeBuMewVR0lYbWUjbApmr7ox
JEmGjHK/qij6oX+ePzQm1aMPikLmkWCxeoPiXoNHapCHfhfk3yYKqxUEl1ZkS1jDZenloN/CHoSs
yJLW4wkOwD1U8FlrSVFACSZipqr8O6bLSo2Ms1oARGzMeqNvdAwOz+paQnsxO6fFyDeI6EVSGjfl
33WmByeLTy7I0Y1U+++YkRhCdp44jgTOF3m8TYUmG76ow+Iwq/Nte6Qobb8mIj53jCEDpQqa3KOv
ueTUa5CB6iD4Au5daJR2OfzVxVuVOoYg4xqNSXQjpItMrKYPJwTL+YuMUaMO8f5lgGdGCf8rInl7
zBMUKvcTCrQb8pSdbKQYXY5UEwDBdNCj4mHtpAKZ2c+Jkt+a47jDVA3ROpvNvMdsNvfyRhATr7U7
95xcEslWdwAyCZHKI7AuHcxFAGcx8CfqrNhztvdtjNLOflyHX0hg+0T2nooe5FrICQmEkZb4vIlC
jvp41lNOwtjHqiISoy50qIsgICsFHPczd2SU2HM9FOLp5vsxCE+9ZEXs4tJaO9i8noiKOm8dFXc8
MsFrjx2sX0h6bBapSqQjlBcCUI1/sIWNamDRXElshwfU6F7x5if6UH9V46uBh3JDN2wg2S9un2+9
O3hddC/BMGyy9dhF9+176wIirc49yaHvQGOiTCv+vGgQIjsr4Q29KPZQeTMdNQBZv3HspHj4Nd7G
lp4ryPI/Dz1gHeDdyGWCJDcGIGN1CEVBzs0Q0YRWGXClFhVWoS98ZPl7W6sfRuePgZh0p0+OXxzJ
6OI6vPyaWjNQ2a+tF426/SBpTLJjUKZXMfJ3SKutT9TJUM7jI9OMR220xnEAQfGYgf+zLdntcZf9
QHpo6o/dUneC4uYzZaV6zeDv24XQaAXRJCcoBnVkSa2FmcHYW+r1q1gMajJijcI+NAb9C12PgVph
3aX7zQJ6wAgeMZrKhDTkjT/WyDxDq/Oe4j3G0CsHwO6KL7DVczkTtDsGHLn7WiDGiw2GR4LhHXp+
uaynX0MoaPnIYbxfBlfHB2MQpLtOM/o1CAUgIW9OtBET9exwLgc8POM+21Q4mzFPi602FkvMeuCg
yANG0SryW9dmOj3KO+tuiDVDDhp2BX7fhLr4ovREX5xpJGJoZBF3XYcvIC816MhWtwY0xQ5cw2hp
y8K1Z5uWXGkOYMEebhkg5N3Tfg3TkmHAs/AXyyeVUG5Jp9PWyVa+rMfoE+/JqAcF7sA6qLfB1gfc
y2HkB4FiiqA8cqet0/NsvlG55ugBh6Py7GTwP/yWmMpi/Y/UvSz+FqyvaFCa4AF7/QdbHwfM35US
LXcS5Ho4Cq0cQzVXR5vDz8cIeBzL75UfrNdmUTSIAQws7XrGRmnzOBS3pRrGLoaJTNyeavUEVYbl
9E8GjQbY5Oomg22rirRIqb3qR6dU7wAWRDERS6CWIpVaPms05sVZ9o2Bph+OHz3jmvVDvrsf3HOU
WrBnNYU4D4KtdJM3s4ry0uF6gwTC197YnW0XH+S1vvnRjB/EXI2KcEey6+wbMd9NymzHBYcnis/l
4gIS+gQICKINXyBV/48YsRPzRaAs9+Cw8+qXtJNzpeQon/zT33qB91sROjh92CqtwI3faqJZQFvz
UH/6jCmzaY1jciffi388tDYvr5jeOtdJ1X1u64UjVRID5utSP+SFmL2hxomO7QyqkUHojUoD+a6Y
C6uv2NF549xRzmLIbvdZJklaV+UTxos3WLBN4d2LEXbrMcMI1jtEhFp1HwNyP2AzQPsPHYbhSNzh
rWZfSC4uqfSBEOsL3JF8YUhAs+s/KUq2fGerxOozcywUEda2zyJOF9ejLxs1e1mclB3dQsCm8qTQ
8bJM8aJCZZbbyf8pC9xKTKwrOaESz2OxZ83c/93ChQ4ufnEKqqtstMQUtLKoh87p5B1NZ1sN2MVs
IzpjkehvgVBf6yiZ0C6wG8ZB6psJajjNtkyjYVlcgjViukDZ8pUoZeNiXtIXaHEAA7PiSbszN9Y8
15WOc5j/6kbKhWA9mDVJ2GWrbA/jSxXrG5kYNndgS9U2Qfz7e5CaORWLYDKwHKyok3e78ouBBsIR
a/73koUK7wP2Qmg+LZE/kSbYH3C4kwx0IteIzKuoetzE4k/7fZMrcGq8S6AKiIH8NZXXeM0GQiky
Nahk+EbpfJzLUqwLPLlopH28VEnq2RbsRdXgKHGppDvFCFLXl+XjglbDw86SCSPWHmTfBXd7hHYO
6DChdD9J/bZ21AlaQlIIwMvEEDj8nHQ+uOnF8tR/Z9qx+ngeuNulTIxP04Og0yrIKEay+/jKu5Sz
zaLoBxMPKg1LRr1y6tJdTMIKW+Z2Llmh5f6LmCST6SOYg77G2ghAr6kceA9FUSY+LrrMaEh8Efb9
wtH2/RujVIN67Rs0nLtzUL7ZQcXvkDWg3OinNytVS1hY33aevpTzi6lr/y+jbJdcMT3BJ2lW3KG0
sGpA/lzlXXc4FFLY9NIX7H8QJ7rgCvBiIBPbBr3d6bOlzpRRMLigAqyQh5mk1u+axulXZCZ0BFUx
zb+hHDDEfX/OHYKkC2Yayi0i8GJWMMbOtC1RQTxgUVQUwWTLBj3aYzSPaE4cSGcQORxwDe3AG5Il
g1Qm+SO3SybEBWwYqzwVLLmGEqLpf/dtvoEEqJLtlLUEbfV6ZP67wRa9cT/I4FwTh0PDyTN9Eyi9
CU7j3liECu193i6Hn7xilFqDtUMYDYbJ8XGDN2L54xhSsw/fj0fXUr3mQQ0pOAijm/fBVcFD5uxX
c0iPPiOOQ2oM9dvFDNwaRwePxLq+IU2WwTayCs7eLnd1sjbtyrXhL4ix6EE8Gh5qjbkLsqLIM6lp
ek0iOGx9qG0icJ2gbHecKphIxon0rWp5oVme/oHM0VwShCdzskYXo547vd4YPQGGdgZhFV1jt9c6
mwlY3YLfyEZsYy2Mpe5yJbieDcS8phJsFchkq8QWS+jir4As5Xp9YEYxbV7izekvwUsgssh2GEMg
aADL7SsX9hjon+D3LBQrNRHJRez/l7yL5TiMni0nOo75Kk5Jv/v9fSNbA5sN8YsFW66B1lZQeVq0
jluqmOpHgj9x+D1GktpOHFNPX3YN8hPbban9pzQBF2+wqiKSbk5lQ2eATcPMoE4T7s1t9qy0smqn
izg3Cd6SZTqsxCGuUGOcIKZd+XSZZfq1BcTxVs9hJY9gOo8Ye+1CW1WLt9nE6vqcU875LenL6Hzi
Sm+Xjl35sNrclhOyO9N/I6vpYYyxw4VJlN+pa+JgSYiHGUf6QphsoVXmG6XAWeOe1fQgAJwzNEq7
Fj36K+B7EJsHJk62AJuxq5cvn7h0zLf3lSGjNDi5lAoPIsPM1wksOr0g3Mx01H9HEtwreFS8qV0k
eqwGMwNARjY7jWW76aFROKag40Gc/V4JeH4KTblDeU8PgB35VRKyZAy5l9FTI3oe8mIUD7ip/bpC
YrKORXzBOVl6lBB1Ww5Y5DKu92ZE9gMuIUqFNHiU5b4jCkvFTvkhrbaprsJcMXE5rek26GzA8oCi
LVHKAuJJyFndNVaD60yjseycfeusu23KT6V0nWoK+QCaDF2FhwY8DdcVfBPPcrJ+qRoVr9gHTfKm
LTd6FtJd7oq81LEPrITCxEvqEFb+On9FpCDzT56TF7rb+uo92sQYFkVh7/WWYj++KWmYbNFeZdK9
ePFDuGuy6qgajDRXtGTTizgBbr8jV+5VNQVsdxzcMC8jRprauKp3y8wt1L95Z0w69wdtDr8ffjEg
MStSnFokrOD+hUJF2uriL4V3hZQDJYqoGxHQcAm3A2WTOHWNTi5f/rSX/pIFB3ZNMwzHiwd1fseX
tQxB1eEaz1ASbCFnJUvPsM4IhgAOd1JWXKCn5MxdQC7CL4E088+tWyEWsU2DInhMewLAcVA7YN9h
9H2n84EuT4kgW6jBaAOEGRA1CKIl5a/EH1Fxt8XXilVAV6dCDesyvKQb9NbOgPQQ4VV4oP/ZiXvD
gyjiEJegQFEnb9IdPRidzPy4R6ACFYZvyOOT6WC92rYDZZE/hrazqGj0OSIyQEqdOItsFwxWkaXH
QMcsjuHfakBSPrxrInwdNOvfUkJVxPnhZMJ/sc6ds3hkIYRl/XS9QN1TnDt8DaNLZvJXExfqC0hn
JPGePG+ylbhkZ+/u9EfH4igQCQkR+gpmTa/rOmCUyMuhPkR3f3eAl+zEyNc6ZqqjtJHeCIdmCw9l
DJrg9zsmzQnFk4bjlZElzbTFZcpjcsewFPF/QaxbHdp9Imj2G07GO984uewMMiUe+1VuwH+Pn59U
EcZMZvNCrKvTMsZIIUtq5u8Wq2V++FrRGIb0o52NlvcwwDwPj2kp+GMaa0kNSLGy+WnxeI8CGbS6
FL6n6c4eAdyXio6PGPo4C67802BSc2rXqN/Dq4jU9W8hS15J2uo5zG3f9ygCzEAA61Wa1Aeo6REo
xocrhuIUB+j38HMbeP7RIhin5dioqPPVMLLqQ+e9l+pYjBLX75lHefyQ8cbrOTy8/uGvGN4gfHER
us+vbIKiFDWIMiIA6X+EFvgvMxqQJoD0Qz7Km/NMMINzXN0RqPw6KZsJjUI6ddg6qtvfqLxHUAVn
MAiPRW5We1kdr7oCRfWLprm8WWF2pQOGCPWtVY44Tv33EGA8/7pNva9g1nPINFzXMo+ek4nETNCf
No1irkj0m108IkjM0alAgLlbO9HbkVXp/TDX8KNECr8O552rqiPnPM9TgYAeN6P7UYGsrCILJEEu
cHg4wfeWEEi+PLCrdqMjCuHPCUAK5Uxx00PGdmlAk1V6WUMUI7r0+PTjZhqky0MXH2oVPBJaD8MH
7Ds5FwT3b9OHAVLZJAh5yYyEoU7JMcnExhQ62ROlrX2LWdn7KR/hT/fZJFha7s/9qxyN55PpgOXm
c6EnHWelirMN3spTHzDeXvTYeBhpOn7guhVbRfxM/SirBVRnQtZ8vDCRQ8sRFVCmvzyeNNVsfJk1
GFLerIaPHUjeImK6fJwzLfmwJ96hKwXZnQMmD8mNRghAn3Xvo6MB3vnzipwtlK/tjtmT+geEmP6A
hJ2ECT+P4aB2nGrlftUtuatdVhpEqHjMBGXjGw+FJN4dehcEu2HOHPfXWNeFREv+yNhOpSm2A9wF
Ife3gIce1bot2khp9snBrsYWN+FG6ZPMtxTjfBADij5k2Tkk12ogLskhFgLGBPwRXdAl/AfoRjF6
ACkyj1jPuoJTrFxx/molkz4/F5v7JN1yt+YY+/O9iimVleZR8bQdahaEcmT8X7heGY3+44vIUJHp
Y/od0/JXo9WUaVQVNf26q+suljGnx3aaO5/f8bzMGYlpCWtSNNGPx5c4sBBUfLschZfSvwup0Xsi
Q9ir/DL7x0qSD2X2P0S4K6N45ydoxaKakckuZz1zOPP77bAML8yVEemVGNjvC5xSLguAO1jgM5Zw
G/e+lL1eYaM5IUbdLzCsET99ebp5BDt91jMVlnAcUjIB2Er2lCQP3+cpd3fPSnxLWNsmZ2rodTeW
ULgdoRtbSY/kfyM61ohFmX3PYmZPCY9hpJirQF7yYvMD1ZJRVDIOocW5Wg/LZ1ksoLaXzLQ2xDd1
21ErHkM1iaAOEFOGtAcENPlVe2CdPUZ/JT6tZCV2NEnahQeoGW2sUJg1Xe6W3k4ftdUI2mB8tjdG
c/tBhjmnYRpxj5vvAXvSw0iVOqgqi/C9J1HBAhk7aLGihQG5rzjtisX5xAU9+E/iP70fUrLpzO92
ApKNFiLyfyrhN/HLSeGQ55JrpL7zMT72lxS6+bRrTjw7R+jEnQEs/XKqVBvDoX2Fn148FJpv71wU
a7+S+esLuaVXtQ2u23dheODrbinAQU/ppbNU8LDiURFoDqpxEe0pXbYiXrOX9nL7DSaXQJXes/yu
hE9khWV+j1RRidNqAuFIxwam3saF+hIn/FOYnmUCujN7Wl+eW78sod/Ngo7OZImB4SjcLhamHAio
tMu5rAR/PyfgZzyy7YvUOe6rb8GY86JekxiGCnlyPh0v/2ZQBIZ3AQ632fLzvRxeEonsVIHPBTH2
7iWHh7ctTODSR3/3/9QouRhlvTnK3kYsWH/Ny+DecY+WuKE8iT6K82X9DN9cCw+2RfiGnB+9Cy+F
RmBalcNimrHvLoP0lGio05Q4+KjstStBguC7j8wnM2vvNP5syL7nCLWDdYHOJfnNoB8fEgtNloqh
AHJq8QMaCjl0o3ANZpvp/yClOiXrs6dmjdLdv1oejT1GNtLhvrHHPZ09woTjyBQGOQ4v0dej+IN+
YgXbACgR9+Z4L78bs+dpOwZ5ALPiAEcE7AZUjiQr4DmyfiAHzqCYZkIFxiU/2UBs6yhTM8ubizSO
LTNxFL4nF+r777FnzADyVeeL3+en/BvcZxR3KL3ooWZ7++oEYJXbyD+uc+ohgYbOqHVg39pAfZKW
tFEqf/q6NsKcKFJY5pmIRsemEiKme/mhNHBUAo4fituwOhtJV4ljuksZt5anFuuEAua9gNP9dAlM
+vXzVVA6PwdQxLD64TkXG1KAu2vzGq9Mc7PeRacmek7ivX4NGTDprIcRbRA1isbw6gp60ekD7wZ+
TPZFBCqK46hyRGdcOAatUxmkvGofPHDaqwmoKDOBBeQH3wZj+nHBVInnUOIt+d058z1qJ2xRAUGy
iOvJ0zNgXcIkneDX/AUkjecmRQh7XlzktlFRGcVmpM7bM6JDSC3Q3cxPB1N5ePODcQhl2njqGYyg
olvyoDC5tDkblW6JGIIvk6u7+Rif7ZadqkNtKAbtimUPxS0xLABKHfAyQqAlYQ2dJF/pLul/uTfx
HZdVc2WnvhsHAC9Xts+xVz6Cx71UPdX/ZL1V5lMoWAv2YK0SngHK2jNCnDM07ftj9sPVwDK57nrN
SP9ucQA7gh6j6VINiKl4/ykp6KHaFQklw8AgzB6FYLzg+cJiz/PaeUEU+wHXG/zPQdTDYykvsLdm
oApgINmFxtxsuMXo2PB6swIw4ZpkOTQFXRwB/+ZJNoM0jZFJbFhj8sMLteGjbzyOYF43eckj4Ym+
NJCTNpjZ/E+FqJUAcrIxR8JD01B2cX66Anpob+T1EH+EjfO9BvmLMdIA0dHGLT7HjanvcaNnKXFI
adSLAIiu44eRViegMG7XF2ciGgt4d3NGuk7eU3rmRkBqTdtLk+t2WWzjDX1h5FJCFegY9mrSWAnB
9PC+cdETOSl1ZbVLGZwX8MMaijRvQ2u0fgZLJkiUqRi5vNuBI3R+lMM/iHnWj+flGrjJNHZiGdw+
CETtBHnUMoktWqvDL625qndZXSwGtjFQbVxBQYXysk57lIQ8OpcfMH5K+qdXAmOi/XqBEol0j6R0
bC0w1f5I110mCKRUrjKQZidEhZrzOA1SyY1UzAG1LCFoGhl7wY4HvyTsjmCJli+UhBZ+2mDhNrsI
J/tCoTb12XwBO5wH6W1C+4FSlRNsYsr8EmXIq6THFIdRIiE6ieuIk7kvFTszQLoMgCkeo0WrhbzA
HEg4fGXm6jzH9hzRcLScRZQJfC6lli1XkUTcHJiSdiW2WMu6YqDKMiBRzgStRbBjo2brI+5wNVO8
Fj64hJntzltL7oz9xqeuaW52F96Ujgx6ImKkCtZDIs2s48OyDxfqkjO/h1AmatByzkPH9LjwhtXI
DYA4G+qodSDzDCsGXHmDcjhALK64gishpffJDWxqICWjkZczvLVXx1SHcnaqDc/qPiFYGwCAzIvl
TRd9lg9ytnqYyXYRk8cPBNntuIHJIZ9BnjCUmXNf1C3NrHUSZJeKSSPWNzwATsBB5W6rn9A0SCrl
fDWYjiMXOax2jBEmfb/aTg3oNAL+CNZHGWYCqPTaJamZCfePeUJ5TIWe/AQ2zcbXohD1uqjJ007T
G/K1HAj0kqnehbwDIJH/qdFRO8t68iUar5x+ErtlDnxLp3KKaxXMURv/Hhrfr6tD81DP9U4jYmPW
6qQVZfXTPMjkN7unzr29LmX3tkK5XraFd681b+xakKzz0REou3gvN8htRTsT+iqqwtehW+A0cMts
g9Q56MQi9GdxbTja1R0GrMd5VWDwhZVDN3wXGPmsu+9/PX77REgWoc8GEhRe3R0OpAvf99zDa2lE
BfnmTMljnTkbHYHwIJMxM1D3oDF7blUrujsTZqoyKVbQkcTz4uLv6c6rtOkEuuYWRgIlM4KmTFa8
6Avpmc59zPeKtdddvfZxQQCGq4s+0wof1ohvVFi+6qcIWxAWcSm/r35qdfNr9okieH72LD8MhVu3
s+zX97Eh+BgGCTA3I0l5GgU9A4fH5xQIM10pOa9i9QzcHnmgGc+b4wrrcaYpECRJdrYH4Z/4PiTV
jibX5+VT1H6YXt3P/prUgSXuX/1pBRE0MxGpklUu57+pQ9jcdMULJGcwg+48LL5UEMhw26E7Ystm
BbrsElyQUO8igt9q5IYeCyLCaf0GQkXoLnX5ifR74YfTsCsbdM7mgLw4s0rRQf7hMEsQVAuEXI+P
N7He0Tuv+yAz7eeukw6lsvZ2CAqh3bzLNn5GOMA1Wx97PT2Er1TUuVeo+fn5zn24z/9a4M5vN/FL
vSZ89IpOmJdGG70XYMyr8RnZkBRE1sMoD+fYqccYwC03C4YsBYI3bDTN95cLgR1K8tFWIbO5O4b7
SdmVqVklrl+TVHmBWFGKvyErfpMAoR7Yc9Opuur7HoD2MThTJmJ+CM+GV1pQhQy9c89RbwgnnOY4
NqcOWZLdc1qiR7zlNCNU4+k4MD62cFjme0Vej4ub8CD1xlPuye2BmEyJYK2jkBBdh6OUU2FXAu4Y
EHp7SQjW36yGdEm/EcEK/49aV/mSGZsuK1CgElCvKTFvJVsJhgDYGVKFNhjcD+mUtvmKarMa7wsh
utIwalqgNV8D+iJy5d8CWco5JI4kcDI0qd/501yo/0fr41GyFRVxUet0uZoD4KxSOdk45tnO3PL8
MHRQYCy/q4vpjAoOG2eySo05FVVQ0Fq4v86g8Jy4FxEWRsHU6UheofrQZiu6DbOOPUgro+h76tGP
Z0ew6cZXVH/R2K41J1DMk+TXAzTCyrwoEf7qYL9aOLX0bYporeXRG9P5hTEtuOpqCCsYcIl+Ie5x
LMxvNvsKwLkgkqJGTvcgsuYoo+6XTgnduPISL4gOrMIZuXmp8GqbuPtj/oKNovUlXJfCG2DiGtCs
McXluEUMonhawwc+FEXJgkZwSXVXnxuo+3Zp1s5+X9u1AWall3so0/cOh+PnPcNmmIDRq6tKJAmI
ztS2AcqNnzVJSIn1LQ1YwX5oVkrNUjaRS4QvHP4xCNDHG54XwnLNRbtZrrFQwk0kq5oo5a7YoA6t
b9Hh9v5LhdUvZMfSCsPngNcNp0URHLd5h+/TCpC8po+/4xTvhPFIAyLYSEKTDr4wI+RZwj8ToXtg
R1RymbgK2HMdDwBdXGE03h5jlHr2ObTBNCAIlGFylQRXJJeFo311cdQKeYTrHTfVm2UFvEx2vYnn
7ydmhCfiJXd6YmDJ6i9VGyeDNXSWXtBjfCvdxGdklwiGRNakDYi7Ey64jDYJrSeQbui0URbqzh09
3fIpcSO+/JZc9uvwGJcvOEYeGHgu5Okw+VE0C05RootB1M0b0PHkTVXqXSNoMJgKyLebl0zadYQZ
yOOArg+Rgc8aFrdIO2+K2IqaPrXGo2YhJYR8to322OFKwjJpt7+/MGwiasSqJvWfHuFMu6rnekBl
CzF0ZSFrr1PrxRf63KDcgcHaALG8g4GQQ5IDXuIr0kgsklbqWbby0LPn+Yas6h1B3sLQptL9g1Mz
4Dd2oLumti7hOi5xYCvEvw5M61DhcK9Mx/P4vy6gVYs20f6MO6c/xONgE24EMRv26eHlpzZSKYne
6C2NjofLdueHJgS1EYxchUeBi9izPVDB7px0XA3LPQOoe1skKAhjQ3ZKQdAOPIKSz6JJZXescfVf
ob99DYl96MCpvVwIEnP1gCD1AcphjFwPDXtiY1ORN0JGO3QrU1qDbfv/gy7j1+NWk4z8T+5J1Ckc
02TaXfL4NnA8i7HlXManCGyeWY3Fd90o+cBBGYDzM9Q2xzgB4zIKhq65npTz5ajSNYyL5405nblm
Rp0sV1jfA5hqNhZomPoqoeRrD5HpUP5tZrOExlwAj1Cs4rg90PmBaZp2JLJETo6RiNy0aJD5m1mV
QViHN+7s5unZrT3OTv5dc5z6tlfRMweu/yFhoeOwTxWA52R9BFPhZiwXT94nCjICG7L9r6DlEBeQ
2daLBxO3Rm5R6bYeufKTJ8zor0/7wq36JcXrE5aepZ64MdNDZhWIgXmA6JDo3jYs/b1PKr+eFHD2
p3Wo4xhbi6hZcUt29uwfjGZ5GjSkqNMgRDTqV/Zm4Lk/tMtAd9eoGmsqEvrOrQlYuC8JT23YtW53
OU+451YzgDRhud10r1RJ2dQtbkqRPp7E8lF9gu0fTYpPkVa4imvexIQK/TQAxx0s5FrZAoXD+WJi
g/uKpE4QGk2CMyGrSL9tGP+a1VtufwUTtaa3wy0jkUFBxUYvNrLLCzSITqatJiL0QvDAwCR/SiPu
3ZeRdraXjUkqfZo0hfYiIkaYoEJayPNeoAM0JNRunK51vGA4mMyj1NlbrovhN6vQhA7EDr0v+vh+
zMgS8/8/lNwI2PCWMoLM5GTrSjrPfx5GEtFfa8wjvmcXZjgnsLsyqCZrWZEvIj0IuQDowbnqh5Tq
sOom/zazErVP0cqdr6q6MJed4rFMaPociiHk8j1ztpmX7RM1EHJ6vxAN6dwJ8z0XO2qyhQ0nTVlQ
UxGuF/cnlsdDzGjAPiG7Ae3EQLvuqATngnqN79AdZNJN7oY9ML07l9U2c5dN/GIZvF3/sgaFUClH
w3LjF7V8vJdHg+n4uLCooAMiTdRw3IWeyN01a61U01+IjOcouKaJKklqE3iVltccJoDAaDkEsk+U
Kk3f4oXPQ9fYwQffAW+1m0TqZu/IQTYIyZrkMALO/t3Qe8vVtEtQFWLPIO3DnKQWcM0GqlL7v+Tm
02Gk7HaU/C58NDOM6LEGtD/DcjvlVxGbXCztBoJj9/huiQn6O0v0OsJDPEhuMiHTiyOjKsoRAhRy
Ie1h7gdDvYYCXPCN4/fFLadctBL9889OgkrVMDZiJnF4wy/i5gKNhDRAlwIp1xNlTEJluN4iNGm4
1MAkqrah1XhfrHXkNvIxdOqJJe6lmuGa2kF/gCzdIdiIlRBBXOHgZdPpSZZacP6v7v2S3w0aA6bs
4JkwiIso1+LkXsYe4I/oEVkvG113Y5E42tyKX6GKupG581IcXoqSdsDVQ/8+RSwZAn35fAZtrLW1
dy2b3VTO3qVjmGd8b7C4AyMeqWnK8ZTmc70WqKCypObYENQMai5axKS3bXa8Nj9u6qr5QUGkwBI+
Jk3NpiSJiKR3MSkKYISRUJyaOjQTteyFiibs4UHRYz5PB53NDjmlFT87tomql7IUnWef/PVRfXl2
/MKjCmHNDLvBZkLsO7h3mz2TdZARdbxJ1RjEYjhIGCdc9Day3NU2kGEICQQ6HthIIcuPWx2EN6ks
9WkmRhskzfz/7oiyzzDni4kjFeBdOLFBzpoNgUlzit1RuZlkxFxxUOu3Q/Ixy2mmnwPYm3pajCcE
WpvAKJw9kaT35xiU7wusD2LQ1fu9L+yTiZCoEzMTxnLEkdSYskyV35c330+YNPwpRirzKAW9+Q9K
Puns4g60xZ6HT5j6MeFX9J4BclrBb4XqzM6Uddy9G3UFpKmYv3EWWVscCdsdHQPfe82sLbDcOSxJ
JnsWD9W7kB9y8jkILjXAMyW3cJg4/akmSutjEnjau0CHyP5gwsovYKrSQPFrGRcqOdbAMqfRgwpG
TpXzMwnNNDvhZV1zpJ5ZnU3K15gQjok0X1PXeU1Oud/vnWBiYBIy6xc9myn8RDJo9y2HduI5iBVV
pIWDydG7g8aOfPz0H5TyU/wty8edO1LXzvTU17NmiV0Bb5m8kNbq+ANmd96BDTUd5hORWY+G5x4B
+Ev6vb5HjpvbmUkx+7l53N75J4HuwfpNdBuauRrzQigyRXeM/pIMKD3ezCJ4HjO+xv1tMJaN73sE
Dkidk0eKWI2mhLtnqxhNsunZiqqoSPDblJxDA3rEUVRIkpVd0m8KSeo9IUe5jxDfzQec+dNuacz5
JB0wEkQjvnUdx5NIXv3F6n3NZTtAg4UUyAjUt8INpyYTy0oef2ixEQjNpu44xZhTA/hHQ36VdPxC
QUnDG2+m8+9cvop/rRofDg4gsziGNt1RoEWPpvWOGA/cegOLd1VT/5NZ3rTRd+PYmMo70m/ApYHN
GB1wNkclLEc0niEW+VPHnkPKkUBd2KQmja85jhhetYst9wbiM1dY83sy+/jfIztnqCEQ9Vp5sKDv
KTy2iwy7PeY8DRndcf1ivRFqAaTjoW0YazGXv8cvgHpOWVWwPKVgJoyOXrO1K5TGOShEIyiD5w0G
i4dDjxYJEJy89/iTdfSVN/6/NuFUbJvMtMWtgOlvmxQae7fon34hX5Q8GEAt5sEka1wF+HS/UfRJ
gSuuQezh8o+TbebjB3CaiYEaO6Gug4y/Em0aDum8HvzdJ1zANaAuE78fMz7XnhRisSucqytdi7NS
K+oL4c99ajI8Pc/zNHVH/WWBcSmu/GGSEmLFV3q3023OP5WLkjh1LDWCWSP54uuZAVIQdcFLQzzD
OO8xs5P1HkwnoK4+HtgaIwX5UdUwOHNk4cGaWdbsjnyoK/cJyyFfdQitank+GNkDcmX0/5O/l/BV
2qLiOTlu6t+ZYz+35SQDoLU/dZZFdOjahFcQDdr6Y8xgyOp9XyEEZMIZmo8xKFlQ/Yd0kyufqwgj
w6NtowkdrcfXD6AlPcrXzZQzZp8+zt4JhgAcx2/yw5h0VFbByT7EhsSFkJgEowEhxDDeTvlhN3QX
3jLqkXZikbSXQ6crPadojNAYwwnKYAoBgVMxg6nJKofSv/GfZKYQHbBjEarXMFBEAz52FhIf+EW/
O0gbNRDgtBB8l7upbAsp6jh/lgBOpg8FoodAu0bXMi9kDADE1gHJAZ0p3P/YFEHXSxuQJGuv8AEs
6Xbdg6OxJZiazFK6hHeLLkyMjBzVz9VunpGZxZtl0Rrm5o7QtxjKlwcjQlKfppaiRyx3uoULLDT8
zDrYkPBSRPxOe+7jRZDn8ulsQ+2jdJmRp4NW8361LgLYBob3xop83i5JW6j0isk//iRjdHkz0eNg
S4r1OOAEtDN6yuq80/5WN8pmnABNYiH+6X+YGGEMpcoYV/EwQUMeg9I17/s18XQuCjzVGK4pRzMy
LkZoomMZsCXrIQGMm59TCD0Q6TmQsCqE1KyktYQOlGnQpt3mM+iJs8D4gd0WPxximg+jF8/SvbR/
8wrmHIpXEamIesyt8pdRAJxBWmeabwNR0TgEBHbwP0teF/NG9DcNPRZ3oQtvBzT1P9C+1bhvbNDq
DGxvsdbLidznrXux6r9zw2JNJt5d8YTB+0lcbDMvayDG1ajNG2nfXpyD46IajNHliL9piwoNCRpl
xcWjw3VA85oNF1r4FdnGhQsaPWxHEg2/G3xAFmso5TdqlPl9dx0ym0ISWSpATQAMEzDSNDdF6Z6p
DRQLybgvvAlzd8mSylkxzSf1YON/0+KR+bBInsIHrBD7Adnvn7Mzi4l8qtp0wxXjz+nnhPfKQQhF
rpDI5Hg7BZSzTvwTciIlQLjh1ldKJTeh1bRMtxv1IvPEQXF+wzKqseFeu4YWmwqmIv3KDnrKxDs0
gHk//w29tQEXwGoCxGOAihFu4W1cUgkFgLXonCWZ98MaN/s42+/M1p3ZRIHUJDTTODOTtUFNUHTB
3QvcDU4r5aPFpFlkAvjN8LQ21mS2fL7OvZAjhzzPhPX0tE0mIN658wZxD6CekA/+3Ee9RJIQFABl
uMr9IB8ZNWCGlEXdeC79agRhUiaseickB4o1Uo1+PevC4SAvuIB/TAecmr4vRomoDbXT92FS3nrp
ew7tWPEoe4vERtfReS7m7mo4trLL4b+6HNJxP0whZWaxRUP/RUw3pNTNdchfZccCwSVLcoWCnJNt
ONmBrI2OTmBq2gZ3V9sbKFUmKIZ9sC87htKEx91OyuesIwLvqZv5F7Z4T7ZrFVKJbEcykRP4NIEy
thnmNFVfIiIoEHV80jPp2nLua0NzYhNRjCZ0uwihLS7rC2IgvtC84UrFGqI8VmVxFvpF2L+dnt+U
JPfoEqsRYMvhiXIa6T4N+xn5zAIs+2kCSJVtT95dB1ZzIKpmF1YnPultmDy5jXwwgRG15ioklEv6
yREuPMD7DK3aJvKOlN6Y7jlTozxAGR+aVkfvk+WXf+bcVi7SYDMWbDwzS5pFdWDjzt74wQWIBXO/
qljV19Le6MZ0ICShu1xYEC2tM7qk67z2hpXxOr0x41nIqDY92PF/4Ss9d9XzkGVpYECnf/V4MHfM
OWyr9NKbEJleZsTYuY3JsCwEjg046ApaEDdxEtInfVImcaXDymKAc9y+37FgM2LeOrqqmoOAMyKd
Y1j9oiuL/OBz1zo+QfWHgpGn33ExJNyhyNQ58X35FpoHKalx1VFc6xmAbg2f3eX/mpsVwyv3WJC9
IpBb6MDr8q2pxeIoz+slSNqDY5u4dbAoOPCenSMeeXNuPyww9VryBOiiOpqgdcPQ5IkUoGaDv8DA
7TM8kEONQx3TC7/O/AWR7e8BSbAHy4usopm0RWPk64YW39OnP/SxXZgqqaU8mSWB3QStQjKXhmkq
sHAUAf6dZNQ2ZNGZHfB3yEft3Wc7Z1ZQivq99eg6Suuh9D4hQ5RrqJujS0D0IhiyHSiwSWX5Qcc7
Dt84KNWEu2X+jYNEcP+HuQc7r8mEBL79QX+KAOmcVJ485iEkEox+MQSGrckIJsTB5TedYZqI0uqc
yl/iP7hoZko+0sn+eCRkcXbuAT9OazkHxwp7XdahODSYG9K2VVeLYnlF2TokjyAqPt44HFtsMfLG
8u22qVqVZ2NJzZVKggOM8PrqJWijWochZhLGzymLbjtFE3d1k/qgJ5SdCD3hqjxU4SVMWHlCpOUJ
0coNX4+hzC3ayn3vwx0D3G7Ixa8sEpfBIzCHzch8+ss6bbrxkV8tLX0OXxwGxgFrczcumrMOS6mj
rLuWntY3Ji9nVfuatyy23+FJlTrDyASBkHxeyrMi9btLjg3zeUEHJfM3MapjeNUAoM1vVAtyNFuG
1fLOlu4il9Ee6+YuNE95dKCxskg3YXb6uORYKNZl2OvcPGcyqvt74laGZF5UKOTtl1rwZglPzS61
oYwyO9OEEWVo+6uAGjynmh0Z/6xi1/WOygs4fhOFGNAAqZLScosO+i/bIl8+XyK7HKYT1P5yptWq
WaKHKyCyh2eERw5RbC1q9ScxvOrfji7xO2Mtcd1/t6A3Cfe9fphGvc+LyIRdpr6i0VS5+ub7S2Lg
ylJWW3aiAbhoMLezWBrwvbjxcxzJKK73fr4gn0ipH3lAkroJBxwB5gpgXaMibXarp+InxH9DjbEn
XOYNDdvVMWw4Jc8I9NtV07zXLQ417PgCcor9eC56WTdfsHzU5hZoO6AVE7H7/jVExHdqbjvCoz5n
kUF7pRjnWsWphyhd7PVANOevZxtbI+o9+6txRqmN0oWtMEm7zB2qE+BtLFA7khiuBtTKylP7RDh+
ZMz1aRNBFDBm6YelVkodKNEMxa9eg4PgaKIjaor90g3mcPkRrco9HpvXMHgolu6FxGeEYsDMP0Ap
Qg2CNwzeRguCncCpyjRQe79kBQk5+YMwvoAgJGFyYg8505WUEmHr2aRDuKgZtbl81qUAnNwNNfhh
F/zJ6L69TtUy5z1H8uGHM7zRMCPXJV+be7NG7cExQSPyKRBHM5LQooQ6kLudHFpxjrpBqN1oN6AI
ElMtrXLKB2LeLgFBfmY/a4Yvdvd50rd0VBSZhZaqEYttAj0OE5tMKv/CQ36LT+rBAH+G0fDdIrTc
8lpoOWJOqrcBR9D3S7MKdzjgeJbvyHSC+OQoNTHe0dKsP69iwQ/Qd3qyeWRxfoq1WiA+b0uQJK79
7mhdWOOfdxX0BjXV9ERDc2n/un4ZYLdgyqJRYwhmGoJpAAI9g7i5NtzooRswTkGQp7e5tSwvWCdW
xOPOvtcVa0tpP4dYPN+In8WQD0ApOER6N0Sp3rAdmcW+NZkNbm0P6+2cJ7IaO0Vbls41H5r70dSb
3l2scIcsC12Ud4Ut0qZfQ1nstiEv2n7WkZdgxLUGmYJLPuRghm7K2NvO82hMMwWVJlbhJPIn9wpJ
okwPPTzjiMtT+k2uM1xGQnku5EDL4s/pz+rdFCIWuOdedpNOddtdHx8AplWQ1E1Lv+fQdCWBeCkf
uCgOhNyazC4zjmkX/RkVsBNkDRB7ZsWs4IjHNxCzeAWrmgefPEbkdpGGnY23iMehwt+hQmdBZJr8
p1Q9vFxFzq/ejf1re1CZmjvDRzPxQdSCKpktILNYMsard3whQ6R5ltPW2NSc2kQOgO4I3wHULCbk
OQzVUo78/Y+Lf0yDfjrmteDkns0OJklTXXJZ+6w+Mc1gSIscFNM1aPHaEb6ALUIczARTfD3zveE0
brIBcznd6Z4C4yuL/p4/nqVHQe2TbmDmhcY6/qtOacxoLApkd/I442bM58eri3iSJzJSe1X6VxT3
1MDM/TtQDXJl6ZdRqzfiwCLGoopPUcMOUwIY8f7JXrohWtTxEWPfHCjrYazxJskBA/16VqM7HVMk
GC2dgpEhYWlOudmvU/b2/HHvPOPAzdH/6q6I65ecGhBnR9xGWs5Tw9kXlVG4EWyl4DikZefkeBqs
TnnwOMMPTFkdImY7AMvsygY1ZjHenJ7W4jhaTdesmNusX+u03FayjnBwgTGkkPZIQaPlxgd4i0s2
5fHpbA2cqCxR3RIK/6I/Xr305MCVkk6SemfurKri+tSkD9sW4nSlrA9sm0sQ59KAg29mrrzNzR6b
3RGMalWZRF0AOLc+AdxxIVhsaW/HQLkkD5lrtjYrRhruYb1Wa0iHwOqji2fUan/J0iRfHXYWNL6h
ebY4GZoe4dOzkDZDz5Rnx0mpWiHzUF4ZnVH+GeP1zZlTUv2cNyXxweVx6SB/StWEvPUOuRm4bB1O
uVz0N+ef2KE0fyNy8MKGeVUGU54rUci1CF3JtLV5Y0A18uUYx24plMJZSclRQU6zYOx2YGCV1iDm
4SFNEZGkMc1VounxPGGDJGHXUlXLtfIJ9DTki3lULSF07IMOfZ7YAIG7XOrPmxe8pFSM5JaRjBJ3
W5Qzk9qmv32K2TuCWJj5V+yluwXp2IgHptGggopDleUyQHJSEszjEJtBiw88DqH28Ta5Te3IsCP0
VtaHlUvc2BwdvN4kCxoSP6FTtvZmfatxNVNqQVsJIQBV0lPnUuf0EbP/U0r3xEN4ysFtUIxuFlwb
E28GQXDtnJDSl/GmqEnb8MufQ2TdOK4BlKUSP18oSQcDMOrGetYKMwdFBP9Ix7XNAzylCal2eOha
pWp65hnemkv6haffJzXpH8NUkAioLYUQ5eirkkB6Ww1QSZOxURehwNJJyG/elA7ZqpORmUnzDN/2
LJIXAsfTPlAhI/BdcYjOclXGBk1etIiUNdTBOJIQNMnW76QzFd7BcW27tITL+jVEB3MA8lREcQs7
7SKdin5kETHB8OMsmkgu3T8q2L0cHU2JCWaqAppEMCcHlnkonb9grZY6ubli5gXbKKOwVJ/No1IN
NoMQbHCPdjM0yWVECy25x5UQiHnTfLfTbBgpiFXB5oqm+mBxyT41XpYiixYh3VkUVTU+J1E4fiMy
uqPptJtJph9SjfzlcR4SvlSWl4eFOlJCppHzY+seLEy9ghW1T2qL+D0T7AaP6J8RVR9idnW6mCdq
QQi+qq+2cRZe+QjbHMXNHMvLcZGL2rXvodJZzytHZxp09aaAL1WP6BA+W1GsxBS71oZxryMQsQJk
tIgT++27Ps7U9iFSM344KlpssNOu3IEiPQDuTHaPnEB4mNc3Cy00t2Qfc/OJDozL2EztNJC+tgqO
6XK0qBlkoA21LZj/pq77OeQe3b77bSKDe5/XUxkFdeq35Z8LfMtYhjOvnJYvR0WnAwxUr11EEbf+
GXwfaP9NsIxoYyvxWcQEi1P1ShMSaNg2fX4yENOdHnqlR1WhGg9MHGxdxSozeYbuHjxvy6Yc4YfI
Q4iXtYCYSMXMb3ftmwuDGAiCzcddi06pGjB7DtaXcd7c8B6pPCZBxiX7abqvj0hsH/cbw1y93BtJ
INz4gIjw/yZElAcacF3Sr+OCPbwwz5T+yWyM4jLcrz7nlMihFoJzRp554/4rE6/dxI4IrSC2e/8D
jCRHNDnffkisbARZPKVm3cTxXzVTGMjf/dwBKwEt/LnN+H+Erbb8onezp2hC4ez+rSJKn0X/vxpG
iQr3fjVJBUlYAZauBuJjyNX6qPIb9FRQZ7R8J/HBMEyPtFrH129p3LUMLtq70gWlbxSikn2y4ZcB
y13TemJGxK6oYqbWqmh/s9sp0WkAMvvaeQFAEP+eyKVM8p2IZV43C6vwak9gHawwxyUAgO1DavLv
XAWmkLhQ1WMFDNfiPYgkfgBb8mnkPUEp0QnGba/hQJwg8TK5jTmNNC/xRJWc1nUnjk4hcBF3NWhs
c6S43qxEt6z/E3ovZ1vE1MGboKH+qQKIUxbAy96Zk9zxjO7RzbKHnBcW9+HSNfpD/o0h/+5E8xiZ
brfHrwQo57n8tlFKo/1cyT1yOQMowDY/5wpJ0xl6PM22MJsuqnK6thKILteDU0xemsomMQIICYbu
FG3L5uCxoXzgMAM6U/QlnYsNpsmY461sjo0Cvw5/4L78BWnKtAGSVHVLeV4mbV3HbE+TDaxxRzRj
VQcuJ4xoHbSAB0Hq+nzOXLd0arEMtD9y5QLHllOhraFFifV7KyCfOUHPfAKvzxvUMaUDNHmN6lmq
o6l8wZpCKgtTzhDPXarf1BLvNR/AZt9kt5ClR9NLt42aa2OBo5nxEpZd7KmpWub2mfqve5EWPTNx
cpLHG/bXOIgEdNGtN6O5Urlq11DNKk+HE7RkKB0IBdR4rzeePw0lYcOu4VZnM+q1XfRh+3thuA5r
vgv/UkwPXiWS6BOrB1k+IFXEH9VRKFN3/7hz9k4cE0EQf8y2qoAU5FuQU9lxkJ5FdOv997ereHog
TFnYu9SffmSfg2WxrZW7fRUKNptgTnn4+/NejGN49CSrGdG38aU+oeR22tRjb46I2k1TpfnLKIAx
Zy6+/fWEjk9v/mNUbQnUSwJLYJ5wyuZUsyPwCPcjNbO+y3cT16yMniqIQX9EjCKbN50k7Uz4l4a8
4SO6cH43tRUWAYWpuE2r8v5F3FxzJbK3xL7X2tclHgkD6lmTft3Ew8ERqdKlBZ/9EWAP0xi3RkMu
bTPwjQuRypsdHUotXnkisUZqdXQmPpKiMJXvbFr67lnbV98fCKjAt9NrolaeMIArNOu+LmM1DQ3i
GT9mNTkxuJHJuM5N9gwxlzj8NfaJxDcuwJfSL4WhgGplMii9pGapFIDRJ1FnsUcbCrNQ/HyzJvr0
oGY5xHlFr2HEdrujfl470daOHV56Yyu9LA9vZpH5i6fEAGtliZMYcyWM29XG1viBvVCbQtMIKFIC
eWvZjuZfoZXL/cvLlEMeti3n0pdLe3k+exdUkxRE3cmLXIQ4ZrtuRPAXSheI8GCN1v1ZoWwhES8W
hD0ncJ6cXRT4iEWXh9XtEfJD7XUjMeankY683Cozaun7do4F9N12jtJJluVmRjcwrW+0kDo13g0v
h6qLq9Biaxtpk8E9REZxI5VLzUCsE2FywbPIdE/HIWkFz6psrTy8QPtHrq86VVSkfpmPcmQKs02X
/oDTyyExBMQoVIT+j6cnNku0l3zs2t8jP47xa3jgFVpcIYJOyt+KhhFD3jm+r/sEMfbzqboirwCU
DDnqaHIRwAlRvyeRoc9o7hxCKnqPISQw8nRkR8njCVW27wQIjuSY+WPimK7TpwFNXP0hJYlksaYG
g3Dm90/07jNk3Vmr3sljVlstPPYHN+Fk94x0GipycJpHZJLPUhZtJqsr8KunM6TH3PyR3io6oH/+
hv7MpNjPeAF6EttJAH9URkD+blgZde3Pg4lUjXc6tPIkycWVb4fwWO/fBTuoCoecCUsjxAnYGNnl
pditpp0kJc7D4kGoQVdOJ2sVcfS20wAmiuJamZe4drnC0+TQHrQCm48Kz+G9mMoZ8UXTy2WpKDPU
qdhsb7k4UDUiP3x8Jx/eBbWqv9a6kcbzkrnBgO4AvHmRbW9n0MwT//EVXxQzLbFgSqEyDSkhAohc
AEkg21LTZF2yXhvzkIj3BKInbqRlcXQG2PNtcQVE2m4MhOLXkMrF+kuw47spXzd+NVb5g0AvBYdI
1vXoP/LJg71DsrU8INGL/kJup12kZeqJEc3V1uXpFYX+AevCsIoQj3pNLDa04wIHVXgQPXaau38N
sGDDmUKwHgY+m7XKlQBP+qecPDWmQ/RYZIYaaoXNij6BDxEdKsBLbzxy3ghAPIEnSPxdy7oZTtS7
1wB5z22ZyaRgl2iYBaDRtQln061lF/Egjb76xt+2ANwWz1TkjZb3kIhuKFaSAkms/ahd+gCO46Yi
KLg+G9ijV5Xcv7R/tR7gtTJSjQjj9ulWz3CbCFDzXsAV/03RoUJk9fSWq9SmwIRUlnHHtOkTQcC4
Fw7Fgv/2KAabkXmBDPkkspPbxuCI4AckxNZ7JKZPyH3+mXMaNzCiQKBe2iZu3XRSDWps1A74kb7O
siI9LN9GYOkoQpmJgWZCX4A5bBdy6P1GAGjATPtrOYMwH/Z8tFH549cHlg/w2vongCx15iaEBrU8
BX4XmdqPiu4Iv7gFtTdkNta11F3jFk7VbzaLCzFjcBS6X7OuKu6+9Avr7tgJSHKC1C3PqcAY9tDO
L2kGBxkZsOR2RcpvfwvmF5HhalayJ761hD0twP+3raCl+HvCx4QI3C5KMBB48Rrp4Q4fyTXghgER
FEkYnPh+O7/wxQxWx6UDzl6gbjoQ1R6hlFnbrJAOqDWm0Atfzp+ehQjRlgAxJh9uMLsXZImoncoR
QYR1b+lao3mEE5exoSJ2Nbo+/Z2uS+KghmrPessuQmiGLf+BasE/cnJZAIfNpVgDR9BSZyVGBZRd
ITiPrWeqXIWNyiLiiSqmAswqnx8ORvSnNvQFnsnjbk04xLFL2Z8YOWF23o9SEmqtdje4VZjvNUZf
P9neIY4wtkZUgCwQA1HUxX0gxIBD2WMDRWMquQIXnwdiCKP+kI8fPhnxO/tAvKoDFw2SugLF60OV
LIHkdbaENIGuwrccHlN9XPN4QhYSQNDGZfOVbS5LnOmshsVeidj1r6H9oHCZIIPb+ioznQ9EOHlA
nIRSxffTH+dClW84OA6QVj6RRCf/1jLC8eJqLmK8hUseFANqSFr12AJtYaT5NMKq7iGmvPoz3fa2
i1fjZ/jh0HwtbZhxIFytJc/cMibiDVBurBjXNhZOkU8b74IKiLBuaCTqx9o05794oLVJWP/RiJ1j
FEXkJExJWySsw0NqgC/8rglAhzrAXL6VehCpjfcYCawj3VqhFBLhKkdJngBhOUHcyIREFOXv6qJ8
q8SaZahW0vUwNdumeeQhutU2KfTIqLr7hqQghV+yGr0cBg+asTTAd+PJzmjvxPRYfri6vV1J2ZV0
Sznjge5ig785ZAPUTPwjVuZ1h9nY5R9c8UlLBronHLV1/BPFrsMi9yaeLJXhh89TjowK6F3nt71t
wyC8te/FvM7pRt641fm2RNzXN6lnl6xgc1l8YaOu6ctP1TvqiiVxTXqHo38VnZGhamtlPAmgpgTX
njur5BTi9JpOiJkY4e32J6jH+GRmBTcylnXfnzn5U/6erJSz5JQCOSdZkrKnMVa0ATlzHeKV//NP
BrSWl2lvGSl9wQOZC6s4XF1HULZnyCFwGBzM3YSRoQ10CNqTQhzXNb3UeVW8hMxAvHUtLkxoNY++
HFcZiDiTJ7p5fvq9q9MnTiyAVX2UUOuvzazmGesGiu61HNCm1oHSavci0612n3GEDE0UyFYizcIQ
hop0SQpPEhBgmwUEFMqeHQhi6SwvymwV0hcvdMAJkeY7U6ZMkojFO3omjVq8KEDkDWzf6mVivxvD
gyfZ30CmaYBVfp356k0mG2UW9GM4Jeof9ZLAfo14EkGHvIlVgHOfCJWRrDRcX7Xj7aYZl/7Nai7f
zSGJOgeE7LMjmFLGqGc+Ps9ddYCMifoCALOpjzPFpL7vRWMLcJWpW8PasES+jPAHk0kydyN7yTog
zLS43+Y9ofV5O3+dg5fJbl7SkU3dcsGhjuUPuBEAZQhMAuA/sGlea0twcCwN1c4OoNqSC9lT2jd3
WOLKkjcL3GDY/5zHha5iCMyYub9LtUDGmsv2hhqFXSwBFE9+LIRndFJAj1aeESyudL6JrMa62Cxk
66P10PC0XNQ3kAfE/eA80G98Zv0Rxqkda40lfIAa0j1pEt7OccR4OXM3eUM5nV6PXRZcRgFoF0cP
ySmW+80KymCBDBopHMH4UWWFbawYMkFS6k1/Y8MDoQDzEYn/qWcwBbUIjN4XcseTckJB05zop9Fl
VVLDJ3Kgyn6LsQwJHyg5s91nfEN9n6ihnoWWj2QCzIQU/vVJM5e1OFivbGxPGAp4QKW1IdykEBQq
It1T1PMIp9Av0pulZuhGRvq0wOrQo26mzfya4Rb27ZUJEYZjzHjLJFfRZvVJr+P7vxxy2CKaCAVO
k8YZTwMrBFmyJa3W3gjyWrVRTu9jSx5yMbG90ntcj+xnLWHXROMNzFnzpebXtcGd2BvelLFbG5N/
0d+I4FZM31c7GtRjhwsGBSPUiQ1UInJ19CJ5/qF8hykizN59pRQSolLB4I/jK0gY8Kmx3yPS7RMU
gfh/S4XA65sjxIMTyoKk5+0nyxvGs4x4PbVBlgOesZAzJ5jCrHs9p6ZvDsO9Ujjxt/KDnm4XYT1p
scfqaQBl5W7kXQfN2Xn0ZVmQzSCAljcpHDsq781S+Eel/rYt0vEnTk0ikJH4hoRxGj4rX+Zp1w9V
+dODbSLmo86wk2Y4ccmHJ5ALOc48Mkls+j2OOJNAC3peJ18exkqTXHUAa/I7oWZrXiuL139X+spO
O54/ATz8hxmdaqXHiW6uXUECUEZ5L3q+9zFchjVuNd7eWXpJjKWNeOHY/MZMXB4UEuiepyJhlPsk
3RSxDibdmYA93os7I6D//coePf9ywPZIPM5oGlooGGKKrSeBIv5JUcxEJj9gvSjtA1TScIMXYNgu
54lllLWqNiQ5PlaHAgUdg7OaAncvdTTA7OtP8xrakzPqqEkDy0dRC3MgKhFReWRSoVQ8zt+8X7PU
ynUTcuD7uf4X729pDf832/6R7XDQuZZajB3WKRAw4g6UcRpmpvGnTdG1oHEfb6KvpbDkgX4CbWjQ
rc8hb9AXd+au5rRNx+whNOaW87tJfPrjSxOzI58nv4VlKjgOuHnqeWZ0LfDPlJa1/N4ZXuFjJ2Zk
5M7xpLSAYN7xH+WLs01zvKfVCBZTYZu9Xzjh0L4sjGEshcnEbMG32ny3MrqMqrxDqAZkjBvil547
vkWGoBlyLsuTk4csS8kTC1VhYcAOSYIqG7WpeaQYxWYOnPk06a1uiqQZHtUOvI8pQ9e9zoujcpGg
oFpFquvi43RxLCthc3/Mz7SiPoK57F42WUJS+raOIwYWv/1oSHbWvFSNdKDBE4FbgxPW8QkSxO8e
YuzxP7NQ9/gOdckonBggNMRJYNK6svjKbXfmzGjhLw5lLcAO0CrMlO7JALzpNp/WnLl3VymTB0op
rUiGR7h5C2dpTHtZbSUHSPkcxO2F1OeIsHMhojN+Q7uabmxg+woW21D/+65O/Ts2TYSi3/Cnkyuv
mf8H1JwjImKSlGhZf0Jjg2zHIwA+nk2xPABnZ0AK/vev8deKglGlq/d1P/iiYM7tOSsv2BI7Vtxa
p4zEbtKX2+plSkO+hoaGzrqfvDnaJXZt9VxVvPABc5DEF1zVO8ILcycPS/bjfAJ7ekq5A65ykWd7
uRzABDchzyuiUfTIOsEi1H8WJqlSmTEcXhl8KEPXy/g6EL7O9nTT1J/v4/f6pEvea5sQUk61mQGi
4UY5GqN4XkunyNBY8hfeWNpE55i1hpq6kH4fLBzlcR+dovkFr0RgSdm9FmK/qekX/uVXW7pPN2lL
iwxnHnG786/o8lY+UIl1a30swU61AcESl/phv0K9TmW1j0AdyuGx/+7Leca2jbCAX61Oiy9nA2yc
Oiu6iUIeqg7LV8WRJ5NbCwTzfB4aAmc1lDEINSLCNVQFHUl6IK4QpggBr79L1hxp6NaQ3YovYiGz
/yfCmtzGORymVwvEFH9/7y64KahUD5CzxLaYqcTNoie6VCwK2sjX23p4biaPCzyGNLpFNvkYyxqe
kIO8+H5M3QGWBGCKtpZmfYU7CvNPqU9xybPyZUgrbUkEtFP9yGgvWFfaF+fp3wwqb3ctAIRj/1CG
x0PZSoKDqrZ1/2dBBMzsp2ta4Rxcq5SUbgq2hDJVkXaS4NSC36gRr6P7alAepGHds+gS4ebQeUG4
wLpzm+GMrPS6R7jRR3rukh9vPro0Mcs7Us6ceuMfWWbjCQ4lvanqqfiVjNj+cRs2MDNVl9hiqniW
nEYUDdCJEyZnzXrNvoG9Vje8BEJnU253TMdaNBnW/21UuiDXBmpS2rZlctGw6BnZBkdDvoUboPOR
17ktVEo0zcd8ffZAZRDgl61/MolZ+uV+DhsAJn79XRHvkJjsvXvsvmUssPQg9F7PxGsLBRbCJzUk
xP0rLYSm2Mb9o1IvfWsghrwElnjTg7Es72kdl78Rrys4k+io032NqtSqqgHuFRzGYJEPpNwU4Hef
uOm+uIlLKlWdHw6E7m6dJ2sDGVHceTw3EIjyxbTHVyPxvHTJp2XB7KNJE0ujsDAJIRF2MDKBN0UL
8xB5WQJ2i3naiOpi985yAF++A0Gidz/Kv+Q9QPQbuhsmsPQMSTpIcDmHuuX3/eG5lklrJAqWMSc/
d8F7w7OnyVwVQyEgGT+N95NFhnm44FsG1RjEtiIi0nfvtMHMOOIThYY/yKJ2t7e6/KcGHfK6qHcU
x8xAK1uvtUM9hA2T4mALboe5D/0kN4TGXBylYZm/3XQiG23UiTovhCpMKQWRd+MXIvjTcRooZPbi
lqH+i84IzNJH6y7ankHTRLsjTDbm1IfNbVAlXlBeKErxtmoPRbtjPRIr2RweRnFnmHV62EmzUPfd
5cSo0vcKDApNi83rgLt+GpOF36uoXn0qk5Ej04jLuHMkDGz2q9UrqtvJH5trf42vt1N7WmM4ZEBi
Lu7iHjhLtCLt0phlkQYofYmBMjejtNvaYFBOe/JQeUifGBDbia9k5Q06MEiBMOVikQKUMZ1kt2sz
WGQt0zsPYTNMvIRCvRhYX8awpkgs/j/yfbvde2FzfP3d0PQze7JfaClscWO50GSfse1sZi2EO8bz
iFoArw29V2W1RuOT8ytwPqVN1YmhXfC+6rBoqmLj1d0bYVVfq82oFI2ISRR9r+h26GFtZLkaInNJ
iMlW8KqrqbquorR7W91HZR6yfgvdcTLfvEaA/OmcdaNEfSQJR+AVnNUB2ddgfiBU6n505cViCsCM
uje4dcR5ULLm/LIwgiPQJ8x6U1EjxTETwSLNvFa4HEEQunwWr177SC4E5nxG6GxDBs6NVjcoVF8r
4QaHVYZvcxTlVI7F2fbJsAsf8j1t1FAqxdepUiZUCgThY3AK6haYVzNWx35BNOEu8XTvqApf0n/J
rOUA47J/vDYCmxevrmjoDzdnUP2oWJ36Lt1dd6WiLPQfGw0bJUTzgIKMKZq5MJ81u/u/KB3oKLYV
0n2M6U9L8GSKLbIHmYk7m9v8lUsX3v78SVEvfWU/5ps7nw0M47/50NTvxrOQt5z1oNbMiUKyA41I
uDrPUvONkyw0QjyKRIUoOi1jHz+DOVjiKAT39tvFb+OQ9YjfhD6iqobCf9yp9TbBiP56nAPZvi73
vYKQaTcVc0CnUhHUd5Clh4Cd5oANvxrnQxIecAuTptvYNkvv+NiwiaA28Yb18FVPTXy8KCTv7GBN
LLpsmN6E9k2tBhkkEk/Od3uT8AHEKPxpfebWJAj4AkIEjsxKT8OmxsU+ROe4IkCRVkAE3bgExeoF
wapFx9D5211cj7Hwb2X73bXZJxBHcUwwEmo1iRTAKZfrtUjIRNalSaztdDoCaVGRwa4IQJj5GPgo
uwimU3grOJplYiJtlxYH5yXWk6RrLw2zNUS/8+/MaT3tFIjSWFdjAN9RDMLKriaWCX5413eLbKXz
j/Ncy5aoFXqMVhb7PWkB26mjjSlKJHbmvDxQXOVVa4fn06UVFuwz3Omj+I9QhNIrBb/VFEIUZq6O
UdJAjdXaGwSvazgefYmyE9Lrt+ap7J4Qic8l5yrGD1qWevdfkuKnIjPLxJC+1kmMwUO93cDa0ija
CI7pbkkVUUiYdf1pp6+VKmm8BXhS6HKAS/jiMuDGqsMr8zGzxy6KT51L8+Z08U1oqSRolY85bIEZ
KRvx1Qdv7IBlx2cQY5vUdObeCoIUfe+SLClh/2z1Sixgw8v1YWeKWa90UVnPyXLuxCnyWx3+eLvV
biKm+bG9ve+LFng06Vi26T7QS+gQHmigis2bOwC2+dm7HW33MNJyHcMJ3GzIet6/SDWrficit9TG
tpNXIID5dqzleYL9ozSiCBg0r8rfs6R5oePQdzvf4LFTb+WGpEjeyy31WXzGwW7X4O9hng0aXPwm
mKPcGpUY4pGIgnrnHjNxQFJGsPVTxg6E3WGjJQuZpTighY35xZy9fp3TcTC8JkUaxCEcIvFoPh1d
uUgHW/moZWWcSUeEb0LhmjdbyssW5JC/VE0mcIQ05IVaqFO27iwoXQYuMVRVTW4qSsbox9H+DkTJ
m/nUXDljazgRdCmbYTjjtwmkW3UnN7MW5uNwEm9be2/JFDtS46AjMf71zMPirH45SmeRcaSc/Org
+8wlDqSFaDJQL3+NsSlvxt8ZtKBnAFq13r06ar36gKWMjgkYDk0aJEJ4mUNUhZrAaDDs88z7u7qB
lxZLvHh9k6TDDiEZjzpVtgSfOU7xeZ/Mmhl+m9bkntelhvMHyGGndrsRvb/lQG1DCW4P/Ri9nbc4
HxtfLOBh9ZJULx5b/u/QKHZZzlgB23t9L0paKoisxmSuao6LqDROt2QG1U2+yWekK1E2nY2V051c
o6QxFcPkazH8HYCCVtLCJ875gnCUJ2mBx6F+8qXLgLOf0i7GQHtfwP250HlPTVUIvqQ1c3TpDtXs
T0g4uEDIAUpreeOwJ1iWi6A1m+AyBHs6XenvsY1IBcaoU/t/nGYfAa9zwOIosSe+U3SzMwcWz5O5
jetnQ76sFPb2FcKaBfhl6i8HYKSIlpJ2gSd/BzhdsnhA/TPihIPCdM83n5ysTip4KIj6Bh945wcm
hwtTlmOAP57RPrUeED/8CT+wNRTuhzniSv3a9ZI6LdDCvSeS/lG2YgTrzaYy2/oh99m5lDhNiZuD
0hBvLCCEin54HzM7MxvKGT9joxcw0+tmmHQDacGkLfdrU0oqrby5Utv6E4eSKEFJRlsI3HVe68uD
nHjAev3micC+NHSjzeu5QjrnARu+A0sKi+CfhQDIDeVjgwdZBkaPELbjN+jWNcoTY9b92jrKh/3G
tYx52gMc1OEgokFuP2OtWcjfjvm+1K/s4eBYKB5h8mpkVDB7Egv8nzPrCZcL2HLYtVlpVI3qCiqz
5avId3BhfuWDxTa/MW2WLaeAdjL1x1fwkuaKl/ArI6jmDNT0qE/w3bXR5FqKsMGvhW8gTCCC5IBY
ariYA5+DvCPbcbhamYpGXJZv9GDODFsWS75S3KOrU5/nAcJ0wTzh4nShe73kKF/o7H8LqZrv3yIh
Ck7hVwWirU2wJIdVwqoebxHFd0c86E+ZW1OKGQMARcm79KM8xmJWSoxdZ222MPUR7/+OZ3h1IqJe
DUlMK24OncsDAadXvrGBBOX6PMAo9gd+MYuFZyxQd6JGmf3R97wr3dco5/etUfRFxbMrulfSIEJv
9Bz+UgopVlVNHlrhgtSTJYs3vXnZ3sIZU3QksdTpbpBB0jX560IuK9hFmVlKoH4MhuRDW5WOAJGr
INVmAjJg/AEvG7s8TV998zi5GYiR9e3YzDEDFvmjtNrLVrILS1gQki5T9doXxKlIQyekMpq8XonU
5tGoQLiTBvGlQoh1FX1j4SGhkgzItiHM3RG/bgD2rYGJNAAn5pwmcAkzRB17jrLdemyKb2N32Cb5
4yDo+fcJOc64krzbUGrP40Po3eogFBJ/0BgwFCNewUQuPpX9cUBIMe1VSOb9BcFFmXYjNGiSpmHN
TtN/FhEmv5Hku02JLuN/wtTEtm6SyU7I0F2Uat+QiO1iHDaAK2ybhypcEgI7/UP4gLcc0EVNhnmi
G/0REz4zIYzev1gAR1MgHlL4dc9NLFjqsi4wwEsOC/OuGK3/ePmcrEa5brOWpPeLypZnKociVUUS
tHDv2op7kZB8MQ6uOubynwA+ahqqou7Q+GODeOrMIpuGAXWRoBc33uCEA8Fe0XQeIKoygQw9fTIl
0JDORF8l3PUgwl5AZs3MTDs/f8eogRMt0sEK0sDwZThac2i7Qyzipn6RWvMGhU+0q4SOO0qynKBE
cJODXtp/Tf8jm1j7qzuvZwKpQYkSRGaysN4nspFThc/sjxiHHsd55tZljlGzFMSlg+KWQne4DPgR
JrtOT+LYeuraULtDb5iM2i3zeODB415u6sl2TGO6EzFKwF/O018Wpiz2i+Hcvc3V0YJSYcIgwfxV
JOrGHPM/8BmepWFDcU8HbR+aCyXSx3HjwCgYTZkt3oDPGwuRNQwP9aUztTSLHX8komDEG6QNVfUP
oYCwPcri+VhfxPQ+Suv/GmpjNCtl0QtNIIy9VbORlU3rpWQ6Ny/q4Hc+Tlzco6H1qldVif4zeA5T
WH3PytvopyusBexD/bv4MMQWtvIyJBJzDcM74E666JZy/R5jraWk7+0zohQgjh9GPmDJALIXM4a6
3Pd1RuOXF7hsidAbxt3sY9rJSjNZiT9XMufAx0HmIDjFgag8w3H3dGz9pljg4xnlxUfmtx4PNBKP
78bXVfX7/kd953sZN3Aw5iNj83xtXMm3LfWZkTqg9n4Vt+i7gvSgDjznOlmmyfS6L73YhkfxdbFB
a51Wj6rR1f5++4WopaneTqTKnWYVsDEROPPr7Fu4QsDXedPrgRsZ5pjGfqKmtWE9QmFpcGii20Uy
Ga3qVQ2O9+FJCH4kr0YrP5/Vz9S8TQ2EjzpcELys4Eggk6MRGaCq1W2YyoR3qNO7dKS8PJIttYc4
DKUKAitA6bRlvTD9iPILUawJ61C26TOVLh3Nydpxgpr4J668/Sr9PuAD3Mwlj3mhyOn2reVSAJJ/
JiyidjW5/oi+RjwOJSKOpVs1QXbXZGYDQGZtJoMGjBMhsXeAtVlwT5b9PQom0sMJygcVJVMEJHIq
NboiA5+lsUOu7qO2Pv889hqlH+h6H3Hr/j893pF53sAK5yQZPXTQiFpy+lEx5EIc5V/cKhU8OTgk
xmZ0Y79okYi9JXOQlmI35mlQYGR+OFInzt1oxBYRkBjAC8L76rOIGi84hfuhOuKIyxN/9Cpu4Apz
56wadx2VDjY88qkYcdQ62hfWuaR1tGotz2WNuuVR4v//jpo8C3QcZ3nGwGecEM6BCrJ3Hhk5yjfy
KEPLv+oQotFjPAoRfSdPSBVuv7BLfanirRDa9H4HEnRZjiBckJdVCZwkMBflp/nPo1pizGVaVzHh
AJz/3GFOnECw+2alLAYw4Q0BrjJ6PWyLX/DGzKoRKgoLNcuVYYUbeoGAp0oUUgjikQcffl3jHuxL
f/YkyrqEdtBE2ALWXr8yslMImTrUzXTbsdw/xczecY4ZNibaZc5B4RnLHHZKyZVTLJrxv/rCS+Qt
sfXf16huthjgNfZF8A8kwMVuu08mx7qrRZpzFqD+9gPX8csSmdEx7a51vkCIaIrTUlodtZKEiArw
BGO+tgldUMICkku8mgOqalLex0S4tyiMsxooA3lK2kP8jPTX3WtaxtqzVonuBXyma54HVWuZxoHS
TbA4U066Eo5zacyVZl/gbSkeLYJFdPUwCanSJSq2oRBZsQf+3k4lr5hy/iQ0hugD2rjjCd6Y+5P6
tpCJ5Cct8z2ZdQWJNi0SZsKbSoFHCPqzU/pcE/MqCTG/HP25O22smVhywUmQ25fxQHX7rfYMc2TF
YxVL2c1b8+H9UzuWl+Xa+HihlvR8B1RDvNiaVGpzJARiGs9ENXzTqoZ3imeAuh588FSFumBwq1Nr
QoFmmRYeG21UQ9/A1JloD4FU4mXFMP4I4uTdk3ZFyMnjBU2d0Y9+pjIzvZvVZNg/p6K52e76KuVg
FEfZWU6+wsffnJttxbN2goq7nAGBXqDZchrHXkiw1JkI0FY95YLGrhX8Dpa/6pnh1dd57rk4X6zO
p5qwKeMyXmNpnoEvT4gBr1jSIqebrC9bUGbRnNac0p3B03atgXxp8fZwQZVWfJuwmHL8nYSnFfNZ
HaT+FoOsT2lySZBOV+ZOV4988rbzTqCeKaIF4psB/Y71UtblttUtgC8jgX71EKiAn97lHBMztzZ8
x6CEZQfzS7ExOR6bWpzGQma03+O/KBZeaMYrNu8c81OMEHF3M8w9kdIrsDYWAWcp03lvf35MWHtJ
9jhoe/srHP8P4ubXPyn5Uel4w6FLHV5R6eFqS/xKSRM2MKYNh8JUKJrCOQd0pHU7Yx78w31Spu94
LN4OJaqj7UOGmqvilo7iqpYiz/ZVhT3elpeKosLYbenWjT5YTXmQ5PvphvbwYlaSuyHwtYMBYZ6V
Yz9gDpm3JdW+XiwlnBf6OrAmApxAPZv3VyqwLXnWIjjrq+AtlvqWKyKXJXIV/ySaJyUTlIcNa+a1
PZL+MSRjKG6li8znxPj4ed0oL15H9khHRNs5T2lSZHkccqYoGaVQQ47TF6fz1/lytP2/JqCb16pw
MuclXBtg4js+vP7F37joNjqcQAtEZ/2nzcxS6kCOps/QGSQqtnnkz3UqajExkDDRU4NivVTU3ekT
5dGfH1NMOw1vK/OdkaVGRPtSzisH9LiAmTIkxC2XWWNcz8GLKRYq+I+l79rqm1uP5oGBGYv4edrF
/paIwZUXx0f7dW2R1P9tNrkkYySyZEmS9BQ3B/STdOkNCvbSEbQiHPpj2H09M8RUndhIeQYQwrlV
pWW/HFpErSMOf07vojkKZF7b5O5aTQYlpC+i0dHEuFmtVOnbvnhooWfEy0Px0v0H6fEkGEvjMLHq
4fCLIYu0T+xUJfcP1H0Yt6ZjSHpahrVgDkyN0vLNugVg67zQUh2o2VK8xhwq9wvL39axlfzWyrM4
neHr96Xt1pPhlVVgJfKJhMLKCb9vJ4Ig3oDohGbiJo+36FCix71urySebY8SAb2Vyqs7GLS1t6ci
+vYuZ7H6OSRIb0T6Mf1IehX13EE32MJZiMJbCgTb4QHwV+uBhA0oTbsFr8nkHau3nW7pCdW5D1a4
yLrrcuykqXMJjIGhH1LcXHtsQcwzWCT9NmdfRRTOkfcS+8DQQf9I0EZ+cGpmxiNcAZgLbQ4cFX/M
u27dQK6o3OqhVj80n6MIPTngLEOnkiizbrij0Bk0B1MwqmUYJQCZ5oI8zW+rm7UdUDPqnZuqpnU2
2ERqxMJ6yx2vaqttKONl2b5g1DHX7jIlMNkzu+IbMFrLGIlmVZZHxNA+2dnl76vuSlK7Xog1TslX
Ic9RgWswyy7HdIf5fUfWQqs7z+imyzpjpU5LGJ5vejORJqLwcR+vdZVO0feJ3kVE9kIkf7LitGJr
WUtzEGDCKK7A6WAzA+zULVpFaIjqg5A3OisaSESN6PDOpFJXj9+8S+RMTjx3GtQGfTlCiNcJ1YkA
NWo8K3vArFQbpCvebdZKVy5JoQzqFiOPQSwY/8QJ5LWgrSCvXmeNXa3O/0mMwM2rnIDUogQ8bGtO
PYNrOGQ39rmqbHHcVb7oQ9M/JjcgaEvE82ZLVm41pYxsI0zWCFjl0tXAT2vhpgW2oIMvv2XhsijM
fwg6LKPSdgIvIidhUlm5tZLXWTF1o/gwpsObI76im4IOboPN3z2BrLsheZbbLB+qiOrshAHTPeJg
uKmdOJKdngDlSjsqQ8iUSzT+tfh5tzD3KA59naetV1zejZk57zR7v5I+HXY9cJwJHNtTl4ZhTjGC
LKLZD1L1sjlApFcDqlNZMEnFNIdznegRUd5gMsqQLFSzWGBPkq+M+cR6hKy9Ei3qGuZ6IVGjayCF
mhlFJNNhBMrDkmgvUJ16HoRNmbECJMlBODV1qMjzK9PClL4Z12KOx/6uGm7fAhJpfe0baYKmLJyJ
VazzWRl+mYndMo1an5t6KORI2x4/2dHu0doBQt8JfymGEz4KA3qpO3PRsAk9C2rKwikvRl4T19XD
RailuhqiWe6h4VY7XHwEpvhLcnEap7bYcmeb4Pq605scbGK54sUM6R0b951PAz5RVyDgoi6VeLNe
fU+irNutZAJX3eaeIYFgdBATGkOkqfY/VOFqTnJJxNzPCdJHy9sEDjUcAKo6+LsmjlP+9Lv+JSwW
idmKR4Ll80yHWRm767XjibWL9o0kF9rX95dfkn4qoqmvrhdv06UzLw8R4HMxvCsMSzANHOyWdi35
FWcjk7xnNMgri16bxNXvGA3oAgV8qEhHvdx3T2aa3wMqm02NZcsn8bW4s5e/FsmlRHEZ6mRjGOz6
AtuircTugijFBpQ84QacLRYkts+kq2rNxLLrq+9urDl+SjGXSPE6nCbIdISyJAiuFCj6+k5EA3z1
McE56Lhlh9hkFMJkUeR5YCrKIEZnydFBkh2kqjQbpmCNEpiOfD6pzlNFElVr7Q6lvg4YoFE0Ii0g
v7eOpcNgWmgVtAy059YD3jF3/6tAx1wnU5m9Msy8ngagtqBakSYvRCx27XjUpT8NkCwomvLEEkbz
LXq5x3vQodp0I/QGw/jOXpQFgrjJ+p55lUIHUgrmI8lGWjn4TEYJWg46w6L9z3WCDj1Cos2Cv6mE
zs60bw92wPaFuSkQGdnWjAycpgGyJREL+YOn0EWjZjzp1zyCxAlWrXikg2EqMkjmu4BITfiywRYL
Vd48MQwmfgU9WX6wFgsaJG/py2AxMkhdpw1qy4eRFWh4P6zbMaSKjXhTTEYfcT6m1/dSx9dixZ0u
zv/HVvMEAZLS1+mvT4hNzHPqUU2efabLGgUq7q9HwZ6Y5ChaOLaLfS/8VyXUWwk8TFEh7wUitEdr
g0CKlU8TMR8Ccf9rjXMk/6/46hilpLNdJy4Wi3OlVkfUC0iXNkBf3Gfls2fp1aItR70a5kXJdbG/
anRw/CiPdJIwA/7V/r3YLRzDid1dlV7qFlGp6ZCE8pNP5KyvVX+sX0da8cyjG4fsONMIf/i6ReFq
FT4PNOhozoJojnogL17NDAwX/jWCND4kF+/LaXRWlL9jPPotK4k6IXfyfwEYTHAMz1dH5iCJWJsJ
aNQGsVvo5IWFvwwcUHnrZKLxTzPC9oKE78ByB/Ip1s0OEvynvzar3eVnvnHUqvcmBdcfRYZLGXyV
IG6KRELcBeHpOMrOs7isb7NDjppolZzbOIgq0mcdLL13RVGSq1JDEzzopDP8MvG2KNHpEhXzVy1F
Yn1xtMO1D3yoo2Z/YZy7K+NUJrQqu6PRQPN4qJC8NYBThc7r+pENSmT5iMJMEhEKgdhB8e4nwlSk
TodIzJ0UfcLTu76idhkRu0I3XGOOU72cOiSOInRzzemb0EqlP1f2fDkq+qm08G+z7Vk2+/FsuOth
DtWN4DYFxk8G90T7jtwy5ySJIzlTI5lXVNZg7qbcy3Qaj9s2Mzll7fbUmw42GUkgJ/3VaP3SeM2/
Nuq8zW6TAAV6ufM/6Jpu+Ase8yzgOFlr8nrQqtDISOAqPUUSIFQc4cYntpILwxT6c5zEB0N34aY+
e0RoT71P9x3bVprsJUR8DRF3fGkRYHOIVvQlaE2HEYwWGJlEu9BKncCivCaTMsrs8tPFqGxUTZjl
JBBzWccrVgE51CseDC4c/KktRhEcXfysAqtBlN2EZPP7EyHihaNVDpyz6vhuJFk0c6sS+DLk+6lU
O/6qM7oulb8LPv3KzoT1tIUHXsxjkui/bR61C7adhLScfWvJ5b3GSELhHxWwQKlYa4QCJyJDqr06
Xni+iOofEQ0xYITS3xgHs+q/tDDAnL1RnzwhrkNLbOZe5c8x4gb/r8AS0FkXwLDSkreSb2LguUKC
zuAcAZb9vYe4gETS+Ci9X3PkA4cH1EU3T4fU7mLIl0ov+wDCJn9nQopP1X/DNag/Xuzcf43AzpF6
BD7QyjXtMPCEI4C4XupnjaIgHTQW2MuPAvALKMVFkrrNBn6m7Qvg9kzMItXtxfNmdFMFPD0MOA1E
YOcbiPcpKl7W/BrAoa+R3ejmgQMI+ezV9hCGtVwKxHdJZ4r62i+BnfxbXzcG7ONkV7uLhUhs/Hx3
+wvkbTEks/VRC96CMFUMl5UaBWFNGyM0yrCXhCJbfyhyHxIwClNsbxe898q8x/DMtWHOeGkHxvXn
SO0+zB/2qHKVl3oRjxp/EMcWSbz24DgK1TUwUEFoNg5dj2XF/IUZczJoUc8VTaRu/n3llCITB0aX
qLtRXC0hKlByR9EUryM0hTykCD4Vu9AYMpAHB17AVxhHDrJCoImb+3He7YDYV7RSS6JWVaD7DHXk
uSNCNqFWKwBYPSzvkQMfsiwRPVbkeDdAfNHxuyy3wxcpMctl7uZ/LUj5QrWa5fWa/RbQ+8KIk+/D
XaMANd/iSy2NSCNH3e7F1awFl/qy2th8g2reZebc4L1A+pEulLj4oSGkF9aGcebbcVcz568WSejp
SzXrwBfx+PIp2SzIIKXnkC3suy/PlhAxGxjj+F7RqZZRBmNyMwPpBgd/E/3ndbA2HGuCNsJxxgHI
3qtVnSe3rdqm3XMPbGJ/TFTJdG4EAIHE1/FQ11pqxBBy0xFBV/wjufoSm6M4l5xraemN0x5I9xUA
eJOlnfTwdtqmeFRR8UvDJ76myaNR2Km1/qYRGvQkvDQ1BYXVYY896QrI8VeRYJCLQrgpKf0f3GtL
rjtpxL1AmGUQPiiAmb8rpBviFPcSjjhvsTYk8Rsft/KUMVTxjLhBO3DW7g6PE2cACvULqvWm3udX
aB8O00U644n/GRQiduF89S7hoLoQ1fmoKtA+ezNRxlMrMDue3MDAS76fkEAOEqCZBkL7yVU3kEod
jng5LDe5Li6pzWFjwi5ASuYc8GsAyJeeaDahYhpOOpZeK0DpvWShE1sWeiH9/3FkcWT5qtfsKFrN
3yvETrN1n9glvArKOlLlBBGu+5ozVZSOsz4qSRXieQZH0kSeZXiWB/rB00OHyI5be3HKN2oi7aIp
CqGZCdVDO8bqqL3ZP6bAKJyQwxmpUALRqvGRCP9CDcPRd9ZMlymUc395nlQVAmMKPtDjBBQuf461
2i6m3qaj3AyN7ZED0TzjpQGQBCPgEevcucRhZykm1+SdIsRUGL/rcM0Z2+bxccUY+fFq4oNVbm/8
0gZRKG7dI2VmxY5uf7dbjpEnmO49hZ4CbU/yschcyVJI8I+SJg8Q87cxrF9Ai+lmrZAVGXvvOcWp
qPGdd3/Obi0xyVyj7msmn9OPV+FzRJcfNS+Tr98xzjxFNMaAa20hpafniRdT9zdqupOqv5d8mhI9
j/r9pNU9jm0a3N7oOzK4G5/X3ledWOYjU9rutuFZWnYo5PbkAUFR2NdTqN0evI11117XgCPwpMLX
xeD69FevG1eYXxCHo/LKtnZ/XLfhQq8uYWL6UTmlxMWGBpzeoTREcfLX83WFzpgw7bKFimtPmPXQ
dlofzb/VPh5jnupGP3emmBqeGG9YzqC9mvmS1nSKleRcXN67qIA/YP5BrTW8uooms2R2cFnEqhXq
mHtfsIX0H15T8pWjvSIcyu2UniWAm2v5GBkGpNwMXGdWtqBaVsX2Z5WBMMz6LTmlMayqPwJwP/jS
q2SxS/0LCo4yWpjICFJlOi3lXFLmcFV2lRZ0dTDstVxxC7Qvv1BIrxv5wm59l+/HTeIJZtQTqbZ2
qwOPbsDPrWpq3zQN7KLO9CET7cHspat3zBoJOeEAFx6mAI6A5Tno3zZEAqzRdBydUM1ygf8KkhSO
Ad1T3UPl+hg0LsY3B2jsc/3Mhmp7aWXfuL/fqKo2PkRVWjVZLSTxFlgTWjkW2Ec78rY3TwMadg/s
JiaTcO4B1Fh8QBGJzeDKKVXJTeXQq/XrBbUVT+GQThd4PVxoZ5bIKPOfwgo/TCrk4qh3M0rOS05K
ndZJ0k9PoWSgmaFLZBJ0/WTvCSiviytdxeLvLfdaGzt0t5oxfQCb5KZYAmC3Isk3JqAIHq30IGtV
FXkdRYNWFNqN/EUUh4byDj+1loG7I1faJbS6sm2dfk9WLv2GFKS87sWucCAsMSL0YWmSVEjLWgXV
FueJ3GJwgej0QAIWpVJ8NhQEsoHFjTLxwUsGBlu3J+bjADC/J4jeVDwZNMZgkzF01pUQu+VN9sei
cAVABdXL6CVE6wjaEPCJgAtWTMMeQzx6JFGAdLlc4deatb8+yXpNI9HwG+L1sEmAcQ2aU2fczECj
KnarAb7yb77QynT0boEPYqcerz0DannBZL6nhRt/cfIpOzuLhdi5+QEfHZJeCi+PTyY7lUHy44/S
hAY7yrFPY5eFm4PbHv3891BYyyD9UeDwLDgxQY1M8vY1gC9Uw3dHzGZHiuM+eQ+wsd3o+ZohtYLl
R1uo0gHsViZV5WrOX3PBTqbSP++uZtKF9RtOpzc/Ve6xsyiwqkD7DW5I7F32se9ogUj5uylWUDeh
1wgEmRyzACYqE8mFNYOFALU41Ezhh++JHTkxHEjD194iIYvPMOWlRMBbAhgGWlhHyAykQD2Tzvfv
j3SCRhjStzoqdzN1tiFXmNxQ/pMT6iyucXNU5lPdhD6r6KWo8ruKknZlqkhR+Lc2J7pUaOe/qYbF
D/7b1WKvVo9sT9J9NOT6QnW5jsb2MxeUSsAnxIT2bnk/LaY3h0vISSCTGoolkINhptkkLb3/ljN0
5/RIt4qCTYKhOmmhPq8rbrHETamgIN7Sb5zfj7HC3PXOOf0t2Q8VRb2Gn9VtJ95swORfeBgtUn7+
3juR/c9+yv9HCeV437ZMpXqABHq3/9iAlkKYurMHxZCI42AyFuNcgyruSMo+8WPrrWRX4QvFspTN
g0uzaRXi/tFI6W11M/mg9qy2F1E9DDLVn9pzHtD84JeyugwuUu9amNWmDOSa4dAMVtKJsHvrYWv5
bV0828bkGcBY/fGRpD/jM8yA0i+LQ9C4ORyJzmrsZ3+PgHsSU6ETD2JA0hYISCXQrFcdu3OzRLAG
QaFPYSHqyJhw2focGpIR4SqBvzjehD4h2ZxpV4Tv6C+Uv5PytjYo7l+zbJkkiVaB6KofuHRGZTpV
7PVTqVn2MzgfVyXPaJ3p73IflUhqmSs2Fqj2vKhtnT0zhxs2AnObYlhxIDXvwZyHDf1OGLbll0LZ
f0AW/qzQTxR/iWvE2cE9NZ244L4RU2UcQuwsGGL1iQpoF8WLcBuTZ9PqzANXHzc+Jh11bU+X2qsP
D2c78KjliwHD2qdDNM34OxwS9vbJ97cNO2mGF8uQ8lCXppcFW7pB5dR5SbdljhtKUCJCfRP86J5u
TBgRhuU7JVHEhiAc4AzjCi4TfLDcEaziz0q1lhE3z3p4/w1RBeTqo5sSAOjzXXi23aBWFnND9I/E
s1/9g+qMGsdYluuxOHOuin1nHTSaNlFBsCequR72AvspVXTYwVCD9f5SGMjwW4n1nW3OjKBki5Bv
4s2kALmP/+7gfiyth73Jf6xA8Nh24ZpOJ8kDfxhQvGUQP6JU8c+t969JjkCYuUmRCPSC4zoqYvPx
Z8gy4LiqeRif+yTVRt/ridf5GvXkCJ4/qZy4XzeUPmMGJEZTMpX4SExSKGQ9B9CI/wEJiTWyvN9E
jJUKig7+IdUv6XMfJD4RiHZSFLZGf+3kYVaP4AqaTcdyOAoABdMkOqnDBiuFWA4Dyxt7O+12RIsD
FPaD9G6Sm1OfjJIKa67+52iw8aonHABV7McDg2IVdzBrgGDZ/wbkQamra6fNv67eNF2MJaBcNWWt
qS/neen6+6U80qrI0IWf/o5c2Ox0BBWZSZScp3Ws+dxME8jbt+Lpanl4+uaKvlNzpWTxqND2SjNw
6lh26Lt2PQq9JLlbvRZNYdkE3ew7PfhGZLUE7nodcQKGt88n1FFHJMEV+dVKGtemov7OhLgSReXd
oRJoqHjlAUpcwZPNJNK9s/RMf7awxcYKo+mwBbcC7D3F9v9FAsQCZuY5B9PM4HTFjxutgqph3HuG
hcDiklevhkIk2l1AWe5A1f1l7hKnBv4EtZXnsAy7p0qLYh8pXXTaxFcv5w+5d6O+CRERvbHiUMfs
drjaVlDFhGTNzHkrbztmXIXm2hH656VpfzrpvI26i8RARDzOTnrSeaonvuL8TcA8MjTpXtaIyrVb
goJmrzOarBoros+hTtquVBo5gvR9btlIGp6OTWRMITAIrSYsbXD35UXjkrx9oDYMOr8wkb50CS9o
pWJ9XPn36u9Q0g+REPvrJN0IwmvVKxviOg0JzjSpDPyimjmxqV9h9kXIJHVS2puD1eYVQBSF5RtM
csrVzjUQzYBWzAqmqoiuDRY6ebWNaJMDnRuBj4HyadFPhcVYPsffP0HS2TmY25uVt5nxoywxe7P7
uiF1u7bgyexv8m/O2csXpPRYjE3Kwv6lkF5KiGtYYH2p4JEPSXs5EHh8J0bTL9hm0j+4iseIIXSV
a3wcIUWe22GM2FM/PX49ltA5Oph88tI4l/3djfqONOSaH5laf6H3nYubOyUXRWLYPSqz4nySOOqb
J4BabsBCF4CqpxqGrcd+4wAY8PKwyzxuQ8cujMXOjqIA6SRGHCDkGoJOM9VJdyfW5i1dGtDz+eqk
q2pNnNMQP2jdOT8QFXEOnEMPWn6Y1nAVYLTccHq2ZBPSBZ5/aEAlnQIyvYB9fLoJEi7adCBydGqv
3Vqf+7YbTWWSO3AAdTjMLSivgTfTULKtBceTIMpejoHNAhRptBxZKaTeBDtrLOoSFLdU9JhqTvik
p/rSeHylvD2A2vg+PIPxRMlGr4l6PayGwPSRbL4LOz/Q3gHaHIKrhHRqKrpzEtAC8oL1vjS93aFB
5jnIN2j2g9sPXiIOK3WuPhGcmoHrMQLgRK0P57xRC23qMpVoZjuvDJp5S1ugak8+TyobyF/922Pt
KNNfA2EXar/HXtEvATrF8Z377HKOmNXECg5WXziN17R85yXQtMyXmTm0KW8h0Zbxb36LG4RbpQCz
TJjvo78nmAMGA4QEIX78r6jX1SmjZji2LzRJP7gCMaDHWQnRLQcb+jXKgBocd8fHJ7kdBc59aK4z
zG/q7MwRBMT7NwBOc3rHnEGDZPcBNuegdl5mDnb+R2fKvLB2DesFnJHHDHAc0ZHPU7LpTJsaHnND
knmHdtICJ+BHc4nR+SXyVnT4FuhnHJPQZ7iD/yNND1YVsftZYVTQy/ZNB0qGWVdRBqqZzoPyYRxr
TG6Y7wbQRgpnHKRr3E//GiYpJRE3+8P/iDML9C88Vc4Fh3ReIr/ckk+ArDEonpVUAVvbVc37KHgK
3SScuyqTN99macacmCUC/ZOk7TRtDtlN8a0gFN/ZDoY+mVd9PfLQHySwuzDKnncehpNe5q672aUv
BXP3NBa/x6jmS6u0TPxhxReS+83adXf4C7korb0d73R2n3/Qt5TycK7GHObbreYg9By4mK1ZO/O5
owgdwcGKLue5vBfr9cZYk+NUTq6O6T68ny53jepdw0lqMIp7tOouxPT1pEV7OoghU00rWmDpZ6nA
0xrDZX00eky22c4sakVnpcu8qnzrmKZCmKfTyXT+WKcNFGU2PJTzXyRQNta/vvv0hnd3foSWkGGO
5mUO2KUYIxlCPL4KRDwMsaaVbV15/cDCNxD8jBgyfzekYCsm749lgMlSLPBIL1OnLtVu9dXOtpqf
NuWLSaXQsryIAqrzT683SNbcLraAGPypX9n25U3fWuSNIqlGZx0TXGCcJ5CGMHOtCw4BIEpQmxKz
0Xf62b2/3Wupt6lH6NWjSBwye/swap5rYYrbO5goCevM27DEcdhSOPopa3pzpV5F6FCQ07IHbHGe
0jPbD+GJqOYdI7wA4px0DNF3YNWNSO5Ist+v0dESEB/q9Bdm1uzxsFUBpZPh8FqaVbK91Q1yKdDs
Z+oFIM8XIuv0I6ts3nDmw8v+AEpHutLpRA7Iqj2it0zuEytX21fM1Kjerg+mEXy1DqDhJidDs5kX
fo12v3wm7Ks1SIjNZANBihmLfdiRg4YH/gS+I3JqRw+cXA0wnzjLtiE14vBpG4cX7mcbt4mSmxT+
wLcik5w9Xd3Qcow/H21AxnvCQU4gdfKnTQgDy6l22G7kl8XXr+uhGDNVL4HTbCfPoiTm8F4a9T3F
hsxOt6rr3MUa6YwFQDAUvKbEGYggHw9+UoJsrFoI3Pe+pHSdqA8Jv/eekFo+TKUjXlezXcncyCQs
Ab7v8Lrq7f97/NLlyH/4sy11dauy6ADAOVEO5X1EzczE38Xsm7kqA19YxLdOPo1VQ5ibMqst5HAw
koPNZTijhzbJDve7Lu6Xwt9k9qKZvKTqM/MZD3+rtOBDcyZzMccoI4NbJ/Zz+U/ArEV7eycTl44u
uTDLxgpT2CdjrYMqa7VxNghz1l1SxarsauwYdYjjrxyQ6cqNLrGzqRf8ggHIyAdJX0pcfd3iIhlL
TYlgLu99DAjjoJtkg8sAoXn32FzlpfWSgOwXNVcRe3Hg0jHsvmcfQb+J0bdoWHyjF3/a1FltPauh
LWrurDXy4p7z05O8KI4zEE3cbJSIc6GBKxke9tuw9wa8cFR5ljizE52Gi6AkBW+ioQrEFtyAMLVN
YxgEi6DWIifeZLFzgs3PbasvAnf7bXkRCrr+k7fzHBh5BhMXw/eQYbWd5l/tt08qTp4jflhAgqZB
G7Vw2DWDv+CFwi9NtnKHzkAWqHimMjvqRWNwR47eJdsFAinvUKlY7tOHOfnnByEsGy1lRVwnt6AZ
87XsQSkKzjxg8jaSFjdx+IC6Xl+JAJD+Al9f9EBsNl1olwOX7RCFdqURZEJzqwGv6YUhPPS6AzwS
LT8HftNxRCj1OXTnPcIdV5uZ9zDU3xZ+YAFV0HdgmWFqG+eloR5zs4f3uFkk9RMY8rrawemIdC2m
7N20kijMyTLgF56rJNhA7IgXcYOlVYUPZM7ueZlnGVumTokSUbuk3aU8YJQvB24xitIcUg54fxLy
+UVg6GNiL3/hfp+ZHftKsFPR8QwSo41+ITY/dHTn/BEtkOvNTSsHUoOy+kHpI/SsO//RDmYJ8RUg
0g3DmuiaE/x1Gv9VjnEUuAtY15fHqT+jfmpbSgPTRpfUjEIyy9n9DCGbwULXGB63Huj5kzQeLiJs
EGvVzLwNu73ad9FEDCLc0lMj+flALvd4kNdpEePBvqaCzq7T7N/j9jbSpyBtKRZ8S6GrmYXkZS3w
x5342UQLToNv60PSDDrLxgdY99xPtfAQFyB+Ss0vAZMxHZ8uHlukTeSRGx4HI7FnWRkyJLMI8O/4
vys/r8DFhlhQ9cEneKvmNKwYZ5ggCUV4UhVMRm1MrleAheRkU4WQQRyVbttaD9vdxy3+TFrZ1sy3
P1AO5LC7q0Z6OYaTIgZMzaVKdY1QDbB2bwyvlSLXAFob4F3fEFuMms6lsjF8ue0kye1tP1e5m227
A95B7CJ6ArJ2V/SN8i+7W1vrr6kMV1mJkdYRmvj97SpWi+ESZNDOaGgpbHzp/OqpaU41uK6/GVS/
mRxSfFcqA+S1WTjsLVeXsMIuJkDLvBE0CruNQjWU7RIUV9rpbxVKE7FndzsNjBphmeyTG045WLsE
jKL/XWhYUic1NRlKZzCQm2MZgALx6NnlL48h1PMdc0VaZi/V6079i81/ZUo+RNlJeRF93IkyIsiX
LMFSy04neLuNNVDl/QBKxpUvKluJLt5xMkpH3aFs72MlKAfK3rPZfpBKo9L6axiqeIzpe1+aR79w
gNdNVyS99gRMpYtG2lIjwpeuFXLL1p1IbUH+lOVpZRZA4K9lwxAsd+y6oKCv+4sixi4JB8XzMpfF
aItH4RQSQ8HggabQAUGIEyuGsMfRFA9RlFvQ0WsY10+8sPjiAlvSMBkkj5KulpgYWk9EvKFD11sW
knv5WSJDIttcF6UGCdujz6pPDohBMNQmPtQaZ/Afn0QSTu6D9MUaTdhQ0mcIh15zfbaldwOkOzI2
zFKe9lEQBwh2OnTQ4c+5YM4dpTRx7JL3Pjni865XmjwarsJjIU9Ab68O3j2XkiMZnkdXXafl2r5b
+Xca99cDJ1bjb7vrLKm69QpbcWB5XWmP4wy1hd+jELsmPARGHrl9NOpWUEEqq0BqBjX7aUe2sHvp
BhpZtwFNLh8r2uITWbp/nZIdsFU4O1WLb7kLrfRLkrWzm4017bceRlHDyP8RZfZeHflZcUteqd5Y
MOifjmQQPXhrpX1IMLxNvGNttVGe8aD4JhbrYAVSG7vK5qTuv8UpCXHiCcbY+/auGt+90dzjb0BP
MzL9tG7+RBUT2Rqy5cHpm7TtFEo5gO/NlskOJc9l9CTVR+s1waWIpBU8ODr2ItwFyf04RUP2Rolx
KEUoUw/F5owWQJiW4ubndMi8o2HEIsJvrFaCvIWecgG6E8LeRtI6ifKeRB9s1IC9PenZCQFS0K0D
F0mgW+eX8o/aaP30fHhSCkijPJPgr8EdIHku25LfPJZCK8nYW64OJQ0W8jEsZ0tExHS8QnUojZgA
Vhfp0UrdL5KtCEDQYNTbMULw+8mPcE69kODSVEQzVFOfWKLuXaaVJj8eAoQIRKQAV9wS7hoo8lqW
oduhUBKNeN6mCaXi/TzmfYPFavPh7AgJdTae1KVyN86g/zkMx90gxEZoiDYAUCXFJ2FdoJzmIdzG
Y7BqFNi/hhwFHMgMwB1zcc0i4+T2M492jDzmSFyl17DMSsT4lh19kFVJPDJ1kZG8TLMlP1OwPypB
mGcFb8+i6CvxH3UsubXg0VcvqbhYtEBCYInCRsQuytlKieXoWCTt4SHVxJczR4KH4taMgvKBIQwc
0fTKy6CiO7SoYTeoYRaawDNgDk2OQsnhAfs/cCh5BFOVSmdZ3oHxGCrIuCUdF61a7O3b1lYP9oSE
M5Iey0qFbJHKdfqHl7kWMbCNiumyQIJwBrwTBjrrbELgRkwN6JdZ8oGTpFSA0ppHRwtmhbLNhKwY
X5FCmV9EjVHsgqZdEeMh9+PoqZCznVKlBPlWuINfL+6LpNqucdnSe047phGaOB4JOaeVuoyUqEAG
KXPUv2Y4fq058sHvqQ/E+z8GsljFB7NV2Rv1gyMOiwNkc3SUDlWgTOlJGYv4lDzFm0PZN1N1FPRl
D/Rbx+TyKamUoaSPtsgZ9X9Lyu30pBYY2REKqK2T1AQvo40jQtFqo0rRqPN8sUBTN4iOoEu0Jiga
/kD7mcthd4+1oPXVxLekPIGolQnKQ3UoxVYAp65SxAZkQFjIv/L7yCQ9s7KJgPd0T7vCtzFzj74G
EaRuJuXkTNqJNdOn465cRNGt0FYHQSRmNNbs3OV+16RwB20u1UrZXrSIQPkcZhmfBt/iYjYiOzA2
IPZCLxg5UaZQ0wNs2f0yXHLYI3JmG2ZjXw4p20DYWd76TMbbQ4UvJgj0wm9Vwtq/DI3JaNjLGU0b
RpN3AtLOInFCT4YYG8HLXL1lOqCqxcUnXKtv//eTfIBWLXz1IyN2beHHSDLJnyrdN48dPbHrohdz
7Lbs1PHb0Ss4yNxnNAFVVzjjK6WHJp64NMemnoq9xgKlQaVY8brADSs6cIuVcGhHdCBjGSc9IWgb
AlO3Z5vFCTM9gT5krb3XI3xMxoWnJyKXsYy8bekdF0//HvnlS94ToQum/+c/+UFUhWyB6l7mfVlU
89RLN3mmHA7wCZixMSsB/KhFemYBByjCZ8+6h3K9bZ1e2DdXTHQxIoO94RaEFhhdHA87v7v/zUtl
ew0Nr0CvurJ3ckmp8qVPAak67aehgLWS6SxNRgDfziNbxPSDKY6rOYL/+lqbajEKxLhX778pZiCM
wCWiJXnEX2kFFbcDqhXSXZbTv66qN9kE8zrSBvnvkk/4K2h9DLSCHM3VO6shbgj93UYZGMsHxY/I
QajyEQYfntLeDbYUy0PM6kLerokZf+0VqzU5mxG4vpttJkqY4FJTinxFRHKSMuN4hrCvfhd+oJLy
oHLGN5QuzkQ8VH/lKz6QlU//dGHAGfrZzVLAQ5AES9idElvwhlfZpVgMv1UiYYoxsP7UwUbqZ3Ou
CQd/PQhWCc4RsT+ihno5KAFktj13UqOdSwaUSTtfE/fB2TNfEtM4kZVWXwg6UO8FS9Mbr5kW2Y7g
AHpgdTegJCOjEk80khebES/BOiZh0sQIawqGWXpERjBg4guaFNsRF/2H6eIW4WO9hJmwMhdyqDT3
cqy/RefJ/ssmVrAAz0gp5gfTx0CNJ/G0rQkI+Vchfiadb18JEV7P/sBK/ZpkUo9L3lC70GLIP/rp
Cf26s27w+VEcBo0XH3ommCbnZb6vHm2ljezaT7IUW5XfREPPR4gPp72UifaeLR9LW59ad3F5M4Ps
AnedPe77Qgb3sK6k2B4K8xDSqy1EOru6qu3iwHkYpfrlYSzrvmi8fVwslqjumYP5v0rHm+0Zra54
i3GIRsPTSAX5hvpyozv0z11up4gjvWnHdyl3EXDXQHNhv/ozJ0Jy+ccsF9rkYA6UAvuF47/Ixtn0
W68tQDvtACDoLZZtVQtX8PFFbfX6Gfr3V0K4WGir+l9zZpCY7WHVmQs31RcrsQXFsbuS21w3PE5s
0BODZ8N6K2zdmyFU+lymldw1syYqvq68ufy2MLIWQIqawtGWRL+4aObjLXlj1FUUAQadAuMFI/sq
bvUpkuYlJld2m7/HgB2yz3n+s9YoU1Bv2HhOgGmILdPkmxs2Oa1IwPFWWqfEohaLV3M/6s4Hnm0m
iTTcFg5/f9yQ5PC+EnH4w07TPkX7p7wQCqJh0IrYjGQUQpOi51pggVY4SlnXPRAmjahmmFo3T/25
AneLWj2VQJAe8bpxje6/i5wSK7ryTT0lCek5X93+C4JOoxT7SaH/vjQQ4aFIizaVVlApjyDAuDVA
hKHv7GIOLs66mBF+eWI1rMxcXsGyLQQtC0DsiqtVFMeEN8sJRESJxRXe56jg6kNwIX2KKAabkedB
0gdt4tg2vxCV5dSPjx4E7HE9KhdM1f1mgbyEfqOvgh4RcXXTTyq+ynQAmMgfAPPj13D+JfKXtZr5
/hSMKcQTd8Ryc1N10/bRcpnN0fSy1diRUdJugVDecMguKzEcWM1xROzilhlCgldhENmINvoZZvlC
BVBJ2U6L1PGtd4tfrvYKx/oN0LJ0KKoFmBT7G9alajTXCaVv6/kPrWazgNmsPAZR0t4Ji2RAbsQ/
VLJICg8XEu7OslWe7slyfZcuQGkj3QAyKWVKOBB7jBj4ILeDxZPw97jYplhwwuYWxF2xHTq3xsV1
zhK4KmNVXUbDNok/aWLSPSctNaXozCkNPU3uOOtuBiIoChNLditWV0Y4yVsg2Q9bWt6koEvxi4dI
902l5EcrVhzXW0EriJlEJYQ7uaWxdPf+tEb14Isza98jjexomFIR3gF1jEHWm3SsjB3na5cT8Tlv
be6gNNy876n3q5puReNjgYP8fDVhauTo5o/M9o/37WraqZv0+sYIuTcm5MXzzGU9Pa0SzM5UBy20
x4+roTWvC2Kpjl26J0oyXRnUeEXWja6TqHv33dgiwpffXdRWPwe6te66K2j+p4zD3beLUBF6jN0I
kHP9KyGOOvx+kHU/b7S4VofILhbhWLA80+ibFdbg4q9g0FZPxlZs7t3sBOQELh8dHgSJtAU3LvVM
hH16YXPZqJ782jUr56stDOI4n7QPFBa7Gy0bZQ9KKgpAnkDyJgMPa4aRlU2kVPqVg8P6bSu6muAL
2+N6yXOZ47TdWM09Jc480ieQaIetN7hQGmdmbGZcMhrv4qP5AUswkhcHe0my1aAr0hkAhuXcZLSB
K5z8l1Smh90IuLUrVhNNEcLbpBvOhREDSMLaFYhL3gmHu0FzBW7dV/NWnFCb34l6Tse8i8flVxRI
N8PxVyllZmEZ+jj/CdxBQ6/AZwbzD6brjt/9LkmY/lti9Sg7zvEY49M4lIeYI3n0gBHUsbCUdcqS
dKFLuORwkmYCQ+j+5qwxdGz86110R8pH/M2l1g6Dh1QKop+lbvfQj1GpqR25iMW/P3uI1RHko0Et
CCMC/Mh0addboPqlC8TOQbIvFoB6XwjgQtbHv3K6X/AcUFrLHdOI46bFHzHANmfhXg63tsKM2jVr
sdT761pQ4BQDli/ueUfkKU6vuxLT8swUgMVkGfTIlpG5p2a6SibhCDUruY7kX0N7YH4NkFGTFDeL
Hlb3xbBWppq9uJ42aXs2uj/nWmOib2mY9Cdt6e/A9SmCFN20nnUZ8vsxtJmA9LJIqUP69Qaqlf+u
HFT8xpaE7aJCca0MIjX8F5IKNcfwaEUwog9sXMbPdNnNosJuBkAdIvdqt4QVJW0vMQ4GCzLm9UXW
CHVRLVBROnJ+2cIcW0qZhBrJD8n99Ec//7npXYBJxy1YFhBwj0pm7pz60j7lS8ThqUBRfT9Afel1
r1e4p/DDPW2o+6jU5hf1/63WX0q7MO7p79V4Ofrq0zpqse+s+D6KSxuhKS2bHVZELZRpJZlVZ4q8
5U0TSVVCnizpj6Z/cjnYfz6k2IlHf9tQ7GPCBbFCJt4LAwkfCPsf3mkkkxpy1VtYciLFoW2nVIAZ
v9zFcyRCojJ4LSe2DrU/tTykFDncdP8FlztxRtmgKTXk/uUU0bzmtA9cQFDg/znun77t3wobqxHK
ikzqhEzfadRmOFgVjgvX0IdQkE4Ddls00a31JAIWp9VHk0NUJ2/icsH9RZr8C3gqqHSyKKTyTeGx
1kjgFSx3njKNsmYcOitkPWRtpRJLCh5EtkmbWBWLej4JtF9qUfDD6UrLzFVmYmAhKGFJlSv77rp2
uFcAeyrY93jWii2VEfx6hmgP2v+dmK22GUCgHOwYg1zxo3iZ0i7wH6sEMWMMJ+p0HWzJeBnSVTRt
FjZ1ROSG/+XmDgNqog12nXhZhqSrI9OpLGfy1D3r75ejurs1JTBHygfEY08GfQt+F9pBYKP3FmyL
05SUODAZUE7LU+0y4lRcrUpdC2/jwXIKz4QlwW+djD3PleRFjNPADPTg52m/ML5qsnjUxOY1NjJQ
DKOjufyHR793VknoSl/gyTCbHaYKn70ef6a1Oh1coGBEIAOJxM4OvyQoYW93KP4+xkuZABrijMT7
R71bzYUoqWJG3JeKOCBGtD5z3OJV8hI9iL2F8FCb4rZTplkRxZdWkvATPz9EzU/OoiofDkmQiHV6
jHJop70g+YgSLrbmacAHOB4kD2byw8o7+PwA5pljqeNQwmgd8WhiAtE9l9xl6mEQFxJmZEbnD74+
otGUih2KFXKkTUb/3xwXu31tbR23OOVbnnNHOSS5oT/SRPxgUntbQosc0rY5d3w2r9uzZmpAAjTP
vD7i9+/JcmDOLO+8DS4jsG/vLoO//UPVtn4301G7iJfuEEqTXQ/KB2L3xB6URbLBxMOUNqRPymR4
B3KyN1tfejtvF61JaR6ELwyQRop2zyKtQT+F81Wkghi0v7oyWo9rbnogZ68HUC+r84o1d/1DqwMf
sgWFFgnlH7MzxZWV63HxyE9ZFsveZa7XS2o2DjdepxwVIBOfE2W2YcaxldXs1nZo75m7TrUi/FSO
pIiufmSLijfe2fQUPWm/jGrx01bX6lw8x7QrXfckQLwBr2wTdqnwILA+nqUyDpWJ0xVk774qY4pf
3YKCGd5IrZkftHFFYgIWvk8L+8hD1Hn4zCVUq5TYcy0E1sldb8B6fv+RFiA/BpqKpxTyfLwuknyX
yOkh2xkeZxxfcYZnAP1nBwchSit3KZ7Yfqne1RKVhoEOR55diflRqCNnhh0Ip9d9emjR9SOsRC8g
7XwEl1Dceeq5YbQkQWLmKTptCYixbaD1C6bb4nDyPhtEBufgUuMsCiJnThE60pR2oaUnkt/B7qC4
AldCjJS3PbwWya5wUQgKAq1dhskLOksue7ChkgG9YvjH7/rym3kni9Ze/cqYt5RbyK2efFI6A2pa
KN6ecMr9Om3SWbVdoWCfq2sjGVNnvPySolTuY16C6UI7Y5K8XMJHAiJON1cLV0+L9dao0DNyuCo7
isMkAvQ+CNrpKa81Yw14XsS/ff5aeQJ7hCupqcP9hA+CyeZRFGy2bzcgRMchHQZVrZAZJ1BW6ntd
tVBCCuhBPNf/hPRGpyDlb/qsBy3kxnMJhVdqCihN1obQ6UM9bfjj1BMibpyDjCcrBk4A9aB+uCSE
YXKYlKCvN8MEQvVVpO20nH7VobF3SNK1txpiIwZ7wInrfr6jADjdV4nKjP2WmH+kPR75c21gzc1z
6HSQohylsJ+LGmwUW8Y7ye/DkdnApcxu56dOHLPsQ5E/uMF6sV3V8czOcIgslBJ4pzpv0pkTmQBh
Mj7F1X+6QdFP11c6MM+c3SbK9HsEO7WAw3Qf0cfDn2sdmhoucRtJYLL2jz2k0ltSD8F6Bslbc0e6
vAvd5pnNRExhQuB/UwOBGrN/lLkYNTEjGGS97E8MamVcRZ0WDxHw1ub5qp55LELx1rVckqiMooaF
Zn1gA0q1bM6SBDbd451GIF0cIiE83N5OwBLvFr8oFa2FZtIqQhMXjOInrpFSJQDZotI06OufI/6p
r8ZlkRg9jw51MGyySCMwmD2zL+ZaMweafNwV5TdtsWcRzFzjRKkBCrisKn9qwkN9edNxyHAZDoQB
a1cMeW25UAvk73p5dsht5pDYF3VvxxJoiwlx8pMqbWfL1wYJiLQIF59qavLrn+sp2CXXPyl9vbA2
PrSdYjVPlLf0wjuKUZRGdnCMJ50wNwQLQ0CMFuB7whIf5IxZFdFZM/rJehg2qXcgNT6EGM7xGsrA
ng6d4TufuYDKqSxdb74TCwyU2ghXI+HNdW+wRISpD247o0qCnbb3zNNRRWlRXSGDBtTSGBPhBY72
dw+f/z1KaiXfvqWPXfSf7+/FvRCJ8PqbpMnW/JC0CYWR7EnxSO8HskCOOrwmwlMv9HdEkMsFeHv8
1oCS2nwA5e7B9qRed2uvFqAkM7l8yBWtfretv8F5VT1fs9a033q4OEZTeaHl4P746X5+FtLadq1o
sLjrTr4Ud7QrhmbT+IAXwbkAM93J+7mFgig6tlAg4LncASuqN2opFIzk3lw2h4iuacFHD2HGnipx
LQhT1Ea9zjOKNqbB7ZrrVCjX1aTMV2rPK3FcuOVmtgLOKEebqH9XkmdgJFBeQ4XANaANasLjwBcY
pffKmjNDSA7pfmDhUA+70qz+hmUYggU4Y6Mak1Zc5qdj1EK2fKZ9EbQ7GChfD/Z9A/H9immPiOJk
/4M00kaFsWzKJv2tikCQmLj0A4eWvFeDf6eeE0VCI4Q1Et5BE6uvBTfp+DAsBrsXfTcK/p3lEW0u
4EcIbWFAQf2NpZKaxuKpqLoTxLOniScvdmUm+wx1v8FvF3BsVmM85mnMS5QnxQtt30iXpQjEPqSR
YejQapN8gg+3R9RvSDEF4diAX+ay4vTffTyhNnr828kqE20hHfKzxtKbfrCSqMEXR2Xcfl+fX3j7
HuLvdKl6menmw34pRQbdGa0DRvjpPN5nbVgAbcPF0OUkaNFb74esFshkNXFNR49TT0lXT2fEzbbS
ANvygbSqHTzXooQha6XX7gYSCGkNmqtFhsTDTXYiayEkZTqbNMHFlvD04ejHxB4JDnMtSUCN+6UT
Ww4lMmmUg6p0gbMJA1CKLYyrzdAZanmR0M9AnhU0QlO8JtYoYs0M7+rbvlYrIrnoXc6na3eVQoKb
IhiJpIQaCZe7KCrJOoYOHpKYnt3jaeC/Yye/xU+ZpXOQyCCoCNG77lSHHQ+++i0TqvAJhJL8gmHE
RsVlKS7+B1sBfx/vSz2xpp5cEU0RGRiYTfqTvOyRd1Lawu66BHkb6UHRAFl/ok3hKYFOCU489pb/
Gs68ImgPiPik3e6uorOSRAZ6Hmx19qHDK8XvFpAS+19/DPAOlHgShOIA28cbo874DyNlchf5i4jh
9uKkoPPR4IsZV6nmsVWb6uJO6vtCMi/4VPLnG9+sdNLZnV0l4FOwo+wFNHclge1LjO3xrK2/W7Ab
qMyTxxX5NtmXAlxN4UoqGF4u6qIw8szR6x2+kPGQEkE7NoekCFYiR2gUUD5Pq5pEFfjXpSVzIdDY
DN+Po48aeExO7PFk8yiBYRBOUVEOlILAGgUJP3TT2OuDD+xl6Lhcm6tkVKe/isplnZbv2U2lYwW5
78yJrK/CZ7yI+GaZe93N4ov3gqqq0+iESCFJ3FEGZLCYxL662jDlcln0OmkY44S8G+UVTa8rhSzc
hXewvNXXPimrkdEjmQJE/xycbcWn0g8vinMVcMOprBxstdINnCo6VWKXV1LoJZb1wniOGXqW+5zv
Tsqavfp62WJvQoHB2CE4EPcGCqG9vuoArTKfopXvb6PKT8+Jud3ExGBYScuEmtKsaUkaOUe8XzVm
gkhNcR6mQUYi6UKy5GVi/hyFgfQVQ0l4c3lF/dSS9rsoFGhy2HvpSEGF/j7tB3mIe8Uf1q6b7iaO
sgJR7XTsY3b/Pxp8Sm5pPwQPsbazx6BR0RSJAwj15nwROas6GY5hUcqFhQrsIsKprkPvH0+nZRRV
qU8QQA5Xvi2niziQb5KWVGX7Jqztq+uEIn4xdOyRFbuhKdpmy6djxW9JmIxEDpqIDUW/xjPSQXzO
eWfKMaatCYGqVQ3CCJWzUc94rb1C3eFlEjpZZzgPiqrHYzf+Q6mTCMr0/PEDpCFQ66obCt8kB67d
QjON9EJwbX8TX7XhRhaj9i46u/v5G4CMSfflp5S56sLJSuGhLBUGUIDMaL9GC//gr/VIVxh2UPYU
fk7Or4NCiVKRKB0BbxkeTNGIJUZj/lVtjpOkyI6srQvdvtFe8DUcF1RRyQt0asR0RrUB8RHRNi0C
H7vsapDS1quilQ2eS4jaRv37PFVRv8gjriOuuCuMLbaWcxq7iST94R29l0dv8eH2lTSNdPrSOjhZ
LoqRbiq66LxgzB1ZrM90VKk/9kDi0OwQaI3+q9O4CSWL85/BwNpBUSEv0DKV59keoC7bIqhZ0THL
I1EdWdtbu8ghvHALgkUWfEq2Lw2oojnipbx80ynzRjmJd5GAEs2IzfbsnOAhH/gwEPdmq1ArnPU4
WMQv+STsXzWr1BQuCNW0Q7Y2j4prVxFUkpVVELlm+wHWHu7em7MnHtyjeUFvpgrqn2aTj8LKD5Aw
9YI9USQkhU6m7EvhTi3uY9OOJu/tS7dysyjqM7Sa+V6tjl0LjhlfVBW0PYXx3iOgi+v7zdAIF+43
uM4vDZMGGhoPpWsE9Aim9SYDSKLAH5Gnd8OFxjfqygKx/VCZNjPl/YhHixgI/kakUmszCpipveXx
ufWR3Q3JiaP01Dzws+kMmPodRT0m7Vu8gpxYcpdHMJC4JtB/aFAaZRq/Q5pidmGhgk6nTJ8ytJXh
WiyvjqaSLeJ1Uig2VV1XqKpR70hGqnoFBhLU5NHUxS0OfbeUAlKGGEriCJ5t5Qe1u4u+drIMTde3
CnsruWzmICaN4i32hxaoy23zE8RtKNmWhNGm4dHG1tFv6MlV1OWQg7fWZr9BLlOBdNj2eHJzV6gW
sV6y055NeY86KCOvti57GnDV8SlzT2K4MjZ1Nay+nEQkbZ1DIDEzHheTSVpUybnoagLhTGmthkyl
DW7EnW09x1YeqAIQsnRuJJqBV9NuoGZCmp0k1kixMTjZTIiAiZis1mky6ChS3YDA39OmzRFFoVpt
Ke5X5cw9/GCIZjJ05Ta+141sWY6WN7k3eeaXs5YttMpJ1ElD4wzLlvS51DS7F4qbn1ICoU57a3SW
gvGKF0CippMjSahlf/1JAFt+jnKTXpN8kqAsk6VxaohVvh/+3FWJDICcibsmkjbbL7Nx5me/xBXB
yg5yvEeB1NyWvDcHD1RIMkoJ27tCivK77X8QscXWo3yr7IfPQAPv3Y4AXaOwzFy0D3el4+tEt+2D
WxW4izzDi7MzhbGXx4IcFAmbDZAOdYPiNgEq46FExpzEh35J5LLk7dNmeP5K2RpoFszcvHoo3miP
wksO5XriBDxEhPCVFpQMRIhpVGD1+vToURyv/5aUbGxPwh6fHcWMx7dj0fEBBRqDbe+C/Ir2sr85
F1vUk7n1xIFu7FVhuxmwdR+EN4SyBNBAXlaVHXW2A7UqxISuQjYSL2rzNxfaHQLQGSBjZqRcY4d/
KD8tnmfobiu7EToCrdqL0TYPM5fp9FTbAaxD3Otrrla9NDR19IyWJvi7TJpa4HlKDHcPa5+oM2Kx
8q6Gt7zZGHWt3llxFZjhoBBlK1W1keh+vTNxMh3Ca6PHdY3HnZrIZQTmCZuW5LnOWhdUYs+5U5eD
x+qWx8qhtRtp28SKIBxQJya0cOmkE8ZUZMNFQj3sfV4fhPtMdflj+s/UBImMr0Siqc3HOrLr4bjB
HqkZxhqbdIMvS5h8g7OniWke4DCJD6WSzWN/lWGfkIKT7tfu/xGPXEDMOpT0GJbAsxkfKfqmwQj6
uS0YFrN4eQDZXFqiVS5yaJ/BxirfC0GQjqjsYOH1fNZKGjIORl+PP8IfDCDP/XYoGTF9IJrARa7F
XmtM99/oJ9BgNjZN1lvap+/VseNUUX83atdTeZpI89XdPP1rVwjyRzNAXXAOLUI5o6GVTpt2KVHS
dLYpSh+QW4ppDWeHOQNgB/ysKo9Oe4q9kwbBwr/ap0MV+HFAVJw15qhxufiCMcLoBP10fhVde3pY
2ZvU6i3k5GGtSZCMaZf575tZwx3DvkQSmR82EMpH9km5tbdLkBkUhymIhIhmoog2zFWuXQUPH8SB
AhoSnCxNcUhujJ3UwU5Xchx1yzfLmFrUALiqXldpCNFbxhrNEnzyV7nSMbTfYu/CaTJsOZCRZyUc
OG3QhNldzxtTOE7pSQxBN3mfzpRohigVtswzuuTof/d2uks8WDRDF07G52ykDdcoDMUu+ZQuqmYw
kUj8jC1dfCiY2RocTvcIxF2c/XuZTPARDxkrXOPiEDpZF0w7gbdJFIcYBVT/VB07X8DVpuUG16D3
kzNysooYhN9SoNqoHER96YHNqlw3D59V8GSvPq0ckstl13nEDi4Y0q4Cxo7yVY5GhK8LNExhFlCv
Fdv3ilXuHewEjLqHU2BTWRPZZOkFqZVwQIGZkWWQOgZQQi5BQokeYqvNqE6XYZOHqxCSArnGkDWi
jogViz5WZ58dW+5cd6PxIEL44Vxb54d7jVKS3N6EkHbK/2aA0Z6BSQt1+GUTUkP6kMOpcy4fyNQZ
dqgoBOQyqokOnVm9i6sIMzMN3EbZdd8AwGOCf+iizYkzAmO2YPOYDdx7UkaWqWTl+QTdcOqEXZIE
9U0Bq9c/SyIcjSz+j83B0L+CaUWjmyx4OE7DSfX2M1GhuRKmJiQ+/RcFBajV9umBiXTlcGT8DvIQ
BM4qg1B9H1tgpGJetGt90qW3BVbJh5+obALQrIMYd4QbtaieOU4t0SNn2xXQ7ArHOOO81//m0vmF
EIklUGBAL964q7NcRStmfzxTvvFmOpE4f+LfBcUJY+WHovx9kDhsjvutip+nB+r99CdjhGqNPbU4
CtRZeZhHvfQQM4o/4fRpdk2RGr8ian8pEEYBFLP/tIXUpj5heJtWTVOeEWMWlqOvYvYVQn58v9iZ
mzrsqzWshwx8FP7ZQu2c+khEIdXG4XS0nso3nCLE2xomk0ZXwYYU+ZJJpa+k/bfOrVpuVuJly9+k
UYeCaVP+TopVoOtAxYdVo+rjQdzCnFwQAJBziU38Rq9HOLcFp3e+vEtELKByt06AS2qm2w17RXhm
SJDYroxrjH+SPfiyb0EMTy45jhzgogKEEkv39iGc4AyFeHb7Wkwr0/9Cb0wwnx4F/QvXbYgDCkr+
MYJx7yvYnq8g9rmQMmS+cQOFDuaCvsfHqOkpxnVhezEsQaE8BiDM/eCTJPt3oSUOhz791cqzHL3N
+/3sFq5X74gsUdLNxyEMKZ5NNzH8Ltcf/06B99WaQMwc91aoqFrYk+Gnl59Ql5EaS7/gFh6q+hK/
CWz3TIpwb9ArrlSc8qckOqcfXGfI+luCSgtsPqucEkadYQbREB5FX+n0lh0EbyLGnjo48oj2bbmT
KXWSbuazjrGC0m+ALUznzlaQTXmOCuaqiKibZpdYW2h0ZOFHUW31zwXiks7H3cRqN95gGrJuXpzg
jOpnh84/xYKijPtMKUq7yhRoDw8UcN/TUDECIgkbHMeQglvXKhWur41hl2bxorePZibQt6Ya42rC
05srAEf0Ix+qayUq8xvs4I3RHc4PbqWCKso7Nb/d72yZ2JwygxDLsF76Ah9unw8yTsX8X/ANDAG9
tf8Hg/mvqr5bNoK7IFERTqX+AYkOd1M/lGj53dZZoaxlw+WfyYKHzEf84bhgOoa5sPsIS+IuxG1v
25bhsWOp6JWgB/JH93KDp9BQ+L94TnWGRn1bsS1dHCPXeDRn55oqAsCzbttDDxN1DgREG39NfqjS
CDzHuQhhx36SNegB4NTfj88Ip8MM0CuWIQ2mODL9M5Xq0zKBYTtJSid8Wl/11509rgoPmq95TUIL
bNpS+XHjj5SrWURWc8go0W3Yc71z+Nv/PYBN96D9vZQMNNmut1LSJhrSPDUuGfl24TGTlzQ6c16w
lq2RslzfT6HMaprTjpUuKYpAGRYcdvuaTnvbdxxpcW8H58KuULnX3m+xsm0tQ3ubkdI84I6Q7c+f
W3rAuNn/yVCuh1SVvofLxuDlhcLsICi4kdrL7fRXfNIl/8LbCPGjrm6XtWNsb4zBNKEKOOpwK2AK
4ZD9CiegnMKCP07HPdx9WXqujPyX3JQVFfnwbQoTG9czAe2GuSOA2eHC9+C7yZgP8pzxjzKqAQwK
rBWhQseU18BZnUYZ2Qr9yWKkXzRZzMk9a72+vKE8tjYbEXSqeUuRw2HXEIRcCNrDxF9008KyBKQj
fzNt2s2lh6X5RRbFPgM5TiUUsm2mO+3/EiyjJ6JxGDXJvIOVO6/j94SDRSd/9x6eBXvD9uZis/Ld
LGHBxEBaEOQ0drnrcvATV9GBT4dNmQut8phJjDIjEsY9x4HbcW4eCwoorcfrvt7ER4vaNUmx8l6C
QUZyRWXUvisYhJQxTbK5IU1NSi6G+s1FSGA9tm1DPdQpUDtPrWIv4Wlq1E7QMB5yhQJlmMVt1FsO
NsodiyXqpksANYixKW50Fs9ktLBsn92LazzEL1M3MM64YCiSowDO4n+WpoqZC6wtnIMuV7YLbunC
rCKDZ2GczFv3F7J5M5pw3ffDuJ96xbkzax2zrbggJ+ZgrgCLmCanVBmLJNtwlS8pe6Rop2n8bYZ7
rx4mGFu0frIZN/arN39puhuS1oNc5ge5KLPTvpoI4LkvjOnKRI/h3hlkJhidFkAl4LHpBGG2fksK
tegCE7HWsIIknGbwM+h0mIUJ1f/3yiDIR1n41w9LMs+85h7af0JDTxZ50/EZiX7wlT7wUGQOvt9J
x8r/MYbmGq6FYvcDmW9se3jRHWOH/UoyKU4fp2lx1zX9NWKkL6Sk9CoJwOAkqRlgNABWLTHS+6ki
6B6U1dsmUUqELwc6H6gFhtrNQYV/PxgQUCei/KWo5BOUBWnTZYzPx2fVGlRUWfO8NjF/h8QZGe7S
9tRnwQWh/MvxyleNPeQyUso1+F6VTqnf7s5fHWc346jzxSz/X9EEuwbena9MvYsPEy5T+h+vOwUe
EwpnvAG/s0JZ0OXBFrykDEoQ56etQpjzTazlnJI59XP/ZLHasMjmff4BdOJrZH8bSW6FmTpXsQUC
5ALB51+vuUofhevxCeHhBJO03BoN0Clb40IXe4qPPgoG3MIe72xgE2jsgzyOjKz5gkeEbFFgweNh
GnJeeDJsOoViF4Qj4D3Xo2qRy8zjf3WqzWSrvCFBghS7YQXE9T9P7b3w4soLOn1oeztOYaT0g4Z9
9iWXKv5708Lr9olJ/aXpoHBN+U2bzV7mNFM8EGFHoH0hiCcxEVWmOFxnQqs8WVCaiPC8PTcW9Z+4
6xC361S7st7eBe0MWWxcmAdvjRDIv/c/Ah+MXbD03Cgc8MYag69qZSNf1hoRK+LGC78/zWSkI/Nx
4t6WvPh9S1JMLYmaS+ymkzgpx+itni8gynx5mvsU6hdUfbWhaiuhNiYIgSrWCRA0cFpJTB2DT0H+
2wtnICtdnBZhWAb9mtWbZ1sGuVdocpjSMYPsmx6RkC4V15d+b3T0aKUo0mtNB9G0EPNiPKx2Dkx2
RMq20vz/c6FdCTKDw9DqK//60krXkl9A3TQkU3oF+SBHe+89UduCX3dE+4BcapH8JTebb05RPYs5
AntpjY6ks1nJ0StKH16rt11+oi3Xc+36/xmBDw7cKNrbFJCmBT1ZJbz1+MUVyPrIs4LWtotOWNWq
VOghF6dxsjtzyG/QH2uTbH1S8DkyJl6TuoUoNry4xL9rB23CwM61oqRkBV+8wPE7RqSTNGiegUFN
T6P1IhMli4Wa+sMFN/UQaIa/+a2KIgDtV9igN0RntzNz7mK++0OBmzZerYrj3HuSAP87Bq13tX64
/QKZQhDnNjxxQ827/pr/KBjAfL4IU9CTIjigsbirsSmVKnqdLBKR+FRkVroAkm4V2TsM7aCIGSep
cSVtqKXh5aT5Sv1yzL94+nb0zpqxNCRb1fF5Vm3AZOBCXsPuoYxMQ/3nLumR7eUMRKWUmTgM4c+m
H4wa/4a19jSXbKovgV7jfKCFUJ5QegUv0UDWGUQfipkryruCt464o4tSsmwCf4qmfcvEOv1z+IND
BnXN1XjN8H2w3x3KlkVBjORXtdzMz7IArHIhMs47aVzDcZRz3guZgReY7+nY1DZjwEjx5PX+xida
k4AENg7i9Kq/a7D+sePj3epUmcpyO8KI1h3d8h/Jjb3Sl9R3PWlHFA6oDNh2jAUrNZkgRm/oqVdJ
xMfbj4QAz5O5KUmdyUTz+hp1hvsIjXmEEfOzFmHp73dVJJjCIvqhAXc8+29Y3qyaQXadTBHzYVZW
VAeDypMoCYf0j6Wg4neSmFgjP7WVBBBVVUaJ6kiujUhYxz5U+Q9M9jWVCCm+irTCIz5LUnLCGeNa
qYFCMIaJtkqQaLsLgyni8N/HIMXG1o5ubbdN8en7O89EvWxzPVNxldkoLqxegNL0nCmLIDp+b/Eo
Jr0zCVx/9g8ZC6hGAco44ifBpWObbSNv4kWqkOHWSqaTdkl/4+q4SzoO39wBdLsAsJ8OD7gIXW6z
YwEH5lJyEDormipP8t6mS249qkpBkceMjHHADPq1rlim4bvnJdPmio14TGmihAyuhifhIAKAyjao
9sqmMBQgY4i+hGjtm0aoavFzdLukmrSvh6+KwM7UiCpDyavFhckIg6XZmg1nGpHiveI1FedkoLFn
3NZZ7Fi9Idr0OJld+i53Tat0JB7rMS+DebsEloI96wDRjioTnHW/LbtQnMzGKBPkF2UQOFs+GdiM
svh664E1XCBTATTxpH1XLQ3ZXtVKmB3oRYw3s/8xO56LjDF9/JhZVPRb1XRIRAmpeJh90cZZ2qRl
gXAnjDA8Hfc3V8r5LsRuikplmafE9WkHFLKcYQaDQMhYWs1KY7Dwzxe9tI5v9Pi982JOy+g+oXsY
rnTlAwXKIwUymIKJUHmpqdLGgnZqp/qLUPkaN5djEpfXWwHOT34iUqRTFVrw9DUIq/+GXlPlxFOc
wbHeRTUW8p2H26aToO1ed6KTvIu5YnMHer56KgUvbNvzNZa1HYSGJtfRju8Io0C5WoeeS9u+tW59
1SaB+ZMfj2zhT9uFPyhpLAFBIptIXa2/r1QIDzEgjCIDT27pOBshk76wNpVFyYh+j4t7TF1iWIKl
YSmf0vkw1OVkyntFn78so2WHWVXx+hlkaM8LhVdhH2+9V8OQo8g9qBhllfjp9oH2z5lI977ShgNe
98EfiWoplCN2rPmYTN6c7adj1tII5FtY4uNquYM7qvnp9/o2EVuu7bXpO9+0zq1lJP2MT8gsx7rY
qbAxsGRZS/Nav/2RgnJT4yw8u9LZh6RAaHlzImJLN53FdnwBbyTNGr3VzxKwl4QXVM7bo69jMR0V
Sw91WquYCPYQkZ0KwRgD99Gm6SRme7X7U50mgXKA2PnzfZCWIk9o1Qm+tyzi2kQUkHsimNu6qqSo
L1z7B/gIeP9bMcZhtUu2G5UGAdWeJvVzUuecClNx6iorBzpUVjQh1c06u35NB0mkmuDF5cCG/7sd
KcTe1m5pwjqXjVpMhcmOK3PlfpezsV88yozcrPRDrRXqoJ0zhdmeku0rVwcj9FCMpZVJE+oN3gne
jZOowsTMen/5H+WkVQRiiSWGm9zQejeLpNvX0OsCfrXX9ifS/cRp9zYmVhBTrg3qTbtQmeUUSna2
MasDxbLclO//eWnMBMA4xx+duYexzZte1d+yYNtzffdBrzn8VvCw1NROsJpQDCTDGRsF1g3t8f1H
+ls2OwwfrU8SgFJFiL12jm58B8OxQuoQe121ysBWiOFO+6o0Ji85vgIX/xyOHHeIzeyyuQw1KKTn
/qQg9tRxuZaiHwAg+X82jBDTrI/M/cvGgc4NsnBIGxve12IPO9mZ3Kzd5TIYxTylFkAqJ7H7mrpz
W/tQO32ScVAVGrfF1CyIhEGaAZuKm0M5nS/3sNfu8lzqfDm2w9bkGCyBC8SEXfqtS5mBpN6L8ylZ
O/8u0D29aCPGa/jMvcERuo9z0k/IqEiGb1CEldTrtonjxgk/SRDr4LjYkCxzGoQyhyqBJD4XEKAY
v4ZBDmJ7l+Kvy7T2Ivus51eKyu9sk3DiW8f8f0UJT/PwI5ixZ5YZIE2ypMIC/78pjF25o3TB/hVv
zIo1qOWUvq6f4D1mdVCQ4csBQ9VVlUZ2PzJT3doP8lkhrF1gr3ClEkk4M3WuH+ySKT4o0WuYtNXw
/UVOLf32HC/vF2bSAfCKvT6ixgrja9icxFPV9EUOEMG0z6Z9n/bm6yD+m81wZGFZxt2svAYdjy23
C3yBLRNUWqkteVKReSA/L5ZhzATkQutvs8o2SYObgaySTlsBY1KPhjuhdb0umX8Xc425eiTvjGom
KmD/QBTCCtLa2Y5Jti4pSl2D+mcI+WvxrWSHbxjBqdvB0YlV+aO1ucUgWX3ZPpt+ABmYHcZ/OR5j
cRgSO/1IzBOKEPfFIJvxHlWNetBxJDTImwpbhB6uEp/TBZZvJDaSxJGnhc6zGFgtFOmKH5qxbkpy
Ya1Af2n/7bo/IM36jDeCxAezJoK8jhVFi7YM0eCOg0yxcjUsGkq4af0TA7LQkV5+tyWQHcz8WdBf
pPlXrzJAXNocuJRoOrvmQrzC6t85HPBmCAlv3/vYkouFKi0z4L5/wtPCEP8q2eOvOpwAZQIO2CNB
AmFlaqnKKprXzxPcddcjadKjSOd62affjKYgOurxBLrM7P3E5Fh9qWzX1bOiCHMoRk7afzAt/Com
L5Y64N9BzDxxQXCAQ7yXt6h+N4BUCU4Ru4eQZP+SqBGjzdytmI1Rs7OAWNmkF+/MAbESu9bA0zsL
5+Eni/73ELxsr5/+qUQweKoWoLTfFESrPUEqv+cgnf+t/oaD/qPEXXHL2DfJ544Mf/4TqfuJcr81
yFl33TVblIz+h20AwDQeXzPZ6eidzulErO7qKcX7GQ/RgklFzQD31Gqkek43HB25QS4+7EDJchdW
CtZrjgcYDU5emDmOBlYNSBcx6fyDS7R0GFH5VeuD5341ZUMBo+nF2zG2dKW4wI4ZRPIOeTS8gfBz
jb8r6oxTyOa1m+qbvFx/jz0Vf90u8QALJZ4VTYRJnNTq95MSauO01CZ9wB6dsilOpzFrQsGGc4Bx
qOH6+8QOJbcrrPo+3XEBjhTthSFiR2tywktqp17an8p4cHaeEGYPF9CPW+lvMA/gOvX+w4Rwlld1
ZA+N1M5mlezyal+kfcAcr1geZFCheOLH1QbOyaqY1U2GiUuJbav4wSLaGgEIN/r1LCTCCbDnGyzx
jXdcHNzNUJEWbHFUtdAz0tQTNds3qZBd7MmxyoLcbuctxsfJjuKS6C4kC3odxjcusvCFVau5ofFo
WBzwsa8+I1IUd3DeV+ovTc8CqcJIPtm8Z4yYlqQDXCZF9RW7jzyHNKS9hsiNOA0xep6fJ00RBclo
FOn5FyydInl2Pwcvzchfts38+65UM20aw96NDwV0AIna49JJSrbauZBuVgBc/RO1n+a2LiC9LQZa
KinQ8SqO1EXm56c1BYFSoyEVxfoQ+tm0kTSelW/B2DFEoMW6ueq3I+D/1ar3sgfmPycqHe/zhyes
Wg2TlWGUEAO14as88KAfoOvg4JHd8a88A4Z/MuzmIlQHM5UpwqooYSibNIfuty3OTLXJ2fsD0tgz
nGsZBY4m2yOnLfJtUnn9QJeygRGgI5IYHK/ofuML+T0OJ07s6hSNpUB/Ce2+CgJn+1FMkOZV5zwc
cpdKEbmhNnGstvj2y19TaMDquwPRaT74ncQ/qhCAb+HFc0rxy1LOVLhFC6A7Hx3XWrEHQAGW4vih
ZjshfICYNN1UomCxPPEp/HXjY0k4v6dl1RF+ysJBf0M3V1da7SoCXpjP+3kx02FrlgMW/6NjIH9Q
h98BHzv2GeEKLmErwWJgMfA0K4p/BKbQeTKzY228GRZ+juOFpCoXhxk71J+ipPLcvWSy2+ilLl03
bJ28XVW1IHW23goab6QfCahisZ/RCW82E2NUYjp8mVjsR5A5UhF362yUSm+PbcctKH4gCfnWNixi
XYjXhRYMglAxf/1uB/MtMh7U4Wg9rsmByWvaMtU+Am752JJNrkL/lQOs1QDX5bsOHRM+6kjapLnc
ixeg0wrTt6sfq5APlSGuc2TOgLEDRWS+WpAmBEOkS6CLtJ+OEUYh6EDfyobMuqPVNpZFIUSfA7fg
XuYKxocGVWu3VlbGlTykL89p8t2qfks+ByjY5bersz24Z7krS/31AWUFF9AJvOOgREUUnxMNaDDx
GD7UzwyvKX8qSq6x9vgk+B/pBEvrxkJh+PRfA8ipjiikckp0hULRumzY+qTwgF+95n6G/j8vAmBb
8c4I1QNtuxFTrwfo3kcI9U7JvRyOSJceR+yXqj0NplCwX8XXBOR2HmyqchrfxQsg25iGc7MB/J/T
IR+kOfUCO6BecdNSAsGHnfZxeP2RD4UJuBO916hC4+O0lTnKxQtyA3+vDErWdKlLZy1F3DnFQBLs
zCc/Qybu2TAsE/3dcP+Hm7n96HFm/5Stomctzp+iw8oI+Sb1BzlkGbDUb/8/Y0rEpG42yqHhwW+2
138ZwkttoEmkOD+Xn8EmLYnUaIbKGiqo0Tfu3mGXfD/lPTwHQIVuQ4U0irXriFTTyzP3N90U7CeL
8+LRNzPdRHIMRxXyUCyfPlyAUfqWvl+v8Oz5IUnBcfgwMC0f1oX3Oak8qy6Z468KvoH75D5N/zRN
hTYbMVGgpteiy957Lh8VUhmtLuYJOYkxue64wuZiKCdRq9yX5oXICvuWCuUCctrUvHH6DssYoo6R
xXtL+DF6nWKSbuIiXFWUSxRkVYUm4Q9r/DnQfm3R7EGCmvtGwADlh3JUIX64T4giNyHFDR5cWb1+
YXSE/d8lWfZtxp8F/h9STbbEYT9CdDwmBO+iZsPMo1pmiRw7/sjVQvQtqa8UZPIhXMeqp9I2P+Rc
O8m79MCUV5TMEPU6DB05F1KZIGEv75f1T2fbZGGhrVBaHSurW8Q4q4vz06FNuE7O8Wboz1VRdVKt
nZVkFu7IRYTpa65gafN4V+vP8bksLveTVhPAhU1Itp6lpGT2oyxyhEPAzGn8TKjaiueLGgRVTeMM
XQyDJ7jz5BvUzKIZcZIGl5cpdMaTSV+ZwtaNUwTIWMgtfCyMP/7h9OM7xTwN6c1oANo/3ysYkZJ7
qfaHJ02G1iA0ryYTnUuodc80XsmxUU0IgvQrCMhkqNYtb6Fj+hZaC2u7wdESuMZmPzWs2pygT9cp
KbC8gKcOdkrOZlHkUjXgoqChfSrXAs0suiclfp6B4TnN+JKJvrwqNXCGl1VCxf8fhNS58kEb+yD2
aAl8rFx4WyO9CnEWLhMSAeVTy51V5H3QxzHSXo2FD4HYhC9VCudBx7LueA3Ta7xu+lPqp6nm6TWH
u6WQIRBf1PvvsHjw3CrtRO61/uoFSrIhcSb42QO8b7a2L8NXy9v5ADt8VqRJ26tFQTBvsB1fbZ7P
5iripKs5q0rHjWf+JoYA+MSuxtxJ+1IY9m4XGPWiKMuRWLOK0WRwNLfn+wuXMhkVX898NQfapRwv
MvZTjBh5mLMPMtM1ITIe+yJTMu5NkoG8P7SUVWRi+3m8cEEvQBUv9d+I4TUP1K9wOdSb7QG9eQu7
vAnQgzryrSEE8ui7N4kp2NICD/ETgTqLB9jGMKh19AwXk3A1fxekVZDknb7ulSWbq2bjn6VM0Yo+
X7JC1Vap8dSBVfale8eqFvCwMcZFT2K5qg6E8Lxw4bvM6xRCy5cX+kI+d9AYTifBKg8KHVLaOLrR
CQ0eQKIRXGUH8xjzr1ldyFRlU5pknVU9h0GvCXaz971e6rwEHW1L1SUb5Oo/v9dBcUtrL3s50t7X
RGWEJzUEQg9KsJq/PC6NSWyjptegTueUDr3RbRDvouErvaKl7JjlemVPme/iGBcT5qZgUUXKxKZu
t754NOvozLp7DNuhNamaU3sL+CrGRiVM6PmN84dLp0N+Fbc5HtgCGRSzsLchJ0lLlSW6PNAsXL5T
kijOAb1q6TGZuPAELLFvLlyuo4jO/EsB5iDYoashCq/fCNgnyIEYooTBTpnMvTUr3f25ca9bbuqc
7oRm7s+zsPXvEIXY0TxZj06DLYwTK9TPxc3BjnmoacukKguxzyObvio3OYEjQyZcP8tSkeUh8LeY
szOiJYvKEbiB8OCFMblTB62CE3tqVKkxCs9a+yAHke/+SplZKTPAklZBo8sAs2XdAKXJNSb+D9A0
W2ezlcGm4pQTuTgyHUvP0WqWyT0WDn/O6kXtTO4eoqN0DFf+TlRf1nPnVtelP9f9iSdPm4QFjvz9
lrkpjJYVpDJ1/ZeRy1PVqXsYEcui5ybibxS4l41eowz0Pqs22HYcvIHfGlSSG5jaqgoTK7NH6GLv
clxd4TKD4v+GZTIczNYhKZ/2AS+9w8E1U6ZpExJiHvH7ARjxLou6o3AIFiUrNjM4hrCYEK+xe4Un
HfJvD96DrAONnqX6ZdY7TAkZCT5w+yM4F1iN3Cpv5wk+Tz9AMlruD5xlfZ9+0A6VRxIoBRI+AoGn
6LCGnFbHBz0K4zcIuNegsn6L+xxP94e+1dzRRnPCN9SvaE+4VSfFu/YvxVgYUJ2X4LHTYmfSieef
UmWBujE2EGRockSysIiqV+HlHqPPDcN8/Fhd8cksKUF4yx0STcmb2zIc6h+m68KqKAw/qU65sa+Q
lQDi11moZOznqqHp6qTVtLIWQEIAkEmQZarZIAMN4EAdBai7IQL1KOrez/yFaWnJzv3bfk21vUev
/btpu42dEECmppQFV6LEm/MCnTnAbgjcEsOL8wXN4Hiy0hjCygYmIYWBbVRSyJVwE+KUxQOlC0O6
1AkcS9hH1ixai0wqDRe6kB5YNb5lJZAJQXLL9d8yNQSB5Yh/vQh+BLuhbrbMT4msM/rI557N57z3
G7dhOmAt5GH39cxTrlTOz15PqhJC0aAwQ8lSaTz9Cc4wSqUx6q7dSLF1cYTFxcnObl06+Fuu3aSw
hFD1Cg0BDgTCY6P2qVCfgigfGhSmd859/GSZYP4kd39MAl+Ov9kRrXaLR7FORt+9JWDBS38iIcKi
mIcypQbUVnt/j2GP/hGtKk+yJGwmCnIbyJh++IZx0phIxEZ8VVAEsamiunihooVxDOmz3PHBgwry
p1fNDn9m56hwgH5pSiA/U963E0grMH0ro4DEMa2Zl14AtKOEqGGEaO273UHTYjXQNosvO2Q/hNYF
+aplmeft1k/tPaRZo6JQEcqP+5oTs7y+y2Spizki59bjyiHiGqCNOlWdvTMxtaJ6v9c1K+zsq/fj
Shyq31c1ZNhnZrVTrcuFxR7byQARhV84FB+Du1Vwj8cvXJPXeBgBAu9K0OtUxTgxzSTh5yOzr38G
MM5YjHU0el0zkbEHu2ov9aMhiWAsANeXFxeo/akx1k64rQSDj2qr4v78c2sUK3I1XSayPGDYYpu0
vz2zmzt0H2y4/fYq9s3eFLKB8Fccvldhre9YWi8o6NMqpPIi0hPn41VUiFIrP20asgFHvVTuAnOX
gM43xcNcbFUIUG5DCRAi5oqu021Sl6N8ccLvUOO+9IhM9gKFbd7v99IRbmFALSvfRd2PiiKrsdHh
kYcaw37+BbP71vLzEqM/D1Q7ChRIvjIpOgTNcSTn4Nm2PjPxxb8QZXZUOUKbcDQoRL2cU8ECfv++
iEDWMssFsEhvVuGt1ke57qUQL+PrnbFFP1eaAYi09rqOCffiNVj25WpfWcXbDy1Gn+5DKGqUvSt8
8i6yRmlh6uzcINRBCcjljRnIr5IXzB5srjBcMYMeeJicaJbstZ7KzNclTrrj5OwTg9AdGETwDCoR
+w5DbFCWO7lOVSgmczykDUhEILCU/6wcaXhIW3Nq0OHsY+TaY7G476ZxZNZw9qyCCA8B+VKrKWW/
CAtNANqU85Ku2E9grESazYdtFlyHoMuFJtWzQYPGfIIvsekI2AGe3b+54BbU1APrh/SezEiph/l/
X3YdR153zhN52RRZh5RgSYW/1mrxkUqAyShS8x7rOO2VQRzPAh9BNh8qX4USmkRXjuwxnEvVB+rv
/iuySX1dOBsYXhjDNyUSH/HsTf2o4khc6AmPSrIqYcUKlsSlppTgcbg/dpZ+J0sqk/uDDBofGHl7
2cpjqXL8cUa2zTIbkFFNG74hqpesRKQSzAuPqSkDN/wnnvc4w4GtMgpIbIlPDYwiGRMqpMUpAC8l
DYY256nDRo8sm68JRtn89bz7/uZDcVhZcwfhwEBfeU3SyjQpfFQPknSbGrbs2vmpBSyQjbXDhR59
izDNZmaRLCF+2PPHC6CWE+QY9so/P273rXMrhqrdcKm7hl3fNgRBrvaPI7YSwXz8YRSC2OGKpNuE
/bfHdQvkRUCr2iOviKgnnsTs17NT3DgXc6AOR6QYrMDiUumdEirE+4RVuu/03sQiGAff/q2XaxQv
yIKlDV/ZC3MxgrzYw6FAe92H6xRjq72c7dFyzgIN5U+W8SBVMKQ30xMvD/1pFL1MCp61ye4CvPmW
W+SRpi3ZDwXfrhu+WOe9p5XGIB00b7QJu8mGEYFLRYT78V/9I1GUDzqrCAGx/nRAl88+l4AIIOhN
2P5LYIker7OcG7UGBTXHopBvvH8wbvPaXW58K8HAanaAvrnred2Dec6fJ/PLH238p8T+EqeBo3+E
lUtFRZhIP8FbjfRLldah3NyNFMuaJeoeZ8TQgtaSlrrr0kgIPJScIwnpl+vzbolbqoJ9Q/edGeXn
ovztQApfjnoAEfh6D233VI/SUkViHhVK0F3zpg/XneXCDpSGGUi50zPIKynborNFIJ9UCB5JKGbW
ADzXPfVBrYwjOvlWRxUjfauUM2bx/jlcWSyUN9nwm4TpdmnmNiME7Hd5xEqqpHS9Ou2fAznCWCIp
Jcz/s0N8SsUq6Yx2oN1imcgXpos/gtJLntc98RP2ivpcBM/zi00/9o9S8Lc6DQZM8hOnSN5RTwNG
oDKjpsV6M3HZvPriV+NVApTL5r15PtdsYvNgXGd5DMvftJfpZOSXglXEPDxsrzvRupIwPc4qd5R+
ky/SZvt6zZmdXyOjtmQwO5sfjtafNg137uLxLznxjLWT9IjNdX5XhKRPjqUdN0gaf8h3gvTL6HZF
iz+U+RQw/SruwhzLa4E/U8JIyWIh0r5Z9IBgSou0tHJ8wCemk3DQqyM1+WrgaaP5in+0fysxSmza
hGjiig07SJKklra/4S7YN0FUkYUQtIV4ydLWdUd6cAKS5BYCwVv9hILxQv2pE7tdu1Hz7oomaEnN
72k2mV7rzMPniQKwTVneaHioOkaestyREQs/NNkwz348IzIqpwLHqZtqAK7B0SEqADW8LxDYHeWz
6sqw5/CUrFeRQ/cxVP/Fo1MInVWhqgYXUuhLIX+3a7qYa8PkQcMtszIC7/s4p5DZtUh2Xp+ahX8D
YE4y/ZBBbpIjTSlxYpKtSHqQzGmrWr3h7yUo5wPWdTSEG7af1NihBTuIKcwmgj16njY9Ch44iV5J
8ca9gFIk0R4w6I2+J/lmPG29T5rMRJ6R1/aBsq+k0sqWmYkzcNjLk2KPfsTEQOyYbuIZh6KuZbMR
Vb3+ybIp530NBWHUFfTVgQhkLBqTlYZXtqeoLDPSCll73KaMpAlOynHI8VlfvmZ4jPo8WIEEbZT7
lUCrcSYE1MMf25KeizkHgDGgFogYHwIxDIGqyULSZ1q6puvZRcHZe/Uiw9uTLDzPJGkVUin9MDGM
oQfIwGy3IVYOhvZwBs2s6/0IU0gIHtupCzWDBCi3Dg/nhDcgQ7dTqrFsHkkXfWv2zNwsZHLrsneJ
fgSIsNJfYwwkN4/RCDth0Kve5g3PT5oVTmHuhN0Jyk1jY7RRylNz6WbDhEV4W/B5CwDktZ0/tRVA
KHeKb4bpOvYTspcjML31h6pxdl3IWh1nH1+XDA91pZQjJ4toYvzlCtbCxd/1Vm5+xD8tvucJiYLJ
HTUV2g3jlBcv9NO+mTS+zB3Xa14O7Ic8959WjXPlwUs3m1HGhrf+Jpq2nu+ZlLv3R2LTJrzS4ejK
AN6oIfdYyexenY8Y4lbbyk5qzI8BshBsapAo/xVKn+peFreovPfsPJXAQDcaqqOLW7JAkfeAzU1b
xNIej8rWI4QzeuyiLSFAQTEHloLg1MFmlXcK+evyxk0uhXkComf6YGEy7DUVm5HLTzPVrO5c/p55
+SvapEL4PwfFya2Jp7L31q8kc27ObywruGIHNa+Irz549A4ogQ0B6WtG//wlGur361OropewDiUJ
UFQ0ODElnr2lltBHM+fc14aR5mY9AnDIMDEmv4+J7h1GmNvtjjC0XQudylLWf9b1DuMKXojwG+C/
HTkF+MddUzyWpx10yR8wjimPMI28tDhdr3GGUcbzXRjeDsh4p/HIluOYTr6sMo8Mv5N8xy+bZiER
fMmfjigikNlYJwqHa2S3xhqfBud4/xLYqjgJ6X5JFVaVk2Yj+8RAIeSnxDO7NEBopWG5/keoeMlH
+HaNTIv35tdIEslYhd5bb8zvpz7VcquZs8EDag/KFhZe59pWhwP/jyUuWlJHakG5yCkBkL7OQklC
t6duT3cf3uaZaoDM7GpNIzmTb/iFDIAVUJ06qGu1qmfrcszyHfzwkvC1nnXE/A2SoqNTRH0nqQBf
gVcmZww9ynUXAaXHENuwAcBzVMXRYNrx4aL516D+pQ2VZunqHigLc8gnk5JFjl3FTEpVVMEd2A8D
6xHPGV6SLef4p7P5Vm3y/qMWCsEwpzCmLCvHHtzR8pshI+eK1Os58lG25D5H/VgD6ugNMmR63D1i
FqoL4sD4XVRJ8tbbgPQBivPXwaHAwYl3uTqDonqDtUP6dX0Cs+9Arl9riiXFtGUICuXaHVcOf2o+
oqeTPyKrpZJbvWKv5kvYQE533eQR996RaI0x1wsqQ9pSWYLfaLOyd5n1aEJ859gOnxkDwTsOjGyT
D9R3fAKwn0bONkR06pYhS8zXvW0PQ/jKRRe8mFdlTg+NESgH3YZYdIKc++b9kBHjuzSSq2lt+fT4
QBeKI6hgtNC0bJ+QhP593XQBAuXD4bcx8JUmcRgj+AS2s7I/7Uc+H5dJAm7iT8A288td6TlskiTy
RwtIeL/c18xU9HnASSRrNTcN5oiTYqJ+Ofv22l1CUaohQ9S6YUCovC4/omUlNK7x44ayixyI2A4G
x+U6CNtu09CYMpKnGx/1P97Py2CTCoeTcjXLeoT0TfmewkguSLeD7ve7Pb9PUr2rJS8KuK9pw9TX
F4A4tIS/8nRoHGZvhU9Oj/NwNJuReU1wMGy7lWZzRkxP+7/g2Nl0t5klCv+tW/OfnDWwtdehkRUc
A8QcmiVvfczwFtF4lU52ASzTLzx8ICUG3UagZqCwhEpOmXcfCYxPhoQJQ8sEzqB0xTap0PwK6woU
mTl9kx5CMTfoa1WFFxAIh1Ri6zi87YYMpGrM4nJ0DO4idYy93iHCmUk/elMnPXmJ6DM3mffqkIOx
ndr1GGlbWwXltiHkmIU5/w4rzqxgIniXRc0AeRPKFw6LQ2Ep+Uvf2U4n9pjfsL1HpRply2Za3OqY
6Dr4VIE70Hc6tadEVAbUOtBnXMNzHTnFODGoLx4N1T4DfXi+MTcIxdcQSjF/SS6Kv/iiAY2B9SJs
rtNArIyWZiJRO9NoABM/WuSkGszLjK1E0RrNZT1kiPyDwH4vuFKKpK6NBtpvKZ4ovWzqqWFZtjwA
sGBWLH/M4wFWk+szFSta1LAFNWXq2b6pE52FzL2dmCsioXVBgS/9Q6odoRGFiqvaDMLL9dvxCwbm
iv8Zk2nvCk3r3pkP8bT8CIElk7vbiIY2Ofwq0Qj5TiPixXGUIY7pg60ISKG3zspRGaikE3LrM7qw
KrtXelBoSaaX9cPD4FxJ1glPjM1ojRNKe/0zToXa+1LHsbepc933QGraSwr0cvLtJgl0AeJbzBdN
5ZrDYut26SUkmRR9JDCo0VKnUOYY93T1X+dJx3C0NPpehc7m24DMW8aDLoCUaAu90dSILsCEgwIE
eIJLC/tXBEegUTlrqwZ0vXjhCSetiBr0fL3BT5bTBQ5AkVTxebcN2lR28HpxXFOTDu9kaOQ9ogXu
b4K+FBzG09r8ZC/HAiNCPo/Rpp92Ie2RBOhfQ+Vqwg/mVCkTUjmFP8HnSNLe5VovUsd9SkNO++iq
Op+rJZejyz7qQW8JkZcdbMgV8z97rKJZJ42OI1024BxBIe/6RHKoy4exlWCoOFdpAc654kV37iYG
HBcgWDX09ej1qZn9fPMA16Zr5r+cZ1xwQOb2LqRetslqpciH9VcrJzGVW+ugrIxN3jCCmdFG3kgO
XSg5EYDOLYR6soYU7rRXnqmKsuK6X09gHKBRYS45h1U2OsWf9YbQlmIvdk0FU8dbUc5iyfg7OgeN
+W825GRqqTUzRnoOCoVK3upP/7lW3Tbvc/UwoAshy/atApWx5IiE8PLRqTMSZHYHaX1HY76/2YWb
CmZBS1V012GzaSiIibpoEwkDeer0SvZklX9/NMCV+Yw1qp4e6Rc0Z2qh164xE1MfmhV+p9M9O48n
uL85cQRzwtsVjMeokzZJLyPv3aGStGENio+4GnGPSo3KY/Ms3OHZsY40U4n9od2wvDEe5qNBEpYs
033BXGQnrRiZUZSpnvCtcfHUmQHtnDAKSBiBEFnDkTFe490xwVQN0D/NuYLD1cgb481XpC0GIW6b
NMmz2VtYfmGpEwtf5onVoi35W/mMIs9qNZ0EaolYktaIgdYbnWCH4DW/qcBTcTlKScx8Zlq3H0ip
fjNnj0ZmH3dLCxUKL5sjm0PlQk8seC3jn/HOEpV9VOpQ++mwV2A4cOWceeR2xnZ4TQW6Hu5S3JqG
QXGTv0ibO4pHxmwcGTZ5XTFj9fOrdNiKJuO1KHKkAjTpBf3LxBxkRYhCqlqM28hgiU/n00mBFYsk
CVqYPNxU/gKgP8dAejssIDL3CVjEZ6TLuF7jmSLLhGN7L4eURkADaVjqcvdAvdd6eu1Ic4clzr1A
1jUdjq232MRvqeU/kWDtzNoMjomkKvC0uax8I2SI8uhlOKinh7WloqeD89QeSInL7PZ6OVLUUK9t
fFJtcO4GrRD974SK1VKFhSYNfOtLDXf4BR2p2CTtjs9K2GabxCpKc+RD6IqA0utY15EtYY+hkYtz
WzVz6pNbmYRxAYMnlBivPyWZdrDKV9GYFqPMvXTTeS6XI67Y/uxvOEVbvtVyverh6ZM/YfNHXKv3
0Odim9040LFM0ANcczCu1lU2vRiUTAze4EmmuBToXNAa2JjHg50u4OsbHcMigjPKBUK8aWdhaF1q
tmLZHy0HDcHK5U/lZe0J2uhFX03MhRSfstG9s854MvUfCc5cHIfqpnL+s/nL8Ql7Sw23/WYfSmXF
SqCrHScccTFDdskJ5jtdPYJzCss8JptnywJW/Gx58UCT1ZwoB5pYUlguIqqRz6Ha5eFB2kJ50Ec+
ns/e3lKMVZLI9JjPL1hqKBSxg3WE4a8jEMCIO0Agn+zAkv+b13TmbdWRQTt0/ehc3V+pBAmI4FVD
hhb5xiHvc4JEfKVLoVwfB25Du3xs4zSZTOTUDq6QkbzkE9og1bPG1wK3wzLGe19Y18POPbwoTNJZ
FeydFD2bW7H04U8pRzvtamd7xcdY/qZmOLDCYUdXx6uV+JQzw5dBlUTxs2dSiCu9p1J9dm/36Dao
mVB8OXrpIm2Uq4s3Pui0P7uIRPVrsAfv4Sa9iBUTelQg4zxMb2KVsU+Q4dFZkohS4TnB9rmCir8v
InBK/1uIo0B0SDhIoRVDdn++G0+iv/CSVEn3F8mrzjJO8jk/ZMFIflS6OHyE2FSRdxrry/qfkhjT
OpXM/HJYel3lVoG6AoVyEo1wAwzSabrbf9lpXzmp5OO+W1F49VygkbAgc+DnbxoVU9HD3eG0USOi
QZeHg4n5gXLGM/jYOzeMx43ej1wlBH3V5loYC81HAaBfOImaSy+NzDCGKxlc0g3cEsvBc39W2yNm
UKjt6b3SQUGTabelKVNHBj/+9qOt0OTlBWS2Jt53S1bfQYF/2S3ee2c47JF6fzRkC+SL99gKgmNd
pEgbJRU3CRq8ELFsiPgBxSbbs200LK6B6/WjguF+CqUW50Q8PDQEYOJEdAnWV2MpMUxgKeEUBoGP
dZhQCg6cAayt6ick58eLyRVhIATIVnLNGpt2sFYZrwh0yg7+7qoRsViDNwNr8V4s53TBh8X0eeY+
7q475jaqTu7ko4ddd2NBVGyEA8ex2koVSUT52XAJKFh0J02QNrxSC4dsLjFqwGxEwhiVZd33pBNK
PYA45GFmZ+7IcVhgfE2uR27SKqF4CnllIsCdxohMsWu/EIQ4iIRImCcgqNCZFwHomERX4fyI1jWA
AgHCP/+V9080mpf+7Fmn9+iyzH9WLmmZkEUfvQo/IG2cMUxCgtSZcWOeEV22gqqk9JwofJmK073H
2YqGm8qNORe6RQM2NN9BcIUQKp9OF53xKoGE9l+EUGDvzzq+29hC9sTsVp1O3hGrcJrTxe9sYpG5
KKKj7+hX2asHCJY/VA0IEjpTyYBMkkkiI+Pj9jsTcdyBjnjFV0r1DwyfYQnfSuRzM96ifd7XDCP+
i1B8gydonEfibrJQYM2B8S6T9d4fRSRh2BaQCwe49y9S6HwUjqnoMcCXAVD4IwdixZICpWBSj899
oVo6bU8SFlIEpQCSXRy44kphQv/uMKqxTOUoaaYxKBMEq8jxqY2y9fSIYPQ1V9Xs/KP4bbWTHee/
1Rp9cLYDTZygvrgpq+S9ES7V6ewMk6lEhxU9vzNneEEEnVk+xLbb2eiW51uEsAUXIOT8uOc6B31E
6vW9yWHECdwtd/GiUnmp0jrwm1w+BjINakR2KDTCcruIxXxh6rhFeOtztpYRl2+3Y+NOw3ck80py
vIQGU0Q9cXuBy9LM7OKJAeMu6Fr7Pp8cWab80LF2nW9sjJASNHsDTIS/pgnwlns167nb4glBO/gX
vjdDdxWbgPVdjtN7x+mpji3SG50G2h/vJi40UnJ1VXTYWxD9eayHwXZHz7Z0+1c1+yqlMcXV3hnh
58N1EBn0cwYbSHMqshhguLMjL4GHKEStVP+2SJhfFcAvqNnH9k6oTRtn8Rno/vFA6+dIw0r8c80Y
G9xdsQ8iwc1DjjNT5a31kzWTqfnLNX/G1xc+3jDTqYvAslPywQyymQS/vPWY+xy3WRvJIEA2+STa
owiqsneNYQHpdQ5lkgn7SMxFhStFAWPA2zgxr4wCpdcjJrB7PZK91Po3gr/6k45qA3QoIQk54LjF
zN4kInyI8L/S03G5H9mNvyl0Vlfi5If2/ZWh5ujT86IxMgIZ9Iev3IgVGQXnG9C9ZKRXFhXY+KPn
iKDxo81FoUv1Icw92nxiaFmuRBNPxXv90jnmnOoykJEP6OCtmPcDC9SDhR78TVdCJ39r243Xkkuf
6j0RMPgmo6UhydhByv0tO3wxQWwg6L6D3XmP7brp/TfLjAxAINass8JPs7H3NV187m1HoGNv6XZ8
QaTrWvPTJCv9OzJKXKDc+nTOZju/KHFRSdLjiohrE5QGS6HkMNKQIok3/id8aAzpaBNX1/7wpuxn
APijwBo1D0W+/mfMZ8yZPlDbNKc3kTkVqEwscVL3ieEjtUIeJsZpEMdYWijoC3sKUFxNsCkEMMf1
TMl3Fbei7XLqVc5wskkavoJNu+u0898zEbxlzPa0YTJ1M6117W5x5u4c6XyXh1PQ9PMOdq9waiDg
RuxND+1518wDDC/bPTGjYl/sbDsadxK4UMNsQxVFnFhgZ0o16HIUxh9c3fOuEChLaSneY8q/wrwH
NbeSWYpr0z5R4E1tjXv13wOmBVrtT16XLe46Zjv3RSfuXRFfCUcoyNyvbDMdOvHwBS8El/2Juv8p
/lg5bUH6OSLZGDSyD+uFEUSQ6UVg8ufTvlcJW9S2Vn1hw5VgkCKcssKhmPNjYAO0Yesh/lsuTgkP
i1FKTnZ8J7bF4ZtWWJmEGWfuNw9lfq84Ni8sjEqpSs2HtxdgLAXWByOBlJkbiLgwzNtDGwDbUCHj
7yjg/pMiXJMTk/VYsodkFMmUAESwGibr2WGnwCij+pL6i69tIRAPY89kD8ZiXzcpCvTLUOfrlapr
TC3/fyU24DQ/sKeXSitWoy2E99990kPVBxqu4MMpc7hGED/bWRHs6j28x8bo4YxX0PW4jt5PV+xL
w+H8JRHoZUX7baD65++5VbQ1tmLxJ2e8hZTxudkGzjm+PUXc68HFs08SfV33Olq3CHcVrFiSyO4G
Ff7BLc7IyKMmO9IXEwXIeoAiuzxtg2t2+Q5wQq/5Iv7vFAOmtUKtXYpfSzjmCqBpM/qRjCPLjVoN
0/sG3huluCfQB5ECLx7K0TEZvx2Trw4v5b/U3fmyTZFAYtAznbsUP2dhOlvsu2zLqIfL6VnXejWP
iz5U273JkRKhvouwpR2TAa0iA31aS7GufyASoQnizd/f/AL099MKkUbRL4CNYeJtDmwXYbBhjk3G
o5KuVKP4IroxRR/TZfVnz23pyXUqXnj8fN2qSfnzHXzaj1VfcOUr2ddRKwVaDzsdPP67+oUHt09p
cQJHCAmRvhmyaY1jjbRENAdey8gyAMcdmEGwhBDPbDZz0iLo0/LHHAYFgom3H38W0ZICt4K24jVV
BdQ8iPIJ+MMy2jsGTazs7ChZjkl5dNeVZ+WC8tEl8NGllfoa0ZtvnpQ5NwRkwpEk2DrK4ZHjevW1
GVKSpQc0iaddcrcXpq8DJaeRZTBvImf4zZpKaVjstnqzMTt2PTiaquow4YXRxf9gh43olT6OvBAx
UX/IlxUTbb1F/lKMyVoKZoslyCH5HiqY9UXaCfhxO1b84T/GZECdZ5wLyJa5/6evs3ipkOpj21TO
cARnpbihq1fZ6jF522dZ2wOY7YhShQrXdCplS5vtK7UX4UyukrowbxnRgbQo5TuzkmRlxNKwNMUn
Tsa6MsPeeSUlAoQ0B2LZOTuyN8BYPHTZzArV0CfZUfcPRxNqb3EJ/U2dB10Pc2PSLXbx3ot9DBPg
oIe2L218BLV14e97T6gOaq1mnIWuKrihM1FFsDA8w+gqDzVlwF88K4nxUxr6a4jNm5Q95fReOajU
X8G8sk1609ApIQBGnxB0iZFd+15EWrzgcuf1sQNE6YvW27U2BvphGMxy2ik6zRgN6jBSe+VE4GAy
dsr56tIeBKfoDEbYtbAAmrkZGckvkoEf9EBrw3MJhDH1eJnDj1FKkv17JR6QadKYXXSKghnIcMqI
OOltDgI/6N5DIjZfZgb4T9mAGxgdF+b/7qlDXBQ+7ieZ6UACqYOVTlfqkkpfKmmOw7u30An5fZt+
8cTrD6TvlXS3lkhUfcfVief/cC6rlE6S7PTce3cMnMej9xCkJhIxfnNNjl5+G/8xako6BgGB3x+v
VpyDvmJEHYuzGUbecemmlydMVLLWySvuRr4XDZRvEvnpXM1NtBPaxoZC/ocLBOYq4XseIP33JbDY
wwrrjKoOuX7Vjotb8HRgWmVoa5iAaojbgkTCmGWqSH8gP38OvZ6tUU6SUTW4oqqb0y3WdcxVpuHR
4Hi8fraFzmlsZAPfD5MOWQ5rNSGEAtmzK5AfPUyH00kHQxduJHHy4C7+reliUjULuWgn3L6WDEzc
8h0LWtvHwJiPnUybBOS+8zHn6ONcPPbx3mdCODthtIE31zPGVjjbCgj7BLYxhqBV3BroGU0s9vqh
Px5fbjIVeOFrWlT9Y3+/yQ4NxaE0lxdvRLFhKuLVAvj6gqX4GrzdZNzWT8bYN5y3cackYVlCuIav
TBI+4bnim5NUU044hGpMRcB3fSJX4cZhQGkzmnJK2cKq20FNAyTcBY3B80NrVaaoTKjek/PG9xKp
Bzi0hZnn+dWlsdyPCIkz4x1AQlUh1Yxj1eio/opCgOQUZzLpGZFB53HjUINOVFcj3RsKBhIveYU1
ThyMgKYbDovMEGq99iswgFDxw4vquu0VuW6sbTR0a+ZKOl9fqkS0Ougi3xQme4hDWH64pgz5206M
lUWbgbVOVJNPCPeZEBQVE5T0rMn0Xe30VUusQddmm8j850bKlJfHbvj7DavJTCLVAu4q7kxmHRVk
u3887j2LvUT3xGlmf63IgS9aNiAnUN/zkZsxPx3wdLwO57o4YTb6gr5TlueXhG+zA2LIF3sNG3Gh
8ByCTd28EitZJyKwM57f0aVz/Uv4DL8WrG/vLgjwsKnei+n+LR/088rv/L9IreZqc8H4QYSp5YbH
pQm7gZceXMnvrCNSArOwq1G86CUgQA9Ts4a2Xsz3Y39AbnyKNr2oF66qj4mVY5D/OuoIqQ5Ew56p
3aSwAGMgWtD2xsJaVUltcN/dWkLTiPHhc91wdElejmBKMs+38wJgaBDYXkSXogacytf0MhDwd/Pf
G8UUktNYWax98nonP2sKVO9Udr4viJ/QogHnhwf+8dHjI3Ei7r7/xFI+yVg7Exgl0xnvM+XmlBPo
+roihmKSUgFVX2lvIFmGRsAAnraCPKZkkD3AX0Iotp+OnvvNajkcNvZRA2Q5MuGO1XjpyIzZKIFx
9tzHY4kSug/M/m6TJKl9SToqz9JSVsu/X00N3FEWzPNVMqguWjrpIc7s5Xv1rMI3Z0GeDUDl0m46
DDojK6S07GZs2iyfLr/n/ICQO52bTxklWNmqz/5/NARTjWK1tyBtsRbYqx/OIxWz24rgYGyS7epo
p61KmhRxLb/92Gbtf4aZplmtNLgyOJ/Nhhrv8u4i3gnt8a929164/Af4qdym/yt3xtn2ehM408WL
lyldNDLhqxMNYWl7mICccxpXjynOY9qjfNY9GwrmeSqISa5plsL3/HqmjZh5pAHzjxyk+CJ+m2Mq
fxJn3WuTHGoJmKIFFbulSNWu/ATxylkLTE/Y/hfTyO7Tbt1SHm+9eTe1jdMuTTfuKFHurGYT1OsU
N/EWpKyxjXWZ+Z4AKKA4OStmeo7BpvxZ0pQQytYOiu11wBTnqlxzvf/bWn/dDNet+x1V3e2MOnwY
ZCvEt6kXZ5OAwQgWDoRL3b5rocpfJfhZXTqfol6VEYTz459KPMRgWSvBugrb4JNL7oAq93WMZP45
t2d5K/kc8cTWfahr06TVSjsOYMNHt8RpXmn52phW0MFnd6zRV8AOnpoHQKl7BZ8X3C2HQc3rsd4K
0gyhBkPartHhEXGGO0zncwILXRjIabnfxXdIZRDuPCUV9UtAIrxQL+2hZ6SLzQgU52YhhfGTjCGK
YsebHBG6uBNduTD9MsSiq1rYLWjLtrU1LZjuo6i6HjnERFgqCGbS5Y3LtLN4ZgktWztFNG1QIc7r
5CZnUzvIrRuvUXF7TMwhQ4THkIEy3zvJDkNyQTtp2cZK8qyOLCfZxnT+WdCYi3jjQeL2SSjemoPF
/nT9DTtHwqn1spY9U/B1n/s2OWVYYhhwfJi1UPJWARP2aAoXJovoXWwTq4UknlL45MT3AmsmlVFI
k7Iqzu1es9+1ZbA7ZDPrIV+OOJkchAgEmpY4wJiHCSaM3CewxVeR3RYdFjQ0S3MPYK5LSwt8QewC
+uOzLZBjhz6w5TunQx6D2WuE0/C93ebPdHunuWB91g2g4NtAgiZZrGFlQFcD0uK83KM1dixojj2C
RMU7Z2PwMkwRRgQpnJw4crl1POZX1jH/W19DgRUPse7we8lHA4NS38h6OTfCAF21L0I93Ihkzfg/
a+322amSyjX6/LQjdFnVrSbanNvf1X5Ye/7DdF3h/R0mlBwfqaAnfu7r6WO+c1XlfPxGunfJ0120
B2DSJdtzT2NtewBH0+TjQxHF5DQUeNOxPbZPZlhnmBUnVnBYccwsj9DrsnoQW67W8JegrTegHBi+
2eqtnA7sJ9D0DadiysF+EqZwHsQIaCO2SITJW8X8v4GrUnKvY5hGKUY7UkrBIvptf6Ze13bs5xw8
23UwqpHl45HHnxd3sGeJqqOtNM381dexFGcynD8zC82iUkSnz0HVWHdMocSiV1XnYQX3KNwJ130u
jU3qRg7nitMhhhmQc6Sg48gf5XMXcTAjq1UrzukYTrY6XsUh5xY+twcahMlLIVGS+kLVECZ5CvGz
dQyA5ABm6x+LCg5NYACqdiHt2Xow65hS1/Ai1QzRJmm+huixoq9K/RuTXzwt6vGCgD3WRl2Tzt+k
F35n29wraiULtuO/U4Xmn+ss1m+xTrRig7nnkeN1vAsYt4Ha+gXWLKtVa37EHiToVwFSCke26sb3
pvfGXckBwcBSQuM51E9selzd7RIFq1LrNLn3brAOBIjRJYePLTDtXXpSQpHCOmbmN1SRP99F0/DZ
DZc4Q+w788FhcV+gc0bPa9vVFufMLen32WH0KUaeESBhMh9lV97PbV3XUooTYEqQokkhFxZttDRp
kK2PXIEa9iovQdL3UtMECm9iOQxLKPRwCaA7VTeor9YitAnb6HoOiN4POR2K6tCIMo4/dPyZ17E4
2xpS4Hy5kKTSVmNeRxrZjFQcSlk8RAl6MLr10RDhvJEum60AnMkMpNzPowj67y6avhf3FGY7bj9J
xu3KT4XgO0QNsOYEhOOc9EjgyOQFu2pc1kHTESS1omKkhzOdJXySaqkonEc6Oe3wRktr4YII4PmY
5aba+vP+llb+NtC/Bcf5AHz3ZzrWYjUrtfmEAwQaWkgkPoy0p2/mPC2Tscv4aWEOrUIBAl3ndGpJ
cvQBDf+zmmHozpxDLhLotTXYNuaYQF4ToMlWrljcKN0XeR+cQwBnPt9eLK9EM3OcVx6WkmJKx5y+
hntVvK96gj+3rpsoCc3D/1yDWlgJklJeNjOFD865bBqdVihoJp6fm5huI8huXniRCVd37kRT8QoA
uyhOJHz1YjsTnXSPgsIGnFJLheU65POMwnvIjKYp8DW6x6ywfWWcv/rb1bmNzU6tvcTgY4fdjOBI
ygdN3h/kUZArSqp4wV2mzg61JGvNtVriEu3zMWBGJ9C7JgijUWermEwkaHNpRopIZrvGH76TGraS
m08nMarOjSqAdfCEyiAJ/MxK68bR8vMbCP/90ywIjYwAHXp+SPeNrDHoJ+KPAHA2ktpsDHyrybcc
p5tq11Bi5EolD+tVDB1vh4zyorSV1mRTT+WloW1RFWRVROgIATNfHYbotorQareEkSHxjueLccI8
wiy+/hfbcIBZmLyLhS7Lr4gA+IPWsUIX4E8iMC2DOA/UkUsWPpmGG8OrkHWLO7h/u5B9bVzld4wU
GI6OOOkVfvCLrTEKslyfcfU9smG8ZfpaLU2iqaO1nT4HKK0Y7n36HvvxzGXHZTRWlSA/24UIeqxc
qCC6uiXQH7ZtIu38qySrboz5wfkxnM/SXnAMTJ/asRPOWmSBP+p4ESMAA4IAo3dHWqxrqV0EBydR
ssdN2hfqV59890yqf6lRTA/4+TcUUm/FayBcCfyY3HUDMJJoatsSEuOLeBG2TQzjj78wx4PlG5yq
9NOk8idXlKvI7cAPmN5jNz6m3Lr+j+ZMHrzuMmNS5Wq2kn5HneDN6L/tNIA+yNquv500XIAeRrTg
6vaQeZABv6fWNXcCNaBG0uPxPNMRg1wc1oOC1YTdokkSvAilWYj2LJsRTbuhLu2gmr1kIRlCJYkn
rlq+BFGTKJjvJv9ki4LcvqOFG2aZb5lwTg8bDlj8VBBh8VX3Bqp9sC5Dq5hOM+bhfr2RMgRh79b5
7QfgyoIYgjgXvr+9r7a2jyzVkGQEcrBik9iwMkZgiAT4leDhrPOJY5uoB0paA5nmbrouMZT+BsPW
hnQ3KpBDYdVQXgsloKsnGzvrLATEqC8iDuMwLFncTei9mpXPb2Y7SaTu3FJKEDdrcDlLezVG2Lyp
5cL5EnLA3d6h2pyYphVBXD76jL6Vso7cDS0s69uGW4sIgBj+uw8Euuhf//6Ff/0vdFA3NN9OChaU
TxQqlE5aQAH/kDS6Yn8oQsOmIohacx0Bg+UBzk/M48RO9u7HPdhos4hw36dxaesVVr0HqRwS1oC/
jQ8VaBOnNVWvXb7p1s85KXqVrsDnXyC94AJgGaXDOtsQyAFoOAnN7yHi4O6XXNjQL8ADALHMVQzw
kdx8Hp+RtBrhnJocBHs71jFvv+KF2u2Bu+03UAOiOfrK4f/iugiWz9fO7pCjcnrOOtrbdvh1dhL0
j7Oy+hGJTrtmuQY8m6quSPtnRo/RMWF7JH/Morz735h6bs8+bZyPUof/Pn8g8FyPRdvSxbny+hTx
AAob3+14B8JM8lSvIX9lDxszdU9DlMpcgxyGW5nK9z1NpSdC2rvWR1lWeFYqjZ8GKuXaKp33X9IH
ijLkvWkjjFrBuQCl0qeDJJaM+eIBBJziLRq/PiLJV2QUm5k9OgtDT/raAy63SdCDpXctfa5AaeoL
IYECB0S2mVgjLnmg6faiw5KoCY1rHib/bcpvU6B+u2I0w2NXxmFWo/HH8wthTfb156OQb86uaq1x
Q5uDQvdSoFVVhXu4EdzNYId/8WQSoGpKmdjDmkzUe/9NK4Y/jnJeZZeL0dWhKssTEGoxjpVQ82Pa
WaU6EK6BSDuY9jvsxWDVJWBh/rciXOmUfDw/d84ZVmxmxRt0Cd8vChfq8LYyrNS3poI9tscs0IE4
HACmHvjIr3sw4Bzfnr+2FuADdTFmEF2/zYQccD+kl/zJ7OSwQclADurio3NUwqodtgVG/30BftIH
MDRHXdWg50VxllfHdZjq7+2IaXhr1P1MQ1d69ddtQMJvNdqNMxNegv/2JjnKiZ0C8GTRph+xj69c
wrEXwLYRdPhhoh6EaAM94vvDBGRGKY5yfEa6onxhtV1jcGH4gyivZVIpAKixngG2Tzn4wvPZYniI
D4vxrQidrOUQDYaHCyDj4/v+I90fVHrZXGKUXf05o4EurNPWW7ka/QNzJJnRpOH4gTQjx6jjdtcY
XPtnLy3vCSyrKqJV68Hh7uSlyLswdBWhoKHrxaNKDF4RhmtLVuDm0I5Q7HLz0F044OhkmlfA8sF8
IBfCK1neQX0neCQFAr80oSqSnsd7st/0phC2iI0nzhNmZyAtNdcvwRKF3FHdB3/brD5O6cyzPlkM
pC3z0Wk9Rr+X7vq+5eoRIMAbOQnsa2lzbEYU1feRsK1WlOBa6NJqo1NFhBoXhTm1jlz6Humqz3tA
vF7UDF4EjqBIOPwzCQAKRv7zplaX7Lzgi+jWYgb+SljJ37Z4xlyef2D/zy32hzeDG09SjBoW33MH
S5tgDSMiiglIPxrg20P01kEA7N4lL51ugIrUn43U/0A2MHIWMcOL0OFAEgE5Ryfnw6BwFq87aPSi
s049GVbLkadp1s8Ff25kMJjgl3zn8xQCfAkECt10I9q5PTuSoiXhNrsaVzmsOcdiWvKfT78yG7N3
c6OuFdTcOCFqnpuSihcdTyFjF+VQjd9+Qoi29bOEP5Ogya4aHFTBzduVaD+twQHn5gpawReN3H+v
2J6B+Rc6Zx2q6Jj466ytJZ+iKG55V243z/uRUwVPR9niktdPQcXq1XG3Mx7tpXna0E86gbDuLbT6
VGCZfP/QQSlK/w4N3WYah8kKjsDS9bI1banWoQWpAcwOSrW46iSmHztKvEtRoLWE/ganICNTvqfH
mKcPCKxRg3jAA44OTEbbm2bMTSHesyZbv9EViFpTBXyDXFKAyZosGQHrLVulxPfln7nTTTr5kKsO
HkGsfXZ/VEXv+4MHZz7xz0VbxouFm6D5B01OYzHFr2fo3x7rNj1sC9YPI6JcrCXS+g/gaBL052aY
btjXL2wVik49Oufm+Lkr5xkGsZ3mMn3TOcE78CbndI13Kbrx/oJcitmSHk1VBW5Z53G4gF4nrTUP
7Mvw8XnsCSdTR1B9B+Ou7QEfMC8upIlVjGM5Ribn8sL3AYxmXBDwsjZ4oqyCjfhAFFpwevLlf72e
nW1/RjjFGu9Pt0o5bWXaF2Eu7DqV/gYt29wow9SGonxugkCR16DGeKG+JRBqd7+61fI5H9EGmlCE
TP8qi2395dIeEQ62Ff5QOpdQGOvQvawu/7Ix2yRl1Id1gF72ayD+TAQxNP3Jy79/SfUEiJxYYDIJ
t3ADDCFmwWUt50i3K8dpfsQZq5v58WfWKZNqUjDr6LhMLbYZOiEPkGgsZ0je9iaYY+6JpkIEVOxX
gQJ75GT4gkgYD3leDq66ytt7/4wg4j8CJs9R1xndJ6JbbTOTQdXEmzJlOH7uwhpXUSJTX2uqxq8A
u+oD+tQm7dmpBDZvU/xcuTTvbZgzRYOb8X2lck0Z/ljkXwavnbG+5sC28SsWjCcLPd8fC7EkZWcg
RiC8isWtXI3FKT+sIGcFOTdgCfIjTdJeD3Q/4nUETyt42gFXdmR9tcpQbb2lan0t9X0TTdAEKgtZ
pTAyzDVM19tfpKLMk54QG1Xev3if7gt3jTlW3UkFAwicMpp70AL3M3BjM89WjQMFzcCjmBT3C/jC
7Kztq1hSMb8OAiaXknhPuA1T9ogbk7A6YOyLscAvyGDfb72/u9eUG+SjsbmPM9MBprHcwKKA0MrI
hNo8aFhwxUMfIubb5oUjT7vSiKHTeXagFGcu8qXwRmtxONE/Qgkjt4RrWNXenLbpwTjlmqwM6/+r
IYo5izK+AoHsvkqpIe2QWjW3rq5PTj4O9JF6d/2EfTExzH2sLK4Y1YRAWQf7onyTCnosUeUQHocQ
WUvVhkL5EalikwwwGzdhxP/c+WJ4Eq/2fpaxUws57N50Zq42THHL34bjlM43Jxvl19HNCfTsoPyC
2QjvregO29TuhE5qdQtJcJvemNXzUzjkfZutuBDJagswqvh2ruodrxFGXXl9ihCVcwqa04/2an2n
aptqwu3y+hi1SfD8RLgMo95mqZiBx0JirTAZTKBKN8DUYB4nO8Z+C1MvJhBEXSF1D60Nep9vHbhG
pXAkY5fspEWFCbyGoJv3+XDYCxgpKOQKE7JiWYIXKow4/FACYb0gy2bggVY7fPL8ur3tW6VCgYCn
2cTbD6X9WhAKXYVqZx5S1yFxJA/rsOYN+j8bEBpWd7MM5LTz5hJBFKmk3syR1JCZGdwj9uxgNRPF
6sA+gXXB7T8X5Gi1t8ar5cVqOpgQY8DWDzdBlbysCuU6rsEQ/Rp9icBCJGczWfwEpS16oiqTTj0I
oYOfgtB/ErGAKt9LowgEQ1fXR8Vd9CJvb4n64kvtufvV751gIf89Gzx+SmwrjHRXq2J3UkcxqU9O
1nuXqDyjZDlTfsby/0A/Ujyd8toOo/AZyR293spdTCi3nQF9BaKWeXBovTQnIUjgrWD6wUdz0hSa
Z5w+Q2u0x4BjQzb8wUCQUBqbAR8iZaJxQumZzmRM3nVzk0k/iJmW+EjlVoFLNiVwTLvJ3Xo5Y8MY
g9glOlqucgI/P8F5+DkGl8Mv/uIb246l7dzewsLeexN6811PePcNmuEGGj9QH3QKvBA8SrV7uNkb
uO7alz29lmlnuNePxHNb/djlUlSpXtjT1vLQ1+kWz/NH0+wlzfg8H6Bcf4EAOfj+xlw+Q+PZDqW/
29ZiNZnCG+pfpDzfV4Zi+zK5TEbr8ete0zA3G2koDfwrHwFDwDt4g2FwKFwUSlsC1XWA6nkwqpFL
T1fHdiuRpDDMB/6y90ltshQo+QoOR0vElTIgNXct4AK2DRYtSQCTLcylBh+aCXM5gZzGCAQrl4O9
+OGRjWq2i3tqn+8Ib/ur9GSNNsVDuS4O0Api6oW61MJjHfgA6Q0U1/GDieHw16/ncdcyOAOAHZyl
PWTLd63wakiZovtAnByMXd3xJ37qetko9Cpq+F14f2HsowCM5dK7+QFRu8r4FWhdDin8CDpJRdv4
4z9R9ZCD14amnYqQ8VpX1EXKfKPU9YrNvnZF504+q19/ulyWW4vpRUMdIlWHO9MhCYwv+fyh2+Gx
2mHxcMV+V+QbFa4L0Jrx6mmyBsrFHUYMktyM63GbKFYrQF0ptowmLQnvuVMTw0z+l/8Y6TGWDKRi
zxvzIm1nsBK5kbApCV5nvlCjM7eFMSkyGVBzUe7OmOpjdYUZ6s8bejMuM1i0jMZlBAEXz8IqGdGi
uwNK+v4ho4jLRUy1rteLZRuQn5ejvFgRknt0mBncPeGkz48ohQHRnTHzVN8v9Ah/jsMLzoeh2mRV
0W62se7QNFms694ieCHOsa+EvGtRQVhQqALz4OPVaH/jITCkiwDF/Dx1504ENkadfI4505sAVLEv
Fzt9h/T/Hbhw3muDjL7CZFiSCw5lLhTI3HglxxEXEEXlIVvt8uEgRQWeLRENe6DFwBVrvUv1sdii
KXewkDwdOKuZQ0UTEm81OEEbQnWpGdr1i3aJTXH8mnYQpZfD6UrhnWgKCVYL4eY+5qbKBdJC6+za
h5URo0N3Uu/kH4YnkszJU2DDmenyid3Yih+Ganmkp7f/v6H/lG51SpGF8GvPLxIXfh8UE6Dkrbsp
H8gnVwkuGCu8tlKLjQtC5AlD7lPBNIn2sKRGoEmW9HDg6Wl8PslhGgQqJgrjEJrVriTovjG04ekg
FlS8qF0e34+yVGgGXVEWcjJQ1zfZL+nAAp3YWJYv1UYfMsIO4sQF/XAEJaTtTg5pAAx6LMDJs645
HKoNTNI/136CfHi17G5gNgwGUfnNJWK2a//WK1M9hs6kX94+xO2vgbTr5KXGG4ex4gKU3eL/iQc8
h367WaA+I3I65ouh7AJ8SUS9ntsLzAZ0diJdxZby1FJuDyYgTEWAoho35I/OqnMZg22sf2CMcpmq
kuUgkPO8MNCPOj9IhHNMQ+C8qFsgIjFqCcSxx4s4ZgXhMLRfArVnOhkfGL9amkahhWxKebnG5jqq
LBnyI7pw3RqXDFmsw8GRSXpkwXDkZHGYjyHqe7FytUH5MhsCbWWn04VoimQ0Sn4ynz1Bl+Dug9na
0QeoIomVDdH3V+8rplNqr426Ht9kEbiteXOGswUplVUD1w+FwEimCDWrts4mihMyTLCpV3CBKLdE
3kfGAh5HxO83yiL1xx0+GFcRQqqNAOzZLCNjteCsB+kUj1dVRMg/iN2GBbS1kzoAcQTsf+UiaZI5
rIihpa3tmWN8ozVyN0K0xS/IGupZI8XX3ne1PyRtBqNpWI2SaBSmXWqw6RcR/JTL95GdT3Ocqyg7
3o/zh1S6TsGYPxMD3d+kQdFEjce0CUEkFv4o0gOu2Et2B1YSEMr0ysp9VVftVX23rQyDdTYjT1Rq
LudBWr7owehgqdmA8h9bzhYpyD4fsACEVZkYtzLE54RecGG3uTlXDxIxqV48vz8/qfno7ZAhSeCJ
O5TmWKInLAEoPpdJEVZdKhAVN5rO0FSccHIdjvogxx4PK/03BmIGzOFgz4mq3ITCtv73z/nET7vZ
29Veta86DIQr1k8XobCp2iIcR9AtUu1xOd3i8mdpoKcNDXxfmWU/j7dLbWA/LchIrO75KMtu/b6H
r1fDvDXYATLaRlb8s0+PpgJ7fJEfaPLLWsr1JJMQbWAZvkb+QJs2kON2nO1GgTtx9eKdlvZ6cC7w
YlmjEcyIrGMu7eavtNsmLcg/K8h+cO/PEwkL/QqpimyyFOI9dlv1cU3gWSqHtf8otJuxhiEZlwWx
5lr5S1SQkFwyYw3f/do/AqJmxiBwGvNg7TJe2MaB+WW0Znvja0aEUgrADYAwP6e67KZzMrrYojOx
lK2J8zG2XGLCO5rkxAfG3RcY+/7+apz/Wo47LMYCgOHibuAyyGAOysD/w/n/LdosmXiJwsFvJ72z
My/0SBY2CO9SM0vD3aksqryx9eBJbY7m61ZWjn2BZZaavjldUPbr+3lAlhdpsUVmd2/JVAqUjQIe
l/jTxgWER+5V1AZXZFp10mDzsvhwaEcRuVJ5NLX3OdwLu9Lk7Uxg9HudaAN9LAvLSzH1A8eQsOvh
4PQ4n+cDEbbM7bg5ZgZb4BazE+Gy7IsHPQaDNdl+mRK4ogH8zX+cvEM0az8bU2N6XzOkErm6kTKn
/TGNEHxLc+kei+2HNtviLDn5ve7J6QniWOdTbtfBcth1r1YNTwirrEo0yviiNstYpLaYSlgcv6qD
gWsIe3FDrCU/0GXH9Ysk2joAySKCbzhrMhwy7mwYlOd1NJoehpnHDscFj2cC/XoP8yav87E72TLe
MwpQ+6vXHxMY66PSYePXpZKepmRw4sz145G+jrLb0J8IA++H4wsawJ3M7NJmM4qsusJtBOv0NGNV
+M/fRPxqDuqO2owhXQXY8xekkKrg8xb8b25EXkyjU0y8pVkgMDqzZ1hG1RM11uAq70GszQAa+OdI
w2jQv1QFXe/ZZC6ylgptrgu80mVVUce4wo+YxpRj0EG/BxfYU9OXCrnHPBxea6zub7gsOFQK+IE6
/DvlWRocRf6tdeN8/u+b/vd4AIuIpXRH8IFDv07SqKKgDQS9h/4s1fYtTvSLkMpWYrOXJUG6rmoq
VWa+rAcPF13FK2GF0nvCX2oALb3dZkEKF4h3BY3F97wReIewFnP/C5679ZMmfGJZXPtY/VgLQ3BM
Re5ky6l7FmxJiJ0zE30Eqc43fU6TiBl5DHxsXutZ6obQhluIkTCUqHeQzPTPTac1gwJYPeoBloSH
JJ8s5aw2sCOqYRF6G6YRtewt5ejnkXG+q9gZkamz9mk1tGjsz5lYHLOJSQEZmSzs0a4CcIsYcC2w
yt9UMZxs8UGGLbW7m1UQEsAcVsDIW17/uMkhXTbWd9PuO1QUpRAsOtZJrkwwV0F+7ZNgDi+D3xFJ
K7NmbwGCiC3fbdifnR4/qY0piPiX1mJh7lVce85PjnMpoBhUC1Krtgr/1jIvr/S8foFPpAEdF5tb
uybCgYuumHGU0L5zurewWzGBMamWSyxkHWIdY+ZWyb9lIqHEfsKlaogBxg10V/O2hf0invRZkX5O
CaS05RP6NSM/F6/Eaew1RPFfX3fUdCyhwD4xwewSE2WlbdqHE7Vn3ks6vbyBbog8JcABB/DQwqmo
NBqfwtN1+AyzqAWEPH3tH89BkD7T7+xKaNC4z9aQxvAU+wQRe2mZmD0wjm7Xfh0e4fFvnESoF8ds
x/uT1BSGlvGzJtDud4xNTp0mFoNwf/FIbtxVgSJCoB90fK8R5s1IZuLWZyMjSnMHBhpjpTTfXvoC
wA1t5Xhehjysv60yS/BNdSXwV8BnfWDqY/R1xOo90+Zq7gzYp1zLtBdm+t3W0vJwzJK1EI5N2yTm
Q4vpuA9CPyORV4TKMsBNO+LxHJ/jHwC3AxVQHv8opIl0qz1pRAmita3ts8gfesqiwkbPaK9+nTEc
e9ZVDhZ8an1xOTAgtoDhpbUYyMyiVs7a0mg0sbcnk51q80HdPb+lA8YFMPolAyZ5G+O1PO6qyLHl
afXC4hk7eDO/P2ooIvOSNXQz/pqQKp4tjZyT3PL76k89fIxFdOP+6vWGwtYbkVapMLvtzUUiPRqU
ja0sd0YoXjWpFcqiil9NAp/IwudDvp2g3/9PQ3KGEaiLXE1UIRL/Sx7qduwVDtiRPgFPpUkjApyJ
6qeJ4J8ljMITnuzn6lZwGjm0MQXB4TVdkQeYBpJ7h8rHQJZ0HZboxHDhAcyD8Ldiov6fgrn2wix5
FME6Dc3VyFs7lVQ4Tg8GueGPCW9C0p3Px8bw/ZbtgoiitJflcVl5eriuQf88yXiX4/o0qplb9QTV
Wn9luxZpaT1lCcfr351XIYJvvEVDSjc1tFdCggnPiTyjOqNTtH6foKFoZoJsFVLDXiNYOEAHQ5Zn
7H9M9W1JhyoRiJ0Vi2RvZtaa+UxJh71fU94hLTSmWyrb9iWTgNLkZAs8NeDfIq5oSUOqoBszJhKl
Kl4ZnhA+iIm8AKaFkivh7QpirbJVYtljnmzCwRP7nV10dJOPbW7w9BRKsXR8yU6Hi16AzvW3H4qG
z9qmw9Ql3q8ZMGINHb2Y7FLzytYZeNWjKgtdHcykdfgi3SsgUG9kNDoIBTb7Q2wn9K6QShjYyGiZ
D1TwBhTrz+Sn41FPt8ENd/HOWlIdzhXpbv7FRLSn+5Nn45V0i8W+JwA0XRQCrZQeQak5FYQRW7m+
AQunzEt9XxmtmyRD8xSizlGwaWGOtVlcegiwioSZ+dOQcHaZhnAqS0DpsVUdMUmNmvmds/wLa3JT
PEi+3yRpenMINxz5ScGCCH3ogzA0V/75VkmPu7b6vqZ3Eq5cNx5rKogFAFHI+QlWidZ9I6Zxm/5a
TH9BO2G7C1A2fGtW7lr+D2P/tYuE5gose+kXUxrN56gxe1ceQLXuwfPrG/ItgMwVxfVI04/SXMzs
w1Nob/OVv9/R0u5HovuqBmivbxDXbta+KSKZwQgRlJ904FqWO3HN26KYfrcL+gRIAOSSMYrSWrBJ
mcjNiZi1MlhRfTqHuuVZLkOjF2ds9zZNVNOulrAOdahVPX0XdOFPf4VBvU6dOuEe3K1yrFvpgoHa
BfcHA1PCl250pzKLBiKSnRNNZ7WdBoJLoA7+HDF4AGwhGv52E8NbV9RUQaUCazTqP3LOq1YO53Jy
WdRJPRL2PAHMutJCXdw9EADSC+14TEQ2sOJTpq1neLxyRtMcu5Gz7+AKqBgVHqCMkahSBV5bCuas
/dcp/jeDi6u+78+mV1ZewOt9nEhKvcCpc02mpN3EPxfWOqssm6slwKS7X8w43HuCWSM4rHgRK5fZ
M+oOAa0DVcG9VWeEKxWjki+DbDu2lLmJlAt5aVmwABCp+wONaCc2yhzV7LPIY8nkTr5otSbyDqgJ
FAol+OvEdM0dvrcWLSpdlxBVc3Eql547XOkOepzzdENbIuL9PvU8ugaPKqowofXKh1cx15X+0nhD
WIM02Oa+zJhuPlfnaFzsmDEiHRX7a/ERs1rYph2MilUO4nVM0Q5icFAaoR6w8WmtX5/Cic5TJ2L6
v/oDCuP60D+A8LuCmlHqXNkf4hXzwGydJsD6i6WJIyj457tBBB5d1o0RPXRtPun1b615i9ehRX0k
pDNA+VEqyNv4FePAQJiXv6VvxL7QBM/W9Xm243zbYMY1mq/1TDNgpHuvi3iOxV66UkYq79HrTkay
7Vv9osxazd0Ef4KH1gYu+dioKTss/JJDKAZOHxox6RBkmDcxLo3wUUl1CG4NrxDSChU8Bc2bUT+o
dfcU58s2LkGoq4AkfxDrQwxVZniEQm0iGPLQmBk7KVN7CxEuPiDsJ0EyOcgDoVT1YGL8v1L60qCN
9lViMRofbnyRBosvt5dfTW4BYWS3FA7k7cFpnNoqj9R7nSbny5X6zVot+jzQRB5J6dd+1fzLBi+P
xOX0ausdh8XIU8D2+bJe7uKU4N3vtWCTyB4dVaf/g/ziAq8bk5dcW1xgOe6s81Gi7UB5LQXQ0wHB
gb7OizZszIGIQrRxgk5LQcOOgGnM325cddBVKJTx78W0pvpFAxGMjln6D/x6aDOc1AftwpO+a8j+
ooEvC+GZBvym5wMHgJX8LB9kHKgFpqCw4Szd35yk1Wg7ZhqJS5rr1F70Gdr53wgLdDVnGHcg6HmL
ebW/FYn/yGfTgowBLuUKDjoGkV39rQuBIsq/JOFZM64jeP2ZovCFaLXajNyGUdkZLVtl36+s15g1
0dqath7opunwcrxQRgoe2ri7mKHAs2szioif3S7x7zgiltbIq1zh5xt9O0PWG1nZ2al4DHlixaQo
kQ7pra/cSIk+CoSQvD7K0ijyNDtLvch4oYhpFsHzGGQI0HH+vlscRJeO/vookoKHNLRuuopXv/Fk
Fofddt5eAZK0raLeNAR/2LOjkW2bSUDrMtoFa92RDjsbsMfR7UBvl8s+7RjW5k6kFtI6iCu9uG4L
0s8LSN+m3u12UsaPcyA/2xUJHSRuBbUQbjWOLtk5Y/f8XQbZ0HGXmNrJsl3aB1hMxUpS7p2OCrv7
rrZfW/k4KER4ZPMR81MJzpl7jC9fVb+sTEoimRNLC8z4hvlrcv/iH0L1dmssRbQdg1Y6STPDUgjX
ZcdhVo9RHUbQmSjDCISU0UG2qrlJIz7qzqM24vFM0zI2NEc+Dy5DuMR2xGmtm+eBgGKETHt5PfF7
fi1yoxysZ41uMNmAS47QMz2ixslX2mUxr0mBAzS3ujnzArQG1wlCuN4mHBPDVuAKv1H1gBJCnsld
1d0OuaV87JQ1+8DEravRHwaB1cQEFjSntLbEHjI76j3ZXLR/BTWaiRrTCzcuCFsThbBGYZKJdhPZ
pYgqhkpOkBR9/9HssIIVnZStYC6fsH5+PETr7XS5f0kW23X2G2o/DqgzBssUTnN7cUq1ljyVmu56
7cTsmZbr1468DexM75pt5llrV78ZlAdeKjXJqX0KscKo2iKl2wSNZ2Tvfom9K3O1fWlOWQEjHLd7
KvsMB4lo51f/oWRZPHIgwKUtv44EelWF+zrmyBppWDbqkYoHTXV+Qyfba/Yk+y4exvBiTW1TIzBL
3PQW7Rgj9vxDuXuPNj7Sm3M+ygoDVvTxMlVGNCJ6QakNEaCh0SS/DBMWChBxT0D+B9/GD7bNbwX/
rsfhHYchIjLVxu11ufSjQqR6xX82XNRjQhb+tXk9ASHUMqC5agoSxJtXSaU7w9TbAAbaulx3c5uD
QBLz/R8DccSRQdDcVc3zXwaYpZWS1LiSsguzT90nw2paAs51F5iHyN0Vwc7jURhhrA+1SFrB91pN
z7TjBSUr7Ooe/d4ogA/uRoYTSCy1RRWLH5Q+PNDO1lqpkvFYHC+Ido8UXQKrpnsrvX3J70oGEjVR
4Ujiko7Zj0h1Hg9XAP0VDsj0yBrdauq6s2iZIUy2OQK0lYo9M1XLKzWXwBqgOWTM1ksa5d4SGUIE
8tlxwjLOu1aq/jKzFyDsBrpaldnHDU6FsqmAcO0/ja3yVAms1ACs9flkbO2hVIA8ajLaxkwZQI6d
aTVLzj/G5bxE5DFrBiKYUiEs2i3DujnwZdb3Vw3if82HL2otkFpxqgTY38lzLwXHqQ5WrfxyXH2Z
8jhbvjnf76CNywKerZLka2L74AsEuQr6kY4dK2PsV528sJTzDUzR6isPUwe1I//WZpNkOfA9l1z8
X1y4JfrW8wGOpfTHrpWKBZWEgia3Yt2EiJ3M8PS7fnZDtOChjMtxaQxXeP7l7OKaNirzTvCbx9ul
TygPWZevb2j+26BC3w7u/MrmiXVcyOA0RVliSsfGToQ00chGLJ+uhUWK4pAW90eQuc1YWkI5yy/E
TDlT8RRjje/nMZgK0ibzr/8uLhVG2FdWoxn6GWut1kXUKNrmaxlYNMSg2UOat2jpoHn0AbLxfZ5g
OhQCaF9A7+mpRpqFK2Boov688OoUAAx4wAsUDHwdIvU+/4JESxmYeW+yYFxdy005WFbbJaVjABIT
4JemV7XTT5oNwRp6fXYetstw0JUNMFaYoZ+UFGgCSPJw90RMdSchYuK4jL85dcspcQA7cXDfHRr+
AC9omEOgU6JG/OjJZmUDnPdVAd0mQy7Y1Wv3JSOsKn5oMx0e/A5GwKoU0aMp5XHSFkQpVAE8aTNe
vPho7bZhHlADPmRIEWLTTl0K8O1jt5XEKXgtR19vDQ2qewUJ40zF7cKniYBQ3cLH3nnhSZ3lkUbC
yL7oIJPbV/m6lmGdOVW9/kKKctYr7pon4jgBJRdNRj1NiPz5uXDAjg7cDSW4ncCvwmLJUaixtaR2
9QETrkfsmuF/MwhlLhs0VGuP2KbX20hUW+BVS5nGZuX2egtMN3BMFg6QKEhgVYSrTJarK7lhVeNM
NuzBd8hhCjOc9yZYCVx3sZSLaAr2v/d/MSbFphnfBXuHxvRvVQ2j/+xm3t+f5wszsj+/bkDp4OkJ
Hda2TUmKEXtwrrNqItb+kKHtabLbdFuZKIhKtmqxN4c9b4tH76y3wMjSXBibWi4Sa42lX0sy8pT1
FsPhfLUsMfBnSbxQJw+H2y1po4XJ0LgVqQ2My/FrkL5Cx42pSflu2boYV8nxKdfEf/opllbYN5Ts
XXjoeihhVRCh5mli52bFvY+UzzEJkTVFR/QhFKK/eS8pQDuVs2hJ0REiCrdxLSMSIkrk/lyaD+co
5+bYqPDHPlArsj7un3YXlATdDXVwj8HIIdxOw1Jge5DOYAew6EnfO6I0OW9WHEE8Ozb7DX0l8Gvp
7EGSXh4OP4zDEsgTQrPZzo3n3OVizpsbKMI7WJ1pUB5+f7llvMsykfZf0WsX3xUMYhUVWDjqkX0q
F9EmVHV4tsGn2+FwdZooZcjOCuWi1QG7DYiOBk2MS4WWXf08iaEdMCxMxmCqj0A0oQDMTzg9/ya3
CuGTM2XVaTK5UQhFf6ucudMqPfvvMydx9jqS/BMCtKotu9AQnLjxcmvdcwTEwtPEFsBoJjKddhYa
2x3C5g17L7+8cFHDDvvPpUzq0SxX5TjnHgC61QYbTzoNRxQg1cy5tc7DVK1AW/X2JvlUPo73Q0ww
d5b/vtxhV0OPGO0IQu9LTsdaZkeoaBCwqOqSIQMADoLXbCXUeckss5qsaCr1KHYnvAh9+rFbXXg0
jm0fCuRbhCu5iSPHNtRa7GktGphp6bQLO/vgMM3AbWAUkHttHQ1JZ6kRjVikb9Wxs8651BDwIs80
ZRutKYx9b5cyzGLDyyFWpJC21nd2gqTnCYoDvbSLPlbWHsLjlUboeiULeOmgNsFckwehE2wrgr0Y
/V2RvUFyLcGrEUkKy6nM/7BsV9qP3yGXvBsD8U666nNqSo1fnfC/Ttapj8QNsU/G2i+PeOvOHPze
L7tAQUZBajWeW/9RRIcvmJ8qZbZJlTSMRyue6uZfsF1GMZUFJjNvaL9L7sCmNg4tmA0SuUXp06Da
310K0jPoCa2HxApSXgq03XCKgz65EVmaYSRFhRokJhON/Iqnq+99yIlz1PgaweFdg0ZnG3Z6akuO
f7m/sDZuZGlyuHolROlsqLJTTZe/RscuOqCs9m4FPsIIyYr8Zp7DMnPzoD29GBZvY8NTg1/mqC15
coaUlgOkr8/PV7Ek/DtW4cZ9rn0FYXCEkVohfDu9mdFGZ2cQWIAhv3Ukqraj4N8YPt8+xcTO4LtE
XeYlMABvJac/zMLn8fnmI1t20MJiKDzF4gUR0zGStqFNYjzzV3A4CMBX80Xhryubv9qzVAiBrO8z
PSaX9A1f3tGo5WGACYPcDHjH/Q/3BbPrvjsajIuSdM30pNTBiZEw4t4nyyoxJ333+/KVTHjOYGQu
xKXLvyJ8KlZRNM+DxEMB8ZGxg2tWoQ2yf2Ev3oeSvV+8ywWhgawcjqklDNOVOJb79nGjrsgwl4sf
b+IBuM9SfTRyL1yfM0s2xWAmgd5EXByjL5ze9QP26eqZWSzxzC11BSafZCSt4CBQMecmYJFtuu7/
7IO34gVO/lwNEt/f8nPRMEcugc/Siz67aZHvWUjCrSjEHSfXaG/g0tBRGGutI3tbo85hObTlnfOp
Zy+YW4vVNAtxJ3NgEM511Q1NaSLJCyktfswmO/ASVmprT8S9+UYEoeBhsNsaroeEyDVPms79LV6A
XHggFdguPIEK6HA913VvLunx581rq8PGy3fgRunDdrPZaJmBzXuk7Ih2Pbemg9+J6AP5DIs4tE/t
I4T+pS3bNRdPfdVzuK5Ceoxicc/LO08l9pk6c1cPMlmXu4sWmJSmYqoiGRZ78YwaSlwqAlqXY3Id
lcywNxZMTdF65jrI+RYnz09fnroW2nyLAQKX2LVgOpEkRMfMYg7Wnqb07upc/l8yRNtQMFw0Kgg2
2ff7k1FqlMZmnKXG3y5wqqibAv1nDpkyPhOmho4X1O1hazDoTvEsMd0O6i2k271dYuru4kVXvR5w
N4mmamJ8Bua8Itylhx5f0oym9JyFqU9YP5QrOgg+ReWwkir+vlLoiRuuWq9DN+XkNg/eipbmK0Jx
vE44r4ujOXaVcmHP+ZkNkTSQKxZGwQV73AdnUbesiGEzFdzAgi92agjmrI+WQWH0HMJGqf/DzVoF
fkFkXLzjaCubZr+ZbFjs1dUTWkJ/yg8Y9afDI3QSE1S5L66FX595KFMmR3lmkIcCNQBqAaOwrksH
G41SQ/EGQ8hqanGwk3rZiKlnv0fvuimIF1YY/oqsgX2V5W1C14xLEAHeeSM/YmZZRFLnZLsB0K1N
YBAFkZlKwl5paavRrVG3NyKEWgy5djrT5w3eepzslydMM0Ik9lpBxQS3AQC9MRHF/PiTTuYIQMQJ
AJ84QPHlmHFmDNKsaIylZDfSsvJoHithuHBG4/vrNdD0rMbXfoGawhkRlDJeOhFEoUuKBnsUNpiX
sh9sZYP7dExaSu7YJ2FtoKHsIWDDtFioSqzFG6ZXxDmXtRqvkDTsPZxfWhGXNjA5roKt6r7ZYjPT
dm7mSiLuYsgOdYLfgzXvnIXQIp7i7F04ymgHky3vBFd0vngcMPTUWsS/I9zajtfndmM2jou0LgSr
cZXvGVpKeBZAWr5QWYdTv6ltYZOIiyxU1lDXXMW534wztK+9Xw9wI1MYndGTAOE+WNEqXgF32FlM
Jxo058/coDCV2138ztr5Pfz03cz8Ugs9y4tlAYhxeBsSUYuOQfZ5rppPsemmAANrQx7r7vHU465O
EL1N2YPNtvUvgjgCpkIv9qCji5899uCFL6xzC1FQb3LlLG50nEgHtGpb1uyjNTYWEv7XjevScXxX
p0V58SpOiBnXyJTooyvuJ55XFRk17dGsgfcxDcUj8Nr3rmWMtZ/8ykxKFMRDmqBM4cvFSQVmmz5j
1MsUKidfHFifmtOqmrY4AznUs1FjwBmGscdkTq1RixYoEiqN1LEBhg1MVu1/oi9I/21mbU5xW+DN
pegMBsG2n6ueoWDZes5WvnHkxZBCX8gx8yMJeDMYzJzoyv7UNJQWBmhzZbSt5RsB8FFLzl97eTXk
Y0ovXN1d2loyK2NdWTWawDyx5/GnW69E01zNZExgHNLt8hEvGvycd4AyY5bQum1wcxK1vCNQwgNI
dYvzzIZW7kj+yfZvq+jasLXB1t08/QzeRsHxkKzFiVJeryo4JPeOnHDnmm0v3qZkv2C5BbOJD66U
aBXBblNtPbFGNprZWsPjHGSs5zgVR47hiDbkdn81A2R28kzXnQwjfr8MwpIjm2KDoi7kXHa5B/ge
TsRbkRtY74cO426GogU12RFj12Ivt8L+5/whYluGmzGs2FkIvR5Jdu4V48Z9Bozieuv1U0ASTzqy
c2R1+2+UzP6iGGsc5ZRLvIULi6/V+hmRYog29ulHvF50UPYfyOPvmdONcGPeJ5xtpMLyEYbOFNll
oFj+nQyXv1rFvTpb3l+c4vPtE/ORB36rvyodWPmX47YKqRWA2ftcfCClZDyIj02JgNQO8qNWqg3x
DCQCvXJwDmzc7uryBaSYYeXSXROj3R5wxg+WE5YzZ5/Gi4lPT3ayKLdFlDZPx0sbVW6Cu+HgQEj+
03ynfMI2Lild+82uEvTuQg/LSb9dDUdSg2vDc9cKjMDTjuUuJFWXPzqEs4GF7/p1ynrTIQ6ERHhK
ww1Fu4hz/6wBiby7s6OhIjuRPjv02tSOti/LJAdv8zlPEXJI/I/l5wvmQcW+9b4HjvDla1inx6wZ
fGa8fomjc89B2K4toaWCcmw0i6/7Tlxo+cn5XUfrqwoRWPGjrgz8iGk/1R96jy7YaJB8A6wOZmS7
Jx7Ok0+KmZ+o4NDgd/Rd0SobG6EJGmij5czO0H6VTZs5Q8BaDyX2GL0vDDYkvp3oy9U6endcOoQr
EA3DFofA6AC0T48mjAaf2ZwgoKeB3yvKUi61ckDf4fpBAXmdZJ10Qge03R+Fu3s5Y3cBk7RB/MLR
+qgCyZ0NEj4edXLC7ID3Jsmh0WVUeQqIJ3JnrOGz4VIjODQXCB126P+Jk5R+4bpVWKB/ArAf2egy
FDhqwjaF6Rrd6E3w5tJdj6uRCFNWREzVXKaYcPd5flumXdKyr075gB6McX6AbziMfNmJrdCJNutW
2bVAEsEKwBWf/izwqwqnE+LpSkeJZMa5xlsaiJgSq+nv9fuz6Wy2J+wG5R239ttho7QogzawYtea
bJwim2UGhVd0BVuT11QfFiERl3Hxvaxyv66ZWqPBw+4E4h1Ybxfav+ObvRo+nNL/STcmxCqqelML
//0myFNMf9X6tNniMSwj7ylkIFD+TIHOJh+2lO5sYq2/6x6tPbNHBmhiVwgvbp+FewFVP4gTBXid
1VasuhITi1Id6SwaXBqSCiXP/P77u6MlDUMvr90sBGAmZzuvderjHTQiZWdhPGy8SD2yYCbR6OEC
sXyzZQZb3bCEX57bg6IUmXtPWPO1nCcgr+5UtRo3XFgizmbwUae2ibI6CZx5TV5nG/vdfNeYRQW4
LpnV89kWKbhZSvkJsVYLbvQ0NT1Uv6N7S0cYIMXIdLgug1GDSlkPX7Ikr7rs8QYlGxJTAzUVc0AV
x9EUgwHt4uuykizNCrVVmhvIOEkrJfT1u6lqifQURgexrx/h7bMHrD+v/Z6fezjSFYwodTX2MoJG
xjJJj1c/qPtLfcVpq0EvWZUgOD7Ew1O2Y3fjQpFqNPyjJxb9ntEcezgdFi4HO9eWGL2PlXUThA+/
g8Q6bmUWcNIKgA746+2B4CM1vCXF+mIbQb97quiZ/SJIIQuNcJyJ79IzrTOBEZOdt6FwYYeSuDOB
w6CcaR+g+DfEIsJ6sUvclwaMwO87S95c3cp0hiSK4ViS+/ZyQfSpXVqk5HycwJ92pAgzOwS8qN5D
9WVHQ6R+k9rR7YOALd9rtR9k7qxoU4vOR+cdOxkYuZZvL9YfMvdGZIGX7eBLM7yEMp//ZIu1333q
UM5mrwtvD9uemR2Wz+sRToHKc/wkRYpqDBG6WBV/2iC0v6cWBRgrrUD6lVHADMM3TdX2GGg9sfbS
W2hbTPZ8u+jfJHsNIjjKTXZp8MgQXdLUikbXrjaYjw0dy4keYd4MGH/gVCyFs05nj61t3DYQzujO
7pdDZy/AdYn+TYPSr1odaJc18H4gr42IRpO1GUT4wJuRVjwKjDed5ny689mVHdQghraCVP1OZU6k
ypIcJzQQpVg1xVCxJ+rJ0QxHMtrE9nbU6Z94xYIw/hfylCXvnwxjAZJ/8GHhKkjXFulxf1Fyz3f2
6daBp1u+QpWn9MhFH/O1WVxj7aRCJ2Qj95pUP7VK+9OxrKzYxvySwrJEHqG1Nfuu4iCbfbnE9Fwh
x6weaEfFY1aIUJr5J6GM3m3gXh7xssVQgze4nLwp7O33BNO+UipzBgPVCsIBNP6jhMjdfBG8zTk4
ntPBngWIW1Bz7VZegtZ55SQTQP9gmlKY8vh5JUxRkUUDktQjntv4dBZnqFiqisA5Jn96c4VloAec
oPHqEPkHWKfr+tQNqoAJYZgrH3eb7HsiqWPiBm/Q/Vr5XUmxf96I15MyDBf5m+TVDisslTDiF8WT
47sRgfJ82TkBQNukUnwy0UgfTUcOKv3AGRD4CS3Y+w5dKKaqByp59JIk6s8rpRWvCbG2CRIkgARD
t5d4t0vynsIgJFttdU5lyr4Ho7nadMl8CabaJMw+WrGoVbBIiSc8Uj3xez6O+Q1g09Z7TLZOVXRd
Nc/kb/ftSBL3ae9TM1YKxAur/Q3JLWF7LPmTdLkCox51zuXxggVI5riZIA2hZ918vk+m1QgzxyCz
NxplqKI/Yc0qKKuJWmkRw+5E6nf/FR1xQVXWVokiQUfe/UzLBAndn6EE4IjRmqx/OyDm5k1aTvlL
Bh/sZjF66H0tAF7NZmHDJjs5q7uT86dFiGv1NiiacgCII3rxGAC7PtaMJ3LQalqrm/MI7SsNrrcm
CzgBxK5HwTMobTuBMTe9HIPp1ryOXZZY9iAxyawndFb29V/FJAJSqG0gk6xZgorNOm+b+1LrX2AT
chWYNKzZ8Vr1NJMWb5LHvUs+g/IsPrdbyxAR44NBw8f/BCqX1lx/1jbSNDQ5EdIMGzDo9UgdL7Zr
4EnSs/dnDnEkC/IEAaH/3CoSJYTPUSh0OIKDqQLPt5xfV1ILyZO87Gc23h8McQj6FTgKPXTQIooN
3BSsjvH52TEGO6l0Prz/xhk8rvV2gZzjRf+TdrZJt/UWhmYU3KqQWKvp6znUdfoMh5Gx34WJPrOa
KHGbSHv1hQELmNXrnPiV4QdW5qedSHcrJ3iW+ktkmfAehKC7CJ81BAd1vmQiAVeqne9lfuIZEnqz
IB9elsTYa5HiaOnG7tffO+UCxOEqblnxifmtCigP7rf8Yh5lMLEtbk1xCiPJyHxR4PAk33rFguN+
nWyHWDanug2yBAKKWVtv0TWpwigiO5tnsbLPR2DqfsJ30dJifEuMhbdFPVjSy8ck9kGgT4cMf3Le
juTNxTYaoV1Pftsd8A4MhEorXSBaow39/ZgRQT/lsFEacHA/txCMsjGUyVpkGjrVvK6G6U4FRrRs
FkALBoXFQRKsMuANjD6EfKy4htNG06Qc4sO9377HkiY5NK9SVppu4h2WztI2wlG4ACtzrJ1Fswnz
NgOBC0pWqIC78UWSe1pCOVXfwHxRhI2akP7++1sH3Z22v4fGOq1LeJieAx/vYD9SrKLcbIildSV+
G/8m1GYCdfWgKY+IvOC6pKCg9VEDIxky25QSHmMy3H+0sq9JfdPiHcLyHdK9I6xjrb96rrZjE/bW
SaOevPCrctyXe6QKkK1qqPexZbN0H3fzh2jWZcnbkpb/8rZmJZvm2rVtFuHYHVNCceOKboGluv4X
eDyg7B43hOetzj4ZLlT5YXQuCJmCCwP7H/uoA8GWEKrxOo8+34ydWIqe9p8RYRk25OUWU9GjklqR
IA8s4ZU3N8vs/jRpMloEwMZ3s8aPkhTDIcEkqFRodqhGKUjarv/Qr5qBJKFUTVANbMJ3WHYwkUxr
izIPPwZJzs8fdZhIP4eIOfNT6fKr+Bv/oqEXyOCRrLAccUPkqsrOb6z/eToGaDdVpe3yvQZlA2n6
xi++3uFeDyhkJtG7inLOonSIX7WND97GagxA6hhpkgHbY0FlCOQh0k4DyWyAGjzNbR7iP6CPx0JC
2gSQITH+UetRBTXwl3nBBNN/xpsd4/IOGkEbOObeqPG+eRpRgIZU1cz9e9/ZHlLak0ESvwxbmtBa
DDL2uUIpmB74Fdfx4wdtU5gp85/G99G1fWFhPvu6R8Pfp7kaYPNxnHQfFcVEpUmNI2wX5g6qDqKQ
4QIKFTgVwGVocifEkh3H4xGZaF+4nwWr4BgkOklEG5cmJNcBiIZSl+EPdYEft/hlThOVaP3WoX8N
kaA+mLgHJE1BxkdAtUAE5JN1uLwXyHjaH7KGVjcIvebMr5yf93Lu6jzpeDpZSwew/KgJnRL0vrNG
6W+kwn3o6bub/eZNh1duWUMpEIZ+qJoHZ+TuKHVBp2NsBe6RUgC79tdVbceUPTSdnGnHHo0tG1aU
1qO/19ilZVT5Oq82ZwjTSTu7biKQJPKF79loRBAMdujz0FLyAF/Wte3PBnR5kGeuTMhsRSNvgkyM
hjKiE465VCufWU1b71g6jl6FyGNh95MGfgnsQx+siIvXttHvMeYW4WqkaaueY2sXCmJ0DiXwLIgm
6E2cUMDKa6PejnPx3k22jmRxdAIBHk3mpQaP09VzYPZwnCmt22j41C7vLi13jFqP/ptQbeiKQX0o
m+W7c8DbjMVHamalNmwnwLIbaaL0qHPjnoC9Nt270JGWo0MkvFC8sr9XY4jEd65yR+unxKGTBh+A
eS2UXAynjn0VPu+ecrLuRCXhPOLp9599t/tEnmTmQursmQVwvt8CkCuJONtWMzsgxIajKVmvMLcS
z3G1j0I8oJcv51XNkDTfadeAH3AN8JiKtp1l9awxVFHpnnqmDrRfV3lopOv0fL05gB3Cz+0qX9yB
8MSY1suL/Nz9m7th2II93M51sviA8jwdNX8wzbB1irMJGlvmLeelIVzcD2qxB6v3iWgTkvPAmT0m
ScHrm8undQT9IY6jhfdBxo9ecERpKKecBaw9yvnV8jOVTnBuKihsYsDXfNmzvrmPHWqNs/EG8wZE
kBRy1FwZyby5erdoqHspvDgcG0HtO+TzG7WKH426saIi8dAnrf/3XkGwPxtG8PcGhZuL/pu9TGtA
TbVFqDya/JRdg1pFcys61zjYsllCVphsem1RBQQMmy32n+0Rsvx1YtWocFwA0uEhyzC/A2mEehdv
2JO+tjVVzlcedSUNJw3E0qRvusD92pHlGdNXwlSWJz1f8dVMIG8T07dYiTfe93AYYND0s1CXLQs6
ftMtsgS3+70wZtVe7ldnzbh0KNVDUsQhRrwSh4dQZ1UwOFrefsQ23N/xjI13CWrUZn/oA11hY6N5
UVHan48mbrltGRa9dTAwXSS6tISW4lYfKFP2DWvd4akWmPSKD2djUH6ww70M+7FL8gz4rts8V9oe
Aad7dada9ULZnOsclB8gDvoi/Tsq3uyr2W8mH64CqB6cpHFZ3GlBuAHBrT/dzEMebZDZrMvCW+nm
Un46J8MFsX5izkkzrviisXTgbjcRQhOT526TWNtKko/TxlFCvNfDp8WszG/eqJPrAf1s58Wka1O2
LQD5b21mbKYqoGrIn+vQtePvdIFP7Z80quCgvL5/I1bV1AzppmXKntFhReh07wtCWk60hEFW9Ysw
iftS/bVAJAy6eN7gCp1C1O5vOmALmImpNfCKUQZzt4ZYXkCq0AYHKH6AY7Na/Ti43O/lfSbWNWFI
QvLdfT5ERqzgh6HO50NP0S17a5zFeY3XjRSYfKe0cQWbivrJMkbB7h7ttDieLhhJNrWXiDTzLQNk
cZf2dfvmV4ZmeH434SGfHuTPHQX/44rEWrTnoPEAag6Ykgi6Thp5yXY2tdRLIaCxI2mZf44RgTPZ
8eN5snIGy+tZ6VGjxFNNctEna62SonTWXnVw02YtcLlcqzAqHVvFyZCefjDbVx+aYXn7ikhf74Og
/TFpJFtgewK8uBi/hlI6J6Rp8W8AtmsuIz6MvqUia/qzgHnzY/RvIqjFSBqsUJFeEVPAeuYwPJbb
dqLI9yVDQZsKcrvaC9Q2EoFiaN5qBXMvXk8WSedjhSoHg5SxU3l3kZHqh3lFgO/QO9grxdmaTE4t
3Vhw9tBlG3nhq0tYJS8Q1G4Dm2DJkQQt6rLu/p2PpGLA3ikMLilLAVV7gkxuRUynaeK6VWHy2FCq
TxqE+HYI5AIrdTiVWrT7m4YCTOR7YXb0otXn8mN24Hzwub1V53+9DpC+pvCbkGgJXPpxRSyb0Sle
eFxkimZAqt18wkbVyVeABKGwlovTozh5L49fhMjCjUTQ1nNqdpnXTM40i6NVncJ72WwT8mbAeEYH
YHNeuPDic8wjXsJOlGjd7sO7it2MhkdKyk008cxUBn+1B2ml6591YOnfU0BuDx0JUrxx6SvnJ9+6
2kvW0A8y/OGLPOlBHRHerHykhXAjkrSqJqg8FpIwUkAiu0qgeeUuGHyWDQUBZCKhlZy+fgg1OJEm
pFuT9ibqsL2grEgzILnZFSqUsM/ECKZyY5TqYvka5XYngBOZ/jQdGJrDeDx0n5/0i7xSWccJOMYN
Jyco+kW1TPfPvixgcaQSDxDJ9NOLPja954mxastXbZsaqOSWgqpDCqNrYdS41v2l4b9PcgGjUz3s
Wi6gPN0DyOnh0+piTdbe4vZVptVpxJeZi+NYMr6O6tqfrUr6C4fKZK40YeWc/xWdKLR3e2LUv/RL
Ei1yDninTVmhyK0EVKclW9+i4BQnvlNVRnbfwPmZVZGDVFCMCrd3984SAy3XcKE/TO4W74IC9+/r
KRIS/SC8hhNfnR5H1s539/y9Wgbl73F9Y8oY/8+PkI3r7IpW4TFfSrXPbm74F+YxViWRzOfwNbK3
aoxgsTQuuek+a1LbUH0BTNU2gwmO+uv+T6BR8xxtXGOssT0Xigxg02ZwhfVgh9J8LYzR9xO8h3ru
AyjNGxntx5JEO8cxBnJoxkbvYNz5MosDmqWSJVXOBYveplFqT33yikW1bjViqvIjI74Pfi3phAm3
tDpe+llO0AuIyNSr1PJeJJayFyqM1Rct/6gmo1toaox0tSey7Rlhuc9nktDvjhxRSbXd8FAgDIK3
pnasywmO2yOytP5B/f2hCwBe2Ny2yCat35uwdYOEKUQxSXLMpTboSJxBPcCm/VwmlhtNQfW6jZEu
S+hrAeBBFRnMICR/99fIG/3Fk0RhTEjjENLhmjiQU0EH2/rlyRWk0sHi9DfAtL2MG75l/3zsdAue
gtHTrGOGK+M78yYFV2vuhrla2unYGV4W4fXBuB2n0ytact398hLhgCkwlxP6D0d0N4p+qzGEEmQY
ZpqKjd5BOyoqOtZY3WicC3b/B2VegpqxQAI2O6pPBfqazSI43RfXQpvRpNvfxGG4iDu4k3hQ8/D8
VffCH+/Pj4MiCHxFuTW6QPzkg8gZQgEBYalYAGNosVpyDR4f4yHp0MfpyEpsJlCgRl3thk5pYtTe
g+5hYBseGGW/7lRWK8cc2YW9PbC/3tJE1BWRKu1oiCo5AGpmJ+9w4xi39k4Gh8X30oOleePd8IfR
ccdKUCnCcIubYjEmKeSWfZ4n2WigbLepCDil0Zim7DF6a8dax7KlHVX4V4tGmXU8j08e93jMz9TR
pSIps4sRuoPk12EukBFTqw+/M1p88OCQo2byN86jE/NOP+bfncCNbB1sEjQ4z9d4TR46queOYG9B
ESJgr1OMDY0UuPL76zGrU5Nqd6KYVZf4mOSDz4eDzJB7Ht2621Dg9hx71/CJ8Ye8qH/FGzwOZjPk
ghwank5czfCTFpzA5eHttRnbnJg8nFy3NO9ScLhiaWq7sNDN4kSzmPU6PaXlCPti5rT/kxFl6LNY
bkGn0jTmAUkHr8tSYXjnCYAL0SmSmJyRcgOQ47Y4dco6v/5rqFzM0M95eoFEzLi7Y0LAWYAVOiOC
7EPkV12LrCLw0HoZcrl32r8s1KAGyuBa1JuJuPup/ja4zVhVr6jSgn4xlrdhFgNExdVobldN6sCM
g/+i/PFtauv0MJQAdeTBrBWlfl4pjA/uW6pyAR2LnFWcG9H8kOkgSfhyMjasp0zz5DTEB9LHKoGv
ZlJRoVr2f/+z0qVCKBzkiwR3fqtCLDul16BaDC10qXnMYlideDgZkgu04R2dmU2Fw/dWj6w3C1A4
ZnI/fdzAirg569MQAk6n39LZmBFwMXYKS8Wi8H2KXXQekRwudplmfYN8ywFzQzTeioFWQtqvs+nr
fc6aS06AduPDf9Zn7p6p5kV4hqGY69bwrzXjs1GfO7vnzJO9oWfcd5XesW3PfzdNS26YWOUxj56t
HXch/kZqHEgfp2yx4/3qNp9uoXLQjqavfF8j2UPvMtRI6hHO9oRZkjzA7ZO4Y4E5R9LqXHumX+cC
gFQQSW5FQHR0vgXyz70B8D6UZCoJ7sQ605Y9Aps5IbhT/Aroc0n1ISYbNSmZLNt5AjrpE8KSVMe6
Cn5MUNP1sL5kdP5lGhmceNrN/6zGqwQQuzZe3VXQrILS9S8g6goa8Lbld0+GQt0pYwTWO30Zupcg
3zrLthXwoMYQaWeSpW+Ux2Mw1e0s/H/N3hj4hcuVopL9BEyjCnbxCVhxfo7ToaYGpEqPOXP42Hf6
gYpj9UJT1ZGsIzpmxQUcWUCNHTaB2EYw/ShW1Dp/59vT2pb3f6IsnvT9TOoyKEFNzi8rt2Q80gMI
F1zOoaqU+3Q5lgelHLFCnDvzfLB47B0IbwsJNaCBo7+Hn2TLEzz/s7mEKZWt9tO219suwC4gknl7
vITeWFLDgRv4WTbzuNXJh6rManKmB2p22KOcfIKXanIlcXkBNn96EKasWUcHm90JG1DfEzY3poES
nbG5rPniLr5L2E5qzkeiSiUwnPU5uvJEmAFdqw520lL25J8WXvXt7nR/fMhclFG0OoPsBXuBUC/a
SjEYeDCtH8Rp77G4en3t9BVC/MOJs2bwzTp3E90714wo6Y6/c76AnJBfWqZdCWLU4orjKtS4A42k
WL9w5w55pyqctoTIXqrlB6QVh2As75785eF9xtzKGnk4lwbr0YZ0xVUgGtisHr42pyComvAjLaok
n6cvSFpK8l2FEiPeQnkM+t+7a8TTLuhyRoll2w8yfr/c3gzlxBWI3SGnQ+6o/GZUKqe5JTdp0Omd
2/HNARM4AlnYLj9bjkoYUNL34IUEdIrRuVUlMQlTwvCooaMnMaNU+i7Zz6TWedoM81KbAOLHqVhN
IWdRr9EkrhXWhKFplLRns6/hciG9C/qrsrwb+HAZsbHsPLVxamp+K3Hkc72PteG/HNDFkrNg9fRT
TmcdgSj2NMi7K6E7qLGLP4M1dMI5QFW/yQxKB/xGBQ25dWcfuhw7C55Gw38+sIzCmMK/lVcHFYjR
h3HrLOpJoB8niVQqO48eCkOHtdiNbHBqVIIH26dJJgor7vhrP8W06AQPFigR0+DuUR/wkd5uHws2
w76sl3XcKic2nyFz3hbNgfYakr8+iNQKsOV+Z3sozHnesRdcNtLlGbX9WLVuiZsack1PWOaM3lem
pUy/c8LyW0peOnrTfq+4RsdTMF8+E+XNiUu1JBd91XqVqTnCB7kr9FD0J5caXKU4u40lVzcBPc6d
x9Ju8xWyrY+31BRrLNeJFCCccyi7812xegEkKbEOUJqUN1dEU72eNI2i1LdlwUfp9r/HAKProZK3
1zuErGAnB2UFfZX7Egjdo6xYm0gkMFOIuLQ7Ksy7jEUjK72q1XQEli0jd59LjsY7Ea8LwnENTK0h
3CMFfC3A8MufUzJq14bTAWuYyEtbWl+oo16rDJCiTB4fZeJQRyxNtNQv+IcKeQJrEjuxNvHK82ij
iLcbPwXC0tVwfsjs+KliYaVgG99xg629r2pxVfIbUh1Vq3JimWPC2HeSDnmTt5McACV4olp0TFjO
TuoGWdVmad0HrZLgmOP/DgzHPR8kpu1HI5k2p8unpku9dXu+MlLrXx2snWl8nCy+Ibm/JYsD4Jp9
xDgtENDD4YUDYDNxBlBFeZEwFm7hWaY6ALYwm1Qv1SnJkedePqyWDkliv0ZF95WsGjMnXPZBcnJI
46qVwx6r26OhP7bEH2sghmmg9ACYDf4wI0w4DFTx1nnvuR3gbKAkxpKKzTNpOXPLt8dSW10NdmPS
rqV6EUj3X0AHxrTB2gT+5SIOsNstx5K/kQpz96PxCx0HYaXdMPeK76tromlfIw7D/xmReEO5ABXt
ob0vToVMmyp79tYXLfZr6z4R6dxNASbjPD9fQX6Qxac26W4aeMoQ2hZ9WW9UUu35rqj8gEH/e9KF
1kjDPZ79lfkxudCJX9EhVpLpvod8hNUdfE4Z3V09uCaAxRs0EYKnnqZaShiy1t1qO8XU4U3aj8In
aNGfdI1xrtQoyyGBR2ITElpbZ3mG8K9K3pa7Hyd3+QIkJz9Zn1efLzscxbdOjb0gvJ/b66NuPdSA
pjrR4DTAEjROkP7tn2pmOHy/HD6CXxLHtWrhaemqd6ZOcjzQcgLFwqvf3H4pXcwIWewRb3lObAIf
eiZrmMJNi8qlH8njxI3KhQZLdTKVrV3XVvnk1NJ3RK3xJ8TlDQW0N6yAifLQDDQeAKhda5+dAalQ
Ini6C4BzOZBREJYwa2/XcDJi6BnX8ImvNiWSt8am85874l9LdTQgrCZMP51plu9hroDDCCMDWA9q
04UAYCvpPt9TXXEXcTmqMEpDqoguwvzrt483FXWCT1gJhN3IAJUzrr1pGx5e7/5ZQAS3JHwIVa3B
lWGoEKa+OhzBuarnAptCkl6ZbnfYf3/J0CQZJGpvzj4q6LeS1LSq5ewN2rOPBA9xJw69863CoSTh
epB1KnIqCpZCp5wM8iv2RfE4S+2UQrqTrvNnepq6FCdWdn7WeOxII8cklW0JcgD6LZRl9KvCIJ6V
55THjfjAwo52FOhQExWWvvvKMpsrfn5uRwUnOawhp2K4hgUFw4urtcHDOGMxuhl40O5dTwUxfPzL
x9fjz0U7moLGidoHVECVNzstCskWOUA2ftuyP183vfo7DoAoZX+rvnvHjI8h45tO//cb6fe+vuFK
Tok9uwveg35p1V7kuqU15lWkWhoVPl2s1743CdV7YsmG5Rg22/A2iGDyTHHaORdOz+b3qUK8OHgb
YdXEW2NfBiV0wHVBT6FovTkKE0Es2ndI9ZAlC3jFXmVW5zsotOhccWgsDDuVvdWIPVi5sP3wHLd3
IHjt39tzwO2LFqLJViAZrKpXGtGDnhq7X02U9t1ach7j3bcMnyN8igX+54ekqjbVU54NiuiZ62w3
51ijNX4ym3p1j/NCJmrEEB9eNqnnWnkyklBeZlZW5ba5DkpCjVoxbNgt262DNKPAqaF8bunNjuMO
W2mo+CcXUGSduxqWqetpvErQGk2BVpEP/a9W1lNhKDnEpTv+QqiVFHcob/Fpcuat06DKc9V9/tR5
0k0CGrjDleDd5yG7fsoi50B+wzAd6ZNzMcLgPn5syWywj5Bgbh+47G/bRKHBN/zHKXAKbE1ygFPq
t5VY2jpxCtXe5eGkXl1V16FqaPkJgEmRWb3YMx01o0BxhsZuYSjmiVvX7dN6n1tjtondIRDVEoqb
D+TjFHJUmP7zRJfEAMhdpiTpStigsT2IRYuKgXsK47g+5RXBYta5ROpTIDG/8kUTaBM0zXe7MPYW
NSX/sY510Bt5lLEfZK+N/OIlUzc99Ik8A9QpTZoCm4WDxmx/6I1TM4XTyxuRHvWlsguLuY8QeBQw
YS7sBxIPkNWnqlJVvI4SXVtRor6dRtH0jlwrkvpRu5khd32EAIvDTy+Z+El4WEc97VQ17O0OpTma
O3sstFV9Up+7WDIoWcXmvb7WEOKQwvY64RxE4Xd1224D6aSbltcFSJZkZAvnWuZLXSQH264XWHFp
SEXrSWrwCknE04+pfJbcbbfbF8kNzCrHOrs+OpUa2WOn9RzpKCVy4hIM1UL5B2hG5DVbDkSfnRRm
BLZ2LJGqXRD5Xe3Bk4WLqzzeK5uPWFnrPwlbS32Vk2ltVZ4rDPnShjZRGz32eZiHeaGeUWYPx+ri
MWxRUW0G2yvGJOzMsO5C70gTl568OnigGGXnjilUY4+/g5t1xp2pQSJ5xlaTLFvAJRTmdJVjjh1B
pUJIPCgXsfY7wskoyGWAvvuW9X0gk3I0N0Us8GnNtexoH9d0ofXDCjniwevc74f1jSc4oq5Xl0to
TPodpAbxTQWSayUVsMe1RZRDRL5T57q0tAVgRcY1e9rhijyeLeQGoYyWX4VGOVaj2tW28Fs3QU/i
agxKgTv8eOiG+OtzbfNqbc3PYzqVuePnE4gXk+3kip6Be98d994+OTM0mUpCKB2asjttDQyE1DIv
0DItQAExO73OdRd2qshlchdOFsSHnozAWWC1F96VygAKsamPzc5rBRODcxAGfmcpY74DRzDTk/f1
J+uKY9unkLktw9BmoBgqQ+dGikm20DIGlOw7nSoFecS8Q2ysXEBpEkMTUldWv/QlF/yYLwko0m1f
lGc9oWwMPF5yDVEyvMjDKqxgMwL9h1U5mMbZC2tH+ZT+q4E5Iq4ha4Jy9vTs1ee0ximjQyOz9F6F
DxJhtGPgEIoMpbMgfqzvlIteyLogHwEpIbbWjk+/LRnHv6NOarwEDZYvCA7ZfbRL4d/eI0nhFcNm
4H7XRCa64tF+FIe+h4h9LNHpHHHek3Q4MGpXHep8oA7V/tWOfVGGkxgEBIjHwgZ3wvmX2t3daew7
VlvM0Az6T1eNx/4YR+V/fXHx1kLiTfv0tzuSMUTwaKLXvSDBllZAffnmdi4N10PKIwgv8XF1Haam
2nUO9rq3GUgXXJW1c0K3JrepdZyZRg54P2bWDJaD+KqzGx/Vuh5rHBCLFKE6yupW7lMzpdY5dw/h
1/1sq//TY05ldWvDF3nllUaV+lVLqTKIDV+hI86nnw54Wwvq8Q83d3VCklTy9hVxE4piqYWvnRDd
Fi99GabkvymeJd8Uu09MB0710QEEO9QxIRYETTBpxQcx/dsPYPHYy0BvMyQ9M2HrzdG+PFmyLl64
pewmyttQIPva6Zwgg+AGyzm3ZciDzh4hO9RfJVXPHpPLh93HbHe6ZIhQpR0ZsjDUUj/poF0VTNrs
EMyY4QwAyLXqFNK7g0WFSt18p/RHdU/C+2jXzV9I04US0pGgmsCsAARCJP6GTzdtxY9CuoElHkc1
g0R9MA6Aej40pZlsEz2IQfybUD122BANh9c4t4uH/i3vWEHlBpdJxUTD/da1npLzSLsDm32XpO4T
sJO55fuvvTHj1DTG3ynvpCLJrS+totp3IZiL4P6zC9ZE1hvoSdujziHTdcUccmAFs4OA8373EU3k
a2XntMHgndhghgtljP+T2bYdo2k+n7FQbucFuXj5mEg+lB2dOlbXersueqIkLDlAtDpwBY9UVeOd
XmVxabpLRRw6XJyjji2I/E1UugpK421y8NzqTgPOX9mc6caz60cKAAUqb5jrGE5ZJQiwewMgjzD8
p4SjiG6qgQktOWmFEXDoxiXalRkN414wOmABFMDh0ocTyTh1kC7o6IfACGObelz2uriEuiCtGQGP
aDtFMaV3b5mZc9NUFQBRoAty3ZmfzhOnYnQWck9vfa/YB0SQRO/s4gI2krrgKhgAhPsimoQc6PoF
C+9wm+4lo1D1vS3HPeqXQjI1lfsA90zCjBUXN4OaukvY9pIJBvvB8s4QyRYsRIuhy3i6/PgszmyP
a6UkGZ9B+j5MSuK/0RVJBNfeqz5CI5gDLGadx/OT0m6+zWMjNrfsjuEtO7IEmLbUPdPjhzSb6A+A
9k0s59VY2HOmN2YeOUZ/v6HI417ClAzPIosvT/iwYaNPvdKDfgL9U2K5LF/dtR7aZd/k44WVPjUD
fiWrT9ek7RlDfcOOJBQmkJgHls5ArvLzKs96yxSc//q2BDziHf/XdD+5cC+SVW3cOfam/QW+rTvs
e5qv+ZJo+1H0zFhp8d/uTkBAW+6VumEd2zkbAKqFooC6nOlFA+DW3RefC+6P7WkI2U620rC2ajwt
GnelUzFdpoOCDIQlIKZcdwxgjrY+r9dEdLWiWXr5uAehCzcbfEs+7mL5UxM8TjD8CK0sH3OElp9p
Kmn1SwU8bNoHgM2oNQoLCQrf7N6tLild46tHeLOlIKjBqGmfJtMnQKpGyWUtPJurIaI/8uZU2lin
0SC8Ozo1pJ/bEWAxWyMkc4AqxGI+SphVvOEDcvkvtPXDDpYLZW+Lzrr1JpjyEXTY8/8z348USWhy
xHsTKZswloXbJ4fSlvjIDjwRGxJkCgBHrqhYy67qifHB+fEsYGVnIr/mhb+3h7DrNklC5tFaZ7D8
cBB0Y5Ny0KqNjlxa1IT26PYgnOUniBetJbTjbVUrQJeuB4PeOer0I18/85MxIPBNa4KYux6d/pzE
sFN9l1HfOS234oHgs5JNNadVk+H71oTzlZw+T19HEezFwaCjaK40PH5qJSH+1JyNzYvOZM+Uibbw
UXjmuLhE1OYf++dIrzwwnC44o6nwlzDROE+CmJn0YsbpXLcBYlEMyiWJFbpPvMoR/8tZpS2OJtVg
Odnv8WYZ9Jsb91Pdud/Le1etWL1B27QyK1c3jz2pg2toborI5MLJJtFKTQdkwuvVywIv4gZctIdf
4+1tFjd4iOGb93KgMVzFOoGnCPijNsnLPzK/aDxSVk70nkpijUKIOULQ/6DWPehiDGdWvT+QFUWn
4T7IQRhnsl/vSF5J3lXGtyFWhIiMrYZp1+3TOkKOn6AXJWGZXQMmQjLcQJx9I8lgCvTuMTl5h4nP
5ZhtfBwCKENqlVMhXQzZQA2yd2lHIMXMoHtkos9AYfS13EiwlTetjieYFUl+jBGZqZMcQhs1t+fd
bY2lSN4DHsPgeyexXg/T0DutZosrRm0b6FWIAYGTtG+oXx8jGpP1cUsJ0bfgx5LllyI7v2kIdKWV
4VXKT86zIIBQokKusmKYnurQWXPV7v/n5/2bBfAqrjfG9jiCOStbFBMqDTK2ss8NfWi+CWUczAH4
CnXKA/mnCTa2gJ0xRlBUMtZaaJICKufPncNBUPnI6TtIn6S30xIA1FErnl1Pl8lKefLXAyeiENqo
20YoPRZjI/cQwfAg8AgzHN7nyN4JhjRkvYnWtqtdPPu22JDmMaFEYRbLpNcs1WH8rKqaVXRYXBKC
aIcS3e4XyVchCqgWCKKKdVmv0gHs8GSiQAzkDlSuSmplc5iWSa2koKN/fLn0m+m/HpjpIVlaRdva
kJwuv8i+ojWh7CHCr+Jj91uido3xvI/vNO1+FHR/L7oU8w3ZQIUbzXynzfxvgVwnZyRGhJOR8BI3
QzKN1sfLyVU9sOpU4Ip5WDR6KNg2VW0V3e+mT5u/PmUlIUMkt8C+Xyw5ygiFR8bQ6GUiKKQwaD82
qrkN8xoppfxJSZHDcNf0Dfou2M5O2BRbSpT8nZchYD37YZSBgO4pog4OERYHTHwQe1QTorMi/dQ5
fEESS9q+6HoPW1iKHKzypfheUTooapEu+m8LcvFEYGUULs6EGh2U5RiH8/w3nV+hME5HYCoqEn7Q
Sn1Ckti7OmFcgsGpI8nV4FEsCPXBhsLgtT8TKfncyhKwMquckosrLpyfGa6H80f5xa/rfTn207OZ
AM/mtccukeKO3guZKG2G3w6AA+LQH1s0n38EpiKOdxzz6wbwGM8m0tDQhlbg4l0gSgWiqlfueOAH
GSldnCaZzQiQCBLsVary7+tnEM4fX0TTrFyRRQGLw4tHdQ5Tg8choS8Ny9sPg/Iv1UMqkkIUcKaG
uOWu+TXAQPu2IyzNuK8C5fynlIdt8ExUoXoRprtlWZZzVVrOaFWJsQBxLJXI6NSgApPYTLXLnZ5q
XhE8QkFlSvZCWM2Ln1hELv5yRCk9hMYZdygoZG+ZwwAFnaKN49YB7mmJMHDKO/pbX6OqAjDOkbza
A047cv6Ad2n6Mog5C6oxwqoMhUg6ewNi+KO2lT3qWjTAUV+kaEhUtejBCuEhihCLodamnBBBd07D
bV4bjkuX9r9TdFUx9R9NrWgCBQn0VojnS0T32ftWOFvqftEYVKQvgZYTFOLiiMHvf4DZKe0ntOq2
CQ09D1xY8I8c6mj4Zc/qAaTT7RhVqf4omHrbN2FyBCln6OhrsHRtHX9XzbicdQoE0dWSG/OUbuDi
a4gULgpxYlMTQwHuEgeO9XDuplGxoScpJ/trOYmH/7nfCk5l4PORs6ILA5bpLroopMXWlBRgPWgh
P6Taln5k57wUBUJe2Ba5KHOORzMzfTuzvkpsq86WX1yl07Q79fDgwin1gcK2hmtJuQ++aSxTTWu6
3Fi0Qc3qRtBjguD126mtvn7TsuaVRVfCe7bW7r6I31WNwCk9fl3SRuHfDaisxYub0RG6bn93Lq4l
pfeu2cUBpZqpkCXh4N6ua2AkqZIdjJYI71r5tffCUhdF5QLcGHFPxB3gpuhtKeYmavquJ/jAB196
FUQob6IMB+0swAC6VHwuyoEE1HKUNrHsFKSU4t1brzJSv7jz4nLInztcI4MdAKHtzsA2giCWA7rL
umhMFZmfEPRWGJCjqr2p74oq6xVW9zR1wrX2McjxluPgDvVOMHwzFhwkIET7WBDKUK84k9iLLBof
hTAzi7SsHrx+oREgWv3Q0qT8IqFiiAmDzHEYRz7mz6iQeDMOl+/do/+EA2dZFmZv+pttA9GqFg5M
MM6Q3WWFHis90YiBKkvE0bF0CRoRmCy4Pn6csWcot/JGpFWPVhiH5dBf/YjC3Amf6U9boJ9+vB0Q
w3E9wsqkR689HXDeg4GhKEa07D6Q8WfG+LEyXlC4Em6ev2tOTSux388M2NGYyiwvRNRyYf73e6wP
YPrPqRT+ly8EDdQ7V0SCuoIqQSk7MqfwKbDvuoFmU2dzN/PJWJZ/mIaIDWE66h6t+Vg7Qyy+NzUT
jIf+fWdp67qO++qlJkMuebmZw7ij6r+Zrd55asfodQQu7BT81dxLCHWRZXwKTwDafYJ8FPcyTux1
h12/a7OFdAivOC83/xKmVwMFzDPQVO7CdWy8b5g6FG+ZPA37JPO569KE6r45LjiNE327BKUcoCrK
kzE37yfNU9YxongKpiL0VYgZFZkrBx4hQSkplMqC0JpeH7Wr9ChP/hQJD+TAMlofcht2YrwQphBf
nSmmJPaOZQNbj78nIY05bO7FqjckREz9DCygI5+VbA5WnMa+GftNvoZzkp1NdQXVa68JnoUXc6qh
mopnLrqAbaTE0eVJKun75S54S4hDsYUnTnrbtAhXBWiLcXEv9BW1B8ai+66RfKf2z0EYXire432e
xN+/wOgPlNH0i65jezzPt2XetE/2OJvn3UqRbYQu/qf1ezJnIa0UwI0Da4E2UxkGgOj5ZAGFIfAq
tghJqP3OsVTgXtEz7CErQgfT/qgyxw7VC7HTJIIApBU1EZlY99HQ0/dyMlJgGMyPxn5e8Evcshjd
TJSyeqyU9WZ1Ox/zXdm0bq3AOGsCV3B4/ZPul8CZ7CawswTjh4nQxK+UbQcbYrq6ZGsfo7bds6VS
dEiE/BSqFM2vlrW6LyNJRD+YqQ6tSpo9jEen79aXW9cAIk343QhlCBGFTbmySLq1DaGwFDu8FhxS
yuPT7l76kFvdi6XB/edFdStJbhOleUDO3Iq7tdiWnkz1Gh8l+OVWzWGYa3CWRHD2IRD/nkkXJcR6
9SqVIBmiM3VnbwbJhP2dm/Y6QqA+5uuSxVihMgTxClyfr4IA1ZObOUwuy0fCk3A//8ipDt1dVYRD
SLnSzM0fKuGmTbiH9tBuRJfV/uit32Cr2WdjMNPRxFaiA06f08kKR2i9+aPIbdXr/w1BualdKaWA
gqW8fr4nQxo+XIeFv4G+qu74yeYuK/jsNOyZ/hKSZ2AsFfPn27DxhYDmWUeI1jRuzKCkGPXjBZGi
pp2ElODgZg8shAqqRTq+O5gkOzhG5iIJN8mrnmsUjTK0jF8xIhlKy/XrTJ13ZePfECPAvscDsqnM
hQ5hx0u9v6oacoClRTeGqyhwEvSgh2VMUNT2VcVg/XqwVVD6js17dFAUdx1l9n7/I2V7dKBBMFJn
62KJazmOFgCPHAphg+URHqwAAir9alixN20TF9+RpLyIx7e3RsEq+h7oGJbVsTLlNEPlTP0eXfgm
aSii6hbU2m5xPzV3zv5InxAd+yffFL3ZxxsEPfCsMtv/iSUR0Sxtqaz6GTQ7U3N/QW0iPV3l6RDH
kXghqpUBAl8+snNGcosBVloRFoFG38J7E87xhbsbg6OzaXA6YTvDh6vEYzf48ZvL1e9LfrsYbn+N
XxgAIa8oRgrHLniL/fJ8BY0Pj56FQtLCcyYvCyKpQL3xl5/Fn/71Zwq+1Gr3LVYD4jhaeQuS99Cx
pXL88K66qI5ZSd5wATFB+XjgWO9ifZ9sZ9k7+Ps5uFci4nW9hvK7RGh/mJELqwkijON/v5sWUi2m
0PkUlxTheWfSfhocn4k8B7pQtyYWPBdYD9Na7iqlO6w11IJnct5ESi40X/Hia3eK719+qwjamqFj
EwiXAx4vftzza+BXwNXwq2ua76LMIv/7hrgLZ6puVCrdWIiJlrKbE2xBBZmHPhZ6x9Y4BjYSV8E2
s5XXE9i6NqZTXGF8EYt3oTkxIGlvom7RZoHFDyLwBx06YPEEoT/kBKA4K2TOQDkE0dp4X1ru6uua
Qj5ng/JAB0RmvP477fx4awLjRAsKbtOqx6a3bgn/UewOmV2dw8K1nJz2rZUvFcJk4aykI0BWClIy
8iePjiU1x1bFnFy9cdjoXb16+5TPRlksV4u9Bv+dQ61JZvBaRjHuo05a7TM5KUcTW0gsxklS/blL
Czio9a8dt7nxcdGQFpFcCUwjgEkjsxipjWigjnyGE1d0+U39wwIroEABTWLs2RZnnY3EEA3egEIa
uRWrR/9Lzr73+Gzpa7oGgfyf+kcWIfxjuMU8vl7niQAKyn6+k2RZ8xfLeRtbu+9TPKedb1+LgNZu
tMV8PfcGbyA9K4Dr4N2TQt2n2qwDv1WPfA/Ruy0dzRQtvD1KPtQKIC1Mli7u5vc64KuOCK9UeLQ2
OHhgWd0zThg72kxIlIyznFQUby7cH27uVjYwcqN5EnuEmLF5ZyJaz6nAHBONwHuLERi4W1ZLwJfP
/oZBJax8uTJb6u4TTT77u16H02gqtrDk/B5O5vGl2kWr9VP8peLKGjty1aiizWz/WMnQuSwtLq+k
P583PyWVNjzFY42lT0YQ2CPu6nRTsi1j54Dn/Da+1QMxQhY4x76S219Qr4cBSY6ng+z4w6B9onkB
axMd+iymx6p8PUfSLX8wJ7AKk8vSCYr3ftVeSZwFN+qLk5OIeUd41fNfdm7hFSyeorox/m4384aL
aEro3VDGUhsXDbxsUOHOC/664rfwnrznIavOECduFQVASjnNYlrunc7pB8uW9lvbfew54uRKd0C2
SYVlsa0UqjBrVjFEw+SIljKyDOf3ppCDGD+xq1BQe5TF4/Zoz90HTR/4gkWOIq/u+8Uiq8JiUo82
gfRKtEij5aix6YjUyj9q+KFXQHbyikaXi8QIDTd1PEo1mNRJwQNjvMw7jNFh26WAu+5m2zYIaIOA
mO5bgT/5lLOnnTxqOJSXZV1hYEBJiE1t2iXEqu+ST6TgZQFdNlJOA+y/1PB5x2QmCd+Ha4Plsgro
eaayw5DuGgKPR+Ze/fff4Ieh5+pzBruDTMXjHCGYlJxvuZKn4boYj0QUWe9Qn0724Vdzs+cNs9K0
nNr79Bq7iRGllDobFkeME6Zkk6cw1JfmdrCmvdiVQUIgs3JsZF4HVzxxnii4EjzDrljVEF1zhuZ0
ImNJ6BaOO7b7tPHZ47v8xlUrgB5mk29Nil2iz/ynt+3/ptn0Xcvz1vYIRG2OXIGgB2EngY2ZbIL1
2v5zge1sxNmYOVX6CtkSYo7MGtAN6vtV6wNwSzaR6+Ay1+EN/CtKesUcGUvNKXYWXcBcweOZRWKW
iA+lXNr/Eg3+i5rLfpU6nf6TukrF08g3AAYYl6yyKVNm61/laOYyhMWpN0XPFn1tbMV8r0Cz8NWY
vRUlSE536oLd3FrN18OKh7pM359ZTRIHKzxNh5clhv+puB9Txq3GTi/t1cBP2kKmDufhp0YiOTku
y9NqI/kXk3Ud4Q7iphkqua4YeVdAoATvx7+5TS19cgE7py6T2MYQATQQV/3CFWNq0b/FwZX8FpBF
Zaf3KeFEgRQwubG9XIIUDLUhstFNcUhD8VP93VIGwh9G6StN9IWzZbyGuiQcO146I5GIl4cNbpsb
ic3Mmt2kBcOIN/5BI+bY/1GrbdKitYF3VKbwsKPg/dI2AGhO6m0sPs7eV+lyh4E9RZIPS5X2AjZr
Pf2QpBN0UyhvzQHiK2aea3Udxji77zviOCbW9+ZSVuZLRkdtJgErVaYvDsk5Q4zgCAtkd5Sed+E2
TT/2MdeWFv0HKhCUoEYbz2RygIVKgd2QftFRdlc7ZLtL4uRArr9uSh09HBViuc8bMLUaLUc4Gtec
CM/tRApIlCEwS1sIKEgkJIoBQ9HBNnQwvbRZ4Dmtat+WXg7XEwBtDPyjYnea+QB0wqr0ZCCfLZTR
DEjVRTWPRAgRmIgALvOczMu9IS9/Og+mknuaPQOjio6pk7VRKehEOW5oKKWDJ2veHlGITXW0azKi
b//frqL41aoM1j2OBkbxN5DziUvunPtTZYAJGw/BSY/3QlRZ53LKjIi2stgO0CizIVcgIiZyhOES
AzO7i58rSrCVEjyd/12WUMgc4R39Z3eb6CVtAiQgWONDUcIFI/yNmf0V7DD2ZPmeIq3QwJ8rdgMR
cw55mmEYx8zJDJxRG+/F1MyPKSVGoAoqLdzf5812fBLlOZlOe5WdFtJbBBJFLOOCRpCTJ8SpfxO3
mCew9EXMT5y69AX4qLw4pHPXP2jnexx8L0agDtrWTTo/+Qnx1giQ7fQcMcuedChMdyUd6PSXkmqq
Hwgx69t2FkWy3gZQqa9u6uI59IVKlXlODsy/aQS2hgbdEtexUsmhQAdaAbStCnMNqmhjDJNbjnbg
Ic+z+awCzzrt74+Avc8+yi8pbux0DxiddwGbSn9yn0ZJYzhrjJ+9TG4Tq3A9/q2VHaGGXhQpfv3M
BbYXHgB9D2L09YEOLXdW7Ip/6tjeGgKvKDJoi1rSqMObWAm+yIJ1Sb1itZpbMRztfk4eOlrnY55T
FUVOf+uSlTPp/PfpCY8EWIdDRgM3WXW6baFEB/jhyjdjEDzU0+KVS/Zp8wPyWU+F/xMezd3LrSHV
FyUne+YdWeSZgAO2JHdiWrMxZ0a42CwM3zjY8FOU18oWayFJEuI4GHE5Qb99uq5c2kSGkHC/BVoN
/Am5/7AbwWGQyFDrIiNNaVMav9DbtJ+qkddzs8EtqenNDpj9FOiIvGJeAMt7pTKpVMOX4csj6bZ+
z0m9R/vzaiQqe/cHz/xwH6A9jSAJevO+anaZMkzLnHzbCYY1Y6iAAGdwh1SUZVwYGTLk7npUxT6B
CpXiyk7uOm3tC7E1yrJSev080+R/sABG0NY8Yj6CWSC3LjCWrJq4NfosX0pyQBudiId2KvNjomGY
XdSjwbHWxtYeFbJjCxw+VsaQRnYml41KvjDw83aQ/k8Vi6BQBEpM56BVXG6BecH+kY5rlni25LQb
JTTvG50QTpgwy8jtzetvgg6Pgi1y0CA+pI8+me1LsHqYhx19l1MSyiTZSfOLwh0YXbWfHiX1iiSa
6iYM71mLm0BjXSBhYblB2b4Pvt4gJ/R6+FJznroT8BCOYyN44k+pHLsimZbuimtgrWgxkwGzhve7
X+pC9X3bZXsYC+YYBIrMdpcjGq8TbJhXHG5zbHtMA3HZJEtgmIAvV4z78xwn/38sZW8knO8L4+7K
Jm9Q5zyLB/tjl4C9niEcSCR5t9jb8vvazCMAKaELAceF3NF1ee2E0V30owdhRd9E0FYIf7lXjOrP
+83SlxFEy2+ZoWeJtobh7EovE/5RpvCj6QyPqSAiER1iczw6iMLcTp2UraXiU5U+Xn+ZpUQUEzST
A0vdLMPSuYXffB/lQ8YE5u/CNo5e9MafFF/T0wHT+UjmUCvPBPn1/LDf7Cc1L2/7QqVi7BY11GyM
1pPxxrm645Yfuzz8LYvhZXlXQvaMHldaiC8gjxAxZrSuLPOG/UUwmDy1xXoEriOss7WmilZqBE21
gAibZnpZgqnOIg360fj3bUBJe2nQIwD5zoqsihQBLSqzlyw/zEQoR+hl+THeCka81NRQ4D12S/HS
iZna8XhV93pSBVrEStGZ8PoHg6Ze3zrjRde/9UgdQ6PC7AzUxRG/1M5cgOM8C22KQyQcDDEJ+Uz4
pI3GMEN6XEm+0i4E5EM+nKGU0lQbneKFsGut5rzeScIQ2PVhE0na41+uaEHJ4C5/St70Y7rj/wvu
1M2ucL/P/usO1+qqYqgd740LZAU0YUi+vto15u1LtAtqbsICI9FWFQ2R35Kp8ckaCF7bUwkScK4f
BkhiU1LUfgXGrWoHa36m/DGJxo86XuDgjzxjdcWXRbZ9l8wka0smDfi4sjFnWemZ4fIgA1ozoJeL
rFM5uQISy1KliuJoAPpw+uKLkUTSTYZpfk/c9Dde13Bm4/PWuP3vEFrcmWaBO59LMLyof4+7j/C1
1oSKYF6wBy87vnoqEIwYvcFTEWeHGIyy3Ll22T0bHeFKQlNRCz1+xb9I8VF9NY2L0Z3CFWD+gk7p
W7HnSSU6XPbx+kBd6hF48v4qJIoTmjLNk0sPGa2e5MfRjqvRsyZQ0u4F3otIkazuCco1g3rruK1G
YDw4iAvG4ruJGxyNq2hR4VSy8x8/cnutUF9+Dz9Y/MCCo1a7eMWtYEMnst87fekf7PQ7LR1f43VY
oDD8EtmJK1Mnnq9hnMuAs5rMq225LopRjAX4LvuXe/tAAfqPAKLPKwL3yTnzs8ACtfQhdD4+VhMt
HfEVV1sFIfFNCg5z7hxs43uY2DRH6B1DKH/CBPtXt2nHZJ+KojHlOBN/DA5xgONifhq2fSJ/8eja
KPT83vULEV0eyruTMOuxTmbz4ORIS1lEN5cCFXYBZDuXQBPQ9B2fal7mRfDXzzOD387HpdYu4W00
8YWj2irKJqlY1vHyobbfHd2CV8WxTRNzjN8fYDls6oLZ3c6RFfmCZ1m3wws6lHNc19ogjLPTy2Tp
qBoZBKvUHr3dwsjQZH+RpU6qD+/r43e5UYbZAL7dVrFW+dkoHXRKsAGjnlFMgKBdDDuaxYKVu0oF
ATHYeoX7p6rooybNM4tUNKx28jPk0BE1d9Rf+RazL5bL3TVmekFlPYqmC+rjP5k1oN7UqywpmK+5
2LQuKoP3r7Zq46sE/xUonGemIOkYXHmLqzGlf8Bcsk1drFQZhEnNgPfICJNlrLpZ2U/wWqWjrivz
PJfgUyG9k1bSMinEmw16KlCjrpCcaR9gwx1Wqs+YsIbZIbmiZ13WMY8FjpliK95F7Tp+r01UDZaI
EqQE8dtrk4Wy/BSkt24Z9wRHV3dkr5iodeSNGrhdUtucNc+oFeP+MS6laXYRe+WFRx38g5mADL+S
OkSdUTCQuGmk5cb2iQjCS4MkWOWU+kKeKZrnl+gTN8hBSNyZitlWpVi6QGpKCn8VprJWqTiNiqBP
WabND+vSR3HnXzHb+28nu8ZlkaMtacibs7AZO/BJzbhYSYWKljZXSUXvgbBHn6A++9qYilDrIXN1
JhrWMNap8LJ6UK4lXWuDTqAFRX6qZRC9OyeUbNWZwHb0XmQMY0qzQYrVXzm6oIaFIYC+/ClTfMa8
OuZ1RHG7YRsHTtKJASikn3bUqS97GI3iNZoEQscp/bdtxvjmyUyf9dWy1rcsNube/Gs+jppb3Mkn
hmZnqd4Su4Tou4cL01kYEDyVRRspnzdxWw6vseT0QBjcNAy+FQh0ArlsYynfQm6oQDJfxjDFaou7
VIMmk+11e/f0ppFBHoZfNtcyzmbP0el055TaamE1GM2SVYdwgqjW6k/eVRhi3eaWC2pXqa/YwDKD
aJaUYc2je2dXRvZRwaKSotHCJTLz6sj3t9cOt/JzMJ6CgJTQCBsu1uieURFolZv6CL07ndJAZM1a
d3CnLBOYdIT1DoixdHEBGKYRfRLSDtbJ6bY3tuuCArD229zsaJznBiM79pmvsWMNah4rN+JaIfz/
ru28fTsKMQwWONrFNSRyDwZnd+R/p1k/fVaqRcco4Yc2FuygeRZS/16C9QUUwfbdrk+Gc27kGeMT
NQcQRyXzA2uMQgHCCtGC4lOTWNRSay6WUV/G7zxQ4MZ3xlxDLAwIh3QOEtifH/GRp+XQr4R/rd1E
zZobsDQXRGk1WDSjbQu/sHmSXBmnBiOheyVYyqVLZrnt5GkDcxRaQd90IrfDJmU3TqV4KrXMGg0g
27C6mdwrhdGIs4oLAn7j5j6dtt9xfo0vOUrjji0iR7BzLgd7JQEqp/r8AwSTP49PRZgpf++pqzR3
0BBM65q7dRqDpdUbP6OyQh6gBD/z72eVG0uL6RzliNznMBvDWDqAr6kyc9NekKlUiJ14qO4qo7Go
I1ek66di1djW76vropgTfvZtdE0Fey+kEdv2sdPyqba2J8WwK1ocbXKiMVpn75hIIBG9omd7GQt0
qgKpHbIEd/QQ90HW9uDhHrfxp6yHkUof57wg8bijgzWMDRnJFcCkKOLjPvyeNGppaA19XN+7MyIO
Kj8LhKrGV0j68gaM9rlU1rajX1QPrWL2GMWkNtjgxL1cuFDv90eSz+G4fGT8WxtZd58Qv9i4uyza
otsEgsCAZczoJHyPQXRMLaBKRaQxycwCQeiblBLXRMfjIeoTSgDSiWCtYtkcQpG9J6x3+wZd1Usa
B10R0wGfWBZXWe1E1JzHWUP5PtUGvGYs1GpMX1Mt8oksy3M7l3vmOuxB3/5wpqSrnmyaLFlddQWk
HtS9VrMD7NgF8QqDf3wFA7RPLiRIGiaK6JToQ7RpdJJ6c+sKOB1KbzOCVRoZmeZTrJyiXZsq3Bim
uONZ3QWqkassjI3K+j5Il5Sgk8NNCTXKrOmwtToY+sqJQfL4g8wevIrUwcbxgHzckgDyH+yfAFry
goKlMD7pjv7piBQxKIKASb4Tcn0wFn2eogEcnmgIjrO88HACmE7kFangozJsSSYbRm2MtYoexqSl
ahi5oEsL79A92uqpbpiFsPwa8x2wLmfhf/tRT6hywQ1BeoNsUL7qlcOIENRtF+svB2EgcvCamblC
DAFgt9p3pBmObAGdpvgfOChAsnQxx7Ggi3VI9vZTXJJ3lpA9vwDfeBVfSNeUc22TCmmynvNz7835
J0R2ovf2O/6jhZwguC0/uHQldWyPecpe5jFipBeMiywUw0cepYf36ZOuMHJSajoCS7+zCTQiWrcs
PMVRWGjHmKmcRkwZiehzVMuf0vrDSwADFPVPq8ClueMlzjkUKxh48Do0wEGmogesGjAMRwZeB1sO
kPw13dj1uRtmjHqpdUmFLhT5TG4L1s+7oBG2+Pa9gfHvGVBjBa8s3/60LsR9/SDpf065xpSLSgQB
pjoLDCgxFn6oCFMkjD8qK4D4bjgzA/5xirof/f/NgjzzR4D56AB9a+/4oi1WC9RNZrQ5YoBCKLtm
Qgi0jEmCvoEzAZ5wT+yqUmZlN0ZgGOW+O+J9K8v11jtvprxEP/Ikx+M1Lrl8gdYZLJP0qFy4lV1A
FbvwakBDtnKXLdoGRUOp/kWGCcCIjRRhCACX1l0mJof5gjST+ux/RGeUjWXOAcNm0qxPX0rv1W1k
W4ufhD/w9IavOj1SsRR6yM3NFkODYDmtllV6fcj51ki+2m3PDTFmL99EvPGBqSgM0AlpBWGDUiGS
x+H3BxAXjPp8HO0kPjOdOw1uq5N/AmTdw6fZeEbpRpILxmnBBu3fQEvII1Zz00BpS73VyTywp6BP
/+24f1ZOot+nnLTq8aNWyJEShAKbjKD27Vyy1a8IuvV2BxcoYwzvfc3SBuNtqaXGyZ9EOXGnl+jm
IIYhgZ5d5/o2ziDDmHrU2Z8RhXkpUuAXvT5d99oKUGUG7qeoATLGHXeZ/bCVbmmzdU3M9+7m/FZx
PTMKH1XieVVvlEMvy2amarWHAhWtC/V7h5kD3hiX9Ym96+2P9Ez+ubHDHA+PZAy0YMmqYChuM1zk
V9GEecgqNfIRFav8T4agRRmt6rkMwsINQKEfkaAXtYjOwWLG3bJEncO5283Gvc8ICKdRlxz2Br6u
zpFlWIrxl7yUT9hsM9PDlzM4C/jCKkLBGpRrsZGrwtsfjpq4UUqVL8AEnbtqDv6LcCwevnSLdxh6
C0Mq/7Xqwd706ykE/e/zYxBkeJB3FCg9PXigs8bzeLhKsYJK6TQVtP6MPP/eJEZdufbMpsPyhrHY
ukzJ5vpfuq3WRGln8prh++doGgxTr/wroO9yYdkaOBFeJvZboJoJ8N0/anmQA8miIswW6/sAuCfO
NdH8/5T9utRnOG6azBXX/lmuC5UVhqucrfTyvEuV3glZ7zPF/6W+4ytAdZIAxVAwAYvfyriYvaIC
2WCrm3yXH5QSyeX5AoFPlkxb0dfTNPRUzEcT44qG/Nt8gD7ZoOU4UI38ux86SnYrZdl8UnrnnlVR
PXL/JhbKjofr1eUy2m7AP9jrm1SAlHQNbzsgMqNJzLw6qPPsbd+iiSUnAmfZ1/skNlK8V1p49OUX
Sn/HgF5JSriEMVnMxHqoP+Mv0aJMWgtajYDbwmNC/zq7En8fJ+3rIjczh/ZeB0Q0MlI263y4sgw0
IfXfGoIvTsJZQWdOkjXdZTS36i8FOG4mX4UOZ3q3jsZ2K6aiVd6khTYrGFKLvnF6brpnkUMPSxD+
FbO7wCV84NbhY7Du/R18jx+upYhBo05qFq3THymBr5RcdLlBWIpd3piwuC6kJ2LuuHvNPfPdaD+A
/Y9U7MB8c6XGg0o/QbFRyOzS4nLrx1xdpnu1JjN/hUh6oeYHQGGtPDpug2yyeetOJna8oOkMQnxe
YADfMW+mLhRngDqUuWWyGQNAO9VsIcCx0WhFABc5eqL0740so3VwiXmwZLBxyHJg0Mhr0I17XxMB
cWTmQ3Z0V8Uadsc2VSvPauhRX2E7HvGh2qyTYojx0B6RyNL1tVEHdkejQPP+2ybHFQqXQslCA3rk
GI2ook3uMyFSYO1Ex2zOQE0uVT74+8M/Z1grwnzsnuOfYhQZGJTGIgAaNnVi418tcIvMWYhY80Vo
01xJVsLdNxskGjBC40KkZOkmH+hiMCgy+nS4M9Fv1YmV1gzzWzRexqHaqV4Kq+ONFH3ZG8PTzQrP
suHtPfW/CAYFcb8XyVcC556YmEWinrUjwyzyfkA0pzAFlcJuEQH911gDjWnOASeDnON7+wB6wFi4
a/eXdPFOrVYwnUDk3LiEiQfOKmNZTWr/h2jNtJgB/JgCx1YsHp8lgBjTBK1lDKkxqePilAygujzJ
aA6jf3CB6zsGAkrhfmy8jLob3Ogg67qGRCspVT39lIYFxZT0WYL00wNbPVFiegbtIPWRtMmWOS0B
oTgVEBxQcN1J7aLAeFkr6hyE5JlirfhkuEqDvSXS6etrIqT+aJEN4NxPvNTliyPd+jsyqkG2K+hB
8mfhWZtCM0SfY00iL5s0KjuLE4EHScoBOSnx9ZQJfcqSdhKQ82LOtIFr/9bpDmwUiwOw2Qvbr3vl
jOxSRalfmWH/Jq+SnLDTv0UWcNcFspX78PFAvgt86gH7CMIzPDfFyv5GixiA9hCJNkCAquTpeW4H
PG6jCJp2rzUwkJ6WEeTtInj4WJKBk2bPb5wDKWDCPUBk81KsFYcGAoJRQDN2R4BjHnMLRHEWXP50
+FujYwKU4hzn/4J2/u50RsgKt69IZh/t50jzbYJF/yT9mmxyklPN3m0064miIRqCycQCQUkCG9/x
zipOhYLUFv0p3LbCxPktWjjxHRPyk3Xpu6QYF8rp/O5W7bT+Ri3Xgcjt7i9KYWJQ2a+BgUj0GELT
C4F51N795xZr4HqbDafOGIlOw4CGco3TShBMW7GlldIXbsD+DBxQ6bTT0DF+W9TpRMCpZtsazbDV
YjfnkBMI/qBcaM7Br+GBfzRIWKF+WDdTfFNPZMmFVQN3ZNvgH3azUs26ol+V0EQjsJiF5VvhlBas
iF6ltO2ZoTBJFj1SVOojZPkl+0Gok+tJJTCdWBZYb8RzvTd/ovlatfbinJXKlXyO0iemSOzKxyid
1UMCtXqjSzUSwcebMAQvJUzPLs6/Y/Ol0INJOrpaTiHUFU9/WMJ7fRvS3OnQjwAA7tPTMAuhciIX
5Kbn4QKV49Ac/dI3GUAxdmNDSGVrJzpi5Xlbvl89JLE4evVYb41SMLQW2vcyPtmvylpFEsxlsneN
27XQhbAR3qLQIsAAljOtvHp7/j4IELsSJAFdhcoYHI1t/ypaYI4d5BmMnJRBlOYIWG+t/iE41O98
u928BzrNL9vYFSAtRt+l6YpsWtr/CUIIlYwh2EHZ3NsblOfl0EbFQ4YYX72JTJtIpC/vf5YSoo12
0DdIkZ9wHlOe+yJC3a6jTsYPs9mj2+ux7X2QwW56I03nXGDTKDGWlNHUVUatylT+vp0+TDoPwLzi
utrO9kLU8e1fN6T9545oCPmuJNFTHNcnFm6oHphGaifOvCza8Op9IW57sZlCuwq6PS0eo1fACW1u
LIuqzJ2DUTDBbzvbwQohwpJUfd+LlZWxx3JbsIM7VfNde+yTcPfDKlXIq57uQDOUKB3Ylt+MY9MB
+y5U5hdP9wP3rvmKfCxMWH2h+7ghlNb+533pzReJxAjeLZuudp2ZTrI77uAOvOQLY66nCV0ho9Vx
xfJvvM51LsG/cM6hqTJxxqbJZbPZ1ciDL3gHJRpZTBSpWLcT6UPdNpDVfcdCIZA+7DY5JoZTKOEZ
b1uQgPuc1TI0ii8lzG/IBvuWRrXQ2SrmlYCGJ727M8b8ZB1At/fu3vCBmwTprS1ouvQ2kA8YXTs+
qVdQO6aFMEGMXwDw+CJK1i6kN6FQJFY5CUgXHAA72f+5iPx/y99caGQliJDObW1GAltptOT4+tsB
2Wd8741OgS9QrSeF/c+kW3oZ69ET3/LonXtLXCyQOkkDXWZDC1DQjRSn4xkxV/hF5Su77VcDPBT3
F5uG17CZk0Jd6paiK3OQFAosLv3fctF2XZ4VTDpr33nTIUN5wf5vQ1fAmULu85pau9Hjh51v4wti
HS16adL4gvVFW4X3cWQjxVvtys1lxtf7YAKgu5w1GTSascohKCg0zVtieEVuMmdW+Lfl6XYnz9b9
mSedf61s9V+vWuJbWCi7QqRvuf5RMq+rMZO0VrM77r2Z75Az++2nsEdTWmGuxt7wN8rzWyrutU4o
hgrrkitgLNRiH2eB+Um9pZwuGzpeM8ZCd2ldIjXJ05moEd9VLCGLPKQIS/rRFnIqBPXaSjeXuXQE
GUANxakAprxIeAGrrpsOwE+D3puIAS5/MtMvfZRVRzEH11f/gvvU27fytYi6UI3BrMVKbfGv6Dbz
7tIPedhhQTl7MYXyqN+wAb9m3tgXJ7USyNSq3PV2v8AWnZIsyz+IUZNsgkcTiSfYMaETSM6HDzQu
wpwPwy6YNcH6KHcWhQlS+F7UNWwhyQTaauIT5CQY60oTG72hZhwBSKk20qZad0N44iyGbffm10Tb
0exeaZwkNZpvT1ZCtuh5AIlTV1hv1G1qOCe9JQwsxZpbEAlEOsxOaEgWzG6cdWUeO1YnScHXTqw8
2lzssgAjNBv2IqfHmM8T5yoqHWYW8ef3QkT0BkmC4WurkYMsdoynmHV5X9raGnHuw5km4PGn2yix
/1XWK8ivsd2XnvSyvY83Cckehok3/L1PI/rjiYtVn5AK6Lj5LXKj+E+ho9hWgylphvcEknLBMgN3
CyNMmBrnxh+gbm6/Ff8XZfq1C06rb6qUr7lMuMqQTokG6mxoB5Lun7adTQF6LiSte9LDkwRYTiWR
YDUM6qNVYSJCXnPqua5FlmmAmEJG+OQsQHh/aCiGiYEfWa8x9RnX52Df8eo1NQIlgEGnbvZMgyrY
EerCSs5R3tFQjF2p+8NdDU9KkGfyXsR32nd1x8neYD9TCojE5a9mh/qhOQzlAvUlbquk+F+NIrkF
sx5L497VMwoyCtgDkbf7N0pgKt7VAY/T6DW2B8aUxhOZvHJludaPA/cwWG5T4giPgX6uLNRFJsLT
FyEogxRboeQmeYgrzdVaHPM9wT/DBjxSEeLatJnNyU3cxaprG30rXwFd1AA+h3H6m1Lpt7IeMyWF
p3nrC4yfaEYroNNqxu8cnmOg0oTzaQydx4nob6HEAp09kQmmi/HAwObhE4vN+4ZCrIm8fw/iaKXB
mmJbAz4txMh6r/yGWyGJdR9toYk5/+oBsIOlUuXaZLcgixDbGzdlHVsiDYoE7wlLIxF7CtgpiD/v
ZTx7ojdvbAhW8O2mf4f3Arm79XYWLGqp9uLEeKLK48KQq4ovmPS6HcXwT72uvAItr/47SssysQPa
ynA09l6xthutVQ2Oncu0PwD4kE6lIBO/3PiF+N1qy57g/OdQYqfjtlJCx88Xvemw7hRXm4tRt5W3
QmfTfYquViKxurBsNsWKYh9jqFHeAaAmcwvewnhoV5EQC7CndFEsOIEenjfcDBwlyloQ2oSoec1G
B20JtRevYLgVheKwmiHoGJ4jlPdOQYJ0y23ZNi7Hc45i1MIusvIgDdb+MPImUyaDEXP3oG4J3fHM
tGvd7X7AazjydP7gYH0kmiabRAUSWdi2g75hwqoYcEPAM/6Fh4ZDxajiiTrOM2AWrDNzp8Dwj4B9
d2mT0c4NnegccEG/ESvQ+Ug9mjMe/eIqG3qs83iaHLOh/y7wmZl9eo38/XOrcYpUqGZJ4k5PiKoS
6aXmgUscrkM/7V6Pc22q+jk1x6C+VRQtdXWDcAmLDOJG1q24oRcRq9wXceP4lp5MlPLJSwv79Kp9
fEEVBe6pACrInhSFKd8aWgwfvhOkoX2nVGX926UyN2t6Q733G1r3Pnd0niQG9vDymIYHqdygb0wb
lwEaEsywH7gJHKneWzp6GP6FPFrMpPmOUo3B9LeVEDOQ3BfBJylve2UvR73ppEk4IVNKZ7wA/PyR
iuyFtybVAgDuZfeDxov0Xbz9CfhphP3OvPtt/U+TbBBHE8ZC+POi3DpPQc3Ciy3kzlv71y+HqTE9
dYhA3I1PAmr4I573/Y84zX+4KQAGYX+FhiXZTvW8PU15WyjiknCjdL2aX5vkqruuPh7gINY5QvO7
ImoItGBQpo8akqdTFQajAnR4CRWkjLlC/VOghEiavnjQ0hmMDmism6HGe2GyobQe1v9hXu0/ybSl
y5YimOjoyFC+uU6EyC2Jn/2LF0JagvfcJsyUwP980k8Hclu8X+rI9lJymrF7opEt29sPtXp3sM/S
N1SzJunPPdDrrpSWhiYoJTHjOGunDWOxe8+6FzvRIXYs/fjOE7+tm5WJCWS7p+z4084kKbzpkb+T
UYk3q/1o0/PYvF73QOgLT1A0ONMiXDXh2fQzTdj/Itq4kIStgPj3HtckhyenrUdyZKXl6Px9jv0c
MuurSChgr9UscXL+DhVtkdUawEjj8luvveO+SSwF+iBPm8G+JrsfadX+qMkpWrtiiUxvswlPz17d
jKpqdpwFKPIPI1rpcENrijyChJifIWwEwyFH8t3IqHu9NNqZsQIyzvXWxXGQDKOKckrMLb0l3SH9
U2Yd9AnKF7NJSN6/r7jk7qmKLBSckS+ZF93k0+VW4UEPbaYBVpfNLNPnL52XSdJRXJ5FEAWRKN/Q
Qupi8TqW4OuQ/gLjZ5yA7ellplcEuZbRWmrAJ8j7YmfJzFAmpGUGdVM2laub+kQSCBoc1MNd7t8Q
dW6qc7iG3W0JYtloqHGcI9oTO4b9llnHgVmoMJXJVrTx6fkbcjIipsfLeyUlDyyRZbKxAWh5uZTD
Chu5vdp1TeZhr67e0gKDjxTvti/Yh6TEjUtu5wIEwDmpZLQ9oaJZEYDk46WNN+DMbT1U0850cwo+
04+5TbEDNgysiDDYVh4mv7TX69tOjdsH3AZuZVwXcKMT7YG9VWFbpr427UJ4bRKZhEhdKsuJ9Uqe
TvOtUEADycV+8ozDP2KccN5eSTWKRa6oXlePr4ewUVcp4PN9HFQ2mgqnKboz+jfuJSj3gYQvdjO7
j63/6ulIIEC7pMmbYpZYj7XUYPzXaBAoHUGwkGW4PayH3hvKcWTPJcOzR8p/cSkqcXyzjcJT+S87
INzY6lYQi0hurQdf6ZabtT1Sm5kdtnVEpfsXrxLcCp0mNygbP4YcpDegYU1jTddEfYzS/mV+AMSn
PrZvU09/8lFLj8LxgePeTMC/Xs9urdAY5QE+WlSJ/yGorCLUDKdZANtbZ3f6juBzdu9RACjvabv4
CFS3fYZiEMggtZgIDaqyuEIoVzPVIpfnorHXHzIlYt2IWahIL8JHhJU81YcDFzmYIr1Om16RjU0q
6Vh7T0IO3B8uJxlxlFXePLQNdGk0l2AYye639BugUH+LpCLbPdkvsKKVkG4PmEB6JpEBayX0E2cG
/I1cwYL4y/fjLvbmeTh1WZAboT//P1vD/SUQtq+QZykJZRWjrfWYHHq+fCcJBLa6qQqeNkTDZn4o
KnXRH8M+VgiHEQJYqXFmOrx9sf59/2O7jd/26AqLvGQW1wAwTo1r5yTHqwDm7k2hH+fBP9ZtasrP
zPd1ta0f9h+PZjgakDfl6Iws5imR+OusabD3iOBeZWLMJItgXWi5XSjBsNj8UGmNCkE5BGTce/xQ
QUP+iuwC3YXeFCm/AfjVeEqPCS/SIln2Jhdk+FGJSqdveXTb8mlFIdUAA6cEqvwB1vQWzfVDAsd4
bT0Sk9e287V1CcIIrVvgZ/h1q/Roqrhyx/Dr+rtXryyst2TQQmpk5oNyvHYy1AdSR4ePpAc9oFgs
yLNINOqYQTI0h0DaO8eHniTPxw9qyTfKNbC+OYuLd29yRRUF3j5E6Db6pCoO+7xGQ2hnzyx2eel+
Bqzc0B6jWXeknSA2zxtYUkNoBWly4a8AR6vbyvaxtVqdhEOGHsA2H8YXjrEVwNBzOMQIZmGQQkHg
fSBXhP2zHDXFmWvC3PzThLQkKmnhMQjdLeHh2srRObyr4QFKtbhnGKah2nYN7at+TRolhFw+Oh0q
H6/UGVbpiW4lLqAh1ZTL/1pvFN04xOEmLjimIhJIPltjVFr58HGny3h55gvB8CPleT37r7rQooIe
rQj66vM2dp/4+9hEGN5pwrQlYJfwOgmpeTRM/iVqQWnysTkPxWaKZ+2SJvPbfId4pg1/rQjaFeLr
xJ8YzliXibaE/fCRHXAUVzjyJgldc84Q1fhOBSAbVxpykd8DltL7hJtFF8wDSQKR4tGrUh/+apX4
9VSA1m36lWGncIIV2kepOafTnFqRpByEZKYnFoGTDdsJePo8E8tHdc9OikDVZnpzL6vzlAJv+lXi
GTGHCBUbKgBsEqH2U8aExTppoW344BrfewqzeeIDLuM1ZWxiDH5OLV1KOLLZR32dlbrATO8BGQ92
jJsWRHBIWI/eO5VykyirS6G5d7kTuAsU3YPVwkr0LIY1Fv8gJUUzt+NBFAURvmeBB6yZPZqUpGy8
HRt7+43rqsUT5V6X7k7g27vFcrZg8OiCV34h5oF0/y7PpZ9eRWCj/g2A+pBaiBIqIespl0KlNP+i
bN98mHFneH20eDdBDH0eljy9LklJ8xanILXF4LufpnkwbqccXaCOSi7ouwBl30556qnwqJaaV94s
WTrAqStUMqz8N4fkulR7ytem0Y1Y8cddQo/7iy058kcvrF7a2k+YGZPq8gLTSR1PQBOo7KzGsLwl
An38UHZH+rCgwdo8q56THAazzl/yPYW+CM7/V1zgvpD4qALT1BFEyvGjtBxR7wgbegpwVfBLg/0M
r9qtdZYWrr00SB1G8jpt0zDQrAflj3P8FPhRQmPhdVC6FfCYg0BKeAV65qQViLForZExNsfpvJso
v0WnGs8M1J1/Qj+/wL83Y+H61bXBVIPBVDDTDEKVsofdjuapY8PY+W2U7V5Dn+r6G89C9lAW5Zo3
V0MeWU7UpUyQfD9qnKTZ0zqVdgKvDmwl7X4DuLlmrLJzQ4WcXUOS/viu9SFyJrxmnUw5eXnsgMsv
1zshaO6wok93vqUIg+cEPDgVdH8JYB36iNFiONaLVvauWTTCqDrwl9oUIOg2C3dqTMltrKxQn6is
ZO1vw0x+ldJsN+DXuE/zWfHsb7tZsH0EHNS66O2xM/THxvYHdpFeV7coS1xXjD/+c6lhGA0W5UZb
L4Mt2RkGRpAHIVqakM97n7Hy8Xkw0Hd8xTOh19Q398xtjCiw6CasGZm1ZIbVLMwAaUlS+gW+qYEc
pb+QbS+nALfsTbz9Gqrj6M+MnADTvcgnPhAndezlHopY9uyU55WhXKhmg5C/0ZL879Jpjhu15r4G
BjI3iMTqDaMRdrwRFqM5x1eIB33ADc6eiQvq8j+INGmEWW6XM2H6/sjpiFfae1YipRRbk0wXVR1K
Xk8WfMARPmsPwDbBwfJtyp3CfvH0Tk4vP9utUT3Kahui9FAyVwrrXXU24QsurWrFdjLBChBc5nf3
i4EpQSDKV9WaQCWQcH4WqxWN3C3gy1rFiBk4xGswJ8h6fjHHHJsMu/GBrV7DDJCAtGAf8OlgGfaF
cGwbdMwEMvOc07kE0tScLrO74dLtb10zNivzfs4uQ1dsGcL2TpmrG9ssX2Noc2qGfPKh5vY/kZ5y
yriq5OvaPKqtR3occwSwC80rkdYK6X9dHgDDkvRvXwQ0HfgKC1VhjnqByQ2LdMCpKGBSgPxJAkki
QfLc8EY3DCVOYeT53rt3/lC11jzQiBbduO968cjQIIFtTWaDOT8OXcEcnCK5ntDwbnZ1Z+kC3B1w
zo/M5POX84DrPt6Hfs+Lh/OG2htK4+0Rgt+qvwK6cyNQ5n92Mbo8of0d4GvXQydCA+fnN8l/J6tC
vo3lerKnIxP39KMQwAU+kDp0rej3TZf25fOautEapFytUQwZsLnbz1BSYBfhI/ugV/9BTozR6eId
wcZ/yqfRKXHBemA5Rgpe9SzZM6ktfQIUCGYHnZWaZQFOoZJG5LlsY28ZU1BzS3JPXtcISk5VK5ud
EkY1bBJ4ztkgO7Q/MgTp7VXj2md6qrTpoq5gUqgNiYm3az7Ths8Y4DcnLfG/ESmgynmxO7BhSFhF
pOb45FEevGRaPyYwyVlWp5cDHw3ECPWf0hPhYvDzV/Mc9dxUkThlnu42VhLshkQ8VN6yyyq524Ez
AKvdEyK/ykf/6z97q9PrstIhun5ZX8BHFsJTfsCrdE+Ah5zpEgfkiPMYJXx9/sDfT6sC2X1H58aS
QYoEtHXzLqR9o0Pde5W38hW5G8PLYIA1hT9nR/t7v6h7KQB1sZrSh6wZqWoUQ6DRMxq9I6B4Hwhf
H3BgML2726MzEdtkOr2ViYjwssT8hL1x1pU/heL7Wg8p98FbwTSAmycsSJbe3xwDEadQHtB8UDtt
+iupBZqSrYBYax4HDBWKG97e4xmHC9JdvksXCzqDy69mmbBDgg0oK4NHKBEwWjGE88TkU3EO0Wse
mJ45ijV7r3cyYE1qWWzNys+thbwJt2nYLxtXoZrvLmx+rK0+7UhBIN0xV9O6W0t4a0xyvM5ukQuH
ev71Q6nTpsjuwYuN67mlteNYL2htDc4xa+XycPk0Y4ea80d30u0mzARpViOB6AB44z7KLAd+kTkw
7Gy81dNuWSuNYyWXW70ST5gcvMfIQA56ZT9zucg52uRa3grdx8TZ7KNHXc7/6haiUWEzZX5CmLjg
cYTIXCmKl1p9DdyhEN75fgYec0gYFU+leSKB+DPFD3ieuUPvArvlD9FIevbVp6ZaXRF86Q1Sk1sK
WX1+rPK1bUITzKg/FguNdbX/6rhllWGloxXuSPS+WWirfS9G3h91oAbWAzq1V1DdYDGyFdk6CeSp
vZ39T8g1Jf/KB5ASv6TQDA4LZAYFMXvxJ/teFo58ct+QjawG3sQSOt/dBnFO328oyh6yMx1HfyoY
TYZSEwNcn0B8JXBa3orq5g7hMs4JMjAYmoTj/jQN9K0aHBj+sTGywWdZnJZ2a5iFVQ2kjdNd0fe6
arJQ25ZZTRLxTcjDnGlesXXPn3X+c9C2MD9fMHgq//kWrEeMHluBWmR45iM+RA2VUu97sSYO61Bw
3xry+T4dxUEpHvxrob6N1aQb4G1mBjc+yUS4emcO8vkn4fy8fZYBwN4N364CPElvM5tiaLEIQYNe
Vil0GVLdu0+NJ1ZjGNyKlVMxr5mtGTuU9lw58Zm+yAJl3PuoW/267eyYr45fhqFJk9ATQiIXVB5m
+comJnpiAUGMTA/2AHozy9Kg+YaG3ngs2pRyaSuc2srYh63naBfhqBQ7e6fgS8thO6JH5NySueUE
0k1paizlVFUznKcg8g6dutMXs9hUdWkG1Pvnvou/RUP+fr1XgMpN2ZRoIobS2KMp9IR+QFphYmLe
bCF3vHcVfWqVnSLaTg5/pZrWKN4d4ytDjDkfAlx5xdDUzmWTKZm9+IsNkUlneJJHhmiDf2fxVk2V
7YPyhfckUvkvPp2+7elzb16vSH1wBki3De6aZpePpefsIIVdeSMsPMzjWwY4qeuXSjryA78FnK6b
K+GZgkdOZBg0U5JPEq0a5adhi49UoOOHBYR2VbOvzW2uw+9QGL5y0hCpPXOad7hQtlf9fO026RVx
7T+6fEjlrYzzvcSEtEBdOeHnMfHuW3XbOouXKZBf6c4mwlAv2b9JNM2t1fztOCxxEEZkus5Pt24w
8dIk6koSKn9kT8j682ur0ox3/EO3YKQ/Ifm7HfTlCBl2q9wpNID6Y+pq2FMf6eSaaTnk2EKRrXr5
Mv1JZiuVmoq7rcB1HJLnJvVKuYLeHePf/p2RuR02NHYGS9yOnKmWKPlF+Z3D9PdvEhGcsY6uCzJZ
x5soqy3zgNytKZYPbGIXJa1S+wjoihU5klWpjDhFvORuMcq8cNrfQZ/eqSKAnT+SRKlKzGvJVYj7
0ixKobXcm9DUsApwRtXQnINdjF2vHAJbv+7t04cb1CAstPE9YMsHhEmTd/9E462heBAIcCUzn10e
bn9aKjL4iQpj0ylb02/abeeO6NwXCSppzQ8Kw3avhmq0du4u23cmmuLcsDl0GHRf9DTViztUkX7m
8PWl1pm4Kg2v579KOppfM9TlFL3JERp0ZnZ3Nbk/+O85TSjgZ6BxhBAf6uMB09x4L3wpF0BtpYKr
8qFEdSG+ajD6VWF1FivoRlKmu7KvWxsir385ahX7GjvwyVqWB0BEBp/8qFslTgmL5M55+Z4/XzJW
y2qmn/9N2hhgdPea3+AOh7lO5ubYRkULcjPmRnnzH7hT7IHFF+x4ELtf2xiXKxpGspV10DHUQylY
iHIr4ZVQlLz8GvXkq87kF5Owhn26pJi8CZL6xqrxltptKQXGE1JiXqDVWLDU+lZuayqdefs3xdPq
LCNq3etuZz6l0vSZ/poigpRB2reB1QeQAc9Ms2KbaC+nUuEdNC4w8+hnW1vj0/nbMgb6cEjnSwpx
WfdZAd8T4zL7TCs2fSq33qF3/b0rlZwEJ/Jh0a+B+1ECc1RvRnOjUU5r5KIY/N8Ses80Gi48bQuV
4MF+j8S7EyI8whKiWr/YdfmucBmYNpFqF/XHFmFqtyTbMTMruG4X06Q7UFzJFy6qevN5+BGD+sKM
vN/NDlstShl3estySrxCl4w5FNSHwltLCDCv0nRM3FrAAFSVHA7mKO9TDPmy7ctDcFAc5lgHyEeQ
DwRaXYjVwR0+IXP85K6PXcV+KctI6jKECuppbu81EvL5RBdZ2K/3SXZANTNOA5Yi2ZtW7KVIqNLo
pwTagXbqXm+0u0h6fVqQe38XQw2PPhZORMnGXU9uONymATjJnQShpz/EzuWk0Ep1YXIsHX64sliP
zxxsFNykl8tVnHHsc6GJV6xw+sD7Ogfgmyv/QcPoNvxBWn+KlZPSlBlWeeBR0DrOTcMTD6z2zTZu
nb7AG3m7l/kVS7lKp7ig8WLbm18+wleDgPQ4QKO8tlionDOO3ttxWpQXtuJLv232liZgVkC12bUz
dVanKpVcs57Hjh2gXzjojQbxU8WR/XSYWfyr7Osl1W+ezM4mELa6gY2cmwNZkzeLb9KlQoW2b3zx
eOlB+pzPtcitahdGGQBb/wzLA0FUbwvKPB5FZjqOb98QwJVGZ8v6YI2NB/MURJj1WL/y5w5/GlDg
JS+aFxR+QU6o+XxHQqjNlCabTYiBFUnU4A27KSaaqD9WdrWn1VlVxxbPFtKsuCJETwES+7pFgYc6
rQppTFE/BY7c6h0Wj99Y4mpaUX51bMLrdlk4XMFm+5rVi6bA9ENK9ienF4nEdm5iwFrpxGRnDTDL
1m9Viil0wDwh+F6hFIXToMEWgMk8OemZlP0BvKu3t+1S8MQvd+WmQufUvXfUgAec+jvwzEra/yCx
jEU2/ezm8VuSZaDLrjEyTxah5eW/OwBu2EdTrRI0Tm1opRFBve0mwMHE87CVfW+fmEg6hEZ6Jl87
g+CsoYEKrvOVaUZzXZPLu+zAGc2tur5fHwO6ST7FYQUenclFxoIxAk7b6xZg0YbFfFb4NOwN4WH/
N2hq5fiQHcCxud206e7YTFvzjao51fNsaWPm1TVc02SzvGccGwYjqPEofXh91pfoZ1zOJqi0z7ja
coaXwF6qImeeWXDcFaM/jbqWUA8xPShGX5PdHJnrj21tPmclHHjdqfsw9XD4920tS5C9wEMcKaq+
NobZFDbiShUbSd/l3DllqcCgS5N3BQvHWYDRI14euAf4+wavQrao9z8h78T/2yEU8fcwidkTBp9y
VDLS/1b2+5cKtXHjanqUxUNTo6iULAWR86HcMtJGsPLYYKP8lJfpI/g5p+tOnMHUJhmoxLlKsb+q
48BgFKeenmFzRlpnZFI3GLbXdOSKwbF51O7a+s65QNeu4AvvZZ/HsW2rqsRSAoE/bR97TokgW3bd
nWXoOxIjJnLKvhKyXJkmcgD3wrm//GmGC9h82gyxHc39BtY0xr0CHmuRsQ6KMCHCu340ut3DHOCm
7KZxthowuK6rkZWI8XrNzlWXYL+GAgN+pbYoCE9KwEX8f+yNb6eXDUtLdpW1VOiV/fS+d63DtrZu
1mc+WN50UpiSGb8/juSoxK8K2Ws8PfqnKDaoGuw9Am+6hMR24cH4RMGs76j7shyqqLY9eX5TOJy8
pJ3JdQ0a8eNyxFyFjf5SlInCDvTQkEnIGKu+9mR2G5v4B43B7/vG07rmZ0QZMSwiv13dV+samdgi
SPFCi9gEFEDyZ5+X76xjQX9Pn7sSTEo1d2S/ScdBh0aWNa84LGczOsYW12D9BtSqeE7kkAQrkJ2I
KPKSL5GfDUsQh6DjF7sTPYCHi3IloiaOP12R56lt6JJGX+5O9cZ2SBbjtqumqxTnbAWvuESSQrOi
9KB/JqFTD/CZfS4wtmt5EShTiAKAQi1A5z5I0d+UolDlHQkgsKFal2ULqtev3r32PG/5hqHZA6ev
LPr4lkfAbkjiuP1Qr4d1z0r/T9I/vAiKI9LU4egtuWsKiFIMpgZxhHcblQWd84cbQ/8pv/84tyX3
7NTP4iDFZHgtOBgrXUCymhIskHdpfk6YJNk8bXDYVuYYHFN+2BiV+sxYxt6WeLdtj/lwDIqfF1mj
Mx1As8QQPuFhV5XVFmtu62kQ/f4M5C1vOSfRawdGQGpvAVf3Aiioji8tcpUy3V3g3Dbi1zQF0wk9
7Vs3sdHYErgBBCXU1G/TJdKf9zAxYm4ZpEAnFqq9Fu0LJDM+Al7932P0rzNm05FT2Y2BKV6OFUEy
9dIEyg+Q4ayrFPX0tcKozVFLj08t5Tg3BlPc/KYi3SBTWwph0XNjuUqvvuS5MVjI6s5u/1NFB/fO
3vFIIzsTBK2qwm1XMlRVc9uqhWH0bmyoxtC67659SaqZ9Nvln26RTNuJtuiAzbtknKDso8RvFjiR
bHxDd3Z/4U+5S19/R904HNIWQblQcm8bt3i7jaGWPccibkbK9iU3gr5WO760Skafpvr89t8tt2Nj
z6Z4lZLVzyUNIrX4QDCEhHMvpMvj49oyE//ytbGjJ0LgeNXUafIQ7VzOEiqI2vzNwD0knWecQ5S5
lQd4F17adXEZ6lJeLmXBX/tTAxN3OhFfo4wPkQ6VvS3mGhFp1vteCl2RE/F5p/MvncsoE2Q/G12q
5rbIVaehAHe1bhKAXwKHGW6SNda8mS/CtapsL6jXmiE1AKuSJ9EzyskJI49pQwX9sXIiLM7CXpBj
5HSwMjieOHXq84ZIYr+oaKvvkso5NoawXkXxCWsaN+B1VqsFZ5NxanfcNntCJLF6WczXTHqlTZNl
aqgNYaUDM723ZS2MSd2ZZ2PuMMXTf9B+6GIis+gBxJQ3t8WbaZ+sTuIHwmG6noUiwUf6omFLMIPz
rNHxJfEELRwsN2aw7GMvzuQsYy/uKzewNO4UAjEozFTK3BGenRZ+/p0sAa+WbUCXTrcrh2HF8KKG
1wlhsNYVKWpLeF/o2Tl7NUWN4wgdknQHrcULFisEmawEZg2iTRp2N8Yn1+jEWbLFTeu2Wv9UeIeg
rhfuLcYQpNpGsRLRrcUMAONcyO0/tHKeZh36lYkI/rAXomXi3FTft9WhGP8WCYKsXrbUub4TivLV
jlBQQkExxPpYatEZIh+4OARjmU6xaNsWH7v7qHuyAUjlWqezzyCFR7EBOx0k5cnF5nl0f9ayk5fu
YHVybxQ7B3bnxsR96ija+b7crojo0feoFXnE/1lobclT0AtC60gjfU7WqJQYQNmaKlXv/AgIVvsW
RJcnnW726ZxIoagNfNgELa70hP8n4cGGyOcF/Pf+aBNh+ihtTCV5XsylEnV+PDo9P0dvLMQ7Lzea
xjbr3csRxXqCdav6YK1/OYO8It3Z4r8HdWdZVstRzo6ICw24Dyn6QKKbAaLZjSqhgzCu92JFczHB
OhB0fbHYqJO5Rnaap9faw7+J7IWZDCKcmdqYaXjXqftc6qUZAj18EaxE1g6Cw40VBMxSa+E2HSRm
8zLdpfaGGJqDCqy1YExjaykyKUfG0fi+laaTGpq1Xv4iqrkf8/po6fBNeUCSPvQOFalTInXwlVxv
3ca/K/nAk9jkbEDBYDZpRr+ls3zu5I9vdszUGIN9/IKY7tXeDySaijExgEFxKvRNDF5ro6gm+TZm
2wcf9G27xULnQyhTdai9FGbOBRktF31ZNLkbffdTj2E2F7hOVTeIu/ozX59Nu12TSTPRKRkVcu1D
eKzjL9JV6ayD0aA6EKYiES0dGnNu7HZS1jhuy4xdoW91WTFMQrZkTOsDK5hRN9nMF9ZiRCiBsXOm
fshZ1z1Iknw0LGdtif4sI9JlYYm+cy2qt1ZebF+mpK+NMbA1a0kncE9yi6LLFH35ytqJrcdS79Ja
+WuUqM9d7lcGCLW7Yty4INsI5Ln+BakiJS3RdoyFK2k8ZAHcBBUIxPVBLeIUDxDrkH3pEqcmRFU4
NcDstSJYhuk5U5nZ+wkqhdN0Ez0w8H8sBp2kPoiRjHHGaV6bLUK2a72ySwIvcjbZ7ElQ/sbIJLUD
dAQtQZ+nFTlv9BmtbDXgUhS0VY4HWWYo7mh8vrSwJvtklf1hXBqUfvjMhgROqUzIu7qSZ6FXus+I
hEhf0F8D+idHYQEwX9aofW0InejVE/MUxwdty9SaHrGT9SWQu4NRD+4MSJ/CvxCTawbWa/xUfRCw
+YlhT6GaHCSSZfvcfo4VACB3nE3ojR/xRt8JA2LD3YbMBiQKbfLBBCjd/6B+caAgp0YLHwGLCBCG
zl5BuHbkRka/Mh5c410FU83uvRejDUyYXyA38dwW9dZgbzOQsQaRuEpbilAdbCQ4yRageYV9MrFM
C/teRj2hbD5qTly2Ej3jeGy1p/440Jkvr3ToDorki+fvZ+45wTbf/6clmO5iGWLAyFwcPVfEp9RK
go/grq/mA9BXVa666UCMxkdo0s59+A869E1ef7bxuO4ntv+ySAAyilxc8jeqx5yjobw7+8xMiQOW
SBiukoaA0rW7wGm/Jc2PAswqOOSRMoPUJ5kxc0cR8sM3o4bZN3rnIw7BV5Jd4g5kSuFbVwR/acf6
csI8Xab8dypXl2llUi49dnylEJgwVQW9eKRwbbo0sN98rikWGEsFHJ0ubu0FxLNH0m99Fktx46H5
SwZHreM2vlRfR31ElHDfFdVUXajrmTyPc9p4Xm/PZv6xh1MmtxVLzWZyeJbRFUU1y/IzzsCiAI/C
yW7fIY7yLCEhgpzt2lIYdjHTmHVzuZfOy3jPrEwdG4ozJVnFJOKsZHRNXLgRHnBMWrLdxQz6PtjY
HmDr2Tc1uKqGBrPFylQ8HupivHFqPmlYm33GHZUXmdA0xKUdv9BZRIV5PdIo2X/qH0hfGGPjEjI8
PXdvVCoyhYs5tYHYCfpFHQdc/MU1JBZUHtOiOfrNN3vonQSK0f+l4bCmibLMWjtoGBQzA+XCGWsG
6VzcjPbnyCjRxPposb40Hg3ePUAdxZ5PJ514iAT/Mo5U0gD+rUuapZ7OsbLcrZt3eLdzZpTopQuQ
LyV0mWhqW59Gr4lvRS8TSsXUmPs+0LypIM7KAVD4OJJHCbFWnzGrAmDcXKutArMfMpv49qMDhMua
ekmayDKBZvw4HXv6JzduQP+hUrp0Zya+QKuXKbnBgGTBXwnHy89j6JbSvu9jotJaQrWz4Nx4Z/kP
e5vD44D/OgMf8Ij5V2leIRWXW9+eJiog6hOzW9TapPL0xrSw9w+SkrDkU4MCoRMSwU18SpnmVUpr
dqx0GZPMPos9KMZ+h/pl+cjvT4aQkwyS6N/8OFixXbBtNH7xFhrBhpZ2wKVSExInorW3v9dFTLW2
iw4QMzSOPa+2+BIg7k/kdiSsMm5130x89bHA6DuVtcKAbQ0KjyQofIoHm+FTkD3f6FgeNhYGLmaU
+oEnynSKQQ7ZlcfzgS+0HbiZeYs3hMo9EE1yjE350+2NwYLsTBkAWG3JVY2ZfUsLL5vwu85VNveq
8ujcZ6J5wsvlnlVx/Z5ydI5PLXQsO01BE5fT0x/5ObybAkpnl767SoSVFQ70sK4acWNZfOQUtAC8
eNWZWbSMk5WS4RUsa8Z5Kz1oETVgZEOdBzAkz2SQ9Q8NQ+iTNLa9qb+Rk7cha0CuZOJkQS020aAi
cDJTU1/73O4XgcHiMCt3GT+QUkykrt9Ys0s4vHbOCuksb1yrJWWMXQmxvl1aLMO+22YjDvQPE36x
hvBLmsY+yudjECa+5FyF7RCqI3Q/rmIJb3yG9DKpXMT7pPuPfE63l4h4x3FrQctZnXBRcn36wMdd
8Xvt30Koqlt2udCX9ooekqmUGmTktlZOCTW99iQTMTmZ+dtqnOOOpBWplozm9qsekc6Fi4o33WH7
n45CGSl93ImUtnpWaEOvuh3Az82UAKuU+/nPyHc+rP4J+4tJuwyZ8azJWLBzEvL/xKARtgfbmOdn
otUPcgM5GN47CGqCqS+t7PpdYJGiQNZsSnG8AJLtLHKG7Oc5WVPlf3lEnx8lAtEErUc0NR52zBAh
tTol54K4AAle+nfMY7vqicaXpBWKprduMUUrEVtwxpO3I9hSglamFhaCOUNiPBwkBCPEkuj0J/GU
8A2ujWN0EeHWg/2c4Jat6XAfRrT6HnJlOEa3HVfgVkaXmG/9AeCG7ovO4UO15d/gsTWXqlFGYvmo
QDZvGtoOaHXCLNmmqeNZp6kphmfjqAHnvivp8pJy65d+2l7I0kmTyy4GZoEB0rg8IDPXfMDF5onY
Rn5ihcbBD3MfJLJZWkk2079vDDfsMpm62CZV9wgK9j4Zw1W2T2X9+nYrZmw/HyhCZdcCCdotDt08
vPxrlbmE+ctVEfrymRai0Sp6/qqfCcyTdufO50yEe6UCHD9PAhMBzo1d8aikbvfsv6mrxZarkWXx
Ur0z9f/MpqOjgw8K83u/Pn/aCuR/dvtwSWwzocBy8F6sP26vOeY9jC1IGLeEFj3A2Zlt7T3nRBzv
lg6l9Z7ccjlY975E2x/jtKjnITXF1LLbGV5cubTdtJlhseUEZAFG8NF6LcCVC2EETF1LfpAV+6Ik
HOWs/zmalWGkcXomeawfJ+C3BXW/gxOufjEvgetZQSGZ8X+g7wjGWkwJDcfQPMgV2xNZoDDdm2O9
vYQeL/gNou47gb+g7V0CIFmEECCl2xcAEkOtP5AWajUjzsOskXflYHifetxcOYFNgstG3xzp0ahB
k+Kd/xKO1bveOHwdiZV/w+JK3C3G0sQ/0cQIBr7WXjgFgR7ldMw3nv+sZ4PHJ7bxZ9OV6oGuP2nY
8gEyC/a2N4P+QJTTbZueUocKbvfu0Yc/k0QO/AcirgD/geXFb+7ybcEdRxu8nloUJPAmtqluW5Tm
MR5nxzR5HHSlByYxp9dxNYE6bwv4WDb5//dZJn+NKrZYMfu60sh32l1SLO2wEa3K2XbX45+Go18p
0K0rB10p8Ee2emYFPbcAIc1hj0VYnpak8YbVPBdSDlpsaJPqRtcfrY156/caZjGnsHPsGj471yO7
CR1+0CApc9hJ+/eoNxUqFRu2iWkrhDi1siF4TYk+I+74MTu4WNKNCOobEo5Jil85JFP6LxCKVxCb
0hxWOUx/n/IV+WtnldnY7NdtbeVIbl/ycGkXZlo0WSzm6Q3H/swwaNiHcm4OUibVi6rfX85/j0cC
bAZdq/uPSOaNkxSsdmn+baVIfU5zXfyT4me8jlrhuW3Vk8YTeP4oYTQwPl1Qd7k5LAl32EL1K1Nv
lk8ECjDRfNpdhCjmXMghyCr8v0eiglEhtrA94mI+HwH0eEw2P6HC7ah0OUkQ8rhbc03y/uUb/mxO
218L/K2sJl9Ne4zqi8vcV1J48gPO7Mb1sKb+cYhhKasfZV6ZVkdO79/fzYEQIMCBemjFSVY23SXB
U9pSrlFwrHgGIxC3Wkkc6RhBfgKKe91h1AAp3eDdrEywyhaemK5twnRyPbPvDjj9xUF+xFEAgrAX
CNWDYzmNBvhDoNnikiklhxdeWTUgLab0gYn5lBYsxwUtXP+FJxZNmw3KuNwoTWZ8jo49Kce8OP6g
IqDduq6zeI6yJIvgYFdf55zsF9N0JBBqAK/HXjjw2gClm4MGtwYma2JA8WJOXA3mNUINuaIM/5ay
rIpSdtwiqAfvMLdX1oz4Iqv+29CI1JzKICzj1w2YIW/SF5cusSYP0yJTvDwQJY3FK0mA6N92lZU7
BKOym2OiWKKN/7OCUWkRj80rvxceNG7xKToTKqqWUTm4sz6nGwsIMB8WPY3YPPoYMrh/vH5cjnsO
kWiveu4UuoDR9Dtayi5UyZyQA5D8N3evDqQHhsaAoO8UO2G+1nHKKk4RND+MFlSJe/XsroElSfib
Ks8LMB4e5MU1U43Rb9O9vMrgIl/k7GAl9GTCpRK2sl3/S3bxJr+M2Plp6XJ7gVOC1Um/h3LUx7d1
Ks9zyM+8Mzd6dlx62YiulfeacX58rzUFZcBo5nayMF41VxwlredQZu6N5ljMZ0Lf9ZMhMw1vwoKM
i4bpr/bkM1kD87Z2QESJwhSKSqzGryRQWP+g99Clef27jVLw3P+7hJHyyWMYQjEU9wydkMbbC3Ex
kfn656Jx+/91nOIZCbHgpa0ASwLNBAdf70i6nq9j1Cns8C1hRbX0YuwM/HJHFIhDMcp769iEbboQ
52snea2+cfOLXDdkq1VDQEHMR0iMLYltvWUH8NIZtVWE72eWOolwp75s8D99ipuAiq8A/yzKtOOg
i0REM+ZFp54LFMjIH/Yiht9TqrcSSIXv5fJVp+K7qc9k6OT4M/55CxUTYJDGsoYJO9M9G5cJN2VQ
NYY0UpPaBDbDs3yfWgmBqo9i3vXRtmyIwBMN78rvIZLzsyN70Ocybs/6cfpjbe5duITir88QIvIe
+jGuPYe+xBPaesWiLk0TwB6dId5lXD/fDdNZJWrs/YIJ1juzDctfSwcUPSpvrQxlxrCM9JkS98n1
5QVmFQgmOdXd7SJ4bcmdXt9n51hlby19zAWFIcuQNtTxU6lAN+CCG3cvVdzx0+oaKePA4IUx/DIE
cusFp85ciLyOSiPZSqsdDVkga0oLR08g3y8j7yWXDUCHt1sQksfc7s2gFlFH6dwHU+duBWZnlf+O
xsAnpLSf6GHUB7xt7XLbTxFCBh3fX9SYcdybBQNDYAK/b+HY22ZbNZtfQ/jm4a3/e16Q+HY0G4ZS
Dxjyx6N3a/ZzZQbeRXdpIBJMKeFG/4NQoUTYBlLKm7dnd2xPQjSALfI1t9QOOBglLt2a8h9mdj/x
ZXSvgir264YfFiUe/RgHxkhwxsuStWRXhQ8TWcabIf26BhsoqmZrp4I8KShjikLS9wQOWnIP59QK
GWLTzl1QiqLLRyNoRdRubvTtYY2bKtxAVJbpDJnVQzSIn86dvn+Ax2oXMOZgHhYgRajT/Lm7Pg8s
2jMWY5s91cMlRhAJQ482vEgY1m4VvzfIYZDf+dwHtMGVptdGFhrv8WkE+/bjol+0RLUq3OrwMy9X
Fb5JmhZotVBGarLHYZ81DD9m3/D0nop/jlr764OnTBB4tKF99jQZStkTwYEK4ymhLJxbh5jJhNoj
qF3pThVjVODmyg76LLMEFA2DjTG8EUs5kxoCdKUEXYuaML/vA3L2D7GqBg+/UfjfODn03g7ZvJqn
x9QIgYbKxPkNGEzVJDlQ0LgrYbKyZU0bRz4kMFH0aNi2oxiGp+yChqvRW+WniAcC0EsCVmOTvGVg
6+e/6q7PBR++ZIK5DF+BaUA/RhMEZDiRvn7/Dsi143yujfkp9eBLgq0mWAMBeKPyi+c6WiJ4tQNI
YvlEEjaLznscunzyQGLN2wLOK+LchPIChfWWqM+aDILgZpxhyCUJf5HXq0gXmIYIl5KAxgiKvkJY
rYpmdyqT277DrFkEITnsxjUyU9JNjXpZcs7XnvXougi3VWd98SKCJcZgjF3QW2PaQsUXDUWJxs9X
7RfN/Sw4+DzYSjSpVFukq6NA3LqfQOlgoNI7fF/tbzRIiOP2JThoYcSBd6AmJU+Nf3mGLOm7hXTz
clJcjjyR7wahYXEG4PIyKzd+xJ/2UxCQHaT9kpce+la6hF7DcuzIJrB66/n1DQdv3XFJifDQ7ph3
qHo4cnnFxQ1VweFpxZWYFAur+xau/uK0Lh8tmU6b7fefGqP3g0ln3oCTBn1PJMxJfnnDzZ9Kgj47
vYNVIt+ksExQoPe1cTNHlMSKyjlkGbpKkt88KGFmEQoM3vDlLDL9pJmoUwC5orrBH8BKoNwf/vWI
+JphtIXfyNJfAvcHwuC7zaa2IroGLjxzyFP+2I4rgRFtO1cvlmQRoNzXZig78qWLeaatAPWhIEb0
gWHQno6HTj1tcGwFK9vIl97dTXjyQkXRDFNZxV6V6dfj3IjI9p7cYzcXTF43Tn/E2AKhb4cfFXDK
hjfVvwuCh+GhQ4pZ42kVEMVWHD7Mi5SE7w4gy26BrO5OiY7IddAPPn5lj2oRyMeLOA+oB38+lI3O
Iqyz3pECsQ50HrsL971EJQ41Hox0aUmsrNJg7o5zQ50k5riL0JX5RTNI0XuBGARHMUekEixnRDvN
XbjuktfKHOAHEgCBEi8C1e7FT7sy4HNcFEEIAc5WLPDXUYdaMm/pyYNnmk+7sPKFMcxROytO4Z7m
Lq+QmEaoQlTZK5PEIF1xoXApa05RfTLqQh5IQiyByJ1G3qqeomv+XpsVaYEcKkv2sWcEC/vhyeRi
1mn8drRBzjiCaNqZ8Hm+94/dUf1HrEg6KPTdLWw+6C0EiLIFJ2O/s7ahmS9J3x1m6HKuZdl405oR
YZ4GMFShKv5dgwe+ay6fo8ng9ki88X8DJ4ikvUZCUtPrRcatqdRXibC+Qlf3pAR93NaaaxHgJyGa
X93SaT/t+ih7qDOLRlnpErPZT8QgxG4vf4fuPswqjtPbnw1loJBmLVMakankLDSrCBvIlQrAgLLe
lTKgyVNz9SneQCuqtd0d0ftvppuZjYjDbFKPSEys05lBstKowCyxhfaU3QyN51UOneqE1DeoPMRh
zG41KMCZMFgdhSurKz2ocTpo1lo7N1A9e2XAMCbNZKGoYSn/qvoQlFsex1kinmRygC6GTzaBGG0r
/5RfgJ7hQC1QOfzN9ZvLoSPh/H3R4pXQeVlXrNK5An0G8vW6wDcW8IXxbL8ykwIgvVF3xx65mklO
7OUquXU7HMZJ/Mo3KHAnUAPQndMZqgYpclA7kXXr3MjlPP7tBuXf7SSD5xn1PNT5NfdnqG7fOt6v
qol+yuj/AzJ5tjLamDspBmN/l8OljHfKmgn2iAjTS51fN/unPj5bgR8jTuxKWcrxm/q1olBLo50H
0NiPjU/tbC+C2EiNaXe6xzvE1mK6TeVUhpFws7b8EPyFLAY50NEhZ2K4DEKZ6YVzhlpfF4svK5af
C1zowMTHqrxbnIKwqdjJSC3t/RSYzh85tYzQl/NcyNndx2SL++btthsslqLtaA2r3tttdJIv3jxS
r66eibTABSG4wr+hMcG4pDt5EdKon805SVNDUfWMljDh+M2mglsAmP60QLvDM+t/FgXfqUvwIzzn
5QnSZw+BAEyVDPDBhXtQYhTCRpXoV21UbwpU3X5oaAwTN9cQyiA8mBNNDP0UfNpIwAK39MPHi4oS
2ksPBZygwCIOLP2dq/2TrENwO7UcBkqMokbWJd6+8/9ZNtLrXUSuAeMshnWVQ9BVu/niqOxQiCk0
6sltR3aaFzksjLZthfmRCPzS2Df4jqADRSY0mnGU/pw1Q7s+7ybzUEegYWLsWdlRFBq025iTXmVq
TVGGp0mC0RgSTcG4IagbXdFMrWhWkTnsUpPz24nJqx3RqblR4y8CxnTakLY7eFeGlFU721cAN0vT
LJ/k30na/8R6DfvwSXg34T3/6bZRypAn/MGvxXQWn+yX/T6ul5+5fdpkDRsZHUveGXjLpKp0TUmT
tvDZ1NXmYho1QJ+kavkNHVbD3tWwBLGH/pDBFiSwEVwysHtaeFJh6LyCYpQ5ZPIinV1B+1c9ySb/
qnW+1/mXlfHaam7Lu/nt4PqZIv2vgW4cP1ts1T8BN4CsaeoOPsLPWefZNUuxxy+Qz71aia7+u3/w
QQt16GFSYsUywSlS/zwImCz+jHy3sELpbFxE8uZbYcb8mpdcwOlm1GqhRNc5eOPap68vexbXhVGo
2QtsXRslMs9xQ8EEAXWlr4/MAoGhbTAlZ+va2b8v3zjrz3Ty4rAKh9B8EhtrAbeh9XgWsVAlixt/
TqWK3ZJrTNLX/49Z3Imkjs0q3BwvmTj3TxFli62FTn2Y8tzA7RPXcJbXyCPV1YPt8aP/6kM2ds6L
6mW9rWNC744lSdWLQeTq9IPIS8QCKWP6A2GcpXwMyPlQebWyNobzP3uMEx7ksF5L1r0a8YSGwgAe
F/TkSj5HPgm5IQnZEZuiPzTwNtweZk9Hk5XxAtLNsEeMMIUxkYDStrEYw7AClnYxci+D/tG8fmQi
zzpSXDoWpQinZW7gJKAZejEuzzfV5gfYodVWe2UpHYwWJRdj+P7zV7yraMSCIQ+yGwzNE0hjzmPj
D80gNmSAXv9xLEe/xhLn5ihOirVSlul3tGSr6/RCEJfQBdmlvULhiCT4aVaE7XKsUExfzLZvJKmC
8qWgZr55oEmQOmKeSDML3Hxqcpeaec4ljYHUp47OT9muUgeQreBpI8M2jn1Cp3eFmyF6U2Ehji9y
N5NbTVQoFcfm01XmE6NzLY2pU7q9mrzM0XRQwd9Bkdi3fjhOwBBdV5YaTJUk5DhooGziaGESYaj4
jMQSonzKiJ+AD/W9yP9LtsStszydrfHfZ7OZllxpjqvMEnCSbs7C2GWcmEXuQPu/zeLyXTJqObxE
LSferK84RsAE8ffaSitJQBi28KPLIDdVdLWs8r11BYP2DhISkwAPXgg+iHArQKfFZBtJYZH2lTXr
9qDQjzJqw5YqKmB+Do0Lz2auyy0FG4ummCfhuOytVIAExwRjkKhRXYUi26utHtnZNlwQ2yZSwdhB
W+L1iNn1z8vVecTv49t4G6aowIa3TxkI/Gcy0oi365B+M508XL/sIBLBIHLOW70b4diNQ6qerkco
CJcIfb8krx1BR0F5eNjuj7rPCTM/bX3pwyt0Ld/6W0bMEni9NCo7+3vF93110pIFRi0na2CnlEaz
icpywdFJ96MLgGrfESIB6LnQkxG16uz8K1E7iuWUMJBDEMUVDAX5CVEEUJu50Uq+JOl2zDu/f5S1
Fsu9r+bq0SKKVhPKx4g4IVVa3XZx9B8AvJeQwFCbL0IG2TCaTi85RVt5G91cIlDAtkj0Xfm3IQqx
x15lu7B7U5I8X8tJAgI3BULe8I6/QJmkoMWXEAEo0zIAPg0zz29FGQ1vCmRls9zEHb8IrMcCSycX
jtDRjU50DeisFYYbk0uqNS9LsaI3OQVPcvTNkrDmKeJNgzdEgLa76TcfRHlsLFQwqdiaARKbUoL8
zAqB28/EHWwRp4eVZTbmNjKQTAyn7AyMNTT6DGVKViBDqSXKVJ8zI4rjkOIIUIm9stVi0K8jx5Jv
8OSRNL9YQ5wAcDBvQeqS5cQ509hB1OGQFEGM2RDa+xnPmsfup2Dw9vcpp+M/ypF0tp3gkUrzdgF5
oTV3IZB58InbfNZbrxa0pU6O1tm1vgvrK9HCNRsIn9srkiIqb7cgWOiLy0gdFmU8sYe/HBREZbcB
rJf/9TzgjlO0rcP32zXLa8ySm8QoAi2pGNf/MZ2Nkh+Ze4+4PewsueX/gK6MX2t0p5VN46+BhH5B
TLYdfIvr5HMwU8paIDz1GJBreYaiy5i9vzpDGPdIWf8OAoINrqXB2nVZA8AhKvtFyUC2vmSUVY8H
9qk/4F9U8AvAW+EiQAI59UlZEPC9qLXEoQmx6LBwxuFJd5br10mpEGuhrrOaVXK44/QEfkRy7D1d
jSGA0NV2UhDL8sczAZy3OmBHjPiVEVY/a8HTNQND7dQUApUCuiQfCc3OGvXEGVoWIQvEYZH/UAyg
ahYDjkn9rJ7D5fdRoR1GBxHftntirnqlcxx3DfF4BqwlpF/slCDQBjuAbsLrZUpUhCkLeQJUy6J2
gGNeH2HY4B9p1lhtDGXHvQtRlWpdWMilm+KWvF8PuzqKMxO4I08bV0d8TwJSLFdCZONK6VpqPocQ
D4s4y3NuqcstpN7cc32hc6cgNcWxzsKk/g+9OZlNEP3RDJeUS/VSHkFW8IniaWv/ZlLifchKSTmR
bYC5a63i0k4lSn9XkWle4kxw6czO+peHHBpmOEUM15xvydeSvN4siZMt9jzxBphfC+O+LZlNlOa9
UPceEtKHSUCcWuEAu4LofKIwb+62BOcNzT+CnRGEii6PRsxXOaFb9tsVdNUCMj9Ye5BIc2XUf0Vp
maGWA2gljFNBqlVsJE2LCgog9J3IF8Y6YUhNrFKlXL8cIMPqCGgjSFlQ2Hs9KbKilaYURsh/Aduv
kjMrqHPobDQzbRMNwqnpmywClkWXUKit8FC3m9gMDELk0rpfd3rYeqH5aOY8VTl1Ya7olzfd0yoZ
DjfhpuB1HLCb11PwiplX24HKaY7t4bp79nTE4dPh3KaHE2lyXyaEL9xe1izeKbnzw5F5mpBAsZ6f
Q6RBxlPFiJ2ivxdC8/xCvo7z9iIQhu2t3F2tT8z7dTlwckVKPhX+L1UItdV3Ei1JgYLEeRMgFEbH
Na4Cga/oyOA6mm/pRFZGHz+s3hj9cHLy7xBcr6rZXKBIZ0M/S0TnzXrUF/WTLG4KAR5wlz34N8Rn
Xi4u5BORtlqYP2Qree95UscREBcRkxf73jnlaTF9YewsSEDYmM+EiKGP55qevExWt8yziwe4eTKJ
ygX1yCngxQZd70ta85x9vqReNR/b9A+CSWOxXyt+iyA7zz+40cx0jLhGa7HmIn6URQcfekmEC0cO
Y52Uz8dM9MdI1s6FAIYvlg6ZoFPz+CViIakGeZnEGOD6cy/3y7kwVsxex9mF3LHRlDBFEycefS7d
8ZXbkbASoKJnxEU/Zid1rAoOzys+akoS82ycdjjygF+EY0m/FzngfW+6yZ1olNevR1RAB/TRSQBV
spPF6kFqkQUiJ5F+XGtO1VGaoZ6uQggaMnrSXpsUqsQ0xi6JxMh2se6BwtFRnljIxwtFPol2zdY+
wKzoiDh9f7Rx3ICq+nk8lffzvzxqbPL+GQ5dxaBxTaV8QxhLy1TZQdNkd55R4FKA/3MuZj1fg8aU
xtOkbv2dGnnhikhzAoLoDAru0XZAZzZ/Q3LIu7sG1jSFkT8Wvi2/QJ1gxsb4FXkPzSV/tEHOQO34
3RxMId5uiMJ671+YHhGSHwcaTzROl7gfG0L+oZCoiddOywuGwvANQ/SNjnXNxkOmqjY+P06b9weZ
3domdfIDCSbRFgiv4etDxRoFFVfnh/233xQNTZzXwRZwj0zIJLtZnPpfhqZeOTVB1NA3PZ3Y/oFX
On6isy7RJ7QWJaxfChN5HYNM9gPUCPQ3LgmhDDRH6Llw9UtccdJpg/A9HevR4bNnMXViSlei1b4d
lt6qUnJm94JBSBd7AY7WQJ7HoIvVJKIveyX7hn3ywNU5m7Ht13XpMxNh1a9HZBZ045xAtTpFOeTE
9nsZUja6iguPLg+i0Ond0j9WKs4OMasR2RAktesTYohMiwhVvAHqQMwyKBLta4MRWxTv0tNSahMX
ARvn8Fu5zrZdP2MB0yhZ7sOHTQ7Wu9Kn+5UyukH9QdmNWLGdXMC/4+e4FTTV9Z03YbTXZrx3xQXA
mrnkMY8SC61jPNkT+FzFTbbDoSjPkvqsrcedBvvfUiH328as+idEAodzUAjdpQWspLWA8pT2XgCE
T84US4d0cijGgaMc2JUCmR6gTsX/hr2jpDMFnJLG5tdtwFGzJu7noPC83NzwChhWGcUxJUcUT3Mq
yt22jFtK768CEG22jcKGeIu9lo9AY/vGKXVgIQz26E5sVJLIADlxFbQcYXgkcdku/YQ7/S1ypdlr
AAzj4EQFj6J6WwGmjkv+CODqNgGdoA23o0ygFyjCPCbiQWNzLSw6fHAObu3UOeaQcudZwgknvixY
AxIOX16nfXuXl/2VGiNL6xAx11pYDCXB8U/zoEm1WNsS2LnLHCBNkbEpKQpz7MLYNlntImWmt4zy
cHRYu8JZzMiqmmae4u7npqBLUMxGHku5F5Q353Br1PYSFsIXpqyNZUP/04yhIN4xuATghC6BCDSJ
JThvtLhzW1FlQB1rRmLDTzgsjXf8S2ixz5lEAHImP1qe/7k0CybJ6d9vs/0h4LzXbL49q1TryzJS
s393D50TPQ0QQisNQjNZ9XOHAl2r4FulYGy81o3V1AyOwRpBDNkCooTvOmFI0GxFz9zMnLi2dLm5
IswxLtJof1TbwWievapoQBEMj9h5j8BQNGzn2B30kGqMY4KT2mCVB1bwr7Uv0yQI/36qx6WEKn5+
6sWZkqa1bfJqeLurzGGEYCGuG6bfYR6rZQU+1lwAJkqOaib+LMPzeyqvmDDN4vaZqPLTn2JAJJzP
3El2zq6dliAWuTbi9nLkRQsXFeoGevLuvCLME17YZY8w9tlnjh6/zZaz7XIwVFCvjdVXKYX4jxUg
f0/PKyP6M1EmhpZWrok+FcN0lmAGqsk50JUgEeYZEPsxykwa2Su5zEml9GABunl0VFAJitWQ4a/I
w6aqXjUEnSFkXjvqYZlA283I0/7sdacq7RIWDrjkX4OiAOO+PFFd00l6x1a96Egdr/IIkEeDaVX+
NCx5FZRPqeO2mPgtZWjLVX4G6CjwNLdbHvP8nv3NE80s5Jxna+/Hw6CGc6+9wIxihN5vUivhlfhO
/TxbEJfRBTIoXObG7zA0bQ5bHAC9pnI7Nzmf7WnvC1y3W6BVdr5BmHQ8BT4chjL1PUlFGln1DUjd
2uLUAj6SGMfDCg5OSWLTB1cgzqvwlj7Qi9ZiQrncaOjdDbImUu6C76YStTxgc8zV123a3d7XRII1
b+72/ZryGfpJcMufk7kx5zEhLOnB03lb0WeEGzx7GQJZEnCgP1hV7KJLqJEDiKMOkyYXsErwvC8F
POQgowmICF/QZ8yOG93nuOBYwIbnc89DAClCxtqgSKqF1fPavoitznJP80wlavPOuxHhDs6LcDJt
Qw6TPSpIX8D0yrVFj/qmkKcfLYItqaT2ZrjkIqXTTx94dkn5KjvmBORlVNUQaZ2tvNKFDsff5yqi
pcdsaL0nG69y4eDKCKx6EN8r+lLg1vu29od/2zbR8f6+I4e6QnQmNH7qnb6Zmoi6tGQWigxrjxgJ
psQNYkL0UVPGF9iiA6KOqrRYCErILMfwan4eTJhYtz030QLUZhAQK5j9UJz56/62vfGTpV9HCjLh
zNDBbTP0oCMgym1yTMxEcj3DO9Gt46I8Ez4CGQHMYTujouGKpk7jEEccSL5ejpspxQVicA3w/puX
ZbylLlRt27CmzvBkR9RMgH0kt2wv82EvrYYQD0cJmgc9AFt5xvpXFlj085SnSB9cAHB6JIzlLny1
+p3Plg9F+8kvW4pAEw/Xo0lAvn2BDjO8XqHmvERMqTGBeISteZcpDyl60Wv3QqVYO4HhbICSr3Fs
cXQD12evxO+cSljZlnsR9dcLN04CbbKea0PgdEgEL1Doq0ZfH8g2e27KBdV4Eu1OpYgTiSPjsYey
hUCv/uGHc4ZzOUDmw+01aa3anhQc3pIaXMBj/dRD5X7+DVz4ziDq1U6r4m4YjN8RfsTLeA1LjQnH
TrdzhRNRswhT0zU5OvqWmletNmwrS1SoD5RS5W+yrD+MRdf3HhjG6JWEysMUl1G2BMPAJ1KZsUv1
kibdZEAE8guCnMyj4ogcvRn0MbwiFLoVKnemYA1TNYRQFlU+k2MK4F6i6bgJ+2bfmCJ6p+7w52/A
v6Nv92HLEZ/55P9L7CsuOtwSHun9TgezCsfqjVF+IxdjYENh6PiRrwNgex8l5lG8hhuPXyg+3S8a
cqbWGFkpQDPSYIz2NRg2mrwNx2SBYms3l8EByhdyayZv5Ejozj33n8VkL6aO6aZWqDcvTjmE5Vrn
NYNEbR78pTiRWKYfM6QA/7IyHTzsE4Rtilx/sDMGVzPM1rN8uw2SAbDz23u7V2OCwMkD0ytIIbo+
MN07oD/Awt8lhAjC7EDdnxcwGG9GfpBuV8TwqA0l0F8fpGO26wR+kPFl44nVsTEBIpdDyBCBYTd7
TFh/23tDtS3Cq9R7id0wbFboieKapLnpaYov0wJaP2vATvcAZ2fLoqs9Q1U7HP2E5wcjqPB3gt3s
YutjxNcWpI1kiXV1Bw5tQJe9So6ly3nmIvuC5tiAubydCWOWBczHWxRUtyGeFGn3DKg/MRqU+97C
h+p0Ejkx8CuVXAYv1cnsoMDPgjXQ8z8RIJ8i2g9OJeAJhc7aGfebzt8vwAptf5iWHb1ZCwR/Vwxn
buqFbEZdFcsqGIlLJwxYghUeAj11a5o4sAPiBWZ2oUMuJC4jA9BZY6dyGrrBSWZb4w07nHMxJL3/
glVHJALIcS97dGrIhf9RkR+5xgrhFQrBHyDI/6PeuHrENpcRXCnwtv00fxpB1C2gWZHgQw9DCd4q
nOhr5FHkpO5khNt+ZaCoZTBtwVcLX+uEizx6jQ8hBBdAndwE1nyERImBOIC2rDC6/C8ZhxssxvTD
5rSIztCn/yDVyjsS/nG8JVToOfdLAYcClxkKEVgGCc5GmLfRWxQemtonkb87xSZNruoeo/zZcYUU
tKKuERGGHqWHtNb1m8SUG5nwKIynUZNC0OG3K3p3QVS00KOq5rSBNfhWRInaRXAgu601KHc6rsd0
oTsj3H9mR8htVsh1gxZ8FAiG+8ux1Siq12EQ8OQCH94LVgnA0CtIAVUapSoCLQZjCsEW4TW2nx7q
TeDxk7TF+LY/T6YF0X4tNERZmjc5LR/xnxmvtjWe9KynHpa0iE4X9uiR0CXbMdErzcYaXDzP3u/d
q4ZdsUxqW1PWOh2pI5BtFKgu+Sesqw7O+1BP4A0m1wZiU6DV6BU+PNx1bHx79FSN0E1vXSNyVX5I
dhBX+j8MBgQH+bbtioC9GlVT+AaWl07Ty+Ky5LSrqx57DboUuaOhV46+w6IHrY78pVe5YAZIR15v
+KWeMzJhjyjnUD0tiAugqqK15q6GWUxaDUr5yryCbrfpoongnamNpfNWgG+/6Nipq+iYitH3tNSo
nsWh+ekMENulwSVQjtmWbm2Ziyjuz3gc9wD7CoNzZthnLGE1AhbL0QYRu82/QoVQpfz77OzkTgWD
tfK8aUlrE7HuKxl8o9qktQkHUk0hngikjDB0ymuh2kavLJ3nnpcyipvfxYiOI/3eeXL4TuB/5gLV
bE749EGPx1EcUZkVgarRe/7OwPQuFnWWOZPeGkU/35LOEU1iBQ9EZ6yovTI5QnUKpk8/yD1h2Qx8
TPJiZe0gdMhHOHcNDaPWtiDOckvmVKMMI5hDSUIMkOwNRCCR8G0zsnGkdUJ0lmrfqlQA+6bl9Gfn
pV0bcb4aG3g8WnBo4uQTRUEOgloQhSd5LhuyLtJNOCNypunwtsd4AkSSAiJfs2YIhpl8Kwl0ww94
K2iiNC9/5okZTF3IG6I+ZT9fOpMdKrX4lb7C0lxN8VAkfQLdgUKVPJ1fBVcaawFz8j0I7E1Cn1vn
/O9fOIxBreIRfQtWNgxjV9g7N5HVwpGC2TU25s33RVwdnC9A0f4EJxYrtc2+OGmMLoXrB/0ybmHv
s3IITvDS9JVHD/+H3Aghx1oX0vwu+57DBMWZPlRYbasSMJ5Y+vhGoHtTpqS7mDQRXnmQhuKeP9I6
6Sciwi4saclfBVXTJ9wMpILob8t+TWBbc3U+BXiS7jLiWjnzoOiWCmaEYAwt/TKF9ofgqC2bNWhv
MQcB3vwnxMQ0TTUirFBhfoFlzuJQowzRDIMCFz6mF2UlgTVP5okXFIA/MIfOZw+pnWMUGF2jA3Mz
TtzhiwwMiSJtkGAeeQktK4q7EhUtGfDT8TPPqGYZhfhCt8qeh3V37rqApDHN5s8wlx6aTVnuglVr
ZCjLuJ9+fhWvXA/bniixDPSEW2JHaJPzgwGkxI0lDNDeTlf+XaLo2OSO/bpzxT5ERRIMehNk84ha
1yC6/I+IUp9OQv+gEHN7l6MrDUfk4kHUr7fnVEGqzrjFU+qd3FoNaIatkxx1HlkuWMGOdO/Caji4
VY1WgnTjtEJEYgeHr9I5JPtR505k1pkIp/AWcI5++zVKzlZCgGiBG9JsOp/q+WH3n7qMahxNSyw+
7kbk0traOM7NgGr0aJ2nSiydTXZg+V2wYg9kDYnpxxHHVwZzkCeqdBMCtpAgttIz90Ofo7bq18ir
KJg8OqwJ3K+qP8alKH20WVmzaqULjbfgzfXh0Wuvu3GPA9GNt37UDSAvrYkjxT3mbPBog5HPGK9g
lwa6h6MfPiApfDx/A0DtdAz1c72YsabsXbokfo1lPof+rf+Co6/nqdVdyT1Y8JeTjnOH9qgNZzND
iIGM5Np3QJuECGl01PlNormyBajP/b99eD52duUoTzXI2I2C4im/yfwxduZA/efesoNNYIMqkZIY
FHUIttMrKUWXmPE31Bbm2zyrxBmCPubjjJ2aHf6nvbG5g6sbD9OCIHUUf54D2twCafUMDQvkIpIP
dkcqPrrZrhSVRPL7hRS2NSD3Gc4f4vTyUnc/gEoIwn0C03lVEbdkQOt0cycIsk3SutSw53PX0FqT
g41Lf3jDBOd68AEG2Z6PQhhtBdnFBMsPVn5SEw2TpDZNj07srlQZ0gRLiPqrAkZG/hX2QrTAZYQS
h1paKQkjKQfvZzQG++jvtSorqZxKWCpGm4aI50Y81jJTT7OHqys+3+hihM2HkE8j0pmANJetfOGZ
YK0Mii4sXjuwFe6IEUqkQ6MGX0HgXOiioJAPe5cG/wil91iUECmryD6ur67OolzbOY7IN0laT20n
6ARSE5sxS3gE2+EUQqjcrlnSPxq9FOz0fsaLHpx+J5fpB0gE+AJI33r7XRfXqRvK67cFKjovCIgC
D3kf7S5Xcf4xdQq9NxaTRBSoaHUd2YnlZRVYzMH7zHBK8I/Sq50Nq9bOfvybTdjLa0+s1WE1zC2o
3hvRXjoewnraX5UlQUGeTZNdLizV4VgRKW79DXdL4aVJ978KYJAV4ZjKrYWtAgO1SAzgX3LfEsuq
Ie6Gd3Uz9awnvN3FDAqMY/h1UitYRqEvzEIPjdF3rlfkblTAMDQuc/06Kzz9Nni4xcG41Lff1Ysv
i2vEZM0i8dvZ7tT5UIdSbtKjScEYE9Rzh8TPBGg301ByvBEq+z0tzZQpDgLbBHJtKw9wiRWPcquc
Kxx+PGh/pvnsNTVLuGYC5U1qX2gL3Q5JpmgjwxAzJxNXfSga1CBjjm7xMI18XozcfamrSE3v8so9
DrhSaedp+lbNg8EFU9Hyx1uLyDY+6GZLqyOEn+YxvicxcH8EXq5HKLQRK5pQNgeNnnI81EKbBt5X
ZSlxlFr9IS3ceesYp356O7DOyRrNw/pBkysL1yYRC9l/EAj3ZvH+3Rl9KLkzFkQupX5oD9AWF7/U
J978Cub5a/v6kMviG5vR3BmDWm+GDK1q586CkUIXY/ROheAZLbN8e3/set+SUySCLGFBb8Za2A4F
5Er2gb24szMjnZwPBbCyxzDU+Ry0W3u8y+48EeZU+LcqtSC2HQm/vSL71DVsBYyLh2A5uucISAzv
1fPIwKIEEkmbbRg9hgZS/OYwwMEDWf0bn6VES9FdoXg2WoXwKEX03RW3yUCpP9kkVQADwIHKVtq/
v/vp37UYFMNDPqPKHb4XU0BfS2WY9GQQ0cRvo8FMPQdgcjMxPVC5J593zTS8hsKzZWAphMmzFIt3
fkRTLjXyM7hSgJUUpciGzS5TsJAUqpt+qGv62csFN8+FaGIg1ZcGmNGkrOUFqbaPivpaStXvSv/L
Jrkll/CRkjBUQJNtC/oSMQPhWdwaHcAxGPbxvCtVK3FY+HvrucBreIi62B9INuMrCx/mBAOGXgIn
/Zmczu8dQmw28ikZ58VX8C9i+ambNFaFOq65BGpUPehU3S4oS3Mmo0swW2cSCgPNPopuw8Pn55Uj
XsFcpPzoNM5O7t/AuJWqx3mOUArANvaLkJLSs15pkCc2/qYsMTQj2PhkXy0fm5VzX4+Agl2+zsm9
kXm9XKL+1k6xnTEknEFlBCI10nTm1txG28KvehEcWo7O6tunXagi4CpLy8T1XnHPEJg4Mx8NITwm
DUwbxvksBcpsSj5hLK7rdaqE21yL4y+KIVYsfWhsZMB82hjSlJSjIcMiWHI7RZ9bNGuRDk/78mCW
ah/0BF8J0XFUrMOI7hjahHO2XKW23VoBlvtLKmQJVkltPWdB32jYlzIfvgu/4RvOUTsjOwHtlLDU
tBjZ8DB3NkFNR134P4M88kaYyH41T0U1HoxBXM/6c9hEP65+Hwdlq7+h5yPEoQq8kAFn0t1XsI3a
hHAuHmo87ONb3r/CXmc1brQAJYpQOnsfnYvdGP3kLLnAnEGZuRMQOmsh2AlQJDo455/L4Cf0IG3g
hhq1jWVrJz6ijxE4Xu9Mgct80EGVthLFNa0O0wzUq0TsSGrLcRD3KclvmTgogqh39GqfCs50+LmI
b6O7e0d566K2JtrBooyRWyMJEYqpoM0jVGpvC1/bISp1ACNyt2XqwPTvoQvqjrt+o2EKq5lFn6Vw
f5T2+5wrQcy4Dl+K0lRP7XOqyqDzUkGtL5jhaajT5H1FdCZWRDNPc7iq49bYzJy/SgzVaHZrmiBc
pkJxhIE8eGxeSuVGjD1aE0/+J3grrRq9NgZP25t48PM1Hd+BdMQ2q9ZZDyrLLtL+zXO6kYHH9JAk
ksaYjlAg4VMH5m9SGs0z4/AzG+2EQYhSLF5YBNUv+Bd26QrvVKNoCKCPt+CxT00FAvqa9cEzx+pq
YzVvTFtZAsu7IExI0Y+EtwkQLPoK9G93lnzsCmczNZpz5t/A730FLtw53bIpSYdnu4GFQUp58IXz
xVlZZz56bBdUZ65X3XkNbyUfBAD48adCwKwPeFKAS2PgklYOmzvPYhIBbrPITFWZafli1cyENQ5T
J6KOVyBobU54T3LhvnRiLpz6mVGu5LQreApMB+4HIqicLplUy0CPlMbg/sqzOIljZ+FJVbxNgjdo
vUwkrbxq1e5GxrUaG5GmYckh08+1HtoHACTBDfabXqn5SgP3CMP5U+SUbiwFd3ioKj4mAg3IAqiJ
Yq36e3PX6ypCRfZkeyIC55g979LL/3jK5wn9zl9Hdqd0Tljyxdvc9CdtheeNgGrRjGFQ4l4g4Qy1
qGDK7/ATSc5oMZPsneIJqgkkyPM647FfsUn0mdoP4DmpcAVZcXw/haDvEUYpCI17CeEdkV/8jgnp
TUuTx3crAeyRCQsd7GGvdej6FIzqnqdQV0P8ZV2eXLFmVmtxTl5f4CxCZ55JnyF6EBom2grqFrxt
dOJUo7+77+rURv+UoRKRRn6NKvs9U2neAPVATuqxr7UyTzYmAr1Q2r3Y6XmtFU6nn1Bup+Ron5q8
FfcCaxRRubkxhSjI9VPkUeJVPyH2PVCM+vZZ2WQihMPyTlAqx5BywECqikS3XeEv6QIP9HOKg7LX
ZGzfldV8Kd50uaigOhITagvVJfmxDjoj7MfYS86Ke9q9MQ8VYlcdebflPKD+H82setrdeQjBtIMg
Z8/JckdKUvXD7mA6fkSDvuPq8WiBvOoEpHubrLIG1+4+XW6iw8nrRrbAZjVSCrqSAp0JhLnfI8Mv
AS/pLlM/dneWGRGRxF0+y691amZEW/QcbewLGCDoAP+jDFuMDd0jRTef1RqPo59O9sO/xfr3tcm5
SXIkGM3UL8svbom6TNsKqQ41RM1lLvhvuD98CFrW6xHLE7vYii5I3YFLRwrNi9/90zGNdEiu9ZXt
S/Cm1uII8vUboANCbdX+d2FlqKKTIbVrW6/58ibOLOvg3tEgLpGc7BeV+Z/Pww6D2zOwIUZZd6d2
esU9qbx31YgG06SoI8IFbL7dmfyrxJcQ6uHAZqd2x4qqSt90Ws+u5ONQ6OY5GU0QCwvEeq6gmofB
bSXWo9n+ghqiWbr+9lsxXfVoQJLWBmqhBeIzUXgzE01Y6Jmq4CD6cGkylzmh168UKMNfx/hpCWZu
BUEZdyq0lmMujfJSfQcHSQ5K0GwKxa0JmnkLf2lMO6s0wcLSDA2PNV6UNW47xmLZzmqhWW1WN7TA
i5w14+DlTKOd6BncD9KUavr81Q9FsNHc6ngJZaFIKHrPwh10T/Q6FAvsd3D48DEWUioih8Dmlv9t
ob1sPeyclRgyakCxvshwE73RsyQVuir4fgbIv7yrjhvyD5KPBKyNm0HXv2ZJCOXKqZfxTjNg0pCY
iLKaNA4/nlONgx08+7abbYQ8QVw+rxwFuozDsYrhom5to4A8ecuKDoN31eBFLmHCJlIsSSevqNtW
1OSLJ7na7F7nGlfqN41uw/pQtwMVxxFoTlFOZo+2M4coMG+i838d8GmfZ+MTa6b7r/445fIOG9/I
0TDbtIiOiORChv/dJre4I8S/B5LwCr5mRFjmMKCVTiMOrN6Xfrstr4anaA97xqxi7HCoLdQLSbJW
Ezc+XEf6l1F4ivJqcEGR66KjZfzkSv7VwEoQmv+Mn58bOI19tA+8MmkZNVJPnzARCIWXZQVF4eVw
rEEXAHN+WmEUIFv353hshXCkFq3Tu1HGnGMMIxHUZh2VeDwQINvc+x+PoVFh7oMdEJW+bISsakkF
2jHGb9BdQanbCoq3lTJRWUOu+MTMkga6ZfbScphrwmSWnu2+GlzTh5PwC44yG3YlwpO8YusKvqsZ
PK99NpUafCFk5du9K1LA3erS+MvQ91t2BS3h0L5M5El5u6Hu6RXekjhofvQvO8PTR5xZ5OFzeysh
HCFD2Ux5PrGWyGmEJTFMshTCXQnPY/d83Jndh8HP/jbgNHvOV6V8BLoLstRWoNfIRsVK4ckuuWXm
hPQSnM4h3pDDHu3eImKwhUtCL1J6lyBXmpiGwLqh9GPQ0ta291cJG23ivkkVIoF6vcOwzsS61x0t
UUMagNpMr2rdPyiM5rBCWsqvIIyH6Uwq0e3I+sP1dvWDHKg3d9EqjvSVABSZg0qdgKV0vj8h+1qj
d9wqbgt9RGYBBxvYU+G8tImiDbMIIOrUuK+y6F7baO7KgW3VobfnHDixfbIVgvUmNGTUhJ41IaYE
nmglB4tk2heOd0mpxR8wWBu5RLDh1YC/WMxt6WRHE+zSOW1OgLzDwir0Y8lLWqvQkISyjPHLOuRn
ykNKhwDqbsLicuon9cfT5y004+yrJPKKzuS2LGtF6NlXbrT0qXKTbQaFLcmygpi9ZazvETtcA0Ow
daWde1MAxYt7ovIby0Jv6Trdh0LaMIwY0i7N01FTC6LjzptxpQwHee+RoEsyANOZCuYRcv5YLvzX
9fEPxj+C5PjRjEsn/oxXsTPtS4Y3/+8RL/HbbZ80wGsX2OrVcY7Dc314vaMk74hvDhZLEMrKqx+g
KVFM93oWrHIPyaUCzacuEL7frvP3AabPrGiAYVtnMQYflIQiuC29MJMB2ozwbjPtU2fPbFOOYgJr
QWQmLVpXOmTtFz94Gq1Sw7p8I6c2K32TbRXVuJC90nWXpvY9Li36WspOIMJGXVTMPYt8dN8YKSUO
MPByvWqWhAeSQJpl2MUSRztD1geV2Bwe2g7xvTB4j1a48wkZtUFKclwD3j/oMdXQK7yekYaNQkDi
DJ/9F7RpavKPWgQhwi+/RNjX3OyZFV3mQLYGpTQs66j13VD4IYVPMxbs/28DFtATs3UTm2ZTMzM6
MHExikI+xO3dh2CckFeYII7Img9TMDy1Y+UupmzqkweRV8Bdn1FDa7neUtbnuXj77fajmZWMlp0G
9Oo71xQCexOzETlxoVaQBypeMokk6qCqhR2bSD9eb96PodEA3vA20YG0lcNDCnYaMQooO0pO+xqm
Xqu95E59oFNqe6Pudl3CtKuBrpFzcVE9bNfLNFagreUHN2GyHnjsiVcxyIcmwsiVQ7FjMCvBLauf
X7e8D4ZqhYfAe2/EWEJA1I4UHXC2bCQPHZFi7wXuWNjzV4mK1GH9a4kqEYUHKUh5OLU79AU9x9ZJ
CdrNyj8KkdWSseHjqCzRMsVMZPG08jt8NYCGGVBO6rA20jhnqHa+glMjWA4zUDPqwY8YpyELKogq
ze5rAA/r5jZ6DZy3af9Crmzsx0VCpU0fa7WLjtJeSJRnMEQZoMWsm15Mo4h0JrNXzCiyHcMRMtmq
i2qhBgm1NqfHjszNEfOiyDXtGgIbcBxZ84qvEIYzau5tOhaVTDfjqfMs3zpIH/QS5GC4vKP76oyO
QzG/moqPxMGsLPRxgl+3VIZElyKRObk2agQpNCimP81AdYbw+Y03qsSfFEkXQ8gNpLCWK7eOkLVy
6co3Awk55b+sRc6tA6wb14rZlttksYOHnEpso1q43hTwxnkEmHTnp5gepr4H7cgyg3LTwMt/3Qo9
oAEVPs7JE7o3F9IqEC1dlgZ5bAmkKKy8c3zwVTdhNUWo1tFekRQuAGad/3QQPU3TK2su+a171cPU
2qlRn7Uwz/c5DtSk25e9+7jn+mKC25Z/7FaikCjGNuRAu+epeYqutVmHtiaXwBuYmLJrFoWN0ROZ
7iqwlwx5sb+/zTJy/wogYoWNPqK6efEZe6zpvTBbx+qVy20mhBNMJC6MiVDwJi5lM6VsrIKsM0Ex
4e6ruzWT+FCNLnfnaz3aYI6GsVtc8IkgyNpPhrwSFcKP3mwlyoNQfIOXGpUp/iH9PSptWmHFN4gB
wc6RM4/WeRPZ8Jfk6pFwMA8lYXAIrZO4yoR9OV2g8QgNT2p7lULo/DngnnNTtQLvIey1mmShdEzH
zUoZRLcMLz5WAuaMTFkRLQHO9JqtJ0xRni5k+CPlDMQlduHbQ1yxNp3TW9ob148+1qBvCuCX1wEy
dub2fRRdwwVrRaaAR5bNbmkFNM1Hhz14vL6H7Lx0rCpkDLfGKKtnvfFtIV3gybaOJL7WgyK/u0Hg
YtdkXL90MQozzHAMAvnHqgC/Xjx8ES0xNMLlt90t4xyDCBqMxKke0X/xCpyAK28yaTaYngfaIVuh
5Wh+7vXzCfcbWDpS+pAtPe3n20BnnMDKwuU/I3YOjConKkmDIKgYwBULnW6dGhO+e49JH4rYvAsQ
IqcJglDNU4gUvb8oERS1l5IllDSfGjSJW3vwjYIQr6gWXV+lSxmuTFrmBYC+XNjQvqN3PfReQifh
TzVkYs75S7rB+SsPbOpnavBfItovZxstEKYEEiB2HKdK4OiXBWTv0nBuZqKjGhA5iAuq0jt27A9D
vo8IIUMAOTwckV02MKmC+NFGAcKdfFw04r/3J7B3+CSyv5m/Vf+bqUooBu8QOzHWV2KcP9PxKNpX
2t3WxBMPXO0I9eV5ncHTY1U5e2lwnkcUa3j/KahUX3LrVElkybdY++IqYDRo01FRCThdOqQ4TgLq
f62Vg9Et2sDyk7K22rcBG88Yit/XRETyMlhONqvYgKUehtkjaHrAJWLRNdFsOxfGTWnu2oyIwcgO
x7F9ZliboObqtwaODV0Zk6yA3ZRcODxsuHzh81It3m0Jnt7Das4LBOZyyNI9gH2qSJ2bQeiCWu5V
sOaEWhINaphk5HtFXt5T4kbQ+UmIq4vIqpcJl2r0Mv2BpK7O0D82eg0qNjP0+Q0zA6/8HKEyWCQd
v3EXOic5EjgGlgI7icv8tnjSBJpkmqUTAH06rLALEtpwt/saH8iPs71vubZ22rRDbVC2rSjxKTlO
W5cOJakZ2FPt1o0g3K39rx7B24rqPFeU+36qsT49/h1+CH8+s4MBbMAHbEoPK46zCkuuoyUCIUQB
LoLq7ZqPcyharPhN4xYWQYWTLJ/Xli+QHlpIN9H4uRiyZaOQwNG0BvlcvwuV715ncbQ7+L6L+gJn
sDBv33UtPTOz4ukDr4792tXvPbvuJJCiPXSdsS5CWwnQSq4IvsY64iWfxrpp3+Mt3vlfFEoUzhu/
qFLB3OSZ8K3/GZxNHt/ytlIjd84RIATdT54LrBi9twCMY7PzaBYQmbLlaZPy9ZKBGoW9hB5Ouf4S
fr9674JbJHBnQTAT2uYiZq881LcXdJ9V2kFrHtVA8NQAiKyj+aTte+W6u8iNsxkf7dCkIm0+sv9k
0w5PoMtbr+me46fO4zW3tPOZdWY1lnaPKbeT/6/ZDWQCOwoH2OqwPVQdMD9I06xKPrvvjlHxmTWR
yI5Jr1p1DRe7irvKZvX7nHDg5VN6X9EUMIzco33rX0Bvk+zglDyDqHv4u+JSD7ihjbShek3wJoF+
zmvqfMR/e/8noAyho0weiroRXMHD7Io7jcNfqstedV+lM745gl51uUbrOI26UnpSQpkaZKtScAmB
LHTnOfSr9l76qrYLyDkmMYjnzlJ6PhVy6r6kXi4UvBzL2468yAastm4LeUoXpvENrbZOGCJIvUIT
oKzWyYYKs1DC0I54Ov+SbmCPMafAOZuiO65ldgMghWj0oz2PdifgFOKuCq3SkwOg90/yiG1FziLs
v9MGrUQ1Vi1vl87iqkqA/qIgu+5iaUft9bjXk+xf6nVh+7WqX76+sR5s+oqD3uPULlWZwEYMpCjf
PWBCvyytLLrig5fb7pJVX+/p18xbMctmnZjfrNZr0OOPaoVIjyeCNzCqHYMhInBN/01+OQasf0RP
f9yh/3kPNY4Wa2SspDI/gjzSGV9C1IpkRS/NZh1yZ+ScZYfPEoBkdqgUi91bBU3898RVJ9bla8DQ
QJYVshCDHbjXICktrB/s/PPIziR+JvlP12pEQRgyVS1KHn/zhlw55Ht2t9nsOLASnNzM8wioCD2v
Aixh9VOieuKXmsUqd/aAwPg+QMNHsyTHhrXj7c8rqkQqYhZpVg3RBGU6kTNXhlISvZgMmPnnBGtf
guFUzknlHkg6Jtqr+DGx8eHgUDiL/nQybVoKrazgEYgg1GtXvptkvUhP317tWCXPY3ZE9IGSVxni
mE1PjI5KQirOs99SPpW/pcLyXNl9mNh+jntTmFtyrOy4ks1MGtDtwUk8e567q70rppp4FynTyqLy
q7501q/VQgfWrrBD1US+5WMSmzuzzxv2wqtZ95gpup4NorvJobdli51/Se69xfJgc13r7c8Ps38f
+/1RF6Bp4GAwQh2ojYoNo/xTQzjnKz5/ApcaiT9/tCNOPPpXeuzw9r2sMaceYz2hlTQmft/atDVk
6eGlMZhCXzWFRLaZxERC1K3CCqnelH2wQ1Z2tD0V7D9GhuFlX9FMmb8Ht/eULBM6CKrGTWrqSJ4C
Vu8gyPYyT7q23v2JgVhpNoFuGjjkfrc8635J93Spt1vE9da6RUnwcPYvc4y6h7ExSg37+xrhBDF1
79yCSow8aRN1zQqBMq4fVY0pJI0pz4q/OGp0yHtEQQxdFiMM8Ho8EwPI9ra6IM1Kt1pIzbjanyf8
xeccdNtRK2XPviHCLwF6Nhz/hgdSQYOJQ/ggKQLXKrF25wyMXnVDqIQdPqQeOu6X1pGPyVnR5wz8
Ij0Hf/qZmWan/drK/2s43boAG9QECxzl93RZdKLqQ7fvxQZsf4mp/HprG+PVS/eAZ5XxwCO2sfpj
2jBsfF/5yWsosVqOFNcFFP68i4/EOT6LbzRBuypB3hg7I4j1+b0o7kTBLEoE+BSeY+txZMI6KT1F
NVLMrmT1NffwB4nUM98peainYLYzwG1vUX14T8wEnVVNXMZBklkwZ8US3wjHHVgYCYco21acqzBr
7GhltQm6Bc4VpWfLfwGyWG9iNrUQaRHkoUPoe/JQn6OBfpnin5n4POgLKMPifyvKD/mtW4Lj+/cw
6NsJgb3ov2YyKym4N7aPFg3p4L1gwGrl+a3gzR3NA9geLuomeUP2einjD2n9L5bZipAkoFOUO92J
fvkm2bDUbXd0HqZJIYHtxHv4mSOTNtkzURNVwuHVzUySKc1sVo6nhsA3c1oDJOJ9mzECpYhSCn8q
ww2wJ3J+u8RcoJMWXQCGgSokOiNlyhZyDnkPqndHQqJmA/QMEVbhfp5tUMUd99BGWxmtQknxUH2T
BbZcLYHju9w42obUkvKS+ytC4sXZyCMWAO176wWIgFECCjWT3c4o9BY3E9FEGGRPuhtlPTsqmypN
LCsD8wPkz/TlFPx2zVTrRLbQfF900QOe3VHo50+kRTTyNILhlaJvoOZWp47YwLDmZykyJ8CmNcMM
qzniTa0lISHCj5Rt/8S/6Retz6HN49vEpInKybb8h43qfZfXJ2toRUD+TdEyxaXol85eW93U1Kwj
0G4aOt3YC3VtyM3/99cr9iNjEVeOLh1Ex+ZAnXzyuEY0ALv1UM3SSEfWrh9W96BLk14hO2nQQTsS
6osZYInhEb6+qXIaYEHwG0vuubDOga/y4sSVGD1Y9sfWqhkPqDpWa+O26wng8Iq/cvBas33Kfy3x
I4apabJAt+d57emxVDSJknGJUWFSsK4lDKFU54664MZpL9lRwT4e92Wo04maYPk+Lxv6ieSiMKuY
E2KofcyViaCGzfq1h5QMgtXRfi0fhuEE0XCl70UYFmTjDI0J8bVE0DfgSU2u+xh8uR8CLaYFPs7e
nLRS8x3aui1Oqc3/n0+LnvBqvVm/j6qySsrZW2gm6oU19k0hPx2zDZ1FMzyLnRunx2ihKDmykT2P
bZpMZDFlnwSHtrit1/6cojoOOCReAUIbLZDb0ekfxwBPmQUn1gIrWs/t7AiQ9QDVRT4sMLKhddAI
dWVbnpL3r74uHIxyb52RNicwchDhesamkeoUu4ApgFujAUanV79ikHURAkPWznnoOZdTeZZtRIiQ
z1ouCHOVv6GbCzpRy1VOYsC82eagoOiHhDjipaj/a7xrY0q+29VCplR1SDDv5pvbhCPr7a7Yb7Sc
xt2t4SRE0Dr19mttYOuW6dX1APK8uZogA2VEApYPDXnoqwhzAOzMBl+25u9gW8GiNQCnEA+cccmr
T7WTwyxTQZ/2hBf/2Ffha/ptgxaxQoB7PoflSzfz8SNge/p1DORsSjWVj4NZtpOwfCoUY401JFwl
KmoZvKLLjHXWvM5zrlocap4PM8xKWTRI3obOncXQJOn6sp+fIEG6leCpuhv+1ndP87Ywhfn718yo
IxD8YCqq3PJHwnglisn1XuAFWn3b4I3n6qJ10UcsqO/LDxtcGwiCeBwpxG2JOpS3XxkbjwU4fqjg
FcvA/Ylnr6SnjLv+lN/Rs8ZoxpoFhI8v+A5jXOfL+UTPtqCnybjPUmdy2k9RTUH1zs2i3B/R4AAD
8BjRcwU0SppS9tYZXw1XJnCErEmQy+7ghZSStuhdL6pD8lqVjqWOjal/W7UKqHloFWVZJ1NtWEWf
Y3+XwcUNBgq6ZgdeSiutcqz5K5lZf0UCsbdUTdNfdGoEQoW9QruKCWr6Cxv25FtT8k2Rdvb6AbKz
hWEQcNizBiTQrnRsJGqEo6F2H3jBStxEsMunjM317fkupusuDIkl2wawhy5Bn8Y1sseX8pcZIZH3
Ltx6yF0MZpzYGnp83InDHKJJfKEqyEE3TrUwYyJb0626ypVpWDbaeHaTQYGcXBrxztdkdL17lrFp
bLSRJ86dTnQyyvuFxTAcBybK0PigONbpPk/SowCCH2Jwg65n7dIT2CSDMbSopHxEa0P69mxLn/yr
NhiqYZAnqy0QaBMg7rxVOmmYRrSoxD+PAteTq7YggFiV4MSzTUlWAKua8zCjZSgqZBjox/9j23s1
TkhAGx3z4bvUgTVM6HLaB8WU260iFJrjMKuNC4IjpEHYYOKVYHMjOV+xaM4xZAFEdI2lcOemXeXU
x158bTA86+GP8XKvfpSUpmvNHcFjvdzu6XCJos+W3+r9W00cZvroS0NNURDCfVtWWYBVsJvmgiyh
Ar5um79y1zje/mwvA5BPtRVlJgiBG+pB6jD6KCcEiZQYbOMpSHBtfhSFpZPefH6TyRPucrWi2GFI
IevQuOPZjO6tHqTRFdoGE/uZruLGo8neSmVmxco1k1raP755vSEu/7EUstwWBQloVeASelKQSw4Q
v3wdlxebhpBZTx1AlqwgKZbZwn666YxJDiWhR3OTYS+gTZA0mbPlliywWqaxLPVxgAOCJp288/j7
0nXlMCzZQtkERZoE370Td8amJ4cR7K/2XtTxWrEWQB8JtZ9dcf0cFvH1beJ/3djYsVwbauPRvHaK
FfSg5l6met4whF4MRL6uf/X3bpVIXOMKjstYcmf+Rp4kW8Vz4fX9WAn9kI3FUu1NioQzXER2lcAe
+RhZYZXjwob33xOcgXp63IlFzVx6wjqgsrXIxXZUFBNloECFsNzz6d0qzkydCfsAAcHXpWtWrg+M
2hIHZEto5a7NgnkYZGP5QUJh7SL3WTHUkGpEwBhSJs3VI4ooH8Z+6QYgev7BNJhSODYLYpCwfoo0
MrFZWImweCbcErZbH2n7fRQ/35ORGE0zPraKo8uiTzpdKwcB8jROEjHZMVlekVA/vBeKLRs4pjar
1NxGFmtiznBIqglYrBv39n24bH09RDgBZIZD3iS3yaML4nR/fdoFOqQWH51dcLtEA1YEOgRg8qDC
PW1lW4P7hj+KjRf+3lBMaa7QBhrkxaLgBZhZ4WyAfcmvgKBC5oVoOU7wWIt/mWshm6YPJsbLXrUC
B0M/vcTV5AAMjvIZPFbgzOG4+Bhs4mS50yTwcK6c8rRyw1Tuo2IhdHohcJX9cSLLKmWP4CPk5j7s
4N9MdTr9dKjXUKjzy3KSi0uB9E+0HvveVJgXpRwa9MjYNSipIZgQMO9OMhvQZ9LUHemmveWDFrW2
VAAgYjIT8XkQLsyKcWedmTV/30TFduTcpYGnl1q7qlIvvjzSEkoey97B8MKWyjN5UmHtrWAZZ4kb
/ZRX0KJXRa8PiaCLCVEz0fDmda+5LdIxrPaDDL/GvVAdyygHPD1MozWRTp5I758RNg2YKz1mCmUv
Jh5OI/xe4Rg5x0ZusOdrzCobNLm8w3PTtid2C3wrTlDuSv93PsHBkJgYiJKDSJuB03GjFn26dgDI
clKSpFMrTw0T6iMxexEulOrj3r6uB5pmYRgEX7knlULOtvx09dQsYAv5Q6gMA7uCibWZo26liLuz
DQNB+oOPmjCcjoyv0LOVgqA7zppqDUuoJoJt7212FvUguWvz1rcJ5RoAxgXHJ6YNWQPogyNKgIs8
HWu/jDNRokVdZEHPEEnaJjAOOuYVPLzFf2IY4UzumzLshSzYVspGHOVlT3qDZQ30lm8HsI5ul+pS
861hlQezG8ENYFluWFf5/FD3Nx0CyXQxNt3RDXWSjP2OiJy4J//LKI6eoAI9P9JFvbMfjMpXaYea
wo6mmPBNcoChM/GxD4Cn7NdGf5NVdWbkAIlcn8lI5iQReAZhLAzZEI0O9UastkW5D4b5n8VmsPkw
j4L93VWaQk9bf8XC/1JNVZDVUva7Oe8MbiTDEOH/8mIHD/BMdFWEAv7U4ATyc4IXqRgrMbZgbS5G
QS7NEO0c/Egcc9d/OKaE8k20BIgWp8NGMx75ZdcItEWjXV44fOYLj730jXH29Nkb4AvgnsqjqLKg
x5qzz4WZkg0iAvX1hj5Y7ApI9KeEMb5YAszjM6wm7rzcf2DYptfA83q+c6nRouIJefJalDhbOdoX
wYZt6IqF8C4kskJVHiEhtjVb1BS5mI9viJ1OeA6gzgwCD2P2MTuKKG0HAdXiGe8r/iJMDyeqrnE/
fbme0zm+A4gPBavpvpx9RnAl559NRnPdWIyTgt6u6EnAgEwRuxXYLmuZrcA/WYLjegFOFkny+CnL
kUpKPHvo6b4ZZNKVzOUctMUiHH2pixxrWXM1MKfZwYHaD8H//n8c2NYMD9GQHrS9p7gEwpwRM1ZO
Oec71ond1CepVlgEdl1Qluxiu2tyTKQ3TauoRx+gKjvmthpK7hPhz/mYsWJuXKvKp6DxM0Jy47nu
+mCbh7x0rtQ6Z3xBNOOSlNB/bV+cwq3b/+G9PrkaXsp6/rcN4DX45T+U7eVhlNEjtRK6Yh8CfxhX
Zsoxw84T+KHaOoxFlCTLIh6DF6JVENJnWyQrUO+sm7F58FjwS+XiJFQNmtCKylGqi7lZTwTDGJXv
urmAfNUylGes5i2pSTBXQhwfQhVoV0gpvCSnI3MTPmmlCpJ1AAmZg+txvzGya8HpBslFzdUQDnda
prgj+n/bn/07jMGudXGnDlejM9ssG1UXNgmhNoTTrBF730715OzlXwZMMQKW73i53+Uh0fE19PmR
eMITCJgRb5DuVaAzoUZZroLUd8t1DZRn6SzmshxN5gQLhNnDdp4XOSrVrtLk4XHkUvuLGGbd4DZ0
TQ271J1ToqkCHPaA7RUZjNVvcx8iB/Uh9bCA2wD3bRsf/4uW3sh2/R7z2/UoZcJB1bZRvEvh5WMf
h/1QPdhzxWU/0MDZ1NuNmXawZ69v4BHPKur0MxdoODDlUo+CCNMUEATcwZQrIoUDfQ2f2qfypkgw
cXvzjxfPCnne1NTpkzG3i0fKHwFto3i+dsgqAd+Q6HVIOTSERp92m2FpFfo59cm0ohu9xvwezYFL
vG9jmfx5+z8bB352++xU4aKoM4jPd6lRBwBd+VWWmhCRGOGL99eI7gpSvxgaXL5YE1i0M/8NWl9u
GYbDd8TpwDUbPuiSEAeznnVNmU6t/HZ1ZO3qDwJY51FTtMjCn81sTtafdyHC3Zvm62GHstCGjS60
gibfkeJcWvnFcCRXmYA170x5M4v2z0oYacep6sRgFU+nWYUFoUJSKS0p88a8NrbcLhqOYk4I0HRa
wBdAAKRmNRlo1rRHGFczSYiLM5LHa/fc8T0r+xVv7b9j6/LezmJ1N6kHJ3szs8g7rPvtZpD4v8+F
43mZQof3EfO9u9Ka5+gfR0C5C778LBJ2SF5MQbb8pYH2Bs07vn6TbJvAITeuIkJ7ndePFdRYU9Bn
iPJHG7qJclUGQLCHW/eJWw9L8dDIzA/gHqLduxuzVBfdAPiS91MvkKcvcHcgRP0ZvXMZoWy/8hq1
Gf0mbvI8adZ8NGWwrQfp12BzUCXMq9X1gSb4cd6T8wv6ihvLhXeZa/+Qm2zOMoVKCnO2wqH76C/G
GX5Y2j/YGiY098DobKG07U0k+pHsbGafRnQnEgya3vRK1R7wSVJXs6GzeS+96aOk4t+KndPy9iib
eITpWDUUiIEYHNSOSzyDwY8ohS3DWoxbKEJYkbeKI8WAsaHKeBJvuUrIK8uVBB3GPjdI4SAPNhIp
4c0eHe9MMkPqblyUD63CDPceazdvJKPoFlZaxQXOleyg/a0WfXL2eofcJgnC8gaAnSzvnTKH63K8
UfE3msYI1hMQA9z/x+HaZ7AAW76hFHiK28iDiQu4iQTrwniW42e0KuQXlPtHu/92aTAEy4T8Z0+V
zmXVwhkyLqB92Z7BNYZS3ItUoAI7uXF2o3lotjVYyQaHxuAqdisF2JkaPpXddEhcbacKGjqv/P6s
LjiSa37NKt62311B2p8C1tScnvKdT060TyIIRMDcXzUQ7jy99L0lNhExJ2F3FzXNtwJL5dsPyqwd
KHwp80zdDwhpSMxCgt9pVo212nul+dLZEflZndiXulloV7KgNqRfCyAOjpB/dk2YTn2ddSm3P3WT
RZoENA121ssLUaz82romGFQhB4bJxj3K6hxEnKr4ueqkcjqo9zHUpuxhHf44t0JwSSgn6wrAaHou
J37RY7aI1VHdLkfdKqTqObTCY3XlZkPndnhb0xfhYKWqgG3UusJzdC0wavkOssbA/EacZtGxlxOT
l1vAXBD7b6p5QefCWzUxrCGddmJSDzDr1vluMyVTjNI2c7F53cPeCgQSgHpZHDr1bOVCxfxuBYON
7GisXfcaDGRakGAM9ejBZy14C8NcfWzEIdEuEcVn8rskhCfUJ6/jivjKNNmwV5qk1k++s4MqKJnQ
BLBVPm4vfX8OQ854nX1QRfHCLdg2lssEG+yY6g8zeAKx16sCe0j8W+uEXUXrrLY8CJ0mbUQ4i+4L
4jZSBg/zYjqL2j60hd6JgRk65+f1hsrggfWcO+UdjskdG5c5Efs/9qrpSIsOral4fP0dlERD91gx
PTNdHtmqN9iPUg++W+HMI5ZqQ+Fa3JLO1VR6UEXMptovbDxPGq65dQ/2pBIOoTQfWMpC7QJayeoM
8YotCO97c9Ti7GhDvi5IS7KKUP30DKWpLhd/kvhVQ66v3UVcPnVpxhbF89xec+OmIo+4nbOM8S/6
pMiPqkBM2NWnI0x5Hkihm/taxkKaAcZx0k+Aut06+oxesfixO6s3JdwK3MfAgo4wqY4I+Htjou+j
oCjCGwuSF3p3wx39fT9cZ6zJjbijw23nWVqR/nRk8W6kT70hUFJWw7e4/VAtRcNV0IjX9XrlPRMM
IPYlYLphIJQngga583mn7564y1yoeNWNnBRvZflc+kzyiaIMNQMjxRs8dPcxm47pO7AvdriJnw5Q
3+DTefOp6lxsa9SE7boYxKJ+xx9cMLL0vP4BCvqQypa6K4MRY5qfzLjPWc+MjxekLzcJwisveJqr
MilBg9qHudYTOdUx9UIACf+bm7bzikcojB7rF7Q9a9kEawW4ADbE5J43/i/wJFx0KwSHrmmUWaUO
IC8TL/uERMeVbKZJfSQUoplLkAR8hOxOBxSMPqi7gsO4FDWRlxHFKSb2xfX/kAVT1PO0fJU1llnK
twrpTeodpXpDzo635VCRfY2V9zfibdy7+8kOiePLNbzWPdO/uZ7gICtOPGoR+a5HQ+xhf0xHRpCY
6oyk2OJeXVUcTJaTEDl9aNWYiC36NiZZ7BOfEtyDwsECdMIvKvcb0uK9X8SHp9YQHXBbjr/RgntB
zggaSN05jW8bfe/aF/idOiv2RpK+nk7zXBI6IJaCimLzQmb0cRzl89asKV0P+ezrkUk4ZuCFqHvm
fs7pEJ7RjC7RUzm6JCyeh4rrmKbN6S2nm1nCS/uwue9uGo7zDAiC9YILUPlwmk8Uidk9+gOkAvSb
KEZ+Nn+bm2VeNLR1l51eK9PGCbT52Lagq170zY+L0iiEFXwboSgOxJQ8jndWrg/wLV2IjwSIoTV/
6Kz0sh4Vwtt31jHBpsv9VRNmGYxXKf1O/i30WzvPIlWJhMgxBHNq+n3iP3heqM2jqWsu+mKVhsjd
uduEi9asLffiT46Oa8DwRoazvVGX0JXpM6HewR7WgzVRajHZFIcac9jwgjPFMu9JyIYVeYeM3klQ
ZhFEdcYUv5LQqylG6yde7mijcrfVGIS+Ur/2ijOFzhOyKadrA+xevbKzwRRpA+pmexBnVVmY0cIc
KWGz8U6E4dDo++9uNzmeVWKVg9FCCNtzVoQM4CUnNwa8rdET+G6jl8heXrDwrJOyhQ1/tVoSu8ep
8la4UjYBk0RuZ8C1d11xrLYWhurG5dIkabgICIV6y8XRh0XnNCRN1piWoTWNl9CMbg3goQIi4RSM
QmAIzwkatRmFHIoz3GTNwATfdOWK7FIjXc4ZBX9SkKSyB0+wmSspScZ14/d525S0hp41JvfpmM5a
ln98emU+Y7moV4tBSOLuc392s2g/UxUKBFlwP9mvYEIuboNJez3UkgUZz7XnACXOLFFWAxDKX7G0
UM1pBP8Uqg8upJqySHLKMnvMDn/PZY6uqbTyeKnSyeMRZXSwVmuS/5Nl4ZTQjNQ2by2B/mnQ6+Ek
Hu9fUIHs2ySD/n87VUWNsz01byIXEwlk0mxBTc4QVwMPOkeVQcC9E0Tm7cJeoWVdTfMAj+qoLZIr
nxHqJWelwdG5CMidzNgGz9Gr4OLbGht6AObdTTatuo5P/IruFkQp+jYvWJAurqcUp0Zka/sr38d7
2Yx7CeTb4naUun9hbAQxGbz5QwrU3aS0xydPheTtQvVCDtwIjhTbzRdaJ3krt6F+q89t73UegArE
UMK9YThhKD1sHkKLbupdf+lKccWzpq956N0IMqN1Sjlk8CMbuKNWcfmTnmJicHGRCu4n7ZqSAk8h
gtuZoelJQfFNZP5IkvRsS6eVXsn6g8QpU2rmOwAgZQKj+HFW9WTSDhjp12dAJPbhNNKs1GXadzm/
GLZ4YGauQwfvrwRcIggHfEHiFzdkLTK9SLV9nUTLcLifYwClaYq66GVlFOGKD3nLvjyTRAnYn7G3
lUkFi46eM8b+oVyLduuNjWyte3/1VOQ3uJVyag/rn3YY2t37oM7EPha6Hfvx4PKAPIY6gDBwfJlY
vv3/0vcSBDJzu217qOIM3vVZszgyud8rcfgDUbzUoRVlgXcq8aJ87BvaJv9DDcGVp0ca40/UYG3h
M6zkVLutztglSaMa+AENNtndh9JlFuYHGHh8aGu6cTKplEJgzpRiT72ha6kYs9ZEecpzkbkVjeWl
W5NCDby8wBQsHvGlSAdCUR6dJD+GmsjaOcY0MqGO3wVY69qqnHYV4zh6gkAzZ4aOJzvIKYu3UaPM
ZrLJUwPs70hOseXmiCtQ8ouYCExAxHo60NlCoefmV7sMWt1WBeV/EdlXqNnY/yvKFXX5gSmmK6sY
XEPEPVjZOiU+dPzmVGV6BZ02NTSUWCvu9YOwLkPfH89actoPq298JqRRLkGk/r9gOo7PF8frZ1k0
thYZHLUs8PDZal3SY3UJYhZ2vMeZdR8gx4Y3NTUQ9aVYGs1AFzmTmcYJ+pnw+Ss4i9SIfDFaX+U+
kmmgMe49swLOuB7jMn6dnTTsuwhGRY/urPHYSg7/9IW5BJcaWSrRtVaPS2mRGynhfJen58ug+TjW
DypJ+UYzvgJKRhS4rA4eo3AK2tNzbg+B+6pSPzGtoKvtzQP6DuHbtB9OO81pMNoKSLCuOCalczYE
cowCnpT7gTypzSxbBKkbl3eJZgOuB6r+pNCANW6k2Hkk3+2GHQr/nzv1adeWgI5pKG+0sNJsPmFv
vMd4EbRFTMKXCRV+iLa/J0SN6CRoSJ4YqHAzFnyr7f6slQEcOI7tHDdjME/cSt/Y7yaj+HxFEc2X
Lwt+yEK4zPBWOoIQe3TMsgy3QqQ8fbpXzd2eQJ58Nrkihp++h3YdGon8ptmTdu2zq4YaVypmmzS8
pyAaT2xdnqqi0NPPHI9A6gfWd+gkNmj5drod/1IkUUH89zKp/zKngN0I3D02efwrgAk6qzZUoRwq
AOxx/LNjr8JUE8/lB44DmWEERP9tkDVjPqA+N6Y4QRK9WNVHxIitdv5ExDfh5gt7GndNhSyUX9Nx
yx0VwSq0ozCYJU31UL9HLKqw+mgIqhwW9xgDqHCOHn2Os6AHqLQTshqx+mgQEQSbQARh0k58bAgR
pFYKaLo6rdFd6EYTXhDMuXl7dqpsXjenFjf2JVBR74PfS2ske4YFAJ3KYNzF5m8xUTxOq7Fqpmqm
r17h2e1UlytkHerVA2qSsiJXByob69WOi3arh6LnRqKwRtMlcsmSKS6QvWN812s9SLzs+uZTEK04
rd/upaQYfNfi2ubcIjEn4Slb2vqKRTIfnWnlzgdoeu3f+QVoehoRqkP/WOCYmvvkn2gqI1yWjv48
PPEWT0FQyA5hw818Rc7OrA/C1XFyS3Nss4ggJfnqpmDuGQP591gawx7h+w7N0MTUPKaOUbbhxznJ
zci/AjS/lwvheNDS+y5b4D2SqDNAVMkbSRD41YeIBSTrs5FH1t6BLH4sYCWuecY1t1CXTmrTf+BY
nz7exL0lVcIXE1VCvjtBXymLhnoTgPNui1oQ5WYbvulcwq//FxkJr4PwQPU/JdsTWEFdF2W3ZWXP
EgG3qFCJsLOedrAvP77x7CxORs4zFmiA+oS8iF8pjYNSfDw31TDp3uHaHImjaqd5r9EHe9waLSaS
/TAjWVjrPd+yTEhrg4PMvN+MHOcxXKl3lkS5BATG4RVJXNU6zrsmhpnD/Brx/nqB6t4HiCMocrAl
DLZF8Pusj07ThqvqxjqJxzJbi3orVXzuH7wqfn5OcBMgiCFBOuV8/yWX3Cd9RJTbAoFqxVGo2LVW
Ul5N9okuUW7rbQwDWPju8Ucsrbu7fYW2O9ahRG7bGijowJd2HYs5ZABoPVyCGFLmcEdXGGEgcHcJ
M8NAVZ7khAWTU5TPB7S1VhSPPh76Opu4FUaYfcjY+5be8CgDIz7tz9FSFqhGMY4rUHihVKvpZ0tU
MmsU/rGjK9j8/oeY2qezcexY7TSbHhonsadXnKka9DATqLB3klyYi+AAxYoNK4p4+m5UUQAH1l+V
B0McjRN8UrJp7GCdN8cEIQyiDreTrlLQHO0ryJsJCzKKpuX94s+nvIa7UtiDJN1D0ftV1VW9eWjV
d/6VY7arIiidZKGMHHVx9+i+60vSBh78CijhKcRKfW5SnhrJcFtajOYI/7l3hAtdYJRqX9XBMXzU
kPYf5//HJY9iFXZ10fptKHBhZR93pYU6kppBhYboG5st9A4o05aDbkEegWTb8LvQvj+gI7mQ9dst
NVVJQisQp3sBIGcQ8EXknq+2ecjUMKDyP9TJAWrJK7K0q/vbDb0Ujk5xK9MTV8JZB1XAx6Dr9M8r
mRfBYwPi8tefwDlXtpJF2PL3C6YJEdEsYBHr0RqzyhnAdo4N7A8/gPNT3iBxZB4hba60Ns+2eqUE
4E+DuCYjnFVr1pIEqewk5TIVMDHC3DJvDo/xPn7D3dVeu9KRbtRqOlD72GH/0i4ce9Erd6CiAqU9
m1eIoeYxIoJ8hNqUze0ye4PZS1ZiCwTaP0lZfBn7+3YBYJtHj++evIk9jQnKRM1pzASv7CxBWGZ+
J5aP+xwolU0/x5ipZxvJEdFiTmmTHTgbXU8rdLqS9BvGesYrs6pV67i12VVwH2cZvYcPbu5oo1nn
5KInW03d879YeFFXFJtgyBhoJDAatHyY5ol57AujDyONI8EZB2d4Q31qAzpi3M4k09SaYzL3e2Sr
YUW6sLPlMgLgWEcv+BaE4CyBQxB4AL7QR77ouN+F7UoY5/MBiwdAoxWJYLshqQ7DR/jmPPbMSXIz
k8Q2nr8W7JVyxq4ymjw0HTStohHxLPs23e/C2Dc9iAWsR0K9DOj92VgZACvAu+RCCHCCQnkGUmXf
QjEfkobDWf+V+S34d/42WWJc3wfJw3Q6taPKTkRip5e97+A022TRUWk7Pn1D/8DCqEVAH3FJUbHK
VXbn+1At0Tok9mDUrOe8kPeuT/HFOo4z/I03vLKhpstXJRnzqz2gf2qxTm4rH2GiPqZqvVvBKOLP
CkLYa9SRbt+sInhBj7KYaztuO21kgqzrSieG0zeNltNNR2nzxeyPfxITVTwJw35SPdTdDdKQUM1z
6W0wSUsUZL4b2exQmd0W5gsRpWZ01fuItlGvr6qve0IyTuPENuNNqLTjdgSXitKCkO+5LvGHItcO
o1R8kC2uJ8E6SIVMJj9rbG06q9Glk0acn47KuN+C9Is223IRcsnmR9ZEZAmx7rD/XdFW/huwldti
S7FjZS2XHZuoltw6nuTrd/V5sK8/qDyu4nOF6mxwhfaXIGYpKh9sJXXd+EVxPhSXRr2e2ZESsR4Y
2qhzrcSp2mVwj0dkPbbhoN/WwAAsVfcjfCl2Msyc6RTSBserX0SWuBUFdhBcX8CwxUyiInuEbdSL
eXlpKDV0hAkFupgqMPOtydj2opol1Ie+B1pEcqEHEQIUfnBmfJvDPp5/G1EMas6vSf2h1vJr+pOx
FMjOtZGY9dtIt0LbozCq2/1GyZA/jfyrn5GLYeBtwdhC5itBq9wOsOj0nS2IpA12/n2nK6ChraqC
IJTNvHJzlqXfsK5qwHiW8YmtTI3zhdlevzQ5aThOxBvQJa4qlKoKr8xCjudIEimV1MAyos1gOH0l
CAqpIeK5fIpwJBdJgZQPK7wAG1i5wqbVJ7/XukGEH3+3y+s1o+c3HTvKqdsUD4yULCAxmAZMimUo
vmObBbsOQLMvjTcy3wCI/bI5g2UTEtEFu/vd30I2p1poxYFMX+Q12d79K6NKUBm0Yj0kRsQrAPfF
TgwlJzAWvnkOAMNZgOl2Y80kmlcxDzt3K5AdDrT6RMM5h/t4E0h+4Z5WKUKot+PrV3jbb82X/a/d
yi484xhOwAnYfGBcGaJdH77qnejRqeAKxt6NBruRN/yv+lBF2+Vr/e+AMuYHEZRlR+5sWiL5k02W
O4CQN+IjxVV5FNj+jFbTL//0iN3DJCbTO7GVUqu/lLLn1bpPjACp83BX2xNRKK63/xYPryyuLOKI
KAB6td7n7wvdMHBNJqwSPxvcn7XqF9ZmKaINT4KgXiZUM9SnGmIHgkYDmniXLDZeIJx/VwkC79BM
JGSKfI7oq/J7yscwLtt6MXYXI6e/rLucaGxXV7kI6VfRuQiO5q6qGy5EXPgrgSNzjNms5MiVn5nI
WVZ4f5fsQuYhh9jhcqdLW3PONUmZoDGbB1JcyTPCFoBVvofQIDMD6rm/S4N+EHl6pHggRxLensz/
kQDx8aNMkoLDutfCF2j5jPknIw2lcwQVXavABp+F/46AZ+4BqRJg0g1z64LGhf6mOj/mN4IuIN1w
elSG8SIEiCtFTE4TkFzbaXoeeXPcpyfGBRtyqVgw6GQ9jz9hyoHAoznsk+FZcciB1rQ2kCNzz25/
5T0YYZh7O4n4w1HdQeLoE65V4tquwtD6urem+Wxt2NBjO0UT8r+CNyno5DKPbhiJMjnmCOUxqlFM
20douAhwFu52hMdNef51uRuzctPY87lnF+rteB65YkkuSWv+iRSjoE3bEFVnFw93ROO9QDFyc35N
IfGTadfDPkyqawQOVfyYL5XuHifdKLTmxONllyHIb47fiKc3F7+DG8eTNQpsCzdtJLrqHbvX0ALS
no/kvXvA2cbuToUnEbX0ZSqbAqfrtV5x6rRTG3piwu/jOUpqHgHnmPkq5MNTf4SxcpgEfmLzijF8
w9C04zH4NdlpqRJ3hjMpTKru6pwIGSklHkssivrc6mO0ylWuSFYxm9/OK/ACzKNItojLuHMaGy7R
a7hi+K6UW/wH8pBmkm/0vNNQ+3pToyaIcCxQwKSQTM36eiwKfXSkqDHrIQUT37uz+AgHI35jzxKg
NpVZoKp/JK/vwQgtP/uFa/5WT/NwsEYZT7E9nhWHjhQ6yZms7WOhreCRvAKLZxVxno0DC3QDFFBx
NXiVx5VDcyoLog73TmJqk5qxJsYvtqDZxxDgZFMP/vxT0sNFDNY7ACT7+eJ97FcGR2Rq64c34x0i
kQru0zaPIyNNI4QraODKsxcVdkmGXNzlGSsA2RxQHIPiVSoeyw+qZlAVJ7Ni4623HF9XHAk2tEZE
HhqrhBFOmrguWnoGuhGm4rvFpjcls1pgedjYqa/6wj2XOPyMnoEJWtyxZjpHxJgBvaTMvMZiGmoP
2w4x8ktMDvBnHy8esKEs91QqdIbL+VrVocMrvf0540TwvsBsAU7TgBHIvdBf3NsH1MQd9iZAbMn0
WJ7r+6iKRLPkeml/bOBoo8t1JvpHEWFitpHN2nIF8evCrpT2Xz7R9yroAM91YEsbYH3OYsK0IsDP
v/ch08F/uHxpSispt1NYNTh9OTaOEpIVzeU/bhYFNXAEM7WRKv1Z41Vr8Q9d2NPawZj+lerj7rVB
yzKk/cjZ6WhRrJfnXcE4S9+3He3CGG0ixJQJg/VIARQM33K7Akgl+Gy0VHnDM+AgXKG08G2kw//9
zKgADKmlxQFgrx4nGiAb9vYqV/eDyoZBF94CR56d/kGn01KwILSYE3eJLhuslsxhMHlx6zNrPUC4
zAwQL4S08c0bcpG59KgPOF6mJEBPVBsN1PrGN9a3CfsYoWQP4Xp7FdWget16F6109gRAMzEbRZ+u
/6HLCtCV8zMEAf3XOGXEzJ4/uvruaMNcjslPmXmEyAzJnuCQgmeHn8Gx8uegDHQ3bOj3KXHU1aTM
puHh+55HSo5vq27BlflbzX456g3oTEF3r1jYb/bv+XVeas9MFKwxQZBqbvMNPspjaLfyw6ARakLw
r7NpJIcTOitAZu6OnqfUAQVnvY147WltLz3f4xNIAt1Dq84+KKrKB3IUNPYYhFE+KsIEnaUv8ars
V4/OFEP5DS17EAJ8+lNmyue/rg41nuN/3FGTthaS8xFmBo3hUzcmkXQZRSQSYGhpO4KVfS0nZl0y
8SKCagMNm0dsXYoryXIvDyb7I3tbzM2ZMnoIH59HvWocMtc6iU1Sl2rJ2HOdHCYCMh/FWqiIR5h6
4LnGFoNZSN00fVXuRYYUgBsEP1Q/jGGRPVbxzYsNHyxEnNWyOTg/g9ysYH9Uh6040PvOsYiFQLVA
rBm4NBdlozwAaEkMxU65B9hDLelmyG8hSeax5CzBv/y89mUUn20F+tUw9plb317YNpYRnhUifxwv
qYD2ZQrKLUkwM3+oYw3862MZaBf6JjROLllidiw3oN+Pmu4bRf7S4JnjkaDueOJconpcsQQnCAGs
MLDbsNxDcqIJWD+Z+u1qn+eBXxXGl9yV1exN5DA2S95Na1c0M8jzD+QjwBgbts/uVRD4SN3/KJRE
E5t/QzwJ14O6LZSzq6fyZY6dHQqSgfyNj9g939aYewljVEqZtqe8LyLXtnfd+l7osuRD/Ug70YdH
xs/g/miXewUqbhVI0NVkse67XOs9pXmfIzVWbtZiVIi7XBfqQIQ8rRaxI1cVT9ofKTEAmZms8dgR
lZyThKqcnIWQICh+qnSgqRXg5VEsOdzFOC9oukPfvLyOm5KFRLVst9uFIhdkLTbe8n67HNLy54Ol
pgNx6zAXIiu3iliz5avZwXbbPpkKq1bckh6XsfdJgyz5XMtnaWXDr3Y99N38o6N9pTknRwJvRljy
DTP+K1dyxqSp40Ey3Dn8ODrGW6qwCRr6NUBiZS6MpN7AQBQYot6g/bOMgc81bC8hfXrOQpIv2Cdx
5ubVWdop8bwljWl3GK1H0kXisAaB+yge18xFqNm9GloETEzD5hVrrMNNX+tJPRKYHqPIajhTumT/
YSRWS7xiDBEsTLVkvWaEUaZ15+HCQnpApBJCXbtSq0b+ZxO/a4CPnP7yLjbrjB96mbMd3rC1g8jj
GPbKEgf7hovtuDdRn+nlUXb0bkJxNKskDl0Ub1NBVihJVaiogHr0miPS8c1/FNa1jhlWKmZTBbTP
Tesoo5mu3E1xOSJTly/n2M66Yzia7CRnhyBrwly/Htn/Ui6smWCWesH0Q0SLCap0FaR5dl7/FyYE
zKhiVGt3nZXEMp2Q8d2f5x3rWQoqR4rbGb+KZrWhytmI7U6jd3NWeRZ8Kl+2+9ZZvB1/BoIZ1VYV
+8lkrIixielxAICocKw8zFDbOYR0s+JMwKo7atnyybtMfMgimk49nRaubnzIJmQrpevm+fLd9D4X
cKD8JVZTnzC/NofWJERpmJ88qCsIFSD+2vY197CsN+8dOLrlUEfJAG7YWyppyPnVoDPcW7xN6LWZ
UPgefaBvaW7BIrlclmRfraDndyRp4UGxcrILmngW2OOj77auGwpTeUZbY8KNRfgCQGXZQXn5Ldwz
HFSZXbFSiTQfrRy3N8DunOMd1o2f4VgwwZfAnT9QebCyU5EIeHTVnoBJxUsSas0Muw1phOdq/hTg
3i7fFtcf3qPZtequIor/MO3dhgpPj1Dzah8LixfHmyvBtG1Euwvals+1Z4++pojutSXGEJWCQQqm
fKPz4ApAXhGrYBWRIG9Etud0kgHSGEbUsM/KQ8QU48g5k9yxouWrZ88c0BsaRwjI3So88ql5AZPx
cA0Mf/o4shz6xhgmxbAB97/+qiPfpu1ixRxrJ0fFxF3cw7ZAfB7jKX9SEwgEeN1f/51go41SHrTL
w2ehAuUCssN6ItyXJRHgWghvSuwAJg5+wR5IAV8e909gnRE0Bfisek6ZLI88vQtHB18jypjtEx9z
H3MmA6etIymrrJEnmfV9AFKwobQJqf9gjl1CnWq76CiB7HsXemqwisU4SIb3ffhQhI+QISGrS8CH
XC/y/wVnxVIQzYdmzzI7wX7ijkv9UeZP4qNzp9MPvv0dgSqglTHw6KH5Z6CevWqj5prZ2cprfMJB
eB96sFOwozv5wNF1e62AGcDMxvs2Kdll43R+mWRPo8qkIrOy3tTl2f7p+nvvuGXNDifmUje0hiGe
Pkiw/IPMsZ7MVWfgcLNuUNCIWuYe/Yg4LhF6zka4kO+9/ga5mPH88FXpv9jtJOaYgA3JFiUiQ2IA
+YULUUQvASB2tP20YTnHNkUogaKolZEwqrVOyEPNSFz9CI0weApfsDJLdTW4yMzpcXoo8gQO0WZY
xjDRmeZBNhBICLKOr9eo2SeHdJ7K+WmLJBwkqJQe0NxXcexOXvap5zacl7QzeTqPBvJhRT1Ig73v
OnsdPO2XnVXZIh1cIYeOGtO8rVMRhLnKZkHgDtMYdjcNvl46irlwog1Xk4tab+Kywu2562TY8eQc
5wj05o+xJcw+lcBa+eV9DAcQ+dIAbH6SQ0IUqJr+WwoNtULIAmubZLVudtwbkwH58b9O3Td8zlsx
3bjkZwMBN4XxwxOuZNWtlNg4Vhu2WDb7lL6sGUNmNYn2t2ztMYIUC17w2eKW7LZym9s5rsZV1jt8
G/mQeBPC/Zj2gOwsyO9cYYzxoHEvghmvFcqCI7Lh6QuiruPfINq2baJSTZ6YErHBziJdo137OLGc
npaUR8CGNh3s+Ki583y+khYlX2KwsDeI3ZUHyJwx3FdOmuHjMDCX1AENYiWiQ7BS5ylB/15Q1KkU
Gx0ZIfUefMNdJD2VeS7pK830Xxne0GxyCYjN4QgWxWlV0OZ+OkniSnxsU5Rm1M66oSg583DQnRNU
10yxhuRzrkX11S0k5Wn5+t10+ybYa4+ehPU/P3hbg4O8ObUcWIv45Ee/QogyGhqCXC87G/7MeNRZ
r2iPusQvhSSYFH0tC25A1lZ9M4jbmvxzNn0I2IVoMEB9qIWlkKBJCXWhS2WQBxBGo+5UA9Vl9vk2
CEvOXARxFjkW60OK8IE3vs4c+GoelrWaxzodjfa5/yRX+G3i8/jtbesexZpWn87MBl/YWSv/hc6a
yuDu1SalLC7iSTk0uk9LPviyvGimmyaiVgVOF2Gq3uTgWfSnEE9UVbbJmlos7ocL87o7OLJ+JQWc
rn3KoRTZOIUaPmZ5aIs8Vj5kVfNjdtB6wMYzZaU3yQXJfsfcc66B7TErIhcxf73q3/NmyRAeTJIG
/APGXyP7Fj43ybWP0E5E+WvdhjSrq5IbNd94+fCh04IYWB6itvZUjUwwj+NqO9Vi6evCESgX7Xfd
z9H3lBRCuLc90cnXJBGCmWqWzR6oWEvFXqFkRvRaWtHffdFD5IvYzlQdBKSnV9DG46uVNiaGtGNQ
c7A2pzW/v1fjxpmIFhRtHZ91spEYHAy/rUEfW8itXqw0pEFvLUzJz1fyzgIJiQgdfOmlHhcDFO+f
wBfYzRk37UNmArzwQVnPjbDJrjyY9gqdp423oH9ZNXoK1IvQNiTRvzn27j63JmChpthZeVTddgpq
3dqy2k8+vyud1b5xH3zK4x/6msTeq235fhR4GMQmr/khbcXeq4QiiF6uCEEqH1Ls0WepunKfO75H
WMyO9USdzTuV+6ix5kxlj5gLMoc+VNQ/NNj+9IS07IX02gB1jhEAPo4DU7OmGsN+NHLBVTgIL8nT
dHuQZ/srWmvyLVbYMxk8XVnjnFY0Ea05GnuzwJRmIXMU6yTWqcpoUdytT19tj0bN5mMOmDgRbGQK
v3ssWAmkTeTtQtXnOkGte1FStIPOs2Krs4eTftrdaV0rJYjY4Of1r6gMN+MDVPOaUv/eIn4QCZQW
BmiKyY9sQB7agvY83oBwGPBrYXVuaumvNlXwEKJywzdAZgRhzgbXQ285cogsUffv0t0ZoHj9BL2z
khCXYvY2X03SPhZ0PQ3P1402wWdVSKQVU4sRrlJ4vjymPj+Q3yWWzZIayn9550SjSE13HkSg3c17
KwyykCaRr5WRQwmBT/U7v6f98v+SzlkozZARkFRkSRkZ6fjGHCtGaczKAM4UKT4SN2NlrHnRmYGR
A565ZKvTikkc3hKjNI5t6VAjsgauD3ACAi/tF0+GjNRENbLHVQ3gMwUccHGNjjMfohJDmEApvwuN
4OiJq2EOEeS7Dkqru4BvV4tRPIlij/361OV3j0JZvKfjS8BhoyxycbjibQP5c1rL7X2V/JUckQ41
Zyy3GsrwzmYoiqbMYv+n5ie2lX/bgJlp6aZGvMk1lASslPcnlRlytEVLy1+dhfyEVnBLgY7JRntX
4kHZzsWQ1l9X/96FyqmpwulMWKQbtrhyBfpB49G82wjOMFoFKZUpOTHQNWJUCCyA9WmwJ7O59Hea
Cy0emYeviTl0YMVJwh1YovyrbrYRE8Azh1GU98lKsm/HiNJalL4cxT0Rnj4RialLWK/E2Xz48sHh
xNX4DqIqild+wDitNNeGUVH/DNA8SwgHx4XkqMHJm4wwnNqOWcExVWdU+vQqNx9dk8yD0o/TQqfo
4KsWcjW//hBkKDx84Mr3kwTRqXDpTy0uqV9Atasv14FSGxtkN9PtzLaNQtDe3ZYLtovwzV9l85aT
pWezZ1gpR3Nisc1EPLbJEtr8vNhFuv5E5h1+ntFVIZVtUQ1lTsmhNpDVUkbKomk/MIS9UzFGE//O
C1WuYbsk11ZJqDMEgeP34Eu1CjoKYSZYiRGMWuUNaCr92I11fWieh3PXhZGvvQNy+/FLR+x/+G2O
8Y+RjR/JU88AcrXBZUuqwqJwIHPzOj/GtDX/sINwPKRNc+wTyQr8Sd5OzPzInCR+Tgwmwlt3rAes
J4XkydluJ59Rda/978Xt9K4bDamwZdMmASSeG6QIIE0W/S1IlCkbPTtbNDYwwgHaV7Incfw+Brgz
790h8u5d0r5epOJxPGbVV8n5tBAJb2m8VOWUOEnMjh5//sIWrmUTKx1CKeeNisw/r/xW/TW/s7VH
Oz1m9h8Z3zMYKgClqp6YIKMbXFqUChl3n/FZTHhmA2XHl2N0IPl6fbVwqutNoB/09tsSC9JhpY50
eBIIsh+Vq6c8IjhNk/Lb9SWRRQjHMz/TxrPv9X/9W3q6L0Dg7+ot31VxFp7gs38Ua2XWk441I0pU
P3bjxGtMro7IPxZOoZDOOqHbabYaCKUKyQAKij+kT+pGsV43yQDj/PUCd17x7f8tsz2O7LffRbDL
zeFY+ese9Dv3v/8FFfLWg0qWPfFxG18HgxkYJ4F64yYq7eTUwjz2qNreYRmhAiX8/SlO9SQIplvo
oEQPGfbHSMZtsYCHUqVq3Epo2yr/aEG6O110Y2/ZhyWZSFG1nUiqMnK5kwai7C8wQxV8keldI/0+
WHxqPOHBv6bqjbWxG+EgllrAaYhb3Tp0IVMSEsgz07AbjwtF3i34xfmac7BmpLn+8dP+K02gHAJS
mG0Ef4NgPGcEYKzX+NObKuGnJhNN/5cSMmv0MhWVuys9pW7kXa4inZiuNyESYnfnpD14zN+nE7l/
t3V5xHEaivbseUzZZuV7o9+DI6kzDo0bM1qQT5Pk70td+uU4i9w5zU+YBsuk3b55f6sEiyEnAmnh
+5dEwOWzYiQ+E6jPLq9k7Mzs37fZgkhw68XyPQkQIX0T1SfIywQa/K5zWxIB1+BorubrN8NFCXpp
3wbqCqgHEX/aUblo9I3UiGQrPHGAg7hnpHND2Y2Eu1iKY/aboKNYlTVr56hr2hNgBsvtV3aU602U
l9dV5VZUntqYnJwcPx/J9USeLaPyLqoteALgZE4OkNLRIT9MkveISpEeSqvezHxKwVng78GSg85/
7h53K7k0CDq7rF9rv8piitIX+lJS8h0aoy284fTp2KDzheZ+4YLE618v6S+XuE2cxr/DNZBo8T6T
Xgh7wDCKQO5AQUdBd9zVgYAGO1tPuWx63K8gH3hAvzb5ILPUTwmrVgeErG0RCPUcVaYPYyttn/dW
xHlMFHLtJ1cDVRWKq6rRAophRaRCduP+ElNr2ZF/ZigwnEchxJuxLyaRzviHEEtiA6VNjKaDYrMh
U2iVhGZjn8IUb6DQbsjDw6VP5NN4tofgy0XcfveeDxRDqlbkBbUY5PYI9v+L9M2sItFYSbB96Yku
MRhwrZB8fV/n8fNsr3eHyXmI6wowOH1CFo/vj6KEk1TgEZlHo1EhM8nifo4Ds1ZV4R/disQoxsax
nKP+PPrtRKbagiS3JfQPN/3zA/VmCnvwokDc38z+O0wsNMrEVBeP6W7dMJTwU/OrIg8DbGxKKt5w
yFZXvmMCQ+EXqXtAPy/n50awf5Z/pz70U2JstBuG1X4tTglowqLByVjR0UpMGf/aR9QUvm0jMq3f
oYFeCj4Tr4UJ+UH27EzMvbFVgcbSmSlCwkxx+qiOhkQnp7Tt9RQ7SuuxN21Zfnko8x6A3FrrLDRv
0DK6OXTPZCtR4X6vFxZuGoG9EAWPhgLwRIZSzmaxsXghIL/8DGJIlZQRbM+vv0HLZyHeOK5i40Cp
1mF64ecMMMh0hpTKsI6jvuGWg/SqDTaFhUKazhtBQfbWGwwOTjdGECksMCuMudgUU+A2ltU0S8PO
BV7GAkmP2LtKmLTExevgai58PBr4CAad0BWQvpUHpMC3ObHpiLUvDyGpHu3Yue9wYflI0oxJ/xEz
oy5DodWS1zcgmwO/xtllwGyLhu/PQvzVYNQy8rHWZyBrRJYdv37lbKpJ2AXzzrmuZf/rWjwHfJDl
MWfIywJnixP+zHejSVDGfRbp+rqOfkB6Luz+j4BzD9Lfpin23hjJ90N8ZRpdfh01qXqAGdB9QiVC
cOGNk2GT15EG9FHa239I84ovs9MSbDrBgMKJVyni+k6xHPQ7S4JjE/EsArlafTTaVoHG6lQAtACU
GUdgJ4J7hoDyqYu855PsBDvYC9kJNy+0uNXA8Spfe3b1wr0h4hwDNZuPMss7/MkoxhGb8maU//H8
xixy7r6RfEudOwNiDidY37CVzVkgoyyhRykfNi4nbuSrsVwSnzbrZfXtk0CRbgDyGwoVAyTbOJkq
46HnRC5b72tPxkDbq6Jo4adik8BBxiAW4QKyb29LJDzzWCau+FYxPU2fNX3OEI2kc4NSMVXT4mQQ
UTFNooCl6toUa7XEOevTRQxxG3LO80aoiW00V90G4bSqE7Wpy/hPZW6yzmpWxnDcwebClmT2uY5D
ryzraYkwwD/vSX+JqUR6S+KInAp9n8LyZjwGZBxUW84CkeB2gemPhnJ+owV9y+d7BaDge5wSheqR
fPiLsT/lq05Tu95yDIwKz7r6elYvw8nJfuU1eNR6d/SGvvy6KrfW6n+dVis/IIijzcjhJ5ug0foq
TEM7bPFI0JQyaSZgcPQoR1HT57/36LKohksEEi85MQoFytFtdFnH0cOzeyDsWGgnKhHvtc5CJH5o
lgMRayd38ewc4YlA5jSBr2PPr5ruFULEv24UeSKIDAlAiZCYSsZAx4bQncZ0cTEk9I9xIXxHVnXx
2ZM08uON93iiHy9cwJ9CwP2lC8BLOm22EDxAbHrcxsXESwTXXD/nGS8XsJKBFppDXUgcjzVM7Ma4
cmfsTjbbKhR5HBpt7d9N8r8h6d2J5F6dBbIQK0VTubCLcgEC3eC82nutiFehx4B7UC8XMAtN0p8T
5VVTlBBcgOkUaE/soSUI/QqZ2SaYBDXIIjnHu6mERSID8bcA7U81qBx1xA0FC2v6g9gmDhgqw6He
i5r897GJUn5Y6I+3r3WK2w7OrZ5+dPqeM29ME/vBr64SNtzOpiZ4W7vmlpqbD6tcxqidc0QC1mKF
ZDMc1zw3icCCu7j3wwnGdfYJdTaS6hja3E/eQUaI53JQP90LowNBwA0mPACRzbcatHAUOu3WF1cb
vQIuxUvm9r1N19lo0RvSJ5ED4HdqtZ0+6oGAd9E6j2Z7B7BFudFJj31mpF9TUFIAD1h9CmKZK0h+
NaVOqh2X1DP6Or6VetY7xz4DJ51205LEV87b8XcAPzNAetT5fcQFnIRVi75Fi6cNf1CnzDTdkqh5
nEWLcM+qvcZ5Zr0o/DWLHn2BmAhvjBV9S2surZBsQEDi6spVA96E4QIPDSat7HXajJ/VDZEuF8Wj
YXSVBPSO7I2nfD8zQfFFHpoG65wWj7NZ+ER0cyd1AC+bpYuX83Da4GgzlE6mhjunh2skAm0Afd2D
P9fNClsih6DIXahQqfqBsmTcwdGkrBBcBenInZKit7p5cJfIyYMFcW5Sg73biBWr4t+qBjd4denn
Yi6oYMWnz/QVdH0C9brUyN2Y9TFUM85KZajaDmrzGkRV1w8oCCjsFZ3bcSb9HrBRDpEUESHf2Y1p
xvJM75GdylT6lDlyGSxJkHlFPKP5NIEYjIx+kgdeyj5+mPkkXmIAsM7NONtnhk4WzvgZmmA9CddL
EfWr6tUfz5dEg8LBvcbx/jO521Z1Ld3GniqSoQflbZ9nFxRNncIxKUPMPuQbnM5IIIVQPNdeVo8R
TOnl2SlyRrBA4Mm4mWUrTeSgxnGp1/kbvvI7Uh3IzmMDzRGzJN1kqB6crHR8I25jVepI/TvNAxRq
S5hKoozy3BCHQAHAMCNP2SKg1ozJPicELqGK2afR3bdRdWXSLDOuzss9ugov9QjDaamJnAF+JRrE
wxreaePYfnHelUvs8J+HnxAIeRgRJXjPDN98/zPrw03ym1sXYXvAylCaOyee1gyeKA4PwGabvNP7
3kO5+nQfm6djsjuELQbTQ4K4EANRNQtOE3lpMaQt73GSxfST8dWd9+gHwrBmAn/ja/1A4dNJHOaB
XYn8wucFX5Z9BW8tA2bt8/t3wBK7rcySX7LTP4chPfNIWiCGwsnzeUvit1uHlB1zueGPZ9JXERRd
B4azjoqtCStbZqNtrKPGymuDeCnE4EWu8FcyQ2C/ccDSzI0nP5Qx7dMltXG9tSFB77PrnqaWIuTO
/1wx48fdo4X+bmm/ttpMgVbKv28zyjP/4dz5D7886rVBGUCsiCq5CYO5yt8HtujpwH3sJ6u99rHi
R8WoKkPpSmb0+oSFi256gXAZVNfCqmGu1omYRvm+zpqIO1ZVpLqY1QlL5D50RmWXWODLCSmt+U9V
Os/R+NzGN59690WZ4iUkEHIG+cGq++s3XjIv5Kl+h8Y3Y/yBhmT2dO8HrTSzGAVWpgK97IqSPxQ2
cbaPH5RUZuoj+AsdjKvLokqE88phbFfM5adVqHLjTt6VWTEC1bJ9msdejEQkjah8MBiGOM7/gb1g
w3iH5aiJY/jDQ84C1QrAZOVrQACgD1ECmGHjkTUg1eXjzB7rjbi+cdiXXZGDiisFp1G3+HejlvFX
tWh3VGXwnmUGjL9F9XLXoH0u53XpxauNoHtSSabzaVb1tPUU64/YfeXb7lZLykHi5U5HmYf2i1d8
2DqwtFFI54mnas/YNCALUQYfb9A31wtvhTBi9r0kr0h7IbpTobgo8C32emjm1vwuvMHxjCBB/M4r
6bA0aIURSPYxMbP+Sqx98uKB4z9k7ieLJxd1s6Dl6DnoXARO/3ucTvL/SeCRPvMSLEl0r5EvD6VF
J7o0ez7CtJwBM3d7Zun1iORUSfmiY8xTdvjq3HNUijWw/i1ehrtQBbl4PGM3IAhOUkup8lCK/9a0
oM6drnFzOYWwr1mrF5TdqnMtQ/zN9xENCrNIrlT9G7P7aCpbPvHSqPeKY5AQ8PWsseL1OMax5CYz
th6Xomt51xdXs1U4IM3E4jbHctoBgjlei7JmtnP2xS0KgenLk5+T7dnwhe9GNnhVEGhxlli2+Hwn
QKJ0yrBr2YhVTdNj6XmJKs082xsw6AiidqRHXSeGOD039tggHec063fH9HOo0O7cwQswHcqEN38P
8tGL0XEQg1MDfQRMnf1IBmx3tj8SVOyzWKWC3XuQQET+v6K8fVMDCky5r2quEV55xMyunmM5uymx
NVv9TRS55CxXVkoky5/EYDwIO1oe8m6fhUXMuPxj8JjFFC1HjuLp+f0jfErFhXirJc1JWLIA2lo0
j/urY5uekQ54E1dzIbS3mAb3etRDZL06e8WO5xroRfnNJcBbc7J3oKhk2xaBhh0icEPnwD7nOfHj
EXScmwkRyPWsrLr+qcNjyatC+mFz5968QUbCQQQ6Dms8fmSiSkMYMS6CU9FA1Ty7b7qeqWR7UEtq
LEcattropx/Ewf3YLaqh021ZpzKFu0uevvxU94MgVJGJbTSIipEd/0FciuYtd357VlkisBRYsKBz
3WC2fTPCy1Ejx5qDAw0NKe3UgPtK4cIDR12csHwcPscFJPnVaRC8zd2jFUUHQ5AWGw67ZXu2BxG7
4zA9Z8Nhi3elcGP3rP68j8SAScD0JQmp9V8D1xD7bk+4584PunlOBkf8rtIQZxrAxxZh36zqgjyu
syH0N1Cl02XbdeuffasTz+4j20OFh5fc0nnS0FLIV82mshfsIs9BlW1ALchC+JaEPDqpKKktXG+c
Xa20NhCkUaGQFzhfFpiEMvzZWLB82KjsQtJ/l3ZqwEOnTL2DyDGK3eRbY8RxBkdBbC3JfOLtm2Bn
HE90IDza+amIgJTJkHgO9hlzxgO8P5fa4D6a1al+PAkX38bYNmXT/Kk4mU7T2RsodzjfyJBxKXBa
Z+e2OuLKPeuZNu4iQ2t+FkUketiU1d/Kq9Pg4U8tm0mCPZ6kqrvOXLasyzOZJ+NWrV9CJ7oMUZIJ
lm5BclwF5pIYK05ZU6mWlAlnol6HVgqGLR4ZfvTQgIEzNEWnTse8eRrdV3XnTzlKsU3ONH3HhoK+
ChRvNRrsWfdB+5tfzKvy64OShehAGuDjpWrw7voIJ9sOzN9UG41mwaCBev61/unIlsNBqutul3vp
vxhVD09pDizB4HvJ+WbDfksuBqYK2saDsAuF+8Y0KvHaKXIAFOgonLWS/ZpNAe/R86t29tnww/nE
BSjGNsN/NO9xM6gDQB3cztUTEMkhPM+Y/xJTGDZ43BKKpacjYwfjidgNZAYZV57hcDIDGrbcd+Y/
jOXESzJqkj95UrBEDjmWGqPp0ynARXvq6o1sz9LzalpGF9ISpWmuh2Q2CB3END5W60Hi82ocOe1a
iz490L/TVSX6ANuFN7slVMgjJY2kRqN+3LxtgpuKuPr9kCKzrn2vWPCHh9hWYNUvSKGFmkBvJq48
AwjcwGraMjrZ94oeUxFEuhBs+J4na0CXUowjbSBW7b6CKIzbiwna1kwfT2D7ZusS2H+cRg8RD1rS
jMAReAgalitLndZVvfw9WE+tLI8+sfGvKQVwhlvMczdnZr6VGogp+LrFLSFRn6tv0TuPJBHB4zfz
0TaOzdxx5HbZMxTZTTuLh4KIk0n1/8dREQucooI5craacCtLH1shba+GMPr8tsvYWPT1sNiQH3/Y
KbYYueSsEr/uWdo1FF52PL5OnxF+rigZ9gMLb5guBoRvHnNT24eTR3NZ1Dv9WQi7u0cR+fuOcWjB
hElin+P2sp+ShaLwec52wrFpb/VUDqlEBhlmOuq2CrhWARD7kxGH1SxbFmPvmrKVkBgxBLGG2A8B
+t50gugbqo09cNbffaF8gY5c3Foffn2mIoHHp4ng7lUis7/QDCtplnLJRyZa/zQ/ggNrj7QL4yWI
MmtN//jR+7CuYrIg7QDyFKUjMI57wBnO37w7AQm7nebPhLR6t/Wt43nnqEWkGcpctzuc4FotEg97
zLLJu+JopC1psT3h9bPLGVhTwy4E9wDC7adLbBsoPdKeKBMDxknw+/h4EhpzYvuHIh9bkR+0Hc0I
F20heDKRz4dBHKVCaU87bRFe5R+VcDO7GIJfgdbpF1MQ34UHoqzHGRlJLC7wy3PPihAcDiPpUSv3
ubx3DamZsCRBKaDVEAeqBscEYH93/364G4OJ81xCRZWxEmQGJwRuu8Qqudd1dMFDb21i+aRPcAZ0
jz6giajwjxkomn2c4lWHK48WMVdMfhnf9EZXp2BEM9H34fvs/XfigGq2Ib+RHyVDZ13R8o/OdNnh
fF2aLzSGRuSLuQImHRq9y9UH3Lkncve53cJg0pnMJMdOzxLtvLhJUTrpDvhSRonB4NsiZeoTZ0fh
ymAIJuhD6eol64l6djOYxCPXf5FEulykKMogMWXSJaPuOtjQAm6klIX1mRyfRIqAZmFV7TqW+Chk
6sxDOqkTKEY6wJBZrdxJL6P3em346suJSvK2rxqDBV4IZUAuRKjFmoMBIPwfcIA3Zik4AOK2FR4w
xsMJ83W6ofQjL6Y8BfUYvrVJV9p7/JxHeV65s16T0bso1YIUdPTxJFA1pm8KidzzVi3nXFQyKxLK
uG0gSb751Q4Jzrtfym+erY9l+FQTzCp8GhzTkNe/zdBKL62G7tYexOUmEonIjr8PfKIpmuwTk1Nx
CHmvwfVPfmrhdVFxQpUlG9neXMLMmUMOcFPgxieox+8KZDPZ3ZsYC9K0ILAwe+vwN87WRMl0kREW
qcofvVDzlBexrPzziLd5qEu9SX+SfZZ33ZGbHXg2dM43AAUkevTQk39Ycl+wXkLdoNKgs2JBhPRK
MBCTqyteElhXONZc2Lg1VkLT4y2Biio4A1gBKBwFF5/du8GDywl0CMFsk2cQ8yMJ7ZtdRUjQOxcC
aGlO5NNceBzTFcSPQFzzO6uc7lYMKV1zbgO544Qya8NShDhKv161grstiT+PovzfYqeM9+UQ2mZE
RON/BMK4lCLGrKQjoMMefOq7zdSqKoM+IDdC1Z6T4/Jhx+VH6gX0jIkuXwMa61Glrdke+mCm2AYL
6Px9Gm3LghfJMFzCBpF7xZ8SLffMSsiaaFgf8pLHENMSUelVhKMkQL7yUcige47cQF2R3wkrPPEo
QQHIZbnZYfPpiF9O4E4UFY0C/ATMtetz9O4BG4LWjDjW/RXOYV1TgUCu4DoJYT1IYgNJQLqNAcZa
RIC5XCo1qjyGf0PKlr7cKO/h7nSyq81pu9+ZQg6EvFt2KraBLy1IlBB0D10DpsgOGJBpmgWbdu/O
lLofknxh/2w7rzuuwPcX5u5JcED6wuYVyOiLEYn00XlP26U5hZZkkaTbKbtvBpgbJiXN/pb27OZJ
8nBFep/Y664hktIDwgW+HoQsfyjxvk80NcRbu0HaevcRAT6nU/y9kgPZ2eskE2Or+lO5OIETmv+8
hlMX36oYS2hf/D2TpirRASjP1dE9qgOwgmXeP57yYU+kcuvP0XeqwVGRPt6NFdYUJUcguV1KY8sJ
eEpKEIgC6fx9AcgsqGb27YPjki7oBP9sGAxveXlw58faczuR/EfLmy7pNQT7UIww9PdYWwjhZqBw
/B5YYNfuDqd7gZRSzcflzlGRci0d7pV0LW53phqT2Twq+wH1tnF0i+iGJUoyHXh+VqqYT2VymvDo
IrNF+t5SricUQOLLgpltNTGBa/9W8osvTjyw9t+ure7e2tXbuTdzIybQfb5ql9K/3eGXJZ2YCIFZ
tIo+vqwCMOdhig01d8D2nNQz1K6HgSL/MXAm/oQr6kDrZbs1OmCOHWcMUo6EFO66piifAxnYTaAV
Ud29R1o60qE3pgPVuuRG0CPTMBxWqz3sNtDAFyC0kEJOqcJwTrlUuyoklkXBXrJ4tqkCZQ9pUgVs
6qgw76SWYMXlmyN47nh/Y9T7js4OcuV8pNf/HOdQjOA4xd76qZVKGN+MQXb0CqAwUeMIzz610KWC
/MpjV1RJSXeju00PyL8JZ3QlBcwMG6RblYEczbzjTEVNi9wF4gGuNoupfFhEVpJUOhUWPzLy5crc
g0WBWoftbGuAlQo5ioZ/MjymfU6YYygefeqxvyBJCam5X8y3Qs0XxP53uq2CoOYH/9lRVZtlw9a+
m+LUxbHJBh3wXqkmhbc1hchq455fqI/Wp/sOfa2Iwvot8ROm22D63d2/kY+JaIU0wRQcS/zjSzAu
ph1JOITmra2iM/rAHd2rYwRBDdcF7SM/F1YLW7xqU/ql2AnqAugUD3UzhS3CER72X4gww71Px1Kf
kDp+xH1IETyH1apWEUXrE1lHB425R4ruO2ahxK5FrmHjIoQGmnr9wDsyVY8Bqgwvkg5PUlTogWC9
eUFCHx3g0YUACKhLt3r2raJ5ZbMMiyIh/EOKqBfQn10qfSCnnpqpHjx0AB8Dz7nDr1kASFXWwH1R
UZOjUQcn4zYF0gUO+hOKpKOWA81zXeptCJlKTsttpZPKU76Wo1o2dQoB2c1SYse8Fx3nRUPWtmqj
GPLO4lp3WR/P4eCmWrADlXEUcRLBI3gsWNgnBMzo4Lcn/O2/nB8P4tBl6U52TTyYR+WxGbRTV+Yk
AbE/XGNrAOimq7uM/+N5yXN/7IHH22tUXp5ZsPJaC6R5xXfGf3Sw8FHG1Nz51BlSwNxDu/Hmy2CI
rIqpwrKCaRUa0z4ikadQ1HkozX2zfeFCmVSHv8iMG5BSvVTSnLrc7sF9i+Sy9aNjO4S9Gs+OaKfY
EPpZpu1ai0FSx4eiiqzgdahupL6jqtIQCOVSJ8PNae0qtfgWjNpxyiI5X1+Wq6PIMnK2gzV//rDo
+wDXrwySFrqXeQ0H2XZpAhCKcbxicY/jl6JGhF7hws6rwYpOCXkgMTLF+fxDUCTDI08UZpBFm10e
qSWofm79hpBHK4+kyZdYqIRscD6QHlKFWu04DXqY84UtWWZMG6zZ8BAXz9srIVM1MP1WUVhDdAAa
VcpwMtdAywUBe8WOFYIi1pe9pru8C9m0Z9xFmnG8huzloOFnIxsxHMxfP9Vru5jmqc103dVGwLqf
H9bedXkvsT80IN82IKyQ7G/0QYJpJ0imQCytvVPEW92BzQ+aPvWGjyvPeomgIJeWpBDZZmyJ0CgI
vQsx322gJDhDsfalfCTsicSZDEKSCjY6t7H2xTiji5s9RoFqIpIhTlZhMvA78aLKWhdifrbAcY+l
c1b6exkoFmAoLDKbnEcP3228ku0ds9SOBHHH0CrP/wYaU/lUvVcW/qf3NE2UNWnxI/TQMZ8tCDod
2k//xbrUi6cZNynC5StbFg46gMtjb37lrANwAuxTq7Qc9h4k0QlpuoXW9U2vea9E9lrAXb4iSyZ6
3Ztim8+ZzP7dkPxxUdsQF9AcodaKfX3+YbLFBwWzkdiLFxCAztkdoJzMa7Nt5dyEktd/sB5h3rqt
fPROZ1Jv0K+mD5UV0f26ixd5tamCKXeOv1EyrRsK1Rv9uphjCrw1F1WIv79ZsYwN27BbXBl3AGci
Cc8JdPvJwv30OCfHLicF1jSmMgVml23Rcs30slZhVBvuSoclBycmUKsI2FhQ5IbNbrjXgcZ1GTEX
H9wgOjSzYb87CcPm+RaVsLhd87D9f5vg3ovTfc/CcBYPOVudzkh8dP4n9cWWlbSCtR5njkSX8hMP
6kbfm5qp++g3UWJtCLuUvfAQ5vBipLdY/HN91mwu9lbZ+pe3dEvCR8cP2s4CEY7hLqdmnVYOSDtX
EkQTciLtPxuoqwpN6ixVbI4LOWpAcantnFQjbbArkYL29zWYOG6BmttYWOtV6z8NLWivM1t85mhE
NCGprbb9wBbNtoXI2wfbHAn9yE3fAC0AVDnxXRJ6av+pRHHTMZvpwOr7+rV5XcYbE8bYXUU6OB+f
np9Xa6O/3M9pqWjlj3EwAdyBXA8XZA7N5wBSwoiDr4jFniHesVTIUU0apUz2mE3kr3i4Ktmn9mw9
kWlhQOywrfzAx8aweofn9cd1EJAs/AxB8M1Rt7hDIXvVLHFIfqYt5Z9E5ON1a0CaxsCp68IptzBk
gHdDvgq1sFw8LSZuKn/XiY6LJbY1TVgS79WMnKRQn7aH2bxBlUWanQNn9GRK+Dke/yRIkR0DmbqP
2GLnC/Kvy1FC9LgaqRhn96uGHHfafF7Kqtg6wb2wYucgjyR08Fo7KwQ6/LkW/93ZrZGKQBnoj37G
0DmfgSZRJkfUFv8GzvOLvEL+Z22gqMnMmqJseptQOt+Ee6+bnq/BGuMZsAl9/GSSVEiKZkzDKO4H
wILQbT7gK58v3QCyNXFq0VGatwaiZNM0MD1BOWHz4EVEkPKQe3tF7CydgKaNihNPtvKI1TBPEry4
xPSxA0ido52u3zftucyR8NxubOKQV6APNW5HGG13ukdzxj01/if9qXTo7RaRcXPLBQCFU3YP5oKJ
UQotLjsGE25bEtFoeMxnCYTELjK5DnMNcZDR4VBxHCg3EV9gg1LQsiZIeJoyuSLGcOIv0mVbk4O8
7dWlg9/55Ec+bdpZZQiltQ0MErsIvJBnIbno5BrkvcBvtPbC4LpHpu11jCNFMHpa8tVJK6V5T7I3
Cwu+vS51Qdap4s0uvetKMQ2JUivl7OsfRknCHpINqZ4W2E1Rrnf4JKFICTN6iZiiL2wln32NOnIk
QrPXa7biGEsZp0UbQiw3d0kBFLEG0YZj1euRPfGEurWQeKOH7L3Sy1jHz78avA1DgUYrAatXhK46
P7j+vtfU9kOVigdm2xo3e4a2zauWo/V3BZ41UIupOFhRRBmy1yeKLVQDrUZfVcd9kSsaDWoj/1VQ
+Q1VZ6cSwyew2p8Ek1GG+PnItkqrGcvFM8Rk5d+4wTQ5masqKxWO7dw/HK6b5al6pdGl6Sj20NyD
A1Yy6wpJw7wJPzDPBRHhSkow062BO0LTv9fGUZh+v1SmEAmgzKuY8GT+kQi365V2dbOWbt6r99tp
49eAJAseaBiXQ123rxuDN+0qiP4j58jdmG71hHoHlun9YWuApZeSv9Hir7bAEklRpq9EknJaX3ND
GDBc9bLbiD5POQ1FQ7rKjXht/0eb+ZMQFimdLNis/T3v/CYTZeq5LkVdhx8WXtCl1Xm/+mIzKHCC
P/X0rnfwvqrT5zThl8uAvC7pMbBvRQ7VWB1q+e880OyR+ATr/wpBrT+EheIAL4Z9xz7wcxeLAKp8
82YsWlbaFhGIwlrhDov/exM7xemT6xQP6gFhJdYJyDrSTQzNCvL2lrFA52Rfr7j8fYLscg6yrb0G
R1dnFX4B3B7hP+/YaC28z7ayFTcktO+dchZ88NeZX/Muudq/q0tQSzQ5G5fTxl2ZgmFxGZTd2mNS
TVhoYbXCFkIlqm6gjtlweKD2WlBovUjA+fjN48WPSYqRkvxj3/CfdrZlKb76/Q1vHG6XV/c7r9l6
TmuRtGliS/kqo936kzvSouzJ+Vjprrd3QKv+Kh2/t6UZmSr+r86CXEqtML8oNCuhMzNGk0R4zZey
aj2Sdzp/xyPkjKRsu28ZBGluNszqIF7/DIdpsFY13hoFzm91TkzMQcr96R3ad3/ffImsmqnGEJj7
wXxFaQWKL071ZNWxvLAJtvL2XBq9FQu96LvNFizd5JA60IKpL29ezOhBHaJ1LE/XePQnw8+Y2cUE
l2p+D9/3X7VA9kvRnKQxY9ueJg0jhnvyjyjo6smqN2Hw2GB+SCZu1B5FFB4r+r/PlHypU6ZYTju4
VoTGUAd7WJB/vvD7QccjtNeqwEpX/7PJOSHxohMxI/b3LCJ0+vMFMj6fHRVz7ABroqySFfdi2WbK
+oE95iJQiV0OdXFRh860tkXkYjqELGWyZxUZzSpVJ2/8JNUfZ2PaxhY1kymjlev0rQe48PnRxDOd
xlmCdw5d5y/Ej8qtPg9ww+FDuRMjSY24lAlfLuT8YI1uzWEjEaZTuBMrcTS0o4v4UP08FutlAP/f
+gQ+ax5Xan7z8aCOxP+DSq0Go13mwLd7mEWQk+Tpri7RAEjzp4QYr2KssJADCIMxytRnV+HjlxAv
vdybe5riw7KDAK6YXsttqZM4l/Fv6AAnJQwgJQkroyjmP33dwc4rfubSRfsxJALuIpc2gI5qd0kA
upKCCxQPk+/noJjoRc2ok085cmbTf09HWItVoNndcEsBSCAzG7O0w6y4u04vsikqJIvvHzaRwimK
Enwt03eCsTuwNYUobw5xQanqTdDOsWX7oxqRcczXbeawXADa6RKr/QKzq3liEAxFXuSjinEiKaKF
F4yv9GHttsMZLd9gimH7sAeTPRAccpsGTuCxMV0ocxcl7qzHJyBFRYUba/Qdh0v4DEn8QtVcytio
HTL4YLg5N5i1UEarKS/03vcFIx+XJOSXt7IeCWPngU+ymkbQhVLVGW9eoN8bVyHnohlTZkuJtvEd
eOxMSnSUdmXu1sVKxj6srXI/qk5295+NHcGCLDsHv5oTb7YmAhqMJqdexAEW+EYcz4g/gxvkZbAi
nfnfRBwXsJPLbQf0bbPlqoH1/YapF94AibUdhUuZhgm5pzh+mg+gLnWe/GVfRRholBUzOSvFcCA5
qR7jjXBKLEGKbtRsODqI66eHzWIjLR0ilqFuqcXSm7SQvELO9e61+IptNvdxKwSfp8icRehsiZYw
sLxwG08GKFxEb7SZ6pKgBxNJpX+cNBQ9X7cH0vaG75ytiSmiC8FTO5XpWMJ83ltxyL78OWA1QMl/
0Ia2DVnjPYZi3xD8OfBar9GIv/iOZ4FWcHVWDNoPnfd1IWBUuwYM9NoBzvguhyDcw4FNfysytStU
FChC4IFmnUKnIQzq6HdsI9wwjzepAGgeNLVlgHNvbB+f7Ua+VZnybQZpCAXqj2qFAqvuP1u2V49G
XMhzg+OnR21GRfmviGyCg22HCIUX2X6RPf4shBlDISn1Wpwwg5K0OBzbl55eL3gAx2UR833AGVlQ
Ws2wgRjG7OhuetWx8Zkqp9LQAzn47Kg0FKI4jMw0YNMZ29FJ2oNNaiFMUQ7WadJvKtjtKVgKGsfJ
Fd4jwRUf6wfsRT1dHHBgbhP/hLb4WmVbSoKgyFqEX0D+BmC5PKv+ML2YFlOrC/T6TOJwCQ99jCzS
55vHaXd1bBNItxtNOHY4U0YPBMldYqFbgZ77CsYFtWZoCN7lllSSQobov9Hp38hWXb+OHfTT5plF
jcnHLvbOIXZMU0oucd10T4dB7RzSmtUziCl/AAEGc8IhgzBuWbdsj/SrP7AdVGbthpqAOs/YPjvm
4Eo8UFwjzRHdDRFkvHZ/1qCTbm3u4iBtdgeBxoPijWR0r/zJbnSI0k/GiV/pbgSYA/dMtX6NoK5v
F7MW54zk6xycbwTlvFEXUsfu5wOFqdvthqcBhG3Z91KPr2l9VYJh5syPTmk4N1vPUaQOD4057dcd
mGMYLe728Kts5lua8P7T0ZC2JpKW2//utX3cr8WpQ5Y25KtJFK+LCE3xnimNC235jubtTdJt5Zun
xEGHONXqGy7BUsk4D7N3ALxRPoXP0gyJsE5w2Lz8Y3vt+2QUsD+xeCH3fmDLv3hT4rYkbi4wJ1rx
tDWrfDRh+kH3lfon3JjEhIfTeMJwq/9FSJ0oqcZKFo02rVjXS3NBbmvsHAj+YzoWNKJm+zzhTt2M
TxjlliGMZdY+yG+glwWIPzccYaza8EO4ghjrCQOp8BRjttHm2X62ptNCh47J1asFOMfJHcQ2w8Ut
ZS7H+UAYFSwwi5+NlIuRm8SwUw/49bQ49K8gVsE5N4eU8zOvXKxcqN2B5+WIX5gK5yHBMyyny/BJ
+KoJvW33NytPSxF/Wh9u8zrX9lywfIWFR+e/hVzRUbLtLjdCfhZXX+oXQeRCpuc23bweLmwBDLMs
evNbmG5yDq6XJe3R7ZVLx/WvFfFiD4a9q88JjvHRMY5S2WpWsyTXHIjEzEHeqThkCnfm+KVUagSF
SjVzzkAz5v2j+5A0CUe1iS++oFXrybKVO42t+9MSXCrW0cuFECixHeLDBOUM0rbC2KkftokZpypg
5NanmUrSVGH25p4jkkCTQ1It3W4Hs2o31F2Yk0oF+eRpOjLWaXMYB6WRwpqZTvIBTE8igOdeIJ4N
aKhQLbMKIQzkN9Wyo4Hm3D3/DuofDnH79UnvZEJuZC8xyVJi0NBI1mbTsY9EbHoqZhABFKv7GDYV
bxguPx22IU5/B0EsbsitobPwocdFKWNV38s6pH40N7FYPTUbR4cC4zfJotZPsAHUlhF9GeBgHygC
oC/0+TwAb56uSH6HcB70+GOTV+e4ioXOLsphrYJByFDMC3RAsW5LB6+GzNZ5oj35qAT56OtBvb34
xE8zEQ2QoglgTmf3N3DBESQMcUrKKt/dm8wO24PuJhZsAZDhA7rql1I6Mbb0TIs3o88QgV2Td3eO
Tz6NKIM7BfadIUES6+CDFTNB9IzFj6H2+qTZYrNZE2MUyhQebF8hDiMup4g4mW1j4eQC0o/dpz4U
KX/HaEPrB0mUkubtygKC+Dh2kiqM/lwwsi0k0c90eZ2m6JAztOlDoUElp4Mfjex8J7u9a9D3MetS
SPNXjUUZR/5owTDzrUrbLLqBWVv3piceQAnXbyG19t8Nxcfq6v59tfD5PPs8wLpoRBm3PKrxjwKq
JOiBgyhdGTXK9o6WXCEfoayqPdNc05RtJ0j4Z5+1+Dilz8AC8R152wzmJCPaz73dDotzEoqVXwqu
I7ZXRA6OlSVX+Huv4A1YU69PSy1Aj1+nd8GTd+lLQm5n7odgZqlHshGL5t/6z/2YViq+sM/3wXdn
+WbvMI80Waak3ef08gQXZYFLiDqw3qNt/jMSPsMpEMTuYpXxhKiMduAtxv6nWwH+geHAQwMNaU4W
LRjnOYtCVBbk+mDYwCDlt7p8tE3tsWEIe8AGJtBJMQTFeOnxbj7LT8+FnMuddR9U3afylNwUz2uv
TkR3bTzFmyhnz2vhhMq0QgWNyyPTbO2OwMHCDKuu1zefzUYEa5SJ7EZPZ+/vWS95gEe98KOa9Anw
OsDZWbRBDmR4XNGIS5szIR+Mu7bWhCa8Fa4nsB4iHuyghO/A9Heqyop0M82v2aepYi6k8sjIrp7x
3go17+RxCdp2IeUQy2mXgfUm8/Fqqb97MAxH+ngj76UFE7+BPwL9QEiI3YEJ5jyzR/fqYQ6AoI/y
PE37jumK2A7doPefgcihaQZ3yE22cJEZNxaP9dDdXCdISzj73wMdzy3OGE673z5SStzbVG3ZaX4S
WQ551aZWs0l64s+fb/MM+aIn4uEZrTb0fvl0DJyHoSLsprnw72tmaE40dKJkG4B7yA8V3sF0mGKm
/0YfGL6xsowOYH+UHRez87lXwGBLtbqCnnSs0d2tzTV9pWrf986GR638K2v3CnZuXVDDr0yei3DB
L2fOrcWaFlvdOkk7l6Q1Z92YftHXIFUFLOzQYso6jKU1RIwhkFwWN1TuvWq4xvn/DjfYyuwDmrnb
iOaPWiHIJXx5Ke1Ptg2Ib493Rg20ftsqrpFor11ucgkdjSrrncEUQHLwHdIgzJoBg6lGDlrL5PWO
9YLp7c+0emrPHgsAYMGtYb/m9OJC1Va51lPkrMC/1w8dhmSV7LaWVzuIylbSosT6I/vko75ss58v
YQTtxnUa0GAbMQh7GaKOQ+q9z6aAvo5Z1djP1PRwsetJnfzU2am8QTGrp2QMP1QG+Y7Xgm6z+Rjl
KDzRTbb5QQPgPcLrEpbQ951nJE3H1GoET4Hgo8xYViP3sRWcuhKRL37fLLP+tdc7xFgDWkJ3vIXB
HBtlKrTWSi3ZNAnPaJiJ60oHdguOiscnhBFZfEO0JNDeMtdpkJfoNfYOhq79J1dglwOLUlF0o65q
rutdM2TJ2/huoGiUpHc2LW20iJcwqIKOYZkSvfFgVta0DJ6+NxrvDPjkvZIAUmTxYmGNb8S4SMDz
FQDalIrAAoGhYsWOr7wc4BXO+qBoY7N9IhhFJSywA4qiBUwa36QkESkGo1J6maaQVscjvNhlz9OO
LPwlVCMyZxPmGUxP9KboTgXTgtQge8TDJk+kISnlg0lOUI+r8T6W4EneTFsIJZ+HHnnwmaWNE0h9
K3fZiZZZeEbK19RPHQu+Qs7XGiHQFcY2499BnGlMN0j0YinHpNORCLUtexn90Lsoi4TPUQLQzak2
o1gfUIeeCo9tOe5R6uMWE412g5p93fB1bdt57HovBmWppIpMbWPJczFRxuhIp4xpAfroMeuy+Lhv
VPYQdr3Q5bcOXGyAJkUaFanrgr6qWPCJ86fTok1+TSPiDUN9KcC7pF8AWDpTtEy8kQd0ub7uX1vr
h+wpPUoUDnXyntb7xCyjFbrfUEY4ITv9Rvot8jpqnxRxpVuuXA3hoY7wd+mN2aEibVRk2jYEIcdJ
iLU0N6DTgUaNoFY/XSW4JBL7iPdxon3NjIEiMdra+5VG7cTOyz3CYkABipqk+9PbopGAtiKMLota
zoi9JMvYV3zA9JFw0MtaMfJql46++Y1HHwKAay2cBxAHk29TWWyf6Qt11/XRV0SkCyqi+PYikU0M
rDDJXDQ9PbmeUh/UpTPfSCUk+S7dDh2UJnWxHpCY41meshyFcSeOL9Ea34bXilOGwyZQBYDzqIS6
/yp+sdivgscNTujrpw+tk67MZ4TKyJWOTKa0+0oyDVyJaYH/Reyk3ePD+wmyAhQ1q/xOW/maJeV7
H3/01kBPtoWkMD0j9Py3dPOjzVcvxdut/cYArfKKZIx3CwftsnTTzg0JZJACe4PP8BfqxjSRc0D0
GU/4/n1oRPFnCXMT2s3Zl8+yNCmb0JLi5DsCdez8qUxztlOr2zFP2RAqORE6zTRGC9L6V24PPnT4
u2uk4/j9671O1wYSCnSaUGERp17KrH58xlDKKryGGgLUzN8utI5bp3YVb7YDluI9+/jXzQbT4w54
5KVqqP0Pj/MU/o+paDdSIFXNW9UrmhHBH9GEpKifgtv6NXiisZBzuPHZRpkiI9ZdpcL9Xljf+Rdp
zd6x8OaCNIBylJoKbEE6m32K8GoIjNNG1jmjvZh1FVpYcURM3xpHg2tVFhFQVSFD/mSTFpuOQxFH
vPHiYE93VO4GLXurMY26K4ZJ2Il4VC4v9sC/m0L+kTNiCX5/7Uo0s5zNBOdia3uwxlG08QoZDGrF
voLGcUtYcULugPyz7MZ74dJrZbyt4QRHVCu/+XqX7k6i4/bWCG0tzBwTlZm2iBcdy2l4swuSBcYh
A7pVKZZ3MnYJOl2+r0rfwVyNPHNuH2T30DtAEbJWA9FOIQ2HPl8VJVkkhHIs+MKriEyaB8T5oar9
aPhuxerTAPJAhC0xBmS1k3hlWAoHHMBZ/h8GQaHT4Gj4/jt8UKJ7TBJhA9KIKef69WvcaqYhDNdh
ZEjK6CfGY87VSbFG0qlv4Id0VEb0IsR4xe0dT/sbN22nN0uNL1MSErIgrGCVN+Nk/BqHrANais/Z
48/zN4RDErOSVwKmbH4IB+NmCRCoNwxO/snqraXhz4tjEmFUOv4Ws/e9hIITb9XtiBZlgfNq5oRl
uNUlc+zX7GJWqX+ZF/n3PScqx8CxFL+CEh8svRUZsNlXztJe9tKg225So3qY4q4ww78/83H4kP2y
18X7Qeh2Txt+HC/mixejhmf8QJJiDPL2ZruK9vkdT+g26y6mNHt8craoIptpN+viAGCqCL/8tGby
6MLiXqkPqvZzUYPHJVFh5cTq1/VGc3INzVJFRvTRMUvuR2mNBlzoKgMowQvwccFqlhs/Zjk/S8Lf
2Tjmraengq+R9cp2GZdWG9/uJc3xjW/tfS8qx/KUzdvG51JklTz2y8z7p3RIT5Q/+pKcucOgS5Rn
/YuvvEbodsQFPr8IyE7Nx2wUi8suAjl7WY3SNcnST9CGSgGiNHnMHoOXeE0fYH9Zck9pLB6x+zjQ
8bbKgPgaf4NnOPuzJo+aT+cu9aeFih9gWVI+fqKv+cyungB7jdDSidfSoxJKpukElm6jUZoAIxDH
zcS5KYT3WMaf9g2PTZWzlPuz7wsdpQu4pmt7vciY7aM/Q+BzILZ6S1Y9WFHrEG++dc1PADfXRBBZ
d64XQhoafKlXoKG3YXN5rhL3AMBNaNyUvCWEsn+VrFmpIKE0oFAMRehn/pXMbppo4g5IUXQkYBaA
Q+xxOdAmyQN8cHRTz+1D0ekzoTjqzdbNAweFc+ZblaWo6NXeLSlrgVY9/Y3E4zd7uivPqVWxZJb3
HIYY0TV3i89T6S/cV0qmwdbjdo5WqFec4c/VcPHzd1AVIDxtX4eYH8xkfH8r6agQH73C/BBesEGY
ZFr3DiwOTK1+Rkt2CPuLvsaVjaqbNJcKW8lo+b1anY2lDa26KF6VS744RTF9eiBlGsdebpBewJmP
uldUCibpSyrKQvAX4hOpGIPN93+q24HdZK/A1s0kNZwMhefV+7BlWS4lcpd0Ms5YSq7W/e9dFruN
AxbEEYEXAX7xvnCp75s/iMLDPW3qaSvPhOr5KzJISu8IaGwZIE/RAy08VEnu2UehWhZCMUynFOS6
rP61CWj04SPEGHzmdinAIYpgzgQULU2/J7isi5istiO+qXlR64K5hyyyNHp/NJsILXO1Trzx+fit
iO3p8YpTGEeM4Gq7yFTBcf38BMoMS8HgVGE+QGgj+VwBfG6FdsGGJekiqu0wQkzKu+/oO9Rwjedu
qn4NysJv77WDuGaEXRf47OftSsuuYvidMlBsQmtO/MtBifwOgr5DLEuqTO4Pb0TWmj4ATGSEVRRZ
MBL9RnlvzEIjHEXN3l1QvnlmIDzY8BeXubYx9n8xthDzT3lDoqb3iGwn2m0rL58kE4Ux1PlEt4Nk
JliOJdKjGYuoXno9LG3dl9mEPAOtOG2BAnSLDrxXowDPmRC68BV0hvFJZ5l+ka9jFNevhemWSSTE
/SssRINahg4J0UkAK+EUoKQ+ZGr/B2QgKbDVKsoqf3xuhjzk3PmEOS8EHqTYytwq4dy4Xsez/yHX
+GWDmrIF0zuxUxtO/icfAmx50/roilxffzPw+ugpBHo5H0MvGItjyyw7XodWeTii+LNLsSzmvo8a
7MZPYCHeyzCeeUzHmpo1M9FyvWil4hEhaLHNtil7aPUUSgoOVzUNNTepyXcm/2he2EX2mbfLmYOM
EMvnBm1RmFoBL6FF3iitEksEmdDcnwY0SSx7khXc466zIa5wM/ULISmt2PRGrvisN709LYXzQnVl
UqhO+TjMQbu7bO3VA9Jkw24ZufqXtinRsRCKuZtJfY/2vqwV4afoqTnNB8B7rZYeJ89e4YrJhYzP
4wXg3hDWEAj9booo/aHvNOpG6nj0lVdoLNVKBUkQ1IAB+zxbh8c4oj3BehbF2oBaoUe9m8VgZk05
0VSc+i5JzLAn56Kwd9a61h0K3LwxFPDtLD8YT2C2ReOsco+NEdvQD64CFWEnFTBJFBZXLn2AqEXu
EInn5HPhZAmeB8FC3TMzifc3maSJOUA2CUe6tFUhaOKJpbIP+2tZnyXnpQstE5DdThSfcnJaMX0q
LfKoN9cS+zBf6FtCLQ9msDnBpBykf2zcVgiV6cOzvP0PAVgiOApQA5JCeBH2ZC2/lIi9dF0v2VwR
OB60oma+aMEuVfxprMAvdnBnl419ao9+v1Zc53oIAsD1k8CKMlvE9S2K9p0f//GXB65RmkOOG/Op
fjbPINC5Uhjo43WgUJb3LM/vzkWR89E9XGtawygIYxzOBHbxDfK+qXRFtauAMoLq2hyyWD0EBNV7
cNhoznwhl29hq+nntkx34dZTgi2DKmQ9MHsNcm57OIDRQvWNOHjEfXWJO/5rT5/dM5Hn5/so02wM
pUZN4E2pXm9tSNB247sLIbI7rAsbO8sl58X8V0RavGXDm2HCz7Qordy4+FlXy46ep898NgM5WE9K
w9OMkmfJxzRUROeRXcmaMx2XnoCrK4Ug7TW+dvLL4i0r17AM7kTRGBEgIkNcgApBbTNFTwz2hFKk
vUVHwvREftRliTREm9VDRckrM34qhCfGi8XrcrNXESTVPUA3ZthlYUsk5klh4oS+6LyWstQGZ3Wh
9rantF3JwXQZLnlRu+9IPGvbmnakrlZ75TEarvH1Mp2NlpXJ7iQqp6k1alLqtyoryINXiKIHRLBH
div+ZPagd8W/iMvLBLPLuwe8S0Qtw32Nt3JyBFbNWVSaQmnBKoj6mKOSDlFKloaHpnW3AtlpW8m8
aZlmqMwFfVMPBntJ+8Ej/7kE3n6SI/ynalTD08tof/lddkr0WnqIUl8FyzmYj4y5Agfh8HT9thd6
K3Tjo0CW9ChFe6gavmsS4VcML9t/TDoTN8lq5E8mEDlkvPuwdpG30+zymy2FuyCMHmvnzdx+Vdrc
oVfNXtmpX4umjH3+HgzZ2Vqetjv62bCxISoohyqkvzWJ+2Hz/lNJRiZu094jFdjw2oPQRzdLSzKy
QwEjfXGZ9nBOGeNoGXZ2uPZUo8irJ9ScL5QJjaffAZVTeXdgkFH0EY31aWtadehOGislNmyV+Fsq
Sjd5LcSYEb8xS7QzSJPbqR3zm0I+Twp3XaejS0jtAhPiguBzcmah/HqFNHL0WTr5mgSegzpLUT2I
z8nfWHezs26UDpDII6Qu5ZuYa5oJFSPtmnjgoXvSKlkNHT92yC4Kjpcqu7DDoI+2g4liaxuDexQ5
8//2O2By8sjufRQYK77b8UIkZl6LOKx0Lr0YkFBvNQrcb6HV5JwAE8MIvF07FbpuhAWpF+LdUa5I
UHjewU7nMfSOsSUeF/k4l8wcI6iCKg/HxdZia8Cv7aLJm7P6TB/26xaKUxX8C1kb6O2bjpPvnMtz
tAs1UDbLbukDkuDA1/zSRcWY3xSH3QiprtMrbdh0atu+OotHfdeL71jlkNreUewwdiZrUN5vx5Xx
6IhHwEmFjUvJUGx0K1vHrvJ94E1ZaSiI652UXArbdRXbj/yXXaEY7SWKv8oti8FKNnBpxpY0No2U
liQk4Vw+vXZKRiSYFz63nw+pXfS4q6Mk9FEJSxASSz8iXLK/uHfonIwDVSFk7bUwhGINc6o8TCns
ZRfLUPPH/LFuBnuFcNOB0eL81iZMv1SxDb3jskKgYlvAYi3vKG1Fn4LLguKIRuw8VPzBMUCymfrP
i4uq1miOHNHF69dM6tJgIMZhwRjuJ8DPTl2YaMvhx9X5c0vl4DgbtrhPd1ZapW4kciFRcDuwx2E+
Igzt3Waa/YKDq7+sReZJbpNiYehCeOgvVa+AH4IMP2uW6o+sCB7OLsYOkYG4/XYJuMO7zTTYZuiR
9QyDmynX95CP4n9/6T5IpyfuaqlHXoFxnPHJ61yyIFWAY2JAkoHUKBOQwGNo6dJ/0zJ4oryXXshV
yyUMKAuYKxoYgpZTge838cFI4j7QadCDAGfLXmuI61b9gKoJZqA+/BIPX2AbTVreP1J5U/tRXMQu
aLUYZem1jDK7rYTT6EEv+Ir9356Svk7gr0Wvq86dW9Hkfh6WXcwiVjkhmTj0+HH69aiYNGpEe6b5
1KY6fpouHfW3P6pJQwwPLXLnsmXzlL/Mz+MhqS1JIYZMEsUWp5SzOkp70l5NACmz+yp7wts6kWdc
LPGtbiqfdJc1m0wR4PyM2Cv+BtbO1c5mChVty3M2Q8PPsm0uy5dpnCIamEHcOCC67aFWd0lzovCK
mlS2onJuHW2u7F2t39z76NGdhM1dXDFT9O8PIRSG0PdPbafplsW+7SlxIUf39rVu6Dt/ZG6WVz0I
KgfSGrFssUkXF9ElIXDGBKSAnarS1F8qNJV6uwseXuQPh/DDhmdszP/Gtuw1ihj/39176SwH5eva
e6ox+r0FTxpLqLpqCdk2Z5JtP+Ys27NSYElry2lXkpzvfnKQXqJWMubDosmUWu+BYVDp0RdQEeRu
6UX0GyJCE8NFmU3eyEUpjAV4pVzsyqbQBnRvfwJxONlrWK4fRgSYa2K7tSE0rlDUYvVcNU2OAZTk
r2XJmbpAZyTGdcUhUas+ANGKWzCcYIvzKult3jP+2G30a7M6RMu6O5P6m/ktu0GrRQ0LGMDMdmAn
O9qFKjpBpNLjGHAdJ2w6v/LWrcgy/ILrLOkUHuq+m8HgAN6iVgteeb5FOgGLQWPCyQxR0et2pMT2
qpcAI6080itEiwnJ8iinXX8HGhv6NZiSWHNrNzGQD5katUysPBNZwa9zyfgBB6Oq5AwlG1CtQVyt
T3C3gI2WSR02K6/dn8k6CaRbGR25ys5l2ca1Bd3IVwJH4z8UFm+SuU0rJprxRYTHMa0xQeSbrAt8
AXzH5aGO3+crh6w0Tey/cxI6Xcr1XDPqF3EUF7S1v5TunLHLnto7ouJ8cbAKt66QKaL7/Lp2IJz/
Yjnci2Si/DqS9ik2+36CV1qukTkrAcB196km2OeZukyiiA1O4flHo2kQ1XNP1vgLCWpINrPCHbEm
13bW0ZY3ZybrbwTtqh+5dSLV0I+fBzwwB5evT7T7Oqio/pOBhfPy2rJ7qIsCn9W218nxZvOtAUFg
Ah1+iJyEnwXyVghRkynkYVdghdSe+Y89KCN42vRTQAiqQmuZhJbnRLtszEcFlChwUjQhguL1UprL
bQ/Xo+YUnxqVx0m4m5njSxpr5NwWYvSEePGBIj0kmBC29JjoQMqYWeFwjeVyQBYS/1EU5IsBI6T3
6BECOrTVVCp0uNw5+6x4wj56KvOaK59hiw1NZNxi4ePRhV2WRlx9V6F7Ly4u67vzEXYXIojnX8Pg
J41jPf7PjsKJ/ZXTsIzyZYJqqFdJ3j7NcnLpewENyfMa++iVV47qN7TZWOUSOJp2MllYCCkFE69z
yUhMD+9LF0CCKuNSnAnp3LQ5VBbhxZZiWS3hoF8Xs1mwd3Blnvcx5NkmNOdkYaIubWOeSPR3Q3o6
jWI+xH2WY7ITFVQvf5v5+Iy5WJKkusvRin3p44B4bBv5qKjndC+WxcDfWEsTimeRQCv7b35peUNm
Wobay7O8UwGE2jzgE2HLcgmvIEY6xdT2mEjMxkA7TonRD3Pn2rLc/ePs+0R9CPRQNW7cTvh1NH5a
z1OlHXpyuWD6RmlzSMQ7pV2/TOIDmEVSwSHXu7aviJqD10g0epji8Qyiyhoq/gussiJTychjS6Hd
ftBOZZbFcS0osbt8fiFliO1K1vOP8KSJcuq1yHWgrUDoAkbaJfgWal8gDt9Tm6Fgyt3F83afzYrs
RTVAxbZvHl2jlny6TjAjBPi0GYEUrBZeFWCrC1KW5/Q6/cKQESFeZTkBvoI+d1xTFO+8CZvMKAj7
YpUOu3MSvG+cS4cYcHqcXIxCEeUDYUfi4DB2hai12cYIv0fpiRac83nbwD6rz0BTSKODY5Kft2rM
c/ScqK7Znmi7S5Ed2iPPvMUq0yAioddRmsIkuRDKT/U5+iRDv9EvUB3eJgzs35VBGZZLwKjITM3u
l2n/G3YjD1kGwfQ1mVAjiwAEUJ5MQ/Zl5plKsa8T5NjKVvlxk50FI2A5dM7CxferCN6dH+gk6YX6
INl6kCYok0DKXXMEkgWRZUMnmPaH2YF8+0foughmnqIyH1l3M5QxzGnFZFhVgsO+gvhn6aAQi6Zg
QIqMPKdofkj69Mp3m8XVCw0YBIsKrebP0YFqlmROlFQ42/Hn0K2axFLJ9EB3T71qAGYkQKbJB6hS
tKHF1ib5WihMcn5uWcCmCffdSjoIv21b4Lrz0f4D+1QaEg9jh6mnxQHdJozZtKIohiZEBHy7zZ5W
yfrY7m1CVacNq8pmjBCnS/UB7+Eg7qxFJk6h9/ZzTa7RL+PP6H5F2RWOZ5FtZGStwxcMiEvsXswh
CDzZWd65FOUula8Zwu9WxRHybWll+n7BueG7ch7ROQJ5z/BKefViKPcc/5E7Z+U0FdFJfK/OrQHz
8cMVaqI2I0nt9H5zdq/NZ44Q4YBNIzfMuTV6LCK9aXEIjNJ2HrTM2P6ognrWMhIJStKYA1kjKWnv
ZiiPPHfiIlSpFZD+h3exenESIlJWGKJxk7C03JcZTfl7gQPpNM3gLlJgNW4udUbJwdoMOWwtKuCW
M9Q4Wd0X+Sj6xJODzVxwloNMTXceoPZkQtVwObRufkuo0/THYpht6P8YHR4iitKHrSbUeFaxRywl
xiK2pMe+6O0cCjWjf68gaM3Gs1sjH/LLfkCnPLcrN/CJfs6MlP3M03DxMfJ5eRJeNp7tZ/PJMi4b
UjyhIjuvzokjboBp8lej6ky+WkczGiXQxJM1IDm+GeRLlzhCDyRMdrZnJlscchdh0UwP05EnTRb7
guOnNweqHr1YnJzvN6J3HLT52dIE0xJJT7uMpTqN4wc2u2cALJybb8DopgbTbCK3IZ3JWYMd3f5o
Nz8rBKBmslxG5kgeYo6aRHYmTRsVQXUU8iZwv4294z0kRH+g5qdOeSen3wpy0fD2RoFHDhZ4q3WQ
5kp3Dsc+CyTWzXytcVkK1XYW7g6YonFipmiAiAkF6e9OCv/p/zdGJgqYGqZho32Av/6Vzt/1czVr
0T1vRy/uOlHe87G0++shpz4FnBZup6iERCeqegb2rBkftSaUS8v4mOI2i1vmXSCk+LYEhAkQGC2T
eXg4rfKEIl97R0QfKe943qjyhC0802QsOXxmZIjAi78T5uM7PjCRlSkZFBLRiU+t29axE1yHaUq8
1bydTuXMihpuOck9KM81VoIxju2agsSuqA/T3AJHuapWeLZsWb9ZBlsQq41WXe88sesxshMQH3rU
26UOWM2opl9OhtD1sJfoTxScdevMdVMtlMVfNI5HAlhzYI3qYbR7OCh/Ni6yHZyZd/71F56zN2iY
lpcLZ2FQowkCBkrLUc0ccv+Gf+sNIhqCMDnABRX0R/R1uJYfEFaRRxVn+0s0A800y3Oq6wwBsgFV
XJ7/Sg9UOWQpGrSs6CkBDuoHLewHRYlzIb0VoT7Zir+VZcQSvkAxfzsgP96R82LlpXuJwq9Uz1Bv
3aG7LFPzLG6y/p2D0vg2OQzCc2Af6+lSknd5hMCO335mXLnIrM4mPv29qyQPbOM/KoR7MhZKkzlF
b6H0OoxF6xhv5QWpXLzCiDopAKWZq5+IiFEPF/dsrbm0hS9kcO9qczgae1vO8BOZoB10wkqmteBp
O03uXVsk8K3nIgjSWvnJVAi4GlrXAU0BQZHtwxuoXwms1e3UTgEPOY0XTROtfVC19TUSAGh6RkU4
fFrHgATFQeYJqRxxQ3rauELdYThw9Gn8nGSITalCobBvZ1oIeuNXwL3Fz5p88W5y87NWJPWDECG1
xqfZdURGIqTv9dC3snOchiw4B9Xh2nW7fcGkuVmD5B3UgKBANLbCGxYqluPnYF+P00iEA8zZLpEd
T/ff4yHywl9+t73Wo7I19fMiwpeGtmq7nJg0fpGVWG1pZ/iPWIdr0jEeV5JrwrjtPtK3HxwcTZv2
cUCHWZCvFRzU45yRjLQyFkFR96ah+wxa5tO+/81ePPyC9t+kj/B/eDKZQYLy0rGd92lxE/erkBRm
n6bus2diMo0IBtYtfCxSS7wCg3PbbOYlLBkqO6aItAGf7+01xBtu4vRL6jazeIrDpv3cPrWgEq2T
xnGBsRZDb/Y8CFPWYxiGrqvvJ8sy6E+miOM5U3Oj+ct51hrn0WMDcs1bF4VSPNZ5TGH0F39hcPou
KcEI/SyfNktu/Bapr82j/pY9t55akK+a8WMmWa8kOV+EEWjKToa3z/4x32YCjxKYNItXKhj5DIYv
y6RfcJgD8vJtQ0JeniFOPwfHHxYDxShsZUK6xOplIieFvb8//Fk3z0Sd8Xhhr1tXbx+n+cTna8dL
pHklcyFF8weuGmM39IrxpL9S8DGldx6D3Ofnt6ECv0EUZsooLi+eQUKl+oH82SAYF35mPVVGVC/Q
e7OmGI/adSOP9RtKEprLahcJwez6VegYBbSsUpeGT33ZGtcSgdgCdODiTSkW+ppOJc3Jxv+mzO60
7z5m/bJE5dMAx1SL2/7uZqrCZZ0aFVDZIT6/V7Cr38JxR9ZDERuOf2oxn6iNRjJXrQUHtW/51qTB
cQ+ypFHnTvLPRUVzz1TH8WVvzofu9HXS8lXKjAt6MxBO4DFOg8iUQfzj3b+/nX6LoJgaOtuv0wi5
Cz1m5JlHo9Q/mXXT+E9I59LkuZNgDQl7ar0X+tXOBV7N547NKlPdaPohwKhOR8BixaYmHPCjLbWR
GJf/tWrPBfdX5tFM0WVp42qHOaSc7butfcBz3mrYI2bN/wXHhmkk8y9VmJQwSbh5HHAPiewaiOLn
nhdm1h0gG8tatbHzunVY0n0S7bezHImnnLHN+X/cuUVcMvgq3xIin+Mt7ES9Ihfxz2aIEJbFbAcy
+eqrRX6ZoTsKyM+9hNLAFiKoNo3eITCjdzN/nS9fH2bfcLdS/x+BKvGfcjtuqAHG2R83iKmQZUlt
LHGfV4pRpavJ355i+bw+EHhx+LBsNAzGWLFdjPLaNLpbM3YIfVrsNRJq7yH+o0Gg26kdYywhzZ1I
lPLQnrkAkdUsGwmG2EPCWMnsqBnQHVdTC53qAQWKf04hzhoUNEkA5pRwuCXCNf6JBObPMzYL2/ro
ApNlCNqeqsYPmdX049edOSvCXNUOF+RgeN0IsMLoLkAQ52vTIN6MiLeRDtZcSfm4XXk+EqBeWCXg
8Sq8JsYGQCr6xf8kQss7cu8bqkpQbEQiQtfHkLD6988C7WhxiZnVFj/hL1cPRCbOdMkChoHu+aqx
1THVGYUMAIJ02THZbbckeIxTjMroI7YIuQz03t7eUYeAP4s4FwRMH0/FxZ5/UZv5Us3fsD45t9zv
4pDkdM20VHCJ+mnlBjM/z4zx+Pm175uPZPfOXy2kETlDLYpUWcZHqH4SXDXOOCusc/X5c/IuDcg/
ltfwMgfEAMpJ+D6gbMKQPWKEtnNIHY0RlSQ2xd1CiwziwDsXVDKm0DyYpqetsa2aqmXkwbc/FEnf
1kmSj2dv7n03/7KhjWa8OVqNiqYmF6FZ01EazV0ynjTIzIPEt+AVGMGLDq+FLYMJOvtTJ3NYw39n
HtSlYgOjKqe5Lh5uS4FT5rYFBp06jgs4EVXFBeGmIXGmp/VCPwcJe2215wxZux63Brik/KtEHDW+
9rptPhB39hdQQlAJCCKaSyKuMwNq/7XCSNSo7agkFm1gSOh7ce5pm4UbiPjRdjfKA2LmvPIonYw1
4lDr/mFuSfsxnl7IxleXZDOwsB6mX5HKgoI2udLl6b3X7kZKknuvCXrdTQ9UryYHWoa8c3tIULv6
iCgaUG2CQ/zFRhuCzIYEKCI4w8+/E9Q32JXGjTDpftbe5ZbXcWBT8VTEdvlI//fX8bPrzDYvDYqg
3W34JTcQlfxUVv39+bLbYjc8SXIjHt84hbgi/7xmiwhrmq2GSDlD+sod1670XyLy/ty/GrPASnw0
byuHRWvnCkZPV7xJqYx5QDrOoHkOnD95ZyppvO6h0QQaU/psZ0B/B7QRK9+x1l9s9RUBrj8v1jwD
nd9uydHmoRCaRAoFfXxvadWVG7vyQau8e2/aDOniAnCthqL2/nVibymCC87pRB+3olUrkmalh0f5
ofzR5yWMqi4//y7L5NhnELBhmQEwkK5vpsAXF6V+kZikPX62pjt7Ls0Pugx4sYuDcay67mDrOyNX
2DfT0OseokPQmWR/0kInLohtY6O8tT68ZGanrH9F6RPCzfkRRpixzVcYjAHzp/HccARazrJ1ew/1
q6Wr3W08EO6ZNOqTZlXjNEHHHOb2DCVko9JY66NPc5O8adnS/AxUahSxSC6rV02vnzmzqu90IZXK
w1jdP1ihlt2gRvO69ZaYT5PEHESfycsPpt7gXAYgj5AlHJm7fApZoMYLylfu7QtoLLKtniDqX+zV
h9ckqF455CnJNBFX1Fg+Km488tDHuH75GK4O2FXA80W2SapP7N1+Ui8M10a//F+aPSCimnoltjF/
SMhBMG3W4qI7Dl5DFiL9JPNpCVOIqQWNEbC3zfTw+e4WUqWNoAjqRxC4K394roJB+IJ/F5p3rEEZ
DRVjJNDjzu07Grh9XyWu9yNJoKEPdg7EoFYxc7i2J2ZArkRyJUpqreZ+2TINPJbP8fiIjH8ZDLyw
x1mmJlW0tUQBgpcqFXVIy9QW5ILKYMHxknzT7liRhmvGhZzQArdL4izj/9kThnZwb0f2BBSYVPzh
hlWFJqf+c1hE5vg7DKJ959WvH81GIC851n+uHFzSgWQO4PICQsye9/pjaHSvBm4hha6X1Ou5Q9qY
Xhyy5pTtusNUgXzzWQSIl+io31ip42GLIRnnR24LiNQbtZQHVTxzVSkQPl/iYsa/wHeKr/APD/cf
9ALAHmDk1DEVQbFTrItY0rBVEitHIYJ0QomrE2kI0OhCjjDeMvxjp7HzTWvyCD9LZvhHVXZpivGC
672bmoBprKI22+ggWDRxXzkp57DfO32m1wnVHJG8bMLTPUHkiJz7CiVy5QVNk/xWGznn3imnH7nm
xAGuDTe4mHzmjMU779QKBPbQMEU7I4qz8qMw1SawwDgy3z8N+7imgxFtxBwa9yuWPbboI8NTU/hb
Ck+Sf8Ii3tDRYvyVktZF3iCxEKgj88vxcksTw5RFvjdZRuTxWLEwVjnFjcZx0eTIZQLs02OLTNBN
wmHBcvyTfzB6vcj1aEkoj4xdu71Vbl3nbJ/WJVUdtXBBl5PZpEVMfo5by1wY8rYgIBa6RPavLLR7
ytV4JIPk9XHuKSRJkgJAuVNSnozeDcnhwp/cpydRkPe0QtK6SQL8Lg+Hhqu+LCQg3VkmCSecl0oX
GTkRzk4s7ETQ3A2FWuFGcWWJzYUYnO0B9JrLenfuXMBIjKKCH6N7+UTt8DUjxd6bYpJsrpReay8a
8SpccLAk90ENubT5HHRJmWPzMRljk9202V9GXlIOSrRQKv6w5OZ0e/+lubJGKS4/GTrovyrBY6lu
ykEE88SdnSZLBL4+/Z46YAuwJoVHi7b3jDJmn0bGUfK0O+Sd4twC18ZoZXuUWNx2XzL0GsweO19f
/zF/le82zLTXBWCKHO5JqQVtYcRAHDLFLfzGuiN15C9eAt9OXmlNVz0vLpxAQcPZ0aorroByWAM8
YboCoy4RMbBK7phvKyt93c7gFO0EqiBjbxHHSwih76NFBfcJdSmIKPKZOtgSuZ25Ea+qntR5SU2b
LG/j/EZcG80mR7Bf01zrLF456udbXczIutJ5GrWW5iUdj6KW0C8Jd1tofeAK7ADYPjkRGlfU0Kqw
eP69FoqE3it2M+ZM5/KfRb+8AD2VmzWFTuRoDompNylaeUHGjkF18R4lu5L02iYELEk072WQWIJl
zq75KJSBkbn8GhmXS3UuS3GequNkBp4dmlrkvII6KvOJYlyy60MYng9oRIXd2DNsBm+RDNLhMPlN
UTPkeEvIRQz4pVLhTIxkP2fk+XMBkDuTg3/MOhelW02SblRpIZkjQ+vyGe7ZHND+q9awWscws1pC
Wi3rsUrP3Gyg13Qsqxzv39EtZ+aFVzA7U86emxz9pQQOJVNRrnzTKrc6rqE28hxFDtqwlWsqWV0U
ZaMKOjcH1aXqjwwoKXoK1yuv5q5Re9+R7ujD/tlpN2NSLMx22NuBeCzgNi5kcRIeEAW+zykNkW6O
XXUFUntOPamLzz7exWGvq9cW1qziAz1pSX/WPBzB6IyWO9zSi2ppLHDsyRU1S+v8rK8UgC4MtNmQ
4xrcE0z6nV5CW33ZWt6LY4EaDqEyLcLs5dUZBr7XHmqX/lAdvj5yBFqfGjmlBUuL/2L0+gLEfS/J
7KMFu6b7Fd8DUqMy8QqdAYE5Hh+m/EveYDeNxEUeExKTt8jPgRipgV7CMxzaoTQwnD6dJ3lFJLHA
O4iy4NPNYppoSnqlxzd5iGbvkJUc/IR7hkHHezi9OmvOuEx+zlynYeckNsQQIqIBdYARNGv+5flm
by9g/XZ0gUQgo4cR0A2laai7e/UgWlJCj0mWAwyzDcEVKJ8ckK+NnuEOgDTNb7UnWIOVGJy/I6qh
banNA1wFmzDZl8VBjT6mzuqspZhBCzJc4N/f0c5Ierdnd0qlKgsrWt3Lqz1wI2JN/h4gRk5QZxnd
wMRdu6mi53Pe1aabZiV6+I8B0Vh8dip9dFP46Yr1ix/cBy+hRcvNQ7kw4BW53iQHDcDIIrhHyz1U
BUc4/GF4Qo1WO9AZoibEKXGf5SvoSDHZ3nPSLkzwxuFkgl6WfmCWIS///TmdBT7LPG88xxQLrNsb
jivqeQzmdCa6e3l/6yQPrEP2Nv/RvcmJ5XKIoylIDjD9GvYj61Gj7Q+KrUdsJYwS+FJ2LomCrPmP
Ypx8wRmnOMsHOPoECAdbnM6TSNk/R6iWzyq5aVChPQufX1UB32X/y72YZVMqAUATmOXw1/lBh//U
a7NuwAjN85Jv8z1sjpz59pop5aK7vk5ayhYyNLBWHfa3Xu6T+mStchPaD4Rj4DL7dCvPk315OvKX
+i/864B0PwjOpwYLtpld83pSEWvM3tRxM6vLxiKjnyNU7ZNhWce1Y3VhbWqkmq6I4XP7Zpy6Sd4/
qUFXxzbcTKtN+ssPenYvxdpxzCDCzMHnyyhGVTabhll72vahY46EhRqX5O0eNRYUF378SVRDZ04r
MwsmFY3Wo99mY7BjvyH/fQ6mJgDWchyXOODCUNLes6Ptu2VHayiZhMCW1bsD8abLqiED7XjfXFex
wQUi/Q3aaYPouD2CMqh2AhXg2NmOpzaKqo/paio5FpfC4DGIV+JI5LzdVzAyMu+xDbQNDne8207s
1fbSzdej1VnWc4dUY/nUh1dRHXhyrvkoT9rzeD/p40oPImlJ4WqM15EScIZTiBCeJs2fs1bxSdnl
KhEHAtkyKvG8Qf26wRXRg2zgJlrQxRsFTAehxq2NZ+K2ZGoDo7sI8RCmrZhhq6c52o7WVgNxFYcs
CqnX0BNMvHTU3VPyYOBeCLwamN9jDSalifh18ySVOBhiW0OGpbiYaJq4kZ+8C8OlmdGwsrNMx0Sf
3R/1UHepftChkrRNCTU7dcxo2sG1znWB8fw30AkCmwomwuvfuJJ9IzWILSRf9/6paPE/PEOQs+zt
Hrr08kGFIs7SGEvAH4u4tCWknZ5q45tGkKzRaLnRCpPGlpMXVpuy4eFlR7CIoMvNLIY2JrI+1ZGp
IumSZxiFWxIO3dpg294LoQVNyeNQMYoBI8lWozbdhvZe1PFWU7KVHSYudsdTQw0vpIT3bWhry7WX
dNXZvZnS5KZ77o4zWwfSZlLFTB3v+sr0OjHf2KL2UOGfWsZlV7enNP3vxObmKU+F/qQMlpE9XktS
+ACiN0PEYs3KX4oWxeSeD8G5aPzd/WnVnYl/jmKvuys5ydXdE+O2SvHckVnz0TrPUNnilvdWUFHW
FaL5hly8MJZphb61seGpPH9pN8HMzXnVOCQPF1KFNrPGcVn7jWBDYepLD2k3UOuHt4mFkFwHRkeQ
HpjpPHo5/VUiXkoWf7Ar9yncV0ehma1a0DSmfhixT/nPW9bTVEUsF711ssoTGxZU7uN/298HGuSO
jXd17TidqQf+U+sfueyjlyK3zeSlMOfs509O2prWLc5RvDD39vyrlqkx+lB36eyGobF4GzEvgCEZ
80LhT23wOe/v+XfvGSGMDnwAPjUQ+ELGCRclfn6yZJEiZj8LHTZ0Xc1K3QlRpYZcj9RQ5zkWy0G9
IksyxzBmJHGxeimf0gMc3CnEedyyAzwp1Z+1z3i+arhLXge14tLPOSMkfbvV2x5TjyomHsEf5oNr
HSSaNc7m53qrwUm+kcgVuPBb1ch6nZKXWQBZgabtEJzZpQRC4p6dqp2F+n0GOyLF3GQ2TZWGjQoE
Ucc81O0klc/Il+s0OVZ0j+PXXrHgH2UXuy/NPEuhMiqknWUwJLUdvZT7ncF5q9gkWXGjweKMnkzn
xIOMrkuVT7IIFYWxReIVGvkXSz8SDhrg/KSBqS1lnm6VQ9voRmBXdlE+A/gEVRuqMp497ParPEZ0
Voi9e4En+KO4z/8JlxhpjAN/MTfUyW7aydIBBnjac/LLiFTBQ1ln3RAUeyEJdQKeBJ6sVpTmjHfE
hFRjnPZZSY3OSHr7JnbKP0XI1oqMtQbMxagZx3owYCn+7VYG2WyXp6D1no2eae8xAZuUYivHQWwG
cNT9I+pSCOXYFhxpE3DYSufxwBF9njN9j6oFfFG1yWsVX4Fj5kJzWQAVJ4m517qQGwMjvP5ZYCdG
dVx7sBsbm7XplGze9UZh0WsqvXOYeezex28vq5Q13cfD4n2QvJo2mrYno89ej3z17Gl7BAPiHUiL
Z4dPpGgs77mCxsfnHwgKvCgexqTdshbOVXyUioMHLbTwJf8GOxHZBuMZkdsh2B6wEIXM3wpuCA6T
bopR0da3biCF9e7/dTJcktsMefLTar0uhPhLgVxCbTmZJOb32dpHdyoIu8zAX4Sy5nbshu7RMFqO
FmhIcZcNFN1kewpYHVZitWmiyw1ey6s4lNFqg9IquJk1zy/8hEGLwDaeUi9C6CPNIG9ysyxZg7G5
PDRgujrWwOZIZTytv5L0CG7Cf0VRX4lnm4iKgBhhXLEZFZJHdmVjs9Sdi6LJ2/ASyKv4LpBST3Vw
xP10emfdkIWnEeD5bGK0OOUFoPmqRvJaDhiW+L70v9g0X5M/p7JwoeIUfkXl+Tj2eQ3o9/dcwdwc
KR5O4RHVLPz1ntEtfmXMoQAB4uYtvloo9zsyqOwRJVlpTLuhZhFiz/5h+PLFoH8813boA7Nv8Wc/
BUt7VpkPY7FFMuFY2qpxaq3M/vcVl6H//FqRg7CttHCUBRP/+RgtgISn/PfuZ0xbNMVmZWwS2thi
+eMY9sQYfXULdW+jhHSmqOqScdKIgtTbhkJSmJbPI9nrahhecQSuu21HrGkO0shT67QbZ2gbLRVB
5pXQntKWBgfvDSKnjmSGh+RJmseuWG11682q/lbWDtEU1OvGCaonmRm2L7FZ+3OktcrU+OysyUm3
uA+EAxBsVXfUAz+ADTNPgqtiQAsU9NEYcYuzOaOyx0/tk1Dr+JJK72B6HEKuvtJNMgQ9D+GAAMXT
LJmkb3ITHacP9LeIhkuC3hynSXwk/3+WKJprAsB+cNwFwR6YMsDaWx0w4jK/fWpYaLCrWf2QQH2W
VELqPA3qlrCHKRP8q3QByoKNSTCX1dzjbpzezfKFG5w5YcyUbBpu8oPa+TI5+t6K8H84OJD6IJQn
CtMZfCo0YgcW8nxHZFnZKfN7lo1HwextB1kEf7k4pX+d/JfiGJYbracwH66fneiKXViaEUUvRsYf
Xry7rbsM0DMES/SHzeuNOOH0yimaQJBnQDmVlfGzFTYnJGyeFYuh92ZDbSdT9S/OjeVQwzGa/h6k
k+f79AZTQUQ+BiDAqOZ+hl+FyyIwo+stuFVQmI9XYBMOQcTSqUj9E/NPbrsz3zKHNOmYskki9e6r
Ei3wqloVOoBZTrGctIdWNl43ElRNaUBhJv7FrVAShFHG/5BwzcJjd7aoOwT3M0+utqBFPfKATbeR
b1P76Uc4dV9K+Aj26Aa4kg3qyZUzcTFvuAgTrSfqSUTgXpuIdB+JE+WaidMJpf2/Sk4Lk3S2DR1L
Uw8tGZncZjYfE2DuHki2Ub17Z9yj2BmD7QqBKDH42NR9pYHZfgEFeG5kUGTnLAZ84Wd39aWLWNwO
bqu5D1cbVjpHTVXncWgpVRBM8rtWUTdNF7XcxlEdj4etDmig85dwL/Zpabr/h0Cd9ep5pJkv7W51
N/EltOwoJKDrWe7sI2ab7Eq1ciBVgz/OvKoizrDRWjT+QdwG1/h6z9KS0RDVlvsvrln0/RQAg0/w
EVYe91mwONRn8ZPkOIYAt64dwYYF3rYJ/d8a9l4d/JqNbyAnBTdKTsXvLEo8iQNOPwcx2hpIlBIE
9JrpXEH0HUs444XsOLy4ro70jwyG71LXn9y2lksYefJ1pm7poHB4SeVi5kYq2q1yeEeMxOIpjqt+
WMcYkWZswaLJEYlk56lF48s0DYw/kTYuVwWvgQei7hURypDUKkWJROAWovA1Qr80ejYPLjZQP99P
f8+OI5QSDn0G8/d9Rhozx7MwsSkSR7rVs10qdzlnmQWEOl6hyL2W4v7cWnSkEJz7SF7UQ5yXGjNx
W0MKBXJteVm74GhvofMsQ4+rxTM3vJObjOFDqs3aJdkN8P4U0VjvBNmi9k9U/GrdHmPCGn71Gg30
A2MtX7O/wHfby0q7KE1OE531uk5APyxck/bEB/11iVrZzMOUrPKX2zpTIo1ZAjCAggYHpm5KsgmJ
whtt20zPNHgEsWcjDymFUqxgALF2XpVpGequCKrpyfawH7XaPJPXzc4dr+myvYiFhSLG3FzITDeE
WbzJKmTsZ3KlVF24pJ/5VPPj7eHGWZarkJyd70qiNx+k2GU1EUaL+p8yk4kOEJM257Pm+JYiPpT2
f+qBVc12uhhWdipnNICk8FWesEjQQcbBpbWyYulpUuYamABP8i7Yp2jwRpKXvaSEsgMO13TVZabm
49dROCK5BrAwowbvIO8pzro/4N4h2Guxtr31ZQzCfR2EhVMfrDbcTRReXzAF+IpOqXIN8oZTix7K
sZ4dwMkUJO11YubEj7juyd9vg9QK/acu81ZUd6rsfm2gm/fBDnJQfdX/2Kx5CyzQ0moQLQIBaLow
cUTe9VPu5nT7TTnGd7R/e0JXU7mHVeYQHP73Jdx2zA2CQnxBr1tOMAl+LRrnFFNOutb0F3r2SxdM
2ZsY+VQuoKPjIn+4sOOOMyAJXglFd+O0IZJWHF1D8l9rKIe21sdE6c/1KN190eYG2k89mAOZIi14
Dy6a4Dseo6aItNSJvkil5tv7AQD43keYzjOQ4FpNvoGrCRmBFB40yB7oFyB0KkyMqfalV3v4nEPg
newxfLwIAgla69wC3jR7slPILnLBbasac9g2wf93Rl9eb/KdZVe8cJcNB884rXBwQAg79sWEF2TK
STiQHT7SbKiMekppKq69tXKF+Kk0riujLWjZeJMRhvt9UnNg30Lmol9ubdlNIOJCLuaoHNiA83vn
nsmEAD9BKCN/u3u8OVJ5ZoIWBuC7PCIq7E6E5GysXjUBZpLlqqVI1v4AME3kOaGHq1Rms47kSLW5
0nAVVytVh44NdeAdcFHsTh/Gs5aqf/fjkTSOXAkkuHj7s+KZ/Y8sAAGU0bsVCYRC7VEfxxNeXflk
Lfqwl232XYk2PPAOXDlEHAeKpAHlXwJr2FVtKJVfjMewl5E2Pv5GpOFBDBK6dKgeh6sxhyAU/FrL
PvdZ4pdFB3dIUkrcwaN4TWcOGlq8rIM6qwztEi2gcCjSDy+rM6V+n3rFrnFLAan8zqxL0F4w+NHf
mdBG8M4/956BcYPPt16o0HAtFMqnUfbG0ROKYDMIqGS86ss+ZJYbbEsIppf4l/9Bv6aCbOJVBU37
vvf9q/8miXpkeYKXLoqbW8RAefH5JAboppKb/BTnB42tlMebX/if9C184KJ029VZmMhNyy/Ai/vp
AFaiXJ2gGLaMcmJdqSDTT4qf9O4v7VaN5TjMvwWhm9BiG5tzL9gCke6koH/VK3B5wcLYCCZVPGDJ
mMxQZx3pXC5qPLmVUxj1lNmf3q7PJJKiGoHQ7udK6lBCv/A26ek3gofZGc79uRVLkxuc/iHZkCOo
jxHdQkAGLdHyUhZ5wImnLeMVK0A/bjFQ3OCI6TW47/0yz5WD2W46OI5ZZSDToaXo7HJQO8+82fmE
GorLUgbPvvH/LpAyL6qnIKS+ctperqp8T7CpQ0i5SwZx8HUy+faoaHx/7Dqbh++mue0P/s/LGW//
5Z8PuXL0R8e8eTHlogyRDIRYhm7G8L5XjlaXJywzkW6o/sQ3sIJ+8ACL8CJc7CKOE9Y9eRR8U6nW
mzdwHUkYmM9J2yD6SsUWR+AHvyUrhTAwunuDne9Ky2kUb4KwvYsYno7ChBZXW0uzVHul936UOCtZ
paK94baexk1D0rsV5yGAnrJyu12cqI3r7DygpcFgW91gUVGdFvZDf53v38Pk2LGOEGYC6m2cspfr
d0vqvFZ2eMWpExpy6+fecatlg+RzM2ff3Zq1HjO7rGVU8bPN4M7ug0fAIHk/Lcvi5dP6i0Ee6z/E
Qt1tsQlmEcbvXmV2stiToTy1JCpaR/5lqdlWp46SAGzKKKWqh6XwlQN0WcBuPfMik9pt71gHs7Sc
DcoriuWlOLkp2bvpW8I6A9gwnwwQE0DjeQl3pPweK7neSrnDb7Y9/ELz2zthREOJZGjSp9p84d/0
O9g+7jEzzC8y1HgDefkubWqzL4F4YPhDF9gN6xfR7vi8ucOsrCtop5uHN70/AsnS1hwgVo0i6Blz
D7D2T8ApC6i+gKljlQGRpunJKGn/Nw4vu0GoHveQ+hdIUm3Rzy+Pze/5iM+TQ7SeIkTakT1+rvEE
2szD9Z1ah5zADi3i+9i9B5qGhtK0x93Oc5/4TT7yfvFJRNOqwRhtvDK9bjXDjlB5Mc3NN4VnwU8j
9DrxSmXvoX1YcxSEEcr3YuzurGqrC0MWSoPPkN24hyvM3JTK2SKrWJkgNQlwNd2UgBhoWhLtJwQD
1WuV5gGqfmbFWhSEwmN44EtomAlPNP7J5fECuecJZj2WGd1u9xRR6jBlcD6Ki8wEtkBhS4CfYQ5Q
bcy+GW2PaqDoXrvWzWlhHSnPIZRVg4UUfdEySp+h4lCKRhDqWGqUL5MOrrWZEL9hGVUb173ruRZ/
dcvdMSRAqt19YlbhuwouDtDbH9U6SX1fmAUOu93ylzpAEK8rpzCQkuXX4aCYEvtWHrQVsOdvVxu/
rvYKeZPfRg3IEC3fN0LZmOTtMDTMMoFpOu6Jy7QQTjABMryTWwXhjgUQF7U3yWFpQiUf6htDlv5V
E5ue2CIlwvTiJ6Fu22/IMu888EejDDZI+IInQUJ35Ed13p79iIA9KGWBcNeO4fU5MAbg0B2eLXaC
SPohbSravvSgq8B+gl1x/7kYK+tsi3o+FoQhbxg87jwafIlFokZ87k5ZwYj5UTPzJNwA+enuZjBn
6ksLo9Qih1Vo2nfoaDoolpaKHwVBZRNey4vqCBGU8ACODl6EFtQTlHqqoE5IsggE0CTd30Tkc8B4
ijYFzw7MJSVPs6EWO68mWycguZMHpEI8VCTb3/ZPR6QVvhukJl1PKrnP7cBZQEKK7L3g41PE3RDU
vRnQ1ppRlLQUoR1vyXGmQl0blZ+xfTEFt9HFpxgp9TlgIYLBKHnsZ9OqbEBsM3OGcigBnc4+qUv1
3nZ2WiyLKV8+OiyyP1DJW6pkYc5GlaTXsyTUv1X4NaELkWApt2bcAU5dmElQBcRONRP1vBGKRlrQ
LtP9w7euKYVdZ1D/L6IHIKyXakrg9W9vC80I7+O1kCNMjxREqwBG55CeZjCjGaQjpQf95IfuTxVo
zD7ggB2Bz3elLvwdVS7E4Tr4gUuRW/bgAWTMeE5OuxImokWuD+JwW5goDKi/yvLgj9T25F7dnZ9n
8ljK31MTto1yIBkRy+T4mKrsKFALfrkKhlWdSpUKZLAVu/YNuDPWDTMR54qOYwaAxA2CdfPOrVkk
svR1EHhspeumBVZGGU69XG4h+Wj0iM/gXLk/18TAVaCp40TFAv53FgmPDZtNUo/TJplxzLVv1n/l
U4BslHfyGB1HjfdhVPhDizBkaG3bCiFJhzG2HDQoqgah959nUrZgJ6UkMFX08romhM+YN7WPJLpP
cJENEHLmWVvHMZsT5DM5SUat7qeu/dO3DizHAWg+6yNsc84O8CY+XNq5AslX7nJSK29c82NqQCSN
0+mNDwr+o7J0EDvxFZOIIe8yKq1JyYxO/eLFxX74WC41EnM9iak09bKvbh3qUZUz7EOh3MC6p64c
z752FI1JrDWWAEr7A/Kxi/wHgPpV1sw321sBdsx3xivsOB3XxRE2QSo/8kUrhvI2zA1UzCipE9wA
6IjCOEB9CViLwws58UC8MqZ5ZgihbMtG71235PWVpR4Z3wpBrAsTVjNyPgiNHPH+JG28nYRVvGzj
WHiSVn0f2Gbzp/zi8Uo1BxZ1nqw4psWlsVfoPkP2VVoHkEXDeHivH/7182K9G6PGoePWfvE0k6lW
DDNQa4Ojabp2ilemF/GTqL9dy9hziQfbIyQM5PMO4ihQPIWW//QJ84u+/eC48YezFK1bn59m5OCk
7wilFJKeF04Fw5jlPagI5PGKzIdLtBD/Eh4u9Do80EdQyJUnE1vaR8Ofm5Nzq6QpLWH+GBQ624hc
QyuikZuRqm7OP8REYOlze58NP9+7x1rgryliVtzHSZCw+Extza9Av3ArmI6xlJ+p4DmMkxnUdv18
DSOF9HM2ncNYwf1mNSNp5t7XEYKWY696UoeOUiersfeeFWbKCFN0XqrxZrYzHLKubaggdyZquoeb
DqQaRVqx1/8cOVanKKm1fFGJh/bW3Xjq3gHeSnzEzKjRNk94BmM74ISEa01NB3oLgjQ9kUMpH970
qP4hq0ynbhTBl0jUQAquS5rhtsLpaC362zMD1mwx5AYUh4j55tWlwTH0/ADw1VkL00oHNueYRyk/
7iV5r0IEkm/4TZXNoV6+mK0aq1l/HxdG66ZZLe4nWGdubCHIEOvrZtuYugIJQ41O2Blh5APd94YZ
Z+6zUEAsGF7NSd8FtZWhr7LLj23glETjpDFgU+Ud5gPd6sve540Wv1FWKEYdC+YWYUoDWBfVxXWE
E1m+zeP4HFs0+KkBMoyO/M/4baY5IY+nAgrQ2uHcJizx/Zdyt4pNmhMAGUvsLTiwdbSjkhc+/e6A
tHME31yB4WANKmh37tU9Lp8/15THNkhpR2hMNCNPCKmDLGjd5H2oXt849XgBcPOCrqypJLLPHpUs
ZPnJ3/qI1+eiTMVlkwcffGw8Qh/MggWx5k/pXBbmGPJuiPX4Adfy1YWrqUBd6h9trrdLu5/Cf1Uc
OAOxrk1aId+veIH99p6TZD3oS1XDC9Rhv0zGK+woIDrmt/Tu0kGHTvfheLVzw7PIuQTkjK0TpSLl
eKLxIGABsaOnG2pcNAhzCEsrxDRRpC4wqgGXE0hV5/B9dEDbIhfOyWuAeNDx2GLh7r3Ja9xCQZ4L
nswCYfYhL6TVgm2kv/XMaxyd0WAUzffmdu+P6cP0lOvg+6damgpRd04rU6dxoh/78nm98gC3hAVY
tm0qpDNR1RVe/571DTq9PtvHrGqY9RbXjl659EevOHynu2BQMZ1kbhj8M+ceKDNEfmvAoGJNz1O0
dV/53hvVBxuZWNIVznhVZFbhV1kagm/QE3FhV1D3RxWL4kFu1vAedH1X/eNcK1WSxNu/ODuDP7Dd
eu9QuDOM66yFgs2Fi/9oqnziq3o2uj1YAMa2OrQoSnAS+Hlo5iIa7sKP3IoppMPVtp0+nlq1ttsn
rWBWn2SDEIL3S64v9sDf8Q9PpLtsGnkGSxIVEFe3zQ9bKnyjfyswyK7nT0/kxwSTCTGhyzQuAn1j
L7tiQ1mEXumFjo41sh/v35TV+FQh6Lj5riUZQAuUrnL+vyQKI2iHt2gAuCgkIkwwxY2bWDx+VTRA
FNSv9xYZQOpZAG866yS+KbU121DStq4LiPCaTfYWMiH/YiM1ZaU8SrVRvP2gqiSnJQspZjhjvLPu
3+HoZLjckBQY8aFkzGoNMfEmQv25Lr41iKuZ90PaXw9hcUYICzCP+HmXUjqGYvaxI6bWagwWToc8
73WyxsrAGjCawHEReOAP+HnFSOZjvKCMnJNgHLC7sXXQVWchV8H4wykTU1XfOFGf0ch9M3zZqW+t
S4lz1pkv9MIK20Yueaiw6iTImyK+li3VW1JfyXg/3xfkTBw45zWE3bcmZL8JI67jhRKeIK9odS0E
nDwNKUh6T0+88l7kW4cCKVlD//+h7WOlrsg7bauIgR8urqleDUjaIsrrwUr0Z4PIR20uxGjsaTn+
VQVAf0JydMlvhbMoC7C+OM2L6SFsveSCWw6kR3VrfD1xBfc84Fg31Zv/B9J5+4B5FgkfzwNTIQNy
/rwOiWApPra31ZWfoMhmFsvSoWjEpYrjFUPEmUM3sP3AdBT43/p9HQnTCHsGxY92AzgXaSpF6+Tv
zZLBuOTsT46RlvId/vRCvghl8L8Zm6ggCzVZv2A1zKk79PWirRY5yD6P7U3KHkd87W78Vp6SKQwG
FDQi759bYqPmfSwo1m1Pb8qeIQU7FKcvIpVv6fEsUKH4ugO8wNCF9eHTXmrb6j9LQebuOZxwNWf7
UlcsXOEmd2NWwH7mEHu1Z5RNPJXDoj84/UD8ta9HM98AAnD7odhKPeDFAeyQH8RfORFhxsQRvlfg
MrNnRTx8/Kmnzaj+eE0t6dNC6EZ2ADcgFCBMKS4l9Z/flYC/AYELUGIzA2wbYIqY14yk1Z1NBkCQ
3MAcr8CId9QZFb8xlmYxjLnNqNXjJXSI53EHRooz5j3teh40YqucdG/HIcmDt/9yX1zOPwmV657o
zuEbsTIuu4X7aoo3acGzKKBYaX3F7rk/21iQo1Z8VuZPqJDtuAz70yD6bClCJdOpFIeFadSGqgXJ
Zv0nVbQSBb0KiBmQQcbp9JOFlHLB+Ufs3Nv8Od4JrBW3ZFXOmCcm7dGsUcDbX/bjJzpsh9UrmIeL
WkZYYNen4m8uHqKWe/aMK2sMe7rTJYb4j8a6/RU36pn+afm9seMVM7eNZrwigCaFvKnxJoogn9ew
HQd8H+sGr8KMr/HhEbCxt1NpdRc+cObEg76ZmRnpgO2/vh0fqXDIQ9qhP0dYn2taQczo84LlFuZq
Aq1gIijV0FyOG61jz6K/HpPFxEYDo4xTGl8bT/NzcX76cegqw/giiVPK4OWDtrf2m92ClA09oLq9
swqCi4uJ41Ow5EgJgcQBjQnABgLOlTa4tt9qWSsvE/LHCxV2xIcE8XzMidH8H0+Xbp+V/qD4HqdC
WRXyzgvyNgup/VUs0eDNzgqR1D1z9CRdm0dj27OBSzBtwZCH9iW83YJV0UBtGSBQkRnBtcemkYo/
wINtoDxJBGVLIRxjq6K1S7xjMgPal6dg/REF3RvyQyp9cqfpUlLJ/HyBsrgI5v97ueilMWlFZKyn
p6nqcsylIIzN458WCsy1rZFb6sNM0bYVt9JdcvOHjNDrB6xrn4ohlUILWjMwsvlV4apMTFJtIAwy
E7Yu+kqK5O5CH6yys8axgDBqXBl753r1zuauH7eX77DH0InpyWFgDSvyp0hBBFkHhnDsNRA33sT2
DN7E3xgeg5zf2KOtHGoOPVkVXGajiUH7QLEa4+ZzSqIb64vW3YanXwbFXCw1hp0lUb5snzOSskG/
EP4O/5zgen+IFFdM7xAJccnjMnHzvg36jmQ/JZgt5dtUy5FrHuVhLAVZB83iZWeAGw2oa9660V2J
6NrdPGD1ykdx0JCnvysTvCqr80vrdvluhXII1LbnmOR6vEW2hXm0c+gArsNGX7Nx+ejGOvYBFAuN
rQQgptYowB8Ge+5W10vwsyTW6hZ+nqvfkDlL4QCCBTtXNB9OHY8bn/6dMAi2DQ/FzvHCU1+IQdnW
SOEVzGg3CnPcrVAW74VgnImBFM0SJTzdi5CYIWI+pF2PO18nFuymFj8Ryc57Ruu7kVqJ7WQohheK
qUffwRWP9vx+lZWGVYTbDhSDhKV0us1dTNGvhUr46+o6XQXRmGgu712b/bb6Cjt4Q6+8BhIGBAjG
D8JarmdvWMy6X7smPAjYHNLL+T6uLhBvjgJbLRWMrAyX7Bt4E/ZZONUmqa6P+r4w7rhV2f8eDvPK
zckBezbcq5n7zW/dLpICEU29TrMHvax7/Wc4Mm2n4yQ+2hn3CRmikRKppoJ2ToAhAMO0qmVM5b+2
9V7tedsVCSaHGxs06G3v5dWYDgbiSxQjLRYEicppHFNccsCmuVzhL6gE3QTrQMzhmnCscRxg/I9I
mDlhTPt4eKUE0iK1BvlTtZdHhT0etyXV9JHB1TBdEw3EUCGrlCtit984/NJIh8D5QHc8ebYi7PDq
foOqa2Y13oRVOupnEBlFqI6q+F3uKj4mL0gUjXXm9AFv+0wUlnvukhKZTUeMHf3AB5oa78RzImkU
JZm+Hnq1pRQnMxUH26acg+6zh4MhIYkU/mb8XFXlaAoBVtDHJ0EpD0lhkWIVG5CQ+4HzrEFyOnyb
HH9RPugUC0gwjW/290dzkWMZCy+nFlqa6VQSTsLSmt0D21zfKfsrXyafpKCfMfMjfoBfrEOTtKuZ
pDg9e1r15/TG7tmn/CKnE0ka4SG+xq21YPEAd5+4UPxRE96A0qKbQLCbmXe+ILHctnbtIUvG5GGa
kKkPHDVh5cEGAikx1KpQlIN25nfPUXG5lIjdywRdi9E8Ppizsb0k7qgO73eYPil5QXEoCwcRAm2/
SPrmzS9Ex+YKRqDs8OD3NrhPfxsyLgb6MHv6IloXNOX61ftiTjNuuIqk7xIDaZvBm4uAkOoaZ8Oy
DoF8d0lG6+TWI5RNzhAZ4eBvfO9gNA3vCQ6P87698ZY8lt2NRz8HOaqISCOfWU9yKppbhWd9zbQy
4i8BVTHKZNB+UmwowRSuihUkNRzeFPRBvKqNW4dzStCfuuG1d3oYJCFanDXp9D0qTeKJ31Z6n9Sm
UElSYnLTSY0GYpVTNz+BKk8hqaqW2zKCM5c60OV/DtaEjCtOkpdotaIXpSGb7f3LdIRwJ7TbSrji
vlzsYWY0FePle3jXp4sFBSP+XLJqKnHG/fzcJn3ag3nUIdfiis/px00Pq5LItfJi8qSLw7uv9PHQ
8q0zOk0B6r+GYcfxTopNMvFd7TSm0bHG7+clzgIkqu6E/O2vreAG2qGPSmj2DSxTTou6Zqm4LfSv
/muk0A930TWfs+ZC3a91fCi9kbA1e0gt2qKeY3bTc8D6+ng2Ejqce+JyVv1+48zr93t9WfdK2hNV
frVqLOKqbtqCjdHaj7+vH/7lCjtDTV40TMvLPd/wiC53Q3sRIODl/m9v5ehwHTdB0hHdeBkvX4YQ
8Ugzbqr96gqdEdu6yNsbX867uHuCeMM7UD9Lq5zv1YZ802QbMAU+OSD5LO+UT3oUOZ+cRiKQnCWH
uXYDeaoQWZ2r0PRLMgl4LZ4riaqD142bFn56ckGGlL3oup+PLivZY+vMmmkq+HDPv2Lsa2j6DkBm
pw67+LRqMWG4FhiRhaRHLF7ZSJxZU4vzaOEkLmZj32k1pvz2H3jtu3bYcBxKUlPWuQTjoRIRC2L6
FQSrBiMsPJf9GCEf2qmsXwey4mcMp6is6bhKabFlUFe3qpaRS9SWfMDdbf5WyE4iihUvTzEERc+9
/sw+TDfTw5Dss0Dh74RVKv2wez8ApkgfcNQE/56nljerj/M0QvUS+vneIIlyPKJ0lv13OctBz6lr
bx2k4Hlj7A/QwnaqVCdUpRZMnb3SW34DNODd6iii42skx0cpmb94ruTc/3XXkmD4gIBYEJUInyNo
ft+eOpDUVIuQAHk9eqXl3ZE8K+vg8N1HLWxVgB9eVABLntm16W/qzSvu5epBK1MGcQKrg8H7Sbn8
Lrtjqgfr6CwHLtZhBr3K3ShH5P+/+axfDHJi+AviPeXe73VqZQIJfwVjQiIbOzDhjLnPLJN266Bj
S2QrTmqbIT5AphZsRUBJPsh8nye4W4722S9bnshXeld9LjTs3vMaOth4y6LKtm6JDUuf15AU6etv
keT1+hEB2DMYZRQ1PZPKkJ6MFjL9hKlnMLCmPg4m3olGUKbpDc9ObdZUH8ko7pjeEIzUZ1ANdQ/a
cuBeqpJclL2lbaWBAqK4VajYdVGypEI1BhSVpeWlGsP9as9UtktnaA9zvGO1Z7yLpENj34UhFJ/e
1/4yGBRiPKXdQW1UQl9VDsu6kERYTYwBMcZbmE39RxWx5mr3aNQDIP/ayfOLPSKxyN01+4jBI4uV
s/wubUEzh3qiGWVCUQJ+sfvl5ShPAvR65AYBwAQixxMj1W9RcW+UeHeA9IAHEppl1FmZpmaAI15y
S8jUWo9B7vUIW0/rBOhyyN72WZ25DjMPoMAxegyHDr6tr9tQsi7oeMGuYPG2kNSshZYWevvVDi0X
/ajDkUHbfaZSgm/v1Ga2m3X4omdqpdar7cJSrcbzR5/78wwvF64g7NHrbf26CdtL6jbnWcZVzK1T
eqW2/WbaA6ygVxqqTgiFnThOGX6fnZ19Z9nG7MHRMwVL3wk2RlDRRv7R/y6q4MuduZCnTKcD73HK
tVdaC16z6GjhUurOtVVrLh8N9a3KTNBA3bJJn0+dkvmOCscoJVn39cFcvczfegJsNXk5wYqqqM/7
Z/LI7Pt9UgUDVZ+C4Xd71zH29Vei9OcfsHDqycSTFCz/l28eURrM7REdW/b5f1v+Awimmke5lT6v
un1RBfnXy4sV6EwSXZAdUcyf4O255JFMm+okhyoQ+ORgC/9GfFJ64KsY73YbFBDyOM41oBP7+blZ
yk04R0Ol0tfP2q08QkWhgAByfEUQ6YZCDURP8D2JAX2J1Y2aVSrgvX9Q45CoIkzuPMPFrK12tRvd
xwjJE1eO0BHrHAvACoCibNgGgfKTZvy7DN79HmmbTspJegO/OivhPpL78Wc1Ic3zx6v7z2eC0+U4
jburoH1PrlDeQ3jKw5ufOGP3NYGbqGoMFbE3YviQeElYCm0WGDvYQ4xovSg3mXOq1LVBk6poDa5O
iAqcOhzbM799jC3AJYAr6W2HunauA4t7kwHaAOe5/uWBtGDmsai0u85EqSuW0qF3GZKAkMn8b39j
vr8q5QZK70fpw5kabCvJExn5YLnZWULCH/2FNAVsRoUOlbNbK80JqX8GP8+VIB/knZjm3ZPODs12
orW4AtJPhFJyoq/meUFe8r1GizzU24K9tiiif2bB22yasYVYbIWI6o8uPMp78hxhUwOb5L2P8WQA
99eKAh67QEbYFS4T7vzGNWQZFLfvnCVFmhHvb1NjqxhYRN92szFqhH9Th69qrZqDAqFgqDXuBeUD
RXLSH0EifYGnDIBHvfdeplKHmjdODEyX+RHzCCw256yLR8Z7chI6m0wbZ5YKpYWQe48GxS8d2dn8
d98TbiYfcpNQsWB3Vz9FblpoZ6k37f5Na/3X01t0NIeact9BeHRUSuojP/1z92LA/cjwRs3+ZMtP
/EE+W6eXMETK7qGFYw9M5XQPdQvo4bMTTiq+B9iMSEWYW2JIhbF2iKB5WLu1oIht+OV2ih9WBGuD
dkI4yDFesxeIwbXpVR7gS67kpTPNHDP0djeNpIfKZPXGR5zkN/OWQyOlYNcbZAL4nQDUy7U0gxYp
UPcVR3FPv1XggzOS9BO2VgQOtwQWlWE8m2BP+9hNSG1ZejDWdZ3TnYrAOAVx6En5G18sU2SAuj/B
F+7vHIwf8zQRVdK3RHk7WB5CDJMhr1rXU6luqJnO6a697r3RSPirJcpLc5VG+ilF59nbtMUlIh45
qjCwsp7jFQq7Sbx6MFSY1acRRoJtG0Gq25XIDafIF/MCiMLd3oK6A48ukU8YTa8Pp961OQHhmfgU
P4ukj4PSRpkx9pdjz6ZTo393BNrMkVLwRP4K9YXZpANs63AdFF405+aLWHv8tuEJPjF7oNcxsKzR
w9cpHMkcOKN09nZhIrEvDgiy9y5IVz98N6XoxAMNXld9RwQZSI329jJuA8ONRJvlvu49Vs/ILnI/
mo4rozzcI6hiJ+rAuOmNpObhq2GsZrwUQtwoQaa4k05Z7tLuzh+J9pANhB2JKhwblEtLHonHGEyx
WjP7DiGjkXSzMi0Gmka2U0u2D4seBp3mzyuz8KKhqc3mZoClNL7XIsFo83M1Zt6iJ4rHtc032IVQ
W6qDlNrPslIR+1fI+GaVd0ooC3SLF9dApdAc/JhwUrU+rKlAwyPO30lRuWW7YXuVqPsXXv31G0j9
5QWHNBWHy9MnAk4q6PL+V+CuoKRwtpKVOCeGHlVEon7d958+NSIy31ZdL7k+vZ66/vUu3DYBv+Yj
PPBo3lJh/ok0iQlkt6gIDE8nrrvHWvd2r2LV7bZxg8jffn9D61ro6Dokp2S4v93YWVEjx/TcfG7E
k5Tk1TtgRQ747/rUoz+VbXV31/3ntwOoyOnIBsDRz/5MGjVJt/UN7kPaxWfMtDeRO6Nrh845wynA
TsydaeSEeZcP52+r1enaMSoCsnhP/5zeDZ5LU9L4/Yh7yKIO470ZHL+YbIgrssu0NvKvOvrknT4y
DF5EYshxCoiAV6ucdyGAcQVz+1vc0haZE5N9pgucYdccRaoijXgR5puxij2n7OpkrYxbn37t8i6U
z3U7y2d09y3C1Dgekn8Vjb2uYmwwT+il83H2olITwo1TIUvNJUZLgpC0hNr1hTOZM+Zew9/EWXTQ
/ECDIsfu9qKUnpnBaDi0an4fbDePLrpo9tkE8PYM9F04dp8CIay1t46zsL4+hJySPMQO/4sPqWp9
R+EXk41kPxSAcwgBTiFRxmWkwKBW54ZRvAQDARlQoz/qFLU4j4U9EngARPafFYqpc/YUNZ445Ohr
5XSoYfb2kbbNaKaoNOUc4DclpNB0/2bSFe2lrsECo7zpaS3PT1nxGRBIoSZTIoBdWLi+AZ/Rgup+
aO/d/FDUu5VmRjgcQXU5jq+5aICecaxzLsvbfGEsZh1RTDBVKAE4rjEkbC7dzqV8ml4LNfnMGkyI
KCkFT0e4bQS02SoUhB5tgeOTtTFnt2iAga129WXWidmIRRRk17enbd7Ejbkbo8N78FYulT45tkcW
XJqtlu0YqxtOLKsfELNjHA4sh+Ln5b18fsQb+JvgYu6+fqwrE0HfcZ9Vx720oUVqdCgTMQEdQOgg
t8pHZiTfQWikjc5fMNmeGduhawHFh/XPDGBgz5mz0dO7TMlCwxbplq+5Vaahc7TMA2YuP74lfz7M
ISR4Yp67jCNQ7SWd2w3j13ElmHfI45qlHYo5hqXx631yZsMTeEkMhFwYHIg8rujsSISmi16Zh66g
op+3wjo4tMrKF+PBxUP0ATIbrIJQAxqxBMQFc0IEjR4S/8UIKtHyv3cF9/zv/WnZHDia7FkaSJ2K
MO8MmTdkGSFR2FBZ88PaPhYu8xHfEc1BWZzGsEs+b9p6D1+lOVUWKS+ngckMPp5AIk2pD1+kdth0
af+nza9chO8DllS29IbGNChwhS799KLoLVYfaiAs830FBRsrlqojmlvA7dw3NxzCqpdY5Q/1le27
RFgZ8ipdR+Cxo05jYINFKnXz9jHnRLD/ArL3EraBXB6CAHzC9IpyhbYCfFQk+dCyIL5yEUYGUop+
vAQNyXdKglu8hJP7s3cBYwWAYgZo35h25DPo6E2p0UMHhAikmLmWehIK5b9yjwBt6mJ29IV7HNGC
A4KafiFulKKzwuALXyql2tHXIkk6jzEHqzli13QgQPfKLL3wPH8OPLzjOt4izUHT08/b4LO9S4ql
mtU2mchzMYoJ4S/2CKxgCy/gB2dEHWJr/R2pZXzR7WwedGmAX6Eei8/ELGG/GwkazOlN4GcBn0rS
ekDrbFi3Q3F/W3LsDWcWTfySaDl+XrvEkK1YohyL0knvttsoJL2L+caJ2xxczUm5XdbYrxI68nSv
E3hCp7U1xgev4hakq97VTxdrroRPcfaROhBRoItdtElVTwS3NqJO8D8XUxoKjixmy1gkDY3m+yp4
Lmu7w5dzFRf6wzdvH37GOp/MGOYofhevwbKF6zzE1NoqJW26R02t9axACdBPW1g8/Zl4oN98a4nU
A7mjtWxMV1lXQy5ZYh9nNFc3rIuIRVdHP+elUnqGZIpnS7LC4/VyaKy4q1KrkbUCFcuB9oqPgqz6
DpLzUP+ADbjT7FImtS9ChatovXv+MCUdvZpAAa8TldHhyxKD14b43QkirgdRBbCiOcgCiewQsftl
ijvoBCyhtyr7S6kK1ZKBh72fmULi1wcZ8Q34n1sbb1pFFmZ+jC5/I1Y/tbvbTzZ93oxJ7tv4N1uu
cCLOY128Pwnjl55bbJIgTg4Vv4Vcy2srCGA/OeInIqqz2ByzkEqbVcdGBr2lIz690O0UlhXmEK+q
LWfbCYiWLdXb446hazMPLt3vdIbfN5EPVgVXSeqAAW/x4durnFVhHWjq5zNsHAu9IS2k3wx4lOow
9LplGUHw5VEg7jXxjXhAwzURUzsRzz5EGrot5gLQI/tELhhUjCN2UOqF/11tyiSbBF97AIP7lmhf
IGIZzkJtvRpa9GnYpa95hfdT86OKjJuGw9f1+PIkQC0Bv0lUCE+uxMsB6xMErM7a1rreEZpjPSL/
dFonrGOrD6VoXpXb3GAtR5OxjdaJC9yueNhAyyXHUkozIHNirqOTGUriWq/wfU6lOuHWQDws9lXk
87P3X98bpvUxV4dYCjkv/K2ulhB+ySTftASHeDS0eqQVd2zJQEqjGBj2GdpJVQLZbiZZcLUjC+wL
k+iR3Rh5UQsPcRrDek1WU9hSbYfyBH1h4VBllv9YtoI/1O/h6MH6s+1uGp6VIHePd4bvTSnFSmL6
ieeu7zlD6jHRIkTbqobgRGGGscV/S+XgFgLG1FpJSMx0lAbmEa/shYqmU+Q4ZQ5cAkofxpOwHJNk
xZqHrG8ihnTzs7aXxWcjiSyu8Ypci2eNmuy++SmLVO2yjx5BwdSJdwp+8qzZZLBWGKMXdl9mAye0
r9Z9r7LLue1+qhJMjrHufu6xg4fPYf8NuPUZPIVP3s7c3hpNauJCwYW10/lstfssTBWBv7JXupW9
ZqQi4Ilff34o9HUNOMEMpaFVqnTlVtLhD+RtTbjyxAf3jEehdvJZ0MLXXcO68lCt+PIAW+OHLzbD
PBlYCmNO87qHzZoA50w6zd4AJZPAvFds9vimHbslCiyTzH6T9MOOIM0gQxmPs5I9YqlD9KuVoNpy
Ses/m7PlQkbXhNgvcUKI2UL9gt7BA+Bfm5DcsvXJt6nX4zyrXHBMNcaoI+zQBItjudOK/nRCUfHT
yJnrg6usvX7oGTSBkrIeHqpCU23QVLd6rVEQ0z3ITncZ8XNpZwEOAxA0fj65WvwnF3MeK55BnXoI
/ZX2pMsTMupdgwtFKjswNfX7TJuH/p6k1opNpCHMQn/DXJyw+vpS+aNwAhySdUuK02OIKNU0S3Tg
gN9bSJW/f1opgjk5tlalBEwv1iIjm0lFC3uRwiVUgkfOkh/iBjIKMTDpnTbMi6FP6c5C3PkQov0N
AmitUeS3PJ1Yjj60YTwim7nPdjjplC5g/JolWjp9fZ5cbEIcTHxyr8kzoEHMtZE2uul/lp56Xd9Z
pnpQNSUTdrfK5Y+4Rjk1r2L/VOHTuq7+TawHxgsop+In8a0n1D58WuQVm2mYFywnCzOO+amK81Nx
V7CTnbk45vJrby+i8YIFlazoQsmM8wn9W98eFu6aNU/m+wU7AHvRd77oy6mhB0jFTyvPUWJa9WEB
9Yg0lk79P5jnp8+dZ+ptZRR0mSqXTkfdfVvlJgcHrzescdqnllES71Kf7ifVxQEaoFJp8hU9tHu9
FpDIPT7eiPbofs+La3m6S3Y6Qp4Awf+ek0Wd31/zAaStzn/6jSrr1LgOrvRHzN4iw76piQEkx+EG
uShuDYyRO2kYxC0ryKpgHJWokgpstgeW0eh9hd022cEpHDkJzwiJiQ4Tuhd8s0OfS+Fm21I71KyG
G6FN2o0mk0CLY4yzmN+tSttZCjscIditGro6RRpcFiQdACTsoyix+1NEJkdQPQsHQN/Ysv5ppkVM
RVv7MBeNmccmcxEX0bTTdfGn8AaJ1uvQV40WWq7DiCBCvj0kz0INVpiPyNdQCHFUm2vX5GsZxCZi
GpNyf/1O3xY+ExK6hAMiawsnYSJxVWisedshFa68QjgWia25iTHVd8Bx84Af7Xrs14kWXriHdhA7
8HGHYwDpkjjBkVeR2nT/x9yjQmgZhzPpO6SryitINaTZWNRWx1z3jpmObVxk+qwvHdn0MsHSFxMH
Opl30kvQgmMvwJi6PKHxBb7UNcCk4IctSTEu/bP9xSnukKq2l4WJYpawjNGi7hZs5hqcE+stZ5Rb
Thh0Vz6XOPfMi10uTC+ydPzmAhqGn2wMIl7X6qwBmBo43MEKiWYUBqJxxZ9fmSfdITreHfop8dQK
WmT6QILpQGAZ5gkAN963L4DpATaluo/qAqvdUz02GbGxjs0HHbE1jMRzhdDgrlD+OcV3lDIKh4vE
X/KjLrNZwAruMC73rJpIs/ar5xeM4nJWZtQG8Wk099ZsjSIhpccnhNx1wXUwrUzhr7XdtPLXG11J
MnjaB8Ys6tc0RU/HO0mGZcOqRpLMn+KGRedb+NgVhPv1mKlAtmXkLamvVnOTb6qbL0yOQmPPIhg8
vDkFWMlDq3y2rPMqlHG0KVtp35ZHvN7ad2LIg1WJn5MghT2InzG8hqznv08z8fmJvNFlEGmNM2w8
cMrqhl2YsajSpOVRXIHmoK6fkelf/kk9Z/4dVi3eixuC6H1XLGZKR89QMLAiYCcP2b5fxJMt+c4b
YqQSHacMg8/ZjCBgnrozvkOR37G9SoP2y2IoeLYwRWF6raHsQ41/XQNfKuUs62t9ZlL4C6s8dHV5
YBIBLpF58i/cOoTYInJoVtl0MVVI78XKtmvrzHRxUJJXDR0iHpQKZKi9oXkwYBSJ1iTVL2SItVRW
Ib988Pc9jffeUKcOBS4sxsunsW0t8cuPNmHcG2K3vUlRNXEnJte/oYYLyNBtK7pisj4vbO+OpYDQ
rQNZJW405E4eEoTI0mqIJ4U2tWdGVyvWiH2sAukso/sQQRYmalyaYDojFRcGPf/nw/WgvXgtRyiX
VkzpKs4YeC9QDWVf9eJNuExFIh85EeFmbWWrCDjLdwPid8orV3aUD77GkJNwfgRK+5Y8yMzNVUDF
2ehpVYjt+6vr/08pP/TJfgY/jcD/CcjsjRG3r7FbuekylUvJuG27WvUE2R4nC4kw3nJ4I+UfH7EE
F2wkEzcwRtRbxfbnwldRDx1p/2GrS6/3wbLvhuZEaK+UL2J+fPTbWQrYwxpQ2Ag5KK+9Nw3jKRUj
mkRTTBHua1BQqCGEvm/LThQ1gaIazFObQ7BR7j9c4n2W+7QX6aflqrOptlfoh+zWgzlOHJ+WSlT0
oB05Y7TQSKxPQQiVjblfaIT05jWQvH/iZvaTRKU/WYz4GsCQNGdhDjiZ9GjNCvHRt5FLJ7OXVQyP
+fsovIxcgtldAZCCF8nb970BGWpR1LmVCooVT4LqWDhl5c22kGra4DBBYCK4lNyD/sXJfKQ2MUwC
tsJWSUY1zVmVDUAiAJ4PotUIWZcuSagHYWtgdchIuncKirTqcoUuZGMN0Pb7tuZbGv1NRfVkEB6R
p4s3GzORs/HRNSo+yNkGCtn3qTzQs3KaLeJcQP2myHxhM1f33pS6Onn37MyIva2fk04F59FDS1Vz
P1EqecyLrWXuIIaHx8af+vAffbGl1arIcB13qNXqzUndGLEiyxHINaOQYiR8cBJE3XMXJxqJ4lBz
awhyQNEmDesnGfJNz17V/+ttTeE7PQKiyink/tm2oAy3JmdxvXQ8I0Cap0FFSsyVrHJc4lAyKoCS
O2nJhS+ez2JamX1iy6pTy09Za14CgXHGDkHg2zEUp2Vw/4KzJNnKkwAOJ2oBfjl0g2El4AwAJDNX
zPGf6k2fzcMW95QXXM75dwp90QExNZ+fCxGQ/tO9s37MI2DnpYUADP86RJ11PWh5PR5JFBxlfRJZ
MhQvKBNcppS/ItvK0/L5tuvZeN8GaIcpGd9MbF2WpNOCk9of49auARc0fWl09XnnYk6fmCPGzwmM
Ur4SmRH+F05JwZjynrM1/AEZhsLaQORzEpcf6auqFqL5Ua2lghZQgsFu3kN7nqTgTddtkOpl29EY
F6WIXwEqQz1rb7evuiJCMzabQTYtVGwXtTjiUqR/mvvKeMN4JY/mKM8PtT1EWNS0jpjzzA2P1yT4
dd3SMnPebQD1YKDA1U1Ayp4ij3Yohm5FxqGj5wJNnoP5PjJbaIsibLHAHelNtnWMf5IaqMGd3PJj
NMDMxn5Fhes/W9PlEIy3P9jq+3nldVIX2m/ZLSSpvzqOUXe/BiCTUQWxLzd2j7y7/WsHGev3DXXT
q/YfLzArKGg1Qzj2FSN9CdKRsUwF6/EA3AHt7idjg70LNI/85jMYWUp9qQpgwKjscGEJ+nrh3vDc
C1d/c+QJ8wSLVb6U+R8ie2khijcZ5vv/6u3jNEWkdcNs1zUGCoVK9qZ2kKCnQhZuBnR8g1oc8gcE
oObEjohe7z5jexOp7OVM32zxKxzMqlG+OVTeljmE/Ths0FUvn2+UkfUOfDe2qyWE1RY667wklFek
JW/9F/1SjzF+gAyHTbl4c+H3/iUHT3k8csBBCpGtnvx9knsxVS7Dx5Sa6ZzuA1j40H/CAOPRTL7e
ykAgHoXSG5cmfs7cVVUVSTqZi1EU+0L8/GGHRho32hQbxbjZxRlvInCNScitmexyi1c4upr3Tfmr
howyzHbDu50JrtaX4LPOUKE1eGPFBlhOpZupA5I+OIKb2DLW0IvN1IT7va07ShSGZu1WHGI5YrpE
tegRZpLMtMzGmMYMg9ZkNcd62Dq1gKlGmxOmYxOYnx9ESZAcHpesV08810lFqqJpPgKp6ihYMA9i
Im7jJBXIUe6x8C6k4q/oOICFqa7q50BEUPLEJAFanvCx7xgzKdMPE51h0Jn0WDZSTthMfXNA9Azq
h1pva1htKqSvEfEGn9E2QeBhiqXATe8czkALBLf3m9Dzm+oCalWDIPZBQTzp9WytMzDn7n7lplI4
HW/trX3XnKvPRGgm2eD38B+Zaokr7U6I5rUBqMBiHO7V27wXYkKyIUFIrlrM5zjXtpo/ewbxZO9q
8QtgZhPLiLkkJC99ax/hWXLz11Fu3XqZ9j3I3QwV7QmpU9O7KO7miSNu9tC7oQejGmdk/CvnU8rM
OddD+45tW2V7kzLjBpGHqa2O91cwGLt00A5spqgIrDo8vg3EyIPbz5nMn+i1tMStqypy+bHBtkzy
SQQJncBRfb9eBfFZrhFY0R684F4qCPZ0XnzdjRkIbkGNNI7U2glxwZaFks8HknMntTwp3S/wZ8bU
ImoBLr0K7YHTYDB1/AUAXw2nWuguthKA3nlg9wq/Dp8pQsHidV4cwYW2su5zYImwVX5BKCxp2KYs
pAjZJGLZgj/55vHgaQ1z4o2jAk4352UM1NnUvcxvIWu8YThPb8H6ncaHsUHWjPFfuQ690ST5R3CI
lcc1w3JbsZocnpM3M3DbxIUVxT69iiT5upL2lCnXiFXCNM1JQKiIddCTjEHHm1xbcdfNtkXSIhci
GFN3HU+dEUSncJn979w9WfK4rX/ugmm1JUHyJHbaQJsMV/uIIgCQWzCDw77ZpBzyeZA0d8iKjuts
A9equoeWFL5jBsDSPA6skOciyt+P6MC6+b6ShoX4wTp9kRpYbRbsFGIhPzyUZmJ5WftXoYZklMtU
hOj8uH8sVwHvrXKJaipLE5UiMAUywAxY3ukLQIo82K0e9lY0mOl1V1ouJe2Vj4YEseANUF9DB7lS
KmeUww+BVy30ATromq7Scn026W4uzHclwExc/6PQj6Tfr7G/Ga2Y4pYAJQTPjRdfL+4p15q2XzTy
24Uq+b/ftcO/hKBbAs4Y44rAy6HtpyNgLjqgRTViKuSOMxd1AC7R74a692LpntZ2BR6oD1LFFbGG
aIou97PNQkcrbSiCbBmFx1/OEi/tjLD9qY+wUTep6GIgpo+RsPBLGvu5MzbdM9P9RR9zjFJuV7hB
LG37w8ckSn8LE9VemXGqGomhhsAFlUgtxfnNZAcMXK1tm+qZ6uHcCaYInzsXSpGocDPfNW5IZkHh
FS5jOWQofgZLYTxwGPyQAK70aeKFTsRgFvjep92FhHDuhNbSg6i+0tiQA6XdSKsxsjYcyMGEGJxh
N7bvsGbTLzTHp9FHSZh7MrUwrKtiyWHghOoU+zvQ6tR8OsV2FKqiRws1t07G8e5SNhrAjbf4JTYB
wVi1NVQkmyN5EO4frDMrkX3iV/bF6wnCuvqsQmMDa7a7GQQQtNzwHcWiKQUFSiMnKLCd1gMdg/qO
LZ4b5U/QOLLSVzATxWiQBHOv4bzJmvFJ+PzU4loo5+AWRcW0LaG+PcQqL7NyYCLgjlRfjPqY97/S
00NEGYUdhQSECQ0g78tvTlKYgP3WGKI1/LoNCvaACuTo0dwuzDUSy4TwOTdSgz6exgnxjttLsc+k
CUZ4kk1bLmJPT9EvpIBOnF6lEVPX5IEvfaEIx7H0GNTKhDVDJLqSXOAw0gAGL3h0p0zQdVmBVlZE
/hyMczy4HvumasUkhsjSGoSuOvwxM9M3WjVCC8hYNpOf43D57QFirrHrwLeYZfkR3h69AjKypK6K
W0zOVcC9/864PKrZuaFPG+FzJhj/2B+Ycg3SrSvdUWIrqFxRjn7vZPtHpzfAGgbc4PtNypSTECkc
hagwMAV4vgOs+vhlLLbpH/fAV7AkeBj0lOlQJa9a8XjSaMTrXl3bhAZoI9AGuHG5iotFFqNHyprH
rhTJQ+Mj8IgbpCeG9g2VUngCPKJ8xLqBWM1Qmx3RGwYIw1cITE/4d43N0xrTcauJ6rCNUEjfHDSo
0TCtK4/4CJUP2iV1pvPMtzLKU6XqbAxOhOLbwtFWaLtfb3JhJs+ItQlT0jCgrQX4+yvowgprhhl9
lUmuN/60/1+Ikiq1dWn7ETOfPlDWj458CZUJSPAey8R4YLmPWqZgjUHu8X6Y3EXcjIv2GSVVn1xc
fRieokASpvt9DOqghZ0rv/4nxPSPfOzjFe32Z0vKSdgainRGRLveA+Iu5PvDXQR51q8i01w28vvq
p0eVX2dih65iKkGGPV4lfpJq6AtRZlXS1sJV8SOCU83ak+toiBWMFjcr+qpRhESLLBnM4B/FvJjl
iv7tMEui0oSG+qP9AFdpGb35uhLapFQlnH4WpJj1TcVRTwt1ecsv/lk421qf1H4n+5gETQuSYO63
FronNDnCwcLkR9CN8yFl2tI7TSzqFYpd3i9VjY0mX2FKBRGRBV/qQY1MRhP4deu5oC0DXPLX9vM6
NpYDgvscNbPcfhuMo1LgL4R47H3Ur1iXzBLbhyZOFufDLamabv4UkkuEHaXWI0UHfGf4Lt+kc1c/
UOMq8jwlUuMEsGyklOFqavOSRYxqNqo2moHlRGQ+iFi1GSxbsVyEudviZL/TG/kKc58C8X8nkSZo
qT2OKhxU+YRSssGzgF+ThqGTj8W4QUyGs8NsHgz6kuC6Af/X3icrKre9wEC/goxteMwwfbJ70VIx
6W0fk4pACNAVE/VzP5yvxFXahOmo/mZi8KABlz39Xq6nZ/w43l3EDTZ9N4bUp+ChlGnxUKVKJGAs
Gp+qScoHtEASO1U9rCrQ79WZ/6AAyLzDHePoUksoDWSMDrMqFdm6X0Q7T3TPZV1myaICT418N7nx
pOmtz9f5luc8U8kjlna/dm+cthPzFrVdmWsGOo7z0QZ5aBJWc4fyVZWzveb2GUqiLtNOU7Y+o7NM
kVC7VHkmJb6acxrBUr6+ngE0rRFyF4UwV+O9Jyr3mLRuxzOBI7Axry0m+JSl1IY0S+nMb4QrtXA9
bTQOWFRdUPDUowf77/1g35f1KKplOWcHM9nUBY4CP5V4bpvQje01X6m0aEfmJJC1ePGpXrNG4OJl
T8GMkZFyiM1U1e0bhiawJCASbX15lQBaMxFMm909nuGJ0soLVWpQSda3L+c7W6t+3VTBqN7fmxyV
1ilpCV6XGhVC5BHNz1tXc/ZXOzXuf+iGnPL1k7Glw3ZllZzjaSApz/HDr5uZxonEyA9NbPcG2Wn4
YonJMa/rCX6J+ZHxTlA0p5URXKkLsUYa7sIrc/VqvV/6uvOfHQ4FMdEWVDKfbRgLmvNNhBYVrr6C
jZPYFKdjee46Z8H0a88EDmyJiVmstR2oNw50WchFUcsqmw2Qux8NeA3JBRxnTLorC0F4lUsju1+l
aY+jSzaG/fUK/uQkCLwLy1RDEYzQZmcK4awhetTI3xp51bGdKDK7I1dWkSO8wSJDxwxeVXMFYpU7
efB5T5QF7ory2eiqkY8vceOrgWdR2AA8popnVDINaQwbBCEniYhAh8FLHls0vIaWx45GAE7DP+X3
icSyJ1s8DRBra7JEhJKZSXdzeC3hnQF+jbI27kafVKuCAYtvtIxND5XbNWIe55UEXKrAPh+QWeF3
763tE+Ktyud8ZBxT0LXWwhpEadXqpQaFSq3qAd6eeM2vGYNqABeB9lHIvLvxIGuQtmlC2Iock9uw
8zJl8NUpB5+5xpl8f/pLTR7MpPejxOVmH7FUIhv1BGKX8IOkNqPktnBCIGu1mVfB6bifMI2HLi8h
uvZHjPKELUunDTPGNTZ3Yde7p1xxB2tFRZ7U2wvy2IqFDnKIOZLDy5WhdfZufSNMK1jp2p80Pyws
30dRsPxJmV3I8ov/TsE0KlFNnHpt0Eu2HURI/rPAj0xsaKaxtRESVlpiA6H0MR+1vN8N2LJ2JWpa
0f3BC/xQNkIX06lrJ7qDlsNOGqhp/Wbs1mIlgiqcFza5l+yKaIyTeLaMH1OzZiidXrwb+OW6d09w
nG623YVihf4Vkl+1WmD1I5CoqXY5p/lL5BjWHiHO6R/+IpHQ8zTYgOs3q903Ke0RidF12Bjp+4pB
k5wria+Mf3B5sLsdbMcjZZctTTCnoH3ZlrnbUeTEuebh2MHQWiyBwhCYjqzp0INYIIKjoVEBdn4D
6vjcsaV+rn6gtTL3pdUSS2sAf5XwYk6WPKRk1qeEZj1vZoQHQvYafhAT+ESHjOCAVycItQAS68A1
m7ifk5Fw0mG9VA3g7g2Do+MG1eqx9UQhrwAxhrBunfPSFTCNttvKXoTY8gE6QmxAGdqo1yRygnKP
vrZKRrAd9SmgExSgk+3NaSSnYdLTYwVLpmd02T4dNIeZn7lQt9iH0KEboIfjlPzeW6A/dmW62rOI
vo2v5Sjyryku08xkc/UhISio/KxEVDf1EB/eObefGdTrHtIlCqYXVZ3l+I6wR975HOX/UOWrFVbV
+pf4ZEadWFeP/1tPHdNr2r2ASucjJ7rSEk40/gvF+jdYx/D3c5s7urdtc67qiECF3TOg/Cg55+H/
WKdl10aFXuB+c0r4ZN1+OpfXjVQdAgnx8qYKL6xe/PcFi1ImukJHJmKeEiXY3Y0p149btFa+NrF5
cnP0A6oTZFu29EQTqemC/YWHOPtcHgFYsKigF1MQM8s+BAAOws8BpnFYZoNwiubF1chj1l0MFaCT
B4ZtGDi6nzedyH5MNg/vA3Lbx4StGfx0tu7ebQf1YPmpqWHOI7Rk2HxVXtO2ukiQG/m9FIrORe4z
Q5p3b/s3/11py2JzFjzvsbBTZ6tRZSYpTlPp8K+NhfSb8JMPDDrkZcTKX/n6yxZbERIpq6wBlNWQ
mU5f/w+knBPTZS57n/JjcS8bds0Q+6lU0NwNMDF2diUOX7tBHbTe7F7xCQrc9EDdHH9HbxVJUSK6
Jxb5zb/63AmJwZ0+WOuMDnwALdga0roDvwgFPq0Wb+Ilb2Np8lmS1+nPAeCspeVnP08uX/DGCVF5
Y/UrS/uS5G9uaxMN5QuiFZUncQ5u88WOPSbAqd8IdeZEx3d8HF5BJyP/Co1DK3USjB9ch3olOnpQ
8C8WbmwfSybFlHCYbusGqT56vZs3wdXaOkf35KN1IDlYZ+rHP4VwTEGmhLOYsWjyRwfB2bc55dUQ
xL0mAteJ7ei60tH3zOFNS0+T2ZA4Uo+QyaHL4PKjnOJSl/wn/KJgXOwELlSSfAPCjJvt1Aq3cne8
BDD3li1njUiK5iJwqOp3hcHC7d4RMMJ5tjD12/O9HL+QavBUzLmnoWQSqFMPoP+dx2PX0AEdNd+W
O4EHfhqs205VigIisMDDZUpxO8kXd6GTqzDS5sHLlcHg/kvF6ROP+WBwnSZ7xaAAsM/YB/APC6/a
Lbi33/djIIJAdxrltG/z/+ZsFcipYJ5UUlXoJ0epH1jC2praoX5NKayeyHXlSVWkTQR8ikbIh1IR
2tqF138vaTitVZhMSmW3JeEAKmgi3T2mCvUW1KZ9W6K0xWdDKsLieWubVGevljVx5xKAACux9oG3
/JCzpN/X7APK/7xninsxzeAt7GA2ZiRz0NLGKH56o4Ha+arK+DqVrgBnvxRuh05x6EpCNEdpmiYu
Rd4xL+hbWnFdm51Hw6FUwLuSSJkb9QdPe8NvqW5s9mAKoKyxn4YtVypYj3Qpkb5Wt2cEVggSqR2a
Gr9z94Ov/kDP0dOy/+6lpm77OFNEWSISYrejHXj+YpEMW8p64mJWgnSkl6N8m5iY66LeyMyL1T7T
FMMF5PSD1UEg6LPUYyopBSZsPRYo/ezRXOvn2bk7TUNxouRmtOJX0vpjHCYR7hjsCGspbr+mH8SU
TAFBU2UzlxI5m+T1C/zMt3yXpXiTVem1iccRJiGzSj1Hmz+PtHd+DdfH2xGg98esWsTtAe5NICfi
TB2XPZcJfxRNvFJPxUQQ9qYyXI1qW/AO8l+qwqFtd2/Sv8AfEmgsTqvx5sP0jCDrxuN0SpCuS8EE
q/UnGfZUNhgYoPmlsTp/641Vok8bPllnMi8Cp5/GE/9h662HS9aJ+be25fuQ44cW6QIyZun0U7b+
B2sN/6Muiqpc91qCPT+gqOUrmx8dLhiOtN2yGq9/gX1s1PC/z63fk2MUpI1dBJ9BYvz4X5i7fXzJ
Z429fCkzaLF46S7RBQSfRZly4vduppiQ51HeMns+VOO0eu2ZexlK8s2TeYk1180LYJk8KN/P2rIF
uBrMmCXvzVa2ieJh9wzdDRSbx+bgVSTx2dcmTQrBMQzD6vlrsIDuAAtsVh6RjItcUmjRz+GsaFf0
S2ehZ+1ZT5NQYZFbOu6XLCgk19X5jYAwUaXLx49gEFl10REH6RSIwUY3woplErKbCERSdCvbu+6b
aqH2JpPLdhsZ/vECHPpMpvqB7kuhRCmENFKKXqouK4+ODWWDoS9ca8sQgvegFYd4kO3iZBchzdxo
qnVZ6Mrz8JmTdu9brw7VTtiQirqeUn6xxAXI5ldcszTu4tMNxcqL401OBMYcW8zGRDS1xc8+CAo7
V4xYLNn3hjd+7WR9QqPILsFj1PimIiiY252ASvJTxLrFFDsB1pnD19BCHboOXT/Nqx7AJY793UV5
xSSbUWkXH2XISnn7DQCY21nawnG6YZjNv7mVazOXuA6/rVPUfzJpSEDgOkkFZVJCA3GO+6cxDeFG
ICDTjFAvijZ1ESwjH5dKTQ77K9qI2jz+m/Ozs2Zif4WnXFOwLnN7d7dSlTikdYEVtgUaLwi4fGii
PwxmRfB3V1zEx2rNvddTV/G//RCV5vr4VlrRgq1b3MaykYmdfp6xRuU2E2ifAPln6s+iYd8FrfDZ
H1X8m44z9irT08JKjE/AjWWpB7cbfX6KI7jWaUCioVNIHB0q02SyITV9uko7iElK6u7AJEiyRito
pTkJoFPXay7D8lQ76KBBQZ9mii7tJ0rst39t2PqO8wUSMDNEypMeQMld15pUX4dlwzZieG0rPFDc
NbTtgnJ/zwl/AgyxnSHzR9PjyJt2/o3CrwyFVJxS5ilH1LtvT8+3xRRHkgoCXz15J7bILArZ/imF
ca5l3MTz6L9h2YDLrFiMFvVXUk/0cq/MmRogcgBTmSsD/ykQ+cPgqA7baxhJrh79e3ZORiI3EqbD
SnLnnTwaH+RQ0CDCgldL/bgAwIULxZMaV3TaehInZuRHx4FUUFtCL3ExJLsdUwlDgK+ip5v6N/wT
lw/ocFgEcTuQp39cU5CsLpiDx2jmRrl3h+kXrF7KTab76ONRFExQ80myBnBbh1Xl5ttoCdD4vakX
JZzT1ZcnYjZpWaLvawEcISepO6CtQjBkBgDUYST52W+ACoqY+zs/b3XcC16dVFiPiLIUWYixpbve
cZV7syFjtN3KDgJ9pmvCnyvAzHVVJA5O8rbCL9ijivqvKfl58S8o+xS3Ehjdqurox/g12KZN3x15
XbT8ipo0y8jm0M3NdaNuzQ501S19ZE4QVxUgKBiQ8qnB0rxhkNJq0bqJo2RRPVwyV2P2PVCw52rR
RCSk5owu+YQxTGj2uokb2ZWo6d8cw7ZXQzah+toreCVK1t3cTUfMQNN9TNcJ9evX2PSROsJySOy0
MYYw1o3ZAvMWZqvq2yZRwj0g2bZ/m3CWUiW5cEM4bA4Hbh8hEutKlYCGx+hLZ1GnFCDJXQiOc0+v
KELp0WOG9mj1GJwCQOqtKiV+biqdwjCpUr7HFcckuU2g2+QC9fndyihjc5Q2ultsOdU9f5SKvYb/
lPI3VvEayAxEH1ppjkDXD2B0w/ombWp1NKI+SdVyPSfOOeIeZzPsycQ/Dq58nyxkXovRFz1Cy4XU
8tcWqkW7nsKtABOUCZrLBfX056TcRQQPMPN6NkglMhbs5VoRnhrIxxrkCmUO65q1ZUacN8HEhHHK
Eh32nPbU9y5OKPXSLuh4mxIOMKF6NS0BcCYR3oat+n8diDY6mnBoEbuQDGUnq5JiieOKh7JtK7ut
6oGw4xPi0NXyiFDH//VcLNBUXzwEBzvV6OtL6S0oeNStrd8DnsVGNM+JvqVbg4e7C353oBlMp2CM
EM8AkUboi9+iy0JBmZumT5rBxpoEOZ4AZkuR8Ns+Cm5hsLzLUaA33cYNOc5BdWD2rTUI/Cjxuv/i
oLxacxtzQXA7MwXLzs6bQm3XSyobf0GzWQDUbwsK2PhQLPkdB6Wqf5EGpdfc0QjX5BkztFbydcAi
Agpazlslcigwm28XZflfxrr7VTUoyW5ckH9PH1YEOLUbP7tX/vxFQfsNv692qq/xWSbT4XnoMGIu
eo4mQYKnj4d3VZcJB2U8v/OWtw+Hq65YOr1x3xmDLilg3kRN6uZkLx96xQ3r95WA1zyRsTPAEGiH
PpJydCCLc8PrI+DP9fWOWxoEThHr5n8NhXAVwiTlx415XVg42F9WzLbICZTVd6eAMx2+teVj84DU
U+GSd1YcNwroxnoFgRdi0c78rnqkGVno9nGdHgIak3mKULggfPbNo1nrUO5+/YL+R2prfyRH4Vv5
NeJa7BZX6TrY+iBfx8yb3u2xXeNIW6dBrMMViq4sa0vtG8tt61J4Lajkwg55rhLw7F5B/J5S+ort
EmLy30fuhS5mVwpoBKcV8XrhCBY7BB9ZpN3dTW78vrSY+2zf6uEXGSzxY7x0iUzyNHN1/l8okQIZ
axo/xULju+JYEypWPNc+TRvyJp8hxJScKevCCs2TqmForEB6Ng9RO10Z/TLT6fe+l3bPz578jTWN
+57ZFpgMygS/r/g2L86ivtFzgHMP4N963JpXtagK9ql3DLm7hkQZg7mbSvC97OZx9Ld33Ds6CW3Z
ZX62FYFZ+XB4NFZFdkadpUm/dQCBGDwm2NJWCN+Pu6dy/pHwgfVuQRmZNtsyvQIWqRlkspiug78O
a488vUQcIq+5B70Q6JDQvfdrkgVvVUcj/ktwpck5BcbPPGXYR3E34qjhCsIIA93/Ou2cgpMzHrFI
VpzdBxzREz/Ypd+ZPnchTvbQg3VRsZnjZdGOxduXF5nFFtsudN3lhw5oDgOnK0YYjmzPN8bR42ID
D2sSV3MYsAKh5Dx3xgHlE0ICfvEopX4NTiEbeEY8sZlaNE2r1Ai4kf6FUqC2FTIzPFXS1RFOcvCd
b6PDAcGU8p/ryjAMeIxfnfSXPc+jAsYTOptkweZvMchbXSaVcrdgB/9Vc3f5Gp39bNCAPW57oRhJ
KQ57ZpCYg9L6pcWo0Rru0onFi9hHdl8fPQFIJarf7sAPTMnw0iozdiu5NINW3IP7tVv9Af4u9xRK
UTSR8vAkUX49JUrSDmSMZ2o+h3Tx3+JOMPqnr8h3WOqZoybd+5hoO/yrqP+PfkG81dcn7HTtffMc
tWDhQkrUyZV01lrSeoh0h9QmW2WO2jxtF3S51+TENCDNcrQ/3RQqm11sclN3HIeiRGeS6X4C6QLs
OqYQN1AU1gsEZKYy7Q8GRi2mjZnJHpvPngo/fvz7gzDwE+gcjf5uV4cevNDe6cZ61De97UIhhB0K
W16uDwGLuZkTcYmuhDaSEyVXohPja4njZf8VyxM1dyasdBbyth6R2d53D4O0/BJY2KCxfb+AscND
NDhMUn9xJJSKjTuWoJ6p/yyf5pvG08TKjR3IfOT0pbgSBXtL3Uuzzj05c1Q2Nr7/3TNY75ZMdZQ/
cYypvFZbNkesYJv3+tH8agAwLi7bNDgNNPhxDF4U0hZUFHhgGaihpk2OHdUlniObqidIU9TQIBsv
gy19RVfrv8n3dEozxsQu4ssmld6kQS77SWWis9RJYb4/+rUqHBGfzPyyklz+SGw6dT2PNRYZHC1S
iwwl88oNsMatgVVbZCd8xB6Kwzbamz9qCtxtm4Jfe0QY2Jiah7rPuswCfteKL0T5TStnXfZcU3L0
NkkQj9cbWevJgB2iuPUE0ZSGH3+gWdXbuYQCQc8Juuj06TWMqnJp4h3Aq8An818R0jna9ToSo4WI
l5gc4HiQcNAm2GOFbdwQ982ghodunqSUfZxqNtbSfdoyb4Uf4m7V+ekBDvjOrc6k+uxknY9PqGvh
URln4d/C/qzn0BWtV6snvw4f3eyWHLMmvuNvw5PG3wPbFfkecJweTPex90anrixj3Zj5XMU2+YvE
pVM2krRzZ8Ce6th4jVMGamw/jnvOTAKJRBBpWqdGizvWR1Yr4m5YhKGZ1fSZHN3G+3VpxTCBhHUx
ZazB9sXL94e/wPxUUQcm2bfqsk+bL1Adg6oQ4469FAuHOrjVNxZZoWBzLBUe+Mef7tLpwP40ewen
snN7rbq+8QgMVElDpfkv5BJIpvOFRnajt/6hX+DQ29pK9ct1LwtgZdPMlRkCNUlNyj6H0BptZ/2e
VdpD7p1Oo+DfFeqUzNp77GehbrPnG1fntDkwIF1RH96/2CC0qLtONP0GsvRAT1wgN709+rYhbAgt
QvLgZmDnZL5Gp7Gxgf/O9onfCymaM3fJcgYaKn/2JO98AQPW15wIUld28DneHyGUZZUnPGCVNQa8
pXewKeMJRCFAMADyXCHURYAGalJz4f30YL4WKULNiZt04imvLKx0K+qBeAj9+3pGC/MEd9QyIEkQ
ZH90MUP+vZu12s7Scl8V2j3wssYLMXF+pJRaK0Tn6DSYaaACfs/DcPAO/QYgoJWMvdfM7tkcKWA7
7UdMJRaTUgWuSAH2Ec5huNjbWXmPF6/sVi5RG0qCJ9u/wCrOlUpP3JrVAoHZUjQSSN1XqgUp0TTg
0QFrMe4/e/GVl7puN4H5qtSfqYlIMjmoplbAEjU551cNc1ZfoJcP55Dbb/PoMOF6HF52xk6eHSnM
XF04vEsr4gM55/N507KOgaKpCdBDFIDSWk43EoPD/ZuiIWYpsmOqLaWRDc/YBUW5fIZpywvqQblM
sKP1cOgIFE1SgFXL/dCvjAGF0IzwrM2pgpwla1kbOXYktqCunmHZrl2MxDoVfYO3FGmgC53WpVOa
ESfvx+Jd+CaNhMPqy95mQ1TTrP70LmGAl4TliV/O5LK4+9jtrTa6zpx1nHOUeE1mtaSrRAsr/HEV
6A8F1mPQqUjyiDVq6xi31AwiZEhAI1J5A6r1jw+oAhlmqivCMODAoPvmHdJDExb5GQKaAWDShfEs
YThK3H5qfXaIjuoIcArbE+dVbqLcuWAkxbah4xV1b01q6ZivRKoZl+QO+3drm93enr+HxjOd/lvc
L2ptogYqfBoKcGmPH9PZNR5QmBcrpXUq3Bp9qkGAkBMa2+ZR1zfAhZSx36mKGwtNVYsKm993V84w
Lub8LCLfloZbGFoh861kFcjOPkpuAytqr0fG/NvcA2M2D8UHSu2mggBex9CTsMiUWVSoW2gIkW3D
2/WYPKbujciUHZQUa6kg87VwiqUFMLUuilKNGE45CLW69lrpaiBdtSfeJKg/GLn2yP5DJcsal28H
46BNMXA2fH+8glGRaMaMZMxccBFl7xdIQnNtpkzopHhFuqy9+BFlP9M5p8ZXYtueeSHYF4A1ZWCH
KS2E5XT5IIG+1qAu9XO3Swz+iG86uUj3sKRWE0sHqO6w4o3OBgSmUuxqxOymLlWdeOAEbY6P+G6N
a/4PMVmUGspXhp9ApnmJ8oxNfujKx+rhsvmtGUypQiF1YD6hvkUyhPqQ32b0xnXj0ZDc01/Zi1Fl
96svtpcT6cjrHi96xpQxP3LjmDqw6I3bLtUHUecJwrRJo+GnB2PN7SuPQ2erdpahMb4zn6WtaWh4
JCk1gYtzxXi22rwfUKV+uFbQ0ucDuU2hLBORxxMTH378lsSlohGtxaNrJDqXcydfC/sNQn610T+w
oFtWCZCXv2dQC5waC/Q0ElOieqpNRxo4vO9MBK5a4/ukkvhHS0hRAft9PYclAagd+nIc/Thmtay2
yBk97osAME/xV7jbOpxiYXeRKk+y/NGVTjZBNcLYjv/iEIna7rgH/iLX+Y/vfjb11Zo2u3qblclK
dBBEd26JqduYtWeqf99jy2ivu8SvsRQahpC2OEJMPnGl9QmuG7JhVHERPBuxeU3T+051kRuxLDLH
G6YRU1w9mBwRoINu/iKlqCzB41KTlWojC1Wr8DsfixOciuSpT03kG3FzvmldYDlzl12qVObg/Jt1
3vWIYpsJOSpRmEuD9M3DUjD3h1hN/qs1VDFNowl/pwLvcZj246YjF3Enon4yoK/BX2kNom++IZtH
/TJKWW5M+KmzZzqS1CrKlAT7cvcBCKjQtBFrB9ylVb04lUkEcNnuSvMm0Enicx1PIyCs5OGxg/TV
Lj1Dqaml9okO9IcpWxNRRpuesIZSspdsZqY+AbosKcBPWqb43mVRxFTu86x3U3NabURDA72pGcpm
L+8cK4dJD/ZEianjielnEGJsR/STzgp8xzpgNnVwlmt8pX/PTa4ljnHvBnw5Wsv7JIFHAVTClR8o
hY5g7ss9ovQOK8DEXRSYT5yL7RO/m1ZnzT9EIFWyqB7JA2MhNr6GoPNtaSpE7y3VHX0/QUOFR3AA
od+k2ZlGQ5hSRKR/JgvtdERYZUAMbeoih8d6ivb4yCuEQQG8mKbJf3sWRhmTSaRTK4rL4m6KN+0p
ULV4b7ebl+SmP8lr3RH4e8SUxINg+iG7gNynqtRCcUeNG8E4jk9/5lNR9JBN427EoOplx/GlhJH8
VyG7n29L/U80+wXHvzwnhy8h21cEaa6trGyNPRRhubu5wfdTNdyDEWLQQzCM4mdmSgNrtI7JBfBC
gLbXsrX+m3Qf/aHuxCN+W6+gQihVihlJHYiFGy/aZlRSs9CE1qbP+NtqSLkwHirHDlS544DEjt97
KwNd5AuC3AwJs3g9MA+OkbEKzAS3xUwavZyqqYg4kVcaB4l8UrOOQW3bBEm58kOXHRLNCOKZOO2C
oR1aczit9ldaozTFL9uUfLgaaWy8yZq6h1AcFbiItE2MDQybTdvs+DhhG22fZMrXwaHaItei8gIZ
03bj5wsZsn3foHLXMDIUjaKa5nHFNNmvjkWQ4fU3sJjBDWpQOZTFdt95t3CIiwL0drBb5zEkz30s
FLmYJkUTizTkKYq35wVEnn+puDCrUrMFIc775LyaVjHo7SPP1V70SPWDZKfCDYyBoFNl3EuQQ80h
JChYT2/T10n0HXbiTrN0nNJrJE1HZ4ZE4heLtrwUYlfjt1SKQQ0l8TGPcePfikEvQmMkQamBXsTv
wzG/9r66T8dqe2FbWR4a+qhiSOQmpc3fH4gmvSL8Kc+fomd+Q6d/OZy86X48ivu46PzbMFiohTWQ
79gBr09mmVRcpNVlF5bDo7gQr/eI2AbP5XYfEo3i92zpK0EwhEtFHkYraIELWYKI8sxRqxjQ/heI
2WtFerbYVIqMy3BKKZmoAw7w7tc8JZR3w8+fsoYcgpoMcrikXP6lTgEGr6y1Ysiyuh0H8Hcwnvor
3EB5chawfpmBQjjfCKiJ0r9FCaVuCPHy8ObKYQiU1n5STS6p9JRUAq+7jmaMCjXdQ5XIT4Batf0u
SkUQlQCdXKNbj7WDk6pcFCW0LSYN83pvNKO1iCtbhPIU29Xsw982oGTdlgpbV+gCay+VJtmYuxnC
4YHeZkLUFdLnbgKPc3zcwZVWxgp4VmXonvHESfIsjkRnbTF4bjONlrfsvdIR48FdC3R9dWMtLtw3
agoL1J8UvlQBmYDc93IYWW7SH2MVQb+aYsQxEjJuR0VFaHHUABass0m1WmUTly1qg+NSnDM9L4P6
0ctE6AImc3+kCRl7MjjOXuQzJ70CLElcUU6ugWIDNqPOtzlParitQUB3RWu0AWgGnRk+d31Nq1Bs
p3mde43ZU6Ia7yhzUtyHpbCxtQRd/91izbwpUAjt8qiRZnKQJqYCN5WxBmlToAS8EkLVYnnCPfVE
TZ80MS2y84MoLIJcAgS19Pd7kuFVV2zpNz+rahWbhh9bqiqUy5E61az6n4905qwvJMTtmPQMpO0G
mOomjGiFUi677BjhA4pWUPdXbHar0Ja+IHjS8YGoNy7ltP6tGouVfiiQqokNaXcunoj4U7Mkr/xc
8q2TzR/qLySbSvO+cdUBsKs65IwrC1UC0lSD8sYbxDh2DhxReIfQIsYyFhCVQR1tcYu5bLH5bhSr
BshdFp25eqKO9c0I0lkbhlKXek/TWVFIyM0z7SqIwOyQIUfoTF2rKwPlsN0CA/Epu6YKTGmK7xXH
FQXVIZUiIuX7pGHStlth4RcpcRYvxNNgVuZIaoU3ytQsO1vIOXGGxL1JbbPhctbvvaUBM3BHDUFM
Sh8ONxlX6uI78fmcpasG6Qp4GOLD3woGLWpaN+A8NgeTFRk9knvGPCd9N+eCnhv2yhBgzjklx6Xe
GmW78XmVC36baZs95GiTeadAckz/L7JaMRHyieotwjVqjFu2IqBjrFKtrWqz9zuhgiOMPF7CkkRK
u1geKC3mWkzYJOa1xQWd+kWm646wyOHX6SoWHNIC/481t3U90cFqsKGEV61VvMTz6XeXm/4WKSM0
u3bRzx0jLoa8XGtdM9zkKHS6AwqzZINEzx3n/mOvysAKbhvuEWv20bo9Ji1wSu8gOhMLirgNKUz3
ByY/cfpc7b6LOZVrB+sT20OOVGjEwn7Nbf0PhOiDuDgYJkZzCXsGKk7Ue/MKfqU+1oZP4ieC16wE
ZtTO7fIu9xn32j1IzZkth1tz7b7vxqEeZebFKXeSfdF8FmrWfnGuew/joD/pUFjsI3A1ZtHdZ/l7
U9F205zEwxeFT4KNfKRlZ3jo/y5wwGeBE/LJq4yY6ryx/zd3jJzU9wRitmKSnIui3ye6JRzqwxWT
8SR4rxDJzHRjXTsGgyqP7u3qMxuppW/gqCQyM1/seb/3I5EPpny3lt6llDnhzNBJJttqWeu8FTZs
DHpP4n/cd6YllZbnY1x5xpt/D09qhMSK3PvV6zgQKcLvW2VxnyM9SwhpgjMrSk3VVFM+sJkc7IFd
PFyXyIMm075i/mDvn1qAU+sHnPb56eFedVtWadnFPKzmlG7+9O2R3PPQsmP21aHTgp1mHmp5fiCa
81T32gi4DlnWRVvoNvUivNc3fa1CZy7ea4TJvnOQDYh2ePDvbyYROaSuQFb2LgzO87eXuxWTOsKL
D/GpKszDCm+NNkaF+C6W/JFJG9okbBdn20j5d92RpuTgA4Pbcoolpw7r+wRDmhAunk7Ra2LRHMxV
6/A378yxbhazxgDyGJNFKHv10d15fMMl18fJSvRJxT/U4nzbwGcrFAy59f5YrRnw1ng5FgNbOccO
QppGtSGpY6UkcEFePB/jXSJLCruurRp3p89qRlFps2OL/hCvANjyy4oU5rpzWR9Clo8GsgbYzAEv
EqGrTicSIwrDdFay21GnPN1TZwEd/47e2BuZ2fMbKePBtvmjmpL3pPhRvJdGhoY3w2Af+TYkDpum
jnkNf+f36IY5CoeQZ4DgA1wmujcLoNBxS69IYuJIFE8CSHcc3O7LVoenLkwlZO5QyLwieM1ktl4k
pQlJScRHzGLG4WGd+1f0vjP6dhA2MWtS/Rr/ONlyuVl8AmrEDGuKViKqn1kChUfo/4py1YkmSeOq
rUYakd7l4tfn0bSCg7r7wZ+6j87Lbm3EK+M/9Uha+qaGDQtBjynOy7ykmyFiD2J2fnOAcuB2gkVo
FI6rgWETcyyMvqNjooAQe9gs2yEI3E8/o6XTDX66qTHIhvbi1sW3x7g4Ng75B4+AyPOJVL9QSdiU
cUD9oMR7Lo6GRbwicfAJTrGuCSXcOEDKs0ZmpjK7re38/1Lv0TzrU/xH428q/5WBhPQoEqx3Rqmm
HgkphRYyGI+KiNmUfpTRoZrFIFK1nnlIJZLp71x/IvxPKMhFHTQYFcjTUCFuKRyyVFU+EAkgMQgO
ItLdHUf8zudMRSgmqlYiz4aNdym0JuG2S8KRUnn6zU4A7gj4gwQN61Br23aToYKj2fkDajfRNDt/
ML8YqMkP8+a/yiFbG9RKOOceuGMJHYzPwyyerD52EcgDubsybQK5vFdPFTA31n3uC26xZPxzqh+t
SAP7WrJQO+3LN5bVIFng01+biiz+H2BLNiBHm0/9fT+VsKkZRjyL4HX58RpTIR/Uwuk94+S2NOfg
nBbFNArfYuEB2zZI5kGAnaD1Ox+z7OV+faRUeZIBAcPUCtZer0kHoBF7PzzsApswzRq/Tx8iU4bB
ZJ+5r1xJuvicN6nDLsQdo06CbeZMrKZSOehxV7DWaVbQ71IwfXRO7NmHNgj65dvY0rSgUMIOShXt
YWyT9g2U/Sm76nOVWHPMPUPTu4CNcDwRu9UudvyoVJv5uctxFtlSm4CG9Y+d3kjFdvZg9rAsYgbd
YURbyH77kAsKof2RxNtTYPXetxGejdqcw57JY+lZZMxzHey+qM2Nx8ojpAycTBuaw72EC45ib3iF
y1zPyISliPYPP3rxQh0Oli8T6MHpDphV+4uGTdskN/4Xk8TDifTcR2Mv0WDLHG35diBCp9ir2xyH
DzOI1aQeDqTj64muFYFKUm0tKEn5DvGU9ZrrfZxAbFQoB28+bmkTiGaYidj5Q2IyvwHiWJCldFT1
1xWqs5sCvNdgaGy9n2ynNtWPvR93hJ1kiidiZA3bBmSQ5ASrHCSoZK+Se98gcj3qJV6VGxJGHaeE
g5LXQ3TDzTIicziVmrf7hw+0ytE2wI0ZpfujyPGwFAVMFR+S9LUiQ3VLtGMRKQKN0RZMJyGk/A94
+3/eecVuzA+Jy7+9u7b6y8JVNnMF/b83Jgwcvq/B0tdozlh5rDp7EmDk2luUxEoUP9lkSveEVf2I
XpJWEP90RJSi1CSg1aiP/FFcL8yH8tDzwbn4zlMLNQG8NPTq8mcGiKaigafpsjY0pblwye/ng+6b
QqA45J31FDKkvUzS3IYEHWEItloFWocr4IR5Q2KAJGADYVk5WObGBIdagrBPx43/nSl0Mtxyynb3
a/SEaeHEQG3483u+FnJ9RO4u0ynqIlEnljM4qxAX4R8EEMEVvMZXhSJku30w1EPT2n5Ua3jF+9H0
l1pWQL4mBjBhZUv8clHPhMpfKeO2PuiyOfiiZDnGI70WVnODl+tL7Ch+rZTe72Pfqzvoe1v174h6
6pcvyHtRjlI18hOCMAZ3f2SB3bOSBAs34u1BwC+e2iNoTjyxNRTzION3359ynQr9nqEsccDvjKIy
FC+9i8wqv2PxnGS4wMPl3sBZ4t6xDhfAe5RIZ/Hs/U+f25KCozX5ZgciEcLCPVbnbGrr0VO5YAU9
y/dp1Smr1QxqQwp+PuUQVLEX3ZNxvJaIyDPsWQQU8X2Fva6xOnQa0J+mt6A/vXxOls9nNE+17CBz
oIK1jlxegn7wN6AazVPDBRwq9C3HDKqEsdZKjchuVylcBvx5M1/DjqbB+JXFIvWGOIfVY6vJMuuC
ih9Hw3MGI01gJjJl8iVH5XyLbpPkmgmdSa4lkx3HsMPbc/SSG7ajFNPiHiiWF3cIaPDU4Fu6DOcS
aOd3Jv87p5vTdFLRWFfP3wbMuCuVCh2mKdI0IH24Tz/0Ox8f7OL+lYO0ysvymoxC4o9Sy4VcX3PC
Lvv4PsA5lOfTn3ZE6Vz7i0FLrYUa4xtOcHNhJn2FIK5E1uIO//Eqli5tJuYWzbsh2xCYTZfPP/UC
+50PEEpf880wmvt/Yv7QVfMvfv1wVyO54Jm3tSW2903qPkfK4iWG0R/J/yn8aqwcQu8kaxaopvaZ
4JhYVhSNmC8XwOwKNjfJ4Ke7BszMwGqEQsl3bx6jfPjCP4uV2gi5NO0mhVmZsCIu8vYXd2S23j6t
QoauyYYBov4UrtWdMm0Jjo6uiCm8dFHYEkIdCcaadZbEAWGN08u8K0V6zBA+56oOzg2JPpIENfmM
KGDDnE2mKD4vzYghZX5JwGvcLE75kaFoPe4kyKfFMVTD9PxXWfEFV0Tvw3XZtPOB/mbAciwPwGlS
4fySlazI09eWppHhHvdCnlR2ePPiuKqP0MxDgPxMUb3EgJyj8MqSFfibP6gJauYTO5gVL5UdbBiL
6P0kWcrjD30njIGTVHu6Q8YeCwCZVInZwzPiccglGWmHs7/iCkVg5vDD4ULRIHLb2fljQRA1u7lv
neuhBlYi15SBTdtS2XwspoNXmefMde5efYsHINZ4g9aatrN0aHDb2A0VxrGCs8gL12Q/sKDRn7dg
WT1K5SFU+WAL1b9zhU6zEooEO4lv4qjYwh0B8K6l9fDxU0os3wTHk1peKnagcaDNRo1gr1u04ArV
WmU51LWD5dkEOSHl4wGwkKB1JzlPGuc4ZhHm/OXySeN++EBHhK0ssGWaZRW9JJHMVG7md30cH9oi
SHNxx8xNFPhtLwDN/Fl3677s8XI21ghk3nkAac1xBCTFLGDJc1Alh1L6GhxjhZxAOah4wLH2yae5
1gPfd9T9TMwJa2S6ccQ707Qlu53rJrNaX8JASG7lNBtoAIserK8BSisMz02onBNge/NB9b64PvII
GRX3hsQvp/ZyjqwB7j47v3Pj1DP03WldzK9gyLljIaraMonhIZE4R+DRVkYood3qrHucH4I6MgAu
fr0++UF/tRUe8kt1b72axJEt650AVp7uizDVY9q60rQuv45LWsfgE38NUd8O+Vo9J9kUZJabNJIE
ZiJQ0pEJU/rY3ozgoJ9Wefg3OB0/ZcLvsNh87+zbB2RX9KDT7FPoaByFSad6DEHsk+yD9ysnQ/L2
rzKJhJWOq3WgAWP2dXNrVY6Dd6z96GErUyKoLSdV4r0Ns80HDpmdpoEkcb6Bd8HfgOw50RwRuwIi
imZMHoa3laS7OUDDCCELufad6/OoSM0m0bpWAT3+YML2aed9vXryscRpT5iw7lM3yUaKgeghDAbW
gHsabJEsRQpV/tTlPYjyA1/uuL8Gvlsd3xVe/7ksQawwAu4gv5vgFAGLfN/vtttomPhyebhBkd/b
uLCGM8/m3xrKPMk/19qeNKdmBeIzhVW0rnQu474QaHllpJP+2z//Y4CJMXqxs5rJtEW1nG4i1C4u
gm8TeFjiz8M34gTbTRbLJC6Nn6pA7zU++44H8RSifq2q8wup0otjt8wtPfht7ZPSrccbJMtBYcXy
DfS+vTJqDFArDGyRaF10TMJKqivVrk7pTHGGfp7Mb/CDo/tSff9SBVTavdS2EFEf5r+KR+Xft2XY
64WW0tsDG1n57MJt8IZCmcnk1IvDoFt7V3SfetbmkYUhYF64YV5DlcvkUoL2nDt+TvA5gUoT74dI
qRHctqVg3HIYuY2/Aphq3+5Fd1PPSldYJa/jNcX5YtMRrNBvMbgttpjhZlmU4+dKnr/QLAydKXjX
SbX9Q9ALpYKNQx0LWVdaYwZCvQBtaMH6KBqovShchlp2yG7jO5YXXMjb5jdwYQN9H2EvuR5jJk03
sJgqK+LxxETZGrUGZ90paRBiO9tdwwmKK07JMalFQtvXUgM8bkDTfPcotI7UcI0Dd57QWGWo/v7g
flt4G3TtbFTmIHjfGwMb7VHjY8uu5E/MLLPEUd7H4KGBR+kOPU6/RtT3poKxV7Id7If+6JRFQHya
21poIWECgRhK4Z69hMap9zUITo+wiP/VKAwaZBhd9MsXnOnwiGTRqd1HOKg5z+w5li4DXK2tUFsf
T/6HfBngy1cB35BCngC0XkzTxv0ABCCmCDOhncukUYkTKwErL12zRgyU4ISfTvgH/ojV357ni2c7
Mv4I+z3/ciO9IomyaxtQ/Sj1dZEuD5trG1OJT2qTJrb8xVMwqtRjOtIMBDztWlcHPMhZPfQKIQuS
uEu5jyXNSMg9DbPF+6DY/KtAADQIASxiHzaCAkRruLu61R3CHj4qE3CoC+Oo18Mak5ZkfCpW5YWh
G1ZBoiEz+fVbV/wofuevxLBbTQ20FsmXGjJBKKdDZCCI9xLyOsA1UsTIaMYF4sk4zMiNXg1PV8n9
rKPC6qbYny3Ayrx8hBmIMnLuLGcvUfvw3GY/W5F76FI5CVoozz1wC1yl0lc+BzyiwWDYVTrSiQin
lMWA/1p17tt+ib8C2yO6jBFXSmvLJWkZd687GxB94TufCj4aDE5tOES2f6qtKr23zc+PnXKJgZGl
owda0aUCB3VpwfqkCWHJ5VEIgs8m+HbQrpLvIymRAUriLXyl3PK7snMVveLU3dLg8yM0LU2XIzko
HOa1nl5HYVciV6r4U5paRc6n7SdpMdzsfj5IKp/DGNjfD2L+QqkjLemJwvofyhFGXyX5Hp0972b7
tcdtP7f1A7gkPEajfGIPVxmGsmBNlWnAuGWpakCgBKUBO4ImSQlGSNMmDYmJnesnnLjY2+xyeXdh
ZBH9M+l/GY2VqzROaGnGFdSKtnPSojzPK5/XGXAoNJqIDtGXnXiEibCyWSSmATjhdC7E63DGEh7Y
vjpKa+YEXdxQGW6VJJzSPgVOlWNK4e9kERGO6d22qq3M0lJTa3XpaVgmn5aziICCY0V0ruFOoi6B
2gRvXw1ugM4YiA+52ETgdM1jywPkV0z4cpTUStYOXa5o4idwOs7a2pADyqfBzUy0G0dLMwKflTYl
GyA0luz35CegwkpDtnRlYqbl2484/AsCxEAHCXCwxKjiIupfxc7consJfOdeb71Jz6hO+D0Efm6S
lbD30Eg9xfP/iNUbYr+vnGvgV5AzSmXcyxxKj8AOFTxYq9uraM6ZWMJtLhM7mGR3j4CGlIlmRzOZ
vrhmlaNcH3paEGb4tTOuNDvzJrafXwAdHiJw+vxlZt1RZ1jS375oZhWOdIHIC7/tA9uV48Dz1P6C
+bTLp/WqiqsNU2jkpfe0y+LgP+Nnc4m3BrXUZUqfiOm4ekq/YaKNXWNUmK0G+ME4pWHZWfMSbK/o
HP2I+vxpzVlC+RWjY8W1kTOQuGJWYM2N6laV+2QemdXs9EsPoF691KMkJ0ELqMVwiuwGuBwYS58h
7N76HvvQ8bQqUr4Nm9YKicKf61mI4HHC+2J/yKQ3rLhL8nZjV426sjFH1Vs5ISC6Gic8KhE+08rS
a16/8qOBGNZ19QcOAmBB/6gqHwT3tagyMPxvO6FmyL4i/oFkAAS5QrtB9K61/K+l+rGANnJfjDGM
76yCD9HqqOlGnRPa4/dRCa49rpxWFlEhbVeAaP4tVvEPqcCw7Ewld2TAcTYUEvFF8qLo1jsNdtj/
c5fZJzzybK/vmUXpiaXJ4tr7ow7+hxFMORGunHnr4IMgx2jg2IZDNzYcz+p4fseBBpLZnoOroem7
BA3djaYqao5g9uxBLhK3TMBdtBWC3ncPaC+NrhV2bUUU/KGfIqXt5PNxxArfy8iKQQJLzv3ZWZnB
wuAvJ7Nl8s+L5ymNRFnBcHWhMOUhsS3tLMba4wU2kRjjEQYRXPl/+OCgDB/IZJxegV04hwdM1qZ2
kUfzm62FBYXLscwRe+Lzi9hVAwjzH5mPBN+HqYMN7o786jeJGGmX88Avwl6jO2QK09mFjdlS0S0p
j4M+ANc9yRF/O6WFgNYbUe78ATYOCnsGSXkn9mWjhyabG5S0UDkc/PDPbXOwrzYZaLSNd1GJ8514
avxkSKvhdU3c9NI5hGfI7BcnNKrjpwl1gCsj5Lz1OAc3IRxLPDFbIqbcbVtS9beUCpet+i9LnLFY
jIm0RzxVJ3CLjFpUHLUFrcwu9jxt7kpPunsbY7uy6PH5RdYaW/tZB8rdHcC/x+DWZNaiHXQPZU33
WTTUFOx7qD0wh7DIZEmjRHrb7dYB11V0T8pjHgmCEjVn7BcODg4ijtoOaqusT9WO6Z/SUEgF0Ugk
89Rk+WOjw1Vn6Zo4Wkyem2bFmJWnKGs7TgEAXTTmdFD24/gz1H7c/8Og6VZk39D9PLOSN7JwOTFN
qnP5NUWtTxcz5PczgOP2T42Y9Dy8ohAmZTCp8kZHBpdqHmJAVa4/lZeOolzZUTt6yxWsgEQ01t71
z57goIhfqeooBEA5BRb8/ZUAAxp8csSpGBPcvCM5ed8hrsLZVFyTMUF+eUDYM4DJRi4Kya90KYmI
a7YEwy8DKlrea/AXTiMJtyDQQPPv17/guWyOOGlZcFW3VeWZcnjIDPcaJhuwYrtD0rFy+5wrAkBg
RtIKaRU535InII+cPeSOObU8ibv3pgXwCkC1vN6m2nn0+0D3qYRBE+70u2JzQ+CpURefqBtqOZl4
yolK6qbXSkO6olJ9T+6IFT9H8VwTUdrZh1qov5r4H5Vn+Zz7zbcqmmDIdtvHFMIatXOxB1Nna5Wv
lTJGpqf0E7QyF0J6QcN97K5VtyM1JDU1I9gUoiAyUvbTH/XErwt+5fclNyOw8yonbh/wOKBKvpsn
tXFylmtjMI83iz/UBpbA8PAGxSkzblPjkq0pm8XJbYtQMNgsHWVE6gQQlQE3Gtpp4FV2DP8B7GMi
o8sGw/YkgZ7mnGvMtZNy6n6fbCWOibD+lB2zuD5d0kqsMI+4kBFmUAgMLFIDyxohezQkUj+xMAbk
7zazAE2LiIyYtMT936DG3zoyN6o64Mhhtdit7dTFRTLsfBVODeBlZSxi9KfF9L4qFlQRIztgjGM+
nh3uH66B8R4OR8HLwvHimC+N7KwcQ5AhJDLDudeha2Po1ooGSI9z7ZHFdnIfA5ec+dQGZzHeAD0E
Tv9SK5Hee837sBDAojh3AEIXpSN6jHj6AkCBBy8tyoxcA+bG70upLPkPZZOwGVou9qDlfp/1DLZY
G1jSKjWNEvwmwSWYjIqJvJHilfYuAmPwm+QIMLxet1heJRlE0r9W7rUCHHBvVbUAKAHz4vqJSAcV
gvXXelGqj3w0mu5cgHrqvuBU3BTNNoG5n094ZFy+anj8ExcnVr9ejqGSimuBOEKuIYtcVLOCQEtE
w3Hg4tr4Ar3MEFL0ud/JtWz16p/DtopkR87n+BsKmRxdRx5uas0yd4+ECiCAdfz5nNVg704SoI9L
y/VrBrbanYG7yjkjsvtxmvFndfeJm6cefrlLa3lm0uSLLojVDQ2XI6uzmFKMeclO00B9D6rcA8Ql
wafiZek5pDu4/yWCwBnW30PxTRyj8g4k0/I3xLZ4jLJsFXyoGZQWZSgLNpH921v9NvD0+teNiCaB
/6o9Mz+1cD79LniGjqZP+ywoFBqIH2+QDTfLYG0TpEg4j5H0sAxoJcNZKRxdZJkqOrGas01cOqdP
20nBE7vrg2lHFKZwOv2ALZLSTJPcmE4kwEVaVpVxSfhlotrFnJkMn5E6UARX7bOx/YM0z8ZdUzE8
9T+VQUXYDImEpd+y3TexioUdZAlzWhE3CdgJgYz42yHhJdxiCnFBUEUHNP9H32b//OgK7dCowZ6v
SnHLx7NTjd/UCIW7dA4dmm6YoSVfDiXlE5mHSoHdANgBE9RCA7tOqGbfB5p44YkkcX7PRtPQKt4Q
v4dFZXeb+HUajmVY3iiESV8f4OjekwixctwPlOLsF5yEwpiDgyoidr6DVAzePUKKEOtn1PKaJoLL
TES5RkFEnhOk63TJQOjSSsMc2Hfna0r+qw6KzMbpSYHFvkGqvnxHCNSsOWm/TZQYnoRh3BkGs/vd
lvgRB/KOJ8/M2S4EtsBb4I5eBIwMd2xT1edEgoX4CkrsjbiD4EyaiIKa1EGBAHT1PIZCBVDxarVf
b2EWKGXkOKLnxYkXeKi31qxLFlRoL/ctWnyAtGRjqv+HnvDGivcV4vSk+Pcou8UWwlUbE6fCMTfM
E45RDyDWeCueiegamrhlLZeefXs9+r9Gy73gXnb8Jl9VLtSUiem5u/T4xZ7+C94nxFhq2R0Gfwz4
4YsitrmMheOlM/+brxAOJAm1zuoRiSB98QANvAVc2h0GwPq15AfPL6ecYKdbCnwBdV7OoDsx+dYr
2EB9v/xtEtHHr7o8wNI/LAlaJhyjEtW1q/okdKGzcCbTwYGJ34kuAFhuz251MqMuhcuQ7Lj5/0bc
sgSfO3KlCrmG0Jbg4VNqXWhmSCgblzvFO6x4mLPNehSEURWNzkq5fxLWovWl2efT9RS5McZeWaiC
ON1W1j/5XTHEWQpD5ttVeSu80BScwRAH6P7Kb3OpwZk7WH8H7OG7ksS12R8meH0tJ90ZQeFJ034+
ly8PZo2TEdEk7G+7FUqbeBf6x6JfsNGJEPV480d4m0DTDn1z/dn+Mr60kBHGg91XeCBCFinK3eOH
h1E3I4Hw3FU+/P6Y9b78chpXy++gyCuPzWCWNwgqZ7hY+yt87x0C9XVdDHIt/1rAs1FJSbuwTbC9
fpZ6EbCE2Y+ObW5VSHu95z9Gr4vCy62/9nrlclwzF5tVmBKPJFV/GDhapigy6uClWjXWFnq5cT+y
UzilDVSRFJA4FkIWdpwajQ/IQs50CgwttcumfSnhr2h9lyrhrFMHj9F2aPBBu6b+GtRgyLy5w8qH
lsphZUWCNUIHMsEvECkVsmUDgzUA9pFkHvZteol0ix3FPl9ZAex4V/IsxKgzEnSuaV5GPSdLKUm0
F2ay2qMWNXvilEUWyAIAzgO0x3UCrAauV+KpfVsmfytDCHCYmVr3WhZS/xaT7QzYQXmR7YHZKQAg
ioX3N9Bpc5y4MOat77hEicahMgGH2OQpt9P5imrR3r1wj2wzcLLcXAUygWDgnyVsBqLFuCPVJIJt
axu1aCfKbO4Kt94sVt06CLb2SQti+2gXgCJHDVLpJcTbC1zChGCmCeRxRRfuNTjqsa1yhH7cPvrI
OptLXMIMYgUYa8haEtMdsOnfnyyDVvH0VMiLqYaZm5bFPVEISiD9EE3TpRGLKhfkW/kQuJOjd8Z3
8qpezCyDqxO9x/wKLSQm9/5cA4+Bn+T4HuT2g/Cz59arJPjiltBrdWysgnyfePmCI5IEp/e04Km1
wmTYOKyRS7eFZktqKhhPsihTqOHelL92CDtoO9iVFavECfqqzApHi/uGElGMOJr5Tk/J7yw3FexG
Xa7obXhvdlcBlgPt3zLBoWBpm6PTsGYbjiRI/SSD5kAE3PPOl5D3/90K7Du5x7tq6reCO4Us5mtI
bMgfG+TzzSi7vrvsseXA+DclPF9CNlWmXDkSdUHQ5gpkdPJ6Tj2VYh+kpd03+lmu85R14sFdzhEJ
PejUJYmG5gF9YeAlEtMoeXZJkODxRZ9hPM+baptqUqm1OA4zxccAlErTI8R7p5B6IuuyTR7hU23I
AvTFs5Fc8IBJ5oFPMA7IroxJbdIPN7RSpNgKgiViH31A5JQ/oIWpDjyMsAyMXpOpKIMzJnkL5SmU
GTU7LtZ0t2jCwPqDNCdo4RRU5feIPRfdPg39Q/iJYwZBvGGXlskVr6P0vJ1nNtq6wOpwd6hIroIX
W7AatVE8LvI+Ln49rNaG6fe/qzF+9vOlz6TKh2nKaxYbdwxR+lRXGmNMwOEWswd9+w/akrX1DwCB
t9qEhqhFOdSCumWQUI0fW9AXcPmAIzvVnk9Fzos0MX+IKacGUeGwtGzjbBQb/+nVswNXo/bi/EUa
fOJb4y5R2LC31PmbSZsQ0tvlRX6/Tu+ejGzSm+nHIQVwmhE8JxtooRL92hjk+su7TSBXaQCHPmwU
AyhWfpsS2KMwGr2W99f6XCFasnaS8l32csh4x/wxA9h2zKTSXWWMPJuzwpYCXhsRE+HMD9LOjwCI
bDcyWV8hB8fyt7Tv1/h2a72Uhj/48BxnNWJd36tL+RP4S18FcTGfwvs0yot0sDGWZ8zvvWS/esnM
2q5KFR4kE3CoCrvh6uC2p0oPbO/JJoir0HAdF4OrUEX47vXfI0blQhKm939IHuqyqPtuo2srk0LA
Cs6+V96Ao/jwaZ/3liYYiYtdUGAAJf3YmuSj3A64nTtD5l13SUIYlhcKDxQrV/+PE7VGGoFtJO/e
qjX6oKbtA9luCo0AHPAnPFdeQF79qHNDLFKM0AWmRzgjebvEraPRqYaJc5MqvJRdV4++BpUGoTpE
O365BPAByMDXQ18jCiG5TF5+AnD1UTTGjcrormlHrivKyUTjEanNUC+wGCH58Kr8KK6qs781Idxj
69jld9zxdTwGMMrUaHg4qogSwqWEiOwiwysE12869B62qK2IfYSG2yKKXnsqZowaWs1CGHWt2a8d
AsMBp0bhIse5kvSAcxf/6yzFnUmdVbdY0P0c0z9jHvtixCww3L0AKPCyuCMy6GBeOF6UsDfRdmF/
CFGgfrO+Pq3jW86d4VcqbXfcbDAdOZNLsL/ZJl4NF20wzpuH5Kf8f7RKQfrDKOD6Qj70mgEboetx
Yznjw8jeOD8sJo7q+dvnaeY9S5epshqh3/NZ74Wa0c1ORacFmyF+M8iXBKjTxMP7/rIVNUczSPm9
gBYOFq3ItsZ4JJGfZGT0XEX77FFxLVvtC49YFUVvCNwIC5sSyDPf4lo8f2TEE7j2oWVNElJHnUXn
gvL2W9LUL+1pn7vrliYm5Oq2I8FQJh5MvWtTgusQs0ylGEu1YdSOQpt2n2QzwgUFrFZNhkzXDckT
ndR0qKAaNVZF1nuhaVBONIptNUJwKBk3nDnTqGLC+CDIvbA6eEW+W2kKTcqvgFntggmVJRHzwAKf
cqOqb08ZFciZZKp8nYNXBHU45IrbfQ4QPqc8/nZ6zybDZLAZxTtRnkvHqYqU688JlVJkF8PcKNAP
JAev3ig8rj84iNxnZ/rEnAv8i7KDLioXwlsXptHZc5JJkGFq4xFyu8J/F2+xreAVfV+owLtUfYq7
WW4VHolgFuiCkRWiWUQOYa09U5L6buHmnG/1g71BWSpJIdhinJcNknkrvj9D3a1IfnUKv9ojEEAI
aNYTKd1LVg6emoEWXhF6s6LVNwC85CmG3GzTpxtMM/Uc0jK1NkEF3AgzZZAVWmJE/5wPuPZA5FLn
1ipC6l2g1eji/ajnxtkoXJfe1N85ysAposbfsBbbKhTzU+gzg3jQj8CGGLvGHZW6TbROwI1oTKuD
LQhSVoVEsNWhbbYM6fp2il2MOBCW4ay0tmwjOUyxlWZYjWTlsKgDTCPi5Z7nvffSORnNjo+JWIkg
lPfxQQ9YhSvnnmzlKW9iBzZKcjIhv7HBM8uJUECeXpCkbZnawbmYDyJvQL8D+jpGdsnl4OL80pkN
CPU7u56NfbtxSlOz9G7ins1rTrb0j+4Yn2BJVQrXvjh6eg8B1vJOtab76O3leWS9KOb2cS50nHsX
yFOPU98eQB37Z2SQ4ZsqOLGP8Ko6eN6yrxPsQ8+2ZZIk5tZLZSq+H+u7E0FBQDwlqIPHsJQD4DjD
h6Vo7uXnRWCgMLgUMKB3b35ecbAafLkW+rz+Tz2lphXIhhmH0voJiI43Yjlcq+yEJGIHqWZWsobb
rBWsCBxsgn3r/nJO6Z57WOXKAcNY7lgofvGpP0d0EpyY3T/2Yypum+SKuCMKgX95G1Cegsm9O3cr
2QzXLz/lYkB8nYABPnsUCFslarRaaYm8nRguYXptKgcDiA6NsXDXymp7q4R25YwVQo1IBTAYKtYs
pxyiB1oFEvtcR361pKBnEUaTNfUGXXk09IlYNA3RMLr3AJGuxRxUmkXJo+/vc9mUojOpVcL0YTqK
bFJEXHtKjC7iqt+zb/or+mCJ6QS+EWCMCuq4UFz4kl6vKYYBztGT7ASXEPrwrdcFVH3M9QlcyEe0
RPnJ95sjvUE8VUiMbms8Ls1rfkWMjA+80XcrhenhNNOo4rA1FKXk9C70Y5PhpdnTiTTO1a+T7QVj
6qKio8Oi1fF3gbqtlAjWBymn7hGnZ5v8ID72I7zFdz1ZVDxj6azACoZNypTG5P+VSR81+ddQpFRh
g4PQ8kd2hccUQWEdbLVDtdg/1QNRawvJeEFMW1NoWqshLksl8rOo4LP3kgCxHPsH1j4dPz4XFpOV
c+Y59s1gJANoJTWDSJWXrAWIg4grY4rGjm+pH0IpH5toaLCXbtuStzJs4BJnflkR0/ov027rzmhu
SAdQv777bX0/vkZXt1jzDBhiMh9Oqn0VhHerRqFUeB4Ty0YRr8clN8FXa/qhG5jkZsrIslGiVpSx
rqAfAwhJes/ITowZf/K9ozvryqO2VbBPYrTttXeStEWrp/u4NOM3nKiwoonhOCaqfXZ0KM8Kl/Rs
4cEeST44fxGoWMqPn30w1PbS8ODHU9L6IH5bSg+/Hdo3Z2X7lgyzfFqD1/zwXgFNax9x0Mc0dXtz
R+svVrKCeBBxFmyAIaIA6Dlvo50hH4l61n6eBLg8Vy4YlvXLatXpvuHcIGjaIR6CMMsQmCWVOgNX
jux9BWxRTfQzaa/lPWRIC4fZzs8cEUqbuiD2Hm7xfAHB9cMsd9xhudZsrhkGQgWz+0jXTNXYWSm0
H64Wzp3cUNgGl8uaWg0iQ/DRhBtJzfHc0E/zD/PufGNxYrTrqSI6VpLkgfLasG1V0W7ipOHIzYL/
vFbHcassN+WqkZWl2HtmPic6fVkH0X9RqxGrdrKSysL/tC1sYcGN8R719clTJdmSHbQRzqjL1MeU
G68KQHJ+U4XGVyCSuamTUKeH7DKHuvxZpF9XR+leQsMSobW5fxa01lDYyIF9jtk1mthQxz0dShUL
7WE7l7ROwOg0wLOQ4oiobMBAs+pumcUYh+jThVn8D4JK0/Q84GTQQ6MeN2DXVzpyDpZBVTXvrNPw
ZKSp6TjwojhTJjgIrg4kwbo1pypga3IJ49ngxmS3Tj921dIcLYiJmg9IenIsa8fMQa9q5QVR9iWh
0HKe8zEgm0IspdICxGj5quDy9xYaT6Hav11i8L/MKknatPVE5tk2GtNGO61QoxmPdi6/9PUnLVi9
fH/apitvktMMar4vtL5X7VX7MyTvvs3LTJR2ZZ9jBx4QXTgFKFe6Uo4Mleq2MRbujeJVkUs7x+RQ
G2MYMQ3rTRaDjSU6KVDbdHN1daMf0rgZck4EV8KaD/L3UHoN401fGM2fxCrQenNEt+RHKSHC8vrX
c367x0da/dgjIVSNvYNntRz7tY15nZG7emjwks5i1pbUYRU9vJn6vW0P77GOBMZNu66Dw7P/PQGA
xVgPItT3lWiTvrjfZ2Lsti4uMfkNOYt9FJGx/US9KvnlSqjwVwZpi+32X2EltQ3A0UWQE46E31cZ
bxPqIbiwAN7f7sCfPvPKO2E0JugCJnohNIRcYwuh6lmeGfgcsN5xGRx62Nr/wl8VVYFFFceDigwa
7dITT3rOqFqoxSOxCOsXeNrJSehE73Ds4/G0G0u+Ix119kartffpgk81KbNrW4cOCpwgGEsLo1m+
Cetgv4EHONeTOhP1GO9/1kFz8uVbDstJ/pWAZxE9S74yj4almagi++ADfZGJHXYdsuW/V6GkTLm0
yYA30jYvmbJkvejqa27PjrFjBJ+RkctQk0rT5Jx/7wpqLfXkzbWZUJkGqWDggl5NQIrK6GGrAJSP
dg4HlTox9N0R5qvfN2eluEKE6Zez3k4N+4fCzI+phHSck0M1EYnulzdETQaui8XGwQetN64uuKSC
h7nBmTI/GqIK5vEER33TbI2a6PTYIJYm/3KGPgZjr9Jly5a/nhT46Px2A4VEjBfKD0R72G2elsu+
wllCyJH6NbiyrFttpY/OqkMwt56K8OO5cT9m2pD5iYUJgRvJ1DNp3sOPyhoBIGHhdv8JtYIgnOoS
aM2qZMbywSFOR4IfOYkkZZ4txynpyYrsDzFmQtsg2xBb0M305hBwYXvyITWvNRlPYEj7UF3Gj9nc
0CBA5o/pQCkoBymmhSfDWVsF2vfbElHXabGSDc6bxfCRspVCsSHUNgCdzbU1W4Z5sMlRl/Ie3DDz
Aq7MogoJPTcmjb1C8O/f1cUoWe+Bwr8XVPDNTaowd/EOIFWhU9oG75sFLHVYj/oFJ4yJMArdkCwf
UyLKcOM1zmw6iT7ERVgHX9EI9ZfrvOdzFRtMItSzrwbnWWNGuoPUW6hAbSOPQT+bh6+Vzk32c4OV
KhOJ+9RLhHfOmzf6CatgN25smI5sIscgSklgJ4D7xNr0xtnxUs2KUzUSrLx/z4i8h8C2H800oiNF
Hkr/Otkveo7wv7t8O+35sF/GcYCK/xfVMHjXJcXd2kDHCaS4I1uBOXiD+s9wituabgv64mLjD+Vy
OZP+noX7sy1QU+3mAp0yZiqq8HBerELreRvbsc53Fxv0bXeVt6qr80YzqcJZwzSqTOGbUYU3fvCa
x595RQe982V9UCOjWqxX9U+OL6sc0aZNNlijI3ajzugkxK+uyuNx7aT5Rjne+r0FWhVbQmPpfo0/
FvZsa0QXttEuHXUIHTYqvvwoCnjqPVKYvnw6pdlbc2IJLLZxwRAU07lkBFGB4/1vcgRSCsu55Tf0
MmB4Ur5AkMYjrwAp8vSZvYHYhdasNXvU790oAQP4xjMXOHhwFgkcXwwqVrgMKd828cU5vgh0DjhI
1VDHQkxzL9d4K/f45hDWt20oFpxO1Oi1At2iEBVPm7gh57rRd/SjDUz5ikbbKPwWsoZyP0+9ortL
ZXfZsuWoNObTYv9urBca+8+uHZ39FjlseYMoEYUEyCOoXCEnpHYTs1iTqWSN8NENujuyYfzyfRW+
II7K8fpv0SvY8VGaLZtNhYMM8wMBx1n/BffgzVCR2pEW9E9HkgBK+qDTb0c2pzrdmo0JubSoxOTl
EWp4QW5+amFeUK/4XuC7O2sKRi0PV6t/4a4yG2VRaHu1wAXqz1nVdQ/oxSUl/TQn6hdIXmxPLlKT
/umqFpk03ZjhTpmMpmKtjDl/VrmcCeLEkqBotpuRzXBEXKDiAnnfcDipmtf0SWF0YFYfuHgegBLt
Mv5IxdHgxlptE5jMUaQbR9ZVPXag03gx6ZGuZ742YMO2fN5Rg37ROO7L6qV73Eme6peilyBjzUhW
CUFfRi39hUBQbbeeOVgTcbXVQbODWCRTySnYjrEnq7hfKdFN+Q+Nd22cSQcEvExFmZ9YCEly3LEx
CQhP7h57fiXLnjzmy8sPIbbOU6y5ve7unlqvDAyBgaEgCr6CgYYNN1QDH/SiXqQ14CDiYPSOILwy
piiiIVbNzF6ZHf8hX0YtJZqnoQfAqTlkbkeIz1p8biA9MsL8By77c6u5EAjR5gLT6DcgwlJHm3Od
wPs+UjS1MVpJTzpaV2JaihvtXXLMgcX0uvqeYqB/GnMZ6urJJgo3yQBIfnDRHsKmnfwaoZx0/8WC
26ZFywVO4GaQ+MlRsY4K85R/G/eJhpMchFz0kY50o2RzxXhFbP6mWClXHKWFndgODM1C7/w/L0ra
Doxucu1GFalLv0CySeUOIkWAcNAC1NMl06y9S8ezWxBKpggv9ZskROwpsF89Dd43wac/cL6anxip
COdKTEPWwTcn5Ev4gGaDRx6A/zvfjvy1aW6BXSN+QFKCQ1HNObJLC4JWJIazJv9NIzE8imqEd1S3
1fGmrYvvKwYHBTalAnRJH0tuwTRrERFhuX6xY0jqPQoERB359B15XNCfzNz7X+ArS3Ms67ei50Em
4KJHKhU2SMpFaysVVM4d2LeHXTe4FDFX/djs7h/X+MiP7rnbUknsLw31t9ppEiiRt0THKDfBMdwB
dsYp4HhbZKmu3V1/nXAwN4HkoAXx/FU2tJb3V8Hz/XBH1lQ3+ar2Y5Y9LdKcWwHwOmGncHxpzYym
TrLKUOW5yfDMWNKqqG+0ZU45ZZxEP0L+8iAgQCXPJ7BE/94Z9k6uoGrjVADmHWwKvZq4rvr5WsmT
pxPFRVCHqEbJz39YSjHOTOYwKOXfgZtQQHfYQMzjz5BcPWv2wpK6xSpG1rNeU4BQxJ0XEOZpOTu2
5AmgCe++dF8VM1dsWvt8asMUa3yJYkllz6st5p8R39YaMp6MueULUH5yWoBBgDfqzZEOw1MUTpHJ
xqP50yYGvFLDlhxm4ncUEEFVfKOcgmQ+glvvNcTv9u06EyFxXZ2vSp9bEPQM7Cb/cmHIyeW48VCn
/W05Sy5hTHp+yGjSWUhihPaDyqVgF7AOfgup/UMQXZowZXcswI4HjdLeS4H3s6Uz38b1u93jfdn0
IpwLRWtcuGeex8kNm63hf46ov9M57xL2CftpLRZi13IAIwIaNrxPum3CGXiUgVhrAJiLzQ5Ti028
3+74GAGF21Snxq3QmPocpJSST4FbrTsmm8Wzb+bx+RpqQPct0i9tGCrjv8CRfqVa4cQqIDxZG4nS
7ezBN3f35Y2UgjF8wlCqyMk4yfRJruqTT1m3QLVW7f1KVtpI/Z1xkoNB6/9GhYzfh5u87rn+oUoJ
cYGBCAVmMI0FcCOAfvx1MeMXUFmIMLyctWd9pRgKBvVlLwIlUCyivaU0ILgmFoi7pYpPoiTlzrvL
cCMOG1lAa+O+yx8YU1bJzVjPjs6XFxVDkJf4/ZOeuefMWFrafa09K4xO6d2XAGVA3zlYBQheEPdp
9sE10N5ZQS4kMAYf4VpubMjMN3NGqUbtU378SusRVd63iTKhrVM8oRFmh6yNmfE5JYavqSme9mZ+
V9fLnnywARdhCaE98ew2ja9Hw+u5cI/JHZyou6DVRIlYAkblNsvWboxJ1LReU0jQeWBMjt2x3zBJ
XdqtGayKfKbMYAvgkdzA+Ak78f6f1sPoL+1UQaM2b6RvzsmoWkr1QOlfSOIMjVU6tHdiDis7WUoy
dHCgI0qgcLnoNh3Dv3mfD2WhODBegoUFdVOig/aJ3zCWaUj90JcOIoDB227Ssff17CK6hp/+cN6d
Ic1tc/vljwIoRfovLc+7m8sHEckUvgSck3K9QVlSoVNICfTjrmsBnlRAZovR46krsGlEVflAwJfU
I9rBsZZmRnGZhIWnZXBmlQfY9uj/vq1bdkUB1nyZtDVZRmNifuIBXOUIJ/zrkwJVxcjV8wWiLAm1
XuiL7ewn+IqXcZKdgO5qUtTWXag/oYcFyhg7GfeNWg9eTXT3G/+dUbLoyM20LAnBMGuWeBAWWjMR
+vKmYFuXL5A08Vxz4U/Mi8Ev8WMK1f7+9d5fvJSui7l76bMDr6AOJSTGZdUuoFX8XjSbeqVCQvMw
poBTVpubnCAIYJOQ6pv5h+3HPFjcxK5oQNXyfMAwC2C0WDzVZEfFUc2pFaDEsjrvD+AoY9z1F1r/
FyOfiPFq5yTQa/Dl4+SVWRdF9K6MSxSvigLzhM+x+RtK2KL48iqFUOWfJG5R5ZpHpRECoNhMfpf/
N13KH6ffMD9I399APmnISt2Oeglaq2a8SIzIQvEYVL+UC7zfq83zvEeAxpr/2au4Jtm0q+9JDQRm
r1D6hwOy8RqCrmuyH/jPYH0vPbUTd5oOYyTnakbRS1WzfAmk9oqcu1DBdeZb1+6OlDpSsp4y61IQ
VNAfT9vdmd7xxvNVI2SBxcoU6Xga2VUf9XVQYX1spIpjoKNjhdCXWfMXJd6SlLimR1s02hNzlAv/
jXXE/tbKpiB2i3Q33+cSjCGHLYkW+Hgcm3SxxzCmX9icIITE0m79w1o7Mhxlfx2AQrKLcPhjcj0R
0jdF/EEmmKg2yno6OQ/QHHQVD6B9ENUBSEO9lzOfteQSfR3gsp1PM5aZLR72C3vdoZpWoMToFy++
9DPixPlGWYH4nlBZNZQEL7W5Xi/z3XTK85LwIkmRXaQy8UkZDqbxAIc23qM0KLHkvrmSSFuRN34I
ql0F6pHfc/8S+TMRl8u1bP/qx4A8NqgEWYea4vfr2PYpBY4+oQ1qcCD0HJtJuMmzK7FBXzXaj8kf
2iaOgJugDhAoDsN72lU6Ribek2AvkUqg3pxonLOFrRyVv/HWEqkT8lr+l+6QspTXIRBKQWfJEJsQ
bQBc4Shc2QcjnWVKC97IwR8CYOve8CivHSzMog2RBuZgP7cOXTVQk6v666/hHlUfusYyCnr+iJrw
+8x8zo5At7LUPZc16ymtXwhcEdloWlpM3wNSCaOzKQI2R/nbSsU8Pm/DGgaJ4wY0AGvCPf0oSqcY
/vbkKUxTSeIMz/HcydzhbxMv7muTwfzdSIIUGmXoFwcH5US7XwtcoUu6YO4rhlxUw7HfzyoKc+PI
XV4QC4hCFZ45tWIbNrxovpRcyiiIv8DsNwdVV10fPs0frk2AypOCP+fcLQNr0KVIUNrK8LnUzOcn
zFdAPs77WngpwEkVwC5XkFmhJ3oGCeF7eCUPkOrDNRwAH2dNWgKC7um9oLS6wWHT4vu14Y4rl0QG
ZgJunTPo576LKNy4qFIQW1mPzq0P304omVQKwBJXatFDcO0LAa4A5Ygjz2R0U1LKCD1OLakrIUt3
pZKsPzrzi2i7c2t8k0daPOQGM584Qmor9l9sio0Prznq9sSlAhJQNwRkmtdrmQxBDcgt7BdEzJth
UEGB/t7x3VfaSRklo8ABnyMbJn/0VCtqLZhDYuSiU89lOgV4pgXpd+eKLcza3sNMLP+3v+yvwuY+
OgglxB8lBlVjFOmmoocHYWZwRycl1NQhehqbctCS/ATsl3MSkBX5XLH3s4d9ebp9j5MP7c8rqJoZ
2eK4SHoFbNiD8WFVhheFhGsMWCYVwu8qac8HSbQojIHYLg1MHItYjPBstIhuRo8fqWCANbmzIFz7
/jeVgJoTu487TUMJjxU7L/02z4h8NOqucvtT9gf3U6CxJxdoYE3dqJZOflQtXFDA1l+rzrdEgR29
E3opjnjsfqfzWiz360WdSc2ZZcvjLIWpMRh9ATApEH9f9meS+/nfqpqSb0hNnQ6VWYgsplw5Qd0u
cBjN3uDizU28OUP5+7Uh48v9aA6lOy2bY5iKAvm7YHNRL+o7xEebWjCb0/b5F/PY4TaaK7tz0mKZ
gey5z/teIiZM0d6gt2XT6Vb7PrRCy5tNNPPhIVqhd+sRN47FiJ344yd5FpC8gC4j/5fpAn99Ct8P
W/2avOMs/Nvs6HV/ySNsfJ9IG9DuOKDAhlDhZs+/MmjVOyH4QF+vdftHOCaTnhragmGGqrsQ6gwy
L31EVaPE1zdmWnWnt794dxqD7xaBKRUAiGmfKttqcgQgtTvO7scIhzy8j5l23TaFFUtKBKD4wbMz
yjn2rbDZjq61zbIBYsPeYCkuv4DfBIcLES6VkqSFNzeIFWYB46zAAsnNK+p/X92jPiE64ks0r0Wg
qANwzVzeOnOovHodM8JdQrp2MowbjSTbQuXjeqL+8shIFK1RBbmw2zAWkZApTaEXPZRU0AW7AEgF
MUa1ax6o1hyUit6FOE827wVJd/spka0b39OCVBUf3fSTN0CY4ku2PImfWtW58XhUECPST6GDW5Kg
F6+IwOmIzeVyTM3obkUtOxOBdcDeo74nHV54+YpUiEnjNnJBEw06dIl/BSrQ0J+H6cy8r5RUI17V
mTflbRyAM8cpnUiQDYPgDCc9PrugN4oZDYv/jj3Q6Qp/8y9pGpwPjGVYqmllO1Rc4msvmvl/meJ/
bNXgHeszoLIRXXxaOnUg/7Yjxi4ObyT/VFhlGC29Je75G3knhHW+8tVjOJeWNOOvkh43kojax9s2
kV4rNGLw5fucH1ehgvPptEgWwCbETk3CYgeXCD6CkMisAAxmC8ShU/pC5YN7aaRImp9dw+kh3fO+
LwoSdoTgEbqsHuoYCa+la6GLISCK3WqGFlTY+DPXt67mOjrrp1a6uR+t7HryoUQG1cNfvS9N3gsG
kxjOI5CHfsyJtXQDSazeUwhU9MzLAxga8jGVN45GEhLnHyYnGEIzWUJ1AT3bri1iCnyZZBCvJyD7
sDv9BRFS5thslTfgQRgYqvJqOMbr2XgDgQdp/FdSkq4xEcoRxAujM82iqkSLlVTBR2B6/+tYlV78
sLZ1n+CqKhVUQVO0lH1f7jGImvLdlXzHNFeVx5Gj2pqmp0jFgPnRXgqyOC+Ybrv5YlJF8aTqA3CE
oyUWc41yUHT5VJhe6Axd45yXQRffIY5t0EHpe4fzbXeeaOq1hCruke9kXQoq4xPgVL0h7/CPOcoC
628kAj+igsiVkhrfB2lsRwlbMpSXq5imbYRQ/fP2MOrYOBHr0eJau7OWBwFvijrJIfhjwZs2elA/
Oz586287ght3BWjMlzWHMD8xaBlnYDd1G1K/pobqNzUTukxtn/UhujJL6StHLtLB9Ctd4tAj9bLN
JdqT8XT4Vbdejk9tObJCI5KGgSkK0mH0piEC5/J7/YHofSef5O7BJppj/ypSaQuhMaCVmTI2AQiU
kfg+wd7TrzefjCaqO80ATN202vXSmYoqtBRsMXHihgjLbk9H5xsh4+p3W9oMYfJABCWEcQc1im2c
DBcI76EWm+BF4pLA+nPx7ABhPidrdMDTuCNY1hutdKecs4xhHhmCcBjVlnxbNnIkOfYqQX0kCryr
Hy1q7Lw4exgq5dUAM8WPQbqgB3mc6KzIY6TgdQfhrNZXC/0gU4gSwr5q0rtgTknoCwMRXnesbO70
b/T+q34Xk4nEnrUxiGO23g+3WZVce0gVSlidbZPZ2O2Kueuj/QqUlT7d/PRMcoF/V6bnCmVvclIt
uOLXL2Qdloo8fIkmRKmztRHRjYW56KqO1FsqVP9D707JZWkMmNNs8WV/EwYBPMTJhq2LR5WEmQuv
irT2blG/04Htz8adry4ecL/LhntE7iPsvkT87fLiKgDGdB1o73y0QJqsF/e65Vsr2aadYhtIyypC
XUaq9Hqf0wTfM3S0h2rFfQNyWcMnrSv3UoeIjfOW5tPgdIP9OfX0qhdzExxgS7bIDjuNakcqli2F
jk8luhJIuWAV3cZgPSb3xHQw33I363iwWZfXKqQjr/qBBeeYWJa8otT6YVNCHRvolrKFhpaTBkVa
agR/dZAOUxa4MjyDpry+sMTc22JllFgDjhM5zSC7icZltezNeOnrZqMoDLc84cNhQ3lZ/rWDRCli
xsk9ytcVorPVNah9XUjMsKvJwG9N+6M4U95SFVm/ygMfeF6+jaHXuAU3dQ4fXv+C+9Jj9QytNzFt
tnCvUJr64CAr2MxhIhPqeS1wyh5jX4dYhYAg1G5K4At1dz0LzAtY6KYTOdGnvyAPmkY4QBG2yGo3
Puci8YPH4aQCLPZqQmN0dOvAlY0b142LCL32BWgc+GNrSK5MWVAazXmeKXWBknipY4sdnXU2MfJ4
JhL5eV7KZRYBhuA23Vw8qPDPyefntPtXHKDW+394yeowCE/KnP3YpXF3s43W7gFBH3PcOg2/j9yi
J2TGCndi6RHZ9xTnTHfRTDOHrPj/WHMd/TbGuOV1KLCbYcDq0Jhvz/vOooNpCWtG+t7OELr3KJqU
HN1I9bu0iL2Vhth2PjeqFsjgmkz7+gUyhAg1xTui5tidnfug7nQUBmO1ppoJCO68j4XTDYykAQYZ
u0tCdCbr5eDEknsEztKvCe/08qNjZcMKo5/miHl/ZlCQ8EVtkQ5xxrnWJo1SJv0/NEm+WWkbslJO
q1sDxEImAf1iTtJJ/t0jf1FW28u9nc496pHPuRYbYZWriotH3cyAqW5FpbSNdrzw6NQbdhe+fw6m
8jjwn0EB94eu5cTP3LmA45CYtfqat1FP7OlSDdKI3fcd/fpNMHNQWYLRcyrFqswxun+ENLPoPTAF
PfxDmaqoewH7VUylCUJbulN7Hz6MRfbaqHc1O0N83QMiOHxzRHY5D2trK9SYeN/+IhYnmahpP94Q
Ys1bm4gccx/kRnelgwE16yxdbVhZWowjMekYsz/siBW7Y6oFFhRZNp+i59syqzdiAkIPeLvpaKgM
fh55hdBkM6JU8RYFeZwTSxXyNBwdg+BEQjeMDqKRA7cKhoio1YGYx/g65hwc49+Ug8z7bdVnRe0v
PMtxwKadOeffeYZ5jdeLrEHcPCmcuTRIEa+GnEyZEZECk4DIn7do5oLoAGiCtdjrQTnukM/WvWMZ
znp2ke7IgAf4+FspghvIr4CQ4C6bQUU0CHa2liCkp8cZ9zrOsy5sgIK/1nM58D5C8JAUsybUle1V
fEg3X+eCHzmrsXRXvyZPOvCpjTtIhGMhQIUtNOvDXgqDTWBp2WYiHPrmxbgOzDIrVffG6yzLX9JV
D8AaVdJh8uLWhlXlCzXcsJW8FCrnXpC/vz2b+zjKyqgxndp0k7qkxDoJJwdmikblFscg6eEXKZZF
/0geOPBiY7IoKjM1POn5+4disrXhKPPtdyDZ5J72Z899+crIX2FC5A2osdR0fQ45BK09BIeRrsJ2
czM3Q6CnydSllIjY7nQnzEu/W815DpaOvnPXwzm9rt5bXBKEfR4ekYItvpCtWuQKzHQMsRO3xwAB
EtrLnyWBWePtuaOpJGcn2i4H2n908+xYxLZaM9PEavJEpp2eJJmi5L5Qoc8youRgu8I47REXxXod
tzicq7gzRBQRewTj1qj8ZCAdCERbJEqs8LLmf5gUjY3ENdF3maZq06OVeG/6Sl6bZI14SgwVbx8e
F/BY4wg45GtReKxNhlXOdOn7mu5W5RY8EwAnq2wRpRlHcVNwAMjrz2XDU5SHnK5pDU8XxVQiM8Qa
/TZVHCSlhsAngCc2v8qeR7TVj6Zyx33RnzG2HhZuFo/1gks/jjXAiBTCnrY7+jNG2x9cVG5C1ukr
ZNQIj5YGMpiCaT9JVzRKvwDmWP1UanKKMdpqukX5a3tUQNyQbPhjQDdXFdZ28wev35mbPWJlrMYY
9Hueuc1XEt3T5IS32Xialeq//5Q80l3URWkDdKaBbaSJCAC9GQrrnOGFWYYRWZRcgmANDTLdyaAt
WjfrTYRzAZenYAjLEZ1qRJr3cV4aV9TAhnRCL7xDVZ8W1sUMw6xGTvh4kHFtIrlDHb91rPyzbUBo
nPOlPzc0k2toZLqaQ7+LAo8glbXlw5+ievwcM+QeXpVYtV/tYeMBdzCIqn42tO4JMjNUCn/1olpK
2kdpQEUHzaTK2I6qC1Culsg2Gtoo3+8zjKfVhW/z0tFxdzLACFscDwNRVvBBUQVr7QGUNTObP1Je
pn6xdr9EGtv61DELV41s1pAX53FGoldoC7Iqaf+3MEvJwOq6svEmr/2TWKdzP/PguqgRmfYLMebW
mr72xN1JBmx5VbHkhe7nMSsWmrNXFtujt3lAgnBrSueQwcekn2qFx5YNHL++duycCkBmw2CcEvWI
U5ZkG6mSOyTCth7MJnPx/GhiwJJueKhBnRSoqY1HJ0+5162I66ENoieoxZZ8w0I1mx3UM4kMHRuA
0UiY4V6A7zGixzArVtVIgdDqUyu1+R8p0r1IoKUWf5l6Q99teGG96tkYJt8SW3mVptN8LNnFjciE
gX+7NM7qTZ5GpzJ61qjOfqFMVht0jw4/uof0nyq8scFnwExEhLvC39/oJXvRHG+wEmiZU4cXVG+7
Gcdepss+TGPCvZIfc3bnwGHNPALxeIceHsLcXsp/I5pLiitzlZbKlgjMXXvpKC/D4AJ7NMe9dr2R
pyTFG18h5YECuYQjz/zQQWei8/kL1DYTPfu8tyQ0nCGexhV75ttmhydbdjAzIUhCihJ55Tw429yE
m//x6+7xuY1fu1gJ4W/gEj4AE5stziMG0rKIde6m2evPwnL3iIEFJ62DEQb9KTT4JWSWy+o4BxHu
AP2+p4uwp86hMGfLiSIoaASkg0IReO3GAjm+72MWKQ9tOnZBZ/eooTV8YQw9jJxylGICM6y7HBp8
/5aSVL80ERWvsQY0sNIwFVtTN19EX7l1Y904NynU93JhglvgfLsQSrF90iUjIYl4qxjbPcaTE34i
6Z9sv2uo377xGiBwM1KiloBsgiQazfZz2Hj02HFU/Y4KBNXNUTUUNBh+i1zaJXjzNAWuTp3lmd/f
kTdyiRyGR/hb97Zc6vNlMQ0Fe4g3QSX0W6RtdTEQt4yG2mAdJKlWooQ2w05i14+DMKbJY3fOvWAL
X+Mhaa0XQbWCQBukzUnqWEY+poi6WK3e/nvZGDNDIzcP+4pNk+LBbFepNbN3WWT+J3re6N/5pDVQ
T6hVYUTXCK5iK0mOTbG6J3zStl2f3CFfk0msdHoHv+j5dHU1/WTZs2haZ9XFfSK9K8iE7yKurWn1
oOROCI2U6T+runy2EZmyn4D8h5l+3CSUot689VtGdH+fvXTlcQspnhcd269hp2/E29JWFrDXwVvI
LfET4yge6IUwahTcIjb11YnpkNNlODARAjPwtxa8FgHzcnZrgZLNpGOmrTFewmvy4uZjDp3frxov
qQvnmrvvAg7LHA91KhKFwVD8BiKs2Z4vpPHbut45xrA/aHl7DahABQ9z59UMgn8udjZPTkXKLgD6
LTXqDHHC6/gDS15H1XcBQsKv6+AP9c06yghoSAGPnow2lJxDxzV0NDb6WFFElcEsML4D+1MWnRKv
tzQy/XeZomsdfsqVbK/NXLZX0FFuc2hPGRtIg2mGyyqdWe1XXLvrpDnTmz/CgFmY9lecHsDYZXeJ
Y5rQwvikTjXh66uJhZ+iZ4GDCcmG59NP9+EyTa4mwYyab28bs/gKfalf02eDZgto6RnlPIMpqVN9
4BhyRdTr+w/sIJG//uT72RlXI8N5htO/QP+yuBgRzT+SLIvJ5UyNaN6BNFMGS3Pc/LwYoUNGxeb5
ekgGEfr04vD+NN3cXu/KjJGtOw+JBfUn4X82WRFxotkAQrRChUXNJ293ulAfLr5D/DuJ8woFEZEe
BuziolFcaX3O/hWOUh7OwurIVMeXLlFa5NU6EYOaNfW/2Skoyds09OFZJnSxqb0+KshWhhsITRWP
C5TqDHucGYHFQdtriXIJ24BrDRQ6RFLHFINy32hOC7ShbZxK32ug27ilDrrmRLD23tRyYhiNCayE
8jPkgSz/uWK0WMdlEaU9iR+XUgMjAyo2Ra4ZPW3Ztva/IQf6A7jNO9n54hoYrbMWun/2YATcyssZ
Scv/FqPZoVoEol265/NTTFiXMMSFCVMl3aiIMca5ZnuclGLhhCX6xqv0MKp55tdm1XcqEQYYVYY2
icvuRL+OtNncmoJWRURQ3rg+lg2Z+xT52vYXQVjAfkgVUSz3xtDjj/8+eB+/amYmg1ih6Agpk9ew
JtM171DuGVKjPLBHAE0B5CyrEV83u0E2s9iR8jzv26l7A/bvKKsCcPaSD3LaStoWWYgIIWDY2abV
olmYc/xmx1cFw7Abxnx1Xp/ISVx4rc4o17kSKBtrjaMY2KkUS87vW0QyedeARsaNMv+dLbAueGXr
W/5QnA+9xSr5EbxjZRatXsS5MiXjFiRj2qzYPzqOsccFr8RP6igvnpxxPCkQjabgmSuj+EIt74mC
g0HCrHQ2demoTh5mgOdetjdFIsFhpeZt+xbE2exrxmOr0+OCTquPpbySOKhdvVQhWGVrSOdlCEFP
u7q61QK0ClH/8y7ep/aU+r9KlMIx3t+4Jg7u5P3KqhZHmMB1QSdMxlZLpzXY17JTu/jYaFhDYkaR
q503fiRFqj/3XSr+Bt6SZZ+rYmiwTomA/AXZdzPVt/eEXVbeKwB3Yx5v1CTFGqtKsHjR+NKaNjdo
b6V6AUE5/LWGfmM11lnLIxuDlJSPOzBTD4DIrXHqcpX2pu3lDz1BOjKhNvbRSlPLwuHE1eFfvO3Z
GwEEjOlv0ZCrEljuDBSF8RnaRgPF5kq8P85YM2nlMlSR1TmlbQ88RSqVmVtE3yBSzseYMgHQcYIB
4dTCdlRzgE83FsDKYOgft7L47Y1evtI44QcG/z61Kk+GqG9q4cJrlWLziAVkpoG97ZECxnvfCa/c
11b7bW+K00JJ9ZXmjIM3c1BcUaREqwh978G5Spbr7OXhq4NRUti/w7IzB5ldcJF39XMoDRdv+Hpk
PJoiWsSrpoHgLljJeJjjyiD/rErK1x1YDnyNb2kUOlqCZ5kqhclQGKHK+H0KekjYuWz0Ezip44TB
HfYLzxvnnjBPcsTHTK00+poCpFgIcIk5pXP2zkb7tmozYHzqstuddtn/cubMWBMPf6Ay38yRB+ih
y9qx4dL3CXr0hqC3N+ur2oZlji19vpIUuL4IQFLKaagM7+gnSu5g/Qixbg5lax+v4NCZppavg4Je
osCdJfSKyPzSq12SQVUvT/z4OM9Av/1Yz0augs0MC2UVG7IDqZjogSUtB3QdStyUo4ENrm0EyH3o
aZ14GvX9ujwniL1vg4Z7fQUfmnh0qmWoJRfQ/Bg/gQGz5DTus1qAg85sl7AuFdYB4k2DbHb5B3yc
cSgfCJHnE21XnZZucS0OTiFXeXiUd6BVB5rbZJIVjeX+Fx2zOrD/NE83aIHXbcfGEPJHyC3KwEb0
YRskt6b4TxsgDf9AdFNr5IxA+Z1qyD+MR/NFjpjOgzKkWkrsze3lpVt9IqWy4OzWIS5WBGAoXW2m
ka5UKXTSSlqm+xile4UB29RM6P+pWbEr9SbfspNv63jx3oxmdKievtY0W4nzDociXYAYlJa8vXGu
6a/Qm9hiYzhY8/aL6e2BGZqgYfRaXBVl/+RppdLJjh7YdSYI9zQ3c6zuiQRE7wF69ZlhoznzdHMD
jcgCgDKEoQF+t9pV+3fakFdL7M8c89dCm1pPPtJCUX14l4xJERT37Rvi3I5uxbkQXHF+jzeTd1oP
wm14cRLBy9MYF+z4B/yhX6RhCF7Bp+y93V2xBLe2x3wF5NNbFuSsDO7JDQa07RiJtDsBLSHWm4iu
GbdYR12K2kW6sAv59uAA29s4LicvJ9WRcvqy87QRIX0+FukZgepNGNXsrFCXGQJaTSOcNgLFEZk8
QsbhfLHTiWcTw62dWvCLuEgeiUDNeqqJ/+rGvczCyjNFS40+fMPakP+n0CoOkhXlXBzly79A4Phm
uMnKSjTCu0HRoDkvOsSBuu62Aw84KiBkmzewQ+U4Ghu4vI91UGxlhnq4k54vqww1XwMTdMF8GyO5
ZI46rI076QIrdqcw7Y05ggP7pSr56vDQGxBy1d38Ezi1LoK9aoADiHkrRjzL5dIj62iC59WXL1i/
tiJZiIvQMME6fhDvu2WElJ+/KQMdFQPCrHSYnkpjHugNJaWqvoaeFgCSSmxT1jjEM88fDkawKp4L
ELtlo2KPGqSe+/xs3VDsCrvnwRJp5nDVpAHfonpym3GpkqY1TrjDQuDDZdR09u87W2LJtTDyHw4L
LVJax+wUAbUNqSkiIumziET9APhaQ8Ns2sp/S/nAnQ5CznLNgUVsgjWPHosxskFxUYdDkx6vcyq2
nO2iiO18U4C4izImXM3khHP1B+31ciSVN8R1XZT6gF5itndUr9GMvSTLvKGmL0L6GbsVkd3+nRnL
mMKPehp483dY5TOwjLGd2tL3oB0bRZkuoOjemRQyFc95aVjl+I2QB7yO+3psxoLMLrTkXSx53hOC
AWJSjCXfqtvcphsufe7Nm+f+aQbhfck9ZkaJIOu2SMurnB84pfO2UR0gOcOpnFGW4Xg+i5jz0D2x
pQoXwlEk+zeJVCFBkqqQL7a+/l5bkeuJzOuYOuajqUfG47ssjjOXkvWaHJWY5O+roHgpbFJhkVhB
8j1bo7hzj1B7BWf6TM/02MV0t3wnPTv2/Gq+SSaKlhThox3x4qX08izI5iPemrial1xhZF58FQvE
TIkCwWOk7vEXsjVsUAP7CHHNajeqqzLWP27sKR064FvtO6fdcETaGGtztzfumUyPUee9V3IYTbP6
NZl5XFpRw2Gin9CsVDEK67b2IwobOIveayvAj6VagVUvosLSFQeC8VGLLoLvGbOH+nFqNyu9H+qA
R+144bqB99dU7XOqqExiz2UvOa5KzUNpEr/OCPjhYGFilhgq8e+Eh4ef0fWDI6LXT+4uBEbFH4/2
DngSPPzzQqXD5pXj646YzLybvQ0ocZT3TF/5vD4l30HGuNBAoDUFEXoCpg/AqJM4ssm6dmr+T8NI
D3LNscj1LtqPWeV51n1i3YQ6sD177nmvgq/kYvXgrsnunO+qfKxFdn44GhcWfQAgUh43QHcIwXsb
gAy0tL8nQ/rcUY0Myysb4q4ReCvYlw0msldHm46Ngo9Dwu+KaFfXv8PWexTU09AI2lYlqBdj2/e1
SYY57NGiy3rxaU929mW04hCEMmTjlZihNRhuHUhrzRPG2F3lRkkp6EyL+xMh7GBkDyM8ybafCr3Q
X2WshchEI0OLKnP+b7hRm/8+7I4IjhRLLpzeG8p0eBCKXa3BVpTLELBqf86rHk3ngYwjAcBiv62L
RqWFgN0BSmBSWCWKvFZrS7byLTPdMxDBlqAJ2L+CrqWz6sS2iS5E0wPx90BJJT6n2T6vid7x6/R6
/+FYYgB22mA+pSfTJNXgHtbzJSEkSFnievBv12jur2Nkw8rwbXThfYBHM6OYtlBr/u7hvDoU3A00
PGzDmoahQAsurROLfjyDQAVmUqhs5lxq+8CXuRQreKl/7UnG1yr3ssi0Lc2E8/XFKzgwkK9Dl/3t
3p2Fw7h9hb4rt412uk+OFAIfm52bvV1vjozPxeAP2tQPHeBP4v0glLqro5amfP7enfN3u74j7bHs
ZJ2lpdi+Tn/IkqbY7ON8148xGDKn/3IWIVZxONfjC4EJ55JZGJ/BpnYy/REC5eQZJ6LJgLMzuGJr
3QGGFabUd2Uz3PwG/5pXkd+GtU4Dvv6sqyRfmUfqdYujIcFbR/6qeCuq8OoitB+nFnN6/vtxtcRf
ZiRGcfdlYYsaMujltrm21PT6gZI89jH1tvru3mjcBzcxbqoBzg0Dfb/gWLVpOhe9RVMPikWgaETf
XjPF2UbTyCLeJouB+rttJJWeOEqV5Wm7hL4aCMexeOJmuDiHpeZpDSYfRi49pLdumfWlZVdfP2Kq
V9E5pEDc8qreEcIvKrr16JedTutStwzk5PS2p+X5fIvPupfNfeNK9estXXqDOF8bEBVPjvkEYgwW
QzMQOy3x/eO0aw4UqTD805MUj0I7vKwJNpXmbYAIqc4rcVu+bHfSdoraChgsuEDozjxLQSGGdAeH
AUBhiqJnXwO395iWOil+I3V1J0P3CrlPz2M9gLhT3TDImOFJmMxK0umTKYlJEmsmDFR7l10hb1qs
ZSYEBB1t1CbOBHLLMiuqd2U1XMfNmjZn7i0zV4K4B1GieH0sBQqzTUbhzDeE+e/vXF5WylFezReL
+nA/7yX55k2oFCHTnLePjmL5nbmGtprRD/dDja3d7NDBfLa4uSsNuG20uHfyzTrBG/Q3jI80Zfqk
7uDGB6jpjrIw0htS+Ag7CQXXXb2Ua+2KnRfeGnAC5p7xZRyZ32rILjoZ76NYOXfCRMD9KanwG53m
qov61GHrB7L9WGiKG6QM9xhREI1aej8QM2yRFRRK+s88AeRxcv/HJMXsYz6XxTFpzEA6mw23LI7S
vVxRF0MWSmLCerytQ0ju1wkaZc700h1TY5kizn2xDxlBF/uLSDYyUL+PHhhBNZTsrOWRR+/5lCdJ
ZKEMzfKMhvgo9Byq5GgolQOU7K2KDJjyf+z95zXrcs5zcVY7tUwUw1QdOddlWRriSFi7Z/ljmsHY
RZU8DZXe+aJwNv0ygjj5kZbgJ6zHuI+agavv2uR/9B56OX3TRoeYq8spXlDh2hmJyCx6oYEahFl7
bKL3iPuIGw5NxD4n0315rgVzDwenTBkHhEKsLb8SwF2WxR2tkq5talva9hbsyc9K6oAgaFPI2KjN
b4o+rOu2r9J5jDV5u6m33UPDQqMjAtk6Lx1xtZpSpPgsJKXivXv2qW65mZQqdhUPsRgGSKu3RXei
BtXh1K74/OI393xdh3BoEJItqzNT70yrslLaqUalRwABktvQiTuYug5AVvGdKBrZLNqHgEUZgLqw
q7ttY6HxW7ZlG9/37R5QO5ZhjUCapfFCP/gNs2u23SQq/HB3Q1EH17wnNiug+Kdgffp+XOEwA0QU
woQ2quoi9KpWf4bwnjhaeltHyTcg8SqHoZxIBXcyyYUP2IVMnFqlKQ+D0owFelkFDLtjEtf2l6Yr
EFqyPDRw/QfzOtHyDCsagUbkRQL58XYx6JkmRhmGyE/tZ2uWPV9I2rrGlQWVgMXVULcsyJKLNqUE
n+d+LmaEwd1B+4a4D+xVM2wIuWd4rlQfaZN1haqPjiv2si0Gc6MA528QWDbgtQbsuQ5pepcgsJgD
Sy32SF1ntqg1+QEGG+umOC6CLNwnUoywr1EcbcZ0J/smhgIduyF+hbLEhPz3ZppYorV2fBpwAv/6
msWWyeZvaNBk1MfWq3CofHXXwJmoU/wjkjhjeSVH2uqDnHl504shWL5+k5PJXsQQtKDgRk8HBKPS
PntMpOLMv63Bcd8iNiOs9Mi2eefiy/e/arSp2bTVs8IQewusyhwoPmf7pUBHa5RpLRXffiT3SZ52
2Q2MSBNWfR/SH7nQO1mYfsrBxY46KPk89e8IhB6EMls8f8hSIh+qzsBqLMSVorZKSQtlDdn/sC1s
0mGQNTR+eDOSawMraVBU1TJ+/DyqDAOkV2q7dFQfwIH2kDxKiL8Zo8iKcM4+NDHj9MvpEb+XjRA6
FoGtxIX8pNVY2lPHaGbLRetlYGS1uXZBA9yWfWfVYR5QySCmuKmUOz4VViJnmXvrziaEAQDpBUQD
oXFtfxwBPXbeUDIYp4Ir6w9r6MlZexPTDhQ45VJpQ0SLYJMyeGvq2Wm+2oB5tvy8hPGw/kbo1g7s
+CgJoTfvwRPILGhFTrUutFLyQx8ksiQ+Qw37Yi4qPvhN++exoHQpDESDNs4m2mx7pTmco2/xscak
dUq1WFnbVnPmhC5dmPiWjAF6z6MuVB+yjSK9e+bsP88X3yhYTQormSwKSOk7oiy+GLbrFrErKxJk
He0wlVKPos8vpVucznfV6WI9Ee6FfAnHupBKZa/Kskej/wsTmf0G1gVkhqA4RpNgxgAN5nGNG8/Y
KilbRk+WjC/tfbFOsHgesDQ9hg34LIcIXqJijkIHCmX1M0x0zTwT37hL7mIGcg8waBDdIQYaSvdD
4wWFarJU8DJW39aK/8msVKipEgenmWv6qW88pkARFdXUa046TBh/P/zKrrXJb6xkpD3vmxVh3mfb
vwgolABC20+IfmDW7Sxg+MsMb+/Wq7Gj1pNGRtoi8KvXWp3MrF+EIbh+/eSoCfgmsj7qOEE7hrek
7RoyZcoj6wNeVsjNuxsZH397ea/0P3ZGJUYJKzWBxzrvLXM5KTqrKFUKet7ksvcAy4ZKPxLYfUlZ
ARXUuAF/Q/PbH28A1NfLGH0VUDH1wlvCU5lD3VflOA9hs6XbakxAXWhOCjE4wfSGgCqkSbVGJjJX
plSX/updyxO7/4BmwgfTG/8TCtJ3LR79yUjUByekF6KQQbDuqtUrpNlrauvAii6SiJ40hnAQgZpA
m2LasJ074tc2OjIn1SRYFO33v9dWq9UcpdyAPT+3XCZyEAuPV0Mk1um8rXmIccqEqMBYx8ZSW4NO
kpr+KdFN3r9/8NbwKiPmmAla1+48W7IvOf9O9GoDoplFNgpvC9yIt4voXOF9pHdnTXVaz/zD6+1o
pcBaEUz7mOWgLNABcd2azz4XDIc1vK6IkhOfc3D6sJirwMK1iOaDO7/H8SMTRYXDvDF5QUnKYC1x
5L59Q0rhaQcCQ5ulFQIOKtO9v55aexo18ht7TyG38pDYrHFKNA5xh5P2StA12kNhL2iJ/Q9xMNFV
Hf6l+L3n2lgpTKoumNBVV0qiBmGub9QF9uvG2LAyI3PNAiv/B8gRTISFRcv3C02tLx+yTwIO7wqD
GweJZoyguP1c+qXbG3Qoz0LKQwFBpDtK/PwnLPeaOuzUFbRtk+epKKzRMyHl8S0/OacSGtrGv4Rw
Lo9f90tsO8gW/AtqOkFMNkfVRKOqZ1QqvBKwAOen615EsQ3d4N3g20wy8dxC5NSj5FDcVJnGmjbe
vBjYel35qi6YWV5r12kmnMy4rqwkBPSUuALhxHUCyPZFu1azPNbNXKyGbjNeOD70sJ+l6vCqglUu
+vW0ig80kHCvaBDvnxQyUtGuPtWGj1jCktYiZwfwbnm69PT0jQr9sbd1BhWmen/FB4rzdlEbZVlR
yW3fWXPJMvNsdZFUIwOBD2Ko0n6KXhR126am4p7LYgSDS6jd4xOCfVh37EqG/wDHlxCClC1fCfPa
WcgtK/HE+0j8bxdvCUMm7F127tWcm8jkOCetbOI8skRFWotwc1jEKZDujN8ZNq4ixaDwDVy+ZO4n
q+Sc12N36cfNEgXtQE02TKKKl9P0EcWLvx6zWI+1utVbdPdeV0P1kJa56G1l6emmoLNkpaScxryS
aa0OFF5PblzvjoE62EbMTx54TRVAL8V7cjz+GnfdvTv+9SHRiHztCC0K/qolkVzakSmOfgEtVVDj
BZRyEEDQEgpKZZDsp686HozYpZmdLJ08LkAZmTli/rAfIbxgifXwLnHUu3nv72/QnZyOxZFpdQsr
fRMCyiuxDg52TXoPwarQpR00v7HdF/4aULOJzUJ50OVl1J0NcNI3ibLF2ITgOQ9i55eeaCLZCL4V
4lptawCpRnVxV13UbEiW592JLC6ubuJcYGJg3Zg/C8X4NK+Yp/j4WcvEV0yigOoBSAvoPkYzobl1
0KdjkSPqX9BI7RcisT5lmCBEftRrGZhOOS/l1hW2GjJdeXVqHYQg5nwKtgfXnfzi9Q6cNb6ntNOR
6PUMy6AQKQhExWOC/PPy2oKdXfpIXfKiyvtVKbRT3aMj2dnMulN1VrwIkOT9ppT3GHoyRy8RBExR
hnbSN8mgIVx4Bog32VsCY6b7BauaXd+VYx42mB+oqJbToLnVxKFKtSW6cukpwP0/KwiwulYMqxB5
AgohO0hWQXjLYucg8TQYseJAJ+kpjdWOlniwa1mIO7Ahiz2IQgOfM3lhhzafu2IRCzuRY7ij+rOu
pkTF2u68kBu3RwOyQO8JWUDbF+fDCJOq7e2X9lJNjXTc76dj0WRxdRkVcSZm62g9lrbM1tpAA9q5
gPeoxL/RFZlAjVdZ8f6J3Jd7i5tTquQTX76d+uDIEFg+WA+wPG8Q11PClKLwBdVAe//0CESbIlQ8
6JIrNEqETYa4L2h+/UzM9Q0im0pHpEEbYJXz9ZN2wrsFyroNS/ZMB8jSAuwvO59rqLZSyDSYIF3B
+QnOjYZNeyNRZWEcP8BTwO5agxUXQe7/B6aVeN1uLrUKM2W0lCPtm3tEynkpfj5JjNiW/Me25LPD
SR7aiIMehERVm+ZBAimfDJ/2WCo/lghYl/Lws5aw3/SJ5pAyGMEpRuaoDcVsl70AtpqwBYdzDvwt
ZVtOLUL/HfTrWvl/nOUFwcrMZs/2pm9N7Zlz39lyam2+Jd6pGTdtMKowsnrgyTvD6aIDMdTujgzG
7LM1TPAI05JZu44SNRRQTsQkxkJUE2hWLP9Z8qmeodYabye+4hrRcCjp0gvhYU0aRd7PjGHs2iS2
2fwaLM0EHFgbKETZaq5Gsj6QPcxr+aXy/fF7NmKpco5olLYcSp/qlWho+xGQ94Ac8pP8Mxs/eZon
RShhIAA/4tEsXPsPePcGv1XX57XnbiR2COkMS9XPh/lXgbT6/PwPHkkPki8XThmySiSCzutqUN7t
+5MST9K5ywCDjG4BPPkLJIkV+0WGqPYtiN2ukkS1yZ+YzCFQrmZVn84R0QLgjMHuKOixV7KPHlCM
XnaNq98kCHvpX8cnLaeQ1aue6GKaopihiIoQJRnp+2Z7c0cdEbwZLR4M4e1p7v0vK1dhng+K4KHI
51py1ne7UpZKTr4y96w4eTQAaOwVHesxUvjZrM8qFg2/5s/JWL94TnLOD0SMx3M2DPlQB72/KIBG
Kr+EfFFlUTfXGTOqdcjR8qdReHZW+o1FLAJh9CgQVdTmgHtDiDDiogn+m5oJXhssJXcbYWby7GBQ
zeWGh4X4busq9Su7HdIj4HPwAUAEVecx2O6cz5ofDZHi/LxD1dnOnZoXWQtW+sMWDMxxFlrbzXl1
3s/t/xXVa7oc/2MWJzVfaan/omj9v3LRtFBudlmYKseNLRZublkibjgNld0o5H5LNgaVcDeme2yP
DEut6YVHmx7OSYD+OYfi6V6dG2dMWVVTtpegjW4v3AzmuI6a1rqUFZGgcCQscWxeQSRZW+Va0pK5
s58957Fu8RFKuVIQ8Mtq/ubzwEPdtbTLS5NqrubyKUjhAgf664Vq9J21P7+YYPk2B31d4z39kPr3
ap55uG9eEey5uUNFwZXp0UKMkgRFWcaU/rKtzU3pv46tPrdWpYAec+91mfGOcammdlkEDImrPn6f
8L1cuB0ospVuCcO1Gx8M94RJhQYCKfiONV3WnlKeC0NtYegpWtlP8bh9dzN5rs6a0HSYoDNc6LgV
EDc5m/fa1r/VTRV9K7iJsiqOcgMdb6ALKJdw/WxwOnM/dH4Yt+U7E5rUAxi6VOsbgVL5yzQTTc25
dWiqot5moY6R0HMcQHaOu5N1NAceYoar39gBoAzghg8lELaRJgvQ8LfgeooRW7KkypuGkSJuwZ6Y
9FJUy+bd8J+8kraTCGEDnJkVvk0Yuul7W6Kmof9rZvexz3T17VMt1B8LIDD0eIyoR96c5elTOHYm
RaWiIvoley99T/oyrRaLBVYbQfQ5HV3Qg7A2NW3X7aprlJsWR+xzk9YVpZZCQZlvn/e7PGY14Zab
5C/jsa6n8wDXyeTgSjov3CHZVcfZIL5HqSdiSmLOYOvDFsyu/MaCG3OOZg8LIIbyPuNBYssj0ZZS
csQgYHqS7gi1wEzAwgZliKejBh6T8L8eOZWYNwVWGX6NzXEGy4U5LIJ4/t393kI3wQLaaBxWx5Ii
YyEornox02dYuNaEKd30zBkhBpv1H5672QkdrlWmN+jWi/dqifWYv96HUsnHPWkwE1/yfc5vnAY8
d/pqW4g/csmj0zdGWqqIubCON1QMvfz0nu+NiCX2ifZso0E2TzVd7ulo3ALsbFsros6QPPEZ23Qa
b4USatSeLmtgLO7wtxmmJ9w8m4mEn9l3F6y5t90lIP9nTJTilUsIVhscnnodZEsKKXYPLdykKcAw
StbLS/sgzmZGA1T16IKfqs5RaI0ZMk/QPFCJI7jDCe5QGJTYOJ0k3Hu1scF2XY31xuEc4nfe6S9d
JW74IXz15l4MMb8P6D52ZAzPNfZ1gZEfVw5gYWo4vgp+jnkD3D7nsngTEVR+rIs7hfh9uVGg1wkL
PSRFWqHGCGhlK2go54/kBdTE8jsx3MOTxHRUwVd6wvFCc08ZiGEFcTg07L7nikuLK0of0eoJceyE
WkS9a3C4rh6EvrCEV+VgqD8XL9W8dICuY8TDuOAB7dingUKqkxOeDaVc+tApwmkRq5TbjH2rnrQn
SXTJHbOVi8DqqUJth0B7uyHjpK9Lm4A8I2WevoGJTxQfZ/wrupOCU2Ope9dZeo+nNGmvlzL+OBbe
vJWS4PQQgo3XZx1T0Eo0UquRgCuE6UR9AkTt53LAssXV5QO1s34d/rHc5hTgWyZyTE4LIC0j7ij+
JUKJl6J8EJ5vIdS2wJ+lNIm+r2+pW3v4aTj6QBzmLBnCku1w7WC1TmZz5VXCuZl8nxSN+GC8lMDK
V3baQaY1AQ9rmMsBD4Nwd5VuIXTahSC1FhUuNyhyKx82wpqfQKC+5A5zphj08rNr+bd9wOC3ZTrU
tnPhX2MOHFquuUY2DRCCAIoL9LdL6jhwPD2jisL13FAoqtGN6nMLVtSeN+NY0bB3lnBAnjU22Hc4
WsOh6l2FgafzKG6saGUAOeE5wv3keI6qmzbrU/yNAV/PeS12OR6a4MHZoOM1VFbz1U86UwCeWlfE
JupO7Fyi6WLmyGrj1Nn2sGJ6V5JIF78FFpSdCv10n9LUayt2SD2QQSzNqJkP8S6zo4iLu1ItC4CR
ewMRLX2VZj13rOa6kMCRYy4cIGt8kDBQv7JZu8w2fwQngD0IrBDcf99uk4+xWPCJDk582e/wGsIv
iiovdYzPccOnBIA70sEsmF4xTbRtV7GmacYYxSObtrclQQQZY8bXHiJfunbPIUUsdvJQW5bJmrZJ
1tF7Ml64NFDSag4jE6q63AM/cHbTffAjee310AouYQaTK6BxUF9rjwkNVPSjHl0D9bKoOA1Ugm/P
/VizhHZNBdNS0VWgSE5LAxTdD5vojdHn/fHEg+IEYpK1AT7U8gIxCcUOGkvxXe0fZyd0hCx0lIT3
nrXGm7UIahtfMvTLUjKklczIJ3g9aKi25bDisStUYxXgcH+IRo7xyDeRy/HpsZWHilU9m44VtO1q
VuG2w6Y3FN0ndv+cADPAjr81YGKA3qPeQ7TvUHpwzDQuDy4Bq8Pr7HX9Z19qInd2sRkaD0+IoyDR
4sKgDavcK068E6DmjXm0OEyWjWhv5bhv1W3JUvOL19fgN9je8x8PhdP/WGLXfsmV4uB0hBgW6oqQ
u9EsFUDaDW3Q5qSXYZkYJ9oypfzy5KlIDPi1ZIolGMMPMT71cabHARFsEXV5FPC5+KRiSwSHpvBS
6syLSsOv4IkEoGM/CetNUOOnKg/qRDArtm6EVzC5L1d/StUj1qqFpOEo0rj7Xl1FwMX6JgGmnmLW
rcl9hsXvdD8wKgiUJr1eJeC9EVmj4JtH7WJo0z7WBrDxOMQF14ijjRVaG2aL6HsrSu5uIGV0P8Ln
lUzvIWOTHwfmhg7F8m5j8MjIoLoAIaVxvPM6Y2n6C/tKUOoKX3GPSUqhstm8avBbEYL2GDYDxb2m
eTXjjXnmws3Qfq35lQ358fGVKfv0/1IUj0Ja+5J2x7YCtQ24vbXcU/8fug4YkbOpYjvxgdL6GnNL
VRGm/QyhxY7gVZFNKfyTXFs+M4ngmO5HBkKIhaT6eLH4WSRt95mgwPVFn7qmye+5JFC93f6nO0uC
QoMty9r9OnTSumNPvfQJd+R5xpC1ucZWB08+00B58ybwo/DOUmMC5Y97HORu1ltIT++SD+fwySF4
tFx//Q72DmRAsPI4UAgKs337AqY0f4Q+2wD83Ss0DKR2xdJSOF2ty/wnkkbRRuk+hlR04C6GEBZA
y1JMCDjk8YXXmKo+i6B4fxSL7nn4mPYSYPZadgBYSFpV+KW2ZZqNTwonQa7ja5JaqmYBr7SRrg2r
TlyfCA6tml1L2nqmdzJY90wyjkZ7OLnG86WtUvTPT2CB1PBH3EyD/008riRbkBmQTSnBrqNgWYq7
tzk/QlBgkw/fXuzYvqbK2oZWhmouKp2hT6voKavqUwCbXs1Pe/0gln1oTvai65B20rx0eGm6FIRx
kl6DB9K3i/wXzFjlLi5idRMTzHWmsoJfC7w+DSVxXc5aQ8mueYc7A9WZjTaazlasRiV4F5Gv/iUx
FZAcXkp9fS5kS44uRxXNBxiM+2akWSCR1dF/2BVbXcltr2Yfij6TzdvIaqqay9YbmyeIk0MuQWz5
T40foYyZgkzJFlS0v16v4o4WPIH1xuAIpuARrjrNM9WlRY+RAgAkQ/0ffLUw3qlukZITz5ssjaiK
DgHwxwBhu1A19ROyXut+U1GY0cpRcYqfLPfcjQOLW5//PBNwBtjnrRViuyIzq62G3mNdG5vpCHlg
nG6kbsee3VC4sfmoAJip/q4nh0W8Eo26NSZzzO2WnH4Xs9la1L2S+48Ll+zj5dQaxZUXV2dhHeHp
QiadjVI9iiR2agthKB1tNQ2ef7zuhp8BU0Dxjy7LB1sNcnIsypqicZLVE/f/jExlUUkAvn1iD3QJ
7jv4rOLZNc5lEID5m+PEgOvl/7+fPOfVF+cqnkAGD/r65SHwaUH1FqFpPJR0OY5DDXGUm+/7TMPx
30Vi3MHSgzVsDjvamXL33tpuNjJR5NBqIRih8+B0wcqPOLVCWIY1NYaJhYCDVwRtin357fEt1Ew/
T5nyELoklq7agYaCPJlfUwqmRMEjcPHrie26h5H8q4RiNEvnigPMSnLrCGQeWWCv/bnZ+08NlY1V
tRM/0/6/I09aO1NpzLJt7gF8WAiwqQsiYGxprRHSaYwcoflcgtEWyL+qQ9rN3Ud6i/9jKIOfC9Ab
3jqacukYHx9OxvMinu064VTOCYDKawzoOiZZ0lMfREefqFRJQMSmDWYo8YQLmJcV2ueBlWSYTjla
1eymWvHR/DsiBW/W1XW36PIqowjvkoXOw/HC3R6bvs68u9EhsNTqQQuhgNOqzD3mosr6Idgw8w+W
BHASTj05cvgdTnBaCuxSxm5oVrGr9fMN7Uu5oRlzxKyFVFn0qyxwOLX2FukoNpW0o3eE9iVHkkKO
o4zq6fjCvPryoBEdVuVfYdMT3Ufl2wtjbjzliC4dWZ0PJXFK6XYaNJMyzEFtQVSc+UJSAx66RtJI
g8tel6OHqjqLfMQOdrxY2oCE0ymibh7SajNYh6kML8J89TCeVGl+0vl/ejaMQw9VpEtU+gEXxkwf
ppjq17KGdNwkji5b3uvRMOTlDy4+9cQB95SSjH+G7Izo1AeJ24sDKvF1wNZkw0yUVvGZkbFWQVX9
B69+NIHoGvzQMqceP1o3IOpXkGFmOsgd7oi5jQDVmiSzdC/+AggkdhYIblD5hAzAA3/4pk4gJIY6
syqNj7EHoEMTD5qGKESWOK/XzRZv/PHM4l8S4oLCnL0wMU1CKSquLC4R27JHlMVeFx2wkk+KXyin
ZGxJg7fwOEVQygSdNujHLo1a+ZbBnW2K/2AM79T+XorCpaimr3WLF3xxD+HdcZ9DAYfRMxXszTC/
e6BM4Mws+f1gF/8pe89Y05oZ7s9xNSUSbe5SwnMvTKZOEro/tjvHi9U7rIqGxZlmWROTl6cOqR3w
O6vXy1smkeZPleNYlqmUfYh5pni9rSKm6U4t8pDdzya+HoyhcGftuzGayVhdCm84brhSvgxaVwxn
7EZoOrnzbFH6WZoEPqjjLJBstaAi4MDPaJpuTNStfQhEF9ZX0y5mkoGD7I9Ie5YcN2g19lXsnjAJ
Jp0Hoaoe3zjethzftrMFxqR4snUCOTCwJoIwh9cStzlS0OfXRntyx83WA9X6tDGHsZv3mQmPn05z
rlJweSjQQgy6cfkE1fa/1OlMDifa4/D7+J8cA49k69m3HpouuZvgKYabc9x2oOPoETneWWZW8rJs
8oDz5JrnA40YltQ1l71uo/ywKM9x0jbfCdid1A677Z3Onv/r/Oo+0BlOCugU0WEpl8aS36EGffMz
gsXLT6xS0aKtkcf86Lx5KAJpfEFnzlnIL/4llVZr9vDHrXyW39lSkjC0aOQoRy4g0NJdIF+6Lj/5
vfC/mKZzoCumcL0jN0kx47tuY4pk2OyWaGjqsxLPl/197/D+fjElWu0IAvD7kmslTZfDYN5J/6g+
bsiYQxumoqbYY+wV73UnIEhabb1m60Q3GsUykIb7WcnYOurlSxk7FSKke+Y86wHSpR4KHLj2xLso
8/2pn0lBB+EeuQ3o26n/XpBUxH5Qi1Q42O16Ij6B2h5mLi0wJTiKmOXU3xv0Pl7uovQKG6hfSvHd
njDwhsC8SPerH3ia6mT2y5dzcbL50fuVwJmClZ/C5ixz0HJ+YaJakc4O+Wu/086H0KGk8pxi4RuH
0CaSjLFVT53/yeN+kEPb96pFFX6sUgrNTAGCc/I/oF0juRTHLVV6TExYta1IdQcJuVFuLEqMwHjK
mWfLpPqTegczEozgGAwDo1/15gwlE1evb+R7KRoKOvEZWAHbqL5a1WkjSSjMknbaJREm4Ku2/S5U
9jYozhwm1v3x0lFxRj+nbs7VF3l25QB0XnX/vs/0UrOm/wUskue0WEo3Ub2F3qZMPjmhPRu7xmzz
55MwD66XNNKS5snp/qsxNDFAJ0POGMwBUBNqwzKPRa0oc4hS3rmMmCzWcv2VGy4J8jRhTCdzmo9S
EECPp5TPg+THopn3f6QqDQTkmuEMmGcIucz719GusGBiVsUwRlImMgYsb7H4cnITfe6ei6I4gHvv
dFkcDFeVR2YAiYrKsM62trILbfXjVGWY/Qy33oeUO7En5snaq71s35Y0tbNTsnV6v9SZo92gYIZJ
uApMd+qa+BOsOa5eKiBEMKqdKqqI86fTqTcGVi2n9kJGTW4ctz5h9uXEWCdw0IYHJOFbXuclaogr
5dvcnUkCPmzcNp9w3j5/zvvGp9jnptVHkE89EfHAfChI3AB+A1op+o8gyj9wtQDI/9C2ytirIqp6
e7pJl9zfZOIj7UlLpQHlam92Ch+NY8zq/t86f2+bJzsGhUwI7i1gjdJiipgHjYes7vpNfU7pj3D9
2P47lhj5/Au2mqIbvlNd+kdCJBwOCQyDj43kLf+d6iMVO9p/xOPOVxm+DrEacRfuIWsQ0BK8Ko2/
Fmo21reNZC8EdracoZIvna0XYAuF0x6/gLIvq2btmJ4Em98dVknVcDJ7f/mxQCjoXld15m0KWnMN
HTMftdnAHhpY+mkL+rqWm1VDDDFN3pdwI5dU5UtRveMljkDSPegxb7Cer2e3E747oqmaXErkPSig
0Z1c0n8/9ZSankDI7/1VA/sxcVHVQWug84BJiYRT8dTyktzlkU9cnvY//BNcwr4QpCnBLi4ZG83V
LHT1oc9knRyrqYsVgNk4BakAbUJGgOHBp9oy5nQXA+gF2D2SIj8tB4EqFbgFaPw2wJkhJGzaGMWv
xYU45WR8v5igcvPx3LxcW1CzQ2tWlklS7ywSPIyJPMe3v1rZMkkEN1wlXZ4M8XlYROkssF3lgwIa
UtdnFVx4OEt+MDlqEm1zidBko4OysSFKoGfs3mKZzTO2sDKpA1/UnAdbhAPAazU1EQwLprwzZi/F
egUIvaX6Z2yB2xBOGKL5PXb3op2hsxhG7a2aYn9NMK0+au0Yt5tNobDzQUufbpOVksMM4fnOMLu+
RlEDL+sAEU9r4LTSNdFzWNElFQ4+J8c64D8NJs/oPtMQwRVLjxO6YmP+0igX2uuqViMafs5jx4hp
LfDC1VirQh7e1TN9ZHxcZ85jgEWzXclGzX4t5n//8lQxVzkxSoNHd3b3PRaqbpFgkTdMP5GgJ+5t
BMwPmyyLOqAKEKVKit5altWCSLYDUXQio9e7zeeQJ+Z4jwUL/OD2Soo93a2M0kzSZjrHpq798864
JJl7r7+m8A/Py/BBwuMlVWbk5uvZYJWY1c++BYidVZRViAi+SRuofvxtbyALMj/8V9rIIIqh3KPn
KajBrWRZo35rlbq9D5UQ2wqWxgUNhtBig88S4uuCocyi6KWAuGnOvHFhP0VP8SeJigwwJIelEGkD
G0NVFJbZajiEEPN8A0FGeSpgqYijllKlTw2api6vjGcz8y8qQPsshl1oEl1V8ks+9EUiNClC/mIx
5hAIry0QuucRRB0HKPR4AuixtN9Vapp0H8LZzk2fvYtXQlpQKpeMbjedJiewk5f7UvTPZTuqzYl+
dukW60KAg2Toz1t2a5F6zidK4jnY1JltPSaCi4J3tXnKxeHGtQYaYGVuWkWyCZyu4Ye9DX+lIbT+
fep0Oezvh4jGAbhdETV8oAjiH8K1fE2dFLQi/NF8xd4g7Jb1etZ6XtbnE4k4esBJR5sgharEDx7s
YHIIRoJYvDbnCASSXpFUT2/ByhGoIY+DUsjp7oP4ztXJjVbEBrgMqnqs93dY0e/5lTvLLQrqMRJu
id0IYWCHx5XIm6Pi6Izy3b+Lyw9MYwUm6VcNBpmM2SbYyGNQyNlyZGxgfupJgSOEvy7SgQB5d8Qk
fbT7eHu4UfA2JvD+Yx8CpI/Tue6xjRd62uGL2GxOCfQ1h6J6Aeuvdj0PHf/DNew56BtPQ4X3lGRn
sEs5rqZrgj9GvXE0zs6L9yax+4HBG85/26Gao/bGEzxqTpfGBai0m538t8DSx92I8eJg4E9HcIXo
eT92rnGfNqqa/o0DYPOhwF7MdisYNfVPTJdzF24UY3ObcPYAE+oeU4KDeg4J+ELbjAzWJ85xTFGx
l6rNeG7wFqc6LKwxQKV84tBFNP0KLtIKz2neOAtAUtg8iPU4J2jGEuOZq+NShgohqPsUvxNubTiI
jbHkmLoAt26+5aNlqQM/H/vv3B0BKhgigYmlhNkUAh9Nf446W4FfzQd8oBbh5qowTUl3TOjdlvny
uJn/45aGe++P08noM5fdNwqol5DI8+JFKGD4ZOlalRIsw1iD21GGHAgv0SS2IznXG7EYiAQRWhll
wREKYLJX7J+1lzYiHBHkhL/bX/gtS09aLmUo/9fzlV4EQQBG3wu7gRm8jxHVMQLIOwxe8CX2i01U
S+s9Bastkha3h+74D2tNkydPIPDWd8hfu9kkrtAa72FpjomdI91bt5NEdPX8KyP4k+6y8nste/3K
i8Z0DcF1q8Q8GPNyH1L3lNamAxldLWshGQWddhV0SOFXykSYMBwD7EMQZzsAG+FOzraxifwRRnHL
+EWdhT/DiJ+oK09dcVnmmJ9f8uD6r6bWXFhjx5Bt10oojHVMrUcNysNTYBUC0HyGE13z+wM99kEv
m7G+S6vzC1GoWaL0r1k0lj65aZNieC2BtMJzGzvKZIhfa1E2WtMw5z2oqhsmplCXpbuQC/kcMRwE
7/dQuQyQEfiCww/AfA6jkHG9Uy0soPH9Ck7x2B65m6frRFkGJDT1omVrZLG1zU70gOHlG8k+FNjb
+rqoeVWu7tC15pfg/vVG58GQ7Sncbzpd7SVOMgx4KGtBjGMs3kQFx27/xMjP8lErwrxoxH76nyn5
m8KWFW1bkiPKHeaftu2iRo4I0r5frdxVUQWdyVDSfcewuT4xCwKq01thY3xjsHGjOuYB9vtjJY3q
30MyFk2u4ArsJi5ir4Sp28Y/1ciEO9FKpkN+pn42OybJnsqjQzSWIks0i7oocsHuBrkDJupfrb9o
UotxORYOLKTWvBEQvhwrbXUTRsj1T3h/3Yr+YQ+wdYKijEA7jeefsK5ERv3xUlQRB1gTSUR0UFCG
KlV78Z6HUhAUWv5Sb3n+ovvpQ4YttmU6KFY0bLe40MSieKlBmsNw2xal/Uvu2h6hKXHKtMdGD6MR
sEa2+LtnWwLl6zYE771qufmupft3IdJ6H+v1MN5Fg1ajnRBHKPycpkm1+zyCtq4qXE4ZYJv16Aoa
KahwTyu6a99G/FG2LCbLVq5cKQHmxjTtw5DeEpQ2XP+vrW4GfyLqoxC1j8Ixz6v5co8JaLjlifLu
ufppLrRjALhyNaNvm3W5ghk9sZI8I2QCZSOTQvCi9UpGK9Rpfdnr9Ewiyr0/eDCXbhiw1gw4j0Kt
KXcNe7DMYMkHYs1sSFMegEUoXIPZU5gZpqEkSthjAk0V7MQvCzcePbn6WHcCiKfovYGuWnZzMB3a
qpHcs/Fw1VDXODGQk7qeJfQv0bDFaYZHgarte8TRwU7d6tsfNG7RVjSnPq/cxOg5eYZebE6j9Q8+
sp+d0xgh28UBca71BtygC8hhvM6PzTKSzC184t5fGOekc9D5Z76FuIKaQe90oQBeDcuET3CFWUdQ
4FDksLQtKuF5T938T/ZiLuInwaXdoewFFdZCXjYwujQzPJbZaf9arOK3UoQN4wMwHfb5C3ATtnO/
Qdx1ZZrwNyOQRc87PlO8VC7zCWXiAQAF4KQluHOQr97Rw0IvXtBUmJXvbQzogXRPgnjM1pP0OSBs
YsJ/O6W4Uo3cJ/19foeoxbHtwJkum5hGUoX4Hxx6Ma4rNIarU/AWQuDtE85BIg1z0dkh/vg2boJx
1fXxB27ozLuJ6cXGBstg77GULk/VaCLGs6yuRQ3epsBDH4q6Hl/lHdouxJGIxcLysYWsdCsacHFw
BV7/78PaMhkVj4d9RXQu59PnQIgGIoh+xI/QV0N0Js+KCMBomcmW3lcRyYkV59al5bdXDuizyasO
fbGYV0cDdRPA4TH0mNJS+5bvtriZuTGZoN06Ah0Kzlob8XJooMIEBY6jfooCR12wGvNhqn/MS0Qk
Z0yGQux1xD9xv0IIlC8MZTumti0TRInoFruiP3RKYbWRi8VIDJawEZ0kvEYg9zNgq3snfK5GgefF
dxhztKCjFKM8iLTtpzlyfbYJRXI2bx3UveAHAO4H3fLYNFDwFk4DjuVOd5nDrkHm6j3Wy2KpwV2Q
d7d90ggg28PcO6oVfTbrI26rF+MUfxt+i6Ofu3y3WCtwNUtetdbJdXY3GmYvYUImqy/5LGCWP8R0
qazfn+Oaat9r/Tytdjny6vNgKiWBnqBrIiVeYTLvLt4Hqlc3xsUibhdL35EtO76Y1CG6I6HkKgl1
FEXKfDqYkT9gCjSFcTiks1Ik5WTlmeM+tD0y0zdpQIg+xx5BdIS813aX79VQR8eiq+tF00suJP8x
pH3+JtmcuIWd7i9dqOzntxi02d1p6O2F5TEi7pjID8QoTICJHkhAD+ZO304s8kcRALS+jgxFwFqy
Q0oc+1gbe54yJ3mWTJguzPGYeuhnh+5mh1S4DSY0rRqBqPJc/7IwGdQ5d46ANIMj/9qbhwVgswsg
a2e5raf+GzZ2aM4OebjkTryRfcoX8lThPfFGZ6jaWEB+xcETFQWtRC4UxVRKulSZsIvXx29n0Fcz
hoYYF1GzuWffF4AsRQpOjoVdxIX+TXhJA5sMtTyw2uKiBxnaOKVpxaEpyvTcC0Y7TU7P5LF2sQXr
1tu0PfPaiVKHiN0w7xmj1eCWCCgDTfo3p7AXqFoXQKKCir7IQhwkynCZ5kvybXMJgbD8OxMW4UnD
W/yYEDoAI0HTFTcWZ16F5oWkzf89Clb53b94Pjlhw8wsrsc0IhVRwczm1gRM5/Ds4C5o3D/keGOT
WEhyf3pH13bybzq3E+xcCoCyJtD+Z20SlwxeTfUwT/Krx+HcvtDFWkM8UOfMxv36YQaQrf+odB1S
0Cec56pKOxbr3eUR4SnQl+OB5Q+hmidiNXVVJU7ik6FUVb/WnshgOvvOdb8+IY/AUv8nx2CPHTmM
GmpB2OS5t5d9ywgLzJQdSxLIqUHAKBXKpjW2vlxv5OU0koU65bQCcOGSPtiN88C1J6whuf1uH5ib
t9uvvc7WG/HCFAubTvIt/qoVSZ6UhLhNbsKrPoRiynKUa6ZGBq06ttXDNOYHhNe79c4QaKlOnQWb
OIC7+Ps5o+7/zWf3NSpBWvbV6SQOYzaI2pJGrF6y8uts4skwxklNW4/cLSRmh3ELKnw0IuJx6OId
GROvgcvn1tmhbuAYShBO8XCTyvGiTlzrb73Y62QrUEWqDB8KF2n0evN6z9GAj3kH49r4T7ZpjqRr
uU2b6Vaua1jiyfB1j/C10cOUvyFjmEvtrX0AO/mUvrbww1HRPHiTzTJ+9AbrFcYwLSl3oWfwdUlt
elmPmJu9BbG8O7RspZQXoigTPlIySq1uF6gd6dykGnpbjJ13XznGDeQFTxcOg6sUqe6ouzpp8MUK
IPR8jIjQnmXk40XkJfXboNEieUfXqcs05oqiVq5/zbNh1iwjyX6+ZLtGMiZjOMqLDsumuda34m5B
r38oqyNWwd3jQVRdkjB94VrJbzM9Y6dd9hYZdj7Gr60JGgAkXEL5L7t4fjWQnlE+ZpJspK/8dfYQ
i++vlP8lw57fvC7IbHQdWSvCNSvicrDzMJg71tFOPJ9pdHnwWdIYvHkiuYFHWygjh0nokeCAfW2U
eugVPrTt0kqcollYvvZcH1KZI/KNnOgip5fW9Ox6kWY6/oJ0gJXzOTgMCxaeqYOxMsMVdb+ttMU4
cGQlcsZ3LGE5slJhTdGy89d8DrHnccLnXxEZeKOSAVJyJQqu0i80qbIj4EFN3/rjfFYkSxDbBznS
QBj/Aw/b9UpgMIq1owPdJ6l5zchsfA8FOEFZ+2/gmtVtlR4Vdy1C50KPFqC5PcyWi1esom2Fp76Y
z+tUni24R0KBH+hqDplR78Cbo8qYrltRPoUd639HfIP6wom9bh3LJzatdXHOPaTuTi8hqKkAp9F9
bP+7YI/fvM0ojnh8ajzA745PyOiuyn5kJbCe9pqkr2T/61Ec28fH4932dZ9jc2JnNopvdg1P5k5m
3Hw62qlRiys+ED70hgKt9n0CVlMTK6owpRvOF6lvmfsrNX31Q+4j5mxU61tP6kszv2yIU45Fw+TJ
yCMXI/6i0nbXC0a1TVR7ipMKlCdZJoLc8RkDLCKYnEjgyV2aUyB8dO9Un1pnD8lIJcPUzb+xvJVw
lcbQarkwWUCKEBcKC9hpaGriZfYIKRmkJvKuIE0mLVHM9foNY8mNs6PppUUZ78i3hQil7n0Azp5e
4F9i/QzFpHQeDgtdFzn5tLbUT59BmDqb5n0ctO3Qi3b2nB95whj5mM6JIqHw2zh45mD2dflZgZSx
UZoEpUCrP3AYNa2R1J+q8txqiDi3g+QPA/FRGTSVdlex7GL5brTI6Hdo0M5zHDU5ebSNoKsbQ7Is
wDkvgkp41sfWw5LqMkdllPrDaBji0PhOHtD3oP1pXr35oXbRIaQLD9vIUhJQsODQRua+ed7inF2u
UdObOcf5vllwuSVSt10Nk7jFIpNCwYNBMLEMxF6facBm0C18KuCVjdrA8pdEf4x/PJ0rmwU7Lb+Q
iAPbkOgsRnwUr5I0Jb0JfCGrlfmyhg4Bfw3jgFFTTxwyktH6axttVgv9qXjOnCXoc3qPp8oo52PM
8v+RFbg6p0joYV/Vz8yHfUYEKLw05gcB/Z8kJenvtVFEMH2nhUWD5u3LuNLMREGKOf9g/zoCV8ds
Lkgt6jHyGhSI5Xif+IOB+6MQpt62waqYsRMdWmj5K/Q9Bpult68h84GuI6rnwcRa5zNxw1A80U+6
PnZk59/c4GsFW72GDqe4gPliISF7zAxy6Oy84DGk0AbYQIJSQNNCMtKZVmDkS63QJ5dbXKO8w47j
fBP8TjzjuYOdVxz6+umztsSB3pFDWeNeweSJtWMIgBx5LMTrVwtcpnB6oIffHIUNiUdkHT+jISCb
AmUmfn+/JI/NfxeMkmV/HOXsVlFU9cWIybkDDckgczR0INLGJ4BLpyDT1SPJ4JnKoEHqZWb/yX85
bJ6QUMGhSBWu21xUINFfZXV98FG0S9iQRNmyhd2Ib+yl+CsWlpX49et8giG+ylbXmTgdIKxO0k/+
Zq3EhFLHv/mb5hbQJUj996N+3JM77BLnohsmzLRAKOuDLXiqWAnMcvWDT852QvXZO72Lebhm16Ss
6E/tMTtG/C7+JfqjQjt2djBZA996M4TohgheEnHx26uiNVKz2B02H4sco7ENAzhXtEGl2bCzBtAa
LW9tOFHxRjHRZRgNelZ5E7NT8iz/wKK6dJEv6Zcydqo4bJuQ5ljhz/3tQ5m4DZnR+HZzlfS5xHNX
zCrUjUAZovp7O0wjFTZZmeCE8tl5aUhugqbnGNXj6qXaAFMLIUIXXmRtW4S9GkXDI3GG9bNH62Ey
bUllDDRcgsx8443rxXyMlpHS6L4YVZmAwhjr4p5cJQwCwkVBiUQbPVKhr8Nvto+RhmdC6wG2EzFx
cCpK15L9Uvw3wz9XMQvi0YalPxJ7wJg9f3jAzEmrljOeXAT5TjuNiobZOloNeJa7Px6clWSl3WkM
4tnoyhnLSN6dnPLl5xDxLrj7yA2IOlgxSNCfrmZpnmxjd0ZVGGcYMc0orlVyOfIFqI99ipU8PkgH
Rbj2K6rbfa4nwZIkxSuAE5qeIliqIud3nO/SsnRlFMO94yuvQs5QK3Q442Z/64pDAKH5E3M2zBL/
Vf8T27MYli6xHru5w1qQRo8RnpByXhYZZfqN8pN1RxfEk0vVj9RphBcL47ZhLQmAEbfvGwpF+WJ/
/ivJBPhD2RdxUwTLOjhibUH08mndFkYeALDgYTw99pKjNRzW67uQsavqVx6cZFQcDjFyuQK4hCMB
fJ18uk8/aZAUKcx79GPz8TnDuyZYrODaqntrVknxMZ/+0rPMBiR65vlOveimlXrAFIA4++eOKAIK
4kQ/DB/M9vS+so8ffhLdeS1JLu6Qn+xKIpHaskyA+AUnX3+FdpMynmLOEz3HaETli5gILUecGxTp
mBkrRaKDWXbCnYI73gkuDHorjqtjCS4W0f8oeTmeyCCnpxkN87lQrN03HgspNMeBMGD3qNLWdILN
GfXYt8yKhGf8p80DaSvGw5FSZa0iYLnKwKnNcc3Ky+F1qa3TQGfnDHKXMJotMB/C7iDbmkXcDakS
pz+mQoFCUC2MTvgjkt+a27A4tkB45dGkNb5E/atriwVtQ9Bq6AoAuh3mKQapKl959Edc2XvsUv16
Vf7LsxRLRR6jeWCIGVm/6sqs7aTypw1OVmKJD3ariZjj0UsKesT+AbdxjhQ0q4MX3duJZzUt2pKc
T2aHMH+NCk7S5awezjYC6aNM2nwDpL4heGP66aHXZ3Xs6gzTrBIoMEzKwFKsZ1bb9vzz5on5qpV4
4tK9toQAx5vWuY8oPFjdFLVw9ePvmAGhVf5HK0Vu4H6ENMVdRYdkzOx2+nNHPScpLpdG+gMQoHvA
ntBHlxs+do7EDvtDXzyIRHvURSZ2dOfeTtfHhgs8dsMm3LMKv9QZsXsuoo4K4u7vwKNDIPesqUQ9
YBok42tFPRfeAjtDc9upXcfaHgGB+OCMAGDw+p5mOot0d3ZRx3bFMDfb2f60xxkbwd3pEDoI9MGn
U/TnIDo7LIKnJDqlL0WytSHSoduUE+8dYxnHD5TxNHJREhqdfqlLuaMDZw43jHMHsLPXxEB7OETD
JEOS9PzD+RrXGth4ahuW7xCGse5WpQ163DUR7m5UEaPNMAai+O9m9/7Ssn5MmaaaoNjvtyLBxpCG
E5jdJvYzRdsU/3aVQsUg/39zoXE1rlQmFIE3HGJUxSXtde0LKn5IBjuGovUdFsSq7juqwaO/sHqD
PAIvJnopldpEQLqoNxqMh2A7W23K9MqUJOTzBrCVaeZq5Vik1uxjA8e9QRGrtvZfIJ/8OAmx8YQl
QxWaBhKxzJlV/CcpsC+6lHSaBTW/dhOPrLuEUGf2ugZrK5iAa2S19pVkYMQYzesx2dWm6G9EkQRZ
b5QtOKseVhoqHywYFxdiE5Nd24I7F+iDRKXnQv6DnSlqZcrsfy4JVpNLb+s4QvwzZkPWqBc2DIaz
TcdzAM0pe8z5ZlIhR4cZ2xMGKtx6JED5ThO3PzPKujYbTZAVnCDfbC7vGJJefgHVp55HT/Yaithi
+iJLJlUNzRxH+6upO5H6Ef75poAJN/2arzHMHM6O3GJ2dpQkNRrp9g/ge3KYjXn5uY3wh+/d3Syv
+lPxTHS0wq+c9xh2T3nr1I9nSfvVu0lp6UyiwoO2h7pt/z+syh2zkvbRo/fDD0w9VeLjXq2ia4nm
luOorjVaQUYM+lL1uD4zIS8DWLseQ7XWR8KAEifwbt1asNak4egXpwrHv8XnRcujb1wfBORveYRh
8byQp4MePTurUSxojnAqVugrBIhNEj23XsBsF93VzEG9c3YbqC2Zt/K+pG/M0j+kdj8UlvPzBRyQ
4XJrlq1Y53FaKmLG7INtTtl+qq8Wr57zruGWJdITzwNBA4tFJAITpyGrplCHfjkC7gdmZJ7UbKga
M9Efwv9Y0F4l/I+uRKDM94b8wwJLwkkmZrXrYT6XjqrwHomXZ6VBsm12KvplL6oiPdq827lgvrjm
33jL9EwhPK9n6tjttyMNKDtes0LLK5liF4NIyvhAAxLtBi8fEK8FmvttRk9CU+KMtlouX3nD80oX
wvparU4+xWQE6r57GdTF/uvuxz6+AWuLFBI9LHm8m4Vxe0rQH4gRamuMy85L2gbrtrNj8g4aTb4h
Rdrns6MuUKuCIrVU+de1UKBJwaHkpUo/ECs3fJwm1iE9BGLVd6ogRkGmfS2MgT8u8TpkWLKQhoVV
0/kJaVfdFLRf3OvRrSCVwzySdIdBsIQlhKsxOMmfzqbSRKx32kXKTjy7FUSyljGP8HO01MWOA0Wt
4IkMCnpep+scFinj3tJ/FE5zCcFzx+aNxFuRMqIz5l2JfP8DWR7pAT2RX0AP59MOHpq4iPJ0yOsR
pRO7wdC6bsvj5L3S9XMj3292f75v67F253bH/qH1lQ6VRMysTWLrgwICVte3U5eN/iuVNjOpW80c
VXx/7cwroZUsQGZqjcIz95o57B5VH6N2KrJlt2Hr+mHzHzErdN3hF6SelkfNYrkg34Qr/q2nvbA+
APuCPKny8xsEUy/DM01arScr6dUHbxFP7opFLq8VLHIy5dXPMdUVlrMhtJKmrNAHjc7+NdOjsJ+S
B6czRj4Lrr/NHJy2Y1d7id/98xWADcJPrCbqaHs0qG171ndAjBqdSknZhLB4oqQDBMMNMVmVwAmF
YRbIEC5/4llDtI/ImpiIBJcHLJ41cydDCrtNfsp0bKV1AWD4bFfFvLT/qKCed8AL4Lq2Wvpis6MB
w+ULvNOePajJ0sTrON0gtcLXKGM/E9vPixDisCjgQnJGXssghmi1UP6Eb1aWru+2Bj9y9vFmPzat
7XM6gij/bOeOQ21onO6PFj5gkPbNgVRIp6mv5c7cQjE4zwL2vhWnu1x8qqtkV05wm79764orMzX8
YcuRZJhjzpw+elrqBUWLv/zOm08O4FIMvRKEA9vw6nGIskF/wLmo1nGz89HRS8pu9txdz40i28Wu
MFj7UbxKw5GUrsx5bx+B4aJMm9xCPTFhbuuWg8um44RriAkRUPpgScKQb45A//irPfht6XH+IoSC
Y9ymrxNHIDtY1AyjuUwJzk6mwgecDqAE2V8yG+lbN1xO2bx5szl30mgHBm6cly9w/CIj+0rh5dCK
0F+ETN6LzzeX1hNerBNQ0UY2nyevMEGeyLp353//ExTtMf1HCjTVF34y3i/Xxbhy/BSUv7jfTijh
hIeMHT/s2aRKLfc1aYqTtNeFe1gTw8SZVqZXRNS49yHvAOZOO7/UMCH+v+L7AL9l73oHjyXBsefX
rqug0+WMR0Sm/EUiZ/LFSXNlvmum/eB+JHB60MZXPu/IKijbwEdM03jy2TzTUHPML6gsFWugtcTf
uf8Rv8WPWYkFfUGB/q52Yqmr4Sy3iXnhYfJazxajtYLNsVR1uUb8jcb4zSV9SrV5BeWVMDT2wnad
pdyzAohP/RaSf2XcF69VDfvyCAFcPPBApaqacONMQYtNFvEoatfyb6YCDO5EPcOeRsOmRGYHbfLV
QMh3IMhjBLqTcMhhNR4yDm48sEjzeKL6y1y/4Fm7BMx6PAdnngppZjWyzTebW7RFYiwxlUaf/eaK
DZk4k/oPksZZZN0YR0WYh/Qms4xIKt26tse0AyGOrIDyXiSnjbhgkT0ONL1/86+AaulgSSgHKIhE
WAb9UnE/lvIZdCZYyOZo8wc72jLZLXxo9vM48C/1FYEeeApUgGQnCFEf6T4BrfQg2dzFD4Ud4oR7
SXYLF6cvRvymSlnoUQGvX3Pbhxcdku3FZmZvBCra+KpP9irVEOtFnfGpdR7r8bSlAfUsbtj/kt3r
iw7icqTqDAvrcTU4+DpvGulQIeTjSkkY54x5UjbjlUca3MoAoLVbUVs3EdWc0mmC9bicfaA/eHg9
dZe0BJLr3o+4fu9ETaQ58DMuxw2r8AJq2wYiPORQgVROnKgxhtk6P7Bwttru5a1Lqzne5/XyqyHU
Tplts5xSkmCKoe44XfmOzXX900OSlJc+Akxh4zDf72CYS1VCeddhHVhxymCltZ/J0bZ0yXev8dwX
q3Lx7sG4j3vn2VkeMfpYn4KHP9H0XLdsMC5SBOXEXn9jncYvZK5ZnuW/aoU7kwMJoMQIUDZHbCIp
n1eOZ/psmfacAtuk48CFv/p5UE5NhL4CZ81SQDZzYtEfZQLXIfzHB20dq+g3kKK0bwByY6g1Ia6r
QkgNgr6dErkAQwl33OUYLCgJb2+s4ejGDS8RI4W/q/nm4RpLq4ppDx2arpjWH9+iRb38KSG84ACv
IpmpOPygoUG/X3AikX3o3xvjCV6Rwvc9oxvOr4tQ8Zmp4dPeRP0cthbT3DJoMnfzTg71QoXeYVb3
9OHgJ3tVUCgMuG8sPlKPHmVljsO3WK7wGLkdWFeSwtLRtm25X3Q4l6VsR4sguGQa+En31btbMqjb
74vg4uDP8gbEzC5S/qtiJ9TMh0XCsiFr3sZI4lXlaUSc2EaKGrAQ+3i4oIVgICcCvADyuthS82yp
i7Pzn7MZM+sdL6ZxV9oWtqbILm0jHKNs5CCJQqOuvOK41W8mdL67iQOUqz8oM6f9Xd3GzvON9gi9
hQ5arwJPwtcAQoNRil/cKo6cVlByd0lh4djwi6TFoXKegXL021eGkDXydxCfvlTn+qGvC3DNqct9
NjXu6qbRCSATPYAGnNfhSS/fSduwGdsCBHR+Nfq6jbTZZxd1mYgvoMnp0kFYnIOSTuwdfT7FGkVQ
7ojL71ocMOWeZBalQwHG3geg9rnEtjzEFY873I8CvlOZokldWCsNqTIrs5KhZ97S0xw24p+/D5V/
P+x82kNWllXGZXE4SnO88Q+EodPJ5WKOESVG+HbRyPLkDNraGghGM+y1MYJ/6bW7RQv0l7jJAJqR
6KChs90A6W6/k0LXtljsETotRcv7/fBgSIaGDoMfHfOlcOJNNS6yW/welZcdDvrYOGT1rmkHBl/8
Wd6p+SdNBXN+9SMCnlvhuPSiKqnqHVjbESnu/gABMq/Mfjf5Rj7kdgbtjmmWZbnDz2sJqBbmOhu8
jHTSE0gYYZYOQxBy+MruD32RYNME06a25z+WlcExnjg2POrhgiCgs05WiE9Ysbv7eSkVwX6eIUp5
ulrrH0X9n5z50BK970pMbKiKyxRWIjVFMbioFtJNWUiT/AFI4QkmsdZ0/Lhu8OKWO3R+iw88WhtU
r10wGFxVv7vJApCsCMi0Qg4LrFKqqWpdktdQe4pkGeEnlKtJHrYz8/Fruhtk/hwn97TyDk7R2/X8
EAn+WRC4BNoGfYUEZgcEhyEKuzJvEP+ivSe/JJDBW8ClGZ79KbCnX1ZPu25RYe2HkjzJcziY7Axo
McFGkQ8482V1/7MS6pNng4oD8xqKU+M38QoHpv4kjo7j/hCcw9m65Pqb/rjEJld9iKibY0UBxBv3
rD0qxtwLPHQpMXkKsrenHUHwPPC+PFoy5PTZFzuucjyl3i/P7y3usN7TzzgmSPP8hEaY7lvgNoKJ
FQI/CoBp25a17AYX5UCQlj/JMVazkbb7ThAVvc3L6HHppdSgynIElKuLXMpkN2jiHCRAt16kiC4w
Q2jyY+b8jCEc2DGsItobiNvsDLBiIaVppG8K8YJzumnk+IVC0AzNdvQPaDFfPjz8pNWnLeTT98bC
TTdeDbdxk9LUyQUWPd0IF1DAF34jpfn1CVL579hAs6iWlze720hefCG4T243hEeF+sAhK7vaQZf0
J/kHRAdpgjNuWCItb8ylvoEg1GSFkhhX/CSSGxrDqhFWDDpKIgDaRNie9rYNFBHD6tmEu04OJOo+
W0S9SgeG8/JUg/dWP7mSEvo+DvmlfCYapGfTCzPvfxS7tQeKCGPUOXHgNHjO7CCIXiILVM4j/X7Y
W7o+X623ZkqCFJeuvCQrbpeEOShOP3CZ8l24rPV6yB+McjwPjku8i7oE/urKgvCt2VevdLNoErqf
yjHUjZtF4I2lgimRPOlzN3jFEUa7djQANqL+gQIj/Vrwq5UHo5pOI7Ja3z89ISVEmP2PGeSXVX0F
p4iXO7L0PouvkZuj/oWmp+k+E5ZcvjObvSfUBWiDfz1U/kdHVj5YdV5l1zkaPX/eQq5tC37zICYX
78rF+Q/Uz7y5gUn/owI8c6FW270w5fNvLz560Kw82SKHf/M9uEfaCU4ZqmkDL+VpSNP8B/no6iJF
JbBEA0VA2HosfUogfBIlTb8GD6xDRknOjaA3KPB5Pu2wMGa6vsX7J0nScgXgmvMtp1n3HrUUdeCT
kTlehyrEAJq0kE4QJ+AhP5Eyv8j2wrwOeo+lqYTdHrH1wL7Z0DP3pva85Yb8TFoAt/8YZ4SpTa85
xvrps8DeyNZf2Jm/9G9+6BSVhdmDORlLvUdbjtdDRvRcc8a+ajnhOtdnSZMhMjetUh2Dv1Q4klpU
nxJwoezW41hjsptGBTwxR9McbuPO7YGEX1I4mOefw18mLIkcr/4I4YQrZvFIpU3qIjJt6CM8yn/l
rpszWlXNVj4cAXOhQnIHPgHwFAzXNKXVS1udBqy4/ED8pLg8QmG88pUO+FjUxSpbVmGkyFmfyv+r
Jn9v2r0c2EmD9TkQeSYPPh2Vo3FxfP//eZQ72q4eUWMnrgtweD9enwjhv4TtYlO1tlIKfyUBd1qz
eI9GFD3LztMRNVAL+trcAcfE3t6EnvJNfCEs86/dD29lmvO5u5GPgSuaU4GPo9ozKxj1mvYtey2t
Dphw1DjupiOkuI++UyLeLAQ/jx8+woHGK3QHv5U67+/YDoFUBV7c6x8UiSDmiHCi/T78OHdCLTtP
hg3DCsaqcqKgs/n68nyftn9fcMOtIDtA88ZotXYJn/RxzgDkr+MidY/CTajYL0GTUuXSbv1vFvHH
gkNXvF9+qAt6xMTbzknPCeiYUuhSn1zalQRBd7+bO4DeJDkudh4UIisQ43nNE9/cmM1BJBPV28Zg
sIX6I6UEpfFgEeXjhbJc1C7GUEEAQpM0ots47EU+fIFhFaqsd3FbFfbrEXtEKZu60Z5xemPvKSJm
mA1vIvd/RIbo/a64Tz69ovYIi47JrdF4P6M3V4JhhDYLexI8U6pMoDmmJz0GmxX0E48ZqUUa+BGd
088m9TtpGoBfAbuzMOVbTw4hTLX+3pIo6+rgL5DiTPqk+VNGd/qJMndH9YaZJrqdobjHoGubXuQI
r9OqTcMuGD4nA+4JXhh9I0Ah7jqHvYTFQ67LNUdSX3GGcvnMUectyL3bZxHcpDuJHLAXusWRC3/S
vv2VEWzX8KHWL5l5LTwni9ZeraR0jPIKKStjaHey22xOffiOn86hWDccx6wgxM45+HVsunPhqvqb
1aPzZg6XE8SF9vkwzvCw+fymILH572mAQMplGQPopJ8GGwZvRJcfqGgE93qw3PYlX7CAkhf0LSTa
W4J98IlR+Cl2XiAfNoD2IZ1BK3zAcUmsdR8NH7tFAFkD8UU2TXrWlwdDTiO1H32UzhmZYTofaeFC
i4KV9GtWjfEdK8YCpcIJuK0fa4eQKc+JnaaAs7n2hBoEA8SMwyJhGIEVVj0l2O5MpRdINgARBqoZ
oaNHyvwN5VcQVyNyp8ZKSYLgzU74hI2Dnr217MNeB7bVxzeSrbfnWn0GavhOtMfl62f25GuwGIQK
5hNFOGB+sfjKCq1kupUVnmSuTZhkpv0FcN07yrPbhRSDWcw5BP+8xBlfxDPWd3d9G859HilNyHkY
CaEvb1e9eUfqB1LkLZWvnSbZ4nCB5fDaPZW57hVm+QkuXT7rNHOUuaCP167Ye32McyHHL/l5NPHF
OKM5fnKCEWdJLE4LyJbLnDI16MnO6dHxg0GzWGAfUQ5MqNvv4SINTFYoZ64x6a//NDWzvj/lSHcJ
FRB5gU8FGQItlDEtUwuNsyiQvdyCmQx2Y68o5mD/YtV12/8vMaLJljTUO81m0M8UKD+nb6bytn8L
gQefSJz8VQUlbUnkKSfKwvS2PfLHdSivw/YddN9fNcmpesd2hcDRsb5AQUGNQenjv0Lyzdj2HHMg
6sNa2EkaJ9gllQ6ls8T8lNwQDmIqyO2UjwAl4lCcqz3mPegue1IKiMIj5YsxDF80MaeQFv5nBu9y
xe4sCbqObl105qfbRNe07MU8cEFSvpHS3jfm+6Sh0MNXH0sYGC9ngMRpt8vdI4rXwP6+eO6vMfxk
r3HWot28T5vUdo13R9nQzl2NB5biBJmm7kiSK8n93vwlAb9lasNimT4R4aecLsVCggU4EYRI2AxO
7wtL/jZ+zPxgYdeuGmIbHdCEbQ6wVYgdMdEQQ0NbvtkvpZKiwmK7H0582LShhe9E7KwSltMcTvLE
V8FZuWt+L0+ue8TVYIzL22rmZynkQvMuDgn0PtZvTs6a7NhnigtsBiT4lzDN+ztYOModZBehSyIH
yEN+zmPAqu4jq7eqvLLzkWHLdaCCfrF9vtmAtBj+qlQi6luKzg7AZTaWphKqQaaBD9i6Zr8qmfbB
tWdNOu+senNmFU/dkUfAKHDiAB0eRF2eSZpMj1m8TwaqPprTPEsiiMrc+IbHzG0aZtR5JMNCiqNH
UdbVDT/oTCnnYVswt9Jk/Jqk4DvmzmYWgp9Xoz1mUvEzN5wDLWu1/IhDJ1ZQVtmhcD6SpA6ZxH7I
8J2pTGcuOkSO8l+z7+nE78yb7e9Fk0WpGvdOxncZLICnobXrzvNqJLJJ6thOi1hBupr29aVDJ9Kf
1BfzQdYhjXr1UZPNC8NIddivxDhZJ6UFfyFhkp3Cyvx/0ONLl/FvJqP24HT49hwcBpR2C8XpaZ7k
aoNln0kLuQQLDTOjeu8NUJUapZ/osfCH2fUoZ6jNS+/cOLvCgrtPOznJoOvDmLOyR/IM6lVbtolB
9uyTrzcV/+JqV170kMjWKR1efX6lvR/ZJ28kn5YVzVIk1RKdHLuXQ6rKRn3N70dcT7RXiiJ/4wRn
d8Is+1jtC0sGUuUqgSx7Giy8H1p1KLQrpmG9FlR3lQIF7h/1Xpq1ZA2U4NhkKH8UOGxzjv4Tewlf
T11IPZoutKzeMmRsOOHqimnO2VMylC1+sgpTB9HeYY7mi3FymA8xfhsO9oi0VwWAHjR7aU2tGk+E
izHVZyKBsiotg3cZB9fTcygHddQ32/5m2XwPG4/AyncUHGzBswmc2kKSwi3QkJWzKcFHXV7G3VlC
1MBKXQwtKe8yBXc+DYUS/2Q8fJsb/iJoqFwgteb6biPUnX2Jpqg/7KhfaIN+JrATxocxU4+Z6cWZ
kvRTFMlI2TqGSKcnGrTOHZyfFH/tw3M91Z323kuyroIuEve3lt3UoVEo9jptPjQh42/cezscbwMk
2o9co5g8lsujFoCYjLfYLivBl4jEYlzBrEJcXDohUJ1Oyp29KQe96viEYee45sSYakup/3uVB7IL
UEEx2bS6elbJsosFx/qpjMOGeks3xcf9AET9x+uCDUn1wArRFQRfCn/RDQa0BdD8hOK8SLJfeoFK
gkf62yYZxfh1awcRp7Bd7EGNTfUYnO//g/+YClgd8jciRVdVboZVoNIkBK9b7Nhy7AAhpfG5I2jU
gJMIZoAYze26q43ruTCAfYq5m3LLWfJc5d8npI2UCXxR4kV9Wh9OcbZ/1cSKwpn4PP+rAKO11XDO
B9i04O/F+NBCVsA7+1w9aUrzIumDGem2ZP3CUoW25lkUlMCqGuLzbTwyzv7BpDzWjHq+W/ON/MUK
Zp9vNKKjx9t8DzKlsydXJGqj/21+VNZIu9kRVnwdeVV5lgEQ4uG/kwkLai1tZtHEaoKi2QzlbQCw
DUOWV0Tf08cVXUmUB3BbB+1NBFvvD8RbXxZOwOTXA2V+WS/CDN1h5il7LvSzw1SnMjmakOVEOUeS
DD/p5Zp+1bRh+zP9G8MdrboQLguG1zK7YvJ/fS7H7pTUhgyv3NxFOfqXh4S0tfHewHpgR6rIj3L5
LrPtSFXAK5JIlrVudmqIENk6d/X8mIw5fGf1+Zw3gX7nEbCxtZLS6OGblL7WO230WFsWmucpsbh/
GjsPEsAj895Y5gSjQxQ+EIncBK7KR9LfowyK1NZU6lqyhkaZ2ZvRDOX1iuGAaRaRFgipdLrFPuER
N0ZgwRmbQ7c651Hma95aiyaRuDpyLy7LYcBjeGMB6+H3MOV6MpHzruzWVxU1oLEB289KB5qDob0F
NQnvFsAX52hG8KG1giQLZTgwv5Hvxq39aCKgFTAP+yc2ciqx7wwq0Rc02aUv4AhoI2uIXAFsS1ls
JeGfM9Tv8hPxaDQFmTfNQCpJABZ3UhiIZlTxk+TVRk7KPXypvWiMhCrJNdhzn6HHfZ5TRQaip5xg
g9uHR60p2OXpilLF1PLHYRZDR9JL+Ou0hwAsIEUc4eZZ1ejsj8iVy+9U12ozrDCgcQ9AVRbc/QPO
7d37Hwf7B9Fj3te0cXLvhkB0l7ngdQrarin9XnS5cKbhA2V3Avwv/Yi9GpEur9G4vtT0p3zWJ1NY
gxIqp+63CkozXWDFlgZ85vA/lbe3seS+gGYHGhpGbBqezo9XQgznrOUreeMIucfOokZOq5y4qXCx
Z9fIyajUoZTX3dKdvj8e6mZfXxNBbvp869nkuXjKcvN9bg/jNfhltoPDE8DPMVD1voIerKSUyf/m
sNkXvoHwF8klGXC6IEnCq/NsBtItHD4MGEGz9WdsaqAHBqmKxtDE1GjRXCEgUOuo+6K5A20yd1Of
9M8LpxMXKsO66xMe1ZY0UuCP2WOn4/N3oR7Btk/rNx60G7YgUMF3vxwlYgmzCTLGjjfdAHtHtE50
PmMklv1TPYTNiuvgBpEeDe7AT4PMQQdH+rxjhoIO4/zR6usTZH0TPrSez3S2e/6PLQc04QA0jYF6
mWzmixPQvbDVeLhBj2KoX6uKTkdzw689UMdqL20ZZ2e50lv1Ye8H1IipdE/YvjCF8XnOjdwQzBQa
BUR4OQ/GO4q8W7/z57NKYjiDXNhttr3JjGZ6+t70cztQy26RVpXnrQDCOJdCgINhWQGOcjNk37jE
3ueG3K3/r20Zl43Rq/aO9Mg4T7GE2X7zevcVYYxPc6sTSjB+96dtJEcUemFKJgJ5NhTWtutHR+1M
73WP41Z2XfBBm+0gWoD7OEgRaXMClgEGElZGaBXzGm7H5BQF8yVLN/JjtKQ1jJ0bwsnrJdpm9+j+
fjfQRAmN02QTJsjYXBqe8h11+WrbvcsftFw4EiHS8YYq0mbcziNijtz7cgWsJGEzIqR+IheuDKlc
DlfW5vrtWxb9L5/WQiRasccKxpnblg0qTRH92RFb2g9zEdPpCdKf+FYNVV56tFmut/aDBHQKXGIo
kvVQD82cjce9HeyiJRHKjTIqbDn0Q4cvL+lV92Nx4lRZXTExpDci9WwJi04uAVWgg5VLo4Kgom4W
LcAPkES/V2G+JxsgGdoPdAElejhlxF2REdaRm7MdJIAoSYfWFrOxc/iQK5beRiPW5vEfQTSK/hHF
koNCAvb/58DTneIqdE6SWAlOZi/5ttHc4SLXLZ/phWFNhO7aOd/4HozrU0O7NHzjk1+M+boZZ//O
LN6gX/bttyADERMJ1nFxrceKZDD448Dzl1DIA3TSEyyQuRJiOhTh6bxs22kje5M8Qrmj+W82pqzY
h7f5JehiwNEZfT/7twfciFaWmDT38IYLD6ou4ZLG9b+G0YnVeNNqLfUbQPGIGa1nrNg31RmFvGog
dJrDBQ2OAO0YXWer9jj4kK+LLbRYRH/2pY2vjJVgfPNp9SasQGuwa/fQgl3ip3F+DLA2i/GnEfem
+V1dzkUNV7ORqahJFy0jCnfE8HC2do8Gtd+aI42IX2N5mYehVR6QoPbrPLw0QRTGGl+u7k1NyoqG
niEAV45L/6tbEidZ93DkduQ1Ho1nhxyhcHGbCYDLBplkNXIETwI6BR3wJ9ftl7xLJR8WTVVYCkeo
akYDZsl9xfgmrRGTpw+fJh71h6t0e1efgzqDIxgQ4t043N8ytNysOYUnJ4Nt1sMVNEHHkpjvp3HH
/T+Bk1dEdd+q4H1R4iLxPZezcMyLckxebf5T7u79DE3RLtXFj+yKddxzTBW9nu0R0rbdZEtz320Q
UYmz+riwBYxG2mhm2IHaP381BZfHOuhAAzCquQVMX016cHdNrb5ZNlJFIJwaCj4/IVMjbMGlcrWM
4qQ2CMP79ZEW5r+hEGimMrtQOdylwIvnCt/4ckGWdpH+HtZX6X/ZMcGYeMStcbjChQGkUb+FZ88n
wiaEXAREzRwyTakWaKMVjeVdbjY49YOen+kWrEjK+6J3pHOaXaLq3rxYFlqdNpZtukgCuCUR9Dlp
5dKd3k5HoTtzOEIoO0+TxoNR14qs6WD0zjPwfMdclkby1QOqK0ul07xY/vFYbM1WPJwVKaliIybq
2GbFwofvlVqwaKMiWvriuDfdSUpaC3Jp5/bEeynRY7j/+3PyAx3XAUOzVMz4/gHqUBFw41ZrVb3f
ROvee+S2xM0VpdoDvPFtR2mWiPPveZxlFRDQaazmcaevC/amk9gDzEiRjxwrZeVmbPCCi8jOVo0C
bvMWpnUvT5s9/S1+cHGCZPyeLSXMVmikkfVO2X2deCF3QCqgAk312JnfHNoCymZFjQMmVzCh9VgF
/TB7B/qBjBpqAZD1zI9M3l2nUaQtgwEsMW8tps00IJKM71gLEUu0NsJCa1yTIFg6rU1m48zrrT2d
Y9Vcp/uD5vEIT7LaJleksGy1CyZ9BE1ySPB8xLHTY087sZicnwXZphEwaF0PXsl3XdLWphE+bHTx
XWY+554/vNidTB1BYdWdWJ1Ajnyq2LoDOkdbfk9FfJb4gFBQGMGCHfjTViDz0uQpkjmlxE6vNfFh
1789onVOv3imgg/ypRLAhj9Dykg6rzmUMFzUAJGQ92wZkvZroZwUCFHJlGFHd2iOfCUCpiCxeKJZ
OF+Lunx/0QEam9RUs15oe8v0wdPtPziLynwvzBv+DpdOlaMkaiQAtoXdvMrEaMUObDWUlRXtjuFP
xcFYW0/vipqsc3VNdJwbLd17rkj02Wky4mehFPcR84pj8RH/HOuajz8Hbvb/aEQx54VD+AlZdymV
GWM6WEGKZON8oBD88py5bGAfecwORKAVtpvQrQsKorKwoNe4Lf8PAOL5ECaMZpy4wvjbI6Dvc1OU
pEk0hG3gqkKj/RSIBuLhVlnwBMD60JLC2ZcW1wiWcY3O/VHBK+lEkzbUXMFvqSYhRRKhN6Kf92+/
05/tc6F0N/x5n0hJ+Ytz8TpJnq71ER/HMW6e7KEfnegMevXe+0wIa0kTY7kLF/d/OhaHQ4ydK8ca
x0PmHmiWmau1P1HBM7md9Js8TjhYLIJ4nXZrv3JmHzZTEDcD+WygDdRdVrmwZzCv9onEl27yaXQt
biIVzTdLX4ZImuWt4+cgAAI9eWkUwe8mN2Y06YZN7Ur6zBXXxk5JVPcPfv2YM3uF5QbAcOFu0M1s
EF8Wea1qZTOOrQnNE/02V1sHh9hD96lrmrnm3qthhUFSFyVmpXTAZi86i84XSTnfRPpBrvj3ow39
NXYAtkx1b06lvVjj+thQhBD3l5ndGh9Sj+d6LZRd5q+92Vcgj/ZzlQfX+JohUKxn1kG8gJTiH/eT
OfY2uVxespmWz2FnOWYqOR3ETIH3Z4c/fl5KwsbD2QDfX4YCBFJEEUryTk3N679zVs5cUlugrVIm
zoXqNhOrSMThXFJp1SlmlTcqYbsL0SASmGPgn4hzjuGRXK2U3O/ICO3dTjSObpROxUZPBw6N2Bx2
y2ZiV5URPNcPcelphDt4Wn4z84XNZfwHF1CAUGKkKKGZcTGjJXuiSotm72xPG8q4Enz0ozSNsqxI
mKT1r1DZjYtkTRAHjIqsPUUzcSyBHylLUx/ICtgGPnNeMlrlqFA66CKXRCatnc4sxOxGxDgW9DFH
UuiF1OviyRktuiahbEQ3j0MzCS1mcXiNBm95C572Uu34seOYEVGShTXVG99Lm67Ug3YrU+AhCp6h
rj13hUXycIPHM71m/FBBp50ZaClUY02d0VUfmuBd6k2AsHtL2vxPFwc7CG1I5HlRvVPD/bBDiqlI
qTur1Fn/SLGdQ+ZXFCaTJr6XAvZE2vt4/Nt0C4VURSXH6GveCasQPqWi3fYT88X/oL9y9XoplH/n
l+NqnUIUYqGnkjgA7fCSHjIao89Sut+v3xjiwO1bePy5kEbps9dthF0u75tnTp7/2rGvtm9LU9x5
qP+R/AWvEFRdZ0AGJdT+Oybx9SoYHn7dL8Cibb3Ux/PnBEMm8/do95kAAGc4FFdjzFJUi3panR9/
osQ9FVUxwPJXH8ww+pV95Ku215i69WIu46Nu3jNcq3+addOWd+WDEhCktNu60pH1BvNe2S/5/a9P
v2jPDcI5ibsId1SNTMybBDACirgT2hYgqJFIywoSYfLOVP9yDg7eM9xXhxqU4bIotk8MiRZQEfft
8zhVbgC051nNwFpHREAVTflV10g4Xx4XSPMcTc8KPK8yKf4bVnAsxmxDhQxX4nQhSMa5dJC3K173
JMX7kIt4ZBH88tmqIV5Ze0IraHctU5eCOCFBSndQ/xWSQNhGp7Auj6J6wAS8XcTPyQeMjBZFbikd
2iTZwKeTqh/Rm9SSVdVdu/4yDduv+R3Y/h8JtA9cU3m4z+G+1SpjppU8tsETjff7Ju4ureYWVQvD
dJ7pdb1zYQ7ipkR0+m1sjdc4uJZjYmAUYyiV/ysSN7cteIYAKSPrEogQEQfFNSar9s6OqN4njCgs
ziTbdfx3A8u6LSLuqcrlSPoY0RdU7BjUK2t0LvsT3AmQcm+4Gz9QtSGaTiigg5W05Vmt6lF3ThAX
gwAQf4H8zb4fjKAP8akxyYdyF3e6fv6kb3u+LDDaWI3/KBuiopnDcVgCgzg5X98NNdSZl4sYy+7O
PhYaiDlcf1Y3IM1Jb9Y5HBxc3F7I+eSelZPiL91iScOOcooskspUFw2uH37S+RwIOwVmgubiT7Bm
wtA4Ywp9OmSaHRnoihqV7LafEso7uO0EwERCzm97p0eG/HSLLBVbyZNM7cfONXE4oSHIh5EYLjKp
SjabOLYaLobMFasEatP4CBONtrZnKaL6mql9LzJO1291IwAauGzaUgX0suq6wS4hae8sKJK7cO3f
OQy7SR1kgfNBjm0nODyKCjuqj06mQ2qBDoONv0qMk2N3FhWOjccshXkomGJWgk9jdQJomlpkSVG9
JKYbHiLiewe/BPNdUeZVGcHOFsTV7ohG6/pOUdi3feeb7TFKGf7C4JFz0f9Dbfj90R8xyQi62eOD
BiSkVSKWncvmhIGTP4O47UkLa9Y5YSKhbOFA78yWYTkSVio+lsEDUqiSl3rvkM4jyV2ik1/oExnz
dYyt65s+23o/oc8hqWPUdBA4PXfLoSP4xNkvw+A4BAM7Tz1D9Qw/fl3RFhNC28EMLCvt3E6tEWfP
ldnxzb3Ox2JKHi3LZ755KxuBmABGGfr3MwjsNpIWn26288DqVTyR8SxbBYydMSJ/Ej/DWwSXpr4D
GvAv8eMtcJ2ptGyVvPb8OkoQ8k74Zq/4l9F2P5lrnqw58bHBq74YBOC6V8eyg8wFSZY9qHCeKROy
h0aSC7L63Nfz2gsy8CPFXK295N9sVC/tWrZJ99waFHZ7/kujOEON9TnnQJwATvv+42rgcNGkWPG9
dg+/mLUA6eYswKw3Yo8zOqfEAFhj8cP+4OLOJFPBWlZc50o6ywqgzlqEbOYU1VTzT6jk0a28T3Zy
4g/ql2mIswmhpKxyc4HmaMI+SrA+LAgTAqvof6z/2DNu/vDBVIF2Oiz5buU5QWeKBQ1FQWqvFwAj
CA6dKv1KkrH/Ja2qz7o6BEW4sfaVdOR2mp7FoZCS23/jjlZn9x8PV/KGfQ97qmPJzB/Qvsjp0yMY
g6okpYgwIrdQod0SQKTeZGJxQ3Bef4Id6WvTX9xSww4cuWSHm/15lX6m/NedPVGUDisu0TduRiIS
ER6M3MFDhaixM+IJxAF0smLG1H2gj2XJCjPzH1OLjmx2XxWjIIyrQ0f3jgu1/0HyariokSHVsjzj
9VhMA1N9vaVPU8+EMBDTSYqsYO2b7Gs7kHLIqrki4Vkawt/J0qqyCGwIZ1dnBBhOIR8ES9XZeD2E
xOHwHHEbBIrC+CGa4B2P6TCV5u0XooU9RMH86dfcoUeKuMvqVdelHAWkC+P815VTBT6tpj3fQwGN
yWpWVNxRMXOisxVSjKM8csFof7KDpJge7B4pXCtQvs0FpQyNdKpkWbcRdwIcqyf42+DopHLvCC1n
fOfIe0QIMXlkePAodEJfEXrqKits1El9cSJgX8K+bsAckcAATfZO0LM4jReOG75KgbVY1QWkxp5U
N841J2hYG5voEQSLWtjuvKpNGurjlg29TqDHROs8XYdfu2/Vfb496jSDWNBCkdjbt1lVPsSkA7UR
204XAibgSAUYxUWfw3JY3BDnIKfHrsZdvX4G5tEPPyfsd+iNDBzKHo0hcqQk/aWtxoO8KzAM690c
TZem22hB775UpVQt48j76Tkq9BM2N0TQCUkikkYrYsHyuI8q+yPv7OdbylpiTZVCtLd8KXUPWleM
sfFrDdSw6v1cNsV78taplRFmjsRluqggdIJBFt5esUZ/vByxlMfm6Vu/GqhQnOyg0PGjkY1zBZhk
JdyR0acPqTPsOOtzThTUuASGB4sv2ixnXLd0BCTfyxjXZr2gFdvhvH8vMpbeCp8V12vjO1ItUDIk
yfhuH5seMY0YbkBUCW7wjjSMmkf49/fHiiVKAu057A+Uibi+KAo8ye/1Yex/iEPZoLuW6oEZXLmv
oiGrpDm7p652H+HkR5oqT5DpYr3RVRnzL/sqTcde1dvEfsG4HAtY0rTD0+JlEqGtlGiBSP1sjqDR
n82eQbf93JvR7r1EvrcvkemkuAkXiUsDsc7qBfVa8QpkudC74XDPeqLLrvk3K5ds3eldJue2tpFF
aQi6I2v7jqn20jzZImkdzcx7xM+vZ0PRR3JGCgOgS7VCWc9WX36IFRZUIWtFQ/v+TllnXefria1Q
WIFNkT3w6U9MWctQhTMMhIl7gAqaGbPwpAyEF/eDpZwV6dGlhgof+Edwoo6pls3Q5RYFiBH0l055
BVdp1zyjUjBj4OKUDYFvifQdugBW4TDIzKApSDu3r1EOl85BRqBu9wmA3fQKuSivwtu2opq0vUYx
JzG76QrFX2726lWpNGbGoMSb/iO8VPxDzlYWwbmx10qZx1V0b9SXCVVpylvAvbI0fqiEbDp7A8AF
PEKjfEz10nhJg+KsvEW0d8cB/+5vRmuD/lvKFN6WMLTIgSMT/OG1JU+1BdHpohCyQHhqsrz7tw/d
g7PdvZih3ZVq/SSos/nq3AX1el0pZX31ZsoZ/FVcLo13OwrQ83WKvO1x8PgNjSEwKr4x7S7nEZrd
2NJp9QbhjyAmIv6vZ8M8Hr6K/RgCzhACSD/AVTdHfJbvC6fytHUPKI3cvw/Aq/aVng5Sjar2cAMv
daTjENfmRckerGI1fE93m5Sl7sbyG/wpVA5LrdpQknhXqNyHU2SgnHBM2Zs/lByjVYWfkq5sSUzh
4roJ4x/EnBB+0dqcNAHRe+Kb4ATw/ct3MSLZZJkx5HTkt6Snoc2CJAxgIgT/LzJSoa/cD2zDjzhC
42gqiSEDCm2LDAHWvPGpzX4OioNxN6XGxiHRic/Fvk74otMaIfitPSEiTyUN2/AgVBpPkKIx01n3
Zx0gdXOj7l9qHAcJs79gK/HCluPsUREU4qWLjU27Env0gAXEwjAFP2QMyPSRJ2zTDy/JHO/6HVM9
NdTg6a4SVpMzSWshcbqR33naHdMrrAxTjuBuwXMnyb6tC+GCg1OmngCHEdBVJbB8QpGSLHzv5Kar
y3hnJunH3AKQdQvrOJasRq9YpYUFOZqT2RX2LYb4DW8Ob5Pr4LdOhaxVGMcmrcSBkRDzTlkGky+2
gZKDLHKTUgd7b8xqAhMPRE3kusKV9oPcDLWZ7qeNGvPkaDOarLbkexCiQtGSh0DdNUbLH+8SeDCF
64E/6Fgu1NyimjCaiMUetp70wjv7dNUK0QhZ5+T1Ky5frNq5mFAS/z7Xk8zAna/v/XQsVVrhDV6p
iknHj8ku3xGzgjjoOHnmhk/y8TIGigItaRNJb8hxCGZz9dVM4XqhY26/z4Z7If99nuKwhS6znzo9
zvuFh/+JgW5wkvbmWbYqIaoFkH8kUdt3j827/Gf4iaghFVmgrhU27Nr2PXKpm/bQkETSAelnEJxn
zU87e3CA6l44CdSK6YugdoUZNIvP2wFAIW2EMOa1uLVmzxYvyvMN4/Ee9789R+cOfqTwC5UYMWhK
DGKg0BsnNR5eyensj+6qxHXQjb32uLydpzntE0pG9nwRKEq2sFLpOyF/qnFoAQbgDcNV7ZNt+grP
ILwXaykg3C3RYQhJ9JV45iCOc8Q4ImlJSVc7wcgAdi/LpR8Ha15x7INv9mDKW+4hjhR3gB4ybDJO
36hhqedV0T9dcjShAOCEese0jpXUcJIqj2NxtScWNwXvmHjexck5XM077A2cGMqqrEGLDMWNfhWF
YxSKBqN6LYeqLuewEwtsfD3QebKla7gvLtmp01MNPjW0L6ZNWS8uuEgz1Uls/uxQP+yGRxpJx/NP
oXHp+IvLuxQ6uks6NvrpD0TAvBu7lm2eTTDUjIp/SE5Pym6gRbAQEQVJ5gL2R4PNrfMAowMNC3tr
AzTOQ1isVMksGJP83h4DH8ksqKNnAv4oVaK1HtYVcdFubDaWm+fukzZs+37hG5kulF0OMhBrzUAt
rKbMC6B32qmC1zsDWP2S6e2QUQd0t0rKZ/7xAPF3wt4NCNNvEXZm8QDd5Nf2Dbug5IF8HxLkGp2B
hEFJsPCSEOS+oNy2xrzxV597X3ndNl7nY/PyETLDNoCoC8QgjrErcB1BdDXynRHT37c45pEtEQDQ
bWbirhVzJAKqjKWPY9qKK2qyATvqeynqiM9mrb1vQcOQAUMblWlQFKOkekMeiqtmuE9eXlK8n+dz
NDYFyvmpdz2RWrM3Nb4HdQV34XsxYFSu3vdqzK2NmEpUgFmya9oMX6VBy1aHE8F1XOZ/650jk910
MnoeD8lS7GIo3usJ8AUDVoyn74YRE4kZ+K/lpQgTbwazTb7wLKnVmICDe6UpDemZ+GPfCmqeTaWI
dgRPOZVWNcvaiW9D0UjoMXTVNBKO6uTJ+l0UqRUd3sVt4FVq5lIgxVnC9pHXtTJqFm/8mIQecscw
QbOte6T8DEFTr+yj25kO90Rus4Ui6RuiU9PmZLcsPkJVSHmPYPDfNpxgoTdI1rFEjFPGtVVFJgu0
hKsgNmydPKk8+qunVQgPQkH0RLDyrd1Z2FU3Tq5dyvxW6E/F+blUlVdtHtX0oA55iR3zXnPuXFMv
SRq0BCWdtcRlCmj7FCpl7b++M6CpUIwjavRKWXEZyRVWoMoYo/4xcDPOyyg8UfDiv1Ey4rPwDdEi
Qe4Fj6v0+KYL6c2qlaHEm/jCiqbCm6r40ilA2b4FatQrqYJTcjezwSrhm7GstJDb3hg67QebgQb8
kKrry6fT6zGBqrWpG/pU7+/aps+vXACWETBCKmg2h6UgWK8EQInKGiK4grmPzuof0onFC5Ie7FGy
pTGhF8J0fsTGGEO9qtR7kxJ/z7I0HrSxYZBRweZi/d2A+sKe+uh9LE5r83ziKP6CMvklwvtkyfOA
ZK/D32aPiBWz8AjWUhiBy5uvUbQTq6/aTltDGFW/DL6wJzyapnVovuIR5UXEvHNE0SsQWUkmLgio
ghY3dsBIr/jVmWO7Djbix349oNsdwnM26/A8o7kgfd/1dAd+BpMcKMltzpmv3KesvuQolUNVJZhq
yfY4NNHm7KBy+CxQya9vklBm5VLKLCoYpyIeUMo25G/or83NlegwsQKSilYbs2dmuxDOfHsGL4c6
ReOMRKkMI+QuoSBbcfihPAkXSwIT+sWfICtqMddVTQGndCt0Xfgl0ZPX5WpD63py+iYg6GvZk+Fh
u7pPx143KaHIUk58LC9Zyo8BIFKbf/LG6bZIYZDvwcq67jTaSPZABr75+W/RuHL/plV5Lb/3zeik
/pFr7FJBXxiXglB3uZUlPJEgsM37YqzLinl76TUjw204E5PywzdXtW+Rm/fyPmquAoETz41yRIQK
warSb4HU7BpInW+2SU8airBotlAGBxXBjSKZXmeAFUsWXJUDdp2NTHM1JJg5c1YE4Cu2wd8FDn9v
7uikC680NcwQBU6ITjBhk4Jymtob3THxNPVkWbdcWhKEEhq6JV3UhORyyTNmZL9udQ/X3I+CyR63
s6UMeflZB63EUZfjd6TZsmhLnvNl1VxkEGy/7tUzrrJ273fISbcxGM/SLSCTMaPM/5+0v/eQ9Hrv
e7pMhdtqnHmSNbL90ntzo24IOvXvyOF/WFxZFJIEwIKpaP67dEwgOZzHLV8u4PSCjpIEtpchNRJu
7GlqbdLlpshCGCTfn2j2VkYxrL0O3fvMAwsIsPa3YUW9nk0lyIendC7k7GweUnE+XCt2KLga7hM6
3VsOP6rXRtXJ9OlcnoYesB0bsMQB3VhsUpZn8LAX/yn4IDzKo0dZm1ArrOor8frrIHPMJRpUqnxt
FI7rdXpoVgMHdmNEgrE3d/fhkRhjwNGUPbfqogGMQmfdPjD/fkk3ukMRQBK4YlOMBoswUCOss5ui
VyMvVIj+a5v0Ss/OCUdB5zzGR1Z9CVzEESYSHe/36RKPgNZMX8H/jFvIk24mlujKUOJvSYzPOjiD
T24VHVvMZBcCigxn+fEAfyMKEiEP+tJieWKjXqCh01JH4CTudUbQJv7Z86azFEKDWtWcPQDb16HP
OerV+7Gwt6L18aZNjuQPC6FNuF+9yqoFek9U3cUBI41oVSJAzedLosUJrO9z3BZQAaqV/dbz0xR3
oCN/Tsrgh9YTD0YfZVMkWvTe9Goxt1B2aZTHq4dhhiwwVWsrqZAeXHjA8GWvG1QMGJDZjIJY5r0B
9uCcxSIAP6jlTfgtJ+M1XkrO8wCMorCeDNqNz1QM9r4LkOLv52Eua2XjkSo09XENPZOnTM9qTCpa
xF/c3hpiNUmsvUvG834vXW6qGWB6rPYpJq7ey0//TwVpdz5a5UUFuqueRj/jQACYc5oic+QzAZE9
4Bpu3aoTeZ1tMMcd/l/q+6SODTF16LaSPSUIpbWSn6vBTV/RcHMr91MQeN41+bByRgEyARXneP6s
28CXMBGJpR8vOBK/orlpEgvDsVDV/F0GwST0HiTCfUfrEAjiquYMjuIjMGp//5yCZDpUyH7ZSLYp
7pvYktP5OzZmJL7hcFDzm64mz3GlpulKgZeSFlHJYkztR3rWlAc0WhEhLR5xJBzNjK2PMFdwVSZD
NwVnkUyCoNyK74GWW9ZngwINkjXIV6k5WCgOHdQ2WZN8zCVb8QzigOPmHjgIOhN8kQTWcZe9u/sj
1IhnhCj74HiwN1DRQkT63Nt2LE2NcPvEvBjYqzqJ6a0YRzhA30SRu6jhj1R/6M4UR0FMx+ZqiGan
8Jb0o2zZVtuIgqNj6zysZC65DpTTsA282hPdILbAFCPI5b73pS0PQwjVfNCy1CededPUoiS+IBfw
RAiaa39ub3ECwKuk1lHWbK5D3maN5fl047VelnN9beIV2fmxnO3AI6qCku9AlMY9bQyYMpSqmgoQ
ouJGuciFHZsohf5tjSWfggXSbueXgcCrq6jSEp9RRU/3+qr/yi8b9pdGBWdT/bew4GHOxr4dUBB3
6z0JCtkaukBqwQ/TAfmTmm4nBpgxvNPn9Nh1A8ka+VkDjKkpaEX83SH5fWFqeFT9mt6ZZCETDXKc
uJ1PCMBXeAwREFKjycq0TahU6W65iT6aswhadsz7l01fdWDPITiQa4oey+WdnvDfKJ1NSXizi+d0
VJDoK3alYZi/xjrDE8E62hB6txk31jWzCgKVgrQSfTtqEEIaYiH/eFaKMXZLmEIkLi6hXJtmvZTl
HIpldaxPmy78VF4vT3Vk9z6iDt6jZEbaFVK0i6Ea0/oqigTgr3KlTDlJUd50i+eE667S5e00zlFD
qMBehMt/j8Iq/yXmsdbOCqzBqijyETFEH7wcVyPBltqw4+S7a3EVuUfAiTsaCChZXZwlXbQ6T+8e
wAtVjg70Ct+UkGuMhqh5gGS/fbAHq8sR2VK2ePDClEC+rTfJRym1Yy0EuOPwIQA17AM3lMr7JJzr
Ev1Z0yAKc410zkJzTAm78qE+kAoS79jzNR3mDNQa4nPpz1VQlF0CL4GZubx+X1Jow4H6p69ztPjH
jeo3hYAz/fySWfpgulBVOEsdYjNXqEVpL3hQESmPBKWqwVqv9SnVXuGWi3B+zXpwyHkUKAExiuAZ
UDzwwr5FjDFKKP/fYciZRj2axsq+n3Abcj9bT1wZ0PKDXssUlypz5OPNNpadaTnrzTWNURONl/ax
jHCO8QDANvPwPUWHQuDEVXWQtrRYd3WOAO/n7Y/KxpUdn47NxKNQuBTkgiksUjHH57JxSGGz4nvk
aFArAQeWfHHqAtADXXxJvZvge/wSF1HukIYi3lMGLUGa/QJwVVrXGLPIdjuKlmQ3OWc3ncKtbARa
FYeZZIVksdlnS1zd7epEaSoyede/xHoCyJmtWSOHzleEWACWEpWKHj9oTFdaZtGTZQguqHqiUZS2
cnqe681+FfImjkMSj4qnslBbUQv6wXpVkCdXmdQO+a/nYM4jlMm6m6/mhaQJi57GKOJ2DNIDrpBn
7qSCpTk92vj9+QIkrXJDd/glRIczdQd/O77WojaboaPZEozsofD2gK6+Zy4kpx+jwobXrpIZsMNF
5ouJlYizHygdMytVBU/MEicnBHcm7rTw0mUgVpDoMGmL86uJNsIz+2lTQ3g9njmTfHj/+911yNR3
/RficBU+7RtoMxRtgBOJ9BFupQ5+z3eBMFOvKlc+T8ZYLAdZlsXYzfLz53xxgRtjbSoB45+VvreP
q83NpOZipaX8J9O76tmp9iF6TAZ/CCFFJSB/1yMzT+I9ppI7TbQM/35GTpXOcmnfNMqPv35W4PH/
HApC+X28rxxJQvYOKCDaFifbcSfvU8XyN2MfRnLMiis8c94aYP3Q1WqWfHlVY8804E2WJspNozMv
Ka28dGcsSSFatnFkPcM0TAijbck0CkWdJRjZuxW+9HUmYV9NSN3r1HVAvSiohwwNYG3LK0tgEM7D
rQnPY30jITBG7QW8E6924uBlwn2nufXNFnrpFjnKEVGcfM9ULHtOtAxhX66b8fryrkeoUZzLl04p
ehMqjZJsa9LSwvXshry4rmk6GqjYztuY5KjP+kluAqqCUqrVRVpsR5+iGcrymmQI/PtA0HSzDW3r
2a3/T57YLLfH05yMSrLkht+NYzMmy6SNvDtQ5b/cdBv7HIoeTjesBvYq4I4lW/nV6hG6cbgmSkMc
5OCzGP343pXAGvGozdsy1xRsqQRS24JngewTNffEIgg1TAORoeMwOxlZVE29R60xOkMay4aSWzIK
W6Ss8lTz0jeGYKx6e/nplSPeYkor9W8Cn6x/kTCAio/hc6XTzeCbDFq/xZCOq/E01SF9HPROjch+
tkhKfDSgkhd91KA2ZEfoMguIealLDNa+Fznc4gRePzeUWnBserSvNeWDR2jJtWd+aR0IMyqrL6bq
GC1qQaj5VC71+OaYAIWlIXSNtBtIi+ioXl+anvGRCt4qe9Qe19qdgLc4EouYeTsi+0qE8xNj26he
PfhpgBHm5ga8dBuZo5LCzxUFoWzT6sM6T6vBEJK0MSJ26D7rhxh0Bs+Wp3On3kqPvrh8VSYhlhMJ
H++9wetkFFRoBc9TzJmDXOc6HqUSvhHuNCEguUdqQTa67v504K+znl96zISu3rxhs4PzwnVtlS+3
qhZ3BLFI1RxLpM1uKSMypn32K5xHMT0qkUPBDfVrdh3Ddr42qaW6ZjlEZNhReMK94yvVS2U61A/3
zI7FI5sf52QcMm9KAOAlN2VLbdwe8LUHHbBdfGq4gGnwmb3HMiakIeM1oksYjE1aidR/jv0tfnAA
Bo0RZPQWFF8bwRbhvkDPtUZmBdlTaB8TP4qK4QSZVnPOW1H+nU/eH3VQ8egY0IM02sQqyDdmpWca
kHREXHz6yc3wwupML0a0BXeTxCvoBCirT43WhATtPQt1TkMiRapNe0t3Qqbg/NnA8DpfDlqaDTex
MTXKQfyYxeQna+kRvomfYBgJpQ0d570KnuFkts3cBpdL6HjC/0vAAo4S9PsQudA4zTAgoxKeKo/Z
5mcQNt9Do07HPf5EdRxN7CGnIHJh22MzpelsEGV5S1+dhWLTFE0+LZtAaFj7AjbXfKo9/g7kh9db
QLhv26b5EJROcwNk8j18pOVF0HPeHj25vkcu9ABuBG6KQrnTSN0v8+9d7UHkjE53CS7HZWT8TM5d
B5Nz4roFiqPYE5OSX7G7Jk25odRG6zHBC/mbfRPpLei24yS6MEvIx66rs1U2s86NhIxyI9yBxRCQ
l159swA+MIQM7N+F+oRtdZ9DI5LgnumeNTbpFvTDMNG8ghYF8LzJWv+TTRIKceH7nQDy+MNjT1uX
znt+RYaKbbumYKNfd75tE439SyhkrV7zxhxrJLL0SA7jTsujpKUG/w3bN2XvvsJMnP2Ox0zj/Fzc
TM+VuKkKLiBmbwmGEoBsk7TJmi1AZjC+nEIpl09pVPSJIjb/DtELxJN5g/ZDViOdCT9N5uruhDPz
juVohMqKaEwJaDCe9hFJ0dwvfvcSVLexeWycxNy5coTNZTrUCjdka6Eo5J0OtI1bo2xtbh0n+Y7C
Dh+++KNxCWTktVZfmvVdeV7rqi1cJxsJ2t5RdBIQhq5L8nEANKQPX/jo6qBkBopWgCfarznbDbwO
QqBEU+XQ7/qSQPAI1MuE8GzkV/fyhixv0C+ZOk/YAibEenLYaSRUO/b3ixDIMD/e7xor9ivic+Yo
tXwAH2mJtNGLvWmldMgg5y17Uk0pFjbxRn+uggqgLNzSuVH/IW3cUCCl0aX6quZRnsV0CHa3a9/t
mjnbw/MlYyI+pNt7xVKEit57ZQHRGQzmZhILKVd9ZSyTSWt4fCJa2BZmnCchPqfAxr8wAueFw7M2
9UA+QrYPqOeFwWR4CId1BLpKe0+XupS3PAGK9GhPqSrguhZWILz/V2S7SUl/6EmM0BR+KPYbJnSF
DHZpPvVq1orWaWXH8JOHaVraAJaISN0glzTzdKRW7aK+nFOwQsZFRuEazI3leZ5gHt37ezrFT2NX
+Aj37/BBMFkZwqKs1v7MewbHyQyrUvjuuck5qgAkMjowBlByrZJaTBwl97oMnmloFbAUU+5RCDBp
Ex8JMAvGmYpOQM9uI5/cMUMNdAKjcuzmdaJYdRvCwQi9jrneQ1zzh0wpSHA4aHs4ycON1FerhT2V
Vs8YcWevdcnDMRPs6qHIYnmnQpb5Fqr4de40gSmV2GgoaLwdoyeFLtkp2LP4dr+zy0UAlhmuPMlt
OaZ341aHcP8hZuVIbftd93vZclf6p3fm2kqdKWfUnkOKXTY/TXgT1Sdznv9S1p0n9OtDIrOl1ZW5
0aiJWJvtYpIRYTGJ2QMBb12amqo4GD8SiXx8kxYkPfz3qDV63LC+/SPKtHsahfE9ugkLwNNrFbu3
lzLe7xYwzx1Yu0+ZCASxnrQUwiZkoHbWMBmd3VhMkaqIAfXiRVWWnpnEnU9dnI9DnqxkQgybL4zz
4J9HWsmNhgifgHWKNtGQfXGdJxio62vsSEn1BGMj0anjDalDQVaX9okRRxyKCrdBTTm65Yf8N6z1
W3qTZszmhx1VSJ4Dwgse5vSFtCCutQJx+FCz8EeLlIi5rqXIzpftTzKEtqu8bfAV/BIaXF6eq/MU
KTWLhIDcL9v3Yjug5QNqrhQ64T+PFWiFfd37VvR24Qb4gbCaLdmv5Kw0SQMSQz2lcTJgFyUkaNZe
U9ihDaNBe5s1fg0lnh5MJ9xTbdwu2Z87qqoOKhvLbuMke7XG8iGJnCVn4XBWtoetA40y7RgER+pF
e22j9oIfXf3y/OnRFsP9Alhvcp4/mRuXTj+Szgi4fo0+eV5qI9bCJJMg0xgevQaFKXXuRxDqO13B
jx+q4pvjn1lUoZFnAnXuL50L+ynYzcwIWjO9jz9D3BTE5NuunG/8T+QanT68yKTG4fGyvvDA5aGs
lUvFTE5n6daMWR00F5naTypBTCWtL5DlnR1ykh2KuL5JPK7ntT/h5VSy4sRHE2c3MP6g4sddWhMP
XYAuf7GTEM40TwKrKDUXD4Jxx4gOTySXUjAP/sAeFLquojkFgbT6OXEzsZ97jFxzleg7MofB2yJs
5+b6RM+AMzKT0S117obz5hFkluOjq5FAPqk6eJQfGuruaQiCj8WSbfFoMr18uma6pf9VmukfY9sD
ylFyiDbRcrR2HmQEar7w8cx1m3GvbsDSZkZOgNEQsq95WwCyb8Msa5roVWoHnRfA0+aueOBK75/y
tlefl4McLexaPB7sC8rbmp+IzyK+vXXY8ssFJsqlXWPRZrUUF59QdrO4Xcl756QTK5odAAzGDJIZ
DpCERYsgDAwwdVemr7w4xTXb/AWyOYyhMX00TuUf/hRzPpMhw4VnpiKetS/MB0+WnC/0URaqfqlS
ywP0SVW4/QsZqacQJmJvFZ2to8v2x5i0nOBKCx3hVlP6yNzw1PuD8kdJTYsofWkg5lmYDqsFSPDp
nnBRjzJSQBctPh5fhrWvcvFtFpUhGdut0LzPhCIX2rFNm/oJuvlalB5gdKfvlvAjJTjlucCHQ+mu
dl0tzBTGtQoqLZkgVU5LncLRezdKr6JFTljQl5An5lVFhXPR0Y/m/ky7Su1ozZOVdUOD112+bQpC
zvWiaFa3BQEUUGe5xgMLEtQfa4beqtiJxtl0StbvKBPDkj3S+DmT0JPv3vDE5gDbcgqfp0fH1eGl
fTNmJXnwHeK+UVlPUYou0ZJJuYj6wB1cCkkteUHJ8yHKpIgYkL5UgvmQC2lqhRZKrp2Mgp12Xz1v
W9IS3/2znlzBoOeKCajJGNs4l4JdgTjRVORkoaJ6dUCf7AjkV/HnJiRfL2dU7xLDCTMR3if2I5iD
Mof2uILfEhduev5PuP3QH1a5UJ2qkiyTS6vCUEzKNLUIcw0olQIv3eYVQsygFmAXyDkQydPY565E
Cv4NOpSczYYHnwxL//PQaV8oVlYQ9erdH9/6swgynoUIk6dq/Ua1SN7znkrTRZk2vB85sOjBs1jS
1CVqHOL6ukRvzu53pEQwJJxcTdHXG0w7tD0sfGBghPlUzyuJS7ET1U/ERehCyJtp6ea6+ryE7uXU
ojMI+Gv0DeUCupveiqLKS7+jF+Crv85p6l2yF5JzTNWwPK8tNdA5xq5j+mFBt1UXUqqh6p8GQh4r
Az6hrvK3AIAuu/dd3HqLtsjWQF95FeA85jyI1JGIH73OsCPRlDuCrq98dmF8gIip0vtKpQ8kzlit
LkjRbFqQyvWejxhzsNF0JH0MTQ1frWM/QV47GMrZeD5fU5i3iMEA3uOQk2qz/4CQmC1361JxroBw
sJWJ6hjazi0Rqy5Lv2fcFSZL2rKQtXM9LRaAih54GbPip8RIFpVlW8FBZrFYmWtWRcJA9ArGvvZZ
l+UWypvsCcT2b2Fm8KH47GTpQB534lPfhkB8XrC2Vz/ahkDTN2rniYHF9Nk189BS1CP3ETfECNUu
jAW+iEBTBHmrQJFQP72mCw0cFJ5+EllSaKe2+HBzwqlOYKfv54Psr4BBI+axR4q15IJqJNo37kQ4
9UupuaFyWwG9R3Ihh0xLqCNQheIYGkL2UVFzmijwGHXmCKA+oKiHqOut/8jVItqQvpYs2DjEDzqY
N7J2yS9ZfPzCDGJ9FynxuVI75zpAhpkqOqTW+v0fnOnYbjz8U3WntZcrzhyUrpHzNR4E7wOA1GJY
vA0u1mTlJV/uDHWStEjuCMcLgQ+G6mZ2nOJFt5LNxir4eK91lPjaHYCbktOpuqX05M81plQ05A3e
XhBjxTISZ9Xd96Bly+Xb/Tni8OnpZ0sIE89ug6UZFgKIeIA72cYbuITW3jUaQ+40GzV3DrnRGaHO
U8pvI0G6GH04HhrI6nK597uw9VN7izY6TZ0090aESR0PSdncml7+AymapiA3DWNDrAI15/jOhT5j
mVzh8tyi83KpyEw5Sgt7cWBHNBNw6OZdFT9AdJ3EC+l8SkGEjxyZIWaSOJMH2R0nESpnLuHUoTCn
50bVPLBYnRCI0LkBVmu9j8QsSVFcHB7aALCs+pOK3/ekO31dClvHUIoK8CX5B1h9XGEjtyvSV4ag
YwoRCgxcgd3xch1fE5fXOqIaPLRRQmotWxhSeV0T8nAV3FzFIr83lsaMJcVAZmIvfoiu4NRErQ7R
eVOi3BiBgvPAQ+NVxW7ntrw4JAisZxHFp7yVJqRtkSaj2uOIuFYLoAoyb6LajgjAjPM/oSC2SAVX
ozRvpGQ9LFRgHNfm8IDExBdF8xDkui7kgGfMwgZC1aUl8kDx557hjz17R2SBViS9saR3csCE+Lfr
lbl9mshgfbkWsk2PJR8dDNAwhFcZXcjNBD4siXzzDyep5/kgmGMQTV/lCF6Rzwmn72k8VcSs3zNc
OEizdycXw2UI2RSBkbYJNSRcmq52nQy42KzFhwuzXB6ro3wqESZvUcTIXRvNHTUbBobqmBvyKmna
MavpGFGFjMwQVX0z+XvDcv5L5rTrzFg4PN+1CHW94BNLcbw1Ea9C7Ljkfy9DhaluRIgCG2Wae8h5
1z+jP3xQpJTu+/+7XRsSIrErQrHtoQG+x/o72Z47a0F8JOqx6m8IC034OEXORhhf28VVty8CReCK
GzBWtn/FaEU7hIre1482DVDC/ObXlPxLcknyWkUfNscp4aYKkd+z6JvhadV2Jc6QV7eQzGRf7NmX
7wAR1SmDthnnuw7vatOtEwTihuTQKqfazHEBGJmYwCW4rYPgrrsAsrGMLd3AfDR7jUtNVgK0k/wX
7VQ4TIVy0UQ0+3iciaIlx5Ss9i8lTj9fKk4FMQ2IG6CKLTv2dkn2HMqd8N5JOKL6DduOZY/kwhjj
ENQTOZpfcN4WBxKUErLEIO0PIwPT2Kd8qM6sgOu4hVRzCIPzSIU7+bSk7OZD+/ODZ5x89723lKUX
/Awe7YmcUC0NL6lAzdGqRLIYW0V0Ly1mAzQGUL//W6r8wtgrJTBQJDMWAc+ZyN/WKrgP+OyoI8xn
soJCdofBsEgc0VDnt6I7zz7JvMB+hjYQCTw0e9Vrf/ZJbvWeE4SQESZWumo1yEKTDXGBQDU/sYGR
xOD46voWk37yPXC+DWlBxXMUTMXtEjlfQX/oN0JZjsryhnUhAJEylkjNgHAEusUrbCekS8pRApB/
FW1h+0dfiMTC8HLMsiQrPq8dGY40uamXKcgqEF62Q2i91uCw9wR2TI8+gnIGXefcw7PVJQmfMOze
TGiuo21RJH8x9I50edinFGHB7ehHb5sOQPqVjg/i8kLYpv4es9YtAbo49AlSSsauSn3kXJ1pTcnA
t2CDdtlsm4bhJY6hYdvhtLT7RArbyo3ws5vp7e//AaQ023hBUl85dGdEzA1kDqFtuV9rbsOmVCT4
XtGkuyob5yBNIypV+FrEYouT17CnC8gUenwFl06HLtljpYZ68JlJ72UzJ4y06BbvXt287a+Meypi
hup7Y1T4Av/YuSe59ir/6EQleQ+vt8JM1rRxGiCJE9xNU5Kyn1Uaq1M83kCeb7ajEeD4neVy5VIn
DTMQQgT2GDzH4+vJpnKruW5QEMVa2tLI4QOOKyR7WVO7DxyzfT28EZxtkMlFHpxJmDPXWe73fI5j
iT0yW7u9uFOW7BimEPRgOecEokwkBFUaJmCE5NalBK0DI66xQIuqTpATnP7bTChsjEaG7X4m5Ny5
xk86iO8mGb7p//GKhGiwxfNkmeFZFV6hW7YlBYCaFi04LM/Z0usUdqTCTr4IWiTyYdnwDWwllPsf
Gb6FJWAt/TQLMbjibG6Q1LoIib0GUb/BNJB3iSMK+TIVhfa231s11u+4KHzSh9sT9Gvz0xwJGjTI
6M636sfChEhmK8b72Y+L/uKIddVqS1mIyei3OOH3nCzpuIn4t+Fyefp1rmqNDTdXSkez+++Aq1dj
dIKARUmKpreQ3Sd+FFiLeYhENGUTh/5aYfm14rLhmdS9Ioq3SWiF93YdsHBBZiNSdckDTNIGVVTr
r3m8vcEJy1CXthQxM40Q5gOu9aG6heESgy9D5cRBw3+NR7NrC0HMFPrawQfd0ryHFSs001NNibs/
lmVygh2Mx7bgnuHY/gKKlRh/OPm8+PYSab3HaR4gawVlGP8422o1a5h22DHQa5sTqWdXYpNPXfTJ
VIK2t/iqqmBnk1m26AZISHFWnNd4bl438JAtGMVx7qJDc18MLFAtjUG5Z+JXC4X2mNsXmjzScenB
5RRmSQwXYdk4Prb4qF1n/k7F5nv/W3AoJSQ4mCd6b1vRMOOn0HvpbXclGJCfuZRP4trgyl6uKEGT
3elBBo5q+ba0sr47N91KY+MLAz6nLW76rjpJZDexCfsHLe07hApz7wD6eHFcnLYiN7+tYlTM4eez
7SCircjiGgJ+1+qByHWj+kjuzjCzu/TX1qWsN18Ej+/lvtUqLecoTB2FcEvOpPujKasxSMPN/Eez
EekHWCK46mh2epnCGgDhgRw3iojBGaBaebRMhu2Uez9GXL3qy2uGyK3PP+j/qz04ETfgeWIqdK5o
GKX+/x9gRi0hIfYUyDED7rxYnviBvNW5Dgh3/F4QHks2wjRyM5SwngmqJvj9F5jVvFWF4Hpa9zij
6NEDv03lWeyO8HXL/SkDmjFZRIIPZyMVPra/G26dK3KBGSJHOutdZ0VwwVuz4itjEAd9lwbs4F6i
Rb/1vBrdfe6Oid6yymsW1oQKpV7qG4VMYFFZysGO0K9DDGVcVfuiLf6/nMhu36L7iCbboT3J3Hzq
/VAjJ8jUQ+JOgVwSmc0xJVK45+DfUYFeZXLbQ+6cm35THHKQpdyTghyxZdk7OOoCI7gevdfsBd0G
RlprPMJ8TG9luD+rStiMN/4WNwTHxZrK/qtcdgxa9oRHyZoYYD71UdpUpfiAzOsac+3/SMCRv5vc
nM5v256hwVzP0VVSwWSU9kjtKgTK7HOKTRIsS2M/GvZUejhPurIFsItd9Yq7K/IpEi8o9+FFu5Xi
kB6qGwiV0xmWjlPWRO4XNUC8ynHbYh6K0wgr/nmSFPwYuCbwK8CaEFbzXj1HwQ1aph5GY+/wuhbJ
tJYooZlYo1SRCOasnHWKM8m99FuODlLbdBBZ41f/clSylEj2YIlHfztGF6owXZj1bHitw0dYKIpI
9EKTOWKfTzznJlq4Drsh5kzVL822JIFxgGKPwKPyZNdyTOVvxXwHbsXcFsBgmepPs+rcv/7iAuyP
PHxh+iF/e0sHD1Rz8e9psqxKa5hNtLmZgU41IXKKAPCfYHYe1aKCb35LUTxfQYgW4gzTCgFdhj73
SyiHwluR9FIiOZ+HlADC1H89cLHsmxZjeUcqULnsVqw+g9Pj5B1abEtA5M51aRAzzWQIWWBCDV/d
1IDLurHjfWiD3rz+8j+OGBArKWYp833CsC58BEb7bBTMWDVZ4ZnQxSaZb/vT1gxpaOCwwj8YAoJi
jZVqZlZHb45uiAHuApOlePRxZ7XlOocGbkzzV3XXBoILDKOYBvq102q8h3L4k2AdLNp4SzuLtD9J
uyG80vkV4p8toN0zi3JUN5ub/cSEHmYv5j+3I2Ww1/agcdAamWhWc5nN6aKhJH7ZllD7pxqtL6ko
Uim7lP/0uL4skMH7tuqBIBhxObEBmp0mj2SkHL+mLdSNLwoMyNkQjMA9IsFBYOBSDIuOX4FaZgRC
UplFs34qGTAdAymzqFoUhmsVWxwPZDsGLR5WaJXdepdLSwQN2DLCUJnk+Pvn9wbAYNGLsjkqc6e7
KrEIIc5yUg/2ZIBzm2tf6pxQVIb+oZ+wWuXgAiYQJIkYlNR9D8KiT/i/6Az9bncjfvvu2aEPblNu
49TsNABdNFgN1Gks7DjQPCo88zw6xBmEzU41TXEFBlrQJnp9ni3VllII5BNHguNK3Amrynmj0W/i
dt69+/tkp/lalg34WOMYf+ru9Ogwem+5or9CHzENUa+0yyqGzag6YRN11tx53Ka9n97IihlBGm2W
w8mwnwPYnRpEVO3aDXtwY0i3153LDecVuWVSr7OYE5jTDjQ/VJxzqZlWH0Q+lk3sTiZC8ksLOgFt
vE7+n08WxX9zvcTCnv/sSJRFaJ8yF2hOw49RutST/E0H5XG9oW70DPVi1v8rxLFvDRr6ArWaycQn
AHk78o2zt3M3WIV0EiouNX2TDfMvc0opMtHvypspaREGr7qv38OCdSZ/DZrCqCcUGiyg2SKzSLiQ
/MADBixTqn3c0CDbTNscbFLvTTUrH7eiyK2nY7g2FDJ6ThQmoRiZoOeSr8d2ySyVR9hyV2f/ZpRo
SIY6vG3q2KVL15DKun1GPfc2/DwEU9zjduxuDoz1LBZQVWLfWg4n+HPPunfS90640YwhZ/FBKO66
DE2XL2o1AEzaYVupZ06+/iZm/cXxMjnX7EoJqZhZgttdNr1Lb145UtPXp11Im08htg6YYWP9hYKb
pygXUZZtGD4EIASkMNqwg6eU4LkUF9yRaPawDX/8Y4tFNrhFKMpCCVkFdl+Xe/nqe3F0IrAMyAUz
Dl04Id2qyh1G2r+30zI29Pm/hjs7iRhprINDoWRnbuZtq5+7FTdMeg6kxrrhX+YQxyqwVTDb+uj3
d4zyRrrl2dpEQ4+x9eKu9jBtmVgh8E8K6SaKKJjU8gKcPZhoHNUBUeadWVcRHZMuL3euVcz42aBv
wnt2hGHgAU5Jj/Uj76Tday3rJNWUiYZ11kDVrUglr2qQoO0BTGD+qJNTonYhiXcxMnBk5OeegDQe
J8aPvvY8gVqSIWHPiwzU5/6LYAN6H2QH8revpKO3cTy1tRiqx9tZkGxH+ihAo92pwZ24Wx04yt0k
BIvHNomhBAGCEOZIn9hUvo+ms7NcUDsjy75YKU2DfrluKCpjaVdq3EtEBjBOJSZkzYJ/diu+WU75
4IFmQy/gcsVICzewz1PVdk/SpkwQIXZ8RE5iQ8ciWGMNMekLMNbMQK0NVV3Da41xcAOKJZn2HuPY
Fojs4obEL8egsKEt8PiHYF4ugN9YJ9njF52CE07e10KtHDsBkRgEeLh4mt+pH2DTlyZ62WBXYNfz
FwZu7FtRAg4xwB2sBtbhomJt22I8KG3jUUKcgFhcInbAvOnG3xhKQLumFk7ZCHAW0cE0sRtqRFkr
Yesz8AiXFYPzZZfEumYMrX1p7K3TItWtz9oG2y4qrJboDot2bUjtZUFJ5Ph2mNo/Kxr5/uXjd38j
tqxkLFAm0ms0GxZyJ2Jb9RYJaFkASqeD3HV7GuFqSfCHe/wvmO1LXPXLM33fheABY8sAMkux9HI2
wLXTh7essiHJ5LXLGrzwP6tiNI2G12LB7UELLZrgVJDAZ8Gmgl6+JPg/7Shf90W4CNM5Rm2hyav3
Ow9dsG+3m1xFACzBKx1Nu9zqEsThUs/SVxVebVf7IMubncUgpm7IzhQLJEmQdphkUG4tJhE4oZO3
AhnvbeyHs+0P4kSUISMa/yjTtBwOeFuHxnBruLSf2sNW2hlYYGUsmoxsV0JjHYu7o2hG+N4CO/iz
NU265m7MKMh1H87255sao9S22R5cY7iGh5G5tzgZzuu5BKsot0vZallsnWbeUu062swNPUkU5Ran
fIpgliGbyJdcMw+owtuQBOprWyv0uDQOga7F7cSeObetZwpr4yJ+ShNF8aW9Cgemwyq9iGpqvLPc
7NXISm71YuRb6VckU6ETWXze3dbV9Toc98cIvSOhsJfKMbo5a7DBuk28wfrqa0/R0EBeggeH+Utd
SjI8ermqr5YEfi6RsjZiOwkUG8PJyU5Un/9Cji5hK7w141yPBl+iXduAk0YbKhdVwa88O6Ozaenn
ujcCDU17U0YCZcz+fWbEqgGc+fHOZPTq+aZ7kdLlueehmOQdhDWxKhqKcuA/+Tb69dytGkFqB1x/
go1jqpue7Z3jAFiYLqJLxWXAQkQ21lCmwR0LpC1HpHjMJXKlLUKxvEBt3AHVQ2LhgZcUjdO1TCVj
BSTGMoUJbg60EDIm3+DZKqmadcuNlfR1CSUcU5Ttq5TCLf+1svqvEMSNXXBcA7jMA6HakYywd5HU
0NtYxGdFF4qwMiUqrfOMUQnfqGScg1sVRl4d9wUJiKhY4Bv+Gdw9xeP6nVvKbBaJRPnQ9/GZBFq7
SZj603k7PgRSU9DVsYT2lv62hwO4iU7nVYHLQ/7GItx3tKst8nhuXCgyeY3jRKcCJOgA1uIkUERg
LuNMK/xZzCoAEO2+yqsWLmcrUei4EpyPZADhFqW1bQ7l/WhogaVIYQLzP/vjsSsZMPh6UBTXyluV
jvwnlsGG2YWw1QhPVpaQ2IPe0Sb9KDQFtJ6vAb29jsBRV8nYCoS9aVXKQZE65sbIpFCuDltktFeL
EndQh4AlPzu9b6TP2HlmSBPnOQLllCyaHGbEkQ4xIr9SlqkLVbJdM8suKLbcLStYgSDTmQZ0SZlw
A+fukQhU+WwGIkJv4by29q6inAkZtauLF52bLiRaPaEuMplpP8mn6JAWG9L/Iwu4Ogc8aNKC+hGi
Io4ifHYLhZdH9RfnsTxenbVWQB7hYuaMeHNcMoSinAUS85a1USyHDYRpk7Hfv0AZapIG1KAExN/Z
DgtVze/1iXZvQQU39EQTcTZuvv6yxgZ62GTvfHn0wU3G/7w0qdzdN5Xh5lNLN6FSMigfZ0nOXmnP
sUyhFdcV+lSL2RDbkXUfT/z73zekezRzkorAjxQ3levqFvdn+zsEGxt3HFuquxusboi15ytaCDMm
hf5jgA7cYBiGJJfbENu7U14IkyTkd6B9z5H/iL0QnfyR+FaM/AfvTTeDYmP5U9EVbhporBH6+/lE
OJ2K+6d2TjasOsZGW6anUf0cmeNq9vYf4XeCGC3PYDcoYIjr07P+5NuaVma/444nJVwKnJ4F3+/d
8D13tqt1cRjnUVZdZ9dsQtAr21142geee/1KoEXpM0a19h66RJYoE1iYBdJjvLc6D++1seyuV4T2
Dz3UvmMA8LxM9FvTfNKppeH28Mh4isIrTVOe1FPU9aY1OgELGJZDka+fYhqToOhMZjoOoJs03Ldk
WAAA1wzcWehBtbmJDQ0YOLZxa94gUuMG4fuzAc9Av9DSMKJPa2PbN8yyy6VW+P27VMLLkjchsRZh
1SgBtk/vAop/eEV3Q9G3l6fBIMLr5X5xMgnpOJNEx/xExajvpahwaEbkiEOpvRntHZgm+TyN6Aog
il2EdFEVzsc76SNdaMd4rihTOP8ZJB5uuwR6RblqpH3C84GheSZH6QDJjOkHEbKgN68qnzfC+URY
OdZqJX54ISN20ht71P3/7rYcDmbSbOt5zyJuFqN8MLBQQPWy6fKCB8yKV00Ien3Tv2X0Ytt8iQ3e
RQG1FWU0d4PjOujr4ETL1hbg9W1y1sQdtJnvCv/eY/39C27glQaTM4TTiLmNqn4nh7ZohxZ3LT8F
d2Nfw0uWlvATt3MoY75pgUEthJs49ZXcjJpcAHiLEfR14UWUF/eKbVIo6NeY9glTJ2h+ZUA29eYx
z5b28EO2d5Z/M+jSD23XiOLQeaytt08c6sQ98myrFS5WDxR4pqlyCYkDoAlHnqqEI8PgFN7pEytY
WsIR3B/jaEY0fZzjv4rhsb/cEoFgzLqTOe3Pfh6QiC5qKLsYM1UYHrSDyb5AFDIh42U/YicrCohv
E3UMK96DL5XL2beYpmrPz/SLim28UJvp4/g1ldBzIl/StzpUV/J/Xc0HI8kCrCx1TQR3wN0iPAtU
xtB8zp4DssaODFJwaxLED70CWZbzic9H6vKppcA0+sW97KU8w3uqnnHWvv5CEMerGr6cPPY5zae1
97Y5Vu7ZalNzg9Mj2H47WsC7ixWniblg8Xh6P3UrDcO4qv840k1JWXP+E+iu3dxluEkG2ROfRlQ+
ekmZ0t8rB1Ad7sNq/181N+1Ke2vVMIL4INzFZkrY22DKpod9Gv4HXIXkxKvJsv7ftpFo12gJPQmP
VJ75fl/H26Tvl3RkkJUDWMB45KJysg0pRlvuVzJJNiKjau1qGmhPh5VYjFY05iYB5cdrqhgvCY0S
xDytJdYIxWoyT/veFv66NxNgqg/XUzSdzZuHgjmyXwpzv5a/J70aGHphogTlSGEVx9lOFC60mtF0
fWL5SYvlWtzNmjlPm9+rs1HvvWQpCzsd0UUbwPhCRrcQtMx68AZBhBJ87Lo1OIpNvCwQX+p3y9Y7
XpsTbIu9kb/704ELTqdTb9+Kl6zRNfg7TTckFFTMdGYKlnlRXvwRFIAse1ew2LmbPNFEuh60/Agx
fzE8BfzqcphQH2G9DdpmPbu7PbGJ9neVWgwKsUMrafbePlrcaC38CI3bbG22UiUXvk3rGNjtrJ1V
OlVRPALrzWvvc9ayG1YUaqn6HxgT1t+ny7lYzvJ+j3pGTHBbThJKiayGExkehDofiKUwdTU+kIlp
/qg4VKPZDdjhz7NGVeHWTkB7LfbQiJekhCepLKH37jxDc3AiZfKb8m1I4FcdSa1Do88v8HiCiBUj
Bezxo5mqSRpnF5XGz1ToqIrkMmiWZSX44QfdfAZVJ05SSGDcIB+IE8yHD8x9GiQoVOflkCWi61d/
/zWItsIxFbiLqJmA5yII89cKr8Edt1d2i9wejC+lX8aMyThyDV/71a+zW5AsjUIC/Dq/yRXa9DUK
46ffH7nH8P9vvj0PDDtGDyjCxmjzKB/GPzrQRR6Sxsk6ePUOwFdhd78ztFWMx9kyCmJqUUWrPXdC
dVx1GgFscYR0NHL+3yQmfFzjj+JNEtpw5tkfMZoxdszPdaXU+gzhDMy+Rx9bjs6XjGGrgrHumNMJ
FFhJxFx1hFxY5X6pBoaOGH5IOL7iztSmFqYJYTrTvpt2r+6xUHrL56khRWizat33Tt6sOJEUk3ij
ylnKMVKMmCXbzbb3TIOCrHQidh4A9YUHyho5gakf7qp9xqP8ws1hHcM0b6GLLSkk1nxPLOhzOb79
Nmz5YOQzv3DhD4+RyWiE/ZqI4mBhUH9K3hzNPfnzqYITKSh3Ytz++U0Q5eenYF47LGsMwH8lHPRA
zMKfPdi/c3gg9KAU/yHY1Bx7sq5mznHi2Zbb3SJZ5Z+13xjLN5eVOMnlOGLooxqURDez90viJHAb
JICnn0BffU8Hm8sj0a1Nxdcv8sqZSbDAmGy1t9u0aMYIkDSyGH63cJ7aq8cSprygB7/ILGyr2BED
POsRTRIwZOMzzh38HML3DJXzdHEPSt9iu8Ad7mNJcDTb1L1+W1ptuX1mFFahB9kiXPV8wwRw/rF1
iW59oa+ao6wZLHpf1o6ihOMD4gvICz+GVFHD2o28to+JChv4diqXo5kyiPuncHqkjBJ2ADnjdEzY
gWicIHtTOOQU9vxX48OCsH//nWhm7MtxMb1nyDlOaNU+mCL9CWiNnbW/ojJtdYWkp9GD1/q+Ja5D
F+ny+vCeoY2v13xB2bFZaPO5ROMPUOBxTgkOzwHtvUNWKh4BzuS+PdmVDJWQ9kmAuM1qpD7REgS1
liBBTs7/s+2chK+HTqY5+xyLnsk+et9tHZhyVcjG3ymLjCAhTGBBNpCXBeURpKns+1hpC4NwM2P1
marmatUUFT89SqFCIf4I/Boz7xL8I/JRVRYJ/aSHRuR2Q5QXyINwIukudZSbUK5vuqJtmetkgy1P
RNGQDV4o/ec0Qj4WgLthI6ieAus+xrfmrZzAIi7iBFpZcF3E8apU6m5hxAP3AV9mrGkRL+R1ABnR
+8hexLzwG5fCrogolECzEEWyVXJUir7Pi1sfiT6oJ1sLlmZjZyCsKGO5GmiyAJkg2yWMdkxMAShC
RFUnydGvGu2ToNGhKy68jZMuxr+vGei3qRTNfIjiM3XosiK1JpNfVxBglNBoI2ogwrOeg+OkS/v+
8Ifv7rFH176zb9AzVg32R+QDS0jzk+ElFbILPh5N3nPNtnjtlCvg1cy4gBLAlFs5Q77mJEklL2ZF
Atd7KOmWDySLcCcTWiGngEJ0A5z6xErKSri/7CizgreiFaNZ6XyArUjGgDFKYxeBhSTXofkFaI3G
OETf8Y8RyD4XoPah/1dzt/bG9q18egKaWLrtAkVghFtJuaPbCG4qGdmwO70coUw8tVzDZGpcCeyO
uk/dak+CK2q5GcMuw5Ovdb2Nk1+7xkxBk8H/7NWp1toucfYbmIhY7Rk3+Poh9uGeko/ZLmfo+OCQ
Vp+k2igQNWWD46/AyCCzqpqoH7dsZfcy7Ro1UPgHTjeA75yxUwhgvqa5lCbJbu4yAy9ALGMrZbI/
iwl+F+Kcy9OqLr4AhYjM6EmfrKkp/1OVMabVZqV3aOkqCM/OMN1BGbK95yJXPzICtFxwYAYQNlfW
PeqbpOfUB8yEx/jW37Iwpt6j2KA6yx8sZkSrR/fAt3bKdO0qOxhZkbg+Q07ooycwMhR6LO3OcGjG
LLh1sEsd3qiG7jhgzDTsgDpt2KP7xMgBUVFbHNqIADAj6h0fv041b6a+z+7p67kmwNBDqRqLutlD
3Vnv8MYIzoy2IZpaTYD80bg6FNkL2zebkGQpeXzzgKL6P3MNs7QK5lj7HpDHI+uKe5/v15U3njPw
ywwMyAuj4ZeSTyE/fVK9TnTFNTDklqpPIZjSnp1/GbdF8jZg4KwhcInOkxtnzhS1KFXgl9g7eR3j
9jxw5ve7JnvCbImMaE0uTigAJGCYIYhch57dod2EvVhbLB1PC/RJATuII53yjyKxto9Pscmp6Eo8
mwpCYWm+4CS+SJ7goRp6eEnbUrBJ9uvACc4ezqMCcfcg12lLkxLdUG2iN6giL/Mt9NfUZXJIMf7M
iETxPYILlTeaA13LI8gRhL7cx9uDT4x3htqKh3MDhXQrogACcreV0ZVt+7VZV6B8wKY8mq4fubRG
7vFmIa8fQ1FWotf/PV0WAZ8VuQnVXh2pMh8wImB4VTUlWgJJPGPkpu5gS9a1m5Jc4kKotSAf/UNt
eEstRIu8tozu2Oe8CLEaCzDKx4aZeefSS8oSD52zBB5Rs+5JhoO1kK0Od6PyHrtumZ/lqp7iJkIU
ZRvdDcPE1sdKQcxlMPeHGB5EbndbmS2oC/u8H1OrPCXt+AX+c8dC5/DXCUUX+PA2N/oK+pfbR+dV
d1kg1fvdX/Ptld+cxvt+/Kz64CW1TfhGwn31booJ+pwLLo8wAvV8ogXoc6+U5FwTFktpsbKhsbHA
ZuzTvEyfGNWiCDYDa7dqpdowaHDCiSPycdsssrFM7/k+iJVYnvgnBaAxKrLawJak9cRe7ilb4z0C
9/Vse0vnq1h41lE69Wv0eQsEEtsUo8snu73oXotVnTGNud5PNEu/8B+H34yjczW5vSP0wFRSN0rp
LDXUg1GL3JN5Zgrt8t8GFvmckO58z3dnW1o0Kobq6rLgal58b+yhiQzxdPzmY/dl09fnp29SbIsu
7aeTFrO0jYfUECWc9g+LziskvYwYND6T2YJi9KWv4lZuFDM6/tM5xR5fwcczD37XjP9YcdYJCBNE
jnLBQgeJ0eF8vgYqJ5YeFcW29Xq/MVnwoezjjwCN1BaGXSZrV59pExfb8Aqz4z2mB9vzXB+y6JcA
vCIqfrrI/2I+D8bJwn8qQgnMVQkdDe4wkK44zr/JZqb1XUTiahycDhYAAlCJ6QdVxSlvV7Tr1Sdb
YJqGSjXnU7LS1FUBXIh7GSjCUbWhopz6iH/feia0DbF4H9Yx0b9NBJIOPeMhB4MnE035U6huSuSe
8mNP6n7Ii7afDBw4cyr5gS2aj40AzBVHpK6DahBCFGNfr1wFuTOQZYf0fEqwsfKxmMcEPwoyCKwR
cn4L4FxQJLOG9WELHk9c8eIScpTWiFCjjDagnOkYIFbkjmZojNwsi/FruwYNKllrlrSAjB+bwX2B
xm+XODTBp5EeTiMP0oOCqTtzIYD7YWF9VlSqTk4AzygZg8UJ9sSF3j0GSKeP2jrWFwg63mpNQZo5
vJdiLkwePFToMma+F2SNNwBgmgroHC2cgiN0GFJyt7R61A1v4gIQvpp00j2yRA/81FipiXfhCHAd
j4kmUuastH42gUq65umSei6fJJO3SFwsdfaCfvdBOHSJz61PBCxKvtTXYJ+mm0KoSuj2/AXiPg8m
FkBxiwWzh5q+cZC4FpNUyTnmLVIXwSz4IQ0l6qEK4ch7E2uXrsW1uLz5WZuLdrz/4tHB3+KReVL/
a9BYyjnjNadwYuwnH+MsTV9mafXnmSruRNAFt2dHJfS6iX3WZnfp1CDBCsk2KWI7Jow8dxC1PsX2
u66RcUwy+wxGnGZBdvDOd5vCQ4OD5gkKA3KuPZfAkPRi1u9iu1FTUjoV2/K1VS5zBLdEUcSRKpn7
N3rA0ztyVCUEd3z7VKymLMedJ1J7w6bBgtKap0TpiN4j9e9vuV2tCr6qFHcr61CPLpBzAhGN3Iof
h7LA9d1zepoDiJsChp7K15tRugg3R2iY5pVMgsv5GWSsyshWNkcaWcBMRwe44GUgV2x/596F6GkV
WCFo/dHx+NqOyt4qyxo1Rywc8UqAFec7W1Lyo2Z8U8RNYUzL6EURp7fyaLJKkkzig+oYosJPpsRz
litamvVgMj/1YAFEaMgxOVRm1zFurdoSNAwD6/J6C6od/qF8aG/pRtrzZfzhacXD4iimrO0Tdr8d
cX9ZAIk0+sQ42E+KgZKAdvZ6eynDBkFQ6EzdikdMhcAdEykWofNv/f80d/nnLV6Oc6p4stdN+SG5
pXygmZL8wQI6OjdxEuzb9mgZ5jIQmsNS3PKOEKQXuHDbTUpHQYVkGviBeeyAYk5DEdYbU7jznEv1
gTyddb4xE1G4r7T/sAf+fi5CKJL8vj3XsSRtcjT4y/vpEqO88XWqBbGl/MVWNloPcAxehw7qOM07
KkmP6O23KvWwT0mMwLSQ4QqCDW57uHl+UgsmgPJDfJgAq1g5XDcIYkvkmhfyM+KYE8q8yQIny2lV
J9pvSjneP1KqKLkFocXZBh35ZbFFZr71SSMncEBbeEPpOPfTCRqdEpPgyoHeAnRcIZqQ+6p4u3D2
A5ewTqfYerSXusQ93lpfVS+RMb5k9vFnDVspxpNrd9mRt7ylk+WybPtyPFmv9LB8XsqVgyNfiS3x
XgYrHDMQlCYx9RpCwF2NaQD1HvOCgb1flWwi3tkYHoemKSZCHOKglD92tF/aDUVIFx7yS+VJb1we
ssC811OlynIkVbp37APXBsjEazs0vhjbOAlvO9QgdseuAslTzZfh+hIiKvA428MGfuzLi+hVMUaJ
1LbVzPq5pEe8Z6Bhf5XJCFB6q2wd97Q7CdMf2I0c6zO3ijchwpIqIC6WZvLbUTZ1B2VQsqFJQn3+
A1KcBxzJKOrLkZHo1VpJ8RpJ8H8DkJyNX2tWOOoO1WRKYNHZM576GbAVtmdX/VFicDCHCJ+FuAQc
oGJYR2gOuKJ3HS7WFb3rATil6AwPwuH7xWu1LRp2koz7gMNkEZMEo1cr7se+CWUHpemqaqZu5kIm
YvJHRUHaytcrSG14rnbAzaHZs5BYdoaWGKU65Z6ihrmYRADTzwOhFanhYRDRaDUWSMCiPZTSLW+6
otTXbr0XCwlfnIwzFXMwc4uI4UR2OQRQPtPgqWrfelxXpfCcFNM8Lcv6wCxKwoTP3A3ABQW8L9YB
5+3eKicemb6lIpRKCXGrncKK/Bj60QcrCYGLS+KNrPBvNldkT8MFd3YaWVD860HGZOtUGKuf6BG8
2dqrTR3+/aeUUQ2KO3J5TFWXsVCRC3YnDRV9fqcfE+1ma7Uj/HLuG1EV0QNX4BwPFovfjyHK0QX0
w7RRiOZhxvn8JVAT3pjinWZ6FbmRbqc4esF1vlDJUNHsEUmNyOtAzWUds79MvT/BV8mwcMV84sm+
NfHf7txl390V4Fcir4Ss7MREdWlHeMWJKKQ6n1G8z+hCgy8hMk2iOD3z+sjAdwpyk5KIrdHAL4q5
T/ROY2z029dQrdfFwaPe5FZQC9439wculqdgvSsmV7eb3TNzKLDwiKBFiZQ8mvX7p1uj6DxZQOMG
e7VAsVDmKjbLOAFoUhBCuXTHgBi0+M+Zc6w9XCx2Ku8g54eVY8apNVb/SARS8QJFc1uFZmp5QFVK
VIwN45nbV6Q4Nr0y9hGz96kHr6/3IsyHFg+8KvTjUdW5yjBWGEF2Hocj+/nlPcQ4/gpENm9vfTOx
RKr4GHdA4JHjEBzOvzwcIvtvJf7YkIp5eFhjv2SxZ9cZnXpmZ5YjQMONwJ5EATjpoy4qsxHYwLxh
LxVqR698VBdgEj8r30yXFwWY8Otp5Gz0TuDdA3zCVLnGMVki3/wd8IEKhm6yd8TOC03kQiGxJqwb
UqQ4ZkxpOUA3SUw+HEaq8OaFZFVx9Vh+R3zURu6ftyl4uuU+bOYv3jfsJswY0LcLTWlQdW+OBJrs
YF/sh7CT8PrzfrfozInhBR5zT2UqY5gjWUeNycM9nU5O1YAxy183G9dDFH39VObZogi+Ghm3opDb
JHeHLfpIzH5sqcnUuMwbaSm30GR/Rukq3IrWLS5jjmP1cUb4M1wYIwMEzU/53o/o/1S9FYnkeLp3
G62ho02NSB+2y7UO0uAYozsxG3pR34EjxJIlm8U09mU64C4H7qZUTs7bE/I8twgVsOptvwgNZ/bD
/XCiZNQ9RlRJiwe3ALJ+AKMKRo23zsbTysCb6nCWZTKAsyDLgXqrMN+OG8sWTeJiAP0FIGaaVB8c
EUXenvJC2TwL6iAiBZ1jSrkHoymEHTz37RkvrHyHoL0MNAP5E37xusITXRBwB7JwBtlGjPsbJSsz
eBjFCZybuG1zHiBxkXxkDPenNK81dsJ4g2cbSBnltbXwo+dBn7eFWiFTJq6fhu8D6kPdmvRWwUOo
AVXMxiCZwbOixwKlODWAvYMeGgwUJE52edFCje0bfzGnSHts72Nxx8LrR0xPP1S9xYeOefM0UvJq
itDATSiLl7qAJ++7luzTYUuxYbSkiNpwwkIrfodNk1CiZJlksDdcgCILpzPsqys4xuj8X12M+FPx
UWI3PbPFusjHV3J29KqQV7jE253AwGZIo9yUb2N4Grf4dpRgR7NYJPvxH1pAzJIsADetZYoS0qzz
m+JILcC83Q8HkF/YaqUm4m0Sfy7wY3ZbsIVwSxcm1raDexBCqClSzsnoL8yPfeJIJCs7mCb++T2n
GbI5l1osj/fkEELbBqOxl4rshYZg3Gx+cSab5krthGKdEjEJ53+NXIci2E5palXRAaSLMbiZaFAe
htYlEum8p5/zu/N6J1ZZqQ+3K7ckxFeLMrhJapF6gSZXpPp1FOdG7/S24l+vJpEZlvRxsubyC0ei
MYt06hHiHNZbtxMAymgvP0/bPAxrYMgbQzA8Fi/mtmtG1A4gpp0pfAynRmNu11F6P9WgbaONqN7f
x+hTLPj9hFWDgEvA80zDgLJyvjVkK4cX7wLes+dCIss7/7MSCb2Fu/24VnrSH3onfQkue3kNXKj6
pdHPhYR+JUBO3Mj0zueujmigmrW2N9D4dH6EximxjkId+i7ny3V5hzpTn0xhaLnHrTqyKM3HDf6s
4/0EVLlRHz0P2khw2nsDAc7YDGCK8mRjsD0s1buuZXZwNHH6D+q9Rk3N+2K2yG5TpZrSNHTiG4qo
ampDrOJMV7xqlYeN4Q4bePCNtEs1qwpJQeAYLGmXSIFtP9vXGA48od+gHVYPub3BkRMk/JGxhaKo
llwW0clNhNHN2h9FkGomAEoAdHF3ctIk2AV0BVJvc4Cl2SNfFVA2k8nvupUtYO4Kkl9aZuvQP1uI
gH73wc9RcYJw88xMBkLbTu7wHqV+CHcX6l7TA/vLIL+gDK7+1Vqu3Jz4ycSJhvXV8Z7jbw+yxhYR
ZVyerfynICr0CNvMjpncf+LOD94jbvpAImxejZCxCn6IHOCeDhaxKOfsu6QAbuYuR4f+y4l67MmT
sxoIgtwGFR3wyHs7vpF/Mwte10SRK0LPIgyOpeXr/U/Iz/U4eGsjPBT5TKJvUxqnq2e9ZWAIJKBX
t3xfpAmUVB1aFKKGI+VuSCOAe7DakRYI+VBKUQtCtz3nHIsVQpBx7+ukBI6Qho3naRORmS/WAUWh
L/JjgMFJTZ9/g6f645QBcqp4BSqdAVtAFfgN7ZFJXBQuj/6fZZxrCo/DxlZtPyv5kMVHTqDPGgTh
bQ4mc2dpQDTPaPE34cnaCNiaFUd5LWPmXodJef5dwxjngJd2WVBCCsbG2luUJGTzN/ChzA1JfaXR
Mv1Mlyh/wwNOD1N0MPs2FYbkqjKqkakBGJXQa6Yh4iZBdTU2OZiCF54kypsTimZX2Ue1VNT0uSEe
wyxi32TChk/QhFeC1Mc/L2KTLdjYLBGrHZQSDCztWWgI0Cy7eUnJ8VPgBMZjj+bLRAUsAOIzqMIb
s63b0lX1MiNrC0e8DJH0pwATJc+P8rMkHfaa2HQLCv4KxrJXzN1kyTFuqhLeEzo59PxuFdB2n5nR
iv1Jq3zxcBlP/t53e3vxV148GsFXXuMvjlWJuApqnpf7fz0+dsiP3vIvmIOgzuVpKtPmgIxesnLf
ivCXWJYK6j7n4XUIfrRY5QXqsa+Wbtb+wYQ/NrVzdxbvmKR/8g0UPzE2ch+FV3WBUrEsyyHXUMQD
VAkBOWhFZMFSB4/1I6gpDCtR44iB8E71PLYSQ5UDIZrSZX1TF3EfcmH9qO37EGKY+KSW2s8x6DcO
fWr5csPn7OqpP2H8kvSXjd7JCH0g1N3MQYSaFmwc89R0x5LrHD4t3vVZd5lQHk/pMWuxhrFr1D9g
2KJiZm0nZD0InrV1Y+eClUzOKpsyPZtxe2x3YlDMoWCcQfMs2IlrEEgkvYND/7sodf3hKqj8PYs8
aXHLUExhMEWrvNg0fOKjATXOp9mBVw3lga5jj2GiGJpTZvGHOOSYkv9f+dFRE76JJuniw9oSBDL+
G+WCfn/X2P+9vTvp7BK3UN7wRUlydAMIFo4eWHCIgVfUt+WaWWRedLFCs4NXurq9Dl4MSj+U+rD/
n5NcubBQF4vc/DryJp0WyD7cUFm+swQWZD27eQk42PLqHmV91wBwD7P0H++pf8Ssr5I2JdSDSH17
SnEjYzelUA0T3M2F12CMn1NtxCF2rSOKNylDS7z0hKLQ4vD2R+3OLSG0lz780xuEnF2zZc2dTdok
7OQQ53luUhfhpNfRBtOJWvqLw8Q/UVO+cZQAErFs2d3Wk5vlaya2wX4AvrsaUytSvFooHNnkHGwU
qsNUAKaMNYpeief6H/IN5ga9oK/49ktgMqPeDakGaqwc5b10A6rTNqMcD5idYOCCmdHT1d6yhfbH
hGFeghG5ENEiSiFkf2pHuFNgovqLs7BfmWQ8yEizrTJ78ltklPcG5yr9nXUPtv+Ae9vwAX+ZRAuL
1icz7AA5uvULUFC9YrKAoCrsNnfglDLIoCFI47SWO4ot/qDtRI/+5iY+D8jnjlTvOQkiBDoTgk+O
KPqpICiKH3QV4FM37WPRVAfp/zrqlQXs1eGeuNHaHbnbtRCRq4JJTKz8Rrgf5ToVlUToh69n03wL
Ru8aPEfSUz0pEKrFv22BklKlY+hrqBIdJPpKHJwWHT5rAh0h2LesuM8u3RyarZVxpsYCkWvaycRS
v2iyRw/olQdq6HYkKQQId0xYeKOYjuTQyX92TNwv02fNahiOWDmMubpVU+R1xDX6V7cxUNZSZHbn
5nVogRPBvfT78eb/mY9slyH1mOe1opk10HgAwS2CmMxnLsEIh2VWDrlt6p8jWnIrr66WV8rKniwb
UgtuWzV1JQF0H15vEZSelSihYeYBCYdHBdSUZyGLsCiiPWIn4X5u2Vx8nQMoItfsJ5B8tggBDvqh
9A8Et3L/IToocuveb6AMza5oIpJA77/xIwSMXi+x1u5e7wFaz+Jy7/+UpatXXekkAnaSllMVzB8K
k0bevaxQdfemJGq65i4K/IWD8g7uMzQS8FM1vR8OOQ1temrg1CAh+mpzXSllSTyrNkS+HnzOcIkR
VS3rUW7smK8eQKcduLhHpKouM7r8tfvFBBKHcyws96TZXuGe4MjGppmhkO9rZiN7HUIFoSgaJk3Z
uN8qRMmV5HqjvTRBuDErSE0gleHcoBLI3Kpd5tFv3jllKdmT1sUibbYBSiDnGskP82lpzguTKkUt
PrEZOemImcSmTh+fHzkngsSP1WfPClfD8vR3TsjtbotnxBj/mVGxLh1z+0ao2tlZfG2izWqUPKqk
o6bsNhOKfTRqZCyM1MRIlgcbETlAkX7FRZpP8iLggnbHNVYMw54Q9qqi1Py1xwL0jGqgxT/ZpIoV
8H/QvLG/rNyxTp+fCErxPKnI/iO+HpfmJkj+XSFp9A4a7pUdz4/ywUZad+mxMbpSP0M4Sq7mXAi1
JjDSjczV9lyHDMDTqDw+gy/Ybsm/tLXBd0hNG90u+ZqVTZ/mE3BNfNxB9KBW3DbJnDRhqUyY4Bl6
bTf1PGSg7KvSdxrQVe5/j7iQezXSY1NDNDJdM68Wkbo2SwVbztB0JyeksjkOjcDLdJWtAm39H1Fv
MlA9WwXlZ1qkpLRaBYtr+gXW7kenZD4/Lo08foBbFD/XsiNnvXMgfd7diGZbAhQP6/p3k7WFwXGu
aq5ptChI1Tpz+HTAkw8HYzMUJg8jAIsPrOWNK5LI2ZwR337qPxAkFBx+GvRQlbZwIooqDuk2dw8M
agskAlzY6qstsvXjITgrm+CLMhkMjSix2nk7T+aVghIwdrDYRNL9EFCa31P9TKAeiCAuUquOFI7C
es0sX33oEqcxo7QUSEAxWWwaK2u1Vv/ZZz/z5/jXSVRQ7iZ8dpNi9T17MoK6K0Pg1VrPqUj4wARJ
HJbgVIjuRjuB6F4QcbY9FosCBxOk6WNQm2N336uRhiJ97np2pOTg4LCiXrbauT/V+mP9g5atLBfY
855Zm0ivGftuW/6oOlZ2FymoQpIo9ZFfwhEVk6z7O59BIDCMN+f7QX9p6OVJ64a+fLMkoqSUPkjO
E0QmaZzA9BQK2e/fPjH20mMFp0gV+vHkD7TjJajJ+pipXh2vVl0ymogk++XTtIaiy59ISaqRB+hN
IagU+bbbTMNfKsyw597xe3zZMgSCoRjH5de5QiQeETEDgII232HCzW65sqy6n4RbkdZiKszVtgzb
d8/G8CO1CCoz6XaUrTFEYuxWmQti6EZ2ExEsLjVKsrBQdUKO4cv0kw43eB705+EC1tzUQUQlosAy
EL7Oo1hz0bO5GZ9ESYCl0G7Cas4QR2C6+F/80WUyePlcTLHX5P3KpGay5N7Grh+C1Wpjdhc3hDX0
xY9YTxujA6L9xlTudelSuRU9U4IvXbOi67Q3ami0rY3BE+d0hS+I5SoBOk5tJ94hBxxcQhwRAha9
yA3KGDMhlYxsTk3YvMgSTT5/vrni10Y0HfcFt2HlKCrs+qMaZiKwjd+VOxCjLuPtS6UXA2yx4CBo
BKZcHt9fWDrEhLg0YlFLC17cLZQIDoO3G446KgIGJPS01FNyKGQM0mtVWm/11+gFChRzn5irDda0
5QuFDEc3x4BYNXhDmSN6nJq5vHSd2/5GeCtIuS8Yq2Em0uau5AzGoWOBOG5hTuIpHMOyt1e2sQvD
NIH5rej6DGQlyUD1O+8kbTZGPD84vJS6rZkmGptW1tYcdti8URrp0rnFVTwbKUMe4u/v8hcFipVS
I32nnKozddhNZQdWAx5fLeIIn1n8P5khV1AicCZYes7MLe1pWX6cqxRuxgYXCh955fJMlSAq0d3W
noZ+euWX5SVBIpgs3LbA7y8+qlcnrGwgEyKIROHGQiowG0w2s/n3XfKHEo5J7zrKVSD60J0BOjXq
RTtBdZVvX/HZ3eUsIO+G5hm6StDOTtPFJIFrNLoyNOduzNZ2BWQBOogGCfvBiPKN/3ZGTgvrbs26
a9pOGbMSkopFkcA4zrmVOx4w8iVpV8DgxCPTB/mdx3xfpBpEP2Zy1yPkcUsxec7OPAyfXgvNTdUk
59vHBNUM06o93EaaitElaN7kdfQYS1aDNL31puCCQStyLyHWq+b3tJQtEDN9xmnsL1+hXHlz2FKP
2/SYRd1vKSbyAlqC5KHfmNtYcsyqeF1cuJCPOp75SY+rr3+rQnaC4hS9mLmvK+QTmiYbx4q76yUU
y2Vun40RTSgJaLMf8zoFsKfguiKf6uTj7ok7Lm3ORiP/SGtfRYohXS76H5thQYKHM2YD0XfClwvE
05x/agprpB/MKaY1WFmrfdksdgB2u+iAZk6z6YR3uMQv0EXogVkN4aoF9NNVfCTxVVOj6pe3CSl+
yKGeI7S4bo60vEm/poL/vqvLdF8B4KMLGDDGgSgrfwr7MFFu/zyRi11JKcKX9wGFp+ronUwSYk5u
fW+oT5cfqLPg0Gzu1g2A67kCTR4xkbdMP3z1hST/0YkvUiAakxcNT2NdXTJcCuiTvduHsLvBj4Kd
rBxZlKHr2mEPtjh591PQ6ZApMUrTuGq7Ioq0l1HiJnRBrO9CPfPb8k6eanR37T29Ol9fVMLsd489
ARUsKjj8ZGBoDP/so+DhnWvBYLyTj1EmGfvUiahp19pws474fD/z0qPX6hWltTpWs0v+uJ8X/T2J
3owVd4NfwvRYs09DPcftc2QygV9Rq9MxIaWO6EvPSP0+ktI4PvOQDYS3yTl2e190EOjGWB/Gudta
+eY2w9/upHWHwr3fmWOPQRDlkRM6r9IIBH6myYDlvEvgibu8LUYlbJqjmSgZ0r2uX6CjedOWnpz+
aLP2wJIUuLe6uIkUxGXQlrzIiJniss9RVNZTpDMdtnxEhan2mVva4+9XECFMgF/jqgJKOrhMfG+0
H1vWofAuZARpP9AA49478xYODY9Nh2EQCfQhEFstFz7n2601nbw4DFxi83ChjKTDi4XBN6PrbOgc
TYWchehv8asKy5grTb3isTP28TnzxZdu7enUMKkqui27U6paD1JE1rslF4KTR3n7PpDwZiVEsm7T
dIBDAGbPNhiL63NWD3u3IVRDgFZSKEYnw8Avw0sPPojnhiaDUdsSE791gtcL/wrKwm+LynJa/m0/
0Bd5W1wunWKCNpl+HMLJm71XUikojDklAK3JEobsdlPhV8lW6V4aoFer826uMKoKNRur3dS5SHn1
eXtfi4PJbqADmnzJt3KRcxnTnqCeUlfRR0zdP7vWstVgn4LLHuUcMiBXXlJSOyfLz7KnJ0TH1uVg
hRCOJepgZ2uON+3fTYVBkyc3vC1BqpEqOTR6vX/6gi4ki79lJVJULw6PqgpgDbjMUgvh9OrG0yl8
P2peSOwXDpkDnxLzoCEiBuU7/fKGmbR0H9tPRNZzHQtiq7wMB0Oj9Nv4H2EEjq6a5wMsut5AFmua
CQSaIs/M2Yo+n6mxya4V4yG26egkGh0IkcjdfX2DcVUhNEN4t2FbPkesCTWR9PCS4Vq3JycJ6fyh
COH6VQTWiOIqkUklCWyCsNEhcdgjjXNvTgW4gprhKxPv6wPyRYOz3lElwXVv8igWpH4jcB+PRQOX
e0CM+iGc15YRDSsL8Swcm8Gh0lmiv+z/Fy3lD/+uhW7zsEuYbK10o0DaF01TIqjl2VeKVWUVe7EM
v9QfMLD13FZC+zSqZgHGxJ9AV4TqKB5VR/uGR4ME4BWeD2TW60bVk+WJs6Lxa7oCfBhGxmZUy89S
IEeef5NTa/5WpV1TXfCGT/Hzx2Z6oSzZisuntU9pXYnNC3lwBXxCVv4qbJgJz4pybgazBl06pGXv
12TJi32EIWXdtAw93G+zu6ZZxHOq2uPghks+liDXMIY4yhkPYIAzMGah5TxsQvPE5YaGAxp/d5LM
bVMMj+4ZoYxaeKeRRkAiUJTQ0dvki0rvYFF2kplbYKOjB7LBS4yg2vkzQDfpLreyEPfqTlVg1sb4
oclS7pN8pawvn8ammGldMjQgkc/aaVqAzJoN0lUEpkSZOjNJYMEqyvjp+XklrbwFEvrFMuU4NMsm
22hCMbk8wLNZaMb82HHDh+gA5iAkxdbU0/U9mAhq58naBjyQXT9gQwB9En1qHAPpVBmBJXEyb2Gw
9szC5yPimGFard6PF1YaQu6BjJO/j2VCvpwgYjQLTnAiVUBD5qS44Ou+LfRToF5Wb/iXYhpvFzWI
1FmBMyJ8egV+GF1CnFy4y4YrdoRc1eXhLGyjWqJPTjUtFezupSv6rO4cDhf3yEpHZ5v4IJMXbE8X
Naxsjkva599y0piwDU9BGOhT2WwguMgYXqh3vPV+ytkSH61owvA9FL2yHB9+FKbYDJy9uSVJuyVU
tf3KpJJ97Gt000b27mmH7VqQJM7iZOn59ycg7IMkKTz22dJoG4mqIzx+zK+rSb+ayGPnQs/FBJEN
g0QRS+QWDMbRuD41ROOMEElgMLjiYYrDIoWVi+NFzPom0w+HuaFs/jhm/9gUUK3jvuMRZ1G88oWq
OI+fMYCATze4YsVRinuMybLMkroeK9DGk0pTaS36eSOlaq0uzx9xBQ4vfbOAl6k3gIyLgMxGLQfg
VJ3zptmi8kyirftfq2nbN7VAqBfVByYplecj5zjJrqoUCNoL2vf7FSXD4IOYaje/J/6ORXRV/GWA
9POnlmWrIqLjWgPjH/Guwg8JoCup78r7DS5brWgz+u5DLAorpSULJkfDoQdMUJFkJwhPRkM6ryVB
pJnqLoq7pZzqCJc8+dRMSIl2Ledug338H4Aceo81rC7tSJ4TXT2vXxXj694mAfKT2OSX85I4xBYg
YLQizHLbIcJt0GDOLiyEQhgxL8xKBRCaNnENA/a8Lo1mAlcTXt7Yn6HNKic1wMfAQjy4qR9hNVym
23964gDM4MXM+RAt4imvbxL9BZxqvrK5kAewS8cpN93WqLW2xaiPS8ocyCaJ4ROiGXaVajKv9BnT
txN2/pZhqnGf3V98W/56g1nwz2vN/6r0qeU9E37sVEQlg6BF/8a35qNJAsQ5WObpccS4iotoC0bK
dgbkkz8ZblxTFo8TbMndJmqXfEbROylaAGNW9tLjFifFxOKeNsdYmEacO3vzpCM61c9uDYkMuqpH
q/NSQaqGaPX5h9wBJV1Xi4tUqzyMFpZZSd/zIIyppXNv9/FRdSZtIGkou4exL279Yi0hiLe0NnT5
WoBBmxaRPCdutd3ceAXxjhuuKneStMP4UaC1c2r/dQxceiMd7XoZYEex5acWCexw3UVm7mzrd27L
UILTYZjrT3q4FaZdLxAYuoM9E7990fv3x4ZlOiVCWMIz86eSp02pDu4mqZFhuMSWBc0gIuWcapIi
OFGq6AlU8a1wxFNgZps1AGqecuQ0Hi6Tf7oHIwF8cG7OHh1fioAG0Ev2XDt7D+d69LF89TNYtJfg
28i36y+lJGJETSYsMe+5BYGJWJ8WWQlUYAoXiWgtfZTcvAjSGLh1sN/fmTpUUL9mhXZlBG+iN70H
cjhLIMa+dlP4Sn3raditu8J7diGp3ChpRwJ5FJpjdaANyUS6ZiOJe24GlUQSNLvmErRVVyynMApQ
0dhdSkqpfOShTUCaOwGNRi+QE3Mf/yZMV91771Ia1zdrv2xLuQKpfJVQRLEl90BlG+E91sqYNbaE
BRKU4U19NrpZVBakMWd6wanqISlf1xs286Kg5aJOmKMxb3fzgHM/kuoC3hI4SCYTN0TDJg+8+B9N
TnFp3hLcKctGlFV3AZ2bKdQ/JZv0Q7sLY8DjQjbsLER4S9NKVJ1kbtQtgvfGA76pj3o8NwcYWFfO
+W6qjJGnt0mcyUnBtO8RncGeqN7LWOtSmmM9z8sBPkMEnMn4v8GJeTQwQ3XtHS935Gf+QaQOlH6d
groRfHe8kFe23sLprk62aoMC/lzFqKdXMuXxy157XZVg68w8PVPdxuMsD8lOMe5WoycXKb3Nbe7z
UtugSWKBvEijtAWIRCAMv0hEvWYc3kQnjAYDm5Xb0PxG7hT395UvtLKYDCgXhf2cWsYE9VRkjV0s
1gGeduB9nJVSlBWjZx+wbLMxcWfLWXRqPVaJiovb3d3ba65ea+Q1Q8gt3qOQspAyNBFSISOSwyPq
AZyWZC9tCrUISvWYL+Zypk09VmQOfVUxS9H8WOWzv4HIqDY4Bqnoz3Ud1I/YN5CQtTs6Y1Y48XnT
GT0zgU9oxz5GKiBBrhgVZ7OzrKLPWiJKFZElwkTWG+EcUWxdlA9y05/74wxRVKEZ3XS5U2QP03ht
sqJ2frR1CxjoPiW3K3GSY4UconKPMU8T0h1VUyJNCK3+7FokqKnZyb/oceYHAp+aNO0G5sjHDz4O
JuxhIYVMbfvNlry6c7nk3bJYLDkZOUXBC2Ar/AkM4Q1cCiD2sOjv8eyg9OCXtNjysQkmSlG4vdSz
Pxb0WON1NjeT0vu0+tgztfeWQG+4QjH4LgFYmSBeNOpezi+LZ6vCjdcwMy1UxH4jbAt96M5b87A9
pBU+rkj1S6549fGBas3dFuI0HsJVsL+y+iEl9ULBgBRMD7X2QiqDvcFuOMi7ejhr3IKGCtdZLXMF
VnenbxBeF+6SqJqn4EZQNome+USmbfYRk65x9iVMcv744AOm44ztNuDq3WpafDe79ezJnzpBZznQ
wTsb9DEnELeibUKrC9Wb9AvMQxcm/CP1MQUjt5nH14p9qGtE/HzwrAaCMcmm5eRRGgdUbVMLvsIE
SvvUbzUz28/aZSFRH1J5q45Lz0nZHWgNHQRtHs/gsm6NQ6yce1guBLywo8o8ZS5elCZ7j0CBx8w3
2i+vbPRj7r1A4LBV9R7wOpD/YV9LfZacjOcuDR9icRMFsTzvSLVQffaKdmKV9Lub621+ydocJBIL
0Ix9hgpWTNTzRNHyTVMS0OhVl0QYbVpTLkOZWmlqy+yesotP41r0pIZBrG/MFIqCYewmBmsZ+SYp
9Z6HFA/8ZmNtv8ZtLZsxfUDI3wDx+eqDVArRASCxscvRkJx8PDesQTpn7k7H8uRjGWp1zkjBdPhS
4BVIPFQnFAYfJN+zDpQyZDBvGXYWIoAWiq34pz3h7YtQ8UAq54dF5nD3hTO8D8vgbZ6/A1mqUxeD
r6Z3ni+VEB8JuPQEo1G0dbHqp+I1sJamZmk6grTIUOJu2Gu/tzpYkZcfCBaRqfAG6JPcbKFZ8Q1F
D2SuKVkgbBqcNxCVBg2fqmmfv0eQUQ6C9CD/Immr9nnjFyokWTF7RIt5LGFJbBXZREKach6bY4uz
8TOBXZqLjwbvYQzKlkLhF1qsd7oQgvBUftiMEsDMB4MzxQakyZ6gKcoOUdjnJ5+f5BApQG/vCxNM
qCk/5aZ5jzQeyhKfCJDUPKI35FE37T8L3Vj74lwnl6oSQDyjvOTXKvR2I+FtsdrcB+mVl3CWGkf3
rv2XZns0xl6DGi9ja7BRW87dTvvhku5+fH5c0buQSi9TIeGoHsccnYfJsUUYiN2/yV2gcZ8etHxJ
vfjdgOrdfxnVstf6U04CWgC3tLub9kX2+69jtfxm2F0BSURTJ/+GVf3rT73qP/MXSCIoAnxcC/+d
b6xsrEPM2ssez+A2AiFyT4HbSy0QoeD+vrsw36RIGibHBRjw0jIG5UU35q2oSzDXQVSS+0hfa9rl
4DJyViyQ3d+qmVQJ/jXny91uq1vPWQcXRAlmr3jlA5dWNRo1/ueqG6b4/6XzQ7Ddc/dBcJeGwwT2
BsQkb1rcvHtSyv+cjVHMxgYS66Ph9PF+c/4hlMHUmN5y2+zw8mXwesjL/8uScdwluWgUX86RujmD
fwlH4IMiQMpF+kdJVaPACM64lgw7/sXkK+kJGePpK6iK2DzN14qxQFJb5Po4E6+SBCVwwo7GBk20
J/M9+ZWqk5NYFdnw7CnFKvMk296NlgqxRY31VB4NveImH+KnJrU7C0Pi+89no9OrQWbcolc8ALKx
DkWGqJbgqbbj4E+HujisT9riBoSqFVcHYFbnyUILrzAGF8yUbrAkkJgunTxFFqvrYttbdxGjGEz4
n+nQCyq+c/t57xWYzOiBRDwD3wkeZl5jUvca23vxojahmnTF8N8qQ8mEsY3lBqo2+gbJBs284Rda
4ibJUdd7jvdQVJA3RREoHXKs82jiiKFeypLxdGVKQLt6reIymjdhTW3lax+ac6mgX7z57okLmpUC
q6XTewuNk9aFBvggWeT/SNh129UBhvuNvOvpdbPiX+0vFboFLjdyloIdqC93QCCqPiKk7a81vjm/
f3lbioT5ZSulhp1D8I/X7lK7ZvCR9gAbGuk6jBMHk8SX3ZCaaS4SsHtqSZ+iu3w0vJBxb7bLvpU6
WSALjtirLhYH2jCygtgm9DaDZRJMRgn5aC+bMw7cakeBDuaQb53/sion3TH/ZmgcKZikZFXdTs45
HqGyl+ZHyVzQt0IzNlwLFAo782A/XohYULDam1GBgzY7wRlmfIWFPraO6JYcqx1AT/+/yi5Fq26o
9emg48JQXtjfJrdrwWllO/Tw02dIgWp2xlKAYS+mqPzLDMdOZw7TkuXurR1PxFWhd9UVCndw9dgp
Gdaq0NWkurpYO1MFklj+3PCXTZ7q/MzzjymdBAFHfI9wd0ZWnQ1t9JZo1RvVgNjZrY0/PTbSLZN3
NjuWnuf3kKLCUM6VIX2AmOGaK1IZe50VIvvrTV2MTGwK5/D7eOSDl1fxNYwvuZwvoKEbGhhDfuKx
la4EWyn1npM+m4jbnhw3QNe23gxTpFtAWXT07/TSZ6wVHfSgRFScqyr/X+eqvzlBq+MYz+7HvCQU
vw+m6p9tU7aC4x6pKDYdENNOKfz3L3N9tiVvCJWu1KBIIHMuYmCvsoQGW5C3AqxFTw67djUA0YZv
t/pPKWHZyCewwidBPEVnWYKsu9rl3kkVl+ZS3RJrXfh+yttgaehBIIc4oP3iSqw+BfpstcE3hvSY
9jMJgfS8KlsYJLeL6fuh/5o11l4yp3kV2/aZLyPu12pY0vwlbsIbQpq1G/V/L1s7F0NnUTXLD9eS
ra/hT4Khdnq/2KlGwFJv81oz67Il/XGafFdwK6ZW/fUVOudeOUBQQQ54Sl69bHc8P46/YuzyinjL
xjg7F4UCmYA5cROBnDJNBsxCGfX4wHmHNOzA4EkNRGYO7NpVdebnv83lTBGjAckZvznXC+EHF5wX
JFbBVoCsAPG9NCLs6ZlMBIB1maYcSm0J/OVwWuk+5V4utMxtcgea5xyJAwCuh9Y1J1yVXXpxIRd+
8jUw7eBWDgX1xmQJx/KsOCGNlQ4RdQ6bcyoo/1xsQFGFg+okwCfDuMMhA+T6TwhbDGp1JeI+XtMt
2s+VnvtTFuQR465r4BYuZTLj14GB0SoDXhwMbZBYTVSfm44lDdK5X72c5S4s99lV5nDX5+AlNgFd
u8tl5ejU+XBp6SxZ77XdQ/Pw2GwtojeGYQWG+NlySYnBQ9fesjitQuDIswRUJWM+UP8cjB2Ojznk
qn9I+hPDSW/jpv+PIEJ9kRHMAqduiy5+RA4X1Y++69A7Rr5xlCwceJqs9UmWBbAJcuYzbwD7dVrZ
uiQF8QjJkNQHA+sPD1mxE7HLTPMMkvw7YI5JZaduByFscty2zzMQujtgx1c92uYoV7w1WwEL2tTC
u4GgOW9jYCDIN351ULsEJQjV1L62E/wJjV32849OsqP+Q55RUA4dzuhcI6QNuYkkHA4BX0zWOWiu
Z1lHRaMJrl5ra443DpQ8T6wDbUPqMBriPVutyuJt94af+ZRlbcdDD+inaJtCkCXDH26WpQ9vpqJ9
mcx2LCtrXKAN5lJf6Z+VsM6FqjjNZ8hUB5b6bMr3w+0y8xaBqcAbieu8tvZES3OhDDLdqwJbnKPJ
j1gbBxmYfnsrGNgrsbWkZnLqHRvZt3O2TPgMG68BK43Lyrkv4L/2xkrkDP3DWTfEr+EJt7U2tlDw
TQYWo/Imi+O1PwBVCCGBt4htIbRhONbpkB/rDxQ1Vq1KklcylXAPn7/wc/x7kZ1wVi4TCG1YBvb/
T5N68349hSq+E8y5p4YzV9yBA4XPs/UjJTM8ojhDnQCyPPb60rm3LUffkMv8c6wMxtiEbSx2QXZC
qcMH8GKFT6yXDpEtGIVnR8TIWtdhfI9CtqK5uEYJj5RM8yHGKCNxkB43enyyeVvWuKmlY89pdZ3N
VFcv7ej02hWTjPzNLa50nDAEF5SC6dV3yVDach0oOxueoR6S/D+Nt3x3KvfsndgpAWXjuclfy+Xn
XRQySeZC6VZd1QgxpUXmFecMmaTHj3csrcQV6U9eP27dSUwKP0sQXorzpXgC1DA8eGRZEyR+nqoI
SMxDzM3KJLy5U7ekbTQpZDtTO0qeaGgwLHvytjUurRPf8QWftHURIOmw/MAdFLq7UDuoQYVGfN3I
K/ActGj1NdH/kIFXy+rIhr1SscjNOIKLXvL8AJ9RJb+KMeVLmiNVBzhEqwJz2hYxxGg3JzYhPkpF
yJTiMqz0I0hJz6JavU2UVP6RdCOI6RTH93+XzdhHDoIIHOfcQMLMPcpl871zXgJVyf3S1wHISk94
xxPq9nT0RVGqYKKd3Ru+J0t2zyErmz0aedG1ShLJoIWw6813SL1uQT1PV1SQKIcoYhji9S1UyxiA
pdKdaSOmZYY4qLkggAfo1ycFjXs0SvERFaRAo/F74Ay3cCqGLO561xcNS0iz4qPzLgrCOXWsfZWE
eqml02uNraN+g2sJ6hIRRLKuG1vegBhmU7uw5kQ/rBi3AC24ozwHXlq0FquthIWEqpkg76Z1yvp2
My+YVaVjMeR6yUNPzfQdUqv8OBhRvm/absqaJFeh4dR33NTuQd0FjKjtiK/GoldZ6oE5Qd8A1z/N
KIdFo37KR9EkVhKNP5oPRhb8PF3MbrPe95Cjn5+c5K33JTdWh9Q0DRUOoqS+gkdsqEekY7jmReQ0
JsnqbS9+QZhyFVBNqnHQ0CC3RA8VSacq2nh+BiJFpvR6zm8pLiwav2w+nrk3CG0913oja/0HFi75
/jwLfQ+vS3Kl2869SWsq7Wm4PGeNI/Cq5mBf9mrV8SgS3jNlLPsFgO+DApjP0+S0I365Y/qRyHZC
BOlLEAWVSSr0wMKq4Kkk7AnketOjkpIaraLRnxtLQVQH3+zBBWxOd56i57OTRMTANqZi+UBPi5Gu
uskJsaDhRUamgnKw0ZVg+vOfPIim/5kE3EslPiBQSJSEL5/ZJRPZ4675K+5V92Qgu9Arj7V3vYYL
Gaexuv5x8XtEGJMWFeR6+Kzi6O/4kH5R4RgQCDjv+KJ8NBAaFSQXyUGS3LWUfmJcCEHwqYJf+6zB
PiUOYe9Ae3YpvwVRCs3WnVk7PahR8kndFTQud75p1MMHvb/lPgcmQzxJuBVzeaqEypMYnWpmHzyO
neh0vnPoAbfSyr26jjRjCYbMUVbmiZdkWE1qdYUqgN24q8RSs11yzkb8mXEr3jfsoEGCZ3UPDn/y
IBh5wqaMmX8OCAIKymdspif1YxX4nH3PSS3qVhb6gzyJrxz1mcwufCf6l2X/nLwdfbrNYDjs9neD
N9b8h4TGcdh8tdUOqoFcB8mRO5+ZDz+kd41xjLxqDcv10buDULMgQyN/mOJbuFUz5E4YP0Fbk2SV
Hkaget9H+7EBIQD6JJaovBjF+OI7lGR5P2WFOv/ssS9vX1cT1bw0ZIXoqtt2dA5sjjp3gNhT6PLB
7ipix+aalpxfYomm4giJDZR4+EhLIHW59axjoiHNKFGQCogde/eMyTesmZ6N5YRmqZhwbJIvq7nj
aALVVZYq6BjDO610MG2ThpLB2FXC3tovEBixgLsQzOy9abv66cpgKa6Wz7Tn7HktNnJZwQURkDMK
yZhlbzS2KN5/FmCm7MRzTVjXF9+fi+lXo0NCSF6mw109iRz8Enx9UnK1NZVE4OKN0i4UiZfeakSx
3gTamLGwAfmkNd/JZWGI3dploYHROAsV9AhXv42U7RMIHK4FY3w4eulwhp7idUybfhFUucP7lrhJ
3yw/vJ1n0hxm3u13w55CtBPAhPv6fVWtUaKbnTVUY/5Re5VfsHz/XGrhu61SMyszpJvBKLfZepzu
eW3RIoiwxs4UpHSXFLY65o5vmd5ETHeDeUGmijOT5WBX1DlRUo0s9S1DyCWbXJ6ezlcBf0H/Gj68
cg/ctWgTCYaOy4I6+xzp5WHwM9U7PMaQ7s0guVOPwqzBrlKi2dBPotSAGf8MuwtADf7VEO77ADNN
AY+8drf+EOuwPCZBo27O6IgHrEn+iB3MImAbKF/q09kbj+hhUCRxm3BHT6BHWmCbQeNnGtdgkGie
C1jSh6bAiOdKPG8BuYuzDFamAaPUFl+Nww6NsRaBa1JfUVP1Gx+1aD2Y0iVc4YJ8PIKm3Qx4zAne
SSNFRV9WC5EvwIQJT28fqrEhAOY1CZC0D+olNRsVLqJ7gvICOzCy2gwAx8dtLAR8NASBsjhFWMyM
OMtFs68A3HhacoxzftgW8dW//WX7HBiUZZK0WEjnpV49pfkyh9rch0DIuD7XEgkUkYSkMWGipue8
Km4CBH+ILJukIQciI7YZhz4D3UDPF4Pg9Em5YvZKwtD3v2nF72i+vPg0NMNd224s6hHspPjLRJ3v
3v575IbQTRn/Bi/NUXxOx52035VtmQqmT2/IFR+n++MsM4SHEg2jiTbm0Ajyuq8oINohPhAx7Xvi
cCPtFt4kt5mWfMMIgjUYJbaEh9ALFBXHvH+Ci/3UB6R/lZl7RmySWP4jRgAmGTlIPPVm6Y60x2PW
EAA6DT4WTBmznFrJ9PUk3rf0CtSBe0Sl9kHfwXZGAtb4XgAwPpQl80PJRI5ousii8Fi6h+FRATmA
IA0r17p9iuj18uj9VsO3yo2XfN8a1ek8UX4qUOguFHn7N/rvE/f2VV1Y/T+sU4xVFnSY1QKEgHAF
aBpHp4Rik8dg5L6TYadzQOvfFyB9XJfsP/qc0cLNzSZ5gkThT7ivudFHJLJ5LTks2nNaSM4ICCLu
uCETh1a8IvxwqIHgrL1MLWzbFHYHgKKGxi8e+dJRLEZ5saGRll+RtGWivNze/rvC439/6WXP8Ohh
xoqZ9UM6fx46kokt4wsSFkdyrqPU8HFHbX5Ps2bduA6PAf4X/OCJmJL6vL9BY3hLX6KASbov1N8c
UJcN5UaBhep0WhpPMTcmSG6rzF3O4+ycaOkVbbu4anbCw3A6JwWWxC54dPYlLi3zdabihsa7OzvJ
tPGSauFMVCQk1vl/CcSRYxVnqibfgCBgF3ybGLaah3RdTcjTfjwhQMk50L52qfaRxV78ty8/uFd8
BoQHDWPbZl6vjLhoKpmvtunHv5vEqWbzUgpBTm8tfaAKpJDjC7IsY3n26dlutfiAZxL6U4rjO9xX
5jd1yWwH8SHJGtgbWGgj3bAOO/Mu4kHSnXseeVoi91caYpXyE1STs4N9uLGf10C9VS8HZbXPP+uZ
avKeYGNZljIc+OZkQRW0EITn8Pr/lerMQEzDbGoC1wA/2X/8+5slCnKHLAChLmTK++FzM1/LeJ3X
X52vLTl8c6XfU3OzXYqRDjjjUSUBSfiOPucBYbETM9yMJbPkXdw2JtLTSHENDUaBAd3lz9Pi+8Tk
18pLUhkY9BNC1HiZIdHA9QGTvLcDEkigzvHzSCaUY4vMq8UG9igmZBLSOOG5hk8WzusIoIuYdJlw
hpYhaccJexNWBEIRsrHA501btkAuZUyErMFOCZ9oS/CF3gcQbN6V2KSJPcFQPGL66hkfLsYh1C/X
rbG9CyvsteJ/WNX5NAauKcZWRfYBTWYEgS7425OpXpDLzoWIhoWy0YELVWO5v0aC9uUQs/+2LKfi
/1+Migha1eWFUhuWaIgQaSGxKTWj+AcYrbttYhgWi93jddeYFK8jUEg2Pf4LKryuq+mg2qa8x846
hAKDw7kE6JIt0c2496bxD1qMaSSMO7MSGHKhcXwsDHiwyAlhdAX7ylyKVi79dAiT0DH4OcHCDJlc
X6FyWJjxY4ucOm3WvB1g0Ml+h4MeinleXh9pFY1g8hgG6szIlUOJb82U1qQhsY/Ysmxipdi/ZwbO
9IY2RG5AaOFN9ipMVAGrtVRCopS38Kzrv2RbYELIukOmAcQCVfzrXDEHa0m/DxUW0s8LrdPXGnAt
hMKlASa/RRSvTc3/8kAs/L0LBUQcL5MYaM/BImOlyPO8VHZh2X69sCqrHyFPDw7GLaWsaLWSiKyC
rZ5Qn+dtD3bl20JA08oKodhLg9cQq6FwrFAbud+YAuND67n52RbEUVm0PwuSzaeVD5gB+uCxrDYG
puwiFDi/clcUsyVCfrNGy/5jvwuQbyt9snDy1PygfFEhDg8fWMQJ6EH6pdtkOlxb+6o1U0ZAl/+B
vnsRcYtm9VOVGtAp7dAhm26w9s7imCY7HfWXvDjiU/GatbluLw4gJjMV1bjG5MCKBaEFGcyCh8Xn
AJ8+clHPOx2o4i7BudzQEj5jbEwwHY5YIzEyuhZrqvOACo9bUaG8Jz/wvuf0F5gL+YbnUgH8iwF1
YgIootdzJtN6lr3S3qGNvZZUZW92eFNeyLZKBlrgdGnnKOaEIDDd5/qfE6H4tw7r1xwq5PLlozwR
2WNwNVerKpQ2z7y42u1XwaJt/SAh4FjMEeeZu5cAIdrY2BxYS3z0IXMftmNf/o06gN7oNlhftD2p
Fa6nM0l1X76ttmTVzzg/EbqlhSwyz2dCSVpw1Ihvs2d/j1nzab/lJE42ObjF9wCkieI/ht/77pgx
4VqysBkCvlRwmIFz3c8LBQHGbqjxkvn/syLVAC/RvN6ehzYjPtBrF6nQg+bV+JXnjP9qg4KKBT5W
2V1yUn22zD5Rh93laPdJUW7NbkfML9AvitWNRDpXZ5CzswifYS1Fp51ErUSBi5UZOpW+bQlxtTmQ
Ctf1hgYsv83BYF3AWMU+SGLEPFH13TvFS/OHRDG0pOkfl1KEgj0GzRoB7YH8GwyD94UrDv5Mzb/n
WWs1nz37hwpZhnJSYBBQfRyRMgXwD+IoyQIvi3EcBZL/pgTThic6MDJubLxyQUV44SEiXejaWyYX
cvjv1XuhcKeB7bWx3hzAnRVIJiKna6J+StBHOTNbLMQWsChKD+pNtIaF/CQDItmiGFXHpK0FC2h8
0mK1zPc/jMCn9lmlddkCRm05ObB8S7C+uY4OCkfo3cNrDcovuv8xTm0oa7STAUkaYPIiouNmlEWo
2Lg9SjQfNo6uAaBLvmT9FpT/NqL6km9X4RLIIWuoXc40NybOsguEJIMBhtJpqhpqgWTVO+rHEI89
R7/4jVS+ObR2NBBcJnXa5q5fuXeBiwnUCfrvXLw2bUpaX3O74iBQW6sXgLFEZZdFbuIz9CNbLn3v
c1q0AYRSmJajn8uPC0nwhsUDC54nw4ReKLgfeHRyJRQCtVU2gRTtniKkUj2EyCARZ4seRcvkzPN7
0DcJdVrunA0APLk5MAGaqs5xbgnWW90o9YBf+f28m4azafT+l+pZ7RqpeFK75D06rNvszhHRW/LX
k8enuz+L7Ox1m7uHxCihylRA6WnptrBqE2kX6bfiEDcxuebbeykky7c0cdbhiSe+9hv3cBVcOd2S
IvwrMwTHN5ESx9gcDO7wvcZCSeXW2JVs2IqJm5anKMkEchF09+giW3AAiKZ9oAYgo97lZJks4r+X
mD8eV94D82mdzTLkk3ZbL3fWgDpuGFpfIRHLmBriix9AtjPgovqYTFMsa8gyZPe2cbjcOVd6bVd0
vTboEEH68l9nP6MVogbWfXEOYqo8K/5wCOEiGKosIllB7Ate6eVKi45TC5w1dIRLIXg3ecieJPjG
HPddA7/u4QyYQkqGb+0GFksmjxMd506adjXavJ6Hoqlj9kogCI/4gk/Jis4CZarDhvEWgdyeZOTQ
m90tZQC5+g2xqyQXhqURV+phnrgye/tbuLdOg9MCmP/wgAnPXQhC8QGzZq5vA8c/bDqC8GvvMw6i
KedSGSZgWE5x5B2gDD5gBRY6YFK+VOuVSjpUQGzP0OFeydbAsV++D8TZpwAQoqtHTk6HaogASwQC
1lmrS2bA23hQRAsckhRWcHkQqD2jwXm4HDejXovTTlEnZjD9kRbS39YcJ45ym0KA0aUdaQgZKCdQ
rR2Nh1/1WqcsG6pXDGU9ObroA5InYDRDNLyAdwj+JoZEPclHhX42zMqDC514+GAOSBPuCpDolUJW
Czho3MatMJ/0RXy+fYqqKA1QpreaPasz7cEbWCLKizEfvBSW67AoBpTxYtxcv9NoBzaMXLAPTvhb
xYSoOtMx6lEEcmikr9zEU2ikANXkRUtcZ2Vu32anKQJMCyrzKGfkcuec45o4sSOm8LLjafP7nKOh
oXiaLu44YczoFwlRpJIXrDyS766K6rmKPa21uNIAEQxnRZAjRTmZftN5OTbg3f3UlcknpZSEuntd
rz/8lurZK4Olc0eD2HZEv94TYDOQIuS8GnXjI+tmU5MR1xMehbsodunIYGbR7RokhoFavhyNiqth
0uZUOi3FVg/h8GmB8YYNEAStZoniPzwOJgzTDGSrhE1e0QsPKPVIPceNZxcFxjwhwuTBAlonKmdq
crj6Be49DWMjqKlZPdVzT1h9MPg0TpySdzKlPiEg5zOg5DwewyUPiBbkSxm4S74uje0DR3QHUeO7
TaQVoX8Bed/YLELFA6xq6Bw98+B5XahmpyW0ib4zbnAM+VRlPWQAJoWYFb24jorRGChrL/UNHPpk
EObHhRoMwOB1p/rv82xYXVxemQObZUGJvm2POxfeopUXg0ULMb6cFftC0FYvB5QLnmaOYTj7Zx6U
fPQ8ifqfVA+kERMK50laV9TMAVQadXDMYDVPD1LY0EOM0+Qpu+osZw8q0IrWcIKERvpm0fng4opj
nxO8YHMS/U70g8SjsDktJOpkYxkCEGZYT9anPE101NSQ9jwAOo2gMO5YqRxOVxKPG5UgY0WtOhUV
S69GjUSaaj4YqsKhzBd1hPcKMHJG+dptT091gBistFuCvakds+XHXH/snZAjtZz9HHdSDM2gs40s
dHlhLRFSRMTGG+2eP4pMV5awtd/d15vbkws5NXUSnFMARzIoO/N8ePO4w0WRRkdPRI9UPePHaTqA
p7X1uA6iGNSuIPD1SI2K8O4UfJjoh19T5sd0otM0H4LAyanrHiPh2aN0hzSnUWB+x2FTB/KiT2Pg
mYJa9UBXGKKt0nnS8FlGMlqFzH2JsKrejaaBCeKitauqAWPRm0eb/fSY7BvzrsOI7rHCYzpMpWqe
3fKQYwinTWrw2pzaR1/y8al5hdKfEsOVHHzsDF6YzSd1FRo7ge2GSd0Pj56S4U9YauNihCaqIYsz
oMd5ww3pAo8J3Fh2qs6oJBwKHx59NanCoLUf0PzSRwpBhl/wwFnJnqKkcm5C4PzfHjnREyqYtitM
kxJjeNhh4zod+NHNVF0VKkY/PDX7AVi2AF8abenkXCBfpF+rcbeCYtBKH1bdnxxNXq06i6RS6sUk
DPkzJL+sOBZL6GozpUxvpWWKPrkTVg6V5RJqhJqMzV56CcH7M8Z5G4Fd/BftyUFdovTXFgbEdeOS
e42yjX6Hn4NCcJH3lD9QksQ6+sgO1N1sNesgmuJlYGxr/JrezpYgzTTLt3W/SSuBIUwVeyd+MsZ6
YuN9MA7qyIkmH/E7a7crkzCHLHpl/Vcoa36KB8w7lFxcKZ89k/GKaKtE2PorABWmOiZ/8ej4vNw4
r1XjnzyZwbwhFI5ElhJ3+oFevNGTv5J6pqBZPdARWtMbQovasqtvy585dCAOWaGymW531r2ChGz3
4F9UCjJc4J9z7NBCxVRIqxEa4rlqzgR3crHCrUkRlqRtLOmcJFF74Nhm2WqrmgXNkGyEUZPW9K8w
CrN9T6KQYk4jAT/EJ6/zllKCjS/rFI1784G3QY4Q+74J462KkL/SI8tWp5eh5TXKyWqp0R8HCCLg
D6z0SP5idgtw2s0HWFCIT4EK2uAesDT/EUjEZ1uqnHSkeEeEwZr6hKUlRWQL8rpc8gieLgHfaNeq
VAM64HoKUWiH3k5KY3gXLcuz6soeYuADQbyoGKDA+n9VWRfd+SfMx9bdw9xzr3/eNT/D/9SlfFBc
OEhOc7shQy0ajVRyUX5iVyPOLrH/3h7Tkdfgz6widZAuYpDLGAAf0607GTavgjATyFZ0YUs7XSb/
AL6BPuMMTnCjOpwT2oPNd0x5c7znqf2wwIyTqEziztipB56VbsZPsjmqVeOyg/l9J8WVtWVTC7OX
qzCR/qNkm4b2f9KVBqimvkD6CcrPvbseAODBza1jbNbGIpuI+2u94wwqhqeDW2SMhZciowapol/u
BWc0u8RH44qcwYqd8bP2hg8tAerBr/uIcXvkJXB91g3WmMabjcysd4v2DjSJSBcAakINZZ7lDq/y
GIjmEpuKBF7UjuPeUQ7EcyLYGZid3TutJqwwCUWtsbFcooXsNsMSVGWOBveBdHIhO7jyXLOm/7UW
c//NoQtqLTJgYdgOv66dNnTJ75BLKgZyGHJQp2Kf0abuds3Tcr81PGnYEic4G32hqq4tAgLY1EuN
kAHPFRuGLy969N4LJhWXOidIoJyLJsFWVRnVqZGkjCai2kNe3LFbNRcJSYdTf8JgsEhSseiX2kau
Q1RA8TGm/uDj9M9cUdBYaMbM8nTbJUyhGdL/A8NH6DVlbtkaC1KGO4jPKiQOSt0k2Vv6JVaDmCYy
z+Bna67AEEmNfvyAl4WEa4JDYO4ISf3H/zWWfdzJg2uh4/lbeJpL6ERAR0Wvo9Xn8Cs7d5nopsUr
3wQqvGJkDFtjAhK/j203gWpoEjdzgVZQS/3l8IK0WokQAn4xh7o1BFp+bBwzjzlfRtxswPu2H6vv
vihF1YBB+8xBm8xJTUsyl5CkmEzIKlskMHGIbqJFSzizwGidUDj8a5CKy0dC0LtRNGGysVQjqcl5
4K9u16UjEEEOn1+6rfHGl+uwQWF7PKRcBDJAWfTuenilEJcmnrX1Z5hvUcacc1rR6F6tH59k21Zd
ulXkafjXtitdyHvXxy2owT78vOMHegoZw6eD53qv/WT9DIV+OSxbxSZ+dJRR3wGL5BBKlyYUAkC/
6AntAAIgePuhK2q9eLLkhUs5OL4wU4XspCaQkGarGvIPCHVkOyS3FXTZNjGHxCb7HbvbNESZaBqR
Zh8wJVCkjoJullCwvYpnH6P252HT4yTuD5yWfOL9bexoSPboz0S4Arieds6Gi/UyddPbSqjV3y9i
obG+IaXwaBnjfYdSbxQ95MBRv7fwEO3cknjwLDwkRFEpt0gwV/SI2RmccwFgGZnxAXAh6xQCQbUv
G/hK4SwD6rXUsbhOTyOKqdSKFfOdBS8BRTsTLn5fWkdm970cPXuAxJK8HPcpqsdia2kmF/ybn/qV
gr9PxCEXZvbeyxhyeejLMZLWoLerVjEXQMO9MXR1Ya3zIZuutnYhnzcPFZpLf6zhM7rAGlnz8Ioy
kwx1Brf5OWSOMEQ6rE53u2L9nrPk0EQLWIKexOIr/A6PHloRXqUv74ZYsanz2LLuzN/TXo0BLgUQ
LyJIrgoeI9Z/dtxEBkY7jQFoO0sGfiJcolTIZIrt42CgqgAR0pbm5OgswOrLxZI3hBtv/9AByivb
GRRqnXNK7JnaSd2HKV7wp7Sp93OCUw+n7Uui92oEAFWrWDZDC2erIKuVvCodj1f+i8tm24bZ7z6F
hqc6fsvqm7h6FqD+NPiFER2Ipx4puAtkGV7uMBHU24Bh0pcfyHJmfk/GHQCKsynysTcDJtrS1c4O
rKIE5+pLEcUjzwcwZCCGP5d9J63TCp7ChuQqE10XSObZ3BUw8rzFCAV66iCCaljbUyj/vZr3eQ7t
x3vQ8uzj+l9rGxa0Ok9lSBzwXUzenp5KYAf5DYtAOkwWU8U+NX3iBFc9xjTny16B5o5f+zy2o/Hv
XoodzySzJCspiXjIyDcUTvhmsLsEWpuEJnz5eUANJC7eLRNAPZ7J9n/lMhCF0qRSWuCwTJ+1goA0
OPBglQ87IZy6cPfSmmXUipkQ4FBgdBvFfdTbl46Ot5lsOVn2Lc6h/7gSZQpfbYyr+ItecpGCdCvR
R9LkR28E9EZy4iYnb/lz5DDZnuXOlnXVbJqSwYx9wvOwmDHPUqUgUsEseFxrs4UcjtzK90xHrT1m
tZgN8KYJJQ1KSOaws8czUST1kMBh3V/gLNO2Rc5XVp6sXdoAOYh5sbYE5zdop5U1UTnC2ojcixGW
m4Tij5g3hf4kgnuLvfbUwfSQJ0+jNb3xvL7k8dkFB4Hcf4xQFqvsTJaKLMcl4YsKG6dCL+J7yNNI
4pqbBgGTjGMOwgOqrFIvruyJVEPbuvBliHGNfol1LcapSroaAfSXHuobcWYytBmtNthjStmWqHik
dkJ0u89VKEudvB4SU9ys9Df0+RKDQxy3oSaWf14QcsoUD3nPlZkEZ0Ra2F9+HcsJnKuhx9TV/tTD
ZdUCGiCq/ir7oOqxcAYZaRqcAvvhkZDe4oRIcgYWuGYMqboNutoSOrTymsKxu+m/5tLcXN1sjZBK
bdM9E/ubBpa+YzFZzCXWXHiXbZ4fkDN8xhu6pmCRR3AjGa2iH9/40tq8I2GdfofaVaSQMZfEvLt0
EZr6fcDrWSCL4jClL90QkWHh3m/G6KMLLYDRhAmtXXYNm6KmFnwfnb4wrLWUya+rx5ctTWA7VybD
vh9Gkd/plgxohwCbV5V6ppnm53QW9O2Xdl6dFp+felmIZ0UG73HPxqGVeTpl22LQUyRUWWO+Hcgh
jXz+t1x5OYuvasUtNl2d6rbYtl/RmVzP6XYx5lHavt/kzFk1hr5CuiqkL8IkVd1UjsVkfc8JhGsM
l6PNnXs9oxQI2l36aKBdY7NrE68XymP/LOp0JcuPXzM+kBKVHosJy0sK/Fp97Wy8ig/o9LuwGLcP
0hFr9Sr7FqJBMRCfGglKalVSZJ81S5I+gcy7/VGN/HsgcUumya0Xsn9agv0BKkB41zMTMT81uf98
1GNUAMZdXXWnOudo2XFvpZEmxpAC6yTDnQHkp5u3pzllJONp9r9C3K8IJL+KQS/h3ukEtXRykqTG
2Igah0n99+6Oib8pPuLEqU4LooQIYc7R0KQeRCIUmXvhrtfYboA/o8/prI02Ik20ZnwZnSfqV5Yd
RFt6PBJeIDVBInabDHFKkcOUctLt0+GD//iQ2VsJEKe7HEWPbLIf5YIlVMdGARz70YhF4X4HfaqL
hDiRsOLwsmJ4tNphayn3SmO5EvD0rEr+NDfU0uHa89H4vmDFl1IHnico4jf6T9JlwZY2xzaQqcsr
pla46HlZYUyjwxdD73JHNOckg8wY7LzoCczaTCKF8rbq1jhJhD7Q27Y6jW+l9GT8H5zEp85No5t4
MsRTsg71rMkIRYT7s5mL/vAguf6Td+faTCcG3H+F5F64YW9fbV0vfnB17QGJ4eOnk9gsOu/fwSKH
BKBTUnTNCSG8W6piuWIpWg6B65G6mqzVQidE1FcfxUUi3M4+q60MMrh/6Sbs5UmUmjwLea2jmFoo
pD+/eUzwL1CHw4/fMYFGBrtjU4PB1Q8j4ULH5uAasNvjUWCL+i5h3WUwtLb5CGzK/ndRuZxTTMb6
RzS/dYtWCYuOxAlMobkivkcDfFairWZWrVDAIZXmohb4xiGsTS6HrwKezGcpCgRiYZpa+vd5WNkv
HmS4jMtmYP8wTkJ+0yq8xczOt6hRb4BryrILELlGUZvVeYuvZR/AtkcX9+8dC35cHgVqMVNaG45k
AHWxEl+NumAOMFBdGEzvgzHnLgL3gEN8ZDFhpCqdCav+uAmmigTxRktSbTIECDqedgISzYgnoeky
3Ei16ifBCiQuQLPc8P00PUJAlYKFmHBVlL/PEF7rz2o5MroTyTbxWnSHJWqcvL+jpdUoRjmmq83s
hqid13Bm2wZFVRQzOLVhX5kb6Lhg7CUr4+VdpFtg7A6E8shBJR/GYBPY0hET9U/S8KeZ0I9jt2k6
z6F4vYJivRXm006dbNAvjUUvydU8yKZJO9+UXaOvreQbXj+lewFlbXbntqyabTAbmSyZToi0mi+b
4EpWXRmjWy21QrCiCbMND8Lqk4o2DwgRXhEg1o9Nu4AsJ5GipN6eByRPIZZWzzoNTF772gyM5abu
PB4anf9cbL/k+xSm/77CPbF5750RoJQVneXH0KEVb/LM1xvZR3hh9gnFKlrpOoJxnJxOLkyJ2UnP
0R7S6pnre1rSZoM1EyQ56NDfqDZ4rZZDMzGxCwR3INA3vUGv/P6d8/UDNa7lG/WbV2O5qtLLgu0W
iX9Wu3sjhbU7HgXT38kAKZx3mtoFwWT0n1xBt6vKWAqckSbXoMxkfVd/x3Bjv0O1uUBx3V8xsaJI
VsFybTYOred329CItzUQlzYDbpfR2AOJKwZZXKcpEoibWjISlmmP3JYPv/+z2u3ZnTu+1dAf5+Hx
OASUnp+BzqIE7Mbg4aGRPPRBugljdft2kfZ8kYevCDpPMxDSSvaPztbRtJAmP0WpRJDxBRAccfit
h6TYy0S211tWv+5GU83iOY2lviy4tyNrVxv44j137ZdLEwEAJnRGHIkGCdc4jwrvjXpGa1ooY3tZ
hEGZwD3UuSb4Zu77j+ZL32n7OBSRoLMwIS80U6hgInGYcRntQY/4qi70lfFGycHMD91eMojIbNJ/
laQK1UA33l7GTlCKaGU5OL5zlf/UDpjzTCYjTZOrKGbI6V8InVHn+2W303V2fNRKYr2eugZc8ycF
nugSuiYFtIm8I5Uib+BSpMA2NBN5Bmh+uEn9HeKIM8I6vRvCoperW/rZ6jfgMr66SM0UmJu9cX9+
scTwv1jHfZ1t/uknzIxY3kb3q+MIDP6AVIf/dzXhaapbT/nMb7RzMw+j7Y9feHUxQEe/lDwgB13x
FYXOo0R3pyEQ56p7iw8PF+++DcRBxISTtq3OKIFX5sTDjdJK+/My51wRem2fEn2TURq9TJ+XT8Bw
R8erSdgM9LuA11s2e5s1e0uHlZua2Pn0NdUss6B61N15Xn9RUtljEK16cS0TKA86c2wLcyLahxeg
qhzBA//82W/CA+svRa3NcF4iHY0Sflsgm5xcDyn+Bv6zu4cvFAdeeNwc1q25R/iYe4wQ8UDVNS2c
KV5TtiTVS370/464G0CPOD6Qk/SkiRqsvLexRgML3yLONFukJYOJ9Xh5ssiJw+uhR830/JWONHKo
SjMN5PSVN7nk0FvjCKmcbsKT0kks5sBvngRcADrZIsC+DKpdIs9ei/dGgVQwh49MkrI5qH3kjhvl
9KSCgI3O7uaPN6zvAFE1Xp2yRhoHspjLGWpMgiXLLzus9iBzM9Lt039JEtAa9iyX0ykygATxPvQZ
JrdoghS7Lk0Jn7UQGn25xx0aF3i0Az8faUU6y+ggs4qgXT2JaOAg1kkAw4fDcWDoayQSL9HIoEIe
20wv3bUgZ7IECTo5i4qHkL1L5FRfahBfogf5EXLNPS41LHcitFRem2HFw6YLhhrxjkYxsdMXlMQA
6X/Bux4P9LjQL5gXMYpEYjmB0Rjz3d6+nm6AnvYiIOtDOzH5Q0fJKSAjMhAiOXujnxK/Qa9a06PX
VWYUPN2t5FZq9LK+oD9yhxqwDWmTHy/8yqAmaMskjEy/blev3vWQZuxNPsnQnX8ujItk8HBvWEp2
B3xkU9AD0bIzg+K3rR8ZsfWiDkywNOTFPmaq7PFr0/MV/HXw3U9GEdosPeXDrKlsRX9C10R6Vg6Z
uMIqeY5KSEVRWcXL5Xrw2HdHLMTb8m7WmTvyZxpB8Q8Jy7LzodAQg6joPrJdxTGVm5POJWqusSEW
4kvc4A/pgQU/VIqdkwh4NPmtjGnKL3K4YugWtW+5gQnsKcYK/k14jWYEl2znKjY/C/QkCXup775h
UOexWxl3tD7Y9M/dTsH9AVoSlUBaeWxG91kMgP+R12DwJJ7CsYZJp3wFDCA1luWUmy0C8rWgdLXR
yY8O/IxRKar8K6TnpzMMrKGKr6Jx1hbubxGnihgxNTHSWom7kvfg5yMCU9ragcCsxneGGX1PWWQu
vOat2EuyCoCM16S5GyFLv8Dz5dyxdKKEJQvygfWr0XPNCB+KmEqPb8IXgZCPfwkQxbA6auqZ+NVS
KjT/IcsEwMopQm7SA+EGbCiY4w1/YQISQSKlkCeVbspqgesUEfu9Ogr/W99ZclVWxCjlxIhxwwBe
LVGRREp94td5Z/dgi6WZDvLw/KvVJ4zFe1K3iheNWL8ahqSlNeUo/cQg7Viewu3WcghtpO5mTcfF
sgOYA7buU1A44e6Kuz00gKB5yzONdgCuWowYnDtlJ4iQOudP6jptxl5k2V/ZLmZik6aBJRKAQkdn
Ed8q5xbE7dazaibTst/toVUfYsvjZD+eJrDvSFPP4jrz4myqdn/DRdvd1L72vGrDWJ5skxOaMymO
UWTjqT16cncefDCyKb/LdjAZB153fXPxLvJfoC42IEvBcEoALjpyA2BPM0Qm1onKiEp6zvIZPLDe
oQB9UI7m+B+B6aSEDXldMSuFTIygiUY7WXVuTLgAZJjOcNHDJjddYfdxiI3l992T05n42myr24QC
N21drj8kGxKGS6iIT9Zjjl/nG5006zJ/LZlkJxyUxsm8VtqcNM9zWfq0iMKpPBHeXoVm/ir36Fmy
Hsrxa5iU9N0azj8bo08xUKKSGNPat/LwXxpWrwhGt7LTIHwjZf7w7s+EY3jD1GmLLFVc1NjSfj8F
xHmB0+lcac1ljX67dlp7MWQ1OX9AViFSMbqN/fIlLDmiwJdzinWAWV+xDHIUQmXp0/EB0fDNvN4L
QJiqF5Fu73/ZdFcR11F3AoQAgztvg/iEueUQsrkZc+Bkgcprc1YxgHWhnJYZK4c79E2Pt7IzZNaZ
zun9gwR6moJUssbg+qn0N6YAwRD2NDdPm+4yOG2VmyRrW0CIfCJQoPrKsWzYlSVJwgCY5Dsw6QDJ
xscvjoSA2xkOpHsAzsl9+afCd2DujvDFOt7roW1X5KH3ETYXqWCtzOaGtAOx3bUHV8CIsp60SZI2
VyBGhlo5pBGOdbjJ7BQibVAgsEbEmbohzRg8qQNl4xJkG1oEygGVrmLsEwCXd0WJk+yjppmSxpRQ
UaU/SxHEhf395FtH9kzalyWY1YTYZWEuZmLGkRE7zvpJ7zsHvS8TKkDt6u2SSV9MRKLG8MmBHV4e
no08cFzlGjvJXrjge49HV114iCyizuwkb4TyW7NdqSA/1/vTGczQ8ks8yWmi64oFTXTBZTvmHECn
/MOZcrVsEVMmx+jvB0VMPsPxG/+UJrvtYMLy/WP0k34vcCr4wsXUIgS+RJ+/bHDOAYnjsTCPG5V+
RPb+wNRsLrOpuK6q2I1N2svMcNkmWVpWb+lLaJqJqH5Ntnx/rfscscuKXDhSsbHIF9ASO2xe4iLV
MKsB81Lz2S6FkmAn6UOfRxQsovVSuVkcSe1Xt++Ua9cxHJXFbIyX6McBweIj/SMPJBzr8NUZXQwf
GKC5AV9ipKB6yoNAz25xbjLyO53cS8YC1jRlWXlMTVgogKMwGhDT3hykOH9b+MzJ6Jgeh8rHYDEo
x9/Z+FzHxUm4MgpDik440YaDfyYrROhJPRjBg0SpD4EQegjAFGvmyGwhwtPM5fL0spr/l/S+CpXn
lw2/ovJTtfjluBZFk7EVo5bBm64st7Auq9P4ahZKPMahd3sB+R81rNZ9ZLooxmzWAD2JhtE/F7us
+54LTvfqc7mWH0ZIAUlu4OuAyzcaSYjnmyOULddWVQIB6c6lJdF9OFRxgLniFEx9kiKZ4yqBTNAC
QXJIZ3Y8ZoaYRpZY/0hG+7WN7tA03EaV1UsFxLTNktFDJkvsgttC+abJMLB1K4m6DTlNdtCVeTf2
+SoEsXemHA71EFVgL2yRL1bxtu5B65iJ/RR0FguaJPLOTANB+2gEHGcPHGICTfgwHSKZCdgDmy/m
IqDaWrVVZohKCu+GljM/0kNvIvvrq59ajXrdB98Ov4uGUTANwMHdv4NaJ5C+YRpTghUz93jT8d2z
2m3Mp1cyxhsYBZwRwfb/Zt31F4azyjQ4O38mlFc7CNqp90tDGO9I2y6S43+I58vUGkubUvDwXT0p
n0nkOK4gjj6prJ3qoyu0H3jya5sqriCWpgzxBwmWVhp80+bgEPLiaJiVHZZcZScbDWxJwXcts1ET
LiIF8gpkmYnK1VoTgvkAt6qEedEaAhXbCU+fgPlSrAb9KhkKJ4xL1TlgmkJMqRymeCpToUZw/aDZ
M4CkIIAjQsBFNyryh99PuNFMWIp5xCaE5sV2CvG7HWWwUtTEGUj8ZNp7rk3l5QAHr0os3CXrmd82
k7txnqSVPdfqb+shVcaoslFSs29cRh2eW3ocQvSDPTfHJuWmgvAjod6teaB6B1970ieyk2KOPYQu
nck8Y68Yp1Rl1+H3Axv59NZXOK0xmJagowqKYi2P9+FLXacz2ZMVQckUIi6RkWizqfWRTHCOBcgc
nCPhuolZTSmM6RzZ4fUJSw4SL0gn7rZIPA4jLsiGnsSmbR8tfgBbzuWqnKh+zqFOlOIWxXucopCR
7GxPvdLBJk0/V+re+Iv8zvoCoSURc733Y4zvE9c8gJlzZ+5Uns+pbEGtMgd6pKzj2289wQ3OE4oI
hIMUKm6LeHbu7bXssRwuKdbgvlZWbSo3F+aUHSBhRvBeiieD32LrolRCqH/rKmNCOiiQ65TR/sXV
gs0nO7GJYk9ig59AVREbp3aFnFmTLne3/rtRKacYKQZIfIWPHYXOQCziGoaVzArbvvX+YW4232Yd
BqGt615m7aE23+blOiI+IykgGrtuE6pe4cljrS1XKTAnEaA2ULqGgtGK/r7jtGYHhqJxW8n0eXL3
9j1vxfkrxSypq68m6FUqK/Bdgy/vj48eRw07jZ2ChCrkWxldFwqdRm4BOA8m75l0ZPWOasQct38T
b+fKV0YyrZK98vOw0XbO+pWBmQWhc2OdKDQflo9jRJRq5qYefE1WJDyre/KEAhw3ZU/v5uh6syWR
qhah3FxaAfdMvidAtfnXM7cyrYBD1mblN1l+eOQDGL7ko+4S+ptA7E2PgAyjeUnwwYcPzDnEZaNZ
7Hpscc6Tzj6h4BFtrdhVZgGoc6EtTfXsRHbNn+PSFjHzl4+py9bWd2agcZ1bOW4jgg7/TMtOVZ5z
uI+pbt7XlG80iaagsECX5RO51CuGNtewgLre3c0Y69Ngm9jD+v078C+pykKNHbGc0YcLCP7MBckp
1KPOGAO0qjxbp2JmGXbyFWgM2GtV0nwABD7cMREoAuyII635WJSDMy7OhajZsg17HwhLaPWMO+9L
3LcuwmdoWj9hxLfg32AVIE5aAHpoWjf/bFkkha8wgEuam4ui9OI8FBqfnPz9mbwpPXImzfHSMw+b
Xrqpx/rqErcYG7RWDnLlzsUuQ5/xKZtfcrRoUdnTkccuI6me8wgt5v9t1+IBWqvsIPF6M8z5Dp/B
HU45oIsCwZOqTQjurEi+iRRPJYsm4Rime85ecPRsEV3J2JHuJo8lmu4hKYyGV2gil1Czx2e/ihy9
XdX4BOJKCn+2B1QiYVFXZXTAOZFyEJLP10bSkXBh3uNdywlEbjOpy2YNBghSN3Rl34wbt6qr/KVQ
xnAy2VactyGMeMKVNaoQmxbOf8Co0JyN+dI7kxGPeUyz4J2EcRvfFbtKc2jzqQVIXgFFnMlREktg
Ps6cyaKGsszMsxW+t/Zp9L1t3bWwq5xrRiTT01NvHU+oXSjXMAyDe4BioqbiMTJMVgIsxSKRM0Zq
I6E5hE7xiTSr0BPOHVOfZg1315kUdXVkdUkzudsykfBOn+6mD7ggKWp29j/DgcAgbrhkAVZq9GMB
TcTwHKfujYYcXjoz2dnlkqNSsx/80oaxjZqcg2z821YhOqC7Sf4UF8GcM3rHVXN74Ssc52B6c5uN
QWED+FYVGCFSTNBtCKCOOrnzIs7cbYB98fMf/T38qcxCz5KSEA/ARutRHM7SELIBfS7io/DYKiuo
3j2ystYanHNz+o5duIUICpmdXgonYAID3kL2xUGVWNoMH4o/sYgZe5jZrK55WpHZe9/n1o/9/aJG
feDmMj+QwtZtNlLwP220qEgl8byGN3YTLhxk0Wavf9GF9rq4UsA8198h55EHSmDjCpnOQJsjN5Xy
AiUeTV5oVDOXCHqk4N6lYadW9fCTXyDD2aCTAS10b8bkOxm5a8E60tsD/JJArrtUVkok+mLjycY1
agXhw4614lDsbhZA0Q/HhNK8iKqQIEYA69cxmG2sP82WpCOVbshgaUz0rkeH096FWiPL38qlH1Ft
Nv2JVCSZl/vsyNTFfu/QDatSAdi1vsLXcSFvS4aZdZ2IG41RMCDHxyg7KJgGMflt4z6+O2T4liHO
MMxQ2qWQSb2eKhrKUrUEbJAmxvniUTVySK1kagr9cM9PuDbxlK9QjyhlZ7ZlTopWKPnFc3yJho4i
uLv3JXGaZIHZPFtNHAAnjyNAx8MlEqGfr4kHtbs8BuwI3JBFkNC7c4vbtxli70d9dxKVcTfkFOjp
cwz8DI3f9hYvNAvztJiY+VkpIiYK2Ni1mBW9+sgA82VOiZ9zlt31LtDh05Dgmg0HQM5VAaOqCz+h
2qI7PR55aRBv0CGSg3au20JMgFs3txiS7DDZg/okU/N7+OhjS/CHKQbyFKoJLhicVXzIbuLb4sy7
a4n1SaGZEghKDM3POIU22hy+tXNJH9y+zr+76uLkMIzDpA0J9JIfH9ZMr0GD5LovcDtJXY5kfxJB
a18kCDvJFfILQl5ZeQgan5E0HTRT+0gEwEY3BjTs4eac1KHX4/g4sKteFNwaFEr0rbgGbhsxCF5T
RTSzBBM3XO8xl2jiHOrPpGszymAyxIYR3iV6rmmWeCluO+LIv2HE0G9tcMC4YAqdPWOno8eB7Dic
cjcUvXYCzx0xj+O4HGIbgYaEv2+EoE/pszPYmRJzVV+V5/cftk63H3WiifyO+RK4ObA8LsIlBsX4
0s6FSvfR3xP1Cyo7ImgwVd9t19IfiGoHpmMxkrPIq8TD7CK/SCGgxPBHYuhNqMDVhqtlxC0A3UxO
oPg+2zR6VhkSe4BS9fKL5gy8I7T+9s1a+FBu19liIlwCjrNFT+hiRunHuosGFmeiZqYyu8RU0OKr
A/atp0hslkhPP0D9ZrMK3n2jOUEaOvLqbbcxAD2uuQtb6UAx3PXFBHw57tsHNnpagGFX3+LUUgCE
UqgT+F3zQo4bFvvlOXzu5ZoHi2Qi1aAXD9gHOJdfI+pt5c4SQoi55Ph1q7bqUQUIXDS8cuud6u6/
wOUa6p/rS9UjIDtLE/3p+mTzZRL2FPcAgsvx84L4J8gnHLhBQfeKIbI6bOQ9YR3Jv1Ko3HCOZobi
+9/sadjUbOsgn5UvLEjZwpvWyQ1Eg+6RSdh+4B39JNr96OokHlP5O0uST6CKoblWO6bwWgYw9D++
xm9SEQED+mvMIZm6eYcuNCR1+IQKxGmFwuhvdUusfvN4/C3NuAJSat8T5XAKm2O+aawiIxwF572W
O+yClwjC9d7WiGUO/+I9ns94hAvBZbV8JNqueMtNOqjV5HnW8kX7e/z6wezT9jA1PiIuUwSz4/Vi
AgF5kM5dE0x72WaF9bpA0cMnc2k2mdJ0LDQV5mhovFy43uOofVqdesY0USwCS8HKDBDFXC/SqEK5
HkwJX5Sr3TDpIeUgSgkVShV3j77J4se03kGfPciVK9JtAPAhqp8KLUu8INCUF/KKnOF2lOdTFSo/
9U0NJPCybZa1rbGyS52iu8RyQL8BEouWjOt6aeKnut6I2PgPohMGfTJgbrWMzlIepN0KdMZoRfEd
dRl4h4xgQAy6odsVtMEBKpkoxZr8yInpbStgHiAq96xxSM7HKM05z+YnxRZiDW5hIKduXgXD4YF3
wnh8dIvUfPE5lGYyIm1e1BK1Zgdl8O6dI1ydAvFFdjRkVDfqazNNZgHqng7szDX4cId+bG7xfiAW
Hxnbrc1KiKS1wslskx03pn7Bmy2kkkDNSnZwRo7xmytiHYYl1AzEhpYnNUVbh7EqC/wbz2HwstJ6
UNrMnch2mCDZxULcfJzE2zlJiRHCIBeUt/6JwnIUFyUpQ/xDjb4NQhJCB04sGWV02F89gYcel7xG
aQtTvPIo8QLNomvLiX82w6TfTypZNu0a5mYAZR+ymvGl0JySyQxbHDaQPJ3nbDmahRMUE5ZXk5ZR
PHc8eC0LY7TqKZCUwx8dmY2FhHsOuQKfziPtkO7zCuHpi+cDa89PuVd8ZQAeYBj9D80XtlrAAEQp
uGxw4qJ8YxHCh3EIhaR4fNdOoZrI7pIG1g8eDZu6uSF7RViQP9nvNlzgs+ljiUk8jCRakm1YuECy
FX1WPADA+WNS4H+3Zk+AMks2teIFq3BwIL6SaTjsF0epoUCzhrJpQhd6Pi6qPN0e4rbYSQ5px0/d
u+Lxq9wDOEQIB5tLDOVHPKItFTNb0Ybc3GFNpmgQ+TgS6bGonKoBKP2GaQY0Wb3rrzNDnOLmFCF1
ynThABHIgaNM0EXii/9GII0puNCsPBOlqXi0HNRVu/5htfGxLZRTcLPQ7kCkqeAe0lMyKbrrBKFX
Xuv8xwxMRlO1GgdvUihL+O1WZYyk0Pfyv2ofoHHqXzn9sUlRsKcoBsnCdOVpAKWGM7E7yXpk72DS
GScZzqtWnK3nBBOQwDhRCz4dyVz9ltgvv39juuMzBvYEfJfuOX5lFu9jbOB7+zoWl0hyVx0pwAI/
2Xn/88e+2+ciq8GmgDjnOrszGkHsD5zmrIdSDZyPsfJYYDOcn4I6Kcj6a0Du3ZJZzlsKZZ/rQo8b
3g98TFwAdB3Uz/OmRmnSMuWDPFhBUb3f2A0g3/oFbRoRa6pM4ysqXjJ27KjhtNTnsw2SnznIJbR0
SgtRP8gYFTFyDbO2DxSiJTPddSpUGQxrBBPGoNNwgVVDG+lrj9MrvsnXbHaj2pttiYHL+q1DBC6w
y0XgPbuK13RgppCFlLOZxSBWX2zv8k9hLt12dmTJr7ACq6sutfc23QduruB3JOHw6GJ9/xgXHH+W
A3t/9Jgx+MiCdG6ZdTyWgoqR9AxFYDqfMMvY/n8rY+FoSYhaAAhQHgyrCkPggQbtEagKy4sLRvji
l1Nf39GE+61PuUSYdqMcwv8Knh5YnEXPXvmyk7Pac1Al4Oe72vF69aRweVF/JXbBNqoY4fCoVZhc
cy925RzzeeAz8COOFlZdQhpKP/bAieFIjmZ1/JUtz7mh2FyGeObQuOG+0JADQHcIpRSaZ0m2lRy/
I+OZ62wNTQ6pMTOogT58qIViOX+KTtciZsmUbcpOrcN2L1YvPPA1oFk7jsk3s3hStPOdiKmkcxcq
ancsaRGRvgGeR3tBEi7WOdmCK/3H4n04OXEy+E4zIAyaybSii0tFY2/IJGhde1hx+Jhu8UFN+Rcz
L4UMHhxrv75EiQrI9zKHg5Gpr2LEOzmmzr79CKS90OKJq62dXfeoNNUOmeV96RuheMgZoPw7jXvn
i9v15A4a0kDx4GK8CyUQWEDT4MeRlyBY150IuV6dWr4zQbXqCrWxRHo/iH18kN/6Lbx70xICqHD9
w0aGUGUsIHo9zWYFn4giPowKx9Hx5uDGXCbT9/0w+JVG+YXefDRHwX/kfrbCIz6cW+S5cd9JBLt8
UB2faw/nBKpWy7Yer5ireTnDWSSPsaVNrjtkpOsMtD/pVkhQGf4uW3jOXxqapUdzhcSl2tlO2e5O
g59X/pxaoXbDHAmrL7pFaaG3v8WVVWc+UgjC83qpKk3I/ioSXJdxVfD07spCA66JE16cr+GgC0ID
bt9mIemwt0d+/s2le0uWkCB1QXb1J4Rcb+AvEDZqbIDtS5QzVmq6s3uEVr8JMD+tl2NL0yNLX6GB
DMtXczDT2kaxoWg6RgDiqP95KXQnfeUT0M7gTMaea7dmi/ZmKv5+kgFATIpCL8oG/7XvCfj7CaKB
ISA6SrnlEru+M810756xUDyYp4f/fA5KMmHU6mjMQbHGjwVjIZWheOMQYqOm6XC2pZsCGupPOZo2
FEJgydeVBBrnjvCoj4EBiN73e9PcyFMJJ5eD0Zn7KumYO202k8ZPY3qzSHk1cd1GAR/T/EAXiWH8
vgen8kD95xVrvthsSO5j1kBT7nEJpK2q3NYIW+GKKdzS/M2fmFksshHLQcx3mMNowHK0ejCfEnSN
QcppIUqPXlyFVthSc1wSzK9xMje4QJ7CkEkKXRe+G1vZ4G1Vy0OUPMo8VJuUruilOzaY6sjD3w7I
NjoHNlpi6eOh9Oim3lzUGlQ20GQu5q9nOOLs0W+ryF9ykYm98Ejrfji52+OvHuDXQDmdPFBZ1Wbz
HEwX2gYUTGHwK5f/AULxjO70jupWVhQaKweaJOgwYOgh2xMi43f0FmcBzgQ+IDVsilOUva34oiI+
Q0BS9OJe+wjv/3MHxYD/+PZThv9zImu762vCfb79w0gUqeZtJ+eo88S56SA/fI9bQN8/+/nxmubs
BNmPSclNgGAqmkAS/vpyCaslSxLehXtebCT0E33gDahGRDrETwOhewb8Sa6hOI0wKWoVD2H7kl/H
B0HPA34/AggAK93AEEVCFdT8VcjPHFWFSFGvtvDig3Zg27GD1SkWSrVo+YfVXmYtm0Ad/Aw7E+1v
UOGE+ETIcQaVOH8j2JQGDgsksFd4m7uHLxOkOEXqSLrtkLcVdsFnsltEu6PU8UDXzoARooqYw8io
cmhYx96egkv80zV8Lz+XtFjTwO8JAaO7JmPpbVnrM7Sd1nYaeLZXagSVL6uGHFMRrU0Bg9NB6LEy
cWv2GdaEqsBib2sXhPrxVbt9Ppvsm7StK6rynOSrcUjqr+2EGEWoANlEgAFWRmdiqrh2Z9Mufb/O
GPQ1PBeU13o831ccqBYxbbehQHWyCYZs5XO1oncg34L3WoP5Vba5GELFX8MSwF2pdt0hGzYCGnzl
0Y7aFIVjUTRDq6eigCboHvMkVs/AaGUdfqpvpeSv5Sqejb6QZOUoNVq2Tai0Ul8qi0tOWDBD62rH
zTpIQESnu515a/XYw8cjpwVXWZag4KYn6A1zZcbOEXrhzZ5Y9HzLfMQ5nYO2ahqK2jfFaEQsPcBh
6Vmt5EEOTLD5j3kVPV00ncWBoGBdAvMooiYU8w45d6skK5KUcEzkgpMfXO/NWTywn0xdlSmVKAo5
tiEmUnvQXIhGn0FAqvQRXP3mh5oiFPuHbtYM/K4WUVEcuGMJ2yTc/sK91z59CZzxT0KepCxPM/Y2
qFT1cv0MDIc9H6So4oeNhThiCBjj/O5sSE/5/HiFWVwyquo624QdRabxcjykOPCL6rhXj/xFQfAd
CCuBaxDaT/P/Ya5eUSi+3o7ReSkp5peBuz4fiW8X67nZXTCshS8BmRJwLULFTo/TZ/qqaSTfXTci
SjGeL++0k+xtKdTh0X43b1PpouHw/MuhR6U/VFzsmmCFx13Zu0y5Xlq0xhSSbTOhnfek2nP7YHfn
TYFqA77idAxEaXj/n9ZtA+h0Fq7zoYzGj59yMGzddDyvMoVmDcKY4lf6h6d8l/OQcYbiKFhgzkew
N+cOPkprclmwrdM0sksICp1uvrkItWIiYeDeiF9LPZ7szAobpQZA2vDMkN7WI65l/sFuVVPX4IEm
8u1hcHuRuJjs7bmVI4hzlkWHpxW3eTBhfLq0FCyCbZIC85w/YU7zAPTw2JStxAJv0/rlmjtkoycw
1YN5XE92o7evEVGWlEUgPZ0genSynv1jabt/JlWbNiFIhsJ/1Cly12aiuQEflv/PtO2i65WeEsGm
8uHbfxhPbznqcJh0yoZJSG/ogC8I1QqwdvzwOf5V043LHq0enAqEe3Z8YEJPEsRdiMt4qnaJkwvt
B+eM7vMd/ajmOBjjDg4l4/9Jy1Ka1W2z36TYm4ok0WZfNSx2mGV+QKd9OZ0PGIo9eJQUhXQ1IPlA
QSrjop3uu2rJi59Fy2GnN6isgpBvXVHlh61dpKWGcoHLu4ahrwNEEMKJsdwCtngr+hJHCsXkC5Aa
9HlV5QbG7UwiNSfr5x+qIqUSKfsIegNjt/YmG+mPJvwNAjg4ydbrTCEFVdfGBK7pCM8mGm86pRe+
/121jTUAchalhJSXGyrEAoJoQrK1D+BCQYKHACxERMS/ndFhYLD0mwzQmG7E7jqeRIwoOWeL4hdS
uiLt8Oi4fybpa23BbpQex9L26CjlhhFGfV2Zil+ybOaT72Tz5Fm2+1HVBqv1T+TKrclknwxhpv3N
e80EbzrfxlVO8qO3ERokIb53YA0E8ercgWHw57IH3+iYYSiefVDpvwLXq54yK4xsOw9KL9YB1e/V
FNcwp1uW0ZobqMxr3823xlSpR3CyVX1fl9kp7SEwqYiY3D36sNMcmNfiLotzsHz+QdcWvfdtJRSm
rSOXtzvsrWfhkYEjEyFjdFPSU9m2Q0KS1NYlx2902t381UlWPyhljvoph9ok0y3I6oTlp8rlcnFt
3EWMdPP2wBCNdKG5oJHfZuQ6IPIs05NalpegQn1cBBCnG1vcL3aioDvYYNZ+0clh/bcJ0yxE2gM/
A6fSw3ZmYyH+XAdqYMetu6x+tuHkrBhSL21iN5B7s0VoLwsYplFsEi8BtvyiD75OaavhN0+PL/4S
zyuyvpmaBmdiIFV4TW/FTDTkNhUS2pslDmivx/hOlN8T8aZ76CiuE/8k8Ahf6wnUPaa7ue+XFNoK
oUSRteamk0OxrKfCyArWKlwoRrLvW+rvK30+2R1Cm70KEvkQf5vDfYUIPhWzAzgAOJRAeZrQcmRG
7eLm3IAUqunZuZes5Yazor1ixoL43izDELWBi0P3CqWU/AzPMoJJUYc1TspHITpVnserFoaW2tpu
ooy5sgijjW/ht27FtyEUVH6cvnmFi7nGtfE03cAlByeiXU7pIBM4ezczxE+9xOwiC+3U/GjhCfF8
LHW96omTKYfmD5cRBDLx2WXI7zfPXXzeEDKugYjW4LUcQZabsb+/gqrV0j4kBS8Pdr6JAnhsikgf
jDJx+64P+G7tewny6HaQYMiEvtJhnUqc+3uZ/UHjmImplWCW/TUh9TIFzZ0OKi5hXje6Hz8e7fTn
xm6srUSsktOV8Xo4PkSR6Aw+f24AjRqxERXPNgoY7dKytBEkXo5q4x51CQB+vHH3lJflKfGGWTWo
0Dl61a+YXeXA1o2hhY8ppCALUi/xBNXgAPt9fu9k9j2eyUCTIwLrQnRTerKCLVeaC0jE1eLhHGo1
VcmCG5JHxhdDd60hwccOzK8aUm5MmQlSiBIRrNbyLgqpPh/W9OfUQ0NKXJTOIqgTc8VoiJziKMbz
ZI0CRZOTOXtTLHvhR+KIydyxjTGXSkvuxy1HC9A6sqzsBd6tVcWi0UC35WUXOZ65NYtO0xsl2o3E
2gaLOTC8lxC39aHfEy6PNeR2CH4PujR+BYz7A0CCRRCUihC9h5H4+k9AG/86WXh6TSqoDSe0oIej
sukPgWHn3hOImdGAD0pHjlrMWiZaYwcaJo+SCBFOjvRoOFzK/q+i6Tj0CROYDZ7bFkLu7wUrDiE0
vgF79zXXagiWawD03niebj/KGbI2hSdnf2V/f0UJ0E8nykeQKylp6AEQQNhs4jB9epyoIFRaJzk9
Ke6nzUOiuN/+wugltN9iuXHf1jVghzQULdQbqXpal2YobnsRw/Ud9BdYPOsW5t9pthI2Z+1h1WHX
Nook1HieAbOPDAcF4U+PIOnHvMsS0m/D5blbZTS40/uKlolivuLkQbZJ4ib1w3MNEWR5At4BzaGF
9UuMb5iRDm7TeNPEnIoOS3BJp81K3Yl3vuRbtnDIG2XnR29gIbHPGOAg73Q9TFIc10NN3L2rVA79
e4vAqTS81Md3VZKY0IDp+ah3U1HrTXVE3C/SOY+rLsvNfthjmd9WspdjQug0uNUyRLOz6ad0tCKK
8cL3WFsSG/Zpuk+k5zIImmXBi6bNcH2JhvnvwS2gAxNpP3901rklamtnITvIoJjJNSj80dP3ivbz
bwZ7L2SbKO1x1TPw4E6qE+Nd13l2JgoaEBHfe2wxbBJWlqPiKoSUNdiPgji765ir9BDks0TxrFXB
P2AgGYVY+SDMaYs5nVmr1BKUGMb5Xor5JjUFa926Sdhop6tt+Y4nMn99HhPV7NIUxdbno2Gl5DVG
RtSWnZ7mexdJS151+gv5F3Xk2bc2GTlmsrhV44vDrP5Ec0dXonyYaWEJMHR9iFoHDz7Xh0DYgAM2
O18W7y1ys2FiiamV/kcuSfKwDAYeXbI4a3liFrjU6PLOV8iZ2hblVG9ait/n+gqLOf0StCsAKtk8
gQpTom74E61iYh3UiB7ucMmfqyI8V/tCjmzhc57/cFDecUAKiho6ZieRFuPu9eiz/ZPsUml7SMs8
5xux7uW26z7cyKDk2XEUXCE9bKutpMaqW1tqUw7DvOOZVeXhLRpZ01WL3g23Ki2PZEdu/t3a6Yhq
ME3v7eot3ec97+4Cwepdp+UtdiZQah1g2OhbpekncB+tfX0kKnoXd+gEQ1NwKhWaLDS81DVh5p/H
FV6E4VhX04+ZzTHfoWaZVqI8arCTEwHtQEht0M4sHpfftyTpEv3x5qLLex2QUi6CtPn7NxX7rwZo
iBz2UI4Q2C2d5aYdRSozi8l8vX2OXZN9X8wrIHkugQeQEpk/aNFHwtma8+8+Ra/G3jjmJ2yd/Bou
yKBaocFfImhb2bgQR9FOj+Q6G/FkRoRjJ2QkVfX3thDiOnAJniGPtpLxNxckzkrnrIL4dlbduMu6
rFMSg11IlFK5ljpqXgSIfptXXOrCrqWij4JdOr65MUHQjyGlVsnFYSpxDNKXT0bMYG5O6fR6lRDu
CHq1vvUztsBUC+vhkyE+aifA4EccLtaajTCfBFk264H1bFglN9DPVNy9o6wSW645ijH9jtOCRmKK
59HjCMDaBRlYbbDlpFNmCx9iyLUcgeO0xJkVRf7FAMfErh4owV+PUMlzB6OulyHh540KHDb8H4nZ
snfAG5Jx5O4ioMKl1ykqATj+VmZmN/FesiR8wSclNrlROzyzZ52GhKRK0vfVqTRkV3folRdGwA6d
XwCc3JrEZkef84UCny48ZrkkQyQbF8j0rFoOiKLHT+/nHjqowjHio0xc7ORHdEJPf+xGSbCyo3up
bglDXT8bv/WnUTxpk7LALXmZDbguQjdOR6yno0aVIVwSorhrE+xzJcDk/NRkQSNaKKHkkGCbEd8/
VxsEQrG0XnjiQ7nZMqRrvbP/Dzp+sLk17GFho4X6zA7orJs68+dc/7AaC62IDvnainODo2bUP1mD
bodYTj6yGHFNvvsoakn/C9B4TRYQOKm0QHB1/tXLUP1ariFwbsUDZ2jz764CEtLmuFPCHpISDHEz
2bTqK+mhJXk+VeyFSN3V+bLP9SySErD/UyIBTDHg6bg2GLv/MVi9J4tHhm5T7fEa2UN4CRsui5cW
Cyx+FQ6uFGlnZiAgR/MJIxQ1fbSNPJcGYED+1kxIS01v7acW9EF9cjunVkFDK8qDo6KiqqiWPhKh
z6UjVxY7WbnBANW/aJ5XVaa60amFjv626es6PR/UwZVBZ83HHsoKdpIoATG6Qqgy8Hjfb0ZzGVyU
Osd0mdFgcp1fEQXYtyQC45w03r8W1/T2LzTKHjNYWCRiZ38GAvHA6+O6vKiYVhzliUbyqcBPsLp/
du6xuCjESLKqW4YGLoNZt/aImue3DJi9OIz4hXJaDCAdUGXL2kEUicJ+4TvjPqIDZoCnBqRWpPyR
KzfUKuKBNzuSjlZj1cf//ZebJQtUk0G3PxNG4M57keyCVGxNs/EWaZ0891irMeWr7MSQSb0z7V8Y
t5pWOonc1jh8CVQWhwRSQNhjd/wKzAdVa7MOtVGZoF5uNUQNJvs6sHPYMvrODji2WOAcUH54jq1q
AvPfmdOfIb6zYHyG6PMiCzxNFPFaqJR2K3P94D9VoITOzJw7fAiZ/epHmyILLCi/fpsiAFtYk/Fc
hi/R4dA5cYNEwo4Y/PghlCQbJZZABj3IJu38u5A5zStt2cDYxhQRqcMcApfDiKAVHuLfpRDpj9uL
XTqYXx2fvxvKuoDKVVKWiYa2qlmDifHHRqNU0B52eYgpaPuKdwWfSkETSJJpEXa+fLKTSZ9SDd5Z
yaw0vSXh0ULPMogI/HRfj1D6gmPEsfzfQzIwGB8P7qbTGEf1KkDYicUdNzwGJ3fMWJhRPNjGrWfH
ZzejqQSiixq6DrN9pSxgxkKP8Rqt4J3Rva8LkAw9joCkS5hvVMQtE+UMug+OeJ8LQFBckKudqejY
/bKS3T9C+V9Y4hPxeVxtchMWcXnuCZloMVdtpYq9NgURbo640cXvJbcQ5QDQtinJ047RB6JzdSti
D6lQejrm7T0TmJks8VBwu7OMgxghZB/qGRWa0W6b859aGIAwSgPFMpsnS62NGKL3t9/nrnWL+3aZ
rztPN4+Zq0U5RMYYkdyvYCGWJGlPkVEW4SMAiTMKMs66F21wgUeyGSGEXxwLvRRIudtBMd2EIC+z
ByB3FzLS7snkxnfJLDjfgG2l3FRRV0AZETyPxuH8+91hfkoe/tQsCXjKDxsl3mhtzXuDILvs8sTS
FSdF3A60H/P4aooDoOzyE1xGULKye/wOTlYg7eNoMNG/wYhrLgYLOQ/2eRlfQXfqWQaWO6OiP3Xs
0OScrZEDDLoUNfnoY1q8mZTBHbBnkLz/OmFUMXZFWA2l3zrFZfcWt+fEGcRH5uT50WNC0iZ1Rc4Q
38E2cPjpf0B6lWB9iq2rLZ2hl04aaLQ+/kLOIu+9SqGsMpoMdywzu2l6MzTKNVrLNeirerFt5GIu
bQEaPk0cm03Njx0zVyPz3PembdEfRQJCpIHNrv54QCDhjBu1wMYJ7dAF+3KY83ZO2OKdL7hCtvk4
XVgUhv0UD8ubBmhmDAEgfwSjW9BhkqmsBjTHEFHlbaQZYoV30dth/G57CAWZDenRgxE0eteGd5Jc
C/LkYWSswuvSHDwRQyZOlSA+xehP70jkQ/8DDZRt2mHHD6c6YnYtwLBVBtTL7fhTFmklgqDHE7Zt
3naKpkrHCq+2y8d/5fdV0n7rEivePj/zT2aKCPy5gkb5yzPgfhCQn+3KRasM7hhaedS0NLMJVXFt
Mt/bFosko1QG+3yN/yX6hydV0/MkU9lzllch8m6gP26cItdpc0tk7JrKDnt1/5RNUT0Ev8mYAqV+
NTuZEkim9l8IYUQDMykngSD06WOP7IFb5iToqCrCbdP46Yb2rFCm+zwD+mDMJPZVbnz+JbTV+9Ph
WCycQkpYjVSistCLMsSlE8rXKV0AhlcDoz+OdH2uTqkacLBf1+4MusL07B5LlS7kcWaT7TTpORdK
citpfa6pnX3fhIFsosByK+UJCP9xr7qyK0m2Ywl738LJSJ3eSSrjokyq20QrOOhshSxync4+7gGH
20ZM2MReS5hB5UoMtUfoReiEfFnyrAPabFlbre4qu3i11PCjnXR0PREntb4i18puzWhRxq7/Zgal
/5drh/L2zduLx3ImKhMuPn6cuk3iImeNNx2GZ3wD1CkmT4OQHW+7UO6qGlVHUEedtvp0gu32mAdF
wOnPXH18L/KDxPDTUR2x2buXRLbdJ0Eohp/Z2sjnzeGzC17gEI/k7V7eb1+rfqHZVpWoMeC5d9/L
HrdGRi4ati/I8yzr9PsMT/2v2QWMGNEkun0bmI1PmVGXovprv1+JFA2ThJ8Gjnc0V1D2zfz/MY7t
aLcf+fHxK/lLGud5Wm/PHplia3eXtghp3gOBOBeLs7YRiFl2HuhYa9dgp7WEMQkwa9f110bRUf0A
FmBHjfnIRYDrX5JrH8zNfd0Q5WG7ZoOWLENz0iPgraRxskfrAEmQ8wTubiLUWGy6zgmIZwXwKEvt
Tj54XCIvhYpf2BhB+BkjXUDep+nR4QugFj43wToMuRynImFXOKuMfSK4TuRmoPZlzbJEcccyCa5c
adFnJUB+i5KMrg3tS0dZY7ePCB+1fpDBlj7E0uoESB3l5VCAaK0+nU9YTYtFayk5rPIMZn6PS35A
KuTye+wXX7Qpp2o4jBaPiDBNuItixJf75ZR6w4yfOZDfC4HZOq6VeN5jt5IV2uizeloWVrHXMiFX
kO/hB11Tm9l604YO8dbt8W38LjzfrOqqfFXcmNWvvbuZuX3yKgNg/+ynZfXUsyMVE5607vUXfNqA
gGOeB9SASqOs3uyuWcbcuduQOon8KW5k7WVpOBM7A3SbFfSc8JOkhlke6mV7JPMVMKImOa1NBYVN
DOFuyQnSjOUPtzzQ9knDZw5t3SpaRwfdDwyyG8pfEHophaI29jErYnmispJgycCExXIhDxFjWSvw
XW6WxsVsKNwmr0pBgtAZRKZAwMe5YRsb6nEIczh0wuDpE7nVjBP6djMuipEEP3Ukdy2w0qptPzOZ
F5+APv/N5Le1SOx9gQSRLIYCFxrSLFoYm40uwLsb7Zs1zG6fiMdQcBrszSOvuzqHx1cx30dmrt7S
B5HwToKNVHVqqFnWYeL6SnYI8sPAk6fVFAw82JHZHurvmP5VCDqYQfe5xlAtx7nOTf5Wss8WNF19
Igv/6e2KrMu0g2/bdmp5UNgnDmGP4+QSvQw1H64zzNrV+oYWNa4Hwb1TTreLZ5sxPm6rDbqg1TGy
eWKDzVfwsb2ahSnaAeIE/4nTq+pkw2GpxhtPJYPHSa+i11NTEplXf/kMT9LCVgZN/Kb/4ffxtibi
hxdpjrvCD6h5ehQ+aMh4S2iFpaX5YwUP8oh+BnvVdhAtSCsnDi6sVAGzMjTSXK8W/1i/9lAWpS8V
0N2Z/Dm8MQHglfFshqC3/UL2o1evYGfhwycyufvUl/xpABEzJDj3F/n9FQ9b6VsCSoLW6cWexr2S
HdPnOcLLgiTxjwq/NPk+nYqe4Qgs5aYPxblUhAYQ00j7YD6vJjGYUPHIwGecY9t5U31+B7xiOLCC
mTZCyYnWyefqCqEQPG8pbFOpBerVsynrAXifUicCvhQuphs2VfhLO3Q9gIx4A1JV2puLhW3pQZ1E
Ly4q6+n/PSZ0YMU+z9GiQ45gYLPeykFPOuSWbQ19WTmrP1yo8ZxJcN1PWnMwC9oIl0nbOUUutrZ+
UkzJD/yp1KoffmHZbuHoGQOLUYg+g+e85xSShZf/+jpNxLUt6hItlX79jc5WzD+cniHsTR7Fs8Do
GtsFN/RGdpo2xWdKifRuXA5qiVhWjZ8QB0nFKMNNk3qExaDDeOrKFJ1FnwlVB2OqWeo0kvWFI95E
DdTNDtZe0seKtMAeZuNUUGO8IKmUlfqtft4CYI2JN3nLhV71bYGQhlWeg9s5YwEJOLvgEHk9+NpJ
oQbRaZLtAacQowMpzaz1EHp+19i/QKhPO3JTGBfYOtz1ZGn7mnGJ87F7u0x5ZY4MG2CBH4N1txar
NnKd0sFLNIWaxKxkG3RaViUK/1FaqsxrfYiOkqjPAikSEcOafDNbDlqqdszO7lc9mRH6ymiEhoMH
saSNimpu5wzrJQ/TnRxPW0XMmzMLbI2o2ML7bU4AOasFsPwZlHL1GEzSKwRFJaSShYUjVVTwULva
lrhZsTEAnZf21t99Of7Tmvq5WYzrgvUNDZ+jI6JUAqzWySCS9UsUrrXUj0UhNWmYmhWRHj2G4OC+
MkytlYu2pFKzx6HfNR6rO+V/H+tWO6ivDR2OS4hd/bTw8W6qbR5zmTKuM2oBMK2p/vRzAH3J5dm7
MR2cBvgrKuKNVKw5N5+44F33pt+TnG5CDxHe80cR4ORvkGLqayBlxzv+k+wcDi1zUxqgS6z+M+W7
GtMB7iHjbgwHZNPmF/gReud/NEVyFLeUl/2f5k8DM8JT1nUngxodu/Wp4gEbRzYjCs3balPjWkVt
HBlD8OuRPTfX7qCxjShJBzWffZdDGB3p9bFdx3AC7CySyrJSLG2QwU5+pNY2rdaLP2EYSltLE101
EF6ycJHQW2de3OyDQRGBX4hhU3MAfz77hlwiUkdaPqdNPJplMLPQTk+zLwKcGUKew2v0khvW2Cr3
sPU0cm7bEqWB4h6boBRvzMgNvwhnOvYhLuKjgi2Hqn9t8azJ8ZzjbEzo4GN+7/rvKFbqVhjAei+3
ooFWKy6AD+44jGPHwf2gMNPyYJv9ZeSqGnJh1LZZCyMaHYL/fGbX6dp+eDCDXvF5efVzqaGNtgNC
QMVTYs3qWMHoGJ6+naIWewD5FAD0MaSbs+s8CnvvBkyZlBZbbLs0xzPGraPdEDbFiveSLCMmou9f
PXeVFwx6buOjjqLoQHAV/HL1qBtEZWRr3ZUDgCyMfIS6zeB3NQD17NRQzb/k42hB8FGza/9fEi2U
RQo09xDC3VSMMPtRWn0bZj5GQ+6eqtqfyg3DsJn1OBTY39nIESwezIqyrS6Zk6UgTQAzuZE5j6D9
KkbGA4RUKGnLRMaoplXn/0ZfHqqLE3v345TFG5mO6tKOAqrAOHIbzlSXKVquvhS+nGnlE6nZ4kof
0dzb4l9oZTa1oCwNfcZh7xrVsrWXhfgXFXviV7N6tK+8EqYBqfsPpt66veETafkvzLQ0GSmSyOYd
a8i6OY+sZTTFJx1dDQBw9tYPcAv07wzSXdgNyHh6X8xsJHWG3dpYutndwldFVnVsQ/RYlDziDSQk
ikgDMmkWOskIqcgWEA5Y9fR02W7ynDDa9aFuCkERWQJ19Ek8VQiadaSh9AjAajD85NiS6ZQZbN6Z
kqg7ZdwLwN4mdjMBxj3gyGIDaDu1x0SX8KbpUPfflp2XToZ+werVxpHdpPqIolSF4HEXXmI0FCsT
Vw/xc1CSZIv+5SWvF4nmgksMWz43lWjJh5pqmntqVwCYdbjOo9S4AhzjXrPq3ODfwrnSBDxsZ+uV
SzCt/TUOFM/mYYb7bJvGoRJkbu25vuR+u68T8CGrqQig5NmCpN4BnnupOV+C++vNs5bbPtrq+a4n
VDh6hnOOOKkoTkZH6XIC56kTWQuB9qnG/PPhHqsaHqCyO9ZX14cFdgn3vXT82vMjLCQ8lZ6d/Zy3
4b0NXKONUX0dTWjABkv96Ek4OKRwEyW7sQt5jpcItKzSUCYiyoc04QXOAVtXA/NK0TT59taKPQD4
ATHI5xgo4DRzIb9U106z167ActRBL5Yn5ndFro3OnO3YekwhuVAdtBTbpt+U59FZwp6nrpq7QUZx
OAdlpQv4bUaz3vqZfxBZKsymunSpGkSQSqWp6XePqXrwF+NcUr8w1fAn0p+m2+YcsmiGfX4bzggJ
UH8Xw7lSLe4VZl8ymdgnj/+kaGxcVIqgGXtHPBanHs+qHOYoMOfycC8705lnk+tLomVtBch+grm1
dhcahd9dFFeLJRSiuBEC+xwGzLMtzueR82j/ffPxIJy7d9AZ4BdH/3/3v0kRabILvez1SwYqGW7W
asrP0h8FcOBiEyxpjBdXp+vKIn6TJG+6ck8nT8OsgBsOsGblV4bLdZUtqXFS3T5RzAPlD+YoUMPT
pa8RCw1+311estEAcCJ5JBHo0mZhgnfkYWnggyfqlX+qWBYD7x1/5ZlHPXo5OLaQyPYSjeePqGEY
XCU5lof4Is2kOrbgzd3SaWbEFzVy47MCb6PYK2fY8S2WhEsmyMYpTXVmytUPISXPuWJ5CvcuY7Vk
7zK8cZ5Ka+V9/2LpWi/3hxB3i5KqOEWzzLc3rRTMZatxG6kvo4I/o2dajtWh90pCltpx2n06sQdl
NToIlD3tnkGzgV7vZ/iVWmhHfTncdyKbOgqf0o0bgVdaTLFosDUaaz7f4uKCwwEhQXKtSeVXkkd3
2CLH88wgG/6/ztD4qiOUWbl6o8hO6KTzAMDdlNECqeZ0xq8pYVpgJaMP7XX5RbPx+XsP1QYYAfX/
sXqnFzD4QcME4N3VaRLJILYfUdneVAEbsm6A0aCO0+2sbKIBZcKKfjnxH1JUX+e0fIOcBKot+UQ9
uUhUKXHmbIa7ilR6C5s4/bDN9n5koTSVbYdmZkqCIYtuAGfoeiLBxKr1agpu6Y2Hge9dg35CbrwC
NLzo7We7s0kbE+VzPYKvlns+8qDsNfgRD3Finf1N/dfRMLNb8SmRFHo/84T2zxWJOzSkIQTqEjUN
HfbBUo9wVgSNmn2cFU3Pbd7ioCApfJ8EFgyWc0XFIlBMmNCXtZ4ApGnk3HxgTErQkKtgQ6iTonQ4
PQNo/sB9bj2D4ay9Ko8CXmPbrUMPdl09QXCedOhcjgv09UpDY0o4tMX3vsmREwjrQJDxTyjeBXv+
p7IAJPwUBQEGVmytKuPsG3KmFTeY9hYCbaD6tHXn1YKrXRyDRCcQkKOfaI4LdAbCGwaFVl19fKpK
vaOE7Q3Y9X0THnKkfvNycVPykFpRo2Hj1xfCzJeTjRaJr/fXo4OcdELqd7e456RrMoPSO8Vvjz4A
krE8aACc7w5VovHM2odJSAs/4uvzquKW88jONxyPZw7ci8J7tTRo0LrQ2l2Hb6ASul1qf5tZgHxU
kvrEZGsgtJEgW6U5Izx+Toeu68J5x6KPeOk6JePaEnSmmJcz8U24e4T8gi+HKcQondllnhxmy6VZ
1jNIwLtu7Fi/5RbL+xhoeGGYfMJ/5fFM+P9ByPVX9OBiVND/+VBQ3MdG2hV2+DaqsGqwQpd7KU7x
MzdJIiGIK5S0aOcWDoorfz+BlV3WgOasMhPhkyrfct/hzZG/GqIYnelCYDqhLkRrVf1EPWu2QHWe
caMysuh6GYNjsiT8wEQK0jALsx2qO+Gr/QnGSU9Rm9RUNiJ7mes2HweheZ7ANbXfuzNB7VF+V/TY
SJQnrYjZfb7g3M3tz1/vYvQ3fxTnnVgdI5nt71a2uXbOZyxBLyEpinIkI/0D8Ht/bVq5PBSeoQAu
QW/s5827uRZrD92dPqXX8FxHPhA+ivkVsv5G8KmKIIx0u+lubDWv9pbjG0XGr2ZPV7+c5+DvVpVV
XQ6e8//5GdP65m60Z7cUX6x0IB5zWmGIbvG5whqjr3WYD2BH6NnBMeSTvkgXtgWyU0S4bem+Ho5H
yBxwGjw7oAAT0YVNJPxroINGQQBg1kY7WNVTchwDN+bCcHER/NmpGJiWCEgLTZbLu1sLATvUDj/R
7SahVOwHkjsSYnz0lRqGNqSGAOenu0WYGliMLueoos4Z0CG/AP2rZHva3COW7DGV5WnvJ/smtRS3
dmg/v0Mxx+6+i2Nl2s3SL+L8mG8JhjKRpWzeWhxwXeYxMPXwGW+ofgpYL7vLcr1DyxyOmlTgOuAL
/Eh5/vK9hIpKRHOk6Elgz3uR4zeAFWDHHGiQ1ecClLvh1TMn8d/IIw5V+qJQTqshnZcdOyIzbT8w
WgDdFCsYa6Zja8YFCSqgVl99QwpS/2cyZECkn1rlj5XHywpRAvswtuJ6Ov4T4IqDNhgHI3VkGYjw
e39xojubA5KBq54Qb6II/E5ttmbxsls07lgFLcqSGOGtLuiniYr4MaQHsDHfvSyAcXyleT4tBxE3
D3/XVwflUF7bieCQLtTjT5jlk+/aZbE/1FtB89X0hsSdAFsjTH3hNoJ0ITb4LUVUf7+xfYAlmMF8
KC4aLRrJNXGilr5dWiOvxq59jGYkjn9iMiU3RS1o32+RJwOIUZQHaL6L/ycUpwl9aoGjuJ8Hmhbb
+x1QvgPuX5+c4HexX9NZq0B/BEF6gBS3GL+3Ls2OfjL/dcsBViQiHGklPvGCGscAh94g615LkCLg
jhSjxFPo6m6s0N/o23uX4qJ43JOkeFmVA/hGHrrNqL3xpRA76ZIlYooe4Im/UYQ2YWEiLNN8KldS
qmdb+n7GUaspY1OFvBl+caSiUIFTVonkKwSj4MvCqVKmiic9oRKOpfJfr48BjgLiw+9UVBS9dtkB
ZzN+vC6IZ3xWKXEyHZp95HXmd5JeX1rkRzwSYKNP5Kq0DgW9NRqQgBh+kWZzkydvjOw6k19gtQaT
cFvpbZFhgOLekalcEdtCPMleMM+etyQjdEhDwLKLXCVwV1cRQNOUi4TsG8fibmE0j+5TqxjJLwti
L4wK8KMi/o9ZzxCPVTbu7oPIyMjAslD5uGUeLpv0PMuY1VsvPluMdYHNpXrUREo0X3wa1M1oMBlM
m49yEBJC/WXWI1iMB8/2Q4sjupr30vA0GDygYRqXjxDQfAazRImjlNR2Qc2IHTkqR3uYVrMcIZ5a
sAhb5+LrYY/SyzpgokXi7/UZS0aQOOkzsqqOgf/aHdJZoupInGGCUFBlnAAmx6/nN4DpqUdfyaEf
kDh1FkTUZtcLcGwsvhrRSJoNWbx9IM0PqsXpvu2yiQnebeRcLbfKiEjkh+uqbl7FpwJvW7iKSYj8
1q29jpTM1RlBgHyOMkDGYKcqWjht9b+EVgzxDHApvhP2+Ffj4Qhqlvp8bNSHPWW6w8wln+S5Q1P7
E4TqK6nKvNo1Vrq732OecZ8jEJhmZyjdNitiHLevxFiPwZuR3GAyK3CVLRzF2ANYF4Jhz0VIeb2o
5o+eUX8dVg0Z0nZc/CVMJJ66Xi4FQMeBq5BmzMffeOJn02Jpyher0/0eYkztm27riPemK8O9ocFZ
gY7i7SaJs35RFIYoSFJG+NZQ/VaHnpwmSnAg4MrqB3CEVK97lxpKZcrg6Y1Fi9f5cn6VczRu4Nm6
ig6pldZDzJY5cZebjqjWKCmMqNGL2yFiEYno+ffM0Be0dQhQUzjOtnYBBklqC/U24S60GYEUxc09
05uKsP1/RMRqvbCYrOYz1NaU5qKp+l1SARyLs2O9uauls7Fmvn3SbwLWtCNKrYwNIr5KgYLai04N
UBGkfAlIW+If8DylxP6NNRGmudZSgtH0jLV/i+69Y/3og+2qG6079wJ62vHbEkfO+lhGx6Uzm218
DmUabq0+R+sSxVsiE3dXRYejtgvQGIAVOFwcOTaIUmGMelHz7ehebq6/wtO4DV8cMFOKpQ6WvVdW
U9KFUInhNrU9RGs28zs2X2kojw9dqCIz42KLSuq+VswCEzNLNh4bcSnYLJL8LpIwDG+WpjkqaVub
9yPwKi2UjPzqIuVBWxCRY8PJez4Wt8bH/aNmfr9wdSVWglISH1nTUvripFouc2QVGvGo8jLuk/h4
mbAbMbMzLmjSq1Dsa5zt47KuRTwbwzffyMCmBv6vYPf5iqaN9Fa1rzH0jt1epzTb/aDINttmvXDJ
jWigmWiedrnnyDL8bliSSc2PqYjxeTo8TGPLweKVGWltHwUDF0x915+7jCs/87WeLgWtbLRcBUyE
e/arj7Sxs1VEl6hU9szh7Ev1jJfeTymsjoEHsrgr/6XQxy6plLpbO5Bs37GGD/tpL9POJ4GH1yOi
YMwab+/5A2ZO+dHfRZb0qtO0b2aN1peSdgCrGiFF+w4f0bTCX9NNWbks3aKTMtasxpq+acPQDvWF
6A7twCUVTfZOMpQ8ElXJs1nTtF68q06cJLny+l/d73gYhGAmHBrcWMWOwaHuPx8iyWc7GFmySEoZ
SWVqW30JzrxT1U9fubVV5eNH/NPtdD5uR4J3604ozD8q4ZyMVx8s0+seTEVW651bDVjzZpvB8HgN
j18tPWdpf/NE7kHNSBy+8IvESh/K9SpZZ29VJoQVf2x3JfV/Bule3YbYtrvIGNAXuunGw/Cu4Nmd
y7KaQm76a+fo/pfoA/XJdaCC5A3QWQjHCqztBhwTks9FC+VY7VkAGFErAoleCZt3czssf8Adjbzj
v56XWVSobr3Cqn3deg1hslzoSxFtGD1YvMKACCHY4wjH99z1AvnEWbQtnj2Wep3xzxaawk7Npfmh
TYLfG7yGzgoypA7RS0bzHqoS3P8WDGKb26GqgMu5ed1u/RQZ1ClCW6Sn5lrAXgEX0SEEXSmxrL0A
55dshShnHb15xU1/FP6fS0c7tNBm7tV5n7eJcjITwiUjUTMQzVNLBMZC0F3LN91cyLctwg/Y6hwc
YIIzRO+nZfGlRlZnmwmByWhTZt8dRNWpmzpi2sMf1fG6hlz7agetXtLIjF2fjfOqCAlr+ujFNWOH
eT/zvcu0OssgIiZhgCkPB94g0FmEDaRzS5xLJJaSJD9LxeywETa4foXmvklFYYOxZON0+CQ1G1I1
8/5/fJnY7RR2yumVWo907m9dzYBtbKQLawZ9sTgqh2nds5CX7tLDEBlFQYGDPXvq3lTrJzo8u1TZ
xlSqDtjx0UKn38WsDt+DnFgBEt9bWtYWEjIrDQgcI7QS+6JcErUCBBiahJ7mdeE/eNNjEsTcWD+j
By0CioB9GGzH/oZMRFjjXCZBLA71vzrc2lQEJPflE5M1LhDRKdFUmwNfnBZys6ke2maYbu/Fn8l0
3RDnAAH0O4A0QHEElYzsmhWrc50cHFa7hdARlbcKNIQ8fRbe3SX+qD37M8ovqPB6hSJLqvOkDbu1
9+DlFF56O7JfoF9dYOLK/bX59pQrEFapnl0eZ8kAVP+MlldX2IadK02066J44ziu3SWGABN91419
7fGrzpy3JH1cVjfPCj1sM7hgD9r0lIG7ZkRhM16XfbCDeiacA3h5QV0PfkM3mE3qsMCyThg0RlbZ
px183yGW0DsAr63qtA7jYBwSJXTqpt5aOXqlq/DkiSlzttUeeuJdMQc4q+GuCZpiQwlFlNa/sMDA
sLRExgBfCAo3xUB8CDrQssvcp71WIJ4FPouInCAicsAQdKbjuK3tHaS2gvCG9YBHsucMTGjTyOZR
0gd2+OFVhiueAwLstdBqfMIqhTj+yRo7c5mUxIHfYi1iebDDDL0VgbTj23Tcpk6DAZOCOQg87vO5
EFHqWGzIX8tNRiHJl6+LIxccB+Ey5OYiLakeuIurIKzdts4r9frUFqxANUWUdZ0GpUMLnFAGzH7k
vXEUi16vg+Qs0qHT1jmrVxRj/UvCHkyUDq5KJoVhWiLybwJNFXHvquQ/r+saVwDttPvHyybS4RHZ
JeAjaFsRfTYw+3dGyPaTzPwembIfekyIWSa77FtMMcuTOb+sYfNG1KZejEcWKO8mli/UeCmXr02z
6/jf8Yw6bPeTqIJXJYfIbrbnYZktP8/x88suz772EnlOUPT94wSHWI8+IMXP+a7tdOB933aDpfQF
s1E5ySvlY+AyxpLYH3WhnnV7RWxoFAb7QMtM/fuhyxkRiXgz7yg+rwKMos5+U47N+WU1puiGuzZG
phSEZJqXGoA8FoVedOjlOtsgxTi/uTSeSa9Pbq4gJDJrdGWAtPdaOx3Yw5IkG3BwVekE1J/mG6Ap
qJoFRBfS5bJX5Mn/pmOZ0jZq1MqTUSDUubG0RKPBX1a0evz2+7he+khI2MNEWyJdigy8mYYgAiwS
gqjKiSiEqfTx4q90pC4lArGBfUydgWKklWMlliR9jplU36dTa3J4nhtwqt3CnnmFPzvXA9lK4iLt
7Pf+hhd3hFBhfXBqv1zyoGLQAjZFRUF7wAaxioiG7JFuACuhMzriaFFQNSWMxVqLtTIMD+EhrnEN
idhf0mviUguKmtx/0pov9mDsFZ7d4bLyxv02hquwMTeapuptpcB6Gk1k2zvpklxxoJwMExabMJ03
FMgM9/7ZkHt7eGe6fEO9Cl2NDSLkzbxwEEPOmhKYSMc3QQSwnnG39f4E5S0V69aXPPq8SLK8jr8V
nj1MlP/tAR219os5Du4p7G9jYdXdKhqPkYYe8+Pu9knNZ0fnPJYbWWyi9Jh1S3xbjpshAR+czPBz
GfHQ8IsPWLgHxkjOOzpy/NFiq3+PFTiyHddCufKycLvgdETkol0zGPK/w7E2j/eN6CywUbgdSsVP
yIFlbWA/LpdR8iiI+TFyz41/yWcQHOL7pVBHgk85p7W8rbY+9XeKAMulmyCQQeFyCqfKtrTaw/8m
t6wUbqIRF+6T0kgnPsfBjW4FfF1oZamVOtxONSure6ZzuRgZ4eEMHfBOKdq23FLxE3PfVz7GH0Fs
cGiDCVnDV9cpOWI5rrYczr2sn5krvOLr8JpugR2FkyRbYDPkb/vw1oOnuFv6Xljf+/m9LnyPz6cl
8C6D2MYPqSNsiHax9QDCunWQRdXAVJwo2vVcD5tRD7ewqeSZ4X/tTl3+TERI1/Dm3PJHiAri+1xA
KtuQ9Ji2/NQyee/WnImdzXr2EAHQJpSo1i8t4RonHVe7kiULY49BKsFiBdMILIx67F/IIYG4+WAB
BXmMMMUyF0bm21R95WXmXwD0rp+diH50pJv167mYdB+XDmiUSs8c4lLwBEOQe7JtIupgyvHxp2JB
h/PrfQhGKusU2e5miKlqUd9wWXlD8YXQlB/aPMTRmBL9WS3exAxNy/8ItnCeJh9H8bsXVAX0Bv0U
/Ah4958UJ2liEoCzKnSAmoztU/jYLBVpzFmDQN0c+IaZNDPwdgK6+B0M4H8qAuyGZ4v6RkIRnH1t
1eVfPfat0bTyRc6qwsGyZqeHzpLHCjKicT8uqebFlhJXm5arfIMW+eQCn6esG3OwPI9A3DVOr1dG
Vgem0lgJb0QtXyBpY/0KFWv1rkwTDsGuLPaSPB7KTPXGXUhZB/Wp+696oQ1qmXzSbqgOG5TTAR4X
skfTEgZr627vY7qsHveSYPgcQ0slnw4W7pADXE6Pl+W5cfXuFP4HgsjcLNRnWgyi/HizwMSDnSgw
rp4r8F3AK42gas+A5TLfgYAbVIO+0TeHKw/qnSRD5rYRyaDkJ8ewQCHjuXPlN5ZTo2mmbbO667qO
gf0apV5fIlt6lGWOhoDMRGlqZ6p1vkERweCK3uxDGtwLknbHjGLK4V5i5kCi+h3X4LSZpG9uj2b8
X++4UQQj7VaSRSwKhCroPdlh4Dd43QBQnJ4bC+smRgL3OPpYr75DMwtEVWP1JjxCM42rmBZ4Toby
29LsFb5oMgX7mN1tQ7RjSAhVD+zp4QaIcQ2vW65JVY1hRkkzIzdWFJSzsrKC8zaku7sH4g9u1YKQ
U1MwWtS6SShEA5AjfSY/y7HPtrQ0EY5SYI4z7hGnHtEXr4mQVCG9717+cQOkiUh9VpNxLxbwQXao
QEIX0vHozimrEuX6mtS+7A9/0TumIaJ506kZ07MiVP0GM64fzQVoh300LG/cNMDc4RWShh5iOtWb
59DSCXUwxFUNclWvD3lqbCjYFVKK/wXN60L9rFowDVt5Qbiwri+5gzOrBM3N3pKCNd2kxeLErRk1
Fg0GdhS+0a/y1t/W8FUVvA4c1nahIk0zV6jZSTfWadNrBlfC8ugseSmg7ihcpQFfnQTnNXoyVQI6
P6FGcIfctxt5/LUYeGgvxzM26dVSu8fFqqS9svkDE3IkJAXohoMgPvO1G3iRlbe19bN7nLMZ8ZDr
O7Z87vtjXzNHul4K17iWaRcq5Qqm/60T4tSUeBbJE5qBO8/GPBGNLec8kMHrIHAfCNUoSA8965Gw
Qc2BnPKU95SQxnp2S7vW+ixm7jaGPcDwyPztsOwvFljyxilNwEIo+RMuDZhxto+M+/eHbI6PtA3S
GL5CNRZ8LptlPh1LM4YwniSGmhJT7UmbuP+6S0+yH4IOse4hExUj/1s5nMimwLiZaUH//73KGo1w
nVxm8UUv01jiAo1sV7/P6PAbIOJNUkju8mfrxbg7mguExHxF5XiGE5In1nkgGK9kDVZEgOIgJqg1
1jy4xlMK/gxBLm8tnp1oOfChDt85gMb1vlCHxLZIV5Wt7Nv3xL+wk5Sl87mDGgq8urm40Hj2E7X2
oFFU9+FVhdPt3raN3DfJl6MNur6Qzc+TVYhrZwzPg7Nlu25QWoFk9QQOl4J6SvJ7bYAUMMSKFApR
aplZ3emjKs8SMYfPf1EuGdgS1UWGr2T9piHDT2Gt+ttM/cAJGmqn13PG93DNnao3B6bfuLOhkcmd
Ng1U4jmq2OWNuXZ7Rb0XE+9tLpyz2KDU968E8efFNWMBo05+lQII25+HX6fYy1O9EAwAK1jSl7Fp
h56++hS3/JP9jhI/YkdppCcFuo990kAdN/fb3RHFugpQS/uLAQ8nSMwoPlQc/GkyqGxuqIzdKrwE
sFVry4WtfhbZ2JgQrlVaNGyAHtGMm6rlJq3fbsuZd7jHckiJwNjIAhUnCNkDo5OPeuZ40FnbwOB/
rDTYcUjUiOuKbzbBrO5SjSo/lzyhZiHMBg8X6On1XGKdSWIF79UAsZtvvtxnebOn+2DCKy3gdrDy
j4dtFayiFbavwpjCoVmVenD90uc+eLiZSa8D4ZZe5XuK51a5HshOb6PCnJyXsvYoSCdgmk4MgrN9
siMN7p6lFjSaL4l6YkVdjmNLth4sbz8zek3u/BJDTvHdhaXCTGCjMcpyVohUk0j257lyESC1R4H6
SJBOj7SmajdOJdNwsdW2Q3+04/Q7HkiBhl9TRsLA5BndYvxjb7R6QwXAElDuYhjClZTqfxJwb/ET
rRGUkQB4EGLuG19Y21KlzuEFg4EzeLBuq7AiOZzQPVKI3XnawliVEAGTxwXdhd6fX+UiA0WbtXaX
ZhJWbpDJTH3rtewXTENH3QIiYb/fZ6jHVdssSfIo16wv9rl6Yg1Ge69etB40aZksypbL/VBPoFB6
5MMP5n49cBcLwyBJiYdfwJVJVJz2BbmuRNd/Fgeu9v5A85jpeGLOrkKf8rJGRbYHoeWNVWDNDY2m
QfaJcMMXgBD3QwcTbIqkD6urMzZ98+IVxuilxkOvtKpfgjsVzaM6OB92c9X5kg+izsmjR+a6eIxL
y9uy2WahtBUkjMRegJp97IS3MhLWK/f5l+af+7QpGEVg/zyfpg0uyhFaufc6WfjkdH9/EO92kq3G
ez0Bw227VSHDwXxPZOqhtCT8aUJ7foSoDXkIMVWFEa4ymI6XQzYSrP801LdnM3JNgK025vpdu1/N
IizjwV3ffPNR267/yiwmOBbiHGr5mZoF6F+8NhIvJ8WgxUUnULcY9mTKlJAu6oNDAB2ceq2IWRnn
X6MwFBFzckBxysnaPvRe8YF3/lzAxB5ur5lLBg6hyvRlFfhvviGIgZHSF0TvzlvINX70e9YFNtgS
9LwEc1503CrORa3X5SJCDsBwn8Emv0Jpw40uOY+yKClDtZYCWBnAwQxva4qpvB/Me/rP8rEBlNE2
AUeo5sHO8AeCXKYOM9ofZknBJrkvBF23uV6ZFNjt/XuRe0H/js1kXDzDkFaK3exwLuu8qXuE2uAK
N0DE4HzyLHPAk3muMccQOF+6LUmckY/OzKMlEHWcetszYbuQ11/T18R++/CH9NUml74Vz7fllQA1
icuUvZG1a5LUAng0eGcQVzgGc9LGDBxhAq379GiEdvIt72n3ggT+0fA3kFFz0o1HR7CNnClp9uZl
D8tsTfbynHvLIUUEkK20rJk+odWyEKJkDef5VZ8lfwfw7xy0ICmWhlzCLZchdb5YQ5TVit4FNqdr
4h3GVTkG9sK6XnW2dxFFV6dySG6XDPtZIbZFdlARlZZqMoe7gZg0WxYMHSpKKNTBvtgDba+TuXbs
041233YNF6noJUl6JY6kVm9fyq7CvCIlgssLAxZxUQ90u9ttTwr0mjf6QLWXp87BHdNyJ+08EDYe
v8WF/nESU+9kEr5xlGAO4W3SfKUTAfzSn1uJZacMRLdNECxbLaGwKLQeAjmbdwH0TNfyyx2Ojlao
pBc6bVxb/jH28wqITmiTIzI8j6waEmVlD//TEUeRm4b9R//IfOkhGwXKyb5PbDX0q6N4AYTdhGV6
vqAXMAIHnuUHY97eo9f9GODyR73Pn+Qf7TEv1gHXokun6vGKXMfMIO7o2eArDPQCY8yy8VIkjHsy
9wBK5DyJqqPlc0CGyWwotmhS0rUN/jrm8D0xe5eiEIDkkSUWv+K20zmuhKhSJvIVQH0i43hnawqm
2jChOMILrKsCDKdBGtRsJBIZpZwun3tU2nYrDXO8S7xJ+VhEk3ct0ncDK79vS1Gb4FiABoziU8sQ
lMd0+00ickqBuKH4LtfL1KcqL9X5KZk+wbPVANPv2dh4IMDLwRJdRXIJqbguGsZViYxVq9vtqO0n
Zy9MnvmtUYqbS87zFQcMQTJUb8cb8G5Cod7x+IgQPcH7jT2x3ob4/1EKam4Paz81qRbvGMeyg9s/
4L+N3yBJXLc2AQhzTyrEB8PUhrAMaj9W0HBMp84m+5b4Eh/6G59my2Ym34/q1jnTeDzF+VyqWpjp
MuiqdiVOrzvYSyOhJgiOWHubRs2q4X0aIuugOh3djWYsYEwwt2ZsY3M1q8By80zfeEwU4plxVGUo
7WUNDhamJd9qmjyK4tLosPhcgSyNFU0yDFTdt6nWJens9hAASqO5axHgV0HLG39ianlqSkjzg9y5
An0sjUpEHSGJUqR9U98iRR4QMYA0IoZAQQgbyyW7nz50O3Pcvb5+ueKQVpDj/obFEHpJn0ByFEUt
2cAlUyJTPOYNx+bj/4J/TwAZtRkuHtD/V0VxFU/303vR5GXjXg/Bgkg/sdo+iSxN8bXir7FGSkrQ
c7CGLyn3z8vH7mAgEhElch8cvMghT9Gy23+c18iOb6PtS4e7AgvORA9xFcp3BFUwBa/rXrSKn0+k
iWsMkKfbcRPDiyyrb5Z+juSDb0juf5pd9hKQZxPMfSJ6eILkATHP66kCWmhtQaYhKjUAGGXnCzwh
iw2S09nKaKRVBYKguuhpuflPyk7E5/kPqzBtyPcsElLYm9rSetCW9vyHnvV6nYFmLaSFF1dprBR8
YCzfFOFYdKJpULcIC3zvcQDPnF2Im9RKhUPr7wa9C2STl8i0ICSkpzidtob0PlX1kgUQE3y0PLcm
CZQDT8VuwDzx+0tagmhVWt+IBzfT3qxYgY52Eo66l7MzQihTT5cTwjqgvfu8yV2nIb6K1nlTW7od
RUG8uWt/yNSptNtiC9LwBxnfiawZjJMrvsZTC/a6t2xkpG0eKZfe9O3lcm9ZEDZaqkzHL+Pm09mt
qZs8ryiFhIsEyvvXePuAq9rIUAf6csd48Lw7IWY3QIafb/8sSOpdrMjb+dt9/D+jetiZIVcIwFjM
+Eg8oF9+DPsqKEyagwjlJie5sF6oB6gbbn6nykVmRCz2HcuKw5WXFMqZE1AN606Gsr5pLChU2NQt
pMkTRGGuDIfJJBZHwG+lQVN/X7YQ5FF0VaTfPF6QxmWVm3fDou8NYHIV8Wynz9TAye6hCAZSlkpf
xJCZQo6VhiIcjoagPJvrEwcN1S672IOEmADj7laYBfFhh78+eAQqJD6cpi0mO91f8VO9XsQF8V1s
7BMo5TaH78DsEAAhtH5ozXV8i2MlK59a9uvq0xTApY1sLRLIq5MWxBv6nviX0ffdoyjqSUXAkStu
alCw5xP7oFPg9F5d92iTse5CnZdZu/5RcbdJYToucvG3iSM8N/L+QuRX+mjLsHvBeW7w/yFi6WHW
LENsdR4yJlm/yZcgp8ajaF0JPWRfQRLnKIRSp7qSCWuvGv7gMx20D+FVPYnMcS6La5o9jM3dZelm
+Iz77IDE2NJ8/WIAeMTV1iiFSKh8DsHP+hkmFXn0ljTgAeiolOQ7KO7YwURVPmTyTf88yIH75Hzv
sOXXohmQg370Sa2/TYu3ZAzIwcxaP8Hamm1id6eU6GlLxFYqPlf6VcAK7dpkWxBG4fo532p0kHF5
rVwB+sWj5YQF5DQWXm04qXS4odNOUPxachSApBd6pQEXtmqOWDO2gYrYn8PQ+7pYcZ1DiyviarWA
vscg3bCQD2YoMVk5U35/NMnPF0FZDgaF0FwSeCYfeFQzIjGHuKvdM3L1Eaj8MTpyVF/NcL6WATSm
im/Fsgst321WkL4LqPRDtEnQH2Ul/5nxONSbf7Gddtn3CTVNV2mpLj/m9EKicNR26Xv5G7tb8b2K
kDSpUkvP7wxvNgEHltBCzgcSal+1/aSq6HfbOikGCDiKAFxvncGBhqFzXKy1fXv94uBYJ2mTQsCn
JT5RzOIYBkIMgf8k3WRLHSmqowMaznnWi2yE2FtaXFEmah4bhBcrwoFDmQrwkEUmCedmfk50EkmT
WsR1qWWlnFhXyh4lGJ85ufQvGulMAfmQ+6qIL9oyLIRQUnkQ8uNrFHxJFNwpOIVXJZWa70nvpvT1
LyGUQS0RZmZwVcUyH1aodE1sqn+kElu/AamDQ97MjwaFO1qbgpar7eVAbXl7y6fWpp6ZNAIGqcFl
knrGALzzMW9Vj6EN15Jsx/VyxiJR4L1VOwbroU8I2JqSt5nIAewbHKW3hx9Kj5zX/AboZHS8orWC
fLKmq4KH3rX7GyQuvLmSLWigSzLeqPppD0deThIDlA5fq8pC9u/sMhSoQDjXPXnBYGlECZ4PNEm5
UlnyYcIpkCqiQ5j5T1XEHl6BK060QBzR4QWM05Y+Ry/g7OLI5NT+JVl4EzFEp5NPJvplCaKufF/m
Ao7oAKURsV2eNwGDN6JwPTwnpW8+5JM5ANXSSUSodvg/NCsd+wG65oR8Pj1AzA/dXNlZQy3AEN60
zptvUm9OCl6n8iKNUy/nH7dZLix1I1v9oyn0xTaT6zik11Vo9N1lRhW+TbgzjW//B7mQKxQatoB9
TU/f5w5UMfduSfco26WVVDEOnFHCVLOCowclv3IDJA2QWi/nvxXfo7lZKdvqpy6gW2PEuxMCs69W
lM3XoKYhlcEHGeZWFE4i5qV2Fhegy4zRr8jJRewX25pLyhSgpubOjGqdzbLKxOcAiE4YVFMoNETG
eS73b+ATAnCvZv9Pe3yNPXIvsjOO/LnOAGSYZ3iGWkMH5xRaWP/c1D5PXFyfJmclm+XrA++KyD0Z
p4uT0WFZ3amTFn23Q40qIBV20D3wZpxIynV4q2rCpFahnFaNBJ+yHx+VxerA3qztHMYrqtRQncjE
HwT46wiWHj9AXiO8BodLpoOJ9p0bfo2G8kRk6wdFLRbmmwqV1shv1IRC1T89P3kUs2xg+FxtGEnh
PkfiqXNFwu3eo9Psu0J/Gyfhwfa8TkM53+L13JQcQIuGp8vqmk8PRp+CIPjy796SXEejmLMpLlmg
aFOyzZTS5R4s80R6pAsUPFxPKwIFMHBW9MdKnAHkvDO7TgBHoYHrs3CIrOQOkaJD49duj2wd0jr9
lF2aW1R9pF4ifA4uwzCx5MSG8XmhArOaM6wAND/cF4N2ilLq/vbX1A7pCLoMKEmg7WdCI9WFdm6G
KV/M7Uh2S+jB1sErAwkwgCe/6psd0JX/JGHBGQpWczy/5QvEsezUbflaU4vj4mDTHL7WdNvZ+4Rw
wzvMgnxBaApEQAxV+Imv09BfcvVCi43Oq9dFcvP+RieVLPAm/JCVxGh1GQ0OnQxXaTAJ/kdkve3i
iCduylgbUg966QQsRUWkly2ZJqXIzssdjk7AK3s+++FC936GnB7pSjy3fW2GLF2ebJ4rp8arcsD2
FA0bTpy0kNrJbWQsEmtTqK+wAwXsSKo4JTQe9+YxG+13LmC7T4ygNqzVxO2w220e2jw5rX69HyHE
SmOlOTaunEM/ZUu3loVArumPaJ5K5VKxu6BOYC2XCogLe7KH1DPAtOZ88AePfgM8Y32XPBBhwaxX
KWoDb2HxXaOVUG4r2EU9ktkfoK/goNipKjVtpIamwjiiK+GSK5mFgEWELFxYHunnYEdSum4a+5WR
i7KHeZ74def1U3YTqQV21fUwV+j9+Y0CdAEC6e309b1EsFn5MZnicfY3+d04b8INRYYee8DLQTbY
R8rm7Ll6acWYTHxjyvCsh7UjadsR4z4t05by2SleQrePwCWO2Pts93lCqpHxZYpGoTWGghDDDIGk
seo9pJ5G1tF4FCbQ6Dmn1fT9thDEFE1y2TweqVh/rilrdzA1o4PVf3fAZSWXoG9gxBBc4W7YNR4Q
Ww46ANsSfLol1hBVvh7V9GS+I9F5gpuI84I0R9NExOcozbUiybk4fYQCWLTOCZ1H1KdWjyKjlqfv
AbJ7Q0bo4LyBfvYXrOw4Vc2B7sQzB27AHKtnyhj+vlSUpjc+KTFjV+oza2+mWDhaHIIveKvF9F0e
VjsAZOhTw2UobHF1GknEYydGEySTWD9reqaN+HqiEaP/7S1NNw18rjc4O2wHmeIok3NczQ/pUaHB
yqsIo4TUQ+XVR2A3Hx0dHzCyJOXzghtdBjRK60EzIVTmP15dX6QnhzdO5rOJfzc+1axj0CtnZVte
IJv8ycQIkBeFFaXzr9xudUsqikUFULve1CCRxW0c6D5NH9D0q52KXJx2s+m8i7NH9EyxTA+eKxE5
0Bw/ogM73iLWCmBlmr7aEh1funawYhUr5Q0bE0+v5f1KApcgHySj5AOgMt3J07ha7RzQZxyYtBjK
fxWkW2o8yUxTupUmIc3efDujFxu+VcOaAGeLsUcGM5Ax9MTjTE/psttj+Hh3slnZeNt11hMRVDy8
ZYr/TRLtwCSkigB328hHiMd74SQJpqhzkrJUIcf9mYjIGAnKirwDkvESRlKK9dJos3tq/0l0ueny
0/PiP0+G6ZnRiFaTzmi406Eu9x47isV9E3mTqbDO1bidoC6Kzj5w0yz2KI4u6RhNR88NH/ZTtRAL
ainOWIvhJ4luMbzG48QTt82oep5PNnPLfo8wunjzpuT6HNOTTiXog9V5qES06ry3H2NFGYVL8IJJ
G+dV+kYWzzjX1RM1oQHsjVp88b4h3ikAN/RfVXkvTixglsgddx0uJ0tyAH1b01r3ZaGtVhrRGrm9
8bYFpaDtLynLoUx3J8AeidGZPGOOzBHQVlRuSiVXGG5SK9fw+Zl8G+WHcRt2ecU9gOTkg60tZpJm
a548UndFCjCThSDj0hH4sm4KE/P5tIf1SwHDSSWD8A+pchr761U9FvcU9anPTb6oRlAPCg8fq7wO
b3SvulefR8nxApm2nYpZ//NV7wEqO0tFJSfA11QwJURRjO22AMnT9j8KwMZLjSbTDRZT7TbNPgbh
Crt3hlQWyvnLB6n8cC678EmsfPQgk89j7EX+oAwTdrhoF2HWQdvqE1NJrCbQ9D0Ya9yIEW/mzZPy
RrUX/X8ie8gF24J7y1AP4+XBZhSKlwiLxl/+cVyFX/imDDHyvwa0d5x0AFcS9rxaixGBrEu/tdCE
6An5GHONE6K3SUVj2Ea7ei7zVXWLqh8cm+JUKIDvnAOc+/xuuS5HqBbnz8JlVEu5fgHn3xD7VWPH
9iImRqrLpe+y/v1ZTgMHn+0wicKK4F/5d8AA/gRt6dh2yui27F1YgsCdsHFq81eYgvMUaTabQawY
HizDfyWH0q5I89LYwBQV/BpxnL4neG3Tpe012d1Mj6+bMxAz3cKrZSS+dQ9ZBKM3B7Ii0Wh5vANh
gUhddfszWLk4qz1lqmuVmBEcPVHlBYqQjYNsz7Ek9k82RPmTVEGjxNNjTT3pDKpkgpuM+ijziF40
s0uZ+FoXA81W9h5AANk87aYAQZrCQxSOsh2WXWWks/yozqAK9RwvL6qMmPTR0LAYnvyZEPf8edN5
9JfEAYmYyEgH0ar3itzjDyu/H5epjiriXktYwX69h+ddXhpTDjFFS7Qjn3gWH+vvn/mqL5kQ4jWN
DP17JcBXpkCl7EKycMuSIFcYrW+2i+dYCKt9K+ncnXZEFSC7a+pgWjP3Mr2puUY5MtSIw2WH6SqH
dwxo9taZBj1fmRpGhOd5w8zMNvP1IgHORtKoUPjEbSKKjJTh/EpowBQT7qyOKVkQqVbMf7XRPnGe
qMD5LFDxpjMrwybwR3G40aNDlEMK1wxehFGHvLoq5b7LRsR9FtXtBplSi8PSgBMVVVhaLo1nwql2
1XZUAw+cf3kGdcST9AWGPTk5ynWNL+QXwJa4GbOK2ymCHjMz1X0Qu0bjBouvP28euoL6+E3eb7r0
O/yyNacCE8nF3TNOr8F+z4iaRJhE8bncxOw2wB+IqWudSQ4JPs//Ek3lpG8TR4YGi5i4o3+4poX0
jbioZl17tRDJ9wSTjY8YjhuyV6hGavGzNYFEbWEWg1Zj0UCYRaALtbCVfqXrEebsOsEc2SZi+M5t
630xIx+SFkJI+eg9TivVoFDVhkwGWOguH9Gy16vXqcWHfj/L/m2f/Hn2mTN5uZkJmXFWHC394PVl
/+obd+xfFYHdhc37mSFY/hDpU7E8twFT4Wj5oMBsXy9fSiNxrB4VclQ71+h4ti9sASiGIkt9Rz7z
RnGGFhTjUWeQMVMvExFB8LHy1fxDC0/8561ucAmonkQDX42cPAHhXNG9+ftbDeRH/SXoY2yHbaWW
TvW6etiLmH+PsayjdRYUv6IF8T8LGCJUtWlXPm3w2J+4DtgJMF6OklZmztyPq/HHYbATv3Sxi8PX
RTtSoQVoCT8rSBtczSFSGGXsjsw8OTnAfCN2gk7jQa3OytXaCPr3SGcgNJAANsXYedM0uvHHpVQ4
pib1wK06rIoxMMgAONbO7FhmU61d26a2Nlv2gW6ovZ7Uos7JdbpGeKbApU+W7IULXevoiwr0fXxh
zhCmhtqov31+rxMQgfzUgx68a+z+UeBZCRZmiLl6xnoQGOpuqAsr/CL6mt5IK8mgXm1cFpq8dJbc
Aus5HkIVJnrPHYHS+p3TNvD6FQ7rfGHc30xFjDjIU2+BmkTNrluQHxal3R4NemtxmQmPOY7QFruG
l/4Feu4ZyiiNz+xs+Q7lKvmjIUmLEWJ7sGVR6J7DShMEGZAw/TNJqIpOQ+7RXWjmJPPeJamLH8oA
B648YBfzXWGksJKP5YS3BGBx/UdWzDLFQnypQ0BgAyuMQajdAHxpTapr6TwOvlXipmUz4L6htJLH
Mpb0Fct1x872xYl89AYkziaZyutaQu4fcN+7T+nQIXF3DaxdM8rOp+iFiemlw+zN7detT6RdEMqF
yeCoA9qP0POXooff/6DDK58BI+VHi5tpiu20KojfbE4ZNPQ2rrTQZMNvvJtn+eiwKsj414rof21E
NodkTZFiTTymJxZFnEqm/lM0gry2Z+VTbb4EjHKbkHM0gtJMz4q/KWx4cdtLJNRj+GH7b7Gwpk6+
aQyVbaT4+aSafg+nBFxDb0M5RO+mW+e5rsNhPDEHOdFFFQUiWtn2PPgrximM/SBO9ODRdd8qAcK3
RWi1zsimhKJ1ei4I2TUPTGk9pXX8EuC1GSa5ur/2K4QLeXIWeUgQ1dXrkCOZD/prfZBuQe1XW+LG
MH2ILKJ8TfA/KfxGVYC1+y5G3+3qMOEQH7siXioh7EIgRczPzy53MZlcf2OKc8mTa/i4ydxEFF+s
HtsXR2BwCAHUVTJGvw13Vggr5f+QBY1dATDcmrBqE2f8zMWSkr2Eq6ZjnPk0UaMFyPT1uBhzraKb
USaD0wuYV5Pa6QHaxKooElKOU00wncLe5dL5ihg2f+06SiMYCVl3R8jAx94oxAUH4tsa9St+uSXx
zmkhw4w+yh2dyyLkKVy2qrldhE3jKDTS/mgIzS/SMIglFHNb5uDvv01DNd59cf2HbvYqGUs/+yPg
5FQ21KkZNPuAKUW78Nl6C27FqMRC8xHQIU+TL+hY1U9hnRUDb8ag7mngkWlth/ldDg6J0/iakWVr
Vj7pIokYEic/RNusTuH9li5n08DwmB40WnpimuJQfBhWSwSME5skpHxX2Y5nImAm8KFvs25w6Jry
ULSNRlLpxFKmT+ufibGduRNPYZWIr0HgxvJKSFdymrJcOb4GoVWJiC4Vk/A/6oC5B/VgIQbiz0Ds
zUWp5JE2ksfJJ3VFhnkQrNGn1H2Ky5R+1cDnjZElfyj9jzoYqqnpb/3qJiU3EAbhW1gVih9xO2dK
3bZAsdPoTJJkVvVwOewbc8V5MWfGKYLb6Dt+EhZT8OAFbj9ALF7+G586phyllLLDzvNp50fv67Cl
6VfkqjsxaCbMKjnMltKKjm2rvrVnymKyucEWIYnzyDy0dTA7RkxrJLXtlN2V8meNutZ70Tiqd4Ry
QZSIb6Wv4UwJBYoHk+EW4MozYxlkP9/C0rME2zTyJJSw8PsyArlWvkNHnZLWT2Px2xhiyZWOYg7A
jFttdL3MnZzXdHoqLOcDSEF+aAjLl/K1+cNxv+SVwKAouAWSZ4bKx0UI1euapuUxJHtUMKT/vgyr
5iJVAHZt2Hab7wB+rk2rUwQ/Mw2v3ACDQnNyOFQ+3yYg2WxZ2/XjdfeIlKXoVVJcl+TNHSzymAZJ
09/5Fl3xiEmuIIOTikxgFVQIQQV8pH5mTA14Y1UuDWC2L0s2sG2M9TR3CHKeaD+NujF64BddAzO1
CjyJ3tSPMErs1fyynafv28AWjnqaGmV6QGVkPWGCO8OtqsRY53n3WEGMGccNXHfBUOmNu0LCvCdW
Q0dnnJXCwMpGh+i/7X7nDTbm2MAV3u2Az/HwNKKmsw5I3fVhDTYPkmoOPYVlc2LBO+Um+tpzEV91
67QkcHPGOzq539A7lTcH2DAPU16P7PY3AGKaSCFU8iznCO8w/9YqfgTH6up+F2CDaPnb3Tb5OPoV
isC6s+5Lf/vVw03dgbIRHa9labxoTYPDymSDk9v0tRQ/ysOCI5FSTjf0eVd51+/Pgqq0nY2j2rjx
eHGxWV9U2c8eoIm/umpGv/bJSW38SCCnn16Khco1EIIpdYniXwRqA1youWERvBzTkG+NpgCKIT67
luV3aYx20Tp5bVzQUxbF0SDRmOTgKvdjpofKX+ID8hpW/slDUVO34Y82ACD4zqBt+PW2zOSyngBA
sIUEt7n4ZrSjWPkRJcDuHkm3lD1hBSEdviWvKvf5cd/s5WV9q8kKQXuna6nzO3DidcPfMzr4mwr/
iDwqPOwcjY57vO7V0eDLK+AUfCmviQPk+jJF5wgBoYrLDRo+8OHyG2pnYxZ5aWxYyRxpFvWU4Hmb
1w2aNC1lSw9Zp9KsYQpNz4guqApEF/Gzn4KMq5H6EnsWkypaQMSN/ZMDoHAYAdqGRTLjMWEO2top
jgrP3L0+DVEqu5s3OlfElAJoj6nJ/BMpDd4lYDRK0X+2lwDtlGiXXMY+FbSarf8j4tP0uKcfJu1Z
TWVrlmiqjGJcOwsoFVupkGDp3oy6nfPVHot5HJvWQ871bBJxSJqT6t2YhvuPIbt1XiMtXs8RCOt2
laKs+2GwY+yPwljRdYotQJmQHUiko6fhHBhHNdiFVHRPKvG74buhwx672LtdNQwjz/ubfxMGpDy6
ULRxmiIzbiEHUMwSab9M3smpCw5gTpWPtSKKDfkA+ZGBJlBnIK685+TYwnme98+MyXbGrNl4is9R
jyYkiy9AK3+OcWlDSP/AGjvSWAQ0L711wUhYFlQ8cCXRnbG9GKm8if5hRfdA9ZBMqsb+wYJsDCES
EyZdpdNFSzClAH3bvRgnFSP2OEaewolpUqJlt+NsYWtK03u+azg3P5618WwGrfj3tKyQBMLXNlbq
BKW9FqGOgWCKJUCOAw4FWW41csxzw+rdRopqSy0duHc8km8ncKATqaLkU2q/QjKXVaWBVeLqR5IH
g9V8hBEUIQ64dTqWra0i0RwdmS5vsGmfvpqJL7sOIelRiOusQvqmwOZs5ZMvTW0moLKOX5FFrgmC
FOQsh0NbAGKK+ey9iBWKWWQRqd4+FvC+ozAp5Q5/HLnNoFskKvwm/BKX39gH0jTjuY/VEleiio4h
RRGVjsI2opGv4VJzm5spvfjr4UmJG2yDfwMI+XhiSZHSYNvtoQm2tUyM6pQgCs7dnkp7FwN5Mo/B
o4zZwhczuVpiqXZahONmHvonvIc0SfCmhzQ2dEuKUPwA3CPvOAP7IrmA+eRM8wvEpgwpIGnDihsB
cz5KJ5s4xQev4n5V6Wb6rgiF+0imWwRGbwpK7wtmcZP7lBRDheVD0ckLIXi0yapVT0UG80Waw2Kq
g/2T6J8kRtshz4gKoib2X268b1gcNbTnftvdW/i9pJ8PqoPw0MieRymNnDdt0gQ7S+FVyTG3i3lB
g52+yZNtg+evFeLrCBbi/vZsRGhXOA3XQ1Q7SK5yyoJV8F2ULfKpWPTqiURbz0CJoJ22zxvgAQRq
42vg2RaOcxFVB1xw3qAOXxA8d0j47/f6Ff8OoTgi5MnMRkTSL3v2xJ0KjYF/ujRnR5G+OtyO3UsK
e3JFgwqZTDEVuZjnHbPIL7XxigDSTSJ3N4Po23OzZEH3mj4HM/Gw8Uzc/WuYcCcOFlf3jmoEWnm4
aWoC1nvgxV0pF1cCEHh3JuoIOXWHGyRSL9OWk8QjtdvmHo3LYj/OsSp2vic2TcQqza8HPFPGBGPX
IjT31SNd988Pd164CyPyyPP0VZ5bbVC/FEI2i7S2v/uJ5BgaPquVl2qgcgIBqVWP0P4JC82I+n9k
FK7uIEVFuOAxd25o87GcBx4Xwn/KhP/Fx7xdVJJxLbvH4a2xf46ovlWW2Ay/ETPo3k+9+9ozBYiw
DP5lgoyTlmLizfxCALGekw+c4pYamPkU35zCbEz5c2wxUdjft4b2vQo4hNn8RWtKnvKUTISbmc5E
qTgioouBWAdm4jUbn4CJ3MTepQ5VbpZ4xX93nRcmNIlaRpomSN/YPm8/aKY+XrIK/GzAw24g0mof
J3pCK8SxnyVYI+dSugvl8/UlCx2qHy5hCOeujb88PFvFtWY0N2es5d7vcbrr/4GEnUyZJ3X1sCQf
qXye7MSsTbXNgYFEj3HoZtW1liphCeIqbohMeD8M8si3eeZVxnyKJFVFkWP/vCEtUg16ZhOm84FC
8s4O8Gf0sY88LMjGLopqGprbTbfulMgISdu5/jNJJKfMsrEOFJghXDAVi+jHmqOzKDPuefkzm0kJ
jWWWaImNFtFDLknpxYBqW/r0FkdcicrOxJDeKGRgQR4FB7BWi0Adnv+EwGUSA2eA08Q968B2uIzW
o3BuqhT+5ZmanJbTtapZR3h46trU0tpY0jtaTu0ijoFpcSz5ibiHx+SBoFdZX5zgb/a4NzsKDwam
Ld3hbtTE//KvZ3Z67j1ikfLtvEd30+6G15vlG1AKg6QTZu7La4+qFeoUgzg83xSPYltcjPCvP9+i
uSrgoim6VvZwkrJWB6WrneHkWzJB64RJhTay2pLxLAAHi+MgOn94IdJdgxKBG8EkFtRucWilWAJo
jd4f7YV86iFW4WqB7r6uD/Lbf0Q5Jq5O0m4gOv16n2ugo7lHO/QTWS/oKcgp+/nZjNFWa5Rz/6qN
lghGQKKFfHajw909muTur8pH+DLaJTr4GRY2Y9/gEzXxYVFly5whndD9dpSZpkAgqziNFhoBeoaP
5xOMArkYJa4D1gHdhe34OpXTBcfpAU7Z3jqQ7pfSZfbe4EH5pCtEgRpJvbqHSHg5SVgpyCa3gYBR
bhf375CbVLy6S2fyNUUTRxjyor2+opkkGzbdP8GYpMd7z8BFOExKOEffGkV0lsfv81Rm0rE8Y6XG
0VbGaD+6uYeaNqI5bUOkXhuO6FuI+R9G9tFI2zmVu3k98frAMwvXA16BVCdOy3ZHO3nvRfptzM1O
BSsoY5STOog0aL17E6pqJ2N+yQCawrF3l8Ps6X7QJpNQ2ghFVTeIZxy3dH63QsIg7hmZZwOvT8rD
yyA6eb+iDPrhiZwXvneW/azKkFLOiFV7KYR8pRFgsUDSO6fKVEaHeoAxCZBT4kfG4R2vUSvfcyXU
pXU+nrPs3eY11QG7+CSV4QHjjVlwznISPdSA+HHkotQBI0fxQuHnVOZKOJ2O916D9DiGQ77WgBLk
MXpGlZuIT76j/or+i4T42ZbAQfPRThNmQW7qgHP4QyXGBcd+map5ZKaDZ67WnrjtAKkDxYoq2wXK
fxpXmTjWtbnM/mgHoDK/S36mJAvwuq4Tb9FGxF+PEVC0Q859vRldy8dLnqtEkcPl5uMDPg+gW9ul
hWAn4AFQDd8WN4nOvbsGKueJpWziNUrxjNW+8owFdamoAeaUEKhHzYCszLu29mCZjyF6TpEVYPkz
VNzbAj5+eWtEtj4XrumgZvwm76+i2vPqlPDQ1mpAQnQEV0oOt9GS7LU9qfE6wY7ydNcaLJBFp9Tm
mx+ofzkfIL3mhQUOOd/Wtw+vfne0EyXRpGP2MtBR84ZELYzBs1lqzD3U9MEGmxiwHMvEHfkvYw8X
2EJ2CPFcDjhh98+0HijMWumpoU+5TbLNgTw7v9OvRMk4n0T1bdxSXRqGDuhQ1McVh/sG6a4kscUr
iTZgcZmThgFr4LjkEQv1i75OrnInAu6pjLtvtvy0I+z+ZlXkEmltN9+COAvMH8PS/msOCf2yU/jP
BgC3UFyfWl7QRixzGd/kfSQief8hPGwKFkX7wvaSiA8xW56MCZpJz6RE7dr9nupK6NuUyBB3M694
5O9jMF/+pTDI6M1Ipo/UmXVLgvUuoiHzYt7YFAeTUQJUvMilYdd1BNu0rquEZXbOtosgLKuW7obC
MgJMHtZz4yPeblcXRby7r4IUlxoL/9rm/D2AEq448IpU1BLt22CtznYYATq7fkxX/ZUYQe353Szk
5ZQ8mCfOxO1mH6gVFWA6YcdCtAH1O8BYtetJhLfcI1VrKnnjEZm9BybIGmY1Tsaa3rY2FHNVN1q/
pY99U1V/73mss3JgLCjsnnEWTc78KjDsQN9PSMNh1U2DMi4m7G/Jz2ZoUz0/o50eINUbyKYblq76
cmDwwQ0Oj+gSBILELwIIdR4949Bda3l81qSpL1heAIj9Ympfklx79utrin+GHXT624VHtEA4QY17
SMHKnhefo9JMj3JqClBYOgHHexuIO8zz42DONYsDWBDFuEoRtvmt5asSoT2XNu9Lezj/c7rDeXCx
0ZKx1aH5CH/Rp3YeoagfoQGRHafp+iHoASMu+p9g7Y584bnwKmaFtuYhR7t82IJ2VXGOYPr+rgbW
Q3l6Bqv8oKbdG+eT0kUexOdZl1eA5qjJDUSvtac68sQA2GyCdFe+UBtxxyjM9g2A45BoITGm49YS
rvMl48fMzwcoHpXksLDT9EQxucd2me8qHf50KbByAvGGpvr6f9R0Fy7OAXvYW2vHoSmFOBBxvrTX
h8fxp1WczvqEAclY100ILU7g7HF3yKxRl2ZvFOHezX3cg/xhHRIdD8a7gzeAUNMKLlrFuHH2Ncwy
OwIpQem7veqcoSlwU4SNl/PM0tOviTdgF5VRTEWFnSmg+T7zYGdT/ITm9UZahf7kvc051ZwkMBHh
qzVsw66FY4ozo1i891fDFOAHWBlq3MK+MyvO3apqvYZzSb9xcWrwojXEeZVScVuRkyN/aJIXDoZP
Kl5gDZF1QKyepN5+7c+SsGtNr6pv+SLKbmIDf2qLjrI3W89AQHuQ9dmTrtbkwmj7Pc8o90S0KW6+
SLUCG12/acjwDxh9D5Gw/8psz1/H4ikDdjtrOz85jwAKZ5nipHP5s9yUYb3+b+VyciB9AvoZN2am
ZnRv2eaNy/Rvh4YYWNQRWqadPJ2Bdvw+qTXc+hxuqVrYpot9tm8+WUoJtIqlU1D3rrz3tBHY1zyF
uLHWCjkMiih77fK/yQXzOia9sJ637sii0qj35TZKgDvJc9LB3838OBk6SgZHy4/eVzShovQAlQYD
iHb3xo77YAI5ByMjghYd7wrI1Xpk5/D+FGfVpxjMYwk1MPtPULtD5Re+r+qcjobtfz2aXbYQo5/P
eAWkJvizdWiGLEhtW3fzi5kkPYqVGJuDyg4H8kSpEKw+9OUivgc5b89EV2XfgPV4enpvD0DLSlbg
TcxczVZUWbZCdqnPi4POjBtH4RXfEyLO3/fIrx3ql5pfSw/BZN5M0tVsV0/kL2IuzMkeRu6bR+fI
Qx5UIPUem4c8Tu4ix3m4y5CXmrY/W8R/GG5BjcfFL0VSlAGOks345bRTvvJt2P9X1jXRwpSu4DNU
hWGj7MQD6X5rORQh1PiTI4vGkU5j62/bjXc4JwRF3UE7VVZvutCQ5LSKJw5hSHcTxzSu+Rs8EOIB
KpcIXqWgaYSoixWIFFgCfJtY6Ki2d1hwoRMpx6ovM6XOQlWjlKx/P6GbFvQJDjvFTHfwO0PGmXvx
+RO31hqI9QHyt+gdPzq30xW50HXmwjPOolFrlraUB21h0jhOtEYKCYDXap/rmHuURxwYB43O/+JQ
nlOVRgz3Wy515szWfeiHiPSoM+a0yu5dpQdE2QXVzixNk1yQPHd6SPouSJr58pR63JODN6lPdCIq
cMK9ty48t+kJodmjxx/SaQjj1tWHhvmMum49ixuqPgxz+AXyRXf0GRKmwT38Gts+azWNRRz9SrOv
v2u+qnULZbQZiJaod80E1ogcsZgQWGNItu0dvF6nuIMyJfaQuULFzAmtyeTALsmCI9kj8LWXb0qr
chaPidLrdt5LQ/PE78SP0gYcAm/JFAsUNBy8SjFmpwALCxQ8Aj7rCHdLe85c76ghVMpcb/yvYUUR
Fz2QP+s8/J+0Zzji3jTueGBCsfeA4rMT1B2vDzyyI3+ZJFvmfO8QHKfz/sPKH4obX8f1zP/786a4
FwfOf7M+HrizQY9U4UPsQ1RpU0zIhcxplmwcnGQYI2rgLmaBucD7KirMsR+E7fFJL2eK88GGoskQ
IcSU/c6aaG98SN2ujZMY9h6X9AIQz88qNskeemecA1MgBZerHp2Y5XKd8eNxE70BGHiWFrags44w
MK2czWFv8VURaqwPPGz0hTJSms9U4kWz/RIkO/CeKzIki3GqnI3eei+YS3mTTHaGM+pujSBSOZhw
+rSGWDxz9/7z+2layv5JyWgoD2fe25xNHQZUagg7sN8n33J6LMQMRV7p8k5a8PFCX9MD9BO7n0YJ
VxKEZTk8SyRdrSVXEQFfR4aVn7hkb9e+ZjpycE8lT8vcMRXBoO1eEMcdYiAE7WDd8khdtdZb7HRg
4ygxqPtcQuhrt9rNIHptFDy65/ydCnqanpobWV3/k+fy8/mr5iOzgeTqyXIo9eFKoDkKdKerY1XQ
4XbRohcDLeFZFDkGOowRw4x3gjyWZqKB58u8ZfTMbn4lAgST+KlAgfbHzwf4gJI+XYY+hE4ovcde
qrYIPnwm6gpRDackHmleNbw99wQuIDHyXzH3Y2sr7HYPFyYchkUTdKaQ/KXdi7B0qFXTpPrVRYdy
kgNx+qedPaz6wxSxl1mUw2CEaTo+rEqPuroQ7ylDdivKCDcqQI/kbAk/jJg6I+n0tRQy8GHckzSf
dQYc4gDRjyq/KKTgcXNnUyM56klPv38aCIT2OmjpFTFzm1WqwXBGBTdw4Rqty73nSUtWZcMjxH/e
edzJk0n1ufOYM1gQNTSxSZKUqpIw3SLKjmSGOc0dFy5lgwLI45J27nnCoRW1WRlbz/Qx9UY9tk4u
ty3txgMl8I6sYPiG3rCgoFIXXelHq7ME9H9mcKFbHg2A30dz6bajnqBaPKfWHsAMZ3yMGeMtVW0X
uO3u9Mm7ubFEuZk5x+ba0+MOqa18PuzMdmQTff4L4+WCwsezcniyG62LKkNBqVpNm+QXQ2GDCg1N
z0nCQrdY+b/yamnGB9wJrzUlPZFsIjnPNRlECqLxHHgGFVOIcTguYj1no5Hes5ShrBqBdi8GZBta
tBz3nJGrbWwGaI3U43LG35NsHlBM82oY0PctkpeTJvMx3sF9QQ2tzGHkfSP0yg2cUX0iUVaLG806
f+AY141IgErbNRktb9y4zLUWNZNkWTJpx58TYHLmljq8BnT8CPPY/Lxk+uzVgkyBbV5HtrqyPfNN
a1UcCnf3tdZhAyOZe7/QilXuwcgWkTp7IvQUoL/c3AOVvuD4dpr/UAEotbhQxxwuCe4w5h5WUiqo
7QDpYHKM1MzHSKGEB6d+HUUp1Y1Mt+p1nbXrb3rqALUPrI5rguNt+0JAfzFMkELhqeOj/8TBpLRD
end/9TL/TiP1DZzfPK9e51Q9KmIYBtkLDcIKAIHxpMTlWXL2aLCXarrKwwzjGyZMBMZ2Rk0hUF1u
W/c5lceP9RJhasYp+gsqw64heJWZWRtVIPIwWsHAbnt9b1mTU/ItZizFZf0KVt7NkluYq7ewgsNV
bll1fJDCsEI71uWhipQ/qRPt0ALwGo94MX5CaQP0dh8mxWa4VYhvCZArq6tgTsiv/NAH5puVsZ2U
D0idjxFBiOLxjDwUgHQ2uQbysqCWHDM6O+/GcihaFQcza97uh2/d7KGLNiA1n1Llm6gRaLgEKP5b
/8IZuYiQNfK1DjhfZft67UJvX8wSaFfqxr4sa5+zNB2QSMMAeBPGJV2PSWQwwe+5sFcEvD7K/oX6
gKzH5/RBa0SA0lNmwd7PfssztdxxYzFJun7CYNGROJpBQiPlWmKGHnXmINRFYApU1UlvViuGIWFZ
9xol42AXpgoFfHpbtZrbJ9x7SJWJBZMmezJ+tkOyC6qDJJkSavCS5qfIzT9DMnxKsfkZIsB0GlfJ
6KgcQbru1oQyjULTFaRrFaH8CDQiG/iLAsbyZobnEScsdHK820mT3qtHT7fB40g9Gk4BWNxu4B6O
3X5pyZ9/PE48VgD6J+F7eJWq8SyEmwUBZPR3xMrmWMbwgh+dNlMIv1Oie6MhMjgPtoaepJRmQiwm
hTwi/xZJXpovISM0CZoJYU4+OBdaEq9PAS3JWAt9dxuwij+MYqmSJBGTY7II0zNbZBXXkz7tZBMM
/K1s9SW9/DH+zdurAiurLitLnRNjB4eOn4KGHPzzMg82SRfR5wjknNzhP2ih8bDAqiUCaOPQbnZH
vqMZhurRFEnnaOochHcG2nXDViPK9PO4nXkyeJFUd33nLS2oGdU1DKbRwh/gCmHiXl4L1SO5J3mq
VE4B0HpKXtjCJJ//rDv/DIHUczTYDgxdMT9wtROzlRJR81VejdI+YSS8+vvqD1jvONPIWspU0nw3
w5WrAgkx/7jF615sWyqPNvv5dl3ZrfSvM5bzUnSrfcvzHvhWscHBy5MXbGeEfvqo3cQW+LD/9C1e
4JO9TkVuDsDScocfUrgLs/sWUbvUoBgxSmWvprOp1GlPyP51xBbfZ8rEY0IGUXvZOkDbOLIfTi6v
rzSUU5t0fp6U+KJJigEZeWKNEsSA9duu/6JyGjKqUhn/JDLtIsMCFTqi6AwCD6keNrI5ABqBU1ZX
vDSZpLp6S/jzPS+GbngVFI1Sf6Ff1HCY4qJsoW1rMYYJoRjkG80hIrNSKuqh6Cr7/ZoQfUqFAty8
Dp7F/FoqCFohFIPc1EoS+fia4iT05Li51fd0icnd85ddveXWQmY32KRTUt422qP6RDvNk6W3GOuv
XrwiVU0tlulCc6Mn/6LD7boc6/ZxFyaejGCiacZOF24bNFqobQtXm+wZ7ginh8s3JCltv0IKdqxD
8ZMR/HdP8EnZXZ72OmXLDlQl8lUIsGP/h0XkTj63lTIKte7jhaMX8A0ETHY60+xud6EVPbwubp+/
04WQJTF6anYblg7Va+L2vWY1NWqCmXy4v/+taYP8721ueMYZHp74JYt3vF7ot90yfYDPl1xiH9zn
/SQiJ2N8EBIjsqLKQp0z5fgRmIIQ76V8rmhZdCutE/lJKLcAX6b3Ct2VhsNqZiJqhkfCSAkX/BZ5
UANh8zTC1tDExxYIPZ4paQzy+FqJvpzoyHqYkELgGRDpTbMIOWjLPaQhftRxsWK4deQjFXJkXyqU
TPV0HI+r8r02x3QiaQm7QMOSvwpTYuhP1rnInGO0gsoCsje4BknRIcgyI9dww2NZ9kFE+pZKjIig
4eAIuijDxNBJ+wG9eNMBMuWZtvGaw3U39PCDa9lL5nh1rGlu8whuJNCmz7LLmapszMJKo0JQtXfq
Dv2t1HMI+OVHQAtFLsePzPwSdCrIzQeSnObfJREK7kEynH5LhSz+t2i2BBfSG+Fv0DKBlsMjigSD
bpWnFTQkfeM82+TGSruoB6AUxNoC5ruU7NRX9BIFKslWSAdYo4sBbaxzuRLsnQGEWMO18yndWzBR
3nFHyqbL/+dDcPesotOb1N2rM9g1trlJeprbdXYG9Vk/rNfPC94bgy5xR/NM0+LeCGHIJyGi7wIN
l6cyvCky+eG7vqw2dtokNL5HbUracs1okoqSqNZ8GxINVoDfzrxCPMO/zrdW2y0xfEWJl2CiKxpn
gkEBRACddzIaq9zpkYK5B3wj52sQr8PBWKXvriM8wTWF8jsJhMW1yxUuTb4lXWpYnEHrJ7cH9jpz
HlGx7zEhtUxqfJL511dl9SRyH3UgJKzMs7Q23LaCsoQlHR6k9ibvSOGIyJZhs9mc6W9FeRaMzGm5
6UJ9eyLNpB9HWIXBAUGW2xwU1ATQmLGgIedeTL5a//DEDgOUXWn9nRU+a4S36LHoRIAipCCY/JNu
tPH23QezzsDczJ4pdxxCw6IR9EgoFDu2Bisqu7u5iuYAlPjXYJYyl0rUckHaiGFP4ZiMhdXuIDQD
GPxvKYvFRM8LmWBBqtLQseP4xvNt+uJj8oRKLWT9s5718qe0QkwlJKfst32hImsaKK+Uap6chZZw
mV0sBACqVkHwtIHRMP5WOz2p1gn3YYTAb4hJF4H08QVCrLYsAzXrm3cd3m+kQKsL0cKc1/tdCQME
6r0pYCGLyT5Bl9JAYkTtpYq9TPMqVcXc6ZtFqsojIwnoFTHXl9mH1HsrB9DzFSkHf7XrjMPxjF0z
WvEFk9GHCQ4tld/M38GZxI1EqSE4D64aBJy8btEPumVgveZ5zwoklSvScrjyjnZy7Xz4LUJ0vbzd
7Fb64hHcRReegEjy1mG1GP6y3+ah/WWZI7dK/l7SVE5Ayk2pggvyOI8Hi6ve2tioYjjn1gyo0zrM
hJwuYrBrNuhmf5eoxazRmy/OqdFZuAYqnqRovcsnRe5QXB6E+C4+Ef/pvXvXnjf6bhdg1PTKsclc
cET7Qr8wTVw7QI43lD0t7rQTEzGw6O9uSb3cTR7OKAb+Tpg72ZZp1FqRLmg/OdivcB4G7nV7E3bu
q8E9gztsOuZB2I0rDQ5jnMrASH9VtCLHvFXafUYP1ky+9mVtv5RbWzHcEl0t8zhr1hhTknCPU79Z
qG3tsZNIGijcdHCvPPDCi9kTQrhOYgKsg7vgdVoYzECQbs6wwHODIGdlfHJnjd8Rr899pGmAaYFo
b8TYWbwlxfjQ/n/QcgRUh/8tfsACeW/k1g53kJhubPA1NtTUlWfaOQbXE9OxkRD4mf6rxxItYJLF
9zUOZeXdnbcrRuwPX876k/02sw0edMJP5Ix4XMKpMOcTx+dz//3llFoku20N26CN9d9FQQM46PQh
z3wiFwWa3V1K5ffgIL+7nfGaoVWS+p4Qh43rTZoBFEezT94zX+X2vHXbVsCAzJZZBy76oBUQ1N2L
bmO9zOZJGRrq3ulUkEV/S4+VaFIwpPySsabXHZpp3O3DpnE0N4+a02axlx9t0weFtAGjbGEbfhaO
47cTQjJtu6pSXtXpaEigEUK7042vPIkMt09LG9vCCTzQjhPk5vykgvFgYI8B+FaOZDIEj5fE2KVG
TFutWYkwRbWvFDiRkIhXpb7TzZhhDU4ObF867LNArO9pcQ2wc54gYtKTse3zbgKkmRz7SxA7c9qD
43UIuixFcGDuc5msJoNggSwdFvmuJw+dWM66hrJpt2EiNgMvkr3wipTLVn3A5+QL3ZsDCLQY9E9S
LMtHQI/87PEtFJYqRKKBfJyLglt8rxy/wJnMqBsVguZhdgraFte1j+DrR9xEYSSiJVuvZNV44Cev
hIZl4MzFDCRfM3ajsrDWS/FThKH6y0OCU/yFQqnIqB1scksYl7WVrBc6zQiVVoHzxEpwuMrE/LVK
PJ1/HLwxRln+glGN4Y7Ap+ql/aUyVZ1+AmfSwHFTCV7sZQ+JINI6Q5bZCiISrOkycGfuENCVdBWP
edSmI/YLGwQrqtr2YWvvKDFpGbFHCbHqus4mUeGVF8CVbsuS0rRaduYnPvyUDN1AKk2/gBLK4R4u
RtavnnXvOMxPjbagmwtBHoTFyjHcxrr6qDhAPVDH6YmopKIK4S2ma25kk87GG/eN7aVBcsZKLZhn
1CaZLwGPLFENeqSHnDQKcm/IMtYI82bqPC05yKpFUqBif5wv+4ycNCkt1qfImdKnQzSn8xXGp1OR
TzTAnrCG9ZfMcjuVQUA4LNU6oxReSucMe1fd+pwj0+GneyRLaKMM2a1wgpwroIuuOPX7xYJCUdE9
3xrgdchE9d+qoFCdsiNVbVBc3Lh+JCVuYPzYdB0DcuQ6kgkoZKhZ7oeI+7WrxuwRhMBvu1/VPzJj
8S/v2wmWiv8iphgDYxyAWMuhPFG//LGyP9OVhIQlPytfWo+2ojc9ls5PguJEd8/GoVei7ITn/Gf5
HPZrpswc1FfsNR7H2RnPYL1NOD71O0O6uVhW34x4fFy263rbnS+Wz7z7/HsctRME/9twu8arIkMe
WgcwS75zWCrKpUaIs5GV6GzPG0MY2U57bG+0aAA0VuaR63/WpturzYrEzGcjjmt0pvKj2BpaSsGH
XvcdtRcHPQz+9oMsXgoAjsPcDGkKbIuo/q4nq5QR1pPtp4SpNxrrxIScEQHKFffeBz5GC1Y+VFde
ufGwG7CXlV8/xl8wAIytGLgSDFdmaAngCsxONEeRJXyyRBUU0gu7vnetisUCliWLvmm9QCt1P9ne
lvRJLgglsQOcNuc9lCH7z4vH/4ycto/JlO/dF6THEQCUB6madrRwUyFSuFu4ZtBA82ra8NsJvXPr
BRYQV/DIaXRVrVzyPlQLz6QCzB08Nd3VyZlYmwyJxJO1z66LLvS6RPVEPD23t2SfdF/ZfXgv730p
V1cnVfVaBPfjQ7cJz5u21TYCbIY28N6Lp9huTGt9JLp33rw38a9nAfUDo2VP/AM0tOiHIkPJgilm
DGn/toxCyTMnxhYV8NxNX8P31kILaXuVy0+r0x1PDXIcvRdwQ2FUmNDRIiarn5+UgMWlqXHWa27V
WdokpnnCFjUePAndD640CZZCGTlFX/1/mEfjCxeiTZOCtjDMRETbn+4YBB4nMybRxgxZ7nQ09VWO
UWwMhS/QI7p/ZS7CirtIIO02jyYm208OWcvth9SlMc16dhq47prrbMc1TXZBLOunKsb3KBFlrbjc
RjPH2MJEprTWVEGzG8mDPStoR6X2VecmpbJk7AUYI4A3UesxJqVAqExpnzjzYgnYnJQwh590rX6T
TJWhmatr9xjgkNlVQHRaOOXmqCYEXQxxZ/oSOf6j+eKku7vzmxVq4PXK1G2Gpziqa+UJCBoO9IuD
zn+cdi6xFzfP67PX5g13u+dJapZTAaKpq3DTOlxOVtQrquk9dkggIDNzLG3PtVzqHqSJWraSeDps
9B8JoYkgu+DQHMVeB9/XC0ys/LWKmBdWQ0Gg23Cp5HLjx5CZ2Dsix9Rp1FbJiMKUR1UsqIMK7aJu
9351Ue1VrF1FEeKet/9N5d6qDp/F8XsoCOKSShHWnBBRNjWuN4Nkt3BuO8Ozrsj0m/4GrNBQBtaQ
UmVx+k15G9Qja/W3ta/XDkpFx/5WGZUV5JIJdMqYF6sYusERVqK9gQqHGpGB3feWBBxiX9KC7NV6
hD/mpYMnUfTH6DXVKm+3Gzt2UKoE4LGvddseF8Y2pdYfHu5/An/nY0aVKFYkZXTkl8w+/pfgtKwO
AalWHJ195zcvtCTsutdWDjUUWptOoEn6NY29eJq8DiCXvwWTqT7p19YnHCx6nXDpfcLlq3em/Pgp
K/xVgnUzof4ebE9rSOxnK9OMBfwKg00srJ8nTS6rNbd+lEdNKR3eBoFsKjdRWqSLarvWu34L4eWZ
VFrAHRqmT7bxGLASaZt7rVIPvIN0d0eBe2ZcAZs8fWTCD9EiUO5guUir6Xm9fXFBaURFEEet1kXe
pVmDYuQlotGoRoPpklGXwdzBwoYNgR+qcf8SMp+5Va9k/VV/OwxGPxRwbrhwzuI36i3jUsFhMKRM
0S080gifzHyElAW2vA7INP4BtHuZ19GPMrEkKMgKN4NZNugHXm2ZTIbUXS5Wm80HusWwD2Ned3AD
9wxBeKnMhCTOE891RZ1HRqePMhkenvcUhMY6UYM0QmgbIbZLBzQj3JrSUULSY4OhEjnzbBLm1YhQ
jF6suZDuyaZkofRiKcHcjuZER2UuZYiqHGKnlTyZ0yVGHyEnFlAfFrVMMlZ1l7DhWiYU48CSYI3E
rM7dHywT/ynenYyhicxFM2ItoCI+TBBVWsGcpDdGXVgcUhxVecrnqgsjCI9WG4VHy7Xue69zKeE1
z2pMPX5YTIjZcymtIQnQ6PBhJ9qtTZD7fquaauG3e2nFwE/0wGkjpMzLeBaO5CCCLDy9ow4jvBK/
8RiwghKckw2aTVyxB/yqKJ8d0HLeQ63YgrCwZiPXvwreUngP9e7Fpg9Z4HHDEleTDHNWNRCL4v4x
V2T60oUwfOk27VzVbLsucgcQthlGmCZWsGHP3OyvRyjS6hf/d/1/OK/JYjYZybMBxslPQdUyWZBv
g5pOf9BA6N7HAIHzSiLKz76bSFhbcGfxpwVIf7QUlj9cJ+K4+AmW5uivYlrqKEP1QVRJ1ifzxITu
J23/ZFhMHhFS+K/sdECHH0ktnReqKKRj3t8xxG790yfBfF68mK1g5aGNT8QlV+p17r3BehxPQZPN
9TMen8GB6ro1MWag6r16jZiwtE17X34dkwIIp2HGtxCTrh5R0CHActkfSiAJQUkiXUBh8BRGCQPa
SkyDlerKXfxQUxSUTHo8yFmdo9QeSNdqZTRmt5KNWOJFRM5Mz9WGwWqPzPfQvZffc0QUA2UBCBMw
4t83ttQ1Jvoa0zZuB2aPT5sLrlf8Z0JOe6EWFno+wh5jdynrnX+RmRPEsxJ0/TIzZXplNgzFNZQh
PZjyocnHuPmmyL5JYuAeTEmWex/VldEYqjjCh80A5JPsX2h9/qocyMXnuQHJUXR1RMIOlKa7mJSH
J+p97EAZmZmMbeq8cjusLbw2hUgVNN/VdYCOg3WYz8RDUszXYe27D/UG+Mh05UaqfWmhm2c8YtXr
pfkn4cAyzKuYZUApOq26jBqfC/PNSqRm7rXz37xJ792kQJWcZSlAV7sWBs69c9ReGafYXHUBT4Ox
bw0TLLhPFy0Mv4LaxBHl9t0A6Bn0dVen0879Cnbd2rK7foauVKbg2xvbqVRZIdOfxagt1xPmllYc
L6GEs7vydFMuYSeHnVb3T1x928fknlGOx8j87uciIEY/8XOgDH4EQFy3RYOA3Aae/lrY9KjfW6H6
GWJ0LJ3X7peEVOl6WwJbxAKL7f5WEzztamVwovJyiJEkgDL/U0Xa7SQL/KivNKEGTuGZ/qamhl86
8dFv2SvjdWtXwMkoic8afjSAB4USaVe3OmLNyzbnV359RRdsrznt+6JqS6//LUcAoDPDcgyYMqPt
i229q6lG0PmapFjqvAOxXdCSUpVqbyLVuKS7ofakYk8lrTILXbV5yfx5O+vhKOLI1Suu1H+VupU9
OT0Uie5kp6LYuQKdLfzSqi3Sa1Gp7C2oB4h/cJIRnwGmHKOYGxPViOigGgSV1dFgijSL39XYBRnV
hV5AGwrsgY2xjOkGP2Uyu6FIV5NXlGvIgGspPKS9VPH3JZ8DoPoc2g07LUhW3kGe2JgfYYmf9m+y
mmTrmNywbyyt19sEPsOMMn1+Ew1g+p2WOStIEM+q8OI6AvFyQJl1/UKjMwKX3abrauOlOyq/mdvt
+21HYcbB8TBcRu9hVls14B5Sr1z0/C4SCOug2uH2m0vFOanQ2wUvwGrAP2RI3x0Sl8p0WqJMk5WW
j/wtYOa5s0+gSZ3KZmWqrctrW6CRv0kOOkN5vKhGoYOwgdkQZCfUrUscXNtETL11qnt9wP95cTIA
LFb2Iv3V6B8JGFczhqptMTT8uj9BkKcTmio+hcP7TTqthPHHiDuul7qS1UINHALCVMmMEuiVIZzu
P1BSVnFadxTQ4mdA6OFil9fH/7kiTGijDEl5iMWOmaGEpfEqhrb+umwN4xChZSWKzoz8jrnrFm8O
Dt7nUZEWLQh3MdFIYQ9Q3XT7d5fmLImpn+0BH6QEo2W8GUQ18VFwWIxiDX0+9ntZ6CpRLkMDva9O
7MjOentiCg4XdmkawvD111/OXMuXs3BBmkV0dvkCQDc+ch1p1Az5kkWxQ5MhI25ClJQriGF6UQV5
N7Hx08aehMZkqoQDNLDKMPi32FbmyF0fgWHyfiViHbnhh+ICbpqM5FDlDwl8thOdyMeoz+phlPT2
uyTij5mn5Xxo7TfSZu4ESB6aZt0w8a7zqQxz3pHICzfmPULR8W8YVqT5DGUaNbh78swF1LZ+eZzu
kT5+tkePrIA2BdwF2ZbufrU1Gl8nVW/7F8rf4rTRNgrhH2KYevF922jffDXZASsBbS5UAiq/+WJF
NIOsRMWkt6zBF4X89vEuPKv/s5M76jffV0+fEncFizrVjjuTNc0E9YKDGblFwMBfAj7X+BvR12on
2Zjx2MFabwb+ajIT3a/l9vGaBuaDLlFdmiyhliYwiIUuWKFNYQzQa8vC6n+2bEqy01bfBi0HdE2E
YNdoJWufuGi0OoHge6A+v3W6HLpqDw5hh4Rh3av5rXU0zH5xhb9Di8ab0MMMINA/BgloMtTLbmoA
tEOi6OkvsGievyfW9BGSyc9HBjAS2fTpmphfrBtCfwsEXjMJpqe2XipySsGF3k/uiPel6gujOiLA
oh/S9RCNmqz2TAMRTn/G3yX9KUJItJEd+CsJn5RkG6q81O4eTDDqopCRa3w2nWFv7by69TCN9Ko4
Vq0zDVVGDCpfR228XzbdJnyxUrdZ1N5jjuoF+HXZX2NEe+ROOBsIjJFCdrkLQAlnMa0atqTaG8II
dWnfQQhc7sMoiri2y66MVzzDeNTctStx1exomhXjtSs8d9yItfqrDmxaX9qeUnicTsvLDkwnviIg
YL5vNq9l0cfadcimqnBfvLPTDYxhHXt+9NQXPG/Xi1wTbStApEtsJ71NPSKXjoaX2JCAwY2PBOg9
2rrMbCgVpsuCmVDMEY/r5CDcZodxDM4T7p4r4M5UoX+Qd4tw63LbsJEdVeE449qMj1w812QSHbUX
hPmb5AoweGOH3kt9zCSWilpmAAbg3n99QXUSBHLJWyXv3FoIzp/TIqPJPz28Lsy3ZCtVZnuWoEFY
OVyL1a1Egbo+VyE/ValwdXIRuZ9L3e6/dlxp2XH6wjilUr8R6Oy58UgfsmgXxdE2G0+ZH6iEUNRA
k6W/qzc5LlNr5BsYuA0rIc1gDg2JvGZqaqk+8RokRB9YCzOp6VWyu8LHNhbTWG80QQsid7iPAgJG
J28BuC5lAVZHt5h+tLo1TKHEwHrGH6hLEgz8Yo6TQVfB7UNfG8PlQTYVtyq2g1jjxFfo+JS2yBRK
hTaKfPy82BiMxwblALFxOGvC2K62JGswY7D4ZmGKisQeK1M2/Otyq1eIIzmlnIezcn4r4abJoVq5
3GNmVMFjLAjUYnKH0cjYRWxsFJxpxTYYcy1HpA16mtec8FyvATWUIppCimQjgPpOQJYy2cFngqqE
k1gtswKoKPElK6ngAIK4AAmFRcZt+d2GTYxBOvXnhP0SCfj1rii9S4MOml00dv/i27s0jzqUbGwR
+lO2zpIHbEDZgPPEjn7CyfcaxcUC+tvaFuQEXWmTZzgpH7Uh270rSsLK+Jw7Ru/ninLfcm64nx2Z
nQO9VbMplL1Tp75P+OasJGmF7HRoUcxoSjFIeygYWHrsnSaYjg/4IoPk215XR4NM9X3yKHT8hFi1
xmGIzL7FNZt0VbbGRZek26i82rpReWGL5b9B5q+gL8hpD553fwbVgEKIEGSzC9b6jTvFVJjjXqvo
G3KSjPUBDyfw0K0W5qzK+NOtttldRpTlP8oDIUPG1lM5TmTG12vngkNOovLixwPk4gTWrnaerS3d
IbNrYiT1EHGo0NUrydJ4+GgEATeDIFilgRJkzGq8lIUscKEOGyIPMPYsDBWeoSxT0IBkhOv8NUiL
j5Gz3q4IRCMgSvOLS0tDLiI7+TzTSeDEc/jKhgXxPaT59qmhukkeZXURWwB3g3Sop/yKOmQoqFEg
yNsplW31bNkdNOYFPhqYFV2Evq6oY09VIhybVpCQ2/AdnSbd6gQpAbzzGD8vgr25C+jD3N7TUZQL
wz0tClRjnt8JC35zr9KCRM9GHwMrXVWSeM8Mk88wn2WEZh8kBRSq9+lE8D+KRIYa/PCiW8WVRlhR
aWCBIYsXinFTnub0CYq+InwCZ4zzFKW0EsVDRD9ptffm9HG0X7kfhg4SZ1h6b/iVQa42XZzauEZW
8pLafWkEcj+LU44gAsu98/TmXwGUnmh+cFN9K1DMMi7yHGvqGQlfDOnc01XAu3phfA7NDp51LwrV
Dp1VnVnQ5lWvhVtxdBPLwZcRukVz+O2p9eQ3O9dSY3R7586pLPFq5oE+AHFyBS1zXDA42hJ42UTH
mj8DGmcHnZpStPZ3Fsh8JnWZusjz0ZTGX0XL9V3pL+Yu8jNazVSc2PkIaxznoL8oVDfnN++n6xgF
c/AtV6vJzZ/ebdY3RNC+C1de39IEZbeZim/PB8oMFLlFLR9k0lCd9CmOMM17Lb0fZ/Ni8YqCI/zB
nx6O72XwuB7m24JVR0LYyBWx7jkZZHHO2MqSiCw8G8HQXN/831ng5aLwWXS335pi/8th/mvOOovz
GBDYWO1jdmh6NhFWYy8coCbZTLIgzQPZ5vXPAIwaHw0ZETgczlo7XLJF8yq0JLJBUMVkUZ5wiYkm
UJtDpAzvUrfV/S+4y6WeaTPY+0y5W7GVfdNstzEA1k9+nKYWjy34CVYchRNqPwYmxhTfHrkPsziX
ZLK4TvFlkRyLYZa7TIyMB3IDUdpmCfO/GY1bmwUJbvVdLPJotL9j0TKR1Cjw1M/J+pRurbAxS5R0
9qFA/QvjnvnqVUpDbsdT/mnwwcewN5/tzvjzAhchOk24mFvaN4Zp9qdjWds/5LJ3JFrNg92+aSXH
eokRuNJm25BOHiC0QnqsLy1CALLHr73eHgzKDUv4OuagT3enlcYxnhtTJ4Dqx3ndogT2P2LUZ05u
4Hyc96IGvdSizu4/h4FuA555qM5s9S5n9fa7kKYhkdnatmkZdS/KBypE5JnCL3M0PJzkOsPDi2sg
SjDj2xVANNW1tCHg1twi1GYHgx8pEbfDWmtgGceC5c4eTzia5rchBI93SEbYXCB/Ya9eFbVYcCWX
jtGEx1aOC8YMHe/3ym8l4cjl//sZxSs9kcjPf59bJBR0BKbck075l8auftTuYNJYgc4fiBtxGWRd
2MLgV2gT9gI4MmXUp6olqtzDAU8jqkKrjV5SEvZnozLNrimOSRI6MiWqprDSMDuuQiSm31WPXyuq
HBcKscpWSDz71ZU1WluDNoynRK5b/+707j1ubtyQvHGfWgvl7vOTtOqeqDjVjqXaqw76CpANWHBx
SwZ1Wrs4+x3zWLsZxndW+ysJYDY4h9A0eUpxiw3ipBfwsvOZK9hGbAtTpbQPmjj37rD4Sad3tRxu
WiS2FfEgp+nmgmdnTs06tKnTyKQwY9ZOGwgjuOnxSKAWEOky1Fv+zE1cPlLI8KLptYfHOQgjsyk4
TVEob+UbtTvxq4iPr6xjWrlnoqiBgg08DNumNL8ynxCA/5ToliKsN76rtNZ8PSbcWPx9webd4p8T
0s4ySgHTgaCZaeT/O164tm9GUTY85++KcpWyN3ywv0meQ59ctlVx30W2Nz3rujvSokOHVLL1sHZA
hd7LkU/Yi1MD/296Jeaw0WDyLlz8rLFi4F1CCxrf2wXw+tJLos7E7wm7XGSPTdtQtVRlFY9ElgpP
LqDjyirUlVqoDEPVEcYayKAI1+bb/vp4/wgdZ2HSPqZcWxw0R/51q7AKv7vNDHT1iG3s10YQQxAX
PmKBhakfs+iGpIkN0HVrd3rePQmkf5oBvbsorLmChMVIO0iyO5nv0LL2SGe35wvAj20kV1FvBgA5
Ith5rwAG0FwqSD/Gml1cGnO3X8r7IPwq5mJPkvrPStLBLjXAJUjGWWb0hbwyvTmLuy6HXXjYCid4
87HEL+UJ2yjmdQIwtvuPz1MXusCM3CbKYmQ/7mUS2Y3ELLEcs6IojTkE4IPKRhUpgkMZz88PkQxz
4adWe8ork6Cm5zqdfJB359jbEwSvD0s+0aJCT3M8Bllc30x1A3xWXsI5AzatsGqwjyMA4GbpH6Lf
9LjZU0bSkqMas9Q4i6d85LzEjzRWtiehw7D6iWHf161XDn/OfhIfHyjSDLdRwcO0uszEeSqGYei2
M8esOmPIlGwENSwUGz7CYKkiCNdDwNryapv0JK6M6jxR6OE5rp51ml7SsTs1Zd4HWci4EayaBFui
xKDYkAbIlHLiLWC92EhfTevlYRnp/rVIYcMt/iiAN98PXHB4npIWOgC26GfKQxXDBFE350ejrE9W
T9CzO1H3qCEEF7fVQzmfUwMCSNpunL9453GNrc2WxPxmk50leIE8fDTrqey3jsRsQiBcNW7JBbGz
3u3/GTbcODpsLYCRS3mA7sSkTT+j7I9/0zPsf8fPfJEg5y6ifOy8VtnpfcPOjz6dfAvBX+p0fOAg
/1C10JgqTjTEVdeJPLiCtNEHFT4FLUbiYWTFqT51cogf5QXIqfTiZU9ubYMBC1a3pZ8oIiDGFx9X
4mCYPLRxSjqtSWfzz5xmfZJXsX5wb11TWRECyvd6Fj9zw0gGLWyLvXY9SLqYnWuBN9eW4FRu3/En
5/Olx6wlG4RfElgdtZqqXV0Zo/YvSW99Fryf/Uj2WmSu47ckdAxRrRavvD8zWTtLBu76sloOfbSZ
yCxVesTsrbSDJnKQIsk1A+VTnUe/M2dbmpgC3p8/h+ubbqlTuyy6xUkf7kSQk7g/CXVH3odbwsjm
q2PFMjUsd26t3083sEFs/QBexQZEJ73N7TLXjJpaNe0o7tWMmLBz9wGr/3Fm5gOsR9evGlnMprD5
LGL3ycVvG/rYgy/BHnQ1MNMBsHb5uJjPhye8RoguHV1lR+uQs4cEwUbQp0WvaBQzKk8xM6LGQIRI
xJ7/L2P4JgrajSBz47rbBpgOtlwZ8deC9KarntChdnZQXo/Zmu5F8s8+ApLXOru3Y3iDkZ/M0Hgl
+SnDl90L8nAIDNKRbM2Os/otRgJI8dpOKZAQeloF/qm98UshWFJKgW/+tQDFHxS+mnzvUPWl0xUT
GhyliC1lmHsbU31fMYP8kSuVdfAeWnpHc+MOWCs0QAx4oJdFo+tIs46DwHuiBFZKRPObG/VTz9yj
8R6wNF0aTgcQzDxwYz969mQxZdZNNbPPjPiKg569zERpUeHvxzIzHtKb1cvhInHoqRX7am76gntB
6iJ05DCQvtbQbMbKX6j5wDSGR0WWvL9oLkvzZxYCk8C0kXYUZlQoqSCaK+Q3lzrZ4+tBIa7h2Jhx
SNS9ZD1ZJBeVVWflo4vpl7gfjfL2f1vl/34kDWFJZyKHOZCSRTnLT7Pc4TcKuhO47P4bdiwKq/xD
SrNkTQbd4mej2avN1d2p0wPzRkps6xqloC8bkqSBGdAp2wIdq+6dLsU7VPHIpJDTEhKbniHZBD0h
LkHJgIzfP6GGHXoYo4KtyUSDkcWZ8BN/LIxTyNJ8hpB1EGzVrvQ7y5PVX0uF6lqe2BZncibfo2hH
7O71m+Mcn05Ro4LgC32qXYKyIWrdBHkLfEKpEqXYVGO+mkgmamWq5E1jnAr304YJqlOYOHdI8e42
wrdHzDtzQRzld15z8wVN3DkP2tMqOjIfvvcS6lElZ/cahf+q7wgwtdkEA42iOPm/pe+XtQoK8ddv
/rDXxKGfFUWgcBopUAXnujkVQOqdUg/Ppf8yqcJ0KE+HHsAH7rZaBlR2EDlgB68Ss+mTs7Fa5iEk
myQUrikH0xLMUYWj1Vi4CN0KXAUZGt3tSvg9xGBL5sbZB579RdPbVr2hzf/E4apuQnTqRz8/83Yn
uytE8ZDnNRUVZnuKaG4/Qb6PzV7mvTsxefdd8ejQmQfhp9bf0JrmJ7aTrvrtFsVo2ZGi+hxv9tNX
KR7jQjvXLXJhi9jKcB+obtCEfU9bTRF09gY38IW9/ivYsYATCh+LRpnl3guR0uDPTnTDFsWOAonV
8Pnwckhnx3PClcYSvhf3pD24zTkjbbI3vh9FcdArwR21XyIhawjyKt0r+DB1yGjG6VLD42J/CuWt
WabLh8gOgGxGpq0EEasDsGHOeEirdgut6o0sB6m34cqxhpfdmvWYpp3qRlla1MFQRGMldg3gJQcf
nexjMDglXxp7oxtAgNtrTULgSVdGzp5rmCZr+wGC3B1bv9cURBokOUYVLLaZgB49+g2KzPzR5//6
E9D3UXFztoksYn1jb5ct+jB8HPJloRSpgL0PIQvtisHElHibIrj0L4dVnyOfU5uvzbTgaINY9kSJ
cDGiFVfujDAvWaXHyDkN7gbdTlbj0NnvWiXWWsr7Vl28HGQFcaHOvKgflAo0Rd7qdVTNCgNu6g8b
rLYTwxZi731UMPnDwZHvNEpyj3dJLrVicvI5eryoChjo3vjBLGwC2iuNr0qpHLmxEM9l8xBEVIYq
kYgGq0bvUYTdBp98c4zCKf3F/5wP0q+PnQUKkJMCuXQHTsswSyhVf5IYPzE1p3Yb7MyFCupiLC8f
5sMoSOlVd1T3lGHQl+A/oGFVjF6KJ1oK2cxwc11POYAODS3VsokAMS+TEsE0XdDgm4BsNtzf0E3O
pz2PqzVIYl8NBGwc7UCO1mmcvHpmI9H+6OblDG9OTiC9Enarwoo3O0zHCZmzG7/bYlblmdJBi2o7
56ykShlQrAWF4bd4mAbMrk1oJ9PAUdHMoJha4MbgHeSSVPnuhXGDAML5NcmUgVq5Bk1kws6nmK2m
JZJqnVsql8Wc4bQ0HlIy/Dg6eR0OMSqxxkF6aNZnXgosGzwiDvpbzJL8bqNrMK2Pkb8+dwFdPdMm
Wpy27cxDJOhiaWTMffmoZY3vBNgOxvc92QChOoUX2Q61D0wb0vW3O9SFEECguQZ8eizpOOnmk/lU
6DAXKg6n0f3rWsNrI+PNquSnw+iC9tSORN5IsYxMS8HCg2zp17kEpP3vi9ipjMhozKjNb4WYhfpX
O6OkZSe5FvA1tXwHGuShJt1dCSY0s8sdYIj96apxc/deMxdu/u2UzF4FIwTSgM4UWifOcyqI3HTN
UgTN7KKTCMQgyfAP0VA06v2Hb79kqofyLJofcjxsr5Wdj/UfmU6ljQkgcHvkEnB1AME3emUrPO8z
u/uuIhIV75ua1I/teh3UBAbFXPNKQ2S3a5nBVYUvPyQD5dGAWE1spD6vNJ5if3+qZep+1IE67yy+
2ollw4Arc2vj1blAZo/pv+j8kzcHB8NxZCvD5HbfJdK+TixruvQEB/7FiEuqgY5/OsMKkSrqAh8j
rnFobr18oDQPS0x0AQls0rbEBEVt40+1IWtPgf1vedwNiSwvQic6Zx3DqCQtC/4ctQlBZHRWTuJi
GRAcJBahvHIeMxu5CHGradM5kZuOrnFnMYDFVPVbLSMDrX9mj5WacR2xBFFDv64bYT+kxiqeop/E
bhjJ02BY5y5jaXscJ7mgelq6ziF/I76ayBNPEneXRRzeF6yaVAgDw9YkHs3WJudcCbWgeRTzxMBu
G781tQ2AFPQQwhybytbY4Q8XgBUaiSiXB+ooDy7Y5Q3pH934B6K1M7KA/NnY6nAkjwSWXUSxImKz
+jJba/dF650ALXy/wSbirxvX4ul3y2WJCDDjsCr98iUd7NkZpsvBA0zC3PyeNUNr/uNQrf6s4rfD
oyf3KeGLPLzqKiB5uAvB+ZXhO+qi2HaBHf0VlrIFl7zfK0W09m1toz4lIj+XuGfKYL9UTnGLPLyF
elOsJIe1e+HhpjFm8dw8+QckjjFah8bWqsM+O50gfkSDduwgiu+f14KT3ukmKeJy4jFxcK7wE2/n
pkJSlNMVRpQ3btJbmTYFbWhUBnrhz1ScT6UVRFJO1AHFfbmSDqLt2OJMdAuF91FvcOk7XVJhKcBj
YecklSRBNSTZo902ccFKRpLCert6oWqedBlu60Vf6kf9Kh+S1dk51xXX//JiDX5llm43LfpkfdM+
T/tzzqdV5N2pMwsPaDkRjb4ktq1qq2woIzyfH98yMGOM6w7wTmQM2CVBL7iz7LCRQKGdVvgMDFjx
DrffdfPGlVdL++B4VOmiOz6PrBsB3GjnYXpcQaeAsa0rxmt/NlCe5Cy3YpEhX3jsiNrKjxW5e8uI
9pR7estp30+yw3jjWmmVGAoxCgeoNoxWcD/adal49hPhThDt2inF2de82ToB2HLOrc6xA9KTg4eC
6ayT2Shs0GsW9W1K5bpRKic9zXpddJIqxwZCY3MQorG7EURfn6p99KEH4yHtVNrWX+eFq8FIYpRB
wXcdEYaWHWge0cz94pe+K1adSE5ogP0j27WdFsLQQrwDE+TpwFrWEqAt/z4UdDp/meBVLjxW6iBC
WImNq1ks2OyCK/Akb6YWsh2D2/LcqJFAx7SVFrH2drH2kGyy0Vpa+0e166YAeNNRJx0h/LhBPLDK
RJnCcZpIy8ed1inuN9v+KL/6jqrY7lrm8o+q2Y0AuGnV/b8c5/2QYE12EpTe9Ibph5vgPKfPMnLS
sOq7ICsZl7kTtDtknWLuMuyIeD+UeM+8mcD8E854l/AtyRt7zINzPMKryLeTpmRKlB7fs3bAIZCI
ADHmxOB8MsQSGmVPaWo8ntIeGesxJ5zxCd0YZlIq35B1Lj/Czewf4y5yXYys7gJJcunTnYi3Q4QC
0ci7BizacsUpxw3CzV969sxXtuYndZTdWnia5eFi28/uUeelAdEorBLt4Y/5cd4i0dtdml1kDEJ1
mAqs3DbcZus1KbDtQnAWHO/hYL/MJV+/13ru3kT8v+ZHvL2TRRHkVLn8c1W/Ooa1sQXFiDmUAN9Z
/pJp2JJ53uri8huyulPSs4QO3jUswQCWZUm7pdIPjpnJphWMr3iIIggWtR6VA/E5UgMLYCg0lqE5
GM0lYKwuzFth6X5wwHtx6dhFQ9DvZFI5HPscS/QejRrLCnMWRz5kJeuB8weeD+KPkOKSic0UpHc1
5lYnzJNDCc50yv/s/vnjSVka9L+yEXUuMrH+safhIUtq3md3y3tcujz6mvBDONa+ekMDDKCUByhS
Na4WdBp5HqNLqrf1WitGGC2VdfopvwTr7o35UtN17/upWLHtAdNxgXQ6fM6mGyoiXNoH2o1fgX09
K9zE1LiMe5uBLMT1OPED4oYg0U+qvGJdCmMzeYJHVYpDQhnLc7zA39lqUTc8hO5EvJd8Y67a/0ws
HatM9/Kaqa1Kshfy8YMq4MBU1INRRRN6QCKBqglZjNLWm2V9yy/rMEr6lyBcosNm7j6oV67emnly
Q1DexGS0euYosmFaSYEOXKh1DIolaTO2gxALgh1KsxrUhGzqIoXQZ+sFpRyDXIZUoUwa+8LEUsqX
euFoPFpgoAWYsCmeIpMYsmsdT3KIm4zLh2gD2GLkSiVaBkWl011bjy1Krf0tOm+0b1CEUBTBU0wH
P32Xs4a6BPgkiJpjsesmFOG9Qlt0UFfdwEt4mKK8BRyf6I+0Z0iVAZ9NN6/gz4lRM7LUVfMZze9r
JvyrPzXApuygzmzdaRozF6Ce+aIpVOmg9JWEQE/0OGlX3hDaSHwuiiUh06Wa/4boHy46CuQnJGTS
b2W+TziiLo1+aOG1C8848qFPklavBtkGfQiXxJIKb5AYHfH9TU/Gl1SJOaZm6bbgcnN75LAF1ecU
PiGUNLjScTj7W+WL2CNDR362bfqrspSNUAWNHhIRjzXCfs56MQJ2MXJ9mxnM5JgeUUgppVnKnXE/
tfPzZ4J+f7u6iV4vE2vAeSpLf+7vYDNDR8rxzvZpZUqFz2e5UaLqosu1gVyYXAXL9L7MuymjEjMm
TliF25qTkM07NVJT4ldZ1+sqn1hJO8CgAld8bZzr8YV6auE9crXd4M5WdklZTCvRjnYYpFlFvA97
JN72HBOKit73Gcs/AXzWSIAm1qJ7UClO3jqkfusi8g7+PGip5GKn6xUVP9eVnSXdFqiSCReN2Mey
XQM4oEt+fBGXy9kaWD9YLzJAWvJAjj0Bgi1IQZEu+As9remCQjS0TlpLx2XGM0hVmMoY4e4Oxbvi
JFgYmyzSSv9n6EkaMpzEynQS9mrjvzRBVm3ZxFonvVzkAHWLdHMJI3eA+lvCsgzAv/d10QYU/Lfs
5yYOExi78S9FXa19p+htFT5BfH1fNkJRESWIvvWkGqXkldqGTIKc/p7ylL6ufO79khz1rCDXNl0G
c9AkuuG4V7PJCO5DO+m5vdcVcAnxhu8oLXcaqJOt3AnayorASOD8Jh9D6/sDqO88X5SlRyC8SHqR
1ZgHAMJNdDsWFSC+v4F+me/QivUtJgw6DDsyqdGstW1LO3qmMJVF+0SBeE/F/Yqr+NIZCnCGLKdg
Lof5OnNtV/v8wpDpoiVsRclsYo0s4BkK/fnDH+/xnB6MnUkd3r8aBLi8j6NI9+7ENsROCm/6kIeS
Twe7+4v9T7tDGWk5dy3EHfTey2CjHAzD+mdkwkatevo2xgHGZLxptzNTWjv4UqRkpCbQ165UFs76
rh27ADx0WhK4RHAUs4t9tq+uX8zXI26u5Z0k0T2nhSBVwILPZFm2dahvqMoFaPUxp3jUkcbrUNUU
GWFCKyDiNJRxUiFXFbWq7StgTQjNrTiltSKLT66C2D2sbStpp0HMa0+Glfk2i7uTzU31DsU94hwT
8OLW9vr1NGoxefgwl5spCaOKJ+0OkJvAf7WYunqvHMK82r1YzgTMwaplXuJqvfT6Oncr7xXWowhv
74Q1J0ghCe9vTo1HLipCPmH53n81uHeCrMFcnxuIvSLQ7bKhnj3ojkGadpC8AQs7Ke7K5cnSg65B
7lt7CB9w+oOX/n8epKxgwACtnEU1e1GFvFHftgCT2IvB5QrAPdBMNKdNbGk3tPZZW4U3tbSC0Zjn
pWvJ8J2SqkgX6qEsh3AhfguWJpC3R3pGLy8WyhxMLhhl4eQ7f+aD72goiYPSwGOW1lYPZJFcxE6E
GiN1tEjmBMbEbji3ve7w8yg/s2wD8UMWPHz0L3ooHthqUTYqgm6uI7hcCD/4SWvwZ8fr0AK00Nmr
kCcV0d0tev/w2EIM2IaBbfi7NOmETxrEBoSEee7kzEuDcTjEubQMB9uRc+C1vM2Lea7ZK0T4jCWU
d4scWcBLKOqEeSKlbN5H8MIN5f10e31v7WEuhDI7b/AlyE8Yn7aEL5eUJd4g/kwSH7/Qqip+17mL
WmQYB+R4hZB5iXXyKGATQ5HC308S/c9bampN53aT077AiKKjcXDPXuSk1lW/rGHhxo4t/Z0Wav9S
YqeEsdCdwuJn3snGNZPDTtaDZ0z9VQKTVHUvqma3s2JODTJIPsSa6L2XK8osRPVWKh8RecWi7BcZ
RfB22LQwkpoGOyaJR8ISTWAVERbYV+lYlQSieW9CqkmwCflQjsFZVddOsP+WxKZFOlkFxGbEB0At
mtDvl4OMoCUWiN7FkaiyYe5+GXsyvY6QKBFl+jUH0qYrGK7SCr7hADZfPgnlCch4OP9HI0e8Z7A5
GP1Ap0Sx74yGGX+K2nFLtPOZ4JfcdOGRT7s7PjhCx40Lblze/EaAO8JnZxNGuZmC7Zw7HZZY31yU
E4z6fWRJdKyJW6YQIP8KVUz8JybWMUbA2nHsxEepcq2IhzvLctZoHOlk32jFgCHBqbs7KPjG7Mco
idm3ETFL3NuSN5GWKifGOzPEA/fb0GcLhvkqOHBpX1qAi3klIRVbiyEFo4yhqnemuPNcXfjspg+s
ainO4RfYh/491rAcp4UyCF3ilE0I2aYsCtxnAhSCyRKsTARWz7Y52KSHnCTLw5OGn8xAWchmHn8F
R9A/Gt1ZxCrdoQEKzC6tqEvzO03ew/ddq7ZKTxNnDn8Q3erUUGqYrP+K/jbMyTE+emplDFVTDoLl
hYDmPGdWEDZXTi83y8tfiqATImNELT0HcxGD/EISSHh7qSsm8IOyZV5KGP+5vLI6yKCQQbhhIfy0
FB7Zs9sakcQrLtccy+oZ8Km8LqHSXQLiQunPH/GLORrI0874Pe+buKACxmaeCTA5fGILIF4y7W2s
Z23TVXvwM5u3e3LF0iPN9xN8d/SdcAxuOpALaq1oxiwTkRFZPtSQUYaBNf6ham5nr8RT8ASMHJLs
xcpUYoL3OzkTrYABu1eRez9ffzt47/HeOEh4EwUZnKXFwy40Twt7BlTcaCMHAg8Rzl90SNVXf5eb
o8hbOAtDGqEeANYIQZK4YDXDUjwccC/a4qIPrd2ymPUtAvMdFsEGcYUv1Jp1GCZvTydBsvqG+fuC
AYnMF0riUGtrbRslNITi/meDyCpR0qSSTUrTIcSSLCa9Sjt03GVc59HD+4zMuoigZ2rhHCVnoAQx
MlXhdfOv39uVlajrVcmoHmxq7y6mw/7GdlDPYpLgRl7aT6LMM4rl84CBri42+pzwJZ+JJk85JzIV
AthB+LuZnIQc4ytVA6wSM3OuXYM3FtJI5mmKbUsEXqkV/tl+RVWU+flbbpMPdCzbqXTxTBtpeJC9
Dqlon8D9qzc2WxEHx/3++cG0IDfacBbEeIPwyRrOlRYM17Mz5NWag0dsL4b8gmuxLMcS81onN5df
L+6bgEus/JBv4FcJlqaW7QfrgNgMOdl/+dEta9vS45a1HHRInCTOxezfhV2S4NejHtvyndaxrKpq
QGpLWV5jteY2by6uGK67Bk2hvNmFtVCA5bGYQuEL9ZXjAu+n7ZCJPSkGg+BZa1Vacw8duWpAflip
6dlstz5Sbx2GLwu4DjVP8FUk9og+HNi2vaPOPb9uUoCbj6jkd1SWdfEtAkg47D7fjyLSUHSx4bI5
srwDLuSF7Z+UwieLrFh8UHiJYzY9LkJiODOvvKtQBl+zVBGCYAvOHwp07dFWK7+ZJK41SeKH02ub
whPOq6B3SkFScfICGbaTFfkxWFlZkX8BKNZmKaXsdLkRIleDgzwLWpbC5msMjDn6Gq8zjSzYQH1v
h/1BEdpy3YyA+AqvfKHVUEUpM+d1QBRIky78fF0saAT6wxttWAzKCL+0l/SQa/s2IOnRh+JwFh7Q
l517zSxGS1PIwdZu4Fnz6qUL7WhUG4sAjSAT2D9JN8jxhPYO6igvAG/ZzAJRqCY27Vzo2qt0sDjf
9I/Oq7qejGEDtneBirQRX5kF9Ixp2MAcc4cp9hZj4vOMw5A0tsvF//lrEDmigev2IMTHMcHihttM
gITk3ZDPPbUjDM2I8FLSvDvBrsf/VOcu1h2ycTkCyt901SD+HyLWpsHMdgoWN5AffESEbvsUXUWG
E4HKANeNAesvC8FX8HXenvDGItXl8C4mMVFpA6+YHHKlEBU6fpr5063r25lNyC7fo+igI5dRevuq
RNRJC9wYsvSvyaA4JpWgHAuNGeizrzu6Z1J/Myjoe33pLIUARD3phd03m0UXdw93Qb6jFgP+dgcz
xfGRQ+ZEVIj3/dNL0/khh2FWCEbudRvg5HsR7e8euEK8qbH+6Q0IbLcKYsv1KFV1zV88iUMprI7T
/3HLoEm82HK3UhQUSWLvl+UIdDqAyZr/NUBVBCzWA7M3ycOj/Q7CVSuEB1fBNiKOUuWw1CmqCpuF
lmLHY5/1RKAeWv632xEPmh7ZeJWqmNgMohIbPIwT62oPtDg/LIaKmsv3I8DBnYm3nxeU93GBzXha
FA7INTNx+e3U3JisFHuXmr/aACMGiTUiDaTr6N6jeyt7DYpGUgaqDHb2tCevGEN0DVjRGylamO/F
Y2XDZksDg+MLx/nNgyCwaPY1kzOHFL7D4QEUiVFZJwxgRY1TlKmgwCJict67tYQzEC2gma4pVN+W
meAvcgbQ69+RFHOoHjoTsn+W3pqnCZfI2tsilRbh4S6FxuCa7nqZy3y9hFQwCBKY1wKyFekJ0gmj
54zSXuWSfrHmavVWM5W7DWLb29VMqR4EgsOGD9b4fdc+BRGI+g5HgSuprNal2RyqA1gQ5CJxs48i
unIpYzusG3UiqYEGaJZIi/ujKh4kkhDOstm+WAdz1Y7xB/gGd3+kdQ5f1pJHDwGzbfLaMxZvSwdX
4l0eMQyIn8U2t3IUGIVTySi7si4S4gogZxc44uLzLMsfFoJ6q8xIU2T/AY0mKwaFwz8mSRPtOiBV
asdvMdQXAa3/1vQbB62Y99bLNJzU6uv6YTscMqaMsmqXelKsE+TKH/MXjxegv+HTabZYLgbuMehx
xWc66QqMGgrVu9HxLtkAzQuUszFGSB2/TZV7WRelEh1LCdn2lz+UV8ixYOfA24Z3YJ2p6jDVGRMG
zfqJB96A+EAu62nHsJt/8pd+rY8lXYoNxmoGZnkhyOFvJKLc56lpaXtN4iN2pBHGah+JuPG+JfLR
/MzVxRTWRbmLrmyzWQ52UhHO84PGbOGPPvSfWAQMet+KTIDvZuQU3sSyYbzGXnpRwCD1UnX0+NP4
4OErOJcUR+ljklPc+G6kII6Dksou+FEbE93f8J8ShZoW5Vuqq6vQnyzduuIbaH3BJ9zP+IiYHqzh
6nAV/Cmw94OGoDmG4vZ/TlI/eAkVS5OiG/vDMIgI1tKQyRK9ExluxOQlw+BRYKlpumT5L76IdPXe
nhG+b4im58Gqc2wPfs9BlaIMY9kTv6GKKlpAdkRFC/ENr1vyn+suBONgdnqT8quKOiNO7BIe1unL
bi7xu7GcbEbbfurmaglipBJ3Liq7CC7gGvOtxL9if4CWeLw3SH1UrJC89SktmqYucFsalHLIBluN
SZ6QWtdXYMMO5yEqq7XfTf2BNRrio/1yT0EVwr2IceQoYiv7zq3BYSQiBOFclogG4TWBkx7JMU1P
MZf8lLLiTjOPmBDxEl7RuQjIFHyVNdLOU+8iSzlmSaAfNnWZkPVNUpCYm8e1C2aO9QpS+N6aaTs0
+H79+QEzLK3j2vNSl0s4JnIGlzfVMW7l6IfIZQ+AjLFpz8goM3BmI4zY8mV1maPwyPPDtZotENuP
WhmAexyG+fdde2O9kfDobbR48BJSoxFKw0kGI1OBlusJWuTfhpXzjo4JiTBQWg/0/TUiRHTP4hag
hd0cM1i7M1KEcfYwO1cq8AqQI1Da07JIoAsYJ9gu4KlCKz0sjMXIczTKfhna6i/ghMoln2+ZraFb
GOZ+Mao+sHkX1TfFTe4KttjsqeVAWcaowQnmub65z5ld/u5OaLCv284RAbNGzDLJG5CW2ubuNaWj
orjyPhl3oEeGSJbI3lhtX4lBGZ4LgYh5G0tfCn46g788ubsT9MA9iwtQ78izM3+m6CwcXyiZReDo
CalUBnzLICtVflpX4VxaJz2Xb+H5DOsS4Pb0JypPqkOJl/vpzEZfJcZe5dZeqGWahIZGyf4J33JA
RjP5mRON1Du6Yesz47QWMQlYzLUTJcTwfffoYsziXxbPkmQK0DE2YVywcJXtsZ1HOPnxsDuZ1CWP
E0vRk8KUh/tBRLoCD80EFwROAQ6An6Hu+mppgeHB1gvF7R9x0Uq3G2uiWvhYS9+pgi3RiCGvHoOR
NNlwdSLbPkRc3JHYyfDHxH1+0ES9UoDpxXdOl1hKChXeNwUtFhJ2ai7Y3VBsaXW/C0vFmcLwNbqE
glkvvVDafncpDazmZe2l0571PaW6hq+WdDwUUsx/qx/SB1uBVKidXgmPlIMqOrMTIMRULjv6gfAA
RQghwJ7gf3c9zOdTaE9nRPPzT4UK7LwAwX1KMviOpA1JX0CTS9yKivDcBLwRTpOgYePl6vFZMvAF
Q7tdzHcBC4fSn8A6EcurOUATtLE+L788bPlxlOjdW/TgqV7HzHYqkKbjYHTkTvL/4xJAm9v4OC2B
1RWmlEc4LampAinwQRnkNiBRaaak+oIhMjtDy8KcssTIUR5X48TkDjL2uIkxB/P/my2F1lUUUF4j
+090w8MeXftr5YIhnJFz9YZDW3CImpGotqx7Qk43W/xe+xzV4ffT8jBg0aXJcjoIySmpVb/wBIRo
tPQl2KurWT/7pN48W23w2wCQNRXA1TXkwfgRRkZ+9jF40rwTd97+aNKbNWyyI3jUMNdEhwjE41ym
oAoYPgklQEqIVtrmlJhwNxmnGRz1U5fE7xXpojJ4xgRUJ7qIulna0DrMfPyARxo7lYjf5B50XX4C
2ECO1f0FHbEakU2K6GHHQMbmORo3BYGHPNKU40oDkR8PYcBe2qPExrituCOpsOoMo8/44vVCVSRg
5S5alO2zVJBEFDcRLca0tby9JxDDdgdata8CAtVlDdAb+xCEd54u6F0padMV71NnEfLTUWA4Z81X
J7V1cgVGF2DqNTnKq80VXviJgrz2E5aHL3lhhY3u/F/djKnFIFWtAXmX7+BCwO3kQLbf97KeWiAZ
2jE2T0+bh6iLlY7XLdGQZaPsTZrUeu3NQLFrCON3wsMj3M+/nh8L6cqKwqjdmfQqISf/Dvnd3/mi
X37NJLTR8R87oDL+jcAsmmeE5lwzfWdVomFzd8F80alFX6udbJy8n4p4Saud0c9acX45B3rq4mSY
2VTIjAHFL6Ql7Ax7sdPODqLsEmIDScLBbuwPiUbl/5tw5FkiUkNbQIarkLGPuGAW44T5avyMdQ0/
BxeiYkG23a5E6bN1qY2apPfCqFWi0OTdbEasHW9dmASHej1lIOsBMLRtpTG2SrRslm6CQFN5Rs5A
+cK8gtl4TTKP0F6dWKa96VAlW4UJXO2nkL4ibMEP2WLQymuooFG8WA4pZH9SPpj/Srfb1aPG6Lvb
MCuXS3BGtoNmiaYHZhpV+pSix+YiduUG9r+mdXNpi5GBg8QM/CJ/vlec3Qx52NM4GPOpJRbKGY4M
vbBqc06bfOKVp1q/06IwVa0UtgltRf/sjxtWO1cUMAZfYJdxU/ByM1kBjg27r0z8acMPB5OQz9/k
9a1Eqqxr1iGGdOXJbn/QDiBbCCgkMyzaSxYzjAofhuc2MVPo+oz01ktd62pW6h7uUM4ih0G7n6tn
Bzew1iLMzfQJP4j8wp+3Ig1CKAL8aUAmP0prJCKnA9SA8ti6BKtjALNPMJDJEYq89BSk8XEjyFT4
J3rZSvQ6k0a8Ble2emkyLTk2m2mk9jp+Tr4DEhWjboTuWTytcr0W2fVH6N5/wecosjkYw7UIH8PO
vktKgyKJRQAVJxNvPg1zoSBjus1oZJQLGx+b45ot+98SVhJ2mWs3aRJBAc+vfXgDZ2fVXDgPlRhe
0q/6Wi15VnytfsbgyjNhR57Fsv6YVOtXoBdhqoVYiplUmq+Kb4j/AzExpO4aXLFQeo9F5FXYI82X
5tNucUkt6jGW7g2BC21A1gVQLZQ2sIWYWOKyvFZUdk+sKJVQ2Heb/Z1NNIwQznMJYS9v5XXe6ToO
6wxVAuklbqaNwlSXcbcKuqLhRLTxldUCyuueAsQi10b6wHVkL8COKx4GBpLJExgCf3OZvl74l+Zk
DRavVRR7i4BGrL3nZbTrtZCP99q58slYk7NRD9Bw/ce0zZ7p0dl9nvAt02oWW89RlGOh0E9TZTfi
DohkrWjjGync0zWvJyrQHSrFTLhNmpGFCl6auVhhOPTofGiprszC9DB99DQo+brKDSAS20MAsNTv
afEM7kmm7YuTh3+vhDRdxkEHTIqZoBKWCR2dAur/uBopJMx+QOEKrjSG6EkDGTbtLCb0eS1197OC
yUb5LVdYthzcD17vzPMTXXHyzwl1tkD0M/wkKJVOt6PwjmqP8xTFe79H1As1zCQYjEHgaSqFZtVD
LyRdxFs4X+lhEyAKTNKBbmdcS6T9BcxUS25tiCbj/RNYWV8rL7/krF5DTEQRKPRN73tNUDU+sezi
VWDbznFfyZopZh41ZemFH7dCE0mSqKqgyPORZC5TuqEFSfFDvPArJ6jCtFsX+Q+rElcGeqf0BBs/
rNTjRu9YA8tJCr3rCAg2QKVqidgq9Xvfwk/Z8DraD1Izm4ptdx3eF7Pm78wGdZmioz9cjmv2EBYc
SS8ID2HLwTYRoWSpljlTWxJaWSvbtb/lBJIo2PE9FMj74rzjLrXJSgAc82yN/oxN0ghuxzfgGZDJ
tzO6s3hSsCZsfvhBVuIBa5QkvPFieaw/N+8ReqBlOODrepThyuH00DxJWkjp/8C5PbdNOHitGJYq
EMYDwJOwZFzPTJEXTB54Pthl+WBIcngO22l3bCc3LnyRs6kH47RQfEobrkjG6xwKA6j2ne4alb3J
p9tAVlsLzpXNzCEl/bQI43Ua5Njs22lk2hrvE3letG/rUwb/BZXDTlDo6qa+HRheaPM1H3/SLpjx
6DUTkXQUzvWXxD4SgTjuGsbykLKo82lzqqFxw+27E/m86t6AsgajT/b28vk16BOWbjRg3rlGcFg2
WkGcLqJuqWFG3okC/8gXQiiMof17F3aS1m916uzrKTiqIF+zkG2XfO4BbqqKUicu1cZ1PyiiBYM4
Q3GkpV5JgR9Z/w0AKPuBSw+7ZHdoL/N6RCKFT45K0nNhQGQ3mQR9hQc7KsjTWxW5nVBxADfXia8U
OIHM6jH3DYktyXlBb93OwGVWIfKz65UUXrcjjFxCVia53QAt/JXdSAIsHAYt3nB1DJY/jaxSQfjj
gKMm/6n7e/u2eCZVuuj3qdKrk+uDtN9/gdumcMsjqW75WV5OziwRjCz3XrTahnHhOap7T9bKevsn
Ebr4aAfJjN8xwwNgWnD1LtAJO7DiPEQTexId628KPWpleTMdAISHcNv+Q0f8nfUtuFF78GLKP7X7
+aKBQL5Nq6oz06jGqR6ZsWUVvcvrTYshiLx5z2omFeP4rWDP1QlCGrzw+BN8XdhgbGFF4Mj7/RUW
mVyMPg9eI0VFXPZJriX72XHcocrRJxOJehzDd04T+gDDq7iVlLaY72q1bi1P1MJ9E323Xq1ZvVAo
bWSqKUM0dstVuYDLND/+goEeS2KwbPJQmlnXgcAq74RHLzhrwMRVU9V5rPusXlQK9gwc2ihNYZD8
3VfLNPXKVdd7Vq2y9oUb2YYG58Oo1PymTBWHo1e13i4wuctH5Vl3VRf3cfRtabc9hr/dbq5kxD0a
djw9DSRfZPLwGd/ss+Mrj5JKf8/7BiWbE3PUcbShkq1Ql8ExWYp0qGg7bU2xrFyrFT2kJTi1aA3H
90kkAjN8iUyr0rmzlF4vzhRfzwxi2NM1sg35KaWbNqEnZsbs0A0o90L9g6oP8Nqw39f5hQqMX6M0
ZHifq+EcYSncWOhGPYN0vocSGcbsMIF2aDOcWggdRCfkvQ6FTvYqO8EeMSZU/iMbjjtjKH2NnECy
HM7Q/sKndofx9cqd3sw1nnjgfiq/YBPPiB58hFYYAzJF4vD40U9tledbug8yLCR9BILkknlmwA/m
PFcH8Kk8eHj3lSn8cQRoiFnFvxIPiFeTh826iYf3lQIYDUeYJeuIg8GXN/gbQKMNxrMY4C0R2deC
ArwWp7YzI9BADlFLlTJSJTYwRdKAkoF5WxuuLbF+dEIyHXuag2Zyof6z2ALtAsAr6+iJKC3mBoqy
/zl3kzoqulnNDZB6rK1NXu6w4bqPGDDkwKnNY9i0wmg4ZSZXl0AkGSFN4i3gPDYyGgZ2WjAr7x3G
awUWAObV7FOUGZvLdX6MJn2NIVrsSP0WrSOnumKfDLyBsZXDLCu7+f4Z9pHvzX/KXgj1M2yjJKMi
uAXHXG9RVieUYbZbvBWcQHUZQNjTqH3H1apLlz08fF8RBlSI8JUq0LtLgDJfk3qjIeSojnUJj5BC
dgS1WGKaj5z7Kysl1C2aJd5UjMG3i9MWXIVcsWTv5HUAi56K7XQ3gOL/W5ARW9uvMYm9yWanBzDG
LxnD+w4mHyCdlmLUaFp14KRS8Il3OjLZuXHlTYdK/bMFmmhhGTGa7RapVb7ztMPULtBHfEhN4BoB
8jk1aUtAuhSPYLwbyNIaZUfqBzq4mTw+7v5zZWWUfKLyixCIa2aF0emNlwTCPycvHca8dXnQ1mOW
RX4mfGCGTaYZ+2FKEiDWk9Yb+A0SzzkiJQbspSE+RD9HyB79mXr7s6ia+uXoC0P4a2K+xhud053N
u2fNoXwq5qfoMIBGVpkt7ULraGaDqiQj6fTLPmWdabOGYIXXZbgn8qLQUcuBtiZabS4xJZCUBIVv
5aOL5ub1tr6ILHxVtX07UTHTe4fYMtf2xGXiZoxdTLat0wB9jpV7TxkCXw5/2rMqKd0rpIga2pKd
ZXNBZ860qOdlmwjjwNefYIT8X3+1efe2RLZXa8IkqqpV1zmfiqdQ6Kz8UwEQCyO+rNq2CrT9sKyl
+4czOfQI+LGy3WpGSPgBbxTrmSzp8uj+ofkoNqFrODy72gEsl0DXW4JIv34+arQQhfXa6dh7ZgR5
lRSrenAe45PbIwd5kB+IXVfii9DvbylXDjQESN7nsHS1HutRHDMRvO/smwmlLFh1o7K0crn6H82g
JluZ1u5Yi5Q1n7vQCMV9ivVaPLDT+0GwMAR5qtnVeICSHyPBfFPsQANAFd+pe9JQeEbr4dvfz+lT
I5k7Kx/qi3HROZNMELTdBDmU2qR3nX1orHOv99yJ/ph4+I8h2JkBCkDYVza3zgUoM3knTPPqctTs
yLhzzmzBlT51R3AKA9eBPbBul+t0lPz8A6u6ovNSRhv+MqZVriC1Y8xmiJOHnbNbNi8ll8b7OAXf
mki5wocZWOe0KBu8eknKW15EicmVqU+tGeDVFxu7+3ICjhlh8nfMYRR/k+J21r0Cp7ECpbW+kQAz
mYTCz//MAIiJ5CxROYAKagj8daxLyTrYwMbSSBvn3kPLYYrcV8cL91g/uhIynSUVeI4C5la/diFV
jPGo3Xg1W2fY990btN1XxaijZbKATp1CsMOYlNg6Vr0R1OMlMuRJjiHF/+2xppJaEc7OzuN5r0DY
quPCqRuQ4wZr1O9a6lPfwrgBFTjqmNaQksmmIAs2neDCQsKpU7fwCwFtNtzGyzeZ/MNR/KUhV2Z3
8Ky3P1XGzLrz9oBOt92Mcg/vAy3AduxWkFclxa9SCoU7HWKiuoe/7BpJRBaMhXpx1Ys/NsWHh1q0
2tNQi0BbW5KQclQAwP7dgnC0N6YsUXnMv75M6xe/YrbCfXjBLNvW/0/lrtnYKZ8Qe9X2upEq8eac
q5+WgkR0UVx+trlxywZNOJgu2ytJbaUgfLz24np7G3dojeZhV4Y1iqxxYYOQxO0DMwX3doq4V84x
v+15fuLAJ70D76ZBBcZQbGgyXo8fIaavhHRDW5TFP7e0piXzns6qaWpBB3o4l2LnmL50A5YbQz+w
wPZrxtHW0JCGpr3b8yEW+gWNzu6Wg7zQh4aVHu0l62NUa2WH24Ot3bkMvorXih7PCbkCdk7Y/df0
hJgC6bo2ZrnZF10rz4EHWY/p/LXxnz/P5/2LE8SLEkRla5UZp72jU1p4jbMEfrSdL4o5AgEsAz6j
T4e3COzn9EvivYbPZdDltCKcDInIAdrIihQskCC5O+MRQFbJtAM8w4/6VXJkeNUzISGs7GpzbpiD
Zk+Wo6iBhKE7jq63ad5i46BcjjTMZcQ6QLDiWQdI0rTp8azHzhTQqIeewFHrBDsyXJOLcNMxxGUy
Z011eREWPbE51umW95SKGKIqfZ/dYjBu2nI3n4SJ6Ddh7PNI+AhqkDsBFjrjidwpLmiMTYuWKe8n
MHTQEAd+WUYfXZpeSPx27+UioQB6lBzsTsJ3F1I8SUc6djSvUTJPGLPeyEvx3Cx7WPqJfjRm/ILS
RFBli2AowQK0PfLi1rjujVPjwUaEcuQveDislRnjumE+CPXkSDs1HvOxm2gUiilF4tswz8aO8+Wk
3OcKkfTKjLNobBmGxao1/JACFYVePMliSq2C/LbzPq86ht490B0ouhMMhz6a+JBn+8HWh4Ij9tYA
qBWAbJMKIQFzTG1xoRGd/fzKKlSJDfhoH1g/qxwUWJI2zOdHHfEMmF0kLsVr6mWezB0NJGxbasVZ
1RLCzikIY+SoCVrNhw1c4Ol2E1GdQZUxewigm5LYwKpeed8uKmpDz4kS8Ax8gUPJp3pRLrSP12/k
Rd9gj4toqUFu/fo/jEJf67zoRXU/eqgEZsMD2304rKTt0CxVrK1J64/6A/2dDKxAxpEsIxpXZiJ7
pBov7LKfazpaCPlF1xWAR2jaPUvZBQrON68wPiMcsWdzXX2Bb363OEgchHEY/FiYloktt0q3O9G6
CnRGN5LBvXN8nJpZqvJ4lzJZgRKL93qbPxFSgX4Rgy7M+SZ554GHcYHUqeqE99YwSWF4A0EzXOzK
sJs5nPB4sXYynRj19XGJW17cOqRH0zUXLuHvLv9HvLiwfdJl1pEN2nmLmjudXOpN9W9gazF0FEXm
Q6mxA7ytbv3Okf6BUzYGW1skXVta4eHsuBHp+fKp7Bj4osTPrljULalz4NPbtlySKvGr7W32iyB8
ur1WnuJcab4Tnum6ympmzWnDXegQaPcBOvH82tzBPH+xVVaZR8qMe7Jw8JaTiPzUQrb009TW8mSn
Fo9VYw7JAAGyrocKRaEqRaYsufpoiFpq9EABFGurHzTqJHtj3fhiZCAeax53OXl6FZVcAes3rMHK
Bs8+oX7hmaUDn4CxzjCcmHDiXALk423nmPZPJcIpNlZ22qUM5NZh4QGnV0DzLQvtRWcsQXkCYchX
+0b1/V3tgWDt6c0UB6+OkXh565ycdsZiSzDWb8QQQqMQWfy6pq3T5ucm5q6oVoiLDWGGbLeQDbEc
yBGah4cCq5Ha+FFG1DXQI+FnT7OP5QOZDBMjLT50MX+bXTsYj8urSpyT3F+F+wnZzcYktCuyMMM7
KcJQF0aDpwZsstzT5g3MALxzbC1Y5HhqKbbNHoJd0JQQhEFdXu7wtIiGBrTc9tdPUhl0jCX576dg
OkhgXBTw6WmK7DGTT1cTdxgZkpNCTpKeLyXc0fIup3xvy8UoKtBvgYvxZ2AJiiwq+YZcVNdxPA2z
c7yf3oeZdcZbl/ADOXlJWpEpEGpeoaw9Jmw7bUKdS+Vkxb9Ke61HdwgsezwefEBi6kPMNgxv2PRr
AOPuDFZI9YdyyRVqO8KAuMB9YtyEJfCj9y1u8/PdOMQIDScfDZlrLGVMF03Ktse8eke8BK3dabG5
qAcq4FzEQxxYqJAalOMh++Q7nzPZ8BXfBQU0XjyowqgtGchCaqt5wRnBWXcwWfQTKZF+Xw06D1xI
DWPYnm66NfXtJblVxaAURhAcim+DsPG+PBxnZiB6M/PkiaM/Tn40/jqTPtZ2cN9jrqUXIS/IoMnT
GeHHMSiqBHAYBBaC3Ftn6HloBQLaOC3iJNUbjLlgxuUf05LalC5Pwb7KCBVc2jOc8COVqHXs5HS1
vhbyQfjYdhjS0ZAvkyCj5mK5O4mS3H6h+UjsFCtxFUnteq7QEBqltnCMMb99VXjrsCDiAn3VFiJ6
WLsj0SZHbO1IqIss2E1KegHNRAm03kZKlscuek7DloRfx7KnTEAl4yHy0dICmAaBM2KWaERPad9a
+nAdkFM8pjNSV3N6Pc4oL8ZXCssxXdZPr2H2BHluezkY5f+FHqdKuxz9lGko+0IkpJPdXH1f6b6B
AS0PaSwg6rjeRDX2azmt74Wp0o5MzeBpo2Jgfyu1V40TDnZanQoDpzELqlgBkwxLOo5anGjSJmF5
Z4ozN8gTpudhsM6rqXb05bBYjJAsb6ljFpFPjvcXAqadQcdq5BCYxACGtojx0+C8OjctFFRV5Z9S
YVvuE0jF5CG/zogkcfqOwvf+uEVk3sk9TxzLnGljYN1r3HZSvqe99byCvr63QGoiVHMNnjGPYc1a
oOMurULpI3zjtyB8ejEfvvKFMjVmh7QFicfv9/gsCrJ9HULYek2/42dEAa/wiZ/muRhQnYi9DlYI
GBak3MuPVastMxAxKcybcMi6Vg1xxX/y5N1AbPzNrKeFI2tnXz4Jmy491qYl2lYTGbBvRtSsxNPA
j+Aq6ia5EeHp+Vm90cyQAqFthEq3+RcZ/x3j4HOXShH7K6VTKv4QjwPlwum8No+zU4bUfc5ntie8
U587kDVD03ZScbrVA17XtnAJJhM0GbWVBCz0HvmrIummU5ibyPe8AV3l9rc8svtGRYobA9DfZMYb
YKCrfgya2jPtIWjuX3+w6fI54ODQPm3YqfBl3Gh1Z3uDBnPniJQMbH9EzfYkT1aEBVp4S9Ujp9hO
YTPd/JiwK6U59dAva8imASsGrOyMMZ+F8Z8SISrIBPk+TQvndLMfo2HsVkAE/z7AMsBH0oWv04d6
MuMZVbqa4Ouuj7ZmlyfuMqcuO2JXNGkgL2vDz/7z9uUhlFg+jxeDw0hANZLPoDTlAONYuYwGZt3B
Jkpodq+CRvpzUtVLm13Ya1Y+LYa1NzfsySVLFUejLAQyZJUzlF7nQ3BotPf6W2QrCboiTbWWzZi6
q5fjS4iQrMinPQwOT/qz1Yx8fo6rNA3KUGChXljnadis3vVbhenAxgG7cKgn9jBtj9OyttDadP3m
HT104nC8HT/kOdz7ioxK26PpI3EJg3ybPsOWcfopIF211FFMRLF0vHhPOJDECX4sEJQdaaIcTYTU
zvuLO8pUCAfGPqlH69hp3zG/aeRUsZQHQurpD2CVHMC7+D0akom+PnqJwcrsstTuO7RpvTK9N6Bd
rLv6+KMy3WXaLFdF+OtMYoyE42A45VzFqw0k2LNI/sH/EZ5PgWNyv3x5KFKJd/4Ecfr6TXlKl7aF
c6wWWsmPXSVAr00+iKUZaV6SEDMTOi20pNu4z+xOuGdhB0MJo0nJ6zVKBoVZbsest1xosK+EwJTk
4TQsB5jR7uVIX2eeOXVs64+/rzrec0aE0oIFd30OF1iI6cKkWPtJnvu/KCogSZUq+qkad8/b5Ntg
35CHvQdmPDKdy9a2HRSdJnnSTHL5/XVcxOuB29f1e3QrUvySI4yAyudKNrsZwCJ9RCPzvMRhHc7j
tM4WK+1gR+xX/nxw+e5Rxs68YrH2G1gWPM1+MOfSYEEh5Fpxk5glXHTAgTQ8uRW1MMsDjSBIPyNi
79nKM2+8AXK12dMqtLWAciO0MfE6sfG9jOvjP/OCOHAAWm9ggWwoLyVZ5fcOA7Ktaq3lUFO1xesh
Q90xyvPJAfJIdWqdac9pKffL0aNNR/mLH3h+zxbfEhSrZfRV9GYwihNVdP8P31C5t23Qf3cqZ2zi
FlfYU7yE0fN/9szSHp/HUvOx3tA6vohJ/lw46fhvwnopcCl/Fy5vK+E0JUhxlhQMcNuWrTGSWyss
L4uaNGWHMwy1ENxbeUXZ5pYSLP8iF3kxKRXIr8V6ZBnDhVCN37H4yhFn2o/Th4CK2uz1us78hkVB
NvhZ0qYKjNLYGDG6pJybLPgpuJosn7/Krg2JCqr91imf9AttqviamQlHiwMtQfF5RZWU+HIMNf+C
nXQWF/lxzQNyRYkgmhGqf+fZ+1k1+W4G3nlG8yu4mwbo+hS4rWWQgX+H9Xk2PP0d9l3U9I4kZ4CN
c6PffJnlZSKnzZjFoU4ExdPOwjuJgfxXKfkkwZN3fyQkr1BJ1eiDr+J6z229seKuwgtEqD7gYt6N
GTyR5edjGrE+ji6mh6JGSDn4o1VxBrDkTwuiL+RLPVccuJGsSQj/QRIctt2lglQX4rrl7P2Yqhwy
A3Cb2x9CPputV1AZTR5vr74el9I6bzN79TZ/OklMIEGsmM30+XG99lvwWG+tMX+KKPrleVyIUx+c
8RLf9cE+BD2WukYJG35mtM7S5B6KZHJpobPTWsnd2eHHz+D/aJ5jjQlIXHHJiC6if4Em2KmGGMJl
G+YJpT/Xgw6H561wdq144pS0jAdp32gLV4wl16f0p17bYSM21htZ7D9p0rvE4Q/IQm9YAyJCLFUj
Gw4ff+a4+MgUXNZo6+JRPWC+VNNnskTzKMQcDFKFNvkiq18VWVTggYZmIL3rbU+/LvpUktt3bF20
3NFjRsjOpJhYmo5yiThUa9BpK4jbOFeEu0YCMXUEyBlZkF7yd0FkZENEgkFcm1mWKm56QPcQ8xtN
f+ZDucOx3bKgkdAG459e6Q/qVHytCwgKb/020OLrgO9Grsmp0Vl7sQRWcbyeY7eXDd5DiDvfYK76
vvrrrnslsClthZc11UYA48VAgGL//FTz73fjTYkgV8H0eT2/FriAKJIZdM9LahqunrOKvsryHdRo
/7NWUPHHUxS5KIKBvc/RBi98TtGDds87BmcYRezd2IZeHnlEw1nTtpCGIy4As7N9uv/EsHrM2O/c
A0iPkUBj9l0bB3d+JIuxNiGVIG8lQeEG9rv0C2owkpubXQB8ynldMhjcK49+O3uMISwohSD/OxxG
jnkIDbjWX2gdUgl2/Cjf2LU/rnWujJvJ3dR9jLT4kqo20/kMRuCTl/uyaixJ7z1yMFjtfM9lU185
T/dFryyJVUwuzcAzGv+rHOEGI7BMJqfMqu9bn+UjeWLMSTBeRgYh2meLg86u/YTYN98dA3Xg6e6m
YPEChNBi6dCjFmHugnEp3/PAAeZQQBKR059IwcB35awAgbVLo3qcyilP5PmbiLXOfK/wVvoOxnEI
/L/j7DWh11florDXmHjiORgwpKzDGP54XoamWAKxlfCT9dXcbYr3nijVy9WN5q0ipV1YJVQbY2l7
rfS8ll6xcb7enAC28MkYFKdEU/7Iz7Ihu35lCfA7K3CPA9rd8ACt3RRikb+Eh/3GzBLc04uyLG6h
O3dWkyhySP+zOuYbfMhm1WD5qijlEfr7EfRFv4fZ+QdCcCFR4NHW1HIU0Qoe3QSZDhRFKyl+yuiQ
p4ZO0Ehzk9oiGrH22jeXmTpqkwbuHaG/YBoJRCuOA89llmAVvouIr0O1NqgITv6T98YcW4na56nn
GtIl1Ybc1cmfeve6a4YUeZdeolXuBybKkxA6Lf0a59H7oJvtjACBRzA3uJyR7K4MIqW2lJwUIdxg
ZwJQDzOat162wsd+6Tqc08wUZkwjUZWsS6st87H/Dvf5wa+4HNRnP45RvxjQ0iv8KHhJdQPrNuaV
5C0PSewfnLpBD5QYO0wzJaZOf3UK5aPX0qxhmCoAZ2jqey42NAuduELL9953Lki6VdgrjRhwktV/
N7a92fphcACdn1D/InOjC9qLtA1dqqnH3x2CQ4E98mD/URYdi6vBCezR5fAG41PYmmS4VUXRsEs3
nJUW0Fjl5B3xfMzQzb+utXqrikpvGwsWhqmoPXeDhWcb/o6iod7kh9hy5oWksdi5zx0gL7KRV5Ui
sGw6NCyJnEGsiSIbzxKXs8FiD0gQUjNAO0SEj5qfPHF6/KlcZDIKAb+nHFnfNNRopXj51KvOtkFx
YK8PGkGJgsS36+mBIYR/MFueX/obr6TVwfrihnFh4ukZeSCE6rvGC8LWZflMXVZ9kvICsSRI32i2
A1beLhBOdoVBp1XSTamwzndIz5hVrdyYXyWq0rjU7pmZat78cng3mF5WQtdx4TK4dE+gWwnKDLoH
RcpABxn3aYzJu3MdcKyvv5THiU74Ed0YpxJasqQXI4Ms37CFx8LYVaK0DlmwKJwLC2myNhktG6BY
Ww/rvFSgXqHoKB7uzb7Aa8kH9Ngibmd6+dip0jStCuHk4HHhxVbKEabEovH30YXYDeVBLTcmU2qs
M/KcYHwOQeRMwcMWTKS76D7jWcmsxUD2vQ4N6w/9PVe1Tcy2+QoudJ6/jOxlEciHWjyDCn2VxK5i
ZURrE6/lEwuLTgc72YPHxAf/xou/9b5IGUb+A8GWNAn+BQNrbST6e2h7NbUDfsbNVz5jeFLq1HCt
1OlHNCm7qSr744BKcvOiWqQXhEBhrssweSKQ6AqdgLZSeoEko8MS/bvJruPChQCM8ATTL/pMrvyc
oK803jIFidDKu0i3sfWA6aQyoCGUP7LOxNO3wg/K3++Np2JuUDs9L/uGM+YWLcOu0wzqDmoLVXTE
uA/BqLUFsz7dspWhhqC+Qz7j15qkIzRsEfQbbDjCt/pNPtYMalMVYOz1ZsGcYZVkjtOdAujW0zW2
Z0F3CwGdw0vdjWKDaveJzdWkIcQLnSC6vtE6zXoBzdWjS4Ul78MIfOjVbcS1CUSFwoUDjM+UhxKm
FdEQLHTAhhYRzEBR/juhC6F2tPdle/L+Pq/FSjS3dE51vWeQLdoyygdo1Uhm3MqSLgCWsjNPicgS
rf5ZWRY+9Hzlzn4YvRNKaJwbJEEMxCa3+shHokPOWcjNY4F1JQME6hKbsIMVDrxa4Lcck3+XhA84
qQr6YYxGKB/+24xid99e/vlXdKNCGDZQAMFh4SzWANj7H0l3wfHRSnWUOZmtBAqa1+mPUqBKHNSy
aDgcnV3PqLViQz6Nnfy4IL7MqObwfWBgTtlJPb9o5tT6UBR7+E1TidQgBPSX64XW0hvXCByHGZZ7
ZvmRhFUN6spgtaId8QJV2n84BontuUG9iMKWYPVccS3dtEW6NA8BMKWjEZT3T/gWSE62kh/lLu9g
zrsUylVVdf7Og++ESbCsIhFVshOAkbrQYS0w6ktr7FHFS6zwhuJQRVKOwkDBFwM1heNo1FY1KiEB
SFxZD5Dgqx8TBDnIuh03mV0JOKAusCcZuhJANezJ9yy/+lYsBJrKLLgDgCY3heXqmFIsnZiV3zqv
LXTngg2Z+YbWR/fmAJUBFi90pdaKJQQZKiAzoknziKVe4uIt+oJxayBmvOJhcCP40uiovm5zJ4mV
NZwIk61TxSe/Y7Yx7r8mqMfdR7Q+wBwylGf/HPbeooRhbYgILP9hBFqbDwQI567WYJW/BzEqd3kg
qoinRjJIDCZ8HuDuRDEeeWsOzaPsViY8eCyeg/RKR+n0pj0+GpR4+tr0G8SwRNhwNJmB6C/BYS2I
e5mUkqe/sPmpTdgr8EYqQJZoDHJxH/kiUVdp1mcb54ztURWBW2e6q9X5FTQM5MQQeWRqiqq5cSo0
gs9iMX/Ncpm8D17xPwR1JMI2X2fehEisdjLH4+B0NwuKoc4OKh75ZSwSpNAJfXFYxwT3lcMi+zLL
n1FvFmFhETrXn30nY5VXpHtxcMRTy/mL4QbMOsyK2cAs1S6UAYQtL6/8XNZ8TzTS/Rmb3rNlVvYl
zqZmOjByA0Md+q6f4Vvx7nqvjKM7HmO2DMLGStSGzKV1ySxAz7kMAtcUiirjWdY/F9EAofNsPcD4
/aKTokevd7JZearhQkhSU7Wg3Iizg5L4YE9juRNbsR2mCViD1rANNsNG2/oEemd0kTTevwqCs+7e
UvjTyHviYXdWfMllsPs0/DW6Z1VZyRrKhAyfu0cI3apFREPbIthKZmwOkqHw3+iEqAR7+d7/oSwc
PvSIx7jAjl8ur3gvjCygCnzeGu8J/hRrbDa+5uZaX6tZHpeeK8SjxXPJkKfuQIT1K7/izskUbowI
Eaepg5so0WwnmALUl98QdBs7Jvbm2919eOAmwFfPv04hx0cafOr7orj0+ype9VUbfcl93QSnIaXj
5O+EI9z6HpEjZWrUpSyKZqp/kDEaoyhvOkh4uR/GyEO15pdRfGZvplV/TEgG1296Vbsm9IAfzkzT
UlnJRAr8qHDDgz+ctSzMvOt74WCwM33O8Xz+Bapb38A/DWNYxsluSEFIm9iJukRa34MHQ1Z4hY1D
qgDRldkZDNKgeO+/qR9y5LdUz7VRXWEz6LgUbj65mp9djm1rheV+T3YPgEPlkpCdnwL7r4dXzE51
R6KkTljceFzq7lY8nmPbVsbl2uFC/14RW6F1KgGFjYw5YWJeN84qnlQhL4RIx5N9qJcHA4YUT+9v
sGd4eC84oIBgT9or2xsYsa04t0QqdxTJyWeLUHzprUHnGJnFIoE0E8N4J9Vg8c8xKvZxRSbxI3B9
NYY99pmwyT11ybJ5tbmmGi78UT+Qy/hEY/fsEUYD/wNJtbNWj1pOcHzkfexy8BXmGOd5ondLXN2u
sFazprPlXR9VbUvRRDkBFjvxRXiLkWBebnNhiAX3Sfh/kKekN7tXoTICMn/vGPP1PT26Vjj7IQ2j
Ghs/jyO4IATSn8GAwJg2+xJiRXvYygC5iQ8aZr6wMPCmTZp4Kk2XYTvfecfy4wSqmrnB0vdITtpS
XQ9pb0/0K908Ey1HLQUjVQACMbd68lAt9IwgaeevIHXmuHmYiObmcQoYSr03Jc96/w8Z+lCe/TZf
nVUwmy8QD4OkZo5WsDzMCFqj0+u503g4oScKXAu0rhbkK1hpVDRVih48AQWUwIBXuiBFJRFkurAx
znv1YIOlsrNNwiB31QWXn44r32OT5i8QtRJAVN4+ZZCq7aq5P6MPu2ljvqAAvuK4QS32YNcL3BDn
fYMsGkKj8UECUVV0mVi0U+mqqco+YGV0EZkSEv9zA4EQ3aG81Lh72Y3nv40qjp6rVoed6etRhfj+
44ggye4o+G6NZAWsLbQKVJtcTMkZ8ocZqcuMq18EQVV7x3e3hQ14a7S+DGBwaR8firdmUcBxQ1c8
1YM5RIyXkPjLWnCBA4JvN/VLENC4RnWfhTAPnHB74HQxU5QnsFlhZjxW7d3HMiCocwQ7Ag3pe54F
6Py//xQVlQau2K2pTTE1Mzeq0t8PVHrCkiTfL7ZabdZ/itFtmPTHXLZ5QC1SDdOcpgqxSh3QniHC
r/NACyLAYA5ANQumviufYjkX7CnyzhjbYSmddpFOa+zFhT6/LWYlNqK2jDUsWscVulBDoEyP3ksG
LrV4B7IKlEYhb990bCYcuRe+nSzkYdEfRDDsCt69DVi7vJfkiAvL4KZiM4JVRE41zpIkRqHdKrob
4eGLXvszSIi4VhJHZ4KcYpYqRYXd0KdWGlFLmyZNvDZ7sXmH92RmSMbUFbpaFzxYBG4Mq5xCD1Sf
PjYE9Uz6DsE6RarxvZsaGWBgkfHdALohvRUlIflIASaiMcJF12waUPSOrkfNcKk8xJzvFsoUDGUn
gWol3IIf7sdTEG1cAAa15uqkH1cdo2DaDg6imnKhHA6lhk0RqHBAmhHgVgjJE64jRuijpsrgJh7C
P6SjYsQVyo000oEj8z9wevNWFXxzEKp5tJdfRRurDCnJCcEXckRUV4uVOQAAK1bWk2721Dy4sRQV
7FSR+bMPE1AqUVdYNF6S/P4rzgOP4+HP9zZ71aw+bBIFerqVMU1xW0qxEiWari89pvhAz+uiDEMS
PQtyd7I+7ZCNUZAH5IPybboUrVSF+N/49OBc78ScQ+DidHuish8ZyENSdNmtPPohUPGZuTbuiauq
fX6BXBdIwQRMNqUCiFkKG4c+QTf9WGXQTDOaaznicLUv2ZuCNItBvz+YQM38gKyIcDmgY+/li+EM
iv87deLVn890Wcs2hSOFhZcPAiOzha/gpzsN/Kr6DLeWaeBYmo7p69YsrHbW3lZ/J2/EBnDp0qSE
WnVH1Pwff53K4plD6Kr9BYo9XJLk6AhN73HVdl3zixKdIXa8W8TPm01hrTfvei/cm7hn+6z3htQB
WJBTHYirC/YTnlq8ERNPVBdXd8isoOFLv+87o7U/oShKk3ymEBE6K+vt6hDFQHbCpwGfL4KvgWlr
j6q8yQmp0xYK+JPpIn7o1QxaEN7DuVtaRM5uc/PVhwhHzQH6WWI2JqEip5TEgFGzkiXJOTWiVq2G
dXXNaH5qHXtW0OgPZqdyVTAdR22u1DytV+dNJ7c7xFDwrhEPx+Y/SDBwXGjRFTJPAoYHyx9NJ7UQ
b2/VAEQ15gkDXVt3CXWIt+6n1TfsvfPqJd8ISKK3CHT1KwdoJESeVYu7xOJH5urO/eeGvFRV1Nde
gSwSbxVKNdjPOXTc4A4IEk8YcYXWA1ATBzBLAC2u9ndRNY8vreBpMvLehn8JyPJZw7JKvlsvC3wT
7TPwMqM55XyQYL8HUHn/SHHGxIYoOd2QiLv642S199ImDoVGP8TZWRLOR+pjcBQULCV+kCFNLwgw
F1ooEOkVlp19zP5w/qBixD0C97szgSKf8fu+/FPip9bwGl0u2j+jih78gUbMrIFMTEo+F1pU/k9u
HnC71YuBMTmX7c8TagoIATtBhnDPlrSX7XFvWVgEs4XN13zYK8Y73KADVbOXkS0WmEcQuPJxdPia
u4Y9gDTElG867odjD4K1hwPqh6UTheq9kbiG6rcRy7Rproad8e8J51k8Q0aQh7qrIetsw1OzkU+5
S6FVGgyDeIninj2ky0qSk3bSClQjqimlgbVw8Fk9opGwthEpS7NcYZgLjsb+Qhr4qEWeaTNrJz8M
tthgdQPeeaM0dckShgJOxTiGt2q7b7hKQ3tDfXDyZzkvvmoYrtkuGeq1B9g+RrKQ5qTBYRTg3Odk
X/dM1QHcl86JmEbzCsG/3DmPfOmM3vY4XfJ1VmcpDZxMP3H1OBKUWrNW+Nuzfi0fmLY82nZdR5dD
rH5ndkdl/0OtQLk0Y0dcz3pZVFe9YzXueFqYuPwZQu89RTgqrBA4O+ieIpVg4UXR5cnK/fvj0h7a
cY2nJiazCqZ63kYvita2Wm8e9gmS12ZXVuCWGKzkbTuyrfRUKhrwE58P/x6LQBFRQnOkuCvTibBq
A5YqJVqwi4WoyVP78HZwQin+rjnMFudXmhkJ+rX95LlvMp2tfQmciZtzEdQ3X1+tsFVnH1Sgo+yy
ptv2eBX6Pyisp79Ly+BE3jdVrNjdkMbeNqWlGrsRfPddAD5g5rchNVs9pU05Jpjuq4AV9DS5XULA
473kK7USztgDwD/lgEXyqv30N/xxVBsdjghdLDOz8qW1+iiRcAraJo8tmgokWwkDrwa3At77VzWu
fnHfF0ZfqaxUKEV5vSoPDvItku4bskdVOeiCrynjbvmH68ZyAMSfMaP6GqzF6fEzO5ghs0mxGxGC
sAgzZQaiVnbheFYuHabwyKfjKx0vtAbORO5EeTm1PowMnJy+YtOAos9wLfNPQYvBaaiN90N/6WxL
ICcqkp83zWd8TZlLP6hCrcduPbYQ1pUUKbICbeFp2MLzocWKxG/BDsnKix+ZZNpbPzVliw2hMyyL
1BLljTLS244xyrCHGYxKVpqy5UNXikAt4GTCDvAVcGC0jyPcuXLcU8T4Vng/jPZdDHuOPkHsJf6u
Oye1IN3RqhD8wt+fughGyT0rKD+E82vNf/buBHEqxxRRughUt6rzfrK5PUQar3bq6rJwm5JXuYm0
rqKt/w8mMLvxCwHrLppIV0WAR8Pk6Zv67HmKb1Y980FMJzpG98mfHAzyE/oZZ5MwXnUe3syFpVPL
GoG68b4vJkqoBUpYwZPCSRYpSRbFlGybLfCRqOvqbKhdFzeMK6pwzWIay5RCkAG2TIY617uft8JZ
mNyONcEgj2bbJKelRLAV0VBCQwMfmFTXes+4dTn18M9OIyFZE2cK9QOgXz3w5DGPG9KuUJ9/LV03
e3aYe6iGOafXB5/4+02O+RzRJ/xOSd4R8/x5IeJAQBpjHXL/5QZZNmW/byweLIYZrfwJt33ZmhdW
zpVk8jhMtTiyVyFjD5iIcP5uqkENPxF1lva2gFmZiY/l4UaMcjCutmjW7JnptRSPKqinWC8WdN3d
jW7vpdea39m3PBNVkTWCghDmSBZZFUJL5KTML3P2F9hKiapeE7thoMnigPPLGL3r6Bs8Iuk+aXi2
raoDr5IiCkMOOtLshcPJW6ofWrtjVEDyyF9znRYYPlHPBhqe61AmC/TkkyrKfbQIC+Kwr4US22hE
ip/Ok3l685pKRI8JQsgv8bd1ObsijPhEwKpvuLQU79NO4mpipAgCkeagWrxlso0fhC3y7fKSGXff
afYrx3k4GqEnHdBKAWh3lHPqFbD16I1BfWstCoRqEtimrcLuyeeQlQYvGMBiJ4aQDh4p/X/NCIBk
exZKVmF/3OHddlo0pk/WsrwSrkFHJltv6wd0UAjCSkCOjIiZPUnELR7Ja94zORAvvVf94zqMhu2u
KyokLo1V/eMifVX/O+Cig6vQwjbvt15V7crd9Y7oMr4vnR4wY5JdRTMsaO4h/xmeF2dJ/5gsW93B
BeHRrdvfh4WZRYrmMUUa4KsBwByi7INu/Jsi3ZixU65AZ09wcpOS/yuUmzsr4i6nMJfUXG73K/pA
5CysqygTR2dQfytPWt/nkf9yFz9516zj/ofwh+gykQpEh1IbWw4XwaNMV/JQp8cHm3DE8v/+Guh6
1Mh7BDukFvoBqsgYC9l0oS+teOaWaLstG2S8FCYFpSSiYU3nEGRWxhGcY7qwYrl3W3QVt2J4n+06
kGaTzK40tlNCz8YKnuw4z5CAvWO5U5LLaCm1BC9bwqSbCy6iYxa5AwV/KYOpCqxWQrN7e/QjJuoz
ZnFjswU56vWLhI8CHIBSH8O7lwvaCYJtx0Lys1JCMCA4JU6fmGpd/i/mYMj7ZXE/cpzN6Y38sFnM
XOOyJBCWYMkI2VP4iz1xbvUXzv97vwpQOb0vSw1jEoPuSrxLHhapen2fSQGXfdD+7TkPxGPVAIvC
0sH3p2G8cLrVPXPVnSxiGJ6JxsXlCsPGN3YeskMJ3Da9fJVN8Hmoc9n0nHYO9fB0U6xY/sjmru62
Z0GN9a/KDwBOtNA+CZ5U1LmtAt78lTxHz2qJt9oX9mQyZjELirptP1icVKVyt97XfT/rPvfTJsdA
4hkFZEMeLSUYr0pT/Wcrbz4x9/eh8xQhYr+mpsfasZsP68po0Y8h2QdME5WiAw42iMykodIEuQtz
wS51olpj0Pe58+Wks0CFHz7zbGwZ6RD7HDM7Dv8Gb/K0kwklJtTpyFgtc6zTW90bu/64yUYFvLkq
jFqXjAzU8fwN2PZBv0orMZApiBcOkgfabzTo02JnT+CkPSCsPtF5yKWl8UyeiNtxzPtxqnUoJBxE
Ae0LWkOrFB8s9XS5yS+31AK4U0dvqlz3R7lHcLey/8Y7SX1mhUoYt+4QFfQCyhNbGy2pcmOByGdP
lyIotMj4LxjiFl4BmLNcuX45XTzTLDWgWGrKvk2EwgicGIltLOKDd2BRF69yc4C1VdGrjypopByp
eDDuc/mVItbe4juxBSIH4do2e9ttgRcz3GN+QukkrkiPcuqxUFDI1n+yppTbUE+yQkESq/R8AbWK
dkHhfi0t6cQot9xTUeWLqIOTLm/E2k/icFELPEy4GJaGD7HgUz2DcfaD/Ot0Fk/OomQUeH5x3+0i
g5Px/kNDqchTxuTi/cF1qXaVKvNVFtaInDtfPQNxb5qGSXKSkDuQDyX9U3brjb0Q7j2ic6/oRpzg
9/3KWEx3qUE46iz29BMvUimEP/ADdKIwCRDoAZ64L8HEGZc1X3JLWWOauCit9jB9b2QDE9eMlgNB
d6fSWqB7BKQyXQH3G0ZSKgMeO3Znf4jVudw9sB669TnaNvzodlJE4QMDD83f8J4lOPq45pHSeN4n
QBzgoa2hRFy5BPqZklKUwxYEoN1fT6dzv0llMW6mr2YY0fUgNCkPpypf0hcepxd/pb1H0fA3RSM4
jLZi5RV7kfnrGry7eU3lta/H0JwbsQPC6P9cyaSpg/uE6TCCyI2z80zeRzYEl4xNTLxFKxmK6a7R
ftfVDODVD41Cl/pxGYy9IT+eYh2yoWAGY0EK2K1tgBl5PuP8XJtGKnuAliHC+yWfu0O2uMgDr2l8
p2lyBu31MG4xlSWGkTS/ONwAiramYqxAys8Dk/yOLuUnCTPLCVOx8EJoscwRP4ZvDkfCd+YL6N5+
GDG99xsb+SeNqKv77lUBgWUEsS0CTpyVFKVae1MJriWvldlL/TxmPPDoHBifwCzdFOIDN8iQBM5z
e8ZeWZVx9DlIHai1YmA5RabX6J3RNRkvgFId5EDZ9kQ3EO/ooylil8xgr1eL5LA50pJHaCeR5isM
eqCto2+EnygfwpIdwqOmQUN8nA0AVM0xv8tw9+BIAhSu2qlLSQcY9c/CUT6XhgEBUejF1EfB/ZC+
Qfvf2bxQ81/CryeuAtXqhSsTWs6bJY9MquiukFYlwFJ7/5kue62CckZL/XDxxfvbMAhrdbcZ5XE6
R02JRYHpDTQO5pR0R5OAit7vfLLRBEET5IRD86NIvFZC3ewRGIND/juvtXLLUxq4rjaRFL2ge5jz
exQZbsZb1stWy6VnwoKPxIRE47KHmiSVnmcIuTv/aZZZnd32brA8SIt8K4Lm1cctliS90hj6nulV
B2KnbQhKHWBtS2d0MMXG7tUkheSdSaHbXBXORbfRjkDbwEjysq4gIvsbTHKBoA1AoqqiUMSBcDxh
42RCB94xhDrqJ8TP+aFcjVGd8DyBtXAsyxcKSLSRh8VSAlZINx+EBtZL3CtpQVeNWI96efoXpoAo
SkvBdiqdpvjiaH6A2hDOu7Pptwk8bU7UmerujLR0hGc1jZOsEGbTu5J2NgSGDHU3p1ZGL8ErSdZF
UEtbYaDoPiXqVaMPSBl3tNxnyuaUM67UK+bxlh0qNl2W4DKnxTrdw14WuzJ/e3TLnORyJJ6hMbsD
clxVjXrKbu6DMgNq+wd4YZxRUxnmOyJgT6smhu2glg98iEFT8g5pNmiYIW616vmi1npRtwDiDegC
zlyx1cSx5vMDS8UNTWMwkQqC+7U5GIOESKoPjh4+JK2r/9i2ZyRZ6RLdUz8Zv4oFfVTZdLc0mmSg
cIErQ0jaBuIf7EDa59WqA7RpplBIAzf7ica48grK8I1U9vAlxO4iedmKiAlAy94ZKMi9vZP8Vuxo
ZS7w4QM9j1HG604u23XVYuUuB5PC+hrAjl97ce5EQRDPIEUuEdyAW5bdiOqUJkjXPV7/nNxvMO8l
8qVwZd/njidTTlZwTneDqXdFZON4bHpA2Goz1fiwZV2Cv/NyqWF6Gamo+9KdXJXU3i0yHWpfKrMU
RXPzDf9wDP9IOO9+ipy8FWhyakjeec+0LBmCCQgg6/VAkR9HGSVGjU/I4qelMNaziphiEvN5fWEr
Z2dylGBWtMPJeWWUzX9GKPEHwMdB+7lhrrMzxnnQNIFGxO+4JLdetWjCXJ1HxQF0nuTtIYNCn/IT
WHubMC34Nzr05YzABC0VthOY2xSuXDzKFSZ2IUNFVr03ZIL3jIdFJ8CK+UcVbZaIlMkX2TP5WkA0
og+slSTfbbuEAvHYnSIb/NnPp/DZaTpUhcOhSM/6Bqh3BCuAaSMOFHCjWu9Tw2FltouNh0MDspJK
hQJ3FA6dEyJH8t5qXA8Vv5tn9iwbJSdjekLdrLfQI3TPntyc2w+NHYW3sVk5WPPyZK/cDuA1v5Eq
zY5KXG5MBIBA7ZIicEJZ1QXODUIdJc3MoOuNq81OLN1sR0qZEeaiive0139alMUTM8jgl5hCTK4o
eRwjVRJcI6hlfNDvUsshRbzass5TOPbZX25uTVil1ZSifQwAatePZKMJAYHqTfY+zadzlofS4AnG
DCy9kNcfiqNlDxvu8RHf6Slin2s3W3VXfgrckxzMXyauYt7OLFs2pNt7W6lAFy37JsXWozeMAkwJ
fXVmQuD+yfkayR1yCSI8RJOEBsPPM8Go1E1AHlUVEhtAFtSHi8nVSfLzvG7kGv9VyMe5GtUmsEWU
BrcHO70x2GTIbKnKf9h7wiyQbqlEQnxCz6PI/D8eSb0fCJOUkplpI0Bwuf+oomnI4Ti7Fn6Fa0d/
5YKPkMJcnCinvto6xPbXsC/YihCb86Loep5zVOMw1ik0uTCHaZLkkqkt9QgfKtfMzEzVEsoW8tu0
0BbzxYI4/tD9pyfivfpG9RKhjmu6nIKqp6Klq3rkxryhToO7Ef1TtO+XeG0F3wmTxsy95tQqtIod
rivZURMlDX8ei7m5ELTSjDpVk0YgSSwK4HAIZtzVOYqtdmz74OmLGSlSkN+UjY6HeoJuW4jmC9XC
utkZlmLvi4mwKndeJw0Txvso98FhBKA4BsHVw0U6cxcUE2KGV5le5LC/hWqp0BaLH9Sv/TI9lJp+
beSHpA/qjyhdwzhxYa/9x9I71d0M9j61xoz9O2Kfqj9Gn+n++zXXJrXuAIkX/0ZafTcwgPuIVtXK
HJC3AYQxRSNtSExjMBvwddCiD4M6oolw0ypltdGzPseKaVjqZtzXTw74dRtX80+SA1XA/SULBK0C
LNV8dpO5s0hYZ/EZL+MHJozw7CCfv+dOsvq0U47gnIoOM4L0ggfDBBXj2IhBn2QYo+FiDRQF0lcS
BIprG2r318aRYp621g0VBXGtyk08Px6Y3l8WY0uINo9j7f6+W7tqzlH7U/4onOFlKeAr9MqyT3gM
NzziswBI6DVCjYiuk9KfAWbl+UXrk7vj/Djf+Q5KBG6G+iCsMk2SPgFqDHtGZLlRIdjQxAtBvvF/
VuYn8V+uL/plQDc18r94nnOhOICr6qa9qhzOto5dcJiZxoCpKMFEdo3mcATWjj4mYjtJlqp5subZ
o8uSWcfMpcI8zhzDji+d/yBsYD/6qkYi+9Qci47f0tI41S5QIA9LHxiI83vpac3/x80W8SYjhqsa
RjogvJXPzdcXFe4SKcqKJ2c04uo7jEoKZfzGRs+aF2E+/kjYKIG3VuKtOF5KvyML59SkQUsOKI1C
tGG8nvoZaP4RxozwogM1kDvJLpB5hlYhxPLlujE/Y4sD9geivVs1OuVyCOnRpR/UZZ5/2V7g/+tT
aYH4g7lUlnll42ra4g34/qqzPMLtnbWVBIuK8jMfjhziBDp1q11WAh5wegGwt2/BH4+/mq4VcrAY
VPeTB1K2O9dmxj+LpootaIcYTORL5OfPuefqz55QkoWPPG0xXOeVFdg1e4ROnlmLnNU9vD29nHU5
hTNkGktTG0E+lFr+Hv55qHwgugTr634YtVGbQKPWC/GBZl8787mzYvWx9JRYFAwVz44GTifsiEms
uRwYanm8IUqG6b8sSWQ7KxkvZ8uBp0v9ufx6OWEIts95KGmedDcw4ujKez3bkBAYqAMNogqiHS2m
0wCGaC6LNrlzXnyVSU/Z3gtdEqiplMcxVljO+d2uoBG9g2Jhp4bte/dDyy4ZHnnqOdHdA/PjoLYN
pJph8nj+M9dOaQ78mMi0CpxXdUGlwctpljT3hKHDaN69+2muLBL7ktoFXLsr3hLL6DnsN0IW4kbQ
bHrP4h70DH0iHb89UFL/R3VkYOgGEXBSYjckdnM72OmV+k21Xx2i/EIXPhngdem710uAHZLJOICJ
zYe/lywEzA7jGUKiEd4hsflaMkht/+KSFd7cGcMX8PFCL6X8bCgZC4fMgyXQmCU9LR+9FNgWHaKj
XlobG2knG3r+qjSSqRbq6jAi5/KVHIr1kR3i3yCIzMfAQJsjVwUNyQQ6Jkqrzjn6nleyjwg9CXOS
Lf/notUYhqnLraZNznIwqnwVFYpiex4CNonKoybGCvuTDXrE+XYRWZ0NTEuvcNtJym1QZY01paNm
Dy+in8GuSXNJop+QVhXTIDFf5G6aHLpQ0LPG8E6LubIfOwKp6EnX4Z9fuc7OmbQ3edlYtUoXYF85
YRyYaVwkDH8yG8zgfZxb1A3nYIJiVmqZps4V0p+LRDFN753XW81MDNWZpteRfuqWVtIvGkAOdr4K
xDG6ZjPhLXINth4p1s6M5mZe6eu0F41eMubglQJxWwg9LFMcFoUZJQDSQmxWR+HJymsjKpd+5ZGu
jUAVwAk3QLyI4Ewslk+RqaJL6PdQef+jNF5guBVVHtFNk6+LrX7tGlfnqtF+s9pU/CCNhCefGcRn
9D/FjMdE4csnODLfo2juJdanSENYGpgnkEKqXdJk47mllqN62yf8lj9NSAAJo2nADgRKVd1H6fkl
HZPhnBNufXqpvs1EhmUXUOThwtUqidBs3j1Jtnx9vRtxmqlp46MytY+HiWBL0CJCaLnn+RuiFjLS
KBGPtoEsWPeg9hOzFSVennBIISmciRz2r6Stgu/Lo6Q8w2+HG2hqIH9B8XTLBl/GTU2khK8S1u3e
bzYbhmEXPSlwYYwQjvvyYmuvyEfKP8Hu/GXsTuXkDH8F/gBOU4IsSpX5ZrRhKtxKe7cN4fWYFCWR
EfARrAFKLfUFDEzmO1V3igQPWLcTOniCXSjDjvcUd4r7gJZ2H6kHO7P3AeL5lifeSgqdStaVjUk9
bGhrtk6qCJRlDi6Vjtn43gIUq+ZWY6X96zzovc5unTl773vYLYb8PBYCmnLr/44Blp9WPIMn958B
PjAF/IRA0k0l3ycM3L3BLdVwKP0eUuW1M6FLxDdfPNoZUCBe8r2acnnzYT9rpXdLIw8AFy9K0bR+
FAZOfaR10oVNsQNAciARGZLcjWQoCg5riDhYV29qc8Lpes1qPnHbleGhaMjgdCXNE1zVs2GqToQv
3ER64fzhvQm6lG/9WT8YZyqyt8wDghbXuo2e+CiVLsUNS9UF3yiJu6KnbJWxtY4w813K2ogaXSZW
LZWzQzWoDSk5rMnWkGBleaiYgZFzeajBt2//PP+GoDhWn84plaOZy/a/rOYXfCk5qvDmYcdVD62d
xOVXzDafz2+upZJ3gw4tdJtDVU/Cm68HG8fKR1lwG5T7F3fOOgX1U2qeqpDC7n89kYPTexUXLaNK
isMM/q8+yXc/qfUojwqqi3znhl96YyDTO402ms3O/YMBdIa5TsgW40pA3aAhf+3biAuWh3SGQwb8
N56LJXkluCy9UW4PHrQYVaf1SfV+7h+V7HyTfBjM8A+NCXLjw05nY3KVNNBqfR1iHdAwJPmLE0eZ
S5drm7jQl6/8MU9+dkA2QmPMbcWxgVg/vtPdLIhrUPyOUDoKHhmxIs3TvFJpEKWNLKBrAVFvAm7f
uVbJK37mtMycjHNs0WJH1iyeTKWvbvlUEnNldXADNTFD1nI6mL2XpMw3C2dbNow+MTZSi2Y2b9Ft
L/udQQKE7L5Uete7Hv/5YP9x9KjJjZeFuEdRVI1XUJhAS76FDMOqKRQiPbMpckEU8tKP9yeLfaWH
YL2Vk1H+ECIx/yioqgMQscElhls7vl+2d07B0520EUaUojyV8RHqkE8u5TLAj3USEX8p3tFQT1uV
zcs2GFyaF1ObZ8kx/dizOJRyKKjeIbGLLQbBM0xZDy/q8lXAwNxja89PLCGZrDlR9v3t42dBDmO0
I1VdEXRZnccCt7B90gt91YPDLDITSYyB5uxTdI21VyAe9XLjw7xzVvj5QscWDMEdVIvf0qpQjX1/
AYpDYa0LJMY5JNHLmMzFoPQ2dUo8Zbzpy3uYIOY///RY+E3LrCRsJtM3FxRbZwNztcITQg3ExGol
WtLTKatYg0YXoy+u+UzyngFYB5JqlHa8QFqxDtvJES/HTHZQ+lAU3MOzM+UPP5EnKNdX74QhDL/o
lCmeRn2wholc9FptML4t/gyYcv+4jHvA5gnQeMslH8kVDokd0dIzcDQzH+yXkvn0CF9qTGbloeOn
SsZKHZDZ+0wADttKy/Y3ibpCtR0YqMqcrZbdABKZSWqkUq6NuBnQEP+LIH7g9Wdl/fA1dVesA/tK
Q3RRmF6wvXGvFX7EIT6Y3hlFX5svoo0czOSfpMnBax3kHIIsJd1gjEswvpzvC00cDE4vH8Q6IC0W
TBt8M9CdRAL147ZJS/3PbITXvES2IFdEkvO4wpJw1kwIPFdzO0LTLTvvfcY/lLK4wQEDRgy5ISAv
0SyyHpVd5DyhLtjcnzVnEmFU+r7f+ZK0FVmlzDPTeJz4IJRIZa3cJEttB9I4cqX41IorrEuNCKfd
J1E2je9spFC1qxZy3PdXNaeGVyEZbXlpGt+WqwR8HrJxIt6J3aqL03QfxIiAh5HDc6uLOhG1u9MW
NO1QIt6p5Qo8O6JtUwv6ZaUgDmnz8AAuqNPW9XfrQM5FuurFpF4OoamTgKOeNeb2EUI3Chr1zlDf
hUJR3V8Tbqeb+e/HJDh+JJhVgCKR2Y9fYSOudRu8zjuYZX5L4E4iBZahfJZr7Ol6bImbJz1WB0m6
bOiXEUYFA0/9ILghBctM8IQ+gCjDpIaOKW1UnEzKwW6ZXEYb5dCC72vo0TnkcIEjwShI59ECM71C
tfg/fwbuO9u54KilpFnT7Y0dLcpePUn2ss1whfAuFJokQPyuFl6TXmZnxots6v+hEWtgNVFgT+5B
8AOsGCQSYdD4GXherIecDIs7Tb5RAAAVT4DyghMm/drjHzQ+sIzsmqPGP5Iw1UjQeH+0ruBJ+JDa
3KkbLfL7eDZ9E+nqy6TV2f8lOSfxYSEfGDr01/Y03MgwCEQD8uQEEATY3jjp8UW5b82txS8X9DcK
9jovvBnSZs5wJ+ezJFQnu7XNi+aWC/pycCrq2TSCfo5b3Ea6pigHA8WI3Lnt12AhwhsD44z5xkvt
R0pmK9U2J5rx+d3yocP6/velkNPU/Jq+cizl9U5pxE/xfZgCuT34n70nuguVQr7MKnkwdDrzLOBk
eTKk1u59/hvqdjB8OCAZVEUVjsDs+3LLv4qjti4TiM2kRhdkmBEmfIDZ5Y2HZQzBj41hVPZacR2U
7cmQ+68j6vM/T1379Vp2l3ks2Q+bEpMrEMfFas3fdPliXAg5dlH82qfpMKnFXsd8+16r8Tu3ce9e
8YF3/aAhLRZvY6HEJpl3AVa8rpzP+3Rk5s3Uoh2Z0EPTj4T3ER+3yNVQgMar3ygN1O+0oh+8t5p0
XnPMTcjWThjDnxYfqfqzY+r5+aos9ErJUHVqGXyRQEKFRiFnc/KZ6eLeoahVxUqZHnD82ajQBqZs
3Mgznzuoa3qGTDzJVY2ESrBNBc/wM56z6eSmKA5oanyRI3jefH4S05/JCT9579DAn2P2+FwwWKbR
o0fYv1Iq44LfiSGBtnLHKISmDOIqAhYd7FhqkoOf9Ylkkjb6kmLJ43gFw58SBsMvKjf3sifjBiRs
Cqyh9cJS85JiIJLjrjPE/N4TtNgtr7ULtXpIDC4lcjdZmMAGhYZkFGUT8JHf7Gp6OwOcnYQirh1E
CaBJ0aIQDZ7DMWpNR30xgYxWEr4lU7+edIGMhofMeYVs8oUlg5EY1uSFsZESKO0TyQaSErngQ+Wg
dWT5DcP4RH1E86FBRlGWtR/R8l/J+R4kqgwvJCrKl7bBAmpAL0nekD1K+8tf2E11vX9FZPhf6ZvJ
vY9ToLTzT/yGzT+VpAMqgiziIXe1iFbEJA/nZ+gxELgq+vH68e5jV+vZts2pt3cKHiJn6TuV5E9K
byIRJFcZtNI/xi+jylWsfBZ5UIOLCEgACe/vM2AO9goYqpcsNkc4JVl8MqpL6EHtIJmcRGTvYmMO
XE8ARS8t/owSDZzfOjbiY87Q63tsUgFoCc0hOHj7WIQdbYhNs5WI1wP/nmBnbdbyUDzkfIqtTU7c
YFLQeOr8+nhLJ0fOS1PH34gG6ejj7SmQI+NhEYg/nRIW3gd8pXlcJ/MGk298Cdxz37OrLEsfvOx5
2mXiRsn4bUORvkeRPdKU32MfYEPjAngcYi7tB4vWaAUS4uYmrhVIdx6UdfikGxjY51F3xiGhYGwn
hxy+7i3ryIaA8PkRchDxMs/iZ0Ko2K6l6pi6W6FpD1iY2UvdJbsmj9Io0zvlocoY5tpHRnDAX5xF
naiAAyi/A4ZDMSAG9KW+PEWLiPgkVUdLHmhwZD1Yc2i2cDylCaNRiyZA4r/ZTbHeIGOIbWSpPRoC
XWyiiUVbjLf5WjrI1q10wOPYmxi8m/IMhX1+nnyADmSQ3hoiNtsN8tX827iDg9/WxhGy9mEk2ykU
UB643O2Ego1BfymVr+EZl+ado8RLwSUqKrNoTOgP946kR832s9QuhbC+nQePEwx4zbTyfiFVoKr/
b9R61QVtWDPub3Xg3xB+bTrd91BQ+JME1vwwi/7hehrfmvN2oKNcxFeDKgF7Hsit7DgAQXNtqkbY
U3gq5Fj1IX2NQpwXeE3sIrvkL5AkeDhbdrZOGu5kmETC02EAhYdD1zGRd44Z7SRX1j2qwRuTAKd+
lHkTJY5WKJClc1MasEDLi3mXavHLzlKPP8QMf9t+tj/SmeU0EieBmsKvDa2+QK3xsQFfEzeXnLT9
haMDAORG4nHgx/mk7GxjtH8nioPZBUkgHj+sw/I/LuvUQB0a17YEUvu0IcvAEwfkaCKRBQGNxSgo
Pc0ATI3jkF4/pgoSmLUAfU1l9Mu1nHI6FEEGsiblif5MX8i++CLrCkiX8bQxGIa1fzZo6E75y/CF
qQyH0qBqHuz4Y5RZ5unxcSqbmHQkmaAMx97Yxic09X6HBF1IzuLn3dXMf6qZ9ce2Io7bOdVAXxVG
UDjr/SliogHn0aJ64Ku1rXKovPuVvNmLQniWV7FrW+2Rb6mDVtcjJCTbLvUdTsJLTpiih/+dcPmS
lvrXn7VtvJHY9hynuHcU6SgK6Wcwvs3O2zRzTLC1R7WfCW4hO8sTRmP8QZUSVmTjM7R9dMgv1QjF
eSlRr8mqVSv+83+aj5k8GG2BCyL01UxcmGipPLPcAVKR4kFJb8TjQgNDpeAkuAnqnxow1IOuQDRl
ZVUkruF1pG0RJUo6O4Fll3xk9w9jwKg1E3Zso9nFWxQ2PtWqk09LH5Guu+UVjVRGZI/IVyytt/YO
2pj0p8DIPZmrOg8jtIBh3m2szjJsl27SRDAQDejLGpKDIUQ9i8P95qV6hNLcCr/1td2NBoUP5hC7
KErAHdpnqyV/DJ/IYIwKaUTg9KuB+B6FsBIWjse3IZ5zxJACYCCS/dH/v5XoZ2xxGTfcHrPiRVcn
d12SD8+WOew8v/qzw3DLwLiFgDK8Sr85drdRjRzWDDp+KFEO5cEpO/Cf362moc6zMRSsHE7hU0hl
m+VT8Gzd+Y9SsW4fIhLmNa7+djoeGX24JuYrMnAri/UVLIV4txuXJh9cpJk7e5XG2xX51mfKS02x
jnbFUD8e0FinG/Br8429tbcOvOr+YtcGuuFIdYueKdNCU/j51uGqA3gA4aZl9LCxH8zKWt22FFeG
pbcYfqBVuhPWGUV4YwFz6IFdWQ2s4rV9Zn66WJm4vO/thEyrHuX2Ta8t3YPsI7I0Zsf42GpL02Hz
m3VV+/SDbbpcQY7I4tnUTPR81I+iCOFmrvRD3rAMKz2l9oanaPzKVsM6FWflBYvTROOFW7X5G+St
x3WDhqQdYmiF0xYw9oHmxgOM/bOsnroxiZGGy0KZp8KViH0D68DzmBt4c9ipxsnsiRd9Frt4KoTt
wTi1wL6cbGPwZ1nF0xAn8HYiwmVX4NPnd6GfYBNunYcKgkxUWJqlDq1aiQ1V2cbymFX3t8xxPM4k
wSmlMD2rReO+ymwglIPgqoDTQBXW5Hud3/CInbmVUInBW8ObiiGLbFwPS/wnIpi1p4rtebTYrBma
gVmvvV0oG4Ave9rKNK1tWzo+9uB5d06QqqxKYUjquU6q36DduZCY9iFooHRyVta9LLj2ZIVsID9w
DxSyyoQUgvyArpKKqgBn1zei1Dd44CaFpgnt0h8ElSSNLYE3TxJU07lHO7snoU3Zjcu96eXkUAFU
wBkDiETMc18oR/G4SSWV6TZoOaD0NTpGI+OjXt16siUAbrI709os5VGt6QX+n0gsbXRYuhupoyrb
zXkVviOv4tMHSpVilX5m4iYzgXNaWQIFWXFuYUYzqCAy7GwYhwZVylTg2xpuZxd11COnK6Pmw/aF
fjezDMncDUbkXqKwDO2RvDToOjHV/jDhqBg26hQVrtSYBmMK5yuZ8wDO4U7u0noFPk43StMv3kSD
XDKRzE1I34hvc//80wTtPadVZzImZiykFob88Eyy6/Rhe1pYPxdw+m8bsNPHXlD0s5VMtsgM1OSU
/ndCDY0m/5NmAsrV0ZrB1ctXOw+hMADrIk58ENrzj43cOTPHuLibdbqsXAU2I03maus3As0uswoQ
1QkLMzUEu7UrPnfYZZvbqAMn73kVqyAP6mz8GnU5Ua6kGtL4024DVovKwzeYnnZWP7Wfm09+uWPE
VebmySOZbbF0Z9xjTyZu0Tv9bNIUX7h/J1yLwsWaN8kUpMzjoZbGobPBbObZZySLZezsQSzocF+T
CfayVAiwSGwEsWkZ6p2xLdPEEEzB5kMqcyxf7exlk22Dp2ksa4x+CaXgi135OP0cN06+WPM20+Xv
1nm3+7J9MycERn8IQE7gSQOUE59RxzTPNK6X7cy8pHYz7tpgf2biP7W9L8M8GVLDSIhFxyIRy6PI
/Hm3gQlgfMjCt5UTAwAm5B0vIhsSSC+IkfFBijLE+FDp5Px/LuyQJ7li3klS+kpgvK/+TP8Wdc/F
4Gf4r18axYaABwSE0gJiNChj+AFjEl1zfGbhDiUKRZlLFm1MGrhD0S/CROvZAr5MOFu2Z1DiKfsB
H5xBNghz8+Rty+swL/MYGr162FDWBYK3jeL+7/bwYI+Ev5OInClikakA7kLMHokIwge2fW4UmE44
otskafK4xSKJ0xUzgzoVhi18hKU+f4xnToXU2HoIezGm/bITyjkNxgA6AYNAU+1eTsyJLZzWrr04
GkTrrEsWXZT6l57YPaNaIPF8unBqBlb0IwciR4qOLAcH6hsmoj2GiqDuSVO8W4WJuviwErLkM2+x
6qlLHAk42SOMRWbZ1KJkbEd+tci2chRMyW7CpCDohDKkgfAkAJGq7YdRW+rlkg2f7AfrinnII8Q1
tRv1hrUAU8ryvW4r0v6XxK2hx7vjX0PqeSTRbTnPGOmaH4I7jsrB5UOlOXTqFpKbB4YhhvDwFbp0
c1wiPDxRHbUtmCHSUM4oBSj21omknqlPCNJbWSb0oVsaYUTsmJkPR+185S1kyfi/3/agX4hI2tAc
FgImTHwPnJQkYvmjGt3hr1SbYxgH4K9J+F/MbFbqV0S/L5xAPquXqscJD+v9AL44moQr/obfNXBw
FZahrz1V0ezoycFI08kWEoP2SiX1yLqv2zNv2zm26Z4C3gYUkGLPiMNeQwihGpXS+xBi6GtpUoCi
rzPC25QGdiC7E+xNCCMfGQyMVsDlw2VdngrJ2605Fp0dfi3wF/TnSu4hQ4Wv1FAJKQQ9KaKN4vB8
YapSmS/QJkrJ2wlAoz5FWphWDAQKjv1Ox/llyOy11d7X2QIJUQgnY8nX/NOxZQlMTzB5KpD8quop
qX+N4AwPKlwBt6GXW0k/CfslaLCQ03yPkxGMdXnG6xxgr8/bFXGEwD+T0onmSZ6omMi1E1042HLW
Hnf/9aAW04ztH/Rbm8fopjkgbXhp87rP0AY5eWHKBX0mZJpwROlzCfplS4GUCgZMJgUSRtmR+4vU
9EGxa0vAnUER3VfSWBJZAA5nUMuvPpKamEWIRILAR1WDXbSfH9Jl49sL+VU09nh+6CqEQ7R5+mRg
Zdh6DFbWAHKNdlgQlBTX0Zfc/bXhsiunI06zUQeS3wzBWN+53fPbwGO9ZM5Ut4HK6rM7D+HOVg0Q
2u6w+bv+afXL11DTPzE5zWrDV8CtBDVklc+iG1fZT6FSv/g9gSmjEdWw33bpj+8bWScfcDpzx7X8
vFrNEpSnIGOH/8iG8R4KdMIUFIy9Mk1eAjbJnG6/wbuuqNFqtCgaT+p7170RuqITsJEenXpdrtKM
Z6XjyVcKx9pfIgKH+MZkh5y8mzBAvBee+sEnbkXuRjTaY0zjtAc8PShlOQhbxKzb0jjIJy6Sl+TX
2AdkrbRcFb3kco9Cq4ZjPqrBwHaBnkkUwL3fPp4iV8X67x30KX++nsQ1MhFvMTRS+ZZBUablVe0V
GR34dhYpn9QKUV/7dXKWdJ4wBWYT7tN9zwcjbAX7ZTbqTV62Ju8VFP+KobB8WPwjbp+byUeF1E9z
MRcDHoYn0TB9XY+oWPVm0aWEuulgCUkhj4dQ13QDIYltdYDt4RKw0bBmrH+HWAkwk64T/vu64dNL
YvdF9/IopH4xa5DCUWvhfWENMscm6iY5kEnPXPCz7olMZbkfS+5u5db99h7TbNy9PLtw1/PfqCIh
i5t86F0M1U0l9gSrCsvAzIN0tQSIKSDzcCRopQ0jlPyvg5z+P5gF7+bn+u79y5TIK9edX5O+nI4t
pa4l3HqLRXyxEEP7BScbTRV2n0jOyW+jQ9uHuePr/1Eez1dJqD9e0bBdaGE5tQyGTPk2ybG77HWW
0cQOfZfmhZYesynZF0+6hv7RPtBs8c7RQfHCnwvVYxYcIcopzQWHyffQoO2sn1K2r3X9my/AiRZT
hR7plohlY8moYkYXcKYXaKg7hDDYaoA8VDbrgEuQCjEzvl69oQVqoGE8UAxsAGiflCb5tYlvHUtS
0e360EzKdatlHiBfRlj2D1QRtwIyt9jDwzRmD2aUP3XXVrAWi32l8hQxXzaJ2LLE2uTxVhNcCmaN
ntbQDXn1eliBOEhr9jQ0DQrJA/3OAWid8mqlOC/blcGlfQ1iGxJrmjtNrdP5NYBqVFTdjjM6L4dV
VOw3KxhnQoZxKaifI/kOhQ0Tel0/FRyyiIKg5LFRhom/fl2n4Dksd6rG6S9jatCwVRg2O8poMKJv
3hHC5fRs+8ZT+5xZlqdMmZi8Vg6pUEatBq63tnwhFhXSCWHwJvKGID1FKJL0lgSbrmMxVx4nXxjS
Hzg+jB+3R89P8Q1TTvvF8KPlI2MPWZRKwGpBydsYRvtaSpCLEnFKTKdxtw2aoeyEAwL93q1xGx4e
S7JJDKboDTwQMLZym7I9MKU/ysKinvC3brwigMnqwfUbghfMffO6JxehdCzGgaZxDbT6MeG0JFyz
KY6xV1I3aMydZdEC9j1SDbs1epmd9JcAGN6a8JT6v9IGk3s04b6ovsynAX7cPDtAJxtv7nh6+E8j
VyUFrtOCBXVofTyCCHvwqP1C+UwuiGHzgFrue+9EGsVWiJzz7mDGB/BopcOylkabth7GtF4CBQfC
PrMeZ2vaCWfYyq+p1219dyd1aisEL+jHLQRVZaIUpvKdQh+ggN4pyxhfkP83th+YO5u8BoRsDlEj
J7MfPBz0Ol/kRgeiEo5pRJlBH28k9oZu1G3PaKaf351sogcJCk/aROiYfBvVrFa2jwNKlBtj5aVm
vGXBgDhgkq6Ing5tfD3ICdQ8qWz08kwFeauUFGQQlwopKfFynqsVq5LpfCvSiDpx60aiKCPJs9U/
DpZlqv5SHmpuYqYhy5lRmJTH023lkcWNcPSfuP1vXKlGg7Ffko1hVT/5/DrFHYSpEJeZnrHcKWpm
B5rqsSTMk0yyH9eOTIome32rA+YZ00tRX+Dna2MelrBWE7NsV0CuUar3JyJ9reryMWFYRxxXqjzK
4Cfd83qqdMHgcuHt+9xmHpgH3nUCKmyzuOLzRTAtX6RAXx/BqAJhoMRZldhKeBl8Iunkj7eCIjdB
S5Ft2ah/l0mm32ldhCmHV//w9x23homqO/JlT9CxcRH6eXipHvrI3ZmFpOJ75F4q3XbIKWQcDrf2
eiItd6CAy49Xh8MLPS7XqOy5oykzSzEzoiSViynZ0MQCdu31ygRS7NF82qeL4qrC6riP0gTRgL9w
vLZWjwp7MuVZW6gOkgdrm1GKOeQKLWY+pSj5sSVa7YQoRk4Iq3/Fir1LWCHSt2u7Sn+VvYoNbkvP
ArsfC/1y7oQ/2+jlmbOAfHKWSWOGLAd2baGEw+lobviTpA1uaa4hfggfIyWF6YI/oMDEoqBQhhm9
m7dHQAFaCg9B56wLVkkeEzABJWsJq2dQ/sbEo3nucJSOmrpKElFjdPA86cChbskT4dKOLYN1EUzx
So6XE5hSt5dR/qtxPTumvFlmBgDOCMYqzLcYPv2DN6i5MXRDigfNfinPLGogYHQNyMjtSJdHrq/a
ZQlyO8OI3rePg6bgHXIv3oHZyt3SYo7O5epIOzdzEPj4Vp1znw82xytQ91bTaDyDio8cM33LaHB2
kZncE10q81xxJYdY3dzpO9dWyuzbq79Sca8p5+NZ0Ojpw0GE3R5I6ljHLs2xY5+pSTLzt8guURcD
rIDY+jyMgG6NngtR05vpibM4ZHpzYyvXrmQcLlc+J6ejr1aSp3XrXUbdksYWfO9KYM2zRvjhZ/Ui
Me42Jm7AdD1c9TWBpn3k0K9BUer8rXgz5FXWDfiVAUQ1PsEqvTqNSR8EQa4jPU/XePVkWazCODnb
qzzho5mGxi76IbL6nWTsvxN5xxQ+/QFQa+mtshOMs0ZCwe43aIKY8Oa75w6XvZxIX1VnFEPZYJuy
Z/UY+iebh9pt9KZjsyphDwfSfmdisOYgk0AfidZsB0pfGj7Fo+FyYWNlfKKt4lV3vQkuEBFBLDYd
LB7CxkpSZnqJ1zHxZWkLzWlSlPvZbgqZNZ5j6Vb9WvXAWP4gomCo5xIODlzSKhavLYxC6Exa2Twh
GYDUkQ6wpcFPzIbrrZS2tJI6+J8CBWbAKCga8GZHi9sfg2DMCr8B+TfbPKgjg0a3S9uqikU6Ng6W
FDd+CNPLG1/gdHtNZcLmHXyu1wPEjbxb50SnNabke6zXMUcvOdjnDNCf5tI+itVAmT4YLwEWaEky
TFk2x+A8xgX/lxSakA6h5yTffwF3J98KNuLqJT39ryKUyivXzq+8JU+vpy/7wE69lH0dcUAnJq8o
4TgaC5kFflm5Urzxmp8WqHCvl+rbxKyuo6xEtMM6Dxi/0NfAg2hJMkLHhnOZsg8INJbMUpuvcCR0
V6jEgGAn+jINzk7qxH0blcx4QUSMPstvciXeVF5u57XWk/lMOXNrPk1CSICZKdDhlTIhQk20tHIy
g5XMwOxUFPYt6DLfwD3/duYZ/AuYGnDkX9AwsMvOEPvAQTmW3zMrodmtHuLLHTBzMpHkUoiZp08L
CQRHs2Q0XedAgCSd9713uPKd2V5FNtXEnGxyA8iMT2UNujob+KlQyZGz2lc8eCz7Zl908mrXKu1d
6mzkUfFZQIdyOEOS1ykacyriWmbl2LRrq54M+xk8k/wHtA5cZnP3NsH7DR7Lxro+Y6DLHIO1w42t
1FuMvo+DatfU6kt18aTC5YV78MVE+GfKrsnqGN9S3XwdxSG4ZdcGzJ1S9ycv4YyPmAjlu6nWVojn
Q2svGbaTc2c+V7R6PPDMGJubVFJ/JGya3hQmRuvq49R8yKvWwRDKaO61nZ9XSJqYj2zZqlOpBt5R
g/rxc7wvIVC1WqQqfdahsyTpmSNo3XnhmdgrW9TKzNwMp1yIYDyzDznlXiIdWIVVEE63s9CLH9QB
yCERqH+rAauSsB8c3MoOkNXMmgpVvZncHLzC6Ohhrb66AZrdiAe3W8LjUP95Me2ugBPd02cyPVbr
W9B+dLT4DJ+VnWMcm0fzXyLd3k/CtXmhj6q1oa5b5iJkHteGHNc7NW8qYUSMsIIBkNjw0NJ25iF/
LVY2dDjlpkVdzNLDdTmpjkIPXxrrLWA9LtYkfWW+el1EPgp+8+fhFTdue+4i5ThFVRZwRsSdkpou
UaY2c9eA0BNkvBtVqU6XSDIA0GlHk+IJ5Kdxk6vqVW28W12Sc8UDIfMTkm2TKql0HK8fyZwyEDSG
/YxntQsiTLbwdipOREqc6U5MM1i5TLBLa+9QDcXttdPjt2DMV1pfbaDrzyHHo8udsykjJRi8eyxF
OpUUhRm3kou9f/iH1uGAUkv6uyZqtKbi/AUqVF9Vs+Ycx0uhuNXTY5NyizsQTvI0Ao1QrYvtl8sw
8Z46OBx3+tDTlVVjq5JUPY1ISTXfKuT6mJG/BgGgwMKAEXaRxbmfYT8hVyxgCDgzP4fcLh1gfPe+
SBI8o6XhGS34s+m/N6yzT2e3g/fMmwYXbUJx3MFLge7A/LQIlHpC7aSzL/PNaVLjbeWyk+otUKqk
Lsu2NPMxUIISsJNg9pNBvETjA9JFTNFSpK8n88/lz2wcFJ+QcouoiEoq6Qsw1UOFK1H8S6gyH2a6
YlABEYRAXBrb/Q2l7BtnXTpDSPtYR3LK4Yp4+eAGhSxqtNnHya2uNr7ZrKIZuIO4R62VOZsPBpDs
CN1D6NIy6EcF4llAg1sxfBhtg8p13rVTzE+oa3/3enzm0GYnNtfRoOBiTxVMv+Ze3c1gb/aa/5HR
uVVBZhPpKXSPiVA5L+66a09/6NqOHNIC3/4yilB3i+6WI8438nf+E0zpcBISaOelgAekMfZUYlJG
Xq7pbN/nmFjQEqP3UOiTpQ2DltOEb+uywGOzMl9Ki2ANXm+n/O1Jmqqt9J2xg4HfzMrzXw5OEYx0
J+4ROnoIzR2UkaVmhX9hJmZTXBSxW7ZaiNLwNS0nSNAtxKqQfGtXCjq4vHXoSDCVtqUeu4CK1mRn
oenFaaqPHSqiD4QMss+7hAOLS7zXGoK9QS4kA7C5bNuGhmjLgL8qSa2+WpDu7X1xxGawr5hzxJ+s
ch/PMG0FEfKxI1sbRgfbJiwGdKjY4BlpHGU6sUi0nY2m+9NgW+1FCc8c98kRIMeG/0YVMVnlorSW
huCM045/pQoB7TX1K+S3vXmnM4WSbGGF+EkYgM6G57kfRWQP3JGU1HDE+zkZZ4PPOu8ZZK5Oy435
3Ok9zNv2EuIoELVqKA6iPsb722E7nOe/U0BnGbHM8CBd7zaFayLiSrAFS3lojVXkQHdBApe3V3kS
2bs3VOgm4enGJ4EIRTXGfv7QZxGO/ZxNN8ZMqpFimBLtDWEasVV+fn1qYy5jREXV/pgEQcabUmsy
7/esjLDvOWCF8hZkM7z5x5xbrlw7m2Cw6HJ1ciIBeL7kyUtwFtijye8H1E7uL3qLJoCZ/P/MRvh/
FA+91W8FoMk6WizcANQVLbTiY8oUrOdYAw4exLWgvMEdWXWwF8xqQoh30DIdKAqiXtmeQWOgflrF
2CcRQdiJaORh7a0WwuwWWRJFxl4N9lGC02LiV2mmVyZHnTAhS3DdNOv65239NOLKKF6SW9UDdyxl
FtgV6ZZ/pt3SjdTQ1+g6RachLAe9t02wu4zn9IOVeEzeoT8avQPCVkpL7a85b4yQ4/Rp2KNKJZkH
6vv5ZOsaw/TpAXwftdy6GmwB0WbQJFh625EjesU24ufEsV8vYTk/wG2JdjRMiVVqukZcwCS452R5
IAXVjVyV92nV9Jvo/d89RcvV4U/yON6VuEJ5UG4ZWhr19fHkas1+L3i+2rGIgxcMYsvuUBUKffaw
OlvpGcUzl6zn9oKnC6D8qHqRt6kipmAq3Ih1nNnXD/YZdKxT2URokDUSph3jUIOOmw3sWypm5QhI
MOZ8Swu8VfMGm1E5CQMv59Bh98LzHP2wGl5B3IWWZNfElTuCXjIo0yOt7bfN56yCnt/WzbXYAyrN
umCsP75VrC5VlditpbmnSAnGRYlg6upH7J7HH+rmuXbhEZr48hn5q7YNgbHdSFng9zEeg1ZA4teY
UW+QvWotU+8FmOQJ62JikBpDDLkCcU9LYBfPu+M00Ou809vxWMGs+9UIG6HZSKHtIAC5idnRolgf
OgHsz1zVGCl1ZtWaevyYQJzmN5qorRAbBt0OcmFwo0xJ4Urpa34kwhGxe4yCnbvL7zRUagoSa3YH
2fOckKKRuyJwEtf95z/RaU8P/MBmWOPG6NOMTxW3jGFasSrJSmnDxFGTZ1E9UJxQYJQ23jia4Rwq
ePD9TBXMTxIb3I30xIlXxgo4gMmynQpQFiV7mjrcwY4DMDPgCoBMvNCeSePfuLIAm86mxXlOt3s3
OsENyYLoWCQTOH8tZ88GAiAYB/l5GE0rZVzRKAgQzB2C6LiMl1xukjzzU/ruC+N5rYC3mtZw+Ou0
5fjixDW+wW/H1dVi7JumdGRa8zEJ5ythaNpvs531KbdN+rhdE1MTss/IQrgjoXtU+RzIwlfpKIPy
cwiShutNi1uNjYHIFNpgpr5nyPUf+Tla+JVkm+kRK2WEC1RyerjUyXieUFC5AiTdOn5sQMghD4QQ
GqYIdRfk6EeXKUjIJmJznAhUthRwX3C3WoWBEosx4qxFFlMFqu4NsGl0tENokmrDqCUUGrMkP2+B
gXtukX9ih60OZNKO+t8D2FAMSEM9+PxZF4IGf49YWK+6NOsC7FMiaKqNklafnu1ezr9UEDe7Tqpr
/JZjK/tMh0gakCgyvK4WpcYpOE96HARb8/vvYrnX9ug4aOVSNqAj6yfse/YCdIP7uf31XS1cxMmf
rCPZRxAP4uyDMKGOHLEWmZVODauB99YtMKpUKdqCzH5CvzmslsK74YPr111Bh3rEAeH0BTIrK7ud
LMt/Ms6DinjDcgj7A5Wxncst0tES9alCwHxpzHIT8e3aifPMJ40A32KgAH6X6xZbK4L5iNzi4X6Q
NvhOX3U2bTHNbNNcEPtoBqV00mSitU8RnTtYo2i5x1xHweEXCwdanlS7PCFe3eM+sGZMLIEHnp7n
fTzmc1aYn7ewhMr44Iol84VzowZ8BQpnpPrCHKuaahiERDc5+wk6r/JJuh0h8ZYy2nWokAQcTvPL
ifr8ivjzzCDNQ4GufnSxIoJYHoJtdaZxhQ2oXERpm+Bm0XRVvWj072cH5bB87O3yAG9sXSMAfSdQ
IMWzI2M05FEIkhvNP64U7wteCIwQORlNrOA+G4ZycERlfZcdrzbfqloYT+xoMokiMdBKVIZkse2o
MJiMVdprXRr08lwuj5sg+XjdET9+SKWv44gnmW5kkpErG7la0G7haovG289zD7viz6/n1C3hxWaH
MA0tqWUxL4ZLJoOTtapEr0LGwrM/hDvfTIbElV+jIhmkMP5xYzRc6wqp45QrWwBwBmzlFPPVfKvz
aLCeNYiMq9WSfALwr7xm/W0nRECXRXgqnPX/xF6X0f8EQaydZVzZQOFNzgeCaLmWQJuurWMyucJA
aMCpEF7gQC5j/4sI1UZS6YiS+7/AmLhUWnOVIX1tKOuhnZjm1czlhEhH2c/VXQOUhAODwvjz/r+8
ZBLivQu0+MDxIUbYQmFDc9xc/MUyL50p2HgpgTXYtv6AQfawxNIKH2z/jUQyJi/kSEq+SndAWxQN
m2QYjfl1TXSZxNC8u5EPrT5uy4R9EWwZfF43oh5kTNPdK93/5hGdmciPzjOyv9AUrmdY5R1AZ1S1
ROIH5jG+kgq306UlokiG/chIZsRGlE9BuT5/A7WvSbwai7Tv65V7Bh7TnOQZ28E1GPIeh4D/yskz
hbISs6Eij/tWxMbT4vxNj9/5tCTY7LtTzXTtdnDfryVaMwD5c9ApL+K82m55PknwYMpoleHOslAF
jEiKY/Mo0M6jwaVwczyrtZTe3q6P65aZ3MiIZdlsAcIP4QpKG35Ij3tT+0yJZi9tDggUs62KlxZE
O4pvo9MWfiFUwqniVcJDSqETgyuqyH/sBMWttcvVEUoi3okCMK/42M9i/G/h9T3MfE0jUN/vjItI
wJ6c8zTS3jws8Dzeuna9Rd/6ck+TCK6kFm8Y4iQ/24QTj18+Zo5qqsGKbvuX0sPhSY70Pjsd0bW4
j796Pf8ius8hpuoaIt5NueFoBdY/CWZNZPWoKnHftOC2LMT6UfNjCTk/7d94IcL1E7uPvdNGgBqT
4x2PYCQo8TPrQdiggRXo0p9b1SBl8XYxI4K+wpbldd6YqwWUxYoaXc7ROPQ3lr2HXAy+ZrplyILx
kPrX6193pQNFKaHLyZwSgfKIYmkv6vqLQvZw/hs3DtxFYt68FuaHiWEBeU8xckRJE9fxSdN+G848
JauDNdY9L9dH3cUAqfGJR40VS61QIo84K7uaRc1UusnBLqv6K4lqxUE9uWeh5qNtFPDjithf4mDP
cL09TpIQZCTUlciVeKCPq/vXjrkN/46vbLyEOT3wL3CGNrt1dLf0Ccp4/obaHS5vuLkThyYqC9bu
VKHLWfvOzIAahD38ejSu6KlPRHUCRV0B/EcOZ7hGGBFvcxTpIM5Y3rTZIVoIyDOMguKzrhb9wvyG
4uwQ6cOZLxY/ZfDLlXIfmwepW5Mz3MDP/WJWnzHmnkm5eYmomidBwz9Gb7URVvjMTNC1RYy/wV3K
hkJlpsLc+wMBXMJsfGsNPGuTZML14r95TqXSMpK+kufAof3SFmb7dUljX+cgTPFW3JWN/zxyqaou
1P4ZevmqayYZzH+XA1dv17mMfSF4N3BgL+nBTfiDSt0W5dPq5evyl0Kkb5ChebgY/g9uQQms4qTp
DtDatPJo1hA4VQbgaddaevpfohS3QTjcZ/FUjatasgfuwiV163SvodxDpMKbeF15m8oVxS5jIXI3
Q5KO55pfunsqkEJNf8SPxPABXKZeTWacRYETaadRvuK42RoWFBb6BUEfM3Fv2WJBT+mygfuvshz3
jIfzA7MMVm4fY26B5qlp2hoEyMP0YVw2qIqKsEWDPHHcVv/xdpR7JBc1dVnhtCSVG3Q/sdZzd94q
ToF5i3YcdInOSna5SPS9Rh9fVcjrPQMWEXDQ5YzA8NTVMP44ppHxOnTNPkzKwDqaQTcy+YWeG+YE
6fwwF0e3tG7I2zCT0sC3cB1JyzahEPIifEsebjV22o/lqjwqwecFDsnVOD37EsIr0xX/fzOgjBQz
hIigA3KUmz+xcHNkUFuAITqmhom9ihWIn/fJaMOWrZ1OT65Z25lRDlNLImzvRyz5nsU51+XWBad1
raHSisJQE+3CrSCOSacJq7fAWTd33Z+vlYhhT/OUp0RltZW5eJiqf1aDr/Dq+KkGpdt22F4g6Ie1
A2NAxFMg9qc4hAXktKL9jT8srypwti3cynBgBYVeGlT+PqpdRscBTzUm6yfK4ziexJg6JLHo1EFp
4ReRNRGi8Owd/hClH8f8AUJLI3ld+w0a9fWoJoxZoJ+Fw+r/hp61859ZSFB8U+Z6+QAkb2k0CE91
NYeLB9k/IFy0TurUPFfvTCkN/nHqZvEGKTRCzPahx+MBLg0lO9tQYYvnwN8l8FBX+3UDFF1Z3P6U
o7zAqGP1xL7UCM/rSI5oP4lyBnnQMD3pfVHbhNb4c2xUlRsItz91VHUWpq8XsnTQHqUXMxe1tDQy
/1RRoRMoKSVh5h/NAAQ9N9WrjzI0EZ13gEvVf3sRoA2lZN7E10GUMlEHWsneYLYHuxV+q6j6CQJ0
9wci6AVgZdcmuy6akcnAB15Xsd3p6WNLUgXeq4th91fCHQ8hzh3TRsmWHFKhX8+T6B1L5uZcy1Ch
EG2upUZJebDjp7QBEG10dmL22PjfmoSj/d3N+v4T5GcNoEIBEgnM2jBUcHeJtQflP2DQIL4+/tbI
MckXV2VMPXVvawcDhzb6UNBxtd4rrOUaFXGb95m6RSlDOppKLgpDhJBQc/OS03DUSqi+ZLN4tUos
fRgG9J9FqOmU/pLERwE5Gw819eUpBLuGNM2s3Ax9OdzvzdxFtKQ/C9rB7ywi7sY3SHzWizVWkHiu
Zlhv8hg2MeZt9e73Do/sCtminT618rWt/yNreCF1VmmPmttAdTmPXlFNL4ikQqmehX697ePXtfC0
RPmAiQjmO5bw/SOP3YsB7myTkP8mIFhJ1O7zGP0ZbP4yxgIyVP/gLi4bv4aa6qlUJ5crHMowvH/p
QkySvCEwZ9aKxkBs9244JlRoi3QEsSX3+Qyegx8RmczAhxYYDMti8UhVIjeV65skaeLFJ+/vCpSt
UCxDHsfCfOpE+iTi1v49i+2TYt21/rl9vOmrIDhaz5Z1K/ZBxCPte2uur/WINLbxLDSXMfpeFAg4
Mp4w6LDnhYIPc+S/308XlGfgoxh/NqfiJY6Nr7KLO7YrlEbZuz7a2w1+dBbMVbPXlDvqOYZFA9C1
4arszdU/yfOPJYXo3fNTYNhyxPX19Ypvy6SorEGU5La2a97RQaTIXSg0mMyLB7xzy5nlmLrT6+1l
QOwK98S+R5uJg5vnRvSvRgpEdsLk4Edkq7bBd9wq+3/TyMmHP32JKc2ITQzkCgLDB7zzWFTcLyM9
uVW2HvRBv0mlIyx2tUXUxFSXJQRdaBgFlwbsQOF2+LDopSim8wkGVO2SPzEmvhel7aRrix4U1ELl
oD4F71dsXub3gtFBSyL0wKlCj/Zt4gE+oKOEhDmuOyd+5T2bY7Kal42jzsQ5Tkf6pEggeSMivVE5
hoYMNzJ9IqoMvGube6vif4kXYtQjev2XDXLO5cn2T23MLK0cde6Dm941T3SODuhfjIvruZ4CO7Gj
8v3rZ+x7RdDalGOvNOSpTFJRKXr8Swl2ZrWeVKzUFYC8PfXGaVOHFMvKaYqOgifqc7qIN62xN7Ra
KueeIrEDRaBzY6wRz4kIluLTMetjkRyr4rfVy0hGga4RDp4Yk6O8G+i75ZqoJEz2rMyCLl9AMIko
ptwV6UoLYE2s/SrRVBwySDh0tuqBlXw9KB9KGKAdx+NrilzRsV/7dInUSVMBVQEGG1YiwWleA8JB
aUyGANGXIIMgGDWmmOeIFhEzKU4k+JEH2qVvIGQT6I5Xc6ZNFt3DOXYpQOOBRNvlkSYKpPqpW8fg
tCtPDn3txJvvQqex7zDGKaVtVNb0CxAy+l95/RJ8K/0ET+oC/r5m7qpnpYZaL5T7a4ErIFDsYTrm
nP41G7AtJ5ohpQIR01LIwA57UvjrQf4Z4Jc1TUZTPeUbZM8ncA37JwMh9I4Z2fKgXf8Snlig/2kV
4tLQ/DPZt0xpdOKmyrCYLqBlGQqQ9lYBy92midVMS78bx0ZIHP3uchdmD1FpUqMJhdrAZalcW77M
BrVhz/iM3XI/cMJse6dzQNof6riu+X9w7mfEOEz0VIxYqfSS1QIx0NPDOjJ9lIiFemjAOEpS7G5Q
skE4MXkVKCTRSgIFNLRLT5PPChu/4MmvvO7lG8tjsQM1cgM1hN+lQr4QR2hFa04Xz2IRH6vBPojd
09DXSEg2/Nvcrse5gaB7mTJH2OGlOjhHdGIek/1TyJj5Dv0ClKfb2T9FyAMbpiozHEslzUbOx24e
DGAumYi56SzBWkorgUM6/u9arErG67GW5DEVxJs/ABDwR+CMcoDkMZU2Fbctz7XIna1I+UxMQtmK
ctfflHdHOR6ytkv3Q8Pb9YvNssAYoiUDfZJXdzR5c16P9bQz9s8K4qBfgpKDGwh7jf2UDWra2w9Z
xqU6uA0RB/gpxqxgvQmikLuShz/p/2a1PSLZK2EhDQBFM6ML5ssIxjiUtAnx5XTT1BcUtUx5NIrU
6mAKhojZMScL8lB/mfSGB6uX45ndkBbQw5FI/tB0sd/Nc21rGnhNWEevvPi9bP96Ld37uDd/PNRi
a8zQDQgH7DRTV8TSieUrQ7CXHbf/Re9jt7pbUxviJeVIybtHu3tV7VXktpLIyNxt+d0mulC7lHJO
5rsofAjwj7KBlawBi4D2OpB7A0Itgi9nGOXeRKxHRyMIPHC//nZwOGLmhm6xzMae1imJhSkqnxfZ
neaam3maBdPqHlVNh8jwrK4OXY6XNNT4yDPzy5XkKES580SwqoGIcPxxm1/Zqvf1efv9qRaP1Opn
kvxmUfp1ZzgptkiXdb1Gd+rLg0K8Rjrnav55M3M/oMHZ/Pj+eOb0oUw8WVwrIEKrleYyfPZVgEMC
wMvg9zgDativzgidbIU9vaKO5vbHQIn0LdJPhjqyCFFLfmeUIyxct3W+F3yeTTc69TdZt0pNwr/8
5x/KeR0yuCn08ztzsb4ISHC1FiETMq4/BpdWw0/z7Iw5XCvYbmW+zHeaSvmUgRLgfksGvtAl760O
Cw2cF8antk9LO85RlTZVNUsMLlhMwni8w7aeIgxlYQNU6F9/ZK1XGZVnl0P7T31zcilLFE6WCtbw
x8eZ+iR/gBFJpjq3Ne4PNUScIgYqQBSqSU7kxsK3kXMZysMDkAVkrpA7vxwWYnJcb++nYQ6ivnc4
/goHwJEEg1R/TNMv0ki5DGvTGYdF/Gu7cE+nLzk32nvvebHSk21aexlRljec4qGdsuRSYMhTrUHT
MyK28z09YXWZwYRb0HKCE1stm+H5bo5Cv2kbnIqaq28hi8A/terR3pWxPfVQ7B/11tSMuV4T9aTU
mJgUV5UG5CtAmcbrdKhhOh7PwubX1aHnmJXXAHLZPky1ILz0sTxIQpwYCU7x6sxwbKTwjjQuhyyO
UbLc+JmKEKlctLPn3LZxwjIYBmakd+K/D6EDSf/aEWOgjqkskukhb7/qVMzh+mRIyBV9ImMiFV8g
LATjPDhYbnomFLraTU6sy+mPLRbCXQMmXb1XirPvNk9CdO/Qyu1TJ5+sXMkjPlg7ZYtTwMk98bdo
IsQby2Eni6G2ktrPMxhmog2XH7WM6ILgurB7lZ5lDUKBXR6gcbkVXupfP+cCU70z6/5d9VOQtc+w
WgQ6g82kN0S8ImOQr5g3cdASMmlZhu5O0aZGu1ZKRPHy2hH/9yiWMZPiXiKuTJsYSm2pFEW1n2uo
YHsvLUjApuDfG01cjbwjHaDrLWaJIY/2d5ZlGIBPQ6pQvJCFcyAoN7wspgtKQpMJcZ8BwNXUypes
1RtJg1uMmJNMeL8NpHAy43aubPv09i7smotQ0sSTzn9+9efM1olq363kDQC6uBfrJttWjYFpKfpD
uTisRodCEQFHSPFCJjclzjSNgjp4M9FlB3RHhu/rKrLoJptY/8MFHDCcOZyg7+pOBaIGz9LSvJf3
JZ09XUKwt2OFv2y7iDYcWBS7GeNZxZxj62uXT0bWjBh6fp72bW5dkQgiY90y+7/CyMmYWH/ODk2g
LT+E58Y2c+0RYtPv+nSt2hxH5Sdnhgk95ueq7uTUsR6ARNvRmvjJviNjAbVfvnrCHU3XVqvxC4Oq
S3TwAofbdeFw+UPuSbnsVCMZg9IKAsJGaUl13y9rEei5Q3qO1cYZxiGYsSzrHcJIiNfFc+c42oUu
5ewXkWXPysH5vvSudoisnuaQ0QgXf1xr2aVBN0KCh+b4hosvTkhVHhjaR5+q+CaLBe6SGhwvH7KF
R2KJIZlCsuoTNPxzqkTGW+Ub5HcP6XRCAUUXgnwrcjQ2ItVLuuzbOHCtuvUG8/Fa61rCiucmnNbL
gJ0aOPKerggg4HSJEnDS45WRwxRq62HMupTgLOdhgAkVZ7AHJPczZjwSaN2E3G6QrnTJtWcPQK5v
uqcQf0QqOnpoUunRjWNV5ZGJs8MvFmr805gIfnypb8DmhRGeLf2mgYKGLuU+pyTLAp2HBFMNo2C5
hTDirh65JKnjiErfcxtnpmldnf4PyCGSsuEa1fDJlKMYHjSkESECX/pLvtEQ3ShRSbzeX2r2AL0K
fbVeidk9qGfV6dUCq7xYvla8N+VqnCUxX4FjG0GnEp3AWKXGRtDWTzO3TzicBPjrsSZShxdkigWt
UhsnNQ3eo8rxsQEP9zlV+S03QNFAncjlgAIBHOCB3lqfjGNZOuHvxbbM9Y0Q5xqD4AIwMyxY3fla
hjd9ifpfuqbKRJtW4ROXzg4aAOVVtlnnZhz7FT/X6dE9PZi4eNL8MSLOZVif79WZFM+QMofw6yxe
ZC9r3rIjoJyk+4gxLkyx/OLL0cZBoUxPhtfitNmX8+Iz9FHMCqysVCUJAzvPxPpYtWoJgnRGAT9t
KKtrkPIHJAtgjYxlT/vRrzVPpwfS38mGZqSzh6jNmYXa9njJp/p89F/fdSpcr4ZRvsc0f3Vwn9BL
MDJ25UxLb1c7zDgGb32XlscYfq//HED0Y+fg7mxOusTr0hrC3zol+9ZIwzvF3wRfSWZAWHEziTMy
qmpvBbiqq9itvNOKbxsKZg6kDjZy1kC6r1Z2Aplj3+1fuqDAY1kQwpjF/Z+Qa5SLivTSqJaxlDtB
61A4C5Ly3msqCgzxpKhWV26vqMsOlZmuvTq7XwHtrbim+RKa7vPVQfaHziHUfEsWMYMOvTQZZeWR
0/wxubZxRh9Y1IG6dgOZ0CpJhCmDirV9mYAAwr9q6rV7UqkT4sXw4lbl93asRfZwSBH/79hWA7Yf
qLQ4wsYoRANRLcvXAqwmbSURiPNqXdF8OstQbfbo+AEvAFP/avmxFGBPy1DtNUTWNmoQv3G0fmzd
v0PZzjwwoUil7R7GdQz8OZ0pLGtCHID+BT2SZIUsLZ0AEm9O8cL/NtBhDgsa62yDbFBKeWM5bUU+
fYNAQJB9P5r622ewfhcmhqGK6EnlYtN11+1lK6HeC9TZcEVv0cgWY07xue0jgojYWsGlv7nmw+en
XI7O6Ia94bcveblVxYYSlgBJdOvAkMlQvFc45X1EafToO89utOJx5ndnb7m7jTu2ae9E359R+mmz
wTALnxoohlohCTJYPFtiMNKpxBnlpcaDrbjqhfpqL0gwo7yGLGESRruSw6dP4KEz1IBRSbmLLFZn
uypOXo77rwzjewc6J0B+IA9iUfdSF8Y0AyiQXLP405q8vM8YPQVfNFUJpqF2mckLsGvkhEO0Ok5b
xWfivVOu1u3c57r0seazwES+bn1gIT8AqN7MJRSFmV7bpgNW+ZMXlc5ZLAZSceBC5TkZPa/mS2nu
FhHcvwKuS06sbeHLcVZLr47AQCzSpvV5YlEVEM/1kY6F1nss8/aEz1f2nE0wC1OiZaC2hFoh0Vbp
D+f4vyufI2OaQwpVAxulOVrP7flps3WVp7Sse0o5hvewOi/dbAezZ4jqjOxsuxklkhSzX++we4dv
liIJExLvTMSpmgGA2W6eVwU7/c0BqFK08jNKh3DFZj0AzjuwJHdlhjBcj6Y07UU/UoVSV6/BxYVl
wdfbfgTiXuKiFFez+hRmar+Xq1LJAud56KuJdmn69CmzqZ32RRQZUcjcCy5835N40ch8sG8ffXgz
guk+8eYe7PSyISBL9JeIubGVGqTOfRW2ZVI4L9SfuZ2pM4FYGGK2qHSCISrKdABBnPLNHvz9U6jJ
DBrTa1n1pKo0hClWIT6jIr4LoeWUckmN5MEdAdock1aTfA57wqVeROYtIbyjL7lveVwpi8QePnMC
GogwCpYehre+cgfJuPhMrLD4Xd/A21eDSpGw3yBNcB019dvTKm+aZgydY88YNjYeUl82gfH4VxD9
/PcZgzIGzHAFkqcLKLb0kHSe9Ys/W1Br2M4zVeuasBbVS/mx8PgwxMHlLvvDiv41JKHthQ+zVR71
pFLxLw+bfnOIlCcpksXJVyp/4Vr8Nx3suhNPHNmKS2SA2m6VSC1daeISCZlsETW4d5qW16MzvWtQ
Uf4S0M0Hn3Emj8o+ebV3Da6vPpod7u+n5uA7Fa1gj1qFwSCIaYHSsJGD7GMT/xvKZDE5YmU4UFSv
RmJ6Pn6A/r4RB1227zjK3C8N75dKlK845xNHDyCn3wyKr3kFqMkxX92XSBgzc9c2QjR1NdoNLFm3
sW1pbH669uWeZWxYqWH/mQhtGbw+fJcWfTp4eoOEmjsl4HOJnR/71BJc4cazoRmafTuXhTkn+ByN
JBTED5Aupf+isMiBUS1gpCq+zN6s7h+1Si06x0Chd2NinLiENZbpevSvHVMfZjEI2tCiKuact2e3
Nf8UsDARPyVM2tNGQOjAIhoFkRHJrzt/c062nzC2PdTP+J/DeJH6gWSbihc0fdZ6Q+2B8CCr+d5F
VwTjovcptPU2objs20GEGxsdiOl9s7y1cQZ8eXdOsxeJsqt+T6pYhZrrYdzSVuJVc4fiQjuiL1QT
YglOVx36jMHDgKmp5z9gLsCiOAUNH2YKyY/ow9a3BXiuHgkQcs+lCYhHTkCc8bi2NOWBmO51HP2M
fWU2Ci661jzb1b1QGRVuGr4G7HLlLkh5yRcAbDTwrCA4r5pT3xSA5kD/XpER35Cpiooe4vy8NIoq
GKrssFkJzInJ1C7bNSF9qXtamny0cqUFuMa8vpFYIbUc9WIX0W8FG0SgOoivuYWcNi+JbTKct+jR
S5RRsEquTaWNaWklr7n7GRykUpU/fTQPMZ1wwO8ny76VkYFOXGbCL/b2VZsP+u3/eB89s3sR/XmI
ZdKSmR4HUaLdToU1w3e6dmpHNeEXvw+ttUrX2iIpS3uESKm7ZhzkP24+D2bNqaaPv593iObLl8Jy
qyovvBntkbn6/3DAcwdHCfUGydyVufnoRXmNDdAd8/Ec0hEDJZYJSBqeL+GGO9/9ZnqYpEKN+DEo
pyRy9nH8v+QsGBwM9Thp+U6fWaGVSKv3W2xoGtZIo3bfcIAty0suyu1aEeAlg80QB3RsNUODYdpv
zy+py6XIfhADpDB52N/1XsuEl0r0RtMnFXbP5Wr/EDJuJJ61NqCFiTMyYSnIflNPQuFNZpkGjWZh
jPaHm2WNDCytBhI3FddVfIIWG3qKNpMV9ShwcjeYBKKhfEzBQyCoVca5FGepohEMBJkrFsvi8XQl
YH+i+B2yw6kXVtpOVqTZI7Hf3inofU9ysIhaTvBkv3Nv3TGJAAKfz33lc20m69mvRxjnPFAgYMl0
fT8f//JeMGIpwVZdgFYDAeP3jCNKedJ+N/9/k0jzLQKKbeNUXMAQZ6petqFrFaEKUY333KRYGmua
jIFcaTo7tWtFpUwwcb0m27MiHOC3BvXNMu653fQnQ/8waGNLEaTzdECyhBYUQU46EAS/12sIqok2
J6eeSpftYvdGI1EPW5fOaDr2jnmcIKUwgys/qEJYVTdMDRNjmPTjred9oQMzZglm713qDtQ9ybE/
vzCBo+O20JsyHdxltkoPm5hPfTuWrQW+kgxt/TcR9ocIWKKKQ0+/9HghqMjFkkBAuTjQ//zexnuw
hntG/d13ErItjf/zw5rKZPcBzVkY1p9GnOk0xdcdeNMFPzXyoUpqWc28byP23DfYZKcofkGbhyze
HkCSYkzVwbjaRY4MugVBQyRK7gQ2+DistiIvJzL4J/yFTzZWSmw69EXA9ALnVb0jomXsUjG84SiW
rPIA90H2P8/SdoommlG9SPdtmFhmrcaCJ7RBBe1+9nouIWGa8IjWwsZN0uTo0FnjI2p4DbL6kNnb
j07G1c8gVaanjatikuxfuos2bq7fJnEtaHfOpWAwPZkIiJU3yVu8b4sLUiZ3JwHhUSn8VnyGmCva
tyvHnD8z6cl6AKFqIDJSmLn2onrZCXKk8zZjcETiqYoDqSgRZcJPSJSGlumFdvQdwmGY489zpnMe
wPZYpAJtEbVYkFdQ3dUAQrqfHWQBjb9iEzK67X4neIcPSkZuwtTNnd+HqYvyN6dm4SdKH2gRHYZD
q4W486tVluqocm5f9p/QmoLCC3tblsc7YSRX6USXBdqKSOnSPEYIzhSt8NDhuSppRcjio6yzD7k7
XQhtYuFJ/KboITj5Hah04UTsrbm/C8+LwQfv0JvwfpUu+JEu+uzOyGsmHsOcQUokyeIKQY7/GdZ3
bBq9eLKPWE7HWOroBskKRqYKk6mmixsEpiFxgWs93+GNLgBaDkTL65tKHfMoZ4CeHPVZTm2ClkZg
yEGbEn3+LFDjnve5lZtZgxFCZtGD/ZxOh0kC+90ernT0KOG8M8A4vh/0afSYlXoN3v5q2mdQgFTV
Wjrbzh/A8lMsWrlvGW8SX9HfFXTdiNAR2011952iu9WFTPXVKjrOszrBohrVEvtngEn7kbPtVRKP
KroNI3FZ6q8WLjIFlsgV60Z7MELM7cBywyyJLOg3LA9cmyxNLomZ28fi8KR2biFOpVH1AUJOJCjF
JZ7g24DqY/PKI/VhcYqZvM28Frs2lrlRTI0WK8CVtenB8EipxMpYLJwZyiBGS25qwppBDV0yI0/v
h+n/sHM5J1iKuCxggw0CUBMpEU5tcuukNiM7EZYf98Zk3cen6Bh+OqXA1l44P+u7LNrXd8wokXuY
ygfsWIpMejQQF5uIO7dmXLGgTxxb1tQMqiTNGlyxz9F5Xm8L7h32gZHA0FN140Q/cpfpS9NejZWp
Bp288mh6iByEx1b0TCeNRkIxnqCcXVXqtGZkoC2EZ0nI7c1Kqi2X8+7dsTJsRGyYhfeHc9kVsbVt
lPkQzoROzS9RGiAMtUpCP/+hXDM3l5w8994ys88V36kPH5uljkkmtcQ1ntz32eUMoadULO4sBQb3
IVs+O/mEfLexqQzS4M5oGRTPeIaml6tjNcpR3eUsJM6OGpK6680X8Q15PWYnrRmE4HJ+Z1bTIjrN
Pm3iDcQdkIDOgVf75Qm4YSdL07v8bRMzIp8mQgEAM3bjGjC/nnwXBtZiBSPgJY5jwfCblzpThQz2
yK0Gv1ODOIdyaa8pEIsCNkOPtxhQPtu/6xHNpBirDzbZi6WJd2VUiq0IrXCosQMnHrYRhil9RnIQ
YPENccSG890uSpSQgsxbg+qtkZ92Nfox6H9TLc/5ZJNrY5eFmDiX7Ytq4gtiQ+lvC+Ggt82Es2pp
v35EwV4EMH5xFWKYFezO2QcCiBDwutU4oXTTqrLnkaSszS2Qip/NQ1zJN2Vm0Zr6+jdy9CVq/+BE
byvaFuMXDmsnuWwu1xlcKOlILgBvInKVqLj7RipbM3ptF4vKVehFVyPF0JTni3GE1/swnjNOCha8
CEW9x7IlPtUMurZ6vDlBxpcC5BGJJo9F0KFss4zrKSel6YvG2vi6k+vdJ41YxBYWFNrwKlkeBLgZ
xv/QYJsu9UAruexd3k+FbFUTjFPIC3Dl30KjCmGEP5e2KTAgVX0bO+vV5vjX2sy8Qhjwp0QHR1xG
knXfFhw7kUzmL4uvPn0zBvv9sn6WNMj4KPNr7kssxYtntZB/cLbKCepPppkKPy50VkFdmXnTH8Wl
uVPme/5Os6GhCVYSerF6BMWnrzQ3ooZgKVAXzkVYfMCd/JkvAmsasWBi9b5ZuTgspNmv3bCD8HXi
JNvZOXOt63mQIaHTaIVyOTyVgtkTQNxx4J+L8ZQLFNNjL+FJfK/h9+V1cZdQ39EvqOmSlnD1lSBp
SdOFQ/8a81ZCRVgJDzxE/YupaTTf3TXZM0e4NznJc6Gyxje/6boqk7mOs1EYrlM7JD5w443zlbgo
o4o32Rcix2UeujjIFZZmY1lIM1Dw7YIHRfnpaOHajQo0p0yF7o5UeRGhSmjaVcJgc8jEKceQ5a8v
911GJxW3IVY7WhsC+PsoX8R0O4kiGiXwWn5KFyKYezyzepqBt+CQUPuEQaVnkAANrfBdp6rDIOax
aYeHjRL0y0Sp9tJmeP1geUFAMFZH82rOWj6nOFNQb6ZGX83xRK8q9GSyb9has7Mr2Vkx6+T/OuFz
hY2ggsq1bUWU/kAjGsm+5YYjPBy2RV6G8Wojazt/hzd7UwKlC0uSAgUct5xKYPwd7DS7cAvySPg6
cq4tiArnV54y4EWS6qzLH/rw5ACIhRWukvk0YZp3jqL//Wix+lqTZYa8N1jTd2StNSn1wacIv7wn
S79JA2Nso+SX4lGj9jFJbNkUM/lb31MbztZobXE7lpOf21XKMrKpa8CeHbulkVvoIu3Yhqdk7BHJ
LrqqbV5OHAu3ixezDtbJEQaNuOraGgm1EpBv0ijfWgyzyAY045Zsa1A7XgsPJoo5SvAgoN9EXHv4
mjF/fBPlEKso6QiLhvqptijPODtuGipn1AJBHAKjgAQZZeUJ+z1RzWL0p46F5S+U9FoF3O+3OynI
vzBDPh4V7aJXA4peSe6q3xoRwivIx72gV8KJ9+xXAzt86Cg9mioQrjWPVbtQuicvkSr86W7ndLNq
wI/9uTIMSkpMAmzazG2Mtn/45HBTcPkxLSDj9WnYnWsYXKkxixmOVmFWfz3c0S27w0k4dtFzPAKy
ey2jaIwKztEHH91W97R6qqE/hFfG40zwsdgqO/5Om3myndcPO2pxN+gDA9sC/7rRmahmayHiLHPq
M+/JKOieuT5vlZVJAedHlx/BtkJixpnxJ9KjXfrn5a6O+PQjGVfsBGlf4ynfxOle/lwhaoxzxzc2
xB7/8+W3aPgP0cJvP/zjbjQn6PrY8OBdysKuuUmGozf5HjYv/1rmVuN/4a8fT442WGXn+XVysGnF
TUdp3ytnY4IBNItxlYnrEn4kBgjFFSW437ySL3cf3j3ewuZDLQz9SltKU6bCEWD7aHBOAmhtkXbD
LLUovP4YQJ0Nw7anwoOrf8x3GHtUb6dJVQGvjNT6HBY4Wly3sPXHBVKl9mQ2zjukyWA6lfutfCVo
IV2FrQpSjvkxcHUv1sp44X71kPOuL2h4JJ+aPjOXAcDV14UkyGV29GjuC+mMGq68VN/KO372QO8c
GueGraS0YqFYseMWqBmeQFMiaS3aF/KtxkkG8iq54OYcpIPJ9bP/6grBiGLyzA10QVaiKM08IW0j
bEIZtg5F57Er3hU+i5YUyokdc7dE5E9KzlMhBsPqGv5/KZQWH68oITA/KczJ8pyHWL4w4g8CmPEO
IeVuUlCPbyGHa+W1ezX1Fd0APK2SQ1KYlyua8QbOnoqOrpoFsEW0Qp+a3xBnhthSXKkGG9PdX6+A
WkQzKsrTbK52zzzYj8ZQCgt3k5D1PFiWxrRI9aYHxmmBeZgcHzvFRqqXxmS7fCiwSEG53rRYeQ4m
JYNUKrezFaW9jaWs8+YhpRna3oXbTSKmgpklrrUtQKhLGiMz/J6riTNkts5s88M/G+tY9dubG8wq
COIL7E8D9HW9tGsffkIj5bWGd3Fm7mulTw+V2bQPa87Qgza7iOwjDXsIqEszKLhNCO16Q7yOHW9E
s6eSlUPWNxbePpyKGIHjjygsnXPeP1vj7z47dAgMc0cghPHBC5Fxv4CK187B9Wb3yOoNlDuplelm
E5j5Ab6AVR6AlPVu7pxsq0xABbKG3rYeU5jJJ/kYpw0vMzUtr3I89O+Vl2w6n2GI/9jr0AOy0END
48Xk5SO4aSTWpnL+aBvgBWLq+VjwrQcg+SB3qJeKoHPOnB9o9mJtzUFk1waKO77k3yUGGwoPj5i/
IxtwtkdJCx4G7u8+dhhGUxYf/P4UdPoPg5m6UF8nJLc8MBsp+cXdMTzvf6mRz9cZsJ6yIec2O9AS
+MVWSrWV+OLPuxzOQZmfrj9HfVRJ6RFS4AiofwGCYdZvFf2Gmm28FNKyKAJiEhZ3WwHJvoheUqWM
xF6vAlFAcXeXlispiIvBY2oqJm77wtfxXwz6LPm/5dmWe4pRTT1R7GXMTHcQ21Qg5NTP+7msQ7bm
7yf7EHHJHtY1u9vMbUqdEwJpb2g/v/A/vrwWEt1vscnG+cxUrmpSRZliTuqIfvpV4+7bPlZUPSIO
HATX+eDl5FJ3h8hsabV8RtFg+yflCqY7uxgPeTN9T66TnyLVbKYTlAN1IZtbzwMJlfFyv9fpJ5dc
5Di7Nfzjwlv9Qu+eUXuat6o/pWf+cV3/3hFoT8hy79eznrlSSCFTWat8owBGoNgbwtRg55y2QXDD
7fG1FyIn3AqTroFgkJJPKJYf6Mv2EimN91Aaupcr8gYKvpBEYqFLzn8PCau3xiIWUayGoQlt16SY
nkOwCP9BUNRgoCimff6IUaMsNTwB7NxtYMRHnFfU00gdt6X/zk72mZ/TSrkTittqe2BIsSqVrw7/
4GBxvxjZwlEgzftZleBjREuNnfWmz3ZXYcjIe5BNeyj+rvXOvdTfQPsOgMgw5ZPt3p2OdJI/mzDF
NUBw5edn9GF0e3f0yK43g+eAxsRL8DzY+B9GpPZ1DlCX3g5lXa+TQ9yYkd/xQ1H/fiBMu1YV1JEj
RIDHmawjFmvl3OIDWMWKowfzacP5uZe1mg0QX+uCSgrkvqUiMQUsjSYeHne/d/7tTW9Zm2CsSmRM
a0PAr7VH/27/SyRLZ5beEcRlXpJBcjjXagxCi/WfWOQA94qZVhtDxUXTY3QhzqyCl+LK5IM6dVHv
B9+dHe/0QaaPEsjtCDn1OIX2uu7CrDZ73bdnel7IfY7+5UkuaGj6QzYtgZnlaCKj5Uo4krlMEMKn
HuabLGi5BRl88XOwxN8B971j/kMw2FYEC7UNK9OtWBZH6aPDR+oozINaISLlOGA413jeJlbk2fwX
bSVOeFD4FO1xxS125PLPycqN48fsj0l6p0tH264jd0AvYbfz7rYu5rkMo8A2FHsCvdNQ9uShCgtr
kaIo5TvyssURugC0x4u/kyAEkfE66QUgRj082krR86hgsX/sdbxGmQwu+iJ1VBaDwsECEnupwit3
uD6W6QcI2HDxOZW7eADdMEB3up71qDpA32H0xxpYF22YT07zLkaKKigEJs+77I6rSmIDr/MhihZt
eqmF8+aHbtWQQxsHKCFb3Tp8ch3HmdeoPVMBDWCppJ1fiJ62y0vQm7MqUZBerZZ7kAkaW+ntlcrJ
WcmXqdV3ZkNhikPNIGSjr7tPoNk9HBCTt8JDPxZHzSWqYC4ubC+ED4la6rYJJfZ66cLTfDTMB7gd
I8g6o/ylqBHCRqlN/LU43mBk6NxaWCLOhiKBnKr5AMpFJ0RwOw2HzXUTvlb50ssrj9C0xkaMPLM8
d6Xi0VPuWns0t15s2rb75NulOgiqv4bFyWwmyu8VkG1zTNpEDdoYZ1m4cp4JQLzJctXLTkDLxvGL
Ay1I412mrNa8w2QnUPoid/DpuOzYYuZYNG9Fu+yb1dRPgmX+XZL/KhIzhqRSTb3lcCGnrkEtFsQt
JW8vvmAydZTtB48f45Kqarywtzu4xldjGS0C+2HnNeaDiF2ATY1bFQO2DFuKjnvcqTvLeVmwWakc
0THuRkouDFBTDkj14kvbLJAtTCx6W/zDeuo0ItIX922LP+iB2JW/9sCzrN+vQaLbnSFN3Rr+wB0t
fANDoa2tdk2sjCuHiEQY5bAYPiHS2dnfCBj3YtF58Lqcfe1yyjSDAE8wFNPQXxjuIwEjTOOaV1hp
C5q5C98Ecp5/t1IhdGo3mHqU2W20EfOz5R9NU5tTWt7uPKaMEzjto6DPvxIceVyr+45EKR79iZLh
wtQTew9ga7DGj79icxL2EMd15jQhZF5qqKFCwUuJ5i32l3YLHVOa0b7u+8MsHkHd4gBUufZ+csAV
tmLTnPrinqk4+UBYfUJpckqM8+AlVPsHu03hgFkwzwzSz264JWspNsWuvduQPxEUB/3b5HqTrOma
6Rb97Njfx8x6IbBetJB3CauW3a5YLklQEuEp3ENZa/F4ZviaeRhFZqymctUiGnAxEDnwtCPnc1P1
XsTGDCekEprBjDSPhMepNXAInjcKYCGMy5J0b5FhITH+VZdicp23ZwRNxNvxiyf4XJvx3S82TTZy
1wpCNudkcGSHNACrSSZ0VqzcZICMNIAxDBtYCyTN7EHJRmG/iOrDDJSyq2BehM+KdPgp2H6SA1OS
ISwgCHo1sO24mM1OJWbWk4r71I5mYQlvLmuelj9Ixgbxy25VUfaC9pIjXjv9by4Cj3ZLbjYMujT7
hNmpAzQZZpEhQDgjZdv9MKhQEuo2cHkbGLqv9lLZ8Pzx5rioVcJgxHQkfW08qujqhdPdrxn7UJz4
AI4rPfkuhvEizGrldl7PnNS9tdcs1KFF5M60wa1deiIyZri9kXrTMXRjgVgUPw+OXxjfI8CnZ4dF
sfSPtVOpM65vMpY4KWOv8Pvfe7wuAvt1vAbvNHoUX4fRrrONXnm5nWfYil6dr6h5lIfjdc5Jk+dH
7q1+L5ln9jXeLuZg6gi5ndGHKikB4lcetRf3OV73TjRjdnGcPO8cmpCm2dnTHaLKiu2k8GH5zEPb
ixXvLDeaiAdCIOx2NkLriEvdG9W7bQZbqYSbQA0cHr06MyrZVrcwAI1JPJYztGekITC+egqluhu2
4hyop6W8qEIlyQ170SgovLGWOwR5H/bqKzMqANkBEvpRjVmJjFmI5mJ4IR75NHbxZo2G28zyrRPN
mHvLfxw049GcRHgc0sRWVXD87jMojc3knATB6BMuoHIb58LMmXJpxL8aF3caQoNeacCZY7ak+Xi1
StGvC1zPFnLLGjnfNfouVo3UdhYlvUAsqm5GUfJ+tk8Mg3tmgx+ASH/1bYu2cK4WTyQ/k2bHkCww
+hI7dExPK86uDrZiNLCLaqUqAPXwCLFR/VzWh+KG80kK066LyhJyDRhJ59EKlqMdcRmQc2ciDkS8
lkhiojhJEuE6yB7SIRzw5ekP7flOPUCMC01UdLp+d0EADGodDVZDDOaT5RlqE4lj8ee4D5yIQWDR
4GMHz1myn+pftQY44UDbeKg3FlZPGr3g4nJRUteuV2ENRcfJcjDsmy1KK8K1tZwebyCyblIeld7c
o1IGNPvj6cuaiRdrCeLNDCFvQajmGzpIBEzS0IPxR+kIiTNEypEFo95ue1NOUnYrdMHGy41m1Wrc
YCQ4FXcJ1evQibhwzPhumEaLNXTpVvEnACntJs7+AGio5xqRHL48BXQ61xkNWndh6KKiNdOXBCXB
gBEws4nFUhAGwF9a3kAPdZLm8i5MgUGLPWOCmhRgS0Yr/feSx/fyW0ZsDaVPalP4nRNV/yuk5e5A
PeyKsqmBBhIZpOG8/EIufn91YoB3/spjBy4BwCbfVzZWwzDNQfnYxxJ2MoukjrblZGYDpe2kLrin
iqTFVcm/GdKVLbP+143RviFs6arm8UTERtgTsBcOJc9D3R35/pG+Pcm0Xzbpaa92QMGth4Ah5D7I
n03moBl842sXrwauG8VJXi6K3FX4m8l+/wdmhIb0rHfc2oqs3aNJQtrNi998A46w3LDIxBjU0tp0
hNZBF3MhPbcunEcLECCFNCw6I5CZieVKJzaJzDDwPaNIt7jMhSu2jaJYHMFvR7vpftYdtmKWza9O
REAf3CRiGmNmJIoJ4wjNtHCNki04Lv20pjJCND8lW7paekHk+wrcFhwxTuPJOhu6FSK35s0QRu4d
0UB+Owk0op1n1NpkMtca0wtv4lIvdCBkLIO68nu3VXzU951UkGGesZCra23/pz3d1Z7hRILN07WM
3C34dkVE8wRmMZSLkdhc3+v8dw/V3TLO90qVJo03N/CLkH9rGVPwyL6M9Of2pdL5GcWb7dhQOR0z
xy+UT1zSQvmwMxkR4OCLobWXN9QSWi6KfqQmaBDQIm1PXJHy0BrE9YubgSdMaILKf28FmV5HxAZh
VlNx4cUNhoePlrwR5EI/1KnaN4bZcRUeWKBiHFXdwAGAASDoPsXy1EktXcJuEABJL9PFVwhgpy0H
B1KpHLPC7ml9o9UO5lfwTxqrGK3VrIOWc+/tHUAGAFFhz3/4MUKb4twndAbkzzgxxEEC0lQTFxIb
XDTtxeAHZY9AHTv1SmMtd2OSZvi2uQ6wdFitNili3SwWewjOv4r4q9h+9ytmDuT8Fe6vsXEh/rQ7
HAU/2ZZBSafW+SU0AJY9ZmeK1KChETpeC0hpVU6UmRIvz/QQHlvkyP79Kj4fOIFKaCZ5/zn5W77K
gcAYYR71OhY+mXTYBVMJ2/ZSVxTr2FuLUTRUA4OCfah9FDoqWPJNUZw4xP88EoRHuSaR2Bc6ZAOk
thWXwrtpgTju0vslVa6JQZn0AYar5ZlvjaAIwnAA9BJc2NxoJ+QS8wKnn/0QmsnfPQtcessRHzzY
9ouIKTQeLU26lSyPbMobj/vtkpNzv84MPdbY9raSPvg8ROehavnq1FeYlm14Pm2ly+Ro957NHIwX
DQBkhI4ro0x22bAIjx6pFh4gbC6BVFX0xfuOOxKc7vXdTSQZV/A6MM09MfoP9qhfjmy5v+F4adUR
Sihk7/NhA3IyerlNIk9C4XJUWlL7/5qHdEL1DcBleYCcvQbdoXJ7AyIL/ERPYPE/u978kWw1rCnL
vimhgY7fT313Ar2Pl2mXR6vm/FFpSBQJbMSpuPvS/0ixgBcH+rgOfXRUp7irKoiUGa2CbB6F1ibC
hUzqYbnqXLm6JcleFK4t95XBcwbke6I/Hc3JEo8bs1c6c/use0zsE1GBWksg08R2nfmwQpbvcW/I
FFRvyq8GOJRYkLOj0kWqHoCyq1f9TVMsOh3KhCNj5COEpoFX6BgaHgJ4Wubtwmyg+Fm5jbyIXXfr
XcKm/+DvoSvJOrCj4Vj52NR1ZWpOQvlGYJXt8TUnQuplD2gubMr4M+nX7IbUdw1LjwiX6G336FH1
5OalzYeYlDsPAIka3nxHSn2TWVwHH9p9ygHt8ssPhtm3NGqvHaP9yfDSQPNpN607QWguNQr0D14Z
WklWOFQ+0F5MH+s0ddhSybobplHb8bL+GhG6KsU3aDpfrUxAn83yDSJrZqCKYsHiVqMQH4Kqbb8E
R3Bo1Ibn/k7+Ys7EISK5oqxDBIuxnoj9bx9Kwv5NjaQ34nYPsCNCOqjuv66sZOSAvpG5+vdNSIpP
Olb4EF1WN7SLnQgDiPr62WwTjgQAJSRpYfkpbI7uphGNNItquBBDbF+4NqhgH5EvazIuskNfD0ld
WrA/HLaK/myn0Gy54h5J2GytBWStwEFQwdxiHNJPyt6M3juYJH5VC0dwXXJuNg4s0MEVHP3LZKp5
RgbtfXxgDu3GxsdD88nnWcZs56n4j+HtzfGHN12MufbVJAsc8BY9BHS190kvoE1PW4u/Oxw7XSrw
NBvJ8ukCnKRBld3C9edIz6r7xa7omYn2cGWVkEvg8LCGcvkeHsubgT5ybRnrDM1nARw1bNed1qnG
mcs2XOPqGRRxl9S9GyGD0I7qkUFo5Ma0H1XC5osLyrGfHFs9aX2CQ7WBVOlJT6DPRGnEhVK7rr7I
QfCEp4u3E/Ppmu0mIJw7bkAiMSLuYshn7l9JWoujCxszdXd6eOSvB708gs/vwU6xp/Cxe09fhAIe
crKzdNufSZ4rV1NfyCJztoNoOPdM50wWb5JPdoKT0OjXhUh3cLgolp3igmgaJpbvZ1DQMMJF1puI
MGlzWlqSddTeJuNenIZGuqbJ2opVAqQkQ08EBnnnaR4F0MiBwZMtalUTaGiuTpVreOPgmFQu4MJ6
nkB0AyelT7AbmrcRwe0EZiaoSarO/5lZ483K8Vq7Lxa7nJcKIvP39n3WbqeXA3L8lus1GP9REoTC
q6n6pl38e4p7y6kwAPKDp+Fs2QAVquzzxG5DDNkYo8BopkyalyAeQdJLiy+uDwHATga3GxCx1sy4
ODvHfX5x8oHH38jdt/Stc8kuAdP8PNQJw7G6qwasdHeC44oGtKw6Wr0SScAEvfoa8FnyfeT+gsR3
LgTciK9GLEYIG/gWAn4QzqQ/s+MUZe+U39ga56vySPipqnShQ6qACjD+8r5p+JszLxG4a5kCcYWW
7qODhJ5M3+K6zajdxssD5aq2D/+VZjx3nulpyPFELtWDLcqc+/XsTQpJaw+YLTBwpyM85pQjVG6M
J3q8ANyCI8cNGYEIG7WW27XNbqo/2wmrX81cDOCyp1q4dIDNgSjLY+tqhdlBpaOHcKuDZw4h0VWu
+l7PQgiXZlCS2mxeywlKjf+GYU7xxkHqcOqZP04hzL86FJsoikpQUiy8dIprJLqLqc0T95+JHtrr
vxYs46MMmbpdL3EuV0vvjUwYjaHd5qjheFeKri4pzETE4fGrXR8EaRsHrQux83hzn+hqFfZQIBhB
6aDyln93kpeqqwPVi7OKeO4rKv7aaaHx+0GbDXTm8BR+AE220zpLYcg3yB9Kub1LdDJa3NwyTTdi
/YX9TcL7WTJQNTcTxEY+OQXQ1Imilfx95jxGjHqQwAcz0t3UDbMbhzB1smO74uXNo+Fu9jYJ+z0D
FH8igMtX7u2bRMQEtfKLFPV4M8zcr2yQ4KHBUN/vW5a1RkqmNWiEpdJ/kNwCAu++R1Qk3tpbN93R
V9hNL9Bxlz3s7Xa4cjUz7cvhSicKP7VC6d7BUhREk4yi9yT7JLeqHiJ34FwgKdfK3beufjafjqAx
ZJJPkZLRXsouxlWzt/VZ7yw6dLsIVOZgsjWTrtvNN2Kco4nZneYnEO5rmEahzO+mkDmzqm0mt347
D3zHsl527lQ+srYIdHXpz349xkeZT+zOvact6269p64Ca80OxO8DXFbK/9qAkJKyZ4uLYV0Ni81d
e5C1VHMEyfw+02rVIAQ7LW2ucZ12iOPfee2z/QqDH+rj+JKJmKmwGy6jZMQN7dDfGVeTqx3CavrR
RUFPfsEIGSQFQxue2A1jU0gneqA32RvSJTH6La/AogLGlGBTJlRNZfxrUrrxWWxj2M+86P2IcuSs
AnTjcXBOki9rJWPmMB/E2Bd9LhPKXYrKDVefUfqN7q6xsLfH/LLR6eXYYRe/oeK5/tgdRRs5/XrW
huGQA1jjcLTeqJah1Xa/KpMJ+kBnUKLqaY7x+tStZoV+VOs50Ngy0lYeGOMDFg6p7XKuJldO53MQ
+jCzdlFTbvnBKJCjQm1HEFq2WXnKPlxzI66jlFI+AZSl0w9G2HOh/2b0J8RjdWIFCpGZzh0QSsV0
/LwYf7w2GUmBVbM/d1f4AmEyfIrpKYQX8gMJudnQ9cF3zRmXBd6H/MDi/9fsO1I41AccjtnbiQHD
dkuYaOVz2aoSmdfJHlp2idmUZ9yMlJ0dsYBelqWT39vgAd1HjUoL5TiXNAZ85K9OICvR6/V7iLEa
wFuKrcdYIWrtJE7iEpvz3sNUSNWjH0uxM016PBqUFuZKDMKN6pLmycfGABwhzUvcSiEtzHEepWIX
9qrtwzYtIxV6OYC4nM458ZBUElUxh2x4bxgOWpwJ6277dwfE5Z+TsqHouIWFBf5kPkmrkytzXWz0
IPs8+uAW1vyycMYSae3OqXULYNwyKozsA9StWjP4JgEUb3sdkH08fGCgm+4l7Uj6H5DqOg4sakqZ
eBWQ+u6hMa3keVNabGA4/av2W7gJXuB9hRdPnYia3rwY6/RVwTwR47iLqNpSsuZu+62G5CPFl0ZX
Wf4RP6k2E5vKS4R1Jnu/g+faa0wI43PqIC0dNnpe4xh6I8QNtBDl7gu2SfZCLo2XeSMZ63IgzRiM
GzPAJrHxSjjSArjuJhINeJH3l+nwERHlzxQdBx59h1abaCPEJNI/g+li01EnDLPn1Ve8OmbxhZuc
XvdgAbtnm3OziR9xh4pmFrP3i9K3R4OgvTKHbVpZOSxpin0xLFHezrRPaAwuZJWQ1tYvzgZuYxfx
brxt6EXNhnjn3vMyOQzSt5juuoTQe1w5peCKgOX/jzYRsFJ8A+7c5x5E1iJaNEEjSU9W2jI/MoLP
dnDhe7XrD876kJfJQiSZCBv6Gr5mErXHEAnmngsvCcxaQZRsjVBEpKxueaiZANOTcBjQy6xcKWe9
LundDAoPh6o8dyHA8BxWtN5V+SPfZaRyhAbk+H9bbn4jXBn/u1KQbcAcGQNuPdGC4Hyk4BTlMQ5O
FWGnuavAiU+OOnf+W2ljPqI8tBVRxgMIpG+2cwoppcBwoUUNofwy+yGkjxFbXV5ikovP3/RJQiQa
BWETPOdE6XzwtZ4F4DA/31FRK1hkICV/Eg9Ue88CQi4WPY66TuyMnA4ksBCCOqncFKnYNumV0+P9
ra+Xplq7WXG+I3z+nlXC1BWXvQwUuMLQjgef3+vQJq/8fEfgEKicjESVT/r9wo2EwLDkD80pkUBl
o+BKJoSltvsZ4pv/WhxZz+MqvgWrXcAaKTqks5WBxHqNbKgWUUBf5enbsvFUF7R0uAH2x7T6433O
rWKnaeM0EgZTJRKqoYgeMBVHTV/QDVzfpxTYtZBauE/xSLrUtCEvSB+Slwp97TqTu0I0wV+dzYVZ
PBl4854lXhcxi4M4noslvVtxLph+mfA470nD8GbuNzKLecC8eNGLdj3FMQdlZJP9HK7h1MYT7Ldg
6Cs8BqBsjKDMqvRcEzEfupEdUnPY6U4wDf9/Q3iT77MHsecrGIPsW79E/djuchhMO/Min4+N1Xlq
mx0p19kmuWg30OYb0N7HOpgnXH9vwUVgy0qAJ1WEX3/7P0KOmSOxUrZfuMz53GpNV237jLwD+QUB
PKrzKsvAA3OjyfgeFhDML/fhGfvxkW2SlYaboEvROGpAmSvuS8LY+80wr71LAoH5qC294Ni3f1uQ
5JZ8TVPhdGxe1zMpCxaRxHRa1WddnXF8m6wlZASVn+yOSyGv4EyxUEo4OQh1K6qtQ3EUtZpU9jaK
SblngJUh4ToooyMba5rtFUqGjkw0kYY00Wd89RIXDccEHhjqtbVpE5yiSaCBiCBzG9Oi3VORyQEA
M3kltCrjoRNRQlk3nal2Kt40IZyyqcWZ5h75LMO57IpmMBdRmdwvsNpNWOxC12X9eaFv+YAL0ZrR
GZh1fWU1nipydnBcZOPHKQInIAGXTLoXUApYyQYeqSGzBeFrAOx+gkJ50cEZJWKFi6yGO7BwZBpa
SkFFMzxW1qcoj3RKscSnJyOOiwkME8UVeAyt+K7uIc7YaCy3zmwcheWmuGV9PuKDVoEdCVHnVg11
Lrbwy+8YFZhIkJuNWpUf9NEkbEtWAwkFkslHQ5xNVOAK9UBioG7UkOsX3J8V/mDVdBcqKnPTU92g
9bZu5d62X4u53TXqGndosw0itJYxmCK60Bel//aQN6qDXn5oSMjhj9sPd8P5a0tPi/MagLjbJwHo
3udegSPl/74ht7jFAgmEpaNVNIszlmj1CoHOC867zTXryFECSfQ14+167T/fr5JT7LWbw4slnsCs
NtAxyPWTxrlVFkA8FANsr+4Zn90yvunuNwxFaGvtla4gdtWzHxAvwAYq0bBD/Cf6yhId641j7lQY
C7Z4vA+24w6LtxZIxVwuWFIQRCxnpbEczgmloKqbCbOat1dp1DEkRZOa94Fyc/M7WdJfCvM8iDUN
wJ/qOe7yTmSG7iA9PJBjkZyz2Ny2umDTXdn2tkZUVgCO7l6zFTEWEgbPSosX5HLDXgY/Ky1dsa0L
ReUVohrzyw12c8GIHGGrKpMWWGjrWtY/w+rPwjiSbfiK1y0zaqHZOmSFWdbFLi9j+f71Ip9lH5bV
M5zPNqwdKG8aU6p4ahHnuspISPkkd64HVF0FXc4sK2cotN3Fouw5EbzakPq8DLvcJQh7fdxQuqNP
iDodyT2ec6iCmjq0V3+SX+My5QGdno1Sf3ZcQc+IuAaBoDt097BptOj0yh8KuTwnhW6LfMlnRI2N
twe7wTOH+VDOrDpB6wLt9pgqrkNTESPP6uj28A3MbMk9rLKYM/qBqY2JXiHZOzQH5tGy78/NE9C2
rhUdyFI0efwA1ZUcnQw9x+scXfF9/+OriHlp1natpg46cTc4MafEknfxauSMJrip1ZuNBL/i2+I3
akVeBks9fhhk8AVOpIXNfkF8CXszzzTEFK/6i1zBLkvgQECu1Q1spQ2KqRSzWSbNAVVu4CLJSIIw
f/0Dc9z81uj3pOBlfyZs2jU5HTI0SB1QneZ57YbzULCs73VJL6kTs9GN0ISJXHFP0ZDh/lkoH+rL
uLOyFWVKxbbJu3ZlCBZrcbL/2VG3RD8KoUAu1pnmKc8p7eGoyjLzkE1UfZeMljaEU1K/DN4hkPpl
+mewVfrMLHyQRlvUCxG7dO8x684OHpfJumaEX+D2gGNzoaAWc8XYE4fOln26/PAodwt3EL8M3FDi
VDjPg2MeL6xl75k0d7A7SKCgdQoEKz6ysnqtSJKNh7ncpy+6/N36nBDywpeHBAvv2tWEahjglNKH
w05GUbSbHbWe2QPcMABMukwCM4GVVSgwBckZ6bfKlxovbSnyum8C89413ObVqqUaZ0AhSzy3uvfT
3jWc3yJFvPrSxWxdih5UUQyWbcR7QI46hrLxlHkZcsSxVWp8qVRePcqgnFOGOHLaovmMkzJTroUd
n3GJBulGcCNR/UlyPT1Y9d8S1XEw08QAEMA5Z6nOSgIHkkMOVcuiNwirRdLfMjEHR26Oxs+dAO/T
VJifc1GreQJQ+lRsNBVaIWtNqtlwnGI6dnYskJTcw54o7BS1tGrOsKd9alyffXxjnHaanjkfjmLo
GLzKBmsafyJVnOhekN+0S43Q5V3KuQJJFPC0OjD0n28Q/KaiRrBNa8oDL13Ae+FlwlUTaCkDh7LG
711a6ry7OnNhat5kx8BMRmrs2JB6HkHOj91NjFyOUb4rZFoQppvrvTyoIYm4tBI7OFqTaZgs/VST
Iy3sSt6Dz0+yovwV97rf0xU6FO7CnppNJHl0FKKfhjpdATt499ZMXS2GjMxa+nJtgviUkEVf+Avd
SI/xm8YXD/Llx3jpthbiK3L0+pXl9aZP58TZmwI9+ue8wcdkcGgqBW82QB1Hy1d2CWWBzz5s/CuE
IR/ogkx29aXM/KQ2zZfUaHTrr5YdcDWSxe429KmYvCGFqViQ0ALpx7sA5v86g1oPHKi2ac6qAz9f
7A+7CHrieiDMaMoY9BfrgnCgv9PpC/jDT443aHgXEbvdN84jMc356uPG53g5eeNqRpBblrna7lUj
4ksGYc2tDCnaqyB7n9ayWtev57cr1KPARmMXL9SMGCs4Te+oklbBJaUBFDV/v1a3eY/ggqLN/VFG
lk6vpMuEJAMwSF2RDo10OB5clOilJcPBWYS6xrjGU2QwDFzCLpzED3I/YNBIZSOf/NhsiFeaPNKh
gj8oKJ9iuTklFmEfMPhIFLmCS37UUmKngj80GgdillhpNt20IC07IpZUSHHKw5JyEce5B3iQtPLw
hK0i1y6V4v7Zzi8PFPWQyu+cQBtapGbfnekldZIZEf7t9zJrqx6Ud3A27A+5J7QmXOc02aGdGXbI
j4kU+ukGjPUIfWNAHU9pOto/kvwavHSGcE1CnSyOh/oNChUFIc7Mky6ILqsK50kX/KdKD1ROh2ez
n7sXEi0f7qOCfA3NX/UQ3r/G60++XslLP5BybWZYw8V9BHhN7wINljnzIc1GvQ13isQrGXNfG21H
+D0b9NJBSp9q/C4HvZ1Ppua2jZgwWt5VJkIrq83VaKU/4UVqp64p9VeInr3ob8S8R5yg2+53rRKl
kGAKV08/WDvgEpDEDJCnhm5plyF8h6VAv9HDWTwPI9HdXCEaYdmHfe3qxAC+PfvuXFaEtaJbPx8z
dJXVchIuVrRfoRXN74Xi0snFaz0TXqC7hxj/Yrovh2XyfK+PxMAKPKRsbyrp2HSd7zmNR8Mt1uEx
KsGIuU1ZorMh2QF8QRQYDkUfJ3E/HmpgDDDKwRpOtKPPctXTUdNgejdHsT+LFYc+QCldC5/3AgHX
Y5jnHgQ+P4bjYhcHlLwjrUheDcQJRliAoqW4UwQ2dDyMqHW7VgFmdjpy67oLx+biFsodV1N04jof
cTFdu9s/rBk4a5GljIthvRSPMYnT/+h8UaRhHEvaICQNa+Qkv4aSgYOVeSCFgQtaWgIqehUMk9vK
5IjDRdJ/sL/smbC5P4NU7Gd6r8OOb702bGTzkhEf372YOGz/K5FV1wQHEopgKiZLLcSrrM8IHROM
cZBFxkwwzNzMNtFX+BdYiYLb3AR1ueinC+6UuldjSKVBO1ZmxTsevFswPTO9058I+zMKGx9/JGJK
aWlfCcfuLJVHc2V3z2Ks1UvJe2q0ORbjh2xMgKDEyGUhGPxA55N714XFtWfk3TBFMVL1v5jrVWQF
U/FcSjAlYTgPnqsIVXAVp06EjBJp/knOu9q9UZs/W7sXVFbnVRpHXhINuVOcFzmhEmpAI7lSPAIz
oY3RDypnHBmYYpOGpYOnuRV/VtX3oKkrAfM2d2nL3/zIDNiM615lwtA/5ykETIdM4//ckeEDkUXn
74mPUQnY6xQAq5UHLHUXBheLSWr1XPjdXSAWlp8ulN0j0n7QurepTh2cCXM7B/AKM/xmRuhUl+M1
OJ3z2rPIbjFdN/0J9hVxI3c2snYD28Q+2Nc1U1nOOvZCv19wUgTRdUcVk4irLQV9u3soTek6hywQ
BEAJ8ZUoVuMglIcsal1rLyEcSnjS3a6aNuIZv7hVmPqbtOHzDpikI/9yV8wK68qX8BD7Uf38hCWJ
RQJFwtNqQ+BcHwlcZpOpZ1FKN0sTCG1UyrBvzckW2JqN4LvAlseJ/CD5z/bgm65GBbZ+s9yXrFU7
yEwn+e+I5zM2e2xYnBNEnHeif+g6J9aF+bjJ0pvB3jlSC6b6WvS1OiZiPuWjosOx0+saTszL01wo
8XBEIUR2kpoO2vsZ89GjOErN6Qf9gwmCS/mmhaYUNiY40/K6a6CaKHe8NoWls990V0+2gugUTRqy
b/wUN8dTccEl9wivWvLEfUVKnrLNva1eq/YB25oUx2D1TJRtgllZ9EPjLu3V+he2XqlOoHahRQxD
dIqa48NJlUrQg5YJ/GZV01DXUZ77XPYWcM8rSPHbRhUb0tRQlWfy02AzmPgM9v5VJfP1TVexLMXg
C+fU/5MjAuOrpausjVLyiJ84Ibuo9jq3keygwAJ+daqP6FaYNZev2COQxIBMamJsT24xL59PpvIg
6qKu7PxhfGhadBjxXuZs250I35WBQwtQlRSXFfAj3IE2UmwrsgFWtn4e77ToeNt4qi+5tOHv/i1x
5m9PM0lhXj5jbccS2tvRDTnZbiMdTK51VWf8VnfRfL6Wmy1mLgZj6Zd9PRyb62nUcufHXomquKoP
cxB4DjLaH+V68e8Uc/iMovJq6SBlfJKHr5UHt06LfNjh78c61/7fWBUzqgeFKfAk0GzuJqlzbxls
g/Ck8DI98UVuqkRcheA8JYdeQTL5yu6uya8H/eBdXKM3agrnW0kn8W70x6qjGSnIjzlQHe/CMiGa
QzW/6s6mudw51QmbtJ0iHbmM14YLpQR/OZ2FWhFYMujZ+BBxJY+64mMVdXZ+yfvbitE38zSF8WdB
EXGtGh1fKOX3CdJTLzdRvu9AtaA67jqCHZ9wzrWIed01ONBpNKvUMJTHjKYG/taJ16kKYR53USr0
q7ZYN30Orh1baALaywjGmMZA8td+xIJBsvCUqBA3NV+0NDVdjOPDDDop8k5GUWkTet5PihxJChwo
rNoEFBc+LHwJK4SYZbLdLcr7Hu9qq+CSmWyfkMUcDkYGpPMjiuW2QPuzDQLTyvInFnrpOrerOpAP
HgFaFEGaZT3Ce1+XXDav/tqOntuOGjlwFRJ5iqpX+EW/tkxTlevTHP3mH30qFlDinc2Phmi9Qbl/
WK4gNPVyYWwwHQwBoVDlmBZ0o+Nj41YyyVd2vz2RsIol2NRMqM6t6EyLIDKHCFaWoddc9vZm2805
VcTQ3ovJO0DWeXPVDD6yhJpabKE2O3Q3AcoQsthd2NLF9tWjS4gOODJDZRSklpg9Of3/pkX+mc2v
sJLeMDx0VY3CRnPxOLFfJzoEBXyJQNJmmyZX7alZW4FKCYSCg5BxNbXRmsYd19Hb/aZLb4/ZaBdh
bsDBhAcotSM/ghEdU9OpgFKnmUv0vnsTMv5zThcImQCC+kMzF8iRMX1RuIPHiAos3Jrm+bncPXk5
9lhhjMvTFTAjTBqRcguMCbv+5CSKARD2EhgBDcEkSdKimUfFxrfInOZO9fe4BV+iVOV/H3/2fKbG
CR4ooYjiu3QXdxmeEXTfxlT/u6/xshppJu4lUa17H2yoUQadtvSNOKAaoD4DiedLi4puGqgtPpKw
WLzaYkLhiF1hkF6lrp6QqSA8qwhFzaXFAWNN5mA0OfeI5FuMl/k7v1ROgousuQvvqjsLTPgQrn+t
WZnt1qVE5j7nPOZrYfmjnlN480Cks8BmiBKhVoYyY1dEKQlMNzBAk5GlfdoqvhpROxtsF+hcfcwf
jXTajTH1eHLursEIcY5D4CdGJ62BA4m91O0smtC5Lgg4HCB7UGA9ItXBV9TbRxWNdPOfT1h7Pt9r
bTjbj6W7+qUjSdyJBhrFh357W4HUkU2ixLT5Ys3CiIxoNX7kN88EQLigf38p1pIBOSzLMy1D2Mi5
PXhTKNd3iCUGgn6IS0lTIZK7y+XZmzbLSPR+SPy1WuEH3CWChvkBpbGrYBRH4Q/QkRiV//zX0LUT
lgmdfr65AXosooiB5hAdvyH5fDPrsRiuT+pOwqb1i4quBv+fRO7BBAGGhA4QXXUpsG/Nqpk/vrWN
Xi6RjpS7dkalf81/TDaCNMXvMJeiXyGtKqH24M/bZhHTd9O7cB9Tm+Ye8IUPkM7y4AgHsdMuThkP
u5XcKR/VFlsRiQOtuuCzQaJRRb9L4TZWTuK6YAdTZscO33FoEow85DynqgKGG3FB8eq4OB9g/A9J
dRgoW2WUCGv6ulMy5OMYD1rOmpbESPtTjGV1f0L83dXLI7XCYcbrr8mvS2PO9zJ8vCSSqL/ub1yd
kh+X+vWWRYaBL35G4gMCC1yfGvsqfmVObduxu7GwNQ5KkUcmO1riFgQ4X+REUQZy41aGFNxVnYbA
DwkMpu1tUotu51BVuWko9v6yZVYWm3naIgrNdQLEOMBsT+H3YKRHugoMoBN6SX9EBCB3Sirw04+3
izqVqxOMcRUK9I4Eprou/Vza5cG4F4xqOT+n/oVpgFS6ZPigPD9PWPhq/VQBuu1srlDjybqcVL/r
65YYrlF/iF88tdCSgnI7aeoFvO/rT/jYkbyC36niJh4iQ/foLZcvWFUNbXnD4MhPx5dvwqda9PX4
9GWTqcqbpc1B3EbvfaprRvxKK6giDQwPdRPOIAqprygPIeZiYrNNheridGUMziNGauLzxvPz+Pz0
EvJFr9TEtZPecrCvlQDZpVxg5yomZsF3WGBNwu2+KP0b0KSy0fmAOfshD8lkz7PEcCpqeSXuUUOK
OplvYKrX6bthtPGF17oXex+UDSE0PXQU4TBQHiGd+zbEHP+JmHmH8LjLgaQxJyTI7xakv895GbAO
eVXU2Hn6Hkjr6WWpJbjhGuyCtZLDQPRxdn+biJi2cDNqAQ3wEqj1eNHmObiB5Z5qDNiZLxbyOROJ
NJNTQc+6KzOoWl5nLbCilUcNsG0lUfIlCV8kcyb2C/wIt2gG4nLdHYk4M+OcywaXvkUrnJVjGQqN
u90zit8Ky6k/g88i08uLMfnSrt/WGG9/L5+xNO+xBD1NrcgF5XvUBKZewiriAVAWrCA81MO+QNRb
v5woq+0qnueV+ZzUBta829B1lXdtOeb+xAxz7wS/HTRfbwVkyqzlH485lhCtcAP4TomsXZNJxe6v
2Y0gYM5PXr0jcqdKjsxQ7M5O4nC/SEBZQuhrXJ3S7LrOT329L6vqbG3Wri30/IptFkFgV9jDjZ9c
3sIL0lCoegnY3biQyHbBhI0Zwa6KN6SIXTbM9s092Qm62F06bb+iLWN5O/qEEeSR46G6L7VebLH8
s/iDtieAmIhtcLYdzTNDqIYLFV4kN5dlw/xiZFLlQfhh6Q5+W7XbmpIMxLXDFYMd8GxFGVYnkT5f
0rR07wscA6OUWj4geVcr96rdH+ktigab0F+8xbCH5U0k9ZzGr+uwIs8qE8R0SHjhSW2Fyl717FO2
k/eANeP30cC391lSFTbHsIEfFUJj7UJovwdYNAEEUEuGtoeMZVJtuuwkytEvvTdKt234gqsO8P3G
/v48V3XOGG7qUXomyDZNGLQoGh0Gh9O7UPjSpxRTv+e3gU/7c4ow2MjWfM9sjqGh3g6GZ6o8r33x
hc2FxYetbIM/8VeGXpSVQtO6tF/J6G7IC/jD93HcRMsPBPCnwUTP++urS0pUZ2lTIcRwDichCD55
hsQdYXDd++MKPETTeIm/CzhfSx+VF9SZUB//PIro1MrOmI9ev0QkNrsfO1n66DCPNCackqeR5HE7
1M1Pqo2dJtcB+y1U/DJDJpdx9L8zgReE1WmPKgmq4ghYQyoJoh9HdttkJnb+mumiy+V9MIxs7OFr
0e+7hofRQbZ9WJWRCnOouHljmCscSXCfpY7cgYxQV7y47kjzoGFJb3tO8DI4m7yB9vBvxrDq0AIK
MH7/AGIy8aRuUkfLSDw3+X8qDtdXUbbt+0hmNuF5zTTfYK1wntHA0LdjifVhq34Sl35JnWY+7hs6
F5P4kOJ2ag70o0emLJKmXL3fnEzbTBhFLZ2ogKri7/finX+xHDGIGYW1vmHtTY4B8AqMIMPvAV3t
IDd+/PA7mTze0mN6qPiQKDkmJ8dkAOWL47r5S8L91IcSiVa8tQXelhNMOZWFM6lIGdPzJ0B3yeLi
TiqJLlmA8XtusVtGSW0XG/C+YUn4OExmXTBu1JkOndCfPrvCfOj59XnwanO8ODniWb6eCETOQmYX
5Z0H6k5dwW045cNhX5i1sVz1HwGbfl0gp1guN7o7F89knohwy/ijVEseejEhD4iAL1UUl0iCSw6e
SpgjncBuSTG8+EdmYu7pMHLKKxMR0dA+lV+jvJXlFy8jYKlsAKJqjErI/OipvCBHOZnr5VyVJH7J
Z6IvWtWDvTsgI/R1XcjQoLmBlwPF1qbQM+p1TQv8qAZoIg4TescUMseo11nX0ebViVXQWFrcVvhk
uKYI49L9D6FCa7y1IkQtGWPxklbg8g9HAoZsnvk8Pw+1+mDaY0cF79Q6Ra/1GzJwGxiLizTg4z8B
nztVAKmT+IpLkNXArXnCToFm7An+rzNuU7u9vWTpEqTMKZhe3wiFxCslQ+GjFqCxDVEPl5pp9vkQ
44V/0rZUKaI+yT9z7GippjD/dVgN1dHTn4fPNwlLpTqfrtCRApoCNrB8H3Q3yMT/DhSKXcGfrFiw
bT8tOMQvL6K96uRfW37npTqyc/Z0TFD41dGrUgnz89rSvWY/E5gr6/6pXySfA7EmU2zT5N7TQ2b6
8aO9pYGaWgLAMcX8F4hxLdVHfmtknufNYmOe2plsXRuxanHXtk3LxO3Hs//QIR9PNsbSZgYdBio5
BnRaURl+p95jt8AJLshHp65zFWT2V3W2q/iO0jb6+xxk2Y41V/nBX4n4fwNtn5vmAJ9mUTkZwacw
x6kz0QXtndb1IrQrd3N/VW9BQoVITWCEMKJa2zBAknPWfllV2a7/iHQGNmsCXJoJSsn6uOCfnDEH
TBxk3w7tjCyQXA/wP0YHQdyMLfewIT5EYdqehjhzGqE3iZMw5lNpRzSqsg4spxFcHNRPU+1ny4IY
TdRSDaebfXi7pJOfibepYS51tbaWEDVTji/elyCSb/PgOUMqW3Yi99T87uiv3kRISSiXwdHyZ/kJ
nalEE/VICq26L1XMFkwGVwivRAVMdmJYoO58VbQlpk1wIW4MkhONDugS8IoxuhiqHWywP+rpw41O
Rm33OVuCV0HwGv2WeJUIInB+Iff7mUpuD3bWFhdbU3QyoVIDYWj28+JH6wr4dlZyLmiulcLjta1i
xk7uXVVsUshucp3zvk4jifoXwBpxOLldDB/Ib64U+tzrS2KKwnj1qkXjzGnSbyRbkrfDvZoHBgFQ
qGjarh7CCWkZlyPEBg4RWta8fSulxa1hDhcXNs3/npst6FzaoUKNFgNnTfncxJ/Z9XeaGgtdI6Bb
SncL4GDqyb1uD/8cLaIiOubLtUpEnL0MxSaqfLxmAzV1y4qTSWO3YYEcy36GpVZNcf6FIHRHs2H5
zfycjdpf0r/1PUJ1Xw+uBSbECLmxa/hrCShHsMl2pfhSWV4jJtnSSKYOU/nC68tibaThYSwcTUe3
H9NLbZxOfjs4Lv/SRY8tKZ2SuItiI28ondyUbd8ICROjcxKW0bIlgQoCEyDtiwwkXhHD/27DksCU
wh1oWQmIWR7000FyjteVClbT092bKOLucrNL8W3rvpDJsDHAvg2Bsqk0E49ioXcdCI5Ffbl/PtuU
0pKcWl5IX40Kt4lTQ/GnO/m42akX2/M9Xu18YZRncDqjvtEI1gxLZqnCySxZ2GJXtM0bgAvEkvXU
CwhdrAFteAgRG8czRZR572ccMNLEboNgDkDV6PhcfMMPxPrbYSqyhlAaOgh9hYs3+iXaNHXngsN0
YCJXhn2wW0Igjzdwo1dZJZajrL7CW7hvMHtddreGeOt4d/MdkygNgQq6lNNmO1YA1WS+OoeglKb7
K6/ry1SjzqSNjoS5HAAtQZ395NjmWcy0vGWtw/k0rKcGdgPY2yLgCBVWuBVNlRh0JBIlQ+kFKupv
vBywPnTsTgvWleCgvf74TEdwsHag1VYKiqJgkArtQM2c2NQ0pPm/iLqoBV9YG+V4En4an5JonqU3
/dXfoXghtJETS59tQRb2rRv0ySMMwsFHq427emqr83GP3zXRFwqhPrlSdVbLC208TR7uYQJYAqGc
riWPgbAIWjUnUhWA2iPTz7H1ouu2lP/P8EntvwfPTfzCFcBsPE8R8MhPmge55Dw7NBr2S+bAvXH1
Mz8v+QR7DZYZrCVG3XbVK32f6ij+4e9oQ2/WnNBJxzZqfyGoHnt5tks15AhGTWOwp2CpoEyl+qUe
4Ov3AXM2fvSjqS6VAtM1OZXImIuSvz2baMFVfLc5FuJCIeXkfG7Gh277nMzSpb13YvtQIT5hazwK
AVlKvaTt/Szk+ofMP9EZenNkVtQF1Z+GC8C+Zle2fD00NcSz93//1+zqrHQ6kQmjU98zJIR1iJdA
qbKnoiYgzPJfI+CSS6Xg/wnct+BJIPaSqi+pCXdedzNAPSFH/iVh8TH6zfx9mLxJJHObPCSUzWLf
ogB5xyzDc2fbdFkDcxvTS2iAzV9bWMMxB23UoR419ZdhiZe5T9PMiIX++JFpWh23rHQ9ISAvbNwp
9W4zkwgIDM0PH/ua2WjkiOq8bz1UzaWTpy6OKZfEvAfScQHmIjGivj9Su2++fDOhlMh3LzlcpMaT
gnuar1daHtVN2wV57Xz21Kb8Mq3JfTcaagiPOtyki4SV1krLk0bRQXV+G21A3F1lDaqrx8P+sQAf
oWVvh3cSYicB2sb33VueLfU2AVM9LsZhICqH4DP2VlpEZ5TcMBIPsvkSCIK1thu/53kTVxv7YjCL
d4QXfWJyLK+nTZcB4Myh4+sZlCsfmZZ2vRwjhu0Opb8c/ZSnyFo7z+/DuW6Gmt+sODYlUqROaIVf
7TCz1N2FsXwaiqtEBKUPq/8t33ES/Soym6VcX5WvHa1C6wBUfY5pUldppJYnKOQhHviM9AtTd02n
fTzPNIGeqdrzvVGAvA3uANtuzLdP5dtSDgiCv81PiT6J7jybsbE/pM4yabGVhuIwhLi8IY2qolDr
/Rs6wwrHUy9uE8Wn5HW2zKtR4/IaZ4wYP4DG7bSohIITrz7YxfeTYtSqT0YMPT9cHzyZcboL0VdG
Y6A1cYyZhBBmlll9aPk1yyYc1nPHXNLvWCGXpbTSHmkeYLK/wXhx6+E3WRcP8+LathW+9onlL91w
ZR+NFTO2vcXYdFYWX6fkEvqmj3A03x8sQRFHPzRm1uviHl6+ccOMi/tobC+8HKrb8kV0xpuqKM4f
XOtYPklhCBlsfTUp6dLytH/A54WORnRhF5rophfHsKaXcS56DV3UZKtIXox60eXvOwoWFa+lKu77
gkxiv62X2epns/Fw5ixs/0smJA1M72Wjs0LdyU2PsxjY5sKbuEZ5N3caK1my5m+4j2IKm6NsGPXP
q8kc225xhg6sVWN7YVL3feMxVq8kUaNHVY6lN0nRvlmNnfkkAeHCXYQ3GrrU1Sdwhg5lch32Vz96
0CEAH+Z6r7pindfjrSBGvs64Tepex00/RScMnrSZ6CWnbzwYqoB12ArUoA463l5hPWNQLM0oKCwP
MCI1itR0MfbKVxCfZ4rJa5zVpv9CWNZQ4pYPhSaAo7s+4a6rjYrGws4FFJDsU/kUzNZxVgYQz3eE
3GBZkbjKVh1n2k07mhbcoeslReN/u2gSLRhC4vGX1etrvBrM9H5GZJqbYIwOyI1/6tR7MCnJiT8h
AAthZ5EwCaNlECq1SqVbaZDJk7aaEHiVouBsfvF0v3is7+ewipd8uEXcOBYUxkuiTEHMZ31gqRAC
F/lksw7NPwc5fu1SOKyK+eubQlslzxFXSpI9psWigRwi//WXCj4y+38bHQsXa61Zh5i0/X/5KnF1
m2R8X9S6TFj2M7QaIAKjiqXNdxvAzNAszQbo+gOcH9fimwmIU+n7A9lre5V4wXpLDXzKFFDy54tg
UgGr1dAW8eDfmNWyy5DwSU24CL0u8kC7xvqfK+zmveiNTobRW2S0o2D9CiwR17D2kUwyAR8YE1o6
VWewCNTrK+Q24wKWkBJZULZ0rbIK5CVHN6J8kd/0QWHRn0jJe5JLX+ue/yFfyELD8vVW+Vt1OsUy
jMfSIRtMeOzfurwdOyHqppQQfzaL3ju1J83R1rUzm3h8hFvHDHitgQs2J/wEqavHrqLTgreyjSBR
EaAU1QOdTqpKXRuiq04XvTs6989AQX2QxonhAtWsEDB/m5JbMTuasSoVf62wDK9hGDv0UZNFP+fE
/ItD81lL+xTnrSUVXH7n5nHcAJlTPsPYChSTD/lUoP+9FkwgxyEXbXAXev8b+Z7NcLE4uCAjXace
zFqPkyXYBcMxzgdeM2fcpZ9iZUxGFXdg/WzRU2upDP+Ttg3pU2skw3kPaGWmOo9uFNxeer4TD0H6
vs6oQXvzLofe8ZoS6Wy64OSwJ9v9hPFLjMHXUdsysUF3+ZaxKAnEUWNYQ6F7GwRGBZXid8mFw0w9
Dj5IevvINjh91YtXrzLomlUR/0xlvMixtEozmEWpU7h0jRvQ2ahMcLXSb6qNGfsEvHpMFSHNWR7z
NANFruKvVQ61BYwACkpc71qMeTroX4KsfdEyHHE9XvUHlCdREZRPLoFFJ3W/STaD5qPhF53Vvz45
LX+E5MgaagUd0CsIs7zUR5detIhDWdKvBZnS6ed5I0jEmqMjNKS1olk5noEwIOTn9Z5dngrV97ci
Oukt/yzBU/fiz4Ap6DETyBslehyw3psKEHurkZ8rjVg6+R0lC7ari41D1Wl83M98L5Pz5f8c1Pmp
uwQ6wwPqNmIJ4AAKJj6UlbSYBSOi3zb7KpeRRCymQNu0syX/jy6XLjicUoNRWTLH0UqztvM8Zhkv
+ek4R6FGH0nxxB/2Jt+1CVuudbdSsrWcEFJq4qyjT5zdRNEaWy6tC8N9nOz/pzrgSctCn+fQWrDz
gmQOWvxq1pOSTnN7tsH94wFbsck8lDBOAwQ4EuKOZyqwDit31pUxmntAGq+CWV2I5stVm8EI3B9m
mwlnUtdg7Aob357hwlus9zkLXVBHHDXLZcn/In8ZPSxiZDJpYqbK01mHIFsXF4pE2jUCF1OAUqPe
hNHa5u8qPimSotLH3teaWuK7jNnSCLYfmQnIhB0VXBq5GE6buMjBxIHvmVc1AwaiGFubPy5pZpsP
ZgfU+/C+zb1MRJLWGgp7wWMmsP5oM4BeUNZATmjCQCVWqy9LVExFvQnggUYqivDE7eMAj8A/WyAq
IuQLQ9OePicyNN3u/baKmEWeuy8Out9VTlPNEfbHd3lClgPklo1Xr+qJrUSbojh+DUd44TvhAlTt
l9+W7JOM1jaNTRtwiYT+An2Qzqqfqn1e2PNlnlCdt+KzWtBpUV1zIH/bn/T41veVdjDb/XEaP8ui
cpG0bedIJ/jAb5FUIp1uOE+2iBNqTxLvbVi96Nu/Ghzo8rJil8L51IajqLGXmQbXjSXUt7GPlyL3
TK3Ss6NesSt+xKyxxL043+h5+uv5LvTEL666qn084hr1NiGP03xyRGUTuDGxW1aFntqF81cLqTwX
IwaZVWE/lVRnW/hKqjTqGBuEaAaE3IPqXICUhFdjlWVKIsNZrZYBaKiMriT3QrYZ7xtGxQA2vLyA
jA6R2b/vlWnjr7BIQsvIysk78pxN28LC4W4lAjY9bZSHyPlNs4I54xUiPtDT9uMT85K9c+pAnuya
hrCK6GnaQHq7AiE3l0KolRpGbXzFEkq1wrIr+jeB4RiR4uaH3uySRZS8jEF3kXwbddSSmbh4HE+6
3LoJ/F6jOo4VozeAGRvIGSn1iLANhPyoBGSqPg1XtcTUBzrJq14QmejB0CnntuFJwWSCkK8pAr53
jcnstd/wrAeCIFSn9wCABpCAbJPQXhbr2UA+Wc9r1v3v7I6quBSMOEz8ndUBAm6NnDTyij+zfwtu
pWBx4kKyWMDY/qA714ZeuqrqDL1GUit/7GEy34Yuxo12gNp580VJAScwLqVyOAzKmGAxiZB+amaP
5jC0AF7PAR4hPnjaXE9Fl8gC5vkabh7YG1zGZfK25JnflsWBAklvFfwkAKNt7nsbr54OVBrtfsp2
pUZm584sMcQ/oTSHJG9wKvA4xRZPSix9F/pwUU/gbkRP5jwAdyw2s0xvnFLCEKl8C/VZcW9kMX2l
tQTSB2Rmvo+7AS+JGqCNAhwrZe9dWTuXHm3E62Ei0G22BF5CmCzJzWxqhMpqW4n7+ujNN6pCGwWZ
aWrgutPc3nY707HgiU1+UFoMeeXSra7Dt8/dsG6jV0b5oLax6obKKWpbNHyPSBJgEXC+SdTEIxFM
EeLqTTP2xE+OusZWbDQ9E2ci9H67bCPyA1rVoA9aRnoFpJIzS24y1B0LBvnC182H2kbsLWrbU7BV
pSBHNwdeXo6UpCtmc0sZTEA0OX5zBIq7wQ/X1UGgLvdgfQRjbUS83OJMme/A3/SPPVvb/uRsUp1U
jbI3rfFeUccJY1yu6OXWWhdAChm3P/8MSnoFMMhBhURK82QUjKmIUlMr0lLHDPs0dDMFSHMKRRAv
Xjzig2u5NuAgRk5cdkTmcaeEynx2PrVDXOJJMi7QJAqIiw8E788taC0CPNLLRhqXNZziyBJj2kai
E2Hmj/GIb3l+dSl11wB3K4d1RC7Gi8yU8xz5um4sZLxSXpFO8RQYctJJQ3G9PjEU5KzCsyfK5iNn
h8Nfq4EwynALr9+zqbneU6WH2yyGe4dSV/HWvM26l76uZfpuGyw0M69GvGS+II2L4J5V619sgAtP
AVZvblm28j/UdD16rJM332xpRg7AFDYmlwddEe84aqe6O1ujfmAUCPcOf+6aF/2ZeJeXTfAgroHN
dv8W0qceRSY1Swm+03YbBJRdJCf0YrA01oxQjf7YOZoReXmIBzaXIX/wQsRQUwwQCttUWf9eM80p
IF4tNHkOkrzSlvOJ8kqILdxB2NwXUSHkQBbO9Szt1FclYjbD/U9YrADiqqdzxgcEfkRktJP2USYW
8Kubwv9yJil49Q42ohj2JUq6FanPHY3VdPZ+GJtHJF266G84DM9pQDgLOlK5hMgaxYaM6jkHLZiz
5ZnlTRUB6fj30T975lMWkc/jSzkqXgXdEiTJDEL9YGg0UT3ah9+kXZ0NNey2ucbuhnj+kqZF0Qkb
zb3CF9SuxoVpYk/EDItTH4+eSCageiX+LFUm2LO1uzfCZSlv0k2XGJ1QOC1irddNn2tCSKNKYl9u
c9aFWlzLzODP7H+EriYwKOwgC9KvbR7Z65d+4G8HR3GdHJx2qEAoR4se8oi1Ndo4i9Ll1cB6CHw+
BgQDBFCRyC8jMic6K/WhM/Yv/s0xsTVP7e8j/NUpYZ8ytjeqT/cme6tAPr73jj+WBF2vuBeJ2dFv
WxL4ADZiim7Bwi+EyeTqLtyR6bzydl4yiNeI/tDAcTeAPlUA8OKYvJ341o4/qWWRaIxLjF0LKzTx
sl7odD5+g1xnM2OvIYyPxu6nqprJHjYI7vS/0RczkJwLn6xzdy2wuWlG0v4lAZ/gOCFYBwaGlZW5
7dq5qFQUbJ7N+caqHzGhkiPlZPx9bzoj7H7ZqddbfQe0lANCg71+g5sE8lN/VtOM7gWvnY/fBtlt
Lbzh+w0ZfUuj4Fu5rnknSjZOAQ3ybwhISbxAr4JywTjkq0LmmNsa8L/y/Yw7OOXmJ94istyG2dsN
EtCXkze/fekmk27EaHVaQ5oiNM68hxZHz5wVw/H0w8vVKrjE430/nVs/FxwVMR+bDB3Dnsy1ryBB
NwQCUD1L7nKg4Ol8Ns9l7sGyyADdhs9D3al5Rgw0pm9ZuAIAzxXwtAFz1S84B72kROGfufssDwsJ
qeDikr9SzHPaFPY6IBr92ibHHkopT5MhcpqttDPFUiM1e4a18Lc1UQMaWIM1MQnNep+7h80XphgJ
hcsewN1FvIVYZKq/9vZ6QR4c7uMSVQHDWzuedLRuqqLwBZf3VNJ+npoPG5C1kqAfHYWcLd0T4dWy
NpR+Du+bfCMAYbweBKUvOU8CIRr+EbgoDHC3KDmH+iZG92DlletoYhD/K8VSz/Iara1OtvZzyJei
tnAs3mf+tv+bSFMPuLY8AWbtRawDyBj7x8Aw9i4W54JFoTsQpTbaRmGllFK5JGrXOBF2usU9rzWS
+r+jwbl/LoJK18D8FjBKsIRwEpchqC1Lzx5dt7LywsZWahekOvYyFWFA2OeiFcA975JUbTDGIiM6
/T9bnTnkebkPdUeKzienANkvYS6xn7pmuBOje7CLGn/rDj95V7x7uF90oXSOxgOLgHkahzaUk2mZ
EYdKDyeUkVpkXh9NfVeU10iYXR2xmN4RpaLgI5mZKaIhBt3UXILSQjQkmb5c6rs35RrhtyvUR1gq
Q817ymF47kb2t1Ig9WQv62clJulrSytSNsyRO3SiGhIa0RlMeFuTI5yfy/fQkMv1ryTokZlqDZPn
71TomhNlt+bLaa47RKHdylYkEOAJnng5PmL94pflgCySdaBf7fNofCmHFxUkWrVnE9hTAoF+K6Mo
ZBZp4adwbtxf/du8iHlKDlwTVRcwqb1KeKYG7mEthK2BTYvizd7nB5RPX+3s+yQb4admvUNUwcRZ
9SPLt5X+eA/Jt0ptWN2uSns6s4ZcExwzVoj2uCNU1qW8y4pKSIlZb5X7cJxN4nUN9mfWy+v0+gQ6
6sthvLIDTwvpZH+oMIR5TI89oo97XOYI97ZmnV9r9hAYApD/+zz+bV4I/zoYu6MzkljnvpEUrOJW
0c47/cEfoTb9GHu1zqbjm7BNnqGl5b5Fmd17oQIjTIslC0DuZx+dx+Cw+gOqvy+yX4KRIwDNzUjD
ZJQuvMMRWSm7Uwr2Df/nRZztC9wOvEE7CxnFNyaz6Yblr1BG9C/grJjSFtCWN6kdf3LS2sUO3Tzf
PFGXTem+aQVGbN1wkqsT5oUrUSkFmxRFDc37/sCFcZjYVXql5KcZbTRXoCHboWIFiJ87fjdP5cfN
qYSfvT29qjS/arnoGFYM0dGiqdCtNs3enGaWKt78mblBPrvRp6+OO67ewLFBmV3KgtYfE/4lTyo9
AhLHIRHRR3gCa/w7E3rmWOy+86fWUZTB0cSsobCamd/eber+91ilmr1tqmF76vGi64m8Jx4pYuP0
ZNXx6/pSWMTJ8HAcr2I9EFE2LtZigLe6TBxkZYALPmcAzNlafxdhdoj97MJRK2DyxfycmM+x+0Ch
+9yohplnOVrQMYxXd+D1Efrt2jQ9WQ6VEw+vp79w4MTlTgXxXv43ZqtleTQhT7ZpV2ElKU1YHlIS
hIoUMWthYGBPp2OIeri8MowRzRpbVf2/rTp0jdmQeziEzKDIa3hA7ADi6ufUTnQA2SZi49IFPx8S
WxTyO2MUOsmSMqg/U0/q72EYN88ac83m+CXi1lDiOatERfYQH0MFbIHH8pLEGVGNrhP3OBMUeVN2
DHYUDroSyj2jQivAUReYtkcJpZWpajSpNDYDk1z0WAdjkrfG7z8cYKK9D1CJFjvBhAQquIk5usKx
RyDn2pu9Gas+wgwBO8Cw3sH9mmUIPEODbsrzRtlpy2icyIhaWyX/xaMnr9HBnXqb2SxkYFg86ZWJ
Wu0kvfhyAKAK69DEakGJy6p9gmSXQ/m5qdCIpOW0ovcsHUM0LzBxutAzd2FHq4oFNffb9TBtnEV2
sbr+BmLxTCtS2Pm0W8OHA/z5n+guAX27yhfMLfGvDuuJzUdSHdgEeoSN0y9Ogp6eNKvfRnGclFF5
kNljbFI2OAWVMvZwkFCoUzLAIbBmGHvf1AFo+uqU6ntx+s0nVdVXCmzKuTT+5VTN2BSIhsUHWFHp
zIdbL971IVJINTq7Dm6Hsa33yP9pvNS+JeOKyq9NwgXCKqD2SHkKXfqKmXqmNWigEFCVdE2uBdXr
JSPIookGoTSjXtSpX+6H700ROUu9DY9WNpwiwLptTjg3Wg8/xnfplNBCcqaZO0sUYcAf4FUC4JPy
MrqxxfFJttjZij2homrmsjNnPuBfP9kTJQcYL5xK5sA5Ugupeu9FWKiWvxBRYb7YR5hoB6q2RRtx
RuMy/ms1rLNbww6OwhdZRaA5dCPuxu9MGi3jCDcZLj1XMXzo5MuRtXs1Yn4Ss9DWaiHfCYtGh/Wi
kbcSii+lpJbd6T6PIIFCzpQspjCWHpvSUaI3buhIQ+uSmJYlJ+QHAgCsewGrskNdymPU16mpldfT
apj1B+lYaup2+xKGYD0b+EUY5O+bRyLIRFgwnGPxRHfhozF+BZaRzYW9gV/1psPooYjEQ7KH1wjZ
M2hqPj36p73CrSe1TqE61wrN3JIgDlEOkbwG+14oidOonCiebsSM1Fme9pBczKQ2wKKNV4tiP/Ox
AqowljE7TWkovg8mbXrLRIUAj0v9kES4RKDHRGFk4DrurblGEJwXsBFkTnGlb/bOBxw1J/HqzVg5
5zluu++TJ1o7bf6CW3Q929BNMN1bst53lyQWIJWFuzzuaLMsfV1wFYkRjPrE9rm8DrzQIoLt4ADH
RoQ7jfLlOv9A09H9dhMNaxmXvO7TG/SEam43RJK6mVmK0AemOUAhJT+22wCMFFRdXc8CsasfAbSJ
gXaFZAQyWkZ7kaGZq+G60uOFPawfYu0k90Q+SZGOJ/JRlLh5Q59hlmcbxSCwToEtJg4I+dYava2e
LIGgxGjytMQ36IJqwY9jxrfGIOTgxOEmphHwvTaDHzB7ecA9xtVXFTJG8rXYcDdkme7Pvi1nyDQ/
cSqVlrNrmbAQhC/XR/Njq7dF2BqxEGRMXhXPnhfkZ61gq+PmvXLoOTSE3TIUNHQKEkzglYEn0dEg
DACYNTexNhvMAe2QNHaTACUJco0I6lK5usQj0IpCXzOmLP8tx3+OE/ttPINGQSj3DsJnp19hBLBN
Qy5SYt/Y+mPNGynXwbZGgkHIDJWgv5M5NFZivTt+3O4qh3gpEAGyYtZ5vN7L9axu/CgDr81Lwg5r
WktVhTp+kUlrenMN+YMTTILZajx8BHGWo9MB2xnvFzepPWNz3wmihKwdI3ekoqbA5ty+BdZQroCR
iRK2yo5STjCACruFwEUTQWEKo1PiJtozSdiLMxJs0qWAK/VYr8kh+pnnmGUXPJxX7AIATfnjDtYt
DgirZ5vCaohrd7V/iIWHK84rXUB0PV+6rDgYtSIPHgenCPqCuGtKc6FpisS1dhqm7t888EgReANq
XfS4I59WmRfpcBOB1EIen1BRgTxkGFRtCV5QiRU3e+mdOb3sGcZDcH1C4SvTdGqwnHEpuUQIpNFG
/ZylNzMYGvi4ZkZlmwepPsGFLVdQKVm2SN/l/CWOB7A3qRZrVMLmxhBCAlKG7S4/X70v2uc8gEQi
PDN7K7mvVp1oDNk/tvVBbameEev98AQ9rcSndOoqngS5YNGqPzDgmRY18mXAp5e7D+OdYj/2NuEe
lD6Sn51G6jY+TJKJT2+Bo4uUbDI49iYtcpegryvz2bamZYsVh1RU31PyU81oUsOqCW4wETaD7t+h
/YnVTwFLZvOgm8igB6Uyz9rIQTd9ZljJT2oKj77aY10z9HX7JiWCBjx8UlsSLzF7VU3zjkjsw5jJ
GUAL+ln6ivUeg1KqfW84HkeoTS3icPSldTt3CFHTDhIsLMfZCTHJiyqTbPlfjn+pJC3YbGJVvhMM
OL9MO1nx5Rbhjdw/GagazcTj9+ZuOXr9B01Nqmjk0aUKPd5MxUpUdPBxNne8jlsv6p1o9TS27Ydg
EUtJ1R0HBEmdKvvkYyK8Wo0JFsaIj3aT2LuUa5nsaK7H6xk7CktGWbFZRZWEovhjlRat+4C5+Gzb
1tu/5bY5xYLVlypb78rbwKgNkHjW0WoCZKtQJ9iS4RQqfVNy654Hg1FC18/WWU0Ul37IOiDkzjYm
73gMDfPVyB7UFS9u1eNYjzrdx1VU/1cbeRvQJUqQd4ybneYihccZ3Ir9V3WInMmJxkDNedfDIt4Z
wOuGiDGgYBnIZvs+qYk7CJncK7m4dawQPqWds3Wi9OXAXx/wX7Qqqp1dMwPGlqBL59pY6x6GzJJf
eff2KAlpN5sXFPzzImkBGGR6w5z/uxrN23phKQHcS2Bil0nJgz/rj8Xl4MTQnRGkFqRSESY0GOAv
/F6lDTyQ/3MvfHfHR3eXW0kPTQJCiGwDkL7GRJcP0X9LeXWwFlZkQMt+pTrXjEa4HAUfYYzlXS+u
fcb5opfaxbxUf12zlGUl09zzpk6ktEsTrBBmtGpQlKKQX5uXari0tH8cdQlIgwCbEZx2ZxzkMwXv
hDnxoZvWptdws3n6zkyNvaaVMx/dlKo25lqpOjZi66hCWPI+ecARnvJoHlRFL2qAdWO9xyXrgLyB
DZp+8osp+u12VyOcpX5CeOOOGLPBgF0Tcq/NJsu5x0yuEUpTdGYSlWXDv99ODT+TOm1bxVhGqvvM
SFwZaGavpiwFliWU6ByiVFtTSQCwm1wlFA9dy079GVGYX1OYiOTNF5EbTdD4As+sKYX0a0a1xfuy
6lO27aANGUUFZ7axEX1IEodsx6G7xSJyap3SYXWeZrP9Cg4haL5o4cbYYvzTHRI0yGX10HBGLtLq
08IbmVNsL0b9OYswY1/fv6eRGdWS2TYZYOoyiwZwzGLz/Rcrb5kqIE7M3wQfAUB7IB0BVkj/6GvA
uQCvp0DWGE/sOocrVPoOtnuJV/8JtigxKM0wL/nNZCNtilchW+J5sKlItxaVfXI7Z98usGfD1Cp2
BvEsP+J377LXyygg3twtR4feODQ99E5UfTi0zFDjYupeyqRNfn/CgFKKyBXyHl/B9RZqRi1Fj5AF
zD0ZsVW14dZMGDRwky4oTFjsEMwRwaVhSER/QLcgRjKf2JN9JgpuYwmT/37PL+a98pL9Y6u8VDsZ
jAqLY0Ri8dg9yadfBJez75YCB6vSpCzVZV6JimFnCon3veZMHEswyXFwdvimInyLL6+ZOjMoR7aL
ops4oLmtsE+v8j6EFNGHFPBSeicFwPT7worwBXuF6WfkPqkYIbEfNlkfM4cRVaDdsuki3soIvABe
HMwU2mkEdWKWIIsWfQqPYGVmF1DVftzXrvGn8CThfUf3+uE3dC9WFz65ez4iOP6rLUa6zQsi65ky
wLxHV/yr6/6UwiSjMMuUtRwn517CLv3i749cOXNu+zpdX8hXRc/EIyCEv+XhqRQD3Ro887gvzrNQ
xPw7KOjKlu5oFG4tOuqa18yRhP0SqhkrsDCn9MtNNU3TlyZ7Abv9JZnmCc4G+YVs7sY3vZJNSK+S
qzxzxbt2iO9aE1CIWYYJzA3HzyWU/u73nOevGMz5pHuk9K0WH7H0fQKr4qdYHvr9FL+0ikMjEgCQ
GQ0fNiMm0FL+3N+NGB+737Bd6DGzSfOT/z1Lq5OHhyxQNrzBYG6F7A276ng5bC2hNG7DQl0eWwnF
CXyvQOBuI3QHW/K4v4mqT1KuFdSbyyta+HRyyIYS5eGtkfvv1Gr9GiDF9vSuC8lPw0xH1JO645BR
u1cFCxc3Az1IDsBM5QoXlizHkLkN0aRTnnHqFBfChmGHRMQAjQcFI6KffJClQl2KBwM+EH2Y2p3r
8GZBxUYm9nt+OgcCctQHmWtDqvFBv2VCSc4rJa3Rul5scsENUAvoiUJfGYpVgiJ44H0gekc9ACYJ
9mFhuRCu7ulzOlTr7xr1l+U/hQn4A3SlhEy5BudDpetbxnurKi74sM2YLJeSSSnOs2jyo76VN0XY
Jbsw2VmbJ2qhR4kxrF2d6v3hOox92PE4i0GzExwSa/RCSrPXR8iFsFoRoavJ/upWlfM+xH+YaRoV
mxx0KEOg2GmjYFDHGHHCyatRFLW6p+MhNZbITpn8iwQe1d5YKxMoYlDyEU4ydZg+7AR487lpDV9g
2vzfHyOoa8gSozuVVf9JWoXAehhvmxSci1cG0s8Yz6gAc3jhQ41XyXAvTrBdEYncQYUSwFAaORxF
nSHDeCOQfc5vWgYE0v9sj6FiWPpqS4fXrt6uoNTVkqYDJBKzC8mrjEaTDdpjiNbStRniecPIX+gH
xbi7Yd8a+QflBDtewU05lTA8PUZUz57d6GHtsKIOoHHTaTXGbBt8q2xEqwSfq8PAAeJmZXj3nDCg
nQCqRB5fdL8PWT1xpp2ClBQbpwPw2lFj028QSAqgUjM6ZM0DNWioN8W6y9/S5uSbBbQmJR8iF0K/
pU+XNBVkDMEN/Gal8jzKieQGX9hkDRgpwCuuhi4GqmFe31ql8CjApH0l2O23pN8CwE6drHiI3l/u
fWQQ8Ai31/Z2uA2VpoPtjUgvn/B7wz/qyHSE+6uOWRnRZLXnaBBF+IrbVm8beW7XyLUHZQH2k4ds
gqGi3tX4vWXypwS6c6kMiBoBDMnrF37ThSqJHjP409/jlw4clqU6GiRyJROr3s64dLz6rzW9uN1Z
SQV67TiEaQxkz2psTKVEneKarYVPWt18SVa4d/qYtgJ9Fdcl9pnemCJqMJVG6UC3VLLyHCWcZ+D2
qT5Z/e3aWlM118iKzKyAHrHGnztGoqF/Oc/wYFz/HwOTAyxyY46d3T+H5aHHUylWE7JM8I6nyRhc
8NqQU+0PGSS7TxZVRYAXW/B67z4b84I/aBwkN1r+ZxOU0mwrJK70eo296Z0Vc68y8/gob0YxZZ06
C7Q0cC4GS0Yl7oiQFMfwbOqyh5fKbUTplHCwBRGdwhFiMKTN+S8kSWUOAeWSmvka7l84nDnvW19W
JCnClel8woi8JQEF0NDGaYlnsGAYxxX4lNhsP1OxQDm8RVK8++dbOt4MIWa6jHl8bk/kYzfgUMwn
/6IjVxI1/0UwGV0dC6WdhjE9WETUvZASkrpPDcgkFoAKpFv0nHc9OyBiOkMMntPmcwgvS3S7A0aq
gIJb9x3JVUmftMhcz2tu1QMhbQAajEc0ZHIXoLYBtSxhy4g1v+3d0FWTDbYPuDzw2xyWor592jxg
JoK4/iXTbk/jmVAmvMVaKyXj/JgPjlGIq/K27CvIg5OkfuAXbjfahpeSnsLfCqvxfYNSH1fqDvtH
le8vQ6dtm0qX15xjcthFWIoTLxFNOKUK7ZQwf9pFdyeJdIY56/b2ZFtI0p8V6xclw9K+nlVPfvDj
aPY00KLyzSXImKnzWgyDrMwWLpJe4dLYt3Oa6Nsf2DiVDCV2xZYIRYEmrlmTEshpiaca883gQU4x
FIcA+nIBUJ120bskAF3ochmNd8Fc9MU5SBlMgPC0ie+3EsvPl0yDAurcyre548qRQYjhd4nNgkNk
apR7Oj1lJypfOV/qm9YqVNGk6p2vwnbm6e4xMyE0NE5dtEx8lLnHYVApMQaT6i/leNPSgwpJuBHZ
KHCsD8XEAmrXH8r8pxBYKod6DvfknS1PgLh/wpeb+Qi9/Qd5d9dYSTOumn8fOMmX8e2AUgC/6vqN
/6nLdZJxEGSLgTcg3rjz5JDIr2/EXADGS8qzVzovt2YSvqI3PaBVDkqKnWcQxPFqHNd4Sx3aRU9m
F83rzuAoxN1zGnaCNJcB2Omv0PPX66rLpYSICdM9S48PFvKU9vwGXlfPF3t3tGU0rDGIvVFXAjDn
mm/JgTrnY24kSwHYi4JcNl4NZAE5Gc0NFl3xGzYE2vdywbYusWQcMceWOMEz9sr1xBa3xDOcCdwZ
hVhMu09OThweEGPfJSNpWfj/pSvZffRev5j4zpSCOUikWsWGC+hgTKj+xHmzWlwfUZzuuIOPVfaP
oWHODDICbAUfQkVcDdQfZLkL3b/+nSPQ9dowqfbZqCdkcriYScACZOFOBtngSTqDMMfVYaiuORuH
KWPhMEUUzQUyMKnuUOVxS9o7/l9lPo/uQfIe5zaJk4esaxMSn0QAtFb2y5vCG+dgfHNf+v4K4ug0
+lui4DfO9nGGWk9r+U6ilOP5Eg3O3RHKHmtwRlNFX+Xx9EPpDayfCw9J43tAam0B2o5O4pgVGcWT
q3XlvIMlYQWOqG0JiHDrHs+sQT2Xhg9mkcKrKZZfq8TTefF6G7p/5qpETBhn6/CUQmmOv5R+yoMa
/kwZ8anKZNocDulpQP0i6ZZBBa+dOoBXEya7/OyLXs9I7xWuNEv5F5zbCADftRVcR4puXsMgD2AN
UC8jkL+AbqGHTGJUlq8HIxOT7ItTyZ5pEo2tY0RzxD2Y2MXuLx+aynlXr9RTPfyn8N1xyCIZp8dr
KJYVwQfRFi/pbRuwXMeACcspF+i2M3TX9edSUyTYJykp7QmHtPnsEwRM3ydgU3YJ+1vq52040WbV
N/vasoDi6fBSzSA0rxy2C3iA4w2XP5Zu64AUA0PsJiKTCgNBHsDcT88Oi8iLmj3nrBfkJk+9qW5J
tl7pdotKp90QI47NQM5CHfc1kBqT/r4oy7CJsyQXEWeW/o5DHeFFUkivnRDMC4HA2n6MM9l7/bKZ
dimNx2Gk8AYN8flZP90BydnUQrtwu6fHIxAs9Spo3gc9i7pTrqFxPg1Fij/a5b/lYYFYdgHyVGQ7
K3r73+Sba5NsHj+OqXNE0wmFymD02/vmM9XnWHZLaM9dI+vuUk2ptvfcllS691ArDD2BhGpCy2oS
WkxCrBsV4C3PYs9tRl91varMpPSYPbumKFJU9kzLLJCMGmC/9OAtUOmyHMXWhV98AmfprrKfztqp
JjoexNn8TTFd7g9Xs3uwBsqLy0E3sxn/Mky/1lw7r9ENG58yHR4HXggqXh3g1F7tmnOOBv41PC6r
fNUAKtufZyuAfn0R7RRpaJQlBh/nApy3OAeoYOCjS9XlsmmPTsfaO9fAAU41Fqvs/muYN7SWHzRW
pYa/DxirhLLRwBBEaCW0IKIUJrEgY5sguWXXl3HTiljfZ7J4dqs06gBmX44etcy+BdZUNeXXZCD+
ongtv5mk+rx8rXED9QmK7UFbDFkFkcIMo7PXucJbqYL493bFNw4J2+7OOhXJE3PjdIr7dbkZ/gkV
RJskACXCAJiduPei0o0dX0eZTt4+YQG5rxevpGjQQctvXD+oJzD7xurlV/3xQVfqmOoEQR/gwAdg
+7USw/VxILustL0QCNtm0Ay+q99IfPo3P6KrwB+vvtzG+SyM5j/GcnUhxEJWSX3tHW+uTfXxZtGx
6Le1iWcTWOuR9eSk18F43hWsoenvBnetpVGEMbVz3gwkBFhJcBM3ji4osWSXdZ1U4+kNk9L+sYN7
AuHSXS6akP4N95HwREoQKVu5wuQZ8JKU9uJJjpCFgMzqaYUdaPoYSJt78UdIOvkAEdgyiuuMrUYW
G7GXTBoUNm1XMKkhfY/wFw4dX4n2mMyx9E52B3ej90WckmAoPHI257KNXdL949cVnkceQWRlqbSa
yB5LbagcaJ/4Q57tk8zTQG8/rcuNeehRMw7wVpCbYCfNiabSffi36EUovXlnW7qBjrEeCjqX1H91
7pcH7TBop1xLH5Qo26E3SR2Qjc9ejHkspzDH3ET+qYBgZkqrPCW+2/YUxheP0TzU4pHVw7grb2Jp
4vS/1TW2/98vhvtBPSqAL5s0pG6hb4Y545Ncvcv3bHg+LELnck4Uwh+YWFm3MfemefTjCfme+xGi
+OHzQaDgRKonnC9eTfMgJzFDO+94f4GaT0jzowJMgII8Oc6BKasZlO1YZbvfgcICQ3dPi12Vpw4X
SJFp+bVP/X7tTibV3gHXrlmc3NvMdejzBNCiuGjdMn3i8g4WSjGTpPo2AaxR1l/0Ds85A31W4aCy
Bj0g5EVV3DVkBuD9tTPQL2qKqIjrl0e9/FZILvnA8bf4bgqcdLwjqth7Clb6rtFju6KZK54Qmhzo
L8FfJz/bq0ydxyDPPyhgy8dLeVGgHUR0b6TMMV3mpouaFhiCV/79ExgZXpYEu0k3LK6Y2eP9AXwD
c97ol2hOV7B0Tbmg94DZS8BQ5cEbpWEpx1cFiVCnALF4lc/py3RgZIsXGnU+JtL0qC4ruATG3NaK
S91ZCvN2C3xlmYRIKg+qJ5hvJ92D2+4M8f/92a6Mvd4wvIINzWiMA4xn+E3DadxGAeRJVZmKyR6z
NdS/v3hG12UeswKtfKq8QjHYlEmS96Ukm72qGQEPNRfbB1mTL0x4ZTyZcz8v5wl4iyiHoODtgjqd
gNYRNzL3p1z6h842kdT8T11LC56KnU3Wp6qaMfxx30PpgZhVR+PtGZH5cKjML9d7KQ2VKXDeG2Eu
kHwNoK7tmomJb21IG3RyT0Gw37WPKQVGMLb0VB+nj5QCMdkIQkVXz3x3A+Lx8uR74UY/qaqGPscP
a9NYLdrkWcIohsbOAJ0lrPuEsZQ+IR+1f1PnfXqLGYZOVGU8/yKVcN1I0UFFKHeHZvXKiiuN8med
iFoGlX/KbV1EZabqrAOIvzrHB57mUxBoNHKsyrpfRAGZa0ifQ3HgWXsEcDKQ9Z14T49FXo9sAl6i
GOLCS+Di1rULwEzj2qFkb5DqJ6+zxvJSGAwMCwdp+TQb7dlQjQivtEIImrsJVBBVUn3MbqwGDh/i
wQSnSuC7zYgVo0OKz7VkbKWKnhx7Bw0e4c0KXGA8Pit1O27bIBZIyvxyPnXY55wQyk3CoWcI1JC3
nA5G7mSuy/+O1v/YaEiZVjipJ6fAgLxs5wELn+PTYK+i5aY+H/L1DFEqaxzSMFfN0GaGCvxapA8d
So71WzvPLQjyNVGDz2SH8WzSr8Q1Sxd5y5mxIzeIageGQrp/S1E4gbMydWwbdpjcKV6fUdYxPn4l
xFMke5jydIO1e9dUf+EkvtoS+fyBV3ihzfJhPu1+VwaO2bdH2mICqPEeS8zBMUX+MxO+Mksre+z0
pjGZ0viITrH8KJ12B4saGWtYu+f3I7JOG0Y5r9lhUxBUaz77I2yimJy60Phsug8cZPNWEajULfn/
LtJgHJgtmynkSeZKRYXSPdBtav/SaHWNz1oYK8orOXkIbmX6CR4yP5gfJLIPO1LcdZRAmMSDgGEW
TZtH4yqBhVHwn237BuXlcvZQmjst4ecGgnCixCySm+VSi2e+ZJFcGSXAMRP37BJ57OnS79pRSKp5
eow8YJFgAgi8NJymZHAeiGQuhuziXi/aYD63S5uq3EEhUGwaGVWAQ+2JmA43uXLW85pfMIZmpNkz
sPgmj55yxOiFzm3RQHzbMgdcjnjUG9QFaTQvy1WCwNa/qv4o6P4n0/8Yq0VWuMhUSdLtuoAf8nCH
Dv0VNuC1zpz69r8W03hIEG7ktm0NNPaQciMP3j0u3eY2xE018fDmvJq8CL2D1zZFNF2ZPh7S+N8f
xG6qBJd3xY27RSN9I9zlu2AEm6KrvHcKH2YLXF2QXq26xFeHzQd8ch+qiT++tHYdH4dG793df0QM
VPylFIdQwuURds5YvWQDz0qGKwTRnvyveZCkZKhsidGBZlc0/EpbHzC71dbB7ixxOLJe6Zh9r88W
FLT1HyAiCJeXqHO5cJ3bHdX/wlzlMulMjRId4Q/Ox3klGjvISgpeoAkJwsLjw/3mtJUrP9p3kmB+
6Vq9snwi8SRpkWbz2DOKPQU7ptmzao3nxffdchJnVm1N8SGvnJQfGDqMCAGfPcS8LaDlZadX8Xrd
+XP87zeRoJXE71m904QkrTtAMKT0FCDi27UJpWQlVLB/33YN+wwfFvG31NOhkJMmNsuPb4Ij2nvX
BbSH7rsUPRIyOXGzVD1QYO5xzmTJ1oMEFUYJA8jMSnXNOtONsbhgCZQeLtVu4LvXjECS4963q5q4
c3hEvD9CQ0OlvUU6lY7Nd4BB22sh9Uppsign+PfzeJuEG+JSeP51sCgaTaWCh3tseFjG2Q78oV7M
2cz9oeQxn8fo8EwXTRJMHD9Sflx0tf4+pufTV9eOmx8pENnHeSgzVOQSSsEKQA2aJJ+RNDi5/GWg
cFWlJ4kp0o0emUZ25sMGLlTn3EqqHJhlzHaiF1gAZHDP5zqNAhE/WgY7+0LbJ3Ro33HL/qxk8+F8
o8EDZCNbai4NLElU1xdqwCgUJ17bnY5sFzLd09zksFLPHVEOrRtSU13yKQmoYkM6TOIC76iVIJPR
Qc1/8f+by80whuAICq9cu2ceeGpL4oQg/TW78FI1Z/aNO4lllZlmJT5JqmSh70wDHdx8UDTyWZtJ
OmoneGpkftOLGYQ3XT2TpZLdexn9SVQpV952Jfhssi+cTWOSXX4+QyBUyVfJvy1wYmHx2YXzA4vk
FfceqppN9ItfHhDykbQT/qGAA/dJKm+6PntaXHmNfqQkQMdWGC5aKNSJA0M75I5WZ5CPFfpxtujK
Zi89kTZukmNQ+F7KmDAtn5mnrKMMlYf47ophUqN6pwo32fur7a7qNYB8VKaJrkHtIaV7sLrpglg+
k/2FGtIPcPanVn8UlRwiLjX2+SRpbpJ0uk6Lhj54YRyMXI+N406bogbUn1R8Asu2riFtZr7M60dV
643Lx2cgZFqTsRBr7ZJgh8IJBCYFLHqwcRl8lU4kCmQvmzE0QDa1qjOuMFxEljBtq4vMIebzSQAM
FblD2TbCQrADLbvllILq5GpiscHBe5pmuTRWOPm+nwPxmQNIrhsbSPD8D9ec/eGAY3xi7XyecAXH
f/OP8jsAVjK/8JhAV0S9VvBfKEKO9EozWpL6xWFSeVXRf0vVFi9B4QUjKHwdShIzDz/gk3ThHHzJ
BJmUcpAZ2CiTWJ4GyURrI5VhHj6uk8TxDaCTKm4zW8B9FlGY0HGQrgYrhCfwpOKsEmvCoDuaUChK
OqkuAqNpH/G3aUzJRXjr70qhz42zEklwRSnG7XQfN7H40K9dTUUHsPBaifVriwDHjpD5JgpypJRF
1jZqE4FGo9AAcjO4DrU7cMKwIDPyovKvyOKF9cYMhdIIv7Kdeh/sLSijoEACKhrOhizpQuX9MOwy
o6hPCN7JhCtqYr3mXprxr9/OAR2Qua6vkcGaQzSTSIpLGZfPgM25m9bmq+km8jkf2aJ6do7+GaX/
PpFbbz56uX5hPWRRitvDU76aKGyu8zIcsSl+chLPfQcqIhhuTdS7brF9Mzexoz2SMUW+w7T7nMQz
xxY5d5Rp3+P91vcZbUuPKpBggactJyTB9V/MTtZ0wj37upoKTnRKhL4VKVKRr2+9UFbCWj5pYwdl
P5v7vrAPmCfC0kj7V4LXlRGgA7CbArx7dZrnuGqUVVDvU8w8bkJmgrWXr9lr7qzEQ7JrLP+xF3Vk
rsTCtX3IkAZ4po20IFv25SHXyGs4fTh6sRaMKNag44zzWbTbkC8Xak+9bEL4yWRigTZ9OZ0yK/0n
sV5hHMQQhkUKCORlhENmehMPGQ1Q18VbF+Bdu1uoFDQr7aSMV4E9iaTzwZOIUUAErQlPwPxhhDyW
8x+ql0KxJK7APo5qPTC2IlZi4lqB1A3ZL4Y2oUQdZImqrtLZBdFCUdkW+Bud/F9jvSIu41d/cgaS
NCMbtDL0JxiHcgPxwPc5ysJxBE9W6PKvhwOJgSpUz9FLIAXCaoY6WUB1iCawVWgQU7CgFxpT4Sil
avw8BDHwUfwXw6HVSmLCK+HYK5bbGxAjp5FtvLVM0qit81zhogXgvD5xzWTIUNGw1gOJw5A9wpuX
sQq7DScoGoRPDwIxREUlcMRmQN85R0X8YbIxzTudHoE5jkH8OaJCbaApMfrqujshda+wcoXDsoGC
kylL6rpoI7RbZmBalaqoz/QAYvKFsspscKZ538uUqONBMGBzmrpt7xfU4fo83IRlqAt2QVCEsTtI
exi1Qs7sp/yGH/FuHkiaK8I2riY7rtcGr/7zS3fyLc0gEUUL1KQPT+3wSG5F/OEnDX/DH7uT7wam
lTDgrWGJr8ZVeXdWUwdypo/BmnWpXTZ+EZ8B4Uh2klubShWvqilq769/6OUYlfsAbqi1tLSu+gzn
x418kbOIpURbYsUaQ1jOampFImPzt5OLaW4yUtu3SixLUChAv60MydGOGW0+I5Wgg82Scd5CiyFN
ROSWonEutPYcTdio2xZvIbuwZQDGSG0SW/Ho6xIbBSIRUgykJL4w8lZiuB2HrWmUZyDGld3F/+ZM
ZQk20AoLqt7ozuDQ6tDz7SKBTC7gD200grVdMIxjYJFNPseI22rJIpD/M3gqhUgNO98WsUv/orWK
jvqZCaqOGnhecZX5yPV/uPxa5r3gpHeYIaykgN+m3CUl4aHRp7A/MsxdLmyO+H4dr6a0QAPxUtBO
6iqRcSOF+l17XbpQI7q0xJyg5z9DIyYr18AagLbIWFCr+nMNRTu2KN1k+PJ1RZmQ5yJqN0p2LOOx
+VzaEGF7Qb9LX1R097xd1kdQr39lCxUzLGy9hdDrejvf+JlSAP+zTk1IuySKqpi9PB/yxOTZ+94x
dbqQdez+R0pyb55bYgVzBlzj2EdiOZo2tLkGyatkMmcymquFmzuHisEUcXsBwR3x8yAKDh4GfV32
h5IE1V/VC/9DY0iQ78Dzd/JNUjnvJZLC92lF03A06+nKqXVvwAexh3GoCLMzSvoHf8k3K/3fkZ9a
YNAKO/zt0MmULMne2qB2WIoVlFbdrzAqsQjyzVDOGsJRW0f8biUUPWTOK+x2dX72FN6M6V2zTnvB
Vr1Ri+00KJxEvv08O3Yy1ex5yjMd/1xLJV+WSHrka9Ut5i4/e85PYXiIuU9nWE+TtZmbG1JeHwwH
RtRsWIj7CrWMkv6HiSC/ePxq0IfxcpnkvwfXNm4r+dKUPWh2eCicT9MaXRAkEQXjOZIhx/okrmu6
A9nQKalSlkCkfMlb1JJtFRo8V47+Oqf4qPSojl+Jx+z98d4tLgo/m1qv6JCQi+B65aX5+fpRf3CZ
aNg2ZGiye5QIr+HQMA2/N0Sh9kjj2zkImywOJQCVkuXtCqjK6ux1oSQqqzDTC1MLO731N8oQ3wka
4eDb2K5dyhzDI6w80lPYkrArnHopZt3sSuWLvC61hRjN7Lz5/kwp4rieG/wJIxUIsD/vD7weJL0Z
VyZi6powXsbXS143qO4E5OgZmhXD2UcvTtaNSKEJBpJPBspKQEV8rp9sEhPINU1xcuJYW3JljuV/
qG5Vq92PIMtmIzCrpBSkyob09Jju3Gl6GEzVzWvHoDQPaKaUuNBEv4+POpoeBStkaaEpQ6QgwPF5
fj32cvQqkR0n2G34FPbI2zRVfqksyXuMDXCDxY31xqn8J1+VcgbT08f5fMlsauhY30DILJbsw0IX
qFo5azNmUKhKOMo2aJBHNOLOpre12d2FVP10BXSTdsiwnGMYB75WdYA5eq34cbfNYjOEzjq0dm+H
h1C3R1dSOuLemrglPCmRrVaxsx0Q7JVYjE/YEY5eWAJ9fsidVRIlYixgJejfQ5CkXC1ZBCTtB5lX
RBBuoOZY/R/QKMbm/QbtQt+rwXXl3p5EzDxRTxnjhHV3zCxuMxnyEAvRja9gCoy4OAJWsJKv1YDY
A0Sp6fsUexLxCQ8c6ISVHsjEh7ry5raQy3GpD6elTkTXqAwyxPLbYI/V/iTaBRSe3lSOI/6HY1Dc
9fNy71CP8IlszpI8KHM3nyoPre48SSvApeUH8pLx3jLP/hA8gis4iRCVGkXMtCAQqjjq6Zp382Mg
p5PFjNsZfOqqvapao7C9S56+iN5SzT1yZJbHoQ9u5d0d8sUqFOcf9qb4P70ap9oMv0284Ijhp+O7
q4UwpXlTGuXsz+N7D8or1fFD45R08YrNatZv0oQ+92yvuO65sVpEDfPomBDtSgnINaOdNIpi3oGx
izIbgzCsFISU8dxABeT74aJzC+XC8fnT5+6wcu6jIcxmBfeHiMljwVsyAY3pcD7MpRuK5bFuxe7s
/T2oqhfMn+BQAZfD9VX42Xn/VWDv2yspkh2XhgLUUjM20ZNH5ZV/1K7h725n0CPDJergy4yif5eT
JW9v6hrXo/O55Cz5DpIRz4sVHPJxat0SQasr5xn2p6Gdmv7CN6LMUI0aKFpEBw896Ol0BWczKjs8
Q6qukIRsCgGw6bcguLAbynWGLRGKVAwBCgk3JEe+sVGdAGxSw8Q/NjCo1fsnITv9u1WuD4/9fo+e
No2zO0PDnVin1Vld33cj1VQlDCilfh4a6Vc6QTXpnImvhDqNoNb1b+MPlZk9T5jKVCdtg03/g0cA
ylPyTUmuJ4G0xJe4dB1nWVNrxIAzkxqTu4nPMYgxaxMxT0WklCu3PJJz5IsNltHBVIh981xsF4ig
pl0AE+T+ZyTiRkeSh52dLC7QInaKL2Cbkbx8tuqeZk0Cr3WSXfwTsm80QghNvmUUgPY0O6sd6Vkn
M6dgP3k1f2R58ICLXK7TBZw5lat/bbN+DQNGETxzKn9qXn/jRnaqRFOL8kZNb2dlpuZ5xKSLLfej
jBJv7KANeRQRSfI2NfXIjAtK7xZfusNc7oUfIjbVqprPRvTagfU2BmYRWYOJ1FFKwQMVFbUhlJuu
gxPaW4G6ArwkeBLz+lJpmEDT7cX39BfJA++aUtI+Ye2EdhyVXS3TZGF6uIsSzeSYvNIzkQMV4EfB
g/gmm+teDQpNQln2d0gZbEbmaAlhi1qM6n5HtlnoqZgVgnwmhMm3k2nwV/NRa2qQCACGFfrIrRbD
5CMHqSDLevHKw3Aveh09RiWz4/b59sN/tYvPojpbrsEb2RXd5aZFLG1AANqldMOxJ1L4TbHsCFax
aQs0uHC1o0IwqwFpEdNwgq9/M9j2j3NVB9hoRVTfD1NnZ9SUsXchL6g2vNsfqktShj0jM8Zqy7dY
cV/KmnKc5bC6VJyB/1lPvqFedN6hdwHjzFNbmcylHSVWLUh3m/SZ+9R9uBtz7wx5zC/3/AZwjakU
BEAnf2iBUxFMT9swYjG+zp34uJcjP+ZkTBPv5ob+Irip5dp62Ii9P1mh4Br6WWBeZHbmAlEP5Dky
R7TnMzaQ5nu5+WP4zOY7eCMDCXwMEgbefY3yIhuZLQRr5ZuVo1kQuowH9wWCdezWtKaL9oik/l+Q
NArVtapvpAzbw/XIfEtQ7yrI2WncK0uxRLvtYpUUsPnShYyCg8hsqdZJBCVfFeC8007W3IWc3Mnj
5uJr9mZyR2hcs+9HaTs96sNK7gKHlGftdo4E26NBtJ7EvXXKPHMwUTd1q8ro1eZlw5nn8/ZlgWcy
XYBArHvg6mh63zTj/UiOjFfzCV6sufqcsEBbvgMmvDL7l2SV6/6Ike0AkB1ybYcRvcdUmWC9WGvf
B5GBwo5ajjixKpGut3xA9IZFnoxNXUR4VvmrVGXU26S9n3ig+p4NvhC+uCOv3k8psL2szoTHpjqK
/pysORom+BJK7Ukqcj3kmxOkneu9rcdLhsyMQWAAX9dNDpfKNiBH6ZvVJ2/VatsOuNtcuPgRlSoL
ayRNeJKiWN91aZRN4MmNPR/DDhFN64Z8GqJj8Qh1dFNis2a6c5sfmHEer4bJZ7i8498+tOiL0bAP
XKXCIGVFlMa9AdpteVLX3vVNeHMFDdRKQa8iPcDn0T6QIqfLSPOx2jrTeMZ5Lyot/eeUBxxmBNlM
anQtiZyKSv7KnNQul1sFoMx3VvWvVcD3uw3anwNhleKRm5whB+EBjObfTh7ZVbPBsOvk7xnW7eBA
YuY43zF986PDfUKqtNm+XAbOqY1odYeZavR0gSSrIfzVRrJphkOkY7SaSXWUnwtjLBDhJ7TTmxms
66tQ62OomXpR8V91qh5yZ4ksMxE06r/THeWNIyQ0ISikcK6UFv5PtbwyaMdGIRmhNACM+uK3VfDG
nOXqND3x7oWaunDpJdDjIJJaMsKUTZgEuAdFu9EI4883KR7DYqV4FLbsofeeEXCNcuRclzr3WffR
gEylO1nTz3wujXEcWXNtHg1srr2Fwv7ZRSiFaf2JuDowSMf11Y13vjDqLL3W6f7fU2PS3SfrBJW/
e1C9TiCKN2+vdQ+y9AQ0Uj9Iclzhh0n/z9A7mGfY7TLp3YZkHZ2IqpOe7J83Z+gOTtzRcbzwTEl+
DOtqxfQnKST5ws6FjShKaqRYJqqnjvN0jYNKZgJTe1gx5lqPF1/e230DTlLG1zCayqIFruldiFae
ogUG844EMWAVPE1k+T9bSS6L6QjcyPjLBFsuAwFk0sTKbPzp0PDWimkyvCL47fKu9d+F2bXgXm2Q
dV6FGT/ZAMUbDdpJVUzUbk7DTNGTRPkXWVMdiOM5CCtnls1jEMK5Ircll/HrRAaELn2+ZOxHLZ7Q
QaOHwQPZ6EIYtRd9CUby0XDG+asepE7YDGrm92LbFe3uBiKw+qQ4RPdT5cXIoHKYkX41eLxLgrVA
uvILy4qWQ6dLc/ObFUT4/9kNJnd+GsQHW8LgcyhhL1sEsx5dI0ZLuuFdz1/09wMRK0gPWV0wrRJa
9k4QkfIZlhokSFca3pIlSWdFeIci3w64KaRPZeqPelMF2j2jUUq1XAXQK0Ewnp/a7TjvaAbkWr7E
VO6yR/KXqiVPTUI+dMmBWzkeJSb5m6+IeCSZ5G5o/j+z/Ysdsk+TxtNZlHilmDx2JCXCJkILk9xS
+QyOEwEQDRep6hTZr86nCBqLjW00q0kLJOgIvi9AQT0hAkNH9xcMrx0DHtAF+AocpreVzEuetQN0
1uXj/kZGgUzc3HNvlJaVBj3V37nk9ejRCFiHY17eBiSbAod+n9xbBM/VYMXPJWN5YWrLW6swCB5Y
+3UlcXp/UjdlWoOgj070YAbBxGeKEj0igeSSUeWNgIRVY6pHi9I3oqAHXy7Z1Fw/3Z5qDZyXAYeh
iVed527FW1g2qbqxqtX5CEdWRc4oYqd0xxFk8Eg7/Bvaj/ZRbijqjINoQ/Z9dc/i217qs+J80f3v
TUu4rHXDXLhqz6NLyTSyf4ilyHq3frFmLlzwznJA3T5E6yquh+OlBTWYqCGEfF7Jv8PegY342nIQ
g1mr6LY/WKCbK7kHT0TbcSujbFjsyXocqVP/2Ow5g7dVsL90TS/r7SV8gawVhcE/t4hiMEZfu5Nc
7ZPcCzEvp48V1J0MTns+PJizgB18di05HTWAaWuZ8bUkCGPuB7gAy9YuLpIrXBHQm2D6T/nyRbYA
lF0bpEls9/+YO+1NYtAU2l6eW9H/XkICSJuXwsF2sz4Scl7MnF8yVRL3tdCSBEbKYFJj7njiIoFD
eY0BFQQwDdEMBoFDLWUxAkcwv1rJAh1D7Ahczv6SCMrYlDNEY0ZL1FPDfVRJVvIEihtMzTIT46tk
EwlX0Vq9GOwvqwYgzIY3tsixO2llHs0mpq3l6LqLiNSWNAKoAlJElNkThozIjRE/nNoQySJUSs0x
3jVrjGFRx1sM7qCvgRz11R8bDfX0xVLsWyiraNH+kcTiGzb59ZOvdPMhz+GiRXiUHU7aDvtUary4
PF3vh32iemkVNOCJ28DpZBPnh8Rc4Xn9W0NQogRSZ8qtubD0a9/agmbTwR6uEfDfDWeNL0y8ohzu
GCAJMdmhvwTAHzO7UYFFP8DPQ3hwiKr8kSvahceUVyutlIPCg8Ts8bXziAUMd45VXDPIvX482VoM
+TX1teb7yVnOjBjMSbihOcUT81CxdUf826Lss49o+4pkiw1Th4PY+eJ9F4YcdqK9BsRLdiVgXJCI
Z9tChpKrrPAvgpjMlGz+2KTPAunzLdZ9Ws319uiD4Tm0Sspeec7uhPww4Zda2gu9uHTdPO229w4r
nnAKfW2XobkYz0m4WO2+NmZWcHIeQH++4xW2+yKB0k9gndJfvLP8zbwI4zpf2R/rzazkBsZFxHT7
L/PunTyvQCt6fOhDxKKKHcXA3Oon1Eyn22/eqIhtTEWXua4YQRtCqlFyP02XXGLAe2dyEFu8Zzbe
kaGAKQkLhlptBNpT0fXAkLb6Zs8nqQ7VO131IOfzTsiEYuREBnFyhd7SgWjfwjszhITNsbgZP6Gk
BB83M0N9agqJC+jbBCMw/tmDCmv2Tm2IX6CEBI7jw4QOBQRofGzrPNVrGSG0GFJFhqPX0ZeKCG3f
+7E86As0D7caq/r1ya95l1qrSF5q7VmGeOM/8WDBXSMz8LXsNy6zHN1aVBiMiatINLzlrIGgqG6i
2iQPK73Qea8Nd9nVqYswdmUE70k/vutGoi1KnHvBoN3ufcUbXGftZ+It5Bi7v7cKaYH66Q7qSsP0
XQiAqm+iAupreLiqjuqPWm12+lxxyOyyXZrF6FJz3AR4JSpxisTVKOZycWFRgBLJMYm+3fJS4R4F
efeF0bN0ikXf7lUzaX9Xpwbw/rzb4bTtO6k9YRDk0im6wNS/2zVobZoDXB3shI/Y2XABVDXSzaiU
wQQEksXbqmsSGxz31H2C6b5tCm9UZMsbAbu6Y7/+KEBQonjLvNHEZW5WrMh9Qkamzqu1Kndo6xRD
cWuh86gagpCRltd0rf1FpInHd6MDspySJ4yGLN5dKR0Pmb+MX/I/8zR0ZTlcWB3KOtnb13ykLRdc
uM9LyErIISmNyhK24He8nzVhtkU6b5BmlPGsOeWCX3gEltSiZnrIxvzFJa+7gq1j1q4eBagep5Cy
2lbNSO6mjvKsEpu3Tqdy3hlX9s9QCZOda1IhegSYK+CAXzjajJ6WAqlMf/HUk+Cv3QQDa1ynX4cv
YHQpYQxFeWLHpqdhYsDDiwpwTZWD3k0O6U0Q+UOtUwEdPztP/DCZyrWNX80fQX9mdWNDDf4ajBjO
MQywshT+mWFyj/gYWvw9h9J7TSo8PZd/6QJcM4ISQwjxUPwaiKAH2wZhXinc+WKq/21lCI3SaBxH
+xYgyKsZNu4pU44LGpm2Yea1MGUce0JQxZWvA/+EgjAD4y3TRgpNwj+XjOfc8HSNpIxSpg017xZ5
NLq4r9oAE/WQ3knTKokN0EBO+8QhPck8X8HqKCJWa4BON5BlCkOeRveMLXCUbXPxRFIINvugL+E4
B6ubR2ET96r5b8zrVyenI3sW6dW0aYwgQIMWGb5wcFQL2+6crRtC4OIl4QiFzOpB1+S7g8ovPqeX
28gV7C+iIVtw3l9iW+KKs4YvAySSLz64XIpdX82xWddf9A1pU8Vopi4b7q1mkpbkKHi4gBg4ETv/
AFa0WORKnNteT0X9XmeYq2UpYDocEGFdrYDQpUSN1LDOD2Nq/HsPGgWtxpMsn+gkOtnn7RVAqPdz
lkL/KuNsjlij7nb+UdbNzOCBh8zLRQ2bdBtpcpcNNsxZkuioR+WT4Qv88sV98E89HJ0Zpmf2cNMl
yk3M0gc1rNppiI5gGMXoQ1mVFa6XgMiXNvz1EsdqV6RLjuqZ10fojrEHunsElxX8YcXHVdCPwHZo
MkM73r7YErj0f5kjNNf5EV+DmR725oWQzP5KAH970FgMgthXSOtF1FIXJAUPE7FByDvp54C3rf3E
CQZHkKm1WKFpk/zN+asJo5GOIxYxXsjFW2Hgjy2bY0TtBgP0FUH/TA2vBfp5TQTFWGtHOLBd6KWD
ZePqdGE2lloZCS0Bye4GvNgDlVzfdQN1AJZQg6R9AJPWSZgst2t8zGHJSU/yL2CguZ8CTId2Ov3P
Bkr1tmvbRjd+WcodYqGRWu5svI6EOx3O30jlNoyLpSKkxfqNrjqP1W+YbNB0L3GXmLcSRBK+3ZrQ
Q6nBjBebRc/YfIeevEpKwB9nWmHoOWpRwcysu/bvy0Tpnj1JbFFSo+GxnWi+d+GisMJeO20Byjtz
PvP8R+vofDGcz+bwGQIfifBbsnc+BsqGY0v8gvg3HqsR1RI7z0+YDNOwR7reIkQ3MOEk757DZJIy
PcqEu/YMmsvucAadZxGWd5w4ghVrPusaEIqrWPlTTpsOQm72+8Ybvgluefiw9rGD3moIFGroVusZ
BLWD2YSc7W+dtMweqNI/Ks7ftV05jKC0K/DlP5JOt4Z24gXFnvHN0HewzsJR64+gIlHaHL3vx0nZ
4hd0lA5/81256tcyT783Oola00+R6xMTnRXFfo21t8yVZlXD0R+3hgn+zkdJ/3AmZ1reO0UbqxPh
bL8fiGZcJbTX8WdSBCh8RHbOjBntfOmVrgOejW2DHWgweSvQPuUmoNdVqthuo1JRx9tHz0jhdSLb
vcRVbaA/77Iy/5ED+69PPQM/GZTCrNwRRGUoHSW8YNZQf4IhEnj63GD3CxSi2a7GbLcCe98RPhH7
r4oOJ94Cd9QaSmlc+dXbtpmG7ajgp230GvOD+GY/95P65fE2Suuw44kMkyUUAr4XP988YLNwx41V
MSHm8A1YlVjmgQ7ryDlVtGbpYr4YEhmsbpOd9m7bsuHFZCDn6wDOreSPacb4DEn+GsPMpjkxk2+Y
gENR0OkiI+8IjEWFYlpyPZMzzqwzd1lABx6uDbWa1A9wxpgwcVfu8Hg0Js9xToYZF1RBM5fEwx9K
UL/8dqoy1CijwJ+odd1/su0JGNjH5ex82cxYlzOs9aGIlBzG+XPrMA/QASP0+R3hLFfo6ljG3P4g
vhYidfc6BMw2RxfKUC07luyexQm89MCTkZazOrZBgcVM9AgFsWOmFX0gLg5NB6Ac1F1y2iR/xbaa
wu2uddnp66YX+wztqndPbhhOD2fZ55lo/HjAjcVywHUVWhe1j4ozzlOWR3HAG/kakFS+w2EFshoC
dlZuLzG4ZHjGFBP1H5pGQ7tlzC32LAw4Gw2wplFYzRI9fIo28Qj/o2r3hN7H7XJg4ZJhvTjky38X
2e0t3r9EFBNNzAOE1kgPg0pZUErM/bulYGr/z6UBBH+PooxHRy7cpf+ixFY2UA8AKayULyHVU6XO
gURZiffvhfi7wZ/HltSIhy1u4DSKz9a8CmNDUskhuhIsNVJDVgK5BVbaancx7e78kZVU0ZkaKEII
Q+GviEHJNd3t8HNABrd2ZHXj2Pm91Sgnwf76AR8FXtZbKEWXTDaGzdfejoBL6tyogzq7BvRInarY
/f/9779D9OX6naCxce6yN2qkXxKHtRWEtH+bpFG4k5Xh0I4j1p/m5GCExC+5SYyycG1/Sa7cUCIG
THDceBFSSSvzjoeqff8bO2U9H7/zzGD9SgXXci5oL3ILiX8jxcNYzQaLc6bwFWZKYqDRx77VVcuH
a/K5KCth6LyHWvR8rRjTdtPj8EYzPyhb2NWERsPDL1PGjSGdwHZj0tcuXyfoCOClk4NCEt3jWVpD
4E9E5ktBzqK38I2kXEsuiIQIXf2/EQSvASkltWv3ODKzxiKjUVEWGpvwF2dA2UpZ3kmJ3OR0PZYv
W+dPnwxMHf0JhYA6nNBC+UjkQOpp19P1yuRuLYHGkXyJAJh5ygdl1UCbRQfi7s3cxtG1Pd858huO
jE+c7oYbXBcgGS81EDoJnT+BlrCLmroLv0IqN62Dci/q+Sotk1yLv1iUwOohOLxD33YGr2ZxVKhp
4asFKJTF5Io4xrp0W4zAfrSmHRoy87aLsjRE80ErHUz7A0+wzpj9e9lOHIg4u3CbAeYLapOOfVb0
b4/5D5qyJQTiWcdc9P5gCidtlWgwjS5s8PgfOfCi9CJXRSqBb4F+uaHHJD0KpbxLUW9QJ4upBHcp
PXJFlj3V+THlJjTUAuzRj+1Gtda3Dk2Wl5XEmbBubXTrA7DYjxW75h9WIdHbg+eyIMgnhSiM5Pxa
sPJzSFqSOtfgmsWN+jH1k7LZ4MxKjXB+nSg+IvNUMbUqt0PzehrNTqWPTNxD2Bjn1dGF66U2daac
Dtwv6YAHHKZcGHJPLnZJkHVYwl1kr/IPNOitxlUcek7WMHa0AHyhaF+eDZgN69qpW0gqJFCIHRqU
aHPFZoBeKpIHDfz8ZiGSAFsfCQJ9CRrb4196X1x42htuQqYnaTcl8KKZEbYug3Gk4IO8JVqu8mpn
ZjLOXLABY9YBdC4zuPsTpucF/QMZOniQiHdFsNJYVrr/0Hd6RrTSm0qAWeGmGg/DXOtn2vcxVrMo
I1EGb6TAQqEZB1KXTulGflTzXAUPF3H+kaqRb3hGNKscmU643+Ylb+gV74qCelbiqvGSSz9NIyJl
DedQWQs222qx+8nGm/b1fPRBQpcRuulztJXuAhTfxDg07Zm009FGDaFxgaBoYcrUxsiGoP6/2Pt4
zlaUVVUQvzrNIILbmfumvUyONEB2QhZEvaTG336n48oE6VZGoDxnxYODR2sTbraO3x0cGGQiD4KT
Lm397jL/5JY8B4o/Z9GnlFRp5qxw1WzvzTee0Ek5K8OjD1ZOVeYTPDzTuXnMvOeAtCsGAFt49NQL
EvXFlgw/u9xu0ciQHXdzbyofOGIR7FCbeb6c7zNOw02B0t1nhrPXzfv/p3b+R8ndxqSRxT8jiLB9
9HXlW4DikYbAW7bIRwy2duAiUrmUDx5IBnn1LQWCWTU6+OBZ9Rzb4dTHzaSoZP9f9Ebj+NzgYC17
08H22MDgTH9T3gW3ugM8Na5S6HmAMnj5ctcwoy3opNq0zsH1wrjI6gM2t0yRY3rO1sn9NNKbo72Y
t6w++RiMXEwk2G6TrrzF/SWNkfLEQEHwEgeXAWcTt0iMYfMSNR9+tnUiGCu+egLyNeTDdTWAjtq2
n6oDirlbHujblAaKdCenBy3bSOckB5lX21v0Bafl5eEHAhB94l0t3gsccVRG9oLAEWVKce5z8lfa
XHERKexDykas5HGR5yA/ANeTK8HSjGrAcIggr1zoasEcbYW7Zrfa2SIXcykwCDPyXYRtHAA7FkBc
lLVZtAFiBFt5+J+16pbfi/kUFfjv1LJrB6uI0gme1IJd0R6WhXlVWslfCBQXVM9OWxRbDnEvbRoB
2ZN+MAegU8xq4AuwaTf768Vu7DRXGqbQkqBOZUPOzW9CTY12WYNX6idRR0AJu2a044lkCVDB9Z5W
DVCgxQ4jGXlhLpeyfR2YOvybTaCnzSgQpYmWyNQ4MyemBy2VUD/eHeFPWZxWxWAcKZp/5MThS6w4
jP/9LdLdsOIuwdKTIWf/yFkNfsIVnD+sItqTFbxMDLHJhHmxTALzeJcIpJ3T43zLH1L1BrpfpH2U
ZQ+aCg32LVubokUlvlCZvda1sxUbinH32W0yfZW1uF568FYOwen3L7EoWKlB5VSHRGpoV3SJREOY
R3uQWoOT9wwAxt0gxQnt4YH4vhd8g8+Zj/JnC0JZplLLt5m9oG2sE8lM/29rXn7viNqp54E01IaY
856Gu2DOjlLehh3s6G7a2mdww0/wIk0hmrkAMb9H3qoni18LA9WivwqW6Ro+MWAz3ieJVSEmVgCm
ijBgDrJ2iWiHLObxncLLMUAatD8w1K+L4pGjLgVlxrWuSv+U9qenMwBD9czwEjVZ30lju6NLHdYo
II4ywx6kFuqbscpkRzwj51dG79/uSIkvxlPayqSSM2Oi02YuTay/7ASrHlxKw30KFZNfTqKSeN7/
6yH3S4Zus2xbl7sKJYEaubVCQEK+pfP+/GP6NzBV8U65AHtc7SaAyDnvhcO/4xSuq4GteGBwrWQi
cPAqLNy1c9ZarcpAnNgnpddVWbf0CHj2AF0/mwXMwefWj5B1oyybN2AnpHW/ZpUdAVwxbJqgiS+K
dp+c9Pf7oMlHH4JYlEJUVUtiPtfAo9ne2t1C7V7IevmWLr/Uj7hEU89iEKh5eOe6BpuWUAunN12b
2jmB+A3dxMyR7/yk4JOUjp2IhQ5zN0v9pWcnguAncDnbz/NkVl20mYg0Glcqm+ShlIrZK8LchJEK
eREiflRHEXHKGkyoteavi63tCVKhEV4UqPQNucFrFsjy/MXvnUT+cYgojg5q9uQ7ma/sL9smdOvT
WW77qQjnNsCuud83TgOk8pQ+ohSdTYjcuaPAuWtVparIR84gYx552DYr/3O9BFwO7cIU+4GQGfUL
0JIIFeiIm+eyXS6PFk/7lJYPxj8tKBU6htpZiD1r54RThiN1Jxn4hPCrQxqNwyBXB80cs47Zgx67
qRLPROBi73ow7DWSyv/3RPXk+LaMiRlqiEUdUYOvmq+WCPwaZ9PHTJxYd6K5XnTHXqgcJ6ddgxuE
FE9NqWnFXudcEj1SXDsC9LIIBDuxP6qfP9vPj7AKuazvYRA6XlC+xKQiflXla/uAwk3JiNblZ32X
PPouoE525rKpjzq2cNVflet+aN7TL7dydjuulc/S+yqK1gCjcotmeY3/M33exX4vgaIJpe/XY5MS
52azgvSvnGsnHBq85X9xl77wOuZVCjUK0YapoJhsuG/s+zQefOd1CE5uNzPeS0BatJDyRjtfPYiC
7j/FDI7wVnvrPjfuM+gJxsnG7O8Bdm/qI8Zc8rJBVgzxQCwQ4JSE+5Hhd36e3fKGO0+obeIwo4RX
dLIDBCud2u0tOkmx9x0/1DFWGjyVYpqKPUfQXWKhwxmD/zyvxcc+MIAlXOvcF04oPf5Iyt4fh4nU
7WuFQG7LRSaYDCF0VCgTiYCNdWDg57KeASnW13o/jIG49q7Z7vh68LsSn1bGdLxZoMd8j+2Mzs2h
pMSAc5UyB2t4dcqWKl/CDVbo8dp3/Rp7QsBD1cKJLd8cEOGTDIPTzEOJ4Cs2VbE85GKFFscL1RYc
hWi5cX8iim2HlDdTSW2uWze0DFOOodTKbzvVfWQrgqdbJk/6M9dgpAM9qboDwAAXqYO4mtKM8OjA
1ja/YbhnB+jgeoWz5KZKyrQ0WiBCfOuJoQ/161X8Ax/It8DTHmeaz8iubU0jRA83u9YKoatB4Q5d
rFZ0Ot/rNjTjkhwH84v00Y8m7SikAq5hgIFGKo2ynAiJspV4JzKD6HSOFXXPm910mPaYJ2YZ2RTE
WgWZjY2/313oXLap5VmNiElMqfXLqQoA10SUFLbh7tj9NNfXx80Xr06f2ogk8zbz3EZOIj+FDKrC
Zfh1chWF829RgCsRax2YUMVec8w8b3Ye7PEv3hCsaTrMDPQKfdwERDM6y/NoIa8fMyqp1jLJ1zxl
R8WZOeUgxuIxmKyticEXwslMsOcWxdRBX4nVHNJiNnBQhmz2Y3FATKWbV7ncsFWZWG0lmj34K3A/
JV8sAue0I1S09FSXSJdFFh9H4flWosggv6vDng5kG80p3C5c6LnZPsZEFyh8bDkYLHyxbV+iRbkp
9ME7+MAtbmcJZz1jf77/62uQYARziC2SxkJrPZJeBxrlQV7D2A609WI0WuGDXgNs9lVxPWqHHtYW
U8xgfhywBfOzWWJ3Bg1OFx65VKCFh0HvkFAC3Pas4KncOp91rEQaYYw45REP0Eytm7WJt2QY+fw5
IrslYndYDFlr5ns0Ur0mKodk0iHECOnQ/riaYHCY1y9WkPgsGUyxCo4NtiRfjszKxHctiRDUImxc
LDdkIPOxGggpR+jb5Wv/02oQSETVEc8l9Dr3t3EGw+k0+t5e1C8jjFNPJfK9TAfH0W+aubxFZzHv
p15B4Loz22KFb6mTNo7lex90NnlHusJw9hmHhWECgJdW9A+2ZEa46zL/EMp17sQvtnO83tBZkJCs
/u2SnTyNQu8T9lbVjIcmDda36Ul+fCSAsRTTX3YakV9DbxjwrNUyvIEc+jOcl1cQBz70aROHQuSS
TBMj8ELpn3ByOTQccqUGs6DdUveyQ6OQxZyAlOcnFRE+RFy5uu/RzhaxichMR4NtKj29pshhRRRX
vMJpu8uNs6v3bVNGdGqJr+bILNNJK15OIId3nEC9QMzJoyl3PFBsRxxNs0SF3lKLc7YVV1vIpu77
6gVFVocxvpPtPXygq+rExNZ+RdlifDSEnjwvEZgOyET8H6DZSbQ/O4urKe+6UeEpWuaIRMVysrIn
H6vx7DZBrUIOZ0hIhiVcDFOY0UOKS30O8/v1MKI7N2dHindV5cZdbxs2NEINbZBE/PrCaGI/REb5
CaeZgvUXbBgh8o/IKM2/bFu9tBiPIqdijCgjYmDnfQCPQfu33tL3Il/mzHBj1TaQkAHPLytdRvg8
HX+Sab+jWdWJ/D3JES+ENXDmS6XE4nL/MhiwfIBYZ5PULjZTKQLIV2FNzLtZniwi2EbwdBf15Ofh
6rTEf79QxV4BhSTo8z/6hh+VQ4iyvNXjOPLJJnDs0dXrFn7u2+hWewpDxqXHLa9dwAIuiVeobXL6
9Q6pnHwg+GES2BfPjq+DvxshvrHbDCTvIgbYrmpJBwZZvEheofF2ogjFfb5sxHcQjyUuK8+MF6h0
/7Tw6jbtMX77GuGjjdu2npk9e336d0nj88mivXG1VEdHfAKbYQrILqXn6vCnPH6I3KDHjFc+6ZBd
uOr463BRdB/hrkKPC6v8nVHRDdjz8bePgzzXVjtxH6PPFHZJmCYyRoqFn+BeDSsV1kR6DrUh6fFX
7oiTf3n0ZICSY/VpuvPqEC1E46GO453jnZbahIQeU5q+XJLqtzdyc1MO+0gcnccqMmhDtdP/MPtf
YYjHhTh7+rc71bOeIEbIkHJXYcT8gCGsmFyQC4+thgk3EvG2met5FWjcEam4yGjcRHhuJRY/Jms2
LGoHGPDOjqrxCUtcSz/yvKNCSI4mk3o1Swsx5fNG8NmQK3fpZdNUeCLCmkJrAsATFdFdL5s7NaHT
U89aqLD9rnlJGHBHyhRQc2WmRbahse/KWWXMVBLOlfKRTWCb7xeLJZXonccNx3xdXpgV2dIWXhDc
8KnODJTP1T4XoR44Utpat1+PEQ8yvTWs/tYrpjCnxdQo97sw8UJjoWb7xCb2v6DsgUMxlXXYfBJd
0IY2hJJgt5BKSElUUuYyn2FGgeUkN9bxd8ai33307l6DgtyQHnGBrC3YF1KH5XOsIPmgi/cZFpxR
mrzXS+PA5/lkqF5I+CiawZuluYs1gmNJ4duHoz2VPXSZqm8yTVtex/iqLIPvHMvO7SsPd5T5GdfW
V8DSKD/UOZS8Ul6EhJ2wun1J+0ZN3seI8fhbMpmAcx8gpxSDvyX4RZYVmsudQg9l8WbMW8z/DvxY
MzxspmoYB1Wn2ouv3TxWeTnolTLJWSkndS8BMFl8ZsgEuQbFOkyMs98VZLQgVivd75XgxcDbabdC
ip90+6WbB0mWYom4qI79hokLc1Wnlw7m+POMJKRb6gbyFdF8W2S/1KWUQHZIxSECq7q5ayI5yHHt
iBKRp06KXF+EGolqPXLshNdcU/5ZTTSQV0Cq/K103OicA0VoSN1SU+7HvOaTlfVp/IWMjYli0oq1
uKcZhB/sBgrYOyXySX69KDD5ooxZ8zQXO5NkUkj0GExjsxffPCfnom0+1OTZ6Aa9foIWkX5bj86C
GLr6SwWt6UroYDDkqJVIik0haYZhIrOACeCZAWA1Vz7DAOPbA01n2pfADZRGiMXZKM4CeYzqxSYk
KVOysRAPbYRm47BJzLMfDLktv6QSUOuOvImBSxlymKXaFd9WvNDFwIyAVsUcrNYzrIZ+TjF7nssL
ZAYjX2455txJwmbBBnebt9kAvIN+wE2RKE4VBDXCn+rEtIGc1tPxMUwLFEkDsL/4QoXTI7l28hqe
s6hbfVz0VpEDoUiKn/jd5gcAKCIoC0DKHc5NawFUcsMTA0Y/pkKtzgKTVnZU6AY4x6TnI5k6HJQ8
J2Ygmct2Uag0Det4vHruDsNXHRDS404mrOK9A1e62VAACXhm3o+v7cfjIdPfuD5iAox+sgraSqDj
M2xR6amwAFKW6p4p/TKWxNYjfU6qMD48dpmyMvzZV/RM6qb05Qh/aPylNbbsTUzUzgjASQIuuuB8
6Ca5O3ABfCunROxs/uXLud9mkHv7r5F8dKU8fWBLISlhzT+3YzhAS5tNhzzQGzezzefjX2O7iXIH
Nus8Bk0sZoA7iywntL9f8hZP2MccHX2/0md5BEDqOyqzCZbGV+0JA3Nd+bGZzNef766jYTR9D1NU
6P1tO097Z2EGzy6jSVpk84VIJRza9w2wlWvzJzF6eZUlHT8SRQzj+Vg4nAdxLQ8u7ucwVujorUWU
gzZ8iQxLixhNUIyISq6ZUF9SrGIASJ4CHN1kROWo+a4I/g0J7bRJTOFbDNweIWuj+KMI9skbfkOr
2Nk80muNhxrXnhYXfrLbCl7Bt4egZyF8RPLv9py/ENrjXOifpgF0iN8/qCXe5nvyGTX+DAZGKXuL
PBMIypnpv9BeQRYjujbbob+5+kUuvdR90SJx6yM1KgHIxV1Z3FN7b1CgVzdvlhgybNl/MK1DPkcV
889XkQNzIiV791PaWAE7bDixVSg/1G1A64doYyNBxJ/XgjX5m+sVW4zfljmf30I+J1KnMBieFMSn
Sd1z5Ye8CizY2qNAY45+MwSUJqsal0/zI+6uHb9qG+vTlpSLYKnCpjgVnpPhGGaELDr1y0v/8tOq
25cekBBSJiufXW4x3C9/VSMWqAVlCGXQ59lhZX8t2jpyb4EoOEpjGVXvS8LLvjRJmMJ2P2Fzab4p
Wd3jc5giLJ/VuiNKPmMtBsn2OOSFYLWgTLrjQEbIs2E2k6YQM1ZkoFPkSDpHdamDql+GkWQ0xhmu
+XmJ9BvehOLIr32QV/W1ilkut3d97wlj+m3iaDCVSi6G35yfJS63yLhX1ToWt7z2KB1eOJGAeivW
WBkafxziUVVorTv+SyOAp69Dk9PNlGHDayH8uYcZeAN5xT4bSwfIBNouJddhSKfBlLRxANaX64tz
ANtlBm3iK85BVGofClVzrdj12jtuyIAtzuwCdEijxSb1VmYSQsUjm0RQFGX+GLloLOxXDpZMDLjw
PzGf9c15icmsCTHTljnycnuiDb112YDA5E05lzjyKdHCpJ2IdQToBl7zMoSmnFuP39Fc69Ya5GPK
UqJpyqvXYHwhm28ZjgTwtUOyine0SK39xCCIujQhfhN3OXboNmLycykZJmvtZI4M/4A34mpFEPk4
1+Pu1mD3VUxQkrVDBw7Gv6AJT0AAd4Yl2utta0304W032piakhO0d+3nkGp3KQNvOQYZk9PobFyW
2nWGadw8V6fcCYnbQ6MTU/Z1WHmOTpkwl9xwP1G9fNJVQfUCsDr739WBSwbWfqVhCOuShAbE/Ljo
wHBFcD0GXDdPF+eCwfK/02oYt8W+Mly4OW+AdTUWVC+GPPu4gAJH5ffga7ZdGqf9b1W4vNovdPLB
T0zmd6XCY836hEzglYMCNJFLDrrJ5fSVZ3UUL0WI20F6MrkHOITaITCnrqWn21uRhitwar58wF6m
K1qmTE9VKK+knQIcSxaVu6IyyQoH1gxXVIme/sYVg80b1WDTiPz/Cs7Oznppc/aVH9bYJnUZxlzY
zuzRdWptHnuCyd2I4MwT9cbd56PZVGB8Bl9jwCcpKfIPjMa/f0mPg1dLfchHJ8yC8VwBRAq4qtuH
1Y98o9tmzkux+6O2MsV6H3Va009tnTtcd/aRPNDQtGahP4O5VSxmYaPsr95aW3U39YmJtHzlT1oU
c5Fsa7LlCM99WZ8KthSm2xe1YyuJkMnvnE+69iSSWu40W8kKyXi+o31A+60GrjCzYHbVEXr9ZTMa
5thajMgpIrtWYz3bOAuMDijGyV9tBCR0d7eefAgNDEBgd9nA6vT9Zh0uglGzZ7RX3Pv38tV7ubEl
PESZMkzmR5hAiKImKZmemw0zGg6FDKpjVz6mQCkk4fDrecvXuxcELQyII4hS2JZrjFr+rZOh2toi
zqjcZcz5qWvCTULih3Q54j+G+9K2x9sWTYwUPIXJ9NFu0vhEvlquZHWxdCUT8QiDTcN/zEyoDXZy
e/q2Ii3soSI2esnL1fM8bfD5S9pD83EDuaCB6ntXau6gKVPzL+9YqKDpKrmZQWl4ZoqOooOn0rBH
M5am6s9GljtoNBsVzH0JdCpIMJd7rO4onBxnbxiJ2mBGG3q79bh92thJV/u7VDiMOADLI1g6GHmS
kWmQLX6AghnmKaKmzqke1/kzxnWKJFx29LjaLsuCWHPi9t5J/0T2LneWBIQrQFLPQymFAD5++w2I
oSC2uMn5pVEyXvVudkklcwMgwJhLGf3skoEyrRYVjSjNSgZeXSO3Rq1k5x6RHim3gPuw1woj06Bg
InGa6ex8KaH8uu0R7oiL/u9A1sZB+KLxx2eM48tX2Rqxf1+/+UR+OCUMjld4Iv90vsXxe3YjHvZV
uMljjfj4uZF8dFaCnoiSosHRPvMzmxkYMAu1zKRo80cUXW3Dxe/L9OdprFNe4EQD33IHNTMUMhrE
7+q/wMLg2f2R/3gxB2+1qjiBjVMuvpOydbQ7CV/X+WHEa10oTqMj9qwk4ftmhaJ9rjzLGiqJJVNF
S0HOKzU4EFpCLQiqWeKPIaeLSCeEPjhXP9JQLCAQLQ1mnIgL90mtP80dWUNzx7k+ht4uMxkzD/vt
A5tBWshCILtonRnUTbR+cMNsjgAVWZBAMC6nfVBsn6zKKG+eYoXAqb3nFFGngOi8CHc7cp6MYhHj
jVoAKYPmIs/bI4/Wa6kGC5EBXjQUWfKav5Y8obnQG+CoZ28yfeGEYBgotrgDNIrMOvBnHHfrATUo
73DZvq2DdfAarYhEcttJWYzVVdC84H1c9ZRf22OP941iAzOkuV2I2A/vSxXQ7XfFKnxO12U3k/yI
fg0+X8prknbmWQOpt9B+g7UuGhyc/9S0fv0pHP1RdZY6/4088SDKjkLQsW7kknAXWQpDyHja9O9x
GOerFVIPW1BdjNbIGO8pj7Q9OkMZh11BsykJfrBZSjxuNVdBB+qWnJeyWofBATX7v8mhsejNqd0v
NbLvCSDLhPVd8iLq6/UKuu+Q2onP5DtJ+BduUkMArQRKbo/4XoCqAw2pRqFLpu2mqUC/K/+k+sYD
dbnmOvAGneIkGqlDhed+6oB7ng0VHYByjBgwCJWeL+enqglRf4uLN6dOWA3G90USlX1cg0HzAt8i
NR0OfepKWWtzKy69S4EH/bQePZx5h7FaMSIdtDL/vViJauQq+y8aUKGHf3SV1w63I7Dys0fVo9LP
AvgVWUhlWxCeuUCeZ55Rcgr7Fu3FKvvclJliKjtNMX7LQGxQj+7dplY6oRhhXp98m/amoijCwOA0
Av4pQyOwvuDqVpDT4XhVNIASG2tRr9F5+RK9ftEAwaFD4PavjvmgWqLHqMey3/MnZWW//7lHdyzC
tBSXnMpDotO3qPsmVw6QXi8r/3bK9KrrJ+V8/VU+NDx00HXdhkFYZpwf4O3GhPPmbT6w3wWPhfls
/dc+p/kGql+bzBcRqQjwvZaXh4QOzKUrwRPK/9RhdXuTg6nlZ2LEuatc8XQGU/3QbqpCd6g6qx1d
ZKKfLyruu6CndDOpEpeQijt0BGpfe5YiacjKXU3v6YyFyftYKB1U8ucoKLAqgswu5/d0uUCn43T4
za91vtI+MhTaAgHaXZfHZPI/gLFu0qgRq7cJ8Jr5Z089iZMLvVkGWHmCeEku8enEeg1loRavfFYL
J2ewiex5YWPFdqdOCXBtN6AyckJDwk8qT9i5aW2TeGFqBIyucFfEp5MdiY7zNgDvppfbfPzMgtmQ
wUKnmzu6bIdWOReSz+FakOAwAS85/OzRkkaJrdiASKq/iSKd22GoN/945mQwNKJGRNMiRyE5preo
XtgurDn6Z9Dq9kE/VBwCe3fFnLBaCiOGvgHma81uWs36xOGKXd9GW10nF88p9HLDVSQBGDxwYUYZ
UquMBR8oI8L6bcAF0oTf+wN9TEGgXh2PfeIz1EezJJNB+XZkIQl7tjbLZ+kBqYBC0dLJMKWHpzyz
6skllUQiBBH+iGkX75T1xueR6aWxDgyVqg6BtJ+spIZPcPqMRG+g4nXAok80rtahBULT2v82c9fu
TzrBSn3SYtvXQGCmtWhc2X4DOhHdwx8D5OMz1YKPnLFQKZKde93LG1tKPzOlXtM13eVBBefHeOHV
RcAhsAwkfx5iiIR07RapRpcfRD93BCgpjFeGMd9m5i8Tf8jO6q1xuEDo40GJ98OjqQibe5Avm5XU
btXExL47p8tPPVyIHp4u89CAr/BAlZ+xJvy7KvDcUFNEjRI8fOtUcWKbFJzL3qtdtf5ucRmHdF8h
8Oa0vu40W3Sp52PNXJ/OdnMg+RWzfDKpyMUqXHUCPITREKLmU/lJiwkgULeH1HBzqDjihuG95tX0
M1gVhloVgWmgZPRb0y0CkF7sLvjpD6KCU7BOof5BJDBofj5c5Qp+CjrREgxkQq5fb6CJw6WoaqB4
G/paoaLhyIa8lqIzOsIR6j09wIPZ+R80d+67vyK65W9tib4NWtiTGiLTOQBrZ14NqGBGMe6/G285
Ryqeqb9+5ZCto6XIoYfwTs95cyA+N+kZ+zdch0eTeIXhtysUUOvvZlMoPykzGRzTsgj6vN5Dsqxj
FnqYRXV/6PQKhspwqPXo4hfsIsMVRp3qMuKWwh7b1pLLaCGT/yB+3/JNxclioPe4BuCFbk666rhV
/OnZdodrSWDj2CDDPDQTMHtQrfD3XioR3Q0IcKsoi6i32sB3hp1E1Y8VjcFxaPQyEARvLVWaR8en
xqrJ16FoYxmIGCdIZVdXZO1HCu/quONc0yjXPpND3O0avCawypxKydy4JtuRytTxgq4BVXZ29jbV
uptSlnzhb1gs39l3DzYPXgLyqmiDyws3w8PJo/0epDwItNig80HOoriYeLQpPQKivuAAEAW46qLb
L/b+ZgnerXhx+GIw3B16VnnL/TAq9yGpMKRFTTKX4838pzH0RmPdvcvJUKGajZXxnQPyZL4tL/dV
REqnH5gA9y0ZM2C3Z3auFUa8hqGgU9Xg/Pasg0hmTbap9djvi+1PZR4GgOBDGz24+fK1xr5VoLwk
AcG/5fwsZLfio70U+9rXHhgcX2K0BZJi5rcIngcQpUI6yGwBVvh1+rkDF2rKi7GwGksNLFvCqvLL
adkS6wjLMr6aBQM+S5X0/nrqkgLE7u8qZQVFDZr/KENQPcPaXHwsTXzZsvNY+aK1+K5C/ep1c5tR
MVlMUzewf5eiAkmjRfgXlCZE4zWnGBC4pJMQepKTdyS4EoFGC3GTac9bpJQmagaBr018FqowXHp6
iScidnWknIQLxCDFraQ0ISgcayU+H0klsQu0acBnb4P0K3B9ly8hdEM839VH+yzO2s/uZ5MZ4xW7
/9VHOWmLvFnYXaELBHrff0Yp43mRW+lW/mQ9YrcN/Df3oY52LPxL5nyYC1y//AW2+Vm05bOeFO5H
VHJ2gPiiGxUtxvZ1Qn4ZOa+fU+mlomM9KJzjs4QCtPRN/Wsmllv/92drXjx+X+wnip3E07XZRsEZ
UspPk49eHQlIUrgS4UxgSVdy8UtgtIydk8b7A1+cyzh/nZzDNE+D8u5JVew/7Yu/NL2IRVdlRI63
yJAg2i59InuhbDSSjQbgZIdGZZH/34UGAB6/rmv1MYPT+t9PlJZBX5BJhRVF6VvGkAKggBQ5aGsP
dKfDQyHnyIOJIUltJrVkM05mESmFLdcLnxQYts00kfPvkukvQiESTJto1F3LO1OvNFrKj3RLxeEC
ytawcMBW46Za8d4sSZ8aU+m9giz+qluPZKbuhJZTikjcCmAMyCqK6khSfdJlY7rfySL7hzccQ1RU
1mnRQHAaiHwBMNwFWpoXdL8Un4LRV8dYrs9mit5vhxNeomYLq/H373zZstdesto5AWo9jmyDcsTe
lZxm3BWb6AzYmpo32l+NWHWbPpR5Wd6zgXnLClHzSJactviTo5l2rAJ7dWoke6tX1a2VqFcIprUb
gnWa7pcmnrplO/ye+8VCDui7WLv3h5NlUD8SPfd4qlgEmWzCBL6rv7rYiIxDFhE+eYi0SDSToqNF
eag7jnr8oosxlv9ixjpmEgbYHSSuGV1Lxmtd0W+zZ9srFdX/J9rodl+geIjSUY7iM0k2+c+zjvDQ
ae7YZ/LxBJfDkR/Ia/JLEp3UYy5DW+sR9eBupf0N33DTtTMAq/ngTIcZjoPwWT+pyYr/rgvy1aM7
fXzMS8SE0ibxThcVpwEuJkZ8hiJnS9T2JopkC/HZM8+KFQrko9aWDLtF76TF3SIlD687tqEh67h2
A1h2ORkCMUsMzPwDphX/WKVF9bwcGOJRWrFUlK8VNu0V1PZdTir1vDJsK1jgRrBU9nSSNIVnoN4f
i/42tLdFx6aLiQrJ2JDK2+Xs9VDeroxftspbn5sGGJ7tYOZD2qOFJD4v6AXn3LlPY/gsKTLg0M7P
ckQIo/FjcQ0mEYLsSU32BfQDW7g2QyS1jdnNP7DNbfvlyvAtQmKXqsYsJI/j/BpTx5EhHlk1hrXu
2qKuv/FPa5UW1HmPqLAyw5x1KsWAedC4HFWEa8NFH8YkTRklYvh+RqvcrcTkpTpTCccGYOW+jMlp
QFZexLM7blL/KlUXmze1URTNCcykusyD+SYoPBNl7P0GTnYL4EFmX+x2SuVLoDNds5stDcnX1zRd
oNOs9RwMIIvVOGD7jw7iyFMEdjhKEr0BTIYHNCBhV0J7jTISqLxr27zCuIf/vKS84YiK/an+Iqkw
mVgNigrndMdBeJ5Qp47ksMf2JBnuZh5Si8r5sTBIMLxWsJp7JVmo7G5LsAZXOGCtmeP4G/lF/oFe
UEW9yV67nEKoHF3db272XG+pFTC7NhRDF+HNI6oHtI4w82e7muSm/KcSCS8TaBjJwsI7W2ixRy9t
VLqQYnm9nKJsgieAjy7Z07nVNA3Wk8Nn62XzMXMYxHOR0Rj8Yik5+IFEYLEnmQoNxqGxkbk2R/QX
2BmoFFuARFbdSnsFcisWy5ThcRHkkex/lCpr0NWn9ebUztP0x5+buTNocwfRG0pR86cDvlWfAe/V
dXHQAR8iKq3WQMRZuPTfxTC622jFjpJCgaRZBc86e9tk/ZoPY0cInKvYZgsGn5v1NwfEWZY0jWN8
bpclzkMWMx61s+n2tt9qMfS8haiGC2brql2SFp22qGUR28GF7AbvBdQTS/yv78WquidRUP1vcb/8
fAKUxjIspxjfcAhCZVyGvfP/exyDA8VNdoQ8MBaLLWj3Dya2HxBYe+Z4N5MAc1E4D4h1GnhicAKC
7iy03EjkM19kgXVb6lN2zXKCOnxwgEjVwy3NOtTx06YboESGkHGhg6e3NcVwuaorNhhqkWvc/9iP
roR2BWTZt46fnctUQbuHbXcMMbqc0ZTpzo7NNcx86wvkiawsr/Bto3MP4MebxeNwSfIBtJPdo0fH
mBplH/EgSFykQGV+e8PYYp8haBM/PklsajMjBSQo0V2OSNIm8ZflNEQBLc3H0+OK1VwUFWNkROPD
Y9pptpejvLAYRTQgl9R0eR3bL3b4QRKqw8PqF2XEfDZCOR4kgq6UkiyOsAoe/R0JuvJcPe/1rfwk
RoVUKNDd/cT9zLCWBF7I+OHLU/+RXS8fbhTWgjs3Bpi9BhEEyRaQfYhrWjcyl0ANohlMXoveD4cL
TCHcA++UVydfVhzKd3rvUDYk41ZazprXkgrLDXO+7UBlwDT90y6TUwedWvS3nn5XDVVynFymcCKS
I2yXzkBXnXIiO3ZbEsr12ttkzlUKGdoTrc4II4ckoVlVy1EtkLyVf0uHEXA7RORppn86p6wGOhNA
PDB2yHnN4osdsLiBgib0jWBLg8EgLiW33MM8bh10uBbO6wDQG2u75Cj8kDv1PwdSIRwkx7bSfQe9
NWzqyZgoUz1ObkS0aecLIf3u6pu9YXRU5PZy2hrS8rIYSfYIWgne9ZVqsRZ5+/Qw4fi/Uv5zImK0
ot+dNc5kU/AleNV/wfYWtg/leZ5HvbOmTcGpsM8jik2UvMbeBzq7dan1M2CAhOi4A1deucaeMwqU
hfAYW5ERde2RVJr+TxbVgdr5HYYc2S68bDQ9UlKqBCwD2+cDuLGujM31AERLSGKOau83o/pTE8Iy
jbtkmr97faJyV2Bg1/u2uxqWqxKgNzcj0rIbR3SECSAlUT2l+sNyVrhnk9721ESFfmB1tEyCTHRT
rjb1uvZT6tY/nK7yiLPvSuOPk1/J5BYVLRwB+hxLYuUIBi1h/R/KQAu5ndDL4KU5vLrip01SJgd7
LIF3fPT/Luqwz/YKQXyBSULhZfXXAssU47bI7xb64l5cb8HOIK4p9JOKq3M71R0zsvKKFan1gk2p
+Yvx57sr56/NsjmuacS9yyKz4rOODmNIv7f13ZJeR1pWFRxYUM+vf6gXHkzbVBYUVBeuk2pSHeia
bs4GG7ENYmLdXYQeGK9XZuDH389WpTKI4fRvH0yM/4I2FMir0thIgYDGBV/VZ2eZ9HtgdlyxR4UF
Db3pfXPkryaaT1AFFh85EdnmiIlpczeKUmBbI3+8+/kVjcQLlYcj0Ckn5GdqDxvwxRCm5Y9vERWI
wA2y09xF2Do5JA2gqUPoQbNmBnMad1Jusvh7As6/Lcxlo++g5Zo926XBKKNd5wcXKbrkzB/0+4q6
NAYZs2xJtPzQX5sotdvLJmtpVHWO4NHn4rah1XkE+Ja45AJ/HsDn9V7CAEentpj3CGWiagqjoSjS
aGRm1MLLG8f4FdDEPOi+A/U0xBu/6MtKWjgQ7VCKK1bR29kUqjKH/URd3wrE1F1wIKzU5lzzGEn8
9+tHvFPcUewAUsh1oYOqR4+FAmsQhlU2Lbxx7FYy7QgqHpkv+jnbmJ4vcDki3RvWTlfMTWxb2CgW
a176Sbja7A/eLD4j0tu8vtcAsvf0sEzBoNqcc9TnieXZejq/RKZE9Crg8E192R6oVVJbvTEhAokD
fyLrgTbPCkYx61fnFfm+bpF2QosH82+fCVb1YyTBxiZSAe+LvMZm+vVcwAU0C21K0qmOoIW0xJgj
ZBHq1Y/ZYvOPpllrtv65WlmTnVtaro886+oJzwlCvwF/ip9UpVCR7y/RcPuVGl/e9LSug2DfPUOf
zoW3iUdeBiOvLg273KzAz3lH/0WAf4zg3xCG6qPVSwzCN8BtQRLhm4irmtPPpsOOp60adM9DgwqQ
7TVlYNdvct85T5dJ/nv8eiY5iHUdQz4BhDWKzqy5+sItOUkJ3VzA2sitRSINa6GgRPsCdJn3f+sS
gYe/aUGz5hT5yRvsTNIZgcJ34Up4prnsqb1ALO9vY+14yNugif5UPg8KOOXeqOF9UHGy+y/GlOxp
bs+WjNjl9jLSgeRisGQ7F6UwwS9CA0WRRuCXZYlt3/4BbQXM/uG0lDOiLvHhmjtdD3MVESGWH8Ns
LR0xIwDMiTh9d1flBzqSj694XUD66wklWEoTXKGaYJQO3gFw5Hfi+3UkppdW4AQLSGrojKKOrSDo
cYT+Klsi+4QlzEzUssge/yium0d5iGFnYf7C71BWvdDbSydLei9uE7qyZ1xv817pUNxxK2XRb9PB
cIh7pw91Fs8Igv61figGH0GGXHn1cawSCoR5f9XRMJr4vh25yCLah5DkfyUEAaQJOM7d6MwyIwH6
s9HejL9kRLwheJHHI8JGIeQU4M9pDTv8zCU9xwsefvVba4tDY6jGgCSsWG2Odm/FapSn8AkoyCqU
41Xblx5QQxqHWc0yumMqbzg8ZPwy0O7cMWWJAQ7laQwY9Q9qPO+7MG7ehXrkD7fl6yFH97EEvSxT
UytxjaMgbzZ32eoe7Qa/aMrdNrEUbX7KT6pUHsus66bd2m4HC9a9Hy9GM9YrQH/FX+38+Lkmd1Bk
dyWHZCNrIOdqrZctCbYoW9wx/NBrkCE6bSV02wCYW/ap6em/k+HBCaR2xtxoQsojoJJBkbjiUghK
DD7K2RVcyXPMpuiILMGfUrhCFDgxMgpttc+BpLdt/jD+zxvR2G0bQIMatppnkOAJX+A2kWzNpuJB
N4vOpVfhD1Pz3iOJ8NMY1jTvKZwKnsGHaoKIERaZWspQmKQsufutF+THX9cdDnWIdZ9ifYdjTInv
kxGDKfE1aKJ5MKyQEyJn9WHWOzKkmqQxYTD1AzRP4+zWIrvsZO/rIkCMOp7+zQzgoyNG0yvJh2hu
4+kALKQ0Bma7d4dK3VNhRVeWzzQrKzSVBqw+mnTqWqH3HZSnTEa4qBynauihUeiT2sts1NBlL5sI
PvZ9imUhjN847JHV4k4zGjeMCyiFLhoKnVq2IxIUPeijOSEhvqQcLObDXKefSPV8QGKJrob1WCHu
F9FV8JmtOMSZD3IoC5HH6zYqflooHpEqhB2zkCGVls9ofA+2ZY9710zGw5ke09Hic7t1zxPDuVR6
gtFF/cyPBWIHtCanvu2AgraCHPmetM15+utR5SuACoY5UU5bHIiVR+ZRz/qILocGw6MO4dF1p1Pz
gDhmDMCRoc17z3GGvh31xazFtIsu3078FkTWyh/8dKXQ4g5uRWdYZAL2xT+02TgBHMgwBtpDVT1N
6hRkiyOvWry+QENKr9FmFVtk2mkzcjIlxpv946dHjVH6GuVi9KhR8GcTiHu3TdUVCMhNvCbboSV1
pa8iH41O1A4YXrGTSkmJ9y4jVVXrxqh3jkIewdURZOgaFtXTmYHEONuP7euOWnaZ+y67GN2d4qia
X/qhM6RFMWhAU5cj68wUba7y/t35hfs06xsYBF2M0tWyfC+eVsk3m4/0SygjAadNsb5gYlDWN8GS
sKEPoIMbaNgJAEmJNg46WLC8Yede8yUSFUEjupV6Nzh7DIcb3m12xRIunOCPDTXc9JFyhnvQ+O0S
fgQm+nAqgidw9N+oCMYGYOC8Vzil3jr4ChXnlS15JEJq3LtS+ZCmUic7WnP7HvFbt6QNoXhJHd61
bT22kOAeykOVyA/5UOVpC4fiPYUAdjQpGzm9zhdzTbYAONmQsvuSukTtejtfWgjzMUlHyCsU0DFT
YdWpoTn1TcUpSPtuOYobv477fI/usReZ/3Jxz9ZtwAuL6NpogQ7gBu30+HBdDxdCOFPeZssDLw7W
SCuFPpWsDpwx+nDDWtDX0GVAz74LjYapo5KNxWr7bRK/DL9lA9Icw8I17ptKz6DDK12c7Dpz4vZ6
J7Z6GaZOq+x3wiCsDPzJVW6Tg4vyxapgLeRx//cmz6G7EaYy8rW39OSRRJq2DxEFt+08JbRjnbnJ
O9NHKrvhMZ4qWXkZ5Ug+G8qDge21BYAypRHaX4+2rv39O2O4WsXJxl54/lz75qb8ObXf8ryq2L4G
Mye2pU833xxiU8EUE8BQepy0XbViDClKK8Ig54QkXL3cmczEiZDDEuaRwAhWjoGbdR1u5EqopX+5
qEc38/kct6mc7dz4SUhHoFpNiiPjiMg5Akis/UWzYHE4ANNjXJ7v/lvKpsflr55wTdADQ704RLbg
MPHFWZlT62MSMyXHSkh9ETD0J9rBktgPxifCNw6lK6DtY2uETE1CKIZidljhfHiXQM0NHarm/wdZ
azb/WzvvtkHDSAb7qzPBbUqPzpitzQNpngMIJVrDbniCzAxNRgPYsCAoYBhHnPN6XqPk92DXn67y
JFG8Faw4eiS0oflGZXgatp38CGQdFXnucgt63O5NsW56uigfQS/LAOe+oHPQ8dDHbtrInVVzcU4v
eiE+W4Z3GAq8A+e5+e5JFj+vD3kzCEqzBdi/X7jnDzz+hL88D0oNIHenaF3Ll7Wir7v3Wp0lJ/MN
d/u+Ts2+x/atIFSWQ8NzTs7hD4V3ygLLs911COVhG1UprAXQp9VWMaAz3aygJiOIBnh549mCf/9/
Wlz2vEv0L44ByTdlHJZi0y6TCd6OLTijDiv6XMtH+FXATC5bI3om9r95IpLlQBqZvdA2rdPRf30Q
NEhUPE6dDm747MgKMeNRlELrX/v66pLkwoh1yji8Wc/xe347/qrsQ5N5yJANJwE6hiF8/7lKnIwx
MawVLfZbjyeAJsSM2oFN7BxeIoe9luisZR2kfSdYmLoIFHKtHeScgGq99tqVJL/IVKnSAOyvGhkk
UettFDalRFwaeG7tRItsDKvrE3z9ilTP8ep43gb3h7u4USyZiyYIvJXMTyp6jBFVyv+VVg6MLLpQ
YKfZB6sMJWO/1SyWll2Np9P1h6vlJ/h3tn+RQz5cxk0S1A9KbuuR7mf6FPTwQJUWtk+aHWgfeU1V
gg2vJtUZMucR472MIvbvf6p8pFWqpP+0WGAP8HxRTZNMNi0K7gHWy0quzaMws2Yq8sKthww/ySOT
i3ZaLTSma+DS61u518djmOIEit9A2QjG/yutjQSeQFZhaAFmN67WxRh8RDWL5Zvyu1k9eah+S99k
kWHK6m+SMbfZsvlScEpC4KCFhufCBS+vXiFrZEFZQaDeMXuJBQmZwwcmv9vY9mkrd3yHR1ETmTTa
Kf9VHC2iE1u8v3CNs7rJ2Rk/lIVfP4en1IJAJM2C7wSnx54ct3NAYX3PXT3Se2TCI4jnnLdmdNLR
Z4hZmdLjhgKw8CTYgZQliNVK1zBpsLU+gudBs2nRIwe51Xe0wqoEr4bYFwqYM/fMdfro4LaCfwN0
/DUIwWWPs/GpYAVDaGq42thw03KsiEQIW+K5XGCKqqoUCYcAuLQ4kD5Hnhb/i/A6HaQi/Z3vfBBJ
vSO6DSTkxwi/OLtvDNjSPIpwEAEUSs1u6BAD5sDdvsIW0zLmuwpVV9EF+QXcA+PtZWx4hQnpVjZ8
/nPMLjfbB04aUrDRohX1gn0w5gF2xLF1PMRE/28rnouk6HFPsBXam8bPCcq30vHAxW0TGbjHU3Jt
h4llScxVnttnplOnhZNHAeMCfZaq9/Fruy/y9nlL1uYkmfEQMfLoguV6YVz+uEEik75usfBiKvsq
S6lZsR7mkdzTwqRwlwTauW9yO/VMW/KcVZH+x91ZIT0kegGFZOtIBaWjLwGfaq5c/d1q5oSB27xz
jYfj5IV6R7VyGaItotAepf7rH+p7bRdVAEcEZa7nY6MrQubeWMhLxyNhfhk4ogmwEg1abQNFSja/
0O10jpQMnZtBvV/1Is1LfOt1gK3d8MGmRcKfeYA2b40ff6EFaElujSrJ9Tp3qm3LAi8dYOOFgaHM
8yZbiSec5phr2T97dZqJ7KS6Gb48I1DCFH0zSvkfl/Yj/k0SGTWk/HLk4Tev8Q9Tx++Jx2/cayko
xFDT4dnH+jWbnlKgX4IUbspLmReJ6qTwXD7oNA9VU0cfpZGNYpKDZxlXc9qaZYeUOJYr6BmYy0wJ
Dz2UpGcWVTCqRjo7YhgLyJWkWx4OYXY66SDJswqiJlDoZoRujaQQPgky9bCovYUGhDy58pAl418m
KLp5bMTqM3pnhYMf8Z8kykuevcRv/D3UZ8XbQ4ZVOtTf9v2WXpuoQKpHfXp05cNZoGL4x4q+RC4h
gcNxmmTd32XJOZjKYOWyfaIa5pOJ0tobk5x2LrdmU8/H4AQMjv2lNJ4xJsx3P75Aj5dspizePLT4
GTAD0OM0ePRZkLRpL+5iuGQd6rSC7tfa0UaJmajEyn+5YThxLTXlvFyKb2OluieY29Vz2c3AG0IP
rd+3s6HFuijS542/rcO/oyvL9tqgsfh+zQLUY/zbRvfORZT21oyzrOvpiAoVb1Iuj610UvM2I4+u
sNRCniXVBwfsW9vhRbtWwd5iSmUFsCYBOZ+G7GN5yc8ZFLDO/B/0OBSGrKLrPd9AoXw9tS0ahXyH
t3xQ49k/mU3vd+o4WpqO2Jh3utamTMT8rGUja6cocf5KvVo1dffrDmbRhoi1zzHyycKRX2zR+fq2
47KwWg8K+1UZL8x1/0ov0UdsX8E9cw0paqAQzaa5LW4l35PaKGP2rro/lnnB3gIo0t7eKYaUU4kG
BlOfbiS/KwP+9v4OKDyTSMeFVVoOEJmK/nCA4yvXy5IpHOMGz3wHIJFjpHoDiZ2TVb2ognkcfe8t
egFP207KJHtWt8YRiv4YN03EQYNVbStG+SHKR8eLhi7OwtrqvM79QsJIO3EdqRQACggfzspdf2ry
hmcu1qgQ5NNikivTPJlM6y+KSwEsvhQG3cM8PsLpmtQ0xCET4v6NTmkVzcK9YroMM0/inkhckpiQ
fE0mbuYraYUPLrCCoeQByIYt+NTMyKuNybQcG6HgoAXsr90ytktWrPjPZMsQgWN6nGjoIEPj65cZ
r7kWLpPITRaAX8YzjXQWId00g812mtoWRO7gBanJf6Wcli4UbYfv8xAPR8MIFzU3zf7jQbZIxr+m
/X727DlDM8D7Bh6UVPHI+/jyyzcHg+zUOIirlUoVduBGvUY2rZVuKolByUt3L32zbBW84XRYffBC
/hbl5Zj+uU7I1GFba0AUKn0QxPY/5NxzKILCcQEGZMTPkAOsGzU4wzAtJWjMGhSGBjGRIbvS9Ios
GFe4oKIq0kI9LVf+PyuyoNIHDTvqLEX2aVIsscUNT+oB8XT0k9PiuYIpowp/mZxrsgs3p22BgYGh
63hxL9GKYFyuDSEmrT2klqElZ7Yp2q7rIhi3S9pLuf7DTkgT6Ak7/GNp6Alxl6UIXKwWvT9TfrXS
7ko/ygEQScPXeRHP5zfnz98Ri7NGXA0U6SJ2IN+eAP4FWcmUY+s6T46suzKUQ6pjpWZlKnRMZj/k
96/i/d5XsO1pFBd465+4YPJDRJ+qftvQjNu78VJO3apGHBdiS5RS+QA1/Rln7zlW6LKTgZN+6iZq
lj+QKHxBtFiAdR+mqM9C6ysnX+wvlQjcXzx81SWpTOpauTYCEsvImD/8Vfenkkkw9deWfQicqnpi
fCrQCGSrsGKZa5/mofPCxfPQLpVm9rNdyiDEa2XP7RIr7yCjV/QPfDpIP7e049zmNFEwPg4lFpbF
ubzM1hZhKAYRoZkXFUk7/mV8zQlmSBc+6Il4IeBbIXlD+SGGLN8Aydx8nYvLtHY33pCYuStVZ0sO
WWQlJYSQPLI/bzR1INyd4tuQsUhqLshxcZyCmwgeu4U4piyC1pMl4CHjYea5umjKYJbY1/nsRMtW
9Tngoj7IUnyhNign7QskWire3kDxfpMMHtxRjYOPy+rTpuy+byTG0nS2Hyuzue53x3Sh4MZbsOIg
yzH/0K9obFmIZxXEA0sU2w9KKSz4BZJJV7i2fVpcfC6fajgBoqyzUt0jSMzZok/sQ2SBwWhBh2Cj
F8WoNZr3R4lHB3ps1V486rivDzwZaIOhUpf/iRM0m3zxIj/z2s08gc1Yr7G1AjAs0ga1xx+d0HJk
gWS9rYuhzZ+SyNLyFkAPvAoXxbicmr3scl0B2lRsapHUBkiZawp3LDFrnyJRVTCG73FNDndPY2hO
1YNJ92ym+7t0yGTGKaeqU9tNKzu1VaIzXDkk2eNd6JduK8GP+kJMEhDlwbvEOhcawfyGjCcWeQoE
47R/9vmPQUno17Cx83dsKjaRdrrhkFwh8Nkfwd0Acom6fwWLyrRh/IGkVNIZSomMz4kGWKeXDQfd
zG8lOFJOQ6wqjESUUbOWJDnoPknfKhMAAWWCX/Lf0f0DP0xAD6+jA2GJqdRU0OuixEBCZijVfIiK
Ah/hGGSjuvW7OyHOrrkzRREn0e1fwzTuHrreIAVdM1odeIJFgfC2kbWEStcqckCkp6mX9tgUNg+D
PAHqQCEIFTkW6gSTzojnA51w5U0MnEYMx4NakToiwMLJLwXej5FIvnMaX91qc6N7Pw0xYBe4DlIu
t7ItO3XVcqnyAUoH7WbxtUp79C6M5LJe+XlI0aSfeCxXjUp6Hlqw5eTkQXGCOz9kwzZRvlbjug9h
OqUpsbw6zKEjldRJkJsi3fTP0E+Q99nFI/QyEqny0Ob1H6U1Rqo3/O+25WIYax88rZLD97bcKQTV
SkbG3LX7XbnPg3m6RC+L6bR9nuJ8zUN5wL/Ln2x3Upv6/c6us/nz9FXXJGGMBplyJ5010scrul0+
QugEXUAYeTlZEN63xujNvxD1ZOLXGQ/PyKTg4o07AS3YfAK3RFOHPNfrhNdITyPkjVPa23qH6GIY
Hat/wbwWCGzE8QhmsysZ78tHcOguedur0lllHG2mQZnevtZ31pmfOJySHMAFpnmJbiRmihe82iIt
9wTdORqFPVIdndejV/3Hdbd60zCUOdqj7WrYdiNtHpl4DaaS85JwRboEB4sJ54uXEEt0peGmf+KG
N+9GJU2ojjMl9IIikOb95bYO/ldxrfquz0BjNsp/iU8lViT8k/nROYTNfCamCV2ZXq3FTBPWbd8l
iIv850IGIUg3qQSrEQAv10tdenyYkoKXZpZ42O1isc4BD42MHb4sRI66hC0q5HviS/I4tsZ7h1AV
q8w6t5MFqmWsisHMMOnwduvVHAU8zXDGK7Ho6RmD7Q7ji8r+0vNzUcwfxy2fY9BrUVGSUH3FOYqu
Q2pMKRRSxmtXC3t2BqpJHTOyTDENg1Fhs5VDqmeLHtIveiji/K8f1Ugx+uJMmzYn1v8nCQi143uK
0jqmJSmU1Fz0LxBLQCkI4zL8SB3ZBFcl7JQEizP9FPDX34OVXrM9Cp4attNvMP7NLcuc2B8aJ0gd
faDJzb/rojS6MaIoyxD9PLhjI0w+IaFg89uK3UHEH2j38QdT7VB95072s+ptjprrIUqofChkCr86
TBemGVXZI5DFLdmM7WmcEoHKa6wpiHyk76626P2z6uTsuZl8zmp0OQ6SJ5o/oDkAfze+zMyKI8ef
Z48aKOfU8pr+GNaXxkTDkuhlu9v1La1A8dJLq88rwrpMAglgMTV6hdfznTCAWiZeiNowctaL5DCe
GflcBY9GaqowB/1FAMKkLuTZ+wj/cshrj6JdouaUNkpngkjyFGXYuulTb6VaB0UNcSGNBPWmhuEG
jbIUZ104Gi8pJmDqE+Lg9X6Hb27fArfAMjfFafK4oo5rZYceJasKCvUGFwgTtGL1NcrmWuOq+giN
uEXUZD8Jymn9PkYr7iZf55scWJy6+I6ojIXTllZjR2C/PAN18wZVkdFHRpDrSauZiPWvtSaQHE+G
fUlzELY1HI8+6Eetw8osrcDzmfGl/R713c6ZyhTNbpm5+pLsvaRQ/KTAyBPnCHcpvHnMxR8BUuxW
RdB4eG6yq5hT5ygMjEClK7Hqn5IY4JgojGnIYoloOK9qiwivEQb9BRK7nyZCrvRwwLd7p2/n1Q8e
q0HCHngKmJaBpWKPkyvj0RayCP3n0viX8h4lLO8a4GflhZnb+M4wWtGbA7IrzwMcYWxCzcD8RUHB
Xk8kNMSyxjcrUPPQtYI70FNKEQFfrlHe4JeM7L0kacey3K4wMZD8FcWB1iweqj1RgqAQ0c5omGYt
pQYMTI4ZHnICKcKqnKq3v0OTLa9PD0HfPKa/s7Bo+MH1wkSTwC7CoD4QtarXuDITHf6295A/5QMI
5wDEoqsknV1owBwQsiy28MQhSRK9CkiEh019cNurp7J02P+GGoNbwyEyl1g4UjnNFXNvCJtCl2OJ
WX4484p4smk0wIr9O3EzivNl5CgtPW7vwqH3wy9NnUre8vi0NpVGNKKH79lis/hFqBtk5dcyS7it
R15g0X1NJ9mjiWln4S+knP0/cCWq5LShUarMgz68/NBNDfXvzgyq5uaT1WGBSWS1nk5ZSLwhrX5p
BgntA9yelQ/2/sU0DkLCVMVy9vpplkQ/QgesoJCahMTAQNxa+MBiaYsmpodC4RuhEVlgK3t6wULg
uOJMxPx4zeC8V49g1ZLnhSruN1PPrha1+fPtEejKqgCgrjrAFTb37t0QQj+vwSm2CvitipogcoZ5
i6PyLxVh4mF7JZLDyJxefrlXzLEMHLKxq7ltX48SWs+e9tCh+gJi0M61ziHPOtmawJ0tO/xdtGN1
Q7tqTfzxXe7fjBahqb/TxDfL8ByPQZkxELYugSqwQjuHoKs32475MchJO8nk4MVeRsYyU8YKM+b7
HiLQzW+zdlN5+bAprsV/hDew1NCNmHAR8QoWu6yT1JHIc0ccQqYm1EzYdOXduZW5zk+T5+OkyA/9
e6VueH42ISTH0iAomG8fFrGKED/Vl1V/vmvL1grFMJgrU0UcJk1h2IsJEsCh0wxjXBrYPoWw1RWB
rW8/PMOWI0/FqlQw9rRoWQ4bTQq8dJk5kaAFrLr+1e5p4zVRZk3gcXqMsviIw3tfihfacVR+sqHa
N783rdTf7e8kYxftfuJNi6osVE9erPbV+mjvM1zJvaVJwwkjoEL5VMll6e32evwvDOXvnmwSf+A0
j91khoVUXnIbiGE2uhDrNu36uJ9jzEYOqzgC33TtdqPAqVVwHExELxfx84vqxqB3gjdyKhx8KyrV
4NwcR1QQIKyprF+TDmn21sD/7qFVbozxUAwSeKhvtQEFFhSZglBYKUqTPkXODfZ91EjVISNIKabA
q/DJO4SKr1vjvxJGXHUEdkBxw8GTW+4TFw7V6AbnX5wxu+clIFgJjOdTWIZG+U/EDSkQtBGrhYqP
oyU62HHHnJDAgVl44Ev3f9riymJsvGE3T/+vJvbrz8fP0FbloU9HPfrL/FtiuoEAat47lP6fw50p
TIMVDWZ9L6htTOI0GdAR1UfNqpejCC5KPPpIeBNkMeBlZfHgT8oqGz1vJy7e4ESs+XnIrqFVRuC7
a+TwDLkMUbrOdaTJYYWlhL9DUOkR8ufT4yvQTh18pm+s6eCUxh8V7m7s6+vVoiZ9P2GLLiF088lq
ZxLGJAB+XORU4KMRrYdsRf9+2s40Eb9jvKiSWYCQG3Vs8b8brrF7a0YwjBrXOs3ucdRgGMDH//U2
d+hNwPE5grXVyRgXa24zv+RgD/+23LOcc9QKu2wkjy6bSWCNkqMlUfVVA0+0F1kpnZOxPXi1yI8N
LHbbIsGHJbyMeE5GKh1n2Oy2KkRELCSzt+6pB+VHYOCjSKTTSD8ykLQZB/iLfN3HFwJs1DUEgR8z
4HkkoOBlZdm1m1k7qwpno3N2qQ1X7Fqz8Mr2kxIuHp/9Gis9LeM8xGAQhuFjNrLXxMB37Tt6M3Vs
GALUMGKOwo9m/8L1wDXYhY3kY5pQFb7cwhLi/U7Ed4wt6dddwgyivrXJmtMtSshIIywBOKnEtYNR
ZzglIKDkFfdFUzEMaOjaU21H0RJlBjkG+5dDa3p+yjJduWiz1pr6WsATx8xlYtGl78FS5FolVpRg
i4UGhLD+9bKHtOfenMKMceVczblQKqojLjDTtVkXkhSPhVvnTpIlhRS/I5ObyRU5/012cZuyk9oH
jF13SxNMGKqEPM6JQvyvdSCan0lV20qzgznC5tldAD4XbApGaHx0YJ7w6WotBSeZBk4IoJvRufjG
aaIIzztVLif06dXAXwQojf1k1wdXSpevDXb5qKTmn5+EZREELD7Nlh93t31b4pelUshq3LjngPjm
RAzGTPZ/jqs9u7RYJhnQyWD9TzKvd7MLnRiyHSF4tpITaIcyfHszRIjJPHcLbUQ5BZTwFKiLT3+m
VaY/kp2qrBYR7oTRtKCqvWHE81sa0+ReN3PqvIWQ9c52qfYmv5rn2qwCjXJkJE1yH0/TmxbQNEzh
L2RAcLz1uzTB6dAosKy6rNQ0svHuKvD5XJ3GLI+V+0apzv/Y6/dQ6dwxlGmi6pPnFcQ2xCNTKSpa
HBsozkda1bzWnqZEFBLxixTIsKbfQbzQIPbpzKSzcO5cWasDYq52GqVfcmtVJ1vVIlReWGQVNNYw
GsXryZshgLGNP4iXmgrcSi9bWNyz1ZXOiKgbHsFOybWoJ5qelbszQamFnzF3++a91CywQKw/5z/6
Z4EwDCA6+uiwM9QO3ctisGVJ2wTWfR5UvggkZUYJkWtX6ArAQqjyCoBGz0r3Mp/f3UdPhB0doZJ8
yAUDlyTYlx1ZnuGdpsd0WdPu0KVAI+2yzLZOfw3g0ML+jHJ/9pkGceBVF5KcxpmDN3no+KwQqtEh
b9f8m/8XG/IsITj8q5/T1OTqEPIzEdrSqQimts1P2o5winBc+0BHLzcee88PtapnEtgIAyK2sWio
t7gbPvk3zUVK1lF6gb1fY1dak+q1DpS4jvIwEpfAT+l3MwR1Wg1NOn1FjnKtHbJoSX5HUbD1W6UM
CZHRmex1VcftWpgA6W8x1blPf6RQFCDKz5byDuPD4pCRelT9YBBsGLa3tCo2CvQI/HwJkUee/HC/
juAAKykkeAh8/hml/xiKh/iwBT3gkopiUdNRbD3gOl+fcIZ90aO/sbZJ1k02HFyNE72XHwe+b0v1
u4jpksxZjf3erKO9vybehXQURkT0ByglIitKHd7gnLGaQT+EaogsxA800QdU4iSVgYDIgxadwEcF
SBluLbju4t3nNzJd0X9QDG7Fl5+0gA5iyoC5sz0jP1f9voDCyqp7Qp3LVhHqYtTnNiyAExNG8Z/l
8P+hUG5ODIs7eOodKnOTsltB9d3b221Zrqr8EF8ca7qYt+vEZPtMKQCtRfpfxFDjE3AZGCL6Q4tj
h4X5y3ZArE3pf7+CY3OEY8/Vy6vfmqgMOE2SnrYXTQwBe3oKL2qac1uIXMF18oXFja2EYzmtzoHL
5CjjTaW4ZFCYHYXBj9woVsGm3XJNGztMdJB4FgPqHGNn4Vsmw7RoXTP+X15TJCbe6xgx5Y9Kn2zt
c/vBll0/xoXGLbazrSZEoq+xsGVqTPeHqHmoROJQh0wj5TNOittbMVr//MHu5iJJhRwcFLlcVQVe
zyK8MYRk3J1Rf0JTfXQ+gW1lG/0BxfRx0+PdYTBw1IfePRyu+FJY7fwCVZz0WgG0KPKe6WzTWy5v
/TKJx8M+OXx0L5oeYMK2Wc6LapGPqYQI4eVN8yCoMR/sfbfB3vatsj8LmPC/iRvH1edL+IcgfBa4
zrtUmyxxgWsppYXDhi1aDiM7jG1Y3FBN/Yp6UJCGa5h/hXVQR9IpLb0JnRxQLscamAg5C/hNx3yx
uT6bttGoKTzE/pECVfFRkIaY9pus5DM0e1eKcnYiiXkZhPN0SaLQgW8Q2b7dS1j+MjmhnRZE55H8
UmhSSCX0R4Np2PWO/gu9VFExQNpPhxMHxKgFhG2+2B/BP+n9cuf2Uakem+WC+wzqvpZxivkOyBMT
SkqetqjSgq/U0ZbXRV+wSL/58EO2F0GnZOqT5izHVy6prEmHUEMkKECb9gxgq8wNU5lNuv0cxsyh
K2Gt1JDcYAneh4RQKOjj/7EU5gupiaC2wwEF3HSIMcTyZxatH6vkztzl15uOtABK0hVOGaigriA4
vUF1BJo4e6K62qCqmngjyfbezPlS92QxvvHTSnGkEV6rsRhSl7XlXosAsc7jy/Qdu6BBwWDJMQM6
OzIi5KvVkPgZjlOkgs4Glrb6+NEQUmpi16MrZoOJ3WPFydUQoDr88Wnp/J0YWCnXmwSnZfvIHIZo
Oh4EF17l6qc72CAlC0kBF0pB+ACzDJVebgKDPynkBrPlMu1dlOvQD37Z7bUbCN0BeaKWKhqPZ4ST
YP7bZntvVWoNEmhfOveW/tKYX0nahtNPG772PNO/ODQVGousY7SfMmmsnzfoeXNO+uPsvm25WSEG
Pkcx6+iuxDuRaKJ1zfir0LJiJGgULHGFHSxFMAlXbgf4lREwgil+8MjXj7RadFDnH1rYYC0gSM5S
bsGsvcrG4CF2CVtagXjZo29ayQzzeETvxoSDUMQMGMGoSF7LhjiGxF1RfkDqEVtKaOg0DJ/0DHR3
pDv6wzsJ2v8b8yU0aiA60CXGLFnDhd8Tbz4ZzVyCXNvUaOpvkf0pm1dFguzTsarvyuA2b8Q5wuST
JDOIA2EdAoQD4hU8BTGMd4qyEIUlajGkGEjxbN/0AqzStOYwALhfKH5eULb9+01NB/qzPnDOV33d
8QG7YEJiwoc4DNtbnpD1NiHxVCL5A0uEWcFPIPclWy4qZR61rWq7SZ/orflwP0g249XOoYGJSPvV
ZIILrHSP/6WGtP40NqNg7R53xz9trtHN1Y6s2w/DHIrVZ8+lYa4agDkhG8Ky6JnC/49cSpdaAqrq
aMFMB6kjLtO/OVs4LXmDjpJp7vqHMt+bKwOVMgbksefC06wITbwl0LmX9HSb5+EKQXejjJeH1lOH
ukzwvndGwezE9U5RA3WRQb8fKeX2U0DRJSaHzlZFm+YKcswC2OWAX52NA/tQR4m6Q2U5Vrts6PR+
blW0lRdOK8yPJ7bpEimJwcaeWZZm/8viiYx6oS5XXz/piuOqKv4SaDGiJk6PLDonezAi+hMQII0b
3EvR/sbh9DF6uZ0IGCr0AVTahhbvALU82VD8edjOJDZuSavQ1QYOfBLNqHTlz18RraYG7sabg4KQ
vk8DnxXbVPDAFzJFx3FSk60cg+tKmB/p6jt+Fdkx0GuCmpH94vQa76T9mwr3qCJ5ssQiBVFyZhCM
8pJoCSmKsjusmteYu1dexKlYkpMbhXGSzLQCkO9khVSDq4ZQ5IKwbn56bdQCPLBsjmzakLmDkBDn
lZJcUErzq+NygsJWYHU0rqxheyGvHWpSdr22x7B/LuNynHI8lQKTd8rOsoOQbiksszqSwbTrnxaH
l196Smv3i5cNWEpkf57wcLSNSWk1VmU49Ek/PNf1qzW2xDio4Tc4B4SC/r8msztXou82XbSzA2fV
xGk/Z7kx0zdOHCg/kZl+Ihhwn0I+jLaQBX99LRP4xhPN6i7MLH9Zz2s1vjHeE88ZUa0jhySJlz+a
qE73V3yo99DoPgeInGRyG1lEF3eYRt67UwrW/62RIxPe56RhNkncNlqemZzxvSHaBsjZnM3UF4Ef
Vf/zAEemGIOsI9aybx14+kC1O6i6JhO0egQ1ifzwYCSC7PRUIEK1MeVUN3S2oyro9UGgUXN+ZfNZ
rbBqglC4EwDDqWsT2Xz1M9XgB88u62R47FjCdb2WsmdXUpowt2ssXDsfBl0LD99zKXwOhWrtYkrB
8UvK52dRrrrDqrh7NXgM5FJBDRz6zupgOLGpjd6lWjz9GXjpM+gfZivoF+MXkKk1SWO+gvzbSaIf
YcPeZLcwELAN/Y87UN0Niw6f4HwJ+GCt8nACRPccjwcBpi7ONei4uYn9AJbCMUVS5ef/Bnw2td+b
h9HyvhO165foFF9GsfI6y0t4Pr6H5XYEqjqz+y1q4lCIJ6aq9Zc3Pbt5FZa9m9r149numa20oJzR
dJuOs6Wu4FNkIYFFJDT83/dlD9Mj/Vyu6XsRFAFZRBB5JC4Db16n2YMXhuSZYkmFoI0khMrcgFrn
uOwPlkBt1dL+c7pmegamPdHSmpUwCRmLpez0l+TXSdPoMChPzCwC8+1YhPF1FPbfBQxM6D6na9T5
Wn8z8+nEwMEDsobtNP/0edV/zjXPMd7/PvG0FOSP61GaJ+jEM1XYOooPY0KHigIMBv46uxzcM0Ov
utRvucjMmxetN3I7G+iuie6uUGdS15IWQ2Xtuuqf3IEfgmDomTXLJQz6Scz+MtP4tbw40wtknz//
xTD+o90a65s7Xznw9ayelmkPG83YGu5txxAbU7qo+uz/xeRiGnkSaTofkwPms3PgD/GE1xC+95vb
55p4kXJ4+eksMtaKuLsvH1FXHvgapcLw2ieFciYkr0W3s+DbEcIw7xzIHOWqC1kDB/aqeUIxGZxG
AapLlL31dOw+H7RvRXjrRb6bWIz780v7mv07riWuqdvxlN79dPDxD6604Ye0Z3aLyKf1foa1UddX
Id3wnmEOlL3qULpptb+vxwu26W2PxTjri63SGTYQqp3sYPcMp1PIZlxR/VCltMECQUV4LxuMDdpN
uhvaGroybGGJkpT//C7zz9ovSw3pENd+5+JzEvswfDc8d7o5vgFs6gskEOQNlp3NDZF5JupWwzwc
v6sRZpsTWLY+X+fbYJvTFLL5UNDkHEDV0+13Rjk483kGf80Cz3qzaR+lquJmyhMY4dwSmw0x448X
FLSHWth5d1y4+utJu1IrlhbiR7JPVwBaL3JA6oxgxxgGjeudenqh9bVZXjpPuMntZqtcZ+ce7P2l
He1iEwZhleFx268HOkuj5fcATqmlCzOsRiA2NFDziw1/6t1UCsg6HKsrjqgS81wmuiXTGJWR/Yqm
/+oE9ru6QG/pSsPYq+qVHBHLGeHEhfTpUy6JZ3SkY/zpnmXW/IluRiiG/11RED6GbGcIIU6tH4ig
61TQ7W8HSspKl4Tnserp4aS1igDr0YNg66Z2XFw8mmYsy2aP2URZUAUMBXBew0Vraft6du6QRF9+
G9ooySCO0hwRFIKX4IH3iyqqs1lUqtVuoxdWzLZnBwQRdOTIIVpskISshBlf21RcOMndEm/oIOf8
bAF2mvqiNqBq580ICPPyF90UN8qMXX2GBspK/zMGpJeryOtjXVJdmB/30v8pVYbiYhK2J1ls05Dj
2tQkC+WqUFbX19R0wDQOV6Le6o+goKJgiRiq2CDNOQW9rsRIiBJ3UhxAiKz5phR0psgJSpdSlB/7
zMxpUPjVQZVk8uiY5PKCfcbjVgH0bg2TdWBLH7YB2pmFmcfFDZpeP57OtnAMT8tjfRzBQPKYzSp8
FEHFkufLRZcE50sItb4z/JZttWzf0AktlFqQj7v5pIGUZWhHLyk8g+qDGNZ5JIQ2/DP7QNZhS/rd
sL7/KbouSnmZRG33od3ybMiwz0hvvzg+c2J873x4ubTmGuj8y2TCfYuUUWb86uFmS9JQD7WyGomy
+zMHQcTBiX4swyi2V7BjBUBluNO5LwaOvwYrHmwzQ4L++MLvxYNKBiypkWOsyFVxDyxT+VwhCqbe
0u1m+VQF1GLsGETZ9eyYrwCkI+BfiyVgh6fkaDIvrQepQ0wgy8VUOl4KA1uUBHRM+5zdiVxhpgt6
hO3oqzpHmLcAhXSuhyFR1/z6xGH926IBH5WEz7MhjESPEgU8I5hbrA6DIZYwjxO+6qZnTNfbSyz8
MRl3YkxcyiK+Ql3CsiyUeSl46yAWnj0rcgyedIJwqPf61BCrgl3kkSIA8gTbo3Y9HxzodXvG3Cz8
SeN6CB5Osqo2PmAnSnS8CSKsdBlnOIvpiQOmgmZBTChV1ualGxiVHNrSewdnHZrP3pVo572mI6XE
+CSBFzzCPZtjo30geu4yI28ybYPe/GvJDSufG9vseOYS1BN8FcpMrZ8xc39wMXrkZBC0zg3jVteG
A8SuB+1J0hHcpRR/Dq+mDO4s3YUaOPdr4PXeosQrcJOTuHG0VSAhelSy7QGQpIVrRjXxcH8/zhiy
rZPcmM1bO27b9ei7WJTRZ/MIdHDjhgkw+Li91TTjrOP+ZJIemVXUutzSpNNpPytdvOJi1Jwe9Kdr
ZV0LnmpF7ebAQ+osuCDgSd3Z7SqFYkkKr9ljcR9cnRa4EUu9xiom9Lpk7dFVTtx7wfaRqu6NEj1e
pV5K1a5iAIy5rbXCfjhuznAa23tdNAtjkG5PPdFiK8F8/8XVdgyGiCMA2Jt4e2xIZT4Q2bOZd4wD
M6WXlE1/dDgqmqtxKM610OsF+aWR7U+K3ND8w3sdn1jbAkFpQgW9aOO9AGOrsKEnF4TuCOG+AxMD
mixLZuAc5VyZfKzUfvPpInPB+05tzPOVZIo1seczt1nXDXshZBDgvrZR1yo2XsAR80ohJV/UxqBv
rL9PFZQpc3d14+DLvJ+wJRdFSAXBGrySh1LLWMJJkTXbmOf1OTi/3KnsSi7LaFZm/yETsRVnzEMh
PFL4HAgmVkgD7HT2CQzoR6Mail6y5os3uOWMxLDUjDu+vxEwo8JJUwbZKkBql/d408i/aJxdz4Gh
VE2n37ebOt+EJtx2ddSvc+HEZpzltskszJhprTEtIywBkUXgUqyiyaxVf7vNW9jjOBFf+xG36/h6
ISSsLKzRmvhozMwl0RwchFWYUTv4RyjVU+kSB4gIwkSyH+5FJiKnlC1BPIr931GXQ24U4YSl1s70
6y0VLfA67R6SfUz5aiv7CL5O56lCknyutON0GS9n4/LxsbQrBBGlz/5ctxxSke2QT0E9eKF6wBH/
szi3AOhFWuaTgTCEJcLJZPZmO6vmwmRPavH523b86r+pTnKOhaPP8dCkuc+gcBe49ZKJXDc3wtPH
XC6tFC07q4PkEcYde5NdcaABNmBD7VtaDQFZrL04DBakIbQo5URCODp4VpQ6p2GzKy2XivUSW2i6
puOanafgdKlbt1zMVpB7cX6P2GoJexIFLGIxww0C3ftyvKLyeTYarf9gAHcM+vQ3CmMtsRbrG1Aq
lC/p2C1ZvwSlRqXnrqfI5wywUwhH9pfvyYr5eZjOTvQnFV6OX8d7255l+QRMlwZw4tjmD6eWy0Zz
cS2AGaKJwEM8YHD6HfMP52nt0Pm3VKaQM7YvFPu7H8OrdZLQBb3zmmZaNOD5bmhfmOoDG6i1Y95v
GYUqMOMhjMt1vsWdKD6DrmVh0eSO/f14zTW6LKA5saz1yNTgPDyz6TbL5yTJwTWF5o6k7NDOmWnQ
sJajV/pzzjMsI9Np6ZfrZZvTU6ZoY5oB5oHfP10Kg0PmUOStl2o7g3p/w4VuMxcnvYwNAYZykBA9
d3BLiHFKaLuYSfJFDXykA8W9YbjsvZfsZI1qYRUDxhbl2RjBFtnCfRmo7KyEqZgbIHW+zLAlmdFw
m4xYJJMR3ZitIy9qc9HqhjHmll1KbdxRR5ZdkovdmdhbQ3NeAv6jecgEH9BDU4/ypDH+Xq5reVf7
M9Q1epA9cE81JTSVyny+/g0++iUx5qwTOiXGSqwN5EGJ6SvICHA3hPPpYPPAKjcX/lA3KP8Jtnov
rn5A4rXGSYO8baOSQMo+BSgDLf9iIyFN8et7fa5UMEFuXmQ2Lhdl4fKtkf4ekOXnd0uHKU+WruUc
qx7lTfku4TS4qC8PQONZwBAGOXgJvD/ZKhJJXO/zNgHVcr5zWxDDaFbX5omT5TxNZjXAAwQNMC5a
aqepkkOnghECHbmdwOep0V7kJddnO7+BQKgx+3kIs0Lyv5EDGO3/x4mjkaLRdv1ly8uN1xDTkVe6
hRmgl2hGUxbzoDfY0i5ifX/w3eKNUasyAawQQZ6pvSEN3xILePKPhBalHFoEWEWSC1VFJAoMJBzB
hU1bISKRqnX3tkftkKpOi2O9w5erInEWVKilRG3MmXHA/jX5eRbtVS2VPXgS7ss7CcsUUdzEbqe5
KGilWPLYqXPIVdA3mktxK+NEe82zjCbQ/BznC9BC1SOjlVIhG4FBq0A1SHzTQu23kFTdtzJULJ76
F1dfpljRkKR4WKrUpZfzqwqBhV/mfY68K/uR++4cYFoi+ll/MmCmo7Tkphx4WFZSMlr8qLROQ/e4
KrzjkkDEnEASec/l9Q9OQ0utnU0lKSVKykOGpMDcwNt00XPR8PXNelYgPqGzj8adJUkr34UMN5pX
chrO2gJM1JfdMShzx+OpNi/+urLXRbRXlx7OFi7lpn7qGKojbnrBIIXxfvhoB/t8FpXTvucUXRZp
LgxJ5Xtrei9yn+DsloKMly7jFHpSkiyE3C8Wovvce3p/nTkm58IC+itWBmeYSPGv2iK0j4WZuhkP
F9Z2NLJd+3A/VgMs++zsne7zoFa7hhOV3L9n9D6U5suAlbukZq3QE1y7Qxaq19TzFxZw0eZADsJt
hqA5aN+SSTwcozT1lJ6bPRc/mrxz60lML0UsWvWQZMjbt7E27PwchNoxYzG+KTzbv/V496RKiRuJ
t7asvhc/H0t/W+i/MBbtURmEeEJrt/7GRlCdkiIYwhYzaEz9xqopM2adqiLAy7ctHY0cT7nkHsVG
Mq42H7+9kfKq45dU8I5GltQ+c0apU2cPHOYX1rnWVnFl2qYjkivT2IwdxjwJdIkmmBpCw+7uJj/u
O/zdcP5yHPcPUgX4Vwc2dUHWF21hVlmLO2xOwWzKtQyy8o1bKeNRLUxhGlBtn9k3JA9jj09PAqxD
IE6U6651k96v82XorkGT6IE0LPVvPQ/oQD0cC6ioHET+1ND9+wczQxOX5KmNcuAd8EUcfQNNeA3o
OGOh6D56RJZrhCAnQqy3ckzuQdE9AOG3AZFKQ8sR2ItlPKnso3ymE0XCVDET4GDYMIQI6D/xnkEg
boLIIsyDY7zRZ00Gpva6oaCj78DUVInC1SXviakQcbrtubArpHY414Fl8XSFrAgo6pGeuxhBLckP
Jpl+1eGrHowavzfjMKY6uYU69bc05IrpsZyr0Yac2mBUIGBwdNE/IBefG3H/4u1IxYsUjNqFwLzY
QK1I+DXbH8eFk/8XiZqowDtkjl4b0VOshBWuZ6IqSQ3veDN6mlM2vOj5F/o8cdkv5E1DGmxxlVKS
n5kHYSmFBwIrDoa/7ZSgBV1/+Fh0tqr6C3VqQi50LgbBZThWQl3YY90XWyfxiXU07F90Dx4oHEJj
+kpfRxnQypLmhZb5PNl/h9u+N7ExOwz0KLvQcqCqj+JLdPfJW/5X4lxOgoi4g4n0IGkwWQYDXreJ
g/T41c6Qdb3CK72bFPbsI2IhFeb8XaMx2H4vGDIY4eJXOC2V0dRsYjrRQ8Tw7EBhqWME6svIAHG7
dpGOVPgFR0H1qokPGmrdzuvRhcPjSlKp8GIUkUDTzPy12W8OBEkdlba1rPP/k5r7ShZnTIzZVV+6
LsnJSZ7GJIA/5owVqgdOwXH5H4pBZJDa/Oqss67wzN7y3HtByb2K91rJw+jN+mBR2y4n4ilA0VK8
eVahUb1C1/VQ7a1YHohCQfyZqX6xwK0n8mjNgYD1xTM7mcABtehf4qUnDLAls9Jny1m6xwEKhUSU
4hpV3a03Q4vXWJ2s+0rzfvZ2P+BmIaQ9yMO1z3FHsoShkK6yqTBE4Te62Y9zgVAzUe/mswnQOeFk
D41eO67TfGG4oV81Aj/F9P2Wu0QhVKS8PSODQcniqMnFhJl+mM7urLNC+mLLWro+mFbOY698ataf
hh/17vb5Rmqac1wiDvLXT2O9Hu1pGgETchCIORUUAnMfhZEIqkV/YlL6LzLkvBjX0HDp2PBJmeA+
+V8TQWl3dPUIP8Qm/du/SIPUXRAnS/fd6R5ZgH7AkPJSTzn1vEX0cXYkQ04s0QjkgoX7M7nhmYaR
GqiCngGYgZwf0+/uXD6oBG9CsED5YSM/ph0GfiDigxmT2sUwWbQmBGp4CDnjtABLaS6BsFAvhS/l
DQKUF3wVZ5nlXZTJWW8KW64u7xJ+jdo6F4qEwoRreeDWimhDnSj4a2tvK7l0ZBsoLBmfHtjK3mAf
Wak3YIn4yIQ5aAvrBw8/ozF2gBpG9/vF1DijswPd8x/5c6Um6X/xINcgGVV1PFeseSobt+P5W04O
rmOl+lBn+jEdQhRotSOSZvUgj7Qm/GyJ8OaPF5b0YTlNorTvelTvcwRIH7HVbQ0+Ty8EmFz4Qh7L
M4XRihG1ajowGHzRLJl3Ct5QPI5SlVINNLUC8T0bNpble8PUg5r/Ewm4sz/GBNoDVz74Mk4A2/pK
0SnYlL7b/enJ3ZoH/pL3DASKfcEkE7dIAlyZYXrTaUiTF6m8j199Qhomnum5qzNoxYY7BBfdmnlS
CF1njafD4kFhxD0WDASaJ/aObBNMsW9Ike+F/Bvk1SaUcAwXhBx/maIIS6qZ1W+yVraUg6PdaEhs
Dis23PdLjCdCKBoxPoK0Tib/Hm+h9HnGsdzL7MJDjKlOPw2p8qFNpkb7ZK/GcsMmuwNmcvkJ+yHL
Z0d3bALAJ5Pnrh8XF7Izsa/rLBmMZtR3VM9rfB/r6ugqvrPp6BzJunkzjAAVTqXaeOdaxStt1ayw
dUKG9Sq3MYFAz2oSnnCysNJX3n5Cw9IwPv46Dzpzp4kFEgkIPdnNjp2f0HWhjai7deJ41BiCGysl
rHwKDFIDqgyWvV3J+piBVrV7fOmOuyIzZsQpxyt2iX49gMrDmMChy5TpoZty2dUHi4sd5QvPmjRo
p4ASRojGyPyxSEKF/06i6s6YjZgX/ALJcO2HmfNbSk/LH9UJVcJGEOVQJozqOpr2IkmdScNKm1tI
819iG+Ah6SWrx3bQh7kua3Wvs+SCTWQ1nv+Yjm9W9Rs6c/KPs+mcHolf6UeB/vVn45NI4Ubvi16X
gBdI20aem/4zUSLx/asSr9DtXjyaVCFdlbBFQZP29S7O2tLLqjGgOZP+aJPhCET5JEwAWVRr8kZi
gpfO1IUM+PBxo4ezq/MmK3WFCX/SmeffcCsDJRFN3fcg4Bi0bR++IiSgahyLfKvjvK0QJ10VHQqf
gt+2VE2xJZ3oM9zOPXOMNYiJIoJy7MQIdGVJqWoiMkTOP85nM3xGJtK7u5ikuh80hMrqK2kdRbkF
lA990jDtSGpL/O3d6ZGA46+ZImSpd9u08AG5IEiW9v7Y5bPBcaoiRQna85wGUFX/CFfprDNNN+aq
ixDiL163IFfAnkJJAXmYRksFQnlumDiWGK0B/Zf1DeMSOZbnIX9HN7vBiGNnwSJUO3sCpwYx8IaC
x/e05B16afN2E+jpPZZCbHNTlcbbeVSZZQ/mgFGL3vapDiN2+xwR2hJwzBPUPYN/zFQrZbWeFlrB
3UTm59vJwDG0Ex12wbj9Kjs3/r5PX9h/W1eUmZ9u4ZhX7HwgLg4BSpz4rOxPIJTyBbzzLLLglWBm
69TBWG07svo3noZGYLUYjMJCcBqFqac2LIMsblnNNmRlwjs+lJUe3CUCiA9DyVaGmLuAk1hV2Aah
TPMhCzBGLJ0dZy/1yLuWBwXtOSQht+gGBqNMLcB4WJS1eETV8XPR3Nt9QC7HxYzC6gZXz23yKdmO
G9LFEEo27VxG3VkvHlPywO3GG3pyaNr3WprQ1VHd0X83TS+rDnBGiehfCWLR49PpgkFdCwePhyXA
TKrcVAiSYKtSwrPw/gmXjhvLtzpmvsvAfMODm6MpgBXAQQ2PntoljXJygJFYJSAs2Cd4ZvgnWRgO
L6gFqwTqbH+L4HMZWWjANNwiii3uAiRgvErjAK424LzRiPq1PZHfrFAybMC158UFiOb2wOoeUdSG
obIq9i5ITUMs+siAOAmPrBZV8Zk01zXhH1EGVuIIYu8H7pRa5l2eA/xUwM3agUZpEdYM2HTywhNQ
MXb4CyDP0elctG9S6JS8LtvJFen3b+IBqf2yaG8u2VirDB9VuFI/fOPECEh+zvL2zCeMLnPNK0t0
RSdGz2W1PrEkfJ3Yg+QJb+fhoRZLDTLrYiZbl31tsbLxu8sYtvpyCEZSyKK1R7XfIp+KzpAMGRrg
xr5/5kGk/ancCUVgFh/MoQyUwNAw8yW9Af9Uy4d3nmbvM0LM1g/7dDznHZ3wxDNdYFAV2hWVdd5V
erDslP4JlUTtQjokBHubYx9Iuh3pyeaPGdLkMCqPm3RYj7YxRJ2yOtvUwprn5jgmdwWOHVIRQhmF
b0vOlsgvW9hIDkBH7qsBJ2g/SOZbO4AUnhiw6IzrNf+/fjq9Hmn0Y9ih868QwxIR/UuNhuuFVaw3
50mg7O1Ve0pGN8jRdos1LBGhvM542up56kv+YgRgu9iHma5hQItntD+OaR5V/tv2vN0AhrZUjfk9
NEIxeUu/+/KqFJQUXVKrkA+hm5129KB8I7kAci4pekJXNXE+7GxPvUbN0yrrSj5Z+XnTV+Dh0pGP
v+sXP4cdKnaZhL9boF9WujQalZtUGw8zy46R8t3SlwZfPNUVSvELRpZuhRxUxn/IRsff22E6Wycd
gSHdSPPL5xl+KF2a2Fr3oIOAv8RQii8iQovWAShvKNlplCrnxZP8faGx/VLjG+LJjHxzB0SZFGiI
m/2KwclZxXp2kB/KgR9V7Pp4u8q2qRLFPsj4GtteuWn39IuSfOfwKFQve0ZdwHMv0AJ2LseWOL9A
yqKI4i/g/n2pMCHZBaNhZ69uAzcBs071tx353vvy2+lFQRoJ4gh2zyWm8td1AC62BFdb/ySZwssk
AHZoRPdXMUMwo8kPGeWgRITCGdKaYZDzmo1IrKJqfNiaeciXebb/whn7i89df1hU5+oGzcqQGuyP
kqaXHfNzSyVdO3FMGWgeFIlMVUcdoD7ARsy3o33rY/488CU0j62IN9/7tv0/ssi7T3ZCLpHJZx+m
yjbne6O/ym5mDDcHBGtoOJ32a0I5hfTUz6RAyav6fz5yJTkH5hfj1BgldjG3h4OH/PE06seggcR5
SPkIjmve8TvK5KqHe29tdct0kDT9vgCd0j1SoL/lA7RBixmSZQgB1/LSg87JXzMjNkks4mTX/gqK
pIxmq0Mvdqxki5mWdCms1+bmBYlqHag4tdAoeOGMahqWU3eQ/HeUCnLXMMDMGavAgk1xl5hPNeCs
yZi4gu/mIsljiplGh9CU+r7H808FKwwVN0bBsy5rh4pQM5NM73TOWTHYz9npVof51zsWdL7/tFnz
kGxcGmv2tiwd52i0hh+BMN++8XuRbDNH4G+PjZ8U8XuPDysNtN/iGTnermF1lYPLgsZQQodRYbGe
aKfdO8sliHbx9QRKnb4RAUWeL7MEgUzLxu6jT/G811vJ76oo9LvD1LmSl05clSDZ5c1/1Vch5rWm
uKuvIe2UFdArT1J1rVtcef1dqoUiEXhfmxVDrduQ8++0uKo/d7yVfgEb3WfA6WiK4Szc3xACYeVY
hYbixokcpNsKEq8/xNwk/47rdjPAzy00LuDiYmZy47aQpY7hLWk5gDwlF7LBLWx7Z4mr4291kn7r
gGdJoQodp0yjAF4XDWKWFscfN03kRdFNEL4a+1qK3jUc66u6ynAoV6CD2273ECwBXaFVVL6qtpZb
yyGFCZLMpdXnKSRHSgT0WhetzcQYBpFDXNYg8uLNWYHwGWoKPOx3RwP6cl2P80I4U5KtyqYuESEf
cPxrHHw6gAg3jDeFpqeuXl8J04D6bIoNl3LtB0P9WOz1F+guV4rYvT+UXDUS486gWWwDaRMMfOCU
j7NPzgDrAgjLaWdh9708Uq4rK5uKvt77tDdhHjXnzkHs2ILvZHMHKJZ9ekDSqjJJ6JkHr3TOSGew
WK5kklukeraZbPIbWQ7K8q/cA33ORXFaG9Aq07RQoYlMAI7/9AduBWSrWnxw+VXJJHtWX4Bbkopa
/s3zY5DKzF7U5LUj9cm1knVN0KGPxF22VUd6aHKKrrzAB2EOXjXd9NP94K615fgW33L0crUVjJmV
ug0u79Tqaf/vmTDnoa/n6U8DV7D13kdLBF9wAFHSWVr7fFvu8+NkKU6f2MPMevf7l6IvMMHBzu0G
fnmEysQdvIs7qn/LmYcE6Os2uGSH1ms+sMSosygadt8D49BSKYo4h8GnDUy7MJHqdeVXUlan5FNy
rnStamklF+bYFx6qakXfSX+liPBwKWiVLr5JE/TTJMfBprXByPnYjQNi3GSBoGlFSPBHxGPUKeJW
EPjDZ2oBg+ZniQWdm+Mf4DodeFEQfwkAOkgPXKI9zcEzxnV5UNwkY7OdVN80jpuiZatpyKwmqNKV
EHl1Sat70umfG58MVIpAnCOiyDXxKHF1StK8Z7nGygo+kYryEe1jrkHY4t7MDzEjFvYaUySSzdxc
+frVCPat485gmlcB3lHEqdOhxtWmnONGKDOXwr4obYGcG4Kryh8NXPvAawFZlT0qRjnr42FSnoKI
Zn935lTNxqqOGrLtbglikXipqKWy9SUIqMGGr/8y2PT7jn/6M0usLUv6zi/WVghzI5xdKxWt85NG
u5KAG7gyCm2vEHg7GUL+jaQdz5qhfE5jx5VFsnAsy2ykIGsCaWPz/YCG63uDxqSwvZv8VITDmnop
8lf6EUyrWPUTTIzs2ELVyGFL+PTuRYJI1w3V3Wfp49DJxZ4+BJKOAqng5G1Uhlg02dE5xtRbm+RU
iKAJciVXFuCsHR5a5PPzi4Mau28CIFQJ2N/KxyIrtPy/j62Qyqz/qWm3tbVy4RDIB7aqFpuLQShM
79iyuBXGKLuuE94WF57wK3AZXfYz5tLeeRQY8M86kVPh73goxlkMm7pKxVRysbJMSLW72nJxaODB
jV5wo5CEeF1HeRtHm0GF4CJbIEXArvTGfqyqGc2HiKPjWHRb0UEwoOZOfW3gk0RBaTHRaY3iQInE
YAARBo/9LeTyG/qPWFkLbNvUYHaG4RmirpymqSJOT7qLkmG9gOzL0QOBncf6z+aupWi+NoF3kOfm
gw6/z6y0hTOGK/YMVqtYDooIFYf1wOulL9AjJe3wa9jcIwqsiaWoJyoyUlW91zBYATHwRYsvAhu+
H+L8ZzEEVxNRPDQDLlOtBw9X3RdRrTW9S1VRPnhr5RF6K5CzyE8qayIYJP+cs/CqHNX0k5wuFmv2
PTxkc8UWV5DitcAiULESXKWSNIGntDeWtX6noawgODnaSDcW/Vi8nEs2Xl2ZEjmzOoPKdqnmco0N
vDez+QmooASujldi9LpDnyOiK1YiWw3F3+6wRcsr4dOyGA/ELpUYZHego8C90rl3aZMOBhnDGepN
caNZW/4TAByluB584+XeEiX9Msb5p4YDXLpka1vjg2ca78wlrYIdSXAz/GoEKcWYi6cc/0eOa1Wl
71gqOgNXez9sGemTUQA+25SfQL7NDvkAcUx9fjnu+ootwYtkWmp3y1HfGKQJHxP0Dk50fPhBUfFD
N53nIHpjfbCGk31X1vjNHgCjM4TR/bzRAJ1AK/B2TuqV+/Dt46KTqjiRE/nzTq+7EKE9aN2Nxyea
rNM4MuiGIIDAS1B4Woj9FHsI2LYAFlInfVaiGkl051eowesjDVZuF3Fm4amhmj7G+Vaj+5cILVqL
qXjQPriZbwqwH2Gdt5+E0mAWi4jmLVUaQE/ldpjJt4tzUy1h6kv0AXQRklZ5zNCzbbzXScWxE//J
/qffu6IxRy4qZCGmn4juvXleQpat+tRZ8iENqPrEoYWF5TyMflZqQz03FKBsKHAr0y264LY3VzwK
NnL2xFwE1H1e56nBpHUwle1qcCw4LJkL8l9HJysgG2CoqkE4thDf8+i0KbG3PnJ0HcelqHN6RO1x
osLgeZNjwy3baqdJ/3fC+f/A8Fu4aIFKuqX8NwsjD/Ytme9vbE7BmvqpgGmYYlFFwqd1huI5HC5+
D2Md4+dWRcyJzhp70c9haLejGjhY/Wbqfoeu81SZIxheQwAP3KHr5Iid4xjChzuOqbnJgkPwA2Y2
RcXGPNSsO0sYUMNed1JzBnT+Yk62eJWRidrV1LJSVRMiUHBHSrjJE65ioQg3UKzJcQnDv/P6iH7J
S93logOZrWh9IQeVF7F/CdHd11XdOQkej9F4jJbkSuGJYdZ60+iR8askODEEchTouje2reE/c8fO
0Vsmm4M2wbpHWzapqARr9g68FRPrCizZkiXH/Kg1jdq8eB+y6oSq14A44HE+sxA72khAqbRdVuzW
MLrUjoHc/4gp8W7pdrvHkT0sMCU391Y8GK1AnRZJ1hhh/FR2Til/TSLIaPsX3rYIn/KbKgcrCTOx
qgkiwmpXzf8nr3mmZ+0JI1dK2zDOk9vJKwj+KO37zbDi79KW7yl7FAfg3BTHcEIYXfasdW1a23fM
laqep/g72xtwsHOBcY1VpyEDJ2vxk7OG+copAtT+YBEB3CVQsWzw8GAI4l/yDF7z+Vh8eFeiuqab
wrRIZ9DZ6a0tRAAsaQ8BAQiU9tpvCF7wvyDhzeBymfF8Cqr+uzjwIYjDQOKkLWDgDxMxdbde8lqm
AtqRetUtHq581Rv0kGKYzrpJGfv4ycyHTh+DnBN7jRtQlfmGskAs1MUE4JQD1PeGOYaS4g/kiaN/
Ua5BmTp6rCp9v5JKGaTXl6XveZGtJv5tTLpFuxa/68vJepduVLZ+qq26vD7OR8SCoalYDj12BHIJ
E28Uym82qpZqstUIws08G7RA7u9RdTCFxLZNimbROK3xGd3bGkSMkthF5mGPslpMDwpORxtW9Eb3
kUGmvFteE5jay40oiWm/R3AiOv3Ar/LJndSysadMri8J38SBkroB+pwcWir3mXRSfcNE2C86FLEr
YBVetHYg/xmofmyYfcbI+jFo8TdtFuXuxdiXVT84HsdcXno+e+uxXm+ciVeDnmKlpd6BmAJ+wbn4
dahZdVMqpKhmhjZ/qp2DTSTPoZNp28EZZLa+gDKW9ZMlIv480UpXTxgC+mvvJZK8z6CZuiI9Z+FY
StBbFvZ/GzK3Ju3MXjlFNMNoY5h9mtISm5KRt/ymLK2w0PZasYdu25EKR5bgiEgE1duxWw97VrMH
6r4740XHAuFtdJCahd3jFQVU3ICPLGsrHHpU9BXk3KagG3Lq82ReytvwHfgPbBzKiZFjVknLtavn
ugza43T/Bfnnb+SEZ+n9qZGZYyAoxmtfxPGWAUNSLopPbcwcoOiqMCKYwR9/GCZZjwgQ0dgzYRA/
LZResnW4fYcBVVF+ywwkrmDkrpcrCxg0Txdl3yvC+5WEW2IpnQQOMN1IuL+5M+lJt0HAON78CW7k
J03RpqrzENdW7uu9jcSYbCKIXfy1J88uhUCBSvDLJiRFBm6PoeyqNFI1QWw1e0Gg+4X+LlFxasYQ
OcazctMMEj8b6ffWuw9f9l6umSOZ9oe/6F27EoNyzHJtK8vM0yN17Du2dVpyJ2BewIVEAZwzkke1
rpQwfjaBneiq0igB8PLvGWGz+dtEnE+U/LrBMtaJI9i7X6p2xS/lujcPV5eL6rYA/UALDsZ2KH3V
T45WlACR2+GEdgJDKS92qCf0NXIpDwCRRCqe9DHwJR8FnGHDC6udn9M4HImmALwyqXLyAwczZ1gw
tJs0FXuyvPLhVDTusvXi2lQf9LoqchvXGNMvThhnXi2T8PUg+s4zCcA+xjy6Nsx0p3t+LQXU6EwR
+ENAnRfsWIFWE7Y9Q1/7zsdEF5Pw9wpVBL16fgZQ8W8997jREwd2NmSQlhKHsVwYuSteHeY/buUP
/kM1THL1NukIa2WY33Qxmjs4POC3vmhYZ834Xnzgiav2+WXSY0/XBS7rGar4Lu7x+0uxz+U0ppPV
s6PVr4IrzZ1pb3KVUK2w7f297d5yFWUCsg3u65Kzuq8I6oPoHc2yfG0Mmix5DuembL57sg8GrGjd
ihKyQoIfprFVJ+3U04zk17qDVkBw8DZ4GjqVPPT7w8Sn85McyGzlxHrC5KDtMbskv5UNDx5ng6Pg
Rfg2uH8sKSVZYsmIoEAgmWaIo7KGPjdFkqs0vJseLiJYO/dbDvFmPm6hisGQptbqcFtVcyiv8fCx
akk4oplxejg23QapwEorXNA7+BwVNi3OS4vzsV3MININbmmvTCKwDHBfslWEZ1WiwocTsEaCRp4s
cNDdnmZ0RxpqloQoPecPQZWnw2oJgp/QJ0OYWLDoZbUQWmITp3bRPU0yioydSFVvN6iDFvEC457C
oQUW9PwGv8BdGcUrGdjIAXRL/dX4cQF6S9aRtIf1CLYVvJV5QNlZSPZoo+wBSIAFscyOBQuwawti
xuTxV7MlzmL+9plonaBVDHbaFGQ57QoT6sDNP+DNQrOI67W3QFAzpKcXBqHoT8E8TugPyJpAMInS
3ozIL0K5gozv0iveH4SYTxPGVHKwN4upKslxv0k31YtS8VGhNXqcDHKPa2BpGhi9MdK3e0xRNxUB
svn84ApJnqxuSJH3rdKAZdIfZiBrfbgOflv0sfG4ZYtSwpPjoX6as/S5Vg75Phr+7CfSGS6B+Sou
ZQ+BNXxLDWvJ0OK6XLziimuvwRjEInvAcGWggUYNZ7HRG9fcsRoD6kf3N51SFE7rsplPbSoYRrMO
C9eQwFzspn5kpaPSvPK15n0X7DgES4c/8cE4GFXlZWHx9rdbpfXpgCTyEadsyrV0hhu9W/URmCN5
l7OdUVZmMNKmJL/+Opmp5KPzxyGf/JL59eWSgF8HvkXS3aBudgUc+wcNEZq/nhfGgSyx02nFctNH
3kQdxurQasDM4oCloPZQxuMqfy/mUrS2TGEwE7gA+7Cuqq/ILAtmfaO1TzgJ9jVlFcHQ4V27YNaH
0fgOasTXX5URiMvApL68VBrNdMdfcJGyKkksD+AurpKMJyURXpqxjukczIlibkR/MywsCEcNxuAD
xMZ+g+rwYFxmTctbB+Gn1EL2em5gxvhbJtOO33CmIppqFDYl0VPCpqEYV1LkDbFNh6VIEnQEn2sp
FGMKpjto2DUjJ5nPU4NO1oPgLBTq+aOSRgPRzS1DAAxOH53gpeTflYqoT9i7xasyRW93ilW4mGer
vZ/lTnhXKD98R6Sp8ZmTZ9ZddSKEXaJ5UGRjiviWpSAkY+ag9LhxvEWy5joo+3v0F3/y5MlUiolm
ug67Xe9yOmY6Ilr0cEoy2QMB72G8XcHCXnE7ioADzj8nb5XiTIw3+oEwZlZFsjQA9ZP1w8p37JFa
V+Lf/gWwVSNDVAPPgcnf8h8FnUJmk9z/oGPwDUj0dDVk9G95Rzjzc0/Mlqeqn8Xh+Lm8xZ2sO4pL
89YgFc8T0uTZNrzuJ7IsipS9aOm/Bwmue7xufnhIlx9uibenoyqoSpFjtQH7rSCAM9dzeibhuV74
8LlHP/Oi97k1RTQrm4OJrRV5MZv/WjAuqOA0Mfsalcvon00s0vw1U8nWdObj6NQmsEkrbMcFyGmb
cnNSHyduqEvQVcYbQ+vG5OkFc143TSPEjGm7+V+pTTzOLHu3qPE6flX8NzgOexQo7hQg93HIQGB8
WfdrmeMX4kGevkfS1tQaYAVPLYXI8iDwbBl9LM2nLpGVGsyYww7m39ez+GWfTwcW2nv38u5/0CBi
WNO8aSaTPDcs9NgDUDWBde2mlg5AEqVM8p/la4w5eUpwPQW6poCvq2tLc+LvzDPv8eOyFjea7w2l
krgKR6pfJR4KSwJYTGg9cn2V7eCU9+QaPPhkuw8N4MSz3hRTO3sztBkTJJomCY0bQzRKzAtl8tqc
Qu6ZDYY35gLP0EFoloKonFqzbcXejodVOxTGCZBU7nEMR+w3lKDk8Zd3az6cgaoUmxzSaWkjzSpu
tZgzw1KhZ2I7ZiIbIdKcczJmQN5F3yiEyredqE8zd0t+CptcQk+wMxDcM7oCqSSCTD/kOtNIxHa0
zhwyMeRWCclBceRbYsfS1pJn8O7n0Zb0mP2tXdwniDZwjnFnOHSdDgKW2tTiyDscAQA6MlK7ZooJ
SMgTV1j6yYq8XKuaaGXxHiFUffUPqRd7t019W9scOazm4hSM9ysPwfaGgnW15YVx/8/Jymy85lKm
9VaBRgjPG9x/+5ed+xSKkdRY3xkyb1uB/7NiCVohykYrdxdePmFyawg74hNPJL7ln1xNM3apcnDj
Jv4Qh/n4ouCGRAOasCRrL5uXal65sf3SQcpD4ltMaQwNRgwrMaCHrT/lFxPW4lDuqLzywXHufsJE
ztzouWMVkCZ9/YQSYI/5rbqdo/SjgOmelWjY2+vF+iawkiV0WHoHRuvQx33QnvESAD5Y3w1AKaNN
AyMxpnJjD0TmqmTTFL+Y/W+Y321yQGWIZPGwEdsKsJESl34r/o2WfJDEnL9XlgngeoDfpD7KInTQ
x1jWhB8UGxjn2lp3xUSLtfs0H0HARyei1bYJtvpacZ3v0tIkrtlA1dUm8gplYFilUnuJ1iPaQO/J
4digqtFzOhxfgRIJ++XC4FmppKHbuQUQN6BZcXCS9YOr9P2kd1OQAIzuoxDdJxFfShTLlZIxqTur
BOIw3heBcQn4h2Md+Vo3ECxi5lEVAUCNJPiVN5xWvUcu850SDnACgSHIKzqJCWFiJ17EGVzQvAQH
BuGlrHT1Zt6e/Y7V1dUUfUnERuwfvOAQxhuHLLoxv5EzshAibiNFzQMD+iAf7ySGKEbJS2iYPmVV
XgZrioaABnpxfEXVIFwYYkUeiKYtio6VuCaNHqqmNRbpD7itvQOlSg8wdPgdVkcwxpoulYTZLTLS
Ly35unZYhKoI8MTIacIaTDqQneWCjEOy5wLjopD3IDGyq8BcBhydpsL80jc0vUPJNkLgpKPyqQIp
2zwskggbsdzWWT0eLY8I2nNYenUWnCipozrWigQTQ4ZCB4b9zECeN8aF7psyZOiGrjjYnejbJS6J
3WEs5j+pk/mNobxfcpTq1bGUBtJ2fKmF4SejVlg0H+Obc9XEqoVRkbr49YE1Ct0VQJ0gUtXDBPha
43QTEohK0G8RpoLTMk96pzhLcKmaDNxoPCRpbjvW+SREp/lNcG0ROfOe5nEulmPqIPgOvyOJE4bH
oe64si9IrOFj+WUM4HFMuSRn6QRn3ytcTIsOnlPisbnlcjtT0tRhEQY3uVUohCV+iK/3KeEquk3L
okNpzU/ORsp4QEKlhMx7R7EFqAeptnBk3UudvBGlnVAvURl5iBLQSfiNNFuAz62jK+a//wbjgM3s
d5GZPUjvHyKlSnWVWQ+qxgX7ypSxJTk2Sm4ZSKuHWSz4UPtdXlWchVTsrO5N5BBgKUv/T3MbzN+/
jsjSfuNOW/Fzse5x/+QsiG9z44YMNQd5iRhLaEFfsg8eHDlbkXhDGa6GBYNM+OmBSVzTsuy0RBn+
HhZBsXmFcRTgnrw1yxFfFL5mxhXNU8CCm0VZ7+FhIqmmFjRl/vCbhAy2FETmGsUFhRDBlep6ABMJ
kYUuJ/yVRSt2eZT2ksvmGpBiTI8Or1E3YuzkAaWzwh3R1H+nle2HRirGllZkc8IuKDe2ymsyOwWs
LRaH7gz62LVb6qguDjeTmayFifzFc0uur5nxWz5/At7uQ1iArqj3QQc9LoM+NgUYDQpXIC3pMCEi
f2HOVmlmERue+/TUHXJ1fXJKjzhSGrIH9hAgusYE8fBEhsR/cNaxvhBO4SYQcwtHsqppbp32j228
ABV9yD34mywufdG30jv4SAA/tyVCtL998ukKmd/1qNStEDHjJ+UzGp/wVBH2I5Z7cZ8Ep+iFO+B4
d7RrEHZZG6bOfNlaaqvTlROj1Df2ZuJ6KQdPnIMn26E+j6mmiSwNvd7Bag0r3hlsj+J0kDYznO1D
J1WKWdbZhjhdoTEFsmMlVpxq2Gq00dl9ZMVeBPh8l/t2hdXRZW4IrW5QKCvHgKqFyQWtuCXXTH4K
1+Lki/XnCb3Q8xWS/rwTvR6ptjBN3zyxcly/yczwCwR2OdZEHnYmkkAE1BHNZbIYJ83XJnuLllGN
DJ2H/wjwROt8k8W0LZVfFEzFeMBLivQt6P4vesNtXcefCtZmKTLpYjZT6Ot9tzA5jRF0V0Pl9F9K
X1YUewkfhth0KSDJmVgVr5txjGYBTQNUMwCKIKWX6UI2Y8E2MnPoqH0/MWYvNbYGO4T3OsTZa1eE
/uqdeum+rNi6v8wcSkZ1FWY+VdRq4sTcsl+e2EWtCi2HeXqboviuVCeFhfqBAjTQLz3pz2mKJLvp
6bdBJeXcazwsh1RleA2lCzJAB4Ilgo7TuV+L/ZIDhWora1QVn1Idy9Ag7/A1RphRVEtNcAu+prL9
I9f8A7jEoOlc14V0gJQZrJoOSef/NKtHEdrNVasflPfkLsL0i67ybbMuwGo42fZPZuprKYOZX30O
wdI1xsG0zoes1jIUIAcFLbooNKOmU7Cv/le+gsvLWM+seBNWVyQ3En6vQYJ1onF10PvLIBhD/jYL
0apmVBw075Sw4/is0FqKEOIEfjXybIIZbjYcF+Ug9VVTYkQmM/FxbPTp+9QB3pAibiTqVBgqewl6
uibx+gFlfOw3WI9H8m2N0Qbt/O288xiycU8XVVYmJviI20rSvvgCCaCoP6dTeb0F+b3N/8euJlwv
D75SJbvJ+3uL0MtDGIuV0HbF+nnQQGdrso9NoLKNNCqMaxGGiTB37+mb+ACV3xCQyj/U67qeAy2v
0NDxjcZuonCmXlmycEep4V/o7cP6SImLAtCpWCgPtASqvmJQSbfXHLwrzZU92kieDCOP/XOUO9wa
JIT2I5ptuCH3l0aTQ3R2MK8bvkxHPNSd7WvVX/Nxbo/FvDBNu6aOLjkO/wgH0PCyVUBe0iCFeLI8
6mCwkPnd5C177RvtCXryNmmy3zUsxDUgCNUnCd+0wzLGH1/vdJ/BlCOhxsDvl4CPzFYN2vI5vkqU
XOe/xxTQzvKfoiCdVZyM4Fx0vEI/H0Y50B/mKTW9stanYg2wbqpcidFL9SRuHQEWZbyAvpQRdaqq
ilcRX0ON4L+V4INxiZ9B4YHqBT0RqRXH5hSvFHmXNlSuvMS0iiD3tCoRM2nqHEQqc/tLitj5KuXL
otvpdhu/aXpHIUIaTIFWqKkpPa0GikDGE/repm3XXdpbfqhey1P7Aets3upLUlj/6+jmkCVfZCPM
8CC+wNRtnmGzuuz437YHb9AmPtiWYsfZVqtON0Vfpy//jiZCyH/Ip9JpRw3iq3MC5nyleMT+/cW9
4TEz84JOK0YAn6rkaGk+4atQ9DO2M5EXQlYG+yCcf+wFP0rbgyZRR7UTjAVcUZs/jMU9fYfFXdbA
Ut3t9f+T3ZfFtpEIDyLE15fMdQSUUsSKjWMF9dgHcD4o27MvOkTluc0irBbJCQMpT2pGuPXORjT2
v0MlxcR5jtYfiL94S4Zq5rQjNHNp+t1r5pAgjgh11VeRHNGPH0RixXkd4i6eVFWp6Kydg3Vb8Pje
TRngO4Lis38R/dfj7zfbsFX+6DF6Pg0E9xnQJzxlZEbEe/FPKG4UMo/7oqk3c+Y/f5Si/k5a1OWh
wBTXgaqmtU424xLQfuW0thTwaC7NAvwV1IiOvNGs3ztjtaygKm/6Z/hMtRy7n9vdHg70oo+nRR53
cnX+IEtXnmhITHMFqEjv+w5K8ornAU5oH+EoQ7bTeEcKw3foc2DtkHdj63LFs7HYbsYvpzF9+Xv3
8hwdaF45msi2jDyDSJPYqmaD+cBAlZ7kRnkvaBzOS2xqHLFn4xOlGEGixMiOzRqPM258Kcltvjy1
s6llAOF+I6sccTeO8qg4Y27rGg55vDdNwVYPMDTKGpFa6vy8/NbmUIMXLGK8citM2Re/ydAR7YjS
hiCWYKdSaMST3F4Zweyo3LOQO9I+bIg7mb5FjpcLhneXGH040X1vMVLbttoqa87FuCcq3HQ2T2yl
rJYv1tCfEzxYiQo0GZsbuiaTCMZU7zjzJW2sSLyR4n+E2fojiWJ+NRKcwl+OODQCzCXMJC8eNBaO
R7dnzAxbkDiGszeuZVfL6VkudTkaGs9ikIdE5zrtiya5FX8p7ftyzw/pNuMM4hzItf+0aSHbB6J8
+XoY4iIrdMTcHUygUtEzFwxOT21eeLM/wZxTI/52hgVlqBXt2KLh2g154/lFO0cfrvtxWX/eeB+U
Nfvxdq7X+2HcFEefNJlV3WMFp2xL8z78ucjmjq0TL/0V9y/7yW16x1I52YNX9K9p8u+wcvFEo32R
Fa+o85gGOFeJvYPLuuNXLhMkb+pE4i6Ya83Mu34PIzBc3db+U2+LecTFJtl3wrgnoKXXd7dU3LlZ
8EOHbAo/uRHcZE989Lq5iimnBkUtZqNncbCNaOImZY8BjZcbMMeRBlPZFThpcfY3wT/VHEzG3RtA
WGEo/IzoVmxctW04NfNZtQHJYr8X09QsqIrjGmWjYqqNIWHKMtnCTHD1A/F8RR2ASzeIprIrXP2b
jpz4D+BtmUnuDuNnfk2PO2qM+dVI0c/EP8izdFUlNS9DcYZ1ISnd85pMaPiMR/JvDT+buRXylkwn
DgAdoZpAaJMEDvCrHJiAOOFUrVC5uuW0Ffb29mOqlEZak9n5pN9encaUDa+QTCjYuWbf8QvFvSTO
mI4hez9+6+caSXG1V1euGMsXHeVz389GbKaHiMI8sLLJW8ASrL51TLSBczDbFYQH59+uIN8amUVh
rfAk2H+maBraf4waRbzZ7YZWXb6vRuAkKv2iwkGpoNdeWjC3TB6CBskiqgj41lVD9wNKRR9h3rKA
VTICwg5l2hQbV+kugANFcTxtBahTZWZ/lw01x8i6aQoW0iJ9SfcJrpyn5wLeq5YyPEgxoJ46pcJk
j3iMMVqI9vPrNp6cqVOZi/3r1qO/GvDVhhb0L1mH43b9nygNAimn2uWyJxemiuYDqSOj61Fhbdr2
S45rDwrlhJ0SPXA8ypGPsP0umlPQ8Px8HPiSGp4crpP1KJ2D7x/EHaTlJ3yph2UIiudg+Dh+vR9p
uCLPPSMMTQCJcIttHWVwS4xGYy2TsOCkXqgORjrIXaP89FTUCac9yK71WCi5gjvoHEmylTzvjKDw
B8RrCOtjHzdJ1NilFyhP+39MZ9i6lXGe0QHmtn0NQRN5XlrmJaMD3ZGerTMV2lc7f3c/S9MdDdW5
DrxOdgmt4uB654NHy7+Mm8KfyY6MJaeu9IYpvZ1nsmnEhemnS/CRU8e/d4DM1F8StQ1vj6Nlm5OQ
KmXE8aFBu4blogtjzJfKZow9r55UbnU49Gyah0piYvku0ZfIJHzkTvE8cybcxNtH+o3xkfqlv5Y7
ovJFuMWoOrR7y3+ZsthaNWOL8PL1az8bC+ZjIn3uCTabV1XmIFlF7JLd+LJKaogQNWXXCSN9Mnhw
xSLseHAowFzulS2Jl3trvbgTmrTbBReZcZoVWb0K/elv9lQZQifpGtAW88d39iY6M0CYvQvIKwQt
L+dHuJaCiTbgxZDadMjKKbVz9JnFXcOofs0YoxMZ1wPFc1VNhwKBaBv/Ntoe16KV+VQo6GkGZNg4
X0ak+cvhmEci4yERbaqqIbY/8oHtHG/XVrrwe+8NcAT+B+iTULAVDg+XRxIWU4bxrodXv/JjM82i
Zo2y6j98Nz0irmKhtPIiRBSxJK6FK2sy0nqig9U2GcP3S9b4VyGb28GeB90Fmv9s50YOyIdNi8sz
kuZpw8IPW8W5OlMD98g5pFFDYbni435sBRvgf9YbPFesSp9VAN4jlgnxq/qsaAnWQ4JNxHCwhuLh
yImF8zntptP8q2gPlPnOnX6iN74u4KDlgYrAR6lLBy20qjWk/Fygwuoko9U5fn4u48aeraNeCV8T
ZzpeuaBRAxe8tfxfiYsdzSdo5ZBDpwgk/sgxq852TsHfXjb302YN43xhUanuoNtBp/t47GF3BtEr
5EkE/1saoOxR+iCei4yUMjoLs7ieg+8JhOvG/vmvtVa3Xta6IahNp/RzQAP4Xoj0fgcEAaA5FKjX
2/amZ4eR81wiLtVui+t/0AlgtOrpsdUslXi9XoEM+IdBOboZdzbmSM7IHpxFFGI+qhr23iTeZhBq
bUYSmT+Q6EdIeAZ36AImdAAx2RHdmJHLYvvdgT3VDHWBnSKcuzqhTNDVnZl6BO9mMGCsfmHRQH01
mhw3CUBHeVbynnNFBtnqEZ0oeAV5oc6fhtnxnR+veywOIhywRAIaa5P5zw1ny4/7r3GAaXrDBp60
/QaDN0V6Lcs9uXNf/9VUMOn/ej+bn+07vL393WZEtggthvgiLUQnqcUD4MllcQkiL/Hbl5M1Gv8H
gJB9U589ZBkcjoUQOIwZkGYtp7IreXOrTQfmtTAjesN3DR3I4WeKrVUzdazLYhca7yZLT5fHau4O
3cSULOYLRWOdCeq0jSMAaLfQ+GiWXoFe54u21+9WsB9uAYTJctAaMWhAuVS9X5U+mIFp8uebLym4
uAh9b2Q54TQhsurD2iBDGC8nU+2wGwYyec6v9ViveK5U5hqwzVHs2k/A3/5Z07Q/yV6BBSpAcKCX
3QLGJ6VMUmzMKWyy7pUYWZKzfz8h+6NoQH3vy13/JVZxRfbKtpC+aATwEi6yTn0A+y2WLUjxHFvT
8ltAN1vpX/KtQiSccpcZCqaSUpumAXISCJFln5DKqYvdh5oaVIAWIx7hLQPztll+vyXh89MgwhLS
bQaGptZTj9CcgZpFEsdVdDMq2TVZoO9MDynz+8JPaOTrLLoOD95sj8xBv2x2n4c+J8PPB44DLtCM
n9dsntS8CGFgMrItEHz+mzJ1seXAvpsrkDjFc9hhQgWV/lmFIK0Nt1DkiXQKmj3CnvwT9N/sIkfp
xvtEXTQC2wSXsu/gCaM/1LpIRtaRLot0sww26f+jjtt/q/ZMgva2t6KrtY2MqBIqqASNOWG+xy0Q
N41wa/qPDukUsZ5iKq+wNbCI6lBLd62678NqPF+jWs6lTV+sqbr13+2ABLe5lQXtcR60VGS7FGeb
P0zS3UxJUSqzTCwAf9XlLvq13fVNYWwcH5SyWp52/mayCMed7IxASNZKk2zJcEkT//6Cx1RcMqxm
1+idLd3j2NIx4ZRCHCVziRiq3/9T4JfDK5/IYN6QNi1jLsK10d6WTaJMkcMvyy29+u2rNWvUr9GC
xeeNCvrSyvMszgY+7J+lXde0PXeQtJ/+HA/ya0B1fEQ8ipROyE0aVNX4x/HvT6zs67cEgghvTLVS
+RJFZ6hSLun1cUpfGSGkzuCjLIhggTdmkNS5uHGRSVsK5iyVQK2wYXBiUAaKqJTL9vRaw5BntiQ1
F2frBGSoNOO9//cJ82RT4CdXb+UKPxhSWTTwDL16oTC7JnZHQCYmcfVLJEfClH0bYvVAwWtMt6N4
irgHskY0OxfyIg5q2MjOMZKcO+IJsxKPdQmO8pNz+uMUtSm++Hei1xK2RixAA9dY20/7nV512/uD
KuyXHDUp1BVLhIqFvF3miazvIQHhfwxi4r5gQB9Zi/2K5XL2Ikxb/3a4B4UQSLOjXPs/WP51WjQN
FSDGDF5oQD54I2tlsR0lG8yW1X8PicWcTyD+rv7+WdXs1MtXE0477IcxtgOunXoVhxokIL0erntj
A60pbRD2Ui/WLmRvqB1doXqkmDfxWXETXWoRk7ssWCWKH3uO2+9GIAny54j+6nemXGYHoxk3q0+0
c/wHOiw13SvFzheTw4d03YI4v6axmkR/lWsgvfEEg+7E7gP6c0DJCfDnoiM+TbS7BIJjB0gb7KYP
H/5SEzPAAEZY/LN0meVqMjlu4ETBY+Fwpgyp+P/JYpdMCoZ1Z7tJr3z/Xj0JeuZ8ae09zCJUEpqG
iQmVYZ7AiVNWPbytHXVgkVoF5VVMovEBoon4k93L0K9SFc+JWeFlSI4Urieq9wcs6tiXJaIck+EX
gzky/mC9VCdqpX+nlgychyGbnKKvBNMVRke71GAEP4WcibtfcRljQWza0fjdKTL0LbQyYSFgHlJH
hV8gyROp8om3yEtFckMN4ckmaVa9Vxs1Gyx0irfehQSP8zG1zbM3lRcrWq2ysda+R8LLIl5Lkmtn
k4By3NSR75/bfhWodjI1+lxUnQ1MyjRjl2ej1YOo04AfbUaAYS4ZW8g+z+sVXripksy2WLOWQ8vY
9GkDX4XG9IQ1GS+ihYaGnrqN5xJemnO7LuM5AlcOCi/aXAPfw6gmBgvVdyTbbV572cNMEy/C/88P
isyw2BZTjBficBfx1p298Dbg/vhYPj3wAwsQsbGoIbOKwf8gav/hs6gkLtqDvWPlX1+B4d6IvcDb
49uhwJxvCykKl0tz8YGgMvyAVRe+16smWLa3cM79zs5F9ecua34FKnNLqOFQ4GM5KTWKdNaPXVkG
pNLQDM4eWcI5ZDtffxRMQEWlg50IvYMcaDBVeI7dn3K7H7yJMZWqK8e87xQ/4YzDNAAW6zL3lxU3
9Zke2BN07NLZAS4uCiDNTABaXkUWyqjeyzSjjnz1oZDeAblbt/qB4j6iMTB0HOv+KzSSydT0TTLY
JkZqm0vdjTreDJpZKocNvR9WGRxrV1IpYgb62MlO+M1DoS0rxW5o7rji942LH3niB+ScA5sW96Nk
jXpKUe+piW1XbhIt5vfHWYhknPTxGKyqEvwLfY/AFh+3wWAITuwIEqgOF4oiiZYSnLDcQKhZ4DcX
d08RqNDSq6Xl3QMsvG+FaV3ckI7f+l3ivw7S3aOp+u5G8Caj1BRrFh8bxvxTQLYtaDaUcO+guCbg
CniUS9pS/QaGCHQlPJszSy+J1wp6CBYT8ukq7y7FJ0RzrupdBmpPkLEU6HhaKo92VsrvOku//rqe
635bQe4AF9JPi2v0KdlksDFxrwMbfMievCJ0D1NxOgo9F9HX7LvcRH66Rd6Jq/6VOoaUpmRunAAe
udzB8FVyjUyqVR1Bx7xNG+H+aB95QuIT9Vo01XLe5EmEAioppE+swbaDTcBPhk52wIDRGc2LDC5n
mLsJOhBYDKAK+TYA1bZGkDHVLHu1kpDDDxZLv+jJS2l0USFhJKilkCJuq/6hCXnsK5F/ILiRkr/o
Ax7aPkcs6HQ8f8vVoBr2xyyLI97nQdFklaSv78IorWa3/Ej1zwOE/vKTxvK5f4vTkojvxZi+utmD
15JH+xiZNBTElkYerqUoMlXvWPAKX8krVMOjZlsyX26MJE3sSAU5sJw6jJeuv7fdLMjv78ZL1Gxe
EXs3ULTU+wMmnzQPgaToEIlBaM1uxJhxzqS+l6oW9zhzLky3MCP1RkAzQDgObNdPG/RFF8G6lh4S
buEdauSR+9ucWWIGPCkWvvnOf/fdn98ZYTHSHRECCLcQkNsI9QugNPpJnePy37brmLtW4ARHLtKE
1btWLjPItB4aOn4M0R8YvI60QVpSfGyqKn2VTaDjdkjvgBsiGVgeEGOog1vrKIYBI8vkbq/iM3Pt
4t/pzfp/3dD175pB2WQmcEgDgnA/j0zfGS6ydn0nkQXVw61PV32UPDQgWzW6q5iPRamskQxu4ao0
jq1wcM6Eq2wTcDrxiN2xQ1CfrEhNcaZySrPVpa0YzEzIyxlafnD1THw4vQbtSl1RCukeclcxdDTU
l3VU80++EsOCoS6S9AtzUvNVfTdrjCMU6dh4cnZmxb1/GrodKXNjzwZTkViktbREr742SKMLT6XU
Idtvcxg08P87Mtm7c/uWqDmnc4krgxsfMdU+UH6LN/xkQ9mh6IRDGzbU4Kl8KPKZoRONscSh5RpL
AnHfZtNkcpjKMzIJN/HfT6JPlYE8JAqFIjexVpwuaLPspXpS9mk+SGq/WAljzZDc8M4ISUlK+tVe
PgqctgXY/yRuYtfni6rIhns+caZtHP6OxM79otTVOeAxNtFGJsCQgdFP/xVYjrBlevExtlpf5xid
uEQCurg/19EJKHrjxT6TDQ7Nsqv53AgMlRENzDD4KhjsctYA3B8nfR92mVilJQTi+6g1Qkh8dR+g
Ovc/YMFAAkddc9svtQdMmy7xfWvmOVvCYfYkh1bGY058xqPohVSegOK8pumj5w/6GN4saFxM7iOX
/D3BPdJHarQExuA7MzDIBjtahXugnomWUpHZqsdoasXrZDkq6EUxcZK5mKS8bqsBPDrMYksJk3yh
o1VsnFaLq7ReWiYL0h8nCI6W2B4K5sYjAq0wV5tQaolIu84hB47Zzg1svSxWvFaQxlpzluHu9e2N
RQty+RgeAJb5M/FmhO2w2IUP39n158ZWW8ja6GHuZO5pfDe5Usk1zFWSFD6rUNKPasFKRirlJQNy
8ZUbQ10exl/mxQ2vnellPwXL4Tc6EtRXDWb5PXeeY1ETbEWvD6bnW4EaIOm584W8JUkPxnl8wZF1
63VVcDRLNhWRf6PzNnYdj/7bGyu1+uQXW0/20V3+5GENpV9qLrMa4E4pTYvGNypXr/bfz4GRD25c
y/yeBncRUXvbP6xEuWhLTatz8TYsY2IdIQrdkx7O4vAuYOMkCb8jd/Lecptgu7kW9Woa5N7nfWgB
Socr/pBpeNZf9+muwt7VCsQr8M4FZYwsNPeJhiI//DxF1OpUwlsaySPaqwY8PNLM1blJK+Hr31s0
hDT8Z56G9yRCgsSOi3x7ABIIOEOpzBykj2SsF9IVColZGYXrwhH9z+P0ehyxFJ2QciLS6t9pYeMy
ntILyNXGbQa1fmluiorwm+KMbHsuiHuO/eCkTwrYadMglYfr2dijCKJXPANxAY8yDb/7UpkKBIKa
B0/EQKEEtdyXYBJG8/eQU7YJKEpseholJO9nQ5VA2amm+/Bq7CeQXSYl/aMkktMG/sDaJc+2kKgR
P1+Y/4lYWNmT7cEpPQ2HXa2Sq7HHF3+8szpKCCVaNPu95UuqNIuN8Qm1m6LlwZSAUqmcg84DyAFO
fYuf/8CMxU0UeWK8HDMKidprHZsZQ74b5yUQ3YOEr9AuEZsuLNMY8mwDeWk0OMy7h5FGcVuUTScZ
Th6n3/MTu65BLj0w5cq2gkhvabq3ExIrF/DFoZ2q+4Vy2mWQPZMgpZaXEWwS+6M7itFMPSPBsJ8p
+0PQ0MlGcBq95Vw9ROieG/B5zAJew8dXT/BSaXocNk1m3VjXP34a86utqOl07NB8IyJOYDdTDAGv
lczJz+TC/My32xZ6bAfzfQsrkcl9VxvuZoFeZA6pqrUB/PSttqRHp9wPdsd7tOusKF+vQpQOfIYL
O0+aObEXwAtH6LO5UCmu5s8ajPUHdfL3v82rnhGnHBcv+XbrmMSHPP/xsJQ6Myfw2R5887yLveh4
8sc/iJnVh5E1QjhD7n380tWNaVBuGHZ4ZcHke8Lx0zgXsvz6ldt39PikLBkeEOgecTzMNOru2WP8
8dxQTGKbmCYc/Ws47d9tlpnxoFaXyIT0E1ybx54s4UpBGVmLIw6614x9YBaf2rL3zC9auILyF14s
5ImURWDwZa2ljeEf+d4ImqieZpY5hnKO2605oL/uScAgBBh2e9sbqIJERkK8YaUaG4COlYf1GkMi
feibriZbXzi//KccD8mfBTWEwrWAiD8gyjQWXigAWs7K+3HM8CbQNuX+RURcFc7KeazlWp14flQI
v3BpkC9SGVBfydDFsWj8yDTDTOqMzXl4f4gCEJtpLsSzM4kKyAyy0i99xDzODEWA4ouUI1GU5aFd
wCZn1JUP7hXFy5YTDWIJrJhZAoxySeGqCUO3mYCZnBbeBIiBJqNdJ+YaG7gc9B047zoE5S9kk06p
mQAbZMrg034QoBswXZA3fDdSPjDXU7UW9iO9Q2RLePhixSCyuKvN//D/Wsn3LLGQyfVeMh36lDlw
1UscF1XTWYNR88H6WdyYoMCzFG9sJF6FEQPa1WJL/o4K6t8TMRwN3JLTFr8SDo1R5Xj4WAw1kxU9
qYxS0HdDDLVpHODx8EOoH0AIT/GylxRgJBEM8QS9JyF+Y2E4TgqQmW1sqaHez+ze08o1FGxlWHcu
LCqqMV25S0Kwxasg49TDeK50e/wW+/sacRrEK0YyequtPr1I4LyAlQR6ZT/4vr1njAuwGDeKZSNg
99qr91/mzRFYWWe3+a9rbYha8jqViBvduRJyPNe7wqLW8r7D417C9OJ5yyQO0cnvvojaxPv661+g
fvfdmTmjC4JaaQ0JKCHdcGsePVPeD7/G7zdHqmUvINI8pTOVQh3pMIvWYMXlOUcBfU60JFaiwkdB
ZYeV+6tPWXW67S3j/pSOfswmZG2etRFtHz3xc6XaBSQjYWefGd4/Ra6QUajSf15XAGmGgRjatGLL
CyT+8oadEzHd5PvvBWqi154pL/9qbjoeTac7bTD/cScCWrHjioWBeXtkxiGQBIChNqSttVg0Ok/F
xaud+5PnnIeI4RmTxmfOn0TMPXns1hcM1tvQdL+MdHkVhF+9jtp13hVKbSKlh6DfVqJH5TvM8WZH
ZQgEiwA/Ch3F9pLPsZuivdyTARVVcMy5ePo5vPX4RaRhbpBDss/DcDY9PqWwjzMjzuYU3glZHCP6
5QtelZr8oVXDaX56tJoOFxWrufTGKxCQ6Sc/Z7f+n5xdkb8UhcNRdZ5LW/tpsUw3DicLVuu3Y4hW
grqGX6WJvgnoRGloxWbKA6ResKt3UOpIRc5M59N2H3AU8n5Yf7CQxyv00xTb3gicutc7HbDYqT4J
vaV1RgWrJC/rcpPTDzSbwMnpD4k8ORTZnqZP5SXW9bERvgFBYsGzfyxILpufMxeZjyL7/y605wQy
g8Gb5RSZU9aVdE3HvXsni2xme7+mUfggO9MrwJ9Ha/KeaI1sJjIuxqmrxYrc81X0OVwaFLD4rUtn
mquWiCO75hNe88FpCqd7dI+4Thx6vNK4iRnEvxaxOQGxRzr6s/ugvgNdZKODEH6PUTIs3nTqrg2K
zGsj4cdqJC37MK+HL32r9i130hhfa2sqPg14fnNEyOdt1h60hx2DHz7udzxoqqNyTONmYIFZKqeK
RFp+F5mgUPlUj1lANHBZ3oYOJj/XjIVexMyipqL99wZNvGLsc5eBxmrfdVHM5DfPWHovl1TAcBEn
NKNM7emmXLS+eG2mGDc1dWKofIqM800muiruqHmaym0pb0L5qeqixjsSiakdiOjgUAXwtJ+0CoGD
dQ9DMcrMpObJxBbH2cL78UT8MebVBmwmgx90VJopEgPIF8sPF85Kc2x0e862kg0M3nJfkEW8qiUd
RbYClSvNb/7PONNzD4SyFkaWB/UhidrZjxSS64u2lz5i32IIj8MjyzgtqLiJPt4r/ZgXuG/8UutT
vYCc//eYjdM294QMQ11JXWvYRDzQQ9dihjY2bfxxNi2gkQIo+y+A1On5XFhFblXcQl68J2gR5BF0
oycHO7kDY5/cdj+EU1DVsMpWr8USoyx68h6E+AERwa5Qu3RrBHBJgmCVaVw+pVjjfejNIRI8BikG
t2hqMu51d7y6nHpCJ72wY91DZgsKbrxj3eXo+GhqufI/Mpp/FXox6wKL0zdFDnS1iUod8RKUKlB9
oZVN2whXJOml0eVKcOKTy2mA3WHhtw/5LYz7w4lEAijf3rvYo3UwyYPx5n0ZNmg/dbg+dP9F/bx0
Wb8k2/c7aq+0P90Age1PeeuvbnkqPWQafrovhOvFqC8CEQ+PDmNhtuEgC3I2kFA1tj9D7KCEEsym
/PWJZ75BHs1jAvRtsQxeIX2itNbJRx3FfnlXm8e4/2AMdSMG80qTMjXAUqwkNdcS628GERkct/hv
Na/29fPWV7VwOhVVGq0M2dihWes605NI+rTTQuTbmpDvlUJ7Shq4wOKtQcqy+BPLAtyo8/Qr3D1r
hAo8EXgwAOmeNHvVhMgX2BW3YxZmr6q0VSSo6pafzU1JoHPf4ZlkKgc11eyGofwZUDKGqV8Hsmhs
QgccRXdWe1vfxnhdMczDA/Yjw5Euc/nH46FTKdrkIUsflZIgcRGTIpB9s4IrMS9XUE0VBA9Kv62H
0TABW4pKus/GLvkSWESTO/fqVCy4aQOMftg/r0cXfoavtNje/Mvv+Tta+CyUucMgMjCBHQ0r4hr2
1kl0Dczw4I4feqyquFuV0EjcGd6inA/ZRbLI54+oAGrwgzJDNzKB97ADbzl5zKO85JXlPFCvC3PS
sV2tdUwoVn6RKOG92tti88ywrN1VQ7DS3EZMPaLQ+A+SHiRIvwpIR5dLZwnwYza8CpUMRTpLbNDI
GJCIeLVt/vkSyAhaNHNDCdp0ZOOuRJoVoDsb05UcC+NcqAI07AcEw9/xU2Y7g4BgLBX/eNJQgbe8
t3mRPNtxvnHXBjHJDzaJukPz0KF7Dc7EA13ZfsffhMFKaAeNhILLVDVkuJJYzXq2sMlvMSzJPHCG
BLyI/yFBgQ1QNut04V7sUKXAPzTiiXFWec3UABlTINxm4uliM3/+RVHinwK9T1dkLMmdA0SSgVlZ
f88Dy/hmQvk1GOnq4hgXj8swrh4gm4iimO4iZwp5esarcdbwdH8E39unrslgMkjmHEGj1htRiVkW
w/WNDEegM2GwOGQzczgBS5Cu6Uh5j44SSAuws/MTBe2yBc9b6Qp0R0DU/EnZ4d1OXTdH7vkdrJv+
Ic/CFsK2Y5IFiuFNP5XtTHv9yuJZ0GpRrT5KVzCna4Hvg1JwQJ77R6VXsct55fINqnGbrCkSt9n8
yGTWagUTEtUb8/EpdDiQEkKzvkXJafL5Jd4CP4wtBUNm7g9+6kYk3vRZ3A2ZB7wJNDNGXycQHlln
zIlZsnoB34FBjsKEm2S6Zq/hvJMJYu5LYUCahz227kNoIyYRZ9M+dAkt8DMHRGPTRlcfP9fHnor8
wa4Gn9beZm8O2YYm49W3/LRkLoOvEcXXJu79ZHsL14+4BTKvx4WpTnOpCbi+LDmV/xShx2W3NEp4
qDPmLIowVQ865JTWjIXdyo6vmaQFEoCjFKSy1XoKsh0C0gaQ04wRiclIP+m5cPpC30KcUrQuFlEk
udki4X7tmAJozlUUduBnKs2iSXI2A6NByflZyrYa6CKFIpY43drUR4Q50Apg1jxTAEqOvbMn3E2y
ikPDKwfjD4Sjmeta7Cgw6wcEB22N6ba3FQPUy25neHOQSz7hfGyQUbygLwDUwe6o4BoTN7KHpeOH
GtQcqriEpM2Zc6Z3G6rjQJBf5LeiG8YfFTBXqQKUj5ysVPdXraXS1kSw9/+BZBWKgTI/U2a3yozQ
MEBKLKzhWZeSfPEPJaDSgsiL6tp007h4yADFzINsidTopbfP4MVjnAxxtKzA/fR/alCEvaBrez4H
s6w2lmJu/52iyKFAzMSbb9+fyhfmrCICYVlyDQoyWs4W/qZqJBnjYOC/gHVOpsuREVQ+OMT4isIr
Z/BPv35N45zJ7Vk8yj8Usxw75Yb2fqIemVCeCjoLrxtDGRdQTRB3RjNuEei0lGk1tSEneJ9tZoP2
n/pxYrLY3udkiTjZmBXTBd6uYIQRzSX7Zr0Zo4q0l0iuwoVVeLT+sC/IqoOIFoGSOga9Ai6mL2Hv
aXqF0N9zbF6EKKaDzjPlConnmE/4dj/vO8gtfavVKpQ4SPRt5kRV2Ko5ibjSDevdym8L0mjYNHHT
bLlL873Y72AlmKY3OxvZT99R/fmzHZlZ2nFWf2OFnlZWuuM+2Iq9X8IsqER+offryeQ/Yv+Glt6t
OgrwLA77+miKXR8CS3609KT6qbVu9IhDxA/8e2EeIJkY0OlVHS2OmlI8slYWSeMpFz8KYSPsj4Gl
yg0eZ0SUPBMxn/1Fyi+mGH4LcI+5MTYIknF05AvafqSpL1zthbguhvc7juLiumh7ZRJrDag0vvKw
5XAFmuPOs2erVfUh2JqBp1OfCimGJW87+y2FUAzNUDl0Whu6nKVl/niAxBuLMeufykcqM6vEB/jU
pa+2xCzD1wQzT8socHDl/7uEKtsE4eoOzaFcY+QhRWlhrw/7+ylJXVaaO3XTjAxrhGN3Ljo1zYew
+h8MqBh3e1haeC3qE/c83UxsiESi1m22E+PlcvsX90ydL9MVwiBJQVhqJZBzmDw/4ArdfGMAK8OG
zHmWeV+r8Ndr59FDoTIV2H4QGAmLlTqvmtEai0OuHwIrz5ncAgr+6KT/j//wa4Lu0XVdrh4Muy7/
xSffnk4Gdt5OTkpLCADYgEJDpHfbTS6kWnuvCgWLYYyVS30oeKe5ZsXrvWwq3aHvKeWwCqCQ1wFZ
ENgGNUQecgXau9uR7qqVItU2RsBVAN1+kEyjNyI019Diay02Rq73VrpF/h1Gdce+ES+SXh/OnrQW
efeeZgzGMegSyPFCu/RalIblLu97gF3WyT8iulPosV9mEavA3iCop6Nl9141ksyH2WmC4LvYPrw4
3ayF14R8LTGkCvMtTZ8gflsBGU+q7Tx895iES9je3yetJ4jckJB2Vlnr9/wnwua7vqMVObjZKNe/
55IRlsK9zkNsn/WdAV8orxF8+3hqtlnO7r8SbwquEnFArnHQMwkJovmj/CClXEC4dT0FeleqLgLC
S4OoMY1I9bJsYRJJ3yzRHUR10fRqsfDeRaxbf7FUXmbWbncYdJQDmvhTSijyqT8bUzsmGe/+2Yg4
UX4WEPAHzuKcIwtiF8jBBXnwv/JloGIYzrbYObJ669hyU0JZSq3QyRUjmqBaxD2KO8+H3HY6yb+6
VdSWG/DbN5wkkGZJkVhfgyK3NnJGOpj/mbevGcqzNuw25OhyarxmK84Z9nMzKFs52nyYjXIUCqlo
Mpm5dC8kNZ0db87yAywURHy5aToUnqKHeqCXZtYH9YW7L2RziEYmFv4IapbrEejBbLvVqS688BCO
LAWhJz+z0XJUhdfmv2UY24n7cm8rWGQ8JJkP/8bQ+4rL2G2g4a7vi2w5SRE13h3+FizB0focZOyU
GItsQRtUb9SwebGr8IydxbFthX6NLJPuYV6BCaqS/6UzZ/LgJVRAuU2zZsgdQVGJ/19+GnVWNT5H
UWZMd13i7TUJkxKsYY48G1k8csq9btmqoXr4VqsSAoKbiHTdSputuAwj4cT9KcZpv1fq3/4Ym4/q
FVVZMN9OiaCWg50AoWAjWuSCnXgDMXLyK0jADVOyNwrODE0FXjapvAQRpCeXzNVI7mCFvYPtOWc/
WRaWILRH6laWTL8u1UwIzpeZKIlG5mHIAisJecQsx0o59h++/K5MPPjEjsjOu8C75RAIdjrWzWEu
/tDZOqpXk1YiFzZyWt/wODuVDr/crqmYzyG8SNyUexV+PFmgjU/uf4TwNDUxuit8+Tem42enoK8r
Hg+XkKxFKm0G16bhZ/efYzfMAg/JyoKY+B6mLQyDYE567LjLYXt8a20sWpXpVVOQFbZhtt6Sb06/
UhtbVoEh9z9cCUtYQ1JGlirnCmRVy4QqWUyD+LiY5rnWWW+8J5S0IhnmhaxVS9C5WUy3BqTboDIS
fXsC6qZmMsXjWaui6VZqQaR1rNm5ZOLzQzpBMh/5aZuFhDy5/3+4tUKwmVzn0TnS0aOItgzaEi8w
y/Cn6PWJ1GUcinvVZ6FA8XGpt5UJnjwQgkC/Fg9eEIiY2bnrsgv+6jOtN1HHzeLU2ja5l7LkDAmP
M1nKWjMSPwDlSJJI5MJQ1hv3/8j+lAP8m3G16lnCemHYnGdTxp/U72fxsoJh5bPWtBxkQP3SDkeH
gjsdEjyTk0arfc8HnlqawGIRRE29fWvhvUiXN7FdqSL7QaVjvFMwSe7XvXFjChkVZCfwBMxdYe4e
/M3LOF1HurhixiX8mqVPo3eaKJURlgjxD1IDyoV+8TWxvyJFUXob3oKthwXABV11vL9JT2NucDqC
RsZKoxYcEvT+5grFFLS/TDJwkcR5EhDGlGfWZWWXq8zBliZNfnAS3oKtYzXZlIamcHEKjEZz2Tyw
MrMrmoncYUdR3zQqt36nX3koUPRdZksUV6tzVRRmP+gmswiWpLgdQ6TUlaFivVBOI6ynILeFpgJk
ConCz6mMLH8bI+dKV8MuEqiGj3On8Y5d2dqHZJcbYt7CYnsiPNIpyZZ3itGB2VxXyelsf23QfCZF
jxGYdl/HFMIYQ3YIPPWjwH3yQjazjePmGwvQm+bj3O0CrgtGF+isk6NQFmtiD5GgzQ6WvWGFEUqC
YeD/m5PBLG0BXttO0xx3C3wFHQ5d30dRxBzioudnqO3fh/ozXGhbfr4Tehu90mAD3li5d6WsFdgq
ujL4cEaSzeZ8WrW9uSajFbzZoCYW7MG5IAwCwhnwHZtk6sVR1vocmswJQtuxKpXO3go3QnSwyQRu
sGOpq3lFp38n3YzOzLBChXju8Uac0ivJmqxWPXEQYa4smi0OBNmrhvjLueMg4/SnSItdqNDapDuK
9HmnYbs8Gxu56Ovd7RomB56NuOSreUADio6DkORP6zQDWQ71yKeswaRulfxSW7FbMvwLS4vevN4o
DHX0lC+7zqg6AOzfXYt90vPqYcs92pXWduVakOmU6yoRawjTGHGho5mil6/SesPlAeVip5vvNYFV
bqo/hWEDx8FvjAj96DhzhKQKa0UKKmI3N+R5qK+++y9TmCJJPQYidlm5sL0ljU9nyZbfV1nic4Jy
vwWnSkz7ngFMGQjkNSk5ASIFOke5uCcylZCWepPMlz85n/ae+cihQz3bvgjprjyAaU2ZBqHMN5hg
lJzVyUbM2IutUWjuaxDdGhg6/Etf4zwWuOyesXvhKehFEMAV91oiMohJObDtlEiDTJcWedXpp9jk
KCGuQwvGkvap8BUcdu8OtducyDo/aHGoQPbiZ/gandXL8jLYT3EZAMTOMhRbWoLdCZo2Oe+ytaPH
MemQ/SokyUzxGfvTNq2msgkr+PgaGRb/1HDxUEIxdDyL/hF1sGtUoI5j4bn5oMBT62zxLDiN/iqf
2n+t1xUSiQ3i3Hg6aeetza23e/4X+FekTL8h4x//sfYibBwQymk3uu7aOrmJH7KNQVVoVkbHvRTr
BcEVSuu9DeN9wteR9runM9msYE1StINRHSo5vyNd+5Uqz1/LnHMGzat16+H8gHGVRC8JT6mADsdH
rPzNdrYJM//VI0ToQJC9VFQBF22PI2FPkADGril0t22P3XeRpni+mmnGAUIs6eMypjSZMPe3NCQO
Wkv5kmzIqPg4FAEzzwbMrqsCjhvR10Vx6zUd3jQK5MM/KltzaXDUQo9kpCCKZ66upA8HGhJRzseZ
8lASxV2AImB3mEzxwJf5vUj0tcDr6qZOxf4lJ6+NIEiBqj9ckaiCsimsrr2DuWVkR39eOkPfoAdQ
xNKy1qgVT+ftxh9ElSck6/0Tm40Gh7VIinUndKN1Vugkrd6MHyqMRq0pwcuFXVAB4gAmqZ0O4iK3
BFpKLac0TvpI3n7EF4RlWAIMrrFAXv0+FIOF9Pgni8AINwb0Gb7BFq1rN1L4RXvWTr7NOFBq7nDY
SUnz7tQp4IaSROAkHE3hAva4mCyaNBOi26kwN5bZoxdaAbl4XeWZUl+Jyq3gq2rd1VQMAvSUA+5y
+C4y4MNGQ40T6JDjC23UdNYmjnpykU4heRl2nzb0+aYxUbSaweMa28DLmwIz45A1/j7L9WE7cvjG
VzGCYoOdfjnoQu0kwhcyrdf0m8dWl6ebk4F29cJkrjTc7InPawcLEDHbQOpyYmI0tu9hiFO5t38p
DatMU+sDe/w9jKesbUBUipEGWJAZmlOPVRKcGdgOidC3hZ4g0swPMfVmUngxtkDAvJuSWNs93hkT
5fOS3TRLzDQui9aXDtRbUcc8c80jcLOb6Z3gfjXiPuQY3FQ/C4SjVWDCqs5yO5ZuIriDZWeM8Mrw
4cczTtlQ9epJF53Qvt4lOz75o4wdNErt03oOo+9BqbsgKe0XyoBGPfoFAYgAHVy2pHCQIjpEQH+q
ipsdURolvjNVKdxG7rawFTfVFYCsj7BKxEMPgp85rgYE5yub+2Rw4M1fjIBag+HSxF1BR9vGUidV
LEq8W5S9QEd0mQK1dfFF393F/0WnZO/hNE7ngUswko5/PTe95UJ8mQTdOJ5fnfvz0qhRKu1nLp7x
5b7Qreva//idGgWpuHVMsfegXWp5mdmHSVMwwPhLOg/CqGCafibhGf7u4CNeF8wUNYu1mTzqGX52
9mPte/wiSmgIg0dz4hBU4c+jz88Bq2uwbS/Zyb2Z/VNAdL37F9yQOdsqNmzTR0J1hpjiDCgb808E
2NWY6GRaNXYjz90OrYn7nOszbu8pN0GOFOkNdJA+gYJn7ApXbV54ARDP04nflhj8TIAhFLsqJaya
WBhNH5kRb+i853KqIEbkhzydOaaWjdBqNaR05cqyMqZxGdjFeWxqFFdZkvW62ICc0FzC97OJOkWQ
KVQFVKCk2Vf4JT0FWkJ5ePEATyJCX7UiNpaj3/pPliNbKOgXdn1VVAu/IcdEFxvDFieRdhQ3+lWR
kO6L7vKfi7DRpXfYeP7AwmW6avNpUsCumfgRCI63aR21oCIZIXNkeK//2EJ5PwE8oB8WgkxzHu3a
vXwmcVdr/8cwaOEtL7fBWcPzJ/UBTgVWAjm6y4FX7gncNlG/bqjY3i/+V177lbImYqDei+UB6Rlf
gxEQd6plx/289vu2fMrz7kDl4Kwr4iAlFXnnr2+j9GAusRCy8/+NK6NPdb8vzDgQAYhAgxHzPKJf
UMfchPxeEJhhx+xCHF67HS11h8Fa+aR69zLA34g99DIu8f1ebAZH191P3yu9oCevn4uadDlPr+kS
FD8A0TmQwNBRBX3gYOgb4NGbKe/L8GZer1Heo3h72l1eczh6v3L2Bh5cz2tpXqGVOePBJTYnldTj
1xb3A+zWffTGcGuV5Fu5eFd2UvsIAfUNRzTVxCusgq+VuVJ3z/fGNMXDoD6A3d1YaDcy7l3LsVr6
dePNKeKrEvAHsy3C3g+3hfrwaoD2tsGlud+umX4xWeGOqd4FndMsuZfxJE9gscXOlLfKh10DxYGb
OknasfJC6Mit8sG7zkJ7fuHeLm7YGAVUnAVkZMz0QP4OUluUKaT2hg5QRhL0kF9Jbge8XO6thP8T
33y6RtjdJgD9p5fIWaPp/5stz6R2DG/6oXAbx81jmIerIxqW3YmBNqFJTKcwNIfq8t0gU2SwQFpq
C3j7vebw9yU+IENGPpZI2JHahJw6JEURYBI0EFChcRcR8f4TsRiycCxqxj8F98T1AHwh/swWJv9T
DeE91pADH4e0/nOe+tq8bRRxFF0kVkCPhUSAg5jthpSyrOEQC+JNvJwb5xCp24W6FBMdmuIVJvSU
D8F/hK+94awsdgLsFC7yX3XN3a7WvV5BdX4ni1xXeoy6prpHpSm9oEMgZPpz3xucrLiTRUjI24BA
fnpQnIKEXHmzaSAgJOlGpqqT4gpHXPSbnJ34H4HErFZYElWyR/H+XzMS2WXbno7MowEUM2iON4FP
Adq8zQYaooj/qOmyDNmUNMb6OBtgdEUgxEt5F2N9CTjnPZ8SnwKA3Jqg8zScVnPbO2wkTh2YBZU/
A2fdVWtAjt6Stel6WZTAr/+Jk4mT60HawRQ+3aJA+pD9LObrfdAGiaHGhWGc3nqEGNlKEgGLJZre
s4HnZuqfj058tsjRlSaPgGpEGpnHLrnpm8qWLLQCJvz9hEhoRqUpGPvtAyyTo+ogaFrasFFE9EQ7
PX2Q3j8x5rIb6Bt0PlZaa3cawzkgrZjwRO+0KeNIano2fCqeBeON7N3y5JtJlJ3qdajk9e+AEJPx
4L+XRV54WXxXL0AWHFVybn2bCWpk/9GPy9QggjO5LDoSwny4Rc3JhZt11itTZ8UXeJuSmf2Ic51n
2mXQmSY8nWpdxJHKq9BnV/jx0F13AYDmCNnHOqNCDK981Gm7OvoiwtEUMqM+biMUSbmwFjjCa+Dh
1W2UrJjUbkWUAeijCzVbTZAE6S8/PitKNVkN3lyGUcC4OgyHqUS4lvjhe5qgsz3AsWhMSP6J4uef
FQLKgbvPCaGqOtcqwsEXGOPHjz5VOEEifBxNrGN27rD1MvXTVKxrnenru7IEwCq5If02IrXJ1j29
IAd8pkfRAWC7WpCLwkHPUo62t+to0mFgu32oIIGT1LKOWDipOOIT7FlHDBz0Xa0cPKCtTkQhTNAE
0MS7h9/oRP+p+TLm7I/Y9pUcJwyQkLybCHIYjLT4M23fXxS3QQgsv5GMq8RvYmG6umVen18fIe7Q
D+DbP3BR6R5KHLQhLhboZG7EP3eDPqDxwujsu7Wnpwv2IhUwRA+3z8JtChvgk1ABwNwUdvel79Mg
QdgRirzNcjK4+tHIoxuJe8HLyl1nawHM597qyxz/Pd+gGbeziry0cObPjM7YxvgvP56kNr4QRoKG
rzLH883zb9BU+W5g072HXOjAzoTYZMHiBlWoVj0vMufz6fK6oZ4cEE3PzVI6wGeTSrz5tY4LN38E
OHhVIqiIiAUMqoBzXGsKsC0PnhC52Fo/ZbiJduOwSChHMuowKd2GH6IyUNC8EQ6fM0/WXC4BUWLH
9bPx/zgr8HEu5X7dhremcqcbPM7XpCqjXM0vwIWYdseW7Cx1e2tMd9ePSBVtO7mK0GIYHHj2PsDt
2L5mwIrGs2ixmvB450dUpyNdje5/Nv6qcU+k77mztjUm3tNTBa8ZHrgS6tzQDTswk3gi42sc/88Y
NKicCVdzZz/lQFZ68uqRsLolrkQ2pDV5WhIH0Hmzjj0d/P0smjUs7P23EkVQgUfO33a+kLKHQvU+
TI0guSyV8gMMmeOTmp19nGksrcJaTF/mwT7h3CqDVgvsdvyiTSHWZnAW9bIP6JtnRvzyzbjdA6yK
ziGHuGKOxDRU6fd0yRXSff1/gZ9owxxWJ9wEoYJ7gfPaWoQtotmyBjzZXqTgthSVmH0mBuMxsQZO
M5q1r9DOMyNYVQrME9lqGeMDEk+1IH1ukxzLHJgTOrV4kirFqjr75fP9c/ppJglk74C4JTAQBO44
eGUhVcgd72LeEIPiQzDUZScRVpnwGnbam2CwTqsiLlczGxPleps8wBTwgZ+JNoYxJgfffRFgJNM1
IVNWBbYgDiDH5hZgY44QdJ/ZdVnMtVAFJ8b050XATzjkuBLUcSZF6tMr2xk5Ifi09o64J4l66i3b
Atb52CmUeIaA3c9x2hCUCQeABgk/xXnJGu/fBRMm2Tpt5lIGmjM2fGIZtjJWw0AwJMiUEswRC2DO
gEXm9yTS5jcLWGbS71wk7qvBVaevTPTO9KYe+qlLeMJt7XoHiVTscMuZ3FVref34RDHWM1QVOLKr
aFcJzG3qgWOW3/jhSqqmi1bmiaBtkpxnACZUPpQz6uncvGgYVOGJ/0akHuUWGs/7Ivi5qfJoZ+/q
C5D5Vhv8CK8ChxvmMxI5LTHa4n1DazVfQYVjCLpPYtZSCBb5Yn9cvtqGWouUIWpvc0CAwgMPhXqc
oKOSp95A8EPc9zrgTm5El4VLhBQvcsMbLS4O/jEt/b0v2rw/aAYJ3/e3HthZPFkPSWUQu7RR+iqZ
N/AFEATl8E8EJTfovuHpX238edW1Vew+OfoF50PcIRzVwCGiLYD4hFIQab5YXFZciQhzsPEcc0GM
50A8X2pwdzyhAGV1oQdqX4RNFh23uvgTBxoWRDWoIv9d1/uBCbUwAktGUFsX1UclE00j7FPalF8u
Ujrl5rISz3PW4aeq334Bz3cwy3kb7pPm+RufeRe7FDTER7D509rH9xwXvZM67HCDlmi+vWzH/beu
W93Jgjm8Ol2eXD7cWCsImLjxNy6iyCiZ/Z+PnNyGhufag28OUewPtsY2BjLGj0i4GdD95YwJGvd4
cEiLN30L/Y+xAdeWPdNHLxsfO83AHwlLwwvetos/5HxKqMqoL7bZTTJ4ROVsXdacnV3YGrSgo6Kn
N7x4ShM0cDCdpUZK+ayhIvdClIi9x5GK10gUv/IDDF1o3ukkcx7MZA/22XChB2mjHkwRLj5djpYR
KGRWrFeAdMj2uxg6m86sDWtt/PuWX6ciTNAXfM3afiOVQ792f5vVxKhqtu95AtWeCrfRh2+M/Ry6
c3n76DkJ7rMo5MbGc63/4HTb4KHYr7KHpYfgwe3T5ZAGt12y2S+bRYeLrjKmi+gkx0tkjptYYIQX
azkyMMrCbDedgPn0wG1xHyKM++ccsXu6DFiq/cZwH8u1BUetX749P0dfFIUDb++XHTuOfuNJzmCT
nHy8JQMgz5wj2iMdZPuKhYv0r00cjxYEOyJSM+LcjqUUqOqUE8rfnSmOB/WmD8ZW3Fy6rKut3/UB
ZXGzaqT1jO23lRYMxhbDt4B4/tnOGz1vu+c8TdiJKc1HuAr9vHXZPqIBV0ahT73qvik5kdTS0vUI
b6Ff+DJtEUOQ/V5ttJl4LcXlP4AjHRMSdoN25wGFPdfiHItgumOkd8zrEjAlfHkyaEJEqqlNBKhk
XprguqEYGZr/t/XgkW5KY8KlD0NrhLRW04yYc8XPdlpUqxTboUTrLnIJbiDHRIVmBXutwyryYoft
fqjLKwAybXErCwbWf9T+jsFtWfj+5hhsJS9CRGR9z51l2Daezwl+gyY6++hceqquZcVkBZzmNLmV
Wcw3MQf1+uqSYyRkO7SoRey7Fh+pdbR2R9eQxlzYa063pMQCXBi7a/D1vDAn5SqXI0Y83QvGXUo3
tsFYCEETT461ZxgqKYufLgZuTobaBRq87o7wJ7QLtt3biEvVuZoz9I6y+0+wt0gQ4YvTV9zhBixI
jIHAR8WDV8pFJyXyUhijL7djqv1wYRB4koIdJAU+MntHAvbWss0d1mrvHnFM2MJMWZZHrkZmdPUd
q+upPo5e8OSJVcjCM5/aKF2EZrHBM+6PoXJ3r0sxcR7RgHxiv9BHs6PAOOhubZuOg/d61hjQyOmU
BuwlvNebZ45GnASZjYWs3tyKnuHRYnc9xpqZl8p6ykDROu7crzYciz6bCYdT7CGdVN5KS76U7ITI
TEhDy419K3h0ZXKbY2FF68m5oJ3Rhuv/d4/k08ho2rwTTTQvADaYjHHAlGWI/cdEVIoTMZkUhNoJ
MhIER5/nD23Fv8W9zaJ7jiPn95qLsfx6lco9sq72LUoLSoSdxJX3ADeMZGfqjSwsXqIO5NpIpGv9
8PSYL+8XKJL9F9HzIGS3pdWBMjinA5/UNqfzyNtwKCbIOCt55cdNQoR5oEqlhufK9Ii26jXaqGoT
mfoPnzvP9X0kwYWpmzLoNmSY0i9Gb+obUByngJ+DtD6nvwRed7cG7MEU6oYnU1mplMIQUFoAYuq9
TgUa8dzqrWlUCsMDnuWPBJVUMlCQleZ9PmyxbxUdcDmoMFZhHxRNg9mGcL+ov+uJOn+Fv5GE5vuv
zuwQXaoLzP0r72C2o/cuLPp073Jz8capCKzUeLlI5ELsSxP87cWgvJ3cm/v+zMent97Pi/3dEINy
ZDoKucGjEkzJ3ATpRFZwJMdDXh+mfO7tS34ryUNY3F5tHUInsFX+yDaBBmy64dDjTj2S33WBkD4X
/iYW7urSqNSo9Zndu8rVDE5D8cNTOLW9WpcaIBndeu58kownWK4JhZ4LV3Tx2PXF31aHRlsVjo1K
SlypYS0bhKjXuGeqrdTKQFycPeGPyRkJWRvNnuFntlNo0Mwwq/8HC/C7Sy8CxHqQUOQ/XtS9uNsX
ASBMIOh4BU6SeZRyJ9dzWSWUtjDlP89oJBc5WWwD1dionkKp1sF8zH0kBS6tEX4JnUPEAzVeT1wQ
CIqWczGqAYbkgrN/nWy+c/4WYo37UdKUQwoZCE4+ixLGuglTEDhhcxFfgaNj0ug7ry9dgg78nrRv
FbKE3WSk4uIeRFGOJAP9ordZZiRq6dGhwovM5CsxZALP4zcG6R2cYg1ACERrwK5azzkA7CwGUthD
cBOl2tiSphOGFR+M2W27RAdOqZ/nJIVQtbIKwpzmcadjwCdH/tUIU2fBP6Wli4KozZSQ+imNGNN+
qNGQGdJAL3+Fl2NqzqMwrACdFnv6zm2hkew786WxVreyWuC82CWVLwozztS2j+zTHqmRbICz+YiH
tF9ltOXTv1RODkaJ+e6w7Z36MHKrT4bxLPoCb5EGQ7s7Y5thkfBvU9QkIBAlmoSlxOYywL81siCB
XtbkqpTNxQyRNkRZBxKraAk9bccPwfW5FZh2LAhaFr+zRO09VzjfSSjjDsA8FFdMiy8h9Or6P8dy
dXMfFaSes1vf5XmYvnv9nnT7o+Rm9WJTomyGwTiUwItCV1/XolRFMh6EgqNsbRlXaxox8M4Q6Xnw
26FrGuct+lILEsPXsZnO8DmXup7Q9jSfi4wSK0L4YkOS1YvS/K7CkNrQKBYpBHtAZwLs8R3BMyxp
JEDckWbpl/sH+RpjPJtPlF8RonHF4yHUmU/yJPW2GEpYE2jdyv4DSDloO+awYw58te1k8qsuS7Py
Z5jm8bLJtb2OPLl0WcQ2EWZqt+Lg/uVuViw1nK7A6tU8Qo2wd4HuD/DFwpv4gnEi6JbB5cqQRrNS
vgHaD6ZfncymdH3qfuy3gSgnJk0es/Q2qTLXEk5+vdN6MVV+zytdgt4VdZCkHh8y4q34wAlHopRm
XVQ5ByB+o93NXBDs/Oe2AXjDPlX3x814zE+EHNPBLy6RyDfSr1gNtzXXfhageIa9IdTVU859M5ib
4z5M7HzS2iYjohC0FyAfaKimqjyT9fTT/qQJDlKVDVFnJE5ki2h422qvDxz8SSQ5f/jB9cbUqIRP
gH8aengTuMUWXPQdpQW7bIJjETsqGagUV1ss7E702LZX4koMc208g6/z7fPcCtdvuEwhKMJbkz7u
mka/WI8lq632jrTvJorZHHfFkWU53MUAzAjylcpphp8w4oZsN62UYrifWgKSerQUdc6szbmsGi0O
t/PcdT1lp4s2UuwKSb/hmIolpumNgxYP/LcjN75JMewmxYUrUg36vH16MmlAcfBZpuaDBAkWeszP
Agr9hmvTZ/yCdTkhXTgmJhf5IiGyNToyHgVUw1YsE4AySgOVGnKuQJpn2aiA3gL+BQit9kREhUrt
I6MtwCfrQseiQVERxE8sNXL6K426MKgZ1F9E6SkSKpE1PB+99D0g0qFsdMcmhfdq/2xm2/GRz3as
vmIavBe3RB8BtOwJxd2h1ylOQfiFQwfpBZAFsQQbKOUAGPi27RNeG/SmM/r7ZdVBBOG/xLqB0Ovl
im438J6E03mUWMLII3n4evm1jt+W7Fn388fzVF5pbniHYJwRkTdVI9MHg7OADc1C7aKqfl8Jh/eE
oBZ005atVuSJts+RyfDVQ9afi35DJqJPruKWVI2Gx+6Qiq7VzxZx1EjwFCylQadLHO0cqbPxyb0d
YjiqqsLfC5RVElWfU+26oe0oC0fLZfmoP+FAyK97h4Y3wmjIvokHyHs/s2xuBiR8sHk83irMz2/O
gnpLc6QxPxUwUKCgFgg5Pr2u6iGntq5QoT+xX4jJlay3L1uvcO0aAsoM3cd/FSMhREHWJglkHBZg
Xo70ZwNw3lNHWGOytsX5WgfHtfR0Xh1eKLGm5i54/wKJSLcrvvjVpQ0gjQeJldDxCDZoWIx3A9qh
B8NFCx5ov8n1n13YvzREGdCN0+nYLxd0rA0CmIio8SLX+e5et3IdaMtnnW4g5Dg6RXZMM/k8hDg0
3LSZP4jaJTkV5Quwvj6O8+y9+UI8UuFbnsqDInAompvHpTGtw+rDz16WoDiKga592u8Xei9CS6AM
6MMPrsn8F5kFA44VBU9exEN1peJgFp3YeFd1MQW6+WHQ+F41sLk5gKLjT/jspNnhX8vHprxSTUjC
jXysdXpVLdzd0xns3Vk3imDUxj59YVx6+UWWR9zL/bRk70vIF2Dt55DOQptB5dw+HyYaMgFZ4M01
84gKPS5cW1Q7sNG9I3Cllznlq8kq9z3VvxelrqFu5Y99SVjLVTX5KsMM7i5YQ2O3wOrlN712P4az
yGUHDkYxhv9MRj4LOk01oq8EoXauTKXY7tWXpJ8CBk3nb4fa/cMuhEw9JHQIbZCObfOR7r4VyOvR
sjT6vw6SCxFKvDpjLTEsAFOp5sSvN+B4oMTZO0pVW5fZFGu96hsOzynXkNVoWRWG5CbRyJiEMD9w
GgHGSrUn0ybCtjgOouIbMSLBedm7DzlpsH8Rr7wHioRmKXvUlQQnshXVWJRRSVqoCe6sa71tepL6
jLN+prqLtvaRv7wnX8LVmkLx8shr5VlEDxVjd3PBBgxDAgbH3Ki+MxMBJGDnDxplGH0WSNdHQV5U
YmyUrtzHLgSEe2DoZfXvhE+ZENXNuM+fbWlSC7PZsVEFcRGIwGDa/7ES/LJ1SiH+UqEH+ABIpOcx
9fq0uwS5bbmu5CrOKvfXHhFO8OkFOQy8Lf5G62+iz257w/Y/Vuo3pQAOvVdU85zd6LzmmPu+Pc+I
dAKMxr0KmElyV1K8h2ntuebk7fsyhlu6auaqYvSTrrbR+8k2mCuYv95veYSZE0h7NwFzZmmojzOk
YbWMUhmluTMuA3JA+l5r3GOy1byKmmdl/XwkZjaNTysMCya7bPCRxZFc3w1CXvyQTp/4ybqXZyVM
p6Auzo3/09IDeygvyRubYosATLtzWarGN79JoHuhlsVQ69tuh+0JYR6hrgaHexVrZAABK6uZMCzy
AqzstYhksiDI7v1vn2HL5jZGWIuvAvo7fTGKHy5NGDDZsiBDInHsnwsh4ksRTMcTZuNcJwUx0XVK
XRq/m1SlgcyfEIBa4r5E/hBX7TxA6x28tkY34jel9UiOZBRdwGIkN2LfS9zvQih5eiHf1rmBHZSc
8md7y2PCV1xcJlhj9rMgke5UFfN3wEv4oYQgiMxNiClWtX0VBHZ6TK2OtJGGX2k9lr8ATdJtfSsL
bLvLgDu2aMVA9AfqvEXn3S6hHyxDcG133HpuvBERM03wEd6tw6pZPNiLmYAC82RWUudul2KsGWMg
xaqYmfio5R0e6a0RqZuFNATkWCb3pBB97cIaZXTr/8xykh30epzy4dmtv9QRVyQMg0UrhCjRmo/2
T0sqVyfH5StQ8sBR5OfME3+e4/DPStw9P40uM6lVCyNoWZdmnE0sOhORe0KCbOEOB8B2BL5QSde1
M3WrmU7EKYBwslhNVxx8xy40JMymTpH8gf7zxjdwHLQ5g+0JhwkeQv0MjRKf/5DA/ZMNfpAOe3+p
RLpgszz6mHY9jY8Hhvqzfwc3+fTgcKJQ99nYaEVpnHhlM56s7R4J3ii6yy3aKrqU/t4Q4olr/XY8
DQoOA3SgQWCKWKvsniFXiWIPr1VEHF/i2/9gosP/E8/BzSBoFonml++EhVkdBIygyjlAyE75iRTc
U9wgHO144ppVgJwxiipFFiSQ3XIgze3U5kF5/T+VoFa9B6QnYL2mtbCMTG9pi8v98Uc1yS5pencA
GJfICAu6x8YwnpuWL320ffEISXFh92ikGRczrlbSlaBoro94tg/FJhSR0OOgPATr0UW3ED+Si34/
M9RkWC8fEtUgiI1VkjGRpOayCgkeaKG19wc3afvOYOv4qBJG6Vd70mEeV0+EFRiCu2W2B75DmkyN
eIO/DvIXNZVy/+D+RqAq2QpQJIgkzA7GEAd237jCvgSJt4hzKhcFypwx7QkIPwNFDuAjfvLFiDur
mPz1Kfv69AO5TbbDb1VvWaz3AIM5TlAxv+u6sWnT7d2/JoDG8D0RvPYdmgl+Hmej6Gz70bZuGAsY
xLRQA8VqBIkzrw3X9LsOkTJPUOzs6Mh1es9ZoHtJg52x329hQ/bMuq5gu7smcDrkAAv61pSSajG8
W1yLstc7qEpaTItmchffmadu6Jvg9enm/c18GBPxriz6YXTYACoYSgyh3lPnzRHwkg8w49fe6gj5
UZZ670nOXqbvXAE51fELE8nebkFAy+ST5xfBOVJIlEBSRCoSTNBuvkHN9FPyRUBTdFiTQKUAyf7F
ob9WFEbE5SqXyUZpr8ubWDYpskoU14eSTS+IoBr4daGiP05vS+X1Yw5ppWgeM0GMiob2rZBs4RAP
ZP/4qLd46AIWt2jGmPQ0eHEIvDzN6RLGvEE2aA0H1d8RU6NdbLVmSl5URAw8v5uB4q0gH0RspTBh
JQSvbMy3xGKfsBHgJP6IEfJ8IMyRxmurrx7r5KvDkp8naFc2FyUccy1zEuqpqj6Yp86yDZdVqmQm
2DD+Mgo0TrDxa4yulH7i51ZyRTkEFd0ZrfOnbIqi1tAIRreJAtExArWPcJOpUzr/OkUkUdzVA0Yp
Yos/ngT0DxqXE5LY9WU/fyWZzDdN05c6MRlBKDwwP6RfTRdA7xmMu49WRUzWpT3XjlU1+6HHxv9P
h//RwMXB6lUDP5ActM8adU4HqLbCYeFPebk1bpcshMbZQGTBNnzFKo1FqMyyxAdwCazmkNeLDfLz
4hgBJh7uztdjqyCQaXI5qAp5SuAkPEOKjDnMQ8YJQoF+1KsNJ1cytTE+Ofho1gXguiKDtlPsThlG
KJNFSPLKrYNuCMHuGwcsON1WaQKR0GT7W0TROqM7wJ1NXMW5L2fre8AEGJ272Nz/m8yM721qix25
NT8dlhazAAegMZcU1Y5f4OQScYumrMsFfULXn6Rc4w7FBgOQbl6ZVjzVtrrm5wS93uB/XJtNZax/
7w4NM4VtiIoU9lbVp6wJOeg37OzU/oWarfu/ImQye65lvv8ZvCFuVYnHqdMPYKRQNYBNoyLRRXJF
ahRb9h/IMbo6vd1rCr0RYL2TKKZjj/WSNYwVgZxco6we/+puCQNZtU4U7ZwUEcX4vGdGSxQ0YNmd
0DQ0pbDM8koxtq7ktg+9REYRzonMfHmoxSXv62kiYGph8PM1JjNaCvne5EMZLRzLCuBf+YaPdACu
sD+2HBTjwfB4wHE3DB9mbsoIOZDL5shGCahm2ZrphXG+O356+3pOmTRATmm39o3Bfh69JHIN0fQu
arRyMHYtXqjvJsoH45Xv8ulxl8Xgh8ZQXgfS4SWhB+T+cVduoFXRJxSfebLOzDli6C3WKza0/a8I
wip9ppqvqq3IergNKf4B1t7L0L3Vl3G8LxTgMveUnFyzYumchVnJ8XL5njCYYF19nDPy4SYqYsCH
ntLd61nCmIkodoY7ka+97tRMhYqWvcM1Cw7QJObg4o72n90SdzMQdmKR72urkukxKeKMIYRlZHdz
FgwZgkshjKaJtymU4CY50KoiG30XenLKtjVuKKu4CXhoQ9qF0M10mevQKZ0cTskpobIwPfxxx1K3
wffEFBJG+MJ3in3cMErGZ3ZTNQXwdoJNay9FIITXXkQLroHSz0ryivoLKwdXfdiSi5PfSOLeFLss
omxPx6Xh7LUnmxr9da0kptmvhth3EC3KT44FOfibqC1v3N38KrgCZfGKUTJ+mjJbQK6yPSNHaYT/
ODTWWaO7wKHryCnWUjTQPdsNCDSW9s3HkoplV16DKNWzPoj4mjyWjhy2L17JC9CA0sMoXm731u3S
gzWkZQGawpT3m/FzMlKxnef3/iGPy0tnn+ocnfPQDGT+6lBFFg1d8HFHmIvMW/zeq4Bb90YaYdaW
wHcBWIPLC8LG9jvfsp0lX2PwZiIuyGBG5uNY8GSrP5vE4y4gjNm7bNLk5TaaQFuVLMEkfhkHvZXr
+yIdfTyLjfW4BNsOF6LW+fb8r1AjXH1ICXOOa2ZrLCMveWUQKje8vusSVutTjItH/1ugiTxk1OL7
6PJGBmXynSDb2JOFIsGJVgQ/aMr9BtmUaTxWMElZss2t65dK1xYDg0QzFpG7vEmPtSv04fKBnjg8
HGV/ZgEpSyL9tHcD+wUBkv5u+7ixMUqwDh8lBh3aqFx2i13ADyDWffmwS3BE2fJqroB/CQ7pepJE
IqaRJMbCxsg57lypfE0PuJFcIxbox0xWGCIRNcF98ReL27Xzd1ldjFALB+OOcI1FY6LtL/5y8JBH
LhjbK/4AuCDLyfoGylqXIM3J4CTrVDKy+jC+buWQfAlaR5OT2cDI2b06VEDqqvNtXqkbxPO5Ew+k
IcXWa+ETPfvG3duNQoBhhStZtfLaPnnR9Pi2vVuT8RTEEcCMMV+Ef/Xks/o8FoYKHvySO6wlDjJf
hhvRUoT3KrpwKrja9tWk+iTj65K7XyBXzkGD5TrBMgEF8+U0dPlMfP8+MPxyldvRFIMzeBftA6uj
xrYIZeT/Dz3b+DlllfNbMZ32XQDDCSrAIvekeYPt+zguRndJmZ8PWqTj1301WfP9sFda+uFug6AV
OzNxVo0VzksMK8L1dIGCllvk6BHcJREIm0137C8tGVItBGARYzY9IzR8mltF5EAx9tdD/tlVx8fv
VmOO05K/8m1pL2g7A3oy0dVuD8q2X7rhstvstmaL+xKVXe7Iq/m3GLPthXu+6XeNwMpd1z5u71dR
RkFnp9xzupVcRZFrPOiE7wGTzMAoNaBApFzBqCCQRygeObCwOu4WxsF9y0R3LeoVzjLDDFIgtCyF
yR29fVn1CE84ymfISMStErW6py43wYvxMBk8FzN5XgI+OkFF6wB+JXt9mHuQ3qsKvkocNslm7873
mCVQYXc51OA3wNYFpe+CS4KWWMTUJAsAlby83ykCFjIYfIR5wQw2jUyfxMSsuFvwTVyj69C1EGzr
u7Ay5/Mt1DFsVGo8rHQdIwrkfhAV+bPqtmLAU9dQzPg4e02xmezVW3VFv+8vVaBPTomYfoGL5I5s
d+7qIYI1qvyQp2muMJUhAQgOwWxjr/6KPSztUYzsBRRV//nsEkcN15LaGkrBZJvyvc/DcH4m1INi
uPRAYT7tEDD2s6dItXK8zPHmd3QUkj0gEfyej399FKNqHWD2TGYGdbUgDFNgjzxUg0hOXec8t98G
8S9KSbzr44t7lIDoiOfgUIqHv+3y9O0nEw3SD3NvMkFmBDIFK76lGf6mCnHCQsDwZz8lDuZtRBPo
1uyDhb5v6h1EDHFPSJzahwF7r7uIBLYDPuxRL1bSpv8EnWFPpWaPRgpMuX67/F+fqW3WrzK+wYyH
3hxA8sfZYLu384V2BLvjN5FgHsfj8UdZFVFMLY0sxioFaNCJpUORbiYZCqqUK3DWcCeYF/H3ZsoK
AyfX7pBKm1ymcWVIcfJa89TDrSXMJchAes6DXdUpLaL49XLr00X8lJo6NCpuhvsD+dKkDQ9qOGa1
uYijo4tOU4MjmboEVt/dlxh8w5Fj5Kl4nHMqqjQLkTmjDqPTNTM5bGAE26iqQvdedHPcEBleuhPt
gJ8fLzqrsGlaGDAsLRfgb4Rh9L9qoJNeUAevgRVDaliHD9h4KVQZURu5+baKNhNRNWeVmNAkmMhb
9qy/L0ItgZZ5GJslmm3w42UgTEIlcjvRfoDau1EPR+RS7ZsWSHaseywDBHPSzTC0fqlZhS3+1wd0
fgbTQDYMaRfpfotkDDNpHqDAe0JVDOo3muXJngaDQskOWB+eMLuoZsN0NTIh4VefnwZ/6i9QXynu
uVgkXkRqfgrVHpo12lRp14kMGKozUuOxjNkxtctTMVlj0H74Vlmpp8SX69TMWeNCV27nLp2LLNFG
5QwQT620preC08bQZdGB1yxBS2mbUJp76EXxbDjyxE7aO7zJY3s/4/XOGpwq3J0NtedHmTG/HqY5
icGffKPHieSVAXGPgjxCKHBUo5N3+Du6rd53kaTnWG6gfbFaQ/stuldbIPoxKQh1l233Phuf5OS1
wKEDYaoKbj+lJhIAGy0cAG5Lqkg5jap8UPmzO2GPKB2K61KSiXpC4NB7UgAaHL3zDsruR1QkvhRI
InFRRQs2MkN2RYJhlBJJEiFPy13mXBiopfpicmBrwJG2Qk6jp+HAWrMKp4URRkm9eFd0SCFHXWtD
jzc0X+KrdeNOUmZDwsJq0cxKZDdiPlfRCoXLMznpNNe8y5ypQ+Kt/R74rbHX+EyawoLx9c/2QZKA
2fWryue0pjlV1uaHARv3q0aaTJNyJUbJjYsdOZOYD7kSzUiGUXSYVMFTrtzq71L57wYmfKJZcS6I
I8ys1V5Z6yocXAEo+MHmE4VIhV0jbCMLek2z4ZdFzk53ejXlr3VG3HCm2eJtHm8kam2KXSBLjbei
9aS/JDfQ9CkwgJMqMTsqr43JZ5ThOWNs7x0kXBwTrT/GPb1Jwq/iMK9MPW3QjDUitYyeVpuUlcfl
RCtqEeMOk4HpTWJfDe22sykvNZptLJAiAfDf84z6ETO1HzzoeMOJSDMrGzuy5YIXqXoY9oX7uY8j
sQITAL1lj3QpvDQilpJJP472PiSuvUlAfqIApGdwQM8Zao98pUTNlhkOsWcUKhn648RR2anHVPCm
zzlurKdMIA4l8mAs6CfyHoMheze34IdoCaHwRRqS1PHu2VaLF6CCiFLUJV/tvfdaxVAJjfTkL/Ie
hhdmtioDE9UVVksRSi5gu+q69PdVZV+CnKjUydrThsCm1UNbW7+gLyHcMrnJTNWDZ6qbHq/W5hvH
0242Oyp9+gstD77GIM2UreVyNPiMJMX4V/i7nilZrdR/1PaTopHPxJnRemYfYjRkTUEuTp5TD8Ix
7wW9gbFcbzEw7bNnK++bOcobWlDiaW3YCq0d3WW714nsXMtkNDs0yIifb2Sg36DyfWGa5tZZyne6
BV/yG4VomfPmPbNTw2coeeyXpCYRsHtaMrr1+8HJ6ZZptaNz6NcsBICUiFZhJCcxZk05OzRNiedB
Hzo5IAO98w1cxUiCmZrUpjlCv5xHKNtTBKZVK30ORqH1EvUqg/MkJDgTJ846SXnqSgpkQiyqZmYe
gDknXaRhAVsMgQ7ZI9oUtVuLzSwTrSxOUOiI2CpKRt3ltJtodpYs91Y7nNUZLdxC7vljOrx/KN5+
49SJ4doAqDMiatUjjFIkj++gcxW3qfgu4FD5kG6qhwzMwDiOMhev2pHiS+ZWBsNxuiA9wWiVGFcO
XZQfVv41hmTUHYit5pI3LFqTpfdyaM+UAkJBGzEw0+/9pFUoyS846FoWa39OgMZGTk4YONyD+s1V
R/HyetvuLix2M+wQEuEdxpFod8e7a/R8bvWZxcxh79yQ+4Bwwco57nwNUz2Y+oFdruE5+9v/nNX2
NU7vVUXzkmSxNKwIBe1FE5s9a0tDhg7NmeQMiWxXV76ZkwgqCWMqL1UJAF4GL1OoFBNFxOsJTxfl
xwmk3CeLJstnU+NFpKoGf/RSsg8xuHIxz5lQC9hmWLOIUyoFMRfBRdXOmhPHxykD9/ZFthvLupa8
qi7wNwnjH6LYeW7wTKLrSmkIDixbFtoOUwNXPUlZSF3TjnH1aax4Z6JGndrEMnmz+c+e6yWAboh9
SPq/mI1zURVN6Ji8832IYaAgvJOmYotKMlfXo/0fpA74ijVFwMHqTdLM9T3OP1nHHm9PpmrFJyNp
bWzN+w0d069keEFJG+/S4D7Aku+uEI9/JViXV2BpHp9n22QBwucHkmTd4fnD6xCvCAul4TvR98Fp
3+p3bNHgu/xDVz+9eLd00iWy+EeZ53VdVfIK8b8dAS8Pv6iZC6Qw1RyDmNblrpoqVzYd0GLC7OtW
bOWRPZaOBDhe7cE7CcTkUJEEgJyIhtn7diYV6TAPWvXDm1K/t+LF2gce5uQf8Ke1/q3EFsLRMSz6
h1ySZ4y+N+51V6/P4L+2XGINXbcSuGWPotDzirVPY5goMWirjJajZk4116rpQvYzqfr/rnNEQqZO
UfMj+Pf/Fqqr/3GApnodCLQOAWwK3OeEbSraLhXS0OQhc3uff/iit//wzxcGmKuEQG9gBLLUE2ZZ
FxJLtHQBJnoazEOOt2oahpgmM7MUtSXTOv+oBjphrwpGwqcBhyL69c7F4XYw/ejccaP4lPheJrDb
PD/1g7U+V3FwMSpAW3IOeO61X2w3rn8EnAJGodjd66H0+hY5pBxIrsdDdEwbP3+JarxCC96iAxU4
lEy8W8UdzUPq3uKbjjslQZQm4vgOrnqaFfqZmtdT9M/Gy/YI72HaCO0YaH8KJLUB7ZbFg/tOdIJN
T7k3GKKfK2RmZbs4xK3pTEEiD2EZXjk5vFzwugapjt3LCNoTK2JuJPdigBDGKWoTrxYQVfGvGtoA
612WWOOhsIasCxHnBx1R0t0uWvryrkvMaW9BCkzUDVRdv53cv9dhMVPcTdHtJDAIYtLDL4okwU2f
OqFmnu686MYDTs9cbonxRxTSY+VjcFRhm9iuDeoUccNoXZHYdPqTh+fhOG3e+GoRJ8waZcQ4BWbr
9rVbDLk2OcWAfORMBzk+CxDCTM1IitvpKndUN4HlYhLlVQ9043w1cAnKW2umKGD+n/br1BseVM+a
SgHeaY11o2n1zs5nPhguX0qISyaHrwJU68ZnkA51LK6ZP6OTXlAmca4m4H5Li0NGHrce6i0ndzdj
UxjU9gQ3dkUETWPBZ5A9ZtZnoTMtB9muK8S/ysiPo5eg2k2GU3xby9Fp65p1dPCJHh8tYGRYp3mb
Ryj1H9V8UKBh3EWGcZ7vJjNjQzhBPrEpeEobW2BzzkiahEcoycmL5l/JMifXwJemx7xChrj8yh+k
ME4XBtLv06vLX3ckOriCPYFXdoKogbIbYDIlyUpEiGu/EMVyYiCCukSNoAczs6jyV0msewSIyfOO
PKjkaIwnxyfic9F+7iajAXdSK/eldYtUOevGlR/hqeOoKxLGiPe4Ff1OZi2x3ir81NTcFoMtr0Oo
ALSqNUCM6Y7nGRUmPgCGZM9qzmTgf88Y1M6dcYFR7Iq0bx3utyMUueu67wMUNnWqDzwecpUk/9We
r8ybshCx+wJOE7KkvqtxsBYEPZ2VHk+hwPSBmoY/sarAXqftzjkW1zsrKPTGnXlTkqYez737r4hF
Bj8Od7dBmbgSKd0XvOB46WfQ6mdC8bzZbmTjzjGDLhV7R3kdAamdNVH6LziCxoW4eE/AcUCmpdy6
8rKMQyxfk/ZWap2wALEbBuO6mU64X/GJH2xck2DYA68YdU7/UBXT4RutXSSoTAIEciOdQjg8cRxA
UThdWKD27pWvTtayP9qxgRAdCVXJ0KSHFG+F9sy4USUhskJYZce+G87ZUDxrWkUBjabJlPkIwd8+
W8I5fvKkKb1mYPHUj5pWk7yjLVMc14sOzJscnyroj9iDx2vpkArruWAFKZuaG7Wm2kl7rknf7dkY
uOUHH45gnWLxXcB3EbymXIMkNv4ngBXPICTxevxuXj5FazCS/be0Kp4t5A9LiczNhbk6ATn8QYEp
naDEdnb5XdXCRSghATMXKhcWp/r28PhA68QHEFOLOpY7zeZJtsFZ0wurvKGOGJ2ecWeO10qk0ZQP
ogYOzSZFnNi4Q7MH81QcKcOEd+ci6kPz9se0MCGKifgPdwlvfwGD27UTRdmIaCJkN9VYAQGjASiK
HQYmJocIAsrrN4cVGAZlhzTpO8MNIL8eFV6LRhvW0LkDDKmleb3rOewe/DZxaLjv2JgqmEpn/hs7
2egEIKPXzJ9a0z/z2agJFc8W4cMPzSTEp8Evs7jnC85q8uelJl09Go9sDs9xG4yRurMVmMxV03R8
eCWDBhKs9PiTdaQbNGAqgbFEYkD+lj7/TW/dt7x19iNph+G71SV8fw0tOi/MKRltG9GlZLk0idYv
Byx0eiR6+1d2+qPvHcsu1gBaElxbVb0uVPqHOheyMi/wl8tCztKKj/D/sb9SRhYKXX85+kZOqcNm
Zo0Gv5N4y0hwJHmPt0HZ7CrZAAaSAJ5UZY2cyhiz4mUgr+2cfr+9SSpsMXG9BhhWxYiRhyRKRGlZ
VWMtgDPELd+p/M0Cj0DxWeZUMJnqTSoZ4YsX3/54DCygQqWswPZGcxgFwXdjIiWw8nhNFFnTVMn1
3blo0KGCB1hWUTdgMJvchRfPG448FBVjpPp0ge7JaI+LmqkqgOX7YI7BszIK4FGe+Eq3r9SDGXWD
g9oGvbYKyijUDI8XNkSIxc5A1n5OpbJ6W8RS3XFnWIGeYWp66WUFO2OwVUZ+E06m0+RGEIXOoXZ4
Q487GFft1FfEdXuJiggh6sGPB6dPpOufEPvz21+RSTstjY7l7rf82cm2P+FvXURX1gU26nIxLk57
PRLZ1BFb2YY7ogvOrBbmpnPwSFubKy/FkjWN+gka3xTbcAFquOTMy2+s9Vo8i9Xrby+9x5545dzr
eUJM1WVyS4yQ2JNlmgW1xu1obPs3oWst7Skxc+Lj9N9ZGfyi+EcMMib9hj+gjUIGqVqq+qvU1tYg
8LFK7F7L+aeAXXfQz6O0qCe69dSqFWVlAjpK6kGtSk3VTgo3CCfXjrx5iI2PnCJ0SSzrsR+HuZhy
79Lllp1suwl7o5zwngKHpzlZhQmRFJNsaL4ZgN+GxVFx5bzvUf2hVsggNx2OhZsy7Xx1/UEVXq4h
eqcD6JNwwrN9QCtwZX+v/nnYosd9IGiqpLKHhQMw1QbmhbfSrrwyH02saaNHdbe2ox+mTlWZS4mh
k/gvQ07tYHkCiJM0aaHkMpUPKXT70OiXheThfg7KMpfA+aB9oRaeJtM/CGk4ShaEasK3naR5bdOQ
GTm7nBmnbbaYMj8VwByvj1AImhy/K+ikePUb/Mq+zgkmF94nAJaXtXoeMyxdyaLsnfX/mF1SffbK
066CnQaQdXEdA9Td6hTnujJnhvutiDDz6sbliEXElglaYqms++oUh40WKtHxyjbLst/8ptnyZhmz
boqEKssBVWCE9D4BF8DBS2hbmlKAUSXk7Hscm7+n0YdWKa3LThE9yrZTKRHvx5MUOEAoqZVtVXD9
5AswK3b0/1P/hQH+QS+SPmrDn5bS93GBvDCRAEZmLb+I1pL4gfiAtP+v6qExKq9xaxkKQj6uEjJr
3oIRgyZnIeaVBDcrZkXWFhziJcblPIyh1MgOZtBpwKWQK+cn3/zhuhMjaUgxguE3t07vYOyprSTg
hwDseJ10paZUlWJP3RBy+vbegfOf9zL920JqR4ZsTRi3/EyYJ45h98grlEgA65wMgxfUMoTMfAV8
UwyOkLFKmnIFOK6GfxPGSC1E9C+VkfZcx3SI3mzIHOi4gBAokcY/A+khzLCsS97rEzi1LzkybndN
+6oddoUE88SC3eJUBgBjzOprrJO4+Gn1NE9PYu04OwT2nZ/Lg6zL/HiXGIm08t6JkqGMJNV9u0/X
26zkJslZvZk/Ok1XjWkSbld1VzVRza+sFcrA0fsWK81ZIz7bCVCV1L5pOieDd9z6GfTEgHUfL5VB
DWC0PVo5VMnH/NE7HcOiggQr+6J2pT6QNlnJ8OUtjrymoCJfImEsTKXVB95Fr+kHx2aQBackuX1K
KmBOMO5VFkfjMqZacHwSYYQ3CgSLzyRHPkoY/YavbOoEQT4LihiFJRt8PBEU5Oj/3ChW5e8G/g4S
NoGZBvbMDSN8qBLdfiGsbh0kAU92v/+m3z94oSfWXV420GFEtT26qmzcZRXlln75ofeCmHPp7LL2
o8nhsH8/ENDrDqC0hMS7ayR9hzQSqeX5ORYb6wgjJIZhMIrVR7ZmT6Sezhsmv2JZ2pguYlcSulPm
xLURakRdgZvAPF02IROfrlJ1042mYI4rR9/ulD2TjvDDQkSTfqHuZnAAD42YqBCWPN2BDhsOqWhv
dNRaFip+YX6eiRE9PnvtUzBenis+fch4onAc1Ymst3P8HROsnWDUthiBj+IEnVk9hf6/3WQ4Qn8Q
owbcVJ+nmThCNt8W0qz+vuaQpRx7lE3zJylbiWHk8ncDrnVzwYMsYDAiaD38IL0KoDFCWEtWfOA/
9ccvR2pSpsa110p+4EhWFG9UI84MmhxqEQoceAj9V5p7u0z8y2LKsmdsMHG1IaF29epeO5sYuTiB
fnwChCT4rV7KDMf4EPa1/zoM/ZgJVQ9zCO+plcsYeNKzXRv0vXvBrrkyJiP84yPvag6iZqtSHu+5
A4tlIRc0NjP2XxBCeCP9tgSS+mOxursZ6Yjxexf/2EmMWVgMjMx6cQLye/R/b5823mgxzWe3e+ZK
svMbYlLeT+zEMpX94qv0lbx8ROfKinHZpPouS1lEt+Vp6CI25nGO0RCbVtzFrPg++5KmGv17D2HU
7xQ6kxMUpD/4wLmivAKmsu3BFSq/lEWOrQlFMSl9/ZL+1JzngDyXZGQs05SiddH/SsXup9CnkPAa
nl3uWW6auym9yWGBK+2oQWDZPapo2+jsB8TjDyGqrpeW+M7OXznYhnhOptBbcLnBpYhWCrjeJ3wj
phZNSWm+rDFORtcUdfwtg54dAEdpuTgMGN4AR9S7m4NfCGYlMuLUeyqQ3w4FXOK3p2om7SI72lCa
F71BRUlKfrarPzmh2hV2TxE73IThQDJEfJzF6vgPXIwcSeX9Plx+sk2wr2YLdajcPDRTqn/skFK8
T5ZW4ZDeL6RvgzPkJdPacXbM24MBVCyWV9qEwCofmK6mFpP9OXAOp5Mc3nv2UqpcL4X1g+yypKH/
C8vhIR7YKsXCAWvLkKay2dICSpem68MhnX77jPkVP/Zk2t3Ni/mqHD/8L1EfB5JZNyBlKW+bLFPV
Bct42bYLDU4rZB4CRHSyHBwWUGUDt0f+zdWQMsr3qv1UPMKgB3u5+dtgCbFak5UVzu4yKsjOAkvM
oO8IOXdorqrkADP53gH0oNWr/748CMvwpYE6VFaMe7AChx+qUizZw4gCajQW+vDEhGqiToTN/4Dp
xwSV3Xs00tXPfQfoUkSrSTK9ait2XWo9o0MeBYqsEV241GcmAHm4dTfvxoz3AEGJXHhCCKQu9j1u
tH9Dwhp3x87gAgCHXHUZxGOsecXA2d++AA98489Z/7PfcFbTsKrbNuG16/1oEaY6Zyf3iIB6mM3Y
qVUuzkmvqbGqCMva5qs1OnMEARJ47Z+RKEumPLijGB7sGf5zS2ENH7hxbcaaUAgZu+G3hQ9CTs6/
Jd57r3PgmuX+zUx0XgooxWOhJyzneuzRTfQPdorOnPMG3N3pem+8OUlPDlDZTMPT2ejagdN1EEtM
wnfp17pAk1e4lqkUn3BlrqZEcAFNjrjezT3KX57c/eXUtyUUsnQDYJH5mkWfn1Gw9XCOhVRhTgl6
duAwGpJPJzMvx00ujVsYCcTdGNW1X3QshTpj0DBxuJgMg8Q5/BYicqFLQaFQJzSHzX0ycpPhurca
GhxtcrYFmmCVoJMM5ktrDerzdKJGpbKZhw1tLTHTxEjg0QdBndKGonidQqUdrB5XBI1BtIbaikSj
8R7Y/YUTQdzKRGZBkUJcrdoYHPUzsHD+Q1sZEIwZt43kv6DRGqAQeebD0OEHLEOlQGXk1SWJAT1S
vs5+4ZyWWfbdTE85o/zCpnXtNBE/rBheWsioUMRAxf1acpfdO7r8ruAq9SqlupzlMqBZcecmBjOp
lAIYkc45HNPMFHl287WolsEk2JsAnqYH828B3Kc/njcnShDpBbAbMExsybPEu2wcz3WtM9KbX5X0
p01TM5cJIld2DXokPPis1NNgp4z0BIQivDHUAiLbagGwSc8ezCAJ5HXrOmcXIBovY3YTpjb7Cj/S
2oD/8QsX0Ms5HpGEwZs6Ut5w5E79vxtESP+8CMdDerhSsnfMQ1tBFaog/1YX7HfC7BG0Jeb5yIDE
h/H8nCprQssDUrHNyyNdx9I/UYABnSZy1vrW0Gif9N/xpLBp0pLcrL7vK73GBIWqZs6UkSJ5JkMl
HA8zbEmGDtuD2AJG5JOntdGlXGgMlifYzzxPFV1O6cXCWpUz8R0++pQL1fSBh7t1EJZ4fetPszWr
gojHw8tvWQu7HJ+2HKb7nz2B6EUS5KHicndAgS79BR9qGCJiB03Y6fUM1qC83eWMkzhy7rCIhXBE
s8D9HkvBRNZbEEaucpuW40rT+EYGlHUy/e9tysEIVSQzxf1J4dtbbHe1SpGEj5JNCQd/lmaKFTIp
QjJv0z4x8ZRtY9eMDj2VmdtwfO57mR1G84EFKTkvj3PDzDZkzeC/weVz7S3zerWQFIC4SwON1ccD
r46oRMhZLop2bMp1y8f6//RzoqkLx3nN54U2nGxAamI1aSJiH9P/xgFp5PiUhW1XF1KLMrbPNvn7
i8tPfoqiCiMhJfgtMCgDnn2L76YRFCTe0qIItdSmS6VpbxSDazmsKhRM6V/uEkOXKRe7nGd4eNSZ
tbgLbYCn+AVZfWICpTU/WRj9oxXogZjFO8PAj0Ee9krs39r7UKNl4y8LWd0+DJwcNUxC8EklxQGU
CWcwnWHtz3x4GUKtxH8h8TOLkQZkmPmlhhpQJY1gCuY129xWx/Xd28HvTBmr1KXCkE0u8kc5HAsc
KgZuLkCuXcrheJL7XjsFWtR/RcZ/6tieEbXQVzAOfounRA4VyC9bLxUAIigno4FTxgPaPuD1RUOO
e4m7dTadtma+8OWhJ29fP7ptpEeQLmpnF1bSX+9ToPbAIlZn/6jIiiAyAb1P1RRaDLqHrpJx9PIq
6/AYpKdk4XzN0NGuUN0dkho8Jl/QmMwjd7HwuGyMuLtLXQtKVD1oVqjgNeH1eDIAbd761j1k+b4F
rT7gh81CicekUjmLWTsC5F54yiXP6IZCa1QpE7J02rNySA1rW0PWl8EJVg6NxwXtxxE+2+DVjLJz
om1wHRvuAL49/1wpAUF79OsCXyayS96m8z981PA0NRdNbAavMf+ouJ3mrQDOfi7m/nUt3puGZvvR
DMtl+JYj2uJB0eZkxvEOcdiwSXX79nr4U/T4GBZ96a4luIxiqT8dkY5lnQm4HoV2Iv0zdC3GiyVA
VMOsvPCvbYcbPnJEhyj/ykynPIsl/O/2vnL+JSqFmMGzgilnOckOLux0a5EYkgZpI+WTJ29bbVRo
l5hEZ1qDr93hB8j+4a3bQXBG6fU+H8IlqbrQtZl8K0bHJhdRJXROzoAWb4uuhUtaajh8aNHRmUFG
M99WC59LzJJpfb7wGbcpM1QwduIvdFv9yMsbQ6Q/zfMYD5YwihCt0s+wsP77y8hTi+SC4JVvEKOZ
SjZIBUn0zQZPiO00c/AjC7ZyncaFvvU3igUTHb8jdQo2e4m17lWIc+RkugRTKFh3V95Qs+E2AZDK
N9t56n752XSrj61+iVgauSx0xpXPPB53Zr6XwWlHcy9uxMRbB8+V2KTReJ51UduPu60+HXLH0Gtj
8t9NHQjKUKunX5B4cQ5mn87L4pTXASMMYEK0/ocZM515TAyAQu7uIIQiz9vP64SjFy1Vh5mfL6ed
84dUY/udBn3mx0yWt8IHaWwZxzSnxPlYkiJZvvz1lWo2nxT4R4HKehw+rt8NCgownsySSceb1mEh
x00prEDclbZNedOYoaVIAs3Oe2Qn5bE3VeRmrNMPYx04IHGCo4nRRmbyuTIK0DJSM3ETZKkh7UXd
OUXSiLpIvIKVBL4OxEcZeQbkB2g9BF80T8s0gujm0f/Gkzsaw6IYo3YLZqPx6Yykjjcew//SyVN3
d9rVdXFQqrePZH8mZ/cgh0XjpFXKlC/VOppXVH1H1m2iPSw47+gIduGCZmYTJ/9HQq1L8thfYhZn
Y7fIia3R8d/0kIMjssx/cBpjq1qIMIdNQb/0mde5gAgR7HT8+FrKPGxi+GdOHSHQ9yV9kcbs9DJz
F7m5kBaZsYTaDdzv2mlOYvwhIVm1wweTho5G8eNqxsafuKgf74P5jyhl2de8jdnDwRA/wJvrHN6u
ILjVj+Pl8DwLunbM1Pptcqs+jVMBfq8U00s2XrNqvTADHhxOo6hecl+tdya4XYeJLgSz3Iozl7t/
2BQItwoq9yzOgYw1icONEdKdepob3cIjUH2EPeRxfL9FeeOdJzM2Oj/0/hteKG5OitLCbYX9OTff
jdxqEktrHpBIw6sAlrsTdYDNR9V6Tvokl5EA7C/QjM7qzcWTOiDgjl1XLjbVWT20fEx2qAtThJu2
GTvtOT1wwxfHExei+WWraYGvjx+cCjfmnrtQriIOnAKS9KAk3CqDqya5Xk3vh0MEw/DRXjmz6gXz
cPBL9xLMrnKR1oevFusuzItVIp8QWY8TeXRunMZBdybCryWVTYEYZtzFdNoE/aWyffkXyYr1EPaK
JjDBkAIySFgejyJxeI9uS+nZrgq3b/clTrlZO56drO33h2Hgx8NnYqha5CQpT2dBLLZwqkTAm8gq
UVGBf22ha3ZWdSNc7FhGDYdZGtqkLavEbQRA1RzhRczjhfxu4hAOPzSPm7rHx9/t0tCCatc16dmI
h/SPGs/U4giO5IgoPn1rOlmapKEEx2TIuCsmsI1poSKjWPv9QBgjum/4+6PjlSocvvNXI5Ocrh3M
BWkui/DoYERA6OZdXo1RgaTrezSeyE5CySzwduH3K0FGgHl7WGNgj1ZXcHLsL/KcFSuDvRpmHGvz
pvhcojw7audz+SaI1BHUh+Oh/mW8a43S+Vbug0JDgm9u6wrRYolMGjZAh0wYNxc7fO9wi6FFOacD
RYD8Fxev+F9NL7prSTYK6fJ+9SIrSkNxzvMUaBX/ZX4fsu43A7dDTswXZkCJ92bFHSidFgFP5e9R
WydqFqbHjrw0ZC7pA9r0bNWZ/mxoG0wQYEFhmSn1IydOYv3vSv6rnpOODn5m9WSItcEJkKMr3ff+
dmi/mz42ymdRzpC6B5TfultHnMJ6tk8r2pqfKXTXi47Iv5+zcizY1oQCgujgmVO4Deyn4H5weWte
8EETIH3PZDSO0bmyjUCc0AUzpn2xXNZAJP9M0sb5HaYvZUY/SzdIQu0jJ8KJcjMAeR8vmoZZ+vVW
5o6v+Nl0suvXbgbwiqLH/Fdk5jSU59mddq5Dhw3Dfeeu5OD0FB1ooiNF4KU9oTk6xhn7oQLnivVt
syYak3+yxnpmDEUuWIv6NOeCSBcqWlwvez0FARYwTZjWY/7e4EQ+yApM+wimecrpOsq95sObhZYk
uS3G6NB1tnbktsxDOfb2Y2IVmreap9rzLjgrToc4bjfsgb+9iiiujfwGQCwMi8UvrccfHw53DYlv
ALebKgm7LYwkNAjfXKevvd5mrFhAgynuMYxchdx4Ftv6AgLluMpiHY4dnDzuSvZW4cZ+BenO5XWF
yAfnRrd+B7b6oxGKc+nzl2yA486eLnvu9nuOW844axkffIYW7SJTNB1spfhhWn84KTgJhiO2T0Aj
Q4pYFtp0NRIW6OQ7bmQsm45vUEUQRxFPthBX1hIVLyXvSnBQQjrItnVRxWJs6c42Oedmc0jjk00H
EJ30JBhFfB94hCLdsUYSOdP/URsWCm+UbKATsUtQoxgMRPJi/WHPOhH59Te/hYALLyc4lr0Bo6O6
Y5M72VyL+xe2OIRVr6EtmbUVsTAIe2twdAv78xMMndWFqra8QQna2kncvFBP94hvP4tINlZQK/Q6
aODbmKmrEW9cXPq7a3pf20aw02DEHwvaCZUQ53+92AKet+nc1l3778H3KHIK6TeUtWBcbAnwKIj/
OqMEwGoPA8TfrD7nn8aIeJ7Pyki5vkMQxi7IWj5x1kPFjWfod8WhuA+TYiizzZyBSZNnh5hq/Y+3
ZddQijuSJzYOem/hjlLqPM7l5mlLrMaDWPR+z0t92PvKFMBw8pkct2I+zXYdORltUn+wF0S0umDH
wiAudG9UgkVr4meX/7+34dfa3/LRSjYqayDkJYzQ2MvTdDLyv6Jd5x9MfqXP2AU23SvhEvn0GjyL
hYnEe5PKChzUlD6LWHLedDgweyGSzn+QjSJ6Vc6us6Ki08BS6iszls2+FFI5oxSMM8W1+kpway15
97lG6f+uUo/ASBlDsLh+pN/9/O4kMv0HzyifU/4xzPWJjZuqQ1iBvf3gYOtEtYdkJsRIcsguGJ7S
7yUtIiOLeEzLn63ytsrgJOuFmQ/1RDeUC2DPtrbhmapPJj39T4AJua60f0FsE4N/Sp9UkYRKagak
A+6rYVLvqaRWBqgwyujuJLMRaW5IuG0kcvNIsgq0W/nbp2Tnbsm1mbqyZmwlG0b7oQIVtpNadlI2
oEOKPudi2EGpxSVFWQbd+fnd2oIC+6pSLjkFXPXnp7gTryG7zDy9mGS4P3Lv1aASuxeaOoWWdOk6
i9k8P4aKG//VrED+EfRtnY4k8VBbCFoLkbEi76MAs0vOXuwV3ieOzuIr9ZlaeT+MTw4Y0epNfQdI
4hD/2LPi38iplhSVUzB9y7IrOfeGc7XgdxJiUGMavGHQyFipd2O23gqWSqSV8HkIpW6zQa+WKpxl
R+dp5imTw/u/HY1//P7mmH69MPbm6S6R7kSPtB34IpLSR2NxGIUmwjaK20tM81zam1riXWdJYnbc
MqGEzNcuyeZJUvaCejPrgv6gHEfB2EG40PLX/TvyNfyeSabc3mvRElqG6MTTsgQCG+B/vonDjkLk
LFwQ7dWjc/KLg6bOpkD1zxvRrAqw32qA9AEQapePhKUBZI0KO1B4DelKn9Sg3GW6KBf4VgqFbUAb
FHWFvknEsfYuqFYzLDvjkHVlWB3D55+7MbrfZX9xqkRjn/adD20dh9jz8c45lpDaN+DXPAXJraKP
tnRSUHuO/8Y9ECv5iu5BFlWBXW2/VJTZxZ2EfcETgB59oXhCf0Ffu18Ulyp2daIZb2Vnt9T3CfA1
9asIaNYF7Gf/p/nmtvvRvHdipzE8ZUt29CACmZuGGyZ4GEFrD/XySPggGIxff9yio2R9+6Wjt9Pv
j1enwkm9eBOB6R8fXvvy5MRhZI2rA9ci92UhnJ3AQSsIHsdtpSSGVM95PuPP1ctzmk/jKfqVL8Uj
4dJVxW91Y72qerGgeeB0oXjv9BuJnWOHeTTKBW0SOxxRjLMAhTsJG/OFlBLpCrn8FyQINeI6W8AY
57WOR6RrlVrS+GwfaCINsCo0yedZB/3g/d2cCer7V2I9slkmFibk+S586Q96vKYkkZnNLtnXxjF9
dWWX6HX4sxmmOSjAu7QKrCadiocFILklyq3hUSQefm1i1/La1fFxrVXBnH5UlG89jCHlJYfm/FEN
gQay75/qIobnZfK28mfFvzA4QS6wZIy4iXTjEoC13fGtwUNieDxXrbxtESb56ZxWTInjjIeBfNne
RW9xEHTRS3TbiQTmKeoN91PSXK6Y3TMxJuCc32Kp25IQCcQON2oF03Zftwv34bsXIhwrxlMTYgha
VAtVXNF1jJW9kbK1wkKbb1WwsENr4m8k1+l1y58xpHyyx1ZUAhaujw/BjT0OpPpYNX6B3HvSUzhx
n7Z6v7kLD6KzZ9VwMFTJig3g1K7Li3uQVqvw0o+ypMsUMRzL22BM36lfpbp9p9GReufSCAieGdus
M4UnTbqQwsMV78rZ6dtojp8sdwL+NLz7bMMdfno6xMmNB+ZxPEWmKmyT0ikHCXm6sNGdW96GTU9U
i5gZDGwcPTJSsxtCHV98mSitq3l7HqXg7SMxOWGr4Isr+3xkRsUh29C02AgHW/OmcV5S8KMQP5g0
/ksqND/jzewhQVSbiGjBbIWAmu3U1+IV993FMTMe/1V2QLZjh4OL/UNPsmo1udwNlec52V1QAKed
NULWWcHD38pDowG/wdI0JeuNJg/U1hlguntFii1jL2e4IhoVxHcaIS6IgjrAez3zdCowb/k7QqCv
9Fhw+pd3i95p6K1CYhK0KJTyo8qjS1XY6P2hRJS92aUhEW3sJsycAbnd70kYh69DjVFfFxRjANIU
y17m55xbNxtVXtzPrHQzZylmG19hu9DNhXXHveKkCz4sPKR1oUzPMYZ0mzZJ25C7bUt3ySSOOmxO
1j11AGocgHSeezXSZ2QJr/4hPaDZiMR763QbUQ25SoBSb5elOpbDxOY/Mp3HsbECU7TAxW2IxOrg
PjPLsHiLpnQjq09npg3cQuSsNn3kyNEm7hIBtxyopcpLXsbmKyYKL/dUVAnh4r6ejMfGWlLzfc76
yrvl5o3Mf9EHP25N56OogAjEXzhumz2Qeq3qlzwOJ939WNdIfVK7Fz3ZlVxGndxTQOe4iUR9fxkQ
6Uuq1N4BzdciECMq+KS8DuI7QOLIgzAFnkBUuff9ddjQPWZDA54F4LYk9IMzwZCWOqCo8F4i0QG7
Qa0lhwVyQHUIyVmG2UK/w09qLPraRTNvOR/FDqePhlYqH5eQvxFJRfcdfY+mpM7fglw6VVDcHjQL
6Rkyp2GkfppGPD5V5Pc693LsjJKtu5uAw9ysqehV4EfndCZw6GhUt4vWyemDiEN+D2en7mIeI0z1
VY9sYidUNY5za1YG6BdIzuARVaE6JZh2/SSVN+XbNL0ZhUoNVsxEce7X/05YimjFSMLj0I3ve95S
/gZsePKlV6pu4W24oh8pgSdxswByDJ6kEU1K+C7gDWeV1quPa6X/p3I4Gh/pYZMBsIklug77UwIy
xbX5KE2N/lGCUmYM67ughs/OO654wBA9hsE3yXr++weYLRX0H6PyEmGCvaQY1CAv+VUy8F611W6X
rOgNuc3mcEPtX/Eo1qL8zK20jSyOoMupGB4xKzWzmgH+wPl4xxi2/8o7H7L8SSpyCs55KEdIveHZ
N5Hs6j0sWhNgmbHGt971kfumWAQPBIto4Nns2E8XtD9tasyx8m9MKG6aacvJ7tfqkEZwRyjm163A
J+o4GaiMjiUYYxr+vSPgbY9o1h0luojGXLLSD3b5LlAlLOub9ZR2l3PbAO27jRQC8wwAMjZ7k0ZR
fVtr6kYc3myC80yjkjOgaIwrPpNTGKoJYMzY4Upw9QdPoPIrL+bzy3DcKeVGU8d1wfNTbxi5QnN6
r36FJia1ZWBARZSLSebpkSLu2ZPccQ4p5JaNTMz1Ryy1v9LD60DRXgmsDOmQaO1p9DezzgvSjZrM
zUepFYYIrODzisJZmySgLqk2UZw/0RIcI99FOXi9zZifnIzDbelOyDrTyQiQpMy6xGQWrypUAo6s
NTIT4BLARCFNjfExtJcN2LWII5J4h3xlmWQeIFJI6DPSnTBs22F+ypms4aus77j2pceipyDEmPFx
z2cBC+mwyonlZx8HWw8jeCVlS/AZR8reGdH15iP9TMz8u/OUHkBJw1TNbjotFc6aakLNZREjQHPI
pjKrToX8xeSgYkHD4RsoDiEcCCr/rYRz/zjsJjgTAZu2bfyk2ASU7OgPCBBk9KkOZz2430hJQk7K
fZZubLJx/ZzMIByx5qYE2pIA8mJqhy5SzQeygkM3urfFDf3QL62MN92z9TPLqa4gS5W4jqCo2031
AUCV+9vzEGspaUF2Zab3KEcBlLprT4oZaewwynM54p1n1JOT/8kgX8/C+occ4jLH3lGp80m+xugz
oNiNDtjWRUsTfFU0ZYxzFhskkflzgqh/mUTTR8P4QvYliACgp9aiueRyUZl2SOI0OXB4Ei+U5V3/
j55RlA2mJy3Yepsv5bmLpGUCP0Kc500M4nPxdqm+gdVRUKXL+tykj9qQIGrDxk5PAzI1ylQ0Ym64
ZazoXGEBCQCYQxtH/Aj2NCWMG52q58Tjoxn5+yfbsIwOq2rUoML9BUjFjPpT0jOLBa3CPmViC5L9
fZ6APiOnvoB1hhmX6h384hOtCN8Adsked0I/vpkLSAPog3AA4s09IkJp+cJN8xV0hvajB/IRqjkK
EwHNj4YXdf1gbA8g8V1OnBc4cEl9mBMe2l7xoTfTC4SDt4EVu3TMmD7mPnLCwfFbkAT4LgXgT5zM
KI0QHgXRRTH43cYlejPZYfs2Z6qqpyMy7qeJ/d2JjNZ4tzvuXcqaXepBLq6/GkJ0XcX2w2o13P/A
izzs4UUMTQf2yIpvdZZsgp2iA6L2yY+BC/qKMpQPYlmYAE2hmm2ktb1adVq6TEs4VNJy8cy/AIg7
kAu/74zhKo4kQzH9gDloPsaTwV3V7PwoQXFjFE7Z2hffXIpCqu0k+yXA0gkqvuIduppWv8EvgRGW
ATeLOcxp4pNlFQ+LC2Blcii2+od0wHN6ELdSC4mksx9oiszSNUTfkco76/89EF8zQUCdfRbGk8c3
e7NbFmATg0Quwo14D/P5MGhwdliAkth007b2rGp0atLuk+QLwAVlUyqUs5Y50SuHuMxVqzt5CXnq
OGEQEQ4UBd6A37UG5NcsyYx1CCMbH8KybNwbhMs2o7750vCM3glknGlSqWFAh6EuJiuPls5282ou
FcBYyWTKkpHPuDMVmzzcLM1k4EAPi6Q3TBXb6KDc6WLaKuH4iomzC8cqzBS++WUobbzz4TjW7kQb
yfKCQKdBp4ReVEfbHz4XUNUsGqZTC4NywXyV14LdjgyzFkTCW5kA135tqajGHRoSo4jZwFEiii4s
lkBqak8PctHNX58NYLQe9Nao/bhLfXwpgIu+Z7giPfyia119wlzFGx4hbr2hNDBGP8m8dfXDDaIy
iQCBiZmfXEk2HUFwjDKTAE3zmaH1y8KpFn/wOux8bsUbil6Ku5B+Sv5xLm55dsI8DRRUFYVGbQJw
w4NEa9usjBWf1EIwOlhEWyS00OmzaJDjpIIUKZ8WcSqO7sW0WgUiefRkmFyekIOGA1E5IT3kHuJN
SzEIBxgcSXCsjksnNiKKhoRP2Fte2aT3PIqE2EDJCOFyaSVT7jnIoOBrzY8tLQS2QtJXbcowsoYL
9+7UrfjvuD2Vsvurt7A4p85BkUPqcS8eCZcTp2XPgG9XQP8cyNZyHJColmOq15bOkYaIWs2oDrb4
BnGqR6okw9Onx9//c28dEV/iHJJKo0wJz/jLbfj4tXFIR1VbQnU7i0qdegWcO3aNB3Z0aiYttIl0
e/bgC3sLRG9yWfgadfTENgLIR0Dnit88Zx84/P137yREzpnYLPqcZAsV+NoOs+kUtK2OaC2yk6aj
9bqJ1/P9acGWsM8pTV95mRFt99EWy8dBW39JAZGf38biQVNUTZxA+duArGgmp6OfuBHZ/QFPMqkY
dU3JPa4BahyL5zZbX9gLAjLJ9fn2XV28gHO8oCxrEZNcdSNfnHm1dziNwWgk+sCyI2DQ12uRlJdi
7/BLCL1bU3C97TbuLwcbJpS9s6yomwR5ooUYRVSQ3/MeWVwz6tpBPlcENsicvBVf5SNKF140bmcv
QPt37YYFkN4hhwxf+gIYQZ4d/GyE8g4ff4nlRsy9Mw/XD3b2RakDbeEA0YxMhh+rGfbLxglJfQD1
uCzocOzdSwTpliTQEOgAYIxir/6cXDnUt4FoUi1tXu6QNCm0NUeppq8YoLSkp/Ichj/LxEqdtovX
kJFzoLgeownXBtDScTLcfq5tS1BeqA2HBjvB+cSlVV6EahkTbCFVpBrq9/6niEBLdz4FxD/gvZlq
yCG+uRUxUuyf1CFxBRkobxihliXkdZL6mPisfc1h6kYcHliQj4dEz2zYYoJvBY7yz+hVAN0qhrzS
v5HMpG9R5P3JlGr1cf2PomRmWxG8Vkru5xSVdCPCEC9u2e7VEVF3I1Wjlq/oMGJuVvIUt+6RggZ1
ykDajC2UwBYZGfYjNf8g5BfYsfYJykJQKGcP8Wbd/64u9l9ZxB81NDxq2LktbW9GCLQgTjTg5ToG
4bjuU6DlQf3wkALumdUiMSNW9XGmsGxNpXGblg3HvM75HlEwxT/FclzDfJnyltBvE3RY12smKfKD
TczgVGJdqh1V907DsuVNP2FhIykDU9/jk5Jtddw99Jr3PCRiNQumOvf5qcCn82VxkH+5Rnc9QEgk
clWWvQjU6zWbgtRDn5Kw1A3OWTKVNQ4rtYUmMW2vK//f7I5XmdtNOnNS7uvB6+/9JyKiv0u55RWo
aNSpKvx47ZY3PNBbjxk+XPWF4jREIhyh4yDgAjC9BVJ/VtqimcEMxF3E3j9tNnruWUtbdYP6g1if
h56FVBJgxHx+7X2FZzu6J3lLSvb3axbLl2xHNwCMZ6bqxdWMFI8vnF2FiKeVln4d8wnOnow28LJ0
Mh7DE/DqAT2sStzdfra7tzuRPTvELJO67PuPCJyQK5fAbOreeheuzultef1bNHZ3ADu8G2w5Fbnq
vgCGJ8gL+8Afpls/ixhZN3hCJbXClg9N5wSsJFFCwfIIyJhguq3xBX/lZCRAd4R1+B3797a3FTo8
LL3KISSlHxo7OpdaHAlF9Bh/rbpJBDXWoFsztaa44g4IHenk+N7cyL/SgPXmFLM/AW4MfebYaSUk
VGHUra/AJKd0fzqxmHwbbG1yfWsULc9y1JCl59Hc26tpw3YmDmBbYD5dyHibt83KNTc+sPDgGFzl
FI6CouWoP6kYyYtueRir3SxSzvKi4aSoQI9UDtvNq477WXZCkQGZH/NSMbtKkObp0eeXDKMeyu1I
fRhdL1ioDMnv1TPlYXyYALoAhHSXM5a4avCYU0mDLK6cQGFDinpYKYG93As0gR1UVAqQGPKM6i6T
esT4boQQyLhbugSsLU8rI1mX/NDhOeR9b3KEImGWy4g+jrMRDU7j7I13dwlTmT+iu0sNOKYKm2bJ
GBKjbzFROKue0SfazV3yK9BylIQd5di9rqVDmVz61mO4nvuxi0NZoNrGLrQPo9dCNZbdNYj09Cqd
qKC68LKqCcYB8+q3jHqETYwdt4dtYL4VTwPIoVoHbjf9r2uVjgeS4RukVTphspbdN++R4hyUuSNi
pqzoD9dmjcEqI35kgK8P/2+M8uJLcmh1TN5Qvee1GtgUPeh04cVww+HF6B18bhGFP2ENsAwIfOQK
xSeVHibKjK91bBq2ss0KPdU7BxAlbLs4aXMn8QBZfpy9KXs/DbvIUDkbr591R7kdEEVu5e0Fxxyr
G/t2EWmrjWwnEGqq0yyWAJNZytLA+EnnEiNqmZ7skTUOsUKmI4HsfYDF3icuYOs4PoD4jS9yNjGl
99kPLXoXLwebG6GsnXhSTmsXZNORDaG2QGYXUc0yGslYzRGBKWft30JhkYXvQYHg8JKnx/v1u3Vc
EMJarfop0XsjEwfXqkd9rGPUoAkCuczOOyBwJ0Q4PfKD/TPVGiolXsGh3ovlMDjiVt+Hv0rvroR2
69ohoEf8Z/aNsIyX0SMRGpIh7fMw0BEjxThk8AiunNBG4Wu2cw4/P3OgY7oZYnSWxSssQZdPUGBz
uTH6RTQdDhKyf2+W+j0xscAGHvz8xXEiqiqoQGFDMHsjmww2tl8HCjLNLsxp39FXLD0W0H+VRppK
2vk+bj5+Ty22XE/BPHBNaxMKg37hD3gcUXi+I7sD/hZ27fLnjyRFQVP8eNGvBWkeV/yQkyCsxhx2
PTwlbAn24YZSi+BtsNqKHpy6ZtbXMOTVJ60poxI1J3z1O2tHv6cP0FoEfXnowk/ehOmPdXb3nv3m
bUogZiA7xUW6DEWUUozfvFeN9qTm1zQMY75fwfRRuuMRbD9AqPP2Z/KMNHI9gearNEgfQC76JtAT
zp7wjW58htGpNBLbNVesRlrcNNrptOxiz2k2Id+PgXldl4IvHcfzknNHAK64Wj5zEtkOv2FHFAqd
fA+gbVIfdR1Z7L1iPTOJ9mC2A7yMwQPslxlmV1/zg0SM6lwZbOrYziFtB9QQcBkXYqcmHuoy31mu
9bfV9ipxVkdRMnzBuOGQyeI5Polxzcqk8yw3nvCt4wUGgvMO8UgIBZW4uR6PmbBe/mHENwF00FAz
gIasZM79NZrMevClDR/WskeD+DnRS6z3y0Cy2tGJR/qVcicHTE/kooxDBWflQql0kSaoGKOTK8iS
8sNIlf8PlcRpi/FIwxEv6S4VOKYc63i4MMyVvfT2PMY7kqMo9mhJ2hINhxIvejoy/BzGFiEjjrk2
MI69fkiN2zcJxMghiTA/1Q2THJ4gbFgIqHawwBWP83OCu28BMEyervNqXORBjun8Lb8t6nOAaeeW
J0DOurYjd2ZotQa/w5ds10tymJYYdpCh+eFcvKBZrj3q59eH97naRcyqePcJMH2NoO/UdLakXDL6
ibO/ly0HG0Mp6usIjSQ8NbjufudB1fBXGCnbQP6wRpkbKvFkZCArnmNxxmcbFrq/NongieliSlBr
E+cpPriEtOnhnQ8h7LQtYfgBVYNCKcDigOjl1bkEupLSS2Hjc9r7q/hVdDINYHzNa6brqbH+owAk
3jyVPO+19nuddROBKbuQqHMisDUKua3+0svBspZAsG/GqOi/5tfpbIBAQxhhsPG+EsRFxr19Y3qn
uphwVO+uhbcyZy8mIbiLACGPKdd33gBh1BOyK0L3HD0boads36dmkYHs2BndOpr3DmVHPylz7hcP
4DsAZ48jjPRlZ5l2DIxTzHhF3yxlsP9bPuhfbjG+GeWFG38plsn+Z8+y57/HVS4GrL+ehrLTmJNP
f8jbDvbqPyv6g2+hjbXAJ/uCHv0CnB+FN8BjC8xuizC2XIeV8KmdK1Z5QnDNd5H3qo5uL0CpU1FZ
qa3hYj5IERDSWA9vTrO6qLMceUJXdTQmsUV3eW2JIAhjv9jfLqb3kzNXX4LVAKGHhBgoyQcIn7Gk
YDxtHyo+58209i7cTWl2gzqOqUxRHnZECJ89qpLLtODGdnc+wiCxiCUxQDQNrZF6Ooj0ZZqVodVT
MvUQHggfQQjx4c4CmPtYvDEKggoRPbiENoOU5j1eA/TbfmpR3eHKGxV2Vs3u24w1mbOWkakev5PT
bFg6GjpTPgf2CO1utP37hTDZa8Au79oBwoX4xOdAIYfsZ5siun4vQW6bkcayMixDRXzapkMzsPI/
bwwyW5er/p9gBXlhPfE6a7T9uFomVgvh9xFBbluLrDQTlnKTJXwoIFfWvHOg5u90PifAxtgn+qPX
D9u9IF+t5GOL6UEjTWPckkDPdcrL8vHpNqRJVkQ44mtLGUz8yaSlHpJo8IOXhN/ixSEBiC7Q+tX7
nZYWyPP2zPJD+RvjNDsdCdxeAbtrlAPvMh6J1hyYicYrOHsffItM4DCCa4dDBquLzmg8IQ08w53s
x4ozhmFO+IUGRHS0Sr7D7ptqu4gP3ltYazBDwKheOK2MuDLaKeZIPsuv7Pu1NqKfK70zPVbECnr6
x35X7K7K1hwvRh6GdnlZjPzkxyb2auL+ko0cF1+r02LemJZ1YaJry1aF9BAKb25Vltv/X+/cPKPt
MKPN0Bn9CkwgM54zJEiTgDJ3RtuVHcerYsmu8+uYNEzYyWofEhBRSCyKNhsUOvOKJr53pA0pGblb
FUPoUTxesMMXJIUmIMkpu/ymX8LWg0LP+mAfuLjNswM8Cmx1ItpU+RSbYJ2Ulhv3UbQ4jLBeZuEQ
kY/+uHWGOQHwb0OgWX+0FiYLU9g7RJ7IRozd74XiRold+bzE8R0+l32eY0v2F6d+MUOvdT1ynlXP
5XhjviodASW2/Mqd5/q/MAZoi20pmfs1+l7j6aXj2DHXhWd9vmwrtGesfzTbWR4GH9UQkJgoAVSn
YT2kcuLevxB7k6jMvk812cOFLAPZxoWqbkjBSqolez2tIKcTPbxHNXHbIX3vpk51B6TXNVGHzV0k
6v+WVza3U4A780RtEvKRgUe+6RYkfLrIksQNxYjntycN4wz/8WOB3H7WTFvxj2Eu3suxeohEDxUG
76JGGOfdod7H8bbHYFg5Gch8XrnuYXVOpSqmP3amTIL9YbQtPyyMUCezyzJDTcHGydW8JmQgXR8f
C1nxxYURUbHiEA7xDyeGz8rUFGvXSI4Zpeg+Fj6x74qgCBQ35eZ7adFY/91+SDw6frT5VOu2tGd7
R5SZtKEZPw/OrgWOliqo5v5pG9JaJQSKAybwSxfDZ1Yz/rEtVRXapW0Mf+eznuTLprfFU9HTF96B
ONjmJxINKyk0CAqqRuWAz5sA0UKMBdS+2hIKyI5MbWv0fet881Kd/JD9lzVw3efAMAE/h6HxLv/U
ncVsISKeFBfx90yvhiOiGYAi4hdiVlDctKXtg2J57LOKV6T/mCiKT++m4dVb8WnsOsjCmyLG6QJR
Vk7iFpx7dKoLHBeH+0sO8/pyRg+Nc3G6iOGodFBSqVGrYPro0xAXraQN/CPyFeRMBX4YVK3XlV+a
AJCpBYNM6epAzN6OAsnRM+lvaqNPFaC+3Z8Qiji2ZY5Jfpn0+h2ThpmtB8DmUChqOXplzu8QcEvm
ysK4gf5mZ7E3oEjBLf8NGczY+X7tzUP7mtaE0ZY4uJ2GP4E1mWQ33R5gW4ru3Iv0z/dLNLd/uVB7
+WuMXdOAu7br5xvwJoOIgKL1Nkl/QumOsreRNG3Na1F4vDrv4dsEZ8hGejywqc8Sg5DzDf5ysvzb
WLOdg6mrgxKFBEq96q8M431OvIhC+1SAUx3zM/8J09FG/Z4Wk0VyzDKxjMAxaCO8thfWlYBMerQv
xGkncKgB6LXB7+kp2p3BPEB09LVL7y4n2yQQlOGzFwCZ4tKPy5ioXdAbNCcZf16UBUzUgGVccm+J
8qGSQZmwEwSLT4+x5KH1oNjaxWfapxuzHTINa7GYO4Q5NqjCRcQoRI9hXzYsOlyhD+jkv1+duKR9
6KksBdaLUIamDwcvLyIPuQjRG++ZyPGRYzZRpV/QSBtg/tsknfbcINo7I3MYWh41B34T8JZ5TVZy
eBxYi5H6GgpL8b4szerH29lldW+G1F2ZqmlnAykNbVV5V7CSITPJ+dm1IkQh0mMcrMWhJC3qaHO5
42QYrlv9IGkYRvRaRoSSE43oNT7qjMt7+bKGUxzxdDrP/s21A4TqwcoNuGA6lJbGNpWot3J6AtWp
0+nENXr/j91l++hLp3L8M22P/W07oCB+0+vYqppWUXcqnT1dMd0ij8mBsEUfBB+bkiXYrmax20ja
DNGFE9jqS7J2qvhNBD8R1EWuTcotbjBoXmLPoddic1GaOYta49wS4SXXEjt0Gy6yn6tSNvuof2Ka
FFyqL24XvCULf+FXACmWb/b/xNiDD4jlJ89CGC3s2pKaW3A5uZ5qICJ3egJlNQmMWY22lj4CLa3x
VcC2/unscnYF7Bl9AaDCMvqWP0/hN9NzLumUfbMnYUG0FpHyXLq9di5bVWg38yH8ibxzinj1Nr6D
t6yGKo0Dg4kVrXa3GabrvzufyAt0aWwi5wHoDq/5SoA1mh6F1D4cAFJsBRLsYbl6t8V699K5I9GH
JqN7El0ci6Slp9xEBbJgFdO3E/bv+rHqJ4SrxFejUC3/se/sMRsm1khcFBAvVjDL2MlMXE4OQwF9
qCOSPKYA30dNOuLcXc+FqyXdJ2rsmr9DL3mVSsLSvzYaNLv7hlOpDNYLe2yvjJnhArGwDV3O5Whp
bthkogdM9G40V9mKpqy2Mi+Wesv1uP4LhwRD5tHQ2IdLK2W8Y5CHk8aL7H7eO2k48Q+cl7H9kA7c
YHn+/tGlVeTiDobhAdmjf7ihkUIrg5dShZaRLbRfREYUCMi9zdsjHsd9gErohese3zqs9dtCZf69
en7FZ8iKPFM+QNrRXMR30yiQu09DDj2OYzKpU3/O6uVCXtNxH+WzJ71jhApvGzR5hOtAaJH+ehx5
0ZuE/ye1b/rQNsR0gGXlqA+wKN+T6QAF4Zy7MwVNmf5M1lKOXdLfHv5mlxfnZMdAuJ9mf0ym981t
IGBtMV9D27tRpxv2RhA5rKAY0q8lUpye4CtRDIyIT+L2RGO5JUprYlPa6vg8XEzvjkH4z6UW1C9X
xmyI23HpA/VXSOjq+r/qFcb2f65jRW+lmOKUYstgdWl/z+toJEtnzjHRL+/0mvCgNfYdQHYsehVi
Rn4AvsbBQoDqZ7X+piPey1KEsxZu/OnLDscrdgpGofN9Kxnse4VldvhVof1uLD/t5UpnCxOaSp0p
PPITao995bsk60W2h+OVOfkEh1vuAiTBneYQdkYyyqhh6CkDr/Gx/GqWVl0Brr29TKwLYa4UVNzt
Sba0Nz07BBMkE2Z/IqQ9/vDK7cZjWZLxn3eJe/5JcIi8FdytAY+sMPZk/w9pfd2Hktr6yBLWUAxi
1F+LzmTMsP4ZLLFJ6bmypKQQwkHB8p018MarK9W5kuqIjHAQ+lVvEXghm7hwR07WfAaBgaxTGJLp
05sjQlbiDOcm7gUhQgkhJgl9G6CCKYR/aqr8C+bgAX9q5uviBD/UcoF31Io+iXNjf/e+HZp8UlX+
3Aq3WQ/qbiHwZ+fh5kfPFnRPz9GAiN6uO3xZ/fZXHFbVENPGFQmaUvbZD2VMbKM/uAIGIuMQ6Jda
0rEVp7wrjUqvQsLpaCTycQyWeA8eEh7855Ftyq29kCW1Ztqw6/fR44HC35dYenwRws9zGgC4Kmiy
PynrZl8TEP9wrc1NWI3IG/ejDVx1SyqaedLQ8/i7DgcPJtMfPIRSfdHZlGZ6Gg0XEz6X0pz+eFwh
vZnwYcz7VEd4fF1o50Gf3def27PvWeOHDUlDHQQfQUDGqNWsKmuiTF1gUltjGgwPl2WS0qtfzyTL
pVKTV+ik42ACCZnEVXoSbjQhnHvMnKp759NW45FhuH5PYlqQF5WRQ2gxi0kOX9wkyURRL4qOoyq7
5VNpkatsZ4GZnlJtpoPCcIa7Fu7TBPIVYqil5sosaXyqQnwP0VIu3rEuzQxYMV12Fd0NreRnCDSg
TPXJO7zfefSwGaBjMGnlnqa2ljQPpQRWnGajw9d+d92AmTLDfbsG8oYn1HwTjbRLHLkf4Yg0WROE
c8e5GZynifSe1bFJwb/T3/KvXS7Cj9XWIIrcESH8TfUijueNrm1P/wyVJDsITbrCbgwFGJQ2oj6y
xUJ4TXs2JKVYHjbK+sKYEBerY+w8i/8QkqwDDDjhxkMgMikHPy0j9k6lEovjV93VXxeIpszgXJo0
fIszspYpLlXko/YNQrk6rKfv26Pg8Y82FGIKQHVHEJglOYAEuKWbjL9TVIRWVokbKnNySa9f2p18
AJVchEDFxiw6/VCSwSCfmiKKljxWP4rUTiIe4REk478kYEdM7fiawkyFm/LpsBeL1GV0Jr0SGxTu
PM9as/n7CwSHbiGDRqO+FwWSZttSzA3ijfnv5wjF8km2yv0y8kjGKqDR4xiDhtMw4JUIWMALRKzk
XJ0PfMEqniuSiPmETB8BgExfQ7leQAdcGWZJkUG30+qfYgtOhKdtEgTZwIHAtO2sbjIZHbh9La19
U97U/D9XpOuvImiEBzXaX9RkfJqS8Y1Y731sjmOlNXIeitDQSwajJbs+b816ujb//8XOwgSs1Gem
st5x/w8CyUQCHBmJvNOKB+a6sHmXmlZRozocJ2ffQjttFfcs1v2X8iMObj+5kFgRvy7UAsnPmo3/
nOmP4EetXF+TuaYAhpiZ4Z5dpCL+ZZNOaznfIR+I9ru9EM81NFFz0GMiVMKDoxmaDQM5WSmtLV0X
QFPvgeM7B5TtoGVa0nOMOMYVM5Q+Qug1wYgNR78rR4CLgU34fZc2sWxWcFWs3sy9jk1XdDP96f9m
Xg8SF8gWeOTkAESDRaITnC9YZmQI0l4yJHZw2XYsLWYtKZkOLF+XCbErVApDXh+3Lt/MYf0OFcQj
DzkuQ5QLZO0do3fVAzsonnhHWYVs+7SdmninQvRDgn4VtiAOOP42/jF+R2HuG8Mq7Cj3JN3XGJr+
xa/f3zGxMU0qcFkNk70HX7mAdzebN4kTaOQR04s/D1RKwMIBv8Mthnsd4aNZTX84QAeJGuw6yh1H
VUlEEsbZ3xdjS6WbaDZYHUJG+KvQD4Z5khDdRd2YvCreOJRD/00HKTBnavuL3SRlwPurYmuNpAoW
s7aFCAWXMvbMpzFNddZsovzy95gaxH9roqQkCk4MoRlIgWQVjoMaMEhXmpKvy7nO6NPNJDmBqbig
gt0IY6rzTupvSVl7PcTe8+aeO14KpBXU5Wd4hL7hg59DtOhDUIgsCdczQdlchAibhnOPQCjwza9H
86goCxkTTcsKAPy1XXc2sItjrK7GrROWZ+ALbpji1oX3pWwMyfHLUb5v9nY8FwN4pvCHJVTmqui0
vYN2+DvSyBBnbncVVXtaXiwVCna7N92cERdTqnt2UjpkBK97sCsDe5tE/qQTezw/ZSPOPXy0GCNh
v63YL6lKtIWdtrkyRahdJFowOuTxPvhxbN1Tgtbx7jyUo+aSyMdoXUGwfkZQth84LmfJ0XzFVcoe
UW89cnm6Z3hOYKwr5ea0Y45//F5V3kCZU0E62HMDDWJI0u8dZrBhB/LpoeZCBkKcFsP+3SC4ckyl
bQ5RTryXCS5jq/JAteFV22R0s2x1twVDb6HRXTU19nZrnwwz3/Rp4g6XKula9KkcisWizdBuoy0m
vcszjeq3E1JTihyfu1JFpA8mvl6S7vFqfViOABNs27tTmZD2sqjcaOtfzewoK6ZlKJtkElwq/tCA
GWgGDcHIypqpk8ykPQU4+YUgOd5DFf0mLz6lKz6MU3PlzxXFJnJ000peF/Fg+PlV2wZ6hSbEB4J0
I2j/2owdIiuax5IGp0Q6gavxbjxJQu/dlRbBd4UWN1keOY93tvY65/dedhNh//e8DpSKhJ6EE4Be
dt978pXLNdYO4RC+f3lL/gzFeDUUN1m5/mxPhFgsjriiVZe34nI91TtH4kfxx+DWqqSh1D3ZaV6H
gPivR8sbE5e/BhJ8wvEtBOucr+uRgA+wQ/3k7JuKy7ht6ICRls2Prd9GjHnMcdNLlmnTBS9BRRlK
aDpzRVVScmTtoLw9XCPG13OQk5H3H+t4bHJLioEc9bFceNBVi7VTVXAMCgjZW66+6FOfT/nADfPN
816x9XM97KrOu5BOd+zH6Tf2pmKKVwx+9wD5rVgrJObfeJe8wDE/eo0OMDLp7N35OKg+pnRn3B1h
Mj52orju19yMBbwvf7rLZoKmvuF4iWPHg5M0pvSa7Vfa34gyiljmcp/g9buY9BKyG5rdYfyVV4pR
7Izvh++Et5hyBoTgenLSMUfSEEOJkWR6Zt2iMo3Oj/ZSvp/ueZKinvuAPFT0h/kwAEkz3RTLiFje
9e+YP7Ng2qKU/biRLqjgWM58eAZMVM1U97fP4aW7C2T0N2Z6VvXUBSHVKB2R75o/a54ol9RgwTzo
n33Fs5eKdVQiXfKu90W8GGBlC0oCFgTZoxpGiOKuEaE0WVBMd1XuS/7mjGopz3e8wxvOGssALrj+
C6nlKsRgVoSjH92BwlWbIAUIsKwca3bqNPj7Zd5VA+c3jN/vbfNVFqkuXNNDVMCPz/mGPaOVBust
W2fPpIz4+fVTGxXOagzqIIGKVfrygk7hOiINtfzyS3mmcIopdE8/uSQ/5cXGbCd8LbYxMG/T0ZKk
Ch3SO7eoUQc3+9pEjzZxdkcUmDA2qEUWut6sY1v7KVi8HfYN3SpV0fi+WnRoy35+pfeGT7z0L5yH
AIEyZfs/a61x4AiN0QiCVBCF8yfmwSa9NrlkKLX450ANvcxdrTF1O/NGTM7jeTRmVBXMXF9c7J/W
RuA8A4pDp8dDNee1/epgQht9T/mr+W7v3MAzSQHRfGeJxzcg+SWkv11qHLQMxFeg6NGQkyEAFVs4
3fxjwg6PhMf9gXw1LCYByn972cDe85kJh2lsfn2a35B0RSy/gn9ReIe7wSb7ULyoOACp/XvsQwGu
tyZ6xfkamrYIwohf3vpAd+/bGKQqAXV4FU3NEvRaHw9JayoMyWLciKbUetIhog3LFNqQ7h4y9dUM
W614vt9UOA2uZRMQQCOEHHRwtaCpzmlyo0okcWJdgR9drnIj+ZI9w+cFU7ost/FM33g6+zwBJcd3
+gzVoJcC9xOYfMwthdnpmptP8/KBOqMcN4gWidksgDAqF2ubv0ZFlUnvxdEbQL6WqgYIMQjW5Mbo
NNjOIgMR9CCQ/eVDN8cvOxJRLBTJY7f0SP72J+PFW+bJdn8Ra4cT33Q0XAdayjbbhJbC2DASgCMe
E8IYe+UoERTynJaCg40xGRMy1q0mXl8va/kxphEITt8s355uZ063BwINStbRZrZJQuu3MHdXDdvU
5R88uCB1c0p7Y9bfcCUeOSuOHMvIug7GancC7PS97Wyef1+DfBFdkJmPhK+s9xuqCQjb8tm15FeD
pH3KFdpcajQPyhl6LJRUEkvgKOGa/DAj8JvYpCYOS09z5EPNcr24g02Z39nPd9sR/HjEoLeRQ9tl
Kf8RfnYP8kCoZH7E6Bx0oBe8KHFaL4XXURhxt832hPIThilA6qG4Acrk2MOGdYl0MRxd6xMAfLEK
LLAsdUAe3seR/pepv1FX5goe7wPjvl94vM+6X2xskPZLUuW/NuN5s1K4whVPzWMoU42zV+pPsFNL
Bc3G0DiKsPsy5LOyALLYxHgvaSQ69ldTzWh1x+ojPPq5Hcd77SCkHOrfwR2jQTTwvXBLpGkpI9VM
4n7Fhfogg66XBU0D3r8QHp6AJ9F9yCYZ5xm/OnlZ9I2npG6Ul0MuTcSgVqbmmCZros9pV9679HOF
afS0Js80kr9y0hdgbXymUkIBAp/+7KxUIe0+sz41RGjxX2J/FuL7O4GL9Nm3DEkMz0VnbTVcez6B
/vOPW7rrjHJuvPXdDM1mA9MRVS2tnTE9wm1NtuzeztBuDgHJlp4+g5+EEARV+bojiuWOC6ADa3GX
u6xdPYS34FeUvzicGf9n2YOq3wTaDmoVaEvgfQvpM5eTyJtwM1nO2QjcQPfY0YkKd1oWLwwCKrJk
iMvtNFkf8YwtywE8ri7GOH12cS9lRu6fMFo3vFJzeQil8xwml1X5qsclGmZKyKChQMi4/VihGOrb
IJzC77QoKohpyBlPv2hYvt+DMNWjsSoyiYrQgTaxDAACaPpwvRzncbWJ/xTAeJYv8V9kAiGFE/Pd
590TZf/oPajpPRZZNTwFEhxpFGmutiH2bUbsOsw51LvpRU4dCm2nmtpMCEi70UeXC3qWuW4YgmEb
lVz0nT2fFYCtVQINUTgYkelq3Y7lC09nfP9mkLTYMNInkkzvqlWJQS8tmyAu6F2WtMesd6CRzoH8
DOJDj4U6LLYz7ctmQ/Ht87rzszJmuBpv7YdDISyqkFVhtI9ekP/ADcLJaZT5Z4KZQR5FWrUNFw87
M0HfbT13wUcei0fBgrh7CDBSTFrZUlipLdG+teEjO4Gtf45TiZ7u7RMKRnlqrEADWug4UhSUaV81
5MpeQYZ9MgLdYkegBmLnZKCJBfinjO35ss4b3+krvoyovP5hWKu3jGTVFdEmPKYC/f95QPH49eUt
mdT8xLCyM9UPzvjpoYOdKHTWzGywHGSh28+mqywjyLnN/lL39Q4arqOuCbe5njCLHPusT/uxkF/6
WCH3txW6NE+ibNUrzIHtgOplW7ryhw1kxlmSUlWn2IQ7pktOkHGoaNpuNKEYKlogdPANYkW//qih
yiJwVBTYu+WIzOXOyhcesq4Htn0vFrutLLn1Mp3AhfZEwlTmlmKpVTi+U6IAZ2GNeDXBVABNaAYO
9ZuR5xCKgW74i3pRBewOtknqTTjKTM8bJuHCGceMMz71nshal3QK3p64j4Xq/PE2NwdH2vBA9ITW
O0JFavzUAMNrYphRc4tC2TglAvAoFwO76l5gp+OE3xvPxsoD5nUlDHOwmlLGP/szunWCFahnysEl
ilgTsM15c63CHfaIKVxp9QzsclsaW0Bve+0XieBaxcq7c15wrZ7TA1hvawWoyOQf/d0onm/RH/74
8dz0lZek/1MU2e8tPHLK0BX55U8N1Oe4QvJ5VVblUvaWuol3GOsjYtrUBcadO0dX6tBzVZeN/Mrl
uDTBTrh1giGj1pwCEUzeo7uHsBh8KBu4MCMSL9xWjxVFFjf6VOb8iTaHFJeNronkrxSC/k3hlvvK
PLFb9Ts4FN2mYPDwaVjzSlk0zOxdszO87W8cSOGVnzwzaTe5jFBFJK6M913iz9bqnl6QB8RiCSQ0
7RjOVV0YlFRRdLH+HmX6C2IITLla19YSayIU00t216Q/wf//hSedZMBIfbh30a2rgyfbqpWgfteN
H5PBAhSeC+KkpuUKmREPFhtUwwQ+PYLvZfSliO3gyi++iQJKaZPJSLeebT3MezqPckvm59MVs+xG
iatbmPFP0YOAKhLYDu6V7tHT89z0bTyxVs8o4AARuaxMoN5PmmP/AnlKpMrGUkpAAdSBYvHxHcGF
PKt1fJBDIP4NKgXaF3/3UrPHZc1yBtRv7xHEzBdPTvEcGfD1yuNY8qh31ba76lP7Al8N2DAhqduD
vnPxYbFNOBFJ0vzHdrG7qGIMrDr5QC+ALXaZl+PL0/Ox9Nt8OYASW8j2clXiR9lS5hx+SY9b4XH2
UmGGqX728vnQ9MeN33D2uvAHiFeWwLTGZde6fUuDQybx79tsjlvZKOQCi9m6/EpEJjEoYIQwKIGw
7lk/PzwmtgbVGvHy6Gdf9Qu843HWgUE5JgV7feneKX6C75VGB3ScwK+rzjxVQaHTfNity6HlAAKV
dFZ/5eqlMYFqLpBM1/PzTjot0aRyBCalf8qdOkShT4I3Mv/wmh/U9nveOJhjSymqpT8YFT9oMKar
wN9BOnQvv2hpvtqIdvXWS1OcEckyD8OPNPqkI76ImZH6Nw8PrODFTjAIgMDTY67cICKwzVGvXFX1
YC6u/ji0fJ1SqHpt7VKJzpDz7UyihFTHDdK3hDLfWDFRdKizki+xi3mDYn9xlstgIC4lWAV1793m
1jvy+7xp1+ke/DiMEB4d7HjirRa6qQtpt/GznCsMQNFSWA+gqxV3zXw7AGd9x3yVYnOy/rISPABN
UVfV1/xUtr8fbd5oZWWzQmIiqPde5DSx9kXnx4rcYZQTHoYwY9qnLfILW1PxzzV2kv1CT+dA6JNy
xQiwcIznkgzimtPkInyd8qxyW6LRn2m0RfUrqkrzJemNwTDR8ZvzmoPO1Var6jMddU0TlITRaNr2
j9pK32lxhkOpXuRiNesrcRgs+WO+5mmIw2yrIKUoRr3ecjGPf6sBpkB0Ykr8ZRzyhVKCQulYEcpz
Lzif7q2QC/m369YSaonod7qSO3j3hoGTDlD2osjEP2DTTuaKNKAPsX4kNWTT/2qZwMaQFRksXpBj
fhBdkh8zpK35th7UGX4oVuCManGtDkJ6ou3xbcTVK2eWz8UERgahJALZiXrYg63DjypUOfMXBNR3
FOa3WZ5tHwBr7nT8QoNnvtt+iZLyyv7kHRzbLhH52qWhGLQIIxiHSz8+G5zpRZj6PoukURSXLEVU
Dn+xfkGcOvS+8oV+n2WhwXJ97fa1YeHE5cWDO4M+9y2+FNYlvq7IHDBOq8+YSinzV1SOFz9w2MjP
69qHbEMAaAODNixeXpw5+QHrLFLM0LV3Jq10yJzDxsuuAXv0yYRB4t+ATVyt9+2lTVUIs1S5ypzL
MethLfD1WEP2BejBbeW3zimze0sp8MydAMmPxeOH95Dpwz34B7XJgQ4QTP99Ht5YtNhAsvHzjNZl
lSID3AON/h3jIhu5iZfBDRaoWHiigq76uag8phm3G3HIfH2iEaTno64GXqcmGSGm71h1gfXnGqYK
gp50UmSiNqLJhBK/EXtWersfwgrXJaj+Oeeo3V97uigcYb27bigHhEKpjWtuYPsppQg9OSDXkPRB
m8DneoRMgZcs0d5lsnLiAMyvvqU83RpqnG8SVsd8FaPtJsv8a+t+19Sq8qpBo6y/r9/B+LWn/WJ4
BgVja4XaBMqYx6+ZxRcBfaboyPegU3ULCNuCQkkt04KpXAqDSe3pjajA2to/lohdWDUFqEam5LuT
raKo2VBCw2Yhl/S4LC0z1PLSW7yq6+pcAxP/U2ev7dnMqj5UOrjb6P8AsdDc8zNcCEHNdhpW0XC9
vfxMUWZ/6JbnxPceR7hHlaizlkFV1kgKzEJKtC/2MgNwGJ6wkqHbFzLEXjuUt8/2JBcGGcA+kgo+
iZPWr9iCxyDpD7GDen0ZMlvJEBsWZOvRnN9Lb5LhCzd6LNKea8nyd96ftZD64TGr161EEN621t35
7hd+m8fMYz2boDfbhFHSVgMIGRhuiqSEBtee4/aEiNW9yskrdVHdEeCOfFhXs8rqxG4WLBQU58r5
isfOXuqC0xVTUQ6dBBpiI3Q3cxNA8rQrZbQDTlnZMOv/NRoagWIZ3pAEOeFn3N7KQnoAf4LxeEGs
vw1+bfriBUiodTYHsjoiV+INj+f5CfTbY6zSBKQD6meSTN+7q+rzAl1b+pXMUgFQgcoYihWJEKbr
dRlQ89BscHp+uQRAzUGQSjiNs/W2Y5ns8dy3bned5HotsFNN3GGe3BcRziUXrU2063PJQ1X60iLr
XziFJPyg9zaGWrTYNVSS70c0cYJNSBb0sKp+Rg0S4zLImrEvFlNN4biknyDtFSKfP9fm85mnPdUa
m1Gdg0RGG1UaKOa2cxd/cgFwUmIUOsa8tYQJSd+1rlzgkPeGg1Px5Srzb32Aq61QgzRfNkbZ9OnR
PYD3sQ2t9jruKQjDejwU/4p+G66JvyIwdw0F/BNOCp4ZGE2mq4vplOtIXfuLhDBu5GVD9LxeVKhq
9Wx6sn7VRhV8poxy+MuejZsC3D95fSEPP4+6ACi0RHidPwvLuXoRIIiFUIZc4e0H7+sPm+hVuhxD
PwscCVJE1XeW3dz5txuixmFbSP6wy3bE5vjzYbG9wBG0zMNKwk4m/YIOZgOizc/vqGTMAREvQ0au
lHezk+axWrBT15n21/XkXINAWEW9+o3789YmmDEav59N7U7mmFFgyoO+OseDVuA6cDxNrTT8YzQN
AbtJww9J0Qf0iz7DFpqbVy7kvh2+aH9iYW3jJm6s57U5hQWUBt5UXCjVz6GV9O+o5sEgmAO7mAkR
vwg0wuPb0c3kLb9YTLaqqQclEDPQktzW8af8sO5PJrlefmXO92APpMbrNq3crr67k/q1tXKSwECt
181qTYeTuB0x11/PbmI0ShJ47GtJxVf4LLP9tQDQFAy7uftnFPuZYd+M00bGPdeUycxvbBlvyj59
i3tUcFm+egYFIf82ajGIY1FpeI+0Mn/7u6il08zJXqexWRLo0LBVjBy5jbspYZdHdo6R/1x0X4RJ
VWcOshrd69XZLaWCjbVdFIEXtNDWy5E7rj4M4HYzL6Fz6QDySSdg65mietvpUdSlpetOAbap5sYi
BUC/SHz7ojXOJhzkwR1J4HuElBPGkIRTryQ3W8t6D1sEr+AFs8sPwZVvbegX+27uKip8GT6Gf+Vk
yvtVBWaQjg3/xHDc33m00IVMSIcRU5mLTAr08QndVsmJWlZgPkifthwa8/o4ebFLJ4Jem7QWGmyC
rh3pkGp5+1YkSEJqV8qkJw27VSg+S5TZO9xy7eYxM8ahwRg3wBBlckBz6d+ANteM+Nv8Rx6SrL38
DwvwJJcq9Sb9/Dy3azl8uLHGsNSFPa7jLfwWnF/r9YqW0eh6Cjq0ac56HpACMeG6TKPDe7Kn9dw6
49TP6cmdVvzf9Bhh8bcHCND+hnMDwVzZJKFEcRpOeq16IIUS4OqIr/mPDMfjh9g6VsWpvQmxTEdY
9zEm6nU1c69z7BaBfHB7CBJC9kgv14pbQ8ZIPj2bDVqNZEWjxdKZ0LF4WCd0TRNYq3JotTvRsXUI
NL7gJYjJInoXNs804kYFiRkjLBgdUAqPLz+GxyXgBTSKFE7ZF8DwdJ1Lixv3c0ruWK+l3A1bHZKW
q3rQWHc7woG8CbVrZLti0dkRWJuNGyCJ1AZt7riHTqYutB/UYxRXRMtsrieTEGlqQOKFN6+44ONW
ZJYYAycAum8Nu35sk3YeGxx1ZrpigOuxDDm+FuTTxL+zqCdEr1L9Ito+ATiH2Pbs9Ko66Exz3j02
DoDC2xxLSa5S0ClE78vfWCUw7juLyBDmnRBNHFzAY3zX5csLbMOGnL10iKU4U6gLrvuUiEfv5CK3
TvkqpqXTCmzwKxAczibahlg+sZozWGeTX1EnA4hGWglvVGSfmcktfmiUSParrpIDe2MfPilEyUR7
XfbdjFWbqLO5cR0MlY/6KUEkm21C70xNQ8SWi74YKsc35Q8rhbOC3QSREIDXoALi3gHlqjoVa6XX
tNduOtxNzGgVvhWyRZiXMvBoX932dGMzI278p4Wl+r6GZWZYWYTB49FIS37Uf6UebJOKywlmK44U
u9X3P6QzlxjkLYF+2adsNtRzfCneJQ5Y2/pFoLbBSbYmpu0KlxcrNjPTWRsiKhEFbQ9yAz5dPBMw
pt/Pvz5T+r5/0CkO8xFSl/uTHflwS/aE7xxT+KQME+kGFHbCn3lcA26vmiy0ASPcTZ+40IIuKdqH
22ddfqUJ5hvmcPQrZo/L4iy3gIGVEPhTLUDXQVtMTTfOv8cgvBvy9bqH3v9FrIiifnoPY7j/CxK2
Gy0gz3MVHpqP+nB5nLhrjGI1nMBz13J/kGChJCMlUGsmAmZMnGARb8qc9opi448OzArHEpPNvXP0
ZZR5KXyLAqNHkqToxlCjw+eZzsEz0Tew7SlALY8VR+iNnZxsqzA1bpvGkxfx8Gt84utNXxwtSWcm
X3BSdithfvQAl9bK3X3x7plCbelaP2PbiljDxf8KikCIJr3cdVufSiHa3uR8FooPGIYhl91TyNgS
tgqPKWEZMBXsADQ3QG+6/A1gkirGqF14UAFpcnIuxSp9+d9y/sYPfTLiXEsPIGOwu3beA59uAVc+
EPKpGAftMN7XsQqjOliKo7EjxtSP1nRkTg9S2TzMMt9mFZc6W5dLAB6cXELPyPgZw38MHnv6Gi07
T/uzuWT+YSnOWTXeNESya93tCKgrKlFePhWx8+fvWktZBpbr7/mfqdupCAicG8zcxISL/99cJc++
NRp1J+x0ArFc1EttapXthE0WTGkL1W51Lu4HvYJU0Efymf56W7VXhYWt2+tsMUrftTYjAaIbwte3
mBA8n39NpUJ6xf7rvrWWLLi7DkuqSeqSzvyCbs6DleQlBXhG277D6ofU2V9IzdmFZzThNxkU5DrR
ZWSBKnXgUE7pMImodmNlpJdkmIIcEMdFd7x3BvNfJIma01Anedtb9dvmnJtIpHFhsO2z0RAH/+DS
KlfdWqGhosD6Oc96/rbVTJYglB77nwj1d0k/XAEJW+vbpHinItIAQpl7iGd3TM/ZryWm/dtKu+D7
x+wCkLZtFTUaDJ1PwuUB4f9lRpoYbGiR2cPeek7KDh5h/3l43Qo4bKhTAX+fvAPiYpvgpuwF+Hka
e53SQlxpho2WnfHrZt95JsnB8dMWLVOVrYWkQ0GJRv6dyO1Jk9hm/T5lmXrdKvn9ZdZ3klt1fP7q
BFhshvxr/FpZkkouVnA2/7PNmzQ3QhA1FlaR1Z1zeanZdBQT5ttl8ptaGm8uey8EBHrKxkurQigk
tFEn0FV+RYG8Vs69P4RVzYebfGYSjryswXgQkuXIwX3bB5ujapuzLzrDry9xaBEUAViVrOM23KsV
C70RdWaLhIhjDxDm5jkDFTqht121W/hxStvjtf2UVym0RI/PGgynfO5dvP5mJJNcnSOrKgYgcFze
FHGN1ykRTJ+lsNj9DP2PzNQTgaHiDPi6CbTXpeDSWhtci5u2N/jWwlpIp71XE8IpHHwsyAa/KMhj
hTgvNhTqzFhpZGd6FtS/gQZlSRnJDWZ+Asi5aHpbBtNw22rlQ+OG7UZP7vfSoDcqonA2Rdjb87lU
NBrmENZ+wwZgdWzet7lMpL5Vbls9khFRsti7sHy7qAz0/jYcnbjwG8+6vsLRd8bFzYiwFzuzUSLQ
spFeB06jd4S5E2BCeGpOyW4h4UC7k/nG4XwcWkfBIm5+fLlkqwunMfQskLJASjtzHbd7D/MIMGT7
1QtWyMQW4lOYOCROtgRxXqtVErJOJKpoODSyFp2aGIB0IfR/V9JrZNYLcOaMf9XFS0+HjtZUf0+F
YQHemo1uNmwPU6kJ+MByf4G6E+Pf7jPFMv1/zvfIWsFULrHgVzMWWM1WJn9Bu43+oZfZw066r76X
7/z3BAXzMfnz26EaFYBG27wuiJBFiLN+nISwy7IOHotDeZP0HPyj5CEdCh2SCUyHFk8b77GswBH1
GT19U9ycNql4U7Y08SNlmQKbrl37We4zOQGBa7a/6hCjdGL/AmM9VDlAifPPn7PSYlw6ry4ixaW0
I30HfHE8EfSsBqOpDNLNdUnJvVPmPevUlE4ZPkQmU6oxl0nF2MArg0WRZmsWanxtpXRPFr99gRLD
1f0IvaHWRUq550HSaLm7fIZ6M11DqQAWmN8Ze3zpIGB29H3OY0ahANUjqrDnMgxBGcAeYoq8oGIP
J+BvFwj9e0fZOqQ/QtcfOw5yTlEtxvrPq+paVs7Mg66/r7x5apheDpBeJyewgf0YXKEHLeUWLQ15
bdw+hoJ4aSt0Qe00jO205VVXl+FTf1JeRpxGEE/DhCsLmhR0wQHiVmKu+W7QHq9ikxLcJBhpavFX
yTWnjg+3b67ImZKTCtDszjYquveSmbqdx18K6bCVW+Uy+eQBE5liGf6ZXVMh6bBdvRgyjlAodCid
ZfkfqErxZQgRAsYFjIh/uC/p1WvCoGcN/aB5NNk2ESFPLcrsfaJKUuuw2nOHnty/KaLxpt8tE207
LDUZSlQfm3NjMSdbB8/+wLjsrmXsQcB0sxElSQ4b2qef+LImIWyt/gOTSfaQPMF3NKbhTWl9MHlH
LtkKpnG/ergRtWROEwEsgwBZNt09mnBIANxtJErcreiJe2a4iGOCRJbJl3rKo4QRt7LAnliSBZsJ
LfHyt4t+pUIvemMJtQdr0R7RLp3R/YqLjR9Ks7LZdN1GTYRwxISSHiRio0bgUCkLZcyjSPCbSNw7
32pAoSru+pwFsPIMZWSCuVHkfn1kWbfBmOycXEkbKST8vyam8ZJCDl5DoBpNLSsyu/wpA4JNkxJP
roseXJ1mSKcVALyZOn35AyZLTn/VVW1gIc84CsjaZ2OzFrcGKauwlu4v05IahdZ4RxmXNcDz3wUH
5JBXVbr8XRCetxvUjLa9O4uDHjvLm/WZ/0cI7b491NUKIlFCevbZnMKesjWcKfCztQZrInrvBVRK
gjUwfi6GstcDtOOpscZT3aIgr4dgm1XNXLenH0UGaYxlIzyZbHAimGbd3ykBD7zbuWza0lYltibQ
adCU26GpZ6ZIFcVQl5bFZfiz0ri/Bdrjt3l2yQT4vjPEOMEtw4vO1XR6/jQqcN/Ka5BF7A3GxJRW
iz2zCL6X9d3shggReWPvUiYxZ+ec/jwqUe/EJn4ytrRLRDRxrwzJFJHB0fPjYsTmRRmH2kFL407c
cubz7Ls+0nh81br/BrY7HOz/l0Lx+PqSagTA2dzJOUhGq9zvizZTRt/B9el8pV0xSC9++Ds/Dd0y
2UAiGOBnaQ72SOjXRnwQC0GIDhA9sp9zTQiPs5sBu/HMpBx4LkMVH+FOKDaPkavGq4WhZiHGhvkK
vorTBMMMQ/Jx5k2ZeiDGip38+QYORkRoQynJhHdtMTI5LbCUj7ZROPGtT9CzzbEN0d5s65fttuFE
unfKElBX1hnFoMb/sOp5kIIg7k58C1xM14JXXzhuRlyXyLUuYnrLoFsDfVPUk+kCv6dAVUAnUoyh
Cf1f4l+EAutiEH/ErRE5aUuhvf3rgK0bzSLofhMQFJv1GaWQAQOc1UIsqzI0+HPJmSSMEptsWdmI
jARDLF49ToZok6aG4fUs11r1Z232fM6T/sZ9Rv78+xhIzLLfSWhcQKhS0xMWKedH/JVdR9eNs56S
uy2wFYC5JS/HgH/mmVJZw5m8In0vyJW5WG1RN3vqJPw4LMqCR3Fvqxibf8RckfUMXvZuBh8/qlch
lMdSWxviwm5QdOaKlZravJzWfx+PkAaFtQJ/NBsX/TRTzRGrLOPJJvWvyubuxEvO5mpk8inmfQBq
LPurfwWP6Z0nmbXg8x5Pc73fRXUnS474l17EWTGSptGn+kUp3DFE/5MBwI9xZUkP5vvRKuldCzXW
faxASsPR4Ih1J7pYiT24iFaY0Yxd/Zr31BQ3JYQ7UxZuMUmk4VspOeEHCADm6yxrdU0ljhlAXsXK
P9YCP1fot1gPaV4vA2eG/XSeKqElQ34YmpLDFLWnx2+uXU7OPqio5iMJ8Fl/x1Coalm3jLhiM5LG
mzW0934Hq8RMqd7y226b/h1X/98VGlYBg6I/Uf9pzpqCRKVvEr/BhibBcPSODqCc2vjEnged3Khc
zxEbNhnYzCN1Hfg4OjY8mURHQdRYkvpHPgqO2zSLqlLw79Ukp6ApB18NFm+ywMMuU0ITsAlAVadU
WgQ+CatSVnj023+UYksaoceitmt6VqcrxPRUr7FWn+8ibFENViJTolg8fTfcWcq4qbN55i4YfaNE
gJRKe+zTISjc0vV3u9tAbOe/OD+vwA5uVLSKGggUjWc/402N6sbZ6XL+AL5i38XbzblYwxbHwFLc
/rcYiOh5xFqVBpnx0JBugFzLq+hUg7Vv2tuTDf5BItX9Hw2tSJdepkqUYHiX4sJg59pBba+WNCnY
DLi+APFF/4s9kWoCaN7s0GZwJLpUZP3Jk94Ixr41GGIi2G3HXsnqTMZ6pYDDynfCafisUllXehRv
h5I4DAlMx3b42cCeYBqlE+htIA9jZFyBdDg+cG9oYzrcOL82Y+YGIC0m7zJKJdh5Dx63vUDYyG5M
C16Sgb72OMEKmLL0Tm0Zzb0cLvraY0uGaIGjGH2sT0tpen8/GdZMlakXwB99x+FVs5eEb37lt2gK
nxJlljBAH7Y0GlFP02qvChi3Pw16dgsGF80EzXNxO0/BPmAND3m308pp+ZaAScoG2SNmJjetL4HI
2II9FRxEU58S0o4/2izzbVnPKoR97HrbC/8+P/pWL8bvC1ud0BqXfu/X5gQv06e7PypHTP+vF99n
oQ8LOEjtD8EJ3y0seMnczwGqbOXXB1IeFoJgd49hHpM1PWr9WX6NMYkJ/PmiQUXFmlXdhCVDqyVe
DfLHm3vfSqPSumPvVdSx9nK/FCyOlWGjEucBKSoC0XHYvKivAd558yTMC9gIg2dFIK5FhoWXvUGb
2XHInGJk+E/90/JyVVCbeIYgKtHnMiMEw1lcDI0SBU4DMyxMwKm+J9I/Knmbvd28ltcnlFoHZLWY
A5LKtKIQBo+JIwEqzPFkQRLkjnwlxa9a8SNYMmvpXUxDErFMSSt6XWErZMJP0x5Y3tY4Eyt5J9Fh
L6xlOzc237aa7fW7TupjE+vnyVslnGZob+NONfJUuqBqV+zfMkiJb2Gfo7Z5bpPv0hS5Kn4SUCv6
sfyHDGzQ4S2fcELh4EfO0el56kga0BF/xtCrGsf6nnux4XLl0bBMgvBpQNA8OFr2qa6IefeeT771
81c3ynA+V/9wNhIkKzgkQKmQi/YGithDkem5/1UXOYMsSydEtioHj7UmFVEBu6UN+6fl6BnC9s8Z
9nA+G24Sta4MONmlcIkIfW7WIPXoS76c98PnEs7PAcLWTZHgCn93A7MDzj6QosZjSG+2KLwJp9bp
WKtYYjd2SSAmEdgkPWRXk+jKawA62LhtdSM8EtxZpcpbSU874imnAq48VaxQjn4yBcJr8OZ/4kVs
PENT2FnjrPix+nUZ3JcZ3KMFLLsnxJl8Fvpqs2lphYi2Q0jtRsviWtDwAsvqQXIgzqD9ig1MkHbj
fQcdCGEXDEfd6cvLcmxa8ARDgYgY+G+sttjnbg9kljpHvW2t88TPvudd1UVMpZYdGxszmxVVMSE4
9O1L6hEF3oCeU2SzpNvId5ga33Oe7/rH2JCK9K1uLoTHjJ+OFxWJtRSsal5ltDa4lG7hXBz2I9f7
uS3I8fYRNATSAl/Ns++VRMnOcZKt0w6LS9Nwhhm20SpoIFNeH5A+LeG367YY8Ob+p+cD1JbsIxs1
wOMyOlrKo53qwghuDgYZM2vy9PoNcpqIQUQaHUJs1rxmI4XZlvgyLHKmjcM6oU3N6eXQhcUm1zd6
k/m9AjTVdH7V7GaAhNSCNRE1eB33SsuL42lv4EINyQ2mlvEGNcL+0mJ5BPNOn9z4iYTjDhyfvyvM
JdOc3Z1j3p3CzTFuLPUwHEjnJpCL0rml7nL7rIVw8pNuuFdnDYi1MJ9pvMYLjm7uwk0YRprzLftn
K+WGnqYeUruQK5OcPgkSZOSh9fhYQdUyjf7GSeSpXGBiB07dvF+IuIu4mppwZA9Fa4fEyFyykOB3
q3RM54vf6fVA3SH30AreUU9MyiecM4K2IKOnNNF7TBAaqMB7e1EWZ0tXMftzzH+II6oaJ8EGsRjN
h4K3ToTc7VjJYPDzz+EsV0rub795w5gFw1koVg+bgELd8U+unva0TuewkQZoIkY25hPqUZHmjenH
hbZlFsZDvzvg3ydQVx6GmNrnviMeRyJycWUmj5Cr49p1Pb4Py+ssMXkamsZ3V37ivnX5wUpQwu0/
6hnKQzbFpGXcgf1Kn2l+CGiW/sMGlp2FzIhD7qPsEJgZRj0qEGBY1oe2J7O57pV6KWzSpLMzPQoc
+hIls+yD7fz8qAAOFK7KMAa9QizjH1HToEYyIjBxW2oZHXjvwKRfm9bplJg279TMyZliQTkc/CBQ
1QMXoQeNf5fMjJ4tfDpkoPsD6Fu/IhImhX1wRrMcJt5b6jebc9MPWkruDC9RrbGTxyZerp4sngwC
Y3bCWBOMCIm02ihsaO7VQ2F1bLsadyIgR2b75w9cdq8/VYDFWTddtn9y7DSJcxmKAfZHUi9cQukt
0UOEsWG5kHvx1VHgorSgtUBvCTbmpkTPFT8ZJQNJffgdhDBXu/jBEi4r39CQvdX2q6gWPqdDRdxy
1pC3XedNmGeD6Rd/lgK5Wz30Eo7kAySrGqcqKy+vqhyp4nMKz3oZmDPP3L9ltx59GkvpumplEC1w
+XCPMzfKmWY7BItOieF0offlQrxWtke62nYt139LSCx9Jm85Rv+fSfEZKMfl0Il0rJe2LdsdZr8y
8+7Mbpeo2Am+G1xUekl/RbkwU9WKpSSIPL138MZZPVK2uNTzPrhFQHxP2nUDRFH6P8I272PufCL/
B4J9ds9cTmj2qxpK8UI7RXQ1RAnsqKuKs2FmHDwnSH/5nAIKq5fr465lzGtZvahSc6gnt6xH/Muz
LpMOIOo2VeJfIHRFC8mydGhjiidcyDj9zIz5uQXAOscnYbUI18xqayTLQot9NSn/onK4Wh1F7qvw
arhmF5zwdoZ8Fl3aoY5dlUIcdJbRaN6knm7kWGxpnzXKl2u4uIINYcU9DuLTaeSXlFGISA8oc3q1
uqvJFQ8pgghocQspeLYFmcmYwk3wXkL5TByZ1qRAvZIW4zNoiVREzOOsURU4GLHzuFrkhcWzTa0w
uHPZIabltsFx9446EApZii68p/jpbK7rNT+6Cgr1fuMjpRdVoktL/4dWIz4c+34i1YxH7dVBScv8
vB6DnR5+0Wy8/G5XVw9pTkWYzM9dUmty/Vnm6gwlNPNd4ivnAYVRK3dJvZrSOtPYPqgq/BA1eRmt
bMDVz3/k4fzxG1rV1R2f1y55AuXx8tqeoW08RLIeeo11CLW03oltzpGOwnzU0wNR/GafHvupuIzB
ufBb6zkjmDZ3RcFKGiA33nDxYK15AqopTp12r7+Jhr2H7C6gTx9B1z4uyR10HuGaBcnbHhf9k31l
xCdV/Tlod8E0T4kjYIYHMJzTOLZkrKvrHJyy8oHpER7AQvGWZROlROsj7napsNaqcBF7U4ktH83b
w2H6Fvq6KNCV69URPltIRwQr2lDzFmTfR52hWlFh18zDogynyBxyJqziJjyGPGgOKL115EklRFHV
nnj+cYuvZNr9bHgw8vnLfQJ0rNW4liGyouXfRkGqBQuhVrtZgkTgQNfS4pDA5qrM6KziUjoyIrfw
BggunkzV1eTtoQAmBES+LPbJ3YmVULe52DlWYInUxX/j1WK8DBGg5S42543PX012zsaveUQ32Hsc
2PkPJ2H/wkiw76WD+Q3LFE2yXTazmzMjB+WXi6ciYJO/5xAUcRyIypNmhDTgj96O3xSdEXUviKiT
lCUJ4lI5xohxsoG6lbqgafWuqMM89oKMAxBN0Q0MBIdG76+fov+tjKjipTAGOfvErjy7mjRBnZG5
L/BUgRtgREPDI7tEq+gw3+N7aomGf4eF5Rx2X6SroAdEgECuIjOsTQroo224IhZgkpmwCNb60Bol
Vq1MkfWRi3usp5dsaVDAkM/rALjXLbZGQ4llrL82LoWrzS3tQGc9CLx3+fZYQZB2dqgWBF6dcZeT
PKCH4/gkuC0wD0Pm0bqJei3nFRb08fBxZgFyzbRU9ZGyKH/w0rzCCQkdsa5/WHsqrZcsbi/Axh4a
7CCqIXwkq2gNYCDQ6wnFqjSdIb/VoHewXR//7IpqNqO1JAdFzmAhJi/DqmVZwzfkstzqhMtd4+2y
21nzMsWqh1wKcwurDoK4GghLdy/UM3gyONWfa4/iIg6b6IzAvmIl5pBakid3Pd6KeWRfThC4oo90
Q4inWMBpKSyeEyutMSo3fpUs+v3rXeBUB6yZDzK7mw3fHQoLQohshcEfMzJ5utYCaU9CW0XtphAI
dpkm3PonnEoLJiEUUOK+Ei8KXG30gUncUGgJpaAEXvScE61Ijf2+QZpBmlwF1EYIDb5Xz1RuEDlE
teNpqzsxPtvm2dg5iF1xvWFSY8mHMEMD7nfKiwhZktR9LlOv39NcJ55TKnxmEFUlzd/jFftyHgQX
5PpPlLnOUTiQlDzAD0AhybigKu6AQS7cWk2fMzxLmLp4ceIjmPE08sKisi/FiEE9Ez2JFp0T0Zlb
HuMqMRhPYXXLbNP0BNMobdBc626PlU7LchnHadH41fDq/AVxq8gEHJnNtuynPAJ2RUvWPcvUXLWy
QTlMSr+gqrcMXYFltmBpW9gBqd88VfykP55CVgHY6KLN62htVBDawSDQLSsBXcyvht3PeBdlVYS4
8gyvFPLKAh5xMyh4SaEWLYHc/uFtKZFbC2m5qZxHzFJ6HddW+4UMJAeggRuWOV8On2okZok5OeQt
5MEMhVJDRaJ2naIZHdq9gfjlpHEEsXyhoh5l1lGyAMp3jsiWj5SqesvuQVe/O+hkDYKvVBdUEjpF
sni9yATrv31fucnZeA8Rsq+Yxt6cu7I2mCQGt1acnTh/WLfNfF9PcGW5JLj9BL1JFLZQcw4asWXK
cL7qt0AAa1mm17ZaDokSX93qEmm+5eLhlYE3mzy7YuDvrsSZZ4MmMnBJ2OVZhPEHFDeExk3aw7PW
+cKiUZ1Gz697SKSq5+QeroEwWt51Kq2ocYfNhpXqIzbT0vraRO6V1SEW9IXwPFW974QisFVT+z7l
mqe+y+nciVzSOMGHulysdic1+YQWKfHbVCksKsACqru9QOLDK4Foqkjc0PFN5exjUUFG0RNRMv7J
SZgralqIgNU3MqWLUp13QoOYaozn18RBecpVvBZinADMMkanytlo1MpHhpGsxnxXvcErgBm4k92r
ItdKvdEEGXoxVYrYEdzYn7+VENNcl03ORKmnjzKIRPgKv58/d69ctoPKdTx42e0ghIHFr+HjJ3zw
tAbSViAMD7cNsW3Wk/hHTm5WQ8W034K1bQW23kurmLncQsPBCQUlXaaoLCBYstYexi1BJtL5Z/Se
3mLEkyOTpy79/4WghZcqmpCCYd5TFEKBtb0NDtjcE5Bjpb5Q1Q2986QITAwi0cm172CeK66KM1lk
v3a3ajWNE5uIU8JjVNA0wm85NVSe+XOvbu+NnbESb+qopcruu8Buzq6oeYsdLCdIl1EuxIr7+0ZN
4nJGQSrEqZhKe2JgGO1XcVyi0dV5DyywY2hYMLzsBk1GfntQD3uGDgq3k48dgVenkOSkV6YvQ6YH
0PaW2oaY3+kzpHIIizhv0qnEJBcRCIptwzcW7GU8dqlBTga4MQdy6jnfUJoz3idbLb+f8HgIXdlX
hlvuhAhE9keIIw3FuNoGt0RpQsI+XnDiqS+Td+naAiFbb3+eMHjLK4DqKl9m7wQiZX18efW2VJKU
d//H3ZtWpfPRi/i3g1Ed6pqSW9zN+5jnnah9Nm5RAc8bYKzbwJlgaSFISV4Fwx3RuSF/x964i5Rt
laCTxBcbQL/1Lj4TLZ/bpXdo9+DBJB9dtZnhWUR3TWG/Zf0WxR4g9n06bdrrB5EQUooISEFqFmzK
+/sn+2sZT7oUY8AKzr2Ed4uZzzwdgm7DjSnM/a+wqPXPtqaOunS8+6dBwxrYJMCjrAmxMNAj9cgp
WihfOZ/U5QtapMadVkgafvkRYTBJSz/r14GN+to3h/HcPwCJjJXEpkp3R3O7jsT85WAPUi8H5AQj
peDMH4zcqigoeVsaIxA/lsnJKyYeBSb5V3k3ZC9dkdR9YMWbdA5Omwn2Rxt0kwFTZibZgz0Hr61N
3MJznG1ylDFKMfd7+CM0p0TcZSehKPpzv0gOaQ1wlKeoVXgd/2F5DUfgiiScr5HlrlmFEjARGNSU
td1lZA0Do1AnWypOsdbZ86EaSdZNPB1PfEnuHell9Bgb1LpJ7emEhX/US8bXRcDDcwpN0QMePVQV
xBH/qLg1i+mSl4925U/YeSQ3XtrTSsSPel0cHx4+fnO17AQY1ChwYs0aK5+Ih/ARxqZ79XQlBfxv
wm4Iu/L7T9S5ZskATsvueLQJbnDEv69s7v1IkfJxIeTzGeAj71uibfsXSoQPn5APUQRL0YWefn7b
qjwDSnnGtxr9m+oXxdn68Wwfd+9i8PWDNTTk6l7KIGlHSFbiEnNRi22+Vp9Tis/IPmzAV6SAKvcE
Odx+jZnMxQlv6ao8rXim2mReNVNzI/chjCCDDPl7hZg1ZQC3Vox0bsmJDKgS8+yQxQqIrHHL51HD
ljTYcE75bLg+yAbFlbg6zoLKLuDxI909wWWnB+LtfGRX4ZN/SIbbFZyye1uXc+kN1eFo6SY4SBRM
yYUbGv+Q7GxcZC6AOHNleyXHZBTQ3UwwcaM3VsUqfpczUnDQeatEvWgRr2tct2CzDHbQzKwqaFat
UnN7p6aVK8Ax1L7mSvfiKRj+o2e1czfN7SGSPwnxpeRObjvXleo+frwcu32qhePbcaPDrc6GRlg9
bLEFkIJ9TGki7AUu+FerEfFXjeu1aenxU+cB0uNYMzQZY4MU8/y+CxFkgk7e7sgmyynwA4ae7yDC
BdDgkiNgG9L2rW6E9zWtGQ/olsFbB/u2VVNq9IrUc3aHMWLW71BzuD6WKEp87h4j+5SrTCHgAEaa
NTptMcWrhWnV80vrLLm9JydcP5Z8suUenbJA53aZQnnP5UJd+BRZ9XMfOfj3Qpa9kxJgKIzKTc1Q
ictFLR4CwM9+uNWwpkp1SZuAxc5HAIbn7CYVNc+xm+NtSR0xatEV4P0v9jT1MYERb7bAqiOMhYTS
oonnazIqZVoTbQHno1st+0vqIbHTrARkW33LU8atSwfXyQ/yl5BTuDrzfXkoYiNlgo91rv+U79o7
c+Q36qw/LRypZ210ck8y0A30O9fI0y19P+sBdssPk319T9BSbir5x+mYK822CowhMira4KuC00J5
6x/NIY6DhSTEpl1V51ySu7irjdixfS5zUyARvtWOMpKW/bExo5IH4R1/vjVjMkGK190P+Hk4Wi1j
HVV58aHHOwyeXp/8BuIpvp8VaACPbKLMwY396hm5ptqU6qUtwSXPOZhJbaSrHMJfU8PV/ZGBtp5G
QM1mjLekr9CUJeWEZuOVL5S2DMzgUKUSv4sbniNf61u3zphUwOyT4tYYta+d4DfbIHTbu3vXEY5r
wbKEphvlKmmfwz66bEmZx1c/Vf1QjLYILu3GNryklma6CPwRYjlxsimtdZpZb33gEUdJaafzyzuB
lIjrwNk30yhBE6uEVfxHUSPB+AdbMm4hhXi+LpNeSN3Rrg3+S62WSdgkOxoOPyAf1lgGNYnHGtAQ
cl6Ia9QH+m9lstxXvgSAEkVgM56L8//IBapi4JERAXuAZh3c9UHNHAuShg2p6rFc+bTyPCta/fDc
xkdQFcO2qKOEWW5H80t7xxr8BUrEVba+U1a7Dqmt9MihtxsSECohLH/TkOBZ2NRTz0bMZSnBDbBc
c2LhQmT0MKvuxoubsI/T3QE4Qf5wjwYXmTF9gekvNl3jhH0mnsS2ktqyTYn3Q+MlEmmqk4xRkOdF
JlixeoIVZaZWSZlHPADFtteTUfSYTaHTQlx4qOEzi15CpMKYJSmHtSZd4LmpkLkyrn3AF5uKz0DV
HZxsWrGHqWJFz3vZj0zRqyQUxVXoepCNNbMEgKMDnszQPSDO8LuNf13b5VV/Q+h48DMUvVgYRDjB
oNN/0lsIgv5qhz8iCZb+NJS//mf703E17q5134mUrkU53bgTB3aL4zuIx+n6Zgar4T5fLzhRLoVY
044+TA4cztfqysMX1a3eAIbFpFH6nRcMHP9ARHAfQ9x6+Eo/WZSn/7eb/UX/s9OAaXpRhFaHTLtZ
clvX75YIWyoMKyKPNPADHWEw9YkiGAFL0cjqxbvKpkU42PirtSu1Zm8k+NGWLFvW3a89MB8pnK85
dCZGxeNXXyhjOKT5mrslQaSyXfTwZK9bQBqINIAAIy2CcgXpY+QE5sJJ+7ALEsmrxxXzXR0iOaCG
XTLoDYwDIcBt97TD4c2WCxs7ovB9zhCsaqrpNDQyHz7/Q5jBL7nDz6C/DorvbFBi+ASZOlZXxdMO
fWVl9dHTR4g5OKwWToefBmZxuFMD1MnyZhQbDaqkpJsJydc6w50CoMgLu85+PDOqFcuCK38rYqsg
r7bcRfxc7KwHm66O8FZCZShlR0s0UneFFfwzZLQEbcjIiHinD0XJ9iCJ+2DKqzG848ygblmj+cWt
29R8yRUzU0roykGrPiRYs6cEyAAJBkSdncKVDLEIyZX7pX0c8JpJtnf81Yp3CHpeZuqoP3R0rFa4
X5/yy3kVyYaLl4GQSRX0V3ovitJ2gvbbij03f5guC6g7KHfwG5e9a8aF8B0exPzO3ToN6wKhOYSM
YRfp/vajK3PDXT1O+cpcq9PLmNIEV31yjgaDxXmfW8luX1Xcg3qV0Fx18gLE9cwzQ6DL6g4DBMcT
X5cM8zmnBUSafKEVlXtkz7ZCeCwqfem0qRXKDVUzndvJXYf7MX1ejpO+covFRVdwXf+PLNHuzYkm
Rjwlgwpn7Fs8AqeNillPgN3GTr80ui6VED2hUuzSQG2F/9VfbpryV/bWu9PZDgDJopccrIZCUHBy
q6n3ciz4lMC5idRAfC75Sg1uk0uf9n2/Gl7lgbzc3pOcjNadlMzhVocJq1x80vPzLW3i04anpy9x
HyEV8Rj4YB2WyPeOBuRjanHQj8/aOm3e24uft2a1UxdQ56FigZmYm0NawXTMU8G3yXmzgG/f43La
0LuLHAeRx2kkK5RDBiFJIEL8MmKBpDESdmlE7732i1KvIuEfEzl+eXNCswCr78tAy0RjNw9az6VA
ZefTJE+i9/Jf9DgRmIvPp41nW27ztwyUDGl+vGmIYBE23/Uyrbao7H1nW5oxkF1LfpX5apAEx0rp
cS3Wrsqd8pF/hg4Fm+aWZ4DQ5wN0Ty99ERvTs08P3mHYjLMVfjyMcdh5OhnVVEf3jTrEzVuTCCS5
DNDOLZrYnt1ccUFnCnk1QiZmHZ2ABmZbj/pnkhlF7gYECXBLJk1oSE44iKFlqXyK0WffCxTcJpZa
7ZfdtDD6fwM0gBySamAtGrAhGESPx1A3VBYbN0w+NUYpf/zD08SAgLBHkF0CKSPvrjCG25hJXgqZ
yfWiKc2QFzleP5NjmU0TSTxX+V/nH6MGYr0WcYtEESXRAt5insCfNmaIBwRbV5AC9wQXRnoyzEZb
3T3SDiF/URB4xlw3vpkUn2G60AQ4qMWiYzKBlPZcWmSvUrsHtdes5L01BqP0boWMfIVdA/MLfLmb
GU6O8U3uNYdTdmCWDPXl9V78jMsrlzfjKjpp8xMghK2yQe6JgLu3u43G8sN8pfiiRiGJpE9gA1QX
AnZgHKz/eDKEPlCLInwKTcJoJ2cHuuhKYLuemnq9/yNiqEzDvVTGaPr5ygPLYY0eMtj0RH1L4U3/
NnGznQV7dlAzh9YUHunwxEgeQeW3WunYdPvwPNWhzmCaJtCkxKdlhVFf+7766yC5Fc3GNOKMtliH
vcYCHZ3zAiDeZWYww4XZti+nfGCdczil2fdNO28SCx5wyTPJW0dM2KeqvrxhRBkZyehuHetWMkOV
oH2BFnzQsJlMnPB9sFC9WZ0DR2Q7L9pg1yo67eJeflX2SbnZ4GeW2b5LVPgkFIGzA2YIpItFmKta
bWKee/ioxg4G64rlzYN+6k30TtlCjZWTfkaREku8xsd5GT58Quie64Wp381erMVktgcP7Vdhquv/
XrMhSmL/m2PgtBJCSdg1/57FV86aFlkt7lPdjf9CW/ocZ6OxDj2nrDW8QrrJw/MoofCSy1ek6AvB
7x6QfGP0uHqtxFY3QzHyjda1vcFXln9n0elzZyeeGL2LLpUtKlR8NCR1Mvggm/6IqODqc6AoLa8+
I0Z6zDZGtMiLoD5GFkLrnJDvSk0y8tSeI/RJPbfyWY1oQjp9/SWS7cziJKp2awnBwDnAMwK8+apz
qYbhdM26+liyLXAnZBfBDKvwt/DexjazaW57ubHuFatKLk/+doH9EGslLWB/i5BlXuQ5/UhPhIeS
zv0CP+JyRPdq2pZ1748GM8pOoB9hg7gTBOj8YFc3akf2KFAsbmi8uQJCIDkWKzLkxkAdMVTV+Kfl
ngbNNXhgScHxgKgOCDjFjosG5YFlFxjFuRkHv32Jv/Kd24DrgPJRYwOf/iyy/tnpbjFtB4Koqq6d
OpeU48bc/N70k+7kBRbiRL5unzxKFz2wl1GXogs20u+HgxnsFXslWytz56ZOuaQ4EwmRetYQsyQe
sZKs9noDDaU3QlXn+bJI0E1J3xq3F2hJaKhcLJZyuEmkYgHCJHjUzvHag57ra2GWhOeZ23gwX7Br
huusskbmIOsISvCxnuX4YbaLue2e33qf5GUk3FfI/2SM/FBErSz+0eshhgvq3/hksjRc3QRclmui
9pPG+aCHwEGwNGycWXxuo62D+J0AZR6sweW4LktaXslIsuvl3TcthZXGO4wTSRRVZ9MrFA5UZO14
4zp4PiOu5tB2F5OWRD2oZPX6Mw/kZpKZY2n0z0r7CgAFZuONZRPuX4U8z/ENEqIIYPgceNPEpGAh
UiVIFNQXRVS1w61QgIVGm7YT68voRFWVX41fWyUw7K51YF+PTjJtX6PuZ5q5Xl/4jNF5Cj7XvUUq
fZMVReR0tC/QGQOQN2EX6Ghdc8n4KiJZskfVxw5dWrz8mnxwih1r6jZvmIBm3DfOWFVMKgDB05AG
1poVHe5Mt0OM/T/rZa1ozGW3cbOnfxyjLnrwMOTkPsblTmxLsElGID8s0APKBpXBCl45tDq28+05
s870BOCDU5tfKYWvtMy4oYzjCdN2IKToL3tDE1G1nb69tw4Olkfu6QVpH2bXA1wdnJdxxTtYZfXG
UCphBQH6SW0CyJRWympEZEg45suggS1VDuDfZHckTiO09OLNKERUCWgWZNmDDNgUaS3yDBoXABK4
9Wyqs4WNVnJjrGq3tAyEHTL0wwKNN/f9/0KWU+tfW4z3RfTp9feFgMI88qd3K3ZsNoMrCBl7kqlk
7y2hocb8wJZFieBwSnTmzxd3Nqx2QDbuSwAI7Pzvw1vvlcxJpeWWjdM/dn2Erj5caH63Y7F3BNnF
WDiBlHqOpiY/3gOmZq1LIdrGvuuizN3MFlMxPotCXPg0OCYkhjUks5l7cBb1fXBCs2ij4lHdJ754
W1i8C35bUHbE+mlZSn5jp6NBwxRwxZYNSc/PoBu7XDlzg5l5v6jsUKM53FL6OajrGhHyLDJDZPig
+O4iG6WzAbyddli5/0xTUj5zUhpwwi/27lb5Tyu9Cmy0WozNCSqxHPqK+MiW21CEr1jrSmGk9Gct
3CaxrKzcaJ1GKGU6yWFerU/Vy3C3E/VAHa2GPGzV7KTA7Qpjta+Kre0fjQqMRGiZx6DFm8eiW9ag
Ll+x74ItPKDHXViLSB1MNiCDq8XxrSAAONMHdezDRK8fEx/pUYkodByMoMSbYWpiDiN7T0ExrbNL
69vbrPEIcXfsOfFaahmiVyUNtbWEVwdJU7ORAuMgA4FevD1xo8xVo5dqk9e9PrU5yQjl3MdoQOTm
xlAIwZTFfEOtOV15wNrp3dquZ1u+gltsUR+9vsNdpBw0R3li6kSNSvksLOstijeG2BvoGr5/37YN
CuNnomGfFWpKtM0jzLLxGVpRHqPsG8HbFvtLKYU12CWNG4g/PEx6htu3tf8iyIW4PrItT8ZLv4LW
SSQStlSYx23EUxDTKlKyy+EQjU2n06a4hWi5nBtM7iP6HUCCHqT5EXMyJNgsRB72SICJTTNbvecp
sz0/lHRD5nEiF635IpTGzPmjbAoxfwbcoIN7Ng+WUVap5mMaXgQnxhaHC3mHfaMLkNAcZWeD6CM8
fOX49WD8CnPwbqjl/XfF2rVZV2uO/6OTgvTOwUUvVJnrfZchhwfCULQi9dciZANFQ4YXRWdg4e9Y
t2hXVY+IztxD03iwZ/Y9d7YWsgLZTl6dpcP3xwK00xUgKfUKVmyHyBGSbEhkWbvxG4mi0dOD+a1h
lJaRsBb5MnG7Xz1nq1SrAyjka0x2JFKVGUbdTCWZ6WBsXX1nglvzPceWVvtDkh4VFU9ifSYYrU1g
bhgl1iZKusn+VCk/OImxSqjlhHEAq04awkpvLIsvlLxcJT02gowyEmuwOUt30TeO2FSgY3HrP2Gi
lbqtETToshfP4zeZaB0SDNE2HyJuVQUKrIZKolGD9sCmPtf9h99UKbUikdizRiwiyvGi+VntRoTD
k2qS6JxiwWuYkV0lLcZzNv8/wFt7Xfno9jvefXBIrNqGwd8luSBgbF/LnTS4InkuDeG/v5+85/i1
wzwOoj++ctD28ZjJbavQLU8qLPGHIjusVEsPGkd1UfSI7yln9+2Eh3lj1Z87MspLB/HDgR0XgRGW
EoP1P2OXQnBd3Pn2R2s1X7glfwhKaVutbTIyU2Vaw0wdH0dDZHGuLmPOyUzKOgft+IgYFZcYhGid
Be00I//FeIiLl5ZgI4HfNhMzYo/ib0QB7NAkVOHfIoMXKDBd7TdVNh7TnfWMIFUdMdUzRyA7S8h8
Ubfk3FESG6mGFhHTJRZnDDA0ZEFeJMAJO6UipPV/BH5uiHbpT0qTu2jmlbbW/4uYwYhX3AOjNp+Q
9zScx4gW05hAOh1PSVMXNkMfCXlHpfxmZggiHNZDT/LjI8OBGuKTuVlEJJYxYS9DSNvNbSsIP+j9
1dbriaajpYvTO/6hZXxUARX5U5l6nH9Qv1Iky+PgKHa4rtJjEzRdZVhhMSf/4VrCPsyT8e5bxl6P
r6AyN5irZlkrqYMAoBIpTpiK+kzVLIrJVXy8h72vtAJb0NkRvTaRJqZ0rBTQUiRrFC/4kR1Me42F
PY3b6mJ1+QyGW4/OU1+uEq6x9DE8+JK/FrB5xtW2b/67Xv3ff6mKVLou1lcdSdN4Kn6Uzya6sPjO
kojf30qpLPqsOrmx3KaMfPb3eULdRs67/MbUiVrTvxb620B6WLO9rcY/Ssp2Py2nZiHFXy04+fpP
v/UN5/jsCqTLRlkd6A2rAyLdLqguKHv1p3OyKuBuK+z7GRFeDPxvATdbBKvhJcbfpBO7tqYaE28Y
PVtdnt1HKHRU9KlUyyCjtTGQhI6Ei8mISFnHgqDO2mhEQoKi9a5Y+i4j0VoRzOVuDig73XJQK4f/
7aZpYEPpMsfxJdlkmkVHsNzeBTrJVzB9L5Xi4aBpyfd1EP70KPZAlOaKCVPlAIPLxsq8y0vpweuz
G5M8LESpfWak3T+wBhgD6Wm80dgMseajJ55HuZ2ecng/HWMoUyZPmj2U2vJwIpejXL9kNJ0+V7JU
7MrMIKrtUlMWGTYf4UGrkCBNISZsyerx6NcCGy3Px7/Na4o3dxhJ6jCBTgGLlu9kdupmzak1HO7U
kQwmwfbK0nJ7pqpkTG9oEaIimtSzNwgNJAvX6TP/xLEg0Tczmne2PUJPBDvtFH2uGrG8IQEkOU6c
0hvbtXeqUPg0GCMavUe2EHz/iydA15+OPHtls6BJmFzzIm3yAuBvgEKYaIDyTYKiIDPXR+9dHZw6
6CTq20dNZt1jkM/tqdhfrVA9vk7dPpCDJW/0V/888FkteGwHrRSQrEfd7om6RtU0IQvP+Z5ga4j4
mqOIDaWpYbeHK+qa3lIrj1to3IzqYuvzVtwTpwE6Zb3p6sIdtr1rJs3zmus6bFET+Dzur6sTetxn
NIi3KRK0ukKsE8MSYxlb8Cn6TWgD1786WbV3IJiv2s7ztCxY9JiJFL50Aea18R0h2PY6/gywLVSj
BY1OFGxiTTmjd+jWNg3QPyUOui+PRupoPTYobnOgw7AlZGj72t0nW1c5R+BgvSD0sytRCFhVquHB
Jyos3cytdD6Jqi2gqPlnphs1XiryIT1HLILiuY85WJ07CzDwMBGAgErQkJggwaqPdAD+RpySeiMj
BxusO9BePHAtcIRSxLFjLL9yGMgfkxUB7ZZi9PEqMdaFJFLuCrfgdda3jxdR/xzlDaz1HSIfXYqT
V+qqEBDeS883+SiMgN6fa1i2lgo9QVTC9U3xhoYBUwU4Ld7BDDY0LgteUXN6AG2Ksu6hGCsnVB3o
9voQNKQ2M8uJHzwy9V/mcI33ck221WVYrLikxo0FzzSWfLrX7KLsFSzZMHXVo0Ctrfn2aCtvg/nn
nnWEKw/7UtZNB2KfuX6wItIJGBIuRW4mvE2AbEpfFul8ivYSIN6Vgtbv//o4hgKWvBbaBNUNjIQ4
14p/gKcYbw1Q9DolYA5AbH4MEf85f6Ba9+Df677aP1WxutlqViVgkQAIDFhiAZxGZ7Ve6Vbpk9Qi
q49zEoieLNuc2Szo8ehJLvxPqPFJBd/FPEKIyKxnkn63VaP+Yxpahy+93jyqloGZ3k2jJNIKujYF
LHmxnnft3cqZhoUYqp1p9ZBg489Kk5bKOc8067MGEBXwgYRcAYb+m61OiN1c7f+N0UhUWopTulvT
6H16B262tn0tcsD9d9xP3mgUfjk/sn5OOgAJgwqY4czzVogw7qZUe9ZMCF+/4zu9oWA3Hn2JjBnO
fEBnrS6wPFIM1ROTGprj9BmRzqCdxotV4ROdnioFwvSn9V7QAuMnINtzEMZ/hZvyTYHXYcRHpjyG
UdppsrS14dF+2JkGOP9F4bObLES+1+djr76AYiJp3gP8gFXwBQqymx3C7ImqZrtO5g/rEEjVMoTB
0cRG8amoqLRsNy22/MfG2eBMgsfkNpkdpz6pab7K3YCgZC5W8yEdBRaIH7TryjfwPY8USkfglVVg
xQqqMgYXuVNkwLjWBgtz09g49SDsi/esLV7JYWYc4w98g8ACHgsAzboZoJU3k48dpCuBg3QWzLzv
BvjHmHFio92MNmRZNnpXMRB738VyHUQ1uOsthhomNTbgeEU6v1MMIUcnomXp/UKUnDfZSEAICGxX
1RUF+Znkh6+cFmP7l2Y1p5qfM0W4Si209HfKwH08jpcQNxO+zgAjvsPNezeRKxNqPn9wG5/NjbCK
NLqNo63AMPUX6GxRx3brmlJQIYlfcGANjVcAzY2Qx+UaKVYkYB2t+mfb5yCohPLyigA2E0598c+5
xalIl/6U0i4RwB7nbz6kff87KScvrp9OoZX2yG7yqQpzpO0MY/k9r8dIGD2sbVSHnLd+wI74l/6o
TEYnx9RYnyA1NCSadStTo2wjpMxYJYSDeDDtDb20z/nP25AZA5TjrAiCsMmWpBBvYqXNP3du5tiD
hNu+QNRt1czS+d0F8f9T6ohCEYSeccAhI2FJwTnntH4YQT0ub64q+i+y59s7v9KTNeO2J9C6QHUE
A29zo1+9kFKz3biTjkXsUfK60nTCABBlZBxS0eNuWF8F0rPel/b5yLnDsbju7jrX3zRK/G9oWF0M
o6uS2eoDIjlUJli/w1UTHUq7lLjbHwRt2aLpAdA9yAvpukspTOiRItRrww4R90PxQZRfuf2cmnfK
pdDu6D7TuAXC21KiCXer+/ikRKfh9jwFKgi1o888n+84PeCPAkhAhQZV2SrAdBmpqufbByxAB6qX
+ST1aZMcpanOHwI3tARPBjH5ExRgoswZeeLXBuJF5OewvtCfVWHL4wvZKieBoopxopxLvhLAyAFD
KYsZuEJ3dVd6U+dmjI7Wy/DpK5Sl3qBpjEqLA5JU2PzrfkhYGn9vJlps0Mlo6sDTVoCpCj7Xyc0F
T8V+GNe8sc7vs7ogr6nuMFp+o++GZNFa0VyDJvr0AkLAh05YQ/DovWcs5GNROgHAxnQj9kC1/gRN
yGdsMM4dh0MkuKaNe5oUg8EwIcz+EVyYneYB+6LOcawz5/6nSA+MiTTGUSf0gGSp2DqTGT4zPPSw
WRtpL6xgI0b6oslAXu1y0JhR6+w9CbQltHDTGYilA9bck4lDNp0LcTzKu6yQqIcdZefeUeZglXqN
6cJ5cq7E09xVaqkPzHiMVONtv0MnKg7E2QADqLW+zn6zDXYZ4tumkU9EsBL8NQlJCUU8ErJleX8k
l8EDtuoMVqeyMaQCbFZjYSRdU7KFGxWOlt7rI83iMwxX96zoRKycdn3R0JxQ3lo4zAnvOAlWe8mS
GwD1cy3gJZeUclfdsBpwfUmexhX88B4swIfN4QAvd/WwiYQk0AIbG+ICKCb36QriraxW/LbTJ9+7
soZEvp+ubyS8j6uBSRy6r+3flb6i1jfeOpho45XmFhAO69tmka36VkMPXl+Zq0a4iScoeqcLnfwX
1WITAggtBXKsJ3WmoyA9pAwXwAwuHNWtIO73oR8A5ceTbuUKVmx2ohz9v2SVk7h8U7d8O9FZaibN
UqAC6LjOwE0/8xBxgJIpGA/ZKdP5BT8z+8AXyqgZo0VoZT3wJ1DSC/9ylaQmDXXxqiZ6zexd/2pd
IEZ5PFh9FsC+XNvWLP9uZfbAasbOAj7CNTF6P4CJk+8h+We4oEL1e0nt1b7U0KlPd/pJEC+zxzPI
ej1ZpdqJzTM+V4/M1FtzPicPyd4D651X98CjmCeSUKZdKT6d4jQDjeIcpRJr0nBM2uuvX9QWhmFq
z5lOymauCUmafylTR+epRsYQjafpnbMCdXU74fdN83lc7UGdaJJC2B7eLuXInzxgKQQxFPdndVsz
so0quB64+0ic/KWk4uJuea9P1wajGdL/BLS7FtNkb2NGVWodLLuLLfr3WHN/yH9sYs84b/vcQLNK
7qrTTrK8wS1sAd+Jn+7rA0mi2HH8V6iGi6aNRQGt9fUtD/zwPhEpzsyaos65alHinan2FDJ9j+7G
sbH8GAAdZcCXi0x8QiQVlvmCYkIn6E3me04dMvtBBxPuMm8xOQxNamR2+GoQ+oM4vRfxCi/hmulR
KujJt/qi3Tb50xgj/eiuDeyDWzPAIKaL7x3YKYZV5G2ul0hoxlCNt7vnLdfqoMdT9/n4sNgwhNIA
tPBlCcY+ebDwS4dw7pHdAob3j+Rvgjp2HXKLZH1QgK5XmapsM+aEpEF0tapnZuioS6ZQ7mhq5/F3
CX+oiW19O8wQyI8HeNV+YHnSfCetbgROfE7VJz6AyGKaZL2fzKUpj/PRJMGquUw1Ln+BEnYbi++a
tzzUKRl/hYOxy3CpIFvYnizf3/T+uCfm4RWTRucZLdb9s8+mUCRs30VYvY20IXPxe/FYM9cAWAft
t8a3p5xbIMxTe+9CCS9UtvNSnBfjU3Zx6m9SLPt4+HSEUls3OQ81/x0eHYNugNTZ9muYr1Ppx60P
dfLVmxA2nAr4P4dLH1F7WyT8OaMybIeFUfItk5fT45TULQF61i4QTEDbBVPm14GiXL9DjOt5i6Cw
i26RIkl1f1vEbRK2dpsscKfOsxS000c0FhyPF4PN91Hz9r2/Ygb2I0tgOX9zorZqFb62nwaAcYlb
u595oCwnyNtzBNgGuvlDgWGY+vGF4S+Wtt298Y5Uqw5kP+yAv5KZp5a+iyRMUOEHH/Psn2A1MSAO
v/j6PXPBHO8fhuZ7lVffPX/20fO3VNsjucigR+g5GwXftZI1QYcSXHGBD3aWHcf4KuTMmYQ/nC9E
1MO6jNK6KGgMgKpe3o6H2tEmK79ikk6jq1Iw9/YHa5qmkaNMYVV5wMddJ5NIvcCXwIBk2Xk9nZSh
xbffKb7MucSnW5zKUHnEryB6+SaBbESf31oKomSBcmNyw0A6dqDXqJU8RmLnSGd2Y+yZj6Fl37e4
r38e0xtUepNmMOJJPzzSWMMn0IX8MDtfJAizizNPXsbG1LZVVifvoG4w6h/rkwJGVHW4y+zQl5mO
Dfic0qGi5kxXgdlEcsJk/qYdLAvFROApCM18vNSlUu2pK164nmOQMNPtnkr9jeUSuVYOrIl3/uZX
KD0poFJDtsV+srG1EtGEqael7ce84WdXrC+QjSTnte6TmC177iszUWNL7lv0cI2jLibh2VedmKZK
FAwI/cp/wtd+YHvvIOqSalpFT0iYoUHQzrrkvUYLaE4Byr4CkgKDzIF/kjJiu1ABa16hWapN3wWa
YuCFF8hGQ2sjObgIdfp/jNNIdTBNNSiZRJwb235XryJFaJqv/hPQBAIMPERpSeYCjS2mXKrOaJca
echJgu1JxSScTFRZ5jHUVh+LHiyFmtgfHmoLvdkQexDcmzBO9POZYIpJv3a8jb4a86dzEtOzy1RY
MnlDN8gzYrdGczHgs6ZXz+yeJVlRekyHFd9WlyssvPdrKswz3f9Bw0Di8lCZ9d+4P1j1Y5KpKu/W
tkfpnrOayJZbUFByJrCdm/1RcXLSunEAdjVS1Sx2ZiH3z3yG1KBrWkbkZ9Oa9JAmhPmh5jd82PKl
oUpvPkys79OqbPqMwJJS6Db7/W2q7HAiWFon6sG9Te+DcWOdlpIj8+JbCb9LP0QNfKKAr9ql0XVI
85lpDEwk66S/8/m1FcItEEOLjKCwqtKZaI/Bbkju8nVdpMkfA1P2Kspik4QlvASS9y1vUngYSkVm
oJtFlkmRb67DvzTkXEeNhtOCcncvyY+Mc4/LFBsfJ+LpjfRCwtsohc9xU/U/5PptgRLOmKsxLNmp
JFT5r/Nc4f4oYNe32kfDqobms0qBl2CUSp3hT1d5b+norlRTPVi70iE5rBJXgpW1pxRCvb4CFGRz
wECCJ+RP7nxloXGgyQVey812yZ35rTHB5M4TEV78dO4EhT5zAPYd5+BkiUG3VK5/Q4BsSsvHx1SS
bntRFc3b7i9VG4OFDVP0WxIWl5j6ZIxFSYlelTWtrlkqeTaBesJ5u4P6/VWU9fsST8fxqIEtxV9V
8SHQkMLDr7wHGIWLmeu/bo7K+sgQngqOOQ7ZkWbH/qOAlK88oIv8OuZH6YORvETfaAO7MQvxY/EK
qnX/4gBb/57Y3fF4c3sdWLmG4r4e+gTgFHLcHZcFVrsSMBw2egaoZQl7BuyVytc6g4BKvF3tKyl6
VungSQnaCcM9u91WtsKkmTNJD/XHZctzuG6ST3V9JEyUkgspgVPxxXUXHOpyLChUoPL8aqyQhd0A
T58wbh4ZlTqgGuuQX3Fe/qRZ78ZvFqbQEXMUCovBNtywjnb3kL70B3+5DPQKymC58yfb+7ES7kGs
rpEvo9oxa2B578tb8USUXq8gF5Q4HgUSnWVcp3nqbr91O2YDP37ZuHUyVDyNYJe+jIe6NQZyBWbb
b3SXTDmj6sgB1AQoTJ6LL+vR3K/7tTzL4dM7qYFnjSLeV05GhHVNNpURF+gtgO8ZEfyQDN3RU9B8
xaZLxIG86tY2zVQ35WEqBtnAiLOjzxlSkGqag2GE8JSZBjVOrJ6hHckzTKFZNlW6kkyuYXj1j8zw
TFLkLr2R/7zYKRF4dv1Ho0Klnk3NQm1HpaT9j54Bu9QMvhaVZ4aa1flDKnkZWGx+10AydurjDit0
OQsVLF2wo7VSU6/qNY0TwEqvqrJmdR6d6u9XKnfais7EuLVNAp3fvw0vyele8ViX94I3DOmivZbE
5edPAHGTn4ysOSYQLyQiaBt5INPZqYSN/lDsOK2gpyTYGu/xDZ1Yl8hsF7iLam9PHQDrc69D6Zzc
8aZE0HHn/t0CWOOEhbKcSYrmRWD1mEWSJI1DOc1NGueJ1rVfH5RZv7Sgh6zpwEDKSQREYjaZ9FtI
F85L/i/Mufw7//AyoXTPl3LyyWV40zp6e5BGaj8+CW2Ug2ZkrVHJ/qNcI5678Z9kSCCQAqb++IP8
/6S492GcjUaCGd2N2VOSuHJ7Y85qO6dJGthBYrHJWURQgDzDjyzUkyGsQQxW0QpVtLmqx6db4VBH
dghOrE3TU/RtZqEFva4qK9SDC6wNPJygAY+ztYMBORIRm4TFlbpIpONZg3ReTkbNf2y5GTQfjuGh
Z1GG1A4VSf2tML1Efag83sanMAPzOxd6ZpBybfLY3ji2L4BWAjlIabHZ4GTRkAiYEakib0lIav/P
XSLEma8nfPpsxTWDu5Oa9buJSNUsiwRUpVjICeIsu/1xVsBMoDtWISdtp0uc8Sb2tjcoO0A5Rtq7
0s6gZ/VpIyswGiZ6WeJ3aDLHHnORZfeLJ+DvBOeoQZi5g4dX4/k2RCGtY7ny33/UWq6+ZUJ5nBNH
XXehdV5Ate8ZZQuRq5vVL4JyUMWP2vyVApE86Aiw33x/1pmocPeCKXHqqdF/vuwN6R2zJlUDxhFX
ZSLUfZSIoIYSHOJV1VtEnSIVyHTyP5IlDosW75Q+zjWwfz70aL0IXmiYptOAB2e5l4nGb3zhObJ/
98d+tIUjlnrhiOFmK+CelVJT1umjQ+ZQ/1Q7FpsXSx3gbHJvYaxMC3b2+Sre+v2nS29+XP8BuKGA
EhGtsMCAoCVxKrHNwBGfUxm/wlvkGqK4xIUgKbTtMZRzcJ4a+s7PvNoKjn7RG0ZSq+d1yRaETx4r
PABbcD0Qqukvl4mG3xbFUytlyNO3xJd73XwWD+UVYQ+qeRlHuvpefFb06Y4xOLqCDTL96H0zIt6S
vlEBkk95Iu7AI3O/OuGlQ5UXQKYOGSDgNxOE1QC0eqrvcqR5oOghfBN5Rm2D4ibi46RojZAhdQKU
Z3DgU+fSUrhrhOx8Use7XdNo4VO8JEcM3uglczGRIhvg6Y8Gu/ioXJIYySSrjHqaIiqd13dKL5uh
2maU/7N69zGEeNtJr/PEGQAh+LhVcBh08oungc6alujI6rQ6nxqkdc+nBzsMFcvYZlTnMf7UG8dq
ZnOEyq2NLQePB1XNQkwp3kLTfdvGdz9+iyT5a69+PN5kfsybkaeN6d6+Ls1x8UJ8pUZLluIKpXmr
/f1vLN393cr0D0qcOG3n0ZpUzkLDsN2gkdt4Zzw03zYsk/pU4rglGs4XplurSXsbs35LLsFgmHBv
hZSpDZarNihB3X6NYrDb60S3iL7lfRyyUr/ePLFxnS5IeDlpUQmx5f7SheyTRQdM9NjaYJ+BloSf
HaaTzknz93nIxveWgT/FBj9yjgmC36QZUyMZ4fTAAys27XKERzl05eZqSMVUcHPhB7qWMzfheO8R
pukY3BQ1qwzqiTRAGwkedUXFCsF7QKXJf5/j90FnPt+1ULlEAm2w52Z1AEjhqP81NlH8983zsdRW
NX5gYumsP59GLB+NRcajG62rfvZaqZSVK66s8LlntiBj5etNkcDAbDHwTpc0pgCwHCV03du/tkBq
1Q4W5GfkpVmLpiPIJvhoOBVSsdVrVf3GcrUjAMiSJjb6hBdkFFhdGh5Bq80job2l9aSyLTaQss/e
gacfpFGVt4yoKJa5kyf42gxZ1X1j5pIP+WYOSk6gUZzMam72G/0e8Cyziwsl77knmW5KGUpPVONm
O7CNSxoEq/UFYy6b9hmhH5vitYt1pFWA4SccwmjlGK2LSxv1dpiuepVWfSJAYRkMWkVvHz86/iDQ
BQqp/u8AfBB5HLUxjjZJtWQW84FQxZA4ABRc0LbRx/Sr1YNFmFOa21OJznDpr9/1cmDWCRZKMo6k
YVCOEmDkOGuSnd317jFV1WPBNwxnkNnKXjV8mLDRSjdyKEhfGdQZ+/ztyLSiLS4L0fZwuYAvpg8I
hd5TewRtR5/hP9TTX6YNnuuNCEp6YUgaVX623ESlyWW23UTdzEG+GM4VgyTaoRlMsu3hCvxtqIRD
/DjNvy0mPDv7ilaMX3c+OVy0uYkVLfwVOXGmws5NJtB+g4EfhA7u+CBviqbTVMjN1n6tCwxZqknF
sx703k0TDuswohiHVCoVR6OLAqWLvvH0khhoKRUdb76RoCe08Sf4FpJX9P682mHUL2WJ48LRQKAD
pm4q0Vf6d+EDEWQQAa8XR+pzObipJ/XmZisuVk+9//UQfj1sZqX7PEqnPQp2U4RHFUNxgJf2MQKq
g8WMIaBOgbExCD0SyLT6ycpVkeLN2Fwni69AVC28IN3yY6DnjiLN/pHrtoQDwUrsoArlAPc2oTRO
Qr+agPhTgFw+sSD1wM8qvD7ci2+s795ayjy7DHgV8VGePHrA8jTKwDqNSqB+vFM1kI6i4VjUsphZ
BX/MqYz7HAnKiqXzJcilQwJlFlfq7/GZQk2S+Y7p/YYs98ETZu7f6rPzP0RXPKdCaICn7OyXZN5g
A8aQmtW9Aa7yVZ2v0jbajxBUwSFixE4ymzKP6i1Kzc1JntPSRlseSYD4Xf5oJFsGiIVFA0RATKeC
niyw5RBdgMT6+fHh3vBc2K+W47jOmjyKDRpTQ5eViwzFvbqTxKLufeFgyRf0RdDkIiiGCi5iesCD
f37VHHlIPNfeiPsvVs/pjH/2RiYtGMiJPZlx5i2AzzUonbIQ4kUckiINGTz8NRSi3NfO1Y6QEyZk
84AbHpttPlUivrIA5mK0Xh/nnYHXd94MZx9ah191novGddWJmF5lWtd5jGLNn00kQyJWilRO6lyt
c/letMDxwKJiDTzNlv4u+cKGG+4JHjyHHnwx6FzJIB/wd14RbSHxz3Rxovtp3IZSkKEIhUjk8Vmv
XpoeyiyafMPppU92SxaMdSd+iu4yFOGXvE4wLIWHTp5XSyzk7e2m/OZ5hReLm3mYBCRB2D5zAulp
kpusWKCcdlB+S4k80pNBBUxZ+3L1oIcZfJMenqM2BjN4Yc2cif1HpfLyk7je+FwVguthPby86rZH
YOIQLO364QylAQpqsq4kNpdBaulG56aYPwjX/IcAGnP4lL7Eb0bSiPXy3IsehIJ/pv1/WbJp3QyH
xvTRnfWMQFoBk8BkHiOjNGDjSiIthsDAERok5j1fITNXLeqFsw161428Yx+wErorymDCWdlQgXjd
PxWSDFNagwMBrX9g0XOUjSymcnyclwFWOdsGwyIiwegJJ5yw7kGYrutP6loRCxzQ/MBkyM/Oepkj
2Jibxff4KK+ANilZ/axpL8R7Kvxyu3kHAEwQJ5MdkJowc3ODPddgRcrRTGZh9rP3/hDwjEc6dLkh
XeObbjHeQUa1Wah0fggReihdL4xRmFQHjarodFFY1kTBTRhs+Tk4qwaM8f48Wam7gapy1kTcie9j
rmoIwdxgYqXNp8QxhczgllTjIT/FwQ7FXDEDB5LG5ePDxhSNTXPS+mvURGoa6FsCfHWxj5/q36vC
KyIX93HNnS2x4Oqp5JlfNQlFDrwf2AjH78e023UbSO9RYgzb2T4S/0QUS1vaxxTdSYtHMP9wLpXy
rkVivtV9hQPxy1UYGl5NeL+R0YmdTZQ3esUIdifWZNDyaSeE+KnGM+Ac/f2tEBm/r2oyUi4BEBWO
D317W6nJP4f/dz8qORJRYD6P3I4r9s9YpPIeYMwJLtIBMnKiq8U/71AUHJZ17vAqCdx8iBD9GdC+
oNQ6evrUCOj4RB/BGLsKVMhcZiTA1eGHniCMOLnUdTdH0FrAhVJS3svpSwyf75E94OUq14yNvaKC
lmjLc8WXqPqCX+PkSj4Vz/jfBD/xr0RxJi+DlZD+qAViq2PBoZJ5VjA05gi5c/AlwjYtY5t3wCKE
PRPm4E2Eo/zlQ800Red3+bu6cZt9Qws3uZXA48q0ocAk3YNwQlmcI1+lDZ6WKck2HOoQJrQw1cw/
cnRtRf9goHXkDllE6n2GT6cdk6m8F8SJumYMqjsCpm3uEyNjKlliFJAaQ+wm6EyvUTHMI8jVssHk
V1c6GOg5j8T0yTaPOKjBmhb1QwVOP7iA7D/qQGn5vbV+cSBVKPB7Si7SbfnTN+l/R50SetViA+au
Ptjyvff2cZJun1NzAjMzJNid8h4CMxjoxMdPSgshOeaBv/FHNMJwVukXDzuxvu6jfJFZeG4YEfBc
fro1YqdOtHtk64yg93mmpoT2dzqyoI+mcg3KEy4qOODBY6pUH7sZER7UCH4jZ3wwrCujEcNFwu+w
XDTJSLmjc/rS3yLIfQjpdBKQz2ADp0BEQjhHso7nCEbXZDapVR/D/MKQ3j8Wsj9Zf/YZxQ1V0ttu
RtKI85dXRUQLjTw+kIi8irsfSX0AjMM/lWq+pKVe6Amn31efj6RuwIQWCxKH4uubxWmsAbJihOtb
SA5RDoWAHO8bSD13J3qsTQiCTE57uKj6rBwIaHdnK9scvDhq3SQ6ako2EVuEpz1KhacacSR7u8eg
GaD6J6then9oS6VsKfIYD4ahsT5FhB5rdbjhdj76c8GpFnoQnCXrNVkk81LAyD+vlRZyiERanQ+L
8CyK2VmF6hNNpaT3kWWsihk0i/LPVp3GMnVLfKFovP79Ws5cuiFimqeLFZlffQZqhiGav92uURkt
FriyUWQIfuEI35YMzWBO/hJZX5GbYwcZNvZk82P/M0iIKrS+Hrsp5WE820zVmgQvM74YXtesiYB+
ww7tjy9FkBwmkHpkoj7ncrl9FfH6i2Hh8kYK28Kps5G8pxIE1diBpVfbpWZmG0/hs80rwN+JRrw+
EjjrR2EYnhm730G4C0vobzHzAVvVvfMvAipz9PfcWIWTC+ej+ANTQwxtldB8spUYw7yjyrNpn6x3
lAU24X9opgs4PoJBgmslWutv/cukp8bp3hIEocL78Nx2SCbjwNmJJDus324mywD79WGAWp4L37dy
XPKxN3/wntWmDew4AYGkzws6GUvoAH3EtTuNc6yd1y8mGxR/ORjXkPPT7OmTJs2RtYXUKv7fVtMK
lTkI0zRnFtb4fUVtDATVE70raJJCqqW+ch9UtGdozpgC2jHHH0gfl5Lpb8dXaCBU1LYG3qEheAuM
NeBrDYPT4TDH+vmsHkQSteT2L6TmzwMLdGTdh0c6FAdarmPCnlovZJCQzP3hUt2dSMRuFO2UUoc0
98l26Yfe23QtzUcnd7AoTw+GRdgrDp1HQ0bYIyXjNwnHR5wTiTy2b/gH47EOFLU7jWL9nlLqa94+
oExTHHLsNYohi0MjexsFx1fkbbU2hLZp8dDBM6tK/LI0VRLHvpUHOV9R/RFJ0FTDTQF2kFtc0POw
hdAZpuVwWIOOv1ZnppqVZ7uAOrf9ZOx7rK++fedGI/bzhVshrsLWN4c2kFhx8im+TisiJGROJLvl
IZ3e3AfpLwgQf60PG7Ybyu6DkisO/iHloGKauJoJ502aTgNh5blHo6+qTYM+3d+dkp12kV2CYfDV
eBHfCcGLzTgiE/wirkxu/sms3YQnAelUori4o2FUfyf5LX0ogsTIsVBuDsXi4zAS1v6+WUsTb4jX
PC2USSDizFABXw+K8mOOiaEcqM8i6mx82J+NM0tjy6mgvCpqTCSo0rMg9+PSV1OPUPw4bPJAc759
94CuN4OlKjXG6tNSaDq/aEyzWK71VJSjhJYS33Z6Uziq6mCCssK6ifOIeqXTVlCFCHFO6QYfhz75
cndm24JOjFro9k1aGCTpi1DcY12msPd2z7qzuaHQusPi5Ht9donRb0ZK6E3dH+j3XykvJ+StAWFc
BTu7vU3bat6b1YQ4B1Avp+ETVEhf8WZ0PtVm19kFTaB3v/XalbYghhDZMZmU/YhmRLA44NKuLtF9
Dm3YfrI5+xUjXw2P5QQLnLnvxWYrbqMCjG9oYPbqZ3IzSOk6KfM+tAEyX/UHSkcvY+X2zoeS6/Ps
TciCi9ibKIAPiE+PQXdHiV3/003dSU8pYzRpt2P7t4STlL2SyrN2Opfm/2m79/7OfVIYRcYNsDG6
SOCM+YOosTL+8c1VN+fu2InW6z9H5loWJi2WYsD3UuH9S7sX2JaGH+cY4tzfbNJcPUV2Hx+yDmNs
53cf0EUc6KVVxzTE8qA4rqX5bpOy2pFasfI0BFJtMVkYx62L/t3YQH0sxoR+nCtgKjzCpSPt/Sx7
3vOUO3TWanL4yYlAo+thhacn04J2djhbVXaKchoUZU2OTZFdsjNDXglZ2m8Ft0nCKznZQRUigZQD
AcBIEpRAFCBTgs8rFt87F/9NasPyBZwQ59sqNAYybeBvznNLxAvURgz9iEzdlfgX7wnw8JFNr2KZ
rMAvfAaipxBzYSc9Jw24m8SMy+vF+ATZg1VNlmGsTo4vBZk4sir5vC0cOwpk3BDE6HmzX/k0wj7S
1G9FadD0+LwpD2URcrB3dhdNMOWF/GVJvpztLukPrKLUn6QeXxIoUVqRdjkS0sdOfTN7WQtXI9ZV
WSVyABA/TW0gDfQoFRbVeQsvzWqEttkcnsHIXk/6WxtCafazbbnrwdgg2d7Pvh/J/opJXA/cHrrV
kdLo+zbtl2oXtc+N2/s+VACWHZSo05x5yAbj/H9aWorbs0kFQ/s2JCIV63mupLYWhp6N7hLRD+hL
hWuh04u57pzDYywrAafrnDw31IzvxBTnbK75Fz1aDBU4IrJbaW4gyW7dIErpmfRDGTD9TRuBOhAd
uPC5mqmiH6/IG+gY9Hi+Wt5SHqZGGtL8hPEmOWseXJBSoKIk75pU2GsxF/J2MOFuwY6XwfaQeOhQ
UXeD61p82J3gJJjM48576d/6JlrieE5Yue9RZvVlHrI9YXsTAl01OIoiGQy4CKmp5EQxq64mBKp7
lo7yWeVpww+uPnHG6C60TXT6fUPcJvxjjEqRcXX5WMiv6pGiZT0+fqNWM7SjUa5iTydL/e8/nX1R
0TLQmo8AVpuf93jIvdk5UOpdInuwdj2DpR9gQPKzONB06h/7ZfQsrqB0WwIhdtYc14Og9yizTJMz
LTbiRvmj9KsJ4oRj/iyOVVnmoI6rU/h47Dyen+jiu3ieRoFnDeJAv5fJWIlFIEZECEelfloXIqom
DHx4WzEhhWgjKqXh1DGBcQkzY7ZEPTe40z32rrb+y/9eqMq7rRmDlorBn1jXG4YBZR52Pl3DoCLS
4YXE5Tz0Qh8Kqu1xtpjnO3llFlnTe2SddFqRRnuMcX/+HY/lEMSuXEDze6KpdGGxN/9Ksu3KBEv7
jc+BWUAkqkgZNseSSAbK9fyMUePFXKUrgxKX9WnMOy72LSusQTuDjoAKJ8gDB1044kSREedWcqkN
RehZgxtstdmlg+5ozV1SLQBbofrkm94EXYSo7XQpOgoi+xFrAbIQPkvj35U2qDTqkotooyaUKHeA
knFvacpU5NBezPPHqqBcEcMgURBO9FAXBTHq3mhvJtEDXyBTP4ya5qUL1yDcYoISUrUOwBakujip
PvEhgQ4NFMLSu/oDZWs6PIHlkD+hLe3JIcZU5WmxpfP4VuMdCtS9nKB4dL5sUzIRt+kAB5SQfewa
msE8wd40aBDJG/8qiF7rrIEfhKX7V0X2Na1wEsE17tmHsEpSx8LO1/F3CgKeMs3TOZZSFeO9JlHJ
Uzh4t8BpVrdleddy/xTDqsc51U4KFtrOrDqImjRHUC2yVYkKcbY0081Rf92SQ2cuXh60YWeVs9jc
VBIvXZYSiFQjXCXg6T3dZtI+C0xZPJXAmeequIXu8NHRB587kJFz42mXWm6Zb5LaWlqVpIfADmjO
Gag3NLyGROJZrSMeeZmW271czxg7VXwvPJbSD4eCxC8o19UYZmw4sOEvgD0Kc1fsg/vnOzqh6hip
uOZrIa9ou8WRXz+Qeq5lte8d363WIVgrBXyU+iw9wOIk+QeYfvOA52cx581aPxm+sNvC30HbyRN6
dRrInYLrpdNGyfSNi1kGrb7ti+DEJXPeJh3VT42oF7hZM7ugwH0ZwmypPKwSy52CLKRUhrd/CMvk
A1m7XqxZb3SSKg/ef5AxCmbmqCyPiWYz4yeTDwE/6RWyL86h/rVblVRjygBLDYULv4LrFIvstLD5
6GSIt1hTbYckqNnvFsQ37w/Rcmm3AY6PLbNEGlsdvzxQIF8MsQdDifAKHparGlOWBSXtruzyvc5/
BH3KFnuscA1ivDi+FD9d5UMM1hdbxbWRb0JJa4D+lHBg0KVYqCE8OnKjqdvl9liWE4qcV50/Iy9m
nCFSLev+5wUPD6sG/n6xquGx8rHj+cYxypY9dQxDZR9tny16XWGqwDSz+1J6JxX/itonnbbARwij
HfypyfQLq0ZP7n4uFzVOe8USsSfsxq3xVJtQCysO6b3MrgHCbJsCbC7Oy7iluu+77G7MB542RwrN
/o6X2KlrQOuDkIAcBRiJ2sI2rYf5Osh9OL6i29ug7ZjHAV1U6OZJYyR73HC9inPN0x04v8jaeqyo
bI9al9BXb1E56ZaZ9gVXaFUyio19hZgAvmPonFORku3qEPOUb2IlE63TdhgfrBnAmquvwyMUcTOb
+Vpm0G+NUVMiofUmt0HH4Zk9PdDhrOIyFwyUBd8QF3fV++TS1Vp8TXCN1/nH/qjP167V6WVWKMdR
fHL+E1ce/RCE3hENMWJcOQHzl7Fp827J9Y5B4rlu7tbUcNHz8UeGN6lMsBQWbKkPZrisSCwjGOOa
bUzo2ZXU5eejKD6kr5me9xfIozzbtYxgQvadm6PX6jvXC668Z7BknLRZuVckE2pDgHL3fZwe+VsU
8tK6EPOJNtHTdQxLpnXAAHZCauiPJUnoIoKG4JWlZfeNjeG88u+Q80LB3/Tjq7kU5KGB2AlGbWHp
6X2/El5aCSVWRQ2DQ5o2sDxGTf8e/93WEnxyf/FI1bXruIws3v4lMHFvdqSioM5CR/R535Gjj03T
zbUdRmXS1GG89COeYGXwWLKubAXY77iQfm73DOWdcDGuCtLGjbvPWXJdVsnozflNWGcUXk4xgCcn
jnaBgnyx3+WKiMLMeoy7NXHJ2MFbW438P1HKsVgQ+TRUQ1yiwxHlcmXTbemug5lo8WqaZ8qO3NPj
UH90nuaHWAAnoP/7jN5r5WdiPE3Fd53IAybQUg39UfTmYUChjghOyk8R4JjAihN1B6UitJgUv0o7
rU6ZFEroi2uyj2qsnQLwA/iegePSnx1Cs3yjpOhylQlQYstIeoxsmu+nly0w5BnktdNMQLQqIuUP
OTaRnMIlmmpL7M79Wh8SoKkzbuhsRKaPFViQtDVvFyYR5nn73/PdQaqgLulbuFedaF4f6ATBhTri
I4EU0JAzYMhzvhDKUAuP1/nIh13oH3YNlVNEDunNshe7WZIHxwMMQE7lAVwfi+1CM5A8Sj4g0TXF
GSQakh+rmgKEuanUYlMcVcVTnMZB7TTDtZbC3xBMcjuxZ3VewuvbwEz5m46ABiG2kuRaS3CMOeCn
hH1QnJ7EG59Mer8rob2XKAqoPI/8/C0fZPUT+fnsBLKsQMMhEKTjiazNC6uJdIwSDEMqs+Nas/VN
VF0T9b51wTAqIGGKL8XwzXBD6b6m88h9dMMJ7rLJ/pEOMTnfIuHYktlt6xzGXkThFclQEJRY29u5
2bnMDeT6ar51ViYxO91JKZybyqMdJwK6t/jHM5RMrpp12jkDdlgipZ7F2ATiFOBK1AhWgMMmSw8W
bk4pyIVRCKIOds08dH4rTthDYtQHECq7/0h5436nOEMxpw5mmbc2obmUTbXjny3kC6UzHoNTNdRp
+1M1N025B6CiFsR2+TNnGGPtF1GDHlIokh8bf8kxYgFYxAZ77Ly/p9GNqm1Z6bEHYTzJtVytoats
XyGXncr4cbMBgqFiX8s4IJCI0Ub36l/F7oqKM0gGYMIXeZwdstk3FgrvWbuqFI5Jxij9DRZscquC
BsQlaJKxGWcCEO33OxJt4MmMvji0uR9piSE7Js+PyfWLWDuRYVFeJ+tRihvObe6Qcgn3eNjjpE3J
eew4FfJqczRaIRHd9JJuUThQlUuhn3lWgxD9qHqJp9ROa07Lmrr610MACwXdYL1VK/kwgqipBq/s
i2Mp6VIYPFIIVW+828S0E7A2KM25oLdCWPInNb2VYODdjnYWoYjC3vztLxZVwvHbMwlr7pG5ILzP
MeDOC1ySii+H7/t2+DB/kV6+GJwGmBk3CjuH9ToWYc2H4SRsF/vRKniCLwuXJqJrZcEICxQJoYPG
PB2WKEPHXj2Hz5PTfCk0b9HIttmV05rYB8fGIDoMS5+s+PnYT/FHQ/KSkMKABhgfZvWmEQDg6OV2
79dRxs21bpGSkGz3yLafRRkiY0ZFjYcKGxkF/Q6cK44wBZOReiZv1eivTJb6u5+eVFyUCQx4tuCl
PR8SSP2KMSx6hsZSwfS/H8Y+C3T3PypfFRQ8esFGU1xoTKrvaNqyhi9XMZx821d6WTefmmktyoeY
3yraGTCPMlg6k9R0eNO1uPnrU0LERUe69zy6yuFByRf/QjIM334SIdjveCU2OBhOgWnwtdzdbJa7
rngZEq2usywAZ7CMVDD12MHyWT1SQYYlPfFUaUvzoM7jk8ma3QM06i7XjnilGuJJIZBek6BslQxt
It4LOlacv2H7P62szVcJprofDvQefs8EuIq9EwRNRWsQKMVD+whRJu3QtbIVmiYREJFkz88nwdXu
kT6K1jreRPaKIT9/t5V7qnld+wJ/iFUbWpQseoDntSTmpiWdxCU5+sdhVf7Wu712qE75n43Q/19N
OvFIHUNS69bQ9Wuwwgg1dkkI6EFgsF3eAO6UEmrF72vY03Sytsy57CQis9sPKgLk96FHIeFqNgSc
P6xaBtCX7nUcp6sVryXlahZCqqbTOepLeebzEo/CFQvn/iYJKIsENjPcwN7Jf9pcBdwnzpa3a3LU
CQiYwRrm6QEd4c53Jsb0PWOxg2K5m1a61cd55CDHwj0xSsZO982+HrIDrWAz+1UmXzdu9no8P/ck
WbsFLHhczvnmZeg+xMNHKGs04QWykj/12K+0lKplp7Z4g4uNjo6ALKO/5u7fMGMLmatdI9Oj4OMi
h6ehOgKgsMm5LVOKEBF/2cEfrqxZlCur2A1a0p5ZTdAZjYSHkymPT3IeR2u2fBuKCWH5aiDy9xcG
iZo0WBESAnJhxLqqcGYLbg+lOTzwMe8sixJjq+Mg7LXkYRzft6TXtHGbsDkz0+QDkwZMkaNuaxVC
WMMPOSy9oqDxs7nTTZBIIEsXBGBXFbb5xTDxDomTNE17dM9MNR/u6qLV5ahhu/noGI3TXvXvs/4/
6z4WP1jSgSvv9ZdH+VeiWYEPXkiOnJ75It4wjhEQHNob0itDQ9lOvHfw3+QnAbTuTdj4r9NfXP0U
c0TPoZjDXt8v9ZHmhuVUJYLd3ki/sSb3dpWuMAS64x/RmGJV0kNeMDrMcVbMqttw+oeqsLNMSmdN
evne0QvmPrfKruX0TagcsOcb7qGAy5363wnTEOjnsHaAaDcAJushBn/KmdPd//FhxW7N4L0z/1YD
jMtwpLdN9O6Z9S8Ydvoo5INTVsilZwrehpl+HRcvHW/9t8zDfvKf++55lV5PLXxt5MI/Ef1ktdQX
Jqlkmqv5RYlCphKn4Pme3wofKL0Z2pQXxFYeyf7pQKwE9tYFyXeOrtlX/FjFma69R+nmbGkaYnM+
nMAOxegqR76eid9W7hl2tD9fIQTivEhgN3rJb6XgI5R13Ld9NpJ6nbMiYAbGI9nePbOUnrfD7kAS
tQtDrl+iXcHmkL1oBS/Bbkzx4/WvkEQ2IDBfT/pCcC9vk3ZzFAfb7PUIggs6HzYEg1iEqJaceK8+
dXWw7Q5f3mO++A/gXXCtld4PWteT62TKxmkbtut1qt07p3mQ5jfsUIzo7RRNdbGrmXmD0d46BASj
U8vui6zbQRj9bu80YEBsHyQ26t7AF2FHoRnVFtAbv9s6RLc10qfrtPDP+di32yDcyy2zacqAGfSV
RQFl0XUJj3VhiVmOrthM6mCOrAbs12Ia6zgO54LZD+5WHzUGwZ07buPXaob98s9zIzwoW7cpGkIo
FfFOutak/b9vuf2nlbsNPU9AQTcQ9S/Q83CrWUSTVUU5Xj/D+kQM7hG+GcGGGMB5IliOnmo/LmPg
ZNIzVBbpQtQGdTxIl5nTkiTZLRaaGQ63DFwlD74g5E5l81iabaLrOhljzTM4+FzBi7mDLid4F3sY
0wYr+npRx/JrRlFA4ubgpbw9HVlMpr2P9e3c7/6UF82DKo18tC10tgt/LphcT/YfGBzzlwRke6TZ
2hMSnzu5P8Kk1LpK0XxwFPo20DYqjMGAJqj8uhX7IchueplGd4SUNDGy2uXNFAnxJRnVit2q1Gc+
zx7yDGvH9hndwjmWLWr8VuMyuUtP8SJ3g6Q79Its4Ez26yOfXoQFg0RsUEhHBbnlkiYSSmCVbDe9
MavyThh/xcppEqKjD5btVOLnIFdqlcmLCi1E4EA9i2y3aDOmYuPXRLPI8dS+GARvNlaZedf60dLp
wJQeXIIZyqcifjt3vRfnKXUuX0+rECR2uUMzn5b+Sy4ObrQxKgdNzGer4ZsSEqZhhz3PI4AZaNNo
AbdUVmm7efJsxKKLAWCd64cEvhIXDU5Kust3pMb+7npq6CTvtwf/xVkoepWDv7FQTczDZZkbSSoQ
kV2PiF7CiiHo3vjV4LbEdpv9WWOyEiahnG2Xq3ndz65bQc4t7h0aHlz1gV1CQBmB6icktCWQJegt
GbV52R0HRNT2K37Cx9jjvUz5Fii7N029uANuKhffRKBBGrc7xXiJqs2RpXG75wiPgy+muD2ito+j
1KwybJsxc+1JAEeTBiHKotVYHGreB72lxqWeGKR4THvkrLrZ0pmNSVXGA/txB+RZex6dVNlde5jJ
NueTf+99KnxH1RRKR8YXyKOBNEotBUi3I1p7n17EcR2ExOPxVvg0WXJM2Cn+LiCiclYbc2BmPbMM
MYF2pEP1SaaupJLKycw/aeXeRe+JSocQdd43rtxgcyFlzv1VljBwAW3vHqaObnqQ8sntHCoB9Gps
xLcyi6XvnbX2phf1MVQ1gsFfQ+OBowEYv8FGcxogcOe96bBpXkGjKAe7iqfK8nQl5x11qaRYl1rU
GtKZ8VDnqRJscqG2D9LRmDSy8TkuQ8awPeBrcINnnDBtvHvJ+KKqwDdB+5IB1MNm+ENgMEWJ+a7e
JwRGfyj40+cc66iQRvL8+jFoCauMTMWUL5EdON6M8SSEQ+21GQYBwVwGqcUygTVxz9s5e97wBEm4
ypldCzj8IXvo3NMYY+uGHy39mvTphgZXnOcplEfOSX54r9k88UcbreB28OazZQiPpDwBTRPNdSBV
8JMlg46a+vmRNLhynhaq+1JPu3WdiJpRoFJ/gz5NuwMW+LTD5cV5DNLSB570nfc91bR1qO81CVc2
YhIY2HrjHBnB2QYvvLSEk1ijkZ7eeLCT+cJvJYZs8NHgL54hRj2i/HkJSZxSRYW1usHWbZE/AprA
MQKoB7kdHjPE7lmiAzfwajZno725EysytMqFy6izGePhSSbSxZHjIVflMsd+kJLAFjk/ow1Pr4lg
5P2P/6WqcRKZlc8Ilb0ywY95tYyNaT4XYRYcKPUCizjgC5KQ5uWtc9Osw3UQsqzKov2kaNL+7ixp
v1kJ8Ip34tdtxrZWxfZyLd5j4Qm9KIndIsqwI7V4/HF1S1YCjDwt7l68NUIRDtYlTVguKuPlD7o8
kl9RixyKODiJXkUzOmI9NMr8O83vkq7TmfB33pg93bPfBRd4NixkI8PenDE/BqQvyT8yLh4bwZP0
rvm7m2bDIRb8rbIQk5GaqkbjMAGxabjv6p+WFJKlnN2FEbwpbDV5uZqeJsUGQv1MXu+UgV2KfDE5
Ix+manVa1cbcN0s3H9xG2bulUlgeuzzuCIbF2wnsxWyRkzWooRdsHJ9r9fqgnjQM2l4bw+5Lokxn
REBVz0VapPfSIcLR77MFaygZE0qa9ya9UScuoQYL5FvB59GD+l6d9a1rN5Ulvd+QiRtBkb4dTYe2
1QqnxIaGyOMxDAz0CgClx84+PlSGjMQGRMGxJaYbeD8IgWlvm4HmzCDK0SOD9172nmyFvTewObWk
vZ5iQ9cfuxyeNEi0ALEl91TqL1hrstHC30sfEBlPgr6y9zQQ2ezmZtX/tkdR4WhEKnNs0wqLf2hY
qS+/SNcMBdBA/+6OiN7tGJlfYjTXh97AHmC3mUMljuBcS6qXbyPxuSg23HH9+/rnIR4hqoYm5mOH
aa52/lgeLj/Rxu4Sl0k0uXcfdxckO4WvKPZkyZwFXsf8O332xpQ+yJBAmVnQSt5esn8yrAk5L8NT
fMkaQ1IQrEuIalym2j8Hgome8iKees7KQ85OQQks55uE+t97StLqXrbKq3KGiEpkErNcFsNzo5Rg
dbiNo6+EW96HSeLndkYgpPoVirbAOIzaJ4Nr873DTHKtORkIJtjZPWX3jGEUwAInMx3MTOul6dd5
n33VcPXb/Cfui3Aj/nOJ4VQp0OXB+LRujwrjEQfNSXIfAOzGYixXc8EvRbaQBHf7N3XC73fnkJA8
MVAs6xBu/AsPoFIvY6lOeGMtlG3HzR6gCzQdK9hOW2rrW5O5QFhbzz3+VYL3ltepwGaHgNcYuxm6
vahCz7m+a2xPvhKfANCRwAqLFM05GSHbHmAQSGZsVSTQzT2KT0xj3wLBKjYHUtxk9zGIFtwRR1DE
Nw73WAqPu/xLBFlc2QDRoVnzOSQH5oiNBlOsmnV7oNJJm1pwsvZf52KvuSe4VelcrgwDOcLazkHI
DkwJGL7z6AZ+F/RbGxZR+x2G7ovvqZeeHqVLoAjXoceAWxMnJ4aSlitIEIkMZ2FpiY9OIIWfDPfB
zzYeJQsWbq6EMCKzxahGTboH9L11d8buZptbOfghaQMjpvcx3DYuuOY4WQ3oNwytamPE5h9NOapr
+CKBWHOYh5ug40EU+P5jbstOMwisPKH9j6XqEt5hPXENbansgArNp65NFutIAcRkVHwIpzIiiQto
s81UOnoe8Flgs55nicBrN6P0I9tg2SYOQBDuVej5MBEY1HV6YLJcxNUODYb1HbYgGJCFZZ6o9Vz9
aFBWqkEPh+yOONdc23hRC+9z6YH3Vi9wiLA2KXfTyraB3Pcg9kmbeX96sqBIVh7YafHLxvkFPBkq
MT6gJGxyWH4qF0kBUfvwqbj1rrTKZ5nRgxOjset+vx1Dy4gleYRTkFsQE7WjfvugEAJ3FwZXbCOd
OJQyckglr5MdJC3ZM8z88c2k/usc7fUBk9pzG9J6FFExhCHD3mLUnHWufacbfMcT9Sj1035XRdmf
GC3al7LPYV5gdaLBFL5vjEgk68lSEmuXjKIPQPnLTCufoxI++BvAIidgYOMALh9OmdhTB0Pr2szC
PGtfdkUOpT/UbWosrltfODMqnlwihpfaZomjSIBQURDi91tli7AavxO5dQP38Aldc1VGqEvWwGZB
tSZf3Cuf0VZ7SomJ7Ntr8s8l4xYz4XYOzG2k0oUOJcRKk79NJaIUdwM93f18/xRP7T1haQw31GAb
c9iznNPmaeVpvFWoRkvnKYoEi69aVbHIoMpHGDyNmOQ3qDZZAqcKZipt1lxYHfVgICWx2+LcqIQb
pZeFsRtFpy6UmgFhgbDCjU4bRJabFwLlNZ51LWMSq5cGgQFFrn0aECRN3irC/ohQX4w2PtokHyAf
+TE8NUtCVNuf7bK5ypvhD6pm5C7LlGIceu/dUoo1q1iPu8oAbFIXTuEOafMzU7KxkA9EGWvpCYcm
LgwQtVvj4+1pN+eTY/+hDCyZQvvvmIqJdj8xPrSOd2L6aEz1DJoxfLlz9TpU2QzDMXccehEw3/VH
1sy2T8IGBl/P6BalIfxKAUz5dZ3z6in5Qcd015YZXwlRxBPn+ghlkuwqTWJ2+y/H8A05zYqTu8Q4
Un3LkEYIyVHZYzyI41Ovu5VDV6H3qehLBzf2oCGqxtUh0sUWWe/P8qeeatQLyaPSf2ZqL8PhI1oe
RcNJjuZoShF/0+uQUyqELh0avQmc+CBVK+IkkVSPljUA4bbEYW8CjgvgDHaBH7ugCgUxDF1ifGfW
2MMk0hZk9LOjg5GGaTkmr7WRDDzGjG9yXzd4g2/vJN0In4j5+xR9cAB7bxnLVOOvLiRZ9NlhlJUE
GlbSeiYYlxNB4sQG4n0vLJpndmdxcorhPt+z1RZPFahk5C91Xy7TAdLslf4QidHOKBSGPuUFDTlJ
h0dmXgHVgO3zkU6Y5nMMWXRMChu5YcUS1a/ugjXU9y04sBcCzlsY988+hRqScDHrg2f04U3gjd2k
JiO0W7iNujJh4CQnFH3fuHcXlcAKrapKc0tHNmYRSb3Jjy0ciZH/zm47Nwed3qLyE8SZ9NjfNzWn
9/pWVzOycXNUT9+yvVp2tOrXhuatAGkyktgVm0VxutJeBTeMECmgcF/pVVHe8mk+0evPWLL9Uc1i
zjyJhL0qT8cJqkSECCbGWxXXfKaiHX8CLlTf3LhQEutOMHtzmlJbIPILBh3yJVnwz+a/IokHCxRy
XLwvvIQ2rlV6K5Iz1MlKxQRGc5hoiRRB33FFw/2aGqwghjQaYjM8cP1Pf0d5E7E2HfrQtd+R3qYo
s/rtnXzNyRV0AKMlXaXFc13taM4cmBdMIeYYTEce4v8usNAlynbjCdVv/daSUA1qtsHtswfggmnN
i6KjdoUMYLK7WWIwKthjGWevvQdef+FIzEs+zOc3UutYqrkA8dTpvkt4aVVZuF0LzOiL84CkeeBb
2VdJyzkIzf6NaOQxco1hCU6k+JklwZUMTEEHwqbM0LnYXk4Re5hnjm80LQIpyeFL1Wgc8zLoVyKl
OThUwMVYQt7kI2Hba753SM5UiiFnS03P97vAUEK8I6MlJzE8YoDxFUKUS8xIUod6FQZv0RFlLT0l
O0/BLNWzZiaetvmkTALWfEX4jQjdycDpZTe6MQHSqhu2wbI9Zp7L2uAy/B+Rn5U/c6YnlqGJXvx8
iJVrCkGVYH+qWkSWBzfAG5lN1m757tmWLiwx5ixGC8dj/JYD/BRCD0C3H6wOUNViac/724uFb9Ff
XbfSiErMJFbaYvwp5gPQfrpJQ2Gai7cmHrPu6h9RMLuwRD8qYcUerijJfbSZp1Ayf8hckSCqLoRH
TcgP3sDqm+oS+QbR0RpmtqAGYQwNPdVTbfu5wEEPgAs4wJPyGgn0/ldHy2v/lYnaCReN9UpNmCd6
V6Wcc/Gl5OJpjeC9zMFCqpNIWhOoYkC702ATamuBSsRcT8nF0Qk4SupQYD1J/9/oOAdIijBn/xPa
IATgVXPJdQRPlRhzl2qUUVZDQuMkoZlfw+DLWS+vvNr1pdMb3hyShnSN0oVdh816wo29tP2np/94
tuibNX6YfaVWOyguD0AG/+xWDf0UHSPl7TVB/2luwK0XoEkb26dC4r3onBNJKkPG+pWZCqm1SHLm
tprhkhrVKjQo8tID1nSsvKSEWaVGC6iqBS6D+0hj0HOVcs/oR76nL0bian2yx/5F31txh1gXzdBN
pF41kBU02xYJ/a/JakVFN73+DGw4ek25N/qDC+BAWQQQzp0Y5QgvIY7461hO676fPSKhf2DfrW+O
X8i0kvYG15xxJAauHUHkX3lB1JrHvViGwtlKXQeo96zxWTMl93QM3FCjssEkVEiZUU+T1qAhqQy6
6dYD8HZcHP1YPRFWosv1bBum+TIVlXrjUDBLzy92QkX3fHQ+KOzLGur2z3tjXdrkBiXt81QAXcnV
s2DXqjL9Vw4chwWwDlDbvn0LZ/g9FJJks3HMCHHogpa5y7s4m0/epvNEdPjBS4iyuPZH6PuHGccH
/39qThxS6KTELiJQ9aCxfyKqJytzwDjFmJ95WsPdSZi+K3CccC489W/0SFGx8HjQvBtZgzP6aPhZ
Zqf1DZZCGbaSNAloItePVT2rjP98/ueyYDC005l5N65Eq40PFHSSHUucXjYakQNOaC88zWlKAZ42
rbSpnHtDwNWpreD5uodMi3R4M31B/WCyPO2QHR0kn00uU/KnM8sh+kwg2632eAsMqKys3G58ud9k
gGGoEJ/G/fIwtyhOQrUjLJ8L0zHT/ioItev2QF9DtLuiMCG2pkTdxHzaSjyS8ZCCXCy0quByNDbI
P6dMN2Urj/145xOjwbBpElLtRwD2QNsolIOXjaQZN62Yk/k4tZTul/W6rUq7T9XzPE6UnTzk7mOL
/dXbf3JT7aXpqJs5k6gaHuedowWiVi+wDYSNOXQyL5LS4gf785otTJGnGtM6x4lOChwtod1GP5rk
F2sbw4qatmJ8qbSe7Db77iF+7jWLLkQNVunqL9RscOfCy0D52NDzm1PTvOBE5l8DPZ7rB3LG58Qn
KbR5WzBu378aJmUfw9I/3S6ijw7BGcaGt1/QQ1TGNcAWuC+0/iZ7GKmOKcUbGjvqhkV/NSeEdpgh
Qeow7VyZvMZ44dUjU2v2TKoudLaUwLs9djnM25kKuIUm0qvSmUWsDcLK2BdwQ3ZpfkFHMuNZ2nHX
B0Nq9YyAfvtZPG7kdy9FqkocbB6u1C2M7izEAWSvvmVz8KfuBZkvJ4iostw4Vtkx9F8wXH+8Kqnt
NepFLJkep+4FGj5V+oNAdhtPffLtMG1V5ezC/pt/u9xYVGZkYbcPs0xqRsyd3bxBbgTnGq8997jD
YOiuWGKVlyGtIGCPsa0ZgR8O6NBnyHKlHy0FgwVsY7zTY3vKS/CQeJaeqWEvWNhxjGhMF4Ynjgjw
N2YlGH6oVcJqM/GIZN2O7tVkVHFyjhYxMKO8ZGa1GRJHsCe6HPujTJtCZdksUUanT6VKiuozbYUq
QS+xIOx3wx3fOUs0OZ9u+9ySszrxZz42/BpU1TOKkaG9SrRZiPJgmcKji70WCXdbjNP88XBoYAhA
s+0VdSlm0cn3WHgGrSON/a1hQ8SbhX0bpRldp/cm9xPTS60KwTZhBcjqzquWvFKRU3xzTH/PbL6D
TdhfbTHJVgm8Bi0Gei0TONeYlyUinC7xi0kqvVHOMIthlU+woxhWJ7oFFdxjweMd7vxioX/oJLtb
uYQulQ461LAvqZLa78QSmM5rkVJNNujHZCNRkPG2oGNW2N8s0u9hgGgB/d4Qprgmm28mlhmLFxjn
25hlCvtTPGa4W//5uNybjP+4AaAnoVtZqZe3/95LYsbysczFWNzLXBGKrN5QNqXdTS0dsH2VNlWB
irQCngp0pE9XE6hzZDChYjosGVRq09hUYSk+CSS7Jli9BfIrVM4IQYKcToRelFB5QCATXNn41Tnx
qlVwwU/7C7jdriYKO1rJv9vFV1wzOYH5lfCVbuEGC14VhvolGQeSsvz7Eu59JyxjBScH0w1mQv8w
c34/wFXJAFKNUI3QvUhaGh3vqtN4u8IkLQ0XBKzBQ73hbLoQIhuW8npKAoVSRJmwyd5pf4vzlJod
BgZr2th15VBIx/I55wTjgI2r+mY92QsT7MSINJoqhmjhXeFpF0p91lTtvRFgzQZ8nWzk219pk6rj
qGjUgeWFr+7/5ewa5CERcec+h0JiMZ6CsV9VCR//cdoY0n57TaYXDmn7A87EJXrc67U2Frj+Lksm
543s0vz+m7WK5rNn6czunNQs7bU54haNBP0gwVN9cv7kVQGywUqAoR6p9CMIGy6yZahQBMzWnkkJ
A84WfwzRnWVHLBijKlHFoCL3ufQ/Jtk939acShbWFk11qLbBuwwJshXe6Y0eubkKC2ngSxKWYCGd
qRuRdYe1l6adoVAUNNRSDquQkYJqYt1E+au5ws2pC2aJSWpJZgk35WAfpy1VurTvtqqh9uJ2ImVj
TTBChbPchDKgfO233yJkqkNI0/gzbm1hrbFyOqB55a9fvB0uGXqCmXhVkoAfqbcMEr+LosheL5J1
6xRAyrbGCfaQpBsHPDlVFoBPtrsKXMXWZdzHnpQJ8FdaFMC3DQSEH+D3JVAo3tXFZqtVIiMUbuu6
lymTjvp92xeciAquZzCMawGjYds28U0xdoZXlMv28OsRsO3RZDSpWeHbeSmNp+7/UsJjBwC1RcTg
AoWryUmH7jV8jN0wgJMUA+AdqtIMNj9sBapRRcBKc4TD4/YO9l7iYIztgmfW5Q/eQhcpV9O4Ob9X
wsEkHz3oDS9K/SfZE+mTlDH4VPc0cMNHdJZ6Sqj748wQZNTyXys/kgav2+X5XfiMqKydRnOv2Pb5
MYQphy+zR+5Nz8lN0I/n/kygLa4Jw/iSGS6GcnLGkDTBIFnLzxUHsJDcFNkYOFIIsNoTTN7bEFrR
J11DHdMEfb16h4IqDk2GJgRDKCcEmy6iVAxBqVSU+lMvTPKgj7w/tiUEmQvmgCslUEQFgkTwa/Me
RV6bf/U3V8ZfCQATLPEEq25QdBwcdgWLyKp8eGdfaHBTs5SPL4huMEZVvwEEWUhr6RWHBIv186Xc
xaRppBIWJfgr++gYcjYN7e0bPNxkLLThxRgF5kJHdlxkTOrPAnA7oa4BmLXb2WdGfbThCoPP44Sp
ECb3aBUJhmH7PrzWg4+6SqCBCWm3+3B8rQhASHMk/1yruXweylL4Ej4EXNW4fDxYVTkG6aSzwFuY
xMdbc9ggRrIb2+vz5GkgqFH+iGDheOJijBugJ65k3FqzfecDkTwV5g0gGZJ+WZ9E/op5bynkxN3C
794AZWAyxQfjso+whhLTy0AQxDUis7+2DmYuSKaBcaSzKgoHDt9TB4y5ruitIAfN8wUW8nfVGeaa
eGTjI/Jtzvn1Z/IowYRdbtDk7KL2GLFYp34bNMp/N2BWxRhIjpL8tyi9tojkf2HohGL4pi1J847l
vKxxdKvesN5J9+oxe9trjSiej8mgJlhrZIB4LsDBZMXi76uhEKydW/eR+tHhytea4xn2D9gwv2BK
CbTNMe+5jRWMvkMwWsIKkraHv7D79mT/4QHRMA7Hfq4FLEaRKJLRdn95uzjjk9lNucSHbjIrePNk
61wpTczkgolrrMbCikMQyN2dc1EkzOjFHnLmAeeXm3URQigxlYU41JKBPngcLJu/n0VxQ09wm1Em
64xHkp03pnvD5iHP82XxNcfNl0nVzMD6h+40xMpAWqgYHiTr3WX8YrfRPx+oEhGf5gaPHQF1249d
voYEqODwAE4/TsOCsxdhNpqABhwUwgbjmT+5HXJdDmU2i91YcquLXIrJj6qKIpv8eZm5Vei8Hshh
SU0auLEFM6ePsAdjb50A4Wrxp15kEdLF7ZY63AqGxlsiqGhYX2oTbAypW5U3rcRk7UXswcFfvbdw
wwZcPOUZ369hBR3T1uC7SIETL9KM9CxcAYe+4SMC+XzWSCKBkPtTJYZHkDDtCF/A0b9dPCtkB02l
qE9CHJZHa0ZweXOArF0mHswUrbWUYEreIorVBkbEBWaTzG0pC4X6vnAlGt/w9JplzhNoFVqM9oPS
wc9HI6dsWycsF/diAYKJGUrMjE+RyA2eRKynkeztMQ35zFyllWSHCviUjF9zC3UmIpovRTYC0tfX
uczbt/CUyQ36NOGy5zixAcwefy1bRaKOr3wv1v4Az8Mx+CI5wcCo4mDA9lfQDcRzNdCKwhGvQEe4
tFnTUhp0Ow+ywd33QfLfs0pvLxNamwcswJW/hhnyGU8qJfgnYmBDnC855pYgXWXpu8j0rYXCpmz+
OOpAj3yYi6EZkUzCnVwNq7fEYN+2zRcQx+ap25+ebmRF1Zptdc8xi8XtPK2ZRn1zyKzF9zoFqLvy
x3iIVl09gx3iID2A298lFBM4yCg+QQf5d31VH+WA++NAeZExFMVP3oQcOYX1EKymM48B1McKZ++/
FAib2Sq0JP0Se5+JpMzABroAsorcR6bUs8oOW57eM8UhVV9dtVG5h0nMvk4x/MrMZkIrtbhZzv1b
b0Xl6U/6jtgwl3vLNZX/4pdJHnOdcr72jcu54O6vaNg5BJoPW5LXoNYy3ZuOwGEYcZKEeISmElFZ
fccQcDVo87Q39KVJtBbJrabzQ5Z0lVs7e9lOrs8SKBP3Z/ahHN9vNaqy6UU/fq3CEBYVbnAn/SG7
HbTYth4xwPQo0CtgQAneFRMLRWZyBnuOxNyeErE5efwJbov9l/3F0ENrOUuq/ZX0NuOd3Zon/l1k
RheyJvshLfntfQ4fs1x7VfS8BCxPXqC/613lyhNqLBSHT4yiS9MrxK56/Cplv3J4ixRVbQGq8hRK
YKYHJ4Whci0aHNw7mQoqgGahgM79GwyYYF4mLm1/ImOw9/7YQYy01DJ0abv0uB5/SSRR7QMRCW+b
9O5gaRNyzX1MfnlRYF3rydOd7dI0dgS8Dzo3FSKiCrxG9fCaVCgdbf9vz49+lSsoOgPE0Bl/Ydfl
juh+9zh2yZVoNTnfyl62gcz081zwZ55ssSx/Ly5hwOcloYqsY1WbAUbrch6FNqJj6v0mxfRRon05
/OZz/0ii8rGkz2cj2epI6NWk3kCrTH8orYZZcTOFdeUpkeoGNuNA4xlpYfKCcX0/jO5haQJ+CbWq
NUABoovkxL08uhYsSemwlvITed2lzMopijveAeixzUJssVIKVFBFdYGru9exaE7/QJtOu7tqFWFf
wRIhCul1bX0UGauG60hruegxIU//q4/LVmz2dYbRgdtyh8KnthnN+o3gpOnI6ODTWLtUVot4T9Np
2uoqKkozbuNLWxaoIBffyj5GdE2AY4U5iCoSHbDI3gQh2/Z/VaW9uxKINScxxwiAyB2a4MHlK2tW
HNjqcpfmq/BuABOOorESJJtK2RBlt6R3qplrBBOcwbD7AjZf/G3KAZNkTcbthQSygymG1YENbWuK
leoijGlDCw/f08bftnVrCXGzQqfRriPO3GIgIfif729BKUpjJS/SA9vVLbYsUNCzCdj/gw9tC9jT
LrMUW8JnVsXqt9cxKKi1nCh7L25RNkprLk3rH/FJPDX15Tfeqk+UfA79VeBu58Jx8n182Gzq039Z
DRcqyuhM7Mj9LuHY3RRGzj7izPNw3cARuREejOGVlM9rbYamt2//hPK61NtueKIz2JnPpuG+gp8n
wykSwsHkoaoTGEJBLwtQolE1tkw647OgbXBf3wt/XjqkLyKd6VBwsuU2l+6B0r8lrraJKpStkzQl
IDP35bBFjzeDLesYZp5Iez/9BoMLVPz75SmVhTlpW/ESu5Qfkxcd9e93QmP4I8vy0zjMtKiVCC/G
00xLlzySp988dcfdCIgX/0i4GSKarJnsAe/39XFsnjf+rEVzEHEwaA7TxYC4ho0vLjDuB3JV2rK2
kXgMB4eO+OCPsMMb7mzse+3PwtX+bjObbs7WJxBWzc3jcr25AoL4djanbBOuyru81S/m59v9s20t
iOsVruC8rZmuUgdURva5oFtx3WC5TXtsm3DFU/9KhpPxr+udXsISQ/+7S5ZvtXkpJMxjZpnOKb0v
ZHMLtPbOSJkdUXSpVgSLA7XfbQehBDgR6BXqB5/J0K3f5E03p6eZtpRZvCdaeD8fyF9523onTR+f
+vPU+ice6elNK3BOcwkq3U5JxCWyup5BcFi2gqKa4Bs3fDjE3y7vxO7FpS+QPrAMrHlqCxqBqIXH
4vdTHmvgtlHLRZOYztViYQRDsz2GPHjoVxVqjOwhxTob42WehvbycOmwnoP+4ozR6bDAZXVZ9VxZ
h/Fr/naJMXld3JD6xjx8tv514GlrVUJVV/P/yUot+Q8pcx7Ukx6xx5EsENJObGxVUosMkHOYcV6e
hG/KuUe8jrZx6r0S1tQzAUKfvIY1lOVpGWIOnNodvVCImodzo1eeCPpe+WPc3fpupNHULhAQmj8y
Ki7jzjdiSjA6J2H2J9yspbhDa2Ld0MAumO7K/svTfv1SrG7YUI6Z+tIE1FFX0vS8drDZfguqRYvj
MhWhyjShiEgfEIstO11xs8xO2639zCyOsf4SCsOSAjGK65zoJflUUfEZ+3GYzJCQ/imVi+AteJ9d
m/nLQF50LSGnDsMiX7MMtM2XMCOGnZ9lbpxwpXycozKhaR2GmFYCdA1YxdsFLDzq3NqOF8RB9s2I
Ft/fl6cq+MCw/hbbIYPkTl1AUU0PkthPluSnEflqzC1EymC5NHVWEvEn8exykPwj1/iCkIekVw8z
jyaLr+qlxzWrauKvpwVW7cyIwzilL82N/8GqO8EyIu2KRONTFPeU9tn8yWEa//ZuWt5RBpxZ+1Fa
X6OGehIDwt3JtpD3bdptf3csF8MJ7hM/QfT/SZ2GNLQO6wrkT0BM4jxa2O4/d3mArmwh12WGOuUO
izNssJ1GEJ2r5ErohoW7un/KRsnAFTy4Gntc88CoK7WT3SyRjyiau9h+YNiiyFMhicYKihW9q2k2
YqkvzBwkMehwfhrFcRHqc1+uJPPGG6S+Gty9/6zvjcpdg2YkB7oKgEPUV0BsEsXfzVyd/59dMhIL
fCppa4Y3D9jtcD0rx+xjYvCSdeN2PAx6BHAk4BQsz0RFlPrZdJswseemTrr8FaHbiJfoRIiEKqsv
62+0nZQ+afxYdhlDIFpIqza/6WlPVmd+7Wivqj3Qyz0G5D65Evq9J3LGWF7qEMtAEsb+hOJ7rYAR
A1U4iDR2JKaei0kt62fv1Ci0gl2F0VVWCrj9Hp5Pr+yAADqoBP1kE5/c5kxeWbH3MJfbm5HyC8Vn
qusuY7AMEjbG9vQPE3gMIan0APASAxoQaR06YoDS8qynD8Syep97ZA1t6u/AaQm2ima0HCl2mVNL
ZoY//f5hrYkfxrrE3CDPh+ufqPvgzuN7n9Yl5mUeuItuI+fLDhAq8ilphFrExyoJCJ0Ju3Su8UKN
BV5e0oCKoccnA2T+o/9EJG4zuiuCEyspJSMjmoe9Tp1xkYtiPNJ+GsH9f3/XLeT/JJ4DleVK/1FW
eKiNnW6mXDIy0M9cRJAZBgsGv2lqoVN+yHGGr4tED8hBm+jOZbIF6c/uf5yyDkkR9C2pk1yIa3se
6wgHmpvCCj5mHglMlgJIhzpLuBQ7yCkla5BnzSLyJ98vr9VvjTm9jFMOv719zMcCSosS+GJHDF+3
rOa/paS2gtfqMHXa4Z/7Ad6KpCix9xF6GnefnN7Hq6mD9UxXw3pBgnKlbTHMi+lHAF5xBwmYmg8R
1hQqxqXJP71GF8vmZ/jga/t3MLIuAPXIiuHTKzLLOO2SL8xSxRkZHluOczjtSX32UM6GBnnIiPMy
5g2r1dWg13I3ucnn1yh+Ve1rnKJlrZ82kVjo1tOi1cGvJjnCpVRCOYIJv6VETTiAu7W+dUbEZo38
NA7CglIjm4zDobGf1eLHneBTx4vproXi40a0YSyXCe4bwOYKPSDHDM4JQykau6FSKefSPR5Oh3R0
tn/W+gHCyFgoTj56A7ZqDJfaWDBCeE9ZdhlhHqKYIgS+JFGnXdS42aX8SbncvF9BGowQ3VdZw8Vn
WtiIx/GfglcTEKqzvqv6ESR8ewB0FYkQloiew6rLaU819Pf4w40mfk6TYNtFGjmtkZxYTUlu2ho2
+g5Vfw9Yy2Y82rdosA7/Os/yj6MmsB3YMtSuuuAmnoRWf3ZxWnLlUpFtxRUBoo/ptp4bDotnLrY9
+EM4uI/c8wJFGyWuAxfd5ZXYOkw+Zkb0eeLKl7YBjTNRBBTXC33VGCTQxtBZwKhlLwZtnpxDBNxe
3/wq3akNA8HKxIu6eozOOgHLpM/IO1ZagDUgD59rvgaKOpffwHH1MjvFZf+HKTJrWIAYq+OwNGHb
zrsTkaJVxB8zbshisjLCImu0ysNvHsOoL/jHct/cyza4dYmsN6MYb4md0qh7nuEFqZR5yWNamCLE
Y8i+E1wY8sn//jNEH3jobhTHs+2YoolGaa7sD2thOrTlnnqaD12LtvGLe0OFKL6n9Ndfve7gfKgW
KktUrj3fQ0onLY6o7fgK+VnxzpvjPgy3i/JA7ZANgx8vteaJKAG2c6Tv5EiHSrlKdwJsxWALdXjM
+7KfEoXCJ/5eSRhecrX575fdoR4AnE5KPf3sJdlAivsCjnoVmsIjbxQbU7cQNrK7QBaDlh/TwpaD
Ck1cYCe4MEPWby96gTivZj5ticZhWnzVPM7Qt6j9IPh4F3QjvNgZp5XLtGGqVPSkrXa+PgyPHImr
VavgQ3Pqbp7BwhUVmZyvUM2AXGgNv6jVQ1rRH2q9E89URZHbY1sQhZLBUKwIm+iYqjOClg8nZO+I
evlmgKPTkEKNjzWTT4gWQS3QKS+pv6aQdbdJdCWtRN4E/EpbsPmf8cTDP7OjMICuFdHscx9zQ9nE
geRd6pSpZJrekM4iZ18R+ld77i3xAlu35gZAP3cyr3lmQCpvPn4Ikrwskg6bG4KKKald610xhZDA
+9YiXoKuoWLKZtwH+jhlZaHztL5MqoQO1mStHTzz7tin4Iw7BNXNnmFK2419o8J6IsS8T+7ruHX2
lMoEXip45vtYfR20ZQ4Zr+5pSDS3h1uS8VubYmSOUILAmdHHgN+naSMhAKJBrZ/aztVhO53aA2fb
rYjVWt3BVn2p0sIIiDynTkzIZ7P39XjczD8wPVLV4fS1bCAA2Gao2eoNgUnZZuSkiDeYavTCMUSk
MVgk7zL7/6MprQikA9Rj48yFD7HxXr8OZlXaiNmUuAWLMqMsuPuBkCS1vNH1y1VBLtCfAHZZWSbW
5mRibhYX5Zz4SoGkDm2BZoKg2eFA0uCsBL/Vfa4RkWbyTGM2JaaJVh0sFyL6SzdwME3qvJL/taRX
VYCixUYd/wvC/nLsf8qHJVT3EBtFuG9Fuxx4g1OQ99Nmr/893y5IvWkIUYYBhV35Pdsp6isYOK3g
3XL0W7700Ei09Ma4oDj+M4OYRDx6oAIHD51igzPkmtt654nR/f9ByckAP+SXRPjeMF8EFDafhIOy
JXTI72TrHK3iLh2rDsBaH0ZMRQ8WwYzBejP6SRzyfo1Ls7y/HR8QJ+Zk4Sn/4JB5B8VnK/QNKw4h
5TMGVq3xNm7cjDIxstreZE1ss17PkKNfNl4ExdRYyiMgZ+hr+lnX620EsOyQkZElb9Ybfwv35pel
7T0jFoJAopGOD88sd2bW/bOvXpxf++xQwqn77dFgSMq3zoFPvLl3WNQM5Xumn2EfybpREk97kbTt
xTigO1r6LHqfSk6tQnqRdL3K+uMBSBJF3mWzaFsyYm88dlhCeOTEgrMJj2tDA0WMoXk8eaEI2Gld
UCpAoh4BHPQleQbrumAyiEg1RaQlJp6aw6UL/vSbH5hkf8amb/qsh50cCl9uWyd68dkduPN0/Uji
eHIXRcn9PZjelaJW5bONO+nelN0UO32OM7m1YgOIX5gqzn00AO1sIzP4Yk1wEcNPP/pysmYq9VUg
FYBTM8NgNBQgSXrksrowwZZpi72eBCb81n2DXtdy8eZlEjUCXxiU2T2ynJ8pSfdeoeK/d3H7Ald7
fILfhlBCvWzL9kvJ5ZjF2a6MNYGmmb7MZIwv41EJH7ggq/32auZ6FqLlzDfkOFShychGZzaJfDjt
3KkBQf6Ky6zWRn/duQgsmzTgkzW12/FqI7M9iw1bju0LYsSC7uexg6UMEv+yOn41hbpc6moi/TYo
Rk+RkFZXX9bKlXBHHHs6orL+xD3w4j9MeDtgCdRJFtT9wXMEywcraGZkv3xTM48bS060E1H4GhgO
wseXmo3/Sy2gRNz7CK4OiW3VZeeDXE8cD7vMN4WAzzNUtp/DOPjabLfUY/7LmUmfDsOuRNNXfxFk
KL9clKRXSsP0bIhLrkbIevqZuA9fN60sIRKLfniNy2j/g7oG/gX34jpOEdU5/EsuldQyJdfkHyLR
uOF2/ke5XVw3fIyv6h8qB0QpiJ1wgjQTRFeyGtiUFQpEfq5MrBYEL5CKqwrGaiD+C7+zCm6vFk90
F0nrMRWF2OcVTRBEiswJ1dhFdzw4JDvZ9LZfFwAgrn+QcW37Cem3VYELnBVg/x82yDLzOhFT4hx2
a8lOsBJfkqHFYogFdKO8TqEzJV6IPBWwy3Hs4Fkuk16GZd6zq1pYVoifdHMvHJdMgNaVtxLA5sUS
ecZ5cg9xvhwEn3XwigjCnRizD9BsO0W02nS5lwjABjeDD8TsjmZGTzIpefaMpr0yi0fVkpHNhLA3
aeztH+bRXNCwc9XNzH1y4+HrQwYqUp5/4fCoGLYh6NDmLv15YEZeiDucSdQFdQY8cjiUPEdN6eD3
KteP7donwmbT7BEjEKcwsR1zAWlCHJBr4mvGwHhcVL0583wjy5xOUsXE+yLIaazhbtC3DzigGiB5
a23/fhSwTPSNVvVFouSnxXlw1h/i2H849N0jxpg+hPCFpltwf0s/+yO2K5UOzSBiY9/yhW9d80Jh
mocfia7V3hq+FJUhAQBT7coEfD2G8oxoBcz6D+KCIKVR3f3jHXed7gP1rJT6VJ/xYck0IJ2hPIio
I0WNCEFXwI1JiPJZncFXIs5Wz8VsbYLGmP7ogVZNnoPGp/m5MoDwahjvsmo2SVTC3Qhf5nV+Cjc3
291BXuJm/I/MbyMl3RNN7JriPfL0gOVrSqHQC/ugXXM7zIsjjA6g2hyrKk2mjvr8htJGvavXGNJc
4DKWGgqFFoy+CtYQUnhzcKDsCauiC692kqqm/lqvwzv7o3DVkNe+QCDKirTz6xF5ncuvLV4kX8Aq
KCf/kBF55VACL8TS/IAp1N3GbEDaR7evWXnozmFaZQ/xmQCDIL7dnSPVhXddMaylg2lzwWpiRAtC
LLrOrCkZOLctMNfmKZV569KCI44ZSTelEFxrAqMYB1O45wXXKbMdS77RjoWVj9HLuis+cuSaqP+V
Fer728XSomEuLpTyESFI7rj1DVDsMvzsmiqjlVWZgi54M9qjsyRjENDGKD069Bve6l9XmE5vglcK
rkGvuf8p+6KvU94qMjrVmog8cPwTVOS27KDXmkwcKZtS+SbpoxEJiRJr22DSqoGdJEpEnuLCp3B2
9na42Q+zVq1H90xLUBkSU4AQQiSDDrGGmrH4sz24tws5lFEisJizklf3FhY4p0jCfSI4EEg0e+SJ
pUpn86dDYBHFAwIFDU2M0OqxVO/n/XCwmNBiyzNyogcCOiv795WYWiBkD0KIrIYuCMM1litlvcAl
a7fcmvOrzWlApEBZWAGYWxaOckQf2mHjlIpCxyHHhC1NT8FwkkEaMn2RB1Ml182rRSWdwGSmZLfJ
5+5Qmu1KSwzSm/X3Ok0k7v75kV7XGQoHX3SMrMmgM0c2c+6lHnx5O8RXKJ7MuKmrx7LG9V7AuzzO
sreVu6MnLJiZTXLwaR0ajmKCjPIKw+g3mHKkTobjb1lzKSlQnC9Q0rcaXRFmIHqeKO2bLhRRyqR4
YyVwCtb516cvwvTdz6m0eKLJtrx6Smkr99QK3U/51F5GGe7m1jmAxzUrXeZ33i5cRYRDbNMK7gyf
/H7c0s+BfsC44/s3+ceBRC/sxapKvYYtH6J7BITMvY7BJf9x0UoQqnvXOQgEP9CLrFr8Y7cA0+uC
Nqi9h0DosM9CTpw+1EXtvbo/6XD3mXP01nmq+xYhz2v9ql45Gn6qCKPw4ClfGnJW1QpPUCXEfRP1
2Kyr61gxhXgVEziSwHEY/EVVWdfKBHISapGRxH57e4FHlNIqKdJBuzm1GCn8XfGV/QP4HT9XuT2O
CcU2g1D3qNAj59Ha/8ehKrLEg1oeCRCt/PHxguyyUG+LE/scV4AYxdD5wmt7vZYX3XjNIj6A6b+e
fGTwBDv+nuT19Yt3dXIp1xQNixfuOJTpA/vu6MRTgVHueS8uT4LrHhu2rJnopxi/j8M9do4QEUTo
LCBJaaofQ/pa69GMKxsL6fLj6CMCTRihYtsT3Q6DLyk1zLo+L0nEM6VNNGZtzEskBzKBI8VWmwdl
Elfzq/xpn9w3hkAaKDjDN8DjwYK/GTf71YpohS5whBIZH8pRDVoqBGeO5d/sqefa+vWypg2TBftN
rxbfYTijvirrAa/RPRbe6kTfXbw/AdcP+H9J8mNynebvKYEAbrzOXcGJdBVThMvtIzTAkUEXJd9/
zZlF4jnnXxcFdgu9ybhIcw2BGdNkh6vve6vb+Yyy6o8ZWhK07dvBO8BUh0TZlHzHOq3EQjXC/kY/
af+fa/2Bbz9yqKx1YE5TiDOR8gKw5bmYu6k4sohRQB4vGNmCeJIpt9ze8nReyyYOwilUm+G10YGf
x9m2ZClXiXdO80zWAipBBUVksAI1jJuHhsRvspHbU9pKdfyip5oaUh90KWqxs7XAzQ/dmEgXq1Ke
K0JNXkvP18mhcNa4g9BQ69aeAzgBhUAFto0Z2esVFA2Ie2B83+5+N3m8lOEzwNLyKsGPrifKzz4A
lRr5LDA5TU8UF0AY/PfiskN4KvmVBZCfkkwiffv21F5KG2+fvR91jVHUMbNFsvzLkmeIiGsKExZy
q+VdNrS97YQ52GAzCF1gCGETffFIB85YeGEaLzyU5WDLdSJDAaUMmArC3HJxIG7VaipbnBIU3hfx
lDADiYRaWM58zwbMKXH2hq9lz68v94yR8P4jAPAuSDD/SZEsOCg7ktL1WThqA+k5GB/29ulU+HTk
vJv3NSAdgTYXooH5kOwCAArcJDj2qa4s5BRMnZFf6BgkoAazdVGCC306uI76K3ihdNnwScd2QDqI
58BfxqDmYePSEvlG0sHcgzj/s7E0MBKPgySQLZhVha+yGhnYa3s0EK6pP3ylKThE6CNEWH9zQhgI
z5Y8RORTGaFXNeJociaxa3Jx5Dqj0Dh6TWYn9qyVy2HNyUhk2oLBSGwykhC9BXqXCLp1FkaMtD7e
hW2/wykwbCvZ72z7qFHf0MHs5j9SZgGjyif4aPo3E7aMrl/va6fn1GzkGiIoSBugvOC8Du9E7tkg
TixhGF6R788BGSFdwymLLW89nWhans9/7U0ZSps/eRJYhcpwFEY7dj+AuQD12dP/UnUmcp+IXTUO
SwrGzflcAUpv/HJ3jwK9Wis7r/R88H3KGJYh05A3vpUdAyIidQ/YDdDZcSc4M1b/H6Up87oLorAh
Dy7LkbLFmINj/bZA7hLBCUEBhTd4yGw2Mov5JeUSJnPkpSfozrif85f/XHLhs3GuzY67V6GhSqGD
+cljd10TGuIH1n6fqmgPxvgeuf2Tj/iCtMT0JCJcrC9fLmJXVKlwUR5n6bqlvaqJWDqrXRohd7h0
6TLfwhET1WlVTCFeeq7E7YxkG0uXjzgptyZxxoNGuHle/e5MUESAJhw5oC3T60dGD2H0qS/dUBHi
NXfsco5eP3WA/p2KnV9AbmKP+hMgcuMHxbGD84MkTo2ShJEM4p1gnAG+gMqzEZqlCk2W8RxWkOzJ
JlS2mKmEL5q8y9pEaQL+Z6QWHkLzN1pUmPgDfiz4/k8GWNvpc4fBUrbJu0I97nKrXa9ETrSeAojm
Gh63h6bg6Bzpk6xp6DbHk7HEkukpFelVfXqHOIQ3AehZwPq8AcxqRkkHaki3nA8jnUCWtLikOLAA
67Lvnret0SwjlVIVM++i+KsjsffxfnVIkXZTjjX57YKjoRlHHsypB8mivLzbbI2OuXz4Tv/pxDPI
wUy58E1cvS16gjAEsDoAB50kjVVCLVcmWoRO1HyOzb8lCcMTg+ByURDjCUf2fm5t6w803vsUR8Ny
t4j9cRw0UxX1coIaayh8ZmR7yCWRpzO+a0wuc7cxxLt9Qln3YN0NYKOmn4SaLhv5a36rJCSYHury
xRmYwO/GL2jwJHe2o4Oanc8m1oiaOj9oNhoFXblVXtKh+fVmPEGGjH/4xVLDLAZxbH+iUJGplUY0
giGRcK4ppgsWt7GLyzk425XOto6p8Z6VSN4u+qI6b0arjSaxpN7uFam+5spd0eAYmGLzv/7YQRTO
6dZ4FVihRkGgvJM2bRbLZnRy2mNwjZL95+mGzOoDco7qGBL8/MvIVWL5OjNPkbOtVbZykCX66QEb
BcLV5UXHXItQ8M/CkP58oYwDdF0489+GTTcjpwhnIqAD4f80Q69516cEuvefRo30Jb4Gu6GVBWaA
ZL2edMSQl6wKQkOY9WnVzPteiCiIC7+T4vq/wydw08i+MgE1UpPV4lSOYaGlVi1UYGfPY4iHqh3U
wPCEQ276yNJZTg3oMdHKW8Mj0v4y9bj0petsaOR9A3FXbkMSIjeJ4QcY4qafLnaeZc4jZxZbVzoY
MOpFqGjwzkua5dSHRRetrCSrNQsc6t5+iEOaV/Ic3ZaH6RXCRaA/QrtqAIVFrJrlb1xNZtxv08b+
h4mhEBYR1xXo+GcodeNARx8A5IXoQXGqOFELrx+Qey/Fvdp3iFzmfWUhTnjeAq5Jve0vSHKtKkUZ
6HBqWVrdXjBNMAFFMMdgEw0cX1dsqJ1I34E6rfFb0KIfrj4LkfJkHKwWKRiwoOP4trcDwg9OhdUE
bRBFXX87Rhj7XFLvuOpAIt1WR00Yu8bYpN8hGSmexPJvbZ1FDCS0+cw1Zo8OTLU1Icxq1KGhHNlS
gNn4qrkADdsV+r96ehuMN5NILkBnWAM9dW6OBWaKZUokg76yPYIZ1dJnvlt6yuJ+ETwa8wBEkFxw
AbkGyKvLo+N2He4CTfDsGxiXh/1DN3ppNMNWqzDzNn4JmU+6CYkJ9iIZWMBl1iUICTrg1xwa1I+a
8+nw95e+TmvGVnjyyz/U9fUj1U2VI7sQWU2Pjgr6Gdt1f7qTpTNpMkl8K4kxKmdhaOYs1INQA9AD
oIk8JJLMpfAfow3kudMe2ZWUxpSdNNmDrrzgbtwIQgluVwZvrhCy+Ib2JzmXKwzyDDNIFFrGVZou
CgztMoqoeiviW6YHdooU5JxvVewIE+hUL/vPuE4EpDrcGxAxvcxPqPN+pYLzRcry0o1y732bOaID
azyIPVOPsVexo+/VWtvfgdOJXJ+a0cwB7o5ENWagHP39wM9erOK31ezRiU67k2HDOfFP3+KnCf80
BeIW2A2dfkgNTA4b4ybJlQPxh6zyHqnue513NGfUe2aUFKBSc3UziY4icg9P8TAxaI84wCfsf/tm
TQTBRgvEzYgJcGe5rOXfL9ctdnv65pqstkpHlnrQmp7Wo/wsEStGhYksTuuyTWaBosnDYSL898hX
n4JmAJ5GOdIE6It4PZA1ApR/ArGFlw6CuXZobohJuHzYsixHB9g2X4/Vngjpu/TT1664C/6lhoTA
tXsUHcIZqXAtJFo62dq5NT4rfYhhHhfI5cNoucbA3dbkfEIkuR2+Ss3yy33TanSXV/L5cNyHIEZ7
xzOwOe0nW5dfMSFdJMdx3YF/KevfT+9q7buXamKbZF168pOHlpPQBB9Qu+1by3LYWomVUta80rQT
wlqFdsAB0oo7XoB7LUI+Nk3rf13pUEE1weTvYfS7K65ACcg2vWWKaqrxmAzos0hmRxa62SxrJ41w
rDZPDgkakLLdPBTNb8osTl7SPyGOBqDyqD4VS0bzlGWG5CfPRS5lO2SOGmxx6a5mkf5coEHQek7q
KhG6w7Aw5AEhS4+VB3ueaWtNgq2oYmQSNQkMG2P2pB9SsluuIF5ZfVn/ozTMgnE5XCbLNIUQvjU6
rLowyr0VExki25k7gcOm8tgP6WJVIZ/eJZNqD22IWbD5VnSs+O5aGfmU6GDzDpRsdR+iH0PpNUrj
lLc8KX1BJ+8bwyesWsCy8g1wcFP5x2EH2Q5lFGbUUwtyxqGyH/p+xCQNb9niL4XEsrVRLhCmYnGa
GzDMpBuHzuKXm8GfHe90h2x6KyuY8DmU7fvRGmrJSX/rMFOMxZ1hD3XSfWZC3dUYDzm+Y0TR0Z8A
w2K801Jx5bweYZYRJkDy2KWGcSz/w5eUfaQ0laSqQeRc3JMt3F2xn0Q6SJSrYokXzwU5yAzJsLYh
34jRxUAMnq2Mt5n7Ss5Ne2tKvrYi4/ZtRHrks1l2NLl+S75VyIouGpXdUwVy8JdSg/O2J3Y2dABh
LweYnidvUX+LPE8dU3ao4NtmizRfR1eDhh3AA3DXBhBNMpqx/evI/Gz4FETNcwDqmiFAcMfdqq4D
jLwHox4Pums01ieFXUlTqB8hfkM3Bj+vQf0uebEHdHhfzOfyaN5W4LygY7B+/UlwQzin4DIwDcdt
PfEiSraLA9BP5TKB/mH2Pw9wRZkGQ6KvbFqMd7qfCXANgOD0ay8rsb3LeMWJUTluWsq8nno8f6Hx
iQWRIt7LUuYVBHSTPot4S3SBLI363/WfjuCswNvmDbcZmg9MVZoW1i+gTMwSmjXM7J9tSfao7QTU
WlAJB9lZP+jM2f9BmNY/y5ySh0GE5FlCpFH2QoVqrDu+UXwfJltiCldc02OyqsA2Xm4C6IkRFqVp
rbOBcw9gIldOkBnFNpLPngbFkOb3uh0rOrvL05WL/GbgFZWeOZu1rUbi9/3/t86wYLUfW7gLNgsu
1VysvkuzpWkVCQOETEbcuIkeK/YOlC3YQcfmCEi4c7DetP6kbScYf7b2VcvaVrdZ+JPvQhtlB+dR
YSsShUoex4UTSYbVhCJIRQLLilZx2aiz3QSNehXti4xQWeOwBJM0vT5TW0EuWCOB8beXwx62ODgo
XXP3C/PdmaTD5gx/KI2Vp/SADUe5mdZDvOnRCHqXwc09iazB7JpW+7yynUfFakTU3C3L+uTSFjSc
2jjpjmuYoNhicgBVYqdoSvLuTbtPQXJ+2KbnuoOURjjODSif0hRxz8lUvMoeCK9rsCKJzJ1BxRWV
r2KBo71jsSfuQkL75YcdqjydZe2UI0wRh88SPaiXNk8ff7keQMeGHa5Rj0J+oiPE+ZJ19nBjd4h6
DcXxKsHAZStuKqguTy1VunQcLdtD0HjtNxcWQcIZuQRdTjK8aQw1VtiMWDrxoeayfknqC7RHBSJk
mcHpV8zpe8DS/yknpeYmDVP/uYz8OPTdDungkx3L5w3lv9AAXroSgdNle8i8gVjf5tppdzqEt73a
ZqcRXA/B6PX0fUYgh2mTIx5YhmqKBWYurXGtyYushlaV/Pk+8XbRyfE/6M0vHysfEO0xL9tU4YQm
IwCtNYHo1/tZFZyTRYqSOsVFc68sE7x8q+3oT/gWiFpAi7/5LGoETvavUEbiWtoKLgeT+yTv7iuK
ya2oh5Svd43Sg8v6LH0i9J1rq2tjqc8DRB7wkGX6FKd+jlovLFQXu/4Z3EP46ZuSKFaC1oOvai4D
L3JVo66o5NGmQEsIv+paIYAPSJMbJtD+mzBQFgHZH/BsysAl3iOKfmMG7IC0tqCh78sfPXNQG0Kn
JxqxvuRGVlond6JdxV6DINAR/K52lL5tbEEwRpqLGnLxZ2vdEZVuFMYJHyHm+4ZQ2TdzyfdfGTru
LLWivZql9DdtWgtCtNrolxa+8LsLN8/rgZtW0MXjh+hs6lc/3Wxg1SKSeXX2lqmFlj/ZLepBX4z8
pJyZWMk9RB8rE/fZV3GPt9XOTeDGgdW2Ced3+XHXDrv4rxBmwzQkgzzxIxMu9oCQbvZBukM+h4vW
vGpLKubd7+UTqY8shsHIC82gAar18l7/b9W9t3NFeFbiLvg/Jjp4SEr1pys8cNuhE7UBCph10x+p
pW0oUAGJxn2TVZjY/lcR8sSgVCF6MlhmEjs4zIzm7IKf2lam/p7kUEwiCElLp4RMtSV7h09td9pj
Ao2ql71qJXxflMC1FSPOuIqtz+kmxH3Ubscv9rywSz55wJgMuRBd3vG5bEaM8Dw/flf+h5xNfOqr
2U9ILo9z0pDWsMTempho4ag5Yje1ClHWHxB/vmHBe2lb+i3h3FAXmqjsklIHMkuUYh3dnHm12UMI
YtcS78KgXJwVkMCNbWkMe3JYc0IjNuId8bYBiKf/L1a6OnU6tv8OUEycZrdBPJfIJ8ZdwfnboRXw
GLnB6Dp0VnIfIyn1LOKDTU1ablgpptyc8q6eBL8bMUMqWGCEb0XuzRCOQonuq4QKDFM8g1mQjvl0
cwcUAYth+PDLORr4k2q/1CkDow3Kq2eR1HIccwB5bicoRHsB6pIBUu+NxU1wnjN3JhnvdzpRpfWS
n0ZBcs8LTka7fxMZnA2HZ6HfLn+bAPjKu/mfUSD93By/oxJJNOpsdkf9yUOaQNwEI1mITniF9YNy
lX+BJCTi/Aua0cMdF2R+6nYdaFkO1FPLURjQK9JDH1glMe5TfD7W0UrKMylUIKC0YNbsya4rq5Io
bkT1038URN54uLi2jRw/EbN8QcvoAIH5hpyKYlUAemAOcVyiqJ8GlQXyhVSmuOudX6JulnUqJ/Pa
yL6ejQmL030ukvll9UBEmgk8SU45eXzvSCswNwkfZwR1C8yZXE/JEojq5oKQEBGcdXB7DqxH7GAO
0aIxKXdqXgMuPOkRfraqmVJEriZNvkwd5Czr8xLGIIPAJtxSZkVu1VuOhnt3rjSL0gJp7BsbfLqt
6BjmQCCv3/gIwTilS7jmcIR+chOR96J5qe0XSCccue0wkTA1kEdjglMr5qq5e9TSSFWw9h0VtOo0
Qx9+TZ/qYBuDzFd5RbvKIkt+8idlyn7hex+BGhxKIXZpDWvB0T6JM6FkOT2TNDp1pnhpPkShkeqN
twwym+XUFsSY55NnncPHtNN9EYNI9no5RQd8pHxTlVBeFkqWfUSMH+wMVhmeqk0s6SjM0nEJZ27Y
SvaPUFiZXeKXJy4aDwanguY7IzpM7uNA+x0vyKWaEFU5KkCR1SbN68N7EexqHRbKvg0E6fRfh/gT
kqHajrWiUvvKky+6h2rpaL/HnzFC7hofj0F29O4h3wxSTO+5eh7sbImK6GUtVXP3RwHxxhuvw3lf
uwKLI3pz6kPDg4yfAymjl3XCBoqc0sfEBTFWV32JuEQ553ujrdAv/UpFhcL8TK3mRDQx1AqDu42k
br5hr1vXt26PddKCtVUucKwWNaEw8EvIxMpcfV78QJzJDhlLRdqueYyhQd0s/1ySBsTJrCROs/Xr
NrqcEvCLiw7jrv0UCzHY0QD6EkgcPdI2Sd3KsAlgTehghC6LRUHptdrod6h6FBOcUpWJcOiH2Mq6
ocPcchCqDosPPUsDDn5sDLpRbyVzx2bADxxwG8k71J6J16OMHEyYPwFHv+B/IssXoyqWIRjVP70m
TqfJVDuG0lZKDpMlx+TIvXDQnWVLP98CF+alGnYWdwXFIeYY/7xNj9aToO7Iruyc1tco/Iz2ISE9
nA62HZ9BcVK42Q+MLpST40/7yzvAca16jMTy1w8xSA2BV1oMGIFxFqiQufDv8SwFyAruHVfFcKjy
91Le0MyYz+uYpy5735WK4X8o6ELJuGqV0HbfCceyr7bW1eZocKMPWKy6P+tn0I998V3PLWNSsZmc
+XQMptWNgpVpjJIBHV7lzwAm2QLODycCKOU7kLrLUUg3U6olg4EBqrHn3Y28s1E5Z4XCID9uopw3
kdsTrqsl6YyKXk++5saLTPQTmvuiq/p8OSzitmAteT9Rl/vN8Fp718leS/oMUKi2xecTOd0LnDhM
gO1usUTcz/jsppV5/6gT/ul3k1c/eluSay46JgSnpXrixqF0MM+ktQ4KNKFrCIf8yHSD7fNsFTiK
zrbgy7E87eeNrgrEFbEnViDB6oddjaiJ7hYuAx9HZvcX6Sd91TQ16YlOXvHtoiM0kkz6k4FQ+Eqp
ULiiQOS2J35rHeaTEESOm76PeE7RLcCjNQvVGwv6z8hJswMnTHW9tV89Z08AZqQpKJLscto6XbiQ
P1xqcQ+R0Ajx9CqUqsYTQ7Q5a429+4/G1n82adaUMAmFqnC40inD5m1K/SN2YatdIch1dYxEsbhE
UB2a5YfHM2Uab4bz+ehIrLs6VR7bAZvpV5GN4/n0BKBf58W6y2YVf3V7WVAEEVdryP6NLLtyVBrr
M5JwVxvc+cd8Kdts9sPFiHkMdWgKlufA6q9KoZQhKAu8nboqqDrzy+HbpfnREP9/sxpAg0Qkmg/3
CDrrs4ktDqKZ6VKzNyHnv2Ly08vC/HRMz9oQ9YBKa/JAMPNwHD378moiDexkk7QCo2TBCqzRTlJw
2RVvUjbmeiWMxVCisk1VcmGuVe25UTFMP0HVhTzZqkLvCR8+arYBVu/fu/ZZp1CVuV+vanMVDvpG
vljvwF47YBv4oVNysc5lLMqyCJEYVFqMGAuxCTIvGUG+JFo0hAPI0ltaGXZvLS9PlNNj+XWEZsCT
edFQBcRE3c7ZPhHaiP6zEk7hhYTA5vSiJ73upnjVtQijaZBqNyg98Ifec/Jhbzu1SxpHFSlvu7Zq
KHQF+cSeh5GpY2i/4gMR47s6bIXBkJjHUJ/EZYT0JLkQutIw5dqOxrajy3035LnILnMWsuoO+VKU
At3QW7hn8FVxVppezB68cj4h05sJeYz/fDi3AfiYBj7Pk28hPxqTh0YZ80E3iNV7+d+PGl/ewOFc
hpcnkZs78S5p+ROJaChEUcIqWfVyiE2SabInOlIi1mf7YB3cbQgKbs1TwJRGs0wUSFZLCMS6H+ek
NQGHVGEQeZznXmtSM0kSlNL6UY0nW41Zw8tlLFekc6yBT4VNAXWj+E+gt4SRQ2FrskxII8iAqiOP
y8f23Emj00zvsoHfHyhF1psbUE69nmfUUQ6umqZcpp3K7FtEJ4J4+43GrchaHbhMPoN/ANqbWwkZ
zPtVK1OxObSpHEE0fvrphUU5Dtj9tvWCC0mmLNrrcvnd9WXlwh8uBuK1Z6t030T3RnSb/3pqd1RK
PJQE+6gl6OWNAtbK8pgnxLNPMA9L+Vti+kf+red8aLPWyjtVc9RKJY6/Vlr51550kXTb3rjDnveS
jOKlSMu8JGKcn9Oxr79tocax2oMo3dqLjC3aRvKQ9Lbk6Ard5+1YVg5eZDJKi6aOaD5WAdlwAjg9
WtIgc2wN9Nm5hTVAdcZAguI200LUJpm/emp6HNpq7EIiOJdBXAz9UKP9TOntvreuPQ8FXCb9A266
YNXmU2e0v7FPtcfKkOZK0lVkQMJ5vE5+puDgJl3WaV6slCE+GJjCIS/XnhZilH7cv3J3lNFZn5FP
H44azqVgO7iDpd7GFyN9a0J8pzV8rp58JRnmKYHW0AT1oRB76IUCHEmGrW61LMJpLGVTBCIgZPlT
papeAYEgHbURIhcSH/zUP/pycoT0a7upv9CZMfhBTbvBNDt5uwWaFq186wrH8HB8NjMW24/DPl1K
aFSrtNY0Cj5krw5cCH/NpJSPULhpzwpjfJV/5NC99rYHMZW6zlo10KTLsA3YM8/GwmIYca1KKO6u
vyqOQLdp4WlXORtuVzb4prFWwwXecOIkAl3y2Jgx4z76p6SGfcDi1y78LWWrnjrNTMHvO70X9jnH
SAkMJnKG3JnHFzWGqdS4NVDyyAPfTjOvN/gCYny1p+5ojF4ayOs/784E0GBmD1HPD+A4/S3GClzg
T/K15iKKju/AJitAZDVW+4RTOkM4a0ULMvTbvlraUk5rmWfhcZWkWCwjMwFe8U+m3PsU3JlHZOwt
SFY8HnB9TCxY8cra/JywVaWYPRRDl8C7Jz7qbqt7UueNcXnnUtQKkoHw1S9zRu7+h9Qh4D2ZpDbu
alAf9YAMR1LNF37RdZ6iuuZz66uJhEk6a8s/dSeMUHVl+oOuuI0hvWwxjLieiP6/zZPOJasDdzr2
+tQBauJrOHCCRv9tnQbAx7TiT4W1HDzAsq3GR2qLQGMoOWGbeE6DSGf6bHS7b0zUmcLp5x/2LDa/
xbu1QeznQmZtLD8C6uK5aNnicj/zHT+SZrj/MxuKxzkodqcqWhH58Zkg4zKQdHWO7h3oqTgH/y5p
luhr8YpEPvHpu7czhXL/ZBWtNNrE4BQNTqEAh34nIJEY915m9V7yr8XlN4H7hrBzOgzDeWK1dqRp
hZ7X/bVpkcXd/BPFf6y7afOk8Knwf6l9dcUid38xbeANRIJdiRCkDSTiwz91afeMyiwjPaD4oTGQ
6jCIM83koL0PbYW7VfYc44oR0w0jFHMEUHNc9NHjiTCBs7d/ns+qjSn4zFIx6rN70bH4htic+6QY
MVsod1ykCA+kK49KHsj7VhTgC5/PyeUerlxjpWC+qr6rs6Qk3XyxSPBWM7QVTxD+AomKygsOqoYq
8hGK6o6LH4TTbmCS37hFvLFFJ3hKdSpkuTSKj4EZO+UImNAwxI7SjpiOAI6f3v6x3ftzu3y5dv9d
OG/dnA4sKTMJg4AFkjUKfcQGQB5xUGG7n4vtNqrREJOaN4Ep/z8HO79j+z3fnM/n6VuW2d7REAKc
MAzlCH2yUY4umZNskn3WvZ1C0b6oYekyq0DwNcV4u9FnuqWDF9um0faHEclbYVJl9xopR5X/vU/4
jRrbYB9u7qLaVJVWzPKHgM9UyaAgfMWd9Ha+8NoE6pprDuqSMd4mEyilCAHgHZr84GwZvWb+Evap
pUAMpHJWQgg+fcOen6YetUvGt71sk2z1Nm1ajFoB2OWlVTJpe50mFy09LAlP9abwCXpU2sabJM5N
9+EafS5+7fP2ckPCeHNF4WzqtY7pLtu75Jhx9p+c2hHXwV6JT9j/6uGMwy4VUW97R+Y0bor+3h2L
JvjofXOsDA+Uo7Yob05xNKdvbvikLepFtx4Le9oO5aAHTgSXS4XQDSqQZK0fNn1paKlk4MkImPvm
EzyRwlci7ADaD0mqC7KBxVAD9oxpolkWznHJDxBbrzRwg/XH7ijePJQHGtwJ4x25ezv8MOaz9+hJ
03x63S3ifxoT+6czc4qA6Jt5tDYk8fpGmXJ8fMQ+O4rI0KdhagetMpAbXvV4duwTwgZDiryR1X2Y
dYucaCFntUEhkM/n/8zBwkMFV43qBOoiu/cpRucpCtm/t4bZApPstTXkncRzfc9awEsiUVfSXc31
xhCMX3KoCwKvwnp3FnLw21qDkZ0RqFej177MPOfEpyZ54kSMbYjWb4dF/hPG1Bdg3k8AAhpN5iXE
i6RDgwiK2KD/F5CgTMljIo7v6po3zauTHb1a1c823Bu9M3rUL8Jh2U51QkJqi6ZEn+jGZTYcGMiu
XEyJP+KpsOmxjWbVY6nMSbPt/a3TBbrVRCcvf9v5rJ5oqoqfMlv6YVXKYV0Zac71V5ZGgsJKjV6s
tHT31yGJ4B3Bfh4KsvH3FV0XuXRleWK3uMoZGfAz/7HSdkkvPeM07jcZnryjr5ikVxx4eQABuWxH
z6dts3V1e++qSq30UXGJbdCeq5CXNkjetq+n3nqiTFGwHT973cEy+UXK8XOj4z+ljzN0aM3Ds7dx
NUf+IQbSErLVH7YLEzEGTvC6sx4IAQrGNluvU3oWX/w5XGreFxuwSFgasWXtsq4e9dd1YU4TzGg8
Qp0GwSpr41pyj274T+mdxjFgVYwRiVagPHpQN98By5nC81YhwW4yNCOkZLlwIl1z13QP1ZJ/fB43
nTwtF6Ffmb/cNZmY8czNU8svsL5349fNhIHJF7dUFpzzm728y1FQMWz0tUL8OYtkWJOJm8AgUcLd
kO7OCPDQg0rEX9g2GBbpSRp/+MOujorzyWDYmYXaldgEjsf0Lkx0v0K0dMpD5AMwLDMG91jIcuW/
L+N/N1c8wmhoiTltvmy2qMicjoT5xdclYem682wU3sP/ptcFoZoOxllyDo9gpgGUdNTIq9NiZ92i
r+fqiecXeR+iKBMEN1G2apvNqO01Fllj7FulE6zMF3M5SG23kcExMcp7hH1aVfBtSBrMm9S0u0Qc
yALLjpzjuD1OPQlQlX09mJB+jaUkn3orC6fS2RzmnD6vY6FKKlsylzk7x2aDmqbZ7bcAVq05QYDB
kGBUoxSG2N/MZKemVK9tkKxJFNFkRGEhFNJrpiqPLAaAY7e2WDXBMvLzt31jAw7qDO075W5qCjU/
oH5LM/GzRCVpJnzJVtE9BRGOPS+ksNZjwQm6IxOAKeKzJdiOoYithWHkvZQyNpbHKf2qNdoWgIiW
iFcJmNVV488Fdoe3AabTx2TYp8jueHbd4EBhMFZgUeJOMLjJP0NG4fx+NjRIPB8jgvagQZasDMXW
1TGmTojuF7xvOO+0gA4hFxhnb83ilAfxqg0BaKsZLsmeujId38hY6V8+jyHng5jH1e73Njuw7vZ9
JjhuBYSlFmcKOh+nMJNsCCcGZnBTZM+abystPhT6aPudhSnHADBDfXgReqZ4wnNs/xr9qCvLZe00
h/Fj9Zs0Rc8gV4euNYD7RQ0rISpEOmRnQNv+bfi7Urnh05//LuZ3A1N4wtTT2S9plbooLOQcKMaK
0GRbYkGqla+ESE87rQ9ysuc+Zq2o/pVIYnZ/sIp7hXLQbEdd11asO+WioZa2GZ4nb53s0ilcy3vN
8oXr+MflLEbtxOhYE9na63GjqaT5kdQEPrpwErm+4V3sNH0vtBXxXGj0sgrnAlx3PXHtA4kXHi6q
xFvAhTQAa30mSeg/O3dRAX7AiSjoWGbcuzBvqVOIOiD0SIRaCr/pPwCvJrPWWuQfP8BYjexF+azB
rAT6dk59yMns5M/LTjl8kpmxgmY4tXZse5mqMG1Yx1sGXa8hwoGFxVAWckES0gTMvIp/+sF1iBLJ
FdxvtFVZmiJ9/0XRDLDBGPqqiO5VOSNbcOwoe/k0xJVTfX708jZEazZT1rj7O/IPJ/TgW6JKMlmz
rVKDaUAH0k+Y1BZLfM9Q1G/VjT4wV7qeSftKj4PXxepQfCwdfJIBz2PcudXqCp15nAZkdJs3rw8s
V+5rvpzuL6azITKaUyNYxNz25lc+7C48j6Pxdk7Nj3tI5sQMJybv0Ac2GWOJROwZTTI/rO8Azq/W
R+/Pn4DiBzp/8A0u9QjmvLjFroFfINidNsNLtfYzkFX9qDtsEIrCRN5hFufxyr6qwX9PN7vL1Lhq
7wg/NiObY9qdy6IJxZzwIeiE85LRTrqEctuiZ+wJoYWF+uIgl4hy5nnUTWcSbYsMrHx1Opva180C
qu8VbJXOCEKvbbZwpMHIcWPwSn2uxMN1F1nz6dZhDXa2GnmKoV1veNpSpaZ3M0489x8e5JKlRGOR
qMSaEQWW1VTNN7H0EfC+sFSfeSm2okwSCSI3xiFlOhoRrP2BfPCrm0UBXEmt45bd3i86ND9O45am
b9rzaO+evVMZ57Q/8U99pnEvOFLO8LZtg6V0HpVBFBhpitL03BNUaAVKPWkPrtBaW9a8KStFgs1r
wj2R14NdJvZNZf4Gt5wtNJoNbjKcCt4JWS7A9b9O9098XbmTWXFMr7y1ZbjGreZ4vYcVHJKlVtmc
2QdkWv+SbB9xqXX2msZSbVKiROSf3wrNdmEn8jfPiWIPq2iZINKpPIfbzokhukN3c8vVW5dAr058
hfbSydYPt7oYmw861LL5+kAaonlW/KgYQI6ds+MZc9er+waKgLUC7lAVkTNz+RNWYm5l2tVFI5Vg
yVZsYv/PH3w+4JpNKu3ofcFzWMEB16cHukoauLgyf+vI13wwCMst+5kd931jP5WDry2GltYX86PB
T+PAvgABN6v8BnEovzXTkG1gDAc6KFQpZ/8sCSKVH33IR3RT+4eAshz0SMwaTeZxpXBi2KWYQlmk
diS8hwsIiN22ZFM1kyYnjg0rriv/Co/xWTEMk28x0fhHzBJjOVE1K1jvBlOSmEnjhNbRYjQQEqVH
GsChon1k6SbjhHz0vPol/mx6L3tlMX9ID8Gp4J86WF3OJRWCgV6u/lQUX42pI8vyE834+w65KX4n
FhlD/qfpokjbUWuA+l/W77Ban+FEhR1kzTFH4cgROTOvxn7cCThf8pBDfD22P8uCEG1vFbuU6FI1
+fvR5+CRqmw51vljQ/GcgwLP1BxlNvMsf5BaJfDvAKl6LaO1RAQJAezgouA6o5ZHI1IsIIAXx6hq
w7uRhuzmF2dvPW9U4usu4sfFy24QDqsS1Qfk4opTsTKBkPqEnqeXVU06DuvE3r/l7z6QzhscmZFg
YTcyRD5D++7Dglv/2T/JTo0lAa4gmb81+KwQGSXCECF2bVXc5pizkufU3acMDBzxuvddBfG8FeTh
RMVR1RP3+nxGd9r/xNiFfoDxfbCArzUT9HXN6qZZNm2rq2bRiBg0mrHGi2ivk23+oxqix32ma82h
X6TAsugf+/1lmKHw9pLf//P2odTQpOhKKRNo/N4JykpQpo4OWfBu0cRFjJ5eO0Cx1ile0OTw0KEQ
3n3Xx38H1jhiPkG1LIJHcOd8EdbAGVmGq9uRM2t7h20IjyHE5WxTTkycjmRRRfATywcpKILKhAy9
HMNQtWgZd+P6sZHwq2S7bxsnSnASxTFJxkq+AA3hRDNnZFCs+AbCvgs1lAp48ZwJ+IOKUb0MVDee
9dDMdlm2hSHBvrVbEXcv8/RM5SAUsVM48GOHR/xgbXZ+bSiKfX9PpQUbeLrQ9kuyO0p3gERcBRe7
Q6aQCoLsoUAilb+b6IWxUgXVTAXfJ/Zz3G1eCzTfdpNZv2OVDeVkglcDKvyTEY8JZnNZL9IkPgBz
SolK46weMXhPJle+Alb+YOQ5BwFIF3nsscKQDlt0OVwTQKOEAv+peL/RW1Es8BBec/I8D/UWpROY
e/U2p190JiDXLRnh9+m8o9E9soRngtSI7X4UkyfnY2Ae/u71NpRi87PW31qosSZFz8TYuGg7HPhp
itzEFyRyC33ZywVZvylLI+/kHSEP/8WDk4Orm9DdsnpSNjytHxkgobOLRBsKqpo+8vBXIIM46PD9
U1TwCWLU/NNlR/G7rzal/JB/VNEipobhBOS1uQJmXxquzq7K0MPLVc/ZWHn11s/b2GxWzMmiu/QL
72TGct2pBtn51SNndVxKbQ9XRv9XherJVoy6FeeQC3v5I8XyBVN+eOZvlFI1WPexEfkvB9PvGM73
DGOVN2Dx9oGQeIQ3RAR9ub5Zj2DP8qB3btSkPaGul0n5Owzrv8S5GOkyzIIUGDjY0M9GTNGqa2tx
lJteEMCdj2pLenKeoBVNuCcok3PGNo/Elx5HgLaScYNiT/iQIJp4JZ1pK3IUIUxHu+1Bm9WXTN8G
tdixWgRxaruX4NgyDKEtSXXm+zVW5XNZOPfhpGnQgh3zfztRXmdLCza5JKdjMZmyHmhp0E+Udn/2
mC7zIntdMgPZvpoj+GmRkaMpH8tuK6E58/vTy9OsVnstG2fvGaSnMWPojP+7Wc5HNJPT4lMGM5uk
hJ3b55xvtBi9eB5rc/+U43aiCiPSmpuSlrKQwXbDQHK5DCbWGYdEc4idPXeZ53+qbTTsPtW3nNfN
oWB3220IVx18vBHcQ9pNY2pZM9O3Fy1Kj88ay68jeNAjeuED1RZthZt03bg8wtDgF33ta+6cozVA
2YwunYAzYBPe2LZ+oiTyLIFYhWIO5RxuUzlinLZf2vCBzddJFFmnqZpJ868SPYRAIg6TNse97DOe
6KzHWR86JRwqe+OURajtUP6SMtX1+HGtrTETyGUbBMJ7qZAOitiq+2cHiCjFEOGiDee+YDjRxBvd
eALn8zGHYkTZD8JE6vVkCO26J5s3MImHZ6RTmgeqKskyZHqcQLTCPrJIbgQVKkwqiXHDL7q3WyUR
og3eRmqDFlFGYv9MCsPBPFQDnS97aYbborGjXTc7UE2WXy9VoERUDMhorCLctCwHYxArtuQp60vY
t8hdUhKOonW51ebOAFYTNDzbgLC8H06WdegRY7VhbgKZOupjr7+CNObP4RxIKo/XwNaLBjVjB+/H
pLIfS2RwPWl37HQt+BjqaEJbEG/2ok+tdgEYfLS030xssa7hliEUrMk7n/aKoGmK4WAjpmbWvAOg
YyuABa0wmLYrw8LqfMj4vbJ5K54dCldp/3ccuuT7ArHfgCGZKtnhacRhed3cVF87rjWYL2b0nJp1
PjXXttGiQg7RcpBgHGTl3D0mmjKzv/+c0Z96z9bTjHzz4i1dy0vaEavHw6hweQdW6Hrp3b98zoML
oIj4wtls1dYL43tg8Amchk1ZrpqyocLThhRKm2lOX0Nv/FF4NYJh1FgDYjMRpX0mzA5HI0I/IG3u
gUG7MFPclvf6ablJn2qzcjSOu02PoRwWFfAU7hE+A4Mn6E1Fl9zX3zGvUNy3v4e1XDnfBY7Lct/5
Vlgrge/8pqwBOVVbRbu00utG/GrJfxc2tPOJMkD5SYr7SL7JXVHNNbRXtQrUpKQnxegqPyI9L/KO
iSCaRhuXJwiUdwud0Oe5fWMUwzak3rFlF9i7V0YTbM0SLWZYBiiCISuuRMCpiOCnO1b5O+gL4o6q
f9lwC9kgUMIyXEpKCuQ4+td5PKe4yqkROviXoqIjyd5DV52CBUMGf5oL6yvjxUTJpV7uX067gJdu
ObY3eXGbSS2eFZpSsDbkaz80dq36NKzo8Gq5mWZFtefXweZNGVjvqRnhHC5uqYPR7k952lYdQvfY
qUsiNG0/a3IkhSx6PdVR0ZHCOU5n4qamF5ohYddNJnGyZKhe26zg491TdHE3NPohwKZvdLCGT2BN
vI2EfZrm8PrOZRg5IhSUegR9W79SyUuv3h4tLKDOrRT7cfxcsr7isYKkw9dNMxYsXVpNvTY3u0MR
5y8BR4W9W8/4YRz84dzX3CyPwHufvJMOj2Y9bARlClN7wZ3qbiGBN+lFmCkTIuUNygqeMykYSGTf
AfTF7S4kRuxzbgr+Uleq5teMa4/0HajCaXdbIvr4JXHVpOP9neh2KZmtDm4xoyckOaRpO2dsb+Hb
qKXJdsTefGWaFBsnriNRFKrb61w8oHoTMuski0H20lpRZ8zMe01MR2oMhKjqyw3OWvTNgQPnvnYu
U/7zuTivHrYJUkp4vbc3Tq6H25aBU2lPVC+0NJsVj0QNMbqkH1LE5gVOHUcfg9sblkGLlgv2BsSQ
sZz/rOrUuIe01G5vVI+61NgO5omu+Wv1/PxjsNCCz/TcUS8T1njnvULi8JkE680GzQrDfb/14ibm
Dn2eKfVEwWyW38u2otd4Ga4oFfsGiaaH2FSf/yAO8qNxrEpZc+wnoP5fjc6vuKIZhRFsAMPzNMw0
5u79I97VHJIOzn8mtDoa4vI/ALaqK5WJjqa6iqaCRY6gXatJWZvYhTIurocJxnAQ4jnyWnLkjWoK
0AvBvrsYP/aJDnWkpN1tzC5t6NuTeKX1cZMraoJznyJGyw72X+z40zne0rNxGOEvYRAHzkpP/MMr
lt5eMEENUE0oJn+DHFvnr8gj+TtsmmtgAMprJXHuyk5mFB0t2l8LZHt+Sy5IecjkP28hEa/j2D8w
mRZ2ax1dA8/gpXXvtOCndyzhMHvkeMHwQ01G8ANcMub6XFzB2Cz71V3H6nkPT0gTBmPa3i6CQrPx
WWUDm/y001bd4iYlRL8FnrBtwncynXa9yq9Jjt2LAkgSI5kla+11+yqO5rilUKgq1bp1cZwQPK9F
UfdQlgmxkO5LtOtV3iLajRZ+NnJgmFIeVnFFt/n4EjF7RvwffPfXLMqBc2vfkUfEZN/cyMhO4rPe
OrD5AUl0CxbnDFNmhD8LuDHroZ4LxaeD34qEUtWmGN947Iu5hTpXYgKHiEYa2Wl23IYojxGJQwZW
o8grE3du1bsfiIszwkZgdzi0yl+6ydkS2py+PqFaRrxdx3QPy3qDSnLVIMh0A4uF3nXiPnMP0aik
QmcEC7wMp0O4FptiAP/VPterll+cpy6nPc3W2VoYTnXRn3GqdU4vRTgxFrPi/9VKmi6oFjAnizAp
5q8a9FwoCvHoh2w5PXZowtIsdCBas1uUj0Yy/iWGL/GrLaE69R5dXG07SNfR/eCfaFS7kjtFOioc
0OYNZhmaAeY9RAqCp6HOxFHD5HRTBj4RX7V0JEKfzIxXHZLTaXEPEAvLkCf7QEHtst2EeWe73LwD
cPN7UCqcbrOhGSYTcptl2R9mVbalkIKycgFNK55UqdLuPOFVrWApV+Z3fTG19x2pSLiZG2GrvaN6
34Vib7I0K0Imo34kW3NYthMaaJByNNp16KtYdrf5Fv+egVIczrZGP4tikschaEQSWTgql2MQEStq
AAFzlgDdrRNQPqhHkYCTrfs71HDlkwmaEzhUdHaqgNRTXjhapon/cFXdbFeoJ8rkLiPguArhOu14
MvRGVZmXHYU0ZGMug9114BwbxVJkgVekUn1ebHUPR2HoMyPgTWBceKZRgfyhNpTwGEen2PEc/+e9
saUUD6dKe57PZWLf5RUQgA1Ab+hWvWx6k/udD/2UuB/5R9lJCDsjFdaRnckHLTFbjPY+XtIWmKKY
DULQLa+QF7X9sqBosUWSWKg6xXWymlZOhMXrnqeAII08mD9KSgjRraty1pBeQquh3zSsXmjvMivb
VAJgchsKYQpanPjsjYMntzUcvcok0oK5tkoPrdfiit/twBhKuQxPMH0E/MZEvsRDA9f+CsiQHs1B
WRWhZyIRBRdvKBz0aXQco/rO6RcIfjLkW8OsXkLZJ06763kVWm73jr3AZvADwES+JEPnY8ooTwWI
YsMu+ktd9a4r6fXTtTuhs133rvudyrqtS9y+9MAlP2V1pmGGbdZ3+bA09Lb+jPzBbfckor9oysdD
xsxJBb6kN0if0yPBwvvpB1nzM1kMuSiiye7q+E/HEr49dR5aZ52Bio/UzBv7iKihXfnH/KaXLwHR
beXNjTNfU2b4OKl1X19KgWRI71Rf4XP4m+sWw/3Tv4Amlo6J+RD6f98wi40lg/2+b1js1Ah5vAGw
/HjN7bD38hx9Afqs2t+VMO4jITZq1NqWx3R8gjlYPyIev2KtQRb/Hokr34UvDaRro7c6vukm4ZRe
sS1y/xieKj7SFE94nh7uH7Saoy/h8XLnejnBYzsUuEh/C4NDc73yLuS3WGnSyJzXGRZ75XofKWxI
K2oW4cvEs4dUQZCbia36bsf4E0qpU9QhJdJG3C0fEL9ckRipy7yjzMgPTo9ClIpIKKtM8S0cn3uN
Irf0lQ/8pFcakIZm23f4dLh1W8BqdV4GTbePox//+WliGpw4NAGPMT78kyrKhZfrEbjjuH7Rz/Mh
1CZmcHCOtjnPz5AORn9/Jiam1oLUU42j7ZAYkHnDbDXVA22qx/+rZXV6geiE3QWf5El6h28PZSrT
plPbTjt+eNuONh3zl08DmHATd+yyouhjfNwe2ZfcKDe3uWZG27TZ2F4Gok3sXm1nfp1FbXu0RM/W
HUNPWXnxyTvIFSkB0aRjzFYdzdN2KEqESgx5nFc1jItwi40B6pVKodrm15jJqX2FWTSprzC04Z0V
Zm6t13ypWH549ZAyheeD4zR9GPBqdDV+TAMMSXVRytmz7saPtTILu4kcMnGWaPCbHA0w7NZ+HHRB
zxT/nrOkPvD4XHOVV2YkY3oScXShbT860Wi4Cvf6Rsh8pE1XiFJ4kVM9fnQrQTQkVRbsEgx/WaB5
I703V3lBdgpgcIGD3DdsbhrqD5mmEie+wMnmMh6qrRlWTAAl9CTTsYcDXydhoP1Rt8UvKkWCiaLx
hV2ay/SOwNas9UpqpfFGRbbs9uW6kx44BhsQ9lCY3lN2plVnPF+XThZGqY2ymozO515zqO0k4N5K
jFnmn3j9PyEizTq/sCqeNApAeoT3/eWHQ3wfzLkGsEMpTRuVwEC+ii8TvEUn4ouC09wRKskLt46c
arAph8yChaFYOMMQ+kBWWC/WA5861quG4pE+n3h10icmHEiQSXdLxxIaActRJkkRAeZHOiA0IYtr
WQfwbc9eqFD0C4H2BqvUCkQXUmXwGLwBCBSd1CkXxiJ0gWxdchZ9qI6ZXi+kiXA24CDt5MIJU3KG
18HeZByAWn33jNBnCR83RRLTdQtLZFwdPnlHtDD5bIoOO8QjniQdRimLwlbcUSD3SIE8M/m04abt
p0kt0bbImi+d0ei344mF2LYq5+NpF4xh5CaKOUgYEeogAkAge+vSCutnXnv8Od+ahRDDRj3hxZsn
8HjuGEJtH1WjPdFlOFYixf2bUK/xV16XZvfwdnuWwpp828O9vleKP6q0xYOUzP/c9SFNqCxBvKux
bUut/fYbL18by+L8XT5bA1MdWH/jNfNIqWl6s+tS1rIVDsagpamXqfXBvmh/RAkyOEG4nbWl1Pp8
1aa6Dd2Oh45qptb6JERu5Q4jgEA3joESWDDmSTW1GW8v1LVl/62+YNJeJl4cWDkGUHwgONS0TBNj
fGTNx5vnjvfgK0WP0yNYTlPPHJuYer5WDQWqp7Uq1sjvgKSBJgyj45P3wECTZxwIt6FfbZb64dg4
/2njJCxBvnYf+0doOqqBmaoWDAtyjIZ90y9hxazS2xs5Okn3ze7tcFdwlbTZKiZ66BWTfNTkQYKY
5hYUx/4VFAiKyytJiiOFSXHcqACmBIfVg0VEZcnxbEj8hBAT/c0I0QnxSNS/gMJbl01mo275DTxY
cONKcivmQsot5+jiu7P0nr4DqPxYI9CcSDSJJsMUPTluiAQAJDhNd1sNMGNoOxeU9LVuFG1y5FA5
zjogjPGdaj06rWsqrX8ivrMKVsEnlQlE+WP/ekWjaCP1f0/36kKjU6sV/8He+lzAZa/lAtOCT+9F
2aQ53wG939D0bD7ewK3HDMI/SOl6LValkNj/R/MoJTbYlGJzCu4Iuv7eZ1ilYa7WoFGQzlcXG1pU
axi78APbQfNQ+0IW/KrxswVGvWk0ZzxDpOzJkLjiMIXI7wiCDGJOMddiCHXNEtiQDhhsZytzJV9k
rKIFzanIhDfpuPJEQR2xgwRTLZXbd7KlPFaXoXV/7xju/EdSWGfb+vjZk2bXMuBht2i/FxiYrcGC
Ac8cMB5SgYMxbD33OYTveVRVzPc9fKQlvmvR0jbtl93i9KBSP46062sJrVGVEbS1FDHmlaqSmIJX
R/pW8zFW+yAMsJmWHNjWIlbnR3Ll5wDcJqCZ6IQtSgBl7sjYoEuogbf5jNePscHTED+ZMXduFnJk
Xi04nBVhcToOSgo4dNjgktMwG0p4RAlSZm5aoGPJhdRlT+Bddl8MWLIve4jXHlpYvVnVW53GuyW7
s+nM3LvGyKg5orlLyRy7ypNhPHR1nTz5Ohs6qhIUs69oj0x8e8kOMntg4ZgnV6UoQVDtMRs5EkmK
epCV/liQSCnC0GYFL3X8nggPtziKOHNjH7YkUOjG65qCe7f8ucvw129uVOMPX+wHYohO/inMDhEK
A9CgbQgLAhikrFh2FvTjxNhVte2mgJe2f7xY2gMrqEPjbhm002+lOxbYdkmLw71Nwv11OUhOzcVh
5FDaiwR+gwwL6W6QMxaDPPZYpCetjnIKSQasr668xqr2D7Kxl7nlqUm2m3LnRlMXdciGvFabH95N
ti+APX+gQCrfiayKi2gKTqeyshhTIgrboBbAckHH/uY0T755TXQgb9yNCKqVAs32D3tvIkt8R0qT
Sd8wSkNREhECIP/+QJ96YstSARv5hUqUWE7Ggx+r+xgrRMK9HFfpQdS3mdiHdTpifrQFdT7rGALA
0etx+bMAka0H/ltjibLGZnGR5ovffgx09XZBkrQdBTam6OYS6S76t4a9VJQMiKx7XF6C8LJpCl6f
wkMgCoiSQREwqZLCJfxDvsK2V+gBCkQAaXdbPSgkKOBBX8tYjN+sp5o3XCzhMBZtmpYignvXBs79
sYYPV/DsgmYNZ6k8o4RBWLGAab0Um2cUsqKbiv8G1c6qByUiSxxUBJnI44ggri9tur9oozVGtJgk
1ZkHMwyqNSWBn6X/5Z9SlIyhvSs514DRQWXdzQJI765UI66bSQ/CRsP6oYcYp9Tr7TkFQnFrNjCj
Fd1pGeXstQclAqXb3Q4bWt1NFDzprt1dEF0Jx7LLw9ZksyzZFGG7zY8XqxX/keSrJCD+j6Pecolf
kf6W2TQljLVzDZEoHhhcjrK/h6WInd1iKBYrB0q3/52UdrEWMPDLsJfBHejnhCweh//e2z0q1Fd6
76nsef3V0qg7tvfWqU1GpNYB1GUwTm/VH4OuGeoR+9uFhzUv1Bx4/x6ijDau5h9k5yMNXWkYB1sO
n2kuMhBtbNY32QCcLuUqzPoYe/Rfif56CoF4Hw/HwNac7CYr7AVZSXHrD03jn5HVD4o/XNNZAUXx
mmlnf3ugzeayTXuG1vNzYHrzY29A+K7Lv4vfMvEQU0Ixbr8iLYOOPoMu+VpDW+fdYSYL3BxHK/Bd
0F/UCQrtBH8zb6dxDLluKSqQo8n/m/IQoxXBWZtu3eE4pnOn+1PXZlQeW+xp3WeVKWd5RgmWxK9U
60R3KcCYtRQ4ONnMiwkKhMp9D9vU3OYC8NQq3Dr6/tY91iSEemzknK82meh9em/s03CcfWKNl0g0
PyYC1xQoQ5cXlUoFXnj58IW3pMEgL4zCvCyuNY+Uznf9aMFs8ZVC0vE5AxptFIc06fDXOkvPwHC9
D2vuzKX1Bc8E8lBwAfdw/9POY39NQ+MXnQWXK1tsajYcCagunPMICo8FTJsdraOX1kpnxwdwxE+B
ex1DruyXSlDN7LLJ6y2/fCY45tDUNg8Ns8B6uWkGrF2VbLfRbgXIwRVcwEfD+F7GX8dtaFxCvnZE
w+Ai5B1eVocTOABM9MkZJYHtfsXgC8taZs84nh8AmF9cRkyS7Pmgfza5BQZwa0sms9lXN4esmpU3
21l0I0T+uM/BvzCibt9WnSsIdbLwG6/ROA39SAQs4/WMx0g35K2BW7URLsYwN2CaJ5Cjfs0ecvma
jt4OLWNAN4O24CX5gnDxckItc2EOlNKP+L8KipPsoYr/DFgGAuPEHpn0TPLLwN3jQSiNSvA8k+wI
DrKB4NwuxxdYWCRZgx3dc+VkGEXkvxEchKLK9tI6S836IESvJ3ziMzXYzstuarVmCLnQDxWelv6i
e0CZx/KubqXpWdtzlU5x6XAbeVcfFJew8JiTPG+gPWqI/xKgDFzhzEcR6dje9n+w5LfeV8kjHbDx
6QNJSdGsVX5+5o3lqpjOXKqvwz94xe6GAaoSzm1zG2kVOBc05z4rXa2wB1Z+HsbGdSe/JyTbPRHU
ZXg+jNidv6ddmOECHZ5010Np5YOsvxp+dqTKznENKRvOj4UaJADToPp6x4OjmjpceDoz/Hrt5RSe
b6051DWXQI1UqKg9M8Uf4wcFa8hjkN06REk+1B1UrWWTVhPEsx46i3ShJpAJaQO3dUftzF13k7lA
iYQ57r7srBjeKJX+CudyRt38YA6+BVcSH8kBoDk3R7FxIi99IBOhPMhV6mhOK/BgP8nlPw9lFC65
omHjLEWkD+QbRJgiHW2MqtjZ5iccdq0b3Cc0nww1+eJ0Vpjb5Y2u5lCZjU8pAs1D7xQAu8nnablQ
XgheeVWPAQPvHsMdrT1BEFaWvaF+J6oT5umUkkJ5C+hmRhpcfrtdYEpYMKau26jVCe3E/f6QQxue
0A7B2UkfLH7sEPworKnWF+eLVeyCKPLE8m0kaZjspvm/wknBd2/khnDJo/YuIMK26nUI8OCGbGh8
JX+09MH9k+0GO5RaNiX0MUIO/g4ca8pfohpZBkyrYXapWasvy1QHzrFxw8scuwFCrYZEZx8m2mrP
XJRSTm5fD/GiUhbec+B8GJiyUbkT3oLkAsONhvv8adPOSQjHkkuyl0CZCeLHAuvz3PO3OqxF17XC
KNsULyIYp9K9yxp17Z2/U/ac5Ph/bDyiKeCAj2KOCvuaRZqO8Gw8cgV9eo+xoVm1Aa3jwAP+Z11J
c8Qnmk0CII/1o6QB6EmeFi9H8k0Ge+4tBbafMPcUN76QB3L04NmsBUukuXk3odjZHE09hJOBpqnL
zQx14wO+2X9M+Z5TeXbpna3kl4r237Q0j8MuMwacpgTOJOXA9+Ela6D1y0LbNQj37x8+vWIhwuFJ
VQpsVlWjW/7vCSGVxB9TXKnLvIx5jLduRdxQ+hV2sTg19XmGnIcNjo/sTJffYio72yAYB8MnyGS1
mFBpmYQrMtghYNycZNVdugcOeQFXnfUEvINdDdueqrYZTc5fxpGLXNb08DDZtQ0WCMYc1zW0c5zV
wf2dy4S6qfCW9TEQh8wNCNFTNcSkVWbZly5ysYdzvmv9kIa01z0nnKR+iTmJbMDgdnnTRwziZ9M9
NBEeeFUTMtXV1NYzAB5Q/8KXW4NijkUA6tH/3wdV8ECcUmoxSm1aGpVD6hPIbpe/4RU1tWvRxa6e
12d1VU+dvZXrQwrCbAuRTir/mPK6FS9CQO4t4An0iUI6NofIDj0Ed4NBPKvq+DoZg29YmKGsSTWc
092KXjYYmcWGa3hp2v8Ux5DWTjEVnGgo3VviwAEgdKu0qkYNeW6eu8TDKv/7bE3j/i8qfyQ4lyuR
ulswmOAJ66fcLU6BYcjR3PXcmSS2oISK6rlivhRO9TZ8jgzEA3/dS7ZaMHoJg2PbAsNDJLQMQMTW
iak5t8NoAkrw0EjuI7/RXZrBhwzQWeK5BoTphoDo/cr2GJMrOwvAuGYyuRyXZ13u2JovQ+xp7ZY9
AhhF6rSW6oEYP/i0hGbeQxJqzoXMyDqF3jypInU3kOsORyuEnpygtS+E9TR2uj8942pmMu6WP1b/
2+CURHIuyHy7Umy5TOS7mzZ9DweSDWVSeq9V1Zkw+uFQ/5roA6CClQAO/sAgBoPzHP4Y8SNGpWRw
KjN6pYBcuMYBIubq7uaZQ56GN0dfFGRtpWNqkyA9oAQDhWH1mtfQMwWbyORngs8IdOTPJL8n7BWq
JbR/A24vFQztGbq5DRCIe5Rm1xUdwrFcZN/qFSGgxX8VEhnrCtVAAeq7WT2hosxXjFB8Ajs/wTKx
STpilPYlbfMamYCHch41O35h0gb9XIAoSUUrxldK1SDKsDK2ZEi+ymujcmhz4wvTpAYy+UEwFyrs
iatQVMdKadwuHLSveDDt3I7Ewd/Wku/+7ZM2m+GzHOiBEtPQJb5iu3rzZaDllJ1C5xJK/nQPj/vI
JNBWtfG97AWIZj/BSu0DyePWjDNtw6DDzBHKk8Hym5V3HaedJbAdgsg+17iDpg74FSEKI/O31SyU
l69W9YfjQqcetcs8PO36RNHs49uPa1cfadbRncJGQjyLOIrQvGeYVf4zfS/9m1omYRNEsgewgGI7
zQcST+FD9+zO1tAdIP4jn0E1mm4YWN74oY05llyErnNbsNXaskbDBaIm1x6IEv056y6sI3f9efXI
Xbo7uxTmPNPvoHEFY81S+iOY7tWbKSQOJiMSwBSZHI4jk8jpKxS9SAPYtQMldvjxJWgF05GeamNL
TdmxuYtPJA6U1CzpEhkcxEdqzZsLH84YJroizdiV797TBb3BCOkHL2Jabcj+uk7/dtMR+lr6+u3F
xucEPLcTMObs1e6GtVTa9DWnPHV7oQ/crcFRPsyGUfV5mrzSCJQJKTF+/XVIaUjC2Bq0Wp6tWn0M
vxmpuB1OVVop8kduX+eu4nrW30gdxbChlbtEMiEDmNqBQsk9FuPix/PHanU10uW4arzbKgWOZi43
jUPh4fWC1HSiS0FQdgcam2YPJqAnhcFAxoJc556d2E8f9YhtcaMWkgZ7eyUMhCtWUhP8qqig09Mx
bSrRrzroG/9I+dCNEu16jglm1rGAfhWwShAajHctL6IJwXrxfFk9javNJyYrn0MKJYZOgIKz/rNJ
y7nVo+ZdJEiyk/ZqbySLZ+2KYd+kgOy60kbxjaDzzs2GdIARvVvuZctM00DFPew2Vb6k7w8FI/GG
1P/tA4DyFIAyp1Pq5kOePbMNe5ETtsV7NLzKyzkRZgV+5PpTBZHvu0YetTuKVtlyHlxX0fYJa3CT
zx/33lpj43mkRTgoXpfsG0s6GSj9NhHdnDhZKp79aQnusSINpakteFC1uvJD+YbCr7LDcKISGAH1
7CbXf9AYZKPi68ZhuiUgSlAHTSKHD9UISZJabpvKaJXl8ZA6VFREgVe367LjPHcgMxw3izo0J9on
MoP4oi+kwhh+E9SxOJ3lqCVAIrmwGQoCPL7WAMPYhpytncyEg8cAI9ZnS7ScRFguquJgb1AMXlC4
ObdzaY5STKcyr1Khy6MT/pA0jq3rLUE65YP11wvbgQxAsRFlkR6BRxxvM2ycPspxCGVmJAxPSHNN
Ug9MIRF/ItgXTInASn4228jT7R5VnY+SYMa407+yQ5Ik36VygVdhL6ZwtYiB1rllUuD5wq6dC9dH
t1FwKDy73KyVF46PbwXClYfo/XMxYq2adIzBI/eJJKYj6ZSw0kZzmV6UW8CTsCbGB3YjnjTCh747
mYmoTAjBexITyx94jzET2qCSitNv0M5R61K7xLjrtehSJuDN9UYMt3v9RYO2sgNJ0WiMXnYuu23t
3O0VqSYLG1cOUCIrTv0y57Rj6SCJ5B+D70rxUUkpXw5sazyVLYvWVN+iMcngL9b6SRDhL83IBbfx
30pbOi8dPHsqNFwABOHSSYMnElqpRvz1yJvkX/HQBdP1qeo7xNTyx7QNnloj+KbJOrVq+jwfNO2C
e/oIp9QPVsmVSD0PGD5c0zl3yo72wxlyggO0RZ0jlKz/G1DuVYPwn9yNLrIc9vHzgWbpXr0fuVCV
URoyYzDraQeQPqac09+q5g+b3ILmW+KS4RSFwogB+4THaXd9Uy3hX/iZeY+geAmmCoBdgjjBeVGQ
Jlo526n3dO3xcCOU/vTYxI+/dYKsj6rJRJXDQPBES83HuvgsivwMjEp3+cl+dAyBw38blKNqntzd
XNfxK8vrpLcO/DQP6un3ErPx2rC2SCNXzChuUl+POpn+SjAbMguRGQ5SDBh5UpPBexAdarNtbOOh
jzwkbgZhEF9eXSy+NBGVc/fKcI9WNyavGv4vW/suiYJi0zVwpsrCnADpt8YhSiUwBEwRlbVVtJG4
39Mgz2qChpEtmV7jHZhOFpOr2QvYMr7nfDyIubF+q5gaHaFaNhxbioOCmoXs0AfCncQvxNMTwxJ+
HZi7/ZuX1Y9FKX0nCwtReokHa7Ilzko9mIFPIHNki3iuYWoXKd4O5jQaC+xZUT1hU6vYvaLxwyIS
nWEeX9sqHDxKDMkZwbWrS1Ja+qHrd9z2fJCain24IaTJAzRkPv9GEj1LVw7V+1SkryJsK91AaJvn
4g0SvCS7biA688kHgHIHTC+cr2mfkdisMYeoGz7PpBHJOU49gJgGNSuvSPPcyYYwdkfizkJLK5FW
0P2V1stj5oh6ezW2KTujUA8c40CGc8tqcNUMZ6bqBJ+Z6yKBlC2n2v0Ee7dTMedazYJU+5JVndf1
QIl+3BQuLxRTDbObXfZctMi9p9T5Oz14aEDVGg/SmnyP7x9+2x2JbnnXbG/ERGauqou4aa/2Prua
PVTbgwoFbUAlvQkdSQi49T7n/R12HqjJjeB1ATarA1DGNhWHnBKjYVjRzzJUSsBAaO5Hg+KlO3SM
S+56ss/oNA2r07OHwfvpIEAe2skTr2EbIvvH7a3u0JROQZtE3jf4Ngl3HWK/sN+LoBjkRVCCCMyV
mElwubpAaEAONiDTvEPPcbHOu+53jmQzqOYB5cVZ+dsptlMq+BgRczx7hpD7+Z//K3mmdFllbYLv
o+NEo/5l2SI8kgc91BLfI2y03Xt9LEjrFuM8uiOorlxG08Qx/qBJv7SK88em+xtqe+cqKWmhoXE+
7GNpIBR+aaTUeEXpNGUr/PVYzYXjOYxsYmU6Xfm8AIjEjezTST2buM3EzW3+awvp+5iIPDUZQbHj
TN9LWiuF4Q15/pT61IbeLUTnoHrzmBZM7IOSE+RLaAyQ9PcguEouq+qOiwqOslFRXRcKv8sLpuJ/
mi/8af9J8N6Dy1G3JdV8qAEAaJHct+ibcXCtDfPOv7a9BDBdbjiIpUaO9Ex51bQcshmXvV3D+4h0
geLXsBahBZbqGfGd2fU9G0UBvHqq443AQc0YkJSSgYVU1vaMr8mpZ57faM6jdYedAYNxhUBs5aGH
NeeCmUiRr7MLyZsc67v50scUChe63U3OfD3bN2g4njn2I9iFMv6mbEy1oBwYLGCW3vFzLORmjBE+
gIB/5ioP2/INCg8HrOieFl+/6I+Lghrnc6aGsh/meNbJ6BQ3rRxEX9ScqOdPxe0bqvEzozeb8MVy
JlKdFBmkfDG9m+mNd69pCQbpnp7SJ6M29gMRdkq2fu28uAKyfgNnzswOkLa3+S0R0JD/MHcQLTS3
ej9kFeE9Std4jc65kRBc1BEz+LVUzsTwll8QjnEizqvgMrO5228MdwufxLVw+QmdMwlRxReA2NMm
LiZrRMYGgBuMFA2dRY+Sb2X2LPc/lcVX9feUroJxxL2c96yD6qgqqoGCW33d4Y7HLDanRqa+WHsv
7DIPQegsQ2udhEDRnj6Qjt3FhvDEnL9erVJwtXbbecioR5ul0dje1CA33Q0A+xFUedBEODYx34b3
/rS/p0Ix2J8V1T0J/y9qsN0lpaD6BS2Lo8iIo45uxgI4qYCaqCb6HyP0q5P6vN8H6xBRfADafvQ1
e6BZP/0Kc95bqmbLQNXK5IY9lfLNwzDXDszdxlt3O/GF1sbM8yeUYnrZFk5Ev3R9XR6oEeQq7BiJ
AzIhoFFqNEZKKErBX8Y6tr6hSMtexK6iFKWfI9Gnhp+whk+N2Sn2Nqnm6Hv0touVWbCcWJR+vBm9
bFyS4wxDAvUEIDd058KdJniEC9VD3sHFmni5LwIDUAlX/vfoR7CA9tQxmH2zCci96QKt1z+f3D2D
t6mdNUaRp+aacFNSKneWSH5j3kbh2cResSqLCDJoDOJu0rz7mtkF3m+MZshOpwlkZg6CanQD1lWL
kkKbAt00m4bIjNL9QALprgndoLJaHEIc7svtlQWh9MjUs0VnBHIuf+XywdnWrIJyierx2IC+AfVC
aJ+xIRdsJSlgbsxCO+UakKujOpDmEKmuSzwRpOR3L5gsBNffA8eXDAZh5Ko+mpCaOfD09DbiqhoB
+Dg7TzggUF0O4F/JzDGE5WO2yB3yAzxj6uhSrffyednIi+BxX6S4Cs9pn6g7YFML/JczjVixlCXj
dO+uMKUcXVs6dc6g1fQBF0P+H0GywR4E1ACQ8G7oNHU4Xl4JHJX69BihgOhkDrBYIySjOtr9aV2p
FdEKZm7gSiJRRDnNmbn5X6evrOYnYy9JlNp+xEm/d6oLhrM64Eb34gQshofNqEfbPbupfTW+Qv0r
cBzn8uLRMiZWV288b76tDgryNxZDPx7KMxG2dkivTSajdAtjyqO/ZqdmRtdl7PY+5lMn5taekuZg
qkRkUdhmAL91TkLzVHEbS9X4l4EKdlvz0/XEQpmAcnOTX9pL9H6BUYz/J4V+wTQQlpc3xi3zY2hf
1yLadLITB8E5f81cZwAzWciSGdOlIqhPDmE3vG78neUwufHlT4P9PgllBscGgznFwLBt82nvku3r
J1+ESyeDQ2YBkrVK2Hi03GHQ55p5tfdsOMdFbIHeFlMqX/xSeX5jikscX22wqSWRz86ndZg9vz7z
YxczWwHVcftY6bDPt58XXt1AYrSyhPeyxfNj3+zinISU1VBHg5IR2PjCjOSC1wAJ4sFIxszoU3n7
32YTs3E2VVQ2jQobpVhOdSpKZLvLIvzPp2zRkwOEdygMygTqft+Q9hMt2v0v8jguGzJWg2vqxhyl
gwXiCxi1OtPgxBfQPCSmw41jkqebiXsfC4UYYJ/ghAB44tqWB1jV84FYZh86TshoWDb6VQRT4wkt
skxoWj4i7X96c9/v3ZAsMFWdn5aYUwIYFkHTfQh3k65CIs83sq8y1ThUBQZAIosDAWQvwobTNH6z
bJZO+d2Gc+i6VyYisYwr8wamjQUVSFTfv7rf8tj4wNfRkVQm6QZEo7gn50JS9DqtdBAcJ3fdwwh0
rLefvTce64+2yKrOeoZoxiwvjZtqDLJXgGwdk+BaWW0mkkHIXGNiQRwsD79+V1YA84rnXmmVSubU
JNSN/8yQKKOSH3bCCXk1GS0RXz+SiG/hHyOIKzbAOHumr3h/1CE2AdYyrHJU4oRYyx4bS8a5KqBI
6NpiliQVVfi76kHpcM5FKXpaVPNO2WJpDFfU9czt2+6oYjaTuQi3ZDIgZVp7dQwfbjo0np8ulw2G
ie2WNyodk/FyboIX4zsIpcjMCdplIY3yuseED49Xm22wb5pS/OXHOGL53JDjKdKJB01SDpAtN12p
uHQMvZxVWJV86ii3h7JKNZ3tFhRLNRaTzcyom0HTWyHTuym/Ak2YXr1FMGYjRnni/p8t04CjTMUE
5HYTENByIiN3FWuJ0MOHeaoBYQu+wgHSVmVjKSolEHhbNk47q9x1t58D6M4CcZzO611SohLl86z8
+waMh/QgaXXt+tlt+PTmdJhiCOSfR05Ho5sX7UHeRTUe+7HxtReJayPzXUz7UcmvRSPLpe4TBWir
t78bZqyoGNAP2/bzqJ9nQmKk70in+3DhG9aFZx7LRI1mibO3MhekA/3LdP45XdT21gFZldAzCijn
0yhL/rBJdqwYj3l5LW4WAdvzct/6anwq03tGukSBg5Qx2Txmy9+RJ62gsklh82A1GPU7y9VfEMcr
bJyP53/PDRig44e1gw1krGV9GcsamJ5gOpaxEyUF+BHXN2/1J79/ypL8NhlY+MRtazcJLsHVerDt
hxWyIfijWoR0j9n04jSoarnzkCQsDiDo0CRPDOLuj1uA2Dr6tsAeGGo6w9Bnl6hww50Pn6zE9A/u
Ydfzn02rgSn25gXbXxCNI0pBCI7NFNDwmXvA3/tPqivjxyRuJjJyD0xaiCm4KjlnwwX5oys/mxPt
JeHbmmR0g9D4J8sGy2vi8daw8WDV65uxTCbcCNpiGF9EJjdqUprnfD22fLtCnfKQ7sKaBSyQjRSy
368qjY5pjR4cI9tkanMvPg7glto4Iu1z81kPJJMB+CX2oWQ/NkBExUlzlkdjhSGVhu9LOshV/INO
2WZSYEA3AKmKPDkDGvumD6s+LLndlf/Hp7fnl2q1Nq3pf4z1Eg3x6ckLjKR5h7Qg2Iq0rtgkJSYJ
LJWTn7E/shz8GIkpnFpy8jfVKu2OVEfhzTwKMnuJQY4QAJPTYdjSY5+Gz0kPkjpkGd07ynUToGKV
P9TQMhiz9hTIfsjtDroM/IZmeEwsBvSFyIK5RLgIjc+qQjCqwuobw7SK2uZA706P78ihrnR7GWal
73WVA0Yt1fCebe5TvQicj6G4iOUWRZPZJzTu5O4Pxj+S4nsbYHrj1K3pxuutSmlbEzSkgDRMAJeU
s52Kq214QH8huKLYpf/VU2dkPorcjUNB6i3duumoqkQWqBTB7K8kibGwCDUWCkMS997MloE5mbFJ
YgrU/toDKkoo1bjluKYhRWiAUFa2UL18Wsp35iJpAnyZmR+xRbo4upkOVNdN+m7CV2PniC9MG5sa
Xb2YJTQpzsIGZkbayytprD2T1Qr67m4Frtota7xx+IRujGYCRuQ4ROvWQH5FI7arBpqSqiWXzOn7
7QuN9pn9brQlXrrbKyuNWNVZw8k/tuq5ju8U2l21ZCCXwt7g2ApLs7g+hre7wlwnCsKk+uzXND6l
PY2oF4Lpi7AiIQcBvhlxRLlNIGsKgWvkdCgizUHjJOrj3BGk8zZyzJV//P2S9czNHUgaB1JLBPRS
kaLCz7CszpWvJot9XCv0VwCrc8j+N/Kn+IzmxjKM4pyjB+bm9wiqSdaWyoimwhF5JT4I0yx1uGqW
oTIxXQG6iCJ2yGAIWtW69yJX2EqgumMKUDYjjz8rCd4TSRk/Y1xIrHIs3uQ4M2nQePmeppjYw+uz
w2GQGZmOfIMfyN6LWVbjhCuJz3mMen0jNZlXtl/W3iKFcXIY7FFkZ1dCwS3nVhFUodreirbLaTJI
DYfDbQ+jW/3NFXVLHrwnqXKH/C/gOy35eyveMSQknovuXw0cHtkwaaAQ2bshqf1hIjYB4wyfHAuY
MrkGL0owWDuqkDNdPzDw8+eiWC17WU7P5XK6K5pR4BWEqfiGRH6qKwA+JiJ1d4J7+LxcPzwp6VbP
ofYrMc4rlyEIxnUMg3QclKLmvUJL7zlCLqyZVDyLQk7skxtGKGJy7XfppvufLXaOdm2T3BRAcRt3
5lRsHVvozNPZ31T5RNe+2Y5J2bxKTgBj4XBkJ0HuRtgvlx9QoQEPg1Bby1gmBLCXvYnK0WHNjVUy
C+2qwqR6MQO9flL7YSb4TvF/LxGyPrqko5nVtSwUIhHVucU1F9owx23Pzxc+TXhSW41xz80H2sSo
9azdjV1UUCCoeJLyIvS6KV3o8EqjsC/+ZQhxEfjFfUz28n0yRJA7QGv90xDzTS7wT5gSYjP8aoEq
/mzKKTsvhw2AYKH2ycixzsksvB4+cehgGjA/vw2J8O+7lBCRByWp9D7V3nhQxSZC6Ji4y/LyxB/g
VyjrVDjmOMPNTETaKmJjtXxJI1QFa6VzzhmMVpSQp/uOHxEPQDyB1bzpnxxK+Jrw4uPWhrfUIToM
+18WlZaVsHSLb3GN9SxxYH7G+wV/5Zicn67yeLFBJceR/E0Uk5g4tcGGs+QrglEjSENmp/rCXpcA
iM8T7zQ2f8Tt1jk5g2TuPMwf/pRSDCgfrz4gCLhLFCWH92taekC9SGhUB4VCpKV/znS0Laxw/4nl
VrKqtGQscpgAZlwTNbekGrYIMXY1LMDslTB7l1mwBWYZjki9edpL9uaGgQxiriCS0exDlFQp9btn
dRigaQKE6uAeHoy564JCKTk3/UQm89aYArrww7DtkIInfKIJ3NOv2gKFIHYhk1JwvVhVsB4/engO
+T/Na6WBtoPGdwA1ZuAlUb73a5GQ3o6x3yw8T3RORP6oKetIQc77PzZyXtvdoWb4/D5K1B7T/L2f
VvUQ/9n9eZIrhpBfCvvrkyGuBT5LGqYuGlBu7+PeGIgITpgzCXTYh+tpDUKsl1wSxmfdw1dD1mpk
7E8D5LB/ilIbJvfV3FgnB577aG8JnwwQhow64FJ5Cgxqx3hchk3m30eqS1wneLhfP+L2X2tolS0d
12dwbYErzNfLIzy5PY/ih+bDkHDV4fJyUdnjl+FIB6W3/CG9u0h6lPZfyCRc1E6DIFV5s1SSRmN6
RVA7RERGfI3bowMEC4NdgYvHwdI1yaCnpK4e6ovfS61fr8q2W1H360BCt80WPvMBwUBl4DbvdGl0
Zj7NX8EIBuROyIn27OZ3RwgAYS6KjxDAnTyFJhSs5+Q5YYo5AfDfnsM//LLl8mF34aRX96HiK5gc
nl5Y6sqjBef4dBKo/mZanXxDCzIZT/7wZkyC5fQOAv9FQu+LWJ+1JKScg7PKEpiRd3efgTu9PybA
ud2ctsFbBzxbWy5je81bJqpdZGGijtuuAEEya/Eaozh1T4O4l2HJH66Vs2gVgT0BuI1/3NqQXUxr
5d2vI21NPRdCipR48MSP07uo49SrPfPpVgms1RxTgpqjrLTcd6sRqVvI79CWyeq3eWAD6Bfx31Td
aBWk9M30z0lo+40zhVkUVMJ1vLjdnpFP7sh8y9yJX6/IGShe4Xd1KsjR74HLIe6YA8KkfSxCVqW+
4JKsX1kPY2ACIoVC2YIkzlErfcvWJjazrLnKPAeB9gH3MAssM1zpU9KsCXozcbtq0hKUexpDXq7o
ARSxG18MyvixN/LPNrA0N5uv8dgOsLoqmK2trEnMh/vJHRbslK22Gi72kDvJsk9bknqjrF/sUjtN
6phxoyueI+Bu80kRUv5yAuHpgqwJltIYaF97VIL66CHkXHldsWwHRhF483S7I6RV9Nv4/Q7VP700
wZjzL5qmRz3CSWH0XR40a5RHCimrqWc1+H+Nwfj1XNNCrjgTVcKzF+UfI9PsoQ9HkbVmdOUOmgPO
GBXTnpcwS3MdZwrYKacaCQw++nVPYSpIsXvBxNqdaqcf2RO9Uawu5ig79HSAGplJquZsGW8fDoZ+
Ebn7cMplZYC5OFuX97wTB4jMODHN6OP9Jf6nmN0SzrAI6vAfklqp8SgzV7i2wQN2wlffxHLzimf1
Al3ZqSbpkZHa6adDF8HcoSFPiOxXTrz+mlpxon9bgMQFlGk2h3dKXAKknP67NNCoOf1l5xiynT0b
avbr1ZnfUByg3eUunUBnbs8ucZRuJqEuRup7tjvDEYHCQs7/kP2mLR9O6Q/yn7MNo6Svs5GE6nRL
kZMPtx/jJ00ftuR00PQ+roG0gn8Rtynh2n+DVp+TXkw4BTWqAl5OmaoipT3wAW0aHYheazqRiG3a
V/hcg3IB3R55sllJdRbl/lOCPxWW2uMybJuryZbI+h8KVUPjRE6byTwO81Ij8aI6ouNqbaxMeoXd
jWizuVgaMy6cqG8vEyMw/oSd35Z8dfjwnqfyuAGy3kbpz8hpSXuLEhNAlkgfAbV11QRksOWL8SpS
hDU7+tcoGa7KSgcYfbvvDNIURvrBRrKFrGMEcyemgUNaPc+qaVec1R+iGWZqEXOLHzYhoiCVYHU0
5/l5UatTY3BkO1gY2nShAKinslInmDA8dDXbL3BTmhRIQfYjCIaGcV9BE1z+9AZ1OaOp7OZ5LD/P
Z9CxGj8fBLYHJruseybczgGjH1S7biI0NrYmBoKLLdWJVoBdKslt9vD+HTJ1Nv/2eTj5eztbymKr
8NLzFqY8iOg/qtTxJ3MlTuwyXBdySO8gEvW4zgRuN0BcqLA4N/PgsRjHAfebMm1lc6xdo1DS4g+a
iQfa5hi6U4B3qc51QGTInt72WTJ6fmGre4/5Ru0mYRHDayHVqag6t90mehW0xIVvX6juxGG4USix
oQHqwoW55W2U/aGP/DZkOjSoi4IoTFeJSxxkEeYsSQAETKcL3uQdqYXj+N40SzMiKc04gwZ7m08i
HCve5r9C9jm3fFLoaHv/3j7sFa5IzH4mXIt0WKiO8PuaOPdhfZueJ75+FM6jdtCNHj3geCTjyH5S
NIDXk6leCLPoXMUFbp56MPWZOwt4+K6T5MNf1VUcH7rX3dLdC97b9OyK15pGtK0I81ihJc55iAgO
iLJJqZZNjKGUi4zfQ/uh1b/BArKne6vQK3lmCQTKrkqBUKK3Ig4b0McdW+4fqjw2PFLf+NTElnMq
e5BJJKxxmEquKxXGXeY3e+th5xNF1ulNrj0Zng/7BLTGh3qLmpBDpbXSh0tsd0X5ia3JN8NTabr5
XJYhdM/oA1LutieEhPa0HubdGHtL3K42NGDrXcCt1GWHwFCwqfOgcz4Qil+eZnz1J+z71285J76a
kTU6tnF5AmqbxOctLlbdvSl5eYe35O2YQ+af2puK0Lj2o1GTUjvSd1HByHSmpQGhvuNVD9rMsAa8
SBqqUVGYW0gU2PHQKqh0yHTzde+WMjBokpcXmEC86C8Qox5rLspyhwZf7NJ1L/IiqHwrBo9ZGGyM
f3mQt2LoTuNGqIMNuVmi9t3GAvsjgDE+G0j0vlykTbvBi7oxzGtBTZFDgs638IeQZr2XorhM1r8s
3jIc6A+HKETNnWmi6uyjFpTtpGjJ7HP935JkCij+Dbs/ieXS/Z9AYyusb93cxXmkQ9DG0k72sJ6c
XeTXhioYj0zRgos9t394OdDGCs27ikd+5hbIqzKrIeaGkfIreOhLpQchT7MfbxZ4Vs3hLBJOnXLZ
Wz03rGeW9aZRfiK2qkfJm0nSnCTFCQIJhbS+pubqBsQFDKFEVmRJomQ9DuP+aSpuEBZC/LONH6b4
r4M2LZwZl99PAIGS1rpczSuAeutnavZCx4Up1Wq6Wc/FLyAAfAIDOHs7ZsW7oBY5pW/Gy4FKOdLr
coA3omgdm4qj5iAUiyKDMaRovUtGTIeNFKrooWYXAtUtOOsH8vKdwbKRX5zFiBNpSTrOGtRg3nhW
4qDc+/L5tYFRC7CPOiS1xrVIjubZrcsKBe3gG2uMy5+4J4ziGgssCyzBOM2Mdexn9NGXPBHsloXB
B6y71/AG670XbmVsFStMQ4aCuugjc/Hmk/g1TvsG6OWhJnaFd/rHTHtVmi34wJrFHeL2mTO/iWA0
MKyj0Bkzp2485guuHJXmDSPVXkgNlTeUDU32owdrX1/IXeYLrnzDrYfkUSI33m+aEBxO/LEe5xe3
t5KGEEDAzXxYaBsCQsa1sWY1rd601t4tN0RHsQjHFaV0NHq495u/lSRLGQT7Jz6B4HU4+RWWfXS1
aVC4YtpvxNJ8FZv3pwUZdLwNbIjzgWGpLa7jPNDHkU7jgm8QTb/GcqDDJrRNg9anXUAnbJATENzM
1I0lsHk2GOus4Moi5Vpri77deCcMuk4YJRR7fWxg8tF5TQZlqAclQnqEbC7bE9LARZvf4NfiNncD
tKcZm90SSt46b+Yp8DuX87S3NN7oqYxhTF/Qus/miZScoQOwcZ7Q3Viu+ZuMWQ2phQnlgqrcwVWW
DAxDdu0OOJZ5NFYcl/fWVui766C9imLBw/7GgKc5vkSApxBFkIQVB3KOBdjhpag+l5Etg/zVQp/K
2YUiKMZzVu3hjQE2B0uxreuOqi44eaO/IqXeKtxPrgF6njXJ+1Hs5p0FoyeQePFDrb8SRYmgyytL
zXkBvX4DHsnrylKWC4VF9fHtuTlDzOp8Nfh2RW+KCNhYIz5ZPoWT1UbRYs1+SPQUPSRjtyGHDoXH
QarRrm1Lti3F2iAFE2/JDA1B+Vss9vEX1g0ON6TsD1WtmFXL/1/YZejgQYG7M6F4VGfZgTBlTcHK
oO3SEExV+SzJxvPDH+RFi2HWqVQXZW8G+23Q3T5CeRucWA7oPXzhPEib6xXyggDG2rszChhM33JA
riiZwQzsDsGPdZTMFCKlJrv4T/rC9LbJSdis0rqmpCWhDflfEIB+iXeQgD8zV5hsxQgwGddcust6
U7iv0n5qFhwdGIy3TmaBcSjQAEVRYx5QFURcTXiOTHVXBW3R3H/f85+88T8eWBWLiU/xVCZnuDFU
Ofmo2a1Xz/hB9CY1mdUZiFqiYc+w2Zvdl9qnL5Aj1Xa1JyBHDFose68HZz4fU9HovmmF1azS3jOu
h3r3cvNqSXJlKnViL+iHtO232GZk1r+oFM7BisZGCylCPFm759T2wi9Dt0GPxm22TRTt1N+9HWiv
hoTqfBPfs+jfU/iYu9ynD4mxwC0rrkkLAbaW7rZGPvo9Vjr5z0AYDJdjiyX4k455vm0WKWIsPG1a
LqzNvjSJoWrsX8z40CacSCmiQmKrMNHKI1aAyRT7riIyLlVVOkk7AC+g782Oc5tG+D5pDk+C7rgc
orAJKHsYluahPXtyCc+xk/NHkDZdCa/t1U3lnyuB14BlGKUiMV8/ZtXIz1aU5mtkVVmzrimghcXs
opdKvVwTWgUDUKl0pjsA+k1FItmA7y0h+oBnWOtv35rHjEhty3/Dpa130q0wGy9jJa896NV5nd1z
zDv8+g+fcPh1g6DwdBDDiY0r1Bd87XAarp6SCEAgBJzJpbbgSpLEojLklY5YFusdJbEJStIWk8Jl
E8LtWcbvfTrPCY6DcsZ57Nt1H65KEb+lB4CjBsBc3zLCiKNRPHALX/1ZZehxsWmkguxTlsFF2EN9
+KwnOPmzZSNg2hnmMK7tr/gYZlO0awJynjKHjz48Bplui0GNicsJ9DSzGjTI2eaANAcyVcc69u6A
D9hubZRlmb7VStFpxHFVF7x7EucQNeovmrOQNzH+Yh2+Hz+9nTgv+ddS+f90vgv+bT9wrtFZA1YG
TbNiiWTbd51b1IvX94xGlZreY2+nGGOOqeq9mjFZBaCbb7JSfTklgSk8mj4+lx5CR9gJ5rncXUgC
d+Dj9uChSdc02s8+RTmU9xtf67h5OC2G/zDMrOP3L1+fsE6rGsfJA4mnLVnox9VBWsJwjsCH0BY/
bhRduWE+of10PyQcC63ksMf6mFuAkIuo5ODoXiuBiQSKF36z+bVhq6Zr9yhG6sv5+X4sSwyLABoz
FYmVxXbIn+lGrlOYlUtE41mT4G1IFjrD0QxzJ7pa7+fc0C4V0Zy0AoHhUVb+1H0WVvExW5hoLgDk
zoOyOIeKe+jigT9+BoaxcyeoEUS1aTqkVeTatovUw3iM4ZDX9pFYqyy7KLLnc4CUk9x2qkHMNoVN
FRw7+E/5tv3gdRvsT5v+wE6VYXb1dTnqDBQst5mQ//o8inksyXiZwZhAXbD/TeMRyp8Nil5OkoAb
ktgOE6RO5bybvgJSF707wt3dX8AdxOmVhRs224h/IxQUkUXXuzK4lZw4G4SbvnI7gMpmSgVWCesm
hmDdVhsfmqnvPsTodjynaCzIQmm3NtkhJlLTu+1/r5ZGdrWmEzSiiiUKTkKbnRGZE+5cRQVfq5vt
fHJSwq09zqh7IpgDEEflCsmT/KDwkZ7W24GaPkhcrsAgkoegAgxxFUPfP7iliGJC3FJ4GWS/HVMw
t1AuYFVi+OyYYXtW9vSfGdPuUnN/X2FA/xjvvtT+5OVtATZ1y+JS2O2AjLRxGh0Udja1QwDGEoOK
T5iKYT0X2rxJeBe03qTtS+2RBPcxYjKzEJ4j/TdBeut44kFe5bNC4hCDN9j21l134Y9BFrRntrxZ
olIykzlNWpu8xJbwFXVRYUynV6ma1XIEUAW8e2iw9dB0dRgwJbPZVtIwfDbVrfDPy2nijOqblVfF
Z1EidpHDzUbVYHs04FfIEWTO3BRDcPqBXQPTx5DlSWs7mZ9CX/Y3fi/BYL3QKyx42ksphPoW7nX/
hQTTcUS3/ZqaYorrkpQAyqr4XeSXWw34HuKiCzxS/F2QbxEIk5RXIc6M1ZQb/SUI+ZC1iL15QODK
Bx3V3/IbLiz6XnjJUgAuTYWPmSsXoL5w9CkX9R1RFD+gygzNnWPvuNtAv1uyWLE3ys2VeGyTMZil
Jy4Z4tdjGkrujjM0DKMMHUSPf4U5DgWHcIGfp2Le7tdWPFi5aPcMTuPiPPtlF7AP+nqIS3RgHg+/
KbWiXaxH7ZU0vot9NqCztxcxbgHaSrp6b9OLNWgl+3G31tNpEl/9Ch3G1xnp1QrAWZj4+bMQcS+q
Q1swnnlyo5ucuskGtL3bN9jI6jzi5bcXWAJTM6rqv7a0JXWNWlJudh9se06e0P3JXWZmz+AfA9cW
0aFH7kwJxmAVr4AodIDH5sTm1NaVcSYjpQEHnCtDEqlYxFwZ2Q8VbSMcZ3jcukusvCbp3mklxNpL
0QVouyV9CwTX+KcL9IsUAcM11J3PCyVFoSnOFvYHRC9T3S0odS4gnzmWYd0x5UXHAPrxLp8HPsBa
m98BD/Nc/gjwH8nemSl1kWVKLhdTC9KqZp9NL6KRrFcPda4LbM+Vf/GJ6ZjTbCE05l4nbJYUWYCI
hSiCR26IEjieRcSK9fqZ5ZpF08v44bBzsIwmwWLfG/QA38CDAcx6B2JSi4+d2ARk41tadv/gnLOx
j2gk4oT0LcqYJ52sHabwvE6N/A5SxqiDBdqiEa/vNTB6Zx4Blk04LEpI0JIHM4NhGf52mPnTqFTh
wuZH0gRJL5r2UYAGmzfIDJGYG6Zigy/X1ySIKkAu3Z+ged3tAy3rPY+2I/syKEW5/rWrtbYWlFV9
f9TKR3+S9lnDM6kYFfBFQwWSWj/sNZWFV5DTA58UB3DFourRM5pfowNNsrGOOIaJSdupMIOiBNkJ
Na8RYi57+aAK0U9IvWaes+u2KZUPL5eE+0oCaWN+eyWT2EOIZKtXOtNkWaAjC5Okg60wQtpaUq9u
Av+VKpGGZ7BDRdRx/MjVAbsGCm2hNl8UPRwfTYWUs6ELp8Yqu7tdD9wpqh/S1nas9LNKVFY4hKL4
cDBUijT35lwSVlH9//Zr0Y0iQOy1JQCZ9R3KwZOhmxMwapbWlwZIFPKs78HnJY7L2NRxXlW+eTEe
il3/DOHMv3iYZQlDB59TCTM21VzSMxUYGPMGoVa3D/T2Lx12X9MeO3exOzPStcW9euIQfRVOdTao
kQYBrgYgGPx4Dc0wI62dQFh4HTGOq8A5oRFMjPe6CQZJIx1Pa0v8coAWpaK17pP6O8jox66SGTEe
hPFSmhSpO1vFRz4LRsPWMUZKiQuC038qlLij96xO3GER712mLN+GXpppwUPRN88RdNXltHh4KbhY
bXFIS7gl3xKqOPH6mH2N8M4BmAlNFdUFIuyW6OYvQA/Od5iO42n7GMM04OzYMqsG13mvD3DHh4BD
6G0HEHhhpctwt4b60hkBNlVjv8sbVlP4gEpF3QKAEAb33b2RYRXFa1ixsEHoCj9LIwhT2TzNW06w
ld50u3RpMt/ZyiBQ/anhBhnG+h03hFxxtcQjUxTGlPLqZZ2m4fTVY+yGd5MObZj2jYQ+RfLfqE0/
q/2gcNR/2Ni/drlBxo4DiQBkNiSvVAOLVdriWl0rvKCVvBHPnC8FvZgfOOEaT54MeLeBWMsNFjrs
pdyYojCBEj6ovkU/rOIr8Was3iBv09CNVdnPTLixgzZ++ini+lmVrp4by45qRmkKQnaGE4u80qya
FQgA7NMM1lILTFyiuQNVNhR2Au8se4EmWe6JEldq73QV0HSMliPBS75SxcLCGWtpKlZiElujNDtM
b6YuetxtCMwxGoGW85suyc6p+kStrVMrV+b53IKCzdjBZe0JvvhPD7sG48F3luWnexxXgLBFXp3v
JAhfk7Obt/jX7AjxFuq+Pr/MPfo+UBJRxR1mf9a56yIUET1S6gM1r7wIId0BGdwu7f265oCt+UX5
NRHqx7v1CV06bPVkVfhAtskyXwHdHOKEsOyiWLuTWmXdJUFHxLD8LEG8T9pSD/fsuldFp9j4nxsT
/tATr0d8BwaqZUlHbnJ7qOoAgoYyTyW7W3zTpSCd6PxV8uygU6NTBn/ZsjXrFO2nt/r1EgaOMQcn
DlYX0t3gFiCjqBJ8qrMKLQHQQ6Z3K0l2SsmFiREGJVSjfTeSojdrxcrKJf3y+Fa99xfLiKKJUCpn
hFYuIXl91JlhZmIyqvqZ/+ENV60udwKCYh0fqhFfieWV8QUHcxNlGpdGFmA7Z+uiMkpK5JmSQGZC
DRv40gYRNQc6r+BGqdChyh4m2fCsRtxFGewby9BhaSHvqy0X/cLXAxDBlyIWvrEtIwhteB881W4l
drp3JivRnKFnASg21VXQNRjkRmMDX0FqLYV8Ej5RwvmPp8Ue/WJbeqHwpyp2twH/Z5QaiQoQcDIA
nmW5tOmk/Eqm9+4FwFn8ti7vKCJiaUOPe8pY0scVZM0DcuV/AIQnFkdAjNumSDQHkkBsuMYh7/Gu
Cx71brKscMwsynKJ4J5mAR6FHPuK53nXJ1uMDGiwvTq90QRth99nt63G677sJg/HLqomGWBA2g0A
3UaLVzN3mm00uryyn3zL3tnVioW8RBg5SYoX3EhIBGyCKYTpetbNwjjUzjYVyfEJaWoyyoXXaj0I
jG9liGE9N+G/UHbxhnuEUppuF3PdzgsILGBEZBJdqpcpYjarM/CSZ55LnP30ZdiiWxrWmes1A5yI
328hiBMac8ElhOV6S71FrWABoo9t/SfkUgQVxt6Ixu0OqLIZG7lj9SMtMubryF84AQh9ZtTPKgyq
pGOFUaReNFXBE7K+Kt8eufwL9xV5hK1EDFMwAUbjAfTEqRAJa49gXMAk4/ghkbes+bGVUA9Aje0f
cOdhP7B2GZKqxCfPf6YeyaxSCINcWcdFzVVncYPUkfKYq7p1W+D89bDW3siPaoWsNQSYBp55Wb2N
IZAd6JtvpWUQfNN8IvDVfAJD8M+9enTbfwaWnQcoJnovI692bIO6xKTI3k4WLw5xCYwi3ppjEZRG
Orl9c7Ci1E4U/8GJx4n84BP5xGDXAVVDbrGZWIBG2w229pBWh9GRO5dW5ZX7bmqStIIdRoR17/0I
q5urw08zp3rJQi8bHRoCwXFU44+QwRyf/RcBR2GwAMx7rtquYGEGoJsbvn2/heN81yC0g7JQ4MqL
1biDv7rAqBqG/oP4nhZHpzl/4I3oJ3+N2dM+8FO/wZP2Iy0dCvqIogzNPpLRssoViqEW6k8W750o
G1ZXXKv0t628k44RShuVR4XwG3lHHRSiucdg/Ani95sy9pHB9JNLl78m2SEuYyL8cBTX3GZh1mbr
s1JQTOFj8X9uV3FCKVq4m8OeFXCo0Nmgvz2mQor/4hED4Dzz9eyicnF9NHYmoP2mz932Dl3bUHd4
ba+9Ty9nikTboUh2fiDrIaxbAIQ6tV0uCRs8XIvY9gCvaISjDV64eUHtNMmb1+nHzlpKwHVQn2ux
hqkALCHQmqxlJr+5pVfFhsTMABfflNExQXDStJhOadC4dfQ/b+iiynuXXQsgTlvrokKniQf6BwpI
EjZ/re2OMzcSFUPH4V9fUrYxTqXoi5inen+ztgxPZ+Rdud0A4Yv1MFvPor366ZyN1Qd7O+isdwEX
nb9d58Jequv8zIUsDfKLrZDIGWb4Sc8YB4y6rigsP5tVW6w6mSeMYA7D4CPMJ8QDB/9fu00t5zpa
sO1nSEShZufp4hQqRsrB9fQ5v8UrGxic5cl7bm10jamR+3sWBNmaBtholCekx9iQ6PkLQHMq1U9J
b/9g0i6cfOxGGDboje6MbdMQnvZG24jKi2GZWE1xLsYNK02OvNKnlJIMDW9cuNH+CPfVale/gF8q
MgSxhV7c3xCOZg90xaZNeRU336KyE8Jq5Hgm5U8FKEAz/Au0i3takSf+vdu8iN+LDbgP8KEJKyv7
dyO3amNqT4YW3JSUtW5DCh8i6dZ0JL1fD0x6992D+jLryrlhSuVhkNgLpxEGFBwvIgEDTHlP2hlf
p97VHi9BNothYKBToB2o6kCrnFLuVQu/W4X1/OinBVWr5ckuwSB4mZbuVg8c2SFvHkgX9pFnQ2mV
u4XdbHOO/tKd0IMncCEulYjYT5c5n3yhTZ95oVnXRXOC+F+6USoPrJ0nDUdBmE/0G1rNjKbY07vl
3prdNHVFoVFIvgs63oKEM/QPadWLf1691+GSPlDA6T1q+RcG2vbPq/Ha+r3oC+sJs7Jy13+Nn9/M
1TeUHTDA1OAzjJQj78GSS/15r1oX5+a0j0/s43YbEpd2ao5OWW0vXqHThRl3wDlxwbRshaDqiNr3
0/yo6l4cGbn8x8pQuVBgaPJz+rKZqEoetHUu3ILstKSxL++qPaYclpWQrxtZKcgLg7iY47CaMdB/
3Yc9Ke+HVISTFUyRs2X5qMX8SnMrwfPrnX+px54/CIpBjjl31vZP3MY7bWKAEdDwcOWo9YIUVt+1
B7+8RbF8/lxfnmRWGEoMMSAXOebbsl3sb8X68pGvzmRHHJR8DydUDB1bosuidQUjrMAe5kzcOVWf
69nvrLptfKnfGkyfUT+X2mHlTKs1o8xOby+Kg8EwxLUo0RzjPbNu15RpMYfhQTMrdRYOeUJrCNyy
IQ8lek4lAvlpPzYSzzi6lY/3rOF9RcsMSmHsWLYDbpZVfiRCVxmRjDN8RR+tCDV7l5KQcQn5Vbkh
AEBEFxm+6mFr9A+H2HKSqKV31gIXjjuntPdOneO0xmLZViEig0/SJIBksgZuJTp7HpgzfLZgdu16
nOfTtDPKc8bSS0HkMaVWEI7HdyvAwCXXm0ckGZ3IygolgAcru/zgU3SJMEGu9uaYvhFPr+9S7sAD
P/VxcWNo+W6uIVWJjgzCBoAZel+qoXHpOChopTs/HQ90JZebBz7QSAhIuux6bqBzV8VqOY47m7V4
v3DxD6p6T2/ex+eiDn38Hqu45p/LIJ2QQ9e4ntvXjdwyOIiI2CK67Gl57u2jTiKAQOVRmoamTxqc
AowFcRjCtnFzDRkkd66xvCgsdgAUhM45U37E8hPf4hAKNcK+KkQ6L172Pr7cVQCgEEWkzUAWHo8t
sIgnjupj3/ZkGYSo7LiMFdP+wM3BhHB1SRfjEPfODvGSbAIxB0/LkyMO4fLn+amkyQVI3Nm8Jh2v
d4386cte/bYm9Jeiq5E6CX6TRsvXSo9eg/UQCpV1NiPkMJNSSJzbZWosWkv9/4hswHqNdXiyzxJ2
IQiU7gqtIos1hb3bNvgpbLcKLRuPNWaXL+1JTCZrWLbGvy5P2PHXiCtEErRSTY82h1oE5Yb6Y+0x
fqbGAUFVKbOc0qLvsTHEiQnaWCvhtnC7rNheFMIh/p9VGc1Tx3qeBnzf85Ef2N8xPUzxXwxR2yEd
QjI45F9e3J6LiD1+9Fad8envzeJzzMUU6V1S84Pzlc50cs0TGcFMRRjaY1ey/xOVRGKEDh4rhDAd
faxAopol3huxDBu+surCc6aYDZ7hhIBY6/CrMLDePXCCy0OlBuC4/x8qrjKmJtOMUjFrIxAiupdZ
dNwAXGn+C0naB+MNLrcHZ1ZtbNFrbpFjMyGWuiAoFoLiCoSUP/FajcxvNyyN98B/Msv+VNX3Bjdh
k8BpPShxFTUYlASmUSZrp1GIA1JkDxVva2mReV2kqaJKxhYV3zPZn7tV9STSAMuWNPmqvHs+Jsis
T+bHA95VIe50GKPryXWkDOv026sjrvP29H7VYqktLmkV458Jxuv6IWVtR+actReT3Lod+jrSrZni
s6zsH2BFjKt4uqEcMRZSkTpxxZx+fVi0X5gG64wCozR8Wrd4LAXU6rUKcZ2l1zvYgrVgZle+G8/t
O6zTenShpFzZJIriqdtKP+b7MRTTafdY/wBliZanxaqXqUpci/U7E6anWFK7tzr7RrW7ImNM4MKB
DBl1/P87ngaHkX0c/NZm3bIlXR9qjpiyUpM3xl24uYVyuzVbv9Ku5i5Gx+uXFw4ScIc6rQ0HM8eP
PVjG4orCRMXl4w/42Ck4pqA/x+h3EmH2hnnbcEyhX6zaR+/7CG7yoRr1XySSb1GdcWliRPAODApX
gjUIChccVZBONd2NJkR/W0ZRfwL5XLJJ3BoPN9P1jxnSf+r38vEYPS7YIrVcJplKQoVwZ38Hg1n/
WOsbeWJqYWxGmie0buAqPyMJc8XVhTx/m+mvaOWM4cfyzqKl1E50JNxRDUTF43gaNoCvI0D9mpKy
0Z4QOZ6fPinH23Vl6yq++sfEKihRjJ2Rbd3ubKq27avSC2e+LTwTS4FmpdWTm+/ZFo+xf2mAMcRY
Ejo+deu9L7NZngcEFT9BSys4jZAPb2wfa+9p1UFtxNOz7QEMyPzyB8gIfpbvDqG6pSHdTa+CcDYu
okRTmD/6pu8q/Ku378C/0S451U8M6KI7Hk5zsO9dcdBjr4Pc++IvVkUZxKk80bFIeyD1r2HMdOQG
f3wPHidSs3BVrNoJQv8z9KiL9lJvOA5vcm64F7FctTejzUCmjmX9b5gnZi9/yJ0YUhOp842BRyQd
ePpaoWKxCZj10GDkvrcV0uvrG2HW6mF8yXORJorn8BL1J9ox82o04e/VpvODr6JBBbuDCjwfCtez
EiMxliBfFg3fSHcxDOC3VuE5xbwOf5fPziu0kuVUPrrYKfDw5tBzj9huOEaTvutfr3yDGcsVD+/w
T0wWx/EhmoBDq9FGZ9Kd5l4Z3mZIMt8n56sb2E5mLLRmR2NEv2f6+6c58WwmIhHAneA1UfY0bAWM
7JlMJbkyUs4GP7S/cbouL40BQ3IaklQRhroVGnZ4qaM0TS2f2o0aum1BxS+iRcloDYiDTkt1tl0I
ILekCbPMO96HW4H/onDeYbv3mu6QGK1AB5cwHH4+3BcUClEnuPSrlO82jB65o7RXrzBWYuZmfEp0
76Ke/D9FKdDuFCA2g9lqZGcuawZ+epsWaw4kkF0ada3igs9YQHGHXdepDKPbbGCQcQv1jbl5F7ve
iIURerPVv8ldcmM9kNApBNwcIS0DoBuFo0Aej/flbU4hyfSCuBDG2IkAlY3ULI3qZj6KnD8F7kRo
flPdjB8oRNj7Z8PaXKehfszYteYg9DDVlG05qnXdRSsLrxOPIAsxtFCJQoIFKBwEalcaqSwOlTJM
S2C4dC0fvH5HeSg/ohSa2mXXOFkHQx/8LxptjMfxm6SsPbxOpMshM349kJW4qB3ZnvMSP1JIKMfO
fpPhtfT90A8YrpGSDyApqjmlUuWivUic6XnyX1aP7l/6zR7O390DeFJR2FVKwoDZw3kF2Q82zCi1
nfpI5mRT5k/iUIXtTrvwN/NyFG2XXvupdDeiaj/RMjcpSebqugOEodrLoB9etQV5WDtnkiKhzF/I
Oao+3eBxJL01aoXs3nieiun1TLWcrQIs0bAevUJXqhJyKbjxf5CTnxTR5wPKjXd7FFehpbUDLElR
nuXY5PiLz4RCWaBC0hwXVS7txsn6kWGliBsfRxFYKIS1+j01ERk0b9/X4Cu6+0Wu1B2wIo0HB+w3
sSBk5yfYoGVcPPlU+RIYEUQnU4Or+V90mvm2szjONLdIT589dk6jgJOUWjhKzsuATp6ALNU1LIIU
WJ0HM+j0a4eUKzNDuURSwN+xxNqsvq4Dpf4tQsSCJ98dkk27TnpRwNEbyWEn4RvIrvX3gp/UGvLP
7yvBB/wCmFJA6vkVEQfauVYa0e9HqX3Db8fNhXPvlRgM3MqV7CWRRvT7L0e0HJjJtrlWV5UaYRKb
GK5GgulDgal4HiEf/y2g+A2ctyu2/woy4JbIFTKyRy4jWaKT1oZ33cq+QWsZwc5Xpdp5CCLKU3X8
tftTsId+n227ut7ofN9FxqV16tWi/eFQLu/usmM/KwucpHHRn2zit8c6jdqR4fbRi4gXX5rmWpss
UC4nxFFpzziWGo7DS6Y+ytWn4CIdriIgnbFdCXWkujuCJZth/hVaA9IezKvlg5zWvcdO1ibwAmoC
wT2JOWnQLVgeMGi3znpu40IWg7fvhsZlB3Sza4kMO5up8PVhsUVt4kplhuMusGzgm/+dY2Qkehab
xuC8KUdiCLqEQuHoth1NA/dKuTVLPOIEGs95pX/VuRZPKIWVeiTZg57CC0gY+WbCVBbgCpck3a7i
XKdQCvMjLjZ/slrXQZ+f4e+/3x/XZKujFUW2JjKn2Tm4rqHwWHG2nA35thdXbGnhzckvmXi59wb+
ZemAR1dZTkVvG8olyts4J7TqD3OtqYzjOLiOKSheIjxauSFILE7P8CqjPY57mxy/txNW0ulHdgyC
pWUoL1Nim7WscQ/2DIdAPiF8GnAxfPDA44OH9HThEF8IjiFO+/9hMDrnIdExzssCWWOlBw+rEcdy
/EoIpNgQFcUSSKcPNTQ0XV5prvV1AfuxF/bMYz46dkZI3PsL129+mQucqKmn1vmsF52igbwD97iY
jfmA5hA7/A7MJxAIG0Vb24JgMlN9fo36RC9Y2T7oKBYphcXn/NHccGkDXFRFxZWWLT4LNHauKZtU
dlrIoXgBtaMYF2k9SJRz8K+Xx78b8obJ3b1GlNeogu7FE+rOlvXGvFr5BEH1isXCCc/UPEk0uTkv
zIUK/izdoJ8lEylQyiR9cn9JynTVTGSNZ+bN7uQWrKsesQnc2kvMRIvZWlHhSvlWw7xlmhdJ69uS
AUyVSSi6ragRy55dVQpdkcrzxo4o/x09iZVIqbdFLN+VcxmyVuuRFog4hFvCEchWPFoATI3Kh1Qi
uHEwIsyd807FcVo0flFLIvrHLjT3uzkR5YCYbnS+Jk2qHT4LaKz4hBWX5pDZDj5bF0JBRAxDJtBb
UCX7ulKyfeyDUr7BwE9BfpqiUf1oBJIbindpHHYKFK4VKTjqsejPBwVkZrcFkej0h7onJlpRKgs5
o05FsWMScQEmo9KO28HfJcjgzrJ/Q+txWJYunrUh/GqCyMXlqOHEIDbF+gX7jCJK36ukAZlI24eQ
1QmAhS9MCw6q7/+GHhxE5dTGJOlElkvQVGDPYahAPSZsC96Q98pU9to42RXmoGPtU/zyQPJMoaM0
gHWMZUf7m144JAJ+JoRZQOFPqdkdgP3B6n2/ntQZeY14uH+G0ILKNNpm2EGxa5j/qum1hbiGD8j8
+F1Peq0WHiCeQhTOAKv0nFImx/L/EeEPXfa/vvjCZnvh6JwTaEd6sTexf0s2YD9Sska3kTAYoTRt
DVlD08jWaWAA2vsq+nbt1jZhio+tDV0hW84AwzbET+oaWrt43CpOKQAx4OzAMDT4CAigMK9XMlBL
MJLpg7Yf8Y+NnjnrRoNjGgPy1n+mQ8++rPdgHdZof/6mcRsFTVRG2HmSEoUF1ovWIaLQ5tUl+kk9
6jshrycwWOW+ajqCr5Hybs0AOyVWml8J0UUS0Y/G/n62wdJMowMKA5QN8Dx8occeFFszPLnIUnNs
LYxxTiPhVmxAcsqcJfnGvjpNK7cYwDSIiVRH6lgHkKMeTRzF88wrTXqk/T5XMwd1j6Pqgm9nbf8I
zUfrnegavgrc7lO4wE0FQ+irfGAzDFRu0Xrc3VKvagR1U7+t9T5CnorSEceiAr69sSieL6H7ieS5
BGgQdD5Gt2+JR7r3qaIT7aeq2UMfvx7PbY3r+DwPd/MDF+YWOB9TGsA82hsp4Fi/65pxWYzlqSBR
W2gkJSNNHycUfDINSF+6CjJFlMIjXTF+RCE9fW51XVVNNdZqoLPa/4pNFv1S8nqvHzGJciZHkNCs
VD9qtI6eQbHGwbICD9Eo47vF9hwH6LAtiV4ZTvm3no8ljm1GCOCC3qNpWXwFXq/1oEz+zGeUwS0M
Q4yvONXSKits7oFSARn89GQu2grlN2cNYJuRkOTSp6utYdSu4ecV1GUDpS1jR+7wQRXItxXXcOOR
8T+nhYHz3OFBcpyzP04EaHmWlUm4PcW10wojM+p0SO6iH3NrPzycweerR1/fFX/aT8mKyuFU5f1H
BFt3BrC6KvH+YJUKCcxYrta52k3qhNZ71DWJKOxhPF+s9npiZolGnJSrB8yxiK13lzrsyWWQPz54
F3GsRFPj5ZWSOL+Kg3KiOJssFhzNFwsSFeMBw9zt4Y125tmd2loC36ymLepH5eu2e6M4d+SvmZY9
jXck4uk/XGvlc1EYBz8DcwzjWADH55a0mjXJu71gpVAy64HYiZM61XVIIBjjEaQzNMjat/js4+CO
CUZ08srhG+aqJm35NUvpMPimPk7yma0KsUdc33ukpHBINv8ptUmfxRK0r8aENqCBm3LNer8hdtxx
ZyD2GW2DmeeWfinGuJAgDrdGHnbctVSVHAvmQwE+iFLXf2p00CT8pd91IgK+DlmoDoX/bDNltNte
X0mLGbYOUXOz4ZOqqLb0eYXqGVp54Yw4bHGD2gtoHfu0KcIvTm+SAzXhSdSLK7ku+bdniuywCysp
878h2OJmg4pTTbm3FCjsqd0IxQMmARFh9ylR+Dv+0FdaWxXBKnBMBmupHYVqOBxrR9oKmpQcOlrF
FhSHBzVacrRS5dAyFjJ4F9rOd6S/HyeanR929FZtD4CjR2030rGJzZGbwV3r5eL9iWLD1VBrET4G
haDoFm4aFOKkCZyVdl76EbCx9ch0DcbACI9jVwRXsjXeCn2ydz59JRwFW9EZ0SciqtUSXWndi1ja
dOtEo0lCzSpekekOCPlWjWLveVPaCqrUooXN2zPRB59VUUfbg3ByKeCXxxSJr/b7wBoZQXCxSG/l
Cvga9uxWr884r8r0W2idm+3ErIvVNbL69j6b0nKRiAH2tb/IEcvkc7SzmfYU0pkOEVoX4Fcil9Ed
QAy/QlK9UGwstRzBeCH07C6cK3gZ26wljlCPHAksS9TqPiUP5ALz6zwiZ0JW9zL1TMS6NA1dgFOv
msXwN95Wna30MQzM/UjmPmAViJjxxHUXsBHAzw22vfJ0l3LTSNIuTr1fqcugs3//0N6GwiOCYem/
C8MASY7bf8FeT3oC4cYZ3+6P0olPt/HsysPmed31WVI/8kJcSzfPqkQIQIEKp8Lfppdk6FxMmXV2
guCtwA40CzjkvQQnbpSttb0D592NF+qFTTF6EAW7kGbjXrk3VnJ41Hv7TXG7EI3qb2jmN9ckgCJk
U5WN+E3J7tAf5gBgKXeW4z2XGO/nBj3n3npCZymVLUde7aCrcJ55j85T2B8qYi3uoOr2eWfufhx5
QFH2oqdYrJA6Z8t3WODqucqiat8GlNLV37rwtIvCDI3vhv5Jbw8TzHhtgdLtv2ZvdQlaewoD2VhC
msW27mPkXHFYLu6b5y+mKYwP0zYWAxzX/gkydduidxZ7E6SON9VRRn2JNW2K407q3x/DvaStafJ3
G8dnh5hJqQg6AFc8kxFrTn1GiMHIdhBK5fE3Qv98ZMZuSEr6Ddej/SNPjupVg4ttHPXgO46K84ZC
ZCelWmII/0pzuojfh3MyXyccYlKG8GaxN+zPeVqxMGWDw5p1j20FWu2bxjpTt/rugTH3WJlaAG6d
ZWmY7YC1vrGQX5owkileeefD/vBHUoKQ1bkbXkKBdrP6pNzfdlVBRZEZbhDDxiLgEnljIACmcizI
p/9MkR7ShQ6FwJneF+lZ4E+LhclJUo5iizrxVS7daKtVIEaKKpS73uEFplkUE3K7lbSt47BO+cwt
gH8X3YBdbrrDce987bvdF7PI7/1FZIH340KezyiDFTmVo3LxIMOSixpqsgrd478dtqF0ZPtzyeV9
ZuWghJA9ZNulj+H+Q5LbujBo8T6D/0fv2gGYyozlP1x6nanCaXic12pKSs4rgJPJCSRRL/52Wtvn
knWKtZPWY6tIp7q5hTbKafN8GPiZZ0pIyipIHBzwhs6MajKxjd/Vf9QTyv3r96H57dZX4fXIzfC3
8sW0haAHaDDAJRt31QDlaDa/ZvUfASOX24OzLdJbhkT21u6CcwmlZukguhn9AvW3xtnN6hXoSf6V
vRakPyihzMfMqEvNceMFMKy8eM3b+BD7sYNz/inlzq6zJ2Hb/xSqLxVgUSk844ZBmBn/GMAou14D
ZTiIaj9Dzy4d4GKbXsIoaCIUsDQpXofJqx1OAzZN6TVjudfqCwZ6wxoBL6S6gw4Z4F4MYQQ+Q/Or
N1bmASCwmQAL7D4Wr/RxjZt+GnOd0FlJGOJMtLCzWKaPBqo8Fzrolp8G+RWvyUdgpRBqxoKSG9AS
CPgvsmMV+XFGhl59we08yt6YLayuGTH8lsMZM2mQIJoSVHJWs+18a+pQ/Owi+YGFs6ZU28uBxMDv
Lye9+inJEruOc176b++6YFG+lHiobvipV/xttGJ4CDe1BKh9buuhyxe/kP0B5YzPv8Wh9D6LkQvd
d4rR72GRyF180hwFMOWu/+/YOPnm2PgWW6awgxAqSKNwTO1jOUXU0cu77l2Z0v1Hs2DA/h6bkcEU
IvG2AXl+R+Pg69IRoMe3kSgHDmr+xKrbD7Mec0NBDR+kqDgC5G/y12kaGIak5gdZNuWR9oVrZa3q
lLeIPLBxfUSW011CYxF7O+f0IUI5DB+gCb7XksJk4bAYw9I1eIwm3pu+UrtydqyLNeMc21AEyeTw
MCvmnobYbmpvCJb8uX/QF5ZKmYjx2ONXLUu70R2/SQ/hmYmmd4smDHkYedxKXsTLAGPCrzusVa3z
akgcOua8dpOUUlHkgZA+P/XE9AXUkpQ2Eb+uveOCPKnBbHvPzLp6qlrYXIljzgQvAHXHhYwBj+ea
EeLhCV/ZvCaUfvdsu/BeWKmpkCTV/P+fvbKc8VKVbIRH4OFlh8+/UUgDtVjUbRbBuRy2c9e3fusI
p0dt9MPFf9TeGe7uATkuYnUVHrafE0oJoS9Hntgpb2sOBKbFiS7ZuaB81Z15HqlApLRfaz5fmiA0
chb3NJQpWIvwP1jxIw67uLF8+sEo8yr0fwwLEEFyF5FqZ4M/2d3h8GHu/Ve2pkitTtQqkL8y7yxz
VFl3qsP76bcxj/XtkgnhS886a813s0GpSJ8Buptu6VxXyyitb36enmvqbMIOmorAZeHfANuhIx4a
bBLK/QArB4RQ+ZMU+47xZUEKhXNuXOTId7vARNoWsxzKqUtwRVKUHnPKDvI76MYi03f8C13XtxVz
DpXc7M0vBagxnLepoIs7wcWd7K/Iz53vAy4Gz4eFPRPs38+0ySX9oEuMCaHotbWpfj8oAQmsm2At
28vmlXEXrp/8slPiN4m3PM6Q25u8RfDizym1FP5ULs2IzdmLMHDi6ARpjwVCyGBcVToyhq7IEQRS
4Ic6opVkT6OZKMparTwo9gF0cNj3tg5vs1SP/s7YFYl/JWQHUrVUEM4Pqd4vJbaGTNF86BC3Zu5e
wCsbaMwutgyqQe7unTaVzYQJN24JHnt1/xDz7M4SJ3+CiEq1caIN5VxHiEMCsE5dQvkO7H3oYy/y
6kPIjmOOCcK62vCPwLoI4PtaSd2QS4Xp0FbSABRZsg3XrVdExVOBIdUjd3OKUexExLEzgT442+35
UvziMp8aTboW+IEjQkO8gefn6yRTQB+ShSuE2Ii+m0/K9ClRpcvy9f4EBWZTzsKeMIINXLSdah9D
WcyxreQsjeZFPRFs8mcDqi9lMUKvqV5fWxlZNDYq9tR2Lu1G3XZhNevZlaNZo8SgAMYwqQQQAVvz
+tEabYJSxJEk4WjIGcmQcSiTFXxa0wrX7m1gqPJiEi5ClMT7Z4AQg8mE1xByYC8TxF6fXCGLB5/F
cIzV6V+t03h7OowA4YUalCcn+lewaZKibhG+toBUDyYyqPOblY8RWRvk1ZquQoA8QpP9lzkSv25g
gFd50pPbtIFvssMOipQK4Z278HttFOXB5JE8bHA9dTOjFLRr1htQJQblYuKu4tYkT6XVuPhOVwuF
T4P+kFWlQqs3t5uDRk+9S9H6UT3cj0lstJ8ANHWVLP/zQAK1lh2BAzZU2cVBr+JAHjhg6+V7Q86M
DtXOeF2vVhX7ATlFBACH070Kcc+EvMw0LN1ugUmylQ1yzTlgbT1zhvi0558S7lDstUDyPXZO9eVu
1HlOi6J9WbHt6bp9wA4AbHv2+WU5TDko3k2WcF3gxzBCH7AASCvPt2rFAyikY/h9q++C5A7F4riI
Ns9GQJej+OisbAyIQPuREIfTOutECvuRzWq8lMbnvlFVBGaX9LFjNHHI3KQ/rRKLH/mKJx4Gsyak
W+0e7YpVryudVgCLchCmJorjL7YXVKNXEqx+rqkpWpD3qPSRJud7MhnTOs0L2F5tcXuYNrjqvQTc
SSLbVXHmpoCLW2EVe8xAszJvwJqygPgoI0Y0pD/PCQXf8Qn2vfGTTRXMtXqo0K8GPwTLxvGgBGvI
F7A2JwwDA99r/M07CFX9j0X7gJ/evihK5OFRNmZmL5OiIFKAxkvIAjCO06wE+n+DpNRq/XgIZua7
P3uS74wpx68nAE2gkKt+wAxJtS/lJHlvk3+vH76I0HWcqmApqdY9KJaiXp2Eix8JWB7JismQfgsT
AgtsVXoF9PwLDay6zM+KzqSxCeeX/5HYvjttTyS6bDLTod1Kan41YTxJPPi251Tepqw/+xgzblIq
QnvlXUK+GMvSUmA2k6bEXMJtJgn9fM/zdVD+C/B1SOjfPfSys3GeVFIVbwi9CCYwOdbS94rd/tFL
nLpriqPK3BPerEDFfKMXXwp/h4LvWANxBBxtgEXEO8VJeQ8N+eTGlWEPD+sCxYjNr5AVrra8RCsJ
YdeF0p0+BCXQGdOd6yyVIKqDmeInm25HIze9+BfTyQe5st9Ai927TgoGFUqRMdYYWJ3pRcQDkRYM
7pqTSE/yhxZeZ0N3im5l73GHM1fnFisli/SSvytiZhEG+GJGmSipUU5Fe6MSNIEhxXoBdoaybSq9
ZdNzXUpmU4Xnc1b9H8l2l7kdDL8NSsLTiyle5ur9SFE6x3PjSXng0ofcmT/eNqAFJrbRxy18LzOX
ugB1aYIBXZTCYz2vr/jmiGY/AV5/1YiJTO/dTSn4gMWjUb1HN3kuP7qTvTKDUw3fignxzU3rvV5S
XsYVEvYL3+HIeqvwcwBKN5zVMicxzZYquYRD/V7+w1ECsxK+2WXlpZHdOwzSUwN71SL+1PxAy362
PqqecvUNUoVOewUzPqMR3InxoAYQENqt578yCird8DGGd8sN+nGwRCtJ9l4LgaM6b4+I3yeb3uhv
3m/QmYH2zaA/Qd9qFJj7P9lEfcVmmOBOIyEK4t/yxicZ3hiveY35B9IC8Finp1V6gHOgjSvXbGrF
c1IrvVj7oyWE7qpPz+WjygB2zOYYkrmxYLuo2IPmHRjDIlIhOVwxv/hlXiLiaeMMFcQTXqpDqlOB
pdKj6Fi1EBM+Ezhs3YIdiw9pKdXnNeGjxhWy/qyQXR0VZln9v6cKn8/tGqOFpcDri/wd4q0xfePO
mkx3FHfWgzLe1LTwGD5t4bZBVno295t8gNdrSohhZRvnWpb7fk1AD2e2lk0SUKJE03jrzM7X6hHG
1zdZkKhDi1ZzpIYT/FoBVG9M8lSpNcvCAvhiqWq4NtnanKxV4dlwU0ifv4+bUfHSEw8jBwAEd5Qo
P5YdU3yOSxyzCbohlwOARk0sP8/KUdXbfY6O7C3sZ3qVGZsw6ugHLEjTcFb9uiDCZ+jIfKkTxqHt
Dujz+SWia5X316KyM6hDFE5E3gHWMdtklKvGUDCvHJQXufj1TSiPTUrlgZzUBNTtdbR7xcMGAhPZ
eqH4TC/TRCHzUl4na6proEC/UgIYLvATbayIVwxNgNTmkWr/kgKEthuklgsMIX3IW/MfQ3Sohmt/
WU2yIE7VAsB/lNmZeEHuALPIjdw3Reu79iZnumSP9WbBCC7brP+CdW3jkZi047OLDx8O0NMjyh6V
MOrVM7/VKEU1u96YBweajUKAS9Azy6W/JL+bYs1hIAz3zzQ7+i17nKDtEiEQQtiKm9Yih9mJasP2
p2tsqpwkW7ooXQWDeC+D30dEoruJD5KkQEH1Z8+E2NDJ7016NPUTZKS/KYUUGDrQnaKT0gQ3EtRj
0PGdcD7l5FiPN/I75A431ARH+nwH4EYR9/1mocK5oTfJKWbLomLN8c3Rve9ltqEXuxBJKfH3HHLh
Sig2L5inosrRz29BEuZ08IXMsFMoTyizA/NVnDd+KMNMV5Cg+X8r9jGbRJTdQF/SvDYE34uZL3YE
ZTzZTvbLL0VTypQbEESrshJxkAesu+l8+gWiRInvkNDq7giXK478mciov7ADDvkpek72mrUckslR
SUvAKqmotoiCmOSIkXzA7rJavC8paAmjGalkA83RiqCueMdOgeaZoMP1FA5nGNlXeR3EWt/pyPRz
OBBenHawWFTj9N1a4kMlOU9T3c+UrrdLZS1vLtvpRtC1vuJhEEZ+Qt8mM7jyk3EY7wyd8Vj4+zAY
0GFcxnIJ2FN96SAMLN62kEaCzhaymvpzsA2TPL8HHFItvqh+eTF/XHU7nJAIOr+tv4tqH4PjF5mJ
tnjL1NXC2GUovfjPV2C/kkOlrx0bsWoZiAATTY1tdiepRtRuqyR2lQWPw7YEFUKpB1/esAKC6g7h
ycfVYAhUFJXjfaxKVgMc8LotrvtzIZc52TpLRXxgRAXJUe+PFwcXSfeIfC5a3Ze0+ydta7MHl0jb
gMfROo7EzuZWktB8SNFW8MXfsJxPhXBjY66ICu7KH4qMyFZwA9gyNK643GKgRHUXU+9ZMIB4kwqI
OU2HXGCfLgl/UkQ7JhRM8lqCvxcv/6RTcaa0wbOBv8Po4F8e2HahtjOem5E497XZDBPWqS01Ysyx
iRL5m3Q+QLypJ9o676Px4IrwXPLDoNX96pqlvAB+59kKw2GEeeZNODgOrh6MDP5DLT2I95VnsIqU
X77P9jALjuD/zoMss7SKsvD4brRpT0Ag/EKFXyesKlNcsWb/QI46+rkAdrhEsmMlOCsfNsVbfus9
ma12irKowA+t7tfKSAhH6S0TaZa7RqD9ij6nsjBN4Ms/DMp4naF7u2Z+0llh/kNzcQX+9VnuLU7x
z4ew3ckIq2+AuqGeJEGmNyv29z8kotzH3TpA6ScZikMOd3xTUgcSx+YHkCBij76Ars5E/JuJkUk1
y0mlPgXtR4zsbJU/0nDqBt+kqAwAmb/9fI+GHn44LxtM+vqXXIjqbN5zm5bb6vtBVZp4sZOJICsl
SveoEpZBpZ5GclvH2KKVKkpp3DYiBaFZfdi+lZfeSsWKpsn0gcEWy9t9F1JHnhVosL49o+un0kGq
1uYFeapqOXVv8Z+mNiGxkLAj0e0apsEs0PZNr6Qi/Z9B+l1Q2TR+tsXLc9jL0OCudjffGO+Kx2Wm
wTIOewv4JJ/GkB/0NFFhH2QBlyGsLuIprT5IFxLX0Voanz1uVCszCaJVkiCPmzmMgWeKpDlCGkhI
mQIOUAwhi5KUssIGj1EbwHvw1HvL0mrx5gMlH/I0Rt/OP27b10XrIKtq/Nvy1bVl4THjcm0FufGP
GgrZqlxSy2KYRhnb3LkL58fwL7sAO7u2a3CW/uN+WJSbdTlU/bu87aIE7tgeMDEpbVKMlUZUkUUp
rmrgLKs5sCeOx2ts+1pIWIQTXOp7XxDneoKGQ2Nk2ZBuBJQr9yEeAlmmmebJ+ssPVLEODtq9Vccj
XpO5su7dcXiy1VE7DmayzjKwveZE0iLhcNGKXcb8DsV6V/NMRCJYZpB8rRstwXbEo9dS9yFwWsMu
jqUu+rGiLjy2gx4eh+y/3JObSdMPK13uNDOULSvPF+4UHSKAqNpYzV7fVZvNgHIwDtvnltgUGwga
LgriATRom9Fnw0a3ZUqhxbjcJmzfikJ5s6fXQCfegtsMQDtgjehHHEP7MqMcPHAWL/HAyCkHlZ1O
YGZfq7Kjs7Hlncip2dAKDGiMgzWaoyvx/RtmLvRuRe/ZXCkuwV8r6Sa0qgdQfATcD74ErWhkh/iA
MyrwMGEhk+ZrQtI2XIePfNZtMRIUzi+j75yPLArZLEou7+MatjfpxaoxMYVcKQZ7QHo9JiZa76eg
Sj2eKVh7TqDsWdU6gZCTqhg0rBpd0cpTbA+03KSUbFao634ybYmwzCcMF+9Q+HktKS8cAKAMrgq1
H7ZA0ftPSlptYN7z40LJbZFfIP+dcqBZIOiapXHk7zGemoBiLm7vd/IKvSL9gk5jrSToAO8Tf5la
qr4INA4+FMh6+9/s7g3xiS8O7/BefaAumX3a8Y4DkprTP/IztVAnobtj/3w41Aj1hxJcwQSM4f7G
seVg8tVRkwIG+g7z+mp3PeMlrf5xmZcon4lkhvfQjCHrnwo6bItnlMD+X8xW1UCufTFIianbNRLn
UBEowPo1fOs9wN2P+u2uyEDT1FYI2sDe44RPxmteynpoQPbFXqPdBc0xXz0SIr3TG6ND1zVmoG1v
SXwCxnOynxpfoVtaf5RB0qzPOrVg7iLqo07cw2pdGqZV161MAChhvUWrXQK1sfCpSl32KLxShAkY
B8bjm/ajorM1VsmV3d9ivZ5x9GXMCiEse2N1G5Ri2PWsLVvn7jj/xcu6OiKu6K04bf1oCb4iO0bX
5oK7q7vbktZSnMFROwz+PoCyuJfVYHD0Px4fDa8ar6d56qUlYG4Y8lJwYN78UQ+RfRwkpBfoagT0
sI0FfAaWOQj5TKGGlNz8L+nEI6H2w3dl8m7/64Gbmb9fEwJEqH3ERJVyVwBdo9KD7KBk5IRrMLqu
3IVCFKJRZWAXRXuUzCkP+KFmSPSPXGKH3x+AORkuhlPDSUwCOh2Wi5iLzft1Fv95Tu0qjd1SQP3a
sTFgr5OzA2hr+vJZDLpCpj+a4JWwPtHCjI01NFHtzr+2tUxSpe1p8fK49dRu1ysl+zzLFoMqNH8n
MtNDqIDUaBCNo5wc0ruAnCo9TwbP2X2gFiAcYBcEgJ1DRTQJnQRpATOqavf0/zPguyZC4QfQ7khR
sNcfYT2elhIKA5HG0MTbsbZj8kvxLfr3Ja8j5AoY3cLJzfA6tRPT229ZLyH9y8PT3g+m8fOs8OhF
SHtE3hpjPx0Hr0eXzH/69RoahPZBEE2JylMyR/NzOZ5nbV6CEZUerzj5DnV/Ju/e5L+zY0y3X9dz
N6QzprfXZ6vwJBj4/adV1iohRX4puEWd15ggPWHdFuOvB6Z1lnhgGDlYsEZVdlLGLse33BhHISAG
mmC7lB8ZvAcWi3+Rjxhs3rXJuHG6TdbyRLDzYAVVl5RuUp9e4nkP85E5Mk7MFevc+a2/Q/9CTkeI
DsydVDrDA8u53s7TfTcpuf56FU6TkRGtAt0AHwga0umtNCYkUkIlszf5I1E8Hr28h2M5pKHGR6kS
6kjIhNxPFMpiO5tKEXA2GCsIk7idI1FQ4/jNZwa4MsMyzN8upw3et3ZL4hi1V4adLCiKdoX/gVHw
q9Hk64sWMd08uuiUbukH2+hDTRKJ4beN7Iw+qMhQqSpOXnOZ/SqJRMmBgy8Lh+prk4W9MYk5Kl5r
E1eHVI20rLXfMaEPGxtmQA1rvqRS/2BK7aXpPsvM0BMHRQtYpYO1m4zdsmtLSfGPqp2Z6uugKJhr
JIZHaq/R4//jPRiEPpNFHX6oKcJIfXeLuy+ZWb6IXHighEXehNaHqCB+0bwNAbU1HkqHlkrdx4ci
FcoVpYQo7Ugm5BK/g7AZ3UEVz7DpQjFgcfbnnF4f87t+gQU6DyXZVBKxPB2BFuqv4cEyjAVqNYWz
mTrFrHuMRwyRgnTFkHH/Bk0o5j+5u4yIb6gSDIrBezdv2E0rAhrH6MbKgpwpoyo75TKWZ1zQA06w
SHWTgzJNqQHmR2hzb2vjGP0hl5HII6hYD2HommwAQUgPUFbCW4bGj2d9xXWB1dVgKSWiCAlTdOVl
PZmtNCQpJEMtHtZopq3kUqwJBjDcM2CzwSyCyxxcIGJLcg4ESHPIrf8aSSq9eAHf1SOqf+0Iq2FF
TKEWT1lk/7t8jh3xb19VwX9y86sEv1wIXF39fXVgIXyWt2wsF2sUnBgJ3RQEFZzuGRzjWfa02ZGh
lIXilvwksh7Pw8rjM4ltgAd1evGNWreUXH0lr0oXiPmNKJ9sWakLszz5bfcZbR0bKGbGFFJoj0rH
a0ax9YELOUqGEXVOJ7H+XM8laSx2ykOeu0y2/Shcb6Hsltqe/LcDcnaT3Ov8n9AqTFqWJQfkOrPH
qD0sy2g3pQFCfIm2zI+oLxiPxUevYwMfC0nO8tNdKvqTcxZqG1OLFhM1MAtavAQT6JU1Afzza85u
KYtW2zop7sKUikC3PdjooaRuy7GjmuPhgP1a5znEhytKHDdG4OaACou1oTS2qaB7HPqVSOHKTY44
NGbXVoIALvcGlz8O6DvtkRu7jZSdGgG/uZLWboiAK5Mji462/q6tc8BPG0/CIGehCehpqMwSwLm9
DEtlaRAA5Tm6y1zrDP3gL7gL9G/gYVfm9oESEEyV+tMYkMfHz7jhlbMuzv0UACSldddUzdPojIB/
zHh1LJrs5XCQ+A33bm4YiEIhJX/b247cPcpg47ngTY/nG9xF+rPg+9roaSA5TgMyAPjfjVAqeWUN
ihn7nquAykq5aT9oUu476DtmYovNFdIGvCu81jwQOw34u+zvUSdB1dMjujK2LScOjXKFO1c8JJ0+
1YJA33rEGaydBAB2yJgpRYPG54VY0FbM970qwII4QY8YGKOiNEPkcgCjBXWO4HRJj0V09PUxVCqj
BW9o1szZZBz9m0EiDHfLW2mLCXhtP01eELczOiskCHNWV/RKKp7GKJrS1cYpe682VCFE0/XGTd0n
CIGMvfa0FIo0iDBa9aVBRzu/VB4rrhHrD1w84QIFcrQIlb/SAZlo1huulEmMUp8G08qLdNagv4E1
+R5ng7T5OHbPf0CrTuYpKb0AnFiVUn/5jl7Mxjbyh/jV2FC0yavIR+SpvWI7sR3J5PamiGbSEqCn
3iJxM4aYBagW6ja5WGSLNCV6pIz6ISBTCFToMgNFqFn1BzgigHGL5y+RnWJGP0UcO7rPaxxpp7Np
vVy1KjT1VGT7QjR+RU1NVRR3e/8XISrvBQtZUy1jURmMfvkyIk32JAlLSfmKxlp286e4cnUInMuP
+e/0lYT/pJCdWbNlClYyaqH+H9FOb9fS1armcjKFxjDeBhCdcKYWZD8DVcSEH5fDzItS90ldSVRP
X12ye0zU/wrySBkaebnYdNstrDoIFGP8iy7/mgtYvPLZ6tSaXypFs3S+ghprOIEf4go+4IjfEwLV
YW2aPjalwLu/cfd3Z7e+rSkgb/ApUpYU4v5EVjfFxsa9G1XbnN7Ach/aGjil7bc0I27iIUJb6HIE
pYDTRDmuvRyw56FdnmTNFxX9rMTVW3ffmYegWxsDYnFF6Jz2vSmhsIZ7bKu7QJ5XpDsR6+ef0MjV
Z+QV+YsTo5j/fXbU0fCctjeCcdsHMwOICr/7+2aMYOGft4dOaY3qpr+NWj0h9Mpk1NpXlN1iiCFe
kpNoSSkeWfv+3DgStyG4Sm0hZL6OGk9WIES94JdTmyUeF7XyKIRJRJt2ee7jFuwHo8foi6pH9+0N
6AMRI4PF2mgjt+pWLTn2Jk9BqckfFzB8+uBaQVvkzSwqFnO1MhcmMEmxI3Uk/CVFaiiw7MvP//Vu
QNgLfoUnKkzARocRRRHQ+FFFr9HpZDKegRLAKGbK94xoAQrT0ehB7t2zEUeVrq2yJtTLEe+8C4dA
HQeFAeIpwiHp3shO8mUGMVEBLTBvqXI3Ki1uOZ2RpcgPFmTt09LFrB0UWrf0XHaxSQMC60j92EjN
GmSRUz87Kxnn09fjz3ixVzQuSnDoeVeQqNvZhctDvbkZfKi6m0Mi+4DxaFzUTMxeoy5okNO5suXb
/xXOvInlRl/QITNfvmyQUCgEp0clofSFhqoSndaFKf66FFuVH/c0WYnEyBul34wj8YKz2jFyyy5m
X1pco0vmmcB4xGduDKvb4LEWX2wPnp7cMi7ol3V2WjrUBnqa8LFCKjFgWQbNKSamAz/b2RpkYCZb
5X7dgjiHuZoIhPqr0ELy3O8a/Q5ikBpg3e8Oh9vLT1UPOVJcHKGSbODVQKf7tmr/aFUGZ2p7hybS
FWfY2yK0lMpgjJYzkOvt0bRl9uHmu7fcurkmqxbkRaYiRitjjjbG4XWv5aXGSk0saX3GOZhS0gtx
jpqlE8ELj0Bbr3GKrET/sAM4dsldLIZ+W1YLwIxy90/6ZdbmqkFGaM7C312yfRxK8zvPqY+tymIf
2ywKTWsz1W26QCVt0QbWV8CRfPSd0GDVBzopUSV5H4ssyeiumjruMVLcjiY9F9HfVDUxoLB5f6Ls
BZwbN1PBuaVUvjqe6Mc9T7KOQY3ZAPUpSz2LcY+T5YykWrR2wK9sfNITLS4dl4+MyUGR6pATFrF0
qBPdHCWaWK7quD2qayFsYJU17W1oYl5WTZdSGX6e+7nOkmEPfxFnkxBYigSJvQWpdYcVeIGAeUAb
rknP8Z6DmaFWTTb5f/4vE8PJ+hWq19tZLgTqnHuJlyQC/lYGOn3TNyKmofuIVmRc78nT37BmwNAl
mW+dl6lF9ad+oAJrIt3DKkKQ9382LHOKZ1UbdLHmMl63DOBNFK17qIbIjvUNyHc37EUs9dp3vcaE
GUul22vj9ZslIm4pX0u8kfIMqpRu4+JYC/bxTqsVv0T3kNAD6htA5aRfM//G+hDigd49qI0G953s
D1CFLcrW6AU6R3YUPinjKz7e7c4N5PQgr1ZAWTBXd1MeVIuDQ5vDGwVzRJaLTYep7gVekmt1iBf2
npCP3t0z84Tn6iPr8zd4FfW5ZxnZPpaAeP1d9unGNnO4M3pN0rg2W99XKtdkff8/U1jDhGm3Gi11
R6PMl8zzAxrxsrIM6yvEiOj6tiPy7ah9txUgabpyWKkmxYva/Zx6ICC19jd0W0mb6KxTRAwAISgA
tqJIg+Gk6d6Htr1okh7mMtRnjSr/91yfsBfNY/TosqPh4WxbxEK/yqunHYR1ca7P+8odNPOLH+SL
0UadM2SPK8eOL5XRcPcagjATtfvpBcCpntABS+sFbALN/yopC3luF1gdtT2SmgcDL4G5H3Oa+WKa
VQl0HJifHytKHClbnw6+p5eV65us4021kX/Vmd+tyYLTrYP+kFGjGXEpeW62gIZ+qtUR5gdoaqz9
Tj0cgd5IxTwupm66pV53a+oLMcr2NrD8xio8osKt4NaWEbP9RtHdKumICYhc81zcXFtx2jWPtzn6
9nw3YBnYn7KeFUHpywWuOApuUVzd0qbHF3vboIA8d06z8oNGO2m7NQTZQtxNX2GxkT6AFpZyTqH4
36V0QJ22lKs0w0S+yo4LC4FBJf1tU51jB4EXCtoG6w9MnkdzWg0gni8cMrJkJHzlJUOZ9C2lb3Hu
yWsnmvtAcAp8b3EfYm2mKKwilNWB3Qh9gBPy3J6Z/a6aYzVBE2YHwOqfVvnLZN0169IaslLFNgXD
Hedwek8IsoXGRsMJTilhbaAAOr6pkG+II6lyfAYm77KVQmt9TtrbAtadYd2vuPBnFGmH9gGO+pzf
NhCsWdKca038/UlO/21/PplGkTbcgMlmzo9JVievuBR4CjdDtKkUmjy8JwTNyX5dHSe4m59ZETCF
nnVWj1S5hGQskYBkH8ZlREzMq0fJwRAh1bIT+6oa4PrGRSmGQL48NI9KCUKS8aRLsa5qRjbBKFt1
fnQe0HT4wcu5f4CkNZPKLArZKxELcaFhT3C0zGtP2iytqjSvxyuzYqucmLl+2Do685mHmfZWGhNT
DzklWs5AsCotxlq69zYi+8gzUpVFpqlgaGXr8aGI9o/DqwUAqzPALZu30+eati0TEL63ch/GnbzI
T+lz9OU4c1igcJWrJLapO5/lh1TkQ7p9huIx6drn8Sfooh35XFQ1hzPcHUum+RP7BpmKRc6eSta+
WSYHThEt/8bZzRpjo4l7cMLkSAuzjpjOGQ+LAHBMi/AeJOeG6LsiVF7T9fyI9kteLZomUUeCbf1i
huP2rxmXpqtJddxOlJwUUVV2X7esxZu9Dg1JwBKpp8uIdg1+KJEK52cwEV0bB1seTI3bGbzMrF2T
k2n8esU+XeGnBA6kHj4OR5UxHa7Y+Ar2Q1Nzmti9cFHHTmTY7On5j9nD31zjzkzDAERBVLwNIP9X
5WLkjRMkq1WJGZsrNxEJEiiSGHg9bmeW0niJ/dJyufyIqavYi4NYrPQ8S6wUQlOuEtMNcioojn1c
3+ZVw4jv7iHB2lclGgo7lYNOXxKuwTv14I16IFEr4nv2xDhUCxTSx39n/oy1SnTx0g/uoHSqjE2h
rMGHvMN2nPXLcK6D0D/2adXTCsfl+jlBSSEi+3g0OIOF0urf8sinEaha2VeRiywJXVs4epaN7O3F
bh5TXR6tZWpjowOngOBr4nt9SJEsfrFoRS0PZdMi4RIbtlN7A/KPAwsToOBRADfYZ2OKvLbuT+F3
AlJlZ7xgyh7yuhID1g/vArvKEzWYo0fpQo6s0Atlgpt05FQUDePMiit4zPHCMLhl9FIyYgplvdM3
2XCIpgnmkZoVvI++VwMhJiMQCJ1LXWr6e7NAkrx8Vj9FhptlxXCHYkELwP0RZSATruTql8bpbtfQ
YAUXq1lpGxgYZvkC+U66HK+nvZwrQtXNDdWn34IFwREwiFNQdV7QST3gT4g9YrSQPiZx48KGwm2m
FYB34nSGjjQQesjurrlAPcWVlbvN73gdNnbI7fghMrHVX62/KcbEFIFZfIHLrj+gBObXtHzvEid7
SgWlUfeR5R6y4UvuPFEfv7eYHRigqgKhhR0RMIi/b+mYyAHwpVMUwdzhUKckIzEBdjxPggCipYGd
TWO6e6dWSED2XYZbr5175b+QZ5/rGkTVClUvl6L22QBrPKTR7oJl+4hnyD12xyEORN2ocyFfEfuZ
s8qddyl9z+g2RMLJ1Jg6JYY0WaG+qwuIUQWZNTMmqKael2+iULPdUfCsuUmFEoOaCwaD+gd2sBij
Godq/zdcC7nK4VdS+wc7vzVMfRPu2fsUNclYSz0bnV9wjQ6rRPk2SEOdWjwgjarbbpIx5Hakvyp6
yR+BzSmtOS+dbwx2oZR1O+gVEbU9ZBHzpiCCkuCVhheUE57LmHL1xIzLwRu780YotLTJJ7kNvUwV
osqtjw2q1gZgFvus3t5fj39BfzkIPQPKjbkGPW7P0AMgtEnEG8oXUhBZw951cosYJE7nBEYqmm2u
ztAmzOKQ3AIh3qIlvOexOOg0HNzWRzxILZgfVtHEcA4/vkMFg9rrRW/fmRdP6g7JVjSSQz7+cBPo
FbdOvYHMsF98fhRmc0zyEd0tI2C2o64SrB6Cf0nCIkT/bK+zS0gLLRTIZ5uV+hd76ll1RTnupgSa
lZmbOyK9ZYo3LXz6O70Iewq8jjqHlYlJiyitgUyJWVoQPVAlvzaIx3f2d7ZQYMNzw+wjdE2hZTzT
edJxuxGPPrEIo07sNmyufHVFQiCoav10kdsvrcfSAfGkk2dX4ZOSNeqCZCrzaN9BnoyikAa59hum
veBXiaEo7k7EslbX2nDrkQCWkLITrYd//wSyAa0eksZjaF3VsAuomZCEP6Lx3RiWYqlLaJ5+4er3
YBucxPJ/zgYtVXoq8y+0JwWW+AtDET2CTr0jTJH95/WBS/C34CQP92DXafTFQPfLHlKYN2FIRdKl
dg2r/OsXnMWnbqOS1Cc+WcIOl0K9dgA6AuzrwmGDv9insNut/DmHTOMhAOU6T1gPRmCHSJ+8w2Z6
ORFB/GSvGReDc4ivRjSGPSD9mouq06hWlGRrpGAUKxmWOMcPlDnWCctjjyix5xp2QqClUl8cR6LN
RPmHtcnrZqfETgajdMrV68oXe2DcIyqteOF5h4cscQwyhotG2ML9kOPpcxicjueI+8ockW2S90fI
DAExI9fWZYFJVMSgs3C+gU0FQQdW2qMxIM1az7lT2/UR1SOc6m44OxUUG6ZltaGCXYU5NJSfVla8
1fNHvqWeP01NqjlzKwZVCC9X2vs5mDbo87lC2VS+kuMa5fuX9L6qbGBxLWVxLhLa6SKtnswnrfwJ
qpuCm08MVlwyviGs1OzhTBiShn0yV8v3ItZde7UbORhyBlducSt/i44c3ai9ndVdcGKyANkHh1mp
z3m3bY2QXihsTwq9bojFOzTIXzJhTlaLGO6V3i8Wu7pBfaFB8u/HGqAm7MXmvZizNmuAaMssD0cx
l5P5SOxs2AkPkgJ6AKfPqU2pilUbKzDyAJCZHEpxQemdb21wesh3h63O/HDVMh9CwE1j6kcIyaZU
wRUzBpa1ODrZcTOer5ZZ0L5NFL5zfUMfkiGHBjIyNXTLMrjcbw7PCSSZUsZ/yLP0AYsDgvHI5KY3
F0Nrin2+LQ9+r9mK7pLxivsu3WX24kg+MH5QD3ikx3JfV36tPfKL77Yjt1aOeZl3QZ06jJwFkndT
6eQwE5V3CCY+ruLyarlH1pT5qRsluB2sy8JA503AiPXDPxlDXoVgSaGyr6CWfvhiEjEEIaxGxkFT
R10aWd4PNkFHh1fO970wFF1NIgwrUfV3eX9HEKp6bnzQJ8IWIoqm0/XV06IP59lRuQfZ/R/266Ib
FUb8GX2duPgQt7PAu1WEwD+kQL+1Vjb8S1N8t4sxPMjuVb58wujpLGJK5FXFGO4iZCqYut34VHuH
TFJ0K2c3iS6Mtazp+VtqUTungtHV0/61l8Yy8m8myKObvVspImTbzy0e+RKr2xQkSH798V3rtzln
RQfnXvVB/4hs8SLX+V5TgMfTP86NJZAXt6RW0zQax0Y6UFSkqGlD+dc0EBljJoT64XEFBX5y782f
ELIUYMMWxtJeN/GaLysiT1GQcYIbxStto7jHgFfZcJANMvelAT5EP4YV5L7gjfN+nwJiSdQo93c4
IwZ5pc68cKN+eSoVFbI5lR78jnjW9qmRC5g6NydBo16BHdGJKH212Mkrp4633wfr+Ov4AIzkEUna
gbICSaMXkgsuO62F4H44JIdflBdHYPKk+SghgJLzwwa9nD8l4ovS35BaPrGZz1II3FEQ/MUbH3rm
ZdygFYhYVonUdu+8pSFSSd45NFrJMMzFYFdr9ZpRgWTtKgKlWC3Bo+0kE2HdyFzlBAVL81aB3xbb
e20oS/f9PMygIDGCDdU+FzCn+lwEj3pNp+RK1whBZowk30sR2heFFdv6QIZXzSVz6xGgGUcSPNiE
kO6cDh4r8MrtPtFwAstgMIZV5F47xRDynXy+BwjkUWHRjon2Dmn75Upi9MXcxFHTjiC2ixGKkNxK
H+DBMSAVxDkw7nV4/VRj9npjVBm6Sn+TXqpi0UoF7cztQ5s2Upw/YoXeh273xkbNtNGpEWcWR87B
3tjK7l8PayyCThWMASjwmw4cEPvb/y+WcQP0C58oPOAuin6arNgQs7th1dy9TTwC34bt4C+9RNWP
plkaQbF1y3ELSbzVk5F61kFGGSic7diJwvkhYfhGVIA5vvDJyZ7U0nF9kymhHxwpyyhL1NeDH6IY
e0pl3q4nALLvdeb9fTdwJm1jxPNmrf7UcObRFNtU+Z4oKQi2lrqdkLWuiCfUJFXxDzGZK/3Ptc4r
kvvsq3eZeYZTQfjHEc2jkcB44K+6ucKBZTBkZgeoiNHmmgay6kgelZLpXK05CgQuHM/awdmMT5zV
aGf00dGQ1S+Wox7SkdXWGyoFJtCWJtl0Muh4eO/YBe8Jjr8Lu7Hp+AK+8utF4/0JJSdHO9wVBGnK
fLfxgTVSExr1DToHJGOubP0RT8OjsHbNl/TX6MRoeb2za7jvLdde8ZZUfVRMeUHr5JXxNA4qZYXG
GndgwWTGDUO0S47zkVqvC2O1u/dVuCYa5d7ZxnbGogxpz7ThX7NvlLZQdP+1uuBgDbXpsuqo34gf
kR0Vw+DbjbQ82aEBJqs1PwXMjC94XkNZyzOSl2oT0BMIHxsBTA1+yODS5BjhzuujXAxHkKRbQMxO
A8uo3XvgRFNuaGdvxOY2oadtOJyRXeUtpgnw9Q92VZsiQdk22fYJyqKLVauBjVA55ZXemZeJECuP
ZI5Y6QRXBJ7KXR4khB6rE5B+VvcllAKHpERYa9ZJf9zS23h3ejPoDu7ks8joh7fmc3DR5A+/JcKl
HTtMN4wENDAsz3L9qtboBecnj6g7kbr2XczZZQO3ohWauycRoUkbWeKnZDo6OorjVqApDDIBoaF4
2nF3RkVvtvUTN8ZaiRe2CWJLqkcxT15X56yi1agnh2ZWuo4DC1tnpB1TjfYc38yf4fyC6C6+HX17
O7fnFPTGOMDnssQcKenzwysv/KZderuPf5jsGKuvYBk7iCrAER9Zbndnl5r/1FQLA9Kjk8oXtwBl
/lQaeJ3yknppVALe+usd2Clhbaglb4039aWd/3rI/JmaJKJLK2MdiZKgmFzh4aok6K6AhnToX82t
U4TMOWgXopEgHFWhIhovENFT9FoVwpeVP/TPlKjFXjY6P709MuMoRqhG5xWPTU/JYal2wDVP/9q5
T5/ykIum88LmupK9xvVEhuoAv4bOdBt7711UFf3TYq97ztpxfiq0HVd9iIlQwK0LvroNI5qpfdKV
1M30KjPFUEmRmTr6+jAIWITFgXlUhEFGsB5maPI4ziVWdLgylyEkvuNJaSNqd8abWiungh7PetTO
AYixK3zEFf+TKyaC2xYk4LB7tkaGrHAcs9FnWZU9CNeNdI7AS1d8M99sPjwWBsgl//6JrDpsdMNQ
Cw0EQLXEhY7pvibjMJIEA7a1XgzRduIPuuxSRbsolCGiC3nRl0dAQcSkr8jvWT8ePsIka22gxhSM
Szktw8nXSQu/a9PSziS6D0LYSFsZqJEsXUfRnB9nuK74DmAdDa21jLUFZGWjXb6tfpqgPttjJaZU
5UgZxN34LkXN572zfSdVBcQPE78hqq8OWweg5V7dlaQKywMCGWYtmN9FnNuTLpXQ5E/j1ZWFELBx
iceDEx5Cql5djy6I7mYhrKp0NbBgE/odh8sKr7/TUgqp4zxfGUvjuPDAokXXaLFT1iehIs/XyK+x
7/OI+qRGj0wiUWPuZ/RL1fE5LP0vpzSqua3HXVKOpw1soMv61z7jD4mi7Q8/GO3YG4Ew1xORmmmK
9PcRY8fIbpZsTWiErRwI4MsZaqtpJC+4B5YGrO/2Tz0YgaWVY5g91Df160cNlC5ITlG0pjs/b2Rr
ygs5eu8JMxvLsNZDLcUUbC+tUmYBzXEe/74XgtBsrdiHIjbnWqQaIopw50yzmvgn/YTcfkgjRqP6
rhCRfwrflsKC/fIAaDkTIepz+kcJNeHRbQIyv+STvjCFDGKU8m4FlXADsQngiRwTpF886Hi7Y0Id
t335s/4g/VyaEPHSacl576r4SucBkg6KGFdS7P8TFzNubT7poao4fo68gy7wdaAV0idIojSlj7uX
T8Unrxhf1m9VTkHD+XLn0WgWuXjbls/Mep2VibI+EacYAeu56Jy12WloVbnz8gy8hP6o0d8aLlKw
+ItQ/Rb6YMePtgoINpaBHM+Y9XhtXF2xEE54/B5JTWcuTepzz34tsT/u0bT1YjPfAenv5/L/gLzc
gRpramkCE8UtcH+J7TDF0X68k4eYSsN/7IozbusBxZcqdu8/HArEdySRFabB65w5hN7Z4IfXTrxD
KIi8hoBcU8PZL6nWskC2O/PgEX6ArmMe+RVkrPVhzzTq2BGoz2T5Wa35oxgF6GkE/hz2gt5/zcty
VcQD7uD8QZ6YhbY2IQc9NEBUrCzql93I8Ul6lRGoymgCnB/rhEowj/BaS5RQtp2akceDGWpKmGIo
qg64hzFGl3JsiHlZBxlEx8aVToSqRu3grudb8iiR0RdTwMJDTKkH6uFkjmCxTUQJybyc4nbV/NYf
UPE6UUpVVvvBNQ360/uqvRCWODI5XSSmNrkCFhgEI7opLmNK3IaaYsQ5YQOeULThcCMGz0fdP7qQ
d8/AqvslM6G8qqPPC7snkUs94Ou4eEXNaCnovxxex/BbhhC8dx4RY+ABTJKD4p++y2Alfht5P0AB
UUzm8h/Gf853f9bM3aHJSLobvsLi+nlmOqLa0GDlEBuR6erGe5v1o8Ef5khAc3RA46uqYpKRZAro
ZuMAdHPdC6j+zZcU6wGvGOW/CuGpdt//4b7w+NhIb6a87qW3L0kA16jds2Kr6cTwc99qNQdzCy+J
+lmROxIonCbSBfLR9XC2M4J85L5KboYiopog9WyJ/eKKCo6ngOjrMPfx+uPso5KD8JTbfz5e6gIE
ZEBUY4+goL24h9Jz6mbbz4KvEs1wlfiOOF8SxPR10n+7pZMW1Igtf/VPdVSpr1W1sAaHMsejdKnM
l6J6YS7rJ5GHz9cS8I8jDqVOsRVaw39F+R0Qo0Lthm5rrUT5kHFs5WBZ+zGTa2fEWpsDALrg2sfO
X+s0K1B9yh3A8CDeyiqRRb2H4twQa3y+/DX115Y66co+PTnyl7Nko6lQ5L8Sjg1oNlb0o20GCUjx
dvgnWtb9EPMQxvXdGGoYDrAVLu0aiGr6V77io87XCBK6BimpZ5idXyMlnGU63QQLr9Gcb5EBd2/p
XWs+TVfx+S4CG4QesSxmFxft6AKq4V2eIkaS9pAWfrdBK7MuXfkGBWx1pl+GJGLUbEpW0ljMGpP7
YZwYlxa4AvXEIMVmLaJ42+OjbVncH5oP/LKR5e8mcqFCrZJ0ojJaw3ZS8MhC2hr4sFdoxDYE+bQJ
1mmgXq98DdgS7rLqZB9ddWk2kcINeOrLifjQCBQKGZ+w+Z4VRtOkmyEIxz08OIasIc5+qW5EkIt+
jr/LxuuiEhl0wTIGzRkcVxlmOYAAuJCuHQqTAz4NNdIfPLfMBNnf6fAWVnouTwjRlqx4xKNoI8rt
WFvdyGSTCWh1t+xI3LpYjYqRS5N9im7rtxHnQwhq2x6nCyfNX1wF9VPXowogHFWIse95xPwP0oPl
0oL6J4nV7CF1wKUBEWSGba00KsI0x5TWsAYb5AvEQF+OxVXabgrexnDKl0fqm3KRq6vjg0LZ7CiF
ay53RbeGu/jiRM5L/Hp08EDIB4R2SXTBn72ODc3rxFklqz8CLewfT2EjqJY4F0lLDO9poag5JcUJ
Kz3St++4gqju8CW2rtlXo7HgRkEmSUEcSHdXHstC1sIeycIqnv4QbyhVZd7itvH9O5tJZ6jIkECt
F8XiZGSRwIf1fC7BhBsmIz+TQuHUB2B59xfuFwboS5xRu8qIlWzmCtNvb7IH6Z++rIoJZk/atq7P
ecYs/OR5JzFe4i07RIXI/0hOudfPOgGrNW9FYnbdwFV98DyH2BYNGCYUVO3SEwrzYHWxHhz5cQ4D
0hq/I9AAh5azrR0EHONsIWDJLig2T09NJPyN9Ri6/u6hVRuSm2P1IaD4GW4Zjv6SYkH+93mvNrGR
BidSEbcTwTwzIHpne9N5UMxokr1Sdt/dCGyb0ZELX2RvNLdzWwu0aSW7pCGbfuJ2XwYihQi8RVn9
ESsJ43AeVpYjhvlCi5wywDbMw5Ja6FSV0A0bqU2/3oToRgPTiyZWOXWk6Wd81SdVeN3zbfcUcxq9
dMT0OcJVsDZCmIn8dMM751dYqnKcfDT/JhsAql3QQPDYTN/Va8lDJXzYHh2tCH3RT71iP8PK6QxT
Sd7iwWpUBwADdeO8BASaRXjBvPBArgecW05+v0MquVJICCfZDGYjQ3Vky+/n1B/IF8oPkl6RagQP
nYm5QtS7S0aa1jFxZ5HD5/2kiIAESYuNhbL+Og/uCMpp01bgwvGz94pomtAXFMk9BkpwMC06cmJ3
qRn+ADOJ+iyORq98ML5D6BlUxYKsNtUut1LEyLd7E68CtGxlbESQSutHGiyu88cUi6m0yuL8v7ho
EmvfVKHBaejd1bLZku/5rhui+iH5TiynEIOyM+Eohiy3mEyJWczeXP1622Gw/83KMTGfv0FEF6gD
DtT3cbqBXsnAE/cJ2cakeFxR+/m9ETCpSAx56WHgaFlVT/ZS4EIDJXfM7bh+3NGM4l2S9kK2JsEm
NXhhRzwpvylieT93qv3ao+srdoK3T63EfopkLyDyU0X4UfOOyrhsxY9PgXjlOFdB6oww5xKkmxjk
Y6/c+fT87tQjpHBGH4k/hee4nTNaBg20++KQLUq0DNeKQC6OIiQh4+ARPId87x8QoejXVb1bRp4e
SOaeRR1ZP+ONcfRXAS8So//e1ohnUHv5EO+r/uqkTEwLVavBQvCL4NY0cpTIAgRBr3UvV5Dozqce
l65xc7C/EYenUpnqwt/rUkKQxj0sbdOvFckdcZYU5ieh4GZgbo8O8/+++xPA7KF2gaTAf47yQvIz
LyRPd36rJQOSwN7OeTzNO82Jr0fCk8X/s8sCHk46z4CwMFO58H5q7dBwGPjKoKw7o1PNKXlU6iGn
9ERJDtrvHYpbRK3IddXeH5qZ1jrsbu0s9uZj6OQB5oopdyukmwPuRCKsx3spzDus0QspedD3PdL5
kfKWO1EBFNDX9Cr8u4LQV19qmjpmJ2Nd74bNv+FaI85wT5yD3hp+ZkAyWWrAXJc/15422wnkn6tM
GXOUdCr3+of++ZqJXO9jhjgVKd91q5s9+0o0b+TDIYTbuckjhl10MuJv0jhUSmOEsN86zZOsX6WF
Mm+dap5ESVKOLRnX+G/+fJtpqu+ZUJLQN0GERAxFguiYQ4Qk8RdlL1TTcfhhzIzREsKKUCRr7jff
ZmIj2Rtkq2AEQT8DcBuuyizMg20hWUgW/1mCrbRsZFbw0a4ikjfTtPYyrQHGoG+qtR8Noqrg5C3h
7awzppLDH9jL1PyW6dgjF/CDp70w7o6zyxJwcjAl+IL4T1619uQz29DmRJ/oQSEApa4qrO0oaqjs
4n4SxRYnIMrI+1RpffTYb2DEQ5eavFYEHiIwGMfii66lddy6zQUbaPQ0u/HW8HDi4zK0XKeNLz5z
lQGdK4vMZmjh1czTnsQ9zi4pEBsDTv12aa7igLywiuMBOAzUHUHhYpMEX12f30OCSgLVBwq0wdc4
a5ynGdDN3G11V/52VMEeJhwFj1O+YcXUoyfpm+zGAFg2k8NrBJOm+us+u55UQlg/MWutYZHc7Ig+
PLbm7bjubc/cxb+x5IcuYROlLnSk69eY6cB7vIioF432B9r6i5wqlgl1rzCnBfmynrIkaFzMUHK+
5VTdR5qwW+BBYkEPTFx5wTWnwdRimD95Q113ozIM64Q4MamAtLMIAAnHcoNI+isgk36tAls6nZT2
VdWn9TnFq7uWtMVJQoJmi00wVAleGqggp7vEkhzlq2qJJT8O9oyAMW4UdzRUZyDnLy41oV1qLhls
aXse4BVhkzcUyfn+X69PweQ/dq1jzmJL4/IxDWTxvg1utUTDHq0bs3QqbikU4tdwFqciNviuFlB/
aiAjX6PMQcQ6LiRlxcFqIcpkGFDxzPNjez0BrK8M7BF/PxLGj7/l7KY/LLaJ8N0uVqvR/hJWjWwQ
Aum6BB2njYyyE0uCQ8AGfj67rFPR2dZZHP5Ue5aQEbYKqqJhqTeA12yFcBHvFRuiPevwqAmfSgaJ
5Uqk+Y6QdkM8n1KIrn4nQMJnvt+Zo/WMf6lfbo7bTVkyf6IMIvV4qbiobLpjwtqOzmd/0Vumazel
js7NmARin2tvbioXG3XOkMacFJE+7TyKoCNiBc00hJJmJa/OgqaG9QZfa8ENr1jkejui/iQfucmS
8CqyFeeoddtyxJF74oCNWtwXmt+dXe0EmxmX7De6Uyn+U2dztdC7kCysHM9OeuGaEYnrD7Z91U7Q
Ha5zwXUA+LPOQYU53qOBouJDB7yW99l9sDkjZ48okjuOG+RSSvy6PBj4jg7bqbQLsVkeQZuG516+
WsuK5ILF5DUBKpzsYCvkFsLCTW7Ws0jc1zghde5SbqOU4prKYjx/veswf2WgZozLNnRMtsWzpL3f
xvOqHZAa+Y/ZxEya196FwWRtd2vnd0Zps5BQmaZWDApWayTi+nanYBuX4BOErybYnepTrxSzxk2r
Adbr00UgvvYvk2Jl3D4pLk7nEoAfa5FO+dz2JUuFUsVkD8m0lJgz7K4FaRs0GHTA4OXeXYMy09dq
xlwJ1QnTpAufOA0S2ywfco6cFauO3LpLII0m7bQppgjCQJNd0O1mIdSx7Wxnc4pgAxiHGdPjbyjB
xkPqmFvjZ93HRTa08Bzebs+tY9dskn6bWVzMZcETy3Z8xA+SbB7wUO1f92j3/oIKHXoUoVVMWr1l
olcZOTZSE/qfYPuc8rOwmxZEZj3fMK7KpeMyNvUPVKb3SUIJvuFDioAkGPlI7B/gDY+BjoSqt46G
pfyosYDS9y31O1AjWDuKn4dIP2qlhNgaaw7Vw3m47yu7LMflZo0vzg+/CKAiQgLWFac2jtrjBQ6T
5SBAgfWzf45PB3HExiXlPLmkPMX1zqyLWRUILN11HU6Rjmr5LT9E8nJA7T4QePZbv6jYmSPDoyc4
8DQ5cRWX6VYC38l9sRYC98kMZ/NFCM5wE5d10iTmuBk/Hp48EtdPgnE3dL1LtWeeQi97a1NbomG+
3grQRZBs8JdCR03UptV6UMg9zbSUf+CSkNENvErqNSh7uOaN8APktcEI8wbmkzPyCcWiQNUlhoym
QproNPPHWYPUrO6QdsQaaB139BzYf4DQBM+Y0FgVDzpgOwkVtZUBkNoG14HT6jaaMe66KI43ioLH
cp2pPInJfzLlN+hflig6Yb4QvKe15obzHi73Ju8+z68ltH/X8qvVDq6ofSQxOEbAblEe/gO9Jnp3
eGqJF+z6IDLMGWIZCL+ZanatcZZtxV6NsZNLlY5BlEwso08f9a7gpk4fGEJbOMVO9emEJcpBLKdQ
j5j5FiTOPbwKiXNt3tHkaOTUnAfW6NxMV8CfdYXwVjDB0y2J2TS57fKABDfxWSIx2D+fVeoPu8aw
aB07/SYIzvYMHFqrpIXhAupsYCUdrpjfmnryb6BJghCawyqXp+ctyZRouEHKtOZNpbnb7SsGb4Wt
OiIuI3iHf6JPvuH7Lyz/DURISKGF61R9Zlco+tEvAW61ab8y9munmFnMB2kVtIYh4cz7oz+Q3pgA
3sMnxYx2aKeCM0KLJfTympRoax3hUxASHVKBhbobHMSojACvLns+5lOXgmi5b9HlgLrm7T87WoJe
91z86tuttGtALO8fKB/gV4qk1My6xe5ONiX+kI0l1rqt+hl31PN0rs9FEvVAaJt73eVSU37gdqPC
1Yhm52Qii6dlT149L0KaRdSMmHe25SyYwLEPas9KMQUt97GgNQDFM6SS4+LkzgLrZRJqAdqUF0Ty
YrzN48+plRFltwInE3HDGZOjTt3tmpDk4uBqP4NY0pdZXxLssnSVXdoE8jAZ17ey/pZM2M66FcCO
x27Nq/bM08Arw/sebk9ySATzOyeQXltQmrSRq14xWJiT02D+Vee9nbXfbSm7L2wB5+9votdRl8Qt
rVu9vpKQ6F6L4NKGp2l4W0m0oe+ljMs3Rwt4HQqSqc2P7s3J7gtrU5L+8JAL1teMAMw3a0uFFFhJ
bKUJLcmHeSSxM5byJBWMOxnjN050jminpfJpEkc03zq/M8buAhqnaxrPS+QroUiSOYjixe6AC9LV
q2LmbVVsgLE22tT4ZYJ6ZGThB6b7sY+lljv20oOMLpeONdLKgHBHG2iA+L6yn2c5nvx4pihkrLQd
s/c3WMAA2OwvOSA9Wj909Q039Z2TwWRIZdHn/2k1v6Au5xdwKWB21KjeJJ1np/z9pd8Zlph1j/r5
6HVcblyHKxUQ148RkL3hgBxWVw6Ql5pimyEIYi9YYlIMeqRsp7vyKKhMbVbynx6wI/QaVZpvKOvG
+0lngvdvH9WcsTsM/TKDnIvXY2V3OnndawvCameLP2TiJUfleDuaUK9IlZJZ27GaSYWO1PU6u3am
kQ5nnCJdKi/qrghkKpCbXVeYlsl5SGDGqk6fL3OpcUAqO7oWl2TqTp5pmZKm5hmV3YYuO+LR5SjP
gKhDs+wngDMCt8loZNp0izDQe92I7FQV2dkHfPQWLTqX8DIFHCBCATBTLGjIEr4y3gphJs1AHBW1
shlAlIm4rJyuvYOFi92mQoX0yUShJ6MYqcIjaDLSjwnpwVnZU2DhfloWSi+QvDZWbNWNWoiwuapi
rkym29Hguc6pV60H8V/7F714fJlNThqil6nQGWCAQmbbJYbkCS0RrLoXIGb/QY8b4lCcANVskGDN
hcKDZXsn4Ppr5a7Jd0Tm6zIw0lqR/up8U06opz5kppuJ/uNLiBlA5V9LIxBt9iPfUfIBmY3lqCsv
qPM4zDKPOMeJxRig+f3dWgoeBfNYIgSXhH8InnM4AcdBoop0/99ELJppqta7DdV9qS5m9DTaaE9L
vt9D8aC3FXAnhb09F8EpyKB6NGH1MnU12dMCVU9+7yc/JRU3guIRfhSIZdEgiw5Wjlctf67QO97D
tTrhmErXa076/fErO0c+bQnLKAmCfD8U8N1J4QtqvmGqDL9waDOkOR2iaX+aavGh6mvAWVxBJbl3
dYmzccCsfDX5yo2E4kYnV3QZF6cZxxdDQ+sAs9SIAjhj6vx/miEQRZHo6E8LNljA2oNSf4ZPEGUB
CIIStadx3ayqC7/DvG/7ChAi7N5S39/9XQeRgiL2M1rKDIQ/N47QKfAanw2IOoir6+Lx690MuxQY
9/3dN79nPe8aLukKMBvA6FYkwFu0UozcXFmg0w8b7XPZMNdOEkVFT4Js9Ez/pYfGaMiy+ljpVACv
DmnIPDO+G8Xh8RKEb3LtU6uF51j7VBHHtVBnvjH+L5fuGGH8X+UH41/TUjSR946SB4Yl+0sAtBwt
u2rURnuGHPyTZ86m8VWJJtXku4ZFO+ADQ32novZXpe4DFGyYTtyKN3kFPrqTNGMj9MUyenCj23ww
hn8Of01npKeYy8slnJ2uasYnFsbbbA82Y3UU172V2tz6K2BHk6SHuEJ2KF9axwIChtzVK6tNU3M/
irt7iefwA+e7sNq1h/7UnxP3w02Byq81ANd1cEA6zjitiQ4zrWEblQ4qrcX211G3wblG5Nz91g82
s1eFtJkbTZnr54UwQ/oLkmy7HzQeTBuvc6c7IlgLprF2c+12pbJWmWkURzkWeStWnVOemPs1S2/E
RfCPTrV+UJjBCq76jyKKdccLO4AzBKPRevbEPiDwJoXEb6qBlCvM/nCFsDxFEK3wBSZIGGydrGZm
j2TSVJaioy/4uf78Lyp84Uw8YZp3eEjYVgw+uhHYjG3pizNKh4oTahDmOL3J5mzqrmASxDZ3v5he
mslDUxP2gjaUCMcftabdeYxp1188IMCRxQZIsfwqtnpxHUAJR32J4Kfj0VlfybNtOEZWLWfN6vfC
FImMpZGsLeMUVESoDH5PbXeqECRo62XgvA/wt9/VrxlK95zn48vmYmYEcz8oChHa4Pc+LtZEvJgy
RR8T2LBx9sWC7d/ZGq+LMfted9Q4DkQ+pRye4Y8PiL0/+jeNKVKXA2wAo9fSpv6seNU/a6UXeGqH
a5MIAqMbVUg1a3ibv7p3lN4wgxOqsYAtjQk31IUFW7Ps3V1eQIP5UxYofL1zskoDACfvcXP4ucJe
y8eU10AL8AuH83+TZ2UXPsml6OdtgrY0LC0O29hzwTZyQPF42QDnoNiY8xp1J80DI8VKD7CoU1ZZ
+aUObAIQ17gBiJKHdA53VWMO2fE8/ELBKDPsouQrvBfw3ZzqpGDhKFGgCD8tJiOv5O8EeM0fU6Bc
fnuagJF74Y0+MRWoniQDkEMRLojaWuvvMXXKsPBOT2PREMRSxpGCxsz0gGgOE05tEgTf2ilMpEta
4tqYYMqNX5ze3pAI3Ncoi45hIM9niiYyzt2KRMdXRthppL7jPUKKcVeeERswff53esn5WFBV/3dd
9FkHOwZq6cxO5AtDRTfgDM393cAHimokYfYJi5exD6D102DMZfXkXXgrRmjxN10xS57iKQpTwmrm
2tpnAwZxyt8/skLoj4EilCUDIUd+OWt9L5Ms2b2+W5Gud4dzdL/SZJej7hYOzKC5OvcFRwwib8F+
RrWQI9pV92j3XFdsNfjJ/Amfajc3uia5bkjPTwXgSt+wB4J0opAILhaK0xZPwmoMmjDiXbbdsR5F
P8/YUIQCF/hJt49DJVmFWU3ORe04OPH1S7C/sbReFg6eFCbhJSk5cACQvGqxsQkp2ljR9vrgJ0Mu
btdSeH+rE2LG+c9M1t5RtG8v8fIkWUYJIrlZgOCFsjYb5VEsU0X+E+/YWEPgnTNaPgNXoLk09Nuy
BwJySWoqeApYA+YbnI5DUHdWmWJCW80gv6OzDY2a7nZorSuc0GnlpTi9rO1bHXXnXR8qyH/sNUY0
Zx41k2Fd/HzLKz3qrL/64Or0lbjrh78+jc13RrXvVkVauSTl8qd0mrfB+c4elDWSrnx/9CKJTHaE
pQU0QCvMPQMq/raveU5yBKE7khXvaICOiziux8l/4NjGnm9DtglIfXJSG+7V05A3OU1X7kRPOIhI
euHd0Pb9gChpLlQLY9OFOFu+Yrfx9wS/65cn0Va08k77bDWHJDLRaLD06KbeXA0ZpAx3TSWC6PNk
Zl8kWRjVKCNRsADrcJdQHtlaAIEY7SKWn0E9PvuFQ6dYwM9/FgdbguC+1lsk3NtCruliTGsSjhyk
sd+r2/VEAdgd/KFelLWpu0naypCNscd8jZd2YROBBccobXzBuWDK76PKmhXVHvY/jLC1p8ir30Zw
3qfdWKAiMS7hZlUZ7ULWF73Ww3LMMQmn/2J6+yzJYmk3YkBwAxj8/ffUHMAdAupUSq6hqnRsNgRf
NPW+7b/ka9mJFZ3d4bopIl7+JDjAaFNwxeWbJB4hsntLgKkNChCIsNXJlmKRSOOISVKSuUk2sz5i
cPbjRx1TVYzh0ioRHAphT1PXCFBVbrtoCMASdN1Sj+5bCiykPumjlfnpIQ0yjBzc7h0LalBw4ZOC
Akhnd6hBA/eEnNiGZqN9HS6901Giq5LBaUOuImuo2FIJpQn4PPdYB1iIXhOcfvWQu6nz029FIX5w
lzvltdtHZo0y/T8OJz5mxFvRPy+s4OA4yFGxsISPKcM8fUHPFgg+8Iy+WtDr+8+reTBNdmM39lH9
ySw9kvYq+V55KYidWWKTwo7yOWsYETRsbKULMAz8H3lPqe4H9wNh/o78B2k9Px/J502Jdx5BwD0O
0/s+QPuh25yPEaYC/kK2BZQwVwbpraZPKUiSqtOO1iDYficNW4TrcEOXqHsv7zAE+QXgCwWyjODy
UH4cNF4dGDY35TqaJsDk+/LpzB/LTPE4dE414TZKfPbPmtkC+gzkVBYwm7yW6Q8wzyHa2gmH3AKn
Lp5hQZ+0cMMqM9Sq6hvUn2PyrcSZiEB/83rA9YmiNYghmn33u6DyFptcpHC4bhMmHOL0SFXEEQKY
1iy8/H27koP1jq0TEPlftnYmexquFPiFL4yg0bHS0K9/0BWE0rl0giksHEyzKDEANASH76itsrhn
w4ERMgHkQWn+2srIx9PmHAUNn105/eLj8lamOEeGmsID1aZ8tXHJojEb1htnwmzKUbHt4i1vF3EP
gTlCAqeZPO64Akea8xp9bQH/GSeRYlLTSb/ZqX2q8h8nAstmFbgKnjV8E9YIyXRlSJ8tbBy9tFcH
6Cw/bXa2HGXOGtet9blFu4gLoOEXMD+4gv7AhGzFwJNVuH+Id0Ci9gQIqi0I91mO0ksWVhWpyVzM
b6yMCZJn5r07+nU/335I7EhY6M99eb4GZcI3lxdXrxmUzaSeE0yGkJuDeQXqvE8tTsw4pLuzii9W
J2xiDaEoc8qYdrCuZhbFkACjTKBgUz7+dsJArVi6otaeLtn1vsm7AiWfS5KJh0xFHn5cvx61He6V
5tLmE2R1/6ZzfR78S3RzcBkhd2jU5s+Q1LA0xf/zxf0NgOex/Cwq/SnqKfYU/Cj6ZAcpXs/Ixnjr
AS+MoegHro3tIrnCHH89cKYGvTVr51EHWAGlvnta9GHsl6WCWwFx0YupvKR5vflRF/kFt0PS7Ld2
LomhyAwp6ZsqibgFjENXsOZg2ezCyK2LcrHAl0gkXp2fV6a1eVD9WNa5kX7lTRc32VJv9evbVaX5
aWOiPLPg3VlbtoWEOSKB63aPuT/8yM5MnZm2AXfsB4x34Lm+CLi2m/TIV9GDUm0GbKbq6w+oCQhc
TjkYuWknChEh5J8mHHoiHjF1Kg4bCkZGqc5Nolm3mRg6e89Mmwmh31zrG7NxAEVGzrON56616t6z
ckXVxvUo0bggDCLBfmS3BRCHGSb1uef4d2H/N2Y/d0Z63RBdCF8uVaBDdnUeba5aI0sQWxcs/Zw9
LafGar+1sbmQNN2Rv7ooFOIuD/1gsNMOKx+luh6ZfFfc4x/GFxbH9Wrzecr933qEJHN+8g3rZyvJ
fPvc1qtRmXOB1MgW/0u5uxlzOSpNyhyvsjRNRyaKz9Mo8w+Nr6nDNUlubnBZJpPPQHhJNCVFDzWz
wCw4Bi3NTqLKhi3qWZcn4IswY+JnNJzm616Vpiu0kGqVoOhQUF9aXUDlvUCCsWOcbMZJI+d5ufMu
+uIbsC13h7plp41lEfUO2ISeOQE+V37osVheU2iI8x58SHo9inoQC4Z8jUcslp5kvownGZe9N4ky
26WLBPLypv4RD2rF4+3hjeWxZLoDMMUdMlXJgz4DeLasOyHRMepAnW5B5HpesU27k8+Vhozfl+8Z
EkISnsCS2c8aFHpqOfcBV06y2sTPNJRvtS3uMpVyWbEpBzFIPw3g/0DbKLXsKb1jwMH31v89dnoC
peTc3JeD/QKeVc/tctUvvwrD7F1abYH8q/xf7iEXq2tdoPRp0fIl+jhogxTrxnJqT1TWsOYKepnb
U0/sB3q0vfseSnak0JJEpBIqyphBArSrVmYjHDx2Me2l4bwjAOHadKToLroNJXZT/eLS+EJ4pLG3
uO9nQplU2snI3Pk3cI6l+qPGxKwI0hMRFphLYPiu/Ai7ESNWC86cDjiFbS+rKaoEQbOy+9IyrXmi
KnwHUwDSNOiVHHu2mcv5r4lQjeGubSYgXU6CxgWjkyD1mFgUdc3YZujN6iV7TPIjhSn3HRYLFb+9
hZ0s0QJlUh5DMA+bELy0gL0FYcJ/NEasng/GhRVUhY5ZAHpq+xheNHGLkXPkTxkWFgeHg9Jbm5U3
xAuPJ09ZaUjC56z50d/KGbljXidyF2ZQg3jeCRnfar14WUZpsED/lH8gHyTHlqtXl2t61Ef2zHjP
feVTClYfjzVKCPe+xAwtkqJ2VAhdi7/lEtKp6MWr2irc6195DkJwvwpcyYC8GB7DykvaPxwI//5I
OGzRDhwG1j2qPBr2ok8Xoc3ooiteDDu+WGBorjAccFRkgeOph36y5sWQ7MQSmXWapAU2GQYfID+u
f1NwE5axzh3D/sOctAAAOqQQH5KcxKTu/3F8PIL0AKg36GaWv1Kjr5rxi3mVMi8GGjBX6DQfvydW
lT2T4jgRn2d2A71+2LvQKXBPDm4b5Yk7sgUQAzL1erClH6MjabBBLoDZbBmErORHKbfY44Kuv8cl
fQcpfoLiPXiVB+6lvFODD6BKDWDvUyUD3mu7nXQXMieWaa7YUTM95YElIPxlf+1SbaDeFs9SuR85
8T716tEnNQ6IICoczerAFeJ40oTs14rcn2D0k5xMMzycFqvcp1LuV9zQu87WjI4oZvhu6XuQKDWc
SAwX6SKAlmhj+JPXUAdL3Waq624Np9PdDJB2Uz0wnXn86HWEm21raF6eqX4/SISyKlDP8udct38S
DuzYVlV5BSN3q8yTXzyUB6mSm9okKiygBUcxjOYAXgGk/9BphqoI1/Xs16RY6WFpc06aSrwXorxU
WPnWSbB+Pwc91Jsx5NgkqtnjTy0aerQMDwIO/LCy+8N8Z/Gm0mdUYwyolyPhGLZ031kwNlFvqbrE
t2QDt3aCjeo7KPo1ubqx2NkNT8JeN6RlESw0cDeavmbAa8/wTv4/wECUyH3GD8OlDigB5DhYThnR
YRKdtYkcHIgJPWg0r/TksbOdZIZACEhjTGzqF5mC2b94IwSuFT9S0jLqgvBpvb4Ti0o2W5pQpFiW
OBQ+kddgzqPSHUqk6g1OKHEl+aQEGwUiZAvsYZ5u8fR0XNcpK0ZwjwGLUJ1GvUwsjCyP/dWTw9cZ
XCGjmuT+exq54vbejvlHsRz6ph5TnNcHSexnhu03lRpuDbilin341A7Z9s25nWytYRIxInyTLYvy
m63yQ0opzHcCQUq/ugJgUS1ki+dnL6nuzKK3/4vVv8zzvfcUQevZTTYJuCdOCUt5z5i5GuW+ookg
8cH/yQkmu5vG7ZwRxSyTj9lhXEl2RKpqIgSLWyas25pJMP+iCpTCNuBF0MP0BPZFnYomhkDOjLsM
o4kGU8PjP8/z6nfha68uvuNpNZa1wE1ZUVT2Rhjdf0BjV+Q3YxHWbXrF17pteopRSU6ZiO/6HRk8
qDQ01pIVBFpEwoV1BmqWbrUmulejuRlbLxyts2KFbCeq2MA0A09+xsfYdqbQJ1j9DZBfaW/ea8DE
sQkTXqzEXO0Nx75zGhbq4hEjrNyA5O1bmNm3w6qiZ5jEd5SGlMSQdTMBJyda2VGmhHTObQlICodw
6n3eOpAns6ljsQNR24aA2s0WPt1wN15yURAPO2x0cUe0552CvUznivFnCxWpc+8nBkV4DzlT42Ih
E5TiQkZUctAUUbIGV04EBAxnKh+0Srxl9bTdkGXSv52RMuoRu7esHVfGh0QMzO9i4VX/FwM/x21L
kdSTF5sl6XvAOzdxJrQHpfR5yheU2djOqF3qQFjByh9fIr9X6kdWu+ZD7FuPM6Kbg0hb8+DHSKfE
gIKimotveEO5v3Yk7bHaCmpv9gV6AlMfiBeK55SV4MMsS2Ct2wZi78I2reuoUPbGcYo581DxdRbK
fP+DDQ1qcr67msKMXO22zz81gSc7Tlv1bbxJEaiwml/2jgv+9kg3/+mxr0tU+S7zYhKaDFH6a4ui
nvjuIcRS1lztESKuBHdzsJY0kM5NW4PVPRQUyp4/BCpZ/N/n54epFKS5T5K8CAvf3Ap+O9F3I5gj
h4T/GdLO7btwstaOjh75yZg1dBoCtUUi6gMNcgG+ccaJL9tODI0pWmXeUela8mPf3E69a2F1xhQ9
mjaY4oJubWnWNys7o+Wsvpsg7AR5qE9LurrTIJLhcTQ9N3JbQrO1+j5zrDwdedaDb5Dz6wiog1Em
MtiD+wodR8vjyHWQRdbLGrQgn/axqRhKLwWOnO3aNEOlJvUCGvPmhyPUJXydrO3Z4JMKPW07v/7q
xY3GESbFKk1gQee9h80+FWa5fp1/xYrH+imFP8yRNOy8TrDVOa+PL7JSK2WKsCXiMvergLodJ6Pq
ML6QAUzH9bGSDdZEOjnm8IbRih1vlRxn/rokDxTPkrCMlZv2EjwH/D889DjrYAUzCWN9u1X+pC7c
ZcOiAfdH/MCvdNmXDvaM+QlFGoosiETWEDKiy6qEKtwmmHRSoiivUSAW9kh6VgkjLtTwiqhc+aD9
8lL69gts+OsZMgF9Mb2kEzr3/q9aY0X/I6vGMdxVVkl4Okb+hhKIP1nKDlnVKAH2KOzv1aos6OP3
USeYf8+htcjTrHuILSip1G/Jh+9NuZyTeSCHyoDT9U040iKbB8nEjk2DCvXtyZyrH5Rtww80yKlC
dOmBJBc0OfTWYN7fXEPUtzfPISxBCPQvh6LjX8tBT011V8UdsXaFoAi3nJZeTngUZHMLqV+htUy5
C2/KXgZgSPElU295VbufKpmfjjM3xNCrmlJALPN7nEixchT1DBDds7SPL0ZPDPrct7a7wi/nqsMN
XAfk4EwX2r8O36dIUg42MdijJ3tfjEW/2jnvxqTWaxmYkI10AAajOWg7nRoM/pnaWo6hSBdc2Apq
Wy1GO+x4PEZy3VujJsXgy2JQaYsaToz3kHXjR6cwhvOfDCA+uU9XGl8v9jsij+KQYaMTjnXhEIks
+coippudZVuS6TzFrOD5e4q+2d3fX0bJREzp+y17WrAIPh1KFku/sGdPyc3mOLhIpLA0vmGC1OoZ
INvu1oFe5JMOprpu7ZBo5juYvm07DUl+qoGXcu6V3PypzEUgsmqgRl+WnHleSGacrUIcffnWfqnS
JWFKfZ0UGqkzkO9HTB7l+3HXW9LfrsMAwm2kgcpFyWnD4u+i2VAy/L7QiNK7/TeeNzHKI0S8/HHh
DIEl0P1L2UFN3f2sQlTdXLHaNuSO+ASj+DUrxWvXebREtO4/zhlzx838BjIO7uyI0dMYLBrQP/Nl
ua6NX+/7oY/ldpU3AMNvmb2+6ulIz/l3qjrMQmXLQCnSQt0p2AvCuaBJ2j0RXkpUgAHHOIcvFwKQ
lK+eC0aTQ+PAiKUbvOoJXeWSdKpOFSY971RTv0zw/ZXdXBTLp2LXU85ovoj7QIUfGo6v9aFtPVsn
Q4gUdsZ6HDFA4Vjxvgx9KgAXkHEwiIzk+KvHmvFgCDJkbKY+s7+cQN3t4gSQAt6QjHDH5jQnggIG
5Dcx2+4LiFi9sdWYT6IJU5rJqSDzRov5zDEA/vgAXEZXHKRFiy/ghMf1a0r3dOLUm/59sTDihjJ7
Y7QizheDh+xCb//YhCgM0xd73RoiUtusyxCLvo9M41fuxkmBdPYC/9MyY37mdEnZ9KKPBWuiBZ3x
5WmQlxzTC9dDhhDYuplFUyMm4NtD3CqHbybn+12zMVQ3RfKmMCCzNYiFEceauWrcNk+pmnlyl1Az
xaD879zz6aKDxemBjbIBy8sP+xk5qIxwuo2wMOX3YfRZ/4jM877HxHQhvZ/M3/zNUPvm3Va2PBPc
CjMZt2sJI8x7j52TlvnoLp+r0szklCIOPvlsFgXbcCriTomBJNsqVxJ7iKpE2veGEnjlAQZzeCps
mv1X4wq3DYku7ZAyLQAy2G4Eu7vt4ELUldqAjSNCklEMRGu2h2Yw+8/MCc2KEAtBeNW78Rw9pr1s
xGaMUSli+5jfpavbrHuDPVNFH495IzcMIN2m/F+SM/DyX/n546RQRcN7JMOUTJkz/ySm9PhVGk7t
bAsx0t03N//MPV2pIWBaSQlgLPERAi/Zvoq68l02dw2Dan2jO5Pib4ze9N1W/ZOTghOe0asuSsTh
fdubEWw2dsSrxFeTVkgpIT92M7tK4VvUDHELqwUP1njUNsci8AzUKl/ilkbl3mYGdzwzIDdU7Ho/
AaEhSc4jGgtaIJpeiMvQcHgpLey7CBgoOg5SWzDhiEMmkxr1SDWML2noPTZEPJUZzilqaotRcHRq
VxXlRMVanhRPW8AlEa4nprgyHNqYpIWzaAxTuylnik7aaC92qm/EkoI9mF4hUnjyWgKsmv3FWG+1
dZQoezKlMpf/0jYbFBZznNRb71e5ckqTKx8/uy/XSc0B1d0PSgcJlNzRTkoy1wclvncxLFCablOk
e2A5JATA2PPMufYUNv/7KGY8jH+j0W/WUwenucTZZFMCVyY6YSMgzb1nr4q3R6J5hiddoX7mf45u
J9ANKtkrWm6RBO4Bc0J6UTUwzJWMWSgy2XWo2bSrojwnrtappGnL3iIHlHsUOVUUEXlrupxFJWSc
UmZNIhMASR7TGtmFDL1bSNAJO5jrUXMUdV6eo3wq1JdG0YmTS8fZi6HSmNKckD6fC9aGtRNB8EBQ
X90vSTxozQapNTBtLxkyzEzUtuel9kp6bV3IB3SJhOWFKBJzCmURoazA4qG8xgMk0PWxgENtAQFq
n5AKjdyQSUiVirIzcxZfAFzprk0xdCZtKBtmgxumCadC595VkbUC0OvYeXXwUeBIayjcfZJ7FndQ
C+eyk+K8od7O9xaQMMN6jU3lpI127dihyHyOp1r0GycIIiWasSlZ0plGmnUNWXwRU84KOyl9pQ1O
jry+ZoiA3zB+6/1KFFlsjy+0dbsgSHBzhjVnsCNw1aRMMYag0fDKQkgKiSoBUjlZu4ihXB41/sPz
dM1moFdt91nFlPSueCBftuHxsZyVzbFs1ybkJ0KRs+K2yi/Y7SlzKu+FcCoJeuVG5V5yGwX9PvUO
QiDRlNUsyPzWVGdrpxZjpDv77Mpi79I4MM3Vdws1IvGwg/UMB6Ae9ulOulX/ktoeAbWlcNdo7yH4
Bq1cSTj3yN4mqOJTY9nn17xsxlzbDITn0EZs6uDGhRt283jS5suS/qvztf2IZ+GIBPOatm59umel
wsOb1fv0Oati82r30oRR5Cm3Z4WPktpKzeeNbR1VZmK21oiqZRhHIA2Fcq/eCB3PfKg1yDHPcSqk
zMuzmwo4MB7yxymcZ7qzyV8FV/WaObPfjJJiRoZsSrcOlfhHm2PVQcUhkwAmDLcnyvHazkIwYajK
c2gpLLAo0I8TGKyXMDO7QSQIkyJrcpOUSrVWRCpBLn8KAxjCOb8VejMkFCN6K0h7saNDx9glSqAu
W7WY4o3WGB6DZLwYTpYvi5D4xOZf93GGNZ85M1/SUPSglZFlEpE1Fi4ys/lvodqjaoRSDAqWLI1N
oEC6X7mca61fBS+Mb6q0+ExtMLpHHjAZDdLr4/+8mA9pEtHjbdC19T+7/eSiuTaOfkLULwVRBG0Z
bc4UJSyiLSFxpQJ8WnZSWE4B4Z6t/XjkpWDUKwtacJFPfAspwOsFr8O6sgDEygnTbvSczrB3JNm3
xzGz0P1l0+1uknbHtOAY2K+bCPxKlsJLNvfrqRfq+nqBEg3JdyjI6oOSq0ed8L2iOFiKnRNv2hEh
URif6Jci0e8y9NLq+0zRi6T0nW1lBv5I748VJlEGttoc37bakKbkisR9WLZ5mkVb9iKQRZumwuGJ
8623R/9k8DiDD+TAzpM8JyHqkCvpUUg6m8EKWZotYg6il8dCPbGwLEy2SSsm+aGvSTkkhp5emdSk
fKeGHXJ4JFT36yEdkpoC4hY4jwBCdp9sWOpT5QBQLBzwsdEp3+UC/+NgvkriFhYIPqFjUFiCDOx5
FANmES1TuGOg9wM10XJWHImzTobxxTOoftdRkLfhMY0hCoMkbwQ1B0tuVQCeZIt3PvYyqjU86EwQ
3D6TwNfi4HOu/hiqTdD7glVvjUrIXwxYNwJl+8nfItc0j8DDApjhcbOP9lVyUjtXd6ihJjSPi55m
g6rP+RNGpRFC7C3aOSxT6/BLIN4CZhH/dqtfN+hvgLj7vYR3eDZAXEB8me51qngC85V9m3EIRPZA
FJEQn2HoxuIVU03NAi5QBsFeyd0SEaZ5OllGsYMGcU9TJu+F/trtcA8xMsVAKdXmGQn9nrMIml2u
6F0bugo1hG/DZzTfUd7WkkX1HQ2bC6e8xJ2TnJmC/yU8HrmfEXvQ4f0OrJTWIhfYD4NXKLtgJ1gu
h5ph8Ui6IG2PFnUmH29Rx4kbcmBlEvb+bguPFHhLIyrUw6kIrAR3fcybxs4iNq/CHuzYIMypcofp
FeQyNfwb8Pbjz+nx0b8uXwL579SJ7eFJn0yjvVPyxDBnzB4HWwaaTVCG6QD8YxLYVbajjDGp/ZBS
at2uC1rY/qA1MB+THGUeiV1vmsqY/ebG07U1b3NXV4V7O6V20+7tdsg6ft8rzMRrqvoGS2R0BqNu
lkFOzWR6CMPserXtOZoO2T86TFZHgDHIjPwP1XxJRK0NX4zYvu/BWG3dxtE3dvX7yjcCJnpc6Wva
BbpAMJytJITsFigJhoZexHkmK0pNQY4KtAvNRn3SvuIrfCcUsPhkNszztD+lIPRdIzynVvirLp5u
ijw3al+n9d2EzArQCo+s0GeMhS4uxN4jk+cHeVgaIVRtyxY3nNJVVQvD3bOAi9Fkf4FqauXowhBy
y3mxa9fLac0HuIeIz25x6UaxpOo3FJKX4CQQV3rMD6Yl2KmqgHzX9swl1EavWkLSEtVTtnfdHR8E
gZWuitGrLInYdO8xng7SJESaGatt+icaBzPl5oG89u8riJtq/fYyQ/0JVSJqkzFAWqI65QkYTNgx
8wWOAtm7WRCGW3ZrWU2oLZ7H8ox2Igv//6GoZAaOUFs/1pZng2Pg+6S5MaYGtqwz7fNuWQ5qo6zg
+bYpozMhyLLMaU9cVjkHEQqNCba3DGUYc5dWR0RgT+vbokmsYs4cbeCL52Znb5fjwC4oT9Z7XoCO
+5oJlMnh15nnDDVTtrsHIPgUKK4uq/eUoRcbAjPPftdts5TO+ejunAA5JzER1y2eGzN1MqEgKIBl
jrkgImmUQMQQdKtDgxDQa850tE6KuSrVLVZ3PVqDlMvpSwq7+oFW9cTQ8M8qHBSb6pHFFNGa/7HC
e4oVsp32/6n9pscViVIxif/d7Z4yOuLl2GfyY+r6yAUaBLAkNucoE9ZCKZRyDe3XIvNaYSmbbxh9
aP2q9g/RTU32FAJU4Q+Op7QYX/ul/38VQ8/A+NrpqjF9evrs9c9He5lqsr59m66VckFupBDRffCG
fdXC0+AI0fAGLpiHNCY7xw6YLLZP2abe7Gb1GzXvFEazkRdqEnlK5skOjlMzPqb053OhSQYntONO
FA6O+AG01TPJmW6kpn0Gg1fztAYMa55uXy2YhaMfNfYq72hK7q2vLy30mbz0BBLGyKsEnQeDX8JK
5dumsLAAPbDOAKTyPHdhQVgI294WHLOFQbaaSvOzkX7ycZoyswh3NbZeMeEV8yToLMtgLWrBXOj6
cSl2XvOUAtpqJQbXrhkMR+OYcJ83NqaOfRQFr/DXXiomR2ZNnduK6qhP9ByJSZ2c/8YuRLHDynbF
9b+4SN1ITyO/hP9ey/1/12CLW85yTMT6O+NCJJWmwMAqrat1t3K9YkTb8V/YUTY+fZR4DQJ7pwGW
D9aUJ5lhl4bceviSNUD3PAPt4gMLk/Qfng5/52V2jdK2Mcmy9SlNrGRBm5HBhHT6FjSp+KUI10rs
4M0Elw+fsRLJgLF8RsNdsntLHWnXFR1KR5f2NYnIyyc9NeHukgBzS7wJJiFKRTu9RjkwJ041QolZ
8hLKBY0bbO/jIbYs85FRYFxkBLlNEmpJoCcmfHaC+12BQpLHqjXi/pHCjW7qBYaInLlusQLcPvZf
Z0itO1QgSLUU4EvvXeIfvTaUmlW2qReYtBS5fLRVPjPQwcsXFg9V/2o5PCrzWam8u5ESr8HxzQL2
chg6Sb9ZF5ysSru7G8cuCHmHFjvBOURuJqZHqyAJUhI6tKg312MZj4/Bgx9JjjSQiJ4gXZEXJmhd
NK3Xh6He2Tyo8MS3wfI05CAZ2ltBbcZVr1xsaShXVdE0KtWoS7Qk0R78/tGoXysd9sX/zum4kRdP
jzWlMUenycEUkB3VcwEcbrtDzrEGhC3En5So4QKu9UJaM2TJQubUbRmclwm54Fl2A68pBPX5B3Tz
bubXCBVDtOceLefwIN27J6jvlnJR5BCeaA/q9ieItGbYQ96onHSHUZtYH+lypfsHD/x94bgdNQrE
G+ZtK5VOoywFPQKLWmnAqCHXKbUiMHy0eilTOZ3Ikt0p/Jn2QE14JsCWlb/lgTnoAW1qewH91y1k
jxjadohKUr0oz9hu+bD9jEH0Ju2nRodTBDttMV+wc+9pY3p9DZJLQ6zsgfA+vC2Ls1BACH/bXy/U
hTeq4w/p2jZMbUPGjg+OLhgCrcPIeVoYcdcKK3DkXuH+8G/+Jn4Zrflp6RDx8tFupOqrULC1pSa1
AGqLXwcvfKcevT0cJeuQ6oRiJe4rWtQ192fJHeJ8SNM3vBWSh/Rk1PfIGb8YMGfYjtJymEU2tSVy
zZLwEd0A2bKu8CzOQYrdaiUiYw5f1nxXwfoTdtfvDL3yB65mr6YlUnu/EMuWZ51D6XxNcd4skeO2
GuEsctHSIjjihOspqZ++CCg/8gjIy3Tf5ZgZzo8Lwwup4ppmArOa8PdJnHCLSnn6zdgpKed8nB5M
4in2DZBsjLp/tJKQOn+c625Rg0g3d42Nb2nhIl9hZz/vVIQT17vMSB81pd4qVB/N+9gGDqNZJVtd
0Qsm1Kif4a2P0Urr9kMjzozRFFMAjkhQBsek8FZC0lh0+iTZGfuBgJac4RlsezS8SL2AKVxkGZFY
qAddGijTTliOfWrkAFEvU1I5ft4r4GZ8VegSO0pOpB3/Ndl1sli5nSmrbPvM7SnZ48xQE4RVIA7O
apc6RRun5hlguNMULMrzAJqfkluvP5oXwqerIweuFFnLNeElONiZbSphDuRpIiVwQRaM5KH+wPuW
SlnLsqv/OdLVsXcjHBgNl3oh3otvrYRmsCuY42kc809P62RwhdiT4M/IZKYsuwD1piraVVzpBrXZ
y5/EVV1u7Lpy6LnfLhX7Cbl7gBomIKm6OClElnBaAgQbqniLuWEhzo2WOCQ6RZSvEWh61G1I7Cul
tF9cQXgbg2yHl9ZRK+l7BtBBnptf4HCuKRYin/CJsm8+gnDilhLzS/ITHmvgOEu281JoBrN+DoSg
eSYze8t9G9vUTN8C/SpEjlZ/tQr78cB2HrF5WlDWn1315rsfiBw3JFzZM9EFRho6DZxxF895Aiea
MgIcRfUaGsQHY9DbQDacgjngenrlBbjMGVvQwOVnqP3ZJ1fe5+rVIXov1kWrAIDLD0Ecgn8Czxno
ojCK9zCRwDVWklI44ggNEHbfydo7UZQy2LnXB3B/Ci6mcSXi2nI2aCymtFRbPkSDRpIBlHOYUGda
wtkg/+i5A/zGd87ygfFHuvx64y0vCvzb5dpAwYO9jbPadwpegg7XzWBYPJWjVIzmrYydUriIViGJ
K7jH7IDeAO5Zdlb5e44htQMXLDa/BuJnrEP/1IHpXfTvSHg7aNkNUo7CyEuwOLGxs95f7R7DzXEx
R/q2jRvyl1KQDg2eClOpblYrhRexmp7sLLhaEmnBwjjHKBrLRkXy2w4fSLN/TMByVI86t1M5jBdE
ymsruyMELhJAOtJPZNEOzPDaTLcW1Zlq6hRCCb3Cs3w/shv5gRBVuP2DxO8ZfRteKIZ5hn79Tgfz
rJD1hBl4S5gyGtJQSAst95zOelJ3I5v5YYFEQel/CEXvjovJkKIeaN7xc/GEQJCEYpa9a4h8PSHi
of7JrdiGifJ/yz8NoNtOPARckL9yGHDb+jTHZHu9p/sb6j0uqwgZr8hh7YXm5k3aptSZg91ffiCz
k1Xf3ZpFsuGAP2SDwSWl+9NzY5GcCoxb+Mb14+7VEmRu9NRCPwm/hApB8oGjAEWoQ7uOZPaHEmJw
sYZ3O/TqWqNLhPy0wBop/ir9rg3UBsBAAKtLhS425HamS67ILXCU1SFHr4EQkr/C9UPeUrEQrXpi
nh8Rm9soov/0V9PRX4T+YDBrsE9mdWle3h0NvSgvoRgfa+QOEACzAfqztSX4rT5Sbg8nhD7nbP7B
/BoPqshKc6w6Y9FiXwIHlOEMBnrguqUjRwAV70kDfO7HkDWug8LmP4ArCr6+v4pybSxL26TyRbrk
VZrKaLKPY0aY1TjsSiDTaXTpi/e0bi9a9qQEO3ndGqbQ1erE+wNfyegWSEUA7uoTedSxbJycgzST
wdWJnaed3l0cA8WQWl5vNcD4s4v2DTo8FsFhHMsaALhEfs1pSNYuo8pzsKY/Q2ViFpPAzaNHtQP1
zcwe7vPL3Yuj5Ybkb//uhgqjHEYIbQv50IWX5dJzXrHjdPq30rPwX3CHl+1SgfFLHoi18FZhHC8G
6A1YfDk1zQeGAqGVw+Jhm0kPRX8XhzczDF5Lnmn0VyBULPe3boBi3q/PY0bzI7OE8DPYnfPK2ZQm
YcemZmDGf25TyJ/RpMEF5oDVTAt1d8Y+/f5gHNAyANSzJYkbyg137sPOQjJ8//Pf/it3SSDWLpaa
EsThSzo6eoykw4+egCsnK42yqlDV9oh/1r+WRrLpCuX9boV/ILBs3a51k9r6lsRATyVcasX/3wa8
1KYM25F/0l98tKeFBWW5KbabdHPq8ymNc+u8JyMBjesB4AGXaVpXfaYPU3FXqI0kJdvilPQAW34L
e+/3xEo51jw662a8KapffXMFlH0jm14siQaqwHexnIMAMPUwu4b/FbQJYOJ70fMtXag3KQMLg709
wM7zCvGeRkByk58d02rLQaTj7wKeq2nz8qzKASUEMgmoOL2UAyCYfZQ9kluacQoT3cKx5yZ7NAoc
/HmJ9barISrhe/nqUUJw6HBKzUtuzwzeaDqfE2jRm4L+HB1Awrfn+2R/NXv7TcS+6cc5IopHWZs5
fa8vJH1yIEgxKRt2r/+SMEx82xi5Gk80/VMqOXFrFkIFHDRXUFckPShue5ylE92Jx61FCkPWlIG8
uBVqF+8o3XJ72gujQIqr+HWoND92ezTci7WP0b9Pb77K8bpDQKSukSjnAltDzDCchaQ6GyR+UhYT
eK1y0+Hdx/hvmb0oud+Si6DGIrUZ1lMCm6wd9DwYOSzAGqlu5JrlDhoPnm7Rg1jypi2vTCRvZ4gW
dGcv19pWcR67FoygSggo6grhgJK+9br8VOkG9Kwj+tCO+lBFvgWqG1f+7KtZHF3ydfshbzufdQSp
mRcztqgMD9SDCJfVV4BygeHqGiMqe4QbWSFGl3CwixmNrN3HKWXEwEZjcWM7IGre567pfULz8BuY
wJ0wDLK4eAEhPJQeacjRSMkV2n7+NNV7/AT/bDNUnHI7JLPZXVANpnOcRvzFJRzOj3DjmS0o6e9B
ZhFjjn6zN4wukAJq66+3A+xbH9Vjw1bNHfh5ZP/AnvO1/WyiH8+6EOhUyZk8zAC9v0awPm2Z6gGX
zd11h2WWsffbBl3O53K1ygurBgUOa0MKdYLfxBJSdXq1wEni/lT8Dog8BciZxSbDmlOMXubcKGUp
+IjLmfhl6ijSqXgPGsYCYQr086JO/etrKI0hHvahIwcVxMh7ICyD9sYHtmyGJo2JTbcb09aU3Wx2
NFPJ088h5fNtWQg4IzcBfhq8CioUfMnCtAzkFadwwgGkvCWdpS70q2brYyuxjRyxRr6WPk3yGWh4
O5syTRlnj2AwyCnj/cv9GIf7ICZ1Y44/alKFZEJjxIz0AEH2BcIX11/84hBv5UOm2Vaiq5qoyVaT
UmkAFUptb3WBf2j30EgZQIS64sjzmkXy/7al8gDdUS5NVa7uO88+xzRNRTDnwn4pALXyTpiiFHf+
NlqyB5qUlEZAEq5+F8BXNNGxjKdA7JKSGleu7/s/H/LhYUji46ppKU5r3KCtnCA/SKRSgyufBeAT
mF6vcrBI+MFwxBU8AI9Q5VWWIYhfJ9Tgk9xQXqwUWvJ95NTOTXOSBObmSqFu5N3uhOx585XN24GG
CN4Ucwco7BHsffJ/Vzf7gcJZadD4aJvt28sFsHyfUS90V6Q9Z1P4xuLbNloEJrb9oKnwIY+PrY1T
qKTwVsyz3IFZMG6ZEUA29UMn+96s+zC/6FSE4/uWRA5anuwcCA+x3ean+ofBcXqHtc+VtNvAVv+2
T4MbWLuXjkIxZ6dQ4VcFbNC7OEoMdEW9Mg88T/XSqL82d3h5vVHHV+H4+I1Lq0jDSU1pPupDFazf
sDMVgwyBUu521el+dvzRIS9mm5YZHXdHAVFQ5DZOWOuMxOguI/3bAgyu+pjye4vw2aWm/1KUypTQ
yqbX8vlHj4jVw/OKly30QKor9z6DOZu+zzSpz3PwZLq0m1/Dxwqp1ltdNROY6Egdrawe1lq/ML+R
zDqApXZqCg0HMZghHHWMymnoh25LXx6oqoJu8hBEjf0XYrhcCEeYSUFZhGsKugUboGKwfeANyFcL
wcWCYk+OykpjNIMJkre2bzjxXaF3BK9GJ0HW6FMQSbFHNEY1+5rkmvgOn1AU9WG9YL+1mhfnZszg
g3e4EoXIppKdC4ijtRQjvjo0GnbO/bgYEjkO2DjvPU0gdERHOgTD8wy8ZYVFd3FoeVBfbAbe2gO6
k662PIGodB4XayruHn4CvEzyE9ZYXHfprQeCsbqP26oYCABCUWJxdNe0NtVgYYR5pufrq6Rkpb1G
R2hiMTvvG4Ir7uUxQegXNyx14AeHLWtDSaI3nGxDpo3FUHcdoz8Ims4x9SMgwmuSMAESpGzAP8PF
Jh4Ipa6g5osI90N3MoIxJxd6rjeDOlzOXgNRN4YFj8DEQYmRje8jgJ3vE2oT2VbR4WJ8Zfk4R0oj
8gk+MrfVdPus9inon1qOJrFemeyUDUgUctjBpRpgr5EHUkwsrF0eRDwSWZcF+vZ+Ez/39vUQzHNo
CRttWSCzgrqh/Zye6A0bhoh0FyjxCN3+B4XHD93U1tufGSSYRNOe7+bTdK55xVP0nw/vNbGXpyr5
iY66SPl5bOqg6ebIkcjC7cREOSLX8fLSdcdGJnlRVAp9kTstk8m/h0UUAuyJII/mRNaLOf+0aaiV
Pp/05l4PE5lZ1+XAqCzMx6ug1+qLXsqG5p77RnYDiHBUA66P3z+eQhgjmKO0S/Z6l8jvTvkpDMw+
LS6FjmnKm/GjPjYuV8cjEZ8SYrhcLd+fPQLE8OHJm7F+T/ppgVkrT1YabMxLPVvVS49aqErSMsnR
xws4axkpoxU0/yjID5LVFjJrPQ8emAy5IGYDYKo0LkqDGhYuR+NYPQG8Mh9TVE8BcKN4v9z3/n3x
QNL3UBXNibhWWh2yNJXDZcEHGqcpcMXY3DWYds9U+JWHYiuRhFLHvfkq3P5G1uXt1sDQI/lI1rJD
Un3H7SgrgBRfmfxAvg4jLTP7QKnQZjmvBCuiAm+x1F7llYPyRO92ggQCwBcLMX6lwQstYYai7Ano
1V4UiwnbQIN+54jGJ0Zkn/aPwmZUeWFecsXIcRPQ8VLxKEnN6EobhaNsJvM/rpHYcyQjvWATharP
/0o2Rw2bSpVxUQ2l6WBzOvwKVsT+A5f2+02Dhe2sETla18DgB7ZGLRzgIxmImavUdfFVahntguKF
9EtBg7O7aU2mgS24XdsW0I0vqDPkv+SauBf/p4ZHLU3bMQjWu1S0oSEV+f5oYoAUL5ArElDdKzjO
hxZtquS00EDYveiL+WJGk4wZ7ZXaKbVq1/9adMcCyiKsit6v4RnMgC0TuBl6XlmgyxdaTrXKqQ2E
g06L392VmBzYA5bSqQjYhUmA5OK+gRTLkwybpMpODHleJhJRlQKJPXDT7DDsWCok1i84OPIeBZ5g
5W31jpbQTRyHckAosQwhfL3JfXwgqg2/6kaEkKaJHzSJ460XB8BvicwWzuvlkkVZOsbLoxClo2r4
S3L4RCnGbkGQGPjEpxfi8/Qbpw6otW5b7ZEyiMRQRDeUJEoVJ9QnacvnprfJJdOBcGgxajgK8mgj
MwL4nQeZoIaXHdvOYms13eZnfwbkwLl96nwUkgQ5aG4RJvSgFEhcXmXga26m3cMYn3DtDKss7WZZ
8ghWOplN1D4mRvPE+ca8zQ5YuQ/Ecbk+ZLakcfvr3SORMqEAq3HifONoHmvJRwG0Ye0n129UCA85
D5CcWVNC+onYliBHmJYOaXMCD6zIyd3OM+XeNFCwRuYLjVAB9WAux2upBIXu9eLVQ0aqiqJUjH4J
tVIzpcewGYMfzwFH8pnlFGBn9S/ShqAozXgb5HfHRGMvF0JSZDebs/NEve6XZcACSvaeyQvodDpv
Z3QuhJtzfUsNIjkLj2+Vr0a2bATezPssyOuy+sxww3AhLGB8NvaEdcLzQj7ZTSNaXo4UsxT1goaH
hQaIZAjCSaIIP77qm/hHUEEiETucV3+2sb/bkfXmx/W30qPs+5vva7QgML9sqYVImyD76MjkOORs
5k9+a6T39E8usNi/Hc9bhDW1kXU7QZYlOm1qKbvSJiLpIbp4PkWlSh1B1nEbB9wQKxDrMwdA3U80
u3p75M243lWhFPM5y591HZ+KyFncX0naHe47JSeEHkO5Hn4VUSHtKWYueXgHMDBJhQpq3sUD+MI4
1YtsIKI7nBLNrZSZH759rjA06b5k9KO3tqQIQJuXeYDGSjJRsmx+zY7RqS5gq9fYrSb39sOhhLsU
9nuzaWqK4ph1OyZCt4G+/T/TnIbfU4ZMODvWVvg9oMYZQmpLp15hxT63rPCtWa89NveotmiQv9ct
Iyfq+EcELzQBVh1WUIXQtWPHRCkFEUJVJQJBYA6x1hVlkfHhStDn7nFV6N+pylsgzjqavmsQgO+S
lhj52IS8KHCjgWNF6cXP7srruyqRCkrmJaE+PBUz3FlxZ9biq7JLYG4JQR1qAieMRO5VZ0Keg5oy
Cp1AwYs9uTjQtP30OHIbUiXpgiOCfv7o7f5m1jA4H3T+e1LKQoYUMj3tXEmK2R1flgbsVzlTEWfv
26ykTm6l+HneimAfY/iHpNDX0AHRnClKZcM3zUxOo4EIb9JrVuOekXNKqvxC/HR+fuD50n/9r9Qk
a0YT5hI1/xlTu2KBLpYdPPTaNe0jxMtLd1tIW+vDzCtVEbZSUIf5FKegkqT0LbcPjX+hYNzGNqdJ
kSLHX18wNUghdUT7GrwxxqbVdoo+Q0PmVEXF6K+Z/3pHgurAF+CIu9ztYA7O7JR8LgK/ABxDBVgw
npTqDkviDrv620+FC84S3eJIQEf88o3Wi+CHSDE1GJt2dkm26Llc2yQZTF7lyPemyOvRs/b3en0Z
Aa/JeQBB63h4tacGnpaHFbwleRRyssKK0l0S3gtBW3f+Tf+CO62JJWjGW1eCzUQn5efjp0xHKYyN
xeiJMus7GIrPzKfdzdZ0xJQZmwOoAJDE0P+Jw/45zSoXBgemRM/hErTChddBh8psx9++rFaGnDRI
aUjHyol6R/EcWvcja7GQqImQtxetHZ/MO4TpTskrMQusIUKHIhl4IVF+yN8yWWZX8euu/FXk1EFn
xB2F98cbOAQdO9S2ya7Oy1hVLDlemjn9go+iaJCKU8EUVtDUxcq7Oosn4P19fEeWP/Ic9kTJaAZa
AFie1wwk/gdvNN8Peu8PPZKYcXfPYE4sLxBt0nqUI6u7wdEHjDd7W02E6lPfrlv9S34eYwB8v37J
KhESjNCaDPcimBCiwxpV4oM7WkYDz2mwdMWfU58E+8cLfEBCclxToO3xNJf6pBS4i56viPc6RgzF
JnEYapgF/suUK1j+bC7PJCD6yd6Sk+PEAKfn00DfTYei+lP/ZwDH4vZanl5awNWJEZCLxHpLJkHc
4XFBiLBGEy4evfemrZlc64G6f3WdnakQ5c4DDG06QEuKJSsUPvzlBXxcTtKf3zNke9EDPtIHTb0g
LhxEEwku8ODjzNF+yuoaD8BwETptbsm0oNHMbY5tdtI12LKs3vQ0SeWU0UqIXRg0UYmmhlcV7hfJ
R3VzdZmLwAHg/aqcAAgwhqe1K5HgsRCZb2LwW8Xu0TwO6hcvplxbiHBq+6ezXdPQQQFIZFC/jIYk
OIlP9bRi1HXK9/HpD96eJNLIaLqZIhWXRiSuWhR9qKmmxxpesCsz6KVsXOBPNW20iGeJuVntqPpy
TeVOIo+eGJHAovL/g8TO2QDhuek3TvAMW1omYFRwgBGWZdktaq6feuVdf9f3W0CJYdxpSvlKlsW1
KOsXGF1cIJcMrLIT6i8yom04pZBMKXQaEKYgvYKT2AtvG/WeToD6J3jDoCqvPVqEyUGasxVI4yY5
Pw4VFOsRKMZbz5zXV+7lULOTKY8LGvnBk4+026ne1ObH2E0KyGejYLrUUvJxJvuUVRt8sH5U0Fwg
+0Jxnyyh0xEAEu9Agvi8+KmroMg+7Qy9QRGO24er47Turb3XT3X3p4rvUfUSSLlTJbLFOVbMvfFy
GaUTgOJaT0IBnAM/1W19XDCtjDMOqXtmpX2Oixk0SGhP3oS1I1kElbCxg6vpkXHOcoE/QVw7syqR
/bQ1aHXscRIyJWpWxuANixXCANMEDdtkcV15eGGO7aBjaNJgZ5aqsBd9GzN+dI0E811k6zefQX8C
4KvH8LIvd3TsQILflKreU6fcfoZzTuJ7u3oPtpidS9/AjV7bOjzfzMCPhCP+QIxt2mCkyjm5Tvs3
Q67XKw2vHAG3trL77tb6bwtYCYo9XPY+JBiXnPU3jPxejQNlsA5DqUacgbBlq/+I/V926eyZf9mg
CB7RwEFOBLC1JXy1BE8PEEB2HUV24FI9qsitYTNXh9UmiB0UB6S/LAzAd4fgoTCnabmKDk8zNKN8
xBSTsA96qjkBlxH10yxNh0m7Ru7rtEqufJnM6j+k8sH71y272eKG0MMSosLXDisURAytOrMi+eRJ
m/QOOBpS3+8IX0AvFzBISYr2UawUaPVDTP75MiNXd5z/4KIfZ5VJyWZsnMAH3uKbqEQEWzph+b4m
ZxDz3bBO312y3GWtlvpQfhdT/qwFNjYVNr9PZ8K+TystaVhX3EbnGoT8NbXntsZiRAI1O/7KOEF/
rp7y1kbnUv0uBn9V1AjeDTDdcKKNlMDvPUtvrqM5694VABMxccUOsh8eIFQXoWeqQBUMqTtzbFJN
wA0T/pWNpsDYWO8rMFjR/cIRfE915c5VYyn8UvmLFysDjDknKyLlNiKeNvjkTwxCy7qWCLb986w5
rUTvuTkoowWkBEtzOxk2JsP9Ayr2ojTVF2Qz3sWKD3ASz7wRJwl3Zy4gbHYmSAWqun9L3gneesQs
t1xWdppNuwISQdb5xtg2dnnnB4yo2xe6WhUQPGTA3nSpP0rv7jvcCcrCv1O/oG7XkPr+61CH6eB4
A1WEBo8t5aDBpRIRsLPLSbFXsWvx6hlGRuI4BhXe5//n3H1WexmnmoyexxCsZ3gH/kgVAy3FT3/C
aKnp6to2aUdCIhqXGjFuKwpQ3nIkVBY33HF4XrcpyV88W1Dbxs6y3Dq+DW5yMXtTOAheSC4CjgXG
7Y0FxDNwoOhCv7/33j4K7YgVYPTYPCalKGmmmSe9gAhDv2IABRU+1zWnv/RqzmjkVrfMl4keK7pX
DOHipqTAbomN4ITWEfW+N3/p8bx9+2ezpXr63NYuRAiIj0X2cqqVi4IKXCFgU99KJ0fB23ae5ERM
T02doN41TRDXZ1mY5Nebb3jAWobpMEYgnLKdZjC3ysdfPp8i8gkeSvTPxBLRcWKa+ufKK2OXyg08
TCf9NOXOR0UY+uMSZH0ctLqylGnGmZySr39M1Psgcn2R7kp005jIdZXhbRN0an6aKINEvsMHF0dl
lFtuYMDmAxJrBEjNDN925/AiW7kD0sifLsYXl1ie/pNvEW2hKwa6jLkVawDPMzAQsNa9ZdVj7m30
7xeFVHmULE3YXndptM+v+e/AbvdxeiK5VoB6qv+k8PrCClat7CY5I1hAlgi1yZfXR76lTxwwQqdK
1GeAcCEt0+tTfy49gMRsZgxPE3tEgKEgSrscXfj3FEOy3wqxnAv5p9H0WxHcKryseQ8NdKJ6gmBJ
ce6fDRc/OEvEkgaqeTbYagnj1co5+5ECpzbd++XI48SnvNbf+7nDUM35N0HAS7aQ+BXapx4bNJB1
QO9viTqMhBllClYZnzL45kIidp1KlUkS70Nqa7/f0MJEolORId7aywF3siT15G8BJSr0NuwEMVrD
LQcdy5VsB3nqpwsBXZnMGXd85xD6YrjGRfgXICE2d3YyKG06dm47MO8uaXN3KWlOPK5nwzNI9BA7
YZWSoVz4YDryjJuuBQ1WqQFEWu6yc8m73mfJAXy183CKT0/SPYvZ6TABUT8VG8cpufz/lNLFGffI
0NOCXUJ+IbqZRBCbs6YPph7MaoLK6zds62w9FplNG9cZhrnq94guJoX40Y4COqPnun+iJAAtqiqo
19YxQMp57sC1J+S3bzNjeIxzJfgOEEU5jwAwwo2NYF06rzY/TbBPkV9DafcHdo/H97A0lT0PmFhR
B9XxbCG8pQfLXY72YWKSyz/DO10L3Czvmd62A2oeI7yCyPNAKSswDTK7v+RoE3taQLsZy7HaN3ss
J0gtScFKpt4lWFWVOjc9YLdUz1JnmfSdUGi0tu1TwAyK82j7i7POYAPpCeHwB+cBOGZzJX3sml19
/6bkgi6X5CFT3BOAAhMrNxrAKUv4rvj7bRDfYA4kmPYJtdTkk7WmHsCVCwkHgUvFBx5ZVWDPQuaY
NRZstWZ9+xKoOpQRGMv+nUGZV8MBTP2wzes5wcAlnPuXyruNhYTIqgDhPzSkcR44WUSr+mNWCYjs
BgD75tvjd3DlA8k4VOP1aaHPnOPzqmzC+syJXxGyKoranncTQ02LswH6wkndUoM0cHSWwPgpa4Ig
4E3OXJepWpaFwMbr8IMqnmguXNxlI7Dvs1UsmpRsdadNtsygJybRzzgXJOZBJqQUbdDn5dOZFntg
YxoDYYPM4tXgCC3pT87PzncXYEa+Tf9aBOrpY6zEwysQIuurJG888Vd6dXTQtd4QfBioFbd3g1Xs
gTtZvPg+olysnJL8E1dLtCYXsuU7dNsG1eaRWkYvZuOFNFzH2cBM1ef9XcT2lGHIxLBXoXPXiZtO
+nPIwl7U2PV57c6hSFN7x8CfnTs9VRuyLYFRsyDCcJOr4fHdNuC4Uc6DK9BDfmJ7gTPi6/bRFIeH
iZSSrpKmWiA0l1Q8pdo6Wu79GfWKcuc+uq9zkdCB7s+emDKiRyUNdp2q+W7t6QMo7EGO95NEnyDY
FvNG6z3u7XTEP2JkHEqDR5N5VJFrU0JMeHYXe6T8cR0kCmOC1+Fz2Pv2UBTSi0IMKabKclxl5YUC
1XBojVerwq3WkVMKeGyoHQ3mhziBOBpsu9vHweXiHJEgcWz5rp0CZTkMA7Phj2hkcOS1jWUF59RD
C8biZ7a9urH3B35fSBEZ/vG5v5M5Ib6hmbU1/5qqBm6r6ZRpeh4K6DTRHAEwDK1t0XZFFmn2yzC5
5tOh9UBlFTQLXbp2/EhetSJqZb51TkMotOg4noFaelUqN77evbR6OdGduKwHNttn6on5VYdR7tiG
UJ2lu72esHlvIg9GoswfviXfzgQEVGSbP4aG2nauwg8zGjxYm9aNDFD5MJIoCqTZG582dk/tS6SS
5Ksm0tlpVv9xSqRrxlGAoJrU+VCv3+tlKfp0WTJFIs5gRQpe7nr6ZNnI4CzZUg27uVVczq2GTUGV
wE2bJdTdCK+ui0dAM2vq+gxzlpaI2BKrrVWDi8nVwSDQ8E8OEpExHiHJbRZKHL1kzgeVMTTzpB9j
PvY1GbZjrNXPFzKz7xV3H64nP1AOMoHrNLLYW2PDmBM6FV7uhpsPqsUBMbxXZkWlrfA0gaReLDmh
EZImGo130060R/qMerA0+UNQITWYINP0t0Xbl4DCK95x4VeU0J/I2235kfesxKoEv/hrByRQS+GT
ArV5LXj4AYZiTm0AK8uSDlmihIa0auzl0ky92mkRvrnQr4Ubi5DJq1gvQjTe1S0V8mdall8UxDU0
BBAJ1KiiQaMM5tl+br1/Hd0lakZcb54mnyUOo2iSZtYQi+V9bIxaeqYTsb0dMJ8v+UK7BZN26wZB
L9OZH0ATcXKSxBM56y2NlGeAsDzAFX2m4jdxvpfrOEC1SRd+EKXC+vQHqV+ejcmikTmaabunBJ7w
XTklBnKYGAx3L+1sHww/mt8q3LJtMabH1ks2xmaaD/Lh5Fz9ADL71/dph/nP5lleiTP0j5qObcjY
U9UtOFjcHdhLqbf4TtBVsjmoUVBTZ0hWG9SrVioaTRdjJ/CphuHqWhITDADOY5yeYqZeeg+St2zw
iJaB2M2aLQcgf1ZXHR/Yt8z4GbPqlfWyhVBGETlPrHYNHhWH+USdhhLQcc7ZbYKmfQQNTgHfVOi2
WJ3wl3mU7ZH9XO4PmvB1+DqalAHiaulWqBPisd+s5OvlPBWKNx2353USUa98RxbbfX7nmezVIHNX
mV5Vt9VJOKCYofnvEwFt3WoDgOd0ILfSxZe/7CesCsW8bumxHF2g3IMBibxL22N5kin2m03VelFg
MOu02jRxKs3vKoL2bT/nFnPk9nqrMySRrdL+i376G9H3c/4InpZ2Jlb4QhiLouSIPqvC8zEsQC7N
p/ShT/u8mUnQjLWg9Olz7TEzasIebqccUv7S8WjKqxcm75VSm7AFDMcw9/Odrt5vmxgrkXQsqpsI
j35m9TQHEfYgmhTc6tUp5q+Cq+deH3SnrS/PJAgnrLMQQxJsHPhNpc1M8YUuZ5tU/39bZ0uWp05v
3To+7Y+k+nNRBu0zKqw/96+YA68pv4EFO+Z+UJ5Yu6ZgHhNB6J29qFgmVMK98OmanD+ZjlIO9iLM
/e4HVjLFbCNThDUQbdNq1AfFBNGMIVpDWgI9CRuyrvsaYdZ1jD/4HRvzjdIYbp/GlGGisplbwE8f
RWnbczhNGOvM89tdTAcG/qYvArd0Rqg61dzriIX5NWeRp+2eIixCw3vR4+va/WRUZykHOOLOZGSY
fOkjei/jjplLGpeZFHxf8L6JpsAvXOh0eeiwcLWptdK0mujwCYw2nTdoQY7PQSuHU6vcXKuGRD/P
WX8Hde0WXZ8gR6QCCZkmXvBlgxQdJJyKxYAa+BKw9NCzT/4tAHyJm3LiY1q1rcDWNZsc1ocMgQ9Q
VwIDdFDugw5bjYroO/5RdlsQkzhRyCLW8y0dZiybL5APyarsUMqcZWzpLFyMZjJiP+XQzQzdA85o
+PoxJAzeO+ibE7m4NCGw67GsZBZc+SgbYW0uSmtym/MKBu2CQET1muChcHz8D+bM41u4N1q5C+uD
vKtjHUQfhGdkJEZWUu0BtBwWQ8BwcDPRwQgaebd9h/b/UFNYMn0sQfEad0V6E/C3gxoA23+MaWdd
1WaP1Yl2PUTaehCoxJUC8tqhOaAloJv65JEnUu7EhcziXRmQdmUVbPTNfZT6o2wDbHCztTNxlyD/
3S26Owp5ByJhOReotiNtn6uDD+RiZaWOSH4YuA7RsGQcnQRpQq+L14oW3M9p212q+EXRu7G20TgN
cbu0qFPaQpUA1UMEantOQ4E1nAkrwD1oWplKQwYtIkLrsnRPnXUpA/9UlXkAZPeKayRtrKcd95OA
obI+jiyjdxg8k4Dx+DPxzOFCv8FA/1jTjCtzT+B3TOlmUTxeG+EnrsUMZsFT4ZfHIvE0KFunRs5f
U48P7vkC+wLK11Aop0+HGLfH/c5/CzLQHDauhj998+jDtxED/SBOVNj5zNTnulF0DDlm7D7uTIz/
mccAww9AZ0SR+qO3OlrM2V1GnXSKbqpUJtMcRZ6GbVUA6iUCPkH7wCFg60rnSnYZuqJAXRFJ/phJ
drimRanOSG5LtKuQ5DgmVxSvu8dkinvirj1Q+yBy6sM426WAnMbTyviT0srgH9DpsBuDY93rky5T
0qqwhpbzPrmqQKvW5cKd3eje4cT3mo9d5Ja6zzUcMoBa/TnMEgcxlstWQtXWCQQfETEFrmNnlzQr
daEt7O05X9FO8762jpH4Nzkcy/1LJfQILtOgOeolX2SzjxRMRpwbTvNEV0mwaQP0JwTAm4acW/NY
Td/nCsRC2icHhEGsSqyZXXY6cqgkAzyHfXLYRZIab6OvWUoubGL4kQ6R5bvP84iFfB63Q768wgUp
emQ91JILXGipqgfPTCA9qRRq3/ZVxLwQPenIfikETF7x2YgSov4f+7hdGBr+FJEnxi2scVuL7GgC
nrnT/LYfD59CqLxtqist/q3BdlpYzs+SlvIuuEcZUDjUiytr7XH+/SBN+2m2JH51dn1b2qJhbBBW
j677hX0snDMsF7PR6e7mJxhRg9d7GWbClM7yQ8S7X5cL01ugJblXPnVkPJ+RMdS7113axtF0AEe9
flFD1IENYLy6YTyXtvywv88LkFK1Ub+J8n9+DvAqOfqQUh1SPBo2a+gZJX0zaMN/EODKPH3d3TMr
JpZPvk/pe/fgt1Dxzb13RRHLW4oWqzEC7kM/H5r9cfMVIINIg4n4XrtF6TB0KWjVvSxR5Amtd0fV
iaGllCs64ohmuW+X4D27RwZwX54jQtuE6wze0PMqXWx6ftYElQhs6vm0EUHD/g+mgiKYNIUF5Bk/
peWoQZgslfKTqxpolhLkbClragvAm7ELtN+m/yeeo5CDAHsNvygxI3hNrzWuFWJ4tP89PBbsDk97
SywKNAiCVqOUytihByLkF64eJcc4Y9++n/RssnXwGS/KBzo6wBZPymt6VLWMnV+EWdHkzj7d3I2E
pE/hvuIIhWTxnKuVxABg+A+L3mSHuLZQnlKBt954L4aqaoeFIABXFleqqFVFMcFuKiiPd71ExKFz
U3gKbwGe0Vzmj4vMY0X+SM0Qqc5/O3gcKNqbcBoa6ZRTbDAMqlqK2lx2gbNjz7JBA6RpekJcwIz5
UMKBOn/fwKBmkT9Y1YUjwmDAI5hsClD2l71MJrW5aXx4SeQ+PuEoHFCr5q0hbDEutH1HSPpAjTqV
rIbC+56UleZUDJABjpR9RvUrAOZs15wL4AqmQYZFcL86dBXSYRpuqYBOOYzAyILu/KDSiCarjijm
ot1mNHNAsS/2XvULEYc1pfUsORekOOikRqtPigYbPgbSJMeszH8Zt9Uu1z+I5ebglaXVIqAOyFHg
3aXer8Yog9gUw098P4kawawtHkgS1zbxUIAoeEfBqiKsLX3JEnexTDavjVi9sbdBC+6Z7xRGMj2v
h89/4zV6bd51uCmAOQzU/l3E2Nl77WQz9cPVjOwffs23gcbRJqyT3DEWf8uvl2iLXqNS1bTBbcmQ
jOA1U4Sex9H7/tmZmCWZGTJJN/c6PA+3/E9cBU0Zv01h6+XGv4uRnaxUHoZNPEXq4jyRCE0IERSx
r11ZA73+WtML0Z1+Hzig6prCgG9x7yzSu1z6sFb99EiUbN7Vzfh08433Zf1iu9RsMizSrsLsrPyo
q8afdvufp8DyuglOiqnlLmKUCRYihM7v84GysInPoa3Cv++ursoVvtzKTCDZyG+5Sfjg0Eo8632A
bNCNmk99lnyP0ehqaZbp+YozgeGSHMfmGrZR7gJIq7MuSXG7nv5J4v9fNTTOvLRD2BpFx9cxexHJ
adlCSwZWxm1aW9PvnSYxtgfhG8O/0WLeZNSe28JCOofAK8jzZW5Y3tD5XGTQKoT/08YGvX2jHyaI
8mc7Wd2AQhpB/ixu64cx0WxzKKdEzwfZJb/i95/0wUp+xpBRA0hJuBfvAEWgLcxtcLo7N3Nun8/z
vkM+oLjXVw2nY4J0tSuLAIYxahc8RWMa6sjVNIIK4QWc3Hocs3izsMlIw9yiiYrspw1sN59dsE1U
NN+XtXpb8PH9pMjrLR8VGNIRv0W388xN0dRhmTBxTrDuT/veoBXxFilsLCP2R29SCH5/drTf+dog
Ueh3woPoVPDVaiYJPePGoJErPkPpZajFxUMG7bUZk7Q9umxcnbZ4YwSprnN1u8nwy2N7I9ExtLSV
mH8E2eovlCQsrFyC2pcTj+Uqr6AGuIpiMmERxoo6UzP4MZiPqEPHEF17lEmmCokumj3si8ohwQ1h
5hZNu3Rbq0xxABvvzqOBPR/FvczMNIE1OCT8x0YNimcS0SCFKpKDysXkEs12WQOX4xnJeLat7x5G
M6byIpPYE0edFWvoPNlM50Rg5qFBClwhG8uz4iEjNUTTZqhuNAJ9mGxllcKYaMeSAqPXsd2KIsMi
GHjneK3Jal5I1y3d2500g8jCtaDa7G4vFiR6lAPcOPKtvqq+HN5eM0knXpaWh+uTpovTlE1MTefF
uCi5MRrKhSbinpXDtFfas8MvHZww4+wDENRjKkfS1gFgGAReW9fbTb25A1aTDY/iDbD67/tRjYES
2HC5mxeHwVr29bTD8+wsuEf/pzcKBIV4ktHK57eoxK30r6yuMqT6H2WUtnwYLLvJZvNwUkNtHre0
i5ikVmITo+LDqYqp9B7GK5hCcYu3FvB2EP/I9TrVSGoJGQXzYI20rJnvxeCeNAGgW8GRDXcnbnd0
+osJx9h0JyMMDxiaDLmv5InCy8KPv8Re8PzUE1bAkdg0c1lL9YCdHw693kb/TY1BtUUtwBrBHROs
cqHu/JOv88dhUFCpfQw9xdMqBlmQhEt9gyWsI7NTIMn/nj96UD18M/AkL+mA9fVuDa2bX9W9mBTa
v9oTZGrwotPtBEfBbmfeFgmzsz4bITIkZI/9wDhGYPNwrY99l9eIQg6noAem2F7Ru7fEr4x3ExfH
WQQkLQ8iH35/0WF2DUSxNaZ2h3f+xNTDaf3PxH+HvLLmZgicaYxXlt0Q2EEaK/A/pLImO4UWNhGq
E4qvySa3sIf+9pRLBOwgNIFydPs/F2TJN7P/KZTRxIzFn07CnseuE7Pip9gJXwBVZ6NIvcwMdbsQ
VZ9HR+KNlqX76hieNVvKzpuCTSSXiE10GAy5b0dKPAu2g5cuh27bW4f2HJiJNBFdLaoiFTkWlTYG
RXBo3E/FqUFXawFjfjugbF7783r8GhqMtdHvvhhCyA0S+cyYLiQXkwj/dT9inuCpKztumYjX6P3g
qVCcNile/582IixJdGEqearraHDB+I/Avwx6XuqYAHwUTPPfYvY6pVDOybONBsW7S6LrWvFZZFT/
sr+npfP7fAttvVOmdwNYwVD+Bdsn19hDP0S4ew1eHY7iGYgEoQOtVwhbt6RoEKg3HlRjGN2bCHbg
7TXX3HtS5+qCvQGdhUENzDHLdlLy+VavPMS21NE5UYvdk2/bCOXC1Naj6VgFh3A1kzt+EoQgCmqK
UrCXIR//JhD98TPRiEwZZunSRKRGauu0sUfmyfILYqWbRZuEAKYrF977k9jCJ5Uo94GUzk5IhGbe
Kddc96fM+v+07WBTF99OCvPqT/ddpSdnbNoba7tlureRIFV1m4R0tnodsJyw/Hs5vvQ+6SU4psuv
wFGwk8WDFGy5Z1BIQQiKobeJqg0J2jhaIFYuSDoCwSLfoE45Dg/vgAR5ykHKWS2fm5M9hnKC7qOq
ZL7XSeyMjaGf1fmEx0vXmi9TyJukyoNA1fOybiwb7rCm5Hiraamv3p6lrUr/Ic9IZP4FTa9QQUGX
qE7e8OAmchz2w/2xquNxg8G6iBQzpgA0n9J97ZpodmH1xHk9ikYsTqYakcf1T0rErwNlxg5cR8Vz
6/RkjeijgSOlUYzd0dEmGsj2WCG7PUlY6FxTWKHd5aNtRs1cQSXIDXyTQKiQ62gxdA73ZSUiePp0
AwcJJkg0ibDdmgnytkQ0dZO86PsKZNTX2qI/1rC48VKFNvA5lgwPzEgI/Bs7d5VrIWCmouHZzINk
z+VARMCUr/rUxN4uhvIqQJUgNXADx9ECqcnVjiEqyil4NO4tHSdl8y6LVT394QCcIJlvX1MZeWL8
2zqT+A7vQdrs+dWiYAv8sAks1BfxZxG+wnXiUG8NNICm6mSthEIm181z89erPJrOTnomZczt7MkL
UE4TuBbJiBE7nNmJM08Vfjdp/cu76xlOzIb/wuTJFsF+EE1e3P3K7Ra16z2gotqC4UOiQUO2p8ac
VJGpLs0w2HgC5/9npATH2oxuji4EP9mOMjmucQJOYofOAAU5y5fGa1zSVIG/PrMRVcpzWnAw4qvm
X9as+nfqCVivj1UbbKsKw3sBt2Mv3j+4O7XdKA/uw/txYvxQWbNvzNRrov4SS/0ZZpxn6Rh6xeUJ
20eP46epUds8eaQkl++6s9+RlmAORjTNzfA7eN4YYjphPuiphMExYIZg+/rkwTuGIC9AJCHQVvs+
6aaBfYcnDdNoVzAmd5f9BRitngkOFUv7fLDD0lhQUhbCKAaAzLxu0hH625HtJ1bFC81u5zh+cjsN
rp23CDocCPuHPXBGgL1rtY8J1+EGpRxO65aQKityT0Tf2p9C5Q3D9DlsgdDciGkDKyRxQKq/MmJ5
v1CTz/TOjbBPF5/IHSNWKs/eyweJM+9lFTD8icwGBeG0VF51Pn7mcRCih3xjvScSdrkn7Ufk3vsc
GjMKWHBb4YvjovzzJVLzZIUH25oera7Isg/Kp5IONtOKlMI2H6olUElD2IZpGkBj4caiTMz+29z0
UMK9/kNubZSMoBOWQhJ5E0YIBiWVVuUv5VE5cK6fsfK4nvIuG5uCkecJMalzpn/RYE0gW0ogLtCQ
nkSECSRYJkNI3CUQcA9yHJDtNMGDw+xvtsDcxs4qGs+7CjjFNu3uXTwIU0ZawuGHY23DGTB4Ype8
n4+/HTpRkDD6vom+QrvLjpBqd3361iai7URyBLVCfZzrRiTAMW/i46LcLY8ycLmcUcxTl4IArHUe
EZENypbgfwVF3ysZ6HbgaMqRUSAi6GtS5njZBlbrf1nd0gsRNTnmReOYftGdvSs9KzKCnDBhIrYo
+MKH38hcV/dUkfNEPqI8Q5Ak0dTrt5p3u/W8hklpS84Safl+sdIeGGWzATs6pB2v5ju/1dXrfMte
rGOh2Po6AffbIj6BEO0DJ/bRDQsMyZNrmL6aws16mZ9bhI90eiJ8+h5ZjsRaJXQrivUNSE0gIsHJ
alEhLCCckNSVmNMswAka1ADnTePQGjAiBiIgoIlxN8SXAhPhcUNXDP5CWCj8qxXDU6VTlhda0xES
v5g1Dz1mjl2R4INkpzS16LUiF7KG79BUM6S5V5BDXU8BjrlXjt5hRH20QsiwFPcUk+/d++7ugAwa
gUdYvA7Z7f9zAfaPSuWM8StY/icY1S3EDJn067TKwJJCHpAFU5GBtRsqiURY3GOgk8Dzd3NH7ARn
FS4otpTjqL0wgNrPOIBD+l/H6KL+ipb19cEuWOxX5S9Fi7lNAUgq/jnvv1kKU0Lyxo496Ud+xnfX
iWxVv3k6es8i4wr4k/AwFZlKQHF2Tcwc2g5DmVBG4ZsoGUF/92tAxj2NDK2JYN+pMJprPdUJn2MP
LhIapH2uMtpUngtFgBKmJK+6bd7uwqlAlr2FBiOy9vWxkOlbuInEwL91TngJapLZat/3XSoqcbVB
62yYS6VLiwYIU7K8R32XPGtoZY4/6VutSX2z92vRnXrazoy6DLC7qXPmQpblQmuWz7X+cgIRynAz
8LMNDGEos6evPAIQw1sl2k5VdVenpVd3r9Mldv1lKTCG8j4Pl/E3hH3WQUW4ilY+hyVX2F4b6cYj
ThZ4hBIHMEZAzuplU1WT3I57u5J9VjcF0taw46X3mik/54xPWs1uQaSQgrRaWT32gdY+gRasWvMF
Grc1n93swV02gNZRjM1pxiZyfvfi8QQkZ05eS79menzuIBbW1z6TaaSuBIxRsoEkR2mh25IeujTw
AwKRXnNZ+c1H+LmlSbcQURRXfnduQ/rkSFMEYKQ0ZuYqOjm3xtUYw4TS11/+JbPl+92ID+EA7T4C
G3MSUOJrdRRgem31LwejAFj2pk+h6RlvtdPLu114TkbkjzxDC1VMPOg5OkqYccS1NYqQcN5fi1i8
iN/Wo02J8TsDAGc/SkoeQCxRWp86ZrVGwocCZMZ2sHa7A6d33dh0pMlbDZUXZOYs6HmMsc8Ie/AJ
lyWp4MKvOOirqPNN/ksSBsWSXZlMGqnu0QAU6s0Vkz6zPX/jdydY47I68rnt2aesVWPlzzLlWszg
TU2YOuEtf2zt+EUYE+qnNuixrtg1oLLMHd5bMEAlOntDV8i3RxNVtLBRW/xU14ts2eCMnW5r6Wqo
Y7KQLRetEHO2RZfw6FxfZpXBPAKps3qRd3NldGyxyVZgF4htzT7zcTV9LXHhlsMq1ADUhLzXkXj2
3w6l3tUphzBV48OafFuGnDu918PB/mj2QdCsiz2eJtetjcfkqd0FxAyFirUmpfMVt0sR55usjPV+
ZJGbqOlOX7ii3+PWjVrsZ2P2ZDTlncg5E3rKtNPZmbbe4Hj1oLTPicr1v+4jgAbDJCPry70LRmOZ
KPaLien4WC9L4042peqEIH3zKJat4n6V2a+YKhLikFLYxvMy9FnMMoXt+hgx0uVckDhhPL9gZGfn
bdrJmvSvq4IySJid14N/pce2wFsPv0mv2XfFArCVTF5nXhcXzeyp6cx8i7ts7LMFk5n3Y3EM4w0Z
WNz72FIEkc3ipFi2mmiIJUxv8t2Q/vdsdvvnrKBN/wyjdLInAn7p3kIvuEkPKlP9/KP52JSKj+2q
HUR8ieNbQrzVRLP1N05wUdsj5RG1JVNwqopdI2u8ALGB0FiR2CHdTb4p2ceeOaIxqmsnTSmuEio1
ahmdZobuKcgTQ5FY5GJH+nPxgXdaPvPS33Z6BNTXb7mPUujqf09VDSHMFfzLnRbIl6lbgwYkrM55
XiJcpBZfLwiTuiul+x5UOpEBUXcaFslF3KcggL7Jc4nXlzo/U8A+rGuZxclnLYfBOuDTvwdq+n7R
y0jxKUf6YBXYXoLOvrg4oc1w9zFhObepYu7zbLKe9vBjRcCVDeTJZ6pkn+Ipow8U34A48xBWZRHm
lLkDuFNBmUPnJhTYMb5sp5IfLT//J+j5ByNddk1O/PPqA+2oWhcYbwhBbdNaxeOYhe/7zFpQhjJS
0A5kIaFd2LiIRXT/+/2I8lVnoq9wpTAqdpJWSHd/5FPi7Ettp88YCyRlxGlX5AFDVhiVip5gq2/v
Gd6JwvLc3l7szyZS8vNJLl4mvZ8zTcsFK6yYZlnwLf0pQxndb45WuFnOcM+vQmGpjrv4xcboZjZC
lsBlFHibEPaO4I5AKHfLEquhbDcR3DUfrWQTwJK1e71l+uXCWlzCrktk27Jm064xHFnLywZ+rfG3
o/sjzL0C4jE0t+rrQreDETHp7J7s2FWELityIpLdbKqStWzylda5ayIPZEknaczEv/XeA00ERPEz
MnvvkzUhlXimyNKCE83lluGDYErPQuwGjzaThGfuoZEilSrq/kOLiDMbcspwJRLYkBugP01yWpaQ
BQOGPMltmznZO3F9r6vxijP7QLFtMBN4NxCKxMkWsmD2hd0jPz19k4eD5hMOQZGGJLUY178eNhCD
pyryyaEezkCq68TntDQpQkDzKk8NzQTiXwW5uofPls4eq8D5QrVrbVy+5hivLXJD72RAuxrEw4vM
zvA7o4/PydusMtLKEFL/3kuxVzD3JxHT6jfptzmm+fNlLMKz/ZMMW2scq2w9Mid1Mb/5fbmxXEn8
1IBByjSldZuWJV+77jBD3HVzrabqSGnPyN+aoiT9VykIMNqSDTCUcXn7QejNURTo3HrmOU3GeC4c
uFsejacCN9oEpzE8uMK2J5Whlz6gU/LqeM/Li5Udh2YvjvLITQGlGsB+P6950FmJtqREkic7KSjT
1QIQt0fsj14lsCUMDv4VC/aeBe93CHlROx4sDZRhjDulUwydyWrhrqZHQZ6zGx+D5hs9BVx4FBQD
15evP8y0EtvF5iQfsDlttAdVOLRfJ8OIAo/w31Cchi3FNaB5RmLJ2P6we0lvqtpIkeOSRn1VfPDL
eICuJZXFe8c/oMM/RngcFNoBLJ/X2KQJK9grbQMyEpMsp8OmisI+8ZdCD1P46u8vEf8aTDE5/y+z
ZYKkOhVOKsZN1RYcj6baScOcF0Pab8ST+9FRvmqet1vn66aEXuvD61d2bJK1PrWjBb2wJhFOC40B
C1/3lU2yiN13E8bH5hAuv9OMs4sb/10+74/tIwnlQDhjXbU3yacvHoLwWsKccfM775vNA802sj63
qeHLS2npywwhyqQT3vCAE65QfuwNu3z00mvKBs2MHuPD+qpAz8+OnM9B+yB/c4vVoPPeZK4VTyGW
+ih+ScyW8LTrjVUJErXe33ZL5JGQz4brX4uLdOfP0+DgqCyrbpKxnml9k1fEHerMlvZNSi46Xx1S
wcfsttIjFArJ3XXteR1LFWLDy8vtl1H0v8ez3elbJ2iFmWGrwH4fw94itU5qdHyTA9rzRACcsMUF
ZsAGN2YhH9gxf0GrFIb8pD6Hc0Qiu9qmHhXipIuhBrNUHXM5OG0/NKPj5wTskTqPVwfeX6A5mRrs
y+1pHnWSpnmDsj+SLefccNxHi2MUsxpzDpLBzm2LqF9iK8sgnE44/7be+w/ZfMvGqMnt45wueFJ9
oDtPC7/d027l7qHaAUZEZ+pR2ilk/iGJhHjK2tvoMKElAEwTdBOgw279xtIOO7gRRDQTNsb3bHmo
yke6eXTMag15sIX+Gf/ZTE7QehdCHVNznx6ja0CkB0idwObY8TLOc/ctL7f17CVl6Dsif9InLi7Q
L8P/RaKbGGOZ0EzlWp8QbNgNLDHOm8kBxpE1as7eP9za2OEfQqE62nc2zkdVWDNrMu6UhzyXiVAy
KkZ5qCKx2Ssa9GcKiuGWf1by84xw5pPvEpLPZK1sMdzo3Yq+i/MhxwL54OoacwERaSHWKxHLU2Pd
SiU3Ftxlr3uktcEGHqp8ez2T4JAWu/y7Vk7WRgN0sLJG/m0tHT+ODr45Y4Ua/A4yvWiffqaKoM2i
Ug3up0DlVpuAbk9PRgUXhnU7x0dWyfT0L8Dyq/xd7C2XrCNk6CKziWe6/KqNc5g21SQ3FLOX+aao
hWR3Gx04emHobyEMCRp5U68Rk/7PQ/8+KLD21x1gCKp0UF33sB12U5BaCeMS23sRtjkywqMy64yu
vKJ2KQ3Vy2XTQaMt5Y0EXP7GrI51LJGJs4Y3WfJKBuxJIg+AYnRxZeBl3KT74vuXvUSC569z8l0Q
S2QwPjk1ov7GBNe3rSLKQheAT2ni6Vde+2sPs2Qve1+oAGmWEbPfi+i3DGTRTurEWMxm8a3zb6w0
KUeqf+UuBP/AESEwdQIoIx5UZNgtA5wEcPgDhyDoq7htbrKkCXusbMSx04PnjcnNi59CGbDBUmDS
w042rAzOnqiwjq2GYjV4qBvnDYaLsJW2BFO6AC+KAs9/rYNyQGeZ+5ffMzSBwnMfwoEYh/GUEryb
V2XQq2Be7prQjnArZr9EwRpCBGLCUD/Ol+5VCbr4cHRA5aa27zIWkZbLTkHTMDF6Wy67yuB8o8IT
gRRWzI8H48OLFOC8DS6yRIrg4Ax1bDC6dlzNGB0fnSVocQFzopEzG6jFCLQ0gB6l8FH1VsuTKPvC
JZvV9Dk7/zEUzEWhGx3AMU6KTWNXVcAQQOA2AdW963eIhW80SWMh9xVKUtMn8uI0vx4D+OFCHhxo
/r2TBAfB2/z1fhx9qbZF8J+KsSASTkjOtjGAloV5WbX5JSMSsoNEoQRItYgfdvuDLSVbTtVh9XR0
aw0CHqY5tLgmCsh/oFva5sXGXWLnwZLpyzuxCsuGaRrhSzPqWDdeUmWhtFHmyiyRoxqfi6Es3UOw
MCGUzyqLPZNu0TgK7/x1uR3vY3EPXVn4uILpH9qXYxhSJohoSqG2UvaXMBtTpLKrQRppHo7ithB5
PbUEx684bG3N7TGUYg29XjaFoJRJhMc3jVYJq/KCRFAuNRye4V2o/1+ZIGB0Z2/KaxUbLIl/PuAf
yxRqS45VPn0NaDhrRV/OnxhsRDwFGRBka0AH2pUS0gdM+2D0VKiNAxnrqZRyjqMzzcPbitp8/6ek
v9L5LJwXcLN8lZqSY3VBnZypP5rtcrrr6AVX3cr7jfu2paNwU2PQQtN8KqwvE508Yf5yTRMT/Pwq
ZaKQWxfLs+yGm+F5FwX7h4j1elkYp8MjF/aXWLNffEAhw1JWA8Y6i6/hzZeXrDUfsb3/7CRGAVtL
EQtB6/TXc8r0mIOQmfTeIFGYKSeUTGR57fqkzHgD+blNojr5xPF2VYtbdL5+3c1dqEpfmUZ5y2qn
DdCSsLBsYvVxtllRf4zQH5QrZZAl74RpZvrGeRCqVM2QEL9l/VO565EsAuWMNinW0Duxh123p0g+
cmUP3IfdcxDFBdSkMaPIhNwlqJJvDNL6K9aTy7lCSp6HEH/Wcafif29wHg0AcuhmzZOhCrG2WEFS
3wFdoZZiy9W+0DBiNgagEy4lJzEIh+KsN4A3XEYUfBZdwuxLP7BmYQK/aNFfpn108WIwyzhtGq3+
iVqzYorPpAqrOQ+gFxs1hYRxDsHXpddYokuuvoxyYTtmN5FurMpr4NVvncM+BZE/0pbGdkZCoC0a
WUeGVelcHAt1/tJXwft5xoxleLsI/tu5YuNL9nZ5qsXH6Rwr6omXkg4eQptXIJvSDJS0ofRNk8kO
HdxECtTFgi7kQtP7Mjs4mOjMacAp7rrmBRdt9vQxvQHjZH89RNMD+iHD7PoaaeZpyYBQ2qDYF8c6
7lIv2B91xwOaMdmzgKgSjstrt4EycviWEGN4vteybrbSOZGpY0dX34yB6XI6rEZDloosQ/H3ss/N
yDw9ey2zLrGk9B3ZtkOB/MS6pSPNG21y+GsHvTO49RlNISCL/420Cmd1XK3DdKgNt35l9qKrSN+Q
U3nTJJwtQeo6I+gTzwM1BgQ2C8ZdMLkdWOGSIaeBjUryek8IB/xiHc1/R9EX4oxt814/r5vMPYyw
XQQ9XwyeWkxmLGzwc0DD+aKdjCPsV9wRXM38SpoNGaJGPEI8NguoLva2W58VxqaCHR5icWaQUiPX
YgUutg0y6nbbKqth7pUTSb+yY37lELBdO0NBnUS9OePE8tUmtCLH0tha950DxdoLc6Qbiu0yjVJm
C+79jbN/0eLupwnOtR7Pms1HFWrvVt7soaCC+wBtn3IfqJy3FBYiIbUZKLM9yBV8DJjyU0+utL3J
UrQgVsHFHN0eN5yl0whI/4Pjm53Ec/fECOX98GFp8fOE4TzbZW3Og/7G8fZFwKQ/Yh480seUkww5
ch1Q5PK/LgY2gynwOxvKpbDe6kKSMuRo+i4TILI3El56ME9z2W55rre3uf5Ub2rx35hgvSbxPpt1
CTVbI833VdvQm4qtWgoIaGAjCC3LId6w2Md7IUQMGmcvJ/gVE7oIJXAPC4eMfjvLttEpWL9MfdDw
v8fHAa8YauH9ZMXPQdI8IeeYQQSBLQMQvW2fOs+qC9fvnmXW3WiEL/M0vgoILm7a2h+joDPFVk1n
eBwgHeZEThS9KFXVIduSu1hm4YXKU9J0sY/WMCmN4M63m2sQ8zthjFlikauMYtnx7OfBvWYTL/sI
gMezCiSIRD0l6EDe4b1pUmyTvSGQPCnBLv9RhQrkSm0perDTx0doP7j+3uRusFVLR5bxUyqI5K+/
mvOT2YPddJSIDwtYeg9mzgaBqG82qehK+T7nn/Ue0zp3Z86lJqMvaoKlmya+G06A590bPIp6ocNz
CoIdiL2GU2g82Blpn9Diy2kMvMXEEIXYYjO5tAxccFZDKH6VBLJRixBds+eD4XeHN3JzO0qerqG4
CC10ZwNbp65OQs/vVM0ucnXmtiHXqvBj77OE/n/+yw0PFve6fVmty10zfWnqBRZJmIqJX8aJMzmw
0/ExSkHCC1FCw6FGrR1AWkMm8p3Ln2BhbNiEJoW3W3hNMRzcCFNNDDtzO8V9Tmo4N7WBocuNrZ48
zhQ+k+38VbrobX5MLtveteWjCx8lX3/rZr4RTXdokmDAgsJWPp9ne8pnCHZ0GLhVvSwR2bwpHyNJ
wU6T+82VpPNtRrIqGq1lF17rycpHrXxzsudGUtqGx/fYVwGGwO/4j40pbG+YgxceBWCJahrfFvDf
iW/m+uKy6CWcoEfY2IBf3vrB9/S/zppGCnc/P9GEK3bEL4Cyr4QgFcu9JoTi803Arz9OROrCsgyy
Xoqefh/v83WpOaOOdK9/++x3nk3Y55lgAuY2slGb5Pst3ZHx73NovTMHC7075GStmp6QA+JJFMp8
xiqL2DYeeE5uwl3PqwxSIRZxWM7efdOVmjyj4p30g4MjvcEFjPlkDDXIaXrdAnt5E9z2+BZaQABl
/Pfk998yFnMiSvjrSZPf3QGpbePugJPZrS8XF5v+K2TmH+NRb9XEsmdtXvhStE5knu11Jnv0ah4w
FjAq6jAn9P5/yl4zRNQOcOpm4MosDcYa2PQbRRvZdlXW4ap2SHaCt/BgEHnB63pvF3pc1mXVe4F7
569Rp+TrF9eexlcMsj9ssKud63AU3BGLhz4GmGP1JCpSxvDWHfCI75m47EHA7npnmHeRFEPEFCmt
MMuqNYEU3BISNHjZZ8KyHJ4GO5CFyNne+L/MPIpju0ZZepPTuAoBpBBxZijYX9mp8DDR9tad7wo3
icMGZAOKwQtHb3PligTpIDBZS2pb8jDbnT3+teZbsrclFvSAr4DcFNtrovFLPasn4b70e4MzLoXM
ER+vlJBJzEsjghDCW0aK+ZRoZ1dK06AdPTjwLHX/z6AliwL/JbMBxhtDn4UD33NSZU6tMsqLPbB5
8/A+m+N31fygqQgWTdSoZazQJ2+05pEL0cx3PHloFdBFAV2hJDEoxHIQkvjmZqvqUd780AI6OeP1
8L0X2qMl1xarhDdArO6G98HB6+5X5kyzEv8J/RiYc6ceHWYmOoPWk3ay9cXfxi3qBjCC4gZsY9Ky
VMiTMGOiL5Zh6dijZ/p5Ds4qUamDjlGPcOnjdQZz0mgogA9GJNDrY9kGmb/YaP+eC2OnhObpXqiu
Jc4vc/r870utj1XHz7ixB8Se9vUTbs/pV83t8ymiVUfbS7l39xDaF2YdfGkAi8L7SaG16GtzjtIQ
rpMoPpNtVu/KHFYcVQAoNVXhaWWwadfJGwvOqrdJSWpcOP9mm3sUCvX2tuKIlDcUzLzu5qnhG4cv
Aq2lL7TqBQgMEclkFacXZMtnbwMXXKAubPXowx1ySXOZ9svGDfpZ0PX4TTwqPtaiR/skX5AzDwpM
vQY6oa9Ebi355pkiUrpP0shkkSjlDX+4LT4vzSOUrb8cSjjeR+m4sDtq78v9BME0oEF/046MVOQU
hIRT+89dTZz9J1eUWFXWKF4zVnFed9Msy6lDROoNHqbt2+aroeeViMcZ73ryl9zs7b6CQdISdhv8
KzB/cxTzgxzWKTm9G5Hq+YI2SrpeCZlSJlIx2S1KA2fkxpoMQHStSwOezDdWWmR4alQ/EzlT6klR
PdZpN+mixJFsr5t2/IYxJvz09/xtn1BmDP1CXA5hzZKG84ik+FJFgN8yKOwwPZ6ll4fA6wAdBICq
LPfCSIHf0e4F92EzCoq4pdt8Z/wULdR+lyuP56S6NQAYXF189Isp7W+eEE9MK5DMiZFm/nud8YVN
0yVo1D/CT65lpzYk1CnHJUc/phm8ER4f703N0aqx+Q+s0DQqPsZhsYyOdFkMz21ku33ki12RNbF7
YcrUjXtHyBJ+HND5rXRNzl02FE5J1X3UFe6qpinnis0XS31tHZGXVrfmQoeKy2K5wWT3YF87NtET
x1aaMu8H6uT4/clisFyN8vmco2b+Xgplt5jIu3hIK0xIsVxlcwToG2LccNsEt5o7PIzeQQu95Enm
YDHxEqLZuNlzrgTHuCzAWbFxKkSsI6TCTGBSPXIeLJNW7X+a9R3NA7XuyahQB+oxI+bXJKLKXdT4
6h2YVVSuA5QGy+6JSVBUSB0gsCi9BIJNSVpOfGWn9x+BGtbcXTXJ1KDeSZkDp1JpKAhNYfWf+eMy
F+0/QMEpIOQFNMbmqttU2HfCebQWz3iXm/YgmVPNaE46U9nCo/FnB0adf48hg3Dd4BSir+31Ycs1
12buzhEaH5m9sHHK8vHRxKKEztRI36+jqdUaaBTgaXYL95Rh1YzwnHAZehTWa5hmu1hjw54XLjhO
fs8CzdQPabesWq20wxX+ZCo9upPF7Y028spOv5EbFbYP3gM6nkhpcz+zjXQigxGgSllR3upIEzEN
mT15li6v7cXOZWxLCs/kOGZHFB0ROOXOv4IXRyFeQyZb12igInCnKsEyDzV9H/RvRbCwhw3CIZXY
Acm2vIaL9nk0h+CmEc5y7bl43D1aytTxr2BXwkYqe6iNYFAMXhIXwvKIfCwRHDNWD9K0aM7XWyO/
7N3Ue/lz0w7XOzeVAqxvfNfVPF8A4y83IJ1riyP21ZbLEw+74K38rrjdblyFAoH5I77yatbE4f2B
0z+MnlTJwsaRsewkO5H7JrwpmGbJtZBP+lQq+rC9AyBOuwJGfNbe2sIs4xlgygvGhVi7H5zZ2eFU
GaQbxoILcgCKsgpfLW07whN9C104YGCnPW7nfWFpBotfkn8qV44iJWcYB1i6Y1SX+ZVRZIN5Jo55
vwPdMDEkarh1ubw7/fMJ0RolcLfY5lNmAQLkVRM0kxJbXhKivwvYCWmlYjPAxa3aDztQVWuPaFAZ
tKzPioHlv6uAtnWfFt75ty+zcatomQiwWRyUtltWfeMgVNUN0vt5SA8g/MFq/kLSPzH12gn8xyOH
57vqK1zk2P6ffamdRAulYnUxdlI9NLn+8zb3pg3FMFQP0RQ+4zUQjnXZTtkUVpsKWu0Zf5pPIdaJ
Axda+PR3yDrX65jv0ouGqdFyD9kfvcIHufSM/9eiEqZRlpFxl/bIDUbqDHdHfukM3nldIT4JCoKN
dRe+3KpFP6bCewYG6krmGmdAZAyGD671GunUav1e2mefTjDo1t4s8sQdbLsaGhVHNTOsCnODkFwY
0VzCxQL6ovkhH1WGGso+rBapB40xzkYwRTjBnPb8yFd4MKU2hvw/SaBP53fPOsPA0K1fYHpvU9TB
6taWuROz2hCbCj1S6Uiajds/RrTqc2TQ75EHIehrG9vdGkW2OS0kwNWKxglzf6DnUllM+tnnGna7
aYzQVE7CdqBsNxrFAoeYBjawAH3f8eO+3JdXm2tIsKLD5tgXt1wyDHkYhSAj4hyo+VaHZ1AUuR+B
3u85Tog2KxjkdnBk2GFvH10lAh2w7wHyVo+Ana3bpj99mgXU62bjNttWA0acFjnm7ATyEIAINAKc
xQe0YHUe/822WRYql9Zz6ZHi3TYkqwUGZ7XtJajdxZP1HPbxCWnFmDxHO7r1h+A8r8ehTUwOf0f/
g0wFTibsN+97Y3Tdaif71aG6jKbR0U96uvU/SxTE7L0IP2JO+lcAdyxMvDvHz56FuUbwVmurzeza
gtxfwyInstR85aLk3VTyxZwz7daOze1zlMF3SWBjeJqITLbXpEqBX9fWTUDctEgvZYLImKCa0vbV
g3D/3vZJjjZ0CcS7GZTeVoeNu51g9qHE4kSQARH4e5hg62IOFcayK4xCbVWNoApGHEKPvFOzPjhQ
Ea/oz95bElj0MFM1YHEKL/qrNqZSmtnJXhC25NC/PfXw/Q7PpqaI9huVJ+ekdYdPVzMyVEhRyxp0
P12c6fAtO40XKmJjyoyq9KjUsBn7WC6LiovXTEkTpdG3do2EPc4OVMeQ6M4ElcpuZhjHngiT+ZW8
Pf0E/qO00YY/Hbo9UsI8gBEvsZe4DKA+rzSi4wuF4aRxUqCJ0krnrpvFMkh7xgJt54QlQUpB5KI4
OVpd168eTrlA9GXOPpHVnNsMWV18cOTkN+zTi1v1YGK7hfQUuX+cO1z3XWUN3w7vlF5JYevss9Z8
XbFnVIzWh2PBFHeSrfIhCa2w2X7+6bLksXdPJ/2feYJ0XJ5vZrtq7RPdHFxTcrRV7JU0cKQ9vqkP
yOJ9S1UMe2/NpZpZFEzdTCLVm9tKv8tcD7uN35R92+PPDf/DSJ4AeFGldymMWGLrPVl6MzSY+NsH
ZJ4VxKTuP7e7e8Bs2HYP/u4aURBeU4BVd9EUNHcWiTFWJrqfqecVBWFroS8BiqPRbjSni6DTkbWz
VzwYeVVaWhT7DLQfjEVrBsV62+lWdhSL9uLPY+HMZ2smA0RdkJYM4WiU0onq39Mt5DAQUqmC7tYm
pUdhllxeAtLsCFFFSnYFJcsJT5GpvGeZz2OVXfbtzGQAynxf6u7X0ktxXMvE7Hed9394OGnoZoJY
MVNoIgvoqKw34GmYRIHk7/aWi8CboHKYw0QwWEzVHOOGfYpx2sJGZZaQHT+io8ZDC6gI3NcmliJR
mTTPmbxKT0lz9TA/C1wDjyuI21j9F01wwyk+xQBhnCjFXW2sPFgL5Fwb/bwgQSqD+LSqpxRUVIv5
jze4K5jq/5zi3JS+Po6xnIy5Q4Co9xe8mpnhWe6Z/nx0Y7io/1WZnf3wiXgMJzS+iCVsZQYfTlQA
8ZAm3R08PsypOoc6r2QED/yOomUI3v/oYrwXMpxBb3G0UXxwY9uI+fIiPbJxsdw6yRmCWLT8QO/7
k+tsJdPx3xI8NW/a82CiuUgwy6wmjdkc15c3Zzy3es+KjaMxn3mBsA8BQrMDFn01n56QBYdFgC/J
EASzeoSTcO/3NpsLWM4HSTP/JGR1qVuQUibeV5kYZnPtnqt4Jlpo/PaKnBHeeoUP0knAmROs6esk
DlypZakmxz/KV3vHDGsLDf/o1MVlx7b3aN7uFkne7NKeA8pSqhxGgsCGYASsIRWBgB3szwH2oAoE
HSaP4IOUeMJEoE9Ypgts2I07ckK7JqK7pBqdTUK2krP4v4WBjAxYzHeJNXKb0CWlrWk8WBumDD5+
IIqC76+bFIFeW0kSP20zJ+e/VbkZhdnJfa4F0u2Bk5VWUdCyP9O/qf25ekh5zFj+y2xOEB1OIRXk
+iUMbKR4gdkgmW4uL+8UNCoUSLDYGf6dzZ4udoV4Zj8uloffRCNxe3XerWNE1uwSgQxlbEfMpGYY
fNyUcJCQJ6D70omYzdHyDszDS76hM1B1sEaLLKGX69vYTrqHg5f8leDs1l+WGlHbdwpCZfcIfPJL
LfsCLMhGY2NOAt0/bOUVUvdqsanv3lsj2Bk4RmcxOCtFeGLvK+AgnE/BXNuKlBWJGbRsFAcDuq2h
yC5vyDWLdoZghAmC1a+A/FyAklOv5gGAE7IF+AGh1oSSiH+kzqWVAKqzJoE4WNOQyEzIQA6ocK7C
kD636wVqN8SyoHiLOb3XouRvlAuFeOKCcpIojGyiyPbMfjKuCZNRJ3k6Fr6XBYWh7ZG+uv/nmBRR
S4bmppTlUF8/bppYul3wZTcGD7SAZTUGAuxX2zVvThY2A+VBav+tu/4OY6osYqrz1OaACeg/ge3T
zPSo1jEACxH2faMBTN4E5+ChYNQ+cc26vll+OG2AuoaIYzoYL5LBb1/HOb5RCA/y0BvGq2DDAyUj
NdxfooeiuaYIsJ6lhl61DEefFRXtf3RYwD9fM67H+1NsRPcEvqxBOI2ohGycsHg6Y/fsVQtQOIMg
avrx3t7dFW1axU+YlMnJFO2f2JphECS+PIx3meQdvjbydWWQS3p4OysZqNXoJsdmkthOfZPFqnCY
XLFU/eNVATAyBiiu6tTLLTOOP+/W52hlEi4dX6SNb/zT/+11+euNrqvcQmDfkQmdv2JcC0f7BOvh
z0uCW/PRMnwNa0SztMrVbqH/1PfZB4FWAQphwB03pqTkyQOxe0P8wZVlKKgOP4Ni64kCWLWIBbOD
utVxlE/CaFGUiFM7KDP3D/tHU7sHLq5UPJn4TT6jX/KXImxGkjpXNPotn4Uwy1h6mEEVVnVb7cGP
W3nGdXOnGVqZDN6wHavFKPtns1JuskkepqlqRqCMhmVi9Do1MJjGkkqn2ArhEDHOR8n51T2z/SBh
Zo7inwN0I9t0+EPzA8E1Qx/Jxow+TbEtUJuz09Jp59DIiAGGYzxU5yMv4+H9WJamD0ua/G8YuYeR
pYKRdJhW38AtoxgPnj5bKQ2T8/H9EtyNBSnPzS6WSVyTYNUrEr5JnpxY89wHjB82ypELa9YqURJ9
/QhNZaTsulXhrpHj7T/YkYL+gtBzSTz5jAZR++LSn7znLFWwLItb02PbWnUfpqSPoChPqMZQsFGM
m6QWnI8MAItNFOUU43q7Nq129x/Uw4dVB8dwGrULxW5q4rxXYFAVscsHUkXGYO+M+JRsRLG1GlrM
zOc+RWlPl+wjpIJhPUNnrcuFeOleYNRCNOEHs1k0vDVWKaeBcsuTjUI28CSXARGEMC3uC7p+hvd+
2WFH5KfD7RvQUkgs4oGqGpjJzzI7cvytohw/lInkoYooTsPfTp4q7qVTzqd+NNAiANoKGauogQah
YyobeV+dmWTQWvD7NfD3G+UTU8jAOfnRj69bQesu/yQJ9H/iDU+WHZEKgsnWj83dRQFA/EMrbnt4
d8MDperE9UI2NmNaNN0VU00fFGLG00OtyODAl0teNCUtkCNQuMQ8wmvOVOBcqmKwOgERRYmlib//
w24yhsvzr0m6RpNTK/9fA3XsQRQqP//GZgjI1djl8HPeqESqmttzncTWhzGwCmMWBOiCghUUK95m
RnqmF0ys34y5S1aCGB09tchGIxgF63q3x6SKVWvZjaQp2vsYk/f7zuGqr+BDXhpW7UWCtvJTJXLU
bdo62qhQfnbYiVKkpREmIn8hgO4CuDbmRMcl8fyz2DBBC7OqPt1KPz2O9LP7wQ4bPfKvFEQ2gtUK
1KgRs45uE93P6arQDhWWrQ6+Rr/JWNJQXt10X5EGEd0T2YF0U7bN1OIZ4M9HJjjBC3TJVsvZyBNb
QDQCnS4Cg7RzmFpgix7OUHCm8AqsI9Ry7Oc5DW93icVD7zLUyA2dZgXhj8pajQ5oR5J2b4O4k1MO
1dAuvwHQQ0Yrd4h80xpJlAtPI2OwA4Pg5aOBqFOk8kC/trxZzjixsIl49DZKwS47t0PeQYRyd2Mc
nXPnGnR08IpYhZ/i5WW6LFPUuUD9APV0b61nFtJWZysWD7gN7ydMYLkPtTCkO3SlQ2Eu+73f5VYF
QjbKPK8DMyKgrS6+WdhKHbujhQkDkQWYNC/I8Gw7//Gsh8rn39dyk63xg3Vr1tLxygkFavytrc6Y
DDl4imayl/ATESZv+T9mfOYU53b/cnGTbcdumA3TKVmqDdfkaLTSuzlqxkuWH7JQ5E+4pj1n6M4U
CNleN/BMkGM3qlfpFKk0PNYIRF/0zakRQ5jLSCXxz+Len+tTl8zYwHK+5Ygzk2+SO3XIz5SpCC4X
8oPd1MoPJo2swVgqgTrDYMQYkKLw3clQG067eX0WVRP8eoHVCZdivV2dzRuVCNhizthJKhENrNnP
PzVLcPhuI/KV7a+3iuimND9nBh/jTmUw9EmAXfS0bhdVl3BUbTbr1Sjq6TILyhcjCiBlAAiSMLIj
W64tAQFmTdnuPS2df34a1NJvBfQCvIf6p0ORMrCE0in1lvB3JWIhFycpRvhPpznS4KRKUlAPZ/XI
Ga4zMT0PvHoakX6RlkjBl/q0nZkIQJAXovJGv8P8N6OChJNJr182BzGCYAuokBzIbBgdQHHL5zQv
m6479FzUBP57emFy+7N4zGSRmN2hhum12xUessX+YU7XbvRKGOiakMzhaf0DKRAvxY6PvQU3EewQ
hWE+LSYo3LVMme3hxp+4BAOKBazh2X6NQnI9PXMhmhNG/1l/rjs8LBI9k9DrI3NuHZUZvDA5rr8V
M8g0/gRUkLPQSS/Vwv76kGhXSj2n8GwaUH8URJbcABuguNUbWko9B9ED4BPlLDRITZm7wMYrElb+
zkwtamTvFldZ6whOpyxxe0Za9Uh2z7QF5Y50q+nXdNi7LLFOep5CnTaTuUGhCaxjI9u9ew//HP4s
SPygSpaC0D0VdQLW7nSKIFcAbQbkeN7IY2R65BEaPY9DwwMII3/lliYFHur4rjglJ5P/74V8TPfH
K/+a3HdOkRFcfFru3nhG8BiU08XT/CMSuq+avfWyOyTdQx2OR0/2zktYd/zyEcg+kTIwCiQ+b9mT
s4/ch63LH3BEUS+ki+mGQwpUyI6eQnMVeCpDR5bjZUiQRDYTOzhO6LLlekkrJjPwGgdbZYG48XUc
XS+hMqnxgfuEvfVpO5ARX7S1gdhRv/qmMTyv7Gf02puUhXio3p+YKKlg9yPWUnWpK8u/LYEzZXoK
hVWyi8QRQyZjCsJuvlnya8n5QVwWit+rdoPOBTpo0hN4M5iyrQ9xK7Rb0+1fUP5TGYbcuJ4kt3DP
3FBRohgYPc3PCApdM9oEHzqmxzoucH0446sVK6ZZqsS9SR47LnhcbOnvaKyowa7GYgXF9e52GRx7
o1jR7gI6r9OC1vGt75ugR2rb6aFFxADwsPNGJK+Xu6cGtfo0HmYu2PNDXvTm+DxnV+mf5LgYF4ve
ah4Cqwxrbr69ahTvwOut4ZGNOLS5W174ZEnV+JhGwAPEUbtdoN3S3PoJZFc0G/ZaBiFTw1gBR7Oe
hdRQcJMI5Px9PKwIL4Qf7pVB2jd+b6O6AfKBccq7rslLzQR9GPq14NxMtzDPe4l9SsggHyB/AKVe
p0+xrhxQPKtkdsgs2UD161EjrXCO4qlsPgzer78H4BTBRVsdv4SYDrRm/u8OPK9Mc3K6ADj4YUcY
U8l3HkKo26fCfzZ7DapHIX4tSbz6/0rSlDTeFbrs7Bcut3EzbuVBNzIDHz2M8F1zCPEq8WgPI6rL
5K9tZOMPP/fZ/j3F9jPxLtnqKikRURlsMaJJoPmQ9TNnGdb4b9g2EBl44KF5A8kVuor4n1Fuhitp
bHWbn2kqiRQbjEa5AzdYzOqWyqvPfinUQbl/WudaC+c2sg7WGDMD78Q0XuOZpydsY3Ih4l/pZ2tb
SlLWPq4VZqHovk+E1nQ7b/4HUcwfEBEJVijyzhLV2nYrBaaDeq4UdqGXdMfa0AUvjdufoI3bJ4hT
1pwjDbOLIYYlBxEpvw9c8RHRmoXJNT2cLBq9VK1zO3kHTv/FPa3pMK5zRmwBnODeYQWYWfSGGbnQ
SMC2ZXoE/r16xBjz+2+kpuSuuDADJm5Msvi92CxMP41aAjUV/d2ceysE+BsYtS8ey9DkS+nb51mc
veQOLKF5BfuCO4CpjaGdu9gTv4IVTnv7txdV60HSk4D1V8j+Fs2G8XAnCmrdnWBB1BEKJrWgEuAM
2Re0MECgwUTIUsbeFMJ5CIsJcnZHq7JNOZiigsGuZxQRRMNETTt0YKhNbjvlaQzpfkzzh21L1m8O
cJCMTJ+eJH26cgIq85jvfVKFrTaoFy1v76ysn5xuBYeZo2woirEKRMsHnR6o5+4huhFDecmMMh5/
hJMuj8ZM5h/VRLuUSLj1LyeGb0TGU0ORorQvGBcz1KnN/ZCS628kB5eMisyIuNSRxUJVfr2f3rU/
h/isR4tqkeFNtvMD+qQDlNb9ImX/H0gJc05AcZ2h+T2CFfLRY+iBAtMqWfUrzxxwtpQ1K0QW72PR
BdXsb4qa4DKsqNFVsG10OSRYbNzcTlzqEOQKaCPUXCdZFTmJeWJlwdVYAQPEJ/sKnJoLi1cA0P44
sKsNjMHBHmgSRMgk/J/U0m1WZMkI2j9OKoOGVQkhSy2gtDiWck5b/dValxY2uXKeCdrG/DngqFQm
Mc3mkuf7m+K8/rnWM5fBfftMFO/MQRJFHZuq534ENk9ROkc24K38rg9/dfsK54zYyRZVadoeSLZf
iXJ1hJKK1ZgcQaSlogMpKaY1dDOSkZlqtuaGCQOEcJ4KJkbpKK9GGMi1BWiXNE0JJqblIA+SHtrY
sIWugSyTyjuO9QJ/N8kta2sGMuzbfY2/njKbn+smgfFcNFpCYFWhPATXaIg4i7NUSQ3pJUCLgdab
2V+fHsmzdMfT8CfwX3RRTRfb+jtR/X0AH/V/k2eSA5ZoNLEiTzTn48xJzIH1OF/XxhYFWJMolrOO
8BoMKNfn1tBcRTN8uX5gG5BBO1XJWKWQjhZsassQyg3d15UfJh++Q4P/cSaQl+M8kX8vX2m2jI7i
rB0z/nj+/lCSf5rAZ9j3NxHCnsh57rBCWLw5N866v9CYIHUGxdtS6MVKuDo0vblcocqQK86qg+Tn
fLUMiSZWnF+GugvCt4MR5MvBYLivwGjIyPDwKsTtKVDsjJpqjTG2PvrBsddTdUPoRUE3rA1eMkVw
vzkxxbfWw2vyLJ2skMdx99w8CQO81Sw9YGGv0VziACdbI5GhSx90Kz6LlGfzgPGdhX3LGav848ix
ucbQe7dYlo87kSP7QBYi2Fp/sj71pxSHuRFvxvZrpu2O8bxy2QwD7zmdNdxBNNwlCR4Z240XOsbY
osj20L+mLlOGMOKu/BhIGSoqQo20ZdePqgBCmIpDbBHkKE+WMa+65RbColtE3ia6ls7w9/8Itv4r
PaWFUSxBylpAu9yTaPt1GFwKK6+baROsvfL75J23+Bqr8YUbqdLG3Da3pzZ0Ck63laeglzuuLK4J
NDnAdLBf99wAar7C1Evvc0IQcgjp9qwyuvO5MyJIzcphrQz4kwCkxdCQiB4xqktSaHAkjZcw0Kxn
juMi7eu1RaXDix06irhF+dpyOqsZUFfdxhFREB6nJTM+b1rPjT2GhVkT+pOTuA5OgTM71tDTf0IG
PA+hqzZEk10HNJDMNohIqjgPfDUbJ5Y3hNnQ4Hs/D7OrJ7w0lVSS0Glfwyhmng/E6VcgnLgOnHYi
37BTC1ADboNmCK+ywjMg+aKBHdGuIMOcekayB3XmkOOOhLMQZ57bH386QjnEB/3xDerGhFOY31M/
kTTSuOXs1T8u/zKyRUk+tK2kRSbM/kmAwet5d+wqeP1g+17aafo0Q0SiHJEVSaz+tUflCk7QZa43
Rr4oaD3TBilLxKMtO178uJPoY5fZsTE58FMxsnS7lc1PH3WRQ6NZEI8fBBz7+XtedkG4NPwwQeDA
MRLCMtwcmFKBsE20iWcQB0QXaymUaUNnMFmM+Q/B8Tav7ztBy3+IQRFFiXywq4yLUx5vDM3iO0oi
zAYq8Ef2IJu/IH77n9oZY/Xe8xLnZ3l5x9j2QH5YVpWVoxma9X0hvmis/P5YmNegOsLMGkW5/V+D
pzoifszSRTU+76Vw3qneRl2sVN7rQj7BVwjal67FJ7wrp5dhyK0ueGcBDjm9xQ2dQwzAknScJqV+
zIG5knHg9WE66xZRT0PO4jTOQqxl6A3/tnm5EMQqqZ3B/1i2sVnccVKtSnYERMypJzkVOYkBTUdg
h08AAuX4ITtHOvE8eUXDe/3gULaAKEz6/UNTfwy3yDURqvOumvjebLGq4p1G1vhTfjVY67K2pu+s
RmEUMY81/ZfxvRIITGODAGE5W+g47IW3NkvbEtnLDniWvdCmYO8AJBPITYM0Qkhd8ArNkPwwWWlj
8ra6fKE6vyXZqcVQPMW2yBcW90gRGhLTMoA5b7SMq7NOey5nXmusUbOkAD7YoYuPC6u5VlJUMwwp
yUMrMUnNBYY2uw0UluXTu9nQ3OatrZ06m/1bNatlJ4xQyEtYLAUN8h8IFVo9YXh9sxvSNSD0OJrJ
nxFtgxxHSlEwICKhoMEcc2JK/789YIsjUFpRcGOe2Yo61x6o9FgEUEk8ZUhtn9krQmMM3AhkvGXA
2+1HyyxSkf5sJI1i9Tx4+dVgGPZa8byD92zUq3obq78tuKBchvcfKCpK5FCmjnWg0U9MFca9w8X5
aPwcVYq2ihjr1+C96Dglh22kPxzy3jKE4+3KKNfCoaX+PQzziwQhU0eWKvXeOMx44zb8wtYGxDpm
32C01D1NCn5Tavh/A9amMSw+TicEe5kIHPBKMfYfMzmfhw/yE8VdwO2eAS04AGHh/uwP27axop1X
aEQLpQRhY4DnjH7sXNlBqyFq7/DwcmxkYl5xD1gnutdPBNP+ny1i0MSp8S/bZIRMQS6FRKPB/CqB
f0OC7Ufz7epEWpiSw56F2ub/rZWq2zs/JQQebWABcB6DpLtPTg1H4L1TRm/p/89vPSbrMNN6cgDO
n0jv4FtVEcZmVNuGh5WD2EP2lOYwAww14uTKPTC6FzQc/q18A9rjs5/NQ9aXOZ7Ddy1sIkskRvY9
nmJ8nPCs/MNea/wdyNAdrPLVDjbrEB9MZRcbCZl8T+fqO5NzM7y5WYyP82zbF4fx0EszMY8ZNN7/
T6+HBNHJLrWkg5DHl2mfYjsHSSWm0IYjTJ3KCyGXAdXsqIDE0YBQb1JBLJmFp8Be4UBKZT5e0KBA
4E6b8wg7kdBIP/pCqWvjWxnx0B4ndiQkFTI0GDY6dvLiP55kqYeFNYjFgaVMnfB6fhXbwO6QsB1L
kgMD8WG4DGLRgFoT4ZQDDxC0OPjLJ4vDZCkG+YY/lvmjRNy6sstLuSssnLc2BA2teA74OqOoIbvM
iMJ/U6FnWCCxs1Wl1htcm7wfZVdjNl4OtSLCZJamvrhKkQ+bastVG0bcDYHHfkowvrZfx7/55zt2
C6QdcqDwZdMnIXLWoWontEPKbMaVsgTbqlFxjdosKQUJZAmqv7iEE268eonuBFClNU8dWfj2ccl+
rpuxK+/RccHG4VEDs/rJzL36h4Pl8GLfVnkV+5PK5laubjZPRdP9YTXaUMK3H358A1x34LIzNFri
xVA7LnbIXiwdHFvl03ClwhQNzOg9Owx+b/70nMq0xH/j2Mhs0zvcekcS2wFeZfIfxU1ZgZtrGr+3
i7kKR74UBBMIomJMvKZNugoJeNJQhmvYRR0Cwq0rKGzc9AZnOfwPTuFUfRj8KLD8JwoX4uxpAV1w
Sn9vRSJGMw3w3j1eSb4yu1vrgEjHsGv5MpQ3NhtGSVYVT7X/zWO3e7PZ9t+BqTiaoDMcP7/UmB6Y
n1tGp2lyJi8/V4WfKODGfg14qfmBev481tZV7fbPeqH5kzguXVthvXltieMpI/2usmJQOyHhUo09
LUte6H6+SYXnrUHjBKxS5HEyPccPikZps61yEQr/cBKEM7UHgTVHt2545Dgd2r++uX942JzM/mh4
IEzX/TsaIQT//aVgyBRfv8eYRSlGJ6wD4t7lOOPBPPQCdjRSEJT4ylQ75QOvhezWawKpnOk4S8ff
97VCFFJPfGKp3gmmPFtG2q8idTw9QPP5kv3Cxxz7M+yIwO5uQlAxa3FXHA2wheyVbMNIGM6HGXZI
UpIeitMZsz/eOwtPq8UVAB4nGxanwCjo2qHYkCWZFAypucdEmBLPAsAXUAmQ4ZIVEIH2biITR8N4
0Eu5dSZsRbq8GGHSYG8NiYGlTr5H9wREMLclVz7PlhiduwFjUxC037tXtu6lPXOBb8f3KUEnbtHR
Kl1zIcT4fByGaIk9RqCAe5kasbi+BUpa8Aqa+k/mDLXSEZ6J9uMeV7B/lKmsV3nnzAXmt6HSYFwQ
OqfdUey8pB2NJRNNWAqNeuMVQm3fyBudstLy58Y66zQUAmUrQ5TioO8HqlS9L6pIbyCEw06qTPy+
SuGU6mY1k/2pOjLA6iTEcOCAXzSlEbsIi+WExKmfQjgJlTgQZOpueBbQG52h5QcBSKtCM5wQHPdq
rnQhJp8aF0QZnRy2d4+MoRBfjMIY3HeV0+T0EqkpAkTdiRYTBqtQsz4fhefmA1jBcFoPWXbGgLcq
v9q9J+RFHOjWvolD++xPU65GJTo8MImIeoeN8cgKwad39Iy1y+IXtDMNPMmW7FxgX89u36CvgQ43
4yn+5mmvmfUnX59M4JdKAr4u25ovfuMbpEJVIL3Pnx99mkD/ZGcC4MMw+wRLPLdUhO41auqwVL8V
jd1wDZS1ioxHlgtOmvzjafvCbp6O88a0uFlGNddUQylVN3r55yW21XVUhQBMJ9N+mrrwvOMSYtAV
3rchlk0xdXL+L/nBl/qbLv8kGITQoFDMGW6yLs0x2dliT9q3wySYiOB1zw1ous2byLMXyszYWpYO
sa6iSGUH2iqJyLtuKDxKRU1rM6lzzuMmtstukfslLktkheTPrwMKZrrwDDxMX2F5VTM+u9dTCBra
1Wn+O7kwO3sJzDBqTS85H9Ry+/oWhqNT3Rx+NO5fgW0LHYcgHirB2TqkdJJkgfMtDlw0jT3rADsB
InbRQIvmW7gTuEBm1ArdgEaSLpyVoKEGXPCvYz2ApJBRFPI/Wuln0X7t6Vi7MEANhxquLUWgBtsa
QFbQJVlcYRqY5NezythCgEkuH5Tii5i4xcodZxmcp01MjPjea+Ksr7vB9p5neaa2uTuU/+EjmjkH
IHNcZFSP+AlungUU2eCnsQq7qJQQF+IRivyrwsxkIPYVM9h4yVaZaSUcu6q3BhJ69sFuvsZOwxYV
NIrT6XovEWcxkHzyT1Kfk1+9FXediGLAqKlAQLXih9UR+cZM6UCONBnc6+z6YJos8+maievp1LHJ
oG+ZA4QjPdfKbHBxfZkpKWh+V21SntK1Ta0mX5x0qnrGPZbg6GymGlr3w5is+mJJ6bFXOBG+WlyE
RMNd044vI5Fv6gPs7EWDrVwpjGsEZK2SRcwC2iC4F/T5PuclD+xGSZ4kCG+3TFz430z6H3C0+uzj
j8Mnd7ztUlYeaaFh2khRxt3vs9PbZrl7tdN04arW/AiBSScYs4VUuVqFO6O/gro4o0ogShsRp7ED
mjo7CxRBC/4iMUwy53b/39z/FId2cl8xO+1k7zPLsSarTdsfzBhymLGEXYvIMYqThosKEBllKNBb
YK4tNaZvI0j2gO+Tt+OOz4tmp4/Of5H5COCfnMa7F6kgQflyKI6/ncxcgBMWDupSCaYoWSNh/x18
MIkYaNLszKKTxgcQ0l9lc393xzMePfEAdA3d5q326ah1aXvt+SDNrO9rr2O+uHt1xAoIUfRqLxjB
TdGFfUm9fxSlm9yxHYtWZRXzrZOoZEaelFB+rrHqy/LSx9Ykqimje4Mj9CYWiqy9eIyCJbrS6xpS
I+OwTDNa1nWcOsS3QvpJkB9tYpTjanNcYlIDft68ddK8I/+cQEAbn9KJOsB4sIXWp/zsYFD0GrHW
zWm/EBxsRXzNhkHRlRZHmCmFbk+rVV9uWYzGlaAR8GyMYzN8hLLORZIAgHLdiM2o2R20+jYZJIBo
kprbj31hS6Vl8jkkkoKfbex0bhGPRY9TcQljS1zDCdxGIL6DN84hyS1vZLZPtR7I797YV/HiPps7
hbg/FSSbuW2ldsW6BFWx/z7QP/Ce23HP1/WM9mAoJVOyAP8fnkSKuBo9EJhsAorxoD+etSdsje9a
CJcuwsi7F+OQs/MvvxHtPjtYEJzuMvbfOI/yj4atmllYvKOqaPxKT+sLOY+SVRL8aPzZ1itwsAyu
f58MjScBdLM0eOQ2fi/o18duKWmFDXt0XEsacPbwL9fZTAqXIIkXg81VSXRAJzLJXItmOZOFhMst
Iamuc2k5PDXuHUYKERNN6/ewfvkjgYl+Y2Gmtu93d7HHD+jdGyQOmWt+SqhcDKCM3wpTWUNkLkY5
Ph1M/qny74xfI1ajy1qpIuR7mWHTV3MG5qjmEDB2ojt//oCBflkNRSSRzE7T+k3yq4Tb4EVmkSU6
WVXl7bbayQFXnZl69kfOxR9IjDxREhwWkM3b14vphS6LHh5eiKmPxTpXgvTyWwXxBqmtdZF9bE2L
EdXKMt1afxikgeud0I1QxmaXUHtVBLx+7CZlNqmZvXqPp3dCFZq1oH84RErU0sEYfbacLHG5o3Nt
O7LLcWdoKykKmD1LsusTqw9+AKeHPiCg8naBQGOxWJQo1jkdxSftTTs9aoDUfggh4xDC8VQS8X71
Ift3Oe0bmbNzcYOYiRnFAygPaT9/9fNQ+oD2wPV6LY1/Cu+XK5umSYHF0zvtG2Bz/jLVXV4dfGG+
YQjYGU20asZtgjTQW0n+vaJr1X0XV3nd8UV2UWfBsFpNNAf/Of8AAE0h1H410P5+Uo5IsCA+4G3M
lizimcBtU/EwvZCVPu+lFtJu+XDpglzXl8WKHn/EzMFK3/cJ8dW9jqPLinIccS5E5CXRvbU4cNhN
KzW13YHd1iXlDUTxVFew9M6wElPsju7k1EWt5TnzCtIK4m7H5T0XD1zTZpr/mFJxq4USfNxm5BA7
B30X/oPPG+vZFUfEOBwxQR7aQJGsudwh4NgRGrdGcTK7uy0OB5TGAzX+EY40rZBo9ze2tG8SA5H0
7YzvKpgFvnyNI9fnkJCwux0TLVVxjuC7emoSYGPTbNj54mtYSAjZHZq/VN+MLNLiEH82Fx4XKc84
AhmuSV8RCiQbhE+gP+uC4mDfpiQHdNOoHqAlOP4cEzoA46W2UMFURUjh3MmFzhA7stNXfbOhj6OG
KJmnlXJvgRvHP44QVDe4t7DnEKb9OuLGzu7h++qHx2ys2AtFhpCsLSUDnJ3mLCoSUcc4IWbT+x9L
bwEsbi0fXA2eb/YnkSEYtc94NY/Ck3Xr+pRgKRDdUZjBXH+ucJJkKNAANhf22KbY5+cCrpD2qqRu
EoTVSw5ZhKou8SvCTeoguvVKdbWRvgJ0CQJsc8tyz8wGdAa/wu9uSNDeqp/lBAFrQIyJ2RjowZx1
BjdVXAfQAz2/OVJXddvTmfP/YDbCBkdZtTwc3tLttWeeNLWO7CCqFM0Ppaa5ejsD9QgDvGegfk18
mBM4ZNruocpJu4imiRb69mZu7BLkubpCqJats7IA7ZAXgqo7EFO3wtbVMAoOnCzyWjC4C/imlDdK
MXNen9mViUcu0zC9kSe0dmff6pF+fjAx5bKwWIhlXRDSduOq96BdsufevuuTRCd6WL1K66XfHYF3
DVqKTucstXIfQngCiUTJeUdxdPBdkEqIcwgD9oRp/+29dL6WcrBgDCw2NCoym/Yc8yySl1Z5Urdb
cawNlS2AcjF4H4CahLTfzz8WOjShdh/jkR7BaszeKjihrh8SLBiDWaxtuXvbOohac29Dr4u3d9mb
8WxfIgd8d1SXNPIHHbZ1cisjOLdgGCVR8ghlJRKmX0bT4j52fds3KZuM8p/beTqXqYj2IX4hzwse
inPjo/c4w07H92vAN1IHxoRJr+8HSHsoZdfFAIz1LvtAB4HMemN31c8IWZeJqzNjJ7WR4puDyG0O
dpsgRMrYIw0b9AbjYVEk8zOr4amiPDIggazWLM7TvXhlRwdF8py6w8fPm9rN0eJKQulys42msWRN
MbEL0by4JgCoTJXjkoM80tUhf91iq2fG8jX69RhTNkjpwOsB6uDfExtJdrHwj7AUB2uMxmFtEn22
L0E3VGaWgijrg0tECWDdL7CtgGQqWk3HecMk9KMR//4jodk72L8bYSEuWVxE4sLShyLsUrSbg5VT
kLtGRRdt4kx1qPHhiKtRBepawkR/9k5G9mr2PhgZlXUbmML+MWNnohs4N47qxWpPORwfq34x//Xa
v0OvHDXV8tjaJOPXtr3h/QPTmo3dmQgSLtbQDaA4qt4mxOOCxLNsPeK0hOL4xA9CuMlB1uLmgU/9
DY9cLO+poyN2bE7hFvBI3ldiCX6GH8rmu2AXwSmKeiIeD7D4TBSVPfGpZwQaAtgHn/Gib+Odizwe
RY9U+5y12BAKiR9hSQrK9Ns8LI3b09l+spCBR4lxM4CRVJRsqVFmCBDZqnHf7MMq2hZUtDniTHMi
TN8QNpHVq/dPSsakVyUYiK8+h2ScnQ38jvCK1fGedjOX1oeD1wmWLQmqbbk7I7Npn5PBGOfK5bpv
PxY933J9DpWgMbkVDO9QL7ZPwkeYbABqXHpfTdzRyO1Y/J2QSfvewGlqa/AWH6a4ySx1+P1lnwzH
f3NFJVCk93l9OSraQDieup+6kHPOTGYlRnpQR6ui/gVMdpo1mEmKI2mdksEA5odXLQ59C3lgugEg
9THESXGFYL5qctKmKVuQYyl9qR45PGdcTik2t4SiSqAdRJWvD8E+LzJO50oE9+Ks5bMvsgeeugyy
DJSZs3Cuo/S2ilf6gcY0DKlFjvVe9mzc2q/VWQ+9gatH7ofcMCy3tJ43HcVSaDgMkcs2vtZwKfTc
bHQTSBIqegO+6awgsMfjw/wxuzdol61/+gfBERXx5rMavpOgvWkudvM1+lI1wmhR+Hd2s02wdalK
AsB9FZTUjmNDc5xlvesed6L1AKqZ/Gt7neIdny0fSqqSAL2MxB0QR6ExC+JX/eo1En3gPbK0WXj/
m1Bb8fME0gntSbZgMML8iY+UvpwLXj/6ftNDartItKmqyPAHkf4sfI22fBKmi3DpyGqCjQR+V0zu
GW4ZLAvjHCpPO+CDRII6UBafvnIrGYJ4F5Us6fOrGBd1uZWO8KWhvgpB6/AXw9Nj7mi/9B75UemR
wKrIV+R7xHvuydbxcuhyFMEhsEmfvTWk1iU53DvIhTCaImHetb8WthUYTXeIAfjth/sWuk7eW679
dn7f3Ober/4OwnAOsdD+em5pzW9PNcQ+nAGK516pOp+5O634SooFAMF+86UAsb7OVGw1xfCxf7nh
W+YPHyHRuh3VUpg2T/q7vU4982J/4c0/JDcx6Mztn1cMNIRZJB7rshs+T6CYsui4TGQ75yJF7Xnd
1MhrffqzKPQ/Sr82YMExsZcFB2u5KRdTs4OMl7jHWku7Tl4opdXZcXqsCj5SDu628E1fQvKU4N6p
uqh2rgAOwdMZStoZTP45iuvxjPlz1YS28XLJByROAKKsC8lMwhvpHoc+WzLs/7Qn22F/wBQnirKX
yhBRbDvTfjsDYiLG7gZ7MZrVOzC8VjCp1gotMA63myzO4x1m++6x020I753G/2LipjPWkLZ7AM6p
rvaT/np6zDDH3lCQXvhhbBX+puY3AH8+5Ya6OGkC8BJC3/FLey6SzynBESbwY4JghcYUe0wjIIb1
sLy0d05V57ak5rkK5wkZE8/1mxF/e7i/Ic+yPCgAFuyi1dDiXlnIeTH07FbG03s+gWLhJokzc82B
ch0Ul6xRpah68rle5QPx6emOUDd2UNvi0RHpqJ3QJE/e0xl/UHdeQwxbuPkad5IWOkiHxBp8TsZP
0VqVqzKrZlbaIf49hvrgQ9UUTTRzqdndlsIe2vNWH+nIlhrd11brHHz8yTsEOjXjIYRh1lPkrK3c
l7Wx6iJxH7Wnk1oSMt4sgdoLv+wyBRSemJBMVWo1MxPXHEVA/tQlpUf9MBSFBsJiBDT1/1AStmRl
PtzprYN5E0dKH3/sWYMb6DVDd+uSt9HKko3T4N2SZK5oabR9930lzaNqjymzXvbYoCgrkMTOFfGE
R4FzQOcxuAbMHC2ZI1DqCNcRbJigwdYf4y1UIcfpOG53xsdua72EYklHXQRJ1dfawYyFvyhYVKEj
IFWrvmUQ7CH/r/XqVDzNM9CTQBCaDK5p3HIQW6Ip9x2oPJfp53BAD2PO4BRAWVU3O0b4qeC15Cy/
S+HTt9gvq28d+6elj/krwI40PhdW8fP/snleMc6jyDHehPFQiy1hwl8k4ofJFLs1l4L24oaEJeDv
Tn/hdPr3fEfje+aZr/UiClG68FhYlk5MV1fhAVOp5I5rVmAklLrzOTzX6R7eEHqDRAdtGNvgMewd
keYowLL4GbUxhtwxQgYdIoeofsWxUlJYesnXaGneTJkRZXiX6v/IMF5eJs8h9GQJno5AmqookKsv
3ceYBpkBMmtggzC297OzOPoHxvL7O5NO/zro/vfqrAubr/XZz8hH0DM5Lw0sIjF24ZJbGauXTZ8w
Ui5HzWpIzNDRilyXjA1bQizHklGeuM0YfohXyyiJlK8lIPtwAUskMIgw8Jb0PP0JAp51BTmXH9l/
yeaXnU3wmlz+rC6q41CawoWXJPKVl9YDQHRXmihUqYUNmldA+DrbTCORDpnNcf+Bc6oETnJ2HFwZ
QAT5AyCGDThxpT0nZyK/dCvDuErMNYsMFHvOotlYiPhn6KsBi/79LRW24FKupfzsk2lGUhWUFU5Q
crkDATYG27JmFWaz+/as8FeUXSj/FWaGkr/whkBFHy7R6lPcGUcV3n/Y7/x7GJHOLDUEChiNJ0W1
RDa3rZK/S+dzZCFcduAZo/V7+fn8iw95kwfaRI4o3QmMhw4t7NFFY7BVNqt6e7aEyHAjraZdFb6Q
zIhzzDEOFxQ8PEtlWHrdNqgmVJt/sO2Mbl7Wp+WCSGzLQfDEPhLXlTm4pW7m8nB8Ghhr51t8yHiP
HiSc+oMsglyvlYYpmZInB7TQ6uaN9BWk4jyhXfvLaKzI+Ky+0JYJVK1wVUbQ6JzykGV/Vb0GsV5i
rZB2JEOjXqvv++7tV5q5244I8/lg/LuUoumvu1soheynBwiTOmGtAXvQBIC5qXycE/nJBYcLfdc7
1uEkzSGa1F5Ogc46KZnaFASSNXmbt3zcLnryShpDpyH1hQmSIC46qI3KVxHEWwNs8KU9UXZShGGG
evRQ+mrNZest7HCOy59sPNRrpb0XFhL0pUORkQYu2uhzKSAAFrhHSdK5pewaq85FygvqT59zVQmj
sgfmojHeYiLVcQcbzarQSrRTZmyCv0OJC6shSTOVsrIJuwq+t7m0bdfH6lWZahTwnMqNbocWkVTt
EkYnH2U3jj1DUXbF1aVtfugU7BGYfBcaHQZbCVVbdWaBi0/YHBciwGlzHOnWHOP2qj6ycc8gXWfx
1Y87RjdY6Zg+bvIv8rFmSW1bbYrShZtYOs86qeWMv01hBkMMzq5773JaeUsPn8CkQBQ+zgeJD62k
1z2xXZLRy+7HeudPnf++GVuk9UfqGe8xVlNZGyw53wc7VwAddaFS7Hg0NepM8ON1OGP2iaJGgskP
FArRZVENxAEpc0ZlKs624zX7K2pk/dCDMLfr6oD2I5UCUID5whZz1HJDd+2nd3LKjaNRhc4Ie6er
Ayj5W9+bqL0aDp2oiQcXBgojB5Z747Ah7X3cRZTDswPevsquWHCVz8GtwEeb9Vn7NIorI0Fccn+L
vzMN6KsPhJh1LYUxFyoZkjwTn4+yKOuDMymbceBXfbH42lsNdUsRpZyWLWS9xG/4Vc6HTcUZDWPm
bN6M+ZPkDlFK6ySZEhPAW++x7PSIRFPxr05uUzaBwwu9L88c0iGJxb844NSJcLQGk1XWDjCrZTwU
NnGgUUTyPsGhQPT4fGkpE14Y46qXhY9hxWRFMOEEw+Ub1eHdBe473DMwQRfOSXrYVhmPPkNM54h6
NbfikiXbk3Vq3rqJiOXEKyH9Tda4vd41nrAfV0l8tqgtpx42Q1PNnl50i2wGaV+gFzDwp4Jq1RLj
YRhYuXi66mxyIqkN4pdOoToeJ7bnk/mskta7iuUKg6QiaipOCFl7MI4B9jibsA3vjZcX75bml6ky
YTflweobGYLFRKE/JONQ2O9V1KkiHFPAcsJ13RfY/G4Hdsk4qX7Mr87+VuJScfvCKISZEIXw97Jc
oICt66F+j7eNlAxzCxW6J48sZC0YaU3XkAQi34g/G6WEHEojW8zjzKrDBWn+PsDEKN/LtticRk+j
y0imJZ3Zdou1rJ/AlCe31ksR1QgavZO1mRRlCGhBjM3BL7qzhldMVVewfhOvTYt0J17FUo19fAad
u5tn9COy8FaG9cJFkZ1VvY+wZqq6LKcqlmHdjljAwRI54HKM9NRYmIp7CF/QEboOttvlfcAYlu/B
2y98Z/cIjyf1p/o3g4ncByFBETmkXJRD6jHl0grmocRhK95RsSgqINjUaFK+I53Du3pRYPcoFpXN
UdzQs+w7t1YjsspSzbfTTViCFHRf9Am+BI0sYNLL7Imm6Jku77NkN6q5QnoY6DkjdqAUaBgont5c
+GZf915awGmd6503Jkfm2nissh1UBz1d+L12qlSZb6cxtQ/e5RMnOjUDEraWD+L8qd/3S9KHwBJS
qX5NVswyAAyg9l4T8G/IQqv+YLBneRiq/OZm0JN7zik7lwcTQ9YBevRNYZTithleZxPSCKScUQVG
9PnSDbU0dn/Y8I+x6zdFiMCLGlmeuHKjbdf9XaXt6zH5IT7RAlYS+QdMWMDjq+pUmzMNR0laFgiX
MqKQt4xnPNJh5T/CRTZHgNvrye4FM9gQUSAJn3D3IB3BOR+MTCi5uOfyZ9aWlGfKyj1T/K6CfZZq
TK8FW6S9HlIee3t03+AeY61a7TpoJB1+ap92cOvm0GGhCHigsQL1TZJ7/dQIan/vPP+H3/wXdz38
Kc4KoXZ+EvcAPEd1FVgPcnY5knvR2DNHqQuRI939TbCKjsxKVgonj94UhFvoJD0oG0rmPMicKDd4
HiTpTQ9vQrycFF9Du/XSMKg5Xb5Y3lM1KQVTH85ympmkkhkDicIGaqb8nUDfRTTTMxlLguEcFcyB
QSp33/om7PW2S1w63Wvc3jfCo787Uv+RU0OCrqBHx6kDxVa71qq8gbhVl43ORo11HiRtHsh/Ms5M
qGhLtp6kj225Zvnwv2AZ5pSWzUISAIeW4qkebXXriQ43w7DFolHMkJZdX/PJPJeLMGbMA7378hdo
22R5PAw/QPJ/7QcvygyE9IyWiFdBQk1N+PdfjHakTJu2/jSvzUMHhGLQegvuiR2qpTkofTHNA3GD
tzuuQUF+C8PolPO0avQ3Qe3otCXhA1L6EqnzsoF/DeumWT2tmKuXUjG5R38mEGfoxildHdRZN4ML
opkpBJVvoks0kGEWmZkyaJPt8E78u1m7mo7xal+nGN9zTye8bBVnAhfuiCoJcA2xtz0A442kvrmX
kSod0MQc8WFjSndVik4XMSCCHk59dr9TfNB90iPU6qQrNjRy5FTzUzjvzPl8ts1eCcW98RxpFC5t
HUIwdK9S5IZNHGWbTm2T3NjoBxBLKVKbXfYADP7yVHMv3ao0UGOaGdvBMCP//MXvNw3LrzIPUrdS
MVG+4y9tXKMh9pd7M2DexOZHt79r4VQM88pkAFAtSjInm8xAUqp77ebktB0J9PD6whhTJHrryoIV
cucXVxQUHcoxPL9nzfa3g02jGGVwHl83ylxTSlKzon569+O+svq9nGfgEsux1ArLFGGmFSjsNgSn
rV5NjfVRCMo17VmtaYWQ2vap0O7y0m6Hx6Zk5124KzSvPWik+GKIQbAqLTqaGZDKFiVBjRCiZTFv
5HvaNhplfBfpc3z5CHIdR7LDhi6vWBVVFfVkt/grUadr0ATR3R1sJ6kuARQ8W7hUgnKHkFdhvL86
g5yIZuMrOqLmcuMA5lJXNGSgfsoSSthZUPXEn86O32WZIPs73HZfrCSfVyVjIWB5ChJsHyN7kF5p
mHpRgdy7Hg6OseIHCjYDVVw6pV7dVYg/40w5zzlsVVU4GA2JDF6nVBSg85DyeiUs86mb1G+YUcbx
h6JBPmkmycdAkitfNFzaifyJv2g2MeHW5n1i7ljEnV38S5g/MACeiYHqImOdL9Y5fuzdn/XZYL29
rtYB8DdeTr+Vc5bMRPxiUu+X1pDOfGCG84vvmx+D9uUl4YpRshfVaJLrBxRi50QOIcVWGB9L9h3a
7F+5vqaV96GQmO+Kocx1M5Vywt0QBNAZcpkdlWh8bErSeuUSjwynjnFbamYinxnDchOqlOluKIp7
GhZ3WwgsN2YkGa4eRTq+btNgWKjRk2kmtHJgPLFyohrqncZkp11UezuzNS6macw+w5fLf3CsfMuY
Go1s1thTiMZMxzSJArTS6/WYB17ZQylFXSmCWo9GO7KI7Yi6q2zfRnKHVHczwv9iwmelALlhSD3c
ZoptQbQRMOXXGGPC2na33Kj2DQ305/uAuwyq+ibllgYJwjWSiO8lV40n8x9uj7QQtxvUKvlNNGgI
kUp1g4Cggeb11Tf+7tsOCRVoK0+BDw9Twchipbq2wiU9g0mRLYwjmJZN5Oo85xS/7sdCBE2kXa7o
98lFgZvj1/JVNxwnhm0wJCgxwxDUIkgT3R3pVo6xQQVIXnFLpXJ2z/MenvsI9TzUbovCJ8vFPNJ3
lG8ylspVXcVje3kZ9QEQafrgiD1640q/s2oeNLqVopsJUHNPZKrTIjgtrwbXVZJsUXJ/sLyd7qBj
GFT/tp03emYp2DZcF3v4HxVwQyDhWizxgNKOr5eGgx1ctxf8qceKZV6MwVqgf8PWjOs0D8zpsNs4
GTW9eOrf6JF0g9qCs3vN1ddzhOaCpC9h9VU9AX4pe0TQnvt8FsUBwTlhLGdyqW5oZv0qMr1nmLhy
SqLnK48s8N/eUTlw0Qkr3G8ynPz4LcgeJ0GQ+H5wxFxl3+9FwKxcPTofYq0TSDR2XFkbQs/jHIwI
mCF0PsmjkrkgYnSjd2JQ58eO6DxPsubhIUCCeRZIBkHoPwcVC6gowpNc9QK+pMvM+km7FrfRB9Em
2uEzHiQa5OLtHbKkzG/CWTjfkjmbEX3kRowgRqFlf5azoxtwBfhfvCGSSae2CZ7YsnpbRzQ9dJ4j
vdTjshGzxC7iCsJT1eEEn2zHQQJlj7FcYKd6gLbiCSQ4fvvI14NEzAIKRvXRPN7xK4plXoP0FwWy
ZX5CzJXghlLbym9mRBIM41e/wNbgF8m2IaBTTPFjfQckit87+KM7SCTgIuPUs0rDSdpPmEaP+k9U
ZITNXDs5WwQHLySyJ4ctqf6OTVuexziiSGY84K+8hHr90JoZzUZQvaNSKSxmt0NDgdVagpoVLRMv
mnC2gj/0TUhKhxq6jWlsZPHpwNHRhNscVkv+jsZprE3K831O8LUWKxAJMi8SNcXsmDhS6xT4cv4k
hCSUD9mpUFrLpbr3QaCaBB/SdnEZpis06YmjUGRBFWSqUD8I5vn6ysBvRd/gBOlvEV3mOF2ieTQb
9CRgSrE5a0QRG7KAbBvLY3bFN4YVFUOM6KHH5Hy83uP3/uzemPakobF3pWEh+lUsYiVZOk3NfSd+
x6hQxcLmyD6/faSMvXY2636i+GLhR5tmuNyAJVXlrP/aOt5VNf7CsHEKSOuJm2QHHoOumgw3uosu
6PCxByqGozMgAwJMjeRgEG1tjb4+gSfp/lCQp7lVFKpKhT25aYchHUPOwbEEVMtMjBqO6UuRENB1
uYwKbxgJIxGC0wGRDgofIqOdkMX/gYwcW0lDtJVNBVutJLxwP14hOxNmC88wZ/G25vYDzce6KRjr
Vh0wlc4l+JYq3YfUkkDOyH7eFRoecFy4BOnkw580WPAvxFBIQd6iL69E53dE0A/6bZJq2g+sYZv9
rCGIwm4pRjKftclzUZ8Y3vwpQJDQb3ZK6B9uw6isusCl0olXrm0zS+eeNYenDeZcFPJBUBS9Q7Yj
uBUuAoYx4HRCCKiAI9UfknCL2A0mLDWFm4KRE7iszsd6Tpj/uFqTJ72/ou9EJkyhvoYVEfbgpKsD
bJed3vsbSoBjwxcrdfK/R/gsDPD3mOO0MqmXrgMbDGqSuRBELNyO6qAIEsCMr3lwA3xujwCrOyPS
Z0A1qRy9KS+wFI5CcDtctFPSPdddvjaJ5nT04ZWwaMtL9Ir7B8Im1ez+oymJUZp10+condKNo/FR
Bjrb/k3vkjIt3yuW+F0ePjZbCv9YOTLflWIq18X1mxkPg9u12pQmTI8ySaBQlHLp0P1AWWAsyxcr
9Q8DiNwwZ8ccZLc4PJ8cslqw7k5GTNYe4ySvioSwECwNtsAR2iqiwxC0b9t5thy128xA3+EJf2AZ
1hFnNXibHf1c9Mq9WyGie4L0/K0w8qTp4p2UYvQ/gL8RfP2FdKePCRWo+PtBeMwzdLlA+yFCz7xu
Vox9c2Dn6ED1tMfzQXgy1oidDusGmp5gXzNhsNDpFiZXQ0O8KUJKBPlPTiizY/DFqVXMP7ZRweAT
5rWbWgC5t4kCg/6NGcjii1rEIXY1FBsZdIoYHTQBsP8geS6xh2QsOs0caZaAarj5/GSI9L2Hp4dF
Z6AqvFgwtpRBrrU8bJoQytOjdVAuzSSwGoXU0AFiz4ZWXX/Xkjl3LdCxUVMtuABky2evMNPORnO8
D5mtU+E3wbl6VfxtxqkiSQ+UkWwP0f13CP09trESbkPo8icR0HzFUEpyNOL1AKCQiH20Iot4iTKe
tGu707PtGexbUKqk5znBpXXq+Jqlzw2POOXyPL2RkFqQZN0dv8KmW5b0qsCt+TS7gyl9at3ZggLC
9f77WQpD4B7Ybyb6JwGgdfuCGiuuNSQ8DbxKZj6YV4RQKtJMVVYKXNEfRwcZK7ujAbxYiIkBJBkk
vCLahWwXdpCt/XpHS6tx+VLyLA4OlOfzfP0RIwVkVaANgyr5mToWYnXF0W0UPwQdVfhgAWUS4fEU
pPhOD6SMqOCxhLTLB/9elmPSx0GDz2sa0L7mA0AhQjZc4spWQswU0rhb5IqrOdvtawF4WCJq5ALU
dQaoAUO0x2tdtoFup92JxjvOxMRS4Uei2bEp1/xZbStw8icDsgV/sSeHBgPYou3w1o+tCz4eBoOT
8ClpDaDYRE/QtLv38qcxsEKNsleFmbS2aNNeyAbh+Rgut+bl/TfcbfcaYmDAZfPTQxWAjEJIwXcI
xV8qxsKXZfv+bXXrnkF8qvObK78HMa+JWSJ58I3wG9ezRf1wSlvWQuOFgZEKPLO32FPJ+oWA87Z3
O/TWScZ6eTFYAdxKZ5/YVzMg8GRAwUZTTvIS4yOafr6wer6PNXkdmpvE8XyQUp8t4VX7jBP0onl+
rugwbPaYwWjw2bNZoYzfg9q63/dMi1XFoXcmHjMGsG7PeccOK2jvB3o+ck3HoTxZ5YNpEJuGKijH
jDAlbWrKo8werdn1XeDVburDxlyqOHl4ZnxhxXxWhpNXKTflnGZPtdZxUptr+y3//XRsO6krQHsZ
7c38f9EQtkHXkHbucOuWEpO5fGl3BNmvVwukqeKEw0S54Mqmm8dsw9H5xiilqsqZnbBUd6e8EqPT
vBndrILgtkeuYWc1Noa7+3e8CiejY7I1kO1wYaea24JaO5sz8Bta+SC3tlmyNhfFAjJya2Ha2lkU
Xf0BOOBPgn231CKuFaG4XS1jZJ7fhjiRYpCa7pmDnSKHII+pbCFepqBUnqBsO9G9Uep3Xawzgs1i
CAl8SbHfGW7DmQqNzU6Yx5Pggz008XiI6kzm40XMlCz6DQLkK9TyujngV5J1uQR/ARto66Ir5kek
D1IMCf+GqDczjyPD7sbkzYmU6My7Ep3NgWGUQJWWcihtHYYLJkGLG4ODa5sOQ/XM6m8gRYZSKHQi
UsXaxkh59UHFGPXJ0eLVDHC7yYTunsfPlu7eNI3DrJV5nPL5SKyiFd5Q3XkRXcBsqGUb02WbV8xE
yFziivdT48uuhHSnpopWTm46h3D3uyys2Tw/CK4x9Dvab94weLnSIf0i71xccV5wTIBJnTiebwHw
R6MXAXcmRsw62lr5yulCkqJQmQgvXuEd2IE1WCVoXh7HilWewv5EA/2F9omW+ai1se1eVJtSf5P4
GAStc5W0e2YTn5x100RvcUlEOAq8XpV5utPTaADW32rla1bk1r0wcTrFykQNCwHh1CNmBZK+siyK
I7sGGy+n6TU1g8nrLWRK0jTg4TI5lscJF7bySGw2XgdbHE+HlAfr90q4l6pahqaZQIoBHP4AqWeP
V38QxF00NDkvd2w5vX0oQntQZ9lc09f86RUOHcN258TMsjMcGXqpPjqLiqjHy4p09uY51p/m/UUA
7kFEIIqTfe2DMmtvgfl7pSwCT5KbJK2VRx1IKd1Q7dmDJXExlkY8HiExkhGOmGim3XS7rgejs14G
f+96Nff6uijZhMSriT2c8qTyLb3rLLVfDdJRinZMj0p7+VVO7uMDsNGyNY/qt7wtQ3VIZQjgDM/t
YOCG6yAlzdnoYrgorVP7CD3FVrwdJ+5TD2N5fWQj3cvp8GFt6eIrwCUsBYKYZBuU7yk6PujoB8yr
d1ihqxUsB6Jz8qPCTe0a4mHfEAZ7hdIN7OsNXbk4pTpTI9Bl2HyGv3Xbqn/TbZ+djvCKr2NfijwX
L0zazGNv4q35qNiknoAJ23RTnKefg6yYpGHLkEMU2bcLB0DNgN8ykchVq98dKGmOMnN+9f87fFU/
1SKrNtw2Dw3e84DXiyzL7zy/tf2Rsf8w9Ve6tfJfitq2Ep/kQY0UPiNhm8WiPRvEBxFT026XZd1Z
M8wZEix4VYlo+hUOPbHZ3rmRfqW4n7gTkU0D/1+Hd57O7aJe6fUNrsyHSWwejC5a8VZNtyeqoiaM
rE5XGdXJZGWLIykjBwOAidTQ8FF5tyAQH3LJNubZP6aaVIT0C3vFScNVC4i0iBp+M6D1HsQ6ISot
yr6hEWlRbgQvyBQ0FzRhfF/LsBSPEk8IEPB9eTjWmXHPQX31Wo+T1aamQmQp4tYf4uPMq6BAPk/T
bgmG4KMhr1aHtApOJT6tzM5N7OtFivL1bIM8UIu8j0YSUAK/LfDRAUzQfOGM0rq9bF4CaysLp5zC
kWq3Rc32+Dh1HFOToTZUloctRrgXHY3mKvh8FGeuTe9rZOJtBzqHXKLxv8/TYRqmyL7nQMZZaKw9
B3sq7siZbwICTm1aRc3PZefwVB14xFkFFRs5+vgpaeNlmHRfLmURGKOvDZuAxr0FmTRSyv7uiDPz
+5HNz8m1wj39dz+QiteMkFNApYjsWgT7dmZ1OOnb0G8Bbn7Yt5s8nVX5ekgPUx7XAbPN4vM5mQXf
bcte2IFaIlBtCXxTSy/wuOQ8mB6orMs4Dcfz19OrqCAJPJBEd/egdmuETXmMezHEgG0ULltwoKUM
pyVKVYh7pGmT5zEFBHENg2S/5MNXzdzlaJ9zDwPTvNCJBsQPujifgQ1leZbdlQTJ/1j1j/eVCefa
jPv/U8CCx4PrCgnbXB5GUBGHURybqjHxoULmQCjpvk4195EOFZaAxRwOltZ53TVJLX8uk11adT9C
ktzTNJ3yHkdE2H0S1Oq0Rj5kUTvYxS0q4cgJEBMn2vIN0rlCs6Eal8TWE53B2rs9E3a8Cfev1udw
6GCrWIcmaNpiMzWPUgnWyT9/QElDcONq+VKyhJXgCE5pW61AUi5BYTAZswe7flDP/lGzKdUaDyvC
02C2o5DJoYb/YkSN9SuHb9kgKiJH1wv91fbh7unYtOvBOzBT2DCdhfFQYIG5G6xyV1ff5RHF8Mzx
VT2jWk5HFnHFzEV4jQA+sXTXmrirxiT5wfwL7gvzueHr47Lgc96+uhEIptc5rFoLWS4h2/G9+cKx
2MN4hDcfKf5BIgAsb9qKO/PRo6GR6xnX1YEpgv3GrR2o/vj8h4MSC0nDxb2TliAOwEs07tRV3gs5
k8GU0Osacja5E0w1trwsxmlvgKF/HUG2JUbjMK03kez7Odf+yQjd+fPRbZtpuHAp0LaLg6EBC7ye
9Lpo9bwuKJ+SN6lJYjUUStE8sFNrTpzqbogp9wscWLRu5C/n3neEpmFGUIdPpUaUpAim/pfMQETI
TMh0iq600FMAseJ9GP6oVlhqFMPyhzAKcGnxz4w64DFF7cZbBrcHDYdAApJY0SLi7/FZGEtkGXhp
qrs48JKpFK2M4vRJW8bsbY/zGRAM4y9wrDVtmhaESLVHogRfikQYhtN+UF5A+aI/MBvGNaX/M2QO
KzvGSm+XOAZVcbCHeZtcRUueYANz9b/yov2nQBMgCJvMx3U5j7FBDOcaZZq4AdH8NxJKtBiKi1pL
zhlR4S4w2Mt1vMQnAXKJNog/CvsAduSXhdAkxj4m22XY9/wnYW9reHoCwLd3kOhnFtuO6GWi8g6D
jZTvSHJzVtMgpFIzqm+Rj/5ntIJijRttN3kMJXSJcmn/doOxU02nj7rZjrU3tcnD6K9kIMCAlv61
ogcXgjQK1mD8qgFFGBVA8q7l0MU6LdhJqvkY4NfRjiyT9wcALEHnVWPIRed41dIH7zNkw8DigCa0
b0oxmRRnbYELYxCHFGXuLNWt69MhcsXeS9PV0hUtsLoEOwhr9z3+MlPH9cBZuw8bP9ExvDoshHbC
YCmJiYtPXBTeNpmgXZlgzAiKbcddDAcCpYc65XXMdKvvxgBc0WNgYq7rctMz60w1etDSAhZ14k3X
o/xvY+nF//fVroWs93K5TlJkBk1muFHLou7s3yP0i8owgHAzAQ6lz/B35EArcFRTxwrvw0vueB+y
vqc6kpkgEmOlhRDDVVNkcFzsOtV27+N72rAnrXlVSQHZJKxfiWDyn2W/e4G5K5GcJvzOLf2ZP/6r
XnswDBe8LvW8wAf8D0OUsVWVQ5w3Oekd+/eGQqZOiB8Bi7xekgi6hEA506Yu5H60kWxrtntizYdm
Z+ZRgeV72SY1WjJVPFH8XBIsVxeBdqWGvniQ1G9Ga2EDU7fSmLwRciVLnINJj0QDHYJlmGKk00Fp
tfUegD5B7ajSfiHLygzRGyFEjbrLweF/VLQus5cxpK5CTrEW4kyKcG1exmGkBPIVlkYbplsAeTub
ZH2yfzESKuvr3z7GcGvxSQkjqnepblcjLTXawuSxu0Cv5IvY7KgAvjFKbW6jIkPcXIPGMXRy47+8
0/xxquLZbBZYpplBLNqcKMjgasROEpVlVKY2l4JV1p6/4ekmxZb8Fm9rKP1C2ESgR8zEWYuvKYMC
xzNIvxYnUbAzizINfG9SCu9E4NNT4iyjeB6/yMMLKqc+hlVEQZG6wt+IeMeNP7TKZwb/hJ7y6Ohh
KNV6yDXWiMT1xFcEUDTvvy9fERUmA8onBFhAEgA2e7WJQWVHYEeNGXsZGPR974ZLetC57Hkm2CBv
I+lYTx3tsEtiencdtzWbZG3cMe2KnHtJHjIm3RPLE4Q1tIdfWfRNHuWRrEfY3U9btNV0QyS/2ijz
jjGjF1kvwRa56wZlya6OP5ob1wStucYnbk7szzVfnygZWOKzHCUTEpwhhAoQ78Mf+tm25j3W66es
Vkc8sK2QDB7R3rt/89pl0oXp/hXf864DORMzdPKxO1by9C+Yd76FKXBEPH1omPrdhkmN2vc0THVl
vOdrP0ww9WEmrKEC+FFCl00eeP0WImvJkjSgdcJtYDKw+zMxPTbKwQrYv5O+OO6pJzh/pRT4BpZr
UHKltrNLJ6ebMjggBKHYhn00RSMIUKdipYc0TNioQ1Du6ZcTB15ob3wropMXUBkD6EIxnycJSdpR
3iocm/KbVQlAt1TC54VUKcXJbeRZHT8POhKVypz0Nk7dOFIIHtXgjZiM9bL0TCfSx9gVfU3V8LBA
IsiF0XYN9N0vtrNkyz09FwEViLkmeDY4ksUXc26lPUh+JqGcMP6DkxIsp2Y8JucoOJVuLUT2RBlr
APEtz8K+nnO6b+PRWtC5OFfC+sFTpNgG/i0NOnv+Vj/L03D0KFBVuqNzgQa9bY3eLbiKOJXoeiHc
USxr9bgnbRHBp+TmWh67rLZSHN5UW3xLzOWgq+yBtqODRwRMkwF4Ku5DJ60fh2x1ah18gCzZP7k7
DPR52EsnVy0JUJLDNPxLdm+40MUAX8bOssmI/vkeoF9ZyokKHjKB6XiEqtGmh6TfPUOUSuSQDoN3
p9S26kpdNsB/gaqaP657Mh4v8NiTexfpsdOSwDUSKBceZmdCrjkLlalhXwneCCYYlFKXyCd1in/v
jEFzkh5ZVbSbtjFRHtjf/3nGLfUOwiKXVjrCHOW6XSI6xNt3zJ1V8H8yoqZEz5on8+LC/4+87nV4
PXjQF9KV3R+w2GX038P4vWNP5Gk3U4vp2OE6zRv0bWw8btCmcv3b2j+0SwyjWoSs8blr3GUuSDG6
FQBhltI9YYWRi4WqCPZKLYmCwhg/5deAGVKHLmkQKn1+a3Qbd48n7fSKpxAXcj4vcWoR5TNUVb6O
3ers6ugraShC3gkV7VzgRmcvn1EtzVu2S7vXK5Pa6DlMWgFQPlhFxewT+mOB1qbhRplNmUGiS+XV
wfxJGXfeLrtN/H1JURWHKVxgQzzHUvah7uFtdQY7h5pUUOSR4kMVgZkhPJH1TspOPI4ZDpJ3HRra
F5Bs32KRjxm6X4lmE+RmYqurbO7Cw3HhkxPKnWBncqitQNKeBo7hn5aRQKsiDyZbR/NHnVI+Eam+
jQV2NDDLeBZKUBE/Y0YBWY5NyOpvFSIi1hdhWmpLWA29FPMWGtmn50RjlCrtDYe101AU5Po4eTcz
PWxM0XHKTJ7h1JsMQFW0q1aapf1xNQnYz8t5nc/PVFzt/6Sf27ptQgqoKp4SL5sE3YupvZgaJI7z
E0KhPEo4au2BFxug7+TF+HCZSqyYcDZAWg2ZGmR46RFoVM8XjaYPowBgWnswTEq3veHnNSeJHyGA
YwIosBMy8yR23XD1EyxpoSEOoYNVjmrjhU5Wz/zcJJrMVL6Kd/8xEWFcZlNGuJl53aL6v/Li29WY
RFmFYjCcTYaUZ5KtaoDRJ9jXjstZrR+3aV8bI2CgekdgvunBHu6P3NMuUJ17ZdpfBSdbhHrINBjI
ojrHB5QpTMJNAPbKN5oJtOcYyx0092MYiURYypsS4wdlbGbOg2J9CdYRqjm/P2ZSuzxUgiyiM+de
1mNgpSbQVAklg/SrK2tnsFXEuuvM4LQUhdjKUIZcOgDhFQtzxQIIEQysQ1AvH9FvIODbz5Oy+yAB
kCK7cxBKRrGZKHzm6ape/vwE3O2OgDfr9vWXfxPeTBmOVNWRpzSIzbFmALVYpz61lOEJdzszEhbb
pmDlllF95i61j9nJiRuhNo5wyM52Hul2TTc67hmcwNMBTVzJSTCZFLIq2KsMNH2mbO34pu21AwBV
FUdbPbiaqn2zLrINa3/DQhg4FOoWfxC11iT5+/QNLhVqXWoDJp3mNgO4wgoXr6s0RoWPlJWkXqzM
MJ85VzW6r6uk+X9+x35dB9Sz+t70IatMOQ62KgAZQdOImTqNGnRuNvy0NjgcUZ9NG/IyM5ltfE1C
IC29nO+J2RefwGy5bpRLyov4wNGDVnlyc68quxRLoVVYp3pjsJoEloU7SS6L/PiNjE8jmFiI/tLl
LGGoMX2jmoswxiUuoJWjPJZ2eucXiTH58tW8Iais5KSVkKijBVPyW9emt/8uAEbveeItNsOEhuxb
YUjiOUYR9OocqCI+KakEyOBUEFXPk4BaETabXNOCD9Bdb2p+gSIaxvQDjEngRehDpTJTWjBY5bsu
xiHuo35+piuhgMmCHOhRnN1Q2EIOeSD1cIfx6skyWrWv+QUnayWiIxJv2xW1UbFGIYx1Xk1lWmJX
ZEF8vrYcanG12veg/t3CRgM1ZMRswtjKXG63AxviSv7RMcwnEAVOQSKlry4wuvnl2YRQH6OP6xfk
72ILbJocfbnQhTls2yahjo9M9mRL9WJECU/drqBsI2ZR0ihhGnfdZfXBxeD0j4Aeu1y4KvbwBO86
BDNCa+/wRQA4igWYdBEHdjmoA1/RZPMPYK4VmNxkVUKktOZPN8J/WTBCxsUhOFyN44JDxOcWYeq7
eRfZN7fo2xGKAPxw3HP0O4SH5g7vYpVqdhq0MqEsCyQAucglV0FRqiDOTkAnJOFCq+h/HaSaGHCo
wzLDDAtVVYY3wndHK9hmriXrwnZtnabxRZtWm/G3Rj0ZWGng3m81OPASjz39DGGuVIdItP+pLko0
f2t1/v34d217hb4FQMf5hMAHQlsYw9CmNIu7VW78wHdCJiILOz2XEyX8q6S1H3ker2544Vf6AaxF
+u+lvvRlLjdjrQtREnKKkucpP1J6PNRJNkxWOs38D5Q5JScGT9OynWVpM7yKu7SW3Yk9ssJtesZO
Fnwt5ecRkipHtmMTnjK2Afngpwwfh3EleMa+xY6+HwuNLgalWJEKmB/RHtPFgzQywRCLVLUvSSWS
ZDIWKoXEks6LGKUu13tKVfJ9HQfMdsDJl6VNCsjk43eGCAc4EMGX6eQktyb3yjWTjMXeRVfmPg1h
s2FI3HevVZIZiIcFt78HFKr6dzx8RcNjzUKsumQe5T+VGXKh7L5j8XRydTICk0cqvSL30OfWsHzk
oVBGqq2bsuJedxWeh6Zy+bblqFuAEmC++PfsUVbE9PuL/9hLrcR7B+UrMkqklPYT7vwIn5+DbGbI
9Frz2Mp/epf0POj7gIYz4YhmQI8zTiUZofpq5je5ho5Nv860ahzCP+kJctAUPzmxGwww6rT4yOwW
Aq9AY+SpPHFMg3jVXG6wyJsP4VnOn4VjCBC/zZlZfshOHf/RBpK3JTlbP/MWDBHzfNbVfPCP1uj5
7oOFCphFKWN4mkL6NQ6PxlI5+gTXy31wl1ffNUSou93sX8CHGadicMmgH9HzMn/5H9iKEC30a+zi
ayRp4uDrfpUMTf6tbXN08Ds/+yIesYypmiR289mHmPCgnHw04sMqQCqbmZnqnaSpCkSEM7z/ZCO4
nhivp2lxRr+rwuM4+sAvDipf4i32g7sxJyOOewHHPqujXFnSg0aS95RCYaOm4hyLPOtEazI3w+fi
rgwrzyOZ3jyO+aXqgjF4rbfPaLqOEkW21aiqmINS751chWLZ8bYfVup0WskuNuahjvpoZMFjkJY9
xMt29c8T1bsvrKXpb3XDkfm+9D9bSYRnU12Mw44jPpjzidktSX09o8yrUwSTHZu8dnTwUdSIZvc2
o+hbiZYxfSPJYZvJ/0zeXLVCwjU10bmWh1GmdwBoVNWHBFuUkrtWobqSkJrZB6zyeOoqw2t6FL0n
9Pa1YHbrlmzDvLxeXYEMPAzQtOua9rHKmrglADXvw3AOhvig3NkawWsqXXFs+gMvyZSIeGQm/IeM
+9fZioNq3+eUc66aM5uVY7n34QNgoqVpK34Wj0qBR/M8RIfD5vRTR+qMPP5ehY/dS7yxs1rOCSaJ
TF1vIbNPd9GvzBCtDAOVnAtQkDhtCpVtPLUUi55Ai7H6aZYRvWvYOEFbxaj6dS47N+XkT2+2ryro
cBc3BZ/T0JkfbgTiJ+CwYXWYqV2Ms7UYltWh5kBVHz16wYkUjVili8AzVRmKnZ2ULU6vpd/yiC4z
xQwDgwHgN32BtnIR4jMnE5cuG7WKO7itvObv9O/oWJe8BwCnItowJxCdUl1DLx7TYlqZVUlYCnPj
LDiBuLmiJQsyHbDrU5tD2ZlRnHzPq4SuPtTpFe/UxLuyuO3b6O6DV/dwgP+65vySl8TFRw26kwGV
PebCZKTNFw88/u3piDsB0fMMDqqkO17q2HXeucx9CLrFWt+jx6JQOdEuIVXdx+oWX0YE0q2l2lXx
Y8YJrKDruyCDMTFcXwpuwAkjFE/Wc2Wr6ERzEXLc+PqKc8USbqIFUtSAXjrtMebq1hvL70YH8u5w
AEHMkQrJe69qBUCeZ0BwZuKdzHVBTpfP3BWB/2G6ySc+0XcK2JZEYmbQOnaZhfiYQkcwqaVICCrM
Er23ZXugMDUBCFDNp3SG0zP3RlYiF7ZP5aT8pwy7WpRLWV90X0sGhZ3/p+cSXbTnQls2oXxO5dp8
R69F0G4Tic5PSYa3CRM0pJZAKj+vMtL3odc/gQl0nO4IU3Cda+7iOJ80QzPtUdobcRC18k/k4Buv
7Rs5SiP0lSqZd2S5wTobpZJnSANeYP5g9AxI1ZxQKtegniiSfKJSQuIbPlIibb99NpKjzCcEa4ty
nv3SpayCkz/IArf53qj/qbo8XJ1RnXEYtYOUgxOCV9Cl0fGdchJ1HmudN/B8XU7qCkbhg1NyxZIK
TPUAftuBxpyYqqs2fThb0AgmkOK3YP1b9SzhqmO7a8Tl3jlfLOmtJ4tydkEO9mif8cY+usu5DDAW
wtOCpCzhoZ3lCwFxqzAjeJGfAgKH3k9q2U1eP1XMxS52PbR1QwvDWEu6zoSsDh5S5GwoJYE/AZWL
EchpxefpoYVeTCXHmnuChC7wd79io/eifScnGEE+PQBXlSk0DLk4heKXqGyA/TDpd+r0DP8lBUb4
caSIqpG4wZa2pL6t6l4iRSq9T7S+EMDDhG7TbsDmBrSDsZENRZUtHqQjJPMlNgLzE15AU5OoYreG
MkE6eCHnVI40te+5ztPzi+IZDaXJLivK3vhaYYGJWZuk5jLo8Doi8TOrsq3tG46kUhX0H7i/DCJk
L9PQ67voJF3b0GJ8nVlV2NZQhGPzc7LmUFWhs3ayRq0W4WlQvzJMMQ/251bdPc9geDihs5Y5s1dR
4fNLZY00GIH9kmwPKhw3r0Jh6PsxiVoFIPI1ckyiPMfq/KxqJi3Y1MxuqKR1DKiPFg1w4WpLLAqA
1MBgfuxPX0ylZQGauv0JCrmVV2d7Dx5eYskmmXzuCKpDodnSlKfNX2MpuvkdlGjRMOgxItupEvPd
98sajgXji92xI7mcDG8Lmhv2vJp0FnGMfuQ/U8cqVJXNTpVAdhLRZOeQi5xKMKRUT2rFntQevyul
m2md6pjKG19Wd+5gOhlpmlOab20pjqMzalxv5z548Qs3s8avvXWk5SVyJT2X32hPWrSdjD0AprAz
QAgLuCttQIKwXIgub2ZCXChH2NGTmCszD+N2jJ+k5ula6FWsNkDLh7O1XD2824LfIZVcJkoaPvCh
mC7UGfJ8CnSHvfHqgHoWToFQmHhteyJ6qDFW2j0DcM5rBxjERwbsL8bDXOd2ndoSpIV+LF5+GEDt
8nn6TsSNiXUg3Wpub5eKqYNnxCrFPze5eaaebqlCSAJu+Gzjligf3iW2bMFDoyWpHE5kDrxGYJo7
wofwlKREfLN5ozReE30xczqzzqnL8p8z1gz3jL2igimy3n8duMeuJoDhPPmjE99J0En+Fo+3xYrr
8IaRfY0BNSX5FK2t1BeHHFq47NlMZY7FtN/u4ADa0odKwUnu2HNJkRd+LTr4xVl1MUOZfYeu1PrP
+9ik3r9EN/ww0TpKYmLvHOzp3vo58T9MyqIX/eq1it78DlB4xMXpGrox7CnQ7eeqGHYGmnmjYehV
wkzDmMP8hT9U3vxH2PBWb+1fCXlHaVKoqyV+LJ5ikUXxHqNiNfnZE7EdvKb6kzfz2DMBYGJ9iy5u
X4x1TjoSiY0/w1lZVz8tbxjmbFqv2NI7W504TRTM5MeDlfNKmsQpkjcfdXLu9RfL1RKqZt+lIcku
Apa6W0u7r90Zxw2mxs4cDAhoLhdixi9ifCW1PDqSOjpYKmJLREdK6PkoZ2KU8Un88Sc9c7TM7WzI
Ma8b8CBxAP0AuuCowhDLHFEPT/4e1UatoGGumtovEI5fC/G7fzSGFeJZhCu2XwPpmwxTbp9X9ujg
r2VCNJCdPOn6a9DZVEMb/YnQ2tN8qoLqY+6Qe6dXnoXuSi0NdbD0VTHW+QRra2kkstuqLsGOPtTe
1IMS5YgBpghxqAgGgsC3raGlyakIHtYNSRvyOingrWjRyPrI/2drpu2pZjwICmHPOKanVQ9XYj36
02W8JapuR1L2oOXoJoglLQrKfcz+Y+EeY++ZZSjlzwAGLKzZM7pZd4XFWwUBiN69wKHetf77CkAJ
NEHDpu/v79t/osFO1QOcWtTO9Qe9g4cpeEQF+5YyfqJL4YIHHmdtQRfHTq0pTibQ7yexyCifjCQw
Ivw64YuBG3FGA9a21JauduyyAm5pp5RTsBjqyVzzyrr5PB9aEkZJRj7YclbqrNFBvQoXI/pKhNP2
MEM3dXqO319pJmqKuT7QY0c5CWRa+t3/tcVz5C4U7p+jJHv0JvE8VlXbTYmHer8c9AoObbWQzoGn
d/U75/KciuqTG+2dPA3/JEeIfc3RsG7VvEQUWSvtwVq1oot4+k68eCypX7tirkeevfyX3rIdBAst
QTWgcItrF7JNd0aPtk2XEq5Cy5tAa0Zx3JP9Ja5XGskVsWGWsMAe4aCk+fB3uMA9BKgyZYh+iU8v
4JUGv4Gd0ws8fY+y7vYMr23IF2Ceu1NRVUsfD2NlgwQe7c3hXoHvcYwOLqixuNBQVUjg8ZHh0o73
NU3ers1K4za5t1LXxJE9fF+gQFGR/ZUnq5B9fNKdh8r1hbPOnmIlAlksFp/EWSlnHBF203MtXaLw
a37wPjdLw5kzpEclB3zNGU7UuBdGuknd2tqnNo/x8SsTna4ljRwatqi/87N7w1mye4y5h1k5ItmG
Dl2vl940czGlKxquiK3iGCDpcq+otyhWC7QRTR4q4gCzZd31bFW8IejaJDqybqhnqap88hqF3aUG
qN9tkkaGe0seIzXPr9NnjckRAhzo2N5n8XqIH5hsjnbtYjBSHkmnuL0yxpniszX4TFX6zoOI+MFz
VrFmcKz08lnEmwxWFN5S9YPMbJUsgjm5ugkaNLXuaOzS7WbmQQMHlsO+UHwACwt5bgqjbnj13+88
bi8CQ4GDNJweTrefiEvXNCGiWBm5tuprXV9EG2EXe56zKV7gWKqlIDDalJsy3I9nu4f0/6fAi8u3
9oQtzCCAWX6OW3l8GevBHtftGFp9r8sF6IWDiy08dAcHxxFxXSMD/PQforO7nMucqlh5zcJZkRQW
9xui/TUKgsDVqFpefu+2onJ6wGNw3QQLpHcv7Dh7vVA4VvMz8biqxBfoG9Yfx2Ecd+jWp3U8b+U8
7FL+lnccChpDa2vT6eOasBQHpeDmkmfGrixa2ZaRQlqB0n2vNFd9kPpaWuLQgh4rbHR6aOuuT1VV
P6y+ha6gcCZKvd32hwL59PM1lBR1PODLCUyoNyM7cNcxTK30KyETY81YvS5z7Yopxch8KwfwTeKM
xyRaasXlV5AM0lJxIRO2UI8qn7Kjoz5mCOR7dmzrnvgdqYc/jhV+REzs6RKAl5WbSWnWCSpQ6T8f
gHAewOAC2Cdl9QDomR4XZDMM8odXc14RALiHjtkqKh8Jeob4wG3XxfBC8DQr6aS1bgn6W7x/uLy3
P0Rgf4B9I5PDOj3eeE9LRsQXamr7h+AP3BkQyJLazJ2NB3OLEghMx3G2g1xI01c7EyW1NeOmfmJS
Q3c3aGrgGLNqo3BfkadbN3RUGLhRNY4gC+rdMj6+gP2ovSZR/IlE96q7GO5Ah16ZRpfGJsm3U8iM
QgyN3VaGVp+ZYAPrAX0X1dbWY6wWsWlPgY+/pOzRWubMa9ExU/fo2fZGYOsuP/E2hhg83hDVTLBH
GaDhaH+4lna1f/x55MtyG/t1BDtQzuq4mrS7aTl8pU7uKxACfFwL+rn2d7zIqQhOUJI2kexyn/nx
6Sf58xlMRdNFoObi3WCUl+dC5upq7/Vco1GulwUFOQdvMpcyOkNpnh1EHgl5v0QUCy2vgzeq00v0
KppEHMeBTOMQ0Orm+8/2gKZWpZGxyglWDFz1/oPdJ50eRxJiDbTXNG2JnWn18c/Ij6qlIBleYcsn
73n77KkqaDT21cuazx1EkQ62ugJwmMwRHckwaeCgCuqNDO4drM36KVwawkS51U6Fm8S7Iur1WZZ/
joI6uDNv5/TwWHTclLA5RJ1dzl8+Qb0RDCWTqMNTDeF3IHQjUbskX0xfwN7eQ7puBgWjEzezrb2G
qkp3wElXoLooUp2F1LVPrg3QTzktEtsyaQQi9xzEfzNEX0C5PDIRWVT2Z5lMNixnSm6ZjdIbKrMK
5k+TFhfhSN1+YopuEVDw9MD/N9pSegGkZCDXdbJYAo61rPUVLltnTKvd152lKdy7Jr6YvGtHocPB
3IY0SfsR2gX5NJX4ilUd7qBPyvfMwfW7kuBglNStM65yqQUj4S1h0fZf11jkWu4bDJpZ3lQ1Z+iX
v11T7iHo4B5QAY0VwGcOwF/uhrQGJg0/b0UVtZQVUAWemm8hO/UdwBkltd0s1c3pLaS/c3LbTpZt
GKBQbkdpkjewR1n4Ox1T9dOvFtBO4iCjcfxg/i6g/9P8owRGki/0wlU4aj5v8iPBEuxnsaM542lC
auXU3QSlh/dQQafVal4JqDDJ6xTvcoXqwtZyfknMMnpkn3tDs316s2oIoDdNWI5hUWZzU+uAKKUD
JlERhS9bjMCRdFxdMjYIDxcGnydHc8llnMydH73K+8QwxhoZ12/blQRnSjr6UYyGypDkXcP6auMs
KmdVM3RgofUd1Ke847qPhgeaenQbc4NRSkYy85nL3la9XawOVRtqErIIKoFnoICYlghsuCcvrvUP
GQrFp+7JI4uA7LI5kAjhE2K7V5OrkLWpqhqTXyn1ftQIs6qJb3Eb3ySm3XdOU4kza3rvOEwALlRY
Wm8xPLhIp+qYdaXdQ86qPte/k0zOlCAH3Ah5KF9O1SQcEHVqWlxu3qOyoHxqq54P8YwwKtQ0rMGw
47CHVjLhKaqLQf7OeWXSPLfaMnslxZXCeVVhw+fHiIzx7fg5o2TaAMeYoBJE03boLacarkzZAEn5
nOoDgmgFpJ2bxZuQt+5NajLkkkIZgZ7TlsgRQv8wp7sdRNAtmiYwS/5qu2ck4TAyzCMGTdDzJoP0
Qk4T1xJMb/T2j+IH1ReW11ciJMLPimZqv4HEi0P4/F9z0GnoEAivvNQ0FIordGq2ObD7Dxap7Cqg
OV40TJSmrgNgVuAF+DjaDfPiFBfdvA6q44Z6wiCafyzeuCUrIrYf9ZTl+w6QXvb2+yxRlxLRdFQF
HYoGPDWVl8J7OiimugwKtGdLmKkOMaSW60tJPR30ssGPyTLPyDnOVl36BPBgmtQ9p1cQdv+y58bk
L23a8GKin8ovUbjgAuLmAiFLxqnhRFC6Ht50HL/6i3wjW6aSAZdcQ++uqHouG9MqnWw/nYWCob1o
BXN9aRCpEKt8yqd4QEfCA8+mIHOp8nw2jZt4cYt3FN/FdvqxJKK9Wj8scXv6ZTFR0zSXIjw8U3JP
GipP7aQMKBNrHib8YV6J08lJN3LF/piB05VyF23KVisdDtB2oF+OulgjmC5d8WOYe2Zz//3bm9wC
fjef+T62nBlLptoTjRKc7hhp6ZNrSTt4K8WgOz9jLtguYjeI2R1rSvG1G34HbUaVDtschZnN4I2U
dGngXGPTOurxa/AlnKwt7/LwPNtwgaFd6+weY6XooIaVhoYGRoMtQ99otG33o5bopKTiWlvrBjBJ
MTwXuBTnhDx588hlkciRyNWTBv9Gw1cFI6OvH4NExDCeYuVIghwfcHQf4IEY88mNAW+vUDuk+Yxn
tozv3h1wvCeeVMHOhGfuV2C6qvL9YY8z1t/4X4aimazN4/m0edmPVqlFleh/cYZmjhx/8CKvstLZ
nWOHTkpjD5qTof0ShYMQyS8q390d6SJDekySFEmNN/mY0pSDLfKN1w9zb4+3AMz71Wm5M4jCsLTD
v8XIqGyTIxccQnQsCqZ7bJLEAaWFO+A2ss4Mho28tvQYElwqnyjJmW66yEvrMpGVLj9jI+wdb0lD
FeRCx5C4tvPl6B1fXpFIDWuZRQviihpvQuwW6L/IErNA36+o/OeJ+TDbX9js73RmOKjq5u4RcpaY
SS4eKbxq4c2HbuRnae0Ox8eMwL9Mah5TRLVZcCzNqlZ4g9gdy625zVaXxVT3uKcyblvt75MPGd2M
MY0SkMEJCiK3iTC32gSEvQjhoF7VRNtD1BI8jIpgB7LcyPFcmVM+muR7Cqn3mtjlEjyjMQyAHtgz
12gUvhBJbLC2rWeQ+6w/FCk9+HD3YtB4Iaqw9A0/zSy0ZtUqua/0H/0vdJ4C3xEzw0NHmtr7xmol
V5SFKbFH8Q0y+pycCgmyx2vDn0/kZpB5nCuekfcUFT/aqf3gCT+VrYw0oldq0IpGG7NM0u46KHdC
Hgun6FlGJ4WdJ5MqjMwnBRbxG8d15b6SwNEbIL0iiXu+fv87ObkSLVBoA+eH0WMnZBBx5YJxYAot
vPKh9PsbasJo6Up4YdUO7kgeQX3Xokmnc8kM+qduGoVLh7RpT/ii6vsd5rpLHW1N4tacjN9Fvhjk
0K5T3dZUvQ2Kq8zg8GD5rKeNo1uszgJQX8qhcCvVROhatirgT2rZS4jIKLhlzjr952m37I35f7JR
ZRE2xhWhdtfb5h85S9QoDUKNIVkXeWlMdbtxDaMXofbIPHrs5YAod4czcJd+OkdlhZgliQ785pXB
QOYpCSmWJhgqaLVBQdRl3TMcFTm2izTfe7finNsd91L8BOo89DvtCjBbDYvNQXq9Cp3eukFh9E2J
VqAZ4Znlr/p67XyyY44Y9xmgsVbpHAhe1lSWIn9gpZldM7lH3A2VQA/MIuHiLyF2kU1IhhViEFo/
gWtZl6GsnmXG/Wwwn9xMpZgS/LkVqe5JmqKTtBsJjCXTOEW2DbbDwuDdsIRvRmKpKy4eR8RF4HFC
rXeToCpei763rfpIfSm3nYoxoEUXGnWGdHqbZujak2CmEL770mtnjBBLR45VeYyy6SzwJ7J/5A6V
yp/YB/09s8ebDEAGYMiyCONEIGS2t28SPqo6/BH2SJlA69J7AoKuB2NhmXkz1l64gGmk06fubIAv
eV+P/FvRPyN2WsKywuAnjv1MlIoxQ/fVJu2JOWrmj0D9ajHtExCewAz9rK/T6ZwKSLekdYidVAHn
Rwe4meVj987AMRbcfbvofC0n+g23nxhSCLH8f/YCsUduXMf5SyO2711TszsI2ttdETOaMHfKLpu5
i2MV8cxxsP4hAf10T0LN00mIczQE8YTvjVWhnTH16YsEfwOmMeCUaMIqUKV1Z98rw3lyxVDNRBNJ
CAXxhVFoius30wcmojgSIOnVW04zj1IihtLTGebB5l7zwGYI5xI+eyfXvNmcDnwOwUf5xFu7EIxr
jKKwo99vsbRDjoMumeo7kcyO7W1vaA+VtcAOMM/3yqoTiaUFWhVxLBx4Xpj8rlmWTLnJo+CM+2J6
C2JS1Civns0aK1msIw24lTHo0biRD1/5SkpSUK0p2YoTGxwTYjK/MHK25clsKBx+JPwb3FE8JNCd
jilNoFzUby6ZP6mooNwwgiH2xcmd1gJIwRvwxkHnIe216ywPZwyAKvZ7l1t38rNgERwn2zEft+b3
2Pd3FqP+kC6x9T1NBoiJO/J3gRyNkkmZyiHeY9Y0rYAcpeFzn9D+JeLSetXC+17rbvyfJjYZx5sY
aebh3Ty4W0VXOsCAeudS70PNdoJ3XjLTJ4PddCoo1Ura8urr9EiwGrV2OVkEJKExzYXNZeto+lP8
/Ztka4prnbc4tVzECyX8gsw5zSaNy0o9S3DzoEuDpm2qWHhbHbcbJfABdRU6KAlKRS2aH5Zohm/e
70cpfbpZHaIovbCcZFbbRkHWbAKZT3gO0Nu2DGSwgcfzeml/D0zF/cesTOV+tV8N8RCMxdbIoxIi
0SIwksJ7DZ53n2roU3G1qpdutGM9B3CaZhn3UoeK6xe7ucQaZrpMxMLn/EQqJTYB5mhJlVS8BJlh
w3cgP+/e1NvKLzcUCWjDxNEeDl7TxbiIjfKLhNmn8JuYUjdmdtX2x0/giv5yfVwqeurtqLanVfA/
Ad8Cr0Y7HaHCprmXMNPvf58cmoJw8dPg/ueiuQYrtlGa5pUfM25CAg945vUA8uZlv6q4r23RF7co
8dPmELDXzYiwPk9Wmb2yaLjpgQECmgSo4+kCGGeaO/KfoKF1FfLpdiMasORxVvwkz55C30I2jHe2
WzW/Du96y8opMAYISr4FLtrujbhm48Vj5Z0YC2bhpkpJTYwUYst9Wc83hxygDN1VXiPngFRBwaa9
8tbOiJPx5v7aqXZVzNhzM13sbBOSZmOJKJr0AZ9XArlmMezEoQ23yqL4H7/eqXfca4VnwvoWcucm
it7LBJQZvIqPU9dTXI7TB6QshRnjUAbVJb2qSQlJCAOSXpdll9PCje1v+m7SfrWq7Rv9PfgPymic
T37RczhhtA+DrW1rvCproO1hJH3d4QFbtAi52zHbWTWIc1HelVUwsMTr5OGTTIgCS5wcqDYL2iR4
sZPF58sxzuMIpn+Af9r0qx5D75xIP52PKf/CO5fxqYLt1DviYxsi7hN3aNlqHzNvnbCLtkAYnlce
LYwiQPvNqCrm5w6zxaQoKabX2mO3U1QFuhV9LkG8q04bx/J789cMxE6mo06cuvEPRQlHc7a31wDs
3yy0WY8tk+auxVGoqGeY63p2oZRlkS++qizgHwNnyJqO5LM0ARtjji5382/RncW0z1ydXMcvMU7z
cEW8PdE9DbbnthgJiB5wRlNpH/tfiEKRtM/YYYbE0TxzIj/J/yXafKRRCMTsmwbtxd07EZXZg8L6
bWz/sMa+qUOMsbVtnxY6QJ7MbodiBNJtiIzrOCWKbZuD+cRQN1dUhoE938AB3MCeORsT/aRX6ie6
NSLG0ZqUtFVzD47FDkn6rEXF7ajIGRgi7qDBb4VXnVrlfpewe24iWeWUj7OgclRjqx6bxDxGz149
ffycBX4VfgCA+x6w8+WKr9iT90WDNePkD5E4fn7XC0GwUtSabCWIBs/ykENP5jqKqxYbjaNyPGq9
zYTbXwBcoN6BOTg2geqHYe2UDjXw22bIfDEa06qAE3/tk1WpI7xoum7kLBTXUHaL/jB1VZTa6igo
aP0bVl0owdLifQ1lvADrh5Mj66pU1Ynp+Wh45tpuhBeFtO5OFHJSWQ5rwE5bTSi0mJeNstw+PIvV
K0WOU1BK32R4GM5MNusbYw7OQPuJEuLTEbmIvJ5VF6LjLErm/maVs1Hb/4RdVOC3IN9fgcWwDyM9
ALFLJ3TOD6UKfsTAcXsW+szVB9EwdjyWnB9E5Va+d0FPQRunm75eGTTpPdoio1ViAXkCBZcYd9Pq
v6Qzur1SWpkQ7V9G3FzunSqbLbVaF/52xmqQ9cS3kXpAqAulVpM8egFzS28RgKjVdegB0z4E4fvn
yoh27ZYHdoMrQ9UnjTRs3Twc6mMzS6d7CLwulAlHcV7nRtSM04lMQoMmhVht05rnDYm7oIK5cltx
Do9mAqVWjVFKBqz/v87LyM+yXvWxDjg2vrNTa/3ndyTRqdZ9mVt737mnKPXDq3oVw/UOh3f6qgEa
iP7fSxd1xY14VmP+sx7aotZ9pVnQHkk1QjdxJ6neohC9j4BB6JcWrV66iooz5es4ipqMHE2F2JOo
85FUGiyeAQK67wVTbPwCMAevcOtxKySIlJrKD1fV8QNNFvMRS6V1KKNe1Ti9H4atyLF8BRzTpFlN
fmAgjT2eku3yQ2RWYGFzCxWGXoHqcKoiRZXw8AnBTpS+RunpG38GGR/EfRbHNQVFEFw4v4LG3qZK
MIJCIhioMEFqQF1K1IMQ6/lHsKdLkDXRjP9OG780co3+uSs5psAqkbmFTTcDjRWHI9dNkb/6t5eB
lvvlhbENh9V5T0gEPYxcLDAW5bIosTbukjq5cjSnnwgcozosfNHlETaAt0AecyUipTY62aGOMdW3
IGQb66GLqtbbHXoDboODeix1tF33RnnMas3O0GjVJKvAukKj5UkyRRppNAc/rc+LciZwLvBPJ9VJ
9azjNrpnQu51FpR8myMkvIiZnPSkIBm2d4XaxpWTiNPmViMxaeMxUDlFpXYhvpB7gxA2sS3Xtt4e
Vn9QDNrZPIyB1lNTk6gQ8lNRAGskqx775O7NKVG0T01aI7DSLZEwC9EvS+YQcFsmvQzX2LCnnQ/9
KLo9u0KQuGS9Qc2OK0mPFrjeNrUxZjpXlqIzo9S6B+kbD8+WIhT4H2DHBS7quXkNuqHzPszuHxnK
yyi9raiOS8CccneiQZVl5swwsrn7FgyNJ7OtwwL2kEDTWDmxC+gxb0OrTjg2ARQUSGJ8ePw1dR49
wo09AiyW3JTg+q0UjrCCCSNjXLXqhxgqmOH3l+HWALdMqoor1nUruOWzzg5x1Pxh9fIaGWsuL0Wz
/z/GaLV8oiX3/czOBQExu2YHEtT83T7hiZYBidllGofbb2Cz5kn+voX6NDZAiYGuDYNRiv/niBuX
XcO+gJUVQCPhhh5b31Y7aYrCIBTp8M59+EaPhlfSPmF1CzLjMldDUUTUKd9pubdYIkeqteeS/M3D
F2qjMSAfSoRpwcpBjDz2RbcfbqF3suPzpqc4JXABwdooEp7HazDoTNV1P+d5C2kgYs5EOPbHWZPM
IfgvvsgRlLB8nr5K8DcsChDY2JIDmZXYyTjP8dQJCSC+GcMTsuUPnkwfTMF2ES7OG6/cF4HYD0FU
AYqVbDFi41GHBTaApBs5wxRjhalXE0QizLjF72ElHGcTqgki0WHXAP3h5vRXI0n05y2ikLGWmpNP
0PW/xpUU4ib9MecEhFnPPsTekkjlLTiz9MMJ2edjC4rSgvudXKxUszVQkIqYNPLaCZROL0r9EjDp
tztsGIgJafF9D2DABVgHA1lM3bNB44864iLwM+b7xbgxQdbn+0LIoibKiaSywGHt9ahdbTqgP+gu
LKNaMJL9rImF+COavFHViBjQBWRwXkvlS6sa+m0FbTXZuvgy8gzKrM216CqZ38T0nOP+99KDRS/N
1DUrLvHMd4go/OOd+oAgl2ESsth0MLzgUZydm1PxOjsOyFXxii5Z57KJJKhCsDIlKL25NIJdrT08
29WMtMBvytu4LH5jg41x/h2u4xHVdKg3JDhjNxdTHpU4QKd43U2ueimufgC5VjhJhdcU0VKNMx4n
tQcctmGlxjwwsP7B7CsgXl4I9p3m3ek23+W2Aj8q8E6FRDwvl6PFmIHWUUBS4ULPzHZHSg+NAAdN
reW9jNomKecEZ8DzT0Jwl5urEr7V7WD/SiBJu0aJ6T6iDAv+xMwfH0DFkm2WbhMwmlysQ4A7Fy89
eh5VobyHakfhYL4V8cXu7BUHn6xaP5sp/UN+r7CK0664q6IZLy6z183NID7kXs/y8pSuhyXNjUgo
rgerfeZnDJJa5wOOor92myKiEWna6PxGyrFZ2I1GGlt0HLuE7x2TYAe7SJ2dwHWIYVKTp+/lRtHf
W5rx/iOywL109un6gdfeBkkzPCZZs7LXdrk1F46soLZ3jj8Mw6dHXgViw79n04No/PabdRBlnv7g
I9dqkQ1+xmFTUTUOY5nfZCMYMC5rQZybTY0j9wdOmu5FQ0g1fRxvg91kAeWQId0FkoG5x7OjIVUQ
cctVWpF4ARbGmEE1woMX3X7dgrvA27CbWTmspUkGpPZ8r2aQjvZpLCu5YLIQdapI9v/YhqXLmnMr
kYwTG/EHfX74zH33D1xEs+h6EqVVR3b3DyiaBPnn+5GFvd2Ta4lSnMyfjEcmE5hCRMqbbgirFZ1j
9bul35Zx3fBGocPnCLHqLqrYM8GnKtDcfeUEfhFJXe4x74mmhOW456LQoU9NVRp1qTVXYj2qoy7C
cQtvGXArxe86tENtcrhwmbS0rgzZXcEobPqdiajxNdfGOv2jg+R2fOL2hWaWvw0U8QdGqih0y0Ts
bnPxlYiQopGrFkbq2PMMMYgS8VWwhPekJcpdtTGEBEm+7hmqkZcz4HmwvBmGRHZvzTG9sZghMMje
v9MNKt12dASJNxDsYrVDv3rsTDl2n4/Ly9pB6y4BqVCrtZxQo/LCcoqTQOPYLPuxZl2euPgZK5J5
PzF8T3ycuC0H4f0hixqw79BqvVT+jBbUXNROCdO/nMPw8AfzqpgeS62bKaiZJR4g6DfPJAF4vO0t
UEdToUPRf9PHY8HOMVISfcTQooWoP5wzWcx5z1Sz3fZJEwGCVufVEaH2OHY39dZVyotWoLZ+lhjG
Q/TFqAfryBHmtML5hk81JtSFzKYrDygGgau8C1G/vwK0GHldsNgxCbx4EZX2AZAQl7rc+Dmb7/rG
kGwo1yvvnzcNQP1yyL2m6HYJKXpPvz2QFc5+tpd8uKO8WkxnsSjbiD8CyrV0Fz1d6WrddyVIOvya
CiIWPQRV8zVqsGv+2CDxLYa/7qH0Ut4JA+o6B5LD+zwDCK/f2GooXmIIHB3CKYcKyyB9nXApx3Ti
m8eRrqSx/k1OCpO3YPkj5NGLKmxVBTnwNsO8e4BIxuzCB6U0GWG4MSUWap2iaBClFj294q5rRXBi
/h33iP4F3CFchziHm5aU88Sj6tfldDFjFHdaZLNNfE8pU0uugMOIuZ39148HNu+KpbPYKgMqQEAq
c3RSmDqUIgfBaoiiulkXxZzpLUgAuPeyWc8Te9Xlmw3Hi1wYJFw/TgM5zctLOv95qcB6VUPfgM5e
4p5QK0/UNp4Oxu9VlXbOQRgiM2IVZgepT3Vewfmdk7qy3BHOjHzQ1V6reF479j2cu7lRDNOuaghl
WCiAaGFGwD3cpmpeG8VB+p1Ui1XpJZ0ofVoWY3xkiwThH2zBflk2AvERDpHJUfLW537vwd79cLfQ
Ci2lClPjubuqcKchHyVDqj4/WoNLfnra6kHfqDkEYHpCNMhug+mOtcr3LuH3IIG3AS6sPlV7+XOE
zI0nmzTkU7i73+49nZIBzBoNEsIzVp+sEVlp5Luy+yskxaG4K2QydmdGwwc798JJGuFht5TN3WhP
XfR04voTZZFOIh1cqtb17h3KHPhryVCrvr2cSkBthxdAoqtxU3ghVuXhLp6cqKGt+e82KAFuDdJq
y+5x10q41wraD3bgcrvSNG1+XyA8X+QfV5M3a41e54LkjqEp7JqyxSm4r+oolfGPSPcsQYjMftvv
ixL2OBVWVLGZK4ispG7V7rVBLXKQOynSQWeXE9se3APVNUx2w9vV4yMDP6BQJoofNAdyTRbDFJC4
ANB4RqfRABsbra2g5uQ6uqy+e7PB1NKekzX51VGZHdmBkU3ykM/AyUY2MjE3lmMOqDuVRsBmkuVb
68Uxvu7/sXUO4ASHEmFqVJnL+XkkQGR3HWgikAEfSJUrZogG8XYCFd6QuD5GHypQL56YSQjw6P7+
wW6MKpxvP2nCj82wCNY6k0iDU/VlDXS04nI/LoPk/DsE0aH8PdZtMjJrlVzDeEmw0mdhGdz1uJkq
0htUqI6xEuY+L+ylZjCKIt3G/ImpXoM4rOF119qk/YBI0A9hwkocc1Y2TnHLjVjpln2aA8MxIDSX
8F6SAs0HWhv2XYygo4LLQhlwy+K3sBYWWmWy8GankLr9Ixe9ZlNtXp7xlzDpSbbBqXh3HLPEiXwt
CdHJ5+YlHU4qG6wLDw5gMnH7W14RDCep0Qv0ScY/hD9Irzch7VpIwPQP6qxWft24sCHqjAFVqTF+
qKyXefx32oab3AjH8oi9x1EdNBmgLD9Mhvv1Dj4Sbnpj17Zs88m4mS/cGWMb13lSVDHtQRygnKNt
W0m6cVYVtyu4T0/ZodmBWXgalZZJf9nIRYK6tBst1ipfhh5eZJlDqLOKGe7dNBS4SCDlQ0wscCLN
2YnWMbehXp8JyQrXaR573NobVtj9CjjfAES2fHdFGhw4+hkDriRW3qrn2f+1tucwsU5Gdw2fbKGh
MehVQ2+6uzqNyGHWkAlSl5HnnbLQi9ZagjoRX+vPKcahvMFfj8ST9suSn2Oq0YSkwL0DftvZ5Dyo
d8gyqGtyISqwrVKUXlvubw/zhFJLab2zfOeYWc9SDowM3Zzv+xoYGSrCXQ6YuGgQzsSscQcc8DlE
kuqsNkf2XMCS2RT7YlXmZtaroIpdjA0Iwy3ju3tEiGU3IUWn2gAowyMzKmX+7uK6R69fn46q6Cbh
jpD15qgXH+c0iPF5JYbfbkOniaDWHToHCwi2+Ro6yLXyXIoPytCS128nNrXl3CmUqivcsKcV48lZ
/2nhhmVscFpOo7OAuZzWtfCrDk52cLXrGZvU79zq4JDJ9F62jeBPITEJBgPkecuLZ/FRPMRLHTtD
BjPjlA0PcIEwN6LZ7oeEmZ2dt0ZOE4hiPLeAEgkcZxMUd0YVDQ8VdwYiOLKXSB0B85NEKQjBeUw2
nR2/WpxYNMgVhXPr8F6mg+11crAzPg1Fa6NzB4uiAtQqnoocN0drsLzgUSczPw5ROjf0HWW4zz1d
4g5p18MnYdGhIv0K/mM7y0SDqxi+57zDdvs8beJ5oKDfkph/G9uKf/6k3oP/W+V/7Hn5h1D4abno
WZjrxyP5dCtk8aFJ7HI2ApQT7wpIySm52mUqPbek4T4GxYEfyucptquFtVaLLp8G6tJozT8FBVoO
dcFrJfoVjrk21j+G2fpbZr7EgC9Y18uVuOH6MyflZUP3WLtjgagKsI+9JQ8n+0XSFLO2lKi0K2vv
Ksm35LU0ZTSqKx0q2IoW61bzmaZLDwIx0Ghctwibv+5F9XlzOXiGoXI4plVdScbdC2GJVOJsO2F0
4BzIjox+w5ZF5OwhO9V1ILPWE+j4OFI0hCOzz+g0+qoy7VSn77a4RFC3xr+n5etjdks3HtlhN+Ki
CC3tUbMdWx7BxQVien8PAdFxshmGszeWBCTfHkKqhgOmVm3oFr2iBk+WY3seaT2DLHeto9P2gDbX
8fQn/deJr6eq3p3+oj5kMalS+MAJxyQpV0BATf/JQ14QIOgsMuy8Qkp15PIIPJnCZu0maABTHG7U
7RBm7FgCck9lHEdR0cyjPOH9qsZfRcnGcLcD0JUIkCoXJQ5hDFm/hDT524I67HmAeRwoUOSKHAoK
VNB84PzoNE62P6tHFNk5QwxrHKJ2BYEytEqf1Q2bCDkXJai/Cctnm0MB3X23Z7leJ4w8WPoaLhVF
utiE+ddtU2BVVCz1UpkNaj/OPJbrpZYxKd3HF2TQCT/X0iavqRYHtYkIPyv8416e1trSW326XUPI
aM8hy2/FPsZnhCqOUtW0wCphRoVtgJr+Kyb/vOj0CQ1HHA1XeuzwRo07SODqfttqR4IaLgJEAN+N
Q0DmpUdHYKAAJT4AcPSg9IEXiBO3ym1jge+Y2vN4mrmGRCVNedNa1xHyWoVmAfkJUf3MdVNxEAMq
Nq5nlQwg61wOV8QU+HfhzYkrtG89godul48NqnFB8KEay/IIJKEm6fMkaKzIg62HFNt8WsamFaJX
/PI0nFo6MHdkXuylD4Be6HmcgYUp9Rsj7AxA05mWnPyQV7LMSUVBUDndapfMG06wettyyvfSj+Jy
23xpL1tE82roXlGTsBD/T091GcCvZ/3RO7gNu92F4BIFXUzY4q6/3t2z8AoMv1+c8Y9tzwO5Be0G
Z5vb+i/OvbxK8IP0fZU28uYoXWlx3I628sUK0TQc8heO/HxaWDp/xr/wFeq649WAQ1lStwRCp/pB
3uAP6nu4s/syNWVQpi7Omj+BaqgpmnDmqtcId7zuhlSmVScWjxhWnn5mtmhIKRJuCDgO+j/Dhbvk
4WKjC0vhx/wKhXRep9OWcBrhWij8ySCMc8/cFY4IjMwJzWqjmD2DRvY9tHCe3F29Vx+rmad6LnXo
a1nlX9RsAIuKzVJGkToaZ3UHm27GoJUtNDmIgyLmk1ylu9l3j4LX8sNuaIeJumx3guPSF1k4Xuog
kiJH/7BoKVgP06PBY43GXyRGzGcaLxrBv+9qR+OzCuQO1hLImf0ON4OzyTRZ5t0m6Xaj1KeVMgix
eY2tG/2yJgcoFos6gDtZwuyyaAAbCptnjWdbWzAV4RqH34JGEcNfS9Ke9zniK5yOiKanJu6OVWE3
Ne06gFBD9yG/cKOh0y+zJvt3eDLDcBiYBE1uLmYYHUWlcEf9R/A9dXvc0z63DJqP3egZnT+LQPey
Pbc48r1vcVUnV3H/ieERQtBWK/fO83K55eKbsYHQf+kVbZoDUCkK5iodoPFHf0v808D7y21Bo3bk
h68dg3OxdhATVy4Zf7mDuWy2r0pMCXSn6Do+nKLovFNNg12hD9zOK80cagHj/A82mUG2cRU/P8vv
+/y0iXk53oQbkbuKv+PNE/ofGAaLOrsXobMDZIZEjJMeTGHHD6PNJRIFvpoO5fCmeFRJwcbKQCvk
HBtmdJ4DvbBvtXEzi0CGBHFFwWbgsBwtIAOpUNYrheRNEBrf5jhvupuC/DDKem3hWvrvLaJRYwnN
g5o9fooGaHHG/+1dKW34udXK1m2+tlPmvSijtVbuK6dTVwJ2hlXqeVuNayroNe90ygKXiln3h1he
/XWHGl/heKDkXBP124nkowD/Knt7bfB3l2GdzF5apfv0MA9pP2eRAlVm78aL9KEhy9IEoCCbz2t+
oB9yFI+DMiv6fEgMLV29Q0mh47kxH+XzffzapGyrLuUoXbcdd5MX9b+ivAKPm7xRBw+ydq0a1HXX
jQCprKImJVSoFACVtSg4bYiaGH7fJJw7i0kQaZ/RzfIOClv/1KUz2Iq6CvZNq5NK+xW3sFU7G5r1
GIISzkXbAXthOJCVVk9C5NlvOy9w6BrBBwxVeArD+EpuMfmtqHiR84U86QEPEC4D0unWyf5MQyUW
l/ilUxn4pcoMEi70W5pf+9JzYxA01166zATfzbowmtc6wvTyXV9cBPjJ4Ie3p2Lztz+OQv7aqIfH
RGmdUSeVZ0WdDlqMwH8ctenc0uWIgT5sEErzZsWm7NhKz2DvcFYP/HokJ6+tm9rOqvjgrqmkdDQD
hIFPrkVO/lAiDVPwuVSIKIeZV0UYg/yZsypLgHTNGA2ph/+v9yGNPR3t9aqMQi7l3PiHcNaG2ydr
vbZzFeBLtjZC3soUMbevTCG+kSBnGCCkZLKRD5g4QjJHR+F1nAK4eZ8rUxQtWhgR029BXChgar2F
rdNvviEOzqLVB77yRHTO5gAcA0yIoz+RtkHHMMZ3ALz6fz8JFjO9DaSpRAuNRx0Y6P1/z8uoVXnh
pO19qmuSNeW9MIPh0YFeOJTd9tEQbqVGMTCqPmgYL2SF0NFiSivTaQLpI0agEoLS16W2sA2H30KZ
sWbDvIYnddy6L9C3n3BdNQES53pSN6/ZEQXmzOCl7+bh/9rlTb2eyLnUzm0SvKRECVLDrWOK35oY
oqX1ckvWjeKKZQDN0/GonG+JBZe3V0yKfH5zLoJhtsHy3dOPIsYN01cUED7gK/JpD3Bah9wV0W7s
xVDNkUu6kUdD0eItON8W4+U1fNk2SVIxod/rMkeydJ0jCPr+zPjlKquveB5itiMrYWcE5EQSBs9j
EHs4KyfJQgOHec12sODtJNCxH/DqrcSthQTfNutLfBfwD2lpdknDBqXyCV17YQyfnxO496qtzmvP
pb4lZMINvBJc/O7FQqhl1oL5a1BrtFAddCOye3bcx+eKXIb1QixKHqZdWV/UlapFM0XJRjPqv2mX
+8GuLb+OcRH2Kua6BR8NH63vZCso4byBZwf+sTtDSJByofHiUozHznlXn46AKHAJMalnELmKHYNd
KrSAyUwc6IjUBBwMsw6BXZ8eKgJMpHty1utaEKnszfYKQp6TXk3Ru8bTZ6CCr0aOtdRT+XzTkPpf
rr13Pcwl8XXpJO8ACAxUBq8tZmejzeec7+ZQXOStFkY/SEjcySCvlLV2sJpsW2YFLuLaAGc38tBC
4Hm2NrV3pkg+6CM+0NWX87mEUUi0SN9Xcbq6Xk7nLpQh+5tFYZQG+/hTFUHpKGDwbpZGSuzMrx9Q
DlqY2GNyLmc+759z9Z2Ll3pQlA2gTYrXMjUWNXmtXUBqc5bY2pDV7yXHF2Ggus7JuRXqza5es4Yi
RcuF8613RmLiTN43SAa9ILr/Unno3BhTx+KmCQkQbYNtprpTkFEEHJPoelymfU48OQUQ/lOhpS6U
krxaQkNIUVW+jLpyUkqgRyHu66AXctH9h26SFk+A8n7WERc2Lq2plvEL73VVachk6Kq5CQ0ZtPEK
B5P9S85g5V7jkJ3odykaAntExu0HTWGDDJbZepVd9vC2Ah3ev7WZ628jR+mXt06MIyBaSEfb/c0V
EuRL0IsU5a/nhRPBthjDKaiKdF6eAeftVExOtBdxXpuJKraUfTyZi1LpZV0LfMgyyrQc2uD7sG4j
Lpzh/XIRs1b6zoNx13zWg5GISHsCtg0J/XKIlsVMruyym/dDvD0JiVZfwci3nUiAJju7CBq9Myfy
DB/MJwiLA4HUxmtdc8/lHvHlREAJEFWDMbrAXP1X+h/I7LBvxb8TtB1FCyPzcLecXx4W2O9lz2wd
DFlxbMGcjK6NK+SynXAJiSy2C6xSvlKtIQtKyMKBjeHB7hg82mDAUXCA+A/Fa+qdr1J4ISr/Sxtz
2hggIqh1e2Ad8hr42gAXeURzBYbaZEXpS/FkVZkNcIFw/COD6ZASZ8jQO1NCJcHaZNJQIATfdRzy
bsihaaMAB81Lw7x+mcYvo1MV+vzEkBI/C4sK6gsJZrwcFTv4t5cEIeFM7IdJldFdWGaJKe/QONIt
1yG8Ro9aj7v0dSPJn7J/V/r0f+YQxkI7tHjm6wSVZgKNGqArM3hiPUOLyUpi4slWQHmZc8slcDh0
3wm2MV/cHOUzvwTuGVEgsbxVOgCHNR0tsv84bcJLXA4CNCd1IzDWCj7Xa9PTZCIiNNEVUp1U5qHa
Iub7R5JJqEOQ1SwinIQWYBpST0kY6gjj8N6MqKZd7EfefF5pOPpVY4CGGeyCBrJBzNGT4Wwc1/eh
q8AWNEX/QBhugEPm/OVhjMjnJ2REIJMs9Vkpl34bDaCyEw7nvnvyUAwe3D2pq2V/+H8mLfGMVuWQ
XHbiyEwVEyJWvNir8TSq8M+CocpKQ2K1hzKaUWJnGhLMVx7mEy8EO42J5xF13sNrFiDbA/0TlqnY
j4BePpL1DeUykcpfOeCS4tpBBquSgctEqezXSvVgn+h38BzzCXNb2XCA4VQVe93rTgpnD+3fk6fC
dyrInDIT7ItRqze7Sr+4LQUNZAGtpTHimtI6HpdEB01h5BK+MArQKBWjTOmTSuqfmxo2ywEaxBDJ
iWie5Q/i7iNgxD8zKmyOGO0UKi8V7dhC9UwkoQqa0Gr/7zR4U7a7GVj9oKOrKO928F0r+TgLGems
sk3NYGAPRXc0f2dkNhIK6Sv+9KGvDvmj6SH3ZD8YJkwj13rxMg3Aupn5V3NgSj9VKZl8CoyGfgM8
XS5weL0Z4V4F6OGm8Nf16CZpu7yCORMAADBVABwzWKUf5BT4FClkKwVZQgi4PC7+w34kYT9g7s8s
EyoWwNNbpfgzs5AIHDLydHWjLxRj6t/ctaHWf3v4pktW3t0VulMGqbmV0kFIvVXn1X4BBBoUGDp4
EUrWoN5jdVZX2cmZxOEXX4uI7dpKqVxLyodexBNjGKmZY7rK60bRYm4Z8j+K+Epieu9l+QTOsZh8
lxs7XlMas+ngXqXL9biiRITZ2s80XX0gnKlKpKnkWvb9cmb++CY0sT7cS5+aaynGDGvKYCQOKalP
kX0nd4fk3yoAyne6PLyBRF1SQm2quJG3L/UwWHT1KMWcxeL/e7RbVS41y39XnRz2t4aU444DgwC3
s6oP4W8f/P36/ALd/x0Tw4BCNuZRIm54S/BGWPE1holbSnQ7+54uf1jy7YnsN3BD4sgekhXTcNgf
aCMSh3LH3+BYdIN8KK2I5LxcXtBI5+pBwsbF8hJiRXhZpomEesn16gnhoZYaZO5T1FJsGE6JSEFx
LSdRbc+FzLIgoXIjZM3DA/a1wgOf1sKkTRFOtLHcX95KuxCeUExUpK95Trtxf+Zy1lcgYTEt6+uu
JeYK4B1+zyomk/5vSUtSV0AoKT0gimKKiBaZDW5/PB/WVyQZEJTlXPVRkw8fBe2TU74Aae65Kx9J
t3+iLPOT2ldIoQaxGkqvCoz1TturDjR1NGUwQnW01lRDeTVxIi8if6ioIkHRp8KkHy1w3DHu5sHu
Jep63KQriQ7lQTqRnzModmBrBpF6oTBA2/k3yctKo+Al03BI2vAWkM9dH5Y1q8hm1+V9eEOQFMFw
z9Ej32l8YAwu91aHNn//esG9qDJgnRapmrnHxyuByfEROm4CQX3xrzgLBJ+09YvVfbKzdUUfBp51
uc+KWlH2WjNr6NeUWcUCyKRddoKtcl1STkzS0tu4i6LaB4d3cpLslO5WOSB4qZVHyuSvHJFnUfU4
QwNdiTpoQ3yhFWlyd3SaQFeBaB639e0evP6bwTfbLpWKIOuyX5l53pVYSwIF+rH+gPUTBpCLCAAA
DGwirs/JEM5IY2NepyGB9RHrEp6SLVgO1sRKRrI+Y6yicXNlKDwhIuHUcDchqzs0PqN04pRK1UQW
0/9rt2jEUxoVf0iYahKoJmQd6ISIZTr7RbMWZBy8y8la3WzwPJ+c1V1oNYWPXMOL12S14ZD+lY/K
CkDHvBNesGmmukUEQmjUm+kSrC+c/z2sH9UVPniN16PXyAVcJeUwMUT1pxfWLEtZv5SCARhcqoLk
07AXx4+nDqxfJ/QVvc1HpHt1Bxiu7rF/A4jmE3TY8EPUcdQ6Qt5qsYU1OVEgRRW2XMEzktc+3u8Q
ZvKEiLr8cE8I49Ypj2L99nsEH6PZKmUnyenGrTdCShCLfJlqX2AWsONWLKVTTjVIVyEyMiXk9SYv
QyhEY+Zq6Ja36zZ5DOWrjM/s4D3asZerUOI7V7dCZz/6gASJrsLaPZVgBGK9xW9TA0d2MGqzj9Ld
vZP5tPR07+wD5LGvo6NAf+qCG5uH9J+1k59YOEZ3G80SQNAP79OlVQUADG/ThUsksbl6QReEMJzL
kXBlFChJRYpnlisyncd4hmbW0p8Db52tiJz2chOyQaiRLsAovXrF7P65MLfz6ThIqMAkkqMNeoGV
XtVtEuL5ojsqmKS2RoF507MXm/uu/vIvlgLyQ40CvVkkJ5C4os96P4O+aEvkDifWTsWAcm68TAGG
H6KdfVliBinSM5vez7gVHD6J8ANtCiIbn0SWLLFF+fKBVf6jMvGYmRIVFVjwPtLE8etTDmbpF7mt
cYNaqkszq2vRCEozmG+BHgFffF+bxb7BkPRTufLGMrs3X/aNehcwFtdm4xrODkkVz/olVdkGxVpO
AILBVhQ9aQJ5Qa5TmEDZKJbVCpFrSYjzX+YjxFrndkqSy2DEuYWsUXnfho8hXLiWyHmXkwFA3glT
sblskpGQw/h7fIIa5s0DOofNPuCUZJgHT0kbNcbp7CLNIUYKKZT3mnnNdZ6WnEUTq1vJGaBEB9Jx
CMMK3F0BfN+GS/Tdyb3vMjffpdxC19wChT8sEuHPRY+xrJUz10MFuy+42VyvOE8UXw5Uooj+cFpl
UW9HrFo09yX93s7uL+T4hxQA2UIuIZuhxExfsnx90NOWiEFBL5Q5vXTR4kRqkX+F9rd+guZdZ2ug
2kRD/hj9NbyWqZGYjWh5llJ3ZzjRMQsoMZwTAsUPbxPaKnZznmXt4sLVVRVetMSz1rf5uhQREiVJ
u9+lB3Pzr96Cf7/CRALZ6V3UvoMgY76RoQZScgpK967HKhWiEes/oFscQ3MG0dpsqJ0HGFJ/rxli
WgQ26DVvPRNBO/XWnnNG7w7KblI93b/55LwKMHcQumLKUD0jugBfbxDYDlooHPJExsjDxuKNXoJ8
7U1t18cLC4EIdD6S+lJ40aAHf+ISQE7U7R8RDhIoESa02L/L1PPrWiQnZJZBQTs6ERdcZ5ERvPWu
7q1TVzl30ITFFS3NSpvaJ3VnmW0YUtKkwIArgDtP5aQY+cLRqcZ757B/V1HtORYWC7MXLWE0l/TN
vQ3quw6iNT4py1VwlYW2Rnu7jAUBBj1ENfgJF2wGsg0UDLs0C1pClaESIdP9JcpahOLv0XxnYZuQ
vg158c9RCqkochsICoXMlO1f+i+x08c7taNyHSuZIk9QYMpo5wAJKcg0djeo6nGnw35lZf1caxUT
X+ippOfysElFHXXU0Z8WBNVfdEG5mUFfUiBcgH/BU8VSUgUOPTeU6NcmRAOcxb0/10vI9wwXalr+
7d8wmDGph2VHt4uS1b0PSubFLeEm5LNG9nJo9h+xU+wWCv7bIK1voKDXBmweVksj4s8hYoF9j7Xa
5QWqYBY6egd/yzW3cwLVZRPrVSJbbIhrk2D3F3IN+Acy+1VzHykf2TmCdH3Oqubd49jig7DMYw6b
xIs+VbijWYmxKEQmr1KiN821VSH7VV7a6kL7Q5znA2RgPwR9l4/qkJ5k3YC+dFEJf9cBRXJAPO5N
jAnsOhjhB7l2Ap1SbZwKYyx7OwSZNYe/vsYbW3pOGhQE8kspSuRBKUeV8YQ3Taus2wrW4lEnDI8n
ez5EzHjlJHZjtdI0fyonjBNQksFqm1H6kg8qZAvHmC6/ZdspFs5QEpSQ+1vvLmsJt8m05t+CiyHm
QwNZzA52B+6EcAtUK+2LwqJCrVo75CwDm+HA9DPjBVpAdc+4ST3Ltvr1WyDaoH6aPuAa226vdUCj
WSmxSRpX1Sv5gmXeOs4Rn9pIlxH3BlWOObUMC3fDCXwWuo77OLP3pk+r8x39pkkzU6ZHumyYiJoN
iE231obGai95wjCzjs8hUeIT7db6wKswLWAB8H0ZRwZESCNi52mPOQzbPzmGQtB7Z7pSz/08J/kh
gg1gZ9k3zonTwQOCUjcoEfRKfYDtMDIaGk6UDgnQNxkzUnuXemF5MnfR/V1mWBYBldEteNpGcnxH
nDWmV7IAnOKOP3TfJqc1JIxSLynxtPsUXkf2XTDHNQgYaUcD70sb5Xv8a11QElGR6IVZnAb6Yheh
zYavfpjoMlRJbmbe90maeYn7jcR8T06SEgvsY0jpkhwxTKvUusfvgCIC/fvAIENti2xVsK42bvVh
Pi2naxeQvXdHG2W4nr/D43ARvXPfS9+E4d7YRaVNXwlYVJDXWs18bxiYFOU7JjIPl2bwVENLEEgJ
AeFj4azHUQPaLKrtwUKIKiAH4oSJCNuE71g5RtL12U3jraCsynEDBMonmYHOytaOk18N2fyZdLvT
l+ykX9eFh9MKUZUcFOSGKcGW/P27g1ZZh1heuPgZVyspbSEhMefWziwrdCbZzq+fI2RAGEjsApKg
hADerA+pQ4oNpwK2hIyIo9M8bTmaqryjkAP4NEsMpl/WE/tFG4UlpIWRA7Ve0a1NU+3Dgx9mRxLx
XPmsuNTOkfUf+0M4+6+t7fhpZYRKyB0UV92DAqazJZNlOivH9v6/Jdq45s0Acj7XI+Lp6X0jMxii
oA46yN9E4z4omKPIysBbcbJD47vhSsLFN4uDbHBS/bNOxpubZXCb16j7aZBNsHFay/5wMTQCEzTs
thcU1xbHMcrws14ywz83KqPaWRlAnHaixiLC0v1bbbDuW25ksYSIMIwovTtYAAfCLXt6syhsB6Ts
q87KzKPF6kbPv77S4WGA/zc2L6cgv+2D0wH4AGKam164QxOhf6x+FhHMrNVNMtpc//UaUJM+OTh8
3A4wU6/PtxSZmh28pHSbAYaD2F/jUhiMIoL2UCZCmsXw0Mg9BdN0OLIU2lQWbZTzVxYYanX3UGmy
WknbOX/gjMRuM2r8yZ4L/caUfs5Yhbz2UPmYxNcb+EN+7vnj7fS9gM5rEB4aROru4HTRuzbi3Dxq
VI3lY/A+4p2jcUExmKjX8kKUj1mkwi2vsKdv0ilg4Y1yqXGwKz2TCcO8R5kfTtBkNB/hCPq71END
X6jOKdF6IZYP1bJtKuUD/bxmMR5HmfcBQEoSnejarXupvZPMW07bX84uVCq+hzeFDJtcaygIUR3E
Q2ZLWu+c3ytvyXcRuO/BBxwONRuKOtOg/O7OObbGIQXU1MOVqi0uIchDT42DFLokQR8MVBuSxeQP
p9FeAlYDjYD1a5J2xeYayweDRrBJeTNiJHtkRUlzv+KgBEGtT8g3xSsQb//HqNtrJEkYiJyLm5g+
xchJ4Dhr6My5zdItmnD9wvD0LKvBZlSvwPclBTP84eNFm2cExSsUvJsqAWe9rAfxTcleupu5VyKE
5pXGULkqhQD0MKXK7udk+3Euh8MGdteAlEKks7m2lvrkNQYVEvTYXkS6JXgy5lp6ULiz0hdEutzf
aspMZ3DIpoLwFAaDrwZV7t84PDbYF3Y6VL8I3povok2RhZ74VMTNvvAegByZn1npVkTUMN2g6Xwi
LQDdyTuDEG+g89V3Y0bcqtZh13/Hx1+Ownr256Y1VUavPJ2mBDLEYuKgm9JJa3+RyHNhDr+nghy1
HeslBkJ5s+edjxK0RFuh02wTYwNB+yX5opAq8qhkbF3rCW3Dx6z/qcSRqg75dWwNvjB3J521+NCi
UP18KWFi+mv0PyfVJRM7ZY4dqIJd+B06to0Rip95YUNqZmlmexH97gjtc2aA4d8M7KBiZ3O0feQk
WerpcQo/Qmq099dKxbtXYKJBj8dYRuXvYJaQm75XiGNsnVS/OpH4RTFSXWjyF9r6i7aQ0gzq2f4x
D41mRLGC/2fd9KCIQrzK3BBGpE3l4S1WnK6Eq7uf58NsmQ4f1F1ijko9ygRR2FhN0C/c5nk5e8l4
GXrYFIuWlT79pyK/XKIKI1Mr04KSTI4K+EvYWLQyj7PzAP9sh1+aMtWQgcC8++CIoiZR+4ssRsYL
3MVH6c8cmTD2wt6JNVmGy/7JZLuQWgzh4AQFD5FVePlehDQX3zDfgFDrK6aPCmFtTPGcyj6C2mnH
CJcKz6GWk4dE3XLvSB80l3StBvYzxKz+JoLur18dgFSLCIujX3IleGGyuDHUcoOzCgIstkRHdxkc
rRI0SPWJlTBliMCu3npMfGG8E66RN9IAt2ZY6MoM0yin2KUUEUzoEmg/ESQI0JYiFxdWES3ToWN+
SsqUQQrtFTn6f9DJ1zPT2MkWrbJIwkmMmWX4MmvLxO4Dd+PxrRGiYUrG8HMKeFe3HGWHj+ok/1Sv
abJMIjoMNe4TcaibGGd91oqojhNDFdbzOlX4gP5gamdIG+TTl7LPQnQm40phtdNJnWIodtNwzutn
A3T0Cv+o8Lm3/4pINp5cISOa9qlN1R5FVE9ygGQ4EJ8+Js8xL6OwHek/1sIC12gBiB4bKGZtrpSK
rnacN2SNf0FTMo6I/DHpPk/DKH18TdsmKvpLiCTj8rb4JdG7rB+zXapehq8ku/BmFxwa/+0TyLjT
bI4bBDzNxOJSnt4OFagbsE2QTenLrbwCCI062NO6TBrKDiYOF/SrbFjymXHPn3Om5i4rS1KJy08V
+lLbpBawPTtBrOa6lR7f4mX7emrRgsPx6TrkgdNUKRiP1cxMrVn4gnipUzdkfHbfc9d++EY9tVYO
q204EVgEbmez5F0bpwMrXI5dzbeCksxfr6iZWLDv/UVhPH7t6dVAfD/CWrp/VdPpNCMgi/QoAqP1
zSS1D/T+UjRfWRBvbJEBmVDPv0Ss2uH5o5cMnH/sohGCVCXzayD8VcUiaaveM8FCDd6vgN8LG+dh
UYY9lRg9gWvcT0ZkDOGSH8/hWmzjN96c0yXAzpeKN47OZyDkH+cxJLTBLwQ2+duzLV0rnVJYsk9v
DNRPxR/thAmiKP0BEKzbrAUo79643guJRO5zPX26GxUtUcH/MLtcE1NbytGRr3C917HAMZf4hCJs
Y0yNFGv/dVqFdtTmfAnhV7vroSBveEG2Kivcgmo4J55Ri1lWGpGxhOtKQpkSGVqO5/fHpHO9wlIN
XN3nluYvv96mds9G7ubVhKp3SNnko2LufE40LaCWgOqLPFdiM0NsmTRmUbiDAShGA9257rWPG96H
jMYAzTLro2rQWI/b0QNBh0a7H4KIhA7oFSKSyLsHoMfwpRS7MZwIrXpeJS1GtLWoeEjqF/PB4RWc
rgBAj4bK/5CZJZizbwQ0ou0J/fg1UY36z3v3mRRSLpVum+D+TVM9DeeyjOova6rU6zZtkfcVGJ6w
ZuT4sJUdr4vYZcjwi2WhYMpnUHKXLtxMIhu3WwGP60hBc56ZnBdO9QaY5I0Z9LnWZOfSzFjldiCf
MT+p0P2BkHJI3xeoyylbnvzPUvqSOVzI7AiC18ECyZ0Mr312RAyxmxIqGe838l9pOzu65R+3JzwL
jtkPglNTvvSTr2dnWP98/YU677xoZ9OPgO1e5cH21NPWebGotTl6izaW400ghWoTo+leMGrEWV4g
dqvNYyz3YhNMzK8POqToqJ1LMhDmhcl3SwGXznBfDRCvpQ+qRm2/H2yp+/qQQpU7jCHtPnBKZVMN
x2N15VzbV73bzMxaXjEyDXmJl1OK4GjDsKUmqdnb/sN7SSfjLTiIPpsOF+bVSCqDNYMc2vC654WC
9YDKAzRfpSFXqqOPf07+ETNRTVD7VUqW/OvVcBUZzLYzDpCuuG7rMJ3EnsMNQySU52Lh10WMH/Ev
GcZGg3MaMjCTyA4GfwvkMN3V+i8Id9B+NnPdIcGidRISmK/B80L5MVni9zuy/bz2wyy+7QexeI1L
4WvYm38BxVap13tWKe/bjPUVxMRnp7qJtYhBxGl1UKNlr2d7sUnBOqEX0Ze2DX6uXSZDY8AmiWiL
O9hhsT1B74d5ha5CW7hD/u9WeEOKQHl11lfAiJ6nYs2IvfPZIP39b2yqeqvNO3miG3Nf2chf7jvn
HK02cfZvFBz4U1aJOCwbOzxKtbS0zQcLn3IOEcgBPsShkCdm+Ocs1JiicGqky9GoQUddVlKIDANF
OKr6hzCSvFsSul4pqhYPcXiL53LfFrGuHG7+Pi9ToBRYz6VFqeLRomI8jf3ZQOZ1+GuHyD6aT5Qx
6dOS3Aoc3KMuJlJNwnTuTQEcuWPyIwvFxzgZ0VcPfScynxObhNjlHCF1DgJCPsjUI9RokoZvOhky
Rzk6pz/BcSrZrwHwtKDwIME6FFY+e5TwTGuKDo4HYrzJDG0tZisOc5sddXjV1BTQ5K3P9qHt4HgC
l1+FrlLoi95uflsv4hKS29GnXCPa8ZRO8l+8bt5PRdmqS1OKBOye0Ndue1PhKurkoo59fQ0vDMbK
YR3cIyLuqgYWZxTRCaFxR2KSYKXGnvarJRP5gZB/iJpDMsbLbSdRO++rIS5QvR8qTvFP5TONGEfs
ARXLE5wQC3SmZlyb0HxlgJ1n0fZxJai+JDeIa4wygMnVuT59J7a3jaWa1f8FVW2xnCD12TjeY/Aj
wU0OcQzv+MT/oukr5WponvrNlb+AVU3oqKiQ9Rw7nGzymdvmlOhS6no8BlgHvEuQl+D60rFRW0ik
21JvPHfIqk56Kf5y8nQMzHM5LcwcF9qLfXHnLtTBJcCkonsU0HkNOx268xYltIsfgwgiCoBvgupW
XQewzE1Ys6GHthxJkYRR+Ep1kU2g+CsCCfg85lshr+4qPVRmTeVPOvHL5NLMEc2YgMLN8jjUThuv
m5H41pqXidi86fHuWpaFRlQT8npCbVb2/EtDPq+k/Ddp949ULt9+4B9XJrvvub+s7wu/zhu3hzQM
cVg43nXAO1GUPtwH1LKNFM4rAosAiW/dERY5UduQWOMI4S+0tbxryrCAFs+yZ5QGZTH+ybTLyodJ
QEptgWS4p78lxNirwX8Ed43j5gGO0N9jwsVVttvI2eFtesIWcnp4qpmKFoti0dwYM2/Q1kjHkyt6
y2TKp8FvPBqJeI8yvvGVPuV02yLPhM/yJysAy/Zk2e2S+FmrsXURC6Nt+IOTez8bq4quBMkHa8nK
h+a+BNbNMnTbdX2ii1cXic7Rctc3U/1an8T9MhzInZ84B1ts/A0zh1NNzGH+e5FavNPOKFAWe8x+
ktcsNucstuaE8Dvo03ctd6QpU+HwvXnAl+dPh5GfTG6hwrcpGpWxq8TpofqGoRp741R2qmOoom0S
mqnYf7HtBWFomdIoqhex89u3jSfTh8z1sOKsbZYpTRwhAqnyV7cgOoooFIGRKVbn5+H7rqI1hdwN
AMCd/e4Ynp5zlufWeEjSjZWaX+d0PVWg0hbzptQvuCWGFoaEY27FuJlaXedd29Ee+j7+UBx72IAT
B/OrW4E7X/4HPXwsoP/l62/tUkq4TPp/CYmBaCq7O0k+38kydBy7EYPkoKrA4RPS5gooQQEezmQP
BwGjPUSGzNrdP8/lCiAd3Hj9EtaE9S1AlWtbBJYX4AebY2XaUFXjUxj7KG8JGEs+vMWDdZtdw9Ho
roPYueyQv+56qSfxK6SgI62ZyTHG7pvcmlbFG4eLyTcUWEGLCK/e1GvHnepAiZ7oex+LsDHZEJM1
HbVra8k9TVe+vqSwqh6Srb+zT8/EQqk0zFm9mWRu+pvO1ChZvGDx+BBaqooAWwAqi2ZTSvxxTX3i
4G8zaXS/NV/Ob/XjqNNVYxdg33OPb3+uGBz7BdXGJ3ruFi5UOTGC9JvcQXSRD2FuGdruLbOfPQGE
7khfeCfsk1MN7PG6vx60kLzuONfqY+Y1W9PEncLFKg7rOJhPCQE8p3R1iILQH8NhKEtOH3RIzrDn
bvv5+pD5r9TohjsDBOmlUuDwicyJHZ7AsPEwpaj/SMNee0h8ugic2ppXPHq7U3jcCy8Sfi3xzYov
kzDAW1RjfSahYHciV5E/HTD4tdvMsjmEPOHjIgXkRWqA5cu1J2UfnNuQ0Yby+mKqAUtW+gegIp2p
3t78kjqih6RKuLvMW6lFt7RydepKVtw/nAO0ULlmIU+ZEBFJk73265zmkozOLsM/LRAl8I9Bl2wW
R6DfWnPHLU3vaGGuCK11q9KZ1VYqF/uRzaRXcc54Dgi6eX7tNPd0cWVFLbAba2FLDlng9t/lP42s
Yb+ni3AfpnAXdA1wWb1EImAuaOdPl4n3+to/uQm6z42lorhLLyNvAFPgamZh1t8BKyRNn1xIXu7Q
VOf70xo5TugLLW+crBDW1LLXSr14I2uifv/Jovt0wYhNVDYAsqUj/oWy5cUai1+v8FYNSAFdBtSO
fS8i1VsKaXj3Lit8fcQX6OIEJas6Tu4SGZUdPsXJ0N0hWlzpXsvcvY6Zj0M6dicFm3ONF3h50fuE
ENA+21Gsr0L95aBydwVB3+657bppuKGSa8PANymxsDtWmReBLoBc33f7O4GNJ7yL/pr/9lYKhcJy
lMDAzJGqm4L8o+G6jVrUtzQ2jyAw5oUZ8qaj7cTDnsjBjCKkCYXPMvW5KGDpZkiwal3GxL9bMcwZ
SfYzqoq7maE8k2EpQPdBeR8G5WHeXQj03KvdZftdIK8BlcRJZ3US1Oi/uZ8GkKE2AyvdO10jW7Sj
rh6zgQWTb2jAl4CkWOoBV2tf0BZvbgQIWTChvGx25Lyyrn3uHz8BUL8Bj98ocHiJ71PWvIoaY0jG
nR+TJhArCCemoEMPc4n0Vmf+UxnD4OGPzJoqE/w2VTzaaGPhoGa7jnf78Qzw6hU/ETlX6A1zzqH9
69RloYzbWqmAA5715+vnzYSo3K0jFKggwqjHz7nvDUO0j1hlqIVv7zUTvE/qn3y6PnoZ92bLRqr9
65V3OnR4CsFk0wjS8n0/sFLUicUnq34Qc+Z4I/gxR6MkruAIIV2YdDskVjekxJs9VYJoSUWuN9HL
UMmDMH5DJ7ADcf7X/KOIccOQqv/01uSNjJPoeH/3rY4MAcjSmlaLWBIkHl2VkRVnUvQZhDjmfXP6
S44Rfq1N0azV7c+lLGFc1lyPhU6nlMEqWnZR40TFqGQkvaoKQG6KkRIGnH/MO1t58Tj1+vqj1Oor
AJbvqsi4FXzT4ga9834VcKrUyBjBeV5YWuUEihwDXQqkqQvzfgm74O9gcFl8ZGrjKikslyYpAmb/
B8Ft+KYJd4MFX1LrdxjusieQT2P3HFhQMVMiT4y2pB18Hf4Bi2LCYVEAtCBJMP9betinvZOPO8Iz
uEPv18kP+LXI0/+3e01FJi4YdBbUr493jnDUY8F0cwgYU+vfU/uEHaeJkruLnX/9Gvi0hEMvPh7W
dVNRW8W5nJYMZs73te/M2qMwlEZ2MNZgF+XgBoECHjYDnf8d5w0GI3zZYD8rN8ODsr74wEhe108/
nO2tDPKiHtnB+uSsFysxwj3208+xviQy5r8FQuGeNnWeaXxV4bhwOE7B5g6r7SwnT4SE8lH19zx/
IHaQzCqiBqzzjXlMVyB8KM/tQZr29/uj4/ppIU7IRa5fSNYu1lUHgZ2aq/G8neB6A+GduRMxIwjj
R05Xsq+e/gyx9EfJqh0xIXr2lq9LfZ+tvR05jgAw4dZAuKD+2eOUy9J+KwP/fzM6GsKDk4X5WpSK
B5z5ToC1T2VQAg4TltxKiY2McvG+6qPZVr02wNq2nfeFVKDO8WrDSmHSC0LXsww8F98Bp2JGHJbF
X1CEF/jMUpb514i+wqj9or1LJzHLh9P0GbQ5sa3yvmNW/L1o/vmuMWXVzzonH9ob/1NWlzP8H59M
C/r+iwuGQbU5vNSytXJDozBjs8536tjySte3ZSBB4ecW9lto9s+izjSZyD6P0b2LWI39b8O1f2ge
cgUDiArCKEbM/17TeR2k0meHc4dgE4/QmeysL+RGQ60XKEtrafLCp1SbrUXS+hc5gO1MUcCSlT5A
OpOr5jQJ7aRynMbPhBWTh6fn93yllv+iMls22O53Mb4OkK39aU7JqM+ucmC0g2+3Ix3P0FaYh09R
b40KF8Pucxvows/DP9HRKK12K+9uf4A8Czcz8BDjKwSYssArpLAtrMMlUPWF+iXBoL5MdJMGWOkP
GcOPUvBYNVCi+9VtbBwPXHwrv1195UA++4qB2M7Q5juY2W5FMDylClVFLu/1GFgObAv4m3E8rZtX
/hwAg4XBuMx/TaLax3viWSU9jEtBV+3liKXrBzXLsPmA1890ZJ6t6960oSGlSJ4eTpcX3fUPBpjn
pq2JkZgp6OSDN9vciDgPVDCnwZ0d2vTqbU5+j9UfMT471Z9lG3BTPzrEbRXSR2MNW0AyE6IgZ98g
JC70/b4IhehLltJjJ4uL9BLE2CsWmGE+P4gNZip10ftvFejwvaKjoQIC8dP5JMJzNYcQK5FALDpx
SWyaDoNngj4rukS2BgPROdMbxf81mAyl75MtL9Qpm4u22i/KWwd/CsagH7931uLcQa1pAGEJbK9Q
KUTGrWBAQmdWsSqTfCxNJb5NCKYJ+8p0ShT24ylueROVRMi4dxvEwgq2mAc3pmZ5dXYLi8kn6yPU
HOvlkEgk5lp0yN9y70ORM+nZL5gazrbjAsQQxk8II3BZcIXREfARTJ2d6qeP0aFVmlVRl4fhftjd
7N1lZvqBQ1OKF0nEVlvdvk5/DC2IJNfD0INEEAt/qIKhVAAatByQyQFDPStbhgFZ4x0QmMeouEXo
nBdx1sspWWm21WXj+aAmpHOVa8IEItsC4M+VTAs+r3gbl9BtpKwgHY4vZWZU5Y2o3EkmWV3KXVqq
895thr3JTK6MLUO4hSm7juIPREWQP++wKEuRFZYNM9GFbh1c8qbmtFjb/MvPVBqjZthRXGmD+Dij
8Lhl4/CjPJcFFe8XmJawrnd/e3/TXvL59E4b/btYTy5W4dtVGa0EBFd+8FTRTIIXEv1+DbUPwylW
wcfWgCqCFdEznEaje8Cf2N0TYn9i0Hb0PeDSa33xmjVr87QP1s5gh0OuSjXaUdYKl5mhqOX/XsN4
bKSKTPb0esD5WvBuF1/twfM82gQwaoTspBjrNsWLslZDgrinwz5yeO8gCGtZm2OjFoyfQmg3VkQ1
080qCHJzf9PBhKQ8qgmvivVXHQzPF2USJSaZ1lFHpGVl95H8fMLKqsrl8gJStghDKgvGZDfsP9Za
yGkKOB4tHdb0xoUm9r7NjdE9ZmUmAp+XMR3o9jvEOHLfQx/hT9WGfvHJ0KemjsDv2AHGOJEHgCCx
8BmqmAcKLXN5R2QudcQc6fCodGn2RLDYzgdGXPSQllcdFJNkaR8pOTVytuJYMcZzNypGgKjZK629
DgbFggNDh7AK+1RLcVrQNgfckkp4hlnO5RwDIEfJkI6HDVY+9sZO6roSdOmIBpy6120tnzwB+48G
k5Kh7vWt5ZX+f5xXUIysqXxketH2AmpEn2NO9sb5uFg/tvlwXYxwq7VFNIuY/15V9A7l05S7ybP0
EGiHqD/I1FA80gY+sYtZrYO53d89ZQ7QROkbufBK9GJXeVgptM55NtPZJaF8vP6dZV1rMTFgLble
vjVRKKQ74X7Zgo+uZQ+rz8EWT/56ywcAFZO/K6ur5YnGJrm7muxxat9CR2JP89g8D8l3PGRhMNYn
GDO7nyXwQuj+Vboq4WT6+egpH7fvZDIFw6zQCUr/wFvcs2JSeGJB8emOBbtt0xA5O9nUi996YcjJ
YyNSQNtZlncSVYhjuGKeRTxHw1TVXiRf8eMk0WzEvdijkQZdSfO6PI6nLvTX+7FO2WnenyfHvoe7
T3GXit4cYbLM2iNC57PF/A2t/EYHuH0IWSaMX/uYmLxRxDYTUILK2cAfj2nG8CwtPuM10077xMms
eNQozYFt4GAZs8jvJ3e7G3Yla52mq8j/xsBstySSYq9grVjWkMfGua+A1fla2az044hFfmk57AeO
kjf7tGKbr9l/UfwNkufKGAfA9yhVGw4jej3215euXnpmpDT3apXK0tPCDBECNs3kR3QCT0zoTV7T
5Ou8r9j0NAZtf/U6CSFuQ14OqG6/iad/geE5Sh+W34s1aOErmttkqZ4FoXkDLBZVBRm7TzLpP4Ca
xKYbSiSxliSZ9HdT6aAxskGsFJH3Bv3mwTun5qgIP7i6ok0y0sSWAZJTBLAJbbTCuET6A2s72wm+
odjVZ8sTz+Hm9ln950JHZJmWGDg+igWe60MG22kIiVuMhYTsutK+uM9+96FHrNszqxgb/7G9bl4/
//9SklWJ9RYVbeOPQZ4/lFnss/8GBivRUjwSIZxqquigBoDKlhlOtHKn76dQVYYcyJZQJPWJwrEm
zU22rDQy1wWYGNYZi4XpYItE+1wIKTyKzmsFO7l7BQVt+khJrRRNkWEL0+BRZYO44olA05M5zQLy
cgTu+MeziTC+BHtItV2fzlPJtsIC2QooCNEeDSKHuCbvBz9PuWo8xfIuwENKuLlIZDXIbXZ2UGbj
ghVtafB9PQa/3FQld637cEWcYLp59VLQUgsRxBh4qaT0bqSAp+Yd0fUBrmMDK6KsNLJaA2mYADEq
jQPk/D+CD48cMAy55aZlFdo6bEuqIUo3EQVnH8nJpRk7bI5/5vqiZq9Aq7arberQOqrrlplyrlXP
krEDtbDGeK6VgxVd/yXAi50w7D7xsItAFz9t14/uhLHGoGw+8BLlu6zI4uFTgInsKQgOH7P2mIKe
L6nZEAWxxutPOp6Z7REJmXkTZwVXoKK2hrqqDLF7Onii6thOTt8z04ASBGTAjYMNwZ3Rh1LzvRMn
WLGsmlApzL+GPjC45jNkHWdeglhbZ0EGijZUxvFt2+0+UtMC2OSrF7una5splyvunPPh3+JttqOD
xMZjg4uOd3poGEy1bzlLpGsF0o5SbMDCDWyMwlkpQF3QUB50Nha79HhjOoQdv+jO2YyRPIHmaMQ7
MG9DxgBb/Au4Xt8ISyzcixNzbgqHW3L2fyH/i3E3tX4/+b+mBA/RXb0AKQhIi6CgSzzXpCOQxO8h
ngPuKBIA0v+FeScJ6jbr3dNOXpOQlqVTcla/hhb3d8p7dAEwkZfZkFVJS9OToHytgzvYO/IzbiWZ
liNYNCVNt/ouj09UC4MSuNAAaR7Pp5rwE6fF3SFiAg77Le+bIJvvhHUEKbUmxHuVrpgT/T2Hkc1n
GUdIiT14zfmhFaipN6z9aXDmXI0XyUnbi5AjTitGHqHjirqtCBRgo5e8YtepXUSjbcxPtB95BpO7
gKN+a/iFQm9LR0F71MOS6ROqkxU+wuBQd0AlLPjNTlpJNbkxXsudL+NH90CGYEWntAUEuJVaLozx
FeFNVzX8t6lpeUkBZaumMoPjROsqt7MTWHd2LGuxXcKYtqY9LLzvhhk7bwkyMcMdunyhzEW46cH/
MlUNfbxPhOVuaA1wIyupi4hY9utxSi2qk2fiy14wqbCSCYsJzzkQ18ONqX412gj7QHQY7keJF9r1
L8FBzf1N5HDN2pX9P/9rsqFeEuC3JeQiHAtJnXOPSqYH2oh1KPKwbAvVIPrRQBHFfyG5yKs6slB+
hj9WxxuNQJGLpt8AWsiSV/O6dIX4dK0TJBxd75SNIkAnwdob1e/euUe9QTDrOEa+SySoW1grL395
3X81f3I3ZC2bN6v7usa+51tJso6p6fjtfQ89W3HLWv5PxegtTodGd3nmF/NuEl4U8dgqi/+pFP7l
LFu194teRsxA0x+ulQik+JZSbV8S5wl0yX4QnJ2APOg5WX0rNi2j22YjRPk/Jj3e+iO+z0yWf0Ww
ODgShXihuSxca15vlbPrKqEgbhqloDTAq0f8dCOsozcAG6XlLi0ovkowiNZf7qpsKRrnVo/8jdYx
J4POIM6zurGx70+JcIfORfrE68nJhYJZPmuW+BhnSoOFHKZqJ+kbOigZ138vrw/mQ2KK/YdTi291
paCEbzyQNlvGp9Kkk3VTJti+qst8mMMxvRNuUoy6+CYI50cajM1A7svsHVt3Z3sk8975r48FdRck
WMlK0BRYAYj/nDo1e7Gyk9q/WLGqHFNKZSyDWZksbB11MEqdC0FnZyKrOY8epABmQe/QBRkigDsQ
iEmowlMRDb3JJO5YH2KekjfvqEiqYk7FY7CUhVYEpz70wiEgj95nCLjXgwcNN33tdyMtxatiI+Bk
zOrexNTxnv3jde1aUNMbkGMYlc+VfzfuMYCdfA55M+hIwLDBUOmhO5SLD2wprY6NI5v9oohSG94L
fiJZP0oV5I6b2ya/Q8EbvoqpSuP1aR7GcbupV7F/uie+9Q2/G5hIRZtZ6vgReTUcar1rl4pjBeOd
Ri4nqQy/yOAA3dRoa6DLGY945h6ymghU0DdUb8+Ilk0qgohrvTPMwAxhrWtN3pCTCgT4/wCztUiq
6ImPwIvkgZzAtiopGcwf6HbrJ9CRnr2OvcUbOzN8YU5LtCR051x1iWFCAoPuCaj00c1qAHHdHahc
oWuVTw2gSHqtjtLfBLCOBQbZpkmMbv5DbxgdsrN0cSiNwf3OtF+HymyyO1Nf4QMJpYggfpSdesBw
/lKcqfKRVSZC+8YCN7N7iL2PvpdaaYxgDHqSxwShbNDrMeto7jHl9kWjQyZvyTzdVBrV57L+vaTb
UM2n0FjBASqLNkYetJosV/BS4CwrkBVkQplmqJROyXCf4/+jyrCUGEvOM9XzqNHvFrmF4C7xFXSE
9twCLgrH/UMOBqGEyb1H055dI1O4zhnX4hXHVZbNTC50X2KhYhwV11eW3Mlkt9ajn3aIvDmYqUKa
kFqkDbNoUEooAFASQF35EKr1zp3zepa2X7yKTILSpQMTWX5/pRoayjA5+UHvyMmeJTWpFy2GENq8
/iwnk0pJPL7ec2gOCYv6G2wID+AhF6x0LS1srFeXmzhwBgmWPpE5ltnfpRs+KuYE2+rkA+ri368G
LqqEfM3LEstEiCzM73Z86Qf7Obp9lGfrwgxsqI42420CwGaZ1JvX9qGrPr3zj4SJuy1Px52//AMg
3kk/G5RkDEj/l9UebUqbtHAtrxz7Ka9pIFIHatLIUaYFMvrDMsbNcfqnHU1EdVCQ8MmKuVmyAIZ8
MjvXQZxmRSYSBRuHhtPE/uQ/Ab6WZrHYOn6/KFvd0puiZHreMpJ0nda6yMdRBggO4Y7UyJCLCBKi
PWNNIerIHZcasKHv9I9Uz7q2Ci3PROM9GBbeZIOJ0ezZDsml9EI4NfFWGJrqLAdkm+hgAx6mef/5
WxBG6U2qY7qOuk+Igm05kYP3vWUDwJd2J1SvnHbjubuldTr58EyQDslEcTkRDeeT3ZqHXxLi06jM
E/gqscnSspFgBWu8aq7BVyKj8gbkPQpoQrYzRpTqirlc2i2G4qO3yfMzbNvsOO3XX5PB/sy2LqJ0
1vF06WOPEbXdUBEAOWraurKaPI3L1emBAeypf6oEQvnaVKlmYuyu+s1TR0DYHlaD206zNYtiP7cF
vFf3blLbWsk8u6wnhKTaD6C8j80vCFInNi8IqRcSfE+6wohwXtXYYa0zOVrMyb8kgiwQLJA3uRk7
u2Jmj27XBT146N6KCB+WNP0KWckS0S7rPyLeHGQUUovSN/q1ZU6RueBIxfd/YQ4BZnhqr13/X9Ue
aX+OA2u8HocoXSga4ZxwsSGzkR2Tj0udUoryXWV8GxXdGhOFKCYV4xiyYoXJzmlW5GT1S87zsAZW
g0LP5P7tt7Wp9ZqFxypeXZ7BS0GsfXyqUV5ibMC1YtzR7ZvZQi5rkM+WmeSNKuVa8nwAA0LbbNr4
EHG1C/Ko10SA7gCAvqHicLMVUZwAOm/ZXDjS7gREnEecRfbDCq+lSnPAb8rPIZuZKnE0QZyRoFE7
glxriNAsQCjxCEkI4lci+8GGcE/Vn8Z++SyUgxZKsjpjUZU6k6OKjpQROyOvwpopV/72NRkabc7B
yPmHUeQ06dDiu4y/tGDQRVW+hzZUUWWBW++O6uo1ePGDSTGBDixbHnYnLA3mnLL+tXDKoqycr0ru
KNUQZewEef9upjKOul9rA6mu4bMxqD+57CL5rXl52jXYLDFhB8EfNlKEwNQR9YVaA5s7/GWDdpxk
FUNj2jPD2xTWkSzaVI9aQ+PPBO8Bdqcc71juzXXObFeQ8PYi/rOLJQ2BXBZL3chJcPrKFKFXKEIL
KhVk8o+DKbje47Y3J+iI1w8TXt6CN13EQFrx6wI9ZHLDh5zZEinmkr5y7ILOEOnd5YigGzHWVAVd
3S5qHc2Ep2Ct53NCsd778T11jLWc6WmGf4gNWPl342FNJCBSimqDaa3S6jQhBrvXoJ6cWHIK7v3H
InNDdi7Avt+O0ayaawjeFhk7D9dzUPv2iDXY6/zLLLEovWk7Y6QuQ9e0sNIxg1FBKt6TmUsJqRmf
xl4NNqoj/objC2m1KLrOvf2+ZX/qBRoTryM8NvHHmdt6+Su/+kJT1O5yBf7DcqvJhl2D6iVeZ38z
cXVIvSh2RVi1fngYU3k/vF4z1UGGzLq0G/1TtUSq7nTBEGqZW9Y7XpWTPF8ArUYn9aXWo3ebYkCE
Hh56bCrnRLR90rmjYdWz1e1zLuE1gllzMTONaY1dJ+KjIndONsHRo/gD0GzAC9jvkYwvPGzJ1JOr
nU87b3nRIUsJjJZ1wSChwe7SEjrdQ3s/crxUqKbEXLgdB6+pUqspDWucltLzC5tFn+RMv4w5UR4/
oliJYQCXccxfz0PGxd1qVESMK7TpK6gYSxg4nFr5XLg66na5J0s+4Xu1Ea53DJLrDSxWua41ClNY
TNEw/40wRxOXukDgfA6kmToKGJxq4bQyz3kb5O7lKJu9YLlRVw+YOqvlkIyAha2WbkrmZaDFKj5Q
iIMNrZjGW3vZRuW/iO/b2sPkGKwpLG/2ZvtypuWYSo2Q84esSBMdegwTJEnw1/wVlT6bQVNN9Q2h
5Dzeb7uoOIKh5u8P2whBQKITG/noINQEbA5b3xdbcNaSXsyooYbGJwUEzFgY2osJEXhRzC7xGK2C
ln7cfjUWjfRFCqpOaUxayZ4+vs23CKeOpTODYjgRc48tFaibGkQCZ19kAMrXxf9g/QmrORmbbp5E
JSJwdTunTLdVvmaquzMqEqbzQ9aqdYyKleppi21w6QwZzDLjG+Z4YiISZv0AUVUau6WUgYn1sZs+
BDGqRLo4PakPXW7Q4EwWmSwIYuKlFalH/XIJm7SLKoBj+ii6z05aDVyBYpZYrIA8h/3Vq9RDBX4C
2m0o2sMTzUEgdWYhZT1hRxYPVNziw/1OYpQ4qV0d9uQzcWR+b4Pud4qA/LrhMhqueB+iVACA4PTk
uhpYctNKvaORLH2EJuuzgartX7mfZB8S+S/IDdi3PylIlso6S3VGsOjKrtanjpyMPaDroTck+tcg
GypIG0ScfV4zyA2JddWrUbZA8lcZWM+b+Cp4FF+pvf6FBQg4+zc5kC2LDaFWASziepInnvXxOD6S
FdP7lRc3J1p8octbLcBdS4Pr8eJjbHXdaCFPm66Cpu4x0+Mc8KYNnVQu/la5kXA1QGHRYA4II6i1
PA0MBvr184DqLRF5KDHSX7KVlMa08GbtoTR28R9iLgR3ncn9lqRH3/TrlkMv301rErefL8N4NixG
IYLMdFw+8z2jWdOxjjSVHTZGY9CpI+seriMLGJhQXShBrR4F6hgLiKst5TTbzZmAQb4pzG6MnL1r
zZGAgbOcqmYDwK4GlD6z288oG96H0+fBX79QNVZiK9uWsY2JyZ7hqV5E5Wtv0IezMMe5HQ4JK7Ak
/tLW1SlLPapxluEIkXCKivOSovCRGFQ/xhOG/YrS2+PscSF0S1rHPKfQyLhqgFhpU0eCO3ae/PLt
vSVq2y0eRuU/k4RM384KVTst5rvUqvRmI6/IAeAfVl7sjGIYni+JrFvrC8vUgCtDiVpUN32XAr/Q
INY1TlNm8T6ykOls0MtqinZQi6PBrYKH9lNXRTAZubpSsKbggHRmXl8Pe9PGyOsHSTRKpDyOhdQ0
lzPg42aFg2f5iXobIJfuLaQkoY1bLpJdl/kRABamBipx8uuy8Ue5je7dcs+en9GLx4CS0P2uIfNx
mji5Jrl6FaWvoq4sTS7jU7lYnP6yzdI3gZtB7FhNM2I74Qp59cvr+i194c3xM4HwfKX4erHo6hfz
jpYYu/JApF/2rHVmJRboimubnVMHH2rryY5XBHk43Dq5E8g4selZYyhq32mPxSWCC3+wCDIqztlE
Yw0um2uiAU7zI9ChOHP+xHT5ysT6hiPx3gJ+ibWxICwNtaOSVTqBed/Pn8QFym0xGpupTB/9QRtF
6HzLmkg9uJua9UBzlh5JYorOppDr1smHE3hoVOAjqzaQl1A/LUSmUXcvGZ/XbL7pedeRKMU0pXiI
WJbfIPDmlRbZOHD2g6YW3U1Cd3UzQijM3Hvl8sjchYtMabdMyug0bxqHGzjd3owuigqdHH4EabEy
rzCaMkKWMRtbnokk5/DmkOdt5aPpUfRChbexnXHV0SNaHU2q1E3L8v8VyH0AUAyrndBx9Cq7ynJx
yPqxlyyeUDET5VIhsqYRmQaFVI4Jn4+t0h6pqIKplriNddKVvjFpGlug4SAg3e0FH9We/7cHXS4E
r6StLLWHFBMZVxbZPebTol2leEDRnQz18rIs+JD6qEa2insbWKSnmphHDAtib0qm7v5c7MDznQZk
HP+1EHZ6zZrU6sGtI+FId55YWptBjlpvLz0UEJzLJjuQC03CcQxZkWMt/l2hSRLVmY9qXmHZCNa7
rfTqqcIVKmM3OmBieGwjslDgDH6j4JGHeIjOlblKF+He5PQid8Nuj7XOn4a3w8d91nW4dtBG5bx/
KfUaDAPAwe7v35RsNDtOBSRt1N+g8V4v8/4kV3nA3hWo/qHCBFnXN5fsQzfI+d69AMKJVa7LbEvl
5iq48CKMftlMHk/+wAyrX0RoO41GQkSFXVQ5aMIYA8KNBPKvih8iw3TT2HVuqUeHfslFedb+Bm1A
q6+28wMZourtHTmCQM4l08VGtRmsxRqis45Qz/nIMFJmzdeQT/n9amV34mtCWBgThEhz2pkmMjg6
iZeCwz/mLpxnf+EV7Bpg7tyzXoS0oAlZ0owU09V/CLtJy2h1gMG29H4Hlpsz3IJ3idYdqMdIrc6x
5/Mnw7ZKDaBiiMEvKCPXBz3cLSLZbuxE+hfz5QRgVsZCWwHvmBlhl1gIy4hbi7eVM4b22MSx1Auc
vUS2SgP5RKhu450TI8NSVjmMTnpF6cuMVzV2OqR5PjBhcPPqTEdMGCOYC+ehaJYL15heXK8gb4j/
MXzQmwC4uc45JBcq0zlTvT3Rdg1JYdGB57cEHRptf7QG+AdvnaZyZZKtjgcxp/GunuJjO+CoYN47
TrdE46sBCySz2i1ZwBmmymZI8bAOLq0D3XbVZXIyQTR+M2Yz8hnDlFUU7ZC0RrvQrslYQmanK4Tq
v9ijuDVH32KD94ajFJdV8vsYrBTXMAyRSpioPHF4e/rWmFq0YsVFMEyiwiOXqRHo2IuqQaYv3WkN
raMn5WSf0FpByQMH+oxHXAbUMxb0nv/dJyOgB0m7qf8txwTEzu5UZRtNqXacB+/oINlEQJELFy7O
77nzQ/Yu0tSDgONpEjHYLGn/wulFTuLm1h3qa+2tblmLZK+hKtk2deNcszBbYOpfxgJeYXVA5QTG
IFjYl3IwYjQfCSh2nQTtjGPRndyaljylumObHS+D0mJdpQ1cF5f1aNQpe9154MnaAWqQq2domg6a
fhOc1lCynmFw+gVoyR9eEf1vOZ94lKJKmC3Y70jLguOfM4mSMS0dl/ZDPTDuisWGSkJFufLyS6XA
DABWm3wO80v/au7hsfxPkfpnkvkys3SmN5Lkb2F+db1aNbJEij7yXQL04ab7whzZLDvCQfewBsAx
bORdSmUKH2kq7y4OZTXCAYmEvtjbj13lA3iKVfC2fUVZvZu5kIrXpz/lK7VY5WwGcEWX2AHbuaAU
HMXlcspIQ0bGeJc9aAGvZTDPweQwf7pZJfw6b6r0eabvhg+NKL2sd/yevt/JNSG0/qkJW4cf9kY/
d+jGJj5thEE7XKwNZGGrbIDrjx4FHN6yh2Sdtrg2Tb6OvvhQZT9OZEmWQKHbYX3eX+i01aRt1F8W
HV1PKqdnEYDzgkCjisA2/mh62fQMlFL+rhwN5IvZ7j48jg3HKQgfNY/Z8T9CNYbezHHle/BENeVP
T5kOwW2K4LU8uK2w5uEsvSMyPHOZHe31LThpX6k70pTw0vwwrrDyMlFgllPdnN9acRIv8ODuldkL
3bLCR4CqRmnqGKfCRykoCKCkOmp/Wlnh6X87pxm1vYTO/irPgmziiRyEHANtYaqGp7lXLXRCy6nD
6tgp6uiqcZlT6Ch8h+c0mzLAOuARP7jBf0FOsRTrUek5PsBFRTVETJho+gYUHbKADcKy33DNPq/e
xUHo/cybpVWUPAMcE7+Wkn0zaNbCJwsRcX01iSFDape9EOMr06l7bo4WJtAKiEg8mFg8a1oaP5v8
5xltn4EkYY55zMGvtzbgRYMcxeU2t8dqc2tP5YfFLBcU8hSA9JnaGn0FZbCAccGNVtsUQWqRqPLI
2F9kMfRp1o9hXxqBjXhFbD5BmJopwk6RsueAH6ALp03T5Pw8ZhlKdwCWbBOHUMMAxDXRYhh2WaVQ
FHyDjDnG4AdIKSWHiWVxTXb5Z/bmGhbhNXDTvha1GPRQRcTN5pxId5eMi0m2wHYjfI6+aYZiXQk9
frZlhBfXx39a/V2VfifrvBQV6ndv76MtvvBv8AWqG1OpwjxLSUIDBqtDlZMuFWoRx/EHIjK8mqci
diEooOi05JSp7p+ZVABTdH9KuwC78sAWdHAlSAMa16MbInSbEe0q7auUwTGUkH/T5+KVEmypOAw/
ErRMLEifdu2FvNQNlGOzkrbFR33RBU+XiXIg+q2HHL5VgvIHAwvKvts1KLQl6vEXRD1Gim5B1Ap5
/4fDFIiO3bVn/OKnbBgiOAL223woTjA4X+gJ1h61hTWhnSBpfHRXw7TUa8mUTQ+tSDPHVAyG/afH
VYbTQZfzbjJie1ir+/dJv4uUEVC2hXlpRsrl2Tr37xLSmlrQKljJ5d9BJFqqM0fs4qpft8HlrMh8
qek6Lk2Wz/smaXHx3vUYdGxmmV8/bHLxOewMKtXwpFb/Yb3eFu77KVnkuOX2YjSZcQhst3beYwgH
kVTPmCZiHwhcnUKtigxXQ31nXjGIuuUp3MnhkvcGSfPaN53jGRVJtm4EQw5xUN3vGmfnpaLTVxNa
qD+csyVGEaZgBA6bDK3plL2YwRDFzC+BGWt/Kb3m0Y4KLXEqRW+u5QLo1H7YL+KMiB0JYA+PrKPz
AMH24UHpLcg4xB3wVhO95BSosnwjdAgedB9U7xLFDXOfdULdVcZcMKWF5sZU970CZ0bGkqkILbw3
Y6xG3sEBQvAapWpjlu0t+bFFs6G9R1YIHNsWCrlbITBcTtLnTQDXjOX5zr0SU0TUJg7MZKYnlHsM
woHNW7IFh+RDiTB6ZvudILW8SIgbw+2IGDwUweYFttvf+xfcnxhelpEPq8kdowehC3XaimVkepyo
zyzjboJtT+6mxQA2logHeBggTJec1b03IPXdLRbyN5+g2kh35c+vpY3vC3HY9nTiI0raichz1RYt
S0RrwSO1Fq5EjswZWpDEnokERWvW9W0WTPZEYuYCuR+DC4R2fPkXx+BXl+948LKycOEComdOdkdl
4qnjWfUTlyV6tD01PMMdfTa5y/3OnxVG338Rvn/DAmw47lIIVzeBBHSoXg7TmSjCXbhacPrnBIie
zKL2yRsG+xugN6yg4lyVvNr5+JU9mRDilX4ngv6PwcQIxK//k97KXlWo/ziovVFgT1IMBnDQi39P
lEUXIFuSsWx1kuNf08GiY5wKY4G5+XCQ0tbTgIw+GQ2eA09Ue7YNSWNLAIqmwlk0gkq1bvYuzTwT
dqqNflhhchgyG3IPFrmdFygpvMi/0HNkaHx45e0ZyAkpEdDoRdONQ52LPLIVqGgi0HxwOSHXPit2
49NLYmAAjsRA8RZYJ5Ma7tcOgXzgCqweXOtIdTsbuZM+LZIiAOIyPXrUOaSPmNEndUM9G3Yo+Ta+
LoC0uTcrCscPNd8SS60xt73uwVWTYy23MI5JYgiHSmVr7pLEkqtUdaEXUPAreY5eFt5fOsbgl6sv
lVEwHN45IU+Lf70KjrQmgLDrqTxlhB1cUPKkQ4OUbFihcrO3A5OBjs0G2EOAbz5kRtfg6Xn9+Qyx
yZjLM42pwufu+MvYa2vHiKasZQrKBgagc2Ik7EE6WEcqfW5gUaHnV8dY8rEDld51ZJRTi3l2C8sT
qdrxr3Efkn2G2viY/gGnX4rQybjwviGC6vsEzXTNgjE672Tnvs2fmI1c+xkPOXRvkNm8cCLxvwWZ
6U1wl+qVEQtZnT5Ot7K7AIII4+VH76m4KinGVC4wq1gsInb6JC4pSjKj5E4GjrJc5IrnqvHbu0v1
S2/DFBymhOR58j6fvE18x1bYD76SpCBMk+0p+R+8bjfds+3sr5QDdWtgYDMHEvtxDUKSdag8qhLT
ZpZTui8zaVdb5jhJS1kRahex/GvdgTg3jWZnE+IdtPkTqjn/49IOX3U6Fv6bH3O9/r+ElH6A9unV
kxCpAP6O2uQtFErVVrUQ0K4kzb+bLIIsoOCjeyh5BJDZ6XQG9YeFl2voR0fVlJ7d6kabJ310+auy
8W1NNuKEq0iagtXQe1WipknbivKx17mWLMm//gchByibSETvzqwMaAZXVP3Uv3XCOsHi/N9nREr7
+UOMXoE4z6cQGdWuTbAR5K1Z8TAp+4Lym6Ovq164vI8cYl6GTCvV5OTb12bUIv+8KGlpNQkPSai4
s7dnWHRIVdaz45/uDeOfnpB2gzyHC+OUWIhQwcvVB30Xt+g3KLI6WivxfCklv4vGVqvBSwQQn0t4
6BQpcV9G/oEdekIvdiaNHTjy3BdZIppQsySVYpM0u7ZI99GUv/bU/KtFWvUROkkm9INZcRtu6kFx
s3uLhfF/bGvYx3xKuaFM5T4g57lwW3Y55oEJDookfPavQoDVSBBm5GQodtmcHocF/uuHdEArcCpv
rPrE10bledg6xx9la96Lrg7sH2yK2AQwMh1Vcw5t+VJ/oCBd6MLt9mZfHsZBgsbwP+reLzE/68WL
YmqkdsPMyVzVoiHPwZZVyoqeWmZYtrd2frMzF7B8ruuQzagM/Iu37O4+LmhgVX0wu8zsovBmx+kB
JAMMK6aJcCWRU2+3IDyHlsmLGNqW5HDWkc1o4IAXuj/RuyRR7up6T/WL9boshoEI6f+QSl+QGcOc
tiGNUp48uYlgGkLFKKTM26EyThn9YYcZGucEToswZAaCUMNYj0/9xW5wgtrwUzhxSTgBjHBg1enk
a9hgOzbR2W8mGWxnqlnu5dWDtr3lXnZTCCuNgsTXOQw9bqpsWDwh7HL9P6YKGc1ODWxXIVCc9eg5
0ZWfg4D7OMgicOMf8Vch3hqrrcL8d2bF9DcHvcA1zV1AARNQZJwaEG+2AkfzOGpZB4P3o7kjOHCW
id6+W8YhlSHMbP+hNF9byt2dPWhN+yRC97XzAVh7sQiPYE4lT3Yw+D6PKNFe8HGKwM0OaiZCZheS
3BOkkpeVbJmlPRLSbvTS3H1eSHMF3QxsKsQENDvjXXk1TYFfD9k0uoyAs+J46nhne5EptAuLp+6n
EUpJRPJQMrK6dydcEVRbr6hdHp6jVmKfyzwz+uJNDSSmm9i8/q6zKNwIiOVrzECJsmsMxmRlfuUc
7os0GqcZ5rooaPJ/DEF9SckU3l88QkiLVZPw3tqhLE7wtAozOG4pyBi7WjSCizczDj0swj/s4ShY
rrOPxmVanQQhlEP8MWNSWXBbH5a/DPvLLesJqYiYP091xzUgVZmDGKnXwLqxsXbq/Yhfii2kQ1jq
PU+TlS/bmI9yKiXAe86RlG6eF0BZG+tw0jce5zHWoP6oQvWo4UPhuuyVMzaazBPNiyZGtt4jaK0H
OE70HeCyStSXL/yXQayoOnqm+8wvYNBculIl+iiQ2fPgSUnVrPaWYSf0IxnACgYhA+d3l83fh7ZV
iQoL8jfP3pyYVAqcGpjy/UVdpI5MCLZ4p6+K7yGdtrJl4N+GZRDH1B3GYd5RlbHGiSV7xuOPwiiV
HYOOA5tnc+RRT45fZPHbzkA10cGZOzyHL6wbP5e3NWv9bv04OZgPLpheqat9kO2HhLVWF1j5NSGY
c6BtKlD8AJjKznsnmIvkRUThsRcFYJPH8BSI0Hkf9spZV5wsOXM68/Fz7SDy71as27vkoE4my270
ZAkFsk8xWeH9MRpzShW32P3yxepeiudBQNgtou9TsA8vomKeP26VgMSmftkRVs04DufL2bYYXLxe
yILMOA4Q1MkFNnz1NlEwxeKQyeS6OoX196H412qMPafIPClfxGmYopKLT7TIT7mUskLKHfupxLDi
yQUp9E6fYT5rRLvnLM4vbDKFlDlXW58Sp8MTciSa0QYxlGY4MhV9SOXEaN46Opk2Q9V32izI3V30
tJ9TIi9UADbrDo875ZE2o5vuOOxxP/E62gfCOm2ZN+ziSAKwFOOI2YhNJhilyrDvJYbDAiKTjUza
g6+BmX5+LHTl9sRhzT8J0HCtg+e10jBNwerZBLwOsWmRNUGbrd2050H8gTED2uLPfKX1eVUmAnFz
oG3EJ0xiy65ux3M7l1fkgCujwNsHPYU3syBVLsqmCdNDn5aBNGeDmaHGPeaHc446PUdEz6skPzek
4X36yhFhWxE1aZtDll4RHCHf0i38OQ+loPHDXH+zpf5JsQlBlPwNkZtnQOlwEwWkEwI7kRrI3t6/
HIjaj/Zl3CpNlnGyQZzK21EwWd4yMYHJlgcoUPeWbyeR8v2w0XQeVVP6DK+mKEx9XakKiSLNwdtP
7SWmhsi3j7VEhVMHnuHdalKbKAuY7gD67bpbRox06GhgbTOrwIBXxnNOKC+rVKtsFvXAgRhEVSrA
6St3MS4bVwGVqaeFuJ9T/Ufr9M95HSsI7LBFjg8RLajhWm1rCwRYiKsl+HCM1w7CH6GceGxN2zHg
Ab5qLucPEgBfhmRWn7Kpaq4KpcewtEhmI7WzTgGMYb5pX73cJXEA6a4qQIxeHYkV7Fb7UTZN0gRo
nBZomgXEV4ug16Mz/yDEK2Ugg7ZCzCjoAnmVObQi/0pYa3GmKbQax7155+KUH6y3a58nOmOwdYC1
w37wDJKO7rqAEP8WtUbpZNLZmgVoHqcgcVG5NkzipnP0rLUAc3OMr2sxw3w9nsimkORpabCOjEnA
gk+cl8s0WIDIUqcEwXl77kseUirsz+izLFIIyEoZQJzby0mdUaaPineeaQb9W2CAwHHKjpjkSd54
DiXpGXvH8h1OB7XJ0NSWdCozsFCXLbpQXUefq8WmIZx0gWNJoCz1lSSU1UFVjIBXEEmcBDvuAkt5
+P35eYuiaX5aXtDM4K70W/og3htlOvyj3U7nRQ8m0nIaPH/ynqIkrA5wSrl8GZNCgaGArIOrf6/B
DbDIdW7hxUzVgdQ16looBEJmvKuGZyW970SUVZ82L106bp8l0AejLJ2FEJNWjrPeTSLB9OLGaubg
a258oHXa7g0f3pqDMe5f6OF5bdiXrr/TqlMDquxiD1cHxnhCowqxe6o8WfLG9QyZgBg8+VRwab3d
DOPAC14RubfkOEzikR2kqIX0kFBddnP8qBRd39zRGBWVxqLeqM1vaP2/DtKn/xeEubA5iLUxSuQx
OLlp+h5i1XnGAFWNEwqbK4JjrblFqPKOemINfdlYXiPyAlEEAns6CesSLqj83jAo+PHQNleEaZLw
2FvCKn3xpSuCZ06xuL/JaupilfKVnouU/xFOqO/XjQrYadneECVHByp0n7cxGtgOIlWEFAhLZUPr
dl7ZwZ/402r0bMZzNX+N3pUNRvdkX+aWXXM6d2OCCMRwluXSEoANH5TILRL+nJgOkmonbp/QUIJ5
q7qPAboO9VOQtLiF/dNUDKMGN/7YkmR/7A9QHe39zycefUpn7YYZC0aIrCO0G30hLj1M0teNppHT
an60UGIIsAiPcAafp3sJfuaaZg+DvC6qh12p0Dm9v3naboh2SobUa2sUce8tsUvGdaUe07AW22pK
M4sUE9zx/E4bS4akcYLItMcMUjME61icp6r/g2lxc2doqLrhraXkq6RqpguUgKAFeL3UI21FyaaM
+AbaxqjoqAIcYPhKUbFMgwS1gC0RjagM+kTo0upppA9A3+Nawc8JLEJFwam1VVUd/qECn4xuNbW+
keKWteMTb4pFF6KPULK20Wn6QJf5keHuxSiP8DtPNUbVFqugInWSjkJS9JeG0Aix85frEBnMf+Fh
6XTO2pMiC9PGgGFVPG1p9biIIonFL1vhgegc281Hv7iJ+1XxEpryLBBIRexk5w6GXT017aZnuTI5
LTZ8OzR5/w716bdS5nhCxMiaWcheLnid0ifYh78Vl9K5//u8ebjQkkVPwPTp6NHsvqIxC8AG7RmX
B3ksIgJWLsEbHz73KDvN6URg2inzI/UgjCwK7NJtfUv0wOJuToY+Ik+3t3E0eQRRAeTtDAWVftMq
DA4kVAX7cQ1BCUagNtRkhKa9Hl+5GI+0AtvMZd6bYdagleSjUBdl1Tv+xcsOdBETtL+XV4nwfvIO
NXx8EvlEBN/Pcv4QwleNnemGwW2IRo74KsMVQ/sZVLrC2/x5FPtBvd/aS2oNlMLzOY+zOSu6MAFY
Qqptg7t7ynwd19nP+dcq0svNEsic+PWc5Wny4HldJdt3oOOCWNIZuJNxmf24PmURw09gTF5Ee1Xc
oYzHYVOLU+3eu0HNkwrEa6Pqtfa6TiiAEKLjem1ZqpvLElAhOtmYi1s3ROGDhwgIHLDKECeLFxrG
jk4QQIUBcpFIOF8WvfWnJ/vrVLrSIaxhWJqLM929dLu8YT+YfbtVDntkH0nxyFijlk/DsFsKK5BN
2UHh0ZlKG0pyQzKh3dLvb8yV/Y6TdmGbGHF1L8uGpcXOvbXVOs2Trng4RwUwvhKEVqDDRK3134dp
qCyFQPXF7v/xkeSda2G/GdE1Dy7OuA89g444pxAT0Oxc3hDQ7qvOZVkfcIdwSN1vJdmUHE1Iz0fW
wueasZzirFpPBuK5yOSBq500X3jhbNasSyNtQ5cHzkcGB2la4v+GWQMI7dbWgb/ly7VoTW0kclyJ
7iTrhBYrKW1yY02QWiVdwiI7nhc3vf8yoKAlF/LuR/7kWsQpnsu/HEa4Tc4Ter7atIOmLO/qBQww
eOtVM3JsKniCkKICj7pJ1Z+zlLb1u5c1OhbHS+jU6f90k3Gq/e8KPi3kIDu+IrcJAKVc1ANKlh+l
4Au3YelidV8MBS9lkrN+Adg7nypGNmlaOjClz6DqfIb72VNS4tKxB2A/G3uFAHxUn1ufQxUzDEdH
hraWD05sq8u7NRVRRUdr5LgMkKOkVxD2kxujGwW8J/jWiNs3GvyizzjpQEcuhp2pDl3dJ/NPcGNC
q45o38wZQqKrmKYDczAR2rhLYuCnkgyLTar09MBwi54LiMJ76jQSw9s9np3Jh+3BG9J5XqjPD0Dv
q9OcdVb1C1Q5TOZbAmzIIekSgLJKzR+2GjTUN+/SmBnbI50gEnXqNsBMRRr+4Ngky8ZJeSSzBTZH
0Ngms7Q3hKIlXjJRpCuSLYmQjE7xdlEo6pRXSW0me1UCCthS4QZAsADXepyLTTjN9Pk2ju98+4GE
1aRiwF+RNkrqK2fl+xvYyFyfv5B7y1pRZYUhJxKTPEBwExpHAqoTf+KMI4vUS3e/DG3nvM13JIye
p8lUIms5AkikRdH9bZSaGd0h2agHg8yyiz8FG89PGiaLOZbIaP/mF/p5OqtipZas7djCSMh2Alwn
2m1j1rf2OliDh08vw2yQSV+cMPUjk3mfhiTF+w0+UmNVDWN1sI9vZvLYy0OH7EOxVDPZVhg19kXa
gSiB0lWx8+Ur8FKZnKjyPIeFphrXAo2fN1AurUct1OQ/d6BhYRiGdNGS+cnOsLkqymNUwyDzmhNn
4zxMiNDhvht57DxynKxbxxdWQ45qrcH2O6Ip9cwYx8VaBymMkuQe/G8eWl3Fle6hlgknVtm0p87L
Gc/WNE/ryTcTRcfma84ggP8M/3UV4DZfANxHFekUAk/P5gaVpzjBM/8lIdlICd3TuMZStJCaG0iZ
840NQ3nY1JcZ5j5uY/KKdzpCm/U3UL7RLA9SrWuxRPeDw0NQISr4Wlan55QUhKVU55xr4T9UyBto
C4i5OLwNlKVpkVxZrIjLide7tFyrK5ssSgexYXrXkv8LPMyskFW5erDdU6oQ4Pj0c+jGu7SddWoZ
806Vo2pWS/wvMyXg4d3JxHTHoUmNNxPaPLoSuQx6jwNhUDhX4op8/x/YUSxkAwanb5BABNAdR6JM
7ieDQ6Yfkn6drzODUpg+AN43DIqdVBS/SgHIJBJSAbA/uh93C2xFVDoIDUfR7/Ubfe6UYBlIczSQ
KaRpNQ0yIzRefZiS03I1Brark0PMfghgcutzy+SD2q3zBOdDLFDLP15cEykImrYyx30uMOxlcovr
8e63MRsRAyCZSCEVus5pfeN+0DMvFgHAZdcybFsF1bh/r6c9BUqWgbuBUXaRu/abLsO9rVCw22vu
z3mV4zfzWmG4nH3KNA86Di33ANRi3pUo8Y0oIJ54owVAomrh8lpkjhbaSUwUgiC6qCNgxCQ7eqms
5vOUpK5Z/YBhaKy1KiQXSlMt8LbKjT5daVu4yUXgDTahptOVgnwsDT22hMQPS/ZivZcDX/Hi+vX1
3f4/B/FSjeNC7H2U0uyJo6j3j3biQs/hjDKMdmuvomh/x+rvjLxdpkQI3Rm8WULFV1MG4Gud/KZf
/uUZPqpyn8kCquTED3lhQvJAdtnyjUaDNmT82n2Ef0r/eN7Pl0OXCq9mGD/XPEA589bq8wW/fMbi
oxkF/Q3rTUkyxFTYKEwpXG8ohT6z4pgMxFKB9rsAGmF6JdnsVHbQkK0Bn9wojZBlyVyAPXcvIZw/
sK4RiBCeROwMY/l/IXrdX7zfQzgwr2kNM57F/DEwE8AvTJgUGHYpIKhpvN9sN7g/oKXE0yD6Cj2V
TLdYsXNw8z4j++ONDJTezLULno5lx9NjC449p0QHST6h2lnQEeWfCwXVDhjzVgFF/bSheH4k3fDE
vaPNbnxauDmlsK8zxTS2wjZlg2SsvWLCbz51RxEjjl5/zGalGzGLuZ3eNfHI7CJqXsIhNk8pR4BO
EHB5tdKDoxu0LPuUBpt3mMYQ3Mv/hey1CPiWbOvDYoC1i6zNC2RI62FLSyJDE8rt33im4/7DbxRE
1PB8oNVY2XvPKjAPS9RI4sQRyxRGswt9I2MJo9iZbB1b1J13GEq1cgiqkoSf7g2MMKsxf61IBYnN
Qqd58OzR+N9+P+p+COoaUurizz2SAgSTSXEeYa3bIGdi7NFjubWXksTULNsJe+aRjDZYQO/Cl4VP
6wbjMJy420UVXZlgK5tAG7ENJl2zDGjeeFsd6Ha9fZKIUknJn0LvLnHIC6dv1vnT+3I2OShrPVN8
EXT1dIyvT8tlAKCgtnE23KV36INwzZEPKNLC5xe5Hpn8nMtjfewRKVnAoPksh481NZ0n9OKaJBq0
LA3GzMu68kIs/1u6WLjkSWXPrDk+cVQCedz2pRuN1RZ8IMtSRq3wxwhdhu0aOXosnNyAJvYTDAGe
XjG+TLaODnMa16R2hs9w81BAPUq9ArzQynH4Lz7P1y5skz9QDDh1RTACpYAqR2UR7pkzP3KVB2Kg
0AVRYUz0jKf16lKKHiEbDWUzBuWxovhmlGKnlP/chwbTneEtOJuki/MiZtmUdkDBeEku30KiNgpZ
0UwO2Y9V2neEJzqF+wiWa/TI+odfMaVPRT5ctaWvOs+lGJztOMRqLX2yGQmIfhSD8RHAmjZHv/5G
gjVcjOZVNHdans++acwpSREtuDDu/GgN+Owi9ag5YfNlHgcqe9xEF+Z/gQ00kVvAcZjpj8k2/keu
FH/Du7qWLWrehPd2eqQ1Nq6681vTTk/IW5M2AP5hOVW+1PUZBwEjon9uuZfKsMeQktlriApBxwiw
UeHPCUeXuLnK3q74ek3AqX9B7Vve8YgKWtLmr5tS9rs1QiEyTwm3EDDzWPPmoCJSV4RWi+UGruMY
oZOnTdXT2A0Pjab9iA2zWMOFKP1aNLIflakWGAh4813LaiA9xl4Gjjz+g9ncm3u3TdWK4bI611nj
V5QMXGaDkaxrpHzTU1RZFzAQ0o1hVsAwCfWFOGVDQGmtt/OF6KedAzUD7C+7NNQTsnQlytFc/Yxt
9WLDB/xOyPPk1i2Ud443lugE/9sEJnYEhResbEnwxcg7VquWHgsyW9xSwyFEQNVhNxq7OCFuzhf3
6yVNpJuhzttJOhpnk2zHMl/akNX+2jfEv6cqEuKQ9E2YndOoAJfjPT0p6V9RwBF8EA9i5B70NQIN
f0XxN/vqJHHsBU5vuZ8cYscm1J01AwfghczS8XmZhT1BBb1E3ZLCnDgg8DFbE7PefKAaoo1pblDY
HitcBdaR/r2lmQViDSdaQe2Ej82Rn/NHGsHebY4BtmuYLCQLnrEGSFhVZg4YqKJss1H1FFQi3/6c
OLoCGbB8cFqnOepqq9lbj2U8FRhxCXohLEzPsxxDQZkdEIwHkC2Ynx9rt93HU4LhXg6vIuXTo/v0
SF3GSZdCj90LovYI70VOEKHecW1qvXBsqSV0kFPM9cCohprsdLvo/BHPaB51l69lAOB8Hi8lxqm3
t4IFwafJjebcqQCF9B1bhanBa7vcoAyAF62ZrAbedJCFJZtKr96txwYluq8A1MDHNfVzs+lmvr+1
VDlF9fH4/Vs8epj8Rec14WVMVdObesYbRDDUs79THtbP2cJG36cAv36dzU6xhKbMaXjfo//dHeVU
ned8xVQm/Z3b/nub7U6dOW7/cDEB1X+wO3MXvQMDsB2a9aqB1e0YO/1Se0+7B4FhLtZqR5e6FmfQ
LYr5WQtA34vR8XLk1tZyWRbA58rQGC+N5D35VH2TwbtQ7qhbTCP9jbSx5or39A25xsxo0TUkaFrD
VUovP+UofE6sXGNCIvMzeLmRtA/Vpi6TolYfld5H+yJViMAtjqiuMMd4Z7YElpaqk4RLZ2Td82WL
VAU9T03vCyu8+yvPpIDnvrHGRoH8ymVQHgZMn1qs0rlL4c5yxlZT8hMLxwrSR29t0NUi4ZU4Orss
T7xRsmxlcrczzNORYlbrbozZeuVj6/90EkJVjDbOyU9lgsX1HTSsGkQZ8INRFuLV7YJJFicNyGM7
1c6ItV5ofRX+LvrvhyNr5Xl4GiLVDetwP78WQ7Jy0xA4sqkw8Ow9QxBqMU2/Mrs6QpqtD9KmguEs
zj5zu0RcM4qDfG5+mOjHDYD9maLqmmiAxptbBnd1EpcrQo88K6IfEEdL376/8MqzEaGhOJCJDJ7/
1KfjG9kaDV0e0A2YzCsgbSXJVrjPb5M1MMRqg8z/GoM4bAzebvByIBjSVLUFYau2VDb55ATeKOh/
g57V1y7keUwcKaHuH7xgO7nN4WS/KGwnk5NjcFbm5j8MU89wWrp5Dt9yreBwY0ouTm/9RFd4mCEq
SQm7pWSpQZNLXYm3o20IvarWw6i8dcT4gOz96KGkvaLB/C89Lcgb50CIeSQyYI2oyltWonPunoZI
YQiz0zSRLK/KdKmkPWpVcnZXG1b7F4gGDFiCL0AJrxSZCUfdGu9rkH9cTUYpKah+DKqjCDO5Z8if
GcnXgSTtcNarGF/zB7tD8eXGjxCNkLKaFUCFJmLMknxfVtfJlL3Nrjvzn67sG1o4pzm+N1TQX7TL
CnPP5/KCb8HbRywYPyxazY4WTUkJ7Ok2D6Elc7MhrMTnH2TDDjFF97lfVOrIIQzdh8EjJWVk8bio
sdjaUa38TQRHOvH2fK7NZ7/FhZtMa5jOqqALSJsmdX5AT3iZ746MGdQ0z7D8a5OAWUgpCBrLjlUo
lnpHcrZy/cYEE5plIRajNbDBRzkKv8MNq5lHx9vf1r8e8OTh7KNDH41ZHcYpslhkd5eaptvSLGK6
tBu5UyteFbIbfMCP3/XfiG3udY29ApVgxi4OibI6mOllXs65I3e+bzkd00tHPLsDT5XCoCZgTwJk
VSdjTyhoa0i/+K/vP/4fh8XlnkEdeiif2ki3zaH24N4LBSRjYQumcSgOS4It7qrpe9X4XkqVdEyw
qyac5IElGUJf5UCbW/wsgUoNuJFM+bXDPWATYMCDIRAZiv5N+Emnd2LXQ++z1g+RoJldR2paj2Y7
e193mFGOY67xS61U+yCQwhoGiHMHW6ffyDmwGdxsdD++G4Q2WbkV8v8Rl4RYpapMxWGgKWHzqlyC
nHQ6Wsvs0U71v21NozQkyg/jS8gXrQL++YKJ1NDiTHSXv2muRQz3rPszKOQXYAhRQn2FeuIMf94s
GZCN8uBJW6YhejZv5+S1qCIDSq1B9AHLhEou3gO9Lkko3qDnT8Etlh1UG/mcoHK6us0kgH1r5hkH
TzcLiTgB5b+XoqCjKz6Ai8fsTW5nmqlEx9dN3qdZLNO6WDisxb1U877tvkAlTW9WQhFMtgchaHtc
P3gih2AZFa02mGF3frACoFP3uvgTwhFr5LXB6wxkSOy5hn1BOFroxDrFgR7CByL7gvfljHlkuXos
ckjlg2zGeIbDEIMoEbeIpHj1RwUbxCwH9GyEVik4qWrJHGlA9ALCt2n630KBmV+i7iMtSIoIJb4m
afPftNinRRzkpPtqwqy6bynkPDRa037DiBWdXVpDcluc1sdRfe1kbh+OPNGj92FWPpcesYRASB00
fWUpJN6i3PbeCBSzhesqu2u1JMMHl9TvXRBqk3B3ColOEAJeScIu7WGIm8x26WgoAiGNxzi5x53j
8e3tRc7BDNb7Bhblti701l7tM0Atc4DeQ9GQ/R1iItf5qCleAVeqBJ+4Bm+KefJWKHjqFOb9RQId
gTEwqJDRX/33ZEZrXIR+t+ZBi8dMsi7D6bSZwZF8CUXFIgXG3YdFQBdcD2h/30oAZBPR9V3sXg0o
htgG0QQua21b0pD5XL4DAvxv9Bb1aQiSMgTwcHcOh8uKGlSX02yu/2Zn8P0v0hGQi1pHvyZT+rRB
kbHDx7zqYOw6/hBOQVJa35NIiFLiQhhyGAjDUOGADinVprjiSLWQnDjYZlbq9uaQJ0+bnixHG24z
lH6Y9k5ZWBi2zkOLxSKnVmembJH1syWdE3Vcw1j4VZQrcRLcMlBQhbXhB0z8cedNU6kGSzwKJCC+
mOkvNV2LX+33MdI8PfgM9KxqWjiQxicYuuynfx+AkRb9B5ZfIRA9yuACwPpVCzA4OQ7BeHFGr3+y
Cxfak8TLSqnusA49kPvnt0lSMf88goSjyzvtRBbPQg4lLMgoJhcuOflbGFonjmtBOgONX3dxwy1R
VbWFzOwM7WDUP0cX5ftp2H28tXxmjf7cy6WRSCiLhizBCGubaG4OumXTJ8bcKdc3/MDKMHVL+DQy
5iRUI8F8kT4KgxA2ilWygtZMo1zQzTCornKbYmvCPbm+++wY3gmqUqhBTGf8zjeOnpbfq2NRB3Wt
oWt/2UeVjDupqPNGpaCnJqXu5m6df/89gP8vzfDqLsHSSYXQhMd1eU0MEzRIQcP3FpdoehxbY/II
gDf+ZH7WlcPoxtJjI2GJTkMD1U/jY1/Ry+BFqPjx/uqrLbMu4haiOKJbx6CDiu/ACPAsreGwKiRl
cqV+H2wjZe2UAXuugYfZ+3uh2/35u77bG2+qWLty4Ie6NKG8RiukY0avcggDwBSgCZcXF4AGcRpn
2R82EDzyWl09z8FRYOZ1uuDeumDvpcYVsL3DCKEfYtxefVig6YeAqueAsnOAxUGRIieGQtaU2K24
3NMoCTxzYCVqWOq//sj/gkbd6blfN1g27WCCTcQQyLrqcZWmmNIS7y4vNwZvEq32uVoyYyUUM10w
lOMY7TJGmb4p4lHO6fHd9waDaJB7CmSjLSyQxNfA62bASWdaNdcqcVd67vAElxubVLfLgVA1kdlK
h7NZE/xL3uFZ6t9iPFWnHy+GPSpOQ+uKmN7eEpzXBGq3CyeoRbP6RePCTYszRFyEnonIq7+sdbJx
AMQiENqTJxXWZiWSiXHZD7l0TLDY/CoFDqkIGQxWj1X33q1MCHm41bNukHSpJcsGCDP0XoiKjzv6
GQiWME7XKxiWjyJLuAPYilixQWcF3ZyRh5H2s9CRVY0SKxZ2559/G3ymk+Icn5E7o6hmtMfOOSWS
57ijYPPlxUwRBM3498H+TR6QLzltKK9/3NGP5TkVv1uphiKED2+n5wqbXNcaboEUs8J7LVSUnPFR
RCNEoj9GhYb5iCx5yMGvUsPp94GMfhgwix6EWhmzLKoBbEcaikL8LVvcyR78/jm3mI2gxAv8U/TL
7ClWS4kG2Bst8b7zYgSWpz2T5mCZAtMerxx+04AsX4CY1L/DCysJLsQd40DSkZkG25IX06d3dCBu
uhe8VwGafrsBJxdaDLk+eWQLUqNMBJQQJCqxUJgoFSZHm5L319s7S2DkRGh+9/CB3jUcE+HmowgV
CIxwBo6hu2zQ6bfAYZETexeRWlu70GKfnOxiLjTuv9oEheFBKG/qAUNtU/DvgjMEg6E5u5vX1kFi
2gAXauaIi0TThvLp1QZBZQn0sLFiy5Uqx6XvEBn4WCTSIYWdz541uDhU6PcSw4FqjFLoS5lmp83z
cUkKJt0M7oAO3WzOmI+AjOsLR6QmKYbTlVIFL0U08S0a6dDWydOQgpKrWry0T6OdE2CgMBzQJuyH
kGVN3VAMm0ZmKNLbFnipWVb0P28ez17a+StC880bn7hZhhxR9Q+n5yR3eisyqtEEggTJLRUhPJjz
ypHcI68iS77yrgXJAoz27STFtj+PwNMoRof2EzFVUKgJh3FL5cBVZ4RQrS4a/OcASZTnEsw48UNy
1bpu2Ow14w5Vm6Mgrzv1XOftd8UdLyFzPy50Su25YNeIZSIjNkwVtkA2+HCJOYcm20C/eYeTvo1g
Fu5J84HL1eXttBgREyTipeTO7J8Ul9ij3pgcuo279LRnKYdj2sFE2Af8MjOIR8lILL7DUYZ9qPNM
JYJCML76/wtdfv5IYsl57yDPhSyQf2T7FJKwOEJ9he1lu5BLHPF+TKkH3yU/hy+wJVPRJg4ATVpY
06+HMhGN+udpFWOX0zLzJ0rXJO1OR6OHwelllG4I0090EtsioaHZVbcL54UxYPPFMhONeSaijUNA
+oxvk3nBDZv/NC4YWSlWrwzl3yMnQOqXO2McqPSdySC4mEcYznLvbgJ3j4U6ptntAHThc/Vq819l
ZnYR/KG4sqnqtvsUmEwPOW/yD0ZupGsHpwsIXYD96lVXhAkvaKya5ogzQnDRe7ofvJv1jfpEfL2T
2m7Cp04UP9rcHIPs8KXk4AlXsMOqopyWzYTBWhTwL8hukgmQqnqGqQ0yDYvpXt/ghz48/yuVC8BJ
uCtclqG9X603iT4oYBn7zQt2ZZ/Xd9VG/ZJDQXNkDQv1QycWv4JW8B5pcgqvH+cEoSyCSSp5VQra
UxinGfyPUR/Ii2yhgI3Hv/cXGvTgvLuUxWSJM7t0whvT1bl/7mE1JQ2ZXCQDEULKUawhit64QcHg
wPvsY/m+4PRGzbEMZBeAUIfDE6coqWx0XzHiCXgx2sUNtbsCIj+mHoMMwwFIbkBwkwE8nUfD9TvJ
GdH6NBny+TlNOtUWcQ7lXggJsVPOJ1flcxdhg16fgYCgiWMrTxcCpEVa74gdD20+wklFbKBrgAGX
JcZDrY3GaBeN9GoDvBgIbIp9AbQgh2U9r8kuSUGoiTCodMiwZrgfV4v+kwldoz8r8OCxZ+7vZGgN
QOS2JochYkO3oLyNOCjpSaZHerRv9J9/yTFwD4qvOHAnwOWPpbDXMq2gWsDDy+ZnFvY5KHIuEPfJ
W2uOOcHkDJ+7glZB0zc03wJgJX7fPMJSBVlyPno3oZK1KvLKzsr+80QElcVGHZxRi4FkKF/LZhKy
6L44ugu8507r0tGEHpCWWN7hAD+InV5rILuFEZEat5gRUp3w+jUZ2Dap7zOaFsryfGKFnQTGevr7
xcQpAxVwDH22l5fsuYgyCCamfXeZ07Ay+Kj7pDtS/s60ShAo7hh2AN4au5XBEmp4WMi8mHMQp4yl
cWj1wqWf6Z0miXoI/GeYVikwjtcYuwpLM/IRBaFniwfRjliwS+VWgmki7ud//kah2k6LT+twROD8
2FyfSB+U8rPOaPtX62DdvS+5NLfo7GLrdgxiFfBQlAlryaLjWECDdzP7VmUr/MZkaIy4woERB/x3
HlwdIpwh0QEP7m4ugd0rsUvjrWfA4JW60+HQlV6Nztnntas7/c6sB4xbhbhe+4SSCD1DHnlLPcdr
7dfvc6fVvQfPJTHiWgSKgcvUsi8TLqbPRVu7Agm+yUSgh5Lj8YCLTp8HWoQRS8F4MaEiVyyR0fm4
pI+ADuIFXFcgX6MMGGwtqUmDlzEnnyNu3xAT/3+ZmYzXfC6hrR/Kcu1eNYg0+83mJwO2nk/ahv7A
eRNMaj36ntmW6iN/9pGN3oGtImdOZubJ3pJsSXIa65jSm5v1yCD5Fq7ScKnwM80Oi4QtXFYFpqNJ
fVFBNgAiW3jLW63D+ily8ZSBvVvNXRGQUDcjtZFssSNVVsugXuoGwwKlqRl7nrGE01JBfRL2q7NP
oDGimYQ6IJGs8KGbAxcdMj/BCxbae0f51q/qI6Jz4O63Lu3geP8Ugt/cnT3HffArey/xTiosbTap
gqZGB8+hNkWR66i5tE5T356ho0FxJT0NgDQEbRO+LPkQWlmd1zlH+UWYr6HC4d8YHFm4Gj0ITx18
9e1IZJsMjECVxY2MqorTLklw+JTSOl4K4B8j/sN0xc5Pmq8a6+Wz/p4n/vImgfEuaMEZpwtiug9a
6j/mPtmZwF/Jo9VJHOFX4TFqHYgUz6CdOIwBgq/by1/qT+JxnE+R+9UV1OcYU1dGcE2cINgQ4+4R
EUHaOiD9fqIfgkqM6c5bWdAltCz4IytkBc/D+neN6Yv9MxX8p7IWJeUtoTrIN+6g0oaWkkRNF1zK
N0rulmukzah47A8T7JFEhywZGgsW2wF0h/P3pYsPoavZidSiVy1AUmjDgd0zhP0keHwXjJOm0L3M
+Z0mYjFJCtx9Cs4vHhPmS/kFl/o1MpMbEqQMpLjOf/mX296Is1hyeEGTK2Qwu2zqoRw63qQ+rKiQ
faz/AQgj+1r0q88jc4N1X25/NRbORK/UdaJD1h9Uj/vXWQdePUiVLP532W9Fh/XgDYuWWOvD58m8
bWUIfh21zHsEGkYagk0Bkc4n7LP5BU94lNpKO52mu1SIisAp32RFmVgf5kDEP1IxmE8RmwFUH3AP
O+Qwws+lllQix5kyZhTOsgEBrWnzwhhmWTSozh2DWNZYMMkIGC1l3s4MCIq3ssscDznB4vjHWIyx
Xw07Qt8yrv9dgJfGrJk2HFTe8lx8DdXfB1IjkogfhEOYQ0iDfj18JoEUdsqY/MNRl8YlNtLiGe6r
ISFrio/bWxVG0tBx4b08faevtizO9WlKxVrKl1aU8S4kH6baKldeMph7rBb8LuJFCTplZSk36bEv
Trrqfz0oTq8vI4MihRuAvP4eshhi3kDBL7QJap9EdMHZo+bmqXvKaxOpwXJn7eP6XLYYwD2409UV
nadZ/Xpe4Nig8f9ERKJBlEjXIGnq7p40h+jNz9MHEg0TMvS33V+aaemRu9QWli6tGWfKfoC8s8Ac
hlkFCsjBGICWabUE094g6fa6mJ9KiTaeTidf2P9Skh43LBeLjO9ZLnhqZhZgQWPpZhhLmbFJV4Ma
4ktr5hdFWDSfqJWFcvIQq2Dua032+GkIt7QUnDV+YoNJonYRv+bv3yQR4QXiWcpy2wXAZPUVhUpF
2ThWIvT7eaAsmsdwjPQahCb4LZG69p7KiMwrnB2w7e0QzH+Uu2LV+ANQ+XazbOFyS87y089ZUoYh
iwvfqeD0pEYTGF80tvJVStMX9n67eHy9ZllI0nOpP+RpXQH3xSvzFUr7P0ftoH//On+r3RJG4dE5
V5J2nQCr3CkD9eb10+WH9y/oAhkoLkWpZ+XdsjMppPmXTL7ZhY25Tlh/OGg5lqFcuZ7KY0vovRzE
CGGi9ahCqt3OWjRx+r+Yge4HxZZAl0wYxZ6CWN3h3G+m0UlCq6v2Wil08A+67xXLOvdPz4JtDedW
B1efxEl+Gl5waOl0X4Xl0i4/2y10y3AuizcHiexR+a63jKjYfhWu27jKv3X1ui9QBM3mghNtb+aO
dpMg5LglN8LN8b/SFENWTP8q+AW5+SOqF0tcSYlhWQ9MBZMLkky2OTj2JI3TgG4OOBZzJa1BhVnk
OvdA0dHpYurhlEVCT/ufMqjHIJjNda1y1pU0l754g8TZ5gOdli77+AmgbBljNFXzF2r7nyyR1rFX
gRXhedIex4bnL5TqUYJXVoKaOypiaFCDjGtTCQTspAeCzYlHVQAk+07G7B7gRgJZ7IGZnkgQwMG1
BAX61BppaAxR1pfkmsxBM4J465chFO3fhOWhKRAu7t/TyIj9C0YQRSnFfY46Yo87t6WlLXs0bON7
IbHvtOH0ywLJ9S6xc9hvQx81P9rro1ulvz4dj+TGQroOUclWM2Tpe5Naa8Ruchzppl++jmpMWzRq
WbyL1bo5eFChq6rfSaBN9hfxBkKJuBsxY+e7cjqgXeEtRBroE9Ty3kzFhCtMR5QHmKxvUYbln6XU
CJ0EVyGnQ+AHTktvMoCI+tys6ICQgMOEukBy/MrdcsUO2BFGtqf3U1H+Bdu35yIWbe41oZw4Cobv
oBAhXClupBlot+UJwEXs5T8mZQ1ZDLfp67ZSL0caRWG07IoXKih0JWflKA1PfK6T6F0zzgQrCFPK
vPo5tUpMtyybSkOQToMKW3TVi4GSbUpsI/loX5UYKsdZc7w2JBWBCXLvYIEU3tqXZ/53uRxiUVTw
iook0HA3p1h3+eOoxnGRLGsybJm7mE7DurM/H2tyla3laCRiuRpp8VQvEAsYEQ9cWgDGAHBZRF6o
JBfbZfOkyxUqvsw+L3chQDHTqkeditGr13MXnCoSjRLfXZ/0xsjnLsZDRssU1Bi5GsCzQfautfUg
Qf4QeZwzhwrHflFlU4Yrr4LHEnxwjOmsjF+QdAolO7t4r6EycvKODTr5TXV7a1oO4Q//P0mv5dOT
Q/aiJbP6kS1s8peOigf8CmzM+38IEa6CzS41SM8xDjHwX0zKwS92STgBe5fctEKXCcZWU6PKRP0B
eP5PsvXO1jqpadiWGDULsIEfYHJ5fKGwkl2MROOwjIe7xQNFzB32ii7F9Dzh4YId4kERoAUkUqpW
s5Ai0IU+beCcjvOS6UUt1GiQVudDCYhD1mRzo9GTG3n/GLJPcgyHhrDuP4DvTMr+M2iiDc97pDtL
sdJJtIIs/+tPgyC+7ztMOngnTxa2NRxATzadvgBF3P6zFJVqj+vrpfhIc1ElEMSa5WKxyPMJRNwL
p0T9OXCBTf7abrbHbVkVcT5EUTbj1qYko/AZIxtWpYuFLyRMODCHKfMq+leN/od6On11w+mAOfwd
J/NvU0Mr6PhFxL0A0b4SG76LiYILXTVEmsW7uiLaXf1ah8TNA6yx7uNBK28V2Rv2alq8dzVhxyAk
mIN5/xWevRROMb/Rl86VDIMtW6zE2+czYNIieHXC1vwLNwx0H8A/Kmo8JkbLuoP0wdJqvis1YLim
u8VMRZAr8/fbyZc0m/IAp+KJmG3i6cH5Ea7oMgcDta2jaF+Wil9Uq5htMj96teOXXyXuRPyQoack
qxJk68bO/EDA7ETpfsysXZ3TR+C2WmBD3k0PWuHtVRSns0/kXnH0rslAsejAezpLEm3q7LobULiY
TW8LtK5RQ+TjS0vSIKG7eiKRI8Fqnx/M5oLsWZy+pM0aurhJG5huJJPrjqPDmIdnS2ir7v4Fqu4l
at4MRQhMTBfmJiOsmOFBIZeoBd6PIUJ++TlCLKPHNbuFnKNghy2HVQIwEujaVtLrtIIbLb1tPUEI
gdwiAIuDTCORr2GxYwxC/ky7EN28J6gqM2JVqLZhKbE1Ik4i6WOctzd34IDoOY6DwRu6xfm+GupN
bUpNWb+DTDERyyqLlPsQ8OTdF5kHHbllyjrZnE5N41qR8UQnF4iWRx1si+ZXjGyAiEZ15zW1U1/d
YsphsuKJGK4iqOZAlcRy33zRQRu0e1CHQWWeoMS4z7NOCFSGMeH0H6sCXNEvJQbgRYpRUFY18ecX
S3T1gSY3PzE/YKyjdYSKG3fWQN/DpZS9VdnC9HRutzM4TBs6R2jzTxb5g8Bi4kW7vsyek43xNekk
YlbZ3e0Wq/vgVf0C3/5lMc7sxJ4J21pkqrnMjpUyYSAZyRi1c+U80SJqpM6txmqf6jP+XjxJJ31r
m1jlQdNnQEHztFRUpdzX1hb3imTvVb6WQPdphu2pzsc01r4pnz71CfacMyYE2TOxnhKBEfdx+cv8
HNxqBTKbYWQG05lEO4CNNFSlSfK4b8qo2zpe/12wI1ZrKpbZOzzBSWfJyANziF1zVBi4k23wmTpH
0pduHf7ZEdA4qNiNI7UEEIvfHjoghaOQVEX5U0bS1aTypyzZefsBMmrlcYALNebmr22RyKzOPbpN
hrR6fnjUqDDIcf1cR3Z7Wh18ZXdF8214QU3XLUi0Bf36f38sp5Mn6vqZ6xTJhWhDyJ/w3rWDk4Zk
dAY2YVvjZFIwj49MRbQ/NEMRtRFt0LUBJCn85DjMJ6Cfq90td8TsESPeGgvoAk7fAcKfeP7whi94
Ot20w6FGmVTn+BvZF+svydImT/08vtuZTV+NEumjXmGAaRJO1GugQSrVOq4OiHkxZa3Xp5FMouET
YhcG8kMGwKkpDeCDuBamxdwviXdB1ZbrmxaTbXDPhXFZgeNwN6iCcXHzVXun+qp3zf08SPq5jaav
sBnSrXL4QTefngqRGiyA8jzd6G9d3ErvjHXkapgPIKa4cxAiC2PaRSeKDQ6R9Zhj3onniDb09GQV
t3Cly/vJBabi6PEB2cMPw9XuXI7fFEnRH8I8vUtCAsfWKQSl1svHJY4tIuRAMklzj1Fg9pZvbeoz
aYNOCUt4Ub1GvNA4T6OjmSIRbg2o0TygJ691OJqUY4p7TDprrlLAhdTEPZzUDYeaCpuli1c5A6Nh
ePk7/QHVvNXRj47zqFQk7scU9yiaDoMcX3iLeG6TzPJJNyt6GmLpGfPBI9e7fgSItLBjPkF/VYKP
LlMiwvk5XGBfnXBLPBgnY+emVHwKYoDSrX73vMqWMh08LwBiligzApESHJMoNaNDKL4vYU+2lYz1
wRVV8vcsXe2dMco8WwBcIyS8AL9flnBkIqeHL63DTjEKK7i3+erWC8n4Ry1sMGVgrYgIL4VG2rU9
H+A/rqYKDALaYa2silnYB5CHf6xgir3mIJ/+I6hoexpw93cDPGqADrVXaCaQZ3gadcxtcoUc7lmE
g+AAPQ46OQsp5T0k5aTr4ukPWRsv5q8DGmjbAl1aMfqEpIUhEWqnA96W9D0bd4180EXBZ8OECF0h
d1DNVdTp04X1sBFJ5GW+4OhJu4K5025SK1MLMrbUZpvUEQPnvE/A8PhUc1bkT9NOgcqcN+l6ZvqM
RhmHTEdMMHjdPy0vUW6sqWklfqR0rs/ZEf0g3H1BJTy6AlgWF/f6IXgPwYD1pCHFttddrLVfBMDi
R/H3Ak/8dqCYwqDpJWWmBWO3zh04HLgSqZkj6fdgLGWYFSwY8i2wH6X2SyhcAGrrGf3AddG8WEJ+
pFYSzmCpBGsHuYw32hfOK3Eg00aR8Z9ECuJHfEo4o+3Xfx+pVT/T8+6zTNX0u0xNe1GKop1gvRxm
wQX6OhlfckyKMmhuCYV34+Y1OS9F9bwSH5UVZQrgNPfBtAQKHgG8+ykc11hFq5JODAw0eUFOlJQn
aazwON7qjM0HpwMhVFGiKg7XVkxJ/r+tDnWsshwcFtuDaw/GzpL/HnmayfxMHly1NMJ9kF4Rw/nU
sqYjQBYIReH73DHkiZGC6akJm/cZUlpkjdoJnWazf5az5DPfcGtGGIYIG5AuAzVLHlDaS/mMcFTs
OdVjFTGlTjq/KKkvOSCVxr2YjxMfk3c7mzqLZV8pposnOgc3mpyuIevFjAlyegDI+TYBDkoveWH6
8CFJ3KGCIWqqBzbOQGfuVm8hUTgO7+he2fbyhXR3jN6fQ7A9zvEYaTQeLKzIbS6uTEwqbVVl1x9L
GIoGvvdsvO5ujzTIpmed9JDO1UNGbCxYN5hzeOWBKJZRWHX/bKGiNcv/0ZNHcjqoZSnjcadofH8L
8YQWQ2et9sPka4VNBJcp7XFYk60nTRzkW8/ZrewyEpATpQ1+ft9UEERIM2Nppd6XSFPJzv+52GyW
qtR1g9HrRK41gApwIbdS0I0wc/JqHgYbxFLqhiiwB/OW0HiCk2yfygwJtph836EoGWJdFuCQNuyw
MeDB0KE7BQpo13LvNVWfGHbu6au+AaI5VPfqTvTXJwFeqjgeTuE1H9iNFPhMsdikGkGKf1++umO6
AQD8FzjI8mvoIuVoZpUAWKvt9dQup0O9UO5DhAaGNQSkzewIrrhc1hwpi7/wnxfNvWlDP9lqOVWV
8GqEKZzgDbCT5VzzY/FYKhOtQZeva/UmpnkPAb2101fZTyAfaFrrmFLDGHQy2QFaUTSZXJBuXYsH
uFRj1A0t+ALLMk+QiCQn1p5NOQVuSHRdA0ng6BcTxMK4Bl61L1IxFG4KWl8vlgYb44fMF5WcRZ62
UIEzD9QuI/2VwDEH5O0jBOnDCuTa8l1qQ40os4u0JbhFaXNmlcKFcCIZAEBGGBAh/GQT7RdyyJwT
PRqv/SvFT1+lhJd/l7yYSjL9ZvbPauoT4mCFcWABT+f3pxidazS1ecvzH0kPpLNT5PDEjq0nuU1c
LG/VN/5ePzL0PS9wXkdSW+DBt7wR4M4vQAU6YIa9tMopJCN/zvuMMkXVDNdgMFKH8UbNgZXbnByi
VThdkbapjxe6shAzVNHVL+LdA9mSelqo+bs7EDNHGjmkct23EB44ocQrsk848HQcozpvV9n9MYPg
MhIjm2HTtLeVxYW35NKXWNv5cY246KL0NPJDYCS92Jr3z89ktTMUZbPYaYP01AMWXKF4T6sLDjyj
w7V0yiiKPwXGk8lhyFboeyJBZqSUD8aq74cDikxMx6oB3mce+ceY64SN284Q0g9cmFjnPqQpkNqj
btqKBxMJgm3RKpM7L3jo1JBxoNXBSOY06BOTVSk7/oUauvPHuxVDIBgxe9WagC8MCffxY6OcSm+m
fjKZxYevfr2inwoCZ4/UEv3RhK8Yt3aYbXugBD+WbtChuI0zsX7xc6dmJMe8Ii8rRPYWYCn4FnTq
EDfg1Y0fPb/O/WyPoUtRbmz5VbdGE+YqZFpXmiPkLS7shBODRmNC/xUWGxo6Q2UndNE/gak4YeRL
UNKKKpA2wdJsJC+Ifud7RGsk+VFu1awz4zavvCMXAmwTrs1DdWx4NzgUYV/Ptisy6ug7nhsQx4y3
YMuQwCM9/Qfl1vy3rs/gmRF/8MELA5f8XYdwQkGZZOqmVRYfdIyWJUg6uvgqYMIjoRJLipBJLrnk
xseHBwt2th1SVEKbLwUMif+AKa8Ylj2yv4bznENoBcpU0HwpkoSz9lZfW2cA4KH8kVUCyTL4y1TA
8rhkltVKGy/j4k1OluJc/V7hXsimCqubYaU7YU6ruERxrwDyz9OTIBdiy/OTlrRrihEfVhh9Kmjv
JaQl5F5neyLR0GmtekVVj6Jkp0Ew5tnQjAsRD4e/sS3REccvFgWfn8UUzO+pHycrkn31S6Ki1h38
1zVyxRVrTg523z37q+v8SmZXS4xd4kAMY4afsp7wW6U9H4I5u6Cyl7FodxSpXcq/mQx414QE45ex
QI1aGwxidfX8k1SR4wgwxPAZNgPbasF9kNi5q9zIF+Pt947S79TLkeEBoxYJDWpvLz9k/m/1zpN5
01kGAIEy/t7mekTyaHWIvQoT/dMx/qpA8We7bkc98UB/sCdmIkEcuC3DkPdlk+wZTWOZ7DuA5xfp
2NKJZgL1VOI7z3LTNvdml9YGtK3rWTJR0jySknnfoanHyL5yJtHAhl0J620KJNgRA/t5WnS+6nQS
1jAgoHgx15nZloblThck4D6oGnGBL04YdvenyJVi4L3oa07Vy1dCb0gcgQH2UqApw2EWqnAxudWE
zxUs8OphKz9KfadBLZhBI7ZFr1Nc3vW1AhHwfENmykiZ+FUGTa/7PKh8g2DHjDb4w62Xrxy1ZnRy
R6f99PiFF/OoMO+WuIQzYkRu7KSoc7iW8lbLqCe8Yz460xY463qCuHWja/IUy57bItoVAsLJbsp1
bo1pS85Xu6g0XBU6nFAtqn3s3l+nMSoTOD7NOVymLT2i3O/8vv3yLD9vrZ/Vrxthav64wG5mdNyj
BKo79vB8AQFtI+7hFTN0MTdb5opwNGPQrYwWY9zGz4ngPjHWE93gid4wVWBtZYP8zfLWnNErpmKK
LL1f3GGa9bQQUAbmv++ECKHGWLxb5LOF+KdFQqGXoEETwhlGq9Gg0tJYZbJQSHVBhve1lUKH2Vr2
FvQ2N1bI0TS0dL7p528mYoTUM0rYWTR7auE5YlrAZ/Y/TxeUK5dgG4pGNkOibj2p6EpEVgIPsvnT
k/dDGSKnnr4gkA7tMKLQXTIY5h9rUlIDV28qfPt40UDn+tHWiQrSXcns5sK6KsquQ9VAyYjSI6ho
i0iZyrVAlGL4HV/3F3m1hXzXqL6Ddz/8McJmvpthONO11x2T9E5bueAdZ+qospUZtzmSNOKSDHjx
S1T35HyjTexByXY0huKjxnEeFFRER/oQapLBDnKsuQa9H70LUl9mVZe6K8So+0f5yEdw1I/DTZXY
XVQ8XDbz4L+9iw+Ge23DrbM1ifKz+vgpKwr5FHRNNWDoJwS44gaPwY5p7ujPDGbQImEulE0S1aOd
YOkJujEvq/2Vw6/Z1o89cJAiRWjIqGy1isa+a4fUMvIxWGDrqgk06Ew6e0FBR1Oqt5K/cuY0jPWm
i/PETljRD/NOulkdDjRBYE4Xan4xga6EYZw2deZAL3PVptg5k/ANBJD9C04ZaPLP0pVCsgXgyUOA
zochotbrIoGMDkl1YsYa0uHLcIU+wq2HNfP1H1iNpnTfgRbxq8YoCoI/m0xsQilFdm0lmOkgv7Jc
iGTy4NrhiODLARp6Zv91oQhLm1MuloJh+7z5Mv6tV5LJkZIcBZCeaQ7TlOuyg47vZcVJYVGrVx27
8+EoIULQqFyAZQLl3AzJn4cfDtMUQF/2ZGbdqNKA7vXjtb1kXMZ9thcfRD51G0+KDZ2Z4Bsckw2U
T8huSiNbGCbGuczAaVriovGaUFzbOnGB2WLLAgMQyYtqbbaHifnRUiien4SOOeBOgmHCxStCse+N
1cgRPUwRB4kvwfrYUanxE2kJDKavhf1tQvYHF2u3dgYhyF02bRVV6Uw8r35QRuA5EzbrBVU5VULN
GOYOKV34hRBVi9WTA9gVpPLkjwQGQcdutPREOee6rWeylhD7RbkNl36JQaYQQ6KRkMg2pAjfKQpd
aLDybrJk8kPQ7ZDkqrPGcgfStsadXWFrLx8jAhAxT7kEwxtT8v3fRNbidnKRJdRRjY07UbYhe7CD
P3mDWwBG7hx79WOPVQKibxcxsqbmpXZIG76zUXfvU72gSWoJWd2lUQaOeHjB2AmMykDqm7+4vMmc
gizTS8N8/sQWKj+RjSWIOeCQotKaEcq2OkaYEB5surcHWivCSDZgciLmn+T4ysLZtXOpmv7q+bX+
7ORDFL69l7RCxMPPlDjH0COV2rXTHhdkfmNFWz2xvaTkFQSTCPIUXrcJ7kpAeHntmiGScxznz8Kt
f+ODKXq8UhqRDiQOQrkREB4wulKMRlDHdO0dM6c8rgWE465yxtMDkVUICabD9OHwCP1Cy8mFjh3h
1o6Qj9CbhZTSTfWZGmBnkR5Zk6GPKZZswELWRd4Ay5KWP4f7RJZFXBOKRoAJHiDn617F/IOxVhs7
QPNIhg/KYTTQoMRhgUT9QtNAgOqQpMWHeu5UALdB0ixFLVwUD3Eblvn0ltUFgagEo85n+RqvtN5l
6cDEV5KtgiNF8NlA5EVhU/LDfRECSB/yPpEc2k/e+L+7uS6tSE59dg5pPY2u02zzeX8JmWxJ5Cf/
50iJ9phcjxSDU2ZyvA2+atLavB4R7g0M+rEcz8zVRl+8x2KfVJKWriNUtiiXsttFgDBwZr2BKErt
Hm38oUV9+IhgccEKXx2Fsz6THzLRuMtaD4PnFgAdmAlT+aBCcC5W1sGHopy6SjgWNUEHFeq2LL3V
x2rNrOh/iczZkBZXvKbWKe9pqbP2o7PwFdoO15/egemFAQ8KtvpFXcuHSxSOOd1S6caxNDkhC4ba
onL7pIZj+meTNRBqTXH4KVFYi8L37y+5cg+/NRHaQ3XLpM9XR9scvFmnm8XYiegSPmkhVs6I2hlJ
t8i29pO9R+X120dReoCIjfbYNXodNKXcgHapMzmzNsdFjygNwBouwHVUrKImamDMTkWsZivJhxMi
r1J1AsHSKsWYKyE62oCy+o9hqkviWvQJs1rURGJLh5RTnEh+VaKnwITRCWrTJQr6shqFcDqWMfo6
A3iw7GFVRyTgUNV9tj1t4v4jzS2yP6SdqXjmPEeOEaYm2nUtaiF+oFxykY9XMCt39JKrQOar2kt3
UIK2glUR/0s4eEcExCfnCgd0QJ4hYpSs23fXnJDS5d5ddHi8FlyOrMrqmCUt5KlZ9c+kNzxXc/o/
AAsOFk9fAcIupnHKtgvWoweNRmocITyMz9ZIPzWipkKA/NhZ4zJPPp/pxO+ApCxuKQvNnXEkJofi
ujNHojB/moKI5CLLBXlfBZT/N0uRQGXqpuVrmjfdNd4INV+58uVbhFy1FWeNfe1lH0tvteu+EoTX
0ryb37MLltoB6EBp939hLZ/xgDbV60+C45ojS+pJFLUrZ218ivtgE7Qje4mV1TZio+cyN1lxjZa+
L5cM2ENOCA2x02rcJwvFAbe1tcbf7bJPV2Ufkl1N68B+q6C3k28FzXjAyZS2KopmhU192frX+WBx
SRxzlrh3jg3gRx1n5UHmfZnL8vI2R3uzOGE8X6me+9EcQfoOxK92uQ48xr0B8Bh0FungiyDnCqEU
UmdsL4mKZcLpwE7h27Emop0tvB/HqQ2Zbe3f3Xu+seAqBL3EJuLL8olS1tBRl7SqOsbmgnSqmVJd
A4Ue+h5jPzd6C/Y4mWk+Paav44HEFsIm0rkwkCJRZgxamLhcJt0SQEOHr2YTKV6Sq3BkeFeutgPN
T4HDg0mJR1jnfZBGv6Doq9J2kIWCvNEQtfYdBK22nOD7bASd/wMYZ11VFXfzWQtcSHzim8ObzMT0
SADeG/rDAKIkPLJeg3wcfw7UqrWfnLyNCSUylB5rTLpP+bzKXzYy+jg+6Z0gahXuVifdjuReNkjL
Hleey2g/XV72F4C/rZVuKiD1oIor3hDk96W0lpNdHhHNCcFPCrDVivhF8jQII8sbFAnRQRI949Wj
G/L7X+T7QWoYHbcMq54yAMTzj772noVg86i7URUmid2wX/b+zMLXzAMsOJNJZ7X4k/FiZAWnIudX
hFS7mPhPrA54cxJcSKze6bwWb54UL6x4Juq3JXIKOGi7dkISEAQ2F3fOhcFWULZd6cj1WabbxgIh
v+jU98BRV7dRweGpce3nLw9cz4V272zA32wVozYaE9gpvMY4EOgHrYl+OlIodbxt0Ti9o48TOgD1
KtPjgc/b1vIpjO4koo1zx5nK903rGh+2UoFP3Vk2tU/pFG3ZI13HnwVSozqvFOrttJOzvOS4a4nU
MWVshA0EvPvRxmsphBbKjZSEN09xBHmW4dAoFDKG02ugFJ/xBCrfvnqMzikpLiaQuP0/TV5kdb3s
9wMiYGuTztc7GFeHvByZv3PpeUwtLKlV2lSxqtc4w7A3sqQEjr+dnGR/Wy9n9zKWZqbiHb2q8Xvc
JpSlMbX1N1DWxU3w/wA0CEDyPf3iR04TD0V0OxRJCVJbVphCgZWuYuzZy5G5jNmjsqXUx0ToPuB7
5EkR4qk19V3X0vbXUFwjCrr4ObYB+tpVNb++OwtkXbh+JqKW9s+8CWoWeb4Mdxz+W+3AseFgcP0/
AzoTeHubvp8ckjfJ948+0QPiZ2laD5v67TGFrZ8iKQ09XaX/i6Lgq54BYVJ39hN6kwh2Zfu4uMEA
wuNUbAn26LPB4FGKCwHsa81oN5wfHYrPQEJ9M0wXfcOPum3ldcGbivLFKS5zWhyhtQurdaW+jBNc
Im20jehiGYbf5FL+T4P7GRXGsxmEEM1VOSexQGhd+UdJG2q0whImkffwu1lh56kXY+E1aR1rvw7c
EXHhJaO6VdjzyxZn5adEYilIM5OyiTwxva+8BnlwalXrokQMUxsbJ9u4Pn/mHajtEbasc2X+/CLQ
8nX6HbrrTysi9Wa4/1cZUWhD+Ml/0+jKQ+V1HywV+8SMFfLA7DjQ/EgtdYiwM7wrw+62ZVmiD3Hh
mV2QP+PI8wcIgDOaHhGpoW2Dqn9zlx8W/7QWzA7DrU1P5Q/v8SlIxG1qwKz88i6ZK6/T7A5NjAE0
TUP7ShvhAc3gFxbMUYfjNfQLQHGZQrBiSpJILXhe6z4IMwHGd78ChzubCvEdcc4ZYLjBMIdu2ubr
Mv45aRvA0lKMldiy3MvvCGaxZXlVivBEK1FMdlX0BPfKy2LOz0IhQy9WLXFvh0hiRRvJCDdiX6St
rP2ml3PnSNMK2LHvRWv4YxFmj1LICGdJNX7Klw1wq0SVtmuzvWlAy9U7wYk3Zj2/BiE6k43pZF3z
0ToniB1IU3h/H4OA2BnpdZUR1BJfKAken4w2ljsQ8OOloK4sja5JzYWVRYpSSdbEoFouZ6UD9CSx
Bx4OBEFaeYn3BdlZR/929ofGeGQeTkztdes4cIX/KgdvxwozhOlOWiRJIM0wE/dszzTlT/AvMjFN
4yG7LTEECgzCRs1d76/9re5KprxmeMsm2dFAqhLtbDPfgQrm6qBaKHdmT3iOuTxw5qfF3wvA4SIH
8Kw7JOCBMy+GLoIHPkN17eOox5hF7b3V/uf36Gs1ZGIPpRkWs8epbpwdq6Mi6oKUoooxUC9kIDjo
K2WH8Yz07lDAKKz5OVxPhMoPq/txx6kqtKvaKBGhIDcBkGivXnRlRRXCykOMDtol2tNWb3p1AvcS
JrEDQYc+ev8EqbduRWrHBgrtrVXRGRZ1F22cmUHGfj7jA5EhOts2DEWEqf9Vw5eYqcyZ0ajEH0mr
474gnOw9C+XoujKkhfjUuH6wePY1PBgAbfIf4IURFtykSN7cHym/3vsalf46fI/IekHkh27A0pf+
WO3Yd/yK4IFYhmIRjBoG80zwwlzcDHtf6cQw3j23W6XyM5TWqbKNuluecLjP0frN6Fea/a/+4cDj
u3Rl7qcOZGhrL/LNrFlShaIzDM5LRCraExjmiSzdBY4jfA55hEnY8yQkesNXQ5P24Lpqql6GS8Dq
HEJ9TAkIYigHIAR9Bf4YdEBYrxjSUsLGQL6MfHrkjiuni9lh3PaPR+Z+8pqhYzwiq5eTEdHGaome
0H8W4Q+caXnkTyA85h3hbk90wvONSccd+4WThau/Fyvu3Gzz/zP8nk9pW2WKmlBBWWYRTiosWsMt
KiPLoPYdLoHn+fy5wZEeakUVe5FoMvJmEwMANj8C03YFgVvdsfub4L19vBzL33CySdFUyyuu1bK8
BXUCSAMnTtqjBavm+jSqxaTsz9/AZSUy8n2owMRVJ794H3qxVqzXOWYm0cLz+J10/uhEdyqdoJkb
pa9T/pfJQP1XN1tCZWBjA9zCYF+2bEuT5+yCxLkJHdmDurZGbKJN/1OQNUPqcneut5b8yUikj09+
XQHknSuyvyCI0aXuquCvljg+DDjPBrXQ3BSdb9k/fsUg9KL6tlEfpS4erjY7RxkFfWyM30EGB9Fx
cA/fiWithQnlj/2pw7cXPWkW2w1BpdCHpTF0vgbKSvcu86OJVlywTxyX39vpMJbfawMD+7554XhY
RafXZqIWt2SVa27jUxEsSi/07hhittt91jxAkRo20Gf2TMtyJrHo5zq7/oM7uJCdoMs75cku5+8L
G6kQd655X8+4jEFd3WlpLrBznkO7nYqF6Ahwx5qsF0NUx3S3X8cqnIZbFj92XE6bZifCKHhwgYOb
KuhsktklcPG9matYyU4SnZm70gVlxDf5YFBrRgpSFSadLYWmElgwfEcUfcXY0tn4KgTHiAEzCUHu
+V20ifMi7LBcb6OVnOD4QHpmJi4r07VeEQNt7niq6GuQmTxEJYxbgvHCkTS0h6wPLu5P5VB6T1Wr
mcwExywlJDfW64+rIomP97zrWtj234v++pRFZD7J+GBFCifqcLUdXVwlxKu0fxgEtAVjbtoioFSt
BPDehXYeHg0QJ097qRc0iH79AsNbq+gqp1kcTfJ9yDGbKWHmwCqqKn27VpSQS2eHNwoUZrOlsj9v
tHGBtnb3xI+QuXKPLRJBCS6Uqgc/+ik81I2vsXrLIdao+3e6phQmc8fNzeIhV1XefX3Kch7ts28i
r7TSuTNsUGOoGkk/xWf25JVWOslmxhMzdWOQPQ65+VsF6xZvFTQJ5Nzj4bG/pI2UnK2KkzOoXvth
INb/yKaJl3pYqAl9T2Fn34blNw5PwEVytGG1FzHWIdDF7LnBonfBBtetjXvORVMj2L0SvfI4wovw
r2pEHmK3zulthYnkV9YUpP0aj9flKKm9DuYjZxZZuFFB1sceZtvx8neXnSHaUJp4UXi7amdZIxiK
B1O0wzR5lwvbfr3JyuTkispwujRmzKgugTK5R7fAwa3c5YQWFtUc8ZbmubKyjrkOBsAE8pn3DArb
wQzgRYAwiyHP/PJ1PwPmxGHtu0DG3TgsCIqY4Xg0SXRfrUZsiWnibY7EeOL4Am1u3K+EOeXYKVFZ
+zoWEvyV7KDoTNVDFEEsOD17tgzIOMjZ+L/4LaLqqQXPPkSUrqc0JqpXDTfhXnMu26C30fOq5m0r
Qa5u+YZYgTxEBGTlmwfvQ1v5CjQO+LuWpjHGKisGCx25Nh8fYo3tscMglHuHHUmMJyidA/yIdMEJ
9b3Gxngc4idr8aNBkGRPiRQgrHZiDMARoQ3mhNwRAm4qLD9PkFdKRnHTawaNTlAnfo7bcjboQCUI
EZeUAX29zBhP5F28KmFjWTdiHFy9386gTByH6lTFngABiDnW1/cyB2qZcvidcvURKQKv359BYPfR
2lWDv2OnzK6NtEUY9g8p+0lSXflfZHp2nSVGIzwJZDS7NoC6QaBRK6YQbZvvR06fb+gKNRYFmfBr
JdYgBMPmDf73OB89VwHacSthQAb9vH+NLNjY3RJSSDOUyN469uCasrEGSRMgkmvKkrg4VAEFpxkE
5JvIwmcQpB2E548hxxbZ7C6Rjm7js5r7jOOAyqKyC366INaF+exYc+DprNpbzNW9f2WCKoSLno5H
87nXiUTs867gxD/2+9X1BMZuCb6P4oTnpy/60MlxYixlTNSRBvgo0BQFKXuNIlNTMOc9e4lQgPm7
OwOJP11E4G4FRsGoeRrfuWbpnIo+JBgCFc891511cHx4V9Jx6MbSx3o1iMc2QwbTUnH4IqBicwXm
D7ZC396dd1gLgjX5t9THRveHtRzcp8+g4O8CN/17rcdIDH9/UR/aG6Sm7SmQe5j3Nv9nF7+Bqo9j
yiL0cHX1VV7E3IL82MajYUF4UHYrfxZrByyQwcGv+euC+UySICNVpl5Nzsioy/Nw4s633rosxJp4
tBIA07rGO4YCY1VnusNA8OIz+/p6ifYwqM0Ju7utoFYy1X4lRFHCezvW8LX7ctqBxntkqRyKCLqv
WHrVJ/rS0YLl3w64sMkfL79TvYoqYdMliNpe7bY25erJRQiNWKujrc4lnRdKhMiAVv4lF1ixhGTi
2uCcb+HLFk2CWX+T/9Ji6g221bdKAi1I+9q27zMXNPUoxQh1pWWegdCcKLVcFxd6y1tmURZ/xMSx
YMgo4X1PXsQsyrONqK6hS0yKaavRWROUS8A7A+VY2xsrJt+M1TkI8l/d+jCLOGu5dtq3hkbM8qbt
uctd3vZvmi79pKZyAXwy3cjsaoPaxZgj81U+b7ba3LTWDJ2jl8ertMLdYmb8bkh4rZxvDLy3hd6E
IT/2oUh7ABsC84i89tCLblJ1OgMiIOPFXbtZPqOGhlWzsr6K6i0+eI7T6A+XvgFbxI4R0Pq6m92R
ZKIWM6shBsqLQjU2uhsVvws1CMkCXK3su535sqAdIWKApAYTF6BzJNWuzh4bDGbEYSaFw2fENRUc
vU1oYRu/TB2+URb64aFVaYSZyk7eGfseqzdMog5xdiRulbavCfnAXRVLDte6F6VpqJUIEShhiE2A
isWG/U+Cw1wJKLGW/miLBLuaWn1R3ez5iPcBxf8qiTWAtgADlFGCzrxroQ09TM9V+oQlzSRwUJiK
wvklEFbUep2x3v5wRYvCK9SG6jYnu7OYl391sAhg0ZgXKn/KJFbR8JOb4S4XFWWFHyz6ch6TEHHO
LoITrDTQZMsnYbTGaiHUqja57Eiul+e9swUHJvhIp2wuQf76/A4akhF37Sw443CtM/1c2JJdL5D5
hj1gmn8Vl3y2SyVDbzY+ofJ5vz2qqDFItrEhev2exOOD+g+TVKVmiEsLFMw09Zn0ZxTnX/tt0iAi
RI1cEuXl6AC7kqaEPxZKyuKwu4b1igxSQa5h8eqdKjuR8cDzutXhsin5bZ+w2kNDustaw24dmhJo
cBQi5pljQirgRewuTpw4yMmuiMQKizgQRF7DQp5m6bd8aF7pyewIPM+8X7Qvi5TSrTq938crfmyp
k6SOxQl/tef+DOpYDRJS51UTDncGOCzLQds+EXEO2t+2949Dc/WO01sR3JMCaqpXGCxu+R5q+JDi
SWS2P3tTaKxf2FmeKu3fjFufO1aXm96+9jgwa7kUYuL5sbF/VUJr5hbwBzSO4bwVgyuyYAQGmurJ
iGNYS21L1moKej2ZBdPln2YRPrl/sMvDA2yXWIju8aNuZZGpMjqb3U/SXJemJkQp/JA2hijDwQXt
Ea88/WvsP/QmDAYPHILA8nZKz1N2TNfvOHVk0vBtVzTshcytk62HuahHwUpGw+ZLw4zEqWcwSD9e
PMz6LhymPn/+d9qcpXy040NJ3WJtOw1v1ElVJRKnmnuf8M48bcOkZyNme2IuMpyFL7UkhuwzGLhM
aN3ccGpP34mrn6ywnZq97ziE65+U1TSVgcj5h8QSTZJlYOsW5RUZs8qQpVt/Ao0iecW9U4ZlpfIa
jgT24OHMMkJV2pQF/TdhG0+i3w8k3o/Un5zgAmYXLVdLPT4H9yquRZ3CN1p23dlv2ZxBNZJPWG1M
G9RTe49ZWG0xS71k0qByCLoe3JbOCmxC9xRONK0mC72xg3D2rNXBrrk+ZGIDqzVnaiVxNpU80zKy
3gVFZoKRZJSSHTowBaNSeVKuAPKwLUroun3nDSAV6vSzzC2MOTnERC/famix1YwEXf6dkNZqgaXX
VNPwTrWFAhcjUC1+QK1pnCVDm9IFDXHeBv2sZHe+7xGTsCk8jEtbLFGbgmVIDWmIhRFWWrmqp7qn
hX65GBf7Z94BWaJWZzVxvqvnBxYILFdeRPS+e+BzCUjjrn+Ta5H8f/ZAzGE4C5/NCJ4qZw9qOYg3
xwN6OxScXibwBL6RKbVLXbZPzA7nLiHFnh4fYfq/AsAFOia40TIoXTh/p0+B+4Vous3qfgI0sqE5
kX3aedNFM0x2sj2EY4VjjLavRufndIxcahAu44gthfSFJPgNHtxNFQlbva7IilP9gBY9jT+bPN6H
lPNwi3TPmInQ0xLSit4Jt9rjg9st6G1uJRHI/0oeY74boTwdokvIRVb5O5ClXjWz1e6D8x/97bRW
+V03ul1eU7Ht/cZdeMcVPDZzQ7zrBWP/TKtCCd9fF1w/0w+WYuhkb6vugKgzRJXUdOpcpuKywfiO
Npy71iOeFxrU4YzX+cktPZXLzUlRRiT7EFrqcmcXHys6tVr/Sb+1f5Z/gnGIBfF+kftO3VE/glCd
DQeHsgwkh72pLtKfK6dH1y5S4CXxtM9mdV9c9tZ+6mJ9S41Ryf3RpJP7yBmm7Uwm0QES689byRsm
lCghnJG7q/1Fno877x+MkptDstABbXE61qEDmfhkkTiyG2URnififhDUwNK43AakwvuQWxH8whbE
VFLCUdHyqo23YuMt4I9J696gjzNHFLEHaG+iXxkpKDq6sDOUAn1/KhP+z16VgMinJG1U62C01ABu
Rr/U2uTcXJjHazLPrcNPSZ6mX9LI14e5lB/XrKe/39ZKRHlBuJarckgXiinBzixyHNYjBmMfc8Fa
bJwwNpLzBbLqUB4EqA0mMIm1T1Lda8VfwEhJ3yCF0D863Y9WqRejDxEh8boisdrQDgWB3GMR0O5q
A2+d0TZUuT2332g5ARot5crcjZ3NvvcaO4p+on0UKDNu8sLD0XSy+Kb+aqXz4uJRXUAF7BKtKRa1
FN999QcBRSN/8FmxOHvbbTfQ1jalN5+08CIJKwO3jsaEZG2lX7V0aE/yjF7fnwfxIU9VQUbwWOVF
3uNxCypmJ0eoi5B5ZWOq3mi6w6Saje75uHeNhpvjaPfmzmEE+8Yr0ySHmogg3hoYh2Fth2sDzwBy
axTGrg4Lt93OgRu218AYOr83jO808FyuTueq5HIB2scVEWzumAkUFvH+eslPkCbxoQr2GyI0XCsa
2ulqU7anDT45m9pZnaE1duq8q3BAeNHtXkP3bUwEiPP4UDQZiCcAsHLYtJVX1YMGl3ZwumOqG54u
+RUT/sKtN+6iVlnwDSdGxe/yqbgC0nXQAtF2/ApM3gV0IBf4POCWVHQkwcRZY4LKfV1cdhF8EmF1
aMOfk2bAORMPdvrhr83LNuNJDDiVZTVC5bmsq6owKMRK50TrwuzEs8Ep7XuGqOXwz843NQex4rCi
6Ev553Idxfic2y88ggl42deBJh9rU9zvvF+xDUNyf4ToNSh+JraZX6XKcxu/cR1WgTt6yBvREGNO
I2tiGbz1Mr7JganoPjtL4wp3YcuaOvKVW3OMeuUlEcUQ3Bt26OJkiQUuuutYJyZlduv9q+WHCczj
k9clCxRgnoLb1eASGRmoONRLEMwMipa/9Ut2LPR2WixVLTplHbwqMr//HvP7eRxoEK5gBlt09jP6
RSkfBeaWZGzw48Nlxy1Oh2YNM1jWQJvqNNSY8dk9LSqSlNK0dICQ8RDfHGsY84CqkX8weDuYz0aV
apti/CLILhagJhKCddBOcEzrdAfAnjCdxsEXBSJvJ77c1M+4udAFThFWCEMmxY44x7E7IR+CE0W/
HQQPo6tygSyV5AuR1ChT/GCLM+7CJNcuK7rP0SP2/zW+m3lf/tuwAJ5TDUOZY9pfCGbkfengyt7H
G3yV41PAOdxXPF2DzXly6swGJpFd2ZstenbDO2404nPyLchUzjDBbU9k5bWat6g9TE+Oa1Eu7u9m
omyEULI9bzuk7BbqpEA47fkw+OtPS/0WIQF/JnnXkLQ2mLqX0+DGWm97nbBYztXyBmrK/FG0NTxn
bPoOHNMnLc/WhLNoFzXysR/JBAnIIg8icaorKJP2lROBWWahf3NbkcRxsYRTB8pKvPaBITWAUmfT
yaGMGogYVdzYh5y6g7mEeVlMmS/LpJhx7e/9mbtHPQHVgNm7bKk3HrpVaZ8oPxB6uOA3s87y8kcb
JRQxrIZQBkgRjB8wIThuWmORoTYy9K2+CcnB/0UINEXnis724uqqiCGGKGKIgUtzEIg+8zhtY96B
CtHiOJOCi3UT8sJOzYMg6NIcYMrZlvID04n+1MakC5tqgRuQo5UyzhzXBxCI6eHQwoTorD5lJyuh
XBL54GxDXMWzelfG7q1xd5D2anEqWl5JcNqHW1/o72dp4svjjddQRZ7NFQYdT1pKvf4vCdTPDuAc
0djuAUNYE/y09VFOggMUshcE9fGvr46zy3SBMW2DI8kiA6Rnp1ia4L4Q9waNZw7Ao0wN0kitodi/
p7TM4MH1Wmrzp8GJ8kReUI2iJLbAyhLf+NXEG55I2FoI+8nubos9E2aISZCNFFLvGMw2aJn8Ku3y
O69Rh1Q+peZfzNvINE96TIaYv0cQFaO5r4ugUKsJnGUvb/toJjtPypdYQ/37ZI0gr11wFlzLLLy0
el6OZ9ufKTOmrjEk4VoBTbdPfFA+jUiRIF83EyXwijLfBADrNDyoUC81v637xw76CfLULIy7iOFf
9Q53fPFQXIf8UPgEBcQgmM8DV9oN2ZGnKOPFL6jT1JtrNmxWTdm0GlhUX3paJPMWhiDpN1zEKjVw
hfAKSNESVbEg2nG1BnZ1uYe8fR4cnruQixo1QJmW9B84Qb76t4VcJeWSKUmdK3949xPIXq20+2pq
0MUBu984lgPNN/BcvYCMnh4LYQcRasNCVFXl94iFgv8lIUPZ475Kuzb/60KpVSrYVnpcUotv5KPD
+m6TJ9qs3Zft5S94MkMSfyHoJcS8p488Iqw8tYyWIRNF2akXmfpAP1M+3EUFBVt58PU6rnAaClsj
DwqSUPNwXWq/0AZSDcRXwF0xenVY+RtyHRxaLJUyrGk6PD+xeZ5boVdZQsPJ+JMcReSMMdsoOARt
G7Oov+byBFJZzytAMm9X7ZueEDqfsqQlbuuRvtVp1MoNEk4IxxR0XV/o5Ri80sxYSQuNZCK1C9TY
BH7CiXo2Jb9dXstD5gN8/vGBFSMMjQ5gmOwlwbcQURDaMsjDiwaXkZN5g70Ao71BEavaBZ+rdqMz
0zn+95z4Xma8rO+7YSMvKnyj2C1xvoziIPG1kLdTctVeJxF6/DjOWUDtBV327m5KFulpZiOTg0GR
D6RI+MgHtn7NARQXRRA76/l5ilACvf9qQ2l0c4q0X4zEU5JmSOnefM+zwR9E+Rqxzhl+DEcnDbDI
ohLIVyWkVkXg7Bh5DWXzALxCJSyDM4tj7AAAl/kZ9gMeeCKLMOoHjQZ5g88Czb/okKpASlv5dmt0
Eq5Q+fDZkJCetmagmTd4FC+4WAoFXhw/RB2wHeouh3NKQfRLK/2kPLiYEUDWFK8rjuQXmUzmzVq+
vVPOtVNX4sfEXI3cV/PnjF+kq+iGL5G7InoBxnbmP357DtXrdiVFxwBCYLLNL6YfsY71mU6BX3N6
ZUPDY+qDA3Z5mM06UzCItXqNghgOxwaaW49XKvPjwz4C5IW9QyUmsTRfcw4rE2Vpp0XrkkSzwgZY
JbdU0iVWOQMgD4IRdDf3LXX0+7YRo/GuFr9JOhcFjZmwVnnafd0wOAXfz2XA3GLb2iVy9ruot48S
0zoOgBIFJvDr31tkQe49KuhEfBuTqO1MKXI2osBYmFKm6X2GKo5/aZqZo8UzBXgMwUyxOOPv1qrK
Omu6+4ArJ1QsOCLDlDCUH9FEHlC+2CAbcEIOU/nYr7cabsKa7ZFe3FM76UJMQJ+XZSuNOZwNAAVg
PM4EWzDwFs1xc39PHEaJeiN10Iw786Gse3RLWvU2ph3Sx1wE01QRz0hvL7ZL6oyUOx3Q/JA7pkKE
YMK5HQ/Eiawx/zZFqlqJttwemOqbBp5OeFGvuhx05aVimCkGH2rEPY+GEbKPD7owR5ZKzbOzz4/H
cRBJhO+yxGk2qWrBHPNCg44WRO6PyBTv5K7KChj+O1qdAxnG2N5D/AB3tYOfRWl7PcKjy2D3mEoa
j+z734ERfZCTT69GqaJv99XUhK0V9zrEai6wsyAacZO9TdrL66R0iwxz8BH9r7T5BYJXZjyVZ7Ut
XSXDn5A3dmNNWA4s+ZcbbAPhOOX4wUDN4Sngn+OX4rLA6HBzsxOtfbIyx2Cm4DQU6vw3/kpzgROR
qkfP6QymEw4n3ZUNL4lrop4OHG32jP8VfGQjoAf8GQB1EWD1BKB5qFRUzzrQWTBwywgZ209klKha
7Sy/wwMgSvxPc5ug2nmqYsIzMXWYnv5hnL67bYyEcdhLjQT2lBZtbtkZHllunC4KAgzDLIrKPYgc
yO1U8aLPCUcS5oQxnwF7mC3AwWly1pnEtuzGj4iakzvlCNHX57smQW/lLLWVYCA252fhZ+NFiUhG
/Il//PNYpWoL3VNXpkuargZiC3X5fCjn9yIau4wcspW5QlLWomQA7oG7xBj6DTiaCXJ0BUtZmY7A
db0rz9+Pp5L+GJWn/FHXrTS0eBFwOZL5WrcVtycKjrsKxY005VhJ1kVYtR/xuiu3vL0dIuNPoPQJ
kxu1MzOF8/s2djQdE6MknXFJjSOIyNEzbHh01g8I0V9kwLv/zQP/0Ry0oBJT6K2EygfOW6RRIONm
HCcU98YJlNZZZ8f1dv9RN3VwiHuznoLZB/0ROXVNleRHi0C1uXEvUhmWyFuhLfDDkayNPVrYibNS
2jPbBRPEGHrLSm+9VkN3s3CXlVqmSmEhHV2MVrbpgV9eLRReEVGap7+DnYKKMYVUyh3jjx6NHrZy
6jcOrrH+yEzWkGNe1p1LEPhkRnaMAADC8R3wm+dRm2IjTn8np0tO7jh0Y/b91teTCD0LdME0VbyD
xJvRICv9hVAx8QYl46aDbn7elh7g7L3MR+HKIF+kniiZ/TaW0oBZcgviu6qo/CwPZ9Jd2nItclGg
zIlGuBhCttbeftExK19LJq73tEP73rBJWkHLwM90bjp6gfT4QvcTDs72+jnrL23DOSaJ3wYqBU9T
NmC56m+hjSqLz080+xJ1Ky3ZweBVoOi0NWrFbs0C55zy83WFngRbGsawZ7lFkRJEspFVn9VmA6se
XvlJzZmdYhzEzW5ftay2wCG7d/fSvOKbZ6Te3cEUgZW++LCgme7MLK0vHHeZgbk2dILmOXVKsucV
oo6ewhTvqASXXaP7JyEmrr0bsINujBrzF9QNdMEZjuIFkpWdNJp7J3Otxbz+xFwix1s5jcsBRRSQ
Hbl583L+mWoK/K5vE0VDPhwJCcFjKWyzPQ6Jv3wbc0zpIhqO5doedueTBRVRubNLYI8JkdKCS0tn
gYucEjhx1VXlpPzQoW+MG+HnOca4JbZLB+Bxyz5HBh/GHWxQeghh/ZZakcUFqRBjxbJM/ytiXEUE
Abz0xFVjwzal1QYXcmiw8GjfrhTJsX2p3I6gn9t3cUkimBHRURk+qTB9eSfDiwmkO4Vj7xWW2itu
CcfPDy/nyAu3zEornoMoE5tJUEtAVC6eyPmRSNKbUPWPzS3zI2gUyhBUf+Zs4knguEBn8RqRjiAm
VGOBeCDKJd/yD/wdQo08vTyRV7OAgb31JAfUhjugYe28w0hA88AgPLC1q+/R9qpiw20kUVr62SmT
WfwPTIFncciw7PwromYDp7h+o7LgV2HtHU2sG1LAzOVT0Mff9+oQMXIRprEPbmIQCW+mBSKJTkjp
/6oB0M+f7yxtlOGxV8h/sGbdfTashCwNVOYeuw3Rz+L7mQhYic9t2BDCELfLHQa//CfBWmcqOVez
C0/kLYwPM0wQevBrjWVDx6T1o2rcNFX61U8etDA5lj+YKZZCNcUpRpEX4+tSlRUMo4/x1czJz3pq
nN3hAwhP3pKUya8G25hh1Q+N3Ku4Cq+cmepryNb44jayiba/LpWVvY3WlrnnKzBuB4W1cwJ3iliM
xIc6E2aEMlJBrjocKyraY6OE2IhEf2C4rpPtmTb3fwPT9RMnkfgWBcV/3jwQ5zoU4z+lk1DtkW3w
L2tPnLc3m/Y5UpXvjXREk/yE09cnJM76amEd4ZUBFQYu6+X79ynWdPV48+uqfdeuPc7Bfpwuxp8/
053DFrHIf+HnK+qwJPa8fG+lnyL7b6qjNqIX7W7Z9MqFHGko+lZ9c+A4lsktpq23oTI/bwcGw5z9
RHu1u4+rGU0Nt4lInDdQlImgWvabjnlWLw6tzMoge07Tr0I5/Dd0nZITXJFNFu+t9eNWLtga/OpK
trTf4+nF1YgULIppTrFgsSupg1G5tBj4ZINzwCVkcmxU8Zut4zC6THb4hHuU3jBtfD5xNq9DhjGB
jX9sX5KQ5++aqgNjd0fhgX8idJMcKASmXfw5VbEjfZcUGAZOWvXNF+ZdHO7YCWLhxdIbYXEGIgZm
yK5/HMgJQ+Nr0Y6MCWiAk9uP55rEv5PYRXWyktuXFsBRVcvV3QKJnQ1dy7oL+i4YiUw/mGm+w+ye
1WZjRoMaR9rFXPzDfQ4HiryOYIaK8vbQCv/xTeizFxzfsH10ZOswltlsTYcZtVV78QlO4GXcKkfT
2L8AS5DETZrOObkU03FtCF8wlc1wcXZ0ZQOEZesxYXtn+wuwmwOts76ySy+EwceySG3LkmgCgIj9
HHU4/aG+qHs/Cewdx8EfkbfTFpnTVtValTDMLfIE/r7s5+xTZvyMXYKNoLnEFVMpNwFGaElDtNTb
KDAoGP7bCIJmummH4U8Id3l59yBjCOBansa/7Z+srlNFxoViWKhdeYqV+K9rYk1dp1sxPt2I1ey7
UIihFN6TlH/9xG2P3WN97a+fh3Q+tBqokfTu3KBbXpSoxDl6UBSciNQKvX6AZohITD4dph0Kql64
4WYh3l07aInAm5ZGE155fk3gsNVCwnOwg+iCp4qWP0PHJ7lYHak6xkMUl+vFN3cce06/YwkZ5tOE
R0YSPkSmfGd8lGRw17cw6nRYGuujALnyeBCFUwJXvbkcU8H8wzPnuQiXZ/kBNK1z9+6Rqz7Okl/V
srhLAXCbxkfnarAuJlOCJK+xxL2cm6LI4Q0WHNtnGf3NiLCvnloEFiivXcuIaAm+gB2N2efJtcL2
o7y3q02RgurEy9xLWwPOiouhobIdaDq6cUEGD/sOzJHtCIm5hKjg57x0hMENax3iYmAAXcGvZuLY
P9vpG+9KGh6sgW38BMXoFE5BOc3o8gBjdCjnynV0gwiXW8vFrem9fJf6mcdT1bd1XCv1ooJdiAez
r9GQci7PfhmLAykVFNdr71C2rBLL/ods/UWSsDNzqYUswEfV8vFvPTt9zGG4NddKNH6M25LfEY7g
+Q/bZqjO9eP1VWkdUeDvWN2d2ymnHqSMn+vx6HmkhXHRh97z7VCTDjkYrBcChT8FT4S6y2XJZtYv
DGZajzYF2v4O9cnc8zedOm3Tpi8W4T4CCcVZwqxfl1rk3XNNjBtcB8Isf1yQcOu2Ug61BJjt4c9J
JT8nHOfeIP0bCwUlneFLA5gpqv/sX9x5lb01nF2yH5X7a+6mTYxrc9EMfgSqNLIep2+f22HoVa2s
QSb2UBKKuC43YB1fJtRrSlf3T96tMKPTG6Ch00FqNi/XZ5S/IHAhG29+hp7l5p+faV+6XWIHtDdm
uROIen5RklRf7hbL1Xlkn6/ugos0WaUvqbrgHf2DiMlOaz+2NqcweKs7bX+2ucyWwsU5tRH+rY/g
tfCDuojmLTprQk8dL7zHS2/wWIzpf2qTLJkI26zOMoL7ezvNaLoAeIMsfbHWIdnKyvjdnN0snSef
J+Y4A53m8q0iYEqwGFFSC7qEUIePpD9gmyawa2zGkiqQSZNczPVDbQG2oPKsMTF+FilkMlpASxz/
F4cntPYBVQ6bZsyxISdld5XgSQrEwzEz+sTve3UjC1DquazXzDgPtXt4m4KijWpcDqqhbTSebkbG
FXTjCH5pMu0SFg61TDwF6gM5Th4i7jx9tSfujci4rw9Y0wlBZn4eu5XYAWrUm4khxPvbLsTTpyBN
UORPP6YpCIZtkuw+MLWbs3Yj659wEmByxN4W8wH4dHgswvYv07KT5rxMxvEBJ4TtZNW/PhmDUrXO
Gc/eyurP8P97U/h+SQO3Xpt4fqGc4t+25UGW3PGstjZXaympXP22qS/PrBKS7knOt2iv82zX7iBD
+nZkm6rm/Ir3iayxj4LUGntNGq2sBCwS8oeaf0aVhpV4PhlWlrs01mH/HLNjIfHKZehe4xWnMOC9
8tgGc/8ndtdD39D1ydC1CjRW4ZDHalqK6dm/FOD8X6nkBQxo1d0nSCkW+0AmWP8V8xMwHRBTHE1n
7aX8d0D0BO+AcTDkeBWXY6BomgWDAOYs5vIrZz5QDqSEO6rVr89HBELPwhftb1/dXfmkBcmTqZzd
2efBfK5q/Z+ZRg2EGvr3T1cE2COrigTChPIXX9EOO5v9CgWTlQ4/1aKUCFlGfojYNSY/EvnT7oGs
zNh0ZZXRwU5M9YgahtKnWKnUNo+fDtSGi4eV4zHSzyZzsRW82ieOu4/7vNNqTJkWv6SfNtWpBdbw
HyOykyQW2UzNgzNwbIZ3RQdkafgyZupB8JdO9JlwyH4opuJDxXpDW7qFa7zSoLTac7J+WGolj/RC
KR/nVEOU+Ej5TZdNJXeRKyVY7QVZoAlQE49oevdtIoGu5ZWZtH6fzK2BZprQ6ng9CKspvdDRuyWj
p2ILGPaDSZRBPvsXFUMV35p2yxbTQpB8Sz4r7uOI0/bcKLVDY5UX+z3zUtsvu1Okuix8GI9Osr9U
1HvS2zl0K3Jhx65zTNa5aCbKECY2hTo+qUj/f/KO53PykImGc8C6EFIpmJc/LlSsH1Fi+8yWFPhX
7Kz54wfLk+N63eoza4GMC2e2Q4D6+5vQUfoSzYXpKKsDryA30vUtpd0vBkK5fWKP4pJQFo39sgWJ
9Amejru6CsOvKUhNLs3i8LBcC0+FjMmnLGwgaLqZMOHS3i0Zg46SaYuo6OUPyNhzzj2qDY0rKSGJ
NiLBLdVmdhSqTDKpb/SC5NdAraewq3Pj0v7evJF2yqgG9eRxzs7fff5CmtH9+mfaxxEPXKBOVPQ1
T/g3c0o1kK/dGpX3FGwKO1z0BvprLnkeC4/3vPpyA+Ry8KkOPaKT01hFpctF576p8BrqsdwsKEFi
kV7vSFEfHZH+mNoVU8P340b8AeO4ELXUoVUAoSrZ8CVrjpfmGxt18Vl1yIQ5H55Ny/EvlmFuFof9
Jodb2GnPMebeqfOkgEuaIY0ZejXSo+m8QFAGE0SNSgDbpXO4lfNTPtKnJPxPBePjshNLe4JX55bY
83Va1XXW5kfEHLXwGKBqhQDTrY61xg/62NaZoRg51aEAZBWIU7JCQMG6+W9Gz3ryVhe9TIrv/9Ou
SjsKtazHYQZ25qZfx2nNEUfr7XSuw/s+eA750Sm+1H2pnA007GdlcVGvHnHsCcfgu+fqUABnPDMD
vsbxuwogsp007zRUFJcLq/eJaJEZTQ316Bd19MsJa2sAGTaZkgbFCDZ734zqlyEubMygSG4//7sh
fo+yfoH7qMDxX19YPeaOhABT406AM6HpArhbGfYUchQJUX4NGLQkVR9ms9Mas52qIXEcJqpyxfar
OZXzbFSe3+PVOaoxw9B92opH97N6e/2QjSnGWJqocnEb8BM9ZUPD+BfybthwrfHkeMcpoGQyaA0Y
qm8pEtY1bUPzGPxk2voo5nw8MyNc+iTe9D+sLJdaxzcQHGauFpTzk8PebuAFri30EwEOSBCZ11t5
xaO3Z9RjhLLiD57/A31qt/QuwKoPgnYnMw+dBnFiNxORFMZdd2NesOi2jbxpecum+ovolrc1QfxG
lefNUole/YxeqqKzJwm8sOYU62VSUMOw40uR9UN8FC3ATuFVP4fcuC4VptcemStXKhMwGuffwVGi
TTNFhpDVaybNEXh2gJyB3Svs4msiacLqpMDipwPi9C59MbbtbrcLgtwHi+cFVwXxQ9JfIDRkzYAm
Vuo7DXHQvwQkNHOkx8Eu0ZTIhSXrvU+MbWXkQz5xyaHy4u1gQG+c6sDy2PY/LZZM7vVWUwJ4uoL9
hhzY+dzphISl20vicTSRBVaL9xM59aWaBvx17Ly0NcRdouui9wmYJRYe2EUeHCK10C81WuRK99ar
cj+claoHnH/s6EjLr7BXntiItS/7fdSCfiMEQtl6NIxnR3wuckjKahyTGGsXbYMY9GYJNBaKvDw2
dQK+APQY/F5P8bx64TmrE/CcXSPGKK+BcKIgdSxDSti+xq51959Rpt28uNmkBm3ibFHC/5dgKLnb
lJEoWU6jwd1yfuONAowy1HoDYC/ZFBFupz8z5qZ/Q6JsmYTExwRQh3PIDPyJtRETzflEzPxloQ3+
b0ainx+F45iaF+LTNKHLlyvj0NjLhqBIZBvuT8mqb5CicZxTZbdxmDxtyfzYt3tcscJ/kpsQurbq
qbuFm5Yv2zfjUnLdZ9dpaPrF6/DRIsLCo8zCa1pkrA+o5AvgPKw678ueu3TPBRQap7LwM3Vy0ASQ
rX65dzuEwMzfpKpFNAdV0tnzOHmaYCrcomgrM2Ltw+c5zy5t8z5z8vVCiS0GrCUHkdYDnoZBDCfm
ySh+1xOFjKSRVZ3w7NlrIf0jnsdodBAHAkAl9Ws3Q5+XABziTufHfAa1OwzNKqRhtpxChi+xVJQ7
bb0+xyWckrKWHzf4zSskgZG+5Zda2AHbMAFeYs/nku5L3Gh2fHIi8wJRFUACxhmPk19bpLklCphk
e2gkaYvGwfLuzIfmEdxK3xyuKiZ65FP/K3vfFuC+emFxZOK8vb7IAz8wim/GJ3MZpnTw7hW7SQaX
DCLYz58FKWeE2RM7RMgMo+ScadmfxMZfNYsAEa9lB0OBSLC6YOSuIUt6f1Pvo1xvecAxT25+2IgY
0CkGco7LuaSeSQqDU8gfNmVUZEIHHAUAmWbPk6TSTgrBA00Os9/uY6hZrtV7BsXThJxDR03Cp3Pl
VbQWtUieuJT1nP3Jxqba0ieoPkk/iJ1BkTZh8Gl87DcnpgahT9hU35ai+DNWwVJpA3eZgtcNV1/P
CI7UZ+YyzPrbIWbLWe+gzlNMWGfvf/dPrfZV22T2CC4+4DSuQZ34jLcXWbpd454TPsrYjYWO9hHp
UZ7453v1NF0cdBC7Dkr7h592LrDz/1xY35LZd2igpQmmkzYy5+BmgqeSpy6p7rW/N4UYmbRrIVg0
UvxyL8dZVYkCLVhdfoabMGSBlSIWwrDSszSO8JCqpM+mFB69kS/MMpnxyTP3ezOraaYibgJ9ztLf
yM0i7kzRzBUyRURhnk8scH6RvRXsZLqUFupPgU64w2LpztpPCflSZMk9VByAyFdXZyxQS91CaWkq
V21gMve+XXbfAHU0docrviVRjAz9O4zs07mMi5uy95UM2K55AMNh7x+m74w51YBZ5cclMiNLV81U
FrFh9ymWsYgclrDKH965qI+JLsZKPh49mA8BSVcLOHvF5jSeI9WYUTdC9nyzuqUSgZTAoRxcbrTl
a8jHxEEC9qM1VC3e1e/c+lNPdIOGl4KX2K6cXutBZVbKp0r8DSq4zJSMRQ/C2wYCDDT9Bt3Kvg+m
xHw9udyC1nNNcnTYgC+TxEMHn/22xhiHVRJRG7RHZRAVilkZ1HyztxyjiZsMDdUNR/+puoobjfQM
xPwqbdvzvCzG2ZpglR5uesvhvMI/n4ogJG70KAKaXCf+r6ZIl43UZ9mXipNKsn1Qmy4LloQ5+PSd
MwYqtaKsKkaRtRnWZdeGNZVxzHAZutjChuhoh8IbMzHuOP1Nm6mwX+z9BTeUarINPqQSIGN0ZX0e
yxzLCcYW6n499H8Z7teC+FNsTmPz6oMpKwxLRxbRUgKBMEqE6Acj4UnRpOXzAOjz6BLHTNZDHpy7
T/P41nYrQRCQ8GgknRoWh5kf0FpNwoYBV6tyZ3PKHL5icCBjOz7dp0OWGPU1IWn2/wfCSdQtQZnj
E1SNPd2LC7iVdpLLUXdUUEOr2tAPS36JCvFp23wlzRiKM1GKGO7mi7bmGUVWYA7O6fpGbBYUMZlc
HGz7FhKNtyoyY7CICJE+LbGApz0oJ/+oYRPDC7mJ1Si0yqyN1cbCxB47Zi+tyJtggwjiabkdcDdR
qw2utIzUtoqiOJ5p/GY0cxQNDrVTeDMMV+BeULzOtV70X2jo8M0tKgnRs2S5GCcp0eOXsrN7urTj
PeMQh9tPevlbORiNLRNOOs+PQ6aeC8YFhTNYC6ECfB1gchkSO2uAAopUwIFwDwoS1Pp4noAFnfqR
ObVibYv4QcTpFweuLkCs9v/oRlIdJU0vxwytYDETH+qRvnIlhBgWr9Yd4Aw0OoZ8xczzouVoEXA+
Un4vq8ek2Q4sVXJNO9mgvnV83X6gC59if1lY6EdQg0mK3OpEixEAWQFU/cMOvSeSq5AVqB88LOfr
gsMcCnzSXaJFmzJITOP6hv4U4uiSjJEtDvQ+4/Ov3tpfl+DtZ2gb2sSlljO2Q7tpRTCg/+MCjMGm
QsMrXiD2+gzrlDk6y/27E1ne4ep8A3XQDKm9PzNgFlVRog2MO6rs9nwNSMJQH5l7Y+FiJPIGMtXj
a0kCSlaOtq18/GLr45fLEoePgykcHqu8RZJOvh6nSM5ZCpzowkDqBXlZm/2FL6c3aqOD3scBtdpQ
97R8K9VwTcOB6cLVU84IGO10owwVieFEPlPhARo+lq2BLycAtAUNg3ta6EqAm6pq8/h6MmFu73QH
fuuWfirfm09odRCAlOBhwM450LjVjc3CfjAP+KsLWBLijQPqpcR/w95/zuTW9hwsk9Cgx+O2xSNU
7QF605mk3gSK3QOzIKB18EriGQcJCZxJ/7nTXkeZ7zSA8tfUa7RsVHlJIaAYotfgdqrBqSBqYQpN
IsDVMEeSl2s3BW4KaNoEeCycnz4diBU7Sr2SFgscSI0qkMLkAi3eRoJIfEYGQB0gE1Jp6g69w3sS
eD2LqGjZBiu34PQEP9xRf8bdXltr8CokuFnpz/HaRL5L2aaPP2G4DBzCdBFB3++y7HkM5QVpViUA
4dVpjgRzs5J1gndpk6JA2oTZMzvduVD47ArGdB1YorppfdR0NUWTugpGngnKsiiO05MLu2COWs09
w+BMeVrUmJFm8MhIXQ2iAcN93SszeMTUqZUqOHADto1ydYXUGkzLN2J1zz7Oeq9YZbWLoe1z5a8i
/pFMwJpPjgG/ZyoP+FxDa1k+pqEZAxSTzXvwY8fcoF1L4Tg1NTMi7bKnGT+pWj0T8mZq7mPjPbZ6
gm2ESOnSajRw4baN5wsh8oQ3fWEctKyrcBmEiccP3c9IVaU278OsQLtUs/5XiyOG6INRz5TUn18s
BRavUwsYR4Ky/NnhQWb9GmjrA0FopT+XK/WOQC13qIu4AzTMnU4Qynj04eCrV7EINOdkfBu81PzA
evQhK+/Qwewg3X2VAysXwRGQGnSRpCL7ZLupmvf2PoCa39h6lVqgBjP7eyRJC6WIT9H0SzFc/3Fp
64uGKpcg+xp1rP19JeodDO/V4/VWIjZTZkxS2qYckygHV9naowmEeFab/PEkM+jsiSUBy2HjAcUT
6T/4aiuIXQeIsCknG4kut6FSRY3C1A7r34FC6XYUtaukGD6eqtZASMweJNXpSFKLmP4SzKV89vj5
6i3jOnMlr31KQE21TfRACwFNnRqctm7lB5XR3iSRh4tGAs7GPwwp2bD1B5W91j+FR0ItMA5RwlsN
e0vT11kXL0ID76S+T50BPLItLayvgVn9EOz9iHL104KByRX8eQF9SNOPdyPJASjVjM/h2hnnGar4
y7AXOYF4eHL3RjLieC1JE/wzItvP4BuS4PEwbsG3TlbN8gfFks/bds4XehGq6EwWP3WkWhPq9tt4
T4YgUgy5xivgvgQB5G6q8tKldSPg9R3F1qCVi1/J+I/bLnqPgKpC9TN/wIQe5Vc0QferU9ZLa4ty
zGHZHVlE9YNQmJzjP6CL1u4e7PBI0R/ifewzsHXXknAgQccTv7yLUUZ5IovlhnYqaCly+yDI3oRZ
VionwhO1K9v4etmT9m11uSozTTvSJy/ShbUz+1JKP9p+bj6mt+KnGWWDlZEsiW6rZMgrZkjh6S8l
CXFKTyynYLJcdonD9wR94WheZ8zJ5bPgC4QyZuYnK1PexJOmImAAbsyhhCTejQtITJjYZp5g8LwF
utl6uZRTNXCyRAb7O2oCqivdk9+MEtRLPA40s+cHxf69GuNPAnQgyh27pGgJC1Ai+By36LJocvO/
IYdAMTv4VVtWvNBBuxi6Xhdyn7TSAwmcArYEzPM9eOmgBMyN/E7UsjPyjeTNN+aeAerEcVIpW1Vm
ICUJkno2a8d7BkCs4xm0afPugGuhtKWVOhL9+LUq/rppoe5kgTt50xHJUIwnNb402kNW52xH+Xxn
avl0V7LNsdWHXVm9x8q8tzkGfUEwo536LbjyF7qWL5iTzefY77YehVAZOQx682SjBpDhq+u/NSUw
A9brE6jKoNU7cIildomxteqtPlXsMagd7XkbpTqZjDR64sDIKr/E+sFM3N/mG5R1siZC+TRVQ1uR
zJsVsEBsry69f1e7MFlGYVrzOWLud3Tqm+MbmyR0vsKaeuNqARRNM8U8486NlzmbfNj61j1Vhv9C
NMhCpFdtgs0sEky4yOsTuI0++EiurdJh44ScPxT+KsIc09gZaOTTaQ1DP+nqKLRQplP4S+UGp6Yf
zQEXLPci9/rKhTTnLGV9JFi+pOSStSoQSFTmPSlvalL9MJy8QVAOREHfFc5QHdvarLu2UMJ6SOcu
TRnXUw6ku+EAAGhNDDHRBt6BxmqLh8ktEJAEyERaQMj/Fo49s1Q6xqLKusAwszssD6AuaHJv4bHT
ay8XFlnv3ffvJT7ONPHfiGq52uQ1hC5KxZBQYZJEmV4czh2YfA7ITlFMgPMJviQjz38SYtC3IDul
92SA/Q+kyiSTPhOfcwpRYq9Kle9+HbTWbdudmWr0HxK0i+V2PrRGGuvZia9ezq3x2fQxGkgcGMGb
CqsYVWNS2HtachvGclYFb8TV+KQB7iVUZ14Rop5HZxxEos69/wWm0OWCosWiFy7yT99rbsuAzTD/
SJoChfxKwMEmjdv0IpF1gqzPgVm3wlh0VGrK1Hey+eAaSlrzjBNo8yW+VuO4IOYK4o+9lhm9ftUW
QxJg3n2jDGB+CGNY7ed4q+Mip/S2EJ+x9j99Ox9Wpv2dM8BumQSM6njSEQsV9192quLoVr7O7VpT
F4rR8e5zEBUzYQf04gMvh5xMP+kJpOqcuIBCBmufiryPOzbaoJFazA/P91Rtk9LduEDgbELO53Z+
ZRVJ/7eqJsCEryy18cq3kGxQtJW5YQDCT7H5IDqKK7elG8W8M2I2RBXAd6b81+iuTAOpDpztxaPH
/X5NS+9CJORPovoU1Zk3YVj/tl3YmlUTgrS3+6TUEXzpjSlpXcB2J3P7HFFV/tUpHqLUIp9t1Xau
L79WWtP6pYfYe5eN8UtX4ezgRcunj1jQBpLtp3RGCuYHY1dvkyMhV2ut+VfrAF+EVksBpLmIDvhw
o2YL9S1D9DciF2AvmvsDQzsaRly0x1lL5KLqFCpfMpBxZ+ezC81bIHum5v/hs27bEnL5xY7YZhg4
2GsQb1L2HtPd3/NIXigY7HSF6lcKtxTsklWdyH39R6fzOXfFTlueTZCHW0uIyaKHsKgORna/kbUT
MVD2hD0eL190MetoPnyrStlKDFZcKJdvSrD2m8Oht+0Waeu90WR0w0sP4gineIoIBGRniqiyLkX4
5c5U2hHQyaARi18yTvYUecfLbASJSKcztTFYNihxGhRfPVlS/PcLzowhDMpxA/QTuOe+XSkqxcje
zEMI4bGnArcACtTQ+pGIXWOPi4ftHQTlDL2KTizun///JihCSQ6vqF6fcOyu+J7LJxm3pzSK8Eph
o1Rj8573JGaPXNFjjfEpaEfW6qfGa/2/e2Hfa8JTSakOPLRYtf01qGefTzobFmWL6Q1Fdnz1Xl6y
Dtky1W50VMICV1A1/IqJYCgs4VUMoDa44ShO/BEbKbUMjMrOZMYiio6NI0VTltc+OvAaM3W01kfW
fCMbu+yLim4Ad/ccE3msiieiw2HJD+K6TaCRYq4vGlbmRA0qTyBO/Z0xnIhsCeSkzwICHr32a9Jb
XRDTd8wP4mjxdUkKCWxQ7vLbJWXlh4VAF6An4d5YI7pyWFCMuK0Ps3wl5Y5UwNcmt/kF389LMGlz
JWMOKvg7JaPFbY5dZqXY5vWZEuZrmF1ZjlzZNE+fUv8Pt9FXDYgbtsQ3PFy8m8MdAFPuIKtGph1k
zkoqXDNu2sDjVjS8vAYXrgN5E2UbjiD3Y75tATqgq0MQeaFSgQyjDzCvmeMAZBXX95zOFKd4ACU5
+UbxKnu/bnPaGnLe9cI0cQDTbtYBdHfhVzM7wFwOM5RP8ZISLJbw1ZYoAtubuCJH1LgtBwEiro7g
7cGAag6JdgG3Q9mENRTuzYldlDED2vRJ29dGpcON5f5TwpkrlFLfs4sM8ypXOw1aF7PLBwdooa3G
HeKFeVKy4zZOWONhC1gXvjQtu7GYtOrnpklF3jPdITE18sMdyopKqmrRgRflUZObd4w5bzxOb5Rf
z3zQJpOruzFkqXYCL7+VQG4H6xDhDYl76WmgF06X2DpgtQYiW7d5++UfmFvIkkJTFGmbo/soZZDJ
T6A32ZzzwIMBqcl/e3Zc3B8ZiSEVxYHxuCDGBYS5QewzX0fp1z5YNtw0U/3luTwBvbbze7gbng0B
JkIE8TNNTDhLLL2nD49dwf+J/dhjWnOlP/lq4rcRmmaJ2MJJrOBMTiCO+hsO3ReZ2MI2VRt6oGW/
K1HyKdeYZrZ2k7mx3FpwY0m5htPcZ6jzMrKCy9+YO+O9uLfOLBiuiy5CVWqqi7GtPGjPT4I9wZWl
KXJ8Y2GIe9hZM+AQcqkoRQ218GpOHhOfVhJIpUwm0Tv6NIc0600VpyxyCamxGojr+VJJhVVMcGMk
NEfIrTyhG7EZGnwcsfNPxbnzVmXWOXjSQa0VsQku6RhSGh6Hc06x0c1lR/R2Af87NVDvdnC4OBQJ
lxRBizvKjb0ITZ3hA4IJ6g+JiVTXgr9GXH14ZR0KjFRi150z22aWJzXLnWEr9JiykqM5SxvlEQBb
yc0bJPbgDXXTydq9R1poICS3sjXUcTYo9MvrBVlNky5KgXrHsnezeQYdebgLhhm0NoN8kNEkDLiz
0ySK379iVrgSZyzWM/bRCymIoevaCet3jtBiNZOqSHQU2UC5v9ifRxBg6WJQmEu7pkAe0doUIvO0
1Ylc6GpoCLS0mNMrIrwZvlM06XTKNtMFqO2OfVSF4Q/grMJc6Q680ejJYHy/deAnDgQdBfLP6yEc
zV2XoE+tsp2cGKnQY5yTxriZDyoIsFW9tjOaX2QQBzy7fpnvrFfuSkx0P+6tPlsm+o3sWl+GgS2D
W6Nv1F7WWEcS5dbejEAjcLqdfmEs6AlBy3wObTUkCvu6KpnSaSz9YKjKTSUVWneTd4eER6n8Qw0w
+bO2e5z/pDY8J3btsiEOhqrdHYGP4SyXPN+G6F4IZCE1ocqYrjj06aB/ooCIhOM8tc5HRoNB2rlY
fwqTmaGbSU9w/6lNO8i8OgyiEWpOtE/g0IKPiKtNWe0WndL3xYgRzza3/d8X7wVXjb8Mu6eFkXiS
TcnWR8puyk1xRlU2Db9ZqCa9VSMwVZ9EPAcW/Semeg3N2X24EWDppulPH2eA/psxSFlKZAInCn2B
PbCARLKGwsZaeKaXYVJIBcmkwrT3KL9LZ6kZ99aS1G0yHeYr1Z4+EIIqZBnD4EolFtbS8xQYxV9q
lkDb9lyxJiXqPHKaljfH+c+Qrqw85HFg1FaxGFpvVxlcyvWdCD0+kAD9XY42uVIdKKpNpVVnOeoA
8opVh5b6Ul99SmEKaHe4cr4E5rRWSP7wADGdQv+splisbyc44yjceUdRuL511VW4z/EWaiFpf2uu
YHtsFs1T/ZqehpjHFR+CNaCZWIx/7uEAQX5brHwcMU2oq97aN2WHUDw8Lfrgb5oTo/PdSMtVHAqd
4t66SYe3wvARVd3VwNX/bEtoo5bM455UWPy06kkg528amalU8GgFd/MP6IBAV5xfypMsUlrvpyFx
4SxVDRbLKtAticmjKMSQ7AAATanEb9j5TusGjtx7zNePsU5+M4QW9ePQUmmW0dwApQUWbvKNK5DD
F83h1mlVuG8W5WWrzYGtjLNZrcl5WZh0p4G2Bn3ZPp6ed7U2x3twwEv1jZRZbnRHlEdA0UvFS6TM
9wlWVIdX0h4Dnh6sAJcO9OhNk6btGIr2265EY3QL0vyV7intbcTwrVzv4NtfQOmw46pfkWDPbeaf
TysnZgk8yu7JXpq9wWkdxTr09gL3+6ux8BLk/twoi1USIb7K3ScXrIsu67uYncGIhkef5uwOKTX6
lzKdklS8jMx3M38T9dUMcB+KsT0G30Pr+754luHyIs9ugpSK/Hwm40cnzTZabpVglIh8zMdGFVBv
unWS158y+EHa1pWumXiF+b/trBRX92Rna6aHtc+tL2dyIj5nHcbMfZBupl8ucbRt7/bEhxebFc5W
Xm8aLemUkDzFZf5h5Gb1iAe1bOCXwdYOGcb49ulH4se9VO6JGLvl+So4eQslr8TRyxtCbmy6RJ7s
QOC3L0G5DBOQvpBMGzKRVPc5IFVIisQ6SbSlnRsHpuA4r6YsxnRL4bslC7Vrbokp/kEPmzTGwKIs
mvZnxu9T4NixDsTQK6lVg8Cqt1wILvkHWB8agabHz1LSr4KDDaLDGjG0Q/PWHfVi21lsTn0e7QA6
IEXRVHv61G8gMCDj5zhqQmL6I3r7a7VJDgFP+3NaxNhoOsVTwTMcAu12Z5O7N/U8uJ4HGN88XnN4
FWNjPMGBaoGcmmWnhhDrlZvjRV9M0rHgBak97M7/57GRDOrdaq1k+owUfHFn9Wv1WXZupdJPTxHP
WsORxqkumjmmc1yzRGt08kjml5/PFYpgDgf4chpH/HMtg7qFHeTpEaC+Q1gGWF4GlROjN+zB5aG7
P5smID3Kkv75Jg0ufClC6o+FydiweyV09h3O59WXYbCAXoj8UkgFFs21Zd3fYHfD3AeLf/oGYR/L
B7/l307aBy7351ByS8gh72MvWMZE+3BRjPaeNNrUpAK7+kQJZz4VY7UfU8VS+fJah2GrMm8/votr
kQUkBYkxKITlFDEqpaqZGxGlyR/Pnsz18N0ussPqd0PA5gKiK0SfLy4qBAaewgOTtJWLBYZT01nn
Obah0AYGovUFFy3MP9hJcq1Wrrrac5P3RtrZN5eP52CkLE3ue+8iEL1ICeIOxyKhwD27p3AUabDP
xfEaKXgpbDqWlaDam8GSBU6VpICpKKQkRyiD/0gnL+KPq0Qr/49SGosJnb/lYc2BaZkqqQrcnQOr
Kkd/Nxh6uRAs4C2A3pSsgSpA4uBud2+DejiPZSEas4OthgXYs4xtrA57wGwxxMv/6gX6j91ARKSR
c7E5k+IrCE1AnML5koH9lVEJ28irHksZPUZMdssLeZKNP11parc6K+Qw7sRoELM2Vpd/6xhuD75U
nA4WC44utkwnzNQVM5qldBWXLDRKdmnObfxPHLcRP0BV/MivPmx50TLbKEjXHhiywe9wHDXJ68AV
gXOHiZ+WyCK+cSS6A9FkW24PvlShXcEvc7XaRFz7WcUbPE4nmmKZV5xcJdrUkgKi58G7/vSbg4XK
QUvtA3pFbZ4U9Jv68gg9EvcE52ji3/R6tOfHIzKrVq+DYfbaEt8nKqKekl6dq6jcQgVSbe08sZDl
q35x10G//LB3CNBGgyqcNMIT0Bwg5OZ1Nrb/GcrYCRBwoIt5iwMibC/ltp9FMToL2YqWK64CuFje
y/0AiikoPdMog0JUFTQ7FNJIX4S285tZQ3u/0WTtuGsqbWldSBHEqYGkye+vYmaPIAGwz96RX48h
r2zYm/B1tYYWBrFJR3UDQtdDDXFMnuLlDCZaplybqfvWuu/Vs2JywYv20YFFLiER0mYh3jX9Oxjb
PQpt11R9oZvivOaBO3Heo2zWO0hRGFUYUxPjquxUeUg8vJAAkjs+JOzsnTb1maUhTDMax3vH+RzH
EX6yYzGvPzYKm6smF5DCwaDOc2QaXGRb1FecrVHSKtqUtohWWMqiFoi1/C/tq1e7Unsm8yl8/ZoQ
Ior6dl3yIXke2jWU2Mzwf/ZjJl4p6HPqV2Ff6YhIRtm1D9BLtzMQktgOiUbD5gvodCkRDGXpC77C
zzX/C4127Lh4sAkDtYdgrL5cXhVJuVWAc5f/R/Bg6hTGljPCYO42NRDFm5nuw2pCFdEVYtdCWDjK
2vmretGPrvagTBVR9Ya70W0+q/EGzG4LfME/FOPD+tUCWasfiRe8bPilc4OBi0oSwaezkRX/yDIz
DD3ZJ3gAjjTnTqrRhSCScmCe/Znnp8xOFKTC4qjFeMYQQbZlYK6W2D1JNpkNtcDb16zjx51vMMqJ
pjk8zWQES67L46g3FTP4tWRDwX96H/na7hqi7zI96jmPCiWBI9ZgpPpXHrP0F5wMHpU1QqiiIbS3
f8MIP3tXhcu8bpIlM7ZcaUUECy4Oxko48/Uu54l8+qqMYuZ3p0Hav8Ycia9sB6Ad897JWljvztAZ
fXUW+CT/zPaUK1LNFpC6g3+xNqJKmox6KCA0BbXcDehqdGicR3M4Mg22v6Fn6be4EL54p65Vdw8u
c2BRF5kqaOz4tBkn9RCYH3NO6a46ywh6PVY7q4OgFCyDlFv7aMpMkVeVExZAw2xeoAmIQOTVO0XL
ulAwDBKrGG4DDSiBuwI1g5acw0Cae8KwBYncDdf4m0Ye//+5U9XRsP+DuNWsWB6utQcRm2DaZAo2
WqIOkcx5dXsfQ/AK5PfiISsUJpv92EQ3dkNLsIU/lcAc6nXARJDxod1+agxV3NqwBQRZ3lHUzzIw
72r89YrzEPsO/k/r0kYJjjuqZLykQwTCIq/e1g0IOzfqy1EWtlkydZit8+Nyb9lVn4sGUIRZgwsW
miEFMl9ErnS6wKhGkwpCjPdNY8hA76aG1x6xnm3DD+YsR0smwNanv6Ds8MLtuBEEH0+YXpg1EU2p
UxeKJqLpge/jMgnPj++rWENro5J116D8Pxw7j1roajPI0c0VL1uC3y0JJ7lCuhkc57MmOuXuBvVi
9vnw7DMvIYincXsJT2bYbTzA41+yU5vD5vcmz5F8s36r/tXxEXSm4UhO/mkTKpjuFevEcSH1DMGW
Gjz8FFoVqU7kPKiEWpNK9DwMsdd77X7jELYn+XjGIblYcZq9mDhe0+UGgfycEk/Io6sBtnVp9vK2
j50pcGuHSWFA7zRRQs/AuVHCdMaa1xbLnuh4+X9nIvvdV01Jt78FhPATANoLnbtjrGGaMDwLMxBO
TlmWRNAe8CFkAgXBo0+D9uMA1FPu+wPxEordBlN9vi3AWVngueAPsjdGDrg8jH34XAAjml9w84PP
h91T/ldpGgTBlV7b/MdgY0CKoZc7CJY1FNmpSYsfd9c/1Kcz4sqHSrOL9M0dZGhCLxAsbwFxBiDE
jBCOiByGQw6dni+YHPwPvhk4MU0Sh7Xuu/6YgxU4gU8gqesE8B05ByKXf5m2skTRZVI6Q3y7ay86
snJZ5d4fFxDTb25R/RMr7H+ato+8JgwwDFs5HaHGkHcd8GssJtVlnewDIjAvsASu2gJ35/I0glcl
SZQAWzS5aXxHYG694EeZGBEzr8VrdnUAvEblYZzWoRaDNu1Y1VVxawvMNy7ggyNb4rvD0LxqXmaj
2q8QAGoLgvryRKl2Ev1WhacTry69QqAZslAU6WZl5zz4P3jApBtwTLcfYY0bd8HkX+taqLXFE2Pk
ANkHO3km5rpFofb7fOvGTLuDbYDD9p5W0RvqRus0MA3yENIsmkPe2QlFuRYlsZ2YxVsLlJjtTOQa
LD00fpNtBOePV2IkbdZsJ3l3La03/ok7n2Go5xkXHnhgdDhanCmcITt5UpEDicpZERmMkKDzUdyM
nGl+GI5PIT5RUhC7wjY1iqxL264Xj7pRFln7QmT5gEOkbs6PMP+i2xNf8q4xTktrfSTjuEqd6bIZ
d2Gg63HKgPx5nght1WqqqH4ymJ6LQHrjmFErv4ZyD0iAUAms4QfKJogmgCAr838n5W1TjuhyStUm
SiGmUOaidfecU8PIDgDohLlYHmfALmmoJlf6AM1iJ/8p3CCGtTu6Ap5y5UCe7mYeBP17Z01g+4HJ
h3f+DNA+O/x5bt15EkjVf2nj2IoWjUhOQMUIu6Tas2xmhZgr//dB28XexFm8uqtMPxfmQHIGqQ1+
DoZooRklIIr+jSe8g3+Pw+iokZk/4a86QYsFijae24tv5JdpaszbMpSUzMbodA5UmEaI5Ux2dX+T
UyMC9YU/gn6cXuy1OOKCRkxEhVP6xZGw1ytItTmGvl7sYB7LieLD760D5FfWwZrTFShyHWYjSRJL
vufDcmdWQNdKtZh3IwUOw5sSqfeZbEhWOIADhWE5Dd78IDiTKZ/JHHahfM38gWy53M7KUjWRYSQO
0JiCpStMWFDx3b3HWk4YPcyGDGfdTb4sILuuIEAbiiMuw7acj9BvUuS0prGG+zZR3XgNKoNWGd7V
iZv66HHJ+zkG7qGYCm2R9O+kF5DWDMw2QoavAHZ9QyyTbZgU9kyBN0gYyuItdmfHnvGlZUD0BGiA
oA/lOetGkrxPoq29CFxBszvdLqlDqbJkAaXJ9tXUbMTI7IloU08LRGkT/Ddbnem1qI+2WS/4XDt3
iiTBUWH54sp08zMLoRyuIa1KxUh0l36TMevcOAnEm2ki3wUZn6bJgumV+wVsdC9p2WXuU8nfWxmt
Ot5aFtZfhRgCJMmQ51vRdC1ygamRqHMmfzRydrwjKu3C4U+YvNcs7nBrM8//DBnA9tZkDIQyUbWo
VQpU2+2k9XHDYtX54b/sjp4ZIAbci2XH8oG/yrYV4XBaekObsfeFL4e+lklcJyoL9w0jzaz8emYW
n+nMvIrY/m4q28/i0rHLXxhCZuncAPCIqRHcKrcd+yshKmRIlzbb+Fh7u6jifchRaXd81N2qZeuy
fpqzDdjtmfM6CTJs/bZCEBNHhLluN8r2H8M2jxYRa8WNWqazEcpzW3u/uPkPsdHDtk1uCVnLBsZz
xotKf3Au3zrZ6Y8C9xrxdKiMHSulrtRUzd+WGtZ4Z2Qb7DifT+SXeL6q6MEo6GjAK87p/JjPmgfb
0EuH29sZ+FrqtLYhEryqOHZrZl08G5FH2Dbtcy3W/iecGgrQZnsiL9rGtjN4xSzpXPqr4Tm09pd/
qeMmX6xwYzGF6q2dfB+XrIg1+ot9X6xZHcWEkPbXAA2bLx/a1Suc4yolQAN4m0VkeFBD8iWg51p7
O73KorZa7GxPVUxIQFgUCPg7zgzUHGuZSlH4rke5LXr7upIZP782NRqMGaJod36XaPkFAfWApdCd
XZfLGPbUxAq0rz80q/Mu5jB6HuQUUvihcJINMA4KIURQ8pv+cFZIvyhFBicdKUn+amkPV1TMJuIp
LFyFzqO5GGJdeRjfu3qspmAaHjVwysUeoZaCAhHa26pqotV0zSEjm02FS13kTQc9wOATG3SJ1xKu
BU5r4p3H1zmxM0GfyMN6scaQBCmojq7qZthJG+GB3IfF019j286BywjfUzFYWD7YWwTLzdzrJKkG
pqJmg7y0tcAVTZRvHPBq61CjZapd5ECKnmoDRomjOe9LgaxtSHNmIpmws3xOGpjpTze1Tkhj8Iic
w8yFqQB6GHDmSuAPAaYcuwE1b0kMq/dplnAXHjavreoHhbnr07+Tkg8daF1lTOojNwMYKtB77mPf
Kni7plekazpIZiqLIc5uGhk4at+hpvejb+uChoqhuTd07nYTZxMuSzFrTKXm3CZbH+hrflsi63ha
wQ7Ois3GlyOmSQccJAxaWaPGI1yWMW/At1RQ12zwwYfBSO0kxN89TSbPRwfl4vpHUpX38nqnwnoC
J9XXoAxO5B/40ABDPMsqtVJFaR6XHSJdPUWSFOsn5DuTg+6Qr0vBwVMYdeXS39eVF5tL7Gkhp/XD
/EbD0iWPBXpfqg757UVm//dHJo6kQXFpRu47NcL/0HsFam/OSnXTioXxTS/f+F/AhgS/RQj3enul
vuwKw9njraLsNojmGPOjsR70w6/h++UkRYGYcO7pAK/9da5fW0UvUv6ifWe7H3QuMfC/a81bA5vQ
CYfS8VVMtLnVjCjqdrw0+mdcpkqEHwUH0ZQh/Lt/nLHbCgPYKv2o4NZNpMCw8CgXKaG+EUKBmBSH
0vVPPWkFRJm82G3yOY/p0113tFnkUy3mRAfq2GuBlYKc/WYBgmwIYiTUQjBW1isZ9Ae76Nc5ZBD9
i8QJ1g4ZIZMrMsF5S/yfbfa18OibP/535EMV4G0/xKwQ1KY1veRLQC2WgYZTDj1wKc6ABKCeKChi
vHcONBCN1WeCGXpyW/a8qaHc5zto7h9rRbgajqlc2MS6GAMyK3xxZ6oV39hqIw0Ic1aRxBQUfuZ/
9i/dgoxdHLxbzJOlamiHfimqR4/a63p375sjDO9FJUDYCuHHPAecdL+DsXuNAbVhlZT6HWskWrym
6IplQI+yBlLnNmkQRYE2U6ZGCDx94XJ8mtPYhyUbY/jMvKZqVeXA1ykzzXucOQRDUX/2BaBTgZ+F
TlpgmEsv6ALWhur7iN+ZgTwSkyEr48vKEuJlciE/J2B/lSyJJYVWfvfxduVj0gzVSC4nikLXMf6c
y6JxouN9zx6vEsYswq7JIEW834tEGs9y+KR+LM1fje3ip6EU8ymOLYGOZCA/A4GzMwzpkxX3s1cF
OCdenAZ7cwbl2Bo7ql6BS4zrG2EnnPWd2wYNU9kRhYpVPoPH1u81S7ud+Qh/MVO9X+JqLWRfOfff
aaKE0FTI+Od1CGclJJIV0UPLv6/PWI/I9Rl118UZilL3L2Y97yyqdNCTucjW6pGJXtrY5uR9U7Fa
pWqUUtNkWqborQwq68N3M+PqOkmB3tlOlRqZqxEZE4FWByMwGIclWw18snVWz8VArxDqH0/jTgqw
tS+ajrWq99SPKhjgpMwb0jybFPRp3qxfEl+0uEVevypwogQ/eY52ksngnJoZsdlPh/A3MxXEIZpI
lUnifoAYen8jhAaMYAXhz8qS2bc3M956iYKrQ8P8DrH9FAWr4UWwWYKYzQQGf62+krzQk7o7A3Gs
qEBRrC7/qjhcAnzixqb56Uwb0QbnUdKe5C1SLOXfLVdDf483trb1uxGDvEYqOusAs1IhRLUM8ppC
6lg6ies1pfbRXl6KAS8Z+GpXbj+m1gIP2SWyyriYteg5KAN84SWNePT9Fqw2AAM6Mi+EPiX/gEZi
uOYjw7ToLw5xw09lfV87lIh4hINXH0trV0Oz/9kQjoBlbTVGUeRHzfRA7+WksHOIaI4v+R1fuY4z
znT2hPsPD7c+NntRS77cYEOaQS7+Zb81/Jm0KPahCoNiSoZLk9/e6aM97B3Zs+Xa90XevkLXTRWH
ogTbQeYm3gKgSuHgJrCLrYpDQZ7jpZ72Iakv4K+FHbHUCUNH1P1IO8/sFyPMr88WwaVWSJdKbUl/
Ka6XO7X6/E/jvA1i9SIaceb7y7spc33g7SwYDx+nU338+KhbJEhLnq7jpeh/P+b/f7kjlXS2bY8W
POmchg1TnlaVuARp8bg44nFJB2sVLGgDWFGKtGzuDreGIInqZjjKpWjJZTdVCt9B0/BtijsXhxKl
hhcIBtVouvn43t/g0K6DK1u243tCFcFDdg+R7fQteJXhr/qbcqQDbGU8QCk/vMi2YfZYisidTHIk
dj3hsj8vzLW7mcZuX6T1zHWqn5lt56pbngyvPww6ttUdfQjc5xFqsgQKw7HqlwaqrORCXTdJ3pE3
f5yVS+OwbEzCcAZYmOS8GNQrWsfra72OKRlUMWrkcINLndLKkgf+EAZGpOJeIfbqAHz70lkmyaYD
VIFtMicq1pd6ycv9lvYsbOY/pDcgyxl85enkenb+47lXJqV8TX+natDTBMvHHvj7ABHzo5k9O++y
/+1kdHOU9Y1WnkYd834yuz74cLe/XxYEM8KR/C5X66m2XPSp9QqEY8nk5/ww1jPqIL8OJ8fjYXll
XZErNT2dCOagLYCy6nWjpd5TR0IhC0jAnq3SNLbsuis6DgBuP3xBWYULtmYGLDqkiAaR5Wdl4r3f
cwo6QzIB0goyK496Z6LSfY8evDgi0iUiyDIXO1t4xurrB3L3U9QQE8E+r/rxO1kY8ojYYjLfsVcK
0BeVtqpUO1oy4PjfCDnnVxTwT2etNNVwehlmCebnEtDVoItNT1TA2zYCi3UlGHTiqHITj0I9LIqi
dwOFvQYeSmoyng3wAlYEyIH3k7hTnkm2Pwv20EQk122NQAncDEYO888RKMj9K0o+JSSQZSr3Gbqo
sYxnRHecuZvLckSQ4ln+sH/X4n3nyxRy00WT9sKjyXYe1Q5ou7RpCFKD1smHv7onDqTXd9vnNACv
Hjz/do/kF8idtYzMZtg7FI7BGmNM+Nlt5VplQJfSNVMpOaMmp4l+O0iImXjAC0aCPBbir0+OPUJ7
MdmOuLIE1cwmysyjriUDbv+MU8eFqyeo4UfbH9d0QtE06GZpe9qQkuc7Xcv94tVjlwEayPqfqZn4
ypk4iYG+mmiSU/UFmRlsaof+8yoWajM4SZsV2w4NaR2Q2uWO//coXa55l4OnvvW0DrRB9nR13Bew
OXcobOR+xF0080Fe2dW4AWOWAmZMoAfPd/C5OPGjcBZHmkbPPImmN+25JMySYnxUhBAurzIKmMKy
k0T1egO7H711DB1dedqMPRAgd98Ifhx5b0s2lQ6zZeE+QUH616iqIuCB/x6mAbBzyp6v0+oxpOe1
ZYE7xKzZN6kQ8zzgTJJ/2BM3Dh5EnNTiI77VN+1wjbdlrP/EdsrsQMlGjKzhoAt67i+iaL/HdCPf
/d5ETOUYfWItdUXhiEMuAz1dNMwhc6Nh3CSYBGNK61M6dJp4dPvLnZhPjyrVszKgBq64n1nToGH+
/714p+eH7BcpYk8w/QH1/SjmLAMm3dOVEN63oyuXnCnAEeA64JUA3C9zhEoCDkdXj6qAqOU4gSoN
+w8C7XdDPO9y8aYlkJuhRSQG2JhdH1kS1vKM128YWvK4B4HXhKAenj1CVMp9pm9On0TQwxLax7m4
gmSl/WoOTZQsPbz7w5Dgr34H2xxy56EcMhRh7MyQjwRc4KMcNZBn4cVz2cwBhuILHkkotucjmZ6n
QgEXDYL+DlDFAz1FGjSitYe1LLoo6LNuLiQ7Sx+tu13LCgqk/92fal0BLZy8q7+AdFzFaWL+QDHk
msnaviLtStTjS70B/rJEmtbtJNpLqDRbZkTmpnn5KghxM/EOTHT1P5dxjNnxwBZhc+uHRYYUwsB2
1o6rvafPivB8vE8g8x4sbUFRatxc52IkeED3W7P2hA0mNMriPIBa3SK8ev+r14T4SaTs3sP6+CP/
Bh9NIR9pstR67AHtag6tBSoUF3KQFXowgU+IETa4NylZWM+xpxAfwWEraWv78OEUkxX4CeK0tefH
EHYm82Rue0oy6+M//KUUWOvY6NzI5Ul21svJcOUHeARiC+dIWo3u1Dy/MiJhuEMLKrEpv8OlSFjD
sgBZWJGWgWirq82BRNnyc62xu6z/0KYAV39El2wtIGFhPKTcLi0oo4heFkzcJLJEJJtBjN+l/o11
Vd00U4fDAKsiUtGN9lwCMT+D6cMS6UMgiLs6bUjK2uD+NOCQTQDchcqA6mEvCUILkzk8IsLMhUdZ
FVX/Gqfrq9lfLNR5S0olQ5QctPPBvG15uGHbe0ktDNKxMO3xIfV6QtF3mUEwG90bWffYDUjnDzow
SJJceJFfFMYpSfixmqYjNiK84G9rH0k8PKp519SHG1QvnpkE1aXwOonZJbyWIfUsob5YaJvZbeT9
YsqLWfsp6XwlTHnQF8/eIRRPs/noLDCrcnTdjX0wrLoodK1sTGrc50eCJlyqultxKjj9x1NVR/pH
2z5q20IAdww7NwoJY4lEXMdV3nLJdTT04uvPxHpP5iMBCxwdbmnyUmIjYKlcU2RwbclSIn1SnGOW
uxZjKbGX5pqMmqZMo4BmwK5vnHwOIbrNOWxnRWGO//Kjy3WW5F1u4WNuIfsKrXSaT0TG2NrmgME0
9n7nHWm2Xysfqka9ltEI9yQGOcQlDHWYdOvknkMYIFksY8428oYr3Rx86TpoUYz2SVM0cIEGAre3
DacsGPKRYAVgqOVEt3y+aSkI6C1KM+m2inBfysu6VS50/dMshUkhYqwnQNSUSeCJyqWaGjJ7DO7u
jqaBJwbdAK3TwOqmfOZA9aLmu+9nxKpbzijFUaq9N2FOj8Dt8/+0tKYd3DDySlontE2x4U9yoirY
Pjh0nVfmq/NExgHCV1ZMdBblMhjwYtwgrE0A1YClHfnqM23SufKgIVleuTzbOsZMDh2xY54F3B7u
ldTXbhgfbmDfIkNHa0FpOTwXMLDfKezuvh9BlBR7mdnZ5EOakH4i0jNALXPkgE6B2mtovkuj81Yt
jW230ziCw9V0p24iFLTi4AMMv7Z6ulxZpcZuXb9ZKJLYFD9ZZcLXip3kxnwRUQubqPkG+UCgtda0
aV+yqHxYZQ4zWSOG5Pmh5GdTA7vRAqP8CmwY77scMoBcOWHQwiBTLSM6wQTBYNeWL0U4vr0lmH/8
SLVJLgVCFqFT2wnQDFyHHhGiTtthD+Koc/7MMEirvFe5gpjRNVv9r5iI5TsuVEy6lGT83IPQsJTB
BGELUALFpOLe83JcWR2iOhrgfAjFZ8hJF+TjSZhEkF8j0unSNHQKHGXUXfJmShmFDk+HR3Qe4BcX
mOWZequjzVjYzgq4ePYNc/XiPgnhmGQed1PIRZ+5Sx1Apv4koMPVRw8cp3oixfyr1TwcZ6rvjAXE
dDMZrhcphZyWpwfN2fBSaCKzPP0X62K2DXtwiLcyL1jC6yw/jNpeC/I9a7bFBs/AfHSIwMjaYXLs
RhhwH1i/HeOkYLtDjF3d6pBbWIYtmvOdrhHA983Z2KNHl3Sqm5RT8EwSxZhQmS5PVhtjpiKYlV1N
evRlmmZX9MHmOzaMz8nlGq7+ZpL2e3/w4yq5xwKsEAEcJr+y2jfOVdy1U26ikGvytWl68dGGCnPH
HPEkziSxE2NA3yev2mG5wIDVXDf5K+Lc/ABWFMOLw8kcRv916kCI3r3yJw78/ViaP/DYsvs7fq2k
bZx6yi+QL9cesl82YOTv5E8pD+QwKioTFkiq87cyFcdDZN/KF5vWpvdoOxMq8C6B0swUjUxmISwL
xI9ZOLe5IlZg/7ilLCZPAqp0Rwc5UrcQaHSD59Mggim7ECRIAS/eNSsCshDxqXMlEXFGjqohCSl8
xkFsRcnNEa/VZ3fBV+AlJLi5zMBsPDOuN4nnZ0rveRrztK9Y/Uza+J3JK7Va//ngaDnO6ew6/cRa
EWwPAgvm9Oi1YGBrj4GuJbVN6n214/xkH3I8ttiokO2h+kI/F5n7gZGo8LUczfG51Gwy3FAE3pYH
MH7fM2+hmOfj7VuyMLmI23ucrWJfLwfSvQ+JCMRiLuf1OtU+JSiVkpJvFukdE3a7UC1422ouF37T
OsCQWvz5d02ysU6WghAM27q7BeLKshIDC/Ucpx1/mH5OTl8HtcAIYjtjQK4LpGZICZn/3sM17vEL
DFdozPaTy29N0Z5a8fTglrzHUauUJzPivwGIWWiCQVY4F2/JCZjRr3AHARQQd8hwYlJ/m18aKfoR
duZ5fBNQDsUSQePo0UICZJlNvuSeEOjokGaa4HUg12a20FFSIHV5ACpXyXiNdZG4Uh6DV40LfvPn
QsPTEe/lXIt0HxovhazKzlcKalxXJM0bgCiUcx8OhoUUVyZ8A710tqXITirU/EPTOcF6RPFmlxUh
cEtUV1/JYVXXDSFGFaW6HEPUrV4LWU2omYm9Hp6MNIBu1/qwIuX6jyJ8u8wsOl2IDksODhRtUjoc
6zTuWh2Lye8GUaRzuN+GhRNtGmpjG27NkC3nIZ3zYo/u2hNXQMEHqZaWlt3OhrLZmpWkFb286Meb
nX58KKsKpyKEO822poG7Gz0tI1wY6NJRhYPu+yc8Ox5aHdm/hpWh8+gxn6Vlm0LPaq9YhaDI2/04
iN4WBRRZW9pO+fbfE4IrI5/lrTcyLvmRqRhb827+U99qv7D7CKwn4dBUfyf/TPUBp1Wgv8ObZAXh
X8U6mhWMOGoZHwv+Gjee90Hpb32reAPb/w5cAnujR+PNoN/kKCzMoStV+aAhEINvn4zVOkEyjvQA
Bq80rIdOGdVx3luM2cd8/fiI8gu4GjAmkeK9Wr8y2M2RRvP2WIG67upNRBCT1oxe0H1HMys01kD/
8TOkMvFWoHSRrqnz0UfjzNLgERcchpnw1oyrr64DTaZWbwSiNLJZzr4z3ZCSfMyVXFfOofAdmOwY
b1sfywqwli6RKeUmNCvRmknW13qo9qPZWkdheT0uBOUEkQDb6Bqw7APlM2SF6/EfzbhtAvM+941B
etTUc9eTpxb+1IR1EJPclK/qNXxH5ARV6SDZqcGEjxnSmeM1j/md2Er1r9JER+R+dug/ztsvqlUG
NZDEKp3AFUPS5GuJFqnzoOWldDA87lO9H+/F/d7nauAJPbUtfW7t1BGV6gse6jFJ472dFaoRxSQV
WRl7xoY1WuKeJtExEjuor+HEgLqCafdogwh+qmr6j+EAw5H259fOYmQOlRetH9H6+RaDCxi6iUQF
nVHCAjI6YtUcT+G22AaI8tEF/d7LMRqxs1m8odJ5o2dOFVc35AJ+mA1wWtZETWMOKEbMcyBLnQFj
xVNuBmmiIE/mSmumQxpnGDhmkTRM0axCWWJnpCdboBM7DRRS2G9lwsR/+yqoYKFlS1s7ueV4fO5z
XQOI2sTN4eFJD97CPFmsyOxV3yJfRJ4Hx52+n8A9re9Nqg85QquB+7rQqmC4ke5w9/Wb9Kc7SlNS
szI/CJQl8ZDPdhzmkZWV/JUopHhG5P1kZP83I0mexOvAO1vTigZ8o+6SoAh0+XT1LIwUJh0ujKY5
pdHOti/E3H7dphdGSudiNCPbLo1f+SsBvVNcIw1f65DgE2XSm4AVvnZXMV6am1TbTuMKvu5j+Pf+
1KzA1RR6mPeIDzoCWmE5FqhTMk0gro+WNAfut7MTdCMYwFXBYs+KZu1GGzWX9x7EMYepxiqvJW3r
3c7Olp/rzGSCSTVMAY5TNJlSen73AY1W29qhfcMEz71nZRHfVam1iutAkkmk5RKzeNhp7z8NzyEJ
Mw3TBibDEQnJh9IUvaUOfvtmF3JTTeP21ntRXP2cKuciZjRaO7S12P6upm9KlTaSS4o7HI80JyKY
vGXP+w6zcqT/Zdg0AVR9gBInfRy7W0eTDsYoMxcAbIIO3SeBZSpbTBzLndXO14/ivzudlr6YEHl3
pCd8k2XYEvlfqpbp0XlgDeo0aP/6pNQe97Cqv7tX9Ia7kJG4SGWA1Wk4aPRUDZNqXIm/2v76oUMg
bLUBYQs4TjUqdLEGt3uVlUSvM2HKmPnN6A0tGhcsyOMM9efCvAoM930SHveyLHXuI6fhvE8jwptG
ccAET7o1M8CprZkMZCGrOCBCwqmIq1Rd0UdFaejEiO815CJyw1RxIJqad9jIX2xJvfJyc3jCSh/a
38MlYq794xaQxY5tylsD928+eEYkPeaAzmOWUAfefYzAUFE5fe8H81vHKONxozPyUfUYI30c8Y03
HgUjhYrsKSrb4/z75Efj5AohVr5iz9Sif4G1+zSksvCS3j+aznArro2PU3CAL85e28GTpstZ+XXv
Ew88I1FIQp5j+frtxsAdUJhwMh2+3jat+LVMUmFlBdL5jfiVpAEySYxC7ySIQ3Qq0zbILQEDju+H
2bA+NNxe63A3XlshhqqiU8gAsxpHQe1WH5vIdJTMKeL9xCYCbMiAqfg5qJzZy+W7bbAK6wEvMn1y
p+5/IzMsJAAmNYQAeJnngrcahodPgSBp/QVqDEhmoAFPboMwKzOXnRm5JKaIa7VwLNXwMunAbP89
XTQo2W3BY2mNbYa94//FcWG/SMSoTWJePFptz52yhyOZzQ51k/OGAIQ7T1Sv290jHs1EwSUjrogH
ok7emoXhewUJndtH/oEz7GCNIT6EQELrKFIV9tqo892l23S25D1GStqdUAglQwRyQ8K0yHUNCier
H3PKrnGyP0SebHCU8ctUImWYZPSGoOJ79jeAJHeLeuPpRBaxz6+ZLDoc6Jq3eBQNsjzuBbF2uolx
zh+gWwf/GzeKdkxpQyfit1t3b3RTMI1GUmM9YlnR+sR1haXwwHcT8parFtww6t6eBFhI0K6FhCK8
dkd8oKgma6ZOMT6ZTASd1Zv0vCikQolJujFCCuzdtloykcK9vV+gKNKjoHdFMNUwkBs/QmR6Cu69
phqP4ewbUMjaQjMMQRFZRfL25PeBngX7mWp77LF3QRRGPX0HiUdGP5mM+ccFkCH2kLjg+4nusOh/
F85clqiduvxTfgh3U7P/MGUQTVql4BhQk2u1H6BEy9+57cQJb8kYY5sqAkIj5d7m5RfV9S/os20e
EBx3RImXVpKj6ZpBJmFDFI8prvfwiICjBRmi0/uT9KNzqCBTFFOAXOEZI+fw9remX6pe93pvgInQ
3BPRrEBgbWQMkuCzusKGwg03VOgY3ZhrjiNDSiKkiTb6SO62O9b9KS8DjySQe6uVI72Fu8xZOY8H
qOqHllSfnBdljsqcLbQrPap05BIuGh2E5PsO73DZ258qJc4dY9Eh7bUWevXB77XfrPGPNdlIRre9
47oy5m4GeEq7KScJ3aZvWPGooGdPkUrkEqMsGzAcMM3xDA6PtanVHW802JOb7z77SiHPM7jvpKe+
RYc4qoM43btRxOn6+snMFy0aC7OY9iX9ybCVtDySuRVMsXTbwHA0PHKlVE0tCxWSTgvM+NYG2O0O
ltXLXBZEgmCjRDoJwAvTJ7W1SgQaPrePN56P69DsaO4kLeHIyRmvJrNetv97eArzYCn+71a9Ihor
5cB+yhbWK4ilt2mQDWZ4cpP2WNTrjcMBjgZUlZz7jBQNH8nzimDlPY+MGYBmynuXH4y5uNJMOb9p
DwODDTwJ++4bs/QCz7PBiPnsQWv+fjD/zhlefGZS8KlAv8wEjd1gbdlOkZr1bhP8eFW14QkbtLlG
FmpJ0dzXd2WNmqhjN60BPU0IqPkFCUgWu3fHvbUc+EoqtSZ5qEpdoSzqrGVrZq8XTzOKI76wwzgU
kWTFFjfxU/I4m4/TUd5aEg2s0r5Z6u/NiRzk/uD8VBW7o4+GhGbpoJj+6AHehh3tO4aADy9fEW1b
huo4K2N8izPpyiuEfc8wqkwq9tOBlbS3S7AF1zGiRmbQhrADltV+LBFVLxIVAFqNwzgPh5oKHVw1
7TneSbNlHwfUPaCpIapx/E+xF1YukkiQZj+xwTOvXePLjQXLkcrY44ssfJgYuDIMjvNii4By+E8k
6xvTj6PxGxLz3Lgl9uOz12PdmhSvRL04wGEk73smRGSG9b/NJbICvfHVgOeDz0kOjOMSjwKNyU7Y
HK5JiP1q1JMxYaDMXUcZHyZ1PY3KOU6diGjmmNlg4K+LO81iIQ/F/XF1yC/Z23WgfQOB1GysONLi
rIRajG1qaOEKK+LAmsDYwx4Hm/y2QRV7bG3QesEceOC275C7bhY5DqtUyicuYepIusAW8Js7SsGu
lwpQTLW1AF9Ha7QXtRSR9ITuvyefg1CeYTyAB4w4X5mDPri8eW59i2Vq51rDwvF4UQPyhoOdpSaO
6CdqqyHoDdeCCoP+cIyN5i1cRTY+NZXEDJW6qtUA4LLRkF8gXQaDDK28S7F0xD65lxk5MODUZhBz
lYT6QreyPbUZoNC35VnGu6eN/Kv/otGV6euLTK7WSmwDgs88AOLXOxIWPUByG5HQQzP5l8Oeemv/
FxPTDvmBw/Bjs5N1r1gO3UsVH2pskC4fSGgsly6M1EuQhvxEQ53k8Z6n7xcf0n2ioOijuRWON+vw
5xFHOmmvie+17y3o77FADAuDHkhstqwuwaowv+RSzelubyQV7flRD+lGHFibKtHS3253euJ5bA2d
WCYFjMoPyQenk7AkO2htg1vRefDXMkeCzLN2dGE0uPKNxTnOkcrtiLbGbbH6Gbma0dcdqNREOotD
uXggKlZXQ0wReshThr2O9FfdOrK+GEONhxygV/PmlOImvGorrcNSS10sR99cCB5TRjzn6rdwOHiN
rwrN4MWWe6AnWgABPjY9tWjybAHIHqaMq7Bno1NYRJArmqwSIRzBAT74B/uwpnW72nDMlXZOEwu2
ayqTuoNqj6lF7dSTBGtx4yQQWjOPAIpVLqSdTfqVrjYPPGvDkvGrnQ7/jFuLJm6GrKgTGvBAQ/Zj
7GMAA5wybSbqBumw8TCVamYAPUdZBmHMUWkh96aOtSKnMCVuYE5J5rjcyFKf239ATTegfvBZbDFj
Ct59JULopyNfS+tTa4sEhDhbKIBA1bvI97mWS0llYs7xU9jAyHP0S+uXzOVKnOHhsnABlgwizCTU
PgIWS8ABoDG3Gqq+HtM7cpS/lmZqsoz2WZ57dBaIIdI7zdBfwGf7gc/pvnCXrgXe0JgaHdyzD25+
NJSwB7x9g1yy/c/Y1qNRb1g0UPatwtMmaNiPAQ4nv0KfBr3p/P2Q+OmN/o6dSjANbaUE6g6tDkJ9
I8uqJD/7ZWdkDPVBJMct8Q8Ho0utB5L6BZxpbE6+lSoQ+j7fdikKjrGgIcLds5tX3P8X+/2uV5ya
DZxAXNHoLszHHB71UyeWcsmWSvezAyesnwfgpFY31DeLctmwHaErm43lfTBIgz7+X+uz9Ize82f2
krzUoFAxejUUbXdhP3ZhSGptvZNNkFlZ9KXSo/37e4VF+RFAszQy5Z9aN7b5OXOEabwPy6v5/lca
j6kjoGbdZ0XRaFKPzEQ30Gg+LWXJqHiWbLn04duTm891aLx8EK2CkehtVJcLbag78YNKaC3FIob8
Cgz6SDWeR0qdL3eu9QXTxmEjMDdhyO3alTs87z+9Nq52rp/u21TYzVLIxFhB4LtD8R3T6+gwmnWq
RlZGao9R3//IqxoEFvz6YO/OvtwwSDalLw1eVNVGflPYhBcWskmAC0Efd3ijZtBr2B1M4PlHHHPc
tDLLNlvxusfa5sWjfMAddtVcuTk4zg3JXhutEa/bGSLtqtS0zCF7l85x+Xqjj/vU0uQ9w/Fn39mo
gwg0EtUqfk58Eu3hewFT91alEx/dJORbj4A0Mz2/49m7gx3Pri0dKOP+YLfGhHyp678dMUDtGKNo
jm9yT9259YZT+BQwX5P3hjrq86ZZ4bausisBJTshzF5PcwivxjzuEJnjqnP0NAT0cxjC8O0UZQp4
6xGkDFh1IPN2X7CSM4ZWg2hjnvgTzt4JsY93TDCdSC9sMn1BnQi8m5BmfmVGDK0tnc6U/FBi1iic
tY98rbVOlWPLORYONhXR5VCHmf0/4tq+mbZG+8WVvt41pCGKEI4QWuSdutqYzMgj8kgw+2TqtMYh
/dpZhv82ef9N4Hy6PltzUaV96tLVK+JC0s8O3njVE+7IvZHXQ7yYPCu71gFfrKij7hWf/eOyOjaZ
vEIopMb17rRsu09joXeb+xu4yRQlRQhLKwGv+1NNJyn8ivpo7TMOlpCGrADtiGbpIfyiFYKVos3z
oOuqNn76xrd/zb3/J7OMgKVsdfoev9nUyyXMp4nYPUrRT/CuXssG52UzW4aw7jXk6giYD6MNgg7o
ki50r9aXr/hyucUw0/nQxo5t21kaarQwYHwYfwDtH5koiOtjntjPfseaqF0ARDXgChEgXDjpHCoF
sX0M58izIOwsQCTY1YOGhTaONTEprgSsQasjlvUdFP/lWiqgqQiwZ+5cYntmdHj2sjkpBf/sIqwV
LNlZUz3C4TzdksaPJrgpGQEmM/kGu1on79vYfccdFA0HVNQfUoKBWehZDRIFKslI7BAi2x71ZL+o
tffem6iM9P8JWvfyHgDcnqprwmIEHh3Zt/mJQp7PsV/V3I3VYO4Zl6A9N8pahPWg/JW9uqJzWLoW
zJmkZ5qkaN87dvc3sZgDCIBVEaA+owBMIoBMwDQl3UWyCknDogpsdhj82UvcWZfiSbWkqDKpDYk1
eRBNFlpItfuyjCDVhA+mlxSxqgf0YTPu86TmxrFULXXx4+x1psjHtcvC4MaxE0UCagom68a/bSuC
j7ukG8/Tej1lFAhROpGLW4gecp3SWy+56oFRSO2MiP2k9vKKMme/RC2XwgGx6u5AZ2bxCphNhyuW
vbTcflbIwMuMqlXnC/zv4uom9pkC/G+fxaj+u0nCw+rgI3Bi+opRD/h0x7W9yegWuk5T7rLbEj2l
ZxIZ+WQC2R6DMqJtgJCYDb9F2BGZClaXzXxuwoDztfbLb6TMv6P4km8pBRg9UIoCUutB7vVrVRts
OZj6w2PkBOl95SBtpMemVGlvLpmfB1owZA3242T2L+zwA79t0dSW79u9aXq0ZuKB8lThQms8nnSv
L34CMlTTsM5DwjYQl8XFCq/r8pYuSaWHrgyA7ev+INMULkm4Rtrgm5dUQfyQZTZV+eP0fUgsW5rT
tTw3EyWc4jP7ayj4E4csIkT1XnwxNtkIoYCPm8a61zntTbPgyLLdEetDh0ORkXrh6bgy7aUnvu6O
WHGs22eTh03c7rzM6qIwrk+CETYlFAKVy7cviuYgnR0N4yWQZ7N/3tSaKZ7hNnx6JDDqlOpnVpwI
BHJr9EpIoxyGtIseZXlog3D1Ti6cmfYX8mU6hHO4MbPM76+T3eSqRIStvuT9Og1rCOtGcoBmqh9c
4DBQ7y7iHx4sXaXd3U/Zo5o7SzuV4ir6olCZtDWU8f4p/tZjOVDL86YWUCVCVseJjbsseCJe++P0
6laMgGe5oqc4jpAM3Fp/Z4uOg8fUY0ntEIXI8SxidYm3ojGCDckZ0PzMLe4XB4WuyfRkJGe1EiLW
WkGC8tGmqZnVcwPjY4Y9rk7f1W5KFYHkq+cvLJZqEQ2cxE+sYDOxgfY/dTf02Lpk77qW2WDBBpLW
XsgNbeKkEqh0x+x2BqaAfPNcZjTqh1gaChbuL/YYz2keecImIUbHDG/zNOm7d32Hsio1ms8xmS3j
XuYti5ZVeFq5ko5A7w1FRMB2PGFJpcCmO/On0SBXOauQPwlCRs+Sn6hRhT/c8xHhzCpogNBLhRH7
6TbS6MGRLDbQ6nKnPHXQdVkR6KA9faA28oI1sQpLlmUvjDU/m2BBw7aB/gzVjPBeFNBnqfsbA+Gk
AVM/Lcd44SQ+sPYkhtNbwjQoluIpbcng2aGjRUFQHP1fMWFFRDQD4hREX9gUI1r6g6HjWI94dA/g
VS8IdrQBUmIyzK6pFZedMipxliPpjJIR3H0X7+/8ziwRWOL79k+3dshR6C8v0Ablih0Uker17PDW
s3Rbm/U+pikwaFi5LtotFWoh7x6s0CzV4RfTEeXhL9YU5qaSWdtkmfTI6t3HuiWoc976dkn23qT2
kKwi9L2+01dlTGRhwebPPQQjJcP8TKGUtJgMqECg9OuGoXGBxl7TPEFkh1TeBKi4K6Gvjx9cLfmT
HNAEG5TE3EjRwNiDBfAwAYE4EXi1T3s25mgM4z7CPZOOx6fVNvoKTowRrkaI9k2Z0+9tT4Ywiram
t7dj9hUrrKp7sMNOz0Z9ObAdUv2UQPmaS6xlu0JUkurISxIAJS590MSUyvBHb1OOugyZVG3RUHbk
z+Ub5x5yrodlnZGyeEZ1JCOO7owr53rtEg+4tnl5ffVNq4mjDBi+JjVuFWK+njyK3j2Dbrk4KYV1
GMn6WCxubLPDYHPRsSGdhsOcp8s1mcsJhyANt1xIiDpVqXy4O7lZBA4FDNZuBf0FQkT1xsOpJr9Q
3fyhjdgKuj7CoKfVvYxegohO1NGU8HzjpX1rXwdQgWu2he+KaQyFXqE/gmCMRUVUhMzodbSdvgwM
dTcSb4fNlf4QGX21BwN6Daz09dREwXw2aTl0Ekbn9z3EwdswQF0Bh4zApMCoSsLRpzwvT9Iy/PHB
kWcukPzrCXn8oE0Y2pd61VmBNJ81kU8+fGVxOA4wP8Fx4gZKd40HkHUfKNnVjlmtciZzD370WqfS
OdGDqhoJ2XR4qNpucwTl1l/2Q1ZnVlI8Vh8Y6SfmVHdKAtFPd1dFSnQUPHbkovEJfDHTZkyA1UhS
SbAGj/ua5RLR3s94lh9WM5ZZVuaKBPol1mbcnZFhnRX+Y295OYVacJLjqMyG4Zp73lXD5IzKo9ew
9wDlKiLcNOuDV0sw8HBWi99DYu2JeEn2Ie5HFB/sw4jHxS++fyOjNGQaZKgCrCvdOYOiOkzlSP6F
9PWJafuhmd2VKfBVaFUY4689Ilj0xbRa+EBl7YwX6752zoGphJYecELjSHXTNp0kIiD+R6iUEKtm
DH1gEosSEEbz2dksc9vxs+Ge0kbxfkSbaBtdwrA9G23ZUJOnfHuFX77CjTvK39BswNru9jfR92gr
tyTk9jWfQ2vmiLd0deb7iQ7wIZZPz8jK5VVP/YQWwvy8iLxYBYbHITcAyxJs61IYNk0KrRTs4qrd
TuU3Bl7jRpI/G7lGbqaMnw1z+wBKBxKLdhOTsGCn6+RGcy5FVibkR6BfWEPzOrC7+pVIa/YC/Akj
bxTnw40/q115kPxlx8an9CJf/1dG1Be8IlxT6mU3n5gI+1xVOcckUsFzGj/GhmLRsQ6OpoA/1XbM
hN5hGXO0/7i2Zh0JF5Ev6pkmOvrdYCY7L9yQTzv6TwKO9HUF0DSqFrpd+C1W72LxB42tW19mY9ZI
0IoopghMLxlkdwq6odoOOExBChE3T2lGDDz5JdGpEuPH4ma04tlc+67kxQvuQJpYZAJx8dDD/BJW
xsV41baQbnUxyoCqUsgFzuLa5lItvzgFMvRAVt7Rpq0i3N/JUFZZh8RnPJU6KQqLzgfE/FS6CsHK
wn/lxWUXxjNMqH77urfjr+i6jvh9tUPQHBx4HuTl/sh55X21xtqRtpyQlPxF+RJG18CuXF9OYPjr
5643yHhHgrXDDxr5vaasCGOVFFcHywZ9jXck/FVpJSXe3P71GDlR1jf9djFzlGGwktlMW0aCuylp
92AlDdhrTTwuAfOrOJbM2i39H07mzobm3RfDigQJh8T2zI/PxOtdzjeOra8xTpRtr2UjjUdBxQJ1
rKauw4tK66Qx+kFINlKNsgsnC1q65lbXX9Q6BahHK3ttFKPmgzsqCo8hg5aNq7VdmFgl/uwjw1Pm
H0Tu3LgsXwFEHIcyoalBAYpw6120X5zoylZq6xMEkiXFIKUpkR2YixVIJm6kExTxZf7Cgo+JPyFu
h/8Pa5WJCGac/T8yGRvDSnVQuajEq2zNvvInQjfe+U+O/gbI7IsqDoCzCcyNoCEoqYl/xREtVIJa
R//47QNSdG0WVG95BGGbPDZMuQXxS/coqaKxVUWj3on/q6W6JWAnJLWDoZFeodNvc8DgBBoqszud
2fPVbAxRjkR2xHOwMoSvMBcQETWV4jofpLi3x0zSHYI9O1DcVxPNlfFTsnvTgyhijjlXAsgx2hGN
EK29TwMKTHJC+n3/lu/lxO1kn+E24DgUHZlPDQ5YWK/qObVTJ1Cp+wN/yJm4V78FkBR8RR/7zA25
iYGYEOwvG4/Qt/WQ+kHiPT3xLtnzw0L3eZoLhdhKVpnp1bQNYLlugxGw0+qn6yyPr6ssBfco6CUB
7sfDEPjTBmlp9jd6oW4h1XbXNQGF5MfIhw+Ojh1F9cbBSIjk08EUmDpE5XMviKBjej09Ge/lXTI4
qkaozyWoAnvL6T09PPMoUebBjy9l2u3kURPRN9qi/+ITfhe/EgVh0qjoOFh3ytOizd4iC4V6I9S5
dUHMwhvx6DSnV+xKivgq2cLYOKDioG3TpaAiHZQCv0rtqzUKGhcfYEfqfBf8pgZNzWdSsvMOx7Hl
8ocpqR9w/QYHTd9hYwuIHIphopm71cyWvs/4zm3uWCPVVG9EPOnW3kM+tvmina0a0aNJKCXvojDI
Ot5Vsb5PguFzWZsm9G5LB5IPhUcY8pD6CPiHr+rEHXN1nrgW0U+3DjC53DIMO6+OTUeggke/jftq
W4rmdWTZHsdHb+cRpv8zyxDX1iCtHIci8SC2T3rJWH7yFvxnT3wzZKANeTCfMkzQ8RrIZfax3Y1k
WtmjAHOqHSaddKB+MWBX7v2P6ORykcz890CYtVNb9ysd6XE0ETylNURAB0XqZuX3AAU40+/ibcBo
FsKmWWkg+AGK+4rhXpxKLAZefJIwFNnoEL0nSchIBKItiXv/QxEY5g02XTQuc3NOZXOQP8JPjVg9
XjBXG8LuuaoRkvrlA3eGNTSCZKE6s+Vs+f4jlMjzE6CvPyhCr28PskX1nbPrfwmlJO0JsI2CZq6P
oxyNo1J33qDS1jd37oxPwF4LyijpvxS1XRe+p/wwj3gLVwZVKYDI1KUEPUmCw9N+fJ/nUm02s+Ek
LvA2AsYhkDdchrKHauUjL0xzIcv/U6yU3/+cSq9bWg/xNB7VQJDDeCxuX2Xzqu9C8sJtKZO0wFkm
UGtOjKuLVzXXJrnSdyTAQ9kUgqhXDHU8DxkVIs9XVS5EU+l734QKI/XKOsaayvbkO4ftBcOvZBgK
sgo4WMul2J39C6r1phMLYWpWwcvKzpZpC0OhdSyRzUgB+aMhNMTcxxs/R3Q/hsJ4d7LsT2p4DoYg
fdFtChNAJTjL0nDRgmVf/uVJbxMQxXiw8s6qmlxHcWUpZvnQsZdE/zlW0zyfrsI6Ff659BPe6btX
IorQ4qRDpLCyp58KOBl48f/4NNjRsTsTvuJ+3+GjOjxe+0IA7Llwt8I4nlHzjRou/nbD5/s5FBPY
0L939o9FGVYocjN/iIEf4X9jgwcmHLU0vf/esVF+TmecmXLNS3aF9qh6l5rKuSFjIuf8T0IUAYbu
y4dySPCOVvOQaLZ0ef62I36qW1H9CSIiiR8uM3Qm7Zawrt1akMbSP/ryVF26VpsVy33cmeQ3Fh2r
rrndvpr82kCnb5ApmPitPlR7cfyjke27SgZuEUfAH1ReAJ/7SJ5VK3HNuSBOsIb1jIGoI2qnocOF
InNYH+Cevh9pSq2TpAeP1e+ZzMxiJZ8KRjb9hBzroyx1Z2H4wN6mo3AVtemyArNcSuoRvmbEwggq
GJYNbHh8epQJ0AtNFfg2EuflyTRKcamn3V0sn1te8uoBTiGGmDO+4kDjyiA4kmXeXLbPzYqV6K07
Os4BJfz3cnap/5hbIM+r4ZjOudCOqRE0WnNe/pIlbyRC+whxU7mTeWSm/l2BYMwmZioy5lypArKf
V8iA5guNHkuNo8Mn9iwjsgk7XBUJ8w6brRexdt6YbDOs89Ybjgs5wZexn/XBxwkA1BM0QAkharOt
tScO3YdfEAxz0F0DLPjnzwuVO03/J46oUZTIBfV1VhZF6ULgijglj96m6sC8sj2MTczohoyeQyN0
14+vCO13mMQ/YBj+TxY+ze0/iow6UC02tX+5fMJHIQ0jsc2jLibHDxzIXUmDCs57CCYhpH4wNewp
MR12sQjFDkPr9L+1xzuV2Xmbm2miZ0mDuzGhXQAu5ognKLOmMswp8115XwiggT2YiKGVmmzyHO60
XW6Iz1sk2tNSOS0yiG3k6SFsF/tn8mBnzuXj4EDuS8Eq+TpiSq5QURbYPjiFze3OcGyMQZc2LhFI
PeKMOkYA6o9okzdumpMvGdFvxyZPkZ+A9ZLQGhbaOaGvsuCH73l8OHGTLNr+ql2kKe22gLoQcKKd
BHeQd/YxJjjwqEqKZRh7aibsL7PzKbS6YXbddSNwLycE9qQCzkfljGGHVNx6LreK6+81IuAfwnrE
ZfEveeWvydXbqCSSwDs1NJGWQLWVXtBHQhBlZJqo7mnlAbLRXnjG0H0XZ9BA9hAzfykrd3FMPgL4
RG4JD/7Dd6bgAqxSfJ7PJfHb8ltrgr1yPBGiRCaSnnzD57RWZ3bYMb0ilooDLr0jzi57v8FqsVte
fbqe2a6JznbmaoiDztZlF0PTizqFhVFwrg9xn10NNsYv9+91HH1FOoZ4wT8zXtXSY5I7LMBpkiBE
bilOrsUQUZ/p2f8fKhiMv56VGRDoxh8prFkZkpVL5AjfwEDnqCusunh8HJBz2s3H0GkTY+aZ2Frb
nqxnx0JzkTZIlTWggrhgYoXrb0ZxEYlCRsF1SW0FBrgd1Rlou+/2RxasF4LxKPD/W3HSci5pXwPI
4j1UcmNcuUfG8NMfGXbttekiQ1nNK7ljLwj5+vgoiTKTQqiSK+NL0UiwrOe+YkB544cx0oq44lrh
K3FfoAnRzGq9AOUrONrLOMrlu4XmO4Qy7TTR4WH87QyeX4guaPjPI1wUDzbYYCQg4u/5qhIH212d
b4/vtVSPwndZqli1TAHVhAAsRefTUFoLall6Z8NSN6RDsj7RoH0CQ13oy9OzsmLCVX4Mt6E1y+4+
s44Y7IPCoVz82YgD0s5XFFrNRTrGCnWF2/OeVSy2mBpbr6bJ/7ZBR96Mb141m7IM6Bv8i7Qc1qfr
9hzZq64IByiubdaphHGLddr3HZCw3ikftu5hPnGpjSFvsWRR+6NhzdTb3uyS3/XJOhgP+fOXzF9v
9PIRPMF6G111N2nzaEIpdeztL24jlwwBKDGmiewnF4PPYX36v3UIuRAJblWHXHmCm1zjPRIx8HQp
xmDQwEq2x+jrP+3CJSeg+jGHcMhXjl2mVVK6jJoimqsJa59WFwf2JD2HjAgA1TlcNXkqcEaXeRwo
HIv5OgAiaTkDyEBTWdy2PspR1g+B5Yb3eRSbBBgQuH5bluVocR8Wccm4BrNSEClppE2YSqBORGuL
h+zWI+bGl7VZx4t3ro9JmvarAM61Vwk86/o8zTPxps9RciFTe6fPiYRMCNBkvNeNoJDuuEMUfQkF
6U5yTDaBGUr7bNN6+lJ5XSc8hndsngHdChLfQONYbTG2jIwDiz4B0YWBPulWKXziT2W5DFXHwtO7
Hp4nUgf5eIyBFSIrrsaLimF9ucdY6oMGyB/soW8EMfFlm4CtxWOx62bX9NWM8gASozb2GWq1z34m
FCxsjo5rHUW0wAFsUzFinvLLE6h2VfG/1SLWzkYxA3KMAP8C6oiZs0nGc7hSph8SMr8qKe0w3plU
TvbiNhWoKVEEKvQXzV+u+VRbYlG16ifqYUJg455Bx88rnus2Y6zRsw98568JDhNtOUubKV7aplNM
GTjubUukidi31me+XY0Lw4ST5jHOM8RdQgZe9c7VE2S5orQNEV7/v4gzYQxh7fciwofmfZElz/Rk
Quethy+SEd3sNIdozTpTosm6O5cp3VfA2ZYIB8m37UvZIhbbF02W0E3+ZBZZjGeHlIhhuC23qKJs
nkwhYXmucEHLiitT/zOdMA5ZlflR8Vu6vym4sZGEQFSYZKJTF09Qg0c2AluBWH0JdKWM7eZND58+
l6SUQvO7XEjKz4rVxcId24gEIeMVH+zItE9Kf0dzQ3shPJnaRZK38uYJ1H/+AtyV1tRSvYNc/74C
rnnpEeTgtUjZUfwKbSBPi1HKtDhLGfBOANvJ6oaIvYFTlz/IU5OzkHFCGlCB6mEdo0dVRriHaWRu
L/6641ztZKWAH/en6R6WNNibY8VoIOPzzEiTEP3CPvF+vM446QTd8A8yMnC+bP6w+QV33SKseMiW
jaSS6hpvZNxlnoixw7Sg7HiuzQsOz8iGHvrmdZ4K8RBnYvgLJenSG2L2MJNIn0Iqk18dPhyVGfAi
L4kmZJeFscBEqP3mkH0COGjDLXfJyH2Zg6qh0QaGU07wdqX0RcYZL5dOKnj/EJACADVXTaiFk/iO
c7DMjx8/CmO+Nf1heegL1rdKTKyYnpRHN9fJdHVRomRujdaXMNwRa/dC5DHTL/zjPyxTYBrUmmhq
9/jkVCNcT9bWcr3fWI26pUta399XiJZsrRtMzDkATb0uyi2cd3i0uF5TOMDuDp+8QjQDjOriXnI2
XdLuxRh6Hve0XKDIYsvEQwKMTsMludk+ur8QWyYUAeA2paEzvaHNE8bHXBt2mu5xlmAQU/dip85q
DEn7bSIOiii0Sxs9e5BWLo/5ZGgt51ajKcctIXzx5H3Aiv9mOhFpqXhe4Avb43Y4zYizGHGM95S8
9//6HwiAYsN87NDrniyIDP3ir/t8N9wBmTK571VcTgpTO1NW7S6cPvTeKKNi2Rb2fwKX/aa+NOE3
srlR3yKeHM8Yjuzw6209ZkoOqgVwh5eNP4afrOSOP+VN6Xq3Pg5P8ZcVl0Lq/J0/ovWNRJ42MbJV
pVMPZrd8xEyeQXKqGSe6+0PzwrLBZMpB+gr/b+TAOayiig6qHBuAf1VKnMTC1G//fv0JT/BPheao
zU8ag3wdiogcfrsemq5i/29vRR7IRw6ayIOyjWE2bBP7qX3TGZzyURA8+rqT35kVdDn3V8CIAT+g
HemzNR+DBghrJg2wgFlMQbD7v/lqY/FlBTnSC0AsR1Q0Ny3u6XnK/KPNDI1seP6EhaBfKhS/r/1Y
k6OZ76YOTjK2EiRlX/KKMBqAV9VDgHpzkuP9HFDvOwK+4oUW3h7aQbPcnTRa/WyYPAJpZeoKO/oZ
lyPL8X/rrQW5Fd6ChNOHh7z71NFS+awFq2g8ktnVuoNUR8tKRk/Gm8wUArHi3dXrcvVsCaa6huHz
2DhuwaZ8e9SuGrYiIaDcfDdwPnzWsFaQ/r9K4S/LFFGZ6Y0ivZQkC/rd6DWgDjFBi2GQEuByMl/p
Evbl/K1h6No5LplNweJ7X528CN9G5DVmXFDxxxYtXJZbWo/cTm+JVpqanN3wH/Y9J6GZ+TU3mQwz
mbX+xcINsM7psXMYH/57zyu8zXFS7+PA8kF/1du4g8sBAwUcAz4XPUWG6m3+Zj4AA3wCxtASGPU/
KMLXbLJmIZz46+iQswg7utZ508si+OW/Qrm3ujpR5hRJBAM681YjJR7hPPFBRHK9CbepHBqHU08B
Zei3SyTgnpCvbXvzN8ekdKSXpHegnKkGJ+hpsp8I0E04N/Ybha+zK4PT3d706eMqobxj9YvLWtcG
Vo9IihdKjZeG9NkNbBMrleojT1+BTE2VrGJyoaq5u6hQ6QBjeqzaCrGpKeAM0JBcAxXE6cMja9LW
NWk7lqZoyI9ya1XNGIDuqR7qsbnROJZNy7bWdWCx4V+0r9aXbxkjE2bcDLvOwC6lZmUeZnUau5vx
yd8gIOgiZNs5Bya7qqasH+DktiHeZxKeQcplrQq2UXEQb2LWKf+YyIDLmOGVN4qE5OUhKy5vDqxk
IrU/ZRu1g7Ve7ziOdjL9QolYkRLY3xKNUjMG+F2/IVDA4yzfuYl5Mc1z3zC5GE5dPajHqcRglfqI
Z4rwtlM7jesgy0WFpp8JhsVg0NfEGsN85uG47OPYYAqkM2Nh7gF2Ay7O4jV2zcg6back07c2e5G8
DfZow3SlMgHcupfXaudDm15EXKc2oSjkIf6n5HgD+CsWq7GwxXeK+q7c8HC3x6n1p7pbiQtg1lwt
0sdaLlqR0TZAyJpmkGmpeBKCtwTBkt6/jrtW0cDc+VSh4HVgyr4PlpHirpsrpabbUXTWH1VEx49u
scyVftfhmttNYSdRnwo5y6LF8324lmm/5GrzmuWf4BtGWbS76lsM2n7uEE/aFopXcsz22iBzP+Rx
lz3G2u541NjfRw70fb8UMwyn+FCeRh0jUTtqpDUcs2lvlMytCll7Yz1acLHAtBl2ir/vLEFertaP
0zz5fyBbUaIkJdR4ubP+uTmCBNAcvWyDhv4VAAXBV5Vy0AhV/nJebjzdfJCskesVQTZ5P9HaeQ27
rUUVQMkdacBdPnxO0rBgO6Fv1HQohlTxDhBdAJbDpVxxj64fegJwC1B+uVr1Qxdo2y47zqMA1NHl
+mJxuxzwXTLqqnO6Y1USbOuRtHjKdzITbzctnbetA+N6ux7z4zAI//EX0F+y8FX38j98OGUAPrVa
IB3xMwEACeYIF6JmhX3N0FOqMB7FSZaH6mVVh7uppM3l5jMlBxigVQr21St/YLDfHYz5U+MQOXyI
90RBhHG6L5iuxdOUw3fUnsd4knwJ2mZCCoS/WCpOWUXDciS8KBFwFDEwoa4eFISw1vL9KrdhOl0n
FLKSKOkbXq+HzrAMImIIlbqrVGuw4j1WpiZ2NzerqxskyPvkwRfj32AL3jZsCFfJscfeIWIvZS/3
b7uXgICsAOzUdcayz54wL79zC3KDFwCE8u/F8NvNiTGbif4UazlmRLGakI3Crit2b+3jVuI1uAQU
vQ1Ft21Srp3pYe1gyfcUrkBiT49JonRSTSKKi2vDhBkUiRFx99PVErrbmK+fBp2zvD4rIKsDWAZG
q/mBf1JXkxmJVrHs6QVAhhmYQ3G3N9+uL0bKnCQJQARZtk8cstjOHOBTqvmWBjqVDRkZeV/dDX4y
eH9chLm3BmTnuOVbx/n0UvYGglt+Xpi/yvJs+AH5uNo/jDJfMpWlwJyYhEtYlSdt+goGxBGMKnHl
HbLsRz3WMFmSstJ9FJ//UE4AMfo034C44P1/knPWUdfcCf6o3zhEMqbQmjw8+o4lqRuxH/cHq9LN
Gx3ANHnZocNLMv00CKn3k9waOBuHqqFT8Io4WWLYHI50++QqdVNYDj4RKRz+3IuLdhFufNgiRpJb
+wQ1Wl//Aw3dMjgGfInHXO4UoyurGxYePSJKOnjfKiha96HXdC4GmG792Xl0rQZVKrHvC7enXXqc
Q3lPXtwZX7NwfICQAFcTZR/zW2JN/PGvw+CPX+6s3UZGDAYdXTjSuGiEdbEX9ywEUYsPPDBnMMew
gUAHoE1s/NoK6lGqkvnfI3L28bpm2142DW0S7t6w56D4GZeZ6azvHA8eFV5iKWuRg/8dZV5ybYgU
V3yfO8jlCcbLfwEVM603aXnmhSQaa062tUDkm2HFscHejFclIw5s/O5WCocuZn1ukstT603bt8jj
0U9Gz4vp0DQY1RsJpBMznAM4ueyIql3+CuXhP2masZNbAK8l8sRsQ5amKeapKBFC4nmfdvxHw04U
tnT0yDvZnqhvidLzJagvUFSLDoo+IN8tXiTc3z5gqcTyPsPQLFlkDA6iqx9td0l9EnbGV5Y32BAI
W3X72ER9CCtILjiWGgjv/+3lkYkhWxCs4cyG4OmTzAAU5BKis9LbC0TD/FvH4tp+InckCbwBFQYD
o8SZ9wArD6qdswR5T3AF+xC9gzUh0+fOK0MZ9sIVmfOuK8LlBYdW465emddh1Ofg4CpDY9ZBHZzF
iUZQM0FhQNjLpuYn7vLtDlCCQ12tX3Vy7OGEOQhcq4Yv48y+rQqkRf1uhyIlwC48SWx8psbu/dSX
EV4KQIh+dGY0y2KU6HB+I7KUiTUCtaB+PAo/gho3hiBo6Ni68e8i6Is4KEUl+QJ0zYUxX7uVIDjH
90g5RLkiIHRRqMGvRAOgGRTvjC6f3vwuRjUm/ag+56JrofsLJMZ2F+hGclVSyXzsyuBvhjTQjLG/
2on+uZ9bHVKAfqdH8IxDqDiiWNBYyymylbkHDOT7l+hewNyO/vzzZ7eRbG5yEgdhR0Xsy9payBKU
B+iuVuf5Eik+YiystRw0uX5FCIkAQkzDD6DRnqb7wcTdXU5wI8/bJaiSAycXXn+CNe/HrBbY0X/i
9EPZwzmoPqreEj9SsUz1xR6CfhGL8DHvcD1kLedLPj9Qw5dNg/rRN3qj9BiFCWtwGz5dqvvtrtmm
qo4cEq5Fsu64EA6yJ07QEBWbxiwvamRnOXRJ8iIp8xnO2wSLRcqExS7sQgwFzpufuTl4Cc+FYRa5
kdAbJf+SHhAaZlwxVhqvgGr47M0KOAbdP0R0jTgqp63tnwc5ne3uq1/HR5gPSFan1EM8KaP5qyRY
hXuwRRlvuaS0ILaIL+a/+QynJ0dcyJTjMInBw4/xTC1CDH/AOIacygqsbPTnhXSS3yjAUyG+wawH
JshpC/R9xQgRQ52reUVCQdIxgsgEH0wS2eCaUrFZsTvtbZjMSWcZV21vjz6RYZcEOe9hAW70/K6C
oiX/P4bcpYrt8AOfLifqGP2FsKTWxrBkrNSTOvioktj7LevHCd7nLKGOtss0nNZv7/0ICW5ygFYu
AXw0blum1bfIG9jn7OmXEoSMssOGiN4ay66EOI4f6wSowXabnKgPNdZP3QBUx2JlJUYDJWHx60Ey
8zAHA8Db9B3RiH84N3ZrU0JRsj0p2K+ShDDFKWnUbz9OIPKotBUNONPcpOuN2J3mBowtpxqyZCp0
PAIDKUN8o7Jv6qvhSxMLNsFjZr152KPuxJyo8TAiaMOOi3N5SWmuzAvcBhdq9uXjPm66C3COVFik
2Iu5zrAflAc7hvfb4WyY8l9nWX2jXqHcOyNF+TyTLhqnMax4fjwrRuRKtwkUyTKHv+ov6xmVnldJ
SrkLy7AnQR+Of45O0yJJ+LgzMsug2sfN0xcpzM9BHpknILwtIUX0be8rFVQVX052hmdSTDZC1TlR
kqFzciTGv8QB7dvAphfUfMq0D1vby28RyTlrZaURBglDa+kRIpqVFav0VFat+W15ArN5htE5nnJR
X9xmI/xFhcfDPI3X2ISL0yuODcDMSOQZs5iJZRNXbyjvB0TO8VaGCUzELw10liDyaYW5iIxua8Av
FmyWTU9Fr9joUui/p5OsN3g2VGJPcThiRMlb2agHDecdEpA1b8R4nGCQP2AlemRBNu3B4zMP1PVf
tSenck2ywwilf5YWQRkNjqwcv1B2aP+rYfDuNxFtUm+REJ4GuadHgOWB63P+BpoGE2z8ejAmTD1n
4XeexzG7/hUiIahoZt84GS+Pg05v1GMG9arDtAdvKwDJfq/kTAwYpfbKZmVzEfkjLlZsuBnMa4aj
T+SJreHT3aFnreIFLqGUm70iqxTCLaXSojhKf6HCSnFw+cvrfIKM+K1+4n3NNX1YRf5Q4iShcCRi
8Qk5hkLpYM9IBU3hOTaZZACu3Iq4Wm5c2XcyC8wEX0dpfk9a1lHqfTYlULSWt3IufAQpM5uWnryu
MTMvUb+IcM9nZipz65wMxJHTcJggjpllVFXJQFo13fQKAKMSjzornIt6Da/9UT+zwCyrMoauKLGt
ip3XBUotbIymxswrHQawix7wTp2P86/Hjlc2aczzLbFDwZCB0+rgS1zEpOmboCUPCyFLT20+/FbJ
yHhyn+6ErlH8VMJp8Mgd8mTzycNc3ol0kU4VyewpJqPSHfOwcr5fDIOQhVHwr7Ov73pusUhz5bZN
b2g2KcpnGrZrCyCAXaH7QOzWbiE5jrwAOd9aTW/qRib4fyhMahZ539o2GkpK0eWWjC9KvCBOBmQK
WceiAuzed+dIcunz+tYk5xWP3tR7kz1hoM2MbuQbJV6biE5Hs8KUR5AYe0xrHlX7tbj+gFyx/pDq
X34OchLAD3GgQWwdi9plvdwxNxj9/FQRmHs9FpObpUpnT+hfnihyNj7J/+l7KwpCNcx6BYZSs4Y/
EoK0aU/IQb6ZV9fBD8OZ6o1iBYk4PzZ9FhnWYaTywKKGxq6LS99SV0oYHdXCepe/A9kc8lehHChI
z5YPt7lmO4JwvWqiWSZicUFk5aQUTU8fv41ORGpT+5/Dem2Ijft+b1sXMXQbPnYlMY2g/Qn11baG
FY/xgHRgfdZLevsJqYGV5G/aXeRg/+sjvMFow9O/xN6lVEgIe5YGLNfUhQEH+y6h99GdWqknm4I0
cNwwjxHPF67rK4gfg0ipd6JL2QlcQu46kIlx6+QkPTfbQXP+acNouKlXTB4oadJtJDPrtohDM9bn
qGEUy6xHKFUlk9EHMmPbYBSRpv9dPwb6GVLoilWY9XeQT2HkxrX68a9lX5LOkTDn6Bc0sAj/BqTy
uowrHqpoO3iz6ideoAAycgPXpuroVWg5o1saxWud1/SKqCbRx308/xk4WqM1n8FUer0uikM1d3Hh
URbf5tshUAkuSghD1bA9zTgKbNqEt/S0G5WnkGWRYvUAh6N+kK6f+R4dZzFwqFny7wJTqkxs3YOh
36f2xOJLOlqqeLgXamhCCqvZTAVK4cfScBBHeFTTz9+xq8qjwBXYUhBMxD6YehkSwEvw/4Oyx8j9
GJO0qDa01CQQ+pU1hLvt1swc5lzULRVIg8xffKs4CUsdF7PnHptOENFSyPhE48Oli/WMxSSnnPjB
/jDvnn4XOLfjC3p3BbrLzcsKyO5BERK3qB+iPiPwfJDlDDEdB7njVmnuR0HaiRPVduQEGRPwrnNX
651FKHfEpFnM3fggTxDrDCULftGG+hfRLRQR2Mig+JBAxh3by4QKS3BANZXRyJUWqFGA5nKVZ9bn
TjjYK1/m8MUvja5iSBq5h7fsQozzMCRyj8f/fjsH8Jeb9EitmKJe4KM4vAWsxAzpDX8omJH1eGp3
6uTTRvrQcXuYG3w2f+PrYlBJwp9X+AHU94YeqqXgH/kWh1G4U4UD03X1Yp2bK6/R6YvOHVlANvtB
dSenhphQBKist2qnU2wVv5JsCl+V7KVwvu5InNx2ADMF6zLZ5fV6Vp0nGYvNK+zDRLGUkEEu+BGF
H8XdQ2eEBhwFWzcEb8Hmiw9VBqiDsWCcZthw/HoBhWjzuWAawMAIpxx2g0VXwo3S1XQaR/y4zt1E
zaUdws3cU8HEyq+oqN6arY3Zy2VYALsxvzwHBf4M2JftGaTMl35UM4FTbhhCwnZSS2NKxLeb3IF4
Ye04Hfacuo+FoBwE9RS/EARAjZpWEqDkB6PMzO30vp6899Y2DsrP4F/KbwgKqCnkoV+oIjdp+7X9
F981waXyCw+0VtfFoZ36Su6cgxsCmPfrBSMCrXwIN/FIp+FUGhwLOkbQco9XlK4mKNLg3DsS/iv+
hkTW+7uwxqpaFwiJLBUs7cZSQjoINuDGoPtJepx5XRW8GH9LXtJYpZQovBQCYKx6H+YXGgzqL//q
DJS40lpWKt641VG01iA8JygWAeKkVZdL55ToAp+gI5hmkoyucwRuhABfyHmnWZjFrVwhu1iJCiCW
BJ0HZJHqsm0VGVY1wJt54qp7gj3GJRHNFglx2SqkylHVyw1e2kwXFUnwajH2YucxCe4Wpw2iLBb6
wOfSVoNF8jJg6/S9oJ6XlkuR3qWEYUjOpAKFGztHKdMn77dvYyoo/kHUZXhD7qu9VVwFskMr3x7o
NaAShu5Owi4VQ97IzxDSES03UqP0Tnmym/Jklq/ubg7OuT4W553G+GNjEnD0X0vfks+q4BWVv1hV
WqbDTi7xbavxf8jGskBSK1E3HWrqHkN1pgUaumIEQMTa2SPr4OO1u/4mRfg6Y5PI3wv/D3fVMBm2
tdFK7CQsDo7XdFCREUWNu3gHiC0pBU/C2sPBUzBtbeNJ8HCnTz7eIsKTiBOzSzfqYAtNLCl/nnTO
j2Ocfu5cykXlsHBMoGDu8v0zY8svnO2uhI/bbOdYFDKsnRaZf3i3sEBHwt1ZByKVLjpCQ5esQcaa
DYk/Jt/ETGu8C04odhMYmIGcEnmK6BB0on9rdl5m3Ux/yZ13Xc7RSlzit41IKm4jKEddrsgFx/sQ
QbseQcG134HLr+0rIjLRDOIFM8j1H7XlA2SnGPeeDC7uFvkK5DHOeJxjKqtq7r92oYsljzI2QN3T
cjbJXe42on6uDDr2xJ73hUBz2eoVuCbjUjcGUzE/8c0qzKw5aYceMPc68snyVrUtKmfETiAGbB92
ECH4AqMHrwc/s8RwtpmMVxpZ2OxTY1xF9q1B7AQZwvrWFY/Q99aW+fhEJAKkoQkNfiB+nyPQza9f
rP1nMbxDrvCoLJiT2+o7S8BkuRly0qPub/l23feS0B/v/bVQPs9gtMgLDf8Zs57FX8057L0FSQ/j
Wuy2+uowzuwFLmIw2qvReOTSjZ36qFA40hjUgYiRclSVVIR4FXEhTo5ptWCBF6fS0KVkNxBcRSas
+47NZIrtrzs3enIoqpt8OfgrEiXOPcIJuuVvjK9x7bPSXn0CpluAPxf5bd2AqneI+9ZShV6JWlLJ
HvOqMz7xWtloDVFiPWrmhgAZ16ssOZ3MoftSYVGwnor4LPphvLFBTH6OxZOVjcW+9WAKmUycmBo1
tpvVAeXO3nucC37Cf1E0Fl3IekE27Z3X86zp7urT5iATHsOX+PLl3hwEpy6ssp14pWcm4ZsOH6pY
oudAm+iqLs6caethLOQFdXGiBsAhQQevhWr0vHOmDNReSVu7PZY9xEz7d4eG9xdPHAo1SStEqGeN
a/Cl3NYUsfeiIxcs4omKHuJFf+itWI3u9Ryww/jF+2FwauXbv53iveEpuq3Mj9lMYIeOjk3anBVB
j0IQZB4jwDKdgO/aMgxI7eqJOFGpTbDPxBQSzsl3QE59TTSfkdRc5atOVXbWiJp1V/tMMUovQuAh
5VbdNBjgzT4ulTRz3G1QB+p9gi5wfW0/855rxIhAWdJJcH8tFrb+vh7LewtHfuy1UW8N1q4d1qad
NnCKrEt1r8a6ZLSTctTCx2Tapo7cusKYiEHC9egPQ8OV7Kk5vGA0KV9Xemh084fdMA/TaavXavm/
QU+HFF5reBM3F8I4Henwggke72pYAzpVZtTZAh8KwUew8U8uv0tKTM+qIT/kAq2F+VTg0rKzS5Ib
6wxwy0in4kqpyOP4Ak/rBe7wumPdgln2AJ65O85MJb6LZiYHbtXhpgz0DCKShZKoKfMpz7KgH+G5
W87SblVW6jl7m+WrVftq+RW5lHvb9ewUJ0EOVF6NtpO+Tf6yrobnwmiP6pe7gd4UVzrdbml5ublw
pA2mO8C9xbF1EjuZnGyShdL0q1R+AzeIaI2pNnvnTSfd8aNWFCQVWs+FaBjPcZhFLXws65U6SXHp
n9GdJHgS2yqhjUVRFshbkx9OD4UGn9Q/ow1fWrx9jUNwUFDOyjS69skqZsAfLxHIZya6SYlpfUd0
q0m+DpQsHsQjTabOOauwC6MvE7RahEr1V1371RbA2JU5mhJG0lTqu4Rr3BlpGig02B8d04fnm8ji
EKHV44KHhfgPxxsy1Qc/ppgpzxZdP4PFpSQ5HnONIviOOld8GcX/QVEqI3AqMtHo0uYq7emCOPZK
xcmaenl0WKeUDLulDiONty5zhIZ4Q9BGg8oAQXMGgrKuAvaW8ZDGIPsu5U+He46LsWpblStRPwlv
QITm1NBvHedo3G6xXYNvzQJn2bwlI/ZO0GFkQbA2JJWjiXs6pFw+jkc6UAZvgIuOrWGlkadNGo0s
6xxnvq3Jx39U3WQDROXNBO0gnNZeeh0dOyxmoU3ntMdrByhSsdGKkcVJeVqw8jfTezPF9Yx23kAt
5w/FgvTY4Xqe8DNd4ZO8NURkRsDapJOWl9alovACjw+KyG46HhwI843YmNWFOD55huoTueUhFTXw
vuxW2jq8McgsdCuiLWItc9aqt49Rql71/d+eZIbJ8Tve1RJ5zKgKKio8HD0IlFO/VgPm6c+ZiUcp
wUiC/AXLiLcKvUUKksfGynnmlTNo96D4n10Up05Ru0JS/lz3qLZcV5b60TLvm5b7fzBI6/WOymKe
/UlsDUOssvt+CIHNRL69KU+YZBi2ETli0M5p3E/iy0gd0VNMMrMzQ4dOqo5Ek94EBu3UnQjV9Zqh
1AozG1XN22rsF7WPZWRVAdpetfMhWQlFmoNuumJjB+e/ae44aE5HHcWfwm7WkuqtlzugRSHjAH66
P1Decl9r7vCeFe8kPsuDgFW0DgCO7bycx84iiBRazfTTKwcgxafXetiO7qZtAA9FvKtCSDbi07zK
UjSp3dla/fuQlY59foRT+H/InPVXFsUpbrx41uo71U2kX4+wU5f//UGqB1a+qCskbJpE7GI4v82K
D6dmA5XyBoHcvfX9uG4lAaQZlROEu3YOAlQ8gnCrRqHB3MwNHq97wAmxUOEADb0DsXiJtaXi5JUG
9Ex4pAm4kxQf0yqq3Igw7/9cJL0+ASq9i2EjLSFLzNOnLTqESNw9KJUv42/9d5MQHfwKyKVdd2fn
iESQbjXSjI/hAU3K/9/Dm1+XiHJRTUu0CVFVXBupYMDGmHSNKxYTTxtLAViUumI/qrfi2IuPg2yg
PDIc6VIfIjUvdmMTzhileIZz9Zth0C9TAkVLD/J/f8OGikNGwWcQkVy6vQW+XMVvzi1edkFC5ww6
ZNGrRAMhAseNfJt0IUcKRpNK3ytp/MKDSWNeFQP6wMQ9HnPCRqqgle/4Bo3dc5d5Q7nAs8yOMVEw
olM3Qs8T9x32XWJMRa60+QnQGDbuhUCdMadm8pTMkcfLmdWCL/TsAV4g83dHkL4XIJBXsUmzQhqG
bnd4tBR4klZtsOgpLNePTizwyF33R39hCYcUyH7ufMiMItXODme3c5LxyktjiQaJzcEd2y+Pn5vU
XndqUax3c7ijf8Mxrx7dQS6OsA0aWaNNrE9UdGjqj0TmMsiNP9RKUWCetbT9RR8tKW8wrF3wsN1a
ZwUA2nlccHlHsSlhgY2AQUjTUAgpT4CYs7UP2r7wNxTVyL7Y87iY40B5kRIRbgvOCFn7rkSaNra7
d1X13R4c/erPQWRijE4+lvtBsAjqbZXkqNPdTHDFVdeimu/9YrZGEQXYfVkzbfZtlaOG1VZILk7V
ChFGD1zayjT6LIYWYl65RFJOCZjbfxmr+LLb/wXWIrtxahqSNEj4QZiBreCg8hr1rdk9TtVkv1mW
hitSjm8XDdBSdFhnwCDq0cWWKRv0IBS376aLrYi2k1I3+LoHmpF+hnA3VXRcBgDvMrjr+I5TaEkg
fzNLVvkwpvHedm45yVei3f7Dqo0Va/mrBBNgr0xlexKC4GdiXFbK+Y8xTahp/4qu8sLQPs8OvAvI
ux0g4sBGnRXkC2IP/qGuH/70h63r/Az1rLp7iJ/rdhEtxLs0v/fOL96sIDrPCVCOQYwfw8RqLStd
2VPg9sOqzlDNRnSi3z+RJ4dE1C90g5Bdr6CiE6tyPVy02LlvzSZEGH1tMAABeyZ/LbdnBaMnoJ/2
cp3jlxSQyZAgWgNZ9U7WqJg2QYQkyAR8BArvHWI9YGl34fPGIfgd4fTF98RQ6t3F323slfquTHRp
OqBbTrUHnJ6N9yN7kktoFhJZFW6AEL8CsmE7XVQ91YQ/2mqLphcYU+g01LoOlvBQ/N95s5g/RXCk
VjoIHDrofxg4hFg0US7ckFhRJJ/mBIsRYA4Pkd+YpvG+TXgP1lo3rRivfvAq8jyAkr0QD3bhE7rO
uyDLom7spPQnl6meybs4YnkjwR5Lsoy5WVi/CHCOJJpOrMN6lkiR3r+FK/2MY8+1qINtRsjrJLQd
casRrkMyy4T7IaXHJ67TrF27ix0wAY/MlDdleSnJrTxSPCZMP9M9zy14p4hVamofVsFM1YBHjth5
uOfOoU1tJsMYYcfcx/jrsD3D4QyQJPr36IZKaatEWk5o40Oj1lx0wI9RbHy3bMSc0dQzsGdQxgLu
6k90/x82xENCh/tS9GgqxXRb4wbs1Y8JMzGShnLh/652xLfY3WLHxa2SeQ+G/RGGrrT+ViV/jrK1
IIxbsLR9QX2mqW3jcN9L6fzs+rzc7s94IYVzpKx2QuTeC+1EZw+BBlmW+qAXd0q7qoQUrf3ByAPS
Y6udK9sYeA04TA5ym7ZmiEi5GrTzI2pbcm/V/5UANhsf5ZS4+EKzHUC9OwneIHq8Q1TBKKt/abSs
ZIT/UJvSBli0gHiPrNsSed6jKsoBZ42/wuqMfTOkpyH/n62XOgCSZAzq7xTSZdp6jUJZwmoOvqfx
smiIi3tfrVFyR0BcNZnBfLAbXgSCBphC/elEWAEmWHxrhvJ/IWNBfF2L+ST39kSQdNhwKvViP60l
IoTFCR8z2ECgUBFDvjmOj3ndBRHszkdMewaylDSEptXrFfwhTEJwOTnlz8kJ7PGQyefBIxX2nUwX
IfH60+/USqM9RgZGURZQ24Aexe3Ygo3atcsNX4LnRVFdcZHGVdq+efUoufGeQGGchkMx6IWXwRJP
Pnv17t7BVChDCCWkEIbgZuyclsVO1XtEWDWfwV9UKnkqbJ7F5XnD6zouLhrfmanl6plGrd9A0lJz
y9rkqavIHizAZ59Dmsrif/G9MJddihnU/xRVYtJq1yvH12N6qMWdTq8i0eKqgvyd/Q5Q/y+IORZn
dG/QrJWeGgt9Hekn6WLFqaupDUbIrNEMQbMb66Gdzwiz/SzxYdoSKqQXNcSccDRZSw9OO8QyhROQ
tQheExi6t9hmN+7u3ZaHk9CONgLSLOdfHWdpW6DbEUbCX0xAJCtQTjHb0Q3b5XBdADeAjar1ymaN
2nB5hQRTaKkGMP9IIM9QOu8DsS6d0FYOzUSRBTvlpIp1/rstyb/mEWQNfPA26YoUnaELaMWXDKJE
pDpXy3bmtUzZA3igXG+ayTSq/pD1RdZxVFjx1x+9qGTcOonPLp+5jINxxnLF8i6VPRhsQX0KK7WN
94A5iXLaGNWcgcmGy840PKY9ubzKrtKakLlxyXNeWophJEqE6GyvSbRek2dBF4aBWSDwcaDDzyZ1
4BHxMToJwQy8X9iA7bBHnTEYgUTSenMr0mwQwjLVBwn8EtOkxkc7ab3Ki++UkwESygQZBkkq6TdB
ybteSMWNEnLkex+Haw4BTdjCjAXfhoKWUCf4QvvD8fsU+stnixDgFCHhavGBLjMjEbWEkgNxx28u
kD86XO7Vv0rJwbABgM3LEGXQZskiUYutCspZyN2Te5Y3wIb3jPJCA0WZVdn+Ea/meYoPbW0X2NwI
Lu+x5CLrnM8lg48F/twzGwYCwn0d8yI/E/IwCQwbsNWXV+P8FFQDhaX9auSG8/ovm5YLsGCBAoZO
PGqE69wGcx+7Xq1za4R+YmRzJGQ0QT1JP+BR564pTUxynVwFBuvljX3HLxS1DJFV9dmOjhO2MM1s
LeGq2l4LuN2S78bKRKBj3K+1dvK8ueRKZ77c7wX4RJChgECjbGmakqSfbYN3KHU8RGxU8B5WVJ/6
A9PNUNYuc5/ghghDUAQSDIAjsNiwN3lz9baAKoGrD+L8QenIW3AWg3ajKG7lh3uRbaL/iYOtJMUP
nS9r1J6bQTrIUelENgZiIzrjxMDexVC91HjeJLg9zYwgfjkNXZ2jiAkS62hED7mLrHz/GlCnO4rs
MFDp8h81kW3ro2tl2l+m8ZjgjEznokr/3f1jOvMG3OyE8prh5VY1slto8JEQMDKrm9jTwrRc2+Ff
RB9pSSTEL3UCa5Kj2mjxGJzLZoYyFitdlYqH5iel3Ww/L7sahPVgnrDKdV8atGClsQmJyiRukl2Z
jtK4Fy0DF8iJxu8HiGOOdE1XCY4qVnGiUNRjcyQKxnZAVl67E89Tfx+lprwwE4BsPsWklU0f0eWx
Sc5zV8uoMCPxxSXGVY7I9Aa3etZ/09j5yXA1fq5J8eIuBQzY14ZEFMYxI9sUSELkUIB9PDFi29p6
6TKVOwWu/u5TIpEJUsSyAlZhXkqSYYW1odgD19ceBEiXXwtUhmPiEPHC97Egrm8fDaH72WkLt32U
An4nmKYQtfCy8lrIfPwP1D9a7ED3bQZxFGl7nRS1t4xIHXszevZOFjG5nr/DYilRBkGyIlmN7uFU
1fjJN0RPJQZMy5irSqNrKGp504eprN6S17uj620wOR8PO+6RZtxwS2LzhsWdAl4CWsDA9/dIzUSc
Bv2C/ViztWhYslGkzEgu64jGghEBEOtqKiSIBo48zOLFO+dUAwthrhbrzmctfAHm7p4M50OdZ6bK
fcFQLfYPaINd6aSg6+WLB8XFbzZTXBBlOhSjbSumlmHcWKEpMaRQY/rS2ho2voN9LWtxUC1yD/9s
aIXvGP51xoEKMZDizGYwQKKRzDfgG6diO0BigvXy5RKbS8Tj6xf9wURUjg19Duy3OWom5v7dxAK6
1fYVI3NNT81h77BBH1QhjVYF3uH+AZ0OGLUSmWqhVktJPhbjVuRUBfyW55fzXImyGUelNeg3/WkX
zeh6f18trMNkz2YTlV1EmKqRzLYiig4sfNaFdlZvT3+r5FZdGIHD6h/lZrgUHdgGy4uGjsGITTCi
iwv+7NT76ubUzPjoaYKr+bC40wbM8Xo76mwxZf3RUnCbAEUTH1cWk7h6KDHZc3Z6uPg4zaHvzEpV
vqJxq628C0KMwleYhHk371n2T1OqX3PkZ4ErYsgGg63orCUpxE7F8u2bwrxHpk514dxsV5w4pBu4
Ca7BTQBqYOY/7meLSq5ELZu9jmbsxQRp5mbpE853LoIh29AELTd12id7lQSVXPqV3wS4IwQK+dTn
pAbKLtjbpKCHp5hO45UU9MoyjONR4qf4puDGbMx+isLkBVgqjYFe+h9TWm1xIVb1KHgGWKThB5dr
HTUyws6rGqTkeiroEcCi4lRatfHnJwIbkN9b1b7yRC3CgAkOgpB2tlIBxiCNQkNRZ1vGx0VVUEJE
vNWLO7YVEf0pt99F6CyAndWnmDXQ7SKNifICSTJWxzSwfu6GSMrqApXZ1DYqdH9c8AWCsCljG5Qa
8+Hg3xvxSikyJ1y8TiwNU6UV6cp4mtTu1G6Wr21ybvlo29afhZ0ao6O7JEpsWic/0ST03+ak+zqc
meD+NiAFcAIj6tY6NRIC6ZBRD6OhsMIBhw70FjoEM7Szzquycx/cFNi//W7pNv0GSHiAAL/hvCO9
oquA/fL6FCyUlhZjoQ03nfK2Ups0vYqIJxDdRB2nb4ZJ3Un/vq/mmo84B192H8LPsZdJf3jCglp8
RxG1i4GUH8p2Afo9vhfEMPOzGqL0/bGedpSYmOYJ2j5wZXSQ+SHYVFY5LTeJNr+QyPJ1c9fuEM/T
az8HEuO8pjb69l8toZFeWkLMG7ooa661aDfnxu5OvUDDI4XlZ7d/bJB+sw4dx75HArq8EJRB1MnT
fBQYMqeLY/+Sfx5+l8H9rmkh8Ku634AHQNm1bFIPDE+rb5W4+t0hDLojzfKzckfmUMz4jmARlhnl
kwq8N9qdjHEf3Ntg3elr2j7j8mRa/EnhB1BHwinM5cYYWuwtvQnAp1LWVlvVhDjHuPUg0M5boD8g
CwtAASLeIt7eDHg+T/NVWEgi2CivnWKa82lz7xfk1di2uYwHJG+VLLBhy0jUZT9jbk47dUF9202n
DtH9iSxn4+5bJTldBd84yu8/xXrGmq9pufTwVNcJAunb2kxrvTNvphywTQ9MvcqcxVwzSi4JNVu0
hooWo/VvP2UHn4diqLO8NvuzV0KX7gYiHfuxUwCTnovxSyrld03+cdY7d3xoZHMh8cYCwT+91YJl
7cbGkYFGh79f7czmV6OD3EafOjIHsXHnHB8W4V7STKMSTsrfAql3E5Fh++pgXBxuO00aeKFTgzrf
yNDJpI98OnoQQKn7NBH7JS6WEYc2y2y7e7jdBDW+TuQkhtkPah+M2KS/mhIJRi925oSSYAsq509h
lxn+yK7n8S7wKJ9B0udhzcgIx89QPo++YHF3XfIC3xN1YtZ7P+q0UURjxRSWxf4v/fCHUNA3+tiZ
to4c6igVZxJGS5UdL7cnpgSGZz1hO3WZTI+65aAFWygutim9uqCbgejBaGy+ULjUxkwl+eXg/SZA
xuLioSFsZ4p15nmJJhLDfb+BjteyuDDQ5qLuAnPLjmNvoKOHWHzHrTzIDCrOGEAB2Mg6bn045dho
wTqhxCBFK6VUC2yWVg7J3azeROP7Vxkzd20M998ztrLUZlWc+3cuRsuSEkwovWtSi2DH09lswHjD
zJ77Tj1i+D0lpbunf8qai66yhhmlzm+JA4X+m2ZlE2+7YpwapJRngjp1iolrkY4oCUs/cQIi72QN
vhGu1xEKF1H0UT7dNU9AmP7W5o+ZvZ+tvVSv4mqDSX0WfBtjROQiPEs+K+o1pufhx8aXAvWUw6pN
uKo7kx8awFUD1PP7aC0uifqiySfzSo1+kF4owe9xwDhTwpq//8m3TEC1r/8PLC9kCOTyd23Rksza
3jSBRbBxSU8kF/e6Zen+SCKKVd0p3+UGexvgYFdG+T6/BJ0JCJsxF26ps89/CcQH/pDsO6syNBYp
X76xD/qkMvic6ByfTVLJFvK+VGrDUcY6NlQt6O6s7Soc8yH6LCOEK92Nx+E6mQDogd/Y0lDy25II
kF8fzgBzdgbJn8/XjdSnMeNXeEBUUxWBfoWI4Xduf8+I/Lgf5Qan9qCQFZkZ8YfSRUTemY/daUBS
vWXame/uDWuRSGjQCn3dO6q0wIh9v4EQyFP/Gfl+mWVZdfoL6bJbp1l+mjSpRmluOs1+NVPKKKKy
1a07pUJ9aTO9D0QHovHZccagNR4RcnLZXER4TdHgHwGlIuNFW5evrkuDN2XDfXG08c4eE8zk+SpJ
FgKJ6IhrM6NxQixjRL6SqgIgkdF6jlWRw4D1+rcGkhU12u/LKSjp3piBD3pytfGOKc47/+7HUjJ2
Hc2JhxJBASite8633yY+RJr4FRI3T95BW1x+s+Ex4uDNu2Tm0sH6HWAMql5wmyr2NGyarU5ygw5Z
dYbdNRDRGBm9qy5lwNSYTAfdPOFxNZXem90OP35VcSfYDKPMoj6QBqiOm9RAHtQKzNOnB4gPKCsc
sT/yHo0f7hi2l/bB/acU5RL7jI0+4FZk+Ql+aDYYtzWiqJJKRWmPUzYS3xcjU1he80IqZj+hd5LL
zjZ1+qDMJpP/ln5NG4b636i5PNAqvgW2n7c+Sp12eR0x1rMK/Im+dtV2v1dmV/5nFfrihHMABlyX
wsu+WbhC7fz1o0n35eQfr749WeiVD65+CwHfMuXmfwD7DElqb2R6pki95F3zyaQ//BdajUPNGLfN
3Hb6sG6TmY615wiMIkIWFizOWGBAWDztRy5MtSInYCeGZstjzfph0BO9XiRfhnqoI8IPdM6VeQfz
21Jl516tqZFJ+PZP72GxslunWkJkbKPcKjhZWsbL1C4IEvrj3283nYk9CjLitQOwAsoWJdwgG0jr
3eNgmzHIq4sIeOx9wenrZwq+W0N0Zczb0esklMb3Xqdr4DfybPKl1j0HOOHAgaPWnbM42uDCiuTb
/GR6fpfaEWzlkQgGpvsJcs1ACpTnMTSpqEqQcNBjgbGJWRIauFgD1r8v2NIaNT+Y3vHK9ghHfEEu
nj7RYq6LVZmCXYJuMLHIxfz/gf449AK742D9GwTeusxdvauJN3KypxBaNM8xBWPafbwSteQsEOmI
jW0SgWjxKqQgtZIYjJyWTW3aJKwJiJvKT/9laHPLmyeFfwEzQAuiZSI8RIELVpg5LNkl9bMTHN88
fA5b1ArpbD3uge/05xY8Sza6Xaf1nw+wn2sAf9jyvQfyQj932CIFEfb8NeHeUGVyfR7Vf7fAzZe6
1rrU+zeIQc8fNpcWTQNp8juU4ly3JxPxHD1qEXZUxod9FPci8Rd9czG5Wl4zXEEoDZkwOAXnu2tI
D0gHwToJ1L/2d6WN5vv6UdccmixdY0YFVX7FbPO6R9g9uqkCFFbNN1U3N01fnj+99VZR3/iMlaZ6
ISInyGJpFwW1NRL4El7zhzR4Dg4ZM+6F1M9r2Pqt0FynC795wq5fDA2A4F/OimvDTWKE1fz1QOhu
JZjWWucNsymJ+FtzjkbEr/xMLBvDw/kKr1m/X3mD79vFZZSUkbi1z4BiEXCbpkilvx7JZfsodvK8
SrJUbxTiONoWX/7AnCVnF4iLDKHXPb2w41UuhBsyYUFi6yaewWBmNaNp6NtVIQ8ccZ/YvhG1sucr
CFFKLTAD62xXcDOyD9YHA+okFq17yyt/iDqJj1tKZtNEo+Ca5DrzpAG06WA/soVuJUbgfVpIfRKb
MfZ6NJCCKFcgjZaSdD4gqRhhE8VVN5pz4DBcdCe4GGh2y1E6CRxEISbxXHpy2PncPvHqRWQjWe0z
PXe0XJAlUVrYcBsXwWWUt9SwhCIjBWYeDHMj/p1stlbAuIAQdmmJr6aLRdjk19I7z5+knWAGWJ7m
6s+JT9qHBOJcLIsK7DRPlNejUopExRw2hnP+yOcsf/ZRUtjPk3torYavCJzoIiF7c68BitBaWvcb
jdtPd8+6ied2ddGdAS/A5GBIwTuZu9GAs50U5Z1xz3/AGZuS/vtwImxiqOF8oqWAuk3OK0x8+1/K
GWKFDOXGhri8Sd/a6GAl0dF+8eoOb/uhgEXJpB/vERi4wCHniY0HxpDo8I+8RWVOlIsEPILupEkt
bE8yh/NAaz2oOuwknEgrkj/6AP9HJ+MCCWf1l1ogdX5KyQ3BVL1MnQKHYBrDjlQCNPqxEKfDR7oF
GNrwKwB4GF9d46MY3t5BwXrCHYWw0cCOb+bOFVRqORJZgiOEw/8pfatZxsUqfyQDT+jfCpj5LuWC
qqisyCocg0exIEzz3OFIIZcdkzGyPRHBrB+HfOab3rfvzCAD8IwGXJo35p64YE8DEdwyE4vpdzst
wnjKz+ghgd59/QY7qm3b2FFNo3bIqCMRdJEEx2qkUVKnpL+yW1vTEwmVJkLvbAC7ADZf36Gy8MRB
bFez3WmA0xBiLDeyYbYM90FcuM4LGL/Mxa2mlHhrjSZtZLl5nNUBTD6CB8X9y8oAt0nDCsp7dhkE
3qBUmfPOf0SjzguaRRBg/p5kHCrQ9XCF/hZ2UB7UDZHwzjyXzMcV+gYDtV/bHch1Rkm4pk1x/7yt
dP3sNLfMf7lYMJAxurbrOtWrNG5/A+AVOf9Eb7ptB4sstuZHmX9GkXwK4iOeTBkhqYyiO5V03hjB
WP/ZYemeftnVICKFJTgqisQm4+lMcSrHv1noje6kB/9oi3srGqtfKZDYekZj+BWcfE6Mn04vdMDK
vF1TS/VwZC3ivIqcGAOsx2nCVpyCAPA/DMGPC5wpK0WfxI1pHyRWzw3erbuTfPNb19FWOadLmY5f
5pKrGbPuj6uPdHNPq1L6TwmcIzCXK4QN0Xc3mO5Tz2hu6Xl4Yq2dxRky9o2dO5UWo4SUzu6QQagA
/WtN+FbLM/PwxXJJiva8lSlI+N1g7EmhicuGDbIzTtlYSkLnSfDcw7o7MPHsOm7/XhN3thIHVExK
x7NTLvGhuLr8LeIycviwhDW4zqQYZX+vVXnVu/qRx0Qi4Nwp/HKYW/If1VMXQ92fdV8NqnapSH40
U0fVID+bwd/yHuVVwXZz7g/wBx+1Zz9l/2EuvOK3ykI2pp31hM4ZP1LSnIwyDHHjF/GKyu7bgSwo
Ftt7Qt+88FgFWAYPrLZGprmwQGsCRXwbW8w5lacB1HTAEmcmlnprd+4tG+6C9SgiAFXC48gEN5sx
SI1CLuZYmPnTY8CL+t0N7YSs+wntItxzCATDl3OH75fM/vhWRlPVpCbGNHLsE7Y3lBY1/SVsNCAH
S+egnOP96HEWOJrdKReucke06WQglh9YL1Q2DQuRD+U75ose1yjzDaEsjmiHr/ZWJJEBMVYxbGWo
NpyWoiOpBKRdqhFB9y34R0NXZylLref4NdwdKsJD6JQPESy0h/Age7YYIeBqnTsM6fXh0Ca18K3p
tO0L0aTBCZ3AgICQ/ifxxkAMsSbiZ1oc38+4ujjEAKlK+i9pmmyZozyh06fbak+BuXfGWLZ/strF
H2/gOC06UcDQ2UhNlJIPXVyycDNbNk4J6w2Xb5Ruz2TE+/dz0UC+9XyBgWHpK4sMsxh0eixhpGET
NZ2hOY6Qd+D0bu+/vi8Ty7oO2nTBwdEKG63FrePemeKON9bT55LgMKRLadFura8ylOdx3FSMeqqK
VmVvHj0HJlU5qVM/VKEvJidRuOzhyp4f/YzlXPjGPkoA9R71wIozhouG8eVzj9448ysTcVHMbFM2
dW/1iuPc+eMT5/ASWQopvZVnxYfkScEgyWnM4DLYRXTxYBiOYrNEVBmL0ZolDS/n/+IUeWEXIyuf
gGy69qvx6iPL93i2/osIjkbYxmNVpakWhkdaRcBpEIBezT1jS3oeXBsBWz4J6jXKKb8f57z5zMOp
X+7qE5KPq5FCWCAmAO2OykCfwqeEXNaz+gKneQ9r8pUB1vAWBL3JZIYV28KzPzWUErtgns+dKSiu
vs8jQaZ6YMaDGfEcKOZgQV1RtsqWE26Ih7ubbCpPnCMUNgHaylH8JDpTLLtd7cG8KZn1yKoQftK3
A+iyIHPWk6GR2haWOxrbjH+zPhDOdyr7bif5oK9tiQR/Jq6oJpJvd7eNlkHyAGdtCNF+iYA+gXsr
e4clxQkt2RG8M36MUaU9PYy2ESfHQk+SlG001Dlvjg3hHukQ6cI6zPcZOVmFZ3crmSiOqYrQxTN2
QKKycqOBu1k3yPSdrS+pASYEqtmK3cF6sglE0AKkDplPNz01LtrD32GylHs/EWkLfnzfYkIiPfBP
mrHZwINNEnnTvfzX0pLuFPRojkYexGeXtFAcoMUX5l8Y0bDD0BX6QRX2+r2w/Ubq4GDCwe912m0C
ajS7JUJDJ95Oq7TUi2C4SWO5MPYSNXkmG03rrafLmXIl81NKY+PoGK1KenUEsZtPzBa714lnemc5
GxoWSlgG0rt9C+xwRTq0SOEKkMaYsURxSmdKf48JVyU04yyXExelfZ/coMMoZe64kczbmVjG+ygs
kRlQeImpbr0mA+IlYvqpDIYLOSyS0v97qpgFEX09B7Qvhka1qUDlO+WnoKqkrAZiukulz928l0Ta
clamYNFiQOcmkGzKJqzG7/AwbX57Bb5kSRC2FVS7cq98+VOcF/3IKrANzPMWRke/arTFWwBjLkth
oe25wTNRF9FZhIhDLPNpAvTB+18u29F+5rYm+gLBRclxIbx96QZAdcM/4x8dl1j/Nr+QlmpYNgHO
f2HXlDirgCeasusv1riq5cG2ulqxKMTXoBQw0tG/InfA8zJFv5s78bbw9VzgN3wuhM+KTY07V/zG
DNUNAukufpl1K7MMKSjYrW/eYNJHAvvtEGG70O96LFOYTSZu78DC4jxvD2DdLvYKBnpmR4DIGH8p
HKy563BGrCo4/E/EGbcvFdcp07EGxtJ6tvFOsGsAv+ZlGBWwFmb4JAhG3jKPLe5Yal4F0AgnaBi9
sTjC+o+YIb70xaH3575VIK3jH7lz9m2qrVNFQsczmihFCSiStrUjbAD34xOVOyLPJIS9gwzAwhmJ
AH/yUGYj+0ZuxXDSjd6cjh9/J9CAjhOrFXtRlI6SJYTdKDKJ6bUFdhmIaJtzvRcGhNpHGfiRTHAW
elgFl1JrBYvkT4LMTFk30MHiPb4UaMPworSSFwC+BjCGMFZzyLE0W8c6Bmu/AHBy8qoRwaO95hVb
V+dnWsbXBuARKx7UbzztIsPW0S1fNbtFYDi/T5XUCIUYrjNo78xPygE7i6giXnvOs0qt+T4vATKC
bfpsLqeHx6TCOcLim68KLcaFMH20wRxsAmpl2LFe1tQLzVuQnDdU8j60d/nzMefwzND+jFRr4R//
2e16ZuQgWSv5WctlupsLvqzDUcMYgHQdhEGD9owNykgVAL13ur9beczLUSjkhtozh4fWywyaRRF+
m7eg4v3pSc+YnvVmon3DAfAWGve8DEI6qxkxJE0Ik52872K4aurcR+vsABRDgjK+ElOFakAPre0J
t+AeVgxcnIfLMFDkLhrEnFu3vSWM+2srosKYaAzZpv/nHbKQWyEKZnEFzWaUAXdqC5ggvM+25Umi
PjzgxeKohng2O9AEQmOr+aQdtUsXw8P7TdQWkbBOvGWclcEjRtlB3YAC8mwzY6mrhK9u+aod377Q
0xzNM6vpNV1KcqY7rwVLBHCBihh4YXzGhsJodR2HB5JVJ9SZSNXF7IibJx9pX5bOBOd6DvJ4gi6L
IFwxTpQc6afQ0D2E+/ruOoEtMvKXj6BxD1cghi+wBCsDmiXDHiZZQiZweW85JK47hhvdFX8ErmmW
ENBfgJKbZPPZtBxnGMEprsnFxOySajza+gei6cU44ltjm1fWpTSqAl3EY9n46K7JcyLzYdwnrUow
LCaRsdyuyqzqkCvixQf31gy/YeXmTxmvC3QP3q9EJ8ImIiupho5HzquuXEtKFbIn44nAZPnMgcRh
zIIRiuSBNoSC3jA/vuugGllqXfyVu4KgyHy3n3MpY2utcArHuxVLubLTPI15KATmPSJQBVq8AWFo
vnIOA1hj3MVhU9LRn93yqJXAbbVV40QKrIN7xEAQXLhI2bnARlZZG1yFijKM/zgbDSjVwDPv9gzO
1oJdmV8AvZie/9TOzsOCeBSeoiAk3Kdsp+eF8xz0EgbD4pd1K1NZ294LYTCtn9nVUHbIMrjgD0KG
86HI6QthGiq4oycNaEWrnJOgjsN3oUMQM8NOeWoCPVF/DFtafCfKh/HSCfCy7iUmG1fcp3YT2hkG
HvX1xptxO3Xk0xeeqmyo1Gw0rTZ9xkPJ4Bz5NG+lBMLrHZGzMk8Olbo5xwCVBm60p2OjyKn8mNPU
VgMEoOI/dCCwvtN8jYapVCAb3FYg/1xDjXHF0GGM65jGZzHEblr2uyk1pc1/DkGvVkYJm2zu+iPb
/lbSqp3bWYsqVl7XxpXUu0UPwPgJbRSG8MBGhI+qsNJ+z1ys4JocsMPD/MM4GPTmjwgyMvFrj1Vz
hrf8j2YvERd8pTwpqN7NnaEbkDcWvWmlz2qqXxr9tis4fZCidjqhglwpWixF+Nr3MgsCTJ399cEq
L0par87PAh8UA95m1JzNt3c+81uILQLpcMD5OPMg9ae8thNWfOU2rduX6gLVNEm4p63b1sdxq7qO
YiRO7eHjLI8k+wZysFzuRED64RNzDQxi6RKTE9ElSJn3EpLLjxLbBSIByRXL5vu9BLIiCkjqj6bv
U68tD+VRDtqeDconZv4cqUfs9C1qsVxrgE2lnY4S7bedtC/JFBHET7Eq35hrKaLkL6vAHCWhhfIo
pAR2fadpYAW3wXULyVvB6wbkitRCXpoP8C7z35DIrgu3JvDkYJTpmXEdH/AR0FJTUywLa3mlHI4W
a6FiK0jKo+NJeXPMfhalnkHAcZZA/yJk8CXSnAKRhGcz7rvwRTnU4PkORvehl24qMHhzJWsTNTxt
C/CyPo51tSjzGxDDGAfA4ERcwVyUKFcZ3EccnDy73UDd99wkCouxdiC/XwN/s7syZqFy8FGercvZ
E5DKI2JNvkU3iKWrwQq7m0hO9ZmMb34b0JkAnA0cQ2y2nkROipYYUA3E3odq/9GX54sNO/NOajAf
4OCD3SGFOpyXRmsOXwMShLwtzp69UYBYSakRk+qOIY1hKUZIYGYDwP7oOMM1Iob/6iNVpToMfejr
NwR8vvq+VL/ITQgpYlFhsP6ZzfkQdXzuPG9T461tVXKqrJsOoaQIGG8hYUmz8A9Hoke8h+ACMxPe
fC4Bn9+JiY8UoZsE79IKmwSfbOl87VErhIbcirkEH04LmOwf22J8fmZczcrO2iDRrUQfsLkPhtl1
VwJ/LA++qidaIwIzzAA4AFEWj4gYQ7fKsgHF1OkKtGhfFxBJpjyR8vM10BzBmMxaWWZSDYzmW5kl
JS+DFS3Y1QNZ5RdaW3Z29bsI3/SwcL/8nrDprHhPQdoc254A3j89rcDDpcJSSHreJYk+YuURa0tl
5GVxWnOlVGl7kjkQBVLwtKRjvBmgHHlcpkGQkNXyqwg5ZAAfRSGUMgCgXW3/e7Xli4+9HNN0kbMI
FvlfPya1FmSxl9FHXlujDYIvPdkjVPz90Q0L5y8+6lX2hAQBC+g1yY3GQiXbwdAAZ2pNiMWbnIdo
dX5gGztMtC6iPA9OWQx463WDoxiR2ohwcSiEPt6Y1eyHxQKCRYxkTM9E+MMCSDYxix4Zki5mTyzU
bCMxwKfzezbY08vVx7GsFz8f94aHlGNC1TPQ3H7/fH3WxKOVZNuRrMkka0a8h+8CjZavPHKuS3KA
CrQXzRnRcDij++De31pDiQ4begJE8Ci3GOfZbCpgXBie4UqcNB3+PXlvOE+4BHtQgXQKgVhZTGEn
3XeHAZnildhHcU8cSPv1IG2KB1JlHNbgdBqkyG+ivguN28vP1Ld9uzwbTStD1Rjb5f/05cOhHhd1
P9YKpX23WHp+s/YX118RayyITc9agzac3mTB60qG4ceSt7cowkeHDFrC+Eqy+i8uy0tx2FBNNF/i
/hH6TuLsQpJ+wlFaZxzejmjoT6azR/MiaKL4nS0W/VwxFEUxIZyhFYF4yH5BI78bqOZrsHr6PBY8
olgf4JK1aNHkcih23CWWprytq4XilQNFgzD6Z0HiyFRek0hdOUUNG3HumRf75w1rraJOjFedEZek
CI7Ohcaa4KtPH72TBpXUWqqEt5v1wEdQbjN+zBmZ/kMaEgufAC+VhCVGA6WxWeyGHV92cjQN9bxO
xnnTRAJWmlzZl5LFM4Qty8AOlRdalETUfJtvUN0ob7j4N8ZQ8eZRnCATZ11dl4V7U+mDq1fVfdfd
5I+BzsTOj+93NYyrx/4eBfSQdwJUcFLPqOs+E+S+OAPn+1AJQ1O+RLJZNFAPbSzhs+mbq3OAhhwq
2efHO6LL6ZJ4/LoIKWug2DYgV6/vVSD40wjD3pPKGa7wlYg3PUwflZwU2XIs3/75VYNfdrhytdOc
v06P3whHV0+TzRrKWuM3kGMYB3MM1p4dEK20qlr8JZ3aOPeStPkAYPReqj+kb1hGsJdGKicaCu4+
/awkNwd6/A4aawsmqNZdfcLgCxay2d8p8gJ6nBy6aoE9SF5q7MyEajIgT5tqYqtgJ5Q+iTPgJpfr
4kkWt2Y/QzrlDgF4Cq9SuV6pF4Y7eSWcGIiHhthJbZBSPvEiM8V8T/hh402c/TDiEzbK23DC/k7y
m7ffo4y6LCfryTk1ouIx0ugdPbATtP7EqE1sU2BQx08S3esPqDP5Gz4Z3LNdS1cJ7fd505Av55DR
V0yBQ9AuWbSZYH2tfrwvKgKgq4fDbBAl0be1dhvP3/Av0O7sSuGUaNNkRfeoZp1S3huov5lZYk4s
cfLeyhPfwhdp2vRMuigW0ILQrtIiRJxinPt43tox6jHSizZlOxcW/7ZCxLgJNI5JyteRfBqgQcs9
2URv1bJxl1dXYcK2CwfNwds18YvgSPFJK0yCrXd3HwWGJHrD2OggyhSzVOw4x+Q7KD2OZ6gA3oce
iK2kg60//p4OOCIukcbY4vgA0g0ZvBK95K0jgKsxzY6CPUbngQPi4xNAZ0arpY6CTMUXwQUXoLZs
ERkLXWSo2e3jnoZHQxWcr01jlTqzeMnEt9xrO/MOc8Lj8cypRzmn+2zAG8hbNM7c/U3QAcvR+hrs
8Bz+GFSwYMfiLWO2Ut9ARQhQbMWN2BCshnoJl9M7Osvm8V9EYHDbTGusHTcjZWdApzyHyIT3G8wy
gXeQQJUOF/YIZ9DM6UngGz2+0RDCekBuqdDvxRMjftKTAxFayIdHWQMuU0AI3Ym7PeNPDD7LaNRx
niLg5pfVhkORQpbas+2JKRNVeJrUUgNBv4TAfWP9LJ+MPBDVwCiBsPrDKgNic8mIvCih8sjuTj4e
0TRncsdmHNRcXJgDGNQKFfl3J3Efz5FfrWVQP2VVbu6g/8OlxAVAWG83QsO4XbWXUvjTqmTb5sjo
7NJ8joXKClRpxqaTUV/Hb0LCbaLQnawpkIn33QfUuSuyCvZadjxUUn3+5zKiTfnLqPAzBqgb0qqW
2PhwykG5PXcHeakqAoSm4Anq6DrXic1iibE0vLJLEN1t96mu0S+6pHvA6q6Fj+nLwI0Z782RS/Tb
qAD5v3YXXGBwPsz37J5WWSEn+eRRFfZXD3Vh0uGfIh3OCBZNH8IqwJDrn8p/33NKUo2scuJM1RcI
boLWW+6bJ9S01U9ZdRaqQ0P1r+4grqvlzjZBF4CwI6ipoYUWaNHwymMUweojoSdUVfW1Gv5BUyrr
FsEMSRrj3UpM/0JvIhi4cMpQyJDrb1FRznjfkRQ844IxSvX94S/uxEZPXUGqrOF+I3c9250hjD+Z
KfWELj6DRdAWPdBwjyFaI3YngQMAFR8CJf2QdcgICz9tPDDSCdZuwSmaDDKjP2YYaetLSY4EW3Wu
JWFe4vQKHRDdX/l7PHBvKYFBsxZaiARaI8veokpZOBy8Z2eDm2CoUGqQRRS3Amuxk4WF2my+0Fyk
5hgfrVmm2kc0qOEsO8Kxw0jDaiwKAZUEjt52AbnvQn9SwCfo0aAkMUNcDVIODjAhgCuYcYwKo0Jd
nuc08Hg3dSSJomBnSI7qt1lVpt4pG6qz7nRLNFfq0bCm+9GLPtlYLbNt6Mc32mx51K+aSPacQmE/
hrlIBr0D9pc3rENxXdHwJ8ED+gKXQAdM+bRaNUHCxzne+gQ0QRmEWYZ/skpF/s8BRpPhbBIfozKp
1ThohKU2rNoWogm34u8papB1dUn3k1b+S6nKmMAPcyR4Z3gJFE6zqyYB22zjtUvaEJpxI69AIxYj
KzbvnsFDj5Ljn2kZkzSRaJOkksFnQDqQ7GbzJjc1FBtbWYMZ+yoyRNQUw9C54FLOObvsZDzVUF6q
4rH6JEOH6tC3JJA2audf5m71LV9PWKv0+kFfB38yueGZyXeJ+qAR7vU9GzzVqlPlj2xAaGkg+OLl
ZckKJLXNDNfLbKSnuXD5IgYf9vTKwHkg7kEMH0vQxhjjRBdBjuTw6L7T56bLMlZQPkPLucwwvnhy
Q4srqO3/W2iwoCdwNgTNNTnr3l+Jas5aVwxAW8DI6NeT1Us7bH68rqEJyVBv3FjWZXYj/YMZ8lg6
9IL7osL3Fpio2Bk+5JmCVhMUr/seGvyOng8hK+Sl6k8xu6JLa4Pme7l/L+qvihS7uK8fMIVQbnDm
zL4A6aPLvUyvDhXSUf+0jPoiB8nNkMiwuyP+X+lj9jivY+dhcWFi7byo5vtCHX6vkwB5/8LxkDDW
+PMKWK9/CGOvNpffguiH9CvfOnX38zgLuHXd2bphsTQ8hf47bEIlR94zRvZoXye435REnVRrpDZL
z1k5EH8rh1WwyyX4iOaNpTaz0yH0/FRIwfXYUzQCexHf6NRfBBBMPlkRztceqmKSiCC+PrHktyNk
hA/UuHQ/YLaeCl6kF2jO7ZlfrRD5pTCa5NAmrzrDc1mqIKDHluNudGqPHYAfoQOsH6ZwUo1Mfl0Q
gSAtKWUSP02rzz5QZfKTJr0W1xEWYwv+x00Jg2Erneg+1oYASiNa0dPOkzFBkHGiEhL4t1epfcp/
95I8nKH35cTttw4/S2L9WVjv0hBLns80RSQkY3ncS8DkBUfor9tF0nxXJ0Eep44nJRECPYdXPEEY
0GOxB2PB4De8FLnEb64nzvwX2wY925rElTxSbpGoR5fkMvNrmRNSPTUeE5zM7dfxmcOoa1A5ys2a
xA8kx8GbIDnanlkYAHbRqK2oq1jpPnRvjc0S2wAm/sv7Zp3uLBsDClLNk+jDAZnnri4nv4tQiDtO
3JhqrbX2w4kaEoOJaz7SX+oGgRaFp/bx6s6s1e2vo1tXUrSTSih5w04ZP6XL2MUe8TXvejmKNNhg
SxdtImjP3EMEOBtSDcYpteMUJW0dkQuOxfzWnXEbZpTK46gpX/kIiVFOSJ/SSSGI7+jpV+38PyX8
sYaIQ3wuRiAjygyVQrx1MqyPKqguU61AZlOIVcDK30zcEn1GrA0wmz+MX/2yobl3grcK3a02tT14
zzf1qtY2o5t7mwDLP1zFUQfT7EsziubyXFjjPkZQMeXdIeR74jQwIg38/RXyV9gQ13Q2rBD7ghTB
7SEERFfCQeMiTacfR+m48mkQLs3vXvXovrq1aRNQx0g/smvD/xJ3uKhq9p3dMYq6NNEwNL6r3FLF
ClMyL5QBESetxwv05/WKDTiU0uUHccmyrc9LsP91kaDLqVYO/myBsjmZuA3tayj4LZ42aEh3JcgA
6RqI86LwVHDm6dBp047MpFN+c/lTeGNMAANRfxAg0dE9sXly7q6jpTBZbG0W5uv6tFGt4vSeGbpK
hm+5XndtuXl7mhjogL6Xy+SMFYER25vqsBoYmI7k9Ag7RlVWue6mZzSIlVW7KoYIS+3KMagsUtK7
4y3xZHDANlm3rGclLRkcAzAYS9LdKb5DDNkd/9PEbwaaTbm4pTCNMeNQK39FUcsxj1MQwWHAXEUG
vfOMVcq1344vhGFTJrzSSV9B4n5p6R9dz3RJSCaVqEMAB9Gt1/wST6uQEfaFe2PpSuFanM0P0Ogo
3irUrD4W1rQXsS8sm/RMs5AS+AsmtBhVi/huOqaNFeTO24yU5nLwWF8/twRYn/XNj3qfmXL6dX0V
Swv7D3M/XRuC8yTTmVqKKmtD2OVrcy9HNndQjoUMPDsHd4BjNsLbPkmcLsC7eAC8E7RqxmLkEnoO
mAByPoq5RmE5G2n5Aeop4rpn3Oa5gy7y5enGE3hsRGqOtAcu+PW/V4V2o/7y/9yLN+O7G4g41+5V
C0ENgWY15BmcAW1l8S6gMmOiQu8xA+4CcPklTaK2lUNSJIW0xc9rS7DtHAuQuhS+vP7urq8n2vJm
OItOTLrZW9F0RNVrw1IuT6r83LHcrmGYlVMM5mk+FN9TpTkcYCcQifqcSymS26c2PafVOlBriByh
f+CCwT/zJAECr2mqDeIG35wX4Pv+JXkQdmbn3tvXpKPXv0p4al+x1TUpIxdm8H9CVyDgIDTEXpmb
skLZIw5TOEcp7yDnSy/v9O33Tll9yXMqHYj0NClAEW96/o6DXHmDVQxyJh05QbA9onj60NBZNqJS
aHB9cUxQE9PO3cI40tL8H62wK5SWcSMJ3uX2MsYyT1bX6LUTflJaQ2SlgM7rIdLCZHPvIKcmF8gX
vmuKwL1b+/NktzNiJAdLLQqgbO5Ve1fi0jW1cF0mldguTTXpAcJcBBhoY/HiZ1ny168Di6aRjgEr
LHi/JN303Y2M1rAXDESkIYC2M027ZW/WI73dfPl013XKlJ6BUvvAP/KBTlOH/ShKCOBnYliyU3nc
Y4tPxVrBNwM1ZTglHYEs8fhnO2UnOHju7ky/7rNeaCheFR1ayEwxZenwaQZbIBdp5eV9WsHeX6mr
60uq+5llcjeCn685/K9d0TGNqRJgd/G+ClmOccyFXbP7etWDZqiUFB4toTTfRGICY5AvhrFX6QKr
gag68yMvDWf56OHKpB4fq0NYa4vqsKpdxf8A9QcYuZspzWVC/tOtWHSutOIdVY3oL/QTExqgMGTC
JpZ4HmXKOPbSouF2XJXvqgYQCPq5Cv0gng2KpfJKIm0JBHD0MWM+2tqQ4UapXnVS4xFaaZKLQDYM
rjaGbs35lcnDx+Ir2LjMtrxOQRna6OgLQxL3xIA8Po31aK04lCl8WDVF7adIFqMFHsATSqsRxWbt
WQVoj+Y8YRLZMfbgtUttIqv/CqCygznRJxlm7wdCdQNTm6/4j3R4xlmpWRzKUnacA3ZJxOVzpDAC
OfEOkOA2T72cH8Ki9RS/O31XXkVfQsGLHYsPL09pAnLcIBkxNYEi+rawPsLGWJY1iTI19VnoMcuB
4Ow8G1XsAoYazWyJElTcRqTl9aguEEf2fYS1i83ylP3XO4sglIWoY8E3x4v3Gu0Mcurvx2wN2Gj8
NgT+tdbLOcJbx0vw7XDklczn+Nh3nPHQOv9IQI9QSTwmVQMT3NSEg9bztR06Qx9UIGFlwA6pTyF6
b4GDXJiBD1XCZpk2t/HsXIZZBesG88VM3IpNigK63MmhgAAUv8R3w7QY0RAv5hcPM9X26iJ6ZNYB
FsD5sRl9/p3faJbBnekFej08WAfRJ/C02+Xd8wOzLaCZRg5neK7duTV/3CFFc08PD0+XfKvujMzv
OKlk5Z6fDTz253UcEu4j+tYeJcOuoBXCIK25jc9WXnFcQqczEe2lVOBKAW+CQ62cHsfotMo6+TlW
lbOlwevzPGvGSdwKG8W4kOq490yquBUq+0ribwWHO3Oyp2QtcomVXvXqlqxxg3JBiVpB8kYnhWJy
4Sg53vVlRPJHtTQnOLoTq0EJHv0jQoeGeygFEKGTsR42UI177liIWWuSOkG5Dhgs3aCXYLMjoT18
NO2vcsq2THOkV3yLDIEokaOxRtOeZatP/4RLu1feR5/dcYIf7LXBLux+5RhB55svzADDgMEoNnOs
6KoHTut5tXuCCvq2wklyqo/Hk4oYS72rKqzzIow4D5rXsRNTMHtRA2yj/Wp3lQ0EA+NyJFaNAYcU
w0dBeg88DyqoLAi9B3qM3nGk6LercP5OeiAevRp+hZcyQfYI4V+n1g5fZYuJz+Ym4uJIOacI7dOa
75XhM2AQjtXyqN+hSG4WJF4ljf1xlMC6P537WdJ0atyWZe9FXVnoRogge5T9YdYfZRhEwBczHbVs
/rY6acBnlq2rytSFGH4ZI/QB2UujOBJPxZ/Lso4kytJ0q6XjB6Ivxj14p8Z5qqLSivjiAX63acni
KSuGP/g9rZ6hsQV4MUkkd+jM9H1dwnKLrIwYGViIJ45xdP5S5N/witanyFzcroEJz34ythjVkeAO
7Sye3fhnMWdlbvdm40sdxDuCpHGL03QSBwQUWXEriXZjwuTjgbUe/27JprVlKobZt82OWGoL2uYG
4bt5nufEvLuY6E/S9WXfUjDgq6nkWkR3U1fsQ2yEujFQYESqlrF/cGMRUecvppHpr2asQPW8FJc5
ESZIT08I1APGGdUdv1IgZ3yIRE/hBR5tEy7YKkoQIqBb2AWRwT1SmU6tUw/DkmbHqLZlBJpRzarO
RPJICbWNcUw0aJeKhPKavuxITWuJGBX5CYN8JXt1d6NdfBCk/0ZxNXucQh6puSDZw6yGdyhuUaWE
0f5Nso1PKtG5qIE+Z5+yEnaWfKqc5zIbLouzBojuMTKX8WTnm1lr3BbR5t6m3pqrSHmD2rmWkcuP
J95W0j2Oc24himfOmE0xSv3IerbEBvu6cwO/r/PLInJFWrGHqhNzne9EfqpMR+88xf0ljAqA2OU3
JDuheC3CSjHXgCYwjK3hc2YCKxzRUlDbWl0c90VIxv/PFH4wJ6PYhEXfR2znUNwq+9up4cvVgEh0
68a12XBmNAoZJ5mkCKCYj3LXnHImjUr6tmI6SABGIrUMIMBcRSnD2ZTGEZPDIRiti8w69Rl+Mch3
KIUbTP04tCl7z/zyQfXMc6TV1kW0Dkb1JjmFzqIPJK+B1+OnIf9sjDCgIk7dUcKkDuRkHH6dGG1m
sOAXj1SLmhJck2y4XNFM/+zd2px1+1j4D0Y2IodOc6xYLI+GTpH4YI+FvDTtKyp5oy9vVh17yTLv
eaEDtxlSm5Q+C2EiUnVISv659bAZf3RSwFmQi/FXxTrrYkC6GzVy7vQ64NNceNwVpLKYKYQmhY3j
EErAUa+OGDWsIg/E9hAS8/UBaOZ8YdxHRgFLTAXn/W7PWV2p6AiiVRr91Ml6FCjdou6vNnw3CfXE
JmocWT6zxBz+o4U6yERys7u4sQCvZWST3xAWkIRM+kNAhVKyXi5muHT6OsiMmu/7rPTSyQVd5Nkh
PGppCB/5t0gKzL/CJeLTBjAiam3jIgLWxSqMVhvQAKLFdJgSz3MeZ49JZpDi2zg0SpsWmRO2u6Z7
T9z71TSYJdO1DzuFIIv+Mq362ZvMadETFaIRiQdSS0MhyIupdBsPuoOS3okLHcaJS525KA3kncPm
fqAFTNwfWGUen0EZEV3XkE8aZyMxB1PvxL1Si2pwaaZ0ZRwHTc1Un2gQGkYKmicl7t82fHbYuNzg
3zoYRZ9DqGTf8rA5SwBd/tcjvn+0F6uqOnEOeme4IxoVIyTB8Y2UT91uc7p0eecEgEwUkP3UoT/z
d+VUwQWw8H+dS9gsFDpfwstywqbJ0yNJld4tMTV0AM+i/8kMNIdOLl2RGCqulRaLtp8kw62ilxOu
1qt65Ay2WuDD/qUjEKM9SUr98YSGBkjXju0SZFZKUgiskAYeyonA67L3MnvEL0Ye4yqSI/mxT/tq
StTbk3D7njCQPrUMm32tfkzOXzuIAuhQmV7ZbEiFCXjYGrD9a3vbHHTrOyHZU3h7S9p9gWezS8hN
6n6BSmatF37+0XXmUIKH+1t7BaU2GABfD7ee2VSUaBpHKCysgLDQf+CQ4Wp5/KCPqCfXfi7dK5yE
AQS8OUPhiC3QaSotUP/37MeJ+IcBGM22dqYgFha0IzKEKniz5j36VXfHRUq2bv619wYO6f+wx+4P
PDQnqgi/m9W4CFWPPWuryxmWxUsaqj2huMne0TEdvu4vLokiupP6IPxnAk1nI8I+2gwBSdvZcKq4
vpQH414V1X/+NqbYLbdnfDe03cGH9qREUkNDVrKbyy/l8Ct4V2w6d1Z6dpQX7QHjCqIzVtkt6hA9
qIzmn2ouiKlX5TO4vk8S7UPsGd4zkr3DV+HroGp3aVa+Mou4B04a1xPVt5JBirZIxCZ8L+wlfMFA
kEUD5ZDjrqEPFBjj/gUmn5A6wyAFt/PPtIX5Qx0U7r/YVIxi9mH8cpqEwStTIAwL+cp36McMrIo1
D+amXmy/CAMG4XWej/1+6xmuThJW7NHvgyYn60KbcS1yj4TeKvWGBMjo/RCp2XwAcZ3c29h3hWNM
h8zILSHe3DOzIbLPH1TffFiLkZvzXojb1OXzD4gM0vEzbaBb1orNLU/CoX9VPPyJSEBRcKILrDhl
HtS0Xf69jCFmkq8VVS6eMK0khYgJPzthPIcQekjhxDzzdWgYQO9tk3w8T+iZhIsViCmo8I3sOkUd
5rzEMRvpKJJwaRGqotHQJCg7WtFhLN7EKiPyMSKlY/T2b0GrheK5rPFIYjLWFozHvrnxercsCy6a
Lsol9nDox6jPl3sifGqgEkK+Mr1WaCHDFnqQPhcS9cw9HDc7gxiIbXtU3u5SPFtapOrPMcbv61pO
4t0TyeKUf2Isr2HCD0g0W4+QXkayNYDkxEig09lCvyskF4oZzuCTS0vXnLd9edghGOvZWPTlDYSm
DLfc+CijiqBguEmb11W5AA1a9HOfPC44T2mbUGPbUbruZjxxT0XbaKd7wdz74dktE+WhYed5D7eX
Fq44GKCC9HyCv9SnOHWenZlS2RiweLRGJp/I8XcWn71kUkHz9l9CbQ+jUvxBS63w8vPnCbgKzV6Y
KDZ1rrIjK9VrqbZ6VHiH4yyMskzl5ossL8z7tmqb36nI24gg9io79OvW5HfGOargqUKmfY8zO4nG
6eEVBqiKO2UwBghYkSpiszvlQcwgoWAiQgyjBFadI7T/CIg9LYB6rOlvAOYBwMfeweKHnoFe/Eay
LWd3A/Vyxq8OOLkarhru9q+rd+nD+JaeO4AlS59FJRHBf9ZUZzzifu6tZri8lyRg7EeQq6EoUVjH
qp7HFVJ5Iql+26o+aL6I83yFtygkfRjxbFoAQAnGm58ajMURuF6bFfT2gnYZorzyDvh9/3XNd5xY
I4nLuBdWDWNqvluMCWn2Vp+rGoYXmrpDa4XMsSRLC/DKRd/zbS1pcjvsjfgZXyQYQzWdjUwfgcuP
rfUNUPfqWlCVZDtL2rxZ/Vso/GsloLPudZyCRnTHXvNVCzMEprBdyRtAXmC9LlbD/bnTTAroUFqf
7D6wdz+dAnpC00zIUONZk1ID6+d0LP7GcuAvlhd1FtAHxzraY2WHxBJJJYYdPzOFtjG8o21bJV9t
mB0lgUNniOvNLSgOghBccE6kk5shkCYYep1ZmPTN5EWJJVrrZiOPl8y6h9Q48F/k+K8V4bfzcRl3
gO7ZInte9H3ttepg7wWnKIRUcAcZ6Js6p1z4nMSKmMkyboTU3tVAR+0Ce5AH0iEAFrxtnjrtkz6I
Vbod+Q4JIEWzn2Sw8mQKSU5RaHUpFxmoif6IWqfoYONpRT23oPSycjkLOXux266LFuSAz5w2v6XQ
OIccshWs3r77VcBj06UZsMGoouS86LRSM9egY9Jl9zt3FMuSQO3mMZIGzULhvB2kmF4cDbLeNBpO
aFacmS1xulSC52QkT/LXz142Z8Vyqfdn9/f0ybPAb0dBFq7vFO64hdnIBI3QxIkzhQKi09MjZVPy
+rxdoN0TzKA5uUkVFZXtTW/cbWG+VOPpDA9eeqv0PFYoVBgoWWJ7RbNxOYDgSXSMkbPeappgJn+w
okiBalvxokkBniA4KjoOD6amwHU2xMI2MqQ86l2gduzRtH9u0ce9ZnC5LIKpah0irzbYDwfG909Y
bvzjPPJSbDpebsUywbQetRt8slrFlazSOr0MMjkGlttqiEACx7bkgM24MK6EQ0dZpLnmQNVURb9m
w8/gxSZITdww9FQLO2FrM9qFyWiEGFM2zv7ALoBnD57rrYlItvguegu07a9BjL6Ht2dGmu6tfxZ8
KEazZHjK/YBl5vU2LGPFxClG0ZYKAWkOufz7xKKHUiL7FAEu1o/dTVfqWyJvDMbt2dojBE0pYT4Y
IhWx+H5rK7fZX0c59Q5dxrgMpXd9NlGFhLzm+Cd+dz3X5LsqhVO0YzFpdkdcsc5olgOl3ywxcmvd
5/WjjFb4M62dEDVI/CzObkpuTZj9oxUkisj6QPi97LBVhsWX4QIvngpa4GiWJALiPZ6rJOURoJqu
NbpcIzdmj0LxkFBCi4pmXknI/+BPOSezDlu2FM7h3DTwaeZuCoJCmIxvXUcTeB+D9/C6ygYuZZqC
L1NTmbu72HGEy/uh9sRLj7HeoN1NQV5T9FiLi0zvTxf3YerzuajEYpm1aeOzvleC0HtEacuAkOYV
1QqRb6F09DYUC3TYU8Xcl1kWgFKfH0vUpDvgpzk2rzO6p7y0sUankBEIUvK/5qPLU5IgJTYWTMty
cQO6Do+bhlIk0ICsSEoXlNSuQStBm0uP3qsfJ7IfYtFu8mcNaproUXZ7u2s5bSgjdSnmMn39VBTq
IIXapjOJw5Q8rTYJ2RCTmGnwhwsA0ic/GEXwmnd0lqgBJWR/HHGk/8RKGzLUDnUm6UFj8qeYh2MS
1cD2BjJ9PKCNNmLlk9mbCb0joUOECfzAcfe6EvGDgrOE6bocuc/ymiSUqIN54ohnoAowOdtdVTe3
3cXZWX6GVR3nZm2LjQFqFdpz+l61HlLy/LA3lSkeWPyj1U+ruBo6/90RioWYb+XFJvnHktR9VLTX
vW41KkDTU9zIvDgqzh6LLImGqXwEVox7IecJHrwzw5KrhbF5aoQqyQc9H6sy6IT3c/UPrd5HMmHx
qLbPjIDRsGJsD8cz+CBzS7dHzazD1UXOhe58oeGHpX59Ce5bVvYWuL7qyqQKGAOYKCpLbEIW7lH/
4tD9mU8T0yIbjkDarsLKtocIK3cubMUSTpZQno2zWX1O0OtZO1dSLTfwIaG8oPl645YbI9GDEXdF
JGOw14jvAit6zAu63JxgeRTHZFynLDyOeBxp2O++4eJw6opDmraZj9dh7VEpPzDh8l4ihzCpXzeD
9/XEswtrKr0v0gC6osDpkrVpphlSgDHwIyGk1HyDN9gX8oxCa2NTtfyI0bMBphf/aS09vCbD0xFp
Xr1ZOxUy9x/FT3RrG3B/nAoMNE5HPabLcpjByJmtm7ybhauYS0v1s44DIH37xb+SwxNUKRSZIjYk
rsOqAwlKVyD9HteS1lg1ZDrki1hTzBWx4ZwfkgB8sCJ15jsDzoT01at1rgITaNFZR5/HT0coxxbl
j2JGapPzVBFnsk9syx6k9rWJELlVmbVpXE9q/YhyoPJ1jO5z/zLlUVeOlkvxm8OeyoFaPeUDinK/
GRu6K3gwIfYxRoY38VQ5/AvgARK8Y8JKJ5nn93YLF/Guko3OsWy838M+A9CGbB5ZQrkjeWNifrVg
S1Cwfxra83TUXpbxsJcILIwK31A9HvJVKFclWS6KdtSLfM4Wk5ViI7MzpsDmDfyUf5il4w6SP2Ww
WqoBfADWNkHLmcO5UEeLMoPREs5VFJa2EUWOyMmd0oBnBvoovUz/C/ZuChns3C5ilUAkZE7+OrZn
XXUXl7tFGf4b7T5wFKu4tYULkwmL/EIgBSTdd2Vib1WbVtYbdE5QQwLw4KV3tqYO1i11xPQ/00b1
SXZJ3TTtIaqwXy54kxL1azKHyK4Yseo9PeDGC5BV2Q0lLCYXhHzalKqxq/x7bWpGogGScOGv6yR3
5uHH4DS9Czr3wlzUKlyeMkp+EMA7RYs/zUGqe7XCt78S7OgIm2BIFeyRaIWz7/1dt7UHGsUZ91oO
s5E8dUl/eqV3D4LS6Zj1chyZSFCjdOVFzsJxYD2kXMe+Kgc4acdBumG2Vthmtgul0DCzvrrvVCtJ
If3nStRT866P4EkK0ViVJ4yKaAwj0GxfBNY5JiPkUikKlZIhWVCQYxX/mh/8m8eSYtIKhjatJfhD
oUIwpl0DuPCv1VDuwwzQcrwNkWAq6HKzNvIqSfTub7zER9u69Q4lhH9say2Zb86YqT9QVyc2dAVw
2M+bGyJN6pvpTVrYucq3k7HnZ9eBqf/iJmy9DxcOsJ10kRnAFyXl/yCC9Uh4E1io8RO7DoUBptUs
fILzkyHRAyftTxVEe7s17+YBNgnWeROWaNJF4HsWUBlwKGle/wNHCYlLWwibLFRFxdjsB5N4rK5V
61sBs0Z+axzru9bSbIxpr7HKGJgDjzUu8XgD08bepvumvMOgPaNrqABfVQCQlSY4F6lDCT0klLp8
+EnMkq9x+iQnCz3/ftT+fo48qGON940cSnDBW1XCv8qPQBu93JENUnnI9++IT2D2Zwx4eDn9GXs6
fPlu1Ld80hzGxUyylT7NCSPqIdt1dDlwJuW/rsnedsvevsC3h8yqgJJOWE8Z3zBQ89baDRSLvILO
YuG9JC87ISbWTcWetYQx0Ts2zQI363ZEfV36kZVdjX99PH2K4CTHwtcK3UkAp+gL6z8BPXqtO6LG
WWoKMJwNhZac9wTCxig8dY6Mylj1nwn1R+JuT1fkgh9jN+Wzt38JC4ANPwbcoVikvdnGDkm4EE4c
hG8K6UTwpHoYgr2/XdOuQn1kNZ+7NrRH955WB6twfw/l7PI978jsN6B0FhB0KP+5wSQ8T17M9wAC
dNV9ycyQGSpz6BHDi+AUGNuhztfB2/Rn+LIOrIQM2b5VYUqOoifWxQD7ZlFCrUvIUJCx4TRI6d5m
+QvI1iOt+1E/p/ltBph9s3o8ZKNEQHV3sEnPFRxLh/RMUXJq4acHoadDbmxjhU6fZbeRJAME3vV6
UDtYzl6chMNXn3g7CVsxRHmGE7fq8hB2FF/LAbweEUESs6w7cg+hSBVdmyx36XeXNKWadjerqNF3
2VKncZp2suSQfspHXm1LjwLAfRUKHviOE78Gl+gsLlmC8gTfagsspoDn48l6bHsDPH3D+6rpCD7o
cRwxsjODrCVxP7/hPXq88NYU0z0M6b4H1p7CpV1Y2bEqx1ZBj+wtwcx0m/dfdVLxgXJALy0eWQIu
zKs4Al6Lt0+OsMw5ICQEZyHEGvuNBLYipv87sUNFlfNhG4vBo1lF7JTPeO/Aa2O/jv/FBv4YnZky
z0a3J2id2jE4RbQtSuB9sdOQ8a16uwt1ZziCYg6gl3wnj3njnnwEtg1atUf6/s+JNJu8TEDFDuYj
UbbJx4sC/KCyNdn+nf2G7yMULgY0RW3UxfQJH5r3i5YJtOCCWbOnm0LJdpGv92e+6uJVS0b9YVO4
GH0cv9V8spYdqExhruJ9l9rzcnvYYGLzW/3dhTnfmL3B66s0FZgP75Ma47QE5mm4KYTFZkOE0h9O
+TBR76R5JqdqdcAWaAN59MUOMOStstlDzPHwxNCJxxKXtPoNgDYiZkPI9BleNdac+C54t5Zajzdc
fLpLAYRT+uVbhBOQNn2faZ5Yk9i54HC4J2YHAuw6Fz7rnodvmHmEVxKtiqEHtL3ejEJKEuwXEXqm
6UqUdmtol/VZK3FJbksEqQJil9RN25a34/2+AnoVIRDHdwJrfSEPLHVTe4mPNZsLGwPiZ8nmXSmS
4+G6VrJt8wAJoJXvaXD6tsON1o2H2NiHZt07mJX9qaIpdt1nYh1mUoeY7lq3KTcIfdraBRBXa4pQ
bvoru3E0+YUmvGGgqfwc3oUt1PvUWKXAKK0IGrEI5ouACE39bCW8FT/i/L4Ddr9O/vaurVxupFbB
UL55816IQggLHrw9YXVsTGFR4wfIDU6FnOtqj1EnljPFXYA8xKDERLnNuxry8iW9wDkxIBfCKiCG
k8M5eJSmCAcriRxlPumi4tXp9ewwOKJY/Kj9FL2Udzxg4AppfbK/95hNygqF6Cv/s9iQQ8KcPAWI
pBW8qt2VGFe40eBRw9yYdXt/4pm67l33y1T6pcxsR8yt5vSrxYDxQtncwofrxIbefDa1Qm+rEP/s
OHsKT62ap6JRWXgRXyZjD2LmP4/ZxtZFwE0yO5qrmzVVLs7Bzh8hj5jiQcxsiFYTeKtPBYmY+IYU
3BqodNfNXcCraV8QQwBpz4hio/QOHPmr4K1mQQaE/UEAC+TozRO59YfmqxOBgLRwJCac75NnTv0S
vesDUqrxayNN9m/bnJx+VT4NaZVerNBexfS9vb0vZS0K988U5c8QDxwgNmkUygKSI7nExpV3L8q3
d1PEWdlCGD/N5vUp4z8YDRZ1hqopm0tVnzEl+LZ9x0405Pxjimei93OMoh1c71EifRLuK7YAv5jr
AY+RezNUnvjYGyRJZbXfI/hpM0Ac1YYzqYHg2RsLBvUjnL4iyvak9xftaWJcv54BuPPe6yiA2F3Z
SsTF1GS52p7eUoNMWdTlvbcNRQHD8aSP+hCTK0bEf6le7Ph7+0l9I+qYHlcbaGU2IuI+QE9FntyC
uW0H3ddGa7j8Ib8xPCtHfQKzmmcsYRXjLWEIeUa11pbxCqwYMwnyBjYNLuLsAJRleHF4fd1S0CQ2
RfOxzlUIyqImVqKpbR+Gi0lkFp7XCjeBbviGO3kTo4DKm3LY+Mdch6CcnDoyuxo9m1Y1IADANi4Y
7BFLyw9JStbxsnDEPxeUHUz2QjFni/NFg3P8/jTcV9IwPgPWsRaqDS/sVvmbOAxE7/5R+sT6ZhzE
A0vglhb6mdLjloAoPo1LS+bbDHQQem1PIRhEzDLf5pFlWxUHnr+c97X594c7gGXVq46fulwk+Txo
i+4a+YbCOHfxczFyjLr5jpCWsDlgAMfCbydEuixtCnwWRdCY7f1uIPyA5CDd8fFbvhZlKAmcT084
P6+NQbqkReHRXN/NEK65gQvj2s6gXox5V5CG/ejaf5hxPlkNsvt9+k8T7NsSLYblYbc5uFB6uf3z
cKk8AmOTZvkYhXhMY+GF8qWkJQLnOy9+MNzOIWpODfdlO9tzsGwBRaPClpANm3iAVYxhP74G6QEJ
9ILFgXcwsXrouy7zSzmxKWFEpAKxW4cVnn0H2iJSbqTqhZhaJXu1306bdtUx1qX8W2bUXOJ/p+CA
/GpXXqGQSU+/5tSlVbdnmBxg48wT0Ky58arRWRgl+iRgNKd3ssytBLFoLPkwZ5twmw2DV3kR5nXf
NUaeOXrvlyrKqEHh4RFp5Xps35gXRxkFm6UGBZaQkyqlmKzUIXXB1hr2lZ7kSZrL6Fua8G22ua7p
iSOHaPvYJ08hPj6Yz/PuLkOpZb+yPa2o/bcahSaUJmCSdSldYqQXd+OqW+qrGXIybmfiRpd9wh4y
JuzNIcYXIzq3Q+ewk9qZM8Hf2CRIjXJ9/rJwiUiFy6uDZW+rHPA3b9BLAX4boCa7tXShkwSpKdY/
4QEcz5maBemmy+x48jFMbywfKS/ClSr9P2h871dUPfnsJzWfSYtamw4qbENNKJNkaBVALEym9Cq3
oDt/V6RqM6qlff16dJrHZiyZS3ffp/l9aRGoI5y6pcJL8SbjijF73mzxN3UQmI9opBMZxTTV1thE
aNB6Z7TlxIeeyBxn2//V0eMNdY8oy1cYPBrJdX6sZqf3IYxGCtMn8xy9k8Kqu9kni3ApLQ58aUgx
QT7M8hv47fhr+CuXRNqutRg93tnmJS00m7X0PYn66K6/XBvY6L6ZCjzgDStizBGCxlyvL/TD3a23
ndpDZ0fQ2di09ahIClJRLumINivXrXJCslegpttZiaAdSSZ527jZ3nGqYX60PaJqfbbJSZ5BGcen
tRd5adySx1+x2KZKZ6HRNcJoRHmkXbWQlmDm+a20YmN7hkMIZWsD4YA4ZpYNDsPXg5CdSDPZBR5X
48da5zzBOF/1FdnUZKyMygemzJUaOOc5EVsaBVr47dhJ8kSwOO8hu4EdNTTkDaT+FranrqJNRvNd
l7PfF4zGz0izM1dGXqUWv6vWDIXGfuzJw/vV9ucQ9Zo7OK9ut5hY6cw1l9yafuutZGgybk0Emt2i
nkMr/2JFeO1BScPN9TjLJuSp98Op6t//2TbXRMBy/WCMXKWj7o4Z6up+yQGqmWD8BWjraUYxGZEr
0mFMXNRCBFtAyb06+uxeoFlXCNvAEgSeA2XdWd5F52goLe0St0wsJclHfuI6xk1pnhCYsTUMo2pm
oCWA9MGLt6N6ZXceIqeZkCmHwJsGTd01TbxJErVz11W7hE20JnY6DZrBsNT9OfwnAdaJJmJXtvSD
tZauHSsJtkJ9PGhLEqZd+Y3i3mADyHEu18YwcbKkPq+hy0vm4AleQlLqABEy5MFksTpFfBDwO6NT
p1S7v9fkoXNUIPKS/jklKNQ+kqKErDcMWukjdhnBf/wZ6a2du5KBSDvLXFDK9LF/ng+69CoTDr/b
6rYr6Orn2RRxkdAnligzFF9lq9wnG4hhVGbUzhXbel8Ww8OU7wRYZAxqOHqUhe11rZzAGIO5kshA
JP406V5/mScXbBEwGw3CH5cGPJUK0BRBxCie2wPmT3ocdNZC58Rw4TX8ZoZqXiY1AszebzijEtZi
CdiQwiWjHvrgFDTWX8/FXTQ1fHPcWUPWlGPqxcpbN5cfFUmg58jAczixGaiFVSwqElLPERD1On32
eCmscaHflPK5gsQxdDlaICzRniYFUJoxdVsWaaQ3qMjRp2+nRM8LdSwEKry6ChuPrW0uBXUFT+Tu
KpfFkMEQpSsf95+Q51XIIjGEOGfrgSyQAERQWbc727ROLTps7lyRtOSjn7W/R6L+28JNAOonO8GO
86YPU5uMcaAsfMm79TSIKDyao9fFNCukk0elofX27OoFJ4m6a9viYVgqWNaUgHnqbQ4O4drj8sah
58bu1/VR6Cu1wFS8AAgE6ifVswkkjhfOerjp/EpF3un7uN9d+Ii43ictWTjPbvk2S59hSU0KTs4M
6Bo81UcqeyIXFEq8j7at8zaosV+Vl0XFCiCrmW4udHi3UiHS/VeulcF0Srm6MDDOOhBOh39AJi10
oCEWCUmk5cfzAoCgdNLshnYay71ogVYiwwyyOmqlZNtKcJLw1dEFIGJmYvKxMOD2fGfw3TJMiXKE
kSX3liB7SpgrliEWjHtRRQsJJtZpSqRRsgSHXONOVkrUEYP0iMOpkx484Kf19lVTzRdi2dJ1lRA1
ZXwmeY4FXW+tcYvoUUq6erruQuE7SYnJPK49JHrAgGnQUxy6BEYfzUm2vMppXZzT5pzGP8N9tffo
VV9qRxYtOludtvd3RBH9txfEPPMq9UsezfUsfdBQ+py9s8aow4OVozEcIJh4nGKg+XrT41Hne5FK
ZuEhFGL5mQyvngprbXk6hTAmsUJCUYqXxnk921b07bnnxJnn3/k+uOo568UGIysLC+3PxloxDBGm
YsWUZiARbaUzLkCtQmTAEW+lqzfJXPY76Hso8E+j3m93PvhjuPIx64s/daEGOUdkuoxapsqhfARO
vg9suo9SSKZJ2riT3qvHoMd6mok4KAVGE2be2e/RDqnPS4Oslo8RhDf8EIP59SQoAGL3BmqsRp3G
0gj78VBH2kNXvre5JibE1pNHh8KyehLbQfi5plDtAOinscsdE5+gOYqzSgAfnnh8WBbL6rvlvFb4
SSw7eh+yM/o6Co0xA9KeFu55sn2zVto/jCptUwO9YQQRHaT4wsQKvQYY2lyUSM/CGYrRbVX5v1um
E5JoZiKu+bvK6YfUci31+J9NIoCXy231xlmfJ/xjuK35tliM+zHQZZYOI/NR7Jtc057FdpD7LHzX
BggW36mAGDhh9XEz5qa5Z9Mds/r0HRbNdfZ5Is9qSXYbEY50msDnAnwWWt5PjhHSj2PYfR1pOHle
NEZu8AL5sE5UkLbVBg7wr1J5x602D6KYt7EZwCxizBpPkfSTDzGmx4vEpNqFTTpQDrzc1v2dFxE5
D1I79GSsl+pSlgcSPSQ1tieDzkN+JZlvCcV0tJ+I28mUqkhMgXg+hAApXtAEpggGk1VFljZe6h6o
oe9TDvOQblpZzatBKEVB/C5CF/Z6hfwBWI/GBafQynFqnxg9o69aOde0ba4HHYKgddiaIDA1orBb
IsDY1Stpq5fEDihGvHL+Co/GBEjfm9eTPcxArh47Oq5hioVL3JpBlNl/u93Isav5CZjGY3K5sh9R
rZ9OhluawM4sgCKH3Ds30mNccst1W+ltuzhzvftzX342auGjHBHo/wdl3vA6NC0hIJoIchKwcrVC
TTbX8umHaBJPKITrv+V9hfMtdFhftUrWG36oNhpE8vOSAoP98hSzphXLM3wu332x94zzZ2JiYa82
jfMGz5rB3L/34I3CW1xXAqyVvKeUgdcCZK8KrleUByARZr2+73fc8IMGGOaKDJWeE+xVZr7gFtpj
9guDwFdMY0NScBHRmtweP85opufxRiIFgPYLHJhz0ANv+oULCPClDL4mIbSLrMDjsU6ceLZovb6U
4NCh5CXF5aHhgruFFQLiEGkwkV3xjNKT+WSs0+9xuCzaKD3BUUzvfoUYYcVOqYuKwjKMML8lMPOE
0+eC4tbx0j15kFAu7QIBOf/1DWCpHS8V9w+Wu3ldFaSFFj6sNYEUyJQ8px95gwqAp6Wo6mED+gaf
TlRRwd3EDKZUFqZry957RP4nl/kvFdHc0mGF2WFUgrvZrXg9xRR+29ltzLmH1064LaBxRMjoo+ic
p/N2Jn0sjRX7qOliRp+AiRD/4C7/v0xg50kSGbviyZCDTieij5F99wN7KaPUDc2R4bKBzqcbNn7z
ri0y89iifCvgv9gWjrDzKC8IbfRGOD3mkci4mc8rrHePzUSIM4X8reucD5Q4pl5FISiv55EjebzU
F35WRhUMYeo6pgos/62ZF2NyfTPi6YTZnKfNNpPmfBK4sUQu/btppLWvQBXRZwKkh+41gQ2CurDc
kUpGaqlU/Tj+z7BQlhqKhhv8O4TnUOHa5A0c6BjYbIotVA2WS1MZ6uQZOmXutYQFeFFYHDbNE5l6
uvhdlzc2dtUJERXTZmqJil9oTM1HAOWS6pk3XBhN/w47bH9sdoN3T/oZriziU4r9yCuZPxn/4NgZ
mk74Mum+P+9ekxHCW5hpRf1JumJ6i2oap64BBok8Pf8hk0UJgAnHe6p3wrcRkMqPxVoyV6l0Whlu
QCcFCqtYWeqWKyZZBpM9kO65xtlYIQkbd7L+vXM93GENl2WiYVa2Q1APLd1cMXYR97tJVyfEDWGk
gMOhxVTlnG5AXbM113a31flLQaUbLWDCM365DqpE1EpqqaDMgUbQi0HVJ3nCi7jcS1aWV9LeWPf2
2wQaD06Qo29YQL+ZDHildDTHLBWyDyZCItILoieY8OO4siQqJP09E/+10k6Tma705PttpB8XobPL
+rM6wRslHmlRBXUkv/qc9tlqYswWIOcAVaJMrTH5P0+CLm06Z+UIhgRv4JPSd4PakGl5T+qyh8FR
aMJawLQ8g6MT9Pkv0FPVuVJd36oFPLM+dJgP5PcunoyXuDkrzSJO1TnmsYI1rgiaGQek+b20BwDf
iOLcQZ6iuy7i5aj+TZfs2N1SZDy7X7l0QnT7GSxXx/s6/8Usm0PqGT5b/qZ9snYJJcvIa+yP5zFJ
LjVWEg9j+Kh6WZkjTX3lfm4Q9QEriEU9SXS+fHYEKndUe0tO7eYBSO3OTzTbaAU9/yBlw99DjAdv
DCzKMsJCHMVbwJlrf52jDCsF4a3/kqZAwpLFIrmBSp3lXSTuBeRHwg1u1+EmGq8Gm3ZH1sUUDBIE
ZpOeMUcqTl3R2ooy3JDgKCHw1b+rp0jmVRSHhb7Qt0nkJZ70GJ+uhZ+E90YaQbRLt08qHtByW0iR
Q5XdAUZPnYX0AMtppk0D+JBJLnvI2RSeTCSbuQRsCDvPRrfdHuyR1613gZsQdFQgWRsLI9b0fKqg
myRdiSTqed9dJmKRPD6087CsNUN0HegpHOAH7FtxPRg35ZvtHDe1mmbmO5wdqy/QxaAmtAb4hRPB
aEGUyQG6d1CoKhSfsyzkQJ5Nptt+e+SaCDHjqhuW6VnceHbeLXZBdNejjCTI386xC3Ck94SPPA2r
ZUZqQtmRq0R48CxelQTqTHwHArPQqc2Hx0v1pIfoUHKV2szlrJgpHOaaZQur5traKhorAhRewQMC
BsL6rlIMDznQnhfJx6Q70Wt3Fwl4LExWf8i800gQHzn3sOnjVEsQdGtfHMQl4mQxwoWzT3ZmrJci
gTJ8d38G/Xzi/E8lkPy0jP4U0676aDNABCp7YDI0OsSNbzDGbZz0PSBBBsPuI0jOlvphOVdHb2zL
0xwR+kwK63P5FU6TiuNomeFmHpYJEN8Q7fnrLeDPna2qg60jGvFB7Lwb8puwYMgwC5JFfu7O+Rp4
DOrHQxsfrfG0VuNA/jBu1blHLvE1YxEt7r2mV234Co4E6gDVdw1wHyAkpCguRO1vBTuZbTcwwLnc
IZwaPI0frDpYX733Jduddbk/jLZuEzZNNLKrsfraE4s32hZ69QGBahqwlni2LiynSVr7Bb1UNwRs
B00zxz8htp+jALwOwtEKqM7k0CSSHoh3tHDAnyf5Km+tW4lrvsCXmmeVUSffO669r6QsrtP6gHT7
VTL/a70bm11oYwtFRbQAcoLyl5+Bamtns8/y89+WecQKriAb+2eaEFbAbfUMraiPLtGY6tts1nBu
Z/5Co61znpT0RqQN1DyYqR/M+5BGcTNrKEcnPQkeAE9GPIJ3mGIAAMKJs+j5NG8MvDsZc62sgm2m
nzlCPeqYGl/0jtyzMU0N0dP4TKMVUOToacqvH1476qKZaj8/lOFKVKAyR0y+31SW1pgYNfe5TPaI
G2IFUlOUwf0QjLkXmdPkYPp9mmXEVcK+E302cinH9OtYw7oRbOSzYHjxYei3uWLK60hBAbxXJ/Qh
P86ugJKrnWNCYFCrqv2YbcJKFi9OwXp5a4ky8iaZT52ssDRRznhNdlZY6oe9ra2gBq32mIzgSUbS
bhTgp/4miJG3p8817yM+Cz51jY6uorNzRaDk/Ad5UTxQ9FMZk/9/mZeNn0oo1LjKlIx1M08yMO8R
CjDaSJGQjH1pRCEjQwLNgQwjocwSRZQt7GNrY6FTfJuXlOTPsofusZ3KDLu5qGK4pW6zrANiP8eC
Dyua4Qh9xQ2gOps/cZgskVUTILPkFamQIBAOvUvpiP3vasAV2uJYwe8qpHAKAhdwANbW5NSR7SzY
we2IcCSjFC0fPSzvorJtsWzQgp+lgTUYupT/UZRt+iCkJgkZGflKFOLhf9hys3r09i3oD6euMq0e
5TND78Mc2TDKX/kRahjnGqKygKKCyDqCN3tb8wBx6erVIiA2ugv88gLB7CnlsG1dHsALzuyaI6UE
8klVGAJqIjY5sUiARy0bifr7pTTp4Lu8e2GsrfET8qvMNDjaCCR7TFqAnArTFNZZbQv6ixPyVoMV
9ODKfZDozzBnjK0FewPdfAEBhJvujMJO1A5tCWYSqnFgxBT5r0YDOEcNsjApjxZOluFx3Cmfiy4e
GqiFDU+5y9sMLz9fKq5T3SxhNnf3nV/z1TGxSe6moDRVfpLpJOCBTEFvADBxghsw8A8/VcARu2gX
tfWQWVMeDaqtHOqXI0KNUVlNWEt9PQ5U2SgDHQnVIosK8nwMynylvQtehKu69/l2fujH33ju9eDF
mMUQQgzKrP7UJmQAjz0bISqOsSewyaSOKojoa/0PEebcAn+DmpArH/s5RymTztGDQRZ1c44y3kZd
gsMLmTv9cX1bQ/rLnKPYwZjYjXZy1bd7AJwXqH5NaFeJebz9cgo5RnLZxY/Jod/qxlFYFC3CCbgY
GlNZUeTwOmaI1T428wex7UzSieYTMGI3qqEEiBeEBl8G8a2DnybvWdjc4nw3I7G0Z18Sgik5FRSE
+rGS9p+cTqyc5J9ZVja0tOM0C5+a7klZF135YsejhhjUxBg4RJsTgaN46+zcKdE1+oOC8BvCOEfu
2mvm/SlQuNHBpKEp3r74OmEfqWzHifFaskj9hWs0uhJKCTeip1Y2QTIyoHSKYMqbt7Vqm1OSm1U5
H4PzCoJlFQ6zWUaQbntqaiN/h4Y4+Wa7angMgh3vj5YAN16unuJPZqIs5Fqf8VOh/xIzpORq0W+l
1bwVU7vJTJXA+/ubvwDXfrSikKEUvx+/o6VZ9zsteqPJ8+JEw00z0w/RJMiqTT7Ss2B0lOVwK8So
u8cMTGwQVrBC6XBguvRJnet/9tP5vViG/h49aSC+mWKWHz9y/txC6ScJPVSk7d9XxEaD0VdXJ9+6
VWXFDEhajT6QLYmni+6H1+UUAjjK6S3Kd7ZkYmt+5A9HeqXSbzLloq7pVYbaB/sdhWE/5AstwJTQ
u+iySQ5eqJAdxhjQJUZxUhh/zfndaP5WE88tB8vzUDT3MOjudWxRelydUyp4eH8/peGghukgeE8x
iJ6HZzmeDyK+u/N//jMwvOuo16mGMpdVkKGoPslkJalBOnM/vVp15c0fYo2hWkZ9qaIbzmZ8Apxb
JhsrWqHML5YEff+NzLatu5HYrwkLkxgea4UfNqqcKjzc7Lzqvubdpw9kiMiZgbRpF3Y7SUFFYkU1
jkOzYF+oYQ/RYdb6/sdFMLSTm9Ii1Dh6EoFA9EZWSqjpdlDJ9uB+z6laMSeG9RlMjvwn4oKkG2ww
tNT7z88fhwttZRyQ30RtDoFF5/x641Da/dXkDn3AYgohNfDs++Y3aqRuotPPHGcfGU2wfZ+uEW1d
qwyAIWaNQVnNSBkoby6s2SX0C3giBSoEiBghWyMuS/29V5t0jtrMoffGeoBPEAOkK5Fqnm4bYMZb
rYyy9z4I1UZLJPibnmG6gBDfHkvGR7GeSy/zF+HgrgDSmG3PVMhhXtf1OSIAZBLa3/+a6A34aKfX
6Hkelrru59DrI03zLjfE94YU0lhWgxS5TuGLPQxGkIyIHr5ZrJKXAifwLDzlvc9lwMzC4nMQVU1l
PBt7MNub3EpGBOiBoCGdEYs1+msiowidO8esGEcN4q+exhr9KKHpyLdeEEKhzPYQhn3Pu2lxy+md
Rg98zoXZi/dWcLeH6rOEqUOXVHttm27wKjZ0SCJ/joy4c/4TFbKYh5tlYjgzldBIRfT9bT7tuoXD
kTbrBwLXmG624CIvpjuGYmROhKf4SaMxe83qwk7+wjeGc4GETrqfWbCMcHoc6h9h+EcKndzEOLH8
7RJmnWHzRejs/6KDNl15qc11vtShPmxsl0ZI49OF4hksNrnAzCtDbZI98kWZE2SX5GPICQjeRsow
ViMq+i2KQ3MYcgSLblCfy4Q5DgQl0x5X5OusPaxX9FrRd79c99wCJjHkbwFI1DXK9/GSJ4WPNkGo
EmvMozdsFhm6hm3IXXXcyahINsuLljKixJnA3c60VYAGVgwJiOQOYWDXxDLHgxRTX5Bk8K35Proh
sdyXcXShpGDt4Y0VP6VAg0OCzoPeHHG3uUWeyJQuHlbNcnXrzcgGhIVNNrCyGDY4ChL2kNM8IW2V
0+wyC3vRi4kIp94pHJU6Yh0YoYgCU50sN8zSdgp3HBAg0O0fkqUOXH4/CgWZ5yyXwNsqWMCszRML
QKe7+pqnVZXxR+UGfCwB+kfJq6iiJvb8TIevni95S67N5v+cXgjrEzQgC+BkQg3ch7Swr0oyJHPZ
Q2rzccVr6EQJimx/t+gNaGkxhewqOxvBBcvVnFt6kr4VIcDMgcTuUgB9pWRXE0lLBC+d9qkAOELS
rB883lch/8vshlojkYcXat3kQ+OyaOb3/v8K4DnvPho7n/mKvfcHnllIelTeBM9eDdihwuv8KIxe
OvjOVrArpnt5hITTypgHHS/8b/8NxSThjZj82GZlrixJx5gtvdRIJuhpSltiZQmL2eqmmCL9ghtb
kQGcibfSGsm3t0dc1X2X3OLDv3apvLqeGC1VS/JhBKSLtHorDFDJ2qlSNb7WasRQlT8O2HM2NUI3
ni3/yQzgwBnoM6/LN0LhFerL234CZwmX924Nh4xmKfae6ae7jP3o5R8kZXeq3GzR5x3WPVQu1Sc+
K2OXZb1jOv84E875+uaEn6IbRGvdG8VWc2TQxVn625poMBPC2Jc4JPIssei56VCbyWE88vVLrc3e
Xa6PGzGn5zTMT5rUmE3ifJn2Z4CXj9OdZ5pChzjXvdt8Dz0jCLJ3CU0DrhQohYmAXhvXgFaD8Irm
W6vEI3ivxWazFeiz2LOhFkPQLD2dhGZoy9k3o5WFlX7K0WZ8AxLWd1vp0Y+tM3D/ZMmyLoHZf3gj
zbbgIHnpmdhWwcc9mmgzaaKOmOdSDk+gcYR8geuqwUhWRKjfUa1067pxzupNigDfkeh4nruf7YTR
Nk+uY3Ld3KlEV1R/CJ5gmLu3dGksNpElF0xFPfDQfqZAFAbJzREr9QAzPhOb8IvJalBV1Ql2RkqG
KFF7kfrQedmgtYvuPZV2NCpP25oJrgyVnHY83Ud/a3rh5hvOP3uoKt/3zSy1qVV5Gi/xSiwCvInu
5q6jkpxPFdockT85IQxZm8kmaGDMuNrlU5dx+MOY99KL2phELB2be+vLFKGiJMTSt+uwLID21cxN
fuGNnA/fXuItI6BpbSl2M8cvmUCqo7CouWR0SSKlX46a+1DMxo2aH4L5kwf0t+XmcH8BlTWFHo0G
Mb0y1EfIirqqxMkysKSTqN3ThCaHXaz/O65Q2j424gTwv9M97E2qBi0eJmVJ4CwsZeVwexZtw2Sh
SmJnlglNZgrGAoZREKvronkOEdMX/GH3PWGuWl6WbIAwgeqauq+v6OH1mPsHSSsSFw4+J0z7eM3U
dR/8b8SaQVXDM+j6qxSVNjCrDrgvaYQocDXsjyp6V6TVgQMK8SU7oxrePh9vVhMl8LBlItLvDQXO
XQtJBE7BS+5MIbIz4iXvsbwgPQ31dC2zD0tWoKCzwyZM2t8IjJ+wu5k8GK89dJqpIJwlipfB14jb
hvOrNEJWQma9p2wG4sYSPLTdNQ3yXHVNrlRLbrnIt76oLwddEYAItGdEkwsKejH6siVwFnHoAcHF
/iVI6GQiqb+ttZzVpeLV4FG04NTNbTfoQCCVHw0FZR65G0N9gvLVOnZiGuwxNsTl2LSsB6FMMjFR
dWNhkcOwpJkILZPrA5GQHWeXpSlpHYEachqddyitpDdNii9Srhpl8M/Ew948wWjwjd3z8OpcB0dL
pEQ91hx4o8AehOz/USNq6hqq5jpKaVFO0tWgwvJUo5eR9sRjFXyuxGR1CZAp2aotmbZeDmPqfBiQ
iF4v5tkWM0HllBbSvICpsbQNS2abxKVeh8XwRniEjCl/0XPRHn8xSFDqWbYmgXBA3wSRGmkzQlfC
AqWg1tKPq7R2OcwlrexsMi/Ga5T9ARbPmkKpf9Fz0Ke8PlxAUBbBdgnug/n4qpdRn6FguDssS4f6
78hEppuYWvcsSRiEHPyVyg7sAAVf3gDjbKvet2L3mB8fGr6IeXzqRTR82ZKxtpMY9cRYgd1B8bJc
SC5eiewhs7Dd4umbBi9wx2MEs8RD6qfkM4d3Q9SqmIn1wr2BvV4wWv4vTZhCSU+cdrn3q7VnyYMq
mk/lWsCbHj5c1F/YOfxf0eiFxbYGQrcVTI1hwi3c7kMm4Zyl7FcR58Z0QvTtXRaB6TGiwqP+CrwM
wg9PoiiDtSl598XivxjkF5GsuhgiIkBXQg1m8yx3dIX98HtVKipV/81EMaIZh5V7QqipWF5YH47O
FAqUGuw2MO1LsMimT4zpzKLIkaewNqHr8lWc9DreN75fHTLMZ2iGc4Ft4QYiQK6qwk/6CV7wZBfd
wSL0fg8gPq45HPaZH2rKPj5wi1ooGpZAoQ4x2KP8gsHcJmxhkNgi9SnFZf/oqPLJa5qrsI2L5mKL
3dpQfKFZwIfnPEDsQO0AYxpFRWwf5GJ5ibEs/lIeWYRi5s0m5bh7o32HWFi1gz1XGRzOJND5uACr
OBd0SG5KYRNVVrqy46UqSPYSr90gjkhmYWIxdwmB3OO8MghK+3Lvb+5Ij7quRKeIJO5R6EChPIpD
rYSV+glELx1AMLNh3s1kEYlMjI2ELJu1jNM5iMTwDqQ8j8Pw077eNI8k6bAkMqI0CngnLrb7hM9b
axkVe4hbPY/floh7teGSsJaH57WmDVeU2sNUpDAWrkOMdtnNuAxvYtr0m22WnbLYAZTbrb7soeH5
KYGo5v3mp4Nef+43o32o9S5F8WNVG4UtWbVYoG5DAwCpcqea9DxPtRKCKrr3HrNgZ8fN29KP8AvT
rFAbYiZKSybUNXPX6r5/PW1XSzCaQn7Hr2TDJp4ns61uul1FUH9UKiDl/bcoZNwikY7YOBuL6fYJ
O585zW10MX66msV11iqoRrgDHy3hC5187kxLni6czhfw4sR4iOwEymTo0q6g71txSnQZSjl+Nu+7
3aK5MkxHwE1VTP3i/I6JCz7ceheE8dgZ5iKfA3hC8nucofqzJ+MyMf79567x8ugLySVRHOfcqN5j
/gh5fREfpfQuTmG5YyJHo9TaS307IrxszDzTVSmjZa1FvM/aFg8RTuT8wxGUnmz3/q50Kij/pvCR
tvuWB9FR7W0kciFrMvHGVq2+mlpiackgRMybgyp3QTlnMASlfaHTmY5iale+QMVX4xuj7LWUt90Y
Ed7FVzZTYKg7fi3oP1KZZoIVGf56vdz4RgCs9yZy1iGjwuKPOgBR0ZuuZbN5713q05zKXlguLM+O
WkkmtyXI70mFsjpWLH2ZW4lVqb5uQzufavOllwSyOm16F99vePPWtWyUZNtMwwiRhPOq4q/qDNcb
GMdmOyJUh+pYwcsUhsVxjy5U7LKE9Ed/HtjXjyH0wU29XmfXbKNylUS+CjTA+37zXVw0JEfUlGjW
pwyp9HoqjFJz/y6wSNl046jyoSk0Qc95UTovaOWa0QPhTelHa60+g4aP3ZzgbkFdb8Ea2KBMJBnk
wRkyBvElD7f1YiiSmKD0X1WGWRPAPsYaAKgEGrdk3LE6G7anNCGUx+FU/n5sm77jTvoqmQkeSup+
tTq+fRBU6q3o0s6b3Da4DB0bd7s4q/xcE0BLVCu0g9UsB0tE7FRUpon+qTpu+YdssG+FMJgQHzYZ
yA4nFPwQLPeOoKGEHeOYKbeWGpjhnM+NnDn3HGWs6SaEgRYqLT5Efwst1L3pNFCFuESaXkuoD8c3
wd+61qh1ZNcsw//oKK2+u7ieCvFljcU2Mt4OeD8jomJQ7VsxjIH2vqf0DNLdnkvRsLd9FvfqMB5V
XhZRWyK+fbg47TMZqtAx/qSpdQXuZfarEbXwtXcPhkds1EZJMsDSvCuGhNVdpEz5t1dzl2TBkKYf
4WDoVAC/J80B4NVcPWIPQCqZFpnc1zeUKrb2VqfHudCtWagAga889auooFJ5NXgDD/uhZQ4JSkqN
XdqywxxTM0ab29iDzwH7/wha4Ze51qdl6KqdwdQ4Z9WERWnwf4c18krzfYm5wbWPFvupNSPPfOFN
cf4wSqRKmH0W00Bgw76VG+vZPtf1lo1iVSqZtwvJQ48ZOU/HCUQNJwboE+xXK75MY3tRda5ZvIsv
gonyt45Ba3gFv3v6q48CzIeI5ZXfO8teGQ5Ox3qYJo1oQ1RrTcyrsPrXAvWa48j3Bo206w3AHiMV
H9qlUelaoWmdxh5ghGDb10lwU8NFYzEccB3Z8J5L7jkCwfPXtfo+EpKAOJQ5dXIQqSjCDXABsHbU
M3UCsjptkpV+gSqcaRT/765ySTxPT1z5TFOPwfjI/nRrSyqADrtvNMJSSadkAn1q7c5Qjkw9sRhB
fx3wEZKMy72dfnnVJd7FNqn6dtHKdy+RRWCPPDrTN++WdNWjRgH/iUrZF4pbD61RI75kTdO0uuxv
H/AciIZtW6pbAl94cGRpon13uxox1X9mrl9GMoKBtgBHhYQbHFmIaKfS6qtRYjaWBBBz6tRpbiii
x7ytwKDlDcSMpYOvQUcJd9dh4F2oxTRKlI+QO6s11nVF+jN0BMPd+xdlyAfOFTwpzeEuuzfKo2Qj
kgp9YmYD+fZK+P/s3ylzA716sy5BhuiWhMWHL3Tul+O+PSpq+Xmew0YOjXgPwHEv3KA05idxIJ6Z
5tUc/i9FukBsRPUL/QoQpHf67Nf3BtlNn4ltCG8WRSOQXZ+Rl1n0C4meLLif+gw1QG9qlqIjwpvT
wNINOPpkH++iYFMLmuWsE6visc0UhuVLo+ge3zlb7tZHZhvA7S42IABrKrsnbcu7IcLYuwj+U2ZE
Zy4myajNQvTglxRe7pP8Cblcs0cBmT6/2NywRG+RZHv1WWE3u2ZNjLRJdhI+RUjXdU0N8j5vlxyn
B9lNb0WVYNPqpTEy7w9zNWOHLZ6ZavOrt8gxgca42DWBFve7wyjk39LJ6/YEcpGPfAdvwkrvHe6+
G4krtI4LQs8CEukHs5NOymtsfaGONfkRChAZV6/9z40BwbYORw2APkIBlCtTv+wxrpR3R7hebaq6
UBjSmYxix44VMynwV9m+dKB72sUehUIe/IeETd+TL3Sm3Cr8YrbqOzapwMC6hTAD/R+RTeoQB82S
Md6FHSzqCiWELW6P/NdXt/C01qeyjyD4HLVJaEJhoAN0PCgSXb+al+EUC2xOZ2wRaUgvGYPyOhxh
RuKsPSpWodhXyFAbMHfhFTFzHnGPMTIDKVsxg/CE5iNsNnnBn1WpHeWkzfmkRxRHf6cK0twsqs1Y
OkdyUDjF6tcr7lYLetdzexOL/7MDUUnfIDCn9wPa+0LwxHIgg6QArwaEgecDGYcTHjI0Q6P7MdYx
bCm+j1Nz3NheQSFUYodukpfYODrQzwUOaYgk/NFcLUwcID8ZN6gq0S46A75JWiJ3ZH7BSblm5NMZ
AFgiAn6HIIqBFSuiILoeMS3jTGDCsmCDtJlhguzSNdPjKb5Xa0wKV98wwkgY4xyPPDRdWRh/x2a0
TrsceQ0G6RcV3OWA9OtEkknUhk8Hq+GAwoDCU9wrJg35cY6bC4x+03xkdTuDOIvynZQOHtYKubYI
zI6/3BSoqcRvfCXexHJeeIQncPhtQEtp65GLB3XaIXU3bbjjVNJa+AxnPG8epyNbyv87LJo2ulb+
Uv+deefv1DWJt2dRDJsdyrWPAocxDu8TrE4R/VRyV+l5SBCnnERZfKvtlUMoiqyT/sEg0KUyY4Hy
+kurHVbu2/zCUhM9lSpb3XQ+u45Pr7byzWyo359CgCX8Xy84ybelZSBjVbq39TCnkeHOa7RCSyvL
9nPYTOjzJbtaWWjLnbwMDdSvp/GC3yzW22hW/lz+IYlYPe4hjkkhQeJmBwwKEzbYxH1wb7+qmaA2
d8hV13Co0RdVfRXR/fTF/f6PtqeerQd72ePKTv70W8AdyQTWcBhZ05YSefwt6WNfegUM/qjX+b2v
cnoLdfLK/pQZkkWUmE19emjSv2ZoQRxHQK4HeKdvH+4qCMxYQdIw/lrWj1lcw3lccPOj6cgCNwde
lT3L0Ru6QX6H1hgu1rlwRNOyc4Mja7jtUqe5pb1rfOKkee5ISoW0F1yqdxSqNBNFEftgXL88zqIJ
TiC9qPOjulwcjhm3kPq/5ayUJJhOejqII+zreVkP6H3zoj5nKerOQXvDtnZnqQy2ze9EQnWw6QEd
bEsphyZSEHIWsqlaFtFIwfa9wQ9W0tlJ5WcQF+oIidmkioRXKJP5iLipRjRNVZy1OJMuP4RmNDyh
RQ8x9m7axXW+hk2TmX18s+Ved4Ig+jTwwxV7s6EGJqMJPbGWYQhDlnU4cvMJ/HI1dxGQLSqesqp8
Sstf9O5tm5cyb8DIdQlyA8VrB0TbOi1O1HPw9wna7UrJqa03OdX0q2n92RPwYVv3l70TLjSkWf/7
Umo70+NW8XSYfawq6Ta9ccCZImCrj3Gk1u+J5f8feuQpye/vZ8hEabhGwopLciFO+5NIZXFurY/Z
HG+SnkncL2cjEwznTiPesx/b/to8mhgHaBuPonxO6PRUmK+u4S6/3NRX8BAGI7FTtZFLSIdywXN5
aI6wUPvItQFPF5UexziuhmvlohsfRNwEftogbHhO3OSQN9sAZhJh5tvbjOA5V41Fwqa+8erRikmW
uAuvJrk2SV7oXXI6NAeoRqtucAWyaEcziJbKIrmmD4f3+4swcCBJU8pvbXnxlx/jMSumGS9n464Y
G3zOdi7KBszWIq85xkKhbG2QfSW7+HcQ4N3S+JtRKF1dISu0IXtfTS9Dh3fwf39v10vtpd3yhEmh
DbKQaCNt9NlxjA4WQoUe+o1Jgn5GxaZPCvSWyCcMq4t8RPfPq1HC+KcmM5WXesnZLYsyJt9WZy/8
UHD7QypT+uYVuHu3oMScHd7uUaIZeagz3vvE7/XMzy3l1JWmVTdJ41MpBvFSk0U0fGjyHw1Mucif
hV1FmhCV3JyktQ1hQMTYvcJ1sTqeBYhGgWrw3nsb5xyJeTOEZLkWi1pH90gm9ERItDVXPtsXss7A
a2ky/VxGtvYFkAWiM0txMoUTITiQi3Za87YHgh0pjc5Hd1B+IJxW6dmpyyG0apoPT4OuftswJmmP
9f6VupCtwNuv2iwht6sIDjcQsbC88zO/DCHvlyKjmwf27VmNXrnoeEHaoZhj44vczB34N9yBP8h9
XQvcAxGMDMIjPcLguOTf/dye/FVGMjdT8/0HVaO5yLwX1jw9kLhtav5coCWLAG1/0Wy3IXT+XhWJ
ylfrgvP4CL9NCUn3rrX4VHR8LjQM+2kO6sMaZ04ITrsUgvUpt6IZZMn2NspasvFMZaUSaXwjGB9j
3FShadvGQuQoy4yM0eyVTKvWGDTFB6zRhGiqpgy9UHgCyqwwTzhW2jqFVaTRlrkIEi6DbAN0pTRQ
GDM+THRiVesDTy4KI0SqN1zQF6y9uhxv0JMJNhh2b9MfYk/nlmxU74FlXq7zf2LxCFkOcnjjJDcY
nMUPTreDLKIAQohUT2mJL3pU7GRh/VDD6s60ZTba7JGqffvXQFiO5XSD5P27x8CRwBRSoUedOmiN
VBeGyaDAdfThsYIaia0uvHgp/ULTPwHnHDGeoszlMbWSRZXQ0qcfqHVH09oknbiolVatNjhM4MZG
YOrStUArR4lVWWQvbmJ69q8FqYmd9dLgejZBaBCeX4afNUX8FI6I5yyQn/dO3bS5qK+8eScQAnQX
Lna/5SfjHr6bLSntrZXV4LIlTuqXgr/we820zohJm3/saMbs3GCxO87BHNRaO5FVloQmY7kk4HMT
ZLO5O9dQ6kkmdrEcriks3yOo4cvmou6KDijVOaRDLbsLlrHin/X0hWEfCl6gmmrrUNTeb2HxBksp
EZUw83WI6VASlr9k3oAdLNGqLqY2Bly/KKlwAmnqNNPLAPoDPFzU/Ztn9pG9sZ0/QxDJS+MUhq+6
Yic63eDp4KvWnABt31weV6GRfxyGNJ1Im4N3MtVrV1o9hhrUmCXR0Tl6vq0xE0nKbX1oMjBtlqbv
gjGuYdL1rCw0kwsaWzZCtBJHLsbqWcmDZL045VzAER8zOeWGhVAePr4GwIfnOE3ffb/MwCygH5Kc
auqtdAkG8I6/aYYKjRH31mDuX5r82IgU63R7V+3T4tUquVMWfguhxppviWKXZE+viuFRRUaNQv5I
o4SwnT6MVqCj8jL69XS+hLikQSFQAcPkLVhVvkVOotspQknCEw1brfxPxyPjs/i8mgkc9Bm9EE2J
hbQJOYjLtewBZm5HkR1Is5dOZJ1TYJZZpaN5DQ3LA2+O5t6MDtgRufnZyC9ZxZJSRLBeAVkzIvDH
YmG/ymd/lTrTO8PSXYE7SOBwfcQ7mwmNREYgsbeIyRsz9w3IKNb2kk8Isl/NljG71XdSl1o7sKAD
x7LXRmVGtAcqX11lrnWOUzhFEWOBiTLazecMaAzlxqLsrZafN+M2/s3sUDlsZicwSEObJYst9XGd
ynm1y0Hsop8RWWxtVFq5c6oehpaI/GvMHZ6vYx9pWweClmB0Zj6J3Wozd/Yy3XYjMh3Kc0ipWoXh
ucld97sW8AdUwOloep2L/W84i2Cv4fVgu6qPXGlO13W0a7h0pLT9GMZmweFBTKmyRhk1yPhaEhMJ
AcxpoxtqwgleHRz1cnD9/0djME/zCSridTA9F9wEm5VJMxtCG6yIj64u+T6iB/wtLvyN/GgD+PaY
0RdRJxlQIgktesg4fihZVkZc/ca7mVuplUyobt8z3Oa0UcG/XB2z54aGrv/oB0Wqk3B19//lHKh7
6tAmq7QY519eBgkikBD0LqYhwxn/hDxF4cmiJKmYSvxGDppp7kJZh4+NAlb2O5MQ6Sm3PmNxuTb7
ZnSQtmgfmIv7SMTqN2S2TESDFbwqb9xx3YCezzl/d35NahdB5QHkAt9uq3UJrzypvj7gZDDgilnD
vWsUcMSHznv8C+90/nmabIBdH43aQL5Hl2dzjAuR/kAybqOQDSI5+QJb4ulN0knIiO3pQQrmFoB2
lMfY8C40EEie8ITt0OCuvUWEv6mmLoYAxTgF9Ybys5DauRTI22qvaFvDxmylbrnlbULjcEVAw2sy
0aWc2+56MKkaGEboQ2ebXC7094Yq9G/Qi9l3T++oQR18p2D/IelZnEfqZBo1ZvTPx+EV+OwFuA9+
sTI/lurs9VrGrIoEslWCKLYMb+EF0rC7feIoTCU/rn9zhXp7BN78Gcg1PPjkvRzUZdGsyGmseJz5
Nl9qPP9N4UryZyCrd32N4TFFhfcGR5nFvoqDabu0le6ez5w0CNzy/nR/rt2fR+u4BjmPLibrRSRs
LGoEaI0p/VFhfGzsHvC5INLKBHAAtqhZxzmW4rVZziJJu/p6xeRY6v24n3PSBoxoR56WGdUGxO6a
aT/OgYNdQzYsNwyeWi/OG5+THjrs7HvTN9GxUDpzxozqlNJSDEXWS/UBlMPvYXYxc0+upBOF1c4N
UGfnsczBKFqpO1Rvn/76OeDP3o3ZXp0s4NXWLt37EgDRBTxGMBiOBvfBHI6ir1sm1WRuzW7LHMW2
3jaONYDeeK02H+l9Djv4XwXHQHIT4EwIlsDiIfb+CqC8wnZfrgfD7BQEeOFhamw2zxwDJiI+8UUX
4yG+Io7GS87o6KhweYpiyWEPZaaiwNg1y5vLVi7aS6VeGzdlsfN0ms5pGHz3e+O2h590gwSuk2Ly
vHkollcwOVHRCN359z7ExbrL2fl1U2E6xeXiVB+iWFSMVV9wrFn9MvxMKJ5ZvdLRfrFvhgoHEujL
+sdHs9DTSR/sFaul2xG+9R7qCdJkm6mokyiP+kgIpCW5fTCaVczHkC9i1zoerUqEIEGccLHk/pEs
v8zg5hwiMeF2VTV8p/x+9fjghNX0cNh9hxJqFJuKuERcoEgW1339mY/ubC3VB7ZZoEToqMSvF/W4
XvHev6VHb9vvxrNuEeIHSnl9lbpuPArTWNfmu9ysgvbkgE+A1/oImvblAmoE2mNUhAYz3jUEbpft
0Vv4DKmCmY2vL98af344W72/9Vnx03Cb32ohlVEejgDomXbE00Odwq+rYgu7dRyau3EpOHzEHY6S
frX9xy8Bxu7v/xP21A7buBbQSW5umFa3uaQWBR72p6VXr4gNEBb1thgbgZMdSWYzXoyrteCtmZDf
1gh02GRwRpQCj4Q4nBgUj0fIZy9umOeEqf2X2GfERA/MjFKCFiHaCIG7hMZV2Jo6uX8KtXMtduhS
g9gAN5f+0GpIsXkNDEjckqoNbqwN7/bR7JLsxEL4phMoH5cdE70rHpxBSOKttb/5c5gwEbKZSvm3
C/G0YqI+Lqhsn7leW+q6Wsmykw3GfdsotDcQZpBH5jNaNSifNqWj0ZjUnMtWB8u8c5JCU+jZqsuF
HKwdpxgRolCKTBxTmkDfz/+1k2rgIi+lrx3sdfd6Ubb83t2qHevS2cGfuNU7loWwPF+NsJ11UbH9
h5idftcd9aAvy903Ll+J0JutF3mu+SyXPmZirCHY5fTiTvaRC1gAwRq0d0lMG6/WLSb9QbwG9Y79
rUXcm7Q8krojUGHxf6CbOMlXuJQVh839qDD9uxc/j2FypPHe/kCqHx6dmWv3BoP53oKqEtJ/ounW
4WgG3J3FNOHMmBODrKcTUxcaEVIUl5yrSiYu0SGsYXr0LqglTDN1TGR2yvMFwhT39Gv+TMB5aZ7E
dPvgX8sL8o4swqYSdxzLWt/wT7cbph+iV1Lm6idz8F5fThCBMS1ldl5SRDejQLbjyHSmm0pwE4Xp
Mh28riNpBFyCs4wZDztsXQHK+jNMODOp5ZwWIQjh5XUK3dKK4ksRShzeXaTM0eZXbh3bAE+LAPZE
uiH34IPlMxQzU31g8AhMSn78vql5h14WdF4g0cChc4z7JjLXDerQqeSJOE4qjZI0JlIo0kQTgH37
Xor5Jus22X2m2ZNkB4c+MUTHBcqV/VRAKZaGBgPFBwR3mDyc+wQzRuacmqqXmkpH5MyGiOzX8Nfd
B63gfP1l4axlNnHcAm+0+MJPWDePbOsytOLMUVru/mqV62IMw3n4w5vjdOlyBJillCWrHAJDWsIl
mzPshYEWyoRhj6eZ5LFwTtgW3UWmjS2DaPr/vMPBSzqPgmuvfPfgcrSvaQCrTyHYRiM2Cs1qdMF0
mbV+B2EkIJMUy72GEo2N8TPefBfFl0knUXf9utgN/KZdQBTQh7t9SLhOFlaPhc3vHaOdA42y4b6/
GfCSDpwmQSbLLE+g2Ek3aMUlTsYMPFc8LNi76xX2JJTUJ3W9eqaN/NbkfbPS0oCjvtlXq1O0GEhY
PFQB/U1MFk1xX8CMOXkiyEme8WkrL2oF6IlHuKI5yWevaBkGfpiFa1D2fv0PoyVgQbTHyu0xd0+d
ljDrb2UqrmSaS3CMlq996Aqm50/SNMQ3l/51A9jMnKeY3TIv2iriz1YcTN0i2x2Dce3/fdadWYBo
UFcBQlYpr001uVKblfTPAsWmwB1GB29m3sjqY7C7BUr265xcl4hJGGKrEED1hO4IrcpEHnZhCfng
VrLUHk+j9SIrmsIUnYKLyplOwRnPw9AzVd8hp0LM1K0GD/yVsYGzS2IAAELZcqUwIwJ1rD042QQ0
I5zQxnscwQfuEahvs/Djdrrp0VA9PTe1yzSa/jQjFKg89Q7NV2iknPWyxmT1Wb/AB6cTOoo1y0d9
CShgs+1NDaKc8oRfgL//dD3vr1nmE5jLE2tLNUuFXrLszBTUJU6FF+CjjgRi5ntFTU5VsuPjGThS
bgJvZ5vU3vfxxD0eB+goq0YuRKpNN1YVyTxZ1w/SN6T1+ylcgeHtPOYufYVGTd6rV7Kn9bibD1tI
QYCZ+uUA++JdsK5/M7bXBOdXYSXq/BAzyV1wmiL2IyrtaL6pzc0ZzDUatKkrghEtuh/y+x/wuw8+
i7XCTEFApnkDX/D7I8fw5eA62DSpIVJ4K8mkoadjde0r6zOuPXEDNizVI4KaXoBb742s0OO4cH09
7d/WIHbyioRs1fXfH3qn1jFfkdFg6CJSnn20d0REw4x9MxBkmU5Cuk1YKvEYfogNNs1xWvt8S9//
eLuRtacMQ+YL3f17qqwfsbfsRFTRr5SbsBJESJQ2NkHFytO1NMpUPL1/0TPAmjx5mzHMGcqhG/UA
KR1AswiMPPSGovLJLXJ+SD4ZUXrD+VNAit9qG56f3WVuwsgm+QL7DFZ1tYN0mIoqCwNY/LpcQ2QA
EhhJcHWU9vZloiM9FWVhuFydmZ8ZEeWRXT8LvlvxiOKwGp3ieGZyEqmqIl77BEPIruFm8lhgS1dt
9sAH9BMX4GnekeuM/Ft3gX9MKTKbY+xlMkhHeJkKd/IZ4eoncA19Zsy74kS+TMJSCCj7yTESYzr0
wbhCRW+K7psnv5EzoRCMJf7ALPWvMTc9ulTY/TDNuoFb7A6rdyf8fSmmlgGn7eovW4etIONqFkhv
x11+ncMuJLtgTmrow5WzqU0xpbMEcgcQSXOm35GIzZFOiwxc/8nYFYhRi1vwsIFiz4ms8ExqcsLZ
AwuqX7jYQo0f8qLopvXCPU58vZlo9GG44WNebcI2ApA282hGmM2Ha+/OhaOdA+4ZD7QoNQ1eOyKB
1mLybuY7KilSqGSsOetne4QVXJrlWk3RwCwBM8JnF6caYMc5R77rgwigV2hCyv4/b1ZARrdMTAdn
N6JKCZ0HhJhFaAq8aUp9n+SfetThJrpyPw5bsojdKKMpVhMHfuq2k0p6aqAAQ2uBZLKaiQa3jG/d
Kt8LrIfODm3UrVuu4XA/yAXzxoVbKMgcFlBvHecxvBKGX97EFB1/lUzCHmGPFIRx6nM3XeQXImSb
OBL0q8cpZi5vhWdZruncWnDSZJxJqAAohCjUS1XZ/NSgESFA3Po7anSQ2nQmJlR1+jRghWOdYIsT
ul9rrUMSoDTiVrjNjUdebXd7fhVsmqaONAiBe6uLfiJhF+Va96LvfRkaE5JluD8OrB/fFfkVFRvC
ihSWa9DeAv+psLAE/o/mXOZNdVTq7FN54CS0bB9WDEihsDHjj2LqIWLFdjZkVNxIyGikfPwgmZOJ
GDEwEFcdxEogLpXPzciezefk2hQjM10Ng7w4735mVvqzL3kA5tpnMMyc3Y3AwPsirX/FjPIdL8+L
DavEhybu0S7Qm3gX4v0Vllu7MCLJJ3qy+MUQx4yExYotEzoRlem3KK0uPvuVlMLEc8DmC098mZdo
v0Ohbnpnf01nvXXLID/ik/Jw5Tv0GR4Tku+70w5RLsnwNdc1h/GDommQLRcJaSyeSf1lHqSYZKc6
kwa7G0bvAM3ag+TGEpeREIWdU87dRn4HVE45WlAa+OMRCtsfTuPR4U7MJydVt7J8k7sHkLMKm9NS
sV6Ygqvgm+zT84VllZiup4HompnC7zVahfVrNMapOKkx6/ZrkH2ndiDi4sytFJ34LHbtDXyessG4
2DtdpviFO0KYlxnF3YsLhd3SrMnJ6twnvOhtWgewg2yeTf4I8+xDdg+bEf0Wv6UUKgF9YkOA4FFW
9SenedxopsTDyhyr/wjIkmu+LgkLomnz+2g89hdbICzfjGT7Q8oOS1x5MKojtnPpU0Vw1xZ04cIY
WboQtjp56ZYPBe9ZI0fzWbNMe3IN8b0Ju5ryk8aPOCCV3jYgB/1hgBAx6JmdotsQKf9t50IuZiu8
yaa9pGmkcOMi0SYZZc28jTmUy2NaZKInn8SOrZNGGTWf4b+jA8HkVIRUIZDzLrbHJHIRkIKeGC4O
geVPosY/L1mk93ZyWl7N815DbiitGP0xrbbala2hhzGmABC5n6BCOt8PXB2cH2Q36rchDCpusX/x
UAxwCdiv2wc2WHLtBL8xS//Ro+/mGnxHPz1XQ11mV2OWrR1+gaiMLDOPIiM6IKQKaQ8b09pW3Fvo
L3c5Vcdhs1hZy0vVV0MI8FesRmr/EXJivC06OwqK+wO8gWXqWR3xo6imoiITjdjSod2R/fbTQidD
LNCCwySlOFGYLcigaoJHxUHMyhLAriBRme4UJ+kg9Qra+/es4cXD1bjjOW1W64RHQeyRcYgz4Do+
kt2a3YfAS6J0Yyd43MjcO25mnoXwKXZ3V9jSchuNkQzQf/5ARxLR4ubSa4LukD2sh7JW9ZT8DkvY
WsV+ks8U1zCVp4k8KNu+KNm2v/WK2NuCyOXmVwTAD04IwHQGKgeLQU7YLuOufsmsxjNT3qmARtuz
b1pwXS7wFf4j0Jag2lca2gyf4+5qJ80fi/nmUzoCAoffXKlikL0QCEIIFLTSv5E2jcYtisG7ChCz
oUkyozrwGIhwKeySkdnfnFhUEHAIf5n1wG0jdmUQM7T/r1OU98ter7RDmUGCruI7QTA69xY8nwHx
pYidSQqGsY75zzLlUdIwf8W6fdC0C3e/vQsUNd45glnL+SxoCEimQWQANdVIpNM9KKmp8XkxVLtq
WHH0jU5rDgUzXjXf8DZMMxzat9cQMqKq/2s+uCHi35bFxaM8klDkASSZhiVfoDIlwDsWIUzJtei6
y4iG87BX/hNVbwcaTAQoFpl213tz5X3Zq2oEObkN0bvtGs789LQ8deWl2T0KBq2FtagPJB9UtNoO
F+sqO9uidP98lKxYOAOo1O5AEExSy6t2ANftRuOg1Z2P0FraWhHh8mHJE+DdIBTP7/RQfJuO5VlZ
L/jblNyVvLuzyFOQiLYXG2stIqMQ/5ZQoGrOMovx0TkYJFO1KcQhes2U82kc2Pla1XRFX3dyGcqZ
7k6+8a8pz6p6hdmVXOKbZx74zSF4JjJZnerSqnqGUGgPpUw3sMnuUQtFWtOh1G8V1NufZgD1hL88
q2dKGFxuTkmmJjtjw1t10D38mPpmRB/GAEH2916clZBZMuX9+iUbclBkbtaztv1hLv1jqia0NHDM
iU6KOICSeuNU3L31ZCVvnfpFqk128deUnqzLMc2K/mJ+oINjKc4QlVBqOCeGUzLIZptQWi6ikLIu
QxCq4SRVGZuagmgAePRNeLcU4bPuJZHPr0tESIkk1nT0WUF9GLvhOuzvTaqHOFPMOX86ZfWpcrMB
uikJcniRtqhIbVp3KOXn0oCMz/iYeWxTj0ZAAkSk76S59hL+n9yI+KZ09GE85N1mOMyS4lIW4aPe
mpk3cel5b2HjZLwKEMSSskkg9EHFeIJX9MHSAAmp02M54sw8jnpAf8zCaKu52PiPL5cjRGUj2J87
9TPDTyxczck9ku3CMlIwWhyqQame9FwEnJgn8ZegG1cqlD9GSonfUGV+N1b815QTVLCVSRXypGXD
dF+DU5lmzzCWok7jP3DyPgt60RXSNkCUaNqIVqyqnH5U21ME9ETDCQGmCjlr7BolGAALhjuI5TWF
VTlBqdx8HcoS1XX9bHoWO5L5H15TjItnR7q2c2NBQhh/x0OGMpMi3UDZD0jr2tNn+JhIkv+VV5Go
HdARcaZCJ8HrLxob4krVNvz+O6745a+WFPBgzMrwN2hDfklXWMJpPUv2F5LO+DihrPYfBVFeoi1l
UKrBniqp7mo+OkB3WNwX2nfOgydqUE1gLfFh5xCbdrYCyGNZZzNSSgeyXWA0x/aeHCAvsvYVCXDf
6oC36TT8Y15+WsGQxM6Ufxl4JMN4FVUk+nxPKqEQvhCOUI0VOLZ45UPUbb+4Ay0dTKtlhGOk3XbS
UP7j9fkn2CdYEulZMpfwh7+d3IyvpdcNFCFTOz2KvD4ouifNKHhG6T/6DlqJ1wb5ZP+SLyjLGOba
HpuOcyHQGyshDUPGVs7/6lDt5/nmYOk4NAKsmevlg2wl8xte0LQSIzdpZLHxteXPpU645uUSyI16
J0Y+HlOtOa1j1whjPhNyCNh3XeMJKJ4wdUIzX6keS7dKdfT0OUZ/cb3aWqnTqVKQ/RFgZm/IzJzA
ZGnrRJYFl2+y1GdX7ag96iboYOk4VuRFH2vx6HJzkE5521jecg4bThAndah4qRJAAgd2zxfTfKAJ
kBdoIC1t8uAMbdIu36rd64+S/MsvPIU5vTSTD6gXwcCG/I1EonUL/uU1cWHtH/qfq4nD5k0QH66I
y9X88tUmbVguKP5uE5qsV0E11UfOQ2Hkz8HDpP1UhXfAc7ymUSBQVWXiayR+DZGWxIW1gRxMyKKn
jAsw1ru7T2u/h8h3wwoqfE8X53D8vjUBoQcQ0gJinfOeT/tPaahQkTAktjIvjFsVWsFrT/thJVgv
NHN/boXAJo2MWIC209gd4O3zbXiAI0m9eVd5MK7grLPuGogUUUU9S/ekjXyZr9hg8ofuzwgPxfdw
MW/Rgy3WcscQRT00Bp84DyIl8DRyySjmZEn68/aYFk7E9Lwo+GHmcLlgoZ/SQli/D+Vi+gCcTo4s
GH/XeKpKQUeRGAVSgdwKqBnbAYsfFLWT8/Pl0wUTnyl6LBBIH8RqcUa2ClYSbaAkNSjO5kDLbVjW
L1n7ai1itf7gC0eF+bO70aowDSTz+BqN/9DVqMcdYe1tTbkfsN9uNcK/EQV9KZzuEfmeLOccdzvb
pI5jmJeKNMg/oRG3c2fvn3Hf326g8I+hekSdh+qEUIZdcEu6oZ6GZd1JZBHjRx9eU79GFghS9/EM
bKeDpfxRMaCxIYAhGeWLbqqXvDNyqxb7DYWHE0smakUMzFMFkEMhNMKEDhbtuK6KwuuqL9YizLrJ
PGLDuzZk/cSP38p+hGRzVwKf0Rd/ugAbSbG2NCwodqpDXXBOcYizDffS2Ab63BLlXvYD0hdUn82J
sodlVZSaZ1AUY0dABOMcUe+fhWQFQ9mxc97DHWJfUvs8LUbEc7GUo00I17IoCfJ4E0n8J8E6GMjZ
dTWLWudcpWsphblFyz6KJVebgS/pxcPNqxtFtD/WETFdlQ/ImKIn/5nqtFViIDlr82dijie4dwCR
3dUKcyuJL9oaOBYnjyqY15d+ip04DtK6GwtoZSCYYhzUPSMxZRwlxVirfDgvsdleMg6Kx60JA/d2
Y509UqLJhjZy1puEFGEnSswAKbGPXXPa80cwCVA1PHUSCABGz3LjvcY6+DHZMnCq+B7n7r7+l2qi
ZyulB4ve2A/SbmxSSQGW1WI5PGsRz4LR8ph0WD9mnHm5qlf8UlXxmTFto2d6C+y6wmOG3O0vQNHm
//tW63HuwOP4A+mIrlX/s1yqUFWK7oZHJkGbKtX0ZgJrwdPaJvUS/SrDLCEFMRA8NS0aPmkBtcOO
SdnyOrQ7cDBKdPKSJLnlWLEDBjE9jraE5uT5XFXFtpDjGQmJvCzwBbhiOEtwc0QIE+aiXM5sW4qr
UsEYd2uYVz6QlH/a3sv9z4Eqy+6pE2/kUOKSW5nBXiELui7YDPUURTrniD6ZPof03FSmmPkiy+Rj
PHCrj+XdVOGYXzzuTSYIx5EGS/mOid/pwX8vPWS/dpuJwNcTOSyVN+fDj9HU84FU2tQ+psE+NBAV
S/lyxuDYDiCiDudibd8vuKgwRv1dBujwMctFJJ+VP5uQu5u6+teXstyyr/rXMbpZ4qQSJ23Ozryt
l3kMznleuvARfELpZB870ChAaVLNdGGHxykMN/vSmjJehFjH0bKwHTgcaWU+XbroxSSBr++jyRLf
J4FgHoqMG2rn1Qve50FeJMBOFYQBl1iM7Wexj8YD6bKBrdxS1aCyyF6ZDO9nvZpjKnCc7zHRQSfS
nY0+qvdYRCGfyEkw5QrUZL51vNP40p6eQf4CJedWcnaQB6w3Q8TOlV+m7aTvEkn/UQv32JmDs7hz
m2ji5sTZbqi9Me23HN5Ly/d/kqwGv4WYUpL96D/UIY2cAq42pRfk8yeS+gIAoMaz17G3uxqXoQie
I9l5ARbaJl/+SoZJPrjIJoDL0h7WZb/5hM41QoGJqjozKx0sa0wlx8q2EMfZK0Xey85Np6d3C6U3
QpCxUH48/zGnZKjTelBrSAC3yScllaRIVKCQccRQ8719KkohFCrDLW+4GmdbdmmiQr4afft38hva
gb0mc/0VbksTmwhUbf3uAQ3sP8tA3fGWU+zOTUFyUPqXRGd1CsTbTc0Dx/UBECvtKlRUs/gaLSkI
VppTHco309pJBmr2fqzSXeZwnbT19O+fBFcxLc7H1dkEcfPeDriMn/RYttBC6usMwBtaeareAuyt
kI+2ILo0cJ4kB7qrlPOb/XuO5YwCTNmhbg7tXVTigomIiMh27M4Ovwjz+IWjRyesIn6TogbFgcz7
qwadF13DHVD87TP8UvBxpleGYNG2e49rAM8VzuDHH7C/k9eH1JMGSh2hMlkqC9CZC3TNKYO0wI89
6/UUufXb0PzI+ZLuZRvhH19UZxlMpcB2HuCmXcAwbC8rPnG/PxNyqZEpHMqJAtErzaOyxzo4w0x4
b/ILzgEejEoCdB12fgnuLaHsOJjip/obGeDh5ynUTwu3jYWST3tQ1ioWKlgQ7Ec456G29SEim/F8
wF08WbZR4+4FsOlHACnzZpKz42MH6YfIFNkBo4ffrFMLKNWmPfXpBm2/zfMmx2ZH2Fq9pbNf7tW1
sOwSt7+u2fghsZu+xURF+GrGhnEod7a93x2aqH9qZjZVjtMA+mqwKa3eTaf1awllp9fr7DGhTA5u
0zvMkwK5LK4ZpOdzF5OLNxgtsXWRqAZcugmkH8BuOHjsb2jv0gmY6ZqNcOx315LPzDNajFP4iRLY
n/cwev1rVgq7X10CndbaphOiIhxFcsZzuTFOJJ6Wd2j+uOG7EwAn8OUx0c4MDnG56ZphbyvzkbtC
SHNQZbPjHgrmSbDelTfIvajT7cpIByem0r45rS4Z65P31Lf1hmbJGTaWMr72dDPhYxo57skgwquY
WJPeCtrp8TRUvkvFefcYtEmxPBGjTRhDeMUkTvRq620fEAQ4AnG+o4vsD+b86sKLjJU3oFuqWPIY
LU8JYsLGnk0wTF008JA1z0qFKj5Z3km7cyW+sA13cTVMu2uXwm4arCBCQLshSlTOk6PkMWEWo9X1
Yaeq8TJhrHb9DVNAUfhTFE7QT8jAskllhEFkJObxTQj07yFU7TRzhSEg91H/V8yKHmT8D2TraxEo
ZCSvA/O+sBBZKV/aBGJKmKS4xoRkqceZD3O9Y3n4MABJ6wZZHR26wWwCSYbXg6YCHXshPN0OX/ZY
dPE4ICYeJar0MSqwsJd/Po7WurOzSUJhm0naPZVZKuYDI1QiBbj3s58EDdFGnsIymSpLfLW+f64S
NshdxmEsPT8paPl3YZJXbKAFGN0wWOFm/fclhMHLBFJXvDqfjQSfpgF07jMWAGtRgbVNvw5JgUf1
gmAbokKn3PEksOE9vmO2m6vgm594fV542Lh4ugGO86vyriECJ0/dCDui+7ZQQwXsRjZJ6GiMNu8a
URIPRiYiGR+FT8bVm1stYjN5wwPeTbBrtKqXw1HyAb33a6/jb42yRXRW863EuToCZtG4ZUxhE/mN
LmPnoVhZpKioteNTJavTAR9y+5p8VxKauC2EL/KQ7fMmmTeqm08N2nNbYGZTDd6bq1nBv1nYuXDP
C1/ymlm3RnzkQ2eUSZUG42dVNtKvOQu31eeBi2MdJ0GKkry8z+tlbPHtFSei7DhH39pYbBQJePlP
eAIcbf8Qj+QMWBDAfHdJPN77TW5sXfOOgj2PtYvEMqPL5he2bCMYduK6Lt5HyMFNil49PZDK0IuB
5x+0ltn0B2tlEXpHMTIWh2JPtpKPEunU5VbhTFImmZ058Q1qe9useU1SfDfihqy5Bg/Tr2F486zI
TRwV5L+qAvpeWYKTQm/SUcH03k/hM9P9RSLlX9WHX2z9EE06//+0WWA9uQ1o7jRuxtPoDdxzNVak
agaKa/dUGvF8qrp6TSX3EhNy9JulR1+61kOLOn3CkfyLh1uKCKyyuWxznNpfUkOd1bPNpL5r0E3+
IFZnxK5TK9uEhoyR+NWHBG0wmkj96pWXPYu/ZtBzzi07z6rzaoFaG4a54hYua8BckwcDYtxIc1Un
Xqbjblj94StbJU1vtk3jQ0BdWEy6JY4qjJVdA4Gc9BB+UzzPI+2LtdaH5ESCRTpcXWe1orZ2rt7G
ca7ZSVkXgnUps7TnISTVFvCIicLgAgI2FGN4wxVh6KBwRaZTtJuGskdMzR7M8A6EZ7dPsGWYldWI
jMEMykq4lVIb34+5DW8xh/DjbVj7nGc5AJIWR8/09Vww/vZlIqeGGi4ke30xTIMa3UEOoNUCrYdl
T2iw6prpV1FC65nO2k2jRyYO93SX8UgQ5yq0bFewUxAhkEUNf+9Oh4jqeB5zLN7Qhh5HN/+m4EqF
TryM+xUqMztRAn8vuWYyKl6tC3Ql6C/hjxDDOyWsP59aWp50skun0wS0ZUQ7jWEkpElMKL6awvDe
LVGKaI85LtFYFJEGPZtsMqhfq/gm9NsRMVPhBs43y9cc9J72vgKbAVxFdQ57n6i3eU9b3AuQdHIf
Wj5TxNlx8gkSb6oTzVnHaixJl6ajm5qv8YJDdRUFIFvMlWXVAUjvZl1QEuj7GLsJXf7F/9NqwVJB
oJi2KG22qJHjYgD5K11XbRMlmKH+j/fV+0VMwRuhPR0Ws16DNPdJBs5uYeta2FLHJx4j1cooqKvQ
lwLT4ZvTRmhaAEMtBuBC4qaOCQBGhBeuC43z3SZWhEl2FgMDIg3PEgOU2VG0ra15GJ2xahWMJHdT
1AIvmZcWyPyHBMjsDdKOJM+fm90ej9SBFr8tz3oISE57sX7g4hxhwZ4pC9TVhz9Dy+V7TC+Kk9NU
7oMOHya1IA5V2gspsCw8Ki3NRNSpsa+7nY4tLXU6SDGR+YNt2VgTOgJHowZNkEu8Krkyw0+7IRuq
PACns9jHIrKTJmqdVhmAQYUZiC4O1ZS2bV315T1t3bdiUouAbXpm/Js+Z/FwEarv+zvM7SCA8PKw
95aKRUYvzS0rOHz8cF836cB9OiSKjPzSKXsbCGqHhsUZAbGwW5i2/HEjo6MjMRlVIBiWoO5bCug4
YsyGcTctHp19+5/2uXN/RyaRAN0LTEEGkB33lXtui/42BlKxb60xjEBjP5l3hTIYh58CAbXg4lg5
RRTnWRosNdMyquMk6CXGYosmlKmD3tTu+e92iTWxPDIToOEfvVgCg2rZwGHBeSVTRcR4DNFpG8/b
ZU6EJaNZBvccxYffmnm5KyY/psD06UWHW5npHPiUW/SBrTIaAq0B/loETIvLTmQGSCNAxI91ZKkY
UQXIhyrdFUmbgYLzP+xPpKfZSIO7mAArBt9ES2CP4Doc4RIm09WdPLS+YVHPzhXSCqZCOsRtKkbS
PyDkSVuDRnA0uC3Vv/GdVyNWAaDi2oPE2yyG09bqAbstpMAeMD+1nFqlYZ70v68geqZPXaj6Py16
VAPaEnSTgFCWrOZZgMDAMy0vFqHm6e9NsOF44gF5Jj2QyAS3dZV3Dzjj/bE7h61GdckGdzSzd0fM
sJdddOT9Tjgh72wA23/mvVlF+g+nhuOszZhygaRNOCiyC3YnnChf7ao1vVOHdy3wM7BZwv0ZMkYp
Y8HgTMQFUR4yS1a56D9y19Pft9s0oEi9CwzvptSD93c8trRx9Jod7/yCQz8U1SVXYL5rYDA+q13J
IJknX5yLFlDdCaUl56k9Pd5cROcKtw3c+LsKaLbT3cq/Ka5bgsigB4dG6sGE+kQUenrtNbFOCwc7
GefB/R5dXFJCqcyq1PhP0vIDvQ3Xgqueq5wiEg8u+B75aLSztOk+TDNr7ziBQOVw/seP/NNrMO8D
a1JyrbqYqS5qbJbBkBUZilCt+xFqCVRuJXchXN2dK60EIlvUzw6oVRbjQCjD7L7UBJfxcTIFX2Yn
PfG6rlbqugihyd3XmvIp9hv+zwIcpWPo3Ux28EvlAi+3LcwT27KtfwSb40sJyg3CBgDftLTFal2g
10DQnE2LhrjQO5YAhwmqu98HjeNPAN20grrh0NulY9T8QYs9ACNvZRhDXuvszbyq8Sn5jg0DLiPM
swQzco9aMv6HTz/uJaRMDrQT+2D3k1ZhGnTooiSlsS4tsESVCC+sAxHVvdB3dIzhbgCfuOD+i20C
1P0Lad/5X6SufSeKoiZD9gH0SuaBkKuJJUTxEeNAcEW9i4nuuEGm92vBrgfZ0QjE/9P2eNgyeYQK
3NwU1fxHQrdnEGgeZS+UgaO89ioka6xs3Jp6GIoOJiRM12ouzwR8bUScxiSG+zlAqLlm0BMEdw04
khN/T1cLFx8Q+5KzHhHuFwE75D6iVckSAO98gLVknrGFCCnXj4jmTND3/UL5yFA66dsOxqSrYo5M
bOdmJBgfOZv9trk3vO8zbCjLIIAMb1Nwlxd7PQctqg+IMeUg73egjyVIczm/wg73kMcVG0oZrbPn
LV1JDIodPvyFWrqKz8X0rabWWRoVaK6buxAv8Jns6KqPaaSe3hDoVARULSmPhzKFqKftPhN+QQpV
Gz0nlMhE0HiL6jMlnb9vhTDL6CnCvoiL52mwkAJlM0rk5OcBdqu4N4WGudYSK/9+x+dp2wtO1FRl
+WPyj5PzhzyhKSqgzI7ss1BdMXCHaTwm9Dlnot0zQ4gnmKrXzjf16w2NwYc3WW1MzMoMi9IhjeMM
mTxHhUdlDzlSeMEWEa/UUVkExWKDPQhc9I3n8cEeirPJh7/sQojBdsTfDxbSARUfcZh0kVsN9G3d
b6RuyBLRyd/2L7Y+dAcNZTAQA+rPB9NPHTrLFRXPBO2mnwaWjSCemnkVA2fnNtHRBepasq7FbKrb
B0w2hmTCY++r46OM3GxB4q8rqZZrcHDdMyYl9y8XKA4qj8EbnjyKGzSak6S7gwYehs+TMrlVd/5X
Zg39RT2R7Ze4Mrw0Bbb+hqhUVaXzG0rp+T5p082GOclRslfr+g+f8LXkeTWerLzGIvzJIy8YI4Lo
XWNVs7qLrULE0dpQ0jrOuanAVnqxJzZqA57y0p99kq9IyUoCGwglk/fY9qlns2VTcbCQmRSdL9ml
DfmpaehXVhSv5HCROaT62Tc2yVeFug1pkbvVnOq6j8K9bXZQ0dsejPfsV2Ip0sNlCilK5Ue4VRdR
acnFPqRaIDwN5dGSr5O8w0LR+TqWxW3hI7yPuRrLtv7rHMtNx4FfflSyXM7d55tfohiq6fg1FQtv
JBvMhxwIMkKkpHfqa8xj+c508ZPZ/atum4zBHCsO7NWtaFYkDq43tB1u9hH1n0yh1SMuc0TL6ocy
XkxEF7EEKnLIipSUX+UcC+y4lb4eIhoE03tk3zqygUGW6NAIIloS+1ENhC4/zlRj6vGxYeh7a3vc
53SWudkhEuqOpqSfhsIEhCTalAFs/axsG48Nh47EURPsvTJQSdEk541E0pL+KUSx7vBmuf0g9EqD
64gKzZ13Neo+1qzNYXf3vwjde/5OUX8LBE8L8ZtCdZFuyaKIeyYx9SJoIIe22X4jEXC/zax7v+rb
B9nieb+rXZTPN/fP+e9uYRtEzCD6d0bcnuUm9SOXSni6iHk88jDNgxvV8xloyW3k4K5U4hrAI7zS
rV8dYGhstGLO0Km+YKrE6V9Y2NMJjr1hmoIERca1xA8K5S76RREzKdErAsrrkzv6/Z98yAMq0LMP
hAQcRoIxNgP3Bbjf4cpEGOR/gQfnpTSKub448dWXCeAv/BnlwCZVQkl4Dq/PkkAy0g7rEQPzWCLi
TZkAtjQ7SLvj9LJI/wIQrISpwC8nCP1DpQDDR5f0cBp33hJAmlcyPhwMvraIz+yXFcm3HRPlwUkp
6FQC9bav5M+ljHzZovrcyir7989ZcCy98yWhCMrULXylZ9hoqhhFA07XnvEPJny6Wcf4N1EXHQ5k
/cFVBKlVYv5D32kMxUpAKX84t30hMCl4l4y3LeHmzWHcUCm+Lpo8G0VxbkTHtmklMWTx3sgrEc+y
raQSTD/TlCrLMGrfK5rxoUAbi4t4XCC156YT8TqH37eTrEidzPkbUWIPU3dFt5TuffX4YXWoZyKu
7HuA3/dvBFab436EKiPl6q6BJK66WvSYJFGo7n+CIT1F9U3f5z5aTgJNd3+MywaZpe6bpVvSrDbU
PKdsQYKNt4tb7/KCwXKYAtMZu5u9byUl7Ncmn6Mj0NPthVXTxWnR2Nbfs6j1oWOr2QdZiv4mmzsx
aIwZVwdj3NroRvdXNuU/nsJZQMiLYpz0sOX144yW+ublcAPYpsQPZbPP1qH1rWbSSyaoFEEz8zgF
Tz1ZKFV9trAF9EjemtebmLnu5XVcvzYAmw+2ujrVdoEaushh4dhz2vR6NQSBjL9iC0T0AcuD2ntF
lkLONnVQ+JVaOV21dWEkzysEOLE/fRGA5uc2LwqeQTIgiPLdJRXQ1IfqgfY7Yqx9VgIEPNYeD1+z
he2nu2/h6JBbi1uHvnfq6YZSJubWYNIYmImDs3rmCRmGcHW3q4axTjNWilxwEciMS505zinaG3+Y
evwanILZ+S7Xc3gy9/TIz543WaZzvFh9CwaSyVQcFnJO/XU7WVYP07ZUMx2qbsKEXYaJexUMl3oT
lNvZETemGqvv6apfBcONmprMPiwfy1ucH1nXAwLx5sZqNT6cQLfYoaMI9J5ftdU4l7DqiSPOtm9k
jpT+CCfEv9X6x6QdzD3qXHW3tyylpECJ9KIOB2NqsHT6oOA+lU9YcVVyyVWzyWGJZSjvKVqX+037
ppXTgJgqzyMH4ehjhxqPj3EVFyZgKHvEm/zKSVNkBHJpikgp8vc38iJgukKm7dQhakPpVnKYRFfp
w3WWVlIhwMLoHx0DtXbh55tssmDLWMJMEf+MJBNitR4jFf4ahK8Wj1abSTBw4JSweH9PdWqIzeaf
g7i23A+vkrgMolfPQaDJWh7m9tpz8DjTF8R+fq7sP6NLWm+FSUirEfo1oAOpoywyon+KHXElHdz9
JNY7cB+0Qr9vojQjFwolD3TLGKhbWvZ0pVNt3yqFW1TOdXzx6JcLquM3yb4Z3DqLhYFNlJRPwSVR
FlkalPH7mcvJ8mpKixt+m3Yt1kRZlDTDPIu9UCg+AOBevaYnPEegE07AgpdaYBNN0bOR7LUnzvGA
Sn6zIgeXdJcfGm/uw6M2uFMsMdqVUkw+PfsBW+mdGdorB4c5C5i9/yu5IQYrrDCK3L0gCHUz0CtU
OW4wvN5IihBNAOLGjrah9JWoyNwUL0VBMMjtRwhC4mhLAvOwJcGir16Vrgzdzh6YXvt7ORAHDQnm
HK9rVSP1w2xCBLDY/DwVNWYo86YuAMa82Ct+bEzgbp2XAYg9fkX4RN0rFbSTahzDZK7+lHi5Ut/S
0gkItKSfc6g37tg4hq0G2JOIOsqJ/mq26gllwnMe7hG0wVejwc86+3dbOfatUyP/MUG2zdBN7lN8
Cn4eRxHvns2+koKVRq2sU8w/Kpfd4TiY/eaDrG6IlvvbQfOzMS9ro6b2eUO5fvYOArlpglKOoS9/
JsiCbG1/B8VtmcXRkO3+BmJUtBFJDF76lmq/AHObdR1ryBfBTD9jqPIwKC/PDvNGjaS4OLmGFliZ
M45f/avkGfwbONymJ6DDvMGMWDhM+plv5SfDefyKOOUsMNsEHK3IWIoZNotiayZ4kfTIxlDwVcC0
FWFFkghSWZPlScZmSv4QrgjzE6R5jXe7T9tRXS0aMm6cpx6c3SgR6O6uUFshDRpWfQMuClthGoA2
fnki/Gnb3DO+VNFp1V8jiOSZJ1JP9EaS9I/idoW8GgzbgjELcOvjaT8uOPPK91gaj2bGeYuAsNYi
jN7UxiXfYIMAlTdtOlL3sRKC/A0t9iE4f3zNxU+Mflog0RTTTV8mG8lTkWCCDrAw7lb4hXcH/IXC
MHZSfEPLhe0GIlYsubuuOaE/1O2L0TJ/RXxb2sWubYUg+t/0yMBg0jbEkqjhzFWari0/HZPnckhT
TAKwYK1FYDCpDtGQGwxnaN1oBG9YzwP+NS/QeDtJxkYORkKsXS3e67E833j/1Woy5o00DfV7J+IK
FUlCSEpGH4cnQakwEeqlT1jtH42kIlFccyMXwSfXqu1w1trO6LGNpYn0nr4g4IDs/ZM/1n2rFeU3
Ndme1xWkHMDLTcnu+BSm3SqrseG+D9Me6vPGD5AuCO0WDHBq+qVYDlcs8Ik6vGeR3vSbsl/uBGhO
r9zKAt4wNBNOSgy/Rnb8BljsOsGQYpL1XcTAD8fCgeDf4RSKZBteJezcz7ZvRmJFlrfGx8SWhtaA
OtQl5J34/fzVpgGLZNnOzRMYSXs5TUCE3oKlYRNI/PRcnIv8/7qmOE6vIS1vMKmVZLLlyoOhtjOb
PXX+GzGbzyYQtLriTLwK+VKFnzwatZXvKGxVHOdfOxUEMqUWmysRWZ2qWfz0aACz2s4xlsGOWDZV
9srXxfDf6e1rs6LjDOhCWIlvrimkJAsjAoDRuDNxndFpRULhyPByXNNBLc4oQF6ne84Y266pqopF
FoxARwCmub/ywcX6DMtrzZY+t/7SI0HNBbXswqf+y8O+aJNuKUERE8+T17YDJTMMdDD9+JYYhXIc
VjhVPOHkBcwiHgVAI0ESSYDw7EZ5j4RlgC1EjuRa9VHyrP65mrYdRSVUcJ1vb3XlSSEjTdvJt0GI
JHY8xKISct/r5ZZVf+4sWwTaKP+D59Wb8FHB8Aekj7SGBjAq4cbMpyJwgDsIFk4d9sjO5RYagGfr
reuztynfvGKG3ixTaWVmvWeWSMM4zZDI11WxnHrckz7sqpoWdqsOydu+Zqcb06+W9pAP5vTx5kLM
KVVIOEKt4HRS/8IEnXQhu1SOQFaUH4RxGApvyRhkzrQlCANuB2vOGUMY90qoI50AVfmgF1X9joaw
m8Da8x/yEGUUOfnbTStkuQgYamZVzfhSGPEJbkWJWdXnZAlFBfLTQ+37AS0NulkLAxHXHDnC8b+s
lHoF1qq7anuU3PX+tZAgFBgyjwe77VW4e7/F+WpdP4qc2g7ageeaq74IDNZDZbFOWPnnEWGOqGJz
Fi7qWaH1AFkcmEfg8Dh7iqiv/0K2w0PvFXNDSFZW0QASoUccoVJNhbZzOZJFBExbIi3XIOzlTAR5
mZIVuKaYAmzSyXqN/nXieExJv1+OBwjJ67P8oq2NrPeMT0TxVlxxpp3bO3kIQrCn32N04zcAeTdn
oINqjL2q2aGJy6UGZ+ate3oUFnXnAPjeV+61LZ8HzLj0E0uDJYA6jR66vTaq4ip5sNInWXh7Oisy
iPgk3umHk/tbW4Wsr3b/Q48Zq6lC3Q1r95zBSyytuToXX8k6ZyrEd3ZclLoiDJyeGN54RTnYk/OH
OE8M6TE2K0IV1erR5daWX1CosH3YVk90yLegGqWgmOuGPfp/3Mqzxgnnqnepzm2hfh/LJ9H+gti4
i6pMhG/r/jdbdF/zEVZtbigtGnKYE7kiPJxV1Up96POfGCREkIbej5W9GO4zdMPLXT/pL0BxNGD9
W44jd4NcbNxil1GIKaacJ/Sf42pOuZaeUOTiscsCaGX195jNRYjVHX3aHdLBE+TOlZWSU+2XB+zr
V/hHAk/DD3XvjAmdiGkC2xNNj7ixgSjVFnQi6b3Wpd+csKggi7csm9pms0V+FxKbYWoDIbfrCaON
vE8PcWWD158+WnUMnYJsV2JKPaTzRTpX6lxmUkj+u9yF3jDhDZCBRPZJXA/QU7+PTMRieEYeaioi
35PFUJfucAPHUy7t2SuCnzj8juxwGALmouBUizO7MncUxzYqzw2kCvb90SWYhQafT/9YAedT/V2X
SdDLDJ80j7BB/tLaCrS+DvOTyyD6oHl/rFd4qXVORqyC9+kaRWaWDB8z1jmfrkYvSLmAmtuwmKrL
R2GVYe3sDbvzNqqSVwXXyjvAhqAAMa1RJhKAJyV/k6O9G7gd3r6qp1xFk187Bm4eipPxYBWqQVzX
M/ja/A6ac1qksI8carGR+pJq6HrVUZoH1a5Pv4wrkZVuXiTJQ0rl3FmIL2J8gEE9zhDyABcfnmNY
jemStXqM22B1nCeyrF/kwZg5xQNZid5H7sRNiPdSbYMbGHZ9EL4Y/3CYe9sa035DP7/JeRm++dXF
nJcbq6fFBxFP1+E8ZMHKZRjP96SdRPrdDJZYDxiQtjUUQwdQpn/yk1wKnyN6XxijqDvXGqSuUIw/
bV61bHckDia3Ejvhew6F8B9OYhyUUHaycLEiwK2DiEnN66kW5kmVGEg8HidTXsm9Zrlvnp1jN/8+
N8oPcMUTujnmHkoYeV+CuYCGGMlBTENUOhd933BLd3eqkJ0P+tgQVjcDV12D0anasREmFmJKpUEg
dr13rOiGGWoMdV1JkTFapORzxXjZ1OUcEdiTR2eWZkXZFpQ8TfabFCaHmbVYUPleOHjz3UL45VHR
oFcpkGqNcu413evGY9IcjWqR+iSUXwHxybrNcS1KIQryCfrqrmRdSFCr5xNRpItx0C+2a7JcOOcG
EOF7QrjogBWN1q7Jb3Q3U74lCeY0QPZPugQ8p2mwuJA4DEu/OEynY9nG5PqIml6Zd1r+RDPkKTCh
UwZwAAwo785QubjwXXCih6OK5GbBiVaqu3B650LSz3z/8P0QMuzJp4xh2wMGBn0YauBx7b3vTgM7
+9Luhxowa9Or6+IohnbyNbLVA5nmhb2g72idmtVEzpvTmjmUAICbbKYV4huFg/CylIUPMfgughhk
YuXl5sOCT+m0LD+bxtbpg6se2YR8rb39uKGn6+L5U4mal3hTyVxgT6PdddTdh8g0mFLwI3SfZmUI
0E+jPeQmvT4g7rYWQHOiH9L23WzhLU3r0bzhn5xMNaIFwA51oc32JWENsJYTIv4ZmUinhVOGMUNc
gfpyHQgkVw2/oOy+KlXXjzdBgseryDtLVGPpwbPBN3Otucs4iTHNcB4Af/0EDQWSj+Gj8hfB1uT5
lMUo9KBoUEJKy9xjhd0nDitHEoK6jhNZ5dzbZvmHJhDhzgDjSZnNT7VH8lRxVVUohb+zJQckeT0P
1NhMks68CxWPzdf2FOpwf4zQHFdre+4HFrOxtNafNQkMomagCDlYTp9RG5tEDk3f/91a97uscIkm
oaarc6jRx4yqnmyFpdwkOWu2M7lhfSYDayAVkJraPJvU87db7CS5Sv0ImBODTQvGwJy68obLCp/O
7iMOl9tt04L+nXLeu5/4EQ3j8xk8Dq3Ky+bLzXEWCb3h9hCTiiWrdqJOlhPad+hSCqjmdmtNegWH
tUWJjyJqWf0pFxEbrBXtimS71vkpxPEwBKHVgsNYMGenjBDu+pzU+2yvbOn8pyRwpiioV7pTt/jQ
F6N6z/2AwQ9WgA2EKDKx7PUBskcr1WMjnISTD9o2WRz4bLqUythC/amel39g5/+CHPPKGCS67nXD
rahm4FP9Ag5Pjj49trX/byUC0Axw/DFGBg1V1+VcznPwrSISYkBUlmEm3l/i99V9q/aAwdDXgR+G
7ckYVwUZSwCa4ntPbAjppSHuCFs4MDQ6G0zsmgfYULU/q+8iYoRkTanh5V/JBE13yuv95yFOc15u
SMKiR4rDMxq0zNawUfMdFl+U3LU7KRSE9u8c/6WGku4OG9GGBKnRS+sHhcif1ZpV+07B7ekyX0Zh
A5GmttoBwpw9rKhvxlGWXWB7wlyr45KnrhvhTn8/tTHXnffh66RWAyHyNCx9wRnreXdlrIEyB1Vs
IgUxJysEd7uU/zzbgPB4Zucy8RxAi9qMUOQg1aTCWEg6MiJj3rt/H3sbazMReakjYdPp/TZzZlHd
xKCRHVSRB2W3mTlz7BbRJrzUuTIfz6Ta4L16M3Bu/abqAhzk0+mXdYJb7BgIVFQlpPk7L90c2pRd
YEzr2buJHxaYm2XuQ2gEz+l+36nQfe35K1NUETXipDUsc+boWu9IA6joUbgCopVdz3MZnGyQJfzg
K8bp5ongYiE1/L930eEJRWE6hLT4wI3f1FYvWwNuyugepJQ3GsRC+tyT/cXLcviG45ms126b2kJf
UNvEHrgKK3kblZQDiM+Pbtj5oMRK2YsvG2n+gZak0BkSI3SCyUVKFMiw4vD7KhynQVlEhFDNqMev
KT6+3RkwWGjf+b2tYBvEljAhh7Vpo6V0o0IVogPPLuNm9x4uT9rLvyq0i/NDTzcwCkXZ6wYP3VJw
LKEu/aL1zLPRuIXt1gKT6hJ+pIGg5QLqD0OSP2ehaEssjFcvQVvaL436+JEjfvqVY9azj+sIpdef
W8GI2dII1DUaxkLah4Ea4nNCWiZWZokdW5PecvJ2Vrf/QZblJUSqc8yyYiQwGNhgCv9JOHcqduUf
Y/juzDvTPiL8skgv/YExpxfQeu2sXWFx99vuaFUNj6vbfD5aqkA7TlXrxPuLN9lKxFGxfMaN6HW6
ORMZXmW8yeF2mrrBS8pkd6QxtOU3fDO7vzTxIINHBPkwQIYy2JAjXXvzuP8bjeD+bJT1hGoemi82
kRvP1pCFhbM+wn1xK7WWDUEO5EZ9eHDTaMXHVcJ6eRxR3+EcKHayiBATdhNvoWtYgxFEO8oZ8ofG
n3iNkrQX13gFdj34e5NbM6RlIGXUhWOdQrADDE137gY3sW8JsfT6iQmvWC1KnwQO+ZVXkY1a0NP2
syUVBovvfswml8S9+I040tb6Mk6l/oFn2ZJvrFfTpTcZhuHAchm8ccnSJLcIVQ3JV3vDyM69nOl4
dpINEbZuE7ngIVSYyMkAFjITggy8TaFfFM5P9XZSVxL3zBSlk90YOpBOZhN23eVMXeaY7g4NLtdF
yxf75EW4A9sErgcUsZtk0S3lcvK+nsCHHvYP+2xVfDdLKyANNtluskgrNALc2vBIp00z5VwkE3a0
inVDG3xe1KzAHgFM/MxUu9U6ygVEhpHQsVMb4YTLUA2ZayzwpbtiB0rhISH6D7aZqWdnW2gGTR8Z
/UI+F32vvjhT2XgqPV6v5XGDTp9js2USMzPUQ8r+lJ7fjqENkZ+6Fu3YcsQEX7dB0b/GG3yb4c52
ad6GlDGqhy6cDTy5KttiUfa0NePUYsQVUKYq2d22KGufifvidVv8U/Z3vy/Mk4rc3Q51aFTzwaSX
MWwkwFimSumbfisX6Ydsnk9OPbCWMeahegNa3g9bIvHMzpohnaTO9R7KzrmEftIAAem/XusDAtTN
M64gcXFj3CspEdyBSG0ZQv2pADbUJjXbYMYBwK6OCJZtbnohC6Wh+4QLRYavRC8XXTemfFdpFSot
h+eTVGjacidw0iD3IvgTwbdiRu4Yvaqo6d9xTFlt/G1Ni+SBK6f/JwMZuNkHmhpMtWQ/gSOZB/xb
2IuL8W4/q4/b8C0WNtmIZ4FHAxawH55cgg8/B2/DYaLwJBUv3jAYw4HQOGpWr1u4g5k3NhQJ/qfM
UaoGZWRgRvyKnlSEWTpGObITEVUvRRNc1q126PEMNs3ftfwRaWCf3QVv0I/4m9WIgULqTNwRBeM+
JQPLbQutZsg+gMGS5jxwd5+V5uFv1GF6ZJZeqVWh4aOGLm0sqFdyqRWMg6x0sxNJTJsSExJ9CjWW
pap704zsR475CtMLpKFSOFmhNuwkTnUKErx4X1zWpcpEgVYn8lnOPY6iCJjjWpZ2DuuLev6QJw3D
BW1KiMkxmjbC/1Ac1RVUFtwnM05+iBMt6Qu4F97FGd9/ZdLRFgcQ+25iTVKQyGgZpagls2MVbs/c
VxXRWU6n4tzObis2mj+Y7jV1JCLtcKRMtNc1iAFd9DSMEnu+zQ6M4X8ZbC2gDDP2KAEXrBN9UesO
YBPZrAgCkPDPhDMl0WlTyVdl9TQV53Yreo5KqIDh46RHPKB9aTKAVXhe9Pp/+FfDXU27WkZECXVO
/5eAUY7SS1m2Zu5TZWhMRQ4STVs7vEHL8hFYsduFLzZcGpAR5YsEp3biYQY/rcnN3dMw4/KXy8ua
Y3s2/BVEn+bnKtozz2nKQaInm1dA8M0PiNBDRzrwZ/9b7swVJelSbGQYumENGxYisSZhX7JXcB2k
YT+yrmTpW44ih/dW6egV7MfMgDrBUUGs/XlvNpTYDYjaRh4Yy7rMy/hmIUDx87lK7Y65BqJjSkj/
FJfERsvkRKxCCi8/I0pSMx1t2O0eA8AAUJmY6gUDNuVSgxuAGbW0vWNkiL0P5t7k5B5znECrl/n/
JQbYZyXxiphRyhDVFdlmdq4TgGGwcx4rHICgZiCZFPc2Lq3JwHOxJzuWCUKG1oWOimC1LQXR4z+C
nSGuzrFCLlcj9VVEwuZp7bjoOBcQP0QWd/Kui0qBxeX5nCgUeOPKt7uZShXJD25dzpDeRe0CWsvQ
ZhTPVOyvIm+TIW6SJhIQ2N18eLV536Vn0QDCzbk/rWxInzQa4R42yH/wE2aeUYzOo436MJ9niNkV
BYp5m72TM1S+VyEk+XE12FBuNd1nB8LnZ0beJoSdvt9MvkylJweTF7eRSZ73lyK3jWj+jHjHfEVS
sh0sV8U6U8J2dH5o6VsTcFt0bdDJf+RPyOIxjlSTg7kgyf4qJMq1PZruSWv5gqQY7/VzZBeYD2hQ
BBswK5g3W7dH9nYNc2KSTfDlZpNSQ/Xt1J4sqzCvqmcWDgrsngLsjSUxcRdt0D4CGKOLOJFp3aY9
+oUY9Uo8YQOo6ngl3RTIev4baLzs7EByO4trxkGXFTnB8eyhxaCCZzXIO3PtFeeuEQGH5ZFItuV6
Ykq/a3ltyD2uJbp7EtDW1XLQ6D92g5ubnUHQXZCOEo7Pm0Rz2ZQPR4IW/8rOoMmseKgox++E3GAb
5mB2Am7kcxb1zmW1FpXpUppIRcPngNiyWn6KZLx8RA97AHvQt39tEuMaf0RwrTiWWnBkow+zJjvQ
FBtZifi2CVUolsaKtKrXx621GILoZTXeV3t3wMnI9I4UZmXoVmCysANtE+2lENZZfQKdEAzlwHav
jur4D8zLgytWDsxmBOezRAKmPixEw3VRsgW8OA/k1aZLRWY5GdRyFOC58PagF97UNVvR15Sw760O
K8HcF+nRVl4vYEENBIwnkUOWZ6+BHacZD+Lx6x8ulJUw/hLGdRG6b6yyb5IXm2oL7c3K8SmLLRXg
0FTv0wr8rrSitbXc9HlJJFqeHFZXOuf+rFN3YI6X8Gc+RZvOMdzKKNkR/lENQWAS8dKjf3Gm4abP
LBTo1yUMRneBORn8j9/5d4bp1RMCIzPI9d5flAsfiBId/0B2imPLQYffKvuHFGPGCIGNdlWPLDqh
jFiS/HQ21WwYTL3cdIyfEKoei/LJpcMhl1IfK//9C1wxQSqRNh8/LiSmaAATs1IS785Oyy3ZRYM9
1W5l6IStt1GESS8obvNAMs5ByUiH9k1RbohP5ePyYvbNByitEd7NxXHD+yyLxZJgIqYfReJtQFuZ
Bax4G0bY0+wkdsi3yLrfthehV5gJpLULQXZ7FVyCGle7VO5EmKimn7EZGGJx4u0yJ2BtWC8LZYkv
GbRKgdPALja3brzCLJRRj3U8Ou6+ujgGRq86XE3Iig3ZZdaqvSujgtX28yrQLpZFEkCpNek1H/jZ
F7waZCt7uQZqEfx2ZfxzQzlz5Jq0Ircsqj8SRjrumk76+SQN6dO7viz0ArDVCEFFM8cfLbQQnike
4Kk+rRQJrdMi6Q7e03hn+TdGA8bXdTEoItDYb9iNm7CUaeMdVuyqiPYYuoHAEXupfCUwIid7YZoz
+CjaQ/lJfzoUqql4wBDPEfzApH+QNuMMxD74lSJWsQehHpHYaQHnT1rykuXKbXNQwpZx01V3dzes
RfAJ8C6D9E87Ko54TJB/xY+kpKSsi9Ym1IqyIwuz7LkTbf5pH3iS+Bke9RXt2/H+xnyrllyy7236
aCh4KT+LxoXoYLC2jg+Ofp4s5iWzG0U3fkOKetYC4uJY7bb6cMhdxGM5O7w70DLNI3OglTo2dCWO
J+OsRW2DCvf2J5Sy9+B61v4mRbnYRFspy44oJKi/oYHH+BscK2OwDjBRA1ZYe3cNmEJF+1tE3+vN
GUQTpcPLJhFLSvwF4MTDbS3oGqSpIoxPgZOzb7meAmKdbR7rf+ofRzDxW4AoWB2vKd+cdeET5JAy
Jf13u2XMioUJSc/pTr9USuEvVxb41/NkRxuYRMGpKO14dkCmzl5hRkKhGj6TQQLqWPikVGYd7sPr
ak9Ks4NvBhcvENutbPe5cjTEqjGJUmqSWAnuTBcA6W3s0V44pCRfhva8yuvUjyb5t9UBjBuN1+D9
mPdoBJRCW4BlW+onL4CeCNTOSF2G8xffNKGsy0V3gplhxGB/D/Pys+MOoEPBuUPyIPb8jSMvwe/f
PBjiey31SWqTc3EGi3aFoDr1v/scXkCULcBM01IUsFQ3ILByF533sMzHik/tNry0VgxjDO0scfiK
nAUIdSR6VuMowunKVZZ++hPXnq+Z5o/H6jqzuayZTeFsPd0lvC+BgLHH7WOphY9DuQUqFyDKf9Qa
iNA09j5Y0jKNRqGuNgkpjzrnYToxANZuRT4ljVPLIFy0De/IyvTaU+9QYzrCPiEpWQ3icjzw6VsY
1C0E1tAm5pnZiSiSt15IhlmIjFBXfWAH2H9DDgXluppLfyxRtqt0GjZutz3FQNzcTMIUsaKlDUMt
spaZIq3FSZij62uoCDdcLb1zycC/D5+oooZVCdfXsVxX+fJpMy2d4CzRX0CXlj/ga+0r0q/46YL1
KuRyDey+6q/pJRpJVhf2lv9+qmaVDK6lfHKT+QexK83nvGRI8VcchapBPeORjGchLLYK85yegS2K
p6hnHg8AMkTtDImpN4ryg09tpshuM94dWizhAUpsVxrFzoDsvskbVAQVHGvpCPn2cw0+Hwy2X0zI
HgBgf+6lIGDimuzMxPtUs+K6GqXrokIIC3TrrdPTvKAdiLviWfRHjX+okdCoKvyW/9lGGpj+J6hB
CwQifXawZBDP2juNT42EKVglO51KFgOvCn684fjZWCI6TBSb2YA3RqWIwPDAYVfhvABXO6bFfqVj
oYIUwd1bFCisE4qRoCpLvRu5xUIdQ4wmNoSnrqiXpypE7smgSZddL1mdBHq3HWoO/ebZ+bcMQEVF
gGIRfUQI+ZliIt1fxVO0eTbRvZY+/OZrSdYBp1VFdJttDpYZCoEPx6JnWDgkYy0lAYyoNOF2p7PS
3+DdU1g+Wi/s2seDAn0zZaWggXXh126GthfwYwLhdyCysajnZEekVs5Szij/bN5pR8mQu1OHCwTW
0xr9vSYZ5YgOhQLxO80/cmkNqAmsHiyBf/9sspSLABqMArIni/srkDo2DJsn7mO3Am8PoH/afqFk
YM3s4tjgSKUe/HdN6AjwbTuFYkzdRkCM3YSZhsFuzY2Z2nCVhJnC+2W1UMrkWniGhAqjDhq50uUU
j/IpCtdDG2pPT0JpLmR2iXQEaQb2n09SobcbYtMDZQ5v5eUd6BhFr4Hs4KodxQ4o19pABRQ9fogD
EHBEKfagvqzZmHhj0Xn4eH3ZP/0ZRhIpacZQDoGEehUAVz8lNwjTLllsOi2NOYMFBnRsj11JPzZm
xbQCpFKZRKDoZWQsyUvrM7EeTvOnC9ho5PRsXG0rA268yySme2aQizWLlcgJ+apOEE+9vL4kHNr+
4XWBMtP9RuSNdsAN5l8zaPQdcnoKM9D1T1hzcRimB3+JK1gm2RWrS40VMvMRxAW5aPWjQZWMmIlz
DMW5wtgdNayP9p1zChYlD5ts79pTnnVaEJUonpP6hgy71N21D+fy3sTzXjy/8S+n3dvy8b7Ni3cj
06SMrlMhzrR3QuU9LyMEsgZ+woLNos4O0bSB0WObdkA6Iv3mAzfkuP83kn9d2aGCiz5a6icwnbtO
XBW+mLdCuIne1oJaEHamXsPVt+VyZoqvHZTud4OPmlDFs05EofQo39KOIg+7Gd17sBQiA01uKiXD
vagrhbah7Hf2hxe13YIIUqMJWYj2/CNyrCECUjs1fNCq4S3UzKnAholzQo4jeSDiAzFmlnzQrLih
GYkoevNXoVlSbqjYoPt/Gdrkj6K88UC6QKBgJ/m13baDTy7lmyNHXOTjjJtCs+v1orof54PgE/MN
FrPfd9DaOgeFiAi+OHCFhX5Td8/D8IP/CpLhJ3QJl3/k0l3bTP/6ct3g7bYlAvHp0jh737/20s8D
Gka6P/k1MJgX84NRV94DLSTSGp+wIgrjwSQ/cFLCIDSuFxNN+U3g+afj0IBZwZHgs3a2WA8A+8ui
pTlfj1R4S+Zj7YgwZcNpjTVvd1+Pz1eO49sHpmeSVSVp3DsttRtv7Z99lDr9+BZ0jt0zHimWKJN4
dlpPbASHYX6x8xKJBCeNOqDVkQVs7E/Qrp7p0RDmzjbjTkuMCbowKDew1EGK5GX7XKyRRbTfXu/e
wYWVdQyS02eKm9MbJrzGqK7DnO9D90QOgIYYVr8XnscGVJP5wkqAZxQyBa8f7D6ZYFt0hVBND5ir
0Xdzug8nBv9SPhxOiPt6AjhjRd7GKPlpGUESEdijtZaapyZj3m6W3BAvRoOXRChhgRF8KGzExOiE
UTaNVvR9yAzyn0/52h5bbgw/LeHF0rlO+VhgJNAvqfj3SvmGx10Eb2/tdIWPxBIXKbrC0ZuIML9C
zCSFvyOD7QAq5ard2bb7OhEv8NHxihJwEl+S1av50ndefEYEETnGFDnpuwy4YxQhx7RH3Vu1SHZb
TEPJL5uYD6s2UWYglRkHidMehoKctqa49QTtYjJBu3QwafZROyeZ+RKfEe06B8lNpuYew9lwvrKW
nQUr5m9h6IADYPShF1x2tUTweUUlJBilnA9r/LNHfi3wiY+G5kFqajh77rB7+4DO2q+yVroKAtbr
+TGD9LZ8AvTMT4e+QeKaYWsjrpAoNUh4Le1/j2b3GfwM6ck7Mo2ZvMmZa9KWTGWCI00M8ShzvDpK
F3TTkuBP2f+YlHvAAsCuLZ2GECDl1+GiH7HnDcZWZQM2rpDe8WnVilXIvR2YhsYiSxrt8XBDOWMd
BMaBNd+F5f6MsNmWJeoD+hFovM5S9hw31NcOT+KWAxXITBq5UGTBIYJRDbe0XD4NWKrU5rtg5Vro
6LM9nm9w8ps0tqHtOtlNWV3cy6BpWyMGhG36XU9BU57W9/7GH857DkcRIlJLCvU5F8GHTIUCc436
hg8Y8TVTZedPybyCHFaXs71cxKApj3UratKzD87EWIt2UvWQMkdwmMP6FsvU3TnZnf5nv2MLAAde
2t5ScFo826gm/WY1SzeOEjTCoS1LbHbolTJkZo7XT/Rqrq5mzZ8rDLVeJQDKPjbZiYbHaLRITHxu
FDLZVPqO4Qq3l9O0yvnu+cuPaE2UalWKy/PHLMG0db26uyTb5tvBNVr2zghAxAg9o04BPHuBNadl
XSb6E9cg8cTx5WuBl15/Epx2AXoNK1nTdxBD1otVrqaRYk0xi6hgn4GlU637rYriAmZiG0MpjtFV
laAjBrT103INytFh62vtWgNqg9JAPOvbndnJ1HrSwE9L91EfUGWp6FhzowopZ6vk0FsOMHoepkXu
NC4WAMJjGhSf9KjmdkNt0DrS2zRl+gpyusWtQgXYfbB2eC7+tHXyqYBcDygV/g/sbHS5ymrLDZGv
DedKb8l2LlTli11PB3ac5sQW1monuaV1SszOlsKnaqiVA7haz4KZthqvpurVsTh47tBc1CfUqhoy
F6qlQFhx9s/YQjWegzS3fJNxJWWeX0o9DY+uGGiDbTYDavp/saK3lUMNxlK1T2xT0IVgctaXoUmV
i5Z/Q5ZT10aKOQNfvJD8z6sl4V5ycJ2U/rSBDVqEWDreA1Sgx/3bdGORLwIQF7VtWDWf+TIk7ZN0
gJYSaveb81zEonUN3iKJSppOXyYGGtmG4/7kpQBDEC+6wao4E2XDoCSUgIj0bJorZ4azXZFiFMTh
m9fDxZETveYyKktK948RklJVlqqnbOU0uY2Hql1UEe3dfiNBq1VwHq8tV5pKebyScqIXrrczA8uc
vBlahv0BrJ3CxPemo3VJsHli4kW1CedQdBFICtBQMzRXUIcN5lUlnPW0I4LEjlM5w48kcTw/rMlg
2NPcHTeF9tS51m0YDpfuqp1GGqzESWtD6NAbCcY3ik2w9lFKhN+ISdbiDj/vkEhAbMu2vNQd/f3D
jkD6/ch0/s5MSgrgXpU8SzTiXXyfxTYXC9PkMYLZPNziYVfJ4PW1BJVdFI3ftpS43NVnMlCQ1Hhr
gFex/dslZKGiwJAWA3Ef1qv3xqZ/6mjrPM5L1J5wWstsSzQpnTqiEDDULKd3CGNKplZduxE8bP7D
6SyjBII9t8wF0tcxxWheERXPGn+TsgkF5/7QpHe3fLYF8CMa6d3w3Jn+8+SDcK9l/K71Ggk5gy7c
CLBTKvJiu+hv/dI86ehoVW7lC5EozfNRWEhOGbB57EHhtnY9lj5HWSoKr6ZyfgH79dlJ17elWkqd
xAh5DBBrqFh7B571PHy/ndVT3ImHA9vEllAOnZlxKGzxlSpFfyFNh8xhS4MRH8WndQGg6XSvn+cW
bCfwCx4hC9+vLzv93b3a7Laf+jJhrqao56sbEnObkiwCDzf1O+sbJccuPZDIDEM3GekrliPMLD55
oRRT3bRjtneEo9Hg04ETHWZMoaIU2wtSZIEXwbZ1teItVG7XaBZoVPlsvjQSIGc8GRqYu7+irv+h
/OX1Ax03GyAdyumcnObtk0C9rlCwY5eisgn3rC9PbSKt0mcsRNjAt3U/xYUSsms9cBLuaV42Y5YY
AhwaMt5P3deSVFJEMD5m8smV2EWmdQINq5D7/Kh23Ypv/4NZ5AlhKRYwYFeAKw8HfOPAASToTmEY
vB/7jvF9qJ/DD8YOh9BUsUOrp7ku01PyPSF1KtvRRwFawxlvxhxxMCkgUA8SgcfC2sut9HnPTglV
96MXOoeZmhzoggCZsiuo2O93oTszUbMl20mOir1eLmwhC14C4YlSoeXqDJybnvqG97GjimtvE5QM
Ua0G0efgIa7xFn9Kp1wJiL6L72R609i70Nq89X2DW+Sv2lKlu3R1kCcnZ2w6hJUNAiNm5dGdqlG+
172r9E3RzerX9FS6+VuHltg8BGFAVZLaBrLFxNbtijDmradCnIAd25SUfVM4nMX1hNw1D5PFyqvv
LRmYOi6ZnRNbkDr8J1z8j7iv4cipt5CHBsdlXOgyPv8fAAqcZEppobiZ8uFPi/mBgmItxOpA6/5+
uJg34kDXKZTWnKpoFTI6nsWvq5rYw/7YgQU/fZFhWmAocu2ajfLqgCsqU/QUYWw5iidsCjP4ePEG
1RTBTTXBZMLkJK+Q5RGyF09FFfn6HoED81PcxXPklJNkb58yzAA6xQd2PowJTCJl1b6LRvMSr0Ii
X7XaFlR9kxVyPM8PrEuHgpXF5MQnmyyl5v4ffzfiE1ks7+DkXppqyAYF2b09W0j/oVg54mXLyd+r
8sg5CuoiLCY3dqEvQY9vhiMzz3sc/qChmb9as9Lea6rci8/UlozFDbfaIQfGh6/GxOz007raoHj7
awDQsxnK7wmhAV5NSZK6hwCYAD8SdbB7dT8yaCDOMH3Q3aBuhdOeI64jBD7zou4moWi5K0OQHv4v
u6F6b+RCZ2comlV013xIx4yat4tuJvYxIYwrMER24Wmjaawx+ONtFj6TWtUYvFaj3quY+qiTsB61
cmk1iZek1pgm+9D9bTBnK8rRGaivJ83f2d/6vBkPIORjZzCBTxG0Nu9zNWqB+TaukWmuJEubBysp
NYmv1h0ICJ33AxDl7Ekwyxc5tdmVtV8fHtra4vr5TfJCKXMloYmmFZtbYoxaWEcOGNiq4QYmy1rT
ytjtl9pjg2sgMbRFZs+Im8ugnFDJxbuAeOg4a5c3mLIFhEHk8N4JXaBSPwYsDmhxxisepzdSyiOp
/j6vRfq5CqTrSuZXIuAVwep0C0J8bbGnNLX6t4y7ohPKBrKhB38XexKeRC05kTL/eF+VdTyY3Ujk
Zpb6XTq67CsyZD7KoLu/Hk3iFqMBAen3Uit1Egoj6MF8g5kfggblon3Bh61OQVYiOLdNIRoJSV67
G/Q8T6m55VdkpBxIJXrF1Me/bHfp5DEoYueq1f8vHo7kUePTgDmM9lD66+VzRf9uXYMkWV2wKkTQ
QdUzeXRnO800be1sifaC3EBrwVR9FtOGdCffCK9xt8F/IOpVQATfKsfiJwhW2byOoOVWOuPJ6SPS
9xWFLOcdsSE3fSeCZCSQOc8SScpNWgAR3SJMoZ4++CIoBdfOLqreQJMQhsmlfu+M82OkMi28k29D
H/8m3CFcDlS92NPueW9pv58Ry61xN2NV2MKQ/WEvBA5zMHZtO9nwTAQb4WecaW2d5TM1598k4us4
M7ytHe5DByvq3Ld0CQA8vF/zSnX0P1Ya2bIti0EJGMuP11Gv6kGJIInPm0SZyNF2EtoPUERDBU1P
ANTpzAwhM6vRACEmGvmEB/4n2WsryLh4R4lsdgKdTfKUSWpoYzVhsLcK8ndkK+tTlS7N2aarEoma
7c1lfETxnmqsIwbGfrCLXkUtGP+kg2i5YsZOw/geViFg9qpi2VTCru3rlYU/GqSFZuo5fNmBeVMD
4DjaHgjqMIkoz3Z29F5tQVO2LsZCfPbF3QtCkHIw9C079OpLmhuYFpJHz0aCfe/AmVqlVTbQiM3X
4ddiUpC2y8xFf0H8Vo9/Co4gjf8tr+0zhAeZ98jEb5+3zcZT0UYSj+Y0tJ1yl7xbvgzrLfhvTwpx
/++549nwAvnl8pfAUAJ5oklhxWhSgtNgz36VugdOGUNNCbhKCVpuuvezX34sQmmqNrMoTRInKk+3
O00nqp2Tu6H8mo+r9yLyXFzNwRUhD7dU58i9QGVoYiB3vwmC/+YBBchhwgcBbKtoz17hdOCJkLQu
Etdsz9DIHu5VPekfBsBIGPSbZzDwD09oiABSr4OPyGgZu1bw37J49cOhAkGwVM3xI1hrklMG+wNn
e5/cZ2HK5wU+OnF/2wbQtsCuNl7HJvW1um32PnK7Ys/rxfgpexdYHFEdh/NetAw2HJO3LaJH+7ku
+O36uBxy6OjBsRQ1gJBsjf+EgZeZchHVAUmgupajRpyYV3p5nx9iy5VshdhsQSTNRlpGVySyAxOz
qZDVYaKyJjc8/IvwmOBe7acRAQx683+XfUb3P749kh0u5QLf+rlyuSGAByVWDk4DZgWuspsV6CjH
E0RAnJZJ5qtaTGEMH369FzM/SExkiHVuWoiQ3K54Z4yfgTxw5G4zqBcn35vJLZS+riZdaJi0KE5A
ARRAHU6+Kzdv/7To3HWeZr0NogGxrLYGOBsCXB4ERHAS8aplatUp0o1Vp0kKFB9byWfWlNwd+YH0
xHuBJq6ZXjZuR2/3tzTZT2gnsiR9QnvBg1X6d1likPXsHa3Xw/E/kBn5QbeVT+6a8+TyhIBxm8UM
cQnGy7xUe6uC9hS5uW8MxtKr4c65ZsLjYALM/aqBuzOcpE6oWtSBHR5fykNRkD/RBc9yIlMnLwaZ
5TrgLqLKQEnfHL8fwAhBYy2t2LcusdBtHbymHnEd0frTXNhBEN81wMQ0FPlLPffao9Iy9Oq3SSDV
433ueJ5+7sxHxV6tBkZnZ8Pt4AODPlYATm5wiewoYiq9meppFekL1V+MbBwcs2mH1ZMCwwl5x4O+
Fa+CN4YZtYkHlxsw73Uw34ou2DTeA/tyP9V5jZI910bALHMPmXHuRjuUgKOdDBqqAT2E0JkKsZyJ
27JDVC8jmLsiGZxdvT/W9YNb/0GkW7riY6wty32SmAkXV2VDYJoVgEkUHMrq6HBamBLTDS8uQzum
MmnB7Hx0rbeCNySAYN7vYBL8QKSP5UaT7HMHo4s0wNzx8Fy6Q/h6ZIffJvz9Ss2piTfe4Rz84HKC
3xsWvlEOY43MTWR8p28FCjtjfXk0T3t6yIao/4ZJyZ+UCcRXKBTJLF16xzvCYT33Ti4LQm/uPJKc
D3+bWzeXHOsZx6SpC/0rfh0mPGErcwrsnQJ3qtgKWYBlzLNvp9MQVRnBSucb+7vps/vkwxdbkTPp
dZjhNDACBZUSc86Rec99Kf+tGQX8p4Mke3IIfcKu+8clBBUj1IF8BXqE51buYtOBumQ8S1jCg8fx
VF+4okdeT6gNpTzC85P2aMzuCcOVBE1Ij0f6u4FvlQzIFKJ1TuJ/52Hddjit8jMscKiNStIajhEX
Znee0xdsZViBC2+BEaMTF9jvmdZkmzUNW0jRc+nHjNzkiFaq6ckc0s47TGjrrRzKjzwck/vHBfY/
+WsYZm3b8fMmbLWyk9FIybm1SGwHCPjyFTXn2c8VvlPgM53MDGGZCpqr2PLo8tlPb5jYCulwQfkf
IoOjnGD7TO5xC0VDiQVUxT9U+EKNO7qtqCKi8sYh2usulmM0xuZ3rKXrhTKpQb3foK1dHsUWpcN7
AQW719BQQohyj7+Q3lENPKyx6ANciKMf3TM6b/7Zo/MhzOVESKhV06hjAz5/jKytfc6posK3VtZK
KojaX8gb2zQtMLQVpVzgeix83wS5O2QLmVhZrJSqR+3mvLqmYhO0RPvXWFIQaKeAZsiTMroquRJL
HyONsiYaKXu6Sr8uwc/beYqBPkJIcK939wgIc7TJlIRUOPfyHm2yTJRaXG+TS33CAyjq1pXLYa49
8XHXvd7YfeKm4E1zS55vPtayXV/7wTonuik2LPmNvGhScnZqm3+aDRqQf4khxNhDDMPVCaqi6/yo
5ZVYxFfkH8ZcKIQ00MxBhCnTD6X5M5Pz343uQwBR4WSwFyR3GGjRCFc73vm0i8MJk4mYhftmvEYC
/KMJgL4lzyApqWxYB9wr9xBLqSiMuuQVSExPN/K3W/H8DwSuPRtj8UaU9sLSFYeqm3iCi0ay2Xj6
gVSttCkpuCBpP/Y7gIlh6PkAMZkebFvDED7JxuGx7LtBZQBxrfngWDy8gC6MoL+Ud+kS91JKFA19
/dB/lU6WOwb0VJ27eMP1t50Y/ca2pJJELvRZtfOsClLGVAALjwmUrB9EkL6OxKdRHm+lL72OAhd6
5yv1DyZeBItUOV3OCTNTJN3ATvPiDdELIM/pHo1Pzzn2rgsH3XM3xoZKX+y1bDM48uA4bFXeVy3N
2+gOIE+GAX+dLyJ/YIYQS0wexbU+tl0HVbeYGkcmZzW/3CPGiAz5l2y8uDgnCOQsS5Pq6HqqS+b5
z3Twa5tF67bYweTL83SavWo4GTRRlk/DzaSm9WWuaxrZGbW/uU4j/tWm4JWF8+dgtfJ6qXEhPsfh
Ke8cdrkRXfdA0OmWepnowBzrkKmqICbfJdZAAmy+i2ABalM21Y2IZdPDGjttN8q16dbA7/O6cYrC
6XixJtJk1m8BviCZMCpJvmHf3jtmxbvk5G3NrJOM9JjXdYO+70CcYWy4a8VDFAGVXAOcFHnx3ql0
7vCZ9kQmDdvl6UzUE8VHXcEkQAxicEoc79t0sFOdj3tvpsbAlf5W/qH/yFlxr/CKOdOsJBzt+ubA
Y2WuiTM94u6RuTbkQoD7plKwDLgTs+6VBk1IkVrsXTKOB6xvpoM6WrPnPf+A+lfynYp5Rn2TXrSV
KU2isYLlw2I9WYECqs4nTOFtxPyU20qXRY4+wI2o6JGeg8suLw2cfDP71Q1lPLRORjhPDFxdzFyM
Z9/5/Eso2iPXUOusJ1cnTKDZcCDqnENWicb7h8mhcB0QhGRVI9YpkOAnv8diG5rR+zKa1+gvRRre
D3oXYKRJQ3xQNBa2vP/j3f5/MTHaWbtzrwUymSAUY8p2vccN9db5VihRGfxC7/F1Y1k1HcEPgjnG
KlKT5aulBBP3F43slwhTIiydIhsfjLHfjiJhBGcsLCZ6zlwprAy+CNaW533Z/f3tAKdpMyrW99DC
z/ckpQXMAl9ueX+QfZq7NB1Ropo7BQPrK/bFQ5T7LJ+2hmTiyB6tlhPBCqwi17MJ4A0p+TrUKrq5
hguijxEeHGZakdwmRprp7CQg2X8M79Dnh3lZqdeleZzWrm7SU3qCBS04a0JBz6M7JqzbnuaeXqWT
+M1qxopTBxL+vlsxl9PATGQjjvpUecFTC1N9Gq4WHkG2NegANe/KCNHFkQLEHSQ57mC83DbRSxZJ
ZRl/Nhiw2ZHeCfJeBO+rRw+0T+bdeCSQim1Pi2qDtYYHjBdOiddKA/JYHg0lDMxlsFfieI+awNBA
Sh0YIgA6xXy2s1vSFhw94/t+8858Zoi7hUgYBBKp9JoUFa9vpTknSUdOxT2VteyWszxItlYCOsS8
xBTddVO+Hl8PWPnfq0zOh30vRlaKW8okFwjhRJroa8VzZUfXjMYWCSRlfn/k+5HAlzTC1UH5tu+r
3MpPSl53pJBoOxHCxgaex6PrSbGCE+Tc/L6fk1GAwAmlSLNLB/To2wpLO4JOfJGkSbUSGF+CjpUd
fZGW7E1FtJSyZVVRhuGiUGWxQhCxZL3QmouNCp/4qadVs+hRww0qg/RNkhfE7OjNt0FO6Nhekpxf
pxNgq67yMphggYpK6RRMgqXiheVOzhMuJrVJPMy02owLWoiZL5r+wK3DSCFJMhpYgmIefOpQZwdK
w4sgDRytQcoLFbXxhRiW9CE5LFgfBjACCXd4A7Lz8khcPRT+PiTi80j2lMDb+cFNGxBmKiausNJE
FFpV5HdDN1sNIAQ9tviKzdy2JMhUbLi9uOBk5iinTfGCR1m8PViwSPMJ6tBPs9XwMSdYiQOcSxlu
RZT834e6Q+173vdMGr7Aw0AAb8xlwnfcrta9libMU/fDdsmq32Sk+SxV3UPhtEddSmDDiHK7k5M8
A8Qu6JF+4095G5bCZDDGtQk3/LI8PG5yTP+FGQPO667I28EDbPPvXLeCvusDtQU1n7jXCa+VvHFs
s6gNwNLm1237l/KCQFL6coJ4ri80nVj8gnMD8neat5juywhQSAguQTM08B2IrkAtLb1GbmtfU8LB
TPjrg5+rFhfRpopVehIGf6UxqKubYiXvOUpzabOv66l07vxtgDNiwZsBk8c4jZ8pwff9JhGUPMdV
mpjYDDXGfkTQZsrHt0Q55vuV8sDpllWioP0n+qRKsX84vi7IzdE5uq2WkWA8U1zhr7XHahcCMiSG
O9JAFh90Lv7hZhfOh6R90LFoOfi9oXgPLPQEDlf+TYRxSrr8+oofvkhOzacQy8Q86c9CjvXJnD7x
MiVeUVhNWc+mzbu7yX9QpdXILC0W1JB6Ptpw0EO1Y2a1T8kwgHRaJMDUsc8n0M4ZeKUAvM7wKmPB
eLnznT9eLRHyadcKZR406JBT+BFIK3R65csjHN8TReA41EymVKkVAD8Pqtr0FcUnjkpaiQ6BXeyp
hSyObfcriGRleRrm8ZxCvdZg+pPxe5cLJSEPO9W3Hld9EVBqvzbgkgLhvHnX3RFkgSR9Ss/47RXZ
nRLxs/aOYfDf13Fxe8MmR9c/OgYvpDb2B0HicuXcNAumeC/6TZT5jBMyIeWT8m0uTd1Ejlj9lN+t
cLrVNO/fCr1ln7VswuxMelrYh4gudF8IX0yLDFGNHtA5S7moRkoQlsbB3E5cG4v+PaMd7bLOvz2j
F2JHasX79wj6lMvZKAO6WBf38IzE81csEmaIG4FJT8UIB+3UfOpNCzSG5bUahXX+ojS6ltEwMlHa
7QAYoWZjOep1z2DQvu9Y7Dxd4hgyONqyd9HssweoQ7fNGi4wYeo5eTaQLfPJdC/y6zOpSQXQCuTh
3e/T/WMw8cc/gamq0dW/1X7YxfpzCr9N0/yQ7fA6+ZQ7VucUMSiROg7aSvnA9grqfbZSMEozNlYb
8G9yEZqEbwYq9uZMzw7eLFJSbTmTRF9+3I++BZy++GDfxWXLN5OD8adk5mpsjv6HG0f3fR7zBTDP
Jmi0wRbcUSt8bVPUJESEgNQbHs8RD9rx7PLyyrvmZYbyD+UObw/Pw2WqbORhKHkN370aWHWX9mTp
Wd6sQBXI3DvuvUdoO4ngyanoLSZh04uZyTCgU5MMszucnbnp5ANZo3vy1v1WuXgUlbpD0avFHJX+
ZY2fa9LxT4syZmAkKnLAEtBc1F9qpewU6/lPtkT31HFeHt/0U32ubIcedEXhZ2NFLdIx7gOMboAa
rHmZTKmmcDTtNvlwhGsep1MqZpPGwWXf3Wwx1yZzV/kIH/j9Ih8RQv+kZB13p+ox5a92MMycEAVM
dlXePaBq9xDbXF6aZTUJlO7E7QEIorQivu7mtv+0nppn1lHoXt1I+iL8Nzf7rxYFGybu96C7Htio
Q9aUBlmAdl0vc78IbRBQX3WKxmoD+FpNiBnqVkimmK/DhiI7x0w/mfN34BKM066JQ5PZtRrEtXyf
OAS0mzQ2ASeieB8MRUGHFnlkaEa5YzB2EK+poJBj08hzp/nELqgi4Zb7+l37VyxDPzBhUpUXdJJm
I5+3P/615u+TgK5R3WFXBEgHxed7FgLg+35/Vkr1MUSahhvYgPT8MmGVyoRC+beruazCYfwlGLZx
yrlCweHzXaH6c6Wx9N1R5SCCHHBh75fnzfp44irUpZ0JzpBvL+LVaziavrapFBAR3b2bCOaCiLcZ
mt4KCLb7VHLRS7cOsT4h4KRoRxPtlgCRzx8Oz1fFI/uqjtQAWIcvfZWrFTEk27DmM09zHJksYv7Q
ch/ePFucAGJ6AdKI/k4Wr9Vaa7XbBdf8TWZAQE5p4Wet4Up/1GvQg88FNKt8J3Url2CD35qaUgBJ
VT+E9jPbNum3Oye/B/TQXXinRESL3gAloBR0OHfGyu/VhJK4M7F3mBaDea1oKAiQKzljQkx1ohWW
YwIKcyVKI/LtLQhi/zEwR5y5zFK3rXze9WNNoS9jz6r6gjLbmIpwtx5+UpZ+ePIV0L3YmOhNjcdx
RPy1ADDyex2+jtvdSHBONpWk4eSgPosBJfrestJfUfkdZpXKRE5fyWtp/3OXtcrbrnoJLQLa74CZ
GZ6xTK+m+HR6+0TJKa8sSLoLDTc/683yX1ta4JA0RmjrGqYa/Ql/VUyrN1UF4Sr/K9oMTnyd44f+
N9aOlY9PJk4vRbh57coikt8pYE9lfQtKHkbwiUFgyNznJ6FSjlcHHMK1QFPvu6fJduPYYUJC2CPN
dfRkTlyFRjEM78GIBZRelQVgBIcU8R3xnNc0BoOawVv8nZuzf1dp/c1gx4GVENIAiMvdiz0IaW39
Oq89dSWr4spEGX8sLAfEGktAGZ9Blj52HMetJiMWaRaGX4CnjwPVTTG9Th+3vegRH/QvDmWmJhAG
UuBPOFDTBPf4K1WHzWHaRFAMUc7DZ6ynyutL59Dxx5U3Dy5RMf4BWrXzbp9PaE714qpVNdwZ2iLR
IrNGve5MPLPeKGqt95bL0MOW+Mwah+24WjfU3XoGOia+p82lo0vMuH8xvZTgnh4dZRj88bnZO+cy
LphBNZ6CA+qZSQfW8Rr6kM23K5uJGGUhGkS6W+sMOzhGRhOTPJrEvcViGtycLimQJVzM80BgGMMv
fzozv1EPO1NkIAHFHNHTq3N2bBu96keTSGd0ypQjNcuZqmVy/C+xwL1SQ0Goxl8Ks3Yg2pC8zEMw
1AuqRyHSBj2GSlSdHk+ccyYr6RRsnqo6sb0iHAGqPTIzc8Bv5hndU4r+AGA4PqJb6Sp6PSq8juAU
GNW69iuT86Lbt9ha64y9U4X6gHs3lxTEhxQV0SuZaXdanGHRvqf7F5oZYsPMgxVw15ZS8BQtxG+X
SGu+e4iJhEY7sGH2ilu024OWda6DgDxYjBwtuUXgz/DM/wwFEoSwTuz3viG8IoL9aCDt6VM3efDR
9GyZJu2RCQ7NKxUYFOs3Neg2wLfzFG4Mf1OIrzESTIbBi1kS6NCjajejsQCQJOSdEvTCrTAOqmKr
kXE9v+aI0Khm3UwraGCNVCJcFJVD6qiACXFZEuhjZutzrHs3dlQUNbI9hKqLMQR2HtkM5c0iCKgK
CiaPPNatxj0h79+Hr4v4HEBbisWZsN31wCx6+8VnmT0kNptmcdt565NZDVmOOGNIGNTwOV8GJxza
tGjuE/dFSmYuNtid1W7QKtxxn8224nouWwzsyg9gh8zv1zL6Zf0WImWte5Gw9nkNaevf4LJMputk
jpid5ieihQi6CzvE763MyOcLqEOJI+ua4jIJdQqYmEKRgps/Yb2ntlxPmScpsk6VxNp4Yh5vJ7G2
Cy30ZkxMicfiXT9WqCntxapfCcBrDYIdDu3JuM0jWxcicCnsO00oXHb3Y1K9/4RzwjFF33v8KQ9D
oNI3UZml9RQ+zRlqMw/bsU3sTxD6Pus3VMFzMIEe9HoDglxxWLZzOVpKsd6epPBHfLfq0CmVSBa+
Z8kKKufnpI+NfhTNLFpC66QHL3gk4rjOfxICVE3xFA4hbuVCpqb4m8eeM4gT9Vi5TFd/XDgQa7Z6
E5n7D/eDciDbW5B7gL9HHokmlwmB4/WRy47VWsVibzXfgHw1PyRVLtKLOnskkrT+G+S7Cwqf1jCm
CsuizriG0NiS2MG3b7stBVbrHegFQnWNwH9H2NTSOA5PNuY0L31YqFex8AgDmIxTOu30rD4DyGN1
Ye+kyw7Vlwbecd3Tima1IoJumBZ4O0GN8S3RhIdUQLYl57Gznbom7houYxhFvOsrwgqgVTTDgawY
TmzU5FOhNpBF/sulO4TbHuXHB5DMS+uwLBBgnODIg2XUvG54xIgc4PnoEH+9wXyNwMP1Nb1sxjQd
aEMWwCwvw1UE/FqCKIwFuBMSEAxEjnC2k6fsUhpxvxWhSjdoTiW2PezYos1G6xKjA6UlopGsxTQR
yYneY71g9Jvd/BSD6L5fp1wm8FEYMW5HkB/pAW/aBS8TVem8fIhJTlNyvlwEiplSB+FveUzF7RzB
VJYNddwfvPYTSoCNyxNt1zkjPGuDExCiLKFWzhLXIcIL8nrpTkgCIv+45F3RlWq1XWfus7dFRQxc
98xW4PJ5nksRxMU7U/7ciVJI50btZXeNgqY+bGlShxeMOvNcAxLxb/QqvT3FapK70AdgOHV9d8jX
+SvkMUCCOlP5NJ6ej4e64tWnzi1n/KNeFrL3EXaxOmSzqRC652+r3GcO8/OtO7qol6QrfUH3mIwq
hBelnElqfA9pVCX7B/PY+/Fwv/97Q9jgBb2I7jwn73JdGS2lnGYavGxA3UZINsnOw0jwR2iMCk1a
YsHMK7Bin2wFHIafvRmhI0xz2XYGXsN69AGgyH14V7dif+qypLHR1SZG+s9jzDTh9luOoTsVsDqL
RygwHEP35XltBa94b3AFNvJi969NTq7XusBTU3o8cmyQcmNmk72nYdi7o3Q47ZtMnrcKlVB9P97e
bXHzF1JNKQgWlC8Tc5YBzPp8kFQYdnBdW+KVg44UsPjxz/Mm4ZOhhI8KO8+QzDEgWPqpLQtg0Kxx
j5FMrsML4Hv0VAiOAfPow3hhH+c+fygyFyBRcTpHx10UqCGTn1R2prLDHyyIOcxtqEvakFS3P/om
v5RufuD/PuI0UidDzHbRX4pAZecEg+76poPBnRwECJ93pdGs8GUdKNnGkHrXZlGzTSbODwc95v/g
UFkaKh6XqOhTDBg5/xteckffIIFOeG7BYq4aQ5yddhB+MCfjmFToDDc4EnJ/DR83BgFMwT5mUSrt
kIZUbQEkmqwwe6aFVF13glR97olGoni+uwmXOtSiE+Bs63y8ufJYeje9MM80LFJEP2DYZQRlxTld
hjyUmgcjdQHRMnnB+MLv3lsxI3JPEVmTlFElWIv5YtrRZKcmSrZRMm+muR6ZYTmhhD9MzNSq3SVb
YtQOgq3JC8+jOIBunQpxyuNyMuHzR5M6KYzIa4xyfDUxiCoH0PrgNIyoZy5udQ+GANTXusLc2SMS
iwi4T+XhYGyaCZpF/s+fxgdFBTgBX+zCPcQoAW5NO/qxvl3M4JWThvae/ZlWusQn3okLVFnFs2f1
P8t4B063MjM/bs9HpHe1azkR4LUBQEnT3rnDP6ZmnCIXLU2q8ZH2UQD8MRl4ksUa7b0Qrnq9qbRD
bOztDOg12d/KtUzQHFp2PciKnxCHKLb8WsVgisayPZ0r+zpW71i10MBsbCjdA5qpcWhWvbn3WJsE
JoWrfJcFSeEqSGessXJDNYQz4x6io8iYokXhwf6TZZ0/iDuhtBs6N/YlnnUkHoMGgdbPAhDEY91v
c8FK2SCus7dFuhj0JPlhyHYnna8mB+I6IoWVoAtIHH/Pab5l1MkrtcSVQVE+zgUtBUWJNZ/Q5WoW
OXDqtd5aDRJHwYPueoy41aXp045wN5jfsWRJIPkN3JxRR8X2x3O++iAAwehEKvx5mF63C8EgNAd+
0ZPdmnahWS90Kz1Kplmnys5qbHwH8JSuwuU3mH4r2h+weYolSxXE6o3hjDdRaWpur9Dop4O7RO+L
+/96BiP/M3LHX7SAU7xAK5tOmMTHQS+0OzI4rNa/R3ine6kM3vZYRLGBHb4hyLgpJPyuVx6uIdLh
E08YQAhDWofxDrBQig8tGCxpROxGSvyvbljgIzrvgHCodWuhqj8OCUWR270rQ8Q51VQLAE0p6gVz
xqkR268Q22Eow4r7XNr7itsPeLqsmhULKu2gFH/N9UOCTDV5bKP/dv4iLVPHO1ZvvmAAxDVKmpE8
aWj9qnmRDZu/VSNj7/CX4DX6RJgpuhmM9oUCxlPQky82seuVdm5gNW9vNKCmmUHvUemHENvP5mWe
VPhZJZlMr/Pg0WH3oBlgBj7JmFltb7OSh10llQXdS0bL6CV3bDAhmFAEG949QOHCRyDuY7Rs7A0E
QUi2JQsWJhoRumPiVD0gvpLeDKnVVODt3baknMUPcjG4Bad6DbodkGIBafEzKRRtMtNT78ppL6QT
W1OeWDMYFO/nOAiYPlcploMODFvhkwhPnz5dixCnYXJZGEYdrt+2/IwLxezkoLFoNr5nDp4wR3Wz
6pPkZPJoPDnhneqng6SJ0Mzd+JE3A1yBxgDbH3fhsrgZbUyI+fQSr4icBi6+/znZaUnMaw1QpTTG
qZl0C0pR9o8IvjK+JeP9BbvCmaQw3mLhZ1OtquZC/hGTu4Hb1JyZJ5MMMT6JDRqmBlJc2t1Ge/i6
PEVINjzuYnItoKGCOmHGrv7Mu6l+rjpGAeALc35DsWHalkXFTL9+3zqVjSMYM7D1i01FYnWV3XbI
0rA38/9L3KzBnh2vDkleOGlkvyCmkXDDB2Hucp6SFICi8wm0Rw/OoGiTXS+pdJ1lIn30jOTripme
AWhfWsnbT6wGw0dlFY/9javj7Hu9fRt9Cp5mAw+GrSACH/AFkibO6tIYXFpbtZnRq8rx8jNA32WK
owfdDEAoWYf4puh+kg/ku1gtIbTnLAvr06oxzN3mnt45GYAnVYL556PBIicqC1lS1TCou0fSWBgr
BUUg6BCcYfGZeoKiMgd9es27pbA5DfNkgwsR2jrUY3RGrLjiXfkMcoCmtOahI1GpBgIWPwBS7EWX
o0Q8bBrIDNisdbZOK0r23tzbKftC7TbM8EvoUml8MDFn/pyTdc0lmDumrRT0Z0T6XI9PX2esXKXh
c3xhjePyI4AI7MbmpKK0V5DtXZ80ofByUXtKqp9QEz2ouIurBCKcNdRecWm8preE2AvYKLiYGLek
oIf78WID5LF9TdVKwE/nn2mQWTnI5zt1k9gRQ4SNNDeRplgBwY+k5vf/5sSGXMhFF3pE+Olcsy2J
UMH9PFLjBVdWLIj8tf3Nr4NYK1Vp7wbg31XrLkvdu0PV164SG6lMu71DdGOBpH+bZbepcHPYk1b2
tCO6XqRa/VQrxm3CWsknTk5jwgFA6XZivdY5gcycE3oX8ZwvwUlcnpntZYIcG0JAcxai0jWrCAI6
OXmBMrB4t63ZA8Lnw6WkwGOU34oD/9LXNO8tHHJG6mnDhRP5quNOGv0LWkpkZcuA72sXJeshwGHG
D2U2b7jL6/CJIQxZXCtK6pfqqk1z2Zz+LTl8i/sjXbCX+VV3qgxcnimq22i9MBolSNAvWrC7at/4
gGON6DLKmFugkwHR+ftDquGKwPz2p24Kke7bdA1CcP6KVUPTjib2SRmr0RPb8rWJqwxWZXwt43Lw
vOslhYEkzegVZVrCTxvi1qsva36oC7r+im7W7Wej/f8/21FTlfGGjZeFaWI/dYxKoSxUOl9CI7zU
pv52mt0XslaEmSMNzjvCcMtTTQJgZX+aQKup2nxYlz9yWGgrpd7BIaGEThWNha7Nvpr+KMV8ekGk
UsVorYZ+qGE0QlKs4dken1mZX2O2gm/KK/+zpzyLvb7phii31ioWb/wcSEalOheFLX+5LmnIxY+d
U8oJgUfPvQFQhnuEFzqBIeqANeT+PXK6n2DCZL2SZy4sBPw7ZqbVcr3Mld1qHT11os+1/nQePyUq
CGGx6ZLn+XSGpknpYwbfx4c8irUc+6gliWB8dhsslAuPmEGwBAVb+bbO/yYzi2AuqcIiGyyv3cyC
Yx8Ocl++chehLvwZlg89UH465i+qCLGUJw4NCF+Od5Dvvl7c1cQhCkDhFkOPgu/2cP2tlj1ix3jU
orIYd0VRbgTtUopYSoMCv3aRznW/36H9tiDPfxjpJoCKm9JbtZOTFE92R7dVMUCiDmm67t78KNM8
m1jO9g8HYL7+/a+A/4vLyh3Xn8bzeBCNj9H1v/i+Ps5VAa3ckbNin9a6KFDKc9ssNv/PYcHjHIwh
Ik4DYH67nwbvUHKGpFd2ZU6x1NzIts4CSF1bwXHXYfQeGBVpWwI+B+ftXkn4DUnPRq/5F7NL4HYd
4XUip9tybKmBF9W/GyQLaUqxHU51TKyxKaytWksv0/YJ01xERBmFd1iKr2S0lSkySyEAktsFdTB1
TtLr7F1zzQ9o6n8nlNWDxn24yhxiPIZLuKk3CBU0vbRPY0FcDa2ONSTWrUAp2o7GJMeLlk5NtTXL
joGI0HjcRiCIWuQE326m0D+SgVGl3eYKn6jEXnvCx1fOuwr/ySG1qc+a/Og2tLBkzryzEuq0l+dG
rhEpbqC+L15qLOuxsJlrkB/VcXBaMfhEjsYU6vanzCDe9knT1R7giR/nz6+9eRFrKgYkcZlw3D0U
hc8aJMm+17gsME58U5Ln6FXZx5Tce2fwLpWeD+Z1MUZcMi7izDM8aUVipmwEtwjgfcJTQ9BELUxG
LFbfcg7ETM4fvDQre9pJZ2qSbqANQNhCmBt9D+OJZx0c/FPPd8j5Ctw+YfDHNreSlR6nXRuqivc8
e7Ln1UAa4Yi41Km/f/RbNTb/tZqq9qLjIfKGbIOG4RpHbRXZ2SFbDOwMr7QZBPPwHURYZbfx6zcW
fyaobrtibR62ZUTONxZADNYsa638wPkG6ULpbSprbwoMZVekwHAHTvHDCDv9JBIAKhcwCJFwZSiy
drTMZST17sw1poiHYEm/VnOOM1CuZaNOqJOxLGR73QGbZ9B/9rjJrDsTJ3vb2dajKrBN90VSrusu
hauIn1PUboK1IMKK9qycWd//jteKvlBGyDYjXJ07bOeQr7u6m0+YVgCwEuhm5hec2KCnfJizypne
NgqyBuoDyx9KL3J5zy6k8TAYTJj/d+5Ujf5+4GD7asaI5zADNIV7TZjIkllNNDpyAjMS0wJ8w6I1
/m89xtyKYeqHhYvWJtHRlqBQU506oqN+Fh5m/UxUKAhwx/E26lLvFvopbcraztnd6Dsv8r6s0XuN
g8AJ0cfnLs1F1d9ivgZieOT6fMnHq+otSeGJm8ftdzAy70bs5zDzHRZRqMfBntOO/GqlHbM25V5C
qPZyiScEsq4Fy+YbM7e8E+S6xM/UCDQupAFT/clwgTqQnfAXhlKmYsagpnz2EqQsmuqBoI2c8wL7
hCTt0POX5lg4rWeExSUu8iSx9xj6Z9AeEGNmSqMzIJNGeJpnq+Qx3VIRrW6adEFm0ILLbLjs0O45
crAXzIwCQwSJOPnE/Ki3+fiJ+YJF19PqA3zaVJCOTXgM5fQJvFjGbPKOH2NvsBZtacIOKfOc4fI+
6lM3ayYCUE66sDzR5PcvxN+dUSjUVjZzQOaKeaFfnLPnQZGXa12dHMrDFLucNfddWq1o0J6fAZvo
tgf1t/h3pAxeAhHBWyA54V9evP/U+rkQJ5YGu2GabtV43qu5Xf88IfJZaXOaOgJtvoW4/cIio0Xk
T/M6/+k6kUNMqnAobOoTUfh6yqHE/MRk6jWLEm12mRCOVQ43FurUGltGROkkX8e89agNm/yV4eYG
Zigv7BDsURFPwiIcI3aExq3iDlHuUXu0P1mYsBOYaPYZeJIimEWJayJ52692q85Q6xGBk0+8Wbin
e0d9hmVRa5YLyiGa5X4vhkFb6xA9cvzXtobKMTIkIX1diC4WrzkV0mrPArWjrnQbJ+CBP0Bafaj6
k724DTV1yvloxERM0BrW6k0I8usMvknBvl+f5rXRR/BNpB/BLXOQnWdyEfqv8MKcNGKlUA63gCOi
Vbglas9KWpf+/zDNGmqjobn0Tf/sGwLuR1dGcIMUk33JDO0mf2KrRDUYaZFcXM28gX2ebkVDSpxR
QNjl3RxxhorebJ9DIgtk9eeRcqd84kITB1s3V8yo/8RpBPLkyX2uklToFHnd1W1Ba377ez1CXT0D
fi7jUXsv/aTJ5xEcOO8GD5D7p86lZqoAp8ldLhuKVBpuy65e011Km4JgE9WDp/g5RgtKaMIvmZ9V
ai7EqiPOpAneQy/giGlP5DPTK6cfJyY+eRrXWN6TEKBKpVngoyNP0kZegDpsy7+SoAfz5h5JrrDt
VlWL3kW9P2biVh67DTg+/n8gCBzT2Iz4h7cN/a2xEQ3MoAEtK+EgHRHjuFqfVPWi3sis2t437nDU
nz2mq/mNpblpFcZZZNV1OMfWzvPmrnJ+P8p3Z/n7J/i5kJoKtyd5onQwmqcFKfySduGFFJ+NMME3
DkVEXcaa9SNxRc5NNyYz+YtFrJXxayOuoSEVPRvJSOoy4IpRcXFWqY/zBIct5cHAR59sEDylCCLA
L/fXytCRjfbFP0PHVWm8mkdKzwDmKYM+cTpRAZzAA0TsDPa8bRMzUUSdISkOOGFyau7ybNnhZPxq
UErAJf35JsI6sRFIZYOdzAhJML86mcCAN5no3cwVDC/A88p9cUHLKvdCt8gFVkDXQIftZzY/qG7S
V/6PqNMhu9OFbMZ/S+o3Hz34o3nJNhP9jL0yNMuFyEG2nVpy44lEqrDC3kgfgJmYtHpfRANffrdW
N2YUmEC3JOdgiFM6MYPVXWtM23GkKKqNO5KfdFpI7XC+gStZ8fWCSrrqR7W0GyoaHr1yC7xDl9Mg
qDc0YIpEPX4Rnd+O+JjuCjyKmIjxoqdIWiV2cA47cV7D393cnwcZVj24IrrKNgnuuwfXIScZnE/n
RjkZUjc0kvuPE55E5i8nyhg00MmzOWGpPMVvn9QFQnXQn1hk2Mf7v8Raexc5TO/1nnvWs3q6YDmc
KYuCTmTSUDgQxtuYkw7dKuYpvt/dpy9ESRIxPtrtqNaqex3WcWTkqzGRgN0PK/+wY45nyw2IQ1Ev
DUk0FdE/FHEATXeg+EMp24zFPdtfQB5HWyRNOOK+2RzgHP90E3BlC9rHO2AkIeaXnVBmTdsIj6Zo
AuioIy6ji35xr8H8NVdEs2/BLymjSrZMcR4dM64+mJ85M79QuB4VbnscBMBdHz3EmQKjNjxkKWtq
x3BkfMfQL1ua5qvbvCNHeXxHQn1OMCCSNjU8cwfq3FGotQcMGx5RBL8rXrfuGZLI6ha7ezXS63QZ
nCUFTEcUtiHiYDa+fkjzs5ELUmTHcMvSBoQcx2VX8LLX7E0Mlo1WxkhON5LJgyJGWUt2iz3p7eDX
3FWvuEi1hLSKu/xRENtdTIzfX8He5tm81/riiSxMXLUk+dO8PVCu/mSqHV5doZ/HdVn8i/OCV5A2
oI/Txb/cDf8IynjSIaobTpO5eZ8xx6IM9cfR+HRKeAfEt4ccjbnSkOiSzk7xhna2uWrtUJamqjXs
feRuPjLzIdHCSFEfG84gfggPPv1AU3fbvN/F6+r/uw+bZ5F6rYJ5nSTNeRBhXSzzRwD3YWj6q7/S
Ow/t8yzvaoJnx1PzcOP9bo8JPUJbvYMfhj7EWwdeuw0s5okx39wI27ZebM6R1qCIPXsOF64vcfj8
i2jgY24aMfVEN7ZRsLT/poL4+sU1T5F4jtf1WVJic4b1YbXujeVT1YSoVHgKiVj1VMtpK+r+M9KD
ZE47Tnbu4K/gtTkF4cOWA43wUNeEfHp3LpD680rgLjxyfYkAT5SI9gVYCockSrFdv+HuOGZcCIBb
KZGhLa03dKMrn14z//wJ2pK3oH9cZmPBysbPT15Sy2Fmmjau0XoN98fJJrvVamg/cK0hvit9Oem8
u027mlaFTylaOHzpaXiocHw/Z6gfg73QSDFmdyw7bIZVL6S68tM0z69d1GDEjJmTZxtN9HPyBa6s
ZTJt0NhtR1VqS0SuqxqZaHGXAgwW8gytGkt6WIq0GBYTTCIfa1GIWAQ7P0Oi1z5/Pj1xFfZT7yvW
e8pMw6fC27O1ryhQoXjTTp4KSO9RLURVvQGl9blcZwAOuszR+Dhk2fELw+Q2F6F0HA676JUu3WQI
9Dj7lsp+sRki8Dvw4Qfa1CL9dV8pPypkuqKGk6MhEJmcwnF9rEeD5iPavoM6Ts+Xjs+stCV4gGt2
tJ4edOtb4NTIhTGP25Rl3xR1P57LvxVl/nLxsGLw2eyXxpd2A91tb2XDleMgRAEh6Ku6GC9VOayE
YL+H2KmXHFNZD3S7bg0vXwK5zTHUN2waxE+cpw8+ha0xN/RmLBZ6jAOuyq4TfCn9lz2gwTtbc2vF
6bzM3MnynHo7UkBLbibpGMR0OD9wkSivVA3CQARqnQd8gBdMkUGIHfLiMfCXFimE0eGnApmhs853
CHfY1f7I0GZdIeKXSezj/zDApzfoiJwu4jQ5jwPptJlh90iUuYiu7Ly24UzjxktXz61Vy05L8ZWO
ophk+HUn87CRitRQugnKS8aOOozqrMibiNoRaAgK/cBINZCeDLuoCHMX8/26qgCuhVvHq5C+DQYJ
YqpK6aUXzkFcvfmaH9I8r+pjnex4lP78VQ9NHM/mwMJX/RSAjf6fixxsVznD4fHgE873hNcCxFs6
JStNWYTF3x/nfZ600FSdCOXaM1NrkcUT1MIcr8qMtz4f6zTkz4VlQ+riadgwg12tVe2x+JK0ZL6T
6KEn7VlfUTGxKsK5mRPOF+sSgvSF9bzBVHN/yAnjdKW7QRTWkHrMGqhD9eX3tv3iNGuYFC+YOdug
x+vbDOwpONbWWuv0FzbSWuDDWidm8y7j+ddIi0hNF59bA+QCZj1ACv+AP/I5ITVRMG213evymoSC
CRG27N+b0Pb6DSJ4K/1ayBkSjp7k85g43r9m4DnFtLSuHYbc5OerANg4xeN6OM5yCt4jroA6Pybl
qZEG2W/BoaS0QnT/LNh5cIC0j+8LHuh0kJEx3f/P0wTOrd27jk7+eGP/Bbzj7aQFoNLWtOdfVZ7V
1+fxo3HDCRshOuG3LYTniQ3EsDlNuvEvzg3ItICjw7k85D2PmFDseA2KCA5VWVWnzz5bqyPeB8qk
f39J7ycT1yBoSDDZEBpASkjOgxrGIias6c63p2/jXteXC2hz3GSMe1BN1TsLSZlA/EmMeVPrj+kn
uPTMKB8Nhv1HlXfISpqhBSykZLW+7gsb7+zJXNG6DyTTGxCAqE6SppWgtKE4Z1X9VN9jW4mY7w94
aN4OqxwCoP66FvKsnHayZ2UaB556t96oit3CMG+01v75Dn2Eecn2kjk/ZqVV3aQWY6TA/m0Gl8EC
mYxN3Z+Pi4z0M9pBDfiIL6sdH9uzct16YzodGKT3eP+Vtq4GGzZgOPmwWUjt0SePIOXnBqgTPvYA
9oAUnQUTue/qcadpicWBavI67SgZ4aSsEeYd3lP5oWLCuXlH5ni7SMMNVtBCo0PpOdxCbxEF2ca8
3vIKm4dc43dG1o6S+xiUDPQ2t8ydgra+FBNJBxHWl4eUcyFyRkiM80xMl2y3bmcqCJe++1J1OUDA
BkQOIOSqsjsEf95RUu9ZPdStYKEyxut83BcqIt6sCcJ4D+fFnx7laq7EwN+95elE5fV9aInh4zw7
PLN7G3TRemGuES8Y4vyVGsfFjvaRGofQLz5FZEu57LOamvaRve8Re2uL0asO69OzzS1BjUsU5bWa
pEHtROyQi0Oy+rJ7li24Sb/4p1RyDGMWvbr422VV9sQXx1/fz0qGfwn9uHKBnMP0AhU3SF0shq0J
0WJBY8C3dhsqyXEv96+MYO5cI93uC1lLPmRaYXXB4ynGBIyn3qujh95qJeiMKNQAwspKU9adc6iA
/xKng/IMW/9ihu0hYqvYpFiYpznfMuxCB49tx8aosdt2XXmLkCH+capptLvUpT5Z8etF2SsJe4H6
OFuDyWUx2S6TMku3V8EIslBXwNyjI1bGIJuDAgs29q4NiBXAcVE3a8UlqHOcNR723rEaQomXJKEG
g7KpfQCl3733aqYGifM91sTj51AWRG2kxPe8JTvbBY+gUjjPwD0S943b8VQ1XHVHEu4kGu98/rNb
Rv7gUXpqxUKinQYTzTgmYW+URDN+fGJpCWuPbnZCGeQJZ63nlvP7WGBKVAHYKKCcWL+UTRxikcUu
OJ9lzBtt/AC03EjAPO0DuPQ7NiSuDPNMJGrqLa+TPZApTlhncZqHRUprF/iNsLsN4olTplZBHsTa
5pbxgP35CR9Qo3m6KdL6uZkqa7vcY/rnHuK8CUT7BJsz4NH19ByqYYfsO3uWZe3mD+8n7LxCmp+v
jAjH+lHLNOj8TfYYhiA5KrAd5S52EPF9L2KAuFGFZx1s8Xo9r1KKDKm04NxMoMlatT24tqEKAXNm
/PLZVp3tJtoZ0XXi78zta4TnhLbyAWBFLAvejBtwyR3k2V2wqDHxk9WiQ630DgQEMjYl3JmdniMr
UZOfrn3FXi9F/ciCxvdnMuLnsRMgK0D45D7c7/FX+NaTZnkb2NDrrW5N4YBxI9Atl8lOROvwcVHD
PRo5sd7VJOSh4F9kLi0znUJ+BPZgmLql7eSG6vHFtiec7uIyHdO1QLjIVAs7nOirDjaH2BObWzyA
vF/zlVyqT1be24CDLkUtMLIGrS4HAsVXVEIqW0VSfsQz+IPRrndhUd5ui1/XYJzdav34QfCld6+Q
OLuJS0xhOwlNyBffzUj9NUNBG4dgaxZzam6+e+d4FA8E4nypJz4W6fuz42tnOtE1q0YqE74ywl0L
/ktCDzHpPBx416taV4iY+Iq1SK8CMOfBkSlvsw/mh5fiWDWEQ/NrD9HCVto68FmJeXFf7IxPzyst
6et/jzGJkZRwQGs2wkAh3vYZM4PCTp7VBzX8ZRTXeQ8dLRkcaeMDu3cE9MXN2T1YENXJsYRq2E0e
qCO0wG1lZZ44Kz8yL/CYLGQ0vnYq8yvJGbKTKXO8ucmdzyMPX4pweX+kM+sYMiNmLJ6QIwAeOqxH
ffBaVc66KFu29Y+K3w14Vgo3gmRN0kaO79G+c/l0hVM3P2uHIISvGkoJn0VSVLYrUPndXiX8smM3
OneXlUyBjfPmXrBfDmGA2+6JToN80OiBTu8h/wu6XLgqlxlgu7E07IUOH48g0U6qNLa8ObPwbzta
ZlTZi+8FlzjFp9y0Pur39Ec3QAfoyHyavu8Zp2A/m3x+zU3yF/HZAPyetbUfe5SqqF3UJJNRjAYF
kD9y08QVY1Q7SERz6FKgeLFyMnu0Eu3TbLSQwdEnGZ69WNiq8Lb3xdk4JMWCzkV/ucRM7Jya/dB5
B+Vfhy6y7tbT6wpxMwx0BBMR0h7ElRQT6/ckDmOOaMiBCVYSZbFFjI1LmmuNroqEqeQtbIiZBbhr
XRasQTHEQtXuPfA3I2ZnfqUprVt6GUhCUosUH0fhzGB6exOpZfsa6BH2uAkyv4NyaOokhkfrvOTU
s5GM/y7afIXCwHGDEKMI169cHv5YWHqXOym16F+jbCltrJ4Ff3p0fcqnczAkXMLh0UFITBaNShz6
tGLNp1praGJ8qUAPlcGMdfO1fLCjpxmKm2SAxX/83aVXrW9ILz3y+jqdtQiyASz3fQ1mTDOY6EYl
cZancmLsadY6xkQJPHP6Fxl3WZGCOG7WGjQRj+h1l+EtTSWidSeOVUnKFaHK/16xBlsbv/zBb9+G
JALJY25kmJiILUYR/fUCUeEIhv5Z2JZQAtMZQ1qKPNWmb7PlRy9zWFQxXIEL6EhN9OUCquGMgfD3
x5xC/fjjpCYbPBCLdmrQCaAkPT3BiHudX1Ocdp9wSt6TUIR2sSxf518hupZk02/MclghKV5gtaqM
AjCCrZQNWPtRkZMPVI9h2shK5abraDhI+CrtiUXJETXOUAjE1096B+beQaecajr/6paIoS4u2cRS
2B0sV4MuzEycXqhjVJbY0ltrU660s1fDyTI87mtlWset3wM+XCaETimSg5K7pHXJzrE2sZsXYSlv
g5UOKnkfEc74THsJ64mppaudJf0Vm+oqD2OmwE+SAB46Uswul7/QNurOGrTowHfbREVFtsMmgJhS
uCyfII3MtwB+zJqGW8ZL0mwnVCa/jBkBC6SiX2xJHgiJIVLofbar6P48cX61G1nD5fO1tromy4b9
VZ7AbDHNx48aYnnfQqt/Sim3jNgok0lPohiobLvSZ+hTQDHrKVSVCx8vp8CLhxucJMZxRd8Fx6Zg
9Rzuj93YrbGlJxFeT+3l+YTXlAg/wzDC7zE0KYoolFeq/3gyfH0rDU0SVo2ENUw42Bjj2xaORw/G
ne1grISDnUGc+ylEa+4EBkk5gD4/WS+TerIbLKMkbvOEC4OD59J3LDp8qSegVsjvpGVcBc86BfMn
RUm/KHn9lGV69JohzG8zsT9mgkeqCoYwddk1U0TuEj3nj78sd9F93ak2qbcy9bUXXd/8PTocl4VC
kvYXs3sFZRExMuMUGO9Hg3U7cJYmJXAoI7TZ35Mq7VAo9GfnwX6EjZNiCJb6s121YzkyG1GelMPT
5xQO75N8boM8HZU/nvHSm6nFCNlZQ3qBiaz+EepKNTMcaqlUo70xp4paEXRnlUEN1daadEzLRLI6
1xojT7QbIk3cbzjbECgVibyS8/UVli/O+qE/3c14t+83YnBYvybkM3kmaZSJDUkMhgC3493KY/AA
9iij+nsDPbjZnds05WoqDYBvV3nvwIVFSv9p+QqhPhD5PYgyc239844WuEqGlgRGEOZNePP2dWni
wl762jCOW51VO4dc7p0P71rA1oDgu35h7o0yp2R6bypFmKQWpdm5oVFYWtQuStIUSaEoL46iCM4O
n53vjB2EWJ+QJxDLI+ifREKzgp/JFe0LyTDp/9Ka2U2bJiiHJ34p1HVvUbqAL22wY9FDxYd/uJWu
sVFmIsjC9vQnxc+ucGrs82uPvEpWavqbK3PEGYFNdcVQyqqeEXgvb965nFAVMBt0/ah5CQE9zp7M
bhNeOOwDOjMSNlY9afRlUsNdtMZL/LERRX+Ob71KaV0MFD6vGR1XlUlV83UwXG35iRCA011eZSZb
+WE605khxyx6ys3iG9l9IJQjWQnOWPhXcXUCuupiIUoHveIDgx96RptAEHij+HKH6XTvJo3GBBlu
suANIbTD1MzeHA0UTXBQakSGE8u/o7zckasuMw8jeeLewnSCNiAhnrgTDJfigKQ8cexjh0ltnLSF
anZNVRHD7EM0k4LZPSX1KFg4Yxf0B2Qk5CyTi+fm5+lMSw+iMxzAApnc47fjp0TMC6GNPnx3+78M
xFnXVzG36AofjUSBB0Vt2XZME8rjn/t3fjX2m64mEB1jw8DoU88shzEr0oEHqCsAzZegccTgstWC
d/Zb076QyvlKoiuxQUcZKIGpfR9XcfLCo0jQbf50oSXxklpsTfp99/u65HDYAV4K68p1edUaJ32n
jTz1aRZfEcNEGF3d4o3VLeIkIgYtJ1phl1kkn9CiAxdWjAjFggb8WmILfxyuVPfSQg/uEzoePe5Q
UD6DNjdDoKcjdm6jK5ngoERDCstjzy7g1CpLBHnEM1LsljdRts7xpsYB59OlwHAcENLxI1Onsogt
ISH6/a7GsK+UIP+6YKYiNu/TWcYgnAxel/4fx9iCIz84miMinmvVzyegTMzWdavXAd2JI0QSLMD/
5CXeoqc5iRwkaIa/B/9IogZbS6jvbmqqLFYZ+d1EpgDnmegNluSXbJJh6oQ/Ms56fm8Ywzrx4BMW
ODULA9yixgWnu0C3Cwvn/tYQ3DS+yYcHwO+Z/IKPRe25pJRflLhA35vFFvfqgMqXpAGMUXpg8dX/
a7Spik8K5h2BXrlNS6pQRuCxpotZnVt0pHYjf4mCFU2ZpBCU/C6T4LnV55fJcHBiJci/Jy5bBXlz
nC5sHMdzs+urcqqwD8uP4E0jdda43Dws0SMscyyooYFMwRW2TtQn1BVEMnb6W9+isOp4rnnGlPoT
Rj5x+fEB+mBmGHbggzC+mAZ8SEjIM7MLfxr843ZfsOgZZ2Wq+r65cGIagKA+P7ELf9+YxDWn72jI
oE7k9jVK3F+grsd/hICZaOrkq0kD+nxcz3nPr/0j26s+MbLqz5lg2kqK8S7rHgWfgbCP/FHKe1G6
AUtroMJubqKOGfE+XyHb880GOPJ69yrhwW1Ck8A837T2K1Lf43oFPKtkZUWYNdPOCUTLKW0PTjuf
cfea6/CDe373yVUKgmUXo9oMNYpp+RaVaqSYnidu9nUUbjF7+2M4fV9vv4A0yKFQ8iBpRYh47u/n
24Hthw1vS+jvuW0LlcjYRDoWtqzlaACxLr0O8mPzurjH1BMozv4lufjU5S0GHmsSXXWISX8+aoYH
Nw33M15/ciKLYfcc8Wp6kHA6TTr/4eUPqDwUjhvO8ZpAufTvdqjgwFd6CtQ9apT7pmm2RcQVHkx/
UhqismSRB6gKPsZgvk0GsMUMy0cI+s0UxGUltleGTzBMXrN2lOE1qpP6o9n/yPMp938X516j2ldx
Ym7cdCnpThmeqDMT8NcUP3IZfgs2b4WqOdFJHeFNZbvnZ5bO6+xXT7Ut5tJsbDXXc6k2XcgmRdy7
XdnLEss38U7zec0DhEKpr51xCFwtVJr8q4loXR1UBYWFPL42lQFIMTtFlDOihH9jTSVGIjF5Qg17
q5F4HREfMQL1mB6g2miDqB2bkNjytT0PkoBPIlZyCE55m2CorSqPOGtWnIE7xzu92hsQkFiVrpMR
58Xqz20rRTEO5iOa0MBQa4odhb1wvTzs6WSlCi4WR1mbl+Sy3vwdFRJ14Xtx8yL0J0PRLRKZrMjf
STNvAmq0K7WPR/I7p+cN3EweSQ8xG9L5ekwrJblhm2NinFoKwsqaw8lkuTalWeoLZBZ5uOAsXBQ5
qcacch9UqxHF9Bd3Jhuz/x36T5r0ZTLROVcihVqdn1pHpipDd/RazZUiWxsptLHvqoFeZbRk8bnO
p6fbTsNrg7jYtlzmLIfsH46Hhr0R1/eXdDMWL0m2xcAN9AVzEwnTY2ex9GRmrd/zOlPQMbIsgCt3
85R2Ncad9c4seFuistZwstLkAO9QYHchLlm9hJVo5peQ55GRXMKJR5iNkXUAhVxllzDOBMp3EVX6
fRjVxixkbUZwBoA2dHde1Vj2gphKlwxCCne6bs9jy3sM+QCg8e8GKWyvs2zW10v7ha1zOR49/hIE
hipPmO78O8vsKtwYlsHgm/8hl3uk3D1aCJJRH/4h+DEcvoeZZAJ0d9pQwyR3gK/jXyn7RKqJt9fC
KH5Kll2j4Y7KQB9ycATS0MVrebm/MhfYLjzudx/jx5XnwHeynByO2NJ/k0lAZwf4zTslcD9yOYWY
5EIKHWpD3q+CDaALXyEKaWtNeHeYaJpxNrcsaKeODMr0YdmhZsJgnpnnYVmcTFOBb5+srI7ReVZx
NBTuOotcfS/kyCQfH+a/XAsXzm9YeWqczUtUtmoAhyh3WeN2edHAxcYbMjr2t3qAeDKUQaGb/NmE
GY5IX35RT7CxLQh8Vcv2LIkm3tIR7gUvcq0P6+PyLjlZetZC+LPe2eSWAXLHgyFLjRxHVqE9P8tn
++BVeER/pu7XRicCcVtMiPb68JnE/0EZooqEeteswwzDPqj7qX8j8eBSObeiSpxOKYr0l7fIZnDs
Ha5R4EsecO6s2xIdHRCZRQHHlM0HIS0YQiXAqmtbnQmkYlWLwqi6Xy+d9Rrvrx+T073Rf5CJzpXO
gaRQzsTlra9O6GPAXi2/iBFv2EwSW5ueDk/ufwbkgT/X3l3QnsAuf+UAgn5MZvdhBjVXduF9HtTN
UuSlik+ixwFxS0/16ray16XIUIWA1wjRgwJsxYWab628KIIYO4FlXh17JuuteqWt43xOM6gZ+Cs2
0MyV0PHz8RG4rxncLTmjBfVDwZ2UFXj9Ef9toXgH1O7TY4S+yuW8F5KmY2lirzL59jzrgDzEtpvg
Bxsh8/VQ8U+Izk4Rs7hcV0yhAJFjBoly3KQF+lbmIVjZVPFrGXp41d9+vCNZsomORuseHSsNmhRC
ozJfNqWRzw/fSaGCUJ5/IZyppBzvCE4pamxLGGQPIM6DFh/ohdZmHBloYq8GuVmBaNCQbKi8/Pgu
m8pJfczhJzIpg8+jV2KtZ0ST4hsIs9NR1rFDIOGWPZgLdhcdWsyFX2Z0czf2gkNZpZ76opp4m1Dv
hz5U5oQeH1F9bSyVgB1spkvzDPQsHRR+ktWBvC089whl/v56YUIN0RKQth7MOAlDQqFrGvTBPdAZ
TpjzzYACkBGjAoEha88mFH+42G/jAWWfwOIgR7HCMPTpLSUPQZHRA/cNyXZlZkzJm9kIerSrzMrO
eq8RFq5II/uBlrz/g7UfPXhOfM7JUM9EztaPaeRTR30e/gDe7UhyAIa2bv/G7hHx3DxUgZ7rQJfc
Lb550tYwkLr/5bPNCbFbiaAhqtPAc3QbZK8QyrX63lzRrpuyoicyVeqmvglYH0Pmvs1TrMTmdc4p
3axOP69qqUmGikxV8gdexKW4DsHuD7ygzSMBGy8ASe5tiNM/bIHu5znFfd0CSQgERektjJntNgRy
BTzoM6OTabK8AszCCK2o6Wh7Hjj2vf5xS4ZFDqsbjwoZ0+b1T0/ab2Y//FDUDv3PO19lZiLeOpI/
pgYcBtoEz/P1Mnq2PnLMuqCTGoIvaXuaCmEdZR+GRGZGIgX7tjOY31wGpdA/tVApQK0s2tw0mApn
PR9kK6rPaRwzRj5/EK7q+u1Me5/rrOXDPM6ywZGQmFqSz4+XO5qCR4Zw6G2byGi0L9gJ8bdPG2nZ
DHburJYTHGl7Jg8O8OsH5L6CFPPDBdRAcwA+al3JKE5TJRwcnmcSbXIiW6fMvNR+Dk93H2JjIm9Y
lZVU6PscpvbRvjT69TkSBUBzK01z5fNSFwNtWQDKQzcPRrGSEy8+9Og5BGpLjB5cZ8s14T2yO8ER
T/9XETcu/1XhBzGleAgNpzCBc1+bYn2C0KHfb0LifrdsV+GFWNeBITHqBdo7iNw8M0EVtqk7LmQi
eEHIQzJZc/Jq7e/79Ge6INwMAoQxRoVyRf2VEFXgPq/pOTQShKy747KuQCI4RlPkKLsr311GD6Ie
0xtcjsPwCX0JYwRa0JXWDH44r56ByVUoH/0cYe0Qi2vk8+lm5iiw0AdqZeMAWtjioOSmkrsE+8iD
/MiHOAuiKs/eRr9plo+PYiCI+AHNMagWowAy2/cV42zLPrAx13tCufCmTb6aP/Om6d7/4C1T+DsU
aJPGiGQ1vULZnlsjYjGkQBEWkQvKT9RLTU4eDz40HeQS+zvNp+r/VBrYBG5208/+PXyCwQsLtO47
CD81fZfQ0dj++CeFCHLewLFnbB5cI2/qh2Zq9hACtapQKu1PC/1xycR9/jRxev9Pl3QHtbcZHRk0
z4dSjAePxDKIIxB1lnIIRSpahqkWXjqtTmlp0dDXZ9YscPQaKB8nMvyDbLoGTFLgZoC5ULDSXzKe
BXcnX0PnALlW4lz8HLlnUoT6mjKSsD4oCSfUk+78X6IatjPZudjm8I9kDjtEB8DToFRCUVBONOoH
fBrKCi7/VRneH9x+l0DYXrzj/L7/+Zh2RW2Ve+RssfmDfrSItfqlXlY1FA1ta628TI0yIois4PWh
AFB9iNk7jXs5FEDI2OMt3T56ZOjRXCZgfuvJhygys0lP2dxT08VlDgKbDD8MZJ77GWXw5cxo/Bbz
7oK4xAsbmCH8baLGuOVl94guCVLOoqlPxEoWuBknZfV2QbIB68i4L1+ZojoI4Mpof9cranIiqfcf
ErOzJKMBvqNAz5el2ng2kJTOg575du3LMyOmp2JHRkLKWGd/ZmQqnTFV9TDUra+MLcnkrnFrHNyX
SqpZefeMmu6lXtxjue1aeNGlYFI4RWSBvwWZ42eCva/oXhPjEucYnyon35hrqBLUkqGoAobdJPL8
swiI4585ul8I7MP4bXSsbhsJ6SPZ5I8RuoyUqsyNF6r1/s72OeL1qdsz8aTGY5k7Z4LcyoLbXKio
3+EKjV506aBoPlbUVdK46wmJ8YSciklm/xgRYLV8Eq4VxdfdovFS1D9VXDpQ+vI/HsVWH53N3IEQ
cuKq4EjXqosLT3AtJzdAWhkhSIsBrBV6wKI4Y8kiWnFNrGOsAGG+Y+JCE+XprVjOJd+jnPJfg07C
NvL/c/1hnreVf7br+nTdMMjZgY2v256gEFT8umudewR3KQ31WMZmt3xXK2yFG7QA4zYLWlyvCwu8
dqr0Xk/jYFzbKYa9tTBV1Mcm116haXzRsH19J4tDLXE1IpMQ+L3BlLvRPtYb/m9vG7T+1vmsBIZ9
QDIsRfzagJpsPHBW6TRidLK1S74emdOp4fKHnzXv3cspkl1y8qdT+WNmr4JDQv6OTBh05ry6kSOY
EQRhdQ8eb0A5bz0gR9zMOD1cpLjqCTWesmeWGtn6oP5j046BFIOPYArq8O4VCD1v9mEDiRpTsPGp
oCMRrATfc2vw7vCLddgO5UYyvRn8SqK9IwixZtHZvUxWVXOhpaDg+bivuSV/Ie84+/IDyMeLcgyJ
WgSHOQtOntjtGsdGwbMIHev68ae01MnLKtSuy+MCfKJry6dABQjq7MpKaBOyawUFBReUOF9EvVZu
ea0gebiII0CwkbQR/rN8B+GSULxhvf/atQpd3PUpQtWU8SeXU7oxDL0irfvpoOYuN0JVYIQbplY0
7x+ZiidTzSeOKqfTsmHusKxRkcDDFbVcFrDdNN+3X/FWpyJo4HM68BQ684ptIWwS2RjDPKTyVMHc
4IzAnBlxDQtLDrbj5X3B/Sc6tHQN8BlTtOi7bYMIVYd53aalfEquFE2bMElbsCRemqlXFdln/D3G
cc4/UWFmYMz+i/Xg+vOrc47E1VuThV9zEaiQUOUoa9Jgvpx0zIfYnEP42epHBf9sCdPt+68CjMTm
63GTw5odT7HOvrEOfhnXnZh4iyzEtMfF1VuCYvMd4DAcyUNAgd2SjcrsgTyOog/F5zwFHPjZ91AK
V2U6sni/7dxm5lRn1bPeHPsQ7ptfA8hbW5oWO2/lhqVvw9Eldh8M3URfB3OQ2xJRlvU+7t3ckRr/
uqowzQW6OhbC7G8taKFwZ7CixHe/9v4Qe54N5ZO6ZG1JX4dYxJNJjWrcqvrfUEszx4cekrrfmDIR
X6wfIaW07tCFtYDwE0Iww0hpD/bovx5dvSUKdnL3kovAhvUh3V4Tp6YgZ31/H2fDiLSaC18YW9U/
zKViDFgOEA8s63+Qd6Do0Ww93vBGyMREp9IY+BNnwPuDYNQUaIDQcF9dyF2wxJkETUNkDtPAc7AF
SzlZTQb7QLvKS2PyoFjuOQv8Q0I8zhx/pf4drro/4hQSlhaCTStz9RWgnsLQlee5OidbrJ7OjlAD
I77P0V8S1Zy9vSqxkaGJyjCIo0an3ICW/z2Wpvzn5pMbaRhjofOW/ah54jnpWrrgo1zPci4AXFGe
iuG/M5ZHJxejQ4qxyzLLKIiVFQIGq0AGv9R/oxYpWRQCv+KieFALUJfxBXDCdCVCXjXd7s7mxWCp
Vq1BBfLpsSoNV5NtFwGbHw0QFMtHTJ4m9r6rmSkaPg1i4sOpFRsFDge58gMMlEUvOp1e1fHiT8zx
f0SzuVJk35xYxZI89rWTc/qkn2R/W+N+J6V1Uw8vAcbpSjcux491KSeQAfhbEFx4saBHG04zJ5Rw
N6NK+6CGFN2RZF+jzY5JpJEXZ90x8jcbA0KMszJa4xzyH1dcoW1j9IaDcwk4PaNU7vSjID8fPbTP
Q/qAOigyDeQ48BqHRbFsIjbqQ9b8GpKk2LMfv7nhta0CYsdwELf/OCmxlNAj19PBMm9H1Nqp+G4n
BTq6C4Zy0bdO5qkx8cc39JuHYKeHV6wu+QyR+Mfl6NwA8qWsBeCsR5zp4f+EOwr/tY6lYIZ2vgBZ
iVQikntrFYbmpWZ3RGFyKwme5gr5r+Dr2eeQXCGpIJ4CaZXwBdxnQC9WXPI3hdAGe47dh76xwPmx
gh1qwh5SZXfH5ek1QLD1p601cGfk5/GAWSxYB8FdgSZH0Ut+OqoVpwmK0Hx94Fp5OFpZpKVQcddv
GPRpF2MYwQceVcebIg3Zc7ICNyY8/YWU8s0fbIFcIcZF0FZ5P22mBFI7uSncgfKD9n8F5PI2pdER
P7ttQH7a5C+0jUfyyx7Jde5TW/N7/G00fMyTj5B9pBhUUkE3Ny3gsX69+sYQ5cjc1JZGTkvIlXGk
e07DKtWf9+SutRzJFPDsrxSxGtfZICu+z9kLlTlsTHaW5jYzJIsB8rRsIzjuXihLHN/h7Le0z3/u
3bKhIo4Xun93mCZ7ESk4pvxwOdS6/nIrSwcTFOxlePY7tnAvK3Tzc49YccXkKuu0+6zwgAH5EdxP
OETAt1iqVIvV8J9zQtE3+modneC9T8r+SXvSDICxVASXUzqmdiREOlqMPdNghQsfCg3e6Fi4c3YH
i0TtfB8paYEaH+hrFa8yGQhzfN0/iMJCQ5nTmcULHNu4s2PtZDqecHG9xpUQeDIvJrz6nzqxslHM
FfeWo0T8KcmcFXfrp5osHWM5P17DRm8+hIHPoF8mSW1b58wDSZi2HCCz9xwP2nLWOgGmEQa3lVAO
vZseGd3V+OXlWYhqegKmQQFJT5/Dwukad7nbAUUz+C65mKu/JMh044OCCZfgAI74njbnu9E8Dyoq
K1J+7KWNVhLYGe4qTfuEzteL9hHpq4OsG9U3pLuo0ogSGcWpO59nr2PiF1TV9bcYHWpBbCd0saY7
HskWHADgn0tjpG+qRG38veW1wdwq7q9OKIzxvbH0tvHVkiPfqBLVxxDpBPLaWifu7aK5X7PtQce6
cqXdXrv89+jsddp+WZF3kjngdw0QhDDOn9abhde/Hr8DF/OYis4yKvmlg6wgGr9EJWjAI1NQxdoU
IGIoBLZdT4dEa8CrhxZvFWaz7CZBifi7bOaq1YvWtMVkMOnCabuu3LpaW83HPHlZ6ERPzQNna4tM
q78fffslJYhDBTQhi1ojlRwh42MaSrAvOPYASesV9qjzrPTgdnI2rjl5HrGIYpHqQVFxOqCcIANe
rNx6m2737EQFuSTBVz8ELm68i7RK/UdCDj3DzDurVJGYj+/IbHlrBU3yNhyK2XKuTh0Bra2Blqwy
T9UMcf8xqc+ucON/F6haQxvu04FrU5PmkFQZ43UJS3Sc9dUENpR4RwXpHXY5hF5GJd/J/8XUsUct
/ouy7fNEkSxN7+YE3lwCrDi3wLpBTDVDs7b8Ppc62ZsiVOKefCw0aKnj8T+JZedKEVB3jy7YabUL
UHPiXqU+9I7QF7B6haHEzc8MMrXe/FFmOvSz30ZtD8PcT4Lv13PuWK5/zk0DuEeNh2WmsKJfv2Vj
LxVjJQKX6nFeW+BqJNtkSCA2wM8tJWThv73wWGObRMMOqpZuTAmSh2Y946Bukhrq52ZLzS2Favdr
vBP5CnSbH+lo8vNmvhhzC58y5fS7F2x+FwEtAtzNwjwUgC9aertakK1XEJXayPpsC0M/M0RonnH5
3i0ra6siwbI6TriW0mLSc87YmrCyiRIy8NLtgzfG8wyrcp7gfPDyPCsTRPWYFu17AEsGpVQ3I/DD
NkrAZ3gmmmJQEpdjOPslLm1oAcE4XbzaZN65Kk6jtgiXTKiLMms4Dh7qBkm6Z2koG5Os7G2koIOi
9MPod/yKnfMwNlokH+PthCvfjjqre7dA/vG2L6rfiNuCl+5c+t0AUYK2qbpHJTdoEK8qb1xNI6W1
PfVCRXEswHMC1/eP/rJKfi2iXzEFqlLAyDEk6aqeahmOQec+cW1TjepUAizIM9xqIYXkYXHiYT7Q
wuf+DyUemXyZpnKBhz18rQNu2e/+Skf8yZePDEFqdxm9KaJHE84bnNqFLUrLeJPnh4PtRZOvm4B5
ywgV/99qOb/SyLqFf5lTapIcwg2PZyIoZPMo/kehnVeu7uyWny8Mv5mMMSLyCbEbW02Wjk8bqkSO
5ukZmvMbs5XZ0fq+qGFsV/73Pu0UM3ESrS59bqjX90EgBpYQgGmBCY2+HAigurIemftmk1kdsGEV
e9DuBsi0FxDrsPL2xtObM0HlKgYnZwhW1mk0cOog/s/z9dn7wRhrLGxnEbA2p64eVX4Y06b2TIwY
k29Ku9vhmjL+J4CsyxEV7+GAWUa7Xu3os3lrwD3rnXri+YAO/7qMguHEwi0ARTWEKFP2lM5h6nb7
FDZSaeL7jtoGhQi45yiieMsakdDXCXxwgbl+TaWGyqyMO7l0Nf0dIEk4C4Z5xTeuYWg5RcXGKzFz
ti9xU6rBowL+Xfq2syHABS8Wz71/CDIYUcW0oUqfJDJkYpvr9LhzMIjufkJU0JkSwUSnZop9V4GE
uqWk+SzRsd+lpOiZX3M6ORvNigSHbPGKhNAIIkK/MKBUsmT0PrgPvlxczIBYOmDzyfG1k11ghaPG
pLnAryIAjbU1AvhFH03njYf2wKYTARhoD+mew6WDDETSvDfpgcSt8Stc+AysNIP9Kr+FMC8mPac8
1YBtfeCSljNPhGNVkLhg85KHGEp/IwBHpHdut8Yi4MjGKw9RDhinUGZg5cZY0sVp8+aWsdXZtqWf
/Coazw0oMSA6bJsN73PfWHzSZ4g8Aq8G3bV8YqfAjunxR8E2keYWd/3NyN9niKwMJKBi+iq02EbU
JNzngaD9MGBWQNXGTSx8el4lSCV6UVv+cg4eoL2u5Y/8EvDivXrgJ8v1q2CNxBkFmoOkajJm097i
lDmo+nFmc1TvqONq447atebDNwGWyxmGjT4DccCtsCbRqeeNxGtup6mG39KKSgTYx3/mqpoyFslc
sc0TZnCRHpnCyewZXkfoy0+JO6D+to0z47hJg3rO1lktSe0oUCOay7DrsqpRXxeeKe8JWz0UPOxJ
d21+IwBgFRTi1TMOKdMBMM2jnGFHikPL4tteI+umDW08KSOoSBsbug6BgY+C+byHQtOVNC1dWbIm
ZQkYDBCvdUtB96rpP7OXypPrwBwvSkYxfSa0ff2hXxtRYZ/nLTUq/q3Nc54x2gzeBiw0CZyDMFLc
IGektxZtBq7NR9FLG4OuZpPHC1uMzgeb3rb/OVLezcPu/HkXv4ciV89aNZrY/AtWgerET2cLX5Xj
V40CJsRwUvt7eq1KZS1GNfi7NXW1SWrnVs7vTGWMuufIyzcAkAdmSYpFTo2RgZtlpBIWUN3itJei
lX2ilE7epQ7Hascm5cQEs9VGzHDH4vzJWPplqUncPALtLgV+exrCvNvEqUnxFjkVYNfV35ny4HF6
GpO0xSqpq3D2BCtMsg9uYlq5AFHYK86pN2wxGalniL0vhXb0bVe3/3zFht5IZWM4vq3uxWrL5lwB
EaCCq7+nbseYMVVZYY2+Y4PRs5+spK8gk4d5hnRCrPa4cEMqvpeH4hSzmSvGbOOcBMLGLj99otvk
8mLy7to2pRt21VOhcmZoKGuprTDFBocjbLVc/LJxaBTsOXD5XlhtkPxwPfJO8CWW8gQdPCPBfW60
L9A+GiyfB8uuePSs9oVYQLkIrMBTbfOFfTT+ua2/AIuNL3pczJkgk+OyEbNXNDn0QXLmdxxKfoJR
eTaOmNwewcQnWe7TB0DcohgGBD6zy/K55/nCThKsEbBbFFiOJWWJgM2zB3dlKvSdztZARurw40hB
Av6cQ9B4nj1MXBn1KJ/Dq4NysZw1Yjb3WQfIg0BEORC2Lbq8Cv0wDF1OGwDC6L1PmNhO1wzz3pAf
JvhgxBFnFnbAwTjOWept827SQ1yO37HyhOTGeAoS4fqyXyQvCEdhxX5BS4DQrGi73pT2GbDSjkQb
Wb8/KHO4ckoayDjXN6hSvekpigklatg8FNsByRwmkVBHJyw61qEKni65Q8T20CEyxOqSj6ScuOyo
WoMG228ayF5GONUDG90yI2utGQnQ+UUDRRAU9Jm2u4UL7yzmlS5I3lUT1/4GNJzIoNe2iugjftlc
tx3vLos4auONL1yEMNj32b1k6/GHcdo7GyRV80RZpg5ak7HN9IbY0n7R3JTKufK5SCg10+BTWZyL
2nXMsoWDHsyRUmX2l3f4LBLUvYu1akWa2XdTJs4wzWvBHe/OHVoMfkdc9PfufF1TNLPISCuNq8/r
VtdtYBALCZlm/nvtlOE0piPftAb55WDz1g7tDWvCAo1uqTQnokOPqnYXCq6JFTBB3j5Sx6g82f9T
i9H/0wmIDq1/LfYmhaKi9NDzF4/o7Z3I++FiYMVmsoZioWUNKRJz+hZ2+aMzEMioGWpUC/V+uZpo
l8zdaZewU3Bp9/YTtWl/4c0yj6Xu7y8NXCiSQ/+oCfk/MarQnTSSoZmXrl0Wa94QVzArg8MGSBam
2I8eM6pXpkADFlqG7z++SCTAKDvLYb9XsNBq+DRuHTVnya2yEe1HLuUnDtJZ9sCuAWdODNPc6G9w
U6RXskfMVsJ2SVnrJF4fjni0YSAKmMCq4SfhEKGmILSOVN/denoPlIW3ae1xQ1IXaBCvEynUIp34
LAu5ayTNa0budAPEeV5BV1Z6QVzWy5kaBt0zX4rT1h8/NOrBtxUKxxLZH/faunHp3P+0GyxFZySP
UcQ9rR920Y7LQKRZnhaOHzC7NwaodOvrQY3rWqTVLHTi4W9kYxh2SN7snwe3OR60bOhFCCwc3r9i
mMyrkH4T/PaeYw+33JtARyFT2n56/zYysyxWXwgXLxCxAqN9YGWakh7KDLy1x9bs0WgIF22xyXM0
ICHmg4xh2VRQ3BUQmA6D+/+2Y5hfQ3y84cxZtanddiMOCMX3n8padOTsEl/AK/QiuYUHyFOsEBfz
UjwPmBb+QtIqqdENM1oiecQtPNAXgvTHvGVcZAu36BBoWqwQzuP9O0T00lymzSVyIoXrHQhVJOeC
tKROUUPBzt4P5QImRUsW0SJ1BJm4ksE++0lPCwGvLK6CYx6GnYBawR2vK+HVaUoG4//B6XqBpNX/
s0ban7KjRjSK+Bepc5p7a3e6Zv8JhF8ynFHzfKHdRW5wkrfA/e3gC0ovHxNI1i2m7arc6pmcooF8
8ILEhTU1pyi8tHrBgB1bi3MqEihsmGQuK+lqiIL9v4DozWk3sdD2g5fF4r1nMs1L3E35LohKZzHN
C3x7RS5RdStTOAd9R7kHiOykgEUkKaPNR1zM17Rtjg1l7COV1nTjr7k5foLypbn9BS0pl6mWgQN0
+JWy4yqB5OHM2zv8h8Vx+83KmC7QKX4b4tiG3DS49bPV02mtxWaAfs6AGFaBRw3mVyN6bkJUpAFr
gQRVnjRdAYyvjGf6EycELSZN2s1ugh4It5emwfAQeVI0swbYiuyJiUI3lqEylreVSy+D5rzlHmkq
ezHK2ibmdGKJGlQhX9751n7vu39IAcXAa0xhu8pHc/kRib/CpGmGrt/p6lOicF+aDOYbJ88kAiU3
aqQI5tU9EhV9shbTe7FLUVzR+7Uf+nfZW3bpQdDf3cRIITR/KKXtLCdEbQB5xgtuXnVvlRTxfzC6
pPIkon9+9TmayT6kDQlk4nZDGi+H4gykDKbG7UYqlTs+1sbYD+jXn8OuIqjtWEWlcq8BbDEfViGK
kuxU8ioV+WdoXdhaDicrfSEnWP9SRkdu1fkFyXjT8kAZzLv33zsAbcQOfdnuD1MWnZYKBypr/7S4
irh3lhAyGUgrn3ynOLBl+cEI/v6rlhQBalFnVZRRrje5oTc1DwJMpq2EV1aLCGXGBBiQhRhPTJ9b
M18QkjbjDyBQaZ9OEm7roX0NUmb4i8ktRumzHsUG2PxehtG6+XHtoU+o8abx8/ZReOmhz9eZz30j
eufeglIUQAIvN6Wt+UGLBZKovjW7orz9S9xg1ta574QMMJgLxo1UxBQ7nvV4S8jsu/MYdBDosoGf
KR7MPoVH+klo16+CeBlIJPZ6rqs8vm9dLGBu1fjZy3WA8XTDbIEFmC5AYIv3O8AzE5Sc8RjKDuuQ
gWiWJ1HbTzMnijSSXHmg/iP3JmWqJcv0zXR/HhxOjKcsqbVMw9I4CCS5yYUpUnzjlY8WDruVUhlS
f6GFP+geDNrlGa2DkT+kWo790IieutegwnwpOKhmHHWUtyuRCOQkdjX8sAE9i9Q6ewnH0TzPwiGd
At+jhcJZk27cUoMieyELnUs3NkD3vMjBmJT75VnthiPJi9FiMOrhs5nZgwmjgyLdFFXacSAMNpb1
k2bzgzP46ud6ZocdbG4zDmVJtEyZzK7eqXOleudcnFGk+ZuDeCR0kxuoYTUd/1usrOkCZPVaASjJ
dDERrCAkGz5hnt1ycWhXLpCEFMagocincd+DfbA1HOdPoC0ijWWNWfxhXfV9DlXYIFFRaYv3xofS
U29IdoajUvRfu6zK7bDj4gt9yqBtDetVosUVGV8zdIZxY8Zu0l4aR84CIEJnoNJnz0Ev5WjZCZu5
y4Tzz299kRd8Ab2xTuMOv5bs1JZ1mlTG1UMMxs0oRVKXISqX6kScsLrojp+FYoL1tw35Zdlh9n8d
aXzgIliy04MB53FxarJU5IiAd8qowRnARPDEftDT2aStXtYCoWCzjFfPqYOHOX+6yT+fr95J7EaO
anGYKOmObjU2A50oRZguzefanLaF49Smdr3a6piWbarowXpHK0425URaO9lfzV+bnHeJWUTJRvIV
Vrfn8yYrqyUFjz/K1iExJeR3osdcwD+aACUhiCGZhDgVFINHQmgGVriYuX3JHY8UaLEkDphbe+Y9
Y73iKHG6yUu7KgA8ArmlQU44deZa7RCIYZqmfHkUlj4Q27+YZ6J559KEVN8oQSqYn3r8pDAs+H9r
RAJbefCpEa3lVTwLncB8PyfEsTkqLQTZwjeok3eQo34xpUkD7tdmO0DhD1WAMyaeqdJKFHy/op+P
kLUIVYGMskuMV4wr7LXKctQ+bhdzYCxBflkjfQZHjoYeAzfv2KtdmyLlm5n/3cJ8fSap+g8uW9Gz
TUz+R5nExfis11j+IeG3QCZ92YeJNbJq2J2Dw/3xroRbR9UGwg7mqjzBUkJEK6mKn2dubmr0mkIu
bQPwbw+WFiwPdxGrZGfCkHuzNIdemCi1Z+KYGoEBkAcardRblYNZUbrLvo+PAICEgW7NuSW8Pgj4
JQpqrEmCzsQ7GGx1ssBMSRQnAYZgTFDIOAf4V6L3IoI4QhLx+dbQsNB2LJoOtcebYLPmv9oaouOa
83UdzUinCUT+wxY52ODt8jpRfYoNd3/wFUEJtgYg8BblJnlq7cRBdMXrNiOpHZEjSjlrHVVUYlcH
sKXVX35RAAH1Jwomtaw/0j9Hc/N0QyEb3hDZkw3QUuQCAiEu7yZOTtQRoWmeXKRp1jjIcDaG3qbA
jp7BS1K5HoCj5EIcnnnVNqs59AkbRc0xvB1DJFyXNy2+npC590jI9rzdp+PLas5yDaZ2GZueVgLh
4Uj+p7z5XGLf2ZXsU2+2XIznwIL6sq5nUykGRbJaAwqZeE4yys/vVjvM5srDORL11ejsMoYiEeX4
kiy/CcNgOnqQU9f17Dzh9ZbzQdZB9GWXBWtJLgYxeDlpFketwqpkUgf6pCc4b4DMyBrlB7E5TkOc
gZdETUTtJ7ANrYgYDYMmqD5PfEgcID77IiQrmJv1egYH2Wmk5vcmC33nR6GNBFYoZcNURSj2Eq7q
JZPW68qAfB6GZl6fXzpXADkkSSQVJxNW4Pr7frgfha63+zRpuzxsW1npwURiDTu86faWaBwAYnSZ
+tIUQMq+m2Zi3NsKJ2svwuHtbJCI/9UWOmxp2DbNLuCmJU35n+4VSaE5sOPJe4QQhoQDdpOhhju/
8Srq6D84GybzosXC697OhuUCtmsE3AlCuG3ZaXPygZlkJDnzCJyrBnPflquDzMukZjhiiq0wYZT/
pobBkTquBFex0EkUP1hHaOOx0WtLDgU8FmT9VHbgq6VyCSatGihBFqgAAfeqn7HKhLJ5y/Z1D5Ue
78aAch0gbh71HkSeF7wqciySzCe2fdaSCvUle/bgIjRdDXZ+AczuNTEAFphnH2pz0WyUTxOFAP6o
wov6VeI6rfudWsR0zg/uuJS1KCt/gvawMEhpYrGA1vStLd4FCPYkl003ZMViJY6NXSSMIXc4UyWI
cMl+PAJ5g1nIoQ/HkXugl7WFhW1Mzd9craTHlLbvbe4skm8VaN/9bOwElufUTxIK71aFhdQk69Vd
XoyPM8uulOZ1G3crxIAN/+TZcFs1hbKY98vY7Uf4GnqWGt/wjIWSopH2SY+S6fDIQno573Bpa57s
k1z5Mkm7X0rSFhtS1aGHtvreV9blnKz5tuLsE51co0QsxC1BI++XNoaY2nGdQhw1jewJXd9OA4f/
CY/roXCStzJXLr8OUebV5arxcSSFeLkBuw0IRZeXl0u0AMyDFFrkXz6aieYMMq2947XrsbC1UleA
bhrzWyAxm+LoVeIf/nmLYRl4vZZSowiXIVwjL1WdQyBlK8hYe3dJBQ/9N2KiqJZNgLutGwUoTJVa
oWzx/vZhQBjgyYkIv4Oh+ZEE7PlBmzv6kUPKiuKhwkAd53psIByK8FJSTSLxWQ7G9QcQg3Yhf4Nf
3/66PKVomvFo6CNCURMejhfOsDSNCwOxlX3Fl3IkasR+boD/byV5HFScDdiyJt7szhUaTbq8jK/l
1LF+Q3IWwdLF3seOIeahD2w6R+qX1hvtUxnPfJYRQLiBRBtHiwnqLgLaRPN3h8A4HjzIPqIgSRc3
uVy6ZYAYECiCo/jLuxUUlIlugsQmxayiBRLzUvnZ2vTVn7cL68yn48rd5lwPokg2SfdSqepU0uUH
PaD35bHmwZ5LrQOPwN7AzyDnJ6rtZL8VYr3DYQKe46U2EbFibNgNTKxtVRtEiIIA/D03Vk1Ob6kl
g9B9zwkHamSVi+uIr6H7XQuqOf4iV4g9ycII3jpCPm89Ibti1WKsP3EJQpQ9q0e7JX9KdIRmDLEF
jOn+cj4qIIUYkA73er6ANXKeYoHPVDqWqurEA5roU9dE3/PcXTFI4XeMgtEIaLGEvOVbRZqys0Vl
1VGr1kZittP6lx1AverTVKW3+0a/0Lk7qqd3tL44ftOoOjYldrjK2z384/KUU1LwacZkMOzkm3No
QjD9RVSrBZOUqVcleB4AQ3eDh4uDeakuCCL0MNf7W61CARQ8od6jShKE47od1KogM8Xfd9QqQZ7+
moL/WHYTFlZUD8wOzh7w4+vJV88dysqDZigZF/xXnjz376OkGUwJKPp/wbJSAkvTiP66b+eoyWfN
TZ7L9ujtrWq8a8RSbhvOfDvUta1qNLNc+h6bwXurbZQ9h8FzkzPwLHGRo029P7D9ZpKbszSO3wqv
gsIQYYIN6msklGtzvXOMG3SXIfv/bfOLT8s7YcSfyo6rw+5zK7FnzPnJRoa6plOvaSYEoWeogDFG
7d9uM4MDYsWOo48FOir1qt2tWKgTK8Nd63eqp2kHDU525UkF3mWX2gMberCqPodMWGu3nW0hCNpJ
ZiCpcKLVfNRq0xcBsKE4/yfSwY6FnvFuH7drfXKth3mcv5afEB4odCYIAkq8X7MWvDWT/D3WB2Qq
5dFhTI+kLsDPJubKaZVacqvLJqLetWU3Ft9Y0In7LbyhsBj6jF15rJqmT5TSLPE43+zS1k0dlqiI
ghl3ZsWrfkAQv2TCA4O61Xuzd098pcYuX1Ou1utfZrNYkGxtrSVrksrJRqSZ+0n4BUkMIOVShIoB
NyGBQTLGOuT7yB90rYO29d+ChRXUTR5kjSwWZYhipxEf4GYsX/pBZnOOBHPvdBCeJhm9PfhlxL6x
Yy70RQBsDD43Qpj0zGE/Aejy4oCMVHd4vSFaw0f1fjNEXfzRLjYdO6vl4akpRNRmGbfzoon+1Kc9
w39m86tBwlp85r01/FDVtuT33FgUHKpTN+2Eol3znU5Ew3IC8looZuk12iMHSGmuwurQhVXOlthN
hIPbXfnv/LR7Eiz1TbOzSXkS2ZTvDljYPydb6cU5szc2VjLFkchsgdOVEtwjKU+fJGg9A8WWsTGO
2zkxcc2RcLDJ3HJRNRUDaED/wPpzl21wMTzPfwjt5F5d3SFs1Ru0CVlkZpGTiGKQkV/N6zYfG3Ji
UTlRqOsUbLJzVISC/lB9x1fke3OE0aOEcxRc5awQncJh/pMbJ08/hPVScnARHlZ/SC7PG5hmbCl1
bUYoK3VNiINMpV5XNezYdDhGDg1H6tOU4/I4yEsBq5XyHPlXHnIZ6nb/lSXesgpbFdGyCFWFH31i
2gCo+YMfXejrBK4f8OmCaDdlMYrEo6uA5eJGYNpaFzJ2ZBUc03GZ8TO2pc6HEAjsd7L8/+PG0hL+
gkbNXU6ZGL6nqjv7nZIeWRDHV4WICxzWSQG4upLQUtBLq+nlBC4DYfB3UzMgfvDzGg8HM1ItvGrr
+i0C3/zKxdEqkSLTBU4hLq5+iqs+T/0H/zwbj26Y3OmKMLybBgGlcTgA15cqUgbT1Z3rmwE0CmER
FMTkTowRALVQr+RJ/fFDqNxihBD1+fdK1TI40m7APTgY/gBb++DpPiM1n17lCLR4YfR7BgJMl4Yw
qpt/Gj9clrg5BRa3+L4e8FAZewE3dNZtA8FYDku8GDd+J3ehb+w8BhF2XVChfUW+VminVcnKxaJ1
Z96k9GTK8ie0N/hMiqbfhuvHBEJVuc3OHX+GHgary176X4+2W26fo8HYJg9UnrmWS6oAqF8KDKKI
XHKnMxTG5RVvAVari0NZrj+1BhZqQot+iEhoXSXZOXMI5ZR5p/FhHxd0S1mar14Jj8ELmHvm+ZuL
AIiGKHI+ZHTtBZHm9Vlxo6E1RhZbBphBMRuOANkn7iyRSJ3FQ4u0OfwKwRLltrKL+jZ+nVbGtdT7
qdnE5YyTiP6wVSFCuVApdfSLOd4nw+8DwDFfWYCGD9L05YhtpS6jSS/vESREBLvlgOBTGAgYG6Vw
/f0md8bR3/BsE1ZC6+EJGtgSPSjYUJ8E8QW7QSj8DTVb3VLeu1bt9MiXp4ZZDqYWroWqdxmlZ5Wh
nzrw9p55hTSADzfq397MdKnR1n4pxeDzgjH9Mzo7V9bKmjL+8A7oGo8SBhI+wxLFrt5N7Ey7pLHX
5eV6y1at7q3VORNmPEyRvhft3FoQqBLOni4i9vGN/zv8icszT+SC0MbsVVQT0j4OUJdyCKhSi91I
eZrslJbZBebrp6TxW+2n8zqzF4YtjLVyMYzhybIFaIKqhGPbIFQe+TaHD+tM2G7BSVAa/pTDItC0
KRiL55xjWe73zZ3TdGgF723OSfdP1NkJ1M2s4sWHCD0gg3ObdHrieeMv20uazZ1F+bbnXbpODF/H
e6IZpIJAAHqhgHGBPYN4UBtZxiLVEVYvYh26NcrYq/LfwXRrOna1lu8TFbtHuAR9FNfYTZo4uX6u
rVR76ISpu+in5rLEjzQZIWQMGkMDTlpOkaYGVzaUAf3sHSrekZktrsr0ICOt2gykR1ZH+49E3nix
3dS8OKlDPgWDviIRBic1639nhOMZ5SHIIVkjmHwlr7GIJauqnVCHQkpJqYTsPi6QFDCEGyzqjhXB
peILEjnA78Xs5Iq70Yep0Q5klGGafIZhNmnRFCSs4vGmvI000IV9TPRpjpkPQLy+J4SI4z2M0XSr
v9HLoNlW0a3KiBRnpmMkldJalAMB2xeelx3v5BXGhN8sTKdjl+MN7LXd5PpVcmQw10xdspo0cpkM
ZUkAcs/Kff4xQnYQTKon6BDvDeOrqaNmWFYK/TADhWDx+KxY1vDiWU3PPN3Uz2E0imGDNNaI2p5M
GMKRJB6RtXyanduHymb4xaWrkmsX7tDGPC6t/THGMnud52LJzxQmEErVCz2EbCKZU3Abg0rRPT8d
wh5RCu5KDMjIcF30/gQJvqHh8EYm43ffDwKsghy34RvxzOa1aimQj5S9DY6DAMVp10JPD6KTegT/
ZMlwiW8Z8pBdGtpMYjQ3a59yOGaJdQAxP/zz0HDfT+LzuvQutBTj7djdRq3M970hY4Hgogqg5Kwg
8V7pO/4+bE8nznh8l2TXkvDY4OXQl1MbQUKt4pQ8VfQSdUbvzBHU4aRY+T+TBK9SWjyAspcJS8gS
MDDI437szAVkhGwHhxltH+5zR+KsJXgimTk3lIv9NPhq//uadv/F5/GoWCyC6PsNni7OP2RAhlbk
oEe0C+m5wxP5xDFn8kPSRJz54mR+nIMI+KVb8Rft9eP/1boQ5In4soLVNgLrQ3SAi12RnTqFiMzJ
CX5tHzytLQ6sER4y/B1b3GrFQ6wwFJv84oUbIZSAXS7UglMrtNlYb2duWyEkC10EOVx37r3hg6Zo
gIk8DbBBzx+TTKKUYT7anHLSOQUS+CI0iaFGPyyyTNukAkJ0E9T/qH5G67QMj6+wDwKH9j35YRGA
DSG3Py+FBHtc7/ngWxdmGEC8s303tNktkuON6D+kgKVgLNV/CZ5kJhT4zH8/94YUedjlnq27JLtD
DTXYZI0ysYmB8f1pPyPU5wyQ9KmK4fJt4p7JGja7qtzenyiXaXzeE1PtqME0YtT4n8C8KqUs+xTP
iIV1L7FkpwMCvjjtOQGzU++1r2Vsz4MKPUy6Q3Y6LG2CmNYb5tpomK9tUqU0y9fYOVImOeXXzAyh
An/GzpqvrRNcqaNFE6Tks4AeB8p2LvbUe59sq9qNf0vEhDlNOFWcUC8+ZY0rcRVp6fDi1stETgWp
dn+mPiZMYX0u7OnLX8zKMLyJ6o5GRdryKO9K7AMWXZgF3fXQ9pGFMWjZvOLZG+cPNHhJ6zY9QVlw
RTGfqbpXZ7kceqLX5b7a/gV2r/o16WU9rX9f9crOyd47LtqePar6yWx6t97qyVps813oQsdOEB+y
W69e4isTBNe/mk6Zt5VsIGBGy8VhND6DPoe2HKTI1VW5gm7PILmllHEd7dTBZAQ4wfN3DxLqQyHO
LGkbQum+G7KA0nRizYDHiZJt8aE+8txm514gZwk95nJfI1TaP4mRkKDSJ6Z/fSJoPp0Aq+JNVQXU
cgAeQJUVHHYemRX6oEPZnlKYorQUmSNRFwSesaK0/Aai4TECBlAXYfRkLd62gmuphu7R7Gugs/PS
a8JqjNj4wlxaUEAalngRsdwnqO5unNKUUJjYfOij8uuaRG2GgcNUu94hKga/qFWXsS6/3MzmtAnW
KiaTzn9sHUbQZvKG83y0DwMP5yIkDPU5zR8+5ODRh5jIA7PNgFQ8t7lDTN/YmOCTnlkKgS4pytCA
6UtVjpoLcgUldJQbZ8+1rnE6GMdEOJlrIBN92JRSCjgxef4J5U3UjsLn9rb71fQtsqUf6jWSA6ck
MoUImUD4wP5SpuR2GSkJ5LDvhNPw9ckjqmDsrz7W3I57huPinNi8UTchI9OWcyGNqhpdmXn4n16C
8AwGmcgz//KbPbcESXWQlOfP3SO22+tOm7pbEzw1UhNq5CWaOeujrgZ82Pfi7hH6LmIxTNmyoj5r
q4cdzUdFZla/gmlb397/fWDEEZJ63caY7XDZH31TOduKjkhbUyVUsALIhoNoQmR41SGlUv8/h+EM
Z5QMv/qh1SypKEXdTO2+rXPbSJxKTJqitxnnZWLR64iuTPuyPPi3ykexyiPu44TZcbEmM4M69e5G
YOdr9ZPk8zVeLwkJQJOTN2jwOB5UlmlknhsENecyukf+01ximNUAl+HSKUxvUf0dvuZ8WR9Gv21T
Q4TWq+WBYzPqbP00sPFJrEgKtJQU46IpHZX9GqNGwJew1hVpoPtSCJgx+E5ju2D9CDBp0ZPwocev
U8hzOwqj4e8oqf+U/I8K3ooY08u8Kva2DFGuafbXq49G6cVWFXtlIqV0VCliPJmyc1SZcFfxNpMs
pcQe+A+XORGW6XxIgVQtBX101z4rwZ/7EDPffDeTBLAVsJeqI7hJz5TihzCQlXoSRxy0O4ER3JrH
niT2QwEDo6LvUaGyoZSO44npIfI4JYbUGIL4zW9813fHMbXQsQ0nQLGkFi+FVUmWaHV85QOPiFoX
9rqYMV6qBGMpUVtyX69yBT4tUw9SE1KMFXvQGwvZ6VUDPZNqn4J7wZF/rVu4kBYm7PaHroOupwE6
0S/eoGLnv/NGE8FrymzNtSoheBWQ872DY7ROy8c/0ikW7yfA/mYeOKJMB2EfApPr5r5oCq0aLF3J
CCMOoZp43xRWFuDV+AukIQNG2l+313SakYtkXsuRrRtjOJ/kzQqzeYpOrtwfdNA9b6MVwdQ9Q5gz
Q87j3SUtOaOrkxrpCxdQMoOnoMkuhyKtGxUEmrfP4IqlrXNK6e09SC/GML8utxGxo0ldgP4ujXC5
3BwHdcbpZ/PXCAg9thauWxvwaN4djU3UCh72MEww7Mrrmejpeiu/W1rH7Ebnrm5HRIvVNcBFqzwL
vedsqIZj5qM0/rHP++Dg8zrqYp83HQtSzFmWsTGdG3b/IjERAtRC7MzcQyoFxZlWucwV+ZugCJ3+
FiTWcpmgL3wqmL6nYfRrSXlXqgjuCtAJ7YO6rcgL6sNqB403188KPUjS6CIrQEYXjI8BD3FBKoXg
GelnkyJmR2sCPP9rc25zvDicbC13TiTVDohoJryO3JTxsODIzqe0cHD48O3Z/G233G07YtAsMdMW
8Dgd3y7STAm/TiK3maGBzV9AeS/46ytJLRPk5CuiFBpADrMQbwC9bvGIG8VdTNK+bxKRPELqtima
uyQfTHcuzuweW8RXS4U204yhPWB4A0zGCUWHM9d+6EfeE468zh6g/iHdyoQpe9G4hBgW1MpAQFUs
wIwG2t2oETd6CLlI0o1r5H8NkvQZIfuTQJxMpTFrmfZGGrvCRgv+YM9svHB2mqtH+2pisAMC0W6O
DSTc4zlBagoKHimISn9GC+p8MXObP3oCDp8pgEE2HmAU+M7JKG8rP+I2n8oMRkVIK4HBlyMOHf3A
4+jcOymD/a3j0Mu0LubsTl9g8gesovh57gwc+UCoSLS1nJdfXANSzm1bHPzp2KjGMrYvTk973ywi
NCNJzidGUUZ/aJo+OkdirOlrPQQ4a21uapAo2iMxPAKo7XZeIMpsKWklsJEEMzAJ5hzJM+pIVybT
gRxOuuV9xsaOxA8ypsg2GAKwPvIc+9c8EbAc8HOsizkJ7jssipNiPOWpBkKy5hbI0RDooG+WfHuL
l4zHEWvgThKMsg87h9hRky0mxjS6SnIQakPVgBQ7gKkHfmwcCRNjSvN6Z4mAYzmKvV17FITgAteM
+VuBFVgIEyb4v1CHbpoIj3U8J+0oziK195XJqOj5qUvMffroWkTlceIuRIo5pgrow8uKBz+Up6Eu
zFTqHDyn5Firwb2X6fFW8DklSNCiEMHaeCsMD57or95paYIlLG2scbhDH3LU/e7046+cvlTZgJNG
+a3FO/a+r4e+VyYhnJvL6yoQrH60xww8a/7VGF1XMOxEMGeMURxLcTEe7KloM3GuOQ/CFM/bzoFV
KAcnH91mvRRLZCJ5gyzL/yq8yA21BYbUGhPj8XI2NlrQpmZzn4194ZMb2sFZq3VRcBqs8u+JFBvS
dGiBsIu/V/e4gPF52/WiOTe7T/IAdykeupmp8SnZgzy+bV+cqE4uj6DhxDvEfAPmJ1prAegkDHji
SAhKG489ie9SqoLwv/KV6ZKrG6CIBEUfG5gpotwSIRpUGt2haL2ypVNHKghqCCQm2Pd+H/HMeZG4
7kNSWlO5pot4qLCMW98/5MrElQPioF7YxFo3Oi4HtiNWwebBGQw8oe1XhE/RjeQ5tUhVGNg2xHfr
PDUjFfXqY7UXMy4gksqQJIdXq5cOR7yo7Vw+cOYDgCedKj+Ku+5PSj7hNXWFemq18zvOEg2c9DxO
2+Uf4FABR8frHpavFgAjOdzQyrONaodqCQvIwHIeyEalSK/xLKs6huFNdE3SVl064TET7ApF2hR4
alkTwO4Ylr9O3Uthe3dTI3NbClWMxB4kC8StLumq0D27v5Jtnp2kHNmNqjzc3TWpnBQmKARDPnu0
wIsXabW6k5bqyYL0UZ8ouJkR07a3Bi47zo7N1b832cqflnH5T2HbCn6fNOV9ICxZWSwWETROFPQV
K1CpAQ8d3Fsha8VbL1MAH3lX1UDmkAfQqIyYMvZXGcyEqjECNrJGPNreINLIx9r3BNna6UC5TTwQ
JkTLuEaPv3djOZR7UB8agTeCrrFTychFvXZh1l+v5zG9mY2ZZHswfkEM45/hj8DF6c17p2PGKVUh
WBROhaPb25pCkJewH2yS5bkWcmrOHnKw9kTs/4oq4VaqkTKmYo/hNlvSeEVqX9r+lTvnaPtZxILI
s9z+AabIOS2QtNw05H36xuS2ZFmLED0FuUx7yD5qggmh7qL+5JB2wwjVetAxqXH1l9OBwi84+8iy
nfoiogZyuADYIMIIvE1KEty4xBPuuVrLA0qWUFeyM/kqUkPqtkQsUQvQF16nIAxNOMoBmwoBC+Ku
ikTkDyNG3RyGXa5Ki1HrDDaFT2cTZi5en1CU7CeT0pi3ENyd4hh01CpWZXyLSurV/Ip05XhJxiCw
Gj2x0HgdLRLgo5nR9LaWZyX7fHTAD7T8PN4uiJR7GYxiQXx/sKlfFj3SkjeVKO7BSTXZkhOQKxSB
EpqP9nkmtoh3lLgCL4cP4MVG+J9jPb5KMSP62tRXR7Tt1m4Uj8Wle5o/Pe3WfHz0GNljVCdNHfjA
YvzC/rxB5u4S021wMQ62csRs2OiHnCG8ocQEJnBlWUgLfOVt1IOiD/BAdcheSS7e0L+Cjc4KRUSz
bh/BvnR2qg7PkEuUM+qcWQ/ztZx1ARdsz25duC0rOWDjvgryxbcAzLlZb2KEd8PjLHsR4LdpIeOD
3pRksujWT1t5uM3/KU48lez5AV1anuHZlvxzfu5NtmVXTGWlxjxo+i1rx9T8zMiLwMxKwIpIuoeY
tMpsfQ+vp6JDsILQ8uMfTi10OXXhiZPwiudQkBtGSl4hfo1x4qQovjBDHEhXAIcHHqppQkCGoxWz
w5wc5SIDfHERgWI7/FccA/U+GfeWJ1xcL6wWmtyEQNBoOcIQ02aKs9NHSlHOG2oPecJ14QwzmywK
93zNIM0vdppymSpNu0wDNyuVbeeZiOW5YNHgY8ozSzWjQOkKewGyHM3xjqP8cDJ/gZbDJJKmTaEB
j4o7M2POpuu+On2m9cMKqqh3krB2zOkXfHOJstT7RzNoKMYMDCdY2ExzaKmy5nvt56JJyclUzX9l
5QBk1ru/kK9RsHNPT2qtq4qk1Gg4Rm8Cq7C8ATRV7j0B/ntTo2FvC4Zlhot2WJ7YSH0KAxs1iK2I
M5v4fEEUWK4LfCs418jBSxz4UA9C5wfWCUWnV4Tfnt2TBqcsP6GTH6NDt2EfW2ERhpzOMnloI1DR
fkhPPuuACNtAi6ReGYGUd+UJew6HVkCnYkLxdHH82J1Cb64qfUUkFntgo4sWuIM/TEiG/mY5xcl0
dezx1feMp30aew+uK0mSaBNeAbEGqRxMePN6UgzGaOf7fTGIcZeCS+2+EiuNjVHFuuXkbn6pYnh/
4u+PpbQ68hrcuYSKcX3an6adlrwS/lZkKttIg8r8n1NEYIXaAd9c+ym+W+ViNXBeWJpt0GxCfKCp
FvwQGEZRojGqyDCRDzsrs9xHpYWBbbXNqLbcnjKOdwKogmSM3GULMnIh8SG5g7eRtosoAwk28mAH
Z21VAgXkS/WemYaKIdivnNpksHupnzQnwRUXrEdSK4R6B89viN0fpr+xq8+AsxmVdEDD7k59Pu7t
AT3V0OpR2ZRMhoZO67iIaGyRhC38GC+GPzC4fYWP4VJ9O8oWx4DQCGv45fSngc0cbeBZqIjqzjp7
3D0w6xsUQeLxx6MHA2Wb5nxiNh59L8tkUYJFV6HCVLwxWHzRMEeVUOZ157SKEZ4kmjc0txeGzoEE
vpSKqjoydhrunAgFrgUTbeNkc9JXZc3rGrKFKWVEwfX2fZ3gaHkjI5FszZrEdjOY3Qrivr+ZdzwH
FRCixd5oIbwDqmDFFXe8i1kl93pIL6QOSNnd9UOOba1hoRw2rph0ZKQhk8vZLAXPYbMe6ZFk5yKc
ZW0ffNvkpH/3WeDKTSidlBtjo3BZ1wQLqZ3r0kfxW0J6PNaUqsIy13qf/3TOZVObXQPu3oRnLVL0
GWpq+/HOjrUYwAjqbQGqoRTrxfFHLN9BkZ8ohrv4i3PU1qfhlAIC8AwF+ePpF60dIM9bWs17CNhZ
AImI2xnXzhX+I37bmwF4KdQFypTtzXy6o7pH9aXW23J9vIq6xNjS1+2oC5ubSIlzTWPxiuyFM/5P
W/viPsSD5j6yfNhUM0YHGdJCZY3QT5JEv4BpgSnAShFBU+CJ2OtubCkPzaZ+3Yd83H9J+os7uFhW
X2AVsSMViZAsFxxwAmngWJin02vylvP5dfBdw6WCp3jCTjzyvx2o4bctCFa5JQIgszXmk1imzo++
ZFTvGOPNMMnzAM/8xXEfD/GZBFpv40dSHssRTLt3aeHX2BxH/LkbIYAuxq57dylMqUAL2zNdngBd
pxjCS97o5AXH+VVOGr4H9gxpaS1aSQrFCH0VLaP6VjKd7uFkcqq+7P9TD8nYFiVybnJan+bnq2HK
dF0bJ2zmee4r6AmM7cqhIwG1TV5mtw5Dte6MRHSGhH4ZrcgueClFx39OaqP1921iimu/nUBudlM4
coqYZ60ICvsLSH4dmCKskYSgGF03r4bSRyrdGgfPL9DspDXAzLEZN2lAFWnUDcqgSsbNZiih9DjD
PLGgCOsqvYMY9Cr7q19C/cn/Te3qfrXBzya1Zs5sd+gtlCLlD+EPeU8CwaILi3a0dBzM9zm6nHoy
3GUX2o4MCYCIppw1xYwuZTpvt3TnN9niKtOAmLBYAesZpqZkBN0mEmKxuPrMm2HJGKJ4R6BZp9t7
eM9/7WLkAD5R65kxEgfE//zxOiG5o+1cd58NF63Nf8vpu5LOCh3dltzGJIjXajWxxYTSjKplIniX
o45y/IMfnjDYiok6CrNkvbzZDxZ1l/VHd8KOOq1uTa14tiRHCDEqBdEgST9E5dBgu4sx9N0FWIxZ
ZTrR2VU1oz7VoCR7RfHxVGr0Dv55yfwmDqf5FyMCESSl4DPSMPbqV79jXT90amlYZKzh6LWBoWjX
vX8qODk81GW9ZfLSYAlN1dh3VFN4pR82ozQ4BGx+XSlhc3XSaUEH+qtVNx9jfb2G43I9vUi7FVEp
l3Z/UjPraCqQfhIjsoCM8R4UQTU8msK/wB6dbFrJy3iyikt7U9i38uXTrwO7TmB0KYSv6tr8YyXE
E8lBRVhYW5sfuDxr3PsKOVY4+Zbn/YtRK+D9fGMs4y9zL1zM4dl9N9N1y+JXy6TW9XpdAd0zhlz9
LxWWptFOQ5sc/AmZtdyHFE0Y+6ZucmdmhB2k98NjQLiUtyJemro392lDlvuNFcmIb09msN+JvYnm
l2zs9uK/2u569AFP+G1bW/m3yRSNcf4l3rXmVE3o1aEB588lELDBvgjmPF1enmV52KfVwHWEusD8
EMHk34sFx8euPsys6m87n5moM8nJ4oZ/wqy67vMYVZmUF1dMIuITwdWf9ATUUkyynOFAadhqttuZ
nNlFyTfSEnukUCWusBOBb8s3qeK8qtv3R7j1a1dTytzAfgr3BmRLL2moY252Bk4Us9bDET0uHEW6
9+OqBgoFYuOMuG+aVqBsJHC963U1/gWBLpLbxPdc6/7iEaNdXLYEwA5gKnFJtb0jVPzr9V84cnOK
aff4rFUbaQEGDPiskiaddiVWbF33dUDa1wGJJ9VDLz07PbKa74atbG5oYWSGWEmXlpRTzQBhvyoM
k9vF/UOemTanZxQQY8k1Ro78Q7/1J4l7NTjeBTJlO+/9UPlVv2ygOudZ4FCe4d7qvQG7EAj2DJQ1
ZM00N86RNFgUXHPbhkmOpLpSnvL3UAU5gujH/87rwPcwEv86tMix55bxUDGB7adBFGfcFdFmNad3
kw0zgsaPSmULsp8ifl26NbxotMEengO3IU3iBQv587srXg0PlKKRYSNcVgjNyRLhPplY/6afb3zz
uo/83v3vE0WhU6Mu6WxjxMghd17O8m+NYOAX0Fstm0ZXoLrhYlsCPc8T/pM/kej8S4iycJ0jbGkv
tKVoFkqci+dtWtETy8OKNmK9XJBSv1V4GYZ70f87p9n0rEO565kTPKTOxonLhQ+OBGxPglpDH8Eo
hsK0muKhmzLcNCtIh4BdToaj0IoK5JmWy12MIB6vDUM5kpMgeGkolwJfAHF9Jp2oW7GurklFnIif
H1AJ+7cdF2vKgJlZemUx0AxDZaTkfk/w6jvMLiyx62ooTtnBJIHu47UdCada3qkslCdBg/LWRye5
fRrKJVa8USRCv6LpHKTmKlACcn+dfxpghge7dPRCKbaXZBJM1t+ZpxTWB7C2wvz/wQ3SNfxBNJMz
04Sceuej/QD+G+Ai8MLz23dYml0yOFZC1nRR0093AO8mcZHI4wakGDbj+cGFtUeryYyJXchvXNPH
C4pbewxse+VU25Spzg4KlqKqBZ4J5tWbBJccmRXSjhW+izh1Zb9OwbXFs2j/PeYAI5R6n3PDCJmW
qnl/0FuglfbRzD4nlOex7npJlkE1QNyiMKw4dU/+hjyi62SwiwFcIHdpVnTQ7DztoUQs5qv7QMkH
vWS3Z5kmE915BwRKVApRAJSsE5LKdeAIyHYUpgD0ArZf4IWT6EN4VU86o7voHJllXi6hVpLe/HJF
fVVjaFQV+i/pufIBeSmq+FWWY17schWT1ddMxiZPNCyiDcrLf1thHNDfBDPbBHV1YgUap32SDb6x
vJT3xMFVHZMyrzcIWMh4xS+alIJOTmS5J40EJzduIDVh0JDJZi16isswqw+9Ea2cK0ArtPRm6Rvm
Qo9IGeckyDV2GqAWPDrldUKNV63/Pzr16OYc517P/qCXQjHH4LgPrH6tbFIywG2D6BwirW7RxffR
HyREw26IplTwOE18rulw13CcFQwdeVFsbgOxj/05DAPnhLQBlW6Tmif65NdBgGt2iDHJEEmA4U8H
UhkuerRUnv55RGZdCO+AmaA32xkAsjt9Ztd/3+hdW2XEVMDKtBYeTPkD4H7hGarfMCOuLBmn3UrQ
CGnzZU8la6yVI2QlPB9av5YwaYDQzglYn9DTd4Fh6s17LdeIunQeuoWmGmmXzO13HVX+8svgQEU0
/JeNqE4vyq/BFgB2DiYYOmzY7Q0heU+EEluDVB1VWSF5hYEOEZxRcvBbUQG1cVdiGEq2waxfO3UL
Hwkb65BYFCGHUIEjJ75wuMufzIDD7bNpT0c6dlpnZUkhDy7Vi04ZZeVpZsQY2CUxfZKLzUhoLydx
ZWxtIJpes8jJRlTwBztlTEcMRZ9lkdHjYy9Xv2iBijX4F7JuidZuCO5Cy4T2pDp1OKl3qZoEdpYq
zRF6Z8zZZPF6sW4lKLCH95QNBxHT6U07k9N0fWwZNnRUZCYmSByHMFaINC68LYQPsArAc1fjEBk3
WJEY2YnSW+RcZfQrRaRvxI2oU8EDctRz8h78HqFQSwUZnY21kTA92nEIlkDPssI1NWz3RMPg4lqR
/9ZnacseZRUFbFZ+moOpLELhmhFCo9mpfliood/ZuOtXD/FTcLwykKTRbeOvLKsQNFXew1PRgnBu
EuUvT9x1FeL6kYAlFU8ri20IVJDMeTB7ab5Y+ThHGeoFGmbNynX3k4oO8GDsP/ZTwJnYuwAMG25n
oHPHWyPNHbwUD4pMPNUMEssYSOaPT+RZ7HQcGcrb1J5/XibmXlkMJeA5k6AgaXlp/qUimNEJj4Gv
CdAi5OtsjQ72VT7tXmYw+o7Hnxue1Cj835su2uz4K0SfE+VQAjN1PujYlNbkob4oG+RqwIT5x/1u
5+aVjlmeuhTLy8F2ELShMqARafwMeKTqk0ph4WF7xmFES+f4j+g8aWDVTNNZV5haNgKlxlyJkdCR
+T02drM2Ybm5a1HkmNSQS1TY5/pQz+EQuriK5HZcHLFDTHVp02Bfjhi5YBw8jO8VG+Lk2jdBFDE2
5mth4Xfe1cnE5wnrSynfWkUfOYRjaqjAco+8pSOcGqZl5jtsOWV4KA9DgIUX7RCzeNGqjomyP7yt
DI/bHyUgzKzvohkK3ZcDKaVTOEl+a6NaArfbHerSgTbZFHPk3nVYgAhER9QLL38vOacBPWz+01L0
9pDdGZWSvUy9YeIjoQiMTZoV9x1TzHkEo9O1nH8ITY1lmSRTvePgcGcKQ/QO5qVWUR2KCL++vfJw
xcTaDkflzqr3TzDZ3t3pdOEktwnC8oToggAYLDlPrty8rAWOfsSrebdt4ZCTNc1cYH0nU3WqCPwd
TUqJDBNj81m8sW4GSClTf2zM9GhwoxuyeEUsbzFqB2XbHDeEN1PmQaqVhX1N4xvAntA5xalzed+m
6A9qPZF+7iBPoD9jatXkVUs3b/Tjn5gJfuqzV1HU+1p+zJ8dFJIF/SjDgbeRUmdIDD/PzEjci/l8
5gF41saGsk8ncj89UeCFMuetbj3bQg2IdgEySGdaGirL0tGtVI+ireLr1VcjMKz0TvKz+vOvr6W5
5uxn10B7h8nu7A7x5ltHLjoh4IQsO3rS4S0j7JH8d7iE/ZT4WxoHDH8RSciE1MAeYUj1VsDNQqJw
69KEfiZkZGE5dZHd9+fv5Jdost67FitsU7aC91i/KUFBGj3uNnr5oz8tJhIajpZ+8Efm+EUnwXb+
7AH2rl0rtvRS23AH+XMRoYP2gvaUeDjgVmXiyiUcnke3BVFqA+M1C/OGaEIktgsuZHesE3QZcaTg
9lAeP3bIFmm9GF5KXCXI+wMCF+irJI7Q8Cdlmw0oj4w9YbY2aNHAO5ez4Yzix14TkIv9SE/AzuCw
YR/r4CEq00vB+zh7OLFayiDYGh/1j1OjVho/uddCjHpaw/BCY9+ML6DgDIPFWeRUF6J6G+Et4asQ
3pqklvB6zCl1lqRdxeMVdxL3Vst1dk8t4iwkk+bpP9knayTNum5EFdY3jnIwBtBPDB9ILf6sM6A8
bP9C0c9eD7gi+GSZCaM8DEQ1Phx4DYihO+cKpFgtfP3Q317Akr7z+mOqDu0pmIH8AhhXCO1Jotlt
Of7Eil83tzSxItQOgMSOmfVFod7i/PolTrA4a1kNiemEUKfjhoVSF9nsr5Yb9elK0qIhHqxiVvn0
ZpyMnaL8d9w7Pu5Hv1EdISjrP+yZ3bQVOPIUd1SqGE37ArMGAcEBoUgxS1c+CUdT6Z6rZS6Vtqll
zncdUsEn8QWV2JgjmuBjxiELyAr5yZsgB4xd1nA57OVjFKlQnY7HsXGEYipPC0/8OSk9/Gq9+lAr
GtEd/m4lUXe2U3vo0t853NShQuv+fnwSSe2QbWQ/AhzJ2XmzSKutkeCtB1dPtZu4jl38hKZHjUyB
M+1EACmTn5HJ3tc6btfqOjk/1fTvKEdVyrhD6YHSA1Hs1/a2QSRfsJVzwtzD3Bw/EbPDMvcOxwec
1BjPfhjV/zf0sDEOqrj2YmbUzlz/ibqY3yvCLLRVtWiUUYAQLBBV5HwIAA2TJol+SqQ9pu7+Ix6/
ZH29hluNHo5ZbwsRfhfzVo8nrvjJgKW/KhcKOfbRdN+Q8MLW6NBKSoDRR/YGC4KgKvqmUJ6NVMyc
U7bitrWhjO/CRwhmAqHO6YS972s03L9cw65OmfrZi00Fij40456r9D3sI8wM4sFerLXmAgcV9OA5
fHrXCGNLOerA4VkmtkV2w0NAgH6Pea7XPiMnXNizhd8xGMmBB7a5/g/YKvKnKbVByBXhwPf6/Zzz
9vBujoEOntaYrPRT+2iINQemz54oUXQcFNsFPFEsk/cpqaQRqIwg1UYA7aY+RSDOHd6sX70swsz0
amNkZgmxdcckVY9wWQgH218WmYjypPM2o7acuFmsZ9Bo2zWp/8AsCpMfBqsQeVXEmAHe28nUmwjC
iTKrFvStYBL+Y6B0mnILDn3caG4S8Tj4Lay+AH4MDU+ooOfPbkgXRBAZL+/2dcE0lMnh1BBQ2caj
eHqQR0S2wNyqoFt52EXfHdSq6zQO8U0vF3iflnoYa0R4IqjJvPSrSAUIV2ah2DBKNIYsYh4s8edg
DCj7pl4EcCjkXYNdh5pTB0rmh0kIYV43zd+rSgzE+yzUrxCuJpr6oiT1Y2Lt3Zvjkwr9cM9wclMM
27G92omkexVAdpCGFkNnql0+uLBYAK9B9tx2e3OnwZu2mhQYNqWMuK1QQA+BNBgHO1ahBDubDYz4
2yNw1gOhH1wz/JBPTC7CCmXP720kw7p8ANlDhdx07QpHYftRL8dQKwf4e8ZGTJNsHx+YZEPm3gTK
mPe2iLNLuktfc1vlhgZfrl14JJREnxfwW27WBhaHFyePlcRkDYfJsRXXZAGIyUvBrCsv2DT9GHgp
L7W5qX7Fu7DlCbycaATU6rQFTcGemabu/SU57E6QKIaANb6qiEvTwP+Pqn8UgwsQqDOUJt+MWiAX
EPyA63AxlV5vTtQ6IufASJ26elMT7SetISfYH2XigXkK5SiePrN8bgBn9aSFmK4VP3CVWJ8gRV1a
OMIG375a1ip1IvuROldGZ9ID6aYkpMCjTPlil0TayyiG+11m+q6TSuuJ8q11VDpvqCR/I2AWZ/wH
ZC3+sXi1zjCl2WQBeYPpnbQxx0JXlBh/DM9Y342Wq2AeQfdiSt2UCNlUBar8okeHByMmIETsOF76
bye9siw74oEE1p5ih2D4O2mZ6wQxyLZskW926PlEy7lGhN0BRQm9WBmyIDacUxQkCKokSk0rxesp
2y4aQXGmvguXSbxI5mKOmgDkYo7SF5FcqlZAu86yDdlVuiiN2SRZJ3dQFiiScPtL4MBXvs6J5qu5
nmEHDUOWIgqEqVTVSYg5RViXiX6VLmMol0QZoUvQ8KnK2mFG9hvUg9DeTusZyt4CEiXqxzK6fyyw
MSUJQbnySYd78BhqETu+LR41ocyxo0o6/auKT7ZykEvpND2knIagrnC1QnCS2+JGgGRoolu5YVux
fGa80feI65l1IfCJevbNHC9geCU+Pwq/vB78yS3FWwXMZpQ0j5ZDqy2K7gGXTYiFCFZJKijI0jbk
vErucLs5h8ZsTF2gy2VtbjGDX32EC7YXVPn7MlWTq2FYpAZzwkrlzt6eM8/b05/WKKWL0SvR6tGb
cLWoTYRb9Ywa57N4zRh2WrYuqpxBQdIDaBsx/EphLHKP1K1iIJm1xDuFhnE146STw5qobkJf1Xwd
5JXoZAgzl+iUJor3Nxeu4TPeN6oWnIuvrzvyYes+1v4mWSG7S8e/vgVUWDYUQzTLUjahz0JN10tT
uEsA/VDLyjerHLsphEUISaBs6tU0InSKEg5rj0UPCdavBPZymE0+VcB3veiS2+jIEAmi9cUEupXD
bDgjEaP0jkSaufiqn91be6yU0vCVgqCP19pGXFZuWWNGpVn5pjId0XhkRwHTOYeqLTIwXrkwgGmF
0NqmkuS2jqcAOldnsJIYC4B/UiEOl4YEqU/XXSQadDHh41S7qMzU4uOw60/Vo2xwuDNXQH5U6l62
1+H5+VxUS5RdXWpjMGJ8l5++wtNu0x/bpfUZbGBn4ar/8DLXBidSql3UdE//9LyoYmtDVTlxsgtr
UEkdJqRCeVFRipyqGdC80mYGpmsCEfGULvExsKNsgx/gjVqMHBPyRq5XRnDno9yIBJUJ0d4F+hqu
PkeUifECo0onvhTKhalKEvzPwWgVJ1sh/8arm1K6LG8XatJySTnVRZVcRbgVmQKTNX9/wi2DF2tE
hudt8ouK3CyPx8OA93QEnwfRbgy6yN5BEo1+4rKS6r9JfWkv8bHU5exHGEiYqNo7lfnFSrT/cGsH
1UjJ0fiwex1ZFj+TCZkgWw5VnpRKHd8F1HfYKMRxdFW7X0CRSfb3obcG3BhrJ1l/czE6l4hCG/Yk
nl0j4S++BB1GBjN4vZbG7O665rIQa/QLavYOEuZC3Oay00P8t+3JdnMiu90cXyPz+3YfEHeYXepH
gJu8Y1uqJLMsB5Up9XIvmdLL81vAdSb2PFdzddl9MRetqYQt/H4T8XY2SULMwBHLM89Yjk+VomCn
+2fykbZFDMvNaUMbhkEtV0yZ3ZozvA9Urg+TlphFFF/4zb4LBY+GjzG1CTkZJchnrexMT8INXVr/
LAZKWcttQ6YcAJdXw2fLj+cg1558l96tRMBlQgUMsPkEAwe/dLFI0iG+YL1Mb8MziFET2ANje+6/
k8A33j/EbgtY/ce8rZiu/r0/EcQwnMqHT459kzq++B40tySjG7WMfRu+eVc3V1/bOL6d+YbZzM7G
zKEpcxJV13q1yqbsr4Xm8Ft45RC1+6v8ZVnKmQapAc3mYjXeW9bIn2CcWXBdmJQxiIsCM9G9PrJx
VClc49QdriXgDjE/3qmpp9sm3q6rUFMUn0lJGyVgzBqYLT4nMhxfYpZTtU62TaChRfYZqHFEFyBc
FnXFpE5sd60lJAoHRvlAFNEjgbyIJ6X9I/jHyrP4Qfrl2vW5IBel5YzptycElTKzwKfC2l97rzDy
ifoXdA9dxa/Ory1iE+cF8XFYkbyNdCLMxSXUV/Z8gqIktk1qCjDCxZuasnB9+H33rQLVSNBhUT7g
CSUqHjqO0uildnCpN+bRn2RBgSjf9ME/OONV7JNejXrC2XalrIDluMm1OAP5AyA4dH7iUqCsU+AU
RbG/0k8ej1s7kwF7w9x82RI/nokMtgbddrP68XhiHBT++MKkGnbe/piOEgjq0t9hG8g5bkNMcUPj
ml8bxo6MpvRyHwPPvN5P4fzE/fHKciVBMJhGvog+jux8W5YD+jpanoQfIzjlDUzlsc7lPmuvz645
gEbrZfXCALCJOjYpiXAdoisDj5QlyvZOwyk138Xt74gDAOQUXOQv6HJEt9lCMp1RVlZZH7ky90i3
Ve7zQ0uJDRiRIzC+FP/MSe0h+ICumfWvryZN2AWut+UPkp400xOXZ5/0+1kmvyqOGzOPBNj6xsYY
vIBxhNiB24dxLbfI+b6tIRuQsxCI8j/lsZxwu4fI+qBvyX2R+HrxjfuzlDsurwaUC45AzqBD+4yh
5OQr5LL0TDp0SM6TyTLuoOJk1DOBjDcRkI2LpJ7cY1+RqchONzfRL5MAzVGxU6CEtq5uNRurgv0a
YZSQIpBdcRnC15nTMvD9QUyfAHTtgIryT2ldmq23fjyhcVzAq5MxuO0vngWGVF9DVjKN8OSc9HQl
28JU7pAsWACdyztr/Nr+LvpYOVaIRxSB6Q22gFbxyocr65tapmwJTl8W4Azd5HiI2umyvScRZiFq
4vU0VWnYM9+N9RdQgIKf4NSHEP9GEyhOhaJ74bNFwACwTk6aYiiegw5KGRb+vL/8P3h5Jp5gPzSJ
wrYH5DBUGm0Ia5R2qVygNa0dO/ibg5OIRzUMf3sGQO1rkOYTEvZex5b5A94wh9DHL1nZVdIYpOji
lh2rj0QUWrHsexbfjK5ALjdZ+aCWz1XOLdjMpVkvce8zJUkhZtAkbyRy55SQarZVn8BwnG4Kf/i7
YAarOhy0fpwgkhg8nBMoNCVosmFWjoBF3xYkj7i6KMXpmSzzjUeVRNBEqTpdGbKM/gXmHgGHPSiO
hbCU7VnARp+iK8x/N3hWt6e6wuMh76feS9YZoBiaSdrUTA5Bdd2Dv4+rKYeveQ6MEh7qc5phe4ty
CRVatxzkBiSLZa9rLKH6qL0U5FeomV9reKjUGoBTZVW0HbwrVVj5Hb+g4x/WQ62p3I9FYihUfTmZ
DgUE2ZwnffEdZi3h3EF/0KPqmQknHNiZ2Fz3X/elAREGA6X6hrUqnU8t30uLSbBvszK7VZF1/3Qc
A3lzitmbq/KeFVcwo2ntgM2zXL6e8mQGhXEOloWeQIsVHP5CfzySQ818IGHb0BNW5p7/AFExjbm+
II+x5mgOmNNimssiWU/hBNmw3+Fr8WCgufX89h7PG3w4nBjHt9XqyVaiyWlA9+YlkSf1POyG+v1r
WC2VowwifYnoCcSZRaP09oHScNG+RlROllOsk6rjQWxwU5Nd0zasxAXqpOY3qkzmFR0lVyUNrLzp
unPAVNGzVrrw+qpjz9rf4yHv/4PTD+VdO1bkRH5oQLPRxmO1UpzGEx2u5KwgNLxFKAslaHKR0OG2
9pqxYZSyXfyQ6l82ShCL3zdydweBqcSJCCBShR2dg5COAkckWSLVT89CwjIDt0WaKWs7NGGqDMGm
bEA5U1sgS0Epq6w1jtJo4RdzWII8dmlUiHju3UI9aVCnoSR5+y47i5EILenXkyV4/UATDTLtx+Dw
FfTIkzBnZur5f6VWOFzr/6yXoKs+M5EI6QHp38pXIIRsSXSpaccRBjSTnPzFEhy6y6JlocckQGLM
VL13Lp2pSKOazoEFgDHgsRpYI/zKZmY9csTWOiqYiAhqzRiBfe6TiCUlW5/fG/LRc+WEjEFvaeMQ
NfVnTeDXfIULZ49xL9eSw04YMGY9coFKAGlX86zckwXEvzsswXP+fPf9tcZBIAfWBqJGWxD4IM43
ePXm7tlP3xvSttyEo/Zf/tPQ1YMQa2wsK/pZRUtOArWAu7hwuYZrF6IdMhR5PucGLni2xEIxf29N
d35cv3dej/d7SoZZdni8/G5PK5hUa4ozgcC2SOUmErtOJ4ZEEbNA7nOouhFF3JxwEfFiItzbCaIC
m2jAOu2UdT6N7SKOOlV93U1cLPzxRWVaxkBGhWfWRfBreP2lmeAhS9JZlBPQdDJJwOjHkemnwxUv
+g+X3U8cLrYHUJ/xS0NGDL3giA38EM0blAekndtYCjHGw2Qp59xCK1dJntbBYqO45dV4qzpBHYri
O6zqunliv9cLpw2NGBJpxdZXD5OuNFq/P82uryW9Ktn1W/4RK1SaA3eD0oFdvcHhGdB72MVb3syT
I9awWaj1VkGnnOy8quWOeGrb6nvqwOJDL7GvzrM3kPWtkhS1eROSYVkWt3iP6WHPD3P15uhk3DEB
ZNl4aZM54C339OaLYFWK7oCVGQD2ud9h8+9s91IyV7askY+89mnfvUrRUiyuEsVRbDUILdUTTz98
MwuPUaPCMTN5Ddl0/kGZWleO/ihnWxjsi6FguEgTRIoy2rZAWswCielxJmGUnlf2rE40L/3rnqFJ
2VGwuaWZq+MzGaTjMKj5Ulf6TtJv5AsmE81VnwQV3XZAFWdzPUs7qTLREpBFfrTgcnIU55KDTifp
Eudb7ARfFpELkaB9Ua2pD72ZOVnBk6Y61VbgQuAwPx29dIFfGx7i1/gV2AFeNygbTGnh0YXjY6a1
T40d5ZMh7+6GcEqSdpKAY3M9JWERjX0v8s95QMcKbYLOGjfUrZxAghSMW+T48mIH4NNSYGSGvFbj
EYs9lwjLzcpsHbm4RViFSPyAEPkUgxp8QayWN0L+LcVXDqQ4dez1ULG9uvcpd+gykeV4J8FHuTSC
5LvfJv8EeWFN09Km6Lz0qArUIbWqKptAiXyvZUGGVWI3E3MlDQTVdwmWak9q+1PbLfxHdYkb68EM
FRYYmzbbxu4Y9spw/03MvhrY9aBdPWsGDSCMWA4Z+QeIj4q8zJx6ma+S60rSIJH92muu2pdZSURq
eFfmMSlFbVVbNx6oHpOSkkm/FtZrd0ex85d6X/zjbxOTmZUIX9ohoAAl9fq6Wy5Vhp4gFNHNhmEO
8wDeRmpVsLhzSvL3POsB91cHfMpFdWatiyKFha12ePhmdDhgj8Mq9eDHyCLSduXjp85dJcb+Xthd
13sl57QYnw0yTwpjsKSR5t4NKEFsH0MX/JT07PuitzKEq5o4GFLdbgw3dQEX8wdpNW2JnRAxPA0T
GxuFPQPg+jQawI6yxubdIN4j5DNh+gORlmd0AKTwbpt6cIy1g26bO6OvBkOceO8Y/HqExUaSBVv6
K+aaqYktl5gEq4NaYxHXdVMfShlV5xOxJBaiHmx12gUJnAfNmh9eafdUtP+vXZ4AnHNRPnhijXnI
Ula023DgrcVDmV36th1ymsCLd/yfosIESUfolj+LnslBJuhUyTotFCvVJpMsUXGSzAtKHE69307o
ezFOOzItizOyK4BgvJ9NeR9v0V2Aa5PMWuq224dc5Na9H/GicKQP/ddu9/yFVbHZ4Sh4dUbTNdjH
+uOy5D4QHMOc4HPbH5DF6nEVKvM5EvGAwbfTbltb8qlVp4CKRlQAMUNLk9EVqBmt/ZUlzguzSX3x
FI4A2vaJykbBs6fWX33JzXXpmND7d2ceNzhV+vuoxtBkO6l8LIaPtun22K8zPu/Pw006WSENMZmM
f+EeoweX0B9mLhbQBlrvTxHJOnfDBbv7gGxk0TzOOPenTnY22iPThQcdTw9dsrF+3BGO3czHKp3K
g9uF2HehReFKS4esELGsUTlgFBArq5NysrN60pBFe332B+KAQh1poTSBzL8asdFu5gAIF0fVc6DC
9LSv31HXDTtfl7G25koLyxppCL7ZpcUdpkrjKQjnJVyKb2Vp6F4D7w3xqTOBA2d9nfl+ZqhkkFBj
iP+MU53rRWDMgP/5mJa1qDu9vDrfeCv5/ycIS8Q6Ws3D265bmAq3ezZ/y18SBOJnIVdYEXoP67Dh
48btn/Tp1D4GR273YAHVZx+pkZaDgPG4Cr5H8ObPRAkkAj6x2mHJJROQ3eerw6AKHl0DZqUWY4OF
3W32wOKb3rdjGt4XQYoASRB90ikKPOzL6bUrGYVOxGJ3J4kjWSVy4QAV4tjr1xbu2eqy5mpUTREx
XoqSO14E9AUwkk6WtoZWcRjteWOZA4fkYq8+mhGdV8ceGEf8A2QJRrlnA7jpZH/R6uOy0hDCU/F1
H7+w2YMwLEMIqQUvL0bipLsEZxP3q537vfkUtirGBnw2iXzDLx69yqs1ZgeesATQkWup4HlM49o7
sRkBY6yQ3mBfP5/yqfW6I/K4MzOEu1gzRm2Bbpw64dpHJuq7qOo2ipKoHGArg4ROw7PnnTd5/2ez
Jy8EyV1fYFVCr3wL2XKeGE03rs6Y7FqYBktDm/Sn0+FFhZ0uhKwcViF+j5/H3EYXZbqTwjCFXqzE
DJym11G/CyyxZF4YpnRyL4E4CgqH6/Jp5cM9mmK2IDn0ehAb8R2QcZLUN6O5tNKnN+9/jVdNzrvJ
ejRFMs/2fI35DVEY5R6opZt+Ih0r3F8ECBuGJIAy/nRhU3IjOFElWh3+S6rpMVzoH7JhhxB7+bgS
jmpf39KkwQPm5koBsWgdnoSrt02WNhEEEMGfiDsq7zFDO6Z0bL0cQ7Sco2nLsyyNBGzzNKTVp3Id
k4RErXiabZGZegkDfQe7pgaRZRGT8+coCEgvEkqLc0yYWZF6It81JiteDKongcebiuvLMvcSM7NP
Mz5mBMGU/MW9P5Lipqg2vowbdQbC4ycuAyiHJf4O0tafnhET5Mh78gUP29b4IZp1op4N/SYUdNIZ
f/WIUxV0Pj5/Il3+WTBITphuVenMfHGSYw687tNrY2i6M7j90UMbPIYzVKmKhRxtxu9fphlyeVwe
UtW9lrELrx3R6OZMpt8bLMaTN5bqXkox2cXdniMchEm/BARJA6FJ7jwSRs64XYjZ8eGpyCkqnW1I
iAz4eLWFOZ5NvVSO8ZYkw4V/Bsz3joAoH/rMSO0nGtHygKDvJQUWu8lz6CwDGGYjgkmn5uOY2IbV
YL2XCDVOCiKnNBK7ShIwdsAY/UE9i0Y+arvvKS2FrBfVokrB2oVeBquzchzlBi1JWpdmF8Iw30yL
ewMXTNwsgf/8H4ozU/6gLTGC1x2PMul/+ioNCRemwfXZWkoxOnWTTVkAvMYPYhUzDRY/1lSq+MEG
2I3FsEcrGAI83ghOeAGhTrbutqbe5TsmMKQfC0rSJoZCx3izsP0X642QucTfEYiH+UWfh0J14D10
ceaPOXAWDRj03Ol9mOa+iieAf1+CTv2/XQGJ6V56i2w53U7FCEKgvfLpJIPlatmBr8BJCCkC8RBY
jfPGbDVyN5OzOIPbU381tQuiIVlHJR0htASPx9pf36wP/rRbo1Kb3NTs1JlCPLhjBHWU3UhCeFS2
zoPkXD3uhuAhEmXD53TO87rpbgKWT13i+v1hbZU5vaq3Y4/GwZuTJ+KbbP77UcOTIUagkL2LfmcK
cjuXDXh7jKdLDABqVT02gSLQ2HYwOAx3HXZRC5cF+ISCbLaQc3wOakG219o9yyOoWn0VEh0umnPM
Kp6KZStzYMg8/f1wJG/xjdzs8oFi5MZWJa5O2RI+CojcywWAS464heDRXxKZA6IUWBL6NCDaUBSY
RhtEqmvHXCkAAnmcC3CO43yffskkT2wlOsP4m1LKsbdNTu+3wF934hzVQIvGf2bzbIjf2lt0Sgw/
KBxCGFRgVvqtel91Wfzre5eC7n0HoJErI2mbiWX61XWZBXNVT9JKrsqnCw4maMbhApQ1ACkvOwSl
4iT5b41G3+uAbs6ACzQccPo4bP5OSKLRYJ7FKemohBetAH077mXBBw49lSlurqzFKTligby2GZQ/
TElvU90knpqFMPInxESZzouD6s6kgDDKVU1teTjbhpRTQee5x48UkZ8+gmnN9gZ6fy85z1+ZRaNS
sLaoymEwfVuexTNYMz5ctrWozlglI+XVfnYO2GSQKOtGBwnkDZ1jQ1C2XeIk72iGcTf71XxF6gi4
thKJqMuSyBE7/EMvkLKhG9soMGiHmf1mICAWjca3MOk+EppwpWP9+z1vYM9Uy2+CbWqc3Sz9qfE9
jDT/ZhyUbRGAo49VJVFe2SOhMmhw2C+0zCJpA8Hp0rn/5dkSkqDkQQTpGhH98yxBzdieJz+eZhoc
a4VC1N4NUg/26BYP2UsUaXYqpI7h4TvdsD59wm2HivQ3pGXsu+Dy0X0wR9lCXEV8UqeegtXBvQL7
Bm9IUsZQ75fYJ8nVCBBBgg+mci3V2s+q3/wpGYRUtK7zkKQ2eCLza8/q7tJhKDsZeBmNlU/tXoqo
ijjfsKQpa8gjAeY4t2pcJ/LOufOP2NK4C1FlDYSFJ7yehn6TP82VgxPUxkS5TB1OyoUYwVUh+1DS
yv8IZiCd6f0jcLaN2kHhlWIMjAbKx7rFFQzXShZyTpMAUfjCUXXyuYSDcK9QglfhBAM6zdJhoUpL
+ufKAFxwlNisLnI6ZoNs50v0OcmLNRYt1tkvl4GuBS71iuEvAYs3OMWs1c0kYzIFoNau7/cOTwD9
iJjd2zKGyClpDW6J2Y0eY7l5GxfdwRP7yziZ0N564FuKwuz5QOnVK5tGrbpmVOxLH/Y8IAQ4L7uy
ZFMSlMzHcSbHtifoPNlOM/4GdGfwxJHilwhzoYs3oi2AUMBH1O7MS2r7MhJmp1skr6WqtdrqnZ4N
BHgdcDeCThOZyHBVcuuAgpQ6Ur90Gi4EmjhiuEXaEZJv8icM5xyzfRtvSPDofAX2OsLiVQlABTlF
BHs7taYZlVEWGmxWYsUr/JQsmzFf7t/7rC/Z9NqLiQ/+TY4RD5QJ6eJfhlyobvV1CvjzfsRAi2RI
qnxbNv4U1o1Di8ksegaBWdvpbROXGDA1vuUUGK4roEcdWKttOxN8wv3ogmpxWFhLiDPVboi03ElU
lkRKRLO7TWtXRXLgHyXZQ6nmRDJ1iwkyNrQZZmuxFShE+nwcpLPVGB6cJi3uF7QSZEeZBZgsslqn
Ya2oZvEuON+TyJEeeA81MeUvp+L7busmngxOL9TbdhRmyQdddJXzG7Eycx6/L5FoqLlFfaEuRFmn
4B2Fx5aVZIjHOR3+Les303pE4Rqgz5zfp1I5yJOz8QWTlSIwKPEPoXcebDemKQfylsbtpxdWfRdf
uL11ZTfH7zVGYbq04QK9W0J3zVhVdDAznK+Q/UpVMgXxm1qbdpCFby0cZbqWieBM0Rravyto2rlY
gqaIkDI4xkc3Dcxd3JcaUM1n6N/ifXIwUv7IOqJDxChsOaTaxYwACo5WJd09oTrZBUrnpV9ufhbZ
UlXOA6rCoxLFOvW/xpIYsjlAJj5pJiH1rJq+Tdr1nMcU12l7sMNWBsndaO6vUI1ICQy5V2u707vV
8v9V7B9gzbyXiISd5MAXAL2OXFxhbn/foxYt5w4mmMaB8tMEbtADVOAisZ4SMuEiWW3RjGKncUBg
Dr26Ukch1xhOU21Md2VUuzWUdu4uxUhINkc1rc+mXl2CeEW21K7XPpMZpVbkRBUVxtZ8VGqpZpPL
vQJSfgQ+PSufT7sFpiXaUJ8pKgsao5fqA+YFZCjZoebp3nOcNCb9NRjCJRvNdwUMNziPR3mS/9hH
n6kBy6HsVhuniIJQ0TlEPL2B/IEc9gpcycqlNULi6AXwdzwBuoUHH23E4YgWLcJUqJxsFcAfqX8W
xrJWQs+z1Kni9LLYRYQUQySDBCm8Tf8IuSzXn3uML+nYMdo2WeFj/4Ip+yTvs74x/yIO2crqCFPg
DblJHZ0TQgW4bvY+l634nSLIN3GeSlvrr7BeJXKbsXfV5EDMEJGgo19mrMCtN+P6SOTi0kc5u79q
Q/S71fa/XGvkzdCwNSglMEF23eAQADZ584GeXUeNIHfmaIjyA2rruesMscBweYrXJ5aIj56Hty0Q
o6NpLQuNjyAfH0+0wmObnW/9IVX/Kdyz33AA1BhH8zpZqMJRHBhfzOb/c72EYPSIvKtIclT7kYGg
Ulo04YPZVkhNZFCjE3z92QFEC0H+9BdGWVFIJDZUiowdPV9LoTMdghgkewZ1jbg1Sq/J0g6eeifN
ja1jN2fK1+FshmT9GLFtatNSTody4SOlleavZp7EharzBzFRo4v7Ft18oRSNKIDFNFjySjm3OEcx
JLP8xn1Fn9MJaqGK9ahfYm/SrkWbYRpuCfWCcW0HTyj6Qk9Ejzs0Q7eOrHlxWHQedyhfr4Ao6wwc
EmAb0JzTnOUD7OwG1J2OtStdorV6JGDn3j1e3X9wdrTCbH2jZyZaLajW2FMNq1C6moJUai7fg4KJ
5CS6tWeE6hFqf2D69Scae6g7sFiquwZICYsbxqNBZGzkluLBMlH7tqlU8MObmoQ7M1C9FEVm/Why
/0CelXZvmrA12EGHQaLHPr6Wv3AYtxO/oe5pdcz5glKlbDXLJFwMwhSbTuL72+v2Pp3c2Q/JTh5i
ez7WtEquIN1tmjGcWhtkldtfWy2HBubsCoG/rdB1xMGudlR6v68M7Y9Ks37WlL1nJGs6M9DvsRUS
1rWTJUC64Q6BaF+RTfI9FAQe7zib3sbbUZ+iEeVbYK+kD6XfjJ2Dj3JsD+o/VKZEGBQjlwMhX6lE
ETL6+bwCDZVnpxCvy/lS4glnuAtO3YvlYU4jTrWeZooaOp2Td8Hd3f5MGmCJZiBivvPcj7W0U9/K
rZtu/LQe35bG40m80vrHVLoodxPO5SuaiRUA15rxVFLSuzKI6dhNy5g9K5rJi5y4kJ5Cri5q5DBf
p3g7cUlNPRIjN4NdwFZjNqHIZRWUwm3Cnb8Dxw5jja3ka6r6Gg2jAqrURKeUnF2UbxwKwifC/Ttg
ZfHnef7CH9owQnZqNJPh2yJCI3QX3WxKciHXM0+bNdpQNIR9iORBxlCp573zw5X4BrM8zF6A1xad
a8hbPwR5Q4KdC61ybHsPnG4C6MNrdx0c+4VZNuRCrfDcPaKbQqG59W1fCBbm/hKT97XHBhEHQfXS
dLdpFa3bm/sudcffiI2uO5gBi8myYPQ/ELfbk0VlhFki6RE4rf0N/8IJ+R43IiCZTpBKAg63iOR2
s3rGcKMp4qRNDKPcYGHnbQ/heixjpw/r4jcRL2UYfZz93KOkn4b/tX7woMmxBg0ZAWNvAumJ8sqg
H/OAc+lvCPo09Dsfop57pQHfXRinODEDM5IezBTx/MNDdMSZl5NoXUogpVxvxcAxP/G8YMzEgKXq
qopoeKuroCt7jU73JBa6XNGPueCo3uMWHWO40zkL1fVFe33TtC4bY1BmcYaE87gQdRRp2JSP+lYP
JZyNVgxMitF3LrkqcfGaqGagyNVKDTQexKHsnAbBOXtPIosywwJH8BU02I7NyNMgPiPFXKjAj+U5
sbhrzOEAweb4tXmvsddGe0zyQoAwPyLT7rQaPUavYqxuKx7WHZnFVJIauVIMVDLJqc9Tgl9YiKdc
BS0q7s7J1Df+5m9ghAOrixY2H1/QgB/tejJXZtzURTU1ohtlWpL3vS88cSvx4DcbwOt/gHYr0xIY
cn1uXp1u/I1vSVRrE1PEX4M8JG6VPG7qUK62TV7uY/TGlzr9bgXl8IGVuDihvLZxYl2FawJ3xfU9
VXnlzvwBt+xDYw6SOQ6jVD/cFFAOo5LBici1r9+qWq54rdFPkQjOolAACuKy6GcOwzfSr6IwlvTU
7wcw8gb9/wW6A9ENrEMBUxM5ivZZRHnjiNtP+1Rvw757Qbh/0b2qAMjrmeXWvj8Q0fZlfSQvwSng
J3GyYwq600wtY4NpbW+2jbfSQWc3SWSo7Rfhl36w1UL0EYOHDTuWYnSdvlaf8ddV1TWeYvmZMcmY
FMvT5VVoJ59SewbooO/WAqwDLDAb5A2tfYVL9jxk4Z84vqb67krbD/tlHWuEfQvH5+Y/BMjhCo2V
6sQyVEeret2dEiY+GOPd+nUsY3Xl8qFYz47hTJOZF1LuTiro40mtseJHC7exY0+rT5SSvxBG7G9s
wfouOpgId/cof0ebAuoNfc+vAmcXetVum2CKtmRZDkWAfA+olQEQPZbV6+K/Aec/ZPJHIt8FxIk7
xBomO/F8c2TJWh6Cum56H+BpVrl4LAAzsituozWCHhTbXmElIVcvWE5EmCUfExQCBpSYAUX65exm
ACbPuPJWn6edigGYuRx2C82rFSvdKfB4iNOi2XyKs0qbbuUkQCrv/GzRfgGHBdaSt5Rs56KE+vHo
TwF7/SMQt9mzXUSElb1EPxuDMHu8kcFi/SeTACMWtfn2eFPT6caDNApRg4STY+oG9E58e5At14jX
hx9NHWZkZQl5WU4mX2tv+y1VHrDRTra5bTuBDsBlOHOPxvkMlxWr4LsZ++l82n/Rol8RMKroTO7g
PsWPlS6JwG8JSPMRybvMvr92ZGM2JsmrD0G25u2qLkCL4/PMnFwj5cetPFxLQ0ihhBNXGksJ/0is
P6d4jd5M/Z45S/AULgq9WSnVzZIF41M9GHe/vjs+8a34JgkMNr4qGlSj6Vw52n2M0jEA0eRTjrat
Z8VGftEsQrCjTPOVtC3FrAFnG/gWLttXHbkwTWuoUKtK7KzDEuyAzRzwPHQMtJ/NEwWRjyjyyfyF
wyPhGy1pOXGIP339WBrHcIXfadVdAfCC0kmDQKQ+96nc7HvVmGz93+bbTChsudjI0sHwtv/j8D3I
s8tCcWlDvsGhAJd9cLxpMfA2sDvmjJmdTXRbSkZoMfVfl8Q5aBb1qRUxYFOk+dxjVYTibPYgp1L0
Ba1WJ2lU9+IDvOJHojkv52xtasR9Z9sVtQdxHPoqO6bc+YZYqNJswi9LSAHSt/LuMogB80WwOihF
E2eU9+i/Or2fvyySjiFXem/yIWJuqKHcU2a72/e0yXx5+VVLd6e+WAlj3ROoowqj/qtx3uU1DqY+
2IFOYY8tDwrkPkzAGw9OSfxiVLOtBJcutAcTA8BqoIGcfeoMCJQpNV+efYk286cvC7SeK3tyizF2
XBGXiT9eATvMx1qEyaKxJcdlIFzuiLD5JVHlqyJKlN/eZw69LCHl6ynQwFsqkpwm9vGCinb95gZz
RXDMqS6J0ge7yC7Pj/U57nHTS5zbH7Ox2OpoNmqY/ti13xLAmb0MaharPYJJpmBhOTBlcCBTYYl5
BjKEAJ1lPUoCzNgoDEKFfWSPwQHb0+EFUQxW8a0726OA3MFdfKfYNmeEBtYs+OzzCXsIDGF9Je8J
IJC5A0mOZZ4JIZfwdQLE5kO/vMo7IcIH0Ltu1r0DEP1Nxs8j/X3f2+imSKqSWj04nDWQa5ZIeAgh
QRUvccUGQ6880j7+f2uItp6Bqtn1uAUrwvbv4mprgvdPAEhLMKambToRLrZ6PcEZUSg0mA7eN8Ao
X0MosDcxkhNrLxmbWiCUQ3qySJ7a24B8hBtjbr2QOojZBqDB30SLsRx3HnqcnNiI3ZfA0FK1JzEv
Vb5AyMSFO0LsWoK8eSh9cOYV1d6yH0QhUlgDAAM3gLfR/2lWVy5mvlCVZm1MbKQCfrw4QYar7QwY
J/x5U6hw1gR3AOoA60SzjOVMuykjfcN18PxFWiNvm7bfXka5KHvzyQRJYXf4+rmZigVGRRsGQzGq
bG+1gMbXWqZi8NG+GExldO8Sk8/SNThguTY0ZwUA+QLbY4SeYn4cupipLnk62wlmWh2SCoyF/E7a
7vVUdNyiyGPCvL1YD+wWpkvPG2Z+vWmUAKXdz6WIZV5tohSZvyq0D7Oglkv3krsQa+WWRUk5nnXq
fL1YRmHnWpaH7cjGh8jdEBTfpiHt/JdbEb3sGo8q6OZI0ndR1EictodY+2YLMIDwXikdrNKJc5Tq
5Ijde8C2l6GVcms+3TQnjYEOwqJ5LLfvkatiw38yKq1XxLiCiURcSaBjbfMXKePxH9/US9rD2sc5
a2G013TovLwl9wYSVXarluvLd1K8xqrejhTZiGJOGKOhSbxTVAxO0kuz1UXgglMTuz67JCBoqukO
9O4pKqtXbeHzMiKr9FhkMevfCRHJS+zJnPcfipBfPxiNaNlunjSbLw5hlPE8oyEjKPJTRNnf4Rjy
kZaRex9fP4IQIiKsyD4mmyi3tqM1S7csfOA6gxNXktRbFksv7xUSlfwL5WqbAe1NIySFfi7scpdM
DTat9Ty+O1fr/Fx2jLBAcj3k3M8qrdCtG2bzIsDcnZtv1sc9KxVQajv8KoGlHY3/xfFVxAtjar1F
Xold6OtIEXY5Tc0N1M6GjMoTWYrJTg68rzEEV7WCryc1niO+HNm1/TT5sHNU+aPJT3EVkrthCgob
aOTTyVxJW9NEdOIunictAQ/Nnz42de2jLARxGUZuwK/y295pKinH45sG2tyf0URDb19YlbUlolR1
Fi0vkWgScz57hw9vMtuW0EuzGWei5KR35qJdlV7i+zqLH5poeVFtzc8OetvkQfciESmHXQD+eGXJ
pzMMxq1F9m10H7Ns0D0rhvlklApTx5gApurWa4sw+8JkUrJ0si0Fm7Yyk+SZ9nES8DakSoYI8kC4
6BjMJry/xaAOa8rNpZIH62zVBbAxSxMOltcOVAFxFmGH4+tfJ+M6Nl4xY5eRGaPoYuL9euADJ9GQ
qzPmfLAhP3fEQQ1v4pj9jY7xMK7yityoffJhJSBnXka4ALjrY8FJIF1gUIAT699FJ1IIQIk8hgN2
UagUOKjaWjyGRVmJZVlH47eoMuSwPiOCxEqsDcFBJJWWsV/oE6W9MK6yFUqnGA5FyiffoLr9/bVN
n1Wylx7cZ9mtJFq9fA9ubQs9CkzdUrJ86/YtKIhUQukK6ZGq5L9OVCMk6phy+xuzB+D8gTeknTzp
OuXPh2xkRkHKTUDXMPK4+T9RaWWQoLNVV/BMppX5dKJGKBr/cUVzl/SGn+Eyp9FIj0GauNibSmrk
15zDuH4P7IA3Y/bMsZfw7uSb7BgZQa6D9vBg8jIFBpMmOk1Jfxwfv4Yk2FxQ61EW29p5UYz6VfS8
ZYGu2h5Zx8iflVELZrGo/7fuWqJov9p8FAtSmdzyjnQHXSdOdOOEQvUky0PKQ9MMA4V2zjV/4QMx
w0fkpwwFCzpK7WGBpmvwJ7Bw5A4bQEhKobNKVGEa0J6j6ohSukMJYlGTc0MZRw+YXutakUKDLiO4
Yv5befBrBgukQSWKwZ13vVopJXt+BIhfrm+uM7MyseUXPlWKDtnYTJth2jKOz12bYh0aozjcDXKI
l4rW/ALw0aR8YWAU+UV3F6jd7oW0rHVJlCdJMwWbDnZYgOYSlFnMwq/pG3mZQ7OR3EMVojyPc4wt
g0rdSBrERINCaUYBNg1Qw1vH+0OtP8wMsB0BOThXQvJEEqodz3sngj8qBWs4TvGsfl5tc8p4SxGO
lrJMNSOyXRz9PRkSLofkd5LPi9lHmVTcmnAo1L1FAqo8KCC/qCU6zMscWuKe7Q+5LwyX2OF1Qa+s
kgrPmMfx/RuacJEfZYjWrtnFIZ8XVnNj3ULz+5KJttrVJcpBk6rxwJDO3LFeL5+mhG650QscASRY
cA5vL8zLVOb+kVpk+DxDITceY6SPYFGVV+3sB0P76k4+uGU0Y9AlF5zH9Vj1yohx5/DpqlsAoaav
FSw68eK4wvuUmNxTR2GP72haaY6/FRYK3F2ZKA4zfo7caHAulFUugPgvlxKlWKA7sB+ENKXXfAls
onH9gj4mqfmiGPhwDBNpyohpCp9MyW6zp9qg6NVJKisMIdLiCOp9teYmwJgk4d+Vm8yMQIZqlHGD
To/TiQPLyuRK6JRKAAsYVoUDC6VKb3w+4TCSyFbmqzm0+m/k4AeiZvNU7Nq0t8xGpkN2Wz1cokqP
8w9eelWRFFP6Pl52vgBQWP+9p10u+/HDWjXDYCwbaPwKsEPLGza2WEqgIUMvhNtn2/Tt93OGwyM5
v4IEZsHZzwxgMip3solJC3pgxQ//iRDLlqZSM+0di/goUr0AcKlaPlImatm7NHIUzmqbuL2isJVC
Oo5op0JEeZCjTQ/NTQBPWqDj3EfAHgTvviO2oRLUSZ3h+hJAxRXCqejeq5csi6ceVzZE4975uwC5
ThwImkUAU0RUjTsngNpQIpzRgXE68EVYF/jn5CCGhHz0dYuDkmx6TUHoGYvJTR9cEs8YVWObARAT
InwiYd3X4UVjJb9RC8qAnSgzDJ61WBsDeXeoE2GzQ0wen0fzRxuMM5wyrUE+xUcBHbGXuwx7vdtO
HvhTTephHX2t7lV/DiVIyvBHno1exh46sARSTHX1kKRvruhAk6rjcogtmJPIDSzz5dIj4i8wfxvy
W7MPPpDro2s7B4OOp2Iy1CWO53976nSXGi9MyQkfQuNoubv6jWbjDFDrqTOTtlofrClzNDyfYYz2
1YNqQn7RO15P9gUc5carjxFx2h+HJXxYrDL0jL66DyObBoQa9xS/U4aK5FL4Vj0ChGgNH/jgmNs3
0V/xguespXRzJq1hbdM+OqO+vIgaBDxKnT4XFrunWnY62XO8eItAKuF8CYy+DpBOgQJpbpLAGcPU
opN5MW/MDbMuF98vUulcoJDocBGlXltVxCYlnwq6nPh6csRQDwlGYLPBLxkamuSlodkoWvH7omHH
HXPx3/xWNTKVVJB4Y6iCvgdGvOkOjlMG/IT4Isntoraag+oTqSETgvu0ZfniI5XJ5nJ4NgV4pulC
SycZmfB2O0+ak91Oe8it1RDRvm7J1TWYC9BRgHeMP6geyLtVbIpMEn23FlB5FzkPH2Nh7iRVrVAD
AmLzxFRs8UxbOTDEdLbsTtDrQL0GCiWiTl+/ES6+Eqf13vv5VQ3zsMXCVp8VnDP7XCmLYD1EmLuS
c8L3i3qUXV4p8RhIIBIHZjZYqR5S1hDmNXTSXNbSvNIRSyISlm7bJbBZ2gMGXFqvcJ/na6F5AJ5T
tn1Q1MAKJE4hyde04f3WczQXzlRqO9cf4Ubsqget4I3j2bU38BB/8mTBGhkFMB+YzNi0G+MQ82LM
ibCwmng/TiZaZppA6xdhYQ+LwvDs5HanoftgFMtDKS4IrcuYF8kj4yyx9XMqhrV8Z/5tBkyzwZIv
42/e4EGHzIM92NiyaqqhcseDyPH7mxZHDAOOvZqsakqrtiCqa0wYPpBB1Cz/ZZ2ZeFSqIALMEFLy
totJyIAKsOp5wpbgZ2+/KYO1qrikjyXbYm4w7rsl4yd/CcQCEgzYYX/mgL8X+7IRpM7Z2TgCo4yg
ackIJam1piTOBQGvzHHgrAm5aMu6c9B4nVI87pGAwHhH69miT8S8oPykj8eRSnq/1lx1LSLUOgRB
rlG5UQDSnRe1c4awbZ3rdiTTnkYDhQlALhIGN922n+sdIkpWVffjmdabEYfDpzN1MdFQFb757+Pi
rbm85q6OOyfQjNbtMNR25OKV+aYFETazFOcxg7njS2UBnvbui4rYHwN/7bN2bDlNZ2qYQEpE/rV6
tZHoqi5WkIcdqnXzxoGru6MWwzF9gfaj463TOs2yvm90PUQEu6nB29KKgNu3OK8CqPB3stqVC4FQ
z1auZY9uRj/Rj5UttqcAUyPoU808GCAwE6DVGDLp5KxiiIqKAtVVOYy/3jE+BV9RaCeiWUUw/UzC
EKAzY07KHBBT8REn+ICaoUc6rLwMG6I0ogV/0XKe7glVBEcMskovcWqK85WwnfykzpJx974Nk9mk
qNll5YFthEVTX6zPXRElyxx8P1FmpIqkQ1/8EK3aTElihDkwbY0EG4vVxBAdF0i4hlvLBYp5y8+g
8FsbzH/qdrWRugtE6Z1MxNZ6nMJTpbo6zxcQ5k2XjBbST9X+Hx+a7n/sBmdAVW5hTAsJv5eiadi8
eTUpgITKJGy8gLxMnyIsIGA+P9WwT04U/Ve6TkVxtWxeGiAsWMpLkT0+5J4Y+1Whc2PGz1/HqjH+
WyRDo9hRBfYhjWEu2J6WvyUeXKi9YIwJiP00V1gK28xjyTMGX8CuJWl/uUEVLypSrX+m+HRJhV5k
kzk6WzAIXeyBr2IAnuKPS0jK82JPOKoQ2Z/l9Z4MLvdnaREOzU8v3/tbEAt4GYCwIieu5nTK7WiY
d5SkJAIW71aAhCUIo3TDNPtoTvzu2Cu33evJ1Dm2u4FY5Y9TYw1gpombCTiK/w2kju9FRj5Xvp+F
fuEeGaUNRofYSOuqv21/+Tl2O9w+auiVcNuFput6lwpYN3QK9yxlDzOhPMora+UC1+PrlZBKuNDB
hbhasc5g9sps8FjYLiFfL1vCu//+QcSgvdNrBVfxHNIwnGmFbmRC/5NbmCKj1nGCanFrlFfB+FkB
EBpy9DLlyqUpRrz8JqWd9Zwq7ze8zLi+54BUfoj8a2HEUuXq1FwMJq4OrlmK9/b26FIWyO2WxCuo
5gpu6bRrJ2+bwqjD/oX2VfPClFYk/FFPe6EQ/UJIicqrsIhKoVYJX9bhYjCx3+1bMFdjZI5suWsw
xlTwH3BlK/D1FRyYKA/FrcIsIY82RLcreB9kZ6qv/k+UiWbAJWDRvDRNYofeHroF1ZjdC8JHBkMY
Nt0CxHxPUy4tXcXg4crCdSBhZA0PswgebPCFxNCKREw3ADcpSL+v2JOsad2UakwzEFTsXej1DIJu
O5lz+/AKbW/O031W4ybNFu4TArkFN/RsT2Mkle0OY+f8WOhbPmWFoeNAnGupp50+v1JbstBjilXc
g3WuthJYUEg38X6pP76jVkLDwweGwCKs7MH9X5Ng5ccaWHgtwAOMDbTb/6w4ZaX6cF+IMbof+YfI
Y/XjO1+EhQcljJl+KL9HGPV72AB/cMKJTzjNdPfUnPflxOQQxgOsFgVXH4uNcvLBjvUN5rUeQosw
5uTKpGydbJBiAiKVcLdl6yytATTa0WV6yEH4ZJQ8TQESu8SDjm8V7/mwCWpcriHy1gGtpcKpDfQq
i5GgNU0SNf+xNFVwKlUBPgpmX/nkOZ0mQ2LsoT4ylGR/EVo5qSbAgs0gdpWiBoO4dX0w/WoQrxwA
IV6sGF40/C6EzKZucUxdvnkr5bke86dz4efbvSGXGIaIWcAF59SFAIwxbFjRQ6HMrRlnKGLWYWNa
e+OiieLQ2Et4JAQQuxSR+NAlyhWZctRjh7uCR9MdbE0dYL2tZ5wq89tEK5DJHoWL+Nogg3OSyKGc
O92ABsExi/5fZqs+w2sD2/XzmRFGJSFn/FdaXgUVztI0cB6u6lXggvwGZxzPItdMHA0IyMrpHqMy
cJ14nQdR10x+uXMdlDeYdBmbX7KkcnCYpQIePwMaXcSYgD31ty7KTfjWSdxm7MZpa1Z2Gogno/G0
wdePlf9ol6Fv8ZvaPYT1RMEkR2v8iDKJQJaiiE+tySo1lgUBr/Rb0j7eCqT2eqEy6BXeeJWXeHiW
8J42LVgAu04VhLhToC/SbXPcs6MuB3cQjt8d7v666EnnWUCpYzydTz3lWuXOg11dUAMGoqt2Jtni
cioEIRpEp7rfQwNYb8JeVd0Gi0g/jAzD4+4+Wb1b8uqk14r21jHWsT1EOV+iAZOwnFT/fyFP/GIh
RNJl+gpwpXDESntK1J+w1RsobYLgiz/0f/0vey/4e6yL8KVHl7w41XBBvihVqQXB91NwmHYghuSm
jFe3/P8VERrWDK4/LyQjKDT6V+QF/nMB3HwtR/9FBieiz2lOzfDr/tBVsuV6rnPAZebZuif0+sYx
owWZ8bD1Y4u265w2ujG180EZgfKZ6a5gpaaGfzwLEn+NGh01JMkjTG7yKsqTVCPYpyfKyoDO0v/l
FzBXXvY+z8qH5KPChhM6Nw7KPrPbfCfpmCDYNJM4g+tJO6Kmxu3vfR3+u/EO9U2QzVtLT8Yq1J0o
x0NlFH+TJYtHpd1oE+jY0ThMyJ+iH/ORjotSbCsQLc5anWdcsmulzIfNApjdP08OfG069X+KqWNk
REGZyvb/rAYI3ZhPYJUe20Z6VCKWpzuL5vHf3XHnvQrBwgPA/2fXApeA8JsxQqUy+B/r6VMTXmrD
EDzM8KepsHhmgT3FcO4vNSjEfOkIroxC0a1B2juUfAZ2+vOAQeEhekGXhDvEVsCQ/tifNuyXEHjP
xJBbwlYzK+9QE5Gigv1MHsUs+W6Tx8hWvTuazearKQKUIwaBbaEGqdfO1MrvhAVBlzE1jSupHOBB
rvZeoq0s7sZonavNiqLgVChGGm2709LjFPeEYwfjkL7YE3717GkCekC9jynKRoVSgcKHNF/5p1ut
yBfsbm/TIV/n8fi9QbfEk5ricGhya4ZUf5bSyHsBoD6PC/ofkf60hF4+fgfGPSUP2UijTBcXDou5
d7Y3KfuhMPKm9jF5mtLvCFAH94Z9LJQ03Fdvv1keGnVfGijaiJyUmZjaF/ECBCYKEp98xgao/UK0
R4kuKIfTdqh1+g/Z4zq/SFYAerm32ARnAydOa3bTW77F+rN0tP8EtFTLDm8akxkQIkrIvesjcYsj
ijmYaaDD2ZZa5ChpTrC1267aYX9iX4eSmalmU43Z0q/QDyctERxsR4MxQ9BjoQoQvd/UmBKlStT+
B3B9bgz4X7sZY5V7Nu4Ef99XXUJs+hm6Fnu/x0cT1921bssazvTfhbOANLLKDgxXOKJhhrJbg3Re
vig0Xw46mDeZzPg36Ab7HSi6SJkKpQ/ZCjXUm1e/eUcmEGHJ3r5N6djL5eS/m8S1NWHQxpifX3hA
S88loIH9i7x0iTJkrSFxwlPCVTSQDjArtbGo+/G55L3uly3maCRc3sLoo3UHR99uj3LH/DClm9O8
XWMPxEpKTlm4myhCEfUZ3+P6cb1vF5wIfr4OAgfBosvbCOUGTFNVwFQzJm8dPyU3XlNJ2VAzi8aP
zlDiv08oH0SVHgYn+jexUr3qxt5ity+t2WotBnH8N6WhpsxdwyqTp86wb/tHxN+RHaEI9abenUH7
v0bA0x3Bx6lJymkTsHBUOAQT15aiAGq3xRw7zIM/CEL3ymKqcsedIHQHhcAsJPszsrGVq+eC3J2Y
ov9kgpflB10RYBEzdsHLd9RBMXtyqXurv/vUbd/OWDM8kehzfgWf4YpB6CcowvDQ3T65Q68POo/1
EXElRwdGu6WCfVtxLt0aMAhcy/SoVFsxqCL/EI0HC8rry4lNuiNoqGYbVVSeK1h4TVZWbVTENudr
3nP0YFjDrj4MBbBarX/3FfN/miXy1IzGTtbhwXiTsi6UBwK3UkfbtU6ul9xjm9fnlc1JwNkpeeam
v7sYSUg7sc7dCgxAIKxt4VLoypebwP7Tf4K/d2Af0V7RKkVJZgADUWumGiGjOS49ukjObQLKfJce
aHYq4iy4DsvUd7EBFDdRp0Q9rTv8kXbW0J5pDfhIaYCZK1femZVYPh6N0D9cdATc2ma+8uX1VIP3
uM9XXWUaovDM09w/htacKm6mE6Tkc6fybXcQf9bV+WTbucPbX1+HJjZzbIz3eHkqpeG4n0vY6J1g
ifughciNsPRcIfzU2QpP5HdMwkJDWXPa8vjOVM24lCSvOyVLXtXS78/cBykGOMuirfH8v6HOPnSp
Y3ZBVBw1fIv5du4B3DgF1MbYREOxogzhxCDWceDrnbz2yTJNhZy5oRPrxfP0eTQW4sFmKC/ewg9Z
w4/1HcLocJpEdwCDjljK8g2NBFsfKGVNbAYVmaxl8M64VtxFFdjUSuwaxLH5MPCtF/f3ePCMFHP8
uadxm5iMqgAVfICfX0EaXPVrCIvd2eNMaHpWgyK2KC5UqMTi8B8dCEL5ukHDM2E7gQc6RmwDIhxW
HskZFHWuXhh0jlrSwrPL0l0eaRS+1MbkItmVis4V5X2vaY1OgqQPpIh9mTLPOVRqcpbUxH2+bpgP
Nurt6a2Yz9wedaW+TziSnzGVHTwpCXXqdShSgE1ISJE0oJMO/CtushES3OrdHoh4Kb2JY/gq5NKu
1K1AnjSKRhq6EDeEDIhVNppzZ6RWgt4ZsfxJQM6/56CeFvLYdH8Fq4OA/pCFNK4TaW9JJJeIU/PB
5d0SiaG2sPBlq2DVTfaXn6SmrfhqarkNv0oqatH+4uXPO54OIVOmZK3EuVDnDU0apivc8YyEoHr7
w9WjOWUyr+fSkrq0Bu4veihg1zsc5eqQ+JR2L2WQBf24gfPsjky/5lx+kNrRAdz8+6WwqH4pQzyw
HjhnV5fOB3djKhgI9U1ZQAXPDAmUomYMyYfjAllCS98Lz9+3tIYQcqyihMkBwTGkU1WXSEddSPi/
/H4G8HnkGtLTn+2cOhzQwcF6qqFysDmwG5eJo1ni72FPnkWmIJd9YoPL3uTjLPpeoW19QT5P7CmR
SqSFaZvvkY9izUAw/X4SOMPdcL4Br7E9NIsucNDJ7pDh3Ga0FDL8qziVEMsVCvJv3EhYpgRf9zxs
qkd2iUTllsbg9kua1d06cNFHbfKA0ekyT0CGX4TdjKmMAcZOTZvDIQzvSzvp+7CTVjGFwQVAzhqp
mxNuSRMzqalUDZCENlitJBfS7I16OKMRvU42A87y6qnI6XA5/LKTpqOa7opQrabe7yVc4PEiaKEe
/pzHkNLDNsfa3IQavWNYy5fRj7huqMt0BEYGkXri5/gtksa4EMmpsIUSDX2Jo41D+x8cqL8ybD5Z
YqrUFPjoq6pLq1LPl8tyyTYdiF2UXQy0twd1/PQGooDm9cioHxONqRkLLxtmYtOY94WnPno+RdnH
HJiD9bSserCZkELzdUfnmNaknNF4esQIeSlXlIlu0c5CJfPiYCrNx5JVJdi0pqWOaXXmvT9hRpyq
zqNpW6xlp3Wr7UVbXR7BJhP0LpZInfGwwxwiiwzGNS6Em1KCyeL/MShXvwC57QP0YI/iyUrZoBM6
PXz7i9pYnntcH99FwLLrSPRhuVZdq+OkatBc0WSmmNXMXj/rnbPWCvg0jYEvgpgWzTCfwaLPDqqk
mcPNxb7Swwws2FSNvWZ2x/O8hNrslihHzXHnM505IjTyL+uA2Ghyt5EOlbJO06UbjNE+Pv9Ue5ju
zr4myuojYJ7/3DVuVsVvaC3hVb7jBz+sQp5lRlb/58YHM3jyiZnnHq9UFB/P43Olb1cPGM8wX0s6
XqALZVKFYDYqIcE6PNowQkx2ayOfh10Eec48B5UV+/1peersTLT4xUEbjS7KENxAM2CPl5BFWI99
LEsWZ/AUv4lFVIX2RNLjySodfWsBcjH8IFWXoEmZ6QZig5s56FzT6QDNHk6nrQAgzjscLh5ZxOPi
OscyFKKckQAkgQPrWZkcWccsJvR7L6ltdXLizhtoKg53h9KTYuNc4qKO8z8C8367mqwUvwkFoWVO
bmuvwEm3YE83SGCzuzBk8yBwMVYyuPag71Eak3C/aXl03D3P+S1uuSc/ORvjfn9JoC1flCaQdmfN
NdiBG7aIWj4voXX9geAJk/lO60RM3Ql1L/h4P20P3N/dM3oSMjHILkB30yo+x9XHhL16ynA2y0k3
CgjNuXIFWdVNhThMGo5G5jOsvpqLB165nutBTjOO+sLbV3oa6pMzOCn/nUqA7IQH63snsVhisy0v
3zrMR/kQNbtyVe5LFpH3RDLPGG3x8RIpujyQHPwPMG2v7URag5mggWFK/5C+AK0iKL8vTLCLhgWL
1+FR8+MLy667r8zx1HtheeZM20C4QmkaxLTiShLAg48Lw2+2i1Y7DN5ERe0mcptjM8Xngxdkzjdr
VeMGPBAxc7oR4XjLKa4IMcWVzadDcuYddP8sNNemYAC3POWwakwg9U7BF3k4m8x1XXwUztHWqqlf
gTJVq0i+LdUqgO59cl8hAVt9yTpjl8wKl7w6wXYJS4HFGSQghuh7PoRuNNnyq7YUxQqUgBT+I7Iv
mZ/7ru0wFwo6jbTpIfqGDzih1877FDssx0yG4kWhiJiGNGdFD36xmdYKkqmOZzV8qeKe2nQWDWD2
Apn5EnKAvf5Iwq9hS86ngvWTYucXUyG+CMe+KF0pQcIO1cpPo2XpQM8uHap/rHLKdv9gt2LrTRM0
4px/iPRCHa2M8k0y46/F87+hM8Pg9DRRS/NlEQC+LXJBtuaVOEGmLBMe4VjyJ5dcgZltQJhLaBsE
BX8EBMV0JY5d/zrdBHFMq1/q44Uebbq/QMl3rMsgN86Ow4dUJf0lNlByIVaw5XCGDt3Nse6gHeSd
yhNyZpQoBPCa/tRXzdHqRmDhDO2rXxw0X/u8LTyG3Q26/POTPiT9wrwXqe+ofGZ89OR7UMa4zNrz
h+tC9PlGBPbtezHFn03euT5b8boFcU5NoMs6zKSWMvjCd3cg60IPB8rzeIss+EBzjTkBX5v9I2Ku
lHhF2IMxc+gZeRIQ9RXhmqx46BUg+6oPLXSPozyaUDACjL8DQtySbsxwgJcKQHa7ur15o2l29Y87
1qll17FhG3HL+Z1iQBKKl+NXSohlTCdmsq9P95vh1q4Dm6+1TZ96NkaxgSPrlfRrdPeU3CBNelQp
SVnodvxcTul5gCveHGeE8eVPkfaJvZDymkB198XPaPItJI1eebMyJ2wQjvAy+jg6NDLxJUuexXkn
d/S3UAntp66gWSgd+jqwYff5BjUMAlEep+7X/+pKYB375+NC4y+Bhfj5IdUy6degJ2hqpIXMiG3E
+dS8yHAhdBzxk4WooVon0wd0pDuVA0FPsSOZNKb/UAxCH3lPE2voC3xbfTT6belxPqr9w3IC2Lqz
EsaRQjf4zhbWs4Jlgv7jvfDnM+UcZQKkF1Goib6CLq4E7F14fTOMsXWAWV4f6EBfrwbw4YASgmOR
Wvvwy1x9SpjvrP1F6v6tXgLpPEZdoaxrDRCxpDD/c5r8zmVulvVheLaLdeXB5JxAtXI4TkAZiCRF
jKndSO/VrPSUwVatLgCn7W7rZxE3GTxqYwrGeNR9ZvngXR01kYR5/rLutN7DoN6/B0Q03KUB4L7h
1a1xVsvY/SudpKQVvdUgWfaPr11QfclZKmn8GWLSYw/SnmuU7qmDgFf4Y8yCQxCY3jtvMA4HQ67O
ghnIIQqzxxXCBb7OCtyKAS/9x69V+3js+2HGQDm8RrsVWLMlMi0Kkf94jqpB9HBRV1wPz0dkuEwL
chJGL8xzntVkStbN29DFhpuoDPT7Yy9riEc6/6WqlqkFO9CT53BGZ112TFC/5+bDodfn9QyuGojl
YEtQNdQRpHAp6uw9LtNr+l/VlKXG+kor2MCisUkeG4nhjW+sdUOJFzaPsVxNJCrDbczgPRXJkOvS
/E0YFoSZdqXprVDPyMU7tbj+Ed9BjttH5YBE7fERxMwlTBVikuNwOt8f1p8UbBsuEH6J3KfG5YKQ
v9sy5xs0rWfx+oK+sl9FFFLw/11J9vYl/TgwnZp2aCj1NwpVI7o6J0zFhs456ivHhxtRz40PFPit
3f9r/C46ogQV9PxZ7s7lxvdO+ZLj8cC3ejlkaNtzXFS3H6dkvCr+4WfIGPs2WPZ3N/ngxWxbOF74
dsD9oeTRZzN7WiX8YKVBL4tr08lwWolb/lQu+LLxVkAxi0P1/+idVCkBR5zxjoI6ZTet18UyNtPk
P4QVs/MBp3ZYJxnduPdLuZehq4Z8eD6Hps4MI5+GfSh7G1bZ56bd1PftwFcXp8XcqklS7x7XPWVx
ckjzjRHj2wO4OgCeNcDArP+vc6V4wi18WqqhIED+pgklNaMszmv3n2JnXINp87YMkta06+GdLU52
+5CRZpkEkwsPp739GB9uKV/kw/4lpMWU6fICuA5YcduNGjsT2Gsgw6cGhu3Od7FGznwv7HTjJYig
nir+ty6HVwuBnC/N87MJiWM3jmrDIcYwGLHDMmwf/GHjUxQO5ne/gqTFl5Q4MtLWg0WHKLjOza2I
k1xup9moy0iK9YkdDSrISbR2+UIAdgGXIqD8GsZHw8kbUaSDFMLUIjSHPHFCOaxdjWxOHGmkDhtk
9mDKrY1hAga4Ezczw7wL/lTM3LTwV+BXkQ1RzKEDZCQuMzXH6lZC0xD6mYAe8dsfNgrAVebrpoGB
I4JmvKidaWTXsn6AJMC3VaVacQucoEH6YQJKOhvMqw9zSwlQ2keCR9aTgzSUFeljaJp/mEowum7R
KgvcQ2+m4bM/5jQIAvaoq28iFmf14t4cnVgeG/u4En0mHndpZ5Ihw7Tm02NwDslRJ9OJIfNql4t5
4thlFhVu6K0ge5npl/mpgCyJvFL1olVqyJJcJrtxsOV1BYsjNVRvh5wA9F7pUPRAmaV/AvhvRh3Q
x0qAp6fuamhEJDklSHw7fcaHd9LwXNWSHqx75CleoAPfy185AyJoemWnJ64fu/dl4ydwWcZzvz/C
CSRgKLsOaZrKE88lJ0wgaK0sn+7rWpYHmXyqv0fZ9kOlgUwmKX/SqgBAQHSN7YLe8SLlUTyjKfnu
Rxj9NxX0HmaElqUU0YTM9fLRF3cJICvq9RRqgyGZGclrUpbfrUFoKbK3vL1HuD6MCCsBOrzGUSEr
fkUyi7wc+ev2w+EBSYeqte0Lhgo5qMNFiVvJSSbU5/54aewmeJj6sZBIcWebxa3GsaVBptb4WPD1
7N0hlgzbmj/2qJB+ch5kOJ6y7x49v7XCJUcwlymmCjepg76Z7xIgOkgfi9QqcSUbJAO/+zPD2ihp
GdjkQZ+KCZ3nNpwrvIZCUtItftOZ1IZoAnmnP8NWoKexXrwkf5pjUtsTrdyjoc7aUoynbkix8oRr
zKbA+D4Fj9HQwmgtbk4QoP4pQYRzF0SA7+Mcz++hCFT6uFzc2B1Y4LQG9A1vlAA0zxgdSmgcKtqW
7P0xnTcbIr/PQxG53aFaS9S5QgLBOvoxlBTp+NrMwTLmqyBruT/UG+qiQausiNhvPeIwbx5HBvHZ
lN5DWUfAo5h0fGYrtsxcX1nm9GUZjNZhhmZj/q5Uaxkkrw8Xpc/hRhgJo4H93olK/jJuR2UjU1eC
zqMm+Cfvp6dz1lXyhp31tkE3qeaISblqPfZiEvLqS8Oh2edFPUkvjzcuunwjP0fbAlR9lmjgycey
9E8dlLSaTE5HR/wTyZlE7Qs1R9ifaBnd8vpBQvOidZIU/hH+0qJSBpfjYatj0ytnM2g2AZlg2vCt
YqUHq15WNukyfjvrwv6vU7ak+43WG8UbbhwcWkwefHCOyPfzu/CLboIkIeur/jhqMjC5Pzbhhkt6
KNylnIlcSubiMgDjeti//9aM1tDQeJQlO1P6R+0EhpGfPQZepM9E6gJeldyZdYsIAYm0+NHpt66B
AI8lzs9R/gw8EAuzzXNljV1bbVdoSbEz3fTSqC94yHwcz4QcmoGsC4otj+pZaQ8NbdtWHrHwqjBk
RkfNB516EA4EqivwtLVCjnrrPVAzbbImCzWLLrEUfIuZLn1rU70cGZrku/DJnXt+ULkrzm5QABPc
nhS3fJhp83WGMq6XD7pRuMvREQDY+JUNt2AeqaXxYBb3i492W8Aa+RlppFSXn6wESyxb7Gx4EKJD
TylEPPDMUUrLeUqh/95IFMSbE/OM9fdiBI293Hc5jrn9mhsFnNeLaYZCznLnovB5JNDILQ+cI7ix
Z/MEiOJN2uSiNW70aQtu5niZUONkUpvyK41MvfK6JcIDX53MGpSvkp8cUnlw48b3asoYohk4CAZ7
thwKr5iH0S4HtsS2svDKhuEeO59NJUHX3fJfkCpRx+d8E0NAqZPRlk59Oldnpdnm/yLtcIwZtta/
GtvNQRFZ4hQNe3IcyIcKVw7LRQr3hlg6klj+tsfSosRzVfpT1/7u8MzCO8RfwaduFdINGs2LHtYv
5BzSJwJh6mhSp+1P6DV+l8Pu5ejhFHH7A8RQygignWq9WpUd9sVmNRTcjvHozsTowx1ZZSdd+72N
EvHLcvAa3G7uOefsPmU2+R/CzU+37mGWpmOCVxwMQGKZfo23AKA8vP3W/d8bnySPdaqzjTXsvItH
3ASJIeUpGChcmEmLVRP8o9Hl/kF2NkeLxNYTzhSvT7RUhOofc1og4U9opECc08uB45yevnu7m6nG
/iD2ntSq2aTyaCobjjLSHS4Nu7SSaRR2e3JcJ/oiG3EEDa7KxPfQ45Qcsm/T5u7aBqOE5MqssREK
kXbdkpbVRy8CnjhHeD4rWjPG5vohEIpYESm3VFEBYdYhU4qzmi0y/u2wkZS9+Mo9r9B1U4LuubGu
1VAKBWfPXzxocAfkWMper6QqjFItZ8sEMLaPOjiE7gcG4rUX0QeCmEefcj56eq/M4aXoORuFVgZf
IHsmj3nmpHIE731lcYWc+hE4Nb4ZmEiFU87XlqF72+XMdes4LEzeF3T81F/Kh2Kfl/ZR7KXiAysZ
a1jqiLiHCTNouJY/ucLMUoERsgkBiLfBvKdkLgHAd2fJg8vQCctNXiEube3UJaut+YVykewSMSF9
QZg9xHW2B1yaXPy4D0vCpVC9V2Wt668myNtsZTFt2dCp1VTRG6aszbgwG4S7mNQ8odLmiDqjr4Lu
0aWjMZe+hw8N79nPmFJmrKDZWzCaWhjgnjk6xf9QBufOWj8mlJnEy72ynoaWvYjaoTEqoXZjdxUc
I0hQYcS+Ktx4oMm3Vl9ZC6OkQ0ylA9fGhyylHq7NZkVHjTaja4G/DGqB2/UH+tJMhSeMi+By8Ek4
aNHUhKzipZlfkmAKZ9PJiNKqIH8FNxnP9eyt/pRLYXFnIr6gDUmIa+klfej9Js4sPTzXdlmkfRgW
TJAqV6PDnaPjVH4EeUA5/w96cC1drn4v+fvpMDX3P1WIF/Qcepk1qlWhDhHAUgViyfceAzVVGCOm
mJNWkpGZW4ABrzXId4cUgC1aowBTT8sHf5O2OO9ShqfGGs4NlUO85C0/nOPlFYpX4t+Oc8ciKdoM
L/xAi8nOXR6FMgpTynlLq154d5r85JMs1VpZuObaP0/Vh/A5lop80UI3TJeN7tj4ApGHRxKylPYD
pSurpmGxKZYy8ZimNn3uoK/Inq7JITI/3JTkvZ320tgE55h1cCGzcnZJTgWgVCC0a2IzRk5otgY6
uX3hKKhNRK7BcfkfCR9gkmTxbUuJK8aEjRNIzjTXy+0VFj8Z0EUJ0nspTvQrrxn+hTOXXbAo9dhR
FkhTThUit+mSyKXEaqKJZQ9Ewamdm42L454wSUBUL6TErhJ5xnD3mkeUOZPVfVBcoikzoIPb4h5r
84ecpFj4hkalwy6nl/F9K/xgVdmd17SP0fyy+mYiRm4f6XTTcOzQjz1so88PfPtw+njQgkjYrhKX
LPaeZJb1tiIp+HJ99V85iEQO6O9qFXjmJitr7CLu7ipxqWERIkfiYCY++1jYEYVYsI8ImauIZjLu
MBzrqH1hyBa3+o2COZYOF98ZG2kUJzID15GUkD2wLgGNMEbtYCFSyBqA4UavYQ4WMfRViUM6CnhU
iCHCd67YN2jUMXZuehZliWqLMKRej8o99GCvRriDqzB27fbKgWZtaoxGv1QVA6MnXGfCPxFDhhnt
uBhN01uUtmyzxvXs7QGuLrwMDyD2sYkVRgr29Il3jmvz1y3jhQXMXdnLJ5jmvs/MetPohj0FbyhX
QNon5w0sifDO9jsTjKtA8ZlEO6qs4GygvoXd5Bbck0BdZ91eONRW8AZrbV8CE0BQX6gXajr0Db1/
9NNjRaMt6q3pVosJMiUAI+jfjXgxvVuQQeeTj8YXc1ppnVwijMSCiwZnPc/57p4gxF96JzdwrGu/
maMJ5n5JIPzqxpSi19wlcO91rsfSNJ08gecCGvZvxDj7fKSCspgn0VuVZBM9tEW6aEsGOvmXVsHW
/MCX22/+HmwFNqTHo+aQozVWNLmHV6pQPOPNOIZZ6TpaSeB2t9+UyaUkmDBOcTjQ2F/M9R5BIbL+
xg4NvlNemLrg/USDbWR3As60BdeYLmhDTcYiG4iZjkyQGyO56ey2RnzDqOdK3buJ2Hk5+qxlExoe
+brVM5pfd2RmzQtxY906JwTxx5ucpJf8FALabdrs2FW6RjWn4Vcjkoh5vFkp3XNKq7OydKVZdhhX
tu6HwtOz77DiKl3fQ3WzVY08o3WldrQWbvNjbGnnRrcbm43YXA/IhSSvoj7Zdj+M8FkqUo0qyml6
idNEwOoNBiK/hLePjIP1WCQ7D1AZCftpucKD/XyD+xHxY+6yeJMOeF+fyiVmHGj/YNZPvyMgRr/c
sXWjF1MGnU6P2VYveZuHwTf78XO+7BNKzsAHuILc8VZX1TPfavBCk0oBay0uqf3CeQMoIEBVdVJC
9fGoIcxft6gKkWu83zaaZpe6vAoNFEM4g1KOVjrnJ/SuDsm+t2E8Uso0AHjPtKxJYANMCMiA8ewi
yNYtjWwpGcslqBfELDQ6Js4F+eyFBkNbabVJz0Je0eq0R3g8jm0QI4R4oAFDzoo0UoPPsBr0MbNu
PZhO8yg4cemG1F4uC6s0y2freM90omFWRurNU+cPOXV+HSGpLXH3P/JeJejX1xaCoch8rr4tgTFY
TH39aPMJi8cheYOUzmlBGHdUz8ZYj51mnv9+tGSK3nfM6HxMHPK+crL9eENb03ceXKcn4AxMxgpJ
5L96OFybOOBHzXATJWOxHwklkYQXfowI9UJdOZ60Fq/S21hgnmGccAs7B81IPamfJYmSBn+mXqK6
p8hFsXFlx86Lq95qL5EykWJxi6wK+IGV6Ke8fEXZQ0EKU8yHL53FjK5jX+IHyoKM1CCE7Y46fzzb
vhOqTaPGmB0M2tcqmvXj2RwHwa/3pdMODhmC4H/UF+crACtbV8EYk+CtoG63XeEagqa3TKurvbew
6IvGBypXBxFhOBBRipJU7LKZ1ZoYQpQ+wJGKUc3xKFnGosxOphgMhpwl0ekpGHYNlzWe29qp8NCE
vc3UQTmQZTSBTTCmmstsnpBgWKhHG5ItUS680imLL5TCP09mMkKIROCtYEACyPfxCsEl92zmQuOA
TfTYKuT49qHaytqrf2lFqODmg01Hr43/bJ2mD/eTPo1OD6c3u0kIxbGxxkLetcX2jmU3kfcMjz+H
5J5H7bKMEVu9nfsBWbpJgGARF8PxVYxlJG2e6ORBQRyh39t0pcU+3avmjvHRrrLG1LRH5Y+I4E58
egaZg1VztYod88vS4Ho2xdd8EQ76xyPmOTCA/BI5xrQ7c6ebJkSh1jNELcPwGa780YFwe7XTdliD
N6LZIQRI6MT+d5fTO6bWkdOn+LAhD3OUbf06HOQj0E8/3IHDY/+L8esA2kXz2YNqi8lryS58G+8Z
hPijtJlWCKz/km5IfHhx8S4yLkFHaBjroqZ1OOmWhJcTztLUkmQ0nXeB9kLnTqFyXywnpKpRBTlH
nvph96YjXjHt3JaLZyc/yzdpTd5gkGAHXc3H5bi9bWYc4NMzNKAVG7lZLX4xrj7rb3bC6MAiO9OH
oyrvFpfRsonvOLe/3vXiye1c9zVaXyRlY2HtdOU00BjN2WsamQCLEBrgYoGSEIieT2rAs9aufy4Z
X0H69+VMcyGf2vnQ1tgVC57L8T2WMzjWU+l14QQxMXBRUF0Kv6G5TsblGcI1uXiEaYE+ju2YEngs
PoH9Jd1zQyrPNkvdC3HDrxmkcPd5rk/gqEaXzjfaokH/0GS3klsCcM+65auBA58yfC3wOcK9XrHp
CAjs8//l5eUUzUW31d11jqXL72XpPdgJNvdmdomNzRfM20+ARItVB0lXx507E3j7CF35LNpCMzZZ
jZbsnC5QJ1syDzE7bQmrPiPQ9uIt/CgXlhgsikvZVbIGMwPtcEAMEBGPxW5FGje6Z419jndjXr3X
b3HcZT389Iyg49H2dBgiGN0x9BHc4yYba3a8cOrGxkKnTRNqv/SNRUTJL8jU9SfvFxQ+wr8mEEcT
7nFzTjI2zvidcD7API8/w6WobojExfF7XufnwmzXlZlk6KixEJCeyYX/SRgYbbec4s8oFt+0fHbX
LvDjWUH1MNS21+xCk7XQmt5EH0EgqMW63RCUtlRdOUkz8L4DeZIML/nrWdNVcJfTAqvLXYVmciVR
49BM44q7SuCGxhyG7Lb7etuF7vQ1m216gHxvkqlLAlvVHLjbIc/9O5aZiQGvb5BUe8oAXUe0m+ME
a6wZvow89A3EyfQw4YfSYM//xIca5uLDxo+/QO25i7GxInIKyVlI8w1elcpIxdgcC4uZdipSqZX1
9OscR4bhsPh7eYpfeuGdFdEtk/2k5wBUvuoeRh7nirvctolj034u0+cPzdzfC5ef8q6ytzKqs+1j
TkKx1dJXs0saus/llSb70cty+n1HsKAoOSLrdNKL0bbtTnmV6kDNc/yj4ob1Cj20U4ingGDFk/Pe
WK9G37vVPYHcMrZLbC4Dsg2pfQ9zy4EyEuDQTUGlEGOhogtkCAHHm3jT/3CqiqidDP5PWN7gYAOa
hZaTpKnohvjA3Z4f5eydTKjwIBtNr8YYXW0hf06hOvh7EvzhgyUYIz/RW5XVAncFOmu4oYtTKMyh
C2fhTimnT4nn8il1eqyJjTuQibKZcl9goIalzR5PXLrkEVqfLC6ZprO/8SDObrJqFez8GfXALxjS
q9TAyRmKavHEZi+S6+HysqjQucQwAk5KKesyiTYGRt7AG8h+js4UOqdiJkXDghiN/Cc4utlneMXC
NWAJO09bZLUW62UnnUa4HcjDKfuD+MJmJMq1OJmvkHH9GNA6Uk8IZlAoyNikVqhaAGpgm3chn23/
A7h9TBTV8WR2NNbuxoARRj357edgdzCjH2rmziUuK6feA5Fc9bT/R1wQ7S3OTtn05Xu6XGB3NH8G
Ax9ZIwdctkYL6ieu//GgLIHX5woGjYFCYg0QTjaVE4GWZ8G/HJQOB+tytt3u2cJYXwigi1/cpXd2
p1ZDCUT3BZgHszcrP5z3tkdTJVDph7d5r2aQMnUItIFlQdCrQBdjaG4ZsUmZR5ILbkAckxieUNk/
7ioyYTo5QAth3tNEj0J020Jw+SmIe3y5uGe/1vYCBeo0yXNlE6g3nLubhjROEja8Bq7O2Yrfm5wV
5a1xKZBMCU0aafFMWKIDwMSnd0qI5+z97n9s8V0hHJjvW14PkQJR77OpDHE1snKN95AnD2pDZipI
hSTKEaJeUF1IvEdI2/mZwZnDu9MqZ9WPWCJ6sjo9f6QHUnYNEl0wvzHSE3GgZVqo6VT0E0oFUSRz
DiNGLK/T1pXhePoDGwsVUNf3W3z9N9pXWfIUhn8L8B176YMcMoZHl+PbXOBNw5RQAkGSxQEkJSQ7
l3NFdm/ZKdgP6LgHmkqZr4szulhW/aK18DaBGxXh+4xU4/FV8h3mIlwmcQEPkNxqDgaieq6MTS+4
VyYxKIDOYIds/SbCG62BKWgzdV2immfykocx8i+4CLXR6B+VcPQD7OWuT+1/ZmWTnLkzEwZKVfLA
05KbOY4FqE92yFXVUXgfj4fqRUIediIMIdSVbRkWZPNRTqN8oUUUy+5rxrvw3h6EyyjZvVEf/Q8w
T0yPd0u/kEHfgjNtrIMIalrDBKAbhX+rAKDtsZz6yqBmvMT939vA/Mojqq6xffV+QBL3Bvzstfik
f3PRDqP3eTXCUbApdRtccNhzWj/GAOIL4pA0h+Y+uiIC5cM7NeMyaytvp3SRr86N3sFL4PCYzPzS
Q4QDIak889XllrpyeUX1d5k7zeaMufiJAiFVZWdV7mYJtTsf/ht9TJcQBc+0/rZ6VDACBORcRVRo
scm1a+ZwWbAJYTHTNjnBGhTXg7XgLaglLV5m2t+xj8JD4/7elJJmw6hAB3y4LwZklMn6G2AM20LU
t+grCSGl1CLjnQ1cqA8BRAgv4YfiHUHSPbmvUi/qKDvwcC5yNYPDo4YINfeeJ83hWmOaHmbORLUb
+CSY2c8Rrq31NKaGpWGU85i6lrmMDtRKczkJtCXP9vtAUHx+fv3nMYc2qdL/L73NzZqie75m4VKL
nglE4iwzSbd3foyM6CZG7ipCB6UVkJu1iglzabg7LOGEZVSSLeqFtS0Fos7cAoxmtAvS+jBvE/PP
BH36N1yOLx1usx9O2QlwPrf+29yIAzYCEWApWf9HZyw6DrNJpUnt+yr5gskm6uAqw2dbL/JzaP4F
8oC0IE2al9cEOeBoXj8T45PHrj/9xpvAwGV2bmD0c2n9Uxd7oI5rKQnfij675i13yq10qiD+h5y0
9hC1KKU1ZJjdbhGBpPU6wONDkojbn9JSu99C3aUU/5+jpOCzTkVmBh7LL1xoYcn9kiDSNVvbUYE4
Idew4HYqUUouJGtmbpwERPnNELrjEO4vm3o5t8CdBDIm8xqqg93DQGSYERQX3FmnlNKh2Os5xEwg
s2whPw7mgmifOhqt15uhYkbVwOYIxzxgJpKZcNLrV611v5c/1NefinOHG3RPFM/qrJDm0ainlqYL
GKiW+WUCxVE26XLBvykzoW0lM3zQIBeocw3TNcH3ie9a0/ffStyYcwJwk9G+DDv7vIPGxjL6KbC9
0GomMnFPYT6iw0pzfZaDEzxeApM8xrFQB/s32Q1ZY6wgciPpoIx27r6zKfoNh3FJ/rqYF3De1kNT
y9Sfeh/uFUDu9fdM5PUoZPawhvXBgFi4G0NEaPtM5Qw6GcHFLAkh2p2ObjVNeycCpXmr08CYbGPp
khv/kJq/htpy0Z+e8crfUG9O8lIGjC9PjiCkisWGFhegfQ4snp6/MZiY6cqwMXz8tcN+lrBnFEkw
y58/y4VhcrjUU9AfwykMud4CKrqSN9cQGixnhBoKmjARANWNxw7Pp6nEm9SvlwEBQoMRp+LahEXE
rz5CzsEVBEmq6oMq2daQO4HDafSpkolOrHa8jiZBgV61F5q8x4dz8nzusNjcXUN0W02mrgF1/AzH
d09wuWQZRKILF0Jnp8I0zlO2XlIe13rZlysXRaLFsRxzm8GVV3cMcq8LJbAKKdvBwa19yTA+nHPO
CJNSNWXR/hfKeytbYTEmkHqIawPWgbsJkjIzBdjPrN4q4cvU+DYtgAImvU796oV/D9N2sPJhYB0E
2oqSzp2kcdnPs8dit9y59IhCy5b1rIh59kR1M3lgwmIN8MmrFlg+f7c2DSJnBpqJNXVjxnaXjkvl
cQZ0vbZW4qZEJoaF7AnCocTywm2Y66HHOTv5Kftv90NYMPVnB8aQBCP3Xz1BMa9aIXQObTkMmhkJ
k1tbR1+4iguiTeDdprekSVV3zqCn6cP6Ajnm9Jwx225qgoyg5dn6plrw4NK42Rw6xcrO7E1osf6D
cn2LjH7gRYoshdu51Tns2cvdjv2NX96zX2oGgE4RyXXs8SmjCQhJZGwruIXH5IfZy6Vo4qErT8xj
JO+K3ekvf1gs3UySzW4++SxXZQax/jC14OKaCJVtbF65XYAWWLmhiHSvUsh7uXr059H4aiD1XDvX
axxaqUNmJSnrA++9dJ6l38Ryr0kXg4M6TVGK+wJTGE9HD21X43FkOpTpRKBONxLCJR9aWgypEUQC
F/u+FLeAQ+wrbIvyRXxH2v9TAD3Gy/gb/dLxcAqHYwgvs71gyU5K9JOzDdJXgPBvl7HYSSXBpJJC
8lyGWueV1Uvau7UlYSmYHCXgRI/P55rx+C7ZPoIpDBswzCOiwcSrZztu6+cA3zca6wnNJ1HqPjXl
C/ye3zFW681Q0ATakUss01EZ5FpnbVf/AoTnNQqerPC2zVsxx7MOdEDKMaaXvrQdt9/gzBlrFZ1d
9zPVadwoQ2HGcA64y1qjCxN93OQ+TXTU283TSti7lyeXGJj2DmDFD00ymIORt86TIu0UZFDF8phB
HH/ww2V4HsYYv41cRIYbw1s+b/5lWu44mmLqDK4OtLYE1K26EljEJPsxqovXwheHQqex+Ii/Z6V4
oxM+FhfWPZnG+6dT2IRDHMdYo1LOhPcQRST9xb8wypleXZYzEAPKbgO9uQWz3DroFLXyk/mNgMqR
R663rXlHu84un0QPwQ8hwflxzxDCghR9d8NZP0kjy1xFGs24zjm8aIHWFGtwv4DUmLagWp1n9IIu
BSbqZc8Y2zvnnJtr9A/IVhv/6OEbTYkviJaODDS7w9eGxJWeJGbhYd77sm1XjFvwRK0lfrxOiiL1
n4i5oG97tQRHehDWcdrEyyAHr3Ao5e5TSVfjhzJ/3VAXSmMJ+JitTw0/SciZYad9MFBlX6jJ6US1
a9nEmE9+K47Twi8NnI4Uxgs0M4doWCRgOKhg4N6+Q6zsTKhETk40lzqTEY0F/zuq9Q2Ws0OiDpgG
yuVxBS+mTovZsnVimnm61yKmcXqRPe/XMN2Td5RW8VqfOJx36Wm8D7GilIero4BPHngz6qfhs/qx
mjRC12q1/zrardJ/jMBY0n7VPMS+M23P/+3YHSqDN5mdVVLlzMpDAp0Tb+87qTGIf2cKbCaSxVfI
QjMiD1lkMEMnwLDjyBcv72IfEeNwxiFRHiN4LHGmivGBMvxvwOpOyap32b0kEofaWDh5KBxpY2NQ
w0+Z6IoM3DCw3P+5jbjt0fJ5JcYjOF3/2pnsPjYLbibaRsCflL4u7kVsqLBZPqI+BrNcyCooBP88
2asRn+KL8fg0wub09TGhka7hA9uZI9RlNkIsWCnvUNqiX3w1u+1Iz4k1ntIM2jImXV+OXOJVsYQZ
d/vVMIBACYCb6ftnz31wd26Q0tRpwPiEuCg6QtGz3lCfl5aBvlmHAGBwxVWtv6OZFkVJWSrROzV2
JFHUESBSrJfVuWE+1bpBAY+IDj/T1jvjTHF8nQSg1PCp4oIx8nGzZPEwccq4pKOAI759FaqHl09e
HSenodkHv/pbPalUTFluVyr30Ec5UPO6TAjmwFz9SIjv7EY1TNhwaXpEruU+wOsTUJRQPZF6YRgg
f/Tr7g0nEkAFloGYwdBeIE3n7ny0xcj+4t17wNE83aqPOkxGpW9eWZ9XkmCTVoXO2F7/ynb+eBLg
LfWMRdMvqanan2xkVg7JPt8J9NhZ8b8l2ulWNPJ5whxr5NZB2J/jGKqBhxwx1euwo5IlnqvRPD0+
rC8VqYDBANEjPl91Rz0k3T5lRx9D7VsKWESpXYKjC2ChFdbbeVnR09bJD1E3BidlNo4t2LeDGGVn
yJXDBcZTjG+zAs6pT6Xf2zyshSfhSXjNxJTx40qZ2Uz65PLTv1qFbLrMv4N+/wwVckyTJ7KWg5gN
AZ1jdzO4EKSX8BHJChQWSfIEiNOXOnT5UQ9JwjKRQ9BfhwNR6Luu7XjaXNMTOz5nwlNgU/RcVbgd
HQUFgu5WL5sSuyfRwiWK7YH4WjnTQZ/Cu0VFYO4s15vYQIBjXmsJL3cDHy96JdttdU8eVa5F6IqD
iqeLU8MwS5DUVBeOM/86p8sL1PGbnf9vL+MliDluwOUZ2GSEsrDHYAacr4iZEisoaOwp+Jjk2oWz
ioUhzBW9tcj6Ohp1A5VrxMfntKYbjaHNl2Xu+hapPe4XTipkdkgcAlFgjHLUkBz5XssGLkFVDKXh
lFwDL6HaoivSTOjzPxmkZUqkwVXMUToKiGRLphaHNcPoOHPt8xwS0wjC+PCFwoPRyp84vzJhl7Rz
X00+EL3leKBlcaRjpbuS7JrsNygsGsOIqvWr6cqu9YYC9CbuoaRwteOdyM14f8ykq5np8A0XaXbD
YShmZ6kGa79qqzaepMnIjAuHhB+gv3Dnh1LtUv5eS4LUJ2ON4Y3NPopZaxXTMznqYHAfnfpwHCmF
fRRPSmazUSAB3LPXfDDOppilh9MJKT95k/2ABsg2EoI/7RZjVK0t4m7jDPPKVPUcs387afvRALY1
9J0ouQHjvjyaa6EcdzGSxkya4jcZekxbcNH2etkBrKXBNqmuMvGURTVcsRs3eu6XB8Y0sTAyTDmp
ZPj8XtB0FIrls6maQKhP2K43Mvpb4jhVHBHy8NjKjE8vgdfk5NP5X7EVCpqauQICF/8IhlptEaMO
odY1uviEQlfWiwuZcblq2t/BsIPS8PoELY9svfiLfxto0/ggiTkpjoOxyVuiprVtrQLUskCkaHR1
aH0WZafb8TmuveuMBhCjHXCPS/hs5aq3hBcwKjVbA3dkxlxExrKFwEkvA0+UoRGcS+6NB49CRy3p
lo4DGG8KKZMflfkuoGB9+S21F11wo9mSMzDaFwdP7X94v58aL1radfl6RySqU5rpjf2VoxNxUUja
ziuzs6ILTMZlpu1CZOrblxUzVzPHVMpuDuj6WGT++2uEul1mfdPMefZA3Kb9UwShNTbDxPL5PaTY
fXXol/f9hFM0EiRAZ2XDgUTVoaAkPq0A8QvCRTQxjB0Ax4ZmNIc0ePJXfxCCvV6aj5MAeoabuEFh
9XP/ZLHBh6Nx85Puw0mNrpm1gZFvMvczYIgzBFvKmNcJ1I03RUzh6QaiXFpw+MPm9ghV1Cd6YTf5
ZBaFs4qPd17jOjCv9wI8fZwVhun//tDJLybK9jgRC0t6bhGF+nr6UF18nS0tteKTxYM52Q5WQn72
OAslYkMUYfVj/9j3Y3dFZIc1T0OVHTwFdJmrVxYyrDIVr12t5uQTZxQ2P7IWc5WyUeW7eWiUAyLM
LkkdqiFU9P3SRSOXtc6C6GrJ0nE+rvo1C3YatVw0uZ4uZ6XZnnwtVBet13q93tfq0//BAxxR+3cc
IbtTCJJWVWOX7o8CehmjrHApD0D7d5mMssVBSnx5dQAgEc1UFUBIkYDM9BbqCxeIf0DMYH5d2Fl2
o7JckfebxZK2kwZn22HLcKWIeR2ijmz/AW3Jn+4cJwQs7v50dTQpgETPDfHwmtjkmWnOFuv/HxAa
eb6Mo+hTlH5PC2OJ8XM5RaClrEvYeIdWmKoLr9yg0IxE3uRYAI2Yxbp0cxpmGOlNXukEY1AaikV8
qAdWh4GwDiqpKVuPZRCWuuesZuTfSfWRKaEwkorkHsBOl8ZYdWuKDYRoGLB7n7mCXX/+mNwLcX9S
i+n33eUGm555OS0lYyLgVx3OTKnfx1MLikZNEipdBcg872BWs0KKX45Xd2GCIzYLBHqk5/Wo3LLs
NFCWEpvXEMdJngs299qAFeUgL1bqPRQP+1EZU6hxbRGlrHYqZ2lrQBJ2hrCiWfF//Gtjy9Hh0WWq
Y+zreSapltZXZEpU7dnDXzUN0ek1XOPjz9uNNE5G1y4dnM9l6fAxc309GKcfqmDGOLbZAaX47Oin
pSJnBglmSIdsj69PNDYxtXOKM0dMfoyAE2XvnmIkSNVRjzXTtUWBc1geTfDQzW+bqM9BhxDM90XI
ez4O3DX5DHUSt8bZ4RXxNi+DSEv7uPsHf9x3W4d1aX7YVbRiD21mXYnYj2rIlk9wNLCL8A31VdrP
UdwMMUpKcNSx7Va454Y9QOgqa8+c0ntCk/0+qNfajztOgrpaTPW5q3XwDTSJkl3F4QfVb9If587q
WsKrTIvpArsDD1IOowxUJAHr1TGVBXsN9N9dTkVu+5nA+X/pRGLteiZjc1TgLc+lAB9Pyg/FjrXr
CTnlevxewUECwQnEQCdr6eJG39LmDggCxx3Qms0euTvJ3Y7bXuECEuFCzmnq5+XFz+A6vFOL91Oq
Wueggxufr2EqpRN6gvchneubGTJ6JQPtgXEoi9Kc7B9bj9dQ+T6E7cVsfwJnIlAjBjo7YQNXnsZ9
XAPn0yl7VFJDwoXzUiJ4aJem69+wft7v+T4njCidA7Rv6ASLG3d/xsZKfzq0qQ3pD3MTfCMxWQ9z
ncs45XmNdsmgFIKBY0H8bzUHT8vJ58DppZFN0zzGNvhuChoNqLbucD1zzWY7rX9MzPhfy0r9yG22
S81qIM6ks11PPgRg7Aopc2dBSEgRXMAvbHAWmQwhkktWf85JaLQdUckhJFwYtacWakyEFqufNyTf
8h/ASJf4TfHb+/GB+XiD1W8zTyi9UxOIaSWn2/npnjIXcE0iMDHrvA9gHFnmXXwbLeVJkkkhRTui
W3kA0pWqcTgTzFQa48qIIvg5XlDoLh7GmWgefrwg9K/klBbkA+uzotY6O+w640r2boWxxrtf3d7Y
NggHtXc2p8VNM4FYrKkaGxpTzrdPcUbggiHPTD6/P6eBLzmkVCZ9610rk3GvqnPTXJ5fZ4tNhs7c
Ny8Oc7oDZhDq3BkoM94Hi8bBUN3+4NFEwInV52r3H0Cb7zL3oWz9o7Il1BL0XXqenJ4Mb8aLYYAR
2/f2XHFmuK3DnbOQescBsRV5yJTaHQV7w4HsfwBGKyjO84hPwScXoS/k9yzj5lN45TCEXedCd7jm
9r7SsJhGjgTng1PA7gMkT1FT8raj//NxYB5Af1vQGzhYpXUT5OY3ldOa/wFWR6DjB6VfVjKiJAOz
c5DNjQ4QyM1PjEWwnb8dXdryaSBqGup7HBcfMnyqPEji4rpXeLCIXDMsUDWClEtU8Go3D3/y0jfK
24OW/npUq2trSDe4LNAi9bhMKNGhBrvyQQ5YC7bqJMg2YH4f/1O+wuhNOpI+k7qks/k82jQ5kVhV
Rt3OAuJX2Yv+2Wr1gw9OCCIEvXI/04V4c2bQ+qnu2i/46hrZizPtPM7GqehHOuctKttZ2xlSTzNk
VT0I6VZOSHj6aPTe4AOiDUbh8W8J6uuPbCXPo8jo2/43yaqPegOnCgTsPPUYYnI9ziH49R00sSko
RW5uB0j4uMyzf4bctEoYVNcjCUe7s7WpjLZKOWwNRyq9K9UPUxrGkFlvzWLn01SSES74b0zTxaF7
yq0HfDNMrRCVz6WpMM7b/TBQXlPU06EBoLGe8dnDqnbJ2qQsUIfDMXwC9yCre0LfVeMvMrABSHuv
yoDeq5ECjKxTfp7PbuqKvi0SOAPAXwxarfTre8opGQ8xY1McXUBCTNVeJZHxvAFOVD3uzyk7kAuh
YsQ2ra7JHkl5ZPYTWzgXyoCuj1uXmjvehpNCcr1Lf+VUjzA7MUWc9rT/0O/+Pc4qv60iK1nYjaTT
BY8x7+TNvtXIpditz7gWkAV9NQM2HQmP2vhCTw8BTmrD4LJkGzAYq86s+n6OkBsJRfKVUrdxZ0gV
OUWwcLU90rv7t2Vxo70xdgKY72BMZrq8nJnbtBna3PjQ7jhBvpTdaJ7jWvy2JWBQmFkQOUWECz/E
rQyygEE5CVQduk3WI50GPnOzChdeZyH8xqzQKnEtyhomgqyie/GNxH+93lv1lzP7W2jnA9ZLnhtt
jYhYmLQQzHKS2r5TYJXLWFD/hIE3fqeVwltJgkHQi0gGToH1/Jb7OcVg6cCkVLULBzszoNR1BjBX
FPjU/L8k/w99lL111zq82hZomNAhZtq4zBgHiUqLX8h7AaV53Zb4SkJBnB4MgUCf1xyphf0wh6rl
IAi3khbR9wwd2J+acBBN2w0/vpytFY3VHAfcYU5M7vm+pQt1+iU+Gd2SRHbfs13tg9O05slGAMMQ
RM74A4whEfMuRKQSbz0+hUuzt3ao3qBQFDRgaj3DM0RAleY8rA0wVrFuumfadOd42+ugi33XnLmQ
MdVTdZi3r6RwtmnD+gyCbyTeXTHqxCFnBge/PRA6bNS7kjWaPBC45Zx3zQ+MjAGMchSbsRQThLcY
JpFXNzd/i6LrtJ8jBD8Zq+BP3UeKfaapEhzUR0J88RbJFZZul89E45ObZ6bbAEEWVKQoaAOiqE4s
8q+hLIcC76qKUdq88OFn0jC4is+osIpA0WTZSm9kb4r+a7qHPuieupv4Ld0dhlnNiNMS5MfVqr+V
y3VN4i2MuZNtj9ahYmSdVC8srn0TlksKtIf4qTKE2daZ2s4FqWznTHGLE+gWydcVZplvOa1xO/m7
TJfZIHedSC0Brz/M4SlPY/S2Ea+2k2smXNVwO06div2rcHg4Rjq4oRPI9h79kzGsI8vdSvDT+luv
g4JHktxaZNgpe9EUsamabmAeTC+14uXY117TsJRFSnaVdbolZUaeoVf7Ykd98SwFXjN036clfN7S
YS6eliUBdn88UU7OrILFm9VJ4i8G7713ILcSAY6ehZwvR2dwZMNUBqq59e+8jo6TDT7KUmNmJi+T
d3hUF1gBfNM6N+KH4/gFXFWJeZdUxL81CkV96CQCQ9DnJIpFjOciXlx+I6Gxezyssj3okaJE8+HH
XeuwvsDIH49LAabqajiBY2XH9B8A7u/69N/yCmvzJhLRKdxBWrqB0H411RzG1ZGQaSfX9zzyN/Cy
0LHCwwB/FjuDs5gErdLOUJGXsqxa6jDVqxqmthwg9p5E7uc5z+Bltv7GNjADzpBUSoI64i2B55v7
3JMdyvkAddZDpkcc2phghaHDQrZkXpOrYN9s0YDVwinZynmev6GJ2R0emgnZGf47m4Tczee8r4IW
Hevn93Cp48Z3OsdfPgkggtouMrWQ6LkgJnOpn367zsl7b8JH7l+XTz2jsou7vynAtZfxGHmNsLmk
EZG1kTfvGVGVFleEWCvYqvOckX0T4h0KM6HU8kfKcYXyXVvjVHs9tfEAl9eHCZCfVqk13Zi4psol
k96Uoh+yNAkia8R5eQ6vHuus9dcamkhLPYsUbnqwy91j4yy+GaWOS2pTNW+hgx31Kmk98jvSsztg
RcBHVf97lNw9Vt2BS1E+XFgM004NLQGuuDebJUr+UqnUxSRMBoBZwD9KQ2sZCRqgXehIow156r+T
YjTKTvvScjr+v7ebjIvOQP+9B71a+xXOWNCD0YPfkZ/AD78Lxy/nXWWNbXbLjBEZ1PjQ6un7AKhB
dlb/jk3cZOVVH2v/4qj2cbQBOzypoXAg6Lrk1tGWSUqbkBpE7Rsqx33PsbHa7IGTL9ALkUQAsuun
eDBdQpxMKxbSvPslB8SZGcpxcsRXEazuIe7lWnGVB8w2VxIuJatucJIVLW8K+xGPR87YlcQb/e3/
GjX+cAG77vOByBlSTb8BTaAPPasEMDHJAb/TYhxiMKvzLFPExhFN/DcyCqcVazefPfBzOb7mUpOk
+URfWVwsPXmJxrOCngJ0zgGXc8ydRlNKllGC1M+C5WZhXBNs9MwVpCO8KB9a3VpnJ1hORWMXJzBv
t1YLPh66BPO6d90C+uAdw9XjnulxdXn7Cd2TZQOJqLVeWMmd96MrXm5xTx6wDV9m+RZs508FcQfV
lm3T6lnFfqGqFNVYMIHcDo+OP2/RNuUV5Nu2ZBGmGS2WFc+JAB0M5F338SXuHPUkc3ThM5TKYtr9
ox5FqXIV5aCOnoGHF8Qj66JAahGSDEpCEqS9B7YLezOHXyv2L41F6og5fjwOEg9le+v253FSCyYW
IR+QGwfxig+twbtEoiUE/v+2CzjMzTpj8LFl5By95uilGH8U+7/j8iCJzw62mv/cSrhiq7x3M82f
qUbKeF08W2hDd9nbt7HCOTn4egjmmGuaYYYcDQnVzuvDS69czzWl0uyDAfZdSodoU7GrZ1oTNKGz
OApXbouq/1GGDPCDBacVhZXovYMrjzP8BxvG3pR9lMrowehkNN3F8Fb519pVmCliPW0D+L5nkvy5
kxEFaLAQFCcwg9sXOBBlSDmP7ezedVWP45f9I0okbpAtZlNvfFWjQBeOQ8f9nyOZLO9OOcBNko92
sprxcNFrPDxSIM5THX0wQiO3PM7aWadYj9LW7y24a4zEPr6NIjXV8dX9TRfRxfXDmd3lvPV2ViuH
lkpJ9KqCX6rTyBvZXXg4PJ0VoCbd4R+USzw0ZJif3lg+qeOzXaNIvQj/qxj0LLID27uoRmQrLRoa
A+Zkbdys7M0EXJ+y9OfWkKP8OVO1JPwwXUfwt6Yk6MAudViS0b2Ac1OITgnJggqP0qlbT6qV4Ope
KBJPL97JrGX6hBJiaWrKullG+qQhPiULZxMNGa27rF5qf1fXdf8gF5/Ort6eRCe+t8i5erxJsxKL
+nrZSZ3UpHiJ5QaflkfuFTHbCsfdRQ3K9pQql+qqZl/tTOjnRyq4ZF/ZkClNFMVCutdOZa26KcU5
ktpujEzygJptA73V6YdMA5Pf9veIaq+qA7xCh+cYb5vyZx5UEO2JayThoSrGyMwYtOVoGsTmuSoX
nIvwDy8U6TwjMT4wvxjQARFmkcdKQlqNrBvSkJK3AGuZRqeFoDpwFjm849+nGyHWGE5KOYY218Tq
8tMgW2iwLmESBWsREbjVcFqtp77z0TIAeW4jQZsTvkWdGU0slR1rf8DTROIBwam72J/Kutr+3i+p
tmfc074V5f0Sev4Y+aDCpQJdoUrkK3Ema1HEN8E6vp5Klp/i2sxVywJZqbbFcA3p1bb1DH1/+38J
6UNKHNHLOwp0+aNgXJSJIGM7b6Zrra4+cuAVz18Y178Drm+9DFaS35amkHUI6wdPurZHvsIIfq2S
WSZPxGUOP0xciVBfJmlEE+RqhDvSQCM5uWDcZrnxEo6hkwPcRBgta4A/Xw93ou/5XKP6EX+IOFFP
kAsIScc2K+P9DLCstDJvBTVlcnFTxyhX2IEsCu0PYotWJRva4FGCgk/d8y9CjmoMH6yzPHonlzs9
n5/6jUVDMvEYUprqDpqeZOIl+FOqUw7bQfvve5X5r7eQ8diYPlZCcLil05Bo4y+YUNDXyXAeNP9Y
kD4QA0nsd4lxNqdH5jtsF39edu6U3F8p7PZPz4no1j52iq9eN/1AwszHzl2RovFKnrHMaIv7C0oD
u3f35gabqk2uw9xdFAEkR46y2o4VBLn6aeAiEy0Yo5wWpmdme+gPLufCRVEO0EpYUjdrxLuVASHa
uNk6UKAN6lXLH291k6qZ8fMy0QnTU2qVROF6NLnE2sDI/pukGN4lXpUl1MJn0mYimJ0Bp6HBdrBu
9SaFCxsT4yC8y+rLRCVPvK0YvI8ZKsORmXl+cTcoSV3hImmuv+gGsjkTN/r71lHh9XDV/HNHERwr
aJtePTedTL9FvikjkmZmvbxaxJaYZlJN4UQOiUh+I6tsCpO8TNWsRVLcnD7VMQkOGcMGQIKrwCIh
H4swXwKYUv1sn+TWcSKH2LuerUIRZtyGrib8SUCs4kggLwpd0zjbQydMx1AhlHDhWfpeP1txsw6+
qFOKOIhKNC3FeL1LUeHRy+wZZAR4v3DJybaL+vP56c2ZMRNfOiALALZT4p+16fH34Tf6+Y71oyPG
Lpzxaf6YNBGm9VmBPmNnTCeVNdSkscIRsGMWwgnfpXl2X/6c+MRp0X8hEOatcllU9u3naCOUDezY
JiK2oM7AWb3uIoJpFylcSZWDOSlJWXlu0h/MKnKqSQrEzx2KR3cG9egbWrg+nywbvAhwnZ8jT0hx
2BQ0CL3qwHivnMKnzedTt02ZFJ+uV7XZpn9zkYND8Y3g6P/avkIQWWLKq5SP4PvEDli9xMPwDXbG
PHoXgwc6qbUWi+EkYvRAeJCK2GsnhPUYTbS1vD5v2KW+5ow1JYr7mrO+yKAWxXxLRDw0rxIXd0eD
h5W1Fd/URl2/xPjl1RWSJPpOk4sVIWSmY9ZMFphbu4Gi9FmDqOOBKO41HQlUXkxtN94+MZZK6Sch
+j+R6JmjeTsUCHHbghvGtXumWyfq9qFjsmLnbg/9fgU7Qc+5ERUOB5i9yIpVshfqonGqgJ3UQbJR
nt1uuzx+HSQ5gzG4D4he7Wy1D8NqandaYJRpBaHrC9fhb09lGuVqhfa+9NW5hGN7j6zTBAs6bgLL
FdAgBaGCclh3/qh2JSbwZkhbxRezPASyWCY6Iyf1WNHAZhicuqdgjVoaWL1/ZyU7glXq8NCDvMFw
oDxTUdcLTfs9NiON+3FX9lwc8hCxsinY16LjSt59z/AG4VrpPbGrzu3HG3E+BkrHYLxkEaYSJJS1
+Wji1OsI4zIsfWi+hy93ECJukWZ4Uams6we7uFMNeQRNh7npQ85LBOAGpM5NTofZdIWpwSTjgL1n
v6ipz6HF/H88giV1V59XNhNEdtVbMICcdyywYYJguJ559+fm6EtZe6dQBdXjaIQYIBBesrkv6WKd
2s3mdVgOCqGbaBzUg+rKwjbi/xfaHC8kB/HQHkvKkPbbqBx+kcBuAA7RQjEh3FVG1WR7KsWMRnf9
mBKo8J1vgIvCycMGkQos9r4TTSh/xpnenmGz6SlXwPA1BdQYlu6qsPH8Aq/h3ESfTo3ahDjkuD2I
uwZ3lj1ovUtMjacPumEpPCzHbz+Fjylxz6LdJjRsVjcoVW4Iw61OY69Zd4X2BPcLxPJEZdx6RBAA
9TOvHTtqo1jOngzO1ceq+H9UxP1W/19L4L5iC4BYCKjf5Xib7kylTMS4cw7byCz0ai+zESxFbVGN
pJMi7jaxFpImRG/fCEHKEM3lxwEcpH7cuN7cfJUGLwBq0Z1lEaltwkFLuPzItye5Ffq5lfewWRu3
Cpc265ryyJZ2gVwfvBBUxaiM0pPRlbpk40jM8i9k/1ne2SblbI4HsrTNWeJhCtyySMI+joIJFVwx
hebYHxa3gtnu/L9b5EkKr3XhHodHRRBq5Tp0+x4VzE+XJ1L8tdZv4//H5F4KZhh81yCg8zeUl8Rp
Y2zSuG3Qs8pnvD/XFeGN+FdKnTqA5DxQkSMFqTggDkRJgdzq1xLfpNv8HjDscUu1mryg2oNXENCs
JNoel7Zd/aPc4qz4ESrMHO2V85WzjdFVD1NtHQ+lItZsLQzyKc8RpP7JLCI2RfP4u65Y0asv8y81
hR5AsfKhMjzjL56m7GfwRLHpC3BsHbNMke35uGLrnMxfGaWbmAJKOXIp0T+8zBPqbmYnTxzmrTxI
Mkjwl5iM9kds7Z5fOKEgu/copZQex1f4LFr7fgX94RDjT7zJx2jgy7hWT0KDp7DSPWo7jUOy2bZG
ARw+Iu0cP7SNQjkWV72J6xRVdFiVCSVtDtDa2+BAeCgieh9JzjE784TK2sWHMrz+XKTAqJ0QlXA6
+NnqwEXKjKnZW7t1nEiNV5hgwq9/HUexMppD4rB3VhQfxyntsIl40Agp+D4andHxtTS5MKVnlxCs
zefiNFDFMQRz7+WY9kY2IAYYru+9Stq6IKEST+VrWZdqGegRBipWS15T5tUxpH330CDL2xEhFd1h
habj8leCS6AkT/Efdd/Z3urax/UwrXfB6brCX+oI66n2na9Vuei3SBWCl2+ryAGjyOcEcIuP7gsn
0OWud26bmRiJebDQ7CnGmlrwp5vRFqm3WYkyXbk9sFiy/fb7SwjKGuLhjy+RGmMOcY/Hy6w4e6GO
F5my+WUMd0+xjrcaSlSRISOeUwNrw3y8eEmnQAW2SzVE2thT27s1frSaWqzWtjWIqzxIA5AdrXdR
zvtCqalC0ZWirYhKqDHZgPTgDhOzsGbAc81nrZUZG2J/FnHjEFDvEFH8a3ImsIm1Jdqzm0Y7Uf5Q
tbBOt8sNJM71pHWGEb5t4PxFzbZ3SZ+9QbobGuByIGirfJ+Wp8/Bx7o6fcOdggsSXygR0n3XG4G3
pDR2l5YHHjUCS65PmoSGjApqDfN/dwe6vUcUnIkTj2Mr9NbK7vBfIOLRpdc03chYFcw3PAtHt/Hz
g1/7yRC/sm7mi36RX7o65Fs8OVqr7tMh6UHpDTZOtBJb1+zqbacDfDdYdJl64cVzTU4eecGZS8C3
Pdi/qombrkVEIIco1Iwb5BpS0mrqcKWctTHa/jXt1v2g8Vy9OFvLkYxj1fiVxyeObo6XRIEAPe/z
H/8k2LqdJDDKlO78X2hqbsFiFAqw5f8kjniRfOmDsXRuE+1PJYU5JbHHDtbfCeC3e2LY4FTWmF4s
JJ+bPuC3zO2sRwne+e3AU0qMH3v5RlFIyQ+JV6BWbn37SHCg8KAJJDzanCaEzdp8dBvQjluSQudT
oBBZsd0bnn4rV3ZVq3DUEscYewBpO4XAuvJL1uPogsiWe5OAy2Vxx+ahPXKoHdKjfYKKQTxeaEyS
PO/XbgthPtl9q0vq6WbTnkR6GIkdEy/fxkqW0CFSxN2Dt5JQDs/enTIOhm0TUUmn0g2Xg+dT1EwN
tUuPD90jLUZ3j7m9M0rn+XcaGIQJ8/YM6xByDsYA9gJqEQun+GDeWPyCxkLADzchv+6CxuS/7rcY
mI/RrSrjeYEvc+u/Oe5ZPo9D5Zh48usIUVzc2KUSxIAoKVepH04RSyiUAdPaxz+fOQau83nvj/en
NeqVuew58Fw4oL9qDmeKcCG1rjFELOdW2VPp+WxYUcPvvNHArRz63ZGC4CRSmqRww40Xmm4XdT03
vELOvGg0ENK9nW2A14U1oMDlRPWRavq39Q+LK6PNieh7wXyIA7ZQBRvWatiJNetYUItrzYskEA/M
/IWJ99sECGH10DSLPRhfm9fKfPTtupSl/7MNYU+NeUgUyWbnN+ilZo89+uzvTwctEmkUFU7W0r4u
elKIX7LmOKVpT6KY86gylqIT8dn1OG7WWkSKkPQA0lNg0Aj2OyYD1IiDpqhJ15WGpBxbM0M+0ONL
nUz9o9FvLz0ksD+L411IBuirsJYQHbmKfUZZHwHZ8ZtOL3RAk6mxubZbvV1VTcN/rru8++VdJW0j
VXaEQ8PzoIinTpop5BqH4pRvk3QILyTubVUCRiaBKLTyYHI3hqyaHRo2jikpky6WGBPIFStJqSbP
b8PuAi4dW+rdri5P3nS6aDS+5R9K4Db0bb0PaBVstcAB/rrC3uKGdKZ7EHqZIuiI0crqPYmfCww/
qM7ARbdXmecRDBF3uzBy+mLzSw3ayJKn2fcJRED2hqHaIWQ+kGbS54QpHsEIKctW0PkeH/OAilt8
Oi8pwOw+XfleUbSZ2v0dnBIQT9fxW+cnc5gkVQ1bxq+90Wj50837SWw9a8DrocNBSyPNkvrXSoyy
U0OeM3N6owjXx69sDUphdJ4skRDngu784fGH1+XiB+17lhVXIv/bU2n1z6lVfczmWMqz5YUQNoBz
Xow/JzUntK2KGymaPxHmcUj40MAL+hw1SNqB9LH2uF2Gq2vTh8y59ObnFJOgNJO9syLxkkLSRs/D
AuUTy49QFD38FpBpb8D8DXjL1osPCGSovRNrr/oPjAWaeyseBtbSjLe/OuyxgGMihmgH+wdXZSa3
K+bSN7rAcvYwkZsCU/s/TuAx/FPg7uQ/TNznBM6pbvdiEQ/ClAce5CPhD2iZT438Tv9Gg1PBde1T
3uYWQr/LT1d/t5g9W94c/N3Q6QJBCgDyx3jYpVTUVkLXIGMIzESt5yx6pmCdCirBBAGMrs/xnO+s
5Lug7gPyDWtJct8n4tVObjT+7TrQdjAyyrk6uS2+BBo5bhMRVKKUtaHiDnm+zN9ZnydUUkF9cv6M
LA7zhR9IbJ3DENawNwz/7j4Bri5Lx1WGlzSn+1yieycpAC2kxKuzaMFfy1Q+1LneVit9alaGnI5r
hMAuI+e5oMjH7rm2uAxQXg0QL0c/NM80u5HhqSesEDmrQyB01QLGIAOreSbNvVW1c+KvnB7BdM29
no894ioLFy/mpTgdx/gypvy1Xb5aFDLblpwy/VtR/EnyXpBGhKmvrAQ6jDicXmSkU5FsFbZ3OGc1
JsM+D+7W+GKmdYTV2kzyMJXGg9mLWvzq5BzAlCqmjQ0tRyqX4RWnZsGyuN+v5613YsgmaKNzS/Y3
KXgAPbr0QuBKBSYMa8Iq/URYqJENdqGB+ZMuJCHnojepjdRXdddZD4tjNGc3BMVIF6khoqvS/KW8
ziGBemM9ENwyoGKY7U9+cHuVnyCLpEDEgMVA5plY52ymkRfx5i353WiTMhnu74mUNyYmDJtDXm4x
N1GnuWuhkFRm+G1Jb2yDPE5cRC2G1Qzr4TmXtDIRL/LuGE2qJolD8jqgh0+9i9uYiRwWK3CnMewK
zhl6EV//gceVPrqpreWrOPLp6REOC+MbCRCehlaPGaglt3DHX89gh8BLnJpyUvwbaq/H1cDNayRZ
hKzZupI/3mCjaZaG90G8SlFSKuHoNZXbREnwvolP/fIjqYfICT8tYWExU0Fkteq4SUPwiSy0GI8x
XIMkLGxbGljG7fmtUzm+LppBcRFzutrURdwC5udY7zKakvsFbhZ+L4Qy7Lon6rHaHdcBEhozAdu/
/IFNrhqQp/qUtw/hAEkG5uO7V8radPGRhzR9fwkOkIzCmJscW+v+mVdJMY1b1k6HsTGot55dsdiy
Bw71JjBMVgXXp3NUw9vAQbbpozbqXASdkCxZqZSD0GiEAbVop6PYL4BJDnwkdp4vx567LfAWnJ25
HJyCbJ/5+rJd0ILY0H/j9EgBG3hFIiTwAbSuhSwHnBFr0SIKELj33E8xs5AipVGRTp4wqj1eRD+S
R/2hFe0fHrZF7ndSW7+yROsea4iUvmoCSWPlvla+l4haNMRPshDjCKvFwLfrpC/485FmPosiTh/5
hLMN+55zNETVSHeRCZKo6/md0Dc/NPe73IS8S+w/4iTqCE6E/r1H4syPbu93PD7YDeSsVzkvSJM7
LDsTzSE8kkuWdRzYf8Tg42ZYkhNAQVXiCNShdZ4DiL2DBruUE25vFDFYt6w72ORuctQi76J0+Ivd
3XSCT9ONWMAjtRX7+jBhUty73zP1u4MnuvAoZNAgz5koqQD816zTELmpUGL1HJS6avWTJtTuvxLx
AX3FLJs8tgog0TqZYVWyuQi5h9+4GPLcQ7t5GxtoLvAoXDov6IS2VFOyFPvlX0y9QayTIU8jAxth
R/xvwNSq+F603b1/rIbzpesPXW0crXj1AmKcAfPElTtDVmw7BmfBn+YaNnAtx6hvwuCzJlQlBHyo
7i6Nn9b/hlYfFCWf6IYgmhB2ZBi0jrC2LIcStk3zqC45HNWiAJYBGNgS5wErD6v5uzKugs6gs/QB
uwqb1WDdC7Pqe56hlThmAqFPiOhWBPxvzboR9NNe4Gj2Wl+JE4oeBT7O3/Z/XqIpJWEgI99Q33ij
iirugvlTcm4eSz6VyG8Jcfp0k2fHUcEy7/YPWxIiqu4YxaNT+sUp0oRqfjecEtYR8yUWfNG95HAo
NcPMWvfX57Asj/HmB1N1vxXCFUWrLE/e9fWfcpwrYbOXhEtpuGoQFrOOISXJsnfxISrTrbrltnz2
JSbtGmSSACi7jmgcbxS/D+NmTxlb+xNTFrDtDC/lf0jrE+oMNOqQecPp3EAn2FBwwgE3BYlmA6Cz
mcep3SbQoE+1PNDRLYi+kqHYzts91UVxVPm4wumAvT+ekKt6j8sSuBR1ndyfVeZDRxcpbuTOqTjD
vlR8yfXsUbqC+7kubHKczcTJS91SjBntTDO8Gh1qLtRHg0i4Ilr/zxM0XcHPqtmZR7gM9XQHxWY7
cUlHjB6SpdIUEBMdDRS0VmF0QDDEQnOTIsWNKaX8jpQ6Ix/sC0JAUm6BuEHhyOP4xp5oqjLwr9CN
i4Zs8fYdfD5bQ4VbZKpKNBWpbSNi6D/+hugJMoMzDi2/ddfzPXUo1gqpA1Jq2Kqeju9uAZ+oy4u3
/lxlbR+jZYs+7skNcx4432Sf8cc1RshvhJ/p2T2psbVO/dy3UWLSR0EPySy3pmi/zQUqA4GQE8I1
F+MjvJCQPw73K9o/VlB2Gt9ZpkmDDE2puad0Psp5mJyBk1XsZWvl2EmJaPCeEDs783xzmIfmr2ZJ
syHLzO+UysQTcbuxfvsgn8NtthHiaVyMTJurNWVnQlnEQTm5Qq8TBD3K5cro0mWa2CQrQsygn3nT
Dk4+QqmKqjFnZkPGPH6Zs9NuKslbu4/3i6NP12kom0gnno/o6e2daQL5ABwWPNwmseQ0NBo7HH5R
jUUFBo4A8DPzYY1I5uqzY8sZILQ4mZsG3TkLRcT3OF41bx+YVXtLL2pAFu2Anc31pW1+nRpPW8r9
vQuiV8fP0I25m7TJBJ/My154uSKUnbVVoIYrpWfmJqtqHRsny/1bXVesdFiMFISD/lOdx2gZO7kc
AVG+DTa0XPu/Dzjy+b8F61YyBIZXa05oFvN/PlWoatMP4lHB0UKtHwlfZoInh8Q8QqoYq8WPW8Bw
DrvCQne/zmcwhEtV53FKuOmjU5TprRY6xGSvfui2b+fSlKQnnBq9/7Rf7m90eZN9DU9NrGevH0A/
NmabbTdUpTX1PbqHdGkRX3dEBWSBExSBCKedmwqJTskJ0LhZicpcmOdr1dxjjOZlJlyGbK35d9Et
+VJ7acLaHwVo9gZzwhc96565MKIxpegaWxgJljSytYyqjMXl4hdnaKI921CQEPnpZLuV+H3Mo+bv
/ogqKcnGX5idBSvt9C6gYfUboOrrkM+KU1w3qluWBt3w+drAudxifQzW65ypaIatmv+8vN9tTKxg
Cr7CAzIY1a0GkUMyJKAJvFxl7/G3KKCrRXFYbih2otVHclBx6HYqodahUUWmme9btIUQ5O8bdW7F
ncSrPOGVoMePo+/Iwi3AvqeNmUiTmhQhuStQLTDGQFUsnsYR9p4GBQ37EyYVpKmBe/5j0PQBdXsx
gb7ADp/lPMaANiPa/orNHS9AKR6Y2AXhAwO3zaOXu2XY0AHuSESOKvEyH7WsBYZ/I5ReRHhZPVLP
+RoFwN6NZPgPMQZrlqC5F36Y9tEfVOW3yiDvh/Z/lnL1NW2Fwn1NEAUvvFrOsQjzc8lMLgM3SHMt
fTUztpfjOLnXdqzq2vk6mVrpX2B/2TlP0KdMw0jHrLfrIGq0oOFeMVwROGBnhHdHtMyrarxI8vsf
O2EK8Hui2NS3zJCUnNWtzkaIc9uYr7ej5v/nTvljeOZWIopUmLayRS0K0XY7dSw+hbjtwAF5kqmL
ZL+2wSF3ETVdNGBJwmo1cTQ32Vo+lUAKIyOzpluRatDZlbo9csO4/mJB9jsol8Q5Jk7JMopJQcIT
StZgNFWMl2d6s9+e+4adOad6EC1SR4l9YfKGDrljipvMpSFZpp1ajJoWsW7OExCDAv6eQp9HEAUw
GymaAGy1hxrQoG0joyY17HO9IaYyU8XW2ituKqV7nLSLpNAwjUWTJF2vli9Gil7Bbu4KONE2YXm1
4HWme72KeRTf0lb+4GaMp5mfCNMYxhtUW0lUl/ZRhUM3SVL0o/lnaKs01vBX3pbi+3u5kXrMnUb7
9SkVj1oFxRbBAhV3K1A/h1e10RRdq94ACBz93UPh9LETF8aWelRx0EVBVJ2ervtJhMT35ZP+Muzb
nw1/vQ1sqS+ztHGxIXDt5fNO7deDxjpYMchwHmHfEFyt2vxwkhCh2taF73uy2w05GpDDXRZr5f6P
pJ9PAgVO7+Hj1j67DupAZH2MjFUoOQ+czaqLkvSiKGtKJ9rIc1a6Woe5EhITA+xGiS1ngZ7bkpfx
FuiSk9R4R3nIQFCKQ7Fd/ZfsbjKC0QBfuALCNjUX2QVRL5fwxDNuFwPRJA8t9Z2Dgwn1kvcVC0D6
L4vkCcmVksjbEzZeKigFzVPFmSiuX9qfuFIBzcBWvf7IDlqwVu61K5PGAdZZOMhBvwB2P8I2zKnV
USWs46SkU60XQfhSEka+pELZ9hyYsRoEHK9mPOzLCUdxPfaNM0sYpRQJvxkB1diSFTHufwui2n1K
gJoBducxYrtmppyKJBgjD8C71dqQxPuvpDiKo9amnojdmIGWuIv3TijQKCMfB7TviHUoEdwyofKv
73pCNGS4AIfMwZ1oYQa5PzaB44zLcN23a0JhS6z9WAnUydK7iJAKE7J/M8qfMx6ewZlYblyLLVZ1
zR/5xSOmCZA6YALmI7d7Z+EDGujBR+zjLJfDhI4+xLbHcxCBbPRdoSP4t4zVQSNlKU2NMjMjphbv
6KrYJY631z8k363fx92+KpNb2q1x3p/q54epfZLEIB+70xxl0DgIoawETLrpsNikyOwEbvE9s0lT
vDGqwfFS+pv2hT4iGD6WJhVNajNOONDTmU0fyG5R1FjSNas9+rYTca0Yu5o8oH42/FLpQVMUsYOG
d77IEaSPiSWzNDIj68bKk4C6JaCM26VA4FLz20bN8tETSun4M2eKJLq/0M28t2WbiMg7/Dl/tU51
RCbrV9X/fJdQ6qA2z5Lp+YSwHGpXVLvOT7aTlCDtUxEtfQ5K0Yj50BBfsZAdiAlwCbMMvbTwdOB5
AgmRrfU0dhITch4odnwzjhCYzVudntHMiB4WEYC4ausgpkpvAz12G/zVueapWD5cyJngDyPC6ubk
mUugMehYduXqfoSZDXsGGNrvdOFaHY9BLBiDJ4YAJj2IKy2bkrLAQjLrOcWSBefHKwlllG43jS8/
kFVROjnuVbvju/2JtHOaS4YwLzkQvTTTQbDlzjcCNjPga8gf0Wp53qs+KR8xBqmUeN6uX3wmjtTY
h3sIh8z2IpxbrKQWPWgSnmO5duhmlq2yeSp65eWrSwGxrP7XLkaOU8SRMR9Isjh3NU+VVbfQaNp6
f6sox0HxxTMZBsMUScr0YksnjNXiehkB6edTOrzFv9X3K1L/0UPgOxRXPm1JjjbzSl+edJ6mudf2
mYgj4M/Omf+I81bC4x2s658AZc+4vxwe+Zhm0FKO4+6T6+8Fb/B/uJNy0L6K7VBor3D6qxz9eFSE
1P1JFz1XhZqeoDyDp+Qp7UAVs8OpqEXpkAnkKH88jNEoyL7ypbrwN3Qg/RlsVglfzxPtH+rNYBhW
+1IE2aaLYyNXIk6d1H/bhKWV8IKd3E0ArSKwMDeUQsWWlGuFe8Dxfdn9nG66IgsG28Rtszeya/DH
XU+PYxQW6P4XXRBDzFWTPL0ThrplCIMaavZ057ilewOlMtBm9CCUkLD4ke24nT5fzIy7Va7kb3Wn
bFdD42hV2p6ilZDAOrgQlDtcmSjMUn/DEVnfGAr0F8JbvEjfO46duk8mMR8cdC6nqE5ihIm5lDHt
klxsd3NoSGs1c+s/TieSwWrBPN1eoiANobfhKO+IEwWipYh3HZwpouefCVWGHn3HBgHs7vNVB6xT
CPooD3jI2Kedzhor0QTvAZR7vExIHyEIrZrTxM6SQRSycELakw3XuMCn0t9Ij91/DGo1wzeU2InL
O9VeDQVYrQ7Me26fDpFpEUUM/g6bN3r5YMekK51p683KLrIvlPCDVzVr6x/Rw9ch5VVnX8SOJrbJ
sRdU3UtdE0mm2FATF/9RG8JanGpSIk7i1B0CZtEY2NrZZ/o7iH/ZjJ8gyawnrSdinRiUYN/XqT+E
ayekQZo/gcrWagRnyGhsWKAsJz3+93gdhFPXXcj0h9NbGzGh4ujTJfGSEPsVpmSQLoVJetiqn17G
0pPOZKrfnK7ErDr5kKKqKfR6WZAOafD0giioNz06navMkSLjB0vlmIWWz/5a8IAQqG86YbfsdICg
0gDux0uX6TrVIxp8Vct4Y9x65x+2D3mo81ohxyAQMC7w9G25oZ/jNIO7yr2DYoQeLQOfwHAO2iyJ
OFwGpROYg5GvqbnRGs5IJ+bnGsTY6gxlkPXBuh/fbsP5amsmQvTLTl3mlngPKCOWRMQkDR64ACuU
PJXGrhGvqJVLwWK7Q9H1G8fTo25OkqA47I9/IrzERPKXetEzT6p5bV75EF+S2kS/pf1AOcI2hKZv
jZhJ7Ar4pUieZXzQI4buB9ghR92wL7mWIuMgb7fOhxMzKbLsLbiDcmJht9nfwX2f8spAxMJauBcC
0st1TIv+TSw30GS16KFAYeRjGnRrG8NqNlybIKb0vGehGmrDshfoDIqSH/KEqrp0YIJZSGW614ah
fJ4eR30AlmGAuxgYSB1F7MqnubORqw++irEbe4tEAepG4O10o3rhfhBCS+gfu1adokXkkX+e6YCy
oJ/q1A0kHXi21BEhfN1Vb9Sf9ivywGYSlIKVv5w61vs8s+gD4/XKvob8uizxvYmhVeyeq2nAWM8c
AdO2FqmI5MVEnJWSqshPpHuvWykZI8igQg+463QCCGDLWiYhbP+XJjkTx6gASHhSxXxpI7SPs+x+
QjvIT5uB4T+Lla//4uO35VMWFxuZk4MSIbIT2z6G/yJHOWiBqrqBrHD3MYowNYZuyZVFBZXo1o2z
58siLbBlXUrbGdOpS0MQWZnKbWS3b2fc6GTSI6x1TpUteiakqynpzEihCLmtjOvHX+rtpd3FP7b4
mLDUDyJuaHq1sXa4vh4J9Kr9dMGqvS7M2eT6xJkB9sH622v0UEFANozt4kziUqVxAKeidK1vyf7Z
5mocEkmx8clcyCfr2MFVTLHFBpn4MrP+55V3m0e2MG+t7iR34ITEQ6EQC/2ja+ztlpUU698zQpI4
MMHOYMivEOu1KB4JzoG2XiQfHh8XW/xIWlohZHBM7IOLuD5kbS8NWp7uq8FH/RmdjkUxfXf6NPbB
OfEzc8AHOfJnMEIDNdgeLQD5bQw/OvrIHLPEjhxE4fBpq2e9MN+b2S2RsL0IKtTubPuFSlQzqYeE
Noaf4Qs9n6yZd7wElVAz5aAoiYAPnpNYS6ZkC7O4ccAP7+9wcUnENGwx+CNZsyNystMARD3ys0Ui
5uTgMgZL+T5YFZh7MBEgTRT7J7M+c2VTi/SsZ9FH//nNAXpGOT2cUr8LEfHOYj8A22TscHZI6M3A
D+W0G8uKPVBpCh4E/jQac7C1Xtw6pgomIjPtHbEIQY0NjOAD0WDYGDniHcHU9ullaEtfVpRViqhp
3s09frONWyxZ0EsNdiBrKgtoaDrZfRrlKxFGPbTsgXllXcS56uzT1I2e8OZlV8+JTSvGlpR6Bv9e
Wlis+A2Uwsk9DzUvYHXMOATKhQynS8OWHVfellkn06OslIZC8uRSMiIVDlqQ4md4YgGyJeZ9qZC8
O+DFj1rRYi2WGCTIWWZDUEMcCmRfJ6Emd5SCeBPoGcht+NLkKDeZ7tYApGJACe17zOY+dxignQ2l
cQvdfzuxYj9Tya/keVkQNsRLg8SjzG5lhrJdHfx5e9+gc/ugtlUG8jFE20XokggF7WI0ijGS4ASO
2oLNH05yrQs1ZFv6yReDoXSSyongfupVtF3FoUIfbvmPO7H0oJ3pwwnJblQ9Myj96P7/cGeAlcg4
q2EF/NbpXVLEWkDPkKH+KhyAXTOYzeXU1htXbl8NtMxCWorN/aXcXShjM8nFo+s6phWHfq3L3wDZ
AopofxOxXt/3sFzbJl5Ws1rdTv9s3aRVVucq+c4XmFyqiA99fC4DOMBrHPI0H+vL6Ly3Z0MigEvO
Xy9KS02E5NSAINK63r1SY65fxt8OLyJcFooVSrTtQ1UDu20HQbUu7fnHS5yKfMx+WBKKzryrJmnt
H8ZLvdpoBZiFNUV3dAXdy03ni8YBDzj7rkFZsxDoo0ko0dARg5eX8Dr3ubRdA/XmXHofPRZ80ATB
GtsIe1KBvbciUNq7iZscVGeAblNSjyfl76IjpbKtzD+nGg2wqCnZze/fktBSRq63gzJVAcmHZddr
95PfXvicNXil/hLxxrNBsLuI4Vuy5FCw1jZK734MmUTuGA2M4ahn2xOcSkSrdgjJJwl3PjdC+IVo
WACjVn7+MN8krVnT+Izq0EmO8cYzPEFnUOZi8rxgfGOnMI2nu4aowNLfRRkb7vfk6TYQLPvfzUcY
UdeFzsOxO6dlN7Qpom6idr8Sp0r7Gh/jJyKsq6rXL0tJ/7QrfAjRCc8LoPr8dhXU9b49OBjnunc1
GEGLw6bDar3xAezKKAtuyUeDWaJa2xkC25I9f/nmkzVzHviH0j9I1c+fxscu5IuB5jSo/WQ4SATy
y2cVE8ZWHh3XOwxLTiowzHP7IQlupfvjrSTGclIgqQjK1XmU7pYwiW5K8m858Qv/aBJlc80hiGPN
WwuRUoP58p9CdawCFujc/557D2E7a6UHohV/l672IMpcaSVr8HNvYjNP/KyYymBKc0hsq3kd5mnE
fKqrNBfFTSh+Na0PtagvHhzageiv53KDe/p/qSATwjIl7UT4pXGGpMbwXIGztFAAB4D010H4tIfS
oa0gqX2Yjtei6Sn7LnRKXGWbFGPmbCBXO/XN2WA4u5hY3G/f1vYKuVe3ZZVwVaqnWo/MM19VyHow
ESauGpTTsGQU4wfzDkYetrgubo6Xeknln1SV7jJxz/rRX4lt3pu63xKxJikvJ7ksqDF177qYcteV
9FuNquEtXmxgxuDRe2rwZZ6cLT1M2ioPSPWGkid2tpbfcCKyb3X8hNCSdxpLxqtxj8LVS2JkiRgn
veDRW+zHYVvpLMt78IDaCTf/ye78PU4qxPZoiHkk5ceBbPJolhu44aU9atMKrpKt844aoJcNjF8V
DLLD3rWjRMEseeEclmIOst7VeJ01C0KQvvTp+CqUc8s0CRjv9CX/3MgLtMQ5/rjYXplJJALm5Xyb
f3H7fuGNPSRy2fNcrywxrF6UuAw1rzSH3vhhcSWa7Gz4DqiGGtCnHBlbOOSWHNcr/cX1Qa+DAkiL
PzV9aXbZUhdUWVObJMaXs1aspGpX9oRRART+2twF/+d3nx/bXLjsCW1IDMw7te9w0e+SJ9K2Hm1q
86HlxP8uH1ZEEq1vLlUjerlRxIEYQ06t+x2nX5F9/DQW1QjsckpAsCFWv8kHkd9FWooE7ofYf+Nk
UTlBLqtM+n9a83LtmXCJ0dRdozUDJK7fGva16ZTl3ysYx7zS7xZyjmSekzdoZ/Zx/lQZRw2rWxTW
xK8b70O8gKdajjdptJqabHFl014S4AFBiXGPSt/AQQAAdZUtz/0911H5Q5VIdliFHJgeQi/WpIiR
VRosuoQb6eIgzd/2VvVw5/Lxh7AewBsfmbyaFyVL+FMcKix5IHgYgYt/Z/mLtc6N8WrLfVGIF1ip
c9I+SgBstd5H7FBfW5iwNHux+FjLqh8rc4+X3oEtA2IIe+VRBnhPPAqAQuG87U9kIKhDbDIchf6H
LeRLkNCmvuGG3TlayvSHMmeg7SeyZzrnMfCjVOrHR+xGotNdia9viO3FDMhIlb7rfPAF0EI9zJ0T
9bLjyX/3eflETgMYj0bkMnAx99GpwNYbuVu26y0xP8PXVs+VUkb9CC2CG4FTrRM3xz8X+NrVGMPX
FFJBM9lmjBK6F1so7+7ZGkJtGO7x88NegqT0y2rCqy+4Rwhgd6Z0od7pcAUtAp57KKipwXusXvB+
1OVnAtmcrfKUo2PSfRhoHo1BMUImGzVT85AIWluaIqWxmtOyoh+yPC4zZ6QGRYxb/pqJGOBW8e6E
HTWc2VDeQdtMfAqFfC84MJWRagbabx17OKhu9Z9wEmzyerwutC+ZQVH4JqTZ1f3/Dd+7BAsnrVUt
O6btYhguDfsE8tYoMZGVB/K1YBD2qsoH5yRCRfCSYafItpQh18JJaiC+p65CWh9u83xhTfvK+uAO
a4JlG3HkDeTAUc0jpc4m7oP9fpbBO4+EqTitMiSLrXZu82/rKzVc0sHEJmksvffoYDfUQKWEvYdP
QQAm3cEWmDgGYojkOwJ9AxhbvXWtkPj+UVKeOGXg4A0F+HyxtY99onXSbIqgk6y2VRTc4Q0t+NUX
nPu+fyj3Y7QndAwsk7or53Id60SH+Uw0UgMCkYyqDLfL7A+C8v03HXr2ggN/ftR7Q1wtautgXA6v
98Qtgbinb5TJO7WBqYCTQNPHf3WbhJrFxFZSMp7/ZFCGjYoYxG6Uo7NnsFG5FDre8gJYm/ONIInA
+gJuTtXiT/BDCbZiMlhXh/KXDcWxxTdqKdIrPiFbGm25wxosEJWoLEkGA3daH5eSn9uInAptfMFN
FWoWmP+kbUa+iCQY02WT2M4Z4CvkFdlv+B92bCxNg1lSmZfh0H0LHf4jQKPbDyIx3inf2EeFH8v1
YTISLPJuduHU4V2KlcPa63FI5ASG8v8jCl/fjiqcIj8zoz668OhGQRVPN0jMaURDN2Es1FV9s1we
PDgtHSy9bLH0K78NAVy0EDKapci17eDAOMjPjHl9RgeVLpK704ZseITx6UqD4cAwjZ7nU7ecByJy
dmbOnXmC2CIVMy2Jr/ep9txyOnwFo0aawy0UP/o602ZgFyMHpqJ7qS8ZnT4TZSIVJBeHGcPjL96o
BDaE/90kAWfCH4PAStLPc/G50zN4TRYZzJkH2XZ9sITypW+F+V+Hl0zZ+LaV0lqC0l5j9C8hwks3
w0JZ8j1hsJdpBLHnbTkYdVsfnpH9VI87gbfuO0lp1v5+Du02Dm3/amqPRR9TiKhT5zuFF6KYIEtj
Gi+OVTp55h+Ipqmn+yG87Bvbb5JCN4j1detLcG577XLnVLDOw1UI3kUrwS686eHv6RvNJCRKWAvA
I0uE69GoSkO278dtTyWUWRNCVJ6CwwVmvQt+MKzhoX/jx/txvA41K9RSV+zU4gYR1rM2O9p64boc
XftFKhkwsvbGjfVPUZEcMQ49gDDklbqbF2L7pXLCuBTWBwOkCYfeCpPnTVhY5nHAcbuPWlS4vGdx
cbZ/N7HAyyfHZ7mv8NAO4is1llZlqh7lsdsdMHBSaR+mE9bd6ZIGu3+OoOorjXPMajPMdJbszh3N
meCNBB7b7JW0eXVYn8f5cAcuxezIzIV3QI2VpvZiV1Bi/MFqnq2Hw+WbTioKYjuIBmBmlcnWFzv8
DELs0hle1NORUuLMpUBKNqghIFAvR3tnGCWwjsznAwt3I6XLiOwSd/5JZwTIPCgwMT9Rw8tWL0KW
i7HroWAp3aFkWsWVGROM44Z3pnYVHIe4lgCHkzf4EV0acgysVGcGrNtTIS+Or/h/gWe+4r97l5EH
xEAD5XuhNyZkx10K+84X1fSqoxsJMNfrWRpyJZWLDnBCQXdmvFFZYVs+X1psnQPqu1cpM2y8GvQF
AQw6dx6TaaHRXQkr92felmCfYD/HU68UBE4xcnc2479KcE21IexgKzVuj/FnrzegEjNL9HrY+ekI
yRGakOGriGqXzOsByY3qllJKGlaT95KJj/TUQTSGWOcDzabyVgb3xyrT1ZhqURPJc54s0OYAveGW
WOMcaiHrRoYWGmPi5De00br9KwS4DIfqU8yNy5TCFZshWclo85mP29NteFZ6EparZ7AxF48xSSFY
kw1JV4ORN7Ga6SqgIEImnLiZD41kVsKwSUQgv3mfLFk0KZO66DoKodiCcncnxYcC2cAMRzIfm8aM
wfHCU7DSehGbuhhzW3Pc3Zd2U7+MIPHYrP+N3KkHU4tCXnvf8fnGqT1eu5k/LvrTRlI9hNFt3f0u
Mf2g+iDxm2NIoMl1Xcxh1EGMYPeVAhylBD5WtZ6siJ23QEpoUp8/Dz9Sx7ZN9CkhmTyFRNDZ9rno
ggYFT7E4vMIKILjAam4UnOqiSt2WZUfJReExMMl51WMUlykvO7j8N/ietotkpNo1kugZNRsgcnqK
AURsC3HdorU8Migt6Tyv4Y5tURR8bcJFNB7n8/pamESqTsoPJF5431pDIFkRo8++5Lg86oIuEd94
rqvBJ7R88AT/Pa6G3IifoHbAUrCU8XPGVXL3vMRpOsKO7+CSin8ZmRengP8hwCQWySXsJ60out2g
YIyplF5pztdXQ3yiD7gZUxHL4pGCEQn8j5NVaAz3BQcy/4LQ8p4Dx7i4hFn51supsAs8Kw+C4tOg
NTkzUOefAYiKUqUJVnFJsq1IJQpcpwmK2K9fj1WpobltCBux+uD/LofCUBjIuvBbkLOLeaddrNfE
0hvINnuO3MbKGDA+o3/ZEGoekeNeYjgV4sgGS+3OYyVZTQXIzvL+TNo826TODO1X8Iflxc/Zj2JM
FMzxvnw2Y1ds9oNbuNT3fvL86JF8meFEiB+YYaWjbANeB6LRpcHCJmDDhz3ifPps0KdfU2ZKsTB1
2j8efNyBP6VhaBZXA+/JRoXv+I3ST2GoXWBy67Gf9/5Z1VjkU/snqDsxC+SZ5FawY9UgnyJf+Agy
0iGYdcODop7MfekrKZOBbwv72EIytycP2zYOYNdmxyB1WJE13xW8CqZLXMga2Ubvz4JQjZ+98wj7
N6Psm43zt06biIMv/XgN7hscI0e5V9YR0beQrhozyVbYALEAzZDMg2924raE6iMJ+nS52V+2qSzf
qBIFikkOXX0S5aYy9io9Go1ISlhQiuKff0FeAauFSLO58g0Eh9Yx97tdSysWx3QgHMz9GWh7o9LY
aLiur1eVUlTRrsNFuTj9M+wFtNX79kqnd2Dju8rMrR0cLD4qwLadty7ewSelQrLYOHChjbczkkSO
0nlImH0gTE3XDakbsIzCgY8MTZRaxKDISPDHjZLqV075GQVyhC4Nx91tds4BuPc3zaKuPL9zgNpV
f3CWrQPurvYtGr2FXmzfDlOWHaErAwbdKIuyYtAJg/KFXGoYl66HxtYmncpEJhJIZNUUuX6zNH5q
YdOC2oP6ds3dOlFx/6yezi3gUf0I7eTigL0OGE0IN6PRg32ckkllphCeExGo6xgdy208HPXlV3NJ
bFAKqzccJMkKFUZYtbyXGRRnnKlOJA9tmEOmWB174UQHqABV9m+kVQOGp2xt874fW8Uah/eyFdw1
D1g43N2+wejfOONjQivHUpN6MN4/edTZwSyj7wcVgY49Aivyu77IwKEYb4pTArYZli238qRFhZ99
N28a9Vo/vsKxwc/4yYEtFl0MjQJTm95UmKrLazzn/voOhYnIflS8rHmScD80UALxa8l0DIiZdV0U
yWMvfKAZq0EpsYK1nohPmo+s3LKFhKoRrguTX1sSGCyyzqO7nvhbrkFFOS/O12rMTf+chB6FRDfK
muCZGU57x+sqTgNQLPmbu9mgGEL+rNhKUOTrsf//s30cNb98rmPUtC86VJrJtS7lHuVr9xz8lpsM
9jCxS4QsiMhLgQ46KnxsIXKyggIoNX4hxKlw6fqfHU8ULfHB++phI4T1WoAb+OP4VMr8Ud7o6EiU
EXdhS+6W9lrBGhV9+iQTZ9N3T+hhL2pTPDxDZ3KyWC7mw9tD4c8C46wI1nozg5bTp2WuJE5/U2lQ
jvN7wcbWAC0MB59rRcc1s6Qx3st+Wrxl6Rx7qybFv9rtvqJ9t1b9lZdc2aE4rd2SDTb3ediWxwz+
CLaBdcQOxbiM7ILdi/9aixT0Eu4mF8FGjWIwDIFAbZlXH0jFdPHnFkLuSw3kno/vKq1ngdGKz6yq
ZA8Xgt9rx9lq3i153+i8CwQh/P7EwQic1WSHxHq+1C8KbSV3hMCl1gYx9JlIMMoEfMQNsMhrgxGA
WUDjdxp3gb4gtsR8k3p98C1qSQWdeWVCzuRJTPGVPXDfOvU6rxyyZdJ0z2tBWEpgP0VQQYra7SqJ
hFnsaJNIIg1PUnXGxtcCqGWrXHjeV0cYd06LNfus0IS8CytWJylcGO6oROE7LOAgiV5dMUJtcHT7
hLEp5AGU/3l89EQlP3KYv56mNB1RLmtKIgaZQbeufY2BP/9lBBlnyySrpy8DYQD6AkkobP29NTW2
1cYN2JywMmkurEFpXeECcWa9l9QUz5tOFRpsXk0Hm9WERjNrkrfkZdw2IbsYTm5iODDL2TMp+8/5
Su9b7nwzgzJ+KMAtxthp3tFQ5CTwaw2/XNTnO1hwRYzwbqqM310YhYeWcJ4WDTT+lnFIPLj/8vvz
fwpcMbtFPrCn+sAPx2ZB4lWk3NSwx3GOQMcoGwNZHSty/F44RuzmOhA+ReUHjESua4uG/jrXj+2h
F/tdQ0B47QZy2H0YS+M8J1SgaQMC/gC5pzOO9D5829QIdbzavz7pBZ44zF6+idawQVkwwqftw+Kc
Vs2wE2/423mD/SbljSX+eB+OWUnJ1mg9p4pKmHuvmUBnbhb0AzuPxcI9ibciH6MQZBSnutoOmglf
+WYUcEdUgNOD7VOWi5hKoSUF6Rp3/TOv2fWxWhRzJhWGkmyZXeOmUvogYo55/+yl3ETry/K43BUL
lmpAr43KfWNLm0AkJO7bLGx/SIsenMeYWRB1LLACtSxYm1iKs4ViBiPYGeElDFOg68bEQspn+sEd
TTdbPwB0MbHeEU0scXofM3coypZd0InxRUDED2lh98BpggmvNNy0yufhFktjLq3E+hoayI14lAXJ
LrYRK+Xb860/7MXynUqYGyhrKrLvR/M4Bi4IhM2/XHhs39uP3GHoDD0levmmW1HLqoHR+Y2XNfV9
qwGeUKUxkEGDzaAtrhtdjQh0ictTg766LCC8BgX82bW7ymCJqriWMWC2XsfP5mNaMvJUJVrt5jKC
VyXFFnS24qCcE7q9eXnflv82720scQKQ5IV4+yCOTnx9lTQLMHXeJF+2QMtCIakYOYzlDvZN2kZs
M99r1wke3cO7wlJQyotI0XEKO/IB1FWT7zmUDEjVZowZuTUSKAzpE1xhhUTNZxn7pfUnaiSgrBjG
PZMZJOiFNMXjZ1XxiwQWZTtl9q5RwqCvCIAlcJEd65vxF6EEZeCyti/OqUUNSGkI3+x/7V4RME+R
lDuCu3JwFaglSltwjhuukQRURwjdGnRCuul13QZii4tPPCwiFXXq4rJjKAnh0fdjhxDZZwur6tkN
4RXvv8c03T09iDT7Nn0aEDMeAmfd4uALNTzWZKJAqQkmEWg3fDVI40Q0LADpdTHfvQe9mePlleWk
2AjNIbaTLmOCk1WTvQA7jcLLDXisnQANDu1lKrBL0n6XxvKIw9N6+ysIXVSBFfopqwu31qtDrpE8
c2/2e8EU2D9WPyjr4dAHe8QkwZuGpVyoLaFiSwVXJS5XrO8JTJGCVgSDmKojC/DUqglSj+aPpeOg
19bntc2Y6RP3fiaveC7EgkZtVRHT+Et1kJNiXvEfxDfYzi39xByTsYmegDkla1g3G9qVkIncGCZB
Pg1rGuC2drYXsJBvyPQz1iMUM6p+gLf/+8wzaOfohM4kjWf6g8q/YHzfxxZYQ2jbBJiuWqPR9ORQ
uc+DiwpsRAg2XMvqkVTOiknKjuHXCQRXaaxgCQr9fkOZd95BxIo98/p2h9LaawcGz2E73FSYyQZ3
JLHyYQ5oNubpwPDilPeA3jxprVjLdWlGLPIrq9RhdwiKbosleO5XX2a4vgRF1YJRbrgNQXifdJkA
UibsewjkKYGK5RnhCSFxFaprVomjm7YdAKfiAeJGE9emtsOucu1jzGmxuqbA1n5S5LQQsSfpHVLp
7qY+JxQ9Z1Zrqm/sOKc/FyvPR3h1YaFYf6a9CIBM3JwE204oHEDeMkur2q5VzqmVrA/oFBmVvY72
JN5hIMIX2mfnZwYINmpwZ1wu/KsezjYdVeJ5P0nlpO/mOypuZcfaZW3p6EB+75p43sbTolRnFGhE
9chfNhyAFf4ReI6Jx6oTOSvq+2AXYQqhAJvH6Ohx+SQGI6m4JTn1f/2cnEIXc/24ChMYqXaOrwCy
TjV0JIh6qqZvNebYayxa+V+QHLugOKuv2PpEM06ZyVvxkP9hk3ncyILcUTZD/+KJ7vVlMR/Ppxlh
Mc8JOuER9pySTWHz3rXC938aBMAC2HsysMF7NTe20/p0iApzGMQJBqwpegjDP1G7FxeTz1uxtYYs
AcDhXM243vqNoryruPY+p6oOnfwBbvZuh077ZgXRmM544o8q4orwRkRPWh3MTTD0eaaiHq09cPPH
kaTePADyHd5hGXss5DmqmdN/Lg/BVttQuqN654ehrfQrkiJc2ew7sLIr21rndqsYcngYA7tbJxZF
hgU10BgvYE1M9cGFhmc3Ce6CJn+KTb6UcdvMXvhjTDfyTC6m4pAXMw4OMYQyf+atlWEo1z89Ajae
DvpfjUJkH8xHQWsbheOqhbE+P7eJNtu3Amf5gKM2oQTLhGV9dHkdF8T1kQczMEsR/fK0AV+B/acK
1CA/IT6XA0Zrt1FSzmSwE669jNoYdE+tjjPt1Fevv8YVWrzfNnOT928eHiczwYmmt7Wj2C4UeD76
gTNJwjDPLtyChoS+LnXOvRHitcW5xtH7hQdqX/szgoA/deVhrL+aATNFLYNWxWLX1R9rYld3wHD4
A3nAeaMedrnJKbxrxAjPQ3qzEed4LUEJ/KMm5naT6zEDCv1j/qno6x9AWiBCOu6X9EwmjEbtAj1B
8c5hStTUzHBSVyNaMr08q9lBVa3zkUfiMbiJtsa3io8Yoxfxq+svdRVmd2+VzD/pRTWUblZrT0Nk
bCjaG+gfMhx5jrZZOXbY43Gm4c7uaq0tuVH7ykwmCqWGbkcnXC4fTYMWEDsTj3TxyigA0D+6Whhk
qsiOAYr6QOgTTwgwYBkPXwO2DIGSw5uyhZx/iVx9WMVxQL2nDZUytTYZZ5VRoHGUPEjeudl4L06k
Sj5Z/IRDFLO8A1T0L6oeuyeBFAokcgu7L94RO2DI/Sw8iT8HR50qkrgE5sSefH54/jZE3LxtGTOx
Ic7CXUZZqYMpKBpjsxR3arChrsxNAcVutyRZ4barDcuM4tAG44vAtr3tkfBIc2KQp182Rz5pBJNK
sQqQl7f2Yya+W0SGHCkRogGNRr0b/WPIJ4BEUCrbQ4CZMsMrSVZ667x6RemkyPxkeTcLBY9vRjpz
D98y212oAtip4jMhXOW09b2DFkRRM2cVmwPq2KkXB2TIlCCoNLSuehM9vjo8cLn/hrRxBdvPGuBK
8/k3sosfq5cDY2B1NQKJ0kqagGiy805Nv0/Pv+UnBKQy0dEzcroZ4M0WOjtTgeiJVikrOdnP9fI6
MvzbTwqxGabF8nn8lSB0p2h4y8KIF0i2mTFIPgnXvEgah/CN9u67XkZJQjdBV5N2FAI0rlw7wehL
wcebmJpBYPNvqqyTN7JwtaaXkVooYPuM9uqv/FpRPVkBi1ZWtNp+ptNKTiLJK6R2tEtbEnrtDDMm
H2kbY99nbKEDUPIvatr7BgB0YhK4RflM77rZKr7tLdNbKV/Z6GC9a4pZKHgYsDD0Co3wcvHW5sEW
VTbPQxCZ+ft6k4NEhrVQnrPPYO2AnK0QWatiJR+nXsoy+UmdRYvkR4VottOtq0BkfoprHW+LORY0
J0gtAYiK+OJiyK3b2T/4/7IHC50RNJwmA/797Qj7nbgEeMyr8iY8/LdSnK5yoosffbU5VYHSVEdI
Yg4oJg5deNp+c/7l1yEWfviJII3u8W5HtKthOggpzzl/TBVByeUqVAqF39Mahi8V4ZjOSPiSL9is
9u6+eC1n/EBOpe++Ba5gwg4WZPjHVQUQ6K73CoSuzP8XZzGfM5azsTfL3JSc05Q57lUkkyQNUQen
kGrzNxzk+PWBLXdmm2xUNROdrkcllW3YoA3UHKtHS6VnrGPv3fTKTSsbX/a/+KcISjCiYArB4slO
Zqos120eQWhtlNi7Lzsf+HK0Be3RvlLUrhZXJq7eSgAJC8I0mrlKmc0NwdN59l1/Ds4CxrkOKey2
fuBM/ZjBTQMiocUAhRCScA+WVJieibYFqnDwG40H0kd+1uVZi4s0Uoajd7MZPNKYRGdnTdKQMA1q
ZIsqxwFwmGUTUQFE8ND9Q3piBONpWLFjmDY5VIAmNFJoBPg4d7keCx80vKjC36e5k5zlylgu4qKZ
SLLwrmfYKUqrLIzeTm4Hu5d6cgYF3P8eooI42/tbxfGhKvUuIGlVBeY5Hhh5yUdBiU1AK7pioXqd
AEjEcGjBz+8xGKahknXx/dyDCsVTU1/DXWVcsHCaIMHfLi9ND/V9aF423WBg0DZuhMRwN4SlEER/
V5R2WhgApSeF5EVT3cdy19B383PQEydp2uzNNOwZ8PsxhrxmNs8SVxBjsEeD0yUJtI/Wr0KiS/D7
9NYa6L4tm1o+9Psb7zesg+2KECexWs/JbjtIICKNr/97hOLHoyxEfQd5FGyDtx6wp0zlJ0ntpgvi
HOhJJipnIaebmj5FGm4VvAMiv/CKBbNZKq/qgHrqVJ7XPz3qGxqhCqoMhLSDRomCoxObQjDgFD/Z
KZ1Jc053o9eKJ2LaR+zbUzjKUPeiduo84o0/fzkeMvNwEcZaYhWoTXUX2cJYgNMjBKR3/HctKuzp
49zappMxTYGRLr1111nZu0koX41X/zjParfis7A8zW85Q5Ks24omyA07telPvME0yb42z6w4FV3Y
SYj9SR/Btfur+4KC8BTCL8sqFhlZ7NWX4Q7RjA/mDq0aruLULA7Z83AmpOz3m5DTjr0iwbE5syT/
ctCDI65LoibvUXwjS3tOvp1hB/4hKG04CawtZru55hiVgwIm7H+o2rxJmUjALMOVfXZkhZGdTytN
o3eyC2ZF0SxwTddFDTP94yMUZX05ZnFkH0qf74Trxf04bmuFuGJDBkVfiVly4LVq0pWLT0kSxYsz
EWeeoOK0cFTz6q/2wjtVGG0Y8mKV3lztb8+DKkpYhVJcjpBx7Qkv9kka2rDshoKjxGV9er/duho3
0nv0OeTeyidxN4Vr+xoPQvWkQDyCGOJoQxGfe56POwLq4F4lXJTDrmnIZPqxzozV7QSglzjHe184
GTlsqYMZRG7eL/n2Aj/H2SARFf+azKFlGtVkECacibxBw6cLXfhuINEigodYZ8xWMsDHoHyZVpY6
/VN6Fzfj/kD6nC1SwbTjO/xeDgEk3BWIAGfoOmG3GvMnOTS6rhcfg0UWwb7oTPLcCrkbkDgN9H1H
O90ZW5u1ZFnlECMoJMMjB+vPn91HyzoUZLeg/K96gtLe0w5DxMt5xslDxIoA58H4LVBOJYR5JYdi
Yw/LOuGEW3+P6x6KOKyEAQq2pDU+KpsFvImT78z5jF9U9sqS0BmBkUEoRjKxB4w3EwajOUxhjRVH
ZBYyFJhjtdieV8d1XBXlAJyw1rMltSkAIHg8s+GdRUKwXmPI7vmM29XJWa41yMS6dGsL/scv+PJ5
OfH/OkJQAz6FKNHG+ccXq6N8ZvCgW6PQB6NwdwdnU/iY6iq6eFCDamF0oNYgHZZ6O7p8pIzmnheQ
oQPGKZCQj/yYMNwj61OBmRa+LtyE+Q7XAxp0abwRwO8ba0OeLrmSE2T6zga3sVg=
`protect end_protected

