

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
R/f6FeJ0QLro/ha58bTY8NKxDKKO+q15gtVmuO+X1HoPKFvrmCJfIKY2+7Y4Wuzatwd/djCDDzbj
Lz/cs4hVvg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lvJVFxu1g3pXdpkq1DD/m9B6mZRZl1z25RnVPa2Pqa1r9owDEtgzfIY4YDwmNQWPtDZsGSa+gEVc
uqLBz0NWoe/TiDsviZj2qMM4pCFiMScHidDdqY7hiOFolMJLOulI7mQ0fiA5T+heXQGYdREM/Qxj
GFB/xJTL+k8zIvuECHc=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
a5PKA7Wq+G9niejwJOtSNs4IYuZHc8JqbN6w2EefAaPj+yqsVOpcNJaAPUuj6cFCMp7VN9w85Z05
FkFSxCcUs7RmQu3uWLGNQezUuGW/d6OS7GYPf4MRX9mK7q0fMkS51Hl+4n0QkyxOcB8Z84+JB4dc
KwKO49DHwZGhr+GGEZQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Jcb8JNchDQSiulaqmbTXpOUYbMkdd6d293bW8sxozNV2U0p6APpmuBEA/7+1IWt2cownZDUiOKbh
vpwDhXEdV3JarZHTGsXiIAWpt1Vb8QcOd4sKL7UeP47aQzH/7PSfm+5VaJ53FRa9Re0Yyiy+xiDq
5WVXsB9CYYUn/nWLUbEWGdBizGZnmhwxGfWdJHz5tlSnRgJn1ZXc9UpXaugB8C9Yfndn1hGYi2LE
tSAxdQ3IeR2usZtM/poSve0h0ybGzEZxjlKK0JJwlaNPwKJMIqwSNyeYlhN7d22YGRW4es59Wp2f
gGsqis3PqJ7NiPAfwd+Yjbzi7svUdzwMx+pfWA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JtZntbd26RdNOdSV6FB7P8Axt3WOPCRpCpwgQKzPy2bHyy1xOosVNfEGfOCxVQ1nZWYD5L94l8eL
17GOiNRzQ89J9xdECYcyMVwbwDQV1nQpWX+6FTvcVdecK+hQyFs+2Yn5HH/kbbObpoIJz9gCxUmF
BH71W4+J+zEZKiu9xnknefZOhniAzDyKNKc9y3UI0pUoJmpv4HVR3XBXMkvPo+wnxzA3wtzrZnpl
ABbEwNwHOUX4HT6JHiiyy8C6BQBDHp/2srtR9XQdv04gJ1JjPTHdrdHy/7xZ4ufKW1UJ666d1b2L
SBegWiCzIFgbSKTujiY2Ob2b6lsDW+W+JjzIzQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
U7NH9yg0f8tUSSiMzO2ZV0vdPTPVgwBRvvyiarSitGa0/REvP3ado3WY4HYt7rtUt6whHqYlgSz4
hK41g8yCOnMvqeHIQnhbMDDd1y7QyRgOUBuZB71vrBBw871SocSq9FNklLclETG0J7Khywsw8So0
HUBpgiZ9bVTO8LU+2SabnPD3ChIt7NLLDHs9/z7JnEqXPf7KiCTdIFM8Szq2mSAw2Q6DTv+cYfYJ
HRazXb4a76QvTIBZbtKXyaOLgRURM4WFVAPBZp/T6h91uV2D4iz5NecaV46d2ZFMpc/6K5y/I4l1
GU+vKtfSH1upfbz5itvG/2sn98hh9hrtmMHXNQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 67920)
`protect data_block
aGLadNnciJfkY9UvX43UAb/CgVzdgFGk5ksst1SyYhmGeeWnyUWRvEESL9pZtOL/YOWM/843Qfu9
c7Cz6GEL5vJGIdIDTi4NlpH5TtRtnlDcEgnb5h7l+tIDTNEOo2thHVrh7QmsEciqpf2YMIAhg/Yp
zqRdegztK5kKRrYzrhnaAFdpUqpY/yECgFVoFFxtfutyWXYQ6+kDw+2xULtXCsUOdH48YKy6Ryao
9Gp4ZBYR1NbFAkygUx288UVXkvwI4kXLyEeqZxm+sySP1cIhBPZq0AaqcGx3k0sfjiy2GGIRbjdi
dT1tzSjp5QS55iKs1QU0HoCAEbV3BiXsxKFRtGwhpxBVdVWRY1o+QtQkVLfAijLMGDS+mXEYMDqX
ww0luyL365Kogjhjp1FK+KhQgWJp4iL192ZEJyFbpP3p6AhcpQpk0rETvvRPU/12LHSHwOHMJ+de
Tahcg1+jYZCATP0uj3yFq2Zn3/E5kudlZljPj0pko4gDOajE18TjZnjSPM5DRmPhVTtzskbCvirY
y6G+Y6C9VmD6nxZCnJ6LgtxMAZw30sdY1KMz9XtlOqLVjZ4cMtSloN93zpD8z2z/1bps9lpic2+4
/fZ+zKtmo9rI3vTUG4lA+8hE4bpW0N+tSCkBVRmOvBiG1kBoQlUK1deE1cXIjR0lz/ach0S/ufJ0
gghOPFpqu6ZBZCKPNmJNtqIfCmhKhbr7s5rRCPA+t+TLJQ3i95xG4ARSkxUOX8WXyx8NjVCTohgd
RRfwFlr800fNSk/fReLgNGdlDMZ2oMoT6veYhhKBqs+ikP+AKkIQi6XiDqbywekT+pHlUhKAnkWE
WREG4KELrwnbr+qcgsRkKcbu+HDiYvjDPCeBuHQhWN/0NoJBem8LdvHAX8yZm84B1LYS4obQXcz8
SL5aQXBEPytHWQ4n8e4nw61o8MtXtvVZwBquHvzWCbyx8Es4U8PV/GCJb4z4XNBvas+RJFghpucg
RUNu0LTV/w0wxguidOJ+ORtUqccHL83Jzth+RfBIZ4uZdVAq/7o93uGKwOAxk1ylTkyk1JCzxs8a
fyBKkCndF/sudEeJ83WAbaFeiAM7GsspHeuetsOUXXgkBYP9vPPKTE48wg4vOMmAXh0yWXW2ahow
NGnNt63pZYxqAa9fMTKyJ2z8eMFMPe2nNE0cFSlCvk0xFrCBVteLf8LIlwF9vvzSTmqq3kIBXyyZ
JnT2743P+qjQHaYd84V/c83awCME4QGbFcaRWbBY2viHsdNr0D/LYSVGvfXUH8Z6wC4V8NdGO3Dj
Y9eYmTbHR24LRPmYJWBTFJeXhryOnEdyRVtqxzJODUeg4JPKNavUAjmFziCkgvmvEtIqtUxAt5Pd
nWm7WkW82YGrZ7EmQrXAjwfp+qGZzXZCKXeKQsNCeV89tb0AaHfD1wKOFkNVE4mBS1V1Bij0bqx7
VedvyThIQvPoMWhhufmfDkRlRnA4Bll3WdUYHA9A0whQKysq8ZxZmyWFwtTTpqki7u9oV8TfK8qL
xrkRS+Yy5OdeXMOGSZdIVqPDH+DposgXU/3enf/YbXDPujwgdYnYO0HyP/yCc7oDBCIqX0wgGadp
QRIxavdSSq4rJ5gSwguESE9O6Ko+2EyTqnlgsteWCqvBXOVbsbCvjC0q+UiSrOlFR8jQ1azc1BYX
PzDS4x6P1Kg6Et61wO+3IcV5i1yapLvQKDa9ZUE2pEtSWrRooeZe4Z7GyePQqAcS/px8NshHaOcl
gEAjApOGoH0m70t37qnGbVrxw89jnPx1lm7wTMk4ld1pZCm7duJdaTjqRAIWjPCNNBM1iQlMjHQN
1OX47HPm5Hneig2nrVDYpyfrOgIM8f4ed1gCCZDMCf3gLHodChTWkFuN8Hxl63CHw8YVSIZAAbUs
bmGqHP5f4GnVperK10xuvL/Rg0sC2R1baEZfMKwutxupSyESZiL45P7ltBec5blWSWVzR5Wpx0Zu
z/4mEwmaqAMLg9QabEm+MmoNi1PDRiILKpQLr8di5UyUm09wHqBEqLyQlCBGIflrltYsRRqOnZ9A
r14nofHYTWnfjgjTAhrrFqM5nSzMMQ0sZ2j3jWX3tyPMFwnCRAixak4csH0m9myQflWzjvn8iHpX
7eiF1T0QDLxjK1xifTbfml4+CdhUvZ8pHhnhRZJNX2U7lB+HABi6f83BDPhbMGNwg3IyX5wkDzoO
AmPPE+vFVHsgsp3+IN+N55+BW7trK4StnyaEakzj1Jxq1L2m//V8QMbf2uV1uqdMRm2vzOuA5N3A
96ri9f79EmEc801uL9oiMLwypdW1dQPHAE1YAsL+frp3djeGV5suvwAyi/1sE8UcSmwvEOFlg9xh
57hNJuKKwfN+0+RfNPwsdzcrK27bwr8WV9C/7xVI8X3GDEIUV7ffHCPfkWvdv4pnOCbWiIjmiZ1z
GOJWtYYgUiD3zRgfSW45/5l4KZJB3QA1Qit3RbYme77ClnWK1MTQDjaPHScbnPA5rvW3ZIBkvbQ+
KKAp5/sXqLR1cmhmV0ZhmIRJ6u5p5md/48FwKt3JQHhN8LsH3q0J6BAVlqkEoqIuYITS1oLgVC1n
PT1Vlni+PZZ8L+aFe1Fb584nkCD+IyfAthouqibtpm6u18T9fQgrm1QhuO+lj2nzHe6wm2A4u3xo
Dh1H02kjl0ecMGvbzADeckzXTPti00f9AsFPyWrqytgXaQeSb2hWCW/rUs0u1zLM8mBv49WVs5DZ
NznZrjQVzE5HN/FPpy3bqtelCK08eo40CYqOvS5Qf3Zn69VuDbqWXTaYppTSqTO2EOW/b81P+M3d
8WAzQK+TUWS8V3AG9aMEQQXHDU1+e4TNr/2g4yrtzjDNHoLR6UBMzVBNhvDRT9LZpmMMVIA/zfyC
kxIMbe0wgZMWnJB88VXSuSTciueDdgv0StWTFC/27p4WveMM3RvDzgbPvBcFMbwlQfS00EBbNX2k
HQ8dK9KIXUPTsWfdMdr3LyygJCxPnrrMwAV4jX6L6Ev2oJnV968Ozv68sIRPp0lwI9/z3vu0rNL4
9dMc3Vf35j+BN7Qkrdek8U7VpnNcluAv48uSFOCmq2kUTr727ybQFLcLKtndZmPJmYJqyMtPSo2G
mEfAVwm5iS8V7YQOWCrR9wVpnrlHLeLcjYwa1+J7oVwYWE/GMjH31MBnpTvXAr4rQL/BjksIiiqh
z110osRWoCoO0Tn+X++gDcgPrWq/qTTE4TP7G5TNdHBDYCMHE0BSLMQyod6SeEnkgjfbT8qTGq0A
Bk1hcxcqGeJrYzOKvkpdeecTUrOjvTd6iRTjlv6df6n24ua7yagY6UGWzx8nAhFug0xF6FV5Az+n
vYJK0MORX+izwPdPOVVgu9/qy+zWrVtGy5/w2qoRQISqd0/XNH/7d5g/Y1BcOgaqIBapbC3itx8m
jESQjsPaaxVkNXhyaM7F1CCCOZ2DsutaMPOVqFkTLku5RsPu4UwnY68k1BbSwf3Ldw+shfXFggO9
c5/sqHFD4bhyI+1zGvs6vd1XgfyyxC8IrO8i1gVT/yPJhFsIwhrYAlvFeg95rH4M++lRL8JjPOtp
PitzjPX9EpGLjxkasjojl1eI1HoKOsareSW+irs1esO4njT/NioxU4nt6h1LMV0Dg5qVA71L95/j
3A/CcwROZt1bxAmwG5Ktv6MRDkGsDQVqzLzc/u57MJo3xhfztFRdvz7OiW3DSmAa2Vvhf6wiOzF7
jQTltWFx+kY5Ybh5vQu4PbfMJPF2TattpVE+lrZDVQJ6G7ltXYrkp7GEXasTzsIo+BtOtwhHtP0X
/fBUzt6W22a8/nB4bhPjbo7biT7fyxWxLae6WDHSzhHqsVBgnxE7K/dv4hXmMdiimfBw0g+8rKny
u58ktjg1EGzPiscIYAhlNHt11FerkLEBaVMPZnwumX/a6xD8b0gnV5AM4BKfRhoFThweExoIsWQZ
ghIlkn+AHe/kp/cI1FsZFv/EKq1Cwv3uxJ1IVvFUT1inrMlgHeb6hrlzLnpbHHZAa+SXwBcU20lj
K5XuE2hM5dAy2fryFs0/ASE86+zBVUAZUhbZ+AWLyq9OYleMGy10iQehioZu/xijKa0rs8doKsUA
U3ydBWDP98lXA/oLjj9W/ZfTxRbc4wsGJO3Fd+EuTGIbJsA00VQr8B0kUlalGaTHW1imXUCbjmKc
EeNkY7HsitW/OhVR5s1EimglR/6+VV3wS8YYd+kUnrnt2E77pZXIMwK0naKV9dbkHfPisgqLCSbm
XzIZaj8OrDDMgELSG5w8wNCSG/IBJjLDytxyMblQLEG+paDzaTi0svUZ/l6aS/D+UmsoZRMEJ/SG
aCTusrpGHQ38bB7fkVyMfLAqR4vKnNcue83uYk+F4hVRfUUUqgGlW15zt51NtCTZZ279syPKW79a
yMd+7krRJhMFacXFHx6uLzIdBclsNU21UrwDkNBP1ZwJUwTtoXDW8NNIrA+QX3FGaSktlCTwinc4
uD0wIlOjY1T+tSHBEkODkzS5MrVGpZl2/Pg6tCiSqC0A//2f3iPkrvZcW49mmt7t/znGXeCjXDHZ
14jZ7yg1ueOmNLlukAaNbiSPAlLwzhZNd8MosjbwKJLjmgeLamKUwr8mZDPfRuwkhqkZs31mlJM5
EVYGY2CAiILiTr/6WbRNn83ea8jlgUrjzLWT0fFykVv0pVO6tzyEeOVIURTmbMaL4FwY2CpojYu3
Pgov7m+nNMomCfhErReLhtEQ9JeYyuZVpuuu38KSaL2BKyTcFrztFSpHINQMgNGo9T8lzzNG+341
BxCD9TZkbBaAUXUNY/QRR1R1+/OtxElnb5jLJsyDleSq6zSC4dcK8BA3BrHUvXZE6e4/Yo5WtqCI
lbRu7KRTJtRVvb6tFGb/G4sOkTloYUChRBFfzGXy1K672EEdKxHkSiIRGXWhDsmbBDvw8P0dYB7M
YZp0pMk6mEueoCKfxwzax+Tzr3uplghILXTGCNOc5nmzoZQRN/Od7gJdrRF+GBtI5ehUz35i1FNL
9pJ5F3j0ahgQADN6PySH1hmchKklQStVHcYKe9j94pf2w8Y/eB1G0SseCjSXwixq6lfpaetVvhWy
3p22mjYztJc5zHNDTMZ0m8LrmxHF74AKXUDBHDXTSMnqGl/bi1+7DULDvcsRp4XxQ7y/A54o7jUj
RiN+7mha1XKuKs6tJWh+GfW+NP9sl3mnMyrH71RKHMwYdzc9wpFGp70UmXP9PYQ6+IaYJ36Qq1mT
S+K7hxX5nbDynB/rQ9tXsasZV45npLcRQhuPgb4ddvj7cBQw3H9ohR7l3ZwtzaoIGop640ZK+M6O
uszUk6Nl7Ph+nDITJG2jpT12pvDG5VkbeujVUbnilN5Fw8Db6oWwV8PYo/alRP/a2EozVJG26CBv
difkdB2fqHieYFBVvpPUqGFXLyNo3donphk104MZeV+Dipq2mszFBKgQwKXWYlyYWm/7yne/mTBx
4xCkAWZzd+ZVMfezfOyBBl8NCLtvgOnnrBuACoCqDqJOhERQIuL5egdWm1q+6Tb4tWTJBP0FEVp7
nwn2A8p1obCvPsyjlRKLHDoFwHLKKIbqJuY1gt169YD+DVLwICzOM1i7hgrGd7/OouyqObIxOIrm
stCedQuSUFa47dldtp6z/v6HfBTLeaoSP6AwkZg92u7LvfU+sFDoI+Pbqi65Cz4FYmhDJmlxES0y
gRW0JOfI/anUR41q5azJk9ga/Tac/j5p9sbOTfHMSdgLxhZA7dzO/kXyenfd+O4KuYihzxLkwXFU
A57/9dAUXp+HGTzqzNl7tA73sspWne1opNmvEH/O2kOgynyAgflVoRoEfuaWq7ymsBTPrDoQHBqb
NR357eaT9rdWRO5QP3pVUHVO8sWRSmFTy1HEyd9CbsB6PZ4sM6baoWwkQ5EIbo4fam9VHTygSDv6
meJsC7fncM4BY0x9iF/ifb/La+2WEbvmWIZkKEw9iCfQ8pBn+v/yjGyKsvWfaPLhY2bdAZHLlcW1
KXjPNDOYQzHZwy4gVLK9XACnYQ5/VkkkIO8A4BFa7Xhr2R+L8aWft24kCYU1UoaIiJaIrwiFB5+h
3XoeR+zbKW4RjLREeGVO9d9EudzsbPi63Ug6r1zawIZ64AGpSvF0kOBycRDJiE2bWaTOCieDl4Iw
e3ar5qpwCD0pl43+7hyX/RkKNxpTDyv7OvGfxbb+XlTCTaxo9jX+6cUbFvJwK0KT6Ykgu2dezZU2
rgoo3pzE7LqZdhJK50mQk+uHWyz0wEgpI5oT/f4o8SQuHU+kj1+nAM86A368Vpx+UVDAzFVCymih
Bn8sXHknj3uqCLLNhBj6QaeKVN9Gf6gzIX00zcP6gCBNwa10yarmQmMh1+HHdj/o1inwk9IXk1nf
WfzeJEsgzkS4rsqIOXsdPV5KH2v2apc6Nm53Wh/PE8ugulYI/jYNNVyFoWueVqpYXeWZPHMnEUDy
trrQ7dQsOM8Z8OFzZX7YSCgqUKlmobj7DpQBo8JkZkM6yxzsSX6arWowwtLiPDdWzzSAn1Rb4Mpt
LTnzEdmmuX2spmFO2xDPJVRLNbRHjRQORRzhcZJrQMhPd9xbJhnQ1DgWIm88k+3MScgzUXEeAYAh
fMEO0FzEG1UsgL7gCdqcwoA6cSifAupxMCHbWBd2mZouXv7Os+Q+YSK6mE6UrUHncPluA4KRUeqQ
+XVV4yMSnWlAQX+FY1jw7pnG3oXST0j5nidaa5Mmhb4Jky5TrovXpvrsyR1aR38iyj6C6jz+hZYK
X2F6/HrZAWOLfuKTCNYFCALnCLF153Y33K+hP+HUBRxhcIC3aqz35HiMAOMxzw9o9g9neuXLCc6V
DVoTbxWFeUMTOfNT7G98Qlhiem3ALg1Bz8vlbfwlIBv8M42MtmC6gaUyPt1GKQxnUb+AB9z8rr9k
PTSR9usjiTFCdbXo7Lr4IkYtmEWhQdxrHDws2ilT8Z+ikrHvhdD8b55CyotIcgqc2xDTOuIFLNZ6
Y5DUafVgJBFhv6tjmHFPYIFj5vdTCK2dNrZ7dUsLAB6ITbREWAacQEUtsDRsTfE9Hx4SmJ8QqcTP
TMm5Djm4Kdgkux/3nZzOv8v1+PQRRm8/EhEBW4PwIjkYXpAGzdyUaRh1roP3T9FkGUuMAZl7tLP8
cICJ2TditehmpAKFg/15cl27QTVji8QIDIZCpFcA7kS/ZNiboplesbscs+3ogDvX3DAUr4LPP8pA
y4TQj/q/d1N+mzMt6Jqhgo7+ebP+J93ArXL1dqJ1/OtBEwJgjGFDa8kGtwFvcFxRBInfCbuUu+Hu
GzpNPuUY73AlQDFQ/x8cphL+SzL6fUxxSuOun8w+sH/BqYjh1Zn3KRlRxlu+qfc2ECCrIFzbcNpM
xu8fKTFmGO5oH3IFQnDAALuLRSh4ElJs5hKG6Wn8yiXPRtKwzLx4cWaD0vrLRpMueBjvBEfl2hDM
YDVlC72F2ZBSXTBtrK9Df9mF86l2sadw+cdlOuYNDjnBWxVbnTl8sZ/S1D06qPa0jHXcMtNG7KRk
7OI2HLhG3WSqP0QFf4fenolI6tIzNPQ1MfWh93hpkQCukF9wEsOmVcdgvwmx3ETS/4h6g5g0zA/f
jKdO+nw3ZTPi9rak3gtk/8SRPjQXUCc0S0l3R16EpXuMcCIouS3CmAn6qmcgOw6ReL82c+EO+u79
hNLaHp4nxdFid5Zhgx0P17zEK4qCfdnWU79fMbClZkC/yQ5rWBlxumIS8N5UZXyvUh0HpcV2N8pr
ZafejUC/kEtOGKMFUJSeu0vOKnkpsctzBTXtQ1RWle5SYYmG7ysImp9Hx2hNOWi65yvnMBUQLqco
2AanhZ7oBOkcLa7bjGh0syjBGcLXDtq7TuAHV92mZo5RnnyBr29LcSsT5G3fHDi1MNsmlqIP7upJ
mgYRhRgkcTjwsq0kziNP6sZpRCTxB60IrKdTnD8Gq2rX4Er4aUKrWeOnp4n3NwyL4DrvsaW5xEK7
dCs6De+JxvWNFFhWUPNosVNR44DOC1Ei/Lr361xrtQiSvmSWY8OYfYpiZqrmWzMaw4nOg29RTqQd
CtQFVfmvifIwgkk4I0i7sL4TTnbaFNZngjKxotZ3Ne9Wmj6rmU0rZcOaC13AxutArlBdFnb9JD1G
yAdSSyo4tDzEUmOo10ET+rHZJlHKCdMtxdsr3huB5pSbbT2f0zxQlL57Rqy6swVwQ1RzX43Fx8/L
XYdsaXs4lffduId4vN7S98zW+uA5qZXDIXtLtfI8Htkf+c4M++BEzOKodZ5nBblo/WA7OI+BNQX6
3PlBBQG7/Pp9/hq9NYazZ6WhN+hvD/LTjtjG9/U8QDlL4eNRQRHJwk2FqibLUPVNY5kMdax7vdSx
HEKRytLB+KslySBO9FmC9lbpmFK+6O8+8eX5NW7RlQjyOWb/R65FSf7Yb66OZSofonc0O4VZpZhQ
4WD3RaD9Aiq265McmDUvY5f+u7kT1x64dkoBj9OHpDDZpvM4hFCxW5IFx/BOsRIEFqPeJsB5ppx2
j+Z0ehFXlY4c6+1V8+YDc9cLHuTdDV4yk0RdMg9K2czmHyusFPlfLI3xD6MY+Kyks+ZIwGKMLhSu
846YRcKjg8UC8iJ07sCZSlf8YehwVOwKA7ltmkCAtzPkUUk7WRgHVyF2IVE4IsjV5hG6KNfRZM/1
zCminPKfHBI5VzNNgQYNBQH7DZ4ELTtjmiZP05Hl9k3yANU3f8qeO4pWntGsKU56/XCz4ejW+Rqs
dSyMi/wzHE7OvbQ2A3T/7DTGTY2tUD+09Ns0eRxEtnoR8S/Xah0/VHAiLXzyEYU/3YwttJZYci/W
GSBYryPgCkGgwhp+8CJZtvmV8ls1FuY3ZMmLtvv/FTU8aB73hs8d/bysdymfA6LyotZRX9+h1Oc+
JpVuzk22Nbr26I1ZtAjvPX/S6GWTfJcAFmN0ncEJOuojzIfbgDLy3KDL0CtDH576kh+UBjoYSyf2
M4nm/jAp61wZEYwZpq1baGQbmZm1+OpGb15oWxB4UtkER9P0mP65qijAa7KBHuV2ptTEEDXcAyae
8a64RCprkVolDM7pRAoBd2rgI+YxDfZ6/RBRVJgOnJuO1a8IhqzkIKBNme0JcoFtDf7EBU+HAEQe
Ubcql4uL9Em98LbEymSuPCQHnH75ZrnKb533e5BqM+FSi7QP/ka4whAx67UoVDWqqDy60h/BCKnZ
VO/WpI1kuHp360SVbITw8MGCGS0ItWmKb0Eq+qUSwQtm5MO+OqJXmPGa2t2z0dENEA/hi56htI3U
BWiLB9zjpVRdpLy2lloKqBCW580Pc8o3KvXHcHqj2sHQ+oxdXz9KrFU3zjkx9DwIuN+JfATE5MRO
egcUguvgb9YcqgfAGP+tNcBgo//y9l8dbPc6e7zDH5flFiqWf35P6rQYB2p8/xAcoZ585qCjnFak
C82/cqEcqNcQbC+pEd7lsgG0zw15Q7Q5E8dL4Csjy17akUNdnXpbjpLYJVCdLtMk7fEdOtOlDWVI
VkCfSe6fyWZQ4KCR7bDFonmJFFgk2LasHQTMSvuM2oUN54fvdP732WqM9CZHSoHTgN+jfTBVl1c1
h92Hbf35iNa6JMyiTGvWri5mPKBz40Rx8+I0GxN9h89cDrLqcUlD1pP6REmUxPdL7GcNFrXugYR1
PTKBHO2b43flrarjtEpjlMSJ6lP6Ifz9VgoyWXgY9eFa7/QjyRd73kXFIo0e64A3Y5EyB0wUTsaA
1oOQnxVYMFVYO8YLvjkaKMJwYsMCpPT/qGjJ+2Hz3YQhDIUJuSWSqHwx3wdj9uio36yFyNTiq0G9
kPimiq5QWEnIq85CabBrzHFe3jIypUL8TwBatITu9WJ74oa5RPj0gwc92TAEV7H31CTzAGunXN6+
N36MKuIlTjoIqyYLPiH21yf/VOFtKXywwh+bfXFl1VrQdMUNCF0K/vOBPxGQBMhT00Su9/u6X+H1
5PHDObfx0ZXEj4Otz6HyC8V/tO1nWvq3vBWDcdg6EXo34+oHT5EoIrST7NhrxPzWFZbSR/Vjb6dr
09L+tgvhZjLkDoZZdthXv5eTvY5Hl4PWRO3cnsWYqlPSNM3xmicuBeGuz3pFo4zIS9JO08vXSYev
+3WroEFn1az6eT9ZEgeSfABmFbB8mqsjlQ4XpbotTG04zvEpHUJI5fnJpRPsNu64XZ8Zr9qfrp9S
M8uSDuqoz39m4b942z5JHi1CbzINM1rqVnR/9WIZE2wVw0kOYDdiZUTfp7zppxel0Mrp69lGmOcI
fXtWUoZaHjt4lKRIoCZ9VA5PN6fA+Ml7AFivXNNK+gJ1uQoPQHOpoXx/BeWt+E2SvRDfP6+A/Je/
lGkA2sw9NuYFbOf/wb7Qf6wWNkiQ5iGNixYZXzJkh2JH8k+EzbWQDOySaIggil0yDoJdEh1dSH+r
fM7GsedxJ+7nOCrK/BXUOjYaFe6Jp82neDgiuM86/i7Ux/wELpl10lieOGtyolfdNwm+goN/c9S9
tt3LR+LBdJeDfX1plcPfCkvS7e6h/szkWd6efnH3t/clAxwe78SM1IGmTsRnCkFTlnVKD9o4E0LB
4fM9yzVvZ5gRTCvaGmQoRJ6Ne0tQnLin1TobhqOonX8pVBc2xVw7dTEcZTgqg2Qmih+zuVSlrV7p
gn4HjMmXu2pQgjEmMQH3l7i+EkW3M0lK3m8UIb1ghoVuWvFoRWZofYe8JPOO0RemE/KsYaiifzzh
Lr9JBOARTc3Og0+jcsT3Rm7Whw9QLfOM4ocQjaSzmlPNLMzDk440my6k+s4wFidM6yOdXQ8NSsoR
dJch5TmZWG9HTggVQdQ7xgxAQouUmOzeO0M7HQ5Efeig9gUe9CjoBIRMzHSUldxzG+5zE+pSCwG5
ES2XCwJIJnfvq984XxioPv0Em+x+66Ij5Y7e7mecIffMqSJaetrip7JbrJr86FAVM/eyamDEwk0p
kK6RfHhu7t9z/rbbAE1lWZk1ffXEgRLyn0LRuEDdo3pIzqG9rrZJ2gtXH/jj97aOMMgbj09J64ij
2+kIm0jOUpFipVMe1Ixi7URP6nnDempjI046RrquCkJoFBvRlMm8V6JDEgJOOSmFRhZmQLHA/NtL
pZSOEjqhiNSd9WIdmuLhP6JbXxh9KcfWGpUm+mAwi6yhUu35ojfXDQGZwIQPMQFmDTgaXdTbuKxi
DuMJNBt/QkPVr802I5t+7/WeOqku7/PCLk1n6rgawos3xVSfKuvqxqULhbvn7zrBJBjTqyRS3iF2
FAWSG0DfAfftOe0Gc99tAKXd+vTFLSOswIufM02ZquDEZIfCOFLWKqiyi3d21McxWuBSGFN/NA1f
OzK+2tU0ji3jwVfm4To5eN6S2dOQ+w5PucKoqZuPFYU/dl2ZWJeopf0clqnnYRXI5TWlp2RWDApw
IRvnXtKWtBZuidgJnkGST748h9tBkbbi+tLEUcvZB+R10vpPY7ij9lN+VgJUe/bVcvcHieRInERt
WdYR/xOCYFNDi9P8esR/AezfKtVLuCEKXAK5/JNZuCtuKUPzmBSx2oX+fKrnfHpQsoq1fRsUeTfD
omn4J0namNeyoJKW/rq4nxCDJXB3DHtKpTQyVCNEwj9TdMPyTZGTK/X+ZHzjFIuFKlqM8RceTjX5
7XLVPWY4D5CalCX7doVwtoMpRYfxj0wXOv52cUWFJ+AZ++KPoEu8a863xJDNY7TcayQIoZoquAfz
LVwfFtHZcA2SE1xh5dBrBTdWvgty+8ZaC8Z2o29H1ewAUJz5RMqYVhRoMLl3Xen3TtfCNuaStu63
LxmC73GPSjNgAkm0hw+Aw0Tw1RsAzKKJ6myNQbWogG8xovf9oNIWL2kJj07FZ0lpiQc0EsGSvKXF
spBEWGGAiPym1kgq4dlKs42nUQRHkscT3IBwYVUPGeBz5eVcIRkWJ2mEWYTTKHl2CGcrqhm2PkXG
EXGFbZTtJA/P0B/VBiGZ2JpihWsI+sfApkhReiJY/NHAgZEzLKGtzyRFrG80b7/eeLKtleve9CjD
NPXSykt1edEniEVAPEP8tFW6OFQLYMjaQEpeTWSEnXOkdK1ntsHSizOnO14sBLOP8b+VcnXhEf/Y
0a/5a81uauYYELYq0ibfTudBGIJV3l7H7p/rDFKYFOWgWi/Gf9oz4qP1pKEtFNx4cpDGgbXA/Nwk
+5rhno7Agh6wwl0nzWsedip9I2KDRbUiE2RwqQ0fv6uMqQ8bxLYL85MOzl2TjRM9XJlbjcQElzS3
ydY+z+NPD7mzXGncV26ngfRyClUD0zqQC2Fa9fXfESxZ2A1IDoP7vKEI+9uvMZLNGvjf12FblOMF
EwLJCYgbo/FfJsOuQOiysk1HkjbS/aPAxKDyg/hVS7uqXnTxcBZ+I9kuoeE1YibkBxLDptpFL7Xz
hcksz+7Saae3655rNS7nGEh6+54cRc/Iim3DheO7J7To5rVzo3qN4WrtuS6fUHeBmoZV9e5ioKQD
Ogo6xiVex3NH1G083XqvvlYCGRir3xeBT54OXbSpwLOkQ9wRg3z4EsUnfpbogxzBpI6FUj+4w/RF
oMdWNtOMf1FCMx0lKW+1UOsvPrbN043PmjQQwVMv1ATuf0KjoyC27hmaNKDCQCZdCiiiq4cjH7Tn
pXybD1aYdg+agOKtVNE2v/TbAJUFwb95Po/COQN+elwolr6tiDQmBywifkHRJJWapBZdaTFTYeAA
bl8z6R/vMqc7s4g3kItHsk4rEWQCYzLhB1XbFrPzSfFzXToFa7BqVRaFmBYHLbT/05IrWghf04xc
o3Mg3/laba5rOTgoH+xbiGQxeH2GPJB6zX/xRLdQervG3uGGIGiEYOkp1BRMPKfbgApXX19jSQpd
i8kluCPL13ZJxPC76TXYXDYcPEF/5WTMgZ/2PsRugwubE+DDXGR0sSY8z4QBtzzEAr52pCgJiKlg
6xx650OVj8ec1232my/DSPBXYMW+M+wTsh1by6D8X6w9rxf4UeVc2/+AO2QC5KBzC8Se6tery74e
MzteBBF77uhC8nbb1ej0Z6kO4QBj0Y77VzCnWmKeGXhb2Ou3HcYpJolhY0sHohhg4UKhxcdD917Q
3FFDmwRjWikiEg637Grcyw38bVNFw/KQtDne5Q7OKGrS0nx84tHWPUp4wcR4esTlJRF0WHYsDZrx
+w5zN+ARFXXiaZznzqVzZw4u/sB/IvWs8xZySUTpm/APHaIzS+2v0c6MQI7t3XtKBf2z5p9cZoQR
OnaqQY0CNSdGhFJHjRmcDFUP9oi/gA979qHXDqhfbQvE3c/+wfhaI8hd6Mlm1v36ZA8Qry8f4pkH
ZKNvM9Xiv0PTWcNfKnXV5tsmqJcIZtq+c7RkqeCm32VHcpOrRyVSmdTmXkX9PRSaHPQ/hfpNLosH
5A+qPVWiarf7DXlMq+6r7yIV5vE7kuwF3eYLObJh5MgCkIzTh82faplK6/jPfsc9p89dwpjcn0se
EBzQqZUoSg0i7CjhNG8rXwbx6Lm/R52/6sYyeouSXhxKHjbrDMXfyaon/rXMvnq2jVS/I0GlHxzY
ll91mLJ9JbLhgDIr8Mu2XqHhFilxRhujak/aSBzgymYzKI00ly5Bmi3B550llqOpBgvJynjwdKzj
dbCKzpkiqecQP3lAnwuwuUI4ddyIbgzhl4l/C78jYX6HYV0sf25CgBlP7JzvdjYEFB1LrMUIw+94
nUow9rRV9Jg7wHGm4elfOEvBqNwSm81We1v/HmTpjtthXH6ty3UdZ2f2TjFA/rB43bQHz6FVZnSa
cn6E370XYueju4wDGNde5Siw9J9aG5i3ZWvGLCX8kWeaR4qcsXxFPo/qbdc9KRdh6PTbvdtnfxk4
1UfCVjp9bBEBbBBGaZFjBqmSG4xceIDhLNomCfmAanb4gs9NtfBhFUNRC8Gn5+jPg1XRvKrFRE24
QZUoxZSudM9Zf927CI8/3RaMOja2gu4s8SpEfNZ6YLuhX1Ig2+/Qt+necOmD6WBWrHdQEi68RLsL
8h5p5VwReEBdnegxQV0IrJmtsdmkcyxzZDdQQ7nu0V9BWS74v7RBtMEyNHHM95fTYEqU1AOeIwKf
h1p5cVPuBSwvMaNbsxAPIufsumz66bdxNUKDa1Jm7Gt/MTpmtmk9Yl3iWTRNIuJSJcAqF/ASmomZ
/m3XgCXYn8tYyOLc7+U6ZZtDKAwPKW5jrj8Jy6yL/VCpQmSZsPROCf2iuJWV3wWzfqlWl4hK/937
Gr/+O4DSfeRGeSGaqPSUH49irvCQ8q5pwX1gxpgEEXG6NdUf0naJd3aSjySJpjNngD0YdccCU0k8
kOhpa/nKduKd0tiGG6Bd75gcd1+Fehs42hbBQeRCzD1WI22TWvv3euMV6OJgxKkDE8rEGDqT5Ku2
jekkaoypTRhLXkJyklF70KWU0Dw3VA/ScXRXmY6Zj/RcwdL4OVDMCjWoMdMwNl8KJCZuBIB57LMD
TzC8XDLZSxhSYa4JfSusYPiIWS4z4KbyBd097OHxRfuPJGJ1uZ82RGmtEAeWeP7eJ1UKi8ahqR9q
0dRMMyxPqRLuHdafzfqa5xkqoXYCFxaBV/gjGSXb/pNejFiToU2CgGp5tqFqqxQ6///T2fKU89EC
YrVvIgZmkChDaMUtGmkdckzVp3I4mdqDSG1DzYMb6t3efjEOR1RiMf+XZk1F/c2ejUC+VDy0AH6t
9GOM48NDhMP1/+XfStQ2rQOy70T0yWNmjMI4fUqwIhYZFkVIuZZrx6J5ftIgjgRvfNK+QGK4FN1P
WqDCiVrnw90VdjMPRBRuFxwecUmI6t4L158GCiF3fyj9aI33da7mOsnWUvX3PTfl8KpYHD8wlepu
wF9Bwe0AH9TmZZ4NTGY5l0DG1eBr1pMOmSPAvjv2/zG0JgFEPV8ncuBEECvQLoEVRPd+5D2UKhIB
dYhMJfTd6O2c353WIgxLUqBA9E104LvPFPbWAnQ/AlYt5GSwhX4SSTxT392vJchDMmX6AOrxTXx7
4l+sFb52d/LgNACJ/c1+17/FyyffSr1c3TUtOyeDnxjPXfIwcihvnYo724Cj27Udy4BrUbz1ARqf
Vpyrr1UZrBqRlodNR+s5i71gWlYSjcNGGU6eqveAvCSMyNKTKSkvMhPbg8Edlb64J10zW9O68Xkc
TSdy1LAPPMz5lgv6Ds+KI0QuI1DmmDlxqXZIhiiY7dk0G4qo4h7MDzL67uMIXcN8eV8tT8jAB1/h
/oSrWHW910IrzUAmVl2tYMvKAj6ULUziFrTXZrTqQSq+i5CPTFpy2AP7cZejwQlY5Vb5ekBErH1b
40FB2KqUhNKviZWZAjzxgdMrpVLmWr+q50avi/CFc62Nf/lGlH5S+TqjnNI06lqkcJrUp8frc9Dl
0cb9AiJS6KTf40bx7ebzvA6ISA/iLSo2mkGkccLmOTLP0cXWLUmHphGrw44Xqjz/0gCJwcLKI/aW
WZAarg/vRoZPZ5pcshZLPdr3DfnAqkRTUE95BTlYp5cSNexf6jIvT/Y3UH9zgt+IDXPCmiQvh5cP
iDxHfihmmRRisco2cUKpZg86Dv6lt0+kv2TRhjLu8T3b/4nfRrryo+6EPIyEDygJBpMppVr8S4Te
4FgUzXsZwBdwt0bL35nWdLgOcE+Sw6P/vuwnz/c0LTtuj8uqA+JGzua1/O062afLu5b5lc4asFvV
WWobOnolkPR1lvLTGvfvkSjawK7SaRK/2pAQ/dXfK7feUKIPfP+jxOD0pklKiG3kiFl+CQwEqFvW
iI1bLA3scPPaE/V8JxMcSsUDCO0XIkETcXYlMOuU2clUgYrkeK2KrvVSTZPd+C9ViV/IG/ryELiD
esFja72jzzGIdfAz7D6AVh1UBhM0obSTQCVFguDHWCccjxm2SHTGFwltCdYtS3E5Bn3o5ZNBrjtx
qGZYKQygLtHDsSYKVxc5qwBY9+52lDuNBVkte97xhNPRgB1yALpHYxH7CELoBSV2YxrdN+VIxuDI
zmihgHzegwLtHO2DfrW0E//Eu/bxqeFh1+ZeqRVyd0gYu5RmbIa/J2Dbxl1QVHUXT/iCJISl3JFb
SnD7paRuJilQ1eUHFpPiWARv6iPFqI1yU2cEWybpg0SRaoGq1Or/N7jDj2kfQRghRsipCr7BvRzp
bdRty3ek8ypYAH4SxbiJGVmxHWHXL50pWYsiNFWBjildlPz+hv5tnRY1BiyzP7QfSN7pfezKO+Zh
nxBt9fs4du+n1K5DtPIHWVRbGFuwpdSNC5Ljkabyl9NTZT8G4om7QPgi8FERKQ+EW1Y5bUSHxjrK
5NLmB99RoRkUm4Q+18C19Lrkk19bhMcO8smeguY5xJhoSgOG6uVMaZbl0bmGIOvVMAzJ6QAp5kFd
yD1+D9kASIAXd2ysBY/Wku0Lo5MWX7mjb5ElcvTV7BPUj5yuZnNpvK6h5bcqUgnykNHZ8rAHVjyP
+RhK2DShvNhXNjuHAKQe8z/JjwU73721p8r1c7HuNTuClWMFFmDdVr6oFml19xmfp7pZLo+GTY4Y
+ps2Y75+RDjgAJXKV987e1LrjS5x2xgjGDA52uxiXBANTDR0WqJ7nA3uo7Hg/1p9eHSRbcaAkn9k
t8SrllVgy2oNbwSXxbr1hFcXuyerU0Dr16/fFOzTPiiyhijvF+n65AMqh5uMebBS0YRdtwENIDdr
0WyKz3PLMP8KcgRWgP3E8U/AOzsrcA1PoitWbPRbJjbPsKUcN8HGexhI+WhRalTmSGOfrOAu7cOf
DoEo1whQRaOmXyyPXuDtwqPSysqMsM6FZ5lWmiV9KDr9GlD26GhvAiSD/AT/p9OtfgRuCbhT4lRT
FdS8KbZ97Eu9s+irnMQM5DBMWNkifsIL9G+s3Fkm4HvEj8Q6qHfNgseLldNN6NG8f2ZB+hcVnMMS
hHNIkwNAo3okWSRO1RinDNO+1yBfw75eFke8I6mX2ctVcwRwbxhOradDDqy5EiVSqfH0jAfFRH6Q
e0zN5rlQEb/vpb+H0krCFweub6vNB8UFwQ816TETDNz4EtRHfoORO0iBa7EvrpOdt8pOo81KqDTs
PRxNz3ZeWKcfssc+VaEyplYldUvLU2F4QM3/avbhC6+GSyB0WAS8Tsa4D/VUsrP5Fbz5LWUPLb3w
yCKlJv6sxJ8y1ghJlKbKJwopDjCuDAM9BCPoyDKpKu8BXPe4RKzWrtzNjlFqaGMyw2j3w0JiaSb1
hYnbaTs2HN3ZqLWXg64hABy1jrCN7dXxetTUhHtpNw9tbwvIjhTOp4wzf5zX0XXBWYj5jnShx/2t
bqBd58mHuICsirmkgPcLxf9cfxrVihs3+iOeMy7HS5+pRJZf/a87K2HZjZ0nErZswtVKKLc10gLl
1mf9MVD8wudZcWQ3XUsoEgtCU3zbFdmUQ94dwxYCrjm2xEB71k1gZiOxNkWjs1LYlQ8M0kPhQPM+
Uu7/N2V4fQO4WuAX0UW/ewR4j/ojv7GyQ/oW1LyQUd3gC6zD4jjrpYCDWUuHRsD2C6kU20THvcn5
9htJOtaQ1Jbs7xa1yzGdLAFVQox3mDCdhBCQjOYQncgjhUYwrz48WRsV8Y2ftffpbaqN7/onCipo
641JGPv1UqjSWat7OEvhhmBMxQ/xx77F1G6QRXsw8iHDH4KhIi1uJlZG6GdBXNxACEBAHLDRtYH0
cYn3Bo7P3calJu7XK06b63/SoRal3eF8eUCrQEOPIDzG3ByEMQ9HXZNhy54nTg+rSPoE20t/uC35
Bj0NIJ5qhIsyJ++GNY8PiVqxPhCD6KiZujmqZLdDUAAN2hlF8DVmE1lh41qTVIshajezcCHmzZMO
4GmdSc/HRbTa4c9yK1+0cpoAhBNvSarFSWSyhpuMBeyYD3ztXyLP/HNHYzn19yy2Q+bqK9a1Qq82
AB6kseOrPRNJgg31Jy2mDpvIps3W0E7rQQwVPZzQHGJ4ev9CHDjlUIZOHZ2++ceMl83LnrFcynTl
Gm7qt9FnBuSD1xuPFGsQKf1VooFZ+Wj3pmyLmOcUbULo+FV1MV+KhR26m7Frxzc1Ylw3kCvattvT
B2CBi1WPudi477rUnbr37JtfoMLfXtWfKNY0CZKNJTKD20obXHZ0IMUs8ZSoly5YYldqArmVYxK/
3NPExObQHG/s0tjdQnkh/W6EeDL5Ti3W+Mgk+9swB4O96Jk4YxfGLWRYfugyu3tmK5beERivfur4
+oP9jxggA8Fz/xLl+4ZlYCjixMxVyQePrPsU+6bUg+tpMdhhOVm0LqmRQRT7T5cHlKQgGTPcoWb1
I13JUg7T1694RAmcGEGXnFR5/SsJgHa3c3F5cjPJMcqTxqVEFHd5KYcvpfz0yMBicv+CDRfJ1/sS
xlf3rP9+4lqyC2EXFxmX9bIisIZWy3mCp1Fk1LGe1NQuvbuHTGxE8Cvv6pYYvlxM0J93yjUUfoE2
vjv2sezNT6KnKewuW88RyzowjflvJ/NmGp6COuvvV0WX98PMCA/N2ufTQ0+rAfHYfA9Dz82V5qPc
goIY/lHIKIs/TBvNLtKWEbaKstpCEnRPkg9VzM5fZWi+hMo7ylJYC3a/QAZ9jg0MvxP/WzReJoud
JbzHxrzC6b3zbQxdOU+EAVulTuxvd48RPEhNxZratdn/TMF1OmF3QqGyu1/I8kPDg6SUjbh9Ch4G
IY9hiZ0kSM/+Uxtc1tfcj3OpKaTqZs3yp7YWtiB29aTXTIZtQ7Yj1F0Wak4h1A4IiCs+FfEt/56p
VG9nMsDoPqoIxjzAXyhz4Vi1+4TWJrxMAvnsUfczf9phKBYXJqsr1xfJX8lNrPWd11BOnQRcaRBM
DPvnx1EvthS2E9JyopDD8DIsoTNbxGn0+xWXzAs5scseUcod9gXkby/zqRqUizGtiW+aZN8sj20O
idReREYNZusCbQAG/53Z+JyqMlnNUCyylC2D+cy99U8f4KDdGGjlEe1zx2KB1dW3U1K5E+AbQFUU
Va22RbkEHCw18OvS3qFmsvicxX92TOka8B4MXnl/B2khHLdb7diiTBWcbp8ULYp15u75Clpeu+jE
bBTNPthbRJ7DQwsKRR6dTsS7/iKJgsUUMQungWvh64fYVPkxvM0JK9C4piciiz4VErGTqGxRgxXf
V7MjSWl4Oy8MBgA+OxofbFwTBOQmt2BZAl8TkAjoJSrD/zRK7WT8uHEMBUfyPOOoNtHnEy4HXwB+
QDfqVJpObh9woEiVVBt4RyGJ7Vn5nHFDOA0x7g2zqGpkepEEpadGC1I2+Mj6IxXEdqeGduZ81G/U
hzJs48xUOlbgZJNp+d353wHqwun+bzyZZTivUf2dJQvu3DNLd7dbp9tynq+TlxgcogZl/tDMVW1d
J/1dM1nI2LYgTJltc4bfE8mlJCuqAtlS1fE/kHH/hBUhBFGO+AcH1U7JMsvXJlOtQZeyAQ5EMtZ8
PNUdQ8+vjP99qSnodaBpsM8+EMYytdVKEGbjW+q4A+h6z0Wriww5mwp1glZcqkJjbC87r8mxgokt
qSE9jVnUsC7LfrpLtoV/Hh+F5unE3jzfcbmSIfsIx8vfxGHqAEvC4t7Yq/V/5ws5xc+U0D6eVI1R
XGjy9ucNAYsL7HXlNFfLtayWmZo3cYhRiPMioiT7s4DnakLIVV6n5uwKWKxrKNIRIaCYUzkaP15t
0tUysYkcFWcYpHzNrj8TCgkj+3ku7ko4h3CI7RHSwrjlsbnIsbEtWmViFWsMwIWPe+qSFX6VdsFx
geGxVh8BRxeb8ycceN5PC5Z72jj21dXj0QLJ1YEERUVFsHV5MQasXregmGpbH+faUSjZ01iyudUI
PmMCXxxpf6yQrv59XzltiSEMqaCAefrefcw6DVX5V6PW5owvlExhlR/UEE1lGZmIXzeYsEvJhwLJ
8jcoDWDAvfb3a9+DoIoNwPbHLPQI8asc+LLMKFSYpHF4UdLSzo8s4+nxdVd6rMKZmeWnKyiVZFhi
g9yp/cSwcgm7NeF3l+1/nmn0VXI6bjQfAOQvFvbE1dKH8ylR2M5iQvCWtLXaNN+3m2QinNKaqqzw
1DWaXKs4jXIITJYsrNKk12i/kJUy+LLStnsUcp6SxCr6eKO8CPZ2Pphp2c0+ZILR3ge6koCfpeZ8
1iC6xp9bFKwVhkNSZY7Jb7KOb9E93FQcwBoMHzd0Dk/WqlBpjfmXtRBvr4SSA9SJ7WMtpiLgpRI9
lLbMqO8q1jbkB+03je4ZYqyUrG9Q2h3BiFwv4YLjUJ9oq1xnWCaAGBbsi3Nt2GDrcr1J5y754zPf
1MriZiAuxP1DyN7oDHMG1ql6ZOOauYRjkPFqNAc3GH/ekaP4hswoNUm9oahLpLrCdjHqtrNhFbTT
XKkUABQnXLSmkAgGkFokn9L8Bq8weT6iNM86Zb+k2xZJFe6KXw3JW++SODggptRySTbgLWI3u+K9
f3+6kMT+02K8EFeE6dQoLNQsMC7ZHDBNlQhIWhymgoedS9cTlb8woMhcUeGfuiEUfDwJDrkf4KFz
v9A+6o0DWvuV64nHnE8s+EYVvVD3E+Pjp1i/u04oFWnn3tGV1Egt2nnKtHHrv/mMNxQjifsB7cvK
t4adqoCYMAXz9hNLbm3nqCUoesWom66JauY8N2h7Akb4YTNZPLfyYYwBM5AFZLrxrm7yKcKKKb/R
XVhkE9qgsx+cAVsg7xjXPJJ0/3y5SceStI8JoMXoIvytaqt2v11VxM5JtcpytEA9d26pJoVLS8X9
NXHLA8LTnaxbI7JpgkFyP7aDbVCVCumAzqRb10xRGRhGKB8TaM1CPCx8lxxQ/QgU7s0kl1kzo4y+
UJjTh9yOqD/gdtMXA8R/zvskSC6+L9SQOQVEhNGTVe4d9EwPap9Hz7HQZRnXPS9L7xn+s4pjsvcx
aaHq7SLOWNg9LEZjuWvz4/7OYrH546Df1gG+sguHId8fciFK7bNoMrTAT5mOOy27FD4A5bH8rOw7
UuG7nrJpOzbTMRoz8mF9ppvl6fCB28fM8dGwuy1AXSGxH5kh0NReWImjJAjRD3Hdjbf5NoKSHSnY
pubLOQdUFt/i42I/F3tK6hm5PUoDK4SeXZ6fW0lzYHVU4G6i5StoaE+ZNeSYMA1qp/y0/u2PAee7
eEH3J34g7uoiQOqlzOaUapWEYoxP5ysE8L7VajMPBe7W4fTZzpQopQLsp56/p751aCceO1D9UMJM
6XY7PDEXtxtvzMnuqM1Gi1fmMJqVk3yK2vEOjQPrccKOH3nXJPUrlLNsPwd5Al1p6tyfM123tk71
G3LV1MVQUwLsDXikd63ciDRhq9vCURulY/1hym/1LfCuPUhPiQsuOo5nNOOzv2kMfJgRiDWGrteu
pvMPrOxWUruMxsxAMKSY9nKF+yiONwUT1obie9FxIsg6pVdnhDfoCR7+uw2y3xADC/rRRIb+7kwH
x3nL+8RZnodFqBozrW9dmmwp8hXvtVNERHDpdlxxqR186wsDHuuYWnR2xdxtjUmKdqaTG4Mkb1Zz
9bNQ0pS/+oQsxA0VI+9gUcQkuJDC3XmURslDKoXfPTdmjnQdBOX1rkBgGONGmfzY/uWwx/SA9+Mc
uyuBvfQoEnGPpJ1KV02hInsi1mNckHvshk35VNnSGTSrieaYC++vkpegyB4Rjlf88BSSPpHfZMdy
dYY5iUA9YoxJRj7qxPMwbleMsL3wsYLKF7IQRUqLNpzEQkhNmuBOIR9542uihASKo/hJ6sXR0FXv
e/Ae5hdaZ1K/ru8C6Zb/FkPGi4Yrgsid6LyByUYpDFOllu/wQIIupdLtuQXoi1fOqH4jY14d6HM6
7yHVgeadB6mCA76NdVAHnppGGy9u2Vg5vF7vqbv14J6+e+J8oxkjj6wEB7hnXXbK077VgO5V6Exd
S3i1pPiQ1PokLBo+1zSRF9Yv7oLTaR67aUtyx0nnjvazJ6yRaLVlhMAUiOiO/Gkp4NMztJtfWhtK
mwk1pi9gKsXRw6gHPCRPccxr004XIkUJWa1WuMpNBx1Ni1h8RV1rr5joDeJ5kiNaTXzstjM//c08
cKh+VVtbsXnqljCZOYmJwnnIZBzMQ+AmGBwT7pTtrnIU0hkbO+Z4wgJ2Z86qA9tSTrOp1VakINWW
rzfhKDtcbJSh1p+v8FdEL/6Xa2Zo+5tzr1x/natUwB1WbtyYDXqHM70o9wCKUylur7sPB7bAbBfG
/BgKD5rVJfHWjbqs28+rAiI8uWma/AlS6jtaMYW+k6hHnlDUPTzGxw7XlGAWgC015PtiCg6yPXQ7
90n0BXzfNUfV3offZiE1m+MoMnBhEsXPzBhqdW4ZbdToD6yCzn8nhFEWKGrsUQwRElcbBswngtiS
s0UNpf/gzNfxA0dpaamL2ahMtI0Mp+DT9CZnDr9Yji93Zory1izPc3LyO6omkOzvKAkw8fRjxdls
dCxIfy0WXARClSZVHCdfSDyqnVRXY5c71XBx2dvBuSvsXr5tJitxUteeiI82+Vjt5UmxKzNJexwk
Yemqf+b4WvXw68fQ2N20VzJApn7xAavl4TgP7/vwa7hzOZtlK8dgcwtWV/v4rxmMe/3A9U6tVXVq
fEJX5NZDaHis6EvPjLydZHhCiEQ8OuEDkBkaWSgATVPLWCrTbE2HQDitHqEEa7G4eyMmdOJtaB2W
tHd0SxQKa46oUfurqhMoNvMsSWeFVue8SCr2H8LcrVrFefvF2Owp1Nu9nvcmFQVKU7E1gmXrgZNC
FuMOLPOd4D/1K8fszfFibhOjBrfnZqoHiTQisLjOKKYOwOFpFb1q7wJOwz2sWkVECt5MU8bIFb7K
cffWVnUolMN6SONRfu85yJ2I2zESSL1iDZtNkhVPxr3R56KeSZ02GSa2dgCmQ46kZXJSUpd3NhdN
lfFH62f7b0Id2BN6I45SqH+B+aMsNRbU3do6P8OvT5yuT1rWkK9AY7hHkSSmTT664oRKr/w1TfYN
y64xe6SQAiu66ws2JCA++1ySmOdngWvhih6zQlby/UNlBLlVeysuqfudONclce8Wyg9VrjDDYKLV
nqkNKoAg7ZdCn11f4iJGK6ZnK9mdQFHALUN3U9U8c16ZOVbY4x1Bc2u6s/AByuVgphwKYJPHIItV
D8pb31R52EDiGEQGxJEFLmXoDVtFZNXqqGSPfkedKYh84vTDHd2FZD2dcsjUIzEZEwTJIeUmoKE+
XZz4yD+M6TwtmSu+p8N+0ZfuCcq6FBv/YnhMVZ8HjTJTI30o+jobwiPMqKXH1NBErCUfJ960BEhQ
3GZmzxR5vlGQsUtbFzR7oSPK0EQDmLXDzW/0HI+8AGXqavHMFKnsYnPakY1jgr9OfE+PyxyxEgfJ
v0lkBxFa1vaVEgjchJa+OcSAddS4doVJWKHkCjtV5uBO9plFueUqbxbMZjc1k4mYOxBwpeuxdAOf
58aR3EmGcnQ2w2OKIMNA2VXTvHxjtyx+rhxjV0GQkbq8p7px2XotWXh4QDUNLqu4EeSQINLsQlO5
sAd5Z6O0Q+PWTLhMR+r5C+9zL72fxrsdQICpu0RLUAs2cAfM+0Q65Fcn2fgp3PFyOZ1QPj1IgeeI
ZUKv+m7Ph+sri6/YXA5CHWHryI3Ay6ab5fHY4CumQZ90/pTQysIjYIUNOugArZoae6O8GuWRE1r2
D+7alWNsAQnbDEHqRb9sph9aq7KEyJp9WZyEhRjWfAjCAclbouisKO2U8UZaDB0zvogJeZI0G7JY
DxKt4FfdDJE4W5Rxo8UesRWISebGvrvysA1BQD/MqrLsmrPOoKmJv5CgKH+lJrS0vU7GkoGdAdKX
3sLJaKinHeo5uoIQZci2HbA0JUwKB+dKuJAX4lDWY3K9ffeA13XRLhfWi1lB5qpCT2Ole/uRq7LL
m8l9C0brYIHjapmusyAgnU5I8eTA/dV4veRp0jyDyOp39E7zsmBylKO4wvrXUSK9aZt0qtyQ7RvV
R77SJMm+zznLpieTo2F9QxSfw0Lv+gkPuEb8im3tZ/srcpHYqcVv54qH1Or7bGZcLK2iEVCIPgA/
hAG39iVQCBwnvdDo46pO1ZkURZD7/dja7b5twqCod/rV+IVbvIto20gdYHEWYI/XuvaDZH6WQ3Ho
kpUSadfxCZZH3JJpwhmuQFSTNbh8ESI0nJ0nVc/Jmp4cnOY6Ui0h1TWYQ9Izs9raEdogqjb5DIAQ
voN+PDXlwxjlzRU59UBVGWY4R/7Fi08ZsHKa+0C6y4QDelNI0kQwD+AE91nhGJ6+OYla9QYjmrBK
V6LnxrBm8JBtndfXPbH9LYiYf2JmFIqjxwIsUS5KvFI9ZQUZoHF81EqfrWAXpvUuzRzeN1OZZy/M
qCcx1Gbx5kzxeNVNphFN/abrHGsHvsB9LLiTE63Lxru78gp1AE/P1x/JrR1SGApzIg7SuZFV8MCf
D8FaSmH0XITb+OGgu/c2xjpwevLmYzD8zTY2zlr4cMr5mgwF8DA2W6nhMtT4c2mKgHenXiF41cAp
x0zlpB0DYF2hDeFJZbhjZvGp6HEd629e3Jq6JdUTH5nCokpWT/PXfQEaKiHN/JuTCSe6kG+xOHNn
MjW96LsdPt/eX8QKoN6y9I768CFfD4NY95tMZyxklTPi7m5TxjBOdCHoEngwImKNEYa9PGJpiL9s
JdXXib2czBZQ+Ziajs9GtMXHdnaWupPbF+t7zc0qCKY0nLJDE6hzKzww+jpZAL0vBi8qAfz6OFlo
dyd/tICnjS8AJxem19kPQtod27Cy16QnZb2+eGUdZ0oNy/yRrYgsvX8Nu1UGeo2WTT4p8Wm0WQQR
X88RY+0gKkoSpqacF/+ebd+Wvw3U2NZm+55nZp9uVdG1vKR7QBygOwGVh+P8cnGyBX4vILpl/MfW
HuY0dFqduorkoiqExmszpe3Jv5NkpX1eC4dbDyk5cCsZDln2nVVp+5QcPrA654/uk1LEPs0Cw//J
fN2rFpUo6OV5L7WME4bsK+41Bxm85NrTw6kb/Y6UgoWX2IWXoBnE7C8S39RK91MLQanFWClxRXnB
3+jCb6ZS853qyIcBm/IsTwujO/6xtJAq7YkSrHk7YhM408AioVM144iPEF6FsPDSeV55PGXR/Cev
vojwV8wxA0eMi7m+J+WDNhhULJvsMCA0y0w4IzVSCy9HB10LkslgEvuY5FAQPLy5SaM6oKDt/tyT
InMYUZNxkcMWDxIctwGwhQKSmyv4ulTQz9CxRl5ruet2X4kfdUmvRsl21UnPiq8xp6qXo5M2QkOz
GNw9W+oqYnisfZUGlpKhn/Qlx02ZiKKtm+QnhNNRnP1uNF7NwQMPpx5BWFActQuzQIXU0rfImv3o
E25sdbn7afoW3mfPM+JPaWbcmcZ33D75K+z1KXUhR+aypLBfT9KlCCk6cEOOWN4B9nyliLbHtmiY
AZODszVQ8t05Y3pmKa/0g20IrMfW6H201/CVdOSUvvlki8qnLQslFfSEK625Y5Q3PQfZ0wbQZzJg
vW1kcbGp/LcoGJ0xHr1yR9IJBMQ3P+5YJu5O44UzOwUGjFDMoe1P1A9OVZh/iiol7wclaOIQba9l
TvrgLmQ++9byv70tv1ph2FOibjvXxiWTS/As6NkIhe3yi6fSO4EcIh9cvnPQ+nrTOor2Xq/TjOyE
ZcopMzu2VaYtMyo6T7UstATYM4gjyGqd3hrId/ATcP+3aITreNlS3EzcXMgrmFgLnGA+3ax0Nc5H
0r3XIcqpBTnlTJgnj0ggwM9CbEtKZI9FlY6AltkKDJh+Zn2cVFlR+NI40vyG8MvHySVpsUdyJndH
mCsB0a6g3s/aanqOeZI9cCkrXttVuZcqQHX2ccCRERtPLIagbxMLyc/h91Ur7rQU6xnSbb17V30c
0LXulEl+xLlxY7yPnG31YIOptPjXaSDJRnK1uahn0X3ngpesmM9T8xT0MCd9EmmoDxwzmT/7Rxsd
J4nNYYjF7r5aDeLjnO/C4X8lWLwkknaceV2xMX2FcT3HvBnPX6ht3oH2NO8xxCLEW2LS9bph92Sf
9pr5k6bv+fhhXb4xR0tU447UkL5zolhjv3dYjf2xtOUFHLDrPy6eLH3UI5jxjswBbWmIU0s7mp2s
PqNhY36TBTkWcAp5O57I+dfluUk5cfh/2cZfTpsFPtm10AdZwvRJmZraCak390FHMqHmCOFqSVTV
lvA4Bgg0wkJvcuJK8Esv1t6hvao7k23pc3311DXg1KDO27AvrIVUHpx+2mrBO6jPEHElQlVJo4tM
LGKjoN8KxkVGl3DlDY42xeawShnyQ7gt4pM2frr3x0AJZWmK/h+/UMASxFHXWG0SvLwBZ1F0RO6s
WQk1weH3EL8VkhIocvwPYa3fiAaZtIhFJSb9kLW0XtFoKj11Qd2kP4BIAh5+yHMoPgvgOeg3THB+
jl2iz5koEfKOXUA5ktsgMRLYDXHU1TNTe0Au8WLTSlLkORv8gBCV4WCMHt3zwWmN6vLoL2f7ac0u
4YIa3QkHSupT7wiay0SNqvtq8YB98kBl6+wPDzQsiv4VI5HOGUJmgr06htuY/QguLY3idb3fWvar
AvHIy6RxGZQz3IVbQ354sr7W2TznzrS16QjG2uj57AnpsuZ+NK8IV6NRjZI8YB5QtuEMWCvr0zYk
d0NqFaFO+Coz+fIaABE4yL8tuLFNeaSKluqI4wCZxjeSVHagnaTKZPe7IUt0jJPfTrjmgDH/lW/0
w3sCHAJ5KmKz7kxpQ6CKZCGSyWdj/ToSfMGCuYulOs1MC5sXBjJRv+kd4O99/IF3HOyyYtFqt220
0sf8AwMfbtK8xiE9/YGHlZRSijvvnLgCOkuTrthc99zXAHaUhPSUxJwHe9Fw6URE64SYiZDy7oaU
5TlvNlbYtxsHLe/vTkgTHhYASiSIM9299ObKsd3QO1rcivvO5qet6VY6yXSpWjSQuumx+9k8XZza
jT03psq4Rj84UtYe7ZBgayFrhACTkR67mGURFoGz5xJM8Eg/ESHYspNApb0Yd1hRlt6MsBJPcpeW
8YvAQcpOb6TU9K+BydLp3FHGwGO5DMy/9O2dvmJV18XTREr554FNTwExpuuW1tkQ4fdWrPNynt+c
qfVQBJGsXmrs64dJ8W0lI8EHmMxdoI7tGKt4OXrMiFq3rXPSqucf8T1m+0y3mdpF/6Y3X7PSScxp
WakcICYvF5+UeZO/o3eteK8uIOXWE0c/GFDDcwg9asCCagcztyfCIY/YheNm91mRkG8QpTSMDIOM
FPI8OjfJYxN5e7ycoZKHjJWyWMxGUe+dfNRpd8/pSs80fSS/Ou+1I7Lqj2KtlRh5Q6LEjfESVWjp
y2EwBHAeigaeX+onkJOTb5kAtyzD3LizK9v8mTmF615U6MQA/pZd1mPngvqvrgiFkDPpJcQKUzx7
c2P2VCuhX3RaEi0aAfmyeY8tfimltDmB9r8tUwZpvujmJj8ggllI+pohdxq9I3k4fcjzRMycE1i2
7gnWHMQtOH0w3+i5OnYtDGRlLkqpp528630XpNQwLOyUq+B1474HtYGmJbRdNm7EYqbn7qOFHIWZ
+fS4M1kKyiaYNMa9hxitAVF+Imu0CZ5K4wICv0fmoCD7ReHSPEu5PbguYZq2C3i1JRIm7Ie02jUd
DTVC8Gj8RqHvL4fgjAFbBLeR0OzP+APPAdfADAYF+QivO3sus/BtSKTNkAoG9CCrRjoCRT2P8MEe
NuQDSCZDAS5z+i5hlEjhVNuBNaU43XCcHPCKOJa25D66NTe/kgZTltFY0CJVz+Uw1BkmfNCQsUkp
mGx7YAuDJcjZ9mNR3sI8/njbbYPYRJakrB6TvR42NduXuUlx/kCxD7St/lV7QalVLexe/EU051/5
s69SuldVH9+s2ravmqhm1mTaRyKPS6ZVqIAZvyMH0f3GCqOWHzpu6UCQY4JYBPKaZlxrizWIAz1O
61WLj3a010yNU36hNhGs9NUOBCOtAGjO3r/809iftIOi21slnPdhwBcqqHfVmP173+r4VEsgq+Yc
HI8r82j01L58mBfmAuHCVa2EeRmqsjjWCVmuSPhWyITamZsxiTnqMeVS9dvpN7BecrUJFmB/XB+l
Ymkt4keLqqZ+j6VKhQyQCU3Hu9JK17YZ0N+ftw6ACbzyek/d/erwzhAUjNC9gVIsEjPS+i8/o/cy
Tz3SgjUSlO3nVMy/bVwJcslvocUlfkvkXDCmwyIV8ew96O0SQ6hXaLyl+Kx8rZt26GQMnLiqxBzj
ONXbcFO/nW7ULWT4DUWW2OmH1E5+DObi5tv5pK4VcuHKhCr7bilWnACJQpTHt1GE8+X1csk5kILm
2GzBtluhm6umbUwuuPegCNouipJtr4+IMq/OC/y61xL1unFokkUvusJdHRYucOxqQpI0h+YSyeql
fXXFNrOO2c0G4Qj9OqnKk1YeH/37lyb2OVvksGLW3qr1a7muafnG4Qky9sXfmwUEsyjAdFtyNVgN
YbTrOzzEzp16ciyI/o+7kZvJtVdoGZki1RJ9Pm3DuvBWdKknpBvh9q0Hu0agTSqbovZfmgXqa6hW
uXjzfwgtOKKFedMNOXMSe0OobY4D+GF2GZt7Amb3RN5ppjVKXYCb1eyJtPB06LH4+VuaiMZ/Mj+m
BRhjQSWQOhp2Kqatc8cUiIIEfJUIVrY9awTB86EnSPCp7H4z3JLZ4FrxMFqsddkzGKDlNZaHFVKQ
Joo30d0suj0ts3vKEDmCPDJXWusV1CWdsBSO3ildjrZ7uGZBKp25jZBQUBRdZakig3OsFbBnehV9
BL4OSy1ZwDiaieDwDTlASVMP7P4Y5eAesI0FVTPMFfMQfqth5JK5fxExesEVBqSm7+NfATmGBeQc
VBy2pVrnfXRk2hP4uuXmy/aVXV04IZQU7AX3Bz9PCBjfzNtRkIxbbk4x2nqNLLGaV5ET+klttSg1
53QV/5A0R96j7x1hza/WyDCtANpt4xrWeBAW+n2Nk5Lu8XIXkX+tJijppr9YBWQCb6Sn+BY84ql5
HFPAvjAL+hW06g2+DBvwmgkJziALw9PXfb4sLEgui4I1Ygx2VAb2pEKyYa/nDp2q4f6KwA8WizJG
h4YJRMxtX8eYcBRKIivxEOH3CPFbEv89hXUj2qovVFoEJmGHMGq1AflgzCSfdu42TewWwqllIMQw
+YHZNjdIJUpbkonA2W6pwofnItysRaAavOA/M5+tKk6UiqN0XqPcATdXPUZJpCx+C/ieRt5ZjOXZ
dJyuuYxw90+W3xRVprekQbSUcRK+XX49HjXYAPBHfLwO60dQY09txNMtzwo7oCs1HNH6pvk+NGOT
9L4TJWOw7oCRVxQ/5YR48YZckDHXBH55UlYCB6yjoSSkl3x9lCV/crSBtz0CRTXoGwt9+FwN8UwD
KGAOE+cfglAWva3POuQwmd9H1sKMxVrz8yRTo+8YK98JOS6NdftN0tkUXjriWV1EDxGx0VQeLYY0
mAy+HSrtaRqQYOpzSRzq2ERkCUhlUGypBO4wDb2rPRCuGZGkSWtl4WIys7iLhcAdVdjmDsGzqNHb
G2zzVGGJCO/Zjx3NbTzIHanNhNgYaXLQ+GL5bkKuOQMQYGFuhKZwwiB801UT2JCBhS6n+nE7Ig/B
m1HlWXRHv5zmS1vXrrEkmSqZlfe8uYNgbmKzYc3OlbKW0DJ5MlqLZmv1qr1TJbf2tUz3NANYCQPR
wGhlCMk/ZuAd6eyJtSVw0U9tzFB8sLmxhoY02NAs+aSrA92VpKpqLHwzwFKf+YV+awMd7Qb1JUTs
lBRfzpvfBdEj3nRmnLgsGCM+ycHs0AcdApfEM2J02rR/RgWG/VrWsY0hbJB0VV2EngmTw1cbxnZr
FCGZOeRSaufBIuFwNun0dePhRNEkslHHJOti3/Y2MYJtETQqSg+9wSQcRwXMQZMjtrbRuEMzxwLy
/WhJa1esFWXygU3PVPCn+YDBS2buM+hI7SVOChnxc1AitVpi9Z1gptyJC13ixnoePu6dWRZaUl8Z
VuEJuvDq/QWIDzWtdzGyenl+i5CVoOvEJA7msM63KKQDziHNPIAZe6dpDgh0zAGRFQU5dmKNOicF
Fx7veARWYJIlAIkZWhZs/wEyt+7OQArMsVvY4/mg30EjlbYo1Tr+0dI6R7ILzuU10pEddN9kLCzB
5KnOkOoTAxm5zcj2Z9xZ64KXG+khH69CYSFodomvKPV6SAcJv3Jn/lr95OarkOP1q/AZ0gpEOZ6I
0nHA4MX4vkHTtIA5iA/YYizawI+1MDMKzf//QncX58S+zdGi3m09/GY1ASd7qxegAMrO26FeBKZY
hY5Ub0wzZbtKo7vTWYS2yqtqXrR5qEHp5Q6hkDMo+Z51sHH/h/gruHtwed3qpYT7OnDcE7KH2ZSc
jpeT9zZ5uyHbX5YFAY0Ff0XKyf4Lc9cTaSUnfV045JgaI82MB+vrX7+U9gSa2yIgAL+wlCmOlhEN
cgbkyIEkUH8HHnPfJ0u8AJmV8uz7Zay6b3jUzcWAkOE425U1Jx8lCkDLQH0Ild5CnoWA/jU+2wdR
He6TOHuPDhwN9GojYs0sf5F/O8H397N5pbpvCMdCbuCcfHsJIJuDIMeIlhql1+2ifzoqXya2HySI
hIdTIvfDyi8Glj6b7SCm+sq4pqpo/rn7VRxDDqrypU9zifzERFiwdVLvma7y1CyUm6OGZmk6pJ6S
rzVHm5LX9OkTWsat3NnMP+qNLnNhkl3rIlFCUO8AK17QIjfsGARj1i8xLtHsH2yIZn2zrUoITVOQ
lKhp8zKbCg0jcGx/RyYG4yI0d4/7F7TPUNem6lJMJ12w0JP+O+OgE+LdNuXtFqPVF4I+EuENs+MJ
e7Cosf2b2bFkBsvz95EL+v5BEOnpOBcsuFT9FaEQ+TboR4mFbTCVYrG0oY13w4z4lgzV8hfEtg5y
n9dXorYMXY6Hjc02uiM7XeUCmOUqRFw4AfPR8L8OzWy5vI8sDEy3Nt69wLy06+q2rncessuGDA5p
gjo7n8NdP+1NJshVy6aqOfvEtkI8A6mQK95ndFHRTXF6ggCKvUb4M/HAh97e+R5K5lngDgiEq9xV
9ebgXfsi0RGNBkPMhKc+qQbtsAmk2Xixkdcy7oJ7NDXdqEv1FA+2Q0wFvyBfMq6RgYl8hWKLio9s
1V3PIoCkNykNJQJw+KP4IxS8fZCvoUqev13ebhXOgsJKtwf3muvSmfarepf2SW3BuUL6++s/SgUw
075UUwHwaEy7Osv0hfSVmRT0f8YtylMLU2r48wdpsW29bANB/YoxM7n7YAttzh8vLn+GrxtVx/Ok
HnoU8vaiwKfrgH5RtETbMMxCNdfKt/h37/ffFmlqTWzFFTAcfkQpMuEuNdZ5WAoZ0EEiQ/xIOc6O
YPwwnnkXh88pwONnhQiohDsT9XmY2RRdYEnKh0ce6FGce1PVSdFjxApu9+LIXeYfw33kVfQw1Yvb
uZsu+qyiPrTCS1Xib/gOgvihw2LxK/TOh0B5e6thxrDn7Kb3GJUZ5GpJ3vvKLYhoNMGHfDWi8Tpp
52yA5cHy5T/r9QflW67oIbwJwY0y6kKxOpBev1E2Fmas3aVxHh0jB9Ik774DjzV6rv5G3fEFPLA9
Dx87H7E16tylGAa7QC3d1WEzc/InQoWkw4JshSXeRnFwqCK6fvfEqZO8uBbR+uCeQQduj1awNzIj
m3J7qjvqEXQ3mo/ywS73nx1V+OkF8KcLZ8sgEJSBOZxKqZlhzuo6wE+zj6fastGUYXx0BYbbnGXX
Xhsi25g1EEjTrQ/P2Ic0oBVwbC96Xi/iQac/sLLO7dS4KfZ9sDkBUcq1IgVJbc/wxolFFIoSTEbc
n/lbvoOZJ6SbldaDqtTNvK4aoUPgpT0YApIRYcZBzxY8i25c/PHEwdXPkl7bPsPcy1V5nMxJxEDd
Z84JtwOuJj+62q14covm3IqFxSexv0XVjaNc/QczW5t6esfEJGZm53QHVKtWzvzAkXMNT6SmecMy
CuRR2iXuujHJ5CGUV36OIBvGPFUnh7iCRXejxGtSyQd8TKuykrdeoICII6t2tZlssYKqXfP7M571
7fGzFSOPuqqfNhvXrzKMmVL1Oo6v8yhnOgq0+ZV2kKKZ+oWlKAy/AcwD7UTDy8nf+89Sv3Wq9c1V
xPiaB8tjRwH5JNtGclrT6XMtgMBDlwEaFIprrnDnFxVbxUe3Y0aZMGvQQBwwiB0e2TeUFGtsYwAU
QkXiRbAHgVlQe9a+RcuhSTI7ONg3L2yBfRPC9+azwGZM7dxL+bqLMS7wV9jehBVYweHTs+rOVlnM
QrMMs7z+O2Pecr+XDHVreyxbanhGKajK34IlXj5JhjF1oFxOEfOBS07G2UXyvYEYUJ2RsPDHSDvO
Jy17G1cE6mOs0vvCv8jijVIBP6AEt1Iz45Sw+CvpT9V6zNemRYislV1KOPrJEw9F9CNyRhYZVtcJ
4LSMnMGcV1sVDkYRWKHi4z3wcmmz7O7GSKQmsuIn0qp2PgzcYEvZjoJ1M6S+6JFqNgYR44mS/pgD
9hY/S6A9q6IWiLSGPbn857uOlcJdHS9ZWhRgdfQMbD7ih+dIKVBLyieLVkp2MKCczOeYBojfpQ3v
e0fk6h3xhI5VnvVX2ZYi8EjdroQZxAkxx7BopzrriFGjA+lq5Y0ImVS9eQLOgliQOtbnyCln7tXy
5k7q0NcPnfnDcYtdFFB7v6RGiEVGCAJrY+Qvx1PgBgrGQL9c1LeJqLR8F/1KbybgxX5/r4Q2GqQi
0g9+12UbEpNAvFZEWrm59AHlphlnXwD31SNYOtDy+2kiDG9SY42ks4Zs4EdDYV4cmAf90a2MC6RQ
5oGSMgqP9X+TWjNI02mWxX3QeYHwWauiu/56GOk4KHC/XFGXQzRn68Tri5DHhddS3+w0eFACB+7n
PPLJhzxyMt5d3pjOKhby1PQyEuWLCy10DwmOLaX+B/OlKLnShcJQG6K1RStUAYZ225wxeyCfTLkW
l9xJHergWVJozUNeXejDxF+Iz5aJ6LaY1KG8CDEYAG+mf/oXGFqoWPt4HRNkQtMeW5T54e61ycTT
84IzgqE9Pz74DqXfRHlGO11Zxt/tqcSqWIpaE//+wVMzh73xeMWuU0uCq7380DpzQpvLX0EUlj7I
LSZY2fyBKLM3DJENbO7Zz8Hly/522VIh2A89xJLcWjunr7vVvTVxLyseBoCFcXRbTGR0fDQE/MnZ
0tVNpPVYL3zTUvVj7U0QNPxYBDj+R8wIdq2WxyFrZAgEY1W4OElNs6Te5mBwiV/YvIYCR79xfSgk
0wtJ9iZBgo6GYSrBoAtOUZ3wh+70se/iEgCa+w/4X2rRUXYkAI1LEX9a1IqsdFgG1HdQQ+M5WLZC
zt8+n4tr+0Jz7xX7LrX7/oSfAbqNM6E6y2GR4U7KfnPlj1npzSv0d4oEeODFkrARE1mCdXy70Wn+
/HC1i+d9P6Gn5V0lLexsZwPa+i1kU32+iFTakuO9Ny+yWIhBARW2WGosUPxK90reDNjMKcDsJhMX
9UX8bj9rQEVVHNsXgvAYzDOnjYnGGpiZaz//qNNTpV90DrlD6Eu2rf8Cf3u/RL/bWNQCJ4NzTScr
UPNifh8FW1SMALTC6QlXqHOOrQrhXXn3q2KEezObHa/c5ShmwEqL876qRmfRvsvNcHMwO0+njPXa
PDruLb8Co3Pzqe0XvsmXHJcfDrH0HpiWZBkSSI80k19dAMrOocnGkddS8qAzIWc1KgMMQFKmCQjN
F3fHH7ETWzfSuHlxjvSZxUFgrxSuMf5YK3SQdbFBQWOBTiz5pPGjs3HP1yhgv7o8ane89UcphZnX
LrDf1EftX2AfSw7jJ2QneCLGmKMfPbi5+s7rgrV+CxVudky1ON/4MTaQUgjzQdo6H8B0Lhbjr6yb
pIlEzldnZKffi2CT/jhnruqrI4pf1znXESdhC7fqkuEoW+x1gnoNVwHLorHcgqTRbfv1wbxJ+B8y
pt5MuxWD8cM5jY0c8c8N1ykIABSLKbT0go3osltb8HrABY/9LJ+/nINLm3yXgLI4EKqbODREUlvM
035Tg4Oou4LUqdpiutpW04ErfA4E1S3yiqCHYgMS8E/PgXDk0Ji2uOC6GMarSviBR/mv56884z/t
NMEjg/0J3HFGcR3C/IV4NUh5hSVYFaMS8xKuJL/5eajugOgSC0hlqfcp085gPCMGJyGnyFJYNz2H
RXAOUxF8L0OrZP7sbAM8iXoWbCOyVRJ4xvbelAjCGKdOJSP07B2ttfN+jEp8dLYt6V4lqgQt8orj
U30PlCe7ySPinCr6E80fni5WVJVbB78Zm23mSrZ5EX2oI4TGrYW5YULMoHmgng6D6B06G+ZJ1jng
Fr5MrsnwO47c1cYsW2B4Wgl7ARzhrx1bLqmkmmRO+cSfPJ/VCoZ+iOuQjRLxQHiZ2MqIkqyMJbCr
e877KdGTDxfwdAIDdcaMJjxCZzohWBH3vqDMSxNPC4TYXhiDO0/w5hyfi6DqYIs+3vcrwfGH4Jrd
1Kkg9FEixrckqnnxsINCBV4GNq3EdmhAnbCjF0ePoygE+vcYkbaMGMCdExrWQ83HuQjnwJExslTI
uB8ps2ZtPlzbDZB12jGmX+RYVkUx6hfyNLy1dZGElT4QvL3ywhQxJDvul8wRkrCAcEMOlNCfVRJq
uKmZft9YyPKcabiCNYGTrcnrQ3OrUDqj0WAqsHfnpchB75KF01mwIzSSARAm47lwbXszkEnSgOFQ
yP95gyYrWraHd/gquGQg4mUhK8cEYBwrxe7v3cmKTMhG27jQogRIWJiqig+wP6Gn7/Fdsdz/hbE4
MSckzSTXf1g5yi7w8SlkA9UMaMoin78dc8T/fxghK/wBTjOq2sCAmxk0pg4/Izc1Psd+ojyYPk1V
SfHQN538FdDJmMBC2dfNo2ttpWwJaRbIQ4ea7TQXrB5esUEB5EzZrpO6Y5y9tYhmRDQ+30TCfS2O
nx8bAfsJ5ownasOgj3M3+1/Zo2rbmV8ahI236CGRmKpG1e4MTwAvw32VZcO8JmvZOaIh2KIP9iYI
vrQ6WC4nM4IXeuh/ClXi8fPc6c1j1BhYR3CTu9/1lB6g+qlcTA6/a7CS+JcHnwZmj4mQhTBqx/QY
L2XT0Slp+062QPkyxBKSPK1B5q4klmamybQHz1oeEwwVDKGEsvaL0711pHnQsj0x3bSJBuuPu6L1
lpMUAwrurdDI3QAouMQmugr9lfwtkIcqS47l222SdGBF6Oc/piI4FMAQ38vbj9oxIzq6/+dCLptG
iNXiQcv6eKiCtPRh3Z7lxukPo5C5RNKkdBM4x/yuQD8/IcQPZ8NFUHNru7No0j7b/4+DK/V3lkub
ObY18UOhlNvVvtVnRjq3LW6/u0N6qEkxRXTv9IEPsGtenB6fLugzPqZRBIwje1zlE8oKxH1Ou0tz
covX0aAD44613fjRGX42ElYtbbXdZgt5E8HDCxDSxe5YJ0uWMI2Kd4ZLfQ2ktPrHxgMysDsuybMi
rpqUXLM73xMub+6xcugoASZTbMIHvai+4AIhX6hdvzKz7E2D9rKcepbHBp+an8H+CIje620ItYja
Q3Oz8cpWCo8clfLpfA++sjIxidREHO3x7Y5CcliyMA1ZzcuudA26h1VJv78hkx+RvLR7ntBjFtCG
eNO85JNe2HJNadt03nlqJ9j5UXaO7JVvU+b4wgnfa6Xo3sMmPLJDekeEmOSqMk2o9DVeY02ynEXc
wypCmTAYI6+wO/FWZ+3EGYR905SQZDbuT+EUmQCKDPGm/uK40Fvdkf2U4eD5t9hh1h2nDnDyhRuj
tr5MNWS1od5VWZhLYOs3Es4fsDWVdZ88kPfvNmw+XHyIsTR4e32hyVnxIkiCI5k7kzwY5E3H55gO
iVPkvgdQlRRF1ehkqHIiv1viE8ZKm8uzrjKdcFb8YQ4nTJY6KCDY3VUo2O55VY7VvGjZipvda9lh
adcR6cghIwnN35vWGnXA4aQl0k22y7Di68ig88di5ZdS0Blb5WYOZuznPrmna2xoVgdBFB4O1cdT
7kqD4D0fTM6qeH1fZBXSDJ5q6hpW8StUKG5t3jNjsHpItTpcgI3cz857yuWz+YG7D9FBywi9Li34
6DBYRAOdCIgQ4vrd2GnGRoeGsMPxqbgrLY5hWNUEkLApWBdLmSdcLnx6LpE2Q6+LGuG7MmF+2+9+
Rp4i5/oMzdYPeb8PuMQUDsErlvh4UHjTG1FZ8407OKhlmRl6yOF1VKmk/oybMsCDFXEAHml17cT2
h6KfpfZEJV+rriXh4t0VjIU1crAGyJ+A4bIQVuOqeMWcbKy8+ImefqSeuskp9WTNxGmltobDvRrM
k7ItZMdao8SyLA3dcb7MBIB9nYezM2FKSJmrFJdAHvq7ZEScocVA2uPKVikdjqCN85275sCtRExj
3yU/KzaAnAvcpZRlh3Na9ZsjG47OfNMZv6QGaPp9zqaOyrXxeRbplX8td838jfkwMyIplYo0AVbj
AaAxptWpN3OHcjsIsWjuf4Gtfbi2Amybo7zoT1IfCx24FvV81jOCVTy7uH1Nljy+HBU+ZOLm/Y4Z
CGyTAhfsjnrjrshbuczsg7ZUzNRRrnUJo3nFNRV6vI3o0kaWdMDauMcbEC1KNcdYZ2MVycSjsypa
+5OX31mGrcSDojXSxnhYeJkz7AIMUYlNM6/phBlGbPXr62J+F1EwFMt7vE9pchBcBnIVzM1/K25X
MDaVoakHYKHlJzDL0hRgULEDD/te5uxfCl+h8eoxUbjlfOGhQkI2zcGaaddWq63aJjCFHP8Kw53x
CwSQqCj/Y7p1U77pmHAuwugbVn0uAPMT3HysCFa4FWAAWJz4H7IXWvgsFCQHm0GnNFrTBw09Ju43
puiG+UdW8DmMPI+1v9HpVSHTfo7jyI3sXnwbqtY5sPvxiYAD7R9xy59KsZY6a45n+yNpNQSpYIdP
njOKHu8Wow0xP7kcSFU/i2cmNz0baHvJALqhMgGV4fuU6wACRW8JXmbDHeDzEA1gXVCMl9QR/ZFU
lwzZEjCxoZiTFLg8LJTV/QMN1lTEnV1/AT6cEu9Ety+48EL/utQ0R993/ysDeapKJJOSQNtTu8sY
cdcRkqkhVgRzmuHMbu8yUrU5QKIPiEjjaPhvaTc6mLVwLzxgxcQyCRZ+0F2VVIII5mQcTd7Xo4uY
xJEfWNXxy9VEWOxxHCAS6MkqOS4Ubdm15h9Mo4f8hTq1PdmlCgJbmG+2+Tgp0fdtaoS8woMgXJtp
4GFe6HXbP5HopppFDjudt7znAbXPJGfarnXeraDLCIouBjpm6qJUyTL5q8kS7LvUIu4nYx41Dnmx
KycO6Lk4ultZg9wkL93WpmuCM7AfwoKrH2kzr5FPc6uRTt4siAg25FszuebObVXtoseD6drYGlzt
zFFa5wi+HnutYX7KNhlluMzHqvj9/w8wJXW0q/TzD2KIsr3jFCAGZwDGEC0wQ6xRLy8aZAtEPFjM
yqKIHArLNAWgE/+gIP4buRDaDAQlQ4nqPFrI5aFvI5/GMxkmzxWtM2WEKU+4Usk4FiehMZRjw5D7
8Ax5plw8SY0FID27U45AgkzFazWsb2yC4FhQs8RPyTcQTy5uixPjebifpRwDcZk+lf1Yb0pB9frs
pgoNf0DzwNn2Oyfiab5mHx90dSqW8eiyVw4+FfSBWNLfOupTmSPUKDw5mDKX/oPfk4TP3hHTNcnT
tjljM/m5ZsYnaxH1u7ue1TyAor/Os0GJTUuIYr27/K2o0wda6RGzYAHMZQ8ro9zy2UOv3HYNNmWO
VGOYx23E2XaJSQCrpPdMD9jN6V7LbUsBrvkfYTM73fvshe1QKJqjo/CEedNadrJm3sKrLncGVP5F
XN97TSWRvDbtl/5gE2g9lSEJhqfDXzX3lXcXilIg03s+ztHoMbtOXXfk8Dl8h9a8Pk0oNQvwm1Cd
wVqNAdSf+EE0YEGPCIR0vKWRTvn0ETY7FhbtH+xj8RQ6xLYCHIxlEcqUU9xOwk1L3NqzzVLcj05W
g2wVjr0L9tpQSytPesYcLvOf6xw4QUwHT7vZnlyGub4HeefSHRhUGz3KCMpvEXIqezTCZcdkUqxL
ETH+AutjsGdtdAQqj/Y/NgDJYrdAj+XduOA9gAI1mdE97sJ4tkNm4D/a3B2neXTc5yV3Sl8iRp7W
qkxfN7UV91n6ZMPXynHBnN5RgrgWGsebhVAKNj+pDSIC4ZdSbppsygqrruuHyWXXea7uUM4AkMvj
EIkCtM1p5mTgeCDg1bx1/n1BVTWgrr/22pUkr5jkJVcZ73tEIN7ZBQk1OvjCjaZL1puBYAph+St5
vJ2nzFX98jZKcw8jB5FNpIydempGd1rPq0HvXwCzi1dL7HvQkHyEPEhluPQfDd/QRphBLfeQP/cJ
vNJCG9ms1rjkK6KPpmC8pix8tT9q/4VQPwTuzq8EVzZO7nFYkD/VILBSI3X50AHdmce+zo9kjNHD
7c7hW2W31SqYXBo3PGzTyAZZXTlyhjhhzrTSoC+g6YDYoFzwd1PM1YP0uYDzSf1j1WHdJ0DxkIm7
WQ8R1uQuVpJa5ybzSYwY+4OaNV1haxJiJNtmCgvQUrxWdMJiJwZ6fdBwVKUGW2jAKFEFpONSMQnM
ZNMqnbXNLiNCnVFCh4fQ4F8FS4XUwR4fC8CO2WHMuP9M4N6ahU6DhWemY0tD9PYoV9jEOsz6bca+
XLjFG91bvVQ0knXkrgefHrz06Gpiagjw/4BJ8NNgG2MDvlDPbirNNy+e3FdjxgARsjMd2gaQPSNS
MfQ+XqvKRPtCmBhuKjs62JP/Gd+6JmSvEJksNQ/kDKLaHEBYLTUqIfupDp2QtJNJ3vmZgLOMsaIM
GAFcq53r9xTShx5Bjz4AuWEgvKPb5XF6Baztu15td9qBbk21NvXSgirYZMgdTPAGEYJA9T9D1EEv
8CqqnPllnTAsq6s4S4GG32n/GbymvOtdO9bKrUNRNk+g2tjfbcAsrw9/p6kDSb2YpsE6RLX+kbCG
QWha9tH/XXOYH5CUkYWH3ZO9BXzQHtRRjM+8dsNYiij4JsvfZNDVWmq5UuDHeqrjKhRWfC1HvKbF
8GMNrq32ejotbXECA/wg/jOEtlgMRUTDTPFBK0EXHO8tOuS4U0mLdz/TRVGEq4LEfpPoTqm2adjH
LxkH8ko43MPEjQUupMlGPqvKLp8+mzy9iIumtBkQeFDjkfZdQJIbTf8jOFh98y+dix425prGNWBY
pFsW9LIevz/kdHLKv1IBzncbUqR452+/Il1UU1iLxP8n9O4gcyIo4N6vVC+LelJ5T/egQGbuhrZk
Eu/sw7eIvf/VmLJcv/YMyOQN100M3CQjgo1SlfkHzFDUebhyK/o2AShy1YIz2T8jQ3xkt1CKs/4L
0LVjREEXxzeWwJwZj5WJn9PQvUx2K3w1NxwwheD6WVugLAqMwdTE2DLS2G7d1ytD/r3S1TnllIWk
R5GnIMN5LeP3PA5fSibThHkMTuO2VkiEzcStr/GcB3+IVHelDnfs+IQJiinfP5oSrI9LN8Rb2FJg
BvEmEMEM7gnKMlNC1VQTNrPq6au4YCA8f0RuixY/m9r8s3aDGUmQ1cElUT3MqrTSavNgIGajOo31
AmnIeQGW2yhCIil4XqJ6FbY19DK2Vfm53s8HL9yw/il2d7Pe+dY1ZCIWyIjPtVqrKFVcZjsJBPGJ
ir4a2prZPhVyZSDq3gUevVKVySBdhe+b9OH+XIb4F5YbUPokYwCxtcEBMalH0ANPUk++XjyVXXc+
P0YZ+4rOvVHOQ6npFGO7lqgb221zDwgr6hIvO8NbQL+jOn05Yb4euz4Z9hRV3iyKyuk8wz2wLDrR
6nhO21l9yU1bZO3rH89CdC6rWmR7FNsQXQkGVMnCdQ2OidScn95vH7kxZuC8pMYYR5M1o/bRkzKP
I++e/5Idw7ljDKEVj2Q5I2AfN/68yiIEiFW2QXKlKqvOhscgS/6l4SJD15v5duHJcE7duB2GYcZ4
P+WjV0bcwBPUC49Z+k+335gQgAZBTol18ExxyVSH5XxUhj3uR1CAHVQo2U8/CBGPjL67/FdKKv9J
3DE6ELq5K7hwcjSzFO6UYe8kTJdibWrobb+m5ESfFlg1TABvJ6UKp8pfIJk/ecnb9Zx8qB/BWeOf
xjeOBmXnyBtGLEpyMXiPyt0dl6dECzoJj1GCdID15XfpRqkeJ2gnXCwYagYWktl3EWE0kxq2MMux
0kuVqOaWT7F5JMCBUus8mcJlDNsHQ/JxJpSET/toH7eGIYEMB3J2DU077HXd4lrlorrJRU8qFd77
klO9+ABwhAoTq09wPLSbCzOBQWmeOocjBnaXF286ViCqqqyZ71GQRARyQvAdo6h8TEAzAOTRnAbD
wZhxKK7PD5igRFtaGY60HRetSNpMzyVe73T6lNKFxiINxds9/3Skj3/QIdBkwgN+urQ2reHYcONT
O9yJl4ifGg/vxY0avR11KN4sxv1aNTiFOBLKlT4pzmLKk5yuZiIVbjJt1AWvsLJ67X0wKquxl3Nb
l19vNrHN04mycMoOn/UKdVD1H33Nth1pS1ZPVWhF1MHZViAkT/fZU0hzWsqS7ENG55Dge4y2SB9I
LMYic3ikNsoka3MX63mdXQdhjbQO4KSrv06vyO+ArI90mMgE9xD8UqsSKta6t36I6bWfCGKxjH2l
qFO/ynXeikeA/6s2z40mQM2vR6sONwx5WwGVhGw8Md5rv9VwokIyFRu47j2T4ESk1b2JXA8Sndaq
x+mttvE4nEglq3qxZ1Z5tCfhAYh20lWbNPqZRrMZHl2nNfGoNUoPE32hkaMB993Hpg9iPa7opr7H
AQtG1rMT1Cfx/cbNHUgRX2g/DJl3j1c7TjAzsNCh/h+VxVm+6WiNinF9esjCip0sPJrS9K2I3BjE
ldH7LllFt8S6T/GMBXCgtEYA3pzQkAosDQpI8iptCM916tKIzZfA+dAuQk4h9dP1eidgClmZIFxs
UuXtXdpCazg8nSc+YU4ZWDhL1toSeldt+5NqlgCMr2JdC/mv3JRoZ8q6pcJsmzM7sqFndmr3nUng
mBrM2zDnF1F6mO8gq+dpJU639FqOuWNcYS3TJ+hHIFajZMalbfUjx91RKYwhaInRZlVr/g4fLFU4
T+E8LfkdFUPoU0AUPuGu1n9wvHJ30t+02KeV2lRbVDLii435RNbFFbug+joiDpPoibuitz0uwFXU
W2utepXUDN1uNZSSDFkHwnHyfmZUK6wWFeFmVODJ3/UIkyLJQFF2aKuVbbCoNhF1H5G5d3GJEc+R
yoMRH97bX60nnIWtJ+l0xR/iaZio5pra54s7nkTyUSZ1/zuHeC83aJqYY/+QEEnA3bW4hcevCVnp
vUtL0JGWvl6j3g3ThYOZ+0rYE+dv4SMEo4j0ggDbCdhTXpAPIo3Gtry7MqxtscuogX9mPygqKvGK
F/Anv2nJDeQgXvteaZX2hcpo87Odfr2IacYPh1Mba0IOxoUeQt5XqylwClhOcZRt0F2PRaxOdC3t
eoHMg4k5jGDQNHvozi8qey9X3rzDrp2vEgca5VOFV8cyTQ4AqQ/c6Ik7Axm4HrJQHugevz5QNLqb
BYCxp8op7JgPYNUxFKXjeJkh1dABo/fZl5nwVcKFsv/QwlTW+BP8r+j9k1HxHYN0sDL9gGJ9nB1R
OJuSKpjuiM2/mHz7e/hc2RSdtn9tUnOJ+jFxyN0NtvqSIb2uBm0u23HBQH2GTH3zrQy67THwpyTP
4pO6/g0xrOk84+LWPwbkne25I2zqGIW1WVzjDG7T7Oc+oUGlR6nbQlwDiVEccxv9zXRZ5UEp6ICT
x8NfeQUjt0yHBylrzLgxOmwMSfWYzX2nGfdbfAWmn50iE7ZgRrfGMRGIqk7wc6eBBbiHThTuD+Ly
vC/BsLlFGiJnJhz2aRF8ccuHKIkzK4V7bw+Of+xV2l8PUnET0hDaf4I39c7geSjlV+dAclt6k1pc
3JbmrQ/BY8BL7/5fst2nwU4wXie5PC04XQZNAdOItZ1CuqgRDzsHM2nMrmShXrrRyTF42qKn/Ls9
cBz7Va8lVtMrLGqgW1AZGwg5oiNWeupCxHeP5LwMZctjoC/zyYMEYSC+uJDZMI0vA06CCwdZUTiX
UsyRqn8+XggtrNpz+L7VYlZWBlc/rJtvHQQpIp2fIpwZ1Z8D7jvTnXVAZ/j7MDeYDn0u+yUkw9Xa
62oFR4/Y42wdRERTV8FXyFvWNs3DSGuXXlYvWBe1ab3IqAJR8nx0SvMNko9NWp+r7N7g/mvAzPIW
8CaEqL10PxRU10U4WLN4Mc6IeSA0gMB74xvykQpjGObELkezHbtqTGLUeDt87YPGTSiRFUxox+T8
QY7SkLA7K47/TjzaBu4BeKJ1VrXwcmnY1+Jk/+WKw89GiJ2GhDwPsgSJmwS5NC6mzd3tdDQAsfmb
xJHBMr+TuYXQCqzTn2mRvAX0qHJ7fKSY9EivX4W34JzMAWn+AXTS90HxwTRyYTq9DmKpibTUstxh
S04jVX7sUr5+47+ISVq1XGOd5CWteRlUUXA9jU+rlPhnSKGiBg99hGHbNWig0Ooas7mzWxZ+2GWh
f6yTqbH8CR+LU/gNUqoOd6velOz5SqQQUHW7dfSHRz8HBMrfgOj8i7p5PGuOhM8c07POXE9iPMzu
HpVYFXb5QYPjpdb7Ys3LvRdP6+paOKLWJfZqDvafxVThIA/QNPEFEUn9U2rftI6S5VyZRbgNehpI
M6vB6oMwQi//jWSkew7u1wjv71Bp4GJM9PkI2x/FAKNPSMyEG7FloRcBAEWkxVVD4qygpmJmrQ5y
7fx5uNWvL+WUkDVXp1llTCE+qwzZmiviB/G7F4gvZLo/yVE/YQooK+FGvfXo61zW+nDFku75KFJK
HTQG5JVoztmOQpyfS7hwV8yyOO8rSspI48CudraaSUM1BC3b/Mp8dhHu9zsLe0jgZ97DS386PAC4
pylJ+cSXGe5GIb+fzaXjhxKCnOlHXtb/AcKisYhCk2noygizkR/LRGOKj/oaHeXEXu7Ej1iepkjR
Tl+mIg17F1tAB0jNp3sq1fwWld3R/2Fze8SLesejaJPmmhmL0b34fojrvIsL2vpjSFyO/g5Cv/qH
dHY8tbnjXe8DG5KSmsQ0SF9BIjw2LKvuxIN686d6A8VwNzfaNVUbSnI0eMp67LavDK18rJ8umbVU
bx6QwWk3+s/mDguOYrmS1KDCo2JUF2IA4VcfVklQjvYvqHyDFW8akBM4QHT9K7v8fcy9LwEd7pR9
1JLL+KWgrRojoy1RySkbOXgXMXubY362bszwvRDv7TRZ7HNm0GnzJPjXLB5QtDTuBIoqSGoSmks9
kxhyuo1oyHpo1guv3UjyxwTPlgPKCjzXmEIrMPJIKS+3SyIXYcUki9dMTes2dqetGSQfAlRUEN+r
Cm4cTJmcqLYxnxIZj3J0SpYRYWJaMiJKmfqHMRdQ//x2SRYvFALidE3K39o20YsRCpUCWcbrXc+X
Mnzue8nTXl+W1NM6P0MpaQjImXmKyruEMwu68Y4kYZmIqLiyn/RHOH2DJl4LDmXtlY1WROpBOjv6
inCAGVyUjPrXwJrJYLXQDWJMpWl82VgjXGX7APFlMJojUSuNFVtdERhzG7jGFtkilRjHyucf0yOZ
FLz0DGAjrJPS7wp804LQ5Z0FbHxtDf/6bQh+8bfKovt26s3tecXlCLfkS5bcqeahcIgnEDB/0yYs
pON4JpD85iZGBsL3lzCnslxu/FNl+xG5EhGui4/f5swbW6SXett291ofMHDVbqe9Nn3jcYD1n3tW
/98BxS108GZLOlqn+BnGb9kXnZ8s2DtOPnDqPEuRgqBSN8a+dnZ/q0EmP4TIc86iRB+jbETtkqMf
7yV1YchHScRx94Sk7WeJg7v2bhhixwcpzUcHNQhaMiKUBq02MLmFZtQu73OtZpKPfTlx018oIxxz
oBJGPAYAxVrJoZUZp1Ul9O+yP1D+aFlHoFLZI35LDF+DParwCsjw8WJMkeR6o+V7DX4CP0UUgY1X
bnJD1sUq+t7KyL/9L7SNmf8HUYWUPT/PzrlzFIRyRszKxWJF+uRPXPkRJQrMGHEnJ/Y1guzCzOeX
MHFUyUqTBHW3Q0XeKvNzKNSaj4fZxSvdzJC/pLEkOK6yik4UuR0MmZZsd1mS9ejlK0rliO7mkw86
4Ty9NF2NHgKUoMFckuZPx1r0JGY0Se2kK//08YEWYPiUaBdMTXKkXvZnWqHfaaUV6qGIPl2mxHdP
iI1v6ulrRcWp8nnmpdcLuBXtNeF7JrZ8tPFd+VOtwy+wHL9bGfgaSYmO0NvUd2QWJcGSKwx3YhxF
t4X76F16n+moz85yxPLdn7DKCGwRonzxlNf6u1LULAs/d6/ksEGhVUOn2jus5Q6EgMg16MXjl8Ze
Ghn8x+XKYSc2M2ghJn0iULEfrGcdseXQrGMlYgiaadkxGzzPaFlHUuSUhOMoQrnOfxic6UKZLgPe
PSaFFCbevMEDT7Z+UEm6OPryxazVxry6mvTu55k45iigpn9v5CWlnN4LwQTIaGmRQUszxkXVTCOC
OOiYGhojpiT+pwY2GfW8GjGPFsDYeJ/CZSw+pMB5dydIBCsTv88YVppRdiLy3+fbBNIZmY07ykyT
JItVKWPK1Ro6kC/lV7DKZx9JKpy0bznXpY2xCDpA+1ava6XHO4zNGAShVeDFeW1LqF/7h2CJINKT
GY2NikK4YSvs+zw+BCtnY9lrA5N6CcHfEEErcK+fwETLIgXI5UrqjNDL23DPF/0FYgp6xaXqfRk/
zeiqKZX1RxAxlw9yMOfw9sMqLcmaP0ayOi4+OdGgwHVxZfZ/D5JOGj4WSAXf7rry+ejMOBcdHohr
eiNfcYCszYXrwApYU+6jvIVSp8V+I8twMmMSpZxyXdx4RnKfP1aKGXUy0foZYmfMS3Sq+Alzv+ij
hzcrsw/4DrEEP6CG6bC1iHL72J+jhjuaI8M7jtIbHDHQJ1IzNGTzzwzGjTQhLZOhsAwgCNmCgnP+
sY5U/sYrpAv2p1QsqWakKNc9SWZrM2RnnPuEAlFF2FclIDp95SGVoZk1f77Fdr2wlsJdUy+ka2vr
tW6ijRkN8C0z2PjjbLkKY5GPqVSobD0j8JYDMlptifPJNZyTkouG0ZyvOLwach3d9Qjoewpbhi/T
Bu9+SPnwfCevJaKaTmXQlKbhBgBDTkBXRvjh3AM5upxE/7m7Z7w0r6wMoDqeCQXO2HDfxP5qP3Mn
IAZSdVug/9Behqtil32XKEE5JjBLscZ9x/4Z0FfWse8b7PSdd6gnlhz1DtX3y7UlyDWbtz3WPZVS
JkJiHIu6BmgQMVolGwBAhLJjSOJX0x7ASDRwKW0m5/jd7MpSqFHfso7bvOiocKpnOEtPdmoarGX1
P+OdIaJIEEGaDkocplz9ze8AhyPenKEU1vYPjXwl3rjn1PuzEVJl4xTPKfp2hmd0LTEr4ZknXIMi
faQoYtBBctTyXpMs6bOi2fO96+expxysHTuFQWnfm55O9wX4W1bcG01eK4zOrqnIP41fnochVlJT
MUqD1lEJeww1F3d/AkYD4+XoR5nMpCM4c+bkx+RYJ3uOxzQyDr8ERbGOq2qJHoLG5jqCt/Qa7gpx
tTKEe/Q6/5BMNYo7RrvnPG5ICuKekWw/ApJpOhm6WFpiNKLhGzWDaWBqHgcd/EMqtHYwNnA9ZbU0
naSrffBwfxnuvNd6vn3h4yq5Ft04j5TizUzTMIRr0EZiucgblF1Es5mrkcLlEEqKvDyleikymS7p
aEmyGbo63FZdk1Wdgs64zPxCzfEDbkMdQb43VM8b6b+up6+Pb4HRXtUp1Rpi7JzGEJ/9vQPQDaPn
ALaemFa0+NW9owQae4yoJWiDg3bCk0gNkiuToW9ggTcv1ygScjQQ2FZNPaPF/rPl9k6XxC4PMfO1
TucaugpO0hsFMwZ1VSABZkY5HA9683mmvzNmh/PfE5DHrx7wC8F66IG9MQQkq+/jlsNYP3pPW5jT
XRIjTmDlm3XNY2Vv6TZJ71U8j4fhn3ENAWfT/nO5h5lkPlQdIXHyGB9KfXD8LhE6XNDD9FNOTZnL
gezTixkacDCnP/TidBjdatg+yEHxMcrfbSNjypzIlGXBBQFRF4mICK+dRsFG4I+Lybc8Uykca9sL
zSv1jHjskN7CkuCVsxqnLpEhOTRWOay4wqE+jkHqCWUIbLlO6GnNtUgMtjAFCgjFAzFUHeVtNd/l
mT7jbbOQotSw9q+gM3/Hi/s1CHymfvpM+9pmd5e+dJK4KQiKyRn66DcoaWo/Af0lyOGKNE4BjCKg
N3QwWvT9UgzKbUgelp0Zq8wOu0IKp4y6euMH8uDsiNhgeM7iPnzrIZU9bBlcCeXM1HjWQhf0TkZj
8P0mwqhMTn1/ZZ+7QV/7KDcyV8sSCt3haaRCrBWyfgXnNIHO2PO2/r+bVR3JHI9M9Acob2CgxK0p
ypIW83eErm1pHN1yfkPHtu2DRpaTQsG9O37I3+rDGwF5jem7PRbHjgB2BIT3Lys18fXC0VblPVt6
dFBt9r3UhUSr0169fK61JlX+Y+ZakOuJ4yBXxaUzyViPQvIvlJ5QBHelCs1cSo85Nd5g5K0HRlTN
az3fZ2rnRkwgs8VPE3QqmhpLwAj0zptUlKZBVZO8XSApPI1rBlMELYIhZ0lem+FvDCObM+UupMUc
ADzKkkEfNbUl/mhL5ABB7IRAmLAiGqiIqv6v5hr7VuID0D2hHYXkvisAHe1W1p/f5evssMW8NeYl
T6cHkFPsRpbI6YERaWNyf7zNVZJye5YHJ3Wr+iKZXJhNKtb1tr3ekXv6EEyH7id/GjsMLodlnRbU
0kIkORUaV1G45VayjGLT0/vBs4JPkpEHXE6Vu/U9l4XmD0C3+GSZuER9fIMnszhLbYYtxlnbRoiW
SMabwzeGQt1PNf4EuOpA6IS//z6O+SUU8VJZ2tS2rAQqTs/vGno/E2F/0yCifucnlFFNRC4rFRCM
IK0wg2RffXoR6rikYxT4I7cByjZ7fdKj8goECtuf0PwNk7TYMlDNA9OHip90y7Ur2Kdu1t/A7zoW
yr1Wsuluz9VLJRxc8bvMuIpFOw9HwfbDdNKz6sSmeC/S1H+uuxF2M2LZreu2PWtuGuC4I6VdSFeV
hKRYxl3D3Uz9VjKLdylp96+cXitiAR8JTUn3J2ElgrBX7Dpz66ZMkiEYP3XUsg3sGqCU6CuO5wZ8
RSVjcYJ7o8JHxaK/sdPylZQ7gIQpw99xqdfXxarTU3MNnlFrADp8UTIej4u9BoyOXhmum+yfZb73
5Ik6vMbKrq8EISkvNcmVPfHKqek3k7KmpqpNaWfQHozmXlUdO75w+dxStj7aut20/ry4ULrW5Rl5
R/mcSpyp+zEq6EblszfuA5D8qZFDcydOLul8V5bcxuoSI3gUaD4+KdVLX2XHAvvWPmosc5eXciTl
22Senkh3hKTlq0yv8fvQj/HZ1DCmA1bEiIUZVLpR9adFrLVu8ZQNyHKD/zecU75269dx06ILq4S4
y/GWYwwAtieVQyUlEVH7UwTy+P2nEwoYinGt8j1FMvqFUPT2cWO/nrI/m+HZ/1R2WGLJol+XH7Ga
yBLePXqmyUsrWsH7yG+mnv2xu7MtVuGE84I8gjdYWCW8TB1MnouPz/lZAo2Wp9InhFaPzyPsdGu7
TiOSZuRUz82ZWc8CKFNnNBw8f/l4jfIlEu3VJQq3cyuWdUTVqyXY7XGOuJ3N8GZAWcUwlnvxNOnI
9fi4K29AW+dsRu7hqajqOFEaCEKQTZVAqybrDKwwu80fYeCVyG4Q9/nTREEUj2MxolM4W16X9fkf
pdyG9v9Dm2EcH4GAo/Trp/n7V6pFLfw/lKl0ido5WZ867AN/YaUGhuOJbQfS/cR3ZNDvAP/OVKtc
Pv74gNVDtnoFF24JZwXvlfEFXRiu8WX21rCNI33lCGYHIr9C0LIqaxzbJ4bouaSHqZLP8sKd6qCy
64EakWz5Xe2s0r6JuEhRrMrFBg5lvQiqo4mgFs2JtQ7C0wSUzd2Ax8DBWYa6irLW4xHjTgNyivKN
2BR1un/yr7tm0UkI86ZaezW9x76bYaBbkIHGzSQsKdcSgJjzhGDqhltfIAcgQ4yhXeJ0g3JnUraU
zUIHrEiHM801e6M8bWddm8xPZ7Ta5SggOeZVi3FByPtJu2hlalQlBHkctxbJ5SNE4LUIQ9ya0u7+
TJFcrgvVLKs8jwQeE5Zaotu/LMtc4orKh2zMhEwK2j1UJ5jC8X8Ok+gbV9sKIzAERzuq82ug0fbc
hGAiRLhuwtELxU6D90KwSFVcJj28lBmzspsmeEuq4oKc6c5HJE1x7QiU8HPx1iQvTtYEu1zRmTlk
01TC/3P/HI2qYLeHXncX9CyWwWDpHRSBtyaoikN/KmWOoL6nKlX6lvKXHQ7DvbCrAHg5g5Ng1zOa
IeGqliT/4wEUJ4iUfq/njlWhCldWFInlsmglNWBNKyOQf/TuIYEjZeVaXgHTHJg8H4RazfTFpGNh
bRP/QqVVyRpITpH3Kg+Uf8WWUtble6OIJ+/3aPf/jU3BjcCa7PjGGC9k5h7mpK4OIK8CxCq0NlBM
5k+p5nZ/LwI4m76Vc+yiST10xcI3kMJVQJF05FnHulN+7iKTT+xMTpiUbiXaBfzgUkhuRMh2LN+k
84KhHRuGsePNcdgSxQU32cj9O/+Mz+jcPmeRJfDgJf2A1c4yNxhxCH54TtzoBDyLD6R7CPPhAKqg
U9YGv6bdEI8lVitU2WMH7HhC1YhC1LDfZk+34WnirHCNr/F11K6mt4QxIWTfymtEXKz/AwIy11oV
6E+Pwx1fo86sAiUlh7JZjrVENz36Mf4OsxK0neEUy/nmUTtqABVTIRH/ZEpJ+793+o3AM9BoGHm7
1WQRgs+k+TXFzLRizIVc2bYzpXgtjgypyP40pvLH+Qd6uxh7z9tMYZhlDQH54SitBUpYlTkZmeKt
15EHJevOoH9SdBRvw58QdlgCQA4x2eCEQ/gvEGrhGAPGEX4sX6Kfkwb0b6rJYN9mnIb48hQv5/P4
exJA4E1PyYwyU4zD3atOnzUmFwhwQV27b/nda1aAVwZKhvlorXFihEilrdi1aHou3R2ZokcKphu/
4f1jBp0n49ueoYVAgyldAE6iShHXujgSg/NeQiXkEBShA3jE0LTSW2U/RSzEOKM80SiydMOL+WR3
cxT6s9xr2Gezh3sdD90F1Hses/hn1dXj3lkoMRpiDFEoYpHyrdIAaJmvlhzoqGKuEvK+0GBLyGmf
I7Zm+27+c6g9xBCyosUPw94NUQAbCkumh0ZJmxwDSLR98ixkLmNReuZOIMajpOXLgu/HQV4KloqV
YecSTMdX7pTvjowFqQldeSyn8+7iSVyc2FAaC6XoyUlbKwGpwW6kv0N7p0X0gwrIlgOeJ7HSIvt2
ymDdDqshJ/aMuvG+VI2Itp/Wlrv+II1olPbsdX4ng82suWdIn/J4lZ6/YEYQYDWIx32XE0DNDeCn
CoYEWzR3aStoXdbLAoWdhnF4ys9JLDedO99GFmbWKiF3CYV7Lky5NWjMB21DUmQzJQxdhMMq8gkF
BAoWqFLFD67ZFO0t5RNju3Na5nX9EXaFZ6bIq5fRh5qp7Gip6K9Xyx5M8ir3eJc8S5Px/zx82ZU8
O/qSUcAq7c4o9uooEzJP9puKFyI+8dd8IAsberKVrG4ZdAn2K13kZDggHgQaD44TPKDT5KchwHAk
h8rNAfuxwrSqX+SQLPCo7OVtZpoqlSvmB+k5Fko7qmI+HucpFn8/8v5rrJ5FiXVb1PqxzlzxEjNr
j/zF+GCokz4/4WikpeAiDuqnZUIgxQe+xjEqiaRhTUHH+vrqiMJYjiG9p3wXD43lPd+Mjk7c7dja
NRtEBc9tyVA+Lma731KQIf1NziZtTgHH0hCdWwShU2R0IZH1qVotTAUJeKyUO/XQZZhYUo4pE0/b
vyppu0PbywJ8fW5FxbTtPA0CFeLscXYc3+RRel5tauTFvBJ26wQuImD1pTEHpXSFnb0Yyw8ndOWm
QG9Dc7o2If2HBmPEbtJNIFUq1TsXZMftrKEEKfI8dZj0jexBAvFgw+aTNUSAEII1PLdGVIMho7jM
umtFfPbTu0VX9SLCiqOEQZh/fqtciGAge/bTsJVadQTWteGAGErwz+Yn9oeLlw4r6wNvQsjzKBV4
a/gVKaiTrmFOVOaNF1ArURSB4iksJto5AA+jgT+jl8qyFFbAY3eJjX/VcWJ3siGc0QTqEQLJLpek
HCbJQxj3ci2Uq+SwM/Agqtqx6wknK+0Q8UqC/jM/s9ifjmNmmNX6lZx801x50Yfmls3D0lrJzf8h
vmpq9fkR58jIqMYwX2zG9yJbfBZJEwEQu2ljXerC8CUD9kAfyUImZ9/vTgAO3xdxk16lFD6PIxgT
qmlB21DbMEyxrOeAUV0E1iIEUn8hBF/YDd1qCU8qpHZXiH9r2Q9TzXMVCYGUOm3MPQvRaZ+RqpP+
tgEjIf7vbjZs43BR93rQ7HWumgrXcKdBionCMB/fyjyALzmKmN6RJzeX2IpPU6fbfUImP6nf66l6
DeksxbYepH+fLxVLJWtQuNrRXYBhzWJHknNTxiYNf2CPR0NZ8ubp+TU/sWSzjNAPlJfcIc0wiscG
clYyf8gljSzxm0IT8IUJlaQA3qgARZNh2h3C9Cwbykm4mHQmElc6mpFO2jnaA6oe5EqEnS7AXfr0
0Dth4Y19ouEUorROv4CEgXtayxETcK5yitMU+ZMfYUxpUXnUjcYGo2baWZs8Ybvl7aM2g3M9v6/d
ZlxoIT+mtvBMJIA0+BqHrtonZtzBXbmvgvi/79tIbFIGcaBviMjo5/5q7//k3cvpuZw89GcyvOiD
x1pw4PFoqaGpndbEPweramfuKntxBMehiLrpI+PCjhvgNBgI8PMSiYiZWC7eNE8d1Nx9x/OtxKvE
8DvNZIu4LyUrVYEk5TUhCUBjVIz7eZufBGWQdRCRTtEuGKS4qeQNthYJ3HdXXh1XduEpbCFB8HDJ
Xv+/KzEc+lUA3zP5hs6xfmPuDC3tuLutR87fzdlJue7zRYa7Pf9OTXuRYlS+NBsnAZvgeyxnYO2u
/jYudDyfCO681y27Tsv/vuqDfm95IqklZq1i9YOfVhbbltJEDggvQc56F+0c+jVJCMtdM6JEWzgP
ku7gjWQdBcMrjq6SzJFkMNoyguYRv+R/LtqvZN+Dzl+zi9quLt9TKBy3CqptBokuP9QbNh3XblC8
dKMoa54SFkztnyNFyrI+TrpwLAXwJyNRbuG1/UJltsHVBdtaCtZPI9DErN8VN9asgOa6wc9xxQtj
2Bs3K+LERz2r40xrlTGQuithGPp29+AP2P5xmP1kCea1cjmH82Z5AFO7vallbAoAsUwtAUdh1eGJ
8XLX/eionZTul2qzosPPC8XUaXCNPeWPWBrDDg3+AlZGQ/0+RGPpgUvTX5oj52Ws4H0Cq5KFqFU7
eIYHCKTaesXoBIu1Gnw0t57kKEUTPP9G4gWuqz5JNjWEguknU3QIFHJxVQPEBq8vMGJDDGggvaci
E7JJwP1AQfSaWwdZ7xowfh2EbqcmUsWUoFpjzbOXTeJmDDJ5v8Qa3vk71OA8V6arEVY3QUNsjEFs
UH8wTUKSWUKUjkIQk6FLoKZLpFZ5bcj12cXIjJ1PfBCEw2TkHu6TlKy/VuJ+QQBnan8gpxrhYCW9
lnhO3ny4q5fjX7dhok3H6PSOHi+WgH62nzK+m0hT25S+c6fz49n6Bwj+ec5BQNB74jQjc9utWVYO
1W7249vxmYwG+7KoVOq+I4p0QV2FkpLrOf6Menl2zU1rFKvh++ogW+/VJJgVf2pKnGjDedGBasfW
HFtxVnfrxmsmC7JzEcrllcicP7fwa2IslSCSRRUdVsR95vCnQniZuwUZEZo9AMeQsnUKLZ+H9Oe/
ocCBNIHR1crNkUcpwXDJtwK+Pwcrj+34+b36fdSsKgIfqWE7WNppbdeWNHFvpO0g1NXqNTFJxDz4
5GAMuLRJ+vT7rGpr6xv4gOSiaSbU5W9L7U4vN2Q0N8XRtmk+ePJwslrq+rhbcc78dYo22+d+RVx8
O5OQTKIOu011WjTCi4I7wCSmMjCG3flk1FUCIPe9ztYuym1GCdla6Nf67E28KUDbKTPrSMav+2bB
+1r+aWNJvnZgw8W2J2jvzW9prWB0oSjUKWoiukQ8YwrivQgUvr0n0TCi1Uont9BE/RJAYJnzgAUx
SoXyr/ZuR20uBLXevHQJ5fpQNEfoosIhskbnS1XbJm3surMAJu1pK0xrE04i75qdyv8Y8l4j38eb
zRgZoI+cmgHkDVO0FbTO/66Q/frw7tdQ0zGl8egtRSw0Pl1UHWD1WHfOdAiHoR0HeMVBpTeMEra7
+jgxDmg9EHTR5zpT3bIFrcb3mh85CfTwaV8tE5MPBdeNMrcsm0KvY9+MUUP6ZxPKO2PcnokAXrWI
bGRcwB4QJuV0d8DDY9dtR1N8V3dN2oMD5teU7HJA8N+Q5nOlmVJEZGv5P4B5wjqD8YmClk+eFb6s
UcurwLrmlcOCL+MXBNpd1RGqlfJhYxeCsnjF6kQyrW7MKm0fsbhxD079fo+Gf/acchkXksG6AK/f
b98U0s1RWbnEjMl78avEK0yf1A0v4t21MImZ4XiVIIFwg7lzO3WTyFu+FVfh06RSrXp5iM3LBpxy
1MyML+jvs++OlgK4b3/vDAvYo3MlNhQaFr+g/QP0GyJJv6CantR62dLA3WyJ2qs3EcHxth+D7q7a
JcJiNwfJmGQXjyWLy+6DuYJdpio5LBOe2rl0cAGOyFAYC1k3NQQCaVdoNWEgbrUd+tINvBaaTUIB
SsJ5oUcHKAc68fwgv75flpDeYYpiVeZGhnEmjo5LTZNY7ZvYCAMxcs2l1FaFliqXN0U2wd5seeJs
PNiiSPy/YzqEMvx/wJ11YoWJgZL/q8k1e0SzpwAxkjDL7hHfrYKCs5LCP6HwjSDLMKROX8E/TdMi
RVqXpQQdMXhKgIiWLsEBelEEC7e7cR3BIk83t2OBMX02BwxiUCE9nSyzulRRoZ5O83hRTBdvM0+R
bR0RwA1L14IKSC9m+Joy6cxCELhh1kbGIQ+NrJYwJCUCXxRczACnYEO7JUz36sjxlByu2BqPKhKK
kyf7XVNIJfXbXp2i0xoOnfAQsLBwkAgMO9L+yIV7RZCmgjjCfI+0/MW1MyA6jhuhb2BmEkpEJcTW
a+rCu8keLnMOqBqWk8vu8hVZY4ZcA2Grm6UgVxum4Tj9nsi/dgiLskP/ZbjgGbmO6G6b2fPIw88E
kprXoVOv+YdZLdjS57iv1K0KFXCJTqsLrPFW77EVKA8puAc35Ig9Ocll21ImVkBi35RTy40SNL2p
emW5q68OxYbxLQnSNFVn29SdddZhXrfPdq0DI76Y9r6oxNU1/bMOzOvdy+IiAeCe5MYcPOvUmZ/e
OYdsY+wa9bn+aP/M+DkJrBDB/ZaJCQkGneoabAWt/v8nOvWJSWVS/FDSSbcaCyIsvR0S/s+9Eg0O
c0ETe7PfsK+LwmSMaZVJQ0utB0YqYF/iYHrDPKblqqRjRxlBhCSdw93Z9os3+9cPs1LIYb2bcoP+
+Kn2LZ79VblnRVOZGNTwqIU+tdRvrLFsPYV3EdsI/N/CLa0gCOMbC8AmDtkuLR8OcXFShJfhSDPE
USy5XZh1bcC5Q7TqE+RtxVcZb0ubekNNbp5ThVbJ92Q/xOQBW6FwZjetrljDJ+cO2oU7kw3dC1Do
eur4fK9L2gn6eY+dIPyLddDJCelv2m0qhmFQ93ES8UtMKnhAiVlbuyxVQw6iecGVlrZ7MOwGE523
tO4bBB1fvnfjZYrdzAiyfDdagG5EkiW4wf82XcxeECBuhMOv3fi0N6PkYTKw1FZvY7if/KgH4Vk8
UFFi4O6FSijxYjMA0+HQDnJWfxKbBs8y/LGsgN27VGS/qXLWSwDn8GQ2TyH93cEG0YV3JoIRugXq
tBQlO51dTqBKY6f8empN0Jg9t9VbURGiF6xpju67hPzsj/33jzb/8dw7rBv73oG5S+TjyvmuzIKx
7Bi4qThGZOBYrk7kjRO34clcLV1cs4sLJuXub3YoNl3hlv5z2RKGiGljnZM1uXeFcYaayvKQKGlP
HUGAfdn/SSCbrKzVilRRx3mAt9hp73zPKQhEb5d5HwHtmek1S+mrn3NBCOubS6ECL9FbzHmQwUid
FZeuZAZ96PjeKaPV2rSCNRZLcTLs/RNWKSn98Fr1p6BhHrEt/0j1tWTdd1lbFemS4e+XdPtOWqRK
zBrFS8wWBaPtlURShXj0KLhixO0Wz4kEPvFq1pcJxCj0G5wVli/sN0djtj7x/um+ZXRzxzts50B/
cT8q6A+e2hQAWtr+h4KiNcmB8QKu4zrfn41eRxjdl/+sR4HHzHlxy/t8vxUTL7KRj+ZhgA7SvZCN
H5SOIrR61xz/GdSpyPUIuSlL8FJ6iwaGXeu6ZN39iBhsi8OSgnVJvRJuhzf91IB12fpuQgApHAu9
WuBVLocp13cTe0HeSmZGGpak/nuIjelZairE0jgEqhucWv2K+RbeNky+TbkdxLVwbeiI3LFgkZbO
PtS/1XI4xgzNEAuw3k7Qu3+n9VWP6WTXEbpxTTIltMpfddt50oKpM51cXugWiUhY/BULwJlGvDfF
F4dIH5s4und4mFr5F+CBata3tVCg+a+FllDB6FWgTnQBomKjuoipgxQQi/0Jup7LgsOzCd2PDbzo
sxGqPi4lmtYXvDHDqcL+8XLCFPiFKCFUicKV71VbSrsLxRxSu3cy8RIZdmAtT4BISmUAL1ug7eO0
KQEATGAQADaD5zyn/X2XbuOzgAsWa/QPETQKZfLTYcaMl442UBoO4EUtbEZwxutV1hQiMZlBVPPA
8Hd6aPiTS1X1le1o3/rSsisS5/zustbEgg6Kl0ulTTxAhabL2nGB57BGlwWSks9QO93PG4YZwI9e
ZGv1yUBglul3rmXsErysY/6opv23X8L8CP6NJwLpV5U3hGZ6JtE6vLd0aAGVdaRfhkLBn7ORakjx
fV19EQKo1MgjPvRbReXmueZvqjCgTQprdJqpd1IAjzDiskuhFGzayiJBQH/WpPEWMimo2hShe2xO
8veLfjFKFvI8PBdsSzXiSBkJ/OAeehzj99zGRqdYG6AzNb3nMNS/BAJOUub82NLb6v9n0Rgesw+g
5oisHsgTS/mFwGpcmgjIc5xjn2SaCki1Axj5PnG4krvFCmdneHMr7QhoNk66BUOejSDrSdkKkuk0
3dtLwwsQGmmU0p5IuueWgWvDXGK6/HBuX6VUt7Re7Par6/bcjVO/R6ACEigVevvf+UusSCBxeguS
ZC3WmI3Ufk8zXPC2ux0StGhF6HSOEi4lxRg35Jjn4kvaz22C6sTCuoRbpVXBwxFnd5wD4l9D8wJF
/uC8C1Te0TrMjkfnDbrif8gAK4Y80VxZ3DHP2c7PsANeT9xTFEf8o0jO7/zvyLB8GWF4hXWNhK/A
4pDM88b66GZn/ImzvhIc4PSU/Fy7EhhA3qp9Ou1XVQFP/K//a+JQg2aRkSpAyvK+/8qZsFMHLcpn
XIWxnEBf+2osu8x9uQLrplhv5zoymPGP4CxYKcF8kqKj+18PeRmvRVNPS805EbckSRYjCKxr3Szu
CGLJjvdHjJZ+ykVhd5jh5PwJ8de0CDLtgzN/YfFyydVCQLE6f3qhSUobRwSulBTqNafwuht6U1G5
+P14iNVQ1NBHlghLZ8WU01ffzdDbCECItTMpx+6yzNy0OPdexNqg8EIZjKTocaNNxw1T389YxIwg
tLoAZ0j/e61DtblnT+Utz7HvMTnSxG7LAud4pX7lrV1dvFlri4+YbZirzlv+XRhshTt1hr92pwBz
SBzogvxG60h0giV8IDjjWqExp6Z0lSaY+sLY5EP8BP0Jo0MfFM0pX6Os4X6XflJZDyCy6d3Pye4U
Zamjc07OaaupKcfVtC8NRZLTHVwR3Ejvvptl/Hg/eEp9kkA5XLvMlW/MAYJw3GmO0HscGOKeN5zJ
5Ncr6wGBDS96JwvvtH4JEMSIfU6r0f3D1Dz4Eyw4R924hBhxvOQK6Qb1brNQZ5nlq5kQakeBaDUQ
0KjEnROCMsmX2emH6tfhtIARn2ZzGNF9K3jReJvgtCwQVkAhwaTx6qCe37PzK4DZiWvGIag5G8rL
AnHyblOq5+721/V9eo1sbpxhPsIFT0Ec50CLVhMFLx1kcx3GB6ZzZYosHEPi+E3EaFiApIGHr42q
6KthSi8GH4g1cPmp11CrAj+bnGw2+5CCa48Iq1sCyLAUkhQx2PldOJEa+YVbLk/yNHfGFyEhmdXg
SrhHRcFSJOPqm6mHGjZ8Zyllb7f1bzlUJ0pU0t8XwVxNDNhvWaGRUnPe5WXk8U04D9dgm/uJ1s//
sCMdXQtwtBsNI0OaNj5akrSuSgnTSOzjyzryPMqpiKHKFAhxr8LZB5C7lsjsDY0U4cp3sJGcXQJ1
Ua5lFlsVPY4iewmDu/KLvWGSEKFo1FYcn9r4K1t25zBbR3MgEXhQBxnDd2EMJMrTj1ZPdaWZzH+r
Dp4clG5AbpEB0m/rcANQ4DAi8CKD16+WH9/SDMbliqJFrh9vFGZcbsK5NU8ipPIrIDLPkfxChZvW
axZSvR33zGf3Jur5njAIeCtxNGs/DnL9arw6mdK77rJRQlPnm8zmIH+EfFqC5e7emCPOAwWvLp9b
mnUL4JaRBHIVkYcIvJctHHPqjV0clUSnjIwMs2PwAWHRSbNKqC0TjurSuHCwltiuuxVV4QOCWqTP
FbLXJkha7ef+tEUVtvYEUm7PrWElwbA/YBOokk90XYbthk4qqQoa/NhkzHIQ+QU94CS2tQJm+U3i
WPNZTnGup1KqbS5ZlTMvHK9HmTWi3gS5W9d/WonH+f/xYsMzwfNBgqid2OqiWeztRBHCgW6DYJr+
09aVe13zTcH1rzsCu3/R8pb35KApap8FTZcfSC/C90BuTjQn2/xhH4t9Vyf086F0lGz4VqvcSV8q
0O07nc/at+imBD84uB+MpLfjylpFLE24UXemUbDBkr/ltvVCWZvK6ALXHLt0aJlMHp6vdjxOQ8x9
F48tReVw4w2qj4TjG2lktF3F1+fh52VplUG8/Ph6AKcTEuujuoCmfvso+XbhFfe32LuNNPf74E7/
BM+pa5iS1TlOf93SyX9DTXfEw0+fx5vXW9kp1Y57cE7Ky+OVuzKKwCWBY3OwFjz7+AHbgd3yk94H
eV/DQLnC+du5zUjAd5AxH6mjRpZg/wZDqS+T181DtVDyIse54YnXAahIITNHNAz7xGYWmFAa4aaX
LWTuT8hIx6fxinANWWyYwX869GAQooSyatSxZVmnBMgP9MHN/tkYnmXERqbq5BqoM9aOFwBABZKu
Hcv5EQ3jQJUlCC+Sl9HdGuePokQvhFwmclHLTmlERItIrnknneQ6qRlLa1JBA2m9T1bd09ZRiox/
v2guYSwnWCcJ0m0VbcYNEnMGpDUseCu183Za6k0EaSpxcbawdck3VGF9IW+okw9boz+5+g3tniG2
hwlPuIMsHYZHtgCI2nNEXtPWNIyRfTz4gM71bIbE5I/GvCWaLXHTbw9e8cVLptzd6Q4mGIHjw/xl
7AiQ8CXlOybBBUyLaKLvAJ1l7ma7eLm4r4SqEPapxCWiD5TGDeGI4j6sVU1p3CivZ4jyuvPHPF21
SUFJjIfNfPTbmJCq3hEhM12MtJu5FwKwaHzGbAHNjn+8bqSOYkOd2aHtwy5tz8d+puEXr72KhSAj
a4rum3CeBz6yIj1eqzEzX4El3QQQL67LEoeHntxfGh0yGLqCWwkCNUuCtNQp5whss6rX4Aqsy0Li
HiRrNYAhof5F3Mml531EH5vWlTT6Sk8f5aVntN0mIKV9kdGM68D5JSyWVI3PU2Kz1pGtl8/uTBlz
JL4H/v3M4otUbYSc1eU/cbObAFAoRXa8p1NgCjehFHs7Nc1MMI2LIGNfpAwy6wbds36dKni3whxS
tTCwQ8CYEOGfRZg/Ppc46Eo6KUO7TItpHuu3kf/BYWKsu1TnjhYbsy9a3g2aIl50CAevJ9mlnGdX
Ix83rVBjB1M714hkFfY9qc4AHTBsVTA6zz8R7gHvoc+qxsUpzAtl0EnmB3Ikvv1TFnO2RvL1LOmL
4ouO9arHORIZ6uBrjACdRtWAEeVATZ7hMILWXizvY3+nETLealVrwhDvIhKV/EDSviI8MX12JEqp
+8xn0QsZTZF9kcStkyKgYpT0mtMwVrPN5WxsvaH1EYGTlFn2oQwQ1cQiSiekX6HZQC8hsde+eo2K
4v9pSf6n3jF6CgbQ/bEaNUJEb4maj6EOCQKpq2aW7yTmvfyqy8Ssheq7CqBGbfXl2U6IhioYbfp2
Ejgz10uMLbY1fut2CqTroo23sPCdtAOg/psIqeek71qTDhx1SPVVIJ1ScI/lEqlw0auqN0ypxHmc
fhAS1uf83so5kEerdBFQw6Qcq2OqwoFpOoIjEhR3bED7oQRG8oYTNVImdgUSWx3dC8mr4iQiCKc1
k9hviFn1LUE5Lf4mJyWNlO0pL/tKVLSMRw9grNEaLELY0y94ysvqor7JXabf4rlHHq0ukTBHwYAL
yPi2Jr93SJ4OuCxMTF3jJyscwHZArbn+wbysZcufHO0Q0bg0ReSvAZSn611AKr1ZK9uRT6rZEJwn
Af/+OQ0imbm8uiZxSUBCyJYouF3Je3NfQXWxZA+MRvAtvMKTuS/DIssKsM1pFOhvzeTRBhu3TIHi
Ja9dCM1WBSInCAXvSyKxQCjeYvu/ToxCwYbt85eauUs6EiH8lJRCr/BhCjhcE7P1c8sasWkxo+bc
SAI40Pb3UqAc7XbbtxsvuAMJEXUFpY6ESGEcJGulmgK/sxzxkIa2ESTfZLnMbV611/Fu0/qov8Px
5oZkIlmWeuEpxvONxo8NCIIerX2cz/psSx+HT46nNj26UYK6Toq8y7Zi+mav35bqFmf+GBzv2Rmj
h+miMYdvFn9s7DR4jS9T86r1SLvT0sGkbVryB4dGyXjVb3fFkv6dSRumwa2d4ob7B2U5eAsFQW0F
fnYljVY3HUWry1r0PzvaEfxWrv2K1bh1IqmUsyTTkVOoiYu3ONMIfkSsDQWYqUUndAHoTUBzEdeX
M5k7z/QzLuyQFIkBoiHNz12g+zqPmueSGIPSxl9VSsZ4kRG4fURLkrjIH1VfuOuJ+D8YPAVUAzo4
X2tRS2Xgt8pN0kZk1rgPDs7uONS3n25P1o3k10uWLb+CFVmJXeQlRdt/MqwPvbyzxvQH9qjc7BYt
8mSqD4Sx7Cx4y/VEPjnDYG1ug374u8HS5wMiKz551PMjCL47YU9FahEOMwZ2SEirEzXNoljAfzfw
nBQQG7yGTrisxRwD7yOlvczCa8oG+6bakB+eXgwkTxCnB9ibYMZZ7GVg1svg4MdX6lj/VG8mx6w9
pe7Ly8Y1baxGBmaOeMSd3tfb020FRclT1yJvUUhG/tFoCKakdyrUqH51nrXf/g6ZtrVecfammMJv
rB020/u92L34Jjvf0sX92OkC+HHOWTDMykbAYhoJyEuSS0O9D/VF1b5GA9R7qprRsGiEPzrfSNQ8
snEgxgaujSjPD8dmTBBgaK4FZVPR+Gfg+fNp4KgxSYXswPpq0L2KMp6kRrJBI4UgAXRGQ3yb0p2u
OSpxCZ6FyOiPtrWAo6w/UYLTb72azZT+M8lufkb9d6mSL0vIzs8e2xK78U94DD5AY/cgdnVxS5Cg
OuDeV+ETST2G50kROp62WP2lM2aIWainerYYnW05TNg2iz40JfgwWlKwd7CwMqJ0l0Mo6B9PlqZV
e7KmWWUAsp8jVUxBIhWumfmu7c7bp7SMexYNlZV6W3Er7GfwtFoCuJ2l2gzSAj8EbNvEZ1XGWMet
K/ZmiC3QxwkjTOnRgAIWG0eDvW+ttUJ/XTuN/d6Wp4zBP6qo/+XQAe3tUK/6SQUCnajhK3KYy/YN
2320/iD4Cv6yBDiBBGD0bbJQm0qJGVqUvbWKE+ctELCFRCZTihZbBlYtMITMmYPwErdJMr11gX73
6OXqC2bPGNQ8RQiogP5wYYpeP/awy3+gCEABqZSFoCRyPRAXtbpnnHMks1WcSxFvPuu3rlSa6vtu
da/G7PWMd8IlI1g9PFTBkx2cWFM7Z0dXgFJvqcW6dHTxudaRGJynHPsh+WDlfh8usJ7W8fiNDLgA
2Dgv9EjfaA3QHRdk+7GJSJlhKlR5Xln4pDuFLLGLFXFYwaixGc+6to1ucT6vYf5jBMSVuhNoPgu0
XVbome50TA/d0FIjacfyvqxmpZuw3SrQ6HGnyf87OwC8Q8GWmAi6dnms5QtaMbDQNv+Ze/mh9qa3
3b+VnFrbyp9yd7kRnqB10U/M8dsA6UC7j3Bt7IZtdehY6jT6jOMC1CvFvxgXCTEIp1vZ8vpfgoTy
3kPAYD57paY27C0jddnQ+WiKlE7cZVi2hRgWl4dayZF6rvQbRLziXIU2RoIybhABTcT0808wrQFO
h+SApN0gp2z6Zn7Sz6sBujtfq6cfjHuIBHWqR4ZFS8sG9HKHb0dtFH/pHELVMhCabeQWzkK0XmrG
aqkMdzZ4YT4TqvEvtnu1TJXJa2UfDf5qmBtfTrCbiZ+Zk86SAJS0iQ4FkfFIbJ1p20A9kBS8GnXP
v7e4B3oExkw4H+UXRzv6m+3sXrNm3+8cpGGdhS3osTl0AB/CcM1/9RjJjZ0+NH4hqo1iFSPqtE06
isAbJClTqAlpeJmSRXw72Z2LAXv3OddSgJR5N1+U6L+6ITxxpRzxMWZ8jN2DRL8OxsDYRscnR6J6
GD0AUrdNdNkNfFueistHZdUqoJYNZ7SoND+86R79MPbgD9BHM0g/iu8Dis60+FNbL3Wg7GQwYBM9
u+fzkWIshHFR1WDllNM5sMLFbRnbxharq9ru9GiejRokQYKIFWVNw4T3reZvs7WKLWYu42CeEgpB
VIq13/I/rFM8VgG7ePw0fvcM2lVJ/xYGZHCtTTOvH7B/SOJReflPT/Wdr92YWUp+611wa6BbLzO4
yd1TuJ/SAmBaXBrb/wHTaWljJPfvcCzd2Y7mTw07d+vdxHB+eWs70jA6E7Gd6dDgORMCJB0QOpqs
uniCVQWeH4HN9rfBB7/oMYZWheGCLwwWVW/K9M0lhGKyLBYQ/nqfVnEe7x+aingtkAX5sLAkG2CQ
31v6IdIY44ubtwG0lC1994Ab6BJ27XteWmyBOSRWQUnqErYPkPjXfQ2wNfw+MBEYyeISHQSvSkNs
6fgDx0QakLLZmrR18edUznVfsDwAYZZs9k8DhgmoJ7nVwb8wRgCJ5wdSUpfpv7SfsxYyE9yX/iZV
2/DxCzspEEMd7k91l/G/P4dowheuZj4rS34dIwRrctOGq//qQNlmcqSmtY6OuWFLHFrUc/FIn+5H
zQTw1RarTwsc6zJ126PTDxlfUSfD/g/xWAxtXV/laaymctniTxINRS6wOzVXycDyfnCscsnx1Vuz
Ol1f0npQD4SJCtSZSbg9VMEuEj7dSdVHscCJf/4sbyzVq0sSvjrZtvlyMTsUBa3+VoGfsRcHXL7w
oNQ4vh495edSZgsVMzoacyVYhS9yo2SMOXCaPqW05z5XkghXBRLTWGLhS15+obWrLPGhZG84fDYu
PrIQkchB7VGgbR2+3sWr5c3OEwXzvtOth4dgGnRByi9+n7Ni7ZCYoyMHth0rs1y1SY91Jx3dsJMu
we1kv8rUZ9D2U7X+CChHdHsVbY5Md7Bc93U78NjUHQzT+5WtgWfSI7ulZTuNF/ZdziSrpNJS9YPW
kceujAC1eRd/h6IJHglkLGYs1p/ew7nzHfBzzFtayRFm5Pb3nSsIhDxuWCd05ns9shn23XRm28NV
Ki4ezS2h9REi0qLbq7IW6egMa6OQkX37sLueYkLL/WD0f9ZyKJ9sEQ54Lgkgtl2a3XpqQ/y4LdTP
OKFb4f+z0WjBNljP3S7QwQ9AJGq/NIjx28HMr1XrzH/AtUP4mLUVRaMgPPklGFEeBzZcr4qHombe
Q6FYssjI1GnZn+tDE3yHQhm/ADcdBRU+mOcPYZrAnSGJIHmkugCI4B292exhrKuW+jm1/fyLuIbR
eyaz5kPeHiDRULzoR9fW7R0D2fEQkMwOANS2fXzc88gJJOeh+/3xjSl7xprvMhL5mV0RKSqcBBUQ
BzhtzyXxfSQOA9FyJ5e/qjImMJiN8GzJZ7RH+qTC/KCodLWtFM21JUns7yTknZALpPjTJoQRbZcF
TwbGdFZF/in+1kJXBZKousraRhXw0rUCE3p7OaZ0j4Mt9suuPIq1wfagt29CgQtItbgxq1NZEzPa
gNFXz6PWwVxaO/1pFjIpqK5kShO2Wkscw27HAtFyJYUGF6Qq0uecGYfj7rbcz9EkH0iJdkvsKS7C
i+2brFOHKlURxYRNwLbTkbZyS22NQuSZy6Tr51Af9/D7lqB+BYEflO6IIB9Euq1oGEIXg9bWZ//6
Y+svcIDkPbhWUdqvH3S1Jw+o7dfhrni2dlGlaAA4pyBPoUTLC6AkBHmdPxTyPjsiARu1aAOTKzrh
se2zFFrvU/PUChwTJn+INgzPRjY/VstbkEv4PO+lnu40waarpG/s+Pj+VyY//JXLD9kNMJIOjpHS
yPbZEDPEUV86RJeVq1jCvOhtjqIcxtXjUcb0i38OzAx/8mtKSYPjcSi3aWI6AlXoi/5SXJEBZduv
cvB2GvjAPj0a45CcZzBNoOgh/zhWBpYFyaUgslVVD+wqGMPJIliWaNOFy0FlPfni04AuTqhq0sK+
L+QhZds76/arF1YEjaZ3KY42Jm9+cEIqv1UniCzUhoAaO9ZmRD9jqPIqj+TNBLcxnUNOK5G4naE0
GpZH7OxTA8q3iJHRZuJ51PA+RxJjy2buDhPCxE1Bi1yeytoBiVB+QB9XiOAO7pG2MGdu2OQGzXzv
Zk1Z3ewBagj0G+mXL6JG3bzf2PAMKPwfEx3csTvvm81i7I17l0bARImwxTGvUQ3HhY8kKC+IiCOZ
YlUZOHauLGvXWWS4JzTOSXSLeQkz5GzlAw4a2y8kqHs3aPQ0wDJKBNQnluLf35KVzlPcPvjWdpFv
c4H9d2211Y5I6D/uA0eMP28b2e8r4YaOOZO1PaHLJiBJlvCleERdNyRIpXO4GnrFmB6VT89HEAr0
3xzG9Y7M2udCcFed2RvTppgynhgceCzQ6TaDBqHnv5+0oatjAnUenmSgY2+fe8xMgXYqtQgmDWvE
py/gVqXwCuJq3Rq1ivVZm8xcFCOTJo2l8tuNX3tjgSXmpe/0Azf0+3bkrA8R/V59Z5mtAcDK5Atx
V1VeWSgJm4dK8GkRTseICACc+jSmDD1k1ZYYE4WDpkVSYCFKZhU/uC4EBB26xlx3kiI7amhxa8lr
8mL3nazjHt8uI7REsOtWTeJsJlPJ7ypmKzM+gFZAaRWDOdCKcSa+CdsJcOGnXknbmnrQa9H2L8BM
x2UhRnrFUWwqrjKy2KLCmarW1Drkvq4gU7N0Jb/oXSCjWS3Xixct381kZa1tsU+8Uy1m2ZNoRCVs
eUczlvoaX2012s6gAdzX0fHZcdpJMSreKpvdvyKw1gxi6fCGoDfSJ3SBIXFmay7LfCnEB+RlER5x
wYgCTFk69Tn/6FFShtuM6GKOyVmDvfE+rCV7XK9+DPljE9XSOdCjWGgjQYG6L2U7b2Dch+wxmZCG
EHovFMuwyyh9ODG/mGNMFMgyHRRix8Lct6o23+MtKVYm8WYvEDzf7EFCaaoBWHiL0PMmJ1vRnm4e
BWlUHYLWqu2IGUg6SeEC/0cKLdd5Kbi3qrsASppwvur2IT4ZTxFxt/uOuVpYMbf/tKWHGdK9haZz
Gn8IrgBkNL2CPwlYoP4dSs7fQjnz/DABQ6DmN0wdgfLvWjOwgX1opzlooami0+Yxr3qMnOFS1pSN
SAVlVGRZ/cSj10r2Y0Q9sPvmmnfAdCLjnYp+zvD0pKFC51F51INu8M0QTuZKiZo5FT8G5ufYkDOk
6tPZp4arsFEiqMwXftDiI4UtIUZGdeIZvx/cdGSqNYlYc+nFoCz/+PSYGBI2HtKlQqaDnxdwRQUp
gMTsPQR0d1codh1vqPgA8z5nzr+9882Ea3WTlVhW53R+9rAOLvzICT4ZjTDO78CAeL8mj7H8f0/m
dCWFPxzptvwLlf/DtN1pI23zu7QZp7UAwU+OCc+8dC0k0p9CHuW8BQZYN8aYrd8kTbdy1xQpzNvr
8XkNJ/vcwitffz+gq9PTx1ELhkwsF0biY5kb0oclMpBTjdMRDmk6JqNCvPfpI+zO0todTPNZv1qD
dDlIYler1taTxNsqUONtgsytTvD71E+lk9K5Yt56ODi+giksiwgr9Xhbu/7W1khl8mnosnGbTtoE
hcBAccCrvQkXko9f4gyk8IpvwkLl3zSVG67CQ30ZzoLAEw6CetfVhCfsdiNCofB9oNbfmPGpArF8
ckROOxU1HZAL5wLf88vaK1BMvHjGaU8Idcq2Th7W5jHWgM7+2aBMYOUjywWf/L5IzHC0uMFBEvqo
14Px+Tny+HORRuvawHO2Md93HL2pP6YCIQ+FYi9ezhFA7+eJAdiq3Hb8ZekqhV/2sTJwPepAhpqr
avR6W1XmDbNufVYN3eEkMg+5P9p9waunsXbPpLBDt0eK076vO+TFiKmRhZyxOayGlBN3/X7RkX1Y
JdXFNmB8lpqYRlYSYw2IGA/4xzyNDgpZV/HcWssBbzGeX+ZFpTLA273yEvNxN4G8cw7yTRj43w9m
YMGYMHRDUCWNYSgxR2FKbFChdv+pCMvTjNI77Tf+LWtYcGhB6NqB+Oo0Ll/1etnRP7LnEFz+Ja0h
7bVNvNHuNBMJWLSyCxhEQwdPx4UqwjmvzkZSe4P9A+8oXGm2Ebnsh7q24p4xzKpKSdR8kB/UIUBK
5faMFPYTLu9/+E6qYdBNMendA6mbkeYpwJPEZlo60av2KOrxeKcMvxERElaRr7WydVl4ki+Toevp
xgBfwQia0YKOrpazTNCZQhW6HfEY+PA8jP+43P/A/hGGmv0/2RuhYOgDj/uDjlwHA71XT53Ol1YA
BiaAkPJ1lUun+NHvr9SOmjeoCTGzeue3+lKj2mZOqNwtjbRvrWPHufJFPIrN7of4BbhnBpIOWZ9N
NFjA6VrejJj5pcmCtOwGTvK7i4vnDoHRkj5oankBKd8gjAIwJGK9sjXfZ1kPfoViid4jY4dr1UuM
yTj7fBeLUsZngbtoMJo82kN/8rrCJ+CMKG335qbUPI5w2WmSuxv7esjDjSL2ATtC7TOrAwovBz0t
SdwoLYmS06woJ/7ShHWgnafvo11LqEPCOlOBCOXBbRpoj54Tjy4BbSYx9m+QsGZ3Dmt0LE/y+FRs
sWh83luzlZaU36SlAUEicC78cEx+zmFyLyDl4UIr1Le1pT23gK7N7HYFpuSKnyj8/BxyyB2euANr
iZ6/vYLbpRzDpR26kKDQtxekQs7mBhv2fauSGravAav9BXfOx5QDOjjFv4QodrLUvIs1L0gveBsL
mqz7k+x5Dtt44YCw+9R6oiNy7RMadtkxKjryoV0t1dY7ULPNf4/NreVN1tn0+otb17TvG2W+t9Zn
MdDLvjj1oHh3apBgbsCi/S4BJeW5iqhc0DpU6AzKkYVyOLN87zIvQFAgASCsV61DP+gF2xnzp3wI
S+RB3N/qfl2623MF/JXK1T38aBcfWukuUvGEnsw2Uba6DRxkkSL41JPnL1nlnEBwWPxcRkFVZZEe
D11Of/8O4tGYJPJyRpq9bnzxh7RSwqTZ46Ui4s103nKT8lL/jQVxU0/C+XgQmwyLxfG4pXg4i2zT
FycGqcbrT3FyGTYHUYMN9HxKY4R4/g17YNaUlzvYK/pxNC+a1BONH7wWgQiER76iZCEDeWY9/wWO
2iZhaNlGMU+TCT1HxNlWjQw7/ZfAbpD0oxU6gtFPzg24OkxtjGsNc37jNveY7iI26BqajFOYHT8W
eswGofLK8h5LYIn6HXZC8dvqqJifRGIm4gDPAKOE+EybQH24oTOxLKCiKwPdVDKcx1bOLOb/OupO
JGYL43ujNaF9oWWmoHHJ/BxY1Fw2SiSbRxgXMP5qJIt2sUO7Zfe+5yuAOZWwpnuKS+DcoyAJxQ2b
HbIb154hUDLWcHlnzkwxhk7M95O6xdUhw5HUq/OwlruhI/UGLWyaODfbtIFsMjTfdbKQRyMnTt1Y
ubVYdUKoizeHHCgbV/yD6qNDyRG0KtN1jJP866Q5LoSHIzgbGFyY3J+y3daWsBWyQLLr/1JQJTuB
rWVXcJB+XXUWV7Bng3F+gQ7OsUSxq1A++9IIUasI5hzZ5xMRSf6xvWhGXsXVgypGwRfsbnIPKmfA
CCuquxM4bf96a8m122WTpzsCx/ixNgCBCI0JlRxhfT0NbnfqeLiwvsasuExfxbFDRWUh/1m5lOc8
dS4YZ3PcVzhlmOAhGWJNQs6Wz6T9BV+ZUUzdvxGma0V4rlrPzKubts/ox638YIr+QSkEi+mQS8GS
Lnp8qABehRn6FIGK9pDwW4bDescL3MSKaLEkYYrTzp3F4YIfTdM3m6fSIeqdREfreaR/pn9fuZb0
hwjiJhZwinY7hWQ7XuG+0Hj1gXhSg6RldiUyOdeqBDwHVzUGTQ5P8ZvDp7ipAW446bisH4wecqgg
Qd9PGMQalL5o0Pf0ZDfCCGXsiFJ6FRa7gig1QNTNz9nsmQVkiAmblO/qVFLLIC13gXvJZ89XwnS9
SkcH6eQDACZl9juH9VAtWtl4YZ4zGz8ABPCcn7sVUifDZTbwsEyaEnXReCoAaDOzlA10sOS9SU9w
oczhkdU0cnVFRKjsE3oXHU7cjjtWcLTkFszFY+s5dQLQFnbzdeikeYyIqYYp3VVjVpV4ehb/vqwF
Fba2oSiKEohxSZDlUUCRcTTQzbUq4cNRoXrpREsNJ4FRd9m9LYYIaELOaP/Y6u7PQpg3LpRJ6EzQ
XdFnircH64d9Lt0ey6c4O2SzPB9oPAButqAMhZ9z3NiymQT8KpjfvULnSgIHFG+Xgn6zHYwAlFm0
QZTz76s6ki7uQqBEFfDI7AXMia4LHfoA+2oF8N41or2ykfnotzLcBqtcFNBSp+Z7KNHw2FBdt2nm
MTK+DUo2E0LqSx1H0bUa37VlU6pvpoDMveIulsMX7FxrZqgzpTJ+MRr7HCvBydwuZ9ioYy/v3pHS
B8qLjozLSdPeGhC8jWj2hZ7gSuGMvpyB8RB7OZpMcnQYM+WUed6jaXfL4EJ/Go5oszLB+61+m4bc
luG9Br7L8daO0LIq2lbpwM3wczrT0aqfYN2RBvt0YfKah0LrY4Kh4WHDVLEJjGjW/GZRkMW6My+o
gppoRxDdIUd+pTvBVBST9l8cBU8uF2Cl0IBfCin90FqGMRE/50IFXGuIFi1+wpPlvkprPdKGf9/N
LBJ4xaboOQ7gbVeI4sHIJlVys+TBkep9dV5i0Dhg1s5N+onJb3KLIOwBduMxrindBK7g9L5jLzkh
C8vxtvhXU9JJsQ08ShM/gmkMDsS7V6LoxcgXZVW9uD83vMkZCxTeMjPd3hBED4gRNSfSIZ67+Sxy
usFPcoIH/T6Mv8lryNr334y5wnSv73Qv7GLiQZF3A4CLEu1nJALj2WGOTbjTzwgIYf62buH5Wins
0dsnJOpkMgdD9NJ/SOdFd/9HJ+Y0rHBgLo5R7v5Ho8uKZ+tNViA44TMReDzVGfmySOdhmEyTTo9I
kZTpCKk5qyQ51wU7AtaYeNeQDN6MJU/eqfYVgb4ucGpF4Sr5NxgiBy8QnWwUMxOP7kqicCUMZjNa
7tfrBRZSwBtbZYSRDmglbfl2Fkhiz9CLmBl54QpB2Slz1d4Fbqm/LT5rhcX17c+eG3IDz0N1SdOu
B3KX7rx5tai7sX6goV8Xx+cLg6rcYtklZPdIZ6jFNbKHBo6eZuHbDtYDRQlCYv33UJlxeZZUQ6jc
VoKIsRsw73KLDegjF/d1/2fx2YfPh1UYpIK4/JgVBu4gquUXDQiYEi3lqN28KDCcvPk1WpR9l7WY
+nMRGjaeFwIHnzz+KkoxFK7k8hGLT3AbsS/taty06/3vkxHKazJsLHDUFpFFFylh4pZf3KjaFGj9
L8YmDDu/o3+SEYHPA2qNJWVqEhWCIc6WMFQSiVh3TNBQGAnqVV1yAeqaIs573oNU265Qz8yz5wac
Bgvg6TiyHcF7pZgbErlFYZp6BBr7lxsC16ygN0PQzEUxwinL9rAz2R4hggG9OOsyh1jG7xf/mjrY
f4JD/eJoBiG35TqlzBrB76el7+3g2zCSlsH+QirXB4MfmiRhmfAkPZxdz3vTTe/2NPI9bxJmGuCX
7M03ahNKelQBCV58iSa20R+95RTKQTJfwTUYcvqHR+IR5vO8Vp29at+BUI2v7IcdOrKyhIzwNx8z
LP9nsf0+k/tlNvkFSc6HwHCSmqJnfb7iCWdPclEc0TsC2H9nks/R+jAkCFBDzpCyXT+4BouTYsg8
hDQZlsZe8I3QHrcmvck9DC6bbcsGU/QHlvbdYj3y/+CD5DYBiBOhpzd2bXwDwKWxPRVi8Kqv2fpS
kVE4Hu4q0JmovNVgCh7wj7X13w9Sm0WmEPfh+i2/Y6+Iso6M8B8vzZHN/cNKiIvTt8k78/WjoTIm
lEcamXh402J8e+V+Xra5ZNro0szGYuyajOzMHw1YF6iT80V3YzrBUcDleUfoPiUHTihTpTvivW+l
DvFISNCBuvI/z3/Jv/LsTXcBpbxTkn1mlP9lcCMFlGm4UEUG9MoL5b9e0jxvZ3KGZrpzlBDDU4PO
0kP22YFQrZe+G4kpYXo2JG7m+ot3SULpXznDByRxHb1n1JRiGohniQvTKSsX/k5ImaJTB0UzZau2
IDXqwiJXaZLtQa+OS/gbV8zmtQMz8QzB2+uZC9bjDYdXyBGXbt5jV3btKXHTOC/s3KbimaWOqzp0
03rtwLn868BED33lnCspvaB3eQPf7njwvX+1OLEl0ur2fZWsBkXjqmoMWReH58cvckHGwWm7sMaZ
mOHNzTjN23aErqsdeZaax5Z0dWYi9GsLHfYXvGjZaIZCoEqRrS81VfPU3or6QpbhJ8KMeVhX2BsD
/rvbQ2SQ2uv7waAQNtTe6HJewV7m9fMaZdKuFW+NB70zKEk3z7utdSk3tO2Lvq3dR29HMnq1InOB
IKxzMd+1PPU8eNvmZO2RgiBjlnrUa8FadGvtYGvMgWfHuUhPq77nm1enbi50uHzZl3ZP7y3xIl67
SPbtS/niVQJMghFdeivRzx+FUuUuQrCXdtZrnwVbO/vrqt8ZWCcvN3fePxmjHY3iWdMmcAUM4oye
0508Y4y+LQ0Zs88y0B0dfUUFEqYav2rfxCkFRQYFFsLkBLP5Q3MD5ni3uOz7PleN1b4XWzV8Z/k6
Lgq4xOnCWtNf5uh9AN3ImCgoCjvAmTfFCrz3QpaPfDlGp2QW2aw1+I0YMGR1pI13yhffv980xnkG
5j3dF6t1cbetkpFF/FOusQxmzWo+NFXgq0198BkcxbPAWKjCom0nSmNDZD8ToNOCDizvnYi3t9vl
Lf1BJvIvDbdxwuozAYOAOW9YnnAHjI/UlIUefP9XT8j5NxsJUwGBDWplvksgFVoIdYtlBjTh6ZFM
8G48+2IXeQtc331nSe1VyqnrfbcRF6N72njvC42aHoFw7zTCUQiB0BA24BLGMC/Hns4yF/J8ZupU
R2plJA4fi9e7eoiFL2nJD6IQ/wwcfy/BZIGSLxt0nLbVs4yDZ04PCUN9SGcmb5XNZ0RTYu+Tlkt5
KxDID01GCuBklOosH20ibd0ZYrJHnMpjwTM1ZQGCk9cz3g10OTTvyGNMdRzE1xsCzzLTNXiYDQ6H
wzEzvvO1umnVqZwcplvYt+j93ZxvD+dGKwUfEdH59cdQBbBfLe919KtVkP7vvdVolTkwDAmlhFrS
dlPQIIrzWLkS2u180bfICzf9eoXfGzJVQHcR6CyjIPZVPXnQqAs71u8z07qtDxVylDPTQFnufqTi
4vtdGZgpo8BcakyyTbOuP22gTozPmA4WUXRv8rT+Y+k+Z++AUhYHP+vEM89Vl4bq8kdROeyKwvav
qJyItoztcQ7Aodqe9QV7cr8JrTkCjW3dLckntTGjp8WBd/Mw81wbXGnyfB0LBuci5UJeCKqaF3RY
vja1OLW+jTXyN2V0JLicBFeuDZhu7Vz1G3XRXoxRTdOmln6rfwLOhnpD1wUGMND5ArKyDvlSlm7k
/gQ1vf4EurFYVjKfjjaVIxZsm/NhMmvwt9J/f8Lz2NWs54TiVmDC+AS3uBjuCxzgaZI/EcubFtIT
tsC5A7DTPNA5UGUmFhnJAoTSbnRxQo2JmQKJDEkgSxdVWfj1IRplq9CbqjPjcaMB0UJWtpK4br86
PsXbTO2TVBi3yznwq28FBPMN5lDvxk7wlojRXKOfBmvVEqeJJw5OxUpo5BI8398v2aNb9/+36E8s
lUE8F3Wc6wz9NniJtvaszDrtSUhWkIHph1M7lCJ0ExpJKlXJmVw7k1aimDfe2pd4dRnt255dxilD
pNzpxRoO9UKxCDS4r4m59VaDt8XGxxEFYFAdU1gni+iI/8Jbu6JViIi9L3bPPkvXJH6LcwRcQrPT
TyuitbNZfqU9BnSEuaR5pxyhYp9RTqELN/IAntQDhkdIPEThaJX179QBBkFe0yakaetluRTrMn4Q
bFpGnzpMoRxFjN4bdg4frduydTNXm6f1GkZyYqk6n38uY/ks2bUXB7/GmnqdPrc5j0ntntJOCCIv
F7Ooj5r3Coaxrmo33+T56Z6Sg04Lzy16oOeKkRMX81hziO78wGplcw+tuuiTbxc4BjvZvd1H0K+O
VeKPbWMO+nP00usSZLNb/ucKKON3i2FxzTMMm6mZah/km/I9AxZTpTL5z2Cqk0CapPwWBFey5sl0
pC+O62JJPBbsqmBFBEsjbaiQV3Iu3hERUSSraU8xfSJUm+c6KB28L/RzyL53Z7R0lctJT9BjHJDf
m+Dky19+tP5t2pBgDiep2Bqku/pkVXhcEl5NZYPvqbZrriDsgUg9TOtPpd3+N/7gN9XuymZPvN9e
fwVB5ZUrLP6lsjb05xD+KnlTdJmQFt4tP3WAgkvpNVY+jC5C0Y+4uc6o76qJI8ZOc9MY5+fYdmSP
tRwaUsh3iI76y3kg3LwxJpvPZDiZb9AI+B2rkocCLfENmxkukb7atiTqzp8lpFIK9VdPqthVMQhx
nqUCqXA665zv9No9N3s6pM3shE3QhZrS22YXa/b1MnI5h4+hfWeOHi0v4yISKf6XHd4C7z++XpLI
JKtYFAkLrDsM5miu1z++gbX6dIHL/ipZTPBACRHiwt0AiGEEkomUf1tQuaM5Bg3w7wFoDPHoVGJG
thEGnGf56w6aw1u+yRWTPbV9TXJcusoJzaCzlahCfxZ5sizttuqnhr5zlt0KOJTfo5xAb5+Fzfev
CP+az+eheqGvFi80s9r2yF8H0r/NmQ5h2MCiR/NKMCO+9u9SW29+L6LEn8GGqvFjdgVOPP/1bkUS
icKOUIqa2u7x1cmZ4p9mFv0HbCX9JBG/9attNLkyXCp4BubFcv1cE1a2CvmvkZ3+gtEnJ2NCf4LS
0uLaf8wLG5MkWqfNad/PlgsRQPM43+e+fed4y17tP0yPqzFY3bKBE72RD7QfDZu/1IZ5osQsFG7G
B88oNLn5IhqAL6S7Xttlebxxa1rOepEp1QzPvY57Jo3k6Hl8jCIF/nHowB9zOWxBU4j9gI1e2OUo
gMUfy+z8tuhSfRBVH+La6sA18iFC8h1NtMVUauoXhEYiNE2izinCRNQvOW5G1lfEKXZKD8ooy07L
WcwnwQEE3qJTwnXfv0FqX5w2S3lsyrZiptCew7AM/qQSE0kc8Zfm73OAzqavQ3XMtxzJItpTOOKm
xWqWf9moMdSmxiOhMF3b0gSQXF+Jktzb2zOKfwfX7LSQdBeWvwgQ038J5Tg3/ZI1V4oVia+PObud
x47DdTTWmMyyxv1nPlyIQZJyP1BnthviYn16YsFgdinZyPJeqrmO9anb9S5HqTnyExvP8j7aE0oq
0lh01zbCAv/8bwXM0/ja6By4E04Y5pcb+tvi2TMme3MuH/L/8UpHAhcua2rVRWSA1e/bRxtAXNh3
nRA60/XmWPD2etOKc3++vpD5MXDBFVhoIjkg544xe7kObinBJ6rLYuvbM0CX6eFyG/Ep+ekBfX4W
KePSuXFEBL+Y075+BN5woV/zxFla6w417w/eUWdGqagv8cXbqz5RGPChQWJuh25k9sZWGlcUtM+L
zOFk9tCmG9XEbXnabpIijLJtV+6OL4JDw8iIWt5NgoF1Va0biwIO0RWPlhBk6SBgq1GaE3sp6iRU
5iBPr8qi2YySfyiSQ54fEHKfcuB5Lp8Wi0rMiFIHKF4jZAKJWEvrk1EhqpmtYDgBlJsZgzGXSthR
DUDc9G6n9O2X/PWF6qma3xeXMvE3OKL5dh/3XL7GlnpAlTuNtWDz6TfeQ/u6lG1u1DUSm8AZ0/MR
VpSdLGQ1Pokf3QycK/6je1JmEw9Cr4wvQUXQzhtGYXy+Obs1p8htlAewGVz9hmcqJqyuYDrbzy5J
w2bjmwQbHBaFq8naSwEZo7zKKaIwMioEjwNB9vBh4NeA6bzQgihi5yxBSr28CvbzNyJ14IHTUZBE
ZbK/UvqCYB0Gq2xx0zPxKMx0Rh65NAyE2CV3ceyh4O1zonjfwe8ghYwy7oLcm8DmBL0RPA2WceyC
v67aG6vMFqjzSLC7ByqNnnNv4Az8wpqPbUYELIrV8cgwGSM7YISdGZslkGhMu352AOkt0A1RMLy5
mrtjkAkDksO+IRFGhXonJQea5Mti8mGcCU8C5H01INSFVdvGdqXqYhGDdH00NZwIc/aPxpy+Im+y
yuHSW+qJUqg90Z7tXl7Txn2Of7kLQZnkOoiyou58tNQYyhRiMNEvUi2Zt57nvMdl4httv1x+IXKm
d8Lxpjfu1olaFAcq7a4xH6Ueqwy4w7CD+NP+lLzn3jdlUAklosSFt887DttHKzNMTD5Sq11WRiAU
ycH/IwUtHFyb2NbcRcDIJeHKgUGE1Pw1Y3Sn7xs82nT1azTFUzZHlLS+kPkkJ/lYrL4atFnzXDBX
fjHvDWIwXKkb6+JKTM2w5WA2Lo2KBsYYTui81aLWqyrcfkVWuU6x/KYKyaoYwp2YjccAFKqBAmsA
rdp7YZvm+8RN9tUU2xiPtoawrQSJzneaKNIfo4K5mHbEqMvmnbX4dySB15qVWeJ2k0yFbMxTM52Y
u0AXLnaOcNNDvGMOxCAhS5m3amhR8KRE2np/ztz06XoSvrOdeAcDKnbo4MHxW/BzWPRP+ghf0t95
50W8bTsooQa4n1OMkZN5dZE4J3vKZOt6QrTN2TqtHoW37X+BqJRBDFQo4JYlKAvqeFIY22CupeaQ
j0Ix/RYNOqgqASjhDiOqUmaJDuSxAip1644Y2+95bZuEykXv7NFLSblelIkN7OadiQDCg0HSKzLJ
0fBQv+jStKOu2VaMzObUFKApPr4Cjx4/j1MEKzrP/GhPtArEzmvm2Y4fS7FeyzGOGBSui69thYjj
dBy3zQOfHdNnyUprJugHjCAJAZESE0R9yP+O48sfP2BLNmHX1xzL0nZaHHVYSSk6bSDJDd9LCaee
AsYye85+ijGOS8G9WNpWuvEtQLIy2pI3IXLoL5tYac+RYm3vPmOvTN77rnSLLtvv13S75L2i134f
ngRJgdPWsLMt8Sa2263ylu9Sv1ZnLYusDb1S0yCs+mLzaqRrWnrLKUyU/ysC4H7uZJL5zDA48tBU
jw5Po8VQ2ricdMgNpRDLGIrGgGKMnNT8ErnlDohrqWatbAMoLy5mKy7D3Bspf2MyN02SlNwQB5KI
lnlqHs9RAWy8CzmrDpd5/aj3WtyhDNnSWXEfNHz1Q5d4i6UhvOwtbHcDJV1gFvnpCJYTL3rIV5ON
eeGorieAaiWelE5hrWr9tl+fgM8QXrRCknKUeoT1vZPknqJgwpFnB/Ys7sV4kuVBNeH+yjonvJAN
GghqV1mu2QKcWjSE+A9za2A5PenVhMdI2SdHexiiJcL+Z4ZjvYl6O7gk7KXEGiPRiVDtw6Udd+ED
+Zqgn6dXDKr3al3tWPfpRWnf2vnzAgggN9dQw1DUYKBO5o9vLt5MmoL7uV3HjWXWoGTxX6G+7JEj
NFdrTspEr7/xFMG+FbHF4w9Xc9MQZ/DLWqOcGFuQVnL/waN/Qash5nqR0WwKvWyDBASqEhgxKitH
S48CpP77LOfKUoE1yTLJmtzpWy6vOzhAlaUPwbWuDXd4iJjVijp+7cGSs8eW13y9DWkkCrcGnkvo
0p1upELj1XOB8CDntuYSRAUHdX5arhW99J2T0lJg76uSY5xKfCP/Lg19X0Axfx4MqfEH9Y7syvQ2
wneh0UyLsjaL+YI7ZjKfq2gEV73HmbtalNDCvXlLHFZu93V8pUOWyyVwnDYcpzILrzcdBBAHzPul
psfjpRqyFXlVPLcMKGGSAUJ2O1hLBTTaUevyuS0T5GkkokHaI3egEfmF/FS2K7E96bzPAfiikEyS
6K20V6dFWlR3k4KkynVSnyDNGDqMR/Etfs+7KbXvZgL/NPR/AjzhGHEJpu8Fv7rj7rsFLhl3kEPT
SJiANLd0jWZrt0bPALODVbXZRv0xNkneFbuBLcVN3HecvnTedWMicMYcWI4/Vl2WzoqVdvR71jpy
TNaZ0JaTYkyB0RxDI2P8HiAe0tCU+6NNaZsROYR9F4YqbJmBghsbY5BUEug8R0Pz+6OjojpqxW0P
EMNmLiFoLCJxvpDVLK7fxTz7buutzn+6te42LzgTCqLpVVBQ1sEUQHLuzmttWcmEegiPYWMlwknv
gxdRwxsRvYFoyoVfPpsc6xhlFRCVp0cEOO2t3znEU+DbxkpVSB4X0p3lJeZgBrMnAFkNpmE9sEU8
2JssSB4exAx66jesgX/1q4T2PjUjg6DX9dHw+MStMg77ZWYqMSx9FOWgvr5028VVauFT3ko1wk+L
eE++X3+kQF3SR7BCX8MdjiIist1b4eodczB+b69LV0jqVM9wMmrSotmitOrAW3PPXzuTloJLu6WY
4vqz722cpVHHthdLndPlwmeZLmWyoop+MbLOj3xKeySTxLuXF/jCsiAG5o7iVGDnxytVH1AfW9Em
8X3CL+whBpPeUqomSkiP5zwAD7JaVtZA7IDD5ZSAUxkUcoXv3ICP+fcU52yw4U0zhZnulq44PYHW
iWRxF6Ec/DTwG3jE+twS9oUijJpzTj9txNmtqdFI6xbRFShLkHpHn0rH3b8Bw+KId6AdEcsQYqLW
02U+6sRwwWdpp+y1tpBlhF1gqeGlmWv7DfTuSKD9Yrarx/LSmB+ZUBZ8opnjEkoSZuT1YZTQHTSm
hFWsuW41ljl+eQSUkylEkIKmfDfkN/7RPe9rbUGWUWrxM35bmipe4S/xDGsYNe0/KFrosF8xhgqo
704HnVmHj8qaiNHQfHRksBXyi3p1y/HOGJWEEEJqw2RA26eFn5wbWLy1GGxKa4SKmPWV/aVWb0QK
xd18pnskRbK1DiglfbbC9HL0xCjHx27pb7gEN0LX3NjxnLhS12rJdlvlmD3rK+o6iw8gp3+8PnmH
fcWBWiLev39cePP5miTOOnE6lRtEYPlsMVE8Tq2oC6iTlNkvSXJFwn58SNmlB569UaUAWuVxJ69b
XqON29hrcqMlwluiLZhQcVTwFjvjS0XbFUPHIHQJn0xP6ydJoiRTGdcuNbCbblVKJbR57unGmgx3
UffEvcg8oaF2Fw0PMVzDMEgU/LnCXnk5KmQGBlpWckx5JcssOlqNFGMFTPkHwLsAs1QZyqwpIA5I
3bP7SP9DTvz2D8GqnFaq6LR24vDprF7PFmFu1o5HmFUNFBUp3MQEI8FsSPOan3RB6g6Nfd0aybV+
lUlITYncsDKpWvPnTIpwlr/PzuytUW+INWzbDwUYW0pVL2RBxdD2OtHg6/t1Miqo+LPYCDRT//z5
akq5JrthIFDUbWluaxfqONTrE21Lr7EN8JKlQZMktnW619xE7xo5KdIbpIpfGqFnTA4+5vfqW1VD
+og16d8VnugForgUIu/bVnP3sLvbElnEFumhDKrxawpUXtueKMvQWZjjy/VFm5ul+D6SSPmM2oqa
MjhRGyInO0TIB269MaGGJkMJut88TC2+FC1JQcOJCtj86fjLDJInq+/Sd5a9e4rC87jJJpPRUvIw
r19qNonlG7CMdrxDjiRCrQMSmWM0z2a51RshWYgkeLWSVyNZ/MXNg/Wg2ri/cP3BwdULMwblD+b9
6GJ9a2u3taIrBOUViG2j+XWahlTm/gNBrxQTgdbQf3CPnh8ji//gDr/iThAsvCF6rQUfUej/xBre
FR5L9Szcz3ERtfGlZKvp+tzWiaNmi0ooAzYx+Kc0BSK13khDxnhpE9iPqP7yFsiNv1QjwBNU5st1
B9oztmmlexPLHwMWVh/rExisE0IOju4Sjup2NcCgj6IIkbaHZ2WJvVy4q2wpng7lIj1y8nZ41b4G
W8tneCPY2CxE/zoKwS28v5oqfLF0YbT2VL1Mx6tQ/w2DWGV7B0XvIc3UUL7LrwYFM2+P+GxPaYUA
3B64sqdQdpF4rbkVHR3dzkyWw7/2NiGYowCfSXjKQxYudEECVYaD/95SMir1DGNStMOtHwpr/F2/
IigQIdI6oM0Zy+NgptxVVlh9uafLjYvbjOjRYIA19qXVgYO/TaU3pJHbtHYazuOlxd0CHvcnbMJP
4yfkJl632OIjSLs+NKO0YVivgakiZFJ+J1bKbfST5EVjKB6PPVHiGwhhD4lPAcJGVNuDLpo2FE6x
ZXUI8X7I+vYWVLaTmVdxA2tsnw0xPcVccTEaT/6mv4wXlrZfB5mBVOtM30QBA7glgUWEhkWIkN0d
ghgE6Mi/BKgOp2pc+/h0GrjGWWSuJkvn/gBkw7HDAT7EIez5OfIfICDO09p9AULydyyGbR9rzCZL
yofet38dkroFcGaijietKsnjmuRYJ652G1TMAv785rcvrPVA6o6PEn6E26AmKWmqYNCpY/pP22n9
XbbU7kFILJIqWq7SmoStV2tVvA5fQUDLeHmuDm257R+/edVdN80u5GpysFjaDdUPE8TgQhjGINr5
QxxG7UX4aR/1st8hXeMrKBFX831gcjpUZCNpvwQrlavgWQM+g96B6gzzb5uGAnjtRoqyr4SWRcTx
Jdw4D12nZrqqG4eTqMgSTudhLaSrBtrJcUmHnHdonppV+C2UwfscJggV9Z81XN3dyDS1a6xR54gB
GsxVqA4q6nKXaqMUvBUhveKoZmDVtUH7RObagaT+0OFnMnF4UvpGyzniGKhojhhpXzhxfcH/oooY
+r9BkegUFSR0Ev5oudiTPaU4HR19KPOfXjlAPqNujb4XKMvhNpESXxQY+zxjWjmuWcoJXzWIlGO/
BrkXtzNQUsaKPiUYy/K+3TS8r0c0wvTzphTzwM5e46SvwJAKq1Q9w+Fx4p0CJdee13zdNL38FlpZ
ECKlGETbIwSdRw7bLk8wET9EGVYdTuTrcCNEenew4REdpyXzHfNCJ2Pw4QNSUCZV9CT5v/22NsxY
KzLE9MJsHdNxoMj+ggQ+5GLzuUBqOTLcI85sfTjeKA9GsiFiAJ2B4+KIY8Slo7eUfo77Ja5tBMxD
rGB59kNPvqmH6Rzb7LQnDGK1XcF01ymGQlw2PggUfvNVN1y/P0ltzkWU3MAf3R9LNV5rUeN9sP8J
2HG/fc3cYbQOGWina1OTOiNkYue7Dns/wJa4FdLisa8LHhHPV1+DFsWGvyiRbIRnefEGntZvCwKa
Q0K6V+B9pgFC1pjBFufWuNRzaN8UUbAWZb7QG3igYmCLWLdtEvgXMaOHXTR2cer25pw0jtob0Bk+
xMGFfRPgvSkYtLbYoxefpLUL0EkWxJBZBor2wFRk0br1zZUg7JNFh3Cuv5Sbpf1S1r9YZhL0SsyH
WJR0izt+HNbxkFieY074eSaAQcMRdn/Q/cvS0EynOBnmXQs2NHTa6o+mleQ2hfhiIzcmgTdxt9i1
VjTzukP/oENyt2ZUp5WhuoEnhoT4wIlxKK1gCmnIWyJMmZvsiCs0/geWi8/1spj6rOV1R+vTIsOZ
l4pTAjcrI5TWdN9L4s8C08fgVwMClRSQzNitwVSx4/ZazPz/8zDcEU2j9w1mfqownSz5pjCkKtAJ
6a+Wy0rnHIM3MKzo2cZ2lIAwqA09zU+V0P4I20iQWEiiL2ypifkCO8a3rEqydX+npmLyIeSyqXVr
ipgzz3mKHw6aYYZ4cERzeedqy3lesNqWQGdfxWnFhDbicDP0bDFgC5HpJPP9APl+qN7gIRuxqNwI
RFxQqm0UUcEyfmg0micb7xzLMhpN+YzUZ3kqFG9asqn8Hq/hNf1xD9JlDqzkdDrnDpHOZIowtDB9
/Iayh4toGH89sGcWOzGRnIuET1RPJelppfJqgp+zSuUrzoYt8QiqJ50RsvltgbVBQQ14lTDvICuw
e2rig3TK8v0Ep0K4gnW0G9lripFjFOorVpzMP7wZ0mxGeun90AqR4FC0QxqqlB50D1FnBJ7T0uh9
6ROwHlbd/v0txDasEnWeGkcYrUKFDKDESmeZWJkfUKSwoH6IB8tDIu4UBS318R2LZaN7wHmjoxdS
klrdMU/X92470YjKWGQW/4EumLF+kX9WJqapMCCA7UATwJarbAyMSybl0R5Qvg6jhJcx0iVAjZkB
TqT4iSnK5eKgYR1vnp8JHVsyCx4hPBnTrUpnKyKzYzQScM5V4TeBZUSZFS4/aFGhiI2DLG052OlW
a7k8JTMWdbPJ+BAst3jbMYMnpyS36F0/wCV6BSryFU4XOS32NsJWZfLPa9wG7Qxs0jd8+GsGmcc6
+xZoOHCq/JXLNY8tHddhL0cmB25lCm2YRRHXEqQjcUvSZWkgIatIGu7DfEn9uKY/HMvyky+QssZ1
qdK3QCHoAOGCvO/P1gAqWM2z0mnJyqppImxeRvYGQLnW7YCZ5J6gky0h92BKMMjv9E0wlfYXVa48
+DdRIOiMr2uJk+9TIi+iLli+KdrcyxQ2mXQcF/1TTMBmlaGCcvJh6kw5EyEnh/GKwcX0bIn5xLkG
W2ObgJy1e1Y38pN1SRSB6bVi3pQje30Y0/aG7IpO29qRTnS6PtRMnOY46FnJwkZjggfzgPn2AymQ
3wpN5zExCzKi706JxkWdz5hJcRRitxh22zRAUVmaPDv8Ul2ApjXw+WkuR5f8y7qHU04posLn0pKq
v1z8kMcGIvaqrDzIiCACY7GMX4lFGPLs5zBbjO30KApHU8PRkB621yewHb8ofBjUyvJD8xcT95dV
Flzns1r5GXfYu4EwZMPOPNY42c8cNGWazUTUx6OnnV0iyNS8UpUqnDVYphYBi3Z+d/OHVWvCMmr3
wRAiaWZCfs168m0YDuQtLexMCIXajbvukCvBtBCQefR2tdHFsYaaHGAK5Sp4Gm89zhLDXyFQYmts
qaC6YWQVW4pWuc9iZGPca5yXkksd0SI5ZIx5JiqiN7cxZdjYjvivE/LjDWjanJG+uRr/DtB6mqjM
mEnj+YQA20v4oOElDEQqvLT2QhGgx40a6gy53+5nGpsZGw9MHj9DGaHsybNQfJrBDJJEzJwEALar
i3HUqAZbU+BaGgFokA7TZhnTf9nf2O2O5Eg/StRjdk/8b6tstr+h8MTWx0CgXZaCh+w9jZZFC3be
sU4WiL4xnUDk2EI3tZBivFfRe2i68pm41855vCGBhpE3IhfB0lDjzgc8F5yvpwqSBa+RoumYdAnL
Ttskzke1gCoso49RDkJ5YwSqqbqyJD8mH36kFY+dLeohR0aCGSUdyxNACHjroIetg+9AmiuTS0UI
OtBuO9PM2Vaem3wM51Tia7ozCKYXYU3Mn0E8JB4tFNBKeoK6kM386EW2pfQmLL6+dkXe06vdkpJy
OD1V9AU83cZ93RdQs2iyfR8BgNp9nrs1rm6DXRXZ4ySFZQXUbCHNFjyfF9KWzgNP9qp1GZEsm1xX
4SBhBH069RVdZS3Q9dNTy0y6aMCaNtZWKvxzZiQlO5/Rww18YmHzWZf0S/p8LzobX5EkrIUxiU2M
IwzRxET4lB6nJ+FCAZL5FuAYYVf83SkKnTyX1EXQpCNNctE2Rp5zSfhBTyq7npj0sVJn7rxV0g5X
uVWTOxuoZ52ZFLB97W8TVfXHkdb4xjWJJ5FtYlqCZMh3TWyjHox+ELW0IGB892B21guc13vZEjjn
i4zgKsKVaY96INYQL7Axu2YSVw7Y2/PgD8p+UuMRIB0uw/iSJ+jwfJaR9vP1S8j88au4k9B8CDVE
Onp7RRr4hD1NeAD61N28KyLA8LF8fJqNYxtmLqZhD89QGLARTit2zXe+qYfgLesvEJUrcekTXU+M
R7Ptb7sXGumGLRQc4mNR5UCN5z4fggRdQMETGUB/XUCq044nEMMvQGdzB5OGGSUnijAqfwEFw+p7
QgPsNYfCcJVdlcUGjcO+EKFQhX/VA6VHKcoTJvjBHTY8PD6JQAxU6vdEFpLAFnDnPazjg1yJGKCq
j9NzQxGWbsFr6nDnktejireKXWotirbX9bIgSZIVwr4Vwkey2VI7hDgYuTyy7921wdYYAC3mdV0z
ow7pPZ24u4jIvIfZOtfbeimB+iXGTZjfOBGyYm9jsMctIIvZjMbjqTrcWSawQGFVrKbYlnY1QsJs
yMyM3vVYu82pkkS9hyfB65gQ0uOwypNu5d1aXBWAURtJ1SOAzGyPmsnsNVaygzUpY2W1zEqP8FUr
DRIHOiK9yz1RNyeuRJmO9G7P8DebSdJ+8fMhdgpHxcAvUXOCL4aGJSy6kEVu0NOAzLHds38H8jCD
z1An8D+7fOTv+cErNK9QmsDDewlGe2DJzCH6k9esuLarBkxtr9Gv4JGmNQR4hXeiLF85yk/5aQgO
ZPLmRAqkuioOzC6+Y6w/JlMi2X3O2+Fbtf7hbfn2hjMj5JDIG1iAxuq0WXPmpdVL8Po2/UxuKF6t
V5dOC+jxOqFHanCVweQXeB51nK14ckUNr1vhPOlOwUXQqrYdAwqUk7U/zXbMWkm59wYoeXNoFiBD
Xlp7E/vCIbKQu3hlA9bQo/SPyFnvrjgkIBZQUXbuq7M3zFAmqgL7Db3u1DWSHQ6yQYXA4wzjBKkE
oYS/wid6fWkmJyRQgggBpEnRU6oTVPN6f5D7VyXj4aJ49RyZKWzDd/QxS74sfqQfHQC9uzHD0H70
Kvb4hqen3j2JMY+5Eo5lMi04fAMWxm4MyYcvjy4lMyZPzuHtYqpz0UmcYf3m4HnPhDwQy+rqrQDS
3tU+0PTKNpe5B16Sf3vBOJlTi4kG4DfMPS8131PtWHpWtt2EeDAnV0rlhnHY0Qna5nLRewW8dVFx
+0JO+GS4gaIJPspjZWN0H/18K06Hs8rxrgAe4CHBt1aeeVcnvA6xtFL69rfc8SNeJKW9IfDzXKWf
H6nGknpqFtO2uwjd/8CZIdrVCfvy3DsVWgtWG2Sb2FlQ7T8vhiyku3LCBFNFCOUVfTASXwKSd6fD
Jb5CshGDGaqtpQkJ+3wr6KMoeZ4QzuSzuW+HxsgK4M6XTPvxr0OYdU9sR8uijTqQl9A64RM9j758
VoLxdIQRO+hoZFSM6cMA3kq498hLn3Q89FuNO2cA/z0qFFV+SELg3ZoYIDGLHA87Luaa5YQGlGao
GOsN7U8oixQqdibVddzfkvYZRMyDc/t7NIN2xhXafWWmxGVKUUihYAM5Vnv2ZYmMNT/lAZVA9CXK
NL70dIq1FoytlIrlBFguEQPVhogkyXUKcrVOTLu8whdisJa1IwCPfRQeKXdEJ8kKTaSUylz7qnE9
FZhW1u7H0BzvmJqOtBb8nbMPWkHTfVx4DUuiv+vHHkpG0g2TlwuY0COyiHX7B8xS7KDhoJ/LWtKL
KEnO+kBLW9y4PiqGwt0gI1xfvgz2wxvG6EiScVpYkT4T/LU5l1dvkShNLvMIzm5pfoU1ozmRFJiw
CsQRKsXiQCSBb4r56wr/w8ccP8RN+EoziRj7Z9xUYFD5P/4mGVRmvfyoqR6JzO8zXm8RDYzeq2aj
doAve/7ndenE1ejyHvh3fg79K69442/hSD+z85C8wkYeVE1v5XVhGjZrsH3UnUjsJJFR9CcnqPMv
Tt4lAzCoUgSE1BshjMCOcZAMjg1TFdMehbpnBHp3JPi7sReh/b3NWul920PN2nxtHvz+YYIPAskn
jEdwTEJ62fjoKodpGqJAySXMutNSD6NL/nW2CSnHxz3eotszneOnmVzrCS4bL6/ziwKcAIF9JWkK
0DmTr9SdfVdpTHtrCz7QQT23o5VWIUO+424MkxbvznAok+FWpEhz/nahboKzIPH8pphUmi94dqKM
er8QGj2cstY3nwt7MVGfiaCK+lSicAIJIZDrqwulmO68EvmbOGpOYi+W5tLZJsFaQ+kvzg6hwdbt
Y5vwbjMltUtz2u6fTudLVLQ9YpA+0VhdZgN5i+mwk47ezn7wxgiXSCsLo1+J0gOrhAibTURPsBja
elmD72uh0aXuglz9nOvWeM/NNvy5d202kDsbvghUHokN02i2MGPrqs6uSuNDbljawfSgtS4HxsFq
cIFszynKD8FcydOZGCiuAzF3yWj/n9xkNYBuQPq2eGRKx53BmXKyJNSVhpwy0o2Nsmb4RRbd1Bap
/4lP8s2gqnBUv2iwiXCyA8r+aO3X9p+20dnXUb5Ry5ZMkl0JdPRXmygUGIxxzItPI00sbZp8zkNA
/Ms6a2OmHpx31g+J/TLXaZ7CXl+EoYRW1aC4hwqJ/7xQxAjWfbSf0mnQgCxCW938ojZOvqh3w9iV
TGN5jkC08AcBWcHcTMtBxSmvazEVUC7ITs5fatIdydghJRhn9VCaEQ/KXDPFhjDJoykmmUFOU/72
o82i/PLyGIqUq1ItsB0DWTnGRNOdM15wyAQ1CdkO1TTijXUgbNYGaoVbnaA8ibI1k8wsAzbhewR1
P/Nq8QZ6mYB/uc9FWL8C31s9hyKuHX2AdB6JUQkJIuoWwGZD297aZJtRFZp7+ER26zRy9Ja7qAMO
QHHA4E9weDWpchpMZLfvij+OmgeTc7nPKcZsPUKahhtN8Guxydong21hCQlXMRgaY0jcHvd7kAUb
42gISccpaFCdwkdj/8q3IHvOL+0Rq1nY/KpTT7DRUSWcuhNaUTyD1ZTTeZS0UvNjs4H6Twd3wjT6
XTuQddREyNU8N0VQQW4qi76CVUp8cRUNmZVpaPT1HF9lZ0QLdqSniHT7N74xuGOVq2ole6FIdArn
A0bztsYOC2VnUvjchkGUdHgZgpnaSXjb6v9gMQIBfKMIH8Bowh4aBcGtq1cvmYH6mSEFSu/Q7tQq
uz4G2S4ZrDD9YsePOdKX7wsvsSahf/up2G40C37GVefsh6zmEqJA6oR92g4Lhu8xd8MbaXbkXobZ
ZlwZHCkqT+fM5uB4TCjhc1bH2qMCZgwxI33u5/cTwSYqcy5YAvb8e+sHTXW6vw/noWubEWf5Mh0/
ZtHtrXz1okhMejCEwyUVhLTZCnxIIBmpKz/8mVRxiqMUfn0C9mlZQTGKaTY9QWHn7aFsJMOo0SbD
AbkeX0ut/UbN8KdZd3zygcNt7vqNOzjAjhHY2QKk0f/pSobBFh3x5nmrLY7NFO7p2nO/gWVo2KXp
6dWuWEA0WNNo9lmYtLseoGXQCLOknZC6qnG4hV9B4keBTMyaMcUWGs8ViHO+TXSOP24JpSrAv1Z6
9OJ745oQ8FGIioABuxiLnVTAKD8ADBw1DElsgA4Mi1HpNFz1MtJVD7M4OB+qfiSqSXmPJ1vH2hlk
6+6aidcVoN68NqN7BpjK7l1Zn3/Obpgj0aCPUVZmwBFeX8BMo7elnn8oTJ5WQTZYIkkVlaX5SkwB
qsyhXoP8FsYNCq9AgX1dNyR4OnTFNVSupzs5I3U6eBXKWRrC8NoSnMC34ri1dRNRb8BdJ5D0Gj8i
oSIZ1RpVZV3opTgHLWPiONJSRKfvLP0EkFUcmeeQ14uwEtVJxz8mLXjgkKJKhTXt5dGu8Rpc+EyF
OyKzCoJWXoZjE8lp01Zx42lL3FH16By2gJSwIxLCc1JMTokeDgzbFuziIQmXw7IST/Vu3hHgoE0Q
qgHhZ3BcFe9vKMDh1UJqFOrSp5IaimlJSOVfxdxSZUFA20urOdL8iE+zzLqH98L1W5r/sxzkhpa/
eR35OKEjZauhW1HTUj/8az3pwCAwJvJ7QoU1BpzEhXwzAZZg/iDO7RJpK3s+q7XDVnhIBPuBISLf
0F3RjawzZ6h+anTM8xw+l4dy79VNuhRxvbZ8TEzO9lNANcERrPPa9VSJUARoDOtg4ZgltvXhPU/t
KMh7Hsy5avJRcSbLeIfewkcTZlbLTIMTli8KXSaHoYgmhOTGJCsnFaPN0QBb8yN5ioGZEbE2q5KR
PFuIaH/RNCxMNKL0BdiH9VwUB2YmcvVAqE165McG8hy0bdE0HoL1MhjqnkQ6D9xC4OecapYu40NU
yZXD8eCnmzOnqD1SSkJYGct4oBgXlCjg4cvSLWSIJj967bC2zlRE0wt49vKCKlzzgf2my4EqB7Ll
CJMt0a3FUpO6ZQOxFaJmnlrVZ4UpFJmfOEez60BRf1rnP2ubKhB9TPwDGU6Te45e1gqNZvM0w2L9
RiyJ+FtgE/zyxJgT9oK2AJe3voSoycK+Fpfp1l1P9fEtytknqfE1MNDeULzqGD2qxK6ic1ZFGwkn
PRphsmg8vyBDW8327Fs+uWum9kF4W29zh2gCWWZiclVJ7G4q9w1uow1ZxO7O6P1rrOIF+/F72YJ3
T+JgJccFvq0WybsZqoUWLWlOl8DDx3QPhrEW05cTo/u9r/lyVt7trVrglgda2oce9A7RnvfDTSmH
e44bi6RkuOp+4VcvJhFI38/pG4Tf2PozTY2FGlHpNads1/TB5VmgZ0+biyf2S0fZjdEjyMpwbcD6
jVrQxp4XpGKx1BrzU5v0jwlQFmnpklQjeEy/XGxTiVg/6ceFM4sfHiJHkGE113dymDQfTroN9lPT
d8abQ4kjQsQk/5HZiT6vvtXkV95BDbBVSsitIl6IK1QW2s6tcqCfM5QdN6nM1ZuvcQhXlaI80VP1
yQatOoFKuVh9ZEeLAVCK9gjTXaZxjh/6y9/XEoelUJ6L9jzKCx415cBsOgSS67MaXgpgXo11VfNe
5F+lTE2+oujr3HmfxF+UTxtk4yLQtRlJRHuEN5VCPTGC28dOpK2rBlXjolfNyalAvUzFcIYJOb3g
cKnhK5nQ9rRcKpZ0t+gvc9GRNDudiobne6wo6cFpAfaPLJGB/fcmFWBlQ9UMOMSXCgvwYWWYdy7j
Z6121CcgF6Ye4cdiGfSV+gh6jlEgO34xlcAzgVPUTcQ+LQDBsv3YV0WK3nrM6zX+NswNBl6PJ3Vu
m9GUnAaMCGH6wpvMpnEh3q+BPnJ3iURa+R58CC3nUJyuBl0izH17Uhnc4npU1OIUMkexmgefIcfz
29spuWeuKBVKAKPAsUv4floyyFN8MZu2qeqUU0ZX5HpP/B6h2Kt9mSl1ajjxRzbypH8dKobp+DVS
7wcuizKhb2/9E8BF9KnXDvwK+tjAtVTmr0nTRuajzgOoYR+C0/02HzJyvnpJx/R0q1SJ/yY3zVeA
7YsqVDweN0rx0yu8Ma7zkoHVG75NvthMYk+MTBS5umjPmUg62gSgwPM5cTVhLFPd275eMfIimmKG
f3u0iynT61OKDkioWWQ0MD9I5HBNqsn669zALRzjKwvaccteX/OsZ8pLiN+em3n3IibDtaolK/C6
lQNypC8A/27ckk21Xovp8xpmQ6GBqxYi7lmMgWsTPA40DyK2k7v6HhWhUw9kxekWAEkhAEO8ptKn
a0/55kD0lmjju583KFHTw29Ve/BcMmA9fG+Qi1s9h5tJi3qYIfFHCujhHrfB5CoDx8smgtdoqU+S
7SZnhVgllFc7lhOAGYjupO7kP4nBwQCtLQkVI05FVCTyBN6yr9P4ZySWf+w3IOkwC5ixkmsmVHE3
Oe9Qh6EUue5L1DcRH8UO6mRjfnYed/u7N0+OnwXZTM+Tv84lWIUb6CANcw6Gg5Qpf7anzEwGOQAE
whMFP/WjU8lUqzQO2wQizrYjJFow/wCwSAjIaDAgWGcJQijSkf414U+k08EtWAPW5/2a0Flcwf58
Xc+3MlBuQ0keiS2+SdxlKAqmaAN3Hmv8NnwPMkln/v5IeYCbG633ng9L+TCtwzkzVCYHz5fhUHpL
uyJBXhNkYcyHG4ZeK7LYStDkwE93Ce93uMhsOFt/xPYaetc69x8kwChdOMD6D0Z6uHvp5TP51xgT
2oYqZVF/mn4jEBtnPgEV8150b3AUw1z1zQn7nu4bDoY+7wllsakZCIPHuhKy3hkoausICZ9LBgk4
sHMT8WEdv3cX4AYUBroEOeaDouzbSRkAUPZuV9A2u3R6SFeNKcAHdwYeG1wbohERjsQHw4LGSKLc
uwH/oGpm3DuphYB8ZsRgTKSVkXrlTrtXUz5ym1ytM8dIWa385/SIh2QM5OLjIC6BFAVWMg/6iIep
2OS2KnwtiZwM14hlCYjBTkJR+g6Qpk5Zvulk4IEmTAEKvk5yMR8g1xlkehnvTqZDpj19yzziA+7m
CUt4qZXQF6KQm/JeexRnliZRyz1LnbAc0OmD+cgdsCh6xwmEWEEwoIqKE6oerPWRVEtECjmFVx2S
xntG53F8+XJ6Y8/zplCoovGxuGI7alDnlsHoCerUg9P9Qr19mJyoEwDj/Uy/0mvVEhNp3TgMeKwL
+adK2DHfnD/F2mTmDLRSk7gORxZFPZ9wXsVabuutue1PyyXjqHKxTN5hI+A4+BSq+YMzsBiIOr+G
rBZpYW8wc90q2lZp9j/EboS8fWR/a2tsOP0MH9hoHnEr1Yj60ZhkIsBDz6RBnUxk9J6KrfSUdY8A
l9dZ5FoCnLElHiCIwKXgNjCAKhcEwUUioXcvwa+hAOIRTI/Mvu5bMAonheDsyYPUzIIvy2WStX5Z
lWTDtOkqJvtrkNEGdpO6xS6OolY1s+zYlIT1BXUJhJR3aG/BohxW5BM9NB0BrT/A/QYQkPQqz8kT
xDu9wnTi4JJv6QjAnKxOgk/ubSqpln+xjHZg+hfKVo5zEG3dvjLKZ0DpjYGKJBZxBXs1o/NSwFN5
f2RKrpiUbS0blAZT1mQPqNJyUVJcBaeO/sTOnI7jeuT9p/RjU5HGUrlfku8fWuoBUpVYkIlmZNjB
gIGqbOrFrNDXOOpxd0zjNm9Mm7Va+Pbe9vJMKV7/XIVLkopVQ/R25oZ00EI6tsabXDKfzoUy/Gdu
kCEBy3/nlUsW2eXTF1+P4yMUyaP8aZLCbWI5zRCPdo7/5X4PhhacQ4lXT8MVThTPrDOhyHGfz0ti
Cdc5y84d/0VAgRlaFEsWqmgiV4hLgWKePy/ijN8xj3EDsbUKm99M9Hkmut63swTBlr/e4HNjV4cs
tS1IpPYGlxdsS53JGpbzvtpyigX4hYjKS1p9inxBrmRBHsd9yLFvj7XTTwWWh1Fd2OuszIhZiiZw
nYvrtSaU4QgkFVDWRGSLKpf9hLcUPJLjeVW9mxBFCl5lpcsv6XidzGBwFrz442kuVwkoIO8ZQL0z
wUWFg9UAWVWp/rKFCRTOk1EFieqqqU5+SzzqpnKL6QYod9+O5lMpg07ltEdWl8iu+FsUl9xDKiMd
dyBkmGGOH72hQKPM++HRNzGPMDOWfMX12e2jl5aURvR5licU8SZd91wqzsShp7Rn8JaRmUwUM13Q
9FGrCDtu2PVcp7lAOPqTOLkRDr49UOJe2DjVJhGu1hVd8Aiy1+ZL5F8ynOKFjm4LpyQrWuBUDcNU
PQeQFfyQT1AOYWFPlK0PNat5tYVV4fgwnYZfgCtUZuAaytK6sYDNJSoLNVMqr70RsxzybFcgeId5
myAkGUe9ItkzHpOEMjayhtQV33bFZuqJRGjxFr3HMD+gln9UyDmKuDJRMUR95L6SJDezP0zbSD1N
WZrGg5ZXFRU60GqdPtvZpTh9Wf1M8UQBI7CttVIdnIRSS1REqV61RBL/5XjHDJKqOgWFJRojD4/2
X5kwjQWj3IGEcr6kjp2DuY/Ly2NPBBVFCGAbzgvLsF4zZiNDy4zkY8QtXCQAyxyotjRWSmrzHv0J
zazWuVlMLLGcROA3uYzST7KQgpDF1iZnNkl2N7wGbnB/rbSpPy3AXJ3a0G3EOBSYpoSRdaFWhPEO
6M1n9ZXjqPtSKuXXSWK1ZuWuNs/tKARz749Bj0MMpboKdLIoYzX3WWb9gRxftDuKU8ODlm6MK7oZ
PywyYZKbYkSw8sEcqNYa2sGjiOLx9ag8dlmqMoKlTCuRDC4U5hcxfhnkBY6EpsuGuh/UplpnsNSe
ywqjJ/FUe3DXDeygqbvy5ZCy2YQVI+SecPCPRRc4HH1hmHXe8JlbQhHKVTixuNktljuTwV+/xxuq
pfsHhY1FH+a+egllNPvBYboO2E0PIJfYsKlTsCGBAvhv8iyrWqvsDbYIcOX3ItSIjh2C/HE/cUgK
RUxiymBVBfZcOLNGHShoXbGSXnv8fVvZs5yzsoLy8C3B9BAchWewzpNdvlLlo971HfzyK9sp1dYU
F/0cZmaE2rehqWTf9Ik7toM4544w5nS0i3f11P+huISaiD/atld+krwAnmfrS26eN6050ci12iik
f3ozrcemZvnYKFleYBePCbpQcm3zXGsNOX3p7X8IfhYi9nqLA7iJj8DXVri8WD7hqCw8TRGb46L8
WxmycIadKM53JRRMeq/+a0YGtkyu+yVd9M8LN0Ia4zyfG7rOTFaB+xXI9zcYUDoWGu2MJhY4WBPc
ptFXVDcMJt02svh6wpxFUXlehPNtF3uBt5BmpQSNLNNwuMN5a5q/HE1oORBczUxf26lIHyjEKBHr
DPMDeE3yXjEY6owHgDfl6YL6OWuJ/uz4+thZ4AjyHp/+5WXFnGxmptWGa1Eocd1PLdhEZjZSLExQ
CDO1ObyoIIlUBcHPo8+Tfn0SLkffG1Wcpf3pnTnjpZwflHDgvAo3shuZE9+CuDF/v6We9XHggVV9
k8najZKXSsoKs823rV+YxyFd+DkOzTOTsYI7k60Ct6Hh3W+FYHuAkigaF6psGiEDDJ0AtqbbwLUH
PzvdVVodHxtdeuhSpD+aumLISwfqN12LIjXu65Y0cnCs4zaAT4aNdnQw+10r/go+0E3/A5baP0dE
UNxaja5S5R8bxWVYtX7Q4dwUy2sZ2Gk4N6VEPDMiuCHJhP2nuVA+/fhlZYek0/4DXjNyFBXIO3h+
mCpcV+IRbG0RC4Ku2a+BQZb75eqH2CXNpy5/Mc97ayGlWaIH0gwn7Mrk3FespQwUnmhA10TFlgQm
S3Q8T0Oc4DFBMQvoYFf8v/fJFTtOkiRl8cULwEsuolsHw2nz6ENMN4z4pp3RdfqlYk7e7/unYtgH
S3TUhYXkTIDiW/vPrn/gWFSozkVmBg4mVGBA4SNXcHpGSybCSBPQvRINAnpzIfj63T1EvshsvLWD
amdgm06nw+1ruXbUzGF9fubDr2tY2zg6xvK/O8ksYtu1qb8SsdttkuLM1cIArg8Kh1e26dAyjJNz
l/ZmK0g09aFAhWnKN6f2mDASDWVPAEqq4cyBPdmFXCtKTT2Ncbiy7iZEthNCl59aXQ3Qt9vn+5l0
boWE6+Ht+kn/cmLODDu2oisqm56IvTzpA2O7Cp4b7llXNdiJRuDY6RhcMSpESAsKF/SwCspj9+/d
J3eFf+s5s9oJZxigGoJi/96a3BxMRNZCiafZ7tG/MMpXV0VdrPC5WVDoIYljMhbOsjAJzPgISUCb
krxsC3SDa95PiW0ryPpsuNct9xfJkusGI2fDnJBidZYQCRYkGrsOEtaTfs70Cw9pZbrVJKSgYmMe
4ierF2OI1d6w7CZ7jUWELfe7osVQSuNa0aadycYaztiGkhUDJMJk3SlVCHrUHQMVqQXLHvnxtmkx
p8/Dr0Kbr857OofDDPcx0AHHYtsXlZDzSn9DiConFGRU3jYcTEvDIcDoEmlBq2NErafk5HJMv4Xl
zeCZRYkLG6qFN2+cPN26vEM9Jh1FSUkDJXyD7F4kW9KvChADJGP67cgwk9Bv7vKdjt5EseuI9zdO
KtCp4016QquEn+WZiEQxmTWOuDUKGNFmLu+cfV9MnjECTWLVZfsnplkdzDJ9Yw+GxANUOuGN0xWh
20vafhwfFVjZxDDzsEGOjxoNQ6N4DWl/vuyANGkLDLcNsgBAsfhMbc4aB7LhWNfQncZcchzJUgfL
z+XJ7nfZZ5NwHiKMNdcVbfppma3x0kwZJqyeXLGELzowuBlL6+kwpv1iy9fCsH6MCKKohTiHWzvM
fuNmmR2zWqDc00PbVazxqMDUCQowh0seaQ9k3j1jblwdgDOYg8zyEkYdvKrcKZ0KYe/RVCeQO/kx
gQ7HOf+yZR09k1ff/JFiMTAV6qdlr16cI80Dw5BC0ugB1fVXQd03P4/Lg5fgp35IbybFWgz8N0k6
BauSRgMTUKMYosRcvjw7ueokFBrCHO4GQoiFx2EHrFEJcIoTu1x4JBf1DbextHhHzY99hD2EsvHD
GY52lTkdwSAZjlH0chY9KMkplqDxjKJUkIDNfkg702tDZnlidnHUlX6FgfVdzl47h4lsKIbgwD3V
nPEMrKvQSc5UKRcgFgehs/92zbYlhvngQosEe/pPR+/y
`protect end_protected

