

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
FWJUwQjBjmpS5fzHVnupSDdqmhC2OFCDg+mGSU08WuN+lNcAeoJYKUUQnaRbuv2FH+Sea8YzbrTv
KaWZZFlusw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FtX9k+Nhr04u1xwEhivd/iYo7UzwiRWTKKkDUDMzXTfSnQa3202aN7pNreKwDtl86B2aeUD9uhoB
uyqh1uV/vjvdtALRZfaugrlTApN+HCnk+zGLSYvoHxa8JSj3xG/GUae2C2DK9/DU0tO6r2Rr854O
RjsemBgkTRdtQNEFOrY=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lN6RxOt4Q9lkXDV1w2WOP4ecEiJbRxkZrxzD277j5dJHu2HqHEP2yB9kJ7DZqiaO/sNnqSJOAxLR
9MF7loAm7dO8RZN7KYbrp8qgED8IHsYzlfwaIQT+CRPripdqe5noccULLbeqQ+9snazw7uNWdMb+
mI4OVjgTh6MUvUKhulo=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zNd88nG6vyShPZz1xT3YuldJFZngkUv6WDSwHyfJr/r1ZLWP6fVqJiMls8mabWQfq71S5lrhKx1e
+o6ver213W7V7sCmOdLfbpHYB5JtqcOIA4WW9k0EHz4RiY7mOxKZGLdrstpLZv4lRs1HM0hAB1dL
s1zREsNpPZqUxWkzZhPtjHD4HOUuh0wGZPmPkvbFU3e2q+Jp+nrDMvOj7DJHnAp1HqiFmN7WwogO
da2/VPgL9vVF5qQvTVGRa5NkHg/XbyRX442hRT3ozJm1tNBZD9uOaRuoU0F3RVqEtjQPFS3jp7eO
gRKtaFU2KIhDAcyYk/LufyEQiOFao08Ea+735Q==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DTIVm3D2Qg2CJm4w4QG4loWB9rWRWi2FI34aM44klha2tzHLFHO/meqhDD1lvLjCqOJTLU2M8Pma
8zlu5SCg9/gwkaxnYv5mkYWytplbO0H1kr01H1RznP6MEp5DoUGyMpK199edCkwksrPmNULxzehX
ky8Ma7RNyOs79sdLwbpKFsa6XfNLZzxP7X5xhIJxcAZZnFFNZumYa0OykUZgtwKuPz3lcKdMo+zc
HY3p7u971tIRBpwxb0FLmBRiBsEmFO4YoUsHGNrWFmehQwXP6wANiFPSayNMPBCH/5hETYi6op1s
nqwwYDcYawr9/A+xGHOb71RqpqtVtWgonq3bpQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Sx5PmlDPJ1RXJSuT6bfbdeQftlN4hz5c8JsYQ/QbhvUbJ40vuDYLpROJVUIYcSEbeX6IH3O18J3E
j3vbfDu/NBXjozPV9IQPyxVz/2wQV/VSf8xQnqFFQFoj3HEAB8Jwq9mM2C/eNWrigp7i8lhdPS+n
RHl+JlINqid6t5hw44UiKqWYZ4QHz9FNP8XlBPPsE2LfTx+vNn6WfVUySiPz2j+QpxMpd46CpsKe
mWIKt+aiaIgVGz2HrsxswXrbZzLX7yueyv6kErZBxbndlDXPVIf/1P77iCaF8g+Za/vI0HfTYQKq
HHlEHnUZpeq1j49KLB5KljK35qYeXyNgBxfcyA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 122928)
`protect data_block
qyvHpc2H4aBJ6HFAzZfGPFKZtuPyD8cS9OKz+xpcvr4vwlXW/jMkRNvkgm9HFOPESM8yGX8uL2ei
VhwMKCgBGTEte5xVAI90nDxK+UV3u4lg58ENT7aPNw1Y0CwzudZxdnTmaYzu7XJ7zANVuC7xnUDW
EDjhLJ1mRhFUpQS9FEgZfphlh4nPHhkWL7iBwMzoTwE+OHywLYrjkYQt5PbTEr2ylUSFYORn+Noi
efcExLTWUpuSfthSCEkjurGD3mfWx0Zxr4bwDSwU7Vo+0e4lCYR8DeMOnr3SP+kkWHNsQePZt1fQ
1ifkEp90qTaVttwrjHrFY7KbTMNgHCmJHl8hLbkWRcwcfPm3I0KAZXwqY5TCwu/QAIHtVJwvqIYk
xaBOZVT9LO/ircMvhvtHp5IqCtbwAnqAjEVtsxrMV1e2q6pA2T1znn2PcySqqCOgSr75oNGFlYZr
hz9/S0ribbI9nAUwqx++eGIrumF8W3zn1leofrk37CXWUI2U2KaaegJ/KbxDs/tuFkyhdvrrKwDj
M2rlAyXEJ4MPY/32gw1yvVyKRWnfgony0GRUObnUEKjptYp2ywgXSgM8RMVg98he+qE7q+uEj2Nz
ttX4STBT8rMhaSiqyPf3XMKS+D6nNG6cxP3Z5/CtW0v0LkBvzeZx/BrglwmYideHfq1Cepuj3WrW
lbSuUk1oPTyos7jDoiiqJW875SGZUs1cA/IzXbTzRP96IELm/5jnGsTpkcPpaVJ831jCITRwaJE9
r5udXBKbSsXXgKqazKqKxsT/urRSCoqIfFaQMRQ4QcJmlGU9KNomAu4smfjRUcBwIgAtP3+H3znv
uxskQd/GDxWROAgVjLPnStETUV2GzvpMkyw5JMp9N/I4yYVhlcM5MMv4rdVLCi8qhZBWb02B/wwH
MOVHk9qU6X0MgyOn0CFif2Bc7pzPh6mmy2zo1uEUpti9u7ttgSjGdtbzp83xg7CD9wagobOYTsD+
yhb7P9a5L83cFUrEWZEQpAoPy1Mu7udkDNtJo3Ocwna4hJcRS1bG0DTwbtogVWow4qrNSewddn4J
1xquWOUB6tneLk0Okrp4XAzQCN82V9wke3AYb/VJs4mZ8J7H4NfSyrobItMV+er9eF9lD/FijTw+
zTU8wxJCXGmWoJdSGp5LpAJKVtx/mibK4CilaNAcFUMQLNGqF4smjy38FbUY08a6Zv3ShaLsmwiG
KVLHmVoK9exzpN96/YVxZs06AegMaoDzaBA3albyEhCzNzljsoQlLrc87cJ/WLkKuDDhrwI40wa4
uXmmwpjZas9O3sZF8Dd0VzAb3Wx+7e4m8QdeN7AEhV8aCIGB6KQ7oYxCozACeH2Bitb6WO5zm/Vl
RWEIgXUk8MqgHY82eMPZsWApakYXdo/z6+ixfLIYovczBrJ4uU5BZ2l7FM6KlbOOp4Vz5bbxm3Qu
Ev8VaEYhedylIt9EVOp3gutiW8uwUnMsswJtjt1MyMU+ets6+eVVjh8Tp7dt+v7ZIPHv4AqSiRaa
Ozjo4n9IwhQkug8VJ8Y5BVHQkB7x1uYmeS/NPQ2DmlpvZocnlYeNNH4Adqq9lnvkO68XHkwcvWPu
35CgmDIuDBDjm3akA3UcbhbtOK7MfX+6DYFTyXV1mHXPw25n7Iq5aiommMRDbXoTHq7oQRKThiNl
tf81YjZvNsbb/7kp77sr3WJXoxZzux64vqY1rkiHoZcyUt4ADtpNDy063o3oFGDM2ylneWFoYwHp
k8bo/Vmh+WchcUYjrvJX/bUDXMCOIbTtuPaSWtwA3sVzK6iZOYo1HLqJeCSWX+Wb2DuvC+oCqcWA
BQfNjFtD8utiqAro33tpicVFwjRR022OfIafFqU/efOgI7VIWPwI64B3wDuSGSHCsLMetianLSiK
eS9s6gZkLY3QqevWJlpa/jXbiEI6swPmZUqCyH52roS8g6jsX2T4laJwuaglbxQn0xYpZYySrLbw
gEqdFUwsHkCUMGDs9cU2T4gmx+SeKyfjC7V75hjMS9SK75+8ZM+QvsIQQdFhsigYoWruaxyMMtn3
TfvakdzlUhFyB0dCvBEwkm2rmfZOgAhhQCSsttixG/qYMcp45w9rVVp8fJJB7VgLv/ZOnXQXJcFb
c1XKCkyKASQKoAP4vbOH1bCjv9hiVZsn4rPBXgXLt+qmi7bdQGxeXbkz+kLZoBl2OROJTMWz8HdR
/Lf9Pv55hGaaSHy8uvCebi2t38Of+NLPzCvPicImM4vTozxor/fYHMCEW0Vnr4WfVwyf3brYUwUQ
t3Mb1LGd9q7jQPOe8EZmeW/TixLGLKCNo31WlLGJIyEY8upe7RXROJKH0lxIzM1o+rvXHG46V/n+
HbzXRahc9uzGx8RLqZNihAtxBzvKWslDv96t+s2AYHk5bih3Dgb/T7cf9PsRF0GC65EICkHrJhqg
FZz1cQKn6ySSOnYuc7H8MijkCs/UKSX0YIT8z446c28qDWWjNQQcYixkoWumu0tbjJEGDbQCrWr1
LQCSZdLnkNwplqlrqOezddpI5zMNdj+DCETbpFnH0HHytU8qwuz5V11PAOl/ZqEN7a3J+wqIEVFe
/sfX/5XQtWKXPM7g/MuILraQSYjBIHRMecc4BAAL/K/TJxoZs1rbo4Iw3tDqMffqGJ4wpMKQsMyI
Op696EFbMitBW7GFq2uG0oC/P0xaSpiLT9Q0fwjVb5TMRgyhKX/F1mADQqWD54L2RCNvF6NqOaVr
K0V3ohG+OE9p7u9ZUB02CJGb+zXGTPEfrjjXPBe66cWdRwFDTql4e/EPM60l+rJKTNBqt7aTGw+H
peDZll6xvdqR7ismDQnDGG/C0ViXxdjtpOeDg3VKGQT6gVip9VbSdsyYsqqMn30tj7FM9hjz0o/p
i7JGANC1YtKAEVnAU/g2yCyPhbaCRTLI35XlDAKZ5PYEKg0GrE6lwv16/LPwOJnKi4YbXxqG5Gjx
0xdsChhaoquurmAWZF46Rz6I19cDdcF0l1QU0vZE2+pa9hJmdDExHlst3JfvqPNVeUAC/4Zt0fAt
zofQz4nWhhFe760iVrLKEuBPW9XT0JtYBilCH16PIaJ2ZG6NdRPTO7o/qgxSBJVTNYJH0SA8eUyK
p3QwUMdYl2ScAeuSklMSTPc9uowMvHuG4R061xVuDAb2Qs2E92T48pklwJQnm7wteqXthm2PJeND
3Mxh2D/d8xElBBhCsn28fUKFH7YMxZqvom6vpYjmU2G0UWZ9McYMzodXvuvsjl+rVdIqmZ57ukLf
jUsbuoINLy06wglviY5pU6jRUVPyGeGDGF4uhFgj0IoiangNiJRkfFT9ckt+UwzHRuiRS+KVL4q9
akfn8muy6SYaJD92GL4RMBx4tcN2ebfXdfeIbNj704d6w1CTzqpY1SdcTVeJK8O7Q77aPDgPPRl2
vHz6FhVQHXTX8D6+hTpYimKDFD8EROTJNbSvGrkRjZCubK2ZU96W1QJliHjlWR5IVZ5bW78GeH8g
2tqTknRpRhRBFgDrfxuV/EEZan9P5mrlWNnXIa9SfrSbpZ9ewIoGT90NvTqZgXogg+ToHZPGeI6k
h2gOC2GZhTUEFwFF2XiVFbkgCVOqNvPqbKX2gtceX3lbKD/AWNg9Mv1v+nKvwc1G3IWWzHajX2Qu
Np++4ehpSYhDO0HlduJIWqXvq+415BqUTGbFFrdNvdhFV1qgUKoSKYhvLxJMos4WsRtMJO6oombR
afPdHlPq7t6t5ByEQ429wIRAwPt+TL9DiQzGE/Aq9ZZQxMFqGYWayBEV5Ra4LypZx9M7hkDImsTy
BD36qJN8USRdmnh0lp/hyzm+a6rFZgl+cmbAj3e1ASBEIHDjp+vpPG2J4k5fAJwtTwWxopV10cXx
r39wfS1CX14agnGUTUh7khJhKetnpBtn5r8xfKEKj1HqOIWEeZOCd+k58ah1yR38pWYa9Ki9KoH6
XG08J9xJoLa6y9Brau+l1+oAO6hXaE+5uus+P4KCJ7bbWO/ilt+c87tXIssjaFyze0Q+JxgPxHXD
OUKmSeTvJn+Juj6oSDiN5CnMARvfJBMIE848wYIi+Bzcte/9S8xm3ob4Nph+qKBDZWRGrfCI+XWV
/qyAmVyl9MVyedxUAgS3uPphjEVqBYL5Yq+8+oVJtFY6WKpJzoslt9sXBOcb6s0wFkWnaxxWkl6c
QPQC8Rg7UjrheAhYgu/YIP3UDX86wNgHKDox56hiC4+QwfVu9YwIwVDqByPQu5Zrb5XGcrDH0dmi
HBs6GPmpTGbVzAvFYPT1ERdFhnj+6J5H5Hy8Tsp2XFoJ73gG88Tnumpc4iywgVXERJAl5rNejasr
PKAnEj31tSgRs0cCU5OUolZ1q/Ua2mYpFphIfsA65/Zgcq/RDqVij866lv+QEg5kpIiQIODx7vF2
iBsNjbijm0FGpDzlT087odyYApt4jfa/rWXqllOb1bPP07ZAOhJBe+Dw0+3+b6uWkKr/PYrnQTwj
rGmTFya8ekbFm+NG8w4Lzj61Qtb+6D/QXcI9vhZ6CzsW2lkXI3jv18A8aZb/5iPOOkrOiimqSsRf
AgTLCLE1vLZMn7rmh2S7yptdIqjgNlqkP+d/N31Dh7Utar899+kq/PQh6+vXCv8IrGM5ycG1FyZz
ks5JYLsajcj04XXeAuWRGfubAW1zpoFUJS/T7EI0dcBHrYvf3JR3opF1MU2vMuuB92v5m0BFE9vl
qT9DSmiqPU0fWre/umk/WqFqqbHS/p06ID1vY2Sy/+jlEAdmstzmVuysQ0uq2gzfQ382et+hLiwl
fgF/ubar6pGHrjlRw1ptFRJHzttKb6ASQBPGrDB72ewf7XIFFZAxx8hMX918/TcDPUfF8l7Y0d/R
UYnZ4ZtzEoyAVQH2W2f6Nzn5SLVC2wUB2VsgLuiB/ruGTYairGF1Awypa9OCMk6udHbvQqzdpA1I
28qTwZuOGxNZvnY/fYde501PhTEb9MsTBQNJ0towq+QBNzh9ydVLq91f0mFMl6KSAkpmnfqo7TC7
dQuDFc9RaD+u4bKnk0GTpfG7E+8qi9sOH6RPsd4T74QzSY1xcZ3EydKnh9POeRu9tszTnd43oKvk
8l6HTpYRp1GPASB3r6ryUtAZ4hOZ4VGXDJCmPQ4KZeqZALlx1a+aKWcc7W8sYmjDkuz5GY7vktig
1SHY9toixfOGmz2E7qL8vSsEINFnHGcpkBi6VguFV9fz6rh+IGjXtcUrUz+Ja2lLTflLrywUTuV3
adF3vrDuqBZsRkiN1/1k4dBhWMSLRF4XmrqNodJ/0lFaB+XC5tZlmtTYFQ6RSjHA9CpAYxkCC4vA
IXny+6S51gO8Z1op7ctdr0knN05yIN5WBHgz3LG5vxcHpc94DGK2u4Uu1vCQpScF5aPMFXonoBnw
Lhh7eTsoQIyb/4qDAFPdhQ0yFMRTXyE5qfAVXSevuw2Mdg30k740clPsoI8o3wzUeNKI6U5y6Cj/
XJOoNtz+jUH2ecHcthD3H+0tYVpnOVrTKqJTMXPP1TJR4P1ePmSNKp4+WC0GW83gLgveaHOG+5A6
TOiB5tc1ft5lYrpXXtLxZ8ZtCPoWm6Dg2lU0iU2DztxUAuCjx6nKLmPFKjaBZuVMGp1LsZa55vDN
B5aJr9hfKp/YNl8DIgkAwTIHpTcfuLMBunDdxPmQx/nzTnPTJR7XkMF2uUycUFTS590bp0gbTHDW
niy0bZj3wN7NgmlQnqeE8Aj4IzaC9UR4hvhWHiQt1/YpFVOQlC27s3YWwGE0N1ej3rqSJZmwIDHA
2DjIV/+MNqexyKlCdvxodDW0kjsfSQ33XVNB1XlEXjL5Vo1cDYzsFdk1njuu0fjmSzOeESwOksqJ
c7G8yUZx/JTdftDqnCKJs/IAGT4OKbnxPz2exxQXIKXaTOvu6U1IjGaFlNSq1aVV500FcvPu2RYo
WXguezGxGfeGllksDs0lT32ZX2W5KMijQc9jAbKOyhpisFqav11xkiLt/U0C9IcQLRO+t09exxA4
Ear6svySeMyBzuOCQD4Crq/mKUa6glH7UjjeFtXphhQjt9tjEn/MUB4U1fmxsrADEMSHGlgcXthU
4ENDDdmIqueHLDSymwNY1sgq5KLLvswUOWmPhxH15h5OKiJo4zDbKdap8DYnTztJCzMKJRuVCe1Z
0D4Xb88Eqw3GXE6LYxf0m0IAHReNEkYehDfRV5g2f/TuW5n9UxpzG2hQOpXcSEkqzYcmr6OMPwz3
adX8IHmX0PvA09NHZMUhtIrHKMJ+/xZk7Ur/I2GSve5HNjrk2BOyS9hyj1pWosb3HlfDCRrkG8jK
DyAcekrrA7+6koVhTOLIhwbNJe2+cvxboUbNd7zjrJ/8eBbCE4a8RBGGMp1BIisvRNi8Tc6A/Z46
beHysTheL4TzJ8bn5FxDrdZfrI0mt1pQMp8ZTb2+NIl0Gg7secRBSXWMMDEdnWDlb5mCX9WRjmB2
Em6yc6mV48uq+1X3/u3q6UvzDPzTvHxlF8VmdogX4COEXanwfZhS3+9J8igtunxx0VDYMnjSK73f
Hq3QW3qG6WNX2/wQnpa+I/62PvH/m2lsbs3JmEw3j0UfpJGle2JQ3mb2Euf3IiBOA7qDj5o/gQru
Bq1RlDxi4JnpQeICEyxKFOWs86R5tv+zmG7BM6dZvDetBy6tV/ZOfj2302XwXSPsbYrHzJtxgLmQ
jpj3WJLDhtA/fUfi569V8d1Qf2ZkCGysMNoYpAsTfOtyXOTtBNH6IA6nYIRKQedB8BbOUn+KACB5
n3axDy7F5GVBTEGjVzjM0nhoSs4K5WWrev0pHRK6Pd8jnR9vh0iqYX0fzShGSVWSp3I/6EkCc+yi
9RnHaJZDrptjPqBmFk8nl2gFk5Ygl1y0YD68SIw9ejJAa+H0xQiLoxTSJZZmVgzCVXvshuK7XfN9
zBZ8+L1ebfEWgMpe5RocGR+WlUk36IfA4GoNd0e4TeOg9yupjRj2kX6kqLDeVXwtpk33DM+8h6iV
SqyN9zT2meNTW1vIfxGh3+jhwrTO9O4PT3xMs1y3IXjToRDhaGfByymOP0DWZZbjfPSb1KJJpjPz
NwowcuJYsYN5ZvJEzKp3P8sD0Pjo2BqPKvdfliZix073fX5DB14uImB1jt5Pacbej3aKKnOU4zCg
A6EnZVNqJvmQds7XW4iCM/gb1gMCpErErRiaQaC1JXXEmgIm+xbsFNrZRbZGJDwJ6QcfukaAYLFl
x20L177KB4uhQ5HlWl3KCFzYZOe5miYAd4cS0ASPcGq4xkc50+xDgdbz5Q5yxURWQZq0NuRYvfLh
mnGzgtYpTRgVz42uqEtzKwZAfVZ+DWSxJJSznBvNovEmao0B4BBRgw/Qzrp++Lvv/awWIcizPyML
V+yl7rtvgZAQBagcmcFxO71SGmarj6+KgMT1NILtmm0LDXSwqsO38qHYvXZCcbMxkSCW5mA4wwc1
u3SUMOnkurE4PjHhWDmFPHzNF0Cxf1OAkT0UXWkrdEmulUjWtmdHPWCxTnY9oqgV97SncrKeAXN7
vdR46ZE+t1ixzWiD3EdmfofNTWW6SUyRYEG6qY8ydcC39De4PImTgvh0h9x1WAuRDf3B8XGgVJ3H
quYXdilXwj7y+v/P5dyzVeHz5jy78UNTKyFCPbpCm0H7ix19hyvulFThmcwayVvR3z4rIBNZntwu
D0VQK5jwWh8NvNt34zLLYDbk9SXjJmIKp3KwVKKAGpnVK0EmvWCyfwbAAQUGUZz5HSbcEYfIiKUm
r+vcdqi9r6eOSZ/Gky+mVRt+QHkUVVGL0oGD0qlzHG709RtSLX0Nd4scigHgFYsSKhN2ynspUTKM
3OXc/XMxakAXh6mfJKRSA0z4K4s9WaVmNT0VXGSs59j2TyaqAZJh6dZKwYDTYuyja7IQu4jPJ/ak
m6etyaxPcDfUz51DPCzi5P7klHXx7rW1Q/OYenPeMn4+ua5PvAuxf5RjWmPD0o3zpyt5R0ZgPFTP
7LBGl1LRrixGgfxCHXuQEHs8avfhJAnnq6TeSHgUd/1pEW0+cikXCmVSj6frelvVz6v/1uuEaEEq
9WcHjkpnF9GNNjQUJ6kTx8TM8qCX9OhKaLFan1t38oZXQNmQ/Hb71RiGu1TNu48/FlW1oiPdY7cV
tIt06HL9djbjc0SQYQMXcj1EzuLVNd6ECBIozrp7detk3PYvlOJZR5umEHRQWuS9yO3KZVCjjrti
ay+JRtWrGWzqG89Hi+1bi6Go0YRq0fbpjB9fT0F9ee8goU0vE3RYvoG/Kz3ApbScxHWsdqHA/iep
YaSjgXtbTWrDQ4rq8Dw2CbUrFIq1VrAJ2PaV2p+FFxVSoIc/1y4/NZohSoNTybgYiYT6mftNscnc
hTg481GdiTsGnANaV6naLm+ALdwsLt+Tx3z0CCSj3+9wMZLusWQn7i6ifHxBgLTQLVemDHcDUT13
YuLDDy1q7gb3F2kdlHP2e2pvjJu0d6M+i3esAtEKzhL+ygjgP7Rqv9RWP6GKF871RBjFnMuPvV6y
SPFdB+hWIF2wOEqOyzFw/jo91sNsnjNd3/JppTyYx7uuwyGJvKqYDoVZGlQ5Tumi4JFHUg8XxRYx
osRuDHbUUf2rv9UIvP4RdAe6/7ZN1AhIwJ63ATXOxDBJSsfx0X1DgKz0Z5IrGdqEkEq0a3kHE/fr
8QJPjkm89xZ9DAY6FklUxChNIyBvu7HDBSwUSNRbRGq3SCLARxlP1df6cXrTeNFnThooCHTJty1H
pvzGG0ZznTMYnk59TD4u3NFXOHkPKh1hGDgFa16CKCYVcxXDpixxZteudvDE3L6Zv2NJZDZqL5a/
9XUJxZIbqyVMYxT2bKvyAftNG00tFU3/Dp0nMCUEPbxXsP7oNUvT/jRfzVxhjCrCG8/hPQfxhRCp
syToeZjbk3ebt8VopuV9cU5P9edG+/dAgtEEx4rfd1E5O3gezChflQewqgBwTJslmZGRvHMrVYeC
D04OAQ+/DsOgmxeCMtCANRMpVfcygOZMvFmrIXIrSWPmdIgaNm4px6iR7Qk1hZv+KRs5lhF4uJkp
Qyv3gJ+BT5U//lQcz1ZtoXNX+vquGVU5VY3QHeg4OuZGFjeC0a3J8Q+EpZvgryNW4BULiIEZj14Y
Jze17yMk0tq69FimiqtMgRievyVmAqxoWdZE2JtbIZt9ebhRGgMWHu9cPp1uvvMcYyTIwFxNGSF+
Fu6108bwRs56dNXOh8L4uX6tIJzpuHQWqAV0N5k8cjJ2o8r/EDymPd4jV2Vq5eDbNHckuoKJYcRB
AxxrZFda34Qz4L5PZGbZDYreoDNp2Nxkrvv4QrmLgLjjnAoympZUIMXeeqnW37uDQU3MrH2kfawu
88PLJuf4n4VF3QVdrL+ETU3lcGsGNCTqGjlyedQKoj/k5FnqupO4FDw0DD8ZPMjONUIIGKjFG9FQ
xdvFhMoY8j/vmuyIe9phOeoxr8H68BdNACLn7zKrGcZdAObRRLpcT8ANztySPFzs9vMXZzIc88QY
oHpjPiDA6sK/o2rdL2KQFEiwAK9m2WBHhMSO++GW5mtOCsRMkBfbamcurgzF+9mD41pHPBVhNI5r
JZLpc/8E+nYU5P2QGa0vP97cbd0b/+5kjK/HeJQf3R7jXPIo6LPecI/+ScePSE5nPuLpFl4MmrbE
WpWogTQOb6ejSAqIT4PpAqHFdrr0Dm8kkN/OZSEXGbWiyXKN+siNrVFRu+CPz9FDHX7lgiebTqWu
LHtqpWSMYBheHxSoxqB6pAsETpGszn/QG7xyYIdh0KxIiAJHcaHLtMN74ufPFG5nyZqENIvEsDd/
wBzJZ6RwNr6AOVHPzyWQGPc2o+dcHoZraccGlotEvFrojs4UssEoEBykQvI/ISRRGSPkuoCIF4sU
pjhl+Pofaj39/Y2ANMIAq7YUEqu+F9iLGSmcwM3IazsabYxRQiOkQxTEK1WUGu4LndDQQXTSpwaI
w15oO1sSu9nYlapL25EJukj3Qh8pP7A6TOkGcIJ78KhqteXIcC5ZicNwZp+Vji97pAVjOHKDp7f7
1hjsUIMD3oBbjSZuGe/JUeUHVmHPhV3+YK2uQUTM/687IuBG5K7KOH1GkLnehHwBdQ7pU0/+Iz+R
c0wJ9HUHmBt/++z9JHNsYhRSeiOeajJSx096ZSfHALyFQZLtQ3lxXqqmkLYYPsPAm3jTcAK1rxJR
FCEITMegxdqJ5GC9bdtzSTkuwlOkCdTFeWS6oYO2BmB9GqGzXhueGTtX2lK3lFztUNtxJGoiehbM
Xvs8hMOKL7yGOcSaVklVqiRJaxN2Ssoy89D/fbLABvyiJYou8ICBWWdyMSq5j9R5STCPqrY+9GOf
racrB3iNFz64VofJn1ouXwYW8heOcP2WK2n45GbHsguN1TG9luKTs2e0/qcKBDpZKKilR0NN5jus
a/QS9ebRo4P9YB7cWpIeGjFlt8qmY3L2EzoN81x/M+k01N+cuNMZM9VGkFikFMiULQEJ5+Dq+6sk
6D+AHZF1PMjjUXUs14/uKRBjGcK7j1b2ZrWQUZxHBsTdkDa4B+hA1KCKWpG6ychKnLebCnv03we2
Q+V6JwsNSxs95x69GU27XFjZ7PHVhOpoqC8aqlh3jwMj+99GfxT5NpKY77xEiPhrPMc94D8nxsqT
5qUBBXELU3qI+j46nm/UX8bshHJkycYc7iKzxZ/mjRZbe4E1e9te2TKzhzNXM5FHb4jPXsFa0H6z
6YSNe/ycKZhPrhrpnapTR4K4jfNun3ZCoNoVtSJazStH7RhGLNtq+FCzTAV98P8sZcUZyKMb0Tk4
3miYVVH3gEAnLkipLjh35n3pwa43iqEqg4t3sDGCXJHKVDcAgx0mEkrULUUGJ/6Elf9Pehc7jxAl
0QNw+AP6cvvCTqkYa6iJUhEV7jG2Wvg5VMxLoPgv3JQ/4D0n93sq0qpx/Z+frX16WyxPOsbeIzaA
kSa2OvxuOg+dSLOkK2TJ6qdIkuGdReRHk01VU2xV8bmYDDcZQ7R/stKypHsvYrDhZuGIqta0uT4A
bp4BrWLLNeCpYKuNjV2cWWNJzlHF+4KzA6tthi/NN6yts5aXNXTWQeVvch5vzF3caMus3lBBMv9J
yh1GaAhk/Q86vgk/R4cEhGYSlqP+/ujw2CMl0Hp7QAA96b2cZ5S3QrFZBzGnZ++0AHz1RzcHIB5G
XH8E/p872AmcOVcKr42IbzsQrZyr9VzhVmVz7qNHC5zWi/si5a5uw/TK+HbyQ6PCNsybvqASJ/UF
HHrB2an1ZH/+uZ0uzqhrCsyIB7RW0XrIw9GKqOfnQHJu8XdF2+0Yy+0jFzjx5FxfVXb0Q19f4mdi
k+hrY5tZWSA7RGDtBqBPjx1464BC1JW6x3T1fcFyoDZFnTOcyvNqAGhTgyHZNbkzU+4q4M2gcb/n
xMsYx9d2jARwY01hh9YKVCJU7wIgZKTUzMq5nB7VXR1/w3Y8PWNf7FoS2ynEBdR5kHkfDX4zVSgV
vAEyXX3X1+6IWIkIIa+ajreOhxlvRmsC5Mxi8cr2Fh8CLQyRUXJGIFB+UmJn9TSuCLZtJhm2Bgfz
QRVI7L2vijRtLHMuG+GUhdCRRc5l6ARvZDohcW97R4yYUGMW7gk2JS4y1OlQWAN0gIxd2hYIm9Rt
FjR1D8KmOUTL8VNDS/ntRxU5jK+NWys44atALj088jxmlYe/k4zMlhkaJdj2j9u0B7z8c1mtX9hs
BKdXdZEzskPgja0/p/lt0FSMcknP9Ui40rsDrztWgGMzDGglCl7iSuEzzw3Ecxkyxrq/v7UPjZCm
KwWoMnAGi2+7LP8OEcxEGKfqCMae8bW4ho4gmnIbvNjrGCK3D86iNwNlYDWFhjQUHaBmQpNhIt3+
3Hx9oMbjlI0VUJPKyYIAL8Yoc3TsUROv0hFxJqKl3lx3aT5/APqeIyHizmC6FKnfIRPxgz8HfyZ/
H0jSqakAPP+pHqxXVrmohoI2/spVuyJgmXdfDJSqD3kWiAInSMbY2uBPPPzOXzlxP2+npHn5t1G9
y2YztNr12eul/88fLRw/5L4BhVP5nPX8tdTRvalFdcphiXJXD0CfyAuFA5G0V9NXpcgjDhQStYOV
Eu+5UUJAMMeZDhATK6TRVnL4EqRu4eA06SIyFDhDPd5sXg+3cVEjmQzKA7JbY0bX+sDu9cEvlLUX
IfD4WAooiM74rMyWghj5onqgNDflo0BsrxIUEETI+uBOcDeF/+SXRi1p5uwDwdEMwmcpFMz0Kl74
Un3prdteQWjHo7Y4OyEv2xeqPON4MuTKVHQKjffj8Q2kDCTJUG1tm6cdc+IEQjtbOujBPRCJ09T6
nnOQowR9EmwnpiUwZIJ6HdKRiXpl1rp8XKrjaFUqm3Qn5nMf5GTwK7HZYnm6fTxrXgm+hzFyPdor
Jxih1R/KfMHcR7R/mE3Gg0IDZ1t3/IdyxuwSU3hz9OUdZNHX1GRxVc41G+e4ckdZ1BR7VdCdZN06
AstplxkG9ykXv5kMI9xEdxX3KuRFqke+7pK+w3yTdKVY6Tj43tEguTNItB9ywiZI8A8EuiXid5aW
IiG8XctJpUXfskxnXKnF4krf6+hzI9A0rwPXh1X+TnICg7xYeGEHhl9boIpDgmPlWOEdoVLjgUWk
YwphdEbj6LBwB9cH2dnogW9dXFpBhSWXI656TGJbUfq8HlrnRihMDkfYmICpv2Qlj1sOViv6Y9Vz
6Bmlt+v3T74zYFupzIhsW6ufulSDAWoJWXqCoeEZlWKoJT3WgtdrAnXHiR8Sf6MaCZDvY+ixOwi0
EZqArDAOFWv1eqLMQYlf4qPbGn3+hk2qffuOAYmQYv1lXxA5hT5ExgSOG6OiyTyKuthC4LiLgXTH
3XhZcrpshZaQY9Qgl35wRvebewa5gOn57gbF8MPNixvqxeUTeo5ILhwzhzIcvqtT7SOGxh+EQjrX
QI0Z/Py3H4tWRJBkL3LoG6Gb15IG6LaGn7LplNw7f1v0g4B31+qS7qYadslXVtNm3oyoa7HTs7l6
hsdwG+l/UQHmb2MfP2cygPv+nOrZnIz80GCMU4tj+2/UHLmExf2NFknpuE31mOJojIT6urDanMK7
ZFgmFoBQqhYkWuAhq024zjvWu/OU9RNvLoJ6J+IYsmdz81HtCuZS6HBXVyDu+2hs9RNgW0GheDAe
eZCj9d4oRmmsPk2fMwD7b5FX6H8YLncmKo11ohTDgx5IUq3e7WjgXTjOiEXUlNkeBqZ16CbwVHUY
BSdYau2Mg1uoJzatAliu0kb5kmn8T+wtc3octvIA5sBWwd+fj0Y9GVfZ5AeHbClIYSwF/JrRCodV
lcj2UJnVP/YmS0zj0qNzHziWdomdCz41+gMWSuHdSFTEJDXMHyzv9KSCnO5ugX1iHTuxf5KY+H7a
crl5KaucZIcZpNuiz+s+/y0bFWuxt8Rh7jPi8Z9R3TeSfwbAK1m+bp42gvSYeXxtsYgAGPaAGARu
JjbLb2jCJRPOD5yUra6X9/Qk26mkRVJrtgAH3bYWAkIGnMPvt54Vy7/1QAb3o/Q1KEez8KO9tesE
UN40egnedRfDa8v8RwEztAVijQ055+Q+lKf1HmAJTyPLdo5ddt8LQ3w9bILQD72ML8q3831Xqljy
u+tmnWS3H5Y80N0pctyJVvp/N4L8fuKRjZMpA/LHsyzTNHuaXYfg7MPSoefr/KVikKpCJDJnAs3/
KuiUbtDeZyRL7aqPyfRwyvkxDDR1v/nQCO2XzKq3yMa4GFB/BLtjf5fGO3/q5hpzLwehPNTM4r7Y
F7yugsx8jHMPgtPd7EPxmJOQ9KJ1bBoT2dcIRMXlNWFZr/h1Al9OKVkzdDThrsHQOHxvxz8cJrPU
bgnZBJiXyNBc7SR5IQosVHt2j/JeZZbgf0nD5GN9tWgfCSvVrU8OsEXnrfM8CAqpR40AAto8WJwZ
tTetXcHe3bKVMUv8B7pAsIA/EejTtiSrP18PVGDgGZN+JJL+pmNsCgmyiWiz8vSBF3bo6mDCoN6L
5D6vQlRykH/AvfExWN+5AjgnVBH4XdxgFYb6+aG24v5b5gcAUlofRDnC92AYjS7zhxsC66K1SASC
UKMHLTltXArsESxp1/+TRCZQKn1lUauURnGErEBCoT8bvzqnLbTd/FFW9dm33mydB0KXAydDW1tQ
A0om59xoaAmKgCP7aL2Yj/YjFxXbTMAPo7NxgRkCyvsDY5a924FnzBdzeJNLZCT2Gz4+6y9EDWLS
afxRvR7AlOT4AW++oJ85i83WRcphLhbivYHz6LkHb6RKtC0q9ZT/onJ+4z2q7EU8JwLNYVvUN8jk
h3k/+Jvix35AjJMr4KPc/d7WpIK/ViBP1O/srU/Yuvw4TQHCY+LM5mOR0Pj1d+NcVlFTbmQHdDui
A11y8eQ/I3OHhevCPEtDOwWPRqEV/k+MLctgmABwQiYPSDGHyiUacGFIOOTebHa3RTGFtyD6nFNk
rg5eZnfRtCP8YiSmA9UpO9iulBgiOSki3MiLwCBFI+J/GM62giJ/ZqeBwe5ltkOd4uTgOxOb9fkQ
QjnzNbykAJ9aUu5ip5N7Fjgbgzu7YaWMUncQlGhCDyt1yA2zaoiNBB6YEJrS1wweRHpf3NxnTepY
wl/HB8x9rbZu4X0nBmAnzWlfJY7Cxub3FhPa6pbhuJO/3rtoQ6Xqg8G1v4cLKRf1uEVdai2y1Uzf
zTFvztCLGc6walNKq6s19nr3dYdXLKsT3ywtD0naZ/NodGUuwRleWkP400QfHta0N1YVU+v2R4SB
M2gguDZJqFnfBiNQ+R8USXYDl6h/YYvH6HaOAK4nVr1WfX521yKtrzM56IC1sz8tzGR3HC7OXZAz
H0WJwLEZ11LZmKhJALPLeprdM5qmbnorvwnfw1743W1E866KMUGq4IgUY5SACGu/ccSOsgwuRHHv
otmr+ajGtl9G4aGcPyAOPBvTsbfrCsuwsytiXmImSu35PzLfC+z2h2Zjxl2BaODlUzaZ1jDsOnVd
HfO6D2SMdnypsab7BO4Bggua7S15+lK/JOthY7s7Vb0KkmQxY88hIisPLcffG1x+aPP3IKHmm3t8
B7ivCQdTbYoy2H8oM9BukTd80H2mcCytJme/8QsqYC3pTns0lTu2gN74vp0xiTginKfn9gD6q4Xy
TWvflBwXY8gvtLAMl6a9oZKXAuGtFUFxnClrFOXE9vcQ1e7YuY4bo3a9+N/K63lOVsEe/yHK1mJO
gfONSY2c5WEVzAAtZDVR6y3nUxCF10PHvqP0r+ppJuehdTpzodiHvmoWwDJcHj4JuaGbBF8k0g6R
51GKuUwS8cn4WCUxwzjjOhUOXGYxTYTkp/Tntcz60rnE8IKGd9GBtScRp3+6kFNm/dCzCmLtmjTz
wgFS4+QQ/idBbGziz5jqNQ584QzmGQG5d0e1PE/whOLoJLvfILDJkGz33Ao7OyIbncrk6HJ4Gr5w
8WYhl+hHK5FkkUcZNf0eJgF6odtWCGq06j35KFf/g8lvOPLM9aCI24BeVGw8ZXYNSpcXsOZPPo2q
tko51Lx4alCx5wtQWWVcbG5jV4ftn/MqWo+OMVq+c6jZStC4r0bG3eMxvBKphkPHLT5fdljThvhN
S2PnrXaYi9xoLsyqEGvkf72IlKc5FjfdXE8w4wXEJR/z7HUmMX40nSsv3tceP+kIGzdnhHTazQXZ
4Uqn+KpFLr2H2IYMWWdCRv9Rf29qOz5LubaBawmu3Rv14eNF/VyT7rLbkljVgQ9XM7X3QpMiGBpy
NnKU0yiIaVb1X1M2zzArpxIRIkf6lOnSg5skxtC0A3u87Dv93nkhGYD0hlcgW1ZDKpX0rhIVcHX3
ks5B40sF+gv6+i2ThSQ55X1N/RaLjEuvQgdr6BwT8H7aXPEN7BJkqMRLC86zBbPRV2jJRTJY4UkQ
jl/g3FC32kkxvfhBvAAzUeAvYuZA2H0H98p6RhN7g2/JGmBI7JiEjJryjkq0KeWLtWNVMUZzdpOK
iX8mni3Rjj9mWTo+duD2jDzKG1oAYnMK3KfDPTRaQEI8XwySuVvriAG9opGWRs0yrSh/qBG+HQgZ
EpYPe51hSySiMWSmUCViD4Dj/PHbzOaflmfcWSTBRqMjosHGxy5bVKxna37MeGIMxvXhjGQqz/lO
PK6MRUuNct7oasIoQrYKiEPgIoGFJhgWQzyp6ceyNJcNKWSJ69whVRXZqkkcdJ2FqrvuXy+7HIE3
fE4cXmIdElreJh6KjD2nFfo0jQMBtr2CI210tSlM1ON3SsXFtOG+3+9Cz2vkUGhuzpkoEWYqhVyD
cVATwPw14yXgim1K48WWvsB/BMMk5OcIrQM436Td9tNI19VNkL1UcyluN8b93iwA+lUWeNmHgNeD
TaxyZ7+vQnba8DYDsxfMZhKmDsmGMWN0gLkdVTYQNCaYq4kJTqH+GExyO+3nN+1MrDrtFMWT0wuR
IzC37jYW4cl5fWU1CUUn28kbk/HQA2l5HLfNTeFitLx8DSkilGjV6uoRbcDae7csRCLYzKXzvSVA
CykQgbMn300tiIZhRYfX3UORHQmJKUD0GygnYEV45D5b6RD4J5nf3V4uHPJZ5ZgiusyJ9Q0pApO4
dYHZGyxVU1I+MF0Q+EoLaQW/WjWABst5gyh0tVKJh8qh3A9jo0wdlFlpj9PEUQxHPvq+yoqlz2Wu
t3Ouc9jA1YIyYRV7sj/PoKvY33K3qh5x/ykFK+NlbeT8Dr8u8FcdYD4kzBQ2pvobH/yVlOdqtvYj
UkewfUz/3mcR7fO/2NV1/l4It9K2d1/m8Q3iv7lhJoYuiiOC02cHUVPtf+tJS6NhZJnMvs0gA5bD
1AemV0EwfPZPYvq76ghx5zmfGFtah2LL/0O1Ox08KrnXDi/MLmE0DWV4REX3VC9ZEiaWzo7CTaOy
DSsUrK3UBt9V7x2BCk0K4/2dbxnqqDadY+BCszUWEWkISDan3/0w6VUOd6DZpIyBTW24hRWOfd5j
F+xJQmlRbZPSb0rMXqBeRgFEGPZICuteCb/dH1wmHKtd0jm7153R5m/ojEgHM+eYNkaWg4Nq0KT1
bPWO0hebGW8MIa4+2fKGhjANmINk6nPCmQTpsvJxScOCcbNNnGLLXa6CGVKN1EYVKmFGOloP0g5G
ZkxkhZT+2Is1LW23MKG4ziveQm2Km0+pN81VJn/PLwFaso1jd5Eg5get42ro05NGcV9zGxYfeVGD
JUnlvl4573/XTygUqfDgHEh0Ap2bCjBI7cDuBxEzovZLHcLrI0vDabRJ+++2vsiamYqTgBYU39BY
K+2D+cYJnsKbRh17yYMG2sBp3Qo7MYN3Ro54tHIJ105PfU7EVWcCJhuBxGJJJF7B3+b0tKOwFHM8
KcPc9EYh1t/mSj8rEL7wGftrkU0TbgA0vuHs27AEQQbYFmItVmZCRy1ak1ldHFCTO8sFvCeoHR3g
BJ4FHn3MtnZ3pUm4RQ12QpsBuQh2Hqcq/hId7JrLpuKoB1rvzHyg1OuxfPu1HjNaQWI7FN8Om2LW
UQaTDLv4BXQ+wcDRxRkjruYpM+iqX2TGeaM78vb8lRK6Vw6mxSzYLtOqFh4VWOYcbPua9Mr5zWnA
+AQlWCIT4kYHGQyxECuHOlTlZ9Y9H4A/nokcIVXs1Q7DQZaUV/1reHbHuxa+hYwsYA1e/9vCi1BU
gNIT8o+D5rcODcPJbH3UEm4MrNAMlW1boZdWQ5QOmuaI4q2wkacx/cqyZ1cbtygrV1d/1Hf0iEgH
YIyvELWskT/Sn2qdnCZ+v8c6V1tgvQduWmZhvoHwv4CEMEeN6cGAr21UlwqzwzL9919leuiligbA
uo1ER9obhNOTgcwuTOsDIdQEnnNYfeNJdCqDiUymv80CmAatF5Gy1mETqHqpaczhcvmtBuXFqxqT
IV3LaSYTD1glCtV/x1htU+MINGwg90mgvYiFpW/sjl8uWkWztxURkT5a8j74bIFvXA22cWnYtxxS
PBhua2I/hi2mfFqLVtubAg03o2/hk3jxsmwjAp4DgIaxqX46FE2TVzSkvUPiut2Q/uUWY87+LauH
XzKy4bqTKhCwPSFAn6cwftgk+7jeuzxVnd2pmaMZD8hr0BjQDOL8tpEdfYu0xfQ/kP8zDGG1x//r
dDCv62po7miYRW+waExJwcS435DCGXzuzhMqHeqQQSw97NH7YLsa0o0IDsCZfuvN+oruddNbkDXS
nLzFvRT6qtTsHADQz3CV/yo5x/eo7da5Gr7W+ISiC4eTvNwwdyymrgACqG/Z2CorZW8aoW6vhRL3
zDvgfq+6pliH0D/ioq0wX8mjzE60WXHVTSOhy5gmSNgg0Dx8Xq8ruhRrCdmLwoOBvsfh+MpXezAI
gES/916t+PHnSgQPFBnM6Ue4VPRDCBPSx/7nYIalppqwJen50Xg1qXWc93pibHxf1uqn7qEQ/p+O
MkdtZFKukm6LqdveK8WJneF1mNXT316nr17Lgt1fiJw4C6aFayJ2DzXOBOvA1udzqHd1mQx0HJ+h
32O9E7QuUQ3zkCv82IXKOk9ju07IReaicNbEFw/1Go7NFLgxviKeokCyxUsuloW8Kmk3e84Efrcj
RJDliw/yQG6AuAjh/2RW4dgvfgOFWlTBX3k3WBvpjwUoVzygWKjI0KafzeW1TcePRCAo2x2aqYTh
zi18ugcHC1kwzHLqzM0OpwFaqYJ50amkE4SmtN9ZajEDqHvFhI6s/nYiSCYs3jD7iCqv7CigMaWH
0uuYf9AOLP1aUzNvrvyxCUHqxBnPRp4nDTyO2V8nfWvxoe3k37GJ02V6pB11qOWnp2nSwZBi109E
2AHa+RsN8btMrQtnv1hU65XvFkGGbgAk7imG9UiPssesi4G0RafP7d/IkXCw63/ZzueVQmQ6eG7H
SWnlATlL5y+fLTgkSPmq1eF6QlGh7PDk9mXoHDfY2UaAgC6lCY2zfDEBrXCDtNcbXmPyB+eD3gkL
3Cehn26Ll1ykPlHQjsfJ+EWNWobhCMNGedygcXfii2YZdQ8kuFaFvDyNNQ4eo68CgB9DWZ9CgtOa
0qw4Lwz1KNIcECt4Eea9zeKRk4qncI2Ee+90oewGb3aPrFE4sFR7BF9+MuMiocp6O2b5XdGLFOfE
R5dDLTL1xWKoy7XrTfiHaFWFOClHhSqr3/X7eED4hNxK3SAeUWHXiYRdvRipyAUiesDs9pJ6N1qp
JjUraUuFy606pDd6hbRdP7Pkg6tUmw5r4oevNC6SA09fIRzpmgNf4bNQxojwQCXnQSI5KhXYDBs6
b3bO2G0+UC7Asb6V2lf13eKfVnTpL4qTLkBa4Q0vyrxeRXVFoOydTS+JfpUWBeuy5+3GFgJbpsQ5
LBnrnbiiRhlFVUpwrT00S3DQPSkTBy52IdQ7STNY+xJHYTCBlx/xAXKO8BMizn8Dbx5/xwpsYO9J
sO6UKUCeZoQK6U9pSNWHon7+uoDcgkH6uCJC/SA7mfmOgOnaoh2ly76bnmIQJrABdNt1yPT1ooQr
KfxOIuiWkxT7BJjd8nrp7vzrDfaisZSB73V8Rk/9FO7NzNdu4vDISP3PP5mNV2w0Y9w2inECc2yr
sVSkONUbsP0hfFbV4oTpH8Kd1gFeMOAoe4IngcC3Q07MiuxTl6QcSuyxXNR8ErF2yym7GVc7b8T1
tGnQmVWissZXGK/df92m/6+yihT8zYGWepGnrcjZSqzcD78udRPgv2mUpjLNPYhV+QMk66QVCyOC
mhj32/OH+7dyW9Uspxp698B6FkWQoc0uX8mpOXKyKRFxxfxgJU4MxDP6PHJtUuC7p6WGXCkwLhpQ
eofe34/aZ54iiLHnP/PqDlhqzvQS7mPnZKysWu3mbqlO8Y5xiOsj4Yb8nkWaIbS4x+EUjWwjR6Rg
5FmBw+Tv1rYTy1SIKC84MVPdstrJ7y4gCvAQOuTkyEsdE9O+ENp+kfm5SEudNr8ePquqEKxUs8uQ
0Z8Zqncg8db8U67MlxMT3lCg8YpVc2mIWgxbLSwqP6866xibBZ28gb52wMoxPN6pJEdiDhFHfpvu
ot+qU83xllRFUBrx3g+TflJzbUGkcYb8KorBOuYfpKVARgfI35qcQ+nTuhwHVzUJEIQePHKGIwoz
jgHSs1y0fZdg+Xehrk/nugh12NVoojYy7AZ4OACIGoCFsXCIjk39QdW5kc2iil7mPaSqUZWoXSlU
VQcDR0HLadlxJ+HR5jr51vLHDGxabbE/Sds4Ynz09PzzM9tjmQhHThMfRSYBVae0g7eJmFw9WfFa
fwQZpoS/80UlhNTn3ZiNzVCrjGD8ad3XGE6Q6NilThjTw4/8BC85xmv9wWGsFAJRTjlEJ1SvQwZJ
gMZGIxffjPOTqIFveQzEjsKfR/Llw7SzhZLm6D9GwMHHhJ1xGPZxWAAvr9TJSbRCGBn8uh26XkMm
HAUNtOb8Z/n+AaoxSlp1zdT7c34tFjsGMRjg/LOAYIBNpTmL1QPHQxefBDFNyEx/UOcTh2vxzXJj
coMzIGCfXmdivREkcCBAC/Sv1deVHPj2dOGgQstq01rqOjeo7x2LT/KfPt0VnL+n79dGLEdOrNK+
HXO725N9xBsMdpcjOaEIk/UqOElA+HKFYCTb3rsCYSVDrc6doEWtxVxlgxQwBZyAZMZ0J0QxNIVu
920UHWnSRwnAlzEDi6F+IgfP60jxR39C/YHnEiKIKwKsWvyqciZoV9cSVgwXWMjtCXAv3As28gsZ
yg75s/SVk+qQAoZMkk0zheSsVmNCdZyPJNBBy8lVmJq2x/EmRtNX3TqF700qfylKEGuTSC8xoWFU
oBuPSNSGVF7nhL5ssrRqKwKYLQJhBM/CuEWBsBUK9YODPxEeDUuGzbA1rMooay9G80dARan+I6Wu
vMIsIzi/+UHQt79TCBzWW//j1Dr+UFpiiByyj8mmLpf6sF6PkXzVZEM6m3QbssoH4enEuSEZFYkg
Km4lrP6BghaaTED518Xpa9frxfQIJGG8CscdgFVZs0QXvvOJaVZD8LZmgpbaDRaGETev5+8ZcF8i
R1nbaYNPolVK0dXy4KGoLD5QCDDIZ3FTPsIgYz7T5PRKX9Ixn2y4IPf48LGsV3IWotqNqmDfQdCb
nTzR9BUJyjWAaIORhNkq5H+IDQaMMIMOa5xQazawLJdTxs/w/g/KlCGiCJN6LZ5iFBtsMAitb6ZL
oJlpU2pxlIV1L6sLcz1uPIVJxBN7HVM444dmBbwg//p974C3fFWMrbLm2N1ZuyK7sl/mXsDPCvqC
RvRP0fBVeEybGpHfEIDG+Ca5V+swQxYSgPM01I7s/Zg8ZVc4L7zZSDyQ0ONOCZJ1Yo41TRAS3oPs
D/+xDVTLk+EUdxC35HtOdZbKcu7/unqR/2diNTU8FjGX+b4lPhGsiSx0T40Rhwvmn5Fwpc8/TqYQ
fxveW2PENL4KYcIyOu0ARAnN/jjbwAGXXAKxa8zgIGpFUNReKMYjum2CMKPlCXL9KSisk1x18bVf
8rgeusuqX50r7VISeXWcR9I3Ibm3pnYGmZ04L1o3YZoE3U4DLTcz1b6nQV8YwBLK484Xlv10wgcv
xKH8a9wEOGBM/CNR6EkLKijDLq7PnP5PbeK/7Gz2xqNTKwjZwYSctSvzAZimDTQQpEfoLRPPKauf
3rcsxZ4jrljmXQ2T+88LCG6P1rxMRUhaNOR4n1HStavbk20IK/ABF/Dd9nQwiJFAYzTJ408fL8Rb
FcqRaMpMA+KPtovl3XU+kyMPkipzbJa0DQZSHIeKkxrkFH0dW+PiO9Sn0KQWu5TGGeGWQXWCJ6wB
mB3B1737aUmLfif5whKIUoB0swGKc0FLqzYgEeA48SWgCQ2zIyJtLaSR25PzfFSvYS6bmr5W/s5c
j8KRtzz4yQEj7f9QWVgVDHksMDCtsrBfSTIo392tIl0Iu5iHUNbfWmXRBLnGLsWR1azmHXoO8MoX
KjPSkU01fRDMEQHo46nQvRn3odAx5qNhwRkXFqcTgKg9GLB2ZxZW2Lwx/13oQTxZOkGRIJ7Rpi7X
kesXDyMSEP3gIu8tFUEW4p85JEbMcbcR1VD/3DLVRWlEOoHJd6i5ju+p8DAuO1w/rMJXHtFLOMo7
XipXN/Xbdn+IYjktWh/Us9sKzU45rF++peM8QR5UX0vUo4+A/uieNmRw82UBxqhqa4lHG1upPuJk
sFPhiyDIjmF7vUJGgBgyvhQuhagHW0n4bxHxC6+3zVDtygSoG/rf54gHg6IlCfusEAPZPhP2ijD8
2sI4/3HD6A+wE5DLXIZiwELUg7VGh1r4XoG36K6eQrvhVy9IuiYGmIff4f5iu9AVsihBnC/Y1GAj
rchj3g0vL99v5xexRxOW47Gq9nYxcK7qKi/em66Yw7iQc8aCke3gkE6viUQicCxUC7D/KnkwL6cJ
eiq71jSEyNOU6VnPgDv8DHw3BcbP7VwA3AZ6N5uVzdYoFRukuEQZB9CxlQhiiOLECfu/iduD6vEJ
P9wpRjWIMvMbMfWYuUEWpNx22uiCUu8T0RvPBPg6Gn/RXKllv8pvkV4R4r6JCdvxE5gZuemWtmTR
DcRAg1FGJUdYs7GsCflQTNZP5WHZt/mBH2ngvC9Euv0dpVJB4TeFLyfJkVER9Kfvqx0aJaaWNht4
6YLuJeerWuP4/lC7yorEKBvJ4mn+IUdtqqnmIEgozSG4HgJhFVwVyeoC8p8jjRMKD8KCwcCgOU4N
JhPx9akxGuCKkbw/oPjZiBEORAUxleNnd/RDw3i3UqXai5VWfrk6oSHKLoh3WwiZGDPTaJn3UI1B
7P5aCx2bcTLXocU6AyWy8MLMU5WABz92cPQ8GYia1La6gDzJ35+2cfvWKFOkMkQXjo6xbwBtHZG8
eyiSmhDBLFRzoYpe+9oDLrX4+A7tTnf+oPbG3vrxJo/OR00kklaYFwOgkH7pEIqNaOdXg3R1ZvRB
QjM7mqzeq7xAG+4ivZSlToOwiVNIiS5GmNxHRLMyG4TDt8N5lqQipdErm0yJfVGh6Jxx2eHk1qXT
L/bvVzNy7BEuHwdDTcNtIbE9Zz1C31t+IBq0uOmQ9nKwClWGdis3A0PVGt2B7gi5Kkqozx/BFsBY
k7Xo54VuhFiuj4Eq1d6cQvAqM6e6CPZJG0HRtMUk4H90qwMgCelUmNa23q961uHtkGp52Npw5WM7
G44eEn0xOzL7jBQLV6xnmM1Jbszx4LclHlzz4bz6YnT627AcBaX2UFIb+JNWHBs+0slM8+ZxekgV
yHf2yj4xa4QiwthxLJ44RRDNkcEFNqMvehVNT7RsxRr+f15J5qUzbD5KCjGbHXO1vkHgQLIEcjSW
+BPV8IGYqPTB5DZ3J3KyrKcBVt0Z0HCAOo/eh35JGcKRmrPHs/ziWjyAq7oyU890+/iIErK+VMsu
Niw09N107RN6TVjt0rZIDAcIBHNw1pRepSecXsukk7ZqLgnuxPz03b0E1tIO+WCU2L6E6gS1++8D
oHTuFQxe4mhBbyBZW7fqgWw8elljTdqSScHImrNXyCpkdC/7j57W6JVTBkjXs8vrnR+45KatbJi4
yvrJgeoBOoWpmXErDxkcdVmzFQzPHIM3STu9hxyNLMx2DBn+D0itMi+/A9uATIbPryRB5aCQy2nJ
8xxqHgY6ObmKgn4ZxYQvAmJtW2c6jpbSAQzGVv9I+gqQzfJg8tsAClS6oYgzIM2yX6prxEAEpeYh
xwpfgRIELizRCnT34312spe+7YzJeGGC0u31w7J1k0nF0lozspNh2ToJl1qYkXJihS3DfgSWeAQX
JMQrykcgieu1rRwTnwitgm6L1b+EYiPt+mLiVVEzHGHQhmxeOiI/IFlV6MDBuEBSf9ZYWmETA+JD
BMxlgaSB09QPQetUP5l/TOuf+coECNDc7Kkya+jPlTxuTH5XGJQBKgP3MMeKln2fPq1O0BXUus2q
z9x491ermlpVlAcLwS2pr6xpDna0+kR5V/5MtdVmvrG4Rw+1fYESvxr3m8iYSXtCHQZDKrVvko70
JlzewixvjMTDmMd9EQETB67/iOyPFTrVngoKJ+cifde6IiV8FkYsG2tyeg0iR7pRFWYSt4+U7zkj
xX2XE9YziDemvmquWCaZaPLPPiJaP3OfmKK6cwwt2MzeSZuRq9VJvc9P4jYeL0OWhs6abaah/6/c
s2LheHcMrespKb4H0Cn3/BHJSIPSJmhd86zAMDmY05Lweizpip011XFnuamR49akq8JpPI+E5PQl
r0Z/0OWwvbITR4ZPusBGkYTdkrrVGMyn+xKZ5qpVCKWACvK2Z+h7l+2VGR6C2TQ18fgi+Mx0UXrl
S8gaJBHZyhvN4PlwzuRRUjIkwYQz8lMXgJKOMsDlYAqe82JMfoOmwpfUHOVyIIwHlBdW0G9rT3ih
/r79mb+D0iZjIsThaAGp+8/IplkfE+f+nYMvYIOYmIjB42oBurtYRdC/jCWx9sj0ZtnEv/lBreKO
X2rn9o8CKFt3CRiLMI0gpWckHKwOp0BgooUaa/hDEQvw5pUimbG5qazAKy9zsstcsbuDxnOraVmR
0xWoqaIP4PVwOYcOWvHeWyhoWDSSMVp8r2HmXzxx5V9CCj/QUG+Mh4QNZdfAigaUj9ugbLyOaKDU
kuZKWWYy+7MyLOgzlQUmglfmWLqttpCwRhQczLctCJnSEibVUEhuiecJa7ENBIIcAtGnVRK053oF
wkNSSykZMmtcz8HztRqU7dTvYNyvJjtijZmKH2H9uztvDJbqg7ptIqIyaHZdbFZQ/uy+r4SYgFRa
limOqgFuGl49/5wuqxDYiz+zodfm6P5exfEc2f9CPFsQPJqiiD1k1kEYRRdXw+CfwxY+iZ1QsEBO
uCIpWwHuDkGPaDuryhmf/U1wuyI3YVVIY2x9VIiKOTCw8FwzOaYC0AfGiBJ2ksEyaEM/lPiX/fY4
xOokxHSBfWBkOOldXMxO+00IwY7wNs0sVb78+PMh7PPVooTQCkeBiisNiJBcX4ivo/ic68SpDFNz
iMNrlUMKJtaLQOFyRwNUVMRu2a5bUfS4MAK6Y6vBK5zFS9LmzjveJnXtUwMm4kTjYD+tl7Prgj00
LS7GzDp60Ob3Lh0u2rIG4aZMdce8OAyEm59+1SistxEr19kX2SKZE9edmhQXoMUSiuO5yTQLK/Rd
rJLj/U7U6gluFKb4nJaPMW79eEZw8ElOlsL1pByTsjL84ItfT99WUo3KOy6n3v8yoUBqXFgeBN64
eMo11aGGfzQeQXpOo5YLHnBrdnWsIPYgGxB4t/sfOdD99XMj+lokqFTSWgg+Q57PMJh5dtQE+g6g
I/yp4Rr5ftBYs6EkafRVLsgZLVPFc5LnINB5aL3zGL73jlUqnWHovKjlXv/oJ9ZQYnN5mb7DD9/n
9ApBR0hiPrRI6FfA97XoKfzbAY2yqP6kWtZ+VPnDtsKyA8Mm5dAUf9nCpcaFvU+RcG+icrkrV+6J
a8lIhrFI8nSE7mqlzN5a/CXDRrf+7b1SKQ84slkhZePAhMEjtIO5n7wLD1hoPLIzLou1vNrAx3c0
SCG61nDv3jjcuOe9jWms8yC/VJfDmFmH3ZHK4poqogNc5rR2842DAxX3/Ng/PZquc7haIMZ5oALp
avIXOE6Rl+frood2VRpFWk5h+u38XLTmXMG3t+n8kz3nR6jlbsZDeGvlkhQSH0B+nDTqCmnEu8zu
9EG+zwRIiDL4sTgDBX/RG4A+/wIylU6g+zKcjeBNXntWCf59xZ1GYhQ0ZjgvUHmaBN/T1USCDvCD
nr9Y3vvMKJcOWFbose3VjxiRh4/et8ENhsTUY2acCgI5rJefKbsoa9YsqJnRBVS5WU9qdl+e0ic9
RE3Ma8w4zLEdG/LLaE30pJakyCl+KMIWSX7re/J9IsUtZbZV4WqB2hESVM+Klkquby/UfqUNoiyc
pa7sM0f5Zaweq4G5buVVhoyCy4e/0doqbrGMIQKlcWlCXeYDb+ZZwLbz/iSDAxktslYkzQENae7S
ptdb6BLHKbQApqvjViANEnxQclaMGRZevZt/EbqjROKaf5Ona1pm6s2FwYv4qmDrJpY06wPTWLLT
uGaBAQPD2jVzTYvJnp3u6n1EUAuMRQE9C11t84vwBaZHqcE1DnoehYBmHw2vD3tOzdEdiBeVWV/+
UFnGa+EbGrseGtspnzvlnoseM/yYjHnswThU+dYPv37l9YwGGcJGq02NYDQi7RbtPBINuTdZAl7f
7xCM2RFv282El2Bg5kJJ0Gjxx+cN6OgNkfGOPRapxluVysG/QN4P7cqJ2kBGWudUEEvcLY11I65F
1haHYhtEIC10T15FtuxMhcAsAjnWuhLvDG4CaNLegYWOVn3732lJbeF82sYopNxZSpM7krQmrgMs
wdjH4YJOy9EdH1A7QYixJzHhPDZovj9Joc1YxK+82nXoNoPpigFjtV8uQCtwAG30AbFlKJCVfwpg
zPFXmi9Bsm5F4r8kCkLJwBSzxDH/vUvDb8A3EUa2sDMOSEg/oL9VaX33xyzSGll3ZCNWZjZWCrLx
lpjJjBhSMWIaTijw9cXpueYp9aGd8UdUAJjDYtEdvi21pyuzIbZ8letfVhnWmxIr+y6tULoFWREh
krxPKrL5LCeH4g9dDrluzFnqeovXF8//MXqPD6rtgD2UPpBjFQYJk7tOpPiyioreTEy73k/LbJcy
DZKM8IrS6s6GabxWeY2Si8yvhv/ayf4etvqkINlYE+qeXr1klAHrtG2Z4dc3Ka0p0Aacea7us9J/
gH3OfGtHMxRQv19fYBN+yMhQ22+zJ5UmNQ1ao5XUWCkPoNU5WDtHMaRVVJ9+NhK+0ixd8uIyY5zu
ZCqFq5FkLTrH64dr0ZFx9zdBiwtxVvwb1yZg6UbeFZsXOfSYQxeF0reblMcb+Kht8w/LOJCKBFjO
gkzpa1hlCTmfjqYtDQzPSRNcxyf8TuLBRD6KC0ch6mgGujdIe4RSe8IMNsSHmHS9e3srFOfOvj7N
EcgBTUck5Fo75fk/ufdpIt0rIzDN7zhQsunx3C45etkQP/qCmYML1nxw6j6N5jpym9ZcP3AxOTev
i9L6u+Tqp/djGzoRWAxr4gVCxokmnkJYkuY7UQHmdvAtmaT5Hi5rhcPijxilBocvPCLQ664LiUai
m5ZmiCtzYYBg5YWJ4fNQtfepl/sAaubaNtGsYGn/Wx1hpgolfKfrcxzrZPA8R8JCFBkGmYtcgtlz
TBXsXdhqDiZhB/ciYNBdUakmnEKsINvT6qF7siu7J6jC7ndocxrxsLgDRgAy8e9J2AhVtn6ZlqVa
FpNzVBr0dEnppheZIWTC8/bO8C3nfDQL/z6JsrnbUyobRbbYeBdb9DWAQrPjc3jinJsNv/+13Gy7
jZQR4W6/gyrFlM4lArj1ejJ4MwbX+yh1PoD/YIyfZtJkvbpghIGFj4m3OrVoy5UfdeeNGArZ19ek
jdCORNZfMXDjtaqYJbikDY3+OBI1ENqC+8AGacyzik5rVS+WmJkja9gScKY4xodG0DKC1B2BQ2Ui
8ee99Gr5T5s09aFu8bzT2PlXLWw9Xl8TBKsMp+tsN+dpT6hCpwMPobR9EBtXEHiwxudK5I/ydVh4
1euSCTbxD1YJCRDmnYuj96VixUF8eSyyaewkYbw6c62WYvOJnu0NL9GHiFIgaYEREQvhtv1f5mgm
alQM4gsxIqgZR7kb65h+wbjC0gPRJnSRxDtDw/LnTVs2iB/ulSmq3GD1adRZ6pp7T+nITK1VhrTP
365n8rwWaCaECFunpXqKMSwbEbDaTa1w0anDXdRZpnYmpn8B8hD+DmkyX5rp88zOBlufJPnQK+ym
wdE28uFCLarzd2U73GGCFCfdP3cwbZ9sE4M/0oQFzjHNdIp3a9wFPQLlrrsSnyPYeTyirc6Y0ZLk
9fFmK1VHphRTZzzUat/FqkDcfb79+X2YmongdE3wLpCYUI2k6ChX2mlAbgrWWH4UJt5f2AFvJXF4
nDN2VIi1rXryR9Uh1TlyxLYklvXSX+H9NqqLhR+1vkp2Cf5ICmr6TODUh4EGeO8GzFBS9mY5ZnAG
CCEFUkwBx7pRCmKPxMyVo1f8u/6lv+C29C6OfmW1Tg9k+wNgqxz9/vBKKHQTDwLayT2bueWJa1VG
jT11nM9cJ2s86RonGwMc+CYJ//ca0m+hg5mvZQg4uE1NId9OK1yCg9tp09FILlGebGpy6VGX4up5
TglDVEmH+q12hg9JZwudu28AmGYKa1I8sRKjNpDkRnsQCXWnjxwP0rxUiztlHsgPGUqoPdw01QTD
5x8ra5AGv/CpI1VZDKsnHfey01a8Om/liIxLGG/j0SZQeTPhzna/+vU/hgH5f5hYsSwxcgX06zui
dvgH97Q9TL4eytsXjmQI2D5oX24hwWM7ofjAnFVeXUWmF5N5auViAQRMIuz5b8qj5ViMj0PcKpLe
FssEM36IlaPA4LECzIXBnV04OabfTA6ypez3NENvG3lxdS3JdrD35STnpBm+DkxjJOhFCY9PrJtv
mPnxbggR9BdU4U9boL7isLtk8+VhEiIpBFvihwTb2EcrI70QijyuWhuz4DDxHafC6kKZd8Ok1tgt
Nd96M5i9KCNBnvUZym1swUQnHU1xW2tdfTrh3Lt9yNFJsbtp1VayM3ymP8Mr3azcpUbEJsX94FGX
MEdCdFq4iSaFaooEKCD2D9sv+ZScdMO0/5VYDZlIGt39acI/MC6AvdNjJUaCtJ4UJVOSYOHHnSEr
NgpDvtWzATOa9yX8FCBqxsbESsESa6UpYHv7b/ZV+QPXcNObgPm3tskWnkqSNrkyafgkzJNwQjfe
z01oSftP1x6OhK5zdKVr9iGyWNva45JDOoQUEO04vaolmX4Y76UMr1WbekTJNg3ojkvODrLG/FBX
jxhQvlpVJVVSYY0DCYt2TqMUIKOt+oEaFDX+YogHZCR6gHiDB5a7b56Zjd9e1HY1ASXAZM7M3xlT
uPHw7mOK0+PCpCqQUpAykZOgi1DLxOZOrSQO2taLhRrenD71VgtJV2YntQcip0B/p9nj9f/vaLkJ
v+nczfn2Os3ZkB1/zBPyImq/BW2KBeykD7uezt1eNdCHYsapjjLs5p4PXkBdR8awLpNlITxLhcy1
0+kmI/jiA0bA9R5UoxEUajjxLqd045JsPMBJ5odYLVWdXDqq36iO4m+E93n9q2kQdiflx0GWIgnu
dtYp7pXP1ibwRONxBOy8oxslF47ap+K/tcEAnzMINYqMCdQCVr9qO1hGR0599PveDWY95dcq+T4n
qlKbmsXNozmvajIGdBgw0sgN/TPidMs3S/dSRfosiyTUCmT5wJnpn1kzTKo2gI7gXZDSSQYZUfdc
uC4KY2txHI39GKyyBiBPUrAfSbFOkLE9KZVwK6aS1GfyPIVHZ22GS+Q1gjyR6xuM+Vj9pO6jAWDy
Ed+HgHKtOvOgwrZ8ViqSTDI02XxE3Zf3eKz2Q//MePpn6HVfHeFeKme/P4sCFvz5itKUkolO4QES
9/1bWv3T6II1MAJk1ymei0R4BrkXwUXc8ULmAgtHxeBlCmb9i4EQ7J+4MLQEjcEtzkhWkZDEBZ6g
6OZ2+k9WWmIjN4bpqWvbCRR4AloDU5lZx3LUlj9HP0bIaJNTk0U0nRtNba5HRafBLk4GsLuLzY4M
ajNmSvY3mgRvzo/yx65FoYFugYnEBkXYmf9TGn9UNpqCm/g40mTPZBbeCUb4RaGr073GBnxg944q
Ea8c9N8QVrsla2DCCcXNxit3YnHLJ12MTvsez9WUwAt2K81R86CuRtvt3RN8kElaScg7O7n9Y/xW
ktUPlssvZj8Jj0sxb0BurstQqjwPLrArMTASWUzql2kUcW8RYgAU8Qsakfj9FD+Gq0Po7QB6FqMl
C86viOc03842RQVnX88QVQgmiVwRPuYQ7ahlhZhgbbf6HBRHpBGoh2XgK7p0dIrVmpIW1dih794v
VhL0k+g3U5YjI3yVQmPpY4fL0ApdVFK/HOs+/ZAjbjSxZ/6gilMDQTfhszjLv8+OQHzd3VDQPFWB
jESaaMUER1VV4hHSRXRyj8VUjFLbmbFlIP0PDk7NnS/VsyLWxdQ5N0jSJuysi9Ww4eqycA8e6P5z
FEc8tM2dHnCvQPaF6H9WurLQa2RVrYSW79T0QxwXqFvdxIozuxve9F12cydROTsk+OSQ2rAe+MZT
w2rOYv8Ag9rLu29jJT2TrtvJhIFnHVPiLXRvCcC+zOwzGXxYrrLuGjfhYrpaxz0ujNHJ5q63uWmz
P/YS6uERFAZvejDq1AkUZl3fOBYs0ytDtZ13RubEdBVM3mgJJy+uE3zzB9TkzamRBDxXD9bHqteH
Y1eihjDzzdBw/nk3op6hl/lNozVQQu3A+mArrlE+NApMBWWbJpGYAag0V+lDKifn/+BxSNb3pkX7
QZMGzYydgT1t2GtmD+ScXLE/PB3BgoFkJ6zY61jcT8sMeUBuIF1mp71wgrdfUIiM8K6FErymVOc9
LVj3B1EeBpQWHVAqMxzs5k7UY8q+hBpdTuwFtZukJ2RO/h7EvWf+1ZYGP09wcUXhK/o+4G14QGcY
LMLsHEpnDH4bFJuHGgMDevyFu+/jwJTRjljbr7QCf8FmyGuYPTayv8aISGtjyJVkqEWh/2PgCPNX
myBEr+jY25M0ZWS1ACytumr0cHZ0AD0LVKzxG0KhHbbZBZBBhGBNy91gEe55t7+RIoSClDJHeZzI
HhTKJim56BQKbva7Lm7B0XdbJjZ5wGZ+iU5C9Pgd1AC0dDLQiGcbnRCwkAJ10xcczcPnMsEU7dJM
XDlN9RhRvpP4/QEoBYwxoj40RswesSRzFA26wkSagR1Lic6RcswDf+NNw3hefLB6OEBQGVSgjRjG
+NUHXHjmyqO4PO9aBjqfyrU8GKSQY7x2FrX4NtZddfQx0qH7PmTWJcHjrMPZtfPdRnppdbueBbRX
0405+qV6qSjT7CmaYW8JsBu49ZU9Rb0JQAIXqB+zaKqdXxYQEsEaVfyB+xMJRcgasY+qiKO5U0jg
KvzwkJEDfpP2DpaP3voVYbVeE+vtr7s0dM/HJGpQfuANtl/TfWqhpp8/kg7Gfinf86TzKmknq1qM
z8FFKJjT+n5X+mRYGdIlpBP5KirsKCbGSTH3d9pLD9s7ItCgXiOkKUrg7GCWuVJiZ6MWbUld8D+Y
CIm88pn8dn/edFQ7Xb/bu+Ht5gEt0Vx1Ojc9O4WWgTbe5DB59j/6A1+RLPtnhAm72qwFukeMoZ8+
VTQOwtxtCBK7WGx/jxvCu0tlLRNxFSKD4yDilC25e5p/P5P1Nwjcj7Og9gKr3LnyYU2iN5SDHYGI
/aUs5X5jcacxZzZwHEb7eI0U4eMvMHM9Hl6yZ1THKeejhhqJ33UpyDgsKvJploGJNje892epun4P
CwdABXdg9wQLtiHY8kg+P+AB/4jg2DcajbIfyioaHoGreZ2VWqY2t+bzZGJILlB2L78S2tERtBGV
Iv7+511mmf+2WNJORNoDb0LhmoMFyfPdQi5G9dG237qYui0kMvSvA2evodZXKwaYrIAokknkjRJX
MQl1WwraC65podb41v2XgUP9jPPPGY/MAPxyKH4Kul3O9y85OfBd8uZl9W/karIY75toLRPVz0Js
o5Gp8f1aCM5bw2XGnKxLNIowoRDAwOG+qz/xu+lGztlLD+K7XqlIzzAp6OiWMhfli8oqyuCzYM1T
poWM9THtBUSYe1mnLLqvzCWwldvr9exZCWxy49fVDC4C5oliftAbpjawrF6lX6gzw3gnHD1Nfoxa
U3SJ1JckjugGvIW87C+tAfBgVAi/CukTdtfcHDhuTHauvP611U9N6PL1uCrIrgAKTRQSKvb5Vr41
ezzWjXXgJSGXeUY2v8wAURY7CKlITAOhfno1QDeIjJiDU2B1QZ+jf7GjRnSr8aZz6J6tAIGEqzwH
8EGC50d1Vqz/nxn15Zg+btsMwbNUQESbRx3octYuwMo0LozvQQwbHGnEAE2kIt8BlOVy+cDptTvf
hAEXzxpkgxau/I1p7p5jcu4K+gm/iupScMsC4VKokZXiMxCHjn32uLtolqfU8qwWbbJkbLYGhAcS
zkN1mxYmGT4b4+vyezMtfaN2Lj6LRxXNy7pM/JOw8GSsuF/VARNnPksEtf0JsTQ3Cv6jwYr7wmvN
X5ZhBcEKGO2i8ozbbfWst4Yksh8wHr2PD76my1LxQHw9LK1u67xPlnQawgzPf35mgGjzlHqFTlqM
fAqVaxIvgww+JFWbpIjXYAL+95o202N96KgycPkIS+1Z2yxQBt5Pu4iE7wAzIRnv1csWiHwYCDlk
6I3BPcCEo2CS7/CPslFauvEoLeRzyDQQEwaGBdbBeDjpvQyDqS/yfSS7JFtFTAjJ+vHm3oW4fIA8
H2q1lta/0KZ3fRZFsYjPB8vpiQ31Ij8S3W7iVQbBS1o9FRAK6waq56Aoa6dm61i4eNbAvvsbvnE5
Z+quLK9EiTwJGhBkUnuxHcJbk7Vwigzj2n3shyC+RaNhN4PYYEeg9QA1b0vpQ9ADIC3Hje37/my6
xFVIa1GE0Hlnl0CvWXYEKvuKJFlwwJfex/vcWFLBwoCRfLHrWVTqptnJ3QDahKzRBRwY7NMLBDiu
Rg43f2bORLyP7W1+nhar6EH1oMdJJNXPI9DjaEsJTx5f2TY6ZhXFhzqYrxI4Y3VoTEFfIEIZU6yj
z9EBII49TYGsPXlJWO0riIVcAPPmcwMVWaR41sEFB7tw6vQ3FNZ7B1ugECyKoXaRc3U2i8eKKGOI
g5A/kupBmL5lCVh0ZNjfBxg08FMlfG3swT+aVf7zczfHdpQ56QfXjjhcjX0JePG+kCWc+Q6O9ZIq
UQN2UoCQi8yf3lvhr0hvlqj5AgLIu5ZSS55v8Ie0uPI1FP40thrB3faMY1AtYn1DsDNhgEQGjmj9
XklFvywajypK5eI9V8HN4MqfLZPcLn9/LSDbdAButeZT/QFd97PlN92PSC/6p4o6tM9krW5ulWGt
NZYBEVZc3b8e7aWWL5czBHACkV7kDCPx/zbC51AFo/RjCTCt2flZgz6VBMmRh/lZqIgUpaHPtI7v
l2ycoZK/lYmNQHL9A6+6LXaGL8MDwvH/9+zP9W6C9Jo2c/fdo4Ckj8UCvNmIiGOtxyZkJ35dne57
hHyMq3WPi5kSWLlezEDVZ5qSOZ/4X8NA9V8x9EHAlx1qIhvPlvNkyxo6he+eIAETzrXF8vrwBWkP
9rAUxuJw4qba4jmYCw5Ije37pTQ15+Em/wfyhPwPB5fo3XGuiijUvMOQ7kpNybQb19O1jS9kdzqq
dxrrUE5QTCOkGU34qh+cHufQYt4H+Fuo9Bc/LUnCB/rmuwuYvXNu0RzC82qPk/Dees2MOtcoepLj
aIxk4yP9NiwhcwN2cvVXtoj4jmV7bJnNrynfXQquubuQdRgm78GalTox+Rg4uzJUPCkC3u6BmEAN
041QjoetnRM9pgw8Ein1xH24nOUK6q8EuPgVXHoDUMVxnbKS4tHpdv4TgEr02xI6eEGrZ1f1kNOe
9yA90PP2+wbqQ+sV70Yg17NH25uUVNMebLTuQsxjQRQ16l+sGN2mTXLo1bujZuf+UPVRGIel6NwB
dounKBf2m7TmR9SqqEEK53AlrM1Lx/GicGEzhs5inoY7Pt2ph9TcdS6cBmMdxLkObdqaSr4Selcr
NrXuqHTD24IAMTZASX+Sd8m9dn2fgfSOVzGz1MtFcywv8ELAJFTiJa87YjhozwfjouO5HmvOqQ9y
zUGs0aIpsm/pus7TL0j1MQkBzGtcqGi26PAuGVLNzr/P0ZrVIxHwvaP2uFxS2OLWXDi/RWgvGWt6
Vcz3TZdtBOW7w23/Z4LKCoqEZLJOeHHe/DXtoZFawazzNzxHq1FbtfsM0zsFCUCsOTXnRESCJjNy
i/NTKQmJ1Ir8yw43qvFLcjHPcYwLJk2binf7rCHOs906s+s3s0qp2zDdzMuu/nSNVL1rwu2JSox9
gQO6ijQ0GrnZ2vpZQYjjU3evM/ouLYZbBg3525lKgihYXNQwDk+xV8Ok4TVgg2AzBGftVPpGOdOS
+yvNtTL/1MhGrVuQkl1p88QMQGvXukL01obYjPbFofzzVG1LEao7Re53D+mGgJjXx6sE0VcLjIXw
/El9xg+K/0ZD3pC1Wwm0V1I0Ry6U6N+DXO5KIdVexDwuXC2f0Z1cozIBbDqwkfb0t2SMSGjonGCx
UdjrpM1qEN+NQtvndRAr7D2RdTOPDnsxZSy6x2WmcmLxovO6S5uIxGqJXPchRCXkSgyHH3SSzcGr
RcBlX65tl8Y7jVO8Fhmwpf7WQJHLEBC9JaS4DpWo1MC+sOW00C4SbumKQSImyV4r/Boe5T2z6zpX
9HEeU5KjBQTkkxYZUeMXvoHkJDPSmK0gqEbDQV0YekaZ1NrWyMFSF23PMxzdVbxk91M+Dc7QBQTk
xgDS9OAk+fKL5aNSTkJyCKJgz2KDsvlU34u4izbs0hy3MKEqvYJLWNE4mfDAYiXZAfYwlPvFzTqn
0Qpgr14oKmo8QZj7O2kAnwH9mZ06q+4QEcOlAEXZsudKn1lMgy7iiCVdKJR6DNbXo26cqXUoOmKT
XEs8L/fGWPwP4Wwuxl74Q4nosQJwmG+2MFKvwx6qtqnweOfM0Rcz5t1DW4BO2m7YfuiOpugxOfvK
bhyPm6LjDjVnsfDE+f+PwKkK5D4mbFocSDC1g1lZpxUEqaKOisoRo7/VCYGtLjpZisWRZDCjK+lA
OuC6L3c5i3yy9K2obGxrQ8eUsB7mh5J0E8qdD/LsSUzTy2mgBjmqIDkngjPDch/y0a0MA2O/VS1m
iIu+bhb81LGmMzqPkjwP6rcbZXa4BWK9/Xcfiam7mosU+vP9iKs5sxCC/IMj0OHVdzNINfQ5Yata
EB+qMIlr/+EC5eCL5mXn+O+G5/gzdBAqB8u6k5P0KDfANaTEYvHgS4X4V3a131I6Uafy75C7emFK
hyPZdHxgpPEF32/2qgkqTz/S8uMe6rwXdigyngkxSpk1J8TnXgPf3oYMkqyXvD0oRNED079euR0O
QvypOErq1I6ZCVXL7TijWf4CtYGhCans/D3DgTtLoi5V+GOTTi4X2JU5uTlWruufEGFSP5PRYFir
5SkEfP1vATTZrLBzYAEr2qbabTqMTLrAN5W29kWnAM9DKrKXrn/b/wz7b+VYcLMiZMl4OLK/Y2Uz
vI96S/5wQ0Qo+TOawHz/f1CfPmDgQR2FQKb8PM5prjVp9yrstBbyB9r+DDCxoSmUwi2EkJjaKqqo
2FJFuXvPlWwu0uEqu8xp6DYPSVfpV6XplCP5qrQ9bbqoy0OOz1ppuWCdHXzHUF2ISgtPam2iwQCU
NSeFeef98mJXR1A9wix5fmovHZXIv15m5tDuH/M9txFKDYOHP7T4/2v+R63Lq6bIOY9Kob93Dkvr
nBqFYN4UShHVgGHezEtVC55YFGU6+8zcjBqc0F6HKThEI6GvaXIcHzZB8ZXkCzwHO/RY3IIfSuKC
qi0g2zKioMV2Tx6igMVx6N3xXxL/s/aJkszEym4iOQNr6d7tH48qGUjttvVN3RPGaXUxCfrcvr9F
IMRtcmMwe3uEFrdF74/bklYrMJKUD3zhbIcXjI8msz9TxM1XHtMLeGYB3Cccrggs/2cf0tnp7Ddm
Qprq03412DXUY2MI98c2faCvWYn6RxkGtg2JlsgDc/C0yAiEvLq0mQKIdg3sDuhoxY27ne2jKEG8
udB8N07jQGEvrF54HGGuFSCxnXi5/ZjtDUjdbfofUTPVEvqT603ua3LcS/bmz7AvfLBOKmRkVXRl
9u+9MYJw4/I0+qgD9SjY8gdVQ6X6FcNlcDyNkUVWWTgqCuCsXODy9q31d5IQN7+KsVP6mHzGOMqW
KglMzmbJMqPyj/Ue9QvWjFRIeDer/8l6n7hBFpNCcCFaULc50g/lZNFRxtHA8e/8GKsKSmF/voOP
Ksz1uXJv9B4Uw8+9PYIuEmsQvaAo1n6m+lAxl8EgNyNxDFgnNuG/cbF1pqnX0p63SWMQXUg/wsq9
d4HoRUCSatMWd4mxHg5bpkQzv7SCuP5u864xnSLE1oLVSXPCUUeA8cUdVp6fOutBDlORgmC8gjAM
hv0nfb3XtawOx5p1CkXfcDc0/Y9jWDYGKCG3K97qUw5aeQJxRmAVCderNTj8nwksK8I/6GjM+pkx
PR3jM3B7/PBjX3Vx/gsXUPA2DrDimzhjW5erlfI0lUaz42guEAtdOCQg2EeJkwS5BPDsG8wdP6pQ
C3GQTd1EBW7UI85j+2PvHQF30o36EKmvCXgbbrnJj1+qoyQB5d1uOg5z5yurCslVOotPKw6DT6cU
R1FCDKCTST4IlZVfqaM+l+AVbpLWLwCJD6nQHTqxgIJcy567VMn6U1jRKEu9Yv8Lmlfb90aGQROU
BNrJjyDrs09TcsI1W+vFSaCHKM7yXqfz9uBppBeYKGKT7uXpLmQLxnozO2Gy8Mmkp3z3s7ZUpM97
WaZsHFkQGgphE1Zabls9tx1fNBAIIFn1h9Dfy5EJA5Jb1FZwIO1dZeshPhLyh2EQR0ZE8oZstlo/
mlTDnC322vQif+KRmDv+ir6Yw8SaXrIuTtrNX4NWR+IHimbhCKL7Jp9/CZUOx/wv/yzxnwrwrFNC
7vCFCBTcgnSv6y/xfT6+D2wWoq3Q5XaBZsNE2rlE91S8AB/zQzUAlUiry1kAtdeLIVVlvtmVcQBe
S5P8mtAf5/F1n/uE6T0A5zncfA5xFeEixmUroO5A/KPI3mtgI0H0m1QYQKye71M3frwSTl2541hH
6T+aUkV1t8QHEKqW/mxbTlGP6QXzJEYVtMxk4XWEqa2Zl5CuVz8Zudpy0iroDddzRfhl4vs3SIt3
J217bEBBTDBHb4YcZb+N72lR39PJbU7sNIoRcIGmc2B0Xj3vECgJ0xcjr3KMo0jdIy6uGhag6WBm
+7UmPnYzEzavqWQTxZwVDEXzgEdsts8WRiJjVGP18UJka03qD3VQIu3yki8yyKzbddOwKy3kl0l6
/+Ms4HR5vE2TwrEQRN22fAtzNhrrNf7FdjAaoa6bLuUKEGoMd88oJK/Syf3pOFKqwb/2J74BY/8g
Mi6NLEjePDG+TijNHem2X38YmzhxRc0jsynAKGfrPrIakVAfo5tKSksZPKYsgqZUeMszONlNmXQF
nthgIxfQt2F4FgvjJUUKxC2qI6ujgWdRqsw/3PFYyQlLgCAyDNWoetPqAUgwEzVEqA8IJa1aT9FB
DzQmJ6eBr/n+JS8Xouy3k8p1imo5w04yVk9Dg5ZXzH0Do7qKOIhugU6v14ps2hVSDHGoQN1NUlex
qdT+6Rxz3gxS60XxnfcmVUC75I7SarxlTdnvNhG/EqC3pT8O7ZDzs6+pA9F1QT17zwiv9na4CKCi
DOJp+pAKD26IILohynqaW2iJSgxSVDkwSsqcah+THdKeFI9/qaKVsfTlF8N+NfoEEA/kkdKo3smB
D8uiUnQGoUuoqFbC2q19Dh8DusxCm1/hZSkdm3K8PH3IK7f2FxC6NnZpCk6PQHrRXN4daSi7IAT4
PrV2Vx/f63PvCFp2HGZx3kq6ToDsvQHlIAJzLcvsMM/IQkMkcs3R75XCfePHEwDoGvHFkxucuier
8KyRXYhO8kYCwwWTVB07LHX1BZBlh2p0R+JHj4igKh0qBdfDhw1j/tzNPb6yPvoKzAIW0I2L+RoU
IypQyFpDfF/JLHdZFkcsFCwhk5Wg3kVKx+v5933MMFueKqrp1nDQFjQB1ZKpgB/a/wM/8ECUrZ9A
z7DUnN+4c/BfzvRcN7J3cgRGWMmYclqNEXH6dYTT5xuHNDS3CwYZwwmbChALSG5ZOn5sCAMAXFMw
f8/WG6mhGQ+oaEQ1zkyvhH2e/VmGYA6NDVv9WznfwtPwl1GLC08XR8KzgHG2zVS2PatFv5fbbJ9x
acgzYS0J1C+pKQfh1+M3wCHvA+tKyyGh8Krscg1QUTeaWWFUHET8EAZuxgeV5Dsdsy9YXJA1PLI7
Bw2kYgQaim0HMlgL2kOsBtIt/xh6ND14VZwwoPxxw7dz1J1CfQHlwrGcDRudr1iCxxG1QdCKPaU0
tRiPkzleVeVYXtmfttEeUgwboBpBNn7Outlocrqm8qv3tymiej0eIp5/AnBR9HCJLQlBSwClpXhj
hW1mvNQGxW880gVBG54BG3oeVphWTKaGre8rVY5Cqh8G2D2KceOdnuTjwQjnCtLfkoynHFukgEbX
7kVa8ILmeuVlEIwfrdaM9YI5PSyqigfh8yza7h8NOK7zt0XFw0qypVl4s6YOlgtMTlkWmdnA46P8
a0E+XUUYG9YnVEXCRGHH3Bpq0gQhgCitmvBQQmED3sFE9idDf7d4dajM2xgayYVeC2BsFT4jIs5P
69po/mPv+1l3DzzUZVHQ+MH6VsU5h8VIfSJJuDWFXSZHIbw0vQsRUCKZNaXkVWfayvSWbCaCVCC0
z6P21aKMySIqo18gGwEWxnmhuUX4clWg1sITffd4MNiiDKUEyLLX3A1GCHRDu1AB84wqW1gx304G
M00XkOBIal01XfBQgnrWpo5NXhMUf86dSheJ063hbZHS8t/U+GGKyc5PMRG8EQLNTFFe1iA/fV8u
Lh75AxZ+S07OMIiPRsey9kSzBoLicsbuDCIAciOZgfDuXD5BWqOIV0+0Q+yEjWVk5m6HRDMZtZo9
uU2is9DoRvEOI7q2VOKFqxrIA0PqlQhbGJUy9KqNpbtRP7AyGOU5NG+3oNfC23KPJy78JnR6y5NK
/akrhtojnP0zi3hbqpKYzKBdR2vmkaDjpUpEiuC0TqfbNiJ8EvFFM5/5dWaho9qIasx78JEDlrFc
2UHZjAHlDi5seKttBcNzzeqzNSNz0XCRU0k5iVkdSf4jS0Vlu39/sqM59mE24dBKW0KgPrj6uFu2
FqG38q+ZD5V6/y7ZqrMnXu9yg2PCV6HErZi2CpADlXOe5hH+niR5p173gZ5G9rTlZi7Lmh+XP8YU
O79ZczdkkXSBop2yCkikbhmD3yCGO72mShMrKlEochTdbANRecozIhlpvFFJgkxlevSKO22Gq/Vf
wEr8eiBG6STVA3/bi8LLYT6Nk3saHlExSmwrCIRhUdEpqd/qxTy3KlNxugEL4IbMmJmEbAs6AFmq
TGmC9jNej/KgjSDiV5jfyZO3I6xwnNVSfI40G1+c6/tnAzhcQaa/a9i0y3as2ELFbT7YHMxFnPMN
jaOVHFZWsqzQPadXkYU5qy5rLX67Ll/u/EFeTJ9uKZVsah7xIiSsvDbX3TG8V/G4Cx+42sqLxWE+
pmsdWHUMRo7XdvKuVfcb+4XBbA7Btj/9mL6GKh2OrSMJLtUbjqqL72lokRtGg4mB5J/aHqovssRW
8LR0oJ1JBc/RUXLSEECZf+euF+imrjbjDOW2zOPnXJo9GjSGb35el8dS+/OwR4Bs6C4PXbKYM3ZX
CzK3tKcbqW5DmhGDmeIVbjj18Z5lpetXt72ybtfC8rPartvtbqKU4JjmqV6FCxVgpujA4eUUwT0G
pFID0dZpO+NTG68SAXlbj6E19uQgcd6vhAuqA7VQA4t7h16Qydd8F27lNOKvzkgzeVyRYSY1SwKc
T7wzC1l8vBd3vE5RznxKazBK2pB00Z53Ng8YDpRyEEFIXFEX+FhtC2QM9VNx8xegDVE/fayZs/jR
iVcxna77wo3PQMYtxFRbFF8I4m5EDkYJeA9+Sg6jmpgHgnZQr5wGE798OyCWEPpG8sAieWsFVbVo
80NqnlztKtiGvqIuYVU0PvPw07y84sjgReYrmJ9Gbcf21BHwAYbpMlxYiCgHIk7sAisW4hDY1igO
A4lg9XWLznx5o1WzLtpMk7KVaIDW6nyaWO6BYaPuEin2mo2uPVxR3XA8dWMU+wWq4Ksq6s13rb3z
8ICtmNupNM52f/NOyh9j3p/fLlgsqrgsT/OgiRx+l6RaUDXKiR5WNgq5hFHE8TZ+SWZXezgs9s7i
gj7kOwMbCuAAwp32ZRNOHaDP573JdHvT4vBzhTPR+/8WNS5NuYURXDtq9EVCVrnrGw21vh8FhMzf
XYvSP1LUpkdMq11UJ4akYU9Zat9zSdnqvDWgLAfXEkIJgTNkSO9eoT1VyL5ecFLk5+xAwm0JOl11
O4f1fBX1QM/3hAOO7QhaeE0CfOwcgWyqc13TPouBoeFrxO5pyvSsC1YOcfe+5IB8Pm8fdz/WJt1z
yUrUxAvm43Kdurem/Spjll3Whzfkek0JGPsK9BNBkugrj0hxgE7RmbDbiXBFrhrk0uqRU54n8y6A
khHX0Uv/FNkOGnoW2HLUw6gqdUhUfA/WHKxtO7OoezlSxMnKch8PSbhAeyS3py4v8dRoc7EapI7X
CowsHImCUb6B/UO3h/af+RBjjRutnkxj8mYia91RGDiWgkMCzQ3X+gpxZsE27dg+Aq6TAFVnY/nh
ouLwxuIfIxan/uU2C1mfVTvq3Okc9dm5LCCMEk/pUtEsiOL0KDN08otVsfIJFidPYP9/nMV6V46N
Vqw/NQLOVaYXiABUlL6qfpgPyQ1Dgn3iJXW3p/5tmBXNpGq4pCVD51dLzC8eURTuxWduA1gqqdCL
i8z36UgQ3CZ/4QDspRNY4fZZTUi9HMoibVlIznOOe3nZ/R8VypHU0Ap+7eTNjbXyWW7rk4eIIANQ
Sv0stnj0XQKsFowL1wiAVGajYyPcum/eLhGwIDxQBRb5yWiyGSQ2RwnIBwqOnI/5uCtzsI3EvvpI
Mgk84elD4yINvrGdNptle/LrjixPVr3ZveUM7RsjlDTbTs4oTzLTXFns/Gep9NPCZgEKwSJCYnbh
k1nXJx2phITxLkb0yvHhC2o43LGWSpco4889o2+Vp+jK/UgcUqXougVJdSgPQwsBTPFbBns12xDy
+RGDMxw6RwBpA8rrC99UF8QqXhdR+bjDGuDuDHqZG5G8hmBtiTXN55eEEOa4PICKaaIdKLW5O029
15htFPEtIM2sBso0AvnznE38K2VU/1nMxHrQQ2A67Vm5T2bcqmeZAmeNO54XDFczXlUeTrISakHp
whWQXtkF2uNudJw1uE/focLwpy8ioLyceqVd2DO1KaZOBEMr16E8SNjdgYjwD220xi4KDD3oFiwb
kjqdl/zrZNpm6nsFAwgB6KNsd/Yh2Me8q19nbaG05eyfG+sXneTjq7lJNzqAoynGz79CaDOHGN7K
y0HmMlmKOZXRt9Jfb3CT+uch7zh4ZUU1tZWgPm9xadQdrFw6BUs1d4uA5Qn9iVIkgPrbNItbdj8C
NAtCUqQsdjSkL4G2l4NDNTbE/IjbTZmpmcWdWslFzfLMNRGlyzuc7kxj6ElnAP/MP/k6PleHG/AR
jMQzQyTDHx9VqyYaYnJApgOOkvk8TeHAh0z0Cc3IgefIyWKCWsOi3HfsKWEbp2QmoF7WZRUY5mTk
f8lgh68VkUZHCP6T/CPzJ8BoVHVZGSY7uLtBwDMqpWFSzEEXj6O/W8jJqAudxzwn27P9Y3yqvkVb
U4nf79iCAimX14NPPpu3l44/cnaczbf/cBgMdkMGErPnoutz992MKz4b4VgR7BUHpMzBtd1vFjRE
6lrwCEA4mACm21OO1y1JMFiX3g8hu3nFRuaqUMZo9qj2H6KCSnYkPjKemuQDPe3vNSnZW9CRYp03
XSj3WqIh3bRK0COKVXjz0UlHc0xBiyC8ZEBpv0dMCUAlkUZcWihWmS+zC5JdjbGOxLcTlchi9st9
KO4Y5YrYvhPYhmSXk7RjZI1An/lfOzpm+y1akpiMa3hE+GjonZ5CwU2BL0Dmk8Kqa0c6HG/toGrQ
ef28z5Zx8SHP5Fl5IHunKnLG5PkLPNnvcp5eGCVKtMc/X38ThIn8aTAjcrJu92T5Fo1TEo5RjUVu
+UAWL9RvPNht6+SwO5WmEfWk/VwkG9vQtVyj5i/BXCxZM1CX0Law2N8BqNxN5U763G/PpVL+cDBu
RDlUupXU2BwbmLs69W5llZPue1XQRrBPx3q13xchGi4+YYitYXxv4Wsi3PoQPf2EeMawFlwjIAeU
DWBmLn0qKiBm3RrkUmK3XFimHXmuGs/S3rqMNxGxdFMBkDQe/okpiWhHPH9HxTy7ONRwyGa5GiwG
KrJTxh+RkkYhYYC4XyhBr3a0qSanYP+2j8JvTpcGTjuoETzVUg7nIjeTj+PR8v6tydBLrE3Jr7Ta
5JsOwPkQeIzDyJIWDwmY3xBKsP4AGbhguLoG0O0S06XkV5rvtgK3DTbvGWQHyA3Nau9Fco4j1Wjd
avCXxFbsr5sD8FPmklGH/UHa9VuFQvKyqGV3+DknjvKSaeiaFfeaI+wqqU60M3HiqOhCkeogkDsN
oiGTShkGNMfFvMp2BU1wEyGY5KUbymg2q+0XfKClofvCS+hfjDlXBPhs0aRmsL95pmdBEqwjZ2uM
dSUR6DctED3LZLgS6v3sH0Aq9+Bd0pU2w5uQncdhDdt8QKmKV6GYe/jEkojCXvTQViP31PTKHuyX
xQtgB0l4uI/6RxnKJCB49cm6h+6bGBqucefM4UpKUwsJwHl/nL8Sc39OPSxXBO/MSPSJpHh3GWpt
1v9af6fewjg2FZpq6w6N9T7K/EAHk7H1kbMuNj962YgJzCzY0hlvB/ZkT9iUHF6Kho7vzc5y0P15
rXoMFRgexVT81vdGlpHY+CbhBaG87+IKyHBt+GLFaGWZrLX9mRbBdPJHeEJmAxe8wM31zBklcM67
o8tLPVqTaXPzFa9HB4xfyAO+QkCAgOjqWRaF2LdzBg58VzvyYa/zOtwXpAbp8yFVxBj1lHnDSZgc
gIe8pQSnITKbyAS++cAg2ptrcjc2JBoWHNhpllXSAjwhUhcgHwxgBBW7rCwkOfqz/q6cozzjBdsl
9Bg3EmBwe/92XoDqRpIjmbM8SWPUubIVGf5lRU2JkpEJsIYjdciU4HS7TL5h0BOs8zl54FD0kuQV
j3+0bqnOfA57CiSNSenhdAlp2uuM/dGQd8HoM0tRisPDZabQsUXSDrsNlgz6Jj+MuAlSNTgtztA8
bjfLsPX1vB4k+osXfevOJ1Nh0hULQl9udadEKXmxaAwEmqR6cvZYbo1O0fhMbFebyPanCHMe2U9D
XvcMOuXxEzqXCLIxmJOE4wsxUXi+43BuZI2NdOHvXjyZ/lbzxjcPWxfB6/GFWTOADcVda57xNIuM
+pUVOMTRKUpCEYbP2zNaYGvqx18W1JkoZBaH8Gq0nq+CbXQvJgP4XRimWH0YAZI15vDNvKNjAa7n
nzZ9BLGGgIFvtQf3YKoYCphbauxbwOl/GtCvCQP68AjgEV5tEuDZN62KFE7FNglOYEPT69U8LtZB
OPrYOCieXny17UQbSZvd25ZjtmQjvvidziC0UoXzThHetD2a2Tq2xNNsB7UC9v3oSYQQ5V8cxMu2
x6s4UL9YPIFGX8SYnLVW0sQyxxYIKHamVkDHKqJiqB3f7A9B5vfn0hICrPTesF2ODNJKx/feaHsp
Qm1oUxhMl6YSqCwTawaQuYSE+JSIdmg7l32BuZhrLCFARIgLEFAgY6dpDkIGcbDMv5UPP4SZIzX8
XY3Xpzk3yhR6yIaEJnMJoAomxN+uLZF0OPczfVFr188lnCVGCz+fEOfj45JpyOIT2xToJqhp8YeJ
KrrBn3HZufAa68HRg92IXZRtzhsJYt4wfuVoRKw8WcLBtrE9y4UtH3vpHxxiafHzkoeOE4hW6s/4
odnOnwl1B02SYG3StStEr38cuqnm2E9RqyAw1mjkMGLDaK0TNupdN6qnrDODxxK1bjMMZL4DyFq6
6dNlxg0kED6sgT6sFVfymPZV5enzMlROXCv2w7dNXCFHRGiXMzSRz7lAsvsmTulnwV6D06TvWGv6
Zilf7jN9pOivHn24GmTFNIv9/34n76NR3xcOEDASIkCFC6qZx06QLWGSOdtZVa7He11wRtgFN222
N+GKZu4qe3EUQUqvHVsL66wCCb/PwHqDcYsXnL6WKMlGo3qKJ4upzKYwRjRDXF4Ayv8i9jDDPkCO
9uiVPHICD4NG+bWhBpEPe/CibyG9/XhXkWp9g108uTVXRLriiVKZYiHzscP9y6O4xAOeZJ5Ktagl
lnKfu4SQNTwyetGdJDrpDHH9mIUzfG3K/Pqdhik8TGLg8LC6ci96YFjHvj139KViazYQqdCu82QT
DVyFv7AUEEYR74+uSgbVn6btPNdKs6tKBqiaVJ71c2mtd0PgOrx9seKDjFHb4SSlPNAGPGzIdpSe
puypLAX4XYkjt/yrFj+oW0aAICD1oNd8snLXUmMOB9GDvZkpCcuOHyQ6x72qv2nLtbKtDiYQAPuk
F13RDfjTNqlnvWVoZwnef5NaVWW2/IWVUoQAZG0cnOVaRH840g163UHnILDOTse/JRepgGMFiGft
ZHBQ2+JuKuDlGQCVmj5PzPI+RRhvTx0bPPPIL/sbao1d4mQEOqXmMJpnV26psF5ltglBw0C31ixb
Eo3Plsls2uUzUlsdcXmSRWPJpUdV+Pe7sUhUvsRWMoeGg0euPAGliZALB42v+ZsrEEYviX8XKcUT
091AAUs1l3+5oBWIVo0r/YQmrcDUw7ao/bbP3CmovJLZ0bWs3ZerinzXA4q1cffnft4DQXU8hNg3
7/7S7seDSUnfrykB/9A9+MbF3nFgWo06eaFyH2AxuSkZx+GdjGv/dHx3pu5ZHeLz+JNlhfesIGXx
lsqTKwRTcA6Xplr1gc4R588WYN3mPbmxsOygwmSfqKnME7OEDAWDYrgOH3Ou5XjrOe2XTY+zSt0V
rz7yN+qXoebHSU8eLUpP3JxLKBFq+a+18lQCg3PfKUWy/cGwPbWKYCInj1IAvPUgbshrUvyZ6i3w
XQr6dKK46dAl4p+cEkZeZr4TbaTiagtloQVneuxfe/qXYK69DFleMYorEyrzgyF8sKg8kbYZuhuF
bkoWmyFzT2PX6uoSk7u6C9fGaH0fUaq7+Xhldf/LG6sWweIwqHOdY+CWesV0cvRfjcMD/4EeCnIE
3QFj8y4DOoBT/85xWzoehq42GU8bps3FL7nMTlgwJsPDvqG9RZxXifZ+5dc90NNeEkmcyqMRd+aN
pwMom1WHWrgZ0oUr0npQcaxQJALW8oYTa+E0DhU12xTIsCXYvlmBQRD5VWppJ3XAmDQftZWudP1f
3BEQjBSBEzBwSzoBqMZ9UCCjUbRN2StkhhujyEnQL9ZdAw+C+T+8mPp30xCU93hW1zcXMBxuZo++
AAl2it9bnqdvXtSQ0zLn5FIflqoinnczSuljc6jwepeopvZuK+vgsKzUak0SdqUQ39gKh9ZSiZyU
fB09dLuttNPElvOd9T7CI/P7+2Ian3eDr5dUwLXxJGd01KURWHem6dzEU984s4BAXzoNKvla1Cf7
msHlheEIkBNHfQ5uApx0eVTKJiTRLH15cVnlnU+c6LrBG72itVerGJ+Hff7iGgR188vZ4IHhJKY2
ZgmI3gn9MPgQLJ6Eor/5FH2G+folOKDdwOEpe9vypNXvZoASXpz23DPiSFXaELYn9UX8EamQaaVY
7lrcUX06YNUVl1UuupsONG4iyFA7m7eoKVyOsMM5OPobVU0AGAet+YBJd2WWl9Ke9YpfiMA+0oYr
HwGswKVestAb/TcuT36DXdnBw/nlTCXOhD4DI95KlS9b2CfQfKMs97/jwaK572BjEHE0BXahgCEh
Gak93llhDpVoBLlx70hbL7l+upH/O8tFg7Vy6qtK9CgBewuoap3vJy3t/XndtlpGSVn7YFRuwT/p
jX/1tyGTl1sAti9QTXWE4l0zFaCu13KNsTVHEDvaX+Z+Bnt1CMvRW5w79zorNq935dnd29G4jCtR
ai+I1QX4f4HFcX5ErM1ZITN74C8a4lEbWF7EYhApiABYzT0qrY4BGOy217VzoNWAWVfblJyaiCrS
ZpzHx7t85UhmnxMVST4vwNadmz75NaWykc38ff4Bj/dUmNU8VCSzISsS4skL8hj/ZdAR3n3BerdZ
j7a/3rIJbWdnLK9yjNT+lD4R2UY/9cAuxXb+B8ETDoF1aTgiuTQ2iyuCm6/4euOQ5JVPNtZlowsH
sEbwdjZuR/mEddF9iVtuUdr2DSj66tl0AbbkIvh0aMSdtGQzmSA7wtwRBvi0ail/dyHgUdD7djdq
Z5lJKxB5zbnCemy2zxYjvvFwJzKdhtc0pa8aJyhKq+koOpHCJHcRJspHB9BYXvOrQPKMW6TUIr6K
C2K7RrPxNM+yNQNtCZ36CKzCcucjcorBiikCilBCU7phzZZy5d3qU6E75d0FCcpiHYFN/g2QkbqP
lvBttcVmzSuf75cpTyyNOs7C1Hho8TPHZojJyrKb0eqKWhXTVALXsvM2TyadceZViET7IzumBki8
7DUKivtMJ9qklHI3xLZ4ExlFIRPfwADzaiSzRu0bGRSvRXlc7Wfy+LaQOhATzvuiAKQn+Wm59hr3
elq5gn7NAWD+Ry8DYU7iKYNbNb4axArOQhfZ/f2gFglustANyeUE9HCAbPNILL0AK9BlLsZH5QwY
1ODPF8Ooha8/if4Po/rxveNV9f9eEXVgHR2s2U4kctrJ7gWdailuXOlQ3lE9Lz6QRi07lUK8DuwE
8XIy0y8j6GRm6LD8Foem/L4i4oCa9JBqTQtQCAd5W2dtONSnhIh7RpksxgHUmysKn0MyPaRoGGuz
nHFin24VFGqetllpFPozudE5k0Sd9kdSzhvpX2dWeH6jiCrqmm8hy2l9W51Er1ULatgkiO1d6y5s
8cXc1EEIcmhYqPknzxRKYcjgU5Wg5carE06IVJyTpMOsl2dZkGYZREIV/ynSF7JPO45sp0NvvKif
r4D58B8QWw3XEUEZnEyzlO1MhKbB3BLQLWtU3p26KYnZJld3DXNjaFChKPMwpSc5iZB/3FaKbjJn
kWyTH+1zra1XqdZggP+Nt28Rp9y31+XzQqNMlpO2/OSmJ3QgUmOmf35hMA5EIi/NF4x/4K5W0EHD
LgaECZnFzuZfKZz55k45FPZT+vcA4WLezTzasNTIiOag0bgIw/AfON71IrPmlgO7rliADGNvVG9i
V8owJlV+Gn6r2EgqIgmSO5mT/uzlFFZGFnTtw1+htjBWyAt0y5+CX+5TEu1cDFj8ryQjPDHYd4Re
nepfnI81XldUE8sfieGbTxcayNzKZKoIIQuzfIQNzyUqLCL05+snMShmgu+hHNV3Uy+21ZTOc8yz
GR2ZtNEgmvA4pH2/cCk6KTExkrldTCxjR+DU/t7YnhCirkx4g+Hz17XCXcLufZU1AJMnHERabVBa
rOnCLwvp8eMck3X1apVFiOllKP4WQUW54JJPLFH69kR/k6FZOBvjAflsArpPulW7dnYFn4Kti4kO
ONb6czjTXq6r+jBNG/ZUBTaoJkbR8gHl6mKLyNjP+4ZL0NjmidptFQEzuShfD43ETyGDaesqB6U6
K4VB0N22+Y5C1501EsQQqyE97QKSVoA0tuC3eaUxKSWHFxHN6S8eJE+o8qE0jSuFMJHGypjyxR6r
opRKIYGm9tZpanYVwvOdRRPTOSO9Q3avGEBngXW3Ta7Ts0UKjoNWAetT3GE648MWq2sOrLHYbim/
m1gzal50rxx6z2FF3lVeefNPTWIylnRdVuFEzcQ6X2zVMZgsWBAIkuAZiYWznGAZSuZ0yIVvp0gt
16GXKsuSDQNchPxz4X9pCvvBhNyjjDG7eOz3CG4ZUkTNA6mRPkwKKkwS8xyffdzn9fAWpa/I58l+
Wpdmf7G3iStbEnvtfyjLQ5ezvyspt9+hEZffA7AglCsQT9rdj+43Gx8hNg1Qp3VXwMl1vhnBlbf6
WmPgODJcuC9dlwzybtwHHnGCZZGDsso+oVvqm6TM8YRgxcLKyd2xWsMI0uzDyraTvgCCzPO2BHv2
iywN7uDVOI2ADdMeDgE2k4bkU0kdQJoyiiJVJ6F5O4h8iYHnujCzP4OnQjp6QJun6AXS8RbToNqV
1Jw6kGwzk/985RAKOjEQ5ql/yPRYi0xwBecafFsgqBR9h2M9sLwvv7ceAv/bH1IVK0v38Jem9/jW
Kj/4uk3yNCHoAkML4QzKZOH4qthnuBZpN7B3diPVjGUY+dL9HWh37P4hnarHN0a5GocQDbZnwYqv
LS/Sey58uU+HLh6Ht8ZDJUCYJF2y+MHNZAn3X1+wpjXYP/ahgAX4+DgYfjgHNLB0AveAY+kh4OCX
e/JN13cXBjAC0F/kbaZqQcIteYdpDE1OOCPRh3ZPQ6X+NjopqDqgyJ2WGn5EDAWB2fvJm2W+bmUw
046gAdN7y08g3O7DP4gGk65iAkFsvAjuWxOR2k3YOkMniK6Ius0EYiFn+n26SgvSdUOB7YFwMFjs
pz9baZLrXtrBMY26bXChhy1Kg1J2jw1fzhGNj+fZ62c10EQbmQYv5Eaqc5xxbzzmMsI8KLjYlieZ
9RYUZ65ASUyPnLEUU5fWZcLWueGL6lZe7mO33cpHl+nDV5cI0zL/3wLMrBjl0BSRqMo1EBSXCVpF
dey4L0V+tzI4PTmYgj/A7CihYNIPufMdfIjuekDfpyqjVLaaMgIm2GGKTLxSJlBGrUfN+aDzVjFG
L1NBNg69/m1MQlAoTdWmMObC2TEdW2Eo+2ejmwOnbTpFiHzhWmu6xNK/p5VW9KL50EyCDchtlG6q
pPvXPh5cTfiQ52dBvEEv/9f930ONHeVIEh0gFaJFu4+9kI5TuZQCc7KSi8Hg6t5iD9+VEWtxnJxn
C031zjd1msb73urq9tZTAUc5Py+ztfoMjh9ue2OAnWMZqhOnQ2Ao4U8qz0R+aCcjPRsGRInlVtxf
B7o+o/u81KnxtRlt7GYXFojlHBfbIPnwjYzTafgLshbzpwEFFpxn4U4wlMw0iyIqohOup+vcle+z
/Ec33n6VHcQyBUJPneInXHvC/crtYmYO3bL9eogsnfzFH1A/N2+g7FC4JklBe3odf9WMBq/Y6wI1
NirAnhbR417q32tYaVp3r9cJqPi6ki/rSPvWoXMEfhonNqv+h1LTHsWRVrK42p+x56r7QYZAWTkM
3nvX1v2m3MrY60p0xO/Qetizi9CT+INcPtZcarZXvddz8GI7hZyEl+x9ofBSoiMXmRaj3F2VbyH1
DQa32NzHHMClmRNSdKigHOTuzua8YupTNYwGZ4GSlgYENq/2ZKUyj88/BfO9u/C+aVDXgK3GF6J9
4WAepLal4uuyRuykmMo3F1RKa+4oQnugCrNMGkOHO/4bkT/0g9ObFsm8yO9EvCfPN9LxjWaPPq2u
t1T1ME90lgzJlbrDeeDhHAUtHUH81vgUmksOKPc3HENmWHe+7arWsBplA265CXb8ndvknd3ip16r
lY6k4KwcqAajkQNL+v3MOFMnNGMd0O6UFCt0VWSadmt7w48kuU/Z8IWzNOslIYSl7V0gopK6IQ76
8TKf4nFtktol28LcF/v7VRcwPONK1mYs1M0XXuj0/oaSHqpt82NVq2uCJQazNDG49qG65cQX7UUa
UjMhSSt1uhwqsjPYEQ3bd/FfXdSx+3uO5lj+Zv/I+8Soez8lHoNqRPxt7Kfo3nHx+D2Vfur7vJn4
JUKHy2rHYpdmbwarYbslzF1I/f7F2YEwvhxsy+CP6HZ4XwqN6trzYGhlHY26hmztPrjlMO7pR4mm
5lYR528M9GLpNiboffwNRuQ/LqA5fy1OlaxhK+ZxzfGkcbC3U1o7Cwsj/HzGRfWXD7M0+5j7Rcdd
NepmbweWLIR7u3/pbiHcPayjIYUyLM75S5Qlkkxi/lsz9AQIk395s1KkuWBCQ5whFA+uxNKvxPFw
tkHljMF7et7lrcRXxQqpBVJ4QiZwbXocEGHJ6iQYz9UWsu2U9/V8FacVsW7zWol9qlTJ55ntaJ2o
LKBnLqV6CCmiATW5yA6pVLkYbf63x4esgX1wBhW8qIEHEZemim0aVFRkVRVFXBp6r/L9hadvhqwD
YqGCy7sp6MYNKzL5jDKIDXwuPUF3/scBKykxzabM103IfCqNV7BKYi8ogWz/bGWLuyw69DOR9j2e
gPV2T7oRaePi9lCKc0Mp6L6a1wMB9qB90Jon+oBNnptkcxL35Ge/O8jviGsKEPkpituRKum7HSiU
dDrUFas4a3iLmqLgnaWVlYZePakpR7FBDJ1dxkHqgLwZDXn+ucUrNT3ms9aja+9SkbR4iwlS5Eep
jXt1VhJtRtfDP8PCcnuI/Iu2nnHaOpOJjnk5zOFPAsQ7fJqj+xl5BdBW3cgcdadk0MJssdOcuonC
CWq1jiGA02e0EnLMghOMg9tbIblHzYH2cXf0qFo4HL0cX7j2IKzGR/FSkZ5a4swRYrJK6FPlNoL4
B3ot+x7MhJ5Rj4CRsxaPMNvhpOBHvAQv1wsTQwwFJS8FXdGZmOYtqI5jyhThFZBF6EhBN4S/qH3W
OEuHqpyLaF0gjkv0w9YgXsxwyBnrr+BH0zyjUuCxo1aaang7Dx+f45dvw1fdoqr9bfpXXC77DAjU
TJ5scdTPtpzHd+NHLdSRPzol5fFflMlfYLFPC6jPAIwmG7fjmxkdMNBkh/62b2WTwgNJUuFosUqU
8dkmcz7j/+2d9WvI860iHCZwUGsznjMnFBZFRATp3alhszIhtEx8dDpZgq8r8GJuz79LB907qRS4
Dfqq5yt9Hujx5A2rW8Dbj3OIANR9GFZAbn2YvS7W99qJKL3E6FEtkHkUXwA1ILsb8KBRYgUg7dUD
goAWAAh+iwzNx84nPIoT52N0t4ZWDGL6tEQ5wswXjA8eMXffav21/bkfwW0Odjeis4Jr6ld6qKrY
5fTN28llJKKWYdfgenuwQ634rXejMe6LqXL1Y5//vPm+6uRqUYjfEONx/3uysKyujcLahzM6fWwK
NQE8YwiNcw3SsV3OTr3SZtWB8iiD7YmRSL8PAeE5qcwur1+nAI9TN9H6ej606MeMBvYTKHRUnbpw
KYA5grCYeXP9zS48DrWla7DHd7708OgqBRdEFx1hFmyXvduMft+ebG5v2sh8eSk0X8GTOUMAZyyM
2SpeGBsAWiKR3djN3OiOGo4MYPcZHPOp8k2BPwsntOTBx4MvMH3BgnyRoDxgKM9OuBBhTNxC2mrh
sTvMZVLDTwkgNutnFbLCguZxY2W/MN4lvInwyPfY0GMirNgZwI/WUClrFkAmB5MMLPu0/o9+jAwf
D1GAsPHj3VXPxL57Wxkt3ji+yIZRtbdedDhvF5/SWnAFHhHyDFC6x6uE0+JmKHNuNRRKgfYWkTH+
ojx+LoYlaFY9S1HjMm969VdFKs1+r5AJY6cOVrwuoETSHnZZU22uWsuGkNTU+09im80b0kuHXei7
8ezwq0VCJGMpe7ck7CJOQwdjnMgpaT0QSFyGpHDLVpQTY8oXjNl861Kzfp/TlMsfOoUanui9lEDo
FhSnahb3ulZm4ch0B8ekGnLfNCvU/FDS38N71/xS/UyOykPvV1hfvXwT/LoGi6rVyQwCfOjqjkiA
XBJNogxNirdsbuhBQjuhigMD5YZDbdB9mmtgMArsf+ZkzcDICvJvRhteWYuXj52I7ceZG9raR0U4
t8IyQ1ryrLmfqQKn4oLqtp1/6Ex+KsLSmH7QU3KJTIh0BRl6awJ5lUi8I22h6CS//3mHZTqsbdvn
33RjvHoRrQwzaMAMPrqlUzFOXP1xdYBswtASWdLwGAbSJ9o2xfafGNfSbPUd0q8amNcJAZ51pFis
qhwo+MFrdkAaNkF40K+fZujEjZnuBtsh15+XLjKwnIJrD7c5upjm/ps8kZmXz15r4p3MLnpWRKhZ
MlNqPZ1pqINQW/yiaQetkjQgZa66xP5hxz0Nq1hJDKdsQKJuPeIalEaUzaA30WgCRCwRlWeNn/TG
YBD4Pz6dO4QNUhWfgLu3RiglYDVcfQaDzzt9b7wanJKMFjjrbADqRlR6jW9HPCvl6PVD3+jzvFos
fisl7quXTX+1006/yKVyyyu1L4oenOBfLFCxFuP/nDn5sa1tLq3eJfC3kPMa0ZPDPwYUbFOHZVMP
g1wu/RccvqznqX2WY4A4RgelbqwGHfCIgHmQ1qdvUdLbN4GE3E5faEDX66QEBRyhuBzFoRjy8vmb
MEafR+ibMkAXVMbNLohRvPmHq/W0ueXLWYkhgywdLANjiqT5LtFs5Swf0AqjdWCh9V3nDUpVgpxU
GzyoKkBw4Lcz1jU5bXz44ButCkNLS24vkdNJ9q1wkFr9XUUOsgA5d7g0uoRMnAaN51GzYqBSMXMz
Pk+wfzq7sipwWNsAJnKuG952lTOjE9XCJOlaR/19HisFs6cxL0QUc11CR8Ccj0oRoN4MrhDPG8Fw
TiJC7PDXMwP3440DoWVj9Eto/o0M/bc7PWoNIt6GGBqOvyzYq8GJkLBtRZNZuKtR0dDWVRZXbh0y
L8Kc6sgtzIRVzZHWv0YJi5031oCMngz+lGFAYgR4qtPniOJW8xYwk4C7qrZrbx8O9G1DtYvWgNRD
QiaUVy1EJ5gIykbah7+PsAuSXWSoRINrUtrX3JOO4jiCARtd0QTr8TwEmKIbUyB9yQsCEyQ5lsZk
hIUfNz5QPEI7EXZBZd/g8sw5wwuwKs24aY7+oLiMQU1JY4vHoTNK+HDbJDXvUSKDMWljN2rxpodJ
oYTixrFVTb1jgtUHTeGSNrTSQmm8Dlqg3A5T9jZ2eIEjY18x3yX8AHrCEdwwlUfmFSXbebl4ViVt
/XqDiMBJNsFp3aOEBh9iK6/qWJ2wxwEywLehvwyRc6Co2eQ9+32TQ3KHUn1uo9ZMGTkoDzGM+5ka
szH2N+z36Axtwumc76VuVDI6fJNwwe5eGnY5R+F90GinH8s1yRtWgBbVrVzIFkv57O8dZPsT97wk
Hbp2W2vw4FrpbCh0Es9jlPxYEys/f+B5UpkEgcwYCkNa24UyQqg808R+xvqjXvVQjbGBzAuY/jc0
oXH5M/NZl8Im7DC3s2D/JvBd7kkKj5xFczyYlnZhHoFbewbJUkFjL1m3NPPAmD1pUESsUtRmFWKZ
mAYJ3PW6jpOzNxk1miJ86uQzc7G9YRHi0IkpMqcLnLJRF5bbFe7X51Wsie1BT2DldwyMfUz1lvhf
MBDmoD814RJFedHCa/7vdZdQsf13H8gzkA4+CXLhUasTMNAKcjmxdpuSfSq3zBDWMeSbKN6YJEee
PuDdzwC1isZPQDcsKeHVzi320vX2bRt2Gx5aTlInZwTC5mrCg9jEt4lXwIFWDDXqrf25w4MCgv/V
qgv+6Znfo94L+9yC5eniWuVV/4xlYEhbd4m00nQBprfELPydpBbCPI1yv3895Gxkl4T7QgDJhsDY
hO46WcyFd+EvBlwHfRkFukRViU3Wqo6pAiboasRZb1cz/t2+j3wj5xoMCOtGxA7ZgU9utkVD5PHg
zct8l7iOKhkMgTcKi7GkS6s/gEh8tOb36IfSHtykJaNd5lEF3XGFN90O1FAOsS54cGBOLgtCoBCp
iKNxSHUFcUsieud1GJ4/yYoc4PJRoPnwq3f0HLzDTBXjRv/cS5dMZOQUP+ZifT3SjKmr2H9xM5cC
vkBjDFzPWj4aLgR6jXAACc1i1Z6wy55CnJ3Go3+thsm3938lNRTBlsMLnihhp4Lb1AivNUbO+q+F
wZZE2ibMs6vV1hVxoy0zZFdQm2MrWTmyk1qy1nN7iTylIixAtEVm/n7vko6ILgi1FNHcuui85syf
6r2MW6X+JHpojCt19zmxd2RHWpNZc70kO9eJYmYB/62sA/xsOU+1shAacqNTqlRCzeiaKCs8DsN5
USBmQrt+3+R/HW8bE184u9rM4iNnNezXgVf7sk13Pzl4TTMir8DxPQPlJViwj9qj8Qn+XLMjed1d
M+i07ty39u8gVB5bHTA6p3BsnIQsM1tpq4e+r+w9CacoBzwbklUT4pLsuG50evaIx754rt4ZdJQk
KzbYDuPtAXXlxHx8z3LCk78fY8L5NI7vhUITbF6a6onyvnvxJ3/oXln6aVvhq9q2bNk2cRufajBW
QKdvDEXBMvmwphX2jlNVjynay1rlzAqr4xyGnjhIgFBxwJ2YS+LHcHhLWIvaBupunijz6z6hEcwJ
hSdHBZFZB+V/RfRROSFRBWaKxL4QHbRXB1T4Y3NLCuEKB4do9Ud9pFf9291orkjgsZ9E0kmARzWk
FYksj5XFo4sT9LN/KBwWUrjQfDid2SC0W/EtJAwWSdF7F3OSf42ZuPiICw9ySgGDIFFdmt10W2mv
EhBo0rJHqd1S/aSWyEgypzQ+XEEhyljXpf16uvn6O0APcVsNg8ngK758cyYYCNd74enqhtcVa1AG
L3m2bxg5n8YBVpgr+sKrrGZIvd4rY1kTgCVr2TLdJxDABpANTK1Gasjb7j1QJ9A+D9H+dobcK6lP
+EyzIzapPoE/XfxkcGDCGpx8yXsRReQBsGBz8JmbBDC2pqf5Q1ppQUL8bwwuNXAgmGCD1oFNCMO2
kVo5ai7hrsGAcLrNZ8krwQD3cDLQd+c6nd/XY5Fe2OL3V/yUWg4p945bP6zomIeIbTnuDflxy2Ep
4OsmliVSIaaKE+aQwvjQfW1AiIU5lUIP/9IKvcawl6vOiR8wAhAM0v9KDns8IohFnGAx/JIuoQdT
9sRenTQsGZdvClVLAHbuvKXXUxrsH7Ewb0u2Vxo/OKyglN6Jao8T39eyMrTnK1rd2GRsFDHvKHqV
aw4V83Errl+CxjAZJZj14wevClN13GDx+UkP6+mEi8MKML+t178K6dJuUVxDrYhRufi8/m0I/E1Y
SV2tRF8vkUf6XwYuOpuo3sjOVwjm+LLzWAD38ayYB4cmSR8sS2WXSCQxYQtYGRtUPAuso97D5Wte
VtZCY8XaSXeZzKfqssK1ryTXhqD37heYQRPVAwIoSLuxQiHvdfQ8MWQ/xldDisG6vrL+sfJ2IjXd
UyttQcwPcAaY1o53S6Nvon/H0lr/HM0kYPvB5na8DfLB8AvTrr2/Aa4eb5dL7uOVhb84vbGdI2Jr
FJkwHlk4rLb3XHGpdaueFpejcNHPiPFty+eYaaau1s99QwQJdJPBnjc0cd2xy9u5oos7dlZqF2oy
KaZaEw0piIrruwEu0blPXZ2NMhWTn22r2vEYBNct8qCpjq9/W+b1+xCMADUXednSC+CW9XVaChZi
zjHzVM9STVtOx5LYbaFDW1zuMNl+ZOmYlW5r6AFGVRZCsZX9C6/jQ/BlabzS+Ble2BNu1a6Vi6Jg
u2od3kAppOarnvVkQ2ITc/XUQjJdWCqbWTVvh+XOlr1TAa6zq+ycGLSCDq/X7ssoH3oCCel+4oYI
h+bdVfOaO/yI7TwP2bT4kpnEw00PygvY9N91SFviXlmRUrxij5lWhECn6b4tDlvE88G6JtZnK4vA
AjlcTmnYTITiv2ij1XFnR+3WjyX+weZSLFRssBUvmwInDK/pPbPdiPbpiVnC/W0ux0tRfWHMpPVv
gcxOmV9b5IoKTk/3SSBs5kKXaA9p7UkmXM2U1MuP/3apkQSn0q1jqu9aeyX2XovmFtsO5jZrjQ6x
U4SLMs+W7rsbB1FKPcZlh3g2jIz6PehRzuJqZYRdpSnmwSfXKJeSYAc2ZwClnUARGfkB94+e2hcq
coCIg6VJy8IP/j17bC1NFGQEydz8y4g/Gf8MhsVIcVhTPhvtfsgsPpflEn1T7JFBC+qKyMWAP8dm
tioUnRqUeiHJOAKxjaoWcmYf2NhGgEbqWBBi5sH0K8quwcvXrEuwdlsQcC5Wn7bpZGflNW2K9E2t
f5+MaFtmZSCxKAV959IQ3deFDptFsU6Kad2VxQkhshsgMkfKAE1c0QGLX/E2SncapXd6qW24me8P
rFtEQ3FSQd5e7mewetVf30z44qKfvzW3DDunA5BxSJbCxC3+CP5GUaq2e82JLQN9zxyCv1xJz+Oz
O4KzJqFnKJH5EpxUOXEtRvCd+n+X4YEqFHUr028k4vuecpEWedvRRKJ5k1uWnZ8gT7brDXBoMCDz
Ik58RraENrt95Nb3Oi3GZ71afuGifYCUL8apbRsODXBWH6wUzx/SlZD84Bemjv2ot4Qo0PY8omER
FtOqM6lFnxyj35Rlnu5YrFXGrxiXG2P54SKZm6GlIO+pVKjFdPBgAUDDJbkaDRRj9252OHttxQ4V
HF6UCWMsHRzPTJUUkecf8VJVGJ8Fg//Srdmm1Tau1mx53fkXhCnvUA7PZGhD3Hf3qcdymTubbSqz
63fNGVrc8abGlPmMQQ1ZtOGrO5vVDHA6GMRiM/i1F6veb1PGzj34YdbstWVtvcojGU4NiLFthxPH
W4sdWa1bBzzgmffrhXUbPkKT1y5K2781s44+z53e6zJjG+rs1e7isaYQZizuR3D8564HnQmrrOvz
mqc1qaE4w/txpTnSqDmDmGkpGpBO59Cf5l3orZhX3E8IH73uMK7TFHmgf668jPwF7bt34KhoNbqr
+6hSGrJQP5SdfjpM92msPN29yVn7EN+VNRXpkrsMEnZq6tFlyN0uMAelFHSeCFjiTghHaW8EbCWj
p9rHaO/3i75xnjCFLSoYZ3t2NHXjpsa4tPk+GlzMHajLJwdHyxRQPu0PCATNc7Ka+B+LAoOZ5d7O
BYFa4xJ0fYD1IkSLuYw6l165F9H2YZnzMRVEYfBfZi+HMk56Bk14909vWON8RZaxnbS0a2KpTtoy
IC88IGWx5xwY29KiZtL1CtVHKAiSkBxNqY0sh0rQsliQtMC55sP/fcTOCMNRGyC6LKYWLGubq4zL
iRtO7KwGycSFhyxNsA4vdGa3KfD4DCTVSycPLaKmRHx7OY7GTthbuburY7IEavrDfgUxAwymamPe
fhR0LFDnkUKlGfmEBq503QMc64FiOrw7yY0kJrd03UL9gvc2c6B0JW2oPBFLpBpC/izIz+FV909N
mGpkUZjKJtUgBzDWtwegCWzBZntKMU5giw+R/qouowh01b1xrLD40hYEEo4NVYtYjeDjzBCOYCmE
SBSa1C3rxBbELvVL8l4i1y9a4W65qiGNEbpAWKCu4oWXQ0BjpkJZaj2UBkzKmKiFwAbnQKNxND7+
VKUMYPSAw18U5jL7Q5ATBxhzK6n6e6Rv2hbS3CZW9EF+SGlmi6aun7IDHAIsIPri1aDCBOLMi6jj
MtPXgRNfczQwo0ODZYcqL0v5YAuGKdLl8SW8SsLpnpiLMAjuunZQxewemZvErJI1uvrrLLVuhz1u
Ix9HxahTuVx/6RSLaFBDZp1om92UNYOqyT7mA5IEHdiVZabkYGVBUj0di9EFH4HX4RNl2AAN0+wG
2WaEG/E39JcTyI83MrZpHqm7TZqcxwWct4mFc8n/1HxmfEl/6cikyMLE14y0ZsAL/t2uQACIBOP0
fiCFeIJI/BZ+231EeZSkZnJcIFyi9dFxKO2F7nur9E1/nnQ+eJC8xjIUoOIRPPrmpqmeq/87Dzzr
Z/YVijAHPRa50KdccPK9VizivnjOPRSYR4i8AFANHNGEbPgvsJqqksB18Tctv7xET3fkQFkTvgqi
uNeXHP4jKe8LGIlQnxr5EfP1D3UR5It6jM5RBB/0WhJEkH3dR2G39FuzR2Ue/oAM6PzblfhMRgBQ
xeTA5lug6YBI2rkw6jLlCd5zwdbL2EqX23AjCKoD8k/xCfNzB+54vlWQsPpYQde5k8hPSl4SqIbX
yGsDnmUj4TTxEePcPbvRPik3fwZ2ynLD60LJvNiv7+zXAuUBEpNgdF1AQfT4nd2wAAjv218NWPii
N26Ig2o564l9y6RnfRd6kvfjU2TQfWUC6mXQpNT0vviJOhB+zkipsb8hT6JrPLGILdUqWRh8tS8/
iIM6CiZdH25O3SvYenG6Xigyf+QpAw+xKqH6KvE7DjGrrlRzKsUG+KW1oiR8zfiie0vOmsPfUecF
zGetKs4SmNgXtDyREFHjM/XZdc9glgTsty2H7YZyTe+wRbn+whBl0iQcw9PnSKAIg5pOzPQlX5vD
SnnMLfLyjO4zTDOrPjRLdaZT8gFD2D1yF5MOVo16+4oDl0zC03TYd5yd0F8frHZjIb5Rk/VHOvEF
Gdm/8iv2QoKDmdQc15HUGtqRWBEZMHSUlInqB23NXrV7FzHjxg7qQ49KygRyLnHIpzlbrtP9vfLT
9jR3mx+kQ3yA5flraa/pS2KcxaNzLg1fjGec7yq4u2//DxkqdF9R2LDJjHLH5qnawW8gerx18D9g
8/evA/j0ImZNvRsmAE/6LxJbDquai8wTpRRLAcIdXg26ZIKi5SfZKhLFCrptpZSJ0oA22sqGhWwp
HMiozs8EE966Di/VWeDk2cFCfiqwndmaAUqcC9ufTyA4/HUc+dIIrZNsx9DZo1xt0BReKv+vlHUR
x2y7rG3hYEfe6B6m6OyySEmx3JXz54ZRWj61H6V8NTLLpVuBDx14qQMmLLYoUY8WWAfknU0c2AnM
/y+HI159EY9xubV1nDy62TFqo3rUTII+3xuIKVTnAnJDkJf3PH9v232jD9S6DHJYAOp3zvoDu6N3
7ora22bRexpgh9g87XLoFWEhm2plvz/aoqfBUsczznaA7s3Z2gQzuDZNOTjsHN5xGLfyLHJEXYi3
WXoe5r4MEyH23OFjPx5reoMbUYB4cuR3GGybZBV2F0ZW4CagZCAuHNsJLdKTHEdyWArqLU/z+Mf9
aZA06Cf881gqqPT+wFk3dyIG9AV1ZDAlAMueTbO/AvyM6zkjjavZLLqgKnmPg/eUZKd7CwxVG8rq
dvxL3Up/dFxNmxTjr8u/ZXO2Qo+dZeG1OO6IN4lOf03F5c+nH8MFvlHmt05ZB2/kY5nSFWUiuNYE
6QA7SKNbf+oyZ6NVns1KrR6ZZMO5HmNtlSStM7Ok0mYDEZFTE1KXegKWGXpo5htRwL8qkVFOgjan
7Yzb8v92pGttEDUnAuLoyOlkm/xP+fitR5H1LEwO10Q3c5IngGRum9r6Zsc4mFAAcFw8fbVp42td
oCzpS7pLtRDgm2bt4qmB1tZpNnKpaKaxoKjRQVLdbOT4VniFuX0MtrVOSkt/8tsGaQ7VD/YBHJHO
SP9RV7IQXNu6xxS0UNE+pxA20kfmL9kpu1svwy2A7RTjQmI4jDXXtidI2n6AXIMtCuTNl/fGTNtZ
OmihOX7rl3JTkAmzdZHrHb8AvNWSQj6HdMZ68Ajr329y/JrT7wkzF9Qh7uDsZqu0R61XljwQRoRV
Wla9JU5+zskWA+SIlp1rfPL11MtRYuTsR+Qwgl8KGLAN4mZpFKiyF8487AH5bcWy15oV7/SnFaF9
3WOdiQ8y6Wo20dQ4o/vGETPsPcdc/dch1YLkG9En9GdHxum5GSbT9uArzTSCQ11kZSrjd/QwIn05
NjiF8pp380/rGqjBIQ7SkQhEEER0zLlgiCeNDdeiFRecUJ7htJwcq3c97wqE8Jygl6m0OzC/OdjN
9mQR5Uh8a0B9Y+/GnhjRjL0x3stlclGcJIOUcD/TZyDE2yURx64nZxed4cb+4Xc12oeBQewuPPVM
8inH6ExsDMt1k6Ff4ExfhfHZGEHcfHJ5uPPjP0X1vGGWSLXL4M1Fz84qRFiCylaXaI3098KPwUgC
aeaWHc7pDDebf7z1kTMByfHSjflwNiJUhCheNTU+F1ikGtMim5BqxS7eUpkImFRXC8XOfRUx/Dgd
fQo+OSCNxkVVnh/r2b/HI8CGQvIEIU1EttQHrbKZLdwtPxiWDae2qLyCzL/kflkTtXEGy0UkYcA2
nQchyrKM8tvyDpea0XSURNTwzuZyZvIUO7jFIVrrz2VjVnn16dZuno2Sf3RTnYscMbHoXyFtEE0x
UcpotXJVOFEjfVeAh8gTqYsawLJKCFQUC42uOEuW0fF6jf6jW9+M5SjptHXJ/IC5xg93pBCEhg9y
MmFN7E2Hcsl3m4xLNyJjaksPnajnnMpOU8DXsHFjWvR+nDfu4LzWofFhUpzOlcpCR8+hQSCfc9cw
aGVbDT1OIKaTkKD+O2e1fryOF/CqDnAIi9PcA6rBnDdsI2i3VL6KkRQAPqE/f3/YSCPrH2C7wyP8
04QPE+EhAX6UJUb0wNH8x4mTHKzQrklgrzM038UwrygQwG/WYI+Nm46AZoDJ1Rjr265VOUG572pU
7sARRItFCMtl6g55ixL7eCZ6e5OIPn8NUYaB1e9d+LqOCumijeiaXIz4fyqe2mxBiFSds3rU52Vw
80GxT0fV4reSqmmcZHRzBD5nKKRCbQ8gLWK5nfX7LIbn5F8izn6DMpv/jUEtbJ4uYAXoUfhtb5/o
CD56LY0GqCYOKSNB54hU0leuqkEz8fwenHnOUTBWaXyNwHU4aHna5PGFIquaDgdBCqpi3d0jU4Tj
lTFohIlLberajDsxkT7O6iCefacFxL16Y4Jz6oZ6f3ynNnXoX7unxlbUWgXgVz+BsPIquKcoFaEa
RK8dgWO/g5TSZAiTMC4ha+rs0fZqbkIJGIIObQ9YUJttI4QNWOS5umfzCYNuxKn+2niZKUQ3mw29
lyNcu+Wh+DR3TNH03vmS7y7fwXPmt1g9+PIeohLVk0ZauJ8e0Jf5J0ep1c+7goJE//PcJU/MXU50
AZ0LcwnogEGf6FJ+3TFL2Umim8ESJ563I/o0ii2gwvHYE4KrK8r+xGoP0pVApcmehFck5BfxJY/7
dowGPLUy+rEgP0NIB445rNMQN2dzIVmsTYQVlZGR9lDOCRL6dtxF14TpvFkyevmAJ+vqlW/xU0nE
7U3p5RlwhSKdMEHjoeLWiKWk3mXQRGslU7CkkOTsApZjteNKwOmabs97gj7odmaCXGxr1k8n8gQq
2mDOMiLMshwg7dvL5RFXum0du597l0s7eWnNLd8Eovu0If89gp/zSsVrHhXZl1u2LLnxHEWeLuDy
VhKFgpjruxena3rtaNw3SruZe5VGOeLnF7WLFhRp4btCo2lf/X51NtDks8BT/zczI1URO/bN+Jav
ve7/WoZLqG2sdgIM0qvQhgwn264TPnFTyksa7+zWQM/gIjsLdWO6HcmCrgMDFmhKvrYGM3XyghZL
yTsR7E+ux3KXnjlJhYSN+o82aFCuFWcrQ/aR93dw80L3JUH/rS5o/NgKRg+0D57NEq7L6NeyHxRi
1g4F/3set/gAVDAUX5RvtDypEgbhB+S2FkgniZdbaBJEfMJyAaXekpIpLVkdhbO+g6RjZFFcB5II
bv7BKfgbXiQsT1iERXeBoW3M2rSgXALQUqHGbjfuGMpfl+3P0PHVckhusAsYvGm8Es1iY+/bSgNj
IALHYFAjlQw18i7ZMQ+wWW853QTxB9AraV7rGTp5fBYbLoANCbWbKPyZvIDEBJN90pmD/m0WqwyL
Ho8XdkoywRTGR90MJVfR8oMNkmI7hvhvZa0k604c8bONk+rXclmAQqm1VXeJ7/sRqqXhuZwzleSm
fCME4USPoZxvj5CQIr65LYZR3Rf00ghEifdwbJ8RUsvgP5i8AR6XjtY2Oi30jyPZpe4oVNIxdMxb
0BB5TDS2x7UWbzfngs7Bir2PHn/kpYBPKrMEh0GFrjs5+dvINfMsx6qX89UDkK0GnUMmomOHoFv3
RbTOsFkSN/0tstY7w98v7CStlAhbXyLC99a/VB9oWm7uZIE5+aSOu+DrFLEFzVrkIBmeDa1304+S
+BjCiEITKN+PgU2sjgMkTAAxpgsYuZ+LUQmp7kcJXJeEeXoyPQH6sq5I0hUcD4yVi3ZBjZewe7j4
/JcXFlZjf7qgFrgtYPASLREsXbnjR2awGqleCb1XTcGYRTODrivg+7g7zHQTsZs+F/lGzd5HNdPa
s3Wb6AaVMEXiAGS11mYERtLJG7F088QVVxTguXFsa3361RAtXbGBVNamQBawWBrvtJfltmLQWEue
pesyEZnKK2rHT3EYoM2hKnLIbInDIQLVR7ILBnYnxJlImG0520YLisRSspJd+NTLqsUh53StNDM8
qExCeGFcbqf2TK10mkRYE3aeztr1DmIoGV1gNx9ude4AtY+5XTyJenDX0NSA5uArCT4dH2zKwWWP
NDEs+Pbl1MHBc6a4XrPTlSxo1wFbAKdZQeGsTRU52gNwnig56uOMPIp4+hbQDGIxkRvlzmP2liqU
FJZhVeN6dn4R4NheUeVZ3uWrXDTBotiB0VB2J6rc5fhMyNhb4kBxxzX8gRSbYu4Xt7+4S2jy6XxN
i6974Dv7NjS5ikQFpXNC7f9qltHlBdpoMmx0zf0Br0QWYLYuXlEqvqFmaGiyUzpSpC0tJMouzrSE
sp1AJGqLEX0vGcbbN0r7LsRgd3UPpv/raxf+sI2G4hFAShwNEWpFQTNs2Q1ljbQHCy2UgBQ5u6UX
w6NSODLhztl6guudFk4aQS4G9Phi2jWtwMbOD8h/gYlntqOWA0ohUAKJpXsW/TtAUTdXp5ZOFQ8V
M+PmjnUF1fJL/WssI70vpMtsZvwCjGVRiDD+07HAhA0z37wvH/KhS6L8x9BUCzl+Tlbtd3iaxW97
h3aLywOEoCR5Rn+X1WALMDs2xUDq4U/gdPkcJU63iSObEDDJgKUY6M9rKP4DkrDHWEbtiw7czXNA
hzvkX/MKkk6srVMth1sTDfzIkx93f3M6sUfTnMjvb3LUXuiXIClo6CXoMcnXird5pnCuFr2QjkSv
pYBofoOaWLlx644K059A7+QQGEjBMpNyBClzyQ6qVeDUtDic6lRELDbnK+5Z1QSc1QPRNGU8fko0
ZqPRMRqc5DISTJTE6kD235lgxzhdHv57ZhpDcjATG19hrDO/8UgkzRHnGq++yj4lTPScXw4VvPvv
tJlIpNkEYNxcciDhLqNNNuonG2zjCBZQDeBllhRXhtZIqqinAoJ/b6dxCfsRiiKsgdrqtYf50sGz
WkVQ0XFuuLC6o4wW7cGv486nuGYISkuZjPUOFUic01KF05lsjQcWhs/vvaZL7xI0L4I/ePrqzAde
F3V4mbCztgBAVHZCPhW5AIv8ox18C8oR8t/1o07KzSUmP2DYXD5QeigA1PH28DtsEiWOKtfAse+r
3AK6tZMNjr0oJTvMfw/H2JQDYnEWA9GouO5M6vWTEh9w4BK0K2sNd/Rp8jTApsosRufq9klTiGcK
d444yBfWholpwOwmLoJY9ddxVumoICQyt6ZYRo5dG3ZaRGq5h/nr1k5llF/nH+PAAM4H8FvUaM8C
albYgnPMvqAGugqQUTFNNXSOYGRbUQKBpXpcat25lmqjAhBUTbR/YEG2pxM6NPAjMz34vvq4MjB9
6i7lGSSJaWD4rXF3qbs1k/aJ2aaKc1LcmkzZdk7OGt3bWG/7fefMeiDM6w5DqHNjWteRQ7DW/Lhu
AFMoj7tbJFmuPjc8D/2viy33z+sKtEBbQLLkP5vcIs6Npt0JUymP4vV+kuyZtRqucvWk0sIoEE2P
VUOhszF5pOwOSAc+d2+s3YEAmPstr+juqBwUgUv1RujhwibGmRivacFcQXYlq7GTsG5cL0n91mSD
rN/7LkkyQ/s1sjljuTXuy6/lnv6knMCoBcyC7Gb1n+X+fT2riLPW5F7QCWhSLJonoXaSSUixHZnj
qSu68lObH6EIrdhnlF7TEE3vsK8PM1YhRXPcXgi/Mltq+Cjf/Qj4EIWH4jdWCBZ1R/ev9xnhn0RU
2PBUhz8phsU2Rg+DOyZ6bqD+SxmREl40h3lQf561Sk78Ke0iyPe62r9DDb+rT1M7TnLpakNR/A3v
BAFeGX9kUWuifppUrw4y/nc/1kEtIZDigCW9igyBlOyLcs5qNZnWlamBQhGwKRvsVWNwwpCg4jjR
nfn5XfOaW+7Zsd/BTXBaiWpIWxpyJhU9XinQoTZDbAr9OtUd4sdJzP3TF2lT8ErDjtZiC+VgmyfI
L5q+09pG/mXROWHQOgZ3M7XXPz7evZrx7W2drzG0XeY33tswc3dvX0duPf7HExoHdaPe6QJYdMZF
Dh3LZB2hdeMycpcDRxd/o9kuwP6PkAMPSYyh19u48BoffNuk6UTEiYg5oD/PlcrT9okfTXiz4fpD
aa/Xvy9MJPALKeRzot7vaYeKMja6djseS6HqNCRH3IDnnzceE060sRcgvvxiKVScn97w4xBLApZ/
rlN8CinxFEhd82ZIqo+JWuY5I4hrEmSVrrYnmr6qt1Amds0p0qukq4nAkDaOXjWw2svIn8Dy9T6g
IaDUzpZU3pOG/1dwNLfT8i3oZjXXgOjqnYMYLT2aK9t7HAxaIfWgzk4ZLS3smtLnZTDwx7VGQsb+
1NOpgIfdFXEnlBkrZlHEtF3m/aNOb1BX9ubl2AfW6/McIiLed6s6AdJmbaIDKSOn6pY+rXdpro3C
B4oLXeX/feSj246X3D6gDkQUxkfMlWqj6AhVVTYRJzptB0VitqVHD9hmFKXl6fdo3FYIU9O81osl
z2DZAn45QR4jle7Qqg6zwiJfWvJRmM2PXtrN8XmREdDBhfYK0RaWPUmBpZyVolFI2ZMVf7zpMjYK
2i0W8rYi7iIun4Kon+4y1yNs7DYPatNNWP3mNtFz0L37u8kJIkvfmFSiaOtC6o5dCyxGAjg50a47
r/Xyrr2iT/L+LdXZmo0qbRJUXTelP9VFfv8gn9cWz+X5PrYXR/Rr4mu9HTZAyesZGctwQINdDpYi
BI52jphuqwx/cQgfcQRpxWDidhrgeiYnCGiS4lxTZRL+JVwSVVjLeVmfLFVUkiFqzfJWEs2B0pUQ
Jp9q6Vfa1eGWdjSbq5uX7bzb/Pi5wEMXqHrsGjYESUtHf9ih7BfTKVWWA3fnF9t+gnD8UcqbaWyh
/2HKcV+ajlDb73yXj83phihFrV+I8F1gprWQ1DV/dfsJ/CmfkfJUrZHHqyGqey7kMzqQ+phr2phD
XsRtC321Fyr+wy3XvHgk0ihC6HQnwJVDam1OX5hDibQ46BVnxc0Fthmm0kug/74paVglLqo3GYt/
cnmU7VjW2+ioJ3vAdlH2XXq6287vPEV38lA0xghADAwcPmgmhVEIQiD5zwpC1x8h2VRCVUUd+bY8
k1uE51voBc1AmQj+Fma3iDeQfnDh190R2tK4N2iYOrR94sPosjioWrYeLxxcE10SENnZVUn0MXNH
OExGH7UpwdjkbQ3mYh6j+p3X7pZpGrMWGOev1NkyGJYkhzw4JaoGBT083OSVGe0ntYhH3kM/Xdle
bAOGGnt7xnVOBqAlO3yG8OOMiwA/Jz1ZXtcsbHnYRludG+YwA/2QkCxg6c3X6x+w7fjO6W4qnPoq
5FSjdTzsie0wknYOyIl2d4v/4FfWw6iP8o1Kw15QOhg4Z9hCALciJrWGLTIWwPfoc6gmyjtz7R0o
1zHCUk4zIkUvkFkNssJJGENjEE7gyXfD+e/FoOIaVNceW+cjO8fS/Evb4S8LNlAOkemnWFF58ATP
zwoCfl4Prja6yMS1CDrHmscLblr83u/kQol392Z23EDfhbACN/rxGTktLwae36uPvObUG/PKBicm
847Spfq2Bc4YeRk7LrtM6trvdFiTjRenzS+dPIt0LAK60P4zmC4lldnAD5oAHggVdhqhjYqmE8hK
KVgij7ODDVd5s+ycZ09BI0cavL1ZAGqSx5vwUHBCWNDTp8ZtFBOPqt+fOM43xfa6dDCF4sQsFxtt
r3rto80aaGzOPoJrqNUD+HC/WSOCWHAWbEqRVZuIjST72yO8TYVjqxlZOdGtrmW5gxgaqNNT3SfB
6vz+4lB53clpGAw8NjUYeITVi2H17VkA/rn3svB0Nybr3mrTC0adfP7DAsyxX2Wxqy9AgI9+pi5i
MYwXZ84JeJRHHFRRGitdUVlGGlspd5tIO+LIKwgvziwwmRtQcgYGmhp2M/IdbcXHHwh1oYS2c8LI
HONHmKSwJGNKfC1Ndp4QECl6NCZC3xRbRaOETUYL2J8Yutfnqi7PxbQTByopULz9i/9FrEiBaDiM
df4gdP1GPaTqXQcUKbtTVISX9MKIhqVyVdUWM83wd1gbUo1Iekkclv72UK4oOm8MuWQtvb65SjvF
gvvsQTl0YW/WSDWrnUbjKA58QWKczyXd9bhioVCgdaXTav8tf3CDnL69/C1Vwns01oItpkcTPMmt
0navL99DD/XjbGzof06BTZ4tu0/dMExq890NTBE5EuTwowCiLQmMsr5Ui5QaNG2mgGe2ybmHv3Ao
veNzaZu67XBHzPx7kWPNuw5kZhzlkY5pwxFbcb0Ooa2nnkD0gvbBvRACBx6bjuuLxxA3WbYhqH48
vnBRsCwTYWYS2HjciojcuPUfFRhH61oT5kfaboM1DiYQHQ+A5kyWTHRgKKtinwMfqyYvx0lWs8Ja
F1kDl340EdWgqx4MF6mwZs7qw7zYeGucrI0C3ZzXnptsQT/80FqwbnPBA1Vl5m2uYp7OZIFg4ik5
cbE0pNsu6H+7Nn1IOOl2SvuHR0QB/0vTbldqAzljW/ZLo+KG2aX0TbG8CH/AXFMLJPbYx0l4x5Aw
5HZY7vojgcJSPnl+/sTrf06Dg23abJVDHqWjfdSROWqPKcg4ULI1WO/w7800t44wBwt7MVT2dXLm
wAech/xrcgiEexocQCqJME85lP6uuxVdUj73vrDXldy2ZmUmtE00fnxmtpEpxUeW8E+5enORGGPr
au/NDtdF76EtXRE84mr6Y2VRka8k4jx6KU5KZIk4h7t1/7uXw5XSz2MoLg6bcBUCx0PbalJSjR4V
S2gEN80a1bYeHAzZuMysfMqS4xaPO74DbpjI8KA7w+a58W3NtsEFAOgnC1asn7Mz2PhY8wcdvcvF
tsyskGNYPi75D1UTTKANoRQW+Tl/jXf4hZrEehsSAi8JkEHWrHL7/EF6ogq+4cez0l3BoXABLgsv
sOcIZE1tY4OYc7Ksi+HENFifumA4OeCEK9N+AgrD4tjwqU6rQxSjj53Ot2gVZm0uiTpBC7tGHk/Q
kE94VDMvbPk0gCF0FSnnCqk0ZDoupoIHjbgg74wHYWOZjtTwWMJcSv7C9RiSh4fAS1TRspLREfzT
+DHhJu76ZhrdOUqpm6fNzwK4TRrweOnI3LO2hA0tiGwcE3TazRrL/7MbfAm8VXs9NCySRxeGXVhr
IOmczUUkHFPJ4wB/gVbFrgU6OSO0jsukdL6raOMzYG1OQipDZhgrEYYgRLKrG5X4fu6eAWVwNygs
lFjMf/u2fPVByaT92oWgQVTkf5wp3U2uT39S105kG73ep+IaMNX4OzzFsAzudOGzH+vwXqSst+Hv
dzD7En83GdA0HS+iOYSbsDOo6Bm2BNcq8tVedUXdk2qLrmewa/Vvkei0yW6M8Yi1UnsUfqbKc0gA
0ZA8nlOust2gsqlU67AYmoecsYcCF/KhjkeDKLwDwyM4XAsTinxmLfLLqXEfYNahHcEM6qkTUFsA
SAqRIMAbPYvILASQpZsw403DWLi9Q1ec3eFKjizwHpPYzjGim3ux5UNCVlq/ruaayMHH/uSKOGmz
pXgwe+92sfUUbO2sbQ1PxiOphSrzeOSz8w/KvAZFCNhCPXMdxpqvMTy1kQxgJFRdRa1lvf5kxBx5
wovztMylc5rE0+mYwyAdb7JNT+tSV0uE3GucLgWvoLuad54VhrsHn4je64u78iVQgjAT4vZ70Bpb
fbEn1RxHqBDuq+OFQwH2+a4vZ9McGdByHcPfiLyOvyeN12EiIdr1QtOureI/7nt6j2rq4F5A9Oaw
ZcsIvGpOZ7LB3EystjcEO3LYnctipxhsAGPwHKcvv5B2XQZAz/xhwJEqKEtSYrkRJhuP4iuBCOdK
NOdEkUyOukkgdrbX18Z0p98m0TDiK+Pg2M0f1K1J2qCV1EMB0iALLfkgO9BBwDvU44CJcXrELhkN
KVLHQ9/U3KgJ+5fJRRdXGA7DQKxjZ1BrXredaEno7R6iE5R/CFaWlyitg1dv2lSZ6zE9uU1IDYf7
3SRK5LQ+c61OikiWB9LBkBEBSRoDwvXfyeLwBaXkrpjKkoCR5AI2j6n9M4AYOSTWxq3AgYXk7rxW
ey6rmIIN2JguedezUjtZwo+ZOaSgfuQH7CMxuvn8cjPXYCDdnyV1JoRsfYPyovmZsKmUrT9+B2di
K5fnbB2og77M9CDs2r7KCfOrDjPN/zEJpIo5KFuJxLttpMBNG2j33AYqTo9qNAhnFT64EvpTwg8B
+Ye6H4aIOZIM3vFJmHhBWob7gmV7dxbSfHsLmLkleP8tyIKWYiMcl2gIN5VGHJHfm65f+E41wP8Z
z7MsKTifQME3elBirpEHIO1Lbr8Dmh0oQZHLTWl41ANL7mJLkmkbTAQdJyc/wA8if12By1EHMBu8
vgWLjn0q2Z0LA2ns1mqOVEuSeB/eb/QVCXR3lxIhmnm2he8N80s21C4w+z8yjySWae9AP7aFW5Vf
ILPqUs3ZEi/azC6cV4JGcl5sYmPa+tOQ6VDCpjXry1RmyThnGnhtV9YqfkV4HpZMByfo5OHdR80u
IcFwMLZlysF4kKQ5ex4vpJD30YQA3MOGCbK4/oYfGANsKxgT0bERpD8n7amK5sq2PVyTGN9Zor1M
Q1UtEhlR4Gq0KcaolfWUdAe2zlN2M6IcMaAvLU+wjt/xzZ0vlA/MTGgOu2ZOBY7rxBCQRc0HKDcw
cmr3dBd7bWsL0a9VyxgpZYKAukAJJ7AU8j1rinShcXx6vpRzRJNL9f78NHeae7ZjZPpXqzF4K6IQ
omcEJX12iu2c/jBqK4AZA5/WE0lSucaCqUDAy4ql08DhSe4io2hOw24mjp7ACduIGtaKFie+E86B
9wGUewijfKxT9hNu2DDcWeGpgDDT+JA8+UdnQA68Gs7jiGNgTKwzQNxAeIiW35Iyu8q0kaex7fuN
KOIUfHkawcZQKskXXelZnooIASPVlXyfZrC66ll8PwSjpjDZJhnbMmm5fO+kK3zF+Zo3f07j32F8
zj6lbJTMSTj8BjwY3w8DDAkvFMtAn+umhMWkbwj71RXmygjkCuymVxtd0JP6OfFWP5eIprAzRaCX
NDLAOJ3PvQAV++0HzdVhIVT2SglRJ7yS1Ysjj1F1yKRyRzvqfguL05S2vNIODpp+qn0CQ23VhHpq
ftGB1ID5LjIXCp/OT6xJFdYD4eHaJ0wiTd/0gHEV0iVQqBEaYxUGm0LNDhhSI4KtXPDAHjz3l79z
e+zMsfFINW+u5onUxP8yW7HzR1JuDDKXsI01kigHXBzCaQss2E0DOLzCl68f9Zerc4YX/0Oq/lnb
j7B1eDqaAQPbkBlIwjd3ejem3V/c92lfdEFqzajhMqMLszl/L9MjbssCYtlu/+RHqONYlb3EIgVg
ZFIph29WFAAXMvsFSxgeIl5eR2zh4iPuCxsoAePh96+9Kx6fEp20hzTDOPjL70UMb2lSUkfDewKf
0D7UJvCnuq6m4HMjc9Sd9nvqFdw/TwZbnABdgqnma7z8IpUnko8pawQMUUf3PhrswYYYOPWukVCI
d0hu/r0RAiYHrRFA8MV+Wys+B0+S7+X87buMiQnzqXi4YqCRl0V6EII/Pd8PHC3XvZRw4SdmBMzD
Mdiw0j4f0nO0GudcnofKKV0YIaWb4LF8QlfDZSOCo2XowuXI6+263Q1/mitP9hOaUUuOoB7mfKZh
AvmNAm3fp6r6YWO5PnzkFR65kc7zjGGtsP/jjnWuytKtmsJTuBbqh8eqflEOxGpFDYo1T3uppEAE
4KyzTmroUrNRJZPcupfPyP6xTVQhtVZLLEdy1M3UJs3kOzVM7TsvR4x2dDCfTbgcUf9328FU5cEL
46k7eTUVW7yiBWlY7pCiU0SOGxANDE5X8onNMLq+hDQnYtXONAYHwiaI2DvKqitniiut3dce2sws
bOhwzFR0CvLhBmPCJBqAkUJ/eVnqQxSgCmSxVDH57p9wwmWrCse2N2UVMvuCopZ8RNP/t/sL6xZW
fmyGjOzVW55xvnT7u9twxNgvVtJWyUwHdrEeKhjvzOeYh/TvMZVzDd7+d6F0Z144qJaGNv+ZMTiq
f4GBMm98in+ziV1oxuYdqs+BFpuHgcy0jMLfjsVq7f6P+X3MwlnzsAakKBL5MKJvNvIm1ndM1o8r
1ehhTptpGu3ROU9yUpSCX2vTmA0xhd/RYbyQ2jT2qsPcer+nfrD2HbJ9S3zVxpY5RBEhvnO0kbJ3
FkodWyDNTs3chE/DahIcNlw+F2IXqAemgHezpLGL+kPbBfT2x4qqvFTVa/zJo4nERczhGQo1iWbz
A46E+EpgVLYec7qHCvYACVZUMTjDMwaj+J9DPVtxbxvrxaG2AiAOylGoMbYps0afbintytcyKqzV
Aj3zfoT6CxsIy0K5aEm5uoclhrbLbjmiYy3USM2pFjYvXs9ZSFUUNd6DqxRgbmhA7YkUe+Vyq6iP
crz0S3uvHPGGlKAW+IoMB/V9ZTlEA81uMxfYSYy66st7Vh3brLc/gu/C24hv/SZBKHHojvlH5Nzq
J50N1gWQfXxO8h6UL03lsitXlBsFRoDXJA9FwD+X2XlArrExycfTPpDrxMAALHSRjkuKnluXd6jQ
I00pvSPJYn+t2UV+tdZycvpXdA1IucaNzZBheNVZHCEvABYJBb1f+odzKwfZkbkzRnCoZBLZ9CMA
M8EyfoZBde/W83u1Vxpa1b+7KudC+OAeb7yO0gFfdUy48YKpIj7M482w46RXo1IGXd9YBOMe5rMm
q52Yyd5/IrDEPNMemjUncKQAf9ms/cPEHRDZ6GZqOEh8bztXf+ttiQwyMmKgyrCIQscJD616CWS0
py1Kl2co0xfUkJvEvufEeptWwRc1CaYzlogWbE8ZJvZvXMPEvmP696m+X8fewsbQ+rMZrqf5fzsV
1A4oYBKTfwzgxniRTjo/yKUSyMsxAX1jySO48pN6hpeEAJZ9Mq7mPFwinPRvBrNApivfjosqDJWs
14HEkRJxBjkN6w33lnrMgHlsxZprIr5dbeR2nhRMq/I8StwptHc7NuwoYZQv62GwHzGj18rGns31
Zj2AR40xJk4O71Ku6NB/tCWCw+qcqDNm3gy2bsPrrbQtwIiqj/9on4o+b/PcQBMPITxD24ZH1H79
LZ1tgJncPqfW8FnEm58eN5tfKSGaAYfaBYEMmFvcqaQ2Oy6TFfdOHDpW1Yxd+udXy7+Rc2SqelvM
I2WQR4cHOrDdGCGN5alx2Y5BSO5ilRY6lwugncJ+EucxjGlfVvipAsFshMfvimgbnfyTqhF//21M
kDmCpUyfauMAFnqA07WGIpKj6euZo2gdgKnUq+rxmFY6ebMNchxVEmlwu7Lgk0gzzHY+Q0jxjqfv
Fb8LMAnfUIqig6PYJQ47Ar1dDCytRvejiZk67FBApZFd1JFmMHzJv3LTF+GE2ky7lrX/IZGh8TEC
uTviXze2JlwiaJJ1TI4ZdCdwQViK37P+ZZZVga2povpua4jrQRb7DA8ZJyHqdzqJda8miXTUxcmb
+0gTMK6t6ADIxLCOztZbgxpS6LyYr4ku9iTRjPJj063WRjkeJ9B+OWjwK7N7JKu6ddcKdUgU5sC8
PSKWkX1wCDGkZSs1pK+wGg0qFz2X3c+a+RQxQuM0mCjFsjvDffYoxtQvmXyOjecAQoJZUBWqijgc
nUhDSGQkPKgWqoKkHZQPY4V3+48AUmIV+1AVTOIHooZYOldzC3BHj+eli2UzRjBykrYImbF2MWUx
520S6STCrLOKGDYCU5TTCu+qFlmEC1L2STSUzzun4i4yFKGwsXTuSR/GCr9bVQ2JPxzdEsZ3kziZ
Q5XSeOiCwCrYs+ImIJNlyJdcO29PzNwCsKC3qzibQ5Vpqfb1kRCxU24D2BaAg3T/5xYfVJK8p3MT
s8LBsN6cdRjLZFkmgBES1uOXtx1qGlFEG4j6VleKBFDzvd0yvnZ9mqOSi7QScw1MAiiOU49BPJdB
pGOAkhvTLjvS+D573GEgYjhPYfKfQxUyv0pxqcCr39Z+FuLYBJaj0iC89h3lLVd4aCfy20HednBe
62VvJUCyuqYzSgBGKy5vWqJmPEriw+eU/FOhY00OYRdqG8zy3MzaQGZp8ZdFB/rfwQCZEIoc4J2q
x/22RLpJKUaa5jJHHqxbRQAHQ1oOXrm1/9vR3GjEGTvryEDCJwjwur9jYEmggQIiBuUai7s7k4qM
yS6Tqob9q1XEJNvCJxO6Mgni1d7W0l1Q0JtH3xrq6L7R22oud/LXxg/rOXNcxOWr+A2L9z0mRfx1
nmaioBxrCtoT0Rt0hn+oMQQNw8uECC66gqTXYlcm0VgEqF2HtY3/ZxR0ORH5NXD+tUwSPyKYy77z
MHmhdCtPXnXI/K5F0HLifP27gyWWbPLpgiu2gzsqaRbI/Zc5BbrSQCHniEZxSLPQvgDupwNiHC+q
U98/8fm3sp4Hzf9tFJRDwR+CqfpfbCDhze7/ruFGA8aD6qrnbhNTJiLc72NPSTCJLq444O2yARwI
FG90QNQL+/ZA59yjSDenBhpaihzb9/DtjPeZuJc6Vb60vgW/za24gnOyWDc9RD2d0NiwnDxNrnra
OAw8dWCcs6w/MEr8tvx/jBHRzwEX3Hyr2ZKWJRq0xRfOSqQFI/y1vZp9XIWO4pW2bXNGJDFGWs1v
SU4EDWxoJq+2Tf1sipPRjgq1nur0VS94KrN3tV1N/PgknV2UzuL7gKC2c5ajvuJOEAOSIrfY61DD
Rrr4RMK2q9ewjAFBrvtLu2/vYmk968HY9ZqNPNOsB9O/PzxnF82uZ72JqXACSjD/osrdk+CoXsXW
40/WtH7QVDd8A/r2rqDPx1tGfXGoDxIgdtbsXk9BZWFKynkYJ7H+QVWRFw2nLWsg4ag9U83Ty9WV
+ZcWB+tIEevn/o2kuujnFtnEGLSrXZyhUiO36BORv45Y+qkZgV5Xh2CjmTQSLnd6vUQZtjhiCJI1
1JDsk2+LQhnFHUewg5Helaqu3lDD/6/dqZPIZfQXSdKt7YBurB5BmJ99j0gAAjhcrkIHFx9JQWVO
pw1ZxW2vomQRKgc79DYnCnyCsdqUZO5LkcDOcBgW77v773gwBNnv+FvHk4mN8fPoPo/edoFib/Xy
WF4PyB8yup6PJFiJUBvoKM7+gEkl5YfwdDj94bQEFHPkFNbrq1JwJI3HMBBe1pBypyZ4NhRXxUZ9
DDcw/V87CVUZSCaEuub+ZxBKXYDiHCtB+xhhiWynzwFxJwqWcP/stc8TYT/LK2MzEkCFe2njG/uf
z1J9NjmaO7S0AinVFhUNEhNOPqNHWvvHP5mLGof8vQUCH+/ezCA6h0NO9n16KTyv8/CsA0MahP2b
uXU/tN4yRBYAMwiGaJzN1Ckz/ICtxD1+RhsdRG5Xhtn+MbcJiaCJWUVvyimdpvfZRyy6w38ZM0E7
JxZA/V2dr9DRT63fL0lIJbulounBOD1A09E3nb0G0YAmRuKQKthexFNi20rjBE7eJ9lVa0jNJq8k
w5saoBAhWiLI1FNZLnJCth7QSD+QW5FyMoRyT023OWc7dQUCCwoNWq/3hEyzScjAvhJRMpV2bUbM
UcBPS0OO4wVLJY8l03kLCsb1iH7Pf5xG6oSOl4NnNitKZ0bx9ufkDLfliMhs1Sdg4OUUhohbKoKs
GHZUig8UPrYIzyH/TiAcobiyrFiXX8JBSm7+Wv5hQ9FG3OOBTe2OW3bCg+Sk1W59/5Q1uFX7Jmm9
xEDAUFpRH8VcVFOfbNkH9uRTpEpHaIaIBLx5IS2QtDPb/PoS/CSjCUsmVgnRyoD+8Y+eDIjR/boH
8FKuf4DVsADNoDb4oR89K4ROaFCsUUpXbsj1DIXBeuh7Pu+2BKDbDJxzKhq5BIf6KcjXTGdGsNPK
A4oJA4KDJ/FoubWi2gXLC7xdiueSaHj0tEjxdfIWeokHiGq7hzaPgRLI4CUZqubo3cqHF9U1a3Wn
e1poUWhVelH2LcqKMtMykBljO73Z64qzdjzQMBnY4vK+520cFt7qgH9ZPfoprjnOXedHNF5Uwpyb
Q/Z8eCXeSFMrecg1zGGf/zGHv0t3AbdOETyvwl7VjZRoYdu2McJjCdBmzddEJV/WjzmpFrFba2P4
rHhsk2Q2m8328TFWV4l4kwjm1+8spLy5as+3PMTg2s/4WYNP1ZNoXFblOO2qZmudSa4ifIok5ZSE
i1zTP4O+8CqBKrrkd3cz44G0kTAe7NZIANSduQwF4d39iGNEHxhT1Xjwnufhmu/k5UOgHsFOxtyZ
otLkvpyT3DmvJaOM9GEurXIIU+59LUqWme3pScdabH1/O/WF5qBHmiEpo2i991ZNxcs451yRvLXC
nruNqweArbldLJBd7pDaAcL7/rbTKfzb7j/rs6C9QDJNE+4cXVq37WzBxaiM1MGWGDhOh6GhvHI4
B+4lQVqHhyU9pexAAtWcmO9K3OsMXpa1ZspwPEPeoD8uU3AvRFl54EbiLWY07myQR8I6B1zWjioE
1nisGgt+tN/4vAcouEu5P1gDKyHLNNhGo/2vIqbTAqbobDSA3BHBWp6YaC6SfRlqp+ayYwxvhfLP
189J8TMcJXB8Mji4Q/1AsbnG8xDc2hCSVhO347qenRxhQ537nJvGfLX1dybPQsQuDsni3+jTKefU
/WQDXzp734v/gOudjTHZ2NZB8KWtuT2nhI6GYVM52l8pHufxnYePV4BsGwMM3/kGEcwcwMH8A0dd
IMh32dgxi3QQNX8B/yk4tnlpDl3fFaXZPLR9TkPdTI4QBNRt9JdGJo1Xy3L5C2QX2J0UxrMZoi6X
KaDpxTYejYF43ud9+f/tppoksmWU2Af4dxVo6nj76yUJLzGCKEoID1FHdgSlVKsxXLKVFV9U7VzW
DmEsbf9ZNA91JuToF1mN7hlM3YNpcN6cq3QfTFr1Bmw01urMFC0CaDSwdrIMw4SnmTpwBKKyx8Cl
Gw2nQg8z5B49zmg1Hf8P1aXgKjJWllipT3GRMyzijityX+YgJnsZ5K1OVGBxwprf2Tjvf621dx4J
jMA7R4ttm5rskIC7pSMrDwHXFGGYXMT5JQEMZmXU2d46tpATyzcbAv72E4eDb2BoDMOb9J7fx283
lF9mOYZKSlb+MrIEwzVqjh2ouIhC6sjvryLvaCYiEoTJeTzR7f1T1PquWefKLczBXVL+IbR5DbA9
uWKQWAi0kOlElNkwkGVbyIKVEabcNcHXFM+b0jQp5c6dy4WzocZZ0QZk8EViThJIQXHpEKgrWc5p
AYlRfJ5vbjGq519rF9LA0+QeFstCjFDzyZfvHD8oZMq4R1deUwnmJT8e8BKJZY8go1ayACtmk5Xo
H8Dj2G38jauc3nktxGtsTZ6czXYr2suWIwF0G2HCyEKGwD2v+PrrIzGVIuxPCbqS4r1XjeY3RFj1
PmqF3kcGnvCp58Wv2zvUGsHon60Yc0oZZbnaE4ZDAn5bl+e6sfzMemW3h1PI6ifla/Ub2iFG0oJ6
wsN0wED2xkANM971LzHhKjjlhTTdkGIGZff+3B2/3HKyuxpHlRZfgczpJ7Gw5ZbPnqPSpcS8QCr+
23HVVeC6s3toabQ8tlPqflxEK1GFEWwZUCknjIzI4G5A9PK4/9+UNX4IINtr3tHGu2bvkznu3KRY
hK+etq01QeoPdl8W2D5OK4+mPk1lDaMtwdUZkLdEMs64XWKb8DOuO/RWMPZt5rS/UK5OaK8I/vQ9
N2bJ9rR2ZdlcujSOhrg0QJCRSlZ97BOCGT/2BXcF36LQiqQpmqhdyXHmRoySAAW+lPCD68tJ3eK5
eCWbdGOJlTIBtqKT5VR78mXAwVmbKk8JW2LcxvJYapz87tEFS9irX/NhCBpPOHprw5N12V6e31/X
BEILorSmR2nJqENXCg1ET76QRflFu9QgOp3p8M3S6wjNSUUTiC8oKh0eg2CC82kntCjvOw/9cl4q
N3RGcAfihtSGpSsw0sfW+2C4VtHrqLJEGU9OVhXVSbecctpiu0dTlYW08955DRtZU4otekY4pcd2
fYIw62vwZjjUbXqoKe4hCsjWDcnN56bzHWcOGIdzi4PrMEcbdQ8kt+hFTSpY92wUbCOXB9tWRkup
ekxsexmYwaMxdzqjaLeU65AQemXmlP359Zbxi8rfIN/xgFR0U4MGi2jFqg0/A8fWjkJBeuzV2+iU
XQST0aZk/ZzpQZcATf82pUXmmFFDABK2QTnTssOVuGNWQImB2MMsWXt3R5Hx+oWt+QtPeGqF2S4q
/LaC1JSBr3jF30ZSIkyHaRCKJv4QXzDKkjANDABx5c3V+270XZomS6BlFuPFIiyclRHo6bmM+6Pw
UxAujfAzrqQvyEoyzLFDnPoZWdH35iSv6HBXiPSAy74yu0eYt0qZnKipZ2SZ7tKMEGfBgRHMPQnb
J9cSaUu8Ub3VnJE0Tm2bSc4aVn4MHD74rH+7tGOac5YLBFi5VAH2JTDVVhUbNBdI0Ozx/Z+pV4+Q
RWSiydlKuTzZ1i4SBxL/pSP/zSrEvDRjc/U/Z7Omx11nAPclxe0JWrP7vIis1IPWUt1R+cA6uSnl
A+IPm3acWUbXV2+gqBGbfkb4MzY2ioP11iB5qkgrKFXomH5nC+ODCqn+M1+qtB1bvpJEidK+DPc7
IQ7pNMzAE345zsPdEafWPKsDlxCi2cHgi7QMioiP/cPZ+hzj754YF6mnw94xF9h2ebKysaOsNUXe
10HMxNYvK+jm+VUF3i4aFuyTik//lzrppc2wLzQW1FkaVvl2XgxO7AIcDpiY+/8xCuOpv91ByFKH
XYIXHD+OzO2QF17sfneglTJfnim6+RoYD/dsm9g0aTw077+I3i1LLlR50341VusjcDnJaxOH84VH
Z3pQIRaxdW39UeOhM0qxN9Qf6mCG/HWLrRPBT7wMBCOG32jfCkBNRS2H52nNhr85bwbOBK+BOG4D
3zGK5bFlZEM/a7Y1XPVjy/k2PV45rAS5s4l+zYJRw0tS5/gQQITSbNQInbFUjFT/m5gaAgE17YbI
+2tP5y2jdM+F40oAaL2Bg24cwIS3v6pxvH7wyCUoxTO6FOV26hXmJfbpRnQTeKhNaiCy1BWMSqIv
pObvdPpGYiXMc4ThhV/x2uvb6dhp/+PGhklL31mCmG69OitsB2d6o9WITeBIkqbkDJYTOGvwdt/R
GukgIw7QF+KB/4mq280HllNoCy4i5GW/XwwRESaTu+er1fYT1LqmGBT6hpktX6OtnXO5p+WXN7XY
q5kFhTvAQugrVV8OfZaRM75deg+VMRRF5MLCowAf00IlFqOkeSetfPvseHZN+HZBaL+n1Z/km/uN
JYno44J3YfNxDs0GsrSvhmVUUQXjPlTmJVz1qmcFRl+rUjv0m+5ffomA4Bv4hqFDedIfxA9mGJlO
MDrOp68qMM1hSo7H6GR/gix5BuEbW5Y5unK5CBZVEWwS0+wQqkE0OStSHd2zuYiXLk6NQZSrxFRK
Ru8H9ZPy3PBe8ZowXFxTP12gSbmrgiCzSg3KzhPIWHLI3Su2/23v4fVZzLa33loGJyhyZ/LhfN2r
Q7mVc/gD0+6cEvQeMC2Gq2PFbQLYzaSJ/OjCXxcMHs+fMqDUrlnu4cpBXhOVMPaENDHpeyhgv+26
h71xrVPRlthR4CKzrnbDPGMSBTcAsvVVr/62GwstHhe8Qr+UlFlQM1rT6z+BHmcSzLUJTybdjUYd
Na1h8etp+XHps9rNcg4PuSD2n90tueYsIxzb04mtRBI/MfxfloX9QaxJukRl30dmLHpSiSmeu4mP
rDbQpAsm3hN1ieRBUMezxvpTF7WKP1K+23kpOVY5aNV+uMf5jgrLA1kjQXQAjVOY8EQaOwb0x8pq
mtzPJaHRF+mKGGztv7dHQjrdPEack4HawJ5B1lecyqLUSUghla3iq3aESqTlDxFSn00hjIJGRHsM
0/7bl7ioaHaqZ+OUnPQ9YUfPDuiVD0AFbcNg7d9mDRxH7frvkhzDvhgCbno+nwPMjZxhCN+T8Mwl
hKsWTnUnxbLt5bF9b9ZbmWXmwR4AhGD+jUnutiTCC9Aj9loOQu+Epj5vLkEbjnzVpKPOPvLMCc8v
z3ffvn4PN2qgBbvP22+XgUF7KOaZvMV46cNxDcM2UkIEXjQ5+vcCVVcjt0Q11HqJTV0baapf+7Ka
VHaVqROyHkYqqW6/XwRixzV7c5Vzdmhv6ANxG0jYrqcBGyYAUh71mdmDzH87CoEx5qpO/CxjFDUQ
08n9/Ll7h9WmA/+ZPLMa+JGHzyIS4VlF1Y5lwJ/uKf7/f9eQNXBjJY/WHOsqKQMOso4L+lxABRe+
waZaE3vXZ2ZfZe7sWid+tedGV7B7u59p5hlQLNqegjHdy6gqrLe/RUIFUUzOZfFXB0ddkG7Ka6ih
sarXUlhJQi+HhZJrb3F4sxguaVAFncWKmyx1a7X0Y/NvZNtSFGhrfxzmgpqNFTq/WYS9qgycMysx
xODfC9xpMGyD+mqq1Rnnyd2dEB/xfjze2BSgt3EXQQSs5eSIko37e0l23BzRBQRTQpdUN6QPHcSq
S7DoGyc2hLzJtrz+V2wYQ1OtRSL3W8rD/qh7/h5Ewco/MZyA9q+KSbkd3fPEczzUgOeYoI1iZSU2
i3MnlQq8N9oPqK/iVi+JYZjTuR7FeHlOG7x0FBokGBfJNo3u7+3bvlCreMCRWGRQzat1CUnVk3Jg
GuPhg+GFNOk6LSFia2WDvs9CUTOlkDuKBGKtYBvyuNwzIjZSJFf/YnkDMUbOy9XkwU1TzXGyp6SV
t4bMOUF1RxADtWpugugm0ORlU78KEc51zvZGimugirRnD5koTgUKc5TuvcXGDuPhNBWyURHYqzWL
PedO8H7223nsTE3Jsfmb7zSqVrgoBcoirzTUMFjN0l40uMjzLOtAGefnfKIzBQL9+M9Eq7bnwD5L
nGI9XO0YxBjnyuicF1YxHenlU1e+fMK/j/wxU165oa7f/cfi+Vyt70hKHA3iSInalFOt6iMsZrGE
dWiVlD4xnncJxrAeelWxyt2Vg7AHrcKWElZsO7v+Znz+Ryh84Dc6eJJQfCMJ22kvy89oZcPy75hM
1oXzFXqwdpmWO1aCOtTWYhXidtb4ZD2zYwdbg0HRUDs6STpPgxDrsn2/pnRYoV9oSQriQ2qXp3gS
5Nv88KKGXZpfsSAErADP9GNSiAQpghBb92y6s27rX8M3SAa1uQQPRksNGkfSq8sxODj5Y6PYZ+zx
Brif6LnJ8Uh2YzmyBxQ0W78HVlSzyCCiFQeUguQiwi1Kuwakv7bBT7PbL0An3HMRqBGWV/ml0lto
hWImAhSlQQu99HbzgxI7Ng6G3PwYr59akZlZKWdkT9tkVDBSbcSD1D4Nk3HzkPxUt6+o4xvBvL3W
j2rj6zVx65pwuWqp/iuYKEcR8fieKioESUt7lAlswK2DGdva7+FauNlp4Cv/IsnbvRjFl2mMC1dH
d47yKl/hu3hcYxQET3Pc1lX3fsZjsINv0jiUnsexLjlvNldMSI9WurLk2pCRt0HqALBnNxvceCgm
z8KnqRnAIWKskYMRczoQHTnRjYUgFy2glyPOcA8IvpRSdQRO1NGbV4xKyS6W3ENkmD/Hx3h+X25S
eJlUHiswZgtyLnjAX0v3l5Mk09vJbVtZSna390aYibzOAiszE4WJ81lRUt2PsEqohwtFupICAWn0
MyPrR2DmCbcgNG2JJWCmaUrx2T5rVUeMjfkGOulVlTgEmP4HZ9x554myB36rmUCWTz0uppn8MJCW
+VrmxJp1+W09rRaGxPVLcOfwA/1mzZjls0T7vw9eO9ccVedk+x+PhVc9YMQaepCwd1AtHJOvQ+hZ
joor1H0yd+/yjt11pPkvczVbVswM3984Y33l4uycaTqNWW64JCtPbvAhISCsnoXJeLmDrUMQ2xbn
Eg9TNjtX1HKeafJ2z3zcV8QCYBxbcslP5D7wA24+Pb4o0pWNlyMSwO55DBXkAPcLZMlCGCpOK8hA
NkhXZa8airKD1ZfMrbK/mPwtLF0y0czP0HX0FtVFjYpzS/XRATRbH94mfCd2ujA+imZSzDcS6RvK
MD3IlCwVVO1ZKbZZdmbNjktR/pYufPduKQgH6p6IAu2zlZ0r5H6ELi04f8muer2CDt2U82HTeDnr
k9XD01HOYkKNvjm8X6nJIuxZnKP5kVi+7h7KeHeZvKsjWP0anaDcOR2UJkNDjjfJyMo/fGSIMkrT
o+xFVbzmsdSkyiWDNZB3FYtLJqquGm6vpEHmxyN8eJzHi/rYy0Kv/a+N7zQerjgQcjhU2to0t/CF
mJTEW97XxdsFGIKBOjOn1voGq5weOQL3TcknbKNyH95v6jiqdlP0KqzpciXhCcb56hmRDtBb69Cb
j7rDNySHeW3Gc+cdBhXCvMpfTY45M0ktcgU1DPCfUxY5j9xFPwjkKqnJJ9189TQa3Jq5s4FBOIDO
Lev+JrIUBqp6KISeK3tfamaJ4FO2d2OSuZzvodkruULQoN04BJYXtBoSrDBfTHJWNn+0Iqebiwe8
n5rbdoforZQAh6CtJW7ZWu+UxeAzSeDQ0tWb43EZM45CJSCcOiHHDE3bd1r0+Y5iZmtsRWTl5V0f
qw6/+fCswZ4VrUxFYBUSRwhmI7mbt7fbqhug0vd3IHmKGw9XtwyatNlWzwPinDLS+ZBZAVj0Xu9n
U4MJh4e3+FHfchiWQxNgrD9/Tsik+qKWvh0IVOBW68ToJxnhq3I9TM1KQFIHdVZ+O+Af7p6NU+iG
F3POEghMBQWA0CHhAW+glCrZCLUEubiaPJMqWElze5Tz/tFoIznsfB+c4y0Dhsm3nZWIyRs5NBIq
r3U2kg6yQOFkknLGfcSZJNoiUs9e178aUTSS24nagxiYHXRVmKsVaMPCyHA1ZHSN2MiYmePfAGHi
spitxp3N77XVPTrboZgsoycbFsML4j99h8EfvRrJPESQtUcaPdHLAybRfxQNYNvvYfaKCmIf60Fb
DjPJF5cSBw6jvsLcdaGfqQ2zcSFIZDc9XB4QY0wIdF2jAleb7sUNn73AohvnX5m/qbh8GkunOxLH
F+iPBUxhNE9lUhNGLxGTIqzj87OwSC2Zw3cqm+mGU+Fw7SsXcKARsy0MvwCEO16hPJHKDSZtt408
Lptsk9y8XaNQNmIfBoWyVZ/nV1Jkbcqh/4LV06YX+Yiy8RvUxbzp10ThPzfYlSbpFajHkLrPkRbJ
FnHCU3DowGdt5l4D25T0PhVIuhOTf/KU4TZxny5AOd9XHtIZkAYrpV1cgwM4AySU66iyWDmTnlj2
io/tnioTqq8RWUSUm3ORpIKRaHjDAMSGFlnGew/PUFkfmYlMlvp4vYE5sENl8cihJU53m1Pf+Df1
b+LFIjMc0GDvpTxnwHXjP3jg04xVdjNnQpusoYU/x3p4+kLQuYFStlq6VJuTcGqpMHT3eZCbsPi4
db0dfE+BQozU3Og7q1L9MF6jwz0Il1NG/ooeIy05dYoNuI+ISRMW00zjUr0AA6zKACb695wfwD8Z
5WyNAUpxD+o4NI1G1SANxiVV76i7Pp9LcsOniPfQax1XfG0VTYghkNBXKx831ZVMHoQNFbiZ6FmK
zDug5FRMjEnUB+tpZj4ByHUpFuiB3Qd4wnPqlwut06g4uWuxhiym4x/QvWP+j2Bte8nFQdpZFfiv
+YavNZ0mMPo6i5YVmPtvWnRJti3dyWB+kT0VgToVVibEpJs01s22u+3QR56P02lx4Ifq6mmzg1rY
iZxTIEEtxrCIkpWS7fZEbkR/XMCir33JmykKE0FrMmA6IYGBE0bYEGUS1AcCeYjuoFIywKfQHe/a
atHbgOte0ybugnw1N82sJ4Q+dJrYjD3tEgdoAoByK+rsjPuoGZrzf9GspRGWRXEsg/nGNiQPEMwE
V9kxvgK0MlqKlEtxCkqkHikccoJgQ+UW1a3spZs1EQXl+Zk0gdXGljfREXJntvzR5gYJOH2amoRz
jG0S21buqpw7QnXF6AX15y6u2DEhCsJqUtAYGVQ2W+WLYlbB2hXmqNUUoY+cL4VLlxDHlNwy6Jn8
EArhnuzJj2V0qeUBH1O2WNZStw9knDoJ9ULUE70Ov+Ubj959+7vxlV7tYip17iTyNUeAdJxlNGjh
rwArHnmhzaIPHNhoLI/jItULE6ENstuEtz/SN0Rb0yF25yCDknfJjjNYtfhZOSaBZ6cBuxkzkWT/
WUgW0RSZXWOpNvKwBN9hV/q3nhvtjpTnlnKRHh8xoJWQLMYEbQpVNg+2gKswnYMezb3VgNrXf10N
890ita01N0fnyXl/KRVs3q84GpGqek9Z6+WYuJNdxUgiYh2I71yrQW4uvr8mT9MIEgL6hWcd0Rp4
QrxTaEpNUSXZosazbtcvbqt1CuzgbUVcHyX92Nz6q4QGr58qubaXQIrO7FVcIIX6ijraIArXm6Tj
oMw3wHYHicyduKCy9xm3cKHnkPdrZU+F+9eF34eTZhnjlaPVUQMYvLTFsE3cW/uRF0kA8+ZYq32Y
/YE6bA/xsJl+moM3dRCu5ZdwS7mVp6w1CCA2hu7S3ZkpsZO6RK22At4iNsWnyguHfivMbd94lq+u
XBmNv/5sOysyepqZ2rgR3B2jf8TMVCEI1a9oXvFdh+rG3kVgMupOVtvo3kV6m2JDWRL15wmXnxuN
NmG0+4Air0SvT3vorR3YtPoLKJicuiu/k4NweNHOVzVtDM3TJ77HJxV83N4PzMb0NubjEB+pXj/J
auWbJkBPmRHjQ7hMVYtxWH0MQ36i4h6v3XuQxWlH55+655ki3qvWV+UpVXVREIraZWnoEWkumjjH
U/M4wwAkADW6vbtoWaWPiGF9a490W4/pn3c2qxbnbR/rSw9EclRrHca6st91axWWUmLVo+kWKP3x
lwrPQtRYpJ8FgVCs929obws4tbimV3fuyDLdQzmlJ7vO1Zp+E2jOjMEy0kPxC6o0a67M1pA27qma
1ywI3ANqjwQn/Dr8qKAkDOcXqb589SeUEbSSzdbBbsJv3W8++/41rzT5oK99effC45wfy0pahC1N
ha3lhS+C7HJvLuU3FDuX1Ffnk77Yq/XNSTXaQ89meLCxM9kZTh5g+sx2RoXjJsu55Y4IL9o2339t
v0/XSPTe1Y7kUAQp3gj38JKjpKRog68SNHyRujJ2j28XlSQbQrXOV4e7ajZXFqtBfTHoA1plwBbj
EqHxFOy6BF36jXCu5Sr93fJZyko+cyfnsv+WGi8Bpj2HiiZHdfkD6deintE7x61J+q+c5ZE9aPwF
bb0zTkMBzODrWs/Cyu4bxjM22JrDzOsLkMadxc0qNGKzVwSdsL1lK1+Yc+vHUnZTJtxd4G8LjpEN
E8PHjk6ME8hzJx3Gk+9WT0Nh2YyrDxfaQP/KHpm8oTArQHFefAc1kjCbmyLx25p3xYDMdXefhbXB
AENR/3dsqOubh2phOYftw4oxZ08a9OFrA9E0abAWCD8Tch6n1eUvb0cxXlseNy50cXQe0XEj/gr6
tYaKuMPRpICO5m9VrDBhrHAoZIzYaW7D0U9IbRLMt33aAQNDE1+UktaOqxew0WtYkIRdbOdbTgHy
gdpoHSEhBAdT6pqijPwBiKX4pODDdJDgxwY92y/Rmv1LpW6gphT6DFIjNJLzytmBaHorKyThQgQh
8Z8IqJD9v9GmdIkNjHcKjY6L5Qpts5GZsQtOez3Ci+VAxi2p/TmVlEcBJeQhEJjzFi9EhD4CjNiV
K849sDUnuwjVMvrd8gEgj7e4BKOw1v/P/t2kUqTMFiquRMy/6NGcWPzMctRQbRqLnLHfgXFjuHey
n412MnyQQQt8Gi3nsgHeL/j90Ftz0xp4zRrtDXMq2JuPlivWJ9NJtOFsk9HZexLvmHAXKw7vPrS8
4eCDm5NEqI0+0EYMUON3VJp2sXgQbIrF93PpCdKo4XBs2hZ+swrzDqDTk4psWeMSJM0NLJwtE6oI
eL4ZdlEUFDBqX0jp1mHtRer+FYnuicM1ZByTaMA2epjzGEj3cDkHJhCXS3/+rJPRRdIPXON75xrZ
ygMviNna9NFDVoyGSLTnGwU6hD42amPU8l9c6bRto03tVT9x1QRyNa1vLyFGtymsZ+yNQaPeNS6I
U9GyUriyx2fa6zSaCtzEb9SuUqLn2cq2E7jTE8wTfyVtzbxii6GzvA47iRrTFdPAh0CHglBEeO4c
FV9PagajyERoQ3Kij626NZ60d0pdujJuOq2vknaZQLFcsS8cwH5iR5NrzuleynbX7I0fP+czkDWD
tLVxXrC/MRn9S/p3FEIMwcf0PTdJQM3H7jgwNvpFofVk5DwRK8NaUQxJX923P1irM0f7QvSonTwS
lZ2AuH5ez5W+NrKfJ9FsxGBjVAPLOCt81pfUrRE3tqEqpW9zSjEsAi4YsgB13+OTDoMnIs0/0eAt
5+et+9dEMNaNa7JEpBiK8xf+cD+C7dmp73z1sURQvASqh1ekPt2/o463JxlSRqFj9MjpsNSqFNRo
rElpRXsidU5C1rZcSmCOAQouYOjXCa9VPgA+MCE6C63BXg6suKQcsN9a0cGe6g2wVmlarPqTPu99
JDXy+wkD4yh06urv7/cN0qf/wfsbNSrcY7dWhBV37KX4/9b3Q/zW70qDMPSYVK3xyFgA5knXC8Ow
L4NFmucMW9lZMfQTEpDwBMFANkBfjDgVTfas//KoZMZ3Opf2oVS1z3wJX4+zyq6hTs6Oz+MpB+Sv
4b7ASyI7e8PckeRo6ckg9tbNuZRu71UMt+/l6Xo0J3+qOXE3XtjAn0dedHMAB6eVOBaJaIOT1JXY
pZXUQyKwWo+gzj2+lb8IIkRW2EXE6PC5jdguXjH5inD6BJMavuXhX19198AUBn2Qo6yJrxPhzbJ9
d75EdsY/W4J3EtU5euljNQo+OJEv0s/9GBmrE+nMsVas35T01EhAwngvsE1P70BFJv/ezPfsu6r3
Tfr7a3j4vg+gwpUebba9kGCsJoj2jAjajmKjXOGT6WLzpuTza1ggxXMoxQpv0eI9fJymt1vTKwqW
w2kv7CdHHrDKGEyUG4KQAA80sT2C8lIlmdQC8qwXKUj/q5oMAtzbpFeCwklT/CYepQL70wJ7vpWn
cA6Ox+KiOoaxYZ6qPf7fGWDl5cOgpMo5e7NzS9IcsO+PGe5Yk2Q6m/wpz0DX2J4cwjl4m92If1QN
HXpepbsJzlY9/UZGKG1j3irXGnVTTXHusmdUnOwahSytR2cj5uLdr+ycsNDwhhgqih3evLnWo7dG
mK4kP2I841U9/lQLrJUiKgwjqN7FVg9A6t2vcHlDVGa5JK1cno7f96rFEdw1rX6gRVaEKoZTz8Lq
PnnnypIsFndz7Jgsa3gf390i8SEQkqS7zlLt5iiB3ZWij4bcLtydj3hDz6l4MfH0jy5TLYh2N4Tg
EAmnaueAUdzUVtilp6Ac2V5rf2BOocG15bBefV1dVJCCfpBVM2+doYzvw/jZ092n9shHy5z3cI97
9iUI/cPQULe9+gcFBfOnWP/YCwQdEqFT5/++Ecm2SIoYkfg4UD7vXeXR5cxM56/FZbT0FFvQ3jsx
QTZMIsAow3FHA98N1DW3fqJ9PxZ5KpAv5HaOmZWWZClluraLRKfqEJ97+O2CPp5dBV/wJ7bUbu/A
xISSSFp7OOzgugvzOqzF4BIeH3csGiTOsR0rYsVX9zcM6jsYlkhMCvr31TStgIyC44hSagyf7Kg+
Jc6f5sFRppIP10grlD6y7X2od1BITCjYl822DZJHB4Fj81T/ppI3dGZ+voLM6McupefNw1Wcakoz
WQXCDf39wHBZSbGKftotZtsxctaMwwHyBoQUgE4bg76k0/ZI6fzsA1hEFKFnioiDmtVuLH/YD3C1
0AN9ZFvx/3/ZsQNM2Ru3eJqOOnFinjmotfhghT43fjhXI5fhFVySwbm//Z5v5BiYtgI5uZWUY6q8
DGW+1t3IwKyA5+lH0/2MNg8hCeAOSSUS7DmNu2hA2xcAUBD75wGHnH85J9JwNkgTl/g2mShjLwUp
W3HvKpnJNadbZOHVcbHRj//lRTd9VMvoc1u2ILKO+puHrjxs79wKHJvmcgHfdPZFhIy2hbnDniBh
m96abqR961Qv1Gckf2nrLi8APgATw0WJAIU/3i8jMbcEztpQDRCHXlOjXLJfhLnEY8KM69WclG2k
RNP/oj9ggQGfjnScMlZB9F4N60yNTHw2pEjVwAs4lEzN2EabVLtU60DT6kw5TkLOdAUcXKXgLc4C
t3tRB1jo00wxlHICEcbPy28K/MzxMDgwJ7/oqsXvFMnBVA2Dc2EMWeCVGVRfxliiYAOVSDeZqZLT
O7z8OyZW153mj3K7OqA8d5ym3k+F1OGHdvVkrQFoErPQgADiKtyVsCLOB3jkRpQIi9gPq1T7G2KW
YN+5hYPARjX7/mlVYGtMrzh5YA3se5tudjydk4w11C7dfjyCjd8XIjZb1lw4hMKA35B+sm4f9wbc
UsBiGDpuy42roOIU2qR+zWwUzjATKAywGfJ3vhA+KWv0xK6GjV4Y6QyeTMLMvt/lwRqmaSxsi/bk
YONXQUPMgZ+5wr3/9Zn8CKx6o9OC7e/HzbkNo1/Q4p4obomduBiTFdnc1X7RAg45F0q6sTjmKJ7E
BIrBRzrcM5Lc8/ar0yAYea1nt2nQkkRXBCHig+WX7zhNJOwXYq26uZVTJs77KM5EFzb3UkRwroWe
XEYXfbQxl5MIo7uAxnkR5IYys4eLXcPm3l0uEBakWlsEhL3VeRDUmYzI+P9JGOSo04xxKpKj/s7/
/clRy3nnQ7W2n6UXKV8SKheOn0YJSbIzWPrbFOrK9qhm9OS0gAD9SDGeDBAsSJsJC3Hxw5ZSjVKy
/Y1IW8IpLuz+jra22KfnKuq+D6mLWzkYoOL1dJ+bRufj/w5/UmBxpmIZU0o1tjXIdeAtMSOjVioT
Lp+d9ghby82ip+fpCd2eYmvw5KMNy26gX9OnI5U4BjBvFJiz/56F3Fo1TC256EEC8y/KTbsbCtdj
jtDxYLOvEOrUdlewpWcIbOm4yrJ+7LJA9lOvkJpqTFnAEtelCFULpWXXjbJ1Qe8CVSC6rGfbcSHf
rfTAq9m3UrysQ0PquubIxfxhH3pJY5huo9E/w4XYxVRyOLjAoRm7vOM+CWxy3Ne9GvawSaDS79sY
WZslosmAHZtvJSwSPli+0jHy7jMDnvKNABr59qWaEh76LmD2atYGbFPr1f7PP7xyd++mEgVtoCUc
F0+39jdiwoUetxmcg8Q7iMi4AkmHFZt7+Oy+mTN+bvTrYWrDFIKfSIXs1e344DKRGEb1OSE67/1l
89gqKnvVsPfnEOiuDzzk/j9J1jfTCTpx4UfRv8Uw92ZrQ8G1KogpZsRao1IoQNVfeGeFLEjgTOm6
WpInLADBkGdf7VwIn/pE/BOPKGi5mcfuTGWSKP7olKdl8vMtrUY9Ki/ptCFafFxWm/pGMfIR2IGp
AVPDgSAM7H15z7TrCxd6/pIAQSLB0lAuLoZEPJiOHThGsj9Sxsm9OFo6Ezvnl732BIPa/ah29YnL
1CrACy+lYp42WaQ2EmqjpHTYfb4z8gSeag4ORrX92OpOwjNcVLmBsifLSTFdTAcTR/hK/kTgGscc
FU07H5lSTSprMV6g1FJ2yt2INsgV5K0dU2FS1f/FdREdq9OaRVUTf2SLRAB6GlD/y8c/NOVBwiIf
eKLPS3LebpCAzTDdAvC4L+++vs6wvAkedzOBGgdDcVnRkxfbNnIEOU73M9iXFOlTxOjisE6iCFmm
/FJZgYFy0zWTGBsTvkc1Nf8pMwfds6vSDz6zVf+3pwBInOWuB2HjFzljnoJTWYhYAzIdXtSfZcFI
1XvWzWCik/NLPq1b3gY4wXgQjCFc7dAeXOFXbli42/T8+u1JNs+UfoKE6QDy6QNkLuHeXFaM+ENx
CjX7nOC5B/biy7KJOjiG5luFQid7KbijrR0mEfjfjfBiETva++6aRqt/Zs6GkzvC+voH+FuYKLCL
xGne/ZqmKK3S7dBd3b4tbuHlrSpGYFjwN3Zi+5hqBuohSoL+5gKCJ/lMfdtNBoUlQRd9o5LwB1di
nR8zKAe0zeJ7aC8WB9MqXxftpw11XLCpS2VwDDPkRLv7mBSxSrPDeYxPlylZWLfIiK503GlxhILS
b8lACeW7bWlPmsB/PHgYql3vGyzsFv7c1ZNZalZHcMdmXMCqv8pXxzkDdmlKhiE4rDZ6XP+c+h3r
2uffjnK4QRQDkNSY5xttfUt3qEb8fsoXWQtqWIww0wckP6MyWL3TLHKTayU7JIp8At1VkpGBDOdg
ju5RgUQd3K9edjvQ7fw+f7e5VHCQNTnF8J4rWpJw0d4YMIDpMnez+F+qkn+/9wW1HL9yL7mPQ++6
m+9JG65J5sDLjsWFkoCrOOMwnd5kg+IXY8biLXocupEkUf7yw+XRXg3CiQvKKoUxwLNOaYKNow5i
KzIWRK1sYixSDfy2x3AheFAqSNPvOKR1D1g8xze3GwltlrU6m0fmBYq2jtHDoQZfd0hf38GU38Gc
+iz+NojNfoREmBFmYK1eWtXYjD1+spmVLeM6uHUhcJbKkbE7K/9AcmgWDvi5wRrYf+HI4lAOPI+s
IjNfwQZPDZ4I/9EZ0MS6gVPo/xu+B6GpfNdayWB5i98k+fr0+BMzhvVWBltFk1YeETnm5Y6ed28M
uoB+OxmQB1AdaHJM6VnebaGala5znFOhI0PuttmTfRYxEiiFcj8sNvf1pHADath6uxVyLIEgc3Lw
+o6fFk3W+/UnLR7gwexKzMw1O3A2AHAVm/4iCSA3AbpoaI2by3Ceg1hEkknNlGahfHuJs4JfEK/P
xVel1EstL6y0Xi721WzvfNhVJxOCcQ1U7CYGvXYYDojBknA1GrebNwYgPYbyUN/xElbChnYVAcry
5jDR/BYlFvzMHkthqjPnGL0G72H6eS/wMQ/PDQRgBd+TfMCvwokdZZnld2/agT0G6RoZwhr97UBd
a+6pbDWgIKOLvu3KI+GMB8bxEcY7zfLFxcB0Dy4HMYYWsBvtjnLrgImxEV36kuukIWNB0sCPgLss
0G+1p+3hiwyjxfMhGewOSWKbGR0I2yORPpNE/Q53agvWM2wsJSyKKdS9lcDSkCgayHkne4fxeKY5
gCGh2/L16y4GhT/nVe76C6PFF67kSTk8V1Bjl3JDlzP5Jom17UYgjFsqdttB0onvEQRU0PsFYGDj
oZwez/MTPgetAllIL11kdpSAe/TLQfEQMQLLRezHe5gljGfCxkYqUuohzuwY6UVErKJzSlzN6SPX
3S7rpzdE/p3hRM5lttFYZG86V1YpiqaekVUSVCZ7aYvjQZR/09z0gOrUJRnwFzptzgrtvrOdMSCR
vjlZYN3+C6XMPlYlGDsTrtnyyXCBTujtSnWIy1ZwbkLE/Kurmq8AGYl4CNmPtINE6DI05qBFWAVA
BqN4izTPmpY/51XV+RCLJWPGOAfwbs9KlHAkEm3GWpSLaPQrri8RSUlfsI90EYxlm5canx2IlcUI
oq/Os2YPtpPdyS1qYnv8bmSIndY19vkFnRBa2v+x1btxooTuxZ+S5y4xDTlHmSCmpUHWkPlUv5kK
isLQ/5Vt5TaewSf4mx4g38PxeShcHaGt3yZ7SxoS+KcQ8PbY6UTh9fzWIgds2xxgJ6ZmWSRhiari
T1T0aXHaEIU9y1g+ubQPryIySRSF09QLXUGhFKGDt/x5S0bwmnzKCShTf6P/gF92R0E4x/ZYTDQp
0rHkAw1OA/FdfQ3usmWMM2SAohflYS6jZVsRxfWCZg51N3XzrB4LhDYlmeYaXAZ1fL5JMekapo7a
6/fONhX/G8JxSrl6xMHdMnQrbhd2Vwq41BUFqxvtLpEeT/Dl5jRZEcAqn4CBd9mlb7ebSh+zR0iB
uh+nYvceJk134X5oNPvs4NPVjOAdU9XSRAeC3kNxlgXkDyUt/CdlQshrM6fOnRjaPEsVnuG8b+Nq
n7cMXXT6Tvo1nU6wBgGz4ERI1DEIaMZl3dLQU6DMimEpWXnOXQqpV4kGNXO8FfxJSBkFPM6+EDbr
s61ZGLXP96hBlG/70ODQdGcUoYpYOlVgLAJ6m1eMWfE4H0qDzLGcqb+Ls5zwh/ANIUGU0hgTz2Xh
7NlM8zZR0/UOZyNqMXLPY/1DL5eExDpRcpfwXI6o7L7NOImgfRXrQoFvXch80HK9caLt73Abp8pZ
7SFd5uWDfc7eR3mTPRuasHjitLxCVI7zXwlkpMVHuDiJj96s/S84Rkk7D+GYpjrtbpAhUEZYBrhj
naBj9chNLqQ19iYQWErC/jXUeZCJt/TKKTzR0vUd+iEeF/yaZ4374Bl5rb/3pxCiFvrQ5cbLyeCd
GpmpWoe8US5SDxhaP0iaNIEqi18cqEu3lUTWARyOcIGc6wfrWZKbMhN6QQxUfBaw6Okb3YueRiiI
+qbwYS+fa99BOS9Q7FH+IOLee5wPXkJuA4a1SOpabh/aMmXwYulBlhY3FbBkeRk6czyviFI6BjO5
6fQ/0VjwHnt9qW3Sm7tvj7VJ/E7xZV/glFtQeOsx00uIycK06036hegC6lzJMEKy7FEppRTyMjmC
yuSX5izrfaDSUOEdXzIQgklCLoqtlTfVGUkeesbyTf53ydnmNypcGwu6KvTJM3uptP3AxcBPAQiI
CH9r6Frpugv2gqe9Hs/gQQfI2KNXVrawBNRShjOHUSX/ynaUzCYy2uJOufSBfbWZ65avW184O5c9
zeXSpXoDbssuOVAlvoXliuK9hQ+IvqvOlfHNCWwzluSsw5nu8S16hFX0e2hrocWrYXgaZ8qGoB3M
GQ8LmOa6jOshS+Yzzy8TfvAaOU3BmzZPN01ZmMaHHHkpQe13CS1kEGqAutm1Z/5LHifmREz2Y7ko
EMHmgF3cankzgZxhZpMSUZ4rmxyIBOdqUHjGr0nRzIYCqNkyJayDRfe5uXljiy+kG19xWym12UhX
CSgIoe0ChPUnrhDvGmGJPimUEB3Aa6Q/iNG/5HakV8L9ZWHS+LrnE+HYZi77tstHowRWFVZVQXAv
BAJByZP45xye0Y/mwFTQjqVbw7u/tm02xXC95Gi+Mu/bSihX9SuM090glf1ogwcWoGW4c3gXzs8Z
xT4Cjdvj3MpZhPmn9ymQ8wu5NPbzPxh0QLRxOOsKI06oJhCJy6TE3QbxtOf2/5cqrkr+L5/bNkDU
CF+hR86ExoaIK43nrAOwaCb/S756bwE5aUW7uNguW0mQqpV7/VSyfKuTbK7sNllZH8RT9zLd0PNF
pbmiNp/UlRYErETTMUrF8JnY+7mh441CDVlnowk52clzFtK4XOUZhYf1RxxMGD1e3rcCOzmUeNau
hjEtuneoy1grQvXCTyc9oa/BhxDeAlXowjrc7ApUtUJznu8Ouryqv+pwm3/24sJlfRkr0Uqfoids
XgquoGA+aFjCLPtt9yr+uRYLl8XHlh8ZFO+R7o7tiLH+RuGW46vktkVaCFM3buzoGaLd8f8uvKcV
ozBiRItJuUPkF9ynfoXL0QKHbwij2of83ag54TyMhnoWG6Gpv2g8QhWSIfrzPVRcTbcgl4TUP9JD
R6E52gyg6qrNvwfmqS//x82kXO6DYaP1MZvI8CwpVhuOuWjdBd4JPR2Jb2rk/fBUKl5iSV2tj7Ln
O4ZUsJaYtcG9Iv4WWygzBsVyOzl2aTewxT5kdMdCg3xcP1lYvpHrIYDfX2RgMbEdzjYlCoESfT4B
cvmdi21weOzFrq/eEGjjOphyXuTVbiFjFRBl28h6z7BZoANMpNBMAcVwVPHuQMAfB+DNQTrksjNT
PUaW54ZxQhQUxG2yrtMRA3vXZlyLbr3/FsGSp7JX4a2Qhg0PrB8Ba4d1oqtw9laJlc8g+D6tEfcR
IwVpz0BERnhla1J5Y4xkwIvReJp+moCDdYJ/+zJQJ71VAxwY5ZMMdbJOGtocUHhdxPguqNmWLIcd
70AI59ZAZzeIfB2ewZT9Wm2lGWHuY4QlsZ1QR4MPbW2/Yp4adygQcrNtu8t+MbdWHa5VDMb74ryD
wYg4B6umDEi2U3d/X5vXHjkxkKRDF1RT7inLoFRHdt/UVaD6D18kuGaCuuzMhfhLJJk+zo4ToE+d
KSnFwEgGCQXIXTozCFSPSHbDoH89w5YtESTyrcDyCvrIHrb5++i15ZxwoDIEMrpbBIJQRr4iqDzG
ffXH3AOoWbgEtD82Ve549SVucAc1SUXmOMpiYNMzQ/U35CoXrbyo/QxtI56xhC8ELIJPP63SHNOQ
7ee1yGJeqUTbXhOX00rf4UPPYbSAMQo7UgpL82lOrtDmM/Jk7ySwP27yCrqzKi7fH6jpFhMbQ0br
vZKHEN3NeYBBZsgWjPxCWYLMLKAM3dNAn2lBbyHBdUnTLfC+ltx15QW/CDYmiQRAr0wia2qaZxa9
MYHlWT+0g15wpg+WmyY37KJ7B0suK9TbjdlPNFu4LtbLjX78Ah/aOrPdRZAiPeGtu2ildNIGi8pv
/54BorSuYNrcQOxG6LteOkfO8Zvx145f4IBdAwVNq4czapssITUH9LWWhq88iEkJBw72aZOLclRu
dGlBU+J2k3nYRfbrXTML1uNO3qDtKqhwZLAHZRVa4iscnI4kbmE0jJV2EPVyAT4MW2aZB79IylKc
Dfp54KuPpac5xhs2mRKpIAc8Nt8Lnx3fW6LW5aBynDILtev19j5a5LVY/QDc8yBKQioENI6N9BUo
bd6pjwykS6cw1nzhwYL6Nj34QDfxWRQp/ASPxUDFzlB+wX17HjpirtzPEP73ZV0ytRi7n4o/757i
MMHKCcbYxmZLLRa03oZgxUgRHB5ssZs7fGUDMOwypeTMAAI+dzy5EM4ZkLcLYYCocCtOh+0SjC4+
pHi001VrPx6xi6AY3UHqnAuscmHEA+4Bnpc+3bbxb9kRuFb6gcFd0ruaaYRn1FsNOfAbvH5SmsV2
frTx9T9UIPv9kZsEhg6tjkSKerdsvmF2hmq9euWIcPLTPq/E8ICXvz7b7iOK1/emiXsi9ChVne1e
bRAHrgDP8E4EQDPk5mKvYes6ehaJ3soUYpW/dBznclkmLy92b9sV5cHVVCg35pI0Gig9f9rR+9H/
dRAJcG3zJWAQ0w5Oos5cK8qOSdP9Yp7rXfPRFA/yHITpfQKPsLLN5e7XzRM2R1LW1h9OEDNp47+S
k2ME3QUqoMXNeNCNXYRLQKU3EZtcvALQ1C+UHQ367l6hF4bZwFy/Wcp07JSudOY5woKxI48LCyGu
X6e2+jhb8OM+mCVWHBX5MptdL5aBAjritvryCDO2Y0XWWI5p6V6qzKPNpCCIgdi1zQ+16h6f1tiF
nBLDKAxUd0PucO9Aei9AYgpAjyXYwRorP2RqO6TLvEtnosBsrCwwDilReMCcidqNIakuTC6AxPZX
5PNjM39PJKMpHvfGCjMUJ1RpOUnDvnJiVZZPiRiPPHUHscxw+DmQt+8OjfLR4gHWzKyrephfGvmS
JYvu+jYToENWDomgx8DM39QOdLvHT0KJArcSKiJ7R1zAQPOXGk0ziZ3JfHmMAO5H0VIIRx+GS6bQ
2XSFqnvwu3SaCU9Aq2i98f60mr5pjeeasi341z59zS6+0bjXDDAN7ktlei2/aqFfVQtg90Z2udQh
fo2dBBzoAHqMbJiEAklTQSMTQuZjRpWtR2zi3ZnohPQdz+lxkoz5NlnAhGVgOLCexA7nfv5DrwB9
gWNwRAPkUu4y9/h5GeJ/E8ywByUqN9GJu+RB+1DFqeVMFnmafD/k2BqPmG6ni8MsYVmC+A8uzuW4
jeQ7+L4JCpf/ZT4kkRACxWvbTFvBzE+wLEJK8GBRNc14anLrXpGWeGCt3JsfGrzSyM03Rc6pq3uI
SsbxIZC2czb6qBJstOtDSbwLKI0CQgnZr7+BnH+62fWzUCID9wlccWoJwdB4r77dTOuRc0m8c2We
Ez62dK9BVzTlTbei8if6gsXxU/SV3eagpxKYfYSg3rZMn8TIpMjqMPqukFQ2Rqr5PE/LveawTLVI
ufIsN16qYzHHZRy6Zho3trAyWgQx/Ajc1ufFXQJtXiI1SY3z7kCvAd5PjXblo8WpIWJkp/3PseWr
lHowrGyoDTmfycanS9ouPHAGOgY0DaCfSdGCeCkgwhv+Wy2rY2zP5wTZiG/Ver7TQ1aZK9wG3Mth
kE2PVgmEjRwhUxTPQUBNrHrB+2UcRBNBGGyqxvgxJsEuZys7EVNB+ARe6STAOkJZbt6d6Y/6RPac
vPlWPyXtisUqLeaCHAC/uzYYQAwzzJzF2T92KbWUap7wvU5cmIvlnTLrbVeRgu192xQmi8qPFnKN
phGDADTzq+qCv5csYjHs6sR41EBYucfFqn/cSfk5xFxqDQjQa361TzHeP0B8eVk6hulYEBoNzGd4
ROtyiTCBwP0Ey6adAibCuXxqu7vylnKQMRk2v6zQlm8rlS+7bsTXSa5QwciUMPQVcIm5lnc4u93l
51BY+uJbiiONpIjWRr+o0FCGXpf+AKys42rsYfkn4WVsNm63finTunTL2ouEjaDkXp8ysf7isb/2
0ctLQtABxImJ8atjT7IQASkT09xbuiC3dnIxX36ruJs9ySgu3dKgcw1PMX3yvH4O0+PrMQJVWPtY
fOrOaLogljBqXERcBxBRgYsQcF6GhSvQ9Tm2WJmCmAU7JN+zRHVt0yG1y1Cvb9Dnvv2inWNzecCl
K2/MQomk626tJmMZalXkV3YjMuxttRF4RfhNoFYmK8tuhdK98XQ5Vw7hm0XrqN87xTdnR3p8hSfH
EheR1qzMLqIQKmJsVWAlj7pBVRxdul6bjaPMDDFntfe9jkwa6JqcptQug8hlFi6Do8veYbX8f2nn
t1gYsl9ZwuS5TdIPHiiBSrhtOg1puqKK30FIbvsgiD3JOap6ud6Iv6vGxY/pQA1P8pPXiqRv8j2d
vLhzRWPIwz32auQ0DMNe2byPcKZ4zVzIYVC+BhOakisYLb28UPBQVeaHZkWMTHpQr/qtShTr/REY
vE0/PwJr39tmqe6/PElKYgKSjIyz6eL8vMqZomBH70sg/YcZfvhAy99vT9pJ3/4tG4fWklIwvJEF
zHd6WbdwERbJdSFExshG5q3ZLiEZrIq6kz7pS7CUo0GKdzZif7PFM2JN4TWwrPtgq+OzqEL7i+F1
37kY3L5ViixeEbPuRFnoPWiK3fedBEvus4cTM4Dtor1rSHoWAF6OZtby0xhFUmGU2Hpod2DsubZY
rVnLGazefYHd3eqp4wSiyzkzjRI0AtocVHvNiJqV03oXFOvJFxNlMWAqJh6PY7FDP67OHN09S534
h9SI1xS14fk8/CI8Z1LHcwE45uJnOBJI2PjBsqf7HPV6siJVAmdOgOUTXowfsthqkcKaH6fkhPqJ
0jJSn3xEO3hEUAAb1nZ8brsrgxThZs+ETOuEwrd/VJjqlZU4Ny0znUdxoEWC161YsuWEy79Y/b7w
JEGkNOwd9oyLkN6OIrFmHKJFxdsrEP5yAri2SgLJdntsZOZfarBA6p8vyy9tNLcJLEEMfQlNADU5
JEYTMLaIYrEBSCt8wguj80/xb5ojFLeMu68qBGcpxZR0FVBwP9ozOYP2WejoF+OlNaikLf113jxk
zhvZ1Ok5y1fCvx1dz7wd0GU7+cRPNiccxs6cGHHFHL97iK4/4K1k31OVMAiddJKIRLhO4qPTSkVI
7V4J49XTYDtecVCWxQoOF1ZRnLilKw9xPv7fm3BgpKwdR8FqhZrd0fmW8CPBmzzkLMa5UKX7FKE2
Q+F8IwLVaPLAgVP4r4yHzcjsd2FPF5Xpxi3kgulyvz5zvI577OdJFR1GnM//T5DqWlxE2dTjjAU/
wGhBj2LOPgXsMw9jCwPJkjp2wZpElD3EWU7Pkve0sqZm0CMA2JJiS6Te7ClZlUOmTrJV/wUIJs/s
kVhLl+QWqEhqXNY/3UZRiP6jctPHVMIAqVWxfjmW0LDwr9/zampm0uq2Ls3NM9IFBtawMeRPtKtB
BEz72YPqG2VEJcWHCMH7ApOeSn2NRAz0UjInQDCkUod9OFuBaTHZZUC7fq3Wvsb5E6qkiriuHNaX
5GmOidOJ2dHO5Voguu8bKKShVoDH2OobQTsifp7HzosISePpI/WzGfJ13pBxYj1xQ8aYx8y1TWV7
OARre1WKdqRi4QH7YZgnRISbwW0kjK1dYXNGQYKzUoyfoOxLYSc0Cceq9ni/xDf34tFCuWpUl17Y
hWrj5EHRZw2Q9iqz+GhvjMcq0nfHkBT9EbS5u7nnyIH7f+/c0UP2twGeATDXOhsFPgA8jF9s41m5
8pxtmSh7jA6qfJqszff1XI25VDE5hPDMURZUdjMd0X002Se5Ra8ql3cF6voUIWnDGxlYQDkM04no
b3KhHyFmu5PzVx8z1Bi1QKnRBKaxr8XuqLPZadhGUKs+5lLn0iByzJVrXWs2Juga/lM472oAMUrb
nr9A0l7IUBJJZKE9ErYW9i681Vre5IifjBcu9nUWk2KMEtkE3DkTD0VdFSWpz4LbJNIqG4120nbR
pwZFi5HMrePuRoP7A9LLygkqHISggiK8kBPWrp7XVQCYN9zh0o5xsyWQHRH53xvg4qWLEhc9aWrm
uJuQmphcwwsLLTIb14VYPgflCEU4dg/Y/4BZLH6CVShyxTcor3gZHqItWWOcnZeCkxb7Z9SEopni
/q/OyCSREkY/CQn/SyCEdUj2p/k4+jee3ourm+8/7oqQSigQL+syuCH+GogxdkTgJUtKs0e+Vyds
91+TsP7SYN/4tX+cmWnra1j4GgwRTASz5a7p4z6YIGTL6fsZpaOe1gYzzYlsqBxFlCaeny1V/tfL
mxmFJv+9ZekjtMtdNR02EZFYCed8AluPrbIMzrEEg7IqsVyVXaVCxDtReofCABq5T1VETIn1Rydw
KgcPSG4WOI+x5W+W3K2FgbBE6C5zVNCkmo/8UHtDJ90jskIvEZUDrE9d6u0VaRQRzCH+E09f+wjr
nnqIZKSAYveqF0s8LvZjMVylKHFCUmd0UXosgIln44dBwON3BkdS//8mdzO7flF63uLZ61LecAL9
3NkUu0burKt+4UwV210UpBsdBm0+BzTnbhCUB/+lvjgZZi/TzK800v3fpCheUvY41OgZy8aucUXU
HCXJ4AGMk2TNKX0ZvsQC4qftBv/DLsrBCWLlsVXytkJ1vXv6SDRes6aQErH/uznOORi6q8RxfIL3
kkTiZKjnuBfw1Ti+Ouco/BbBmyzXvHssdJmu2vT50DTf9fZbVvRarT5dg6HGUcfv1CPhu/+BYGhf
ZAythwGQlVsQMgiQn5/BRygLqR5kNbhCnUHZAQlr9lI28yeGOr5khwY/dNWfb5c4aZ2+c84fwwNb
dddUS+YUaUNdsP7l0IkXqILBjpcL5+oS+FI70Gbep024qZ3PDf7EwKUwplWT7mG5+dJ5FXyvX9h/
wKzbMgU7/nOPIMTJ6stnSX2LvA0pEalN4ClFVuJw9ED1ZxXZr+J/wxp6E7w/j0ShYG/RbMANMyle
23LKwR/ZyHq4jMBAtcI4VPUZpEXC9BotSpsnCeBj3NK/S0gbg1uctb7Su84QyilxPuoDhRn1FbJ4
b5feILrxr2eR+gRWeSevgpFpHImXWGcaB5JjQsbREZQ2cEa/eeKKx0+iVLtD459qxUgIxEeOuvSk
6KwZUsVxxDNw+f4CrzPwXL5OKI1gWG6wkoGCi3fOcwnr95t07iPp8YSSPzhIfBZCXtRDhM5+ujSo
IYJFQmsLTHf+RUCn4WM0INPFIqWyPtQD3Z+STOhEVp7j+V01yGuqcHi/Kd/0P5NrRvPiEVNeueKp
Oj2EIxp59BYyJ8EvnQjGr1bx9AbJWWNJqBvnLdefSr8HxF0tPOnP4hYi/R9rFUY0YR3DOUr0/fPR
44zU8+bTns5Nr1ZO6UTEBEc5XVAtyvkQBbcHqpNXCMHXxamROInhIjdUMmhYRsMNeV3GElFwfbly
Z+/Tn0bG7x69YDKggeGCHr6xPcEmLtGL5fJobm/6S49YHKb3u/qjpyxMimbrkQ6VSkw1H1CR8TOq
pazLB5FMqb1UEb49YTLna7bh4Lawa68FwfZWrduphFPf5n2WzcVOslmX+h4C67CK6PVjRQE3jade
M5zDPP+08o/uoog3utu1V3RyrAnZkX2ZrIjbdj+No6i6xO8orn7EypQ6Z/gZm4JML3JT/9gBqgPe
fanTmn8zTsfnA0eglJJo7kXNgFWvXi/6jF1nv9bT8thzH5S2n6r6H0MSijzBZQMh/NgWLpcK8ST3
2JZuddrPywMWV1d3T2T+/Uk/b1DcWxdQ8z9R1mB/jLY6bTHOMgHhIseCsk0VbnncjQZvqm7kAZTr
fHelNp6I3hW81/S9FSrJWKtPiURGXNev4PCvBhpdlt4e13kfKn1fGS6EWgrC1LYSPQJsGZ+2gOHE
0IqGyQ1j5WSaCdM8yAE5HQk+AX0jaN9XfCT+Wt7pwaa7gcuujPBe0hniGY2V9WGgDUTIUXe7A3NT
OIGfFcYsQFUgcFgWzldr4b+6s8oCZD7fDfhAV++jvbK8asl1jd9p/pwYt/CzT6mGGQr+Bc0vNgE0
dyUH3dp18Xob1gLw/mxmdONCUNwJwwVtMtrE0LOgXOYQhAm5FiTsZcwn2KfbLh4EpBN6Hccz05Nu
LNryAwIypA9xleZd0iq3tZbhYuRiDgwHxJkXISpq/beevorpgvKNOXqTb5ZwXD/LDvletkfbDK3V
4mkaM7yUKwMtqwW60qYUqTWsejwZQOItIE0ies43NTX1WdpPE+u9FFV54U1aYcg/orPO0OBJOyES
HNfQNpb5PZqzuwbFzSBdQP8nmWG50TvEU3qB3BZxs914qAKMXm/TwnMgh2Ne8+vTfVkTP0uky5jT
cR+HI5mUSObxxFF2MtpDR6fKbwADfdqVlDelme+kBZmLvWX05sV5laWapDFLI8Wo8J0l5nZjs9Uw
EDqaKX2KJXpAOfjVHJA1rwiQKEM/bnEGtps5wAZ3hJzWdd+xWQDlF8Cy9ALmuXWS7WHR2x8aWfHn
KTmQPH84hmExPWXAGCnyPc4f4nHV90UyldMvINBIk+hHNglajjrkVWRw4NNQ906paB1SBUr4PioN
lY2ZGC5wmh17t4m85FXUZ9cGYAG9xzdZOuMZs5G3UeuL2nRuOxf3UWGvGIDzJFnwSK9eAp+DRSQW
hvvFBsqdDQEBaAcUGOHmku+hJFbF60rm73WhvcYJ1ZVPPxiCWmH9rkPuOxESZ/sjqctgFjWHY5XQ
54aLGkQC/Tsu4nbW+NMJbpzhj+SjBVFt55UNX/LCsDcZp7jL6lBBs2/4eK0p15mP8Fid6x7eM96k
HnL3XfWCwRL2KYlYm5l/YhEWwWQyll943KyJPn6PWg5nURMnsWoaX511t0OZOX8gc2UN+g+neMT4
dzzeOFOz0Fdu78Nmvd7CmqHBiTbJ3N336/2SqbLhGh/H3cItOSInriw0OJBmbJrpDSs5gydqjHW3
iMZ+WFnSwLu8OWWAF+CdPn+vk5P7il96RViw9xZH8Mv0o/D9zFToMVew/TwptBMqLsvgsRv+2Jzs
7nYAbarUjgg0t7vG0wo02oMWnx3CfR/+2h7hA5gFMaHL0bYkzQXSmGtPzOEEA8Di2txJcaI0LKjT
Suxcehy6kUhwNpk2btM1R+PVfHL7DZudXRynSWQXtIlY8dfKIjBVfyYNgjlfaLduzGC/t0cKv7j2
wovTN4XRdNXV8hAyI8RE6w/Li4zUjPoMxDt3m4yS94gkEQxRXcyg6BHAIdrJWRDZ7Qs6jmyFNxIg
TJsCZg1bEpAKOGXgsxTn8I4RJa6PTBVfa6u+wD0t5hSLBQzYTQ4pUJ+k2iYzRAo9t5B+2eQ8yvzq
91ZHXW4MCxomaen+cn4UwDOQUcSp5iMLUFPPC6yENoq1iZX3/B6k/pZCc0TCxGhCykDjYZwHqK64
iKI9c8Fy0dY+J5gh/7Aw/T9j6FQTrjnafIXIASYjYm9LIXtgnHN0w8vt7DAGFzP679f7kqpZiRo7
MVPAyLJamAnS1LwabetAD67vmcFjpVWOKnTPXCYGMGTJicxNaGCPc+/plRo+Jfr0cyId1aV522uo
G0WAuLE442T3EUEq13ckMvT6kc56vmNh39pEfEEIzfTUckzmx5+KIi0pcll9qNQCG0yYnBF9PqDL
Uz8/PAcl4Ky3GsynTCQ70AL1zYsqjrvq6koubqMi2rz2QPoNWhzd68nw1UtuH6DpJjGsbT+HkhOG
JEc2g/2FUK1Uz6XYbpyxj55wyeTxJRQpVsWpi80NYd91vj1vlM1jLXupUIMCxkppuzBzitlYdmF6
kf5z9bctJf9HAecjtPSRSqs9Uq0r2++YVP0Qh9hnPSsWy0FoWHdRO++tBpyCFgGkPFMgntYYa/wh
QzMOfbazW1nPCknZ2TnaXNJRxcFRMq1qnPNxAm1cNSlnXQRTwwt/anUeVrYNo9O6aGTUMVIgIQOV
qJOXaJcuG/NBD0HL0UivC+MWoRwl9U/5e6jGIvPRDc+DHHTJ0MFghtbqen4FlTc0h3NVtYA68TFY
PlPuSJIT08Altt89RyZPtuNw2iVp/mfWcDEIK9ikJcEWxZP7XeC5piovWz0uoj2xfPlqr9mFssdi
UxX7Ck1p/r71JQLLZyXDP/QdL0G/uoSOI6s6ixhi2mPS4IbjB7kGSx/UelrJwuhdEwi0XiTo/RZQ
QxyAbwwBr1I6wssdNnvyfKFDvOqU3HrVPEp+EkjGJnrDXpnAzn+f2SF65T9rEYcDEqxweMySuoqx
Tpm6s08n3rlX62O3x93eZ8gxWWeKKDZ7b6bo9UWpq7YWfHHbzh/ub07ApMUhPBtdPVTOVnN2J5mY
JCIymMWJgGcu0eRQNzczoFr/GlaVK8evwZ/MZwADEKVWx9uWgDsA3Vwh6+AvO0Vu400KX4uW6uuD
sjFeoKSG4G+t07pl0BEQ+Y7BgIBll4e6mQHT8G62++L0MuQvm4XLEihvt0bvdm5G5a/ky9ws30ia
/IcXqTzbPmiyFtK9N99R+ygQjm/xFm/fU+Nih9iu4txBhDnIH0/27/MkcBRzE34ouDY7FzG/566Q
+VOF7Yq92yGlbfnOLdnlFmQEIWzI+4VJPSN5U+VryFg5F9CgHCuXu2j82G0RduZEovIXPWSpmz64
kWvsb9tJu5y40nWjAybDSfgMRTFFzVmraCd15ZNXXyD8D17m8A/B6eVwpTaLHfkSe2D2dUWZUbtg
tnhDlu8Qc7/CvvkInd8LiJepo0/msVdyKhe6egOy/AKvUh4SzkFPpdaoAtpsrcVAbdcVBLNO8Y4e
x+60VRyciqwT032Qhw8pC8hWX/4dgwk54ECxToRwMYFCA0kaMj1p/j73sq1TjI+8WhG6UC+kg64j
lvQEhydkRkgSaiIqOMwsww0oXi9Tq+Wt2ASxetVGU+klAKKfoJYirDODikDdubcGm/ob2Li1FXLZ
deFvuXeom55/GvnDlOePI8M/qq3kfD/oicRR3UoeB10yl5J/Pfd3vrWISlEq5v0hzC1fEFwsWW2x
fid3qAkkJQSud42DZ7fiFOBw1HHUp76BA7Yehl/aEtoJ5qLo0F4PzmW9J+WXjysPJ1Wob2mrzfwN
xaVfRc4UXvelkgJuaRcwCMgGuqpXiaswbdKxiGzQwLipV79+wodTIJsSE6s7sInAQ4DZqBKJnSLO
QodWtZsmc5IN2rL+ZnPE2g8htX58HY2TBswacmGcGX9Xb2SVu1mfjfPHHXaVIicnrDJWrWkmTxaX
FuZfLKavlbNS+h/8XQzRuYf+VMmUHjGYt8bsprvHzPs66J/gPilhFTFEX9GKfoSROZTCmdsUmgAY
CEsMxhgi3jniLoxWiF2zhYGy3Y4FEjuUEe+2805x7vto6GRZctQruXJKGQzExfp1t/Ybs0AZ48qi
kYC36Kv81DV97CYjOt9ljKzLUQny113vTrucu1a4no25UEr448gceDWg3lpcR/Nejz+bNRrLfPb7
LtSg3/PBhdW4jLT4YROG8OSLRA1Auiuqi54PsrnXqd9rvq0GyO6u/oH/PlpPFs4dpUxKRabVQUtK
f+IsvSqHzc6UrdMrbuqXcLZdvr1L3DObM78BlauiC8rIddf3+9wspX1txEEr3EkJvJ6C505RuBNN
/IXkrOccFK4hHD3BPNUfdKq3JA8luT3RoJsHo4E8+i5Q3BStpYO54V56V6NJloAU1u9Yva3/1dH/
UMKVhy/gOquT3PE6GLghALZM5p/BSGHXBvKMxMgOh/uTi0qbvtnHLdLKJNXmrCSuxahnehEK/vjG
hqpBcJCLaGJslQW+N9zZsfX+V6qvcrW4X9CHVnDuJRak+T4FcAoTDAkUV8bZfvdbo4AWlOQzNehD
ZQpIg/Ty4XLJ/uZfWw5lWB8ijtFrgMkIoueXSMxF/8cbZvSRqTZhmzwAM6JYCFRlZIpd2n9utP/o
Dmi4WLaiYe32F9UO06Tf3XqbNZ5yOvw/wl2o0OudxXcMjQRw0sgwRE6VX8fu3UnkbRIBzfK6sce6
Lu4pcV9BNs0LbPoGhMHToUf/1Og63Qr3w/AKdKm3aQ5VrYqouVN/kgG5TIRSsFUEckbyZwGtRoLJ
9mpOa1oohQNDIKgPAlbqPr66fs1f85+U9nw7yYfXSszLFgey/Yv+Pde2L0DNqTqe6tycrbDgGJdK
M3MP/6kZiQgQxFGDu6MmUFZKHq/X+cK8mvuQ+wi91IzVsldywBjtBxxiZf2fanDRXogN2q47SuNh
araUNKCm/RMgjWAdSTw/61G3j+1WG7TyefI7SV+/TRSnshBtUb5zUldOnrBLdW/9H8uUN5GyP+74
JeqSZ8zhyroqmfLZr8WyzGUSVgzzHj4EUCGoAvf8dGlPSiWkc874ebCSfg2buPc1BJW9Qb8aXCU9
tRMv+2hDFVDxBs+uXVhnQoIlRoCtJbJ8VBKiFiK2pbZDfZUbfqS5Xr7XJ+CKab1FfsoFI3KSiYSn
JSOKCG4SkDVWndYaeWg90hu4+jAmttlerNxCw3msqqusWYpMNZPb/q55LcVv8gbDibnJKg1TL2SH
9gxv36wq7G6WicQ9D8gmbwp1wFA1xa1W/Qyj3rUfZV0CjNfb+WC3+dpuidWfGSpUgYMHr+5om1qs
1SDQw5/om/bCzQcEE6OTPyoMcBvq9BmTu1lLeRoafNDK5YsIakaE969HwYUNEegzGoqxCZvdSzRx
13HqfeRtIsjPXA98nhAsCiZveK7kA9JH9OjRBdI1Hh6g/SuDMy0/a8ysyNGKW3b0lnYDwvO5xTBu
j1Ag5pxk5f+XId5CObqE1gLXf39kRI8aHAQmzol9rHuvvqyTg06VIn4UZPkZuIrIoIJlWjwkLvgU
CAO6PjZOlbLBhNpPqIU6V7bt0/FCLbqhX1X6YhC9AQeB1g56oQEE1UW0duMt5rlsxFXehxtaS0bq
ldx9YGPFtwYVOAHmrMNFzbyhfLEapYKiDXMOCn3LUJQBeHZOZKRHTXIQxOC1xAqyYhGvAMa6WgKs
SsKxVBsXtu0GpOVuxJF9eLSNGLKtEqvYkR2Vd+0Z0pE3SVq3ltpnncOlJBovam3niYmICh+Ti+9Z
Rp8d9G5f0r3+H15UXLweoYAYYSJWeYEu6toRRqYuYu0v0KNVSvcI/clvnuy1tOc3PJ2BYG1KpwJt
iw5GaAsTouWe0dVOSlHrf9Yx0+fCWqkL1zckQM2QsIr+b7Fj7S0mCF0QYz5GXRlvXjUG2yvwYfed
o5b8CQoh4mD4gsc9J34M8gbJXNr4HsS/TXq71pQUX8G834SVY8Ly4HUbm5Ir1Q4LNMOzR0mdHYFM
RFhoNa3N9QdUZvt6WiVGDPTQOjQYqQoiVSc+PwyjiU1570zfGcVj1CBJcqIMF4W9itnFZxlPrA5L
HSMFLiGa0guLFWFX5lMuL6TcEGi3cJEv9P3TdrcUzxk9f+0xXYwHkFm3hkfAoYwmGsMJ7IwA7AzP
woyW868VcbRXICo5iyDITA0UaARSHS4adrzQsO8P6ob5FiwFeQwGiq3wQiFA0N/kSDRVpM6J5887
AJJx2R3h37CNRswzYu6Wxns9pIwb8asMUkg/eP5yfYgzuoJW/FQUlbQshb+41NkM1OM7eeG0idoP
j4hGw3scr1XNeqUKbETpwJc0MFYIF/NTgihIX0aLty9v9iR8incX7hA1d6geDL44ofEGFdu+OUwh
H+wG9ckXFHmd7/FNiTUdULsZ4hu9Fzc6hc3b/EnE01Chv+RR6CCYNJQTfM/ethg43lU9u7ajfwBd
Qv8eV7y/v5QK/f/q5JfkrLGgIKpwVSkf6r9YvF2Ulsd54yElzt7UKoJZvg6Rf5ZdJHVfr86QPqYo
ojaguuXrRl9qyr6MP+yq59PB73Yl6UHP/gBzruJNkhhIrYFCpIFb5+9WLYGpiJk7n4hJFsx0k5Gb
dwb77PYVgJCmw+7ehBDcqe6TorI/lYUkCBLnPZr7ITKfcshzm19gc0fF637ta7hGoYvI1CraOVMB
HxD7Rh6jvy2+XH3X/lCNMokhQPe2zbjXF8hnKvEJ4kBxq/iKQi3KFwrZLMcaLo8OzzafW0Or3ohy
5D/ctv5AC7FWHNTIyzj/74pra8l+zC9f0hlPhY8AlVuGBRiZ65FFQ9YfPHMaUjhZ1v1HCmNPSQI5
XhmpJOKdTBIrFX/9ePuMumPaFSTbd4bNbfGAf6nAwNavIfiTmavc62ycbMgHpGNR7B2jotccPPq8
FHhlBA4ai9X2zoARW2oKKFwI0sWm2iYE4wZt9SdyeLWMifuE8NiACpLuvl95odh5v3TYJ79cdAhE
L+7AlYCqYm9mten8JBi6WIN/f3JCbbFcpqS0Xm4duz+r254AIzGfO4lucicwY9oOvIvyIppPTNeQ
1CozTzIYK4ZMWI3dE1i0iTLzula9EzqkaAsHlk2dMLQenRNYXui0WpIEzAg9xAK5ZzvfhZVgEUad
pI2DRlcj0XHMwd5aICTYuLAXF/tWGplL3qGitXjm94lazBMBtOXsuPzRZWRgx5iVk61kR21d4km1
CkaOhSskcJ27EdnjLLC9GgTaxVn1q+5U4438Z8iUyi+YD2iBV/+i8d8a3Ehfa6w8OZ9ENUrjMl3K
FlOYRaCQKgOM25T3eXzAyD8t8f9upd86+ZeDI5Fxlys/R3hl3F2eXMAzOIAUUL5jSF1rAp2bIS+f
P3wT8rE/qgi7X8NicNWwM6oubSeZF4Z3pfV9LVv2wCjFro1WR8rVm3sMJoxZdWf+JGxubUjCXlnJ
jpF5xqzytKRG6lfNoSDvZG++052x1SwwGEKR/DUXWZWN6XX4K3g6L6s1Yap8/q97EHa2QtH5aLnn
REUjN2DZsq4Rkmeh5v3GYRBVvijzMmOJLdBiKow1qXJz9nNsFMjWCFm1TfwB9v43NkpBPee9Ym8Q
pxgoQqAJbiopwpyKZtE+2knrZvFKLXmKuH4oZXhs6oI6cE1AngqZx75rPJxIAy0nlCG6QqGKqTeN
iFjadpij8GHx+nsWyptTaHO6/pg5rwWpVxWqjTyW2N2p+9QyY1gplOINY3imOp5LCNsmdoG4XRUr
UsUomE8QOZl/bIK4JC9jCPjbNrzDu0RK6LSrSu5l2K+W9HA0o63iKVhTrkyLOtD+h6tZ9oGmiZmg
lN7amW/PAYpF7b54PHOU4ZK2CdIPSDjOsm60NhppxBKPCNF+ooa7PG9w9oPmTGN2g+r8+eqNT4aT
H0oifchKk0aGeqdppVVMnX+tZfUKI5MafYX+8S1tE705EBHfOa7ncEEHQ+kCJhEXO6MKSRbrRQWS
DESC92Dor9pjTLgRGzJdtHJ85Qtoo181egBx8GCQsWVPxLoAVra4CSThVO046kalEdwnH/1SN6SG
Gri+jH7Fyguti/jlL0hQBmMLn5OOLD97iqxGM21r42fS7ONNIcTKPF5ZtCAeJzdvxOX7Yk2x57gm
pXjk6/MZU0R7x8ESZIozFHa9uDW2yuyZBEsXijQovtTmcipRls2E8b3FCc+xFaN0PtQZT1ESp4sg
4VZ7z/2k6Hy659zI4i5wzP9V0S7ZP/x4xFNQhJakMZRJ51UclzEfAI/LO+o9tzvxIY0s0seMTJ/W
KyzdQHHinVJlfrPp97sOYeKVFvsV17tBn6a1bjCio2GZEQVZrIowGuPHmX9vZi7eQGyQwmB8SmRW
nexPXs6qtbPZyVG5thbPO0r4WITBYdXtGLQ92X4kSL/IAaDH+/IyJ4nrshVhXwXCjh/Ejv010RGc
FO8zwtnqvD1/eM2PPc5+YQBW+JA9qFwABfW/SHxyqkwTXfevnKrO/ZtWL4zKUzZGRWAcXVyEYUJs
e6OMZGU8PfRtkqXNj8mHze4OjEqZOoGIejAiPJ0hexM2J/05x45QXeNdfStFdw9LTfSBFbfG3cF7
9aqAvF2HS5yffvCWa5A6ZI7+XQ3btWXDGrLmcLUCSpUNDuyjBSG+MxWi+ly8+Oe3RiDDyWe8gPUg
Yu9crPiCmk5tro0oPBnmEeVg3mR7t+c5Bh7ltjRAyLSEfKXifwWl3kWvHXGgEsoyYO3Haf+Ptg0z
rcB/tDTD/nZAa59gPGiABh41AxZgVpjgVNTOipKjjHKdFR9+MFgKeNvUtya9eI2Z1qN3fWvHSpXu
0BMHcDaGJjAGtObXPHZBDlUge/gtevOQLd7l8qNA4HkRojd6on+on9ra5w0T6TN6cgZgsmBJm+tU
JlByQCO8sYGNHSexL3waxTkl7/PKCvboh0ehA3Totl48v9p/H7JVrPG+wL4NFCMJhftC+8Uxk3Hz
Up8e2xr5T+pseddN7G01R5ivrAvkBelRwVERiQ4lrvUXkfwgGtSgYpXO9rmniPVca18+xPT6QzmU
7umgW5HrT8PTXvaBVEkgXkEYCK4xednWjPRJaK85J1ohu4TZ2oe1c9M0K/8vZ5NBOcFnMoV7FuUp
WSnNUOUS61plBnf//9ek/9JYY4+3kZO9AW3VfUIAyg4rdndl1VDrzepRBXzYBT4+8keX8c5tBn/1
NQ14+1lv5qn4yJ9QeS7B7EtvGBA5Hmy0sLtjnk+BvyEcuJw3smTZdSkvtnTWUFrvahw/mp/xOKxL
XTy4R4Rb9KbnhFBt8UGYB/ZquSrtDoNiEAKIlZSNtAsm6VFl4M6J+TILCrVkHpKegylUFatsUpfb
4UcNI0kLpCs+DBWRMctPHV4ltKRrRffErbBKz99JmGa+65pjp8Lj8HSofzpSiBRnv+p/3bilOSWX
2oHVVOGzpd8yQ57wGjDroJb0hjDhZJNRq6mlYsSLzaDXpJqtzNH7WMh/cc8N2Bfz559lhERSCBfM
CX1XblaXDhujJwuhSq5oDQe1oWtqbw30knlFv8Lzvcu/lofhAqqzL9jh2toBHNmkGjrsvMtolWdP
BWz6HYIO0gXaBxMlMB5B0xl0Y75LvjfvunqHTftfYP3NE3j8Ku4o0taN5QIblkkKP8MQ9619m+UY
fD3xfWlIcshlHge12b29+IviGmnMnsO0JemWmtpo2mHEGGTeH6vXiAGCdk3ZH1bFDqgwBxEiWQzl
K4unGftL4vWzZYhKJjhHn3zbi8tYp70AaP4ob6RCHxRGbO2Xr/5Kl6EK94JhhhNxu/0E4tvPfBxl
gb5Fj3GpHP8NEczaMVzZ+1gpVsgAQ4w6QalwI0w6RIFtAcc2ijFxqP7t55n2QXjZh/uR/StQFAtu
xEyRDhfaLX2CIoCJgYcyKH7eQiZ4Ou75pkI/NDqcupqcSaDxD23zxERES9l8I7xx8KTrvYko9m45
J7cdzCtDRt3vwvwTruiagQBl3EPuj6Wx8teqVgBjMSFLG947IZXnTb04WADLPlLWOH8Y3Hj6YB4v
Iy/ye+6WVV78IXTdGrv+DOBR0kUwL58xqlToQBbbm28431ZZYjXxO9eDKdxfYhrYQonzkI5gRiNX
v7uhM99QPf+7q8iB4xzjho7upZrP80xlD0XPDiyYauyvzJfIOqDcioWDvYvzKLCsRKgZ97CZWLDL
u7cHML2rbNBuCim43Ey2DlPQqkKebYx7uSsNuJWH/TvAZ3xRm8bXWS/p3293nqtxm/0d2bohCl3G
LIVRGAtO15Na4QswQHzyeJgbY47TtrWiW0VopQFqQLq2GMLAsAW0sZcaYEEBRDlFXGzBVYyY6+Jv
PEdEPnffpD/myxdcDnpQ+Q0HrQ8SCAdvNEln1mW3FW+7oTAaV7EByQ+U8B7sygfyCH3nVDXSGfax
zluGxtbeVZ/QmOFGOp318ljmIcOdAVCkNV4Ux3yT3FALsXQgZ9isuMyY+rT2dDfrUFaGMk5VtkzZ
DSxMkhzamuL9NVSHzUXHf7S9+VICWlSg4hRUzDQi02+9CNZF4FMBSG//4yjXi4UVGmy8n0WjXb7C
VODJwaeNjlrOhZrkmnJKLwuy9uxiRK4c1o0GuEE7PiPblIDA81cjAA8/UI1WgM4WnVzsyPHRQm7k
K+HfcX3cBzixYO2mB3GzRzwhElYtE0liFFXVAE95bXVjVGne733bT0auyo9wkhreXekGD8sqDlYZ
h9GH1aoZ6CaEmlMECk8rAmfuUkjSg/+rAD7qtRgAkvWHsOjGjjeFrpsBCTsOZUYWjJFrN8hC07yS
hVgO4tP3iWlHQbGX52EJW9Rr/oKK2XS+feWNF6BUfPON7iGSV/PCr1HJF7r5ijIeN2f57wqdd4KA
U4fvabftt18zGou931/n8NitSBIWHLBs4VTd6ivgfclGobWwZ1efCE/TeBqNyHvfu+1z+El8vZOk
QsRwd5SvGXvvlQ5E2miFxUAlS73sbO+VzC3QScfP1au7rjCnxD4anmay+GY+Zwq7/ujABQfu6AwZ
0uyPK89Cakk44lifohLmEZ3Kn9tlsYRI47emn0Pe6mMTygKWN6WL5eFM0K3PauLEE+lE0kT4f2B9
kSj7xVwr5SMuN9yws11OK292Gz7NP1TVe3W1FBGiW3X7kfATJuuCoRwbNGTpreJfvY/Da2Kl1qK5
Wzhv4AJmUGCg4AH0QlWRwuSRbC7PrYHMtwmn3IACrF2FM0v8qZwLDAFIaBJNnb5kckMrBKNZ0/j+
PjQIRRJwdkXYiH3MSvmSsi/X1vwtv3HUX9Pf8Lz+M7hA725FoLGupsOdBdFm4FMl7lHXrGO6CP3h
kMSCNC71UR3RBPBqm88zuXYa0+F9nbNouowuTtLf2fKHsloMbqBsuYfHydud2n5GaGbBO33epKA8
nWHGM8XLZqxpUAHxG2HJOHcbVM1NN4sDb9rYu3xBEYzMd+5vffIGUdKlvJP7+90iegXJP+Rr4rP+
VcFFLf34Ek5mEyxRpmQL9RChMO9RxTXUF1fM0f7D1lOCamWqnWmj4ThanwiEm6pvRxrquVQiLPTU
t65iDJWESCb3FFddnfVGjObb4x6iYXjTOWTcXT4OUGBRZbQSPRbMyZeBihowl8ZW4nHYblW4EfY7
oEaaItypiWuHuXfkmp144l4S39ow9YN5ZPuS6jTSNG0PwTL+Ak9EyX4wn0+SNQoNbp0StS8Ata8n
qD0Nq26Aum4SrpBWdGAXmD/ioJ/dRCx68kJfqHHSxGCr2HqadXCCNF87hTA6Wnci3IB7K0zZ9paB
XDrYcCwkPVv0ZgxVCgAHzR3dyQdOr6wf2WYMUruwSQP2HjQ8wSQ4SreiOHmhvVHVqsYgxHmayg3g
w3dKiOIP/Z2KCVYDMAnUDU/RN6FZL5gdIh1dAiEGQHtukO0pMlvreCv1kJqtbpRN7BdpmiC4lSB8
UfB03sNzW1nqN6RvDQArrnxDerF0+4g0+7CKTejk8uC/BQxdVZV+9ePenwoSELHSyQFAzMq+RWIn
flBERlsfwlU/Bl6b7iMeZiuPZoL1O0rrHQXuT+EZlYMbkU9D/1qFSR/hw+I2k2hl8UJeDaNHS7NG
sPWUMH7tcpBEANeBMRuMRuy+rnMwHdPqTBCYZ89f0bQGg0JcbwV6+DkQ7/fC59KbnDBXVmFy8r96
Y/Pmq0X6IzyZS/KbpXf6r8GvqZnyPhqtj6H/I9BYkwwUbjtORbcf/6jZEj2FEhi19nP/8T07H0DB
YjnGSxjXVRDEgGd7HkRiKZIUvuvApInoHZmtIV36DQtMxemhRwezpMBesZnAWPED4EmUBC13gMAI
oGz0qLSr9iGOMRSkPHY1MGmHtPa20a5oMky7JCB9y6BVj8BxN1TGp+fPN2wEUtGCuVtmCSRrFo/L
zK3luxtRJsJbqwAs2ftKTijM6FHidHVh120tKvoTrnYrx5bt6pAbiT7elrwQqx6hVGwTlG88QdCI
OE45W7fHOdcoPRmQhCWhyZW/L6wBiGPwSGgsUZK8Og4VwPWl/YmA159r7w6DqN95PTztpjA3Ykmw
thMZ/kZ7tSNOcDzKDUGP/ml55V7T4QYo8VlpHXdGsAwZDVTwnb7Ml+4Z+JS6oPk5m0ifGlqDBHW9
Rf4AYMibId56Z5/bxNgk9u3l2XhkxPnDOM8Nul35rjvefzaeZlXD71DOJ43j9YISxPxfOHiNoqIx
oJDxi6C9tL+iuJMaVKddzKCkbm+ZrTRRKP/pKbxuwyX579RqFuPy7ubBGaTgekHfU0nJAt5sRo9N
EX184P86uMqx3CciVZyxoQhEF+OlxDLxnKAnX6YizH8mupXEDFtC7Sonasmp+qIXiT52UAW7fxjP
mTpWlhw0FcGJyP9RpIoapnaaKNx0m0cuq30w/QsDwDEg8L0GWL2uhw0We5BQ/yfBmH5LAcCnunZA
gwsS0UuRQ8vJhJJI9hDP2hxE2f3Oji3vkZM8TY0QijZXkZVMOJZRmt0SNrEZICojGBciFeKwUVVX
RzR04UKtYku80pu8WsKb1z0ITKhAotRL+6IURg3c3pz9ejhxBlOe3xRskfkkc2yeJEZFM/DcMvY1
GUydPFvcUyplvGoRFnmBhJ+AO4ZWEgdTZui7UCgcg9FkU+bg2Sg7VE4WYZQqkezha2iFBDVQZ9Sz
qv5fscjO1l9DmkKFTW+LWFMNUdKiQ0qDRPiQ6CPSxH3jkK5mj/MlhHqMUMShJ1TT0+ezxXF4TnrX
T1zejClhIDzuxX8jf/zEuB5PaXDCePdj0cuAs2jMABDt4nVHrTmWkaoGEBO70mPhZwjXXhxp84n5
IKMJKyDgYCC/zmmBmY/GeJz4c/YVJP7A/yFNkl4j5ybTdBgCEhD3rmpVYGsN0fLrcUgBJQ3ickHG
ZbSkjuXf+2CQ3MDbaKvNJ9ZHdu72uHMnT4QDRkwDo4amDKbSniSHumKSDiGEMHpipgm6MFrPMyNX
OkL2RlbdGohZoeY9Sl1qUMLb2XJx2cKqVMyLs41vc33JWeM9iLKsBYHsZgkbS/MRSX8s4CTwpdQV
NwRuCE3wrg+10jzZsYviZ7v7nj0RE+bSdIXO93+6ZhyKsmp7u94/9BdfZ4LOPfEuiKvLDC+xAKJz
DIISm+Fncf0kR3hlFObbolM6uQZu4qGF3VCiA+W2Fc708j2n84qTCixkJm0MFe3xAzWaHE/BDQIA
1xDp/2FssAmDHa2CgdGK8pH7L7G/dvsTCKAAbbXFjDFlJ7CHtDzAOKpFAVEbwNJIELyeNnGoEklu
ltvPTE4XiqI/Tvs51B+KJnXFJGyDvGkOXxJP4N8+QlgIB8DIiAbfbqZjxpCnML2to7ElZVMsRoR+
ScGoAxyo11lHdpONPNKCFyuOjcRP9Th1LtAsxTomPgQRx3ileKUGkxhO/5y0SF18dl3Ny9IVszHL
68m95gIKoGFZ1K3yzay1llsoVTFKcvJliL9/mbs5xiz1mG7ZYjm+TxAHoioy9Ng8mXix5dYs/9fq
/aAwEqReN7ixL8HOIK9ZjOGwvwxE7fL9d4zoulTTor73p9Hs59pBsy29M6FILHdoFuMjx7nkBI45
DvbKtxDANi+pUJLL2cxnR2UFM+BAhp3Ds7hs0ziqOtC1N4bvBYq/FCY7Dju2unyPPlrtF0EtJW7z
bMb3ZJIp7QOo4xNTAvasgMGLwQUsHv4XW24c81BTNXDdHC7lfMzG/za4ovMSUnHcKy1cRnuXsfuz
PeSj+PcX/9Vg/JWWQ7my1KQ/pNfAVzdg4zOQzAUxAoFp+ntae/+2uUhmslAgVj40K0ObIgfmVyh2
jLT0YVcG+8siggLxf2QXxOo7MqpGshcmp63NU9IKeWjbQaEKsR0gqMVsvpEsTzGbAIFD92664Y+/
qfLrI1mQjQPnFeno0hnVF7XIrT3oT6Fq8DNKDbzsNc6kwTO0ZN14nca24yuUpmctdBBAhFt8fCDL
xBNoacSzImna4bLaWntHLQzJdcYMQuxsYIxxcxIx0YlsgV3cZQzRcDfRQPGUrD/0RPGWejqL7gDT
+i/06uUfSxaiNXYEmjXOoQUMKwqV4IHS8D+DdPSqTUafHdaoM2pmNASj+8tarTUh2HP49K6fEkXd
tkNgeWwcr0Omkr1U8ECJMPbG4/06Op2Qm75N27iOJ5wdcRY2d2SvHG/hxXxTbNDZFtIsz6AjpOD4
iuzWKM1eTI2ypLSBOZWzjr8NQL5PG9GgmxLS+8aM9OSOuX8AQ/3ZYefGZ0S7lJLv9ujXraqGcrOH
x1aUFi16cp08fFjfD5xlN43DoSWx7/Q9rMNg0PYKKPL6qcPMKySZxiVRLVjbELjF7a2Q14U9zTKu
i2kEYvV3kCM0NyE4WqqAg6+gEruqPlMs8GAEuOHPu0VMMPQx0FaZnopzxT3h1YyvCsoso7IYb3Xs
hXemsGn3ht4sJfJzl4Og8QfoKwsAm6dY+WRd7rdTyRKoPw7b9ZP5p61kVQWszYMHxRoVrqpJUfNt
fGWWsrbyUO81jPmSMAgd0gGLKEEvYu5nb7bvB31DrLX/K8n9sZbRrvsP1ARssgKEbY/IyYYIMRTg
q/bIF15h3humwkLwXombEHq0E0DARl8cYH1w5f093m1DbXpRa2AxxAA+1Sa5Y8BMcExIYzG4TCou
2FPWQV75uJ/s0Vp0kTtXx8u8EP8OUyQ+qq8dRB9+z42GBsVRfgEwDP+JXjh8G8g1P4y0CBAkOtKz
89kON9hZgKRKs50+lTQZSsJs21mrNqGitRjV8rN/o8N/3proQqD8vjSMfTvvatfBZGBrvWedlyVB
RHFo46ZNJbmmz58lr/HLY/RMGazHhgSnWYyTbyIA6oRAMHnuD0xO4JqdvfoWxch0H3Egl/n+PY47
Vr9HlTpelLZesCbPCUIB1d9CTbaKyc5S9hmVHMkWW2k0ejXB14e5gGuMAi1s+dGRiq8GKtmC8VOe
rKleqS5weFhtD3voKd2CDWnbzikEbpONvo90hfRB8JXBvw5sNHXUS/4ntuwbio6DxOJljXdqK5uP
P+qm6SvY79ye75PkVUYUKuQbzdd/AKCSwl+OJUhkgU5Z4fquxVTP8LlXgqGURtO2qlP7aElNuVms
AJvnDCCz1kh5H8BrF/ajoyHzCX5nruwWh8+Ki3smA9EhYg9KZVidu+L1mvgc9LxSQC/WCHHv1ssw
5l/akVjzYY55k0Ul9EYdnAYgiN8CHxE8zoaT16EZkDQ6KPhU1UtlUdI0krrEsI83kq4Xzkg4tS1Q
yQPn77er9zQ4VV4RwUC8kxbty76bFWm2k35L78MBOq7t0oUXnD0fgzIWThODHQkMOCTorC70CJj7
VcRrKsepQW/vET0DHIJDbZMkfWNpv/M3r0i8MX3sq13V14zNc/y5PQDOm7pTCmtuBU3KZp1J2rF8
FwERaINz+mtA63DVJJGKHbLx2WPqOi+D4fFOJ4ZWVvcFhFGs9wL8uPRxCMVtEVtZCW1hYIUryopA
9oqz1WAhDpzLaE/lzDhCVTmMLSkSrfQhqgwcRmIHfF2ZOrVIbBSlc3Igh8IRDI029vYh1dqFxSud
k9Mrc++PKOBkgjPAPdZ+8oPak2rCITIVN5eU74UgGlDt9uN16+s/to50GCCYndyQg1UHki3iW09r
dktmQDZHBnxUXmZOEFVZ2DQu5LE+k9EvunRXyBBRigu5KASdupnGEGXC8Vj1+UH8arBjdOko/rr4
W4tUnfMXKLTu4+aRkrY3kSwuyH9A4KNF+nA3uca4sKGbkY3v2ugBaeZZjN9BCn3KeVLRD2iLniGw
FUiaBYdNQKK3vg4L8ip6gF2rt036WyRKJQ5VZhlQvQcbBY0aylaKAlXNIDtcJnO+2DTNYsbaqltR
Xb7Scdxj3WqPzLxgoY/OBxrko3z60c/SmLXeIucSv6gR3ZuusPq7/tSnsFJwkS3EoXW19d2vRe3a
N0jAip5G0pt4/0+F9CByclWXRzoWQA74qEbnAsHVu4k+X/lc84Vy9nuoYA1U5KsqrVkoFq2tqxoW
eoLcTItNYtc7DwF+3SZbCGkqN/gATY2WPjE2dgktmtEIIMDNCfYf3m03wD/ZeQAKaEZutbGaTuez
K48pKlN1zTYlLcYWFzwEus10/q8QmgGm62Y2bCa5K0PD2kz62mE7MeztzLqLoiCXEmZHgDVPRWrj
HZHMysCjrB3bqOxVQh7sgx0+u2Z82BySeyRgiIHw/YShqBYuygOWkb47uk2TketZNhkwRmWVdu+7
1euyLQn8D2MNzXSS5XX5PHRsvepcbiSmMoILee2HuDxSldI1CJiajEvpbUezVbrVBzxsEnOMMrI8
XCVjPk/YVByt2Tu4k2w9bLd3K7aT+A2ZQ8OXmyUQSlt1sn97BZgLrlfiyN63X7LTcaT25HAqi7mE
BYKgVOJoeiVD3cEjl6NTgc1+nm8VxCmyulG80E3vVJHKgODu+IkuRg7400rN0aqyHNgYkmGNxu0u
44+DvB2DmUj/6C4VrKs73MtItZdnK59a1KV8dJo7/wuF9saUy6fLScRaNcKl3HvTWcYlpWR4YcP3
HcQR839WWvrFVcMvrdmQbFPIBvfTPvOU3g0hkAyXjL1g+bjPax5YkhZN26Sum4KuFseH3J3wgXnd
KfAuE/HiP1YiRBLPb5opdRWtCScvgYzLKn4f1ZtkrDo+CHIyjEyMPKTodrkdOpNmy73FoNPKEwbn
oN927xtz6b6X3WZCpvu4Xr0Sx0/W1oyGenKZzf+iBqqtrouZy9rcwGyELyZy+aGdCM+T0vW8UPrn
dHOMMAgXabGT3uutetDsz3uQ6NYbMf1TzeQq8TFhJ5fHdvJVW3xNWdfg+mk518qICXnAD8l4pD7K
sAINnTiuoHyzrLlJlLvyGA86c+baK+Ud45VRrLXSR6kETYLlrBktvLLeZSqcW5rzLiRBdJXtgSlD
lCs5+5j3s6NXli+6i0Hrgmw1oDcMYiAaq9V9oqLgkRTS/op/LSNR+9/+Vw2o1HD+jLxGfDkKH1jD
ayCFs8AEM2pYIb4T3sre+jMZ5uOfRt7ngGWb//lBAs/ab96erQQtGnf14wwkV+k2ucVNg+ljhLxA
uwLlpwih/4R3v1vxnF4+7zhmrLU0fqXzPDmVdFDb5+vM9ng1Z6LQqW5V4gHD9GM5At4er069ZFXC
29No8gD7VvER5bMmv0vTreVWtbVOyouzMX0agG/X3gpzRe4wG7nbpDvt4SefOrIYyMDuz3NFyFbE
8WnEpTP8MWRKyCTH4jq+BUvFlzR2YhKhPyAldmNsnum22gitFW2K3P5QacGKW1hqDzn9iErbTfW6
bgfCSs9o12FbZlV2m0wdIeoqY8ck7dJKy3BcKAmkZVtVtIV6Jrboi9lIdvK/aubPJUx56omRWBUD
7Zh5gXzaLqI6yN/duXPbSC0yqjts7o36Jjbao/Iq2zs4f0+ImrPaxlrheZAcRHnIFzuG25qYWZw2
wK6wneTUcywOTxcuVKbI4XwqXwEgJsRDpQq2UbrJAk0LM4FVVYQF/3PWiKRuQ74idACQcV/g5fv1
PtU23EkB0/1urmYuSJQ0vvRepEZZaPKR7O1dbxY4Bc/wZY8MJIyvqTsmCrGsB9+bprp/5GuQUZqU
wAMwUHg5SCDefQg7Zl/Qw3ZJELDTZlLarJWDObOjNjkXioXfErQgMH3pQRPE4A0quM2F9rS0YeOu
R6fVbpM8edfa4n2+7yLsEsw6itTWx3w+tZdSCZNDy+SK9J3dD3FKDrVDvO1bGrYc8k70MHW1g1+1
QonsSNGzDzeLm7SWlMHTRiz7U+opsuEwzdUFIdez1dx07oePGLHHO4QmVlCIkT6PzWKOOCCyXxeB
gaud6n7aOGhLCASmx8h8RwQWOXOCjbaDjQs8Ri2fjjuZAfk4yxJJ3Bp1Gecbl3yoO82+6eM199QE
dJRM1mHVYuWGzEVtgtd+drQx9Lyp+DJyhKNRr3tyXYGAU4mvxP0R4yAzKr+NI8RQ6inPisvaLuwz
33/YHyxJK+4ix92eQaS3SunbJ6MtAWgvX+s8RUupKCwUM/+afjx33KMgxKwqITeP93PdBY6PmHlI
yIkBNLgEKa5XEZPzOEHTmZJYVWfP/liySR4u88nfHb04WmTBsEyYYu+aTHijzYxkJRHWwpwnbz+H
KUVXLYtdOr3b5fawHrOzeJWR8zhGE6+ZCyOj1ze9Voj8tnu7AtSsR7Ipuv7lTsAtOiWN0Ql7uMA0
AH0fWVxGC8ohtpRi0kan3yCEzPajglUn7wUTAA/mDJ+YW986ri970CsoVdUl9mWXuzULpg4XsFlU
O4Li+kaRtCVrRFfD5O7LSkhVn972TErY3uBEvH/bMFeLmUAnrySIkFmx/E+sBDecJpqM5XuPF5xa
6BxvqFBqFfX1irNDXLKKJt6SIPxs5Ep5/eTcHGJHko3cSsXS9bStFNPnRXebF5pxXDtAjH84jYd3
fdUKa8i8ZOEM1EaZwnzJYrtzmf57GngqeYpBar4SMhRfya4Bmx8gUh7TJo5aEGKGCBMe2hkv9rRr
0kvjDyE99zE0tmhZJcT8MpyYDnzsWUgzjI+Xmjxv1y/mjC2k7HWUSBvuIHPKdUu9WfeOpWKQp/V5
AEznlpRRFB/6KgsFpW7jUZ8tnXxBoSv8JJE00FlviOag42cx2df5SNv3O+k6JEvBi8B0HmISp/dG
vK0O5Jjj6yPC8MUuIS3b+oU6oqezC3JyhEEjSYX03oYpMz8a09J9p3yATk3MO2mUngU1Nc7k72gL
SnOYCLy/xh2yt8f5p1+bl2bDk6RYKV2ynRbUXYkh8kWh9TbPA8Gu5aBuzrHvVpFuOLo1rXPlApty
ZC3B8c5mcz5M73TU5NjkYc9idzzntrnkZvY/AzRhe2wwck2IeJFnGDMCZQoyxBJvLBwFeGaX6GoB
pGAWVLHtNqh0f490esccUDTQ9TiNnl3j0wEyoly566UzVy8zxP53C5qqfV0aye10vI/wpGFu7q/L
Ln+3i8dk4ndNVFJfRQsHiOzThgKsH1mwB2DY5p6sgNZigUB10riJkoKhRjRmPa2fbSRC2nNivbG+
8jhdyNMS5ROgmd8kY8QvbrVyvwONFFSmMBmHDUmdYb8SVNFfUuYziEscDodq6xtnj1eTY9tGfB/c
BwY/3tJkf2Bn71188QcEZ/9QhfH75pHDL1hvUsaprFtEM+DyKRPRapoxR8HELvtkOCmJM2UCsaF/
0xn8jk7OsdGVj26ZhDcYLWMxnARBCvhX2iFkDpsbfmrf5sPek7V7xmdYN+0qqaHGPDACDKJO5Nqs
Hpd7e2QL4VSEPxvrPZiagVjdxIizuOpkFgDn2sA7jsCO+UgJAdMn4ihwHhpzV8PMEI++mr0MW7us
dMBQLX30kRgu4JSSScovxndBnmzhZUq4yWsBNtTXnSHcOkS8eRpMKI0X7OVZ0aq1ik9XB0eJInLc
KYQcroydu3La3u0FU3QJmjlMs0ljyAIA9T97NGrWIs+QGLRqqA84ICTEsjEgOwuxPWleQkKAAHAc
Oe4pFuhshZY1yOQ4RHZlS/g3Fd0Q2/PxTTxGb/SuQkXPTAF/Oipd90+9qmscvH2/CejYrunecLg1
96Ar3KCXF1YdJ1by8aJ55LZdjlXnEnAjL9mMHZ3iTuOkiDZS4Qli1NabsBioB5HcsYIphylvEI7E
Cepy0u4qVdSGMQO3fgyyGGjIwGhRFd7Ygap2bmujCqITRELNoSVo7RO4E2gnaKJfQqcdf+NtbD0K
BDZGP9avxAhixiVOGJaZeLyBKsnfGlYfVu+7lJS9QVvDtTAqoe8pTxggcNTSN2DTYRU5PJ2HiamB
+2zvHGXJJ4Qc04UUQ+lQCt9+v6SqNUpkqLNewBC2m1DEeEbH+0+/YI6P8eoCP/hm9m78WjZ8row6
sly3PeCsPlJ9g8oxFIrsX7m8ZyGz83RYKi2hRJslKG8pu+hiB9TvVB9avS8mufR7jxex7Rl9YPGv
fZFg41nbwn/X/E8ISZLQueJlg4C8vlXNNtWVe8W+faec/MvF9ObYtczyc0xqjQ7ruRt4WIZ6Y7Ag
Nm85WWBDe8KYgmlmlzaQjJHZ6e8q4zLmwhV6OkQp+wBoiTfRxUf7nabSSp3XovZOs/86v0iAIL17
NkzKJLSP4R1Nmkvd1zor8tdKcfZ4Z/oI+cmcEjPvjOwlb8Jo0HKZuNGqZ+eiJDjnCjJrUciMd7Tm
Rt4OUqk5fDUehCcTkMYpmTKOgmgOQoYvXx82Z1IeeCPRC8eQcCRfO/bidyDHCKjjeR5ofjqAt28j
+Nzxkvx438GqXbcYMbGbDuvhHpCAI4qCHvA421jNnOlgaq5rz0q6v5dlnJGqeR5gc8vrWVCijxvJ
iaxjrxzLXNaOPVF4v7NuFfddj4ULouhEG/Z5+sLFsB2mr62jDjdse5Z5NSRFO8SGuZwLFEQK66ff
YT89iqvVLdu1lyfy+GAr9HmDXtpTU+5t2rmJ+Jt/uPl77zZ+J8D8F08JRBcIV4A1IZDEKOHtDsn9
bMkrBXeXkGnpiqjrxiB9c/2OQDtLLRPV9e1YARAvSftXeUXKDtETEZTotPPmE5Fatkb8R1sWEISR
tVS7C21IkAEeookV/M+vTpzgR0YupfD6fS67vtmApka7qExQp+rFbZsY99a47wmgZheVxsblQxAO
4XZ7jjfB7GQY6EEq5W7gq1636A8k2ohaDJDYxmgZIHxqhD1w7m9k/YMuBuCgq/BNFUuyEME/IrRr
PuEgSEvfzTG32XDvft29tgtWitx3dXScp7BLeay65MnL+hbjAyGkloQ3FB7EmxrteYhCl9NQentU
txv9aor2JvFW2oJIAJzk6JdtFGQIjGRFbQsjr2Nk+cTf/WXcd+09h6du4kbJCltUksINHIDjppy7
QP2qJ7NezwAZC8Xk6fO5s3TepHhuj/J6pcKsdGcCqy79EikVPH7qDXUXvJfNg87w2UJ7o/K7ietB
8Cf37sWopd/QpqcE+Pprv0W+U2r9DtWQYdePNqrXlL5eHwS8aa5dcH/Po2/M9vZKuyrPz32zDOVB
WJTUKTMj41xdvSD2/kV/HvR580dpeYJ5bwSOFiFOJqt48Cqyejl6gHwt9Muzx6iAfJO70dL1UFPi
1Ppa0s4slssQAPT5rcPnc0/q2G8ObY7EBv1uqa6SL3ON9Tej/+IE60f/uKEIkppCYmuqKlhE1R/j
YCe8O+o5DymO+xVOkkThT63jXJrausP3erjeQ8tnbBAi7Gddw/6QuRJs0gKgtyHZoYTGiigzlQE0
bod6rtOIaBKJBxeUFOZreNADmNljYnD9h/j9ssRjFjqRneW2TlvSKS6N5SBUAOwt/3Kf9cpdxS5j
1cFj9Osyn3ub63ufbYG1d7MV3ffghRFk9pjT81Sf+q2+6urBVGVkVVcEBE9PeWdBKvET6EBuZ69W
bonMKffd1v5jcelOSpP8U0GRvqkSFz59hGvzlj91+DjjSwLH2krt3D7iXupnUxl1L6Q11hkUCc/G
H/nKkXYuIxNLh4o5XmwFe+N0F6137SojAj4Ps/OXY+i+t0kPDTo8ZkEVKmeS8pI6t9dd+XHI04xR
ZuPXH23zInuoTNSSJye/7fdvQ9Po9x4WqxWudBnHrayI3AaM/o2lDz4c9MrESwOsRmUXvJHBTj/N
eMVj97b1pb5sjACkW82qjGNoc8x02TJBWb2lnhWc6ZKYGkehDkpuIifwV46937mFTyMD/qg8rpLi
CePs5DBP0KflQk/8sAPkHmcRUpGCy9ndCbXqHGyMuS4Unwjplt3L5QqtBDggha4qBdiNDOIr41fk
Ew3+NCDiFVSzggrMdbJTUP8Kz3JwtXJPiNloRFX/wnzc3CYqYyINdlTZZpjHuUCJr8iOmfw4NI0P
ItRYY+Dl5CwWhH2uzzvfCHlgWzUsUGsiLogLJUDK6cEOOWRTTioUPhoLCY0HhOiv4HFxPOjdp5D5
HMpjf8gQTPXnBC4ndkfUkcVQTaIzYTJXcWRr52Q0L+1KDUKGnLdMDNpR9+LkzYeOIGzaBac5gs4C
PvFccCKncGW28ll5vqU46UIOhkL4fRJfo7CMIKqXVJIZo+GjrvYznD9lKg2DtuzVkISSeLqAIkw8
nwJTBsenvkWoIL9FZ2pwbxp7Z/Y5VT2FDYqbvpwly5sAPYLMHeC2Cv69L5QurepTG+oh6qZJAVGe
24TF2k5cuaT5OerzdJ8oQJaU/SErvWI2HxvzXpRN/y6+CUeQhS8su/aELyrXT7EvtBIxKMWwVCdb
AeYIZOIZAQ1I5FzJxpFzpDAgAp+ZHQc6NREpqcV342hfrPg1KFaujmHBioEyGTnOx+m/hmq5CIJE
Qf9gLJ7teWZlrDHurxXmnxWz8WYH033+NWNVjwbyCNCYkcKZi0UnCcz5Vzdh3LHaArIwqjNNhG+A
dZu5nMxmmtcGSeANe9MKKNTbH9NCYGeCVio7PxncvWvm1tgYAQusmKvpauLapVIzR9BVRPwqjAAb
rq5mpjDa0UgPMjHh86tUAzwxEAXRdSiqK81UlvMposJIM9FiKjXcWBYk2pqaLVU+3FiUWxnH/xmC
1jMoWizua2BouE/KWFtBY2Sm2mn4Hu7qqkphxtD6qSHqIyKhjf+Ec8LJMvQVxs1tBOc1DLuu58+T
MwH6zEJBcRWCklwlsR/+JQf3zG95bcQqAcjSgUajrnyR7V7jzGj+6MJ3pThRjI2sbAnd5C8SIhuI
Jjr2cmzMjCZwxHdcHAsQfokFtyjFHdnqmUwzsHsw9MuL7gJAoRu/NwTLL678Pv++u3qnpC/JK4Zn
DyTvPYnVDrVzB4bVmNO9JwFPMKwxGfmE/kTARIRtHgePtY+l8haaW56BrQH6X0lE21evXHx6jdu0
EctcbviASiT7sAC3w9KJvmcKDDbt24qX1PipNHemuifq/liKt39rzIGoJe3qavIYa0eyEXHlNF5f
Strq7XZVRf8PWIcrUPfyfWMn4gmVjv1+N3v/bKKubFHjLMjygfSQq6Pt2uZjpe9pnkYZEjjrQ/Eg
7TdTRF5BMW8Z7kHCsIv7H8cyAElA9NmI4Q2l/JZqWss1nJgkJC2XhZ199jTddaa3NyL7LoCpKvG2
erQOl1L/jZjNZON2jKkuRSSBAOeb8IDtxU/lTj2BKbSqj+b2Pn0b8vNpNeFt0bf8R86OCI+ulqd/
B72K9B1jf3bNa1MmtnWGtcvvYAMsM6f/jtgPUjj++NNfwB2kXEPyT4gAbAxZglsXtzqrvuOaIvHV
C71ZOz/4vgBdztOGoH1WzEpU9Id1pZ9E+Xpv814BakaQ34FWplY8GuhqkX+nftQ3mByZ2vMoSuZF
KWB48uOiZhipjAMcRbwm3QBc9OuNyQ8ATcasJMCCOTJdSZEymPEkPGCONL85Td0nhAmXxEl7Xp6/
8GfLX0H2ZnnHNs+YTSd84RI2YHYPZ7ORLUFgzA4a/QbX4QzbZe8KDnsSxhyYVqQxF47h8L1DCyzC
bfGh/p7gsBdiNpftcJI8ilAcP7jXy6ASXRFw7BV4/ut8w8zqOpe6LGMxakUY7AkNlb8pcdUJ4t5Q
YxhPsc+6JD9F9n5dQ6bK3AUMQnv9tOv4SNptUvn1I7K7VXAMLEJKXg1JhV1ezax5vY1LfFkbTrtW
WErztbDVMyUga8bfXAy4x1dLPf9belCOPrpuCm6pqi36UfoTFk1J3yGFKEbzqxtv2y0Seljp1V5N
K0Xr40/D7pYT2sD8DVQmZewAdo91oUzcMKHPPez+vnIuCIZ/cxWC+Ns/Sp7X0Vcmt095Jt5wIUxN
xn7GEC0pIVYT1dbfpmKABm5VydKitdN/Gh1596BWBb1GPK8+neCoPd8dcY4ZQ36YkWF8I5iVxEpY
uuUdtTuD7p3NfBP0OPDgkA4M0QKAMKHFbfvxu5XGrVgb0ckLKGvUcStXH0ZVqMLA22lm6uz3O4MZ
zGfAeCV8qwLtvjsXVx9mPqwTx+IEGKgX2BQyjx9x8BttpyWegDbXbxhlvv6vzDCXO6t+3xh5dHtu
3VN4Gbn0Va52FQ9o1U/QizDkYMdla8dpMzV3InllegNYLHypK1CzxrSDsRx14ZhBC16CTQ84m5to
fiZOVM8Pi+5r7KPJqteeJJa6KZyKUpPXPj7F1dreAD04pP/9wEg+wP4wUFXqAoG4C4JUUH//+5PY
hlL7jZiBOPjj2j4NyDh6XtAyNLaYVt4xUt23/0ABOLOKexj8PUnjd58tjPJQXQ/jmpz5fQ+I6VEf
eJV7JfFZOthoLInmIyNKIFYLisPvXDmMirGgDY8EPOqlpf0S3t4IbZtyn3lw8bJIg29ndzaP27gs
VIhw6I+on/qP4xkOpZogsLa3onY6BW0/kQucQNqnsp6om2lSQW4AJYXQ/UZbmOaEi3DfFOrdLS8D
+uQT6GGxG7rv7ZyxzuQmOaLIx7M2ERdNUh6B7Quy86RQC7GrTQFH+4qY2yLJ8khyZjmAPoHpzvEe
hy9FBScCLG63tI8Upj+VxbUhQ4zgKkdjHLFsECmF0y5GCmoNrg5CmB/PGlumC7plqZvU/gWnLHbt
ny5t2PFQ5RcdscEebTFpr5Ka+YRJEjA5gPFCUOgXyrDbEw6sQB7eGHe1rturECYyvaMSGUD88TTV
9WQIoJbiL3fnbNeMfsZ3IfOZebq/4Rx1N48fwn/syaodLRDWfNGoHB7ojEMXk7prct40z/Z26oMk
PDa0YGkmvlyPH/g84cc7Jn0CSUWVZdNFWdR+0uboOARNan5JQASwfqiT9awb6wWLNEoIUcdYAntz
wOyecbSkLiLlTsMtIsn7FOy8Ir/NFi1OxzTC4OStVwJ4z6B190M9BEHd0TktOErIoueYASfPFuzx
GIoVNW//ZK3IUurqO9mJgXHYnH/2KKFY8vZBb15MUA8Czeu9pvFqtEa0evlw3tgkuObXK7+AkaGf
coOaCCtK9rvRitMsOk9QyP+cLPzPoaFGYHwvDvR1hkynxYAlnzGfI/cupZTLCxeihOTxGakjoWCP
p3b2j7xvgLYXWEibC3u0+bGGopHaHwAwL95bz+ZOGU9j/NjI+XrFZhiv8Y+uGLrAsjmUYfoYh6ie
6epcbm2RaHu9Q5xLyEu/nfVNIfdfFxNOET0Q7DaW/uGJIz0aU7ipegprmy0xfYO/xi80AypYZ9MX
7FAFNqKskE2VFoY6Lyt2cfxkz3OAaGTihlhf9/ri5aQIfBaPH2DXpRg7KxS2raC6eUDAoHiaGaqD
jvvvZ+iZT8m/7UytMvME0g/BOPv5+7DMHkN7llnDpdxqQvnLOI8WlCEREfsP7zF6en6zToE/0kVr
xW4w2AtH5vZYX3xOP5dhDWElcbs40u3EyFWQ6fKAqXWM9lpDpFqiJurvaHQdQhXdyF2hfyyzTDpa
fJ86H5BKtxOMQLqS9zQvPFYnESvEglPWNLSsZL2DELPbyLJFYnEfBSJ2EPoU9Q15O1HI5EMwBKLp
N1HC+lXoQtxXIAjfXXhQbp1thA8m/Oj6aqupJmArAX6ADE8gGZvm882/gLE08UjmgcA9XaGbSoOI
zVpqUlgJMrQawd+feLDdHcbLBLuhy+mElBvdiMXmb4hh874yq7Es60dWZZF2OuBxIMoH8txL8UrX
lG73BEPJoyWs1unA7DPDkbsHaRBwIlMW9tDTq7FqLPfSxjXzbfUuZfaeeKcD+ECYYT3ul9mcQcJU
uEDfKU/EC5fm2N66LfkujODaTJSC8EBo2NXVA0HBVyUm5IR+umNE0f8A/PZuNj57JQGsCPctV3A0
1yBJEYYnPZlouduwlYYskdA6tNuFyT2orBFvTBdnloc17kFcuW/MvtFPhJ7el3H5Hfzt2dsyBNsb
I05Xk0jYhffU6RFhr66kM5agRUcE5+6wWHPAbU72+jcCk8gfB5icFe3xt6OqAPU3RZRvdUBxZPCl
CddMrD7hFTXNnYdaHgoPWGgGeCeENptb1yCFwB+BrzAho7giO985e5v8ETYtLA1nSLKDTOFyf7TQ
SpayOLGdHjfTEFQSu5c08fAbr9g86XqYTFneKm/PKfEkJROqoCEu7zG/ntX03YRhH/sYmcH8lpNq
My1wUN80Yt1Q5c0XaW8YL3rqZOe9Ptbc/yi8nCGCX+PcIc6j/NpzT8tRP8cYZd6eOhD0kqtPfJm0
QFVQoLsS0cZjT9rcyUfsUHHelsaFUd2AMH+CLKfLd+EurJAwf1odfec6SWjzjhTfvJgrCv0XqxkN
4YQUssXZa3cigeG5U0QvhE0HcAFcG7Y84lvi+UkJyaijl7uOuTqV5sjZSfyFjwoLWiO2FjSc8OiW
xhP2J6FcRleJfZCeWtHYPJ6VAFcH3RR6Mnqsh4JICuoVxAE8+fkIxn96VcG8fJEshDvpwb9gJ9u3
OYklsv59DAnH0aDtJZw2vjSEl3JwAtByFaPLd+pq5VWk6b89vsVwi0+7+jyjmf42Y2IOEOJ3FEX2
nHvVZLRCo+pbCsuiDKnYavxX/27ntDh5LhI+hWQTvjyVCxhD1DcmHIr6AKW4Bs3W+U1CFYWpu1ZW
EyYpbsZVaIQODDFcS55/PQ0gOU0ERIaFOo8zPY0gcf9/LNuegtzK7Drqdx/q8xFI8bznhduVuP2i
oTXMTCu61a8zu0BdC68XzsCPrstGpokTD6KPmBK1hNow6tKvxUp3j6kwq7Yyu7MCBrHqD0hzvCaq
gr8G84rOqyfyjhV1lzwgYKhF74IGNzjdVBUysZZKaqiQbm4NuCohJdJwndeQPkpPIMRL9WvJ4F58
oR9PoQYwv3BaKsugYK+HB1xlu7UnTg0A2VbHITHNz9sjnOHlHzFMTL5l4QYsPeDK0BrE/jNAZsZU
1iF+W9O3fTYHr6+jScTc9cUo7GN5cp1rPCjloLKfvStjQmuACPRnV8szt7zFhtRcl9avcaRBAdwJ
ZM8Hekicqx6MjpeXyBSUwsn4OgJFabjJpS2ljwjn83EM1nc6DQ6LYjAX0tQA8GDbaXuAYp/5YRDh
9mXNsB8z6+vH1O4EFvXHhA+7OYuxX4RV2DgQhSbK0x+LV76cPNzuFw1KaQV8xgSZR3t3cqFxBS1A
mMwcmPTX7HS1RmqA81LZctNBIgkgKIE8t7oYPKycwTVHGOQd549JyaaPKmgGJXbAR6H2jbMT3bLA
a8OHTKn1LnutJKO2yXdu1sP47sc5lj5vpvwOgjU4iVucANiigBZ7zB1c3XUdnbrHM7m/C8NkBxbS
iWh7ng2/iVzE2+KdSu9taPidCaomc7zeM2EErt+8qHt2yYPeqOItH1s46JDgBzsH2dm3PzRMpPVP
mk6vHXajKLcApv/32P2OuqiF+RldCpxg3bqZ5WuQO9yf0CwHPGcVRnA6nhUi2d/o0AfvinxC6Q5/
pUrWWe2T2Pxp+NW7smvaR4ZPX/DMHyhwHQy5RrLmEHPkvL4A2WaiwXd6MbIN4XUCtT6ob+SXRl4C
NwJlMkADCr/wZU8Vu3xNlc9g+2E0Ane20Zetf5LrrjyCS52WDqlycY1qXvdNHKeiPepn3qLxVnL2
kACbn8Xosz6sJlOaLQZ8YY/2vt+wa6c2CgBoch+huqfsQF/xN7gi7vv+Y3IClPjC2UhFkFM9bhz+
z4P1ITCli9RAUHgpL3KSQnKaoH2C9wlxqOYfT5hUMEzJtWlAeii+oGyUPHhgx/NPXWsVTeZX4Fsx
GzFisAuUgM2HVZRWlX9SD6Xn/HJe5CZSjhVvY6+9Ohoa+v/jy+6vQjiIAaPd7XC3VA6mjs84RPSj
O9tCHrQ3vHKVCzGpCQ+8XLLSrTJOjGqL9GiEiKJkICvXfrEn2CzQ9948+pgwSozx1rJXj41SUUE/
B8v8sKy2D7gKs5GRn7cMC9V4Nar3RJ+I9JjaBYbrdfrss0Ujj9sBPNE2q1UZvk6ix284dR3J0MXv
y2/HPFBXUvTapN+LfeRUgmsnI3WjBdHfPUMyh3Trh+r0QcwFKR8XJrTXz6NxqQd3IxfHaA4j50E9
/4k+IlZ1btK9KbPKKXNDbnZ5U98Y1Xb3Igp0QzNpqybLyptHLHN58dRq/7Q0teuy++VOGoEenQ4y
TZBlsNhXRcdUQ87pD9rkJsJDsz9M1PeXF44WcSqJes79Gy27bGwyiyg+DYzPSQBXDNHTr84O73yh
+ot6Lgh0ZcnJ0doY33Mt7ymv1G8Gg4Az0ZFBkjAFnantQyc4Pya05FbbuZ4PoBDDhmM0dGPTZseX
YkbvuTF7CujOc5nK5isOLjsu1hUhQ3OUj2jKtNdbeSd2YwGkMtmhBh8x2M64aPgfSuB0K9/ydJYb
0iKM4oZBnber/K51CnOpZ9IhIzUDkz8SfGG6T0IEZv8YQHtFeB+UUhVhS4sBue/8sq5KSYGtWX+r
/OzIgXoSrCpJx594Awhc0yKXs38JOCUgK7tDPQWRDEm1EfaXzhgjK4+Vd/sbiBZxwCFfLmUNsyCD
cD+LwwL6XyGLmV6eIn9PtDUgrPZM2PUdzoTHlWDQgNgUt96hNJPe52hwKjfKX7K0s28ceVzQRTQS
vVKJZ0wfj2Fs6XwwTAGH5fqsDxCzkLMY1qZXoezwmbDvAuoYB5YHC0VYkxwza3928P2hA3hrZIeK
6gnPAiyp9t+O8c+s/eBvXD60irxvu2TVkkJk2xGaz6Pvlw0UHxbhCA+TErSlTMh+7XRrxYN90A6a
U6QH49iMw8mM5t76/kraKh0+0BgujWNJCFvguAtTXKVul87YogzuidUhwmu10UH/KLwdM7QgWxB4
vPB1ChpnhR2NAXhOd29sBaOAgfKrq+i+c/4NkPb5bbcIf66YmNAUlteENpEzyL5aCBHccJjOZuKA
U604VEiFk9y7MO2o52ke1y7P+nhGukxSdTe/eRdXjzpAGp71+/qeHgzoT50FLQO109GvkuhclcCC
dU7nm0cogSNZ13vDXRnum+WdhpQOmevRsMD974CyaFnVIaK79OwXTEk0BdovKSw8pqwVtPTwuujO
ox8g4zI379XpdutXQIltWGWt20xnnBi0Oxw2hfB/dhTpoX1XPSDerUplmzHNWwSu54R/AVe6uUP9
XWIGmclan7gANlCZ71yqo1ZBDDlWyrZrhgqBbX/ltFWgGD0wRV70MBLOZ5cPk1LdHUPZGTd9hyjs
C7Hi+5oyABL2mw9HGogjAgEnVqM6+csBGbfKhDDj8ikNXVAqy/rroUnxl0CtjCyI0lLiWKVBy84D
Zzg5K2KUY5zVdJoLlTezj5aV0Kxlcj7+IEQdqGr0wn+NjMEA4+9dOPVLsUjcusY9cN/khvNJjaPn
Zl+LiRlgJM0ZGZ9e1O9OhnJbph5Q5byFCi38rUE3HtEkwUX5xvcTUw/MjkH/ov2F7XoE833M1dBr
guc8ZVgAdA2znU0xSjs1nc1A18YYXBYaKLhGecTFLDWyF6+i4WihlhQgy+LjubEvvI/vFx0if7oI
00W7gC1NJ2CxZQW/OclFmyTn+IHQk5K5VtRloEJn1ZLESleXaYOVA16+k/Obem085sjOUaRJxsWB
EMJCGELNNL15Y7A38xb8pnKNXJTzyPkV/aOg5lbDhDOa4OfPyOjM38oAB9vwF+DTLpQwzXW8r049
wqvqxaF+JRUBsIEvKInOUiGVPUKGx6yjkqdrL6dE5qWBYKys5a2GYWl/IhycZCs/o02oPkWqdPBm
TdesX82QZMaoObVLT0UZRkeAPGqj5qtLRqoXqX3iw54MRecrLSw+CNPhFmKHGPoQUdqa3V550c+T
fAiBwKmQmyintRof6MagLOfP+/FSdfkjOlSmZqW2G1yY9sBbiftEfnb/6ghp+CbVXT3HTm6NzdF5
/6bHt1jl4kWkGWTyhrV81VIOmxoRzygrg0iSfcl64aIPQS9csQKyodKTNulPdOxRYvmjumckyaSE
mm+6hEf84cTqGabyYTDAOkH9lEzs+ImX+t/ug0frnytTRig16Nvvln3UAOlF6pIoL8RfikLF2mnN
uTAL9CObNGP02ThdhrykXFfEK2lKJHHxRJftgLh3bpD2ePbnzVKXsYUIU+P4Mvwi/ra146podZCI
H0JIAWbuYF8PYfLUl82+aW5aM5qF2G1TKW9seeeBFYbiQR26VuMo9ABp5pwKP4KBvcKcJ47gO/zQ
y3gvggjCmqg0+U8FgRimKU0w2eTz66GkW8J12SjC1t0M3rh50PX3wQhtafqGHImmJMDG+bF52djr
IJ2ZV3NtiDDEgwZJrBR4tr07Wx1QywbicgzXxETYDEV5p29j55VRHPz5OGQQ0g0uJITeEYBRddKC
VV9JgJa3idM33V7y9PnOzSaFiIaAUBgbmLNiViTsv+h1VqHdN6AvN/lBw+gaAmceVFoWpFlfogIs
WTkF4hLWTBGLd9Bw3fqMhdVHq5vKMByX1g/KNhEwcmfOwAWq9fWU5ZYKaq2DOCLunw6w7XpC7Hzc
T9oTgobh3ULMlz68CZwjBh8l3Z1F3joP4B0F1nvOor2WQqdNVlO9OoKxQ1KeyaugOlsW8l0kyh/a
t7PyUWy/KCBJ+8r5J5vLR3PRS9rNaZj4+HUUvQLWMwnkLzszIZTpRIcdKXSmgg+LL9B1Buo/nAPW
iXwViCMWhR6D58Gx3hRIIh5IvJfQrJ8MouMW6lx7uxX6R7XAsxODYkvqNJpfQoFGW7i9mu/Y9xjD
3cFZyW9G4qZkMTb/D7EXYa36pC1Ijl/bJWLclK8g0TG3oUR/IdBBaKfOrRfWuSXYdFrPM95HUJXo
Hpr/DYuxeTcY33qZVBjvLHkqPy1MvuBhog0nXEDytnK6nPMx6hDiVlEla5CDf+F2pr9iR7tHILxp
J0OUf1ZHfcphj3Yfcjz1eE6HBz9ZYQ2fDGgxuVweN4AG5lsZFM3IhbtgdojhrYproQYl440qBpai
qCry+n27D3lmiN8LwfrBCqkw8oNacbtBWKotD2XbzGUoF7bgmAn8r+yJY+IeAaem0g2Pa3bAU6t4
0WsFl9mWfCi0cG0UeLHnyrsB/Tx+3skTGw0FwDEgnR6nkW5bN4+nDfRTb8jnI0hjFZ9FQP/Ol/ba
3Ygmo7qkik2DvcxqBefG8gVFmvEplwWjPKH2Rhcybt7WPt6zKIlGNxqwRwq9BSxVqq1YkTJt+e24
R6dfoGNBhL3F3X8MrwY1KNp74lTU7F62Fd4Ntq3eblzyO5vnO7Z4VzQn6s6wvWfozvVRyyYFGUDs
ly13hNoNXo9cH7f2zzdp/UtFpAcFEWZqIx28lF3lwlxXUlTnpZw28FXJGJObp/YBfDHndjWaGFBZ
m8+KRzP82CORnlYVYZ53URK/YT2d9gH7KDOnF93t2z4HARMWK5omOMpkofn0pmWg8WFvdYLSJpJg
eRhBB6A7U0vkFfp0+9hGbFQ92mljORslB8z02MYS3KfBh1rE9I1/TAICiwwE9tqspS1Bo8/eXwhw
abEqIGutvlwkKd8YrCG8rAGGuzjK4DsMKE7dZ9csfwzoNAho31qvXtYaIUf0of/V7CGtPCJ5TgpS
zp8lu+SLCuCGKd1n9IWy36oD53I/Wvj7KVVNgjxpubdz+dJ+P28/4rPb4bzgdL2cXDGwHkuRU9ox
md59T46IXH4J5ctkqq6Z7ISQtjpmAev9n0o0JBe+mbKq95i/Cu8SGIhbEd6eP83kN4VMm6pTrc7V
7+EsgQI3CctnxT0XslAE5J+1CrL50TWfIolFCXWMh4KEcCwR6hX/055BKUGOIVt1H8Pn4NMn3f5v
CDJwliWpKh5rfwPl2I3MuQhNLoKO9Sp3k6+gCwXaaXMLxsWIIMixJke4l39RN4QEkmjzTQnR+0UV
WYYCmkzA/r4LUvTDsAMye9ppKOCYRNxBTbVe4uzuNHqnkWd+VfucAG4GA2rJueS4k8tVp6L0xF9h
7P5q5GBmjVfXs9eCRq7XciiJbFmcl6UJf2ihWoh8UOVRoIJJu/CcFhwEXngVBKDgtObeur3h/IVh
IfBcZcdjghHNK72TdKiBoTuQxagfBMf/mn3nk5Si6k45PRamM8Ah7YZFCKhXteqeoXabwJdLNd+1
ADfJxNFcVamjqWD1qNYzzd8QrAXPA/cb9afKL+hVwl2QtEfILIt5vQ+N53qg0y6h4IOW5wAFiaj0
NlFsPu0cQjggBd8q9CT0pba9g9A0XhhuOBXvuf2hBnrZSJTrC3SL0E+vx8k6K57j/W1y7c2SYek1
pTkJqrpyiL4H1QRap27VEkSkrIiMoTNGBDtNV2RwIOX1nVsVNJd+7m2DU8ti/55ZVVmTRIFl6QrF
wd77+D8dZJq08PBRR/28AYdo8MWSxmQ64J37pLC4fjacrbsEbMHAPw+Mns8op+csJiiVCs2icIRr
jqERtaBU6XzYy7e106aG9IGr0emMqXaxIwGHUWVo3kByTs8OFXsgzzwNDCtXhw0FUbSf35t3TBES
PdSMJLsL3R9MVCutif9PzK8jMfqSSuGAWLV5gQmSf/+PSV+UFOQYqo7yqfvr//ckwkdO1dcFXW+P
svEvgb85D1B2pQ6nIWC6MTQmBSLC6zoy3YZNzBJ+kOp5oOXDEY0OXKwb+bu6S0zByX4LpRosNqZg
kdeiGZ0nWFzS8Vu3YD4elVTXcHoDUACVk46V51hTzkJui8lpa8+ujSlUT8kQmPaLr0d+gEaAayDw
ubaGttedPBX9J++gMuJhG+nZxATzSb29h9wk4ZRVWIJfv7nrqrYj/xkE1590kpLokubTxxqKmQtB
TcvlVtmT2GoyoLN2cGrVdJSpWW47ydoyfk4B27IX8fNYhVsOOvkyzl1bkj5AkxdHnbzeHw8HaFSV
FT4q29ix+Xq7GGorf2OOGwFWy0v935QQ6nWtT2C8+VL6aWIkIZzsx1m8xMKixhtPkB//LB+zE4U+
MYga1BuE+dl9dL94QBWzCi9JNgqMtMN0knzngnwS+X0fpMhKQHJx9QGGHq4dfQ3U36biMulYb2rd
M/3tdxAAL2lhgqJxuSIjoMDDDhDo9Oy/UmAzdGcw59g5ZVRpz19JgzihGktWsWQolu5sS7ulTyPq
c8em/qzG3JGspq25Y2mj1n8KOvOOjGnmgO3SD6xUdkXpZFG9IP47T5djoCh8Og2+JVdX+1lZzdvL
k5EMDf5OdCcOLulpc6z+bPqgA4ccwCj/XASeyaVICrp4Hw1vsuDbXEh9bWChkvwlxcs85flT172O
C7eigbubz83Fp8gk+5sYC9PWn0B58nVedEGkni9VG28G/M4UzScH3dlHUEbwCgoISjQG+FtHSP3C
0N/Vxut5Vm8/MJuy0sblxWRC7Vbh0zBD2zAI+MiJk7dxPd6f0h1v5mZ/QX6FfaMgqMZQ7O9yyPWo
QwhlUP3UvT4kiuP0bNPfyCQ8Zeaa04zyBxU+/svfetrPm8RamHhqveTDhLvDlq5lvlWc1URUA3AV
kZbTKlXeF5BFqxfEdbdarqJuiOfUa3TYpHM4Ecp4I2NckEF3u4tjp1H31FR61wSPeZtgztq35/1q
jyJSKxGI+dUUA6gjHazptymwJ87mj2rixBJd6cgrPt/9MrqYCRbt6A41KIePI1LAhbsylDlQt+np
Xsnc5ULGV1r+u2vZvlygwHd9pFrIvRVolYu+I65ntFKYaL/9DYSHAacWw+N9feiVSZg/f5ZS1oI6
cOGr4MRqO3jXybYmNbGN9q0NbDwCaK32hDExdbeH5JYaOqP+8r1z2QCmFfqKHK/f44zNDujEhYpL
P7mN1tJRJycz3KQSFdGN90ta+H0fB63CECJGeKlV+rqBmVuNchnaAuV7gJaZVHP8f9yOyKwWJtSd
rbovxgILEZ/iuZavAhb+QoOfOvETGynPZnEmod56zz6fydaWMisnUAQ48wQan/TlsIAyPVrBqrwa
dgM7tiGbcHSAVPw4WU+M2qT2hzrAMa1DLQS2bq/oeJjsLRc729RSNj1k5lw4fHcNul/Ad7lfAToA
do4Xv3kHKBjOnhwN9xi2MAp31N9VXC+dbRrfCqtbPD/NT7BbhJ0fIvfsURMvRElM6IM3JMs1+RL1
744/7/2nF1BldNajd89zTHbjdxSDk/NKbQpszVcrYB4K3bxNGg3ku3+dblHiVaNamH/UCvkcHt0D
kdSqsXGeaEzXMRM9vyvHS6Aa6MSEPoiC/78ODJcY5ODMxDt16pPbGZzBYXbZLTxairaCYz8U6Us9
qRAK/CmagfEw/mgIYqEI8xrYOoArmDlFSlp99ZGLK8SbHAxAJ2csXuVqlUcfnnIlmzLNzpP/MEkp
b14d+cXEez2Lqtc00AXvNsGXFV9PkJYOK+Jua+R5y+g6+t6WVWxkYiiM7SArT2TqmHKS5F9j1e0J
/Zxyeb8m6b9tpFQpjHkVQqcnpnZOif2grh0zuxONd6Vf8GAuxpAHNa47fflB1N7+s8xwMPgDetLy
2JyQutEz8YVtZ7vcy7aN6mhM0ZXMgkAIJ4eo4Mzd9PaeWV5RMHKOcX2wGhE1C3s2vg/2QSLdiVPJ
8lFzyJWhRt28Q6q8Acj4wjxOXm868q06l8tY/3I8A6X6enBEJelXXEswiw8+lbROWhS11StpAbiC
OxpYlTA5DwojyQzd359qQRtOlFOK6L3QvKSFQ17uEDdtU/l0T7inmLQ/kK5G8QYQmH+ybRb6cIPu
XKLcS8O1nIZrAQzjnis4gzoSBqh3joLoqxuWHVPRnRkb+EKNQexpJAyIRop0EHSTOX4VfAhkgQm/
gzvxlC2e0WW0J1ekXytPx9YIdtOnJT+jXTzsFxe9etDizl09N2jK2vh0Vbo/2P1+CNwcIcJEwhYY
VokgBUvEGElWLKah9X80z+tZ9wteVuQXcrMIFBRuxtO+N8eGZaDs3KsjK9000h8NXzB4HqgYzY8p
Svz6rmx5d+q7T9SVrxV0qGmOi96ny1YnHIJAnAn4eD28ka+G2fM38HZQ058LdkR1JKLnwRLIGsFd
rbzyxvoKjY4AtX5To0ybO1+DYeVMpg90IxwlYjf99EH2K5u/KjfXzb7z2n+2bJjhgjxPdiosWzkq
yaFJvNvF8t/jvLhWkXx06fK8ObL2JxFVATATEFawiIGipA8A5QjxhjovDrhDKQYjosPGWm6CZFSG
PytadWnqZc1pdxo3WLxUwg2X1gaFLdwKvGIDhQe2i66fNvy+8cCkqK0GaMnGmQduoLCfFQT16SRD
ApHemv0aQnruzwN7nOSKasDn9FWStUoIwC5I/+OGHH/d7OFRMI1NYUma/NDiTgSg9DaussrnLL+1
euR8IkXr8/9Q9DKGwgB+QuN1bPm949mkfA4In8bz6KmnPtYqjmSa/CfYNm9P+QOVb3yQKuTL6+SI
+gX67gUKCb9sZgVKfed0aahM9w+6QrkRPsmpwEOTgt1JbjVIDgqXxlY3srsTGslEBxx08PF1zZU1
TFH/0DaW6YigMeoAP+SN91Gkr317zrt0bHqsFNjpXnJUhfSeziaT2eJ2Kv7yhUaduICZ+YjB96SK
KTN0tSq5wIIu8lSlJpNI+sxl+tC7RfFX9N1KVjpR1MBUTKQpg2WNLlbWQnfGDA2B5FFu0VbCX1qF
I+OJyXA/wqUv2OeCRZE+sWdK/5m1fcLQFqWn2YT5p9c7pfyvBVchyPMkurvCoKwYtRaodm2UUw+n
4mTB5uL07xrYNA4uIjM8cXa4UZ7z8zzRl/YG30UY1A2bt62fSN/8izWJ9pp6Lk9SNO/F0fLunknO
4va4J3JAk/IqB5IN/N+UenuvUylQvk5yz4mmRb590Dxz+VjqgX62wvgnNL6436Be7gNHTv5bNaOe
O44cHa/hlEHKOc3N49igOAxh6yVZUusQQADw78/z/TTruIj9lwoahc8KvZuCFxsWaFebh0qmHcLZ
510HsY7j/6OcVoIIiFc4bt0ASHvPrPTedPCnClDXChETW9kXrsw+nM9CM0ydtt4T7TKhH2/zeUoD
0Iky1VkugxqUoRJR/WzBNs9CV1pUwJqYjOfKTbXN+scezjORctiYeFCcyyWQ6HbIT87ycg7+5cU5
2i+n+CgYLREVr/YCAaUluJVUDciDDGyZe/IIkZ6R2jhG6BBv6DvpvJEJySnyRVSpkc/NzL+TBcos
jJw9AOe+VjVaCmqNaAvwcp1LKncH4NW8sgMUkOEmn2Amwij4X8+2IowYsMtBjjzoOW5fUQG27/jF
iy54CSn151sqodkB5W/qcoII+/rwyzHKd7HGpJnICsyvxOxiz00Wm+x4LZkzcJYRYwYMEV1UlUP2
1m7D1ZR10T/jW53c56EKaMIpl5MTa0tNlAEE3Xs6JIdbWecqU3EMsIn83L6tgt4B8q7XTbSBp5D9
o0RonrZLVWE9IN06UuzzvFJx5TOQeOF/NMyl1g4Yc+xPvZilIyJ8b7WuwTD3hTGXlVEAw9p+WQsJ
jfxOVP6ne+K22XJuheBoGxoW56x+AvPnfJyCgqv4PDQWk5h7AxD4igu3nyLzYD+tdVmpFiUNH0Hh
ZEAd1BMaf+lZ6ViLeQ+lc+8CKA4mSrdkdTp9PgQnxNYB0F5R3IVvJnzZKbpE3c3MGTOIPf7cFK0H
S6+DJgCCnHX5AdVEwTwdxVJU6EJzRzO5bmunl3NccKhkYZX+Yzf/yRbASz1bzH2ZNcoUoa08W63b
f4YvmAtNhh01qBP5Po4met+e8vsT1rlv8Pt6WuWltGDT43ugyzFPRIgB7ieFaR7pCqHc48I111k2
j7J+4y7ySfRYdScFlgOcz0ius8omrGQO/BIhUYn3ARS2khZh1S3hrBR3E9LyPJSDcGgNdPHs/afm
v64Wv6JsMVFElbbHdzGVFrZgxnZgsLSFGNuaiKMn3Xnx9fO+0FvDYlXUSEYF5MWqzCQUglVzm1tD
w0wYNTtlpis5LaaBFPbuPRUyI1XmCgUMV7ZC00IsMHj4WV5u6CNYWB8yMTd46pumptx6bScdAaQ7
UnfOOUodRZmo955nFo5pDvoJV5ykuZ9OBkAcx/42n1wOaokCHqBE0KcSDdbYr5OTGZqQZom6+IKy
7fYCaxChSOQcQA5kukLdjQISwGa4fDz3y6ZybFdp5AL9SIpvbqDGSW4ftIL/egG07IdQLyGLP1IK
t+xRtGu1d6qxLfTcStfeMAekpy2H9E8jaWNQyoMvwdFzCisjwhr9ugqrLuWBdr3c6G3vVB5h9s29
fHPKGea9ek5SzaP6weASqWA7CNxvSYhjdQn0SY0KhRSVhIvdlQ/y46mwOhAWMeyvp3135pnXCrpS
6XMJgdaNaEft2BHxuHcbpZOJ75jpiMd1lcso1sbknqu8uKDcGwgpGcB49C/z+/j2rEi11I6Y0GxO
0/DxiL4C2oZrEVqLyJDEt1SBL6W4MFiep5AC+dOcJOYljCk/thL+q6WmdEe8w+k6q52Kk4rK8KDU
h6A3mIPhQxALv06amX9HFvJR72DMDpyuv7wx4lmjrN9PNpql1G8jXgxBU27KvCKiEZyG13iBpuhZ
wAoVed2mrKKhcX7vl8qmY7+GXyNz9Ryjc+pNK4m8lePduL+QcC9B/yjiUZunI/w2I6Mf8IgzAzA8
XcVxbquzi7VpGQkrMccl7wNagaptB/dimCox/S9uM8aPBL0uzHZxHGCrcoRPW0x6FOrCGKS4SAi7
SuOHdVd9jIU35AKUjQHI3dgvSeh0wA3WjkL4Mm4LV2kOy5GNjYkIZxvBjIkZtXhuJZ92HKaCZkJU
Xw3Y/+nVsRGXsQs21mKZrkqwvL8XAnQXq9VtdwmlbESZasCjaDkVdgoTNd8O67z5KyVk8ZTWN4QW
f/AugxI0ESh6proXOOPdABdeZsK65exRv13DI4hVBnoWcV4eZZeTvsnpGGE7zrmtAi5a/8kPoP9K
21aOCI1aUtf7qpclTFEPqLTTlMFqMsjMxiXCIz3l/vFXMKefouB0tdcywET3VyruJT5M51RYlwHl
+4AqJiSEgXNKcduXwtW8OuwWQ7/BAOWpNyNnSLScmUS3mjrP/WB8cvd4e74GibuOLAyLZHuzebeE
OCQVdeQ+vMvICETKXCB9kWosd1T3JOAuzdb+QH1JQzu+Elu4PrQcZh+0gM7OJaA2nmMDmLPi40db
PHun4yGxiSKC7MZoVvpod+YZJsXOK7LdaFRFj79H3WSP1uDXKVYT/EUF6efon/gfEvkQ9kHZy07t
COnBULzqbT2OU5yBBLrnZ4vdcksqWkteC6mtasJbAwmDVgzX3QHk+nAjpqYYy17ZMQp0hAoSx7cd
unBemDZ4cRowdbsdr8s+KRbNtwVQEyq7rCckgHtMXGVgx7SbBnGKnCBvrCG74ardK7RtvVobOvBe
0/N7OzpMqGrLEwxaQ9nyF0liAaB0Gx69vnbcSh+BBUongAB6Vqfkiz6zfSdk+f/OBZ83Wr8Bpyon
eFEswS5ZqFTalo6GCPRIBztkwpUWCvuTqZ0O6j4RT7My36/zIn7WRhqtNTCSiLDil9bQNc/U6NTf
Ej/GcmtAFp3lCl81BTRSqj7E5Hchfo2fLgcroH/9Tp94q99knuMCLSLCL4KdAwCgUV1CvlcB21oH
3IBwBkQ/CikfziTwM3dOyJL5XIOxjE3z12UUdqMbTdVEZFJyJNmKeZxjTRO9DlFTZZN5BSxhgMYu
X8jJxH6nivWc+4SX8aTGpbfplBvnrnpqcV73H576VL1qmTzbLs/7M9arzn2GwbLXuwDjzhAtF9sx
+yWR/6qdcZZDVxYRiHc920v0GIm9iuHnKv7pCAW0OslOnsCFB8v8OSCfEcQLTNskCaMIbw4ArhrY
ZkugebgZtCJVLTth6Ber4mDoYDVEATSigT9b+fWmmaLD6rHXZ1zKDneF8L+4UWK6dwUqHnRgMbfD
bF0y3MbKJ9RSdgGKsqraYnyMDmQYd0AtRtQWSASKv0pynFBe7oJ++a3T77G/2voRjC8RzgLh9bdO
cqMD29hmaKDKFHMxVihqEXTSF4MDxbCdc2QecD61yKweNysm3OST8Bz9Dp29kyJrSWP95XLINyLE
nkDZ6mqI9yv+N/V6IQ/lmeoDfOzmPrl1HrpaPoCTKMWTOOSSKkqId6xV0noY0O2OKcQpK/VsgyMJ
r42x2IaPD+rS9/2AXnvGDbHfEE/hZQUoVbtq342mz+jDoKbVMIYa2gzngIXH4q9Map3YWvvCOSxK
Rf3cqh+TfNXv9X/CVdQMptFt70IQaFLUf5Dlsc3jhwzqilCS8dHyui3fIjBvXG4CDHYNN9qzkSI1
5ATi/RHAQTX6yJP4tFByfcahgeDQigd/gfhcmKzjXNmQs2pYVlSesKh1J8fQy2zzD++tXrywJcxI
qL1S8aAdSI/+VEvQhKEGFFgA4eXa0ABhkKYrJ2+WfeobTwoRqwC0sEeOo9yPM9Uf92JjZB3tNT3h
TuLlKzIlK/a/C7YG49a7atrtUGp3N2eZWu05MG2PwKVi7PVoVaCqU1+giwPLpJIEwRDaSya45hTM
NMhulWBQoApfABKKRDlrA9XkChqyFHd7CL1Um1rtqrYHMnkLjdkpcUcET78bsfx2iJRyiz/pZVSR
RRw/43I71tqAerif1PMB6AmMd23+cbk3z0DBk5XuglFEqcvioQ3AY590duhrUBRtw+lNNVf3Dmln
4pSZ1RJgg4vQQyXn8ApxbBwqK+zkUt5LZhMSkb1zbT424PB3obYTOMLVyuZx9TTnhX64B46W5ZRL
EF8bB3aykkA9MsYJjJjtl1Wv92IHHX1wt8Rn7/YuZyGWFC1oRvpVgekvwAOgQOeFQ21+DaMuCiK4
YlFRFPZjlWNc8BJ7KY+85CKAljm7jhOlhPyd5tOElIMUG+CfkT3XnQotFKyWCrRxWDuhdb4XdLsH
8FDh3cwyni6SOsDomqlL6SQ8h6cfNzozUC/QEIwjQILhgHByb0rmuPwJ1ANkfj9ETaC3Hnk1h7Gr
ZFM5rakuYG89NAF4rnQmkk3fC/8e98eTXyeLFdz9edwpkTcSdBVP+HIkC4qgPmkvS4iYqgFiAsU5
aoORENQjGMPkfImPC740tFeyI8Za6WiN2tdpiHtoduCvJBeb8Vdq6OWkypRlsTZ6EPqBYPOuQy8L
acXZCLE8vCqn5uI0dQVWgciDeN/8FPpbcGI+DHW1Bbf2/1OUa5GKTF768rMHMnO/lV7gT13HTZWR
Bf+vXcRIl1fKlVTRJ66pRxlEQs6sJCcXkcP4vHjLOiWW7G6XdGuSrfhM89vfQ8WqTLRrbk5uB1f0
cZIKE1A0h2J6PYcCj3RLW9oCIxvsly+wweagkV+VmTXuoyD2bq5KipJSbQHIrwJtY0J70roNXP09
DiY8dH/eIkWVaizo7+sw3dTxGq7ka/lvk3jiyNMA79+CtrD3bciLL91ZWPLpKx0zkmTIWKt3fZzO
hyDFt3WjFd41l2xobH4oICoWkFni9TA8nDHjy8aR9RPO/03Z5WIPcZdKumGBB+UDj8aWZPFeQsav
Ms9P6tHzoyd+mH645l0qHBAW5yH/f6frXMX7nJuyXaVLTR6uLCo6F1lzklCYE4/1UMgOGXHejMDI
jyyDe7vxO4Tx2q/k0RJtw3pyLZ7ZRfcJUO6agiPoDDjIz1nZ23q43Lf83Y7XPZZoccegfLVwNO1K
XV2fztl8U41QCnJSrpxXV95xyzcRyk+hxiwMyktWa6XE2ZYjoQKSAZlC3JyyZm+Drq2+2Fdb35mY
OzMn1IW/EzMvCoFBpmBI9krJeFWv/aCmVBvbjqxnO5bLj8IO6Srj3CO4B92jHC+xbqZlcZZKR+lS
QJ2ZHz1GrjcMXLX8bTvD233M1wUX7LTgzv2DoSW+oIAqrt8nKMYaFFoAgLX2ISy5wxRmHq8AE/+k
O37O3ciHDHBtoLcuFfWnk1k/4yrhGM6mnGafQPgTt13JvJrOGqfsqQnE+cfqDS0Niqc6bLbuoZAt
3Zbn2woEekP4QmBE2QDjwXXizeSCsLmx/m/eA7GoD6T5ErkDTjsOs/Ii8BAdZCm3c2EGUxNBkV3a
AaMB4xVKOV66M9caco9H2/Io4IySxLY22PKEvkuCR61dDAmKGY9CfbPNSqKp06sf03tl5JKupwiE
Kyl8PeBEB1r+ECX3XFXiUBft+zaX1xGxcyB6YTJHnmhWvsfwRcAXGKib0e1SreO54IQmXXGxELPK
nznZNvOfv3UNlhJkVgC5CPJsuwTybiVCRSd5mM3KIjr3EjQJsa5fBXsVSdOkhiPC6MuN0a9195UW
uaho8/rsorFPyoddEBN9ok5XjRh+9kZMmE7jldrSO/mLIaIWxvXG1a6BwXeGsSalhoPkSqQOw+1X
9YAuLgBdiSWxicjGvZmuOBfqGKnWVmVTbXcjMpUOXfjXlLnUs8ByNkjN8NiFp/K3RxVP5oyNTOOI
jvou4VoZsH2zdFLdeR7VSvjo6WJVEdBUhUQLXLAB+nWXym+TlsfmDdTtRYVX/RE8ZC7BWyoQfegn
+GdMPxLF4FLglOLN+/2bB9TSlMZUTNcm4muAwlhwlEKOQf+uhXBHc/UlE0W+IljLrjFMbesNNdp4
5c5oVy09EmbIjET5s6oN7PUcwNHaFPhSJNLbQsV6N2AqWSkh5kSch74ay4nLqwPI3Z4a8T/18ImT
triOxQy56c+jyGo6PPJbYYT4aPBJE0H7Ot1zeuHJb/M4HU++X7dhNj4Rbp8GEaZxUFPTg7Kstk7W
7mXOnQtfC/Hghp4j3OZF9GRGlEREyf8bITW31yXvnXeMqNNSS/PapOKg+5PRj3CyqXJyPzdeXkI4
FZvpaHiJGqFFdqbxySEOrxrBaUZpvf6UnIWl9wZFqLRW4v5zrycXd36sZpDO+LIuFQXW8dym5ujN
WP4pzTWRsRCVgbst6kdNuBsLgqTOsXxkicDzcMmWFtqMCYGw0u/mKMFX37AuttfExPLjGwoWDV58
ubEfQk2obCoqS2dmAuMhMRznQEGiI7NGpFGpM+mO6qoo4j6PLxIR1yKt9VxglPwGSSXi6hyW0vDa
oD3C7TCz0h9uzQPK47wb1piIeOYdEGEjY53FAsRHVQn4UwechxAGUtUZVi55MjThjp6O8/Qstld9
/Oz29f6gyGn3D3spIXRySOt+SCzreK+762PSZ4g6hKsxDYRk6QrSHnRanCU6MCV/NU8bdrY7RLvX
4Hh7UkVDG1dISday5QoSbCNZyHm9txXIz+x3fkhR9Yblxm9g0DvW2OOCY8DVOScQHU9TNAEor/tY
OZbzPBo1A/a0xai6gL/HfsCK138YZysD2Oopj6zoTmWDWx516iPKRYiDCDLMbHCco2ZlkdT4mRGs
Ria266gylTTGTJh9AvTIqvRLuf5oew9A4H1Ct7B692dQxnHAhzyS6NfYgnPFd3mlEr7bkq2ih3N8
f5riJ3r0gw/mdhH2uvA3maXJAUeHgxOo/h+r6SO2gCCNVwwC6zHaTG/f8NB7QkC7F8+2p5JqmWvg
V0o6eH4jiApxSIi1nieyFtv2N4pDQn4YQw1FSNr8//TmJrf/b5J5tFLYVP1AIgHxi+QjAKFxVkjo
4dtgEb6Hzdch4cF8Bu0Kpeq84kDTGno0dRw0zAtLuLfQY48CN0BaCCq3LST7vxvDQPFZrAcFApeL
8DtP9YXIOtLQf4a3zrniwPXbm1dZE0y2CZDZgwC57/CRi5mldt5wUjoLe+pHPz1ykBP2ofEgwdJS
NEim9nE62teTI9Mn68DS2jsXu96GVIzt2knvuWabi0FnbonYncl0KyU6MJ54GY+x/y+CqjqTU5QK
G1RToxsM3AHZCbD/XJXaWlX1kpmGT3U8pswDzYzO/8jBYJzO9B7JuunCSp4HE5ca0f+YHA3mxG0M
aYbfNFKAbPr64dLlDYgVqPTuAVGZA+ilbRfK4kY3U/YulsoqzD2OiyhxLiyZ3b4x+xQYX3CwZhf0
A1IcOSVYKkRfPT8H+hPnd4M65GBd60+et5tiWXONZ+5b7g2h4kjT2ipHUoMFxRBPptZ/9awqJv8R
7ogwpi69maXH48HZlIFCSVt7NdkX5QmXp7Kw9JBbEY20ULde20tga+Ix9ZFt82mDWrHmFvefMovV
UY3tr3JbUW+seHv1yTcuAZB07pl3NsHyeqg39dFZIe+giPr+TVBSgrkwgE30Dt0PP14FYNmltq4U
XqEuM+dx6oOLrZidiV44yr/GNheaSFClU0wosR3KUzkvyU1UNTom3yQm0P3olss6a4YMZ5m/LDdV
cpXZDprAVT8p8NiBMjG75okvvtpMVY0bswei9vBPk1o7SQxCY7//umwiIaznbZisWDpP5eQNTGUq
Q+n5BDQcolNWfPa5kjcalXwHhQYMETRJWcvgAUmlafMR6iFzRZTkVLcKLg5KCTP59tl0hY1uAwwu
vUwgimbyHK0YbllsS7PHsS0uG6e8zBlfYKqj9eB3cKOjCk+0l0ZB8kLEzC79u0bvcgBZqh5fx8/T
I78jYCNfbzw0HIsj2XpeR6oc2+s25QhI9bY8mH0Eed0nQkwbZ2Z/2SQpwdiql+ea9LEFCsiPKYQ8
N7Y69CphtxCCtKrgcU3TbAyUMP3d+oD3rpmLuZ+fKS902J+gh9jd42BzJsd9b4iNgEXIiEAf6Qw8
wyDx7ykEhoX7+yAxDr4rUJo3ESLnItzy1JTStHJuR9lf+Rh3EEnoweqYkaE5Xej5DWeWmA3DlRJi
BqVjM2srZw2RMaxTDQs9kTFyW235iHlnIAriiC9ZsdsiTg29weBx4JDv06jEI1L8xjgxpQTQsVmB
AW5mhshiG6gY5UJP8BFx77fp2M0QacM+yj3cD4wsjv2RuhmoU5gxtwDlZruedUoC6euKx4ty85Wv
Vob2hnIdmD2Duq1m3p0U3EMvMoofHRRy1GMxMilczDyFbGt8dYINu5WEIGjaVdu25dunrqubF8mo
4kTwZmhTYwe1g7d6fmH2q8gq1Q9gQoAMXneONKg/VPiy6uO9+xpvB/sLWk7PQi1m0QBuzik9lm9h
6hhblBWmH1rHo5emkT9sictbeGk3JmQhJKzrMeVT+AZ/O8tl/twMuQGpc3lvBAM/BV5xrOpjMkJ9
DrEygIfvMXF9dWslW5Y88aM2se4A8IP/di8WGPACsoLKw6WADukgZU4Hn13numD3/Ooorkkxzg6G
7GA+2JRpIFop6TfekMZ/7VfzK9rP1Kr8P1FwGm6nrVdUx/Cub5iYeeI//pi7l77dE7wh1sSNB6vu
5I/WZ1s9g7EwBf/EsKQ2acY1phm7ZhlzO5PrhDVUZDGq0sgenLP9mHGTZdNegLHjdim6VzrhMom9
dNpMPN5U3dgy1pEMQRuu3U0MLNt5Yf1wIpiOCbfm9mmkAzwjfByriKmFU3LHmiG52IQRPpB7fFlD
f4jNZLr5kqpnXYrZ7CkfoXhDlLe9shVplaDlPg1nYv0/kGqbi3YdEUDd/JnIKjIBTfseJmdwXiPt
q4g1VQ6dDgDw/HVUD7nrHGw1fdi/mMcH90lVqXaCbf9pghOq5YXg4rsQwdHLmbWJtjkATlJCV4wJ
as5yxywSBVSQr6U9y4xi4t5/ESfWsc4tyDlBJDmCL1SVODf8xuxhVP9qC5DWni+vFnENLMSPK8jw
FnkPXn1AUFWHeuE8Wx8clk4V4TdMM/x9xT3FEl7RnSNzHNlXZY/NbYRDb+Vn3c4O/xcE1TI2zBk2
mCBkCQIvNNIKcLI/dpGapRLkDV+YHbnGtNlmxJp+cCRh/ffCpYXgzRKPANt8uxcOEpqQZqrKtQx4
MMgJUOVgT4WNQGoBMztA5ateMXH9DITyohONJl+hFsr9kGn6JeYpyZ+8hBffCuIrVg4xAYCV+duW
KXWB/IMjrPF9S8ZZAwzrdCDijNwC1zzNCjKKGDpTRGtHq4weaoHw73gew1E9XtJhX6hlGgTwftV4
HepqiMyhQqhLZG2w1MrpXAAWSL8gzA9oIcsht4IZSrJktaCDo8TJhOHOze9Y2bKM8Eb2ctwoKt2X
wvS9auSn+4Ci65RHg3YNN+Jg5M2oxK/7sZLLK2aEl3u6zS7rKQwIkst3cOallcsubJ25FxaE2Tok
d3Cf8dBeiSnSC16MED9fj2HsbZrXTAQa4+OzgjGoKu7D8jJ9LSR9KORRmFT0LVEgNpsNRhOCHzJl
Vaxh89c+MWBm0PeeKCjleJFuYzXh6q1JmweFBWag4Aq0RjKotBkUZp8n46funM91UmpEJp4y7TFA
6NnfB456LFHIW/DUotkeUBGLIfj4178lyCmue9Kc98WNerMeCC56XBZgAwOB3fT8TiPSt2bfHVvS
KmQ5RttaoIOZ6BhCRZV3cGT3+2bL7YNxiTBdI2Za+iQIMnrtjox2rj8nhGXJvno/UhQYlvjgsQSv
TuZEqGjeC8jlcBGJyLH9A6n+WkvwuxIqaBx0/CRnKyfLJT3ijPWp+DXAUJznSHfjPSLMO5yTWqUI
mPXuyfI9CJJDslt0D1A63w8t7qLAeGZvZhqz5qVzLGI7RtwS0y/RTyPRtqa2gUcfMBFOF2F9P+ai
BPBZEXTosA8EMYhOeesdnWMsdEV0BX4LnsM9Ti0gKR0xAkM6TOUYwDLkEmKG7rW5oo902ul5ipUJ
7yNfosjqauEharJS+FcKqSEfbxwmrDT6or8Zaw9iT7zt1mGe9LwZmRQproxaXIVxm+DYS7t5Ik7D
cWEp7M1fHwvZpO2mI+xWricDJ4ngZBD+Co1jujR41RmvUeFHvkdJz7TyUm6CcH+sF/ahT2drs40C
f2v4SpK9tuxkv7XBftd9HP84Qn5QTWZ7rNtmlgnXyCqR7+7Sf3v18tqNns5n3BG6BDnxclpwvmZp
BlRNF9irOK73n57vCfMa0skRl9Mp+0r0LpJHq0mg2pnT//5d0NACjqK0cFLAc5mrAMJLvJf4aXRW
fPaTRRoFL8JH9rFzBKWXodmzNGP/ZViFOfyCm3rdW2hi2yEPdn9tRBCkfN1Wq7h6wdIUw8IfrKCI
5EHE+FFa4jDI+juAiamg2qAFFjv+M4W9RuZrl+aRYewl3bpU0AAuuJHs+AZPAgEWqy+LEoJMEjPX
2uEp3NUHJ02rQLE1oFRo4McU9WGJuCVqUpt4av9JuCvmjOePduvouusdZRvzrU7EDFDjo98vA3bs
yGRA1AsgDlNCFCkks6bARnF8X1t/IcWTZbEdnEL38FWc5lIySKhvpg+kVOEvilxYa9uqo71sYvTk
pjFox4TWkL/7VvG0WgZm2vOrw5GS29jqLjmeRDqHyLY98+/rE/5uksrADqNrS09Y8MO0ihYn767t
tb3+xGA2KhuLX9dBKfQPZBBolx/DGQf1EbeIpQtIUb8fZXVJsPJE+1NrGNeuW74SrVt6MsFSEIB+
f/gKOJaUxJ2Y7ewH1vTeszSRUn/gZrf20+h79aU+sskxhiY2q6YrLiV6GXo/OtNo1mGjlx2V+GHE
JQBGWtmlM0z2VvfMg+2o38pUQxBwbI1S/FKWC2xWzMLHxfzEasFL7vrWin29g4Rb0x06Drw0h+5d
Pe+TkgizGjqKIF5i1a0cuUeBgZdDLOXdPlq3aKUD61txR+QjN2wdaQGGl1fZKJDpP+NajrtZKs66
AQ7U1tI74bf2W8QpaGcd4imRK3r62t3QBa36B5PCMi73sQqVBOYczJLRJhNcJD2286d1+nhSkYui
y6ZTNbfsmJY+bkmc/gQxvGYV7GYqaVShEzpl4V8mR9wMgJBCS1Ogl00KPIgVXvQLUptgI3g90b/4
xJcwU+wyJ9hd/GiIh8I3TD8q5fMW1Q86S2cOHDDsHp3FBaZCIx6bjZpzcO0JcDknWZZBbe2BC5kK
3AWLbHMsITdbJ2/WAUXS8REcxGtfEA1qN2pRCV5XK4CYMnX5kLrqbWtZ1oWqSidYcTdpcjoiH/RX
fF4U/c2cYem8L4XE3G+Ttove2e3FwbgLHqMP6IaWUYymSGP2QtWTxD4aXzrkw2z6F6ITAbBCER3x
nFWwxzE9YzC89IAb1lX44K69oGtNXfgGD6w6ey6RxY9LNHHFzDjGfRrfCLgk7whYILljai5/ILoI
CYuaEudn9qd0WbIFhzVZni7gms0VyiKNcPPPYX6uphAZzQl31DhpmDEgMQWBoEkPMkq2W3/L+8uS
N1/djewcAGZR9Mo93LMQ1DBAf5DIlKfph0EmM8KOnITVwywbMXTCYTyztwdRd4Ugd/n8P7KB3nix
j6H5hXjaLxlmnMHpMTfl4bBbBtHdQVcX2PMff2qd91QKd7S7a7u7tGwtbkNBIuA0sgZcxHpKJIL8
6zpFlbf/s7B9rpXegU7v/r+Ex0Yz/n30Vu4Q9ttqlKAHlk/G2K6PE0QcrGsqu1zQ5+LCbGlz0UJZ
s7eh3rkJjKVDwdLtvN+KhF6Vek/4S4bxzNTsf5wW5gaFEorSdOhX5Mrxv5R4cgMYvXjHys9mrItA
3INpNk+YPEPBYYVJxiHQ9noG0NgaGg4tGc6rB62KqyknKKWiXlw4Vl0Y+FzKAR/wfuW9qKKx8Z1G
24I9bWnJzkOddaLNmEPqXgZvz8qUWwKHLbGNqqJGkOYJsP23Ii/GBaSVWElPfvtX6Ej8N/drmXb9
Lsfz8j2zB6Uw0usjB0dVFcr0QWgoWwlGGU8rPSFW/efcL1R9E/qHE/u2YQND6LOwpThqkHh3AmXv
9x9gjrT3QG1cSoWToy+67TrWZIjx9XEbNlYPPs5Zt4Iz/MHtia45itY5kSEelMe8+kwcMUvJ4gzJ
iYwRBP3MjprxhBR0T821AEWOfbkA84wYYHJHVjIDj+iO7cliJQORZdWoOMtAdRA7wCmAJM5kC51b
HKQbJMVR4HmzAxUJAh2TXUg7HPJ0fAF/az0g46uHvQoxNe9hkJMbZtPlLhAhvL+7tO9AjEv2pr4o
3tIw+SKpHMJdl2Ws0guCZF1i+YXpG3Igc4rg6fQZ+VogCaPVcNvp0XsQlbqLoOtN+CbbQlZmvyNF
Nh7cqm9uu7as2Ko2obMDtknpcymQ2jtifuuZyNVrPr6lgb343jf9lOEK2Y0fDy8YMec2apFlu+If
9qdFzz9fATJAzUMsqV8y4awbUdC13yq1LuiuGqPAgBXPcU43bPQxG89zl79NXE0o01kdTwFRGhP0
33EOJyxbvoxUGe/0uLsY3E5AwHL9BKNMK4hrbZ6jI2XLhOoqJrEpINN7HKiU0DdouDT1koVdH5ac
cNY6YI+qseDZmbH+Afe4TNWxn50tHIQLRvSKaV6Y+AdMZtJr9zedWW6mcHwL395eNajYXUpCCGqF
Ge6zU19iH65CE8BXM9jgYTIUCzdmd6qq7SOAqmL7VrKjmly6HZE+x+2II0niIEH1UEtStqOSH0lp
KB+aO0aQFlay81eDFPUWGgjmkVSvLkAR2maloUFFf9r3equZqx9+Sa8xylqqaFYv/O7/LCGvTeOG
xUEohokOQs2WzCewMVmta88DW5XVOlTocN3mNBUamLD98P61/g/yr7dRwu+M0cS4qP0ZzbTLwtEs
LfAzEUhbaR8+TecWcpHKLGDhyp/1+6taWpp06KsOexw8/z70pzfkrzLkdojpreAzurwk431v+m1L
6Vf9blEod0Nn6Dk+CRoNBi+BT/EnSLllygzxBZZtHGfJL73q66S4PsawtBI2CYGEnsdV/DEFMfcX
ZJVQXNpYY2tY6zlC1hDRen8GbBoLY7tkxybxPHG32Kvav7DalCCqskcJabJ3fK+bhPJHqzdAxIWW
XjvW/yyS5A8ii08djDH2TGmSw9G0Zoky4DcJDrBUpZt6hWOxrKw8txv3iv5ntvqZ6foxuwENdEY2
w36lc2jfsIQ+LXTb+ymXUgI/QG3qSeXBZKM54JS0qStpoJwW9DJwtjPUTRKJhx/cdZv50pdBnaPw
dOqRmaQRZqdjfJHLnSHRsYRqbfoab+72dfxEWpVIRQ0ttkJ0ngev7MzdD4D2w+cMho2TXCH7eFuX
r5KGJbzpJNut4ucQps8InCxjsubRN+MvM5bWs22E5CHBpdoFpBElO7lgWf3U8BrUo283+ukXKW5g
4KkwS2afficM7K+/XKB8UBvUOVe4yg087AUx0Zhk8qu1diVuMHJ/doYyRdfTjEwOfblOV4ykq5K9
0lqX+ebkltmGba0VkwDMx7C1kFY7sABCK2Ywv6iCD3M7f/0v8lB1BMxai6YWhVFzhiWbdYXGdZ8U
33/01yN0XQiuJMoxW2yAhkG3em9upD8wgF0zimMQl/e7CrOC2WNVqB84fmafgorBsDbViFJoZ/Qy
EPVoQ/FpZrJMuFBF2k3WVAw7loOblcHkW94fbRtXOam6XOoLKCK6NGIqNWprfZzUVidxyI1WpPDX
OShBWuz55RlgO47mvV2aRecC9hKSsBtURZ+VjIjvIU3uZYNxUsavbfVeTFxdCr7aOzex0+IRK14v
Y+waH37viclHVFjx6WA9ZSuEVANWCYeRHl7I9OlRmQg19zQtXQVlA3Q5228v4NstiRshLW0AWwC9
JE6XlHzs5g20JFZbv4k5U0BVdJuFUf8mRSFyTB+SrxLE44rfrgxJLqx/vEca9E0o+G2B51U9TVSH
uS15blyLs8Vly+lLa3cMs7Hgqnv0Jqhwi9Uv1nxtmN4YNpTukuCG5SYaf8eHDP7hM6rWZW1TA00Z
qe0tWk2mC1y+18FCtMxl1jZzTkTgdOdOBBfgmbzAZYPMruRvfD4v8CQt4ouyIbp8JZQyAaVzat7v
xYrlDxkteL+21FMoUXltqP7IhuppzbU1s5+TPxLixgTmOuUkgjk60AXk6e9TUH6OuTah4fvpce4U
VL3pO68Crkl9ubb1U9+R9+I42vfT5FAlErnlcLfgSmiE5veZ5ldNEAbSa2Q/3frbKuXIYK5y1P0g
J6Lj+Ut6dboghbCpvCHJTtoO1qWlbr5fnZCbVOQ/Yla57qoD2JRqYy+H+bSM6sNRgJBNRoeBfgws
65I9pftd2otTkbNwPVzf5O353wmiB2cRgnj/kahEeT4arYBa4sPmns0uD5yOkeOy907H9nGLV+4M
fdrVs4G60nOG1967Pr143O7q7BJLySFZE28PNdHY32rZ3ugucOQVrnebg7VFwohKHgtjGvqCWk89
6FUjyRzR6srYOBkVMKOfsJEMgsofe2+uFGR+hobD+gkLUJLXlJ0GmgwyfHe6X/dPWEI7BcHe4Nh+
jq/fXxEEw554ZufbtJzMt2Q/VyDwCRdUO3lZjGoWjFUd5BJKJu421FOZcWDUBxW6bf7suq5j7IE2
825Guiynj4ifUrHIidWdBHNtkddUWaVFJ7A7ChieGUGtc3ahqaq2N6LFaQ0zP6cFoyHJW3Kqu0ag
vHr6JmeOCDoesdqEg3sZlPLyJFeLrlM7yl+MdSB7/jEPVwPc9eephbrlDYhdaggcph9TumcTxP0A
XQP/vJpy6aAQaENFXT3QHiW+JqQYBnB2riQKwmdszXDZKsaZWY8q96mfvfw+5Ma9F9t/Am5HGrBG
/oK77kUCYHNxASFut6vs78cCgZP0WKbNhaYPBmyUfiCz6beoOP8SGxVbxHdswg7isVDhwSmBAePb
JzpGPmZHlwO+AeZGshJ2w73GDP+nDwbWi/XScu6oZGlKWxv0B5QYdKFrGV4tmtcNPZXswN0B7WfB
f+sb1D7WqhxdLpR5rmNcn5IB48nUqvIz6n5bX6ctN6MbG73g8fO/f28e1JskNsB5443yYGHJ/P6r
t9vfsr+uTouVv5idCkYlwL/uqztIX4FR879TGPjPEbRqKMHUHpIPM2zJpSQ9alqmNSyuwOhPDzJt
vxBgtlKxETfo6gZAbnif6oRb6g4viFymZ5UN/fOBw83H/XdHL803lMA/3Fot9QMJpHldIc+hZbK1
kOKurnUH5LLbDkgjl6rA5Sx090qWuW9204NplkPx74CT2LnVFiHIjS15JsglOLeMsJI64RBY5pTS
QX2NEH1qNH5cYmtfeMTE6BJMesNzzp1gJZDSzZ3PgjtJq/Mwe/afVBl3TF+vAPQf08XiejPIK7XN
e/JG5wj8bMna/nNVhjRqY/pObd2WQjHzxOOzF93gc5HO8xQooe9Q7xR6BJWvvxa6mv0HZUAEiY6Q
feEa/C0terB/SDhcn0cfI3M3Lgyob7i03pQFagn4yxfrgEoynQ/XerFAQlPE9OOBR0y11qwpqxRr
/VQk3gWjhUMQK3VQIsyPo4GXSyl7+7PoOub7xhvHyFMz+fMToqH3or8IQLjLVq2nhcWa6Bh7BFWy
VaRQsFpP0xQcSfvWK5Lt6uRzg/yZQdgFZPTT240aTF5FHs90s5SQZ+RRhtSFuECGuZsvO4+lx9nx
iwff5/S4fiZO0z3Y30t9u8knUsXHo896tjRIKjRTC0YPbLJw3d+4V4AEP/1HlqagelsF152Y5nl5
GuheFZNvZGJYKogXqRALHexZ6uO6rTWQiOITswqTyf4wArQiC5tJmWENDFu0yWqxL/Ls9kVHd757
HwXBbYRxWUgAn+kSKjZoCo6Bt+So/atZRIqacLcydj2gmdOJswRD5weFeFEnHlQZYY49cCE0Wb+r
JSx2iX9ONGGaZ6sR9XsVn+RsRXXpR+RCYHD7wIkvpQPdoxq/OyaHDeT8lg5IlLQkmyqQagxr+964
gWHKR6d78dvmY9pr/u0y2rNe1Qr1srkGw6WAuGcWbomrrUHoCsbChqePCpVwLTy+BqwB+nb2L6Km
BbZrYx9XYm1J3MLx3rrraMt5qKDCCY1y6/YaUZ1Yrl+8TYN+QtAJiQ4Iqv61Efcg5VQiXP/dNrhj
AlRKlPHO2KSyGfC7VYDtrWNT0f7yFqUvRm4AcnBYNwMz9/JuBD9oGOvtZDfGcxSmrNanMSPcGEYb
7hUbeHqY8jozwhTyKV4zkUhq5pUbLCZvEbntEVA64GeRR0K744FUjI6pD9hA9gMzLz2GbKW75Mk3
PAJBMhSto2C5qXj3+3zEO6oqU5tLXj/SC3WE5VzjJkvaIXb+Oe8GKz7y6d++SBLdGoDDPMyD8EGK
bUGS70vMMdfM1Eluh+qPzh5aBQBAUUVtdegs2cMPoKan8ak+kArDRHsc7bw8FYRdKm8GNVvVuu2D
lOWpPfd2BflIx2Ps4QauUmeK6hPmBeeCj28idtRzSKa2Qwgs3s7mcj9UUprLQkk+SBi5TkcpEXs1
zf7vVWMFPQM8YxQAaAEE/jHViYvYDng0+BmjGozPEtVcC6FOWYGvnfRBNwaAaEUnxotMiFz35B4T
IV/mqgYZwN9Zaf3UOGkA2/K/1/mShpvlZKtYDwkHMiOBbmaYliGMnFdez8WRCHjbf+veZRnmVtcc
ORZugPBh5Vo6sw0dwTEzmU5LrOPaOuciwvgGT20Rs7Un4OvrRhbG/fTGK6Da/z+RKTk4Xor67T5k
I6J6nZMfTGcXTA9L4aYdDXox2wnKRNfs4r2r5QTrqFsSCn04VBs3gk3ji3kEC6AuQeIf7753hpB+
nnr6/K1WQj2tNFUOprNa0PeL+032acW/li9GcDBj74+N/13Wr8Thv6o/ge5pUOjRb3xHGhAFfliS
jf9mHtfoSzz2IqgM1igi/VNuda4nK42bRimqMUXidokcGPpgacNvHRdcWJQi3z9E00Bl4xCL3HVA
t/QnKsR5ol1U6GTRJXSiFUvCh6N/BKe4WwCtemQoXmmhpsGAEQh1Fy5/IpTplRVEkZlzPorLVeYc
A95DJklgtbwCeT2fueboij3FiWdiouBkDn5b7v6eKjYvX6Yi4nO1JYH+qbiJBXzrkjr9r7pPleLD
+a9DOdsci3OGXKfh56sFZbn75QXUrzJ6X3i7nQlrbb4s+trr62qFX9sf+QhhM0ohTEhvzjt0CMMI
lba6JOXWv0F/7brE8wSqf4V4ixm0H/ME4QSqSUvs5iYqCEVLGgoqN+g1mawwocKTRndxAFBr0Jub
YNm9xer9KVZ3oLf0EqCwM9oQ1ILi1WC71O0HwevIFWp3Cy4P9T754I1Q5QEtV4jEiztyPD4zwN40
al9Rd2oZMYpriA76v+HB6gENJ+FSkbhgJnILt1+TpcVfh0MSzmKWQCSuUGLP4b3bbG7jZr2/+4aH
/rECsikuDjwITgcNRqOsn4ecdqk9VZ8BBiJE8g2HIcw+QSM+zPI/tpJ8wmlXcgRTpB8nTQdftfIQ
2vSUHw083MsNFfHKL39JYGBwiii+bwa+dx3OzWRPUcJCaUGc000mZ4PDnR2K4SrwQNf5cFbe7xwq
uO+7qYyeazG6cKQOQfLf3ZxSV7xg74DkD8rvS9hVeU3/L5QS49YucL0mVfElIOqano0IrBP7r8mO
v3ANhhW150mjIsvsM8OLOM3LT707IIw++gvsx7KbITowwvtxr6qu6ePeRbcHFuyA9Q3ZrHpAS/ck
u9HcXDRwxQ8mJwZh7i59vWKr5JH8PVLilPmi0uEe483i9nAE43z95X6vsGUpIuimi+PImfj1ZV39
Bku39p4WXovKEmahk2aFdUsxxsM4ZqXwgODTrjwDoI7e0ZJJgYBwWiGoM3nFrtWQxwjFYbFpvwiL
0LCJJ/dHlEdS3OX6rsBoBV6LST+IAltljWikHvDegHYCO2vES1PyUJYR3bFJToctQPApv/SjUZ11
dBWj0DYEEb0EcSz9O9IocEzmKgSqldbnzX4z/9Rh9EMFSYn42+caxDoZxEvnT3DR5q24a4KvuFhc
N731F/ZYPLMjP53TszV28uUk35NsPjsTfrhOdP6sUCAL3MnexIjiTaYfr9PJU50vB8q/IK/HhKek
yIDrm0mqeMJC5h1Laq9acxMix5aoIbLFRHMUR2UJI2bLVI0hOv0XUqd27z/7PrDGuaothOljGMuy
JIhCZ5srjAzT2IwDJYDceNv9w5w7HQ/jnnmHbI4kG0B5bkjJLW6HwppK/SCgxXr2ID4OqpJoC3a+
mFMQFO81qFg10vXteaRL/kV5UGSygnR7+eP3jA8f3fa39pTw8+0y/mYf6t3CYdHjv9nOzsF4nl01
DtUOXXtSWG45ZxRr9tWRrS9kih+fNcJWP9WGOzzZXPFEVmpKAXu1l64fV+3w4FaySYJovNCXtl0O
wPC5omM5lgDxWccgmA5XX0subsfTFDdO3bm/sFPQO0mZderbauI+UBqoy7xhmf0LWsrqxIhThCnf
V+eLRYU5qtI/utnZi8nziMu2wl4SGPAPhtgFjdCJtPtJ1D0mT0yxK5CJU3FX3lgAdGsHh9CroDek
SofLpO1/Bb03xNeCmqei+IG94VQe1EkNQ0E6/9GM6liaLD3FA3bOxBnqBNe5EogwHaY0FykILDPV
IjnZu3VGvHRvTcgWwhu0UcVdsTAYgzDRSXXjEyf1NbUqG1OxkyF7gMvehDpUl1SqwZJtolAmiG5H
XKNiYneWAmn8LL2cLnrO1jSPofhzBfCjZeYgCREP+V4XMz2g3DdaCNyXLy8vwB2vRSeqYzBWKHDi
keEE4ZDZtjZb8WCxjCeQ+h4zLpzAD1F9C9Fbk39LmDoJeNCVRyW5YwdjZ6upn5w9WXIseMzBvQCB
Mc1zhsI0Wwhut3vWRdTul0GOYagIN7emJOxxNEDnVHNk/dfvsC+ggR9WIy9z9JhrZ/1SJITM58of
bCahXanrEFaZxJRpdnKqNacDV14XjZqBDhYsiwNQOfgh+J19FQOpbb4vmHZ3oKm8aVv7NpNxgXtr
OwQc4jUV9DKcFx2fo9MpXNwwgLzuBeFL84NwJcUASEjFgjisoQt+jrktHkz+oZ/3bb8thqvGcabG
mf90oeB9J8Xos1FPACEkdwP+xJKybT+x+CP3CHyC5IBhlIsCzr2P/Qusrdk4agZjqtMbjdl2blNW
OV9ephcZv3Er+o+kGYZbhf9poW8KJd6xih6rT7+5PtbAwLVtAkbK+DPW+vZydXOPAY+qfWrzMobS
8zi9IwY5zpvOjMbPOa14H8mBOOpdYt6s9NPF6+H3a6IMiYtTN0x27vaA9xTvv0OCzogm5W+ZoLQk
5Jxkyvw9++I8Bu1TWuByc8nQ7xsj8HAtF8ZHnesjmGUpkCuBN3vslGfxrnMM+I+o3VPt79I/QzEL
nXpCS51WRaH8nZE2Dctsm22uKldK4l5IteqyJgX3UY1fkfsX+ftOAmMewwMWwv9DUGmrElduamMx
d1ItBpcFA1qF5fIHMBtfVNZnm3hkkRmIYA7V3lH3g9dBHa4D3TnX+wJhyfgHtqpqmZ5WHyCHGQnK
pcAvqozNtt1dYbhtRIuLYHmSNr9udlu6jNKjBohImymxZealHS9UoktnwXRPma3tNVhw7s9LjDb2
HTqsY95pFs6AT+1Lw5QBNZirkwu2tQysnrMxFzAy0XKJA2lBTe1S70Hqt0X9nf4uLOIbTOtlw74s
lPqEzsgNSyienUFR+2T3+rFr92h/PR8DjcAuKny+1/zbbalrioZQKP6EWnZATvCpfx3pp2413hnh
BTA6dTiioW7ofgCFbc7xqPNPmHUsjRBPGK7BAvGt4d47gngFaXDipRzy59zQu6CBu8mzRlslQOYb
DBZM6slpdXx2bl/qOth59cN9xCM5Q1vl/JViVhJkEOl7aT4rvOF6chtsYNj77ZZ76QSh+JZlggog
CdbEv7b2hkkKRCqDUV7GuArb7cpxKh7UfIHSlCp1zR+F90ObsDSb7ymw0u3mSu5nexnuogg1rfoy
q7oA9rLfHiA9GE2GWuG2Oxm29SkWeNegwm/7DpJx33OKvt+2okMnnLhSuTHEYbXCpIKEze6A9ry6
xvpFHjUQhVge+nHl9c3aDwvY4MXD7nhT89FkgaAEAzJywnvYKCgnYdKm6G6q2lmOK6weUAr5eLeA
wgp2v8gHqZj861/yCn1KD7qdpSgHXW2jeG1/73uDI108KxfDgHuKHYRRlbihgkJpLSELxM1CEKRY
JJ6L15groBLTUe/kD5kLqsx/rNLC+YJu4N3unbY8m8preNLjp0iR/nY0bJ+bPSrbOpJ7euwZzqKP
4HhH3Gi4ib2eLw+A0esF4kmWKTPesHAARIC6DdKwI4AQUp+C8K1NORtIvhrv0qsqulT8UIM8+IIl
K+S/mtFj8hiLisfkpHjunqxwYXXsXvyDbqjzbevLoYD3KFdbVboafj86P661tjkisnPgUKCv9cxv
eqYBlWrzK19N+NLi/yXt18TA4XYF9ZoSEoHp9NAUH+uATOmhuBLO9k0zCbZYZZMZwLGRlZn8AhXC
a+oO5XxX54g4gg1xpp0UfWnrCwmGFec17miZw9EQ8tR7fGVDQPt9Z8+kX8sT2H63BSPn3G9Q6KGB
0+gf9OCEIVrh71mvTKJjoF9Xyp3UyManLejIZq2lY54JyKWKtC15ISotFRotL73+ao+X6Uto5fBs
00/uxYzR9G8OtfgKRzEjHEwiHeikJIFhRZTx2Gh8HbKWxNnZJ8SbH61ThrdjuacW0AqG85TNh3pg
5a3KuyO4AsBA2pOGM9VZaCBLBpOE36FKqwW2XvQsh5CHoE5lv/Guxr/ciLu47419pXjRkEVMXA/s
iwUYdXpr//5KsGD0RbcIIIAfYds9342NzRN5ORozodEKWdHkC0kAd9YWLzlL9COIx2/dAc2ZUYoX
mZckBo5vJO8dloIQb6osNslkbNxMCYtqpQDLxhpnv682n4kaJ9mUX7M3R1g/eqxhiCmc/5+nprqp
xHmhX+sBu5PnJIxIj5r8VjO3G+rZx8yX+5AiM44HZjAsQhzMtTGCQTHls6QjmvBy0pzvI1qCSv6p
qc78RF7pdFOnWvxbqXsCskwKeU4NpXXDSqaP9rCEE48tGUIMyYZQ41RP/hXG46oBQzp3oVdVFlLr
7YwhFd1SKu5ttonQw4NXLK7+9jEhpFTWhnvzcq98ElBBbSuDPWpkLAZLcFOS7L/KZscPYcCDwdRO
FIQPxe9akq6Qlq9t0rLELmgaKM9cCnJD4uhmt9wxY2GIjyzP9aHtCpByiJqro5mCHLVeerPsQOUr
ks95gP8Q23J1fK/lhIkQaSKLHciFr6Bk5qhQ1QABQRpz5P6a6Gaq65qVwiNs4Da2ehRfFV8OWf8F
4qLfi4Qzlxh/Szj2TTdy/HVhv4Ep0aMa8hbYGHYjSNCIaVwIkUuOf+7v5mKxAbtN4JJMvoN3rAgG
rClDWvCkp7xhs/wPGZ0B9shDOdiw8w2/14L1Nce8YF1Y6yqO/tv5c6agjmEzN7rD58KTU06aMzW0
3sUR6O0ARIxwitgUF2ipzcqsEqOj/ekpDN6hyNwBGAxRi4TrJb7da5vCpbw+VtVHqbUa/pHVQC8Z
E+Iv6lKsZq++hx0WX/iUrqLNzr4FagtcaTlOnjktcFntDV9lLVRqjl0RfS5fhRTT1g8tsUfckIi8
8r6JM3lx473IglJmnSwrtjxTKIh4zBAtWHpRwHCW6Ji9ArqTseVht1XlZy41o58zl6Z2glsh3gN0
01RbwU4qwWkmP6F9CQ8dePNcZMWrG53yiosiK/hHH/TzcWl3FUZ7TH3BNBEVSS5RMbaijXBA1zPO
G9DNlqCLSDSga7BaeSpZ148mf27I7b18hKGd92lEWu7X9h+RvtxE7K3QIG/p0fOyG8EovXiss3ER
pdS/snUNVzJHsacc1cJlxUJXsDjCyKv6W21frujnjdsbTWZWWCJzI+J5D2SrVSFTBkjg47lpvMum
aYIDnjowjM1KoZmxGFnYragQ04aIb0NQ0vVtY+YeiTZkSrpqAFCrZ8Nsn0/b1X+3O5tGLsma+J6J
4mALP48I+wJwxwmylc+u4etkff324kyqQWRi2HwK9qk4mtTsHIjjhWrZfueN1MVMO5MGvb3Sou1u
xMeFVNVONF//Ge6pKdCtn2/u8EP00+IdJAchY4iCBL65XLz9MBVwAhzzOC8nTKBrZ4dAM1+uxOs2
VZTW18WywkfJqGYEevEMgPcQk8vvBlLt465Ud+dwzqMl8R46oQpoOsgLPXosbUcJ7fLPXcM6Zd8G
L20xNlNAzeArxbh/DwJ3QJ5a7dMUJQ6T/2KDDUHAdCQJQXumGHTrCpT6RF/US/7BOvPSnT8elUco
oLoOdez+w12sK94rRN8WeY5+J7AroQ6o8LUAVTZcC5+lElMZoHeDYZPeDCDxTRrxU1iVfOOZuWI+
htYdpzrPkB4xk9KA6y3eTdl3ro398w5zuz/q6d88aSPY3NIFnQg4ybcyLDwdWtv6MQKCmhoWXzhD
QuAdPLoTi1knQeN96lqxUv0ldwiFbF+Y9KpzHUF5MSHDhXEJm8eftUNMDOBcmkKZrPoNWb248fHL
an3r5InvrpJnb5L7HBlVvor91e9dGaAtVe4K5Jom7Nb0qZZph2TU2E/LOclMYDvq+wOWZBGk4+mJ
3CAZpWutSzXNJRxPH9CB+NUWb9hPy68hvsTgtlywVOeWCWV5Oy/nD31HD0Hc87kwQJVvjEwM0qMi
6IV49Y4vqKLoR+eXDl37aYlQifx1LTj9q+LgRFsS0A0HnIlRE6ZgvS5aU9mEaBZ/YsSgLwSq2+J/
K2MOtjOpfKzWzBomdw26gOh6iuAXVA/UjY+38GB9m4Je1IPGO2ZYg1WNF9HZdFDttT3ke1ZGhaPY
+k7gHnW6g5YCTF9tUWzhv6zD3vnm6Pl/9mwlin8tW8q6yDMsdTCXbUW1xbU27X9oKM0E+fXjZXFu
RTHX6h6T4pW9jxPJbKCFsPfBv51Ioacq1EZ+WV789RIm4GjISxFSPmNRC/0GDRtA0iCyr7rMGPAc
tu2+4WPKDZ18jHIwAuJkUZL++fWePo0Lr2g10z2vjvdfYB1fcPtI5Etizy2hHEw70g/sr/NPwYUh
MJgLZ0t94kUs/V5nnDQqUCYFgonR5HKuol6XgiwzKK7IE3Hon8BbQ/b+xHshsupdUpLC3tm7c9eW
i0iN29oljnGNT3E360LhvrBYU2D00dRN0Rm0p3fXwRKYd2pDuKQSAsuOXahv8Igy7Qkcor1VNmGI
+glC2utzxALHW3yPUqi+hJWgEnjuKCFoPZTclb/39if7TaoXKWEVjBk0VfajVzqS99nVlp3/fZ0W
XlKvs5k2lQS6XhKUTKCOreQ2cJ7BEzaiYp6Lh01t4qpCiAvd/dNS1Ivi2ReY0WvQ/Ui4U1uRUazd
Z3XfAOu9ZTWetvR7Cpj4IruyYjivSPRJov21YffzWBngxfBdOGRAjEvii2w70xNJI5SDJBD92QOs
PvlKwdX5P66ywf+rG0ZHyqeA8IoQwMDOnzyzDTZHOYCrTbMwVf51kXP8ouHo8ZErvvIWljdomwm2
+fkAm6FQ3lozJwDfXn1c/3muKpm22TXo61dLCT5tj8oIErF/fJczUMuHVQKOzAmqXwShapTC8Vmb
Nbz2It5go15y0l05iV83ppmJwrVP9GNWvtcvn56kMH6qc917P+tjZU+7b8M7cJ29nP/XYAOnqOCg
GgCixcZl+bJseZ+o0aDBBy3Ms1eY8bB+rfMlDNmSyLLRwAB8BW3AWdqCT9+/F8kSnecFR929YfFU
H6II3F9EO8bCSfRPHCOef/0oES2i8JRYIVq6w6SCAtrOTblv9ZDd6VqXGl+pwxUtOEXroMnnuYrh
bl/YKw2T7hRD0bv630GEnjdZHpO7lgJki4p3OBuFvZeuVtt+Rii5TJzxf4dVvbZsPaaiQkkz4QSl
wBPpx8sKBOEfBd0kQ/58AUzUMRT+A1IexquWtiG6Yrkx9wsYo5AbRUBdkrpPbxP27Jz/csjb2jmy
T5dDC+BKoJQC5Q618hsX90giB41etxB6rn2vGLWnnkJXJ6IqRTi7k9vj5Ehv6clC4d2B2SczYws7
QjY6MxF2sMeAmo9bl5zBkJYjv7PAsIWjxmWJkmT1gxVThwGCg/6ckFCyuWAfyWzak6U3t/bm18bD
KrDtdB3wSB7TeIyBiHUYSlFMqwzMBL5lPqlE7k+GT87kORCGjHIJJ6y7eWtqsyqdFSBmjvPUKgE+
k8IUFYNqMLPwe99po7PWFHuHOVv3cUmhPjpZdrX9CZYM4Wd4RkJqlXW75BTp+nvEwL+5oJApnrLO
5ZUMviOBUSMqZXVuYdwwgXwOncfPpUwEAcOJmRy61S4MzfGC+3zcKH/ClYG+wIUSLGDLi3MeLYun
09ocVizF29OHG7Zen+Gcr9S8GJAnvJCkkSmqWZbypiMTGxeBjUtxe5SKHXIhbh5bJVtlNhvd/LSw
DV/II1HsS8TV/GaQ6qnEvFHnXZVmv6Mi+j1oQrB7fo2ZE6muVWcKh67heuLJz20H7qh6RtITzzUH
KkkRgXeQeq920GJ+ND0+Cq+YeZlLEtHNrM3ZGPQyAP5PmTYhMXSe1P1UMnPbl5sG0Ysf8ZyjNrJX
3fvY3mPtjaSoIfHAx+1sFMklE3Rq5XbwxXJNuDXif/eb7e00bHdmX8O2kSivpGbpDPue7wWZ0D6+
cQrplTB4sbJnigx/kPgIsaH89d4Qq2v0UIHx1gB7Lw8kiVFXaRi50t32NZA+mSxkZdqPEKsOr0lL
cxHyiOMQl7y/eZytvoJY4K6uSrUszhBgpmxqQNnTAvIL7qKIVVnAs2HS37wiOCJCccbg5hJtBeve
SGPJBNRux9g51bAer8bn5DcUEnIBgv1cpQMPooyUmVcuLFR5b8n/FiJ3fgUdQ0dofzSJrk/c7CHt
TPEOEkJ+/Fp8Z911EZaWbzNqEYyXrVKTArYdeBYW3ONDM4m/ady2DHZmPU+OLSthvEPe/PQ1lAcJ
hj/JC793cbZzckqns6eVG90aS38KQc8XCBBM9BXLMmrSngjjhD5V7Mu3cm0osBcTDLy4BzbxYiH3
xaazRRBVaPOGwwkFYY0G4JB6y1W4/jZN9ltIdHUTVpcHeXPi3z2nVsDpf5gw6i90HjeH3hLVPuYd
JiZQwTNOMmRMHfpksJWVglmjIDcF5D7l6SYTfC3w06xWUWnVfIgFeh80cxoOx3s8fgXv2Z3lh9Mj
ZBfGqooaWN5nnBAwmG8xi4LfLx7KvbIV/qbPnRhAWx4NwS6pd9a+gN3Kr7qGXuVUrqkptICsYisO
Wk0hPXDv958xQ9RP2tIH/uvcp3qkz9Yerhu4RoJuqLdSHEKV9dcblgKF+d1ke2coo3h1xs+lAMeh
uw68PO8C1JKKX10ncUEDIjkt9+Qj0Cnzii4OMJyFBvojocJ+3dGj93ewqRWRzZv07VgmyFGbKg6U
4Dt8TYTWQlOBIw4FIyzotUBkzk+sF2IdqHa5O7g+va9rmFvv0eD83d9RBKUKpK5jzW3k+OKX2WQW
uvFYKjC5BYfWc/WPamNnZEXaXNq1Wj9FADih8QjwF5dvpcAbHeNk5keXHSGMXweCTlKM/SEo/rPS
DKnMkH7O8KuxJPfsBtSNL4aWVtrSxR7r/5j3NLlYnSNz7tMk9IDn/e4w4DLppxGhUHpg2ErnHEqb
CMEoTiz3vNqPMyPreI3YCJv4ak9PZQevHxOrRhkDdVueYp+VxOscBMipFkTnBw5yHZ2IahT7UVim
NnOSN8I1RZeZ1RkTFdGCkJulPvZhKiHlYWqQcWi3XskztY5Hfapsno8R9Odv/HsI8UMtPetDBUtB
2rULuZzmSDGJbtCF/rQYQyoLUjdlYIr9sa2EOgu0zEeae/xFEHKV1GkZIbMiHjLBjtWg3PArxfHq
SMzh6BywcPZ094PPEZKxcaVxIYTQ6hPJku3UBRqWX7Ndv1CmRXeMEdlGh5MUepMDevcL9VVGbFay
v7VZdcAU/ZyD01E+25HX+oEK1PaFlf80lRTVZLFKudd23lIYBduLhE5F6IVTLEQsZpZPV6hcguBr
vmR1N/pBCgs87N6a0V4Z19iNDnP+Xy/BJvIK4C7WDnHk5qlWp690ODrO+ne0Vmfh3ssyxxLyxmqm
I/EvYgJJRvsPu75kw2q3sdTFPb3rXbC1LXlx/gmGACgkhXKen30X3H1rCPfJCKWnJghW8ZMfHqAz
ffpVnHBH0tM5bEwct57BiVwC82x7WrftH4QnzXXiRYIa3pzwK6BzA+2kFPcta9BViFplzJ4jOM8N
uPYlIz9bH8c8XXd42CajQIrmyeZDpB7AUQ4hMvXoq3HOntT9DVh+vDa5EUphv8+bJmC5S8iLWCua
lkJTycZ9ey4WmZYnEkYqtOxEWO5cdVxlbjC3zY8G9VQ7IBed+NrKGhQh1wYNZGUJkNutO2acRkwc
C920MXHWF2SBYBgVu5RMxTFDxJtHDsbvJfUrgZNScFGfgLRlK6RbSYq7BYep9cVijkqS7ZKKBnKZ
/+b+ncjItd64wYwqH3L7BfqaUZRz57ESYUNXNCIeGbLwreCwlqL/oLSWCtH4dg6LYCcvzM/gGif6
RHjLxXg5GfcpUBwwJNbX8JzTdICwn0e3ATNJ5SmKqmnVKYrK+/d7kM1ejFRnI1NTqqTL6MzAcoKQ
BjdfzrPob95fh+L7gYZ0A+UyXmWiOy/o6aher4wY2FYJpQmxvj1n0VTWeVEBRjXneV26hbQIfmdl
CI/+WBUelbP/O6VjSJ5JCB9MpYNeA0jS298ioiUC6yrzZl0EUo9dtBXSHCgcIfaDGwpelpv+gQrQ
TB7ZYIv2g3Evx6Di+KljB78y/uQD1eoSwXc/XdJaE9WVA/jZFS9MUXNnzbdHLdZ+LzruvZKXv0FQ
L0XVx/RpeqYtbjs46sQzab+OqNXcpHNrKC+tkEKPlxMVaOGqpALbzGBQbQAeLudYUl5Ibpbi5Eev
pPCdUSzJAzyYyD8DLfPye4KAAX7ASwVfCJequ5X03OGRUAUXei1EbRfmktULiO9mnJk1VuED/haQ
M8ZrJAbURTAkhtM8NnsaxEDRigi1LlEsL1jW0rbIpx0rH2FSViDQXi8xpCHl187YudkdLCG00tmL
c+P38bVO5vTle/TabWI8dP3+Uawx576mhNfqCtWZeWRD4Wtban7XVfMFKAzJBys37MX+1Nd7mYfI
gfKp34+yE2P7p634fFWSzW5wFkyHEhP7Bo4BEcNPH65L8uW0bg448O9MkDftVoCqdOAibP7cZJ/Y
xIt90vFTRMKQDok++QcA13h28W/m3M0txVXNnJw6XAwK6keUc8SZwhKO5qG9AE0xK6XmalbgQ9+S
U6TtVD17TybdKIuQS2Z+WvK2wGg4SXaShcnxcabuoB9kvxZnZawwAoeK5+Ox4aU8n3H/CiaGW2SF
9cTJCDhqGi7b91cK6eXnYGmTKjhZeziNas6F7bqt5WhDRwE/dsDCJlej/DDDXIX6sPPEbGcDpvB2
TnVuVgEo7hrYHnPnTVA4kVFMlWp4CxNFPZh3bc1x/E/XkM9Xdz6GPzBQJWHDe5+iebA2msFouvn0
VtyJ+8+ki5y6PRg+A5gOjQCVH7Nf3wuyXfWJuq14ME4WHugeDJqoH9eHymXDtThsVK7K/SzV8Zee
o9hIzODnqOYg3jDfg+PxLuQvcsaU6bEknxu/1c65og+alZLNNcxge4vt6dVbHNoD+uIBFtSz6OqZ
jmeLq27oVDdbQHQdzcdrshBn7OMHZZjFkPGivv4WlV+me0pdAhZ1GTR5E/pSDd3TOsjTbO+1DSgJ
kQzLBsS1CweQ3v8iU8BeqVbO/vV0SXguWNQ06sSSvv4SXCiK0h8WFAzccgsQWRGGlcSs8hP2aw1X
meYlQbfkCQQ9Z9At3FE9Jx8lF5CeNwVlVHq230I5jTDvHKxyXaRc/Aom4HrmKv66z2hrFcUUFU4e
m25u+XqZac23F/86KGN28nSwIp5HDFikyH783WtZHYUp/2WN1c/hEd4abdV1sF9bx9jOzKFytN0q
780RP1GfeZ9rdvIDfkESZiVowtNyGcoDPbJ9DWKKnTKg1Sx3Uc38QYyxzqV/DbKe+koePXxVsugy
/srr4a2JxD2Y1LADR1OqakmowuLFk6oGr2HJZHvN8Rh4tKTsUazmhvJvlFlOJCeKJvtgIEF+UVkd
9LEBZ9zrtdK9BoKz6WSqzojjCtn9Q0HLaXg48WRQ9ljWh/fRDO4L1H8hV5d2xzJmQLZqlhy7rvh5
o9dJ68BJa9ulno7vVHtsYbDPzsR5R8WR3VNpl++Duk2wavqmygom6DkJ0g80UY5tCjiIvUqLxVO4
CExfYSikwzuXoPRaXLHcj6xfZZpI2vcCB2M9UNqqk6t5HXGZa5GUuXz94KG1ZmvT59MXczCoQhop
jTNtj0DX8C4FAeCBhvMEwAcsgmRb4PLUad0LnHzghpDI9VyNjQbv6IWf1/gmsVZpLO3zlDmDBVwG
NrnU1jW5kT4u/3g3LouuWMbVdqKEnD/Ddz4C/j5D+kNZhlC9UwxtmwIce5E2ERA13aVBSKypQ38e
cYcN6nLCZCiwNvsset4RdcpS8gx7GUb6c8/iF1RbjPQUagjyHA3Co5bvh7ssVFTNlcSQfxnHuGHN
kQgYrG+ChuDAKolicUjjokANDusgfTC+ueh7aeOz0pKGrAh8qZv5rxe0DNpkpDi7WbKb35FWLyTL
k//NnYD3Y/63mWH5wUi6IOhdsBYL7RhvKDXb41wUdvA7QLuneJHEF6wBhd/uKZqsXyTwbVQn9BIU
YJsXNTfBpohQGsML7+G9XV9/UbeGCYw2FuRwi5w5MI2s+GrycGHjcq4ag0AWBmu0vaQLOtUsOYsk
d6LbS+5g1fuiDlum1KE1o6QlEpb6CGNmFoNHwUSWf68NMmIyKBXesB43YGBOPSkLCw6eGoZbKc1J
VAX3vs/0WiRjLiYqu74AGGMOa3Pv38FS1RR1E7CnBO6yt36bB9FvgDSTtNFCuth5yFGKVEsuum5T
of9O1Pg9gjVb4eybNqJ8OGEdhXsXXf/4zcMBHTzg1wJ6VmRw60Z6FoCL8gfLgoEaRdrG1z9WRAvh
j5g7GEvJ9p/zhAj63pNWnY60TChv154zGljs4tCokPNqCvgccJUm/5xFla4gPJG0PtxarLVvN5b8
85awYXkCjDVyxQ1oXcihQmi/k7OnWiFoP1hvBxVqqDPGc3BgJcyDiDwCudMAmqj6d+Nbr+/tIO9A
t7EWS0XTqlodzGos1JWB30BjbeLkxadVmePYPUJgyHwKH3JJbvWNEkEiRV7zpvRdN9bsxOs2afEN
wll6zCv61ajzyBAPSgaN7RgWBukzCVfDugJVSR7BATt4pfq+bmZUsNjngYJCCKkI27uESQQ0S7GS
VMhwVea0zNYPeMOybxKkotRz4FaDIcm9V2mxu/YchiQkoYEnFRbVUzpZg9q4+byUECgXpa340A+E
fcCOP+xd/DiNUTpfOV65ZwwNb7IhEHRM3TKRC5Rw28pMVCEpx5QdqvToRqBNdeTf40VANbv+OMgc
SlTN+MSS2GEGVSo8t+98SbBjiLkIWS2PNQvhsciK0hOqqqxpSutMSgQeNxOZorlGs3FygqBvqjz7
f82inL9RRGk9kzyyYVPxhEYuaSY1FIAc9nuesGatgXtLAPS8onM62rWSBe+eETrZk9AyTUOflel9
hV6L28xdqd4mGdP3qjtFhZ6iDDIAwfNPQPrkLzqv88VfJr8gLLBKFI2kqiESdccEqxKUJYerWs8F
sAJYeSHgsgSf30LCP5I72GvnmV4sqoG2dZy1otbAMiXBiphKKAjOHGJnTdfoSirQfABBU0cxGlBm
CmBNERxVVTbZk4jMBqECU8GsgvcqS8CKiCwTIukcobl9fhcMI+UyQFDRdv1vWsa1O8ylyYbC6E7M
4TQPe2uYYHycv4S6VvuMjr1Z/s1BN8VO9yad3IJUL4WYPFq1wN13K/Yt4pc9/bdF78WlCn9Tvbi7
/n9/2kISIGQhHnxcnBmkaHbq2Vb6Wesej1ypg6Nard/chPzWvrU5FrRNv2G/CDzxnIvzfXlLtHmE
kZYlc5DaMOK4A+tEHTIECTOZZAgFyVAMV8OiDuqnnvYOthpz6WlVm1eIbLG+TUjC9Ml7KLE3jmrX
JyvhjuQQz6zP1C4wz/G0RicIxTsIBGSttLq2PXBNRPZHsI+aYSuh+SlYQE6NxulQdr1N1kv/MXcc
Nf+/ficz1pu4IBiA0YRD2EmKbd9oOvkqhK8d/4NjuWII2lze6qXIpQ2eEC9tARSZKI8foyg1WzGN
A+7CX9eWy+JOnVt9IbH95u0LJ+SmOpnmEqAREYM+wgZd+779Xv3Ub6TBZgePfXyvDl6G5vtvGZ80
Kho/5lsNrUL6dX9NPcjziWQeAj/QPjVRgiaE3LmEh3/X0NyqkBO34PGHNLpRZRtT380PnL44C4rG
0+D8HSsMUncUH/FYKIitchqH6T16VK5VkrvwoJ6Sd002BoFH
`protect end_protected

