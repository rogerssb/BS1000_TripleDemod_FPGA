

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qQPuRISTa6yTV8jVnjDSkAIpWnmjwx3kjaC0UCjHjlxURWKOpytjCpREdB1AZ3k2rOuDKh1tFF8z
nITOmdZ+PA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
FhyfW0Ufa/XiVrqmx03BtroBYCuU/mp6sR3FpSaGqyKkZFDoDRM/ihUn1g7Mo5KFKFOSABJonGsN
ySOdGYVbpdRsg+OrUW3RdLHpdOFpZU8uDR68eu8kg0+zwNjbrsx0HbvIeLBtwr0KoQQhu2pBS4o7
mud2ji8nl0taVyBozi0=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BE2ncq3uF8tnDn8h9h5fHM742dMiNCfhsDawJ683Nw0yNiSjTQ+1d/6HbLM/tVbYYXmmcE4vOkkH
Q674koQDlJ8wgf5EsB3kCidNIx+3gkuVo5nM1zxATzpwZECCJXm83EQnDH0Lv6xY/E9Yu3j3QKGe
+7xamN1cUjgh1fWgZsM=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ud4BXsJG+kTHw65pOwWDRCb6uxLWdd9nVaHEr4rkDstKTWriaxV54Z5dRu1HvPL5yid3csZl5XFu
Dqt6IrmXo5DGMSE/fbJ3/tIWfsmL7VpEq18NRtSZf+NsiLguHJ1xMfSMr93PXkqN3FYvQTV2lx5R
Rh16G0TpvTTy17sU1sJYtmrI1AwLDEOv+ZF7K9m3CUqcSylWDzQSikoB0RarzW289igUg8+5Z31D
oqM3r0L7QkcYsnW57Aid2cLxQYI5RWvSsUrIJI1mGRNl6n0jKx921ScNSQMdLfe2+GECAtQDrVVM
gFAPQsUaNLZFH42qTJKd5YumFlRihpR2lJRYkg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
u57iRnJNC65201+394O6893mBhn/gX1DDYraiwctabLy3auAGT0lhkyBcSKHCVSBcnA97F7TrPv6
Vrw5DVlmCk0ORpBhXNgMCbU38+FMxsPE9rR0yV2mdTHXx8VB9E20hL599rFWWdRK/Hpy5y+/jNSk
FHs3zI9MPUzpQTUWQot8qn9ytAI/F34u54jpTCmeTrde726xdwGDLqSwa34CS4gq5jC2MvL4XbWn
5lrObExedvHU0nQuz55iOFW3deuwcJUptOVLu7xtao1T2SzCY+gEsIZD8cVv/IL3i4xjdgZAQmMT
k4olqiQEN+P/sz+tMSCknLWhaI5cPk8fxGQx9A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
N4ZPkdFwfTQ1lL432dKkSr0WfcgT2w+0TqO/8gZgriW7zwcrd/NY+iISaE1i9Fs7OFpmQrowLGQu
uH50L8dpIcahExL8zepWhTPy55u1DDTRe98Nx+AV/o6cN/RKUJ4o4sSAyVeu6SJaqLbMk3ZJKH0h
POekpClZIjwMygSY51H/hIoszQ1CirRsBoYpS2LnEpIBfX5zusKBh69V9rwpWTTku+HkO+vyeWaJ
Hifp22CiFzTBTyGscknns2X2jgjH+lpcgN4rGz9skAFqaRqb65f2HM80biITmgE3dh2UbVBu9Fck
wbHuIImn+BU8qZkUUBcLw1JPYKhdfQR6mfTk2A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296032)
`protect data_block
p9T/Jaz7l2Pn+KsLzMZb++eH5gHkyJE3ZQ6T2z2vb7Xlfpj93/yRqjvwFfpTDRdptFuG6AEmJO9P
B/xAXZU4rUFUJaL+cfUW4aEqha+e6JTJk8H4sg1g6PoTQ5fy9QMUTj12yeWOjuyXGwUDu/8j1cSs
XKhkmZooeRS2dpkQfa66+txMi/dN2X6u+jxWhlM0WWouSMiVnLTxHWgLEqhqIDmzYk0Tv/fUC23/
uJJS6qGI8L6F7sdIr2jf8iaVvvYbUnfhfQXlLG2njC7bFiwwPvzX/m+k8PsQvO2oQXuVqPBIGaay
7UaB5z+UQ+XMCujqo/yNgSLOHYmP9QGNe9XXNdSwvZUxRT2UoVxpQGiN/rrGFuf5/LGyH/H/Punr
XcLp+cCg6R4jFPhf8pWr3goqoyctGxeRdOoO31PHwB2DqCQYalIh/Ltmsm7btDoZ5pI0knqmvKfy
HX7qUQ/osFZvhziejnp4RkV5dIoKYKCTw5yK+2gPhauPX/3JXasAtn5CC4drp3SeBOXMYsp30z6j
XXVTFGOY1MDekVqQCWUa/ouqfvH9bKlvyFWLOm+pM/tYNmcEnHz9Xvia0vvQEI/GQ8Nj6z5mRShb
BV63tOqaOyIw1CL7dM7ElsxzCEaVBhxT7w7eVBk/aLiHa1TbbVZdAEWU7tqKCXzvn4Eewoad4Pyn
bO4ns6sDHfQ1L4Caavm2fn15i+USj493w6MxJJ6FDOPt/lCC6fxZJkbooIpzTZnLMZgOYRJLUmRq
Teg3TJX9Gf4ih6kbGvEQ4yPlpBr79ln7zQ5wR07O2MpKvKs/AAhzmbQDNB33Eto7rAn1OLRUBAa0
d6Zg4XJINGt7sCvXhoMpihx/afwBBhhTMpDpqlVg+PoZe6RfgGiwkksjhFcE+kU4gqn8cWB+PiV/
VdV+xaEWz2EvdM2u3I3ZZ9KPnmq2TkTo9eBnwSsybqbeY/KRxvDjChFCKDt6a7gTMqQS5lKN+eNX
CExixOd2JmjcKD8HerJk1uDsBj8Npl11YR6JnBUYc7Fg5A/iHSf0gxxjYQcT7E1n8gjEhBoUthmx
5NmcYjxwOneIzrx5mqoCqQnD4aaejFkGqJ0T1TxRqha5HCbGmPRrhG2lsgfWc0+wR8k720dpy2zv
aQkz/zpk6v/442vlyRM8GSWvDXBGBPvbt/2DkKWn3uURC/cPmssbydEGj0qT/WGlzkBhhnMAX5ir
aCoUwr2DeF28FDgneFIXxQDIZj7qXUwhje3tdcNFnHZ3Ufqw9wpYQNHr5v+/3ORCZOo8CqoEjnvn
VA2yfMEEZOqzhm0o8zKSPcVeblREXiu9B0VnfmSrJr1r3Sel6HE/Sy/YOIUfjNU33tULQ82EMf+J
pYeib+1e1EIwJXbNwnmhsah0OVR7PHYGSYOf335l1M4wRIVHiLKkLxB5oZ21KU2UuYQ430E2AwYo
dYHCip47Yp7bDRe5nvStZCVghfI++Z3IuCw5lp0gp2dLDSJcFZMY2qPvrvSnDyW5ALySsJZuWivu
aZCWenRWJi/maQJ7iUC4Novy7pcL2dw1dG908/1A0iq1zX177GqGGnBGxVmLUZnK1c1a0tD+1Ihs
EbQZinRPwaIQ/PDC2S5DguVIg0vnyXJw9belDf20o0yjQadSveX/CsULjjxfjPgwN0h2qe9IwXoQ
bTjAmu9x5AVGV+vjiB+qxeNcvwFbA2ju+L+i7vsHf2fDxagvGcNIAM0+4FHMstMflAffiFC433oZ
drcN5W6wmox+YkN7XnSYOCWTHggcR/oceFDN49HxVd5UMUSv2qzeyHhWkRlsYrbHrpIGFo6SjS/a
dWKK59qNwHKZVrYkYqOOO9u5BK8sfvF7usyx29HPPNPFcQmLobrHeWlm1g8d1KzB27jDwMsu/AVF
N5NekXjnmf0WB7PJ7wrWCNE7i0EqyyykGFlwaUTvesRae2y9kFKzwBfJbFs6kGIPuFHu+zaa2HFy
y670hKJZURPZD64jyYQJo7CdrjnY4I3vg10icMH6zZ9JYIfOV/eIFZFSXZBX1FxCMz2rspI9+ovF
fx8I2zV5e/5f7BduVMSChZR7ddjVxgRmTZcYNb9HsPlhxwJftmSxbxVHNF8TpS8+RHohdhOXtvNs
1vZDGg5jiBM0bP2eactDU/POFfx958soJOPPG3xtUT+PGnHDkI3eXsgsBDytM8RCLzEO6uaaqPun
aMjAzGSMafdQL/IR3kyNEHm6+OSp/4sinrNy3Ypf+SizMMYxJJAvMCItrCourbVtJ6Gc5RSfcGQO
eIEjcdbK0EYeh97NZTrK52mh4in7vTENLHrWCDWg4GyLtmtJZFNiyH485sdbgYKMPNwD/t/7AGzn
VpkMAEUT+pKdMBepG4QvBlCuV3/9QKIW2JGCX+EsK9sSS/EffSpfd62HxOuqQpmczV4Db2tyJRcY
9Et89zD2CaJCmy6/YZ4oKHC6OYztH714ZjbCxQoY5X0c0DduHCJPgLruEqUUNQd2GVEvSTRspHsc
SVPWYabjExSSLzwFNKOO6GjcunaaK3hm3psFjnjrsenbsKk1fv/y6hcy1ryuVIc+dK+T4+4QZjdp
NK6aAi/w9JF44e2FNYgxs3YlOizgPM4gPm5DBzPmqSW+Zu3qXv+wKTFqaP6LHcXca4nMxnDw6TfV
hGqYa8AEtMSy1xuFH2SLmcbEEK9n4kWXSc95AjwYBWYQloWu4isXMksNY2YlujpO8x08VxvsBWPm
QTlGW3jNNZ32lFVLyu/IyRTLLfEfaiMwPXxJWvr/ODyfA/lL5XOUsRyn7TXAduMxCfg7miguHFKt
zkHmsBoXQZPFN2MoZqleh/epLxOzFQmJs3kgfiT+BDqZOJ8fhRfnXYU4G5IAqoaQSIyj5GMcLta6
w4SfK0JJpwuY837PLgDKTgeo4NuNxRVk6bWYK9FTY3II6JMXC4OACSijY2HF771gRTJbOwpOs92t
TMaBN9arOHqssHDq0TzfB5Tv+6XnWrBrjbmsP8mbe7A3ftXV8vMmzGtkXGKqrsas2M/MIjGQWMoR
OSNbGwaNACfLE+9Krb491n0R3feief6MNc/m0m0Bl06/BrpHTjLwvA/xGVUT+aRPQS/I5RK1jWnl
O0uat9I+zqx6Q2RXvQogPw5LxWRPg5XRH1iwDVQT/53dz5kEzmPjJmZqwTaXYv1zpiJXcZK9yTDZ
1YUcuCFOkheEumI0ZD4awRfunXJLKA+v8thq4/TNXZ1VcCwfi/8EJHaSSe0055nt4OMJeXhdop+P
xciADdN9ml7tu0e+5SajFuicciKtbm+fehC3K7as3meIQ4LhkKv9XVC9vK1fN2B7+TYRG9153YXH
JiBoX7mWBJhxswp/Bt/zZK/xFcsqCa5HIV/TfbD/hOwWfgkD499o8Fwgvj9Z6qIRDfW33/Ozi9EW
m055h/DljlXZNS7sdgQrEwh7VGssC0+YXGjmyCcW/VJ3l0QpPeNMvMW9enPv4CribJzuKvcn5jrW
mfaMlhbkIcVLYEyYjis7brxjFdz2a31JjRFNvWZZK7AzSvzr38C/K6zHBr/Hoo/gzH0F89Nhk63z
VVvW9K8EbjXMFmiFhzRj3zMgqVvpkD61Z43a1QSFjRebnUh4nMMXjALF3v2yVdW20e5vpVqoS7aJ
9Q0+y2nLM83ZZRgOCnipT5rl1DWE1LIytCSwTW772HUb2Nook1OBVnrY+kYy1zOBJ1f4TufOpgXH
FTVFqwyTzf0X2e+qvXoTtzFnF3oYYYTuvx8NVropYxX7JGYRF/MyLUnzK60iv4Q1qC7jJb3uoulm
Wm9MF5mlipbVg/8SsCUBpav2qY5RPizjPtPq2n0VIj/Z4E+5BdxNzPjdVsWjf32vJB5NBCCB2y2w
C3Z0RqwTMvE0CenCfFstJoK7BptRpRxrZSChb9qYfQdVXjOYQYeGMA9VdiLEmOcjgF3RDbgVz4Yy
Dz+bG/J9qQvxDHsdw9NxezG0oDnO+/91pNfr/oLCjyiiAH/YUIFVhssVJmpZyxQKOnK+IWJxz70/
1sJvcSh/mDvPGwGeLP5RVzISaf/QvFa7KsOwAKWBNpB4Nx11lOiKtkAYC0aTEyNxZSDTnw4WVqi2
uQ4MGLrnWP6mifUjje4H6vmkmRoG+ZZ7rOB+7EVU/y17LKF2hAFRXZOHWJ0jBeBGXwAA/Dsr6ptV
ijmGh3GN0q0vQ4XLWdYMAVnXMdg8n7N8zIpd57TEjY1wLUwFOuG3hRbBnKrTLNRKUv4EIvR+U1Xw
SyPnkWrwYE1kMLOS8OBwKYGCs4Sl95H8nJPFvuVTV/U0v2hcBElQPW8WjX16gxDU5SPV5ZnX1fRC
346KFr9L1kG2XnzAijm3/SJ9QMNXjIblJGIuZ5Q23DDb5NPVaPJkRinXbpPDWOXWCQ8CXIxhZavb
h/k5ayQQi83PX3epSBvp3T93LHZ6tDPpQ1ivYHcFwGaXu33MVCGhHqkvkdHGAVZtMcKBS/fNfhwa
SdcXaL2rNLylkFplnqrK9S7+hlY+2mQc3ElmCGgUp7qZSFdSsjEHGmZ1tujmkTn0Y9bphk86XsWo
fotgom7Y4DxacrTzN5CG3YFNSwPyVZ+AnmQaCnuwKWlyxC0DR15K3XwoHDxzr1tZml+XNTEw84MJ
3/9il5NIxTapSXiUj15ybwxUE/qL3NNeT3XZ57ondmVh6ulACqys9Xu8mlYonznpH+hGenKqPuxh
eBrvczNtOVuPJ6pQxGpYYUJjBs/+czYKe+UPSaayHKZmiLaaFR8K9fblNjcI0s+I7qhu5f8Ru31L
joKScW0grWkRhabdv20aeFHwMG5g2QVK+c8ZPuVfm+QV/b5o2c+42VIImg8Ai2+I7W4dHWxnhhsR
x+zfjKyhZwptJ2DpJduFKeioV1Er6potzv66XDTG01LnHJbRdWCSN4FFJwCXeYA+DMb9TO1MeGSc
hYWQOwaKOg/6O3i1Ge/kybDu2MVdBbj2pXqppVt1eRSyP4tu+tlq1stXEWLRI17RdA41rFvgC0p5
l8N5swxBp+BawrLHxCPrtEWA59s9tKED12QezKuLsSrB9wFNcBfZFPHvZHUmvCxrxDB3rvatZcd6
kAsCApj2n6cLOGcyuC146S2IOvGpC4YvrvWQOGVMnCjApwdWmU0Ncx3ZscV4C7GJDk6DBK5Kj5lB
Rn/EnmwsyxJaoZJa1WaN26a2jyjCYF9HuoeBxrF/TVadX33z8VDEXjlzb909Dj/mm9y0HROP8/4n
366/fE9zLXlNw0CfOgSDaWi56jOZwl/pDOj/85N7y3HqyCpfmFAwibg0skOudpA6lVrQo5s8wpGe
ewQKslORMCqs7dZUW+lQz0dcORE/0ezYX3a6i62c7s9O3Vgb5k5QWe0Kduf6EjkyAi3fdAxWnzhn
66p3ljvisyjL8nBoynCyalYavZOIfjZXfR7Jiuk4XPKWu4rZTbHmD0Hxt7iKFXFlHelH9zpGnbE3
GXlFF2e2k2hjO8JSw//vy8db1O8Q5BjHqO3UXlaNoSKWSdsVHIkTx8oE0ukcsm0bP8h1dpio1YqC
QQD0TGCaVJulhW37/pqyChu07EJQmxd5B0v+q/TD7mRmtQmSNFVFtHAsagi+CsQiOi4EPrpMERY1
VSbWtUs6K8ylkViWZwar+tk2bTL/eK+bUNjcug6KodRbZd4xyelsai4+Z8sPXRBLP+Uz8eV7VM1v
/bgiQH2/O9J1Dd4v/AHcsbQOpVJ49e+my3XKF7VNvfKQCyClfQ0Jw03Ew9GeAZnqDfCnS99Bkonm
PL20k9tSQK991JYUZBXSlzC7gxl4/X7zwIXiDWKUow/hhx2YX88TvJpBVwWId8h5uCx0VIx+bdV6
JI0q64rHRJSazaP5prgVGI7s4uwhtoZqPEQyylq2hQwa/pmytIML/0ssN+9vVhTfnc059DYsFMVH
84g2buECcE64G7CX2kKFLnw16cGxF9Bnbh1KTVqlP73AQBzN/x1QrlaP+rZBd1CZ+9dtLAmi7oU1
hMUfBMUqJ7t2jo2ca6Lrl/Y/E5Mi2nJhMklINTyRdiwndoGKg2b3KqRGBIUSMvEeMh/5YSNTLIEO
Y2xmeILeCcpGu2fXSGDtkaxMjdKD+/gacl7OgTRDIzPAcQ3CtouVDhrSCWLbKPbPjxpiriARUfA2
cpyFZ1YTwMDMVO4q55JK87Pvbw2maVhQXONv8rNj0QAQc9SLZ8ubgawsPcdXrEvHRaV1DPE7ZX+c
GE2pAsSg7dhQRb8ONix7NYsOEeHQrBSbwZaFKSsSysF5zsYU2hvgJw6TkJeJRVQJZNT25oR2klZC
J05+kp0fpoai819e+Q1e9+anwj6/RbDobOMUxbz1z74V4wZ3Pi6U4CbjqvZ3o7+n433Din4SWFDo
MvIoMVDTWSLFSSSm3Lv6GmQUjI0uXK6ctk2vcKElyRsh1kygldZ/8N0cb4Du4atIEzS88DwzBgbS
KIt0tziCMepkmkNKLZGqzI9rP9lfgNrpF6P9sIbla9rVPGw1kS6rIFMqtbelv9MT5y0oB/mm3a3c
EprpLjZyKBWgLHajuGS2vToX5bCikZocvDRkw0zFFXEYu+HgVNA0IGp9ibV8aCPj+G44j060Dlkc
A8JuvYZ/huyB6+jNs6q+pJ9kQuA16HnZl4bnha7Syrn4VlqbaVgItV9bEYyGhCmrDye9DvJcMUEo
tVJMp1thiHmr5dPvA6KD+yYqfJOtjV104CxOzjx5bGqT39DqCmne0swJDCyJFpEiFSdbf2uqeL45
yH9iBiUMwHBl8/3GGUn7YK5ObsVr/X5461W09zgMD5r01IktULHR2iO9WlQxXYILJ2a3COpqJVcw
rZFRIgYKKV3hqvk+5pVsfZPfhs/rmiPgX+HpC6t3WfjV2D6YIuhWKiVyB3fkTp6CopmcSAezzeJ+
kXhbWYUy3uP9PqMhbfGAPKIWUf9DpjSHL8AFr1AQN8VgCHTlNCTKmDWbWEM3rGCu/s6t10ptZiCq
nOhaJey52EdQiFDQKaeGvau9bi1G928TuoxlZsPvIPw1CdjqPFAl0Ra24KFx4ajnoLEY3lG8fuqa
Dr85fOQ1R1CaKbNx4RwWn1ItTOLCMm8pjHSQR4VWcfE55OKXJphI85/lr1UXy+WngsA+hcr9CpqX
LradveKC4uzkXmOHcYDxJCbPH098f6FKxEBo+L6bGNREemfpzvWsTsSJq8fHD4yQ8DBpAc5Ez5c+
lq40S0dcZYAUc2tK3qx7u9fVEOAd0G51g1DSHwPCI/Ah+hXEyP24kaIb3pyKlee38WzIxUln5pCv
B6Pu6du5MKfRK8IMRq43NLVVh+MmNFkcBrJCp/jQfD+139u+5jrUhz0sujWN3fXdLyjxodMoggPZ
6kuxYdQgrmrNcry2oLwsmKl1OwpquhQzSdVJ4EiLvccTKDV02BNS9wk6YVwFbsGgFsnRFIfSnr+J
b1FoyVSYItS0ixfDTwBCkt0eYKvdBdTe7M+rR2ADqK8m6H/MogZLk4L6Miy+jr1Qo723vnTSeQpI
hOuPswSoN6ENwuQVsKYPA2bmJlr/7Hd9M10V5aZU2snEMrGy1UqZg1hBUUN3vpmPFmugnGRcwEb4
kUmtRoUUooH5AGgyzgk3Vnyfg48qI4To7/oeAA8qfonrNE4c492ByLmQdsOsL8n7ySO0pNjRTTgp
fjuvfTmwcc2NPDz1O+DoqGGWQJ/Mccdkv2OQV3xwR7or4KplKHlwZ0GoLQ7vrfr2eigLgezdbQGB
IcyZcN5A2ido7fZQmbCM8M7iuECdXpfxQrm9JiHKyiY7mJ150S+dXpl6EdG/vxa2O4qwpx4RUUdP
VHx2MgCHkmGQv4B0DEnn+LKgJKS8TpGM+bDjBjQ5Y/Jfl1Oru/kPOeJgyFQxlAnvuRyrOje7mh2l
d8XyP8/ORKZD3uLGwK/JLhRGjr/WVKPMvbZGirlhbyTFobslBL09DK8r/TDwn46OrcsVe63ytwSG
mMonzhiOMfZr5sI/nVSx9gHVIrfySel8r07Kt5ntUGv5okuhKu1cKKeeey1B8Z55ZcebIWLjQ6NO
f8RAHmlZX8yO16AMz1R6DAKwYXsI4ElNV7Rg9IksGWOtYHDKzV+llhd5llGfzquKtggvVLVObpOw
AVHVgG1C0xDLmqbzJOq+wg5GCqYVTBlxdZOU6mBk3HKchnJJjG0Txb53Ce/deQEtEGajo93umAYP
9oauXpQPs2m2Pt4cqn+w7lQ6XcUqx0VLQgaXC8NcCTxbt1XndyvaRi8i1hqf0oqFoLRhQQY4cAF4
FhMnOr/airlKtgJ/Ly/GPQwFG+de9O/hz9xEQA/EzJUb5VOAbLFDML32s/N9RhjLE7CCkNR+iifp
cpRz9zWpVlkFYEmtExL4+/KCor22qHBne/d5TgwMIAqMZztbtxGy3vLrLSOycz0IdrIL1U70R/NO
nDZ/DseT9PG1AwvVzX3tV1YEdEl6oIDP/N0SbIUNtFEavMuqq68+GU3M7O5PZvV/tosK+yGW1qTc
yq7mVt7VdhExawOdm+advvwFukU/fK9yz7XGAMedR3eTGDYR/F8lmG9UGEA7+TGbx0qP2X9DnzQU
wG6EOdFTPqnhi+3lyNja4kiUhZ/5NCWLg3e7IlqCbht2vbnLyvsFib7FK2qXOZ3/DOB+LKKpKO7j
zyV2wsNDr8/EVA34rFHmUnNupxacM/YMBovZMxP3j+d5wd0FXPcQ1CDtCCDtqFLjhUQIeVv7363x
b9Ny3HJ+0iexQawS/s2S8+YFDvCstXaJ1gKpues7nQRHTzjVopW1RDmEtFAjt6HouxdzzUkSm7pL
Z5iTAadVZXivtiJYeOnVnWGLbIhQkfq/oAipABSe+fL4Ht7smwUXyC/gacYoIN0Kwud/EseuJT2f
x6nzMw4VDOyih4XuQhfxRHVfrieFqMobbZ7HYWiSosDwtjdLoGpBdiaA2faWZrFezjZ0+z9ySdxB
hYWrhWvgVi+otq+j+STx7dHkk0ehz1nohAvZAG2Ta+dYuZjIeqjiXAiMSLXaR6rQUcCOYHvJnplu
ST6RZJ58LxU7B1jokpDQ3dM9rnAUu8W0ucf3PAcS2uIOt0M3JE4ZSxtHbRTe7j8GkZv7ldlmSBqC
SdEZwWAXDvcbQGrbfIBzNGTCdqKGULG/kpTIhkLFshWZBj0JAtry0YBib/3ONuZXcOL2OANyaGYA
S2oOwq53UCOOfZs9EWAFQyO1nxyfQd8k/LeO3NuyJlcSzMl/eS4JVQq+i0CjVaP5THf+++NN4WLK
zR4vN1rB4FynIlLjOS12GmgWIsgP09vxs+IZIcK/aMPnBebOl78+ExNGsr9paKYdAH/TVXXlaQyu
Gkhbs90j6sCdFqYa3hVIHmhgxTidRr38JM+yLFJvaCupY+S74zGWlQuQI9EAbDTGFfxXMZeq1Z6k
aPHPjjxSTtPzE2sdot0ymCHCN8OTASzS8RS2VzhLVKmTg+u1DAsPNGztlTT64gFc8FdRbOCBDcMp
g+znuFSS9+CcOT0i6FvrNuJ6v0Ag2/lIHGL6gyp48/Q1saRSQi1X88ky97c0f+KQCGog2fa3LTXf
V1HkBNY2ikFbIeaQ0/dwLc2s0oeAQIjFuQlevqtB7c9nGJQDJl3y9jkVK/9u+CtO2wr+0j3tOrmd
Um9jSOrfoCw8nsFi5lOn/nhsUOXTPi2coxUxkt5xNGg3wKYuPOtoyYesSc3q1W/ETD8w5HDHGOoq
BEaF+NqQV0IX182oU+Q2Z6skd48O0irjm7evmhLVTOZwAXtci4kalw3cZ/MoCZrvkMJNdqAJbdfI
8oKTV7722RyFqyWu6TN47kEAZJAdFjyZ2IYCQnUuyOlL/Mh+0A0stOqVomWl8LWiFMdEaWf7gyCI
8pN0OnCpP6AGcsXqOuYH43e/+/L+rkyuD+fCVcbLqqAlnRP2KwWECPPSIPbdeZ1aCTA5KfKWGa5Y
03I0QMazrdV0h+b1tsC9ZwL2eKrQcugFQM92Z7rSofEVFLBaSM/bSHhRWk+U2hRdlK2bUdiQOP2C
quyRv8h4yhNKCyaPxGPlvgJysMIYJJyJRiy3Rz41l5+A3q4HQMjL3vLjwARnMdMjyuijKHlkWKZU
1WQANvzri8pvsyzempZrx6Nu1kcRxUw2QV3rBnOnhH4+gbGrrAB7IjaudqG9rAhX6uz4UctIsCx0
e9kuAB0VX1DNQf/kG82hYwwbKbFcGRL5MGeJmc49oSkkPM1OLa46dni1ZqAdNLpe8X6KxE1P59l4
lvLEnCOThhb3gU90NGONlWewYZzV40P9+Qg9ZPL6EOgquJHi2lDBaw8R/de0vi5RNJtB1bzURTm4
BnjcupwwKkmw6TBz4mWN9vC+2tg5xexh9vbd5twBelcYQ3xHxPi05RRZMgzteX5U3KQvKXyoHrvQ
WkDlPSv2u4ZSJgPtil93kAQZF+6K2IvHzBJED6kJJ0YC+X+xN7csxjxHe+Y3qc7o5V/UsmV4zfWJ
plg4cX3awwuvpDGVWUIkM+wVd6qnNNCLL1BLCFlTUD13DwQ+EVTL66zN6yTV3OLj0Jv1aojbeyVK
T1ga/zkWiwBxF98JUgQuNN1s17mFflsPiMUegXAeSz0G/vy2iSMIXH9gXTDwkwltc053GaA9jw8X
Npvt/cV+TYpJs3cDPrYg50QQDneQw9A7613Bk1E8TV8mXzashzyJbAiBHzHGN2Noc0Ulu3VPET9y
HzEt5upWYRQw8je2QJ3vh3fXFpNecfYuxuUmRAnp1TZEC/6k8maERbFBaRldGF+TnG/yqRiPczJG
tSnnnpFFUQ5VeeFYpKhX1eyTcDgg6HJdwnNQ3LGi1ffK4t1rWb8hWV9xno1aAfh8s8Oj7FHdQ0xE
dh3FvFo4eS2iwueeMsVz7DZxlEMFoel8xN1RlIqKZYwYGFXZtDoNNoJQiMsf3kuQAKsZqsUuCVHy
pbHqgXilSJo9iTG5haKOUJU1yGsAls5fNYjkWEygBV/hkWDJCV1UDpvIT+yAgX8cV3CWdXonWqbo
X3TUvyOGSnCrTIHMCPNXNBlkBPU1zCyzahv0/2PZbq0+zqQyuTcl788suUnpqlvqulRXOLuoC7Ac
lmRtm9G/CjsQB+WyqX/2GeBYTW2bYWaHrkrOhArlXUIlXVswuXD4i7tI0XhxTdent/o08gPWQRZK
6pSOfF1K//bFLvGL6J3pFRDXL4cfj+zQXsD467R3Bx5JUDsBL3DQV45lqxOLFHh/5rpncwnPKnPZ
trhP0nAszrS0DX2/hmRZyU/0jX0XftzqnN561Nolpz5jMFyNiJjANfOr98yUb3x9xNviR76rerVo
hO8vPfkyTVHCrnUFhBBvLTN96qdqQN+9EZfL4HzAEgavYn7poxs5l3RDo0HBhwhDffxBwQBouRuK
7L6bkCzgVhnxXZV6HNelJQCh66S/L7ILRda9ZFxsZqOTa4aJSgmaGyiSjSjIh4o1rVo+yrZxBCXK
ZkGdZw3dTaKJQefngMK7eyEgfqSrESizRPxfaoyyBRUwZJRlGHyE7oBEpIC4IGmQyUwgRqun53EM
vPJqIXs2VNuTLYhI6ot4HicbUJHkFiASrVGefPeG5jpv9t/ZJavt/wdORwlNcMmlMrSvitvwvk55
Np+f8MRw0Esiy6HmJc5j9jNbr2RPEzpXLa4gwl3UAncDKvfySZUm2GNCv7rpDR2lYtjwE67OKZsg
/5UJvxzRwOTmk31vCKnELGEOKLdQ5DeWjAgzxAa/cnrQu4K1kZvxtGbXa5PMBf9Eih8pz4WyqoSn
WMjL9t766HIlcBtLdYY56xgrGJHsjigiMTbEp54tdNjtW3gUi+G3tKLqLco619tsw24klXM+n9kr
yzze6TkRIgKEnKjGRu2hn/PzhLAchSQ27/tyhK1+RfBf+bftuCsWyEYhrxnei6KVRItIqQfrICgK
4qTgWwUF8DbyHr/zBdJhy5Mk/bYIctSJLUunR/H3oXoSqBF2cBsSgnKoiCPC8IMSjao/Spq/M7qx
Xi+8SeJ1RFNDxbXqYiHHwpeVi3Dwel4lf8QeCHftL1XrtqEWJtKcRev9mfLM4aDpfpArpfjGyKC9
M+wUaaK7nEgk0E2KbVaH0xyPHG6NruQa3UAedVIyFlZghjyx/HlmYIzn28rGo/i1uu5DWiKWOpsk
+Uy7K28TrWSG+OQH3RuCQN1glOdGFwvsvRc6vCBmfcSJqeCL0Nl9wCj7UrByoSSk7q4k9z+PvODb
D/8TPDVUGTdDN4D49Zb1aDhxm7vwCUSpWvnjq8WLSptw+QEaoCb2oEzqjLoGkozT47v8ARwKhwgS
O5ioUBGCsDlMfbu8si8DwxqugzBZstDWcyjyDYAh8EbiaEQc8iuLIzbudnQVdi1i4PWHOeUmLNHF
pdCHM2OhYDnwCaCOURNHa2ZbBHw8SuP0YJbnVe2uwScNMPJ4K46VS1TAlaqzYvV2u3OZwszHcR2C
xRj+Ipat+ukVNvek+JB+esccNalCvDlnk/WPKHJbfnI29dxU+Hy1xUna84GK+bBj3/ygaC1LKFYR
74ODXo+ixhUcrFlit9ADEir5PVb7dvnojRV1LovIAjmflfex+fnp7Z0nnN7ttO/eriL6wEVLMiFX
LIbImlgLrA6tWE2kT8xgBGyhkhIltxwxjUpRcN1oOAOR5N9o5MaBlOiRZOedceC1dNXE/j9Ju5H9
cpJrTDj2BDSp+JM6OynmCTsE2dzBJw3e50hpTnaWyvtFYCwLrfeR0DqLK4jnagXPh/yD1CxkjV2V
KiEkpH+ekAnVakxuTV0EhbBkyOgAphAeTfNfjDG6Ee5Ns4N+xMcnwltdoAmU0XKeWRFPgfElcXFr
UL6htLz34YVa9xDbyUM0tr5Dt5ANKkbfP9UDU8XQOgEsRoue3sBvZjjId0GsjoZBsOzjT6O0EXvG
WNvi8vpRg4YCpKwHjkZJjbLgHclXvVgSBI47OFSzhDpSeKrlmsPyvmQ1pchrtYYH5myAzivNWoLw
NwStX6Zxc/VZ9bIUSAXJifXSty8m8Q1fVwMCIzcEiM03wLuL5FY6tBGhGcbQPBqfjr5ug4rgYZQO
cr+QGF1UIOIUWKRxlCzjltkiwZYqGRxQPlf9KwuPg804z2xB37SAiLJeaDfMG2TCbd6fmkbh5Ubb
rwmYb1H1nHkWKT96CM6TlY3USYI92FBEQxjLSMY6HguyHIrfqB7Z4tMSlgbYISTANr2tlnAQfJGO
hw+DxaMiYPiwWBfkmm4AKC8EIFHaxRu9YxFklYBvUR3m4Oa7TN+uQQNONR+tjtywDpAqI43LgPxz
0x76aUXJ6XB030cAJbSWS80eUT+PsEYHwpTJniskB0bGoEdFn01k4TicFnJtd54qVYdD1viXuU2M
203BwVsC47FcfnrmYLJIzL2xHPTCUPuXK6qMzEFNwZRt3XwYsYo/8Bj7ANHmIASvUaml+ZuGwbBt
Aum2nvQPm88eXdt7Yt4TKlErrtgW2g4Y1QuFOr/FsuAOaOaEqypmoSdVUAdpEi7KU0a/kalz7Jxv
JauucVFjZRFs+lpeVr9lupaGbS2Cac8ouVS/4tq635bdNAF2Mpzl8k4cM+WapwHQCFZzvDOu3Z1q
pAQXFIhQdyRALGN8QJw5fLaiYDtBzaITKKCSNvGjS8EhuyDYzAHvpHKSzxePL4KBnRksSViRxiWq
gQQZFeYfNDsRwZXyIvNJMW5q272+6nGnQz5rDkZDhyG+CzpNQ8Asox2YaUJAyyaa5pX9k2HZXnD2
1hl5fDiUSaZw+hIYMaXhopCcfqxRJttt8206j2eskcaClzwaYrkbaclv1VE5Ke4EZlhUcT3DQpwg
RG/SaaxqTIaisST6kbDd8goMI0TOaJq6qx1IEDfu52IsURF4Fi3C9BOZXVyGs77HfErrrv/FVPTX
NF80YGnLYcFTEpM4n4SCRg6yvT4q54dAK7TVJnRJloOCjAx+R9Je8SqPi+NUajufSLIID1/wpi2U
e3nm73uPXjyhxtiilFgCFzSACrxxWmNUMo+8tiyP7SIpp7ibwKlNX7f6rP109MfexjxxJHS8D+H2
rRawffr1CsRkZA19lH3SJnPKTVmHVmf1niSqtW9M+VX+bzEFyX5yKJEirBwergFdFQ/L4qDiFjkG
UbHeY0TNbvkwQU/AAAzKy1HCcqrYAED86qBBJ1AM2wftxqQi15TzhU8i6uv3XpN91ytraZaCpu+h
Fhh+kcIBDwUeO+g4I+qdaZdojTPLD8/dExE7rTgsE1sIL+xSuK10ee61twyQUzwr+O18aZp48fBH
t0ib1vCZ13GiuQQ4891fe7z8uMAPXja1oiMr5Pz9ypjLlbt23duDvhD2xL8xRcQi3RfRYMlQbhiu
X5wuCzczsLHioTto0C6QiyhCXBI5Wjft6isqNia1uOEAIhc1+WqJSb1fhqaInO+PAU+v494zE0aZ
MwDARUQ1QB4Mxuh+HEpfRT2D/fXOO8PJ8Q6Z8HEw0udHatOY6hIVw+I2p80Sk6nWqhXrl6uBpdj7
CnGuDrTKe4mCkGHXhhLtFu2hXWf229ZO65BSmknyhnc7a6lMM6qmQ0IDixGJwdK9nm+YChyeZ9Tm
ugkUiLnUX5UldswulbGTNcpOE/RXAeiqHEMLwRNxD6yGN/kP1JunfGBUpPUoQjmq6jEf2ZYfG18e
6CAb3eBpmdpMI7h16UK++w+ub3lCxAItj61Du+YZuP+hGFAMQYo+LBGFb2odEpR2oKFWOmz5gp+V
Ipp9OKjQvIcfQANE1Yfas7cz51w8QD31zrWsHs9CjDC3KTdNfBhuI29teMpSC1XdACFjSVJK7vY/
hMwKmJ2nft269DVl4Cs0kSjdbwsAjLWFCO0ObwF5XX0Rfe8kwLd8N7k9jYFh81uqE61l/Y0B/7CK
taEw9PHxSmlr+OkQW4UDynuEroulCkinDa4jpaOZpR1CFjYKmBNAgP2YGXXmcHIwtRul1lQwvmXi
41Y0X61ZbjwufY7SrTeXcHViJvIQqnF0ERggbK5HQQo42IAkm/5wRprQ53+Oj+fCDv/GujkyXbJB
r5iFjwqHPxP8KFz4JjUDJlUAz1P/eu0NXzwXG7ZJtRM7aqDhmRXU0/A6XCKRBqB76Xnp6NwlzyJU
bMTdhOBmT0U/flALOrYyPIrWCkmZayR2zepxtATjjq9x8Vgp3pqyJ5/TH5UXp0FyqhgXLVJNbH8L
PosOUzxsJwWOFZCTGLKuEXnBnMDkKojGivT6c7JJ9b5+2j21e9/ZwryFxim6yU6mVDf4BTMrZerz
O0wpv6yuPqqAi9Prpuyh8lOAe8ORlyZTzaEYSz3XXlx6zWOjAG5knoF3RYBQxDUk4laFH1t1IEp/
4SCQ9DhfZr1SZw5xUPn/4E+VpEMFEl28InVWb9JMDfq054ULyPtZ6CXLhR9ECvVRld3MS8TSDdDF
x9M3uz4SKRmwT1BRVlULjYC22ezRbPgjrF9vx6t1DteBIIlmPipalPkxk8+ccMnU78QNsDf002oV
MYylOaxk7fq/5NKpG7jWG7Xykw/5toWvVL/PDr0Agmxjwy8N5Rr6YLWwB+hjpan7MoOMSa41o/AL
BiVz4HT++mI/AdLeusRY4VsnsQF6FeHaEqEmjA8zK/iIT8ZUE09lAlyze78MzCxzRYay2N0tPdj1
wk88E8dP8McT+oegXjszz77wGMU/q7O5t3iyCym3t5zmQCEnnlXRxVaPWdXDHHS+Uzn3ATVLx0TJ
QCkV16nAFuOky/FzvtOUGRdUwxlrV1OJZrX+cTROoxNxQu+FO83aS7iWuG2oIcfM04CHzas8GixU
BAI8q6g2j+7jE/Xt5KMmR7OMaWRLhJfU34hxc+mJssV2/PqXaCB2lXpkeywQsLD1+yENj5LKwW9u
tV6WwWx4jdeOmstViAvwKa5ZlBL0pDitWol2xqtnziL09L7dLLNUWNyxMQA/2WlPuJ/cFeariIGO
iZu6nzyxs+smUPs/HLhRXmQJvUJxSHi+s7GYa6O/CQeHsck3LKxgVDZE3yt/1PbubaQJgDPyWGtz
M7Z/Jsv7qwilLIPBprj1UdczDn6c44OS15t/BkutiaHYC2VnvRpz1/tC3wYu1tbjhGaN7cYeg9Te
WOAl5pH+vauSpwHN//TU0x2AT8vK/VthJsRD7533tzXgzrEOcUwGDSnaOfSRyZGYw2JQSnmU8eqj
fRCbNyh8I7z6ftXJaUo1iI8xgVRSQ5VpeLtwDZ98djzozepVzkknyND3Vfo4jXt9M+cCb8j4c19I
/hkqM8ZnpW4x0qF2jaJ72WhHbbo6GH77r3Jgaxch+b9PIE3Vf/m7CUMXShs7Kowpphjv8UTIKJYt
pDylohuWeG80dwrtR4K9gQKQBJtF+/8bFiw9/MRBN179LaCoovhwjcrwm3Yw+jsnKllSbWfayoIT
6254fVv1pkGU5oClkSfDfI+jx269NbqYfdCECdPK1gILcOPhtK3WyOPu6dl+n5+x46sb41RTdYPg
bNPJ5waRslPL2PElUByRYXS4J8oaEI0rXuwt3YEFPRtbOf6e10xNJPRjUmqJISmYWRnsXm6mFi6B
BNPLZcRwdwW63j1ZtQuJ9a7le2aFBlnnLf8CdVg7fIznrfSypgtRpSEUa4GnEC+eY4eqOU6dNCz7
Q5WKUv4NEMNvAvkBY32RuPHAw/F9T8gih3Xc5neuWVf1T+iChIDFP731h7m5FYaLmc+Vuc8XWpt+
qhWHje64EsBZzd7Sa20qZpChDI0W09ecJUywLJ5/KJuMC80XHT7s3S0IobAe26l3Jj9QJNE1RbS5
CRFkP/p6EJL1Gufk2dHO2Uvg9YMo3IDK0y1c9Hz8AnTZ1y+7PELqbIz0sVONMSXPHgoUqwpsfGLz
Um3H//TChZUXZl158lNFeZ1DfltSPl3+upQE3YeWVQFziJcxQSG57xjT+xQXS6tLINFFJ9Y0FWbB
Wj1vFR41Dl4H/pmB63lbbwOBlUBTzeFUNa1c/yECHfW0zzrgPF2Q49hng/Qve44wcprYmGWMlMAx
Ekr173XvedIkBB/4TWEsk2kH8MrZXKf0kI+zsoEvYp2odgMWVceTEzqOhLesqWozAbOf0FuuSVzY
0om3dHrYtqFVYf91zUXLnQ4jpEb/SbGBbdzQ1qtpSDD487DJtsP7bIn6DCrXAGX89+jIITt/BlmG
ANdSaM3KvnVgWxMqi05J+9Q1zxzzbOGcbrvIx7D0SYlCjKtgjEj4NUo7wR0Jnv8/OtDxwCwxdbwh
YjUl74LBX2/IBaOwZepu4EudKRHPYQwm/u8eFJ8kWjo9emeBHDx4t1jdB+HXMEhaPNsUfihdghP+
eGwStKRmtouvFTdBbttoWV5HarVLZCD7/Xg0KhHD3zt7MBh3sM/0C2dBE00ftMSBmzYgZppo/tS5
CIxt0PapRF983+HY47BoGdhw17Q1HoT4kedyrOCyvBSisrAoojMPDLqQNdl/2LnHzSfbcnbwPHqt
ZXSGzM8bQh/T+y/mdPzGMEpvfdzWbbqh1OlzssqnbE56c2qUZcH8AaIrwky/7Of4wKgMkIADd4jU
fCIleIm69ymx7fWkGSk68/XCSjNBCF0iX47ne77l5rwE4R5JXB/imLDfKMeccIljuiQKK6q9jnCp
S6ar3FuGekoS194/K7a3UjdttQ7EHvdS8wkz00AGCtF7gBEi3fxzN1WwTNPnkdTideSri0gQD7DV
cqIBxy5abjyWw3H8kPq0wTm7O1GQAc8ZciPcNuXBJERpv1ou1Pwdiplc6zFg1EG2GoqpeOcaXuxu
fhSqJda6qWNn++w1qHTH+9f32FcBnJNETP+gTLCW+tB7hpTd0CtTRLOu++qPo3aYQxEIUWuIclCD
furFeiEyYMeHUcoHMEfeOVQcQfrXvToxxOn3mDYVMQuSiugg57T+vjebOwXVJDcwoXNY8lcJpyEN
/mQWpDZsL/J/PyYG7EeiShKiuTLIaQ4KCiMLtLUnjAa4SxWvQSpxwqvooo3k4Qguvi2b5eD791dg
QwNYWaBMt7BpH228fKWt0fPdjIKiHTwP0EFBMurApJvLXcO4Y2syjG1xWTlti2kCQsBhe0NxQHc8
3Y3Ln+7gSgknbXIuzv2+t8aB4S6AbblC/vONiPfW/wVXXqNdaEwwnhPoZq0F9degbLe4uLCUnumx
gh+G7x3m0mHfmuZA1gCo7rSsQ4un0eSz+YoAWmFSkMxGcpTOreofVUv9KQ9u9YE3Q2c/Ygqf8bEy
PpG9HUrxvs+NG+cwjuo1lOM8K5Qeywo1wQqV0CRmL9lQigcjcbkjl02bFCje3srTdrozJMlCOjH3
nZWIHuBe8DkF3wRII00X8TA6Na/ty9JjN6W1sCvM/E58Sof+M8h10myqMfMRr+VdCmCiCv+Firfx
KhEw1KXJ09Hif9z+cTgaSaIPdAt1rrUFC1UXox4YtifKwBVKzQHOzZCnhMfuAFTlKVrGVz8flp5N
tfKiWGZ7XkeuA8D95lJkCKng98tb3y/ScA3Yt4OYh3/39aI+mpPatyOefDR+/Dg3W6eDIzDHJBjz
JmWsOVdes+t9WBIp42khuNu11iDGCcS6dNXAap2X/EYY8ndtu7QylbeLIQ6VSliVoDh9ojUQxH6k
nELf/ygfDdWpEYL4vcViiCNrDalmbLZ0UrEQ+PdJdAHZhSgQx6vEwH7YDYc4vEy5pizDgAHBti4l
T287NhUK7AV6YtxG91ct4SnTG1B+QutdWcbLvbnf3tRmqM71WsdqNZbrfnm6B2EU0+Y5CstJwvqf
qe++Wj/R9OgiVO951Tz04fGH0x4KzEkY5IJfynSSTyN04I6BWrsiQRE2X3lZnS90Z7BL5/517HMS
texbUoYNbar7KDP9q+35fg2MZ+EOAnGY1QwrnyCxay89ysHVdTnoFdkpTn8TrioiL2BE7igxzIcy
BPbwTZk/CsvPpmI8k1Z6oS2S+5R6eBgGnjUKksFJmWPSYxONO7GNXho5CGLbCH+npaceJnny95ca
Pb5646/tSptEXbdCWLAUaop+klg5kD7v2w++AE6e2jsEtE4dFwtZQ2G0GIRlBysEC6Cvv6XUyxum
LcY+rswg6+zMUJqOTylIjjcDzRtaWjGR19Ji0OZv+vil1n4csw2nam7HQfo3AhcyX+G8XJs2L+qT
yu9eV8TYxg3llM5BLINSKc+deIRYpKesVBKFQhwBy9r2PrLfWogbJIxrPAY/bIpTIB5wgmreKexN
SBQEaTB+z6d5r0bOHyv8KnA8OnuVU3Y9dtruLrNVJnoa5zma8s0Jy+Ee660jIEzY8ibqHx1IEwys
RTxJGtfG90sxZMelZ5NdQrBz4EusDfQqzV3OxtpMOoyQsXEfjJNqx+9PMxxgXG/t4kawV0feCRYe
Wthoq7lxiop4BjV3Xa5ZsO2KrLg8ThTZ99GsEAeISAxCrqdPDrhB6aL9iFyx0Yjpk8rbU/kkWoAC
OUKxUTqWxAgn7ACkPK4sgZerAaBazZEgI3KDVG2HUmlnrouDeJw8se6o1GEPp/2XgOiJ2Z3r49r4
f+boBl4m9DPk5APSOsbwBPe1NmBW9gFx7LIpxIFrIeYn14lH29/3t2kZKI+HhMCgJ2EIjovhXN2i
EZvfjw8QlUi3s2u9oVphDa58bfdmb0JjaulWdWcUWGN2fLZhrSUaK45Ubm3kg7B+rV2hPCo0eO3P
SHbnvXHBIi6xg4zaldYJA88fhiMvvScYXcRtzn7CPdzAQMzZE5azeEDDGED8bKBmPiX6cnlTufsK
2+qurKdMqx1rjZIYksV6kGDEuRIz3quT4YtnWJIt0qUKDJ3op11TL/+mwRk077R9F/9JrGiCXN7I
uQrQj52QdUKhMgjZZvqbAjXbmCgzpLIBYWbo2+PE1G8Vrc5LWLfdPRGBRbxEviYEFgVkL/HSqeTF
GLrYaF7ExlvRVruHFIMsg0dDSgkd4bYrdsGuQTq7KmdbCebJuYf/rc/Xx60vdzudxYxl1+xKfYmK
OotkpawPHg3J4u4VU6WGUThd3kqGKCpW9Uc9N2kw9T0LHgvAXw69eqb6/LsMNztugPtaT8dceR48
ORYxUI4eIP3zxrm+VZoFnxXu4zgJ7CxvXlEugPUoH7k9GRHMW3AQIAIbJI9PlYkznXjXadwsOiFI
WKeUk2iHZrraSrLD3W9JymLHX3bGepjiwGjxMlSs1N7LspjIprmmxIwPl9w4v/AgyT1MPG8blD+B
tvFd29+V4OmbatRSelwmGcPBoEgOV/E9gWfv4+c3F6u3cbCo+QnZUBBw4ifIi3XcR/pk+NTW6U8K
pWqmz18yn/K8ytefA4cfYFnzu/cfGogyRYs9buaYb3ilQOQ6SwCSg5yjm2Yqe4J8Bz15khNt04xJ
mJ7jEDkWt4MHLxvMbP5c5ONUCObUcSIOrali3GETRRVihgeQU8GOW6yc6vhHZ/90F7aZe8P2W1IB
ghRStIJ59O+5U73xpYgJct2kxiL/j3DyOhC2z82eHNHS0Dmp8xU5rWPwgjXjSyqjHhJ7MLFC91I2
4iRHZe/E2rQy941GMXgrNLPY9DXVNAQrZEW9QDlKSnhE3C1tUCSB7nNXULmv2w/MbdcdZgUQXDIY
z/oLPzNdFo3XA7+P3KZmMvINlLkzc79lEGsIOfpkQU3MKFOIV/28pv6caadhNPlZy0spdh01a9ot
8cUMhdACmdggvaWG+UFCueOTo1YxO4wieukNPNiXqZccqYpZ2iNbcNvXruIjUtzw0Et33Ffc3o2/
G0BbH1bkJrodc5PKs8WBS44S7L4gQLRX7rD1lJTpQEH6jurciDhLG/nfZBP1oYF7oHgTUoTSgtrI
194hyMSei+d3Hd2QtrrV10E/paz8s9GWU6o6FTBs1D91M4bjVMi6gU4H0Lt77ZblYWBUTCqUID3/
5KDtCZqzvwBZ7nDzOCtvhYjtoSo8/ZYMq1VoCc3W/9BCJ9ImXNlL1lRaILW8NLr57OVlz4kiuNFT
nqs3iFZT/aXsXpRapcdvVky6AN5YskHKiM8V3DwLkCVRflVndUTxjF7kIr45nNf8eZxdSMzJJ1AW
iqCHkXc/ZcmByHoiC0ArVysEtHHyJJlfT+qClwAWkMCZK+CIoSnPb1NPecSLHnlcd+KfJPO/VPgr
AUeaQ0koC86l2dkdhA7pfp1OGAreg4i5ZOrCm4YjDg3FT6LK7CP2cKS9qWVHBMNiYSxuY8s9MfKi
Y2F+o7rkqw4ahtdII0x+vDTKh3SELGZ8E3EsdOLq4z54OGq/TpPKnIxaz4PyzxO5wY1h3XO4Sl8D
g2+FoJG1raFCK1H/farGsVh4z1jRtlyl132fSIi/5tP58yMVxUkTpmk9714ABFE2MvdEwlL2/rDO
4sUStD522QLvcEsL5GdNZax0wVBJZ7wfTnTgBujHuLLl5Njig3wF9tKbEvgj0MMUaJ+MRrUgRiJ5
7rS6+cLHBtCAOZ6c+Au3nJiEmjLJFVKrmnP6maq7DIAYhQxcPmkh7ShoF4tOyRBIHd2X4damNAr3
91+9hoX2QK2tucDjkBFsjg952b6IdCdPRHoLJyZBQmRRbprkQL5SsZX9DuIvMfS/13DQD+Wavmr9
6VCR5c9wQX+ddpdGuOAMuIkbZnZ2wXx/tZuTL/622ru8ZYN7KrpLulWdHtSoIpdipn2MI5c+t15R
W7DcnvmWziWvW8itmJ3fFBjtgmuqJ/hoMON3EZOHJdYKUxpctYxDjysldJxJztZUcX1e0zGM6EPv
i2CVii0LeW2UEcgzYqnF7x8KmLkb1AJmn1eJDKKFGUkoHSxrjr/dysCXEKnoCG0LhgiV9lDQwHxM
YCNXWPsrkLQMmiNotn1hiOzOzs5dxIusiMAqH24gkIIstBma9K0DTpLOrcK2dI2TeRJAhLevgxWJ
8Zl6TPkCNJc36Rw7ct73y6m5zCnUitwRZ0dTZX8KlJj9sR2JFmuElQTwiJQepEIOP1YlwWFQaOtM
Df2D7EgiwbxCp4ZHHU4QMHGgsJssELOGBcbVHCYJYusgM52a3iJPR8ZWHPSD+caakzfgEw1FAiwK
I1zVU3Kz15hzcD/ftv4Iolcx2ygYwyiUsW+lPuv96EiOSZY7eiUinFUaXSXJWSQbI2O0E4YCAKsE
DVxTP7O7SpnFqYr5w59YD1/5CfGJaWFfQezcrXPGU87LyLnoeLtX2D618ezfEO3xDiw4J30C/K10
Dxc7PWrlbOCkl2tI8VO6fT9As58ZTJbdBVALHboLXtJ6hyRWzv55osLsMpRRRic0vch2ne0X06oy
vT6a7C732bUQi8iptljDMqMvzCcJU73tsQpfoks8wMasmK9CNW4nJxMaBGp36rJbVvzz6WrRdmzt
5WJ+rtIh8kxZFWWhLBEScICE+OveGEVDRpYIlbbZSM768UHQiMqOjs8D4j3j/Cra4IQMUPKLGwjq
XDNlBbEwS5FsgD0YbcJiTFnE0SUqpaIIciHdoKwLeuPP1uOku2S4LuYBj2J33AfeInT11WxUTrhC
P+hLLG25KEcf7FE8oGOkpIFhWT53i945/IjUr8f3T8cL4Nexis9P9DV/sc7Z6husTTlBA598KvcB
grY51w2KBbrS+YvQH67eiZS5LFUAdv9AM3/Mr7CoiX2Pyf0zWTA3lOe0cuFY9Ry9n93Eky0YY5EV
fyu8krQlQroBYT/f3eSqVq+y/ThrvxrkNa3ZRnnmb2m4CQF+QhIXQHIL8pkUUoOOor2yUHd6qTer
riARENtudeE8JPx0ObTEsK7g+ZC1Lfslcuuvo6FAWFSTZS1th32gdQz7hm2gyVTSxPDDVCPWkuSf
XFDRUm/dC/geMTtqsO7r/g6B1psFURZeh00ew4eF1LiT0kpTQsIDUUN8p5Gz+XUAhmXxaxjNBQRH
txLrcYuzpnFE7n2QGUaX+1McQSrfP80tKEWMi9s5kwMpJxrnxF2so3+v/ogLa0lIpCSh5PaPiv3K
SAwlf+lxSoQT8G0PdTkF5a0pDslhygDLnG1Mxlq7b2wVgNCihT69Imtuk/CKbgmXtYop0+ipPZCA
CV38MjTGwS/IxiZvgURDTIMDnjjVzIuSzPNb8DZx+pdbHKwO99igO/gwfNNha6yTBdu99yYcHZJH
vjJWIWA7/pcZWC/b5UzAfGW1yvtZZVwZWH+ph2OxOesS11OJewsTKL+m37zbSM2jmE+VVURW5hcA
DzgW8ANANnjkVhrMXJDRJUz9Eb5mAhMhiQuSynapdxzYnFFFpehxf3KL+P3oDsXCfynbIDLdJoGn
/nXYP5nFTTObHeDgMB7dOnBqT+SE8GF7NwCdpUZZrfL1wg32BX12SKC+LdBYNAHj27t+eqNcRgdD
sl8Lol7xxC8v2PAwpxwpGAelyRrf8DVvGhpQjhIdExpYO/2n2Rq27ceMf9mccZibrkanqJ908npQ
5KnnPii0W6XF8Qan87Z1g1raupx//SSyJgwcNsU6VHtjjyBSoQTIogYa/cCDU5ongpth8lveU7wZ
BIpJdBEUpkQjDOJX2eqLsZ4Z/iVBsywCgpyhPTNSduIQKBpNCiSXjaDW0ANZOFuwEjojBNBTaZjo
0pR5wypWy2AuN2Vr95MFjXwQh6UfHr0ei9CmTMaWF4ByIJyYGwNFGxPh6lMnKxZm4f5IfB4rLlgE
WIzWThjMH1OeGi8qBGuLgSbrx0FeiaYRcxtzK2B/jwMh2aQ+06fvG7NUgCET2hNbpdn6ks5gB0jz
RkQeWBdIsA8UOabL8IQNZCSpDWZvpV0eFp5LTLYhJEj7jFFIAlLhbsrLMWRUiAzw/G8Skgg+yjxE
uKlCXEL2XpDXIG/4zwvSWkGQSGTdF6h+aF2H90NtvHLUu9B+ODjldpBcjOsbFKvI9X13aAv9xSei
3/XZGVHbYgouMo/Hm/3XKCoTdYEoywhqO0jmKoLc+RDFnWZ/ZspXFqkGejoAatAhpx2gpSP6wr+L
g5ff16YXh/vFDcaBh4uXlEdQYxlkbCB9wBZ1jTgo9BAsli6fuY3bSH+itwd5d7jXv+d5zIv0ylYk
yepnO0gSeh91PTrzdiB8oJ5CpEKTzp9oqVKdAlZHtyENQmxhCVvPlBncz85N7UScEZ54VnN0und5
oPepkfO41pn5bQBCxJtugLUZwsBBH0cpPSzybPUPdcowiyZdibZjMQv8d7n5cr48xnlgE+Mywpw8
WeT2foS0R3nCchfD9Y11ZQQntmTV7oSLvMxn86wgi+vc56aN/OnygTwRStp4zEUnMV5QbKhbynHZ
eAdwMbeTswfBJK1iipzTkKdPfvkQ5+5eDqRhaOJK2DfpMoyTTXTjyl/65RIgGP7YBPlslxMp+YSp
njbKuEVOaI/pOfjmUZ56O42DJRtxwuWLuin67N/5M8fkgx8Xxwn9C26h4X22jaqlFJ1MUMhwqPGj
JcLiaqh0RGbnNqvETRgbrs5QC9UJFukgDzwi/YmaJM1NVWjxC1Is9SJk8ikUqeMFbfShZf812E56
5aRxvVIHPFyRfJRkLLlFG+7toPNW/FrQixc72JY64Rl7rhDA/POCpXReVd/SOdQbJ0ApmXtVAnXs
ERz4PsORFTg3Z0DBTPIjJjEtaD+HnMHGZkp8A7YrYr7p6nxd3k+cUi7MlgdERVwX2SkSF67ZYQjq
AQisC7CMalPkNH4y3U+8FobS8COf0G4qKQnI9pi0xlN6TZMh3Cdg8ZBgtC+D7a/hikkngnSYqY/W
ZUdH8m6nNxe2lAkVHYibGgGXAxnuIPX65l4ZZ47GfLVVtCFyaWZm8GNg00b+Gr62EOwTguan3s2P
1f1Z9HbY9W5dLSUAPVmRQ3dMbUMWuzPxVnPxaK4lrUiOtLec9bS4FWM/3hOkSwZSSSgGajPVFykm
Nm+DA14Y7Kt5SHvu4yoQXG3zhlUt5kT5VdKJC9pE2bnmwDFUJDOKYy9pnjJrlhAhSyBByjnGRbx9
RZ4Tk6ukmEFlIcj27O0UT6dXz3osXCSr6i/mD5szXNFJfpLhVKR2F63XtYW3mrTufZXimdi4tdD7
pVrhILVUnMVbQUlAmRqgXBDxG+DFhlPsz0whSNCiWFU63SgAQCsggoXb6UFQblluj2zkhWIB6EPz
CqNU5jF07kEmNA9ctiPTxM1at0af9lNa0y0bsx115YoqBykUqi9laVDO2KLQ49gjcOrf58QGlA2G
SpAGpTiAVnPegmzOFC0yDy2S+f9llYEt6rZrVnnBIo0qLP+TOwtkMXZeiNuT6KWN6tiDXnyvHYlp
hSlHt4aCI8Vhaha7JbYif2A/oU1oy6UXM5AmWit+w+fSd7GUsWOKkxtRJaZK+2n3xbKSkSV3CzoP
ex6uOqKdGQ1WcbxAbQynjJW9nkCFgO/pyFPD6L4eop1kEbZw7CFqzBLFF7qvuKZ3lQnZ4njUWczg
2cPSfTu4haRVV8h76K8VxWjX1m63O0V6ckkKpMvSGn0NLVj57nHBqj9D8gzrMBkW8M28RXEDWOMV
kuWLMaIVqXR1BVpe2qHDlBVmJQty98RxnP4SPMmP8Hgby0SjjyYbt6r6DbFH+77Nexlhc5Vssjci
eVd58bvNg8in9kT4FxaqsL39EPE5+IHrFYVgLYktVW0iE56oGd4/mWkGaPAVDLcz9aSZAUowm/Wk
uzpPN6Dwu1jUMGdQXZj7y9/avp/f4NDkmLYelXPIhlH//jxxFy1U+p/9ZfGtkepFi4SePcLjEDEk
z19HuqniDlKkRiysrmKDoI4FmnkDrS7A1rCaJ7xAXKlS/32ooPLdnkFocVE0BOC+9UqXdLOCW3dk
UN3e1NAxylMqm3wxsBFMv2mJVj8OE/tzzFE9Ko3ZCfI7xa3I9ls0LpXMwgwfPLJKXU9KJjJF99In
SbOkQ842svEx9g6gh4GmTWL+lN+aCRYL6zMdko2AtyWuDZpukM81w0bhMWt9eZxBeyz9p0bc2ojt
j+nK2eQ7u14jhU/8QMZ4KDXXaR3CGWy0xUdIWNYj1kxt+YHSGASucL4dPPlHAgRNINjabFp7jhkP
j7xTHIQOl0ANO+RU7ydqagbhJkLkCr74CikfcOjXXXAbl+uDAYoCllQvw0RqcnZVD/UIi0oHjVG0
Im+XAV3K/QB2/caQ8WQ+LoQcSa5YtV3UuwpebVJ+/rkZL1cNfI7zeU1Cq3D/vjwdu7kXGIxtOYSR
hEjtptYgYVvPiiJ75YVayUOSMLVdQ1kCWRzvSRVkftURah0OdYzlIeZnxkkLYubrV/1I9nvRl+z3
g+4YppPdMsR51R9Scl0WjgPGyFl+y3FGHU3zffHPhMPdTbTi0QYwAd/H2rhMsyYVHAWTQQ4Fx04G
6nJmdaMv6lLlPqg9vzu8wGqBRAv0fWn0fVHhDtpX9eAjLOCaT5lWx7blmYFGhmbnStY6NEHieHav
WEsFUO2TIvgaFXO/2REgOiclEZ7WJekqzq706BKe8jxQGirKfSdu9T2VtZ5qj1BRFun3BVSS3BvB
qAQfceN91WIBaJvsM7AH870o/mj8T++YbiUm7+ZDX+UjiZj9XO9f6ziKJv5OhDmcv/TYy5oaldER
3fxXZrBuiGeL6e3PhmGEOP1g3/KTY1QqIP2ij1+nR4jr/WObwqYnN64LknPNAV/DZgUlJMkYtKiX
q6nBgSkPC3VfmuXENJwbv84o+ZWQb5DNspGxuKc0BxRE74mxHVCC6hyEVh+Q7Xk6T1IlJ6R+IaEv
bTRT0coisZ2jsGkhVn5aGMuE2GnMac9WR/fYw4SGWZk7dwexEnQb/8ZvkV0iqluFw3o0Ltyqc7Mc
Pg6SGSMF3An/aYPdBfTG3+Ww7f80jp+q6+9SMis6PYaWxiUn/Q1RRd8O9TXlfN+KQrBfQUmYBbGc
XO2p38ZhMsI9nARc7u3zNSJLqAEQQ1+Cn39M6aVzYLb28dBtV7QlvUtCaBqaREW3EliB/b77ZFXc
YhP/3Z4tT/0XiLgVkA3FlPaqpzNAqiLUIFfP9jfhilNu3/1IdrMxKqjFe6w7XKajhKBRyYJ0Wodk
qMnfM2ZPczFMv4+wLMmxU++M+vr6gARtJ9rbq7cJFJUxlGYI/ujPzrxbSeBBtr4HTngLY6V6EuyA
xNre4PDWKbFtNAW5pozWlnXw7tqOviiy8yRREuXh88h0EAg1nFPHqT23dfC290X+U4HFr+418vfA
VdIeQ4OorJw6mSE8Slb1us7wmoHB3iuxtm4B2a5Pj8iYBp0F3i6dIMzUhgKoK1BmpfuDmjJnzIAw
nUBV+xL8QabWvw/3sfLThfuK15dB6ON6TzbYjn3Ov7jl8IxuXKPf5VQGbyS5SQAtD0qbCwsvmEr0
DIwjyYnBSDoT89vhoYDVJuVoBxZszXeqHDQTpG/0I/v/N6vWCyRndTTzflr7WptX6bU+G2f7w+wZ
MSmUxopeS9HeFqfXoTOuag7woANbolQutJkW8Gh1yAjzPi9V3XSjgo6Cymotbf9ibyl5+eWV+moo
pS7UuuU5GxJdIzY8+UP4vfgiEPkJObYITgjqEn/uwxin8GuJ0PrXRzpcR6RGtjrEvEerUHPY8Kp4
qkJQO0bEY1V+w+03C/ulJ6c1XS9QU6RV0XGt1m7uv+FZhzQBjVUvEeDk3UOSC1Z0RdYew4BNP96F
TTMWuSipbe2N8z7cmiDbGGgllIqQPyo2gFrC0uavjqvVVbsLwykxxFztf/35y2plRatspfdJ2cio
fZwA236Idhomdy3xEkcj6XR0HHEC4j/6zEc2/sboMKWH7fwR6AHg2w22JoagFXZ920G1wLwCmy03
/0M0uQ2/zXb9odcEJlAtJMsYW4Xap8Ko8KhdT0MI95rfMHeVby0AUpycH3wOFfR6LddCFaUQMuHe
UkhVNDAa6QvSvgPvz4QDcedcBbC+t9p0r9B0e9GZUU1ykr7rvD9NyGUIA4k3Vo//lnBt8bUURXdO
hi4fBebMZiGucB9vUCPIiPop3OAj875w3RCPakLnOjwGEKzcr0guxMPsc6tcbzLr+xMn10teGaGS
hZfo35sVvuXbYljQv9olbbxaXmu0O/Z6Zuv+0ioqkmmKYqLzuOUemxWFAfn3/JbveuP6GyYHtQeF
9d/6UzOTHSijdrpPVdbkCxdTGoL6b1eiCpQ5X9RtGEq2yFeKW6CcXJjPIEH6mqCHGv+Nn9fmz44Z
hJUVxzHG4pxb8uDJbo+I6ivNYpUqhAb5CyyvbwSDKj8BgPZVjMTS5MIZM3jloHze+ZJ3dNXyPUzP
PfoZYAMqxibEr999jM2ZYZ3DStAPi4wIUSx+3oiJeA0FH7v6+dPY1sCRXiq4Yft5tmP3Ea32kHP6
csMsD+tisl/5os6KlmjwzsoZLyppCrD3cNzb0M79J0v92m8iMP5dQ/mbqeGexBn6/1CD7YmiXM1H
qxDDacNKWkZMhVbZ3wiVoWpK/9Jls7nXkG5gVbEhteRMFavZ9hGWbwDdabGXgeyaijeb/hD2EPPM
lTuVJX2RGSnDr4Zsooqe/AyeLAVhDuv1H+UOGpwA1dUYnXHnROg7xyD/4QrH2wS7/0sMbCFFWHCt
2NPKQnPlnInCNfuuXCEZnZaRWearJQ2gTJuUclvzaBvKT1uDoB6E7PoGfz0hi4TOs93UMHIMGj11
4OFd38Tbr5FxRPpt4qKDvHZBor9F1AKn6Z4H52pQEWUtXwoc3LgbUKjinngBnZ7KOwDrt8BUae2H
Gw6CGdrVJRZ/spN9RuVxIlMXzEQwtt/0GX76MIB/vzCW5kujnMFUW3l2ZCwtHaeLwQ7X/HPlUF88
FAsd6qkAiV0Mzud7h/h9NVf1+DUfkm6Ngs+5oOs4JsrgePfhK3GzpRzJHBAknsCJLpymriVwu89f
YMPjccUn1gmD67kO88gdbkUlbf8e8muOvSfdkKmNDnt+svRzPw9h7bhKYrRbTFtvK4aLCt+AzOWN
dT8I/TC12OpBLizW3fIvoXoDJ+eajvb3V51M+EzaxdDA+6AAquAa7t0BksZxs0OGqLerWKKVhZer
SIwkgFrLQ8elgdy9Za8Lmt4XdYsyV7ikmXZVt0mjKwFc/a0jNYKH+CME4Cap342iR9begmWb7B6H
csejGximmPtbK5Gro+ZFDdzZNntYM5RyyJ5+NS+zFrHB/ZVCK5xvu8sn+hWgoW6GCmq+10pDAwo8
MoskqtzYuYbgg4yFo9ud1lZ0zI8EOCfyKcdMd9X0HQDmr/VOFByVpCMvrpDUxe+5GZdgO56TRwRB
9uyvSewEJjybXLugtdX3LDR4MDaYnfUemt3LjekQC/HoXlckAJFqA4XG+dIDPfKo6Lw1IY4mQTbO
fquhUp8Qhzpe0hFION3c1iAUh6KXyytmZQ7jcfhnTVYyzSMsE2qHPFpb4H82GpGhJ9KjRSYwkHst
qEDJZP8c1v4uYKsuPPeYdR8gFu2HXO0oLj71HchMifF0UQd+SlMwNNPEouPzdhzDrB1bP5ZnGUzl
uvUtfbEKzfJBfqLeKVytLAhQUymfS53GOZyW+wHV+p3Xk2Q5Nu5mA20g16WBlmKda4sa+1NoB1aH
Fcuiyb+5JiJ0+xgV34L5G/E/pT5QsQpw+FmUHykhYXz2TmNMeIsaxwYqC1EpkPQxGJnJ/H2JGv4e
ZwLK0KnfCxsX4qTbeIg3ocwY5jK9WVFdiqFMCephrH2TTGBo6Ihug7H9ZWbsfBnQgiOdiIx2j+qN
ymPHFnIx3Vf33gwjUs0txq/wQmMcciyTLqIr9nwTowt+7jxfisXjR7ivXimNIXAhOPAvvPKuUUNJ
S0raGk2DXTuXIxh/QpwQCWvRgnJbzFFlBC82nxNOXn2OHArW9RhLNUlohS8AV6W0+QbHN62t+Fze
/my7mbRMJeyATF/xmBDamurpjWpPJbVe0v/jlzwLgMvdHEIhaBeBTyI4zVdthjFK31QOr9pKc2kb
vIeQM1bjegOCljHFN043T5DIzDZIf1ildIBqZYImJoJwD2nbFbSSUTF/UOgHuM4VK8+rDgcn8CTt
VRsrCHH82lSAVPb0oz9sNcSyj2+55510E3EaXyFYx6Bm1aLM064AD+TNfL0Byq0rniTKwLB7cz+W
JQABw8gb0ygwTvD6Z4WN342mnIDygp+WXr2Qht+PoRT58+Jt7xQKGLq7NyVjzfrHl4BI5M0hCji8
te9mP5G8i2KUl9LqlUns0EfANWHzZ8NFyc0LmjD441z8Cwjy+TrEGZo9UixGQlSpPeYQsdiBEJ2i
IL54S4sPQldU5hdDW+6WnIC27tIL0D8Is7vjTfrJMYY0jzo4YVZ56TNt1dIlVPMuoTnWDwyQE57y
CPWoBlkIq2lSXGSMMnUn73BZMgY0NdQZ+DAkvhy+H8GeAI8kZ2XbZtwL6DBPUXHYoUVABASjLB60
vGFQtvHCUaCYzlz0+NPwV5XYYV53mlzqeFvtircFXpyKQrEJ9/EyLsFIai/sz/TgQj8ixNvDx1Hk
ZU45K0QyKFUVotHEZS62q/8VpVhE+8ktZ4xN70edZzHLxDmyEd0Rc5XPskRnkn7UDnSG4BcoxluO
4FeLFELIz/qgA1MYmyUugIC0TRst6meNY8ND2Ptvj343Qt4PK54CTA4oEE30gwuTJrOIBd34TtU/
tt5CFyo772dvB57fPBekdlAQ9FbWd/OXfzwehtfjnNJ2vpFJXTgoFXvV1FamGYrPIx/BwNXKHgEE
uFkb1JKqtLmSCyEBxNwOVod/19URs34LK9V9OZ4Z/yEpVcLwT/nQ5W4ygg3AibCETDGdgDshJBaE
RUBBRR0bjGenb7OtjbrMSUzLVQevGPGZaqYqBRk+K2bym6YHH5RlE/Swwmn4cAqAJj2FjTYvRBtD
gkUq1EdhP05jQUNn6xs+HNYC+/QCjWK9dhWVY3Fkn8OVhGiL/Nv6w7l0X2Q2hp+aDRECLnxqM0sM
0/2pgVbQ8ln9Yv2G98Ee1w+L9QwupVy2dcpcOgsP4jeBb2qCWRnsZF4W82pDh7q9lCnTNIr9i/np
CcKvnXKcw8w3BQ0KEPIwiFCdGal65QA+eeHPE5MEPgqHI3KLW07T4r288Q50L0UeZG5Gna0JWMN0
JtztS2wnC690czrxO0Y4EX/8rAJpeoFLUi8kiQFxqefjUnI4M34cYVjdycDw7uGrNgCYyZOqpxY3
UntZpnHc4yhx1NaiZ+JD+Djk/9y1rrdcwUJEKPwZHtAgLGakhOlVIRc+V4vDJOiHzqs2DQgfqmQq
vC9CctHyCGcsF8DvHx48ldQWYXbX5AKMEZSf3SgcRSYyM0ROmiVPGbVYvCxk2g5XniDWE3DXAbLv
NEs2OCZLwJw/hhDa8PW4LP+lj8hplBQVq0GT34uO27rPFUKDJO1AXRc/63mr+0mAaag0S15lq1c9
S3UPb5/qHeWUdH4MsT0owxDOlpFeHb3txl0hTV9mxwN5rOtBTMlFvokzVSo5Hyon10ejD8OCdA1f
DDC6prXyT2mN/9AkhGnyNzwz78dfnsjPh9Hhq9tWLM8lQMgYNcb9D8AamalPzVdreIeIxqi9yOpM
r2FIzrg6PPbhps2yYRtT7jxajFEgdhZIwWIA2bEQP4oVGZsy2bQkI8LWYiDdId17rBysYCITQQjj
kZVWASGR+a0dB5ttIH6HwlGi13kDe2Vn/LFrpOJDk4BYEmX1khnCEe4/46A7JDhymXuUUDeCZ0+F
pny2sbW455ip+3gWgZ4tZC0BOsxcKFkJ86dtgf2WV7rFMMD1ePFQqHYJJFe+qwA78qXLe4+PjkAr
C6TL3oH0j5wtVwE8qVSFEwNUzY84GGEC978NsXW/O25+jD3WqFYajjevnvJi+qe5yboX8FOauJzU
qPLKsv/Taq2Wt/dnrFraqc4CQZ9cFirEjef80dhQjBIuNsAPUhFg5a2ZFVL5+QUhnNIFBg2amCfX
szrPNoaMy++R8zOq1E5sCRnZqAnmF0PNGEgA7bce+4zUoa8rYeS7KKRmNFXXsHxqZ60UeZ6PNzwt
IoJ8l2n7kmNQdKpXukSiLSSbl3Aw3PnXd17OUcG2hUJqhjfqV5k3c2So4JRhRJeEOSnrjmeyhZPb
nGzQsHQJ5ts15zdFKRrjsIJXVneO+Ii5iC7v23vvNVm6OlSnnZPQx3b0Sw1DkvepIOwIQFK2Xb32
9lpOoN07QzHfiz8WbrLy+HcPfRqXJ8VGYGEltrXUCuUYNAxmP7jyg0f/Gc/I0AF3eUb5bvWrhwJ9
EwcdQSxKfDFWUcxW9N44o086y0/iTmB1VVl3wM5Tv72+EGl7O8tPhzjr8SYK9L3UZcFbDY0U+xDx
dPryalaNeGtJE0CTypQN1M1BgdPQWpkKGjlNPiCFpvwEimX00j0Z0x/2welBVLiYFm2BKFUBXyhs
xN5Gy0cMyvx+979K+r/hYABX/OChgdfIbvVjnJXx1P9t19USn1HEKNlyjLIsAWrnuuYsyZHhVMvU
wDZWqKHZ3Xne3/BGQtY6sMM6ig0/5YrvmvdnzwVrP+IVIlWr92gP2qej5iNg2XjCEyW3ifApHPS1
wHApimNpJuFGeHOYZB+C1DKGTIKiJWICgxfrOdwNZmrJgH4XNboR1id/aLCW8iINrLGFbU8FhNhk
nPMeLwh7HkE2MfA6MKD1/RAgRwT9GX/NG2cX1/nymErJml4wljdWhm6n3uwKFFuuq0B7j8Mv2TtX
D4uHZKexVzq4wAXvROAAooi47JNvViBMcxr4nOLHl8qiqv4nXpLKz4qsoEsQsc8+g6iIqT1hndN3
QzDK7DygReUlpYpzigWwumhhZEMTd5KuCW6OLkKmhXpgIIM0XYtKZLsdOWliex6O6PB7a+wO6F4z
6QNbDSSpmRw2w+e4C9Y5dNJRbJ/sX3vNGo78jXtPE9cVWYaW1nk3x4t3tfeVM9g/I7k186n07mqf
fW/ctA5S3WlYd3OSFx3avxZ0xzUaahRJY+NDwWULe52/dCbmqThljbfEBDEqf9wv5EHUWNrDipXn
0f8M9vDVYo/tBZsD3Ht4zgf6+FbNXhWYhZZk2739QyrW79iKJTSFp/im7AC5TTpIBWHkix0xxjnU
5rF7kUAUKByAiBl5jSKXtUddZGy7KFbF/Jt03BJ/n6pe285e2+po2ZxD/Nag7cdEBEKw3soMz6m3
9ZD8AevFg3+SDNYpw3vjzf+Bz/DznOTS7svac48BaK03KxI/WYzXaCJYCDN43wsKBBWudfrNJOgo
EE9hsT2fmPMSgxq7z7hxnDkIUzGmTKUA5b3izYNOggRs3BJWfnys69Zmhzpuv224sp/q+NE9EN81
Ln338ut3Kd0/4tmUPEaAZxuBEknP38sYLHLRG8uaNQu5gfVJZ0uVjErBReiTd1CDGsOQUAI+MYRn
vR00xj+hJRNHuKNMkinWLp8bGEvR2NmrGg+Ew7HtTB/Xs7BFWxtVKFW4ICA5SJLc03bbrMFXcmeL
baS5fQrzfo022mCJvyUGydcHDpdxeCDU62Vsp0gJ/GMMgIHLD6hVHGtCnzLrISgImsp6Xz6DT4Sn
KB0EW11EiQWriYshoT9XTl2HU24a5EZhK7aRUDucp9DnJ/Nr7lB9S77T2c255pRNJC20JRGy97gD
Ep7TeKI1GCanq5N+3x97coEMIGglCmlCJRm+yl2Z1rbgEzZUBCugjy7gzj7M3u4IONehqsIl8DDD
Ch5VWyUyWXsn+Eg3mOAqKoF8xqsCxVfBTvNz5QN8OqN8OfMs6A867KTf+Xwt6Z6nfWsBGYwN59xx
RgfrUShRAfcgh7YvVDaL5FqCtcXNEflMWhsWGtTErDS9NYp/oR5fQDAG6kUK9NCOBNMzXTeA+fe/
CSEpnZLjPOI25stO/GewJwT6ExiP/hO87Vzsd2eSl5ZJR6kkZQCZSgPOQmdB9d4diyBeiPQlNP9i
TxCDBU/IDrsREtcmeueW+iorU5TYYhbopwQ9sL0yQjD1e7df7PICpqfp3LEQ+7wgAqw5Oza2p+xK
PCeUv2esqeQoYFFYcHBhXzE6qCbHntyqjcBrDT16IRpzr4G2s3D6NJ2oqNYbDiXcEG2Meyb9fCLi
0IVoxDQUgrOF7HAvV6mSCYcUPP8PmVL4FQT73jhZn7DKuZ38QXKDm6nM62LAukc/Tcl8NEFVPD0Q
w2THtEHL8goXmuIlf9xnuapjozjTq1ABWsw/EQJQdPLMfReZIBu5FhuyiLQWDH7ECNmksm9PZwUN
WeI2RpA9q41YiVrQT1PLJGIWMZJYhvT8/pgwc4J3vDnRllmLg6DTCLDcOZn7nh4NXlVWpwrGke0h
my1PAZxDuIz70K6JaPRfPKq1Qo5W2tyvGN8Z0jNjukuo8NEGTcPiZYvyvbMRJPi3nQqEJCkaxOF4
KfCIegoYoVp7NHgZijcqRQJNWs2+hH+mtlqW6Ho6L4wW+rheojB2d4B28HWD14PZEMHxPa62iSCA
wSfBEjIRNdby5Ni7snoZO2v+NhOfhUe50YYQ9o9uqu4kyVoPPeU7821PgKPBVudGVewdy3j1ORdj
nr48VnBimdwRn4Yti0rtHg8Yrw/ZUtmCLahIe5DmnIpUdPcjU0rsrdYedyzL8GiFSk4YdO9Jlstq
Z0Tc64g885myJdq5WPaYurt8eAMHVPcZ04TglXupZaDtsN81lqR1X03GNIR7AwHvW7i7nlbjQ704
nZyDBy7bMlMYWEUBuJMJ1g8jO9rB1j6EpoCfrOpd+9UX5MtXuuvhko2fDhuI2YsjMu7qB5tmQyr8
EYONY9coXsHxB2ICQaJN+BhybkfOO0bY5v6dvPr3u1+tgM8lsAKdsDhoYctOeFLKYT4siEVzs+X8
sulI8MI1de7Io7/EGuYgrd7t4XdMBf6F/xKMnSWISsdgIcRiPzVieTzF/vpOzrYAyAtW4suVGf8L
5oJU1owv8pERayvD7nuD6hBNVuJnnLj4CcKbmFsLTatx6CjyAo2JsbKEUDuebZLe0yrTywfPJvI7
aEFo8x+P6aobyRRPrws4FS3+WdnTbH3qS0omEi8rAv5Ds1zA7zZ8DLSRVqii69S7hMXM2WquEniO
fE4Loz+pImTdl2kLvS1lcPq1TniVP8rVZxWPumBk+6TJfvzeLUntlwm8CT7WNFHZoU5bF0tm5YPQ
+psBgRI01xrkAwX3IVMiYYEGFh7O5wxql4PnFZi/CTLlnN5lPSN36982R1UHE9HNiuw/2wvYSJG3
3DrHDOR8pDUZo+qtK2gI8VjOVF8PcpdaSMUXQYGP191gRkL9oP2eIeOJcxo48lQ6dTvANcBT0fOC
KgIPOMkVczl8Bn0sY4bhi1buPNjXrbcgQLATKsxlC0zabP52FPys5L97RoRpXAadJD4jhC76iP72
Y/LJ7PvWF0m4ZZc2/OKAQA1S9/QjYW/frOYtPgX5gtO4PHygTiM6HrEotLDyyf80ps8JvGGjQCnO
1n64iqCOQpLo1zxiwevATA7eKeL3sr8vBLtitdz5sslCcnfj9tRBzfIyP0WkBSDrFepW+OHyGMAj
NBmt7f/MT8VVYJE5SQvLHiDMhdFMUdZkbHd9O0+vjMZAHDmrKJUvZejpZu+lQuQQVZQB/ZkR/Ksd
gJDQb0Upc2pibxtg2Q1w/uFI/c8Xxqr6we67aEon4Ec4/QfQBQ/t2KahobiJAvYKwnx45ssdH0yC
e24/62/xzJU+KShGGNkas8uS8W6llPX+OdzlizH8DDt03weyGWPHXXxC457aUg/E49XkCr8n7BDr
AKnKwDWvoEJs+X9MlvZEhAjUxCnQftwZRfWxGSPvpnm4U0D24QMnEPcx1BFr9Y34da2wFLNPSewr
7NM+7J6tH/ZCesiS1JCcXRKX+eoz497aa8a0dLjRi6jbec1GHGUrcnGCPQbE2if8CyQWgen0tgo/
HhEYzjdC5wg0/gWEWfBUG0lNCVOaYOijz+7yKAHrg2WU1oQFXt+Tsn2MDxzsa9Dh8R0yMfWi892M
/AyvKN9aCm52UN50VRyifDJJqF1btF7psddvIypdRi1chfEeB0CXE260ZXo/1JPiuc7BuD1FqBjA
jS0e11aKbSX/bw+J/ob+yzNKQGsg73PHsPNYNtyErSPxGgv2md0nRMdY+zQoKWKZuqcSv2DbDgAj
q5KOmwjeD6YjoI4P6Yo/Z9ZE2PRudKTHuAcFwlOnHlglfc0Eq0lG04tvC7+oa+yq57auFiurdSrT
y/fRDyZEMCRJoD1Jdpk3ugnM9IG5OO+danosFOCP36TTMOg8EFWryrmmsTtV6GhxV+sHM6IOmnCl
cz0uGP5KxdwdZu2LeFOnC0cPJ2Ty2f0JpizeSXZBhK8h98mxOK8UtYd9H88RSfso7RX4TW8ZQjW2
SigzShMxS56a5u8P3tBvrac2DT9ts5pEgKbzuI7XKrNRbj1d7aetUUMZEOD+y6bNeQlpo+sERt7/
VlUCtbchS9Yo3rK/Q2hS7OdPslzqUvQ7LuuMqMoUYITD38IC4lDaaTc5XvSGTjfLFGbmiLkMuO3I
T1/CYIbM9MU5b81twjzilwNB1JNBpsKFu8PojE1Zv4mGDGJraSO0QCj+qvC5HJ/NeXeg1kcY+qzO
FF6aNaStFVSAsu9ICCNk+pJVq6GLobs/linRFX0U97pHjLq7InTuffdHQbhkEint88cuRhTLJ/TG
43Lp8JyYzbGMdtguluA6Rr+5oyLpksgoDPtt0PsnvbNCIr+O3Yi5xGTXPHMQh0RpgKyoCuNQxtxq
srD2hSwmy8036nMUr7HQveBHjmfg2D8U3hP+sCOWtrTpeY/G4L0Ymqt1UC7qBfsh+cN9sppsop+G
63iwCNvjyWLA/5PgjLwmTDeFUEIMCR7Kc1JX3NsSKiJVaTPB7KusGfEc2rUpvJAwkBElV07xyDlb
ApcBMAzhcGZu1n1sPxdRPE9rswB9L+mMVSSZ6IaKGIgDxVBIo3j394K5kD5jPgV/fR5b8sCxyDRx
BmwoZMZ4boMmDPhHOivh+hn7/9+KxU5oya1yMK2N9lopM8wLlyaMQRTzi4En13p+kIpELxU5HH21
X1v5a8+uw8sEss2AHg6GHEmu2Po0895baXCMYlKCEpjPr8O4tJwSKnEVhkyWudMi5yZHVwg1Hnzq
GfVTYE6eirl/LzKclXLujTcUgpe+nGuHr95CVUc0nGQ2KiRLcN9DXq1ptSwxH4c9BKWA/t/8JFRd
qQfhwrFirIVKVaY50HNM7p/uwA0m7/Q7DGMEJmzeXUpB8glFEiOse5LrwphWrkTyI490KW9Ny3Y0
/t0cwl00NQTTHbRfwUv2W3lQr9wjnov6uZoDYhxCPm7Ow88pXcCkl5d/ptnzQF3rJgFrm+GXfrbH
JX9omxfGHdw6J8KyqTjceZ4sfZWF+51n1TAs2ROOOD0MnNH50902MpuPpRNvR1l1hqk08OFexx5/
ClL/1aX0KGr1DKt696pAlz0Q0240EQVqSfL/5KObWVyqu7ntFejOmPgHk57kV5KXz96RXCPNwdCJ
uvOL2IqK4XHeCX/p+daxlI6CCyJQ4uPwbONrOAQeDhlG4Kx/bTTF25Eq7KNm9wCNMqIJz7PRCwq7
CbDRKrQ9KP/icFRr5eByHZut2e4Y3lXL+SDcivkUocm0rWAXOwtlXWgrpIOmzEmSIhqSXgcZj1ib
B0PCDUGc/YGEnoNQHy71nJV3McV/SPRqXtECrUQeheaEasPuB+eg8mEgx/xt3tEmWWxbWFlT0B/e
yHR3PwUdHO1BvRjrWGwnLogIdcvMU42GEzFH5g/Wrpft0H6nkW2mTG7kfgqNSBI/1PvWO3g1blKX
zY5NSunMaZagpWTakt6uxAA2rBYKGzQhus58VOsL5HoDeTO7kaFX8qyepxnWmFpsPOl7dxIaZ2zM
f+A2P2FK+Wn3+JAONuSWLcPNT3EjkOz8Q9ZhyCy9DLh+3AtJXI1kZ7wp5RKt1Fms5/62dR48eQsC
wPTgLaIugxTaKMJi7s55Ki+5DAjSxTHcGqHhlWQlpAIWwfWQIMosp8lersVdiBwCeJNIxc69cNrW
8xNBL4e7pdAxEsacmlDzeXz37zL+IxEvK4thGSifKZkfZ5KvyBxic8yE7yBf9Ua2jFDHKeHCTegf
UlDPM5/35wKh37Dswhx5k/Q+coqgDMBUIJWHRv4lkR7zWfxhwLQ/z+zooP0yZnoJ+2HgD1YOoFfz
RTf2KbSY6m/n8aSuGgVzYJnLe6zrwbFjRA4ND54J8droKZNyOaZOFMEJoOivuFN1qTk6REEq2KaE
1kpYfEiiDRYLLEiGPEf3RAWWOmBMoV9+ZsCMKTFI+J6aQxf2RA5qGU3waO2JlwPnSJBROfvKPUDs
CAt+VD7vbXRkk6Yie1MKoaN/ntNXPGXTYtnAYvjl4MKrIIS/tqAuY4DrMjpmaFxdVtKq8/FsUt+3
q3iWRD4K8O7tNfAoWMk8kU0lPOR1UsEFLndhuVQ3v//iVh/ZYlSIk5Ha52YfvHqILX2BFyX8pg1p
INdaQJOg363y4wt/tEFL1CPbpwC/u/m5FJo04jD4DYJY9TxIbCzKOqvPs3+wXzrIVfqAQdg112Xp
uQvAfS7yhqYC4C43xxOsFVNfNK8aonr81Jqrxckrp6+aqchCrU+u1LNkUslOtixv2VJgyfN1wund
SvZGFk4MOYj9S4pTXsEr6HlgOZ7/h12DfX2DSRIlk6J3PaEu1xsYpiWRSyNKsg1iOsQ+R35Bpgmc
KAM3FL2WX2YxznikxedSBC6NmrEXkjAJfuALsJWR2wBAaPsR9+GgY4R33dhC56V1AuTvBsWVDyxX
dF87/ZhzbkBvNFkHpsElzcAAkRDnXcARANvI/Ue69D1c4gvGf0ri7ANEdb5xZE0jtFVn60s5yfYx
97CQPTPxLeUOQeFk5stAhiFgd2mdl1Rsigo7m+vAvl57cr8KlA3evFf3tK7uiwSG2/R8lGGys5nP
+X21Hl/ZdhjB4/jTUxTvA7oMn6Z8IgCKtwh6NkzOWNIp42kdEVC13pcPCMTPDI9h5vkatSWDCu09
K5SQXQ52bP3HKq1DnE6rx5A7e+NTsxNgF/55jPvXIv7ZlXQzTP9GWj65fAvl3EC9L44wqqDoNP6v
eH95m5jsOtz8u1x+dwpmkovxSTBFSSX4mNop6J9xxdsEkpdOCV+upPhUh4ueFStFgtb/yaxhVq50
o7k7Z+qfvmU72uO0XBNLcfUIPw/tQLHhWxHpOda/UrVSXHuLgVnYmXC6iJYV/v+8nd/Da3mjA4Jm
JVv76Ln+YmgzKXZkBtZt4TwZhcKuf4QfW0zAzz5cJ2UTVN4AxkeqGk25DCsq6kuVW3ADgfgDfT+e
lUPmuE3bUu0emH3orhUlJC2bwRJfufUf5HXQfpuLDs7v3aWd05mYmZSUEqVJ3xoOpe5Oy1SU7RQS
zOnxAjnCoj2cxqWwip21ZNsze6t2KXVMe9a4fAAELXDQyMvXGv8lQQrTdKhUWO+BhjtikiIWhfPL
chenLX2yRd8bx5KA/Emn+dHKGqlZg0QjJ28JwmNu6QQ/OCflAHPYfw6hWQ/sY5KewSIExB5hmyvT
ch8nuoHXr6IGWomZJwVc95F9Nl+OLzknmcIj6VP23+cWPiGLatL+9NQK1rbh6KprZ/C5VTF5cKBB
Ny1wJwtjH+2EtMvVze9GfVEuj17gnhVGhb/v8skGS5RjFSZUdvjlIHMDsk9dlEinBqAGItdGmYMh
vhW6kmGVdzh4b+BYbcDMk3oc4OgjRS1gVb61e7fuEQKVnaGPhTkUWOZk8qyFujs0J0bxGiwGtRSJ
nq2Z5GFFcr7p2Gu8P9Jt7321JCGlC8tdZgAHyBtmaeAND1qGXxORa5VK4axj/pHpfzV82hV4C3h9
nf9MNgeYpn2Z5dhN+rnKpG1WwJkP3P9SOmtowRhLm4ttbM7aUwyHnUt08klODWl5g/0QhYG6Hh6q
rupGl09fka4z5N1Pi5rReRiZ4lRRvgGR6KKNhFeW12e1PzYPrF1HqfXodjjgyedvtrMvy9jfIhGZ
GK2uDHEJWT4BV4VjxDr+hAVQkkBuRb1vSdtLKGAtfthsxRjRZ8cvSluLzIgcg48rlCa50G1fg0Mu
LdWzh8lOT3r2qQ0FaXCvmI04KYUv/pFlChwvzVrzRvpOF9jqEKxxb2B1TVCdgSs6ev+SdZ4KvYfh
Dx0MFrc4pOks4rCkrvUVmd/mCteCbNOD3pMACInKciJvW4MRuY4VPyggGh+jas5hX55hPOZUGnHP
B2OpznwonTIAZvnwHChm1GMTFcWQjCAlqGIC6lvH6NDUUMTZt0cABwLUpk0BtZnBxOPrAPnrb0nK
cQZcqQWh9bC47QBh84ZZEQJrfK4rX1elGGVBCOJLabN6yP2hAjPpw2iCC361BFgmpcN2Vt2xntOe
NMJn1kKMrhhalbIQ/sCdgDKGiGkQdZD84LYV9MkwtmrIX/75+hGLQo/3SmptCHi1ohFakDOpbjFB
tfHSwaZmHNjzzfTlW2HGJqb2U173VJIJa5HQV9+xQo9N45+g476WFnba8PzfZgwtoNdnOqQu5k4n
FWNJSdSBKvRYZya2j6iGPjbv1asEyBvG7C3h1KxLiyG5shQqn77BlDorAobjiG83koZByhnU2kzi
6WDEDXAFGYirXErduFlCrglePx5M8iy5sg86tmIVzuKRXxp3hw8vIVZlWLeLSGId8wJlmW3D9okq
VbY3dsrSpBNB9pRPhEz6VWfGeKmL6vDYMIxsKWZL9wIxsOA/Bo/Kw+wYpaBhKsAB2m38m8I0YNlw
EnoKQRtKDy55LU3gRBH03vGZHjQoRjQ/k6LaUuKgIkkkWEeEiPyDVQc46xcEBDmydQtYFZet79tk
8g93gCAx1IlHTdIBO9l2K2aWEjsKRaWB9g15VNbfzQ/X8vfW93hQP5sZQD2D3oemXgTetQ4aNiZH
aokNy+6f7b7msL2HA2YrPppXCgDUaSiN0UdoivUvqIvn8gF2CxHFSCEXyqgSdh5c7KjGkzoShT5w
barcRDI7g7wTjj9ZoyuzPIbXNP3e+yUfuamGAqNqmxMOh+MPREgjiEihHu9NLBBhvDiyfkVz7qqX
whpHX0uupmtbxMcc2xpRRcr7tfnKJyJwXCtTEOIUGw8igztJV27rxh3CSnx/V9QETqMFIjkXp4XE
VA4ggbkGTliRqIDxRZEtYL+3e4vmRq3i9+Mmg/TexJ4rGGd1PRVRvBd8e4HUaqhxtPnIbPJYwZaa
dmNZjlhAxNmpCB6l5Y+gWoR7qwt41XzfmssMbandaqRg4CbvRuaZBW1zz1V0NGn4VvJSo+0qrzsh
BKU+1vQP8NtxyrUJ4MUAsHUBBFpMuzgRNXhjUsq1TZmI7X2bS5v3d5PvgE3K0IO9PUAJE485zH4Z
LMfugKQoWPS3RrTJxUhTCRD4fbnXLPTlnOVsScxG2ciaxHOnf+y/Szn+wzCnmbpBexKMOajt4uNa
Isvv20ClkC6U7+HfIYWfgbFxn930UegdEkwdRKouSlD3o0TnukYcIq3OzstSgN6PlogkMpHQRi/Y
7pfuHAAdJcn0sWAwGdOMX5TbGnX7JM0n5pOA57DCQdHlOJXQXajzBCQeFtQHSt5Q+i+96XoD/Uoa
ju5eFEmOE6/vBc+oqmHfu+W2N5FFQa4otj4aPOR4uZ0YFIsW97fc1gMwPFRKtAnU3BaRdrcPe5RB
IwuwpuRHy4Yq9lsayKnQnyPdtS1wPpM6bKRrPfrvYVrVGEfbotalFhm6rVKf3pnYjnVuEwPPR81x
alRTw9xibYHQ5gUty/sv/6lDnPkST7/WTslI0zVQZ0lDG/Q9ud14WwzN5k4iOHDUnnx+9gCmiEbO
YHslRQPRZQ/+rnhL5GKuZt7vdVo0JDnfjXu0sX9/N3NXviEcAezv6UJQgxuR+WFfr5iTbp76LzVU
r1JKNj2kWNwBqO9/K8GeXkYRGLphrppOPNgw83pEofMpyLMdktHmu5UyTDtv49MftHwnx/QeJbM8
QnwMGA+FSJKddn/jxzx3nHzvgIk1tAe6haHvYyhSVi3t6U1XoX2JuSnah73/LiBAeaSeDu563AOU
QociKO5Sx75au1HmAC6T12Y3BxJH1QyPZstx6rMH647G3EwGP9BYWGD0KHgxHsGIEqu42LZtxilX
pKWm7fTU1bdvhDFHm7LrnKmEQP1PBxzLTu8egzgBtBS4pjO0466xm6l9WQxfY2ST8RdZGfmI0Ed4
zPnAqLq0KaSwOK5htXxieqNZUh1KknTly6GeUNnfK4iI9EVgTqugUyOl1OabGJqFkNfzh+r68s6n
V9keeKk7vxEX/zVxuKCgLzHMfDcS08f/drTzR4VJtszrwswPMI7GDYMJ0ftPJA59jLG/ZVSrkygc
m6+nL4BZaZXWEE/Owq3yeQxEBKO3FjIKQLtgrZYMcDgax8AWEG7CNyr74sc1gAJePo1BxjCdMtoe
c8CPN1HarWAgDvVAFIfBoJK9FXz/0o45Ew3F79KVhWW6n+IKPbChW86E5gDEozKKv8G4kcARXKiX
Q0kEwqmPR65Ka+e7ULsHl3v9zDxqVn34RG7p0TZsctIEtZMgRYLwGDDwnIcb7XEA6taNh494LDsE
J9untNZExSFkI3kFbiSTWvE1joT0OGu5p87t/mfQIMb9R8i+HuJWcLPCG98bai+AMUVyJDLNBPtJ
dcglHiOiDZhniuKqW20T8ynQr5ek6652N5i74ECM/nlOJSnlKWmVHF1a9+QFKok6Ig5NBoR+hbhl
O2Aw9x3PjpJKbFOMsfHSopMQSRi11LcXaKm7MnFVHdj3rmEOYPjBkjxkaVVcWit8G/v9M3I2iQS1
4+UHycwVt8MXmkkwzQt08LPBTQ9f5QYjOJ4606w4bwl/n4ADsMsTAhk0Cb0TN49XFa/24dWbGW5A
VBDHGCLHhE8w4tfM6boQX7Rs1gmHLpeQ+HV3UwMmnRdffZAuDF4JOX0bYFBW9s5KjrTVZNAergoK
XQs1HRa1+Q9z67xlGjPdQHDshKpXizpTCGluOfajbGEa6G9GbujaQfJUTn0CFN3mYtfhNl5X9BQM
5Z9RC1lPc8KsWnsSeunm897YuWk8GeD8FiOPbp3jjPMEq5zdlpG5FRpGhlK/Oiuo11MFE5HXho6e
JbMDKPjyYltMBc5lIwZOEadADm/s/vA3c0G3DgmhSH7404P5H2n6Kc52g9amgdIbjt+el2rrjLYY
X90L0Csq56Kk2XeLrrXuCSwVBYqGcVdzP5SsMIFt8JQt+INT6h9G9WellP2LfVeCvo1DXGTMw1Zx
x2F54H5LyhOjg8ha6yFradgFspcBXLUYW6hmJF7g7sOuMFN/nC7rqAniE6XQyscX2/vLjVZCyONE
Lf0YyqwhNwHt6u4cvblr9cPn8Zqf3VvdrF56cDcQcj99qzELM0QcEIKZoNxaYX1+oUK5ios+3n3Q
kmq80nBpZPGS/nkLf0b2FbHR5eCVxQFP9QacPQWN6RiNA8U+XIko6vy3+WDxLT6cempAQt6ZiDng
tO/Ktw9+SuDJ+3u+9SGAn3kGGBHZNj2w/vurI5sug3uVBLJUAtQjXN1MVn3CY1KuSZtBEU/m9Mxy
aihimcyBtYNPPhs98ELc1WRIcJCj5isRrPRD6jsH17oERalc2TwlsK+SGVXagLIayERqWXnaZRaP
FIsJCCfXUSjRFxEQtBz+kSTACp4aqXomoynv3IYJ0KkDmZDzLk09Bj1m7nku9NZkTl0csqwqM93j
9/qgD/vb+5ZE4Gch+YS+4S39YBybK95kiEcp2vo6I60Z+VJ8CMFFdDzpegqIkQPsdMj4IsLvPpNG
1gtGE++QeszQlnACywWMEsoX1jWUFh4GH99S0RCwfUqaJNRs+04wnQZXGWKfM0K68zqzWQfvPFIp
528f4MMi4DV9dMWigXT4/gkz8+A1RuIliQnasbFQilzIw4/rB3NlxAo9nYTRAXY7liB73QpdHxQv
xTYeZIccovS4qOFfIRg3JVLLpW/QCaLWcUjsBymphGM10lFMPKIAkWtqO3Q8fVy0icoRVEKZidp2
KWUMxI+W98F5lXg4EwsSf4Cc1SnU6fS0qg+F5PgnyuCBy1JxpqhcgxXc5JDS0WbVxTUyA6Ssmlej
FoY1PVmyOHan1Hz94LLlliWrdkSDkBaOJ9fYz3Xti0byv+yoMqjYrOtujDADQI2Gz7FJleA9eG4/
B64jZYUbuntWjYj0uUXDQGA6uIxbyG/GmzR8CCplWOnIsk2RGg2XZxLW+sGKIZYZAtRFs57gpELx
D9a7SH071ite6GrrKQzbYkVLqndkgRynOefEAwVCU4f6h04vUkPd/Kz/23pEHJkE4BaPVsdKGiIG
q5+6ob7NRAo7nGUYOY1eCev9gYRdgOSD3NOxYKcDcCxDJZU2BSyK/31FF3jk4Iwyxp7LBajF4sP7
6GxbtrIoeqG5gvCyveh/XbHIqRVymGF+F7sdAryp//9tLRYoiPJqn4bdi1mgb+YGejXZ8zxi80ta
tBQkQRxII6BjH989pbYa+KPrNkeIgXA6dbkP/yy5k1PF5oroRbPCA7g8V3X7CSzKwxjHYMMR3U4v
UPbBTz5WNQZOG5hworAzmVlEgrjlRHdPWtbsMDUt+xRE45T4Qx70ihNnSXpxkk5rbmWgF8dWz9UH
4RcF5euZ7pCMGGpibND9pcHwc1crqSOeiXbX8elEboEP2AoapOpAybcDXIp8uc6my45UbXPL+4Eg
IyrHIurNCFw+V1z2KIXYe6cGMgmYJJlrDZJ+d249YVqG2VTkeWGCVZoftJLOmsyYyI2EK1kqQCSx
mm+Swdm7iYf2+3tJyIDjURZDwqSkKBWV7by5ZtJR1nVzU5188Jp8mXpUgVDCRNvclYm7C70OK0md
3mvJ/TaNkQLENsThkZUIk1bYuN6wZJjT2p4q6l7Ajlby58vPlVoJVzhE/aAlMXc9CfN0gY918O96
9dsYMGxkbvjvQbxFvxXaHMfV2ex/UcovQuuyTOoAEzh+kP5hKWiE2TXIEhG8D4pfTvHjOc0BzenO
2JFAl436NLHizoxyxhzsRAC9rWi2CcJvCOuxYM+ZFQv8oBHBCpu/++UgEc2J0R4aae67gaNUyhNu
m6GMxdbeTS2JtXQ76Dvepclvjz54B2EBeVnJhJXcacOMTFNTG1dIDxZgWSOHa263j+hmhNEVoEUK
0QVRoNKX0LroXi03tciwAJCQfTTTm5fKFjDkKTNU+voBXENv3KhN8YeywUjfth0ZCyhxDIeCeIgc
52jHaLTBOiY5p9CJa1CasrXEN87aYV9sCH9DkeygDHK3StUaIyWiD3MnTs9NAO7R0lBK6P+jn5nr
n/rwTLR+SECWUZyNPm+SqurAHnk3pvIp1ZIm3T0p+UkBuGfI5a1nnlmdMY3KmVPwGTFbkvSN1mVZ
rR/X2kjjH5BpZIvjiiQKXCMGXNqPbYWXuQHTJOOHWu6u9J8LRhSP0GfqkIEQ1RKdpvhKxKXYFwr0
tQthSd2olRej8chp2i4umI/FQikAufDDXcEIQO+8kyrvCiRTVjnZ9NdibtLaBUma2Gq3oRu9Bke3
zX5U9nZWi7FEJSDa3PYVXUsDl/avKUxzoB95h/vIyRY6zSVmZ/cSzf8hEgzUguSbHXwBO1BKledl
wd315azO8kk55epT37BV4QykOd158yuCYmj2dCWm12vZjNS6yyxCzQCYWCwAAzZA/1sAp+qsuC/t
JWcsgHw4IFPT9wlWCxf0hAjgKsSM8mO3oX8fC6JdqUrqexV8LT4DrJv0MjZ3ZpORm/92AJ0bpwMc
JXYiGtDjKcON9uLMJJeIR6UfjsnKRfBOGs5Ewkl+LbFycYvqpob5x7kbRaaxBjvsRDelIcKqMcSk
SZBm25IC3PEkQlr/VRYSP8zSI7zMzbWcpN9XI520ejjY7TVu7DIaHZUvbjB6CD224NFPMU4mIkId
53XVqrA9oL5TnAyDNnrX81tsgxgLtcq7CIdAPldloCZoDQ/ChEQgii7P/h6+I8Yed8SK0NxRAvkT
nZu3cnKVFTYVuNnFr+q29/mPhrTaybiwXEnkP5OJT42yPHYDRfSvM4S//b5W5KO46eHJwwfDeAAv
SCtWSQ9WVsDlJOzLCcgaKkv/kMBdtM/1Gj3Edy+UFA43srXVevwu2nWrM4u6Gtbfoqjcfii8OB10
lN+YDX7HO5jMs5yIOg8+3h8RVNQU6PjsE8BeiPaLqbLA+KmiN+7BADs67WymtKYn8id5PpNYWLBB
gY81afZmXT2hWEZpiTAzBNHfgUI7zx9jFWhkGh+yMsKLBGW3qMOE+c+rwlsKwxy47ArxFoXtcPNR
6Cf2yOtHq4zCuD+1rYkEEJ+DUfe4caCVnZmMMjwpNiUPMFDra8rMco4NgsB4mI9TxJUH5BoYNJED
NDJihPaRxVpImeUVQy15ZQDVVr0VUwa1MK7zhtJKuVwRqKlxLpALzLbXeahOR9sdJ8t/JxUrcFai
tW+sdoFG7Sy2K41Gxj85i84gi9LnCZ5870rzwN/MCz1vQOdlcj7j8lbJCzyVgpbGrljr97GzW0Bz
+ONoMCPam6Nh+VUnRmSdN/HBmbPWPBRI+taK0OcZ/Y94MMKhlDsbuA7RDDpfSrc+FdsiyLlzj3OS
Po7OE5AcfXCx/WUN8ImQaOwQyuxCHObR19dMsNFDs5JIgOp3acTeWydL65Hf1ZwNukApTus/jUsw
sP4oWo8djD0Hr0107z0siZByKOcxDm43SsphIpOhf5xCYsW2FG75qhrxY5yoxuyVuM3vuRx4EkFt
hUjpYteLg5d1oMrhHgH57eEHspMdItRzb2SEK5+W4d3w/58gnDwkJZHxak0h5Pf4LS/xrqdRSZwB
Wr492xCWFfrElzuEOgLUeKzfrHOPVchhGp/1a2PCv3FnR7+AaOKUeZeuBJXIqm0FrGGRPnodNhbU
r8yg9AJCvBjJJnoHZ/bNqcgabkW5JVnrhYiDNI4N0ngMRiIWmcYY+zZSAnOMAtDJpOWTxondq/Zb
yocQ18yUdzfs5bDKlyMWUI1hcNyEXwn5aekvSQUIMpsk9PpTkIN0RX0oKKWHtAbps4IUYRd0j4FH
U7lJnbYOBexLwFlf0W8lRrM05DFE3CY8elXiQwLhv5z5pExpvoIXm3qHclyASfuqz+2QCPMKrAN2
5Ts6CHAAEOxGaRdLxcwJK9wbTWvjv2e5yMjxWHH4V1ckVnKgFL8Gpjy7rzZuMsjUtglXYj8UIyvl
V+zZlrtOVop5lt77l343eK02lq0EdInQcQvpMJkawVlX0XlkexYXxoLQC5z+rK1r9J+n+O3JtiLc
qLhNqXV1FCa4BpxA9m+/m81P2PvweznP2uk3HKLsshFYW/vIL8/7RCx57+DF2kR1Sx7FId7Bsgiy
3ZifnHDOEX8rWcU85UalPzXhltCKnGs9GUG22DVH83DrkuOjD4ZTzESXfTddWCBY4HqnX1P6fJBk
e8jg9WVjLZgvyNxdeduRjj1n9M/BkxerIBctlGpE9n+YXQVWrx1guOwWeAoguuT5KAwRrJ83AOU0
o7oyoVAJwh820lrXUSj6OEy9KKLtBhHRvq80euh+hOdNaB1rvndlG7bs0xM8ijE2TcgEliIcKUAq
Tr58PfnMP48SjpWGoxkD0EhEtrd3BNMuZv0+7MJaeeoWsw96jQMCGCQZmaHl45bd74rG7jHm2DwB
5a1t3MH21M46T2DhTRUUoYdTMxTy5/jeo0iMzpNUeKVTyULfnGrzFU3QTjDImG7Ywwo0FkLHDJ30
2eeml37bKCe+PoUDmeKXpG10JehrAF/Naml601JxjYq4nLy3PfK36fdYuDZ9zqdcrGnhfSWeLRqQ
oyRjhve1wviJ15j21onmaCBlvgEKuMdk08WJCiBybUWHTs46AnYBoevFGTH/T57hd+TAZBY7+dma
9LJKixDKCinUXeKFOJSU0gAFpJO6jmabxOzdq7nUPCtvUH3WsEAx2v2Ae3m0CN3PJwZfM8wHjR8E
CXY3oTojuibsrL4y6Nl1GDrUePa57MkYxykjnAxf+n1Au3+uyN7UsAM7qvH8TwhfcE2vljIPRcPf
UzDWWDob+QDfnV8BQKHZMLfjrFww533FRfEo6ljcMkg03OyBFiY3yrB2dnQDx3+TxIT25yqn+Nzz
AuY2R+fGTIOjFWUO/BUX7DPvmOrngHVmRLigYgfNaG0ul7UNAs2h9niN0dm8yL7wg/aen59KpUBP
obZrnfKD6jhJPMHXlxOUAHo+rUqTySrWWhHjjwQPsWnl4eTKg034+6ow0CfrCasWpG4FxQvG08cA
fXJrNLCl7mcDlg9v4cRqhjgN9evqB8oW1T1+51rzhxz/C3QdUXEb0oHomWZ7Fo4RSYVckLlZDtuE
A6eJUOMMOhFcYLGdXDYobM2UrOFcmNwyr0xNgKGXWgClQothIrs0pEdbLX+vwvhkXHQe88rIPSO+
5zBfcmTl2OqCR0Nm4lzN5EQIMAp+ZAHBhQEJFkJ39nhuKsYnk1aEXsoZeIDkZB+tzn4s9zL2Ji8C
FYNFTM00TwTOCAqGSBNBklrvYSNzIHxiGaQktIr2YuWEBjElgvNoXuENmTXSeWEgoxhj9U+bCV+Q
A/2pfRp48oaL2R362A2tqTnwt6sLbjAXaXQIWKOlrzzs2WiBV+C7dg3bhynSTvOD8DcjA3JH78GT
geL28wl2drHFy4Sk+57LECNo3bZHRZkzPPhW2/Y/4Dq+Cia6uwKHXajhNzK5OPJRInXJqWi+zwAw
x5nVUm7zJ8ruH3XgLXQJxUFAQs8h1bMP1SfnNq+CPeGrKdH5R2b3rB6dYYbVmAEOu+M1TmDvAwWX
3o9q6FH7y3GCAhQTN15FNK/JLO7GlltD+crIUZvVRPhKkyF1M7ZPuIhxt53RtNm5DPvkPvg1Rflx
5vdiwmvjZYzGzazhQsigQtL29j2BdcpOmjhyK00dgHtqrji7wRTw6ArApzrL8HLfykJeBdQ5N0NA
1PwuF/yMmi8O4ZZcZuR+mh2UpQ/w2Qt7jSiKbU1zFy3bYhJ2utXepkzX+p+y98nVzM396fEvYRPe
NMOWOwyaxlwDdqjKSks8uawqkWYoyEWXe7TgN0Z0d3b2P9QmveXa0RCSS31cg88yC+xMSnOBPlP4
TChkoyPs+QlHq7pcx0J/DdsnLmd/NC/1fxLB+TbdZoPZF+04sAesUlTXJJomgwhhlnmzXw7ZPA+L
I1IgVel54yCfAp4TuxE8eXXCgwuhn93wfSbIlXk2dKOJRUpxNc3pIvbD+yu8YCdAlK6iQnMWdd6O
z3uevoTMG662TzkpDuLM+mgBON7cdufufOtpNUsHaZqd2t7PPVDzsjm6wWO7frZv65bhxdZ0s3X5
Sd0R1QmZIaO/ugcZjY/mlpf+SMnSPYTUNBUV8oiJpClFQHsRilU4S0HT0/RGEv3HghDnNGFGqfbC
cqO+k0A1AL0dUVhvZoBTleJIC4D6zdVztI+QCAhK24QZfsksgAo07AGVevna5sRFs6bQnRly+aMX
zvSY4bZjQm+XbYw8CL7v7th1zswgKwu9/8UfOdnOeGYJ4c4HpLbMoTB1Umo9M0AfWWeLB+TPL7uB
fJ3oVaD3PIdDowy4lCMivKB1XKLtVv67jk2YWbhvrcghEsfgm1Qx2qM/7oSal4nxyM0n+d6RZ0S2
62rT7KFlP4oiMACLBksfXWgk6fvPgvXt8iSLJz/7anU5d9wjgB2g2KzuulRyCQwyOkRZiECLWtxL
PvwyKSRX6SAYH35LQOKGextAMnuG7aI0boJYcJ/Ruq++/o3Ma/QOspO3Y+zrgvcWMY9Zc67OvAZX
2r0BmVivfohKHKjq7BQfRBZ5e+hcgAy6YTwX/GL08+LcbncHSIE1gsWI7LhuH0jDC0Wl0qHEZkpm
baXeQDofNmdRf8VZCXvyd/gQHrBjsUsgoqKE33AhJKxp8GQgpmga7ZQcnCAhxgqhd3cm7hUi9zKT
XLG2xKIFhoE0+txvMFUqYJ8BT0IfodWvDsF/Wh24kdSBMSRHr+91wqrwL3wuY4lqpThY0VOUbt2S
RJg4u+DQsVwGQrte7TA1aiksYOpICAlkzIiudpUexad8hkzH7cDUs6BMD3Ygr4hDz1P47I1RBOYj
0+Q6K8Ip+qeJn45NMN6ST42aFGXiO/vxRYJoLSwgxTKhXihqy2keja0bFvSpSv4zOfkNFt6Gv/xC
lQCedO5SiegkfUENsXjGXRfvjNOrLmNLXay2xHDqHOJqoRoeLQQwLjnMa2R16c6kfQ8oWJFPU/ck
lm8k0ETubedlWUzQk31MEH8fJy1IZbvbn+edOUHnzqcbMl47vAb+LFmnm3loicDansltej8vqMhs
e1G8pVtMshURK0eiTCYpGgybs2P2milhFB5Nwsdpe6gb0sUPtQ3x/TxpOS00n5b2sbfnkFXkGqaG
0Mm2WVljQG+8udlp38B5r8rx7u+F/2uWhIIB82YZ4UHcDZTN1M8GtM5MmeXyK869LL7tTNpaKyvj
0dRVuf+u+blXtSi+kzqKUfMvFpT6Rk99OfXbpL8n27i97DPo0OUQg77W8mKk2OK4w23iro1Dffs3
3ZrlR31tsHpYvRWVHYkgoFDqDvikWTdiICzSqvPfIdeTyeShQY2xZQfvHrjrdM/fIlp5DOuHjACB
vShArMxLUXXRmQabM6pU09dUJ72L1yUTZrcWM+PPgTZfk4k5KGA9da+EDd7rWypOSHWNeGfO983w
wuKc7BBKDWTIQ2hh4QRsfv8jT0pJY4gyw6Y+sslcLp7cyZg0kvwkB+boU6eCJqFIvFt2MOEbPd2C
aezx1VQoS9/Ri+bUSJzXUOrfIjXC6OK53ltlkEWZf5uxdrwtjIBGmfzll7xNdbB6/+uJwfevV3mA
0CIsjjVBzEr+9Tywz8QFDX1y0XHPSgiBo++0goO3NWC+uTfJ0wN4e/FvUjaXuJLNznPZVR0++j8M
A2peNhLQvvoTxMhPAxjliIWPAFcZFnm9gZh1I25L7ydhgMFouwiq5WaukrvsastYuZgUnM/QvIwX
lcBRpJLUDvi+bVbmSamDj02ERpykpnu5i26SOmAeqgrLVt55To2g8aNJG5GcLsnEll5ICK94q+6q
X0QCN+F1lTyBiYSoNTmO3bgEzhWKOukYObOaqQRjFTyxBZbeXVmcIFU+tbLKhZNa+aDe8S7M9gge
ZE5X83+218LrAysfxYYOO1TpiWrloCGhAjnMWSGcu2Y4s1bSfOBESh5vprbayIvfDVMX18c+5g9+
mvMSd2mGis48hKuasiZBzyQ4XYqu224V5SuvEXVuMx13RRunjznn3UoXa1W+mEhUcuOLvwaz8rD2
uaakSn+SL6lsxpO9X7wlol4jJvFYiH5Lmbjpm69TzE10fsDVfohn9hgzYrP2BYHMfPBrXyhEk7Eo
DxBOZPmjzysCDaGKpPHql4aun1PfY5J0bXMzCG3/bSA+SgxQo6Q7JvUUq/w6CMo0/IOU1v1WEZ7k
S2MIW3BTo1GTRGJM8bR5GjlwziQ6K5DWt5XIocArtvf7wpLKTimhX4T5mmI20lqHXdOUUoftCd5X
1rHdd3IzqxWoZ8En6Jt6GLFz7flMp0g1zkWgWiibeWmxNwDlrgI+7yZ21FSUKy43nbmox6AITnMn
Wzmf7Dtqse2SK7QQALHue8ASozLiw3aKlumsDiXptML27EcS5I6ggo80Q3s+3wLKddOXenTqdje/
XvzuNpaS21ylDPqd8yxVk/JtOhf/g9OhxoMgCHkp/QZEi78xwHZJW6nbIeRVVXIToZvLlU6kpIdo
kCWXpK7qJ8HXaO45jkJTWNyfUKzPZmw39KTYcvJmfIL2lncspJQ6L/KFosuU9vZNoVQKkUrcFm10
q1+TKq+jHJCMXyPskWDXgsBI6jWudLPxtslKrgJ+xeGnhfMAAqK0yD8pYhH5G4NK19/bn6KwkKdm
7TqRXBjskRAjIr/MW7R0e2FQfdsiootPc6bZ0WrV2Dq+eoP1PjZDJUv6UpjROFCpyEgkP2c5W9Gn
7/uO93vLY587OcDIT0LIdpydgC/a8kVRrA1cOT3epdHPpS3kZawXPRyAmSxm7IW1uNsdyx0kGM5q
O9wrDNKVqafvipPrrEyZ6JcBKnH0g24m9TVb0AAok3TEAh36hsUUCTqe+bjvLK6Xb8ARjzsCzT8e
wFdOZ7VZO2fUABFMgjmxF9raVSQ0JH/3XDeaInQ8smBg48CyBu1eYwGevyz6iKRAgPDCJLGBPi/D
V4+SgnfRD7nJP+vxd0+PdA0cfqjPBz10Nia+EjM3jlLaL9JVeAVxVqg34+E6rsZ/a8FDKRwojZ5C
fmxZZfOKZ5yi+19/cNa1Blu7nk/z+YKWbFlnftKbe+1X8X9Y0EpQmseENWRox8Y1e/i/uVQNjglI
YipNiMW0jE0PH79718z/j2JFJ2gPmSt45CpjKfhzWsuk9MtXZeUMTFwfFBTlJCNeNzT4x/toxmBS
/A9RnKey+7MlBasxtO9b+HghkhWvgcd5hQw2EFsX+p8cqVE/2Jc3XacdkSY3q8pHDL7XSLrXerI1
zwfpc2bKc4usP62lHCMiuT9hcduibBd66mvsyLLMKPky3LnZBGiGQ6vt2lez1r8nLjjoTNt+plbw
VQIOlgJwtfqJkAUL0AR6sJ+JGnff0tZ1Sx5KKlcGLkzUS7okYCcBNh6MsSi5QDJMfsPKpmYkuAk9
STUoSeM7LukWj4eOQLmjzu6DWarQ4OAtCvENPQdcnn/MhYyuiqB99rgPHd9S1QetY0P/BBdpgNM8
/uln1RGaz5DKuLnxJyaWFfsYRz2mjhYjpWwYzULkRcZbGifqQvPpLgKITVeEulse8BcJQx264Rll
rdgOplKMReOSCZYWFVfWaHxi/1F4F8UEPQ/E5QnVjQWIP77pur62XpzDiYgEx3FG1nw/Wl6lx7aG
BZyRc8QJeopOheiIvTT7aTpOBb5kBffryc1M3tRIpeogJN5D3hZEricuLEqG/x9/XWwtkcMVVzDT
zKhOIprtPU09OVW6zsFIVKEqv+jefZE/kbwVpCiK7ZJfltnaLC1ogC/ZpPiTFnFB1qLpfemJ7wN0
LWKCICx6S9hY0Q0V3DwiP4VabtOrHtg5m3VuXj7EU2HxpohTkkElZBf1b3/Yewotx8t6hqugnZpK
zi582iBeiv2nFaWxuCjn4ODyz7tZuIkTw/jLoWE8b9hvRdRRDKvDbb9N8p4k37j9FqZj7v71Fqqw
xpDHzvSDu9WLCVuH7Py67wIfMpVHbzCm5Inr6OwHdeGhSR3rrKfNujM1GNF4YkO81+mv6rqVSUIP
LznDTNm3h3lrtldZ/bOh3iwIg3wnS7oq6EZrb451iKK76xwnd7U8hiA6wdhQnizaAdro86+Vxg54
bIs+85pKnOmcPtoWJlvP2V+dmSiTSPT8bSxTkfpFpmCx7xfgNF4BLyBW/UVLLRJeXBR9EBmisRd7
qKlJInALPiw6aRah9Srwg3/WMpH4ECm+Kztj12YHSatYCKFGbpWuSq6SsixZke7LZadimAPf8jNg
qlizakDXImG83DKA6VljrLbNYbCG4ZlHlB5LHFqZ+HozDGAdj1pNp6kppjRFne3fa5jBW8aD+muP
xp0OB3CUqdwYQtOvXtKC38nxMt5jcJBnVxkVayH0wrrtHeGINH13tl5fFXxnFJEt4D4I7xwHSPxP
dEKc8+Q9MFauXmdit7SX52gd6xgcWXh/aUO04RlcafapqMmbv1jfwTIUfosDpGY/M8IgqeD+cXPr
y7261LVEQpL76pVNorpZiVPMNPDp/VlNW9NA7RtPe/+mQ5Tzykum/6JqEHhOBz6RJRkX0LeYIB2O
GAiqh0XcxFsYZDfTVvWerU/Jkqk1Aqc4kkNohLZ5q/Xi1+1RSwDPgxv5jTytVgG84MMNPr7KbXac
NcsuUfIuFdTj8Cwdr1bxhjw8Vb0BeObITlrdRECdAfYbvSRGSHzd1S6qWQpM2l+Tyodl2fOalv7F
1iUlsDk0aIf3yPGDIiIjzys8SRWbnSlf6Q4yZL1O5wJaC+Nmi37Ob9qn7dyUIHYShtUJzx8yWasj
Yp7UT0ZbT8D5pBrk9Mj83n+dhR5YWCplfJWQDmdxwTsXkO5TiUVOnUFXgbWB7QPF7DGWlyxEhYlm
EIciojd+EKIwwgdlU6EjU60UcKnRN3qK99/OKDJavy1T2ZeWGm9ku/Dyo4yROtXx67kuGAipyjfI
98tQo8CRltTKtfQXmt8txVE3j0F01PnU2zxkrV+9QQQpv9tk4HzAypMOlU31wzHXygXBc9NoblED
JQZW/DCSI0EvdSZq6danCO8XqbRZfyuBeWRieVoQLk7ge7kmjkdCEB51EPGZzLpJF1DLEY0w9DZT
K48TAeI+1PsBmO4+AWSwQ+FwFSxjzYAWVzbFOE5CJB64J4nOrk1SPabOzVfUpVL/y2jmqjllZdGF
c5PyP4jIj6S3J+dpH7j+kLu/7wKeL6sdnbsYfGxZcttPTH9oL8YJgF7r28BCNP0KFXNZoBSOJZgX
jSSR6L1Xjqau+GQiFwLEeim9I34C583s7qfZiUurPIoQbume2CFmBnf2c2ZuGqfvvjMUF48Ndl6o
b9cGCHZmvWnlYrHBrZ1pSzJB0U74YdvwuvWR8fPh2cQk0NXNaSqxox/tb/GmZhA8mDiwuB7srG21
zOMRHXn4nNt2w9l+elP/pz9z2csA9wbKCNhbkGsUUpMaBQW4AWCO3v2PHDQkDzR/ZLreXv64Twtj
kcQwN/KuSs/xu+Ma0ZGEcxmH7MzQERv0mMLgvUZpY0ZMIOUWxpPsfbJD1hPVMIl0qCaQMH3/TJdt
NSIicdrGjtGFOO8uRHpsPoEJQNysjQ93gpieIgtXdmUr+JOQPpPlnlicHkr0JMsmgzVlpzybBMDu
B5z96qyQ+GTW/yocTrnbdKfjrJUJfIi2f0u/KUfQuFzHbOe78M1XzkBWL5DKGjFxOZA0sTXWlIlc
2T5PdtdEbV1+8Y2dZhcODEp+J1KZSItxbbSEW3u/UNVAAtNxpCnk/Ljb7KM8nECfqN5UOu/ta8io
HHLMhmf/WMgGPkCgoxBz9bDr6IrhDUX4asy+Ia5RQ40OzrnpIGcqkMnt3VGW1sdKkgensfLf8HH4
h8friobslhoxC1uk8AmdcIeYQn4VxeoxA3IGAaeVMEHtbOeT8qTiWfcRmyn7SHyCr7lEof5sqM8S
jmB5qt8wmEKrDZdN2MZZuUUsKijCQeSeoh8LebXl5wYXo5Kpmx//2yg4arqeSlvmKJzJ0ArbwIm3
TzgqaHCWJ7lWM4OeR48AI1130U7W3snRxG2Stux4cmI4sKaNqY/9fFojw/OhNlNbSuxOPj6FcbCz
AyhDzC14XMx/RF6G8cwPZNNeyxxNzwcNtGnjNDPG5PDyZo3DGKArkOaOWUKmzjB2lVgtZRXtYzQY
Qwa7ERJqtKcM3GywFImlHGqzhqIzZy2xbkNtlUs8xs74ljJnkB2sZ64g+08Pn8IWkdpq4R8i4F/a
DqyjmtZlWNL6cFIUsB1IJN6rWkH7Bd2i8GiIGtCaewE8x0e7lelRFxfhB7BvwUAe7uLWld32Tisz
Cj6lbxoamMSP9f1sHd1NuAN+qs+efcKkJP7PjoqhA7TnXK6FeDXwXlfqpgePDOSieikueLB+M7H6
foqToHro/ylxIhjKMXKK6O4xdLQLh7Ahc3LbZ9XmTxsD9wxTfNOHkzdeCQllSD7MeDwJhyJgzM/4
kNsGvkPp72MN8dm3H06fSt2Caq1boi84u7DCONCEMSKSr/kXEwm8rxSOqO+etzGOJB4mkE2QUFgB
AV1P/n8ai89LOlpWVXGx7O7rDdFB6DA9E/acYyN39H6EdlZ1LbYZRH0iusayQo+HFX7X6/Au958k
hB1sH0Bb2y6ZkrdSvjBk92+Dwsol/6Eq2bWenWIEARkpYOCv938Hc24SsZzuJgLGosFbqo3E1uhw
bYHGGoKBlXAFNoKZkX6IWk1O89sGKE45xVAay78GHVinv1eT0rBd3b9QBEx0YfeIyMJabAzu+GSx
rSGIADcbKp7cB3Dg5zG/iDm+mGRJq2Lqb8V9npLkhpyLR660B5swwKwq6GBK9rjawBf7qCcDX9D/
htywkasafe7ZEixPlljQLDmCkP2Z1g0c46+CYBMKMPWpL2DE0PzKTbRtcgtQ7vsRnowgjlXLunxu
7m7vYe5CfD4jQBNSfJECLl1UsPa0ZVPzrUn9o7s59VVQXDdsFae6PeHjHVZXRF0po5kxEL47cGxJ
ALhobI2/mnvqf3eY3P0L/4PcFekMF0eNzWYYFmSy3dc5hTjdJpP7bpwXk+mC0ikgkrK0/FGJ0YwT
UgpAw8JKbHwBHIbhBa8DvGWu0uVaS8J3HD9k+1av27zDxrCS2mBmWqgdrna7VWrjNN56oUFJ3pf5
meiUaid8EWfM+tOZRL04OyxOJZbOVopmU8vPDh3EtdhfwABnbsQWrApFE6RP/hmZY9Ihu7d8mu7l
YE7CMA6W0maP20E1om4NyfftTGsegWKGboaiDQH5KIRJ63dTxIhMR/GRH8OjKEVrtCpCswXTkAbl
OdR8IZVVDmUTn1XUm69NvCa+rof4/rN5NnOuVdU5ffDSmU35bLPPazrJs9iTKi/tD5ir4ptqf2tj
yspXXrNmlxP4IQETbR80bDLSuwQoNlU1CYndFleW4LNmp3VKwjwTHPSalFv680ab/Gp+f2dfuaOR
RaoxPva1w+F2DCt3hhYIJVNh0MWlnpb9DnBgVaYlW5Sod28IGn4kIBKACBtuFMrkGY6TXHcXAn3I
Lu1uOtTt34gY0yh9NxyS9Z+K4VjqciVOeHMLrFcR8pfwJws6pBGVEq1q5KZ5+ASWFX+6VcOz8UYJ
4UJRTCC1YoSRF/M9FEj6fC3iTQBLpoO+5D4hWYpMy2QCxcq8J1msu12HMg/ylp+G2ichkxn8XITO
zpuFRPol/M+TJIfk2ObLxyArh+G6+2LgjlfN98WIICLMytfXZYWSNfRL9fKTp7dPzK7LKRIpz1EI
wqDRn1DZGLgfYpdjBdkCaUMZq/VJnPyaNJig0PGLpx79+ZwXJVToNzbl39OrgRPQZGae2czjJ3fY
85S/amAmua5/Tl/7PYIRdAwvEKnFtzmilGNnVtWVoo5soGTN74sF5mTo9coXcufvkQ2qEoUgkMjr
DbGc0bU7pUYTy5JE4dw3IgLhjbj7cuujLlnKGcXsWEbe/2+SHIUsAWpmu/RhiXyibaPmTlwsU50m
YdbJWE9wJyerQBefH5VoTL+Z7SQCoLbEexJ+5dLfo0j7/2iKnN0ZAQgg7hujZrLOl42CatqkKf4K
YxjdknH8FEC5BgPj0pHGLovg8sjCVb1ZQAhWbgz1tCo3DIDZoUFHc/U/nsOETw4tdz62/DRKT0y8
FNiVAtcqNBUj+LMl3McMcbarcskQ/ltBtLSr5FrVTggjGFz+MGC1udZ2ZZTkIyJDAnXQnRBPLdyN
dxg5cE8k1n0L7VzYJYfe1Tpqxp0yNKrK1SFehHYbWnlvbC92jAFKsQmP7FCz6k1VveIW1dUDckWK
S/FLbpDS/weeCNq6i4o70dOwwwIMMs3gYm90LH2GqHxljAd/A6KI922lxA3rOTy7g+W6aI+NAJOM
w71JW7IP5dJLQval9a40JonK8qvbJxe/19L93zpBmb6XaCHgZhLjEL+PL4SRL8+ZdegIUlMtn8l5
ZY6nC3+/iMkFS7Nal3wdWgxstGpNm7KgoDiuN5KzRTrgjv1wIX1jBnl0Apc1mAfx21vib/AEo1M9
F2ahnJ8/6W3c360ysO/zPwoRM7PN1HmmtNTagXP2k2nbQ3+J4PziwmoVJeYaS2l/72ujsjRIDOGT
9CWRaMRuCBF1L78fXsQw6U5XC4KRhxeu0ZfjjpNzWyewph4A6WSAKuPc+piKbrQ7KYak/OxMO9Hq
OcSwtk9kbY154UfOHzKfx/KnJEbGUHyOORRv4J5wfKNPnf0IpgjRuVpOiGu8e6YAX4or6+PZCYUN
Yn821oTph4wuq/9Qu8sMU4on+QnefMb1y0ng8uVauuAvrzco1c6druzgYVvGoLuIkSoSzBjsmTsO
fBxnF2BaLh8y3CVX7VI5DoVpycCoB4kw8EyTNIG9/m8VD01dmGAOjEbFTp8h7jGnCZQB1bNL2usw
E4Fg2nb+oR0KJFrvELGuqP2jWeKLFaPdRmze6n6jq6PRhwEdJhuQC61Ls8h5MYvIc5gqmI0FB9oC
PP/g1NRAJib1mZMM/+LYGErnOCGn981SirlDQjlCr8XaWv0+5btFmLZrDyqqehNdyYWXWBg4XkhV
WRkOdQrZFugU7aRY5m0hbn5tAQl8r7cS4YDF5lKK4Pg7ZDzdjncqW0DoV9AVCbo9nP3E2w8HzZMc
q0UTZmMCXc0yNVf/FmRRysaevUGpXp9FUS+dsSHalK75SYM1NsB69cjBTiXGyHDjWcy+Mo0lYgCQ
Ogifvg8fGgDkoKZy6LRnGpbAnIzfBp/QJ4MigqRKyWp5mUnx3orcyt9W+Y5iHf3tQ13e8dpf4CDY
qLZfYvEfeig9WvkI16/AkJABRTf8f2aqE6I+qZj+GQOsbKIGz0OVSPgE04OZJzeWL3Q5kcwaxuWW
RDt6bhYvXJ2aX9YLRl/7l7tch6KUPC9hijpgMLH8WTOHP1hvh4yLzauHpUcswFqZp/JxNBvEktVK
pUZbc39aQIs+8NtcT/rhhZtabS1xECrqgG/9aD9JFn/l3YczEeKMb4S0m71LBKnSHOXcyynnOdre
VmIHWuz55YcjlqibAq3dSoiyxRlpUnjX1w+KPyChRUUBm/KScBy6ppbYU9fN12OslpAEPPMURyDv
j5eqOz3bEMowBTn1Rq3FURoN5VBa74g0azR1H6IBunimFODYkhomsS+TMou4Ad7R3+1QhjdLRZ/6
B1bhD88jQhvbPVLYQGvqAyaNZaW8R6vzY3wsydnL2Lj2PLCAMd9sw8+1n/LsDPvBf55ABAPXhyCp
xxUtKiuc2wgqMTTNzeGm1Tb4lzb5vHcCYXPNP1SlSOwnVyydfuoVxXCyEGh+kYQr7KCBrpxqsu/G
S2ISUd+7pvMzZAGQpvxmZxXLisJUfVGOhvxK6eRlu4kbn0MQJopX/GkzY0gqw6oH9uue0bK/bTaC
WzcU6AKm3h98rZsFI0DH+fNCTX1Gmap1jv/1BOrnbvswfd2hqm/sJytvhGDcvgBSMBz0TU/trOe/
jfsAp36+4FoK7XQrQwgGeLyLLOXLrZiZ5XibSkndkuj1YVEGxOb9IScXgv/gs1m4Wm3cCJlDayfk
rNUsuNvwOtQP48n1Ysrfj8k/ELGgFtAj5CRwxipBeRfwu0oIgo+kEO2tbqkPvWlEiJYi2kfOi2xB
z4kyG1tvDT3AafYDQA9fzrsegaQh0FbSJGuFdcRfrhbKM2k2pClEzyWb0UjNaI1oKP7F0CGQOz26
wtW5TZcxhVh2vsureJkSA0WxhW2eh3HjovxC4Ot7pYYKRtWE3hJk82RiwROhWZAWoNWPhiv/zfkP
6/UZ0CMuL6Iv32oWiAFjeKUFSarNk12YJTzluC22oEKCnt3ksGRTyuhFimRfsh30G12LWA+lHdEC
aR0PsjhWTjANSUpCJjzaaj6DL9qxIUspje1QXd7Rdui8OF+3Oi/8KCrda8wrsZMh9uwJpNVPGmk4
jNGVS4z9UrRwr3A7uDQgfoloQede2o29MDYUWfXX+uFYdczKaof3syC+Uga6C7iUnOxjqJqP19tW
X43pNkhS6Iifww5kwymMTMRSPWWL1zWXb81Qto+0hENRHP0XOHPYQXO6qZGjNUJ0vUFdbXSlTLTS
hPjVLfaIyjDdsNHskhtkcicT603/65CA3VxSSr5796QsCkjJVRFS3RGeeSXP/JMplg7Pr8Ltv8LV
dAa7a6Kvt0JoBaZSISKG7A3A4xfa5EPfxv6LbHz20evsIOegCJOqt+QnWCvSHMxn895fuaC13CCY
e2c3YjgCGD/ypM0rlKElI0gHy1IZ2FwrlUUAyo8E2seuUGKcYX+Renkz/IzZGd0Y2gUrdogmbn9S
0eom3QoL7tOh4in6JptfwFb2LJ9gxi9fPNseexLAk0aTBwPruLtb2dnKd69fbUPcK1kW0ie7H8cu
33AYmYaIua2do482pBvba5BR85JUtRRgHIIwExYbC7c4G0+hnhF8g7wXG1IL77qBX42XWkMOzucn
RqLKDOzaf7DlvAW7vJmAg3IhSAhS98Wt/qitqGsGY/FtxOVYo3moSIiAJ2cMFeKGzcwoW+Qhg6M4
ZqWr1uYR52VUPmxow8NzPfqtbamcwAaBPSxqXnEzWFNt70HfWh370zwgMTg3CB5SyYxTJ1ptcW8m
RZlEdZL7F1b0zlXX3OtXe+zVHfV1crmn7jZK997J/5krQh7JexypJd9Vk/U++G2TFvP+Cy2fd33t
FaLyXNzhSyd2lR+ihhKtQcIYh82mc4HHHYwWVJhYeCGEbMEE841xdVqDRyUcJvz3lsZbyG3/zaa4
EKM/YPCPqVUVkrW17eQfN3tGj9w23AkzjOswk/BawJTdj29D8Fn01x5fnyh8b0MKHfUoNFMFzn7t
0WSPeQwBbUEUr25taUGqtTA/mLAzixM35PlTtjXKcdiNd7RHEHS13bKFSFjWGD/bCmi7DPAqqCtA
rrypnLicTwTZsF/K5PMq0Sn7XCkgKIUhPlQkN3SYnKDAcVEPKSJWMmNEEqx+jzKa7mlPf/nMgHI4
Cdmyiv6h9GLaNwlGq7yJaqnL78VCYJ8JAIUlx6Mt48jhWWndfhTqnpF4tXDbcIUQg+BtI08PKebl
zEl35ENAgCBbwENFG5U7Iyx1j+d2Jc9FfUTpL4HeLwKx1tPIdUPRDSf2MmFAwkwhuuIisMozc6oZ
KSszJRlJu6PujdWqMJa0YjmmzXDdnQK9kiBN6GuHSCLBhH5kx9gJbg7iFFqvUpTXt4aysXajF/uu
Sbz8L1watJmE9Q+Uw3xoEzWbQjhft4Bx1KwTvYCXMbGtV23ZKOHbP2VPtlAQoEnF4nctdettnuVv
l6SKKmQSFgiPvw7hB1uYupcjCX5SlkjKhvVL4ysv7bZGV7RRe9VQtwnBOyt9XI7E6aitl+yhAuXM
xnWMSlYcwo10IHkErvfeb/qmZQt26OY1yRogDvA695jXLp1XbJlTAc+xOMK4U2xrYR2/7Iq8LOlk
6nHk0IJn37KNNNjY5e68jEhQKzfpa135rZKRhpZRwK1k4/yqRcQoE3WEyT0i9bEprBnraDou4xb7
0eCXUFu1/RnHBEmLq6ZS/lw3qt7QBGrxVuGgFKos/BWeLg0cVCFND4sst3KaTNpK+eVaiW4EPlOo
PB4RhtcFZpPA4CVK4K2OD+8p8TCkMoHCadRXYAywbcaeEvzv23Of7NMS9latrvOykQs541OIIhXL
Z+x8YH4V3dUfmNRSLVB4zRokivCQL79PoHNnWQCEf6jYPnff/tNrAd7VmQRmsog/XULfDNtxEcze
HI7SPmtR+i9G3CjjRzIk0urcOB4Sc+enHg9L8E/7ETUNSKLWH7aKY2XQLNiUPkMLnadqOFlyadwM
4lfHl8lah0wG54aPpjupkfUbjoGVBJ4uOnYtGrdIoCek8KINxqjFZvnsyh263eY4AV/s2m4DmzLO
ZzHDAP8y4oyaK+ljfjmgxLJOuMrLbIx6BUVRTAD3SWoZKMNJX1YhFF3GU9DYm/68LH6c6/muVuV1
MwYMXw/6dSH9q9xamP6IY36Nh2y0evyo1Mw6IXvbMvLT6mjLxKL8+jJg/lPYsGctbvVNWf/TtBav
eX3Ltt7rbRoLiZ7eobiNlT+2ASs3M0dwxahbIneAv3EW5XpuP4QJ/1bnMxcznc4hPJ6tE0GjGIEY
8wobwMlSKGP9Wk2+yqQJScOT3UzjV19R1xPSWTnZ/bSYcqmILE6Ea7LDR++tHmqf4Flh+sDOE2hk
Dhxfvy3GZT8uGmI0aTZk2hAfLTt3pUV6aSFfrYl9nIFJFU74RfTXUADOgcdJldzRk6wDzPY+Lz4T
3NT3kHXph1aUvvyW5wZTC+hPod9mftwUDWOwnB0NMaqBhI9jf2ywbY42Hfegx/rEV8wZ6ibIqCOp
B6kd0Jy5b3o/ZFnw8ToLkkhvNJWZLmQhls83BKefQx/VGQtdzwPR4m8eVIVboWNQg9LrjdXbeYVw
YzWIZP+YvJX2l3JSUEULHZGaPE6zY8NVNtav/97lD7Xf3PCZhBBMJhiwk2Ii+77D+vsY+7Drx5RZ
gGNfDzEgJRtDuQpxVbXbXASBLdCZDZefArlFDfKhN2XEZghtrbaKSTtBIE/1jP+AoEfaCfflyE9x
W2exI9WzICF+5kl9RJ25M6WhCO+X8cTsE/FJljekCLei/mFDpldAHkz1KdmIxoGBMMaeoKjOIQez
EeoLPgkj/Ae33Z5hDfOVfv4lXc0BDejFTAGkhPP/vwFykaffmYstjDKuUy/5/eZ9prlEIYfiI9y9
8CQ9SSj4RtML8n33NcFDuQDw78ReYHKmlNOKxpqEoiqF0BAEBJDHcz2rlGkc0JJntDJnz7aczNg3
mTqW0g2XH8bp3bYfUtRvu3Mdy92vWtKcxjkkQObY2dX8MKfE7fP3XywSyQSTOjXegzJqCP33ebZu
NjMa/4q9olcbD7lECTfQLFieqNpYv42VFWp4TNXhNhc6Yo+WXocHLw+BU03nBgIrGDHjGHZknN60
5DQyk1bDc2koDFj7xUBSUC36/7ko5bJikp85SpnTvVsE3eKtZk0fEHGBS6CELqB3mf781KR8QldD
bnqsc6lY7I6dy0iLquYO7L/VNve4HleGUWvRvJKxxKxL/mWB7okVQxlrTmPUt0NPt0i3VK+nsgu8
hJVNPP4jJIi9ATcHSI51zltcn4HJNLeikJWgMbwy2KJidFmmpomQwCfnUAZHddgap7IEEiHQ7Xvu
i0x8MxMfQ5PiVcsX5eO2mT/PbtDIEz4OhFVNL1nClNdMrCn8Uafoovxvt/XH0TDcDIa2cqGaBVtt
sQSglwA9j3bwGWpxdIQaYvrqhHtApHbkg2rjYNLTpVm/eNOTy3EOF6O/qbhjYqJFVRnuxGai4nmF
aLgwWCikgM4rgdDlrO/1rDziDwEBlWs819J+SZsX8OXgAcdyMvb5NcBu8E1dC4EIX4DAro7rP2fX
6zxr6znpwS6azT2Pl5zydcqg3p6gAhmiXmWIzDHLFAWLKR51okpAkQuIWbwmXYsYzrEBvf8rJ2aR
CJaG+XQfc5cBr0+XXVdFuSgeMKNuf6jWkpwnWRNiQOlzVrJXoUMZduH5y0rj6pLoEB2BmKj5YS9I
vLjNxx82xTcmG08WbLBrJPOL5eb5B6ihYnXDAfcimSiEuLgrqwk+TOu134FWMxV2IgY3RA5QPJuz
A0AFf3phPmPTdzAkju+vbnrc64n1l6PpHL/5tgh++tYhLrCPUZUakqzEhDn2KAZg6jufvpHKtaJp
wcARaPCbsL8BhGpBKUlTWfxaB9Av6AW5jJjOjDk06qgiOLAUyxY5lg7B7R0YliH62saFjFwKP2CH
B9PMtGTQRqg5JQb1W7SiPcr6dwn5O+U/JQCzGTqEmDGBQmrW6yOCjP7JtEhSbL5lBapfl/IIOWF+
Tv6fvc8unh5i6meh3ks3d3yGF2UEHCdGegMmYvfwn29thHpA7gi6rJ6LC5nlkWJRMVxFepuhmS+l
FSenARPCEnE4IsV24sWyNv1dLRMFPQYZ2NWQlDjisknj3mDmpyZaOfDd7wYpTMRWGylmeeZneUov
h09v3XSDnRKlcJ+eNNCg66dJjsMmULpEamDWMzLeTHnER2w+WvCbpiPIxxJVPoOfEaLj17UJExUU
w8wXOxhyMfVPOSmuqRV9CpHXNIOYcEfNBMJmmF/KLbISjSHmxj8TBTC97+kqPY03+cv9ERGZSuJV
l/q9mruAElZMg6FveKcGD46u5HET2FpXeGJjlqpWnkL5UR4PhHhUQqihbPIVP7ascxWAVwgbnPXL
PZnXwJ8Ih6ewm2gJ025OLTHBeDIeIomiuGPNfk1jt2NlhJAyoN01N/UPxNJDkqKtZF67atIrejid
PfOxeDgAnXH891YXR1jROgyR8QHCbTeczMscci1CcWpp6UsyAl64CgtElP86pVzMPoZ7u8F2cfJw
WHpjj6ocYCZ2IFXWduxI2WlNtcFxld3bKDLSunUK0hWlnBkk2r7aGAXUnfFaT7oE3cx6+VwMubCq
qvNNKdc9Mpwq+CI3lsOplIjNQkl0CXjpj/m9jAzOs/EPEfC4WT2+JqRC3cYXGDrgwctdPPDRE2Lr
3aagSHjGcfouo0WWdUMb4jCzFdooR4v0lw75zwidbALWt1DNbjv9pozrwWt3LoLRNVnGrrbT6gd3
FgCHXEY/i+l2DxeKLgiWHxFVWiuAd8LbSlCmocBhkXEbltUCrZnXkrBhqTSbPw80wnbNGdEn1uBp
P041qPBNQTodwh/jn7NQDtsDxzgwnbrdAv1ee6L3fbNjIqVUVS6fGN2cvI4ylTWg20I07xxCgWKW
8tDv26N+eI2wx8wxlU0HtQwz0bjY7oPh0Oj/uHo06H8HLZffP4fWPEBby7NgZNlh4Ysib9DOnRHb
mFOf9ig3Wvqjaw0pp36nMEM/6OkR6iLmQp9wKPdyJaiSpwB8isKvdRNsSdSBqCApZhMXIfWqHMRf
DcFwx1VatxTd4KtWchjZq7gNHnMrA85ADVcOCbDWXO3LEAtYgEAv8HsaxJVLSh0028FcYM3bOe2Y
skSJcutr1RN7jsELCPxLSo/Xg7cTvf9F7LDSeTtwLCII59aBM4a7cS8EYtXQMWLOr+MxrANamRRU
4X1BF9bPyRS+PF7l0RiLDzEvsK+sfgg1MRKHsddDEte2jCpL0DnTrZz97GKHpYJkx+8EelJTZo6/
KiM1OUqLukstELgyDlWljs/XIyhhkDqIlfth0jLiN+sxhs1AtKRzXjQn61dSWR7G6r0UftB7N5DN
GV6nvXOu3qlx5reaqePbYC7ImXOELn4OkHEYYqUIw+2MopBTgL2eNrgid3Hu+J5GwLOj/jrujuue
1yCCuBZdHwVl0hs6MJ0ot/JTSN6Q3pnUs8Zhff8sZHu4CJmDqOUn8bt5YjLjyxVV3aomxpBUkvbs
hf3eOFkKudsCq3dRxUutEkMjIWp973CYmh3v5SqbSeHyc2FSDUo07apHWIxXDz40WHH0BlzJI8NS
at7RcjYgEq+tPmGvme+HHVMo2hCGMfYl/FTPIgFJQpRcKiFD/kol7Uhb3q5hn/+bQE8ihwtEyPXY
+0V9gm59KR8ygKdizqTK4dtzkzV4EfUdYRrYLVH4WldLXfU0p/kJ6sirpuOBghFyjWltW8rJHp5g
nvlJQ+8T+t9mSabZ34824w3DVfrtVJau9wSdgFjPek5O/xtciaG+6tfvXKKyIfJEPxiPBoX2l2GZ
mvOIgm80Fm5S+/Ey+P2iVdozcjkVWuquKdJlI6o8XEpRmgyLuU3bPyeOZOs/XErq/AZAtdzIhX0v
CcvNbXeQ1OPWKDzAPnCAyDQjHMc/A7EK2BnL9dEoat08CTIWHMJMoSdIE+4udbqWuPuRxPCn2jyR
V9A0ZC7wjy5Gq/wSHesbBn82u2mDu8u8ee9BcqIk3jyatekB8guLzb41MjfylzEHnWTYAamRN9d0
CFJ8e3tNK0m+mMl3SLyac1SmWc7RIIsLVM1wWo0f5Jjgh1O4X8qWvlcobruDgidJF9toRT87/u5U
I9YRH5b7t64lA6aiEXC4N7Wi62ONoYuTgGkM0RuePBnJCZ56PDhx5f3nI6FoMBuvpoJqf97PPZyy
gbkzfJCtXzz5FwboVmZ8RdlmX9dbAPHVhKMN9XwbASVjkyXg1V9aPoZ9MlwqVSH1c+8OHfHFoy+P
mgbYZqWdsAz+nMA+sFZShcYUing0HJJ6hqHSPQXazj1B24b+re4EfNf+7OYLwXbFYa1gykKpQV7/
HLGiRb1WAefISVZi2o/tJfMSF+VNh1b8htFhX2eZb3aW1o2pAXa3kDsDvnQRh7QUuEcYY9L0TI2N
OzDIqPSAYKiwSIQrS6TpSrB1LzjeX74DRsrn8Acwjbxou2M6O0jqvVqyvYNN6eOd2sAk3dtSBBzY
M5CbtlBFuRtcoEakcNUV/Yux0Xw5Ihz9oux7Ctv/MWghMpCTmIzjOkIGsrBeGcidfWh4ePeR8sZR
MFFAqUgQi0pVum3ER5ApDIrb87GTgtPMpjtWvcKgA9mrE5tyKisRwT0YwqeIpzRaw4Xbv/MHpMWJ
KMT/MsT05OdMnovEvSRDsMgbNWokVeTwVdak/QGBvihRefnAclxbenMF02A1/iilH0GDgPwP1jsJ
PBeTOzY9JDYD4c1gTFUUrtPvi0FOaHSZBqj4LLWjnHBEl1fkcnPDU92qivvPSLv/dPBijSMOTbEf
jjh/OjQ9s93LffO8WbbD43ZELLpTYvcKmdc+SlXgLQ3pXJWJZ+Qf6VCmvBk/s1rP58EPlF1Ol7eU
RD715QMu86FFjPSRDQFRjZw0we2IstShj9RvhjBqHJ00Y1pEcYE1QYj/r+qpghWn3B+zH79mKuvL
qh1Xr7PRttYtW4OrmHkVSmihpKo6pE0syMWeiAAr2khf1nG2x9TR8eYe5+mdRunIPl+qZ6s1FqM3
/CvR5mUvIjXy1kzl24FdBo/N/cy9G6Bo/JayFeoV4yylaxKeq4S1oTcBYbhl+UVtkY+rngV3pwaK
5HYtXazyg1qA6soyIjhcaT+sBLJmAod8LbuwOG6fCfsCsdw9qfW2XM7tu4ehwr9YKonWOXH0RO1h
zTdXUgyszh6ihe8Uk72YE32BPP2w2nV7fUWz+xnOYdDK4Vc3L8JHlNtRAXhw9TNCE//h8hKAXhxW
s7v51BSXAQXU1mug1ReY/czGjh9CnnvqPpmcGBY2WPa/Nah9an+3lkzcpoTIcgExmMiryAYrUtWR
lmvxlZKcf5D/Xl+rrGdc+rsHeuCGEsokPDbs0txS8Ef8OqsngLKzTDr0g8mkKCi1NTBNrpDjhe4F
wsLifjfcM8AiM2vjZY67No6TDmJIevbf0c0VXZHq38YJRwPnVMvQ2YavbxNnELu9Jmwq+B+ksuqb
9vH6Fay7X6JjEbIT8ERfTfwe6+/buAtuSSy6JISLnU+8oYlnGYVF8b2TPs2FT1hpCYH9i1Ca643U
isM4kGbD6e0hkEA5rGW0j48eTC/J6z81+RFBRrXbt2gwFfDgA6brMhmBatvbFhRv49TFcKAk9i1R
0Kv+Aa8hz9ZQ1MUNfAeyiBBmvPdVph6RjCdih9cXZVO+l9+o/5OFG4abHg4KTdHwqHbyU+ox/0us
4UdZkEjMM/fVWzh06pHgN98YXcZHYn9FBRnSstd078k4gxvzKyVn0SUXtjJvqA5SsWpcqK4rL0ce
TKZ3qqtjucFc8HgJGK+MjzueZfpQBOa0nJiel1lF/nAPDho9TDfspy83Zeeg+PZUoSoFjSUspQC5
zMzyEsbf95vEnYNLEDVNnfHn4WMCIlwl5dLv0kmbhjf5zMA+h/5wlbYA5A+s9uG8MxGV+Ziy7WHB
GtDPw324y+ZT6ZlzbEPk3QPH4J6ikf/2Yo385Jg8XqSxyUvfmJuQNrnHfIZWIXrnpbACBTtT5g3E
TJv7AieIJsEoNCIs/jh4M1k4J9gZsjmfHGximFiqc8qOU0FZ+jsvpqmqND2eORGsOti1vDl7gPEY
0gbPz3gTIFyn3p5w27kFmEtT3r6lw7+v9QmvQgg48OmmiyK46XFf+AgEaiwhNOI9JdfGH9yv1jM5
eENa6O3t798tlXIpn2Kuo0KzpZCF++ab68xAuawts9cFVJcWxjwpWEIgVa5k0Q+E/SmdjcTqLJ2J
fBUo9U3sfkwfdP3EqRQGMZlbn0aSI+oRnODBLqNfesYztKH6+JD+1YB1rnKzW5+CVKNzbPvxKAob
ZnQ4H2aKsYRw/ocrj33J01ivEIFiFVadkCjjUy8YgCAgJpMFgrlBiY15nTWFlg/XFFmFKFhA7PnS
Sc6twXUQ0atzaFS9lshqQSw1Oi5zbn8IY6wOgxMRCpIvkkP/94hHAVOnLIwi29KHBxdzJIAg/1Il
QU+NMegWbjShdvoOsu/QRgpk0JD+99oKUT3+aaEE3OkLimj4UwcZFnrFGfqUOQFuFQEn8N6tn+TC
9WSheaukjScSCwRjer/+ENtq02t3waMPHMkEWFGwuHrlpDhAyg+cnsyO6ycPWdZVfzeF1nFZVVOq
uey13CFXSwajPC0qfaGvZQ1JR0eJNnXTL//4P9BWaafv/FZCc5Fl/yui9X66A73+PE0G7jQ73Jar
5VWwW+8Vsc5X1xxnH4bZvSFi9sCD8E75+9UA7/acpRJeG96AvKBfchg9RM/gckZdMyvwf83eFoB4
wXr2xVTzbOPx8o5/Xn+SzXKE1Zr5HFv5aUKyTBmjCJPhD6UENyylicaO44eXvzZsgR2EBXdx6Qnm
OOORocuxoFgFZOCOal2dCEJqEIvws1TWwt6BoULD4NrgwkpKy4j5hTe+lTpvxyBTWP9I7whJKaUR
k/fEQ1Dbq6RriXRhmIGUahQeC3vdWobnE37SejxR15ZJDiWrSYpz4TMFxXQ+yT12xaLk7VAv0q3p
nTuE4b54MdWhsU6nCFocKCW8gChp0QXwHvvOiITbAe81MYP4MN5zw9CcTBEk0N9M2y1ILUdr/YHz
Eg+awLDR1VE8eI+h3fk0YUFyOPY7UPKtutWg2dpYaLRH2PUBNC4rpgOTSiXhNFCtlaWHGZBbBX8h
fFH1QxWuS+hKwFshtslheFn+7xt2sEgGucdE3iG297lq4KBjKhhjgLwPHVnnoyZvddyAHOGStoD3
1FCs/3fklatOP0gUZumJSgbaTamRYr87ZS3YdLa1328TVbe3IbLy+YNq+jYOhx3kSnqmTmwJtmXe
MyvVGAKlGQaJsjzTz2SV9X5QDilG59+HhY9O59xelKmYyw5G3Hb8IUyJp7v3dN/mRE+DTMWziFYf
XhbLCfOOPB/hyCHeLvWRcpfciJHQSh2jAMTdZo7EcTOXUI3jNQ6jA1TT3ZaD64OUhe8gKJ45XmPg
xkyqQAZkpgh+hJ0omNVLquUDdMxccVdQLVW6FI4nsNbInB1sWNOyIJzhklEQ3UDQI/BL4DQqO3Wo
8iSR4/rl6JS85crg7qPod+QEs1T+8LKlVTirGGsFmswb3WqrK2d4MSsaFbDG0m7n29XP4g5VlpRT
GfjvjR/TSEH3e2NertnidzvJfXqEwss3o4/t6Xm+Ic8b4mYWe/wJx0fFGDjmgcGYwhp33KrP+j5X
yUlAuQcpXc8m3gdkBUfS/3DQLbs7byREO4akHVUKXeI1uDHMThuJbdvTyuCL/Ru/Y97PmlzsGxIK
RX2i/Kf4zP2pGE+FtTDvdOfUpgaxKRVFzKHfPPrqW9ZApeV+qUjIYunCuDttB664Bw7E/pj1S5xg
DHuMcM4HfmAXreMfAnn4yaKm1bEfhF/MMi0QES/hmVNUJhBahPv02/qFwFvMOMyEO/CXkO9pGGyA
kpcEnwdhezG+vv7lRuLI5x809Tosz5bXwG3VUq/PNuSykAxwGVKl/Ry9qJ9sfhRuZZUcfXQVK8H1
tjhXij9TuvMQMR7FM5udyTFWy80mzEd6Y73Quddc30tDl8vnkPPbuW6FjdSZ7mFWLfODK950z2ll
w1t+2hm0dqXGkJEuIcRr4zY6nalfYWbmIoa6FEyIiEON3kwapZurkhjNY6KgOWGswde9igxjiMra
cSynsZ3jno4gcHCeuIuzZMRNxW1YGJSYc9GdZhLUzZZr1ZZMjqGyxMoUiGqhXori9d1+cUt11ZNS
JNrl/QYqIgeX7vwcO/gdNSJWEzhmYs82dxWKP5T7AaxMbdGRn6n/iquTL2ge5KLx6CHWDFmrRUSd
bGDOFIErjtWnf45oVeEPeh6KHQGGxts7LFpEM7yhtRCz19Ws3swDxcj2Tuzy9CC5KA7b+X9A6B1Z
H337SdL4A0wZy+MAdwif16FHOYHkzNfMfifCx2jH8cQktl2pTu6Z32lpfpP6h27vBwhZBiIjxYZ+
5QOngDe+L8iv+/IoEK9wlkDZ8cGTvTtYMF6NbM44Wt+0a6d59gQkLIFNCMUiJY0Qsz5c3MplFhbj
XwsPk5DoOVuNz1dfTt54gSfif2xEUO9D18SQ+pR6uDT9OKdQnDuyRkQmPAUwEFXwlaktqncBLbXX
ZFPr2RR9gY9uUTlwYkX8gp38kjvej5P76hmIofef1yH+rYR0CiEUb5ExGg3vWj5Tw2lh+kcKE1Gr
0dkpxUNkx3oZyQPwDnS8u+0THTq6VitrwCOqUaInkGVCmiSIBordMTYiuVm+0YzBeS7JBfTl6W+j
TNZodfV+Ayn8ULDK5JXCVwjoTxbFdEggipJbgxT/LQrwpBIiI7wGcvSaea48EaoMzePFVJ5t/hT5
EHTf93ArYkcB9TdQ/qyuWzLtLO4U7QljFMQbCU6w/+rg++MXO+lCXEDB12UrFLAjVuvldwYFbmvI
QvR3aw0xvln6l+iTOuvcE7EUMHpDmruJABC7ht1EXlXK4lXWKd74Ccs8n6qnqjB3Pv5lBGWNNKb7
9e8ct5pQs8jRRHeuDx6RAjO6OYElWNgmiC0+o7u8zW7NEs4InGDE0T0OGIEPPrWGMlISeMq43D84
sqzTdw4hmGAb7zbJ1PJhuldXwnVoM4LM3n9M25qeTpJ67klgyGIRVULA10uPSXlOuvK7g1kO8sNL
EQlB6OkOvfqnTnbukFyLnEd20IiD9bQGFoqwWwk1HldX+5z2Xx/rEQYjVnD1sOvxF1EWSlTVrlsL
QyHaN0sAXwoYf3qP1nmu/OUDOpBhPDUZxGV9nyQ5UXKke20vAH8SwmaoG33+ryHECxedsnytJrgu
Q0zXfDETVy4tDOlYRoVdhhKS5IjNryfS15s9rH3P25b1pAzhq4QbRmIgqPzm6IetneDaIEGosCsU
tL0voUfE8m6G/bZVqwuhVVTM2y2goTrmYNeeCQB3NqlhdOLXEO8/9mLw1JeuGAuYSuaPRjEjU2ep
Tl/Zio/1/6o2oaN/JSRBAs8BmxsSSxyPlp4gQnjnHzXiyqH51dr7aMysumXrH4kXKJX+CQRh0sst
O8bZOyn7CeLl5lPaaJEwDfpgDUE/d4mkHIT0sWdZiE4P4hwmoYUd5ZRyY9MGV22umh1SYnuvlAGn
h+wTC62x8OgR3nxQYs84CrH2fHPw7OhYCns+Z3hMSrnrlkVMcoJyBcc7vaXHL6yGmnSXM5ok1LUC
pxxHXw3h++24zSHHImdwUIl+O0mUm8d9mFgJyMWO+Srh1Kn/ge+tCR7Lruw27NaolafIvjKDXs4Y
8/dVmEAUyHkuHAr4mJkbULDlkIHdJbxfkY43UDJUokG07MUXmgrMBIlUyUpFKeRVbCQ6GWEWv6uG
y9gc4WFLBtsryP14YbVUPB2/DvNr0EYLRurvJMtIYpUin1APnqyrjIStlsJzVoshNfpceqXB6j5t
Gg6mpGrTxcRZNGwVszLBwNnS27cznJ9/uDD/cxr2tKvMFKswsiUZKiNvRPzv80oW/FmIb8FKcNqd
/gmPC6HmFkaBh5+1jXGa5EuoXmrKu9fak5PkbQqNUdweIaGqvaP+6yFYV9f8byV9GSK7vd5UC242
tEwBmCajpfNm95wq2FXUtjZecdE4cCl4qGTE5Njt+pAi30noOY6WcJrXn5Wd3s5RVexp5G9e+Uqs
S/IQs+1hYB7xJR3mYQ+tHX2YFFoshlPNIZkhHy86aN8wwsQhO3sPZ3oFMuG8FYbKk1SAWVlnWEvv
kJmbHA+LwBKTayiCJjx/jWPU66mNOM/nvFXKtL3+7q10owB1KvfAuPj0O+JizSwKlCATH/zVfirW
dBzGMXqhw4CFlCt7VfkL2ZTHIL9r44GadP1paxcm8CQ9wVhhk04QFnG6eA42/gB7clyKzLdHslVZ
38mLKFC1VsYZzIBSkRNGlxF3p2o9F/BgSyXipZn350AIrpCxuuX5dVEeqRbMGV2/I3GmLT/xp3Ia
jWHnqlqFAsFRLGdbqkWSxjGKJOjgL7slHyAzGXJihyutLYWPY8e0wcZMw2/QNCNwb+Sn7MVd7wUg
cTJvofP42GfrbykJ5rFbr/JJMVDfyKurOH1GofN01FqIBtsK1M1AOBPsVxwD3BT8F+HSloBE6xIF
U8aF7NH/7hAsiMMJ+D6oIIw+9zn1Hr5T4xmzM0o07evHw9BF0Fh2td5Wf0Oo7O2VVKoo0ghYkGly
fNrVfmQKHBmzu1xUD+gC/C/wnV8cgyV2tIvYY1c69zrifIa07dUtsKGoCNh1mzsPhYszD7yYd3QM
lZm/Uvk3cYSaVoPYA5YGoJuL2bMFsyEZ2mfyRlfR+nU5esy38ka61Mkm/pOnTlCSGZwt7sg6mHxs
fOE8xCaS8mEDNxWG23VSICmomkskjWe03DlOid+ytS+Xdn/lPnWIqrpZp4ZGnoL6SChULkaj5mqS
8Y7vEJttI1TohRYew4VHzSlYry2mf5nwictrcvMJ6/TAVuMo3x18M8B4IRA4Qre7K01DtT04m95k
5D/mqbBC2sQrikool9PKmgB74Kxslhcxxy84hyPbDKYvmX800Lyeg5F55h4ldzp9Sq94ttZqfPDt
uXwtjrV16kYlaQ9im7XIfB6ryBMrzQuT0Ojgwjhc1OzldLW8qZh1plKmPdDjWUkMdi7SxwHOWwod
pyQKA5PoUKL4h+qeXAqmGsMspioQDPxuCfXef8uW8zOwYFkYoDmnI0K5I4HmIg84eBAQ/Qu7Axw7
EqR0+6SixLUfyQD1OpUSar+ZkEiAAeDYy4uASqG6ronJSVPlOxmmbX8hUgH+aygLpdNRspnDa4iO
7Ppxc7CqfzIcU0JIGxbpE+yOVzdpsFZVHt4GRvM7i3SsnFZIf7UiLoW9hP6PcfGvd7sABpOyj+fv
F6VH+bDf2+o6nMEfD1fmnXhnzQOzxvoWVHUB/xVVAKbPl1RU/M1tEpM5yuo++on2IDMt+3d9NKZQ
PZ/yZv/8jKseDKUzabml+1P/fjKP/qu2PmVE/MpesqwWACtUlo9DGjG/xHNlRvuMiFnyfuiny4Lu
xE9cXXSHDDSCCAH8SY+mlYjxLaDetE7blIHrIwNw4PHAax+eOiZXP/Q54ccvtGoS8TvVHHj16VX2
XFr9vuPiyovIRXiuLbqHgDfl0zKTTZj1yFWxzUMq5o0L/u2KmEBcmHm54LBjWqr4DvPWySeEYV9U
e1j1s9ku4pb7e9hXpcZD4UQWhxpPuvABKpCKZPfy0g+KnkUTpdTBFtEZExhsHJhM9kX9hQjGn6Xe
cyJuR5U5SGLFElpLX+lh8HwsGnZfK11WCrxrihOW9MCOpfOk0G/w7hbFYKGXA/C2XFIvU0N1Eysj
fKsjeFibyj1mrhsCaUFSNbPCnAM+JfpsW5gIpjmOjkq33fdsTByxexIgbIXcLBPPqxeG8fdBLz2f
pV9e8dVZ7RlQnJhTyhgtlmO41dAGs4EPXmbNXoUFzOdENhu+fzolOrjSFOAQdmLE4cCBwC+8qD/7
vDaarcfCedMSuZ3RYcMtY3+SvS38R4MWpMCkxGESTjN7MbkmiQkE85zcoETvfTZfd7r6WVoUHC43
FtjQf46W+37D7T6QWwI1NTUD+mSxPHIk/pffjPuDGBOqKDrBbcpk+NpczGBnqpxXiYXXOrROyZIm
uDTRDGcKYX9KvzIXRmJ0eaJGHTa5NMzG0M0+kHyvar03hZFtw6DHNdigVjJ3QN0Jh+FPAUIhvM7A
kUwah0Zl8Ni639GjpodpshV2637PeYYRMSTibQE9fsY8F2vnOzrWc3cEvy4+MNL/DUmrH+qlqaSh
XwckY4nrEHftH9UJyPybKu9t2nTsXOihBQaYvs+2CBxI5Rb/fa0BP/0duiTtCM4n/r6hZLmGx/WE
6F1lA9Tl0Es1FcqlN9DetNoa/9OHuksBTy6SrZfLnV1QjSHqpe6pQjmg3mgtIzZYMFdYrR3A6Ko2
w7POJeYVouNW5UZ0gGKxmnsTvrqruW6/yeaLvTMCxY6puIPDc2ZQyMNNGOHQyrqN1dW+BQNi//hN
6sUOPlmJQe2YMOhYFffQD9DVrmISn3x73y5jmZEWuHx4N2PnJWvpHt7xrjUVLe7qPGbGQ6E0U2eT
atiXfbZnZGQWAsKzTUIqk8z2TjiaZ1zExXlWuxR4YW7Bq+aU2tUYg/I4MlNwluH1W6R+O1dVZT7L
sLT6kGJECXNbDzSm4uPnRrt/46cFdQiFaQo/EABybZY7CcI3auKKVs3tuf3tJ2YQyivaKGq3njBf
UdS0uKyMKfCQGtdBji/eT2jwRqFOpBCxS73A2iuqrzuBzh1Jgcs/V2l7e+x1TTzH0oCsecf2JyTe
KO0yXdDIg0WghxGTJSeYNSgpiFOHVWlbRI/tjVvuioD8xbpKDhrXdm+j1WS1tSscMnfTM08AfkfQ
/29ZrT2JydTkIWfRM7/uT5CVa3mhtuZtzxep+SmgMJOKma2B6UHzg5PcvElmSjLczIIzDWYkk0kz
1vs03rLcbmeLybjViJrbYpj1ZUOYFl8K2+8FhW6+aGLqEbdM9dD+eW2zYWAvT4hf+OhEDmwVE1Bv
QbDiG6TjRZ4A4C8I1VN5tX5g1Deb/M4+iYjiJKZPxoH9/IyWXZAY+QpvZnx3BJh4ZsbsbEwwQnlf
Fj9dEMtOcA3zgArPBG+3EY2RA80cvmVDc9u9HX9RZzz8JGReDvOuQbh9TgtwtoWTnPLV+MH0l5UF
IrrUa9e7unKNgdlvpBRlPDO9xgyZVzh3j3TI+ppt5hVe/BwwCGYLQHRUzk8m//Xir3hAkJWkWyTI
SzlpVVkeZBuBkB1XkfnhgZdw16zmmgbL5Cq4B1wW6HFSXAPGVJqrr7Z9ipKicytjyzJSv7szKlrW
3yCO9fPvdTBmYDIYy/XVesxKJYSx3SAVUPPZl47VxLngnFvgHBtpbMSZEJg2bK7iYn/MgDachiLM
6fANZgV1OqXMjKDIQ/gS9yXjkrob0inuCD8fucLJIlAlofHzOUjzjbsJ3M7TubkTxv8sK+KEheDV
JYcurUpzR0ex49Xo3GB1yNL4SQ5vebfGOPNPnwgi2FskqwaHxYU2IAgqLjOWuF5i+450TXLBPuwl
WTi4h+TZnjDc7wlxGuaofbCbEkGfkku+PseAsL7ICjX8MXc4tPFEo0qE3FDlguEsoZY4ZZMbP35c
P+sPjedAF6DGXu8t2r0avqC/LWhvRkfYVGd0Sn7lmxNHwzm7FhlMK1ar04ofjMTzkdg/pgYvUEhF
y85LZzEotNZzhj1FKeh9tzAXfWsi7UvckC8RJdHqTsryinX7ki8kd2qZV8e33GbjRmHbDBmCt81r
mDprfbIJr+01Ud1ZDicQerA65Q/5ZpJ3/FBwfI07mXw5oOvmhjUWRDjuAEuR+MW6irNdprtQcNvD
DZt0VieYx7PCsM400JwArz4vFFdu8dcyMsxBVKWGYubed7PXbcopebJ8R8hr4gf3N5g4z3iKPbgc
Y+BERkID3LjHIguSvX8c7gM/OiZNdvEakmRUkqV6FkMSJG0iMqPtiYg2mAoilVI7I05rCC9bDFnX
U5fEqTpusjszumVfyzLVrGauAmd4WffVzSoNmGpFAvNqauiZs2+ogyC1YvFekJPlBtCHUJ1fKsdj
eUzbNl4EPGg6KfmEAEswEIWK6Rl3wPN84Dp2TG5TA0pBQ1LLpONM+Oca856f8ECjPkxb6YqU/k3B
N6wfsGEv65J9IdEYwoYd+YnXGSoHyVx2Q59NPbhARnadqDhMXD0oTEX+y+b5Vz87RKUGlErUMIc3
P1ZBJ4nCIB8twaM9sgeUKrDWJVgCXXfRT2vXCixqb0MOuZkMruPVpI4SSmenVS+2m85D3UHdKC72
OgtF5k+nM9FvbbTUkQY0YVA6oRs0tg4MYuouQWCcsqTdeGgOnyoBz1/kQH4gGQr+ml/AVLzcO3tm
zTAGPGOjl2sHa41qdZkJv7AXua+RmGqxsYeSINCK7ELRvLRoZB9jVPgyvC9s9/tB2WXhrLf6GLir
uEFZEJz8nN0+jmAtpjp626BenOLY2M9xh5/FX+a6I2dkX0FOfdRhRYkHdigb3oTCqEA1l3mv+ey9
dg0nF+/NbcuRrp/Lxz6I6Pn1A0/Axwcst6IhYydo+zKNpGa5SeDQQmZbzoJrNfh4MpNUrfMiceuV
xrBdl/jYjoj6JW9xTmD1J4vcphEuhsXYcrEH7xUdgsPtQBNl8rvL8s5/vtaO/JJohtpRyZZsTV1o
MndjpfDkokMAQT2bGBv0ttiY3lr2PHkqF/1zgc9euAVDOM46noyJ+ox9RNKcIJUOm71kVa7CvEDY
FvJeGUZxW1OEwbXOIG6wbegqFd87Z1d8SxtIEkBwmTUtXHIVYChSM+vPbdxp/SWZEioJ4Pinbls8
UZizEMP+jCzl5aFSpz0G9l89A+FzlT8zav5UG0iiBiuACPZyDfgRXLWsFGG/G5a2WK2fviuNwaUG
zGRktpS+pJPZMJ6k5n2D7qo8J0fzxwNOJnuBAkZz+jOoB1aSF6Pnggs75yWLaQ7e241IRp9G5KNO
o5Gh6l75wcCeU+v0x8c4bP+zm2WLH+cGclXFWdyO5XKvf7Y5l7G7ZsfVnmb52/iL0VClGsh4fEMc
XFGJTdY91jZXYHfqHnO2F6zG0fNONqq3LxecGBRS/Mzr/KDgjf53VxT/bhKrbBodfW5KvcNxkTuL
sgmgM0J1rfPeRQHugNp1hjzdmwSHzGAqp1fsDsZTYbac5Nrr+nNhI3UOetRjBCDcetWOWft8km4/
AHmv1M0rIhwKhdcl6IvGYFPycOe0IhGk0cKKVyD7ktyWGEqdGMzCWi7BuLf9bzAKFCQ10L4DsVpw
iJkH3RKj4yGWmen+xObXbF6/4ZPM6o3h6Q/UtF6iT42kGsZUNkOuUUaIYSyf0KiCXKI0uZ2l2811
+xvI+OH01UMC0DaoKuKRwSk08jyM8o4+9bZsBjQa+QantTF9+Igqr8ksjUurnEZsWMd8gUDXTFOu
IBlkj1Mem4i78e/3gdfhsBybkmKCyMA6o+1vWzcdCvm2DT26j4nF0Gdq5h4L0TjH0TqKrIVmFEKx
ulmozc2E3Gp1ZzSghux1zwGDdNMYIj1AhUNUpKZnKa97cjFbMYqx8OtUozsFc749DOKm+5lsI1+X
DiJpcMvt2eCSAOanRiqSlWUTtANgEOsLX6TCPPyyWb29pwBp+wuvpMcOM9RL7HDrsBLLF3A53a/k
TcBMl5Y1xHDSZgOwQsLT5HpfGHw0V/MpICkT+NnZCE2otDcFjBIdEq9YXNt9l/+zqRpUYXEaAj6M
qrVFvrSbm+QHT915XxzbF7a0/52sJePiSZFHcJpe1qeLjBb505aR8/EA3npfczl8aQeI6WVU9FlI
ZQRpWiGr/IYWsdd8XCQqr1CgH2a6ib+Ys5rdUOxOxwCF/0mNJm/j7mXiqMr3v6hFxy6AoLeka075
SympQnZUkhajBPepl6bsmKO5PeUTM/08wKPvmHDv1XYw7K3NdzfqeR7cxvEYgpjFLtkhKCxggD5k
lVZN3oaS5v367OOiSgRtE9REr1HPp3XO5j/iEIw8lPVVAFYPluFZnJgki3Ze5dmTsWcEyGKOd4nK
BRN9k+7OvCXVY02XjdwncAdvaj4sTUXik3zz6rGtvTHiuxpp0ixQvrD8OR2JrggjwUZ/uHisWKUW
ur2afvd3R13IWPSkQm+Q5jAFdB6aWy3B82kxzJMgpVRkNYk/ERfe8VvkcWo+Mka0vriGK2j6keKR
8cYjGqFKC7+ALSSxAuKfaas6PA/Kuu3fTTsZkimZu2gQg3IW5jztkEDtoMR3110uu5MCnQqefdlU
ytaNy+WEXA3VO8PXqKdzl4QwzkDCH5/QvEYR1WyWrQa8y9w7aHV8NlEi4YhCJH/orJ9tYZKh6FBM
fyf5Pb49jmlLwSGbRmtk0+R1XZrf8iNNAvnMfyaFxpMASYQWanidbZEwBGkujm0OTGjUBbe066pQ
aWljcCbtJ87as4BalFZ6VM7j/iZ4c5CQHc+yTm3FJWalNZhKC1V0r0FlgpEXZD6oCOvpQAHCT5F/
MAkn8grwBzuZzMXUW+4l9Y9xdvLuBifgh1kCFvWoGQEfmysYb06M9e2O+1VeAokaBa0EnjLPqDZm
NVQ2yvRDgEZW52WPGt8OHWbqek9lqnRMy9gPnZZKjV3dj0y4VrVWz/Web0iScjcdCC/3ajWSwHzi
hx5ddZH/9jGTiTzxFtbvl7HGYiynOHLHEk+IThSb2pzb+9lLuC1UENi7bPIrD+WzBJ/52AqZ1NaI
E2IVmyL7hDjRk6AthrVzpMmCT7w9aL33ufqI1tvpNIILBpCwrIPRYUsWIJZAuHUxQRyhPITrLIeE
PQTiSp0iKsr9SSQXgUhP6OY43TjKyqEuXacYjv8hB/ANr33tZImAnJ+489O3LuzW8XyZI0m64Plf
d+h+e3K0E9j/k0rI5rYEPECMWTq5zWgZgXqUJHRCMfxkSu1B4rLODiQTwtvGnuMvbnOwYyUj9yjO
vuj3E/YC3VCtKUgAADTdFThgDmKizpdeRo6MYFooTT0KNTwNCYfC5GxPNvQYf7zaSWWisPCGdxmZ
CFbxjXebx/QenVMj8O5y2KxJF8YDs9VRbqb3xpeDLqgqCJG78TJDQQXj9LKaZ66fsid36lSHyUUt
7Id1YkVoEF9F+ATNcRHBjWdyugWk5GGHXSDNvEvUNoc9Z3vjrW2weA91M6VaySfvAplr471swdhD
L7xtKJJdctlMFB358YvGNCtIgvT+0XAPMbVQHz6xYO9T+xjIp3sAB9tu2hTAWWAeHi2HbEDaDSdc
cExcsBuIA/f4WooxGFnjEcfcY4unOrjuOYgcGtxGAU/asf0E1dvz+WHsM3X7HlwNBBkFKdGV4qtd
Szxp53TttcrFeyHE4YZy5VzRnBia/qDiCUfo6jwPlODNIgzwdN1VQFd1X4mMqbp5OgCk0PHXyudA
dFR4VnmqEaVQ+axJJnmZ7OGZI3g6ulBR8ZW1aPaWSIYYbR3E1bAbMcrW6EOpEVEmXf3u0UewXPyH
S1Jc9JjWQAYqBFZG5F4l4Svu99bIgTsjT2WuBXa1w5VkaUEG6zemlczZKRrkmh2w1Qn/MqCAVDQ/
/8YzulKtiPYnCcE+Qewz9PjBHkFMW3wdHApDYxiM0UNSBGjJ1TSkO4xn3cnUGBQrg/Myj5KJO6CF
HaXSdTpoFQmU64t4i1UXogMPLkQSyU5A5WZTts6YzfoOlDmBhTbCqFOx3K/ZbGO/h2zzNPJt5Dpr
gTyulT8o4ddSiFO9UAmsBEvUaR9HqSk+oMtLwkjvoJiAycGJH3ILLF0YwptmEm3XZE7IISdEMW7j
Y18cXhnd2koO4QaVXQWIkIz1y2X3vkMYQyXdtDEO5EwcaOx+PtUMTcpUyMAYiBly0SEQSc+aR1hk
T9+KmMkxER8WVdy07+Mo9KYrTiU9DoSL7a26hRd859BHAxlvKW05NWxs96MSoRkA6MGf6dIC5tbL
mbpX3vRdCeQeZF2EZiCGZaMJ/NLZC/yjsNz8MSQh8I1ONiMv6R46q9L2lHGOWbm6BRV67IkMbHwT
udUDDZRdG1KJjGveZ12wzwOAPPUX6M83VwyG4EPrauJqD/UXAXpUt8zwUzJAJXv3GVT9gRPd1Kl4
PcyiCQNm6GSj33a0Z6+bj5K6+bHDFpxI5L1WiRu04W7uAkMqFWNj9aHsg8s1saheIbbE4QZEYmuA
wh+xOzX5UustiTjcp6mIzY8vGYvjsjZfNNubNNNcX6jpkLpGAwId4ljBosnQNCEyffnc/IUvXevF
LWbsJfu/hP5kSsLCwvbMYk3eWDgECbIpkgeuUemIpH1Fno3AY706bD2xKm0i6vFiGO3y1sPmiTHE
Nr6Ik8/AtSLxXGzJTCUr+4YSDi58tnV+TDfUdVjTvmu6pULeLxBYmLmw42Jn8SuHd14fJY4r9hqD
2DAd3HOATx2rTOf++gGzyuFE+nydKqIxP0TZKx0amxzbBLuWgoB3sYoLfEcDHOnle+rTjRWxQhEZ
hBom1w4j2b00GOKN1naTnParRicYETlMFgZO843fIEfAsXD0NHr3G6Amq1Qn9M5JhrdXYP9dkFku
TpX8ugnFb/860b3YyVbVLviCMzE7aYrgt6Nm+JdPOE1gHygppw2dRfve89MQRWc7438Uy09G3ZZ/
VcRuw+p7LXcQcfJM4/67b6XxaW2t9i64ywAugZtBTY249c5Z/NT6qiYL9YpszaETdJGXbL2L/0kw
U/UerzN8EpR6NpJ6lH6/n6m2tdM0SOe6mdQD+jH5uKqKsZMtciOtwxMMMNkEdPWX3fx0g5HcO8eJ
ireB3aO0G/XfCBPhsiL/PO6lIaMFfilCIJzcUbBwLeTJM2B5+XVTtPkaIWpLmECtmrVqbu11p3QK
QH9xL7bFm9WPdRQU3YVne3cMg5AME0V5ajFn0g66oXY8n1op8I+eFaXogpyplpx2KJuusQaxltoW
wT5RGKuH9vlM1zA7H7vf5N7w/HNl9cgcZfVAZSDQ1lc3YWKbdnCHxPCfVL2FACYBiouYOjV5eWlM
NxzN8JHvkpd5tfhun8OMJtm29lk2+Hhdk7oEpqBQ8+60vUEpNFrUgrueGuDDYwgvgVG9q7W8quD0
VTSN5Om95lMUcrC71tr+QaFlevLyF5bsebqAA9HfEVpbUxldXGik4U62NP0HZek7IHCwy33PsrPF
1LL0B0XEXCYWJ7JJTVuCQspCA+pRily+qv4+4zFgQbp1bNOW8R8NIRP6bbUBs2Nj6o6bMeiEzv0D
y1LakToU8aNsffkbMQsl0fqyokfISzrfN/21lyD4gu587q122bma0fMaaSRR63DsmO7kA/HqDiYJ
sbXfliAeebGS/HZF/koKhv1jUkoBZSUnLJ43CBDzhd5JLlFZq74A+08P3o1m1z6zeI/x+HzDEmsN
9RaBikDV14LYaImbYpjBG9jLwyKFMJpBphzvsbyz4gyngWsDEoNfV4i4PjAsRjB2P3Sre0+VU1Tg
oKqh/oYweIB5qUbChodK7Sa6dd9o7yC6DTZ4D9wWwEFIwZ1CL3N5hCjn6K6OXiscZGn5xhBLx7Iu
RUn1WIQAAV2eh/GMDUYbXmrv/HRWi95esMHDySVOALLVAGXbX4cGInwznvlWigAhKd06E9hQ0ASh
ArxJyxv6l/hRHd/R4OLlLxPohxDTmVMr1jzbQF35+KCUnQYHXthaTLVeWg0qoEKLn4kyXjbhYs+r
syw0ziNacLZH1FGFifL/YLo7zNb0ZQmZk+XBa8rSP7f5RxMWO6HH3QslRs1RkQfbXUuGD0eHPOeH
BC5FTNJ74QRHBOgws93v6MDI2fQkdnJ5zR4tdhjWX1iiOBCnOr377s/0fGmCP6Zaps2Xa6UarIob
drQchfIztFrJmcDKyrpfkEKG3lzZYISKswXGGOXEiBvTvu9TJ/vqC2Z+au9v5sFUIAy3xlJLknF1
ArYCnrVtpy3yLqNYMX1FLsWmQ372ZCXZsoY4CF0SjUrLSnxWa3w78Oi62xIZ9rE8BdeSwi8CiaUG
9GmJzVc8PFcxpXuT5rCjapvy9PJMd+JefGqohweVEtVQL7JgHz+O5qTESDLzJewL+90KbU9gFgp2
zEoQBvzHUixjIjRFcd0w9L523xTapOMOby8UF/xxlv5u9Tvp6ijep6AGfXUs1JQK+oL4wkSZzILH
AMEWmNLfL4KvT8NIC9ATdUFb3R880PH/Ucz87+w1cVjEPJ3LHQeg7bYviRmYc3noB+CeJdBqfHxn
RTn1hATP3S/4DdTHNtvG5t3eP7E77e9czTyTGJrFNDEhxEpiNd3Ii+0luXt96nrMbBngZl86ioYb
h5oIKKid9VB3m0dcxwD7KMwJgyepLW3uMhn7wg7ajbYyEUFCiLFd7sFUQu6H28LPeLnV+UdWauRR
/3+gnwNUAUOw3K/uux6NijzTlYvrzcUgn8aEBbFt7T9GlF3iG8XdzQbiSM8dwzop8VPyrXiryvQ3
lIuMF94Q1Fpqxprf9MoRXvXssfVQbwPg2zoV/0amxFualpoy81Q8LmiN7jnWPbVFX9bt+w4tDnJE
niKTW0SpYgd3RVPlzcEG3tUYNDW6O/MotgNXHhKQNus/Y/QvjHOtHf0dvM/I/ZbFC3vuerhYUWRT
v+ZMFtdZye3Ga2qCUZCwmwat4h1PeMv3Dp1AcCE28IxW/p7WXvJPbVFmdU9PWKQiLk4CCEC1VE7t
1PVpucH4ks92fMgKQd0binbQShEg0Oncfz+hX80UljXPtF4oxgQ5SwF/Ip+6dCE6G4UDdVqIRpLx
t5TDTfPS79kFTiTCJZJsWi8qPGdO8CF8LgiqZ10sFHdi6PH0DUxAO4RkQk/tpqxMh2yowEoFEhy/
eDkmGkVlJBWB6iJ4LA5pGVMKLAusXYbmAxlTryn7jxmrJeUTQrfFPngqmZnO3b7axarXEMVhZayr
bXlNTqr173bF2qUOyeFdAEqkFhk2OPCKaAWm36Ud4sS+DlCXHW1lECtI8/PUJzzQkLBw4jQRJ8m+
vI7QxfKYGP46egZn/qti/vmh1418yTivYhKLwwAJ9t9CLH1Kuf24nVI91298MalZD98qkl2fHXQw
OcJyDDa/a+pEUQ1lf5v074W89MJluKobSpdYlJ2FZW1eK9L2bNHeBUdCmK6/OcW4tKwElon0QPRn
3Fle4rd3umfNr/zVoqC34l3IzNGFJQqCDGKjdU+PZ58725OWYaCF7I6VvGVqv18S6ehpa/iHhz9s
QSVsSxbukmTGTc6YII1AXNysTMNTg4rbvSoU2rFh94FgcNZ7or18g9nWqCH1UAgX3ACukMD00kbQ
QWlQUCAXHCTZ0uiKQ30bBcdvmbcXucq2JZd4JIuJtCJR1n2g9//SDMrcvQ970lN1vDlyh2GpPSsA
0LSonmF65qfqeil2DTR61Rk7xzsOYezFPv+/BZ+uc4htJ2NseVMxleVLTWHnOwRBNQhLqA//GnDe
SLQiTCj0NpaEqLRCrLLGpDUZoDgo9iyw2bj/58v2GLBo7MdC6kyT1kDnxbhBWuEi/T/K5wUYW8mO
J7j7IjuPChSYn0JrwzOsj/2dXxddMEFupm/C3Ekz6lKMeqKG6oTN8hVtaqAKSYO4C15PcM3+1AQ3
zPZoUF6Ssp9fJvVJFFb9Z5x6D5YcTN0eWThvImHjwxPyKO//qvgxa+Y/tAAk+tAb+6wVLnUTJsEQ
h+j5pA8eF8UTDS/1jdTuRa+P/XSUTPm3ktWMVGwNBxb+gi8N6tNGA4vclVhYlHuD7s1mvdgXDYv1
kZRW1/VCfkDXMSQkSSF/6Eu/HD53GSgB+7lWYx+zg7PSzWS78jeBnOL7ltWbStX0+S9r2HjdZDhd
I6gg8bY7b+oiCXlfPpKx1jmuKEHilr27WFBFAMxYclbnC1pXPVSh4pfJK0KoL76N2FL4fz5RU19i
aqbLWv6vrINwroqfvCBTx0xgm8AKP3rhhSeWg0qyaJ2y97B3pkCYZ7nta2T2KFwdzi31ivF13l1b
VVs+KCvw5JV5faCTYqncLlxnRKMiYj01M0iNSvduA4ZVfwHyo0Gp6/TlkrEQDcWB8gPsfswO8V6q
Dohs/5TmKe1TH9oDiLC/G3UNEKx/lxHrLC92VipvbBPchE5lvFffCqseID11MgZCQqHI3MUMRfu+
QgsElZiNbWcPh+qNY2kgxLweVBFwftdaQp5/K8JaMLef1ATLH3HcAV1t/vJLeXA9q+c+E4W8ZzwL
pb8R/NA7Zl1ddQfNq/3ChEKJVmSenLXbpN+pys+8qy6mIpVE/qEkndnC7a/4iOF3MImRfTYz5UYK
g6gMfUe2G7bboiwLPmYjmRUFGPhivf4fpvZ5JC7+soqSE5j9mp2WH4DrEOXtFj6wZnURTCx3MUFG
Hm6uvF66NDqot6RtLEpsqq7nIOuOtRZm2PZAt+3+5LTYfr8UUluAApYnf53pYqd7dkWLA9nugY4g
i2j+DVrz8pt0lGwPrcW50sLHLtMFd5EFvAZ+fzijTmEyEuNakRDRpZfc2WhUG5HvavMx+sCdiQ0h
GR5OKC6sW5OJ5ZVu2BdQS/D5Aeul/bNfb/Zijv7Tf8Ru6/NL/c5+Gr8h88wmt2J9iE/Ip9s83Uju
B1ZOAr+arM3ErYyVWZSmZO+KcSnf9LVKzGMT9C6t6d06vwxT0KMsBHNiXhR5o+fX0VS3gONAQjTK
S56s0RbUnpxCX+EMON0/SE4Rk+6eYmeT2ae1A0eu47lnN2hUwNtC8YOJmJNDMosMh/eab1cztaRX
iTAihkA9BFFKObfPHIDuJgXCtJIdbLHellH/xfG//Ut739xpVQ5uHF1zXPL1fQHOVTU8GpmpD4Oi
Atz8cIfM9ZyXCRrp+gI0lCMhUg217DU40u0OKlTzkj5JJbYqyq6/pZ3HbwXZMQzcJKDuMSpUcF/u
WNGGPpxWJa/S4j7/o86taBN2TBbNz0ElvXdY21IeYjiI/SOjn5bPLqxWrJgJ59/7i16pKUpq7wV3
cRUg6yun94F2Bzx2pw4D8csFdE8G0H+oRj78BG+YLSTqM+9R1FpPqkarsniCt5jWD3cFaw7NGGml
ARCPtsA8jsjedU3kA2MCCfivBdBUFK7yLIKU7BvInkEftseqIUgaqhFAG3M5tUuzpCWpaT8iAfB+
c/J5hgByLR4lYH0UeksFlnHRHGyH0ocaWdzhFXfJqUZa4O9OBQk7WBWc4P7HzimaA76LHFjDyT6E
hKkblPG65/hMN6vnlEqYdyMgZCxNV8UJxWL05CQah3eZmbBgun3JbWa4hp9T6E15iWQbO18PqeZr
pLE6WY4qQyxn2EOnIMyjxTuPZ7nw7GOn9prjkz1Z7AhNTa+fRSWV09NgLR/aE0Me6s2YGEzWpDQr
np1Qn51cFKmeorq31L2QTtNKa/sm3puDMDPDbPfXQgBc2ic5XbjzsjkSlFxuOp2+Fq1eIEM+JJko
yopGjgMgpX38X54wA7yue+sYZbmFeG6rQwvN8fz5cISNojc6qo50dJ38CwNfBA1i38T7s0Wm/qVW
onE81hfdWV/Mv1FZ148eLQtqtOTfpoSsp9xMr9cB1ajLxMZ3zkgvqQHpYjaIdkcubvDIiOvTot0t
GOOVouLNUIX+czR9DRSm5bzAnkuAkkyFc36FQOpkG/N01O7uvTRyyfv97k+ztkgvgeWewrSXbHoe
rPz1+fiCIqk2R2Ssd1fWefdD6pXNrVBgVt/iWckeRFlU9ZNoKbYT/6AEOCdNzZj8Y4q9kvLvcLFk
g7a6lRi+HUqdStZ1ZlA1387/nHFav3/Uovmtpr7WNRs1DS4Lfq6nuOJNyJZWeSAlvcputSQxs6wT
TSX24XEfLWjpynP88Fhh2hrdLfbKMbkXTcilHiQ+3xgAWHqqm/qDM48Hwum84nylwnWXmEMRshgZ
RFab63TvCjbJ/qjLnfReqUlldRqlU5tOzlRu5Zl410usivj3wDM0dIbWgIeWC1E52PYm9tD8BSFF
dop8wlwpVTyX2c0c76ihJUgFAG3uEhckBinLwEy2tTTNfbbMHZbnHSRtNdOnydwS71WKP2t5i0ia
Km0MKBiwWYTnYDQ4H6PzbjQTeSMqzVvQohbhvD8hpWYfCnFgstz3nN0PEMWXCKp5YRAR1+Bl7bm7
YRH9NEc3SQG8dXNB/2VvWTMoxi8KdRmQL2QayPurf+ZPpM7Lr28/mFhfw+LwFStS6nHhJt9UWNEg
fkW2DuEjzNB/fDzgy8LW1zI9ahOQXrUY/cQDpCALweDVxeY3ttWZsJnYY5tyw1TCEFKzLB2qhXO2
VaW2XIhEGTAvLyUBciJyh5Qg4MRxylN1FJOJXtNiht7ARlZgkEw9ou62tCcWnWruBHFATFpZEeqa
Mz1AVrF0Qa+juyHHKxt1l/yf8DGuyAUiB7fOmoA3B2bmSj5SMzKRpbOcQYr2bxYOgR1LHo/0LhDH
EM7F+QL/HHJXiEKstZtH7fa6Y9bc6piUksfovKB9IhLoRFmXjxhKjvQrjg5frci6ruEbkyMwRPmH
+D1mnnB03N4KcnLnoCUKh58KEOE3WFbj9TyQoq1saHVEWXKcNl4yjoh/gMpJFlDMVJASDlHwc8vW
cS0TUwYthfvdI4KgeHOn45DXDLRAwngWKhhMwmrMWU1ufZvWxdcqL8CqcqY3FTXWRiKfgNpy09Ml
v/IRbtFYdrn0S1eLNVPIgReCY6id2qaGKeb0qGJ+ZSEYX4Y71IchmUxEdpkVZ3MXUI5+SW+lpCRn
G1qW/Q23AvWwIohwXq+bS6bOJHuHKtgbJjvKsy5q5ePhra5IjjVDcprSr31d5CrkoEMbWjY4Ygkj
TuYVcBgUB0mQ7nxPLNs8YxL0i5YUhPpoeNZO1ap/51QMUYdoktpfOP6doNKJBRvh39GeP4Zq00t3
bFdy1T5YW97ltCFbdBTixZwlfFqvPwTaLmhCE6AyWej4j+3orXylWxj3YXhSy4OsSNKCgnAznLw3
dziFQvGsniHBqDE6vM7h3GQNWGtp5xnjJceCNLSaITSm9ZUKcOUnS6iZRWW9jgBz6I+MLKthcljh
dDQ35xB/k8Nj/O/DK/sO+ePCKxbT4Vs5mX5/QRb8rNaaIF+ep0YRhY/9S88BptRI8fCCsEpb8F1z
Z8956hPM3uMGuKLmdm8ouU/mIrVuIrmo58rTD2ASrnMKcjFr5EfyW7yfcWY4h+sS+ejnrrpAj317
CZJFt0tX9ZU4ttfcDryVYvkz7W8dIV/IBP/DpjrBI6+YC2P1cFRy4gs6OMqSXDXx8Jl4XBK26qtK
YF5zixk2Y/kjAdawT7fjcbzcalyk7E05JAssB/UY8Nz4EkjQmQa9OTIzOxLMrfEJ4xhs6fNx9aMx
HwhFHFwUaa6FticvR39QDkn7swSTyJjSjlCzg+yM8hvxdn4qd9Uo8Ohv4KiPoyjLsQ1x5NLPk96c
+NpblAdFcVEdlV/XC0YdFpTMr3yHQxA7UsnNPjVlPaSuG8zJeDx0NwFF4maZFLsgUxv3e33ZliB5
mYGrTS6MAPmdBBmahCNuQOXz8Q1ICXIqO7aiRAfHvQve4hrpv/EXQG9t6rqnlOndWZHvsjjWvMvb
kj/7CRLLd3TVE/rQTm7oAf0fTDi54ucZL3YQ6EV63leF9SVPRdNRRTfTkGzM2A6otUBCi9I8szB4
ewVLDlydPjzsPAQuUQ7fVVg42nr5/Irkb3qJtQYz49o6RHHo1ZijrpTGVOTcaQHsqAoqiquWatfu
+e/b6dCyfYN1LkdMVlgifwuC/TicmXoTkB8JJDw5UmEJHi6FTIRBe6GpvQj83wRDaOBAoyFbW8Ds
fwlDnYmA+s9nUKRcuHw/vve/7N6tSNSqfgp3KByX9cvL20GieysHrpz70P1CAvABfcgdg/H/7D1A
VBB+ncmiiIONiexORqtuCNXjBsdTLqB7wY/qb1TF5aFb/pmAhw/j9pfk9vwaX+TlDHKkO+TL4Y1e
Rge9gtzQ2eRMfIjlXHP6jQVWLJGHBplyEJWc7mYRUmBrN9TExbVscGwrahXSkLpOtR3Gs6yn4wbT
0/GrpTyuscflfSnVAnSGgkJyW2LKEBNEB+onRFNXi/pw4fuPYM4spJ1fAQjvHIIR7wjlYTcLVEZl
0wDQ653eeFOVH8mGVgJlLkd7ux3fXhOrlFhU5yiR+GsdbOPBZw8CdE9iFf8K4BBW9EerOQr9fXLA
So6zNVR2wYOkt4mwhUMwWlGZvDfdY+rXftmPEUARbqw0u+qW2yNNdejtrMx6nHZJ1Hzs54LxHRTR
Plz+0poiEvOfnFl+KVbTj6RPeKJlcybpNoFGo+x/Di5ol5q3Q/GBFpgNCcG60ZO2CNYsOz4JT39q
F+B/FhdvT+hN6dglP3nYsazAcdV2KjlwpAbMWWycSCgBxmtOsQiZ0t3Mw6+Rw1OgTnBRl32raYCU
j6CoAUpMNmaTeZggVyampg2NtPwa+RZniso93mMnmDu8Z/wm+3XAUqg2+m3yXttcfXNmtgnV8z2/
P+2hzJLLWEDLzIxaiv/LVFS/cg9IWHYjIfeA718TMc7nVaak1N/ZRep22OYVn7+EFlw7ymDMUKyi
zbpVR5/cTcs6TgicZCzpCfkBBl93olU8LJyUx8ARIYTl4WGu0hRflxfw2liRUrKkbtnIbwUTe7f5
KWiVwTi3lBE2cqEmaHPjU3bd20bK6gvm43dFyPtCGaibsHHm5jERGICYMdlyATqSgnzGHw6dmtE/
9xCPhp9Fa+DdILJuZffXNcZrmlf4Prv7FtitB4fBg6N5Skb1/lenGY1T6zBAQMVwGT0KTOozalsn
sxLWToQs8eOelqEjs+mqqLz8C8pA+UqKWcN+wz04jtYYdoy5rLgKUFb1lolUewc6p3xTOJVHYwKN
ens92IQEEGW9626/zETMP3N2UH9kj0uvhyTQgFfxpOjkBTtltQnvkEWu5FAabG5XNvrWZFHrSkdW
a8rwbpx6v5hwl2pYUQJVmx2qPVZCZ8VFBK8uv0sgypOYl9MAbRNsAOaLiJtJQ0r2Bpwy5HU9mkmD
2R/xYavQRiai/XnEz0e5bne6aJULXfIn2kN1XlGPLWJMSfKrfCYhDRUdPatFMlGEowhY+I3yxmkc
MImOGzhojdPmVFMHI7Hu+8/HMfmW3uUHC4kv3gYRF0/Lor9aJ1s8nCnWBt6PvgEOD8Cxaqry2/6P
cmaMvKt/jxbe38Vri1D3Q79wEmwAqDBZgS8W5Z/kM48Jmwo5ZaX9Io+kCnfxI114ESIJpEwbRUoM
rVAu8WTKfhhTf3XCgRGXgJ/E9ZpqNfo4BxLp+JSJC+wxOVKzW4TBcik5guW9IvIlsuYU96f4YiX3
XncO5b1nGS+u5+39w4HRJF868as77E4ezZPDlLy+LfwAsmQO/l7OA7KLI+15/0o/pXaE+1+2QYx5
FuEA/WS7Pq6J0MSXxFii5g9Ye2hcEs3DqGzZ4/ZqZnOKJOhpp++81QC//K/dwnmwy7NlsqPOF7yd
pO/FqFIO4+KGIDwpuWE5zpTHffcFEOz2ZMB8Uy5lE6iYfYpaDn0ujKneE66ZJLqUbE0SNAXPMCv+
jVLaQUfHojpKOAqSw71rIyreB8/84ay28X+zzsnV3Np+NRk+QqfGN8HRwJsCA1S200/6PxKDY1Wc
vy3yowK4Tf/hLU+5+OvYkzVicpvtIkrMXWw4YBzW2P2KPMnkbfQPzqgtIB78AT++CPhSp6ukAnIO
fNg8U0aGIGVjqH3SpNavKDfyGs+fazGGcrQDuZhBwXBr7Rlymvb/dOcKyVPyKvn7b4+yxqnuyFhv
k2TpHWEsuH6//gUk/qhuG+cE/9gXCggkNdtWBlSWfxXkZqy3H7Xa6GhqS5C6FluQzK+Be9YxSd/j
k4cnxiU8xyUUJ67VJkn2GFpHEFuwZRl0ZxRHY4Jsp7Iaa0bLCS6njXcqke5Kzb2B8J+K8Jya4/TS
6Gc1vIL85UZcl8OUZLI/Y3PaOYGDcPhrBRaihMKbhEE0FY2HsK/o6pWl8Vasx1K+iH4rKtiYEdw/
Wx6qQrj8YYG56dme003G/M1JINC66iepGLvteXKnG/68ll48ceTXT94J2qgpaQLTBjzarNqBnCWw
EeIw6YwhVEuns3Oi2MHQimUvy8HXlo634eg9M51p/yyjG6LVVKoPZ1AUMPYgTdYo8ShvgVNw9TM8
Jm6QsdNJoDv6Vcug7o19JRCwcF/DZBmQxm5TUNz4sMUYBlXOYPkfvaPP51ELdRd9P4EIxDmCNKwo
gBoEW4Z5P4lpBXxTXF6HFJFKodUSVnbZpCodcFrGy0yuCBdlJCGiVJip16lQlst2atRfEojbI5Ux
eKWEDyQ8Xr8pmj8250hWXI5ORVue1YnB4bTCEuHI8XmYhlP86p7bhePqytaEpd/XlUzbQkLNS0z7
hFCcziLLfvgnMx4J2e1ltnvaOrhkF79H/71lZeXm8Btx6lAocgTCu6cIjQZtpt8QK0lBq9+TaJ7Z
P0t2RcpK3bgObVnYw/vcEXU9KgptwmKElgfLgXmF9d74Zmg2lELsuhA/+skeBYmGquKqsFKcBWP+
SZnZRgs75UmOqNwzW+V1n0PqOb4VwKRbfHUOsD9KhIDp8q2t30VnynbYv99QCRCqv9LOonruy7WJ
2TTgig33NS822jhGVF2JfkvRTt7z0AmsYyoEB9V9qFpBvME+CKJEylVq1QUBLNXdkdDMriwqiqY6
2jtDBWJsjIlZ9QByfuTCqzB6yZkr0zjDL9HoANDBVaJSKMokCSqkU4ryrfPGxVz1OB9k7+aa1UJ9
Vskajc3CSMk85mS6CfXWV8Es2MT7pZco3KpUIWSqj+Y/+aEFZ3Ty3ojTrV1nTfSnFRrWczfidFKx
OLLj4RbVZvht+7td5BbVWKfqOe/uzYRr24IZkLZy/YXIpmZtkY7nEsUteMzUi7Aw/ehw+KWF1vP7
GwJj/Mgfbcx8txqwiX6epyLq20G1MrRifnOXm65R1fTt3jCwfjtiGo0h96AicXCdsVH4EqZz5kML
EwGY/i00EW8AstmZCD6N0rD1CHaqNvZw4oXG54OpdrHqMLf5ihTccpuT0tq6qSYe5rosIJvQALdR
qr8z4Ul0rp8PNo30S/1kB2i9pSCIO/D+zkXwFUlsgrlKQiEv7AE8iBIZqbYQtRJn/bM5ucuFSRCd
LwHsfy6ScnhE6/iznMmxBV3j3GR66p63Af8MGdBc28Qxh/dVEk9AO05hw5RE8Hq2Hi0hWFIfLyQf
qw6UrNRHbwte8cWrgnPAMJiG1sgX2ihf54MHY0iG9ca7Ecrl+0FQfwiTYxdq7zik2Ga9DMWou1YU
XyrfJ/UrA2dt6WZitvtsSZiBVbqLTkI1OnyQWWmx16ZKxxGuvOWokth5Y4g9Rwzvf5lBLxeMp+CQ
FPMPrsXsrnbulWLYdvrB00MQE4zI8J5nBhf2IV1qeIP0rS+B7hnWAqJ+GSlcItHmLD7seDhmkcL/
IyYZdluwDQBuxArkUi5ot72R2q+dE1YK8h4/yGHzCHNUR2aTKgD3g1Z5r6hw78jXytc5i68mUVuk
E2wZ2CdNYsIPFdSJxsI1ZBzSaEoP+ypuLEKZlHlmThom7Iz2EtUTfo6tpFZhKdDkYyOtBT+jqUDm
EaapUGPbfQxwAc2oGIWgoAt36Jpu1gLvuJhWVby4YWscVgfpAsgn7/6CP6eMfKU4l/xdf/TlAz+v
5jJsv6LQig8ywz3NnCy8pNsMgHPeGbdlTonRp2YD/Oq8xkgGAYfBSJVO/ZoGBaapbRJbMdPDQgSQ
WVxiC+YigaampEjmJU0FmQ3vSrTACuiBTP7XXFOqGtRvPMqBoF00YDvbkrmwUP/KzrGxv2jeqaG5
p4ATnHkdzD/cxiNlbSSVpuuvPXmf8EwqbN/fxE3WR3wX1lwCFEGgKiW8Enp1EK5/eAr8ugFhNVrY
mcA55Bm1/uG4gkMuAKz8bejjRkI031Vq++WikoP1B03xCf1eDwclwCwZy2PMU2wyQOqnDcNbMo/n
qlET3cTHsTdvbM2KHxEsq2RqzHdu1m986IAgd49RxoboUDqOhitRs2XFrrXDv/oZ1LH0sUstr29t
I2H0xceAbGfwmTy94fiRtqgjaE5pPuPpaMGSAerIcdHfKdeSfPDdbvgmp/QB8zXR/AvAxOeuAOVc
vywbeMUC9SATwcIuNixCjJ3C8Mn8xo+LuSKKfs2XaYYS4Ywe9kA8XrQss4XHyHv6pB4fLan1G/vy
iaL8bZQPj9m789SKAEtr66t67iPiHwDersbcEW0aZgMLXhn64KsE/QYICZzQ2mo47XgccBka/0rX
gJxsijzdP8LQ2XUHAOPd+roZ99ibA+DfPtKJqSGOdYqmLUsSdwLAHomG9ELcownDb94K8VsDLeNT
eqgC8YpWObnfR3ATjqWjevyfKy69vOIzsnTsRI2Qoz5wZ2MT7KaGNQe33jKoTu8o1DpkL/i1iw4t
ZotumMqvsCFvRDOw4E70AcAJ1LS1xRZ/IGhFHV85r01pjLJxqhKOrhfH5dO/N/ABgS5UowSbsMC2
xmw8l+fd1F4Jdl+mPnJxODjSh4qcQv+nUPjzEMiIb8j7eJpbE0zjW4l6kz3mBMKKF5WjXOn/+Qf+
OT3YjnRyTfDKpDWHniJIcIF4XcWJmiYqjDkVjU7nFc4x0OxTP6jvVRWVAGu4380WSrp+NPyh2wTq
bghIB1cX7DQTa+jJaSGTYa4GJBPoS5+pCjvRH8NvNJQ5fbevx6OApCdz1EMp1XEb8FYDqMUxEYGY
56/iAT9frB6xRoTxRAtAdz0Id7+8/k6MmGUK+m9da5VfLPNpUaSkni6hMQEXQH8xMnj+E8Gd7guv
JsT/YiKHhT7Y3nCRyCrC/SYpuw9k150VkmAmPqGVbA8jDfcZIrxXlAEaw8RDDcNElbWiJ5BfKmPt
oWXKN26kB/FwNoQ5PSgv1YOAPhQoBYV0LMo6ImgbeQPihTKo5fv3jPuKjZnpuoiX6sHWD3iWG0+b
J9tA8j+ExMtts1XawdBNHro5ok3BAyhg2nYiEFFL6j8SQ1SesZTfQL5IN3pLN0+joRC6bP0O1d26
aZ1buRIbF2+jPkITEGfH5gnfpQ44NSQ774wxVvKxpngW+KXYfH8WonGmzoG8kB0hawc/+CtTloVu
oO8kaz05vyMxTnvanREZ27qKcXlgMplyEcPry1K9VOE+tzs7NZ2XkEFgU6z1yrNQwmGEQ7MFpJ3e
JAdhuo+LtDBU6q8QkXLKd20YCuLUvHxRcByitiISpfsYgkOh1YVZjjYZJaUYA/SA/wThwtcqwoaV
lzIw7ete9vcu/icRDPIQJAVQRtNysRG440XhWD6rQ32QamWTnRWGdK1e1OblygwGQ/sQJL5bScrH
g/EmZ2oOY6RdHpBrn8YZUtufjZdwh2PWCV5+iTt7yWlj5+yZGo2OfMTD2fCUmsbHeuIBH5IvbdhM
xtN+QdHie/KQ9SzkiqmU8p2a7jsx910TWYsVpWSBO/blAvIezDz+mzjCFIMlVPNkOm+snTDMgoZz
e3pqt70BidZqhrL3tVzTtXelskv6JV5GM+sy8//qZg//49Y81YJ73n4GWjAfbqUkDm8JJ54Rx4ql
xmqjrSfpqJtqLldEd7baM8UQExBc+753iLSmlC3oqPlTZIeiIDPwQuTJf6MZ+E5x65CVEKaQElCd
hqF+sM0Y15v+OQPAwBXhyGigumPvAwcTB9l+7BpIZK6Zt2WGo/48xsS3gfKSqrXruryPn9hGu7zT
j2lLurbvXFLVCCM/Jfy9hccKdHhEVbZNCHT2/zHBNAazTdHE327ACK2/mpWLn/G6a64DxI6VBGS7
Y1gwtg6fgZrkpiq0SbYYl+CaDdyOmd2PlnFbspVh3ePgR8TEu4qEgOHOOxe1a5TUnRZHRIVTad87
bPjTPaezeCiQb5vwpKALvApKEkqZ8klupCNUktq2kXaGqpedNxzfjUsGiGp2uxP9xSWLD4f6wHzT
zJnQnWOE6c0876NelBg7vzVMUSXR2+HLYryXdupOS/GRWk5sMf9yOMityQ/t+J/CnDeiFDhXr8uq
i3f09YmPgt40IUlPoJJwqAbhTa2rbit4nEsanqltrIX+zdsSVkUnIznTDJjV3Yu2QGkWrdxAseLt
7O6V0eY54EVgBU69KlErjZQEtLB1iUjDrLdM4v7EXB9M/N36EEljdwoihhUyVNC74x7iUThl5HWG
meWvxyB00rMGulK2fjAR92iabB5Go5BH7LuA6Sr96ZZZAORKIMh9jHjhHKfmMrd+bkZj5JY2jO/T
8pYvO9/5lEE9qk7OYhBoU3/mk1dwoaHoR5jhmKKdC7+aZwl1GnePxBxmOmBK7fFUeSCfh6dl+G0m
oA8KN9MralkWuu9CFgTKiqDjKjlapOT09qjBDaHw9FuFcx3lVnI5Yv9BvN2U6VmCMSJRpNtkWXq/
+YDAPUdwVUnPdKQw/TG0nSlRxbg1KFemEBfre7tcvR9UrXzmIB72bIFYoF4omHQNHboTDAkV9H5p
nKvAfkEER9t5Z75meD1AD2ozKlouLyi53kXso4S/mff+kiATZKJDXWZdIUfCcfAGRROTUy8wNxZ6
TB9OUmnD8LUIoVxVy/q80oBaGjGs24LJ6LiK6opybtb7eTM5uOIO7yhQpt3g1Y8JkDcagDxjWMZY
Uz0SjQsGIJv7NaNRuT8qVUXDvKcWaJb7+ClAgVQ1dnpsizcOk1PlPMA4N0Ek71X9DFR5M4uhbZXB
pAvLDb990gAQH+mX6IA63kiOSh0IEAIoYclt3V2bOfhSfanDcmMtA7tVnT398/Rqo/yzAcO8ci+C
BSVMBnhxqi1lXZ2v/1JfaAt40VQM+LDhoRc3N3gqJ/PNivDCHYT1zk1WDb5qdoiwUFIvmhONbiV4
8e8DywPCx5GcmDY0tL8hdqpSy71t60kuH25JjdoqagMGfwJQNJc00asl2oBWjoZWh8TJk4N+sveT
xlf8qlGncAy6huYcyvTRzqVRpoiXzu3h0Fuz83U0kfpCZ9erIeX5xoj0BRNJLilgyzSEijsN94j7
P+sG5CA67WbX1tEII1GAlCIxBzducIYnGLBpByQgVvTVtQ7LWba4ZECF6DUWOmejWtJjMdRzRjul
bG/5Iok1KXLF/F9m9A3hhaIlki53sb75rqhh1ON1yMvDBJMQKsiR972TYTvWC+a2DVPUyN1I4RGZ
zKU+fvttc4MDI+XE/zw7aurc5+BbxY+qDUXdmDm+LKS0OZy78AHvSDo4uraboJJEA4OnXcRjK9Nz
wouRXSpa2c5Ef24QvynCB2oeOlUtrSixhlITETDKfDK4op7P4tU2R0gif/4S9APh4qeKL66kTEza
TxQYkiQ2MMV2P8L+R+TjjNgtypfv2nmSXaBun5n2nHgeXnwqTvhd93wP+RqZ6h801vVAzxdd3KKU
XlEsxMFjsBj54iVu/2x6MYZEMYCq9l5uXCK1rdPMYun6ZsJ3XuamQfrEdH7v2uCb+B2VJlILnmMl
AAUhZWdCYmQIHeWnLmiExRNOaaXaOUXPcJVYm7xqsZT3gJzm/nxC53S62C+wVHmSYmKFzOyJl3yS
KOlWP9pmOdut7Jy6uhloy2EWCJcJ/buclMCUOZx5gvzQpkQITEsKxeRnSOYsgSP6ovkp83vc/RN9
fBDJ45iQfb4TXmIS//ni/5Ivf9PNT0W/KUlKzm+ZHdtR+ClB4qPL36GLswthPiXb/ry4mZi9be3L
jJe8aR5xLALvyi8tqPM1Mw2KPfTeENzZzHJ87Bjbrgi5s5B6asfwYZO+pqap0v7InNfNm8fzN/3D
SEwTe9BTo+c3D3z3Pc9ta7dmleaXe2vGaCnIAncsY219WqINHeSgtkPUU7DZpTeZCSv6h4+WhUkm
2utJ7U8BgOQtPdhhuowKDRRsMjT06buELApj1BKHWXsOAzGfrQkZQQl4uomuVh/bxlApRkOkcja/
7Ee9HUwx6Nkb/6tjkDyJkhKkWz8p6pVVZQ36RQq4UVkiKEY2xLb+uxYI+U5a/WO+M+aUt8FUXfdp
YlowGocxVMS1gkSj/guf0k21BMGDdWKBwU9V991CyFb/cJYc1E/4TS8zvoEyOmsT8TOwIaZgCKrN
5uvKNWdt6yhxC2lhtLncNFgIzjiwI31yt4NKrQW8BWCJiYOGI0WHWzhfvz5Ceoi7H2nVIgExu08n
GzVjI6wjd/dbz8GgbcMfuWjopjr5Y6AKYKqFcWdCxjuEJ85rVhJb+UT2YCF3vEJoixS25aJZJrKP
dwFRdmXCXht2NKSsJwNcHTwRs88y8b4U6vXif9k2RW84O5cLCQKFyt+Vg1k4qpDNTG0BGoGRS0Fs
Y5gKZtsKCQ8aeBdaUVbTn8oC25gkaFvLGuGpa9lswgweCkHarsvps4GBJ/62m/v1c7EbxBilRp8F
3PQDWAR78dAQsIm3zq8tiNJi7dt0TlzyFk/wdD630Cyl3xZjts54Ir/TiuccqsA/krpz01x5NTOT
YHitaVqzePK3VbwgHlBVmfIs6bq13AMqZ/kvSjYxtoKDUB+neZkCZwhb3juVzn9Lx1/JPtCFd9wc
xT41qEaMcsunzeCU/ESIJ92r5UOaVsMMmyGUllBmLN6yq8tBLozPaNKPISP5B+RZlydmOe0IRiLT
JMsObDM5ENuMlvnbKeCAPoSxzyhH9t07JxXidzM0hpaMpsjVYORbzFph6Mz0TIm4L6jDzHEKi2uO
RNdtAxHp0FFDYy3nB0gcNrd83f0LqL6SWmSbHqznhTWqE+c+4aLjQXyGtrnddfsIZ+46juQqfMey
SHm8H00N4UTiigrSGChfPaMihEBOUgaVjgtETTvCi8I+m2PbM0U0ORS/PFh/yNd2D+7QMpVEKeDJ
Dx0En/cQAHKL4oF73/807rqND3PTcYW6X69PfzIlBktq06EZhGL7gfoKeaIe2wYWqSQCBjIr1C38
UWCIRK35+vqIMCZwTfgo/P4+9AOCLwCASp0UAtuzPMRgkLOZpYZpG6W9oFPXEu0+lMaz8Tmcizsp
RUxdVu0u8Bwz2HWbdsy5F/YvIk6hroPcwMj5N4HedqQC75YnfzqjZ31chgh580Uyn+OxG1v4tWbz
vwsb8HNjVbySTaYbjYWGBTCCdWTQHymVhJyzt9kRsDzOxl2IBoB4rRjAM0QCyteSdu7eHriSVEK+
dQnH2srFu0oj8Unlc7n+124PR3Y4aDtiVxcCFviXavz87NY/GihBH5g9tbSjxGu7uSlxDdAzzD5K
kVtE+ihVIVeqJW3pPV423NUlaH7O6b4U10ELNPBwwLjD4JJINuhq9ck+F3Y1jzh6DFnAgb9vrMfU
YQsJUVKJUXUJMlmKeY5suFHhmpxM1zZafF95f4KpK+VfRJ+wtqofqUkL/58CBO02050SaZItLga9
4LpZ9LKzhIKMah8PjqW8BKOEZm5wAdhUZTxQTtrHJTFi2t3Ebm7Fmx5rCml5AtVoqVv6tyDIdVWg
yRbOB4IiXPDHiUzeFkolxTVaEQ3yt9F04396mycSDpb+65V5cOguZ0TsSmkFmss1gbO60ZwUffUc
eBWi5YMJGf7uXqJ/H4B6tljPXf25sMRMQAO2OorhxwRjAvopSHljdcuD7w4u5lAgLm/pkwzbmAR3
fwMVcSSOTV/eFc5BfUiSEF0oMrzzLrVKyKGTUNnazrtQulcwrzzv85yAVxs7zoK89hMqMO1NKZZs
BLK41FTTbJeoXEOxApcHXcbz8HOZydAtiYaPUopyBslAD63XtZA9buaVZxWNiwh+sNQhVsm1BjgF
2venPdOxZzwgPr4Hk8cjcVQbTpHe6DBUUutY1FJguK/E1ZCaTobP4TVjSy5J5x3pm+2QiQOn7pfI
yzTAmj2a/uB2RToMviPIzc6Nu5UKRiN+UH7mUN8iNS640IABJd12XDVx8fKm4FqVL8E5uZd3FEGs
A/EnDbGOA7eLRkI4CtuAc8sUOKBmPZUEcUR+vdMfhjoP+4kGV/57YP7kqMKdWoF8/2+OpKu+I45c
2Mdidg3wz+kIA/jJQBOqY5479t6EDxMj9BCau3QMU/MaQuzPuvcNi9H55yAU+jLnXCDjOwrwG1fr
tvldmTeWcG26la2L8oNt6t4y6r9r4M4tvXACFKFrlERuuEA0KX403ZWTuLITu1otujdgTvjzpcCB
ZjOzZjsyajSR+zQiqErpYNjY1MSG6/LXFwcK2E/7nVAJ9mbrJF5TxgyQmZg+0ExhIXhpc9ZYrA1Q
ma98N8eNUSwTvLq3XAUS1mRaeWdzOsGM1BIC3SnqLvG5TmKMuaPLfBBIyJQiHusAMZLc0K9+Q3yQ
XwKEuJ3g5mrfXq9gCGtlkagjeR8FMQt/Ex0GXq98zTrNLCi2foz5PZ7kPo8mHdFlvoUE17E1TV9H
2LPipsVzwEQIwEQjiQcfr8asQmVtXnCCgw6WLTQWaQDuRlHoeroAT45V8rfisM78MuNOSfnloKXH
G+EBWCOZYILVaq1asivNbAC1CWKFpixfYPzlAhqah4MNkuU/q8w5oY3eqJfeggcnYrdaFAGxSw1M
Mgj0Sh0MXB05pVwUpauHsVCvnBwAPR/Awi952EYc96yxPSJAP3F3gAW30gavCTxsmPATIbqDJwFj
xA6/GCRl7xJoAwJMpddNpffjmYpBcdm/+Vv++GeQttZdHNy5k3Q1NmnuN65sG+UyLYsN10UJ6C0a
yEzYDgOeLznyHD6Airir2Dr9uV8YqpjUk4rj8k63cny4uW06Y3nAtqJltGvx1phY+TT5JhlIvh+l
16mqsOoINVO/BI4LdlgDWfyxc48C5ya4pXbJbuZ8TqzivR/ed8QN0GWN8ho9U0qdgMAKboxep2Op
k1ErA7Lm0FGnWulXNihZ2/xJjIrdrHluVwlZKazJ8/SnKAGUXin0BOnLXarn4z1bP1Q1NcAVGSVw
WZKiX+iA6X8cctsF0xVU9jp2uuCZakDyZ3jmA6OkREVQHonWSvy1i2FgL9Xws9jlv8Bva10MsqWh
jWNQZ5bgYcmTMIIvW19S0DTc4Hf1GYC6QiCEOazxeJ0bXS/lCzVtdp7ZS3VfKJgP1PK6MiV1w4pe
3jkQu2LpPZmOTZize+vB5cB+pBa/KAHgcO4vNbtNwI9hzFxTuaaBK7KPxpKljhGbwv7rUnYJMaCX
uR7kBYf6cgsyZmsq25kGjGAV2sC86dL1nK7J5TUGxaPqpMaosYiYzKyqpcSehMC4S+ifMlXRBYls
eyA5NMVS3dnE1LdITDD38M/adBu3OV7/z+INtAWnyFZjF35ptSeik+MpfZ+jZEFGF8/mEKlEYInZ
lPZm8ttTB2tQ3k900EGy84ErWnHNqHAPga6VjbYW0/gHciUzpxMexEDjlQVFFYbyACzcFoqfkNg7
YrLBZDMiH+S1Qi6JLzJZuQvthT6MWaO0SupcSWX2GS/wn0ikdt68iUqZQKebypkPmQ2pfLD94/3b
c6zOCKZoQZ+sDI7JErAmh3Yezx220I5G0RFFVJx/NZg0rujLKt3lzSw9FzSYli9WfeOFIUFyR5UW
k7yqsgCUAWove4R/IGmCsJWad7LsG5Z00GlhbxSPE+RyAQ1+nfaxpplOtNmF/Y0ShAtT5GQd7fiY
lytz9bNg7NnFBnPs7XrRMjfA0CGDS/NWXYh3n84EgdJ8OzYFEnN5JbbxvywJdkv7nI7qUo6bFAsR
p7uFyxGLiJ9c2auHMdyhN/5epjlM2VH1JKsLFBxeDftAdb1Oqy+sXVypwVmPJJibZC1iQWCgd2R9
HwsweZDmBJEfg8y9oPdXXdTf9Wb0f+3l1eSK9dP1wsEBkkVHqPdNkwgpUnvbPnWRxyC5E5ma+dH6
zj/lE2PZyb5tLl2dT6xJ+PEPLTzCL4aXMHQLS+DfZlW14piRCo6Ca2uwJ+gM+SzLrfX3WepDYjNB
irArXbkKgpXLzlIEZm+RWdmSAniBK51GNEMyI4wiIkAUcl9CpOkrX+4dGTyTgmKDQDGdQJ2Fh3GC
C11BSMK33ZF5ViZrdlRPH2hLQihNLCqMuo95Od4eYMIpWYWCudMjlof0EWqcWesUer6bkU6wAAVM
zd2bguWm1Kfu+Nqw0G9mm7o4mBb2F3jmqtODo76hapQcDOub3gseY4XXan2xIrKLSGkfwUMhAfjS
0++zjKm4RjYhmqfP/+gpOsICkUMVdZENx4ZISV7PsaUztWZPUttACFPsUUyvzijYFYg+sRwixZnI
2A9NlhZasRhDvXg4Q/QWhpFFizNdugataof1TPQYFNtZHr+Epu6N5hqn4q4twbQH+Vee2I0OQVp7
E2rCrFMZQdGDlYxh3KlrI+23pzCwsKGcq6XlPzyW8Ey64G/LHun4Je3nNx+xKC5WhurW42HwHEC/
jNR1HUOBR9DddpRY0ItgU9prNPpM8POEDmbTbbuaTFjQt0cLNw8n4SnXv9CN3kGv6Z5HnmC2fhvO
B3KYjuiXBWyB7xi4rGbctavE5OVZkIs8UrDf0wuu7+WN5ryKXQqT7xW/ZxCUiWFZGN1uAUvjP4lA
HOb2AZQ6pHfxdfgwaI8nCqCrTmy84j4bepAiKQICg9uasLSKILdPJ2q5rdECh//BqpIXYEF3jxsv
fOFJv44tEUowt9i+vDLPVAbrm9vXK2AStGF1nX45XM2Lxz3Dn+AK87kK8i9d4PhfhihRRfBUJyy6
8smUZIbgWZX1fNlmQqxeQrP1OqpjeHVAvHPUXzZv/7442rsAQSf9RPs/HZNL1YgF58CEt2AyHLhA
RJ5LJvsTwCRQ4icrDqrPdSeQmZNcH51UNF3UL8+UUVopdzWDVrnV2KN4RCVkEggWD8UtNb9CDP5u
ljLTxigZcvijUlROcvlDIgyvsGPW74sxPtW+T6lokr3lCOqYiFFwRBs/cUXm4zVwu4pUm/EHEk8a
5G1iDW3QfhkrGOWvw2MCqoHdg4bNi7bcEuOnRIoZ7bGtPRgjCzpfpBauVzb0JTK/m/449Njp/fiC
hibXB3CsqoOmZ+wvtDWHF45uwj3KGgG1/MkYP8KgrH8I3CFJrBvIS+Y/Wp4Pu3t/n6FV7e8nVm+n
8u/1Uv/vYUTnUT8DzHAfjSB1AKVMmLyWFKp6F1B+YCcjXK3FMkRlak5K2hAqSQ+cb4aEC1eGJpkX
N/Eo7OdWKChLTYq7gNJaKIIMV2WURQ6+EBC8Sqksf9USbS8A928cTYeOoJzOzgx95IF4GwPcUXAq
EF/OlOlldA/v4YvDGbbD8Po9CYwfwWKYnEdjGnGARH2KL9OsR1kHwnaw72ykh0CJvHSstFNwUq/b
fYV8bRMS0MpohRHpgdkA8kKyX+lLQBKqwVI3fbuksnEoBlyunjJvfdDgTsGXz4KqX6q8gDhyGghT
HYHdRWnW6ZTe9Pmxw439PMh60FA4TuqIA41RMh0jCCQRGimTrXKdhv8DWxhKVnIugwb6x5FjFzSp
gyutbyCQ8v+VDJTkydIBPcg6fEIaabu5ANFyRirqMGMAloiQBCTA2u0CkTD7OhrwhSN7HaT3l8Yp
p3wh8+gXUTYRQs3jaLBKC/T0QIg/6c1csHjJYEJZR6Dkyq//55SkOByoTlwI7piGLkmiQSoGWRwh
8iHdI9J72Omsr7T9I+5bEWTUjdn9AcoVZBOHCjt/46JEGwwj6KAnwOftQWh91Lg3w3gXM0J8/ze6
AmV3ES/Dry50HYXcjJfZM3vAqJVSUCg8J/LtmIDRCqeRTbeMX92iQGHu5nv4iT98ZXzXWmzvDtpQ
8nm9+H+jNOurGHOlOhSs0K+cizRHeqqjonnjZQ7EzjL0qBQM90CoYs2iNLjVa7R27wImwaHkjUiN
qmV2zn4peKemw7KdjtfSS5sw5UTB62zKry/darnI5QwwQmm1O4VIWjLGnSdJhUC1ZLGGj69Dp8ip
uSzpZY5KbzTIjj8k+1JNCS50Ope1FWYOtiDhX5e5ztVjT+aqUezcL8c4H7gu2HK8qSpV9FF864MW
Ono+L+ITzoqGzwtw7ubC43bqq6IP9mCYt4UKSE3/Ibk82RTJdFcwrtX2km+0NCZmhlYcDMKIU2I8
OCTsq1aGBSeRMI2Un6INTLB8CDRr07Y42rigGSp3czBxW4f2pAk9Q/g/lYXCwzvoQJIsOWOMbZmE
ZbnLS9fh7h20hbEE4pn8VX9A7vOtTxi6Anm8NyNcXxcapZ21Q51zE/D23JMZqLb5dz2qZoGPwOBy
PCVhvc0OmdYO4ZXf9oIkYf2huJwPO6WESVYdn0YeHvkU4aLgILGri50qiAFBgboakI/aS0UDNd8A
pHquWk31HUYyfafoAw1zO0VSV5rpuC5u9LXBx70dApEBmnTmSGqo1FDoxAvUXvo+wOHXoUUzGxAa
orjKctmUZ/+AehBRh+lL2W8voJXXMrQGTM9y/oC9G96at0KveqDVbbos0gvzqcedr9dB8ScYUcAZ
E9DWYdsG1ueaTaijj0i6AipaRZJKLKwYmDBNVOoLFNXBUsU8XsgdrLr2pasjIwbw8/Z0V0K2wCqu
VptZH+KymZsS9gVqTafzlQnkcYZoNjcPb4SB4tfBSIWRePfphSghsAEPnkkwJNO4zZXV7+xB1pF6
vXAnHmATN5i8W67+l0RA2nQuaZsON6yY9ckdx3ieNIIlyx4E9PbhZf1MBXsPLGThAe2KJONPe6sv
R7lay4kr5VVNyMuRb0C6a8+FPO6H862sTcI8QnwJ14mkvzZ7f3JzeCY2aFElYfjHqfXyWE/QoAG3
R8o5WIPCGthni1E9G0dhSMfdxukPL8aLwHMxMu+hqxaoRbujekDhvsWkCzhfbyzE8ndTgkhWr3K6
ZnIohPBodepOu0eLc070ogIsIlO1Cc2qCPIyVOdKYYF1sXQ07hujWplOwWDbYaHhYKz/hXYBBmrE
M9+KcW9/yM74jB2VWgxMt605Bj8fReP9fu9c5ADx27YZbv1GqU5d8muNrg0q7M8ef+eZYvD3Htrd
/2Bp0tNhxmzCRbKITqungNyNKmA4w9h0lOOmIiogdXxuxRC5hbdKgwdpm3So7sFE7AY9U+3T1cUQ
+SR3vTB7xzM5ERscqnd94BB8GizVYr94XD7I5nTddOowBEmbwqwMiRzAO9BUtAF6a+8y4l+ybJBi
ZBQie1M0r6Yyk/ZsXXN2UeLyYJfE1JXgNlufQPjo/r4XZrJc4g780zkxUXW/P7nLXsUBlbXO2ntM
MBW+P041/eFIVNUew59dCxDSGAY6aSx7iwYsNJ4gMJK/iWHGafUSxX7D/5PslhgHvjof/YNABIJA
ABdJgekSxDVX7v5jK1mFzPDgHRe+GY5WlCKcJ2NELUS0kF85IfwK+nM8xSjhxVMj5LMlz7ECmUqb
kD23w/7/JeEfpxcgPKNaNmzPPUI3BcwRxB+9AmEoGv3RXCV8F4PVpQZ3ont2FPMt3l3eCwNAm0Kv
HJvPxUK/9hO7gms6hIg5kGsvzfdg19rjQ0xsERgxqwfgVwfvItbnHnzsEP6l9r+8/CU6rLhz9xOQ
RC2Qe3SgQAQINqEeb5BuxYkKY6N2nxKXi7jDWIVCa2JyiqRbD4QMgEOjbIRKW6HfN4w2CqaVZRk1
uMHbUNPt6pukib00DfR2m1VgQ1x8iOG/obX7lOqpx9lE6DyaB6JKkN85RzjEOrHueBQ3lfeGbsia
hJs9OjNBN393fD09drB4qh+rksB9XND+CfnENnMgq1BnKPk0rDocqLFSiem7+pIDmMIVyMYKZH5G
nhZbAQFmib9G+h2cuXGHW55Beb+bRJtZ3lUXxISE9ltQUcnWMQQEv+XY/1+LkUmArY2a83KSXWVH
CgM+W2lwiQx18STKkMIZevYflYQyOUQqKYEDNVqjTCzdJoT1JIo6y2SF4OQpE5kiQ8wGGokVX/bx
tdex0h2B01SlBiaqBJm6uSYxX9nDStadEWQx6Yfo5JWCMhLhJpLvz3uESFT6CnjY79l72VZLg80l
EhP9091J9hW5TcaXeiIBHOSGxVIeWKvuz5YX9jiirtN79BMB7WfDyE4ZO0QEvORTbZ9hMUmoUMT2
20fdcF6Kt7Pa2IuzUO7IrZhf5DAb1Qs9Fgm9IatFalMdarEZcwLVIvqNiJYo2pqBtaCXFq2ZQfFX
b2cmE6WL4J9etiAA8833/Qh2nfr9uxVoRZSHFO8ut/VqEFrDr+Las0dGNml5NVV6CdsSLO7OPw8b
HiYhV+JVWVyh66iMtRNw/TDFXp5UnkxWoMAGPJIR/vGyUPo89Cg4X5gh+/v2so9JCgI3SdyhVmHl
1v4Si7JcIjQYkVbedPpKjjFtftMUQg/yr1JpFIe9ww9rPlFGpnwM6rpSuyS9n4i5txEDa3N/xu8x
Lbo2fQj7mNh+5kX85lWEf6d51gtoK2koxJh6ksZJ2Ut1+SM70WgCfsKKH9aIewVNNnSnSauvDH1S
spvWNzNhus1v6F1F2LL/pwvCg1trn7t47xzKcHizCC1OPgxn2QGIrxkNMfSDfXJg95+zrvtbFqZf
ufnV1x0GnM2kygPCgFuJ6K0O25JQPb5kIY03VbSGngI3vfWsu9c4pWCD5gANbQbf3YVB8g7Vp2fX
tmU0pxC+HG/nRZCqYTyXfy1Qit7U55HfLkiiMClFdDRH2cDU1AaDf3KkbQF+ku2iPTBqpb4966GY
6cRCU5VT2M8e3PTG2nOeQsAvok7k6CYBW7N3YDIZTN4EEGvBwOhsOhyiwW1QjnL+qRWybg7hXfrQ
wNovz/465c9kC4ziV4oWD0+om27AZ4jg5RWtKt3ejVwUadjhbH0jnae4GD6YZFqZu3/i2VkiSy6i
qSgLk07bhNuJdXDjkfqNJ+gEAK1FFW8uOVMEVGzwKBhSBMJw9KtUAg7i7A0O7w+XUccQwmZb+Csq
o9rxofWnyReDSLyy5VZtXFcQaA3ReDqxps5Xbaog8wA3X4HCstEC2H/DOfGggkEaVUWOeE+1gO36
x0HPA3YxUOKrEnDA8P5hhiU5bvBPB76ERkGDckdCWtANyHtg1/o1LuUuEYUShCnKQxcPmZKlMPrK
sA8PyzpyJp6863zeRYm/lgm8K1bvyJC0gGemMpEHfbPveRDg39s/Fth88WxKLyMduOIYvLl8GgoZ
gObNKOcpntjqmf8rtnE+IYAORJuhLiDBVPbp5e8h5EWdZkscUmAhxhiBFKKuiR+E9DxJ8L0UI4un
f2c5B1bD00P17NH/N/A0fQ4iOTtzNdoqkfaWpZQPTONupZXQfKdNOkBum5H0439bcvNZ0vwgK24d
HWEeTwpeM74OiBbffLS6ng463opeze1Zx1Ck6FHqRDQDcCIvKn0tsZ5uO20GSJQ/hHFs30QIOMWh
aGLuXPDzOgKxrrdmAzBcilkeWri1kfS0LrgcrOmwl2bAZZvMURYBMKWSqCqehRWEjN8es1cG71Ez
wYMVV81IpBwI0UtVq6PxFy3SEUX4UuY/uW7cUFeuL3oZxIU/5jWYYlEih8sEldRFkmLG24N7JwZj
Ue6H3jHwI0gB5Z5ad1ZXqkVfaq1GNC+VHFNGKWbaA0oLpNPI7aIic4ziw7/IegDk7i/V/gVUegQY
V/jRpYBlW3CKLtOEivhTCWYYmyOKDG7p3Q8cw45kitQu1i1n0JjXYmdBaDjAwIwGfRJWUp3e5esV
n13QFr/P2fvdecTz7KuFJLKDmeZPpK4ZXHlEcNaeECUlXNpYd75pq9Bu+BiMzWJuT+Z2aSlNRHgx
ua4obWjr98w1aZmNsnMraC+EB6W5rfEPqsuVz4KkG6iPwjqVWxEQ38wun04O26bMHvEYnJZtLbD5
lV/QMgkZCtXDBq+0X6Nun0P15pA+ASkpeqvhKkAjqKTHyS7kPnrGBlgjHtU/8moA2QAnUBH0PUsy
vREheXmsLc6XOiL8H73wimsOZOQI82OvQ43OElzkPl436a5/tYOSK9AIcRBjB1uP3m/TxmRnWBP3
iCHaWf3rNjP7XC2hglwLZQR8Ukhw2CQ1BH3ghhIXIM+kvoa3hZxPJM58QxTiNnAFEb+eVhcbG2Cr
jffu4Z/rr8Pu4aYZU6604EF009uGU1ObV6snks4f6jC0TxsGoR9e5oNHyouHAaZ76fwJho7iwflo
pyOSoYp1GRRkYiZRD4GfKqyU+ANZveA7w7Y+RcqYE5OFExQkszPRNklf6ck3IAESCRe6EOgF6hnK
Xun74qxepA88SKWJBiE4NAM3xkg2r+5MDRc1rgcG28ydSn6hc+SO88cd0r3nbQfaWtYGYKcQuDec
OJ8I/XQAkza/S5Aj6UsbHdlmGwUL9On03cMJHZxxJ6CG7oRNhVRrQVgiVNncBbggf9rjJn1WGSH8
+OGeI4vT7BYdjLba4ATD1ilGfddBQB9CXlTdduyPk/kqcpR3HLgFuKWDi1aHYnKCdGkKCNurP9af
8Diyh4LZxccIYNPfwN2+ctNeDKwOid7TbG3LiEhOXONcaq6i+PxoPlxlQPqv8xE+oWRnNSPcxIlE
UGdew+qfYbBvGLfCtqY7rT1qxfS64E2R38m9XiHweqGt1CI2IqT7ktOpPmh5+UcadqD7eSDgXrv2
M35TpbQJfkNktKTjlx2/mJCZ2XV+E8ZK22iKlIHRqb0TSeKPA2ootd2FMBjhkWkOzsfZiwna/aFu
PRYv8cTAL8AeT6yKSdtlQb4Feo2iUBG9HRhdhZMferjNxn2XA5jgCYBi27fCkORcMQ8GNmVDagbP
rjEgkKqJVdl57iWsl6JYItY/dA2Im6dFG+hqOdTDjSetTq87Hnijq7/eBDsoF5ntw11+ur8rZry6
8B2uQyaYlAWA8F5GN4x0oul0vo3HtAYFMEyqhk9pMJqSXccb9nQMy82JDP0HTIHHO0qG52DWZADQ
SEFt0JFuS51nZJ41ip7C93JmohNWuyQIct3r9yKMoL82SqnZriLZbXBk53dO0SPjBBMUknwomXC3
o5DSw1gZSS0vrKc7bJgBZ3rLUYN0E9ilbMz2EXATCxbvFIbqwmXry1Jc5udsjhoBueZKHERBtt9R
H4xJspM1+iArjCnivtSJZU5ymNS0Mcwh7lWE1oNFGsdq3EfA9YvmKfA/j4xrgksJDkJ46ajKXYAc
y/SmRxZfSCnZUpfeWKDLgHozxm38muvslsZGZ7qQRgo7RdmM9K6Rius3Z9IqMfAof9Ha+hviBTGq
rextB9tnQ4hZwn0EalsbS2yyzA+tBCxn94YtN9QTJtrc86opGnk43C+Dk5W5aZRwfMAQc0W+FhPO
D+tXop0SMJmK9GHBZK5WhEbjW2zGuqmSRlb6awLhfhp6RsGmWLbevr6OZf0S/rj0F2wVAAZHF3q1
k7O9Hc9mJyjGlKZqlnGMrJK1cfGb0Jnq9NGxMGe3gYDyXLxwj4gVdetYot7MxjBxoM5jnZU+fCZk
eN7VCUEsiY0t1PlitNtZXkxVosAVEjxNeznczVNgncDBWZnd+uzSmGRROzy08CZYSuDFi7djRCh8
242KryePD+MwoCtUmpuWSyXeDWGnYhlLWgBKEmes+c5mYNyUzO/w013sJVae11lxbZ4Z5tJlb9f/
ao31mYxwd9flXnELvHqz58aQizMWdsIDpwwiTGj43K6Tubgl3guHkyDw80vqa0fBeltM/u1U4PxI
HxLQ+kMSqmy/v4Fo72At9V7M5wqe8KN2DUMxwjQ7FReBpyUkZgZJARDeLBzgOuBuudKeRHFGmcT8
k8FHRqQN9WwWD/Pg13ZPJc19wdYbNuVOHRAvaFdqDFoPW01lDaNq31EVr1py4BwL+beAhHPMYRcv
whkXDhDP5VSvmB+FH2ndn6SKX5kvnnkrEArbb96dNt1CmSYz5O2dWYqS1H6zioeiK73ldz9N6ngO
cTBcpwnLEt+Uv8nkDJcJ1ZT71SudN9MM4LCpEmFoLfaCk3iGr9WgFW2T4RMbhlhZ9EYjfCbn0/4f
7vZAFeXhacDcnRF3unrXJYu3zkgosJW/nZCL7PoBW2Q/y54xZBC9xsywkOzkUdw36vWuwLJO08th
y2we9/lMbqKvPFtY+UxrENAgGB78iqFdEfBv3j7XAL8Wrx/I97qsEFo9fZZVuyr/7QNGENf4iYaH
M9bMuk5pGrDdvUYi7O3gvfSSf2YPbJW/3p3AhNLayItI4zd2HbtfZOJp2rJgi5a6nRwadjNV3fO8
3LipEvJJreGr0VCezreY8Z4gcAnmp+Jh5ErsjIhLArtc8G92jbW4gYDtCMgvh28b4s5qcdeHgW3e
uStFfkiflOyl/IwSE2Fk3yuVOjn0pNdKbJT3HmEB4WRUcrAjZ6qiONY/f1u0kEvPypPpD58sWBrJ
71V/5Ta4M7VL+lFRPZpSwcgLxGz8Bx/VGilEhi2O5qhBrXz3gnyBAmwKJuP+1EoKE5AObbpwOo8D
XIfeyV6HwGO9nlM8sQ9NxglXqLwnXb6jKLG9oJ5YFF4nSfeXvmetJOr94IS8v7fW4raZ6B9vO9im
bOChZymN6gArNc5WoX4hGd1JOLgVzfZhYqpQbiZo5/Tn7kLDEguWWHQiG44p8m+FtKod9jnvrpN9
TkuEBIM4RcMO5jAZIECJx9bqeChj93X5THCRG2HOdLmBFKFcbMWSthB+LijlLF1Z3UOsT5Me9C2D
NCSJLTS8pf9PSnCU/ozi2deBjRbbeuzqXpd8iHtMBmmw5pmBP7U2mofxs+eAgjm0SS26l2zrbk8B
gwNNR2rFo6r8K0dh5y7vpi4eLliLZreaYWer9bm/De1AAC4pfYOyluxNTHP77dHFxI7U7YRaeycB
k1JCIsRGjU2oJrKbizcxhyhVMdixdLQPAMgZTTTNZ3Wi21J3rp8x3gUXWl892esx2Hsp3HxM1OZW
Nz9MV4iJeb8AsmJI7sK/KwkiJLk1GLZfqifH5ioWBdbraG0mTMfBo3gCnmxBZjXSbYGGI1P6l/Rg
Fr7dLvKtCVMXuEGStVkTYcT3ikr97d5EGL3mGkhFiUiKVNz2dVEzcT/PLglI6brQwPeHKoTqzRKf
+U6vm+PHjXphVqD7PDraDqiRviNk6IhFraDVOuH3KZ6JkrEcQzizF89BmFS7FEOxTVY3ugODWtEw
lzA+r6RvGkqxd/ns+HzdL0LrpE1B1liW7EBcBc20R3fqIWcCvUDovSlYy/izSyzgMefvos2D+ml3
fK+DuI6HpVKwyJUh6DBAHeSAVFwgCMgw6zNmV2/WAB93m1f8AZHYGhGGyLBhAbYD3LCi5jhTq0d6
CWv0MDDEPe84ZGoczJUuzyYcubMVqvFmEA4s++PiMENbtEK/Wt83f2Jh7YYAuGl6lhFTYSFg4af+
DupNRK11DBetC67237lHeZ/LeEd5uU0r1jXy2Hz/KOiWMvQgacrurNJXuBBdnT5lvoAUuysBOVdK
ptKisWzhYDI4+n3bIl72T0b6RlyVkY2hDKTz+MU8cRz5mXzlTsqe1z5vnM7XL3I1fSyj33YJHhga
KWEl26rvcyBKBkHn66e3ihIenGPTTCAB6HymL5P4onL6MIgM5OHDJVZeQpm77sVrUf4QBfgdfKgP
YA+OnJm6s9rQo8YhF2ZL5LfFQJ05LGvI6FGjo/1reFdn3jD6ztJ9c1/p2OEF24/ZYuJpxppusz87
xB0rZalBJNKqPWNMMmIwzeK9pAK1VWd0Mq45DW75VdjJ5uxb7QH0VWNFkLNxZ/z+eIlKaQsqq57v
1/e/MxbpSxEqVp1PSf5s/4XiK2X5j7eTVdd3EuRvhrqOZNlXKMeVS2gS9R5Ofq7eY7OnPNxDcZKx
dO6LeD3jLKLbZVittXlmX/q0nHWHiCKibXpSLU7eJSfKcgqGMkMJADzsbKuqzoPCZnbF8G9loCWw
NdyOPLMbV2Pq9EvNFAZEFCJnQ9oT5u2e1e1MM6NsDoEffULAPFJLHQd/6cqO+JUMIEjoXEhAvadZ
hAWalKzLeK0u2Gbe08ei5tDWHeQ0A+L5AEB9cwsYwHl41WWIr6U2ESpnakVBRpIcf0Y2E8f/WbK1
qO4403phx++neZuqhh07FjhIhQzznEGluttZGaEPRND4j3LhMLN17UKD+xduVTxU+NpV5USd3ZXk
OFF69/Rtp6C/SPqzd5fcvgpNqGhqmA3sR1vpwv4iLH6+TsrrY+QXngTlh9laU7ZEPkr8PYeC07IR
u7lm6RQMJdnp40fJcgf08dXdDRVzupPS48L9mjWLu+eU4K6xBjA+Q/cC0oBXcWSD33oGVSF3aSBG
LY+Wd9vLMNr0euTJTjrtNlXAcQHGrCi5c25HLKs4jBdz6o6NerS5pbwlxQ7eKFER+ZA84mM1wAUq
rmY0zGHvlhJSU71obprhbK592nEvT+y9AO1oUbG3ZgvsKRt+Akgc6OBHADtscv2gYiVAn+IzMDJr
j+rlU1JZz/l1Xu+LzmUcf+MMy6lvCCiH50Y0VIt1d+zg9Hq5VMAGhKNZGUsfIEBMZ/LFjcHOf/oD
SlMWJqMdmFp6RXAUDVK8b0BpmDVKRoPdpoUz83Kk8OmfqqAKGWU53QsRQA/AvSvk6kLdTGFciBXa
3bhw32dC1L9bw0hjLSBb/b+BpRGRTGOVTOJYU/li9HmMgzWMSyTQLV6XYYJc1ETgm+zViaFs5bRR
snbT3+i25M9uZdzVfIYP19YYVtDA8e2TVJTgcf7SjtNqqG/nEWOxV9OuLX51KZG4hN0eGCpKHOcs
nB8UiIp8cQw9ED7JoNHxIJJsW1+lIu9x6JmfZQjLNHirrFHL1q5oJEgS0pB+KC6VRqvwMgWQb0oy
tsF8w8bVfTzVkHCmo47L3YSIqKxrGlib+SdBvJyVxeV6PNxcYDq1EveBv75H8inNQ6O0VLFHxhrg
kGaaGNgn6j5w2IVWirRcMPYJpcgZZUEFAdloV1aNkUK6beQ2+ufBRGB/1D25w1LACHreFNiGRiQ9
SQPci2lTxSMhbhYMVJ7+WNh90RQlv7OTj6z68Ez/AYkUEYw9CQwkhsIsoa3vG+t1Y6W94B6XdDi3
fvFa2LBfsYEKNSlATlZmpsFESBjc5xydWMIxdvb0O4JmD5+RE/njMpOZLryhR70Wli2URc3n9uDI
SN9c1mF28fbTVumSGMJo0l1vdO2aDQ67CM8G+jykRWgrJvQYs71Yaf2EIj26eYkcC1AxvkyTqZzn
Vv64i4h5RWet24KFnGPyx0CPx8ElUNetWwB/1xu2yTzaFw1gRrZUYVWETRROOm6Pu80jprj9zV/h
+5hdzZVkB5hi1JkX8HnprzPZvgYQ1n5Ls6cY12UMOCFkH14qzy6uq0bNRr1WrWHcdCnPxj9ZKJ72
mov48htolx+RWlAH4rqV/WwqPrUr+2IFMlOx3wokq5Kd4MvwwF3aLI5v9PwfGiyN2X+L3OWIJCvt
sqeVXbexw7PfSCkJKPbBaWrtVJ+Zu3Fh7SPhc9YKyVjEGRFlNNGLrdYPsC/qtMXB+S/5adRbfSJC
waqlBPTHc4M+11SENNXjrJI3eeTXyxDNXsvGlAjBFQsTIXosay6sZ9owR1XnoZnHLiIuLRxzd5ZI
yrVO8VMrayA53hiX6ttLm0joq1MRpBzv27OEpZoRACZG28bWFn3KxsAmffmdO66Nantfc210Cozb
l/pEOKyf9fRKeAF12XZqjyGkiLFmYEHWAFWJMQ2mYmtESGjDfNO1UwCv6JcJQ/OtQ6oqv3i0sNjV
89VUpSu6Jhms/t7vvHdplSq48J+FWxdHkQkGH8z1qJ7P2btzfhCbATl4j+zDCM46d1Dcguei/X8O
6/2Z+UbgbAw36vqqg2lSBUELAW61Ycn/1vFRcfgdPP2Ulgc02IsACfGBGTiNrVTWkMcigVqJtvoR
xs2p1I/19efVwjzrL3bR0ydGYOhF0RDuCTUeUefpe5Wm1FMZCap8GS1kK6H5Ws7BhjzEhaJrgsOT
3QdI8gvMGlPiY+DrLzWO1Un3YrdFIbOxlJAjDURtP3gJQePkATPdTEr8RsdfxhDTMpZLUaSTdPgO
t9XNBbvh3xRFCM5v21FmLRcw3D99ELikVOr6FZVV/h8/tsOpnoWB4p/Em9cWaWIpftbUY0c4hTNe
Og0X/YnvbYF1kKOeTQjuBv9pqYtN9dnItvOZ86NdbPEdWHM51ZiAi5B4kypV2366aVr7Az1sT1eo
Pjvo+7e058ZbcDdUTg0i4HlRcVCcJbarbAyKuqPr4aJcrKfbzGb0BMiJlh9HkE6GUg1uZynN1bey
q5b+5lv31M0SSTYU2rZTuD9aHAcb8np6ZOp4zXCVraKPRRFJB0v4LyEvwdmkCChLH7pwEPZkHsUN
QLEGmZWpNzmHsrsw4p3mJVpqrIVuXiRWaqm8UhMo/cu1IVv+JLeX3VqqMpqIzBJ3Bg8dBsQLhmQ+
hA6aWERhfH4WGmUYk4ewIBoD5DR7MVh8Q2mk6942lECCW7cU47/tiz7jmb/fSfgqQdYwT/mOMPPY
Zrd8BUMGQirbimAPv3wN0LEvvSndMRBGMPaDKPlnN45Bvwa7if1Y9mrsuRvMO3nhpBk+BD/Nk4Vc
96IBFfEyeHpyZLBooR/ZnbvO+m3Uie4L1UfszADTtzopiT73HCaq8bST7uZ+Gp9gMVYNIFtgKLUW
VAMzs+26vHI9KWrkKOMWLBZAh1s/NAuIr2jazW23R+UCO+vkImwsRL2Mvwl/OMHutS+ndkgu77eH
K93XmFGnetNyXstxHbKAjFooP4dF/xyJBj/fNqc4XgVU19l2ybHPrz8igk62LZS0lIWTSOgZfXc8
8PvjAztQ/ZikS4+om8rt+2GFS9uOgAOqrJPKRyoN1kcpolwf0S2b4MFWabWHvA4dyC857tsmpfeO
eSl9c53NsXcZ31Pj/+l780x8GhACmabRoW9XlBFs7arqvg0wd+wb3pHR+6NdD2lpK2U8SiX5xK8m
Fc++v/bCTkfdhG/+FPAhHxD/JLqPqJSOIQRBScEJpS3hEWa9vULdv0hFrEIqqT2LHWI41f+7qGJD
1AcN3YRulISA2XFJnapjWZfOj6tfgqV5ScjjJHMahMxVuqzPbstus0iCioAOrqPlIDsOc5Xxm9gY
fFMvQQ+45PQGcmPYVu2NuBwkwODqgD7f+6N4W/LlJP/7Nq+v59CC9TZ0+kD3sAY0suX5P8/FX05i
3qpjDTTqy4IuWRjT8SpvNXFGwZ/QhYTdVi/+kBz+c1n/IVo+8y5yzOeAK2KUA5p8y0J1/OGhbAp5
u8v9VY6jUUBluBFZvRgekTv3M+6C8Y1pg+hi2UwOPh/Dsv5yFBZi50KSPvaw4ujHZIx2LcJsDbfX
LCatkcYLhmtu/8nN3HjXzQx/go19n8F7WOfllRdTu6/J4LeKtmqLA5FARobqUMoBAks+Hv2AjebV
takG1Cyeew0DwlJqH8y8UcD49XCRKaXRvqclbKcD1SbznzZj1RUHrETPq0bWJC3q/8j+bd0LkFhv
zeXwU6w28Re6PgrxQ5G2P5OYmkDs1FdtUR+3FoH/X6FRCSuPhKx2oZr9Izr4QRx0o3YJdfHD5W6q
L8F95Eqdg9Fgtcn4WYCicm3hJns2doiTL785cSg0eT4vTfA4pfKm06lFKDu7X5jzDTpy5HxFT6rJ
aVvXCkfO19GVrHsdAqyAtz9QvE8xF2cvRKPxgstS6HgXHznOS+9yV9C+oWpWHPEO7KTFegNkw9Vx
1OjUFqvk0v7GoHWjrlAu0nd/oTGQeQyjyS7M838AMtyWT2WbJt0OASNk3JguiJPYIh78DOqDNt7p
fENedU1vcOr8Qh2D7BKEvKOWrVY6ZHZ7I9oxnd1EYBiSi39jT3L4FalC9OHRt7/E4vAYmB9VXGA5
VpkmcORg7ie0lURVlvgI5VxF9QpwKJergjT+pVRguPMvs1JoVWQvJKEmL+AL6YbpcAx0iEjX1nbl
NWqa5UkVpnk4RkMX3kvhfpz3x2kDZzEdlr4TvsHGuUlwZdPXDzB/3bKtpHvoswcIVUHqTP47/Yq3
m1lqmCn5UVlUAZZ//jfgqolXEX18p0bCqbwWI2qQDbGJYrDczyD1CLxYEjle71w1iBQyfC6bsAHS
ERaHRdqYAuSil3SUhe2UQ7l6+ULK+vo4cl6neWTM5XPvamRJ9fbc84DpgcU8HW5KETl0STYeRIop
cHwo73M7o50X8wrkQRiOMM9jI4DtNnKEV0HjQ3AoDvxsAKf20b2Sv/G+A2kK8H74H6hFlVJvyl7J
a8h8/7a9CRYz/00zyeaTMNhc/RCRYhJaVAhSNb0WiXCPJ/flFF50NICiUg6Ss3C0bb4KNneiuq8S
m/iayAmYFS3+Hd6TR1LbM7fZbeZVr/01g4PB58Wripn6X02Q+ac97abp9CdVygPz57CfqsHBUXM7
j9GDCEqfUKBdXf31vKaxCG+tL/9uDf68sdFkiHFVQKwOAH3BHIjrPItHZcG7mKYFHYR/J+YcmQB2
QEtDpoDyvWCRkocBUBDEqRg7EmyFsX9cE55E9q/chwSivQDXLZWlZP4R4i+QafNNXwpIZolkqpRQ
ekcXwLJLl/eQ7iPZSh7CZvEyw3aCkKk1XcJxPQY8up2YyEoiRtdX8ZF+WmXugzmTT17LIgpDJy7/
qSkSV06FmUmuay8xEu/i8jd0bj2gL8J/vQwcYktb6qwqng64sDe+MqCfaOJ4jeqcwpXS2uJlenX2
UH+La7RSQKm7fVcxBAC2uwt8CDd7q6ypcmU0EWUoflYZHKeEw0nriDPv9hdzAI3EkapnTo8nyzF5
5y+M7WtH5O3WwYSwCMD9Ty60C/R6MmltGb0poDfyUsYgxCtBNDH2gjW0WvNON2KIwk0Nga5NTz+d
yIJx0nOxQajbKikV8uESDBS8RcfQsS4jnExAhs1c5DAqQ14p8g3QpmkTO41eUhnb1HJinjyIVJfM
PZWIMVDdJAbPGk14icIElRXHHuxHWyFdBo18d5CvzAWsRD+PUB4EpgBCUhcptIt73+SE4KwgAwpi
AeGBQRoVBObEQ9i5yaYyj3KLvtMQw156sOqE0wm0qhPeMOZJB7I/XpK20rAQpFU96eEKJiewdqAK
c8Abl0tq8vkPG7xnhSSCjB4zmRSSk7fhnIzOLXQFM92oQGU8svo1bUBubNlRk6X+c7d1l73gI+Os
djhFy/kptFHBPN+lPOPY+GgVjrR4bYbh7AnIqeI3jLd3VF9r8kTj+vOdjqdKOacu5ubhBVyHcAxc
YZ+71TRXeb3GagFXBx0JfFVMwTE6GiFU3OTQYQt2KLvmBLFHLdi9IHWn4D7uMxVL0w6ULvVNrrJi
YfDHk/A96/z80PAK1FfQiWa4wML5PPmBV/1Th8jwWBkVVXSflytCH9bSSbLOmlr96aDiysZQkKx/
2TRvJpLXbeSkM0ydbnIdGQOh5A86ZkV4p98IgkBPbQU6nMtX3MGUh/dW6gE8erQ2Ew1kVvBUmdf7
Y1sT18lVVCnuVwMBGFtr8Aiz3oM2ARUCEAl04Kp0Rv0MYWDGFlxAcm9uTCk+qpy7fAJMfQy7z44d
eYK5uxczDGDRiMAqF7tmglctHFMI/4W5TecpZnAWeQbL9lo7jPWuI6cggAaEKKy6UdWi6gCX4+G1
sdUqDU+Y3B0lrxuFzWQOi8BfEIAdRZ9z+d6bbB421b2F2EtUOjaqNbt4fsKzZCKh3jpUsTvUwE9G
tQf7uD+5BWc3eH+8kiE69Iw+1lJCimQl8m9kURnexDW3DHpoyDJvTsz6Q5SOlYfeuQflRpM9ZGED
7L89GL5KX/kyFVEx0EKdM4B/vDRh+/7lszowImt085zKCuWY8tMv/u1JjmfZ/oK08wcCgjXiViV9
9/B2DP+qq/kICtYbdFUVKHdoeA3ZIroaQCjSkl557xezZR6vcaatsbVNE3lDOBI0R11qHH7eg5Bs
FQES052Q260HwKEun4POrvw5/qZ7pFlFPko93eqYpMsNW1K1jOrgycs+Ie35uLxyrtge/6+xEsMi
PKNMhVDfV4ExYSzxEUIKt2YdrwUKSEVuiBxgh5G4Lj+pB5f6Bk/n3FpM4jwB6arTAtb9x+O6Cien
evqpPTChn4sM55XwCoCgrWtivEt7VZU1WQnjfYHNZCapn3ah0EnIzrD9q0FHd29hLuYLkDPEbiHR
Hb7JN/2U/JL/w2+bmiaUKDmxfxuT6YOUE7mJDj4QVlghd5Kl8oVWtqYpI38Oj+v4vw61kJ1l4c8b
NbC1Mj8Sutc+JsJief4O0a1g5OoDAc6B4Aj0GdxnuJf8nIQS/AnI4QGGrDMSKyajtDK5ajOSOYyY
ZKP1yptvQAWCdbuLlI9BrWlY8wmLa/7uyzxCxggz0+dKIujz4W+6Vs1pPX66FvKRc10DGlmO1qRZ
bFEOoLTw2J1L99RG1U0f3vt6FMVNYXUwCwsn1z8G+mOxIiGvKa37N5jj2+Qc87tXUdMWtTPnocfp
VyCgLzUpuiE683hDcpYG/jx+Hv8Zv7tRs/kFwgNRO+Anb/dd2uqnjnqhxn88/5baGyHTCcUrqN41
XTlo+DCphiKfoIps+j3U0ZAUTVcYA904R1nuVsYn6Tklt/lDj7496EOY2QB4atn/G4U1JB3LQT0o
JksABTb+Dql369cudlHd++/3asTBkffBSh6RGs3G8Jy/05h/xVqPgmtQWGqLVYMH1EgIb88HYyha
Lh1u+awRRQyEPsFkOobRt3nX/HW2Ba7LiwacjIEKAfoq49KBB3LRPKA9LOmUr8ocjQ6KylFB+hyJ
ghcCNDqqfP7WUmmg+n4+ZPaw9u8jGn0go1s95cKtuWgq9E1IOKcJIJv1P63aauyUpbotEa3gX9Ln
RHRejf1AMvnR/OMUjjIC9Qif4JjXc7tFrO2O5APbjrCgL6r42OjqOmKKI5YeCZxcu+G10QeIzqPC
Sv8r65jAsurJxjir1sevNM+syy9aYf2FpfGjjhuP57jo/jK4NYQ0451hyRjDRv1hBK689XyBL2n/
6RE+WMyxcEv0bi/mICKlD9U+whMmzzNZ5jISacNbiKSj0V23lCxX7NEV6Up4uG/Rt7CcXv5K6Jsz
Obqg3tOUxPIM1B2dmA1w73I1eeLsXJ+WokFPGM7sqeD30tVOVCuuj1K46WW+yBUKdTiFH0i2s/7k
E87+bu96pz8ZXYZ2dnezwF51o/gpOMGv1IP5Xul2OAkbVYZ27PI1T5KrW61ufttdezjVXXFQN7L4
bzudQRBeyOMshOe5V1HCfEaTUH5Y6SH41ccD6XLTOTbsZ38A/YYOV/DfDJpV2L2lxwE7/311TBpG
QnHYlSTSpDOq7BMICxFU262N4YpkbY1rX7q0DuJXCdYoeU8uqr4f94R7zOW/qf4KirGXRBqnJhbu
WKs3x6HUyNpTzRJpmdg9fRo03Ih+1Jq1OVGgXuKSnMBY2SmqR8XHkqElWKcYJU2Xab63qGdHRMiL
f5kGH1Jqh9saUZxOEOoh8JSYu2ikbWuA2Y5yi4yFMxORgvLqg4xZFEx4vK+D2yuouyz2YfnLS8Kv
Ll+Xm6ppuqzE6H0oPCc3gr9QCmenmbbW8f0iOmgWmscUMqOi3rLZ5B++3ft6pH85AYggpy84OErj
tn1uMEnxh6CnMY+JCWKBwrIPtPt2bMd+vo+nDucVzM+7E57ybtQJRUcWeAKWV7+Qk50LgHwTOnSd
lO1RNmnd626JI1tF8Ab2eQdLL9GZLYm5B7yTLqzBWQPfXqhlRFT2X6E5BPFORcBUkZbaMnzfocgH
YlAlrPj6+xrG3Rrp04A3n2yZaUNuRQWXqCUp8PafrKgiewP+v6yv4xylDblAFJ/F2YeJibLOtCSY
eZLoKGHOXVwii6+DGVC4/qFWmmXELcE4cLiEzT2lnkceCGwiWLjHy//u3ozzZlLqYG9+gC559ppM
OwfnxQqJ8RvV9pIVQ62E5rOZEoBrVOBcCY+dBJFfsBpoAG8cwL9c8qJ+PeocSJ/z53mpVTMPS+sx
ps3vAY3mDbXeSwdGTUIax8GqkKeWlrd18eRmzwCKuAhIu26faiyGaQz3933BaLREBrK/jzh1t4md
/x5UDAtFVSKOD3WGCRP6uOu7Izs/VpGk6r2U1Wdf8QPvZBqIbvPf04fxXHIoHE3PW1B4Ofwik2Nd
tBYI2oF2YWNKOHTBOUpPaCIjSIc7WKjGittUl2jkuZCZoyBjjbZYYQqwWM6Hf/Ix11xKC2nMCH8y
+WDeH26jG9TinODmbKck5WLpOE3XLYPFEUUulsEkQlP3x2rFMzsr2bCenmKl4lGeJU5PKVtJiXuD
OzvXy41zsshv77CZ5iUr99udEOhqS1hC6pzw5hWV1gqu50OFrS9E4UNAmBzzxOk+uHbgGl/AGbgq
PiuMhx3EfY+Rh67nTaLbqslNpqpohX4X98CFfavLwAOuCYA6ic2kYa75fG/3f9MoNgPJ0KVqIiP2
FKNP7ZtY6idcuJc8BTHO5wCIGAIqx0A+rZA1ONyHC+XKnnJsFRzv4ZrcsAGoEM29DQOWvYbCzufY
Fs7hrzWw9v99LWSAMmhigQo3mDSDGHzsxrmtbGVYQiD8e0TdGYTEKxvNpVjHycso4e17j1bty23Q
+BNqeWRUaQBcwixb+3hB/FlKCa6HYETLLFjTCiFilRS/frQMb66thxhu6ACfaH3LKD34A3oE6tJw
WJLFqJDGL2rN48x6buPtaAI3yVLKtDHMjktIM8hpj+HJyDgl2oYWPKYNwSD1WdXf0vXlIX+5ni/W
bV23yLmPNK+QzZRCbB76r9uDiLL6DnDiaK3GAUrWwg6sRdedeLk0mzGlBDa+BUu4+33lMBz4GExk
QhW8Qr3RuAZzsaQztN6H1GbyELiPmarHagzby6iLpOqNQX2EzezjMvCnatZzGiml2HIcSkoEaIql
zz/yivGfJ5LzkYPYJ7vBLoWEniD1B/429bzpBUqbh/fptIznQQUlc+e9cFv4KciyUK15Ut2On94t
45tcCo6Bbv1jZWnnELO6UyEJ/XweScvrzZ341/zMTOG7SSWJPHUK0okA7BdkON9QvoKMPEUGcGvP
M7z/6/3m0ZN5T20vDdLfOsCS/gy7V12Jq7fVP8Rbf36z/0ybbk3THOhYa3hcJv2AU89hD8tj9nna
PzkZFCO/iTQYDUSGHrF/aJvAB2EJJ+QVeHmw+rwMKmz8crmZpOPCClczPnR1cXIVglFzctdWUFt2
V7vSpztqHobE4VBwzpHcJCLOyyCECh08232YTrcY/g/KY2VGB19P0Q7Z0JFTCemcfvklX+Z/5fZs
EkjXllpuhEe+QU8665kUD64FvQLBSTueXn9LzYCbEJT5hMxCJV90LxBfdhZXukdYejzHtIhCOEd4
By6bjS8a4CtnQhS8PCyQ5V/Wsu+wRZvUjxN0bGPsp58FrgXqRIMcOZEKZfIVzgvFdHx8tof0idgP
LR6nKHw7S/H3tdSZvp8eAK/KSNksZLyflEgRVxYgYsEKQwP6xeArnHRsUOr3gkf1+vf47QVswsKM
4WbcYemQSWUcDYboMyXdNLDUAfHIsGVC4QMIJVwZT2k34XO6GI0x4Rg0iGVwa8D+qltTywhuv3RM
pPfumEE/VSh9S1oOSqZUl7DciLcH/ziWw1xCqNoLXPuDiabcLUsLlKyCuN3QXBc8wEkmDR+iOUqi
f1Ez6cU67FAWZCUBd1N63NKP+qs9q87pDpFxWQcvIRpJur/wts4WLh4xs6EJZ3jno693uuu0eKwA
W+fVr4jm6bCcLecueOAn88tTycYS3SQWq94/LIv5i4UM6sqLel29hGed0ZVfwTvHkMpB+Un51YUB
utDsswHsNm6BeN40n/AKBjcLm/Ys6Z/mqhWzNK/AzZSjU30itPTBV+1a+b/DvsTxycMiq3n5Z+bZ
vkYnDrYnfa6PWWk96WAntnnIxh6CNqdJosPqdorurQE/bhshyXfWW+f7buJrhxwwsGJGhqY3VgtW
+W1DXl1AXgtEmuY2S2SC2dcfpGKd6dv6eUne3gMv3xCz8dDGpn846utlojTKs3FVKg6HRc02tcgv
M/eUikX+hqjNvKyYIXdofLrTkEn10wIJCwCTZPYidzTP2JC8l4jpHc1ZHTwh1eW6HtIi92nNrlOp
QFaYHrY3z1vQLdox4Yenzx1LY9XhlYPEYR8B6LFmZzxmeXqmSMdsS4viMzxo95lW6BgJUXZCOhAh
+ism0R/ZbMxHVCSsoPHe7R4qt29O+rkehQgeXgTdOAC/ZfgBdlsRZ1nVtF0KTGotS3K4+Xv7Lei+
fm4V+gowXfBoig+ySSu5IMG9oRr2NxnsE7EbDFr3vC40bEwjSMxOyx3/n/h0SMKtzd4dpWpWR5vZ
2HjVAvCV/kahKoNeYKFU809kzOQ+SxlYHd1mlBocB3zmvQLmZ6nsjeHYUZc06+YDusaBTGwM9T3j
A6cjqTYeXBp70MsJpilRQMpQlUG8xnh/eUHQod5C+xFxcmSv3RUW+uRrmcXEyNclcmC1rlxh4Pis
BPnOeV5l2A1aoMeFv4Arihizvb6WwzNR++NUhO8uf34Ll4hb+qkrH3ziu3HM0gMA3/qd+Qdl39aS
KlPJaR3rclpPxcwL/HbPpw5dh0oiix6of0TCdNjqNBugwTummPq6EwwtiPDUcEG99UZ57ELSJTcB
MX29tHeEnpCg2ibwjlw46OnGYkE9UJJEsdfOBa/JgckVU00/RblTDlH8tHLsup5Dh2ahRk0ab50l
DT3GswyUJpZyy9egB/xL2SFWL6Uo2VBX39C3dQ9K5VeDft3V0D8/GKnoIQrpgGn0SDzRYRjZN74d
/j00srFWn5S+8nvbcnSXfsULBd0LKL8v1E3PvlP7RVV7RB+7koZnQC8VTkrIGoEf6sheaSGyoF/i
8mBmpQmNXLiyxNfXtV4YYKso/bBvu58kGglS09tIU6BGmnvdLEygLUHQGHldiu8cgTcI40MfRNlX
P/t9+Gj77pZ9plxlnUl1Y9Z+NmB2eySOibACmAWy73s6FG2l9o8LxywL00uKPrVFusr2SbsvWmze
HMHcyi6vRo576U4HfY1NgOMZ9qQkJ90FDgQwXl9okToRGktrLhLsZKPGOpFieg2rWZ96Uj4/bHFh
sXk0dGan5wMRnyumFvBocsoWEYU4O+NPRIzNay1LQKRmEfP15wdN36EYjD6Vl3iot7taYsp1hHpY
1rN4hZaJS/dBzOwXZ90gVFe2J71g2rpUgMv2B/wvvn1Psskobqvp3gxOf2/HTtRaGb9hiNOwKoia
108y2OJSdgFaF1kkaowMB47T0+Hi7IhsjROx89g3eraQeHu0eabHfM3ApC1SPP/Y14+MsHUZv2qL
Ele1LsEgqRjOEC2/+uhiEyuaRWOo0LcqblGdk5cnplX2fKNubVCOyYdVuGGMH50v+28ZWylzy4Tp
YvMDxMD82Tfu6vMIptoMS6y/5fWuQo4qM6Twuv6uTBxHYng6rMpJWy+5GlFyWJDqVJHT+kG/P2eQ
lIGPzghSYkMl+doTf4k99O+ldZHuLrTI5WxYsqq0San0JnmOLMY4xLGtAlN5lljeKlENaLiNRK2f
sFVa7O+XJ1i7KMBz3iRcdyGl/Bd8YYAt0Nyp8eQ2qFT2gc45f765JZHapMnTT8wb86HNX4o2Fa2X
FYCHRyfv7BV1DuZLdzqoZds3+OGmUNu9ceH8P7dvkWLeWnhBkQ83yV/0f9+IUiwGIRBz/U1wpTe0
BIAbejypk/bC4+0fphKpUFyd40hzXyEE1TziatIqZMMgo+6bzISuJcSM+qV4BI1DJFRta1/Hknke
8mDIfwV53dBYPiIEipe0p9mi+sIDcpwab6faEMI/gW1ND9nD0JqIbpC9QMutajt6c45wirhI58s+
wY3oSLG+DMiGYSXlV+Kgsj/syWMyWZy3TLzTcqxirQpzRNSmHE17vrR+NOqo75LsKoXENxCMvIcT
zYpGf2zLPZpexTHbSMHhkFOtb9ON/pKyvcKYwX2tcGANKzTBN+tswDQ/brq4yiBUpV4B6lAou6ww
aGpb6lMTrIYrCBbg/Fcp1jxdoH/SUoUrSt92ngQUdYtnGT0sOq177TgLBP0I7d421LRlAxLBMkTL
EmCjCZlMmPLhG1kwmhtJIcE2eREZnL8BX7rSNAMpeOWwh7tL7I0XPD7zpx5STxL8mCiPRb69Egu5
oYiMfdwuqsG3cJqoJb17F8c8TbAGyNUDlCiyWYXmekvmwUQ1IMV+6hNvdK55s+FD+jh5yWFUh0W6
TGyzlytWwFhdi+oYozuSlLj+QO7k+yXQcMjZ1CCDYMzA5lFNGdJS8BhfXBv3h5fVakrjc25YdhWO
3VCcO46SAAW1aLorKuIdioJNgm6GgkES+7sbS9ZypNNhT8Cxww1Mez7mAeJDXxaZqb1DtWhWasz2
xB4KSY5wVppWP3Ksocubz09pDDePjtSZoF9TRs8QfI3G/H6fgY8ol5FnTp4oRiMefX9vIDOTUZkg
/8KntwFbBREbzTYfY56NnVmIcmuwY9suu9LGxQPhrAFMKSUwFPHY/m38+CFs2OEtumgTzXqFFMhL
Fsfhx2gP7+PvUKPCYdK58PY55dQ9nfF71RQSha+SJXwZ4fURvRCAwttW4ns+xTzMMRxfSjNDMlkU
TzC9BdESN/4IkjwVH+UV8Ley/tXC5gukjaaTgTdw06YJFq1FSsAcgF3h04dV9zL8cNd2xERV44uh
F8LR32K8xjwa8nKRVhP3WIfXHqdsdvm6rQOJqlJKcFgMnAB6kM+7B4NQhtyOp2r7ivLzlwePusXT
cLQH499731hHR5uz9kcwb1z9afU+fkkjHJzXreO55GWJgA517yYgDcOCxPqtxtBbJOPKo7AjEWuK
eiBRr9gk9KlkkQ8PZcmtZt7UaEDls4ZgPCVDwOz5f2sm0C8mqQlfCzfiI0lHvvBIqWnYZBvB3E78
NDZYafD0Pc95J/zKzejH2OpP2DOk893OVMhwfPrhRQHV2CuFTYDOpVIdy1ltFUMPPND0/uX51qa9
pFGhnJIsnlAu87oOe0ebXbGtx6VBNr+PNYaxNuYqFX5eOPMJXBVHOhm7t3C6bsLiN5i1AOM6WUVI
BGs34h9P9d56FElHqNSnqFrgZFzynKSXPbMaLgpiJ8DZKNzmHZ+QdIhcQn3dqNSagljyxoF9MT4e
3L39JQ753iWmNUOXmnw3Gn/t21sz/cv3vS4lkEKm+yL/8ftPzXI6RRjtn4WWSktinjBEeFSBhTUH
NsT9cjoAXPKlwbjdfnmpFYPF0l6OEvlT2asudNYolWoPrzVERzxJioNVl92L4bresmK4Wb/hapli
6Ku3o+WGn1G4d0hysQWtWf7By9fVCIIWA9xazViUs0xZ7ldsiJLXHqhj1KYupFqPODues85bC28O
Nda1LGuArWd18b1VLT6/qlOkkH/vpzBoJeQQoD6bVzxZl/O0mG3WIlrVPRsE0taltBNxEa9C//jk
1vW+jLcljw3Crxz1Ao3Q23Dqtjvboj3U+JEu/M1THd7fVxzeVwFYljKU4xQyZWLiOtXISVor0/92
edFxQ0B57Up28t/0uqYngvcGQRLhLaSuqNNAmvd4ZuPv5a9tvTcbPMNuml876E/jM32A9KsLOqSF
W3kDmhw2C1QRdv/pnEdMktUajaxQ3UyPzajScMgxZXab7Su0GOn4CvzYT8uW2I2gfbhpPyrpS/1P
MEhcEObcGKUx3krma/6hTz2Vdwwada91wcfv7BghUD7cqPf9GSp9J60V9AU3YKrVla0wLElzzuDx
/MWHHtllyFVGlYiDR8sxQJl+UF9zyf4EkPNvsXOlKG5PLmNT9YKimgIKu6YiNIARY1aFtdgFWCO3
fG7RUh18OJle2MXtjNVf+aWuYF87/XhQ1OU8lcxjP1slWgq1rd3wwgGTfkfd6Kkj8r8YLjCq5/eu
61wdF46HCSmpmWikd1FTSumeU7SVcqYc7Ycw+Mj/fF1GfG6rHRbsUx8QmEdjQysP80nQBy6s9EEl
DDeeYljYAtvIdaUC2fJR/rweLHcCR4rmJKbAEL5wuYnA/Dt2JCKoreg2kU2y1se9grwRT/eisVD9
BWavm9Zu1c6dP5pc+oAyun9XTazLZIwjxft6PNjb466IULkVAeNErkuGEX+HobG/qglNcGDhEdtr
MudJ2m/dxCvyJE6NODDGZwQz+dw8TXD/V/n3wbqGS9F5A1nz35usMTYSrKEP1DUyYHf5MqoRwSMb
61yyfD1jznKl738d7zN2X1uKGXf27EjFFHHM54jlyyhD6ndw5cB/nNO+seGhEN7WjwGmkS8kfc1i
EjFk7rwgeHYRiJ2EvMRJsNBbepfUw65I5AbLQNexlf0FWRmIMa3tjh6IqOSMLx/3aZq0/fSobTMw
5tvEc+ns3nueTOPWzeReSpVPsLiA752GeUXkYx0cqnMWnXWI9SaYMojXdILsPjshsGszMfkpYx3R
AQeYqJm25Bp3uneliwq/EmvPN73ghxYcl9VdXncKtT3em0Ssq4RNIHMYc3YvOee4z5MA4HYNp3XD
cbGe5TTVJB/bIy/7p2nkkYALnlSI/oDdIZJb1uADkCO9it+cZYr33+78z4Qqv0plaZvQqm4TDb2V
RDRfcXRgi1FBuRJjkPztHu71l02t08g9snbUvWPIj4Skzikn/vTerMg/gD8HE5yjVo/+YhBqcz3p
y6sIWAb0ZStyzkYa2G6TqIC7p/j5szDsdyp7N6M3L+1vhJkw9hnjEcpfqv56SvFco5OyLQW7cpIf
rIjYCAhHtqL+D54+2e/S4JMnJ6gnuONJqiid/3uButbL2zJvKNxJsojV/Z6LDkxKhN18gzC18KUT
WsE4Im52u/xE5hQ2A7ZrRhHp7+rkixxwWQuhwkPPxXoadinNoqDykFqFWgpc+Q7WINYrKLKryp7R
GhyB5H9U79niJZuBCaA0ZawttWQ4Kil7z729cg4JPLEqE7t4L7khYul1l4I1vwnWIUPirT91uLL2
9JBwi4fHngNeSXka5w530jq+UTIE7J1XQXDviqHZz9GfybMrGK9j4nKfZDD817DrMX6tfxzacCMk
+79fDv0Wb3rV+rIRdMXlIk7SyevZhb0ewUCC6L/Xppb1SQi3qV8sYqmr5yWKjfopUg7AnGuJWWxD
KphwSwc92GG20sTecV6K8Y365p9EQzGcIT/xDFIGRRBlQcWtK1f9B6i68j8wdoXhxfQvs5djtP0C
dOwXarwECzI0YD1pMmQF72ihb9w7cNbiEmzPBHy+bbqFgYw9PiRvI5apuQhvva/Lo07oWvMqjUMe
8Mco3O672fd+t51BVqoaoV+I0QwD1+UZch9ZtaUN+6eiVgPfp05wc3BI2YXZfeOV8exOZwAsxgyD
7xF/SNTUkrXcEUW5KOP/JTBfrwz0phq4IYRi2hwGx9WoR5SZUlHt1MYchJbcO4DvbzL1yvHCQP38
P/r2NhSZsKV79jnZoBXVXT1aQMA8XKS725qrmAiZobyi9l9ML/xy8dOcu71U1BSv742gBDooxRey
y8jMMR6EpDQSkqlT4sSlj2aUg16M4Dljc9tSpJauqgXLniAvM5lTgoW/G5wkuYzuV0rybFLxHkkL
B/egUKM26scKhsbQcLYDPIP8S2KJbY6LDT95Zn8bbu/qsZ7BJEWUB+75lc9EOw557aqHIRt/iIw0
us4nJX/ZkXvB3I9GfxnwLd/lb0d2xvuhpE74SkVHtAmWHtnwfuiHpR0goq2PXe4ws+4HDMHkjw9V
zqjaApka4kOAl8Q1JG4BWtXVA0RH7LvpnNt8MnRFnLAE5BgCXYBvkswE/HYD+fF6wCBxdQGC13MY
LNAYvB8D6wxESQcP3AA0xMZDZqBBcQcj7ZvpFtkvD99+QQLdPkw04nkBYj640FtGryHJOB8YmWrR
Vbk4FJCgdaRWmxy2Z/SbKJGT7HTRNmFNzGH/bNvp97hASsEp6cTmWngK5bcYA/lU4swhO3ptdH7W
FTnjzeirUoH7bK+en8fJKDbZjcrntJ175u/MDnsGO3ogODGMlqGIHBeDhhH6SY5SbAs5CPgOe212
B+Noc0ntlONiApfyxLh/K2lhBLwMx73P5D+Ch4NpT/PH1wppJVEZkyECVqE03f0aQqnxDiWuDaHS
HnYElTbtNWtFp3HHeM9+YVIjvaBh9ZozRuiljLMSnREPbf2pUfD9va9vZSLQg/TuUtZyD+Y3x/XC
lkOaWI9/V0gdmSXHrXd/R9WYb3eWD7/eXqYemD2MghjIfPxbpdnvaLsify849Ct/gelqcPRW4DyM
KTOWJPJ/Vlsby4H2EZzahYIMXMq8XjjPpwy7S5PDagunYXLn2FVrwiPy1yL6fIlpDSDtfaYbyoOD
rptTvbU5m2ZK190Ig6uKsNOHpZ/ZHiBdCkV3HwqT0J0dCJ3Ey7r8xLkSAwdLTWrHaoja1BSIzrEo
1hZMAi7bAhxb1FtpNnf1zuXjD7fmaX+4Q7ayd30eMrpnvQ2f8eLVt1gDpJwfFk9qBAWur/N/0ESj
qZS0BJlHaXY3Y4y9hHuS55YYYpSBTzoBvS6J6jlP/5+Sw3JxI+98WYlY7NNCwwkaHIuJMay/b5A4
Yu8Pd6se3ssVTAfWq5XepSuqeecPlTePZq8tyTrGQnB5Dwlg+hNPLOf/9iSHftiYoUUn5pJ7L5E3
ZHyexxPQUAOj4aM9T4GrjdifOF4wbVJtrb32JJDlWTl/ZrE5c7BisKEgrJbCt2QeLCLKLrzbIJwL
oK75ZRQoerkbOHF3W2XVeELABUBvhZ1Qlwq44eW0I+7SZvBBTtCBxvL+f8rKcFma3XKnL06ik7TO
86rJGb4qfycaG8X489KhZMbPMH7qtwCZK31BSBT4yrYKnPJ3atgTzUOS9e+2xL4LNdwe1+LznfKs
tnubvvrrCXFSRWF9r8JKLuK2M44GtWM34vAmaiYPtd1jKGxyCYjDYDZroYdvDAw4J44OBECh4FIZ
PntknJWOQ12idSCeheqqQM4IE0DQtGPTiUktyDugnpWr39mQp1bki2CDKJwLTjStI1MfNOq58cpP
QDcR9XvWC/XfElprZP4lZ8JPbFSLTlFfy1TJ4qcvuAz8E55+thsfJ+mbGvQjp3Rto/RUM1KTsV50
jasTl8XET1qGYNDg9IX8ROmHISx1/IRCkfW0h09CHK+j/CxPMymHAmHSUYVUqJ7trdYwKzd8myX5
6y50gUwThXgtMsDH7ZsfvrIhtWCvuq6FJ+N2w5n6/X//HA09UyC1jQXsTOw7drIXeAMrQFKYQTTZ
u3Gkyd9B5sJLEk/66NraIqamY83mFzK+oJglvP5ePU5Z9gnG4xo0t2e+m/BOxJSHLt2oN+APEICG
JSTTlUNXTFv6oZtvDY54/7OtKYa42QxUKp2wIO+ddE4ZN9GhxbI6+c0eikiJ2Tszc2EY4uSlo8qa
2AfXsjwq827pupllJsOnA9ZneTebU/HLrqB2ngsFqzUct9jrb9V08gl4dRXjop+SrdvZr/Bi9F3n
H9tWCIesXmbHGZRXLspoiGsk7VuuplhGCghkqDZR42CuTdbbSEx7OA3WXMEh9+VFlpIpfeMDt1RX
c6pgMbOZg1rwKXn9Bc0bNkkEiF/hDip2wu++dHJOzZ8KJwc2tjKso2klKWguoRBqbfBz1+Ekvvs2
FJL4dR4V/VJlJ5JzD70wwudIKRDJN972vCyzugYlZCQegG2Xv+IGaAVmDLEoHxEtNCAi3dnsaJKm
FiVezl1QSJCFGDvAovi7pLIqAFTzfe6aSyzS7AqSZzErByS2gJ045NkLYUUg2MWrgP3b0KI6EThh
hk2z/PJ+tznsg/7Hs9Ni3Q1WP9nxL0G8OUqHsxZdrkjL70w5iWFevn0Y+a9ko847iC4zuHknjIfI
qaPGqTKbx728GJUTCBFjR/1B6VQ3x0ThRqYzU4RsEKwOqPlOPhcletax8ZZKmAdBzfJRgkD5lbz4
hyRpgOD5EvemUwShK0MLFaNIfoKwBGF7nluIvmmw1rtZDZKpj6E0djvBypz/4oB10ePnNVJFXN8Q
CSd8dM+eaywu4ednRSVGLvEvDXOkxqJ2FI2k2sJ2tIFaZrQPjT9s63EV738WjIPXz0am2qIGg6DY
XwhFKersa47Ujd++CblBCEkHa573sOfSrRxSypkFnoHVbGPsI2FcNP5Q6JLkZUzh/ridBlgUU5cK
Hr550VlkTHJQNhIZLcoAp4zAy8StcNPN2YBC/ljLdsKYt1OkiUJU7eduK08ojyLmGlykbEP7+Rtd
yv9x4j9HyDI4TuUZ5P0fu3CBtomeMw4SYIzxGPWhtSqdDXkI0LMb+rwsigJFKdSVCua4Gv5QiXMS
AeoZzaw+p9HM72+zf3LJokSD9h7KK9dieeXar1o3+XFxmvh8K4M6IScADyESEZ0EGEb0OMc/19Z8
UnYVJ2XbjWs5ExjIj2Cnn7HKQVu5FVXIGDA9i8ACJ7bJD3RgG5qHPFdeByKC6g6GSN35xlSEb+yr
UgMWsaDsj8jh7JuudQIJ62qn/512wJmd674bmlmbxvbcz1EpvAw0gVFmWGHOHbxQBLBl22J8p+9o
9fCVGHIRXH6js1igRIbhViwJhS9cY6GKnxVGWjAc9r6TlcSXEvrN0nbUniYx95EDTefTPdb70eGi
yUYayVoWCULDxfaqAMUJu79EdrWJ+VwyabpsHwt78kI3aJUpp+GopEbe8YJ6GLZOmN8MmLOw8YCS
K3YRqcmnvz6xBi0cPmOVKH2jLB2/WIp6nDYSM+NCar0T/8o0tSOWNjHx1AiDH40kTgzHJUlC4i0A
wGPgzuuhU8QIdtPznHpwZKPNpXzYM7v3+vCSrEBeE8f7mVqTdAhfgtJ1gBsgkH1bcQuTWh+IiSKD
L5qfykD2AeaHKoDjG6eoeHkiLcsqBUhEVdneqH+cfyf2Gn6iaxisJDosRAJPPyeMQzoHbHKszOjL
ukbS2AnCmHXVbH6vvMYbC9joxq6FP14qD/MSQ32U5GGBXvXLrakzXtWEsizwwv2mY7wFQDJWWEMJ
agsziQ6/CyFyOsU2rN79EU4mM61OCtfwEyb8z6MHVahlcI0Ffiy5tejM2ukSucKyfR+UvKUwFBXB
sF2Q4V3bK7DHzOZip/HAq46GUxJ3MdVjVGTj+JknkdGg3+tZtKtINbUIaNNp1OKGWW+tr4DZ/iJ2
ned8GGxXXVqGjZZDsBR2vGwSYO/Vd1gRtbQq/QO3ZfAmo3EMh2h/jciO+YyPc8L725wccBIYt/mI
90pj9MfQsLBG0+6M5+9DzuuLZ1BU3d0/nnKEcEwJCUIVgvsJLVIGQJon/B4lKfcjqf8XPD4EQb+m
KEPe0BEvWuXTpOjvPOK/+cHLiCsLtGHJn7nUCfvQjEQCI5gGaROWh2IxJhYLlL7bERG2lC3xbl+B
etuuYNg/muv9CCQQjINIKSvcyXkVZSaHyBlDvlx+zPZE6hKQtmZIUDOgaBbfngHqd44WzlM4jyqS
aT3lJUm/cZNm8YgKaFW5/dCLh6cP/ggR38p7cqAuJyvzNFlAQyWycR2PPp3eQiZ5oRKTU5pw+BNQ
jtgPqyWgYHDS8xSHs/1YWAfulu0ARGo0ZVXO/yZztAAz7A+AnTIaC0vVBE0na1+OMMWMyMQLfjpm
OTt/R7TejLht9pVkO8zBZYTVryOeoow+8yC1FLZeqS6GvIVIeCi6PGm6AF5H+ZvDhmlfNdGgU6kc
dgyCLsRqA5xashvTPaG2UlJu6+nZM7iW9O5jxtY48s070WNz4lyP6o46vEtsea9mMI1Bh5aQMPij
PnUhLm2fhlPrKqynLts4QiRrUvXJjA/656pYBkrhQxloqd0FNNx+AUu+PrLk1bsJbYqAvm2GJUbc
Hr6kM2jIDEq65V38SyZctspzaKs3VwLss2pM7z08xA2Tz78ixsMTA8Igq1fBLm29Po4jzlVLSC68
XDU2XtEwAbEIIoxAXKvBtkl7dIqdo2TvBpOSsTmzoAkfZCh5zoAZgGREW4e/TjUYJyg2YneC6seh
x0obUUFUblGL0VvsdEw8/4yfxdMYNCMdNF7nKVoAjsNgxUZQnlUOhK1PDRW0Okd7QV2GNH4SGMsi
vk6er7yrP2piOHpS1Zw+M98mbMVqyDe58HIFnMorqMF6loMwf4ypZAEGB/0jUltoI4ZGYHhiEWXC
pKNeJQH9AUROUDY5jcqOjOmfHvL7w/MJ9V+BZanu80lQJpwISjIgzeCrVsM/+hnTQdfyO03vi58J
18K5BmXsDMKi/1G5Fa2LZvKaMtv0mTe+JsPRaskwGLCawagSxPy4ZTqsSlalyqzaVHtK1tpa5rJm
XptxO7Lo7SMpT3HwXCaE2bgcXYCJYXGhgLQasHDkLK7brbACfTySwnulG4GMFGkUFXHr/Y3CGvU9
TagMm8Oh6V3QDFu7B55n2YV3omI171ojrBa5I7y6SBW8ZRFtBPJ2n4BQcEOIvGfkHr0vDHh2bYaU
1ttaf1f9uKmgPVv9oaLkIiYJbldqmLghnD6Ths0/t1pjE/9BKv+LRVPuJ8j6hQxSQsb6qbhYxit4
AI46/GIL7FYmubhtecvieaLEPKIo4NagdD/4U1JjLyi0XiS+ep2nk1tDX+ACSpMVkJLOahF2FPg7
YaVlD7ex3e9Tiqc7roJl0JjlqTSUPB1m006iw/xR3A7RWB0Vz0hOKbEl7otm0PZ9vPTORuMHcqL+
8YAy1TFrznTk0m/Sen8I4Ed/9ulM5/waaRPydcrgKBdakgo6gTZB8RnEhfx9Kv77ql60lRV7rV36
bvezsvS7eTpbdg+pXb/nBqtmA/5Ri8N9T33CDxu4k3HqfuPX18Dd+JE/z3DBFUjRy5dK5L5bsy/n
nrUaDMwVYiuACRpThjo4Q/WJQHABDpOi2m/4rtPGqOi3imFahk8stuM1zBRAqnWkEsZnp9sM68bX
IDjiP1+x20JgROQZcnnBc3gem2eS1uYaXTKXUDL2otMLbRB5F9GXOu/ADbJM59bUsNj4Mw+MmxVN
ddhXp0ALinXbxxxp9MGbKgy9q7TqDy9kQ5KoJd/lnmg46eSZTSxfRCL0xoJqZNbkPidsrPpglI1Y
4BEuPQ+3R6xF7YXP95aQ026bTwv1DYJLlNoRbjAMWplBqhEeEsH+uK5oC/7TK4TzGddRATzNMHY0
/Wqv3nXN5eFrnKYLDKOHUH8tsjD6yAQCUgyePZKNwN8a95X0chEBCAExlpqrvk30h3CulCnKT9Ha
oc/FhoQT0J2tXNxX3mFzkLs7BtpgGC4RVsOba1pcD+OSBoe4ye6+bVbbGkwd87/GvyG4iYmLRq2F
Xg8AaySdMtpGIBrikqN5o1EcdTe8w/Wsh9Cap+YmKunZjZV4pAb/dX4hKcfVkN2JblpNUj6Wwyh2
zeebCbKScMpEK3iYNsLXOONFFXVy1KKZ0LblC1f6QiWe3zOAsGT5yqo5HEaGHwF6AC4KOX66UL/B
aBnuvjjOQJb1ZAPTYgG8g/OOft4DFi8gRlMjxzsaToG7Bvl9kHWIFKYAdpnamvAUU2HAshrqr9ZA
3ViUDpOxrhbljk20W/Gm72D/1ruI6WrUmulwlFot/a4wdqpfEYdgYq8YSDL6nbqrFBdait19GMoV
ozYcxXqnYE33n0AM56L2w/NAk1pKc1IUM6xleo2pB2wYnRa9LWGN6ks7J1qLLrL4a8hCh3crcXXg
96ypWlRU1TCwRbBWt+9rFaEScuFfsbRBtiTBS/o1oXadTgJ/cZKYhduNxA84A+ViD+9k/SPDwT4d
Sb5uYds86IGHzRLM8UWTHZmIs6juIkf6MBzhLFI4qeogJeeAhoL79P+ypp6AlECwmlJnAJCktI4K
oPTeXtfz7bihbOWs1Zr6TfsUm4yVxh8ODJoTZT2hsRskiPIzlfkb7lpJ2NMcogzaX3FdSt2guGkr
I659zJQvtUCSFO+bcB5KdOkgZuN2HS3aaB4ZMbw+XjeJl5clTV5hY+XoV+wW8UO5NojJOrjEUYSk
IcbuItI4S0T6JNnPZEsiIXl2SH1FXr5yF87Dt2KY71CD32nkP5PF7d9ALaGqQUoCu58cfeQoyVvQ
U5Cm9B2m/LtJZP2eTs5k9ragnKYhWclF94a/EDZc5XF/c4+e3whmHCO6kiM4JgMUf+4s7V4TUjNy
atGRriceeWwQRUeFGYxGYm/vrKUz/GUjnuvEY+nda0+TIs6+BFsu3nWQfHkHZfyESbQBlVilgBQC
fOpKosTSHSl2ltjFfywCBVjJ5FAFGdOVUxNb2hEkpvJY2IiB7tVKAnIj6KRFowUx4n5odA5f4sze
0rEq/HQkE+UsMZD8qKTJNa3lJ26iFWrg/g3q+Mb5a9QRiAPgiqurKRi/JS8ZvwSOy9s3m6gVXs1Q
LHhog2IibkAbX463lXmTKu3QHZh/t7PbfnYu9zFm8LFAbesLVXJAvMLCWQWG53DOFAPrLsoyYvRQ
JbNZ7wsmsr95Q7INGo1ZiCkPD55z4sA4HhFXIjQsnOZFnhKkTQN7Si8sM7FVUG4FvEWjlWteIXmU
wejtIb5gKDpAIYLf3hH3N+QnPjMRHqbVEz3RzlsC8y/xRuZNaNlwmlKKG0SyUSl2Zqsd7ThdRiWc
0u8zNSnDjkSLiqWr/Sy7trixWGq9EbvHmBaQRQE6wQJyPhwKAK/E+Zo9RrxaqOGTUEglG46NA6WQ
p57w+7CCXUugEuTVKtAkSGQ8d5S6ObzEorH2nBTOMIAVr/Wg2IW3/4j/xxwa2Grbhi4VdQqPgJwj
MMAP4Hhw0ik3E7gF1XmMm+PBThHaY4WV4Sh2emahqbtegV8iJq+rWdUAFwpfuNfs+x0hki4IApif
7jotRZ50M0Hk2ijedYnKFqgKTvdvCUd9iP3P/2/bGbamiOyeEpjgYhqxnAFd/vAoWwYeXNIfkwJb
BsEdzxhNK6WTh0dvI7rJ3d5CjRCL6uHo2eT/LW073e1LRPmqTV5bUCUC6zoUjGLj0bJp3JSvzOnL
bbqIodxrwO8Jd4EI7r8y8tUF1v2tA7tteJILaxVUEf9r1U+Z5n/xfTb7ZnVSw077cZg2eSysyRqu
KRQmYx7lqhtxOYNlBhnIZTFN0VmLjsR2U5e7cVYVCkCKdyfzZiv1yxgKPahnfCukqtSw4t0f3gMd
uhR6RrfPMhSkRBvyeZk2Z83JTGc6vO8/uX+B53+o5x87adAzywAYnk/gE4yYE7GwqVj60D+/Ua9L
JsE9hBSE9f6krrcBX/vn+VPXEBcUXaxDMNUTHkQabXUSMBz2UTRMbY9alJpwJCcW4Jz+9aU0IeEF
OyRnTfxgVsnV84UBNAzmQ44y+jaPulUaD7UKZG9MacFm9r3rm06efHXffSrJe/UAQOOIVwhz1xGB
RaSFd0rM1aX1rqo0URUAwU5vIzDC7sxs8u0KpbXqIuWHabkfZ4s81tvT89xuUhT8jyJNvYzmIM0z
E5FY9oa2OPMAqyuCoCImUOyoVtpHXRUPd00uvQ5XwSaHhQM//JhHWS/2kStq/TmCCRHdu9WLK3B9
WXxZfx72HWWyPEqIRjoga7A6/8XHsufSp3RM+5R5igR3CXTPwhFZvQz/EJiEbH3XYiJmC97M0grL
bLaWRtcPii3zTcAYyPvpxiiMllfLC/Oabc4RM0kn5JLsfEjaAsjlpzMjrn/twmgLbutimzmhCneT
EcUvbvC8SZerNGOWx/rLccMqha9ki6WORCOE/96WYwnDOEaA4hErqnJRNN6gelPWPW1h6OLCQA98
Tvk1kMEH/HKoVsohtu0ahkqWgDVX6ntsYkPxkS7Amwb/ulH1QN0VrfNDObKwfI0UHpC0lUdRbNmY
3mRVMFGfQ/ed9IV2OpW/PgMr3tTEzdgqqEPzaF3RLDOLPy6ZBYKZlzIjWkwyVuINRdb3FYfjVu7I
NvYxWC7DkUh0OR9A4NvrukVAYX5lb/R3iOMU0vwtD7K/BG3p+y68GxgCYp/esCf1UCmJo7Q1848m
8Xfyt/dXpROkhIRXBHiEYjUkvJruQBVSk8VY1mep4//cgSRJmi269pFcqMVtkU3wwqr965eMsKi9
+wqV73E6FGSPspKuyt8g81qP+EJx2Fv+EkHQk2wj3FeTNHcBM1ILOpJkWtFR/oroJuFiQ8d7YJtc
B71IPju1UpvfZVbyhhdtVAdNf0G9clIsJKJEL5eBM3VBpqSFOGsS2Za5bFJZGQMs4e/GkYHFNtwH
CLymQXNwmzGyDpHoorCNZirMJ8rw9P1Fk6w23c/u2OvaKbjvpI7t2ah/7FGSSHuZ8K+AR4wsRE+k
sPAHQ91aK1+QueYo4HQFd3xSQm1lRoPJD3L/62KoeSMqrMeSUw2h1VgHPG2cqWh7RojVJGvev1XZ
7cc1ipv8kNxTOoNuQ+59X9khCeoQYYwTjT9MrpDaJxc5sCD451b/ubqADkNSpQm79Z7GtT6dZxrz
02uj2+Jb8jJotwjmmvODToUGEiMMBVJOi/c93rZ0qxVyRwrbRoH/0XUZLs91dJWoRAtwdWxFAppS
0r2nm4vWDd5ohNAxs5f1hxjZXrsPASgqQ0v41O3Unfr8I9nzpfT1q0CcwWHTJnINNwpDMzwa8yDV
dUrPOEadVtQtGsLkPRMlL1/x9bK1qE+Sn+aqquTVRe9u0oZU4mbrxQkMxkvJaTzNxTCo2G4ocYiC
53WwXo+aFR+GvjEmhW/hFHy3PnKNjKy7AA/AG5hU366qvja6cQqkCNo6W4CDZYCfZYWiv4Nqcw6h
md3kGAgNC3VpYYfsZWz/+dUcgIV3bIB9GZonvRrwjOz3XTFFN7ApkvSlrTNSVrbANuP3oCw37aRb
pzCbHOb2BsUQ27Z5u3oKmwua9EAUiJW6gn6mSZDue+dUD/nW5ELYL4/TlXLGYCfNrbsav050DnOH
joYiq7kX3enkCaow/X5W5b0c6SRxMxVpU2xf2gTmuyUl+llAWVxwi/AzjrF6IvEqIcJBtZDW3ZhP
6DA1rylOzTIAUGFTGoK1sdwaiMYie2J0HbFHRhE8g2+DWtMlZa8jOPiE7b7lGHFMP26dfQnwqfAE
xRJuLKkv8QAJmRGLeW+/CqN5Gs6bdmCRe7QkCQWCGFKIywxaTa3iWuPhtyBQqCpTfVJ3vy9HVQqi
xOk9EMZTKr93FAQv8a0nmbOWJpv2FCxah9GCkPX8Pvst0h5U181FKRzc6XKc29PHBkQ6065TvVlW
Q6SvPR2I1c4sKzLH8UFWBuReWCYsvahZoZM3allM8KTOysW6DgQKjYCSlzDvDkffpd3f9cIIibj/
oIuGKPC41uSbULI+dXi5L8PZasmndsW1Ixu+TVYMHawR1HXn8im2oVeQVqvfVDWSZ+x1+9NwGp2Y
04mDGveaJ01dvCu52F+tLpwY8Vd5X2Ve+jJkTd9xEZLRIEP5gfwJf58s9toXGW4zBJu3fGrarVDy
2NDErolTRJJLkb5ghSBzLhzyEB2otC51UABvCD3I5biyon94U1Mo3E2p19WV2l/VTq22V6TJqhIA
SilcP+uZgfZdZYV3y6n+cHt6oB63I1kjn5JPkSvgPVS75SBvGFLFadUpIs4uCD+1KH8cN/Lmhdrg
oJjN3TgEBeN3DQFmXdUYT3nfxE0s2+taXCHaQHbOvz1fN/I3kMr3coj8JmaXNtwEMr0kF3T3W9bH
Xtslz7WNBwFhjfNzpYTfFPwxxMmaXYlr/n1IHB2A3i6Vq6EptQw7rLUSyjhQC2kRybwEuQXOAt47
aui5u3XDhQQ52GdQ6+UN4DybS1SYD5XScukOHdtTWp1+Woh8B0zbqvszXuswigeheE9+xLzxxNVX
PMlup+0tMXbIBcONMZDuEPosGrbakT+DUihjawC4+N7N2OPPxjPHq/iI44sqd8S4mgO5UmZ3aRyR
qEYYDH1fAIjX297FV2g1nZWAAGfKR8N3QXKrUdAMR4pBpfsLedTUI3euSpCWnZys+59txLKsRZQt
XhqPUBtwcT205nVtZFNJ11iJGCRwkVPKuASiz1eSRwp/+H6Emib4JCg8RS7wysKJl1yt7CFUCp/Z
twYnG+0VMQFg13/HFMnXMneyKBgAFzI+XxP6D2T+GGAl7m+4stEh10F3zeofaAWX11TwQoE+s2AR
xXrHgQfj7GU/+R4OgGuZB/kVSxQrty4bFXPfd4sBuxLFcZzs1Z74grMJPT9b08zkcVrpqIYSS0Yr
2/ZXdhWLpvlaG2AyrdMZz/zE1RQsHH6CrGol3/69AdHzJKeDuMBokHObOby5TDL6Ak2GZxNsnpAQ
VpsYjYPKD8HiVico1/Fp3eSrP2Fz0NETzzi/2gF60/mss+qoTiLgYQJO9KpcML55HfwFesd6YWbO
twqL4u8OIuvNYVNSUAIB/F/+Mfc6z/JIQsbgSRPrI8Snb+vvKVyG+5Us4sDtY0MuR5b8jvljBHx6
ayxN1KyLauy7YXeRN5jpoWhPf7I+vQqpF4VyE3IP4CYHl8RmDJ59rqishdEEDtHAaMr3fItcjsC1
PGgc3vreHHeUk+0zeuqQpY2mK3h6m6hL85t3P+/qTs4u8dL3EUX6Uf6JKVWx31P4ZE/ocSNrpyhY
g4tWNNHuvtF52EZ1d2IGrumULJ3QZuD5vgPMfgtPqzBruBsp3SfCERN5zEWbiidY/lX/WDsgZqgC
kohBVkVrZFY0uWSrmdBSDJ45fq06PnRhg4NxoMUEvcGZrHp2LcwJ9K5Ls4sfvSYOnXjDYO73puXq
BaIOmGIup1Dcak1JrJeK/waoKbJmA8z1MF266XVrCZe4IpV0zM6tPPOYMuN6wFEM0+nxuTBLqmZo
k2BFO7TSroznvjNnOG9VJUyytBDuRTT6of8v31aKxBdk0teuLCiIgjicyhiCCQJf2cU2Fgqe4mVG
iUgFfIPVim+Pw27rEqgQmkGVfJHKD2JNkscHoTk7fNbtjWK1CspI2AdyBeqRyfYkJCvI/E54ZEZe
twatGmHugruSOLh9gE39CLuL765l+0O5U6x4zLDWWXp9mNRHkzj+sa0wml4EWNvTgkQ7aBE8leDD
hA4C0KxxtYObNY+E2WD2B6mafIvkE8cOEnptDK9a7q/amPgRCehvdVf929wpBLLKQ+D/S6Qg4mud
7Z0gSHrPXGbGiyUK4BZHvUSjyRhwrHBWgZIE9C/p6rOyrjifhAogxCbtNhNGa1aTo9NfpxA+T6gw
jYad974GD1t5jrEfLul6PVE61Em9WvHj+03wjBGTtSuxtxfuW7H3++53zMz0EquAvap1nOeKFhAg
j9wC2WNNs0yKHOnI1nrWXgiPseNwg5j0pOtNXZGoeHe3HAOrwuj/YcsClx0mtN0ONj87MzQSFMwH
iAGsVRfM9M/Ir0k876YrLtD5vGoOTvqDqzYN+tPoMsWXGsA6dZn4D1+r0E7i4sYj9qOqWKXXlgR+
QtQvPNgd+pbEvzYeLGMcEetjNsVNCQ1ND4vJjWWFot5RdJY8QSSN6voOzN3JzhulotOtULUb1sUw
n15fK8SI5dNaxe7ZhHdTVj89rKK1973uHwUbCXImtdHfFT7v/m+ovx1gvshLef3hWyhD72XinRjG
394E3ifgvD8auwYCiMdhJPvuenfM3AWxHx/3EoYR1s+y92zovVfIVt/7FQeTIKJ2YIIMVekxwnhK
QkzKkwqDuFFy46OnO5MuAGFjBwVAKa+kt61ns/6LxS8qj9LbwUsGHsTwpkM63lM7PgpYDS2j/D5f
kg08JICOZ4sFHQV8CzGtaciTOHD2XhCqa1cp50tANFFtSsdMTLSsglKJNOsB42XEld497i3MFRRm
xLyyptuSboNs59RHHnaFDSCImxcFQZnEMoj0pv4aNpRxvVj4fqEp/nSq2qU66atmjxW8Dv/WFMxL
yG6gGQDOl1j5h+tQeZY83jEJwCDlSMZStMnVwfNwV1qVQst+7x8rjQ53BeezLYJpYpV6S/K0PPfK
GVmeaTxc4GJVaWQ6mrZSrSkpKyfgRzS1079U6ICFcW/BHHwM2oHcijEon09EapXU6u7dc0xP1nBa
JVoMLs0gzieDwULE9FHtYPOXW9l0z95GesVFGzjMOHX3Cxp11cQGu7Y9MHl7z6Wpljp7XdaruVY6
+QFXKsD1/tQAeQyjWI945imQGpOE/VYM5rkURaHgz3aczDkCpR7is93fOiGrTt7gDMPeqGDd9rtA
UodS/O8WgloR/1eDpUeKbw1GlCeTBbGv2/QU+0BZ9btdoohev34VjEa3eYegVA44eJ47DiAuk4VU
1e0pdzFzqzoBJUY0lRh6jC1vj+mwZeCDQHBdbVExLe6o8eLt5mg3xvmUnX7NGIB06qYs5Q1FvXfI
lQO9hEzv2JLskAsrGVIkDEFVclmpAMuNUQtCbplQHXfdl54zLLd7EWhAMiP+B6SqtA2sdwETLSw2
1PQO28/a0RC59OxI+UoekWNVKDKhM5QRy4lHf98dBhXX3/OrDFcJDHbFy4eHjzfmbTvDw+LREt/3
G80YniHc+YgPKrnAMq/hqgw852k8vjiadluRgXM0IfsfkKPtmlY/B3I10lWzy1b1ZLtR3RYLrVDz
TyFvvPrJaqjgGc+zQVgpwYWq2Fr3h2UUGBhXgaFzbehrzryzG88+n+RKqa4w1U/Wb6lG0DhVJNKr
HDYMjXPI2fZy+pnwjnlE/nXhsqmosfuXBhEmEb3uNRerflDp4Vddk3CUILi9sUSafkR/JlT5Kldg
/+i4feynjxYO2bI3nnAeLZHjOXXeSpuW7663JCWmxUX1No7CPhksZWrWJmQ4sGYBj7ei0LrqNMLF
v3fTZGxgHYD+ZzSetdNJceWgWV1GjKYOF5Shd9sKZe2gU4LkpRj7xPywCKZ1NqO+PQNb+OqKHEpK
GzFU5eCw7Vs7gUdncmTLW+DcA6Dt95gZixAvAbtvAyS/P0MmDQ6bxtUBNDvAr6ZeQTdlZ1o24RPH
vI2oz7SjklOMe2Do972u1JHP3cU2SgDXZvVCK4RdmVvwsz6xT5zItLHuapDWVhaYjutTgcLG+ciw
xaEqUSDZbFd+ZNY3Kdd0yTTezuJrhmixdVNZ8K1SFb4u8ZBq+jx/vnAqz+NXtCXnzH9AtMbvnXt3
trAVBpwckbh5iAHFqmd5mHfkdnTGcsW+m9ArChdSnQeaGi6IMwD6rx/4Qw6iN77AJn9apPTyBLSP
EJB2jJWqGNnFhAyLny/sqGceWrq70Q5z+5h8I4I2qDaCe9MD1c6/rj4cjkgZg60NL1esXorwVxFA
B6Mi91RrcQLg7pt3M2/Odi63kPQv4s28qXJ4VWCIjOiXqwyUg1VU8mvCswAEj/DUBOZ0csqjdkxW
VnHCd9f8jbGUorreFESA83xf3+DeO067EhYPmptgFIoUAdTiWaYeHTepnRG4AtKmHetYr8MnfToi
CmxFKbPnxP0ykOQ12uAv4ZTKZo0diJCrO+/IEaOnu8IMHFH9GeQJA35vQ2neENze11apn/0rye5b
4yY9jkYWJr+bPPqgb+V0lF6JhxqtWBKBKPrI4Pnp131hrxsWKLMnbLNsa195bWFok4YejsBWJwXD
W3wysNpF4JlVpjvoYt2Vb2eMcPAmJ4TNgkAA2ik4B3YFsnyjT4fxknp3/Sz63o6XvIb8bgMlXvBV
JIttPeUejw2W+i+AV/q6Kni9MTWWtHjVkHUxW9Hx6YbvUwTbWuHsWrhWwFVjSXATPvjmzfTWVta5
gY0wFoclDpmTfa0s7WdXnMYg0K0j8puPK7KZH26Oal38aBNCSC+kFYaf4vPEuKUqkxcokyGHB329
SPI8chPbrRU/Yu1yvNZNSeVOae7X5EatERhJ/KwhZocJpIjOdtujMG0XCDzrheCRx+kMzcyxItZn
vpIVXsmH2IunSWPOtnL9jIuZvpj2hlQ5cqubr2rPtuVJ035VgD6BJBSCOQI0SRoSTR3bYfom5lZf
N53DlwwK+hNPfcPOv6kQCHaO2al81uJt5CF90VXlNK8ls8Ih+gNrLIIWDB4ZAbL37Q863f2jZqn9
w+EknPNLVeAQPl5F558wXNTLhAPbJ+xhia7vPWXWHBLZytRwj8RNedkNWKswAs+afDLN6FfoVI/n
CZU2Vdcdg0lTastoTa2eFA76YFjKy/9Kjz9XiH+O3vmDcOhUcqP37ECa+sDZU2hNlUlh+p8rap6m
0Z8SpisXu7oJLedlHlSOYwp+kjYZPHkEsod1/T09J5rwNRRJg/MQ8P//MhCnM9aqhlFjCnOOqImg
1MCg4ZmsxcScShZIuNGjE5Vrqny9YuJSmWmjj7YmvF9vHHjphvSziBHy91QeiMF3cntpvKuZNnIP
wMTxFJASN+B3asJitPbiGNPBLqkNlA3vF7Z8fHAUQ8rORhX9ZVfXFVOkSUSc8PCA19WivkPRMlBC
qyqxX9Aqcbb72qZXdNwjhrKbTzbt/4FlxcEa16OrJfSAoZHk+MQ0Gt/gdYR4qNRAKOxW13KdcNdp
MUkDXLB80Cxp6uNjXH8XVEQ32XLVrx9Om1mS8mIUYHRnOfp5TbliU5XIf/43kgsxgsqDtVXQpsEL
+72pFa8IKKmlAEt0nG8cbT7cqCUD8T7S9dJklPqhdS3YNWZTalVY6FMRbJ2ZCY1+ASR3Ryw7SfnN
BdEYssZ8mn/DPYeV5fZfZlOTZfnBIMEKUDzqMzCU35y3sityVKvw5XK79NWTK78FwaGhqrD5xC0e
Ohn+T76ImsfwcV71D4XcrQMyyHvFSDXWEAK6yPq7EIjcrEMoPBh+BT/EAJTOsHEfwppcwc2YbYwx
jsAnxcrOjYFanNqV9am+c7tREwB/ScqO8YBFU7k3Tc/qV8ovqfxxd8YSgBEkzQhGbG3SuoYtVtQi
DzqYhaGhxFzPhuXw1jEpzOe6b+1YCLrjqNfmL7uwW6z87c2QNkhlYQC3Pb1trSgDmTPuqYLBxne3
BfHu9BfD0XMYCgcPLyYM0mRIc/uHYomSBITA58LHTqIK0lDPzLQ412OhUYhlbCypFQXQOBuEWDDb
TqMg16EK6KC/6bH6RxH7tm6/TKvRqcLD60hOA254k33M1o2sTfmm9ahiW/epEO+eGeomRSEU329c
8w9ATYr5L5kZ21YUmdqNp4IsQvBhc5jI5wsWiUclyAduAiFb1V6So5raOmC9dhmiNQKIlDqTQHWN
lXimjAa3BUaVl5jFP+GpRPjwZKuY0e1THO45r1Fqt0g+p+uL3IL9gu1pZaTf2NjWCSrrQCGwBrON
pt9+dUSR4RP1M7N1F8KH3QQg9XY3vPFOgXqW5KSYDZc4JFqyYxKey1OUt44Onjw9p5aXz8Yes7WZ
fPNxeTA9OtlbyF2MCPZWKFOocz5lmwPPkiYNsuqqUv3Adk/+5cr4xKLjcLK6cLL0D0gzIWS8qQa9
lnNffqxe0c0DtrAwB4/u3coYo2tVgSgw4M9g+ti9VoWgd8y7R7WU9EFQcDrPvLAJ15g+ORa9WN/Q
0ItHal2U0yeMtPX2vHzdhI6abGvSPL36spYAgaZdeArL/N8FTd5R3tiBT/CxFYp+HmgBab61ty2v
xCUWMEqxPErKHJuL/96CmNqOZ6QdihXo4I4y9mP0utnK+N2Ed0iG9NC8pDx2SLddHZOpJhxsVwH5
SzS4Q0dipw1UDoYuLadg/YL2fOf4ooR2uuNpRFd1X6TFT2BNA3znKcgTW28APoQAeH6kXEZNujKY
goKAfraS/q0m+dGYmhSWAYfAMuRnHOJRspXPexMZlbT1Xd36Q6g4/udu1waY9iPLCmc932rwFhxG
/z+OhnUBmG84nZmoyQtJSQMkzHScupcZ5UNVY5GN1uh/D+BX5rU4bvs7wZs79V6Iu+BdO8AgV/yy
9+0tkJ/ZJOmHNEbNagHCt8SeJKpGS9NBRW/+4GlEVHqyxqRTCDXtY2vic4E4oFUgVL2hcJy7qyRk
bAbUcVEArgWSgwnOgM8c7Z0NR+ZylssRJOj3tBhzRC2vQ23dyTIOBqSvMhnv7fNyRoptNSSDuqY/
k8ayabq8qDEpPcmzpEy8iObbRhry+LRtHzHE0YKCazIjffI4pfFilcwfQzk6q1+2uxkBpVD49qjs
wj6/d0l5JHHwFof8JIJubdQemZRv19EKLdYXAPgBYfG+SxBgSaOM//BbB5H9zCLPK3GAXFl8Vaxu
QvZeeZYc6VJxZPTEgweTBps8Bf2UzHobX2XZ0WwazSBeOu4sLyX1sDXt/1cpP+Qc9jQ1j/8PFr2V
R+KfxHS6PcnSt85sixSW53RJDav6u3RBzeIG70pz3KGhlR6MSWSUncHzoHDBGMJROBe8fWB6tQ6D
4Im2xoPlnLdnBBjh2gO2A+kcDpe/g9m83D0KOiyBybdQ4FoiExmw3oDy0sBVKMLPiU2015rQase5
qVT93EKbYqa1WNXCdZIpioCS8l64J1asdSexKZ70ayNF0hnObQunpxodGg+CCFtI4Sd2OPbzK9tH
cijH+6mMtXSuBUhjtm3c8bF7qqJKN55jKw5zm2u+NmcGzg6rOHRHR3HetuYTBL4RTMpHGebZhBLS
IJXFJk+gfhgnD/fxdBrIaEwQtv6HzBCoCLf1NH1WzQMvxqXErrw0/RKcgd/UuxKwYi1uXQWiCa2y
4Ah6XzGVUYvaM84djIxlnUU3gDCXhF+7d+TpW7BPmv8EvYdhlCRHJyXxXZrwU1bc9tlk3AShXT8j
W6joWiuos8uB0Xkxh8JWjVnoJFz9gJAJL/j2ovi0GG2WkM2fuxt0D3DNBHEM7Y4hViFu9PvrxGGH
ez8xdcsJ4ctTFnF+wPVsWjoaPdLulhoy16HVWd1tLM5w5UugDh6zKGqSygwRKZtdj8b2wHc2kfTl
neeQitJAVWzHQ8BSbLRrGESoYKtEPD4D10KEZRq3lGHNw4v53FaO0nh2T9YiTAY93HvE65dLz7xy
uqEHziZeTPAeLTGWkMH42iAUrCw0Gycj5SJIyV1GzPcY+MtV9grARnG12qPmsPVF+cHNUFn5WD1S
0k5EmTkOw7RtjNeb7lGdR3ZRSmKLu9axmfP1/j7rnzVkkw4dCn+VEis1jsrFzu9Ln9w7rrqevCHO
qwBACuFsbt2l9yytp4Mj2YuvPdjdfYrCwCQbuSWsF94gpkwD0AW6HzFPl0zPl8jRgsDDrJjZbixr
TodADsLJfipFxrjS1naUwSbrbVoUSfXPNanEpMmmhAOwah3CWHXgz+v7fHmBuudwvHX1Fy1LAvBT
iBacoh1MW80hDanQ5lWhTYYVFBEJj0Qu9t++tErAzEvjMhgLE2ju75Cf406LGqzz6+TuGzgr5E9d
A66yueRu9pFM7lmAJaBze74TgDVc7687ygtQ4rGfPgz5sS1cu47dtMHADW9oZbzzMP+vvajcPEFg
r5L7adelNPzV/2VweZQGh1130Q56lBzYdf/j81GLxJk1uvB9+ixnMO3xELHETa0S+rAaoediWsxu
dErWO7xYJ9/8lcC4ssaOog7g7ujjuNuT9QWCOdniuEHN2Yo7BA2+KUUQayDh49F4sYSkxFwY3k6A
nwhebb74hIak2//dt1g06p5p7qFNMHeE+UFQDN8HDQ/suokElBVJ+UvSwLFAGSKBGPKP/cU7yw/C
ovYFt14wTpQUq5RXhS+Eg0JglAc26kKmvQUh0oQt/jv9ZIuXNJwBYBcYueSQXKwfk6YSuFdIgQxN
XcSGoZ6LUrpNsNSUd/+IyYiL5Rc0zyG5YPoGUBOJPtfmMEtJFzVQoD1IME3fkfvmbvlWk5bTe53m
zW8q/UAO/Lsqs2A615TP4qrPPVOmIrL7qOqemCridnC1+5v67PRWzVLCpggZUsAe7JIQubjwOomX
N6s/SsSzsGF0GvB5taiBkENm4Qfe18X/Zm6CLNIsn6nkuBNAvi0pqltMLXM1R2NEXESGw4lc7k5f
WZdE5IoOmzjDsUT3Ey1HKQDsdUDTO8SNP89ncJ/CQV/BrJdLdeWPTSAP2kqPjdKP11yVsu04u/BY
mybAUgiainblGp9fj9WKD7TjpsyNx61Bo/dZe1Kqh7/xdwbpH1aDCXUVlnKR8od3NX3dzV5d9MS2
/IxYZoMEcPhPbbjJGl+EIRQJ9Kz8bTSGX3NOW2cC5AAb/o4kirAxZUZRLPIEfhPZVFsdnkxaQTkK
OIwkClaPXDmesaDxRHvk2YlZreDm5p1fQJEaPgDD0JL2NXDFAdzp+g/Acn2xqBoX1dfSuHCxURHg
Z131OgfyWgaur4LyaGi0+KYiz0ujionX/JtI33BCAn4Pg0cGSyACVgL6m5NmRS4deG205j7NXskr
2AhGRrFSuz2NEEZMG79kxeRhBb5U6iB7RxaAwVtUapJ11VbdQUmzw4aw7dh8HhkdRIu9GXeoWW3Y
gxPv32EABY0+nK/Xp2RYf5a9uikKVA/jBCVn+uSSjn7Z1rFoQi5TLT+H5HfivsUuhsVpB3qOX0+Q
U1yLIkkK1NwgXUXJ9nAviEw88816Y0gCxkFJnmn1EYmfbQPvH+FpYMHIsJXhH5Aclnr2zB0RrMHJ
9QejPlJmrCvxFcC0JO9PDPCR0ZmPhsc7v1h+wuwigeCxBgNIVSlmZdHmoOlQltF1wJ7sR/atYo6w
MqAgeudULN/0K3yk0YbO0tY4o7RW0fFbewxjddRqJ+tka5wLpOfaqdrNLz7Vpn2VDpg/vvwV7kyC
ikrNY1xTJUuMmk2evx6C4Jmyv5SgP2icUODVCPhFR6qffnCddIpHdWUBqCOglJr2x+MN1hfZ5UP1
JNa7Hktig97sjWXNTpIwWQ1Hh4dUn+LwLIcyYdRpQJTSoYEUfphig9vAsvI8/yNi0C7LsK7HGW28
SyNQwWkm7DiEsXfdDXbgl87fI6SCpC2cWT4dF6SS5heV37fLNX2Qj6rxWpx7GH/R9vvd6V9cpNnK
5i08SVh4W85mus5d78zp8Q6Y+P7CE63Zk1+g9GDpSZ4DPvqY1ybhx5Dw73NlTfShDpWO98TsBXJq
+oDLjZ/hHjp+6jqH73iLwrYLba4dTUMEnx3pV/5QcFsstPYawExNYDPY4KSF+3GdXz6kwASA85HF
iKDcagszKo0JqWHROBVPXBR2tgOhXMFL6425hqbKPzm8jWtHWUSAa0/qWCdCANpfP17hZbo87AKq
gr5PF86nnFB0xFXgwgQExuMBVX1LXchM6mEdU8sGpA10fbizv89gkZqNrSHvH0r10AKz6cUxXIqS
JLlzwohTLZ9twwbpfZMWV9o8Uzb385tWZyRRiDyXi2QkjZx9jYOPM72eKGQ7iJ8H1Ay77kEDHB2u
hu2u0ZzwbFycPraVOWgar5vNo19f6tBTtJzOJ4FCX6qhuwAJVMQtZMHFgGkNoajPqf3yq9I/5A6d
4zst7Q1wzVds6Bo8jtNeHcTdbTHocRbiSDz9tA2eDbGEIaAgp5ZmKFQ+mWwW+OksayDR0v5z1KLq
jizc7+4yTNvKcxrzHVqMRnBBpa73lUm7u8inPW8iUmqim7XE8H8GU2GfqCOtDScHPACO9B7breaj
aR4R5Gdyn+OSDlAwB/mMm79HSzIG498FdOne53v9YJG/DlAGfTTtrBXyvqVBa+KM8yxHA9VUVzCb
ifqVBt1e8q5eHbrXuziWser98Y7AziB0wyI3kGcn1SyGmOFrvPtAlejkrVnkaK4A2azEEsEpW200
BulnwoUP0Fi/E4Jbfc89Q/JEKFLEF+OXs8hAFJ95CWuTzjrVLNtAcC5X3+whvd5VTpe0cQkOY/sE
f8kqcMscRalg6sha9OexzIrBWUkP6dEC9bBzFgGIWRZj6O5qBAUYThrPYGieHe9huTIEahiBqB6s
3kgJ7UQqCMfPEf6myFA0/qQlq/Y3+5j9eOH7cLUBxwYEdIKzR5MflRGPzEn4/rbgvqEOqTb/MmIv
Uwuu5WhXcZtICrytH75tqtmh9PmS4TeCqgxOQi23USgU51ajcTsTN6P6vuBzMzp0WZ4DhGWI1CtR
RejsxarZI4phvtTthmLL03tjqMTtoQV6U6ZsG5p0f7h9PCjG6iip44uTt3OtAMYwXHqOIOhWH4V3
o9FTgrQO8JjyTM0LpjGud0LzKljCyAscycX3DzmJAKxpFwrWbUTo0dF60L2xpqFMTw0TFBPRDERO
fej5FdPK1yKGNUBdrLU58UpHgue3IXI9a8TGzQXnXZdAUkRQFqmQLh1NIqv17sjTi6zjYi3Yj2BL
AjyAmSHhoLrT3wQP+vtsDFmBBm/wzeQGSBd+8RyAVB7w3Evz+C43sOTsEp0RDkNvLDM7jDoIdT3i
pMx4UOSyW3Q7DbqwQrN9E+umGJ8R3lsfgHuo4oJr+1x1xOlTIic48bhemrdfGWKGpPvMIYqSMAzU
hr1Umlsr9TISYwNdND+0k3lfdkagCsHlAJZMOAjkzHRrAEujMzpHijWvcOvmtgZ+dHFoG/BJeyio
XrTqqLf4CNLr6+/jRe3SLarVL+Nxg1iZ70V/jZUxK8pkFvBzKnQUIYyUOt0/VL5sUXGt0VZgri+f
rQkrRGIcxmWNKmuOgGwc3HhTf7/2ygcF/WGm4MZ5KGe0PXbKUkErCObF2XsD/2FizMjY4g1O8bsq
nH+d+qfsnv/l90rpVN+77w1V04iIk/upO/Ee7gaX8xpj4X+89HrCrG8DsCR9Luopu0PhOXhI93fn
9pxYZoiWUo63qJu2CAdQHBQ5vJz2uEacEcJ1kXz8w1NGpGYZ2IXPSrk7PVjkMXYkHoPP+rLW1uOK
4UHqvD68KOhy7p/MDukLmeLyPnKTfk8hE3hGVfrExgFWZpiFVHBnV5kkMbd+h6zlwWA3zYVzx3p+
471SuDpzsCRkcgUOSJqe7khnZZ/cbSwQFEGe1Iuk01QarLsnV4idduSTVRhRuVhz9aL2zuhCw5lN
A2u8TZgBMuMniF3TETFy6CleKokcirhjZ+tpmlixThX1hbAqi4/xwlXk83a/ZkdmC4rXxW2SHUf7
lNG/sQV+WIiEKzfQy9/T2yQpvDu/GTF5qf+2rqnBJ0KyNi8ZEwfdYXGMDnjQNPOskpL+1zaBB/Zj
VflJAAGXdxLhFDcJQ0d7vl1EbDcnY8B4J4MzvGgVLkSW1+sHjFeadYrDbbfEyC0LETh2vG1pf6gh
1fpj8pHQgfm5I1SNLbSiy17vetI0h/8xBQJ5WIEDgW5HoNTty4hXbHCqq9Soneq0ak3Nw8IrFCR8
LGvgfRQz7KFftTwswOWSdx17pIU/hZguMSndii1K424ZH7XIqhbuV1REU0FyMnQc/W9XPK+ksqr7
jIqi/ndqt/nZIvrkPhmcyQLH7RVsdmJco9NqpAG2DAE+AFOgQgn4dT+roQH0oYNwsBnREaXNt2XK
UknJbZCBtOWmJxn6kmJiZEz7RbgmGwiet9EtIslx1D8NdMZKqdE37wcsaV/l7POHeJQ/0cfDm5DX
+9WQaJ/CQpNTeNfYClPCkDRy1OKPFQY7LdAYxRjEV0FZwCP5PZ2uf10TMiwWlFac2F6ZLHz3AypU
zc2D4H6yBIgtQSiIaC6mwVz8CxDj+nmhgcN0eNfaxtWHfrElXp6lt6eRossGeN4JxgNPtuUbtXf0
zmVGoAs/uI6lGSNHtiCfMMof+ytIJAzVb+WjnD/wIKxvbKKHDRx/Pd6knNbjK0L9iFhYjgZHQFkw
keC6ih3iEo6/gDQKb+Gqc0V47npayfrl4L0Txvk/12sjIhuAs4uBJoTo5w3/1/5oJvsp8eX/T9ZN
df5PulHYsPF3x1auWhOPAc92M+Kc5OtoMg3QV7quytDH9/8uWIXGqK6X1toSgpm7LuUrV3OghbhQ
vDk5TdMg29c4Xb3NjeGzmSoSxU2Sq4fDLOt0wbI2P2qqBuSy40K2IgKZEzXsJeXEghyKJ3t7Mccp
8WZuxBR5SaxDey/jhBHjYdowZfJ77noh4pa7hBFVCxiMVC4l8c8kds/Mq2xsDqhMRbXXvRXG9Aap
140sN2t2JS195+3lSLExuvLxo2UAt1p+eoGJKakfMNLHOwDzxuz+/c0c1dyRabMt3EBEmRZTifDG
AXa0H+/QqAwdHsRr0+ResrL3XpLBYdtSMXLlYipo64lnhV9y34X65ShkumSwAJLNjNBSfZVYA/30
TSv8HFqCJr3JSwnT7X7tcFiQ9vIYjTmNchTS2YDo5hu1wwujKOTkOlXCJI7mwYNRdmHvN5gkrSHg
cEQiUXmfVq4Xk6dTMoarF/5Aw0l8VVTMCGONSwdtHYyGVVlyAzCIKvb3p4bNGITu4XG2y6NKjdu6
VuZsG2EZvstcQI9W0/DPJCoSQeaQiMUnTtz5MWQMOGlyP/pceooK1hfk2jNHEvBgHjYqWSc9+jvQ
pRXYufXvo/gSmwH8BCCpRw94iGN3d0p2AyRlkPSCfiE4AOy+s8/KrTETPJyVC66/DBARKw6kfUER
9n2fuULL4FiYtfiHJpJ+tfBc6h3Nat2nKIhpwjfO/QdnKqLMg5AA4BhPTNNly8TeTrcVwJ1tHiyZ
GvD9V/7nrAIFNrwVku7sINCiQAuvWfkuch0H//t7Ey0ao6hQBN1Gtqfq1TlX9CNd55LEZ+v72Ols
y3a35+Q5IubKhsYRkxF/2v2HQxKLiKxK8ae+x/w63XJhA8EVlBI6/K2LVQ8jKn8hHrqWFI5OGFlL
LrFsoSPlJH7p6rCv3Irzx3ihVoFxn+Y64fbxyZeeq3M1MFT/vNB07S2p1rwgdsHZLId9jQgRvSfB
J349qkkk0w05AbS6ASYq2nc2PeMgM3dzckwefuJhtJ+Tletq3I2oXcL4WhJyXZru4yrwdbYNZeSQ
le5TZLN8pX73eXOBzVCjT/pVycI7sXBbLOq4FxbVWE34Z84hWSkNH1+85uw73ZroiGiglECWhaEj
Sl7sY/KpAGQOfG3UY/s6QG3UOYBgBViH39upiNtEpIZ2txSBCiKeGwi/i5YXgwhGSx/vL0glgJFj
soMQ1cXL6F91AwFBeWg6HaTRFqTgUUTTAH3Iv1fHPz+e6lsETBP9AWrmNcOQ3OT4dd0usjhoBdYc
tm50Gn+IPYvP5dnOwvQMOo3NtKyJgHWbJ4W9jv9dDHQESCCBHVCRIVU9+DGTc9bcG0MzWIkDULaM
U7NVwuaHRW41InqIftpm8W8jc8rGD8puWhYolTlPq4VYi1VwnNqqD9pipmf+7F8ZqzVjQrzM5qg4
AaXXGjgGn5ocjO6LanUPwfdJw1yIEbJl0GFvDEDGGbqu/ABLRnoaQGBf3OXTkJE95vl2SgosLm3/
pYmX5f2xDMNJaIqvCU6a3A7U1Wqiuasc4mQJv1ds3Iq3YllP1qinvYn0XULVlyfbh53l5dQ8yf8h
6UCSloDTqJ+nDnmgo+z/IhHTOL170GHhUXxXMGaEZstqhcqsbs6lrGCCRAwE/hKwKVZCHeDSio6e
WhFlygKYt4z8vrA0z+gxu6elhbQy0m56J3PFqK7Q8i0uJuokiJESH44hrD476Y83u0qVr5XdvbjM
pqazPNf0jd7wf2d8O4Rn569fJ+rGf7mjCtBD9Q5tq6f/8ZOtEPgVOfNaCCmUDY864fu1OZnKzPvK
ZrmbSkd3DlUZCb2mql5DrzmzOGKAqoj2CFl8erI43auuSCYdoJi3nqOh5ESsbP/5sMq+cp0hGP/+
mlfREPaiPOpQX1gYMaTj8yhPj9md4t/XjWds7REZVPknBkXlCpn5PzOR/A+b/MHaCMi1z9+bpz83
dMFROaGhTjwKEHzwGfFUui/5Gr6FafHCLoSW5z8QZnZFMTuxPxnUM1Tz5SnuDNwet73gdKxKN0Gd
PEg+QnSYlkhS6guLDDvcOXkEBBQy9rp+LTKihXxcJ0Oh8xz0c1N5IfFJMUCWk2J3Ki0ea/k39v7N
QqBfF8orJ7r3REX4fPmG0Bj/n81MHSpfR+bgmRa4Dm7vswvj19kKYl398LdldA6c+UlDRC6fgF7b
7XxElRtyjVkRhmnHmyxx23dujvSD9VIyLvK8QLcwo6M/pCnO3/8boc4t4Kt5VU4IhplQ8lNodR07
m62x+ih3nGlk3uz5cNlun3TlFdBEJl9tn8YPq/lZ6SuKUOXJfkxdXzIseH7sfniMlAWWGM//Ol0o
pk/tz3ql5QQ0cGUjdPfBG4Cw7bb5YlFRFSuaTFHSHRcKjTBw9Vep2TL7fLNgQIrTZv34E8wiAnd1
QoxoEvhFn4MkvUIwPraX1NtbLgeRJLFwbWvlKU7/2eLFFxNLDCX8DCLTRW2LKaFn3ENv40Hjniud
sUDogAxKus7kIzcsbGfFpBGxYamxfylDm8IlS2YS1a0xevxSN4XB/HSWL9BcH74uts+qb8QN+AOH
ltH+w6yrTuYo/dcC57wE3yycAUHtCWYrtmsUNAEEEdHuI4gc1D5sL/4yynd7r7inNdR4PF6udw0/
RFP3aHTG7cUHuwvyJgEgk4+BHZ/NJdmkyr4Y4mYzP+NzEdDQHQj4da3M1y28QKNac5J9uHrL3EU5
e4/FybXv1hXkYe2EADDK8jg50OV5umAJkko5vgp5I9Cx5oDnOE1ZEaCjS2hyqnm89Kf1cYxa8+j4
66JVYoOeCWS/HFkmCMEFTpbmC72U8EAhIBx3ADwrKjzARNOfGKU3uj3lR6r7Z8FRSvztQQBaHqCI
cZ3NBIDWXBrQq5bScnI/XQOqSjSsudIUfbBHkTIcH8i1ORtmDir86gwgE4xBZcweuCQy3ubkqh7Y
Lmi6zXabk/96F6f+X8XYVFvf5/+SptFCKNFL+zcgBGiHG+ywB0VnAfabyXSv4p07A5ke3RBsTMez
pVnlJKhk88SndLbruefrMhA4GdQA1nZSkWx6BIS/NpvUPEzYuVpDkq4/pYnpUhQjQoWfgZGI0dyk
aehddIpRilnhdnp91WD0vMRCQkc3spRr1ULxFLRi2rgvucm4X2hpRFP6gLfkb3PKby+S2QKC7feu
biQUAxpEgtfRtPMnrdw5RapKNY6PAOCINNzetpzB6uNx+RZcQHCtYPIpfeaQW2BID2QxR61d8HPx
dxaz4yFtLbnr3gEWaakmfA7inRzvUbo16sXPP4UShOjxf3JU3KbZZUBGTKrCm+XCEBB0DAYoV6IV
Qa23PBnR5LkGY7ljuFQrltBPolMCSsEHEPfsvCL41feZB/PBG6VGmXz/W2IjDRrQKeLGP/YQp2M7
KMBXuM8Cjj7vB2Qdsn/rRt9EfcRdkPC0mKN3pYrlezv/PgfLFxynsXqHkRo2FiiifaXHXbFDM1cY
Tl5IyZ/cbHM7hzsQMRdv3qwgT+A3hhmIgH11mSv8Dk5p1b/pyvD/ozKY5jo9WtgDQZRhNOAgP9NK
UTdWM3VSu5YPpNBMbwQrhC0au40x5O/bjAGiC8BrXO5agAdsxCPbwV4cM8kb/ew+H1dZ5/24aBwC
YG5vKRytZ7P5hSH6syVY0/JoepVGbKVLRSvbFJ8jnvsRI41WMqQtOmNZh2+3l+jLkeIKFWbZESai
OcBbJkUfZ/jq3zPVX155WdCWzulW/YiNGP/8a18FtclYbZR7ZhpMVBHZiZwJhq20z0Ofr52kDa69
X3WK3hyzIA3/RdgJElHsWmv3aPiFrbCqOeWoz6IbzPoQOfTH6LZ9SKWhCiBCQVkXYWcCCVSaWQku
CWjxaalWNJ3XKpxuRJhReEwi8gAnov/dUY0ApxGrK3a90zY6zKxtgYDVY7+kTC+URCClcyCSJhgS
VhuptjSyu7JDuMviQKfTZ0uE6kzd6pGSpKP3Bn4uPpaw0ATk2yxnReyaNOeBaTsZCvjLGHpd/x99
liyD7IsGpJo3xPvmvMTeyNb/xAUqT14205s1IbaE0dJ/OtZ1S2ZvOKBy3WZSi3U9Np7irGE1KLvf
irOG6yysg+dFXMnG90Uf0C6o4P7R/KkcGZiKPi+/lYI2hj04GTzmZo0WuZJXpA4LcITv2CI2eEvr
4qJl6OHfKOr1X3/3YoOd/hwV8t8AFFa7B14bELZU3s7AtDBBroO+ZXnPHIRsMfLzVRAYv6+TURN0
WO12eySXdy1cQfR3U9NY785LtrLU0YHhGeP7aWtOQhfCPVwdlCRmA8ZRDweU7iSDbtiE9MNidd/e
GOrrCISPhZyJ+nI05Gw+bn6DuaeQeVqTTrurpyLWTqfH81/nuh5gbEeSXKFC3tXap8FqZgcHie9b
hkpxYXHB11JkDdp0ZuqzL4w75ihfyEOM2B4jQMnnlMWBRLOjqJ3u6CnsZxGzORP934bov5y+ag6x
uHU+lLjTle8TVOFcjreJnKYzZ7LzXKZg7u5ZsCoFt4dIlWmwPn51MasGEOBZf7sY3VkYZkHxqFMP
P2drJv200p1idRrVdMWiUttKWsQcre1HzG8E21fOzmEuLBV5nRIqmgd/KFXSqxqjkS9vmealMD7L
FhVVME+oh1qYKr54tOUjcH2jEWA4zeoj3asiFZ7wE74uVOhyGy3SMJehIkYNFkWzUX6XAm6s7rvj
lLehNoPDEwfGCRwGTDlyhFxwQSrTIqgoYp9ocmQUfFUvB7xjGGp45abkJJgM7V1AnXY6mBMVoJ4h
2vu8ug2IQk0akNLTXMz78r9W3NE4SonHejzFsm+Sy/Fww4aoJhc2qhwKduKRGXP0LZFAlYGi/00S
fLPd/kr7xZRceN+RW8nzKH6HtxeGrO1GZNXf+4UDTmvt0yFd0Z4+stUZuplvVxK5N3C/NM5A+uSr
3Mox6cKBM+WP9EkAp6qdjM5+JUQBLvCbmx5jJ1NJbJnfI6GdNMBmcXhWQBgtfMmaLb0zKeU3t2DK
sditOrN6FSH8AVDdmUeKz0vcrckH5QvyQ8YabB2/Q3RmfLaKUDpfXpTBHWKEbZ7bmWlsRozbby5N
beHM9Vow+08KbC920Wde/7OOJWVt/4iSCgiG4HqHngCxVWmQ0UYRdgA9aDVMjem4vbcTBIgwehJd
ob9j3et2D7ajcQz4q29jWNFzaFYubIQHYlkSn5E8kT57A+RkIdJuGzffpH+XTtCroSWlMwuhZI3M
SW9OwcEghFBjygaNY5JPgwFFHYFwQK2h7rpMRIn+dhV3zahNI7jJMq0LsSmWGQy0LKrcfhgU1Qx+
IUB1SuJNynZ6ftA5CW3GZHNmDFq+XwxqGACdGq0D+aFEWt4ITUbJ2dd4r21jooFwUguJruF/Y34n
CrCjx2bLREF7a5Q799wzHVanqhzFSVeC1g/dUHD6a/kR2SeTy8erdSDwyXJf3ZX+8tHKUDEJNFtw
IqDCdrME80WMBTa8V5NI4Kp+T2TKd5m42duBI+ZFXbsnkxAE+JcPBSAtrb0rf6eOUENyEBMypOOQ
+YoQIeZNf3Iq0N8ixbS23awXUBmCujgq9QsrB3ZdTNlZiZNrqDX4++oIDBuI39XK6AtAqRYzjDUA
BFRbPMm3JzEvSkVnpm4VqCKoYCdfFOTEJ8k6v/60KIw6diHvIVA6h/DS9Sx+rMCzO6VIDwBuzvu/
Bb+XHgY0BvEJflHuC0hwNur3DmZVHKM/4u3E5548jqYAtLlVAQhm/UqeFcmf8rv8ptrHLCQgTfMk
jjB2uEReWu5iCLw427FTz1pW/XEimfTSqmGsPjZr34LGrCUBzpuNmPZcVQDehNF9nmMmGqb5/m4u
WidH0TC4aP/TaFfuTVL4iYs6HtPotKKmsGvn2loVOnqKSVWrR6+OaI0EG0X9uyPpAGFN9TveVfpo
CI+WmR/78tN/AYfB6uOAoOWW6MI7YKbD7eawoFZ5cg9UI7YpU/rtOBSKbx4QfhVSJP7YGFgQa2Wg
rpeotKJaz05DQdB/kAp8TsWVtCccUAkvrJpidD2xrKlfCLHU1Y+0uSiwSr/PFVa7u3Xtdjq52RGn
QZkl0BSH5jNCbi0aShfiU8zxkadDQJyV7SHtfD1QQkHT1yOAIcKazAOoxKJMfUL/LbGarQBd2VGq
hjbchPhxjotHuYIBohMQVLDBQ7bAVwUwMMmnvbXQp7gwey70AP+MgQff6cTfabubvlO1R6u6K0el
BZG8VhBV5N1BY9l9vDK1zWfbOxIzvcwbdm7ZNHoDrBppgsmiXr9sJy9od/48cOg/5DtBKogLrJOO
G2zQwqnXrrAWTU6olzIDRcLNt44Kw07pFi+PDf+gJMuOKoAayVwU5P+ugBNXv7NfwiPt+uSRh988
gSzmL33n+cjAcQdQJVUMlFCCimCqBznz8hlWFP92SYfx7gZRUDGlo/+5vHUIeRVFAPg+grvRMEmN
h/lXUiioHz9ZXAqpnbrDh/qEHKfGh0zxXm8BjR7kE+U4RNoTkhtrpm3lwjonMbX+XPEeluFbsYIf
caZyQ8cSE9T+BxNl4LvK6W6cuzPtNPmkEX1pyS/K7Ks5K3nqgsQR1yitXlZY/kCyYw4Ty0UnfKIM
a6HmNdOm5QySqtq45K2AF5Vs7VgQDJMV0Vhlw/QSdHQW3UV67Bcc5NccOR1BmHtVMdvxdUMhnf3n
BB51s/a6QevouapOn38DpvfArjKWrMp54Bc+cNLSyYqLjlpo8Yb2vkt4Sqzl2KCrqYgU8ewXdeBp
jzOjW7KsbdtudCcTL9JeX+01gaZSGXlzryr/krC1xniDZo9HecFA4TpVhjaPgSdo63HqYHVgR/SR
yYw6r0xGfwEq0Pbbj8pH+WMkPahc0GYZOjicp2lGCkH4xLQxPYarh/7h/geRcTTj7oyW/4Lg/sX5
EkJe5K9JyLVTtEfae7+spMzN98HaRrBoDlj7PnE9E0R7EudNbR/jSfJdgCfVHV8AXltcKeeDEaqZ
OJlkzDZGpfg6d/SOtOE1bwFKQ/AI7HM/mlpO/0ORrRVkwrAUCQZdyOXn0xe8bsDhXm/pZHrlj8em
q8pxX0A82ZA65+MJhsnPvT5Hj/IjEv0+LAROcFWKnVsXazcZgR0G9nJOVxqO4qSSD4Z3y/vBGwZ7
ZNAiBtbXM+I4iOaNcaQjRYY4XspDAe6XHUghZ4jSGddTT78/4/HCUEbNnXD5tTFgHajS0wlQLozD
zoK8l4wslzyH72pyewMdvHdECEjozsWMfEc2+MKVv//FtBogMU0L2+N6PZgHU6BoygeR5oSuMkXJ
MkLU0XMnmIdKAuOb3rG3TBzi852/xMs+53WGNGRpjlpBla4WJ+BAIMwF2lg6zamCJ76Hi5OvEu/F
aXobGq1OnjcaOV9PJkrTifwZA6waaWpS2CxjiA/vffDi6vNmEW1EcW7iuos10vgyusPc1Obh3nvF
mC5InclxS0GhYI0PiaTM9J1Q9wHSbQGHe2HQTNrOzSK7/+IgbKZTOoyHQsCtZvwmK2pESnU634Nz
YFIkCYTLIq4bnqQvrsW3e2QEgHNsLV639Eg9hhku12rC66ZNbwKW69qBgXBbD+vXQXLI0rYpXDdb
5qkOMx/4TzFEjjUkXUoQxddw69fGgZlRMghXBpscUSf0mB+N6GbYC/E/fw6T8wa30KfNv05NoVL4
rXjST4zZYqvaZ1OU/48z7Lvw4+KQ5k9PMOmdJ5a5wh6kvYrtfXCGbhHKLjytBYSiBB/JZIYyl+f9
AtGIyeQGkSxlGC7ITVuDDJpoTIx2bMIWnMKWEgmUALTXHuRVGHyZ62jb3tcFJfT38bm+dD6/ntwF
e4trIQOwDmEhDZ6+yfsNc9dSf/CS0FbsGUy/t2aznCxpbUQt7RW4+FjfJPsvGQspQgDrzj8GgeAq
WaOTnqVNixVWPbL8DlXnOG+0IXPGUJKyfGIRBNmVcEkToRP1bzBuvuro1ONeZXf++iAJ0PLISzu8
951JlxB9Jkb2daGCqkTH5rB5pmyWECc4QgnyKBE0qaUIkXvN8MHcX2axwyBizMp3oFK+xrmaqysF
UYpzw8SVVt1HWz6egzSIVvrQzeyrboje8we9+PmstiAoC9VFrFlirRp5Imr2HMp6Vr2u30r5MoYz
iP4W5NKESHdDl62UjZyAeA7ejsnNUaJH+CcUtDXCnmDnXd6S5wvZh4e8LFl+/2SKWoPtU7pm2rzO
KJBAr9FvItIOSEFa3W5W8wJD913AR/c6C0PgdRtWIg2nvUcQ1YWvUmvrohCi/20WAKqyhv36Xaug
+9cOWugvTrV5cGswKFa6xyxeIQMfiI1Fp8bzmenBbUlNXvN9ohFzGWU/eqGj0dKW/7Uoq98K2HEi
UHalsF9mzQKvLxIKLNu5/rPQkfFrUy4uLydNv230uOD5DG/ijEPdsBwGcTvljRWTY3CU43NZsIwe
DqPpYr33ryxrKO3q1SkE2lXzVg3400jzFM/3292JvKIPysOV4Heawe7JfhKJ2yGnhvk/6Qp5G6I9
h3ZFUWbbf6KS+YiqwCZG7BUfDTrGqG7EUd5LDy1w51lVa59x5ww8wlhH0m6aA60cE3Njyx62vVyt
htwr0xA6Ju852EdHko/CLJYkV1mM+4VWXAZFtcIKuDiubtpsIYnrJbdwh39Gh8Qo+4xyPlFyK28F
qGNMijz9mU1wif/q1yvRPIqZF+vs1e6C8I3WJ4rMiBLu4/PZpkW+Mz/ZeAPwC15LmWIPxdi/+5lR
aqM7JBq2mxzbV4t+xK9f4fH5cKSqmnNhEa6QxBHLoHXG3z+eRawGXXArBSLs/JOD5KdQR4yiXR5t
1x55FGYCfiKY8BR7JAcLk+7iLZx9Y+4y0dRYq1BSVrvxAXVVGfX64qNdSSKPJYB7rY7cJGHFLGo6
hckr4HlwvkpWpQMtJ5oYbC+KTMIZaY7WakyMj1xLbfmb4DTWivtBRmtBIu9TTy5976JrH5d/zWFe
Ik9d5DLuNsItBCJKriG+nh3iJ7jreULw97BvB9isZY03OB7x+NkUKldkkaynnkO53625nqqwOSqV
boUo6JA+gC6T82mav3xd5r22xzrqvy2qgyKHyAQZM1se2ZTvsQExV84XggOCgF+wsaMpDXV5loe/
Dd+yiK20nqgcMRnB8RyZYTUJ9vvqY7zgCBJtoY5W/wyPr7wUwwtdcGkmH88zWzfIvSi9DoTcKBdl
IP4vpYrIBXIPypVPQ1nqlUILCmJWKfbP4XeS27B76x16hSZe5qQWoUr+k5/2v4CzdGIutyQTL/Lc
kSGstno1M8JGTsL2sjGUsr0mQLBoZGL99aYDKbrUJ3Rm1JVR704vUSWWwAlwSPvcsH0f3CHHaT45
BI5Qman7pvSUmKMYfJ9PgOgOr0GOB+TqKxP3bZhER/kN+DfA3as2ooq+EdJqRQH6mKe15Ln0OVko
i1ORfID527um65tKhPQGagiCPfDfUHMB6Nf1wfHJfGrMBaSXxYmdgV/HTBs2tdGevhTAtwc2pON2
xfEQ656eopHT9Jpi4SHAUPvBtoZHlVB/MxL4geGbWsW+FqiMxpzHnQn0y1hos41HuEI76eSeFcJh
P+ZRVz74C/coXspDcz9WwZeM291eLNCgs3qW86ob3QRYoTPOA1yxRvprZOTuzha+vYUiFRPruA3P
9ikJ4IKeZj19sqhgwpjLI5A3I+i8+YzJnlGKeR79IFPZgiqZClMs4wbnbTwB5iuygC1k6lLvaGZy
w/ulPbNAgw9IsOCxgzBQ35i24Y6mhjkI79RV2AeHkLj83vrMjGVpz4TSX897gyp2nM9BQNRp6YIM
m7N8T/bwtLNyy0XDuWB2jfqQL2TdLGNPOOqCo4YH1MCLdDgxBd/jHGP3kYONMe5WaBn8xO5NruSp
qR80Z96Usjg9QZCXl992QpKMbvI2dDCHEBfKLYYql1EjX/SiQqGYa8CudkHcloLNYrfV96omz0vZ
P8RMpQ4eMCtBnO/6RPIwaLODifVushBVOFCeZVzKy63bCFRgjvufDBBBNl79zA88ZCEOx/In1rjw
enZZq21lraNMFiVtd/ubVGUN/YAw1a+H+v1CSH6qksw7dDzUEwlcM9a5M/2YeUx7jLxO3ShFooLf
LOdS8TjyI3H1xAi4OkozrYd0OSdK+4AgcXhL+p0/3xwuBrg6Nvc2VL4o7PGjax8MxvU1oSYW9EU1
JJe2XfAUweqPByr/XmqJdthn80XztI8ZqqQvWG0P0OIf+YHD11TrEAXNegiAz/3jb7cY/OkJPsu3
5n3eFFCa85lWgS6x9cohcqb+K+qG3bHKulngqZvakGHtzuxqfh9jSxBBP8U8IozCZUMZUaaFFGZ8
JgKyCaD2HxDI8Ft/6+abovtZXaIJs6iPyufBmImEoxufAbFsSBxbqy1vPjd/aP4C5SEKtS37T5m0
0ZWdU+l65br3nBKbMWEK/YHO9maQr44obMg+Ny91+aaWCzmUM5JjaBOo5Yk+sGPEEUEZC+eonO4L
WNGdtpYaq7AG3fI2d0dE4UDMytD7m/uZmzSR/Bk0vd+JKKPvPSFSHkBNwHTQNoQ01Eu1EeiDL+5C
7jLsriWiUIb6twy5EfmITu1T/L32M55kR5IlrG+4Vp4kSfnjygqh31bGN1lXRAZ573nVwH3C0GEB
1p00gV73em2+9wSLT5CwTm87r3g6CGDlV4MoZIX1zbWZMXb46ObT7bTAxJT/sMFnQW3c4R4CrvRf
3ZGHgVdgK/g3xqHdXaOGOgiTt4ncd0rpBFlpYg8LJaLnJnKIfM1q0jtx9vqwACLW+nUuW6Bzpf8J
bNiaAb/LmSCP1aGgDRVR59FfgInAnjakOtupr9pv0Y129TTpvPAr9nVQXBU+HTTvsCmHS+K6AxM1
ssP1YNjqDK8n0UjxcluHWopTnrgvoA+iGqL6083eBXkwAGpzHhiEIigqmVz4Sy5urWs5t5/e/2HI
PjwIdTTl8q2pG5QKEDEcv/hPNVnOUAk2Enosd67hJPAYUm3iWsl6PfAIluk+Ei2s8cdq6W92TSAr
wrX8pbOhJn0a1ZQPxDUrxIBqJvL6bDNiGozcyJZLomj8ZeSQ3kpb6IXvtG7sXMUqaNVs4aspTdn1
EGS9eWYJWaVitHwpaRQiTEg9KBShizQTOx6C6dvl2Xsf0dDkHX2jkNylnTfdtwNyX8CirOC7BNsb
UHL6liSuUayuF3pTSBIxWjCPqspkeN6CYhIToSI8oyFG4POFHoy7ws4pj3W70+sJYVo8e2hFwlvN
C6tHU4FHOn2ngliDWPJe4eA1fxgNXbkad2Rdtz9ntZ4HpnjFJsFTibR9oYqkcKZJ1T+ipvmkK3Ux
oTU4QsEPqzsqwI7uL1LSGOoNKlSqdJI4dl8zsbECIrITZkyJ4nFcXaCVTtZddHJlkrtpfBli/oN4
NvFjxooWgGYyD8lHuss13l9Y3c3BZ52d9W9+wnFC/2ojuoWICIDJtE4gaxV30GyqeLcFQxpqNKVb
ywtNfb0tx1RtLdzfmAYUpH0MZQbZW2Uw+PSigvegefA1ZXLHO0N6+tpaIjcDG4YbsjUW/xZfz8m+
wupVHHrWiPoLid5ie067qz6wWIn9qSMo9w/NV+Sf0shAIQviUj+F/saD0+ccQYlGygFj+fV20IES
/ssGb+gHcq1JSlgestxF2C5rKGCMtlmZZS5f7lQ/z2NKVxChLJnD06ja+3HgfZRYrHBLpX8t9wa6
8/lWuEig4lS+hSSaAZupUcZJSPhhn0zuuTlBad1c+K3EnGIMNAw3cPqy08Zas2oCwdx7O4ZA+XVk
+igKK6wL+JE4ivyuiK69Ngp54ClDu3wUe+6uksOuhtTJR6P78ZgiaumwVo3G4U7M48TMI+Qv/43X
AAn3XDd8JtlbWbRS3JILU5yr+Y+Pof54nZ/Zms+XorQr3Aeb/KpEgOO9+uM2lipHwl76NOA/w+CG
sfr9Kn56hBwRLLE7BgWS6PS+4Q4EOcVGStdHj6KXLE5kPBwqVswKT8F4SaQ4MtBCblPCgBzeUzF6
5Y3ThAE64gFQtX5mdIFLr0l/2L1xi3xkL/5PaAsytTbyriqRxKCPOztQg/sg7putPQ+xlXA6k0LQ
ovU6gT/Z2zLVL8MNgRiA7cohcIFA/OdtNZS4ri9heAOy09OtirVLGgU1sD4SYSy918f/DJnlntXG
MBD0sWS2JihBtxOkGk/TboxNp+bynopOmyZdc8uN+IyjohG1RIY8HfwndTdmGnMU3KCDrqW3fsgI
omG1DpeCtu8U9jDXdoagqRmq0sxiNq61EGdDgyPmFmf9Jz6X5vCkXrBvr+42CeFN/YfllffZzPfE
GFEutL+jJ23C0ErwJxfdMgpeiRc4iQrptzZgOw644JBL4bjNajb1lVCkIuWkxxvBqYlcA0Mysep4
hWtLoYraAXpOteXYLbXmUlfE5wLsAd5XFQbMUswAE1MTVWTgjavDtFXTmHfGUCML1t5HYMONiLrD
Rx+DFQFJOdtIV3xdf84zd6PWGJUMGMgIYKJy1rfSHlfUib8bEw1WKPh5N5KJfk47TBZjFfrKl1PL
ovoikfSETbQaFh22fFR6MM4ZREy5XX1Ei28VYYTAA6I8mj7ml8p9uylHd34ZiRW6GCJQyhpJNCup
hfxZKEoZPVVJgGDJs90lVT/C98QSp5xVYvmpATkjr6OZtcrRGW9UcMWO4eNNqcxO3pCrcDzioOLC
ydLgs7ahWtZepjZP9Ujkt7J2/TgOe0atPUPtWdcbIXJYM5ASdUloVHezHh4FSoFWYd6caX2Bt6J5
nYqvRix9Pp7RsUFBi+aP3D1sXDWYb4uH2SPJOWg2Gz7YzYQZ8ouDoqxaK4zliLgvwbgjvGzXtV2t
69DvkOo3VeYvUprb45JWZbMuS+Z7tcNu4I1gLUr2ia0un695/3ac7L4lXCJ+dcPZpkkt+pgh20RU
RYlCSV4XRdieRI9OXaSUtkMgvd7Gkbwr6YlTSRF3gGsG8o41h0VkfHBHvh3oInqOHxRqfUKOCQHU
y1luDDDdtkKotRaPdRER4hAkNTevyiNoX+KVGNsvG4TVLT8Nkh0iKmaKKFyDYpTwzYfApVBjvj8A
DPyt0jlvn+v7r7hMiCNzeOfJ0DQwkI5WRtE81TN0emj0zpnddSqHWhFWRIup4k2TpSPr5XGLNUvi
voHKpYqs+SHJbWasfyqWMsAbKIHst51HtRo1JDTBo7BMzc1z8DMmd59oiv3aAiE98rnYT+NappbZ
t7r7xzEsKweraEBK4GF+V+FOxPqQvCr5gaSuyMPyKBZffkUURDUvTR38P9EC6H59d+pwCqTGvPlD
wxOr+E5k8q1yWeXbguJCU8CeBn0btqdxPQdqTBnxkIDzw5Ky5q2ejDliHXjal1Iu3i9FzLLlSgcs
yHdVpHpwroVb3kNdL8V1YZgwtMwkCt9NVLSYkMnDYaOdwQ7PGmiCp6seoFXD5evzNDJWTc4WvoI1
QJN11BN0UzOXq+nKH+WS1zHY8ZXX+h84T3d3lPX0nbhAlA/K7IY2Dcw9p3NGo7PdP2m+hwStCn0z
FS8eACVROQupAr8cxtBlrGIxMihAtE6iTolq4+fOG8SHq21ihMYpeXbHW1Tqc5TF0FvAxQDl1NEZ
OffomZ+O3hbQzh3ULOq3m2AFmpCi6IheDyVEl03hDXoZcV4fctVLBsPhljK46jBTjomwbMKOahaf
oK3msH79GAWnR/M228+GFWX+ElpLYuH59pHznxI/HUvcVT/s47NNNWDBmwi2+aDwhdq29Ks8bW5r
PF1GR0xj3xts+Aww5FIET5ey5EjFYSuodzhbKoXoggXzotUZ/SiVKiaTL41nz04U584LOYTgR5A2
DQC1/jW6zjrs68YMXaHMjRDQohZtTWtwJ3ploJsy+b0g8NeIPvauFSWb9mPhxuJyOSez98wKltbj
aOHVgr/mdlq6PdbfnUyAd8l+cLN+GS6jcz9Ib+bIigN6/+sAKxHzCQOM3dAj5UFJfq8lktst+WWR
jMYt0z/pZFRwC84MUraPXOYw1HSDat483grWkicR0MKvd9kMachdX4j52Cmem5rSfoOqOBWnNULe
rENXSgpfGSsgmYdyUVZ24VhhM8mmYnFjWtsbUdnws64N/0lLvZLyNJDL0w7se3zd2B43/8O228vw
3ZY3z022pkaA7+sU8fhiGlZoeiSJnmfBdlvLwGUf6O+gFVNtL6V/YwLv6YEtvS484t3zQCXtSnCv
5AK7y27V7r1/uiGX+r830qwS50Rn6c/+CJC85hUbNtYuWIQ8D3ZgVkb1I+UYL/T/j0WPUOyq0qx1
3wUlvclwD4Y1z1XvgmKX/5Oc126PUYxLDQ1X6QwpSH7+R2wAKvEJrtIHx4wiEjsU9IBOJ0Yu/tI9
c0+DpCLu+cmrfr6LtGCmEuEs1l9ryJepdDBNL/Jz/Cl/g+6luZ4q8soyASvxM+/u8AcKnW92INs3
m8ttr4qDPXVlAagIH+kw2IwcgEdGWcaS7c1Cfu8GmfiZXGtOFV2zR+mr4xwxyMKJvnXZ/BhrOreV
p7nz6sFsf6+ARNle5zQfCkDQdPsz923Eod7q3QNq4IzEo1vXS9McuwhatFWfN0Tk5ENVHIWJVAGb
cThCIdDkyxRaocpIJtR8z/Bw1AkmkkXu+BNWEYhoh+IahY84HGOsAMUJKnMNFY+bngOnrs9yuIJd
+4LYJOXJOD7ce4Nw9dHEA2yKaDbjedBcKAaSlXxBNo8Vjy73bYD7hp0plpFGMbscp4Hlx507JdQx
hxSfXGGXkKZIxFGgZc7hojkAhgbRfqDiRZanu7keoh6y9T/be5AY9g+GCSsHuSne3hWJQzzKdC03
x9Frc15Pg984odl7DyLogCgR8PdG6fGx+p8dA6tglh4S1ydM6YprsaIRXUwrqOQJP3VFS+eISDpF
3nICqL3gvfrjUuagyguNRFLY/iMSrqB/zGxMolVrKJ3tr641ZW5Is2rnkD0hNQQu8KXGZt4g0ZyJ
RgpAQ3eLX0bLaODcsueMd5Z4F2pZKUTmMr4EDqsyCdSIelGcBa/66x/Q60LImUztIoJ+ptIEHw4T
hkThAwFFjjI/ojde74GBUe3YvQ/tQZMbcj0cInWauUXKvFCHHsVe4wBb8RFq6kZRg99psPAB/JA0
fpAd3xPT0VU49oBbCaWu0e23tYFUB+lDnGZNqScJ/0DMHmmQQsaB81u4lNbjmf4i/C5Erui9ocIY
XiW9TH6mHeF8Yf5k2Q1Vzf1rPB74c+3prCj4qP87jmeAJxPKE96PuIrKqFHETrg+U//QuuUnOEjP
SF4IP69IEdPruWgZggNScCN30MezxU725cO/GQ1xtx4CDJkUNGxJr/SELqJYabltJ8IfZGLI92kp
w2W0NMBcFVVR2wEaOsq2xJ6dEpIdscQi4Nqt78cu8e15ODv10d/RoHygNeJyL4WnPqJDbbU5ePoe
shOWZDDgqfZeY8vlXkEB2AkQOJ9yAGV/Jp16tur0evpry1hF4UTWVIeJGAWTvrnDLUaEfEQhij8v
tyk2AZFaaniaxj8YPerc1tmFRI1UWJrvdkTpBRO7fCkV+oDyGU4rEYNhC7+MdvTTJHja7Qe9Cvfc
bOUjxzwIsFPMczV7Hxw7K/J31ZWuV/lAHkeAOM4eZLJSgRigZgYN0KkJog3ZVD0NAZUbXGZ2k2if
dY/LXH7UBZL1oNIjnxVLU9hpMMAWLjeBmMGsLSI1ZD28cM/zXq6/NUdFUN65LIYiIYURFSXiu6YW
eWOBJz+Zh31ZISfRVnN0mGsmbSPAygrAih9Tqmk1vAu3+zOFL41nvqw7G6Qvehju0nP7TrJ0AK/p
/LbwC5B6iM/DEM/sVjK5nK5kQJFrHhXXknabbpK889tUCOIbxi3UsqyoXYJnUH4L9Hsyuk9xn2Tn
r5zJM6xDSLV75Yvi8e7aDR6zZhNSSZ9hG7WmHyj4tK30u89aqJs8Syletkt81l8vC1Zgoa+OjMHh
9c8QYycGQ1xQdAjXrqShHlIcu0LdF5n9/Kza1nm8tDkNdFETTTy6W9ahcvq8JmvVdvUu0CR0nw+2
k+qwUjFYsbkHaxCEA68tmnjsov0LmGXbFCdwruHVXUHdd3P3mcXdXWiq5k4d2nFTjOw0aXNfuiRA
eeh4wBBKfOFT1pQoL+lDYO3yXxaZ8CxBSMwUaFNQOMfWdznjRGw4PZ8cPgTZT8hepZJmtroRtfu5
QMAaPICvYwtaIcHFuhrNh4glugzEjB4Fq0wmryS6RZsoCRARJ8uOZmEhh5vsgDRGA5YSgBy7zUZo
TmWE/frx+ECLfVzZRRW9bdFECaDiINfJxiPvQ1+lQcBdgxBuRBzMwCXfr43rOPsGfkQx7ujB88NB
1RyezlraT+PSd8vMUWOXLrK8OAvhz8On67kN+rw6OI1x0xdcdCWIALC7Jyz5FYwaocf2MrqvsoAX
cwWeUH5Kp4d7PHWkpbd6I1tTWwAnB/HQQ8ctmjb91GAqy4M5EFuL6pi9N4cnYdt1iKn7+yYVQEYp
swEnaIdcXiLgRQs6tdGiXQWyotO+c8nP82LKSLvzgJ2/b8XFJr8nO46IUB5jOT0LL03QmN/qgC4q
zjcGkxkSo5c3yK4E2O24pUNi172/OySuxncIBZ2v6KFUj8znIqddPAqBiCugheAmEGl5cvM1/Qe1
/q8wazHBsZeo7kqs2hYDsJQ/Ss6TtV2lGTHwyZ/HLiKL9BPSsKn61V+enSaO1GVSB3vnmT70ckoM
bACi4UzWb62bs2WjMHBeJt53A+8rz4AUDEjYEprPB+dOdQSzhOu9RtqqkJIwcXvmKzaruFw8Od0/
qo/BkP74ToKdTDqHyZ7KeNmn/xE0pR5iqNuh+JzEieSCKWRwT2sNv/sPcwXWJrLk5CrFiIj0BPMu
j3R61mPJY28AmyVWrydR2RCHTLwgSZCJfUBMUikpwG90lWYxnRdtvceceybIASOdF1V4lXCsyLg5
U1r9HYNCgPnf1WDTBTW/pF1yt4RVfOW5uTIsihTgDf/CEXWxKH8sjuhbKdxogAkjpxPLbcCQtMaV
ViMuzDef9iajrZuUhgGiSsf/QKGgzF0SII7ZfKorIwN64aACTeGzWAL5NdqJjepDOZ6ClRBq5pRg
tQpv4BxL74LPaZsUNoGhHg+o71PV4+dwQfJ+z+CA4F2RwoFBmKyaNCmtE+KqDBx+ijKHaOxNO4+D
hH/Y0W9G2d8j7Nr01Ny3STtJqRFYbqAKpY6LrDWN8xhL4sFdQkzyx6R/DNBD3HhIzH/GYw2NVISA
QzdRjh0oB+XkjSI5WS90otKC8U/SY0+c53IL9B4I1vru3GPRDJpcAaxf/YEeHqbKTuoNXCs59CJO
1KeT4a2mpTw0+Lv1z8ZmltUhXtptOp/Oks9r2tIZw1uMDtX0dv0SH21Awg8fFfQVJ3IcH0r0/cK0
ovYmBqreB5KLJRhl5pQ6wBBaVBD/uLC+7+zCdLlpDAT9GybNGdm4FPSVSzpf5gEWGZR8HaF5l1ea
VaIyLzVtDD4iED4ySHFMNKK4eNbIGhajnruahooybVY+V1zA9Z1JQLOpFySpN/9gbzJbsgdlFE8g
k2K/ECA+uwH8oIdOoXmYpxDSilFxxgNEos2ijyh7/pre4nTzG/EdXjWMQlsR1JTwp7cyrl5G3MnS
+F7EQtuEomN2q7ahkNOXK0RC1FXuqs1oT+ns0cVgyZSKUrC3eKGbR8q6yKiyef4BQklt69OJaLdZ
DBOjCPCOcUV5hmXTzyfI9NacRl1M4I6INgUVuuQN50FCS0hbLxVOX+7eeRVWRpGw0JSdX0ED5xTR
tO4BHvkADeuH/LjzdkzScLDL7YUmlijwxeyhKq1VHetCMBnsvLwtjobUhEaA/bBZbDamEgHrbdfF
nwFrJfU8QTlCo+HVqzDOzv3s/Rz5BTqsJ7VfVbWUmdVSP2V3AfsbLI9mIB2nUyPAASrt1qX0nb4u
CqencRCowmOFNXYRbM6OgGFiNbi6Nq/mv/vHqls7Ff/wo08mXV3Ce6gCvJukFevF3b+36kqxQQVy
4/aBEYovvt3eKCGRbEt6ASxfTMKWQsdauHGAW+6yCwKqK2yvzI7OGmH4F0bhG0+q+gH5iM2Nw8JE
Jxg1KXQBzI41BHZkUFPNtjDYfcTHTmtNIX1wvSIfNjpGVl/97ozDqk6LRYNDOF4xTloWtrErnqGx
/ekL4XMgTHNzBLZ5npyog0CT8paeTlKwkyg0i4HvLZbD14J5BaIHNnyoNoeV1zEz37EVlzsfnpqS
7rYNML0AO1QcB01d0M2sjFMABm29sfmrmWkkOtBdrFW0PzRkdSYCOJmA6PzCNj7QOvM9K88E5AWW
3yvCAzLQdR+MuroScmx4zATNB6Dg7Mgqa/Av4uhY0GpTb6HD/LG3iTiBgIbcJgUdZgxYqUTkar4/
32LXzPk11ycKPd+CD6BfQT8ZT9ngWtcKRgqaqIkhdSWtdvwwnLP04H4BRL3qqaP4QSISIFZMdE3r
kT85ODyo7cRhUToOg/Iid7KS4QHFIuoSXlQBn0L1ut4XpE7CYaZ+t5oDaFVLoKsNVxEeMI/uUzF5
7T/JUhYhUYKRdXfb1PlPctiZKCyAY4JmRttwiBZBMvl8f5r7g6uxDSTvcqI/zJr5pOCxZLi3i2pE
cD5gldWZspaJn83imCDlUaFit9E6NOYqZcNLnP0srpbpORU2XEwROV72p8qen/ysUhNDv4yHp6Ti
VsNgKOveZOFOlafQEyaDHVXM1SFAfyqMKr2ZQrjRrvtuVWiVHfdipKtvnmyqdK7VxcfxkZdEThCE
w5P/QKjLnw+gxkQcTyxeTGeZRujRAMIOf0OSR6zrzicGMh3p10UmMSiP94WHwa3xcMiFzhT1U4Dc
NdU18kdWuR95uBuwR5FZljkRM/W94hPJG3meS98QWt/Q/FqXQiUqRtPU1FEb/s0xVCp7aWh/0JBb
l5Ouy0zV5Rt8e828AVsYBmzBlE0KhsturkBw8aw8J4qepU/6wpgozYIxOiQcHSAOmG8uvpbJG+qK
JeKQqsAKvmGktfXmfc5gLa/Sb9gyAgGTNDVlusNsU7fCF+QVPULRoGLVkWaF4CaP07f9Vl7dnmFc
S94j0M9ay+5WfABV1TmZaTpkqXZ60XLSN03M5xJ2S+GCwzmI8AGeWiYEUMoY2I5nmvSQdQ1yadZL
7EQ4Ycl6xAwbCwd98PPGMFE4m4vSVlItvRSwwd+mnMETrlwHatYCsEb9UsFNqh/m5m6o6WokrowY
8SZ+Ei2D4+CDstfiIuSJwlgILRnvGXvTpx+TXgGECr107F4Cq//eJW3jS9fnfQxQqrWE95yEu5+s
d7N8Tbb/PHpJ4PHuG3ljwgn+1X2egYrVi5ifVmGjahE6hFfoHcYhGvbDVfM0D+YQMnyZ3s7t99le
zrKfMA+apgs589M0eMK2K4GSouVuktIiTBkD5W8CjB83HCLs62u5qkcPPHIExNIJai/TmdWLVZUn
SlcNdY6+RN4JA4Loby25TtpTnv1kkdnT4GbnnYyXOmDtQUko/bhNAZ/X/zwXvQUL5wnJpkSWNU9P
d8Reab5CkOXO9E17gCqt6Rlkp12nWai3WW6TdFL1TEfXU1tU0AiItUg0v0DDn45diuv4GIl0TcKQ
hsDE7UKGowQ/or8RJXC978WWml+7AnrCv7TDQuOs6yHxNBdJQV/BOx3XJhtV7fWV1US1hcltrMAz
gyvncdiRUihzljzPi33MdP7GD+5iFKhV8CU02Vh/EkTHlXY9tSXComHydwOWR/CzFZkXiNNVfMMC
aBcQTgHgD+wiSABBkbseZV4CNj1CempuMZM+jjr8RHAFL58XyNSvsr/KQjGla8O5aJQXt19yH5ok
xRA42Q4bOJPUfZpUO4yeYpjyYL9MoYmwp9NoeICCXdtc22voizf8nJOk4YgZXVVGeTp/7xJqOH0z
6eiwFIrrgj5Gd79+doqayviBx7okQEu2ypUNqmIVl48IrQTTPnYJpB7vMsb93arQrqZhrBhCAnEm
xQ7vmhK4nnmuVh2Xr4OR2g2kTQH3vNVyuUadmQmBdQiSE0118SgAjeCh3hMuIsOU4HhOtY5ntKH+
ZqZKUd6kGEApZV0OZIp9P56cAZU5gwnp5eH5J60d4Ggj8FmdD6Xiljg2z+GV4K/dEY4fa5v+AByt
3WAsLFIWnch+bMytg6RT5EoHVdmBnm5FRpeAj/wFBsAvjsnHM0ki/3oRXyp99OYx7oQmxqpnsqCM
8OHwKfCiXMa1P/D72nnLwg+mM3iRYa8wEFO1vOMvsZ02qNigyCBX76SbKGxlVyZLsERh4bb97bVx
sQEQDM+Xkj9UBF3zmt6cyhi44a5CnfQaNa1ArUPZiLsJLMRC6z64mnaLa4Naef7fjn2TA9JR1lnR
VJ6P5Cvz8DV+xea0H+pQ8A7ASo57yAACNlAY7iTYIACVgGYiN8kuuzg79/q/HV9ox50RhCCyv94u
Sr9jpHeOxiBrubI+Ae0Yt5+HoJVQgt5kAk8EA0FwHKXoQ5i5df9HHZ8uQzzxw8z3ypqkL9B4bY1r
L+eKY4zWp8u6Bx6w3/7yrkt8iYZIX0oihesrghXEopsHEQh/tdx4A+/15X98EEM7SgijrLLUFBDU
MOS0hoSbyY+hL2fxjbyCt25njkoqtbgUHXYpIoa+luuH/T90FrdB35H4PRMdKUXfmqTz4CDY0Vkv
e8FH2QkcSw9TD7ZH0npOUpnFetkFl0N7mAP/Mirtu8x0EEmIXdDqljYzH2k2DETrm4RG7kelS15M
/9lu77IOxnTUSuQiyw8vf9gLJoSLEfAOYFs+gRE2melKQ+1so0WbxfQVFVunxWZa7T6r+ntqFytD
kLC/b2kLYtj3KNZ2IW5gyDqli/UwX0nTN3uda1RxvUL3/VhgnP0ZVGcU/BrqNE0WudGpWt2rR8sY
ZWBDTHbhwoMXAs3N2F07YpdrlarHCcB6V7AkDUhM+nOci5fYcw1yR9xpOmeajCwZesh+NzBq1fL4
y/3jhI+x1C5r5iOShDgQ/tMrMPyeBBkc+KZayhcjb4ipFBzZqO5wfOR354Y4BkirF6pF+dVIkzk9
yB6eF5dMu7NSx3Tr94X+dyYpkJ2RmwcD3t36JMpQDPA5GR0SpRfA6xUV7eZ3VHT5L7PQ84Oa3f4Z
kR1o01HDdHyWzgJ+Wvk9ePK57wSqCUGb0GmByK4kN/6at8igt04wgNdX9qB9SddsCR5NAg+DHuvX
QEj7+RxIeW/Yv86vCJ92+6MJ/eD9/vsAAq0AbzAVPq53GPFn+BmTZlNmii2AMgbetyo/SC+4uIFw
bKC+1I1e2SFrREcfTBmyQRgTyBxwQPFcn9wGEe7El2EoKM5+zoDBbUSkLZDbQ22w2s2KvY8PjWvR
tbQzDDLHIFKGV+gEQeo8r/f4RMEZwy6o3CdFChP/MB3DkDO/RCfyPlmdxhExT437p7/OYHkuc7MY
3u+Q1iSF94jDMPM4Fsmvzt5Q0kqJBULv8gR09x2EK0cDGLl/MPy9QNIyySeJebiUF+w2/O5ilUpC
qlqOeS25LfbSx4oOK/TbDer6Y1d3j4aEhi03wa9QQVw2WlDuK+bTd8tNhxPvahZ3B5LPzJ0k4QTk
wm5nn4uuoyk/ExcgOyNG3XkrvHA4N+ut/K/rVGpTUXj7EKcEifMI2lzSQpYHM1ALNlyc2Z9zM69C
elvhd14siRmA9QqRF7PzoUDNfnsoxzPRJpuRDTCP7tRTuJYBmI1KROEfu7K/J06YC0R+9/AedSZB
DpCc+DvucjnsYb4tksIj398sAy03qSu7hHR1zcA5pS05x1tiReHAUgRFh4PQX6JucDA7BsD6+DpZ
qtHqbqxF7XCDvHQ7d15NQ5YNxOOZmPdzkq0UwjlhbfGgjNO56SIlNdRKE93tWwubw+K796qK3F6q
Sd08+8NIi0PclevzDNU8ZM23DqOywE+4Z8Qx+cMxIq2Gt77rPvBKHgqTv43trbQpeDP+fSvIeYMR
+7Xf4lkrXbNF4+69hljxa7rYnRndJmboFkkuFRZ+P7N5CzMh9o0Un23P09b/OW+oYEYoOt+EHTqP
ny8zQQEjb4altVqmpnBqk2+cXElkoqio2RIfyuSiImGOhSAlqakT+tvkx/wPtGrXMhfxFVJ5/1BG
0ZVRHX+IKERkUYwlBl+RJ8lVqBeB76V59CfsXr3B1J3EsC8v41M4BKU/E+cGvi2zeZtIll0n5CYL
DC65ZtM2sPsN881fVEfqy2FQvlGRjTCSZI5x6uJibTI+PhRCzChoKr6PO7PzYft0TFHv7XlsQ/48
zRmt0vAbdG5ACjFuo7CldSe+/ng4VNnQ3p3v4FI8tvkYIrkmQ4d7dyspzVecWQebBYHggpYR53f7
vu8D8+kbHN47hOanqQrtv1kwJyBojnVOPEH+yA0DHnoSeofglHW6iM+DOXh59VeJNFxc56Oz8sjR
CnqaY1w75GODmMq7JRp6/oVEqlkFZMptE/FA3/B6ONrqrdX7+djwuLQxylnePOWJ6Ibj/WUdGO4u
SK5e7pLLqtb2bkAli5sBIw20NjacoOfcPVtIIWpLsV40kXh2H+Y31N+zjDTOTG8s4ilucShyGxrP
k3umHMhVd1t5nHj2AMs+UuAGAi20lgwpiOT5RnSD9URHQhM49LQfyNGdDR5wmrTVFVyhuQov47JJ
JjEGvaeUMhv07slshFUoaYmeWj4qRF13fV69LfPOE1yZZfr13ZjOuCXPWiWwakyl6/NsxMdy8eKL
h4ZlOqEdNcliPEnUj/S/DWHrWsdt9+LHOxnPQxiohpu/PGCoL7EZwDSeG1gesrR1iYJVKo8VQ86x
3mPQaRvdnY30vAKOopZYV691+/NkBJjpTwBspe1K91w+V6sb59yoEZ7tfKl0Za7y+UlOYYvEyzd4
zVkG3lzqL31nc5g4C0Dw9EsJw+jOCDZu8NZ8utiuEm5XWDzm64GkXGuLI6hZrmJmSCdi7wqVvjYy
hHwnUEOQbdOyYmr92cPCMTTGjpOFCggjLlUk0hIXnqftLZpXg0KOCnVJD1nF6zS8xumoI/PSDIbf
BlMKtkDg84svn9QLTdGd/ki1KoUM97N8rruXyfUF+oHYzWOsaqUgrUWYKUyFspXiOpABVT3tK6Fr
Eel7CvKeys5u1Y8kDolWk+Ikf9O3y1Y9dKlCE94X6WBeUd0XUKu+HmUZSIPMp5ksiMRrAs53fd1u
9cMfH2pp/87cQSaOagpx7A6pbxk7zTnmHolvSUlJdjLh7MkS3CXcchpXEhAAA9FY4W1mjPrn1J7y
bilr/hF6Nbunm656jcjGPGOSbA1Ln21QU0/K7d2839W2S4lgsXS8ccqVckq7u4OVgQyxx++gVBWt
15bX5PokPWZuzcfsF5X/xXGDIJxatmTU+t/A2yAPqVuAY4JIzUvJkDt+R+DFuGcPYENIeziVkq6A
dG1KSDawwjO5VNfjWtGN34jctVLXmOMfjafIIOnGfXXvU9Fdk0n9qf4QaZbIR3AyY8GrnREDthzq
4jgRkAozDiV926r83tE61AuluiK1gBxGqptGut4VftSkRcKEflPqoWUEuJJuXyFl8W8vtNJIDYND
1Tsbc7JK2mwv1pxn60R6zRfwFLJq+CPRc0d0aP0GRVUgESYOBvSOAa7Hga7il22vh1Dn3D7ZmSce
ecR8DH9uOjN0Z4VT2e/wiyPG56p+kXImlVUnTQheRNbnlGiotNp82gc5dll6noJPdI/aqE1diOrt
oZAptxhkwqQrGxuviN0xuWLzR1lvaY4SeH9tkTYqqbHLT+vilYPAwC/B/sMs4pC8QNEnbL/fF9RX
wt6kDU8jhhDCx02OtHm8GsMgvJWfGT7hv98CWm6vlsgSBUwExFRAa1atmOr16SjhbTcN7kGGiNJ6
vhCs6jTBWeDh7frUSCwb0blChufL5sOQk3NxnOav1xnJ04cQj67sLLBRB2mkSbmYO9U7jQYD8z5g
BdkLZLYMealxVoVmTdZAG6A+oLDAv2cisx0YUmK9UMfJ/gsbmuuiAFDtcuO6zY4UeW66CMjub/5n
gczNAUurS6Bo8mrg10qQ3mKTE41Kf3O1by9LMdryQ86exZ6C1DlqFdZtZwhRIH7MBH3+dCLN761L
t5nYLsoByu3ibuxvTEPixEB0Yz+rKdbV+DmCgMirU4wd7ekS5InAwDbBA0MZ/HsDUFifIzM4ES1C
QafOKoCBhdTZ40/IKlu3wKRQRLA9USJVQiuDF/nCXOEnX063WdOHci/eY2U7SnjU+r7S4Lunn5ex
cIaQJuJh67FXoS2ZaQthfvQve396vMeJHSi3aOsq8GCJfzmMCspQc6NPk2N6r5vKnM5zo8kvU6st
LBk0E5x31HiTVBOwvdJB+aeBJCzZXU2Rf+lXHjbX430kHmf5lFL0H0U7P+4l2MszyPS4WCqkd9DL
mGwCljAcSo7VrQLd5I6SaLyLo7+Zvb4bJO6a9gkrKykdpRPMsKTGgxviT5aNxcc1aCc8RXcw3HqJ
tWUVlwN0dJxYezBVYu1S5w6CVXqkrbnc9ntU6uvHFu+Kk20krg9fhIn2B6yTRNdJrrNjH3Qp/XXR
nAO9oSmRYCT92WgvUNFKbK02WoXKYyu3V33NzfYzs91Jb/ls4rWPdkBHXpXPVoAE8gIXQpmXKxb5
ljp8i2B5k3BDrqnXTbcuEo16NcTs+aSdIO2JWu422DuDIzv7LEi3AJT6H9uS6X0k1tszvSqgTgo8
l6z5NlhPB+wGZJgCqLEjZ3TDe5Z/qsiGKcRE856yhXmPYFoqBeXiKNYZrfZAmolwVDJRGavKxXi1
CSnS5qj00Hq9VL2oXQKP4VlqGx3ZpqVJRRSwLjeP1xwkHK86gtg9EhAIV1N0XaV/p6+hMDwXCgyj
QrgEyIW80ONR9FQmrgpRsbSDuwmWpN+a6sRVcpj8NQSmOQzwk6X2z/v2wIH0deFhdHaTBb03v0jv
d119es8LlyY23OUyQjDGCVjBSr5IMcOtWaWFXYO5cPMslaqTF8FVBNlMEoWvgXeu2DQqbs5DMaq8
6wSuH1YjMiyIK79C028wcmVJn96nazSmRkd7IG0oDdqyUpmg2s3WQsJE8sC1vKthnA3EKCrEP2G+
8RbEj/zFj3n+TKVIBaeCVNGFmHfMMDurQN29VMn52SIZWAFfRYeGCnXXoYdTBTmYmI46iSyZXt6W
sYGR12UMQJwn7DVLAgSPFaixVa+hzV45Pq+oDd5W+odgBW2l5eZaDJjtszAiv8zKCxdtgP2KpH7U
VJ2B/yMrfUrloGrQlx/lWaxrB1cvSCuCbYS+0bTZalKoVWpYwgSoeBbWlx7BttLMUAtOPY1zp7fY
3SNafGrESJtuLwM7Er+AR6U66AVKQVrB0DGYSj7MnMEtgIePaA4lwJdZB79ogdnm2GXXCKP9Vdcb
3+voPJj+/DCip14qtFjmQuhrSkpqi3Iv1ZkmEjMvQEZd4zKOyy+puJWFfIzJOogIB85kh9wvnZKN
d3D6Kxqwh296RnjzmEVHyYUIhTBlJEQfsDxjmCzo+iFxnWwP7aaZtL59Vb4EImRD1RaRrlmUILal
ImTUDjmCal8TneiCopKl5ve0D/CilhjH6T5qv23TH85MDs8+UVwQFM4vf9EX/p144zvWpGTxBnYf
se87sr+5Qmp2dSuDmr6R2jNriOCHwhKNoCCPBDafIoEE5M0LArZn7MViMIVdxpMcL3KmoMb85miy
5ra8pF9PJ6OpusG7Sf+Uj8NTqSl/wFh0LRzwcHYYeJEtJ2nGmCtX7Sq1ExHVESNeHWKwko37p56g
hxpViX1QDyloYGOfT6nU910y1N+wX+6tsYvz1wOMqRIMzxmyoU8FGBKeixyQx5JPBAp15sP8asT7
fc3jGmv60dG5U5QQgghA1PhhPseCXvFlGNfVJskx7ao0hKs+G4HHTB0vM+30UQKd5AbP/2ke+a3e
bkhyrQr58k+kga0iDJuBC3kEVX0JGsFmkoGeyZQgYth/rdQd/bDOxKVq1xo4dEbPOQj4d0hgycQh
vbJDEE0Xsdvtj5fo2WzKsTEH1TpkieHyYU8stfa44XO3VFoJ0XUiDYjOoQnQUJ8UTwVPX5WFagCQ
L5LABPqTNjUGFMbeDsxB6NesQzTOklqd0lMHeMC8AEEpUNmiM/qEUW5kIgrCKtjDIivnMSfE0xVD
RPC9/xT0JVeoLQAulvmsfUHCORn7y8u5aTLzQYTE807+9DS40MtAy6c8gc/ZP389oSCkj9XcIfyc
PuUBZsHj/7tLJESW6vsz77K3EVmYp2w/qOOiOmKvyIokvmOcfCVOkBfuaR4ko36bG4H+jxPQ2Qbo
D4xfLY0HXhLeeLH9iAoXFcDFI8iTYhnxYsIflw8YNJzH9Qus6ysdhhvDpYrbr5tBYGxx+rIoOHwT
QW1pQz3snnBMMlr+ZGDerT158Oy8Ds0M+axPbSPAWamc9BmULzNJ0qIv3Wxy4G1ez/zeT/EBtiQE
0nwyaEc9ctUlZ96WDnNXY6mX2Ro9hhrq812fO2MhplqoZW5dWUqSxxCVhr2WjL7tTi6hSIip0jzx
WJd6ZczLnZ5LtJZG6TQym1SuNW+AuOn4OghQ8ColJuYmbjr6KvTnyv89jE3+ncceW6cgFnDKozN+
w8IESf9Oxmwx9TxNwrKWdLlIXhTo+BgtYQXeCObcY7FH8rVuhAXsZQgtRCCv0tOqU6NZpikqfrI6
n0hSMnaFdAR86LgQOOqhJaF1Ya+3KyRAT5xtSqRY90JxmkgwM3rjx0fxH7kyiYw+n1eBwaIieMuq
iH955Z+aAmb51VMiaONgsolKbkWefIycW4nL7jGWpyXr9ylByWggoRdvxhxiX8Y3OAaAF3IMc6rB
PkTpZmV2rceTH3Bn7OCZbhWIPkUihf5AmxsI5DayaEpj2fnb7bd8jz2t/PVO+3ZPO5DhfCatN7h8
OkhNRaRPtb43dGEJ21y4UeBsc5EVFtECahv88+SmJu3hXmfefUmGr3g5K3d3U0FtZdEJ1HGvJb96
rGcEidgly34t+a7Yx6LTZ26lKgug6Z0zQ6eSE/Xkml8zZR6G3uJlICtG3qEsi9WMUzFcBk6txF7W
sfbsbzWQhoRrswXKmX8951BA3CV5BH03r1WVd7r1MWllseN7u3Ivr/ahYlhfoSg9mRV1o44NJ28P
k6Sd80eTam8vIJJbrW/D+BnMf8hQRqkdM1btLYiQVKP0bNdufN0r6pbB/cRWUk2Cm6ElR5wN91mW
hkmTHZnp6rxacs+R3emG2mrXdJxswhPl87XDGUhkmqv3m4yOUJwPZWRs9ix9h8knmeK4W1btfZ9T
RbjFUlcU6FLqRNrevGPffIOqp26B8EF7wgfEiYqKjEFSJL6LR+/kSeSOmuQSjvrZ2zSdhwrhmd+I
IMOCcYzH3GbmfRhLJJm3emAt4u0FZ4MLTry4xHc5OKZbrOLA/s+Z4/0sjyOxm2CO1PQyUuIOrkaK
E6AYssdSRREfVGS7G3L13RBBmXkaZN+/bY0MIHYUmxJ3bpz/UfdUnCE8zdIRdsUko7i51gDYCOrW
sPjOtAD0nFZkLTD8L4UH20jKT/RC6ZCH/sB902oeAuLAHcWtKf7k9KgbpbmP0BXMcwrPnaIFPGwO
X4tgrxWAAnS3YwqBphnO3Bn2Ut0FeYT3TOYbm+Yrrz2WrbNLGRizQuXda04EuAYb7S2KvTWahMGX
NeUOyV/ug5ZfT+Tc/wNI9p8NIsU0z0i+tB72IRMlDRM4jZo2mZKv98fxG4JARLgUMUPrIgqHi9RO
aKlM+cXxHqLiV2TgI4mSkitkcfcluEPFOlE1qDvjYEr7l5Yr/siXTie+iGLljP6Vu1z+fpYsxLqU
7boygb43JpVSdNqIdEzAWNqxKC/O1Dbaj/ScCNpZAl0ZqfBYCVvkkALDzCLkCnFlj0VYuNmh0p0o
T69PmRSII9ak9cIrhjOyokoJZLQJ2ZMwqZk0fXSHGbMKa9HWqfrjgTXCrSWp0jVDbIbErE5hZkY2
BPGKkkb13Ppt5dXNB8Jjtm8Cifzju3pl8bmlM+jSPy70BjK1XnzLQY60AOfFDLKDXjCsTLnIox3y
TxbY+2a66N9oJWmA0TF1JCccl+08K22Szl68G0OwGic0QjpYRENp4pzLPLIMTRS7+pNAJEBrszEA
Ek7VEOEroEXJIy8VUUz7Y8spqFUVQUNF+eI2TtdPF7jP/YqdooMqf/80a35dN1arg5rbDBuPruf9
Q1+lSYuK70M6VFooBZhuuWUmf+dHT8xUYJ/g+JUoEMsFFm+AVcvQddNk1HwKECKPBFzpieGS/Jgu
8mY0aNBk5RA1GnZa8MQLQ2f9DpC7wdIQTT0Wj29MsqPXr9XKpMnasWCt5NeSyjJNRFTESMHQYFRv
iQM8LkgS1kkpp6ma/ZJLt2edzLV92kiIMkwgzghsFeXOV4M4OLkwxdvBgW1cYWtcUjjhJucdN8/G
JxTlnRxFMIcE9N7Pkuwp5STaQ40ob62bs55PymTcqHjL/zQazOHaEyo2WsVNBcqJt+ftASWy7uS2
BfpsfAYBT0L/9J/M6XTicqv4YfjvyoASWurXfqEKC/NEMx4ydBmvjmQTxElnTUymqbYXNovqMicn
bjfnXSn68HzrOMMc/SbyCBqXpc/xp+P73m6potGmnDP8tUXBqIAeupYvxfUuOneArr1504t3nS+F
UT0bXyRjc2Xb/u26MvWjq4RQc+6y9Gf1yCjXCBegDaQALZtmEMxzOgzcK9nXWpFh40QN84aiKNqV
EudHATedUd83W18ppTC7N8dKuQXo0bk4QpVfhTDKDY2Hz+ZH9d0CBm7nYGlMbG1+DDXlV5tUshjT
N3Xg8GM6MuQ7gph9Ucie8xdvdVj08OU3tIzp1r2cENrlTkKrrTDoKMYcP+T8fF5ph7evpGfkp1Ya
rmKh4DeSD6MiZ0k+ezgK9ZvjRziTkd0zeJPdS24WPgkWSRstGBDd9NAsICJcjIt6ZJcYY+D+/WCR
Pj/sWjkDEcdhwlUHdwCGAmgZONeFJ8oilg28fVpBU+aDEO1egjcYXZ3yhZzgz8sMzdQs3TcJYOGJ
UgGfG+1zWhQiHMFLjx31uW0ajCVA5/5uhm8mcP6eCD000VdxzB+4G9yT34uO/u8WCWOZGYvCjwCK
cYltpSiLBtfAZadZRTpmw7kdqb5dOeUTbr9E92O7TMondXkNcEEHyBhxypQk8lf6Tm3s54HbQiP3
9tM1Wop3KRuy0Fy2fujUzsFI29T8+1hRYE5CvQu8+7M/Zn1JMzOMnDZXZ5r+BFZverOwDup5lIxw
qOCRRYTWxNkLcjnMKZCeWVfXDHGugda6+7k8Y0ILPlnUtfpBqrYJyWBzqA+TPv+fw+2tID2dod5B
vqpa+6oRn0OFSvbjIAVx/qCNJuMd0qFQD/rTL9pE3t9AauUliRlSOK08YdVBRIYHgXor58HKr84l
y/5VBOLkjlKmJIfdDTbiLgglbYZQJRKBNn+6UqXANju07zooe7cp8x5eZJ1BfA+CskyZ4nJXIY1o
EhlO/zmX+qGT/JLQSvj5mqfwKwM4pIOwDlxFnUrAJu3mQ/AoWUMGx6DXma9JrOwl+OfujvXAbmCs
LMUtNmK/FVcm75y6ERaa0ZRNCZzieGwiLdxUXni+YKGU6UKKeyQRAEb1hrJR0Lrc1Sj/d6bREZBf
JkFf8aDcAVcrKuV6QT9So6dmfNIy+9V90OO2VpXbPyxcspVeJQGHDveSfFHXhzhh6qb7Z1fUZcSe
0qxI6c6VaxVFJQBkUMHv+WpEbnl8z+9aw2GwX7WnXjd03oE+1CqdQyDnqlQK1xaEsVJuKtBmLDRG
tkObZsyS2mKdpHBAE2MOMpNfp+8E2+qih1d4fEfuV5Fal9v+bbwniVfNoHYYVR0DDm39XsmhRq8t
wpYPoR+ROWYpV2iSh0BEQhitxXlEtwA8mx/4Jm3fyTzPkIQuv2lCcCAwYNafJf0nOG143Vrd7Q0h
5eJaySty45HA2B2RZlesx0Zz+hJL5mnwGhtdke93XP2kU40+OngFTLN+bDd5GEb3RshkWdIR0rj9
PRHBu989EDLP5Q/UHP3xbbbDPdeybt3mbElc7SAcbsDCM9snL8qQAJVBCny2jtRf200ZG4mHgw1t
rtoG5lHELK38LNpn7aILg7jTbwq7bpGoq2tVgyLqZiaYSHi5r0zc5ytUyybroByP6DbzhzdjHiSU
okaebqDtO3PGaySXEDHXGB0i6Rko5nye4/zrjoxVDGoPsSk/NBxJnrVNXiE6C6ZuCpZaFS4zzJhF
ViJlSQIaVwmre/Hdhf/BD67+y8NzigBatuXTvm/4whRyduN66vxy8spJYTLta1hI6fC6wSClIH1F
riUI3MbJWWcapvXVGruRkYcqEhJAnixhtKht1mdkJERwCVybjW4TZOQZIcqbsJuGbUb65d1kw/Fn
05UXDeQScxJ64KN0fsY1sxmSevkdH2bjoPtoPbwP8TQf7krkJw5+kEG3xh6zgORvnfSaNmDm42Ts
D1OrM05Gww3X+o2Q43Hdy7Gi9jivy9e+YbQp/KVNyzUrvKGwexT42dh1BvxrpHbk+3rz1zj2Wm/N
rNt6Ev/2wR4Dv/jsXuqTQkJ50Dve7uM2h+6H8Dsyv2OIekplDPD6BKIhqqjxXd46TPAdTkXzDceX
yjrlC8mWCI7oV8Enc527NalBWXCKt3Zw96M6EfNAZIHHuZ+hjuCTJrICN6pNrB/53Mz/UonAqcSG
eNBpvG3Gi1b+D3P/YK6wpFS4Z/45ayf6nKrkw6LqVOQyCY4pTvhB+o7v7ttna82CFCohUpFcUoBB
D8zjVCH2eb8iRo2FHzvsiHicxbsITqcpmkYzqk1544mb3OzePVb3J8cTxirSweNqoRFChF7KnAgd
L390U49Js7lL13g3n/uQ2dEq/Mo3yg7+gxmpdLNGrFCGT68N+xUXRujpobX4uTZJvzx5cFf4lR5D
A1isiTL3WAkLW03YtjVbgmJmnwQYRMju0GJEsoOurWP6ZpoaDvQwml1p29Yf5GWSwN2OXdD1xjmA
OSvyU/IkGgykeSqF6zi2sGIaCzFo1kfWR2B09ez0YfKltf+vOzNFk5itffpmt3k7vwna16o/PkAi
3RhrhaqqU/bduO4SUIm9BknwJSWdC7gwshXrUnKNyd308eEHx9P1Ed4I/8scIA+mxDNn2NRNP0vy
yYgSyw5UXVx2XL81aAAMVyRRQMqpQ2SdPxN77BuA2eUHHhOs6+XZ7G1AVJ2RcCWSTfyTsWqSH7Xf
jb7VOSk/Lu1mzHLURmbat93TzzWm+7SfAPKYcfjlbRsVL+1sEx+ARPOvtf2TFmqF8VIEu363zc9B
nRkwanH0sW3+dv+33ZY4skxqjCiYYI5WcUMInOVKdm7xWUTgQiSGfH3yGiN7F3GkCtxscYmxncIN
IiyVAsbB6A1gYAzU8sqq/MeEB+hjb7Gx+43aktc0hVtHx3kMlxZFQZRjsahPJlkZf7YDC0THmnfr
kZi+57pcpsO5YMVMcn1GQr1RncMzIXsXbHvlnXyCwI/0ElCqpQASID11XucQG/DN+PtBnTlVD4r8
8ex1039tzTKu7aVkxUoxkj2vBt8bF1OMFCRfaX9lezZvD8emL0WhzDpzBJ4vpaTbNpYiRPIycA92
9qEsB+QewFvVt/w6o1cdgq8ztmzTVwKMn/0uyjXQ+tKrfgLhNWYsC1l+rOH5z6oPjENHr3BUBHDK
BsUV+dcLGcIC5SmH5SA0bGPf372yQZvX0nmaRbMzZJqiNDQBvNQxvnBcu2tb4AK5+5nUMotm4zXb
v0nTUBw1cTN9BaZ+xZmjNAVy+vDhrEfrGmVPq2pNsV7QKJguasFuK7Wh9FKHBruFHBMUA2qnVKWd
2G4S5Y0MJ4/p+NsWUi3yDvaY3MUj37huJIV0iVRi8yJbfoyLCmgGU7Ju6AWRICBAGa05ohM4KWQN
owfEKz1QLLB3Zst7j8vj5pM6TFau3m07wE0whUCCrhR8skZmneL03pTbnyekyyUv4HeKRNCt+S0z
q3FM25v2B5Ox3OcppyfJl9heTxCmUwYDUSq4+RImmgAIW3uG0N/XMQ+hF91w1SQkIBvruEWzUvQf
WRV5Y0rQqPLmYDbaaIZPX88/YpGL6tvMBTRPDxkRXiGmZTG3qW5/fRiWO4flGbfvVqE4TQ7/l936
B9CJm/u8Qddt/IPd+OSjXXNtYRwFk+BdJIuE11Wb8BZg/N9HnWjoqiptpeOOzTp5NEq5WGiM276P
q7GvJnd2xttg4EmxLPTRnIkYOopIX4m8ZdkVhIzT0hkpmDPA3U2vJHO5M7P2zTHOxaCzi6Jm9Uii
AyNe4HPs+d3eHpyTR5TAmGNA76yMaaZ+Qup8l5VvIuVm6ti22QBTHTF49gKCnx9NSZkrO4czpo4C
EfKEe/0GyfP+U/+hD1ApDHsFxWUN1uCpzBRk5v9sdHnbuQOHLgQ8oIHr6OyEJA4YfFYBwI2QqT+8
mcoEq6BJnNb9je8hwThMFTm1x+0VbLVPvYb/1eXW1IVigt3aDXLZlLJomezd42BO+P0lmoLdShVD
fivgXEWYGdRhBHrDSQOc9F7p9CEmrd8HsMnxSgLjer+sSjT+Bhd9DDkuEMnHlPSW+3tOPSAqAEbP
YFRhkHUVb6ZbtO/ZOEHbFSoRjOdVIaG4k+7wiHhbWbLfeKsBwx5kkoJxdVKIgSF/9W1RvshA3gQU
N+NNS4iI6RALmBqxvRcPjplbVM5FWZ3bMxABVoUzGxQlyLmedu40L/qotyyCPjw4VTlXgDODjAsI
7A4YqsRSx/J0c0zhDuI504eUoFK0nlYMTmKQ3qjvaVn8NiSoL2Jt5iUeqKbFZIomy9HqefrD//rg
1z4keivcklVB1+r8u+KOdvPk5DofHr8RY0ywtFzcKXUiPDVcUTkcBnJYvmzWxh6kCMVZMMmwptu7
UVB2eSOf3DPrlfR2ne3OKUpTECVV1u4p2Sh7rK3lVzG8UwBFlGlhVIeyuplKCF0fqhfoUzSsSZUv
l08mrqE/u3CgMc7fNREvuc48z15qxtRkvqwmJjw5PZMCWfy8S+Zlld3WZP6uVc7bQ4dAVIvEurj2
fbwXqWKujYuCRmSiPJACzl20A9XXaw4KDotGFX4TtZt1sPrKzbcgZ01tlxYhZaXn0co4HpTFMVVd
u5frdDnohUaf7GrJdg2ofRy4mcxYQTcPgYrfyN0gGSrBcBUvKf5auBKLcLp0Kh7j4sRLv5PdU22A
cxtBys/XrLrqhxkU5c/QqAFxj5bOM5qC48tZe/VBcLW5tMGReegrnEJd17RS0pwdgsVX4mgfYx7D
POGY8Y82wMY7bYZa+EKwrogS5VjnuTAwKtIiIGOgFfxNOAWGPBixsCZSEelI1MScxXadFKYi+5Fp
8b7icNJNsb37bchABaf2ibsFas29vCPDw2Yhe03XTFhrcN08JxnraAy2WvCPfwAIxplR731oBRU0
GVym41J4ZU0VLUeK6L5rfxMe5tpu4rHMJFlFkkNvVlXFdclqzB87rsnEhwhHte/AhxcA+Uif+xjV
BsXpdCO7YazxmmhtVvBn1Haf1EmoNvcLCuGJREr0FuJ0Rp41QcEAshwsKzKHc9mU85IYhxCMbC9W
RNu9lc7qpDf/yRV5omokIwz7r0lxTM73QYUGmqmT7HxO260an9rweTQPIz/V7Zj+qf7XXHRqw1AS
YER7L0lq13wz9o69H7+7l//16xybusIwYkHP++WvAkfDKoMyBJKqeQlo+d1/hQxlrc8mmbw+gNEq
P7V7xAMPFJZAAR17hgtGZMaAWLTC5NVnD/g7TUvBbH7fTIcZOHIZYoFs/ByqdU2fV+4Mhb/FhaGD
EbGMmuswrSOwLRF5Znnsl/NnZ2cZ/PlOm2phFDmGs17+OA56WHYKWJ7l8v/6wd3J01HpyQw1PcLn
pUTIT0Ny9wtOGKgMZW6oKTwcpNT5MtCJzZ7t5nY+DohusqnEeYa3jdC4RqXfwVFWUhxt2yJJ8F5M
DnH+3zCUNTk1CybFFvR0OJL9fqsKddqT+0bbrWXa9/fDH82LcG8liS1yxdR6WMRS7ui0uv5jUb6L
Egd8oDkXNDS8vtLBzpxgujfYshYQ4fPEz2k92z0U9EQl/vucpCCkLszO3D1u6aBgCoxT57/fdE+p
0/KV+/cw834Dmr5NI3ZbCdxjxwxLdi1B36xo1/PpCuPUxMdGERwYYwacrI0PZeDCktu0EMqIiRed
mN5J/OxaEzvkYn5Y9sV2j5XIv1s2q4S5YKPskJJ3P0eTkj4ciyeKy/ppCqIX7e4f7GX4Gg7KXOyu
nJXS7c2cfB1qUGCcv0NaxZJeYoPxXBw2246l6wrmUE47oKnChn1VlxvZwiYYwq9yeW5qlJyEj9JD
nAzy4sUJnGNseYnCYpOs99TgdmZ8mp+3MZr+NhK98yIc8DpHwrANlQ8iM+Mi9q8gJtAd+cb/lYrt
ULWwpm0EFSX6arldO6DVXozYjHZuQXN030J9HUR9iVUJ/HwrGAfSVVb01/DuDmSlZyu6oR6S6JGv
HoHVxd4lEiHyHZ++6K8m+24QuTb/X2vLfp/LRREk0sdMqXLFiJVOVXGrvjrIut9Aiixpv/OzpVNH
mxS4cLVDOS7ff0LmHPwcKjdCSC4m0s8XW8w8Le6NJStboQ60+PDUnpcBzYySa8CwibZ4qOJVu+6z
Vn4mIRRCvFFopHvOZ6wTL+PxN6nGrP45VHBmuJeW+k66IcH9h+yr2QrcFznDlEqEfnE2J40ikOLj
YbdYBohUvNbL1u2ZLlo61b+J+VDLteXxW8SelV3nfvas1vNsCTd78TR8q79McFQ371UOsHTxFmCO
FOJAAphM3QnPvCF0KHpWQN8BavTLnem+l2lfrw4ncHlMGJIwjUt1qZZIIvyczQKr/Z4UHlqAD3xf
3lngXCU8YKlk10/RuybEcnCT/SkuondChw02md9VxYGKTUPMdH3xGmQfvDz79ulCQWgA8pRzUQtG
qfGOMK1aMK1G0et7JvxHEenPBDipbhGrSnLL8NIe8STVO6CYxr+GazN/lLqASVyrVmoNKDPECv0N
SrED7HeoZ/pasceHvSJT+mdAyjQPPyMUiL7h1WezjPBSlJbZaCBTqtxiX0/JCToOrGguEcO8LGm2
GFz4VKsyjv2FR39hSPjQkBW4iHerkPX8ZGcFGrbXuERdiDRgQixmZ0Djd+uwWLAgN2LDVsw6EPis
0cfuU7Uj3XsMCf3VXB1JFUESuT5o7rXEjh3sGSt4ityz+grr3IHa0YPiVXTjVsLgMYV50nTmqCHh
ywQPTi7eKKG8mn2axlVmKZWdjzh9diFtnkvyH1REHUCh3WbW7SuuNRtL5eGW4l00PwfKFtVYDtzW
SumxilNzxN3IKCgfFyishrh51uyVfTq0/rtPUU4Sb30MHL5gdozgxn32sEBOuYzR6tM1X2RID/11
Ub9RP+4PCRS0oyAN/nOoFpnJ+1X5MUbqMIask/ZzjuGybTKO6oJY4wog9iQslxC9eC99RXFgirlL
OrJ6FGvuKJyF8Fadw5XmIjM4pjb4snR8QqtmZDrxFWtCbC2h1I53o4EfduB61V+UBbL1WXKSi/JJ
BvSqfnvfVOGvCtfr1wLGe3iQpsgOVAbdrDcJKdM6/9TPb+fLGTDA3fEFaqLsTj3Aot6IGek58O/7
wlmPVwOKe/EcsgX3OW0tDJjQgh4heqYy+P0xjX89inMxBLQLzvehBI/DhzVlXWtZFRT2axxr704N
KTLjT3+6J8Ea7AZQyuYVV5KsD9B/6j9gK+eZtMNguBAA0+fWrJivmz5l/fnndIQXV2wdAp/Htm1B
TPgZzjjjGGmK2WhH5iynYxPHpNdsiuS+QqLZwslqxAxlITGyYln6nwSg6aNJe8xa0QiKtc7sA41u
t5wgRHILd6fbv8EiO5SVgDp9POlb3bSIZm1zg649zal32gH6JCu4CYlQD1VT9tJIB+iYwzr7EkSh
b+1mycybZQmFTvQZ//QJTYTYP9fHprFHMy4B0Cr1AS7xdYyDb8cJxWXh7d7Aav6zgjQBwfk5OuOD
KLfE7xdkbarq4MDT9DR3ta60iBumVhGd4bl00QhHrbJcI4zRazbcIv+l3E3TSBD5ZC2aWjRreRWi
2SvQf+ByjWmlU+CStubYtd/+Qt4fXhaB1EFC8b5irhE9n91KADDuSqvtJjeNg1l9WFPZZOEMXevI
B6U1Bki6nkDuLM/l1u8U0/djSW9ElWnxAcouUh5UMteGROfVaOSRHOJWKbhIgDgZp8XA5a34K8yq
415ztkbVStxdM2k4V/QFk4o3lLISPUpTZPDe9P8iqScFvaLRsR6zOrKuKecpy5WOc+hPxJYg4CI/
oNUg3ESFNbyWILPoYznPwCUeL2SQfcSSoQD8Fvn39eLsgOmCGQqfphLbFX7Ommd8MBsN2SnmWFlI
QJmDjD+KrK/ivZNMi6H+f7p7g7QwabetNN1eqs5letOl10pPTaS+Y+uf+q1edsYqQ41SEn4y8V3o
Y2Nn9/VItF+b8gZlS5135mEFvzYBrnBxkaokVMibXGUs5nPuWyAWsqtkfvNyLJBayziA1jvYc/tj
XTPSAEL1rYt6pvNSq7p0JaFPYTU93EoGXvVTUcsxpQCiliN9o7fppLg2BspFBe5DLNsLFpNMro3g
YnKopYFKgeJ2HeXXQ0bQt/uZ3FiuXfhzjgTQ+5YRlXJX2prQWDArF2WjWCpAb01vVXduqJL23R/G
CgaPyE3mszmS82LghDWa2zfakfEdH/M3wv/LaDpPTfS2p6m5YXQYUd4QgPSmBZi/dYBoK8sPdQJL
Hx3dHWItNIYU9O9lM3AdGyHQr0EdKaYDSq2c0SmyZp+sEfwNEpQrEeGjlCQS2BxZXCbDEMsrmtGg
l6ELRUFK45CJLfCdQWsHpHLSb7ggU6RACaVl03vMKGD9Dx0LGl4LFKEirRf+XoCgtWpzDuHG8NDL
q7whvfPHfAPPbKaevEaQHn1iFoedSC7jdarqY5NLqAexTuxGMWrPMgb4N5i3zgUYWpKaVApyeyAQ
yApsJdwHDa1Ffm1gP7K6HhWhcHZRcWEwVpqmsS1QYTNsrjXCjWJkHAhTG85ESNp8iNkG9GKBXpzJ
B/Ghk2T+pmA9/JHqAT292uS2gp1wY7qwZAaJxLgqd04tu9mLFMDKXAHHF3Uo7lsc5DkxW5NvrFij
41q+xo1Fpf9DalHYz+Q87sYKVACRv8T0gQZ801wCWdpAz52f3327ZTffE1Dbjoo7OusY77pw05xK
aEOcyDAeDmVaoQheGH9BYNFtKFkwDRygkfUyKZnRyZj4/aHXwYvbb/+LimzwZzzXwSjyFTXT5SG8
AaoCgFrc1IaBPbwGIab+w5wf8NkKFDaJ7lfPZbI8vNMgVE0I2unJvmvFZNDEuX253yR6s8ZRlTHw
jzwryRTbDNL4NOmkfWFdRox9YcMJMtKB/WKs0T0r3E3W0PT0gBwE13cA6CWYfC1Q6NrDvVqXWbjt
LFzjZ5YTtsgMxKdEv41p6ec5r6dPgZX1IGdzbgGbXFcMOcwuxf13zh0Ftl492gTFaIMFL8+ZQvC+
n/h54ppINdPQc3vBil9iFzLvqzJpbMmHb0fdCLMcQebJ26A004gQpbqhhE3YxJUM5JbBmUyl0BOY
VlJI7qWSuqjg20qzJS18ci58UePMsdxBn4qfJI6RXyZMqg2ivDUDaUkqSIMjD28wOyzWASaS9iEL
YPze8G0yYeh9NB7C6u5UzLLUrD0J4Pvb0iOtEZeLYwsV9WhKwmsjqidVZtF3Rhl0U5H4XtkyO14g
r+Una0jlDacnLhXwnf8DrO9VuoXJJ+fsl+vWC2Wb6BZb4/Wrsj5Aqy4fgeiuk+EJDfUjEF10Aw+H
eW+M0W/PpIKBijFrsFnf1H9PvYJzHvrvUlapRji0meKvzTvGFM63nNKhDXhjFOUl5lO8SQyo2dTj
WLfaD60AJlCL/YW/1ZvTKraMgO+G6GwhtVynEk0H4BxeVtClqQPwUhPPZTZecxxo+vBvX8d76nfT
yme+vl8HBWgJQjlio5uCvvcp2/7D7VdTS9PpAOGeWTKdlUGrRaqTmAITzqFM91RH7ji7k+tAI5J0
Ju4RpQqib4EsmSFAyF4JuEkpm5r308OtEnmkHMSSn2ZpyPjAMRqfuPnFAxtigNhzF5R4NNbEsgWs
LnZS5U4Wz9wQPVvKl/o9706OrHtorl6rhDJ0z1ThPsuY99iQNY7rUbAUUP+RuBKE8F18/zyCIJmS
QUjqV7Dp+JQYYlJyUDa3melatnwiPeUZwqb7jx0T3JnTXxggLInnokS/hsrCKWWd3F0vy3qqDdva
DcJnlUU8YqoqwQibVTAhJ/9ArpF6r6i0ZH4sAXyfPUlYIwYF1v8tBAseNq1tdnPaV9TLLbQacGPR
Kc/yWBLGjbc1cPa50gQbr5yJk7ynfdBtR/OGRfQ2GW48omsRSWyvr+SAwCC3hoWA612Fwbwtku4E
uNwFTDk1KzbxrnHkCZ5eCPf84JoOjNnth5qwaqo2h21GqTQSB5n4i/H5zMUsvSgXTJEJo+tr2v80
gY/Pj9gW9VbtG10RjTAcNgS+uS9kWO5AySQX5qsy3JRullmfc8vSqR1Eqdw9XlaYOT90085rXsVr
xy7of8a55GZN3XKpbWgBOWSzyL3zhbobrd71pajp97Vgj0IvrmctNBCFJr5WAEl+J9UzeuZM/iMv
wgiofCKrfBjgaYRSNT/w80SJSIldQAsNNUy0LPyZcYBt97+fJrDsPstZ4XSkSNEBFKQtYmUsPxqO
ssecRy9I0BDlfKv/QiBLHKIRTGekNCkPLL4wJSgj2bvOv1NS+s2GOJ9fS5R1KcAQjGpZNq0yQKPv
craBFhNNA9yuUqfw/AUjNLgMyDrFGhcXVQhsEb8AseSNT3+b+kbX9/oCQcUl+rbyBPfritW8zEf+
mPzMTFywesXwQPoCpMc39ZcHR+Hn6WmgLJbtburzuXHF76RcDlkFkQtOP11nkMIsX2Vza0fSYnog
ZoU6wzAX3Iz+7Pq8K8v9stBt7NkHaxiZSy+jytMRnqx6B/nQUDMwIIFeTPJAPYTQazOqmJpDGKND
9ksmbi0ozUaHwEiAB98htoxP7KziiQq32RgElpJOXMdI4/byt3GfgjVwexZgkfCCL3DVc/XGLZVj
tycvTgKfmH8pu88U3g2vbs0JBCCfxtIpjgLRZoQGD4wsgAxWqRgULfUzmFIr+GprIJRSWGFe8ytO
dfaejoQZShlvXAqTPNb8ckwwPolEsjubcFeDABYsA13uKEAJQargw3Mglo6BOgFywGVJ22WD2oeX
HVCmLchuMPiCvOHRUl/DyHvmYBb2hECXJNqP9CCLxzUyfZIcg48gTgXtwlaMQlX29S65dqupI+d8
ROSTnjz2LVZlr4RS+pE8TwzxbU7RnXe8XdJswJmJJysR7LuCzx2me9vDSRa85lT+9Q/jgK1FPTJs
KFASROrFjUnwrSiM/dNUslrackc5GY8lr/z6e3LuFy5okLQeTBwEthoN9LIEoJydCrKLc3P5c3aF
B1SZmNXNxhI4qQWjpH9w1gqEtp2jJIs8oBgEYjx7E3ygv8AJRsCGO7PFU3o749BxIPwr1fLfTyet
xxvWaN4ULZomNjwUXVr6gYO/f3M0KAOg6uAcdblsB6M3xuE+KNnY1M4CZm7sRg6pyMDQykuQ6wWw
lGJ8upnTstPMknHWNq7iEubM+A/1+mpVfQkyi8cwi0fc9dLCbqL7OuSPy1NejUWe2A/cIGJKI849
nJdKA5vRIL4qc5dZUlek6h3b6HHIqWZWGfFa8CYSVKfACIoDeVGsL2HNWlo9JToQVTcAxyyOUVzb
4FV6V+MHexjMdkbcWTGlTOqdmZqgkVTXYwBpUuAfLscGKz4T4jKYbs12PZ4B+fGqI3D8/NSCZo+F
1UMGGo7Iimk87EF9vHP8m66Qo0DvkAHvDZ8+TRB18VOoP0gGztTX5k42KLkm9KNvYfCehzw0x2zp
QWyKEYYel3/nh3RYkINyFxVofCiC4S7FMac3t3Ks/hF+WazH0JMGVnxkfNa4m5GGq6pwV9zEZu0j
U9OymUQyzGjvkjoNwOGIkuYyR4dN5xswwyVCnObrFWmg5aU4Xqfn8k6aQgIGJ1pDQR8eRhqLw3K8
ldF51OsFZg00MdPOq9sMsjzw3uS55Kf3Lw34lrU1D9F27StpwGG5274Z+vup8dK04n2Xy0RcUYGo
k2EYjPi4AxELG5/1WBbcGNxw3vKipK6udF9XLftNdDcAZLKOqhXnHPMFUzKK0uY6CAuPPxcuaifW
2wpbYp76J/TtvuaOsnU8JnJZwG5CY0ZYyzNY1Cp6vCN78S7YoRPdtiz/csjPaMIODJB6Oo7wkkI9
zNNwqa3pEbs46CMzTG382CydI5XtRZZakb6lhwFjfjcyO/8geCXLnA/aXAPhUcoc1B5Q4obEhdrd
kZfGbrxr7/zBks4h+z40YSuf3Hai2VN5VqU7GSFSlr4L4MZnUVT+BNaxGLLwXt75ZV32KW/FOGxN
pgU1+P2G4lGB215wf4gzbNc6CynCVUbDgeqFCRdUj22snu9V1w8wMraQoiI0kAZKzZT+VncN7a07
b8YAcHATIRZshVQTEvc3MaMVvj48o4I1MgKrh++2CRwjRZtyY1rdXt8O4estooyAJJ75jgwEFum8
UlwlnUaalwtS+FSI+sA21NzLjQ7IRloze8YL9qgNMVPMCMMC5iVK7PB13PbYZKWUDulc/YYAQk+J
eiuZtMZ/g0q9wm3cRcNUf/T7zc4hjtgOglYF05DX0taXkPFxm7acNuD1Fne7iQderPvSONIxEsyG
kM19XGzhklF4ImCmAa7TdCW5X+cINDsCGCwzNBsbbGCFz7BRXjV3RA1NCaAHCH7Ldai69+yKRluB
JIDOZoMb8RIKlmrMAJvTI+yxr+1tfTxYqWqADNDtpX1RbkEiRAPpbHbZl6M0/lpacXEVBjCasarC
lE6dxJH6pLdVdah4hoR1TPbNHkBR4b080v5BjZg6avriioxRuhr7Ho2pYGHMkGPhpXh7RWrsuUmQ
tLj3phUFE6lglNAXeHblCgjd3SA5onJwqHjBdfllJqDbmNnN1TnxUGUHPZOUKqtepPuP+7CuLQ2i
pVd0swQS39NGLu+1Ir1jkT1QqmaM8fAj5e9/+mPFXOK3xYPMcUM2Sz0Uznl1fHqUBSbdAoR0tkfn
xXDCR0z+fDk1inGsIoTGQpH6IBy5rOmC5196K9LruRy55jxjn4p3GCzUmhVV/dMmAocmUDSf/yuQ
NxJ58burPT4NggmaW6gupSPRJLmgIAMp5kql8o8rXkzpvM3uK1v/fuFF2VUd3ZzjBaCw7yqoQlOg
Sb8xCGhDjimID397QF+yVdrfmsMHJyRAwk525KzJmc5k+OYaVXyZ4DYlvScO+3x2Cpgy7vBaVdo3
zcQNgn3FkrYh3NuWqqsBqruAUuo79SxCU1CY3ldVfjKMwBiAcMcke4LJzpi5UvbXSwj3EpfPwNM+
UpkfEN4cTKSF3taFdlBnjs3w0Wvud4+y757a1j6/OcLW5Kkd1vxOvfIdcBkQ/HgZuocZae+45C9W
6PDOD/kBT1QsW4szQ8eUiDy4G/vyCzZ15701ow2USXCFHQxBvWl+YC4k4QH/MGLannjxHW3m2T4+
HsCXCOGahCxXf6l0dpqijQVuMPFRpajiHssKdH8LAoJBJ2aiNIvws5ybzDPRS3hJJn8wZzFJx9S+
rLBTMQonTnAiMkpTe8PkhkPnZxRR0/9A0zR+lwHo+q5HeBgw/4zThAqsIMXUDSexmc4+n/rfsJ6j
E9X1ao1lDSbbCiTWxB+lbLX550Ns0GiLKtbkDqrLQByea+KXlQ3kkhSjc+gGu3j3dXZ71nPA71jm
MADNThcAbYRv/6OG/EHRHb1+VHS5pM2Rcx93wBOFfXN0k4izAhOqkHjVFwp7C8Ck6+n99lJVMjKi
4TmGO2bgU1+NT2GntYJT7/UVwlygkPW0U235RX8WGL2+U7sMCmZquVBNv68ILvP9DyAXZUdq6Gle
ZrSo4ZBncTxN3rVF3ct0m2GTzhoK0nYel7PkgaYooVLKJafNYbgKK1cJoGBPtUl18u+QvwVL5Ttx
+oF+r8yvWTbXbtK76lU8z2IoCHhIOEVadGrGWjFVu+9nR2vg/hPv/aPVGK0aAjuJr8kFobg+7h0X
DpLb0yTypwM70qegG3ELhmekXIexCEr1PF7jxU9/2XGtRC6jhWwfjOGHSOn1l++rZis0vhY/JcW7
Gr52Swx9/2tmlGzM6RiMGojA1skkyopK/mR5vBTqyRJq33JYWyTVXcMykkwNj5HiyldLwV48JMT6
fVCU9uIXovDTOA/DZwTbN7+jJV/i937n8NuA6spu3iNd/dpOvh+p02ON/Oc0lFYA9x+uq9xQrFTk
bq3j1qhrdBsEkG9QYXIWelY634mOlCQZN0U0CUNV6iphMrtXdBklc6AlxLkI+QfZ6SlRuEcUE68k
Pd6O/FVYDqyLwJlF61SZztExggWaM72azSPaaAViDrRGImj2GguDiQOqGwxQtSQgr47jXsEfunSM
EH74I2Go7i+nXoZYMoWKlvNZn1NWYwaSSYbmCVosZ35UBCnUBIg+M341Mkq7ifimr4E+tEUf0hSG
PU7iqZbOPp9TjG9grg++SXth4nNbEVl1qEZCcPss4zP4quZx5eykpSRxZhkZIKBhG/j+uhpWQQac
SUOh0OpByh5CgCjjZfnBy8Vn0v3+GcKylk9exKonQ40/2wzFxesyZWCK93xajDyJOxNWotwtsMuX
fmrOZTjjldwrSRCVpjGiINH/JPnF+zzLpXMALbH6H14YnzK5OSmcdJGnQkBIFEtpg/fq1Dzw4Una
cHGm0700tKmupqjA6f9NhiBSl3yK933fPqFIaqlqpMHW6capbbsdO1HmwwFMKK2Tvt6yw4wGsIkQ
Ztalf435ZQgyXB64amAK3q4jVRXnuQPwvJPUkeyrZ8f6k9ypzQ8USGaQtv58T6+uKNNoR0kOisWb
CThxMiqbJG0LnAyRPnSRT1I8WmRT6l2DWMom3x1yzUwWb7wYH2IgIUsuaBtXyBcR7Xm2Ms3Nb1Qw
BH26a55/wgvSx4KOabPz0BUtz2a+TEEX9TZuWASxmPYjqtNtARvbvcLVYcs/c02zSsPyJ0Vro1z+
Nkw2PgfsAavTXs5u4M20JGyx+NbdHibK0ts+LiKEg+SDZVW1YkMkulJ481ESEUpcIuICNs5IhY5W
/AI9ySfvXsMVvUrrfkXdz3f72gSB/rfZCdVOPIphjcuAL3O0tbtIj1HOvCOSpbunMybWiBvqZNrS
04Ex74L8SSZ40OQZCXSy4I4Lh+yN3eAIUBYaXp9mJSFIe0zvtM7NDw69LiEudrGZOEbxsmzEGff/
butOruriucd5/RGHI34q1Njyk+e7rQc87bbVNPmoCYGWeqIbVLc1Uu3kf9wLRLQ54VmwKDrT5Zq+
j0euO9S8fhEfGvTp0E+Pug/hz2O62zzMq98JsnOUWt0l4uvI37aw7cBeXsxcakKe3IoqzJpjCbnm
G8cxXh0WD79dzxnwGK91RFE3nuGZ7sBc091eeeV0P4x0T1bSXKELAzL8XO0yZPcujNJ1T5INJiFB
i+ya+iD3/PSmf1t82k6wmJuoOaArAAZp6oWdefuiPEHlyitAtG8Y3vjwFWBYY715UKfBmts5STr1
imevSo34+RRvcgK7FQ1IeDuOTTHe4Fw+MU6HmXYGiBeVFUrYmeUsJ7ciT+bn6DlqKtlKbqosbKHg
UJle3GZvyYwLQTyS6oZgXS+a0QZvQ3yIreEd4FQ/vr1L7fIWpBeCkmPTKQTYc9raQCp8QdnPCn8T
8cbDzL7IZpmgaYOHfp22SjZTIiMIUfQnm9Doo/x3K9qz1j+Do1cTSUeQw3KS5Au/mr0Zxatf6iyv
MWBExf/KTLkVs7YWrWuQSUVTR4z/WPoeFSboywQ5jxYqTGWKfTtyaqPeEDgQqEDMZMlKkZ1REHUe
q4wa8s6hANGSdQJ/Yrbcj1bQ0aJbUIGNHj8/NxFyzewUN229d/o5nxXXJ+ifY4vjZ/APqqIpq53k
yBzwcZx+FWd2Z5KnkJWOmxJy/wa0MlgS6qjpBXRhbabfpjtj5JNH2dHgJTXCYPJyNuFdQohRuMvr
QXOIEtf167CkF+DwQNplvFRa3eXNekToqQtWDQA1KluF+kAoiCKrV1A6V8OUgJ4K0ubrJ+DdlWDk
cq6ITaUq8+paurS+6flyFhnkeCcMLqKBLsrcd+ShMNjFKOGPOl9V2p/QQeBFtsP1uEXa38rnklVr
SLLWKE5lWXCM2yLVA9rRc1HGF/VJJ+1rdtKCGMNQgmeSPmFwnrL/XBzIux5ILDgrjufS/aAhfBV5
wMcFHU2MA/LHmtsFDcWulzGCFCZMqtDxVnjWasgI9v+ov1KjgDgRApaeRL/JhbWy2S7xiDoli0Ts
PFZ7k14bjXGko/lJsRlgmyyUPVwJQ8B/Oo1c1519YBMCK3bJv93FNSUG3y7TX4hiS0dtCWxoi9wn
UfonK1hpk9y3NXBnj3RWvgPAsi3qBBorXhdTM6PMhUSmc5NILZkTWHyo6HiMr5GZk8JysvDuktmv
0ezUCgrj0svkrqbIw/htYNXEXBsZH+tzJ3TMOMKKLqT+Q026FBjclF5d8QloOC4CIaj8hd3dgqk5
nrpknpZFAfbUFlIW6sa3XzrXr6lAaNJbMBN+qkJGqy321LVBxZN4lGT2TMxOqyZa+yn/VulNw4IB
r7NLo/6OftnKzFIgsW5UlGDxh/W/5hhsR9J7Tqg6DpmwCqzSy+PnLlzTQf2W4/wuUtXzj8/4RKv7
oXbUohmBhemD/J/OHByVh5UuT83Khv8oheNmVUcz432laz8XRYo3OBvbMxWAOkW8FrZ4NiCsqLWR
8c96QxADJO1vDLl4GsssTakFhPJlzwgdJNLk8BlEHfpz4f4rd92HW5qjZSkhqlmtSipjntZtoh/r
0M8uRWe7tNSG6PRV7Yg7peLZptty9k4gJ8IG2mR4b60iKdmL7d2SYzvAFPxYFIEqLGUjSgz8iDTH
wM/pc97IOxneHkA4YzMWOd1WLgjAPqxOysEgTEtOwrPVjNn6/kBLV++9WHoRYrwjolVmmlQzypVU
p3e0ceynKlFO0XCkEuP1x5a//D4asnWfMBeZOuxUfCF28gTWJUTE9v9c3kGtiksMA54hexh/ULhj
e1ANtD2u4O4cujHAlUvUCPk72L+ti863Q/DnH88FxwtLs1DKINu1NK8TLdAkzM4jJ3TOJyVxXoqk
Kc/CD1qSjjvX0K98m2AmP7fHbzYRcq0reVwGo6igmB/hr7rF3qw8QPgFYoZb4BZRY3Uru17tkcc4
CDXGkACLqHi4bwD70ZkVztTfGDgFAGWUT+z8AaS0mOZUYFfk53BRA8oAeFg815GRR0xvAoXXI8XW
JS904DKt9oXrjdBMTZ2m0p69fQe3biqt2kxxQXZJ3LX7ZnID4CHgNWM2hXqLBNSf5vg6xyd/cUEp
EgxwqnrRZHNjo2Gkih4UexPFxsHkxHa7oCK1zZi0tp2s+0EkqiTUirT0vmLQKWaYt2Kss3SAZazy
rN6mSrvDxX04UQa3EebfpPjjy1ODAnie29BCwxPuKNei29jBRJO1taHNvqlEZE1AFtLFpR+VNx0R
j0/5F5mhGom6BwGX+hnLEgChmyfss3ZhGqO2DdotKdtkTtv7WLTsaow/PO2BD4K8k1AHJ98iSyYH
C9R8Gu/nzVFlnQRQM/TjdI6TQeRY9G2KBgTxzHBAiTVV2QL6hSgxdG+h49RWltjmVlZTbAXnz5BP
Sd10tXXu2TRJrEEUsUtm0jfcGJ9wPBNH4sRvXss4y2v+VM+FioROsA6jXE2KTYtndLXNprInZeC4
aSf/s+e6qxRt9vZ+EqR9JyINW0pgA3c8y+fqKAQom4iZ1kXavmbn28cGG62sI0+/+Afa0WH9r6kT
zKPo2jMG0Kqp2BDJ0o5NxZ/YlyPybGhreVuAe4bRlTPMcb2Ycl3Z4odIi1u7WDGqAKEt4cZTD5Pm
xo+rzkO1gHx4989sAjC+WwQRY5Kgt/xYK/rAtNfbBiccLcHpdNR9CG7nZU+NsfrwOLe06GIBvyIC
xgZ8v8y736n7Nv7S1RRWPTwr4JSVB7g09t5S+SDVao+Q+nWeHvkhaLh0stfXG6VHmhmXRvs14iHN
GaIiaIEimfYWfK5zcBjJSWgRaal3FRww+mwCLHDEQ6zlwK3OgF87iNrUQVdwYJiMDC7/isJ4/of5
dL/fTldTHo6acE5fc2rGX8auRKRe2lp2Dx15Bb6I4J/xNSjTwr7dhCZxfRPe8nSUagXJq8Ss+1C+
QYrwaC6AZPjV9w+bNUfcccuujYdGOArN3+gN+ovaOJCBEuJa0KpJ1zV2TbIwyqVjX427HuLejFhH
ga2oEUEkUN23tXUN3y8vbv9J/i7u7GTYQQa60ZQrSTnol8JXxYLIrSwKQ10TfJFDKRZNjr52LRKx
puSUDrw13chEwIwblaaFdCK8wo9vX27QoF8dVdam0HC9/3Nr64W4Tl+iM6RhMYvHR3Vh50wAB/4R
uxctNzTjMMwli5qHw60ozD3XWeTKuMZdvecIltkBH/xHATWVk4GJ5EGHZNyNUB0MZMxDXhPbxbvi
LZQsQamI/jbV3cj/mTdP/F81b0DIEagdKgyszNHrVao5Q0RpF1qvcFq7YKAqHAky+uiaY4dUU/+U
9d3crKvf8qU2kerAuxvcw2YwqZjpju/8dWzgBJflDOq8/86gzQpQYRpw/J6ZNwl6dKNgHrsRcPfB
FaXdYmmaAnwZj0IGhafoXcL40Tznm64WCPepeqCFN6rHjxTbwFRGuh+/KObIZwTFhY96DH5jl0DK
2190CTV2JizPwIkqb9WeIfURuAlTiX5a97YVGzWmoZd0RobxqIA9wUmnTbmbzWhLI5oSS2YhWA5E
B6MjCbtQyn/jV3Z4PAREOL1wkg7nHRyXuoFN3i+poPScm91K69cIEyv9zyTNtopSfeB5cbvJpcOB
yIyWQWjiL5jZXCxqAZGKCkPnQiiBFzDDAC7ntIJPJashZasfv/qQIWkz++kT7jsp1JoKGlk00vpD
GBW5dNegCCKFH6ppGf5VDoEdKLdAjhm9l98sX5tbC2Nyu7VW1tyB6mvHbDN53ZKRKYWs9Yb7L0YI
00z6n5y8wL8sIenUSTl0P7OsxE8Fy9VsdiJ7SYjk24HPivr7jTCS9kMnd8GhHu3kESrkye7k/sKJ
dMQebvf6968O5f1Ai3Seu+kWlYP5Z6kvWGBkLLb3z0a5RxQoxxMvM9EOfeOCiTthaqiT9D5pjDDZ
w4UXJS9DaZxYS2u+8nTYOaN742t0Pah+apmi0Letze3RT9OM6lbyUZYOoRwADEL/MSEVzvYNWh7i
JVyKPrqtb4YaFr86rTyHem6xgxNj7hwqu++6wSMpmyn4PCTX+lQHfY0xfmjpFTWYtfu3tG7MrAP3
7DCrfcJDCK16XeIYBnRO/sD/aTY5+Dyx6A3tcdJhMyUTSq4Xfrc+D6QaUwv5Vkj3JWWUV8GpKVzv
joGllP8zMsP5hoVYXJ87sP+karA60jrgaddbvJiqaaO2DvUbSkSyq/LqYX8hTuMv+kTiUVgT93fL
y4CNjWV8qr5jf3XR/bRa48B2JfLb6z5AqXZKMIAjteZzadsnBlbQWDdjDRb2DWB33kCoZ7YP5J9H
Ho9bgEzOYC25KQKAybjIIJ2dOQmPUssjeC7gUHRxXgtnuFOiL/ytMDCsUXlBA1bs7MI7xA7qXMp4
w93kUwVs8b9lrTpkWj9a2Fzsk9ifIIhTt6krtR7pfcXk4VdjKKoLjjAsuIKmFsKges9pzIoHtr7N
YcXTtNrumTCr4FeSPuTyy02bkilmb7dOCULCtPhQnJj8l1Fjn0rTMbcfn0xDsaY9rRUTqR2bTuRq
/ziwMCzu8z/UZgPCidfhkYhQtzSwzT8JhNTV2c6i8Vf8QxrNEIBMBw8zNZIuVO00bY3X6ZnHkIXJ
lE50zFFPELG3fYhusZz6wHZA8/0s8R5KSC68jdPZm8qSVQTd4f2KXLFi29g/KKuxWMPu3G06iz5y
abWfCesCsweTS5r1tl/QFMB7bKkJYF73DviK1+uD2iGklBkxVYh5m56bBMcGqQIYfmuriyvflssC
Cyg4gUSo+qd/0z6Bt0Qj9eTTvmhpmSfltsajjEXuM59UhrBoywHqX9LHDf5+K19Z6j0ZehganVSP
GrtunknOKaJ7L14jhC1cNZVTn39ZoWbTOBf6CTkCoBMGrted7u94h/Zhd4F+NFwdqIkBbx2CBRPV
Ql7PBCyhrE/9ilPXrj4b4UqOwOXROGESCvsn6iswIYmboWLRbJHVR2XELxfc2V1PIsKkP09SQhoc
wq81YWcZV2HKkNFXlqqBUFqv/IFapSqBXfVG/2f+v1sRZB+c4coXsd2L8s4V27JNWhLBZUTOCpOl
CleGy21f6Ayh++g3qqIZs7D2Z/wECO7+iXKaR9K1vZEZzbN2KL8BDmAJLGgan8tU4jKMtIGY9lDU
qh3TlxmAKnQ5y7eOoBgU2HVJFd5DI4dO6HJq5Mfa4YrvOUO3vSTb96rcvA6Q6E9sdp0/LK/Xox0M
LXPs0IV1c5VFeDG78NuOzR8hAVImAbf1kbkdiIjNju8ud4O8VAv7UIUE6SZbFc+iwio+2gT+h2GP
zH4B72/fdCzHnthqlR4FTau6BeIhBgkR7EyTufn9cwGYJ7Bftg0/DIuKbKGjQWVeNG/HhNKHUwaT
Y2dkKyZ0SFZyGlcHazLn9eR/dACbqvp/TKMkhsfxJSmmnF7T+ObMjriKCZg06gLi7/9acM/Duepv
Q06lX+eQAx5bKQTyOnVxt4QMKQrxY7qprzx/UVCNrbchYlOx7Zd+cAMeRVhMedKNAsNpU+lXD5j3
AfHqP9j381tHvMyGGP2BbxALBjZKQj7bccBCk2dOXfyftoxLT9iZ7j3mS3HOLu8sn4FP/B3TvNlt
RX3lCB990TlaWDJ2SHZinfDtfkpXMAO4gmuXLkwtSDm48KEKpj6ZfR6eBMJA+y6AtJKnyXyoIw7Y
oSnbLG5fkrp0Cdgs3yf0z6nVWS1WsjkhP6PPF55MEtEcS3aVAerxVPvQ6cxrZzkS2uovLF6d2ox9
4vdidnZuwQKfQe0lrrLJAQd/8oMSCMnLl98xgz0vo5HValEfkJ2XOYVK/HCXVU2GtfZE4/K/3cJR
Ehnxz6Y3WxHtohyLHRzlmjPUzqtEnFJato5cgZfrdjqT2EVcTCyynBbXpPSob7OI/Rp0xb22mTih
axh3hpdfDZAmAaO777FfadObBBo33U6ObnEG2xd3kHp8/W/Dt3drZ3vE0uUMGTX6nFE0vMntNHL9
BpyefzMM7dAI7iugLZ/lor5Sl8DKUj0ON9BgVyO+XPAvRydE3BitluahiYhdN6Pr8remNqVmyHYO
q8uE9HgQKxHTnhdiAjRpKQ+CuaewLmIu71u5TmIu5SdIG4YLbu6ISHZhkTW8/KABh5OyPHylQat+
fBsifzYw1aSM9mZ7wJuOrPva/3JZ/uDEwcDrUsDs4/MZgCx39+dEDDVkwtehVR7ghitYn4pCrGON
gVDEx4QRTpt3iNc8m+AzSyT8NeJ5fVG3oSAdgDcEYl6f3eZeZu6a7SfxkMfisgioy+LqzxU+2gs2
szb20eRaA22ZV8XdbLQ8AQ/FvnBH+CnX7436YgGyK53cYSf+XtEB3kY1CDvQI35K5z0AzvUq3PI9
XA2mOMa2bDwA3NEJ7N+TO0KVl93Ho47oVcYYFU/EeB/5TXcrrT5VNBmq6C7uvPiMQYZvHPXAI2+I
zwMM30wxZVesenkPccRZJjZZvuazJo8HLIWis8Nnj43E/VlomEazX1GVxF97VPAzNgDBoOomKhiq
MVHk2AhJD8hKKus9D6IA/hDiFcYmcUIE340OpEhKx+dr4BHCpzfMImvj/N0DpbjuabU4g942T5l7
AL48I9Z0seJw+HHYGOI6jOUHxhIN3rgENqnT/BWLgZVmtaR/ExwBykFOTwWexr/zGEujwjdJ/EFR
EvghGE0jjFIMzcEEhztFroa4M/QbnM5AnkOmZ2sriKOEGZrAAEqnX/8qZBy5SEZg9Kc82nb2NkYb
leYtO/hED5+M4dyKcrQs8BUVZoRunC26IlUAZD+FnYXQxU2Dwx4Ge71YyuNCmeOXpIkb7ge82A77
areuuMREoyt8ZZ4r0O9mz6O8WX3JLsXl4PFNVTzECe8OVaRpua+TBK3o4cslnO41tPIBACp+/msz
xaAdihfYHVBumZ0blnVeQEhE4gTZGSDGA/eRzL9tNe+57vlod9ecty9CB4MMBsC2V03OpdiyEIaI
stoqsTaVr2Kv4Vs5HOhBBIHK91dVCflGe83poRgVgaGgFRlhvNUl1VQBLaxXGtlnfbaMYMsJFJvl
dFHS8Dyprsd6ifPyIp7uAFrFG7/S+bHk1em7mCyhnNcdia8LFITZSvEW9bZ0lymUTHwoQh1f6RvT
xGSAGY4rNOWXRCc52j7wNismVnDT2p8ZKTOHK/pqyOefLSIqzF7FirIWqAY9r+T1zNxD69h7XIFp
gSbgeSM5Zom9hcWnnEFPPla347mTfPFMjzwNhuQweOnRS5mQuGvZhy/sMeJ2Eid8eo9h+Yy5dmGC
A/qsnFC09yD3pPEgNg/Frf3QMnyxK2tWPMKyFZLlkiwRMGqCCBZc3G1Tytg6ez9YkFzr4B3ejllL
p52Z+4uXtkjB0JdbCoAmS4nbyQvZXKqgqgXO0GPVychGz4GAWApFdl7lNcyaCWmYt2iY75rn1BFd
B3UaEOHxK1FLV/ggUPl+otWDBm2OCtuu22cARI2ILM8g1+IgNpHue3LIJdJkkMSLLsJaebSqxYDJ
khAX7Maeg53ePucK/qtwB4oYqMLAbw+cuzWRe+g8ZtT+UVcJZHov2UOQ9cs2APrNYi3XLoojzat9
aVreNIoEo9AjhZGsS9DJddyttU9GiG502WMZKt7gct0g0diAOEYlIoR5Ge058TRPl0Dqs+kz4oQ5
7u1FX6DlnCzbNjgStdL4VmyTjMoQKOKAN8OEloOptie3WqwnB1miipT1i6qh5KhwKwTtV0s0hV0b
LZ4EzhdJc/ChF2x9Knm32Y1wBaBvBQx741Qpi887HSRzSD1Is2jgr8eMoa+okRw80Hb6GIv0mXZR
jmjVHouiAvSj5l+ROXvaV9466wcPiZnubC7lRHLIVYu7PC5hL28KM0U5lUF7OjTkZN2+/JM/J+ex
8nlenQ5p0oN8brOo4IJV14/NQpVAvoQhGXjVtTPOYZ80oTYBsx1gpIygiZPTQuOKn8Q/PNtuO7zM
459l+45FPHruzDehZAepzj1QIcTd5YlL5MzBmgZEquUtoV8xYkq6b5WIsdg/mVkmryacNZnuOTRH
D8O0cecy9dUCkJtQXp7AISXO4zOwDhPpGNcFlSs89HS9iJk62vqbsGQCzrDbFEjRZhKJEr0+zMQb
81L2uIw8Xv6U33r6CJckxRmDUEBNz8Bsu4jAawLF9gvOPjM9QQNghRr6sx6QRrPtThc4OPn3OjHb
WZUKF6S8HbAT3zT+/YIwSU+Jcz3fIVx0A2SsGJJeSqM8FI1l8NDhPaYrxnolxTFs+hadiQRVaMax
A0eRAERHpoOlQiqmcqoSBYkKaSCoJtIvj4SddiSA5teWeQSiI19yJetKJmfhOKZ4hayjmKGT1kIf
tLUFhivzr0Bxq8K6bBwl+AIdQFMcqJiQ8pLTF3S6T8uYkeLrKvI4Ml0AbfqyOyCUSrCJnbiUBSNf
RkFP00txrnXGFpGHhVzuJldzDUd+dDPYXmCp+jYQ18QajUVqlCtNqgwngWx0DalCF5Q/6cPW/oIU
6Jns/+34GYQnZSJUxudwEGT8+yaeaKINVmoCAYpAswNna9W3nFBTvDj0jgvvVJksZqUL9Krew26T
4pcFoxZlWVHQBdkpucGdBPhGZgJEV8tteEI6s0yS/W1SLkfgNBunhdYVZ8BMIxw2V3gRX8RQHbRG
94mFvI5R6MQM63VqtuopT0TvgrDZIvqyuBmL1/R2w4KvwwxXZXg4GggaT6grswV1hak8f916leDP
9YcI2tVJQgMBTVVmiqp1uYpCNCcWRPFxX8+xAqNo5UpZM6jRPTH7j/0DQ2U/lO+ilT+rRmGqeE4x
+o7x5hp6fd8tvyqKk4YbI4JMj/T88Urc7ziohUDcXvqHAD+OW/GfJXU0bxlvUGIt5n8pNJUgIqTj
ZO47JiYw1bAlNyPRMkAuKoSj+LwT3GJ4Tb7jPyAl0+z94Od+mRCARllMHMadBOpMONFT8vSezd38
23r4yuRjmeM9+yXnFeHFAfvmgbb9w1sItnPV1vfUe1ak/nyP+lBEh30WNWGFx5hr48vWp3dKtX2J
thM2ajctTf1ryar8Nqc+Ipz2fY7PZ6djL5C4I2hFFg1AaTB2pDT+4RWwcr397VJBb/bTXul3PvA0
yf37EbhcqzS2uL61ZAe9aTRzivnXJ7uKnSJhpVKqkYAAhMw/ABhdRIwvlclYqf2ZDHI853OFwZRy
Ar8E25zdnAwS+SRPw8kdYAC3jlqZsAOWFw+zfwDe5KgT5FrlIbpQmIGvb+OzMuJAzq03mikaJWPd
gqRDQhfCd8OAcfLvGfirlJE3LMjbsGrbue4IQ1ouhdcUyXkSry3smj5zQY4b4NR/Vvaa3Hpi0Hcw
bSdsb9Y9WD0WXaiHp2vR5bMDJRVboVmQ9ZzzZe4KO13mFWUclxaY1hOZiYGyBeHNQylP+ZLoL8ln
pmRUv2k6DxMA32jw1uGYM4s4KgE1mM+iQ4UEGav9yUUjQ94X7110RQQnMVGCfW/CPvgh1Ce9/pHR
v/hBOTBvRKR1kVzi2xP0SlROoteYQU8MCcIW1Mvz8SLEaW/0PV2g7drl6KSLPawrzXk0+UK+nVmz
8jRqAMDpt+YfPB23w4LRnVGLPAC7ATj2r/ugdSfH3/GTEEIFplhA8pKKJs0YhrgE4Kafd3tWh8PK
nkJaDta0r8ltvUA5nbtFTNIaLeS3sgBHVKualfzYGAHpd8s1OfhKiTp44+S0zagDC4bzt5+8VJhH
7ktu4OgitoC6kb3d+jlHiT+Vl0O99oDECLj6sAPWb0qVJ/Yvb6TAFZUFOuoAkOTrgSnFxMXAe5aF
pySc9mcJs2ghQrzJrWIalaOmFu9btNZE7KRpvZchmsWByoNjDKx7kxlc6edJ92UQRGPbOxr5G6db
JfQJHnXyU5y+ZC9hoqjdDUzJSYKtw5goN9CdNb9K4jsw6Tah4yv4NCVAWLSboyUNcYGni1bH4BM0
fcb0sUYIe09QuUs9/7w4gBr6qKI1bhOHokz8YxOkL+CvLQDfr0Qu6ZJEcmpkqDyXIR/g/dLZg4fx
rHE41lG5OFBHYwujdx3fatKpfJiU4/eI8ZiAA15UbmItvGhDtxjPes/6P+NLoVb4SffDpAy4C9XJ
QMhJIMDKI9mmCU0dcEv44S3Eio9h+tyxpn1Q43lHYXTAb4JmeW3NYQv9SeJFGXYkFg5LHZ1WQpJH
PRvEMGUn0QbM7gPvarAz576Egf1oqfD8OEK7G/HEbwNuQnGVi/6cBmg6W2ZcW//6OZR1DRcmGVtC
9+abepQk5INODuNuYqgANW3LJuQA2uDvMuKKOJrGCWyhuz9q3BpKtrD2A2xF+qizY6NUkgsfbAIl
1rcM5wU6PFi97Mlskthbm9NCn4lGZN773MmPedVyVM3CGm5dfMlsdAHWyGzTWOvNIU5DtWT9ZiHe
jLr/a3eT4mdow8M4ezOS4oWNx3eLUiSpBEqZ7yvxHtTCJgl9CA7OWu03xzLRsRJkOybGs4dKW9ZU
nsUH0eSg3FetBPP6AyHN9BlJjzQCxjOkz+p3W6nsCMisBqaDO5sd5/+bENqET3J43Ax12VYp3Sy1
fYNIAMQFf4bEwRq/3iLqhi73K15mAkTCxlx8CqGoxpmTveghEx4txZI3lE0nHE0Komy2eLb2VLme
ELaVy5s8uGJLIjnvIyPnaha5Z5HP0EBRjCvXIApLlBkRGBBo4LPZyzAWCbz6qhIDoUmkXX0s8Zlq
+oPCMNdHkJ4A3qWMWuOgYXXKgbbl/vqc1bZg6woYWtPUA37cQo14D4jf8vnwhb1GXiSei8mLVh6x
fpK4wuRWefq/HUKcom7YxqfYIS9oTHHoDGtCmPrzQVUCGK7LT5JqiEx5qyEGt01m0QXnZyprrhds
v1fQK/5zemFu4PEk3Ym94ENq0Jvmq4tigDJmuhEYdRaCFrNNUY6B3g8+Ps2GtiQTVrQFF6ef77gr
NFkmT05CZbcf1h01Pz4J0XLYBrhKwMFpcov69PVWhao6dfgpil4QsYjVkx5aGqrPmwFcULdze0kS
IQquLSeANE/kqKaU3z8JV2XoerkU6sJ6GYsSHQnPNq3WSVR5NA3z6Fvo7HvXxSFVInPnYoRGmUP3
0TdyOcgvjHKv7Ivad8CiP5Xk+h22MP2oRdO/NBU2r62PGsu1RhFQ/u5ru5tLeehSwxNecdsRE34U
6wIZDsUJ0+a1BVqZExR5tRP8+6mZlDcubEORHz1DE/ru6VkRAe2iSxbsheRMdbGKezQpdagf/JBJ
93n2L6DbMjiKFExzs0Iy60heU5J+eOK30tsim9u3brNOSA9mKOMMQCDd6fc6i7AOMDO8dYrriK+I
gTPYYvumipz8fMuJ2Z12FLWE+fL2dXbVp/2uhkLOewBAIPngSAieGudVyZFiSyOtyxpi73CupAty
OeB8TGCGbbg2FUbZiCVMckdTlxtij6GNO1sLL9+xiYacZBtYXlzFN1c2DFswQWwwVrLL1tHaZcvP
61TCGh7Dm42/+g3PRqQFJQv37mpcpflvULrmS9o7R8QHsEBq2aOSxIKeRTPU8sOSHSZpraV1gM0O
OvJ1bh7V3aGrbh3JGcgWtlZcNVoCNvAGNOKPBUBtN4Askroyl0CiPU+hNwMj/Fkywr0n5pRDch2w
JHXkgFdBX8GHOfVbbU/yYIu8hQVhg3iiIWSrHAv43r+fEM3x+n4iIhDKt5G3GZvxRhRZQa7qfiyv
F8QngaMHYaZpIP0gEFpmINDio+dlLmDEwtO1o7NRNvmeJZQDJrKD1mKyn7YLOU7LWCFBQQ6+Sxhy
Q+IMHmjTREfj0niclHJfzLDvrZTMtZbdl/7GuTImsaHKrqHLTN8DyohJiIRnyA532jzP03484qhs
edWBj0Bwe04XNQZQN9laAyFE1zziMtx28WFbjsXsl0ScdpuQyN2n+ZX4/V0KoSbnYoT4ENbemuf/
I+LktHa+g+IB+MPsUttUPT5qSl5+P8+S5cBgfG0wcTPYSZ3nzA9Hse7+DjVkusXZZpzXQKFgLLdb
HaaKy93wBJuTdOpGud2Oxg+3y/Vo7xzlEPqoROKAfiGVyNtoeQ5+cBPhcnqW7iZS2uxUYUKx6Gyr
DsU6kqdIJJ4CqV39gV8fEvrpFYyUfOiU66rWkL8NVjUTeJU/RXtfRCQnHzbvs0sW8IwvoHqszqty
1XFny0hdwNSgeUC2NhWc2hqEilGu1583PFQDG/W6napn+DxHH0GKMEhCQAt9SXvlLvxayZskCbl5
ebxkjOz1CGKaECX5LgJq/vrafoMQOxqeSWZ492zWZh5HUp2+Ojl7CQNWuIfewTMfLQx1eC/zbip9
pvZs3J/HniSpjbwcueCpmRDiQBt4uEWexhnJnjHvpubMvNwRgffS48anOiV6TuuiCtZW6MKbfszA
rk0375b9SHEHiXGMyiiZe4URL8xDWjageWLTjcF4PjgCJaXEDh2XDT5CwU41+Icn+gY9lm1jNpHk
7vvAXVqC5FHxosD4Y5+XtpGS4TyJZaaIj+Jb79nA7AzwAbfE0DjSCtZ8sO34kySzVAE8lPSMmsp4
7uscf+dFRzFDFNahj6n6w+6fwpDgBA7EwVcfOC0QfsRPd7klXGG0gGwRrFmIW0mMve/FSR3MDqJ5
DWwNZ+DMHvVhUoM9F3gY59xkJUxZ7xZVZPHHTspaIe+ygf2Un0wRCY21NCgHJECcSLjojLb0P7k8
27BP3O0fJ2fYdsDXjtwg4RDJxUOLocwbCuHT53I5l6Hzv3K+mNdCzxSfSPZvfApNRZ52zfIVZgLW
XPWNbEhtCdagJX4KskaIOAWmg+PFk1l5uWzL+M5lavPfaIyd0IGGUgQrhstY98qqZEaRhSIG0+5z
ZH8bVE3lFXQAwjNbRl7Xz/dRB6hn/u+qtB07pt3AhWH7IPtCsKIE3FVY/ej5M/XFp0wFDfbyjdxn
Y894rhubrpJ4dWnt9kJ297wpL3+lFmEPA57nxVfl6hAk91z4hGTyG3fgkOGeuUwdElwrLP7DKxZp
bX0LiB4SKBSp8XtGm+w8woJpPQv6BbBEf7c5+I3AX1u27Zd7CQ8ywrHegr5pLOssefUz49aV5SJs
ozioD1l/3+6qoyNkZWdVR+QkKSZWF8fazsSUlocbsfMiCbkbUctjm0DgkQc4PjSISEyvmntsnJK7
TaVPiySiMNTJUfPuNMe3t1F5fhzSbwW4rlmjqcHVv6ANbiyqCZ0ZmOVDjQTJlhRitRKA/9iZNDWS
Ssh4i/cTUwUJzoFMXXm4O1uFZRxxoON9x2xe7Sj5K2sN/4N44T9jgvD0DmV0uRwGYexT4p5hxF2K
ZmK9XxJ/ooiMvlyX4wyKauKsDz0kipbPkiuiLV4xkRgNW3pG9C9+UH/c2wjMo2zFuZ1JM7eXOAKd
eIuT+JVl1VshkzuvJIWE25rZHAWSrS6ElzckhPbJYU7VFuBdGYxZrF1Pw4OqQdYnB7CZ2o53k6oL
VJKTJJrosGmGMLzpocuWICcmfAJn27KQQXVnx09Bwhegb96ZRgidJhmu40+RX8m1UpCLmJtMPCXW
BNoeoKalykxVeiIdKxRYK1h6uIUsY2y8v3hLZwzfXCPENCHKMu8QcmBQxRvLc/lEmZUqtY7N+Yl0
fOjH5dnQiZP/bmYAQfyWabAkGo9JyzfEuHfChota+3pFRDkAbC0rvHKMx4QMqGKSC1ifF6GjnYlf
SmrOTIyLvI0jiQqy6i5Pyk2zxHSTUBea32nc5GJ6voEB01hHBhSEMqRqvWsGlV5ctThRY8TI3b6L
JCXuOl12VZp2tLmA7zjFjz9OkA4NSPBkP8kVjs48lYic75Zz2GG0QtGELrca81YK4YBArwOigjz1
iW0KzzWFHDa2flFk0UIVcJPqQaYVFlnDQpNAqxYy+EPXi+UZdJnluwrmN/1x8YOwL4ZYLe63J5Md
/dSPwOVjwoInuXVCwGrbXI0lJdwViQwkDYTHwv2zTy3tHw6oOG+yooyOrCNqEeK6UMa8SwzDdHKv
yhfYpClDjvXhAE7jMHd0rE9fyAd9yJnJyhu5QBtEbqmOWv2A9WtxNeqlWKs0qNQl1s6qG+dhLckB
RuBhMIxZfp2nQ4TgZR93+erJJpD6MtN1ZQ4v1MK4JOQUWrpZWaVV0ShhRU+1uaaWTZpBpFYpKfM1
yVy92Iqjd0w4UNyi+rwHuJ1V+iiN01VcT/0LmaO/oK/dpQwJZ3Y8H0suvAJX/W2izS8xm7TkidZN
19WvaUQUs8WTsMoB2ASi1INqvb8UaLLY6hHkTIQFdmfdYyN++BLsqpjYcpOnn7YYsEjn4ItcFYNR
ki/xecmhg8bVsZMwjQN+fQzCG5mxSqwBW6qpFIGP2bCf0Hr6mJoOEwxT1gh0Kdb6E6Y2z8W0Yxlo
R2shvHEFGJ/PyNeJ7JmNdzxZ87IV78cPJNAtzMiwc0X9BckouI+pgCwY0JL+95GSL8Oqk1zjv1+C
7Drk7E+oErTZ8fSZuB4TdUWvQWLoJbno7lZwASe/EXlfQex4tSu0TtmJhBknfW4AzRGvQ+zY6laj
5H0gtefcfRtBVT9DA4M1kZiJyoPi2oIJBjeLP4c92pz262/9ddzNTgiy5LJYGaFhsE2+MkgBiJGt
OYyfZ+fciGB3+x1dUhJXCG8OckbaqCOV5D2gklyX3m/DQOGZNC6+DzcJVnWylwBryKszPVAbmpoj
ISJAklOVOJ0YoX7IhMg9XsXGvWADSl1q/o9cvAxhiWuROU6GYL8DfHy/f7uywFc6OxfxmRHzflZ/
pBXbaou/wGSUJHDUHHlaM34DqVB9CxzdZSEl/M+6j6/B7Lnh4JCNEWHOBXQHhgF25rSodh6U31pm
uwNESUDTwlVY2WhQ8fvdXJ8Kkpjr+XUcKjFs8DQGET5oqCY/aiXY+oFOhQbhd0AhGECw1GkG9HJc
8y0iJmseYvxtxlR3e656+rqy0DPx375pDc/+BQhAf6B+o0FJsr47hNLbl3nJc9edOTx8ZWSWMMeC
MH+p6Yg5bjKgkjOU+/m8+5cbZ8vYYDB8vw4vSRxecWNlQ9W792UHnUl9zVMhtST+FeJdjzDbf85q
4RwdRr6IrImjDkNJYYRwIZwKYNqqKntEK8YIOA3fvh56O2gqEDOOlTNYp54amFa7Y8M+u+qJ6/Ax
C0P4D3KAKUf2tA0b/FZFKiT347ThvaCBA+FEGKPHVJ/EaxPqRKXqKQu7rJPBZh1P6mPvKzQ69S+M
ryoP9diVczysJeCUM+Tz5l90qL3Kxirdo911DJFG0ndR+Y38+PnNA/BfCm6nthbE+DFuMD2pTGuc
o0EPG6fYZdGS9HHZi475EbPu9jcuj8etxIp5HINpqJI3SoVdPikf3Ux52pakiW1jZWgF3Y0nA4BC
+cI9q3YQjdeGEHf5aNfFL4Tko6aWRNciW+Mv8skvEZE5zQoayJiCV9nSy2mQs04YA64x2qOu7vZd
IeHcAR3QMdgU8wCqJ3CJwAqe6fBUJJFglmX+TEtDrI6TJnKgviq7O0tJkEv2DpACBWndAq1eFdDN
Mv1AXhgTM3n+j5dFCYf3P/WWcYRhwo/bJUIdGtbT1Rd+cb8DUdQupNYujXQTfcLucSrljMJj6lvp
1rq5+6o08fqrJ5scgAi4/+zZFAgjeosQibY/3QliVSVFCN28KOS16x3qz10wkag//iU98WJtjBtE
/N/7xSt53fmvDo4z0qKo05kUIr2w2aojlSGMTjnakgAO4nziQ5U+kVy48REL+hhZAHCB7zl+bdy1
cc4r8r8JyDXwgDVgwrw7eKdOFYtsiB4YBffxx8l9lsF5U7ZZYvSuNWB/jHD8LaroZMOrmFZDqcEB
Q31cBf84Tmd/mgQTxGzM4+qVxvqEjepVHnFiSEEebErE3qLhN5BS7qWfI3vYIxT1PbdtOfbaM9IP
Dkxu/t3+QCdyCczJ0u9gHHhpF2ZztNwcpsWM+gu9ml3VrnRBS9qbAs/fMendsilZGC/baZEog4SI
RqYS6lsYFmB6O74eD9JvIz93onVE1UOpmmizX//e46DJEftGhJWjeyriXeR99zlp4MbGRWqjcQsp
0YmLA8+kHCq/RarXo22a8ct2Zz8cXJwKxl/bxj6Z1uXJ8Gci6lcjvFEWVbppU0DrhXwaFjUv2iu7
6Z0702vBjyX7LTWVPsiygoFXUXxr6TBSmm40Gg8+5T2vyemN3Dfppd7d3ncGJv9UcS04oS4Yfcsv
DqifSyDCU7TfLjhf0IL6U6IMXvl2pcMAAXk+ory37+yBs7wxn7FLnEOyHWjAMsxL05XzSyLxII7e
y8/y+tKZjNkWUdK+YEHXhbIumfda/XqdZca38qBQpBTMe/gZR1enmIybVaSE55VgIQ6n8aVUXjAl
S4W8HBHBI72+t07lKaojpRgvcRf7RQhs4yLSDF3S+7R5tvxnfotxymbmjybUnpyQCU/Q+8Tg5Uu0
O7xzJPdHLfaQjhNdVzgTnSfCwfWCMSd12nvQag51fv4th5d5ZILOdvljhbOUMz1eS3PhusfwsQ4N
wXhTKgmzgo84ov3oiz5k8PavM2weuWFV/LQaqsVIrZP5Ls8DLfE+sSa83ketlgVU0CNExA/uuhuv
DN9a6htyi4Po3GGxzrQ4HL4XYI+9I+pNxVxbfi73aZk6zjFCk/o2icx2tBspmz0XnbHjrnvrH5sA
iY+98AVSSjTGcN1phXgUQq48AfWOTelMVb730ejtu9+EKMCNBr4rXv6yuqgC4mqWBKw2F55FvsXj
ho9mp2X6/MrnXavPjf/Ro75C9LeAXaHOweCPDdRfCpadk01Wh38QNTUhmBQd198bRPE3tzBJ5+Cu
lkWwB5dPMZuYdPj7VJ8pDyNqXpqYuQbED1e6m5dlelWLNzX8XvwOLr9EusCk8UTO2YIZ4uNceXYd
EPWDAWLEerdElA6LpT/Bv9ZoZGfe7nM4AdQc/y53sz2i38ohkqNd3rSgsLOYyAu6iXoazLoWUMw5
tG+0oJfLW9B44R82P2efOF4t47YoDAFjTudOz7IT4WHDHzJzCaDFQXEv3Z6qNfMfq5zEfUs6ghcm
TGXbt0kaeqbs1s4bDrFGN61GyN39/tpeQF7AL5aKolMSNo0Jq063jBLWVfazaFKNBSFthm5wLOsy
l0dU9JZjMvYSm1GNY4vvyUu5AX/k74az4c2k3T0YooIuR69WNEDsSm558JJu8GOS7dGUqmGqoBUf
fbfs1ro7f5VRcfgtilXzfZ1KiEVe/oe7crhyUVtOjk5UIMvgEfuMpritQwIWt3lo8FQlz2wUJrau
u4ogoUhzx1ll/WB/XI4FTDQYTRUmIQOHaM4DKWJSg1HHewjBhk1Lnzpd4EiofZ6VS9DDGrZhOJuK
K7Je4haWE/L6J5cJaNpihPd4XShP+FiVkTxoBwr+BxCT48KukNaNOo9rjgA3Krxmj0fsJUjRpXCO
/CUPHdLlEWHxJB9tuioEzZ2aWjg1USCKcyot1grYfSTmshm8qkFup0Hl9pseOdW9ztKNvzttZubd
oPEYVUOEr/TS4bIC6l+f5LFdquhjWo2P6iyeh955v9n6ptn0IjyAA+5Cd/JGErRIVTHgYgRNzpE5
rPu5OMkt1DTr84liaVKDPtThCBmkPZPQOxhNCbVITskBKtXlSZJs2aFnzcIANngW1GmaeNBu8Y3M
+j/omHRwAdFBO4Tdl/UcJJjbGXSJ0mWNPowRM3lF5T3I2aCPV9jn/WXv5VochBlOAmBEIG9wtoy0
wh82v8Qr8dvmmJ3iGDa3OUFZ7l+eeUu3MErWGR9EaJodX6Re4h80QVWJuAyBN36XkwJGwKoxeg7B
ZvbXr/kWUemL5Mc2qXess+fyjbWbHggb4ns1QdiwowY5tU/7Yxi2/nq4coTwh2VPXqFAltzr4EJT
mT06kHYwfdvkK/6m8E2siwH6aPkgR7e3+EQpzmT1SVgEybX+aThEGy+l+kGjch/OVzQy/OzgMRZn
VXZr0KiY0EtOS0jCaVVY8Bzdg5eI0h28QpiTxioOcFBaaNYiRTh5KC51fb0KcoMbP9wVIjBhkeEW
EgoCXC1V+zOUZKkBgwTHCpnW07cdY3FLGHq0BcYMcGWTkzOT1fDlLto0354G15V/86P4zEqL4yiZ
nKj7QedzIKxgknjU9iexzmvvX9iuMfIeqHkxACo3iupMZjLZgnr6CDni7e9iPZEOPA10zxX3vUgx
pqTwqNfj1EGL1QBElMs7oTmwpcJIoK6rXmNLqMXA10HVemY03RyZuU4Sf3w/EmTPkhV+ANGJ8+qb
ApmTP47VZ45/feFzLT6xnOEi/dfxHeeS5cu8MBfKV8qpCMuQkH+9JKQ9U70ctDz94j20Bp4VYzrT
23CUc6awYagYOnL12NNvF6AGLsHNqwTBYBIsiTdcHYqyssFCjC/jt1FmUAHZMbniRjF3v+uf9vK7
tgQBHhQHdT92w3JB57sq0pO+bcUhokHCgqsBVlVjLRv7RYMks4zYGEM1I6rBEykREUCMGcKw7Qyk
mi0aTxYPg8P7kw9LIjS9sObvMQ8WTOaqoWL0lJs0LpOZSZZprP/T/5M5AKFrua1lhi+elolj+m9K
qIO+nuH7lXd6GEK9ufkCGTqFtXsX7JtKBgKpBoCHdi4zYDyR1z5tJMapxIwDGnCzZVpIgRL3tCbh
NkGEXUof229PJN02vNyQglGK789s+kzMgO8OOCjiY1U1s34PSw5z+WnnF4HkJ2FPAfWhRZq/o2O4
8wmrxV13Kavyn9M5Bw1Ha3FXXExLT7TxVOznf7UGbKg8RGfkqYg0GqMql0dlEtmmAQazB4PLWAA5
PRf5U1BZnASb44XG7aSdSik0Od1CEjHaQrUDFwllgTqwe0o0+m02T78JfsU7hdvY3Hb0o4Gk/X3z
nJDLqgrwskuv3dYDkRj+v4obzGX+mYevwbSt4mH4ib1jowCuYac+0/ffs59p5qrP9udG+Ic6jyAU
aiYAwdvZc0eVExk5DC5ocvpW4eghSJQY7TBZ8QVL+7Iy7v4wI6NEarFuagfHkmxIrC9FbO29F0Ns
eRF3LjoHHeezrdZLSEX/oOoirn7AuljA+ymYkBWb7sRgVGDx+zTSRWL6EFrpDuLSwQ3T9UA5Lyrz
y7D72kiVdRw6aYmp7kxwr8RrqL9K0PSlVGFWUqFP26l+SiZeSday9UK71nWhngIQh5mlZfP66uN7
vRDZyDOPQKZvPNXdyXckMMP6+xvqtW6dKVMwzpnBJ+Umo+ozZe7xWYu1f4SIQajAr1yu9hz6LtfM
GhieDZawYoj7HBqDLGfnkgFEeiwnsOTdZgXI8KFzq3lW4nj1nUEfyGTO0sujGjG9c+3jHFON6ya5
a9ujJ71fAdscIRhGBeolVHUWAQWBD+pRbkTSSzBUqRyOzSI5VU0OCz+odS0zPqE6Gc4cOGfTFzmw
aWX1NftpCe9IWcatGPDSoEQx/wsLgYj7PVHfs8y5WZfK9VmwK4dEX1ZVqKxN6u3tBuHmxG0mB2lO
Ma+VfG5WArgGSvgEvW/96AjOiMlBtpnRRBnETnxMCFN0/mE235r4IkKO4UErbMVxKa0HuhPC5w/I
bCuy8ErA4xh8Hfy9Y3JKEGDccrOD7KLYvysROVqksRpYq5kduv0QOXX44zZCZ2Ok33Wpab7gX/MF
I3mTCnIxXPp15Kh7OJxJmKIqxMdlHpJR0c9cXN3HZWMlm1VFq60xpEgfojSLfM4FpDC8s+/9W1fJ
gdAg16FrIC80HHW4o/4pTnjz2kZvUf5dLLGFS920bU0gBJhqO+MqNT28fQe7nUgYMrlqjeAn9c+T
X7NtWGQ6MAvlbseec05KW8ekYyB8RTq3VnmPShkj12RC3ppXev/xhOxo/iqPAh2EqfqU8KRRLYdo
avviboRtew3AhgevQ4ab6bQkdM0RtwX/diGGx2a1lEj0+DZp0vCi2zzVuRzfAiroXfg4HEg9hz50
CclTBc5dMIzQ2WLONPe1sVf/VBxFN63HP6xhuvvNS3A6uCEYGRxOMlRbWcJjTl3FSIB7GgZq8ZEe
gxICCBw05BI8USaB1wZvIh8bSlhUR2SwWi2ykyWuxTv+RA+Q1uz+AVdnQTiuFoxcQMGeIyQxMFaP
z0PWmmqZmRAzRNrrPMwHTuxjcVXlDnfYPgvfYmwXRh8iMIBaDL34FJLCzf0yvAacxoSADu79O3IV
GOf1tQO16QOLUYeMIDy97LHC346KyxMMYr5L5lnEvAWvkCTC/wYu019fnr7g8mCKmnqNm7eHpczc
S96PJmZk0lrAnWr3t6QUZJFTYORMc+rip9y9e/NWBA22jskB9oLh+0UxjhEXtHVIUIMygu7dNcd5
8DBb7PNBFpD8FcRi3uU3C7Gmh11hm3gBfpprgoeOTO5VkaGegaT/DylU1/fdTp1quhM6ow4zgvvw
zuVF6tYkWzyUWT2zyBjAoPq2QJuvDWtNOS8B20daR1Md02Iv6Xa2qnuQJSqkrXr04ium72r3Bqiy
1QA81apgKZnpPC2haIO5UO2WaT135wo1OSsSb5wJozgJVD812+Pe0gRrGIfijqahuoq+ewBSuWH/
CFCYB5IUEZtBl4L2nZxiKU/2IZ1sF7kMJx+8Tlb0uUq58CzjRaMii53O0qL5q2kAXY3CJ21kTojh
Nl1871vrkVQ8m9I7TMaUCsJXx6xenGZ+oXB1evU6oF3d+uVCs0Yx+irU9tYVBhwiV+4SaOkESJD2
golrXgNPoYmCWKNSZjSJCTZLqNUrAEcpCxyqoWEddAp9QUYENv1NOUVrh/AyN2XklBYuIEzAuncl
Zg8/vo4pOhStG1cMZEfqdblhV2idCkvONYMV2j/mlXyDbytviPASLf6GHmiuHOrbftDCk4ZOSm3a
yI8mAGozVV0AoSQCqtOmc9DDzLcIVKLX2phD7bC3BUlC15sgiQ+HIjX1RcsOQnok6tpx/jXR68lu
rrSh15Ovhz0rAqZFPfnyY1ZTDFYFRH0ZIYAOg4SN+6rb/KMnzz5bJuN/lCGJeYUBzW44FpgWgTsz
JeHdATMAt5QfNePlEOhP8ORuFIyc7SxrPluNKui43cG64wBiJurHS9SAXVgLCJRgbguOPiY/aIrb
GFwoL6CwQixw1N2jPGpRT8RMUKGz7TJ0w3hElzjmocrj0hZCoCVcc0Ig6iPouHBBeWlPnU48z0Vl
7pqZMOioNp2X7aHgDT4AaTcUL7rvnok4v0nkyVEFJzbkNNU6SNPNqoEoShiuWr8l8jDukyA1RF7l
ARfAp9TZg1MNignISVwbjVV4pLJgNArHgJOCD8u5SB9ce9690o27j7jCCZQM5fwyo/+Zf0A2+PSH
NVpyKQAfI7mn8OO2P0obKWchSkEhCzjE+9LJSbyb0RB+dEUkP5Ld1iaTP+ArJsGp/6DiHImjrZDK
ay8OEbNl9Ix00dbEryaPWHgEwd/majlc+Dch4sbWfR9lMtsCdI0/pGjxq2Z9ua5lr64Lj9yFkT62
JFO3v0bBGSvjUa308JiwIQklq/0aSekFolGv5ekF7BnpDXNM9t2gngsyHFo1supqf1WxQH5yONBK
xkDApqNTGt8mju2F1vdgsxH8tjAWc+tzhR9JCg8/CzOeY4FY6LGnzUT30Oho1+dLejUbmVAgvVD8
W7mA+jVDqpzw0mHVDyR06+A/iKW0jeJtxLjZh2GACOCoWi4oXHlyZQX9QzW/jEwCMChIRBqwaWsa
LN6pCRIvnOHXa3FH93zcI6DBY/h1xUb0/EcCR6kWAWHwPTEbfPeBAEu5Gkcj27NwAaC87otxHie5
lHn725TsrRJDbSNBMxFautkJNoxCOcyw7VIeWGoUJGkiR4itLasWj0ctFcW7MIuCw0suQdOeCrB/
cxDnyp71XrUbR7M14uJfzui13RksSuffzIgIhtJnQVK5TU4fv+eaFrxzxeM4HHeboFUzfjvCzelh
3I0gtB9ZK8RqGsYSTGCLEPAZAdunpg45SpbeSCce23/p1YcAoSWlS80i0rgyP468RtGtR6KJFK24
QnDppGps094wAAJALOfkVqUp0oabF2TFK5JOnc0cr+xyCeLIYv/WYCpvy7Rv5kGJ1OM1K6qzuvfE
SXdOJZ5s0JTgabRlAdJFsSuXj8ewT40Yapicb8gm1qW+e5NTBjGOdQMxOIFpSROejlJJ4PfW40Pf
9sDeVfTLX+Ny4N4tQcGZS6rQBHLhM+kXi8bH3t+xyzoFeb2eT3JHaMgkS65OKgBAJFyu/maM78oJ
b+tyqmmqIuh4VQ8QTuGCfjJGG0fEWgZ2BiSrIk53L0PUeFNAu9Hp1FPJQ42eBU0LHPIs6zJoGIaY
Yam4xpdaLH1iDfouKT403tThhfRr4bdtyOHDqnb0FJlaRlFxkvifLObOt1tH5F/c3Dw+steu6NXr
4Q8U/dNWenoyfeBeWhiI+QSt8fVe++SvHTP313zXI3bMc6+TP24+7SRkpFZi+XKXtqaOScFTdaNQ
mGG6NbIkw3E/3IKrvIEDoxa5f+9Y1vummUmyDMmh09Bq49IjsI/bUUt9S6oPJCkqrnuxNbpjxcX1
92toh3pC0PXahf59U5AI2EzAw1lgurcNXlYc3fd0+D8T3cJSrdSEFwEzavXh3XXEfQBi7IVTMZTk
sJaH3AGHFTkJhJMTtmkjn5Zy/KHI0FxrJYODf0g3gIHtqDohCgCxX3/YnTcmr0RbYTKPhalOKBjY
gemDfSxEF+RF5RgIwDkMfg0Ld7xPEeZxfKygjRQzafpMqSK0orZdsHAXM3tTVjcramIN3rfqLg5i
Wvhm4L/QBf6wbfRR4Lh1zNKR9m0/bYOpw75C7Dgf+ej+ujUkWh4L/jaMhRHy3zwdGBBNIZp6QcVb
L4PVCwdn1anDlr17+ge9QWiNJ4irlT21EAIMxAmjAiRd8xr+NtAw7Qtu6CdaYfBflkakXXCbGfWq
nkrOTExSVajLAF4pc0aiYA8giLW6/3mnN1nDlMyJV1Vj/hhroAt8ncNgKNuLym5L8ejmfU0O9TJg
LxoN6yR74RCRQC82u2S5NslxaurbO0fDVOh/csnbyoQF8YDBafT3x2phhVAZwg3ZLlpyDc1xlkOy
RuE2g9KCNi6vYNoOvQ84evmt305FUsDdZP/nslfNRd+esXKBbOdKDtpPJF64WzHo7ndUcM/rpwG1
zCl88Cv1AbJBQAnJuet5/S8SqEL7V1iWguMz49HBNaZhFwG2ImHHjC4F0Lg6uJgoMjt+e8Qp+KRG
qMVYjcy9x+/org/YG2dTxHm+00p5VNZEDfz35Erja05yrQeAb5XxNyG1dCrDa0etVxuEIdQ3nkKg
DptU9vpkN0UD7dM39JdsYSK2KR0pBNzwGdfzWD/ygGBQEoF50yE4AiLhIp5jWn8yVCDhdebJiiWk
SXEAEilIFP19sSp4VRRWeWc1YhxvCnfyqcnkNZMVHG7KpkxO7A9dEmAtSedKGXhcDtGKOxjEzPp5
YofFS0iCEc4qpsettE9gJvUr/wY0LaWEH6eF2caE1lDDvDX56gjRvyMrPQz4whnBCFMOGXC2X24Z
2s+5P4xB7QZEg+B+yqZx94jFKhQ9QbbB0KMmJe/EjWjPiKQODYhMIGkz0vKp1w1INLyRnHqRKsmB
ek9mvp++kReu/TdP6c99PYG9fztZ/s+vtSIb8Z1jFJMINTiXyTIxK0gTcoLTm+C2ruGUujGYyeZM
ORtr10d09qEZAwNagxkYOSUO6t9jiQ6lrdPmuNvroO9FHzyxRy5CGO5R0/em9fPza6aFPaV4/Wdu
J/OMgemTg8bOB7AaUTIQgcTONgb1iBqBrg44qBbon5eCKjo6IrpNpFR+diuI6vUx8IM51UkE/v7Q
O0hJfhhLwzyqA9Iysl1yrnY7gZ8tk+VJnJGSBnUb40cxCWfSiGinY3hvzpLanMn5WmNkxcsZ7wGE
QfzLikhk7DcpMOC7lEsenkk+oHk4IariXezaiNoCc8Lf1wqNZaIx07XNxGSULY61/zAXbrjsEw6P
YPyQbywHTZeW2x385w6y/imE4/WWayhzvS5vBCcC7iYuzpYMAvF/5jf0/kievVi82J/pO1rW8XYw
0nshzaqUf7Wa0dLjNWomF4UcA+/ygghtK5w8eSQskE5mowP+DUk9NJ8P5Zt3Que8pmweoyU4Vo0H
V0Y2a9+fSmiPcExzAsJJZuVrlYRH3y/4Oi58Vwn9zHSnTryKknYquF2qwGP9jiCYrEXnaOvA7B0p
dID5/nAPO5v+yywTfEQthUdjf76HahQFRfM9lqTuDcCDuxnJX6jnc8LXte7V4aZ13SZ7KTP4Smhp
4VDroTnb5z69KHltL44mRhvQcEK8BBlvZrcHW+aBYUtCwptY+0Zffu+q5lIc2ZW6VxcIeFuMcXDp
s2ec/QF7Jk9+NyaBIl9soODtN0js5y69uFq+Umvexl0QSxQmNBaO21CqenHJ5JmbDqGSze/7KdrH
4wA+devK0PWKLqfz66g87Ok0gdUjvzhmMM5wdkYfK8LbeZym+PuODbjJ/EsUcBH9SO9YX7S0pV0b
5EDSK41N8PWUqEznz4VvZk7Rsl/haGlfWnodCVSCLNs2nh4IU3TUKBgyx3HEp+rFZnUSVlCDDa32
yqNVy7l77cOBqHX78zWBk3vo+3WvE3id6C5Hj7LAMGFPry+UN3SdoBBIY78C2p+7wT2TiKml2/yu
3QWB/w+AY82dy8Utk+Xzu4qBshLAsYZEpfzMrTXP+6izI8c6q7LtlAEnGsV5jCO90sZrwwJRkei7
H70Rt83RPq6jWYiNg30klORN/VZCn4fY9uQjQlG9oYW17y5RWcuii0eq2oOOffo2Dr0sVYWtqMEW
ZbOEkg0qsS5RKKPVbwIXNI8lIoyX/lVyYx+QtpA0hr/RJHxpmWB/GPm2FgbAkbwUEbdW+AzK5DPh
yioo4f73I3QUu53be55UfgPeQJ6R3yrLzQ9o4x1mGdukfDkMIfVh/EA9Y8aBRSnAj0WszyiK8ID/
v5mVao74iqr7/hCgEkwAP51ACWGIc5kxVBDag+3XK3NmadBEnfO63KgUEC2CL0U0+weLh5X4hDpO
1/YoEhGrjkwVkRKjVVdE+Sle2juNenqYyYjJtJUgvyDjxILfx2cgrjJ59C6w6rJzmTvqifFKvqlZ
moYYdNLle5Qf2IvL4tW0QFZq503uog0J+R+2WV3TFfbQb9bpiF7FGl7WFahZsTYCgNp1J8MhHCVV
kZ/u4j/Um3+2BTFrkhRhjj6O2MxDpdINn1qk3mnaM9pk/WEdwxmF7Ftr514hYISstBZYI1lzh6HA
BJtfb4LBoLdUxrJxpttBjzG7/F/h7d2vN58VdE9+CZisORoYTZ4r62aiSGcPDdfeNkc56p7d0Bsd
C2vmOyULSVacQu6G5PEfjh2vzXtwhyKRIXiPHtpmpuo/qhS5s5mxaknWvaAUeUXgqr0pK/1vK7NA
4cw8c6NC2VssLaMzo32DYDjbg6CzViZmSDaFMSLHoS18at05PgKnBaZIqa/mJIaD31sTf2kpryp9
Wc7IvhLivSlVwqYtdkefkd7Zu7xfy7uNGoDwJvDD/pNB8TsKETEZOtfM7ZQE6a3ebgdIMK6gwmQS
G53D670qTg2r/jrCx4MyHznaaWfIiyn27GOh304VLv64pyVLCytfkz9JPHjyiBKGXBAG0qAf8JVH
iBInkSDprFCOkIxoCVxTuc4pwOWxw7XDG+awYKrglmy6qKa/bSMHsOc5NYhWVbj9NCzxqmOFF61Y
DUpiuita2Ok8Yg+z9GO/XuWn41rdyM9zEFgG4D9B6vnXVX6C/mU8g3dhHOCraS2BFN6Hpt7IvQ/7
ZfAWhbUYfeyQR+BPtRlLVZxyPffeyMQG2gsrcdzTsfesO6SbKaT+WhC8rRcXIw8CJabyKZIv0Hnh
M6Hq9GQO83ApCbIJVTPfRJhZ2YI4n+nZcGOl1QWsWeS+vlcs7CvVQzCKUKM9Hpvoj/UBuMSZbOzA
uBRzeRQTdmXq+aqNdeMwzLr5hvkVLRF1zCdTA24Oln2tMUJk8YPAFZTTk9qGxpmy2ambjYUGcjrg
VlWeHUwgOmxF56xjc5EF34X/Fid9AMD8YQjxkF2kamluBLpmftPRUb49ZyZbzZjpsn4IANgvJBIC
sI6etxd4Bq7ormthMLpRB4XGimS3M0OBJ+H87daiF5MJEqIe6HqrdEeILqjm115Efsd+HorOLezS
pDCMMFlFhnD9ZVL8QRjnVj+iutJSQgHEbmeW8yAwqNwegNMwyJhe2maV8QhfXU5JBFXVJawRKrWR
4hblQfKYaagey4YUS7FoFfwDPjOAyZ2gUBUvR2qR+IY4p3T124aK0ynO8Gf8Z5/G6V30pU2wn13b
Xn2lSi7PJ8oLiPkaah/ny/DbhzU9zJRGZlZLTJKxwiDL3l+lpwG/Pca044YZS+dA3E7pX9Qyk3/l
JC2CTd1xMZbxTGnWKul78iM/pVlqLguT/iwC53Df2Jq1617IEpJ9QuS7uWhbgSSMEDK4PiJbIIDO
+SIzRibyEGdK85FuRkBNWPrPlP5po0tZOGYAYjKK/cXVJmRgAtZMctJH+eWob4kCgyar8QYErK+N
xa0vmFcl5WQoBSvwUO0FMNZO0olPQbpB21haF3jWQHsaE1/I/9Zza66jawUxPVz/XApYDoKCYXJK
4OFx+kV7OqZskoi7Lj2JLMpAjFzSXL2I7Y+Dqd5skp8WzWj51oiDb3Ctu9+apZgDxNrFJRrEf5rK
UxCngTRVQ8JryuTIqIL4ddJmlWcyBc3Uw1RNWzkTiRuljBa94hxGDV6baqYno8w/qFCu2owD4X4M
RcH3+Q5ngYCw9JKnH3ora6qHz3oU6Hyy6UYHgJ+i+0TMjTFOdEljIiOyHnAEiVSOvA+F5+OAPBlF
M/gjrWMb3KaAXkgMhZjQREaaY5EKL+8MLV8fLw6hpWNyaeHzQZm+w51QZFc3vUkk+UndkbLkIojK
0fmv7FOhE5m1/LAKnp0yAlK6s1MkQB9gp3ZdetBXbvyYvS9fl1maiZH1sbBJ+SAbGRJZZ6x0l2+L
nWMdY1NRt0JNyDGD5RgUXbIswL2ErRjksWBfOa0dnQ28URDdERC2qIhqccJ+So1nWVCDvVQXSOP+
qRBwKYchF6uFuyZKLvR9T5k9o244LEYamcbnvND3qTl3gxB8LdH0Y9DDa9/FmlL7mOXZ/B4iJjSc
V9Tp+Qjydi8H1RQIa0Rlta1Jsk1yb4HKrHIh5cC8+lSNFbU3Y0TOyKymtQNhTe1S9sQi2WrtkphR
duTsAqXrav4nZsIcetGZu4LMluDvD2zikOC1o+aWYe8oy4ybazK3p1u8h4gaaaxAaMT3Vxd6uKmt
IqXncUsld0prO2aalQ8zBB9WKrRmPKScX9liUqu0JUjzJF/KEsp2Xre4S/Jmlgf8R0wPuCe7GBHP
exns8MTsgaypKJO10+JTL03qdtovveFeXlQoc75FC2mx/aUHA4sSu8AVwDtMZBaXhAjGaPOuDVXH
qxAzbU7MfXh+U4gvY7/z8NnJNDkF20sH8CcZU3C855wdJbeHn48ZFaI/tc1w4K/HUEUSqP8jfn/S
0yZFdjak+rt4DR2JRw5QXxG/pijRvzuxaUwt9vjwGOD5N41kmQYwQ2XAhEUx7OhK7BVn9TDmolW3
ME1DzY6csMve9yiNEKx/TB7ywI+09N1rldPpJUpUeLAaTKzA/zpumzpzDNKD1rfwyOSCeus33y5Y
AiLVgtWWJSJycJ/tHvsGscYDq15NQYmlqTClh84NCe6UgeQ1GDeSL5oHTlQtURhmm7tQlx/1vb89
49JtK2vIkyB4MFLnCEMbL8HQ+W2bd2xDBHOI3qxAmA8udzT96ZJ9ezR8eBWsmNUoIRIG2RzH2vTB
Sc8QhTk5jao/SSP8z8fjQ+NEjmcHjfDPGOoeJQNqyGPkozWurSJq3vUPDsPgOR3qOI6C+ZWfkc8j
unmdKiE8Y9AGD/o6+qiS+yRZ7ieG5kpat3CTov2513QrmhXJs4QwxnnLCWt4YiGOgqlM88qLo1Fh
z/eBjVQdHFoJ0FVqzWlUbpTMi0sHD+CYZLPFz9lUeWQ+fJDikX82nz5vyeLmP4twxAv0qGXnOiYj
U3ICjkXQZJWFkSmdPRZhim/Vpobp8puLIoRKDpFq7leLZGTgNBRO/SnhQpkcn9vQODWuFXesuBc4
AqFtjEX9jCVA+zPmFYocV/Bh15ao589C13bfWCTuPaO9O3Hgj8CiGb5232GYVzOaU0xNmdsyfZ8J
jr4OF386S1vC4d6Y+xKvczxFH9Xk/JSbCeIGFubhu38WHMquzI7B7K2WAdLXXzJZjkTfTcsoTOY6
BM0uTdtvvnTh43VOodMny69fpBl3/1BrQCPoZFpVYAA9nm9lNxXhULShoW2jj+Q2XcHHjIS0HjnF
9iYRs4+bUHnTFVPyxgNRVlkqIMgLP++bctWJWzngBb05JMtQEyTlfuWL3xO2OUOBsc7DXI41l42k
sncrfw1HpwPfahRmTFGwvGGqJ8Fpn5WoRXpbys92NJEKyz3iWTZUPcMyRA/udmebNrCAifqJvptK
2Cm9YhKazLbh7cbXpaYfptHYGCa8Nxuf3dwAOWRUJAQdPgcZxJWcCAjfmKVPN6e9ZB4g8KwBYio7
1qDFacGTCyLSni8Gp1vGbi0UGicf5NHaUjmBr4kgjYmYw/Gf8UFp3758cBKWsN0s+zpFtuvcTmZu
+7RtJrfJ1W863CEExISmBxZZWxCob/OOwW2Yf+zgBdAx5+ur2xcovOyD3dn4U21K3K3xHoU02XuR
4TL/0psgTurkCMR/0Ojfg4bQ0EheR/mRMCMg9TpT1chgd4izWXCFVsoSc4J4QLJ95Ta02Z+Y6OyA
Ucq0UM5B1wB1oT5kKjpa2kqfnmKJZYeBEt6lMuT1oFX1gf0iJxEZYincktH1IiiRCZuJpnG3ycdL
vpMRojVTSxQbf+2qm/IDxbpKuv2syhlWUcpu5u+pK+MRskV4ufIdB/09N9nf82s12ATQZ52Iem4c
dyxWUDRxcQnNiSk/OUEV87DgL1Wzu9e0uU2rqLkSZlplgM2ST5BBS6NxwriJz02a2yk3WIcpPtUx
4OFxxo3Al0O4QEv+kFTKpJpIMZCbG0p4hSVyu2WyAcf4qSOxvCUKqQiWVPKhfzFtG2fr9jBP8Rwp
aKAtNSKyzGahXb9UtQAF69Sb6aGkgEoaXPKRvLSsMa2hBQscFxABM7JEziio6RfZlsnRiPmqCnY/
ZsrnCb8fpkfxBAUV4ESYNsC3RiyVmwgSmVpSjGmccBnbeuohksJHaJNrXzHQjLmxV98BWayWGr0p
N9UoKNKLhnz8GHbnvppdgXEPFHo+u7+9Ek7iEF0pQ+c2eaiBKpTEtzfzdx+b/jkQ+KtEoBXD1/Vf
LPHQVP/aSABsFm6x8/ZAzzhXQPe5CRRzrinqRoKAOWzvFYuxM52eAJmVUHgpgr61sw09rTgTUya/
LF4zPf9ZJj9/zbAfCKHV1derYA3n31NAaPb31xzHExSkEGeVhIU+bilVD4IfShnvfejRfabY2oIi
X91sTo0CSZm6rFZ54KZ+8XDxCseAg5Q5Dnj2sTFu3oV+0/3AeL52OrHc2f6plRSjBe6qzAF10N3h
B5DQc9LOR1a9Y3LBuNtuW4P6C35p19Qv83scGJ7QLgZxal32KrFKlFDcUXgylxSyvpcBL2YtDcjE
dN9ny5v0VotwwI/pCxe3ZcxRm1Egcxv3UKvIc2sMGLjNr9JDbV5mlbK6JKbYdVozFWXRotn4dPF0
ojtsQW2+jvEeg2RbrM9/ty1Qpf2XMWtvQ20osRy4aPcbb1tyM74r8yfyIfccvzV9+wSqrTw/cJrf
ootW17GsUX3M1SZTSpt1s9LErgdRFNu6kJrS/1InkMNH+m8dQ3lxP5hbAeY5JQzpSlm98FNq4Ln4
OEn9gpIeF60WQF18ZzXIMKRcTCSFWEC3N04DaYXu4mrmdwuc0J72bIWskZkSM4cR6QDUhqqyrOf9
M5FmuB3ceXtD4Ae7zy7sCm0/TR4Q78LSWPhkrXtFTQT1G0/M7ScwLaqfCb62vUrZYMqwwobSq6dG
RBhRq0babqOg7ORm8WLIPY1fvQwEjv7gwT51e9/LAvgrIR+7eocJm+mQj+cBgjdiPovuW6box+yT
6Dje+mtVhwD1zTSpFE8tkbK7gbJqFeLQ7sNRP2C2TL3xAYlnYrVdMw+Jk/bcbx7zNQ2hirPKHbNW
AtjP4cWc0I/NQBfG/vg2X9SyxqWfUmp0X43Vq42S1Ow1tKigEUAcG7d/FTF61s4FBgZ8Agzn8/Yp
LWM5wXIWv6QTvt7wC6QpvoQX1f1pkdWmG6x/uSopb++LoTWM1pkOLHfFBV9xfIC/RS4EO/1TrvxL
TAtmIvSmH29RSOQp8ZHs24tjuohrK+yIpB1lEdu0iIK1kMkvWFpXoo/nffiTdi+Jtpq4olhtgENi
OBTlE6zTB9jZcbfAWrjQ9Sc6wI4Odt7y/srwrH1LhhoH0z4cP1dtdskPgI9OrFekinDmbwglbbBw
Ls8xEYAk/2cCHZChpYqn91eJJGqcxXEcNmvDAj6Qd4BwVGEQG2c2ktKTESKQFmkkJsPNTwE5JWQx
f1bCQdxavloMnGu3/N0xAm0tFVFMaUvjOHV7AqFPTdziV8+co5hF8bTBY9HHZMQVcuUoXE/vc0wd
FdesNjr7rhxXYoQ4DfX+sgjRH/8yVeYTjvbLv81mRfcDQJWdOZ32WUHaFCBBkNRk2IgMUX1P9Wli
chBQ5FsDZPNoXmBIMyJrT9yMIrcjC/ErHsRl+skdDTsWt6SD5iyGIxc2CULQTFuj6kZKbmDqHliY
70qWkTX1skyd+/5hv5bjsjlp4G2t0rt3WJxQ89QPCG29Yr7lFbnCPa93OrzlMb49I6WlfZED0VpP
LSt0sdpyHalbXb5H5haeV7KVLtM4PSjinJF6DQighti4jfg2zVI/6jNoaVH18vx929T6wB329vr5
OsCYuVeVt+KpkJd+4xIf+B56WO/5pqgXLYtpozxaRl02/dO9Ybdpo7mYKlF3r+ZtPKzfXmVWlJ8D
uAwEYgKlSAnf4kXpC9SO4Pls1C9KXNZGis/NHPuJxbiaZQ1yZWkV+r8MAjI+ZkL8JhOaosEm6ZlO
rdpFNZfOIEh2He+AzYujnq5BFfXqog7oS17hzgM7qcBzmeJk/Jy60L2gcQxPqEweMFhUNi/I7mZQ
0aX8moxGl/xZvtB+1XvpCvTVQ+aEATMbq3wp6QDOSP14HSHbYH516m4vwZZnoag/28VQy5y0a3qj
UHIAOa2e/ukUxgF7vhuo/YaQayQ9ye2c5P9r1EMk1B3BETnJCSxjxvrsQWRlbW2mBV+9GgAu4s+t
s9MKm5P8MQy/t9B5JmQx/lPSBgVi3nOiUIgHy7KEwFlktROZ6G5lXI9aZsQ938YBERcxH2a65p8w
P2235eC+k3Z7ZfbrTl1Pl0l21gw9xb4K8fn8IRzZ1et3EELqtijklRoex3BmM3uafDePilrlGwyd
QbhRwlWISpHtONJMgbllEfhe7w1zRUTiglVjh35ptSW1mm4pofXjabB/VG+jTGsFJjZ6mL4REZ0n
QXCcYQVADc+Md1t0CVjY58/I9Vj0RhYMImTdTETUbR7iJYJ629WJSO2kyXLCLXGLw700vOKwPFMt
Wd5w2/hxZoVxENnfjqpNAQRrDu5OwO5gGQ7Q8wjUkLxt2CFuifJZaGPEdIDoYJtSOj4OZzM3cg9E
5XdQ6Wsm+HSDoDx20kI532/4wcM8uLL55wEDaJ98sUc+zSiGA5yI913AXX06KNArAcSU+HIfdzEL
K/71YODiQvTE3HbLRAY8WTvpW03w4osS/wohOnnu5fl85qUf1ijSuSy8KcsO4fpqPZ5KyoT13W+2
D8so0kxagfVzSEGu2XjumbJdpdIkUrP6Exfcv2xkEYmKY6Hk7ORSaC6auubRcLvXYqKB4Avvu0+x
oT5ypbKiRhQCcPPl4/uP2ud9/XPzFJ5dUxgAcWHiqlMmI7wkMFN1JXJfyBsQMQHNQX5m4Rw1ZbTR
rYVv32czkvvQivpWmnsmS7LXErUIGsy1nwADQ/CLcEHjUniSxVLuqfUrW/r7UKzJkAIed1l7J3Uo
r4DMzuYiLrwqyrEBTGV2oRuYe05AB1mss3GITpO+jiAT1r4LuM6aCWfyinaQwm8a5RI899N0dHfD
42m5V85JNryOgM5JL+GGpzQ/sr//NtPdMt/qIarUhvUIHevNBZDdJNQ2ZGIrE9PjFPf1ZqQ43Q0P
3ayUTwhECd0kmDl62z3XlZ448Hh9+WkMVCZL+XI0mAtYi1TmnSs5VueX6ARYGkmNnr6wiPKEJp1G
9wFu8h2R4Pkc3CsbofrxSnzlSlmzj1UBFH/v8FQpyAJycIHVl5S6NAInMYp9qx0Xqf4TjbHWIrv7
lbHS8ljyYhCQBUDK3NPCkb8Ht2/iR0gb708VcAWgAX/PXQKCKrH399ifTyF1a1SvdOyKJvZi70xh
AGBaHpH7J9KatgBvW5NwUpwK6qRRS/Hzq+7MIcQ+2bmMiJJC8p+9P9b8j0MLO5ZjGjkYMtvjXkX4
yVbie7DkTyFVXNq+tOHrHeLayf2I8khIIq2p7ai+57jzWNiHOFptXv1msxPaHNH9A7xgSUVFaosR
DsooyeX1xTmo3MjOuY4U7oXQb5kYnEkO6hfh5/sb8cTBOFA1GJntbNQ3Srrk9LYKIPjf5S+6UneZ
SJnvlAuvkAAysnBHOpAJ/UptgT5IUkPIzjs0AbAQM+ClmTkcLaoqF4JOfxadtIZoCJEA5RsTDcMk
URvIScQhMGtUWnV+z5Y1zAv6cH1QH3d5UQm0TjaVREV44I+lUGcNZmd3nLUGlUzjzTIB5Wvsg84z
XRj0E7kZ2WywwnSvCD4Z23J3eOcbQN1jXZchlDqsWte8nANEHZ4DBmPbs5dJpC3T047wD5fjl3YJ
8kWCfoiQ+5hV8eqX5K+BdlseSzdLdwsU5TGcgFz+ZVpKI2k+Tv+ww1nrvmfTQu7DisVp1S+83jON
A97Vpmw9Y1hntnCfao2Y0DRZYtnly7X+9Xmej/hw4Y+l5i8mSnSv8NpUWUyMWN17IbM757H4n/Gx
Aez8JujymZTWB5s4w4Iza2oyFRcsoD7SlSkhfl4XAu01zwHQEKQv7uZBavIl18KPmWlcqsqpxXAH
JH0ylKhAypfRaboOrAWwyzqqcMDxgN5Ps6FXPOm8OdjZLyKCfTHoEFl/Ue7Bcid6nUZ6VqO+2Y3M
FhhjpmN+QlI+3scVfnkVyg1oqzeKybHzdH2nzNP8ET/h/Sb51LKrSAlS3HfabaT9tKoaFkjrE3H7
W6/O1LOvwQK0FBinE+Xm0sB9AUHawmQzBgyNE3ZMr5aKZ1koP6fjw15XuKIG5rSJKWwDEtILRnqm
MlxBlicB5vgh9x61/St1CkOJ5OzrV0rZ7iENzHbtXegX+XkgDA9bhZDIUK8HqFVTMYMDrBXeH6Rz
sVDwtua7psGVHan7M04zaaInIfPjcTE4HVbQvrnG3s1NYs+8P9cWz5pagX0D1vqOJS3bWIM+8yPo
XTTe198zYctVF4xYoEaqK2xtx/tgvuYoUen9K31UumkCXBuDIYuwCGILGGexs4Hrtyr5W7649DN/
ntJ6Dat/GByLLP066StKoq8ESACf7SFb59WFebxj6uuaVbVL7b/i9BDY0Xd5MhUDVVLVZXYwCKiX
QdOfzFGaiBwogDA3fXsdY0Ebtgu3aZnPztZljkrmtcwKqGNvXQfGvZVIRloPBGOuyFvVUz5O0RBk
FebtH55HIhLHQ6/3+DHpLawNbIG+/s+WgtsQ6rxqM7L5OpiRiFTwQQG9EYMcqWsR2CpXSvx1FzHP
QXxhTCrD0s73mQkK7ZenTvyN2B/CVQCA2KqAFSOILJA5zF8FfJfNVxMvcYlE3vVH41RZMul3vXlC
1qIt5aKYem4mlJvdS8danrTtZ3lVRDUKdWLEzNwDYes18yYp1kugv7f9hvb3txQmOhL1C7hBpS/O
TxLpZqANbAhzmPqTLqaEcl/W4odj38dwtpHHL6dwhdxRm6kzwmM5R6TNCZSshZhzn1FdWh33Hz/k
IphlYY7apjgu5lhxv0lB7L0Aq4CxnbJYmjpRhajSyVpmwmMqkmD6jw9KDDxsAeznce97J/G+Hnt1
sq3aZ+djrmyb0u/8JUKgqdFPl6eKU6iiZccmf5xhQSAIKRcgcvG2N7O3jQI4oNsbRWmF6dRgJWv4
HM7tCCEslZUJ259jaAcNoRAdxbXlD0kMfNageDgCvgZYhEjGaB7BxSTMC4zSpufjtUeZmb6b45TU
1f5x1KrvqiPkrltv44qUdaRYfG6EPp53May573mzWnz7raGOk9OjoOYwwtHnwGs9FtgjbdsjuB9k
FgLyhW+C9ADewElIbk8JQSmrKxxaR92xHZSrYIz0HqM/GQnTxrEbJ8uXzfQz/OwgV0Ybb1kxaJyL
+Pa/VAEmo+jjPjbrxy0+2bQaju6ZJCxsM9bUqIF9TlLpPucEOFL4dhPiY1GobQRUEmAcrfqtG6rc
rQnSvYGj54124s3TqQ62uxhuRfdAQr+dZXbvQGa9KdiD8CR/UzsGoPhAO/5zSKSJgax+Wp/0cyB0
MnygoSAoo8h+IsqLowrtq0a7P1k4CTtKNDpCsXea1nJSFjrSDFARSurEi6aY8dOlVtQK2cCL8MNx
LnRydACFLYVyQmZE70Io/wXJII/X9UVVWCDRa+Rq8MZlP61Wsa0Teiqv7e7DGpPhykbS1+tkNzuz
IiL/EZEIJzy30oVOVwFEMAN07nbxsww5uOWxfKsJdF7H43dhD2mGt5iWTRfbr5z/eEkFw3XIkLWk
KjQttz9F9h29jobjHBynjJ8QHzyShY4rUGXvQDrS6cybSzQwY+9fGDll6Tw5ITCqol3ViHICdNok
ileTrL8CKn3m96OB/OWqGAnCoE9iRV9z/WCwx01IS1CVW0SOX1BaJU3BsKQ0CHt1v3WyQpE3wIH0
K4ZfBxsANdrSBpgnHOaicsz7749w+MVXtiW0fYkUMFD97vn9S5oaZCOYSyCv4bvJBTEZRaG6PdIH
uFs+Ywk7Eyx/NQOgRroaklfclViDkvy8jGIN+pdqPczUgKecHa+G6jhNGjuty6WKwmwLymJheDlO
rUKNu4h7iUKTn5bSh276QtUo5SZLHN7oDTkQvxEJhWvLbRsyw3PSqjh9Pj/195gOfoWe0F0nDFuN
EJV2qJWhWfFakgWJERbtmcq8Zstg8jsB7r+x7eFLAOhmIiWJsHDG00wOLZyUNh1ziNxViAGxbiD+
41o2cpPppnReiOfghYJVVq8hm8js/m1PWIZhoNT7cnLZNf/B4Qn0OPzjR+CmFsRQYpYuJ0jJ43wo
D0YiR+SXxy8Mx/Vpm5ly2PCtavQFV6398ha6Hx4zsTL84UdM8wBsoWtU7B4u7wWm1eIsevWWhsbF
F1Sw7yyGZLiPMxz0I+rCThjYI/y1m/vbxUEeSEXPNZZbKD+qeFAnp0BaIF0uK3xQAOc4UPJrBGZw
D9ANAZ/DqtYTbJ2788chDRbwvNw+9gq553zs4klRwNOP0doEqA50ylAqOK+psGsxFrkvtOaaVBHE
lKp2uc7561UR5lbrFUriIQ2i11g2eqAPOu9XvcXi2Tw5T4itLA0MmcUtAxk7ccq5BXS61yE0332O
3pYRmhz0JFkZ8R+6IwwScKXARiWE2ERPpBPkPl65bUJ/o01Vnjb7PL2+/k2jLWcdYZbTj0Cw9BK4
u14hzvrwzzw366B476Ekp5zfYJo/AtsjHI5rDOSvI8tVDgEqB4UJmlwhWw7098n2jWluVK9hQLLJ
hQVJwGUPbAyRohk8rcbDDzZOKaP+PtFlzRUAaJLmqm+e50ypPYNI5UuBE8tARn8/fRbncHvipR7w
RBSo4l2l61IOz/YJ6jOR3zaz6yo0iXo9DdHV3yxl2PCRqt5ErirL6x2Ry/HxSVP/Sn7aUiG//CyP
beKW7qD834tUk9fCvgZ49vwhU9ohTW5MqRoe2fXZwjHegChB6iyPBDYNBYHOlZwi5MVUfKRN0OCQ
9U0xvwAI5CiP4P9TR/PZg7YkLfBI9oigETpxW+ajDrQO51fHldX696W6dlnLc7fqjVvLZQnHN6sb
sd8bkOc9EBxEXGVYB9e2zmnlsgasNDYNQ/w6GP0Wf4wtzcdwE0Zfxy7VqLaMBzIKnW3hbHw0g0hK
mNPOlaEjgzI8uRyKbc/YD5bT174bV36x8DN85GfYIwy3m5vwvBj5u/AQ/KJJ6Ts4LikFmo3lOVE2
fDDCcwNcoqDiHq+Vd/7O8Y1uk+K6YRKeKj8nxVaz2Cx9b3x0jfetRgkPmekP1UrY5yB3l1WEnj6T
Si8W7edCgMl0IL5fCZwqmFEbE+Kxgg+poSSCfzpQstF1m8969XksFbOt9sdk2bYRRmJbY/QNr4j5
+kBvYJbwvo24+ziQuZBKDJgBzkqoZa1RJG7OFoW/LXF2Bn2XYfrbGn2ZB/n3NzsNWAko/NaPh5bJ
B/a48vJ9AZ97OlHh7NlW2zCwCHEzlUsDETeUK3c+1o44f1To5hjCzkcP2F26EMsse+mgBeJu6d6k
CV9HVy+mvjSy2X4mXgO1QcXeSbkacdNfjBi4Y4RLjDh6opsTJkHt+IGeaJRhVc2TO/M0agfEEVrK
AdAnix8/IeTzYWBAvRCjYZm8Enlx7RZw7+YkcYe9gIs3Q3eV2G8BkkgIYT+hU1Zx3Uv29T8pKyw1
CpOycCWZ/bHlZfMGruLRVdmXexNWcJCqwfTN7C9HfHTqXhWQW1NLaP9dq3MkgBUfIObJXCw3jFw/
a2pq6jJ02S7w2myzQB3Yce/8F+Um4wqck7GaiM7dDgJe6bHiz98KmshcwdIpZQa3kgyiTwlTXRLB
fzjnM3fyopLruRCbdNaA9L0Y9Krb7d11I6sxb1KGokQMFOOZrCGXMQIhFTq333CB1/lw5jLYf7Iq
DQR8/nwzjK5Lc57FQaDLjwBBXTPtRUQHJCgmTr8hOPiP7AnKrEhw/yLEnG50zKxrudqMpGsbxFm0
bl9oP2nF+XHrVURZjhB5U7EXYes75PEQPBu45k6C2XDrjFk1ihffJE/s6YKcVdtbVcP3VNIxi7a3
CriPJg6BMngd5DQCw8VHvlzFCepE+zENe4cXoVjdTeAX5+WPv4C/FFhFTPTLKk5a1fwCwWPpF42N
cKMEsYqwhrUW/QeOP76kpEyrkCAO7ZpY1skrSt6xTz54454KBle+A3SLed4dRvcSRMNSBUk30Tv/
flMSauQlfIvpmc80VIDEV5ZxK6vJqPQZk3G1qU9HSTNNy2ODjzXBjDktNw3w7kJniSNdPndfJ81j
+n9omLcT0ToeAa5MvhrIjVhtMkvKxt2xflZ5nIFxvBiVRckcrU5BzDbge0dim4ibKsTJRcYNZG/b
9ELfh/LmSdTMTeCHONr0p8EE8kzzDvfGYhyApOhtXa+b40cpQOghlJ/nxw5p+6C0Qk/NulPhQMf6
OGyNoTQia9DRhGgu+DY/e1R54bErahS4jx6y2w1hROTBT3uwkn0Esi+4GqCn86Feeb72wsQf+iuP
KdfhqELVoVrhTve/CycIz5CgOuW6E8xwofJQDog0TWiakYXbFIP5VEJOzjAKEwM8TNOyQY3PlqgG
j1XVQmV8rTL2qt1vXds2/oyZe6clYklrbOwZwwjM7YLHrbTVdd4SimmEx7QMqWKknkwzhz8qbJa0
XFYsNRWmPaNijopd8uYvJN/qZGcAfeQxD8d2lRUwpkMe8P1JwfMg3iMs2MQIGg07KUvCasPIlUGV
0eIsK1upuCez/eHuBqfVILfCspQTy8zPY+B5MpJsifRo6K0F2TQPt2ovkAw1sN4cMFUOG+lcXJZ9
5AkwHytLy8gHDriAUIL3OYYjmIDNXNP74kT+BODRI0CyWi0LQrTkPUdvkTyeWTDI20V2sGQnJuZ4
CzBklJMIo5mb0Nor1qXz1VBwrBcCsutDntSBE5t8sj8jOYtrsEsGPeKRRoSy+g5u5R6RO9w9awsq
ltpmZRd4c0EOghHQxoPXux8OXXwWoq+EoxSp/34xS//w/uUn8mSehcfkRv/OQkMBqiqm39vkCI0U
q6tSCfgn44IK+UVh/XTvhpSjqu+orzBbVosUhavQOBXsKXnDetTlh/YQcds41U5pYs7MmzQ4I1us
2UNX1MyIn4GLqV8jiV5ouiIzgiodm3B6ljdXl/WKeh4lhHlU8S5iSpJGlQqB0tHVR9c1EsDVIHRB
B2EFETOnilkLujdEz+KJ39tDlndQd8MCwjOA0aEaeqCW3N//9W7CCwcKdEcCRZaVppgcM7OZDSNn
S9qb5cWk5XK9XCo/GFHCvnNL3tPYLZz/2Ol5DMB5YsOF/wdrWsQbMXw45bmcNBxO9SBAxLnFfesS
R1e/Ey9cdMwD2d2bFD31d7ym5yxtvaDZVwRFhnRQDmpuKmGDc4IKdIr1hlzAqphmycZuxSogl0B9
bedFTUnxCrhc7iAyPr1pxlkOpMyhpUsnYNsSNt60AWsWuwNhD1tdT8fiFmzds5VltZ0PcRImkIka
aEDtD0mH0hHQ9sW2cs9PPZ488tavw0a9NT8JDDtuePsf9ICdXBPDZ9xGenL++gB9XiRbybAQfKzG
Jzw4vepscN32FhNjKPum6ymI2SeQy1pj/Bi1NyaHzVyh21YO2r1rndfS8S/XR0+HgW1g0Soer/Is
ZfadHglzRiILC6cgcc6Guy9SP2uKCcn23RZx7bMtzzdCxIWprZPcKhdXEsqxDZOjLu1yf8syVprS
Oe/MxoE93TOxvFscln+uDAPlueudxTelVEK32uGymzWdsKEUNOJJu6yJqsa/bAl3wTLqqkRcGaW/
zVyDkngjLt8YoFFo3tQvyj0G2aQZ9nDiXzl1V8sgT2bU0HJywv6GXGRJMWqPxr3vUDLDbTO/uV2S
J/A5vYr7cFWn//gjcE+Ze2S1vlN+jph+Y6bENxDEBENQfkpWjCvse+b8PfUvtBElKN2fF0KHEphH
mL8jxEaV9M0ly9IgmeYKFks7yCO3Q3kKp5/g4N7Ffia+KW15DhdSkyvlbcjD5SKDMA9civxEPV2R
K7ICPKKnxDmjVmGm/IwLaMHxb9XQ6kHse6e2KLzllE1hPQkctt2UI2ePCWydkprihYVnu4D/Ubx3
L144YOvptz+eR08pC9gS6MXDAb6DIPVXDQ82zUXFLSkes1SnhMkYjWAw/J8IrrNXmBdkUbNMk6bk
hHL9D6OoHxBo2BF7VnvLJxVDu7eS/EQcuZIhllxMol8BVDmOcBcXqG9VsxAmv8cQT8+1ldc0wQkc
M5+f1SQgJV/z/UIEjB8eRCLdz4oTGVX/yhPdhSwg2RyEBus2laBJyhkRZfdoJ/wo+JZ0ayKxI38s
hhNWQP6rcopJZyHPGxR9XNxUFg/LeTRtyZt7VU7zxoD+h+nMZd5NDlNIG2TAv3l4cfIfRX35nepO
wLw7xXhoNBaCybJAoiUny6AfRh7XnaZZ6Ht2YU+iukfCxKIexWj0fwj6B1Uf/fEfcqKgfvyPhbFc
wMR/j+BgNbfYRhImLAmm2dQici3gNh2qlv8YMyaxTht68MphPOYtGXcJ/6QLXJ1Jt3oUgqhSqjbF
MkegtU/85Rsznz+Ersw6WOT7G8WLYFr4dvaV5uR/JokuXsLUbzHJUr7coOihAkd2/Z5tEAkIprhq
5bciaT8Vh/BWLHuH9OYYgalcUKCyIZpDVNJA4VFnQChjVJXcAzEUzwr93EFohIOrEcoTWNVtUZjn
xcYm0mFA2QMYOCarx9y6WCXO0tiT7QX4WN5e3jOLf7s5DkNiT5JR5aVgsSB4+l1eQdE/uPuCJJ5z
cTiXwGSkL2Ip98cpVmzZvx2gAtA0qw/DgPYYv1DBEwlq3xU6V5FQHcWGYGHiwCk0CchDgw1vwtkC
WGomys70e/bAgrdNzzLwiBqtUi/kTcQbdGcqpJedK+3tJyoAg+IjyHS6GTC4n/TlUjAUDFIAlusB
JM9X2RYF8Qt/wX4PVE6xw/OxHK8ZlQ5D16C0C4utVtKxejIREJ0GQSZo3ta0l48xgBwltHHpPTkB
E4ZK+NWSULW0/gvvfDarSxI3NH6yPPWAijWugKUCfeorRkoupM18n1JNF6QGDg9jq1zT7M0VNdbO
AiSAZhYhFRe0NKV3HJ0Qs0On30KTM2ZvrIZ5qNz3l3mFMC6/GDAZEviTWAxav83E/s++R8zE6nSS
7TFUTCp2Rp+wMoq0eKy+Hlo1R85SXKdAO6gOW9zwpovDWkK8bdna+Ii83CrVi9+iLpFNBZz/LrR3
4nFNzM4DgQijmWqAkjJRIP4SwPJpeBsIxCrvFSDE4jNqUYQSGpphKrentGKrttPaKPq5xR3QFDPK
iaVCr5qdQsKVOQE5MGKllQboSuDi4dEXmuahlgCGjGsczT4Xu8ymYwhOAIwFwh0NkbVB1oh9KO6B
MADB8KVVt4RHl6Y7v3J8bqB2gUkk8hhlBlOGp9tT0S/eUANbeBdb9bi3yIhJcaewMGEoGV8O+Njx
LdlflCUxoWYqLmcpagLpQ+aOM3jlPhZMFRgdmayxqSA4QEGGyNC12zzSVvJfurmaFaOvmWtut4Z/
tTNhWMajPuGwgK7rxxqmT3efzF1sRFWjWgEROqzI6MrVrm01o4WvtpDsilGnryxgrL7oW/o7+BIv
yZkAYxQI5m7oYTjnku9QcgNPo0Q7hEJ5HJc5havdeiAhNhbC4jqkg6UuiBZ19YftjcY2+D/SyCS2
R5zrt1tVqslU/ZWv3qofJKt4s3xHtrpHHgvLNTvyDC0PQ4gi9Z5kS42NM9Nkc3okMearHSvUPSEW
hj6GP1ZZkp8N8Sw/0v7vGq6BWM8DWSmknpysMphQ1iC8DCn/O6bhwW53maA+D+L5fY02lP4pMQZk
/iNaJTZvuyd1tXoOMjBaKvsWu2nQTMMAdCr/cK98vVL6fKdD4wXU59uvt7xD8pPd180xcI1M4/vi
m5icZMlhpPsp4Y0LmUXQe5SnZo6y+LbrUhv8WiIqP1yj827e7qrVOTuDd/gHf11NlnAI/uQ/7dHd
cnTb/c/tNTYAdB/w+uKJg1rgNn1gyGzEudeosP8bUor9ZGUD14Yd6esRrx2VWb1vjXtYl6W2KVpV
GfI2SqJsHLrns/aVy7bs9eMqN64D1hcuQ+edrU1Ishq9GaUGYcCr8yoW0BnMv1SlOkQLZLsSB78B
YZUNYnUF8gSg7S88PuPHk0kkqf18cdTrX+fluo1Yp2z1qz6ARkM2VmBb7Fwazd/leheHS0OynTU4
lS7tyaFLdbcM5WvnDqpWkHPf2NOA8rqYiA2W6y1OH83wQvp+NGFPf7KmQhLzefoWRxzeolW7TcBF
peVteCIiik+tBFrNmKDCrhzucowHcBWyKGQMldSRtyeDS26gk0ZXD38/SYfCasZW71BaFhP5KDA+
7NGkiRIcA6iOiD1YWWvI73irxjSYD52GQ0xyMEOD3XIySrhknocTl7KxPXTp3/DHlFYSXWDfrfQF
IkoOMzwibyNcXxdLUUPAAknLNXc8ReZUrdfDnxy1Oj91q1uM3GLgLqsL/OVlvB9qetIeZiSjbjFu
NKqXZENXWCqW26b3GJ4dmcSnRiKRJnJd7Q76/k3t0gpUv7+DbI/U8eZjYK+dhDrN3bGNMDnsgx1B
tkYx5R0nLDlSSmZ/TRMJmlE0kM6WJJuG7AwO7fxT41Aw6P8szrjn4s4Y0t6AGfBipvDigcoYao0l
XLfFHu4k2aeZIpUUys6LLld77WRfYOJ0Sxdo9H8EEFqqtLjuWksMRnvkxggvaPT9jM+jlBluzkMd
ed1UQ7x2AeVThm0wbv7mh6lkSKbZ8wZu8V+kuwN+ezQAX9errWdz2JltA/h+FiNn/pGrG0PiZNzo
4wSfuHY5u3naaWIAlF2zE4IuMpDOd54aPoupmBaeOS3DpUCa5FclxKiz7DZCXmruCcJr1ywZ/Xen
z+hJKgzuHflNp3zyKRP1bs7gccHB2bKfIOPVWiKhBhyvThtuByEWOiNn1cQBRqtUEo686XDw2r+3
FKL50sXQNgp32Y5NAGkviPp1SilGgf+gdlwmGbZzpq6RwiIrxCiaeRqJJc40/CPKXCOW/38UIcBR
VPUcSvm4PFpBXOWSEv1B2DMcW/DfiXe0IQsHi0iYzdL41BUCZrFEjYUO8qAGJTwdNX7A4Boh+zpw
cgLvOyJWN06NGmc3KjV92bh49Y7AgCGJpLxHoyfKe+8UK0oanFbA2I3E/OaSuezpbk5S/mYe139G
0b8wtbK5N1+StZqKfTwhKw45RjBhVKUGs5fHWGhc3ybRVQeWOYU0KqN4t5iySoP9xfiI0zFNG/pq
R/VcEEv5E2TDpSG/oO6KYa7ox6+JPb6yqX5n3yxKkxz0RAtoCMCVxIDSucUZ+dgblwx2NpSoxpoj
wodo6gRpojDSx2I3W1WmynvKkOsHpepBbBHhEmdZiN0nGXSSNtV/yEKsoDSC9RbFttN9RHeNwJ/r
IJMkcNcv+t+XW25D5ZGI6/yM/Gcxcz+aO65WhbbAuXYyFDCoGKFtgZkY7Z2YuQuHmcjWKI0sdWZZ
k9OW8439Y2ybGFVMNvyTc6ODa/lPC9b0NCKegcGH12UIb4Pi5oARWVxWfd5t22SQbiQNNmeDNrae
TiHq1e5zF2rmsGTctFqIBBFXbOwYQ3RZn1SAwR3EbDYjr7+Eby8isBbUo7SVBxd7p80WVHK/VuEL
zzK1MZ4KhPaMuiJQsvV9A8z9uHRD4uzf1UVO25I897nZaxMa77AIHJ8jfu2xZyevK9dIEmI6SEx/
+eNSvBjDevMy9TFsek/YV+meOir+2VLgfWQ6hjoRKopFEDpUweEeuU72z+q/pO/UmPehfBvORWae
NlsQczNC1VqTkcG+OtoKkgb/ln8IY337AVLPjOxUZzyYdY+Gqaz8DPy+wOXiSV5ZnTBESAt7VkSf
8q+0Vxcajq/gshVdZm661qymaXg1AR3lPd/wiDafPRNlis9Ichkdh6/WY9k3ReMUlmWF0a/cnIjV
U/p8lde2lciHhjT04/8I61aRcwo/qYZuK5yYr+dFOzvJoCh+jLD7Rp3sr5ZSdliFfRclrXYdLwux
i5Xet9RQBRT4+dFzDkPJ5niqylRcMS1K5LbT+Y7LFDeUORLa20ExWoEgsqRqHOaU8SbniSfInaVv
xXKgSYIIR6Yzn8QavZnoTUHgnrjhBOd9FQzTR3a9t5MoGXUqCLawFS1rPLrZQNxP1MHtJ1y6tz8Y
emO3pODBIzkeHc8fIdAxTYnnBw4CPefo9N20rkKWT8NGsDsy5bCjuHIGxV+zBUvsFHySyViovj0d
U9LMiH7FaFFSyTQMiSl7QHN1Th41m14ISNfYyakmEfdEoNL3NDHeLx1NGzJkJByd5kLm4KSCoG+0
UtYpcJW9IxsFdHoEAl3Oa/EdiO+WGiEmm7E7tHSYyaoGnfrZHrHXOJbWyZFrtOa7EOjxQ289V7xW
0kFLz/L1ADeaN2Ut7LOKakKsb6gtBp4mqFqmPoi1moSngFuW6u7CDAxGkq7x7R6vOgMavQyuwNtd
U9JtYngUubRuRvsjeZTz94W5FkzGazo5RXmWwL65ehqHdoRdxXJoRD5qq2ypBnZ9esJO9kSbybc0
26qtEhIAhzQ3lxDSN68qHWkqlhsUpavIveLUD4qrFvQ408A7mMpTAne0JRbJrGX5ggdbh59ZH/P7
MLd/L3YsNpZ3DGNTiKevM9RWUj45nzAU9HuYGNQe8GR7QvcL429Y8bsNUxNnL8ZUqsRzZfwN4SmU
Rc4stv/jkRhjoXAEDVe4MFKOhcILFrDEid3YC6iEvZBJFBh54P7og9oXP6wrlJIHtA7YWCvTFJJ2
1qUy6Z23awePl8QEFQfJSVc0l3Voj0f2GmJVYALPQnMNXJhX6FzaDodDnjHQIosAFOzQ/ECnMehV
JGoru4xWBGbkNHSlYLjA/xTPGYGZhCnQZzCms0fD/Qy4oQ8/CfHhsKs2JGCZpRKrSkkmVIwtbmV6
RcaBKngxYk0y9ITbGAJqiy01p7DXKQ/GTdUosclbuASQJxjBD6WX287vGKbQ+ceV/YHy4toPA9Br
JIn4fftoZYLE3ZBX99XhmS2g626v79dDRQVQ6ld+rMPgmgStivQScowRxENR06DMjFljM5MLMd/Y
aZa+i3o1AjoDz5BgTuApAaQn8uiVZouO2oijhWb90ZV36NVi6AqCeTSh9ycmRFTIpUi0voyDfqz5
8q92QPXJgd0lIyu8a8R8mMRtHVpka20EiymUYj5I+qOY2Eqld+lFFU+g+mnfg2/kUy9sMvGwvCcb
f0vZCU85d33wVAxlGMhaGFQ6ATs3JGboCC5mW5HEM5VrdkcHgW6FDITWDrmPgybOU0GGD5ava/Ea
SeUPpoXGtx6qiKFkna0L+SZDMnd1kzp818y2I3FXy2VFtbiJywKM0jLSierDDW+E0uf97vOTbc4z
sSjtVRYEQVInJ57dbZjTLtgh2rATHXrZb5updOjQDM8nznmNlTK45oqdlo2bnBM4VsgNtP6elEOz
tdE1bhU3+5MKMuNQs9R09UqBGb49tWrC65QhiroFBDERqwtcYSy3nsFbft3sEI7V+ro2eCFrk9QS
0VwtJGwY1KNrLKBSKtmvCQ2tho6ta85XNtMv05iTM9LQlX7imT2gS2gVICL7RDjhJu3m4YtgKTLH
daKRBnsX8GLTcsCYBx7aNl5exjTT9Jh77+Mxg9M9zZSocb8EiuSVmWClYOIu7AbAbxrmVYHKsL0j
FnEjByktZ46Hgq5x65qQNgfaaeFF8W/2KoIFtyeWoA2R1KX3SmWqXUtWL/D6SZelMCeayU2cmOXN
/Bml3V042sSEiwXaSnAFirD1HcYV8O+wyVQZyqqIPhFrhCxcao0Z5+CzUbZbNRdNWyexm8DNSMOB
qaKP3ZBAIis3+5+1nnB7eB4COqDMYx65yf1PLcFT38aJJa9D/xPb5fSuj0WjvuDfZY0p1ZD+G0us
s65We78iUBWj/i+Urqfvs+PSiHFBdKmP4Yi2zyFUkUBjh9LgT4IU29lF6zdfSjx14JnqrSPVba2e
UvMXhBuDfU99kYs2MjIf+lQU3Qj8jEq/AUnqZftnDuuklnAofaKuU1DsblNp4ogm1DRa62NlfLdT
7daa+HoLeRYMXfXpoYFvEYPz6iGDq412Q4jIqVrzyrBQy0csZQ9TujyqvO9MySDendsI36hIkEdR
9+2bx82Ls36xC163vjy9Jsq4fsXy0xcJaI64JrIc+ndG7OSX6T19HmLE6ldYvV4A8GrUTSsSQpsE
ndXD6RvCmAe89tliSklSctdP1DhfuGn0kzgPsir9yL8ZsUfMxapuM8zFqGFAv7utm48L8qi/fa33
ymMcxPAci2dqzJuaXmwsi5PhLvkE7J6X7o2mvpH6HUUmRWYLktsYlVVLfRYTppgHN6Bal878/FNb
3GM05jxu9clmBRN8c7mQyybVBHdvg5erVPbv8Upi+2UBVxNcTjnL+z08pX2X6tQeVgAYnrAGwl53
gwxb8kO0NFkcL/r08PdMWHb1dNz4vMuvjmwXpQ4a3HZFDrMsih7QdQmyOzqPtNnAQwqvgtDf6B7V
9jcmxg4krhcjKHpIsSKXAkryI1tIHj7hgPC9JnzHXetTqxdQm1Gq4/oz9Gf6zjXipwKdkU5fWBsc
0ehmmcEGeSDlc1vWG9wKvvK+g6uVzU81GcoWS1Gh3Eyxz8sVzRgK0vdSgtgXCvX7G3pvDFHt0yOk
BHoHPK6bh8PhkhHkHrlj0f/boaaHT6GouWeaaDg0dwp4wsgLY2JNdsdvujMu+5qbbl1g2EliHOcB
cWUMmlM7l54Ym9uMa3/A1ZDSid81HN3fJV+rzhVpS9anr6ackssmofui/sZ7kV9pN5hv/LDzoJaZ
vQfWSFzyTVi/XAR4uC0bWjiXX+GgPBYgq7jYymertbmbrrBBQUMmpcJ0Ymj/XtN6Td/hzCET8WDv
xEQOvdxI0vxj2HTGT+eKlVtmXS/aiBmzwPEpEzQJxYbqGpYItBrTjNa3XRmRbCswcW7/zX6iVR/O
/3ozCcabRzCxsMgulCl/UqYQacI7M/P+MqHCYEnw2HxZX25e6FrkyqW4TEvN7R3juIhp2vY4aARN
Z90dQN8c7aF7LV1fPscogV4FOn+5aR16iOrWJAYYe06mLRipZxqKWRSxvXwJznREPbXdrXH/q4J9
bAcWPiO6WPZEmKUI3h5Z97Xdtwnc8YDcbD3+RQ/wIGjat3xdLtHUqC46dpWGepGlZlZ03O5xPBuL
uDp0BiCRqaAglqmVvdNiqGQ3q40p1kKCf2bokoMWvfGTkJeYUtQuwZ7TVTUXmovW/jAl8fpD/Zw8
5cZ+kSb6qTw1npZFflrGDeG8HcEEfgDmOKg1JNdb2lr8l+flbXvgXhWEUnYKnNQGo+OjZmWQNmfU
8HiSfHVXaEqT+7Mf8z2AbJcNfesDe+pMi3LHFkhFfVRBvhgLdQOheT9lQSZ3gvusKmtL4stD/0Ty
nklOr1OdGVIv4qAHSYgecKD/9MLi0fHsP0/AECD/yPwvOoITeXVTsWrWxvcBmVZfFx2qN79smbGl
W+Tc/QXCwTuvO9fH18xklQWu3oNZ3tBbyzGEg/JyNF84A/9gXTM9PJKTPBVrEjlypUxN7t/J49Rn
CyH2tJ5Be/etMedjMMcHmdNo3+81GG1tqvKTyb/H02ItwV+KQJIkRmDTlCV55mdS7Vv9IC7/3VmQ
lVKMQ9I+ZVd/EMSh7OS2DZ/WnzksuznnYXBGKnT92Q0nq0jSwzDaghEWsvFKeNZ5hE1GiwuArF8I
+oFTUrbV2t+mLdcKxTXY/ISzUSWd8TzHywTzJLRhL76rLh3eZ7BJjmDkCaxVL+Sw9fSxwUGy1bf4
7sNK5Mcle6rjONBqL+kuQTxRLfyPtJCyn7ZtOif0omrzKM0QZ3uQa9MqZBRuyPXLFS01oIRTUfKY
5uvLsa9w7lK8Yn578n+b5wjDIoDOx93+mRXgszVzDtcEPgsdb3hTgNePzeXTWd6Lq+Xx89k6XNnP
OQEP/Zt3SY6p941hQaYEKRg7RueW1cDB0aeucjQ2GYd671sSRgkcrKjJ9cSVfZJkhd3UGeawrbFW
6Oi3jRuXELWm5LFdKf0rHSb3gx3grwGnoJOs81neWJYffb8vpUDnrQsE/8OOajd5igdEGAIYUtMZ
V0deBJ+t9bUjvR5DG/1CbD4QbEwPxl4vtVRB34ZWQVgH1Racwr+UiVxv7bXLWMDV3S+DTI/10ITx
ZHxu+uNSzEIe0IkdqeH+e9ZXEFE78iLC3nzZo6PdmwG3nM6UTIQ1uQAhJySeobXslX9L0F9R9R6x
OiyOq1+bImsVVLCEtVVVhH53OAZQXuCdHERmO/q4yilFBfIGaCHjv1BMSJSPjeUIFeaz+EPv8Kr3
tPa0yQkw7Gmlydct+gb/sNr73ITrrSF2ATLOnF9McH9EBPp1uo5PW2QRmitvIFRyaA4X3LkIPxJT
gJHulooJnzkDkHGbAvSBC7ehTVZbrihMMrgO/YeqemC9lnnGDL+TC7RVKbom1ClqRMsv7PyJPnc8
fp8qzAbEESivO/NE+b9LeqkPUNn1AStNOj3DjsQHLZoqUz0qDSZtlfixkBm38N5N2X/krC7uKX6x
awzDrOUHBorJeZMuZTKwGpkTFlyO7cAcRiDxpvYDkC8usayROkw3X8SNRfWi15VALAxhyzF9Q1WT
M2RaOU95e0odttFQyrxj+jidyoFqfkP3vH5ysrutQ//IpCPSGY1SRoBP5Le03ipFm6szufVMRp/c
FYdxZBD01M28p9jG9zRlZM0Uumj1bXmcIctVRItLj8SqiYPAPpnAi7X5ktgaKelyWenplpsfbsIv
XePTxpFEbBSxN4GFkc2csHu6CPOkFhG5i4AzJjxgy27ZeFfieofA4RAq40S1GmdistDPLeQefe15
Wx/qFvuoveScADnv2YtFKltI4ay+Qjm0JTzP27F5exdCq7GTn7KpNGNLudlDgn3i05U/CvRvRa4b
8uqb+r+7MLOtKOAqZM+DRz8QOrA2yXx3U/bWCf69qnEpl5x3+dJuksSVqXaM2t0fMOCW4gBwZ2Ps
6OhqAHxso6Gsrqy14Fvs9eQ9Q2e6qEEW5QtEr8/7/lpOQRU0LeJE1QVAq9VjC95N14Kcwb2N0q7L
4/L+7Zl1At1KnNQXMRw9fAGXO0h3/lUkGDmhmQQQAwoaC3qYDd8ayQigXb5TKB0o2oehp8R1Kro6
yCTMNXMumSajHyfJSotndPEFWEffsJBLfhUY2cNX3XYuCizIb/Ciw0hz62HS6czfkkaT7g4pX3rG
sb13yXFbR7HUcMeDzjxC8OHrX1gGTpOFUUIkzo9q8b+sv3PylesrHhrAoyee1ZeaC5RSgXPurt4m
BPh0hUS85PQLszfceSqhh8R9Jqw7SdVIKA5QslND6EVfLfUb16TJH+Aupd4lMbZ0GKt8aNGpDVgE
+Lby+4ATWH09U2+jOVHP6fUZPKMsRmuqFgy5I3Bw5XnwxD36WCX4pxRLy56p5cgTbxUimCul36zs
dYydMiZlAoE3ag4iswjOf018TGJv+OaKmzKP/e18ZG2bxyO4D6PY9kpn2LoYroICtCw4swSrOl4c
tfWPiK7YRXa5RPBRXx4Yz+D/WJWjSrKg1i/vfQ5cPvei8NxbdLev3xkkItKclvPOqHVgSeYIaQwZ
cuUMURJP5ZwG5ZQ3iiwrJr+CdpuOdWqRFLri1ZvQVqlVbRTnK7pbBStzCVYlc2hkC7tMLA67LMB6
7CyJWeH4DC+TpaE2yTn1YItTjsyFie0HxX0jIyOTDuT60zTZ0MGGxKCggjIIafnS0bqpqARcJLCM
mknnd382eDBBcvDFiqLTgmGlX6Vl/p7EH0ndeU8aXA5BY6cm/uIsalOi11n0IpD9JJViupvBeUJp
I5Nsu5QPFVCpV604IL5OCRQ37hDF4Pc6MPec2gKBGZ/d+J4GDR2oza/X1mhBmyS+aArl4o9H+uko
eUs5w2euSlwNdKRbmP4sPGk+wAda2CNupU+gqU338nMJv+I+l8eDPetp3MD5FfBSb/+XFtTe3p3+
BHXtp4QFZbpZ6NlDZ/zyHkXYug/PNMy6gky0hRSy2JlXH6Uu7bfI7MS37VbyPdWd20IFq2cwuvus
9cB9XFNu2HzIZoSb4DxO3B4wWPvO6r26MjOQMo6h4vzLrxjorvEhX3gF+xXXl/mQ0up4vIBbdZ/t
rjdxlxPUEC7L8dPez1/vrFpanZtMuDSOakKUnVlnoe7dAEvg37MbAdtwYqsFi/daK1+YR3zo55sI
TnsNqxqsGnLZJc3LFmQsXMcCWlpzLCrt/EtHwlILwoSPdiU6vukd+XehIualWwdF8xLV0kRLCREH
ARY73OJI5q0yidFQdhWR7fVpoNjeJ+sKiYTSAzbpKuR8zW9svBCyF3kAsC4yvwXGUUzFZ2qwHey+
tbD+RLPOe/Q8jutL1w5ZjKIC4fQsOTOLF4wjZl+dFs0t9+jwacrZm5ci+vBTyPcIDifdvhVRmIgq
AcBDptEknCGZ5rC/xht97QZ4XfINCNcqTa12QT48MOEMs7HhX3dsEyTIq5TUPAqgFRtxGI/AIFix
U1eUBqlAFNWagBEwIRlaJRfIx1sitBsME/a1nkxKCcOnjMNKxObJ8ukvEgVQYnH9iJlI2ZXxZ0Cd
+zaaxpCECM6OlRGgjP/XLMYyuRic0L/IMVai2LizRi1AAzpsR6yM3PqSdP/DEskvfLuLbgzMMhk7
bb9IGEVVKXFSbrrVJjcJnnGnAlpUVtCrFKLtHaugTWqDKxJSDz391V7t45JtGNGTlJ3hnSUTyuqq
W/1P4KCE/DNO1dhqDoXtHAkGmaIavJHFGeFDTmjZjX5sj5/kFe2Sv70JMswLn5cXrnfyq1oWouis
TXxlwRzUOQqqAEG3OGMEXpjZqa7sI7MdeXs8XorddwSl2Ef0wbKUci4RzrcbxMp/CVhlTCXrZOuH
KSjGbokIFjoScxpbnz9jB4SnUJJJMdWLHWW8djaBJhHOenSp9DO87L5YqyK5Hg6rtzNUaTP6v+8L
Yhu08Cx//sccPFAuQisQP45N3FDRok56nSG0t9CHWt0IE9UXjGFZrJcEVh4+AoOUTHoWlOdOQhVk
vF2e+ak+5UVn9tahUmMj+2bxO8BbBzHI8daA+JTEz0C29PFoPGBZ706UihQE/XOeyaAMPQm9nGuA
Q5H/OJBJkWAyW56tNHMvEckO4Yv+n9gIctbbweb+swHkIqQbZu0353urSx8/deOX8nL/R2w1utuk
T+bLLiRZCtzoTgBh9jXVhlr+7Ty6Fg0ZRx2q7KJVXTPJJCIz6O9TQKL/MKYkJXiF6M0Qp0tK7Y1H
kUDI1+cZ9g20DeGmuz3KvXWnI9E0xBTJEXPPTlrHOg8sNWiIVqcHOhRG8Rd8bp1nyaK9tdJ+Cn7Q
aL3ylS4xTHyk+5oMfPvKmIs1o0falPhGd2QEg6g5lVSj4zTn/7PxyUUhe8bbIL12TXN8OZVb4Bj+
8nXK8/tKen/zAf8qLe8PbuiQh9s9m+anP2mch8NirI+mEkJcNHc/zu9Cy+R5TdgCQmj+406Rj1kk
C7ffqaguNjEyhRzs7PUmEPB7TM26cloyxgR9aXLyACS6AoD3EfwrM0fNr3g+BGAcIjzipB+nLBv1
SCegHXzPlRkoE6vCGG7H6fxTI12O6DqngkBgMHCGkqqB0liXmZLDe2xYQu9DiSFWQeRTg5qe9Nij
yI2nvfcwLFsX3GX85GlFHs7wLepUfSF4q1ss0B0NcQOhFMZbuJ0vURoJrNqoghC0zpSYTyeGriNd
rtcAjChb/WzdGYgpiTDQpM6oXnQoltOwd2bS/xf6M5QOQSDihBpofLGDuJvdEfFrFh5kcJU8aZIa
77lB6/U7TDDcRFrFZSY1wMRRdhz8dNEj8zJd4Fu0ZwpUijA0qg4LEmy7l7xfYdx95zVN4mXr4Qog
8ZESIKACxQi6r1qpsrv6EAWVsJgaBrZgaJl77lA3ZCC8Jxrs8/65b7cqOLXRKOByRF4kacY5Xn2b
tGbfg9w77MLrsdjLAhp96KjOatz4WN+NQFBSB5+g8bIDzLGnI8vt/E6jO6mVoMmm97CwrfzuUkGS
pkklVzJspk0pd0m+1yC/4Uoc5cmEukfvRSen9WJ9Zrw/5rWN7qiP9EpAUbS23nK22ED+Cid9s/oA
5AMes1GHQXEMRMDEx92+syRVwRusGlF50ZV/7qde+HuaVFq4+zWL4xqezK0tZ8MZK6I6KtNBSstA
czUCE8t6lqdfcIN4byGcEUyplohxrnBBKtXFKfbOh1/eRyQamSsZ0fHIDjL28wDX4nhyBm35vkym
Ccct+87tKwOu84bbMOrpo1oKhQiEN4cQyz0O3TvUdEYZe5cUVEfr0C0Bdoz/8rN6Ctu6BtHbR7EH
19eHaaq7fM9K6yzQ3HK7RtQcc2FLMpZqMuDT6ACzBPgBrIgf/7C6yvzfmyf171LLRU6H7p8rzb9T
jc0NDiG13c4T5VRwJjQRihsclpVydkRJDk4I6oM6qaPxhdz4s149GJ5lhh4AWP+cehwUD381NNbA
bMVP4EB6hf1E+2YQz9GtgnvCxoj9hQ/ki/cJyRT1KDoyPOgBHpRIkGYRBkWsV4kYhva0N813Hs17
y3SQxtDdA/+GRBn0epRaaALy+KyQyZIIk4DA8EgreVBJgFzjfoRxDR8I6jOeyQpwJzly0311BPzg
trNh9JZ5fqeUIWn/r8EpLLENz36RMDdu7U3f6cIC3V4LwsaQ8gj77He7T8zB/bQX+hTkXdpTbmqk
uaw+qYUe19lvuF3fgDcCJXZxRDmHQ6SiCI/UII4O/g6I8drpzMNiwWQ5dEkSQhPEvSSbXhX7Fkvy
SQgXUy1sJukN2EQSweeS7tkWT76h8FWs7pgEbbjY+cq/2R1sEQttYDbuUAuwCAm/qeDnjCCHZ/Lr
1sGayGwKsPTcymaRgdm+YiHZ8F1V9sJX7QWo3pNgvv2r+tkrYw0F3Y1wir6g/GZPJ3RQ5mlsZAbw
F9ojmLLpPXLs5wA653mCwE0Vnt7UKRyaYrtr5O4yundvWSi8aO/gmO9jr3yBdBK6R4MoIHO3LS+g
DAbJ1+HhJp2Pf4k7QAVprGVk2KUjtoGuiP0/3valmEB6AAgCh1sPvzr1WsuTIpVgRqGv13aXNs3K
3/tXOHQPrfKsXQl0TKbqNFzYYDsw6faCOMQZ1wvZLg3Yuy4TZmPquwkEvg+HzfTrmPSU03a5E+ma
S48o9nJk7uYR1ipv2ixHHAKrSejbmcBJ+Cw22MUV2ZU1EdvxnEqWChnolWAbKlRLGs6fIXmxjwJV
Eqx0ubtp/2P6uLU630FDAapx/kmeL/eqyat0XVO9BEtjuQ3eLh9svG1TeCtqhXhduoftq80cBGJP
rm4nn1FgbhADkCELxxvqC5ALgSedq6hJCrlK//85sxM8fbikzlhRqpAQRw8/6u4sW2i5ZMuh0zWb
VICW7Jg8CBjJbIDE0EkR0cpjG40aqPG4LSlAZh23tugA+Ma7noyEHgz4FUC4RYvcBVLAcUsu8WKw
RgJ82/9IdNZ0PxPSHEEt8aGdD8hSxqPS4aCzJuEmYuhjitHnmcxOFeWXZ5lysUM3XS1MNW/4a2X7
OZ6qH1cxlhPjVY5g0rndw+xp2NeO/rIpkVSvXaGPAIk5MFH+nZNXVEyjG0YJxUa4qVj3+68ocJHV
TryEK3kXfg+TSd6MikkXoDbIhpoZP7afy5ssNv9dI+Djxviupc+zmUgBe9vM8XAoP1dmHHGdCDE3
xjAqBXF7CMyqFHxKO8M+D0dIy1G/uq9gS8BeuFwL00tAzgdMi65ebIjugFlOaVn9Ys/rSQtHDBtp
ZQ3oZLvJtynhhLIGPTZmbH+w3TcyaZysSa1ISZ1Bg0IOIPI13m/lIwPfJtm/cNP8pqGT8MX6PUmV
4ssqFqQIjf8rMzKDRazs/TdhYRDfuZkzDP0eT1pEL94MPMz857irc+4KLUztkyekREpAIP9/za8v
Pan2bZvmk3QvX6efJb5dmxCJmB+x8a/aczhPRr/GVFjT+jELozNGaA61yZq6mWpqypINUg4crW6d
FrYgE5vvmZRR9WGtRZMG/oK6nSnQmInyn80/MpmzKAYxTxZj3i6Bi52CqNbV2UXJJz0VUKDn6fc3
dYMpgL7tWZxjltYgiFlDDkbcvweptrQ2ECwxx6MXst4AHk3OcVNDAi8E2yrggBSwX2+DTKMs4dXs
XdD9dNzcykCOncoHJdR/5iFCv17JuLRpSSoBacpm1oiXgOzzYKJ8z1r9rLA0mzMjPK7eCtVy7lKJ
w01+hLr15UR3dofaaAgs96KgVNLIK8NfwwvYPi0XP2SMJE86W2pgczq2tVQfJ0w2sBzeAc6eeBiY
/0NnZZ/RIZlG3yV48LkUkynhpfvS48v22BH15k1G/3K00a/z5hfCAjj+RH4t87s+HZwdoGznnwR/
T/hGegybX2wBX+WL8yBmNpbBSGrGWtNc9qhW5OMRsEysCMp1HyDTh6yKgnZQUpe9q0Ef9FLcCdMa
W8MCkSYwXKM5cFenD7KmM/BMse2K6PujhYBpQaJi28I5A3WPmQqxKvtFSJYbfDjC4Tx7zdUF7v2w
VftBeKK2MK9qIakTnL9duOUbf/EBsQNI8VSN3mw5CbbsKEBtONnWWjSwphqEeF/90wVjEQWNgkdY
+ctCywflD6T8eQzbCNa5kifJM4LQtFvVNPeY7VsV2Kmq8uKovO6mFU0TSyFKLTGphqojesYsGwr3
aG7tEC8XsKiAOVY3wRZOdeCmWgoCk8DJAN6GxIxJ+bDcTEzPY5fDb+a46ZIS74q0AZSq6tP5l0BP
TDZw0tQnSoc+RvQT4q7KM491ZGByell9TCM1OshVF7u6Tv8IW+phv0O6qGaEAMBhGolCyrA4j1Sz
HNw/DGx3POcsy6Moib8PSmi2gu7e5/JGo1HSpMFPtkwOZxOEcURaOa0q//55yotdeOqpDW8nPEbp
vmaOB6trUheeqA1gJdDXoWq7HUnrFGgH9kbPOVOAEKXOQMcznbftgBeEw3tTAFGFOs9D3kv/SCUb
LLChBK1fGseU3snpIsC2g3PemjWvie8CkpCuXt/Wd6lH7jV5OrkrgqRcrYz1hXvTGndO/wvJ9MV+
Dp7wmKaeqCcIyeU8OPyNosjypiUPE/zcoH5+b5bzNyErrFDFyzDRCmpcIPkqsKMns1uR/kEBnBRY
RwJ0Vg39HlYVprqhoEkLnbZXRcpL0JSnmXXOODXC0U/ncp61AmMH4QT+MoIm76MDDyPUnLDsMU+v
3O8bKSTRb/O29jSJxMaF8DgmKdUw3gwT1vml2j00LAW/R5XsvnXdL8B9a/M5SI7uWv96kb5u9Mp8
klW3fAcDdI9Ez7kqmU5MvKtwfWShZL7sKqYXj5ZMN7QfwaHHMwfuhDEo1SVYwriqu3Xs+B2CDQvV
CgLAa6d66frCiqMEezc9/dZ3zQ7R0Suq9uyD8WAn/7/Q8NiY/GtWcZ9rc+qJKxOX41r26fn/eypQ
Fzo7BWvbvGT4tayvG0d3MBcL0+W/YhVF/r29jndtBFm5kj4HQqfKXmhLfGSCuZJbFSbBYJ32h91m
rNUVx1sIsML3hYvaGhAvc+FPQ1XN3PcNBu8nPB91xA65lKAi/AUqDuFIHMT32dS4EUKqXWduI9fO
0JYf/IRY51Se4jq/Dwu0a3CetbS5VBV9USHJH1D4Qt22k0kmTqRVJUxi6Umgqj4uJp/162uKyOvP
+9ZkQ8GqdQFjCp6q06Vr9YJPUxa3Lg7EX0Q6oo/SxV9QaiQjIbYPnxu5JJ0gfk++2z7UyuuxGXF9
FIrDmBxX6xdioOvygxi4xgu2sVQcI34brKRkFvs8EfNA7u1oTC1AnO2tczg7R4Sbc/6BLrc2eWcl
kc58VTY3LfIrD3GcFM6PNKj7Xy9TyOOxkPHMLG3/mgruohsc9xYvySZtd8x71JqAFcn6E9ZgVE1b
SZJEmR7oEGGIoAFjPUCUVWJx4wQOSoUc4sXgTtld+sW6FJ1puW0tWU6MLAD5Nro41WvpGk04IcVO
gRjdj09wXCVGRZV8yDUsH7pMek/bdXTKe0e15MKigh54Oobg8ke+3oPGARzJfhv+o092RmokK3B1
fbiVo9rHcs1/WEPhZL0ZjTVQ1W1aKLN6gMFYqb0VTH6pRzInxrJUAPtczBDS1lx5SfJ/cflnV2Pz
L/L7wzGiFYEkbfUjyOrGMwuz7sEh2T1SVFHDnnT0iMqqo/9G1BkedtVTaV6jvSg9Ba9o9pC7NmIq
cvd+KX4AP200YUiSCnthwCtU7XnPMHqGAMJlaeBLqrQPz4paz9LkDSaTet1rPThQQ1uuVLWIlNmO
pCAweypb1iNbsAaQMC9furynsu4AKxIU5kxITZTQ5Rcsl1rdqKgKlrYO8c1wm2MuPMHDBKTIhXvz
eqTAA2IK16pnlL0RF9nYQU5O5HdeKz9uhymyHGH8CjXGNRDwF981jpNKTIBwdbEik9i9Pz/C+Nrq
1FTeHBpg5c9tFQrHxpQ3aEAJZv7MCpsNADAjP0FYKeGmQfWAdvISMwGKyI4ZLpdd/dfu5gJXDyAs
9oykTnpiRfPPu4WXO6A2pnB4/UwgBtpfLilAkl7qG798ixMZEoNWG7NgNSHLZS+4Pg+eSlbk+yZV
HFmvcnHkgVgsHMRHHJ8LcrJmDspssO76z0FLawhwLAPtCzFMaxUyU0Fey3AuzWjRoNnKn5AyEMFI
SvLZIiP8+TW3fj/dKkyP6YE9ex4ckgSsLEhVs9iIt/iL6OAEnvamao7w4XYrtFmyGEtsgJ0iIhSS
eN74rvF5eSDvpglzSMWlJ3dZRQEcH85gAoQZrXp+xt7H0OZgkd4HR4Ni+TAnaMaV2vJ0PU3RBdsH
/UKi+ey0iIgv6AbaLYGa7c60MrKttUFRWi3uRhFCuCgHnVEzS5dBWNq2OxIamhfVsX/F8pGghIJv
AttGVT77LIHqDVAYwpmm9Aj2GHrLI2CLGPSG//mc4EZw7HMbXo0r+Fj/4lPZFQUsZyu8hs5AWG13
jf46CIizmYC71fLmPUUptukVQb4MKUbd4REjMjfzQj4g64PqhmeW3iQzLlNqx5sELDJHdUt1o3Jy
dlyiqImF81W3HlZj3WClGipjT8UwUQRVqu+xNBffjE0YsUGSn3DUrs1a3w5g36uZ20m3Aiqnj25b
AjLht6X5L8mCzFf5wZw7oy6HH5JkZzzYJWn04CNAsQjrDhUbZRH9o7vngcmb3ywamCc6i0a1+9so
6g+n32HsqX6iX8NrtWXx4nbEkYkFL5NRyMukjlaGD6HetybP0eTz2my5yyO1mXjYUV/ILhgBNBGu
F9Dxn63khfFRDb1TkYT5NN/FDsx69iJnrEJRtyPQZY+ZOpnZjC1F+9GlMpC2h62LaDncDJtr2PCF
hPo48+uGtsVjPgc8ODnRvym+Bc6bxft0ea8UfTZ+YBHHKYuS3+pBwNqhJkJr1c1G0OAG/6vEwPGf
xWKbNZVsqFo2WXU1Iyy8dQ74xIL5ANTnhLC+/Aqmott0ntZQTOxiIe8yOpicQaPosFDoVsXPG9nP
3BWXqld/zRxdK2ri42XiyvX/GPtyKQOVC2SHA549RE2wkzEp/zGupNfWft+vuaeu2mc3JPDypSfp
ucxRRXuSCdAB08s6gTa0s+jb6mNvaqg/KDhRiW8Vx37yk+2zzicvaitgzaJmEKDpwFscmzVe2+eN
iNO8pQcWckK+Dr0ZFWK+NMOPDH5J4cs8hwHAx2Uo+/Zd1rpSzxZxk1fx4pTuMk+K7L4x4xpE0jus
dTPJes6QDrFUYJPL9clDD5nnXPCnmtuScmoljguNspep0YPF9XZptP98YX0joX566wtfJ2oJtwSz
JOn5XinkcJqbimJuqKalrCDVPBdNPcwur3CqzFx669st5uPdN7ly7LXpEbEcTR6g4QAtzupTOL2u
GlCPuD5jYQqFOfTAGjzopRfJAoBUi4ogTCDDRJM7y/yaAGmfqxuuXMKruItlI9hILDpQh+fp7kLf
wu/6frQPkXdsHwaMPJPynMMhDQrHYhYxoAO4Kl+BuULUXrClUVycLqCdd2hRtNJ1j9Ac/zmXA0R3
510RGVVBzRqMU/Gw0P9VXBcE+eQvLJRdoP/RmvdpXkLoEA4eL9sg+IEjCWgxrYn0LuY1g1OOUH5C
e/7ul/yY39Ih+44y4ZiR4V50NXpzLKrVXbqyyxNIpcHtT2CDaw0XtShT4FU/gCOMux41zDG28l/c
6fQX9V6V2RzI3fhhwor1kAA4lOn2i3FzuynDj8IjHoQyZ7jj68PIt8pqQUxTp8VPK0QnOjpLeKWU
c9buWe+AVVXJMerifEw0G3Hn/xSHm9CYkF/YU5PQVvR2x6rB5o2tGjN7JYFmuP/K0GZw+xjWGsnc
rBxhQmJ8P2ZEjAAB30YgRZYMLsWggZBX8IXCsNSeNRSsMay1SIucETN+u/VULP5lT25mIT1/OA/n
tt1xB6y9l07mBgc0sdHz8bVodlc84pUL/RPzpE3Ef+LCtpifiJC83uLwBIXp6SH5vcvRxHeeVUeu
5iVE0YFSplvTi4GKCUovUrEiAMakZ0Jjb+JOZKsOU2dyvug6r/L/Zg6QMjlVjqaLjTbpteY4ve/r
yQshieWVqn74ECC1uC1MPlEnrTQqYJ0/0oEyCnyeYAPJHwq4ldGlbduU1a70oQfc3WVROBD9muhe
iRuACIJIv1eaR2L3OOAbZWIJpQW9zncvNNEfONbspU3D0Lbq041X5IuJZn0wmROdxerAUYNjBkZP
FXzL1FFLkN8kVmF79BVngNxGpZD9x9pLE1h4ede7oUmS1ORdxz2WHKjlIhrW1MIpk3cShUjiZcGk
QStkiNDFuCmONGcH9f5tp35h3fRqtCdXWBh0hwR48ZiRAsdWNg9ULOvjr2jvAop9o/JRbKwpl6Ta
5A6/SBlRluYGuxiZ0qjnukm1GlJNqst22ci0GDWjSQXKV9FA3r9Ec8qeznepLINuiinzlm7GwbiO
z8idGIk6gpMD+iJplcvbp4sK3GTMOT4mwN1FiyR4syX5S+XD0+Qu+/gsv43jsPQ/rES/qWlYixI8
Q1CJnfMtWuH2VrN4165/WsYAJmXA5gAJgEpkLijQm5U+zEfaFH0Ahz+wahk8WB02cFB2qhL5GVXO
z/ImCZYgm2eSIYi7r+UFNck7R+rwYnXlEJlitpRWxMnISEXlniiWx+CNRkgrVhrovlOciWlCZpgV
UwtdohK3vB1fjUDKfMt6N6GFwMUT7Lv+jPTp0ZMhDHqR+sUpPRUHd92OuhFOmQbF/yNHWbHUY4Xa
ySHKsVXI5D6mTmPiZotIwnTxvKQrK429OJu982cbZ6iUaDHPqbLEb7BY/27z7xGVPqSRB7fjNqVi
VhPJaWtV8w9H/dmmubdckY135djshrhGPcx6S9D28sD4dGuBvYTDPE0NllEyC4uA/mkADR11GjUg
8BIKoOsoBubgOyctPSZQCgUIcFA1aBRPWwFLwa93OJqi9aPeUqI7c4o58G8+kozdRIi+DK4vKDRE
my6jvPGc5EQBX3um44BcmuTvshxpIkCAm7vzUommTBcCe5CoMU8GdLIx/N02vg36Y9UI8HoSTo3E
2uIWl/+kAvuH5eXb4Cz/mPLGyHL31rG6/gw+0MWYm5PYkYXzmswAO6GEHk/SezJk+948R1vVrqXD
7KChU60YbCy21AcYgZTKhrvJRM92WGzqZvim7htQ/lZyoYwaO+UGBXsORUb3FPJGpcHVlPKmRsMX
xjV+8CgpfSgt17HOKs7YbSHoB5HQn1ct0vHOsqQamoAnpYkUnl0QzS+S9NCYuWLGOIMSlrHYZaVH
mjR6DCofhFx89FEiW/reZc6yiuGvTBk/cP5ipkcrp5jqfj5kp8/cEzROk8aZBP1IIX9W+/saOMB0
5E1h0NpJcZ4ukDl1Xcga3sVCOvnCY9pksKGyUFzckiaodYHm0jhUJ610OQ3OWoDrRihJMn+nWO7b
iuKvVPBZcpFUwS6plY+iVnSqXNzd7RF4Gt+n8hA0MLONbRmLGSCxSykIGDO9jBuP6HE6U7a/1V1X
CDch7ttBAAAHk0UScNFtR5hwyMBWOR5iEDkLgjUn68Rsuks7LPfshebufIFZrJ8l1LKNI49Un48R
xzRIXqBdugNBJ550AKzvqCCYX9fkCYlHNBElYsuzhxz9d+3TmUrYIyN6mVg6veFjA6L+PisMVxtK
I+N73yP2nYpkF8+M1E/sk2u0aLUrE0wikMujxKeAmgkmsEBLG4J+nQYOa+LFl4jndFFNL+MbwF7w
Sxwu3MK/jpkSErv7iEk55gZUH1kQ50xLr1/yNdlP09iBfI0FwBp7LnuPcsWCqQpd2dVMlCjdYonc
DO//A8jFA9E7y/QQOrahHTd9h3oNivPuRtoYzAUYnCVTF2gZsRXCEKCqI387aXo0ykyrERejZsj3
alBG8c7cOV/r9DrS/K+ewHLMD33sx/OgOKoyBmCs1QP1PSvXz1qJxjX/oEzzzEl/BhJjnA70N+Xi
pTfH5HJGHM4fXtg/1f8mGhW027Tg9rGdI0WU3PmGpWam58Thrawsfg4XVNqaOfiE0blyFEXMV3Zk
Th/Y9uIWTakKGNPliASwCJPzPOTVPzOcLfdBNc1ltFPU69vOzL+/bXgHhuqV2jOLyk49t3h7yQeo
9tE4h/n5g3fyVqxgH87QE1+/544QUhUbibUKHyA0fzAvt8D7uD15rQfabCe2yCsCSLB9n64PuW1+
OYHzX/3ANga8F4lbpmgRCo+AXK7WSZqQA6Ks2n/5fjInGBQTDR5NasGW9MmGJ7bN8XtfgPVoIdN7
PTR0+ov/vz8fhrC1ejCDHeBcc0EbEyJjtPVsoWvb/EFZDCTL3pqcX43TJv7G+K/Qll+Wa1KaxVf3
O4Lch9b+gnnDUUe88Opf/R2OXlvuX1dfB1pae4YxRD2zaxRbwDjc0HYEM8J+QbvbdKEWEBAysr+Z
SNjdP4uHecx0kZmAlYHojM/FZhQM0W6souEpEkjSKwPctrsRyz86GAMa9ZPovYHouWxIZ7w8QUWz
TJ49FImm6Tx6VgtdImimHg1C5HVifrBodLpmHAh6NJu9nXAPACFMlsV4A93V66SArTLMqJtbv0WG
F5UQ/6i2kE6tg8T22yF80vRR24J3lsJTRXuQAg/WZUtDcfoxYPGJ0aRgJDo3Z7wPenx4KFnpCblk
csFI3MLNBZY09jOkDjtBOawUEb2erX1gjsylvQ6/GH3MpG9fUWWU/jxVVEch8tEKqGXonzQa8+ug
nLMSLX3iHYiyyp+fO0UoRwORCWKWcYJYGS3eNE8fUzNZ8aAqApFhrBqwCdIyATWzysSXuDimnUeC
j7AOsC0VCvX9RAg1CO/3L3PNCCljEpkrkPQjxdKLzKbv5NK+2e6h/ekmApstLarBuDboXA94NFSX
mzlo05hskhfEOG6JnAwDUEALL1Vc/AlDw43lQ1pRE+xCtBJDWAlX1ruWtN9ofHcT4xByZQroDMdV
/YM5pLxddxzD2iZJRJVBrERRIBDk33CVuc+pE7tyWB9aLkuNuYGDns/u5JCfGxY298dkQcnR0wyT
svCEuBEHOyfzkBAZcW+MAthLcgAz/LBA0OjjlOmGD19xXJoBA9oZep3NQUBVt3y1hxZM0/6RN69q
eU3OJCcfXY2pxo6S7ja9SUVYxt087epMFpRiK5Phs0oib8i1WmnXVqnq2h+nyX9eKqm7hc+rz8vY
YEnKeBqMrjGDX2QUTnGuPH2pURcFoa06SGIysgG/um46aIwm65qRW2lF2V5po8MjrRdJcPaod7Df
bQvjFj4KuK86My0SB9q5hNwGFGAqE+csHBF2hAjViYNS2IoIt3AjDIhTWLEgKU+LwgX9HzekL9+K
KaXAff/JFtTgdUfIzv311DKaQKdub0nTVMP2XW7YzRdsbXqD7kXWoDdBRUE6hYfqBSHIEpalY6i0
fi6OVQrntBNRpP75jifWPCspAmMmkrJO4Llbu2J1POQRv/QGVqsoXR27dX1+zv8Ef4SQytYVdRTG
4AM/sdMzLC44wQDBJhaK9nhAxrFccc+U33LuEArYwvR5B8JcvfKeoMIR224PRPurW53dLxmq0Fqp
g3gz4L3AJyfQLylzhauuVEPG3LZmh4yZZf5+b+Ld6JhoH39VrglEMVREb3jO4a8XCnBuqFu3yZLE
LKpY1d4XJFTojBVpaCIY19Z30QUVP9fW9qfDwwFkLeLmBp1MJtEatdsdAoKsWoJmSq5RRCBvTPt3
fwYhZmoZ5IL1ZgK9GbOmQzmamfetU23SXwxITvHJKpCUhNM7LgsnfU4taF0Br9MsvIaQ/ydqu4w+
FrE9tSj8VfDkHSB9lK0qz2/YeT7EEaYVltL5Ed0s3RckxOpAjRq1IOOmueHat13VRzrUc3RDjQIR
v0rpMBAoLkB6PR+SU1Ijdc0bFRAcQkiKZ1h0gz/95Ku0lDA2V464SqtK4in16QnDxB1Lz87K79Eb
Ss5LpYIBEK/Y+TNKo28q3o6bNPahAlSvTgyEd5zbbkJrY3CAoJLv+aVFVN6EVPjAw7Kv0qguDKyj
cGJzfNByc0Gx2786leFgCYTOTOar8I7E46iuX4Zk5vsD3agwD9uA2KgUba9isO8oxNadMMKwKcZE
cLCe4whJdvKVcS7ZN1IbbgFKF4gaGxpbWFlvo1OXilvyjGrgXi0sUiYSQWnSE/FSrUWt2Ha0NbXD
G1QUEli9q+QDPf/EJl5wxVF5jOm38aI0JB3tnQJVHq9knomLjD8nhM7NadvydUOAvFmks6jhlutC
wDybQ2mdL3IB8ie5tv9UIlbKazchXfyalWP0G9Dx2s5+lEQISEH+iSiZdlJM+RVzoKW6fRvnFubP
+Xkhz2L7lTb4v9s/ZizltCk12ozWiBnVSwTW69N/rSlSinpuvCf+PJ8VYcdAUf2Jn9qx5WQfj35j
KmFHpWRF4VNe3kRsws61Z2OCuQM2uJbucX1j3bmeArpt8GIZHIgAJR0ntyikzkuEIVrI6eGMcGvQ
53OvF8sxok+ZX6xrC8O1vf1cYG3MA27/jHrRex4+Mp7sSNkp1QMlYf4AH1TeSLxiNeMxzUOlxMu2
emKzgOszERFN59egERjt6yZWdlxMIjZ95PCy5Pc1sq1sjyctV263tU132mZbNbaRDOSai/CTuoM0
lsNvx+FvluFORqD6PKjlWA88Yc0711iZf2gphc27NoYHYSXlqp/2EiEhCYTJzP0z20OOAaGKl882
mYdRf0cTNR9wBNDFSJouNN2/Dw1mN+uf0joNCfI9sTEvU91MeoXSLDEl4Zd8IlRuXux/sefE8CHu
y+Gg4PXcWRGzAGnjIkTsaMt+gHMtc9g/QMyFwsFWkbsXHKomWXYwS+De0rxF4KMTiobqZIxGELWk
J9Y5BfZrVdZmHCp6FAlmfFvHNM3+me91kngoD1Nx9oQ9QTTr55f+zsPX8MKsE8Q/uX4v/Y/EAHAJ
0zqyt1PClL9VTA9OUcMz8Y2hevPIKhdlgwtXx4tvzddtVaCka9dr00JCx7ABYZFeyeAodGZE7jc/
ihPTnfz5sNfkNA1+wwRIL3z61SkfPWN0F31rjmOw9WudJqDULbQjs7jGa5xSm6y/zbmmkZEhwdr/
HExRq0Xgf/jQ7ESZtSWmS7saIGsDY+bDLJFzoOnXqFwFCua0nmMoOtDi46rZ0cKwRzEvvbsJhpAP
PVuGzQ5yuuweMT1JXGu+lwl0rylcDEQzy9Une6pZQ69mGefjAblR24ih1tT8b/o2jPwZgKWsJhFE
CiaETinM6FpsClGDvSa0N6rmq+j9kJUtvNzxhy+AoznY6HDu1XA/KlWQ84LEi5+v6rslSUK1SAEk
XWBWDg2jqrcJHiMtMvG+7r03jj5kn1/6KcOq15ekqIUlhwQq8uDfUnDMMf67FiCNpbPZ2RC/va+f
N38poGZ3p/8PZh14DT2DCWTqwueE5lw3x6+/6hSy2zZ+fxrCO5/g9uMusOIt1z0pxwy4PGZvpvTB
OhL9OW7hJ2QAG+1JK/3ZgzN6ToltBpJolc6R65HTzMo+HgEdsrNnxwa3xex6+hcQKE9LgcaBWM8+
NPp3o3lEPwOs8G/Juvuv12K9YEjltIxoHYg5ffo0J8cvnB20RXuDJGuH6BplneQHNgFkTSL2epRM
KSy8GRZpNIhzLZ+fs+od5L/vU82DePToCbEu3iEnGCaMoHPiNdD6xE81pIhHo0knAK3DzbxD4AnY
Go+IHHfUfLDWz2XLjGhxxULbPDioSeMeVUnurLAZ/15SIA4Xtmi1uvqQu5fe46MF03/a4PnRyysS
hZHkUhPucRYMPEd8IJrNTZvgNLEr7F3IiMgiT0TP6eSbmFjxZii6uwt+cv3reMeTjbRcPdPctHK6
s9P7zlzm/37a2nKfgLEihzyKE0uPhI65mhH1tJGXJZa47sfGDFURXpjOgBWboG8FSiKeWTfk1oPJ
2xnB3RnVUrg24gXf2Vf2dTXXwV3dkhRGbr4XxttVjBvqRbQcxNGzmBNSKz0X19mUAeWunQWkExfE
Pxnb+STC7nbS5e6tr25vBInS8ilfj/JiljvAfSF88HLn0WO4Z91nOD40af4L9lXeFMBCG6shgraK
7eqcWhFxQOwkuIU9nlsCCI6AIzUp7CDj7DyJaCzB039gHhlnm1hvok+hWUsqcMOCd9Ge8YxOSEbi
Bhf+VQOgmgSXNZP+X4EmihGJu0dBR339xb7iGZf2cnDI1QUa8XdOpjwYQLa0uzYCZ5Fo41cNNCJ5
Aif7ReeeanpHRvqFy25DphRYkCX6D7bjiaBrKYVX09Dae7mISCuGyqNCEZDDnH7i4wfA0gliWenL
T44nRcRbYbui8Au4YfscaHsdWrjZAI/FcTQ4iW6/E7yLdjQmoD5WTgnjInZfTh4qZL8bXPL6CUTR
oGNftG5NYqTuD3RfAemZtx6ZJbf7nh7xJ7BexehcsuUdFf9cglILdnafbW/cz2adXIq6jqDhqbHf
FMFQWxSYxv+xWZpxic8V+TiVYTULzFqfJrfXTUEPx1JfXQrrmqKflnCqOxt4vqLfXZFDSX9+hY5j
1WUeB9cPlBP4wVOVAGupA5KyJ5aRqbOGeJhzbWgk1kJlzVGnbrtrehWLfm+BMIilNKwfgUzAsBde
QJrHI4ubVM0SQOHZllPVaoa0+PkWC8gfzpAOA5X8fddQKK1oYzpn1Jt55hSKpyNJsI/sa2KD7CPx
KwBusHHALVXKfLmUu0J6rin8z/cFUbe7xFciYVG7G3IsFsWhbphapVr0cAnPn3BWiD9cxuyluUrh
z35FdBF82m86EfqgODWJtKi9nuNPzupvrpQVy1McKXnHrEs/Wd3UlP8U06ej0Z6WeTF2EjNYfxQs
TZ6EPZ+e1X4vQqFcFYcLc9Yxqa8XK3Xagt6y/qCADIzUkMEZAxdExjxzPBrr58QEkkBdnsObM6hj
Bm+J3CP+Cgd1Zecjvn+mtLesG/e32OXxbqMJFCuqg/OjnCO+6Cg4Xu4vhedjaixoRMM5O8cxRZKr
8UT0L9nce4QUO/vraGYGIcNA1EZW/pChhwYv3C/Nf3WxNO05SSIw/DJFrJmkNTRLdDHdI4Q00Coa
yRSQURaUKIohMarH6abQBy/xYbRqmFQ/4a3sF+yj9aZU7XLmNltvJpp5QxHt3kc8t25PRF2oEw1b
g64N4RnjmydNJRPS5ZBEe9VhlJFFdIV58qWH2JEhnP84WZ46+4NT9wQ6GrzhZwCuzKljZhMsOOSg
ZumLKCSNkUQdzWesQxg7dfv4PbmGedusPnNssSsvtNPTecJfhigpCFeya8x8OaLgZVO53KkksWQy
L4hpGd4oY3voK75bd/RIv02J6u3xaRA/bsppoS13/n22ZpmrFS10/Ru1yh5cLOJdXqrqSL6IjiQM
g0SQxQXmaAXm6QuesysrNmPuehzIzQ/nPgX85kdp6qyNzaLbDy+qkBoPLgu4ig6rikDtjHcI6M3O
Uyvm6qcwxbPlZrwEXBiYdtBCQO4XjOsmT8tmklEPLLe3Xt3tI1dpZVH8ecarHkTLlQ/rR8cCnL0D
6Z0bf8ulIAwd188OS7xuu4degl5dKe5C011mVNRyJbD4VkJo/j1LFEXnD24mIszX5vFUkcLIrrgh
s6hHomVZxpgnicwKgHwCHkWR2UPBfxBbNqjQtTWJ4xkRabI06Y2n0dh087OZoGHOcazrGPVK5unq
PYESzyhm9rO03VGSyf3XrXDJVReQVpcQW8TCAo1/gYzoNZ/8Vnfjx4m0pNOW7no1Y8NbuVkCm0Br
cOnfMmRj4loVZ5lvNqSUfGyAX4K7/gvehAU69a4e5MGFpt2Wp3d8SIRV5gTW3MD8Jy1CvyAs8pOA
SM0nEXmeJx5vAE/3JeLztamnPSg3H3k3ZJg9Uyg2C5Lr3RdmRsJx9lZntPC0F7NzSQ20fYL1CUPc
aUu2tuZmfRwM/cepMiPyw2urKVo+SD3O7VTwRkpbKuu0R6oq7eja0HiO/M1YV1mL+rX9tZCfRwX6
ej1m4gFAgPjXMNj3aK6I5N0nKPejxtWiO3uJf6FwynTyMmrdlHLueO/TKkJY6XfTr0A2qoMRxOYX
lNLjxU6LeNEG0epfINOWzF0IF3Iez0qvzgjnS95b4s2j9hoz5LZxmrsKJb2BN0/OYXD/LV56Z1uU
U37Y3M0WX6ThvYRAWDV49XqdHLiOyQekGq0pSLPSpVlGlRsYBDWWXzES5gh5Pk1G+1aS4OqPlUrk
F24uyZNUgEeJZI2TaJbqf6Smkf1y4k/XCxy0WyTMKVhH3CtnExc+1pcARQd5l9ZA897IOQdgD2DY
uvOEhyY0hkBTQPvlqy9CGpFZGHLzXRZ+SfWd0nAPEKKdTGVHxm0dsOLMqpXLxVPriJFPw4R5XUy+
fHtl2p7aDD4Btyt+sBi89en5r88Xqb/j9vmeSkh1BHogOlvl0FSeaF8lB8YSrdBQqBKky8xi6+Oi
J/CR7Y9Mk6AItbCsPVK/ZOZcMdGz6MQHzNWfq6fx0n/JBf1yLa2NocqDFhreHfT1Q/UvK6vvJoOz
ub0KG/a4PIgJw09Qkrl/h1o/7DfxQlqskZukphRRwTOexsUjkJZp2oz/CAONxRY6ozSoVlSigITO
Gf4XnTSPBw4RRtMD03J85ciJy/Y7bFaRv8DsVE9/qMbzUxfyT98fytG4XDc43n029DvNXUk38/yA
n3dS0f3so/mwvBsR1zwDys26hdbN2gd+T5V5jTQP5+d3Kmzb1xza56RJt4egOpvQdAQqe1VEzXN2
jYUGubInc0sM4hFScMkcFQopuib2NMgOiiz4pYWfcVYheblHq/NIpM2GFrXn007O7KAjHiSYISG2
0xQUsMjp3NMeUfXpnSNLi/fnvpwCEnKgly6tWnAoKYYsVzqw4eG3SRIV6uwSWYrURuVGjqcusxeJ
JNR9ktE6/FIY+mohAi2meLPbWEvbBT6H2SOHoQveGVQ1knEkPprC/3BAxVJ/jpJGwRzoXokRKUjV
ApsCrrOiUlWwfTpIGj48lTihcYhWAo/TlR6VlEKjWtU8GkI/vL99AbAddTedIlWBNOih7cmz9dBs
Ypb7jId0geOqWX3FNQDwjEZxyQazEg2apIyj9IJMwW4jLplWPGWK7C1iwbfqXRwcLiWX1MG9WVhw
hYjwFTgnFJxQaYezaCeL0hU1dj1YaeF07ac83jZrHvWmHg3CQ3dX8o8rLvNEqvw2hvCC9wHbyB4j
vk1P4mmR+exhVAfo4WwfFoBAoouUjIMr5JHaTZUhY0ryAtIN/0c3Tqor6e8AqMpA+asYqLsurBMr
4ceplhl5F9RvEJF27gSmRSBqZH9ltJ1Ylnug9v90W/aZyalpKrDnSvewKbst2v1YQNp/pxe/hyug
v+BgO7CLkxWHjOngF/qoQPYgAF2cNBqUrX7A+i9Jb2e3+B8GNg5n2kmDuSGKaTiR8ehNbDGYq/hY
eZqY+wvvJBwK8s47WuLvGcAbYqvKa2ROu3dgTkAAzOs3O5CP1NyWuYZNt+AFt7gAhLea/Hg+GcWz
xAumWtPTO2Cl0+TDuioY0A6nqNK2/0A6iP0ma58kX41Ijp96kMj8ZSlBPvEAi0FzDH1zbc5KF5Ap
wJiMov2i64CC73qwFTBOHi3wueBL/LCaW/wBV7VYVpnGnJhvj7AH25cWdSA+mP1X3ymRUU/qKIq6
eoenmkkVPKniKmaW3Tz6iPBhg/GdapYtvuEB60OyEa5oYzwvKCaeW/ORw1DfwCd62SELG5p0qZ2A
5urIkNJpGyeuHV1uy06oRX3SIhDzShtDOxIKMJ8YbXRzKbnJ2CSPvyAvwWTtCPfsQyuihRVQFsrn
9riqWlKD9LMVh4zRvBjPL1jq+RxTD2QxpMMzyMTlsmO3GSefxbjGzAeFiGYVaIE92WnhoCHGrhbw
T4XOymT/InkYDPaO7G06I56W3dTS8tXjGMit6lrsxDxxoE6CCw1eqaAZ5BiGyx/J5yreRd5e9GJD
HHbVF4VY83Vmwj1ipF1CKNFdSQ4jYGEvY4Zz34++0jVCTlGANBdxwlLks9/C9KGwMWsjM740VdlN
iuqfWceC83phNLQM/kd6F864agFu2yRl/1JEA5hRO/Ky+856cjlMOSB7jU/9R2ZxseNGVSgCJ2Mj
p0zIHGZsnCDx4tpL8BUGTJvBvMxKU7GS12fBE6jPEVAXAmxlE3Bbd9p/uiakqpB0g7+//gshtZv0
eNvi+gLB10FTre8kQDSn6gHzotQqLQDMlLSel7DG8HFcOaEm6JE5jx0UhpqcR9lMMZK1tzm0zf4M
zKrF7Vr5FOWYHNMjbFauTi5UInaQXViFpp+MAvuyR2eKuKm2/nTPNmZKJK/WL+p3+wsXnB7k1e+s
UxRW/XIEJkzFMEIi75mJhPdCHzgP2IRRx+rCh2ehsLnVUOVcEuFnzL2JXC4I9FdH1T7Za0P7EZ3K
2RjLaTNamXfTaJgFofZ/1Ea4NLyZF8kAiC2eZsgkCP5aeZIjjBb/viDAPsAc1MoVdzx0w/I5n4ON
InsizMt21b60tRuOA7DQBfsPTZuJRO+DnYEI3QxUbYCzhfqFVmDhEMBHfrsZOFyNMk4JJu/Uh8wj
bHcdqwAp3h6K7vfDJWQSsKJyybY8NWtaxOngj9Bz1OlajxvLxLtnhyA3myjOicxM3l83CCfaPIdm
8pePH5z2okF41lNgwOTpWhq70Bvev07FjGjAmJKaUvYCz4/bGWbAskpIc+sE3CKEAn19ZOSXQJXw
ERSwUdyybjk21uKLFi+wu+CCzBEihGdtIENTs3LzyfaXJt53nw1MsYNmiBnis5gGYom9ZgV7fT6D
IEWNMigtMn3NNOlvzLLj+4UUfYdJFissk5Ggn6fHwowmI4HcGZSuPbEwFX5sDJuPDhydha+8eSs9
vXzO+kexjQcn1z2ATtDmc18c6PxAHp8LFw9C0FDNqxEHtJ8UdFwjzC1J4ry8rDv+IwXcamUd+rLW
raygAikB9RkkW3I04gxVPouScTmjFtkmLZ3htNtsVTW96c3GWM7kVJGxa8pxj+9ZDEU3SpCWueSl
kWfLiuNFkUIHBChhVLKaO+K/Q3Vk8mMPCLDczx0viCQxdAawYLFfMSBpQ7jeZ2QgviAvs8C523qJ
otjOwpv+2PfbN0Yz4HAkzyfbGjCq7cHkzqgTXZCbTINUSL7jUvZ/T7c9wfVua4wKqyX3+lNUwFB+
lRUcJhiAqpi4ehZjzw1uDcKFWh23DHKMqzYK7Sl4p3I6NJ7UHQmqLHUwPAFDGcwNLT/jQvHGrf45
9sPSsMwMsxh8gA6icGorlZOCZSvVUbyo1otqECbqoOp74ILMNSsWpXclcXssi+gU8EAIE4aLH1BU
QGQLcWfzF+pdqrjN+pLFlqGmkje4zQFYohBprLnLdgym4GT+5QuZa8eAqsBvJ9rgwZuTHqWR9IiD
pd3ZoTrAnhKnG7/TZXzYAyVn2/FEHXT0p4804mRpaXL1B6iAF8E4njlL6JmINkMNYnF5eraUu9bm
bi2kjCTyBOVKjLWcOZl34rCoR917eVzkr1KLihITgYRDaZhVa8B1Lu+pWyM5x8ibstC6QQ8zT/F+
uEayaXQ32cU2xPvkxv0q2kKX1P0l6bZpikLRTpZClDIFwfFvQfZgQMxKxlnIqpmVB/Bp9P0GW+3D
JV4ob1Bykgs8wqO5Q3moEJC4GcB+mPr/mmhwVAYEr5u4Nn+Cf0PipemTYmCQ0k42fH39UIxRvI2w
CsorLDgTA+GsVxtU0d7dpEAwrPzaJ/epATL3/rqUGnFT5L4WLT+RdeoSpcFJSIOLJLP2e1PTVsta
gwSX7/Wh3b58gpoIXGlwAyEsGOj02DHcu4dQX6DIxycjDdLMINjWpALAQWNCSjTVxY0zgNqvhIh2
ucX1G2MUF1oyN38Zb9RPsedS+JXsOwMpXUfL3dKn6yzAVjmQZ00iL/Gzm3Oq78cGGX3hGCOxTpHO
TkUioymWe037DzyDzYplaLEh51+IOGJqiWQe6nUb/tF1DyeHG+2C5zjC/pRutq16aGhpnAQ4HrBs
NfvHrVTtpiipfx/3tKQEktIbM3AfCmZCjt0pzzugLxXwl3y/RgVpySjUk8CRBcFSjZCCM92F8kOm
IxWt2G34fYzGvCG9eLOvsgr/IMCik8X9RbIexsid6hCqZElC71TwlN1QOxGcyTTdfv5MvexL/brP
9uMrCCnvXUHkz7ZemYpSjiTWO+XlzG/Qu2sIgmiYxTghfb+bUPtzuM4I3VD7K/b9oCK48dUiHMZy
+EHvKcqA4gwgLyDwUHbqRAZmmjoLi9nYkdTBIb58SF2ozcZD4RhLNbZwoIxPRM9wZZgSbrRlp875
xKpVbALJ59KiWbruvPmd3bjxpMxkSBORL9/H9bpMxZhdLdIU/wWLED9R0/HU+Tyg24+vRhjvZuHN
hgbZmCUscQxANW3whkE9XgD964xzh52QA4uTSj39MrZpDk2q2SupJKoejcp+RRfuxQf2rV5FP5uk
N1mV/uIQtr8OFC8F8xqFgU5z67i4BGXpZZLlwJcR5tE2/DPao8sszgAAc801s70grjUxEKJfFy8A
0G8RidB8Em4o+jiXYzipRu4HLh/Fm1WlmcJ7DxTkRQW9rp69qnt/7dCy9nr4d79hDF/qwaXCBUPe
yLXZ8VUUBYFJASZTpMBiZZwJc0e+ok8R0qnaQk2+nGAw/mgck8NngBgsD70D4Za07KZTfjewe5f2
XmrSaAwRoeAgSS0U/2H7bxW0X51M6t58scvKKttdmQOPZcPHGOlE9FR1tRMfvTg6W8sDVIBhUGH7
c38Bbwjs87rBoXEEi0TctQSzbMc2TV9TaSalVU3TMgjLgho/ytCwR08CZGuFKH7wXkut2IYEsdHr
/GNUaZVGmNDAnd0WkSiEUyjYsTbK0YLFaMLpYt7hDT6iRQ83LLV20+rzWZntcFTpM7lrBkwaiqq0
xn0mYTpSICYgcqk2XAUmYDuG1EKVijuK7Uyx00ufChB8B01fCaKkV63FJMuWV2Q2EShVQDfoiAVY
FwmvAMqaSoO/jH3r+meblhov1ZHLAFAnSITVHCnZoitJX7cFdLa1WQ5iocugUnE/4liPIi7haKLT
2bwqHQ33CWHdxsCeSxsipGEeY1JUDP+AfJ5ggDoUyO5N/kUlOtX2ebe2pkPPHqe5rhhcSTiCOlCx
GjYUjmZUAkkz06PNHB1fXjfgT8Mv4UwhFS8rdMLnwpo/hEgcav1n6Ac7Q5qbrOM3f3/ZZFSrpVtE
XdzljuvTrAHqXGOs8VBLYwGctLVs07/+QgQtrP84n7tL7WGcjOnPfKzoEmW7kknBkHpc3wYXrbLf
BS6njI+8AGM0t0dAPL8/HdozQx0SxTVFiF92zmNYb1H59RXQaUa2VGzy320fUzSXcBAHPvbL54kg
7I64gwQYOi71n3J23HV18F4o8rQOkuHCPjS30UyYhYxQZMl8tCKT5SOG+2NzwvdsdqFiv2jKx480
xnuuRyGZYsoTPV69C/UrYOzGtUnjhNCbZHmO5uqVxl4HHuLWay+eXrtqnK40Ts13W/bqWiJgWY3R
h398EhOuMk5bNV8/XP84N7MHke22RnvR6mJ0LIZE1hU9Udf61aZ/ik5wqMVr0LKilRMebd7di7HW
1O4HPtbn8l/fGD/6U2EYCCCHVYCZNCyovywjS4+WN4I4LBWncNA+yo9+/SIE//M3RnJZCvEJsWBN
I+6bZlF7iWYxN1S0pOGL9X0cqCMEUOuUBK5LVMzejK9CX8OAa8FLqciRbG+ku0whLfyntszOVMJR
QlW0rMTl1cdO/LXHaJiQGnB8b8UcRpRAfIwRc9kzoo3DmlBF8Kz939yHup4D0f8TMyA2RkCcq4a9
zQQwhST/ly3CVApzdz9xXg1IF9Lec4eskGt8s6kyvEbJlUryZyphnb/GeRnNsxWRYd0Xgv6TwdRS
iWKgaOipc2yN5xReBzHveJtnyAS0vb8PNx9pEpoVohYELpk1KwyL5YCbMoxeBE2Wk9vRVrxZ9sOl
bqvhy44fvGRtrb9FLlYCDpvnShTfSVBzvoDassJuQBrT8tSN2SkQ32TxjvFWKwL0xDf3i60a60qN
6eLr02SUfv4Fajt6TNRc7G03b823U5iOROEsD7zWL11dIQrjbGmWisoCLNQcWzaCGhOFX2D6jxqR
uquW+uRVjxdWzx7wPhjVZISp71DUa6Z9oCrghE33iAYotSINNytqAH5NdeEnRqLoRpJsdMFXMDLy
mZ2t5aI/Ugep36ZHmW1r2G21oSDvNpUJL62Y8m1IdMqYj1efeZ8J8JAyDfPiwDYv8aHnOukPEitl
jnZxHuH4W3yw3v/HfxWytiqXi9zDUp2fRH4WP3dwQjNxMXmwI0kJ4PbU2jggO3kelLs010QKioUu
2sBytzCCYAFffpO51Hbcm7qG38KUh1k74mwHIJCIuUFMUZvlVrq9OL8nADhpo/RCoMUrzAj1Wjls
HClAFzAWQHXi3O9Ty8o1dgazO9a85Ri/QhfaDEguma5DZ1JhG5hu6mQLhUW44xKW5f+b+hQndEKk
RRCjg+6g3Wd/osBkiMqU3lpm/Tng0ER8jSC35SaY09FLNwsjkHDKPE0D3f+VYnYIHtAaZYRxIgkj
lOjDywb7ndes5kndYU1ih6JYtg1AkBw/A3tZHYWlmVP6GG1rAZPon2f7JWtZD2Rl8g2liaarC9qC
SlLAVsOm4lCVwqeKCcsYJlT9OlWJtuII1LKCYSQl6rzoM6t7KA8VIR6IU+n4hqcL5kQ6Z/9N76rj
YVU8JlTjcKMivZZ6YsXlHLR6d01YXjiNPTpbdRQL3R+w7+HDHfE8yeHZy1i1zTZTMsFbSB/5Y2ll
N8fRrALnLB3xQpogJoxoqTQyGIlpv0Ez7WWU3mSWX1Uql+yKEUl6wdjey+WQ66R1SJHUXEvTyvhM
hpV8T/0dwIH5DgNlIBtyANUVSddJraJV/ZhA6mx4AVYop/4+tNdSZOPd0ryfcDjqMcL6gW/EIUwM
WC7klCX1fxExNL07mHs4GXtA6jZA+FrI34YIEtqHrfMhuWjDIcwdBDc2eeppNgkIVwwxlHjfVe53
jT3IehoIg1xRahQRdMjXKn9fMhmf3OfMQxfx9jVRIFatEyndmkCNBWEcdGEz/UwDU4VQ23yj/vNu
Z/0HvjUsuBcb4hP9AENHVBD0UrZBCMC2hbAVRGXK/Et7SMFWCVE+BBKeo2zo98sVX/nT03xAn4Sn
J4+/yGYxN1t85AnXWrCFEM7sMRNZBSBSvAKF5qGRijdbCBzr3PoLC2CckvMXbhl+OB58cvvGsPuC
w3W0d5UHdtbBIPU3cLgJiVTm0qZei66epo73CRMhUKDI7pfZsjdau8yg98TgGrQqJIXVMWf0LfGB
STBFgRu0o0wgfx74GPw85zCvRr39pVF4UrWzGI+coKPuTwW6lf5n9Gidb1jIWx9ofnvOr4TPIL6I
T6Buw+A/oK8pPYryFhPphKMn6qLfYL5GrndxvAgRaENe+P8aHAWI6AkoRaT0YfwHMVt2rH/Kq08L
TFAhGspx1onWNWSKaxnczKvpuZXXQFgndsmzUOyVYeGKf0ysMB+NxGZ5RX4Zje93GYJl1AscnUr9
8YqN/LpxS+lbBVgLnzhR0IAbXHndHIC91um6WfAg03YqmJ9Gd+DhZY7BhJi9HwbiPg6hjFjB0wz6
AUe8wkKvpzI8IgMzfcTiziIpFNL1xOb/5D6w+SBmFwxJqQjpTltaZ47i+VRGuyNRniFbbJf5C1v5
L0tdVw+kFQDOrRbt47AezOlaBDqreu1TAG0tqbla1zZyvJerPRbGxFTnnba9taq/rU4XnPFaXnlp
Dh07qmhJVtAKt1UvSORIqp54tBw90Bx+f7dwupnC8tp22QotnzUFiQoRLp6ChG1xJjvEGf1m7ChS
/qd8sHYxAZRuaN8pMYK4FsMNtoxXVLvY4PgF8FOtwEtKJZ8cdmzTwKqJm3edVNPk+eP82DF+yjr9
tnD3ar5rtQCnGHNuDpcSdS8zCJCa65g5s/kbBavPKhWDICeYfjm5tbuuCbMONvnKjuwp1vEYkdeI
7zPIA2D2uVf+bSHQUHWjeQofwOzPgRLuLxSwSbnlXPeieRZG6ugnprJ68q780LSxtpvE7Xoi/yeu
E6wAIlBbdBkldp8mJg2Utq9xI7FydJfle6VXHfGI9sTYrk0G6F7w5lfoj43e4Zv/XP/I4z2D9wNR
by4QSj0Cua/qjD3K46xIsLEb9Cf22l+FiFMVM15iDjEz7J32K7r82yLrdsGbAH7R7TGsPoucjDFe
oAqO+ZgJ97HoAcnJoQlF7++l7opdXTos7Ha0GGZ3jw00uhbIz1VSZMuZ+/BwQStPbikv1LoAmSwr
qD21C6Cm51jMKEVFgWXCrIMqUAJsg6DNmlYgelFtq0LPK9EiTc+seaJ6LXlztavH4M95jhGuOChK
RLaYJ2P/Vtf3aCCRfcSiZZTJE1MS110lb0taIBBSgBjQoJnwqARb+ntyTN+dpbvBJ5XH3ZJNiOQq
b63Keq13bvUoMSFxBqSAMzSTp0Rhgld5gTxPZtYL877i4FZNP10oIvTGdj58Gv23ynKo7iCqORkZ
L2WE6o31mNFzjuSHgE3NXHedZkqr4mJlqHfTPZsXwQ89oE72LxAqRDkrDKL2+VGSFzS34UixiwTo
0HpbDEf2owb/15teq3mjBZApWaOrQuZ5T9N8hOHG2+/ehI8gncL8terP5d+o/ZpSh7vWw/M+gko1
qMdGS0dRsNxd3pBgT4TasI8nI4bOGanQhJ/Til1HH5iR69DzwyDsLA+wkDWQuc0QhdRGk6joFkU4
u6G9rrEl/1xKAtjPsksrOTInA6Hb3CxNVBY3xjVPCCOtQ3hl1ZI7CmB7kanZUHvL2XxD9xd6sGNY
Ur3BTNfd7H0IkPFfaDGL4YhPDfh/FM5V4oDHZ/UDb5ROTlp/m082uUvVLczQcAneRMIwUL0Pdflt
Ze6tWO3Nwp/hx04ndwnObp7fWBzbwEXYXSzFQYvW9JbP4kXEywfHM1hlWQ3J1Ryx3SH6bdPKzT8T
aKriDd7MeV/PeJ0BfrJS00krEdOwmqK4Jh0L/NXp54h25QTyYEUVAF7FBg0dMq/thqhrveU6FCF8
/aROZ/IB2aDMcxeaYim2Qmnypdzw8pSOVpWvymWB8oTs5TSGKbmZsgwo/Em8T4vYrDNJGjsPrXbA
52ZyQXQuNjkJnv9cGfyA/agW/tU494dxBJysOBROv177++Gl8GEctw1wokgv96ezNXNin75M3Amg
RBX+PKo0fExWf0GfWQxrkWkMV2OgQW8PIj8Jvm9TQnsTuRfvYUjNL3f+b9FD9QUfy8CBF8y8UPhV
bN83OJ0ypq/Js7oRxL3c3EN44TH/OdQF2xYzYaHoxtbigQ8Lw4TQdWUT1jDZwAi8vlb5K4qSsVuQ
KYat4uZo3sBLXrmXfVN/uKW10hOfJm0EWDyPTI5SlpqQ6XNXHpfm7Xci2IBywqMufb1WRKieJK3W
LtEUE/isAUV6CGiSNn7qKtT9U0M9SXJgNePla9ZBFdvgxa+YdgSInrTyB6bUzsPaa4ckUOKJEJBT
s23/9BCYi0/5mbV0c51o+nQRVdMY+roH3TZtl5Y5r5isIIXSh6Vb5c2JxLDmthhXMI2k1qrb/ILV
9CY/raOx6rWC0pK39cMcCgcBus0/SNnnNxIsA/6BgP/MR8HcAqVhB317akEU+wHHnCuCw7FwGXnh
k8LhzUuyQbxfGt4aIeWXZl71dwtdEw/y+nAk97CH4XYvcY8FxE/DV2Me0LqvzG4nQ4fqxMULYn95
10BkJQtQBb2egHgMrAoRDZnMrhQRApxt74JKzBobIERzwmgkw9NHCPQ8RukpJUxXvRYpI4+WoAds
u7V/JtI7nz6dOz7/soEUYsG4R4G0NT/P5R7u6gOOdLqwMz1j0d4lExn8Zt8Ph/mNb63D08Sp1XZb
rlOFWNAXHq5qkRWCkhIp6l+InrdC7wmjzpKU30DSE/pU4OMfhV6gIRRc1muTjEMPNR7dJ3a/Lf3m
us1k3w/+Vll2DnNBtzAfDRiQoHktBZEM3gS95N4ye/VD6cq3U3UfZnLvaHfRHGKPAtAUeEM3cp0W
3QK3+Yuc7n2pKVO26LrJJqfWLIQPXLTUEscxnZN9L2p97rrek1qeH5xe2raoVPC6vq/F03WO6efI
Zy01mUsjgVsWIUCDt9Li26QR4HmWjWrLSOfmBbcfHUPinxFRasEhp/h296HbpIbMvjcPqyT8zqv9
X6JHtNOQWOpo24/K4327zURuktT4JBPOnhJbIfdhfhFbA+6rdqCU2GA4N7CHz2M3YW2Br9Yuy6SL
eOZl4HeWlrzktgevNr3p1z+II9rZivdOzdurkPP+EUA6pMCuXlIxy9Z5ZtHuzuFK8hbbyY5x1T7K
eKaElnnmran9M2cfXS/kHPl0dkzgPTg1evg885ehQoFQtBi5xTNRHNVgMfA8F21xShNvkKVyiUEr
9XQk//fenaMr6618e7BYv/iKrjf7blyExlgkfSbJokrliZU9ZH/ECUPnJnJPzCJPsFb3YXivOuKn
V/aaQmI80+dy5AwuwMC9O01fqGnO02PRcdkQYkuu+m0HfmWsyy0jcYNu0PgA6UeXFabUge2h+Ya3
GyWheF07eqJHD6PNA6C7gJP9LRs9jzrBVi5hA9sapXSC03zmfge096s1SUYuRcBKPwrceSCQy49c
nFEpsEqRgNkmlQ/axZIuCpyC6vdmekB/y0alZw2r7u+ylhSc6N2cNo/Irarti5pIW10Rt7QXVJyi
O1JOLwXt/vVOadaqmqLNC1BLMsixe9AySIG0IX9BEDitFlZen9cgQkrpm/CxISJlGSgCb/nN/RHr
gYo60hiL8Z9v0Znkri/5THlSlpWG2kCB4XlIlWidmRx5JiqIVAgRBpKjxNbC/Udpt/9zu2INtknE
4pHLMpWvS48LU3brT/8aXYySKIIICRltWCMZsgAqEvfkPPNluHyUyfhjwS30qjl6uk4Uq/HpgXx7
ABFffIjy4z9C9Wba7d3o3u04HIp0nRtypXis24hOfD7S8WExT81PYsOiX5/tJ0eF4lLI7pzGSkNn
F2sYz5EINNsfETnCt7cii+aPJMjgpjc652Ps9Xas7xt84DHs7nvNxRDsiLfT/KoItuf3KxKvdSTB
ofx6zKG+cLjbsXI+bhq/W78+IbXHa3QoX/vMkBLo8eBcob6xQFU0CwYxCqPAVxQDCnD2c7TmF6Cu
oq/O9aXhRfelF2rhkrRk51JcD8h3ZyUk7s/Qq9EBPFiqzPURkEpunqviByfawxnOHpRWDgKU80MK
Mu4XeHemAVvwYsYyPwtXHYtAuSGMc+g3P7tKp5kUeQiQZVXC4LM0Fi2mZXfhp+6NYfFT0K2lCUGl
KrsiyjMcZm8dmNYcnYNOB8+vRWo5p6bVNWs5B37SYTFmq16HntEcRvIMaARaiAbEU4PB1V4kr7lO
AlL+YJQ/deSZkCjHHz38REG/+T0Et4I25z3V3sq/5Rh2/Krb7ywSKLHf8NgSvBNo4lRbkLt1fJgR
uYQYGM8NcdCrODFKvYMTD+MSEVfICPZwkbEaKgz9lT/MMu61B17tVyY8pckz4G/6LgEi6lPV9AS4
r+9l8+k9y52EXdI04+K2Ssb4GXqQrvFTEH0ql/fwZsZ4lRxY70kXpeXg+rXt25NDzgGkQ0kgqtSG
3z864EVQzspEQAxffjveHjsl8Vi0g6s4e3eA9g3cN6j2mhECIogw6n8V56WX3cTCe+/LF3+4W5m7
bxcmJbs4CJxLf8Nb5M2myyKq3Ux7n0u6XwfsutpU4k96SvImfxe6TLxHAS/lFzT+msA/h9kq7rZh
lnSObD06fk8suYfeGma2/uOPQ249zExvfTJ8n83WVmeLJoiwUaiip3L+XyZ/cy4tD0RKfpqt//Uf
zWFcVhxAQyT5esBl2cQ8KXzgpRj6NMTtttHRFX4WSSqYpCsXrI1xav0bdrGxkINAHJMQtzLBTIWM
tMl0yfR3riO/BW3IucGAsWjOjmqRiEIONEL1G4pEdm66lKoS13f4WBe7h22vZ63qlxpKXGyW3BXD
Fp+iDucEHtHM0RW2uuCiVmvPoBYK5/gvSNOlVxQ0EQhm5yPkaa8w/GhFxu6FTePcVDQhUE1a8FHL
z9DaAMrQKTs9w94FFaQJ+Rn5hzQ9Ei7cXh+C3Gbeffk5B0FPwcx+IEVDEZjG7Z3pV1P513DRk0XT
ynRqIG+feKiXTWgXQ7BJ9uKfS+eS+ZcwnV1Zv2fS7SMR7driCjkvITd2ImiIdTlKPfniU3uC4mnU
cIy090kiuAz7BkPky8LD/6OYZUVNJ6Xh6ccl+hHC9paeX9M7eM5dv/M6/QK3QCY2ybrrhEOo+LZF
RVYL9xG0zj+OkCgBUxzmB6d6ZhQySnduPL01THmNdtQpPTu2w0hpprlaFzjUjvDrL+7BL/B0au6i
OOEmuft7p6vcX3Zr/Zi4zFwWDxavyMbiOWZ/l5viMaJY5ZojKWsqCnInGoLSYsA/mPbI13AtCfJK
HSdvm3ZtG5RPbdb+GFEj7kIvli592e2wiNa6cYkUDrx03Rv/feXaggveySxSoLwvgy1+E95muTqu
P3TZVEQ9rY6NzLJY40mnMN6HuWGj7Gintgkofqf29DljNlqhVBigQujiJQjoL3f+hh0cRFLMfnlA
my3fxGLURPBGU56gZTWldDJvWGna5H9VwVqu6SVuKHEDiQGty9FwE5/797YMU1dqD5338Kpm8AtF
WpnbkMpyjkASEjUU1+nieam0STXIW26fo/uzqFXHCM3LslVmRrTP3T9GmzB52U9AyK9GjvHLT6/1
WjUjqur3A520VSdNIxPZXzy5+2cTg0dBKvFxENlovOkKUUUo9kt0r0WywricHV0ekCimuTmHzkTr
qPEFYyDnkSzfZCRTZNWjcW3n1VawFhqvNKIxDhLYtqH4KgoirPNofmct90MQzZXysFEmdQlbSoeb
6b/T8FGJA3dEcRGZaq7uPZ0vsSLc7+ugLEHuq9fDWxWZUXgdsdvHZmJlnbEeW3ixUwyTLmELJSaq
58WLZEyQ1Ajg1Cgt1SwHqFW+0yiIUKhF2Ov1mqKAMx8w52kA8L4oDbu3qExkJT/1kEzURr1CsWlP
nkne7K+Mya3qBf+snpPQrj55QME5jkxibUG3Ot+51fNXFADC9iebsBXV2bvdmt2D+4U74sN2vKCB
lyr8AbiBJfPAo66cfOjT6juVfoOmO3M0sa7Bwdm8906hna2jm6E3s1i5JnkeV7YAKbbOh4esKl2M
DfjZKCWEN6SOsCUCGKCcLLWS1DZD2a6ZgDwb0wpJ9fJDrlfp6av0bKKUwy4eKdhMyvjzJWv8Y5vG
Hiar8wtsKNu8QBXrRXimzImbWRDbXc78iQQN53m5oUsjHDlNie+CJNDEpRBYZsD5U3LNXGCbDorj
NKKSZaOacojUc+cvIFZvwdMYP4zQ3xi+zSGr6ACii+swQ0OzTs9hRpNrwpsAf1nSG++D3ilxNxy6
ZysMwPFn2SvG+xmli/gzhRupAdyuG6We2xGjDk6bHarpdpsMw5cef/4FPXehpNyAQcLdLp+VLCNl
GGzhJIrvZzqduGbQH1mFt8kJq4GGWrdhg/jiVdYCWjvwy7g1/5ylQcOVkWO5KAnsZdm5gkL6AadS
SffZnE1NlKXq18YXZp8ccYc8SITQM1cSGEK1obk9KXB1mvN86ioIz+zuC0m6SSh1mfeIqlusKwEJ
ltmprxDY5K7iV9OjGrEIA11MML7/jCopUcnFl5rW9Ke3vlYl6DgbSLKv5qYlWuZbiwhiRjq6m3m7
lKkd92+2PbwtgFqGm3XDeNb2G+Ca/lM81OuGjjP9/yEmu7SpQ/GaLlV56qCGFmkzs/p3a0wRd5nt
pklPOShI9CuPdJ2+kLmlgv+al4CcNHcKt+NhYiNEqEOr0mOhNHwhhmK+7NLAD8e42nv5Y8UZMQdd
PxgijxpwYcLcErCbEBTKUesQRgVdnzJnFfNw+TzhIej8F0AOooo0ZvieA5eQn/R3u+9A+/jsi8Ze
FOlKehq/gotdhK1sdgKQfdx5Mh/iMDuMy4OyAWCcoxGxGXyZthf9Q4e6YRyzAdsQNhFmcLxlLInP
T43aDeYGL6hoO7X1U2vyeGsUTBlKkgSTd3C3AqjdvD7zxkwaUjX+LbNiFTLPOeEKUAKd2vHZPCwE
oHQGfgbVOQbBKVF2E+KEbc16+Z0FDAMmfrtz3mVz4dK4EkQ6864Xm0Sep/aPXnmaEVAz1XwEZEMC
DaH2/sg150KWiPD9fP/5PdEGM/IupBTcTB1CVW8P5EINvzTQw7W6pg80asEl8iqHNhvoWc7m7onc
TBTmrqX7Z6jLchhCLSWtwYmiX8qBCJLfHTdjO31MDHnoBXo2Nqyq0j3zLiYBvTzBKkW6hfou7d6r
YIkbDqRwbb7RM5vuzRVGGetuzHTvpzQDOOANv0EWjscXMJaVDaaIHL/UGDRsyGjWru6fXU14McPw
IJ4+dwGfyRyRhsvOhTKgxT9kY+COIR9Vq8frxp3b8uZrK3i/4oOPEAgs8VQ2d32ocCmSRi1KYHFU
TBRWcxmCLfJtK4vBRFjXBf+1F980PcPi4NcPuQLNwG452zbb/aAV7WG0CcatKIrEVKYD6M/BN5an
TIPPHMyUGIMvWNIecqS3WtIUL4LMrl3sgEfKD05p4YAI7UlXUkn4M3j8ypymcMgMS5WKuoShll/S
hxSwnoI5AbNH+kUZKG8WvjZWZcpjuSIwScy3jTfA1cJsgj3uckNVjufoclGOdN1nIW1zgnQif7J2
JvwJ6xmner+NByXSzMLrxSO7Q2XsAbdTzHBiVzY/oiwvxOUumwxc8Xjmpb+MSgXukdt9rw91N6N8
tkMg6gDNUv3ZHADCdvR1JFTgvNfjinnxugKDGtVzozNs8aEY/vH21nWZGZE+n9z/GM3VYZC0KHYH
gD6OC5Ky5mvEpNOcNo5sn8/Hu3UYFgM+3zPI68RF64G1eqaYUV5sOEkgqo6jvEd/mLu8kR4WBet2
4vFuZebxL063hTGHMpP30BOhNcE59Jzxc6arv1a+F+ftP7Bn0jg6hOyzVvXopTfErbtS6aZLDXdp
L3WTlWBSxUJaxMUzaN7YULkeieFJn0rJ1IMhjtITTxmKZR9IpSYeUVE5aXRn/U9egACFun0TK5W6
Z3f2F43iDsXyzWlTZU6rjK3vKHyKp1LLsAgS206pF3WSyjXNLr1/XsjqXIXQejwiYJM1VJ079OyP
lYSE5/F7pzgiHZ1rOPL6CiBWA92H9M278RnbZ8Z9ngT7SiLwwfRjnUwxq6izu11FFgfe5LCtqbEa
AasV5XQZg1R3tnQPtXR8tzoyY7RxF3qWqUxZ9bQ0kRG275eLFXLwbYIZEgeoeXcGZHQbWB1ffDid
B9fnLQxlkaPmJY52cZLVhNF7qA5IiSsUa+GItcXsSoohcexGGMcNo3zZeh+f/OMaRwqz25m96Cwv
TqoDY+uvlypppniSeQkOLYUXOK28XqIIVmSdRYlvWlZaN3s8oUoqLDfq8czaeYvK31tBReIIhycO
yQeMMNAXdMRwmYBsmLQz0s/wscoVJ39dE7hZ4JM+MjxhAjjRsykzzjGfGWSJ3BJnR3RHkM4RZ7aJ
YjRWLTQMfNQCVhKJXwwbwvlK7Z1xfOiJC2VvyZLAArpV1Mnb+wwY3rbqmqsRt6Xf9puWcgdEgGr9
1PKoqmWRlwd3mveebiTSkJ+XlbadSoGfGXfCWTcoOtrKSj3n+5BkYf9wBR3EnUqFtTIpOpvexdFz
ckARpwgWax7BlwVoQtR+NG0R/KePt4wQhbxC6RWzXyOFieaCuIUFEaHk9br5wv/s0A6FgHXzOBp9
SdJ4rjhqcJb0u5nnAsH77IartOwk/yn59pKgWmVHzsHpSnrU+q7cYHrzgFb2mwNOgWf3zNuzalq9
4oaAPAGNWA0Y7Y2Ztcy6tz2oQZamWHwd9Jplu/n5XfiVWCKxE55WbdW2QPaIbuZ/vGfwUb5q7C+E
ysMnXWLxmj8Vu4f0xP5SyO4oMbQJwELLMwXRKxOjqm8etUPmOYcZzAPq3nHgUEHJ2r28FdkA8UXq
B/TGQ9IgNbWq4DMObVKRRNsDyc2RuId3vtuOJ7tNXTR0ZCLnnYRgbm7PcNhDbX4ud9X5AKgMOySn
B/stmGyQsTBdwzcgMRNveeOiOE+IQ/nzLz4JsFtcMQP3YpOs7O1hdYg2YyYALMzi8yfbzhG4RwCs
hTIQUCPiwcjrhWIT7sSKdMsb5HYcx4o3kMf5dfpdW+u6YK78bFbA3KUYdZLhbacVvnvf3ygm8Sb8
1acZE78hJC46muhPo3UZvorYw9QcdeA/4ng+IE5TXJILXdc8Xxu3ZpkMEhWAeqcr0Xzrq8NDpzVS
2sBu94r5/IxPVooFexSYXCrOw53/7dSwuL8iwMliXByYFVYrE9Q+acvoJ0V5yBQNeyw3YC/wfEcv
kebwYLY/o3brapNUWWYnP7IIYYk0zoPw9cAziP1y4NXudGq+uJuEE6O3eNlR1r9smGhptbw5DwBT
GX3qZoQq5ILxShELZfdQ2tUd9T+DbrD4z4qXQAy1gLYK11Z3lclFzEK1eONfaBcl4fybXS7wMRJg
TpOqDNeSsI3DVVgkGHW0dOZs/6nxnOads9IxtBYz7EIbnfdvOkSr4LelDxFXLn9wEnlQQErcoS3o
/mUtW6+vpDoee0MU1v45j+7VRC5JaHUabcnIboyVSK1iokm07tOmfdZAKcRQP/x92RvmiAXrspMC
Df7IbRxB5MoR9GRvFm1FWKn6AjX/kowopL/OVD+HQXd1hMHSorChMLsAaQRaK1YdaYpT+bIqSu1N
4/b1Zf8aTiDLgB7uS7JDWuCSwDj4BgL65PemWTBvB64pVtttydYss9GQc+nEn/X5hqHLrorxUlQz
cb7kjFqkNehlFvqX9BMi10bxyttwoojmSsXVSOSyVCMiShe43dqGTeLhL1J2ivzgpZ6qcpgyTFGi
YDJALA9KmQvJCPgE9dMZTCeYsBkIXU7kRUtw/IAevnP7ib8RQ2Hnw9Lv2dc2sh1KI1f0lUZ9U5bx
sOH7NbEBaOYnF+V4lsoinjYPUAEdmSa9JfJAqzusP/r503GDHfTgfDNd/hzEN320DOLvCoCDrOoR
+6KcEIPfusN1Va7SYRKq0A3TFBrJ29WGWB8rkRXbdek+aRYTdtUhSAkuNLvgNbTG1+G/vvXIwlcV
bh/bGnmQ02EVT4UFfvNu9HVtC16UTkzK1jbrQ6xkFJ6NXQiibGJGTUP+GmjOF83CHtd7wrl9biyI
bsv0Cz1wvxDN86BpcX0bMM69AFC3D2z7z4MTeWibIuRSYCQNCcKhppT2xEJaiXbfVAckL2c1mBFz
uQa+7viOVP5TIJwx6Sfii/Egg2RIMBFPy0u9phhAjh1XT26hdhWnODIpXLP4bd6CWZedIgUu6w7Z
WvHXKd2zGana/xHSREuk4hZMnDCwoscId/PL2pQZIbu+cM0LsWoQzPj6r02SpK9Ox9r6zF13Y+jD
zyPZlLS9TEFBZFSLAjlz1bLDsZAdnKTNxBg1RKku39KHopYIewF6TWCgWIWzMH7HAscKYHUELa2r
h2SNHxFJCJ1HgWja7T+HsTuUZ6NuYLRnUnnBGVT52aULDXymMY5GjfWx/+7GR4BNUFBYxL/kzCHf
IOT2Q3zF+IDj1F3OxqjFe83z//NREUBJdE4W8uleWZyCT/KgZLCNgnE1K+JJDpJjJwQnMCQqjaYT
Up1mGdgb1qXxNsbmJ3DyHwKcRaithl5rs78qmXV6B4diIEOdaIULyTVp8uTzYbUl6gMK4XsZd8YO
EyaEg+Im5K6Cf9IJQhpMLJt9IXKq0eBPTlp81ZcUUCahSx3/ybntPkY4y82r2XO1ZKnSflETGwQ7
UpPmSB77dRJLAbPYhTOeSnAEXfRdXgwU8W7FpxelGHxBPBhx1wcIw3DsxFVcXDb0yTqB0lkgb5nK
8B13LDOmFiOxEuiSo5XTJ1k392Ke24tcS87fjpgiGAJVuXg39uLoo4Gzv4hMwfM7QxVuZ2XJ0c3m
MPXxwGzhtiUCZLBDne3FvuFQ6KK/u1ZKaj25lzKaa0DbK6jdKMyaXzwN+HJqSiKV5NaI3Auc9u5x
EgaXRf5iBquMUrdq9Wgftx0FLUSwSLiKy3AxoFbyOOXAjF9OAOSfrpXa1v3W9U9UXtzRmaYS3hrD
+/HvT80ixHE+llKMwfriYlMN6mJD+XtBikRQDh4lmS7S6LocV4b3ZV5IpBIM7KuFvIQ/faSFBvSN
+eCkHVVEWc7Vz3/IxHP+4prwnqp68njLXUNqoMh52YoIqVnoDoHJ1OcWEKHRSV2QwLeV1rOXBuVH
h7jefAOSY5IgQdh5TnlFp1IVFxosaVX8IixYu6Xvh8dCXuZY4KrCzT6OaNeXDhxjJRNOcDKliz2k
LEy5arHBmpGC+rbDUm5JejvU7J0FTgTutlQQKRyvc3M3MMa0W88T33ppnpbR8ihUQH5anglXzMN3
T8iz4RW1ZbDsd9Pf3apWRBrXoMsEZs2hArRfeNX83P7Mm29svlEHE/WsioNK7uxEcsCPxghEkd2H
mHbj/msy61JMBNgdMog+Y1AWlz3IXO0gowJCBJcPEEPsNM981jmii/3o9Hzp9J4d7M6GuS4Ei6Qq
2AVMVbQLNf0FZa/PMDPISotBeLctEm9AtLtnSuQdWPjXAzd7p0dSft4lBX1+DfUTNgHCeqhTiSO+
MaNO2AlmC4n+xz/DAlLx5WAsnQRp32xknPRSC7xJ7t1cp59pBbd+NhSd0dZG2c8htbUp8wM6YGyr
fNFJp4NwM8ruworIR4K3ycII/Xxfr7ENbP2dOQ/Ysb/waez28+OVO0PyAwWIDa0ELytRvmQ1Kyxo
ZnjmP/e6mJLqMgWTcllK4EFbH3B+3fawBxeqNwc2nxoaSKR+N4EGZTVNbe8aDG4Fgq3mqCWhqpid
cxIT6FEf9bFB2S+BydccIv2/Kc5s1m5qs6U7cR61HDo25QHmoL1wZfjmsm5VvJsUjDmY7QQUPX8L
G/gMIKvY4XQCfqmvdV43ninjqNe0mMk+AOtkx17aex7xm3bh6D0X1kNRUr1FiZ1DAK4kPC5LkIwX
DPUXDqP1YPtC68WbABX5a+yYMqr9ozPckDBuBVtYH9cl34j4D+HkhOxige0M6tZVw4T3T7KJvFx3
UR6zNQZ4Cz2ioL8kFWg+8d9qSe5pBj0YjuCVZWhy75i//kpnig+4WmKjYLQs7LLn4mhAhNL1hWr1
mQtigZTx1JFsCnGvPoZpXQ5efGpvNJqizuyB/q64XPtzRUI5gsnUxRogvGf+ZlshvmpqVNN+DbeD
T43oDKO2YCMuOzm9u66a0JaJVGGeA6W37KYY+mzMH/gl0f4s/E+po149iTsEcMoFpNVwEQyNsxpb
6aQ/RMF2shfza4wFTQU4AmhiMByfnFkUa7qBXmAvZO61HkHkJH4RyYiInG+Et1nFmC4MUYkJVvY+
AIbk0O/CBE7rS1v3n2twdYELJ+RbdePGV5YrPRqk6XmUJfD8AV0wXODRLdLVnEUqs0h39Z8nrM5J
234na0eWvR4XYcvrZ7EStYbSFBBb1+Q9MHGdk7NaKbCnc8DtdHHU8aNhxTxmPlFkA0wy4xuoLI/5
rbrSwMUxVyC4cqFdC1kL8G5Lh7GDeBPyuPczuO8r++IzyVJJ1f7Vb+qt7fbfIPr9+6z9JsuDR8KE
afS2/wKd2gSb5xxTtv0dkG6HJ7tXoIhcXwrjtDQlYLmEMQwgBisMFpv7fdN10cjc5Bh7JXIm4b8h
/sQOdOKJN1PDyxMwQ5Ey2LBvEJe3BfM4+/QtLKn1i/Dh4tz1hrFWiDkSo21PomqnmrvJjHGH0bqg
P+n6oFemykC/ly4z+MxxdLAjHT+nqRyNnhZTFQG+6cL6Oa8EqGRTeaNMqj8bgCnmJqU8jG9A0Zv0
/47SOPFiU0M5FJw0KkLzEIRT22DOpMOTpXjSsf9axoT57SQ6mUQVba/YUHg6UCYBA+/5RaIbXmQW
yHm9pCMYJE4YohU9ePXnLqNcI55yBDCbaI0qQ/iz0e6tl3w/leMWmdlze+1mDNYb+fRMZbHXD1iP
UyJj4P1hGu9DmRazvimZgf6YI+p1SAC1vcAKr/T2mSzhSRh4Tu1LVZjFRV7SvLQUah4F5AfopNrU
vx+TqS53R8KYEyaAFm+qZEgsRrI4jXabBJWYLzysz2QHGvLMqLnRPSAvUdQeF703/GKckviIf/yb
PMN3i+oFA3ScMDwi9no2ksO5OKtX7FSJBmnxLdOvnJ8aAAwSHgRRQemm0BLnwuFDgA5c8ZDoopqu
0avqsSfU1e04ZdOxXLZmuHs0GDSRXMoRz4OhksEJzxU9Q4LeMzE2ZatRsiOtaFGMHpj+VVydNx/f
qHIktrOI5DTGhMIKHwvjpWTWSus21xb/PTQKT/1jM3gxKnWPl++wxPNShl2W7Yyf4mve1COPC2Im
u8WQwmsJMGYiDwUl12rkWalMX4Bb69OnWppsHxmmf5d/OlMl1LegyZ7txtM35Hb/aN6cuFnRPeK6
kymwyA/3jvFuQrKmlRflcc4aEIWrs7ndmpATbGZsQclcolaPNWMXG5UvasmahoFlXmoJGTSmaIgA
GUH/RxI8ITHugV782AZ8QyoTz/1t1+HyhRRnGFgzfDcJXa20KV12SMDlFPwBeRSAlLpEOJ92n2cL
frsI6o0gR8haUFCDMM/IFRuMID0vNVfiKzj6SlmG3x9rXg7/+yJxBTcNSb6be2GSau1+lbr7pMZa
Tms+PoUTt7rdp2IT5f0/VGJC/FwhsTuaqOmi0a5Cw9oJCFPUBn6Pq1slmodCGo8Kur5ED6NJi132
hTsIYJ/NOuMdj0xqmG8f8HF6deXaqdkbFQUo4xMkozSTtiT+MdPSVY56BbZU4zOBFxMMUHIkybd0
SdJFU4Hr6P392kTz5bobqkKHL0tWqrV4H74+MXqcK4A+2Zgy8zqbgCNomTDg+ZCYJXp+jqguJpNo
DnVtuMiNvitLzlrQzZjQlgLkd92gu4sbjR+M9sVWfunNAeUwTkW0KM5Svh2xGmZjhNjWvOApfkXJ
fbtxv9121gQxHPlvY8vZUrh7DZPlU34VhaP3GPc43N2Qr2PRAFI1DGyd/mhYUC8yafCcIp7tVj07
AS2sCdUItsjuON8d1zAYTVtxY5Ou8nHNLCTU2MoE+AYNt/QtHPCBVBNKwaEV6weaaNVCEcECMTk+
W2YbQ9Zo/i+k3uHQ7tFyO0N4iCtn4mtYAM51LqiOTMHYzKiNYbaEAECs44828llufESKdxCTd4aM
niWhHH/XZkl7KPXsBYynFc5XLh5JBmwv+ak29IfXq2pnOt9fpV9ia2BHIAD4hc/krf0jInvKwdPw
m15oAc/9hQJkrj/lgEjlmKm5negB5PkGlZfBBpqDIgcNy3viueLvougWRO5RkJyw7oBb3Zt8OiTA
LnUMU1qWMoOHuCdArCY9kXgaUzTi2f8XtNKoph2jK0zz+RRIMcQQFrfuJO6VzpUdrvHZoBKE8xHH
AKxwDGghKTiVq1aF7ADYcwsDEY33QQBJxJSbOohk+l72ZUbxNucrhPhL4ffAtyGz0pBKgwEcCtSW
A6hIUfsHQQQOVWwuUI5cQxyMZ+ALZrxmC4TydOsJ2v4CgJE4eHBbKZooLEsCvxUg9EApkzougGb5
al92b74dEMGNwqajxIHZ1TlstrDPhmcZ9v5aosbEsQ7qnBGKZ4FlSP7SjHBFSCUOXbJN1z9zqi9M
z3Ijxfkf8Ijki/jsBW78MBQaZQU5YM9uch/cfwuIbroUMK8K/RkTtMwftmJ85YL+oge8aEr1Qdrn
ORyAhwSz62EBQLyhGUKfmHVKObC+8zV0r6ylxCUEb2eXWsW4vNCcxiZnMlG+TsMRVtTX5rz9oAKE
JZm2dF7hO0OJyNLQPUrU7vRiEXKzw0r8h0XRpoBTS6wHMfdlgdnb56OtrVGaubI1REvDHs7LQ9qr
XsGOuDADBedGCF/tcP2+D6GLQ3LUs4LRHdGzSAt7UUJHEez0N+osO4DRx4u1f847rPrScJ35uQb0
YDIX1FlpOGmLQkNZv4nYd3nDanUPvJzNgYapUHQncG9Yn+W11OV9kgK++qN1QEZCehPYzmdDfTSS
ng/xa2goT9fMmir8WQfo44jyzrN9GaFrmsMYjbYlUvKsjCyYWtbZMIRhjoZ8TiJJqIaHWcL9dYXq
FE6TPr5kWX/sJCdR2YUC0TEtEReBdVvsOzf8oLOC+w9TpGFFRIFLS6oakG5Bj9n9IBOawCUtmvoQ
CTK1sRiPFKyS3NONAcF6qH1tqT+3VyiPx1RtcFnFFzSIcTvr0TRxEqlse0URGR0wFvUb3wtAiFFD
zwjD/kkKCfJx5UiXfvQh5KiWNzxjT41QcIVyvELl3RCYm/tVxZPGtxYZ7/kUNrWXsOAHt71z3W9I
EkquFUaGtRI9+I2PmH2yDOzccJYqWzL7LFHrq903vxP3mPJahQgbWVO6gnpqh3rEHX8Hcvq37zBk
dYdOjxxNdWEpH5UpVxScJfzYFqUFXYG3ZP8gN9F3b5aen4VSRJAqqAeZlC37Qwt8uFzH52wIjn4+
4Qg3Ia14vgX2ZU8I+3NvrohPPA1EQ71mhMykVrKdVYG2aHKGhrECJPckr+Yhs3tooexC2zXGBqz6
+5d730jm388ZJ7d6owRbiP480NLV64uI665SnjInK8/Kr5qUwh64aR1+fB7Y1eTPVLnVmH1LltKW
ao3eql4p1jL4ozBIsmvgYVAELTC724+xZUsc1TRzyIMmb0a7qBB5Jm03WpEOWQeycgTlh4H0/qcP
mTo5ReTJ/GQxYrY4xhk8ZAqyzRjzab+eyNQ/k4fgQLTtvjlM6h0PvWkEBeF+LyAOmj3iHZcHUUoz
ZwLMztitPi+eA0RhgnfWBWSr3Nei9HMtwLW3AAYQa5qeYlnKpsnGovZ5lkxNnPy35zllR+MES2ki
3LBeYXA/M+RxQYvwYqA2nvr4BYt2lzhsqR0rT0uTn/0uvrhVWJP08oCRPq/OBIGg9QkJDKfebIca
TSEapqkAjcFTqH0tLWTnsg9H21uIF1lh/1k9qzgsVJn5baXWPGQ9cDFcn+sPFE2X0iY8jENOwB1j
HLiifjg0CHH9NOp4dAHg6InkmQRZ9fKeJubDh8D/DmD/z9KUO80UjYyIruSjBbEUCjRVL1ezEocm
PuiCtu9/1t6+2uGFTgsBioeYkklUuozLgKL/noQNOF09lIEaLq6wNMAV2pSoNjKKckg8p4jvHac6
pJ/hv7naQc23cTuWgMBEkIkKJx1+Z9VzvA67JZCY2D6BJB/FfPuy7TqBdCmON2EzxkTGRUMMmUJe
R70dK0Z9en5cEUEhvrLwYX3Yxf8TolxeQcwY/99gXX9LyS8Lpo+AoOrm47SCvDd228lSwD5rY8QU
XcrKvmZIJXJ0QP6N3aU6/nJYRG3EgshL4a+JiV9D4il7WSWZMqBe5gSX7jB/UL+Tq8RjKeoqTjXW
NIsaAOoCs4ULzKjEcgqlSibi6LQob2r9pX0rIITufu3f7r8MQymBDquqjxluxLXf09rQ/wQlQ3Vv
mAkVytpVOh84M9Ka1wltJTUGi1MkOMXx/Pgfn2ldwhfAmELOkE2+R7iz93Oug1P/LjVfoKJSSVB/
mkfn08OV0T9gu/Y3IP3q0RfMkZviLmSHrsHPm86eie2hDUCmTbmKFc0HrR3S36bFwfNpz9m/shYj
uroZ0A7dxHgNP2kMZBNCLc/AViDJXM+09PM3U+6ru3QJiS7XfHVidt0GRSe8HnqOm994ApqTUmVb
s6SLaUxdCvYFAB0vHGZ5OUuRqTjhpsmKFqHeKZOdNU6HCbvgSFBzcjN1kkkOXLaMUBBXfSGfmJGZ
7eOKcv0ZGM53vsSf45nhxk/fLEkksJ2XQbYSd/rM5SM8o0hOEt0HLkN8l+tuemMiZeUtL558SmJV
UuqFax/N1EvlbYarXcIbCL70IqMe/AxMgqI9puHOmDr0SGY9ex9rIEwYEK8RRknZrZFHK9RDvjJ/
4u6e+yqdMsqMHbJaKkfxw0a665KTyJEO4vy9jRS56BNW7jaJQF1dR8+CDBf5bHGAxkxId8ecV+AV
BRhKqaHCKd0nMEVsDxLrid5f9+mmq2Oc/rIGAzuAXUED2+qpniZSeumoRvUgi6gPzKNfugrxKtT2
iOo6fd2EWAPeEBDaW5hEkABKlHJ4yAh8LkSWw7+P6OK0Ulq0A8mR0g7d6cdHQlGJ87PMg/6ZhbYL
6astjQlNj3s3ss5nh9aZVd38bRRN+IDW7sLPTkbT0t4c8cS79cY+Me7WVJ06haEaKalcwg+AfJ1p
WqnVRKZ5JojR947AtVsKOCEqiYObHupXop3IyFpueGc+Yt/8HdVxYj6hbmtXicq5PjOd+FSJNpvn
rXV4+0/oyKwhd8aIyX96kYaQwWCT1hPt5Vuj1iOLshy/H4qlOx/3r4FC1zbRhpSK6en/FjVpPdfs
BSftTiuY0g2vVYGAZ3F4KMBwTLF1Bq38hbrx0wnYdVWi6/HMNYMFOS2VIlWdOIza3iyKrnqqXr90
pcOvQl4DAhwMHzsidKdZ2lXP+Mp4vZHOhil9JqyIaBeUesm6MTjzZYv6Ll0b3YgujhXwDuRkvvju
Df6WT3t7X0PvIJ1YX54A6VRPJuzNXCEGdzqs/4mv54Geu2vBpKMOQ4FXVa576AaCUukmvFXcgFyp
lHIw55w9mahBVVSW5qDhr1ZU8Jq3DadmxlfmBz5KQM0WYhNbrEzXIKmD3WiRDo3sNwZc16GvxS6q
N3jpN9ljbrXm/K3mYNsa04EHFOrl/oaEDtDO/Wu23HClwmoG8aMU3fwrr8UERIihO4pdfw7ylWv/
yXZDfbGNaK1JOdO33y/E72Ff/PPs/ndq3wYC2SE15TEb55M8aBYfPslBXkKKKdM7v27p8ZIfbTVA
YIO6i/5P2Frdv/61QMGuEA03gxBarWv35tBT91zOv0FeCXcvJlQdZaIdm0JmaPCQJT4oG3QDr5XC
O3W826XeLpeh/eIYqlxRD0eCT8sQmHdq11iY/u53ID42G2OwMvlOuly134uzLJaVLn94JlBGu9x/
ZKXVxP3qSYd+LBS6zfL/44lshXfhX0+4Bqa7LLLx8NPgSnHE2H9mie5RZiOdG2LmZYurSwoOFiXr
nKCRVJLNKyD77u01lUxgWlBepQVBINAZFk6jSW8k/uv/15ztYv1tWLZ3RasVQAIB0T+/z/Ed521V
1FFKw56GnR1ZFmB9tqeq8/FnnK5TfzEF+clTfKGU4+HKvenNp84bVgCw57y4TaKygGhmO24r2VTw
cSSMMMqVr65bjCByvZ52azj+E/ZVWjY13JqvVmRQBQPXcLUru8TUZgNJQkwU/drF+G9DwXSkJ7WG
fPhPGbDUjsQH7Q4EJIOx43OZrEd5leltTOL/y6AA/BP3KHHpIntLgISAi0gBThnBK17VZshfkd0H
cqqgciZ9XBEEK5OvEOFEQYnKFwP8tbv1NGuKTyMeSlfWGRnbApuftREaHCTKonC1UqAA2N/0gs42
Uxp0eKTsQoepfrt7DaIw4m84khXslo4lLjLkIqLQgPZC1GmsH3L0y/vw9xIoS04uE7YhfzSHthoV
M2ySmN4Z7Jh3tRIfkHAKEDCIvs/DlysMDeSUzNYJ5gBqyUXVO2nGH1uoApG6b/DqGlYT/9A19DkW
4BlZRXWvvJExvH6rK7G9l/wVNnqRwYpNfFHHedBGViePOah9IPP56EhBSoqKil3qGvQrsqxnui1g
FubnAAZm6JcF3opvUckLBK15xtEi2Ma/xuS/PaIOV0LODUvJXG5TSR8yv6XvKai+qI4tJ+hElq3J
19pvC3zmfhjxfa87y57ooxivGayAtlRSuzEYzniQCvs3y+OzAbiRK4aKy3gr2EZAtbu+q2IqMzN7
88G7xVRChiNHWl7uZDOHPIiUSvoVyQ3HXQ16ROIukql5v+HEnHgXiPuSHcRZ9jeKBJR73QCSldiJ
KjAB9JddGAkXved9FAJgshIr9YvhpU00Y93DN5vjjIYW1F6lzI6wPNkvmJDmWoaM+O5Fnwl6SSUK
KcTw5vGvBtzJasPKwRWlJuUwatnEQInYEi1KTJoJwAVvn/ojXf2cgt25VrcO1Z9WwYddOB90LnWh
J/dD2Jd4u8exmR06wqvt3/kzpirjmiXRXsc0ab1e4qqUjFvnCqEvE6Wl4Tn5vGgH08Mbsek+3ekV
6t3dzBFXMsfdm3qBYBSmNBDwvOGsWO2gxQve8dnd16RsesKXgyISutuNDUrrA7BfdCb/xbTpvemT
BkQjV220BDNuxlpS8YZGsJyFEXRS7aqiyD7IGbVW7da5CQVJICJ0zzHkIbkFpVUaWgGQ8MdP5z2W
xt/OFkCdEhRFlyk+1/Kvm3VYctYSHdDLVf98ZOSBOXMMEYegFvHfu5lxiYrCpQdkH7oBsjiVCOvt
OBT1yjp18xa8EgsRjJdgAurAYl0MABMJbwv77bIf2D2EVVl7PLinsjMzjXivVSt3RX4b0P5T0SOO
029YoS8vErEOaqR5B9YMtWIqk3NwOJglsJ9bxWFpsqCgj6qaccfxDw+81RH6nGZViv+4lHv/QB6/
UPng5IKy/BTg51mg+M7vN7xpJwX3rGLJ3Z8llchSlkZD/UFnaRit1wbWj9aJtNO9MQ84mOlXaoEQ
W+TSLl2nhetAtnv6MlfK+BT54GHgWodApuSepPgsHpW4KxeCk2u0qhuOBeZPo2VNNBv9y9IBir5V
WNBewZDo0MYHCwruIFgwy0UrElHCQGkb6eCPze7Pl3rnCXHtGRqeHEOjdHspOk8XN9p/K10ygtHR
CItUgtgx6CkbdMG19xlRG3dvbM8xi5fwS2hxxoMPvQ+4W6EpyDBm99K7qtAoKX4B/q24vT2tC8Gf
tL60cIeFwz+FlTTFLphJAfnPw2nWwrEMaGM+6QihZFIxGAmq4W4OacfypevuJGMNV7V1bf1cg845
2lxQ5zTJff316HL6D0we5AFCymGuzyA38BxtHvZiu3KfDx9ZyeEIWtflth5z4vwl0HOV63Xq04fc
JpXygpRxKIr5bQvAUMXnD0hc+AFzRPlK2hybvwK/mKqpDPJ4fgdoIDX8rZ/TLGNdFIOrVBcAXHq4
9saGlUJvQxw+/i0XTIjW4EC/qv7Y/wsbvDywHxcOc7s5JlT5KNcLejQIn9t8famLH3sFeGWleWSH
l7V8ek+YeP4YmB9LQy0UKPIqt4NsIvEKmsUKU5EEucGWbL2hbfSN8eUcHWSm4sTOm6fL5u3DD2wz
S8lFtRI3d4t2pYc+QGyMzbbYjsA8dQTcu1Zhz5jOa5j47FEpBQskGDvJCTx01yXUDzRQCKRrXsyh
gSRDC3/LymPkxYsVq9b9wHQHpFzEbd1Ju3kU+zucfLVBbGOiRZTbgvM9snwXYzPDwV2rdfgaz6kc
ZHxU6XN33D8hk7EJU1bwD4aJPcB6V+FGqGEdyJE8bueRaJpoOG+Oubp4k1+xoacm98rf8GMbPr90
c/COkZHqu14w4qOMnHgDqxHwQWEPU0aWicQsXZajP+axwQoz+dBKMbuzNkXm22aaescVTgvhwFEG
fnYU7u6JuDWs5RrxDJ0QftB3aBPU6zB0YWmztVJdWHi/CQ6XcPJP07yHvm92StR+EpSFcHsmIJm0
K49sojLcerPmySBGiddPOcACqN0r6hj4AGwY14nt1auaYPn1goCcvnc34DCAOn6W8/U65fiQYg6D
lC5pWoC9MDO/1xy/tBK1zYhSlxTsoROR4i+U/tTPDAQmBU4EVCLueyv1sjoW5jzy/VL9LYG4irer
P6JmXQQPp58N4nPzaU7PyC8UjVlQB65gZY7rJdfGlUXg29knQBjXn0fnyJO14PbVL/qPh4K6NRFB
l/iPyy4fmTm3OvDud0cfU5qmbvW+al61YZra09FF8sGOaz947/6f04/oRy3ILszwUVUAdRVDYMiy
1ADUYoPak0iZ229mLNO0ZnI31Ehh3DV1knEW9MBq3SDxc7+gnQmUNKzLOtERwKKSWfYGieaL3DuY
8gQ2Kw6y41scC1UtNOkKYhHf/AQD0KGL9yqTxP0XlXZaz1VpH6/ObkLwcwzPRtiknYiXkbx6rUxF
r3pEblYVXc7gds7NZPW/DLJ6iS3foVC4H8kBiz45Y/YxMe2uW0AeA8WWdRkHiuucKmEQWlQwZOzt
4YpwTprXxm//Fwu76Lh430Wq0R5i9oodfTFWSSma8aSLF/bnhArCA8TaXvz+WXStHF4m1SAUoW7S
htAig4BIkQPFAFD2Eud9EXzzAJDF4LIPqx/9oxsCwXHhMN+UaY8PjsyrgACGxIdzsY14l1XavTzc
u/AjVd+Bm+1vo1i/mg5u8EKahGgwK7ovaY2NtRkrUtmmaDE/ubEW62qfXAL/Sl2iTgz+4XsNac4/
RFgSxegopYFRRb+1C5hZdEUYIPxfWWtmFioG1xgVHMs92vaBfXr6aiLHlarY+XfOdKbbfsnPjCTk
moUO9hHNZx76M45+DU2HzsxncEj9HSM+1/tYW6CLsE693SCyKmjxqfObuWe8JL19nVrE19ZZVPt2
3c8jnYFwAE0gQMlkSXovCExNucMSQWaGBkwHEF9fSOAPxYgrKiF4fgxTz2s4FJtWCVE9n4CUSwYo
Mwzk6GL2EcbLgWhfWN1rOThG1xSnCYSjUaAAFLQo+ZFrgZpL9NCTVSCVlff20vqtcOpYzJTe63zR
DHNS8i8371kcspwiuLlfMx17jlUTPn2wHusWXslFM+O/eewF2POiRZwdEMccX2gAy5czt1jLwvJc
/zjQT1cabCOq74bTuOSttAd1VRLNMR4CLKrCelELdVV3UF933Os+m9gH5NniexBHqFVdpbu9H6CP
RAkijAaRWtNAeUB+5/jm4lA2ukv2RXrJk1YqhV0kVg4JRgOHij/0rFJU3boY3DydFpNbZxelsvgw
0jM20NdnPhbsg9eO8GeeWBSCO1HQMcVzlIb5BFcpYhOKYx3E2JXia96f1H/m6SYHhMuJOm9c6hjM
Q84pvK+2Ze0O/RLMSe0il49a2O/WEPeY214ESmQz0xnIttwbx16MWjAxAkxAug4SLObaI2+HNUf5
UvQJiDzVtkE1otxDLSkp9UgvCjm76HTr/XSSgHZSBMy0+vFwDZ9WYsOWG/cGMUARmmx3luCLUnyj
jjobdKtqTMrAHeLyxcJzm5Xt/QQ8hbjcZDBgxgHt25RTaUyBUQTnNZ02AdPRbusuV/R+yyYQHyNS
75yG0sciBmql9R3/+biR4bFSH+oTcQAFzs92cvUc0WTWbalnF8ec8MyPMuAntkCHjC6dtKJw9FiZ
NI4MFvq0DqyWdsyTkLb0sKmyvr9qhEM7baWdQk8pP5YadWey0yoZ5fhCP1sxZMYhguK8CxYfsFpr
tadZMDVwZ9A/aZCVAbPYKREwTThdpy7Zbxof9FkWkQE613fYj88vK+D9XrV0ovis76CVH/hFCInW
6q0MyIt5GgelIGpythn8W63HfWxwBKmpB73lI7ZRTYVAmW+y6938LJN0QYSjxv5QKFoLzD1xCfrd
yTWZhNKkfVV8YFarVV5o/3Ew1MzGdChLfFCNE+yS5HW9hw5x/5xfeqm7kY12RHM1QEPwQebmv3le
k9NWX2obZ5L7a0S2PKz9jZqKHQOR0GxhAAZ1aibCaETBC5dJT4zxZDIdZYv64G1v5BXoz/NWOA19
4g52jp74pYJejxjqq7Zk3KcaCywIlgkCgvvFdZ7hMami7n4bUm+y17NxlGfB789VByQuOrPnBlEv
rhL9PYl76/0vNEyTbxkgZASYq9IVHjE9CSkRZl4bk6dUwTyAqmCIa1mHQdIv0xXFNUbwjlOYEiB3
V0j6r3QOBSXix7q5r0fw6cDSznSQn9qXpKwRl6hFb7hHPvvji7lKXWGpeBsvmWcwhQeeqSha3pmQ
GmESJKBiszzHHtWqk7mEec8K5S2M4se4RHkkl+1awQ8DHcwlqn8QhxLLSNlkZTj6rwnU+3PUw6fM
ST0H1ASisfPfxkOkI6LiGZGqW3m8isp354CUGqIGQ2ZfXQj94NnlBkwohtdySEiAiS2IcbTNHAV0
HN2gm3AqTGVG5gENr+vHEqJbTbI5aUAqPv0cVtPoeJ1362W0w2lH2aty3DhHbt27yeQ9l3KSP9CD
hN3yF3uBgxEFS5bWrMMEuMyyMRSTgUejU/Luh4rFlt9iMzhG+iNGb9ynUhhqMqqYW3FUHvEA/9TG
hV3sVgRc5ZOR+UxPWM7zyGPAmbi0jgLgE43yYKqMRwNT9mutJ1mTZu0ZORcFbA2GUbn/nZV+9n1H
t53Rdzsa0e2qC6c8yKe52O0bDOxggSbp/4oA7i1yambNFmuH/Y66MKX+NOBpruvsRXw002h1i3IA
qXBrqwKYGndw23q71XZ4cTSXkS7CL6BVT7VLkukOzAhnBV9ltAnJEe3rV86jjoIXARQ10LLDFamY
/Mp81hLSKy4gKe/yM8IZ6ye5rgtsnIvArj4F+unSHcLE6Xw5YuZuV4gDk0XI6RJwleBaXeNCFAze
wjrcTbicnuCeB5klLVWziWCNlAY5hFJFzr987M7z5ZHdcHwPR3GIPPk8Ui0wZ/n8sx2+XpSNJVTZ
+WqjIftdb6wABeKkRSJoT1WO+wEkUDUYnWMmpVsOLulNXv4Ygo8Pvshf6vMJz2IiBOMY3Tc0YKix
s4/V5JZV+NBPlcXq3//92/9Zf//KvZW1PNeSPdQ1MtApfi1gIkeTPEQVy3Tp6mlU8cj4taqr3hgb
7azRHCQnr2UPofS5QDLnW1TUe8aLFXltvuD9Jrg/ewtP+3nIiFSDRA8NfSMYU9hPNNUM1jHvjdp2
A+nVDuZJjuy5994j1z3jKFKti1WE5S+pSWd8Drffvma859sxO8QLHCFsmX7J2I7kvIYPTNwfHr/u
rCK8BsuKdHWwCe3WMbR5sQ0jqKZYtTgPHQS6Xo5+uawJ5xON+zUDxei5vn1P5VPPW1PyprDRE50v
Mab/dqF2nWFeEY11lHJeW1PhdrHmol7rPDa9unp9Kw/mn1/VkMBnFHzIlqTVyG9z4aqy3NqaaAjf
G1ARu5HBrcPAAbmO5fscK0ZC8PvTyrV3mJ9Xat2TbP4RAFGP3sdAAf4jSgDQdepsM7/l9LPAbC0l
/VQc8klrTQPKFIrwh6ActXhYRjv17bNSWFt+JNTT17eEywGkHDKXFDKoPAwnIM358sslOtGbom/w
xe4kjvCmEc2bvoKw4lT71l+Gk6DW7Ftz1yF8m4yjxP+sEee6aOPUIH2hEpHOgAm/uXReb7wYJ200
+RVyeX94Zwa2j/LHhv6Cl804FJnBA9xux2uCrgi73f2L2opMWh6DbN4IuEAtCLTLEDKM9nJ4wufM
AO0tIcku2oV4EwMwKkUhPltsZ1e9LXHVuXlFgxRs//4tUf1OP/14b2CgBqnXH9prLEC9+SfJyEWL
UahlS+yIMmW1woHBWaDf/mp5VxXPQhV3UlBa5BrXaLvAbbTa5/n5KPC1czkDJgV2hkZMO7Rmy4wJ
mwmQg5rCLKBPBVsikMsbkxMFLODvU8C92ptZp3jBbxv2i4B+MY0Iqh/nJICpjv2Y6XiY8ExHTVGX
ezVHq9ZVJXsb8+owczq23okDxGG9Fj7vi30SoK38VeAFC4WnaG4+u+EEHdKdXplsT1wX0HhEr1TA
uhL0jJSxksLLS4Vi8svd0yzvVhPYflkatdBG68ZyFk81UKwDaWYBU8WqdUBAkHSKEMAXrl49H/+s
OftSn1FJvMPtyt+Cj+t/Vsa4g+djIPvciY4OSvhyMGxFIMgmFuEurQQlxWtYjos1GF1QF3O1oZMN
vt5EsPLRCPgR1SVtlpQ84t5jTiQRllhKl/LtpoaehRelJ2izaqMOsXWkica5d4f5FOUJlcP4OxWf
BPALNsHBD3sk7bxpSNHcIVgXn8hdVPmV3OmfOfwYsJjMCBEuL7d3aRatXUEYD8rcExPj02tCxSXg
cKPagEKWuJm0DeyIm7A61IbsK1iojhJCPcMaPuPza9+3BCMIBugYzkrKiVI28s6ldAV1lD4GHzBg
EVtdwkGQz4PlousQoJUOZdWq7rxtmdJML4k92xouXHPO9d6jBpeqD+8hKx95w6NnCK7fGP2r+EZ7
09YjObBujeIbKMCrOQIJOLXqRpdz2S5QOuS4RJbndTF/3w+MWTvfuW4QtboQeicAUWLYuFxH1vXf
6ay9H637yqv5UkP+0fXr/HV9XSbBIBEzDjSu34M8Z0Kja4afvUXi1SO/FHs7VTdjv/6JMbcJ3+pL
5U0KP9p7vft2PB+9WsofwvPcb/4hWTmHHZlCuQjXycBTNwrItKbv2FIlxLn6ATrmXAE89rtXt4Hm
xKKURmulpXwBvzz4WS4n2TeLcVRUw9yGHT02s2CFuAeJwy21n1HBE6pn1bF8+aehv1ItrANBKga1
HchmDNk7mC0VcaGt4RGoLkpwOEqK/UaqpKbpyxMyGeMRla3Z8edWrrEX8yCeiAVmc/CVecvPfpjh
g0YH6MJJ5+IYy2POY1kK13T3blLzwp7bjVzEby7crXPq3J7yOTdU725B3XP/S1HooCiZnaMJr+Mz
VZULyuqOlq3E0qnRS1cvwZ/qhZ06zo1Qcn69dhmBHey0XvxqHnH/50y7yDDwsHNZ1/nBri8+ungM
De78cbZe/cf+iGLMzo1FUYY/9sFksTbD4Ku42ctck7kCAPq11QhyxiYliHbmVbBmFvgsv8AWNZP+
bFJ+94+v8qvlTGsZnQnAfhEfY4Ylyqk7p6I3VUQbCu7RjvEqPyGxnkvw0FhdMS9uCCctTOKg/oaZ
t5DNm6QDMBK0qCuNlVzdOTszdhUFWmrr6t/RRjA3mjTE9RxWw4Vk3Nh5196e56XsxuBVa2nM3C8S
6bsyQlvzHmh/9j3KYhCwd64PgdKKjy/nB5xwlFXghB07+YbucOxEq8wOBDflqszCLIHvTUXYj+I+
0GmqBCNEQKUalwjq8dIkY+s5zi1HNpXCFuMIDV/1TwEJDpVFfOC8wKPpGxj2H0LTSmpMRDfPQbUl
xDrajF1ypd4qdKVxMNC3KtS8fd115ePxJvBsYSn/mz9kZCxc5HfP8l2UsvBEw1pyzok5cQ5vj5Hv
bdN8JkLPLx4gyOtLc64Q/LEtWDvVkGGFB07UHutblWvpkq8lzGDMFAPsHxGMEvImRFiYNhVcs8OG
7FA0ISXCtYlhydpyxU6+9F/iu7YFN3thc40Jk4dJknVNZXdB6uTno5EcGsuqt9w0ntZRb2H4o+FD
7dM4AnI8HZ/rdCKcK9eGbSKBDMx4afnI2xeCmHC4TzhaPxRDiHAJLodKRA89bzIz2BWxUnOxR9ri
tjcQrXh4Qlni4mUyL971IruqMUxmSFD+lyN1KrWQsL9HjVQLavbZUJsbimtSNPSdgMsfHeIwbA5/
342arvPPMYn5NTkdYP2KWgCcvEJ5DHtgCL8BD72LLdqNtgaxwCbgGyGp5fslw5vMddbJaSlw7WmA
1L+Fk7y2FjPiOLCqigTvRDQqETiKfCWO0DaUUr2OJ4FY04kg10krRo8NfVRPU3r08w7jotDZrwFa
9fBsVRcaqwoWKuf0Ru/3RU2p+UuAzn0gGwZ0wOBvajPh0r+Ic4YwgZAdxzQg4JJipxnvtc1N+5J0
XGImliFAeOR9BA/QKbe1w+6DtgfW5eJp39y3Y7Jw/fgjksz9VD+OK1mTRItAtHd9NukRGBVvDBpN
FUCCUYNEnKTLmWlgJ0pTnS+FF8Jp7KSZdwFzAxL7u0DU1IsODrrRIujnHFe5wUIet1iWTkoWgmf8
7LBRMUf+zw1UqSjye1s5CG4ayzcDiKop+6IZ857UrJFfVL5fjWb/pryGyxr9K6jCBmu0Na5tP4bM
RDR/1qDMaOwKHRzwpyC7HWWsgcWPce8XYnDOFJQe7kYQpBRjf2/f8jIHdmdDjUjRsvt0MJoDe9Xi
eSHM/dYiEEeEU3G9FlJlDoLo5q9UhFFVSPVpy24jRkQItMizEtL4Nqvm+hOEyEIHpwjGGxppsU4E
hH6H3wemA/xjjG37Gt4B2ijI9BgN0rWP35SFkjrlKRRUyl2VzHTuSqGWBwv2J1BApWlSGFcG6ycS
NBC/jpawKyOiy9o6kLYNT36PCcRRkHRm28VTs4X/2pBHsXDIAOPsR4zVaRiCBlJaCiJDcTS8N0rP
XXfGEqmKjXz/KsMHH+l9rOBKzi8L7uuaWZY07R5KNj5ryKQeSfNeEdqcXZWuMjL4THPpuAUmz35q
POGYLVMvVhtJMcxHf6+GQvyOCj6VNVd5xcMHTPw/tcgiXnWsPzNAVfxviVdotkwCo4/N59ouhXCw
hGVWkOrtqBG2ubvftCo+32WBvkr0ZRnaIZnFLyPvdRivH2KoL8VdaTsK1Qw6CvNJbZ3qr5R+ZedU
SPs98HI9d75na3e8J5mFVFwQf6YdcPr/a3VbcymR+tc0bbmhFrErRNEAYbzPfFAgmcf5OSUYqCZH
D0HKIsV9z0tYZqVjxrJ9EXbRbA/nVZUQwPGlhbzU3Ix2rYbz8A9QNu21IMKoWnLWnj7fX5vP2NuM
gRP1jwZDFlPl5X0KhfQsWFf1gEDb2nyKYQg0TbIMqEkJOb+9JWzsQbToYaSSuszW4WMMJG3IbcAq
htbcM7gicLQbl5665krWokoLsk21SD1lUJi+/Me9nb3VrOJ1m96+Hme6wfphV2AckdJrQFxE4dRX
qiOERy7bUvfLxhKekXYDDpk9AZ2HGI6pjnkg4HyXEFeHi9QAhESEz/TFm06nzOVWCh1CYyxlTZys
vhE9ekOA8MPa3qsEUHky2OkjXnxj+G+cDU/oBf0LiwvVVBkbfJeDbrtITq2WJs0OU+EqvHS9Oi6O
b649pupKPx0y7kYKITOuQCW223jqzjTqnTWBkF4ui+blSjGU027cE8YDOoWBdw0JTIMIwpuB9plL
HmUnt9ZWryyV9sRNBuYpS7GYaeeM8FfDzGAh3j2F98ZCGBNUWdZ62Kq/2hzVV/tIUUKIMyyMu8cs
K2v0iw9ShXD1whkHnxYcNwMK4E2+qdWtp3leDeZEQSm4WEpolfsg0Ety41A8dVOk1dD8H/klF9zg
tNSLzfxvQw0vINef6WpYPQtUkLhcGK65/n4mx0thTMHiMriFqrSAr15f2f+LTorwp+TsxzG4Gejr
eEX9HkKNyStuM9wq2OOItw6C9nhngVIxCCQjaM1qxCawH3iayBlKpZoKw3Yy+tVFOaUDHbtLH3Eb
s5yk3NlfX0miorG5e3BPDouv/xFatJsJUEXOKXjAduZZGE1QOnQBe+AbhHylQKiMKPAJi3hJARAf
DyrAMlGdZUP01g6hpgy7AQU7lHFgTDpOZNjBGxXfif9C4ZLSiAbGCYJ6VVDiZq+LIIesV9Nbr1wy
iD6a6rkLUV4Thsp2htmSfhEo0q/m4UbGmfcJvE2A/sB5hD5LlLX0Rap6sXd4rd3ZwkP5/UF0Bawp
Vlo8cBFTEw8nKyb3MxPeH+6d8ZPZzyOtqsoXgU/nIUG9rOIwzqcKZoAnFv+PETm1EV2ZukiO1/IW
RBhWv23M3XymUwRysQkMaubvziQYapgze+9evvo3O7+/z2PSyq6bnz7iw/OOND2t/EfTdoDjQVsP
w9/E2FZJ8mFAnfqJGJ0HEWUGvWRn6G2AutY6Xg8vUYQpyvxk7aCp7oLrlIAWjGejEm4ZKRRTfdKz
5pfR1Zc6E+C/ZXoblRIlfm0IY+4JMkVSUqMdJVklZoyG21lLBN+eHIxRiAVuHtIXpzsXbU9S1KAD
6V+1YZtiz9H2WQw0a1IBwei5qTMpYC8wJpvMACBbdc9OJMNdVr/2SJWnjDRaX1Cptb54X8j/sZGG
HUQ88MTH6Jo4ljNZ405yz4h+iUQ7zxj+G/VooUCDZfiWRLFI0ARW/FW8wmFEWmJiv3KJOG6hgR+J
tz54bOqmUwwfx9chQUGIfZpPom+GCARr5Pg+M7fOa5XklqgI/rphnCOeg86wTlnJ4xFeMqU7umUH
FdyflEmO73fF7vbI4knyygJuF37zybewisJu6MpkbyFApzYns1AL2/8kro+0LkqyA9Xg0rspLIJy
cxdNCz7qETMDZpZS5+hIdVjRpuND6PWJ6Esnx3cUkumZFdysTaEUMCcBBW7ZZjJD4isHQirG0h9U
gN5n6eAk9N3eyh3doQyAaTPwdcYb/ma5GyhCX8amAkdHNDTRCRBpgEpEgKAWrmhNDH5zr9XNXcIU
lYFgbl814IuUtQNYqKWw2voPMoosCjyFZ1TOMI1gCgOp9emXCPj9lOBKid6l/ct4KJ7lUeBd6Jko
cWQ6lNG05xIJX66r5sNBkiigw4xPcVv7vM5eytjY/nMFK7LU13bx4y9aIOVlGaoTwP66ge6Vif5J
ffCyuRHBr3qiRLqREIb/ksJk3IYkFfepym1L1KQUghED1YDZFkJBa3KWDhbScajQ2KZ4vVwN+zBj
WrxC+8uG3AcSl2DNSeGjcfzvRvTzdlsne/hr1ZpetISYrxTWqF4bYbRZlgLj36ef23qK590KJyGi
GE7YG4U2S//Hhs4f+IeNNGnt0pDRkGeGi9ttsih6q5COCLbbJ79Vv08wd5H5v0AJjVe0nIWDn3I0
Jne+8cKY+7SuT4wFFh6hPfhxV8GyVFmnHuY1HbE3SDkGSVYahJ4TyyTfxUomBUIfJHPgWJO9YMNx
74xGEa9eVx14C+aYSrEj/8WIqANVIgdDVutoilgJYBykGqanWYhvp3tHOEr9v3fJvCT+o6dgctp9
FT+5eiQxnwvkXcf+wOy2ImdHlI9p8BE9D3LlFGrvsQvBkRknE8BkOZWuzTI3mAkvxkJJOpqivib7
Kp7S6Jq3qYpYX+7lLcrYpLOKEsdPZlI/6nIGzfQOUpJ8HW1fPF+Lqsccz68tS59xA3mH6aQ4kLym
8LBvEojwTbYPVMZvtK7GG+ArrnMKB2Py8HmActBvmRVjpeocKr5ZuLXYtrtZ9C32FncoVotqdz0Q
YPfA/PacErvDLcq/hYgE3Gvc3SRnrN7GEkBorNTzxygbuZhR4zYBrLskVXukflqsfEo6CMKKPl2i
eTgbUnAuAMQFNV2Ejq7Ddqa83A0eG93tkV6pcOdOuStq39f4E7c9Su7gmut1uei5eY4FqstSuPhO
smcHXgv4+3JAV6+2wFlovqno6INhbFg6qZViOkjRtKoQdWIwSF1vEJZRQnH/CdaBZojIzjQvWR4q
D0E26zxvwapWWc+bxDKPBzk5u+w8ghkYc22BqZLbFw88wgKT3rkO2iYOBBVTcu+nox259mSqhRNf
2CWbpkRp7Au4Bfz/oFb7khG4g/iAWvfNvuMPRWb3cSL0ANz3idYuzWff2VWidbiB+3SnXeUCXLSM
3ThKb88XWfDxbqRnmNQapkI9xlGHZpgNGVPXcxo7ee9gs/MnEcNhP49pqfWDqG6Wrrc0bus5I7Xs
2PQM5MUJ4GFfhlieyZk1YPmLApc03/TpD/K3QL3DM3w4ORToLr2wfHCJxDpjsJoxfLE2mAbK4HpE
kIJFs+ksJPPut+voL7LNrxxqmmLm3xj2mxCf5lCpe9ehqOLJWerSBg9LSZola+olB54FqBu9pVdn
E1OImLlmJ8QPWindyrwLXDQgFUKKk5P/HOlst5uBt1Tv3l1qQlGin/0mrelUd9LMDSXYHAXoYlcY
nmm9Vt6T71OPLj1e8Srsbcl21mV8UvlnjyN3Bs4d2RsiunOmXt5KlhQdXFzQ2g2HJQZ5xEKPqXmO
VVqKcYZrXYBy8qWLrT7Yx9fRJuOCHTD9YEJTBWgtYwH1+c/RrBEjtGI96Nv5GV3dvlwMI3+OvbCO
5rB88qtYvvMBw9l1VB6JFdsfp6UFMUDng9TAAA8TEM8MjGVhl6SAKKwJJ/a89tZkoxV4ajy7uFXU
CnN4FrAcz7rEUymHt5+Gj7434erh5rud5a5sNCBtmrQNzm3VqHUJGT31zfJjVWFNFA3LbzlY73DK
vl0yvUjWtl1MePH+7J1XD+x6z3R2RxxlIrwKdHjZvm4g5eXf5jHJ1L0wxsg+lBMBHA7BjKpYHe48
8ExSQV1/P6FoIr5XujnlBuOEFPGO4hjjrbEgqT849RhJNhBiM8WNG32at8/vPYlAm72wbs+fNQyT
nIv0fF3emIQyqvSvmCZj50fb+WP7XiHIt6pDerCGRaSeRF7L7+o5LfFjRdHlKv1uptYwhrVkjaXs
AYaENvltbG6RebtyLiIgT/7ZDD0xLGVZehfCMO7hwSd1n9QUcjU442ZQp1X8uAHD5/U7Uj5Zp+pd
Vuzq71ovNO5m7gHnKgwpV5CXZzMQi1lRgLEvkHGK3EZq4EYfE40+liyx/52gnzQM0rxnJqr9p7rz
l8WQ1rw5MK/sOB+Ld2eL4Rov7qJ0sMCzQ4KaaH8vlpcEWbDDFtsLwl71h6iB7zS6evq4NrQQxpp/
rIS83LbBRBXzSTMZ/Ap6sr2mO7Q9xuwrvRi2lOGoiOtMP4jppMkdQyN05BJwL0xWFzeujMxt+T9+
Qn5/QUGnAHoPR8Hs1pfXLvXOtpH+LNfp46dhN8I2zWDPAPCNAApgWHUPNwKxt62U0NRTJmT+2eQn
4XLh/0AugQQ2Sv4joDkbV0rJTctzsCShEt1G4WTygEGhJEP3Pcc6f3WAnKWfEPe+8Zpeb1niSQ9a
v1nGfVNOEuffydIcAuZOOiYr5AbsqJIKg8V7Eydq316jh76lDKJCvuxe/vbtNwdqzBtaX6oPDoAf
y4frd4vLz07dyzhY6gMvuakCzCJKkUj0T4jPf9Zp5X/UkMhUkoiTAmHFKwaURTsIeHSJYKmHed6J
JbJM1lyCVn0rBUxVXP73QEpTCoULejsz1/zsphsERDALLUYB7S1BiwqnXHt8iAveYWSbqCjFFK+A
K2wFC6RawMBB6rB4IZu8H2d1R3pZZStg0bQY4TE9fVT+OPQYBcIiRBrHkLwfFcsnt7MJ43KJ/LrB
4aLlLaCcltzrqd+jPoN2r4GpaKnvCNY3KA4L+pi70EHbSt5W2ZYTj5PnlnAQobir9mpX4cS6+h1u
wa+EwlFEwd8mQWE9UJZQKfex3wcYwSARcgpqb0Y1DLUqBh+XmDHiNG+oFSan6Goy98/50x3aTZCX
mvM7g3LMHHmStDCUgJ/ZCSRNbOtXZhdwfBaDWgvoubfkbWCZu3AgVHf8vNNpSjXUp74G0pc1p1k6
+M/GYkvKueOJxtgvLsxYqLZHoNYRa4yPsZbGmFTtO0M2zmMLEnXgl7OL8osxZ8RSddefKST5kH4A
gd5o6uQHebaBuX4sPLVw2imwTHtMgm+bxxiCImd1C9kXAaX6DoHEKVkMxdduohq5R6NSJfEKvG7a
6dZWzwzhmOhZqFFrIZTYbc3buPDNVLYfAP/thw5aXrZf1ylNz9u9m0VcxpKDE0dTPifLmuyJK6vY
1C5g6p6ctOH40AZCz/leBUwOf8TzXgOJwykWtBailnPAjgcZ2N6YqGczHpPuxL18JI6ePBKpJqu1
r8rEy1IWyctj+Ns1Wpl3oKwlg8RWFxOJvdIR6FV4ISE6SjEd1M2O/Ib8rT8oeKyUI202wvpRyWym
/bcDaoeqDHNQnTp9BER8QAmtIRHxI56HoleFYklsQcFJddJ2DZFwVMx3l8kWXwi/gh+nq0mDkcoe
i1xmSAzcOUbf3rFEFkA/dZAKRei6nuVKs3TLstaPYg9vOHOamCtK4cEFOvZg+TVfbAoeROC8bx5S
CW/p5rF9gr5LPhZq83oovCyjuqcaiPDChxKcj4KctGlH401PaeLXDmv1Fu25X3uIDWV4yd6D+cBL
+wQWO1ofUFzsNJq5jIL/oAZ703/7lQ8RpFpgLMZ/MXprF5PjYJzUtdEn07rXZOS4n8oSJ8uC0nSu
yndiZQHv2HzZDJrKvwBsJE1R/f4P9BHbq4u1V6AF9rGVnyiMYLOigq0xHpwVdOY7PIltW/SRWBqb
ABa9bsq52up+evDPGSd/aZaUYx2jIjzh0H8tNhsPRSLVxQRIt3mtjhRqX1lIGFduDqAUIG5xZ12X
py/LTOix1nsn0ph+oaBVi/8esG87mCL8duDpcAtnXWfpGgicOz73dbqV2gumIiLsF9uMfF78SlEO
xO6DY0Bi4MKMYz8ZSjfiHRlF7KTGa/oyrf3+hw8b0NuH34CvujleuCt9WO0hCyEdyaRNi5+R/Iu0
vApRqCxGKlSH7LlDROxBkF/PN7O8xNvTPuLUfo3h6p4gmZDeIRvCxxwphksGJ4UtcqZPGwKurlwS
gtQaCXoqNcAXHqL3q/ER61/Onc3DyB99MvNCDQvFjtuZMFdHYiZIZ315f5yyIKWTrdyvSBoq5wgI
e/W8uXpM29JYrzqfBhvoZfHlUgDPeE2udJ614PjKlkI5caHbbpP0migTZoiyIOd3zBhZdlJ/0XRj
HcD6uN3E5WqzCaLSAoRGBGxVbtk9+SyA8Z694plnI6fZLN0W8IRXllaGZCkpc6AmOl5jF/tfmvJ/
m1ay4jFtQergBmxmzQ8cAHlD5CRFN38dj9VTygXTpjjUIMenbQkN5RIAOZWh31gmxrZPkN4LRX51
pkxnukD+rW0ECmjo5DBoV0C7eGZ8mTITzURMpk0PmDg2CDuAedgmbMUzQZKTy1Z6J3DcFu9SWnpE
N7oU/JDrxGXIHkbJ3SIAhErvkf93ASoxGTFgeV0AJA9T3U1GclHf5g5I8vr1ghL8EpCDI/VjvBLO
G6q+IZWxR8NhBYnKxj4UK6X2u9zQPCPqvMrX6UGUrNtilOtETQkwoMn1ElobaOviE7xvFqa+CeOT
4usQl2vLtqUyVI6pskiJ+XqNKKUUzDuBE6Ig/jDgSxPh1TFQeAcRiEi8dGxJrJtYSW7aLNHgporO
TeDZXQCnd9+ZfaOoqZNXkmGNydMmLznCYcklAAj+uDa9mXWj2N7ToAzovnud48ZQoZvKXvC6Bzxq
9JTbDuiP7eE45B8nxyNYvph3HGu81xbU33Rf7zzYgTRmm2Y3che8ULoZUhnNj3PzganDLTbhhLWj
vQCCT78xl6QvJM2PHmm5duXUK+TWyAO6cYu8zWYlWzsNc+8NLLwW3gEFAKiRf8sdpdOC5vQ/Xfhs
aLYgH5iXKyr4jfTofu5N0MP7d1v+oZ1H/+zYWaoCN5HEgtzkx+lIo9+1T3Q4DRVba6MHH7znS3iM
cXcv7CpGoadNTIMQhRYtsuzWoa5lNpzGJMzengmjFQSk84uHW+9OBn7Pkd4Nve91LBYAg34XTvaA
5QcJ+hI/HldLLmEycZK3IRdkTShhHRVElhhbqbvq9PosTSgnZq8Cb8RU5JB9nwl4piOKjk/ySFsp
XplxRzApgAGuLHlavM4drcI+ao+70E/GAlObZuSCF9qlMYntV+PBthTeeuRrs/sCKZsH+mPPxBB0
Dnwf4hfDTcspnYfZ7zdAFwW08c28NTfet5c8o07xAHBrFsm/CAwCD2uXd+37XJEdrhJJ2o/YsU5k
Hf93QajanS5TzJVApKdJCVyX/wwOIvYB8oIYW9hbiGPoqfuZaO9CPCCrLo/s5EdPcwWfepQrkien
TETVCpv80hTlJi4T8LbVWq7ZabIA4MSeMPmMcIcLuqS8ehHBJeoFZJjBn1QJ3ObUhKvEqI8G1DHz
orVrdWCd8sRcuqVOrELdSzEN5xzak1kDa//eynoMhn3NfvDohfUN8ckKb3SintAe5hhOnbQLNxws
cWcy4ffS5TqYPUKkT/iI9Z3xVgJHr2RK4jKmTEc6J2li89J/cEE5eUFOwotTsG7nLZCcGO3+xHbF
xscxgEO+qV1IQhi+SO9l84khAWo/UK6R3GKSjhBGwmS2RaSt2CZuHC4hRDPPmCq3eyvE0L2Mcoc2
OjSykH7dKf56PZLGnBtQGdwmXApuDXcJotAWDH1r/r2me2ONlXDsuE3MlFDIJX3hdXKpHorV0LDK
dBqPoSUM0u98f9y0eQM2SQcWYuf0oDAWnnl8LkcVHSCCbjGAv81H3Y8wzjTLEHjOggQjUWvqflm/
yfUCbuUR4JSkPsPSM0+v7kLHpTIvUNiZ1T0a3Dfz1OOTcg7pTQJ2a13xrrCoeKjIrT1DF3JY6gmZ
wZTHwYWOsj8BfV/haedRCx5BgOAALFSAz1mWTt7tLJDt16I6vW6v3guerTUNnzVx9+eMn5H+l1cT
KNiRR9qDj132r/s9Wz+9wpBLf5wXtQMur4jMDCzqRD5Q27SjaVjObI+1b/GuAj2dBKnuQdkwzQEE
J/doVIOrd7KnFGGMaTEkFnQSd1xiSN58pVuVQFiejWajcErVlKIX//jw8t9Laz82gASEZZ1Z9c+m
khdtodFI7f5Z/GiS86S/I7fF8sc83nfY+B/PxV59TVzv7HY1mWzjWq68hZ81j1+bfbOLAIaFSBcr
3VgLk/PEHH7G/6X5i+NFybJ2tMHXSEZ5mctKBfP51+FQgviCLXpw/bM/Ny9tB14OdF8UDx5ZsepF
X33QdopYIWYxC8DU4eX7PUObuesSIw35BURt2AUSKFyRqBFqbWn0uzsxD3S5QUvtaMDa8FpQVu9V
Ose5JiTzHrd2SC2pxaoK3BMmNCVUm+fWnir/xlAa2iwGWJeoPG12lrd4jHnuuWFLgZXX5oOFAMWg
luTaEeNhe0cyqKSF9aRkgN3nb282sBMMpgrfEQPSOsaaKfUYU6KRDEo+tvcvO+n0u921JJSfkmfk
Mm90jEGXeSJBavLDaapuwE5ogiss9w2cMRor9GY63oIR+YjzAZbci9IWDDmAAPA6p8pr3bNKLR9G
tkbVkuOxqPer7bDpmklZd+K3uFuER7tk1pPm5ddHDEm6Ya1Ork3H/sp2Q0XTFns5TYQT+6id0Cnf
2arKTP2v8i8nH/o/SjEn4I+dCE8+8JRpQ+aNX3I7LjwECGzggXUWIwOYpQgi/Vd9yAL5gzOCT6Vs
sC4BaPB7aGXgl9FosbMRksE0h14Nil8O1UXsdGKOx22x6GCYmKSorIsLBIQzliHycVyNIGod+ddg
sMrHirKvg1mn+VA9gy9Mn0fkkzd0ptV8+OeqrhWxkTFcanlgtw1M6iRjcaRHD8fr/IzEUAyb3VbT
jKK5/QyoVl3zc888vGK1BFkAATNcLiVSepOyVHMl0R8uh5Oh9MlM7B1H3A5OXHOIFARNPNsA8q6D
Mw+EKPczn4BZpgZt5B5xJmKQfDqn8yx2jTtPnz4+vLWMGr6DVQK2FVPOCuRwVL9o3ovzLtADCP1H
RcnrmNU13/++qbjEoIgA+DsXnJgtpF9SJJ4+2NECKjY4caL71tvgRtWmLO7qNJkplRO26+Hdu0rM
Q6QhgWMwNmM/DWTkW0PiEuEGGze9PW5PZPqt50BarQ0gyowlshuInGW52rleAS8J14NaUsqoF309
qi1fvn5VXayuhQfvgYPs/ZSfyPABWSzgn+6lnLvRgIG/9oJSDAzdNRWjK6RnAHi8MgneBTv7BYkn
fwCdymAdKDzWoPb8i7T5SSA0TbLt0FhJ9eR6BnzdKaF0/uTiryL298NMbJJo1sipPIfSCIvfKsEy
xoDJFce/4NxGAIv0pDX9Jiir+UiRGi5NAaZS7J/+zpSfv1ncC7cO6uNjBVtyNpC0fO018oJmPtua
P5oNbHdN4x8wi8nYlWU+7xRsyjPEeb7xu4PtE7Gv8VnDo1UOLaIGeMz8ZkDW6f/RaKgC8a2mJ+SP
sdeZM8yzbt1Dv8v1rsQmBzaScS6ZY0tjerEVC5ADxhAuK7kakTEcVYtrR1yPcQioB7SGZow0tGut
vtRc8FfxImObk9SvnzIDAbnrPYfvAH8HzjfY9Xpfch4Pvu9+UHURw9BGOCCIGdhPVAfDEgSz+RmV
EabyRXG5kLfFXfTXRfLUMxrB+yIrY4ZH9KsH5YtTS/DIS6VcAwtFS5IoUDijwpYocM+o00QTLEk2
ECcCLl0qKSnpAjqynFkMIwtf7qmgxmLngDZeopTi1kTk5hbakXtYaR+S72rorqHcYEruyuccy7CY
syeuq/KvZ0aO4SNY+ryimefxeDZbDxVevhFBKP9O/wkm7fGV/mF4iLeK0R3ZqoQwMJ6Cpi1UWYE1
Ad9C0VUSCt9l15AnQRTahbgWZJHl6QwMV200ooZp9ubM9RPa2Q16yYqi+5WdhKmnZUG5buQQkVpz
++9gPKmAj4qxgUCH9ICpy6ejtPDWsK+acCbSym+zpyqXwUzrSLc3YrgiPssDsJ5lk7PINNznL8/6
Q3Sps2AxDUH/knv5MKWIzH3ICTNWRR2WcnfPFEt3C/Z0/FlC3PTNsx59GO1JUQ5NXE6u1Hg5EzGI
Og1n/1jzoEp+g/4H06wPXaQJHEZQXGD323QM4sx8bxoQks7wBi9ngsWCi6IE27hGFfL+nuc/yMz+
UpGu9PNfvETg/P9zL1VjdCnQhpl7Q8myGjqTigD0qodko3gRFZ+52OJrcXsFU50KWUwXJMb2orkw
X1mk13oVboJRxTezkMZ1MgEKneJOLJSO6otgNupuIYD8ECJHv1GUt5jtK4EU3nwWsd9JjkAcF7oq
g6vd/9JS1X5NoOlCPHNU/AU02zM7vEtLLwdyqqBcemttTRWkUzBG78cVkMt8JMeKapVUkMotCfAd
Sz+M5Q/lVkrD5lSGaRcROF7NLhtXiGh6qwJMxGkEAFK5OAi3vSzmAkLYMH0OKzTzp75VIDheOnUQ
L0SJr8/++K0hO6IdmdSwCrMhfEFtZEbfdvIZhaBBTh1nd33V2xplUtfVVtEbY/2fIXh0DoWdIqJZ
gBt0qF7yOovMqSGRWlCGaz05BVcIwaym+1+umUzFirIBk6bEvmh/VZNfvKn9cWwmm7TDbS/bDAO5
Db23ENfU1jqwsGxCA8pg3kgr0rAVzD91sGkf52Ze9mlEKLjFb6qSihCfIAGf24WS7wPxnjgkFZ9N
qHVOGG3894SbgfUyk6jSeAcTeJq2ZgOIyuYU8x4okFPtbpzNPAmsZLhoCCPWDOj/P7zVeV+nWa5/
69nah2VAYaqBCLysN+EeZX/YjkfCqsPkowDjJCAEAzsGw8AlP5UUREDp56u4GOwZP2UMWXSNPpq+
HjfXtY1C9HTP9WB2p5bCVz0Tc2/a8mIOzG5DGpGgxSzzB7qUYNQDcqD7Gogpv3o41vSfgpnY13As
HWjBiuCX89RbCl1Xsw9Xt8KN10+1YVYRNPOXRzi1EIxQbMsNs4ZNixqHZRcaxWDNxwjehQiEH7ki
hLy+199sxZ+2IO9PKVQglWYxo2jo1AieqrVMWRMGdxWkSAVDL0vnPt8ULN1gCi3fKR4NQc7GJ7Lr
Ipqe1h9wjekw9zpXsJhPLhxfHOl9QnBO3coCipdDTtC8Ao+iG5LMWvEB/HQgoT23OZG1+SnGG2+J
i4/1d3cucylAt6zozAipwAR20HIBuTVViMJXSmsBkSOsLqW1qrA3ZpmGKAd/JSIfujzBBn/Z02Ct
4La+ziqvonolEVojSkimsaH4DQj/1Fd4D+piRIXgQ+AfkpNFGevGcBqtaQ1Y5m4Qe6728+XMHzqY
+s+Bp2IRaerpeJrmE8IdDm1XT3jD34hRKrmXdqXErgFzo5YLFhgvGTd6ueNVhApN+jWV356OWHpy
JG9rIPe81tit+ICqFF3fR4TDU4N4TCMLzvjcK36Gz3flxEqvYjAYhv6lXAQEzopiyNibCrT6WlU5
eEjNx2WykaAbTbbR1hPkTTSPpeq8JStdXQfem61bybQguYYUuuNpioqyL6+/DDAn59cew3++yPyZ
YIYJmsEJYUKh0jj2EnotMjz0nDs9695woz5id+oCc7iMnrX3sUoneM6ec1zE3pbfiCNh9Lo9QbIo
7w7JlJz0PmUgFUsjVUImi2oE5lT/NJQj7LdVsaJuY1O+1WuqB3K/MrwU2JSLz5YBydLoEtQZoqY9
1tmdWj09ZaPyQ0MSzbbDy0qQD+Dhxm0xn1SseI4/YNeXSEe0VwziNu7W9WW93g4HpVa1s6a41uid
LEU7ZMIDy6fiwSVHEWKRHnfdLxPrq4drw3YGEUhNI9Z2SSA2Q1ygH2WRnf3RpzKZbDZ90L8UMtMe
0KSx8cljGuPsuyLu3RgehpjY8FiU3JE3zhDjqQkNa8pARXzj0PEqpVtnpPcgNQ3TS9L0G0JPbcB3
6NpDytivHDo8VVODAJpBJaShp1ErJ7fJ63mu9/LbE7ctdBay57DFx443RGoBnWn0HUzm6KBALL33
VcaZeDoyOwndeyj2E/9V71B+u3ZB5uup8lHNyq2AP8pgtizZYHawaNb2YEH9am1iokEMDr/MQfum
0iLSLhvseY/m/IjznYr2BSJlMV3GA60m1ZIJy+tX93JMwfAmWPQrQ4Pf8F//9zBjdGtb42NJmvgJ
uxv6E/U6BR1mYRSHpA7x0F/VqV1LWtvFQfsSvK3q31CEeC6pEz+GNkAgNtH9sYbAVGOPhoRiCm1L
WCFV5wHkFzZ2uZjCr59Wo16nVd33NiKY9ZvkXqG/qtVFprivIzpcn2MrETwxWDL91jBXh+s4hkVf
AOB0mwZoXcnJki8RqDOduoXxq9+xIX5i+i7+Rpyo6WuI4r86GR14uQ5L8TSUK96pb4NsrxM/GJB0
m3q+FUviOvrwTf339ge6ly5AcQaxTu1hAps/uKSmD13vJUJ/1+EFXikIIPsd9lGjmjQIGJ0aiP/G
75B1UK1cWcixABhc/f3TRk70ElOPrXm3aaN5bfLnd9SteLRSr0UZ3lGBC4QgV85EW3SGM+r2Q/oE
KVDVIVfFjwFxr4iLxEiq4RxD8KWV6q68l8lPSibCm2AClJvIqXWxRUoOpljWSr3tPSwKcpAHISjU
3A4ZpWuUApuwu7OcsGEGXon/jZ/EWD4Spy1y41fv4nPEKr8vt3he579WNSGh5gyNmuz1Gxp8XYEO
DV+7GGxNp/K3Lp39acpoy7rBxIAQt3GfPAh2qAMPGtkjG+htDAb3Cwymgvi524dRGYhXFMdr7ql1
nAi4h1yd75GJy1zUmCnU7mVPxW6mtV2m3m7v0OCGK07Q3frNFSyzagM2gefgX4NcxftD0L2gH4ih
bMwT79b6AyOtEjFMytcD58eqVSuGBmVwNSjbwEbZciIKf6UeEui+qbXm/vElN1Ttnd79YZZ2WQI4
jUppqGUbsxbDQ9SvHp5B7/K5jMTNz+k6mhCxxLUDmKJVc65bPVdKo1ikdZcBRh5NM5WSVDdHvOXY
PphoOT0Os+5x8qz1pn21KNkwcRatRIz52cuwX626hdWSc77IkVXeY4W8FqGeOLT5HtififAXwo/f
rjnoicaG0bT7Pbi+zkY6wxW/Op1M3hEhlCSbinID3s4oqeyKRe822UKXexkVtygHMpUk/phb3hIB
jo/qhGxibfBrL8X8Fe4MtqCPSW7UP9dMlBu8ABTp23J2DQ62Ie4Zmkeat5KmPPUv95L2Qp4fNktj
gcAK0ubFkdXR63B6t/xKIl+3LoZWghETb7dICxsopchYplLltdnoa1Nzg8vQ500OCjyVIAVvTXBa
LYQS4laFvdQcgzRW8e0a9SIL8MmpJIzzgqqXSXcjQl4aZq6HqWFybX+6XcTDGqhN/cKS20TuaeG1
mUdqUJA60uuD2tn4n4bO9cxM7uqYKp7YvpwvoxI7Lx43pgTFYkGlugQhUVldyh3RPOKgKzpz5OXy
Mo+OEcORbwUdVMHJoqNUc9s5Ai3wFxYeBjOrUOzyGqptKAR1hQtPEXh15jbHqK0W11ka6h2c6pkf
3g5r/Yg20gicuBsf3v4z0pB9oAngwLEBpEUtsg0MTJPJzMpAyR236kY7hZ5cadTYhJ0OoHefGd5P
2dUupuMGq7DtHrqdf4YOpVpBHZGF50A3KPlqcc88NZYI0n753nLrRP+cMaKGFRNnbtf5Ghg1eEIj
29eYfzyqsblMKrzbJAwmHB/GKVs3PFSEtGErpgRtf1Vg+TNyatNRBRkOM6Fj736BNtNFO9YSpdkB
gk/itScMP2lABhQNRXEd2tzYaMyF6idAUXktzfZf6fKG1zTHPhyjjX6FHnUnq4BfKXKknVCO6ppd
8Un634sZHET3nQc+eIiGx0KqSSfHX4A4sPBStoQlTaC4bjJ4eF287swYK7JsP1wuXnk8XYBBqJQp
rlfsfFirRB7MjdMvWlz95X6p0G/VLUD9rifObLzd/PCDhlRlfIXOoZ+h/43C5lYdO/ooIACpnzwT
QIxuj3TDVLyTyVs127vPUu7giqid9EMrqXxdhkEGZJPlBZMYznTZmOoHEWq/y3DLhVZR1ftwDsm1
5L7zX2X4pkRCH3ylWewl6RKz/aNlGuNEdciHOs93b0GEPjsRBmYiyf42Zc7Y2TT/Lb0Ubnui9xpg
QC4Ms1cM8B9K1A6OIp0dBygRvFB4hZ+pJBI36C+LYXFIIjuk1RaDDsuCNTZi6DblN+N/cD9oJW9t
BC6RvFVagNQGtXANXN16fn5m5omtxjcKFQE3en0QtUeXldcCIMTwuwq5YD0a3ooAybs/3HM6Pp2w
tmo0u9n/hkO94Q9TbmhIbjdHtD3BnUqxcRLMS3+GmtbJtNiS+Nxlewy3e2Qd1gvIgC2/K9safU4X
jirX8VHkJxLZzxQuvi8947UqRl05hBX8sF7fj0HQ1KscokcbZJ0OZJLkPc7jRwrY8N4GwrMsZB2Q
LqPDb+Xaqbq4UDd01s1QabeMn6TtTgkGfl0Pe+MZOc8a5WAhGITgCtbzelzcIFut8iKfGh7BhR7p
RAPwXnZUWQEYiTGLTIPKFyaIkjYIipeSFoxu9JctEP0sIPcnQAq/dEQMR1Rh/12CtJNZe5h9KBQ1
SSlkZJNGVuM52IVi5982aCG9ss0p9e19F4ZImkjM+4co1x13QfxEDP4lRJgxtVf/glJ6yHSW4Vg+
/2qHaPNE1xxX0PSW1sZIv2xOM2DTe1qi3Yw1Z/iQQ7+kEwHCzyspHjTLw5m/jxverCGQQGH5ROg6
F+e5XSM7Wglntu2V2W3Kx0Pxcb8K+dNUMdl2UUMgbB2sewbLxnFMM9XjGiddnjpdD58M6jolMeH6
vB1Zo6g/eZPGbC8yXuFRXzgbKEyXAEWauW/v3V2Q7e7cNPX7Dig3GwUCgzXCsQsz/i4HVJZ359P5
KGDiSh9KuOfxYinhUmx8lIEIV7JOZa/3sA+lkFF6b5/NV5usDT6kYAFwL3SXmVmkY78tvTgovSgR
OcO5Gc0sJTKlEi6RJT8FlreCgAlkA3xSYDdlWeAYqLL1/Oqn8VkBMxI7a+5dH64UAx6ZWX/JuKlD
uZpVsc+0DGPs+h+RBeMnNje9MzEC/2oL9k+EB4kEoCODDBsuBdvak8oSFx8PyG2qGXIe6u+yFYmq
yil+bIhNvdwxORZKB1dfCf7lfnofg1vyLJHTleXhRy1dIZY1RrHV4uF30c03aBuFlVben18eD56K
mOS1J/3IkvJSCYqJaghZHpDaH3mtOMxwpbJjD7vT7nYMsDD4SEBNuNxZ7ejZihAJvdQsq6le4Gqy
f308voMqUZjaYV7od8mNG3fDQnYDA756/uE68f6KDnIMcTTmla20fSpce8end1w6HWfQQPrhFAux
naxw5L9xPqyMMjEsQNhF9TQe8VEOkfojj/7rah/DXDbDGmA8cZK43tzQUDR3K3mFuIPGvbrbkHVq
pj7zWTiGJbZ+X2Z7YQHD30Ho5oLO7WHdH1eL2MWMAt7XKJg6opMjGJtSGeOurgLak63u6iBmL/Tr
HuB6snDNH3a7nv18YhlRXM5sLrbFsJmZfsQ/CJ4flQJ/1Rt7dE4IPTEchlFV59Ow10LW2Zv4qtK1
rBFnJWwhhyD5dkNr2WSaDsi+951AeD7K4PBslJrG7YhIQMebgcJp31WHJHQ/v1h7RI2lwZJlOtPy
dEvBGlbOkv90pknszKx6Uu8O4v+cN8h7SYjwrF2hJsoMCe0ptD0zMlBmB6ZFE+i6GVK84Q/p48h2
PkX/QsSH3vkraUS/EZgM30o7fJK6nJHoVRjNa8lccB10pL3PLTsf29APs/cuVMRV2CGEpaxZD983
hEU8RYhi/E9I8I3Tsv2WTkx8EGkwAC/ef3qFq6lp8y94GrHJycjeGmsxok5tWyBa7ls+L00BPKT2
/Tzrz0b9B8tuYa6jQ00iLDdDHbCT5Z0Iw1OBU4rqSJNW07ZOv2aCvM/vbTmbIt9IdKcSb+wCjBO3
Wg7ZCvrZT+NgG5d7OsueB7VrP3XAyxEcgPVirHob8a2A4gM7wUKf2g7Wh9psNQDiq8F1NKxSYxp/
alyAYzbw/t15LyRKmBsmV9mm1QzDj/Mms//fzHXGKPsEsAohw3sgBDvX4TeU0//Fblg9q+J7KPM2
3LhWCDirCfbW/qh9eE1q1etUDx7Ba+e9WtMcFYrMsHWAbrt5CCC199nwiTT2g1LBUtS28T1YpGgT
50Vx8MjCfqBqfBPl60SqYyf6aC2H3+nxMq4Jy7pSeAad1bTek9YUAHf+wi3GtQZqkV9uUZaxc/Jt
8sZAlzSnRTgZgbd0cgC3jeRQdoIj239Alz75U+eAGn78fTxgamBC8OM7wi2ovFa39uj6goaOBmoO
Hk2pVo6cCNTXZ6MtIKyfLOXww4aoCvrdtRnNPxL/vc9j3jwrcnI9AHK831TK/X/rDNnp+77uZtR1
itIZVAeWmOAGAJnOVr0gsDNaybvqliMbIDmz8OrwdUgW+9SGY9epTPC/gonvtWeQqHlTEsQmnuRY
HwkjoPfWwI6phX7XTONrbn02021ERVOt2EYvUwl+Zw5QsamI41Toc12IaxYYfcJnJCUe+fbxWSw7
tHs+ZHTLx50oCGvaNSoHCuYF33mYMUlC7KxOV6xy2Cq3eafTkhUhq4It9fQ47XWo+pWW2+GZboz0
rA2Xc/DFczKSNid3XWb72f5x3fC2j/L3vYkQI+EqaBCPHvYJFhP7iZhXYdBdwptaFs/pnuyc0MYk
BQJFaBHaROHGIAxTXxHg0NTD3nm10C+sVX2GeTfdPQ0QgkeZ6kAIdiiLHop0+xB4xbIrtNkybpd5
RwRkWehFo/v1XooDpPkQegFUJBOXilxJZxYfGnebXS1+d/CO8ASCjRu+kpCPyx+dPw54LXZke5HL
3DGGeNToGmkg3znIaWddk69MO13qMdcVhMTNKTi5MAXFCbXuUoYCJ0z4imuo75ojifP4Y6qX/zjd
gw1aEF+XKmd7QBAZtcF7jKUPWtV98PDeYZLp+7QWqMXrJmD/Tid6r+nhjc8J9bOpQx9O9gZ3fVVx
lj18YuuXdy16VFeA1TUJtYLAhef+nGsT4IrQrZsJfJ0hrf7v1NBqfA534ZTTZx60v+GQkgPFuW3U
ywzDteHJxQFeYYtYscftRIxov/NLscCparnziI7GGClLWAEMO94+KqhlhTOc0T86QTTwfZYousLf
Zv9fALg75NY/JTxZctitEV8xKc3/kIqu2s0L2saMoXP8a2aK3dP+nk9zDsRwR28KwObWR2D5asO2
xO8GN7SN54X19pg1N7XzOqIpPL+HCL9dzDvJwxFTV1MD9ioxWdr/WtoocernrfXcboNZOStkve6g
1t9QDAaXfso8F7M1smfZe6o5AyV6rx89B8Ex0H45SsC7LYsvPkVkPlWMbNgxaJJ0NClh7GdN8ODb
033FQypCQbH6B7Hj7RUwy8WsfiAcaT7bH1dWeaRWSJ/C5HXeD6MVHh5npK1gaZtD0Er+utNqoImT
XMw15ByWxRUiIUzhG92zukXktx2Y1EpFOgUYey9ITBiD/uwJ3kmD5dLoG/m/FUF8pi/nPjCaO8ke
Qs6oFzQ9xFnjDUTS6I6KdT0y9E3HKmJKBZDL5CazIjbgyucMezKoh+avjj3gskpeWjFj2ZY7W/zJ
OWT64N2gRSI1L59PzYyRGk2cOecvaB0BUaulngpeQcNJ2t/+jQOdgXADDSDlyk7sWrGniDTKuokj
TMOKnWlAbEQyXspTMDBizR8IZgX6a4tk7V4qcXI7h0fPFZre5kMpxxmlUurfr0TG+z2/SUkDV8b1
Mk2Irdd7UtKkiznd4mXPOLm+RbpZgqLC2faILO0KgD65KFUknTI39sGYveJaf3X77ddCL+djeMhN
yG5xMhHrceZuxuk6YIrZnrgqgE4W06fBeJGQ8fhEq5WXldsmA2Ny69rkINhMsrKVHdeJd1IokaEd
PW4g6bGFDeZLN0WqqafPqarUddJnXdTzeBMeu1VBSW3d7vRYmwF/D5x2CR4ubru50XVgfZA4tO49
Nwy9M0GY3k5KmZ6EE1cSwphCfagwXw1xnt9GJYNHroFf9AE6kjqOU1HsnE4MCd+7MdV6BKtpC5+N
xyEPsorDyI+SnmjHd31KYdy7c1z8QdWzDxR+mSgh0rHYNtTIB6Kf+mp7KZpURNANcQ/K47hONbFU
EC4KHnSDfFkV5uKA3ORgP4QdtraXHbnI8YGTfanF7sm4VrOqGjv7/iJa9kcsEx0FpsaCVxjNekuQ
tzbj94VARoJNDdg+SmgkfpSmlK4fMY+kWlR0Rf5I/qOgl2hYOGblfDNvu0V+GyROtW2j2TR6Rdc+
mWczDucL6LzhJvK2iS9EEUoCFTHyO3YaipCnmMnmmL0wf9kv24uUgLHzxtyeE7AfVnP/fd+mrg4N
1wpx19033PyMd45vtphyx5mEBbUyasiAVTukQxJ+LHfMi2xMz3IC9eDHhpIGPEwXsxxIb79Kjz4C
GFFt1X/H8LrNwqskHTs7oNTKiZaZdb1/R6r8MYq3Bx8IADebZOJalDu04CUtPV8k2oskZeeyWpwv
PBL0TqQA8iW2IOJZIa07lL7bMV6qeugEyL7tW89xP9OZ/F+bI+zuCbn4bL/DRJ5xGMO1lT6lBwpJ
s4FCP6mYWQGeB0uBkwv1rgF7hYSQV5/IzZwZ1MMXGlmtRvybvpFk2UadlnUYJphL0N0DBnS5o5Br
WISTTTFVmaSdBiC13ddQf+Ymr63yDOm6PECic3YYGAwjOMyw+FgVfppDBM589xJ6/ykspFFDZbcF
1sug+wsfrWaY453im7MYr4Y+xVUngMaGsfT0yJCeyOjN+4rQt9kh7EP1819A51EInKrECMxljYiy
GRR3heQsPEMVCTPb5VyO3Fd5svObt2PjKvGSP+cllF88O9O0VzlukThuX9BtmtQWjWTeeEtF3Fo/
SCVrgHvZCGtNCw9BHp59sWZd/AXqhr0UxfgqW16vPs+wEadX17FK38Ta2kO6Ex5ghrH2HdCtEV43
w3LJe7yRvttxbFLWTFmy6LoDxvFRkvV8AvP28QJUOOSnDqTTe9k1Dm6+p1SQXCuhWxx/k/CaKyZc
TCLy50oDaTsf1eDN6SbodQv/7XR2Dzm8bjqKS9B59R4YAlQvibG25K5BehpM8c3XvPzDwfdECtmB
567e/RWBtNN4/qTJyVppuKYgZT5y1589ZywovQCY4WjaQaF6/SWJxGZWLeioYiyh/lWKQO0UeRwE
ZIe2WxvuoE5LuPF72luB+TL1vfD94xvaCygRDvUIMFIaVX5SjO71473qlLdH5DBy1SGlEkxdsSZG
98TVh77FkLmCJLe2l0Kcc0Z09HM50OFBrTg0F1HalCptS+U34XIfMlaSpbQsedO15qlqtD6Cz8ZR
L3CfAmIKZPWDId0Y25cDTONMde0Hn6ypdjLLUA8aL4ETL6uE1rySsish1M5MpxFUmaFovE8O3f25
v7BxFudMoTEewxMh6egwo+2603X8LlbwI5qUgmKoYTbemoIdFfXdr2Wwr9CQKTeE491Ea+0167SF
pGFxFH/yXqxVCjAg/xhHEEQd+xuLx0aI62f7JVwVbMKmo8BCKNkbR5piwivH5XuIBZfMpe8OpSuA
L56a4XwJMa/Pxkj73r60juVuiW5kLleDlc9EFiaZl1xQRNdX7H6m5tKw2FHpk2jSlw9wGj9DOhMk
ag3X4K8fpsIIqUOKbYyE/qDvCo5eOUq5JOt9V0a0YxaWtiEZkWMjzuBZA0I42YOULdalGJbPSUxr
m8rl07Rs+bEhrTxIW9dqdoAcazehAqjXXa9FW/0YdLgVxW5w7qBVB55PPMDT3dF0y0kcG+S6lFNV
rEzofRxqmiH3v8PDDccDO20ZUMX4uOi9JB0D+xgN2RmwK0GjX4BEB8PLXIRkkEfbBdNdMqUngrMZ
kkRBNwhBly1FJL233zkM+EB6AB6NNCTlilgO2bPCAmxu6M5EPYP1+b9CIOetM9KTL4G9qz9lWpVj
ebbSokfXB7Io/ZpP9xzgSsU6KfqMKmE28YkjdGG3Ln0mnOY3ODj5FyRsgxct6T0ra4yosb0EJOWJ
LyXvZZzgtYFfSzCYDQl36pkkoHc8sDkO0xdUqE49rPVPtj4ybUsN788DiUUXqcjPRYSjYnzjKbS6
lKxcdOc9RiRMqhwKuUM4jXDyZh3l87WDYz5si3N4KIbiQSn1cRcD9M/y0N/IOE7RDOE+h+gZt2Rb
iAB8rA8d6JJutTh9ZTfcxPwmAq1aK1VuluNO/NWwHxGKdGlssWNgMc1iYbE4GTK7ZforK/Aot671
1TinhQ+4Awi9xWcIf0ms++HBK5Qh5f5HwXG+I9+EuzIO0jEFGBPB44SUqPvULtS6o1wEM2CRkW3Q
WBkSFP2EzRwt7ui18e92CsvSTvI/rysQ1VhieWnI5MGqaTHPHGno3YymuNEEE8lOBiC/BHNnkqbd
pFB26ITIBpXfrMiJPSl95KRvGDuJHp8B1qjQlt/gvMAXf4hq8pZKLTD2FsjX3Os6vHuiI1UH6Ktt
dp/uIwH+ZLzyID9KxZC2q7Jx5R8Zt3/AuKYuDBrV1uNDD7JXC7LAG/+FBRDl5e7dN6/LGFj/C4J5
rYgq0P7jGHKXm4A9ufttODVkNoWLLYXGl0+6V/Wr5GjV7tN1ga/pwjEWZUgcTBdT/ZLVAsB2/ttZ
w+hMuOnIFcu7n7AJz7IudYGh226qSOFY1ZoCunm34arKAXRkcZ8BjcQcUwQ4z55h1/sd6lqu0d/s
vvWF2Vcjdd+a7IrvuT7S4vNopj9YmLyBFPeBrswKu2iY71zvreOUkmm48Fp8nF1fdjTi1PDK8d92
WCeRPV5rywQ96nIwYxwMeI222sHQI0brVGDuhDwsNIDD7HPT8wskpg+GwQPRKghi6aTbKkIkU+Qq
2gLC4N80AQ6CGJsHBeHHVNRRNR6rU4CrGl2pQQ961HNNj+dBjjpQg9AOVyytveEJw6TUN4tf6JCk
IVPCzNJIzAU6tiEUMXwu/pKpOZFmxkx7FhAGbNhAvdh4eKU3HFjnZhvAcDCrvAMkEJaU8y/1dI31
DUoZ1o5lBfmM50Cx/t5YJXoTDR6YI1CQ3xgDlIO4r8yehfdWL1GMQBYFwBsAPA/VvxDN0EVP5fSE
UqsZZqwAbhbHjdz/KqpKzgzb7qg+HH0h3Rn1a6WqUx8rgPQE+Ij4FWWoX6BMG6NgnTN5Y3RT6++W
XWvoJOI/L+wE2ZXos2w28HkIfcodSkAlc0Iy4N9DBGmvrnMAySH3O9pw3bH+qBhNLnWy5135a2q8
n09BKjXSwy7DVv7h/OvY3kkbMrDH7vMZjh8E2HQTffcl/SHlMMgmlG9QHu1JJsfbIuV96ga9MCNF
0EtA97cfV67rWVMIAiqaJUWsXYwXcFQZ7uxycwntGVs6IHINvsQZidX59zIOKzYF1f2Y1+E7YvBJ
mH9iitAv4O4HWBA7OHn32EkgQyM36mlAYYgRb2dhoCWY9XnBxt/bbdGQ8FH4ImNycCWADILn9pKl
vg0zIqGoed2WzLrO7wIZ23+bfeq4GYPq+ZUJb6z4kDNGsgEjtY4nb0MSMs8UYobJbR3R4JSHOmvn
vyakg2tjBjZBbe0ZswzPRybWMyWXtLiksVZVtPWOMkX5ZH9oWsc44EiU2E1SAQ6Q/yWdr+OIkqpp
J5CelErpzeHdEPj6P9vTka7qDjez1RBbRqOvcWXxMvOp5UQ2qVD/gOgqNzBbf5JGZWQwOJN2p6N7
9qv6grRu4vOKh0WGEJUmy2ZRNb30VnAw/WX0qNaFb3kAxhEVt/Ta8JmRcg7Gqf+m/w8K9zChWrUO
4HfMNJFVugEAMSLc3p+bwdG/lYqoMKXoEVBBRtpQbIzbTsyAQru86G3HnTXVXt4hDjCvAzN8dOD7
0UbZwV4nj7zJ8tCUl4CzucbyLTj30i3XGqtDO9w1iGAiBr/FhHYRvJ+NrHLUi2y+spdz150DC8LO
hFBvwmHMstOw9nwzSnwgPpV3gpHOlevf8akX13NkybxGCeCd5IK9seT4LKo4xWTKnwrSDGXOSm3r
qN68ujLpG/hmJ7sphdBThNhDSzsqpanOtstxsaVPy4VfD8OfvvcuSwv9IFIm4Ph7EZno9V3HED2g
2rCqbw1FCiTPl9JL/c3czeSBlk8Z6lUdtivZKIQJoiLVg+Jxph08/PWHXDt+r+ych8V63/8lB1a9
nwoJqtnGerbitO0uvf8CoeLJM93I9/FHDuT2bXOMET7sDkOGqKVaBZR8m+WEfainja5sg+uw5FAz
8LUtJoiSC7Iohc64TIWB62Zj3AD+kHFDUh975CiYa8N/OX8zaXhJSspwIoNA4uZF27+dtkL5qVBQ
+3lC1gBas6kjtIlezCmpFAvLHaruN0M4OOk0/P9Jn5FMuhx6QrbEWAhO3VZ/HT2yvLL8W393kYUX
XN3TLIA34NgygpCWS9uV4gbzbwJfrzZtmal9Ikk89POZ+NabGQwttewUCj9gqMWRkdHlKWtc82Nz
iYY4edt5DSgsaep47xig46ez4zb6XtCoYwmXUY6bkdJnTII93VETPFnfPDsU2q/KzLReDx3ABcJm
fzZ+iafb4q3ah6vO5gz1HDEqJ9t2oMOVGjV4yi/aRb9I/KFo0JcKgAsSSBzdPqKHtXhjvhawhGWc
LMC9LRvMKJOD1Avah1f+74YEmD0e8Nl32GH0zDPXZbsbSFXb6XhLOJsRCEkbA5ZND6NoZ4RWDGZT
SORnjHcBrRwLYdACOuVN56e/sh8rnK7szaSdwhX8PTXEoqt5pZ1uc/tQQS03TXmRBC8o7jip3Uj6
IaI984kUnOlA0NGiaHp118qdZLhr79jWHvbBmdH9UW4jl8rPMQFY6wV+ef4h21adYlqyEgS5uUdF
U/Oj9Xy+votetxzGvOTrl42nTuMz9iuBepTjLpz8DCKVII552etshADZsH26CuBeYpkR/Qf5BS+x
j13n+MIb4F/7s/R+DMUFD4p5ffzzRko19vata6WWq5KBbMhHO9AwKI4g68f+dyvROSt8QdCw7+Gg
rFEt/AffcrPML2erqfC2aGYUSUnkMb3SjO6jb/WqTE5QkBVZf0chhjtqMEpUEVcC/TmQ8TYSPple
aOwIrBBmXqxAO2eGl6gaRvaGk7WO9sS7cFatu/OYPGpGoT/JPAXFEa/T67y2IEhVORHoF7idd7ZA
OL2bo1/OQw5IDrkFX8iDsZsXWkc6qktwsy/NwkudOlfvfpp0Xy89FailGOWcuFJmkXl8kttny5Jb
qApXOmCZAtG0bR8paaBPAKYQXcRkhYL3nU6URpreWntHPu/3g4ezc8x8AAtK7UYIysFirBqj2Eup
hzYLpmLBNivjapoKiJtw+8UxnJQeyXkitdrz26BcsJ2D1BlSqr0TcMDuz2Yxljvv2TenL9wd29+O
tBCdVC+isavSw7PY7kOorI4wVIUS9g2lKGi57emfRunh3oMd8Mi+lSTJ0XW6z8OC+LGCY36gddQG
dFQiZ4SVTT3QjOgRZMkrDVfyz9xStTZVfsUc8LHNHNHGplIS9LcXMBNYzDCGQK5Ld1R0nZcByE9z
ZZXMlSkw824lgb7k9u4mp9PsLvK9ujVt1ymvfH4Xz0RQIXW4EDFkARrtM1Q23xGljAwEUaEWG6i1
KEmmt2pCZGkWKSP5ZlQheHP8h+Ec0N0uu0jM3edF5Le4ooaLx9VNKN4HOtEG51DNCcbYKg1FpRNU
0YwtFBT8oG9gWw89aJH6nkMGoFyIMmMyk8tpPrQHeCY2IYISZUGey0i6xaWK9uFhxfOyCH37mq+F
ZN/yolKZRi7KCCpHkjAngvgLB51UVarC/nhw9oMKsEWO2T0HyZmJnxpPWM4kJs+Dett301MFuBUr
Z5mJM7nWZbRDAN10ZFIEL++tq0bO1K4ne9A3t2WV0naQczJDS4rgV6nTQUQlKMFEPZubiZ9FMiFk
BupwCBA0PmaGCOkAVskhq9d23m/zRuWpdrnHHUh/Zl9Xl3H04hjWWUKQCOzHAC3+ghrHUVxIrtN9
C8HINhOCGz4be0MY/XFN5oDmWM89T4WiToaDQN690Kgaebf1x8NFXjGfzJxtrVM4n6hjjkfgEwi+
TgRU3vrzzRLFHHqdEzkTJ6JU7VLDcikE/9xbARrSlLEhtldOjhdOooeHmtay3dOGRDeLNRvucrC7
AmhIbWaAUMCR1Nl9YZ5Eju7RPcJ2P4SM2bZPe0S2FptmqSQygVfDWxwMHaDZrydmTaMniGlxcK35
sk7Y1goHp0wXyvIHy1uhbhELoecIMLJdw1FX60sG51Sl14YQvw2XNoUoUev/0YtHtjmtOASeCItl
tVhRxMKVzHYNZLnv8SoWnRIL/Dv2n+mLYn6S6dG16JQO8jL6FDZqES5XfliO//7cB2fIxdEnhb92
UQ/w1R+BQvX46ogqxvubytKHA2qv4IJrqBfVlvfgZ6cAt3v3mxLP0LXsaAMqGxjklmZl9rcs+snA
03Y0wsQ2ym+Ro9DEgdXLqx7pxwRrzQ1XxlM8Y2CaPHiR7KALUGMTyzxDetSBrDtiYCyvvRQaG1Ec
NH8OhRH0/UB9Qy5pa5M5znYR9/7Yg/i6PyE9PHYvd3tGtKik7SWdMI0YQ0jQ6eFcffT3MXwowwaJ
d56ZI3O1ghtbAmvDqfYNkAFnL4IZckkQ3eeDxMwHS5hbrwZW7CAUkP86Mj6lWS6fsI2JJ7jAZhrJ
so4r+gv22KTSt77dbi2Bs0FPzlawEWD44nDvneZshxToO7Qyr/s8jCtCGY7qJeBoL+aJi9jIiVJ1
dz6h2qiYo3iQCzxOHg/fpwgxpByg52WLeStyPGbjQL+m8bBOZzmFo2JpYvog6ih+Aq566VddNbaa
LR4R7fvQIwCk3kNshLDTAQ0aKqxJRwgMksmyLEjmwIAB/+7ImwoTrUdBN/0fsFNy3ULGEF+gmAsc
1wMrM7pzP/o7+1VQPSMtiHeN/ywBcKT8J7hwlY0A+nC5rwt89hY315rLb4UCL6OgmjlfdWnOwFkj
+BeBw3j8TGkXlYQ5fAqg7oBKVfTOYQJ/UeIGtmcxtYgTU/+hQbN4IhiajZjWX9QLxN2sZ3czLWL0
58yV+WBC/XZ7aQffIE9ioyKTjfFpC5c0jE+zCAOcqRmaRGq718dpo5SMu5pA55RPlv1ghf4RhFx+
vbWRU0tNkLjmT3/b8CTsXOlIZWxaxPpoC5APyeW62eJlW3B1Pb2/wyeha8Gs4wZUnCESUSUO8VkD
A2NBvf6M1FUm7tLzgr1TdFVxw+ZOJgPXBCbJ4qiz2hRjCF8u4WJp/bHhGqpfniBLAIk5mM20TDUA
7MME4rka3GHocadZ70fiOsrA1LzKf47F3N/FOCbUYJZoKmq8rAmuWgEChPpKM/V5lYkr7eaM2yZ8
CsSpKmLTfEYFgsuQ1+QB8tgeShbJ6UB7Hk9lZevdWrR0mdPQQKyDbFE7xWXy9reUuPcn0W1ocIRL
DUmZvhAqothNhyfTsnSYTY+nYqXFDAnRWXuaXcp6sETX/gmvYZ8cnOB7FuCdrKSnLHk5JqNzs4HV
AvgEgQnyzVMa3rpO5hn86bj6fAf4ML8u5nymQGPxVG3TI59ZR10lojmHMfU7flZ0zSaQuw4o3mWA
xgi4dwyHyqGzSG/TW8gxpgGu6Dzcoq0+vgF4rBnSJo6dl6IDL3+aSBzWejOm1AQdhmPmoW0+vpgi
L52PNZ9TlGaeGxYwqvgFa8TdTsx/c+psRnvKApF9I0jC6BjDbP/gu0lpXx019l9Cy/H3HYHQWKY/
CwcfKK+RDdRIvWHXjaQfjno4rUw7Zr3UFJjP5F1ZuJ+7vKGkW9uWFWKy5mcB7SU2HhcTBeIccQNo
jhABO2U4GrmykbbR1c7aQ960cRYVvmopj4t9A+nRBy657ETBOTbztxWihwaJHRndPkDng2oa2Hkd
HJ3vl7hSaujP+GjIqP8uSSCJ6Q/88zQvB173AFzxTClFjNnErRqk99AuASfUYUrInwqVE5nmbNqr
w7bj3P334/g3nQmId9k4KAf62y4f3kumwHgjuopHDjufO2GRrT2GbHzg0ix5AFMORT1hm8suMYu0
II8RDkfhPByJsNGWhym1ERrPNcJK+kF4+xeNFK/XumLmmmLQ7OQvEViup1UOaohV/MeWEy184ObN
DJQhVEhldp/cF7RveYj2LQg8ixYGkQua4ch04DJs1BynnNN4xVnJAe6bjz8cvyEOr863qESDWl+X
ea3VJWWw/gxb3pQRdcGqgy/9jvMqSauadDcuhN98soJclg68Rv2JJMadXQuoiQ1tgK6pnBfKXYYL
OjSUAWBJH5y1Hk1kSrcpP2tXcKEjteMnVdt7qGPdkBI2e8Mrcr2O5xjIuYcsiyDbJG3nWNWJ5PHj
2OXZ89Jn0/kyEiseqdF5PALefWQU6D11Im0RZQz5EJ0J1ZkuLSbIixMjHpOwGIQZncMbE4mZF1uH
Lk7ITpySyeALUtfIF4Ayadmjnq2Vezss8XmWRf0W9YAZ42QzaTq5f1iR3CW6voGJZ2jqlBnEFF+/
C9WpRQyONha1d0LIdIn1M86HjtRQBxrhEamf2Clf6ZE/X//W1d6hno/EO+HU6xdJGznRyKpxfhjT
ZS1+M0EC1KvjABhwYuEzC9w40F/aLx4VxqzQLXNsKXVJcES5cBbJWEXyJ0wl3E3X0uOk7sHELmAV
Znu16MDLB5z5v9pRM09gu+8W2p/1AeY+wT3O+5imeX59YcwsFT86HyRiJhRN4k8QRdpXS5SyawTp
OycMIiKmg6lxZ+0FPbt+UShg/jpq3UzWHPn3/eKy7MY7Vn5WSdp42CFnkv1Motz+Wwco9qWHZoJK
efCmgFz1K6drYHnLXzci4wVzLgXszFydQN9n5v1+grhPuNZZvK6JejIDsirINfEitXIoXjIcvaQl
UhMDJeAC6jsWL2ukAj8mK52w07Du+fn9z/V/wJMDM/5OewgthjcJYKoQInNyLStkbYlzszKJuZPy
HWzXHWjvphhvusFo6tATJdt5I9WKDAOwOT9aF300S+6YGAeKuI9hScbyTcP5SkhzlRognazi510J
Bwy0HErL0ZwfnKeW4EbT0VVdlqj81pmwXyTNgtUjS5jXBAcU7QzDVHXmN1e4cX1DgDbdbiVNvhNr
E70hZ5b8J1y62FJAp8BYGEui/r9qgkc+mkmhBQYAwcPghaSrsq4VVkrjZwOBeUnGAM79YU5Us3Yk
NQkcvFfxfGztrAo7RXolp9aN0PXSbqPB5pSAq2wBFxM/qF0qknNZ6kyTizdvWketOfqEfk/pwRRh
Cc9huPLtnBUlNUvX7mqy/wteXuaTqO2U+W8g4RCeujvNUNDWA+7S9a4dfLdDoNrDuH3UCmsm4Fj4
Ydp8Ikx6r+PjmmAVrNbQnvAnRbE04+71xV2sU1cvS1CpchiIyNC9taBUG95S+T9nDDjlWYmtgDeQ
ukHvv2uSTTVDISFwSAwaeheOEndmPgVuzvFxHQ8Lb5E438sW5xGJJ7KJpxCuLiJl8EHcMCCkCGzV
Foz4aWEQKI8MuY4LbBywj5gIcmI3VDQK94ozp7A9wPSSuaDjaNpaiM1jCQE/XJNbqDOOJLz3++JT
nJ9xbrvxPkO6KQg1rApDO4WL4yDpt81yLw+fhg5FYgT5Dra7QFgzBquThBahTiucdZDdGUa4stlg
7ax2zu91zg2j62dgBrScqH9S8baBzMPszFRbFHhGfidT1/MXoai1hN+P7I8Qrb54scSJF6du/fFZ
ez0aZDG0RkadDaz9O14HSrckN/7VE4zVofuMf/QE0aH8L8uMlXWn7XyMRASYSca13gs/ODBrPjwb
hKRTiat6KbqFtEAL5hMMTTEj+TVx8nVhcJnVnBnhriiXjcOWEHVqL7+AOQESrgW6PgDI7w3PtVxX
uzkOY9MELJBqoPPtNRgX5HZq7HvZ1wEeMj5EuXKV+XQ9XWGWb6hHQV062AINk4LQpNqqzIjS40Nh
0BmNpZ914GLkHFVk5xyTsRWZGujHK2Lv0IyWoeFu/J3SOl+2kOPm8LN2GAR/gTH79u8WEhcoXe+U
dimi58EiZ6xS//f3h8gjdLoqyY1xvvlMoKLT43Gqd3+OgPG+ZUDLYfg+wM+lK6qgBoV1q95gvNyf
7+VrAU9B4Dyl7cw/FBIJDqda68Zg4PQo2F/cRarbDJYCNM6DGzlp81T9VMiKiO8ix9qby7ygxC4Q
1QnmSc2Gakk6IzxAOvjlCm3JV9cnNJ1RHzaSZKDGcd5gsC5jk2KuQtTK0TPCQZ75VVxMsxDf0tMQ
VmcWCQoeu81UZD+AoY4PwgngxqNeXAuPgLfU54SfA/XJXXWE9ggDgeVLUOQXtqTOca1yu10yXTNp
cc0QLUYxZftUrYP04EeRlfyBbco2TQfQfOF4L/2NiL4lZcvI0V640GitMjliLX5+XFwog9AMmkdL
nPXq8e72pLUxxx8LMzCh/1LOpGRq81nxucI9prSbOvsKQoKifC3j+lY8xVPaMf2m1BNcYoZfUXdI
KokamiuPzaOdMKlfulYwzxLdNP/tsxgKLeneeOVgHoKJjKMIwPovLcD7XYy4BvT569F4ejtYrmvy
1jEcUovwxrQxA0enTPBAOwpPDjM7nvODiJMZFpEfLP3KRkL3T2FQA7aL9fxmhzQHxi00puxXLydd
Adpu6AbBQRPdmwHnvjNDNA9k+x6ynliZlYvnuxOUVxQGXtlUas3Hzj5Sym40568ABMtKwK8cMod1
APNO7ZsPGRC5rjxhrOvfRYl47JOzUbcnUoncT792PPRASj6atWo7nj8fJrQrFV9ErYPeI8XHUve+
rfGII1riJGOare7J32Tb0oCw2qFp3WCVOzlIXu0rP1xGN7RrHiLcTCUcvGEKkATh17XbAmkZ+m+/
IW4KKonlYfXYHfsjeRQsz8BSRwSvvqN7SSsayt2goIUEnB36eHNM1R7+ttfwLuvdhsjAKRNHvMfj
U22BPAAwWu0lkS8zRRmOOg6rrTTpqHQeDTbCoYVNGRcC/NoC29dXlKgMf4MBMbXppnF0c1nmQ97Z
BqyT5R/Vv4YdirQvu3bn4D4XcVqSiiWcALqMs1+wh9yyaw8ubId+Yd1Oo/RApvr6OU37M89FLFPQ
fOZJPHNlVjDZ4HMcY+OTOqbP9OQ7aMuWiXX8DOS8LeMqKhKl1K2M6LoAeBEI48knzL7e2QFnib24
VyBjJ+M1KzIx3yqmpB8IR3e9ZgoXS4xzh4hq7HKeXkq0twE8Lt9YHLokPaMqzR5TJ+qYlQnfeDPM
KQkOqJJ18tj7GsokQ5/gT5dIoV6xPHYyZZ2bgaRGm0C8tHIFJZrQrpYxSfk+OhmUzaOYAjWiznV6
Jcf1pvw0x89rwt8M9slwhb+a32LO+rJkm6HNRnijYI6ZG1wzvvjuz9brZMObrLNuuSFZaF1J4F6Y
BOsaINS6OSJVH8hAFk7YOczKSZIzDTGfnddALPnZtOJ6D0uzYSH4a9jR2YgiAnNaoyVOYX/yFK6u
7wPpaqPH2e9nQq5Yghw6GN+2Qq1bPdBnzdswbaFQKbfB7WJonoaVEurAIiLHe6BmhabIvN85ENKU
P6QxTxVoA6Pd43ZI0Nfb1r3hfihc/2DSVbUe17qijSlR4x7dv0Ct1D76vFdb8pzYAV5k/uIzTh01
D/zA2OYPC9XjDg3/2Z21likDr9V+paGJj5/ap7BdzTzWVnKOqjPBp6FVFFnDQOnAhZVul3iGUpCA
yGqrbE6xRbpkmlrkGwVkiaF0AQ3A58axs8O6OkIOxoWwEqZo8kzMe5zO6IjEkbPloPE8POy0Ig5C
sZPqHVUEx2uTIr+oKdH3teHHWsSQutKnEJqBUoAiQ1kU9eMlAc2VbbRXudewa0uD8vKb0EPd+s9l
Nw+VbfR1WAqPupOUHjKAneMOfG2NzyKOQ47b/f0kyr+ARVjLHVIieCPfavu708KMu8scJiKDdQ5p
0Kt+3sIu7/Q8Oy0/LEFC5h9Dn/9hTXniHB0mBW1+AtqGFShn0//G3QWCah0c6C0IxNEB5yW0TbKm
piLvdh2Zb3CXW3OdvxH5TuzbzNJZawvF4waqNfPjkUk9ckyU9x0aB6DaltzudUBIhivkqvMQXcVa
p5CvjD1BgmjWnBZN47YSAYp+LjfHcApH2udhQs/5zq41oNjwkZFSTjCAPiwbxvLEoJbor8e+3DUQ
SdMZkSGTR8t858ZxaFFdL7B/+pSJAgzxNCvOBTgvctbYFgzmS9c3Q4tyXCpO4rhpN+uybMxhbnUt
gujyymVGUEaaV12s/KKt1cHWt0VLT4WQyRAeWNLaVVUVkODvtkiglOBMHkspTn+wtLwIgfm7LlIX
CP3O6lSTqTNITJAmlP2fgjawX0Bz0v7Rih+hqL2jKcFGhBOfaVLqEZnmQ91G3l4dOatpFc4ual/5
kJD1v5g7tRCuH/Icj0cNiNOp+I4xbdZM2RhvbSN3ZXATNjMQXd+/5pUOBFgPkAmJIo868HWggZnk
HCZb6RXkVvjKhQLjEEQIUgmUWSqISmTraayFJ6IMPZq/hhj/mf4WkDR7+NsfEVMms0I9zeRznAFt
5Pn4/MRk46MTTjbq7JxG9IRg/ZnkXGZUfxTS2KK/7fED6yWbNZ/tRvMhW33XAXLDUTvdi0T7fCqN
B8AVbUrtTY1qzLRlws0JnxEjqnJrUFgpWzVo5Qyf3K99VW0nqHNiYSi69107Gk+TEo7CLcJ/tqpT
Oooq3zYi8QFq+q9WxDJXCqAT8m2NAxRyG8HjtOUxLpP/EjTzO9LPF2ZMErpO74FMLixdQJPkkRxp
tZwkESa2Oh9u+BJ3glXRzQu3Ig81TOUchqT35p0g0JELgSEtZMQ5jjhKX/R9lCpbQ/DxDVID0+/A
48bCTFLRYd5XN4+9/yj1jZK0vbV7S0luHx3fDVcrKwUQ4Qmm0mB8XsVbUy8zzfpm1mTYC3BVT1Gh
uwVRRVkxPXYBD8KbV5A2xexPFoic7OEtp6w3zQTFX+7dnSVS7Fsoxs0AMCzBcmnYcrUjBeiHVEEv
6pYmzaIkB3qh8/br8kiUlgA4avi/Ip0cb2x8nIh14UFzG1f6faJKNPkRkM1obemBJO1CCnVJDrlb
stkkvFTsc5XY81qr73UuakKSaeOGvc1D5CRyLW26JFowTZQmEen/r104HpCaO5d5fFD59ABdpC1M
nl2t6W5k330arUvF7HjZPe1+55gByIx8EK5P5/bdqWmzjViEu3jru/dtTrH7yT3Z2MSLmSTNXvLs
8eYbrBJMJg9jy2rDF8PNYIu8l6blKUpWzPIIkZvJnfRyfHgymDXbqSwp+t0Sgsk/UG8U7tDsOdbK
wsCOKiqqfJ0oVn/NqQEVz9B86sXdOZkkZ8xUBcrapzDutqwOMYamb17hyKFu5Y9w8tMDPEVpE+rO
6kvyrN68cwpQdBGN0dJJOzr36e0BPT/DXQSK9zx5XzNLNxB9SlQHYGISw5TXCsIh3LZiuaHrZJT3
tcf/OmFQzUjTva2OXzKpd+K/J8EiR7S9NpOysiHyuG3XKf/J0/ctHX8xvJxK5YdqoYbMBbl4oWL8
db7VrE/L//QiPy1XH4tz0FCl2s8enrUzRAcPvhKMDJ/ga4xrPib6wOtj0lJu1TKzcUEUig36xJd3
GwdTMLWQct1MPE57p3CoR4Rcms6yNzMvfeQg1VHepqkgsDLf1veBCPN+OClf9uehrVdGbWdKCtWb
82qOr10RsVGbQq7nUyC+88DRLXL1TkHpu+bqYoq/JZOc2Tt/cUeS4VlXCfgrhx9BPxh7p/hT1mqI
c9wJoAbA4zAZtNoszhLecYS5tBBHzcw1g18UlwBCrM0I+61JG1g16fvIworVjGnR11pOIwSnRjAb
dPNj7QjqE4klerql0OjX6ymCCGbTJ3aoXaqn63WK+zTP2UDV3QuEp15efzsmYG4T9TRBD0OTTCtv
qlG73KH6iPaE8H1z9IYMCVYcJgF6H0vXgeq8aEjtylHaRkK375y6CBkiEuH0rIrl9HF/3V/YY2O5
2c4meowGjiDqIG8j/tXwxPOLsFTDpFOrLIZpX9soaJUH6CEki7NNaJ4BAaEe4IWDLc/3iv0aEzDp
5NwmhioLG8gT76CmwznIkEGouq2zbZ/dggxdltLD3ekbt/6+/srYwHc5r9EW14/xsUxfeEa2GpkI
dFcafrHRGhCfky8K8Ca1+JJoDvMGMnU5RUH07PHjDAjbPXOopNKlgbHNW+pJfFvvPXOzD2EOOv1L
rrKRITbFpbSSH329wyEbPt23rBx/WkO4CngIyYycs/lyEvKROWpXTiPiqXSYdUc7e2ROEr4P+X91
Hv231Ul3A/Aaqia/BFNoq4VUhfwp3rnKwgGTsSwd+5Ag23FoVKYQKjBtVdrzr1FRFOUwDQnw5jbO
MkEUbLi8q/cJ2SrwcTitGTDmnxB1VLYg0zAUovd0vTcx+lonaFAdittFe8pFu1nnnh6bQJC/hV86
3UbyXhJxrEYwwNUBxX+8TzJelcA0UYB0azFUWmGn72/5ljEZnrJWkYxk2AHbWUMBQnkQ1aywNNCe
HYHKjg2dMdkBgzdHTgcDfQPI69QKFBwUVZ/kGwJ/pUfuNEb2W47dfIWWFIXmVEiL4XeiviRvOSEQ
rq/VBftKkgXKInQwdxz9CVfSOYdfiKKuwcRX+2mw7P53J4xy8nA23vtvYHdnzV5je/EOG98Mzh9v
HApAVsN9U7saKQi9bKbxkYFfJCJwsrFz1X/74z6fGKxNktwbb8H54yh27b5mhq/d3T+cz7JL6Mms
ZMqJwJ0yQ8RFg89IBF0oPOGZNEQstY4PYd5ux9OliKtPMDXGVJ+qAp+OJWQqjQZkjLZhdOG4R33d
jJqwZex8LMx5CcbY0jNCjCSLboRPS4sunyHtmKMmS+uSaPNk96A+xwEVNvjf3JtKA/m3RJ1RTUve
USXtVAkK38bKftCbOTFTre8hwwMDFaxe+862tWXL+LYKjXIW9u6rrH/90CmcmEDgxnEx8sG3y76Y
azZX83hwH9B1uvu6u4shq+m14G3hmaq3gRuqTPwlpr4a0/cRWQl0VxzQBnIUysjFgT77kU3jbLyQ
/TEc5aGeTHx/rK5QAeOcygQpvMM2rzh8sm/AlS7QaHLvE9GV06G5w5XeEaiBxWVYoNH2qp8LKU5f
Csp/sUPZ7411zm7P9ixDLG+W6QmrzPH40i8VoaGQJ3ZKbLFlktun/8sEKkYx8ohUIcJZBJOVMTG4
J78gc9rgeahsaaC4rk+yQEREcAAHgA56ooE+2fRHRqqe+3W0H2KULJ+IT0zl8qgaWLYXEq+aF877
6PXr7nfU/n9Hyp4Fx79LjRegmZMcBYk3XRxp4Y4mjF7PTecW3ITzpsObj0dEBTy3I4IjmBSsBjJD
wBK+AGQ1BYazdcreQs95ZO6nxjREPiA8qtNdra1bCqEuHwcN61iz7Ncw9U01c/2HsL+fvSt6CzkD
EiLG3uyzuSzcQ9J9RoMwCz61L+Q9TFmxHo69LvYmOa/rclVUH0qo9EK0iEn+7IJmtH/JWuhvbCsp
6qR/nIBqFKdlRSDpHFUJ/1f3/DIxocO+/SYKg+MTEzcZpS/5/KLqZGL03O3pszgOUqbm8YK0RUCM
krVf/zFVhd2nsE91avbb+KS90lu/X5heAf6uwTq9G2ymxyAiRnVWdZ178c7tdp0qGv4LKT4gfNsV
EQOAuLJxepFdOPdLdXOxySlel865VokU+D3PaGMICzIhTVuS4y6Lfrzvw2DoqWICM/UZwRCnub4E
MDJm5GIkGV6ksHsQWULfUygMtRbX7enIHGEd+MNt4xIq83rCkhm4Mwr6nfaP8UasEK0olCRAQBjR
OcXVGGb542mo09PYQfASV7eIYXgsxATpwPH08xsvX7UGTaEjLXUOiKAwtAHbY472XASX7EbEsRQ/
sgfCCa7I97dbI2v3O8SWu6qaL0oPpa0mGijAs/iolvrZIWeVTxUqAdeGESxVVW+0eh/r+jxniLnI
nq8R4+cTvUAQFaWgxsKZtuDM+lgvQXSS51Tq4k/y9d642fSSzMsvnTuxZOkY/6nlsr2Yu9hQ1+F4
0FtY5a+PCQ4Fy2M2NtTCFbyRSnoUgEMS7a+WL26goVN475xrvfh2Hx04lciGDqqmt/kNqt2cEe4C
L3CPvKFRUqgfcIjALTGNWt5tJrkmRU0HwRrqGSVYp9hebvP0vyqw+LQRPeMKrHVKRGsmCDfh7I0u
rqC0JAsQo7bFhYMxRJJh5rBDkzi529TE/YG/eaKS5TpwgcFApvZzJJ0wRALxtIIfGmc2ihT4X21A
yrDvJ5oDnljcXOqToO2cC7AMYqBp9fLlB3+wZ0D6+V7WihOMoyCKr4MW2/VyYVKr8fuanhXZLCLz
78I03GlNMnnnFmnz7YfEdn/7RBzqLccUi5ysUKvciQX6SsBfid5UCxgzWJtlxK2/DSqNsMS8mLYs
UVodgXu4hdTm5zUemsYlSV4B/Tb7lgqWvX6qRnDp0gkauaipwcuqU2DdPlYZkcIY8m9AhGqsZpnp
BLanYBAcfVlPqHl0gHasJ6RYvss7Of3NKgl1lEbUy90OqJSL/BSuqrvHtqeCl7ug8b1dN4QTg1rt
59CLxnnN0LCyihH/lngeAizvy6/NQl4ia/zHW8EkcHOJf9CrYpU8x4AZkEXcqbZ7Uiqx7JyzuIF9
wb5gWOKRSHivV4UomIC3vWFJ3u9i4ff9MLv7szb0ZAICeuCDUc6ooX6Ibi7XitvyC1zyMIox2b7h
0scPpcihfRPfVjWuzJub56x7LGQNpRydLFMTdpPpyHZTwGcWJRhu9xr+1DvpiT0nbI8qOy8rjs5i
Asi+IxYhTC5WvgP9rA4wAWAmR936KO8xbaOD0fiwquSrf14Bb1hUQIO1QIfzRA0tmgaAn5h7mkQE
ERqEQgbp1LnY56Hey+n6KtoT5Ow/QP+WO3CZorHiWOtTmj4JO9m3EXamqjrGvfs/ISbvyNxuREtf
qbI1oCL/87Dkdw2+bEMYMlUXDHbrTOZ0cm/T51A86yLIuW9L9MAowGTwo5ZEMVNsK8HI53WD7GZd
6uG/TV7QLpuFd3ocT15IxOspv/pGtz/E7TBnKzQzdZqrJ2M9Sd4AXo5lOmOJes8w+HZoJKhUzNkq
nWKuqD6fNJcBdZLvy6PhGJQKXhp2gV7Ej2Rios7o4uPcJ+5zXtNzXWHb/kouXsdGsiWpN0pYuAsN
CRNXuL6E0YQRPE5hkbR4+H0RbLTtC6zbRLOTGuadgH+bP4+abYKG9woWF6918BvRNaA8VhFoZPcr
j1CGkNKLgt6wc4GDpKm90DNME/6SmH540ULaHm5bWWCcSeXe7kItY9HsZwMA5/ikqO2dlzmOEjpS
8Dpp5FKb/ZyZ5Yala3uL0EhJpiO7P0sXw1sHEYg5qUxuVBBOVcNgaskfKYsvGcy1pikf971hrw1q
OnZv4F4zxk2B01TQKuercTq6atZbbpXvsSeWqZQIg6URW6i8VpRnVwgtaWJf55VUmEUz6ew7eD43
wWs+dZIxOlWuz5dyKdI63S6GCOj3uvnWTVF/p4/+BF/vR613nqZUx8Tel6ZeAaQsJVSF7iYf2q6/
AABKvSpA0wV09vLn0geOhhbVxTpNAKr0ATUay8594hPPV58Y6hA/ujbvMwaAjg8rITI8csEOSGXz
8tb2uVU3D91KBGo3PmBxqed39ifxL09kNRnAvxaQ4Ic1huOcUqyvSXPMPoWPd9aVrRTdB9mThp2Q
zMeaqNkbkhh0dVxEDnQEEJUfB15/2jJQqMjR2OMVQZTgkB9fkeN5oG+D5zZkot9tusHkLtuN7f1U
wnlhSDmf1G+p4MqCTVhJ7SJklWrpcQnnjsu2KeiSsoogxsyv6dP+grvHn9S5JKNNlKbnmzKBUj+n
ZNtLZQE9LZdGze9I06Y75ARgHTiHVT2ORBbjPNaysCjs2QHobH1+aFeqgaUKJZgM/c1oT0qeSjcV
YXIZWWDuEELqzTbyEv9rbi2UL/RtcWqLcnHIq8RRPrzHzKfC2zLjH/f00M4arLxKkhZdPt+239jO
/9+V8P62JxS/4f357Rh/LzjDIasfwK7H3e1nILgap4+CC+g64tRBiR/gkphlFQo84DJUcy+dgZHv
nk4+y5YHQ/+NrnAGFYC7l5m4vrgqPfLf4zXuo8TQpKjf30s+FFtiNSFRapb+CGdv3km+cWBm3CKo
gcTSooFv47qpsZiymJjqTdP1RwAi5zEBYGN8BNOCGB6KdxFapDMh2C3z0w3Ps8Vqo5pwp30ExGc8
KTFklas/4Lm8bkNKI6a64uyBckJ/N9KPA0DU07dwavGWnpMUMsnL1OkbSYH9riIYuh1cZj93kISx
nQ4on3TSpr5G6gDDeb73bML19jMvk7Lyo0EbX8xuDuowMZTFV5/mED/Hm+Y50F9vC0kiukVmuCSx
aK0z6oQdYkHeRAv4gGtEH/tImT0SkTxzvkDEXslV9uKu9Cqr7jFDUVk5uyleXM6XceJkjDClFif+
UGzdV7vi3USJx4LdECq5XwB4W0sON0HLTWG7T6u3VMfE1o+/4N5aNYapuqwCQYWeUvKLq8q9tOuN
WIatvGXQmlNI6uChpj5z7UgC4+w/WnzAKVIFxKtadQk9tCVDjyd/LyzpmgaEMQ9u4A13rcK3sdwA
mqgROK1upSI11FauoAhQESr3MVYXLKZCkPrY92qPX7tOz12VgFDLrSe5roqcNDv/LO5Jwh+G1HZe
UaKz7O4y710Inqj/z+bewmaNJU8xqEyd9t/SuHVrFuhyXDITI7BdaVcJT/zPybHWG+OPqeBtHDyl
d8Ntd4fs+f37zyIUYyFcJj4P7VhiTvHrWkLSOvh+ikm6e6KKvrUSGrzlzJ3QbubdEoNehkH43Zav
Xp6jHz96gMwmJUBhiOnImfPX7J7eZUX0pDdNcD3D8iCB3cb/T2I1xnYu+ikRHqYYmAtHiqZ4OV7V
ZJcZM772ahY/bRKy7sXGj2KcqZDlYmlE4l+anaRMHMVIMPxx5AVwo7nP1SHDo+dOIwDYxtvv8L67
I7HEWFmiYdHxlnoOYFWLWgW/pbjud4oKjxeqkMjqJaE0LOQK2fVraLvPbaPlT7uTzbV+OsNZ4c34
ELSlozp3mt5y9IjtX6iAqyxYj2kMhBxJ3E6D5s98jjZWL10i22S7gal4iQtqnDfjcTXvfJdTHzeo
y/+ChNX0gehRZn8r6YPlZcNMJST0WuyBCGtv6gZ7VlbLBLgRChbvLN15z19sJ1FjQrkciVgvr//Q
UdK3J42Whdjtw+jTAmnx0YHlPCoyuGrxhk4mGdUy587aSK1+iRHL9Qk1UyYlW+Px87Q12COVWZIm
sO+2S1ejroLAhQivJ6mts5cbvUBtnVSPL7olOZh17SV3+5BNZOx0d5jxF7t0PiCDs3h//TfAXhN7
nbG38SfvC3oXgnSDqW8LBqpzJ2nx++NJofloyB8fiNKeapAoS4LolQdYsydV96c1fLX/ZqBylvbu
xqrGOiPt7mucdYKgBLhHJEFfWi58206v2A1pd01WQnHRkJONWpGDaS58zvPWHd3AJ79BEKszLFUp
z4a+q1zwlNXfhR6EWoONYgD4YfHbAz/Ou3vcu+l1iSuRa6aF9YA4CcfKR6WS/F86XTn54C6c2tII
Xyv/Td3NIVBOmJGMwOlDk8E7dmHJevjOZf2EeweuFtvyjw6DFC80pGuJoQ00/mqTJmPqIC/NuE+9
xfeDgcR73D6x5/xzEumLuLn8ZAhk3gk2GH+VGmZgBoy5FzwonnncS8eu1T7ROzjWKwGaUSmv+v9S
qJWAhCOh6DznoScxHi7/NepzTlzY5NoNztadCTaMSsMVTwVDL6sFm+3a1CsOjjvsvWQQRDZf7Fjd
jCwJ47DwAPC6KzhubLBOeNgy5Ig265+22D98St1jt4cgUmo4YkJkGvwJTT9xFsmNSETwkwGWFvpM
hElOUNU7bZHH0kLKEo061stsSo0WUnuCzr7j2XdNM2U6AWesgsQAV5/GkiDgjXuBbMclYQgQvJHu
mEyC7W78JGsHArUzChkGBUVWggWOGdv5md9ZMYFuzfw/GAPa1kANv/ACTGhNVhGkPXjgcwkw7q8E
HjDkxzD/GrBanLDy3E30gr0e6KPawrxAP/7LaA1Ny5P8qKjcjl1xBY0+BU501ESAdedkefFyWkhm
EV7cIKG1lvi4TsBHhCqNmR5JS3es0DX5JM7lcZ+tDXzW/TssIkMVLDaIaW3Ks9q1oQc2u+S5s28q
xIFyTnmew68D5pMwN6DeS0qudZqY+/MfU42npphg24hdhjtdPzRR1QPCcz26EMd8I4jQZucVyjAP
0v1pQs7wVyKbZ261rr5VTd+tl2HUOI2BewJ47/y3UnrXmnQd2EhVSsatrtl9doUSiDSmYtruc0Ul
nsQUqClLYQmL7OywPeRbK6qh0nPM2csGMQ6wtn5he84dlBt6muDBX2SEQMbxx9Yz3+DSnyj+35jc
h2w3t2ellK4IgqoGD1yXDIIQJXfVmt+dbIOIHWZt4hEw2Ivj3B1YYa6jz9ZmgJI/eVGVub9f7Wod
QW104jXTuaViCTZjoDUU2/eQxd56ddXLipO5c1reKHEKzecBcvbvoz+MOHD4xoxVqM8bsWwYcZHH
b+q30rDb0aQjw/e84Y31YYWzv73jNtGL9oxCXGlJBT7/P2XX2OWFSSvGBBuheqU7ZcC26fIFIlCg
JbH6/tudRmpo4x7XR5YzD4Eu272GNJdkZmXprk0e/jvUKz+0Jwi3CRuHs15j2r78ro8Eb5xzSC6X
lU4PcyRTiNoQLiMHU9pw6sopFrH1FpAn8GRn5IrDxQq86QGW1w4AKCK6ir8nOP72RQPGjxAU503Z
igxhO5LaH2XcYA5vMdwPi00UOhJPd5MezsHNHApPugrH0Dr5J8RoEQwJyTZOCH+sdYVwv1bMubHs
nUHo13rZ4RFhGHBNFfBI6NV73XeeTHD4hCM58je52WVaEPihasVcKvWZX95VUIY6O5iTcqoluE+j
TnYfoVUB/DqxjczIfn0YdfhrL3cyew42YSsYxF901+vmW9WkWkYjr08+0RNmlddkjnOdnhIRpJBR
wT2LPQoEfDajQccslVXptddpCElMO4Qm97IjrWAGJnVWvJ4o7XNNve6jLEYjQrt3FplmLxKkIlPj
UDND3DEZ2qdofT4hIZotJZFuHEg13c0Sr+X1NxqirsS+9I5avjASzpWnaqBo+pAVMcrt321G24R1
uQbELVXUhW29wZhHOskcFzrZ5VC9jnZy9IowlyggXwNYQ9SmzbkqjxvCZdrDKpoIdNYWsk2TXEGE
PXFrMkwUnl4Vfsh/5mraIi9tLrRYx99TCcjOdtP6R+24aEhhMX4uyXtq+R3/4ioulMypeBlzQUk/
4yqeNeAKcUi6qsfrirybz5v04lwrNWNW2fXHkn3yZ3qJRBm/WgwiSdBEmXozFERCLkGCNl+uxp24
+v320+IhdybFkhErMOo6BcVgzfwRU9P+DMQw14p4taPi1OUQn7pML3Z+KqyeJ+eP2/H34FGdjNS9
Adv7QiXCvyIDLGtC/FDAFJgU9gbHM8j/ZCXLYXGvTnTVryvlnyfqbkVZXlWvp8ul7+2955nhYTuB
h0dk+lS5CudENBaW8ZUShs417izyTH8D0esv0zDLX2l4uqT5C/wxHjPN5X8CEq8m40etdIgTXYPP
10kVOyq5Z0nmoCfbDlvSxSJ3l8daFDol1sVfVXM8UrHJGlozjd1T1nas9MTN3LvJoC3cUGXwEIi8
1jdYgNLtbXypuY2LH35QSCBOqtMoHpzz9ODnqsFTBrAxptwCXyQdzdO/oHJzC3Y+rf/DA2+v2LVv
CzGaQP+nPu9tHHLocfMz4WDgELEpywI06C6VaIjwEonfGaTP6OpLSrvAxUe8LiwlFqRoUgNdGV5X
vZuzKyFNrzRn93hsjcUwvJaBu9YGFO0KtJpeV0ru1JP/19Qjw+E34Jdh1KvKJqm5PTEclsMcYVCo
r2WhYC8wsCMq6aaIuEKACrPoDX4f2EGSv3OxVUfA7RFIZQ2NF3aalKqXdUOZuWXo/NTHKmsMdwGt
0OFNxutCFSt51yJ/eHu4o0/ZqxBGleupKmzItqsihPuBgqgURg7kp8ncDXnl33/1iRo49YxKTG0B
mCfzBsDSVEyclW6rmMxvenu8oEnePnhievJW9ZzxEQuVQAI4OvF3irNhDbtAA1NgJkNzptdyrLcj
HGOQRvnUBo67ajm66L01HKoLQAq/cOvFIqg9RUyOfcPGIaHewvIl44TjtziPTp3TEWxUKdZsbxZo
UC3YfRGtAUyMu1pFWvcWXVmGpC4lyToVGElOvAI1SL2SnkT6bcRUqMhTmmyqj5cIkImmTY5UUJbA
b/heo7ojmGaa+Gcq3hYH8aXqO+lqUUIcMdFEmWJYpbZoXtBLnevgx/xvQpK86Eh6j8RH9AsnGU1M
u1vW25NhVb58SJ8IzOunRZ1INZHhdS5gaRoUuplrgIl/E4NTEgBEcwu8W9bcTEgM9whsj+2D04Jq
viYd5Tq53UtR3EJhZ6FLZTQZw1cSm+YNPbcVYV+yYjXNfhSYpnhhu+WJPPpirDVBMVD4Gi5KlDFa
7zxdIW4hFV0fP5UQKdA7FJH4an7vcI794/wXD1EFZl46TJdogQ8jHGrcDN2O6154e2RCBloZxbD6
GMFH878wKMapxjIuCDoYsc8HokYvEcDKVPsFQSHq+ApAI8S6WHJPZxUQ48Waqx9m/gRMhYzouvw8
yZfatcoX7TXfSpavOxPAr47powEOMZcYSl5wipze01RTBxkbj/IqRSPFeqDikNdCJc7K0A95++g9
w2YgJm2/4n8UC/Q+zT2Xh7NcNnR8xqxaZWN6BFYcTqOK99mBnsg5YM84/T39DPL3dS6JS8yOSODm
Brs249gWkW5oW3aebczvlrw6wv14urKl3XmUuI3s/Pqkg04HmQMxoyZOfjkDNLKB8zR9hH1AAby7
bPBjlB076wVUo2oDyBvPrUtH/tyLxTN7Y1m1qZtDuhr/dzJyzd+ibSWNDYutOzzutnss07Co/+HQ
xs+eWbD0KlnOKUKIQt4/9dcFNARe0jfsC7EgToKC166PESvwk43CMIdWSuR+YPY9U4IPNiH4IN/b
Yw+zSgkfiTQsyYJZcBKvPh0FOe8uvHb4qc51N526v6QLRoC1Ht146N5p31UKnT9XXU7IKabFbmla
JNPC/zVXuXgOkS9gaOPs93u5lXdDcr6PFJLI2RGHbahS43Wj1/VzLH+nu5xtiSN6T5oUQYGCgyw+
BHVVZxqp8URfq6TA7aZEy74EEDtmdWMCffHLi1zpjvn4nv3DjZqI8ur+W4WNTx/ujvGHzU+sDepT
oNamJX6my2atQxn5p0vj5QHnYBPW21LpSpFNGxOkJxOSxBCtj/vgQX/7YcjWGIIGgkS2024s7lTC
U1diL8k2xEg2FIUPoaon0yutFWBY42kRe4bWvYu8LR7gYtKBJI0Bbov6UZc0esKkYo6QJTx4eoSS
earRJNc/Co+3vspz5okfLu7B1eJsZb1ZTWfyXF17FvS6A3rLG5EsbMxRPcJ/SE2oBGLljfikYQS6
UjBAxpJN7VkiiIp2PeL0/NfgVGcOsRUVGHLCAT5YGGXejfvW9faPyt5paLfP4k4Gu9mIzludZAT+
/XxrXtgsBUo2PMYAYP5YDmA/Kt/dN22D7U1fUSvj8/lDzG1t4QOWzLHLrySPG0HGf8wtpHFmxwf4
pE0BS43kInksd8H2PYNelAyPv77BaKdjWEHZDbeK8zwpJSa2koN/3pQ0yAoEwlGVdW+YdLEuBuNo
WobywvszKb5AEzEGRdpNEIu7FBevxlsQ7E1XoNIAGRlGIJcyZBKyOxas2P3JWtH5firu006E4ad8
utw+4hs6W+RUQfgHdNbRM8umbYDkrkEAvd8Cs1I4f83Jsv/nNv3cKZ/7w9HHR1+q67NL3J/g1abW
E9Fl7Xd4pHVF5TXQ4mmjHsYv6jWWGlxCNewjwCqS1i0WPi/9bozASIGthzVYBAY4+h6YbAcM1zIv
pKDrJSqwkANB7W9E6hilUSlKZX35b5nW4mZ/oc9r8SgRUN3sf9bp3aeEezGY9QRSrjLaDZy1Heju
SmhpiVmF2xRYzA2V+0aGsOra9Jf0hcuIDORyPU1Ru7f5e6qF2Qol4O8ErPjUyBG+gqly2E7vkVgv
tea85C/fQUaL1S0+Q8m2SQx0P4HANtGhGrcQK2LGYbOacLZ+BnZ3va0E9CPtsNbWeRn0fTWQ8qG/
sNemcWIdpfTxRXPBMnQRe2uos9+a/XepSkTDOtSlcGHT3ml6aFtwOF+XMcGcRjqvdgPQWwyvdoLF
liteG5QvPxLG0bS0YGFehNZNlCEZbmi+HIm3fI7q3kQFC+YOULCioTuK5j51NmCW8y1Td4oWn5JE
9gWQ8i7F8qmUOlwwmt61q8SuzgT7mpVEajDm90WdaOKxC24ZdrG34z/SljufbAE0RMeAwoNPbgy9
DNboCSEFN+5RGLYIwPOUoMp/sANXDmYiPwfaaQNE1Ei6aI6NpY90yqhty+6ZbDrtNWzXbjCHaELV
V/w2rHZk+QmewHpIVFtk1XacTG9Bf0ZGDslRArqprCFt4zxD0xFqdcabqA8RueK2HPNygFLeClzv
UQyDVELWvAedozpwr3lzgbK3n6e5MUMiw/rF9m3ReEygn22wnYNJDUKctgEQMzBBjiDXDanZr0kr
LCmKWCDrW1p/91DVy2Lkaxc+ZrPPOTOE3cL3NZ6G7mJSbLH+3lV+pVzhFGWvLJFEx3FyYdJojj6J
LX4h9O0QgrHXMuyIyZn7OQQHFEZF+Uk3Wt/wISHlcni2HW75Ef7ilnH5pl0MdCqS1+LA5Mu1sTUG
vlv0AabRnVTeLt+JeU0fpEk67K/B77gxB0sdOAPKGC4KnJnsnPX4iQQG5KyEshIzPPPzAGcRQLvr
jSOCciUc5EIFZuioH0Th2DzNDtRtvXtXW7w+gtrjKYx0++OXsGFp9ZR0tBVwH8sYEkFsTD8ELSNN
dn7Pne3ih+QnB+RiRRDvWncZZ5ebA+dZe5vmXS/E3C0OXe/E9O3YYFqjay2+VWihyNyZrVb7o6fM
epleZicF8Ma8dFi5vgggTLZlVFww2MtoEwUwO7ek2XdkF5ayQXA1RCROo2weapld77p8FE1skAGG
fldW9I4jfF7gk2urte3OO9XAMkqOAWG0Y97aFaPTW4CAmHtlDfeMIZlpprnXQxtfILkj2K4WH/Bp
+nIwlX87K9qA0IrmnLClBxAz7KrfHN4GEgtgGz+l9hvueLsfYkV2QGIPJScPn6IJ8Lnlh1S4KejG
tir6LO1gDqMcHmoi1fo2GKWjRkYhWvn29q9nyv/IzQLgXe+HP/PyuCBN8J0VVT6dMGskV/R2gvqy
5erblOmDRGTG//nwlp0HUKXGFKrw8RBT1gCMP5tHnuLoKml6JltfQxNyC1btTkkMItyKf9zOYlSa
4dIy5t4FU2RLT4IZd4InmJ51eCUnCSLM8lhiVAGFWkOySY/AM2slE+WlRMNWnLHcvswh+m8HjSCd
onwpc7FrW3JzY5AZhtxSJut3DJmfbiZT1jUEBpPlKlnaK3CMsJ5yno+mqbBqFP3lDtea4+PJPQlr
LQe4gQ0YPFT9rCEeOHzZvI/Qk1aBIQwvDifaj94hNghZuCwyQzb85Q8rsye3XLB/Fyrz3RZULJi6
cIZPwpcI17rADMrBPIXL7lr2gezajuH3mnt2PYOzpBWKsph2aja/czv+Hdsf/Mq+UCpjIX4+i269
+ivza++kUqMa3dQn1lgetnMZrh7m0Y8qVuy9WKwRw1CPifKylzNZ00JAVPonpIaUfJShuaCp5IyP
P42X8MTyst+fjhCph9Uo6ipdOpSIjHJWZm1mpJTdbvG5/X52fWpIJW2n55f0NqJMs2DH60UtkyOJ
xfYzLfSrkEpv1pqFxWihI+dyHgHyJ4r3hLHx3wA6zG/7mKA10iity0CmT6Jluo3qPTMg+c5mD2uv
K8hISMK3ghtXG4XplsOamH61/6dIg/zl58QkUzKSA9vdPbEeO3TgAJnopSUSRKPwAeGDTCF5x+lS
KuN/O791Qrcar6sNxyZ/kb01KDamfO7OK6bp+NbQl6zuwIOpLG64Ape/uGu3vUewdkSTf17l4sb6
LGrBlSxLG0HpTddBi/6M05dhwv69eOQtgj7btenDAng2pZ39n4SHlav2BaqMur9L5Qq0ifpikPDp
VN02nvjWi57Alza7KMYizUI/9VmAGBsgzPp16bN/chsyKNRhkgaFHkPKW34W8qGr0pMhmYuCAK98
w+kBAxXeF83fJofTtZk4gdvMgC5LKr03S7CwLJK9Bn1wARqB/sdbs299U2gt6DOiY3tJ+h5AOuJQ
GIOmFIPhLB73XirfYK4+cxFR/dN4e0aJ8iCfDZCley6pUeP4pHKSG57kG/wVBGkCWA3fhmxLy5NZ
uJe1oKW/xYQR12HqIXst3dAfYQTCcjMDEmSdwH+0+RDKbHwxqkn7zwmp2CS2Pi+fC71/BKxt1Pku
/wAO/4TojTaNtmqZKDJLAcjPqWt3dp4JU+QvZ4WSbZUD0xSxbpBX4pitgO1FySSqm5ik4SlPTXFc
WqSpuOdQ4gxsr82j3leEiKsIKNim9h9KFHvtB54rFDa8I0hn8wIfCf2oby3A07cgkxe3Z3OvRbWW
9TULDwm2pzgPAZmGm2TSqMFQ4pYmB0FDQHX92OLdtscIpKZeg0dnbXCuTHTiBZrB+C4GNzhPJWg6
RkhszuYP+W3+7Eq7+aJyMX+qrCY6e+PoH5PrRsLnybWGHRczqhICkYpD2Q82JBzuhkiMTQ25HMmf
xcjaupQbCopwurCnzgyt457Ssf2mpLZkTHMy5lJOh/gsTBqcNk2MUUhTpiwcdP60m46NHYq6lVBK
e5ubyK3tQqKIrb8Ojz4+DuzWFrBiDac/EwJcdNNdIrcqPYJuf01T8baQnQfYSTsb57DpwPf4NSqx
6pn4BHmgjgMQW6rwwJUpVV0kizkmDMBNB4KdNRvsZ+TbrIiLpl8YekMcDlfyBJLrcZD+K6yhZO68
Z06MPzx0Ewlt4QCIFmM51k2repfpEshl8SNd6P9M3IzcJbQF6f4dsSiqQozuNZo4MoWdPQ+hrXu2
RC2Bm4TramOACYoc/Ju8Oe7HsyKYZHzFMQVhcj7ik3nlyhPthpYlmfMSdcGBl6lCPxRh1DB4Tev5
UjHRc5nyVwihE3GOkdDGQD8a/k6Dh+B0G1WdAmIFRSgUdKbgRrgzGdA9iApWdKvSTVnp/wi7Zlpl
dNFghk19bkcnHze630+Dvo4COWgqLII6nsYoa1xHrfGDmQOOt4JfryyXOqIK0TB6Ffkzdrp5eW3L
95Tng2g6wvpYQ/CyuhVO8zS0zanQNs4yXVs2lAbBFW1g9UDV7MjBhuRiCUUqzj0pOuxeHJ5yMuc+
UCxXbs3F8syYptXLadNC5kXzHFVZL+rByzdwV2gRVwW04YlWvcjgFsXEppSFRF/DosjlxCkFdiV4
BTaiBwyDjOusxPCVxltaRaCj4tul9O/aKN5dBnQkUGMBGw+dtaOl+pjl5eJrM/VfmFC6t6gNnrKm
1dxj4dAP4DXwTsvrFjNgDzja1ftuEwpj+YXwXS80RbK+VonnjMDR9B7QyXwhUGrWk9CTClhEGE03
faHauoiRmuhsIzSospiAVPdsn2PEuUSJYtq2JTSXVs9y0vW9ON59daINFPSTGqPAm9eCYHJX5eEB
NCUw+DdurltHTh93GmYuTnrSbCM+9BVjdTlwwvuMqlo3d3vZ23YY8ZMhU+Tzna7V2F/k3oA/LZ42
VzsFnX41AFFg06qHC0rFUoAuKcTB8gBwWjcEyU/rFaQEhE+d+o3YZKtN/OXvpXDrijidaiG11Eur
O7QUbV6ErFImcAfdvd+xw7aTOS7SLhTohm+cQ72s9DqV4MJHw9QnyK0JnCzfMj1AjT6i0o2bLFok
kwtH0yrAJHiFiihOAJVHIYq7MSGaO96zADLHCYOLVWsuqBdfT5J9+Q5VGvq7syooAxJuR4D8mrgI
qm92m49VITTLfdHIl5ayObJ+xjqYWtPmGgfd8ODQT1+MwKdYd99SOmjYjn+njkzQ8N2jpVQ3sEYm
pydiM1Kj3TnzRyv7GN3CeK+I6eNn+NNv/jKD5fpHet6UKj5lWF0102dazrXRDmoBID9hIZ+zj04u
P5JqJgRDVroUvsrleYxXMRfQnVvTuvTAabIoIeqxkoYGYtsctJqADN6SazEX+L9Dur25Yb8CmCF/
FTHAGmi4MkQ517oWsZytdtVq6rroDsnLWfw3Y4MZgy6rqtRh+1QjLLMFYAt8SiwvvcX3EKwhq2Zu
H+RwHOp7k4CYIAwoFNupmLdj3GI3cr2NPaVnc35Ad5Y0FxS2ujdwWyl2f8Im1uQaCvDeeXhgHlba
9d/CLk9k5GhTZJ8ItLCLkdLKmzwhnMpmK4X7V6HkXwR/24z7d3Fm1rkCV1IgYxSrAPzQYqQXmMDo
YC/GF2lnSc7cJ/vPw2MeiPT/PJiSquDWA2bapmZYOWRbs0vZiu3YUeq4kcNB7wg/4rALItSU+TkF
K1GGEbXP0wc4xRpUCy1zmA9xhKhmC413ZUPLk7UYzp6M+2Wlj3C78uuyOaOSbKYgeGAA87c0JTKK
py716B/JvSBLznKHVKU6SqQH/E4Vqy3OaZQJTQ8LMKqBp2swRur3rGoO/CkOtOuuzfcqwF5gWVOL
JH65iS0FhdwLVWVMQHm4LKHLHxcYpABf2AJ9XZJ0A2DcNAMIUmAGtlyqXRCXtCU08/kRqPF5kozS
7aVOoVb9hFARAxSGhU9+LRnKbz1fG0sb/hnF1e4JAvRd7w0cbhv/8RJXWiFKQI2SCTdnnKzsbRYn
/q3Ofdu4c6R22NxtcRvk8GZd7eEo4PK+AFhIAA7bhOXcY1HCo4+yKtUwHokcNCmqPqrAZ75yBIAZ
Ogy6LqSI26Ok36G5wujOMrZts35AkQdqDLCR2NXLzQNDqoD3XY1MVKmaueOOB0/N5PL/v4Q+hsIq
3oCfeKd7BR1dtAnWCftc491whdC0TlF4W8MCmpDjiXcyy4+bzGG//I+GwaXBnurZy8f5lWqvh97+
av0kAp6L3nSOHBLIvgG+F2HdZYefv+cU3YSkLii/0mvs3rVcVW3N64EYYXervQ5NXZshlEAIwRbr
C+Ce7xrO0N2yzCdhthHYMihBwgOEvimbgVB4iWfSCLChmByAW4rrbYNi9nxcq0gbPn89fvHCbeWb
QcmK3JhU9W58SSjjEiLZhM05Y3bg7Nbhdcu7oS0MZK3+My+GVR4rSwxvC+TmFsCpV7jpovQNVDp4
XKN1b6diKsFXvsvHpjOMvj7ByZwAV4mpdZynx0gTW4hxA4lqvtcoP7YQNvagjCA7aliTMtVctMRt
lDptTD3R0IzUR1hbIN2RBxetoWR/tijpT0n5ykkzz6/BtsnUwW00H6AgEoYGowmV5v0lbXKkDpRh
sqpLLC3n2QPKfMdmLNDyKomESZHnfaMm640/QLk7WYO/faZk7UAN+2yxcOQtUB0PCkiazZqA8Gzd
o2yNHCxwS/jylkGvvHrP8NC7NmHkeGWLqzIn22k/UYO1E4tG72O+wyM+N5a66WjTGkW/PHxrW8PT
tUsnjggl6eCEG/IAGocGHSeFlEmbtv1sZp4RfEudXITEaLEqc+VBytKQBeffPL4VxXPWFHofhXmY
JPHESs986GBxcW7cyQ+4Zvd7SoVl1woUnKm2nAnKn35AccMR7vN8D1RrDlU+uHAJRo0ZzgxTLxUh
DIT7gxXEWXUh5GTqgefDCqbY+aV02ebEkHmJCmwyar5YLHQ+9u5Cj5+87+1FDz5RfIg6qetL4i4+
OqZosN4UoWroJjLGc3NBGdJCY0nDefnF4CTKjTXlea0f7THeaNCFfV7i9OrWHsQ+nmt64xwEBlxM
bn+QeMlOQ8YqVYuwIHvkt45Aw1HBGMIqzu8T+cbngGTJtK8tfDaQIW+jycqmDszU90GQky2gXQBA
jH7FTF/03wxTvzMqaLnQ1B+V6AzY1pY13HU6+KY7997Tc1irIk6GU/9xTYK98uXxlK2rMbDnHkcD
e2NFr8ZG9Skyq/wd18lsLIVLXanYRoi1T+KoMJ33u9Bt5wQd1e3/zVHxDWT8nEDL6iHa6BGtqfzQ
bZMZzSKwSg1ezB1aTvedJopblIHO/ws6nchu09fRy1mPlN3ItjJoQFrPKb9nSzm8RFEL2njLvbn2
qW42BY4TgkmC6IIQTXPeG9rORd5FNqONJ/Cnpso+CYQpxJFXkqGDm6SqZsqDewKF+zDX2U6NGGVu
Aaav0xlYnAHQqpgkiS9/kvwv5c/t/jfqb1KxWl/5hmti/H33tC2RKQYHEjPx43HGbgU1fBS7EQiL
BFj4EqXyvAvQwxj3Wt7kh71bDx/TEZ98l+ylov0Ig1Aisi1qyaKZQN+D98qPPue8zUjYpIu8UHlA
enqTDMWYmePhni9BxPPY30/5U/Slz8YHHxMojFMP8wnBipYos/7ABBZG630DT+NBAkKCbLZFhzu+
XUe5y9m9CoJ0HVBXIKDWqjTXWiWf/U0eOtAB68Rid8v2PBoeDicgJ7XZ9WTCxhrnsh5tDBqnJTNI
iTKv0d+K43TYDEyOLJOxDlKqPECp3odz9ztD55TayoeiosDu5bfKeBF+0yEwtuH/LyzR+YkEkTv1
K6mi8bGvNOGxfkYKvC57jIyOhyYRCmyG6ew6nXgRr9YF0FhB3kdKYJj7znhJ6WPKJKY6C/Ljlmns
FibY7C+54//grPBALWXJiHiu5RFx7pXgihuId5WhgR1zhJ05mLcWHisD7FA1AuJIoanf/+ESxA9a
rs21VPl3NjB+7oZ9DHb28NrEbPS1LWhekAnF0DBxkAytqyB0bsvM8BBzIbSBzJ7M9Y5gzzmMdnl8
9Awzx7Rn0zxxs8DoHU0ZXf8XTJz1BqqyNj1bNwiUNLHvIX07vGl5Ro+ZaU9CnzuGHH4ZhoyS5f0m
OCS7QZYyhMeOy6H7Bh7BDCZM4VPy+VOL3BeRhJJdR4FBTIyexZA66vZu5Sgkp/JHiJAMTcZF4WYA
LTcMxkDU/BBYKYDpDC6SKrHe8PfwMtW04ZOu+w/eVyZ2D+ZWvq0qexknNq/awbxBafAllwSw7/J/
6QDWCzJDIdQGzyB2t8y+0exNUezPN2Dec53ikF/sYl0bhPRJF1IsQYuA7+QSFjHsng5CNsmaO0sQ
/W/1qDT7UjmvlO18GU0aOsuItxcPTFByVbNUjkcshBVIzOzkb5dhwntPCe/RIbkuy9tvUDbAinrY
3PZwQurC0c49X1SVkYi4elt/KwcpNWSYtSR8SP861yncsLO9LcJ0lc4EVqdzvZ3j9GlRV6othhWw
sDD+RUMv8pL1pHHn94n5HGryzy9e/XY4ldmlF1DdLh/lyko7lodz+rpvZXZLbhcYrSMJydqrAYBC
ih4e8n1iaqihxz/4ZQJCss9Mj1g8Ik8Md4OgZTSpvD6RTbOVherPHQi1/AXRGogmAswRzOUqpRto
iQDYjQsaSYW4picy4FrFsKNYlUkS40nsQRD9wfFNQvk3C/2ElCSexA2M2jjG7sAz6W8CKSC8++it
J6/Sju6r/egLtR29BLGO5H93e+F38BdMkjb+0HarMHnmS25wxxjjDBfU5xorY/GkVYLpO8l/MVSE
Rtu2r8pfyC9azoTGUaVHTpVLtf5knR5slT8VqZafXK9TNOP3Chq6Y4KUqYW9Kmc64+vzEg4meBWU
HMt5T3DBr4Zw96SXAkQfzVo7NeyA2SYM/Lrs7nWaNYE0OLpNCfzsHxjYsN8y+II6f4E+yrhMtLGo
9mE4K/f7M2fEVka9Z/VWkiI7xTf3r4JLyVBBIzIWtmy4wk93J2tGAC7aKjer9gzKjE+JQAumBhWS
jMVlzG88PpqhOuuxooRxY1XEKHxaTEgoiHteZkZgGgUUBh30KHMjW+0oXckWtsVfrLQstxeamtYG
gWjhIWta/i01718f061+POoZkUWlmp6VXiJja0ngwLi05O8t/8VpLeEtGHJpj1Bi9X4T1RzI7w9g
OPGj+HsxdKTMbihMYYcaPwkBoa7AFXljUYuo1rivMJTVWWSWhoxouz0KvqXnMt7E5Fy4CJEqZJoe
JNkE59CVe9c749QN1T6u9IDmE9Pk5+c1G2bSWQsBBlfLB9M+x68CpFmCS/w3hZilK0dgQqXHPwEw
dQ4LiD9Q4WRb+tYiEbNTyVmFVQ1pzPR1rjzcp4v25uI6xf5YcLx8zZfL0rwHQP7ZM9eLOGUN6ggZ
St/YW6tTcRUqtrto5DUT69KHwHbk+ITvbhsElYPVpZD4rScgRN5TzR43VVfiLQ8vD/+azJsHFbmS
NIPSAeuk3aSm3R1RI1rIFTNzAuZMjvPRAT7y3ULEr/MGe29AS0coPxFEBHhICGlEdm6+faXOdgNj
W1umsd6Nnve8SswxCFOWUd48EGBJZQDZ3cO3JLJucL20RjLAzIEJam6Nm4Welym5DquhcY9DLY2w
pBeMowhTYkCqVZ8+EPSDRBMlGjcc/7yctb3vRbjDspzx7fCcA//HT1ceRK0bWecQXVINPIq1LrtU
dxwwR5KtQj6WQ1rbr+nJyEcVSlAfY1KbUIG7GjeS54pwtNtswLM/neHh+szbzm3bsPsfRZRwqpWU
iK1UZT7GOrpqbwEDgCQIUE4zwwdeRTep0aCywyS9infZDFfxvQmcGjHtxvmHjoI8m0PGMAzDIT4z
ZfUtZc4w8z+vzt25aOFYMoBwZ8pcOpb6bJCgaWf5hkH1NbgFIZxVNItt15XIn6lmcpltmBuLqWl8
bPQuKazvuIHn5KYOUxK4mMtlu2WEQ43B7OvvACUsKwDNDC8i/YLBE7HATVHoHtu2ha3zCfwO7iDJ
Lqp/6I7l/gUS+kQv2FdKbupXSDbwq0iUOV0xNbUbel5HVsU7eFivXg6vEarrEwNpRxqZaULf4Eu9
PXfU1n1xQi+/xC+2xImsb/F0EYIoXzrMR9oljf0OZ4ayI8o7oAFOmd+slO2iz10m9i2enVMpnHjq
Sy2It+fiGOIusE4OB4p1YpvfoyQmlaVKgU5mIJoAN8dX07kXxfWZpv17dyGcY4koTT6leOJ1sPit
auXiyAsYWM/DNfbpKvZUZyRCnm6a0ifbosaE95eytCk5/Utr5cA9shGZuT2h5TkbpWodQWwG7Ldo
sYTW8L0gD79N1oCF2FJgohisJ7hfQ8iRE76EHPQUVSuocR53i6INt81ymy9BdZT7mWSI5dTDuBpW
eGYK1WpqAl0bkqbBLiXi7niqK4pddyF3RnR/mG+G2x2RbANuvBe4psOjOqCGaheDr2qCItWENjAC
c9SbIgCcQFfDLrUhgk0th9S5D8fWj1c1poJ14JJQ1I+PPv506EPsX97QZBDoJIQ9QbquseEICEEc
pCNxpe2XgzlXOFlNOXl4AqwK6jUvVdqNQYO5qGg6s0SjA9kll/To43q1CECGqoWdKXpM4e2Zg5lX
LTQVntg1kiOJUlnTtJtzkVXk1wNC9CvjPTbJvLdihNlBbx6Q8J/AXcCKXc50e9wd5sOxWj4rvFUM
q0M/TFGrEm2j/2scq1HsIUTYyg3VhuWHuJPTv4QhnfiYhmDObgHTs+Keg1JFuy/YuENvLFs2J3oJ
UOB+6H/M7XbW7nIomuuompjpUquWQ35F0l6ni3eqWG1dyITFGrTfQM3RPd44uNnwzkko3qBpsh5L
OB5gK1n3ZOWIUS7DSZFJUztAXyOk2B7RVyvOrnhC2GlT1TfP9WSdcqdyme0e2Ox4z7yEeu4BU3WY
A69O8GJJCu3rQn7MjLSZpovtJSRECbsFuVXVbsB1p8OzFvVJfGN/958EW/7eeutGk3U1xgGowFXV
DAYYKHP7i0aeibpAgOUZGe8SoaWoCnUolnDFzb8mWUCOn6wiKDq+JGk/jxf8IJXX64iyP7ovwj3T
oPxvhQ4w1JCs4lCC321QtcHKlhUBaOE+RPH51t7TcO6DN1IQtZekoRmMJ4aqdyS2hxsDU0HRMFog
nO46XHhJW6+oO6RRKOJLO/WcPd4gSuatEL/qMv3QX0CKaAPDBZFocXi5igcruEVu70Z9vtMoTDWx
lmEtI0jYiwlYlU1rqXXIrSHm0un/mNF/AXsKvPGuiD5CcDF3MCfNbToJVGZSgHPHxPtNlVGOXmYp
Ez9ImxegXNTU+7bDRiIJSRtBN3DEiVt99y7f2JGhhkS65LbMslQvDR7iUzDTECjYRq6ptlwPlUC8
zJY0g/nfELlOuZc7oZe8cLPOsYOYKoOPKiprw2wV3eIypXCvSrEBXAQEDvZOmLDm8Rzlh/wAYIJK
xpNYfRCIHssMrvYuS818mmM4nFmx3f8PzsDWp6RcKS51Q5u0KYXW/Sy8SzbPLFYZZY6Jq447JSJu
e4MZKgcVEBGsI/zhb1fM9ooUOPxKRRCrTN18a++a3u6b829rVQo0YL5LTnm5vhhCtnIiFGIrQswD
+3QAZPGH8a4Lr0v90Djbbo+1oM2HdYjINVD7a5e9wnKimSgEbdXIHKc60GrG07L8JAPSYQS+uAR1
LVvDIS9JwXNWSf5ti5WDAa+8fKeuUn8NlBhGarWLQGMzu2Hrog4JVNP0VpWhADSUBF+NUbmNTLss
1M2WSynZ8OxUvqDBUN7h3BQCTqmWaAmIqkUhIWh7Ff78R/01Dg746+J1nuUfIQgb6byMNyvzVkPt
RUPaWJVy3kSNZj7qOxhb+8YsuZy9uxD6NlVIAL888AqxIZ26369hHbGHRgrCEwzFMLDMJmLTWhWG
V2hm71L3QO1PO9k0+HtG02KWcVM0QXpXif7VKpBlp8D0FIdvrC1A8PiT/MybapDguJ4V178+aqUi
WVbFZalaaSrrICCG8hnq/5sK8zcSrrjpSximktTDEQOML8oTcooVoEGpSMuIsdFWkJSAm6h6k1jo
WS0LYwBFRg1wolC/KtGLko2gSR6uyo6cWP8EA+bZADREEia78GoXtrkBmt/hHOwhlAS/Z409o5pU
nKGFWuAb1f9Q0Akrgktc7fLXt/3XhYeu+k7UjoIdQnYoqXSrgBPKyZE1CIXTbIBy0E25GBJTySUR
YrXKsrrySTo0EhrKNAfVGoN3oHmy1KKEDaQeoIhSsMocC/iYbdDlVVNF2qfwakPM6m8j+J+33jxr
sz9G9Tmd+4Bpc99gRr4/HH+6SZbzIBnXJbc86nYu21q1bbcnSL36W9Y8K0qaCm3Ky9VfsJgkeqv+
pjeGmsHGOZ4YuwkLzrXd91ztfntjBvAu0Mazja0x7KjbNbdmzuUisl3xwUpKHtGe1GtkORbJ2v6U
qN6r3Bmg4C3FTVaGxCZyHcoEfqUsr2cHMLPn54a6nVD5nfSL7CCuc46gevs3J2704eaJM2JRISLQ
4gZwuFNTsPVG50xTz/j+Cp8UQefQokIwr75M6zpgrG1jyHxtODw3nYFu042kGbarMXZoxlnAYJA+
3vb3j2/ObIIucjRLhUXDRbxse+yoF7wiNqgbPvkwENw5pHtS5NIYYFeGnsNR7C0RG0Ox5VBxBMOG
aiUyDCjxAmwhaDzsMGYQBwYIn2BvXJPiSX93R0UEM7QyFEmC0t9rLVgra2ZBQ/2axKR78suDACQd
AvfJj4Oo4UDMzW50kwvj+8X5x64wYMe3cy03eCvvRgnIBa0qr3nbFSI8+uugqKCZSxnYa6X9cacJ
5L2F4wQuh8Fllb0k+oV5bZHIXwJ8cjzUeHNYZgTxdxcJUEAdJq9bPwEk6gcwnA0XFoWV3W5c2yBZ
cruFiRwf7oz4PvqKFaFRW8/VRtHKNuf5N+tS0fbCLOzNJptEgWgKPeLUeWq1XNm4jImUr3k/Zszm
ATlHC1HPFyS+Nya+M47BNaKO/w8fYLC4eR278tCa9Ryj5cSQpP/XAATBIPWas/yOf7iTl5NaF3tX
BeKtXPAsZLZOC1NGGcvZibKsymYhF4cWf7nqbFapV2aimyylipjJshBrG7gGjuGcFmK4k0XPYgSs
xNr4wZRitTKZjrDTK5Vt4YOcRi7YmCDOa0O5vtpKy/u6UzfD13qAdWRvAzMjLPVT78xzA6ho0Qwi
vRr9OvdOh4LpCHK9DVL1Ganjed7okhImZKxkkelDbCkdAvkGBnp8yMmtlnICo7/fVKDpI89ORQT8
Gq8o/xldptI7hrUE1X/7e4wX3QpjfCDcKF0pID94ptvNniD61YcctyB5l2my81LCG3wvb5nao0yN
GeRN3SM+AWVsexmlpj2gvnGLwhRRflpi1BlKV35CJsngRb+CAYRWckFC0RBTmz1jbnyMB+csE6PY
2VH0YWGb8LNggqSfGLoY3dO5gxm95PEHZ0Y+dKrqbVfoDp+iwJXNbCvpf2p/wsiA1Y/eUuH14C3k
MifdMfz+iXQv2z26Xb8U6v+KK9R7L4ykLTld9Kiurqylqxc4S4o7EfwejVoQdM091hGvCRpNAgM8
TL9TVAxLtuqFvaxwVtM7sjYKCuJRkOg3WkZaDlo4g37stO0bSNDmJq2zIXwZAfb5jy71hAYblZmv
qqJVfacsZIrZDVhCBHv02ocOVaoAwf28EmDt8y0pMmctuV3vhhvXb+lNANBEuBCbbmj5hyjQafPy
UtHmjactiWhX17gIXknK5DM2qJv/+CGGL4dgZyOvyk+uhffTWhe4izRwVI/bReIY4gQlLk0k+0cL
bXOvsGCMYlW/x17/Ssj15UPoh5QG3V1tROtUBS+XhLBSGK4hYzocP4cBEm1OklyHczFEh4ocYxyJ
s7SPBvfGk1fvzuYL8EhyrOhZZZFLtCeuu7xaaYz0og7CrdUS4ohB3pHtq7orITLFqglPWlwi6ufq
FSuNBybiDabnHk4pgbLiNbc6K3n6LmuSumgvjSLxqhOHkf0r8dmu94RYjfJ/z4wBkoX7wRr4awYa
NfFFLQfnbuCjjGkmoQ7VWYsosgJ2T/VRuER//UB0u/8qcdLmK9N47uHg16tohPRB3j79qhOG7D7h
4g23nNOHq3cMqhNJ5vJPWOnmxx0xoURsSxR8tuADqb1lBIwNqgPGTUurtWilzuo+VkrJQC3TgU7Y
JgBkk8eQMd0f2n5jvSK4B14ZcpgKjojb0DEuH3mMbozP0ewCTSRCE5d9fjMQ3XDRLISX3LiefUwA
mE40S/uB3bCjdMi2EeTWwEj2HfXDXSzbefcHmLeShRmHl0YuyjoWU4YIyLBkdsmpRjn0HBWUG3jC
kw5nvzTKxNydXTC9s4k3edtrUnOT+L56seJGbyMm18EofQu+5o4qXW4tTGI/3Q6WbpWAMK23CGm/
MD0qXGiy5C7N9huZpCq4UDsHdHSDkr7pRkTQGgtUZ8Bqg5mwXsZTmtSF8w/Nka0VugNRwlSijVMO
8ClP2FBs/aea+vA5ELSsQ3Y73CobW1paGtKymhuySmEHBB8Rr/gHw+jpmm5+EkdYS3RKKYMw0wgf
WMrXoKcO0fTga+4Fh692ZKqi4IhTGhzfpWIMLsO42tcWTp++5ZYSzZWq0x0Dzr9oP/XoXXVxfo9O
1S7hzmYbsNBz282W8xh9dX76VCWRuT79EQPkvUBOWUFoiu3bBM7ZrC6KzPJ/MWyKp9CT3dKkllf/
m+lImJzwdJv0cgBQ8P3/sA90ETUkYSOsEWq3ahYbRnBYDD/gm4MVEVvMvtoAog+X6GAjPjXeyREv
k+e3I6E4DAiT6fGD9wKBLMIUdeYNK27GUCkkWzmzjrUbJQzWCefX+y7af+LMJrbqmJq53GKIFC+1
5GMSfPPy0vEt4LxzIp2h2ULCOYZxQ/lMKLYvTpmxRcQ5rnHRbkQ/5hJFahCo+gk+3AEpma7XThKC
eu3Rlz3e7Ivl2DFPxFcmbzPZk62B/ae9nQYaWNnniSBu7WsW6M+r4O2mR0Rwq1MYEYwQe41gTbAy
MkmK5n8cNlRfaykbn1PCiAhEIJhkQ0bM2LnfoW1wCQYrDxMRFnvspssC8LKpu80X34V9mR1KeOIB
f9VS45v1gajW1zW7ULhWd5UTII5jaTeXVQ8uxZSaDAdaOJDl426HBVO/Od6oLh2hoh/+2n6W79AI
j2bm68Jnl2BYWPQ2cDF+O6f4gwp0nAXk4YAjsqBEsr8CV8bJ08kp2I+MESUQO9wsQwcY7FV3+Kp3
l29N+/WWSuihp8BsfBDwy8VU7iGHkK2TYZh5LuotuthE8vxTWgOZJLmWJNBfvz2n+o1hR9KnTGRL
QJ122pSz77Wp2/ryVzI09Pi4LHpIWXByVQzKY+xAU1m1T54+bmhMox9SahPbfec2q32pyUNsv5hN
I3W/mAbbxTSkXEMI8W3+HlxV1oymMdJEYMZLvJ75yMlLxQjMOE7DrqAzVxdpoVM4xFqAIt5HRGQk
shpD+blY6gtbLUBzHXZS67R4viaMC8YDdJchxnZxXehSKQb4MHX7WUFgb63cpnsGPuwwpUwKWaQC
AcqADKzr7YQC2y4CL3kXHe9QV7sWUZZARnNjXgpWivPZxmmlxM6n+sfhIuQzsGB+I9W3ZN1A09t5
EGfHfuSkI4O58ZrjCMBfYq35naFn5pmAbfu3L5hQ/0ilC3dmeC65llnDGm5YcW1xlBwXMLZHYyVk
lhYo7dIDKqDqTS9BTRMSk3WSkH/h8GT/sprv82nrNc8uhJGmA0Pp1rlw8+OCMPG4O8Gvdgpn3Yzz
zKjh1oP0y/TKzDfyCrUgReDv9IytBT9Mtqua04gIcMEgvgR46oTNdZj564e4jyOuSv84TtS/EeuU
BJuiodjn0L6TtkP93/yTnvaeCDeRe+x/WI8IaFeGvnOd0x6q0UdUCYlcFzX+4iJV4nXOYvSoLM5S
GlItm1NFarBNyZS27dJ7+Md4np/3t2d2mukcSL1j2bqfWVZzyB0enE9+RRTDEWvNcsKZYKbM/lmk
15SwLM6KBfsj3d0SBVrfprtoQF5yyjIhqykCgVrjYlc9JAR4KHL4eiqgPj2jA7I0ligAPV0OdE8h
IM62H5nY49IJ2xYQSkAA4eKb3vjmTlDhz5vcFUa0A7rsdcctlvjhDKEfgJl9bzPWW/oFO1q5ehdA
KS/8uKezNwEgp53O2QASCH9JNmaz1HN96Ww6L0QFJsqGWzeonFPH8OlU2jZ3JRsA/v6PtlqSdT5N
okiuB5yavgDnAci62Ob+ocyGiPprre+yfaFVfVivtTCHmcFGof7oK+IqDIYXuPahKzLUzPApnvNY
5sBFYXt5C54TLN5YtyldsmtEbn2cmvppjvGG0E/UkHDIq/1IpU+93iBP82xn12lGwB/OyX0joPG3
ThWa33O62m6APWbn0y1793A4uSJdM7fcKogrG9lIV0zYWG5PoXNjsMZ8zhUAUaZKDc59VcUW0LvF
x3H4UkAYNcLp20Xna/WKLT1kagsernXEqBHXZFsyxsUqusVZTcBiARXPilQrl6kawo7Csth3TAm6
oDpLMg/vMKQS+pwyLjOQ/mTyKaWKPogfxx3ohDiWr8nrHRcKE5XtT5bHHrEhyg85n+4wkInA8Rqm
U/baGTGtxQ5Qzo0VDnxnjwrgnUkLvTkbshaT+j7axDWYK3sxN2DRny81NufQHA+piVkw1pOjIqVm
ZzgTjCi0/9xD7jRqsisfbh5rzhS+SR1xs6oXXd6YH6x83QfkGneaFWl7OgRKNEa8+DL8Sd0inWUx
pQt/J05gfXI6LmqOjtZX3JBQQKUBuSrD+QYIBFvl1ZksLU6KL/VuTdLFRfbe3oUnYAdn1CaqzwLW
OR+hQznrK0p6f5sscpnbBSc4mfjEO+F+QoTSvmbHC3BRgYwxP+sK9zvEAE5BS6BLvkZfPN7O9sAS
mDas309SpuJNYoKP/ucRDntDV1bOvPwBz0PpXcSeeEbLiRjnzCp0p8rGH54fIPfoB6J26yeEXm8B
BjIjJAbAL74e2i4R6raumIl6cUxPHgY3wd4PMcVZe1Z7hvp9IKL2KNEuC4G0Y/Mz1JPriaFyTbCR
DbWkcJnPkPIUPjQjOQG2TyidqhzLspOVVVdytwxj5IplCA5nAGKvKt7Hd2AoFc1526Zu4M6Mv5QZ
Yq4krsrBk+3tzKXRlK49COIGPiOAVS4IAvPsqk3CRAJBPisrzwK7BpsOHCJK+nbKAxRCHGzKriyc
OOe/Rvsvy3j0KgJb8/9yKljTEJYCZbmD0MgZJ3z8Cmz8QbFg7BSXtCKR87fhmGTjzo3QKjm963qU
lrpba8HB9rz3EYYI/yAWxUd5ZVorFo6cgTZ5AyP8HPPKIBULa0ASpc4nMUEl5Yzwt8+GbA/ChDAM
T927mS0oVAFOmjjWr2MJ82QAdZP/AZsH3i2OtouzbHJOIVJ9oisGoqZ/PHo8swKvL069BAG1bmVZ
GYk4EZLgX2o378h9GIYIUEjVviADW2p2O9QaIVoJ06GOY1jwCTUK/rYszZDneU/320F2FsjpbHUv
76UIZWT0Pg6cedUKpDCXudHES4EVe/7G058e4/7B1HkE8sqYU1rKQS7D7iNEkeDqDF+KIbOdC+Sg
aU48xFigqkLGMVnYfbRDNr8WqnxbKfuNpVVL7Vnf28etKlCrcnfIrIFQz9UeZ1uSQSa7k2Zu86yA
+2bE3hPdQS2WyIhLmjv9YIJpBtLH+XwUg4VpkCKtaLMxv0SVqdWDO9LnPL+A4VCTcwtXpJBFZztD
E4D2uJL4lrwZOzE19Jg8nRZEQpPni596qb5dwNaMVt/LkIaRjPRD0KE+cW7Ht/2XqF57dwuJaWo4
B9MsGtU23MMnrApRmyO9KbpeX2boa4dWD2G9FBEczOrp7V9Zz9oTn81VjggCXRk1cywAC7TegCDR
q+F1thLDgR+qlMZ6BHJ1ze7wuRjytLnP/Xa+NgojS9tJZcxN5ZrAsdZ+9fmYC497wOJjSeWGLyOn
V9wOJ1yNoKEMfSQPnK9ymFpsF0HUuzSeF+dmDdzytRlFmA4250BBVcctJ2zysVNAMnIEU0b+Y+jp
LZBAXaoBNw1Ev0+GcrG0A586dXV0ZMqafy/9xvRqx8sv+0ulfJIZvkyo1f3MTn0BPij2ilxJaOX9
nywEcmNkeOCbG9IuA19vw61eK3rGtt1Cyl4MRlBelsyKK+dC//jrAQRR120rvwJENkEsHacUp2Ja
FWJp0g3qam8+ptq4kMKNou9I4voTSqVyRiWHFO2i06VYOvLbsK9bPxshlucNfZhZy57Bmy3JBn2r
psiszUBL//rtxF20ZB4pMUo3L0UhNIwyUuBXFAbqcdPBY7Lq86RFvRrPbdiMZz/15tgDsP37o59L
Z+AlZm+JucB359ggFvxAHTp2Z6j8wMerS1vLduDnUdR6Yp86ZXHw7DhvViWosRgfbxT1jLNT8u1g
pGYe0U15iDZIyBIEOErGvYfkIIFJCgmGpsWc0I/oeWsY0Xb5Z6hkpHoqYcPTu/OodCiAr8KhwhLX
uqqFVE8heS+fbL6jcdV0KEOtajnrpYLl5su02WZwlKOPgoEphKriPFdY+QXe+acSzoDwqkuDMeV7
DqDC4TyXgKwnBET27bx/cAYnHkP/OiD4B1kTYHjs3LPxhr2PUOCi58MwP6FG+euWgKo7/mM8E7cs
ppk9TBeBcm/XHEaSaDiiXeabpTdf5OTZzQtZgs6Pk4KF17dS0MuUmmRwCR5qzlAqYCdYT5YZa7j7
hgyL+SjSAQ7j8Wl5zqucx6kGGK+NbNGpRWostBbAy/wnPesn7YPQPrEuI03q9Eb+utLnmrnbBaCy
fUp51wMjjza1phBLzsNRhbEz9hvjLxSLJMlG3OMU1GgJxoLQ9XF3/lkMfMnAQTf/WK+U5E6zW9QK
TuzYz581KzMSAd0pCW2m+Rn7UvcYtlS60z7qts27j9FDTaIcZSBw5RjzTKr/vQ/u0gIFrfwRYpTT
CMqRD1ZgZSfsETQDyEJC53B4zqUBgbcGQlnoh0uAm3b9WmerU4iD/1SDdaZjdjNWY/fllZ7fNW8Z
qQ6POIYdCu8ZkTWH+JoqN4KTtnbiY4222tX3NZ6+lrftuyqX076zX28nrCFJZ2qLgWmjD6R2OUQE
q50KFnQeazDydv3XJI24o25mbgkqTcX8g+4gG7AJUR5bJ8A0ovJw16ewtfqRM4rDBP5+iVi11IOe
x9gEsdAzlfRgUXArQ1jPdUCMHeQgNOogBjkKYf7xgYAAiqJKIwYpoF36viWZ5G5/IdeLEjCI69Uz
SMrlEP2aVCRhNA1OsR38/jDWPxJIHaIffnABW2TNivdPj87+9+CVdfPzEUMq9IHDHK4sx1w1Ixjo
Txf9Cde40Fm90KMiYL1iOya36+LzGuP+SkKlhlcQROkdnbWGJdqhm03FQ9n/2NHVzllQxa04F12f
YH2z3RN3BfxnyekSdJ2saP5/4nrc9/IYqU/ieM6ot6xcVWZmSs2MwEiQBYfd9/28wPKj8lqZ6RDO
WkmL2orjrU+eqZNW0PQ/DTbjn1Zpw93KUEgK9FxkDBldQQfp8MiFaTDCYSe2b6qOsk6XS1rF2Y3w
ZYbMs8Woh8xWXfAVgJwF474hAFiepT1RSJ17b20JhZZJ5g1tZfo0CJiYGLNmzRA1UtqaBDIRuNAC
I+9U7c33Gj5+sV+UIqAtB/9LVpp0rY+QVJ0EGAlz3fJwC3VoF6b4ltDpwSDJe+LTEpKv2ApteXw0
DC6C/ciQ5w/xN+7MkSibwAD/k5T8VB6ke6m3cCmlO3wTaXYnOIgAxoGN60jdY2RHV8KWWYGalCzf
gZ/HvtTNDVxZt80FPy7gYZrR2u7q5Le5evlNilMo4/KIf5BxxME2JlV5fpPDMhvVU+ouGY6+/QMM
UTxHaABF+QNVmqYnLwpQnP93nfpAzMlLPyPqxt0jYj2j44I05fgUidRysOM8TWYXoAxNkPoEAaim
zwBD4nr4LAve/Xn2OTIZNFWqbQTUVtWe1IM7+5Y9KdW9t3duHo2dd2c85wMLyOyk5Af+ASWapUk3
my9thezKQJSgZlwUQrEd6xFgIU7hOQyHKWvhEGms6dMNFj/7UrEOqsHKqPCK5upTVPLjJLfohcK8
5Kd0nSHiHqyhkmNjnsCuxT78QpqEoGJDMgMOKsjk0nJxS1PEE1zcaGU6Z/T2+2HlKCwf4PeComod
qSfPPc4CCgwySjSsv4fA0Jpu/EgRKYJWx60a6gN2ybZw3MXDe56OFE+j+2ZaPoRWXipkTmY2e/WN
uXsHrWzr9rhxnPAdrfWvkqAEbi1yjQUz2lVsaUmRlS/HieAh3mNNJ86+rHoUyQRrZ5GF6n0fMoXX
V/yQiJIHNZUYpC10mvdsqlO1WXyqN+m4R17oEFpzzHOIAwfm7v2h5sQwYVWL9m+bfeC5hJ21kCO6
rLuwqSuD2YVYJ9bYAeqCVQdWgEjcj1KYvvwibh3/2oO5OGTNNZaJDnwGA7VKjM7Ctxw1pfbf45m8
MNDZ23dGtENZZqGBiVisYaNswXjcRDxsTkQ4RGsM1cRu9fvwLozdRl5uuIhiD/n9f4u1C8wsZPsa
xNwSxVqeVRMIUMjg1ni2VOc52Fr/KqE/XjYYUsKFndVNfC9Q0Kqfh4AdLREx2YzHzgRhFni0Ncay
GYx/1ZBgR8FATeUFprTyfbL9yxuEY/yP8PuuyPwjOBYU+vLtn4NqDQ+Zob6sZU8nOl+jaicCbCJN
qwOLN9d9DoN+GH2dH8CjsMV/JJzduVUov/jeIDFvefdhKba/47kQhXnU4tPlfJ/Har3hF48jbILv
v0ZXcBN2ebInlznorDEAtjyacPk1X/PhbmJjCNTUQO3he9UtFj23lhigBPC9GVkZtZiUQCjaYxKx
EY1CbHFPabcizWnSk0Wjd+l9BiYaNchdkNS28a/11RwXSlDXGe/6AYVamIJYVu2PFISXF2a5ZhYW
ZlzFfC5ZudiRbsw3nY6Pllwn0MJ1xr5xrdAjdrO72jeqNvIdy79ncv+ST0sPFC8w5/KVGILUCVoN
foEwBT3OV36v+1sQQEwN7C84rZgkarGerCexzzfQHXYi9D2Yn2f/5gI7/64xUl+wRXbLahnr+0W8
KMVFuf+3Wn8R3t4dNbAY0z3V7vIyatxy4M7bo4YIvH5Ie37m3EmckwfWM27fZVlm0ksHptNFOxFs
eUaPeNeiDjaIcv1541rx2qnRCBUeHRUj30uGVm742b9hwT4mVOXd5qTfr2JeS4j/7AwhJ0Knk6kY
vOPYYvgRoAFEOLMtuuPyLuhAKHaEX94X47EKajVIJvyUzyID41I+u0hMOI29T0C5ST8Ej+cMf+q/
bVq+H0wTH7j7o8wzBuZXt6EOpjz/NkahTfj3IHKSPtItvmbB0Qgu0U+RjRuuSWyPWCACUBkFI6cT
juWSFKUtQHu4qt3qzVBZPNoWTKu/SQTvXnYip428rOKEvHQojKfIIxq9MdnKrkelYuiw3/2IbWlp
FQZ0EngAP0Dj+u6byWYnYooSUWEpw2r3FMCLYgvH24mS83JWL/tIQ62CvgJphEnqZyiogMSWSZbw
iB20qWDbefTAnX2mR6cBWdrbSkDS2WpWsJ7guE0aZfYv9AgB57LNedgIlfg/DYIU6Hu8tYEKr0Vd
QimZ3rEIykBCwHZ/md85XECvqMmTcnYH4QdrAaJHTVSBTwQkpSU7l7xY6dFVW36ygr8cK5F/y/Ax
5pRZ6t/r55qL/DQ1cxwHoozAB01zRjcNh/sMgz/k3Yr2atS1G4+eOvZNk4GKd5wZ/1ur7joT4smM
5ySQ5GDkzmEy8L0vBWipbELdwUdu+ZHmcOTIyOQJtHsvI73PnhdZxnvNdTpRWcELISK8wD5ghjJN
LaC3iM/x7zkJI7mJGbkXFrm84TkdfQ+u84i/RnnLhxxlwdzpKvYEELGdT3jqZ5bX5843Fwm4kjVb
2vxqSRmb1UsbofgdMEXvfDG4AYXSujxbAXd+h+AEZq1AufVUyhWcK9Ms9Huy3IKMktUPe9SfSCA7
VSJlGLhWxvWOToLckVXaTV72iJDPKvP1Z99mOjLv+uAvQ0dUsC8RTsNFU6ojAQ/DnC8CAez9B5A/
RKhBfzD5kcfYT1vu8l0GRfVe1N6Fx0vLEDxqZZT9GBVJbGUsvZnx9UBKHqPUANIrQk+86X/rz8pp
DKi1/JuvtSU+aM/phW3w8xLFsr6xMhjA+tyJhN+VutiO8Kd/DyMY4rRQZynWFWf4yfBv7v7q0QCS
FVaOxgRQv8DgiYewcBSkj4hJECFa+ZRwBgjPaLcGnJR2B4a/CPjGua7Vc0MtH0+acG+LhhyifPYh
8PCWTVTuf3NBYHz0qIBiPMDDW9csY6wX6+Ybjb4QY8Tbq2CrKJpsjkSeNTqCTK2SfjFmnQcGH+34
9BeOjfy1rcoIm6SXUFAszE+DaYnWkW9LaxSDQOvASs2Ei+IF9skfayId64Djvezr8dmUuGnD4abh
rd2lKBDL3gYfv78h8OqnpLDdLidICyN3ZvGxH5Qltcp711W0wMlZBVxsrP8jdvE8QcX31Zrt3o3P
dSr6c8rb12DXVm+lVRH0NRKWtz/26lavA+XU4JT98CHI0W9EApzDcxvdA/sdx05sQrLIu5k23khi
zMPqggdQbvioix/SSOFhFtuh5O4iUoOvfuU8/i0NbWyxOi8EtxIvL9o22losWPuvl157DH9QF+9S
5YMdebB5Arx9QD24lLnx49mV8Hc8Dn/mmBnGJ3YelJgzHfP7CJ7V0ZtnRuESbDPKGJb0Dix6iYKb
RzjomZj4h7aMjr46LptJMBvUsPDuklJ94P777XqLi5RlyB9t6vQmvjV2i9IiFHbyQkXEp5iVy+Qc
ytLc2R20Z6qnRISst9aS01uHcngY8YGfzfY8z56KPCkGXoIMT0DQfkZK8i/UQnSpmWt+CIJ78lhT
Y6vq2Ym5AC1W14Z66IbN3ouMlN63vQaDQUaDmrb9YHLSl5yjfqePr6pPqPiAUvQH0BF4KiXzJZYI
84xL36J1DBoHL+hEVBfrtDz6fMckPgrZivFK3fzQD3Rrz95dO2x5hrbOZJoCWlZvmnoymfuWZmwX
fFXsLIUIxHtPVJDR+g1ogT9j7O1Ppkj7COrRW5p4u3Fst/CL+7Fugd+lu0bvsqWD2Um/TiQT1QL8
/WOFPZ5gAsPIZqM5IrqAVyeTr1iNLsG+DVcmesVZ3NtFKsR189AW2cPFMO/IP14FmJ+vSYRHNWk2
/89y0WUeIKGuvNCTKDkifzTr5/64cAB35tddyxJPs9jpI1xTaaTVGVnnh9aImCZLsFZp8vYBjC4p
H/RNS2xvxBxiOlhU73Iij7nWoN4TDpKh1Ru5OraPKjZFixtX2ln/uE+w7YyeJuInfq1dL2RaCTTP
hFthN1QpAH9PxJgd4It1/GI6/Lrie57kOtZ+DyLpbTT9b99MvL1VKbzaDk9glv4H6gew0BW1HUqg
mR0QNiyVT5MsK8EQK8rtT4epTbAKr1XtCiuGS13DufMi1O81uijN89wFn/b7/jabE/8muHj3q6IS
Ol0ytahbyr+15UwrfZrnQu50h/uHmUY0DzH0FjqZ+4IMHnqp2q1sQVG2y0hjt7fDbD4dsIHMu5vZ
Ro0zXwJLC3cj5gUUmXFcMYMhQvmgmNwEc59PanoqSA2n4NQdvvBovq4YGJ2B1FMv5DGY35fuu1uU
MQukiGNq12m/a9rOUnx6WGR5PBxydkXKt4iubPlaQHuk1BRmrcT8xCocER+A8G1c9gw3REodDWaX
tVy9y45TTwmhxzH45wgC+cBbPXUSKAnVofX1CSxnhRn55bQwznhNm8lLdoCBQadNH6io9y9wtLY0
QUJvbmbnh7gSBW3BaLB55xfZmNPa+sXBU0xZ70BXTWnXOWvBjmmeopBGJq4f/q1DeNg6CY2AFGrg
BuTm7Vbxzk3FnZeKWExvOceifsPPr4+o4/PprZ/V1CfJARJpN00qZA6LivaQcesuT7UbhsqC0MGA
Z7fxFF3il3ZmZ2j21SllQ75ILhvrXj+RSwecRp2V6WgGBQKwIyRqppn1ZcliQDVK1kiNJqDiH47E
6Whyciz6P6PxPSJRluVAbE3/MxF0KTLfWCYPM7uNIano1aGBrirQLGwAcRzzs2yXUVqLmnN6TZI1
g7s3aTgR4pc9xLyqHZnaoRjVDWHeiT9txDYxcjx6uePqxKRugz3+hHnWLxD58nZSIDOE1grHyCX1
8sx42HLt5TZP5a24isz3bClTzqlXewSqXEVRjTSBTjyJHjpxMTnwbSBjVy1NH2mlz4dYnPYrYDdO
PDCpL2LeL8PODoOk9ncBecyJl2iZ/hNFFFKj/eax8q/buABnj4KsjdOrYoVP0lTxqGi2ldiQXWWD
RqfX4cqeWRipuHEOtHwjX2ijiXKMSHzgyN86QiWrtCn8IpR22CSoO1tFM0LNr9zlqFNDoDVD2hoz
BazdYVS6ioneSvZsAJXE2ETWe2U1XqzTfBLxETTl6XM34qfISp8Z51O7a4dhhj/my0kW4ZFB/pqF
QvWoOnH2+cZqEXCvuV194ydodDBlQ74heoEKkvh8Ev6fGABn9Otq12r2B8RkQ1RBJnhDRejP8BCz
iHhkkucXSEqKyxKwHNLQZgDqEs2eyjc5bJ+6aEIaaY0R67d69cqWUjxA7tM2HZlUTSbHiuZcbHTN
QDpW/4v5DqTCM4y0OO+AYQYpYxXxgHKHE/LdfMw2UphRjkDfWf6DYVx8HIWAqmNHZuNEcJ+g04VR
H8cx0dMecI7UX/FTqvjY2d3iIim+WrP2ttyvvCzRFuRFkbYEQicmN03ewsWTIr/aMtqkbUGSOJlz
YG0SUv5pVpSmenMznWKrGC4N5P5JBkpufkaaHcqhWs9w1mt8U1UJYdqpq/wS7ebuJW6k4i3Ae6ug
nROSgoqiDdavGNHlOAWOPz8O3TlfKNGr6RTSmrgsLGA9CdYMaKKEtIM6z73WMp/JaJEFatlQXK1Y
/mnS6clChrltLLfPOR+a7PLD6ymkIbSeRG7BRApNcJ8rBCK3WfON/lobuRzx2IPAStaD+rWDJouT
o8eSNHlsvxh+7+RxuWuwsfpsfiJ965ySgAl8wU5RbsmyBSmvlZglM4FDJxhtOVZTlt1R8d/deNg+
8HhrWrlHjpgdldUwhqNuX0hHbUvnX8iRrl1IR6q4pDr8WKshCralzOiCj/0V1zMsAuqK+HXgprDM
1JwfDmK5NEX5w8cGd0zcZE37VYyr6G2cjRNeZ0lwHCuFmzetA47QgGat6gCBrCfDXeFufAKFj3+E
nf7qhWZxo9goW+zf9lRhcl+dRBBYxFcwnqugPHsY9ulNoKXb3pQ2bC+RZQ1t/1SvqGq3F7euDlx8
S6aNbjTqJw0SUa9SmpxPcIfKR46xqrFt53H4duJ0CCRcW5UkwRYnI6wiFcNlTGKIe9bSx+sATpum
/PoLhS+ENzScdi1SZlhlcQiHU2l9eB3alO57D4mOjmrR4AcU7SsnF5/8oI5fowVU/L8keDriOvwy
vxIV4iVDb8K9anEFHFg+HS18N91P8eVregcfXV9uRRqRGBC2DoBPGbcjyYXUBvevgspA394FyXn4
eZwJqHnt5XMtZ/py6YKacmemqeZ3iJ5nMFh5JoVIMSaSL3U4cmD55rdVYN0+3ilL1HfOe49jFb9p
gesmowivAkRea4rKcQCZjg7apkXxq5mx2XVS/LjZV0qQsJI9lJ2QxZcc+Ai0263G6O7NHUkgioZf
glsIcnXnxs2uAobsz2prXk/zpfCCS17Bi1jwqzU8IZIKxr9/MRkz3zKQeNwFqusWiRVYWMWguj3h
iuYyFCChkjcH8Iy2Moht6assgk0gOG3011asFm6poDJ8uBZHV2YlgkfirRBgxS4jSXXVGahcDurz
wuemsU8FrxFXRBfg82c14+c87bmtLCGuR1KZgpCo8tFQ3cAm5Km6N0J9OhEIGHPCdTH01kK8na2G
j4U7AR1iJEmaI0rzotayRuaepBZ4UZ23gLHpUranKLUPwT054e63jNrSS+kWfMQiYE6AvX7Q1HLT
LetXAj3u10NHU73acVfd2z9i5MM2kZWT+kydmzfSUt6vu0wP50Hcdf+IkftTeJGo+EqtOBcDgaDT
Mnlll8xHj9HSl+G+E/T6WCzKi+YIO8+Ri6pMZJ7hLAwwNSoHNPziC0j1uLWS9l9pWpo1sw84fwwe
esLz8r9+AFFOxZKzmbfQ1LY6z8t5Nf0v3NHqRg0IYPzwD7fxuci1qGC7rg7C7LrUXIbd22Mm/bCj
JdxuJaBlpv5U7iTY8Q96w80HHVJ43AVAMbyvmmsXPknRKkMHFxqqjWIsnO58zOTEQeNWDrqefDnT
xES1mUi8asw07U6Nyb9S5v0V9EhG+8D9Y3fsCkiN30/ETL4K3EZb7/fj3KPT1Bv+0fOCNQvH5UNq
O6seq6eiuDx/9icucUr9cRt0NpJ/FYaRRYTinAS0ehJJaLBKCruxvvW86Zq6gtbVhMGxzQEJJ3d7
L8zejZOVemdves43kXDGKdcyMsce9sU2wh1YKzYGEYgwiy3qnmRU7FvvMx9SHOy+XkDZhFPAL3Vl
ZYnQfm4cbs5AdIzCQgVBVyllkM6psOuvot5aULcuLiapJKx/X93eXu2WzEvSD2dBEb+SLXlcpijV
xeFE83xe9KGa7VSzrjv5Wn9cDdu1v4zOGb2m1tP+WuA05r9rF2ZY8PYrrFAMktANKL3poGM9xCMS
/0vYQttYszxeLfX54TnPD45yIOJxEE1AUrsvqXN33zaM55s6nAm7X4NnIiMDTsRbFocXqclH0eo3
s0YvTZqlq6M8OOfWZtPwNy4KsS6zjg8mLTfB2qyvBgjS8WHEqjKlbkiPHERGbkHWmrVSvOprW2cu
mMZ8rVBJRbOkhwb3BcSulRI/yoBxfQgYlR07Qs0nyOVBc63gBFvTdXM71UpGAOVmpCeqv+ynVChL
C3PArlyjdEiti6vrbbyr9mvjPFnos6O2tI52qy53kkP9Y+lp3XDzdl71JlB/X5VYtUEng84uxi8b
8i5E/5EbEjJ/IC2Xfoje1qkOXFrDBok0nr+tzTcr9EQL/u8y7YYT2tI6cPhQ4AtotWvxmAiAGZ2t
k/bz1MiKqxs/ttYiZFyqhOA9gO5T+tBS+QRHnKzZ3SgSi4Tm4T0aWfatfBdplN7fhOcSpLKi3y9s
abeYKE9Bnq2ufHukAka/aOceXscTv1X2pG9hZDY6TOk8vgsf4XkCWVA2FB19Dh2EMxtMEin70HyX
tfkwvNODAI1qDHIuGsNJHnC7tmxC7d/to4RG2UKlpsLiZEn9Djs8mWd2Im25dMfVVxwHvKlG1mtj
ApCmIirRGKczh1Xd8I8Txur+WuBEaEbVazFFTlQ3vZ7mBTZb2Aau0aN61jOhyX0gWeqEdm9q7ONT
QlRxyNqZHhbgv7W49lqp9RYAr9+JV3o8UDjfi2RSjW7RzIKHDyST8l32xx9J6GijjUOTYzJX3etN
Gd/AoY+IiuREuW6+w3uB1paeUNI9QdqDl5tSQt7slypmCiPb9OrDUyq8i1pB2er/0ZHWRCp1wdT/
RHXIXv43/PZUEEczc9uCU2FJGU/PmQrX4pvWMbYYVQOcsiDKpetnnkdb9lHzEOiT/OGgZLBgQTRz
v/lpHaggz7+ofbr6/Itd1AcSPWUYjVGihNU/Bdqpdm/1xiquwfN1po5uJW2pRFM6xEBNiabMMMxZ
TVdMd6PxSXGHKVf5Fo4Atd3tF7eziCvHgN+8Q64/5++LneKLS+/aecUO0FSgm9yVA5nIqYvWjedi
a6sTLVa4tAOE7fEJfFzSsuzni96fttO2Jxg1jLMmFgfxqa6WpGLzVShTmbcZqRxDDhzEq0Yc10lV
gm5q360Rt9LKMRgVsn4Ruztj577FXUQwH8aYCnlmFU6An0xJjlgwUTXN/g/EeDmlCj3y6ozTygvS
36qis5SxFmeGL1Uv+y6jgp7CbGCkMxSmRKc3TFhJMoV0xYrTLDBUGgg8bNmUI8sZxEpxnWShCPXJ
UJ9If/OM0Lk+SjBnbNsePFgoDRHi53rqPjIHYcMItE8e7kegrb/+CxjdiB5eTron0uDemd9uW66Y
hCJ3DGFJBFtgPQ9ocW1rpsovJZ0FGkjLMFCnwVJlfzaHlGn35Lrq+Kl0wpth8NFB/ax9tgmJPpg/
U/a4SVThR0/W5adlhdTPaP6Y6OOr7vmkWyBxhu7HeYPs124XX7nFOvOE+LF2OjsaaAoxLLHoUgzY
buQWpWfTOiICCipQdO/UUE/xYtlxDp+be+G6pqODxdloy+Iypb/gyz3H2W+WkSP8IaA3AtYa3YPj
KgVrSwaEyfmkUXKaSrT/1g+XMM2N5c8JtaUm9dh03IjYMhz7s7jBpeFUt2HgqoK0NPmC2UxArqRb
2Mkl5lpS3higp7sbALK3xnti1fJYGVQAHbd4PIXdRIAjWkJK+t3VJPj+7igDFE1ygvuEAkT5DVPO
hvDSpXnq5Muv89Ul2Um8+UtqJdEu0kaKcTaDCe5F0MwsOjivzwuf9Q0OLflCzOaTzK0k29SL1dp4
V8gP1O7emLvuerH/oPtBUaxFH7lJ9IJeQlWF/f200hOoYtmGjEZbmlmf+GV49Vroo2zgeTmBH8rI
Y25yhEu3x9EDeMfwuJWasIXuHhPECbSMoh7pTfBEMSNL6Cl25rvFfaCygC1Oy94iViD/r7FFMxyA
8JVp9+E/Gs2cOeHCrVTmldp5UTRa/Gh5c+6BXJvfdky32mAF+CUPsQribYVQ+jPyVjTstpGJ+t4B
BHyK1VFO+w1uOvkx96Vln35sOHgfIK1Qq1/tekx/b8BGgv40yG2rRC+K1xIYZAgD12MUAnUcAaR9
ItY+YZZE+JFpC9P/OTLgLWqe0jbAnci5AGF/dGznqUf87gZFPTWdVO+CmURFsoRZkVo8aZZ5MRqs
6YXaertrQdq+ZdKvflK1ciXv5/9hhUAfgIsVeml2mJZNcK4jeHiZyhgV+eJxlYmqVXBvWK9gOqsC
AysCA2jZZiJ64HQAjzFMTOGUjZCswejVh7o8sVWhHbAAY3vkPufEzXGJRRKq9lRK7GuNd/laRWpZ
n/UgEXh2ENxGbQ53teHg78WNYOsHYv1VnED8QkejzWPcZfX/Yihc3jcq3JFxkui8CvpatmI3VfTq
surywPlgvPwKvJOjDHdiGnb1YtSqQcN7Z2wA6vjCqnjWFM0b4U37bkoi4pqtqJW6TF3BwXWWJE/l
l+qUoU8AVvLwTytnQ7DqG+WIr9clEloeaZZ01KuZwhxPDJ57tkR7ql3US3SPYvRw/5NUn0QDuJf9
kFX94vuyUXuGZGHNy8DWW6qugp6/N6CchRj/8EsEgP3c1KKNVxOMXu/ZfVJ8qQ7eo/GOQN9UQ3OU
HatEjHpHsYopVwtkc4wx7gR3ctPzZxBFuOXPXYGlcTLmZPaCfw3lIsy+DissoxnX5dbgqDyWiYtB
lAJmasVQc0YDMajIAKrnLdrMP8yRm2pAzAj5Br5qGzVfxGmv5SImRUvCbqRPU7umNWVZyHGnB5+0
vJ38yPYbGd8lZVwu+Lew9KadkYmBqyhWKWpE0PgK3h45DwlTATnfs0c2GNBec9hflnYaxodgz7xE
XPx4tCl0lPbNlx7OGt45vLnm9EdAZRIaNE6FeT3YnF4cLai6gEN1OGmhmrcDhaZven3G43Kefxal
b8GZytVgc1aWxEKEoezXY4jPJSkhcu2nK7QvE4+ybgyiNMk7AR1crkiMIi8mOg69P0RoKds0ugQc
uS9YGhp285S9Bo5QBhlmBIEMNdUfLoiR0gqCMo+mVS7Ih3Ppc/xHa5zDyrkcFoMeBFnVwtRp+3oI
0laiBVzPfspRuTuvzVZ76kGoeq2uJNbkqVPQHxX4p4tD5+1cM8z/ziRYNGgAP/THaPTnb1JogkGB
MxPio829w3EeF5SIgkMMSELGj8suAfGIzNkLJaS/5aZoNRfRxg69fFRXV6vniIrRje2aR4Bm5qqw
zr8XjBi0w9oF4jmE34OcyntwmoimCC90NIoKfsGvBCIf5/t4CYJiAmUzb3iUDfLjv2e6o8S7R6zD
s0QrTmblh7j4iKMwz8brMhlChLzbs+dqAkK9nmrbcnND0cFtfq2Hwt1fID1IxYFbA7XNF+dFFbX4
s9jsaw8bnXaLk9VhTONM8lZypOqeTgCL/dnHcptlRJEyQN52nJVvpo+zUlpgKCTmibOPv6wMBaxC
Ko4Ve6SdlloxPVreeZR8Zu9YyKXcGCNA1n2f5/2wta+nStxlu9ss8+Tjun3nNxc1dEzWeyqd5PLs
hbmjRMhttKFFYleFMVV7J+F/5KpEjgzT5tDJNyT5WV1WSPTr7VLYg3cIYKS/gf+lDX+y/2yjJVey
FpthMlPkAgYrQQeuThby+TLrcZSiwWvJv+c/M6IDekLY7h/h9Yl++voWWvEQo3BGmQE5jipSv6gB
zKVE5Ge+KuGsBu/HebIcrqbAAVyBW4+9Tk9xXKkvlPWd2lYRCGk7DQ0wybf6LrYduPl7i264FKuQ
A7mN2zPPVLWHxh+bBGxWxnKnvlzbst706SDiKy0nYHGm7CbKHkPVwn5cctyD0RF8K5tvgV2dS+xq
wLxz8ZDKsWcN581rjyTgvD2A9/CnLNJX0ZYAYTVuyFbEvUP8TyTPLiR9/SeXjk8aDB5btiKiDAeJ
+TIfs38aqCyqgkI6LYOjsNVRBsJTJfzMbkgxGokH5ffaqW/WO4eLGsSJXqSTsVM6zTfuw2UnBiO/
/ghJwntM175KRzgMIY0BdRNZXUkg6L0bsMB9aROqRQZCgHWbi+9sG62ayYeRX+RzYrKXG1mF4QDm
7iLnBwsMw3mjY8TGOduowrDM/IRxrn64SuGJJjkwl5pKcUln/9ci5omIY0kMEK3nnqfc3ikeU5nu
1GqvIJpFCp5rQPt4SbbE1p08v1OJAqq2hfnLlZ3GObDdOhLQwaoHZMvs9aUa+EzVjk3nfJCttSsd
nSrJjOHQ3w5wbnc4L/cwANP/n+fAwyQilqiQXCmXVZzW/ZIO9vxPYacpBNZm9CByqiq6TyQVCgAU
92GqSBYUi+N6oyszfwFLY2BD/Dx9eGgYqvovufIl+p+qFlapZ7vIiCt2dR3xFF8TCoKJ5HJchwn6
CNCfhGBG7/1jf35+4wITECe33pe77Mkml0+cXr/mcJOi6gD+XP95SiCyz5ND1XN/ayZL7C/BliI+
wpuSJcCdH6ghQLOO7bywz5GRnYh9sJTgdxCvDi17i/zDnrSiA19yxIFbt5BIvoIgK82wwdhKCvPm
F0CJiTR1lFO6IeAnE8XPoaDR67qTqUAc7wAT3TmYsdi6zMvWTL0PaSTxO8snYGt6IHaYb5P5WF7A
HQtqSrVaWxNRSzAeKNGs9jbpEyn8NV9tkmkn83CB40WNe5IYM025xd+exyFOahfbvnv6/egZcAdM
qSoSInY44FDpZWdGL/8p7hGhQzmiJKo0l+u4QIThQgpRdEkgP4Nk3RGzPCuF2VMaAItxGjcrOoxO
EjzyFAnnwW3pXUgNBcMVFchkGDh0TAS8iigWMeRx40/vIV79bkf5NnxC8T9L8WdA+mt6u+MMclPE
P51aMAOhOPdA4zv/ORciRRnccbdin7yGtRCtTKQveqN+DHmciT53v4qIZfvH9BNhi05GJvbQyqIz
OGE7NlgGl18C3Pxc8WkdUAn+vK6fMz+E77SARFiCJkWfVjludMJCtaoCMcLXtCzA0lEGwQ/HgDS7
cAfMhF1PpGx/XEkw1ZjCASh3zipzCH1O8Idpxp7eLWrS7ZCd/z3MMDMRNSr5PWjl2f2HUrD6+Z/I
OcUUoYXHAdw32LiYEFEti5V44/T/g8DNzIplHRiknHVE6rwncyTnUGvakA9CV8mtmGpoEKltbqny
IoLZgRBZUUS3pLsrpFD7U7UMt27OD51kYoOLlqdSsrqNUmuvc+4p+AHibzCHV3b8JUEcEEF7novm
b4w1z5+5tYZYdTXJlQRg1YMGCPMA4D3ZMSVEN621XUUxkMf+PolSq2jd1hvYRxVFrA7Kwv7qTlY4
kcBrtqVr1m5VbGjvLRprX7a1+Q6VCAJOZeaWc1gu0Nz3Oz8ztosu6SFZJiYEj6JC9zyYFEXLy7s2
RaOR+tgeP4FEbEoNqhilYPmEglQMMDPIeLSVi9l1Z40fHTavB0auTkJ1wLkADZVkCZkf8cPvv8qm
qAEfgqkxZhx56AMVMj2BUNvC4z/8O8ExehhW+vzrLJNwII/rFn/QppMKJ1lJmWAqWRRhtOpKcp7t
wonXoDGBySD9faegtmgfH3R6dBrTCaTKZUNIgiOKP4Yj21bAwoQuQuSkpEuZ0yFNu+sbbs3k3N25
2jLepv/SRy+C4leX27C+bVbzw8czFXlhfOY1jzIpfdUsdFaMuR1gfqilMFsLEb33rQqRdVG9dq6F
lRO+9ig4/UyRayBufdUHhxHQ9/MJV/kr6NTdagIy4SinM7In5OklDZvk6sIjT+kvlZAnEaQT2etu
FldD8F5iKa0pAvTHhahGTACqXBKvjbhrhWGy2arolAgi3j/J0DqgxwJMzKypcXUz8Vka83JwxTlx
9fWGNfvvgwYb7eF6oKuvkH0Z9Sc7C4kyS9yCD28+h4/KzqkD13dHxq1jeRlFqQzB9W3UBrdyZo1b
n6N4Yjk9ENAUFxTuyLbgo6cKA7tCWz5UklgtbM6bN1xCucWzdHVw/T+HLDkH6ow2YLRvLTVXNU9U
mwXF/oHoWWFvpmKzuDVDWUfLDryDnJfzB5kF0cvFnBneii17SjE/mGlwT0nbGCcamcPOvNjqeXfL
QHBBP4MZ2LJnvNz01MngRzHzNvy4smu7ZxmMLG+IyGHy1bdWa+BijBw0JghZDoGnekdSGc5UFiap
xr51JfMxgPpncDiRMqFATrzIbUqyYEnNY8q/8gysFFTCYSqbXV4JjvJg+ooJKSt5lRLwyF01eq/v
SN5SD2Nexfu4My3KeKUTOwy625rSbzslJB+puuQR+aacBoDGckAemyTXcbzRnlGv0FDTVcxkMeDC
pWJW4wc7n+6lT4XKGqSLpKyxCicW01dB1gPrNNLRjt8blwCjmHVLxxI46E4wPe0TAo81znw9HnXO
Fi+bHZMMOc0LSMyOvOIBcEGxAIzGszhKbkWm+0sy6BstJQEzDrz2sB2Z9PRNWWiMqUBOYOunCHR0
GonbOIY2Y1ZNohACVCujE7QVKh+YzeZ90D9DXk1ClCW/pcjo89MP2XtQtV6aYImKElNYYwGveSzz
7BuiXu5ADQjc+IuGuigqWQTitQxgdFaDi3EBRUSNnClwp513wfEzKYSh3JImLSeXuw/zTw35THzb
S7N72JvI3bTuUfR54MVL/DFYgPElzxE4JWskakvk1OWwKEX/Oq2kNKANF+pOri7qWjV5I6bap1TC
mFupxosdF5c1xXoCATHgT+W/Mxr/WfUMVkSingDuSm2Ig9TrtLPs2673skGaK/lqQoIvJNqS2KVq
uur1rk4Go0zh+7PImt2jsNWwhdED/hOcdG1Ep1yCDgZKQyztG4TWUmmIrel7TOly7mEK7oq0J292
Xb0m9Tiaj+pl+C4k2YMzCc2QcHWX0beh3M3TuLdVHioV9osspltYaRdxAXAuYvvTza8wwjSD8orf
Y8SS1rjQ/CuiY8H1Wz35A1Oznisl6mh1qNOyKBAOnw95a6kDSYqaiaGk73TNdjF03AdP2w00vTQX
gBkkiBCagveqT402Etv4sQ3uA+TeXSZ0OwHcHVZGoWaHcJlVIxeF3Sp8QUwVajZWVFj/e1JN0OIp
3ZdbZID11jhgM+X4xhROrSShT8qKsi5eBaNd3ijfIfVQL3g87weBfJ7EGu+o0pRGKLZMnm2FXO7w
UPRoLlEnDCwJquSHgeaD5itWWqp6okZ1G9fy1uksYZarFVyHgfsnZtotJsHRQxJSBdEX8dQKktxv
5WIM8bqTCcxnGt/xDfiQPdqJ6VAOlqdu0JUfPJOA33kIYp+iyyb4g3O1TmXhf76pZnlcDYl+CrAU
n2r7EPdazKJSeCc1UE2d6HRy6DCHU1a9JrPqiiXMorl0BdiMdaFPyMchNheHzv0D/FDoy8IOP0Mx
K8WQqg1jyRuKsOZGTfFqZH9YHb9ojUzH6YcfpBV3QVg5NXHboHb4QAA+7mpgk/KPi8/F7/VSayTI
IiTH5viVbmysUBSCRPs1d4x7xM98v9M59Of1CD6enaL4S5rxkrfDE+XW1KLFWzePRZc0R103qu1E
h5goO6QjLPQLAzrwSEUc1qRjRsk3kiiufB7zxdQslUW5mxy7bgOVQ2ksXgXntEZ0u8xZisENsI8h
gpse53RqSDgCCDlAOA6zsEVVQDyQPBtSA0pEt0f7zWPCvZOupWNbygxa9kK6UAOn/F3ovX3jhnQG
I+457vI18HKRo7MHUk6Ec+bBwBbevPrElfdMyar8lFzBimVFm/c3ANN50jOimmuIGOuYqRD3N3fk
Kwq4ZhQBvaXiS5gdh+2ucW6fCL+kpIvGBqKB/t0UqOvd6hW12mY9nUoh77Ra60MOAU4Xy5ARajzc
uaGOnTU5XMBiJV1tnz7m8AtaxSRE36o9xsiEuEnutzgp1EM9wop1qmVf+4feJFjytIwTnoXGjgsw
8fPW5EKxPx9E5QGDLU/r8dJZzvZ6Vd1Zjc/hpLyS606CXWOWOSfOK3lGV0RWq9J7TEVcy35uW3O5
UtwWUVJ2WLEi8aEkZsIrBfM9k+XGzwwv7UwarJji02k9LNnKu9Q66UqfQ/kqAQj5vQW5Qc2A59MV
M3PNJJlZj150yXf1k1DjLPquSHJInBjWnC8nD8kqrOUAsO6DgRxCtZGhGIsyM9F+POn1D8mGlqaJ
cLj1fHLLiL4GF4R/3dXyYj/Kr+4br37Y7FK+/fi74qIXag++NZGVdGhpiyr5gqYwon41OzuOnC9N
UGNqVgF/nRq78rZWUyAWjPaCIiuzsjTMA5HS8S0smgh18GgA/8BG0Ok6YxItKM7kSsjEQl8pTpLX
vqxMqJwFFeniLwEjqalrGH/xavjRvORflXQJmpDMvAHzD6oCu+vRmtCRWtNahxQJ9hrNu8dc1x8o
0X8z7VUrzoL7JflM5lIVBggdsBqrlmFdwRjA8eI9aLFPVWq1603hTZSStC2EIyIyxQGPSUI1tnhU
lMgzX1CdrgJhXOE3qGCvYLzepuBhK+fBCNaI9DJH+IEDldQkH+u2abGofkDYjiYMrY+8fQWpOfjI
O8+Y1z9Y95WcOt+sVM2o2S5QoTjhCm86Ik1vknb4hXeXa4CwcoGo1S9aNkg/nA3PXH+mA8zavRD6
vPg8wGDwHOcFnBBrNUJMSuqATId2GEEDrODlyBw967H7Wn3fPc+A/vu12WQEfP/okfHEI9lYpAkS
S+uWx2ds7Vt14jrdl6xFM6XyqK/6dprQsWT3tJiXQmVmBeo+6YWotmRvRBKPfcKJMjlL5Bypdtxz
CTj/c3p9rYov2c/nvJL5D4J0gdwkAHWdG8e+Mp3F5KERHVYDK++BlBU3JmRLXryorLYjqcpuCIA+
r0YTUi8umBVD7x0dYPEs9sarFd0cUfe5lMo9PR6cxclBBVC6QUEGPr8u376nL75OrYq+psyRI0KC
0hIH162/Z8odMR5wKgm5/9tctCjOxwmSwI657xfy0dAvwCRWsTsI24llQgoserZ7WLAT9W5IvhHt
xj3IZdpV9Tzjd7XXYPrK04k/lPdPVpChAKa2KyEoZ8rIono2hJl1wCtFxU3fLFiUvsp/RJEKvFmh
RaJPzIEAGmonfVsf7+jIGjRR5Edacwm9nBrAWzRnkGLQ2ez/KTpXgyncjxcMoLycP1WEfJ8R1klo
IYPSJG7NblMEansd0ifmw4hsQIqe2oaz+C20JHvKG4OfRbF38gkpq7dsoXwTPkKxzy5C9FQU/17f
LX1G0sRyIrEbIJQyAwNyXpULMPC7VuW9iOOntVLajhj88mbyp7ryynrd87z53dRi5+wxyvEPDLzF
P7YW7E4L8/7GIcF+htLnrH8lE6aM6t016Gg8l5xL/gkiYCmgGHjUnaXz/EoEw3BZyycq5L5EGKrS
HQAXtUybztc+sB8UeVRFZCmSdicxQnDelBHnWlEvh0TAU2NE+UMXlu2oPTsee1P/ZbWSbXLWQHSF
qaU5suYkplzymqJ3bjKvxghJbVyyM5akXjCoI2AfcGc6KPz5YDsml58vmMDBoyTWtqzWjh9pHFrw
ltZLNks/bwOeqz2pbhKz/fpx7gdv/YOuUVW5jWXYW1qO606/dFLMrpMCZ8S5wHNUOtem+2SY6yEI
nzJOR5r3QKitjYy/aT+mcZlDZUcMMf91I4Ea9WLJjksNkHFcTy/686o0JrgbkTbDdL9BpF7CZVIq
Hb7egr5a6gF6Avxx3Sx260F91dyY420JWKDz9L90MEvSAu+fAyOOCMCPf6pvNgMd4dQwy9Cuwq5K
cblfhor4oI/ls7d3La265XtApM9K5cHriC5QWhmPScSZwDaU5iNIPeo++MNv+gwc+lIXWDoV/rdG
jHmkffCYVl2sZpHU3CDnNNNyNGTTtqeD4/EAtxilzG7w6OKMrRcXoNuXw0U+8we9j8iAtm9nO0IF
xV2G8HBLr4BT1DxHOfvRb2k/LUTjWB3i4s0ZBR8p+Qr2AQWx3bO/uVdnKI6rTH7AEiVIfb/4yxTr
DI8MArs70256V9xyrhUGnIhncEj1cN4VZakhz7xY7QNDoEm7pO69k8HP+9M6f2Wi8u6osKy2YQ64
iSd0eSVWLFVptSZQM9hx5LgBTFfXwyQc4nsrvQWDydE6mFwqrD+aK8ZDnQIm0eJd2kQUUwH+YEj5
rjEW5ZXH+gn5xmb6KkPBOzgm0KKSqSCUT0Wn5n6n0w0bFHkkuwcdJPsIxX0jM8MOEgyGaiZ8qtku
CZbUiq+GtXnvBYfjuINSBPDArwES1fHkeWzwFHE2O3l3ZhrDoLRmpEPjXVsAcjIJSN0xah+kUman
ad0g6/GdjuQcGQ37xA6OcFNCzWJvjwSsdPA3XJwFAn+WGVEcJWT2iMrkCSFshY8qIIHW3RAgzKHw
DH1D1+/cxS5N79K3hHQmUvG7vA0vBjLwaUGyS2kivU+aE+DO3euszS37CUqg2mC1ejnh2SO8o8vL
x2ni7jccuLpXkr8+EUeRkcMsyQhlavfheWkQakuSkb0GxMXXei+PYJLCJ9z5WNcn96g5f8yWUK5V
0H7BU1/FuUCiNz/hqL1ClyszmSh0UK5XEmvMVO31Pz0CBj9q+8EquuEJF2gD6abUU3Et2eu/toZE
ifsIv/ay0HZiXJMvp1jMN1qaIdKl3jg/B6xJwfmCNLB3AdMOhJ3he6RrGyplJKQUK4Ecf3gIqmB5
MBjucAVa3ZTExP3qrX1nZwy7lqvs2TeL99S0c6Sqf+L9uSOu01q/ThV2LpmLWaA5m0o69d0K5kXS
96pSsNp+O1xBC7gZPF9Lfh6Nvelx/3uBIOpUc4hUwbo/ioDuNpxZEsmkZAZtnCSeNjDWb5Eq1rfC
Am2ERyUntVvzbrByCxcnTDfjZWEm88foPhYyPcGmSwpdmgtwBmaDzXUY0qPsXJ43O5AHTk99RWT+
edtl7HJRkFM98CkuzSCWJP43BWEWKGAjHWYsPnDL6LyXPDcVK1bitPTXJNu6PvZDQXpjwQLWlyO9
UPJluuYN8NeORX33vpzqP1smogLahshPyL6KrcWe0YXnhYgDGgk7giqzYk+YyxkaxS8qW0zORQmR
VXcp09ST9JzibXoIMBbC31ibasROBGJVPhU6fuFYTJRKMowaap5W5R7cpvaLZxaO6xHXX1bmOhRQ
DpZCU4Y82o3cEnoJlG7zmOW1QSal91bYZN0n9xLRgH+noLAj5/DtX7VT0FGH4r0MUH4G0l8VYN73
Y4ShHfU3A0gn9TOKwIPAtxSsINmqZgsIyUZlg9zgTW8F8KBIVxOj8ryYpTev2KW3Ga/PWTBPx8+k
GoHOTan0JAapUo5NBVUjh7TkUlVmP4VhQ2c7+6TgiUjKLrAnH7xquyYuhioOtSKtY8oKG0ppU/nD
nHAMH9XW1GWf+bWx3sJcyv+YJs5vQfryAdUycQTRMjrswFbL99Xd8EunJ9/IRxfFtESOmiBfYw/Z
ugshE4UfZiO5KrmMfprQBoqiPB4LE4JiNn7th8yHiDhMXN3UQjtES2E/XyrufSGuS5oNxHcvAjx2
U4d77q1K2zqsTza86WdWIzFFI15mwqho0fKCbkPFCwKD5iDWDyWliAHkysaH+7CJnc2F6j/uX2xZ
q0kBQEiJIqsBqvSfM+CsEPBtv0x66h1q1ea0ZNyHRq6ciNjBA7DCL3lqXYMGMso3mkYnfbVW3sZA
8ZV2HW9LJoZFKaHhzgvZSI9jJ5c6eLfs1yZyv4n7b6ytp4Ul4o7t4FgOVqRrNBBdEyExT0fQwpfS
rxRJBupxJ3TuR3b4M8uPuV2zLPKF7uqyAwfrW39Y0eeC1jwzoKuoSyIo4qTnY85KZWP2UBswyoXJ
cQIH1oL4aukfMa2EpXRKtdHnY9aXa/AhMcPLEFzAO2D7pr/Orbp+zwIi5N02IRvXlI8L+1I7Z5NQ
CtNeSXdr/ST4cDRz9hF5myk1N0w++kp2p+PfKllqa6vRPd6uyWK6d4LSObYkunIcFqK2BgH4QWXB
BO9NptzXqpAt97XbCZxb1KQiXZ3m8+ApaqIwhfu4IJxFsLFoBBu36EH/4+Oiwwejm9jAuFASeBpV
uVMm3HMfcWqPnKX2PWKOVOMNqvDMVaTV8wO2h4s+sH8gsJfSEegn7Xpm/Vtfu2DMBE7bdU5Lbaaa
DR4kiRiCacv6udRfWYMviTpCN8708UmUIehBpJMVQQ3IP1NvYGkNpV9bmpjZVSMJr4wDA9OLmv2W
6uL7NBtXBIRTigxRrTelzBa54l55qdoyN3MyiggsIYRrl/bwi/aaUBf0ttol8M0k2AP7N0v0rYni
2paGPVfLieKTaXyq+InR/t8NI66ON1LGXU+WXw9X2Njs9YMPZvkSGzN+v5oNC5Ep6kckeRGJ4dGC
6mn2sH863OejPE+qY4serf/yaIdrvHZGwxHtU1mdGXYM1y8p1nMH3zybX3AMeErLaKipUWeamlf8
zfXlOL9xiOiv0s8Kwazhr/3PgBI82TvJ1VqklWk1HErKzzrqq9b9qAy7odK4DbLh+5mV9bfd2pul
qM+eGi81MXf7/U6i4HqHPoA7Bsor17klOmqLhttd50w6MFYt10Tzx2BC0jYkYmlAU9x0vTQOBhCy
TuK4ePyHOmAIIVJR7bWqbqpOdNE9wMkdQSd/QQ8VkaJyvC1muSce/cXTfyR4AnfICXiS/2vmFgZq
9YgcjAvtgG2cKiZvDUxheQZ16vZkcNImuUQkJvAoMFlO45BSv1sBPwYl7yeMEkJX9unqFeS80nt5
FdSTxwA2TnyxERx2oywRkLaQlINV6TtisAc9WbrCclEwntfNd6TA8lpB5aoY3HCogZ4HBNKeeZCn
1+a3xd/uhznnIDrwBWfRAfXdNfPZP06ji8i0WX8lJTzzx6uE9mU2+wNFiMcSPrYyKrFc/a0zDVZU
sEMbDlnh9auxeIo4VtRlYb9QIxb8H9M5qpXxsDGmdH7Z2SRKdsZPBRV5k1S7mCIWwBYbpFLH4fCK
FRYhbifdDWFCWR+fqz12dMWyN/vghR7BtC/EiB3UgLmyY/9K1cBXz8n8IacTnNTvPCCwTmx5/dIB
T/flF0Ma7RFkm3YLfKWMKFFt/PpKp3AgDidqnjx5ZImGYbJtM0+bx45KnkBIb33O2LNhLRF7Gaox
3hBilK1VKbg/6mLQ+m4iZvRYruarJBeZpsz9YAmsc89VyUIcq36I5R9zW+8mOUycUhx67af09FDl
3jWB0fhcpu+ZGQlr+edPxcfyUynKQ72c2fK0ja2YZkzzjGIxu5ODX1e6hgl1BK2ZSDHud9UnXxda
6FU/GTtluaKBGXczBaIcY4ydbQ6XRXv/GjPeAvqfgxr4ZhKQ40RJur99xeW6vqZeYPzQv45ksJ9u
pZUV0cF3UqmKHKclfmNzv0edX7rtWevbyZw266srzaKrkxPlJeLOXFg/Ys0nU88yNW0B82ltlMOZ
KTusaUVIs6aaw9xsvwjZPxAnYgEZeVVIKxFe8RGuCuKFYJ2h1xvvrb//yH1thhr8ydItih22eQ4g
x/On+kxoCoFGnTHzhb9eGzOWkvj1QTVlDueYPYXFGaXE0orj0Q3SUy6KmL6QKQX+D+BGx0sRHZ3/
KCKmYjAHHKkN/XBSCY6veUp2DHi7qmtyt7pWkIOwbVZvembeD46aUOMRaSYWVRA5XClvpNDe/++3
mXKKLzmcCBYKFXilgRrlZzxkVOAVdqTYJrpeId7O508etQIcgXz/iprZd8B7H9NhDpn+ugY2mXSZ
ikWZpvxbR3Qzov6qOTZNb8JkKtFTvEmQ+J8nZgppwOjaH7wqFudt1lpiyMaFASNhagG6d0LcoRfe
p0bm5dOOvUYN2adap5XqbC1e86o5Mrtdt+7oluHcFc32wJ4Nao7zrK69QXudIZH6pPNsY5P6xtrf
1tU8b9qJamGHQymn+j3n3HsHFt8P8CO6S5AHKXIQXJZA+KbAy+PlpWvGDxqe/2QZtMBybNlByin0
uQz/LYSXfW6w4Hn/CX5OVq44QpAITNt4Rb7bG0+uDl4Cj8aJ6z+1aW+D/iOaDKspDAqJhgwvjydC
OJnxNRI6H+gr9yVBUHbnr7e9Q7b9anlr8jPpTEWDBCSh9cFyARTX2sE8s8EvopsZa8SziutZem9Z
tlNwYkKVeJY/4SARd/ig3n9Z8fm78cJ2RfdydAUZu2bW6iUzdCMKVE3TNSPUuq/wOjW/j8zePU+m
cgarmTJC2BsYD9c4/jBFwNbM6vQa53IB9M5LV0aYSq7wYbDL6ymF6QpDw2d+XB5H67BuS4wThppz
JFRpJrNWbs2Ll+UUY+1dlka8AZYqFYHBf+5iMTM1n9qPiCfh0DoYd1HHq69ZVQaH74HK7ktNaN21
Lf7tTW00++1NUF5vmLjla4Q6Q1dAiq33DHJtXCrTbcrvt3pgYV017kMwNsC65rJNaoJNf5+m13JI
tTsQg5+oyn+K/czmpn859OAnnNZqCOq+yy0SBiMraWwqH5VrC3YyVHBwIyStH7jf/m4qEkeQ+SlH
UVHKp1/GtNOEpZTvSbCmk54MVi48FYW/G1U4Tj/474M8pNk90v6SxiTdEPBHy4e8hneeel72CXMs
YCeVTLaYAt16J4VDQOesGBySaRlGmM1Cvrzzbt31GtA50BReLfX5ZanogqYqPFd+GKpYh4YN7Iot
uUBzRue/dWBnyS4Q2Q1nVruRvQt4FS9Z8S3zh4LjF2FM9vA+lZJG7AXQow4bhGZtE1ADqQ/n/Ulr
5Me0/cdVyM3n7qgUe25OFyPr9KK9hm+L/DMtyo3hP+Azb81ak5uYpUGR8I7ige6MPBhO2xyRxIeF
u/psdv3UtYTdzUI64PB4FHAnV7A2sv538aMkx56eb7MeQQ2LXqkde7GZWRwYOV4PR30cDtEKAyjk
Zsnx7buSXJ7fz/7G6FCtcaeEnvlhQFsR9ZsFP9geiSXj+l4Q1/gj6eCtHhGdy4Xx3qlfk/6Hc8yA
/1uYVeNIogrVDq53ym1oEkzm4b9joETuP8moilSpmooZdoN9IGDa7h7/9nclnVXbZFWNftaZP5Jo
xuEnkR9p83R0PPHGA+rl+AT7VnD+jqfz1RpYTTLWuOjUtrMVPjcYonVe7bR7BdwEbVrAgZD0FCyn
dWrOtn2XxbcyLGUAUgicGLl0mlW2Kdogy63v2wBHI/kArSZ36usbA0hZ9KsryIV9k0mj6Xr3ZeWh
3m3THP/KK9s6I6LnHle29UElGt922PE3EiN+FsvSOr+BV3Caxt0jlKomeGJK+ZAONmBSUCdlwbSI
lS57hTcHgNoYp8Q2aYbP7uCnnwZthyMHBM+EEUZ46DGGLNDfLKu7DnwvvL5FSLoyW9Ga0Z/yYHaL
nngO3BOeSl042jHEQifgRiOhr8KzVjT78e9RbeCm3w/utQU9Hf9JVxpn4OoAU1Hz3mbriPtbiXyR
cSm+5IOXdBBJjxrz5KIHaCwSwP1rz6RF7WDbhoZh4SSvD8QJ4pk/Q5E6XGfL5kdya3qa1vYuosTT
XN62X8Leh+HblXpq2887dXEXFuXbT/116TxUhtALAQPO6kbBW3N+NY5+t6gmqpY2r9ZMQTTGoF57
UaIu8q1aW9+5X9fA5q+WHC973w8aOslpDFc095eLqPh5oFxnFBmJGbFNyjqwpkM/Kx7TwWBuXK3G
IMfzDP8swN5K73pubtJdjy2PWq+CSsTt0TlNnfWTS6mIG9qS6qONUa5ho3MwzqLpMd5zme4Jq7KD
xYICnwo4jcS90QVmk+t4mlYwJdyE7W1WYgP0T7omNiCCUSiYXn42Ow7mbwFWwSyG7SLpUpDOyU9b
3TjSbFFUKPATvsek10vQlsHE37CS8yel7AATFQ4gnOq2x/zLgIFZMVzjVF4snVBLg1IhKpne7kYX
TsmHyTx93IIfZwr/W5+MdiUlVd3/7qaATqsLCN8VL3r2/KLoIJGQlotOAg+l2nr1OLdDcNgHB/5U
U/cw2jVbmjB+Xhu3UFgEsYUhpctZ9Dhnf9aQy1NcoJkfRcboSw1/tzVw66REAqDUybJzFfzUGjxF
IUp+BNRq1HU9SO3n1eWeIpF2hr5Ahrsk2tykKN5/U/TVrGmgkB45MkcjPiDzdQpQdBXWMM8cEJdm
EysNlfCdabsnavMCeKDKKTeYZfX5QaQY2K8yrDzdwnl9AqVXzjq8P1F+SDfW2xYVKyWvV+CQCiOG
ouE0+VfwZ674ZHnuKzEzLZAtsVV7dgAAlPcET5Sc9VBPJqivzXN4ioeDlNBDkWozU1KMyv/QGtS7
CNZHPri7Op1+zNr/qUusqrTnajNd/+ApAU9Yp2YSIuZVdTjmd5Q3H4Pch0zyNQh1B6MqnD/XzLBv
2CgSOfVqXwdvKgWqThlDdYhbtA96s1P7Jyz0H6IOG1/XkRrKth34ibHb+0XRnhQQFrBBCaJ2yTqm
s0kbMLbN+g0TagsowMYq7B4WQyxeabtsuuXsD44cAcbmke2G4tKGsU6sBMFOCFM/yRxGVcDysSD2
ki5cvcegonFO32/4/SIkhKgwIVJcq20bz5eeMfRhv09UXj50ewsL8Bg3s+AfVUqWr1DKr8aMLWIt
n4T/pK3nGVW90oSXOtHIGzmR7H9e0GmZC/G21sXtyLJdiHiGxGBIOVCZowlP9ef9Z5GeRIpDq2Ee
SrAD5Ow8EgSOZROOLO2XaKAa9DpWr2RUjF5JUL2/7OQ0S5sHsqLtMfeIcO5lbAWjMzuSG3t8WUb7
yLA8yL+We9O3XMZK6EeE/TUFe9QVcZ0JwbZJF8djCCO26IEPh1UgfHs0RIW0pY2on3HGp3kPKaVk
f4shcC0oBamOtHIK1jdQ3trcQ20sWjY67eyn18+jNB6XYiKgF5t/Tr+aHxp8d9xP5NJx7v5cIyHN
8jUGTxprhPQ/gJN34+fNGiC83G99vVyZETzToSj6VeKS8EXlmKjngZ3/Oc+eNVdqXsWO3FBZE93R
OJk7K7ARTS9DtjJyaaFDAjZTADKxl5Qv7v4f9rGI6izPDZ6UIgitZBsZQLsY34BPGK7n36sYrHAq
2I/aKOnDr7C5zwibXe86kG67MdT2DWM6bBz2aYTyddNPJvUwWMdwPxsIs4Wz06LNy3Pk61hlRW0Y
TOLGxR/3WyA9SjZrnVb0QR5RDfMC7du2+hHSNHk3JoWov+Ykydb8snzNQskyuUG/tMls9QZbZOTG
vIQDBmxCMTtfOK+UmYSz1SQoV5OGONdBhyi6PAkIMJjlmTxCxn5Cpn0/nm0sW59YyUFFRnwxRfdo
HqmVVMwPl2u153Rl6XY+ehEj4HE0pEH1z9rFy18dW3z9u5yqkpUbLP1yQd2k1iSJaf72kYXQkjGZ
RMpjNJl9xE0xw45gq0pwXBQ1ECoJV8tVCcfmSi8qQrrKEDbYJLYcQ7iqlAWry/OW0azS+CdP8Krt
Ko4Y8WAVeSSkcNZK8PQul8+QJfP9kQSr4hH4zQZ2rTxW0uYwSwj8q1bSqp9j39irWozoAaS575dQ
aJ20GOx7zR2tNXx4xsimdQMZ4weGbX0k4xM4KpS7uOI/ytGtw0wfg0fUkl1Gw45eRZyWbaYcB7Cr
j9y8WomhPPeIjVBe/JMDy73LNu7DApbz9AUK1qDiaxGf1NCRstgfoUuLwe4PxYqX23xwjTjnSbHv
tYswUBbxRwmk89mspCbi5RTZhDWzDCqD/ZxKRMPtDlWv8dOVva6Vv4Vo10qagtWVM6V30uknpIu1
XKcJy0Y5VE3NGiScqdYTWxLtbrQBRrwbzaXF8i804awGMrvxnPB8735Jj+Q1KYNc8Uv1nnoLp5kv
3btQkCuzk8+oDHJQc+awrmiDA+vUGH46POm6zGU52RJbLX2YPQWNf2nLHZrgfw7fZpDA8+RJ6ESt
rtTKgE1D141sI6y3GL6a/XqxEk533exLG9XNHnXWnPRmKS0YZbMFFzchO4NOd33xHhnoqwVyrEPy
J3cB/2mC19Hd8FxYkGgXRlpqAY2V2L1RqtPvzonuisap65DclOT+/UTWkpGZTfkIGy7/E0Fb1xcT
2CNGvxQBph+/9H+HRPPCq1ylM3CxIKS+zSWxr3GUfrqpj0tA21MfuGWfdEHS917JliR36BGWDKma
JwySUurLyCFN0Piq11QmHL6lqVyEPe5S5pXn+sZE1Ul29NrX4J7Wt8zl4WlJ0i6uNV3qOBrWSZjD
M+y8yrbejzqKQ1Z23TboRhT7yNiBZn6m/qH0GoNqP8DEDzSOFnBAHI4YjLslpyk5YDMNn/Ynt1Tr
ElOzUNQRVFSpvhBpa7PizpNkFE1AaPTGR/QfIA61a8QY3x/0tz1bKO7kw2Fky0w43wX5Y7KQ8XbZ
IihhsMPNP5V+wnRbWInm1JmulLCao3IJT2SS5QKKLKN26GdyzvJCgkn1qdBAOJQSNxvaNJS0F2mq
pug/WVlHDp8wY03wtsV7nm3ibX5h7/jZcgMYIYBRGbU3btayCJB13tF/jqc3nW++gh8K6AFyUSWT
l3eX8bm7dVXWRH52cYzE9GGfua/tDr31aoXwrUrMrj6xPbnqrfIbVmfFCln4MrzXifw5nmHjcWfx
/vbD43QKhGLJ16I3/IG4Ewp6GrzwYLjXghSAQIm4frh5ey8IQRUT2a5Ty7BQG+2vWPvvAExQFJh0
CA/cML8JSHJyQZFF4JISXklrJPGV6VxsLgbDaY21+vdH9H9JanuzwM9mHK52yWWQ3HAVwGWuT5lC
s8vr/yov1pWY9/ik4ib5/D9TRnsVsRGG0MXbfxyRfLQtn3NQ884e/o6wnbLH9evWkOQ6e3w30VqN
ry76PmdusXWV9wUifE4nhSmQKUf+m/Dl3DX9M75Q9CIz/h/6LGMtxAlkNlTWL4UzGVjnNvxr157o
/lahYt6pRqFLcVrqtfVFPk9/bItyLgZKS0j01jMqVPijPpArs3vC1XPMPjvJPcNEmgIQEkltD8Fz
LTWfIoqFXBtOXF1lredHzCYrclcKgx/kKbdrhl80Zq6nMvTw/PcutLNilmvb21E0DS1dxhlyYGDb
2Ger43xBAA51qDvMng7v6lBL4Zw1Ji3Jo4w3o3kKtJ/D8Z2hOFHnDrIh8RLP90y1FqmEidJy7ZYC
h8tdXbUKcKexHlS+1zBnmQbs/z86gDFVWywNmfdQXKl9eZIik2oxFDshzIYo0tpm7GiS2fy8YKrm
5e7YV+hmppurDBBxScO3y7mnBMy2//8Y9lZ/iko1ww5eTTodGWi8nY0s/9ZdVyVH3zSzySc6EG2z
EyxgKtuan0OYpZHyWXBrk6NivLyINzWMX/bM4wVcip7qe8NIVJZEJmb04O6Ex71qW9PlQ/i0wp4G
AuDx+ipunJntstS4zZe5ltexXXCfA4OXnzz0Ra4UQEKYwCj1dFV2IotQt0vKCoDV4XvuEoh5tPwz
yrqPO/2AP00inwklZdmXta/s/FOU5fCfYASVHvj0r600vOVP4dzxV+czV3OxeIw7cTk3qPOBJnNC
/5HDPNLARaAcksSwU3AYUG4aM91zX37ghpQVwp2m8OeUoOnsAaxo7hdzySV+4OwmBzzQOFYcb5UH
XElw/TlkjbzXWoz2zdZWNGJpnaxpV5Y3AI0cdovKYHrugkPoxxHcwzTq98hCxdvgp7l6EggCrWp5
CzYHEJEgMeoJTp8lNNTY9kfl8iHo5G8lpS7JEjuVmKTipoEnCdzxs36XfhGgSIYarpYS+lypiwkH
nVIOCY/dpdLcVv0032IYMmKdT/KI+xO2ALYOe5IZdy2U+xVLBkvgGJlGBxW6allWtUiGVAoDjmgh
7uUfDsMSaJ7wtG9lbfLFZ4x9EVpsfH8D5/auSXuprNdo5QoQc14nbX5oJfNd9iIKoRwH7i3TMpmx
CxsbBwzlsThaTG58L25g2WlA+8gXYmbbSZqNnlbrosampl7H7RGcf8gG6np+/hEO4FNDDIxaFXWS
ELe00TNbLH1wLrULaQB3SSHe2X3jSlomxrxytu6+VHRtusTN9MTWZy2iFprA2N+HoYyi7VmSQKGq
a7uT4SvyX5j/dzekk84+WNeg/Di+m2PKH6W33hysiP4iKlYM2UDpfHIDxUgn4PAvv2AKA0DhR9RP
Z2B0saTA5K6itS3Sipz09gcPteFzQzHhG+HgNCV/XonIUuiWvv5JPlBrSGTt1xPKyZsVUUmy29rS
gdqpXaMNCTULLHH6umdDzZOFV5DvD/OGfd2rejgju3/tQ2evbzXyAfG3a44g0rUIsazM+eWCGc2S
TqPpXO7WaGQ0BQ+bvhhVUNdCxeWJX0BxSN8jrsuiFIV7PioQkdxg4mBSaglWUFuRB7ILtIDTsgQD
rKtrzo18h7kbbVK1CAG5uTAty3keCUb21BVMYJa6dv2LMN9kgPG/OjAQZGy2IIbkGwDxHBzqpjrW
xTCcZwKtogidx6Hli1KHouqwD+JBNFvFjdtjcavgzXt/m3nQWGihzF8qVyCQw9rsUFBcGTniOZQf
mr540SWZwuNizNQwlXRtGtb8+gTXc5kntRKRZ+rQao7x7DXa9speJeOXdrEQyzf4XYsIN1C6jzZQ
Dz9/2+bMdKHpacvljGHMTU1XS1ohMTKjcNqa6nz8l0hHq6Yqz+QMojRoaSgl9toTtJy64OqQae61
T/eUuxariN4cfI52kGz+9XYqGRSx3eSgkQAmNY9O++GzRyJHZTJ77MUGGa6j+Uc3v8vhQu8XjOv4
rWWOwvhDhYosrgs7DXkBiIkuR96P8Ihxx1dDcHNaI3MKFJK6SE9UF8unw9wgRKlxEMi61mIkJBe8
nqfZ4NiYJ19rnhcG73ML4tAy6Vx/dtRaB0RAlV6ZCEbJJwB1RNME22YP7rqdHw6iVmTmwsdgOcmt
55Qon177dhNRIp1+gqr2EVnBNZjoJd3t++8I7Ouwbj7kC/5Cx2/BCW+gjNw6InzMEY2pWJn6w6jw
l4Y4WVmBx4CWOwPlkYYOAKz5EjGFW8uAtvXouIzfETXLxJNMI/0HvmhQIWapFl5UG00On9OKmFE8
D9sgud2iI2uMf4UdEHxwi/5v0h8uiadxmb1gPO7Pq9mgSLrSs7xyRENKwzAEedxXNck9Sd28AjQF
AWgpbNzbo3MT3s+klhucg6bmSq92/j/lfgXB11YjHYHcY4fKXbAsGH5kKjIuBNO4rHg7iE5ht6ei
r942Fr272HCILceLLahhdKG1zx6r3wYryvBGHCSn0UYiqfn7vIj2uh/bTgG7M8yaubm12YV4VFyE
JJ19xntrWdsD9pw5lkcpKtWE+fBZPgPRhItZKGFzwNpKiUkvVZU64zi809Serbj91yyVfYHkt18M
fIQxVlGpG639250tkzhmIpk3Lq4tEWUSI6Psv+mF7bU8Yk3yWHmw4Cd3/oSlqnCPRjXB0hNpPUOK
Ad4QkbCijNFUKhxWIW81aVoIJhX1jN0T5Ws7IG1xEkSOIFDvbROhCOsWaQFZz5c+Tk3q4c5qfErj
vT+vX9fOk3cFTiHi+dT7beOPsN9O6j1sA7sv3GfGfsE3fdzpi/r1n/Mtko/QyQdEbepp3730nCpM
QokokPEMAAMZcBFGGqrWithptWBRzzDCrUIlzr6c4ogcRMUPN0LnKbOdvRbTpDAghCVRMGtvYUa6
b2nbWhgdSM/bpDldpGt+WVii5U7h0HnDCR24S7voT3FNsS/x+xUV3GAG2sSLwOsYEOhNKmzhvFhz
dDg3pCATMhv8UAgp0tb26r3UQbXSTLWpE0JkBRNtMLDVor14KWmkics5LQ+HFKcueb5xXbrDZvC9
76JhGcqVKLn/+9hMNJnju5tUobSYzu1FSA1S2852n8CGnePIa01bDMPxkEYZvfTy6zB5iqRYqWeE
JoZjA6ufPRd9lV+ccwyBnmozU58hveTwpLfzn1mY62hhlXd321uBp4G2eo3AwFYvT2WjbhMBciMa
cn3q/wmSV9FhWH1XrCIogdWDo00QlyXcS4U9uvokFQ0hwowIHVJYg7n86jNapeX+hLeH8AV6bNKD
GgvW1B3rBqBctykrJbmRv5ES28pcEFK99si9VaJ7/zlSM9peTeqkrSggSK4p2dkIDuoLFhfvB6TH
NxUjQ30iuFl7sQaHWoLYgaN5x5gyNhtNdZvCqrqd+TiiqN0OJBF62+ZQXDGYt6dPKAv6fXvGouE2
hclFIhK8obuGq1TxU/WKOxMxyc2ZYofnha/AsF8+g6J4thZQnN7JUsdKThke7U6K4tgPQvDmrfVr
QujGC5u6VdGWJKKDBxaKp7dqdKTZXVN0LI2qhsX4KTDMCw7JZoJTUFxx64owqWueDd1jGjdSOnWt
xH2nSE8LL9JhILxROUDUAi3wuhNFVPQA1W48OGVPWyNFx8mU7MBNN3yytlHhLNj4za47ij/eLw3k
yXRfdmwBNint8nhGnTiOsJSc8bhh1eFmktjekMG0TtH+pP4KXv5MUQej6pCj0VrOY0aWV48yVMUu
HhudIN3oCvxtkcTy3YFhPO4w5i15irNRx2gzF3w+flqtLd+iN0G0uN4K/HGEiz982uClCLz2TElX
P0QSpSMZMeXaLsQCjg4ExI1Q9LPv9Mumy6LSvz42+5MldFtvx2nsTOwX64RwP+TS6KAsy23TzaeI
iLEWlsi5CD5B6koAFKrlwQvpxwK8evtq7mxHUl2RSHl6z0dWSyFI0irL6Mt/Are2gpVySmMf+isk
pd8xuk8ZC1In+6/9wYJxmO3f2jXqu2Hz7j1m8i8y1mtvGaEXIeqEsvTnQegedlTdM6M/+3dipWgu
WkZlBqgaEG2L0jNbCeykxWlVARyzYNl77vXif+KWJEeERebXdn4sfp7O3Aui5llkn0HvdcxAFC/2
v6GqqX9h5pS/zSH0kIbtEmUIn2cp0GAcPGbmqZJ5p5LpCD46lkKeiP3zEd81XetR/zSg9p6X1UeB
L7/Rxbhbk7zrxucS3OlV/Nuogzalgh1o6V3P9t3v4mWwRyZ8ynp8QNZEufosaPOyeAk3M0SZ0X94
opDdXNvYfsJBFpfMMJN7CNKBv3rPx1nFq5N3fGZpRdPKlv6j02kK5OYjSJYfNdznmV6T1a1J2kGc
UfwBNzca/xl9v/P5oxqubjy83aoOsTv2l75F5z/VB1/ufnK6j7wGo2MEHe2kPk3C5gVZt9jfwsl+
jQCP8hNCyFq0tYGUdl8/TzUv5aBpa8vYayaDm4VpOBQ3DEfla4EyICyVWhtcEJ2zE5QcQTFASfrO
AqqV8GjfdqcbT+mnuVb5oUEJzjpabG5gNWfVURHegif5YfRskroXXKtVZvOUJLZeHuwRcG6OklX8
yFMJqpKoCUTXJaogWc0mHOOHfZ9ohnPEoGA1IagS8qaT12MHPSff8+Wnp8m23Z/oXxyC0Lsp5Ywc
JgBR0LwEkAkjBbuDBQvyNGi43y5G4UNji8XuFYRXlJNCpL7egYd2K6S0aQJAV2tKaCFdjQIpbvC8
UFsI4d6Z5foCaLwUhuPXTTfHN7ZgVAcGKFCteQhfrvZ2Vap0eVTVeVbabnINdQ1TvgfPbji1EywM
DnQ0wMTfjqo6BwM1GTcgz3liO9vhMYPZV9ruQHikzT7d2TiIiaKDZ5FQgtQagIppOoo0NKSSin1t
0QsdX21psmI3//q38vID5CIz0bpL1SMYOq5El28GauOo3eBT25pnbPpWxmmWWF8B0iO9oG6jn7oY
uFys8P2ASrR3bH/qHkG5wbSyw6NU2nM5hrY5ji8Ia+nlrEHvSMtwhCiNrK3GB1yitPdw7boBLXlD
59Qei01TdyGFEzLPMWPWt6f3Zwbjqs/rDoCCPeBqKJRTa3tdZ+75D/SgaRXiPXwcxWqmoU7wWBYk
kfCKjeGftP2r46c5mR1I5fnVCoyoOc5FpNtHdqWwJTXdGlK65x205u1HJRdngbXXHKRDDx5V86G0
FULhg34wyt3phWfqTTrYvMrc4IDn1OUh0o5yKeNomv51pOjtPGm1gUuAyQQfrKGkh9HcRRWSaUL1
eUbUOC/pYb2vsumOI2NPtyWwaYWM7I/fjJiLkoZogFQLZnnjKftrzbgbqZAeeYvzStL2wO/JjSQ5
iW979MU/0Nk3N5lAQ7/ZBc3nCbtI2yKxAV+4TkbHzKy5fpHtRZ2caQCGKm7UaoXlw9BvlPYvlwoR
C964LScEFHlmVKkQvUin3xuI7bGGjllX4cXG5mWpY1gVUrQygoJqd5VIUhb6LnBge5Qy2SrbATBL
GQe5V7GRXLbgsFV1GFxWYR0aOIIpd+P9fGEAdFJ9rEHGY9iMCxskZOCpqAiX6iqDZ3NsuIMN5dvs
mMtSspQQ5N7NUHua3vze18uZxLrYa5Xb7sy3PGm1w6j/572ZXOAj5Zar41dVvrIV7ISsTScRd3LZ
TB5w4Onlqo01z6pSULoMKsXCX18KBIppUX16y/7KrcaPxnGh1GSBFdz1YKPe0lfzkxASgeQNGCOP
p4RGFJMFOJJbU3+yjLCTTvNapzy8sASQjGgfY/9xGvzwY2oVWd6TCotZORGnsglv4eowsQaTzaDf
qTKv+rkBngiM/+8PS7DE2tnj2kSWHByLg0Jkiv/Al1RrQiSDrCpEND4cxF1RsCJx5UVQHClpYuaP
z6ijnrtH4lW2+gsrxUzbKtEXz+YxClCikbEJrqEOtRzROSqJKD3Q8nAhdutRLDQ6qElegrNEtl7N
0LQd7yHdtIimHby/G2iDC+KiwcYiq3lSCmqr2ZoH3RF8CN62lBI4HbDIXJXq3GES+bvw7GTs8VKk
PwJY5Vi03saEBWexq7cAJwgwF6D+5+CKN9lr5dP29bQU8bXIn5ic6Kd4THaWBSwnljNo4HlZSodz
cY30fgjKxgcUAikcPytMmjaVIjh5eTHn6xqitH6nS08CY094Ai8PWl8jPdtaTA33RdR41J8aWRjr
HQH6qhj9/JV3P4AQJWN/m6mHefygrnfGo97gyHW7u8UgyD2aTeXwHKwB+FghEdkKBxnxuUM0KQSj
BA/q8iT9pdS+/qhX58ya5w/LlBuL6gwdtGsFjxA3XO4qA10kCUsIbrBtVPtL3nx3ziLf/wVZCBlY
NwAfTF+GCElcJp3xfV5C0jWoR/R9TMvsHBvKD318GgEKUJSMWTZ73BBahsAuWOcdTj5G0nHl+UhG
LNHskjlgq8KTOF/rxOuCH6Mq5CS7PHPeHwYZBOoaFieWNvyNGCM8TVHoFG7N5OEJ3rfh2qNojP/8
HYSJeOZsLpsrVGNUjGzlizO0H6rwf+g1rrVSJXJZHZ5k+cVww5m6rdJ6yQ6lUAbWuayuJkGkbVl7
nvl+H10PVfxQWgs2pBtSaE8IOFJn+XzgAcBDa6Nvtof0EMs+e1LrI73UFLxsJ8Z1YC/zsX4yPA1A
f3m3w4hmTymjlguKKxeLDAp2/MCA5APwaWoq6MGxpXkOPHUpImVfyFgZkbCnZKwnOesRumezU7y/
Ll1NEy8vUmjm4EycLJTCfbait+lpSe/SEwxxejRUt5xPOQi6/5K70vADczFepTdVt/0s5nJUDt87
WiSlvcQSUHbP7fqLV8XSeN22UXtIZO0NpravFZKA1GQnG3BqrFbNpp5Yr9RuHSy6l1akXHeNWyro
DU5nDf8PPaPIx7VknfX+Tpdu707aJiKsEqOWHghfEbvCvLk1oz68l7+mmX8xoutQisR7KWAvab+8
IdmrsB3VbOFYDMRE3PdEEFwhLxlpWBu9br+utZLgteoFWraxhkqeU2m1/BPlyPjxuNZN8BnbgZO1
tqE/HwZcDXoqmyOgIIOqptJlZR+CF6o3khH/b9N8z4xkZgu5lY7UasZkzUq/pnhGVC87yz6/l6Ju
ETYcLeg6VTDR2+4yV+LZqYtzJw64nSifTqI2JpDAn8WpjUu45sfZR6/sk8pCOMQG0uFEnG6zANlV
B8xuPbqy80CpnT/QjIxEFW6ZzAhvH6CvCdI8KVTYoVCYxIklffqMugQXCocIssw6k/k2qojzm08K
PHE56V+wvEmU/+RXpVUPVXnxyP+S0YtEob5bo6xinMMppPm8L8K1U6dpDucq5Cq9gDAsuOnDOs8B
JcTagfVFeZpSaP5vqU+h4P2hvvAwp3yx5btHsDPa5jwbaFR208VK/a0SRZgCJL0lT6OvneOhKQ9N
BlgRdoRMiIIPBi9xHfEZMlsQBKiR4c2+OABFJzuxd34kKV8JJ/zDLlStFLQR2Ik0kcpq1FMVLYcb
ZwzXt1l+9Fioi0cehSW1DGbf15rHQbFjwW8QJ/VE/6lufVccZ9IJWyvfNASXJmyHanXYCFfHPPRz
1wdrV7WFT/GikA4HUvQ4xYxqi2TvZqgl6T1/XwWaLGEkx+a+9teQ6UEvuR4aTiBs09vKFidGS81Q
JVEeD1h8ZRTwRaPDuRX+q+uOPib1AbAzZhbSjyS4wErEOzdYLuQbJVx5O/pjfSkQslSayyRiSyLD
tkBSPqjVTfd3ZFq6S9J4vJeh3Nwu5L7f7zH4hzqQvR8GMxoGWozSQTXFB1pLANz1qp0da2rPnonV
5A0y/HChdbEaf767y3yv5Qqr1WpoJOw9ik1l1wwi+5RiyEP+Y2groi1hV/SWlQ5U4sE8nWou7yli
NdS3+6w4aZAM8+oamS7xRhu1rCj6FJr9Y/I+8ps2k1TeTkbhr/SNQ2bKdQUlGGWjhRZQ+SOdVFdV
kd527e94sl85PNWtTBrVsDBS+yTNKhSkN1UNenbmmXyI279pN5BJtRikHyWtjpllnDNsh7WZhZ8h
zuBm3CUawE1ZxC5Bly0vUWHdvjD/50L+GHbHaVPxEutokFQHOi2cRQIK9P1QKC7IdhEnzArt+XVa
j5VfTNmlZwPvm27Vsdz/bkENcOkdF2XZ+xa7CasymshUSBthXkX4K9YVBFSm6e/1l1pmib3R8t4/
+Vin2BUP16nTjG7rtrtfTv5A7yMtPPuam0ZoNRTW1ADOBaV7ApfVCOIiVtxTpb/XgK/2b0OoDhvU
JwFOKccrE4eX4s0a8VWdyNbQF2Jin+PoX21WnJuzf7GUdxiF6dXLN0+cjzgwzb2kcrElmN5e9e8m
eBn6xB5kdo7rTobaiNgDflNU3z3PQimj3GqnAeK7DqRQGTbOqIywZjMVmlR70LOdR/xN2rqU1oat
tY/7LDWIFGMFkL/HCzaFXrCytcUvOmMCYCKZNH2BEiycf2+2jYRGtJOilJ9n9m+ONN7rvtLKX79t
hua6ev+F+bvmuFU/Gp+Eb5pqO0VpuRVayX26fVvRqvwyWzB5hugHo5WdL+KXB0ow/FtXb41gEK28
F8eJ2teKzjRORtZq9QHnNXZczed8lKG83YkN67RrpzPIqi/JYS2iGo3Yygk21rA7WXvP7BNrxRhA
dTzdw1FgNJyVGeOJ4W/+7cQjGuLz6SyPmBSgjrqIgwd5jN27tJWDS7XES3RFkohD5R/B5Mm53+D5
D6s1fuA/1+wZKvl6FKQD1/8WBd6K8jmN+qv4Ko5iNhP6cGZrZJ/H+KZhKTXTkKH8aL4/kSh9VwrP
U0Us5Rp3+2UosUvywcbgpfubm12p9F56/5j9lg8E5jULjjsFqJm/3zZpq5S6GpteKQK9/CUN4orx
wVqaEgvSoKGpiijqZ77CnWTTGI5CDdN3lAgXDKHrS/Vaa2FwzJzz8Zy/4zKcJ/RoTBDKuItT+4Ql
Qi1W2o0YQY8eBCvskR8Pl9n/lieb2/jvYaFtXnJVtA1gRjfOsHmpwYsmtjO1uu4BBtSisHiyuZQQ
2h88xROgcIK/k72VGqkc9qXigKtkFDWd6hHV/UK5LyFIve+Jztkge98Nk9i5paInR0/EooaExOfH
iF9MR5zYgDewpk5U9urVPGwKfX4s30G89xfJ6gE6Nn6uB3PoOmS2wjjvvGzPAbXgqFkKNMVQnoW0
E/jwg01OA6KDqx7w2k9kDpWedVURjTJT/4e6yk/rDWU7Nx1hOILOlbU1uZ9/UOTAhl3XmTyrDRwN
VrpPLM85q5IVYaw4MA/dUOHDIVEM5kYgN2TyCRFWBD8XsOY/ggl1364V2jjFxPZMoeaBEBS62e2t
RNrzwowOoLHmzHDSzy2P4PMvpKbl4sSuHibEH6erb336uc8xqYVPXpo6B6csT9kcWAZTyzqvddXV
rnm9uS9B5F46lw3iEhmvJtziOhVKhzFe5xtp7g2I2lKeZKxNNhqF569URziKo9argNMx0JqZWDJg
txDVSjNTu330PbvLsMeGrPGSDOAUE6daJrxUxUeVVnBtDYGaS5rHfbIzxuM6a2oJaI4PqY2j8vRU
DR3T4YvGujBXqoSfWnp8+uQAFOkMn63twz33IJQfL7TjEDM+EYdgygm8D5JZU7al6oOZZh2qTGeT
YZ51R22dGpI8n14BSzRS2h5zy1PtZl2u+hBZ9Em9bihbtL36GXjfLNomuwTKpw4hRofAy244ooWk
4VzmcY0yzQ6/BhtyoK+LA4+snp+7x0xWlKFTnajWX5YDuTpQYzOgzaYdwQyqFhB/CPymRNrHLdCN
FkR2JLW9zdb1pxwiM9Pn7+W2aI8iRaWg+EBeZ7OPkCvZ1IoOkH28bYzpZ5MXjCTyGBh/xVaGsEhB
4Thnjs3epxrMjdLbrehowT5lPgSX9hnrngtdIv8UNbBhnHNsLFPtMnJmjRIqMaa1TabdXto5zG0V
YTNyVqIZsml3BrXvv24HXbQJn9EFN+VMn/ErhjKPTUHOkQ2ghbSkpT+oHj2qIfCWAtdwkPpPi7qY
LVJ0EUrDixI1MSoPcn9JHlZwihFr2FOOY2PxdvRv1CSRXNLBSc4nlDuuFgQoeGg8pjWZrI7U9361
VQ8DGK/DuGcVLTdII9RAtIgeKbTNCwR9z89MtyKU6piU8lzArOPwfCJuRGehyfooCVXyRs7xIPjH
MQSz/w2+IQSB3MrgfImis0IxJKFbBKMFyeMJJOPwVF3Lht1xdLErOiJmJ42qhN6TZkJNXGmWEt2L
gzRBGjoZ9YcSJUMvJ+LzZW9JTjBqC6KWNgzHoLbxhorvimyjPDufA+8w9T9LcGwx2Knr09m28dV1
pa+G3IuucKiE23nt9dMyDlBZYniqp6K+u+mRHC6uif9smuj90NZZZp7uj0NNXmJMrWMZVEWdjCno
dvj/jWRcviv2C9M1SFoha7JIcpi8TVOv7P2qAOM432Gsq9VnAYdbNFFDPv51d03lG96DOlZ61mfO
A7xWJ6tsUnFhrO5CiQcU04THsso7WFlOqGPtSuK8I9n6EeCD+7YYC85ENBJkv9VTcyxDiAthUxwR
QNCOKkm/349fHyZaTJBkvX0Gpia9YcZvorAEG/3fLJPgcDRNa9G2DYTouScL7aYbFje20iQw5tsg
//8Fnd3lk7jIerxKWC322ljNXb5P7YjQW/QrQLjQRZ2bp/ZhKH2P3wzeuaop4cO1lxvOAYJcKFN9
SIIMeQqbyHB/YEA4sBi0PMjWyhpmSWtEV6YIMWMzm7zER8CLX2gVo5RKChmPduM9MIvlnjA+XZ0q
LdXQIq639iYGzMM/zyH98Woy/6R7FYqv2CYhxW9mBEX5yw30ghXlxVRIKtWwjyiSwZ0TU16XOIRW
chDvg70jtw6iEFaBxpwXyyiTr5yObG1CwYwSJcu/VZ4/GHsqJr172NUE1mupWg4ACF1/sjuHFBHI
eIOy9oJaF1piCx1RSMwVRDmMRSHZGuj0pOJC4BojMDZkoa2U8U9Tzumi7St9u2Xkz/BT9ZvlUG1I
PLmP9kOgPuEAhyyPzjQzyyOMjQuOVFfFU7CC+i63H41UAgUA6mpXRg8bSWa2cY8mf8valZGvvkIG
dTSMBaSXAHZJCft1QBH1FCmIzyNwj+ZoFWw0lLQhdw/4koSiYJfAUUwUI3IxJoFrHxINV4hriMCs
hodFw4MUo+0P2IVvbgRPyqKk10o0u7WAg99VcDBbrh652JZ2IilMh3ZQg6g2t3YBWK+9D/cRycJO
pFEEs8BXVz2TIoJwHbjQC0hjdwyjymXaK6FMWmNiLbuGSKcMMArtkeIpQcSO735lXt5nd93tw4FN
/RBhZ3HuG5bgeLBBNQClOu27k6hr5zaErePvYtoQtKcDyreo44FxLVA7Ej5eNA3Q59P1RiQj/HRz
OpMR94Wv1ojM8anZM3o6jH4Yskpilze2t8CTb/q4WO82uFnpVHm3SRDOHR+xbEGrs6xWP0MHhtnG
zABHMFGX4CQfCpDWOChPgE8eI+akQBrhutqhw63ELVPn9xuDO31Ws5gw0VjZj9Bh1yVKzzYGw4VV
JSqpS/WWIj/VCqpQAAJ0J/IXR0tW/zMaDBkDkThM4KiI78wybXpW1juDPoPnfXrI+vYhDF+jhH9L
lmaq1q/AlntvMqcppkSoiCprtyuyCH/bgnm8pZlK2znj+w8NovELe/fVV5Hh8q2zSML/qos8GCfp
amujZAdqw9Mt00qkXBP/uzVKlJK+FaJrQp4tcqoqc04rNRhesfhfZV8oumgZi5NBLrdp2BTUqNhk
eDwoE+RsUUOogwSKcOnB0q1Ss2x0BWA9CB3+cTiZeFJNmQiHt2LN592zU0T2Bq1Ejvq55I16DIed
fpWVp/n0ngGWkMTCtKq0KpI+nMXKLNhGjABJreEN42rZyHL4qQv/dt3UX9BYds9XHiMJIVP1EWIj
yK/5B43vnrjGYncQsJaRF8ig8eASDp1k8w/7JxwoEnDseOsE++SLkXY3Y1GVNKbHLBM5TgCsaB4M
wpBuEa6gFuFFJE4fL9mOtyF5gbp4M2OzmVkdQGJsg1lhP82tZAaLi1Czi2v4h3wGhUqCFAcKNH8J
sPBvo4D9SpFSwdA6vLSR/9ns91V+ipqyNdaDr2tg3iInngjjzRhZvWV+EP0NzvLgEv4zLJ+sazCU
OUU3K+Agh2HMLfkgh4VNmIms0Y7F7gwUwx4vAIXA8HKmnxQ/VhzV74hbm2VQ3tWGljFO6zz2tnE6
wU4bQ8BhQzFACMvbkgF5QgH+G5q6he6hBahcjrrPfufcanyiL59wj6USET3Xqt7NWWjsNr94Rwqe
t04nToRSYHGWSqhCwF1UYX2ehsfa15dTGyvHQQkVcnFOXm1uB1/xWfhC+Hj+pOIbkzjywnao8gqy
HRmHzJu60LoOIuXm+csFT6oy1lvvIfcwMBZF5D3VXs+uu2yOEVUXsc3h4uiQf/QGgr/KTnVvqxek
ytsM33XuRlp2XBPhW0uhVRkYSWF1GkqaD8SwRqvtOqgvTb8o3WS/HhkoM+vfWzzLVg7bvxBr7do/
TPh9D/n7+2oDrGpS3draNvX1GDkAUzTGL3urAVXMHeOJlDQcD5dKOQO0QIXNvbr2CXfY4khleSp+
XPi2coe6aydD7C2fRdGhTAaFP8PMFCqjmnbaq9GhLS1jMOSCRHLSMeWPmmd3e6x5rn3gxis2VqUK
G92JLqRsco2MfOiLd5EZ1rLO5cptLpVuIID+2j01uTUnxA8dMGGqUwmzsFOXLyBhlblOpVE3Zw4b
vrKkiUFceC9Esup1DSxvPh8H2cUFp+SNO4TJ2UzxfsQ1PFMCngo2S5SjcKuYUYcc4GqqtcjZxwjP
V4wQIslGdi8HxcoN076RzezwzZ1T0xQiEz4ZsECrhH9vTsf0dcIFK5qHpJjN3+QQl1UW9/zxCE6h
hrGw2wgGNKw/bG4FisDwl5HXSfneY1MayZWfdpaRusjj9s66EWeMkm9H5MnJKaDea0p5UBQ/l11o
ILG7+i2NoDHeCCLdaUxYsoIIcSLdYU7OyzY1WRjw3IbEPmESZAhtsbX1rxtDqjH30+d+pMgXk8US
gJ0XGcYgHue6PiOocuYDBHqRg08SUvasLaZFuAqMLmSLCSM56C++cPn9Jw1rvp5ZxQNhMar5RSgA
t/HiFPbRILljj74+P88X3LVlCm4PjqbFdmXpuFnEqQco56ex6ff/kxaABaGbiETWbMdkQKGuFq7N
+mevvvO607WT2fyVSxaZ7G6mNzHs2ERANRGmGK8NI73F+IBKG6u5xI+YZvcBP19+0xdbU8KBiKcI
cNUIC7D0g6t4drRbZe9I5gkMonTgF7FgMceYYljdNQWU8N776p1cjnQL+eZ2MhcdddIasrstamrP
SDQkQRr6eZfqA10Actj6b0sLtcV9qD5TG6bNJWaVg7zZJoprBEy1zCOKPFwIQ6iTyPpqVo6pMHGv
ajXF/cZJu6qK4bhHLeAGEXUYXT8QxMkjaPa2RSyD8z4DkjO6BL+Gb5FwaGX6umuWgTqbhTlZfSZm
Xs5s6MYENVhD6xFRsAMPGkAjR+mRzfND77zSbN1OwNidm1J1da0ayOcmpHu0BRSF4W1QFH22I0iy
2nxVH7+nGvvPR/xmPXSP7eh9SIy7WCMIN+Od3QNBBH7zO+xWaZctbKH4vYaozDIET6DnxrCOtqcb
km7qcukwi7qLhw2tXKFNLahwTNWC+Rwb9STbHF01E5Mx6jNYEpAMHjpVLvncMSCt4r09FFzgeX/b
OFZKW+cQqD6z53RMM8yEdy96/BHPLIM3A3SE8JvC6GJi4JQfRpA4lfYfnC9gxtbZcFsKGi+e1GP1
b8YAONBw7uIPg1mWp1/N3sjeww2mr6D/BOSMZ7lB1Zz/KwwYu7M87K1Ub/vRMXXJzq+LF4pXhIsb
4vXtyDuLpuHBIO4cu82awqq0nILrGPjq2qXViboy/RYaVpy5in67m/fSsLgjf2/6qKc+MP0sm7xF
9UoCwcGWXcwHvb1xbU5rhMu78YgxBQx5lDyep60nUFEyiFQCwkWKYo83r9hnK2RifykH2EIGvPKg
ukzozYOu89+neubAJ2YIt5jdqw84XEfHdvCcGSHt27zbGJso0gJn4d/s9Qdn5JJH9yYYIhff3Kzb
MiAUCbZlbt7Grd7jvu9zStHFQ0hMSxqFqgKcfRvktA+OgUtcgr1GRdMeA98eSBARTVrt1SMMflXX
b0Y6VQ7qAqQaKDjLPsfCAPBbOL5YsQ8yD9R3zXlTMU1vk9vojyRwmLt9SN8YQQlA9ZtriN4MPXMb
ei8DMmrRHR9HucBbbghKWleXJTLfeeoUf/KvoqIgKXF8WHX5G/AaX1Jn8KVtUjPjRjoJ3ySXm/aH
Df7iqwaZeRjhQAvfe9O5M+9rPSyUHv2vXtNnJp4gE7eflLS9oL4ahF+H8SVKoU3G9r4tVZK8LF+L
zKdzXkcfhd+CCBwtK3hwaZQdKL91FS6R5Ovg4YefVzrEvYPLCmTYRcGifRW+bv1NDF7acQVcPKup
wGmzT4+Im5qltva5YGvlzmdUh56cQTppNpdgF+NRMuJe586t3AEtX+r+vL1NtRipdhk3tJd54z+u
ZWVFdRJJ4D2sYgRwS6Fp2i6+TaLe/Xh/etgoEQliSs5r5CcHNRIKVEBynpU4azm53a4Pvd+XZdXf
cl8tw5tqJmKQD8BRa03PzwocmJ3/5Yg8sHhHkx6MjuWzKmhBygR5uIKuwixPf9Li4fr+FvW6IT80
w55NGoA1y28oXF108K/OKxQrw5UPyZUTAMHUL0ZRy0n3nU6v/gJ+5UAlM/B0Xr4ylUhoznZySnfZ
ao5Tq+WdmdPfR7ij33rtA4c35YaJuegVOvulu2CWuQRSXtPpBCIsy2xYxHiRQuzu9gL0+L7MWlM2
peggbOvIWuKoiFlV1Tnn6W7gDEm+yQ5Ho8lzlA8EbcnUnTrWvp21f6d1rpmJzCqlqthAjaKUcCM6
WUnRptiggvQtuVollJ5uvx8qCAPj0TiawRLwPkXLiUsarxVZ1kEy632qK5eFVD5QPmtFZnEtp1qk
YntWVmrkWBEqeZ6OeBFKiRX/VmPGecmS8BLK8LZ4WJqKF1ZCdEHuJAjgJudjHuw7JBwn4T0XwujL
qN026RPYfAAULbyaO4bJ14zotPYAgEcrTE8DSQa0nFoBw6Zwyh3V/i3qsYEFK0dBVohQKN4x99Hz
goFXOdYifjsgnhRpQd/Fh5ndFGfB2eBx1uZ/rdAZcy4VmdCusesnV4OMP5QXPMD7joxQdW1GiLck
j7aSJHbM209ytcJtDw40aflpw2CZGvr6BqBqOHd95msEn8jjSBk3T/CP1RreXSgUrJevhx1rjPAc
RrEJzM5jGAYk/0GvjmBXNqWfZ8jPcloRDZqSyFdzPfpdL3o613ZM6Wtzp1eA/5K0EVk+KbT6Dhw4
ZoZynYXJZ5zKefavm48XzpLH4OPm+T+34VqFvTjMJb/w0S3ksWsRc9CiYNY9PTc0vOsktlGXIMn3
o0BTH8wAzgRZOFNwB9ns9l6CG2GsnsOYhcuBizpiIFNEWwFGJCv1n9AKCIIrgi800O/yiQnn1UXI
NSug+j0tlBcUfx8PrqF5lcCLT6Hr0o+dC8pPT+IrwbJrZNykkclIoxKnvwACIx1kVkIMQfz7unJ/
/ov7/kyCd8VJU8LLb6BaKl1JAcMf5i7Qs0vP4KqRR7NUXluASA+Cp4JL7J3Xa3YCL7HfEGDWLRyr
A+Vp/u0j6tJS1LFsht/IADxrWizR6SbdSrJbIvp/q8UP2Bgl5sIboEQIhiVEaG61JJKkR/tuFD6N
QnYlKXZLvNNdYdpT5CtyC/Jzgj4zRPkzbFF3FhD3Q1VVR9qEN6UeEHjPAW6f+Hsa5ZVKI8ph3Kn7
62Ig/eVwmkOmj7dsQ0FTQikBq5oPiamveG4ZHJtW0wsxOllpk/4SGkxG/D5CX2hYlM6TY2kf7vAG
E3191E6LCgCQ5cmeGt7zTsQoxAm+7b5z7dP+LQ7OoDxllR2LyxgfBSjVpxem8Mj8Ziu/o0FcLTOe
1bkuiBDeSHVDEyySvoqbh5ebEExI7fMZXz7xVL7lK1ea69R/amfZAMqRq1eshSqfKVaEvQfuLd85
8QcWt/+mPOGo5rdkYn6OZhuuGPshB4a8iqReLbhvs5W5WwlGZBXXmofj7iHoFAuNXpGSFDIqiRmZ
6xhUzztEUh+6za1FfUkctlIW0gKP4qSvyGJGylqcHNGX3Odp1SkUEsqy307SvWBvNGVG/ZNGVt9f
ZceOJFHEAl08NRwEYjXlohZ0D9Z2L3HWgMvV83o4/T1egSCj4ml3R76wSgJBYC2qHq1gDesg/6as
ymyweRaklLwpa3COE4RwYzi408ZGzXHwVy5LEzoT2Nic+4fv2bBZ8ph99YoQoOgB6B3C0mbEFL1m
eXw2wZdH1IX41Styr2fJOwCH3F2Fg9Hj2Qufquiygm4tQB4P5MvhC7c9tN9FWPsxDTHbFtl9wHCS
sCrNqdSyLjXQDbcOgS1mVlhTWgu3pWzTMSeL1qaHSTmpVzYJ6L8mZeO+OyhXQ3AEdxlZ8SyU1AGC
3tjxe90AivO2MghjIrj/Qx6YXXo1tbEnFpV5U6NLFizxEE9q6alugQJGTST2Z63nGZ72sgvMXUHC
D7u36mZgfIjW/LaAWuK9QoYSvXiKL/2EfEUqTUfp40MCsIZWrMcWQS4z1dtaBZrydvEQVBSp4tup
yrohICDniMGjyotFbc3rsoILZrdKRdXOf3CeT18wCCDs2Id9aslBUJ+dK9C2rxa4nCYO6Rv6PR/X
LEs2BhhNyBLNQnU+qkDkkVyuL786aaZVN/8JB81aWn4BY/ZBP22yKTAKp/8pulAdUrBM/7XmYXRa
m3cEcsHpFPsbHjnmUu4CYDYnZgRJBRXelNftLod0oUdSAGvtGXOa/vOZruLtCyD81vgiD0V0ABkg
NcGNs9ryUke4TS389p6YrK3p1ug89ZSjLwezcuiaXvsKKdeQcl2fiWf4cuszTfGRrkHrzqPXl+0i
cjFA3adfNr+NhRYTUjV/FzUv2d72jwYuD9LRiWs7C1zmMmkPFvpc+Omj594PFSPDzwdaP+JdvR4h
H+CVnzBcXdQRYaeXe7O22i30OuVRX7zlcqTE20UiR/AyDub4YjCBU1rspl381abXjDBf0SN6Qm3y
QvfxSR7A4GniyX3/45sq3p7RWSqwXQfwnrfrmAa4yP1LsELdroRTg6R3M8sGs+EFu9Etj5zYyFPz
zR3NCgqtGW98XTqpP9MVdmowF86QB3CVKfKhGyiej5n0MgJJQIFRBWkOFxaQaLiYwqBkBCmLJN9p
qTtkqvEtxsFV5myfEayHjFVlaXsQPCIR9qLATSq61OosvRnoaRvKjHYwtK5gdOTD5HOjUe3jMa6z
ePMXtuHZjhoYFF5v0lGfU8rtcIUDkXYhT2lWAV2fwl0bqlo+lzhw/oCBjtWV5uE/M2hgYamdbulR
iVCyULoYJ48sgUhRex6ljx7khy+9nZjLvbxz2Q9hzFa9gcHaB8GXtITNG4qeGSg7foQuJRSFaDid
8VyApRJf2+rj2+17oLZh5r+CzUOeFWFxn0i8MRJlCUQ/z7zCSGI+EV3B/PSXyjywBw58Cmil2JIK
F+3k/wnrsmCf3Wojt9GxbGQjZn+12YBhJO5T0I+FbgiW2g5+PD2iwAsOkJWHjsYKwPCriR0oqhw3
1AqYYAyywJ3nrpWqYVr3mOvDDV+YeM+9maaa0pakRw56byAxlAMglZjrGvlYFKz+lkANCbmSv/Le
HbCnzlYmov3nsmUKoNnEKisX01NsYPPh7vqwXjthhcSK0Do1PLMvyyCWAcvjPZaQNTgaZ+kevi6d
yXf5GF1Cq2f2E5a3sSgYAG63u5+ApXoXrY59A9phG9TfRDcuP0wvRFaWUg41YBwDthc0Syp2qg28
zfSXL9qTR5korQr5dUUURa2RkE/ibm4+oyzvpXn94uoePFsrEqID4chE77I+XfbPkcAwqMw4ief0
qhVlJEj1jWvLqv9pqnmaOg9tnau8vx/1BtHxhYefJSkKHRkfakbQOqZw4tHpaSnQol7dym/qsazv
JhvorTBp1YVSUfKZBKhrJZ3U8yRCvTmqPzQgtKYbzqqGc4cYQqq9d8XCMg7Um1mfywrtRYiRgVzK
V405pMRflxy8pcgBRCLLaM/pR10AbYhMM8BPeMT1qoR1LjjYYCkeuybddPm433rlrO6Vfew4DmDr
C0VjCbaIbI22P2DFlJm/pVC+QYQTIQ3h3MXuV5z+8w==
`protect end_protected

