

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
nFeCAmfGYh679FNL8x3jS3knawN5tfsSDW4InIdQZKBRzN4kSVkztq12/tMe1NyjxAi0cMi1p1mf
v6YsF7gSNg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nLvd2l9aDcTJcRr7PlbIbTAdTlqSll7rKgX3KRhTm6DJ6LKnYLgujWQn6ykfJMZcvIdD2hQjETEl
AVztkXcemle01ooF9vTwBqEgni3MUKzB3M3gislQcAk8dn7agiNAvn9Q2m3tmAUg8FcsXPvBO5o7
zc2EBMZovl2F7DKN8fs=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TJiYU63EGsOQzcVki8Bdr9VkW2GiYuYjy8cb5Z9/XG8LgsGJYrBmLZ2ERU0Z/ii01CLvlE1YydJn
WIDOCgh/1WFJYRL1ZWB7ohWbB1ugPLKV6HJgXOpuDQoJ0rQ304b5xBjSiLH4X+LZbHURDJ7ORm80
EFq7SNptkst73RTgLss=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fx0xQjMTeVb9mxjL6AhaMVwdj/PIeQwJN/xbL+GV7FQZ9+GRX6zMNlSaQ+s5iG23Lve6Wlz7+6jy
3JExpduc7cT4EK8HgvvuFvM9tBzkfzyXFid4kRz1yyfZ+22KyEzv5nC+jGKhBwdyJNTpZI3nBpBT
YlCbwT/wPFwnbooZqUjpksnu+YIODAUJzuu65eAi1fVwQVd7gEjv5v5TvZJi7pKcrK1ZXEadock4
fqehxkNd6+EzbUcfbXjgplHoevtQDecguFi8/Mwa08S4rFQCHEYRwF7ppgui6vwEZdLOlV0xwkTM
mTnDaR5c9k2cM6UiOolTWhwgxnMhk6bv6k1PfQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jXzUp6BpOygpeAJ8nt5CMi66bQLf3O4FAxzNCP69YWp2qZTZKkN9Js5pUdYjEyq6+T+hvf3Mcsm9
nhmM2NHgCvzt/Ua2sR3CfeS4HmlbUdnhyhBp2sta4UIVATLo0zBFA+I1GVZxCk7QB57WoTaOsVUC
PbPyAXclgp1VhJru0gjc2pDQa/fpVpchYRrm3ofLqy9j0xrV+SWGpQ58OpjhYkUlrc4CJ2UwT9eh
cr7rW4qg5+3IG/og/qjJWObQPgMuXYPtUSSA+xTtAWAvYzTRkirupyuJTtHfrZQ+vLfxPyqmXXUh
EMr2dTZM8Ufm4fJtapsCekBOiCy/LFW6zWUUaQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ir+GtoRS/s2W9kPfZ7WHJXdlfnyH2nh/Z5PLPgYkiPBMa1f/xwfEqMlF9oi3mKWj5qvsTMIuL8Fw
4jIMwjxDs0vpjprQ/Cs2x505GOF/dlCpTBARO1ObdA3UH4Pe0q2oJZLBBHdCJVxqytG08aSsgO44
9F30J+4EcZeFmiSfP3YyD72W1NtIqzXS3jeP/H8Cjr2wzBxNn7Srksj6LVHHFLlJI9kYqqU/I7e8
3Qnb91E0H13AsPi1J+d1p9CxhEzKdeCMq7m4kioswmioKsqbAao6cQdaKKbjyPutVjpZmS0Z50Go
B7ERgW2xb6/18GYTGqr5Mt+lpbXxYZT2Y9k/aw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 175296)
`protect data_block
FT+YvJt7Bjrl6FYiNGq5OmTZCocUUabwN6kKSR9CV0yAntcVVZTaZutCGEuawUpp/NfDJF8zNIHp
b5eBOC4vcUIKxjmmCH1KomWY7k4ZUf2Mj5VHTnYtlm3qFYthphZl113zxCh2e1PdjAc/FXVN2GsV
NvF2BLbXvR8J45YAXeDvXZpDWxJ+LHHUjKhbRhgaavpz7Rzo7psla4QJwEIhde1IGugtuudoavpM
9TGnFnfROhzkWy08BgI/OOQ8wvJDAkCQDELJOETLCHWDDPziMweKXxeya9ECkaesPHliVgilcl8i
csij0Th+CyCAtb9bbd0Agw4c4sQtLQJRP1+LM3Oqt+Hpf/InyU7mFH7zGWVu7ecBqplyve50rluP
bhORpThkiKcQ8QHAo3TFNLEPstfNJSNtFJI9c7sOkcnMskfp+qzzuHRZUvx+zycQJBQfwHr+S1cN
dIRO4fYrut55/LPK3BNIQ4UQ/FuVsPbeIevLmMXyrUXL2rELITGrJkd7Owu7GEnlpTcC3f6elkZF
93LOsd6/WkHCidDaJ8rbURbJjvrEysZwQ5Bo5yA2+CsgHvz99h1WX7ZHm882+ylVqU6ELD3belJb
zEMPW4JtNXIRCrSb5Gu/UzRgqdU1I660Ve0bW4bIZ2NVPk0bJx+aloAD5Q5jNqT58g7i+areVrR/
E+0XrCgmahaPYIFQ8blleO6IkiXSmKLfXdQuZQP5X09+BPKG8qJlWn1eG8pg0/TSq3IiTALoCM1l
ZvVmx5ojTvFUG9hY7Gb4Jus84WULCXiKqaLHcXIFZuUjY/Kw/B16mV5VDLGZ3qJAXIH9mwqITblh
RKF7o78U06yH1UTW+IkFUoHz85n6oIJDhVSd2lax72vdjEAZNWfoCWWu5xuGE2FWf9qBLOIr5woD
8aPOV60ZjfaYdKavGe9D2p9a4du/fMi7/tBVs920IusEaAaXu9G/w7Akr8lLwplEJpkxDlL8GhVQ
RnQxsw9MBx0zZL8AKcOG8dM5kvnKBixtBdKHtAd0ifmHQCREDWxPXxr0DezTffCX/ncaE6+Byn4F
uD9uiawAW4K5wx5R+IY+DMklbcvbUTWttl58I+dddI5L7ioA7WyufA8KSCCjen2nwr3aFi8VDbIf
V3Dv2W3mTCGrEX91syd+C+53YhVBrT24j2KYNwHQlPszs2mRlNNuqOGQlqIaFErOaAOruK5/FK4Y
30Kqo5/GlOFf9gy7n4vv6nBFyM/b+384w13YY9l3X1+QXJzwvPck/nzQoF5U9uxzeMain2UM8zkf
D4jojEz17ggCKbqbn28CNCbuxkK7+OFpaWU4YMV6T1Ud2mSEC+xXijHPf9vR/HxukEgNHjkFh0aA
uQFXBqLYwWCAnWjyQcR6iYofzSehlN0jhTobCJSQ9wjykSAxdoNFiqEOdYODyz0bZTodyoK/+iFo
5ZD8UxF8k1eYnusHTVHPJP6vXr+/ZjP+rVrjNhdi5dYANqpD/xO9pvL84oL40T0ctt3HGjAJoGO2
H+heER/Nsuhz1GxcbPUp9ITanNukJjHdphGirNGzK2IEexQbhsk3iIsokkaCWBpTpnxYqfpPLNm8
kzcpQopxhN5z+i4IEpemAScA+F2ZJoxRM4YryUvcnu3gu9Sk7De8dFa5JlzQj/FqvwLBu3KhRIyi
INRVlIOjc808WdP3576o0i+EdbAciA/iIW18AFj3FezKldrMZJdLt8tB5E9z7kQG05MovFGMshuH
+ho2LAfBTovyuJjtu3UhIUJbI8Hy3iOAlVkD8chpvdZRa+gJj7mst91ubj6ACSOQx+e8ttfV4JwZ
QHyOr7teI0hewbmqQ9qWeNI7a+gJy9MaZQQb6w2WVNkYk64AuWWZ3WNFvIoUAi7BndBkqzbgg6Rh
QIzs2+XPp9SSwpHSFIVEHYifdKzZ0bmvd1n5+KxR1XrGDIOKsPeMRfNUgcbu6W8g3N1KPLz56mDE
RIpE2OcAdioKGI3igCEds6PyYo3hdltnp1Wh0chwzpKeEXUdQmm1dPD5236yA1jGNpOwhAe9Mrjw
aPjaz6r2qjZegwfsa13LLq1FQBw/KfNWQA6ReA4+RJ5N/bGNvNAiikIMHeKfrad/YJ39TbWWZTCF
duKeHwEZD2Kji6AZF03/n1cPiTtwfPIXwPQw0CIwONkb/jvCk4LCdt9Z5j7KmYn17teZX+oG6vBC
gjkE/dolxyfC1Q05YerHjGSduiAgP9byaviA4H16ucgjFWwHZZCcAGBpesmFxC9+6SQJZtUvgH0s
XCtlUGjcyQdD/zSPXbNmY/JftY3Z9rvnlCc8it0L8hIKpLQY5wYRrbIVEMmwpKqCPR/9wMSzT3nw
vyhlI3AdagwdgrnNxEKEuz/np3VjrGoLQEBJSJZMXF4EGpSmoJWmOwwtBwSmtduMoUgbohXG9Stq
1UZrtdvZ+dnuoxQKZ2Jz774cHUC7nFGH8iQQbw41aIAD1m3MlYOwcr6j64fp8+PoV75NDZ+UlWeq
j6TZYn+xxX7IEzP1LMsU+f4vFhWmUPd5SPaRt7tab494OXt9WvNN0gEDm0X3POraEQlikxfPULhv
vM/6pjnIpFf5b36lfEP9BgShS1vaXc/kRjgy0rNyme+QJqxXObYcRs/cXlDcm4pRGoS98bA2v+IT
xOn+z+XiPYpI4ejoMpVB8zUjUphxPA4gKqpUMa4w81rZVvb9UerkRPwtVMD4KlinESxksNgGO8dA
2DGpFnAk7GGLMPunLwinHKkxJcMC+ppYQuXRdct343l6SuC6fJkUiH2ysYjw0wrcGaviONeF7WSb
tIszsPKUdTpwZd6r+o1uOaRA+gNp1loO7rOwlOS0gjpTTH9+PRlkS50FHazcxlP5HsCKOResQJ3K
96oIGeD8vE+9Jlf63CGrOWwIu+XvIGUh6BDkZJPWTioZN7IxoCOMXlE7mecoLcj6HtIO/4NC1pHN
I/LnVB00/iWd057AW6iKaivftPOrzrID0DlRHJ9+2WU23NLVlaNWT3fbdzIo3F47LxCGTA+jtMTt
3Yf2AVscMhibp2UamWQUjB+/M81KP5ffMj+ZHP0l6wcwHmONwUuvQ7jzydD224m6/7HsZwaB1JRZ
fLlfJJbLiB/ldKlDvHD+7Aqel1oupcpLGKTkcGeedD1caNj/wWAW5sSiNEQVHBm4GXMXn+2TU2WO
kod/rgoKXOMPBEQ8juqIUrTlJUPiVU9xMJjFMzUEgcFZ302nzy5heE/AeOFOVWxyhKKkz9UTxnJL
/SBo8rdMCtQb4xGSSUSNli4zweZbhskQ15JW2bIy/Rl+c0qM6MFpihis0uTPTED4RvFnef23APrD
1pbvfG+QWasbB6IOrO45UYuyR2fQ2xr3uBW8mctSfw8tr/VQU4A6dAVq2KXRGJBZhPF6b5bDxFG2
EmEUNkDZgkj0LrpbYSedFDjrKPCTdeA2dvPFIXPIg1KG0iNE6oORJIGL8s7mbIn3bqAJROSEJ8hf
TDNe5ezhmnn0ACSrEMnnKbmQ3dXg8MhvzOU/bc485KuVdWqIPyKyXxkYiIPo+BEqCkbpJqN6pqf6
XBkH2uIhMFgiecjptFwngUC629qZVOG1aDVZ4/pJHggz4XhwPDudB8ZRKtTipP0/xqOPzlLR//ti
HxWeiFnTG6NR/+d5hjTi7CFWWU1Cz+Z7vwLVRLTFQ8/fccVn04lC7wr1luYerKH8rynT1368EPXs
Lom9rrOk74eFSRjUE0PCOR9B6v5zU2X0a4aKLFbYg0Ttosya0DCSYuhCU71A2rFxnJDrqYtx4nUe
Sk66P87GFYPFZNr14RcX5DxHtl/xyvtJFEPqfC7V/PDEokqZjZ6aHP3xUp3naOb0n0cgI4LflGnQ
6PatTk9luFARTw/iTFban9ZDDbeXbkDx/aklwQP5pg2/gVqXSFz5jquNM/q689qgMSl1T54BMIms
MEIjHxW1NbEIPOJhE11S18py13ClTqdwVIfioETAY4dwytNDWEG/Fz0EyPSVYf3QW80CM0QZoAS3
rn4QuxKB2ESKNloiqhbq/ulz4Zj000QDim5/rGK4VaslsEGQru5cDKdYwKokohS8PpO3AMVZN+g/
CR3zuOWCRJ0wPyAlDb5TPxiseDfNZOK7X9zPdsq4YXOZafxE3FYjvsgIdwSn8Q+xNyXXOz72zeSM
TTxLR0kBjlyO5XhUtTzNu8jAdwdQ/7XZF/Y+iBMwrfLYGf5YZzjRzJ+WdR1Kb92VmcnVNFApENe7
Dd3SqIU0wa5pG9HCfG5f40XswmBxE1STzXASPERuKwgoZtQbvD/mZBlJ4AnhqLMptySaUJx60Vci
oH2Fik9yVV+hSG8lu5Y7ywiAnxz74/aiv0+EFghsOZT+B2SFQeKbFw5aUQBHsAwXJRiR5lbvTsy+
50EwiBspZ8QBcbEg+ad+1ingpuBX5kMztVk4EjX9RPmzIhFc6vG+aL7/VcK2xw14wSpwjBdckP8Z
fR9VQb3CsrmFj+Xwrz89bPANaF+z54WwI62FAxk1DLj7BKHVNMssfvsuqOabUipVIQJ6WM1kZmOj
JzA8EtvjZokEOb1wKf1CT9RzTOS6ZEgQZTvgceqnUifuWSBL2RFUonx7UBLHhGLnMDbvUTY4YRkv
Smo/kp7E5dABdNXwA9qWU7qL7HuYQ/A235z7JspZ1aPA788FQWZzaZpenVZ/0l653YFhBGt7CVF7
C3UohDhi1ZewkTObCWI0Yfl+QvDtiJF8j12M9GFKgoiwD6pCzBle7hTDMp4MSMbLpSfBTUNIjwQ6
beGsqrVIbSIWFnqWORMWpNmCq5qJdFwYAXDonQ4wom2bxhA9lpGTbypIKj4RIGqb+3LE7NPXmRTu
T1z2TpyqGjNO9MS0HJ+nfdniadqDFodCjnuUZdniTdwtenG0+YM9uvD/z8nUdUK8sUbCBHrvcXiE
f1j7UACodc/OKRU3TXWcIkXCRt3dN/CjUlxCZPdxl1ZN2QJU75GnIENuHARGHSAWhk4TLTm42B2M
q0TFngbiSXS14d6uL8BtsE5kXKXFXVS+1dgf6xc8u7R8b9itSgdmzCyYxY8khx7kA+JUZT47fah4
r0nli5A7QMkNosWFH3eHuUp4bDKDUJWe5h1AKPXigBvIVyOLStTO2YNc/HcmCAYN35RrhYC0JuQC
LqXilYD26A8Gg06hPqEziEyNVKY0cBL9JPYjSRrGDZ1dRQTCQzpfbYQo5XBFwIEdP54WjvsGicqs
qbX57dlsK/7ACCRdbdhNv7hIHif1v9kbhLAtDd35u+EFCdvGnhl+jyQ7vVIr/8mHb6e2NG5IA/XF
ZzT77bb9X8AdMWT9qHUJlGG3f2tjPx7c+EFLOji1fNcPE8Aevk8d6YpgUGmAI/Sk8/d4gqsElCq4
JaqcLEXb0Gc4hWICMdOKv9LklYN6noswGSOwTQ5JoIlRVm2lvw/UjI7BFm01b2wntTYsQkkOB8Sa
O82dbLJyO5D3owroVlYUo0wmwhuC2+3IOOggUGeBcBVwtz9N0G2p9A30YWCS7u0fVPK3IRDLpHfV
aaPcZ6lKdxHOqoePoDJgvmvOj0gcNrD5QiScWV4QamMllaQmxna6XMyidIctxJiMWNwd+nQDdE+a
U5eIzJgjwfunNOrM2g4ioXPoMXT4NFdSz3Xs8w+W7pEvtVR34ThgFfv0Var/1kkqzlYaaNjC9c5W
GeV5ojifOmNqO2w2x4ANAqwZ/tf1PnWXfgPcUZdl/E0SPoJuoUGcIhtqNevjroVH7zERDHyR/seV
knFhItua+fYM95CzBe6lOP3Q4VO1p/4NWAVrGGQNOQIZb2oNXksVt9hdMueCL4sc74Sr96TcMDpv
0O8BbQduYUXRsvb/Pj3Hra95O9rs5G9QHy23Aw8oXVrPvtLfN/fEwtJhNkmUuKEFOq+MPS01qBYL
uYT+BkvHrJGkEg6WADA2yzktKAJA5nEr225DiDbeJbqQ4oo2kzx8SJfOyOKPTlOkLKhuKnGxdElW
rTVkq6bixpnb2Feiqso6VZ/7IMQECY4w56MIPhk1+iFzeWW7mSN920PWuicZpPsqvM0gSlTH+7Z9
CQ/XF77s3Ajyt0LqD1ZYId8ZNEWvI6E/cqpIwkWdzd+WXLuWXqlmdrQNWr6588w2xMYaPSBxYj52
XS8AGdOQvsSMzaRLTWvKCRgRcsDhfYiO2Hai7aWfUx9gs0OgWVU5yazkLX8ZAympSCLDVw127EXD
ELvgbJ0LvE6bdbtilTzwVrM3xmBBtxJJrHtO6HMqR3UjiAdGeY7rFp5hEYiCI0SgWVbht6SOR6Rr
vPqpkN9p9Jw6SLM7vH229Qfal8dNYQbrT4tlvZTfAA+vU0aYpF4ctFynlXBfbPuWncDdkDMc0QKi
1KtXHkoxUvQQBF71vALyZ+jOQFvLdxaYaWmliGIRmZQX/Fx1tv35HsX5dDjkUncEsZ9CaMJjohCq
92F+KX7OCpq6PwlbuTGfJfBn083zbJLLL6e2R7KZy8RAVMne4NJXsn3yIkAyhSQp8pjQJAx46n2T
5g36kvb3YJC33Fa0OdN7fwBkh8Y4lzP83rbe6s00ArHRmcCQWzEKSjY80O/7pqeIZvpBZPwd1YnH
/tO2OlcGPoKmN9MOBYx6NUsi7WrVODquOjp2KyfnkAXmKYvI/EP8eMIvaQRw9327BZExo6NkTLf8
OWcF8ZvyL5pu9gvnGDtn0YhZqUhS8nMqKIK4b0pkUfpWGhKECP+jWLwBKdqx4eMC3JPtAsESoyVn
oPPGbc1w/IEO2St7/IrTJhaD6U3O90Lh9uLsY3P+Joce/8cFCyptC3+trhEffdd2GXKRk2me6Hwl
t9P1mEl4ebTdks4HJtq1oXK0kB73/hnT+i6KVptaT0XQ09xEMApkbH/dMkQb7W/2ZVGCJwq/X/CD
yvVawHussoQ0F/L9hqAX6yusRMghBH2ZVh9m4l5sKpudR+xEf+y+D33ponjO/VTi8UgV8lhzucXp
ixSchwzgQIJA4SUBjCJDaoq5w0SxDzx3+AZ9URkuQwgYr3/7hQIBPuRs4TNBseFszZOq43k4lPhc
jqXeIsv7/HdqqdEPnPUW4xRGqNdmZ3mizcFbonPh4SIby7rO/H9Lffsj7K7RDRi3h/tzF+1LW80h
59e4uHr601phnIigTutW6rgrJpSZt0zFB20Lia3QDGj/B43MIkcDFvZDfXn0WmcbzVcIavmTfEsN
Iwu6r0Pe42uClzDRRJIMWaleRPPGfDnv+twY5yci8G0coywf093XfAhPd74WuhW2JmJHFOVrjEcg
GuqBWq6Ruif2FKymjsMDACdprK2bC9MN4ggAv/rJQ8S8n9zUVetey6o3tgNUzdBegnx+g4762nT6
jt15u0Qf7384xM95GZklK0191WpfKne8snPe1u7gG/2zsUmDf9b2uH6bit7qojpNQxriMsC3Wh6k
+0XvaEwSjBlorlgcNPOolOKLqIGbNd8OIKLakSGNTRL5RFK0uh6bFsUyuplygsZWJSrfvvsqnhyv
TnvtzXf0pGaPQqlvd4UkUao7bFQzO4YQTikFK3SGk5eTX8YeUAr45MPZ/MvAABL5UkP2auUO2tnM
uAQsxYRk1yc+jR8D7aPK6q71t7H/Bcd/UsR7XBiejtPcfF+ZMKz2qffwbkkFSUvqZradt9Wk2LfG
XQ/jkOjtvS96devCD9eKQMP7lmQRs8l7+AL6Gt8XXjyPYvam8ACwkf9CVNaXkErYfau1PiQAQW16
EwCH8J8UoSDEcSzRLVI/NKMOjy4pds3sIklpEwUXgaW7bF2qaCwWqciloOp+nYS8dKe8LYfdZ72u
PoxOBRn2ims9wZuQXnV7v/smfeLWBxqlXYg+mleQ20R+q+bfspRQ3sGnCNnccGlTbFI9+NQ3fj2Z
SfPF/MpJnMt49j9kRIR0YVRVQueLflQIts6hBcC9nk2Nba2HGf92rwKoDqOrcHZW2xKxKa0CcDXz
jGs8lITKsPhA7OYrROSq2grGCsvDH9CFsXDcqY5+2LWNGyQ/o3/MfNU/zMOjUNMOE3gxaJwv4VD+
A0GQYMnLIFXCsJen/KHNFcHZnbnW6+i/fuV1lDfs4dGjD50Rq/6mqUuCFrD68z17FEqTLgEa4Xlt
8aMqnEBvV/xTKb7tjpKsgOBZahzAPUIanufWVx8keGUYTIAREabFqF3GZ+3d+bo3XlYEZHc5jVZO
185W275oGnBYhlOXWr/YbfTHKBv5X83WppX/k9Kd/XBy4/61ZMd96K5RqMSG66SEwxnwqfFFS6C8
ZIHPlTa9rr8f3aWkto1HMM94oW9pnRei14J/TM9WyTRO8fec2RUtHUBpUuzlYdq7o6Uk4KRQ45+v
fVwOxgCMnWdBFCNVWJ0zqKc5pN+uYBOw45mLVfqeMFBJ1MEmpjwo7G7RgwLys8GH31y62JR8CV7t
kPjr8CwNeejyISqXc7w0cFNZDxEH2JSVFrh9UEEid6aJ/+4YDkwFxF5fBKLavtbu8BUPQqGgDNyI
bGbU2/uqyEFL6GglXF/xnD3W9rY1B+wLYqd5HJXVOFeuo+D1S2YPDuOpCfIaf9RcAmo01w5nIJco
GCZnTvvBngSYQ5seyXMA1YoPH5W1u9EvC65peY5tvboTIMFf6kTeVQQdB5z+57whY4kiDyN9cwon
AFX/iuJV7Svr4lKzber3rPo/cQxFkwsZFjnTSc/HXMmizOgHYhCzivcKlRF0ZjqFSeRFhkuu3/qm
P/H1z3K+mrOlwJ8abp/t5kzfpnMpPtgk2pv5HSbyiaBFHzm5sSvSLXLIwoUXChHJnJqymAMwSmFy
J//4veX1v0k7b4USyaN71jX1ddhTCRDleIPbsvTf0qW5Q03EIsFIiwGPG47zKoV0rhwYxRAMqnxK
+JBYKTmkMlHKVr8gBZqzm3JRHNtz49EYXWWAH4fZiuYqTL8VHdRUE3NT1R1kON/0iuWPtLfJpwVr
6WEwE/cq3WwsPgY8pIkV3zRNhEXOF5P/+Adp38Eq8hA/CYDIBK6bOxu1H7vnkocLoJAwPYZf8ikP
XhvG6/i6vZCB4yO6Cri9Kr8OaJesQ85prcoLZQzhcm6R0GMAm2Iek6r0mwik4eT07XjuxOJGGrVq
xQoqSY+LThFleej3cVUdnCUPEXfLGcDBQ09ZRR55MkZjmTWfqwaHRXtTHwhqLxaiysHOvQ6kiEFs
Fki4yLozQgBq7fVvRLRSWd0mG7RVRhSZWE4hGNh+2Cxij5NuZ8MECvKgdvfsQgMsA07DJwPXztM8
NEVpcJfMk3IKiPhblT81YRyozyLk7TR/Z9UG4YGE7diZfMBM9pSLy6qL4Ih+45IqrGrSMIIGGtT5
bYiV6sOoKmLcAukv9s2AYByhYamqstdyOeOLpETJUixffL1pkykkHOj7RXKuE553IDk6cfCu9Nwt
A2iFfeT93m8D/axHiJTibUzJL/bwQoliM1RXjRTXa8qiC1E5oStOqZv0wKy8BAc80SlIBLOPfw9J
yJydmu+RRItwUe68yT3CCy/rL0ouUGxe6yMD/8+Q+p2kLSb3BBlsjC9zAf7JMmCOaLBxGeTudtby
mkLqb+dHnbEijgzMz4cGDQj1nAQVxId/LP5EVmnI/opOS6IP77Z6EnFHNe8v3tKccprtxO6wUIuQ
2AJQrd0YP3oIRGZPHCciY0dLa4jzKkhY4TBk/3z/EvaIUar7s6SuUl7zEYfn57/iYjXtMW2M3At9
jgkhu7ivhO+TckFM8zP0JuX96N+abgT1kkhREjYPPsqEHAHgqoXNAx4Nd3MQx6K+CPgVHAOdNj8w
nplskRIFr02zvWPqM35AkrFdIB+U2qvx/c4vT/ZxVuoi8OKeL4rCt7R/pfGnT3EkPj0mGpqh8MuS
YQcB9ti3EWqntrX8qkO5L5pRV5v4Y57qHSC9JIPHOquikz9IKj7JMDNw53gd67YaJNnViyfGgbQR
44lXnnBDuMw3BqVUiDC2n9z6cXS6QrFWlnIGxBUI/L0ZT+UmlwntmRremBoCDVfNi2B/gb6k++8g
7AvSPZG0SqWKFfgxiVs1ml8CvvDT6UVldV8Hd2JY62sonB8hvnFvciivAN0UmvGRj4fR6nam0YC9
5kCWe7bG0td4J+N8e5dEl8PDfL1vJFLvOkYmaHd8yCxbZP0jh3oi/0SxWUiG4o66GJwmH1CPGsX8
X8CGh483z5/JpLH0p4cWS9R9uiaXfd2bZib5W5ZzDPOAwo/BECdUZxaQCgJMq0M+89xCsDD0avnp
XcKYYU0L85hgKrBHuS3nywqwY2X56CJ7K55Eg0Fzd/hpG82qgTSBnFGt9rKdsWjWylF/Z6Rw9K/S
vke8KliUZLEu4w7N8r5N4af7OtM3Yq9KpYXSyP6EvpGgZkDoocSthCSDG2dJ/03YxXoOY8kyTmAy
ZX6JzBdmRepfz31MVYRxsIcMFjjEZssUYlVM8mOqxAVKfnT8kWBYwwSbFXLuu+UExjWk6frJGfMV
ZClYC9IKUdTyv831zG9ngs5hdcdOn5tQk+y5j9iWbO6Uc0ABm1d9HJVsNlkfzxtI0LVH3UA6gehF
fLHHzBIdSi01gfOIArPQs6dXRrhITFFkSt6NU/ti1Ay6z/2pzmGXXXIfRvMGbEXfVui0xpkMWCIa
5KZ8OR5VfdNerfStH+R1XRP6SyH5S62X3qqx4jmUhWqr6jOHouuLlOo/Srpr+ollLYMMwbVBvggy
2s3fY0Tre3TrExDRHeMjC7lR+Grwv9BTJE+01OWt8ijxwkT+ravFgUIWZ7tgKY7tP2DISlgW5UYQ
asmlygGyoVt7O6BNWGp4Y2A4pWtnYQ23Xs4oUNBpNM3d4K+BBlaZULyhKj5sfTsl7fONOl6ea/67
s4jwk7WahQeJwGR4Td8VV80FY04dJBEl8rOpqtlDAr3jDTZSKidxarJgE6nXSVcvlUGofYOyo1eK
A085o4TAYEiPXCe6Zl5k/M3l1e+2Kbzu75mAy3PknOVoLeKDmVen+uZKt2USXKw+DMFmzbUqainz
Me9setxlpAyBKqCBwMAq7ej2osvyxmwiYhaj40VwpJ27e+vBleJNhdgIi0ezAFfDiaxsv5pSBesr
mz8M0msQZUDFZM4Ye9PSeTilsoghQRbDY8McMhjGW6yarSfDbRshkC8TwnvZwpNDox2Ci68ghG1P
+lA/e3s9TUYZIGb1oAzH0UAT+IVy2CDYdfONk4idKCh6UTf100fMRSo1EAQs+bOcMK4gBaUxR5oj
rz0nLZ6XAzV/4XH+Oimg4oDj8FKs9FQRAN4YvjiliRL310xz0Tu2ZgeaqfYTpJiDoo4cg5cfoMoH
A/hyAavTQ4/uXqw9512nCnFppOB1NTOyErgyJwyYenB7+IqmgrvfZEzmEgKcTyBFTcsAfbhqMyfS
FHK9lr3DvZUfyQinCB2Kf4SJq4zdlKKap6T+mGU7B8ROD/1clmNW/DTAN8RWRJEf/06S4FHrI4W7
qhrg5cgEMojcE3owj7zbpyEmPlm56IElCP3ZlJhrecKWWHlMTn6YWlPacrkq0QaxnueenSqS27OG
/Oq+VAsLfWVMX4/uvNiAPx7fvq4zulTPWFGapv4tRyFyE47M4PqoFNRkfR4zF4ejqVplN88L0tvw
5cZ5XWYjpADudFf82bk8sXdnNaCGi77T/ucSmViBueqEI5XEbj7eJLVB6tytXuxvfEV4tK4aXJ1g
n6IRxDC5pfvqAcnziyWqI61Jq37GPKQDUsdGbLaFoLc9USKI9HRC+ZNZDhMdATvo/gTPBt/gdzwZ
EW0QQeWC35gpBqsaFVD83WQynOQT62MJ6c8xm0XLGvgc+1c1/zefzcU/0loIygE8BgMmTPv6Azi+
8B6dL6ncEnCx2CHvsZ9DFAj8a1Nef9GIjkhw0KjKWIVISbAgYu+uyN9MufOum8VeeyrYOVA002Z6
bjb23Yj3KV/rAZSeeM6ZJGeRmoeoJrk6bttXI9m2m5vvlycNMc4CjK6LENEG8epHsqFPS2xYasOm
ztcxSyPUuxVTHLKVw49Ea4bGvgLwrVbnoZA0C81B8OMKzqw7CrWMLTUV6Wftmvk7jfZMNcTn2/uX
RES9Enuc/8fFOGM1NjWSKClLCY+coM7o5GVcgzxjH40VbqnKW+3C3eolYKnZ43C+3/sz1vZYW8Ka
flHaXEGf/B3yiM1DxfvVnqfpc8nVHJklojHzwRtna/0rIjsV6VyoOgja+9LKfExyixW7zcDaQnFb
RVSTsFjiV2nx7o4UR+I69QZ5XU6gMpFWqMLJpBMgKdIaquUTm1twdkuyD5YiuGSeK3pO18ow5/0R
q8jchbsZ+CNmtLhK8etnPGZyjaDCOL3HA1GakWfAvBsJLnO+lbUHGcoLY6GfkZmQ5CYkNKrqCOh6
hVD0UQJCGyxsgYJJjQBMRhl1gIf/cKBj1B90QbyviQjCgTpLR4yO1z8UruPLUBvwyoGhg1oPj0Dm
P2JqcqhvwK7mlH2tEW6jgoH/URG18YxftpPMxK9tVP4W+9g4cMRrD9WR3Rgz0tLIbOkWhLAs418l
iv4XCSWrcFevlphKRXn0P8r2d+LkcsJRlrHZSZ7796k6C/l85SfZ9W2fryGz5YolWJQfPz/Rw9El
INBSq3vjMuPNgD/+WElbn4mgsY6BqhRHM/jdwwnZAfCuVtspqVFHImOhkd0lrHB0GIFCD7gx+Bjj
+8vZNs6ZWZK99hp/MrbR22w2S3URbpYeG+5Yh9BFA7Xc1PmqBsY+bUBtAndm48vOkaPAvJSZ8Lr2
NRpRziDLXiLdMezilO4Oth2hCEfN39f874rViWLeUBgKzjt+cobQ3mSDftkbEznZcY5zrU32DaxJ
MXbr52N0zsbNc6zDY811V3scz2CrIQoLkaXDkGMSDnEGTmLby7mQNm9uNyLFV9gKZnf7qep6LV0o
t0+6T67FMbCLmPYHC/Lu0J8T+XxtGF5FKY2YjEzVCEbZdl5NfN8tITW+6O27n9Jp8kBgmVXBmeCB
iUAXORGqTYrhAqLytYnm7ek+cAhF9wVNfZNp6C6OsBEIkRR/oGnTE8k8sJtvrdvQjXyOMS1nA9bI
kVPDNOoGwkVijqn8+Ivs936L/mnqyZkdchUWSO5Mk4LvswXfQiIWecB3ESb0c7werg3VxOR6vvRq
EZpfHaiIKfpCFZSi44jABbH9Y258MO0vcXT0dpBmu7gaKR3HePrYfFrsijg7/1AcGJoUqT08AI4b
59IuH3hKnX2eKHuNqZ+CVWbTx0BhFx5opCAuL+aHoabF1QI4XcyxyeFaNti53peP8ghw79Kbhl+w
ecftMpSta2nJ2N8MgktdrLAkdC+GdCZOq6YeJSf+T4G+ei6v+mmBGhm0Jssp5QqS8vYLf3VO2/Jq
/qetc9PcMgatYWbDl5OJiNMTxjY+N8EHXy+ttvLugYZXAaaG8TIaruluvjOaV/TBRLyFEI/BgAOQ
wjVzsO1VIVNiopB0ZachAzFI4eIloBRWP2uDbuqJUYyfOUCwKAzx1X8cgDysPU3upvUp9KknN2nG
OLw7R+vM5lp7AfTstPEG5kU5JXJx6XGvaOSQfM2ZknaSpyl5gdJKaqc/J3IO4q2pYH6de5G7y0U5
MQ3x6J9piob22idK9yoAoh6PGt1SAWhy3/1MHVkhZJI64CxCtkggap5VqukZc1CpDDa2BIssd/S3
3GKkz/28iP8XjIXHce1goVmvYuJsenQ3pEwED6eUSvPj37gi8hsIhM03qLo7uAM84LWYyM5RZ0gM
ntP2eKNhXy6eoBpvgXlgYQvXDXFRS6vEhCqJGn+3pdyles2mveAbhwH05hAMQEz6foXHJkvZbEYs
IAhVeOfXRMpqe3WRUMo3qSVPPMd+QwFKT6P3Z+c5TYHSrAKfW68/RvASJ0VYG0D8HY3p4xKjxQ62
GH466aTr+e79aQAy1NL5XaSbGWK/Nf8aKcI2H8KfTndyA47AFnrHIOPDN64AZ88ahveFr4GjLKzi
8+PygDuRyQnhw0T3WkrwOcrMuMGmm7jSHuvC2JiAeWOpVtC03lEQC/Xsl5cjndK4xPmTyuD47Hok
4/rVyV+XMtAnc+RMfspmCrXQwbuHCZKfgTpUw3kx5NOVxT1F2DEhI9yzewyhhyS/Te6cvp7pehYL
2eSgo87wDdOerTyX/TyVsZQnMGH5ppkhix1n8SpedKtoZCFa9hAKH1eKoG1zZE7NH9NkZsUxd776
GzHKZymOr4SusJCdMrz1e6Ol4vSUpfjAomVrmEco2ht0PafUfwAS15gHgdMoOArO45i0KDRpMuFr
mJp9GlVuzug45WXmbfxkORiWI20fxEvyqRINrOwpVhoNhYnyItBhqo5ujoFzxTWhEAL+LEFkVony
taOfmj4f6Uape4miNsHWGUvsC3eHKHF72WIKH8Ch8mW9p3luqPjWdgG1gtuKhaFMy4/UJpj5JGQd
hkkN95paDYfWtt7YBPUI5yT9dX1QdWU292sK0iZdX50Cnn5jqQVy6Izk3yUOm8ichOnHTYN/yzcq
5rI6+9U1kGtYkEFkMnzG98hceEPTsToqH5VK+U0MDAOBfj014nfvXfSpvk86mQUfrrkDNQvNSdC3
fBdtv8HcD56Q10YYjrDB6sJ66JQrgHCULwL0aLeDCjt0h/o1fsSPemgynI4nZfxTyLyDvTRLpp1l
0VXBvmXRJmHVIk7K0VKIFii0wmIHmEAaxY8HecmCuNzboVZnEaLrOH1N+g4ZT170n8MJfzFSdz2o
tVEUXFupmO3wCAJceiTMqT8mMmMQfsMQIY4zx7lXzB/JTvGYFBqjxtEv1fSB/I6EISCM3QIoZBwW
BVXuBpYjYrKk+qvtK9UMtCUQSjUE0Lf2AXtDVbLe185MjIqzfkt+yrK3Sxe9GsdgyrnlaC4BrUcF
lZwqXRnIgXX2vULGcIVeRxdiwwyTkF2wqx5U8jw5nKncIFsiZJTnn8G2Fx5yKDrfdSp0I2nODwzr
Lfv+F/wpCBYH6IX6BUuPI4/gt0wEiKFszWH+Q66yffGnaZIDJk793TIU1z7YWY6qpREGQeSW8oQq
zvwJcMD5o3ShCf90lJbdyLID5JWQyeY0wOmfHUVdlcUk7+H1n5nWNrntBWuBlVtL9Oh3Xr50y67P
Z+tAf21ydJtjvDbX2GbAXQ4jil1079YVh4P4ql5EB7oYdMhtG9luuEhVfhHALLKVH409HjYlKvJJ
T6f5HscN747PbSsfWWf5BNx6h7wTcs2qs/0gvweGI4u0/V3FRZU/ue3vkTtrmPiE14JhlW7VLRxg
/cUwyjYToot64Vp+nIKCWeA8nNq4N4fhDa0Tcy5jPXzmnIPI4h+JcRWf42mEmfgUS5u9iNddQoBg
Ru7FUgJVouSiMDhP1rXgvaXE9/ota5pyB0MfxTgi1GMbbBvwO4zX7wgIZZIFfZgJ1AOGydtduy9x
iuoWMY6giDRi8ZqYvQ3poe+NabNF4I3d6eM5oCNh01pMzLuuevGa1wvQXaR9aomBY3VmWkYJea+T
BiHJYRZOqSO36UIvhc1rMDy9X8aTLNnWhjvTn2BOryb1o1CoTRq3NV4ZHWcmABEMvX1zZg4FYjfs
zCBkMpUN1efFrHtmZSr+DxryQyohpJ+8YHt8QHXSj4DHwQHrEqEVL6Gd+9WZyUWKlGoeURoiF3WQ
P2yVLa+lLvNvuBPBh598neoVd4GdOWGVvBpoGIw36KRbUOqaYBCR+eCYHmabNo9ZajUDTlxIVMoW
I3ecXwO3TcL7nOMFpH/C/afJ+S6KCCTqfh+B0kf45nQKdQjdKNb9Ngyc5Rn/quQdIW3c3f0RgW8I
ct/XY3sdFOT179Ux4Bs+G2g8WhsP2DI1liFws729mfJS3MLclDgk9PjbVZg9hRQSrWW7t287MVAC
c0UcFwC//HnrYkA6XxdBOOlCHKZTxdiYCBSXAGXN9TlPSaErtoRQvHZQ/mxfo+lVMhU2jqZTYo21
LAgCjzEnoKNaUJMnCNE/x087CpQuP4A+uKq5pETMWDQWKtyx4Cln4ySkc9R00vQagEgQWdb/Y14t
et30nX4rCVPHxWv97ylmO5div438pzSRHkfdIQ/3WoKqQ7DcJ9D83QeKSQXzrQQ/cWvApmKZvXBX
1mfhmrv5hk8RjGv0rdgfwKtzSorVY8DccQDg3ESPtNnJxhbBiKc680+Yh8Sv5WymdD5zWpVRfVjq
4yaCAj15MMnqfw6pabHp7b6LBaj5tUg/64UM90XISqfEWo4T3WttSKhFg4s9eeS5fcq0kMGZm/nG
NgBeWxHI0lBsiLR/ZiWZNSmklh4l1n3rGs6OAryEYVib19zhWr9BtYZLQebdowPW45V4pH9fR7LK
q86oe3xVJ9Pl8svz5g+qHnKwxRHQWyziX3zmoXIMD5oR5aR91xXFGVACqZMPvcONhMIjtkBUUcY9
cl4VyQnK6FKL+68btyKGwV9GYibQxoftdI3LZqVBsDKpZz8iPmdSJrNC/dgJ314gX70eB8JvNzBE
h8+IxdpX9BnaI6zSoPQi8HrYLS1bVRjJ9YhuqtzR6I5rUeGmaBacip0KtDh/pzkLauwtpacecP2h
YF1TKzqogmyxslD7eOA+Hx87I5e8AmQv32YtC9bRS3C96nR/ACeQKQUqBtcUE9OcQKDvCYIvGbe3
/DlZ648228S1zhqPOQLIOjg7ilVUoTgs1EjPDeMPfD2NEtntnYP4nB+HGImDYtNSV82vA7tJZxIf
nkz3I0rb8JjRGuRcR0XKmKDBVV34w+Pg/2uF9P0y0emYxLakUjhS+oP+28VCqrvB37NSYwvHgukQ
9AeROP31SWrothaA/puFWnRZhU1B236avxbr0ip5N1qBc4YvHhRI2pOkl57v1XyMWeNUgKVFqxOK
86ladz3c0tzPoywfwMqdXo0Q6Qvx4WsLksOMWocZxPGNQzWzqLa5wthaxsf4padpi43R7inSzS3J
KYSdWcCi9AT+ap5Okg2ADcJqcTTBqXWwvbxmToADO8Cd6oX4OPEURTcOzjjGfFziqKUeasf7qUBn
331dWr/sAwLURHjJr1GpI8tT7blBnQjDep1FeQUJE6n4nzHVx5TARgoUWw/3IRgItOhS/TnYJyF0
Xg9tGaxXQo3e2LnL4ue55doLM1SHGTHUd2TaDUOweDz6cJswn/EShNbpNjgrAwXa8X3zdIeOExEN
EplJI5Hbt6qfcszP9rvwt5RtVSbh5ShrYjQbo5X7WmZxQmDZHSZoXGapOl9OkL/Y7vlzggN9OpgL
TVvPiHOBq3C0YYfTmqHxooCJGgDF9oTe9vJTqqxFsd6HsttbtrGXTvjDkrA3LqWt1ZY0ZVSOjoTs
wzfcg7p4joCS+Pslk9sh2q/shDuluXbDWNw4aXPGc/cBj/lPcjMTuNyOUwuIWira9mKytTn2efJ9
Nk4RkLLHhAcyFakkillRACHexXTasuY8PdYOHNigMRKsw3F/o/e+TfalKgIAUb/Kn9Q+YIFSMUc7
V9xIwWWtEsGLY2jwtqI0927/bfY6tzausPsJn23ZARAoeI/RJz3e/ohgDCxVyH6i64g+g8goGRp5
TELFiWvwOK8gQEJ+tVGZAvtYK9x78P1PYeMREz6+vWGBZrvcdJ/odKkb3qyAzSM/M/SG6y6Awbot
LZ8vkGvvIt2Wp5vHEaXZxVfX7BwgANpdIhDl6BOHm36IKP9yYLFyMrWqHKJZxQvHzexHYbQbylif
eUicPRMIvdqNstBYMIRSsGdPvPdQxUbVnBZWYKMCEXhc21I4aCSXsUCQ7E8HhwSI21XKhlTqSkSd
mdmgFnjUs7ksRF8pSoxMKuUvnuL+r0rrbyzAu9DvyqiBRU9Ds25mJyjUzj7dTNeWT6n5vjOahDrQ
cfk7DusjlELhHZI7DqdGdV7/Xdsv+RyQv3J2cjETVmmJgIer0CgynnTqghOrGnkiGvpE9foxJ72V
HpQTH+2lUUELmhXeJmUXS9SRyMJgDGRh/gfPKtgr4GAKNeTFpu/MsRuvu9kYchl7WPW0VFtru77i
Gg6kVU5UvwDuTWWX0QN1+Z89CgepwsIvwDSOrj7s7AcsMLQB4itmEdfCWEyHmv5KC4ryd7vqo8MZ
WSr1laqu6mR2THbLWGxOap2Fm1rH0MjRHQz83SxwEY6LC5fTax/ideNMZ8okM+VhTrCD25sVadzI
DgukoqOFmWxkaMHBZ9IMlkIISwiPIt068Cau4wY/rAYvdzVgMrWxz8FFwbfmRvUDxk4b4Hn5nMw+
6yzqvoFq8PSuDDjl/b6izR/TiDfK16JmAbl3ubwY8KGWiVcKEBsK8KSpYK4jYA2UuR328rz/QSCV
HCyCs6K1KWgzfRSPaR6OSL5hpjIw3HUHdwj1zEgRRLvh1hTgPEcXJGFGcqvLSmEanK3fj8Ke2IUW
BSohPLwt34C77cNz1jJUVMRQNKD3HjlysbkvpnMLzUtXmEGzgt6gkHbur1CreMVq5I9/Yp1/1MCi
gvAilOsF9lr5fA8Eh5L0caKimWolUzunN9L8mdnQ8WVdqYIp3ZvyzAAEIw8RittV3UhYlDxTV2i1
ywdBUFGTxjPZun4f5rWWIuklODWp7SqabqJISf6K6x51W+CSpu0rb1SyJYz1m3Qc44192D9DuLn+
6PvzhfV3N2Q1KkfqtdaQ1PAIKyNRnlGr2ErzpUNlyWhnolLl3D4gbgZg4KxHqvqK4BGXldZab1tH
9umcgf+5jt1CcUSLbEataplGzWuvH+IRoKOWUZOOspq9YNlxW1TFkYM7tqRyQdYclRkiEYIzKzaA
9sT/ebe4fJUxtsB9mceL+TlM0T9HQ0v3GeTzNDayQ1gnnKCoDzaqvFIgJleryVX50Nbz+E2E/eRw
5RXSivdZJZF0xfICLziHl+tZrQe0PDB3DsjTwkjyf4P60HsRXxF1kKUQ2AlCXYY3VSUdwAwwUOXu
nJ24n5N9MIxyV10er/TYEOaggij6Tr9CsVrCiFnv5XhxVQe1G/yMVxTtV4ig//sCzJOzjGHOzSJ1
Ps122APJoveZSv0R6n774bTn1TK4ZJNz4U1+UZBJk3FtlqGgVjjahaL8IMXjgz0RelthjI4Rsdzs
ZJLWvCAoirXmgbePye1AkT36wrHPI3xZz3DspmtFF8VhIVT+O4xaPNbtdOc8iqc3bDqTpAZF8grb
nNlnFZkAoqyYy3JUmdXoeGCpmMaEscbHGMzKrAEcgMoo+MSmAU1gMA5WrqqUUtqdMy3S9hGCsN1H
IBn4Dkndp1KIvj0Mh8j0+W/4I/3Lqa1/9pEoossZbDpcRTUsv/P0+7FyjqZKnVq2Jk8p2eUXHVKf
pZvMGzG053k6RIHlHXj84dFWjtQV/27MXBDTCClJqDP46iDWDs4ATmR8KrX2eO1zAbtn4gcYX0wx
h2mtQtcidoEiUkJgyltBAfHozK5Tb03+ouIxZqwGSGBP0UDDgywuBKhm4cPpAAISzMFP/Qbmf1r5
Lca/azzfjKCp9fDo1ZzT/HMBV6K1ml2eo/GCiftYYKSeQAaMxQdOnSek9mriOD8svvNbBJW79vXA
BGpYkT7sl34A/lJAJ/Bf+9OugiuyRfwD0/Rxcw16BwC10ma2hILRm7i4qaU9qVF2sK8utiAIPDou
vwMfSFY0LrgEf8Hc3nnS2FezrMxQYnA7RugW/vApzgeQVoMarLELVJ/vBNuoJRBHz8chG3FvIMaG
DXFRx6Z3TAwVprS/CodZxtQ1Q56KV+cMDc4wgcaW/Kjrbk/WGYPggJzKmZBZx3dDy69gKCbbQZHm
FJAh8/j2fzbpOCLhZXvkUmB3IqaugF5F0eKjo7Ei0jSCF5Z+qMDgj+q4wKbAh87H7rBg1rxFTG+t
0tIvKWgz2F/0n4APz/TMdc42rsjQvsJCGkSNEV9FtVNc4j98gJxgM66Bpwrp4/3b4yftjMUHm6em
14OBMGin9TNtnRCBBxCtSqlWdmUM6XQl575P4j+Dj7if2VR1HRqgKmwH6Exu3dOU4/V++tjqchBo
iRL6Ro2sIzKvtPPmh6d3NQij7rniSOUHD5pGR6al8NWUKKQTulcZrI3+0ek4EQ1DGNLfaxrz3way
l6KOC4s/i8maGLXp/HR6Gukw9NrySuGv+B42qoJZL5HV82njhJzUISXGp0A3/Zu6LNRNf7+Uqrl3
jO9Huovw1VPKuWgJ5Ky6daVf1WDVJm4vQDD+wzwJ8xVArEu55Pc0XaCoaSE0BvvegeSzB0st+7U+
+hvRtJemJHMP1Xk8uHZvBlNhkMLc+4Qv+x59Qn1vkdqk8w3rmGNsesKm/kr2EtX4LelAhGID9Ryq
bzczuSLmZaVR8NTbxO27yCfdI0KsaeU1Gf2/7WuzJFRiSN/l/TC4j+MPXH3hfcyZ3NmfQ72/2ZMI
Jd6xiPxbL7FpF2SAxtpYItwLjQc3CXgRwn80R2vbl0cqYYd9+Kz6fGfxKFeczLlENVyAoE9kTj2W
T1SoMaMxysx+s/DaDdD7vogeVf5GwkDsY72eLlEcH0dMrMk//ud5T4HbT9quIta1YgAWLHocZpET
c2arfWLkjSRlmVbtHyO5hc6Iey6ngNioStP0KvOQkiUeulbVYLoBaFFk6RCi/tR9/A4Vhs3vPf9H
rPew3833cUatBgV1MKa90o8Xuyct1IwXxCz+cnkqTFjfHZRjY9XllNK2TYMlMse3ht6G51doZWBk
Ny+vs2vsw4Bkr5dqWTyUzIMCMnLfWp/ybOQMVWteDMEwS1cix6GgRhbfO4JkJFOayBpz0gQFAyZm
cUIue6MaoTRwnjEj/Wo/UPWW2jHpigXjg61/E3INxx3NbGW4Sy2ViSudJZ+eeYur6M+avjniH8sM
GebU7xGl54DxuwQODICibzTN7PotvzUYq2k4hPxQjk6OPXVbqpxGOWVyljstMcal2IS1/eR+vXz7
GT/xR+/vLsq1YIQ4qE5sVCYNrPWT5mDMUXpMvjspxLJI7ljBQaqzrBajLRijIWyjzUYBomLQU+cl
g9bB9Mmv/mLynn1lhrTHOVLpGCRCZRT+L2U0bMavn/r6gVyDZSZ7F9wCWFkI9lheJ4tMj4h6Y8df
/e4GNBhIXvzKdofVRGviyXArgLY8iSg/+bFObk8+OEW3NXO8c84W9nG2Q6nAaboCHhI9GZ2rv5mA
R9JJagwE7k+5nwSUtI17SEbzcp5ITRC+QUEQl3ZroIf3oxAuqP+ZlRpcPnAj9s3vsLqIfGYZEomU
MYvrhotTmjcJ6hH80SAGTP3LvTeh5+HF9fvyybg6/tTKYr4a1KLaegrVcgN3KzUMV6ESj6SF08Cx
dQ/mY4wIHFX+fRp8bf9bjKZ6nnIHNbTQLmje8pbsISB49X16bh9xaeI/L9PpvFhG7sDOV5oIsi+8
SojC90YDj6F38W+jO7dk6FGMDJ9Q0I/j5vJ2LlRDAhcP4Lz+qWgiL2+D4Pxr08GrbDgm4Iuao4Rj
/fZGV0kcvKS2gzrOIzvomEvsCOfLo7BSDkXt4Gg++PceeDHNhvz59EA4yR/2xAvYqSBb8jH8udvY
nHxM9uIVZvq8xHvRAYR/z3sXf5wfZyNJer9j6XQQLbdM4TgKP2jl730utzRnsWoQA+wf7Qxush64
vacKyCNv7G7fiT5HKRCoJqygRjIZgPIu9JLhEnhcXCeHk1xTQif0N3JnT5DTMtudb7KC0Hi4GPUZ
CYhoydbQuHNwGHXXS2nvo+Gu0mtdbxzZzYu/HsHeezdcARfZQrfepSGD8Mez7uhscKI8jO63LeAW
1mHJXWTTUanG7AguO4KHHZs2jUGc20HyW1+JZXeMAtHrGKrKe8lNozPjRNsgxD1C2wkjAu9KbIdB
0sJbRH4NbBdrgHGqyvSNwxTnyo+Pmlx83tpzPwX/rh+OxOGSWarUZ6OwHfHfcc9SBwD15Q14lpEl
wH3pNdFX7F8DvFfRB7L5Nd0Pv3cyAwj5c1XIYVrm4nAASDGzom+6ayZ+2Rc708qB3eIEzn+VSv1r
Dpr80Dw4C8gfmt7VbaFIgRQROOYMDTNLwYT1Sd9lr68IByOlGvfYiOG4Wsw73y//t8DahQyUPDs+
B9LDY/01XI3icZ0wzDFfvUnYV43o+cTqqYAPvYtttRzxG8Q/Xnl4++QOihXu8bHeFejto+U2qJ2/
z5tPjKs7SssgWF6wfw0TCHyawf2CU8ixcF8MYJkA8/9x7ByGGZ241tOH9xGpSYaCe6+3jkq3MosR
om28WqyiLwoM+MP1yleoNHbeCn+CxUrj/elmxkf4mAY6ite85e5bqu8Sy+QjRJRlmGdeDMgBLthq
dR0KujaaPp6VQdRXsgSDZ3zAsp50IxsKK8eJAdM9KXzDn5AK24XYSoFv/b/9d26e4aTxFT+/dwDw
SvZsfQguoQGIx6nQhxkBLIus1JJqXPKOPmUcWeEmtG7wgovnfSF3rH5Fmcm01VupNYU7TQZNyrBv
pa8lXO3cHkeOBCCAt2dIHYIW9DdZS5iNjgwbqL00NyEPb8lrP7RkGPp/IJWucX4zbmQBswzr+Ns3
HQNtg+mzf2QlJYEhgxKZv5gUn2j9q/qMIyjCnXk6HeCxUbHk2Nnegzh691QLrW9wC9XD+kdI9T4F
whdVSnyjYSKYVY32vYDw3jeEXD/buT5BlSGFpBl7s9K+yjYoo6aIQSNXBwW04pZT2fSe3QAnubpo
fagiQh5cWduLQnCowueQSLbL7NIREcn3NTUDO3gGB9IKeWPHLuDcmWtBZjymiXmFHMSjezbCjMY3
cICwdCzENk+fXiqmWo5rG/h4NlJxQx3kNmINneTcEabBrz35Bb6jtrDvIwgsimEJ4ymCSeeGMmJ6
aQtFK1hs2frywdbuD1wYcSUMGRc+RuEYTCf7LhB0QPxUy/tAspNxFqbR7eCaA0bTMwCjh5L6g4/Z
ASq2BJTplRfEOlwiTbgwow2yukO0NsSyEEiRRdVt1LSgpU+yBxsl9dyCXRH9Mlz50G5jU5R30Lpl
phvgF3J7TyL4hD0XIlPHz2uIMJ9SKZOIomP5r7F6p2u47xz/BzYFavilmkXehBkfNzK/LefyElhY
QdDBw5T6bHK6wGeNqL4WirNX7uCrpW96VnxMJUFfM484i2DxGzz+EqsY7sXrUQ+UrVrqAwqIsbX3
FOJBw0eJ77swQebl2HFQzOOl7HMHVXQVniyK4l1pPZYmshGKnDQuYdLmVk4MXLYxhtdvLcQi0kqZ
Cn0dnGrf9ETo2hGEJAu1xqIS5PaFO2XJ/z5dx0goGmifA3F9x14TOiiLOZ09zIts4qMgsWXk1/Tf
3du6PaakcboW+czVJSBBlG3m8Nd+EEXw293yVAywzwBFbdkmGF1r1P62QP2M29i/6iUhkMcnxxsL
zXKWQrraRFMlRasg2wnWFGO13H2tQ5Hgloj23sbooTmfbuG5KDe1LRwvHm+Kp1y0VZnIojP5lBbG
wi/LA0nGc9sSyjbEUgbvOhZKR9lwfD2B+Y+BT+44lljHcjEHYQ3vMNCzrYU4JJRHyaxTCIdVlgd9
hndV1clvOeeLkgfnFG94x16bJK0nh37KwIosjOI4ieVprpEKERp53qRrmCJpEqfzkFOp1i+7Ph+M
Qx5pfPiEb9pEqq7ox2Pi+PhnXusQ/G3koWG5aOd1H3M4a4RcwRXgaRWVWT1rI+XF97GzGqAkWIP8
OUWbPAE6ZcgrIFjuObwVswQRxvzJH0LM1f5jqFfWEPmxoSMPUwqUCcNocC3uPRpcjrFIeDvoGS+L
ymN0ELXBWbKu4IqBgmHIZgqPtMBWDWHGgxGsn99M3hhEl/VILW+9j/283b7n1No9ARguFab+/cgC
tLoBsGjelx8yLy3TO9mRBkSEK2FPHRUflxqtbuiv/0ggDPpDc9DWKa4BGhc0u04WkTgnRYJSqqP5
51Y3KI0HVISkm+Lro9wI9o07YbnjIN6sLQU1pEGyvqLye+SVXWhwg5o++vm9EUlKhFbJTzK2+OJa
k3J18Z3kzJ6xIXb/vzzdcHgWNjNOTsyBRIEQ/Fh1TpoF/EhmALvCZuIbmC27klPbSildwL1ZFhyU
12zUW4qcJbCnlqyVE18E1cakL5AiXiiom3xX0aTPVxMxBzewdru/orgwKCiqGQyqakUC4PSTZKwa
brO69G2ASpltcbR3iWhg6+dR1d3MAKmov51t06Y++GyfoQaPr2KZqiXKdtR4VOOy5I4hn/nxicVi
hQzK/TM7vs7MMOqgfQSOuUCL/+VhFgs/bvdoBXCKFrboCJZeeZG3m5msxys2d8JTVgu9JNL0owb6
ahU0tLSRKDdP9iWbrofOgarwsESUAmq6IiQDIeNkah6v21lc4VsmqrGXVblyaVkduVFVPmRqcCte
0/cMfQmr7seLEZ8S9f3jknT2XvdtC2e4v6dckzmjVEIABxk7RvGpcLEcsLyT4VrvWzdGgKMGc6vI
9x1jo5vQb5JeUVvNexMKzBbFCtR7rjQTgBaSloRot01U3tR2b/w0J6p1Odf1krfSiZxTCDm+z4km
RB9cDX4noORyZPjleIlMcHqrr4I93PSQZ8h94DGdBkE/AiQ75d7BzgmOfd2AZW7AiNQFGeapcXVt
X0o6fTEju9GpXkxudBziHZWsRcTm5DAHI4SbmfPUPz1tpw9o7Tv5grNAxMuD5zbAyKxI5WNgU9LI
lxyj6FsiPOvCtO1+h4vuWRxKaL70g7khJk+rcy+M5OCEDqxiyx2O6A9O/gz+ozOaCOvUk4dC1wEg
Nd8V2ggOaqmAasdS9HWMHQJUOUQE08KXOPqSyCC+bnNkUIod0EXe7i6PICgeqvB0QuRSPdvk+hmR
yFa/N5f2Hyl6SMgnTjLSpCESoA6fVPlzdD8M1KmpRhClGCnS9z0JYMoMIrP5QqtwH0e3TRGX9r2R
GTM6rwc5QnbKJ3hO26NG/D2bkVH9HHjeNMh/kjRjtkS9wWYFSsBElegxhGbJyprvv1EFP4V6s3qv
wMN7ZYauAFg00+i0DDqcX+v/LO/fiZ9tpAayBQzuGHCmv5HO2KCjHSFkraIiZjK524MH3D0wgAHG
AjVlvJM0QwH3vcW4U/sHM6IUh+c+yfN6XHBsQtsjupwuRBEpiSQcbjfbGUQxEBaiFZMhZ64nSM7B
ZIz8s1+zdLIXmHU1M6OKYeAWK3FKAX87Xln7+EuMaZuu5WR1aroOYWMKip9ekOcDyyPzcvwlcjiV
wsd/twn7NTewCqBsxdkDQBNn44QkGMaD+YZd7X0fPxw2WqATTpE1udAlHrBD5heMAyI6gRw1QDih
7CLfIDUrSzcSgGs6gKvltM87zHAoaiytxgIrpaHjs52IHEq5dFXV13ejHw24rnox94QlCu13YT7j
xZ3CUrp1MHDmbwwHyR46NFWE5ZLcVFP08LATOk6kVFIon9fqVUy1GDXhkRQS097WkMQMN2GWI/w4
wGK0kOUwrGeG4kvFNxOB6wVdM7gZ1gr7QVx4bTytJ/YSVQAX1LMVNwU0XDWgKMtwzBFPrwOR/gZk
++BaMigXCEP7dQ41xJcXNWsPbxv/o8s6qe6V76d7h3Ir3H1Yzg1tWeFF0nzcmYEkQ+Gen+0d73m1
n0FHWWbBmjs8XHKWrkLT68Drcc6H0/NAppANudWKpatU+3F0SWtzpwjKvDuPTd66/A8Q2gTeBE0i
G4GnjN6Ce/cj/VIG7nGfWiGVXh2Z3Gxs3oz6DA9OVZAtI42n9jAEVaS6Hi1XPr3rj6qbYFRkvvCA
Qb0zb+r5B+T5vd0J+udSkDHSyoaSFkVerh9ZCl/PoFQGkjvyQr4O50/0vnJHO440kXkO8WZhLH9A
5WXv46K9ixoi5H7NiJEtF9Rd/OF0uPecCfmKrN20BQ9iUi5n9M85ZsCjObX5+iA+/ZIkExjiWwfb
7AoicWC1ggsWTeej+v0q1E1HW3BCBGuy3Nuv04serniDpRFEXyGGlslTZDFh2sUZym+Lv0eIFy5U
wnAghYrG1B8BhFz6Nr3EkxR6H+oN6ByVscwCrSODQXG2dqMpI0x960bH+t7OD+eQ4rZW/PZJqC1V
9460pPWHxnGyVqD+uh5nJ8idkPmSazRb+8HIZwsZ12M94hQhIn1Xy8SWB2+cAfEPnaNI9k/t9qEH
wiSyjbW+tP4p9yYWH18+fEd/8U34oQ+cu7HrVvToIkkIQePmlwsBDbuOoXTo3azI8QDI2r83pM4f
WFVBzZiupJkWvD6TNaPlic3ZElgfeRxDqubbiBbaOxCLBYru8HPnCU8a9LPqCvS1AHEMv7QWjrRM
O2+x4va2Vw+xb1PNbndk5eaaxMy7XkNK+UZehufKoZiOwrvHEeuW5SLRAgNz4U5L3qa3s54SCHJT
Yv8PsWgxJDFFIDZB/EqQe3BrA6vV4htqVD3jlnGetD+xt6Yjz+6X8+cdhDaKLRj0C/iCF+wLPmez
8dXVI2EKDAPBZE8PiF8Tzss+7YcwcGAQdxibLy20Vbd5Vd7YctEMX4qzRc7R3muZwbGCCuMLrAff
fzBeD1hqz9L5rV9+3Efh0bogfN72NTFUzavNvP2PGyJgD8n6FCUPL4RQ2fwSgWWZE7Z2/9JsYo4C
fnM9RFKKC3gH58CP+Kd4vhg/edW8lr7SFBp/6jwBHyjeBnVlsSSDYB2tFf+cIha8Ooa/k28iSn2J
cF4zvWvlz7qYt8GjOk/ALaeTsQHACeIiuodjo2l4xmtpX0X1wJ1lCe7vX1opLA3I9Lc4mew5ewoI
JwaR2dub1MIArmSCV2e+5iY+B9tVnHeGl1gOa7Ejr+PgjHBC6VgqMVz2cvcCAZZOnI3Bhbuv+LKd
IQKX44stgF5fxWJ8dxnwmOmo2sI/70UB8dOlbmB1UTc2xuIDj6/V7/06OjHtdvCHEvfTZxX/INzB
AKvYVAYUjtDalf5DGSlPlAjNhCpJAAt4G1sPWyg6EbDj4cLa+Zm+6B8d9EFWqI5MLgdqTlRiOwvk
Rz6Dd5I9zJrYzZypcR0RyqavTnzF5gGlHGG5Yp2YykKcTH9s+b3MaD7uAGMtkICTvRow76dmv14x
ebf8LgRVTzrUO6x0+8HgZJoXG5AbrVxBan2/okEoaTlc/oVfgGoepLJiKA504k4w0Bs1PDtWgrpB
wQbpRljql7zkt9FaDZqNfwHmKpJZ0HOSixIG6Mp7Iyc0COcETFSY4Nj2Tx/05XYttrVofVqGISps
GzOnqI9OBrAtkDs1z6qTdhzz866wKB96zdIRvV4Ia9/GNYKPEgzISGjC6EcXmvilX+hq0ZlEOD+m
Sk/rReFuga/41l+TXRJS+0zgF19jQxtK7P2EoR1rZGE8pVIkLXZD3/BpIXLfWsfxIwtJuAhtEExf
sWnmESrYwiQBI/jfzB1PHL6GfXrOn2aRoHb3EzWk/X7Pmf8Q7dX0xOEnl6r1ERGszw1RZMpZwovm
tyebhtUKfrCdhKyXo2p1DhronH6mMcWVA5n/YK0kjWpe+jPj5o7qQbcKkqrBz+O3vTr+h/K9mMWD
nBP0fXiaIWDpfILGlAD/Fypk3hBkzKx7enR8DQkoR+w+oi2e3pxccF+4zdLEAIUjg0J1I5pkh5l5
3AFnt/V+ppCvVNtW5tqChRjJVV0QcIxa8L/Lcq3zWvbHI6OLMsi31pI9vF6svBinFtWnZ0M3RTms
XB18AAh1A5c9+782m+ayBDOtGOwDQzOHMmtHz473gmCqr+ZT6ZQHs+Fw4tRLnumg1FrRwtWxjwou
pkxmXAml+uBiV0k1xj9+O6PjBn58sPejnb2jEX3GTvVbXgeTKfkDTk7FaZhhMV9BGFEE/MFZ36wA
2Te3cTfp51NeklusVS255Urtv7pMN0QvodffZfhq+bX0REnbiFHs4UkPZkozL1ob6nPdpgQMtKfN
NQ3FcSt+6RQxNL5CBDLwJXiSVyngaT0Wk4K6pWHlnabxl8pJs7f0xoVaODxLZS/YzS7gwL1KLHjx
JOZ3oqrWc02c+ViSRbDfbsaw0GH1nVTtlxpDa3J+arQjgivcO8aXk+/9T7XsKbmoFiSuJwdPiS1p
bdI/ZRATRoEBkuhE5jigUIuNoEKOhEb1BMtKLx9dAgLiPLK4K2znokFIWdooANpsnJC3W6L2qs+K
K7vqJe2N5FCYyqnhpzkduMFwEuGEJmxKr3DiBHkZeyTLlBnIu8l9GM2783HbxBHBXhw1WBiFMR9W
p7/LD0ATA8udmUl1yNsx3vY0sJtovsvpLizzC6oSR9/Xeeh7WdwApZrzFIrRddrGtZwllK/UAmJ4
z8szkTivS41smWrrohXmz17F75i9YsGSp6WQuM1CDn1ufrR2wNZpPwigEr6ZLHU12jHQP2VNA1cd
QyvaaIMwlWrLPUne1oICjDNNycLByYnirSx+Eu7qRXflZkP3ooAhG7jQf3qDAMXxX+5q/j7fcygt
oDdrRx00h2/ef9pWmDh+qw6eCacYjp1hGPi0FoRLHDOparvEmL74LQNlEWLc2wBitS0T6oGgAR3G
nc/7DRdw1WIC5o5xYolH068bn6f6yKiz2WEDVuZ6pXp6iIMg6B+BKd4yaYKtjouRDvArbsHOgHu6
rScy4be3D0W2K56PrX+Vlm6nL0Fk2FtlTncyY+k7dM3wdA98w8hZYS/K/pUHQkmiSSJj+6LHD1/g
fCXHL75iGsQwCVsZErBafV9xtBHZE+2XiwETQ9WGb9UIjYLtL6rV52BUsyeXqQav8ixG0nEpDZta
s3iwiALC8yk1fCoFw21jeGjNgBqt4o1r1g29nqT78MUKrSEPQsT2OSuWyKAUT3YZUjxd3HVgITg9
ZGQcj7DtO95gfJa204gcH7daDNPPMfhUqdPfigmO4pjYyaR7dDnXpU+5wWEdj++MsgnwqGtrRyh4
HktQSH9eTrAA8Frdd9pKFzWeIVxz6rG1FJ+mwsuvuP2JQHKNKE2bf0sMV3AhZxQe+wHSkrP3+1NI
UAmJ7XQxNqMB9d3y0m7AqtyTVOAEQdnM+k3V3kSmyNAV5lqohWa9NX231JJzcg9IFxo1ENVfh99g
t3UHffmmXuCbIMXsYHPHZsyqnKnksEMEOCFBE+MicZ5JKFSKgSxEePaRsJNM0UK15jg5RYIqEqm3
KM04+1va+duPgkrDq4KNc4sFtbXeFeGR3HWZqU6oWdONIPY6hpo4Nw56UOZqjBi4kJsPl2sEgeP7
iEIQcyS2C8S5yyXRLmmgwZABFUfwkcoP+p9JoH7UWfXZgZK3TNU4bWri0OgeNOAUQM0JCR7t/nWJ
9k/48NjO0L6GW5ohffdlF3HEo+G9WCrwejObnKPiePzAtqspiH/cCkI7qmLzKAVefED8RYGbovQ9
MDnGtUwwPqQgI6K6w/8rxiaAybXd5CLpWwDq8bzpNmW4ZXZikU71BJ1vpz/IN2b3CghN2g2bweQf
cUrZ4oPc8xqtHWaTje3/Vr7rUyjHaVjTSHayClxiX/PaYxFNzhYiVFwvCBxmphm8UFRphG2Clmjr
jA5ztu4RpW6zGbQSeAp0W0JZMDuglf02Xe1Opr9U8MSvpt97TPm5tg4PWc/GYHHLhOIlz9yNYaAy
QBWmuMeu8lM3L2brd52XkRH4HwX+2iXp7k1mMxlMR26U0sWystB4vb3OgYwkySy8I97DuoKq+RxM
+112Jm3Jqvz2+rvrgvVcUhZ8b9NNM8u7bJ+9/t6rhBvkUYobps9+r0KBiDmFhzNfV5O1yoZRY12+
cL3TLy/PGAVGrD4VXUveEuaWvRIBkgPWQ5PltNVpCrU1rHx8vAKSA1NsGKvcSQV7vyVpMOjAZ8et
MBEIBbJ7QXA75l3X+UZ/9MW5FqCnH465iAvFfkpdhUfqBYIDMlx2TRHi8nMmpym2u+JqJ5juLBcY
ylRU0TSrlypF4zKGXHItCF/UBDtIStDANRVmGSdemRVus7tJhkiuDua9vovLSOobhWv6H3lSQTQz
jRjBQshC/ItEVs1wLLCERIz/jLYC/NZZZh4vnz1ARUPZunLCI9QYbGUgIBY9+v0wnWQAO/6RRo+j
B+k4QL55jjUEzvHPkEgWK+PaMFtLDzwr+tr5ylpZp7WUwjGOSx+t5pZr3eOm3jolVXYBvZ/cXgiW
3f3yV74NYINBZ7AD+Kt42iduSPXLkUxUlJUH+vg8F5fr5yfXSDblcFiAi8xCBpoF0nOPhYi8BG7P
h5dd+4+3C14X0TH5D6u/m9D5h89w01zsCqVhOEyfJuhxrz8IZV69ONjza+HWKizLcFkWQ+3f/IvI
HldNLZN+Q+kFco1EP/UJt/Aig+OXBq/6b4tEdrxIxZjaRDJqRJ4UABHIaunVXZQEQGfIAm0FHcY8
+tYnoSDrL6Rd437gzwze0bJK6Tn15XMSA6azKIIOiko2vftJ0tVG6Vn9dLa5I5HMd5bEJF6v/g+i
tkekPsJ6lDymA6Mu5gPcWrmwBaoU6j6efUnpNeig9YQG0cMPT1ed9PPMfYXV09yoaw2CkuWGrASA
QJuPdDwxU9sCIoGSMk+vIf73sMVRm3swmTS9M/Pbs7g655CT2C6Z9r88OIuUBLsO+t9EKnLfZNDG
hwrduI9oV6ydecGfTv3sCOoKAzBtO+Be8HmFmL+79mLTSgMxehVSiOQ4rsYwAsmKX4W8Rj4XlrAy
tmML+Bf9qyjwW/X/gYIJRmjYO14VSSBzWlcWxUIbDcnlYMVdzaunkMYMwLoPCeNUpTmJMW3jWKjJ
gst1L11C5LUIfjDNoVtoEEAwLGZePRXlXjCziKR2+BMLP6iyosng5gcLjBR1FlFBD+LZomi7eJwu
cTCVTrx41rrhFUVrsSURP7dViUiG7wbEt8rwUkv5w3ng5yutkLWnzK1JId9lZn15DgP2adrY6IQy
RTkxzbVFfhAyW+zHIyYeiBLAlQ1B2sczcx9FGX9nuj5yfJmIuOdlFhDZLD6klTqIAVSmjdk2VwII
D7afcnvAO90LVYC1xuVcO4JXTf9HAHPKNvbUcng/Io70zhewkR9HLp6A+fTjW8waphwHsmb91VUy
dSelWoNCqLK6xqCAOOGZZw/pdJpi2x3LiFE7108Z+lN+xvQ1qAUjSkcOOSZSoq7Li+yzldTAIYZ4
i1Ao8Jrss3bqKrY1KfWKbrXaV+fErY6l2bYa/CVb3qrh151O/Yqp7EhAaynh76YMx9ecDbEpUqAn
ZKOyUSs7mt5hB6Mt/1wUIVNTALVpoAJoOZwAKNiKGg+URzRL4aBdw9TxqTY228zz+xrKkS+vrQDR
iuHQK4QllpRuntF2WrNqDDBUZbTZawUuWWWWrnsc+IA2Ryh4jrnIBVw8V5jBCgZo1aMvXtBM5iZg
ipfrwv3OagecFBv2Rh9RWZCYBe93uq1nlFtRxXx7jzGncXpDEta3zXl/59hVl2BLhbnzFXXDfvvA
eX3JTOWMzJw5/qtJ/KXQ/7+CjD8tZARnQdiT7YzgCnC9OFejfZYE4Ezgifg5MPjGiMkzIWAafWYo
kFKsXxqnxzmITACsSstF5/tO5VihTUAL2TjWr9MFBVxMfgyFTqfmSAxs+l+PTUHJbdh8+F5uidLF
MwgZtBBkThnI7O7ItHeYPRdBhJXOm/eeBTBTzwijLrOsaAM0aNKhmEKzr24xfzqIg6LeHEPf4MT6
jrhENg+BErRVzMmR7R3/zpVAufFvKAfKe55tB7zzAkiHZr9NfjZ7EZE+A/0WYVnFxnXvXKyz5j+g
dYgZM1bz59F785REZrwdjTR2lOmpczkG8cr+ZJ8vN6TsAswP2hmkDKlzqBJVYvm6zWmGmQAYVvtf
y+C2gEkCI4c47ASx4i7MtRpPCRyQh/36onypSuZX1vmp6dweqn16LIApLFErJxKj1Nbo2AEH7+a6
Pgd0/bFzHC4GBT6dN58sVGcH+05DL84BAChHxhWkpLnu9ZMjGbCfGKXGqUs3ZtFucI9GX+xYSsGA
WMmouXcX5Yt5mc7T1SA+vwC7BXdavz9qm3+LTg3vnMr3tJe+w4rSvj+6oLcDnDvIdZYbrJfztkP9
FKWrqnZyEUg+2Q6Lmf9ZZlq/20VGDii9vkwN7OoLSPLzSCgV2D2/s9B9qNgb8BZsq5+SJj/rJasE
secL5ba4pOp4Qp8o7RhsRrJ6Atu/pcnpukNWoaJ+UXQnlAhimG4wjNfDQxC7VoD2Ib7Ev0P/NCHr
h6l3rGAEjGeFksvnS7SoVtNXa1VvvXZ3d+3hxnSV5RsWT+AzQ0SIGkt6dXZ5N++J7GMU1tx+9AEw
jLAbYIDTAKC3vxLe49PdrBDHKtwciZARVbMPwnBFs4hFdnElqjlKXZo885dkZ5qL8BFR+w1z9L+Z
8E0M1/pwOn+kr/Qvt4q8zNYpIwQxM5wmzztenjWroGq2xy4GLOKUlRbeNIpl1wRrahfdV03qSO3H
kv1px7HaynuaHJFMrJPRpsnZDm7uxAfZ9kxLQpfes9ui68PT/O2dRuhLwdSUbm5L5U0hu1U8awFS
ElopC+cvkbP+BQBxZWRn+ykEqUkeqItn7etq7R4NYCEth/JNC6IWUAAnlB8EyEN7sL8RKndSTUwL
I8BzK3masUj1mLgTUvwEleL2dqH4oFT5ckjBeU/2xBgzXvDiFqaiQzMgYr8PjDBQFsSgEeXiibzP
4d0sGRhaSzTMKWfMPXXE/IWFYvZecPC/MWXRItll7qIcSqWowlcMzGjUD/2MB5RLtFrw3BOZCG5z
qrMynmuya2CM/7hR5CGk9YCSoUYvSh3v/uKxXpp/7nwoxqMKHk5kv7bz8hQpPrI2c0QKP/OFw7wE
nvI5XSeKpQ8rDIJ+G25L9IdMEN2tsR/fTuZnZ5V6NeAAfM4zCQdOZyjfADo9jsA7V3U7Y12VamAj
GJ0ipztbilPLCPJ7W0JALlqF9PTpshOAWACcxkLqVJf2Ofg55sO2rda/SKGO3jm0X53I+CtIFqvv
jTty2yB2j4XYkc6b2cyzshP2ZJW8F3bl5ZDx2VX0XHxgIJEaOQbi1Q3sZfaDeOTq472AFNL3Cn8f
pF5qxjdlZ1OLHmeS717FsnmQcabXXkiLbsLcoOJJVZJjdBzoP6VdJzHvsecWVmiYsmxgLc2OWjxT
ei8tVbFBwRXZ6rpIW0Y0wcdoXHvohjmGTsfJBSxb2H0Ofxuh7NnRK/678GRRMr6YW9AkxwrovRf8
dirb9qHmAutxk2ztHq9jC6Cg6bswwn+iHK07DMZA2Bqqqo84DVIfCFPsCJ98ZiYylYAZjuReF6HG
Mies+liMvZ5W5iFg0IbWVO636jPHDbi88+eLSSZ7LHbYqSP7dfS1/TMA6PQUXzf/QX3mhd90DkIC
2ZA6imKwsO00jkxOI6pDwuAaWvH5h6fhpFSmmnhVR6OFcFMMCylmZ2zAs48Ph5ZnuQIKGPnplzoE
HFBwDtngDQn9hWMcCG7aApPAhQT628z0hniCK4z2UsiG1WL2lXjlnV1xWjh/OrIFYyBwzL3u9rqP
WPwOMEpC06kyOn9622KQ7dO0GFlolvnTZtYqV7F0RMpjnopz/1vxS5EwV6daTiGrFDRB/9LY61Pw
KcJW3R2/IMdHoDMNB64cacPos3rn3ISGowS5AcM8fL7I1hBonFFaMruHuYQcbqHv02LpPEaxt2pD
8V6upTMLeOxjFQt9HVQK8fqCvDp/Jhjo/jNyfbEZPR1ZTsnIaRFwPAUMRP1WDqt/C6WfYHgA5YnY
ZQvvKUf971GSnfShb6TqlGvY7T/xPWbZWC+6twbQyDjLnPgJsxnOPdqfl6nm3rAx5RgQnTu0qY3J
0vge/3TIGYjVF52duNnGNFGlOHG8wj/IwzwcZ/K4uznAPgm7m9+yddp28eCw1CnxCHjJ+acp9WY0
D7h9qREUgWz67GkbUb1NU8D5R5MGn2DLmwzZH4ohlEIOFsI6UHOwcBnbROEjCiDvWGoDPP3ntTn6
VQq6PSck8NupNn3z7BfU2zHNewINu8M9tzGBapAAE+gLXWWYg0d7AKB9tZqEqLXigkMwzj4lJUyt
sg/sRmNS4fJmURVSs/A7cNetfcBddPYI0zcZFQWxttz3b6/rJV4lEeSxEAFyTci5/JjJpFp+CIdx
DgagtY8X5ckpO2C+LX240BKNAHcqQs5++m5sGkY2CXQWZok1kOPHFwOXy3tBS4uVEcy+F+wUgfsg
6tVjEFciwNy9E0KX4iqZrs0RwuQo/p39z0281xqs4SNWsQeyiumhLzswz3bydpFTdeIpsFCD23El
Wmu44VrK/lSWgQXxMchspMxUuMjFg201Ax9FGSA+YSoYzHLASafaTLwrLsWSdHs/TvtcKtxWrtYg
IX8WlGdRrQ8Jvp123l/+0uB8JfaEsj1Gwcm34c+NnPqQRLqlTtagv98/lN1gSJ7bUHQNTAdXmAAR
E7nFhrrgeKnyWAA0wr40SE+yMO89x02rqlVyiRZR2dKlHloSW1rW23laAoRPh4cF2PBkboQ2PnOP
jivhY8XAq7KnZKUsfvbt1atOpBcejFs9jWCnxYtcXpDw38uWouEdnXiwSIcJqCsV5lGAgLHCEU7n
8x18KbtLFHmLQHxxAx4/043XVqcFMq/4WUdgb0hADhlgNw4f6QqtL6TKyb77qgUgAOUdFUJvtOoY
5/5R1XmqaI0D8G6dPs4FnwJxXMQcAWpRrA99MeADVwX/w+GfHKrlbNq/kjWKeexsXTgnNjRDyBBa
c0+aKteeFl0KifrDZ+bXkJ6625VQ5k6D4zSpqbAR403clkabAsbkdx+dj8OjQ6PIY00ikodimwTv
wUxoaE2kuJYN/6zXDAxsZsp7g/N9DgT796KjE2XsVr+YkNY8r88EM32K2q1VvS9G/k22wwV0w412
++vwnxPxvbLi06JSDIBz7is2dtx8DfBsblX6JnLh/GI/kKbeLVrrpjg5Imv8VhWCQ5Zsvx92zaEs
Xis6HnEwKgQYnesUX6IW14dHF2sxn0WdPQ4eIKjJOX6P6ScCNSVdEExAUpAS1pxQQ9zHK8s4bzVN
YcehUnDDT1+xTINTnrUWOYOpe5buY9GeRKIBPP2soCk5f1Z99qOPhRGfiHgvx6g2xNGoBuB4F1KK
s/sEQ/kRDLbZR9Lpn2ZJh4qTSDj7gbE3Piw+xiPktpgbB33ozfbWkFwExeqr/Grut3UG6yYesJjs
craQRkY3wY2SuqphZo7u+/Q5JricuBXeGZXqPj39Hdp8VX3EDNpWD4kOVlCrHUzooR+v6v86RUaN
8FGwyBI1VRo3A1EmUtwGyyhWcqTf0JuMt99xXYxs2ClN5ISojaC2iysyr2qqzQ9e0F6VwNKZ4yoi
u2qKJ9Cw1B5V1MrhVxK7A9BYwumDMQKIk6pBC2Ut8BT2B7ch4HWGvMYSkFn/XiCPNes4tTHN5nTd
7k1LogzogrWxdxr5cPad20ooZAir1pIxAMPKDSHVJ+SttEoRIp+VchBVYo92YdpCAjCxyFgu7kVo
WgFBKH79/Hv7/i5MfylXXCCya6Hui1jySmGcgDLdR5/2zmGS3D/xEjWyMdvmIw9WJSrnkwD21mzK
GNyR+7bSH/XyIJ6Aa8/vlqgEhJsanrUsHb7K/vzr9QrpSQF6DRCks+DbjIph7ca2SGJWr4aC/6fU
L30mDzZR/zA0CI0CkOmbGsspv/t6GTknDqqT+wOD4PvPb5znO8ZbYNNZs3kbK4vb/DePRHfFPNNi
obMyv5y6IpaH25jjNHzp3t2dF2SbjC+tDYP5zOiuobKeT/CvYVi8yjb6+v3KYJB4uRQ9D0CaMqvn
aHv7xDRMKrf1rJBc2FSpgTKvScvj4IQV5jHMpUu0UolG+kuLtaXjEQCQiilpgDWy9Q5p+JBGkQxy
gKDLYgY0M9Pas08YDbpE83DTPMiypdCs1qQaN3Laq4tIFk7JIFIUmvbRdmyzU6HXsTV5MuU1eqNQ
TjflTTg6ZlWtdPHgY2qYd+jIBdQCy3wHSkcxlMV5NKYjsqthnPx51H5LyvmWi22v8LQEzcP79QbA
gRLfZ7lajAcKC1TOZ72k2kRUwN4XqdTC3ArQpzGAJ7L49Z22xGCbZ2b2q96jNIwXbVpLrsBs9ikg
GoaVwDphlCIqsKCAdoFQBDoaGinY5TIr3tfO/DkNmyHnmEkWFn3/wTLE3tpz7FmHt2MYBZkG0T7y
FQC6ZQjkuY4ySWPVkzt/9pDzfSybpIUAWJRnxgPlfCJ4CFSxWPVeWhzfyE/7IGyM88/5Srp6I/ts
96TlsFbaOus3xlbPrw5R5DnTgatDZqzTOKoDtOVFdmLe6mOb19bHP3RCGvvtDAuEURIgU5IxLotR
ssiLvc7ZhVdJRAuBFkix06mUaS2NXmwWuiIBIK9tkfGMoHRkPwHnqdbxG19X013lRTzXpUP63BVM
A/WufiPzrNMDlvaG9SqJP0VlUbFaj72aOChAfJci7wGwYgBWESCW7bssncvVt7pjVGVqX53XBJXH
yW3GTtuuviUZazzZ2ynWn9DWiTSoufiesVXhdII73b+VXuFPJrTqUHA67WIcqx6AufWSdmrO8oke
0Pcp0f1sCwmgPEn/R12kcR6VbHFYkcSu7MoizlwTH2VMVyApKaJjOMHEP6fKXRJtQ606DKjLzaYg
BQhyCe/ow4K5TN8Bqqg2UDhJekP03LRHAmUbN4ztfRTjqupi8pC7TkQVNJWN9y1Ob9KL2Pl+OCrt
V+G4t1n/Ylvz9WdNJacV+YMOETKcZ4ml58QAQRknEhLGxv3qTPiuKwbk8TgYiT55Ui2gmPlCZu97
qxYKydQqKia+6gKoEM7/sDl0i1qICps0SmC5DwyJRHW/ObuAX/NsVZXAAh7bIP+Os/X2V7FZjK6f
TedVFbt0fxELASrjeJL05s6KAodwIiUQuuLgbMuc/98jsUfipaL0kT9zPzHxAfx9sHe5N+QmQ26C
saT7F6LVQz0JFte8CJ7PByQOpA5JmDFHPeld7yhLeGngC2UJ9ZSofdR5N7SD4UQvyHOvoCTXCh0+
0sHk2DsWo2IFnYP44QIQ+3XdhAKbzo3hwvcft8aY9tmcDxgxQTFZ+BIg2ATiN6O2ujrFHbeS7RAJ
8VUQf2FmEWIBAeRGDo9erUb0bXiED3tNV+joEEl4hCcYTRLcqdNghDFtYD45HdE2ArUkJSo5WOG/
CMpMKYHkOqdt7lcPAqYq3zn00y0qXIwU2lkaBGz5Vcusdq4/D9GBqmfXBPNcaFmkfcnKVJyKLl1i
xPrBCt6KMR+pAiywAfHgmvonnn1RJJLSAyezBVSg/udtHoGdKacEUyH3GDBtxCGm0Paa+BbIttzk
/g2nsmezeNZ2oZ1jnIoAHnVQp+NxT2pI0Aw92Ig2Tr8tbPt93MjeP2ranBdyatVTpr0YCngAlP2S
ToNUqvtoQUT5nJqDJx20SgN8j1QwHZLKzR6QjzgOvPXJqUNUO5Knc+aSX+bDnPb7rOPFZ7MV6Mtv
PE+8eQWHcAIUlb+PnSxzD9o5bjF/w9QAEUFS1n75PTHyksyKsDfuatzYZNsZ9gu5cydoamV3BIxy
Bp6iYwCrZjTNL2yn+pUAKAWQ+MAO0QwFfVqTXXAhaHutGJhxM/+Hr4a5Wbm0HQzVZY4B9obogPgR
GMZ2b14OttMZDVJGkiiUz11nwVfx6/ALci/eD7UCoVzU3eFmA+KgQ1JA9Hts53WQejzs0Xu6NHy4
2CfgryqbjYROfMGTuUZ/MitG+6BvXEulzERztBl9Fkw59IJnJ9faQGAxkbyNe8cnV8AE5lnciAn4
0WFb1rRqAL8k3DFRw3nRH8M3p2Vrs4HNyzT8ZzAZJJyzCxVcG5Fj1hs7t/q7GDB6k5pQRSnl5vBZ
cF/oCdYSSV1f/5W9SWc7yQXvYOLp2u8/mqmQ70oXop6jVS+THpLupP4j6RO/PTfJ+SMJtkB3leIJ
ZGy86YDiL2J0kaXx/Y7GHFZszvCMBP8L1c/kGPwr5lutNuRSVW45cxSfbYW38Rk/gbpgktx6xh0E
/qliSfHh6ZTsv7xML6lG/EHQxxYvvpMi/gg0fDNtvAq3sg4Bx/7Sc1f8Lz8wHuowNlFaBtzTW5wZ
PN51XIPo2OEBTQ/hWSYQYNOPqYNBhBQcumoCPdvWVp2aaq+k8w9QSHfTXkiGv0ICEn3kaaPHK6eK
bLinN+atGAoG5v9+Tm76h+s5KpJFOF4TLJKqFyZIEIGfc++BZTsezHcik0rKncYgrWLOs07l0nFP
xZp6nIhbQWUPnmtZ5hWPINiAV+rVPtF43eD6A2zLMO+LwwAhYJRlpTwbx08GL/F/0IsRPELXtGlX
KqPT2rOa6GeXqiKgYt0QxYrGTPTNCr41TV/OsKOvql4xOmS4i4iJOVuP/gfmOJX4xXdoq+1IO8sR
C5u/HgpjZbSJfKQp5acEkKCG9sretAIsvn+hKFaErmLawokFHOPhYxfK9CpNllkxFmY+bl5X0qgg
daayq8sO2J62c5rr0Mr8N7NP7SJIqXEP7qsQ6NHa+G916VQIS65MxZLvhfbPdcclmieM4CIc+yGP
QUuSgZOudy524EyWFdp5PkspBwjpfaSi8UBoSpQatE15XP1t30LPz4aQg1LUlHUro1iCa9u1Jmk5
hk2soqK9pJlUt1CI4hTQHT+OjX9vlbfE365lnr0S73It3pOBaprtHb3HF+TKJeplGeT8Qq1VYvdK
jT88SzFNS8TooA+efNC7DPUhJKCfDc5HnR35+wJxfYwef6EriO9Y9UIn+Xz/6QwOR35/dcqwuk+a
HbSC267S2HX9duIzur7FYZidjKJmFIeqhkB8e4dyKWPfxzZ8EPecxtTlfqP8oq3oeoP0ckQU6kYM
J0MOCTvEw/URmIwkC841jgU0fRttMU2IjftVeV5KBrFjkp5h30/35lJ11GYRZCEtI6LejhytGk60
SgyjcJ8XVdj0FUg+YsXEIEYt1jDu/tPkks/iVzP3oH+xapAn9svE78xsTKJJMshLj0MCaplZZb7y
DTvanKSE90xWhacYHspXmEH1V4tKEeswy6zruT0aeQpp9qxnEb1PJ1kZuigMtgR8QAIRYyafzKoq
0azk3faKvMMzSZbpxfRcTeIvP3p3mwfdsFLblb4rrPgVAgOSRZILdjGtx3LHMyd28XHa/FPa8JpM
j/6jNXJPO1m8oOLiS/pIWPIInJGaBLWfPZZHknH12B8fSlG0Jazk8yCZt+dH3RFf5Md59KlU+FLx
1tpKwoLTxdFMWyQ+MT7vlWPbyNgze0LeBBhCzpeCHaDAZgqkL4Y+IqtxRDWHS9v7KkTy9CGX4vWY
4ObhivVrKCsuSOtAj2cxOjWdglN9YPp0yOSB5lSHIbLsbuxgX9u+MNUNGuklembSaerXTaipl9Ju
92pQJ5+3lFK+9IOSr+4pPfVcv2hguSAzZ1nLGUFNWf0ztgG8qM6CBCQpFtumYKHL5HIGTTgvl7Ee
HvUwxC3zA6COjxPya0h3PmU72aCyfYzG6Y92L2f2MzA7ExB3pyqhm4n1l3lh0EogfBAb23dUilqr
9fzc5vnBhwcgXipoWbk/AncPSqgcuTJYETYT7C8D5oWfo7qF03vLDm0hpl1PaWfggniedD0qCLto
CdBOF2AZUWg7PZp+UM55JQ9v16GVfWGQKjueCDUXD6gRaYVtdhzIchQr/YHBG9lov4hDACg2+eb6
vMp+QtPIugDEzCoQCluazuhwo+e0/y/V4tLWOrUQZyzwbf8/p3tcejiM2uClSRkXeAolbvaDQT74
1nMg9Mj7qJgJ3iVLUQzo4lcXEOK0oTj9/rR4PjzVBmspeQfV0O3EEra+O6EwaZ8nwr9fYEl0osPF
nfgd1tohhYCwOamtpJeASjQxoJhkVQOZx0FgZktPr8C9rWgSJu/Xcl8N3DKfRWvByxrXALmuqc77
ta8YbXPi9R4PadgDc0EIFhOaZPirzrYxC9LSfrFVV7iBKIFlCld4B6a+AigpzFdQ+8+LDsNBxX8v
6YWWONePM4hTRCeiLEpf3xV2Guaje7DuQz5OKOhlyFbCAn0VQr/tjeG+w97LA0HOofMxRhZOjxgB
nvkdRng0xPUyqkd3tqZTwukffgL44PVbX0XjFLNunBDrXsYcybFVWm3RVtn6vBpsbhZHdDOLADyI
PWeCvI2NPqeHPa0dlkGNloGjmsZVtfWMfmnVHJU/oaoygdPZLhTs9UG2FmwwbAAg2scnDxj4IqGg
xfpZyn7DmJysQvAqph8auCDO0UCQKDqn8lPWE+nZKjJJRjgzoPWaqMH32dS6w7Swl5VzDcptR47U
Gcgn+gHVjsxYsnU5IcDDzFilEt9HHBjCLyW+5FlF3dsMW9Xynj0YPyfDteFmcBUqVUn/jbNY24X1
c11EGpf7kyR/Iy6Qtr1IX14X0xG/iZD4FUCIMJis9LSelvDTBtTMOZvyEenaiKbBmeebIll9uIHN
jWYc4NxmO9YmWjGCBpqfOMKGS5Ac2tkf1z7O2RYN5KxzhPMDP7RLntYpi0gD559m2XeqRcp1PqrR
cHMfaHgKCCUNIKa21+IByFqcpEoH3Obe3/neBzPB+qHCftlQIZvemQN9wBH02dvEiTXVhVzv0OON
Yqq+7On4h1WiFHWowRs4fae5Cecud4BeIOcG8MGmSm5V/80OaQ+q0lT23lgeLVlWVd9Oht77ZYEu
N2h8kJdXgkFA+4ADPV3o0M7mpC7LK5ShjtyZXQ/Jo0prVOJcZPEvuqHEd3CzgeqJIE4vsPEHXyA8
b9k039iaKbzZXAEPC3MhY1xrMKn/tqILYz8Z6O8yVg1iNBL01WR2Wpo5YQSVTM6zF0O7bHPPZsRb
HhmoK/Rq1VMNsKFsu8tT4TAxRx+36F71Ml2oMrrAbvlwHTD0YyZO223J9PU9GchuAXKa/K9kqeNe
qkd7Ko4F8mcV7JrtlV8k4v1SaVO1EOL6EPAQkTFKvIK6XHBdl1Yhx3CCDI05bpp5bCQyLCDxRzEe
KjI6nt+W+1pvQmnWQ1kIpLvjgxn+fZTgGu3Ur2EVGClTABrvP+mOoL1jn41UDfiiuKARLcXZ79qU
DkICg6JA2sTgt0kD+kB12AWTdPlkjH1Km38kMh8SVEAckVpTVfLNyTP+z0myQD6mprAfZuGlSQJh
RxYJugd9dKUym1Vk7VZ+YrwdP2fbLJloAzfZE/HUvEC1YxsHF/LM/ESnV/iYS7VRPQ/qW82Fk8mG
gvgRl88LNyYU2a/ZEdnrDi6kTGz/VLe/LkQ/MOmIB5mAPp1+EBBqs3WWEWRU86pCgNRKcNvG0AAy
X1N/iRr8HA2DAVK/aaMpqjeVyKz5TFzfTajJ9n8xtFdg51RBLm97pQMMwt95q1fgn6IyeT/qy9ZF
7oPhLmEFFzKT8qvzWjiPgZZ2TlV0T9I2mu0C//pDZXp5iU0Fn9vkpf7/Bm5JMWIEM/tyrq0hBTrx
Kys4Ds1m+xXD6F0BAQmSKSYBOXvvIRcc3X6KrS/RLOWo+3Ss/XMUiLbdm8QB18bLO9h09N4WbZhP
Up4mH4VsC4L8maIrJ+YebLrCBOXChJrGsm/GdCh6qsXr531AKVp5f4BF74ufUDHdYKbec97QdQHt
rfz4eNPt8IpgAXEu8LCjtYG+ENNMu+Y0O3wwsB/Zt8/GMIPYRIY55hSz1o1A3kaAF+7IvyYvNPHe
QVqeZei5bd3RieKwXZgOdNFDgIdHy9jbzIWiyL3Zx3TcpQ0qLmnQN9hP/jF3/rJKnzdcsrmO4voY
YFECVJPHHW2eIb8Ru0W1QwDLQUtmJpiRsCMJONJQvXz764s0KLJech5c1rYLWg31GdnVfj4vxIwJ
bX/IeJK36jTo+fn4974hJ+9JzsyjRuzzQ7kHLCweJ3PQPHPgh3btbYyGgL+myLALRD0HAOM0sxrm
tGFIKk73Vaow0MkFxALVuIyv+ohCXjxz+Wv6paG02CLlMcnjkiEjxhe2RO1CZjr3bapJzuQyOmHJ
8/g9iZve5TIir1auAGDMNQAm5XisLzEWUkCjQYoIh0jZsJrl9w90JxrExeLtb48aiQqHEA43sPyx
ATszSQArD+NL8KucCVfPazHWGCEgPV0he+SsxXnHdcEz87EaOF6tCy07gOpuE41ltzECMGAXvZgg
Y68Ysgd889XoXdw4l6AGGmQT+rPl+dsGKGk3WmK6NNmgUQYMRpi2nOHfisJq406yhljmDhCtZb/M
CwHY3+ClvOzLqFdR78/dvFEsa1wpfAVPkMUZmXALYzo8lWLp1d1l7wAe/Knm+78mN4kjXvR+y8Rr
HrtB4UamkXSFA0t5OQf57NP+gxdR9Hn+vGUADeG7joiBQDp+eKjNcayRxfr6zjNFqTr58a48AsQD
sB85yLmqaTmcZc4DgFdnA8KK3rxDv6EjXtO+psyjyB21I67hbHntRuQ6Hjfvu8iQOgtSF/cC4o4P
RBzGpdRHAs40k4uLG/jPUZlBy5AJfyq+aOAHgniX1XynG3xqRoZik9FM/+eTSbJICAcxsyJAnFi7
mtJbiLX+tGVxKS0pHwJqih6Q8cc8bEcbSQ2lJv58oWH381A1N5rGt3fdRLfP6QudTeGqXIv/Y+pL
iyU5pzjzZFShhHLm0lM3RBAeIaQQcb6vgAKNyTlsk61k9V6Rj4vX7O83xQwlgKszeNs784QLNsSC
0JPTrsig51+XhG8FMC3tJFWRD3Y1qaEypcAFapGL2haoF3394QPzCK4qwI02ah2RyeKh8vmafE4T
Ch4lwsOpY0qkwSj+5DeqCk2M9ukr+lSpHL80lcWNKIPCRQGUYHZXA1V6SqmXoRl9Yn4ChI84xFIO
yeB5VF+0iSDk2HR/DgVzj82brccuAgPPCyGObEgvNJU2jNGo5gWHEjCM3FiFubLnjbHD9UHf5sC0
6DaYWLookyIWR+Y+tKtfQNXUX3c7wepAf/InnWO3mbrUzz2IBPoq1A/Sx9FzG/kxsn6NO1XBc5al
lwiihLYzvjWKQTyV3E3rX5MqGt0zi+xwXlU6AIMfprMB5FiTU4PdSMF/3DYEE+fp9NT9ozCkjCFR
dI1Yuxmc6h2hq4M25tGLgHig3HNbjQkJP+fSInpf37lKoAY4LvE3SdIKCaUiqPEFAeX7669WKGeb
7k2+rwC/+BeJ0quYM60jZNp5CiowG0OkbFoVN9tpQemJvjib10N3i4ZD1U2XXbp1TO8t6rCFB55U
SD/h/3OV3wtUUhJaDn/MqpUbnhgSG3EN/SBY30Ox1fp3Xe9hPJN48uu9yvg+Oc1eV2ieMRug3jja
qr60I3vi2sbSyga9WcWdKDnNU0WgfQGLkNgJQaWcPUc2COweSb4Lgetn3NcZfO0pJZmtytvFmTq4
kuKZNz3ePoALaP3syxtYup3Fy3OWJgPfI/JIIFkqTZxyKrJOYvowLdCqEBo+ny5yymwkiJAf1Bko
YuoEe9tFhFR4HPthKqr2A3PQzK8BGJAvBpDR1bmYTpG8O0rdVViUwpGYkwmzZDYOYJMUyzHzMsE8
fNYnhdUqtP0wjILTSmPrpcathYyU3yZnR2GeRGKetHEyi0NSrJ+h96GhcJtzbz97qG2iJ70y5+F8
/pimzRO61b9K17yYx8HHRgy0sspxkQo02Ta5e6G0Zs1Api5s2PEHuEP39OC0kCwkpI9Sw6uelZUW
OeMGAAazGNE81ittx1tHDPghz0dJjQ2y5cQY1uAF7K3etpSK+XduWDpHx5Kc68n0iiUUJzDRKuh/
Kj3gbux75q9R2ICDl+aMvLUAPyDG7qq7L5Ke73wc1YrpMZJAUz0Kt+zQdcjxLlnxJa35X1gShZnU
Q04TKQF+LLoeZuXHswXgJjdk98uORTv7/AJL9Dy5KLa9D+0SvkSRDMsWb6YTI6RhxKaRM8SGPmyZ
bWUxGHYKB6WREkotyaEqJqhDs3wbZMRGD5bxT6VcFXKiK8h4L6jWbMOrG5gEyqf8yN14Q8nvMJM4
6Z8xDunhniOBRrE+bbZsbeeTdBOHmLaSSSrkapxeKiqpDaRhYOtJ5yaLbftQitddb+UQ/OFdgUAV
jTgNQpZ6gdXpYK9gbmixWIx0+ID031Y6ohEMGW4fl8+pUYXkb59SqYxASvKIcr0jIRIqh41C/kMT
sD3MfZ1KHPn1ygQoPJ0i3+rxKfRbuNiabugTjMC1SpRB4t39/JOHzlopCGqCHy2ELylBzYAydjH3
NeUw7xY0QxGfmRWkG4NwXzGDQPJD9AQL8AKmpd+dQO2rxu7LF4THZmJ9F2dUdR0+KZFj49nHi3yq
avE1POlpsYOP8tb2hX3p7hmRYMJXHaJJ3skbJzCo7CQUEbCPjTbfGXQG0D3Jdp90Td04MqeiwRVZ
NrzdZz4BouDZlOk0vC6sUcIg+1Feu0suz2/RJskBUBzriy3AJ2YdLHpAb5eyqvBWnV5E8P+u9ptp
+axfCrLnWU/hruMiA956R181u2IO/qkD8UvNxfC9XBwJtlfRsiKt8u72rWB+GJGgxpyquKcpJfJA
2SU0IhUXkHTzTSGcfWEuPRilMhx2wMQqxl3suImC6pIS0914/xKzhdtazd8RVhqX+4tVQZ1G36sa
evaNu+5CEQ/wiTp0BUw/9TzKpdFR65F2qmYwnNKP8zuiHQMRx8oNbJpOms54sWRd9fKC2mPgWsNm
q71XPjRJ72FzPmGiOAJzbP0GEG8Pvcgyd+/lphkPOaA8lmuaHSFPWs8ghgUmFNTdd+cli4Wdj/lJ
IYYNOrtpelva6xq3I3bUcXc1a7bwa6CW8JPnhqZ6MBbfH0uZ5odPnKyYsNMMrBc11W8sfgVsqise
FA1915dcexQab8cJrHU1tkS5P/Y4Fdh4tEaoJqqCl03UN3i8FInUTqgRf8sPUJjCXspF0EZ+UZdP
Lb7t5TvGpBSNG7rjWw65o+kkSiNgAy4RGxO3TTRXEYsX4rBIIf9VePVZh1fMgFlCWvrJTRURoOxH
M2eO6CSVbg8wHj88S6kA/OdU55L9Bo+/OrE8DomXJIxxn3/CkjIS9zZb1xR0jCc3RTVMSPBSXjmh
4W3hb0R29UtnfFMe/jgZHOYYrDbnlPUy/QdTKWyV8FnTRRKv2FprIC01H0DSPkYRp2yFdLZHxORI
b0YyjB87Cv7YSfVl7+kqG6TxYSTyN/dmotLMejlEqYPMgkqzrZ4OACj6q6q11SUCa0Z/J/XtlQyn
DYLCVn+7eVtMHZoXv52SDgH+GXWE6evxqhqrJISuX3IqVccdv9s2uwV+K/QuFbih/cqSPB0ol/3P
zlgELfAxxd9D/2ydm4RgQlorw1BAYf6cdNUhItwUrXdD/E8/devOH3252+v6Le5GxqtPuhldqIfR
uqE/SBx++3/1E/0BcOnRy2jZ9AWemPQwHs+wsOs0jIOjjUaL04a/FnRX1rCHDxdFLounGaEIubVz
hIOpX0qVcwjIofMBOb7KrObVjlwILQ+ScrFdjJ2WtxK7CM88rJiVJ43RxtLqXkzC98XFnpZe2qCP
yC7jRdoEDu8LfTMxvFKYzV02NCr/1gSDacF0N2+FyWjaGzduHyd9DRSu5/fv7gxGrlgGL6NujbuP
schJ6EXbKveVoVzNjKTpn37Amc9dP5if+UQxHOsICx0ekwOZI2M0/fhsyMEGlcHDqmqeoblBbqTG
QTaLzSEmwgIQuWPx8Q42RoDIET3ZYVzRR94V3pfMDkZRJalv1+B5QRrLhkW2NC1Ztrwwvi8zn0uC
Qzh5+mi6ASpDEilG0hwYBin7UVGzFuEc75/PSsl16H+001LyOLyS8xyr0frt9CqItWAzdsLPBuGL
6kdgmK7jD+kGrml4WRcMDnSfss0wYEF6iYT05CWQr23FyhrXImPtOoEfRIxCATEyiuI06WXt/HK0
d8dAfBzDxRkBsluXKzL2cB5qpb9Bt3NlG5i7CiiPAcmdO2azwqF9IH0UI8dKvD4xZZG/VAYFSNLf
15RFsNJG2z+BCjeArJsUI9FWN9ZKGZ3QXZ39UfBHPytOwVn+BMOQXjtaKV1pvByHykFjns6UwxJB
klKf6h9xrdMhZaEmZzyrlK0R9wrByO8N0j9ngE5cP/m3Cqi19Q4dKVlK706W6S/9huuetSdHlOwG
ixn6all4wp8oPvhsaP3Cc33nQRs+VZd3YQ96APVsxjZVKk5+UXLU3hq0cD9PocVY0FyXcwv2obLd
mSCctG++0pDAxCQzFj+MQ7bbNf8Rlohql6ApIdu1ZnLMEOQn/8uOyQsdJAwpmwIIoBzvNZsI7bAE
2pb0nttqwWtKSDCph8tQ/G6bWNin5s0vabc8BTHl0yGWTBm9/Ppzg6nBLeUXh7WCP3yYWlY+RXxs
oe4gqrYZuSrw/Qb8XCrCH2wsir0gT3mTec3PvciS0MRpzVTgtvPgq5Q8SUBURit2DjltQyG71mFC
LR/8P60bZiWAcM3231iEHoIKiJVNlgawr3Qi5ZjiYYrBCfc7M8D7LtMPDQQu2cmeGl3mqxeaZ0bj
mAb4gA+pyRVnRzcJTgv+Hj9qr+RjXz1FnHMTWr3rH6kBYdQKkhbXGGVRkG7HcCXobbKYSDyD0atu
gSm+JXYp+7yT4hYy2JWkezzUFrt3CMyJDlPXQyPZDZ6V3jkgOGkM90rs1NbwAzWW5rgsk+DHBvWG
wvQencdNw9vMrFj8ZQP8TSQ0UbPAZjrvQNWl/a37473k7hn7vzHoH5Ud9ThbykXnmNHsmo79aQdI
UWVqjKNcsXtiPutfVCCaRoqRM5E4NXTJAeQ3uVQS7WoSne87YQ2RpUYR9a/MnYytk83/HF46+ON3
E1yXBQwySTCPGZYyIDkV+ReurUfzFrXhyuY3pHet4ZPMLgnL5/6B+j2n9c799Po8tS6CW5CPQ/Yi
97rQ/95cUAs0KmLWUWIh1LNXzoFot/Ud4UWXSUwkHfTY366e4NA2cytPhHh5WRrk3WVopDJvwZMK
JOYUpGp3euE0qAOyWTa0N/a95XT39KYs7Zap80R4qr0RyhrKp+A8zZDdkc0SYCvZwUuyHNCIN1J5
h0cAaDiwFxCAMaStAh1qIVE1gIE7ED6tDdQeyO6P7m6jbBbp10in1MrHBt0tFezavtLWIVbGUOy3
81Eeg0zrlw7YKtT5T1VgxdwV8se6qvs3prPFzGDNmQn1gIGfzz3Fl/90ozbkWj/JqRnLNtdFXN9S
Bofo4I0JyS4j2YZp6zgyt6NgI150IEgyfMSsAkr38+shpdhcFwS6H620OczucwEhKQ5nF0efxHwz
Qjw1leyJYoYqlcgbgMr7gMal41sls73d1Uqm7j1d6GckYo4wdawEkw4ROItxc+xJzy+RAhvWjPT2
ML2X7ifVJ6RwGioQmTwvhqz3OE1BHYxByf8m3U5axIp1jEBaPogssJtVjgW8swqELsczG40edEWL
VkA+8ELG5wnUCOihBA9QsvKgZ7c7Wt7twPu+jr+YWEHPVOe4PZ/nVL8jbfnymVYr0k9PdmDP9+WO
lmQiphJGXiq8bU+LcAb5hcT9aS8HrFM1X957dkwB9Hd/dYcFOv4Q2r7QiBXJDMywWqyWO+fOxVUg
LEPcR9RCy8H5UvrvaLFSs+dXQLlRLljVYpIsoeJLAkuWpqzG2C2JCTUQncSiTNDgQpENa0HRX8P4
bfZe3yNXxY/NvA56N7NuWoqqtWLRS2u8OTvb2NIueYy6nJ5T5YflU4+YUEYCaJW0LJGSTCw05Dtt
3WbMx19L2iZHvIzJwoPtdb34zQjI7NMPFfMEMs1Ew4LLybQW8sJFV3qWXUVWcaIUX9B8pT70S6XC
6Hb/LUQpHP/FKfjVvZtFUpqjOLHiHWcEpxbbIPbRvgaUhT7oQtjIs1ZiF1Lew1HQxAYMxDer453p
HTyYO3UbSViHAJIZeLkQuL7k8wzgakZg+rdfrDBUqQFIa5EhGU1lgwhC64W856GeblcKTxftndcn
rdQw+JcvVSxD9+zaArL2xv/efrUAYjgM9rk0Dvv12gzi1MBsQJebnT+lvvClcANQAq0Vp2aNKEH0
N5AvoFwkZhNN6HQkXGnrloSCRg+2uL5iTIZgoXeQgOf9J63bHwvg2q87hD+0CqErj5KIYphzhQdW
ju9waWyiJwlCQGm/DQkHwgdvguZalmwF0BuZY+Xv0G0j3I20S0FfpMiCiEYGxvo67R1D/sd5AIL1
KweTdiYRXaeOQLWAigxCeEBBZ67zZ2wUJU3igch/LtcHVgqLenajRWJes5NLb1asztpSzsH5jR2z
we8+9FTGuNCMScA24aaXBWUtGmJRKDadhtavw/Pd2UrWuNwPsYV3lSwwMfgdaf4obzNZdYUAEioq
bl6odThNG8MSL2qV0Aq6iQYl/4A9Sqm77Y+hAfKbiHP3Bad7TCpBeHTHFcj4AJlHbyDZM9qVFze3
3Ye4OHyIR7PsidVPJhDk6qAlruHsPhyyiFID11WuDLTWHNrCZB/HVnLe+cAWHbKOHKDOd94a/Na4
UuJhfJYxoizzlb04TlY8aQwAMffnVKlOoyTT0raLIjt/Nyj6WE8QQq6K1BO6loBIVOWwFuhY3vkW
kEJOBy6uu4NHICF6VbNkg0MaxdBTT7jwSqEE4gja4BbNhzFkkfdB0BezVjjyqJd1Lzk3CCARs/a1
ve99TfBm2xtVhZ+Qdo4vOZ9ar2zOSe/hR+hZJOiXd0UA8tkkHt9fp7YMeO0LJQSyszGV2xSsXcw8
9kFZjmK5JuQkEYUehjmOQTmG692gYnXmBxzdJpUWwbE44akJ9C/GgbIDlYZQSeS1CxOLoK//6jXE
1vHsG95ODZxkuHCroLifSjQhRMppgGsFKE2Ruj1gPePv6Yi7Rfjhj2yEikCXNcaUd0jUR5aMLVA5
lAdF5wzRfdWhgC4z4mwdPclL41ehF6JUqINtJIPQR21Gb7iZwEphI+bKtm8uYAB035A+7v7ZYAkY
Xa/uxy0fdCxNZoMQj+SHsRyKTd0Jm6CL3sIZ5lzNV+2a2ypnXQDRi8YGaBh3GktEpY5YKa2AolAb
NKcgGxg4+95LaCkzgX1sCmN0YP7CeCva3RprtDk4yxDvN1G4RM5CeYIZ6VcG7W3P+fJpEwBBTvNF
WxJ9TZjm0bznyf1frUkuqTjK3Ez+WexNcnfQ25CDTaG/z90gZUiXEMuN5p2B3YzEpFNWbeDYjGsX
/u9N1ZZ1TojT2TQgxKOjrwqE7H2EwjNFGZ0HaxGERFJphxkN9lliG+3JPE7LZA5FS/xmczkCCjUh
zQv4JcUhxVi7DyuS87CYIS5uj6T4+Q05fNwbeSQNRXTRYX8/CDPpAPrzjpFWFq/yLJiKTTRv5FZ9
Mag7lU+GdS25dhlqwmktpeH07qPbZphheC3nFaZKeTfd67LLhESh2UhTCWMOGZ8VASKd7eI1/gOV
K1RZz16xBvAKVLzbELn8u1Y3Za+7M4jGkh/1Dbrhf27A4Cinq8ut74CCxU5XdurB6498BZocWiz4
5h+3O25vvyf0EVREcjEMemWli+I3Ngbh1nMrO7GHQFJ7fW16Klt8DTHC4o5RGbSfeZclvLV8JyHR
HQDSHyLha7c0dUP8LeCqS4fjUB8tWO8Y41Oykn2w5D/XVnn/j3buc9w9kJQiOUO27IflxsK4dJdj
/7ibwMVHpw0t6HtNXwDQ2CbZj9nKpfJAvyXxDLX+7f+UPlvx+cDI2ECH0ecLNWT9jOA2NqTMQcK3
kWgFyBzyz6ubatQ1qIIXV1JqAvvTCcJ1mh9E9Z8Gz+qUWHKWukbcbddDVy0eDSJ+T+4lVX4OD1Aj
PZpuWF4e2SkZD1BrlYMjTyaXQUiPvNpHFZI9vsnG2TPZBJFi4/r5oYaf8IohP5yvSaHMTZfIxHNj
7I0KpSF815yTbHoSzGWqcKwmd7od0d0M74BFGN3SFO6GJ2QLm0Y2i7rbAW+uJr5RlRuNzwjG55Zf
vUQqf0S4s+FKQpqxi3N0WBnBVdvkefkQIlCPPhBc1Iwdxbn380ABRmUOxxeSJBB8rFEeZu4mFHRJ
oMoRJxIXN1zIVjza/tParz/2QrlnVFOWE1weNWzP3C+OYKe6BFgq467mEaWwTWDi2lguVGCK61Nb
a9Gkr8gIFBnyJkPyP67Vcz2LzYUis0QThDj8lNwM6iMHbBqYEbGGfQzKmKeiYscuKFUkpY8cvgNc
uFOaP1k970YUEqhc9laoyH92S/EfQMTJ0oDNMwRRM4jltym5+yWUDtH7hbREXjbl8PCVfNpk3fgm
t3Ez4hhbmHXVMEJuKkTuMU4jHxp6FXFP7HkyndP7pMdVVXWYOs1JwtP+dXmzfUWEZDrNgG/L2NzK
nEVhFizBUd8M1V6UTWdvqORHrDWQaeoDY0/CEepMjCB5niBjNj5kTthzyXUI5ili+xvpoPDsKUN5
M1SgudWBXl+BaQiAKksfbGwokVPL7s6RXGjXoCrxU5VBA8sf6bUrzWm9BIcu+Jz07UEvaBx7Aztv
MTH8K0nZM+iV7qQl8OZMkBuzYFN5vh65MmpQCihMu7EGRrk4F1pgoO9zZlLCmvskoWT3x47oy3tb
cTZfcu+BMhrLWlVkY/9koiUKvfF0OJtlQ0jiZ1Q6TbTcVxv+TgVPMf0UVNLttLN+2oLyE0Ni73f0
rdh4Kv7YVKJSh/UqufEyVjEuyy3TaaDV2I8XmCNhxpAuLyQd8CNwgKxJQCKfyMZuUMJ+jhEYMC8f
3bW2iJgtGf8NpN3nI+SrGCPoWDzEDiW43qpYOFBsq3BT2Gdp9YyHaER0EAMvgP0jEihl4gXw0oAY
8lOiOi6UaTv4ijJkHhtp9f+YF4ijrpb45iYzKtjiOw7BTF4B6zZXdSIw3OMyvrtd//oGzsPv4zqB
rOzv6nGOBkds/FHs/pBw4JfR5gBSeO79YUq9by3kqbrj0a5tHScP9TBexOCDiIdfKGqowItpo67s
cZSH6wG4+MYb/MLA7/OeP0Ugt4DeUDz+dxzF7dbaEtWsSzKbIB3xlenD2dDlNx+rgdBdV8z8iVNd
/LJTjQcgZ3UpmgbSeDeVqugTuzSKR4ukPrgFklD+PBBRK6zT0PJ1LX12w6cD1rorei45hshrQqk0
on3IxyFXKuPnuEmU/ykTOv5r5eLWZ7lmiEaFNcVCjSxxioQQ+zO6MbA2BDJJh3ROZ0cfJS6ZPzbE
5ms0/Kd/7nS15kBSGdS2TO7UL6b7ykeAUsLLaiPI5clMLeMaAe6s5vxtBWYDj5T2zeS6lNq9F7lt
XTpE9OgdM0vdPUVES0K2AHLPbRwSJVb1mR1qPUvM6yWjeuzke8Sbv+x+L7SuEOfHBKIXLltIyA+L
ZtgTM7VC8Vd5qlw3dkEQEqHEN+YYHNE+q8yWqBQCtGhlxV1bdUSEZtcgmDD9OSm4dMTuwAMigvnN
nNbIJynKyFMFz2uy7oxvlt0PgDiExjQ5JjqmyOyOiK9iNn02j9tT7ybCGk5DBUDzAMpL5yfFi2ON
lUYal0FxZFHBpnGgOhT8AcjJ7Dodp897wnacxcKZFeCXld+L5Ora0IVM6GyrW61F6QTP6Uqvd/e6
xWcjhlKTY1lG5yPoB5FBqpWUDN0Ay7C8+NrWj9BEKr+1gLLIKiLwJPfgGZTohqVoT/XvsQmxFjZg
gWfF2qyrs/MzmQLkOG4iFRIH69zprDI4yKrriKWFKjjPyQ7nBFLJDL1obnoym1AG3G2SKVv6qzJq
p5PykYr3sQCOgJP+uURHoEnTM7RQuqs5ioGeJyD1VmLBuMLKRB3Bd5iZXjjnlXK72KIengZN092r
206xwp7+5C9HTwMLmt4EijTEEhDnci0VFpqy/KYUpLa7R3ij43nsoeEDa4KFzOGQdM/xuTBQswmy
k1sMuXSCvQ8nzLncLzaEDi5vBUoD9Jby+Bni3/fd9O90dU0Zi8mvb9vB+ik6E74tWD1z+Z8CpwAN
g2PiBWINXnhG4JBvo6QU+6kEM7avYMrZokmMDAa5GJm0zNdiPP3G6gitF+eAxRB46nIyCqr8IPHV
Xw+y2aXvRXRebuC2zOTPqnfQbyNJA2zzSLviy43SO7FrxbuILq3lHKgfh6ZYGxZd1TZ54QoXH82m
fLxj/1IHe6IRySoxp5Tb/MJmf31Fy6VsP4S/VYMj7+sJjmNuOXOhUVa9jc+YrS9/18h/XMVVTfSL
2WniFaUoWnhDygapgNfeKQIXgptZ8NQeKNUU4GNThgAadSGPBEYIakIF4aH1zyIvqn73K+r4DyhW
5rMIbi/IFgM6Enh+FV6WU7MF2GZa0xBU56LHMV+F5Kt8vB1seDyFVaME6DmZwSWIgRHOOgL9y2Ju
9BhbJre859FK9NKU2C5WBrzv9bF4jsUBY74FsbwCUmsj5S1ARFBWGYv6ONH4jfzWSAPZzm/QvnaP
GGN1fr90/sAC/L0+pX9/KXm8WAstxn8YE73AS2EH+xjsTgsXj/ARjUFzW+okln4HczFvV0k+OHGh
wIQADa2G5qi9mnCFZHUE8fOxrC0pkPPzPmXW+ysv6/GqVK2G8jilFNIt4rSbvEcFtbdfI64StWqc
BKhG+gQwCeJal8w5BV23duiFb1bVRkcvN74j71y2gzVHZFfo+QJnOtv1EMVBOQdKqsC8ytYu5t8O
zHuoPQjCg1p6U0c0nPaX26WFsE952SlvP1ZVCTwY4jg0uaOkdM7keEqSxrWyhkM1MvMf3bwjTsAT
yMhFGiKJnfWNSe0fK+z6O1wiWgn5B7hlYqhBcPHmESCgwwpi5xzD7VTGg0xz6a2WYEzkGUJ4yXQc
onARvMkAAMVKc/tY4nLx3ARNgO/66k5SL/8cjUBB3glgs1TxXGXtiRfYYshuRziSnV/thDfdoaiL
BflNt2zGsB3ijbCrSqMqbD2Vhni/d8X9/XpFPUwFBrqI/R4YDMmSgI9CvckhTD8Xi8/GSK6fk6eO
5FLFRLlrCuWm5ALXmbsKI+1Fo9khkhK7IkFRHlLhtXBlVq1XtBZ+wnVM5RiocxtCDaV95KhNkE6J
mnW2gngdCiSr14VY72p1S7MwkFmpVAS7VYtYxhK6+fnK14byzjdRM+CJ20KEep9ZZ/ughO7NXaeZ
pZ1VrkWKD4juPTqf0/6MGySdi8i6IqTLAvExjawBlof9cQK7Fxr5EsDBIatEgto0nc9ogc9MiM37
mo7B0KlIDXXz8nI0BHqqaDYa/J4ucb5TAsZolM37F+2rFHA9o1uiWTdsokmDlNULSbNXgYAHi59x
hRM+RWmAhmqHjO1KGemiECNDW5iO30N4lxcwj2YokfgxKQV+r9G9NBS6IYzCKq5j5Sa5MvcXDCs9
OaJUdRz0kLnsZWJ7O38pOVoQVmG/sbfy4+YiO7jHkYZPgecD2M1iA5oowZ80dKv8KTOJ2y0KoJJb
T5Bo0Pmf2R2kM58t5RBuhZIJMazcGwUhGNNq8rUzAFr0ZFpURnoeCW9wYoCXYyNXPrbkCVj4SG5d
AApG21bxjG5GcD8xtGCzQQGcEWE5+KJMZGyJTsi3tj/k/sYmfYXPycwUWiPKbG8I24hHyqNVgNFX
IjULh/h1kDECuB0pdp2Lnsx0bmGdgaCPRASin1P+vrO1TeufvbHgD8YdCULWwsZpDupxJt6LQg/Y
M1AO4a3b+h3rn6QWFV5QxfeUtG4CMPGF7iXePOV2ZdCxs79+5zBUIT9xkdC7t+qdpVROC68WeF1A
9QWgIwzy/cdWAp82humHe8XjENgZPeDj/NcpJwI91LVWqqOfLMfpknKFti3t+uqvfjmxg9LE1IZZ
iw4bbmfZwCf8ph2Mg+8RSxhWdl2XxMc23HRvew4NEJEjxMLVbG50NLrn2ReAC8rgyRX8t7hIUmVv
5j/Qw+3Q+eESftFNPbacvjIpSE4FJh/7kqfrEelYNsNxmMtye90ndRKoTQetk7jeQx+DuXUURpFq
gPwfTwmQMNd+Zmr4SOB+QSuqFx1bc8xSX8c7Fz4lENwfmH5XJlzo+T+XMGBgYALA+nZjXG00nxqx
9feUSbGOoId5Z7fzrEbh3keUKaxevFze5yD6oFK/7oSUKZSHik34D0wZl3NMH98kuAHxB/9/UhKg
7TXTiU/JIhOOYyvLbS7Zl3y1yq6hNVvQ5D87UMzVwn11T8SIdQ3VWba/jExESk4PKK91Uqc6g9GN
EnzD4hvG2Vtlqz+Rd9Ia4s6HC97OtFDaCxI/zcpxb4duOVLTUJTCSYTjf06sfaeNo6ZQCNGXy+db
IdllYHiudB12Lklc7dIV1uv8yQT7RUB03s76uLyjkVMeLtx0UPd1ZJHweOJ2RJIbQ7Z+JgcSZmA8
ZgV9kTg5z8JihMTWjTKKykkxKHQ/dwXViS5OOX4Ywfz6lgwmBB3y7yr5F+sTGdmo0t3KlWOI2tZf
hLQsr8ePnRjISqqf3bE7ZQMLPzfOPxQrFjOkxCKRgUZrikuCggJyrAmDGbzDbjz5cgkli6ud/lWY
AcVV4Kc5Z/wwABWdXpn0Lv4tscDkaXvhXZCtYRXJdtYZM3o4d+isHi4D1l0S/GXATpp02FZyjxKj
xNS9v5rM/m8hiSVhnJHl7tLbG4jg7kgZ9ETOCmtyPlf6B7oBTTKYSPFx3j+MqcQgvJkqfuNAhiES
DaK1CMRJJ82JmgBLxxOFriAwafnb+HOAGokuN+omgqxhfvgRCIzjHWcVv6RXzSMB6biSbKMi6tj8
23uKHpH4O6Fi7mD+k8Gd+o+uVQxjrmugpINwWHoKWxResZBbnKVDsUjIm70pmeMt2U+5WEhWsl7p
CNfbdFWJSP+DbZqFRR45a6F/NknDDJB9qZ1CqNhdqIej0uJJbnP8aiZ9ic5enMpf2AZDDzKjAMWG
01gNTbL9aHzR23intzPowAdzYuu5Z1gyEidqV7iP220Bgky/tFTaalaVMH1tlUGsH0CYAKmccfwT
qj/QeDyyP2IlgUqkZuDLg7UtR/s9ZhOvJGHSMawmrBvrpi7M55dwg2ska8vKUn7SyUU/u79HVDA3
YoJh6XmL7sD1WTOyRTVt/wNd/SUUMS6cjcnJtRxOS77tgAhf/PH9iChLYAA6/07ji5JvCqSpEwN0
dJdpH0pVsrsBVYyBxnXj95K+KSfAq57dERytMWg9vCcycDLFIUJKnsEkEWtj7/ZQXJnvyyQFSoIR
tAwe8RYGe32s5twWPjpcXfXRzuc12+7FEsIPllwCiDFokqy+X7jSoonx3SNIHD+mtei0p6Sk5lHw
01Tw3HhL+Oz/82UrsgZw7QnmRFZD4clTuJ7zFubt+6kVLOzzZo7SJfjNBSWLBwEs3WHdyMVaheEG
VtylCo2k+JX7m1eFAYCQ+PtAQ0w6Gd5NBK8O9eURNHIaS7NsS6Z8uzHhsup6X5WUmapqVCO4zybG
n7BcAZyU5qPi1PIcxJObhJsYB+otMfwgqpuMyDWyeON6vqEjZmolrc4LFAS1duAWIaFUwfhuUEB5
kv1u4blfpzfmTevIKuPwz8kda41D1jfyua2oAzG2dUBRNkot4QpwLZcJ8ukl7t1W8WahZjLif/l3
xpZIcKuBbe9Pw9QxUFtzbemXjvaLg90anfAspHnLQtGLSYLt5aW9D2yLH8n5xGBiMzSUYYIDm1n7
XfRKv78yL7kvU4CzpHjmYXszz4/IWHMAB9x4DsjfRstdCybuCaJZ2G3rWUdtDmuLv0SwcG6a4Rrv
73ccKphMmvJjkDXdrinFX0oFvwcicn5TsWMdbF7BE/VjBXHEVX1ca+kZzpshCNcD3kv+WuXcHiAq
/4C5OuQ3IV/vCIGrAC6rkQa1kQSgZpasDeQNuW3zK/pNgMx+0/RrKEWxsjqM7kPOY8kNCX3YQT3G
Z4cYmBN0qPRxqAbuYIVrYyJLTwowYHqdKp9lGDGlhdoap+BruOqeQ9EVOtgL9K0BfvKD9SypDG4N
V1ywAqQ6LePX/ghU2tqI/UXMmT8eOfvLLcnVp39PoMvJl6DkMqOUmwSOITJf7WFIicS4TnP2luSe
y2Sr+C42zPvkOvA6QSdMlrYkamFgfCXcFiy67fDhbzrPPKeAXOtgAit1LmcIHhphg/DPMWn6Jz7E
h3lNcFOKE8K+uMiZq2VFsE3ZsCxW6qeHnQ5qF99YfNtL4fiaxSDz7D2MADUVixqpVYKP9gM2IUdC
jugfJWYkuzoqWWcbGf8MXl5kadHW6hhtFcfkUO4fmEF54HLaVGTT5jO3e3FKIPZROFQKf6yslgYC
LBfruyrBfu21lVAwtihq13DXA/YaVhJdZ7vkBj/FZeS25YD/oTqiQsQ6yqfGuffyoeE5lNBgsJAI
1Vh258kFi5UfC1KrFbZCF/CCFq5A20KI/HWf+0Utd5dC++8GumAp/80eBRwdkerTPlxKx8ohY/w8
miOQnlml+tODSsiE/FX4QHeRwJPAc4aHKLdDR9xlk3Hn2vzO9u+VlKEZmpmqQ1FBC9zpO2nE0lKq
jezR9pvBfnGJ7YEDr3TgvuV//mn/ihaoFsGeuBi9sq8oko66uT86dsVe+yBGIfXUWQl1j3o3HVFv
CvnRFHaPBuQxk+o/PIvgvsCCuQm+LdxfoZe1y8i7yJCpjaFnBTUlI7ioAznV/43/zYBKR58iU2ip
NkqYy/lMcSvab3SMSgX5YDSmNeWKeCKCEIlWrkt8AmmiFOyq/b/kbh6pPDi73n2d5UY7+hCmCut8
g3kSgHN9uyq4IYGwjkpmJuV6KvBGxbQ7LW5a0MFrgWNeDON6ItejJqRc4stAbnFgzsQbGqAzk/9s
L92uKHnhHUxfRFYxeAPA7PVkNeHbzdJGEQ2OUlFGG+bLNWJaGe1RXS9gs2tlALNMJw17TfSeV9EI
WYzZ2swZAzic1li66ZRMuDK+FxZy3NFDK0+zP4k10pQgiynz2hcC6k7VGBI82i9xU5jb2Qi1+HO0
NqredRwgRjvpDhc0yVNNKv/SW2ZhIl8eC8A6/0aM2AzalZSGHngMUI0aW94m0a5wnTn7mCxmdSTU
NyCcDLqsiBIqkshOYy8wcTsJogOepBxCW5wQ79t+EiAkrqBE14VYnx5qO9tRczwgST4VZhkQToft
wAFIT7N/RcEyZ1tVokZmR0dyvg2/EZarYcuGO7bOhiFjb+317ACuLPHAmisMkE5RenDkYRpRLD1b
DeHK0GumySOjKqNyLTCZZj4Orvxqqc8gBIfjM6uW456mBZMLQCdMayjc0zGUQzk4KyxdXFl0TsWX
CPNh7ykssJ4eOQDRUMC0JMPSgnDc/+BFd+86MSzHNQSpENV6jNA/79GexVRbcs1nz5iHRTfc2UsR
Jx5tCgWJIGsuRWyNIEhOUF/Q2LzGiw+nz/uXDDo5ZarWSgCd5xqci84Sp9VSYKjTofpR3jgzMdRI
l1PEbLq8nAUv0/10wvCE3fV2VmcWX/wzXA6McrNu1vlnAY11dTgxjThE7pV13LQJQkmqhGsRI/r9
vgU9mbYC8b6yV0velamBiOEUIdY4i29PRIBThQuLLHOJT4nLAgYe4UjXqAElksgMjw546TIzFBlV
dGBR46IMnTLDyCP3GO+Ny86FCRTD2eVwIKmGEqbTMXOXpnPcilfGs6s4eLH4Aac12VF8tCRVQl4w
E5Gt1chFfxyhASYGXXQTS6hAT90VKNKHyEsSGLN5YtlGOYWR1xpNQgl0LzJt7xkZDxAub6dD1ECn
xju0+Yp1UG8kFxDv3ufsdNeOUNMM/GYBsx40wrQvdcEl1HaANKNAqh9RuEMxUxvnxx/uRETj5gVr
KdvywRNf4Jyd9BcdEyP3Omn9oQ/bp98brIaC4xFRR20Z8uSgdjSoruAEtLcN4byeCXac3bzVvvO1
J8A5cK6SCmWTyiTCvwEZ/oft5acUdvJwjrmzMPnan+4eX1py8J/6iqa0p9IwYq5M/mwAg5LNIpVV
HJZQ27FuO+zJ4Pc5JxRYopKzowU39ST2COP/YndlyLivx2lrTFCxMZaTcgnjz1N3d97jOzZJiiFQ
t++KFZeJuFZso9u29GZw/oGXjJu0L0V9fXxuVp546al18cQpSjPaw17g0q8ZfF4wd56Kq9qU5EpZ
tPvtOvB+fJRgHYBmP66dY/hq7d+8MyEiCMf5J1b5B3C0/LRtNg9c+0vsjZvXbuFeEv4awnuVqviG
eQnDZYhBz41bVjw8rJ4o9FJlH5/Jeq3MIDHFfuSnc0XRyyKGQ2ngATUSQHLDbw7x7zWG8TndkQS/
ZxTEWzXRVaGIC8QoeF1B2khEDfkhPLfo2ZGRMm1XjIDSPKCWud3v9cGRZsVworCoUPGq9dBI6gq1
LVIv7j2DF1WUMj7kYOD8kuNlSwregVOwA4hyt9IehkKs35XH576Et0Ni2ZYCJntqLTZLtmcJa9sT
u3L5URw2W0Fbs2nvK4YXW2vj3Tg1CCVzofIQnrE6hhc+Dt2PqDZg66/oS3qG9SJLiD62o81yTUKb
VDi6RzFG90GNUFOmxV43OCzA1iUfuQiJ4csglMsDs45e3j4uUdx7fN+CRskCIWMQ4hXyy5QJrTAl
KwFupB+w2JoTNOGATkz+ONFFDtCGKiVCfmFNLvWUtYP7SkgZwGriqPojZZTXegRN7g25tqFR828w
uCB0jwwQNVBFg2Z5ZLFbgVmba3dZv1HsWUr1k8o6EL24ux3Nmd9M9eB3vlYexL+ToO2bVUMwuoDd
r23bxIdZUeBXouMxpTjp3GppcuGGwvzkNDHN7G9mG8ylS+vMf8PWDrV0fomimnZQxhnn5UQXejtZ
GgTZtC6soYjBfzSxpEpaP9deTkOah3wEpP/6b/14uJpxoDr9KHegMvOsGy71EBghPlOiT0Qk9qQl
pt8E7mqNfqFGwzA8cZdAPfJur9xbh+2H8veDqfUjkNDryHeILqRhAoBfe8kkX+jrPOsfY4ENpt3G
GS6chhO/T+RWdizadyazq3HcIHl8IS2eDqdziUpgBAzftFQvQVuVVuj3+JLSLKN3kER0HVg6/P0v
t7V1hiN9t48xPm/uIUnCf322GETvqOY4WQzpULsvDTE9bvWdDTPTUA0TYN+izeQPlrcdq+Ws9yPK
MutNMNZfFoYuJCVnhPYZerF8q6niv+2XWV/j2gh/Owj+ru/xGtP1P8QOxCJ+Af7BairKT/Ux1IM4
ii63HH6GQynbyazCn/FGG+J7ND0OiJVqoUwlK7R/xIEsdWe7HWSF73mfq6jxwwWJ6Kh26mmu8Fmh
9m3E/egsgcpWsaVdesh+idT8+skmzHyqryY9NYg+ZoH0gqMhUMmeLmTaJLOo6w5myeTNCOD+N4nd
yuqCdRaxNUEAaUdokboeW1gG+QKho/lYokl9B1uGdFM9EX2FKo81J2vKqruLfAsDhCcxbCdlXoyq
0MbzaQfk2+d41HlraBCL8KhyVOpVKDN3emz0CBfZVpFm8ogRBovgjR/VUlGrbpBl9ENvrCWl6RlT
Uj77Q3mvFBSnpEcFH1JSqM5li6TGoMIUdDC4k8Fi1GvW7ZtSqvtMsHPfySDe5pZIB4O0vfdXPlWG
lkL9bcJWmL4R+wZSNBkWUgM5BMUWB1wUD8z5IECYV9DM4IrwwNFkz186qq1VxZxGWdhJY6Hf7zf3
3gdu04JyvwtVWhOqdDhNC/UT1Yg5WuZH5jKyj6JGAEv6ve82EK+6HO2EtOr5x98tU3ef8Ph0iGUa
9VAZHMt1SdlGVbfwqCIcHseJO1DCh3oCVzGDPbZlKqwUoqqsRjPs9jORN0sioIXoyDVUA4KjqxtK
f1Tkshrvx5KnKa/4rCckvRoOkKY1Th1chtRabGYwCEJT/7GUOAFBma76AITJAzViHS5vHKLJsNGT
DuYlqp8WmrNpNtdC++2FImV7Lw1B43h2dc4gOzbzpH6OT0HHseD9pFFR7fY8bQ48Shei1MEnb05f
nXsuWQGh2lkU6LhQ7D8F66ifDQqLBmG8tjDw/69TfdBQHO8OI4f956zoKpQ4yoQYbhkB86sZw6Xo
oCsGREM80aJ87VZ2xb6Dd2Xd4bOj23421tbkLHziPeYXWmyVzwvFOe/u6cn+PfJL/T1LzXEJ/zSl
10nBUJoQvPWoz1I6FRs8QUwvXSkd9tgyD2YxC9WcvZLIlAJZmn7hFIhVNLx8kV10hTMPlU1ukiSw
AhWuUlj3fDVoCwaXg9VmHya6t0AZDbls22QdUmdptYjebv8MN3ESteq950t4yFTlYk5tdMlctYIP
YWu7naC7Zn75Aky+Xf2Fk/ZGiGGL7eIrmdzIwzKZP1YAckOv5td1+1L6JY3y5sMebhmLzraM54dm
PxvdVuzdCoag6nXcpRNSx2bu2ZtG5VWrsrovfz/Wx7q/pyw8jeWsNV5W5P7iT3HoX1TxaHknEEIX
pJ91qVG4SzeCC1LpgKziiEi4PHOLnGxoryHytMybRj2Vcrn/eyRnd3XJEoOJycT60rmpmI7yXWRS
LqpU6cdpIE09QqUx7gFF/vYRLTCvS1Rwr3QNkl8N9XmCFIKf7hMjN33xjSUF0IZNcPVQ+03+bHcR
DuAk0VrRLIkWEQLZLfRUjbM0DaLJk4EbPOhvfjKK2dyYTgPoO9rJ+Wjj8MR4EBzDzHrjtrZVXRr2
IqaW5WrXNYfzltRL4OtJDZBNrFhXEI8qq4bGIhy99LZxsmTune/yXjtzsJmWAYBD2s5m90FYA1yx
GLTxC/YQlXoG3Gf7WGmwjMVHOqovieSYFBiX/mcKCffPJWoFSxjXBFLgBoDIGOjCdjeQbQeJZOlJ
9w0lOqZcY89qf8hOn+wljBooqc4A9MW+a8Cdndp5Tt4MguTgLGhYsVZZtwwcwhFkUYcEIaiYQB8k
/99yLVKp6dIQq2z4Y2YDfl474pppAo71apZDbx1wFjy2K0i2RjFUtEmxxQ2HC1M9NuJ4Ppeyu/Cv
y87/MYl6IAwkYguAzOT76gakn0KqnFEK0x2JFglKOeBQuFwRpLVkxW7pQ8V9nCoRPkyAgdtc+I35
huR4aznyvzVVhtu2IxvbvI+8Yb7BHqxCcyN1Xf7Dd6e9x6vH9wZ3E39Fe/p9rfKSdDdZ68PqrN8B
B7SyGc6C5Oc5WQLjBdGFeMin/qfVZ87Gcz1metuOoSqiAxFAZR1b0rvuz9KRlxe8Vc/q3+uFR5kB
22+wd7i5BPXeDax74y4lTX4/+5csoKZRv/4q5OFpi7D+llZYklhlHZ6Ic2Jxe7iiHikeCjoOxXKQ
CIVIC3h0YSpNoXfSgQ8RnRs08CmiTznsRLm3oNDEXPYfeh5AfRsfEtx55VRYXSCGZ90UmuzdB7Yg
GaODAVVB5Z68lXz5oOOo7+q05ZhqZSUdRIET/tYh5nO0rwBGvWL5ZexRezUSSOcV4dHKAbt1t0TJ
fzHgH5F/rSThNFGZ/L+NmC+LBQqMxyH5dFpQlrrDedyOM62wNlF2Q+AiI8I70+4CYCQMTtuYFkaU
nU7sZP0C+btLigc9w2h/Oh7Gz/817eo5f+oRqJEhvqE+Epgd3QcgGwITubERb4Ge3vkI6bU0gzyi
pH4WztTm8shbFN0DxkBDz9pEczGrSsoPh6WPtzut4FBBXdymeZi7HRhDoHP9ZB859gMCVJNCrxkI
liF2NNoyhu/vlJpOOUYhlsz96Kv7witTkgWRYd9mDgYjHLdrGBZLulIv9QDLgTiCUM2vo4LlL6ss
2YFXz3iVUDzXEjChTRtmhJmpa6lFkKmlSHgwxrjD6dfB7RYL5QcYOG2mez1mhQEy9bRE14TZjR3n
bep6d56V9463AHwHE7TqVvA2aSaP124NiVec7HwaHjEq0dsKBxRT/VGVFVkGM3MHeIff61vw9AMv
vZCj4CTXh+pSCvkctAviP8Z+/YEjcL9yQt3nI7TPc3zApyaR3EUkjMW02Hf1OaXwv1ola1Kae2tT
XmuXAnfuqqQNytg+VKfSNcULlAOm12LCFvs6ziggh/oD1b3IrIhn4NpIiLM7tEzRmOy2EzZ4u1v2
Ykyxba2Dzlpw6pxmzXO09jz6pZ7OoBmM5Zqnf8t/lfNYQUUAwRwXdi/tRLdy+3SjXdj9gcFaFYiF
pts4zgv1nI3LzDe26zBccrNobf/Rmz7fjC2iwX8Gl0hyBx+Z/FmLwNDLBsKVdD8TfGogqpBuQ+na
Jcy+2AHqHU+czqisA6Q7JY7oukZP70HXPLnL5JR2AAWZxLG52OuvJp+FBCgKXmuaZHsO+fWQhaQD
UqKetqXbbnA4rgXMzXwwQess+LIb5zT9b8ZOSLKQeEq0tPrzsZMJ7g1ZdhyCRfPkgcxkgxLr5fwb
Fd5prXqY+JYJw4Qb+JzGysd/NUKSkwh4zgbXot2ttYla2BvnfUBfEbTHWkyg4RJDsg6hnRxJ6X1B
jGK5OlfAkmRAjYLPxf7irlB5+nrtZdCpa2ZWU/jcXpjpgx+dE6MGzACzl+aN1WL0BBv+Ts49nimy
OsqPCBGvRRVLothFtawD0YAtTV5OxS5FG+6lcZa9Ky8jMgEQNCRFQUwu/8TsVNq0s30YL5bViVHN
NIab/7aQJKpV6n+xi+pScQPf9XgyHCN3JzanZ0+XM0pbQCPprPHHY3/gyBp6YHiRhVJuMnLJqN+J
qm4UbDNjG7MMXVDNaqXQuTwyYkWmagg7jOfbQiRygUqRZKfN2BJQNtrg45GaSk/PWllQSw62iVCz
TvYZ6cIh1gu7zPtlu/NKPFAcahgUAS0R/8NNLxasTA0dQAepr1Xp0kTKYeDeSsuByXYCqYmkyc/9
iZ/ULpG+dm7NqKDViZAqk4XFO8rSSk61+dgHPJNrZAJz0jS4+wmUY2wh0PRkBzgOTzoEjYQdPhHF
jz30LzRIv9b9aJ+YBaV/jT388HMXevG//2PTfP0Gw2+m/NJCjd31TY0Ek51tZ4tc9RIIBGMCdr4m
1UyIzaZzl8F+KQAnFXW9vySXNT04AR3PonvQYyiF58ApDuglLYIN7EQYQ/ta5DNatYHDljp29Ge3
1pX+SvlKmPZVVzWA95EblhjX30Sk/CgIXsZ5LvrB2t4U2t0bUkHUxIsm5r+5x59Fl9DSQSzoU00F
IAAafYFyh3sDr7zhJhN9Dv8/a0HS4HQjcF4M64r4wPQSvZH2da9t2HNq+GbJ7HG++8nYhmZkbacS
NmqMtEvy5+l4sDnzn7+MrTJnottjGcmnSOafgtaiJVehG/l3cUPnqdDHBPUsEexzH41TC2QYmivg
EGyTj1kAjsodILfTKSADquHwaLO3nhrVzYctAdh8urPdpaDO1IwyXREGTbKdcP2Cb2wfz7M9Blfc
BFINcx1X9xjrTA3a78Vq5ukRFW9oyUxqY0Osuss0VekBCeWUAE239luJh1V5POM60opscWXTcqr6
BPs+XGRKAKadTAX/rtxYKsTMbosSa5HswxPZ0pKE7Z0hmNL9ZsWo0KqviCqXG784+mkcJZoW1zXH
0PVXrEQVrR9a/A9LEay3oyEPVj/9D78XvJ53tHVsES6kEvT5N1MvF30+DZcvbyNWHrOoCgOm0TRH
A12LBIsBW2MINk3X+kTvGfx+hYuWPjJGZOD5NOeTM7+2Ts6VrQWWpOZxAwraixXM2rv8HYl/WHnT
hCczKdM+OnKk98NGF+w5CrCXF+pedfnzFX59JhEVlc/BZ+RCNr6nwXQRqd4THhyMG8BXJ6tS+JBQ
27WN59IK6cO4D1CL+y8dFaH+Gtk+vOFC9uQLV/cyvDC2dSbaTM6umqhoWnfJajo7zmWjUHhAWeT3
0nN7z8pAfJ6k2S305RSXA9SCZgVGOpfS/ehf1YevaZDm8j2Q6PjF6ew1MVU10JK6Mpaf8OhVNn8b
/Ute7Azup2e3pmaZ+IGSjgOTIOyhJQ1Q+wAhdOaOA88k7YZvXgvp0enbcn6HFe1tj2a6+KNp+rKc
j0+nQy8vuwkwS89FKQLGlokdi8z0i8l2GByhZRKNETXHnLAEF7GR+nQWOtIgABH88sLumrHQvfmS
oBpUD8t9MsMFFmAGBZbE5QOPKu3GsoPx223u4dmAEVjvGDLVmLkimFofbyfLFrfEoRxbF731T1bP
zfioWBZmg8QA5VDGSrljpKEhR2rVZCBs6rP0Jw8ZEE2ZivsFM/kddVEblEyQwPdwnREujvQDXnw3
7XNVBS+WkbuB36EWa1g9Dq6cM5fb5oMDbBWNVTZ1kbkuw9AR1yKuWOEzOszwDsmdAmWrYmg2BrGK
WTegj2Esb5TzWHISbKb7FJHLxwf9Sr94M7TMqhM+9VDtp0hkAjrmwKaTroqQm3+zTJjSReAsuJYh
SSTq+twge3Yk6iYRIMHJBX1RYErtlyqeyI5OH3Rwh2RTdMaa5mwz+bECw60Wy0KssJsGQlwerp0s
9Cn7I2Fqtxd0On+Q8qZj3sDJRewKgdKQC/IH5lbwOT3DefzfuGJLVwgjjbZE/Ad8ZsqzXwZHq4fl
WD5hnUv5alWa5X1WyatpxCkjH03F7mzSAUxrJnGkr6Dv69AaOqSB6TiPlDSLSeB1yPAXYCQO0xhH
EyhJD/j81O8Ex/CElm8+kXmchxmu4W3pVzSb/LwZWAXpVUBYGnk68e1Z6CnwENvcqjwkd7z84bUP
YpswCNEQAVEzAtK0C1fxJiVgSaJwws6wLMgGJTpzp9qWCI/QO25kXvOmNwPxa/LYj5OZ4E51dPnv
lPrDgvp3mQwdTFDVM2SYeodz4F+PIcVbOfJxuUnsKItvgzJJCpNnLZPuGS+uPTDwQ1uZY1+nE9fM
ThzFew2fJR86JwiUwUhc937znR9MtWqr5q02cqyKO4aYv+g4A5BD5ocOOQTk3ws3hDEC7JT2ZDGM
bgARfY/JftyRSN0LOmPINUv4WwtNZEadBSaap6Z57h8fUA3kT7k5LQjQNbM2QEk+xZdj+HLFTUhv
awjKHbLzDrY1siyvYqAxZWn/ft+cfPF6n2j21pbD0DaWxJhFiZlwA2nviTy2044KLbOOmB4om1/8
R5M7h2/smpg1BSnC/5UbQSzu5Vz9ApgiBKpPDvxvUhRjwk+KZWZ+FTFzPifEfa+VrhikSPy3Hu1K
Q1HnYgFH7sACsNGseGBp05LW/9yqRVp+iGM/8KnDHjjYCHmKJoW1LaWAnvd86tRxqs5lPGNEz63T
Hohv6gbnGrvJUB3zlaNFKg53ujMXEWIugcjfwLIZqf6Yo1fz1WTzzR/0kBFkYmj+HL4OG1A6ezRs
ao/SQ40SAAbbma+uI01dHHXHY2vuB5jd4xXqkJ4gh3mn0C8ZxWKPuXZPj3+EHI+b8GlTAH496AEb
qK0i4nuAdI5DfCJvwU5ZV/hEWiTwx3xbmJVTnKZqrQ6ocWVvpTMCXvw8Peh2pAmBc3g2mNuq0m1C
nkivQA6zEMYyH9vE+IHSZG3VJKupaDxX3kTM7ChIAP3XzcUEQtiKQhQCH3AMf2ya7iTHfNI9KgAX
yf5W/tZCCiAd0fMF+wCWxeopWuT1T2cpNBTJwzLk7Rwn+BhSeqaJXgW4e4FiC1giU8NQjYlUFqHR
9L0SguDs9hKCOcIwMN57UZjajAsFQrKs9JYKeHKY4ZYxGcZTKIma3xUiVc8BK2FciYBQ36r4nFlc
5/qgMUd/nHynwWMn0/M0bHLAGyfi76WdvSQY5qGa84mFHutraXkzw4p1DqJF6A8fSq2hqPZk+YUf
RMiHt0qdXdDux6vuIvwywBanWoDY42OItK4Xmzlfw/kLOTyPC0RCTLqvDrsbmPd6LO3iQye0C3yE
/fgew8YmWDT4OI/NEAcgtpsZEGm6oNdZSqj3AHI0rdaUqzms0QGTc845X10xSwNLk6BIhOdRV3lO
jBwBLa+8SEBfhdloA6szTfdhXox8QgkgAsB6XEznlN8B5ZIAZrtE8NqnQn+OoTMjXIn8+Rb5kkqx
nuhljk4bkW5quDZBweSSDaWfDZIKExDRS0UwTnt1/kq1tf05ZdSllQFOdqBhrWwuWRKyRwkmUz0I
m2Mq6e2PT7twyM4izjmA0YYBe0HTlFw7FatAPSZTUcbKU1TnFv8JpQwra4kK5n/pgUlYt6rk5IVg
HuMDcEKVNF70pudSX5y4zB9wUrpshwcSrkJnd0Y1QyGJgE9wfhOuj5F02yR9EOE7mpJlGYr4yosN
5qDF9dDB5M49XSwGDUFQPGIbemiEFCEKiyPxiq7BrM0mQ0UdYCpysUmCBTnwLfd/mHHGptQOpFZP
M6gauqB3R8C1rr6LbHGYikc/KJt6d+NoPgJ3+FYjVhVFQ3sPVvvF5mSUwulmpVx7e+5mw5nfXPLg
QYRXctk458my+c2EtceVxw5dDw6IWH09ZczxALiPVxgfINJUYC9iVV/jYvuMbaeq9/f0mYZ03kiL
y0h8z5EwPcRtmBrPpVCLfYwnUy0Wxw5o+QdJ1rhlr935fPV+rznFv4KCrF/qoSTbLc2C4Sbpna/x
iRUAFZw8sOvkmi242h2heBK8GBQL8mYQNsnrYLsVZb/aVzbnMPuIFTSD1r8xmc9fmb2fI6HKWiuR
va7w9Kb4/ukJwpqZc3kk1X9Zbc7+ESDR+ZdUxPlK9cWWJtHx3DoE1WqEGw56USQdutvLqybco+lz
h89q/XYwKqqV1SPHLfsEZ3wGtsKTj90JnfnFwmoZToSBmBfrCRIV/Mi4S/qaZukitYa6XjUJ6VUJ
J51DmizSFFZr/PFrbFwqCtvIHBiXaVg0OtxhSbdEKLHBtH8b30P8huXhFkzQh/DAGg3twbbE7UJO
wgt30wMfIjvZdpwnqQMLGpWiGt0aqtgEfjJ9C+PbGl3NXpYfQu68Rlg8INDunI+60nNDLnz53T9S
g1verY1GW4rNyGpPmXxTj+/o3JX+7igWzZLy44QkKBDxcjT2Lx3Yr1kUE7r6cH5F0OeJhcN7F18x
PAbZX9RWzpNtlReMydnBrI2KRZSpcWmnCCNDWxyEvMu/BugyUflzo02rbWX7Mbn39P9AScBD05zA
6S+gDqjsRg/X/rdWxtT4qlDuvjeE7JWHKZPGVPgz9eeBLcHlRxBLz2o6SrESCEHErfpNbLyLTDVk
hTAgRbHn4dmn7IYjMRIXxfr8Lp04Jx8bb96zE0nyqvAG5pRupT/Jt9lArw0YSjwZiwdk6OnYPLk4
jar1+wqugriWV9jo7eJTkenzaWU0mh87dCTOvZXqFnh7QjMPB+jHcBKSCHx9EmFJM0ZpnuTLckPX
UEONUxrzC4tCAYPNtrVMidvv9GsmaNXa2eNk9f7LjWK7mlJzllaCkGD2Js67I4oavLiG19tESENF
Agryn+oDcIRoOgwfbj37ZLJscfZ/Vkj6MSZlTkfUKwd6XENT6OGgMQbX6hdnyRybSKe/lhsFFi1X
b4ebuA10CC66O4i1HTxWu+aiNrwnAOiXjWtzpXBmkGBteTJFSPEmk/ymW3etnlDyO0mW3r7GEB3h
GXRWZYJgjVb4waeYKYDOKxcpNMdC9RsWMa2fdr7cXyGZFBNEfgk0e0JuZ6Qsto9xdMezRPTWFN+V
Iupu9JybqVivlhWmbmA3LjDdigAeyVmS+Osxl3DGixvCIHcrAJaUc+9dAn8JxTkkxQSioPoGEcYE
443G1rZAJMmYVuQh81vU//NzpQoAuhg37edU7UvArv/vBuOpl/YT2QpVvFXf+0ZAesbrt1Fy4BDA
Vw4QN/OlMPkxZHULN/uRg4ysYEZz84BPLauq4CsLm/oJxWhdKxTspMPhEf9N1rGKRBQbQp8o0Tyx
7VW+SQU8O04afj9uJuEyTwt8CmOGx9/LDlDXXGkdKdgH0S3GcURqFJf7Gq/npcv+OccTdcrW2RJT
8jznhkqsm56kN6L5IL6OCJYByybzn+Niys1RMTwF6UWBA695moWgwL9hTjOKbTynyHaWNizghnBI
Gbxkpw70l1TQIY7nWzsy9DI8rsUgSOEmvPUWuvUPMYQtkJlp+j8jsfD/d/XD+N3MccuZ32RX3dlb
bK6oeptY0o8E4VRNCSn4gDIlGcr1jP8RbRMQW4P3H1yHxttNDFY2kc4zueuhyGH/+C/BX8M7ZbWr
9a1h59uFEvtP2p5qetDS14D8x4oaYCh5PJpfxrAY33p3QjsMpMB0DDud11FjF6NpcJoRJs5EFUbG
P3obW45ry1wKQdqFzXcpfuzzg2qQMlh0zSZzIfBFR4iIrHM+h4uGknnhtx15hiDwQPV6vS4KBKA/
haCVNs030e8CAPTIi1Som/5Q5vj6dtVqOzx891dOMUC321YBxe0xC+qjgv7tnJC3e1VWrVEeNbwe
eVEWPfId4e+6zLfSzvEzGmb18ZAwCacRyjy1NC6NSl/Pn855xxyOVoVAP+nkPGj+xJLIcUk+25/G
l4Ptm2wP9sU7hLspxeEldB8ssRM2dg+1Qb+dxYcxdPD/07e9I6grmdAYnZjCQ0HwT+8FDcKFO2or
aFa5NrmvGsU3UjGVed6r+Rlb48FkiZBKU9O/ffSgnKSK25hRSOFvwCbUhfd2w5pEE1/rxP+hhZB7
pAIqH63dKYIC6gCKkudw/s+TLIjusFBjSr7QnB1gLy5+y4POiOKJRW0EpgbItm2N6UVSlkawY6JA
ybXLt6nhbM4gSYDoTbY2DT3LgVGhO2eWaGy8SL88FYwY9WkT0UEt3eCGCm4RRihKOnGKi6SBNBC4
2X0tmcM/URpvabT8YLy26nDvkYt+VuIGxj2ZjaOvM0iP+ojAuHfSiplqWCmIt08t25pTy8w5f/b2
ABxxyXd1xCJmrjGZEqF1aDpXATi1Rn54JLfJck77Ti9RRB/wbsbemB+/m0FMdR/ie953i0dL8k7y
OuQPH85Vtcw+AWEmRMNbLAPvibV0AUFhaslymJ8KiII3LenUuJ2Ffar+6uYLci0Zx2ww5DJN0NgZ
mIBRmvElJnA7s6U1cPzM724/C5I6+fZROf32EDza4YsndeU0C0YduHF2ewSTZ5+1VYeTIxAFM//m
38eNh8Eh0oy5QMzRkpYgtJetUXD/6A0vwDiTXMx7x54Wb1WwGobf3LnnD6YRt0PTnSDAQReO2V2J
NEPiYya1JyykMITsVPwVf9xlL2UEnpRXpjJ9lCtOmNL8jpOjegxi4BvcRUv6ns1Pj368/k4rvbjg
xlwX5CJmgXUdRS9BEuwAYCaRgVoyZSnomQSS51iCVntXLxd0EoCRvl9CRdgQwQRi9Fmgotjk7b5A
7z4A2mjfqsUIazopyZ2dSm+YSmEdf1i4ZrgL0D6HBBAQT4Txq85MtLgJeTvhsBEeoDObESFyQiYe
VdsbYgylT0fQfRL2a2df+Jk4doijHwms3+Xwmz6z8h7jAdCyvklg8KiritTATz3Q79C325AWYsUe
nD3SjvncgkyoAVCsb/s6IdJlhp9IE7M2KzNvnOVd2epaBaDBt0Fy67qNCQ9czBgRMRYHiSwB6c77
i1zziq1So84l88So/7QWNpindRAY77AeWlw7SYOEgHi7/HZehIvn4qw1oALl3PaoDtVUF+GtMJRb
Er2AifNA2H8dGsbrY2o8ZWu2leOa8rJC9RKJNxnw3I3xNG0tqAtOs/tepXqObbSswmUQd+fxYRct
LEUfdmD1NTEqCHOeDd6FlKXqNvi9XZIEWxnkkzAirpSr2+nRl8e4BTXduTedgJHiDLaT1FTUCHmX
7kh3Q3hs9/3NRPEQauDn+5HYVhv2UHI08kADsF2OzmqY7S4Px3WArXFQu2bGmls33oE5IhcR6jeG
Pjx+GPU/v9P8uH52p/khHReXtltNfiMJZeIxBqkDXELCQp0w/K+U0C0QY4CTyQkbAhwtXFLL1UYn
+dHawJWabR/hpHPrK7tU9ryIn+dQuPbZbaPwi/5Gu42ZsPoHVTih5oTrFBcVaDnD9FrqgAjvpemL
1opmMb7kEp1olvndT4ckBtPUvZIUea1O4+5M6YJXgNZWfYJKe8Knefq87WRz6oQC8m6seWXu0jgf
FySKRKR2vMLUkBWckK6gwgpQHZArXKk7VkgyWVbeGAHahgSKv7DaC8jNNNdT2gJZbDSjcWWnJ0O+
eY4dLCjGpsurLziLJ/Dy5Zx8u88vsOx9VWylMZMSYAQmQV6BjxV9aDPnWhaJqhLRbvFqN5AIHNUG
6zm+0uS8DZ5bZhIwjADKkA8AGVsYc0m7dupnoW2rVsTovqqI+tdASaYlV/xwwOLaVg50zN/+Beq2
J0lWPg3Z/+h2EotSrJGsghHPu4gnF3LjhLn3IpzKnbPKREMS0MKGgnwbBlyBZM33x5ebjP4UknJz
c7wKjDmR40q4Ck+byMcQExejb03YtkY59uaQKSBcf6MYs+ZdD4UoaEMnlsaBIcX6cLpjNAbQHyZ6
C7qW/L86Wsm1uOy52y4wg9oADC9Tp3X5LxiG5CMMMxP8FytpDqWFNAJY68awfWY7tZpHJwDB6bLZ
K3H/tCD69+EvA9gpHsjsHQ6PpwBRabw0VjtfYnptT2aLtw2IR10fsVPrZY5MEic/ccJPvBrQ/1z6
VzfLvvBd/ElQOSlHPxetpvhPcx1QK3fpjS+csHfrT9aC72rYrYpRPqidcaCjt381UX3XL32pbzqI
AIcRs3ZSTsBsZ1+EZdtkZGmwvgRfO4+m83eo1Kzs8pBpuc1qewWqf0vyAH6cFZaoWu4XZJQr4t8q
TbNgkbpPm8rgPKeBESNHjXyUQu339LSiUUON/TSJfoG078lGh2v6e2S5croP9GCFQiomvpIAXcdy
Xw3zzX8SmGF7N1VrIBvvTp4kxAPFBRTU0WTGsGuQEysFF65w5+xXuzsFWV9YGqCxc9j7DsbvaWYC
uCkziNfvJH2QunirRBYb59pBFsJtK1ZWnoZQqHcGeglR0Zg/NRYPzgssNenjpuUuyN8AKpXS0xPn
1QIdRe+wSt2lkFDgblpvyuYGZmXd8ve0LMtEAzIrrcfEl37IHLLbN7eRZJvsZa6GkZy8kKNlc1IU
dIWPQulKagL/O5JENM8GNwoQpPanrOB1e/+MVAMGKaP8MD3HlC8arfTnJC2Q66/wKBbLLxT/ztpQ
9TrYzIQQmnRK+JNT9n6HjDV+NNjxzA6qRKKeMUT8kKz3IlwR4ON0+NthR47nyeXtgYTvI9493jNi
d0DibAVvuq72p50WbsaxYGk0MU5KV2HSs6RxMI9HvKTbYUuKT84novCnVlQSGfoDPeqi5xYmRogj
yjL1wEoO7tz5iwsT4ZK77HvF4/pGij023lLwI/RyiP2gXGUzacuCnVxyQu+a6igFc1AqGrEa9an9
wVu4WtCGplXz0Ooh8sgQsN1Ph6sqC67SGnR+E1qMCnkIJxd985cV+68r16EXZ7wZPlwXoxFNK1Dl
BP0PTXj5SQg0uCqBVyqpzlY+6v+XxkoTb/OL+kFh0NG/5McJxMPWRLXC2VpzQwT1We43AZmrpox2
axaPY7WQQMb+0SjA7JcdKQnf5Pe+8+Lm/DkqJaqPgD/Cl6oaPDktJncRcK/Ni6u8VEgQod51ktRP
UOad7YQI6wgE+GI3y5gUcNl5+oTwGwGPaPduvYOelaBexqMYcgmSEhvcAEWelLeHk17okMg1vvzd
BhDaOwoiX6kJvEpWI72+lyj1ZpQPA1PniiZFJLY4rVpYyNtAPuo3N+62OvYdSEnj5DPXENsYGN8g
HE3n8Il/Bve7utntf5hriyp03wGBSQb345juuBMUKKUwiBgVWAl1V5I0hgrUrudXjAiBbYafY9Eg
iaDdqak//nYzE8qp2z2ry2QB85CxoNrDzMeTuAlPfmDFszhnU40yaBDnezavmQ2x/POdkCaJbv6Y
VVJlPmhWDIAYMYt72oXc6u6or9dnk4vB95FDep/6F8Y33AUxLPR9g6fBjCT4lme8Loa0LWVUDHyJ
fSn9KwuRn0hA3s5ljeoG6h52XxOPh06aIPq/32BELdgdm0K7+e1XOwUa+v7JZ54KUV4xDujK7Wgj
9Ga7nNhn71I7WoJUkY5lRbpf3HBKkBZGT4/ss1EurpghkqM0Gomv/PMQ8zL6vgzxuXwd8RLZwkor
ZYao3veXG95HN93CQQ2WB9Cwy+Q4AUs/RuBBuLsWBRSyf2O2Nvhviz1xM8d1ImKJp9HaHw7Lomfu
VJTYuXUBbg2FOKLUVc0ET7HA++WHMf4R1Eb8tyKrCbm0230sdCPnUda0xdZLX7tRhl+qKQVXl4Cu
d1LY31yM+OqpNgE1xyCgQXhdOOc2tzjNx50PvGu5AHbWUPu5lj1vORDJWR4vhPWjgZ72d8LacDH4
8JUnzWmsTkNKPMZP7i1opbdgkAXN4pNg6n+TlhcJKhiHANG0ZzS5Sv8I8PvbANtJ2hISUMrUjndx
Jj2mVz0C7nL1sdUpJiYpkHqBhvy5LJ9Yf3wZN4YkVYj4Z2xHbKN1lJBmpCe8q1Zm5rOa3gPpOr4l
qok+M6RBwIf+xUytjlVkUonC396jrYFEvAkLCexV8npVmGxr7kSQTCGhdo7TYqw2jBmojexJRjM+
wz9Q1fnW+CIbU9CyZSdi6j2vXAyo1Zwq8rEvpgYL0RlkMHIRQga5FJJXY2S3BJEZCmki8VumK0s7
G9UA5jC9MSg88JkvnskOFi0bX050ci+VLFgkmEYQIxRH4ZVxZ3CnbniM1Xy+p2PLnmmFJchPby2p
EKMZmBkC5m6CeyNvl0EjIsLeFo/Q+vmw/B3NNh4wlCfpGjRQDZ9zvcmzKri7r+6HAaoN2a+9q0Ix
Q1bskkFrYvyp44jeAVnbdThwAlazFmwMPSijlUZcU3Z0KPRV9lIaYngZtH6p2Fnt0Ou0nkpv5c2U
JHc4Itl2mblAwicy25PjOYaVG2F5lcz5u2nWtUr4bHhhLBJr+ouQ6SlQMrsstcWjdGU1F4bzHezD
HnAtiQOWDPxmFiVEGP8HXM6SWfYDrTPwb5G8FXI/P8rzkFQ1h6sRGauEFVSaljIM3rozN5jIAnkt
clbElOBF6fN5exgcHn9yQJVRkNWOgmSJ3E6vANm3o0kBRrW9C0+lLIsYTa5iEI24Cyra9op1liH2
eafAHCxgcu66dwg+ZXLsxi6TNqTi7UPfEBALxR8yPr/3KCuOeSF8TPg4j16bFlP4c2YXq/rVLog2
wZqEehVQf//ECPQfqj1jE98zCtvBKwliMvbqufe5BM4hq+Nr1eTnEfIuViIcDij8oI1W3aC/N0l0
Jvb9Fr3e2LCilWsz4WTJjKbopDaSx4YxeSJ1N2IgxrDRgQnnoMgd82rE83Q41v2LmTC9f28hMVOJ
GdVP1hVgR+I3dJhIVAWqG4t9p2z3oRyGOOuoXAMInS2n8GvxNFt9v1uzlqs/idgQu5b3QotRfrL3
K87X547zanu4yGNsP7vgla2K7GsimBsxiqa/Fri+CqGyDVpdld0UhTHdVBQa+K01qQwcclxWwmNj
gTEfGCA3sXEkJG/CnMb0xEQYMrJ3Z2AqaoC18AOPG8fpRebmgePKp7X78hXq97Fre/VvCHMnNPci
0coHrUHhwM0kNZjIG/hDMky2ukJw95ehlg7Ee3BkW1ICawjksIZmVlRz7uusomJ/YvUar2Pw2dTZ
Ri2T7YxWBE7JaRG6ek8k5KU2wN65DYxGQtQfJJKmaEagKjOMhhlQ7IoW3UfWEPTuF1DrwOJTqKsP
+7ZEsWr5DXaXOo/3qrHy95FxwF2xwVX/3BNnv76Tw3qpLOkCPifFyJASyipYLRYmkwZuWymUzUKz
QzAEZ8KXKCOewaCe+J3CxBZz0XplU9itwB9KojxByQl7dFm+HuDfj3JexxcxsrT+Ez7WL/bYDR+7
+CA24F2D3LgUB8mbHx5wvHi36o2NIfnU3KA18d7QpjtbB03LmZrHIRYIrf1iwUle1kIJRFE0Xaol
7+GcjLcSQz+PAdc2PNNT7Iu6p7vqMMJxp3gUOSP5RzzNCQd0BokzvkLw/6DsWxHoXkUHFH9XVgdn
64/ZM5s8X1pRCNopLCb1WJs4+CxJvu98Dhpc5FST2hbbbcBd/VZLFpBcMbJAlYvh2lF45Zy180nS
vLFmOgeFE4P94zvwm3TLNmYOzijjeweEZwFPfbFsTJI0yDmFheiCrIJuphhoRbOQdaQPu+3qjBfE
B5Lrd+tClO/FmXP649tWcHC4WmmWo4xTjT8/OnMR9tE+Llu9EaegwrZ2wvNhGr6l/rdWCGzuyEke
/m8RTgGV5AHAllanQAFQACiLX8ddELGPwhEu8X1bifR8d3BFTi3+CpXtDfiLfuqzav5m9hMuXbEU
gSTMgmM0vr2HXtUIPAL+gNviMJ91gNPs/k5g1lEPgYoFKbb5DCbHj9fXyuIa+ecbcaLcEYbcyfNs
vkx1pqK4RmmnpVdLwQqOmNw8D/hsXAOW54kn+orAWklMddC3df1o4EwVsb9vzgVLPWqOtDTWDtTv
/gcoALXnE7hGxc1sFiCwcqj/dMON0peMcW5uHkffdApo4MKf+C/0rQIzqzH3d+fBv+1XepSeovjB
sCG2fmAudeQ6HUF8l2xyaM66iEdQw7s0Rl1Ti/Y7SWQEptvC+f1Z2VeCDBzuDQs7maOfF3IMG1Wh
FQ7CcSnPHaguR3pg0FlcPX97e7bN3COkp+SW14Vnr+MbDHnpKkigaKrfslQWT4IQYLzDps25D9Da
mC+zM0oAAY1zypDWgyZvC+D2Ms284aZu1g6Cvm6wOhfzYcyN+E1D4e9l0VyZTf0pmblgwYWOvElS
dZeNuntVQ2xLbIMAy2+zv97tkDGzCxizEOVnk7VkwHAr7rmQekTC/ON7hq7GkQsFeZ9jY9oU3+7Y
2FzkTgWsXq8W0QxBTDSJ1Zd1eCsEpxdQhexGNrJaXg4EBVJD/h+PrdX9qSiz0hZBONdm6R8/RIzz
CV3+miTUmRk4O4lp8K4b/O0s6rXPRyGDBMVIs4TlonykMbIwT7Wt9ZAErvytwZz19y0zqSx62E2K
79dMEsPBSwYHXVPlZT81eXb1rJphp0YKRCMe5weHlJMjKHD+rj9VXYGdpBy34L3geUygxH4U7xbC
stmqZVpHl5OmUKB5az6t9xOCgoGvdSgyWVHRXTCwwtIpyNWWDEBc3pTLs37sjL5uvRlBgg3m6YKc
nBf9lVz9b0mfMOfQLe/ttRn21ZY8UgV89DVFDwCnrFeYwKkT2t9qRUsZu7fH6xgexDe45PHQODR+
Udmys3gDilUYCn1ZklAcChfOvVMq09LPTGZXe91FYS6nuy5TYhZI5aaSIqY6zIBinTYZLWXQOF68
mavp+GurlhFwUoAyZEJ+C78XR+ENgOGF2n5ox5L8ptXyD6+iZ2HbxvSC3jaxQ+0arEwABeo/b+cA
C3rJJfXCvfnWNH6t3n1+VOI/sxFUiWMhmtiGsseE/fiOJBMgwyrTD5aET+9sK1Dmy01XlYf7P9FW
g0xahbK9D+uUBQ8kAyeRfnZl5hiX0iP/znSOk0QdoCGs/yK6uPtI0acrcqWXfHVoBRt0+WYLVd0i
16I2XFbajFvX/OT+9i9oGGmeOxLZYfmWw8XS4TaOmw8SKsgiL//aGVDlKxfp+rXtchGrXaNJSNVT
Fg+mt/g0E0xijxMHmNzXyPTMvTgPmWdMG1Hhju0cSBxymDwBk2ucATI2v5fPypqbTczOoTW1TBB+
NTwcYm4KI8Dj0O89d19UbAvL/0FTWONQE5oww21TlM1M2dBUkRIUsnT/c9aY//4Yd5om8QAx9JVK
BEYqI4m8rNpYUG/lrMWtPkTkXh2FYHftO2Iupi3d/hXffWPOzgzPvVhyROXOQ6iIXYtTMVfihWSu
/JD2etufPmbmcBgJvkLKbWiwOxs9sQQsIS1l2uS2CdPBWwfz9UIKYjeNmATx8klNaDvD4+D78U99
pEDwYnevVQ4Khlvz0ptyVflaCHBp6xUgYAPBzRRdQ3APV9Iu+XeVH01HrKgS9R6HMHX5oFvacU0h
wMWQ76w1YTpX8CVvimgSsRU7o0l6u5su+wmujk8ywzGHRcezSAGj244favdnpyczvOkqVtgNvpL3
MBg6w2TqC3CovUvhzlIqggHO56I9T7PrBWbhEUYfUvE89lMEx7yl3zz1UR/Ze1YEXDQCsXaYfOjB
Task5lXIPDChVLJK91XM11P9SMSmJIkK+ar/bRXxH0UufDEQ157przpn1yMkEmiez5/bAagv0hjH
BPUAR9NVQ5Q2nOKLmy/dzyQvRXCIiV91tw+8TXg7SjbtHSZBVGgUa1wDAGba0cTMsqfoA9EYOH+x
QUbEREkWG43CrKYaMwCbA3v4JL+6+WM19wi8YqwazXlNEoUJFT6EuJbe/1T52Hj/07mFZZPbCrw0
S6Y6wtvMmRLJB2lKQwMwZdEOjVLAaKdEJpRSn7E3FPvvWYvYe+TPFmziWNyCIjP+2BqaKtC500wt
RhP8wkcknW8Yi8ipA9WiMHYmpsN8JtT1in2XkD0BovTqFABvS4+rRe0btJIvhzjptnfdfE6YI+C+
oYfgFEDPK8M+Git5BX8fvVKng09ssCBmNGNDaBk/wUsI4KGjzapkPNZGlWwQaf3kM3RAlpe9uAag
0bO4CWmiHoZelSCk/mQ4ECYhHGfFI1dpp4ZmDWUJbvYSDzhOLPhWx0aDLP+mkq3RAtUQ8YjGi6bC
tUEf+VnFtPt98LW1HmUFujcCBc//hnkv3v+LY4GftgMSu4M2oaELx6rWkDS5/M2foIRE+D2PGRlc
0aoHJjSqydPq31uayvtQIqu/FG8Y2dsJKB9xc1JwgX201i1wXyO5tct/ixevBauNGjcfsOjStKER
vEviqJseIM/ATOMTJ7ktMq0OFyU/tmI0wMHk9zKbOIia8yxtF4TJOX9WuuZs05U4nvLIwJrwwDVV
E/wFt/CHSZpCgKVhBfjUKtA/0Wo+liY9QqWFopHAxvKEibUseHrNhc/2R6+UrMRt7hnb8GPctDXr
jIuyJ6qP0bYzq9oi6dZ1SIGFB0e96s5eR+nFAiONRcq/anN1UU7CY/+5lUDTVNinwV0eIncDmnUN
sm72LDzWvIPz9N13uQife0XB43vVxAf+K+t+7bHbHU05bMxLxaW1kf7OEDF+mi7kUgtD3aUNs06y
ko+fRlfjrdpmLsAmo4aj6oKd7K+UAz9q4KzCkk/vW5wIJC0DzJw2LTvtMUKe/QSrVvG2Jt4vxBC/
IvFxwc0Vat9Z/qAtGKPxtLKwqArPGeY9Osz/3scH24DZo3ZvFUWC931vdEebXVv/ozDAKnOs544i
YyYzK+TFqhhxddEYt5F7rvrDiav1nh/HF7lddBvPnQR1Z4IPC3DdEhsZLrVMx/2IgQ6MLaxASz0a
gWOkEGZ2pyRxHjkBHi8FI6jDayFduh+3f/I6QeNcREUjglvwxUmzLbHXsI2HkCEuAb+80dOzVFGr
k5OAuOJrlW28kIcz0Bpf8H5C+f4bbp5MUOiPLyFZ05mbBeZiv3anZw6R2tFl7Y61YWR/LNKc4GwB
E1EEl9o6xF2ffl9ITgMTxRFCnJgBitTwYAHaWOphuwYZmRusPyNJ2f9+z0uCVZXMShTZw6hiX1WD
kEbEHfqmVxgypMPJcIs3rcuqkhGB1WxgjmM+FulzYYdZMAuhWxUDRY/3C6bLS/fXG0pCZ+odFfx2
pMkgVP7XYr2VvFHMrEwgWKhRxe2Dr4M3lQl/neCShMtngf53S8JvIqlCZmobR++nJy+mC6xBMDkH
xUOl0SI7iMObe/SZtt+IBWgn4B7pa8lmAZj8m+PEj/mXFCABMdwb/hfMA0xKtZ+gj3B9qd62zl88
CKqzt58D+cQT7PRtIpDeIiBGS9d/tGfPpXn3lC1BK+zsWBcjBz+JzPTVHITTcIZBQJRoX59kyIiv
IyUcBIw65hZma0G06K0RYMG8dsJrB9ZqSnJkt7+OhLeq6n2n1N437icmYSsbgtiUy9PHnSI4S1K9
Y3hrugCXvxRyi1V2Q/C1QRjlWiHZ6ZC7tBPn0QW2wEwHQxHB/WBoQqZZ3hATygozYAKfvVxkTShg
Xpfm4zWId6H085pM24+QHmIu+UBwlywqbeInnAZ9t+Xa4cACsRLbAxcDv5/l4UbTAx/YOpCot8i5
gRi/Plin7wPM/FzO3FulkI6gElDHIGL0N0UtPOv5Qq24S08L69zgbYVMm68Ws4nRS7c3aFJIy9TI
0MHeyDTUZq8V0ggydxklNl8DZrrMdPLymxJx/RllNsDeCZhtun2pi1RnTqNGJ6SDwYFtOr4Zrgvr
HPEtzNN7X3KZMYMDSWlSn9OtPix2mRhAuIDm6R8qIhK8Y7/CZ9GdAyLx0xYSikN7/8DY5c+e/TB3
PSutP4LrGwtchDsBqXqlIV5N8w615GKxgprxpeUGQxctbvALcvt8OT78j8sK3irviVMkt04li7wP
YTL5byO6lzh1EtXSJ//uLCjtU0uExegfVIlSIveR3Lvp0q9HIh63a+dMWRrS2MnVL0LHwizRxHOQ
I7mJ0uDSZjIythZLRiIetclfFS7reEp22jSwziPL4ocH/ApL1COUoRVGjYApZbA+wVSDwbUTkxTu
Jkvpz/H2Bq21iUzANSGN+5YEiMsr+SFFImaRjr4wHdiW+g28hyAAMb9U/0bnqIHstVcsM5pmqZh6
OVN27CWFa/ssnSs/7Sxzpva2gXyN9ouwnh4w1/x9INSUd+r1eVHH+BdyzJX6rgFNvzAJtSSxB8et
IzFBmigFkkyyULjkoSOCDOk9vuB83eaUJHgIL7KkdUN1c9eClTgjDL3AvzWc8b9MxefWfefDnhOZ
xA6JUFGN+4SGkr++8YHGecKVDxLJGvytSt5IHIk7lwQHWZ7aKpCt1dzBSWoJqJFlyaDSYO8OtJwx
MlFVXrGE02gKDNcI1/gunmN2wk5q9KZ9UAxr6nUiLfomk+0gjtOEcORK46nBsWDPB+ob+esKsjya
tb2bfOnp00GkvEjWEqtj2T0a/t6IS4uKLZSk27s1SrOxEkYUbfeO5G+9Cl+bCUHzt+qMgMHbSKDm
VIS+HYc48U0vkWpGpTEOWz7xuPX7E64/pf8sc1A2bvRPsqJXDuXnsQcjmj1/hAIGCvcbjuTLcLhQ
/BSlcWvteDM0iPf3g+tAVP7BzW5kDE3ck7jlrRxexU4muw3pz0HYhVHlOSFXkaRxTOn8tHbXD44s
9uLrbltgcwUSOp8RYTsMwOeogy8EHxygLMIeUupnwQAj7617Z+tNjC8BIVkEwqoANCHCu2wwoG/f
wX/0N8v/pj72HaxJqD0pFj3Oebo/NEhGNY2QrrlB272kS5nvFCgkZOg7p+ZX//uiwX+72R1RtcsI
V7sV7Pd6v4IIiCnnoGzHp9F/IhrfHJAfmonRAZQl0cS6bj15FhaPZLVIN2sJn1L/0N5RmegRDWze
o/Wxdz6i9EHcIDax/26xrfgKVHrZyHdB9QbZdonivvK4jwxDstv97B22Rox90toC7oxOuR7303bV
Yr1NMv/2fviOnFqlMTHPP/XEH/KBw7t1N/AJqjcn3Fxq+RSjpgfjorgoA8obsYP/v+bD7dz3PhD1
1kWAVfqTrNSwr45w1NX1A0aKia3UMK4kWnJprCZUaQ6RTN6vRsJfrwGWew+MdGySRg8AMnVElhTQ
8f72JXgBXAXQztvLa+NzHVLE6vYSNaMaPGkUH3xJjPPBg+6DE0rLHRGNMemONhRuJa0q5bAygab7
zHYrwSpQLgasyXdaak5CfmvMaZ2uc0xlzCl9VuERR3Ux3f78Xj8dP7wBfMbBz1L93tNqjmVVuXns
phSwLLwIz/wZyRNmvH3TznIGqo4ZLAhP65vuc+aCpRUFR5AL0PX6akNNm2YbGW7RBR6VHlPslxP5
cbzzXmnFLqmLfkhGcBB0sVQNfoMzOMon9OyIi6IMPWZBPOLvu5nij5X+fw3E+d9UaQaoaatKfoKw
yTcAewIRqUm7+6MW6oA4Ud1Gr7ZZUOnas2uVB7uyxo/vf7SR/oaHisGltvrZHCLpn7oSwnXGy4gI
MBAk+H61VhbcFK2OKSRT0PQASOAxvCyITGpZSNYzzroU1fmN/sL21Ky91B/tTHO+wfm8zzMt52tT
X7VZKir6ygdWnIyzl5KUMybgIguw7pYHroW3lgMHAuDqh9efT1iaDI6Xl/nr203X29524cPDf6gB
uYZ6B25h0b/5jEM9eN0ajddw23pC1Q5l2xajvFjdUV2qmjVhGnK3xo96XSf4vlZkheGJ0y0ptmJY
Xsxhebmcem5lUN33PmpY9Y/5GddKbh2OVhijCUg9NY/gb6MyMZhkKgDGvWm94mZz28so+YAZYAFt
U1VOr56TXYjQxpAfjbVAosenhFYJfxf68a5c2auaX7MSURLWq5Ukp2kqizvGZDP5xSkqACoFitxJ
QXPDsl6G9bKis5AQwWAcRlFf8y9slrAkVfLFSW8v3V6Mh/8N49cxEBOyOI1LgGNt1EdQUslZTOW9
RHJ/U0BPf8dFCqEyR+jaOHh9mufZTcgYRZ8sj86qF3dV1euCTRcTAlCzUhIhKGQkfvDgzpG2KTaQ
LKmv2fuZp6wQaExrws3aU21kwhKkVcMv/TXCkFhRX4JE32AlZ9nnS7Ah7lzF9OkDB0tLaNem6Yg6
/7I23QEVjMljPdFxUN3l39AiVBUXokDz8YVVypClrIil93vzN0M2puxyKmthSx8m5MWpf3zzjipX
XkQA9Hxv5ZlM0cjkS5CihywIwVzkbbE6yJgY6OjZUNEj/1C1FLrh4wG0zp3mel3PpdkpAWksgrl2
neOCFzbkDOYWBURjwKe5ZdgvRafDwP9eNgAa35XBy2nDOjop+6B67/i5zE/v7I8YAmsgZ76sLtRR
0mBT65qoAr9/NlBoqcG67PZRtttCh8A3KxranCfoQw/bVo3i/oO2uqc4u4JZoFbnh4TuVi0tqvz/
bAzYIV/v4otu0wpYHwH3v6JOUWA2Q5/bC/NSkygBeiWbXlZN2nCzsOj1M9KXvCqzr3ysikbhw0Ix
UACwF4vK2Bj9slihXSI7Zf29tNpHzY1pWsRPR+jfkiDTAvmpfetc80fEVAyQsKjQFw3F0Cu2HTXf
wfX/dBwx4havt5kdTsLbxA6Ci1ci0uV4MHoR7+jSP9cEI0onL1lZSmoU5rzdgwNcfekFB5xmGyX5
Ed5qh9LO+KloRLOHbg6PALqdW0R7qne5rZuontDoJWTSOdoj31mtE84n/+UN6eT7Mq+yedsgliIR
QwUaH9NGwqdKiGtUT0Uval5zvxU425CZicJZz2UDnzVJevBPPWbi8YffHCAU+dV4sXRxsF3Xr48s
r4RYXn7LlEIXqetJ5aFVRmKWwL1tXGWKSQD6TDQjdPeX7usDnvT4xri4mjkNz0sWzMvhgZC+PFVX
+qlQASkI16Q8Fy/R4IqYlcJo5hoBlR5iBoc3Oe7uoKAMKDMVbSh3PomBrVNOuJzzwLmkm5oC+8Ls
y3OoRrzxaSAodojw76Eg5b9nCSs3wVtrb04z9Ky0ET1rrs4gAJNShzwyPbHYUjFoQ3mIH4QQlLB3
SQ9IzXi2Bk5eqCAlOWrXLxDt0lM9/uTiUmHOkMLi+DCuSsWSNitMpuPoiwHGhjH/CMEfOdSUNEAG
SAQSjztaSPHnkXIPN5OgyApvXeD3OYjLLpmipuK97VMtGbKzUC5hussoSLRSC4wCozzrk/9XuPW0
8ux8BMnt5NqZ/fHG1UFg9j141pd1JAZ342Gu9bZWie/1pGQI0v0oDL3ZFYTUOpZ8EL4W3dRMAo0v
nprMx9qWY6YJoep36bCxOgi6cayQBUD9p97x0Ngdk2Jcp/qKueFe3Pb0OYOJt9QkDdeiJEHYGLzz
pdkQlWTbRs3nA0MgtYpyNwQw5EwzdcfOTo1Ua6FiZWI5S75m23uQARG/cBFv2J/JAnp6PR2CPZEB
k1bCyLsnHtX3NjJoPwXqjvdSiovr+756p7ZTzA5nku9p+QjsSiBlmtc1qzyfvP6nF5QhcMwkbHl4
sKQafKRwtoruJeWW5MjkBkB8qE/SoFaLj2RyFoExuVGiBQYcYlkg5H1T1L9h6Qw+U44ayW5x3GIz
WRtFoHc962qvnH/o6x8ZSQgZ/21xdEYaUI5NgblAULCf6FjrupQ+fYIe9pUK7NMUbQpVV5zXnjwl
tL9eCrrvJ+GbNNLQFUcfBNzbLQ/nC8m426JScOd2MllkxlMi+zD8BljJbf2u+rDw43J7Dj9xnxiX
iVTunTWBsvqn9W138nm6ku8lRw4xGLbiAtQF8U8laaY6AyrcawrEL6I2Fk758t8pdiumIFzEDm60
ndnTwh//H6XePvnPg6ywgQc6H0ygsGYVktV19AT4hG5XlaePaR9gLKiRMZLXWHrCHHOJA01sGhf6
wwtlt7QgNiJT0JDPGG5n1K9LsI/Znl/Ot8Fs1lVPrsaEO3eUjObOzaIxPa4Hw7CukR4qTz5J+8dO
f7Md/rmvPD5djFkKk22ybvymPPptfh71jEcQDdCBM/x2QUYE0YpbrmKrvou2Gi6ngkhHPZCx+c8z
8oA5uQsHGNt+HmBs6o8zSGI/4urVnXXxA4Ff+uhjdHmOVnKHqTQng3NbPjTnUu04NxNBg+bQHq6t
VWTiNQ7FLHqF6IbnSuvDrODYFNLfr66cozC6wpDW1q6VFZIiN63x/IYLi28cIs4Pt1DbzggMsffb
Q6dsSikyD5iEoZP3e7SKyP+w87wLynL44uQON/GBLNjVILtZ/MlYZ1ZRrpCIwH4+/EohIzOQ9pqV
xAoajvW7SRGTZ3CSH8l//o1qDai0Ij+jIcqbtqL8fMQdgKCA8eL9qI/iS7Gy+fDYj2LsafVPoaD1
nbGJddJ5KVxAUc+NXtrqae6H0mGAAfvkx1NoOGDwDlPwu4sqcuf9OV+Jib8cjJ24NgO+jnQdx6pf
jlPmpih/35TJ+rJv4zPZBjCpqYiIBvIRYAOKR+aqOgFbKwgHTUCPhtf8eT6dx9CWB3bGwbD8cjZY
inPql6d6Vefw0HhLdcJoNbeB7Qr0fLUCy5BSSOZGbw/BhiK08jESLAgO5SdaOYF07glHL0Pw4Dzg
ZaPfHUJUEAhypA08T6h6993yxRIP6SjFnDX09aRG3FFNd8u6nayq57kono48mEAfuTT9sdTpb/GW
pstOavwm15bW7i5mOYTS1VVk+Oe2Vd3Akx2G8etpGPTLIY9l9jzNS8qpgoZoaOSmCheCFfz3lxYz
+kNMtZ9nqIq950h/+KK9OzPq0HERq/nLXQOTsmbMULEeCrUGE8VfzdRuum/brHIqXkJiQsp5SjZx
apQbPUFO6E4+4hzqpA/rpclsRM5Q7dKKtNIGLIKZZpv7WetOG1oFwZ1gGxQRBcvbLsB0n7++xKPg
AIkKVOiT5oFid+iQVM+/uSnvD73iUrW6BoIi5mJDA+PM4rPdj7JGW3dULxEj5+BthSZd+4ujtOvt
THOUY7T3z9MuwxTuCXb9H122MTPBVtaSVnoMQT5m4L654dYymknZtmcMRN/DOJLed91LcS57saA/
GUjRrd/wPhT0INQR4AhwkoiEbBhUpdafodwwpRJedELVd0swmQr7tDH7LhXE3mHFZ6Eu/5oy0dg7
zDSdRrV4RRLifkzeZGNoCMGC0D+VgpLdhydudQbDbqXYJlAOCGz7OCIx1SEu1Rsd7mVQKvsFzh7z
MKIOA0NRSPf67nPVcgudcF1ofEPJihhT/Vp0uT9tEPThd+4pgGtVWPATvWuPRf/qcyHvZMCjX706
nKVwgwhDc5czsMY8dPUFEaXP/AHgT803/xfPSbG3b31ROjhP9t3lKeAqaHnkn53MADIcRdMEX5sd
9aK5gbuqIub2ia5YzoqHDrjsH8quxDjqz3+9QZeO8TbrikREi41ucKxOrvFvpwCvD/XUEM2oWe+A
RxJuBFyXUwmfWRjwvM0OE4fTL2/ErycCBA66xTQ0tI2TJuqNkhBpftkHPEMV8PR61oeTU1dgGDNh
i+QANdIU9S7aS9AKbb5KVOcJrHSmN2bc5n1yc6AWRLEAqiBOae38PEEUdNg04axeWG3gnEetjSVu
dVYoDxhTACMbeYVzhiPml9GqY39N5x7IdhiiBBX6vE5geZHpIJY6mISFgCzN2VH26fSksSDm7h4X
vaTgyTtCLKGGWaaqdZCggdSbv9QKQHAJwigtot2jXzpVwI8h9lp4UDlsvByCNOHu525EpjfT2tDC
S0j//Cfsv+MNKsboqM4MWIJBUY0TCINTvNkAFQrUdSXkjuR+eC3koPnEV9lWCroJZykvuJbgspc1
sGfly3kXJbageMN3OG/1aSuK1GJGBnAUbCSmiL2/oIjecHkBQbfZAVT7TBc53lXie1cWwlzZpCah
GRtpKyfpCXxa3WxV33xKxcAJiuZhIyoDa5NfuKa/0U0vLoUZc5EhIRc2j7MV/P7D0+hal6DZIhvt
1QAKQdzW72YrrxBHC+gXOxjzZFmYZ4ah65+k68tSpASBpH6DlA0RKzhbUAR23zShm9QwKInwF7VT
rYnG5mLu7FGHsuwNHx48qzGzw+HNKPULAumVnee50tXJJovsJGuaQTvejCxCLjyvUHl1214SNVIU
YlXwRBDMBHOS3EXvi/zmrCTDXFKIPM2UfJHD+v8VKUS4PmZH3uLquNZlEPvxOJCI7XddzToALMzN
DnHVyfS3lI07wTg7Ur7FrUTqMMqKnm3IK4eE8XmB1nWqkz7tqcRVm4AU9Vrtp0xudP9Gb0rCPMcm
Z0ABNlxRo79Jgmqs7bH6QFw5ZEREw4TDtRDWL+aiagqyWMNz6RXW3qa3bsoZdaVyW743i5OVJ15D
9mKXU4m1OnptGDst+n83m1afR+Cw/IuYqPv4lNnaqSkT985+KbbdG7Bxszbvl53md5/MOXg/tnCj
cIMmBfdWxecGkgvY/EhIPj+UhIv6426a1yv8Ym920ec/gqcLkHZkY1/p9nyD9QN3koNl9V9tAC3B
J1/w0CDNZujkZBqIM2VFkLh7GYsc2DBKE3R4KOA3hGOGQm2s945705iTgkipHIqm7tFYG9eJ266a
9AhN6xw0vHgHhYxbJ/RyZD4JCubUTwxRRqvWXcFdE1t+jrfrb4XtP5iBwRv2Cvf1h9ctiytyhHFI
K+t8c5MhQJ/MCEFmdXn1YDDEga+1vhcogg0rb0CWvqx1hSsn45nqRB8erHF4HCJk3EvDxDdGAnA5
p0BmFD+hf1t38rQQ9vgHdfAQ8xG6QO6RbMtpZ7K7aGi43PgvDLlRWvsMci2Pygig4557/dxKW+R7
LZU4lRpM5i6K4NsnCvLc+4tJhurgIdnWAyg+RYiq1qBU5ZL7B4bbDaXhnGcNTlk8qRtqbf/k1Ymk
8eboXluxlTiH1n5UcYsuyWCqsessZ+tdGp8QY9962aVeeVnY/9tEzOJaTcFka/eXXrcr/B9PXdgK
9w5SG6gc5zgz4fH47UJgRSYRBmuncglKaOJEW4CWgyHGW21YqlqWLfJJpzjpZfEbhKTT7cuZcPKM
rVo3ZdrO4EpC3byuceUVjBc4OEiD/1crdWhCCDgn56KoHVXXhH7BIx9Vlc5kpZ49V2VG7svA7IIg
O8jO5xFcQEgBu6K7vxXSEdi6HYsNo0eux16aoJrcsdAlsmdgOTyvOym6q9jQ9cdRl1xhVdpyQMzw
jMRJz/w33ehstKsb2JTscu12ZSGUaoDbt4f0+swcld3TdXeoMmh+Gb0iJPrBwVWEBL5UumrJ/F5s
hWic+5GERLEeLzqhQOhPl/1/A8+7pv1hqM9qn1H10KskK9W68BUmhJhRh4+Us9I1AAFXgXlFvWAo
yF/6XveLl7vcOYDcp0RAgIY6o0r4SET6wTR7nioiuVWsPhGs8yIqJOcwNcypkozoBMZWW6gLEchd
IATBGigqViOnscJHioF0AL4CBMXZdQwmaZko7cDv6ldlbnMOmBQS2d7WlFCDyxJ31J/DGcamHqI1
fwDX0a3LSdyYI0Wf/gGktCow0n17zosvUkeHpvhLJmT1cVJeBE4+9V1JcVaNrpBs252HA3cNEgJ1
l24rddI8hEZfH5A0YFlV+sw3C0IPhnJbehk1Dj5bB54Ld9KWCLPsYGKF75agkGG9vg83UW1vBydH
QCDjVJ+Mj/uYgeG7UByhW6pWC3wLnyWrPf2bvQQ/Nz7VM8+BooFoqtzavFdP1cdpI/6lfGQRMbUQ
H1v68cih0ZkC1MGlk9Mz2FNTbVGGbYmrIK3LEgmdBbNONZxSOYnheDQNvIqbwiVlpqSZs8HIMBP/
K1JPAfIkPV+eBlFdnpaVeaAkeNvjOkMOcQKsG4lY4IhJsMb9m1qnhtFWfiS8GqUyIKoybUCpe4fb
cflZcXlWxkwA7aYCqhGfSurF34Xqt88Pdak44V/S7RZed3yQ5htaxo9kRh4mcvm00MAftkMw2mGN
g3goY6uq9Mdza8P69RpstwUlOhl7JJ04C7BbMlY/C2OIpm/ArsQdkJ84/p5PEsFPL6Z51Ar9dOLa
Qe/BeYSv526rYjWHxOkFdAaPg+ImKJfMPqOdC7KkjwBuxW05m+wz3ac1WTLipPYqCt5O8lyDeJfE
VNFzLVlvrOrjcWz2Kgq8+Ql+6BhmL7pXEzZYACGRi8fg3fkWvCTBx+eW19TBPD/w2UygQ5uCa18h
9wJQENfCT2VuCqSgK9oiG1v68XOT2h0fSk2DQmntltKd8BP4JuVyMvhvZxqdrcLTs2pcWsV3Mz8E
1CGkrkmPIfP8FzJV7EUQHjvO4PjE+XdDNMJCIMWKHKNGeIGwlSX7LSDHVIhLL277kJ4Mrz3lrnJU
BgN0yikvE7fg0IOi4o4/TVkSpur5XXJ6XMNMEbThE3H45pRd3EtLGdsTDRqUlFrFkdtXVvZKT9Kp
MLnJCAcy+AjQ0Bme/fldAyJ7Qtxr/0+SpeWtTk51zBNKNm/TQkrvhPugsdcLOIoa5116djivVECi
1dTsqXotWSN2prKLKf/0WG2lzIqYiLpNbgJEuMVI1h+uyTLVOw5bAvkrKAMJPSbmDxaqiE14vWoe
hWRZWEphySann8xxMbXPS5nc74ubNZ6dUaNZd2zCxE6aocMX86y9x+vpTAmLi6hsxZ45oibzXKQd
gNE1IipAiLCD20TXyeC7ZgwGdN6GFWdVccxaqedUo2wIhHtzIc0eSVsvW4JTZeeWOgZncV0+ReGM
VjS7NG2bPTo0yn7YcOHl/JwwkqqlBFKCVjCXjCa6ixHXA1AqGW0gFX7H3fFk4YMIN+RlWEikyWlC
cHYo4CwHJeKmHeU4C6ifXNX0wgaHGtPIgNugrUXMVL+wCx7OEGluIr0tRju8cFXjB/qzanW0BsOa
VUWJcldeBXfIh+kbZofB1+d2tm+MlLa5HX40Pz7iGRGoPggk9u6Rn+H0sYc6uFZRhQe1VLmyn8GW
VGtWqmXsHorQHq5mBkUIr+toEp4u6DnSbUwBHKBEWo8t4D8LB3Gygor2PsIbuZ7ylwt0375xuE4c
zf8PumI1kF8u7vMyohL603FCBYZAQXIG4smyJjeSW6wSnB+dw69c5a2aG5kXL6iliqhI7BAn31Se
ki9BuFLiVPUYgtKrF7VYz/PZCSQGXGXm8KIgf7zMpEMvYk2a/frtt5ETBZzyr4bWn3wgEV9i5ZoK
ZYo0BH2BVJVLuvmQ+n4yzUnX/L3QBf3hRFK9SE/mIzt/bzZqFc13Oi0bGOvqe46ojNo3k3qPvQ5m
+R+ZxKdRWpCbtWGx754DIEOqff7nCOpMIwdfhHkVOMQq8yin5RFX7S5HV7++MfnmXarCw5lTeVTM
XChRf8MRhso1suqZCoSjmGHwCPodUIYn7kHRQDwpRqDwSpsfNAot66zh8actuyJXiwE9vDIkNkC7
bH4BikcjLSalPLkQLATL9THkVCeiTjO4NmSaNOEEoKntW78CLDzNnCu7rpro0CGRAR7DJ3j8Idoh
3QxsGXfr2dJ6yDtpFA9RSLw4EkrKVClLIlyYLMe3v2cSVPrr6jNaPG4jt564541bOyexlIB9HRpJ
+xauZfGQDQb3JPFbChzksxJCv9bfGTsmTBa0I3KXP0E6ai1qkwKyq03ZGf09JEoAbnd/O5+vDEpI
XMvx3WE31wSPxyPSv10aS/RIwwIzVYQWRx4ydNW2Y2WruEKBoJ1UQi+KKRbDg/gw+9AxwOQfpGGK
aC1z2kExJqNrZnpLwToJG+kXbndtPHqgmGJDJKW62hCUUcc7QJT4UZbOAq2fTic5vtfhecdaPY74
8v6Ycr8xd1abtQx8xOu+Jll5OWUScnkyU2HXtnSCEC5mNxkOGv6h0Raf7mJhX/9ArxnIXb3TjjF9
P5m57uFzmNJn8NclMc4592JdeFG4pdwXbegUucoxdoLbSAaFgMyg/WILul0Js8eec7aQYN5EPcQ+
VFg7ZHYgYI5BnaQ38txZdxj4Aj6fw5kVLLU+ZBgUucc1hDKepiHseKyP/Q1kMiydtg3MSZ1HfUo5
cDJGPMw9Ik2QdwFjG9gJMJ71JNKB06VGZblAj5pKnwqjQm/sG5CYOK3x+LFtzucwwFnax+Xok9Qg
U7+EzxzzCfo6r8oXP6z+Afgua3iAGiLD8w86n/NQHQpVPbm0LZ/Whn85o8dYZc9A8drhqfHfISBx
/tBwvwdrq0NQCMjEJnXC3m+x1gFVD88djxAFC/izJEs2lbP17C92kBdI303tAkIpyyFXq8s+AuFS
3oj8jPIYt2t7kIwS0WtZLIZ+pLRzmYA50qfiF8P7TyiaKwcu3WznA5KrkZvV1vxnZoCfKgUlZ+zy
h14fxVP+TZIzSeks17IPNqzdtuhUmhI3MnBGQ0NWnVRvXXAp4BDecxOHqBmZevV6FAO8dwgoQoJx
YoVUxqgxJaG1r960av2vWnv9osMrnPNgV6gkFrwCw0zlu5SA6EWbsAv19LXrFoJuSMpufInTxngm
n5sj7WaYRu6EQxrFuyNc/Vg6HAyEZHfaXOHUqrtQa1+2enB5XgUXkwAawLIQWdJs0IUvuSdMHKYP
CdyewWumQf8OM609mFQvN9RC89psblQTcY6Ojrfa8Yb1isWcAObCdqWvCA5lbNq7eGQwddBh/qku
L8o+k4KwWm8Ltn40TcUVzHwcYsBrBzPjzQzulqW6IUIhXP+LZ0x87ZzR75AQ6rSDOqgci1SPOx21
mL9DmSsdrnHC5HtOyNPe0iySrq1ZsCywS1XtqHpAgDXeFx7cyRto2nJRqPpEsEtoczb9GdHr7V7E
+zEMGHocCXjgTBy5KJX8NwB50PIgmpXLRTKxqYnpZja2gI1WTLUdAqxtjD/YP1x6O6fuchKdscNq
I48NOItYj+K9n5iiX2Tv4eS0p6u3XUqv4PDxOpb8cIxHVlRQyFAsViUzGXwOY/tfgQL6kVxEZWiq
JYQsChnBcpjDaAEKZ9wjuBqrwkP2mBJ5McHEVT71OMNOya+Hmoz2NZmKFIiC/JIYc/qyf9yq+zSF
0nKhQanHbd6ExAC7ZEQFTqRq7HmmuASlwNFzdIBLH4ZQOLBWtegE1H/2oCMP1Fm15vOAybqfJk9f
hOyOLYXSrV6k3Lx1a1ieuQ0wnOjiPq+hOvxsPOTUFWzDF/vaU6jDLcYJBybSxZAyv5HU1FCgJUTy
RSkn0EJjZKqZccy6CsSFGFfLHwY7O877jWBudwMtSphX6NcJUeRhvGjuu06vr/5KjvktLEilEFPr
cJ8SV+kaskl/Ogyu+7kaNSPqSl3ppUytGr7IgzsSwx8hML00eIVtCqRpaexTAL1wzWulbhGyA0fK
ux4eRiWiLlFwiPAL8xANwZWc3FcmV3HNm+vREv9sQDhuYPRfLER+aPzMqI7XYGmBORAVY1i4a8KH
KGu3t1mT03Gg2lL5w3+SRCJGSvUU84nzbgA+18jKfffuvjK4bd7oKnOHUUv9TerutT9csYnxC77M
q4WaPq2Hgm3hHRqEXJOhxCITNizBHz3e6Cd6Bm5NBRqgnI+615muId1R2dVRs/7X0Fxu0HchH37Z
HasfTvgSmz2vxp5CgJg8q6ewMqtUaDB43PUfgGdhTxl7yU48LHNq30KZLapcKfKWUSFj8tvuqPpE
OYK3HSSiI8WZNc+RcMAP6hJxmANJNv0tAH3HYXMw4+E0x/l1YmkBgu88T1/Szgc7wDx36qxV9gcN
G9ZdnxJPL3jS9Ty7ERVKO3yA93lKXtJ8xX1xbYD3FPPnLOo6kA3TyKwplyM0dW+UjKfavKBLLMRa
WpOgzXSllk+rMM68NK0GJhx65Vy/sZDfZ390PxnjSkkSXxIpK+j+XB+8pS7dOe+GcRSYSH6v8BNS
mwYK6mivv28WWu8kuyukvnRor5xJs29/xCDKjlxENPmo6HANlsa7rW845bROpnrv/EzG+uon0WyY
eXG7ObXL2G73VBsy3AycfE8Gha0WRLQEGIg+ikVOBBO4sMTmufj6lK/bJnegaE8NX3wTQdbHzRxO
9Cmf0+5BqOwG1CpIfLtXdZ2aFj6TeMCPxphW+atWGRTmViRzJieust7Z4XX5OD46gjYpbfVP2OYE
XSnBEjuAWF9WL1iMQSC8omfvNDHrHJAncD1MfdYW0K4ylZaPCJSrxVJRoSyhYZP5LciST8Qv1A+O
YeqHxjR6IRGLmjdkHY+WZVCOdTNbeHHjx7pcjYrpHufz55UTxsjmnugFsBGOfvqWBq+l5nRrx2oE
j07yHfS2GNBsROesu/+dkNjZidJ7reb1PWLswj0a9JM+MuCl5kpA0EmBmXgjFQLez1s2BT7vC8vU
sBqGqNj0EXKBCdN4pH6AeC2z6LK+WjrMHjpLCosUnNtL9c2qU6If36yT212U9FbvjwNLwrJEcEw9
J1OwADHPNF7xvON556j93eUhML3p6+/trBppf/BBG3Ix/VpMkHUzk7Izz9iA7uogwckdqzLBfN3R
q1ry40+xFRKLxOIU1Fu1ljVt8JTvV2yKpbMcKRUkSCE/nY/IuwuEy4gF1RV9WRvj0b8K/N4e+aha
nkRC4s77sx4HOTq5leEFaU+cNnKzxQrqG/nv6km7m8AerTXcSHFtxcxr+od41XEK5/qLJEAtxN5a
qYZ4Et/TW6ypxy/CRl8nn3bSN/qXiOIeiNPmvCzxG3Zf7UbHVgfOfloTFYiEZxtJVV/BxsGQ57Lu
hYgbCODPBVpzSmT40zLjJNje0SqAVZomvZd5kNf3moWXR6AZNRH6Bzn0z5OMC3KxjI3PgMisujUC
CEQFzANfFNZHWvk0KOayNqc0YLcu4ZJkJR8TibuYm44CZRLZThQYl4LwD6dYZez80EJj6cZo6Cvm
u2ljbCgcpcGBj8cmZhsifuGkvtdKYrPrRR0ONRolJnmClEdznzlSRc+6KxiXWvXaLwUEXWB2EAZQ
I0a2uVweDIwCjsVbLqurQZYi7Xgpd2v7FLv6NW7Ndoz0KFAPkOi44YDGIFuSNWJD5PEPlAh6JmBI
XgTfR+6m8eG/eRemNaTVk5fcXeLJ8dj1bxqiUTSPBtNBjDfBAxz2FqwAXcf9w3UXvNOtQLmtdDrr
8qIT9cTpRbke/WjqWCDSg6WWNHDnGfMu7bOLGL1KXw8gV63UTAd6NG0l2P9ShtgzEki/AVEv2S+r
Dv1opbCLnPVFEulYuArZQnni+xbeHqnq/Y9znuuFHaUbSzov6zz9/W3G8vncmuIr8K9aO5NYhuh2
80amwYU22Hn+wqIS9bEpcd0YJ2JqfbYKzTi24Wtw39nNfI+WZQsYL0NeMfVIhDo44KG5JW6D7kTB
cjw/UtAxkKs22NsHlwQvDqC7/ml1dyCkA/ZOBgXRhyrG6K8zNSyLbtH1gZlGCDEoXzpUJQO2PxVU
Zv+uHzSS86OAUxEzShFteK9VYWjfZoZUQfjMnN8TfMPox5pX68euFF6eJBM+yhEgzypFD079cXYW
pTsyp5ggMexMP/Oq77pJNl+Z4ZnkYsmq7wWW2Pymee5Uif0rOqSwNI1A+mdaQTCESUP/wx59lfTf
iWKklGYELDffaqaolKIa0mnR8c8AFyHiYNeeGKl9f0uUWSomHzJF0Ye8GkPQ9wpIGFITq38jQsVb
8lJGLT86BJbOkMnrQVOvrM4ldbhIj2bEPOSBS1ClRC6vaQPPKk50Vp8a7djYZ4SNvwNXHQQbzWse
PRoThLTal3OgsfCnaw4UO3hQxRqdly1JVTHOneqGWuYduzk0P8rv6juAvd4stmVwjcOdl1EAKTNe
RNkgpX6hkn7bmf4rZmUerC8eOxVampcD11oBj7AUBzxDmj3JGMgt6VK2LNkWyFST03be8PM/ALjS
ek24148pD8hP8H5UBtKw9LFu1ONYIX70UqjNHuAqMtxmjJ1peygGPBNbm7k5/pZM19Gfz/4m9UV1
hiPEnlLZtXWPQWKwsSjAPFxfs3F11sRi27ymgO5ID3BXZeu+RJgfD4lyFlSak0tk1vOR+GXY6g/p
rrWcLqmCir8/Dk2bDT4Gp0NsRW59UbiTvA1xtePWhIFmuhjM1OXT94xwwGQvbub9Ow2rfZ++yhH9
P/5rZEqGG8MyqaD11tmVVp0bAYwLwKGusncFMoT3S2JzAOHxTgbIKn1NLryxsLwn5XpjTPQM9MKs
foqZhh5z/BOME0e7iKeCPpeW97wAEbWkxinBNKmsn+ulxZouNxvmuyCfho5UeMnx+K8LMCoixTl3
4wwZagHG4h47Niu1Bg1tn/dy25XAVPPLS+3f9Jn9Qw6x+SSkP48wkClbwUGTIi/M089RKDnlLyL3
afWLOfU58wCRTEcsBPQ2SBDZcPy0YmbGyqaBNwvNnUAMUgErNhejkEd0I0B2bZRjdzpZjcrSjnJy
ACuFrBJUbQxifO1A6df49PdxKHNCVWacsWj/v9DDEIqwJ9ktjGxkwrT8XyJvqM+B0NM/4jZYXLnK
NWHo/pmi6UvLDQq7aDo6SV+zCdZJThs+SyDA2hyXGdBV4xRgjBdu0VGw7/CCqP1MeUgmXB5AT2iw
lYcRqneNAeDJ6jckytvAVwWzsLeqEHHpXBj42BDQ6MMcRJ+g2+ZpAqTzyAF+tB03eBGg4sN1IHm1
r7q0NQFmUhydY417uf+FqrHIdrLAnS2qh9m0f1US+N4tGmab4jCZmnccr8CB+4OlDGP9ncFW4dpb
oF5zuHPONFxf/LvWyVjEHbIMibGunq+Wq+IC2Vl/tnB5/7P7x4tIJbqfn/LADXY1WgXYSAH8/Fwr
W9sbZnKZ60cKzYBUuxJI74M//JvzQkPuLWtrGRuu/ourmpUigCa2AaMK6sCQgAI3RGkMXHmy2Wfy
W5mkavwl64i43nML3e1l8jqdg0ZKkbKuhhfcG6W+M27j2zZFypB3UcN8SVkZpRgSWf4Wff/rXVzd
+4Aj4z4qoUhA6qB9E/GSWXFKXaEhq1GjE+FBMLrp1VSET9CkncBj5xxAb8J6RVYQ+E4kVudzvIz6
+aT43YRsGEcGpNSXGWIkS2AltxPHSgLehYBzRsCD5T+h2AV1lTv5a/kPW5PP/pKQ25bgiGZkIrEs
xnXXzuF3ZuwmtGM1k0AEzzM8lZn1rDW9jDjZLBTRNLHsmLO1GKJ9DGeI4US0dgT6IqusoNwjnOMV
iTZEr5ntiMlvij2diwfIEdoeTrBKvWeYmtSnv0xE1CGSsbOhvY7p1c9/8+NzMkAK7hJdD2Yg25m/
PGUBwGaLtstiPlIWxuoOH4ysfAjlV11Yv/8Qm5IPJIYxUgX9WqamqcOtKcBvPumYzbjfTnZTKAzl
hSBhAh0aRC9W9mXYtGjudOpAw8NdRZlEky+2tzYdWQxem0FCcFnSioUhToKw1MOYZFtjo+ulEa/I
qXtKJmb+VFEZgLibuv9mtf7BJOisdfBXg8Fwb7x0kdhWBns732xj8Rp1lrgjGecJQgduAe1J8LjY
xqulnHxmQcyZi+Vtqsjsuez4yoZQ7ItV98AaAyM9IaLUGMra/TVVi7PneF1gL5h8BoG84p/a7nrg
3hELZ2mDcgZcUi2ay99Wpe4jAkXOTqLuXLwZB+hfujGYaBrnUQOtcxdEQoVCi/KPSkKqME4ASIGx
mHVH5nd4mmFXEGyYp7nikomZUDeRWdqBgurWldXlDg40nIN6mPVPoNx1Qb3J7VEkyjpsqq6kUcNC
jbDrhw8F2VkPvHpu2z2zwBVyhZomItCVGnslgNj0pj7W2TG0Gb7lpzFZeJSt+l3bRb1GBlg0hbqU
Aos5x6kUci/aTZaL5Xc9cKwJuDlbQ7YUDWXFlIsylX2pzX5guiHfAMNcWe3Igk3mJjaqnyOUU4dF
0DLGXeiRrVCN/YYo+4jfuaJmbGr1B5xOFPQG91aUcHSfjse5lpnWz7SZylch/XnACgvHFTn+6yMD
wRSwJLPQbfuaNCO6B5sJhMmpadc4vtk5xE3fpDhg6tu5jZAO4qpbyzh1XIDOcdmFGRF+zOrJYMkg
H1NJ/kS4pr0PdGtsh0uyLavRevk4EWh4smoSeDQkNQ87VQdmWuIKVzWFKoGMMefLxmJWSkY8eU0P
NpaXM9X2P5FjHcKOZ4IB5odoijnKFyF1VI9p1D86x9Ye/ZNJA+wUOGhbJCY0pVrVaHtNbMx8VOdt
tm5jJ9vc3o6y+lSXSq2Kp4XjPMJbsgWlN+zgIlZ2OqKcUUp7YQo389juYYhOEZWisFityN1xf19+
MdgtbERnLCwX70azwyysiF2IZ4Z4Azzbi4QH9l5gM82PWkx4Isw1onAUDtNBfJWx46/+PsfNMX0i
Qms7HtkHNutq1YIOuXbvz+FRbo5nFhYm6r88Aa1ecF/F7OM0Q9G0VUg+ZBj70Ue9nRYFaiscSjNI
5qPwpai/H9rsknRZmlGGo897ZQX2fICo8ZHdTG+NwCP4SNyhOw+VER6NYVIWS4jmcTeoz/z59w0n
2yssRNcOzY4SimNjpFvz0ya/5X/SikMpRzUANNrW2q/vS8YXWARxaJM8gO9LR3cyDUtKhfm5pd5f
vaSu3WneioVSTfPMDNnd0aLQaS9+KbL90QPaM2bbJrlcZLDkR4B834PRvQMbe6BQl4zI4TzgciWm
QXS3fLW+/UtG04cn74ee68QSKZLmq2HKVxC++SxYraouvrTswZ84qXC70Y/HVe6CYz4WpoGBDy7Q
Dv5hFK0kvXgVLkvjrsLFVV6gtikm8zNs0TateLOZaRUOe2oYq6TQSSvTcN2yj1VaVImO74Shbgb8
lB5wrjLNLuUNddruezlCmK3LRELJ4SalZA80BpypA0VRYeA7MrnCy+T2b/W2gkvW5Wla9YIXvfji
xnj1syvwvZwOoevRXwTZj3MIl7lrumuPoPItG379EOxLnW/5JCTxkcTEBPNDlfEbTyIYColD+SAL
E0gqHS3KA/l6borENdbYBCVA4SOySyFYMNbkl71H1OvXIi2XL0fwbkROlnSYjEt5RtbeQyqP09yV
lhIBqxSJ82lgpA3udKhimTSJwIaEwVmHQPXIBGVRyir8ZAwAFVo0CbADfRthmjpLsbF8iZvPvusM
MI6O0/6JW3rnowqJpW89czQdkXT8sQG5Q1sLVcziEA3uDcSEMCbspb6ko9XBaXdpk0i37GAuexv0
l/PWt3JPA28wKulJHhJWWgQ/P3NNf2gLxr0AhrBrGHkXg73ioIkmUbRvmKfgcP9uLhpQh9Sz4cbL
KBE20RlSryj6XIt4/f9hFuEJpqo6RLv8Nh11visUMYOpg2D2iDo3AKldvBDkDXa1hjfzsAI8MeFs
mDg7zHcqM96xuciRFuRFjZ7qGtYBqMTnrAr292qrIYH899ag1px2vC+N/wKJXDWrPy/pXEkAPBfm
bjn+jFKhKp1tOrJL3mQYIHSX21IREqRgSYlp33cLi/gCqwFfWdZYubL2Qbb7bSLDJmT/f58Bn4fP
mfp4MWE3nP2P8TRgkpf0SsVYW5Q/xU+A9a2QoOKXyapuqR3QCnKM1Sbn0kOWOpuObbdYtI6uX9HU
2ZuWdRVYO0Nc5qyZH27wJbccMdGvSCDN6tC0/mpQWhctMh8EkRtLlZu2Sv8hkMcQRXoFBu/7KXMb
1pBwDSN/pIBY4mqiyMVhURnFqHW8j53a12nLA4Vnkh+dd2MDx8SBechk5YQ7ExlElBAcHjvFvFBu
5ASINCwCrWPhJvvVQ1Me8Il1OGr4vb4Gg3b3GaZxAPz6rnfrBHyN+ERLHC8SEGrGFbJ9j8UmQLKW
RO8JAn5fP4qD9Xs/1PD3HlsnLkg+OtQQXZCRKCXf479lxSixbcoLi3aJ3mOXCfAW1lRNad34dcX9
IrXi/Ap4bIL/5I0NqvhOXJcD880J5RLMwu/SrKUuIWKiJZeu6QPN5zOfcisjIcf0mELA92R5nCEz
xSK+Vf2cwgP1l99yfarEELtR9SoIUtZYKIqL284hWz7OiC6kQjkJuFpfa5BOhMP+IaxN+EQSvhQu
/IE0hRWorkB1AT2I7WjpxCjzzjw+5es/GqxjORgqw5nnlQ9Gms+u82gI8U28MaqoTc119Ubqz9iO
yPnuiavAfEv7NJzwWU3unnHEZeyOC9IxNttnbfuTuogr/LwxLJjuBtMLeojLHm/kNB/ZYIEQiKxR
/XtxbIMzlEGMzlBf3RRka+2bLXpjDM5waFTICg0DaYnk7BXrPGdZfln+y7rtt1iZopptoeGz7dTd
3Jy+dVvJrQ36csNyYqeQN1tA3VzW2tBK+7+J1lsbnNu29nqkh7QUkI8nxv1Q5SuO5IA5zHsB6w6P
DcJY6h4LufmOipjb6xJS3JyaLlckcqaThIN0LZ9Bw9F4eQpzF7H3+gzzHiiXPcNN41iy1Ml8lAJh
kkGP9TJviKKh/8wvhmIydrt/qmNfRj4cuk6o5rhyRFzXKl37M31XI/H6piKY6mbXEvqh+PY22fm/
hB9PHWyabFnGgRpDcniB+fRg3kxqrNfbV+pQC77aE9GwgDsiyc3i7Yw8gGRlfgZTsVOzi0sq+bM6
ozj/ZGzqCQTTurkTEqHsKoTBXGMTKVkeDKaS/DQb6+rLNM76rs3tasrd6pSbaNMlp91Vs9KA2Cx8
vjNG6OipWPSF7Iu2CcZriLCu+a2DFuEMVbHfdXIT2LCHZE8+2JUtr5NU7VsS/5DnkbogBuTIXgHW
w6FFZUyifgqo84y1u7b6lb0mSsMidK+hgXroBzQSdU68OM8d23PqplFGu6jLRMSChrc6NZUiboG0
50f4f2xga+A80uLCP3FQ1WyZ7ZqLMlM5Yi64796stPU9joQgu6T/J+o5KmsV0la1pffVaQA9vFLe
3l1J/m98hyaHmcm99gwLuYguoRUD3Kz4UVw4UN/kolprzObZ1aYwcaDBBqEl5vMF+XYES+u6d8bm
yJ3HVFadHbu69Pvlp6iiN7NflWIhLjK//1SLZjoAx1I619ISKACc7xr98JaTIvrIiFUA406e8tcF
mw3+jxuNhyM4slZOnsK9oFzzweZs+Ld8/g+nITG4A5JGL6foOft/zyJA1s5nufWDxxmA7URWUFP6
o3ct8ZOj+2EqJmdjARzC/ockxsevg01oqz3ZHWARDhcWg9CCjI8wKQojPmUfcG8RNJFVLkwKki8D
s5Zj2GtoQf+B46gcnIe7tivafhpiR37Y6Sr+vFCe/zsUpHEhecvCW43rw/72BqlPDpWm0P/38F75
V9bQN0f2zzL3IgvPcrIU3ldrWTW2HBjBC7q6ZOsZQGjs0FoMdLtN6k6n1E7buFhuT0moTBcsUAM5
rvaKkP4HtCOoeSoTdRTWo49mmj476zv1CuDqyr8KJUOI36ZAKXUp4m/LyzmyH8EoMQbUFdwQ836v
FZNj6PctHYW65YGDWyxcXftJcMADZC66Xs2sOdH7kxMa6XRg8ZDEwAkPtw5/iffXzIouhop+LvaU
KZPykWIBdxUj25//lz3HrO+C4+PYMgaam4bYhF61SDqk8toCQMyiqHQJP6KcQ41cw3Iyt4jz2RaY
JzD+c8tYLBq6v3i6UfRJOP1clXNAbNeuAxgGhY1o8laAA9Aet1OA+rMN3DyPDqpPGhq0fCVoyf4S
y/oT6gz89B3zIUAttWnJ3hucZ8xJR2XJiRhOBlEmYRWH+p5AwD9HtrS+hiSOtb8XmZtpOAe5UUDp
g06b2NaOukuaCIVDNbBDq2BBJcDT7OGD/DL0Ggy2ynrYVIUjv0QWpdScdE1lAoq8FFQMzS/OrwoF
mmyoXqYdY3fwwuVheX9DSs51qLc3vNrNbkFY77oDFMBV/h/3Cl+l3AvcpsVE2vjlGPW3PbJqABy5
vEN9we6kBc9B6PzDk+ERfIwuVKWYC2lPpyWTyMUITK1tkwpFi1MOAl0ft28M5gFmRcT70NlQ4Dvf
F9u3nTsiKwJLU41qhSLJyaLzRWw6jqQ37kH4FepCsW/Bp0sBh7QV2U5CFXo3uJ2glk4Y+pASlSNH
vM7h4f5GkBPtJlZpXsFylVvrczI4rEGA/HmLL37z6lhkEhy7W15q6mBPXwk1Fahv+qowDSOk81Fz
N4YMZ/j9WISpaY/E+TEG+xGI3LJsxe/K16UlcSF6c705KqtMaDYwk2iYQ1pl8KfmJIR5785LiAaT
HqczVimqBgpqCnneRC03ppD4bz1XssIpg5Sz6nwNd3RsKIMgtd6c5u2zYKvUeBqLK79jn60Dwwco
jANFznB426ZEXEvlXQpFbKrv74qvvY0wTlTlhnpnGFDWPgESHTmc5cc3aRZjtjcIXSVsR8QJP78C
bYI2TgF2KcRvrjzYUbzluFXwPPSWNIX2ACct+oZECzKh90WXHh3EUPAmcNoCmUGa7NMl2Irf1NOS
NQXTDpeJgBGLezqNZIEy1PhCfA6NvMxgcXIcMdSnMHg+o6LFmdz3Ae0ylcim0GVAP0VIlqOJirGF
fkdh90a4CFgvGEsPvPFEoqB4M23ZyvV7L8t8AYKPfO4WmS0zrPB4G2ae8KBTSogbTGJ3LxTsiFiC
n41laASb0PhsZph4PIHzp5J+9ATz/atEAfTnbaCR2C81mvkZlVRf70AqtS85KsGlN4ou3c3kEyPm
+vkmXqnjF77Xu3wqf1OWaWAx9LTHjsNhx/qDVHfNbFErOSBUcz9xx3UD1YO8SNUO3X7EDXXSxTTb
msCOMVqdC9qxHqdWDt5i5zoawQklaeU9EhiSxHBTiOLptP7t8A25vXkMUVmmNKOMjNAyzxEQAqo6
kNQbPeA29QcZPGbo4FfBIzdcsYbTfCqL5Qv7wkuwRm0i+1RAT+H1IxW+yYw4qxkPwzGIN5XEByyv
ouJ606qsMB5znMEYMRGwPzfKCXMjbesJ0m/PBnorj4wI9Cv6NxMT0Fv76HELRXz13IqPAeHl8RS4
dwOyp8wp3vwlxJwpO+PjcqH1Z4v6fiN3iv+cHR/UTU2dqVGqwEqF/YUjRH7V0v7Gla2As/j8kyxd
IfDBaYNPp3KdFIql/LyZGzWHjG0WioTkBcsfuAkxEPPynzi9y94/vW9Q8nAcQ7T+3kPhL0YeYYUr
OxEbZduQzW01LqulT1TyPfzVeU4gLinJtNmOT8GLLQ5DIDmYq0A7deyg2TSoyj/IKA7OLBealxXU
91djHlSzzjyNFRK1Vj5fkxElwYo2ZsQWX+Tw+NvBOM84z163LTe1vCRuTT7eBtGyTd+tnIzr5be4
jXhtXGC5JdVHp1pPo0befHPuQiV93ZV5jQSuCvt15uqsOzUAa/W5RKyYEcqfIetA4XmnPmP/G2cl
bS0n7n1Uw8JWtMI1fIw9iKrlFaNBrGWMEWAeZ71+Ft1ijAXHh2Qjjek/vi0RpylZT1Rp4TELr+aM
1abjeageVAjNNflDMuQlepylk2WbnLh1P02tbctijcBBf4CHM47tnflXYoemvjZ7zycr6jwtey/H
bfGhc0rydWkUAn5LQSLmUU0RqVcdDazhI7wRPkTMm+7xQdmOnUiyPuaDRaxu7GsT0dKnLXwB6X3k
A9dTSuKX6mG5Mfm7nRXrF7hTEJkB4rpRz6VpRifv8NFWbO6QDOUVHWoHTLdFt8tBFtsLFNKq5I0m
3DDKhmDOxXgYiytEIFa5xozwgrk6OA++MK7Q7ESxNajEurTb70e37H+4a49FVDYMMUHC3BtFejER
sp2hWKeEyNieKTmUNJKzWzBzQDCJA6ztWGFCo2e07kh8kDF/KSCU11HWrO4aJuPpVYdAYOr04sUT
bBnfKTl/1WbSvkuNAai094R+HB9uypneDvR0P+yVVC6Kp2bWU1Ejwidclb2MNnU62bXEJMNLvgTb
VkcNRyQNzBbgnAhQec4wJbj2FdN6aerKyGjA4+hKmKEE60tBp2L5RFXJPdRD1uLKx7YntNSTKOAq
MDdOvoM1LqlxSaX35L39PCos9tmrS7lHECEGnrJl5bPp6L4pYa78A+yE+6uT54/WgxmkvOqVBu2r
D0gkqztgAiHmKrWAqJuUgyxexJLxwt0uULQ94oQL3VgT7ADekEs5KxlOp2blSqBza2bLemR4kPD0
za2oEWKOKRtyq2NR3GV7Xe68bT/924qK2en+rWYeeTnAbUTBOA1BRHjEzpwrBdF0ou+Sup6B7uAG
KyWmY4DamhDEUz1JWcmZiPLlJCJdspUrURUUkjaj3kqGKFjqU/pqdfVZ2XRPH18DpRqt4Od9KJs9
tqN/Qw6up80kAK+blkr9QBwyqJM2+1GNlaDg/hR3LUR5tfsf2Gv+1qtoRVENYRX0wVXWgPlC5/Kf
QPdzzHiKi3trceSHV/AUyg5kQkefkVIwzBEORDf0BOSLhD7Ng/nzhZyeGQoEnKfQeQfFmoZ3YdQP
JFUjteYRxwgnYmoEXQ/UBc52eErVaYwuCnS3AmBwHqQNxDMhWNZri/e1jYdpIH0fFL+FcenmsBrh
gG7kgLrcC8MYQMg3BYB0fCSrReCzoWXOft1x9iEbq5ZWXyi9GxYhaqEWvTulZ1gXXyY9JBgL0Qhg
LFpyP/tMwcMHQqhSurENGbsPaN2aVjnhNGWxxtYIQ9DQvx1p0cojXSKIpTrUCbi9lodZs1B1ylWN
pns6UhysR0i8oRw0ZNfRAN0NgV87vhoTccgUl6Cookb8aVxt+xb5i0g0eFewKRU7Dsmt9yr2gEnn
j38Xk5jNljGcVcwGUOPXvKAArcPjhS1ysX4/DFJixG0UIidkXDl0h3RMbCguc2lIuNC2TrQFk9Yv
bMwlHgcE0pbzL+3CEkv7l25wJ/phPIcfe5Cb5ACGx+AA+RgVwUp3qSmtF5qjoa6YD6JczcMLeCBV
xf1EW3Z12TU83Zvb2VBv1lQNebgqIQWJDFBehy4yKQm3YeGN/aDeuoq5wQvJCB3QRkeq4Vlm/lGs
ZT7P4z7HXG4pP15BESLKeu4QBx3w77Zgf6l00JxzxQYlHRoekCsM2uIcLYxx9uCH174UaNKzfoZC
POUsuqf/1p/AGRoVoN3ccGP4YksFA/dCIXRQl0VkA2+oUzZpzRUWZAI6c0N/GwXcgGrqNFnG6HM2
Havp0OQ/zhczJwLj242W6xE1ZU2V93PFZ3Qo9hzac2M6AHlouQ3nXMmDbPghdjK8a9vchrEbp1u6
a2ExM4eSCJtVgwPgK2wEzt0utng3EiG/9rJBeKH2LCS03NRqbrs+KO5Yn2nltyB5GCDLzqIjxx3y
RMAselQ2Eaoo0htgS0YrCsy6y4TLmzMPQ9YMU1uo9sxwMRlak/fURC4rKrQtWVXUV1VYVvpVWLFL
jk2ob/+zhoHGSXJI+ZPL4h47J7MoO+h4g5/exG3XnDCnokUYOL8qX9W/wPAz56Sdp/TMqEk+b1KF
Bgt2UVGPAGN3TNLjgc547zgV7nGv9K+LUw/M0vGfYqJGB3UsVDKydtbkN2dfegpZHVAc1uBaNlbU
Dgvjr6a2pLw/LFjPpquSTf6N5vAn47FoR7IApb8L//ziVw0pQ4wEbvhcR8z/44PBbaOxkiYiPn2r
NwggHcPCzR5tYkvThMlAbYa0PSgOH50eaVVQdRqFRcM0Es1t0FaEw0zq8m9QqFdECFsfPwESLHka
S9Q1CrltCNlGMZOpcwBe2ywMso8lX4dEC5cIQpiwNazQ6ojr0LKeP/lduLJ9D/bNgeX/9K63/QgU
PTz3DjmweAcGmoLV+gcBqhs3kpqVvslbIzNnrhsRyrLTpJqRMAS1qHiEcHr+seJa2sszFdwNRHlF
bcjbVgeKzPaZPb2i72slMmBv41VMrnDQALmaUDTVQaPesPBXTS3bK6Vylr8yLB5AfaF/F5jM/dgW
Dy2Ildx2EjlSyKjUwNq6EYIv4NpvB9/9nUzEwzJTktmXW4EbN39DGl9H7tCTTIYSUgTkDUzEWsP5
NwDo7XabqrKHQg/JKDEg6/qmEBA2si+LYEJXjbx5B+0FK5dL1SGhqTwrf/fIH0MgbXz/4I3fBfg5
LY72DY9txLyBkfPGqiokQ1JMZVYy6IcAB1eqptQh6LtrccgPQPxCbVz85rKym6wxr1WoGgBW9Bv/
O0p2SVH/PPYocqf1nQAQg3HyxEI5HHpwA2ROcz1X1Dn3iimAvgqoUM49SDYWi8yHRzgIa9LmfG5v
DqA6q8pHUm/Y3OCeB3Ga7Xyzv6M91q9bzVFc5PhkPPfC39fQjrXG9EANsFc8rHzTwXfBaZWmrGAG
mvZZK+s+3q8URfhvKX1ffX+Pt+/OHgMuc0Oq70ohJTvmEsrEs6J2uw701552kVTXrsafr3T8ZWEP
wZjnpggH70XZQSEnIqCQ7hCdDYpMhYMB1VZftuRf13X1GCZakrIJIsVgamo1oUagXl3eKE8h7Ex8
0L/2cKCtUgrnprIg6xQvO0FbBzgXXGN1NhV+ItmyT/SMA25aOvLTZxvSSxgjOfjGmrf6jSh5Aw80
flpMV51KPXRsxJnFO4rWdSQMj279VddgzyH3EBvX2auqbkj3UEiID4wsRtqsLWSAv1LQcPi8/Rcx
EANMeQs1/6bu+tSstLpHHNfoMAcRydX+mJ8ZmyRr7hMypMeIpfC7m3ION1SmVI563BiRuYkA0PPj
FzmyGTCH0oWOsiVm0e0DJh4JofaSkyivgI3+uyhHe5vp4tAeyHBpRa6TZPCsAAe8EDvWBmW5Zg9f
mS4TwInJtp4UCeNFzjnso/jTO3iK0teSsq0icP4l3CNJHPP0rlnY8zfCrhSooug5IQSR1JNJb/M5
nKL6nlUu37trMTY6alyhPxXTrxKIjTmXL9aaS1bUe9WMpovTTgXtbFrCsXQU05x3Jlc1UBRfIcmz
eC0GL9tkgX40oXltZ5DqHXTgujcGwkQOjcKG+k0m5WOe5UF4WTQlcbas2tO3FOBoiqyyY4cQYr+b
WbQqENbHOXrbqCW5qgKuHws2yGXp+yExS2j9JBx0MbzKeEB0iakqq1FM0U5PaIDoatKDTJ7yyktf
nnVGmuImK/0OFK/u2QaBkdEpRC3zXLy6pR6r3kWRp11bovRKW0278YvH7lKLmCoPViyKuitUtLJ0
CWR8X/o0Q/6Ytu4LiunHoTA07L7aHfbNBea3JNUdL2NqZPtTxaCm0PlVv3KmLfmmmmgDPtoB+EHo
Id0Awljn0yt31uvyO+v95TONElucNKAKqiGcDe3r2LEpFKBsdcbwO5Pbt5l1Pw74br0dSVw2FehT
x27hQRsNkgfylV26fT1RquVy8SB1YwB+fsQwnUF5flhO/y4O2FC5/bmwmCHymd5dqEF0q5pm1W/U
qhfHJDX83a1ACUpQwnBytRg1UJz+0syyNEfE3OluD2Qcat1DD6WnLGqi7hSX1EhXA9TKFN82B40J
r9L0Fe3P3O5GYbHyq2sAW8kbCvL+657DKqXkh77FHvABpOAVACOtFWVfkNyd2ZkZw4MHyqH5pDNC
l190W/mnFKgDVBJ4h2FuRCXH4ZjlRKxH2dFI4bG8dLdCVm+cofdYnnmkYyKTK5zhjMy1jyDREEuC
fWQauvbMqp2YULoFRwQ2yFu0xK/FVTitN5jlVA9XEoQi6R0kmgYF5Q2sajmXZZzXTOKj/2nLsubq
LtHCPlf3YWPgMQyznpWY18vJSWhs0NuUVBLotqpMArMn7p7K2trHUp+ppYFtMJ7sZ9Q1L6yrx/rh
YtBQGR+k1i4NS2RFamlnGZ9+8DESJUXvXtG+yrpPQpmNZFpat4jW/ALEAz9sbfEtuht3qOxdm48S
SmbgdwTs5X08MGsdNvWQN8LPl+QTLQ18ctAa3IwZawkqEC1kF+diGqL5FNRg5Jm3MxKrgPs5Xnan
CYLow1iEHkB37DW7hyQapzGemlsXVLTbInWU8Xfzulrc8Jvz1mLJPFKy6HdCpwcGAyJ3khbosRY9
LYBzGXhzjh4Wx+snIMwnZOPwuXjIoyZS+rAnATgANz6nNWlBFWz3V6fss8NWcXGP6WhDjhvFbdyM
DNrQdJfz47uokW14invKdCxWc+hOVnfBxbA+hXcyZ/2xWMR6Rf8IVzBNLPr4P8ImjnYBOhtQ0Qgg
BPyo+hYzl6QM2DhRJEgIJOKUSIVyV+iloAitxi5awR4EeF5nnj0hJMBYcWE64SIfaz1KGHNHMqos
u6M36cw0GQ7/e4/cW0kj+bO99rHm6z9KRW4X/m3+8EOxqEgUiOZZ4kBk2w3qrmQanJsjqGNiersF
hohKIvnnzsCSl2MiCMBBkk4jCdbnb5tkcOpJGrVrRcjU/kuhhCtj5hYLknjk3FPQqcdLO5TnLpxm
u+K27L7OecmLuaVwdST/ezBj7B6fvL3rkmlcaQQnBRWQUQvrDoLKV5/GXCOrG4hsXeCoR6XiAYeK
jVL/dA5rEpudPVLjDsIBsOKmXY+02jz1Hq+vdefq4natl2xXV7L3roQPgtxZFlp1Y57PP4Q6vUjd
/1rIRSbAd9zLEV7gWaKkHEtylRfFcraAvnyuSrRegnqOsMQgrNL+OhX5JqECIcyVcLqdYB0zhMVo
Iw/kfwq/oEee6jorUtrAk/OHBNoxeeTUMwt5T2cQvra/FzdCgzi0DKlJz1I9aoaHZ5M/K6HiA/aH
9pOn5/ujVyCzYvfxPaXPZZScNuZIcX4Lhklu1MLj9s/El0EGDNYq7YZA4W99+j8NH5iUzHWFxPlC
WJn3GyyCPxi1hWTATVVNEJLxHAuPIsK3q894dovT2zlhWfnw/7hJLpjMdlFLQTbnc95id9xud421
3dEMeIZXwz+K03J3bJlNJEFp39iY186+xH5+6y0Oqyxq2Unc7UlXJwCuO+72SZ4bLltre3Ail0k0
XZz729nNCqf4xkvDkGEx5gBAdvDKj9xEglCBWAFC1oetAyt6NfJrtympMHb3PJwouclimWLOREZa
99+8dGHnR55skZ/fsCNqm8iRz4ZIVZgmfGqWnEONv7ImgWgR4UhLxgxYOB5NWkrx/psIAqowGfmn
3CUozIB3GKZmlF0c3HFCErxg2scRehKr9sWd1/TGStcyg/iuUAkAUvFXLYi8JwaxavsmySRsDaBw
NVgSGSegWaLkVtTg6HavcMXJHOhLGeKAtjacvxOefZJMxFTy+WwHAp+Ygw5hhcAE/8p0f7CSDAyN
ygErfMw4rkTF1HP8gtgjkVQV+BFcQhjeFT7C5apJ6EUwH1Yvmk1H6n0E0efoR5+2CHPsjM0RKQpx
EdnzcpyEOyEPs0uqIk8zWB6lCOJD2u7aIB+wuCu9OnBMtgMfkfcOQ1RYERexXcaIsAOuLIYF7JRR
97OiLMi9hkrYN9zpq0xi98FGyFHRpaEoe1y3WPKzUNi5uW4RclMiH3VBGs73QHczmRZMRbHlHQG9
xbnpFPsLbgKGWDc+tk/eMvVrWM3bzmH8CFwEHHVriwxBn9jiR903CMzHvNpQ7aHGoxdE4RUTybQ5
oMViQmr8E5riMbVT5Pb9w+JkPVvil5Bm3zR2YZL93fK0N+MvWWdN9lQr9tLcj8mncIAbh+PV8yof
zylNAAbZz9chUrSVbOevMuZJGFkxbYHO/NiDFjeP9GiMaZduws9I2Z13SxtNGoAkvgqa0IT2ZYhy
kTDvCWv1lsbxGkiivmCjGX6+br7WYXaEEIhuprc5SjmzOtbBFByiW7bcSizNHdNFTd06ah7ET3L5
S50+Ya0bWjd0w7BDeQDICSqPkSS7MXoyT2plZBlQxoU7JPaQ8qhX5ywM6M7B7w5zubK2/Ps7XyWL
0BkOTDy9dUpuB0sJlww07Fs61/1znj73waSbmib04ps9mez+ymu30fa0SVwK6SGYMETVYuzD86jl
sDdFG93QTGxNCpljNtffH5DB/BugpBhdQ+K0e4vuz3Ja8knEDYzh2+ngWiqplOtsg2kVB4Vk1TmR
wnocb+fSL2aH1UdklfKMfM9oPn9HZ1VsHuTS/eVIwynVBWlzxPVtBleJWMs8HFqG+4yZ1RW+oRjg
C3Lx166JQ64ySNd0OJT+rxcJqxuQbqJD+0Ml0YJt5obhQv+PtRo3/qSF98QulummBAnziJpo4yCU
wIz3A6GqJ/My6Bu/Z4PEd9von6Iy/mvue8nar4k3gx0qL/yjN0ykRE/OxBmTZNEbcTIcwEDEbEND
mZ79P0J27UmMdP9MMJcK0zt6cBGF9uyDwGS4i48x/TBooInQ/eSXYkkNrSGmJrHF8aASCy9RJ6V1
e51mLyXQOc2FV9k9gHKiTkeD6di/JTzVjsubqYhA/nQOmZ5SIEMnh/0Ly0Z+YD4qr76KR+8JJtOz
cC/+booO3uDbdI3hQPKqNlW6BITYEUf+cuXnArXqRMUh72FNzeh/dx6b9yh6U2Y30D7VzJJ/Fl3Y
EanNduXBOJzQchi7jm0C5SOYvuk6x5DXI0E/YGu+k6C1R6wcBHePK/+xAvwLHrXsyftonM3/sM7+
VNAIudh6b6lp/jkwGmQKrlDCjhu6OydQXbxZxnCRXGSZLlMG5epuaYufOnLk/1xIfC9Fb+wucJdn
ojepuHxdAchlQ/Dkkga7naWfUaQfG1JNiLJpQnJmT341FKtTX+ducoajr3HFlxz6bMBPa7qk9bla
NGRnyq+muevQssWBI7iOKDpmz70PTUcJXhWRVSGHQnnA4zAnqKkOfIVWxO88plHFxWhhTqgg72eP
r7lw8cPSMGQFIS1/SJtNyOCb8diLCmDQRekQJ6PoDTyznBNkn9aPdNWFCkwpFGddy51LXTOYNVL0
NFsCE9+EEap/6aymkeTluBmw/glKLbjAyXtj11jYGQO4yKSuzh6xpLUwUDDbTvxw93+qag2mNib1
P34KSn+6Q9KmoyPaiSkNM1P5hf4iulCg3MakupbEtbBd8SGn0d4KQoAZ+LoqPRWQRjETg5gKceIL
+pfJqBzL2OwVtUdwkos+Ac4RBTYYObKsEZDBvilWV0isPnFigG2MtUldEHy15NSEFxE2NigjZJxf
0aE4D12H+B25Jlb9oL/5xTAYQTbopeWsbVslvcXSj+TVzBV6fZ8nuLrZ8heTjkqBMDTyJWPnPzk0
aiX/MFAC2/+yAwhTCucB+CBMBTuF7iD0DZoeXcKVfSsXQc5LT/TlBlZ62XqyUNhDZvinMf4jhpyR
QD025SzLjP4z2L56uLYQLBg/IPaPSoF8Fd6eZ5To+yesWnuU91Us3oiQfVZlrg1Eq4Ey62B03nOZ
ulMMJTFHCmzVVFRJ3j5HDwf+eLVoTdN6n1F4Tk4dEySTLFg1tAI7KBm9aaFeWqxNajYCQh5fTQYf
0/S4MCZe2kwpQCBOg3LA/AgJsEtLmCYUiiNx0Qj8osvzyKeKnfGkLryQJIbKvXThkW8S0uBYa/Aw
HnhwOMmAlSMsy4kR97BB5IvMlqMAl2aaXccw/Y8l4QZlH3smlgJViBUsAsBw1NXjl9l0Zucs78sU
KukkwOjkp48mUyVCzjBCVkbxDu17dJQNzCOiEwMFRhkWOTbHDwhVNufQeWbtANbN5DMd6QshtaEu
U3elwbG0gwSN7M3cn3C7Bm5va+G0UkFSNGmlmtKV0IkpoKQz0LjdS2c7s/dTwLY/btMvsTWJrBNW
1nrWHZB8PRA8pbk2zW557TPndjJ7yDgsS+w33zRNyHElfD0wmHCOrFSCCOszbu0FLRpMRNzI8cC5
5XUqsk7CJHYAeYpO5yXziGpTKE/Mygd7OAOdPWRkrxqTLK3EDdtvmSKgzmsfQul/KjO4OnfkoFOQ
O0xPei2pyfQv8jxdc1CUlg7KXncygP8Y1G2UYuYQ+JuobH+RAMcQdofG5CWxHpZPTKh74PMwXaWK
B+ZaOFUL9KUz2q0oX54b7M81IQ3mISTSz889GrWbdB/QmbKCL22KLyNOLua7dlWd1me+ubtVXEj4
TyQPuK/mopNKffWgE6q/Meca+fdn7jyTUPO4laBkDiQsOsQJp4wE+xWylc3ESlXZ6Ti5RCgBHefg
lfKSoewQLYN3LEi/SKGY5FK1HNmpkC81KXcBktxQEQzX5OVyrmBcimiWtKpk/iJG0mWB9fE6LV5R
EZ71WV8pkMYf1jZOqShpQ+bdjd0MBJ9wtPpSRN36S6oUTz29ZddRILEZB3sVCcOfIRvz3DUrBXUb
KsaeXW2BaIid6DCqZ59f/HFp8uHuoj6lZJ7ffyBiQbwseuoqDVGGQM+u6JBswJyeRAJw9tAeC8QI
Dwujk9DtS84YQeP3Wk6vJQPX+unmS/wuKO+VFBO6RiRva1wJRm6kugs7zmNu/rW7csZmxs/YS4dn
KFeQ5BmFnxz/76qe6XWZ325NsNqylafBUC8YWG+nvWpi8cWK5yvKOU65RY1gGHjtsco6I3qp4Iwf
qRxsvDwLZHVKLWdndvIh0N9WKe39nPeiN91mHymYEFQKl7ugqtaHuEKxaau2To2R0S03IAIg0FgF
GJ97CLJV6KTmAGaFzI2tm8dzv8QQP1LrBuwXBor6m9+3CJtNuQGT4fWda+CcKlTXt0aI0wC0sBM8
37aAH/0nlL5Hnn5yOx9vp/Q9XnnKy58uzsNCj4Iej540goLlUNYKs+bmKhgHvB3Nc6fgcJ2Lqcea
VOJ7ijpNlp5W9YRcKch6CQnqpWfsQ/qOKRo6tPz5QqjTmrpO1nTLv68Yuoio4vyHFcTRqwhg+4F2
21XdvTVKzVnehrOIV6kr3TtZd6kCmZy6h+E36wfbC4gGNs7cdfnipLxqBhxZm+Y1wiX3ibF8KR7q
gg0z4PznmTrxThROotLlZI6HPPmjLrwTTMKN/vr0UzZjKm/77SIUXJPkuSW978ixZRiYov49YqIc
thaiTNfvKmMheoXl2JJh7w+NlpFa4vMevKdYUDJUnj0JSXHPK9G2uIj9RZaK3pGf9ooNChZx7NkJ
JIMxmd6mP9odL2k5c8kAgD2JIpcs107iViUQ4ntBYISmeGXpNcAz0GY8QjpzRkP/Sgl2/QEA6zwe
K+LU/D+yTVG3LcvR+xg01Gtw9VA+auVL0rFUOw3aX2pva1mJTMSD0pEnnJnmKyaJqkTztalTOGYW
1Vtjz4xEQZqKeiqM/y3slo2GCBrE685PwZ7RDpKhCwXxZxo+gtzPJu6NppwXxv6ZPdFVdavfgbf4
E2fp8zPDZzi7KvoPKMAXNl2y5CuKFWhMSa7DuQedgYRjBOYuXfO6HfYv8Vh1wdXqyGhVxayLEPIH
qHEujuefkMiv+mVbGL/sRvDkBFGzfpb/5egYmTN+Twye4nLYx0XC9tP73OJnPHtW5xdloBK2dGpV
anu9BMKZIvY9l2qHfJL8A2FLyoXDTSjLP2yccSIsXkq9B+ucG8xvv+qX6nxBYnleOb5HpirCEOnu
DoCVLQ752hUF1wUA4qDhLyyycrzaxz/fFNvUOQ5EV6yvQ8VAMDJQHL4wAIP09NUOEk6To1gs7gA2
OgVMuiZDPrWzXZ7we/h9z4+xP3jDaKwk+PitY4m8XheKKwUa5sWwbctfqixZAJGAL/POZLG2T4+v
If5mqB7naDBodv2JA3KgMtpVAM+hSNO1PZ3u9Kb6B43sJuJaY+JRA+5e9UQGUQiN5AhL3AT3KRIt
it2pACCCipgmZ1nenvQ57Uj9dCkgWXoTUa7bKhMj+igRb6BKV8cXm7Sd4m21PxNVcTrwUdpwor2Z
gPdrKJYUaZgl0KxCOi/42/91qAZXVtpvAwGwg0lTxuwIARRyVOX1+GSEBf9LKO6icE1N4FlLcoKi
fj3Z0Mmjez9UcpD10KmB8VQXMIrjXEgid3i0on8+O7wsys4m9Mg2ChtkgnL86ALbWSzbUfGBDJTs
QvRWM1oqOCyu0nj0Gh7hTlD10STc5J56fOAY5GH1UM8c8NayZwZbgzJ5yr12FddTWQ8BnzPnkoK+
7Fvsm05WZdtADNIbDUu5tonfuCe4TPt+s2mv2BXWN7IV0GDshCWTitlU9ZC8KSF6hMBvw2jdUYgm
659hFj8EJrRBJg0cq6SDsgCNHtGP2zDJIQk37ox7QJF/aaD7chEOBf+0DhKW8hciWagYTK2qWLLf
mfrh1dlhp8KSlBrNYlDIMJVGMD7+xCjyksXMrwZOfXsfDniSeRivE+sqhyDE+RFK2rjJErnZea53
0sVn0cdBKgehpE0736U+0CLQ3AiV98RyzMOhqSlUAbPkvL3vRPYF+R5bUdOrZ4gGBFhd84db5UaZ
l/ft7RYy4EjJlNAiUY0dmBlf2XBVyAtWX6oW0fGTzdDoXSqEhjnxDf1sX6N/KOhaKnZML+kQeEHJ
4PQVks3S/DjwYZS1xTfkf/c528rCiHAw1UlkAsbyCN7t+lVzimU2Kcirl6MS425131OxSaTOEG84
9esM2G/laMtjbnq+pVaWP5b2oWHgk7lqcmE1vDS+zPqjTG8TopmQXA1//njQ2TrFD4LT71/0Xsr+
uJJjVvKMYuvGHrHkT1fKyOTp5cwBOMYfgxuD5vLWQKujNccyrdGSe0e1VJLtExnwG9x746HA/Lau
KSsqR3E1j0W2g4fvh6DGU8Hpz8ek1K1MprYN8kMqXqnM9oDp0KRNSj9Jk8fk/bRhD73S16lq5c5M
DTdG0c+VyXMI8WHsyyY6inqELlkHOPQWHLg6uASi8b4q/EauPqhpT/7Az0BuogHK+gkmr/7OTqaU
OTo1sX/ArhuAcEseIRiA829Tv3P1oIkSMr5vbA284zwbT1IBLQ4OA4nGClEBaBv/uifaUdIPmXKQ
HoThaLl6zPHlH58yVU13PKeIwalumVZcRXl3USWQmJ2c1u4c89HTXdr+quQa8ATWX18l4iWb/40t
ezBTPslY1HS5Ou64+0OrG9TjAE2sWeZxrDZ1rYu0V7IPJa4tDVSkzEVdBXYPX0FmLdjq6Ay8zEoB
cODGLx2cg33J5FBZ2ChTswf5FppYhex2qWk6VMT9D6orSzMIzN+yJUJsSOOvS8BuMzrO8jPWMGMW
+J+mKXDFQGT+LGABATGu0NmzyIZRXS11lgzWk4i0O0c7++KGMbE9oYUEmhNWUaM9QzvepMHZUk9M
xb9S0M8YBBDBax8eCpENi680TcsfxfZrSP1Ou055/IXLqKSW77QKd6R/ABboxxTpfbh0sAHmwZtY
T88r+JNHexABsO2Qj2oFk5gGwtO0nyF5g60fq82iLqxQcbxUDqa8xUIQrIOHE28UwoxbjTssKHDS
lMfNURPy3a+7jE68YHp2XZBVeJstkCp7sMMRDFqRUOQB7xOO579B1AaSjaKZM0ddIqCWuxeHJQgm
cIz+4pJQ5LHuWaKgSJLkasJFRYRr5ctG6xHoFEq++Yy3XdNMNucdGReBRzFn2WBMIiJjFXIl/I5g
ISCoj/LaoHelaWXxtXffFtDvYuLl8QSWR6hXxdGp5eY6Nxf7E/CeIXil/x7ncOd1v9fFkZkQ0Dpw
g2tikzraBi0jTwLTEm9lXdoopCb6LtjEya77kZdW8yIQeCdVyoHT+vbIKmqF8KF5j+c8GBlUgmNm
KaydcMC2MxmFFmqzgsaxqDAq5StVwd944PnyF1u3NSv3nK1snxvLf+9Ywjf0Qb/TKN9RwLPqkpBC
3hamMQABWaYHU1U3ERrMb0oRrf0GK4MD+L/HID1dVLIaf5e/z6FdrG2RBe0YrY7ne9TliK0sEATo
ZXqNeDvcEz8Zh1FJqkfadaVaCfpBtYgbbQIQkxie7RGsWCcnDXd/WDZqZbUhq75+tE8f5dIsdMTg
t/gGh0FD1wVo347nwz+Je7X2GjIzdu7KHjX3EcXpFEqjRBnFdPP8ibr94MU593v+rcDElH2BYlX7
ZNzx4gaf6SCIO6BMwOdY9pxvd0Q3OnTI67CMjdNO/JSsYGVKBXe1fg0QP0apNmQhPiyT6cPj9W1q
FWdT0GFy829gnlwOU05ctoRXnZvEE6oImif/DhZMYc6FCTmPLx3iwEOoFpwD+8FzCLQhIOsFj+eV
+Z5U7Ad01/heira1i+vr9IbkLYEiGqrNznI75kKykfhrCZX0Mix6swjZgijY2Fzz5ttxFeEH2M3V
rlpvqTdfSUm4Ql3oyqg1wG96ie+V4QI4NQvl4/efVvwxPDe/M7KAIPjdpROAoujuAyo3mM/qDl9e
LOfQs79QP2OH7C8Wv9GKgo7/CNVYgB6D/yre/r8lgL7O76Icd4y+i6mIFjnQFbwcc3460v5Ut4nz
ckctWleOTI5rDdowN+SsFEvYc8xsBYZQY/v7oUJkZ8iPbiF6p1hVOiyEW+OX/oI8Oh8nRR8VnUds
5GcpEiO5zfBRWFYfS3szuoRG2IM0K9yMWeVB8RiI445Hm7KQ6Y0yXmIBOXyaI0YNHv2nfeWdpl5P
va6GdZhEqhBV7AAKS99HTE6jqk9ScRJp34BN8yaW27FWrt9K2KvkEOlHBKqaQNZ6CP1YtHZHmKKS
IHM8Iz53G7Z3mffsKbvus3/WWyLDnlsmQL2TAY8+i/2drK+xbcHJY/eimJX2criiUuNTYLpH/t+L
nQm1F7GoFPKJ2RivHY6/E36p7kWkd9ThwB/qahNZiovxAkUzu+36hVsrWzHebwPacG7GSnQ/fXf1
7YGO7jwWvjXNlpRd1p/9+iFkS3G52nURMgwg0Pr01P2wYJO+X19LIE8xT2CtJh7MOSE/yHZ0SdSU
92LQXe6q23TMyr9wY369a5Wdsr3dPLm2fGQQrfrL0vX85rNXf+iHDGHUnS4La/5GrwEg01VH1yna
tX5BkkDfg6MvJe5x8xdltpoR3JFSF4QcZ5VH0oM+Kb1PsreSdjOuuu1voCuc4GMcF8yRbCKh+TER
9Jp8g2H8fEnvvWd3fg1b1EOWymlCjuyzVxVExHs0psTDwrYvuIxgF3c4rDbFhk2eIOY//RGFay3I
3hd3g+isjBuMhTxHyVULlI6CY+Yy4K+Ntbvd9l0wW1IwDBka+/V0BGMEwHvmIUwSFgxhBN9aizVo
GaaYF2v9QS3C/0yT8MPVoped3OysHkUT6mwOBovmrJqhOT9pFdpkwNuTQqOc6y2AScsy6KyBI8eF
oB4xLU2Iapo8Hs0TtKhrWaQBCIFT4Jxd80Ew61t6ZnX/EoHCh0ELzCkOMyPwNnrFEHS72tO9LPQU
J3/qyTqXnp/A6a8M0MDbz8xOhRVkC5kkelf8kwVOvymgldan5nZf2VAcW2khdlyJTPgGSeVu5S0X
YCktk52BIohnIdTIJFlcFhLgVO9QGPwxT3Dc+5399QDq/jIWzD+nHkX25RosPXZaWsIR2oQ/7OBz
ckFmyZYf/tPTCLi/Qy/xFtPacth+OMofSBpn53kh/ZfNTesnpwZ+aI7vCiNHfhylahGFY6rZ5tui
6Mymscd2JJStICNPXze0P6wTp74QfbFOFo0t0ctUJeEmcAPdybZ92l6hAKWWFU8tlEkwbP1sPuq1
vEgfebF3Qt9zWWyMwBMaFNVrxiWByY3+lI8Ur4nGDv2KGoWd7ZApuB76GZkKyLeN4Kr0j0Zr9x9m
UfBjkkTSGtYd9zY5+hKUEJdmEOv6UF0ikKb0XO5/X/F81BiwBLtFB0xYn78wyRxVqt8jK5hCtr9w
Qdfc11lGKtAxRfULsEtEDyMipgwUvAI797gxm9QOlO5ITCxjyaNx1qWUWwbuFksgrfja8IJaecZp
TAdHQhCwKq2PmhHitrwHHv7n3fbStWlahvgqsslFPExhNeJVPJYMYfu7/lWLn3QjCOAXMMuWpz+7
jbAlfym3XZyiZ2r3MTVrPEE8jh0Xo3sBMA/8qV94CsXjTUQym/xTuYoFwe5rqrrRYO2SDfiKo1gQ
F0YMEDrl1X0nZBIFYHLYSnvFAFAsSinDS7OSZecGRjWC1d3s2910MqQiLUk0FZwM6phoTq6tvlKp
pFuk7gkdQbv0/5nl1GUSFBMm+pdvwUSncTK/Q6ucIq+7ZKMOMd3tbHwG4D+5Yk7nOaVesToZx+WO
tNeqaZsPteaASQaWw7JLWAcZihoMEPYe9BiX6VA5bEXZbvi7iIVUcngCCjbInM1ryLSIVlwYsAhu
2aIO3YAKepr6ruI3hH1AilHRsyjQm8ki2t42GUap1uysoP8tHU/0JrBC9r6csb9uEEi87DPGmcdw
8a1q1g1VoNt5Mg39/t+0dXDrFjC0SZrnM3g+URx0reIvYB6QWLbRj621znAOtAg33Z2wdDH6+tTr
0d43UOKoVErtptE8JQWQG2YTXrJGP9/WaodUd58vX2DebpJtRRAk5/iYpnXpwwceJjUEyUvCfJlq
4jw4TCWI13CWkcU63svTrq+ucMhMkAzV6Ajz8etkzMpyWXwiXo6RG/wPT3gwOJjH/9E2xPS+dP3H
+4D0fdkmKU569SLlJqx8xTDJfRWZV4ux0AhWNVLhb3bm42IRfZvHbudX/wRoyW7bFgHPFs1Ews6N
22GyCxT9V260AsNcYerLGiwvcfWTYuGNxb+lRUue/rez9BjeKw0j2eDUMYOQjEdX/tCarFwVucD0
wl4vA33Y6ukvCkOc+cceuA9j9tde+Qr1cY6HlcFWElZ9c7+ro9tjr/M+Q4DQl/ZMlwZwYlmZWFWu
dO2b5J8H1a6KMYJPHgaQOeHjh2j3aj8j2HsJgaqn5RcIjt+thi5IOOynqkEIV0Jf4eJLsMJLeYsJ
TUq4mu3QoBDNSWLGpCwaLcg7de3WiBWMU4xBTRU7afljQL5Nk71idr0WPjnCK2Zqs/J1nlwG7zh0
I0akky3LC1uY+tcuM3bPBc1hGbXeEnLVQAyqyairN8Q/q7FY1UoSWhdnZs4It+SyXmuPF6E6domA
/PrYO3ToE0icCz/laXh0KEXFAO9jY7pSzHjYTwXigbXjZJRW94En0dXoE8RowKRyO7AD19ORk2B5
u+T2YJf6IUJA8Kc8qyF0kYOf5u6FtG4GgwcITjeceJur9ygIBkxYE93QE+SBk9gwMMqLpI5pxmMR
zwN+W7YyVGwZ4koLmVxtkFYCPObqf+s3Tp71uaR+pkjuF/4oYLnMjoerpGcLxVtb2uuaXOnGTRHd
1CaH5fYO1pM4EIzyO0Gj40SwXnsuD/eVPzTipKk+kffPjFc0PaWMEQzt8AsQbfeKmYmeBONoLqTX
2nC8I1EOiHFT2mEXGM/ZOBvG2ENVQij4Ixf3vOtacwHHjzd7/4bp11P31wPHaQnkFHV868+NUa/J
ZtJc7gQ4CwWz1LSoKKLEdP6Zsmp8VKIEsTNIiRQv+OS5BS+3gQ4udyzlPjutOWVybAQsPoxGbcLp
QtjbmDqVZl/92xFTWKVqfAbCj/VgMf1K5WcOr2PJDIneo54zlUPRGdMvWYUJyKD8atmO5nGdiKuq
igQ3ObFmLZeqS7XmjcikZd4mmjxiA/k7qA0kZdzPyiXvtvaGJcIUIxWaM+oBGNI6ytahXefW8+Bg
Z7gi+MpuX0NcJa6cjA4CHLqVo5lKUi7X8a8r73eO0qyUng25b7pUv4/O8R72TlFCVcde5+rXyj8y
Qw6T9+08fLPsUexyEMPd5OvOE6Lwfee8Et8mbkFhC/8tbDH5qUwY7NFLPfbjaFg9pwic6Hr4p/LG
6qmVA6JmK38tjd1qdijOP1H2TAcjefrVhwnsy5FRu2A0HFmiz5c03s88CndYplIF/uBJyqppQRfL
oXQ0pxF2MmIEmOAyYN2H/KjE7J7rFwHBHOMjcmJ3CtK26MTDzt4tnMygR4yo1qHQrYY2R+HWqWyp
M7Z/1QrSUBuvGKI7ufXWXXfYeN5HmwEArnTn8IRTrSu9AhilVaakFZONRcq7uIuYddVH3u1M61ng
/UPtWB4Z/oifQzK6qvxUVK/82Rgdd64hiyKlF+b+Q0xkmlFh7Pv8qnCOukrdqyRF+SEcUTAh8HVs
wbfGaDE+bAyG2Wx2+TlyRRwq2oEuxVVIkq0J1Y6Bbtowdx1lQY9xYZh3x2MizYUrRX9RpwUZYSk/
ldczkUYmx+gyS5R7upkf7M75g7Cv1yzFCJ82x895EflrxPOxBRF98NiYKHMpw30Mm0BacBmIhjFK
XprPvj1lgpfMdNxzcNz0jVM/6cqZCkbQk+h+Rx2WCJ8HjnPl0CVkvTwZMgA0Uf9R1gmcUss7d0Cg
MJl8b9x2YsZrf82RUyy3sxb8d5g68brG9P6dbd4xJ7LJhVx9fToG52sBw9l1S1fj1ocX7eZrc52O
ApBmyxud2I1vYzRJkZLB6fC2cHqPkkE7pTKflZ5jq8rwklLm4iD6/H3LwyufsS/rTCgrk1S6dLS3
6LLF+IhyOKLO3h/qt91QmkCCGUpzfScmsmR5BIst+fy0oyZr0sLP5BNxQhKZXLif9uOYMARKEOg/
g5lLpN8jsArc/lRIPe7e+Tg23Rw9xV6N2lQlIvTGCpl4pmPt3zsGqDqxo2veW0x47ffFopkvuJxM
iDGX0sex522+DB+H51d7DJAEwUF5m08pASXJJHqluyLt6x17NDGLhHm026GducZ4wDnxUoP3UVB7
W1N7Gd0qBdRNL0gUoNrC4jyeK07dCq5RWVxl7FFn50G92HFn6ynLCC7RNg+oF9dIUTV3P49ffX31
Sx70p9vYe50YiWXfLh6t39Tyu2ratlRgotAoKQI0F6UEmMad0Q1SXd8sjAQnn/BCg+RBIEPriYZr
97gONFTQ2sXyEEU4hh+0cAKre6VzHzOUmlvY5OhmLoCm2M+CP6hHNq0e31HqOPOChlxUiPxLfNlV
qMA5kKFz7B5ahnJde/MC32l2CjwOLSREg7Kzo6pGhHkge29UKMYjYQJ98H3SXBb86V8xzdSwQShU
lX+bRAxhC25cJSLK+hvn9MTWwBdrWRHOgqzsw//ZSHaAkQdFgoNY8IV1hd5Kptob4omFx8/lY6NZ
91uEupSKYPePBKMKwvqRs3ky1iM6fwy+TBC0RS7Pm8DZiDirgOR8YqLh23lfs7SPBQWzB67PJi3T
4NFACMyyUvKf5mADHF5nIJjgmnSXfXbjOFGsejL97IbxYQvQlzbnNYPiQr3Vmps/TSsQlQ96xlZ1
MXIWiLmpFtMlAJJGWtLzUfoaky1iG2DQOLM61Khoj/fozoMAjvSWf3cN2ZrRKA3A22jV05cJ8/nG
nqzGnO7oYEr3gc2C6lKVFI1SiD2OraTTY6VQnppKJPqpXDo62UUHIIS+E6wkF4hFvUskTt1XTviQ
PJ/7biXzGme8WJ0hMcEbe6QBTg9NZubW8Dp7yknlrEk5j7EnkGxAMp0Oo8iRJOH/hnFITzUfg/Zg
Zmi2TSDjZNBklM/oUD2vUpyRSnQJGXv6E6DUS/eNkGqu/59mBTf2yD1+2Cu0q97BgouLcnJ4XEFv
02t5hX8Eb+FpCT9Lmi81j/zTDhcT/RmgdUpOc0rd/6FECGyCXK5ydao3BnMbM0g3HqUW+dmaFObA
b/5Vju0G86kjOaY9gEdPXrvbZ0TT4OXL/+ig+2CesgrXz2X5rHINlFQw0eZTwKYQ9OKBbtBynsMb
cisnc/LZpGlKF9vsb/8z5hJaXbTsyC0yvEt05cppK6SPYnn+MUFC+XTfGLqQiUQfuFxz62YCbzIh
AeFnz9OwfXVJz3IN7fl5WO8BUmyof7R1tK3PLVvjqw73/bAjTFsBVzLBN5Xd8kWhUIbI9fYm7cUz
Q8tfTHyZpsQqP20ZqSEtCquoq1MwytiZErc/QXlNuC2Tv46MTpa4noLVwR3Rb6oxz+3KCuU5XJbp
8Of/dWqVNi9frR7YV9UTFsgMZ46+yqTunBbpgrcYQWBVKjoru5GjQND5+Ch/ag7F+ezVsDnpUFNd
kgckp1hEx7XHuM5HZA3McVdDb6T/0RUq7Mipr+FAnCVO09McqcGtnAzCze2axwejqPlJT+B0EhkD
y390c/jpeCtF5CH3gr/koxYcXo9A+jge4CA8s/lQ2H1GG1d+B7OFf++GnJxNdqbgHhoicyu9Xhjx
cqN5pZ0ammUOG552hgMhceO7q46xxAetm3OmcdRZNSoL1fVSP9VQXBOqiq7eciHDKNHaO/GlhO1s
tDDNyTzlXnrHQWbW21wY1paMnvXAdMOr7EOIEoDEvdHA7N9mBUl9TNlyLviobw+2hOzyJbQxJ2dU
Kc3SY4PmXMljdIqzzKxpCSp3Pv+7QjBzBsMIm0CR8aOTeWNxajbPZ6s5LXH/Gfo4rgcmxNSJlXz/
dMVdBGfiLwK3BL518e/DjKDz+60INJcKWjtt5Bo7xBGriGZA5wOTfHVe3ZTx4QxzHpCSM2Bjjl4B
7EwK1OAXff785YmQH5glMNfzmR74TqtGG5baJv0SPxnzBgxiHhxle1YeCDyOAWFeAYrVFesluLb4
x7WOmrYDcv8rZ71Noe0Z8etSi8hHQ7bWtQ+RDUXOFFAOMrEKqeTIwOd/f2d59PhR2eN7eyVCPwh9
81T6RHWIzf/aGQcM1Fqj3lZA7qk1/1rC105ShbBkB8j/TlnOjTxOG77PAWq/G9s+RMi+OnkdlBZj
KHLAiyCVagKg0eQLcpl4xqiFkJhXzrNUR5kUkXaXbEdVZ+c2bjm5tf1ftk9opp61NOgSNH7mJCix
LfzarPag7rXxW3qTGC6KRnpoDbeK0+R8VxBwieeShWtJVEP6C2a4ejBeT5mYLIYW+Myfk0N8chGY
XME2zfR+78uVRgZW6iKiystYI0Fh+3RqA5ajcUjBpntFcs23+7JFiYU8OrlIuK0b+iWbydmNOIGW
Xu9KOdeCzagX728L0qGB9u5G76noPBRyNwTrs9DFzcohSpV1Gq7rof6NcjSwy2WFu2uA5YkPdJDS
gxWGxuHW3hSCYzeQ+JVg48kER+DXcAjcNx2VXELdumiGa5gyauoPBwzzJdOy8DTyDbLGO+dQ5Ptb
KPO7x/Sn2/vKoGnuNr6COW89t5S/xkK0/xciFxxEfm0mnA2SgxYy7NICF+4PbQXl7HYvxYQmbYOA
GBJ0b4qnjui6T2+jFuutnwVu4fR28CRaDx4fV1wEYsq/PD51QUMSMdWm1qmhGxa41GqjNARt2FPi
bxZnQaCjSND4vIYp/0C53ZJyrbL/a//6fJzDv0sU8TFqLfaJcyuWjA7AhsYc96ni9mPy+mGkAo6N
iaiIRNW9kx9xDdYrI36CbWUaT9PGPRqF/45FWVvmqDDQWQtqGu8QZiHznif0haF/mvXwoTMLZmW0
KpKpp2k+A/2VbMGMr3WhXAfdjWkFzpPoDji+H83Am83mtFo2ltsPYfIxxc1R+fjpkGU5Jg55RqlC
ptWD54V9vIWezXWZB/IkrHnZ8ieXYWbLOHc/RHWJvW3PaF1X0YlHZwbbwTQ1KVWd2uJJnXVqrdyX
gW3HyWYdvG5omq//7LssF3IDcvIoNOeZ5H2ucB1LC0s9VrK+MAno1/GzvOBAlza0MNbjDxxU3txZ
rJYd1d7FWqWdXlhqfBb+gQ2AJr3s3sBEQEbEchA4R1XSc94JzsCfq4vP7ZgCc4fosn1t93nA90fE
dMV+oCU/Efgqvgf71QyzrO+HKCpZ2c1BbbZjw+i3ThNARze6ZJvxAaJqnjlwLqFrxm+FJeBDvh9q
g6mUBdWhygW97VQ3u2eKVlzz6Y5dMKafqK0HxMK5mvfb2g0Gjse/myL9dxPRG2FihkRWC32LGqBw
s1F+XKwUAr092UghxfZVzq+fn4Lmc/rL+J/HnKO8nM1EWFrLpFw47B/4xoJVWdYpam4eXS8QchVM
9lS8WECDobkbHR1ft9aTkbFemghYoYNY1Gyq2yKJEbtw7VpqoJcC8XFtKVgK/ApsfqQlqD0jBtHv
vxeuiLAwPI1JxoiUplOEkCBSC3N4H2uF6h/r3QnKVBnr/K63stgBilfELSl8dmjRkNqvgiy2eRal
w7//1gc2K8b0YMU5ZfQIiB+Ln39Z/lXWzhTLL2NqhXNJfGgtECWeo7cEWD3OdzhGjlnmTWkt4GCd
3xvsR8IMx1j19rxDgUQWkDRIvWQHm1qxWxBzk0ZT8YyE0Dd6SgU/wiGvkI9im6Q7ygun/nqVN1bp
y2tZqKx+mk58+SxWK9Sd1+DY9uQLLkXgiNOqMxQtNof5rFJJaQoRjbrFYa+7KaGSlOuZ7I3eUqZu
pxJp2B6q8pIkwrFyw7opom3UZnn237euXShXtxej7bR1uwgqprFfMVaC9V+qb/pnQwF0OgjjMeSu
LxS9dNZfT0n7L0Ib0Q6uvbL3SCth18nIpGXvtSJkY3TvQlCcWQ5qFEgN+QRh64Li6f9RfAfYpuzF
semuFcGZZHfUoJEszVW0M7q6dYO+Wd4zw78wvr3cVzaTopQGT8pQCth/tgBVxVyjfdRsIN1+8ssO
4U+H/b+IinKhfsE3ZmM1ECDbPZNfw3aJsaMd4c/CnZOYngpHcY7fuTTBrALdL7J8kBSjaDGx8Zt0
iS1ZPxcfVFb2wmA/fqLHzrMeU1lyh7rhnQfrBlt4+0E6tHOwEHaT7laKZx8UUdWPshrvVDEb6idU
ijD4wun+apJZSzw9v7Q+s6Bqw9b8JeYYmu8YNJIXaEfCYD4/SsKMgZnrFx6ZtAnmQG7zQomcJK9w
ONo7J5q4Riqgukyt8yu2hesqz90S0zSIBKs/KLDBnomOR/gBUnSZzKr7WZqLhLrndJVBsP3kGuLV
REQFg39Sraemgr96CiuzDXQ3K/TaZTkX5cXtgwtIhI0qHiW/HpvNHf5VurB2KAwVF+XXB8UK3SaG
VObxQ/033zRa7VuVKO6ZSBPyuMnYjaEjhaJ6te0aBO0wzB9bekF5Zyyg+vivzz2VNf+hS8HoVrzp
5g9ZFaUneuvHJvsH/gsVNgSISwdNkJEgMFdW8V4J6JAVmihW+zG3ZyKJLzvMPTcq0eWqckN2HIOm
edVdjaJQk4LrIePyiG9+QhcfmoMgQ9XEASwQu9l0Bjm2/xQOUtNgPyR/M2EeR9Sjhuuo3jp0gajf
6LcH9Y8lH92NInEiU330Q0NH3auHilwCU2NQPXhM56sOrnJgPCpjPuM2WAb0u0I0phLHIfoBFv+7
vvGc08qQIYgvb6qGbhF6/Lp/XvOaVKFGVwn2illAODwYTshaNDvLBtgLEJ4s5UhPNm7kGJFxTOwZ
bLLVBnQy3t0huIXI+7A8b1FkernDIzpwP1v729PQ9fQNE5gGthyFip6SX8jAMz7ePhcj585zMU49
1mX6h1KwUy5dLLH1/mpVf9Wam5/8aTs4b1aru0QAt6ha4x95lSh9oocoQHKsKn09Ru7x2LuEF+Y9
gnEF6sTLtfjwDnMtfBzvBi2Y1tFyO3H+gYHanEy4OrRBDaeNBfpMAkxrOOK8qqDdvAIH41AUcExw
VA2CSTs9hwOsYGL98NpLPDd2Vp2tNfdXNCDsAyhVrsoMQ+eSwKJdQYrRC+LmeYGZuacgXukyH39I
veAFaG7C+nhG+tlavgXJRLLHwgCD+GUrp4TZahTBm3aWwUX3vgclLa7/1a9VSsa9IXyvaboURQEp
fsMBXRWkOOpJbUlWc9e1PzK4DPaFHx7EiLQDapEz4ic5XeXTs+7P3YK7HXEKSQXPysg0asrvgqGH
t2SWqsBO+p4yq8APCzmr6yHQfLFmN1ZWJGUTJgNL1ieV1L3D/WkxNaTuOIHkheITnVKp3YSAIjVR
amLKh3jPxbvY6HRYSD8SoNreIfUW6XBD8PNNeQcMev1g4FlS+rqQ6bXjSd83z1SMGJNK9im0QZ9A
TUhWKv4yD8WUtscAghUXO43+R5miEmHVQaZLaK7yj8eZ3O3dFi1//a9F/E7rVioLpdlKsy5CCqoa
U+hbr+sjgcMo/uGJblAObdmHOZiet5SXbiWCSZnJV677L/8Ye6kE1ta2uLCXUWhunMSyJBfaG1qJ
Mmpi6rKl0iNsugKx60P+PHLtygemnuFvq0DzzG+6LMzbHIdVXSmgHheWeblKp/yPDywrfChiKIX2
qjdX/4g7vivnxOHQcaIS+IhsP+2VHVfAoIuoaj98C/TGrSBl30Ymw2/n31R7nUsNgJW89qUHv47+
GJOKv1rr+T4Br7l2u99Nk3W3cXuzGx5CV/c6+CHCLK+Ug1xt3JOUscG0GSZghaAcBK557EUMY9tb
c1uWgbw7WJ3C6AXC2AI37KxnuO0JKrGh81ZA/j3rezRKywmkXoKqNDc9EKqn6OvCew9k5nyrFH70
wE4Ojn7FVgS5NpCOhfqnqoU3P0QoEVdG/mJMDlYXIsU9DV8L0cwma7muoemRHlj6Utd2oTYztXU2
H2LsJTtvWzT1ZS5h0pAxBRVBaAjfSRGb1jrP2Hx8esTlvQOfUi4xGFMrWjZcsuSHlCkCTbOebVuv
h3CQIXRNGZB/YilUu0Ox99vR0SfD0BDwlIw94Slwo3mvESxxTEb43ZXLbgibzSbQTMpL68QCLNya
+ILkbAwIk8QZBhT16jp/Lfzw1UUkNQ3e8lYilUEE55ETfOiI0ZI6fJ3rBl2NrdjQnBO46tlaiq59
cC3CyppIrwb/ERxHe6V6Agr/5+MGZR2sgli1QFN4g3wxOxRWh+mPxikcIdTUqvqq2h63Ew3CD7PZ
DX3iR+rNcM69+8xlPbgU5JZjeRtliHhKAHBjAcW4t6HjLLhFq4FWBirBSBPEhYbh6Ac9zLdzQlsh
76dD4d8cu/X2FSxKcz1n5iRVWfrPAjFYslXIp4J7qgluYEAR1teKLuk+ncj53t6sr7K84L8ksXKl
v6dKS3DT3YVCzjJAuKpRyfhjAq8EeGdfMJ+P7DAWeaXHei+e/cbFThz5JsuFoqbTLmsMHSqM7Q1g
NFre2cE78oAcWApwAV4DU+3e0D6qjA2vfBsXOEagFy88A6nA7JoozAJvhUTWdVfy8Il//Uju93Mm
MfjqqnTx7WlIeSyc3zFzgix50sKt3AAH9oobS4OBvnYXn/ywigOjL07hlUMb/ewdAW4izLDRqoG+
EDeL79eeT//jU2e2v2EtaCubHe/Y4AEvsCn4I9wxSIJLs+wkrYI8Tv9hWPGNvN8lN+WiTia/G8Tx
hHEfsQlfrGYOz6TXDMGTbvHeIZxZlDbpr/KJBwWR9uUG6Gwb4IdflcHYPfeNhiVsTubkrADaNpfW
7rFNUgS1UvTiPFi2rM+rpiCSS+5amIsMOBlNCF8HuL9q8ZGs8C8yGExW/da+Lgf7Px3ScAF9WD9s
Bm73vZ59QfGAX7xn0dCQJzdSyl0Ntz0XjFVmkTV9j1JXpYSrUmrlvr+YP7RS1+DZiTsEe8E1O6SL
JCqVUlNDGkZLDf09Nr3nNVgESr0x2XCnZbrisnC764DCl2V4QuMqeks3WWOQP5nqDYRBLHAyatSy
zb9nIRhqWxBzGtMEQumFPmtl7lKUCVRoxIU2vfER6ZakaUgSM/Yx/tGIOICtPfbwLj7NKde/seFK
T7VKlgWowFj0q+XT5sPWKJBFeDz0NbNxlkeR1yhbkrFLPShDa1oUs2TRibH/jQpJy7sU5oD3jIk9
fpx8kZRvwmLJh44B0iqYGImcvezR7++3kmAd3VpL0vHZFzCotvHjef9Fy3U/J2tvnIY5v/hSwNKB
TUEfu0qqZlefIrKEzmV2y2Mdz9W1hNYZdmeW4I4F0TWKlH4sCv2hXua/p9xe6gC1lSVwi5x9t0T4
p6c3klrGWetiIupDlAXFt82bA3r78vrBRIu6+skMcMcer3ozhtJH8ZC07sfVyYtZm5QkKT37D0v+
f4k/vW8WVUrsX9wkFyrGoqVs2Lo3oSOZ8L7Eynr0qqiIoYlAGwh9ZAVhYAHKoAs90GSJ4xxOMwYy
OUqAXFK3HHryHAYRqNhO04EAKXCw5rgzLdwMV8ie09JraueB+VmsfMQ8ifSfq6fobPMd2Yvvp9OK
eHUWdhni5tZaJvZRyCyLSpgHwHXQ/1b6k8hy34Yg5SbV30oULfOedfNQo3lz7NZhRj7FSQeBpGPF
ZEBdEYx2Kls13oHjw88mRf/K0Kk1ib9sKNLGNeqGTqswlTD6924teoDvDAU4ke2uhbjX2H/F9+xI
zYwc4I08ZU8rkDuvKYkIcE5zpEuO8KwvtAdcirktQiMLINAqEvB+Bt76/h4QFeOE5wqd6lZmripn
WZWWEAteqOV85D0YeTP+N9F68uaqm2s7M37dSDfTQ5434p8/qtf0Qwz8RGyJpCAvR6HDTl4rqVh0
d2h0SSWPISe7LhsnOfr8DyzqkTxda3x3H8DppQFLWnDukkW82WqyFIY9c2u/xcDBGzmB5euB049e
ppW/oPXhSb6sjDMhLkYYgikCwbvSELz9OCd+BA3ouimyC8qmcOy2j0vpXhwxSJItLoWf/x8//Y9Y
Cl3bncq7hZAdTHB8F8qbeNLQXq+FIAehgbU6orQoPN2ju2DLw7Ehu9S93QaK/bnX1qX+/ek4OB4z
Iv2OqGkmTnATkekzRRs1GknohMCw3tmqlCRqP+SNDw7gv5GIixWwUJcRJtn2k7TS8f7EpoN0qDv5
ZcJx0KXYS5amjuzZpi28urTzzrsl2e4VhI1AAOLkxh7kYWhII8qOymySzvgeJX9RnvZd0rmtRajF
P6J1lz+IxpwYoepnf/G8dR7xcNSwhVUhZIcjJ3ZXmSBmhNu9J7d2RGHoeMNY22b/qEeH6UOaVo6+
j6yzczUBzbuh9VQkDPFr+3AdX8YB1UGAsD5WMomZYt23BFCRgf1/nRe9emRdc+2wKEdEF4fmGNPB
/PNkJD7EGwrftKbJCXpJsYl0tEMedL6cvyPefRf+ynKN1w6xQmm66D80QLiQTC+8IuxIjrliWZT0
ChYKVdrAnvNPVV8aEKYCr22zRml/G+mQ3rUPdOWybAunn46GU8euczxoDUthqLcKaNBFw33Pljx4
ylH795zLWYm+QgbifVYT4wrFdyDNX2KhJXGH/GOawLYdmY1B505LrlGgThpD9TWJo3QkFKbHMhjm
OunN0q8/MlBL//Y2yw16XVaPexm87c87oFot2qS1FWrQ3bwW49QHGnnVlYmFXqE95W502QXG6Cjm
M2kqsEuBslWgUB+bcxlBt8Dps3ZJ7x7lQLMSy7ToXLuIYXq9Tc+PRu3oVYWCIzmu0XWlVeO/dBM8
XLbovZQzxDyWKk4zcMzRjjHq7Y7q0wj/16muX2rP4xy99yXZe7vIyKHC1shUSxCOtwHuAhChIGg1
YzEv7jZP0p8tYSYQk+P5hcmviTs8gkNeZ3WB1pVJfVvkc0Y465+w2ku7oaF1OFSttyy7ECUYDRMQ
o0cT+gPjVM90U+j/4jVEkC9jtEaaBLx5HeakonOYUqAvs45W55UlwXtTm6+QM4BmeEOtnMCHjIHN
zeuuHe26n08rHguyFBGjDe2/BvAKKNY+FRmYOC3Jlx2mGsgjXbYHIVwKkNSUX1FR+6nqR8V6mYQ1
/+m4fgXYa/IHrHTddJTjubgXsuX7OnfrU0OYOt6W7oxdql77rKj/OW6nb94J5XGDDx4FR5mcAiVi
fiwDs+hlRgQUWdsSdCgH143TXlPSKXLL2Vm8PD4kiyOWt45AvLNSRxH/i/hl9lT/nOX3/DVLSBPZ
JGfptT7JCnLzF5sqXldE1A1i4OPwLsUY04u4uG5/9Zx3ZQ5DpLBtmHEGe42xRSVPMRQlG8W/AEVj
373pMJ2IFRjbIJhzL/IAc6Z+3MREOymiJ+MjanNPcDXpCGfGNOhUlHGHosrv9pONONswo9wkwLuW
GOvEb1DbW9XVlCukGGT7WkF4OYox7TXYgR7wjyL68pgLdAODQt1zP2MwxbNTj8zc9wm+OVlkxuYl
tbFFcyUwxTz6wm885G3yMnn8/eDXvUor3o6RIxJdqSGsD4+zmN51BALs/3YCPYo/yZRrX71WkQTw
0//AaAG8HZN1nZsXgjV9W8pt5pRa3hpDSJ31KfaKzqsbdoA7AcZ8mOBOsqIYoTOM7KaI3dWFumgn
LznPpvJ5qrtXT51uqjnvKYpAGp+PAHHOP8zj2wR/aMjQSZrLUsrGClRy4cHgyglYhOCpaT3D3eT9
WSoVc4MtJ8a99m2MVKa+QiGDuj2YonarLLOTkFViPlrZr8tJAGB1Rbvb59o0P7L/nMGcpD+AR1DT
5vc/lw0iV07WgbBdWH5ES4BKxGK1Ps6guAeMjcz6pRkW6Se/P5kqNc8nE7G5ucCAkT8Fr8R69w2X
A+v54KLbFN0P5sgJ8sN30bl23q376pZk/zXZjrrqlKJbsVJt+TcYIq9IHlFITwFzQ07UG9xDW8VB
Ijzn9YbiA/YtQuPqEQ8y19S88RoFXiFCiEmFBYqgTaR6Jp9VV14zLejUPwmmM24rrlgd1JtIzed1
C1gKfct5g7Dtx6QKYOjrYwjNlU1Hnm702eaTE2cRyQ8RCaJDegNFBjcpdb8XsYNq4NNYFoCfKlab
rypFYzleriFPB5kmbzT4ywFDtDdlyWnA9UoDI+6eZepf/Tz9cAZSdlRWBpkxHj9A3s4qb2VvSnH5
vQV6SGJMzqGKWM6jrSAUQ7LKxfWfHqudpBv8/PgbouZrbN4yh/tLjgl9NWVWfPFdI7XpgHX7s2zT
Am+jyMuGzksEC9ddYmvDeW+LxZoWHIL4N1ZF+dzZoBqHN3SD5TDzu1E2YlaoFdwED9TliYgAinkH
f/K+ZTLP6rbEuEmKTQUzdwpWj3K2oYDG0ZdxRbtYgjzicw62xOI5NAhpgYyE0INuNwB25B95fCkS
St3jxQr2OxbksoWc5JaHqzZ5B1G+hjjB0vM3+TIhKl5Gxb400fWfC1X2WzTloWl1StgQXASZ24aQ
ktHd+PVttUmu2cZEFnqbNFSk9ukECOWDPMrKo5B/PmvnpVCsXKeP4uZCyxhPEkBIvkyPlcbKA1XO
nNk2QXJdTNt89HsUa0LKl0OpOsxAuZDrTzd53Dag/2+P8qCaF8R9wkoA/1vmAEcqzW7r3dUHSckf
4qk1GFrLI0yduNbtOlty5AdyA9SSDO4IeWSHRmUrZAoSTfDM5Sgpv2krSlq8adOUIvF/DHVEGGxg
2LiFeXVfw8ii2ml7a/NVXt4pq9NjiMsEq3zK+hXNcdjG+QlSHJtFUon+CxOv1ixTRacPQwrlT5FJ
IPngaITrWgx2DT6HRjFcnBI75+PW5l6IoQg9Ewk+gt70+0HVodSm5H3n0NR6bXGfrisg353wIu7m
GfZ7SzyQPVNOHVYNbfYEtfdKEUq7ORDbhy1cmOnXAHcznh71V2YU0am48Es0r7d74ea0l8v9CyCB
JCvX4PElY3HJUZWqqzsoYwTJ/VG++zjwEvbzKNFrRQa/rJ9bUpH6ZiJP75LV6F39MxFyzNRHLG3I
V//EJDDwrZpUPBDVKyUmCYUDT9VorQqvJOdaYhjw4lf4QSGKoTdJ9rEgR5Y+iaJ3IyRoFYYafEEO
1XFUWt9cYufbFLzgsIjpt9w8LajO7mflC96lCFnz+qfTfzF6Ce++bvmU0FVuk+w/b6hyM3Tchvav
rGD57dQlglIerOngdfxJ5C9xeYd/Npf+2p1GAVU+GZ7TK+bSzZeb+ZfTsxC9yE9CnVaeKayVBhFI
RqTzz8VJtJMX6u4KCECGRyxxV6uv74+l9xdXAEs1ceFyLWuhtzibGsO9qaRDRahC/Imi/vcxOrgO
xQejQvvaPk8CX1s6JX18mBtUTI67dMSG+bE4UhL63UowWcADj88l27lAkSmxfCAclsRCCoOPo3AQ
uYiklNYf//OiHTGyOGTm6NpbabWRlYlVVq6MhlzeiYXURzSNRWBwN3ymNJdFsTOkGcleU9ndw6fa
RWo2kc73YI5peNfRdR7Xs1/YvQlxGpbBnUlExmTLErfz6etf/+hGxNsDJ8R7mlRTrypfn8JiBpuQ
wfFxgPZvDB4nGy7xb2oiFWv3u5gV2Dqh14Nz9vRnsxVTbkApLjPKo/Kgjpu5j2unuibMuY/qyP1c
XaZqAIcBzpEsuBXGpWKgvuuJzw2Yf0pKvrvoDrbzo8ZC/hNunLpdu5vZoy0a8mjzpUwKt7yHd1+m
vVnx+Tsh0gJZS3Blv11hQjYIx/hUpIQvynrEQB3u4vp6SMYXek3FWAjjuJRb2IkV/V74vAMu62oF
kH1CeARxyuDdwGHcztBKjSTNBQmpYvwDmZEL1feYHUy6fYOSdih+8/5Iep99vjXhOiUxY+r7682I
kmoYs+XasbFClCee0b7Cb2NnVTMyBtU+IZSH+mRm7XZvUpQeeyTIwBfjMICuOFCkcpWNHuF846Ik
B+zZ1NQMPwKttBDOtuP7ysSbDKNJrHzjm40vsEF7ISOWyVa9xdw0b/ruhdtpQ/ZWotFmow2jOyVq
WOtiSWRV38m/61at+2vkV0M3CX/sH3u4dh4QduFOB9BfFxTrhOWGwHXZgboAcRW2P71GyLISu5lX
JeLBHNtHyyToDcyPAniIaHOhZShETLwt0HPR701wqjsMbhK8K2oo7Gi0lSffDcpL7FjOq3Mbno0J
5u5vZHJTRG3OnBz0/Y2KmAWk18aiJmZVgFLX9DPaXVVDxvAjZLfs3V3MUuEFM/ANoi8VVLOp1VqN
mATCnm+h9kve26VmrT1lMFtUnzQV3NqavL0udD2CGqcoRb51X3fYmFb7SoNZqGt8pMqwWfXrm+Ee
+a/NV4z7v9wk+gGvAzQ27i83azRbS0xgNoBwIgwY/pxViUX0Nn2fKcLSSHsgSwyhSBTAhpH7dVGf
+8fVKZjath4gjQJnqcl1wAaGgbl6Cj2tJT9SUOEtckBp1QHNmCB5BYCWujeIEYunyDfpYet62ESq
AC89bWFMT/KlyzXd7quwGGsBsq6D4WO5yqfzk1spAwtUNGE5tru3iMEJQKiahaOhdulaxGqVFGC+
Us2rvm9ToRNGDKqYlLdIyH93eYHrZCKuskhozuTbPxjM1p8Nqn6Y4iZCo3jxaIQpUdFNmVgfMfZU
zHf0aNAbF8/uRH9XbmVCBlTc2oGTIDPw9EMOOe2DZJ7z4k4HXoO/Dxy8k2zKvdNjOxxc1Y2+/whX
Xtveh5XO4kUdL/ehze4TvkrOPY0LKnYL3wOmRHAfBT4kjKP7dIvntq/c6nVwSVYVQgnuXFeKdR5w
h1CBRCQd/r6vGehN3lcMcpwSqu4davbPWEuMp1RP8jlDVAtX9gaDJaWXeT9oqPF01qVZxDTDQb+G
GR4+2VqG8LUxu346KU3OYFl41ufxzrRDp33JFMchxzynYYqI2oe2RDFVK1aaHuazJRmggiCFeT+V
FqF17Ui+DVUwCFJ6bhRCgnvky0uQ+Bqi052x9Os/jJefXY0RADmq5noTUrQZzvvrC5bD1Kqa0VhB
5t4ur18YkvU7D8sVjUmaJicKy6fCMUvIN4EyndZhmoje1DWhaS/GO8NyqecOxn4wG9SJ4djDx18I
CAFcBgqVlVKE9ORE5m1jxEA9IdK02fiHPSMWMDuTsNVyLG8VOecJBZU4mmh7jmdtHDuS1OnokxLX
azRwjcv+lb6EY4D4lRlXZ/WRiRrMSKXYmB7iW0jYHFvV+cPwIXOTom9RrZHW67FTz3nw36VbwvF+
4cU5Aa8P5BUNTI9TfOEAY9/8QZAXoLE3vReQh7gf/z5cPrmD3E/iY3yaWrFqWe/TlHI2UlBoUXDF
Knnj5IaCeP8SqgOn1L9P4BhvpDzWX3CmcBZC3hbMTZQTSyhOSVQkRWPxntydbLSfxtDj7gWm6TP1
+1EKQnb3s7/lOL2qZfLbemIZYzfJlM7gssWtBaD05vqyeuc6UJff9JDeuU2qgM6f0IpN1tQHJcWC
jsKe8P3FXjyr+FsqUSWIitBxbfseewHuVDPWBVSrwzUD8gwHamDDOyxGJzqx+nHbvU0gI5dVYAqA
lpSaBiu4tLAbZTUGZHL3XbbEHgY0clbJANtUcmydxTfQXpIqvSDwK7+tRZy3/fDvjXWs+bhVprEK
ivQbX2nD9TBjufsApbqVKpraexwSGtnj1b09drt0Sht5cyHuAPlkUQxpbPGym6qjL0CM+zKLG8oy
nCPj9PzgUVaKFRpUGHlm8tWfUo2ARdNA2hxuJMQ/dwSjUk8fpjg7t2vFIg7GXj3txqqbHlBnoeZF
M7d41ve/93KbHCfYLqiKp1b3yTuCkVNkJxAaJuNwMcwqDNGNOpnGgn7jTlkRa8DY9QhGy8SVAx4O
/cRGBVENUJvSTiHOZ0qMXyQ1QW80fuAtkGruwNZMscYTQucWY4zvAbNr0PpQU+D6eF9EMWEcgPUs
54sadI9hgDoafzady9/5YtKZ019pYc5hnZsYmYU+DJiEFG08SOSyBzhlj1fOsl/wB08F7bp/ctlp
Q6aNDB8zMNUgxyo1SezuKai0Ck0i9lR79gB471ESGm0On9Vc3CLfLZURHcIe2IdbepSPACaI4BRy
LFQYzDZBeXnH+1ZaVtiFRlhMKWyhRO92qSDe65Rn1rCN+a+czoK+PVjF83UXZcWx3lCWECAXvk9Y
i70stv8O8rfeZyVUYSY50gF4ot3120SNUHOS+L5+FlHi4JAJbsGk67FUw+A+2WdtFY1aycuMAbRa
RyauVht3LeedmD9QRPqIKv7DZsozpzATzLKZZndL5CagV2pyq+xigrXzNEjmVvRj9MCB3d5l+uld
IzIJi7bE91b5LriIr1vDIcFejLBWduAQrvwYIU3ABsJ+VxmGB6MRVmsZ2PmEyHXwfPD+vzuWAuol
eSgHFV9bSPa/gxeX3aCI+o2aJ0vnMfStUim9wDwIrwCLyX5bzDBoH6CJG8gcUD27J4+evkHdZJI9
dp5sw8jaVozrG8o7iHVnLd1VTJp4rUO4gwT2sR/DlUZc1DFRfhf5ZKO9h4d2tIO7KZCZU5LCn7P6
lAlDsVf2JxXru7BZSnxTqHWUiQupS1ZAtYi4FSxv3B6/rLo9dBASsgIvvXNukCYRi1RTaSCgxgpn
oahXrnYE+a14SOVL1DFLI0FqIx7kX7Pc1ctRIcFp3XyWRScqMSdVkq0/+pMKevQFUzON7lZ4wwu5
a4Z6+Q3U5JAYbAlXHkU2YgQWRgoREhj8TRlQTxud5eVqiszEYvHG9Bh08OULjRXi0dFSs18REayv
09aji+OqtGD+AHUBEBlUB98xZmUkIGQqM5N7tESEkzWcj26torX2KtD9asgWklONL0pRI4eYnOgb
opkDifHa26i54MswBdMPgoxwxPkYEN7/1zbnIWyWdwi+FIKYCVnszLFJ/ptjvXmV5DO+YPHEu+pl
R9JYBjxJQ7fz7C+6WPj5gwjolahRSFYz8rdJmcdd0ywJW1BBUoPHlsMZHhqcXFmiqfySM77V70ZJ
YwIHhBsSiT6+N3YOgNrR+esC5mJtRSpV2xVtJIZ+zHZ6/WYUSSO4bBF2ejTHRzrrroRPDJvGJn6Q
9OgQsgLHEwxRThE0Lskeg5NMya9SOP3gxHGSpy/GN8IyAr1KOO9b9ryzqrCoF93ityiwej18EEZV
16WNMcvApHRWM3Gqr9g533EZ4Wjc6pMgk3JqzhnTaQiigKjm+Os9Q9spv904f/DihP+RObKMMvtp
QAr+jHOYLJYwbB+G9Uxn2EbTBlijKCrRhqb0v2kB3YaqqxBwx9j2YcoTW5dy6lT5lMymvUWRzJiR
yWntuRk3WaPfZkRwTHKA/8+NkO3jT48/6OneOHrgSKQscb25CYO77iQ+D8Pee/RkuNMKlkyg7gkh
2n96JnyU4+rwEzuG+OC/bO2YE1mH2Na+YiPcDGvjwsglDqzf27vpAOU+d7R3rNqOuluyOraTf+GN
NAV642XgIhrgwNhNfMVPI1LIp4T+ThVIM2F0uA8keFMB1lZWz2rG5iT37PeEKvzPPyL/M7h9HR2+
IawqILu/JsZylMGz28ENXtG7drlwt3ohJhncdZq8SUT+EeCnsWzXLzW/r5HSHe69UW9dhBObiuWN
UADOO9Um1FzISOEHsJZcvhVqVKTblpzSqT0u81SWxYy5+YqwHKrdGTyTOBqejyHK053Aufwn/O5m
JbRA5/UxXNa/aYKGYyolLmLNUDS32JQNeqN09QrZAZZrGqVxIp1Q9A6Lxqin2fOoCa/srj87OfgO
hRL9HDpvS4H6rcmEDDInVCWvaNYfXULA9DjDsu185q5IMars0gtyh8tLtuPTOKHH1g1D41S5VAJp
G7Zo3QQ3Feb7md1Zo3CYlQZctNg4Nh5dZBGhLIGLGypIsfS91o9YzVySsOGiIy764xV2897L4HD4
StvGNkdoRk4XkEJ9r8xN6ztS0oAshzTZja2dU+0hX5aGSP+AbL6HHo1k2FlHuncLbglgnzIevW01
iykAJ2Bg5YtIpfhHY8JjgvMKxo4c5/EVVUdXVZ9VwfbIgMFf/88xf5SxlxvpRiwAxhMDfw+o6KJ0
mizFwnaHcbuYllx5MPeN2/6JDbp2tHj3wbfgQw9EhVsAQD/h16CaAxMy9+9Th2TxYh0Uigut4hv8
u8inQweJIcQWLxdCO8fWjkLNqR/0RvnGEnyc7MVnv8SsAKmOY2xlkYIcu5xV9mxobudDPzZ4MUQL
AeTn7/vFhLdWmo4wUqjuDP/5R+XutuRHzBTgOWCmaS0Jdvc8PxGY+GlRkAc2BCMPxdNaxBkW+6I8
LPcO2onPDxoVrVmb38E0D36RExwSDB8DZC7dRdQJYk2wCp1kA7PaaX5gdTukSRS0qT00NPo+1h1k
L9xIWeewXWQoCgAlmibXIL1qOiA0KZOQjH0INats+3saLiaMA1l2QDTX51VouogaqOcLAAtxZ1fH
9kyySl0tJ9ydfxkapT4uU9Z5Sp63d+HYIFo5zpGNb/g4neNf+izif5yJ5ReAQdVbQ8hxFMEH4JnZ
y3ZPOrAkKmC7pUVTU/2eWUt87dlv2MiHWoFGdiUMn50j3wD6sAP++bzkQXHHoQHpp/gQQAykCJxt
44kpJk8q+CwXcZD2Stk9JoHf5w8aGyQ02ZGcSHdWQTW4Qc5lDYIQj/ZP275Kb8ZtAFimGwegZQoA
gFh1l4YjDXRrdy1vT70JFSfwJuKq7SCQLvoHek7GZkc0cPsSYn985LOfUI0Mmo9+1qSqIfoYh+Nj
HFap86ngOMBtim7ux6XzfjmIgNC5NaiTflR+app6TRvWtRnAazln37tl3ljUsvO0zboh6VnGz3gF
wY6kzVIzuee7aoyoBckhzHbDXDF4x/T7MxfqWuzsCpipjXLwXvGcwDUB61Q6/7AyHT/9GzuPP5LM
Gdl7QOX6Uak4dytPfStjEi0jy/HI+zm9QwD4Q+ZmIgRhewgPTQQp21I5oOUI4Vx6peORVk+3Z96n
b22GqolONrNOXgarhg3qGzUhgiHo2QIaxU3KT268k3Ax05gCQGcCvEJA4QHeFMmhbi4vonlmSXU+
lZ+dHjudifq3kMmayuu0KJoA/YHAjcpRivQVoMxesRiyH9P5yzu0aPUJxUtPZT/LNzTzMrcPxoqA
wP2Oz7oENVhihBKX/tPAOd6nrlOWDMLhQEcOh7Aq1XsuJBEu6I+irAJAk32i++NbxmlCGRGsbtF2
V8U8iaaOvhNgc2sB3TLaxdXJS9BiSQSHx0fNOBe7Al0SdvyQYIlIJ3aXyFnz9gqN37jDNvA2y6vm
/FXj44vneNp5FTzIOzfCbBqCVXbH/M8SlkkjCeVfMixE9IOndD7LA74na5d9NzNoANNkEbJFSfjt
ZWvlscinqa35ceZzE3wyCyk+25x9L4pATrhwOCXVYQVYlJL8U1Cc5eoEoyUZxadjHX+ObQ5Wbfic
bqQQ8dVZwk1Hsdmv7o9Gm+cPdV+fZYYRMuGqR3n/k5hmtWnxwkUW6BNgseMmBqFe2lHiA3Bw/4In
9DjJ3vlIxZ9HfX4W+H/dnllKfB7Vfbd3kywuPQs5wje6mTJuO6I3HJHTaGq9zSz3n8HQd8vOieTp
OoWIegsGUWFM1/6t2Aoiqd3NoboDspc5Ugmo0X54c/G7wgJ3x0tdOMAWlQ3K6wkS5F0R5nukgfQn
Ge/Oj/gPcNfaRkgOKzAUjdzKzfuNg5uRO/I4ePBnzZ+Pg0Mjg09Lls9G9LOZm1F0SPu92dwqFtpG
awB97NPdtF4K4GTdeioYWO9Fm14EDXU/UcDTD0HkxaNpqPf3inM04Z7goHHRBLa30ALjZuU2gKHM
hEFKhtQA1KHrGnz0My92nJiEni7JMXM63/s/bka1bOtZ4mpk7hEVa8vgQclUO7ZNZihrmwXo+TfC
ymcCMHP15yPZLPnzXjxrDTpttydedIqMOHhZhSWgThlBPV57PhYPT2DUwIMl7jddUI7TpIhcfIMV
9xSscCdgHiLG1r2aiCfsw+tohxq4XxHnWtUjgxITczRy5azgBsx7znBUDgnkTFv+kwL66g8jTkwL
WXe2UlVfv/oGUVPoMGHnxe9RapSxcmDGuR1uGPPEAJhsgDkCq++mUG47ub7SO8ABoqHK/hynD4ZY
Vk/w2m5X6zqokAyccb4jpAEtwHqCZF0uBmpKPorozaSBOvMxUOpJ6yKOkbumToXbN5xu6flBU/8c
H4PSNn91RrRuwRXeks9CCCJqiDWeITtnaRTBi5eyLchuf59uYcjp/sRmupF7+6J1TrclVJb9YqjK
kyeGTdZyZDq0jJhV8p392pJh1njQhMMfoaFY2dGjD83NG3M++Ul6aMN5lttX2DbCSXZ1jP1C8rr/
VBCaOeNhu5qaHJbpHJC1MUbPtIHjI0SXOcpdS4Vkz+4wtr8hjs1SNPEX23CQkM0CjRMS6eJ4OOcv
Aizbxd8W0G99nxUPt5NEeAeOMrtartFx1rNWUBLxx0W5YU9woA582QkUmMHJKq0MOFR38/7fZhrj
pLf/sFD0A3b3pUTMfCla4WdtjmFEhPsRj1aJ8ze4FSkOMaHFWTD7F/kn+RW2YuzIOCFh9Rpg3Dn1
v6OKf+n1fkJa8Vw+lT+O64DiHpgXcc1mhjn2p07KDZ0HPMqHRS00rZx7awg/Ot4Gb8rOLzbkQHYv
/g3xQz1wrbTQjwVKgxlkfnSvlcId6y+bgPq9aLxfrWhnCacuHXajGlm10h2RRV5dDNmd2uQV1Xav
180GjsKkfittC9qjxNeZUdRksqEQKOaX6oHwH4ofsoyS3TxCpi7ZBPX4qv63Osdhcbi3xkPr7xPs
/t0EFjT6No4lmZC/01CD1mr2FUWQoOFiMQftvI+9yqGpiiDOVEcTIRYU0QpCWUFnZ1eJ2ML+C2Jq
BiPLNvdUElSMKSN17uf+5mGJkU3W5WAYLdsGH3rb1e4Hk292SA6tF9mUyUECT7iqjWgcprSpCTnI
TeFUtjq6cEMf/JEvWQFjTtLCEzalVyZECWKprL7XGhjYqyv+5g48ENeuGh0VPZmhhBPVFwKreRuE
g0Q9KAaNHRFN7YlV0Odvo2D2oBW9D7p9MZibCdPngY4DVUVuWwIhbivWxyLSnIRkGHTAfj9hVyU4
S9QpkVxVbFEZ6k79ags/u/wXzm9wB+j1pAFKO6duku/2MmF3XBuh17eTCUBHdvc9Wj9msWIhnRj4
1pgH8JHpqGixti6zveXxkH2Rf8L5KijDtAo7e38yvaKuua0WPHeTZBStKSkMd0aiyionDUpYeRhx
Z4qRZazwq5tYbFpjF034W+Uhg6yLxmuehr9gLs4deo7DrNyk9AuVqo8C5PkbiUv7wqzsUD6nXTjo
27ZEbGanINbO/91nOlpex7GlZPDYi7CwnU+R4nlpE+KiPKuIycGzV3YFIT8SyjrIcsbZNVBFG8Jw
KLM0rCXdWsc4MakKTMRgpmcItggR8i0gUCQ2LlOFqw6o6rISufnrjnqEyWhmqtBXESHHaBexDUyf
F96vcLYu/1WuYHFntKv4PUdhdGbxFbQq+lbISGNi99CylZ1uY+Y9PvrXNpvFts+F2hLi3mFbcCIE
YTkMbHyS5FHVeV5MSwZlEDZcJulLb3Leay8Y0COgYHOJ5sjInmtfnGPfzlhQY2PtqkmUwpiN107l
Gbku1pzj6xjdSgep3Xl6L4FBGP0NeA3CFziPOQKcRvkW9eOj9XKSh+BOsnnz6xBsgXF2W/EPXvJr
UtgnZynVRP4BbcMoNBAbLf92+kOv1LCtNTF8QpS4HKbnDBv5c3UhLfcmcX4XSdIByY1n7qAIO21X
WhmX8SLHStdt//mziKbXu7fqWjZobeU2RZiZR6ZFys5ct/zCh4n4KvSpFm4Pt64Q5Oc24nFcmpf9
wYR10Xi3mRHLErxGqvyK5EhvnU9LLkRnPVwFnGbXVRgzCO/ZQ0VLVNt5IsSbDzyEu7xQV6Bv4ktg
B++qb9sIPNqEbOeBtpbkTxrNK29aDSvIJgvjdtpqh31xSbhqESqJb3I+pG9ajMhQIxwpmBPaJIm/
UjhLs59vuqJC9eVMaK55R9wEqQk47GokTWNNzmJqRyKOVR40M1LDRlkSybJSHJQK5JbEEQrZ22ZN
DnQczgyoIWarbDn+/7tb6YckZKZpgAkqjtwuBeVNsInwbBCGD3pOV0ftP8Q4JvHjwZ7yKDNEnlK0
hFqZ4dF60BYNp6+jOKVOMX7rjHjaK7vrN//p1f/wR2nkrBrjdGjINYxV+CUmmz0MlarIPtzAGtEG
k0V2ZEG2komYxFiUoPGc2uINV0U1pz3LdPJkh/p9MtkBBRc0B9cEpsX0oIB2lkDwReIg72d/5Bna
2wwML5LDnOSNZTp1aGtOsIYkZ0kNaARAd6mBuAtgJO1Gw/r1gmyJJVAsGnAewKMI4l16hXGf3Hhf
zfKPwPDhROflX51lXClh1cjuwAktQH+T9acq1Hu5w0RLKy2gVtFGoTMvQpOSrqRy02rAEKXXmDbj
vGt48Cc3wEzZq71/jbd/ZMKHqzA4X2aeibp7E7HgDwjUwvnYz8TgaD5D5DINKgQXQxTUsNMMS7mX
4B2u80kxkdiD+m0Y07jPHv1GCtJuamzoTlPsSWUuq9ZkZGXsLyEK9s/X3Qk1MV8LGsNzFpy1ez+0
cFLTHeRTiMuf8Mp3zZs7zGIMVbd6K1xQrbXmglU4I3GaXfgqL2EV2/X1pYTrtbfkIKITadLx4D+G
MLqYtSBVUe284xqXmfIlOLVsAAhTmkna+og6H27Nvg5aImJPJwMqSY1ikDz8B5+FHeainqYsI04u
lElHFd2SG8AcHQcCqrhdreJSDGRkUO1hUVVewekuxNLDrskoPfi/4oXsK+vobvvLtaWRbolSInfQ
bOniYb8Hpfs/TDFGjPbjXTPsy9zovrfuq0CkZBeNJHg0+5t5XZH61f5m/eY2Vt/YWAx0ehMZi7CP
dlcIm0IVbHX9R8oq7BOFRPnm8rVjjhwYc7E/5oIRw67fvDjbwHvDrW7Uyr2jO7k2tvcnlRE9HGSK
WDmbf6MWCpKPUbsqAHSZpKXE4ogQDmT9Rd4wF23jJTz3Y+vl8YPydE+Vj20v8a/dcTKgXd6/BL8n
T16lo8JVBPqodgv54A0rRl6kFf3rmLJtos/h57bKDQTaxodA6PM4ykebGDy8+gcydHPWXik+vXao
7/B08vw1+79lXa8ceehEBaDErur5wWQ9whxIs+ytCqtd0OhA/pRWR5rMwFauYUJLaNHSi/m6sh3o
XJA8Gvvk8K+SAEq3zJaVE7CoKHkWMqzR6aJ+x0ht+xDCS6Tm1HLqU7D6fPeiCzShyWri8mdlNgKq
kjtiqzPD0jnsBotI0WT+q0RYhLYWhdkg8H1PxhPR/sYOC51zpriQMVB9oYbXsSSUDU1E77OLBH8X
2ZIN7+BbbuplbFekUTKGQu4sUK4wLQLJagHIaNy8/c0TYuRPsMaLja71RhTryB/U4+DdvHQa6xy/
ng/2d+g7UbTdW8cDR22sIDNXJ/rILplFeYoo0y+92cJeaPptWDUu3C+6oNxiyNo09uih6++o+YGY
q2Ij1aWID8UVSa4X1LIFIF+PEetiI0nLLH8CJCuh5IB+k1wQEiWJ4589q+eQXezyTiqipHFBaKwJ
BScr/3qZ6OeDkEyT9GtJlTJGrdrO65jNW/gmKYOHEUCHmdIH1107/JRT5faWOxNx196iulUFfV6P
EV6FW8eqxB2bG1+sMs2awJEfo07Xmsd+VCuwxNDb0DisK8C14IXb+NgHL05g1t95zaSdh6uDgLSB
QLLeuiaVUEh65LDfQepsFGfYP+gRTb93XjA82ndvcpiKhJhTeW50O4YPmYo6mBh3Xcl83C1ZMR2d
7DHpscBM9fKxfthRR5QTlX+qckhiSes7FgcwxMk4N1jh1m98GnOCiZkW7Wi270xbhVA6bT0Mx02A
qtpRxHcIyQRi2Z0a+zoJUfDBB4aS9cYIKdR0ACN6k3lTEWJyTYIJUoS8a5GdBAPjQ07N4sUi85mg
JWgFr9dVAFfy2nHTa5GJWDLxkYziMGynTMujL7KUF8iq+M2PuOCbfYkHd4teKGn2zWPmRVRSLHUY
Nv0jvo6G7g70jC7s6DM6oOl9ggdOT9ah0hggROROrrnrw4/26rekQOSQ4XWhrpOJAXU9RGpVmAfl
xG+Edy/HTt2bwz6cO8Y+toqlU96zaZvhpsh2Ucecc+Qbdai9ctkz7FZmRyzJKJxrN5r8AteNjR0D
Kk1oAXweaRDuVLtJXIejIfE5wk9IThpn4HKt4qczXdL7KBQI4Q8DqFp/YBayeDRyeTmIj6z0sgT1
gRif8x+mZAzAf4WRdFn1c+82fpE9BARRsoR09Xy/5kQhepEX06xlwCvkKaEqR29qKBlNnsjH8gY1
3QGTQNzDpurOzp5+QSTF3pskWyBUbijI4R0ZRDuqRDMPeKi65uwM6qp5b+rdM6MShsTbXSa4QU8r
7URiAvFai6Q2G8XiAQDBtzB59D6mU9zdtabgM4B1j25EWBsyrwf7fNeGszJijEwlQrGxA58h+2xV
A5+mVyL2zROGHw93ABPZIJ0nq9Cm47ydKTGhvoMDP9vLyUQu26xzqcDXgp+zk8bz75o3q+UE7Xy/
ku+SO+CrrXaVkd7wf5F/LCje0UG5TrVzwQs67P/xod9eq09KrQg3nNM9cnH9mt3iuA9pJ3wixK42
KwhaGBRWo2l5XvQpjfqz3BASIrHSmgnA2xlVAZ9eRa9yGDpN8vy70fBrrLw7JTGsxhbMUlntzIpo
tNFVmH4r79NVm35i3mfIuhgWWcwrgULGx7RkP9wAaUoe/kGDT2wbuFqj5JVY+o+hDhOL2qI1Dm5N
6WLUtHhn6VHTXU58fLv1J8OJzFVEmtYd9L42Kzo7bxhUBZsXZKUAl4SIf7Q1AAW1+BuHRm/uwMWU
ozxW4WRL1FcrmWhhAlzwY3Y9lRQ4vYlhGveP2Odd5Ih8FCyKf+WoPq0eQZ8KlLbBIO4XyL/TWUuz
oyvTOZ80vpzcJrf0IJ8ru4AmH5hVsJkxogu1F+F/KEunzMcojU8F1HjumhSrTXZZJXuAUPQXWJJD
QDciPGk5AWww5wdkAB/+IcVYFK2sjVD5v1n9/KwC9O81hsu7HQk5wWcxEOCikKMWYtNLUDBFrJ1N
bClnOsXX5aoCNfz3iUWFoMNM5uLas123InHMNs1cF6z3pgYKSgfQVid+FDoePFMBWlpI4unT04UY
Ms8bvSfHhxJij2bS493RPwGJ85WLRYPg/g03UgpY0CXLyygVDRzLPeNlw7HSga4KJKE6OyRQldT9
TUPrUUK0SjdvUseRA7P5RL67TOuReOmGzN+XBk6j7On/7EGJSrPWo1cCxffo4FUAT/+ES8Q0riI3
ZWfWN1bxryiG7vOBmLtRVufmlE0Lesy/PVVOL+ngnuteA1W6LDoHPA+clIRWN2xJl4vmGREed59F
/WjfY6jWKiMSCA2fS+omS+ABhuS8kOPaGdFO3xc0nYI4ExLqsJ8kHEwMlb5xtmi40APH1ZgViXhl
RQKrDga4OAKI1ddirLUvcntaw6aEyiNmkucnXGeJQBCS/Kj+e2LSpzvzPHAuLeWmL7eip715ye/g
6qy6d91VfHoqTyXdtYKrc/KeDHSx+yRX4+Mhf2Uc8VZCKnKzmDrDUJWqi0uz0OKIOToGsBm+9IU+
XJMtp1wJCtwd6IZHzRg2X6WwAgd71jkkM4TdeoBuOMAjCqhe+rCDQf0EshBzHWMqLibknRQUJRbx
NbR+Lupw/ZHEEhx3HB/JqCRUEqmghC/GEx+lq8MvA10PzkPIRGVLbB25DLFu4lqj4xwW6lqjyYe5
1C+a8Li58mgcUig2LjtJbbdf47+Y0oXNcwBUKX7tZfAC8Zi8vuVLVZfjjbDV77h6/zksF66IoEfw
C+GJUThE74zbtF8P2M9EGXgxE+WY/Nnyrk35ie6xw4JxARIIEUy70StO/1GcDA2r1saCMKaJdSK8
+yopN8hKmXck7MsR/bt1WUElFY7FlvzjbblTAyWvoducKRX0QUdTBQvw9uI8h5AayZS3I2mHa9E9
FOxLv1S+LmuukEsdgJwWqQUYdr0SyzWScGcARmsWPBQU6Bo0IPibDLp5DUAt8f9V8GF1PG+z4Lfv
1uitpiKiTe24XpbYq2c3vcQF0g/yRdSdNMMz1dEJJVszGRp5ri2VNO/6xG87XLKZ/kiLuFIlAoaU
D7yEvQdk6ZoZfiMIN8H8WKbpItto3KRz6bEc+hl567s/72aYL36ZkFyh4R6QSUI2Db3jBFGgNdar
R67KDMupSenKNRHg6Q/ZuH6gjjrVUkMr5enaKNh1D5esPNSAdTMdbCQMZRNV82KjUhMRzIBS2fNg
UHRSYhkT3ayYWHYTbGU0IhJxjc1kW6c+lXHVL9Z8gYyoE5ybZ1jbULptVGW4r68K4xCh6z5teMUT
4tkMsSr7wOOA/hOLXiNAJv8yTyuER02gYgzrHs9YXCQ7rdECdUR34AEi5KnMnmFZ6lm9Zr6SId7H
WbTOypMEmt0m1QFm5B7b9erchAH3s5WOX/om+IJY6/IybKUcw3Bu7iQCAE9X5aFvKPsXVhUYN/Zz
MX7d5BFrKgq9WoxFW4b33bit4j5t8CFP/Zj9HtD+jn5kqZig2g5S1MTnFzSHnPu8S7aorc7FY1sp
OJnCeENoqUVoghX1sqQH6gJoSwkNHi7Ve7OwWdwEVaTqa5CLRlu9u/QPYOhGzSKTQOeKukw7xTH1
2/cijs+LDTrt7Oq6SG8nOotS+Zf7icJ4QmoSDoRgYWzks7l3kHklOJ4JLHw5hAlx+ajvlXwrCtZN
7IHDWsahlHQmD1vgKrZP6rrFFPynZ/ENnbYqjjL6ZiGoPNJMaR2XN3dK2fzhulnbYk1f9kxR7Exi
9ZspXw7g3hgxIhi/6CJPQaN0n0TBg8njiYmK7TkPa2Pkjv5hvHpgEn8p6jnqe3nF+1Wyba4QCKsN
EOYl/QUUSrTTjbKrh+OY1xHk+l/qZU9kCMbivIQapx7Y3gJlR7esXaus2Hw6AYkIifYPpSPaMGu2
KXdJej+d3K6vqiOv/gMvTVJhtsJSUfFwj8KpSSPLbF/eG58JOMtWwqk05h5MX4qdYRJchDVwy1Po
5BQYjMRpgiarDxT07qVNn2yTmMxa4dhXTE6c6gcI6IBa9jmVGW38lyH4Q20yvZ4ayNtYnqEPXLyM
ilpq0ghtgmLfxWHaaqTYQfu9LqHiEFkeZ4cXw4vgIaBjOEfmG2hutJicONn19r0yOA384DIkmmTq
cnqWOcszIzTnO7fA32Uk34P3/JbmyRPQGdYttjcH6VeaKayc4ZtpNmzTv2W2YVc2DzA2LdMcVyCa
ccCAFp+PRX/OuoUE36hvSPOLj6RksMqYApenAEF8ozQw9LPpJ2UyQPi+k7uB7H5KJM72ErcKTD4d
ibuzu++K6yWcErGnrk4+Ile8uFTDB174Vwt2KB9XiJe7ss6O02QNOkbHg7Y8E1rvB70vClUV54BG
Tit9sGu1cGvnO1VaKGjv/cyHim+6maUdGRc2ihzHoAlnF5ItYTa+EOzPH4k7KLGRB2y8NkVkPSBr
F+akauydoobPld0Yk1wDq53rTB2Lvg9VFMKrG0+RX2qdRaKHqirUFgHz2ZG7IZTSnJRPghocS5Wd
DTEkGBLbXoXnloJwy6w7GHKg6OA+seVehmcR8U3vbnM9R2u57wswLBBEl6edPaNGyiy5Oicgoe8g
acc9y9KsiQJzCkAnBW49yJDbOawAQX0kZq2Z60u8mbttRNWz7gHi9hE0yvZacEuIMA82q0sUKLSO
J047LPq0l/zBdggyP2CcIzAl8nqXwA0Gu7GiEkdZD52mZlVPlBO4prDf4rqk/JLUXdmdD/MiV9eN
m5N4ePLhB7fwpmqABzOYbfHyVqkYldMXFnIq3ZeMfAxlYyxK0BQ12xnPL59VRZKxGKRgo6mvelv9
HkTARjPqW5V4BFP/moX9GG19VJjfeitPHDwelS4J+TpKgxSIpGwzm7tCPw9s9JnxeJFEdME/Opm8
FInhyHNCC123l7/P+RgI2a99rZd+veMEMPM72HzUY2E/VizPCeq4yNr6E7rkx/x3U4VvspSRKcl1
iM7r5fq2FmdkSsVNJUaJLcUyZjivDnyzqviQUfbXvB4/z/W40WpOil9oZstiO/hDfOtZEbUbnv6M
kIQBo4JlqTRxysUW35yCh3dvhsRXPIztqiwc2eH3ttfy8Bj3PrF9KS2tlDsUzSgAP6GJ1RuNF24n
0f8usNGM0dJzgH91vbZ/WyfP6n51HbDgyzMVHsCCLJ75J+rnkisgeJKUtrt26LwAKNosvLamUi9T
K76cct04gn3rF/a7s2R5wvfggM2G6qqG4KvJ0Khqwk9bVS1Z2DJ5GCtfQV1x5kFT9bEg2cL9xhOz
auixLNYBeAFRocyNlGwIJmoYJtv+PZOoIcdtO6xgbI2bXNBGxkg/TXSaFv7ucuucm8Kza8r7d9Oa
aw9UIjnOiEu8c+hcPx5rPz1KpvB8qxsnofgDBkuTBawwHAJGL3IMEamQRj43hMqmAfwXHFw7aM5c
VIsGOkM0FnTkuu5qAL2XocaxGVdv7lectiEhDDlf8IhShO7IAe3XeUuH2uv75jwfQlWFBfrMdkmF
OMcFW88qLtk6pABxNYpuhXRGlEsyIm3MWpRG8WMnKSmfg7BVRUsj87byfrKuFaD7e2KzvBxcZ8nK
lphMnFn3IfZJ2fRgpHUu4gllCzX3jZ+KwI3foXOJM7PdklXY5F2Bpz934w15s2pYD+7tSe/KANxC
2qsnos/Qb1Rf8aK13E25wlC8SUcfzDvcJvcEKn9wEJClY69iPreKL6lm5nwdIt/lqRkvLaTFEe5K
KcWSw/8FyVYkVOS4Ooc0mI7tCVKtyUYjIp6qaz0vun46VgYRXoG89jKgCOOtlwO1AzIhPkOlFRL2
XMO8pxYCL4Lo0onxmcAWhJFFRWl9i8Hpjf6MzELAapaWK3M9nyUxPTUj0/2VvD3yvrOMhz2CjPqe
0bX+5PgfMbxld6/ZD196t1r+FQCwiYtpmRXFSwTImYfUxaET6w1mvkSEzKuiBF3ViHwVib51bc6a
W4B7HZm6ykYeIloRBGEMQOoAAdavqdyhCpJPOC6yphKBt71rGcRS052cheK+MPeLyXY8UKuAbWL3
NbBq7sx/qidplLeSys3l4L8st5eGd4hQYQAKbumkTYa+cnhfqMAX3HMTMjLySrH5e/PlntUl16A0
chxv96mz8N/aU2pTpvEJsm1rFUUp2vWjD+wbrK+lUFaGSKxarMhX4nRbITdXedfYMGM/4pi3yI3M
4v+SYdBv7AEc1jujsA4epx8S9la3rRHLc9oVoOZzn0EBsiEEgf/rsXkMQVgF1kEooX4BSCn0JUKj
aG5wXheK9tnMkgZ/lkOP0bmace6r2cDugunLUIuyybjwcQSeMJaKYT+ITBrtHijq/slPc1+JJd1Y
oQUhYWeap6IRrdOJaYEyXiYBRwfS49Ml8jD8veyeyxWKkCpCrwazMA2WTRLudTyfkOQ+icUi3BTB
FkD9EIC2keAMpJkBqR90HwS21F6xmuuAWStJoI3iYMGZjbSxWIR6BfIIaStGUhqfClp+Pot9Q4sX
FMqRXQioLI5T/7F5OoD33M9DZSD8c0fRDY5+qs+Nz3HPXwB94H7EcUzZPXLim45uTTKuKx+cYTZz
FLT3Wo3tJDmfx6S2xp+bUib897zvwHtwDhJUFnhgpBBkMH7OsoVXaVTHh6Y55fP2SP0HH7A8a2eg
SCeXJr0nswqt77x6cDSPArgICW5lywUBsusMqkaVl7Q6/OmOkf0xhz8mHpew49Fich1du4TR2sUa
ys/0uLWcqtZvO1Pk1w19nHU7Hk+a4q93XzgiqTE/49aPzuBa6Thu5UAOvr5V7nhYaweEWrLJaVup
Oaliunl/2aBdSboAhBZFPIpB8E0d6zmI5TaQNMhwmd0I+XkRTmgTjVXFQ8cVhiSJI1NYPc4z8YN/
IDgndpSjcI+kmlOVATIaUdCvoBvDN5tzx7SV1KBRAmhPZvPoclK3D88sh8gS4s82ey43NmuJGgMm
FJVNWS5ruPiOn8pBZfo7hbqiiDRTH3CqSWcgTIeHXyf5QREHg5yyP7/fKdj3W1ywtE62VhFdQmc3
DlBMeltbTyxkEO+CHUOrBPkkhQqkVKGbeeOjH5lLfZJ3aWVGd+Hcsm73U1z126tGMT+YhsXBon6/
rA7WquXw+1gGVA4TVHO0RKGlIxmRAZZlM0vCd/FSJvvcWNHVKohZf8b6K+lHZt2/AG2NyZ8ThhuG
uoLBocn8lHGE/6422mfhmi8URUmtpDB58/2qu9ASV3NatmaNtM6z3ggursTXs95gQkNxmD0AnASZ
z33Zd2Vsh/ZM26HIi6C5+aRaLx4AWd0pPoWQYKCJqb9fCIhhU9HTMUfIfPJtm9yGIXpBz5+tfsK/
SpHhrWU/RdmUCM8NCJ6Evr1Ki6wGYms6PcYEyDmM8KbLl3r9/MaEN2NEohP0FKi7ehwJYWHzySjG
JurecrmNfO+7VoGtNM7MraNWVNIz78jhYVAEaySb9eebM6NygLE+MB2ymZm+iPztTAg7UwLKSVOm
BA1AWL/acJ7MtMxLWmqM0vZTQ2xJJNTSa0ZZ33B0bMf9U/Nt2CsjoriIPp473TILhyqzOe5EXLVx
ni7rWSVARHD39QOCrUwOCLv9vkluQ7BjRwOHnVLz3CepzJTj6vMCUIIScc0TjDUaZbCi5qXZ/Kq1
SdHXiGnHRtW/7qrP0Dx0SNHyxvh5EOEOMiWKUeIYNRwC5bYMHhd+pU5gU/eAz1djlXYA0tBBf1EH
aRLSAS88Cjd8sdQwLPHLLIsykiB9GCmXjKB/o/XWMEHFx/7OabnFOpEQeTMdw088M5ZPYLKh+5cc
FJZJm0+mFPPokeNAITl5nEcfLY74C/87kvwTaBzp0qzxPL69LsbUmrRE3FmArIn/wYk7QGdPVYiU
1KV8ojz9ESH2BQCB4yjK69zFcvG8cAUy+1E/9bS2gMJNnfZmDhH8PHUwCO7u16RAA85y3/d6KJB4
5+OY+T0tokNVBIXqXEnPIpbXfAmSgP8JthTRlpWhZvBbZiCC+8x7HI2tU3iA19Bkf8z8IjEFmfLW
yXjV9by8imgfskblNiIKQlo+EOVMKbn694Q1nd1Xty6OnR4y9vQK0ixYsXQgYvdH/oNFiRKhPgnd
SYy6ySUFcUR/8KC6Aq0nxCc1bPB4yf3J1WgIqYfRemj0ocvewjcC+sR9O+ULdbqHzHrga9qy2/0j
UA9Yfv/sgRvDHfQnWZz8dJidomOc7yREzS5KCXhUo8LVjCwaAfXmW6bLeSCcYAvX0wvNLdJZGX3v
fwDHGlnMPcG+N5J4IrtNKPuoN4rVo+OKqC+P/IH3Ty3u3ea+lZDaOtPXSHbEKqDMvyjg5QTTkKLz
JmPbIiBRg3/so1Zm/SRsMeeKK7Cu3aPrhCh4G5+lboPFUlriFIpHEyCBIn+7fbCYH/OCzPS5a4dd
Xfdswgy7eb0rATObEr4yyEE9E+EIwm/im8tQbY6GS+CMpGHRLc2iQaLO1YeR7mJpvXxVV/nleU36
q8i6p7169Lbpco4IVNOda5nOPQfB4OCcMWPr3WzAqhM7mfQi+GRbu+TTszKOSiw9c84R22+l3BrY
c5WYbDqjiVYoAy8QDE7BakNNr7BC1e8HFFo1yH3HSfzPCTma2zNEPPxzrpoXDoPvmgYyMypRmwFq
7XLQALgRzlZbaVjYvg9QxIAUzLilGOZtddY57W5FsRXMggwfqb/YNEKr0q5H4FFT8R1sY7m+dd6l
4bagkkV344sAupezTBTaNtPVp1yZ0wpZRFBGuPrwpljG2dlRt3ttO5/k91Me35WU7cs0K7SmtIfC
fialf/39wtqv5UC1oiUOUvCNCj+JgffD94k+QLU8zphC9sb2Xs89Y1i3iJ/EZcMatVZLXCXCcjZ+
rZwzpJv9JXzstZSCmXoGj7KDSpXg589PkK9SQoEJwU6WEtx4yYm7SWLf7eSujYBDwtUFU+IVLvw9
mIDVHkIQwPsWNAUWZnO2/S7Fc+QFgYQZOtowOvwMdKusunxjnReOfwjOZWNKPzn3xmiDutdmdt06
nqU+jbm39DVPLiRhM41pjXjRKP/dkttbIDMMeo6YKvFSRhRjOmVAniY89P6Ez7HpKIJaoz6apEaG
NE0dzYg0AVDG3518ieBlClygB5N6mb0mgOWPvbkdyR86yavwphB6qAJ4uaY/4Ec9N+4ddpngkS11
9hHG6V6Mhc/N1aB44ErR7L61itkGBxKa1uhlUFAtyOAdzWlnogZ7YLEZpkf6hV50SEjTxcZGE1ML
Ss2wNpanUffhDE3trZNryGFj0pw4ELrd2OZ+P938dIMxdfmOeV1o6Y7kHsxoaokcI2lsxo3oT5Ya
GtOXO2K/Zt3WWBLIb9lCl5/T2KkzMObJxXbRcDt7aR3SWqGp27cZv1Du6PVc2H2lqV6701QmwUpS
zgaFuXBDtaxVHjWtJ/ue86XoiL8Y6OdZ58I3RYTWUnEutQ4+8q+d/Ho1RTRjcNTvrFMTF22cFeMQ
FrVigZ5Chr0I/BRyqPjz7KSKcXDjHWZyvn4GbTQp6UDzfnSdP90pJOOxMqiVfERnqT/tZEWEvvak
HhIBosMJx+SgOvrdTPzezhSeAku+VCD9LgvVhlOD6AyUc9Uv79aNs4byOXv3shaEPFXdBfbnJH/G
6DQ5lqoCtprphs28cQoDWOhdZEvaJKIRMP2DtosRMN7p5oxkAU+nGFWO+HcEOYa7sSvF1qQU+1iY
I9L5s535j2HxaWx14wbyWjTNeMwOU6+aiJ696uYT8TiWHPXYK5uScNXgehDFXRC5f12VEpfsn7jH
Yv54pqNALUpvWMu9rgw15q/i6v1RC9QW4zGbZQxwqyGLVlmy7w1N6HNNf0o7VTDvDXt/MjbZzI07
RsE8N1yVKl+Vq+urRtDtiTRf99csNBJ7SkoDqu3om+yGcrTDrsLfCeeoxWP6sO1iybiV9dTjFrny
qXj5L26Bj31OphuNCuPMuY5/GTFhi1dnldAOaxjlCgH0j+TTN+zS3z5tHPZp/58MVPskrpB6agjB
l/ZMBGSSXaBkELCHN+99SsZ4l4HOUoNpuEP8pZU8o5l9lTg14Vm2nMs8EyRp/iAVpdB5hn26emXl
ln1Lyv6sr8MMaAyuBSpO4CT3jP8lfKBeZcuf+fzgFxum0dIv5syPWA78WH2fcB2wNOVuHmu49ma0
Eg7DVr5JsYM3rDyXDt6T8i8dh9/5v2vB4xksxnLcFsirfcRM/y4kAtibsF9YPmehrHrhjhRSG9vR
OBPW4lZmFh7E1QT++PHkcYWH+AX8/NcVv73qBJ8Q6pX+LeOJ054Iq7VXmXHYW067K9rBXN6zlwpO
r7YMIMM6uERqBP1aApoat+WmkSAJP5N+yp8QMOA7BG8Vh5PiofLgEEXm77Hp5flVEQEgFY/WImfG
MAAAFAERunNtcVJvEk0YG9HORgw7s+TrBPsMswjtHZganZxykxKByY6yuy1S81dRZE98Waz9wJM4
Q0MIzfTRp/HKCQK+Da3hMPjUvz6Tt2gNZJrXLjFLCWJsEw7aIXAopHdjz5w7yrVCmcwvw7nRApQt
BR2BcRIheJt7uvwY37ufp3iCTmPAAtR4mGt+B2/xOfN/ci+w8pLSXXkO/FAGdkxEVGY73wpypYvx
vpKd+9Z5gnuTfBTy4abysDxfnTKUfYTEnGHRrmnsnjpGHrdcfbuIL8QOKPNs4hr+7zqGjCfEaNiq
duBwZ5FZpDG3qnwj4rfjLDajYN1oSUXEfGoP91HqxI/eZhuBDc7GzcIjh6ugf0PYhGgK+T/DQtvJ
tw8Rc8XKiEvZZ0ZXd4j+ToVq2cuDg3hrR+vZlmuyIW+KzHZvdbVySqYH5+9Lb0oFIx2THZ/P0yBj
PBesQzfKpE5ZXC8FmJzBs2co1YnJiAIOWVUMPt3gSHxI7e6HVDxRndkIOgUYZ4TdHDWrErHa79U9
kn1d3pFDCVQAmu84aQBaVXsBKQ4Z1Pq2ea9o/cx9yEen14VVOF75a+Tn+n6CsTPLXEwqF0q5Gzr/
SVgN/64fjWPYS0ONXy0YrxB7jPpOSqr+k0yNUgSE4BRVb2+1z1kyD0QS+EviR4RTNQyYjwWKy9LK
E7NvUqefmXnWZLTWmpWTYRbyr7HhRUseGtQbwqndVuvcJ7v2Cn4vx4w5eb1KDNJT7+aiPuWnnTdq
XICbZUp3Sce/GA4gKbN4XPM1MutI4wuODWj+0xx0RZsS1tzmD0jLN5qicTHm2LawsYcM1DxWMUKg
P5HzKjgz+jGP4M1U552wKFaJzPWFcbFXEbZtU4fbvtpLV+ufsNT+Bp2mPmPyNu3yq3EAEpvfZTh4
KtU5SfekvDOrIAxowAxLzuHvwODyhu01pQ6ic7xDYGJkV909u2F2+nl4reIn62/IL5IA14x8XTUt
9v+Qzkx6VDE4YvM98xWTbGu0Un1V3pgDUbkoF0D6PoX8ZynVwl8ZPFniNPeHeWmTBnOk2FVH5DeR
f2LrgaUi5bJUn32Cvzcvcz4drBRpND9OpqjAO/71fSMaOi2TQFnbMiQ7YjvUMJqXzEu1IdcqieKE
+CVQ9Tb3bYwuiAV0zUwj+h6UWJpkabrMRbOgzR2dMT936mfTaWml4ThE/Y/Q3z6ZdoouHyXXb7J7
bsrp0mjVOx6waEPD35EIQSa+r9dkCSwHFRU/M7crXmALFPyqh1I4jejJAw7EszDI9wJwhNayOh/T
uKhn/fjlYQJJbeJ5jyEwfyGWd/TNXf3wDQcTHNcANLCnH+riNYKNGuO/N6bq4gjKdSUnDT7aFWMa
y+oIPXTfdUzwVye6ZOzrEkG27htrEzUqLVdOQKPAOZAnxmZjJ9dJgGDsdmDP703Bv6wNyEt3eMUw
jFoYn1tXTXcAyC8OppxIa05EOyPlhvEMyobLKNX+lRYQ+Bd3OpSOyDmiWRzwfxEr67Uz0gFkXuj/
KFM6GsHfJiOcwsLiAjGcj1D5Dw1aoZZ4XO+sJALnuhMkkFaIQm+CURp6DGI2BTT0da0Fog0KO1Av
Iu6Fqk9ctiCJSKcPbHUX0/VWjohFuR74u7Xzw/ZN9buwvwNzfPN9P1Z/ZGsK2mC2C7YIlnvmOSmx
6nIieh3FfyJrd8FrPmIUoSzfCSVc6tNrmfuR9EhNk05Wf1njy4zIMUb6s40hLYMZ7n+i6qDxtY5f
MjFgQ9Da1ITZ5puGWMaujnedeGrTXH15Zo8bn4IzKPB0yBqtyYG78r/IRCo7248zYrKUeKqod9F6
YWgQhZHOEDOxP8R8Vw24pV9Zhs4Cni5mWhOODeLPj+a3n6KabP2cXhluiJf9Vz8J/Fl9aXNExpRt
ohRya25HO2n8K9yoJO5Re1VqbVfSZkF6f87U1adC0cz8ZHOmwXmQI45nqQ0fKz7UL/AVsxGP432d
dXDSxW+c1nAhBOx8zPGv9VApB9kBpzgWEkICcw/CgvFyaQ+/bM1YbwS44xoiTm2/5zbyfIyUvvKU
AJ2i+kXe3rAAW6567Z/Y9BVK09bS1EllyWQCRmMTnKq0aG28gC5LFbKcmjukkRrZ31QTdkxP2CRN
udSwRIAhGMP72GmR1nxDJOz2H07tnJ1GdyPl8jeT4UiCykpcrAXa5T3plem6ktP4gCqHnDj8ks9r
5i9x+kAoUH4nG2yJ8ttx0BLW9ZskdAmDuoywogO2JY/O/DsltRrnh3hkgVLSrSsu9wCLk5QUCobu
jVaTH4ITp7S6iFBwmc01oU9BK0r+6xfUmXHPPS3X+Gg6dzrhDOlCa9CJleutxAkla9hW5nU0r7eZ
LewANeQyIXU33X4KLmNKV7TMgFVkGGJjluvJwrI9ZSi0KAj1uL8Rq8DpB4XjqGK0ycBEXhBEDEQJ
ZqmqjzC/4bATyh0UtaUsNIa26+hzOYnmGTE1Ea5RPzwx296dPvuFt5cYacCLD/O+fKlf3YXATQIv
iWcHJMNkUsBE5VQ6PywQ0qNZiRovhMVCKuav8nypu+K5XSDq/qjNYEt/ayre7xsFb2S9mtE0bY5I
FONtiCJWRHBIWTHYw3bi19Zg7vG3exDvkRUaXZybPwegCZJX7bPYaoXst7qcHB62uaR3EH1sfdVG
+x0LB+UiWCogNQ3Zd9f6TfXIJkfOeeNGF0bAu9MX9MgmUbjqO2fL82+W6s1IUTBjNYeNA2YiIAbV
aAavN4HnTgNMXRlbs4HwuxA1OiTW8HA9NlPgD76gd3G1x89aKDpfetSl6fTaE1/ERFO620uxkbrn
+fSUtGsjPMY3esTH5CzwfwlNOr7x5Ft11cu1SWoKKQnsXbcPVPO1oia8FQYtcC8SrntC2Qj4ddvj
8MXnZ8vN8bbSAyH9u8bQJjYGZrmX4/TSTSssqjwbMBzTO8Eh/y6SCgzWW+CuRV0q1X98/gPTUTSJ
9SpzjjkiljlDNGL93WXWxCYTpC2PppbQ/Zu0cMhA7to0vKjA7hOUuKsYlIVCQ5qFvOYDXxfavvez
aa23z3x4wELhSeBLg2eKr4BAtuyDCuxSo1ZKeQlHl4CSnOg+Ng8NqVBAXbnRkDCzRqdBFSSWKEV3
WLzbv9Wjml+p0fhYCK4NXwp7ESkPDla2CASVZoSDOqz/QGIDdeaxYdSMoyA6zE63k1vCu4p6YR4c
go5HZbpRn/Z3TaV5J+HqnPOFPnr+7/+XuzJmqXx4HKpLSA6B0HdtQAOLfqjGFKqlVV8NLvRNDVPK
Q47ILSku+dx6H1/fbsZ1CW8EJk86+IvuEG3+1DPokiyB9gtHMqAEvtBbKL6ovYkVp6e16bOIpcRl
aJ9zAWRZJv3A5aRcUUkYWap5hPXWFFsPaLrL37ru8H0LSIGlIL4ouf5QfoOxJUVMixxn6cS0vARK
DR83woQtxAdMb2a3uszrv6M8TbQcZcjaQGSvu1OBfyDUHB+oBqBbzvsG7ZZEo2PC3+rIjMDWQ0lu
iznYzRuDi0+HHM/AhrSAvPli7UNiHLIYwKZapQkFqlS47jDbHJQxLFA9VUqiivR9ZUK/Y8J6MkHG
RH3wmmkWqPkEXAR6+YL3aVDltFMOgE+bJ2i1fvTW2xyBQmbkrxVc+FOe76S9gAp/JNsP49rRqyJO
43P+R2Ipc4Syt9LovQLESdhH3kYTZZKPLkxPXr9HdoYXaqk10kKJRPDusXB7+PUwpZrofgq4FPv9
85B6rtwBAenpthmlEkHXZ+fciZU9xWdr811sdSF46VLLaLy6rGuuuSW1d5p8/b0OyYLQOjBHS2WX
dWRa/gEzIo19Gv4YAqr5pud3bEn9gvzAz4ThtThp/wCIoclLhGuOWZtIdbsvLx+Y5nsZeOGI6oO7
uboU8/UC0kN8tZwV7SkhgUNgRAZbP35Zaw4ncttubL3bSynQzeRzfxBxwxNVYcaDQ/1JqitKoEdA
dYE1ZJ4JCFc3Q6xNZGBTCA94KrtnRRufHBgSFLAuGW5Qsf3RlHQ3q+lBQzcwcdoqLhj1wlBZ/e5a
8WVwwzoiiAo+p+nKc2K8PzJJ3aTtA4F+cxskQkmN3GtlhpoI6Xb9rh6x2hkog5K49cIEcHyFdF/o
/L+kfcckm97jSeUabnk3oDEzPXd3QY1FBP5mIDPKsJdFQtQ4seLMZSHq5YGVe+s7CSWGitkjuNOl
PNt3xHQ6iyGOoq4esI/VCdpLU28RSeU4NTILJz7NCIA5hUwV6mnLLhQ54Ca1HxOgDMIkQirejNQW
jjT1spwJpqYQYd67+2GEuIbd3d26vcZJ2RrHWWNeBPd9H83my9KAfBYerhLuqHuZsVpkYCBEFV6c
JaHoLH2BdxXtvyYH9um+joLKTJiH/R9w46DpsSYZJLykzg3wxs4fcJ+bIZtNJ0gKJJOPKehySIi+
4GZUf8AgTuioeiaiHR2rTZLWL47oRcti8rHOCBlmSDz2jHrqIfR6L2LZ/luAaB8whht5YImufc23
MjhIiX3kQNHP28/4Iy6Gb/XmE2DrAQqN8LfawhAtWSm88w+qJznfk0qOfpfthef1nKLTKkjRc7m/
gDv5l/S3cR3KlO1r4bn0VMNC+r98gnUWLazpPNRc1vlMoQmueDVhmiiZw2C70tu6QoW8JPUeAV/r
HnCQHZnw8dHKmQcZiWtK4xPANW8f9fRAYIrmS1cawYrrh75cyzvGlbLEcrwn/hQjZjogv7Jn/nd2
VbGxNe2GvM60lmD8cOuquT69KeFdv25jZa/c7+yxMJOoiJji+fMkALn5VklevS+5rsrNczSDGT4k
HvhGof1Btqhg/WsPDe6fjI5KyFY0uRXd60y9J/IzgAWjJRpH4kokEps4ieLX6oKsTDzbhDM5hEy4
7l/zv/x+D3KdyPum12EhtuRy3pXrtho84+dJLrUlIy2zj8rawtJqND/FEJY/5Hp4zO/W60RY4C/T
fl+bJtDTSCI3sjMWKK5w8E653IPb5qnd4EZyCu76EVysrOlkN0oikLaQZ1LRmhKyllsb0Ijt5FbS
OWhDjasZHUA0UH3wtlCfhuMLS/63enrnE7wAGIKGdc7E7WvxTeNcwCtVEJa8xDh4O7BgakpgnDkU
zFPJmzUDBamdsJsm8Pcu1m75vuqRCnCDNkhwjs0TdU0900jYy6JToEQlCMxUjsK58OHpiak0Guna
EJpZmJnQ/cViwKCJkNLUWMjLtbRHh6CdEuXdq8EIQmkh6FD9uJ2f409xyZns8JjIzlghzD9+ldAE
1OLcEuNHm1Ls+XFPAl8fu5SvgPAdCm/WSLM3gyE7q+dBau0THZbYzfIYQl0Qypd6oh50MGrseTOv
WVkycej13AGiRJ5/w5Vtdywwhsv7VUf0zeU//9sPgck/B0wUgYTraLTGhzPp93n9oigzFd/SfyR2
6jVytDjMG/AS58Qt4CoO1FzEqx9aKpdKpNTKR4r548wNMPDFKdwvN4eb32dpoT7RM1LL7+ssAuVS
dSyBqAbqxNnCL95DnQ7GK6cEwKwDcLBX3zG//UCk4I0Hbcs7Li0VZYDnCl3gkwQbnrOXsoTkr1cW
4FCWDpSd5AmXT+XAjKmc4pHfiPpycXBMiQeBCVxe/ssvOf1BKkTr3DNcyPK178q5iCnGFjKpmCpv
D2LjofkS7euzF+bAU7dIAJib+PCtSJr7KX7kJVvL3ceQb88EO9OqKToNX9EFDPtkAGuZfPFhrLz8
EWQBemPwFfux/BuezvSzxQyBjDoj/keyTdN6SFrMSDuQ9I3qGezvI5doJiznPRjMzWdmezkjV4dz
xK8JRjZonm8eKBgctxtnfsqRnUVrGZsgp089Zwt66YeY/vVPCI29ubSeobOFG/A+6HnmEKmleY9u
2gzq1POfCbqZfgL45z/g5BeCxEgequUXdz87LNCae5FeW30OELAr866ObKXtTNkjqGLZaWLw2Vfr
wKpVPMl1aaxCCZywgQK1AQ2ZVJjdfuWkdn3H9wKZHB7z6ZCTl+aPvk0uDu8q0Erx5EZL2oNcyyfk
KqyLo+oOVeggt0YFnQcS8wDVmcHth6cfxYsdoecHjFSKVsx+BKImqKfIU8WcFc/1Wg8Cnz2aRM2w
CJ0dFuryxxxahkxvKDQWhsd60htyCgmoCLWTZo4KwRxHuTBabpm0Ta/ZvWFsG7Z0G407Znf08YlO
tE4QByLNQlu9fwwfdfELDwyoXRsS2fPGqhEjyU078w6ynHstW+ntYCFK7ReGxxGMweEhOYrAbFgg
bYS9B2B2sZzDNt01JMZdt4opPkeHFcd/GhsKhkTQn6eJTd/MKnhQW9xibI4AhiLe0SKAo6uhxfL7
GTINPe6xC4lO2L8BTNYNtniedFwkgsazkNIa0Ijb54ojewzxNXS6iAMGvE7CPJ9TFULP1tTwLtiX
0OVAzFGAZZ9+W/eWDOlQXu1jinxJ91slVt3rCEgvHpponmyOlAGu4Cjyj9n5ulDWx1Np/7jcAyAx
DZA5O4LI/64l75oywbnysxYAPHMyHhqFHnKlUXnyDNDTpWdzdta9r/yiqLIBtPC3jHpAW7J8rWna
LZFrmNQZLpT+uJ2Hyz7y3HJun2IWQ4Gd0AWw9l05/uUb4ZU0tU2xIJi+4vL4gwkC0oPm7NZbbmum
aHXHXfELuYWiPaOIfhWh0Xdgh1qwg7lNjXWALfZ5/as7fYBJZ2vhfsgW3YUwFH2s4GPY/N4yaTlW
H5QeghIVD0PT9G/igrDj780mEBya9WOSZMWvY7Y6Tj5rTzPnJ0mehafQNc0XxYDNKX2mJRZVi+Wc
RRpzsdca0NQ2o8uBgJ2ddRvDcasaUTKVPyxc8jkul++vwE9w8BF4FKijdg064wh/tpOCtg13m9te
YVRlO1sT2WL6W0WW2ur3qpfyE+jkTqx55sOoPrFi3tXXSLFtyAovQsjDG19CpLHqcY/byZqnlcWy
UZtqsYhEz5Axd2WqlGJbtBNMmk2AWrpxmdac1iv9HNOJ7lKU3IyS1qZqdjzXJjNKkrGsylp8RAcH
oFNzhlXpnArx9ReObtGRnJD8KGTF3WxuKiBQ1++t3atEFpZgCqRawlLFzKh7jE7MqRjc/DiqCNPT
CJRmhEION55y4htAD+pBsjeIPvsjHcewvqZ6zQU8oBQt3upGvjKFS8qQSD8HDMjHF1n4Yoi94XgC
BORmr6gJD1RpodSKYL57jN5PA/+ffQgR2LR0/+KctFQRubntTULQl9Z/svKMt99vwU/pgeOyh6mJ
8C/2mHZjEYdLpmoIPs9T+OVwDE5nftKDZ4zuK343SZWI2UbfGbXqlWKWW2NIXkgyZDTM0KsKpPEp
tpbQ7ozRaK6sXkTDNO+UJY9HvHG2lpI3w5sJkvbBroxvZr4l4adoajkK+R4uhSwlSVSQy1RdXX69
nkBN2e6X7hWxzrkPy4yNKGvXQN92/d3I7lITZENzJCgQRNXs9UakYL2YuMs/BRhbYiqSB+id2auv
B6jU071mF405C9IzLuMgKAmHkC4NQV4diwqovcNczl8wHHO3kYS6Z3ftII7uyhZ9/PZtzqOk/Pjl
2/eFPQaKPHftCRtq5Rnj/G08a9V2HZB9aKqIjOiFfcZArVcis1NE+RKSxQqSFabS82HwL8WsSn8U
7wZcXSGXZv3dGdJS87YIF7UIz6AYdKpF2DYro0tso0Zktd9EhR2E7fS74NfoQHAA71HnJAzdSwIU
7GDmcb7Btv/YChZxKFytQhEb2LGfzMWf1cVFJpfs6XLiUWWKebzzDMR8JCKY3gwRuglHlwv1a28I
QPsUbogu+BKk/VLNGwXdydaVpWVUYW0bSIJhpl73LSW51uxHUnRGze7FdJmGwWSRDCTbaXGWodbc
t1m5oy4QtuwL573oRKjrKYA+ewHBnr+Vweo5rUfG/CihXze0cqDOOupujfNxsa92P0U37Qq/BSQl
JUr97YR30QP7M1SxoUkuvt/VEVh0s+Jw1ViBsNjHHcbMmuMPjhWMz6Zxp/uMfc67dvA2Sx0RcePw
h4S39H4guY91mETaRyTuJEw91fC63+B6qqh6tk/eLugMuJT1pvbmVN82NQ7G24ggKmvvoMNE6FTs
d9c/JhnO5f/rGZuBoX0bqjWETRT+w2nBNBa+0ux1ZwJYmgBF30b3L3jGDD4PsWr0XqyK4NHy2lR7
YuVTFovXjEiBWdzbgUevY4yLrpqw3aX6COeGCaK4tfZYEQit5Q1bm0lKj6PN0uNHpLE/AE6hBj8A
BMRcmAZQ+X5uKVOz1Qf3KwRQm/k3sz4ZGSC1xVvaB1BentNgYxyQMhXAZsDhfPl9YGNk6Fx8ajy9
lqbq1R+AmFlL9dr/QC9R47p7Ulr7RLhhB1mKFX7a6KCm8PF3/+D7ToHkMO2CmXtQziPr/mCyXVqg
szcMU5zoaSsmhHH7z651YZZGdGkS4y+8FutpBV3dh4c8CbCxah7BkParu5+O3H8qxA8LE/p7AMPm
MHHEH17NmS/IbzmJBPyocv/850roAt8L8oTMmYabnoOrCb4VSbl9/prbkPlkpE447IWt0MyRYFQH
5DyHOvE2ue8cvGKhpAxJrHCl45Eln9idAfhQfspizURAvO0Y+08od1cdmYIRefIJe9Qzd7HBHSrj
pZ9PLOqS3SrEa+KR9rv3l5NJGu1bMvkdk9eP5VKgZlKyw3g0TdlrfbJOJ037KA0Kve6om2lxR1Kb
eAu64hWYeOOujg3cc3w4/RbPu0VVSpE3QHceIAXo5hvFiyuQaSaDuYmrXPZ2/UEGQr+hrqMfWFta
tV+YjIKAe16DGXO/Gluex4HK0d5jLDx0ZzbHRRBxOzSpFAjA8P/8rm0Y+qx/Kjp1etpMJDEnaqya
n/QGPKzUkq/xs55ILAOrF01s4fW713Y5Vt3lGouPaUYvABFPBtmAucVDwKVdDjMqL564AoqJPVbO
lGQSAcZcQmkleyTlMGnz62YaU0hv9OvN5OihPo/TkQkMut+Mxk60M/Ui5db7upeWnnW1vta39xt5
JzCzohQz90ccosU37mpZ2XUwK5LV1pZGhryPZk5wk5dw1HP5m1d9sAgVtZXZx7nRwcn4wlOXzo1V
u/YTOxjpo0pxue3dy+OQQHn2T//8l0ZOrZo1b28Dem+xsdzzPwYy3MRF678nuWcBdCrzhd9Tjowr
xXrQxeRMWNQIX/moLNgHZ1fm3N8vkrDM9/v4ax+a1X4+5omSrm3bGYERiVwiPtzYgvS+pl5aZ24S
dNOhvR9FePbumFy5Lk1r20zTPdcRGP27x+iGPWlXOvKGB/LSvYYBAqNXPjGM5ldYiuNL5j/BX+rw
sX6txnQmnQ3MORVrhr8nsiD8TYjTn8OqebJ1WVrGl2uZZrUVKC7o5B4wwEc0jX06uWCanisloukQ
yYM9XVCmAqg0lht7DoJxLMuU7MHvuGvdSkQYHg0MpVi/v+AUKnjyBATVTO9mj86Mjb0P0AEekhPl
lnpSFclJqZlRr+GU365Te3S02IqCiPH8qd7hDQ179j9K7JaOyyznd/OUmLgb/PrIrAFLtb8VuPmO
s33wOeWVK4yebmwMO6HEJbPOzPWBuZTLGSWeGJFHKMj6s8pUTglSMOngQQQyakTt0xJn6uEYcrt3
I53fBXOiJ26ruInAV7XkJQiyk2Y5A8eMG4Ffj4cPbQZS/TRYVCKRpJpLwR8hb3WHiioPOyUoUzvQ
6rKu+Lqz/l9iVh1DNxn0yEQneld0eiRjtEa1zVWzdz/u9bBl0K1jcTa1yFUxoCvPPid8lMJ9fakL
5X6IJpFSr4AQxGEyK0RtY+sH926GGnEssCpoTPthgHh++dgo2YT7WC2f5woiUM5sH1bVPg+1XOr2
SbW5n/eYa3GSQjzBjukM2pZH8VYHhHZzo9Gd2RB4cXwKdSFW4VamT879BskRDeBU1+SlMy9eZpx/
WIPS53qvxZRXdgLtXoNMSU7RnR9HhDzSnPL+PlQrUqisnSEb5N97+es4UOXoDuUs5glkzz678jPS
LWFxXuj7dUMNH67I3EWjU3CmUXqmFRH3DNfwkMFfxzGBDbJITgndhmdHiBnf2opxqEG1LrBUl7Gs
Ar14TFelYb27ce513t/PYR/gI8Gy2okI/r4ZxSh1LmbAmXxN3/FCy3NAypkhi/6bHb/RbJzgpUnb
PFPt/E0Gwrv8GjOO5vRzFVcgWRwJMPq7iHYlscmx4uX8wWXOcrSc1Ca1GO7p99QFDdwIWi6I3Cru
PqpyPXhwHbwfXm+l9azHNt2bCFaOoaywy9gSkARyLKJyE+i5HZ0z87Sof1XMW4A5Xvtpjgqi+o3o
dP02CNtGKEVW9AgdsdZwPj0sW7Z8aDoFxNVQCYw6twpprdTSRZ9vc3BnEPE/+NYw9HWj9QGygGkx
ltxwcSSGIig8WlV/8nOwM/eIevKZQW5qw9QEEdRKQ6kvro07RCN0wH7EDBT9mAlQiwHe5a3AjKir
7pSE2Sfuj3v2/oXgJ855Xab4PSj0N9TYf7IRkrVMfAsfgXTcxE4GNTW95el/rxolXIwxDUBrf690
rBwlDGHFoS3PbLeOcC+Ak5fEjBKStb4rSIXeeionNBfbmkB2iHNkz/tklPSTIq5nQ6zWpRVyiVW3
g2cB3kL24VIcY2jn3UUqyOdVhK7ytRip7dD1zJ+zDbnuerlKT11e9np+jd4RrVHwk2rWGo6ebq/i
7mu0mUdV1L/yHbeb7VhRtKQD9zinR2Dz+dMLHgHVg+4w/RaCq4Ye3cQ1mUb8CLQBtQQxLFBAlSf6
e0gK1U0KfbsKlkuCEKnbGDEZlpP/3qEbcn4RZjHXGBZNd9SKtvd8KtZLCntikv0AfyoluN4zsclz
IsPhgsvvvULn2frARtakYCJYxup7E1g5jb1C8hJbOw7rNcy0o1ZL4ijm9WC5S5uSLzHgKasJq0MF
4k5gf2DI/uMo1eQeiRbdBcT6pT8vXqGOZ6VlLLmfTStpVSf6rui8z0HscXykQ3GndsUved8QnUrK
0u9GQwf0+x91pO1E7/D9s6sOD5xhSDAr1ubcCka9Bd97dTn8c4vSPFsiEL/8GgV8j/EKfeh6+vrW
uv2XDDRduN/nKz6xmabiUC+rzv5QtAqc+FGmPZkMwuq02LGZQ8Rj+CRoimaXJwZMjLN738hgSQbb
Wm1hLHHPZh1Xx6RMGMsA+ZoqoukvaBJokWD6kuSPzG02y4DyI3M9mwoOrpUobAxAOj8hug4DeeqH
5R5nBSF9xp3HmXXPIDK9xwyo9Q35mfk5JvDR2XlrO51cxqc04/Y0VNHlkm4QhUXG9XbxOhvXQfhC
6sMcAzUQrbvfAyfZ35bxP3aBVdai/SZziYN1uxo9keJcIlBBQI7DC/G50vEqipgRdnAfbZze4O/C
iRiRsmDSDIrJvI8Ndvrt32MjQkDNQ+dDbyv5k7Y12g5fifg2JfGWbE9dgzxlkGpvdfkdnFObN7I8
U8eGTvfLv/AO1Dhl5SAsJ0QrjgX6+FDOFVBPWOxTzEk6BxpRM+aTRFgSzes8IqeoF7RFXm36xvxd
28ef/J2Ou2YUP3gyUhqRbZPSn8hdKwWw1YZ3vp+2FtGDxDWJ6qHev8oV0pjyLAfDDz7CIRuz419h
zSweNQRndCZqdJOBZR8y1KbI1/na5WafSxAQwkirm4gfgI/BtCXc9WPx0iBtK3HLOAF60nCLHGCt
8GRcYGvygw5YlSlF4vWVNPvMqx0DWY2/Fdsc2tXTkfJKe5s2XwsRnW9Tj18V40ljXRoz+96EoG3y
eEnTmxXl3b+ECuvUuL5ykfSJl1wrfHGVeaZnH+/+4rYX87x+zFpuN3y/XM6lyCMLwHjyybI3E428
v8eM2v1vos7KXs7uGKJNifH310a2isJe14ecTjQb82w7u/59ZTqE7SvSZn900eUIvpGNdJ12gXSm
+nxh6DMUJAYLgkmxHZjO83AAIHwN/sUuTxdTHU3XTT3NUh4rgl3SC0XkMc4jO10kAb5aUZ42endu
0rgVohp5/LeIxq2pfNRYktXFZvB3wOlwlMlLcHBihZF5VmPPZ2bl+YaBimsI6KNnYX56hK+Sx9L9
0Oio1jqd78u0noUJ15qHdxL3G6zhq8TgJmCSrL407d9vm33tONeRYxikwnq86MHkQl4PB/M2R+ET
GxikfJ4CcwkbkKddfqF9SHTQUZOBqeGsH5lvXYNSwpZtZtPqaVWWjlqmMiaPHBf2+kqTBT9EVuHq
7QqR9ZlmWAAVAPDyAeFsYVJuwY9sT0ZnbMEhPmZhCQMolt9wmufwDI17ePKTut127y7vWHxssbQk
nz+HO8vpHKnOsHj+HQKCMLyIpyzyXdgPUJGGkaw9eaN5VsUSByG2X1bP9nJWQ8N0WsKEn348tEKT
YXC86dkCoeiE+02l46mUbRI6OGtd9ZouxZYUfpBCLifDMHPSA2VbQvSvkLDQELURfwrs05EEi9Qk
Cge1Aza3BbScCYUeX8a8mZST/DH3iUy6QfHWhPVt2p8KnF1AhZZLNi6xY81xVZ+o8CVXDv2VyxmB
D3S22n87Mr4NtFB7KhqKy2gLzaT2k429Bahde73hPoi/6YJbEbM2hju1fxL4cDArGh0MCoyJBRGC
rK5sVvBm4gcO4E9LF2DTHCHk+tFI8VXiN/AZrhW4uqlJUUKAZaeF1Wfo7uJVY3kVPBy+qlfCaxSj
xbRYY2+ndKbpjETGYx1o5p62B5w24TKqpYPZyI9yM84hCi0GoovOsCVqN9/f/OuVAp6odGMcjnJU
w660Dp6uDK3dpQxbi6fxBZORBt1B5bP2cSvZm1PjTPNCsVv+D1xWxz4Irzjbr34MoCOhDfhO8Mt2
PHF/RcEjJkLOG7bxBIFTq173WAHPHH7g9SE4+ZynkjZ4li3313Zd8uRPb8PQQQNa3Up9907mlbfg
EsujvVLgsf2FXIinwGNG3wfEx7TlAK5jzvW7wFxabA5Y/wg3EqotbI5D0vzuLkhOzTI+8Ty2pZNH
FS74/QQsHqvqwzKS0A3AgL7SXSV0bZuVLa2/Gg3iW4PQrknekjQMWlSOmyT2wtHVJkH1DJfxgEs+
akXE2LYm8ebTYJc2YLpi9KlQnLuLyvSwtb61INm9pUpEzgu9LYWFATHE1whclXLh6hyMF9N1cqay
hmxIqcbT/ULP0C/f5q4rHBE8zhVA3j5Px4PxMqjCEN89iUWmAdK1Hg0Kv9A5e5QvdtTKkSBnv3KX
awX3r4pq8GAZvffHcZPSCQOfZT3rIjZebw090GTAXk815NOMnU6ARGFVkbkPLajj3pgJAyP1UIHT
KTBV2GMYN8LHKZsH5zKFi26YCuYsr/lrt0ngTShsjzFChAjeEtWGx1fWuUokbrVfubOztisI9yGl
xc2feJACrVUt93fsepeOxwevhh5sP6YgiVnPU0l2Vd18vhOg/PIN0GfnbcqWHh4x+9VIyoIDvToe
esltA0XKzvyvPjz6FeQVA1OUX9kQqS2Wpa/G17VZE+oEsKR5hbJj3huN/rsZGovV5uY1d8LrHqWl
xqe/WyMAuaoBz1lQIU8HIEFHIlo5f/bT7cKZvRJgeDdNmFcvNggcfmY30tTQR4JFA+ON/FXoDQ3D
gOVq1YTDHtoboGIda776oClFVfH2lK6Yf3FwjWL85r3m752utIaCZmxZokVmm9yJmSfEEFEdESgl
LW3Cjx0NfM4XIu6J1YcgIYxrV9MZSXuNbsacrd1C6uUe4cYtGnqa67TPFDg/AHjx+iuxQOK1q1t2
YqPQWwOkBIjs1jbyZs86umFkD/ak76ngrKk1lsqA4KZqw1u399GXRhYAskuTUflfQWT44Y3FoxDf
p20flpjZS848UwmuUMpjrl3KxfrCdA6OWxUEnDQvSBwlbL1l50bm23a4IZZTyspEIyl3BXtUMfAy
kWFENmh+bGMh6Y0wGEe8F2UypRpL5VxQbZ9Ps157OfFiiTh+/6tXOx7qo7S13Uj3zrOHZnrfSsHQ
eTMr/CXTv2JlMO2clLIc0ouFjfgrq7r4WpaMNvcPLAP1uYbj8zgHBl45Ex+1KEuSljJuIFq3Iegd
m+5ffocydTKhxdpgqmZ8Uj+4/pO4BzzlHNBNmX6BrA5NC1D8xjuFy5HMhxNmNZQFJ3qoeBomBjc9
qXn39VIIo76WxSGIcD60NN4rh28hXzyTu3e5yGkj/67z6B0zOcwdqOPIqUvBGhXiwVTQEu2xasPB
yMUGcCrnE/ATJzQKvzdgGNdUeK3oq2UIyVEUeShjc5FI0h6VvHOXtOAOJSbNOx1KtNQk1eZQfUyO
GEm2yvTKAfK1q5HBaE9KxMH22rpaf7Dm8jNl60MCC45AdlkOOLQW5mGrDdS+8+vrG4MQbHN9jToq
uR/xrg+/Yn5Hhpn+rJDEw6Jw45UBvGbbX+xm3JRkDrzZpuP3oaRfopabLZMJuQnwJLBqLFssXIAb
9jT7/ArpGbixmDdXgxxGT6UK9qcN2tgsj9eKnBqLD5A26bVBR+kVeLOo1rwYBbHFRh4Iq/1WBRsA
FDns1sdODT93nsxX7dG/lSOuKNWvzt5ub2ePp8W8iGhnsuT8Fh+9IR9CKRvKLUTeeBhiMDYLZMWV
VqNF5LJuU2XHs5v3Yf409Tb+UaOCitPxalL+JRPEcrAVd5M5ZjGSW46Atf4CVmqhcaT5+r6WP4H0
c7H0wWB/kNcQJrAQEZ2MktGh8Dh3n8C5HOk6WhQ3Ck6po/0aqkHtXgYn/pLUg8zKlivcCMV3AsX0
3EiRV7t5qdW1LWk0pFOT2rRolZIj48wONjPrOk6Z2ZCCtg5JlfPQQMufYUEHPfb3fiWFXc8C5Ss7
NJqR7eTnqC4qgxjQNiT9SsmxRunUTmz/PG9kuVUsggvCbvrKXeuCLyJVrWFDMMwprfh53CCwKZp1
L1uZY9XPzcuzjDPUJlc8GwgMQhR36IiW7hM1MZ/6+RbFz1K610wO9YufnNJs91vZAAfEoMsswLAL
1UzYndK8+tpPuc/Fc+tHUXQzOPGKA23rAyGpExt+Ps86rnVB3msPYuej+7/9qU9DQrl0dGwOtjEw
yum91/MvlhRtNajZwV1nDLJwlbzgsUTUi8aYaIRxp/aKPua4k9lYmqregxMI3AmAjqasDMz1WSa2
62zq3ve66QVzSGPQPfKQ7dugYYdLR7YG96+5/O2S6yBvA5WzZktxsm2mC6VusgQ3VyMEE5azcqnd
jkQouRPkFoVIMpexXTZIyOmQ3+ufuYaplhBDb5H8MgZyvTAgyZ0Zv4cJ0ZZ27QZ7gTSCDGnUPA2O
Ns1tV+ZhJ9HxUHddpxJ7iPJRTuS0LaHzL5T1JW4+uS21hdKU5KQOjBq2h/l0AQKhvoo8tWS+g2x7
MM3jyx+Yr7XGxZNAJ+Kx44kqgOitU9P5YelPZTg/Jofk066yPXCjLYNtqvk9Nno9QUq7lzIX0dUQ
5UYZ/TBxz/hb+3n1zq46lgYFdGH7MB93orR+RHRJTg0ZEozYdq/UTsYhWKp1Ffvmvow0Kk+DugPZ
Le9XuC6iGSAx3BgC9hULWDi6BRGmGXu5Tog1rCW28HcB/1xvDI5o5B+9naWvgoJlt1dP/vfjcNZL
Vk80vL1Oa1pBXdynR3IsW0bLwCoWdBb7cYbTVasa1HGHOIHO++xPPw6VS7jI6aHVZU1c2w4wPRqD
8zpPXOnCBv0cuZHIj9uhAhcGPeNdpMHqh9/bssgWE1OrKXPord2MPjq6m/m3c8H66SvUzflH8Fha
zI0hUkrdWkK3Ue3QYkzEBheoEaBfoQMB9BrTybTr/gyqVmSpgxol92dK3yaoVODF+xBEfzp7/7eV
VRiWOX3yscfC/UAohUDVgCnMMcCLN1MSSCsl6p71E/txkBLiOjVZYFAXDuSr3xphEe6Hefilfu+4
yhNpU1aVRAAO5Q12kac3p69Z1GTiYcQ3KwYsOOqZg9KdV2t92hGD5JfrvNOvBJLjJ1qzWhZgUity
yDkzYlBSN3wTgiA8bYXS56NdkQ4lNsIH7SN4NmPMLX52CL15BNBrpX8EW0OFeNc5LbLNPB0PYTzs
bxj33UPQnQPcWcEU/xfs/SRij4R5Y0gA1oSJBO4H/gD0FjBCgpc2PxkDp2ApQZxb8JSAjyotO228
cu4SLcfgOLtLMfen1DKiZ3GT9VoHcRCROE1JcDzz8JTMCz8IltHvxs6nbpEhwQMdKeGjTgBmP6Qp
o2ksjHvonaQisB+fQuz2kp7JQ0XBhyMkukhCtRMRKahTP7N14Dswgg+kjtjY7aAgXv7kVCTJgCJ8
G0sPQ4atusX3k8+1OoPZ39v1x7aiy2XIsEKrF+/BncgsR3hfOh/wROdAAXp8Yqe3ZXH1+2tqi51S
ve1lH5YGCSblqbXgvfdLOMzTKpXWIKKZGaUap8w8uPrcQsrw53XA+YZBaCLfBA01emZGSnMzX8oV
DNAkYwBalV2KOfmG91Fp8X2X9tMYJKh2QYUd7CtURESDwGGx5kH1/FzOvxhQ7x5FMCZMgM2JCRob
N8zDUoYwJXDn2wRnjAnofq40P+mZGJUeNchmjcu35zM/Phssf6bx/gWbviMtCYIYkz8sE+99ohoM
iUV/MoluhN/YI2pQCuZd3OY6TuUgHJUiX95EdoYpNAAuqMQuGp35rmnWChDb9NEofZYSzSPBX0Zg
8spXIXocijRql3EVUj3AiN+P/zTRVZ0pRX84MOYFg9UOosIuojj0Pw+cWDKp6AynaG8lsF5cVjrC
Z2j/BrOm+ks9t4riu9rtDjE4pYR9rXGI7AJ+93D/2OuENDZHJanYROPBvf5FqQOW4nJSeTqSPkpd
I963j/XeIv+21kXbTfiyvt8UvYDHitVYZt3sm3iJmHZ11NJIozaxC2En/nTihBdgTtotSiu4I0av
hZhLGvTnSQ0+Ucebl7sF3BHvj/0uEtK2haYi7nmlhPYFvBNyWXJYq5mU1F5QwWGD/ICXq//MJQI0
SMi5H6s5sdOMA6oADeNf4fGFoaoQnQI3jA/GEdfifI6BVx3d7bvgA7jfINVm39LF89dgLtP7zHkq
IGaRCGgKmYT9g72yHGN7WBGrGL7KhZ+ethtpg2gDZwh0ZFdZ6OECrsSwpUtIdC0TPljtXrvHOqRH
8CGelkU23Y415TMB/yNram5aWvzxiPsCVUjLfzeGLkxXBy7Fetni523FVEUUUrO4mfDMQb6NyO/c
SsmXtmxRqI6dK/JgFFlZEqQqHZxklO0P8SHtJ3XXs2P57LwUr20U0ksx6WXmSeZN/jMbF5wGWnaf
Ej+2j+tzzLZx5fM8jec4hxCxYTYama0+VzTQvQe4mXgXmfKvXjedocziVbnaRJuhMBDQqDoqZevA
AJXQdxoRbLhiRwOJpWvlcY+BVZXTLpH4hnq/hXNnXRpBLfCqwgwQL5QZX9ORFVzpehjwDoH/pI5E
9AymZyXGhv3o4h01KAbtsaZ7Cx5YEDKoKpVbniKH4VCusnqLYBZjxCovcYx/oTXKlIF5FBw6Jj0k
R4OFQ5FrHDv1z89C2Dgi7i/2biymzZwa83jIUEx9yVnigtcHjG9CHiUBHxhGhxH0+/4HwGufQhAX
g+wPvZGwUo+IvnhU8bXmV5m518/suADpqNTUmwme82vPDFmDDr5eFMTXdl7bHGy3zGPHllskgo3s
7XpEQRYF4Q22rE9D7Uyo08VDeVkREymsHqYm2DwZ0OtOsKvCIcu8B6MOJLpvYg/1Aav1E6KVdLzf
me7SSDKneWuaHGHVHLw8bcJfDOH+npXmmcH5Tu7+q2ntfoui7vulLPl1IIucnnx5gfePilaTvMM6
89kVgO3unbkT4YW2+jQ9wGj1n86WWoITZds8NwAALeF48y2i5I3IUks3DSKInUl6lggIoZG1HO0/
DUY+RdBTKMs0uv0HuHboyqssZGXxHu6L0iswUtQsmopAEK6VuBGs8r9oEpag7ztUuGP4XyKzzBoe
0iOkq5Cd459kAv4f+eWFYTfqALD4xHvxVQgtbAk7pMI2vbxKPD6w1793HIh/+JSgTBKytRfxVqOD
6qs7yVMFjtO5DqXuaL4Z7X2tuuR4pS7aWLp14gQHIdVbV+V+HNzQZF/HtJBOwvwq2AFOcmV6/Py8
Xe5zjrJbgJsHPcAtPfIhUKEl+IuXVIK40T4aWLbHZul93rTAu0o6O3jQDi/+FwHFT9Tvu7iCHLqa
VoVWqwxNb1nWpGhA5HCNUEVWqGcqrYtiMbW1ukKuk6Zs/PsPX5rJOvk4HwiTb9k0F3Hc4hZu1XlA
C9VoGzdbXIyizrh7tiHaE17w3GSIumCO1Wpn4f+jTil3ODz9toDS41y4oWxpelwbCUJc9E3EEZNz
34bnyqU08IrLks29LW9L7O0Iq0lrDVOjBgAUT2NfLtTjw7ArvMpJVDkWjNHgkye4QLJ72JqoyBO8
x2FZGfQUMYmLFjeydinAARl9cEkHUAyd6NN5wZQGl0QM2+ezbcLMjarQPZDPHKk8tazYK1UlQi+r
O7axLlCnSPSi/xHkw2cpW0BJ0f2pOjGnNg1kJP8uJV7b0+mkngowG4jRd5Os4IU1q0NSwCMLekKX
uMifv0AzZn6tEFjV4+3sATQfgpSQJsaQaCGwxjQueRCVlJu44xriIs2/ATqumtvBa/5HQlV7qWZK
/e/xIaVqFKrHmnxH+Zl4WYcVyMajeIzwf4IRu13tog9EOss4yCIW5804loOs4zfQkgrVA31NojHq
fKP9PZNLyxiBYo6eFvXBQcthyNzXiVFHsfminz6YDh0Sqm6BcVo4+5PLyTGIhxzTZyPgiG6AWW9p
jVLof1hjVKcDUNDUPVlvm8T6xwvQC/AG0xfqonqcNilj3GQcgA6gM6ovN+aBwEamgtxEEu4g4xOC
e6JP3SulPSpjXMyNEa6ak9g8YKXuycUJKAt7smxpjSp5P6ny/eSnSZRBFa40FnHJ2/xpfziq3A9V
lQ0Ue+hvCobC5X9+jGE1mh+i+GW7fH1e04rV7WUgF/KGZPrfdMWN4JBVmSCB21Egm7VmcCHJZuP+
jdej7ctfGpR9dMrac+ppeesL1YRcTu6nLc6hLvqjz7tXa0dEvIyr5BiRCfCjh4fk5JlvtjCK15za
MnY3QCcHCa2mdVnA8SZC/6SSvkn2wmpt8XWR1QJ+GU2L34SNT+X3+Ri0uiWT8g61USnN7nAknSgR
mhMtpi5CiOUKFcEtN0A5imtlvL54bR6ZT0nHYydMScG6gpIkGUp/HfYljVz1xeTC1Zk8WiItF7Dr
iwWMwA3jHCtt/DvvgDpdMvlBXL8dXwsmJhYKIDpDRjuXK8HeC5rer8MYbzW/F9j3RME0XGBwbZJN
v9JrJHNdmajbCV3Nk68GmsuPKpBPcNvyGMI8jI9IVPFg1WPAiCopaTHoy4uC1FK4ZWn0+Rceq+pQ
w2C8OAvddZZMBZT6dvTIT9wkooRjZBrqPR1DAZlrXoZ6ogRIqIvkwxURInC35pflsJqryOuGgy0Q
kFWhzIQlkpXaG1rt1FD5t/ARQ5WfAdaj9FulMBSioWmou7eQv42ZZKaXD3qp85C9IBZAmvLD3yA1
dgAgIrVuLtneE7ReKzJczjXR+FbD4iSwAwlmHPhKNZDma28Nz7ueIr1IG1xl4KcXvWihZeRNbpXa
q+mjXLfriZNmxLSjQs3zF7FXWBml6CjX0+Lhy9J2DyyCEMVWLyJ1glYjVPUs+WA7oWAFyS0Ft3mo
3mXJto9VxN2Ucn7tNXZZcvzE7kCPJP1WQD4YTcP5N/jEHKNNY6Zc70szzCLL+iUzOiiQ7qp4enN3
tHJ19ioP+uqFj3OvovREzWRQ3ZmXT2Ws5MpxAPlF+u5cU8JzPGTiesGbHvBCg2dEKfaPghTpgd2Y
o8MTMqPO/BjR/jeif7R8Xz+ffDFrcn1RuSb8ShXo3HPXbMAdoThyRoqVNpTUVRzQp+8Yz7Z1+1v8
cMxf2MDdFCBBDLVAUDPJbFrSgk4lmsXDXFk9PbUPYVuZ4o3+z5dP1S5X01O8d/wEtB28vR9H6+EU
WDOsfAlQeL4kPQA9FfrAu7T8PtdTo6e9NF+M8cDoyGdmenXAEbCq9BfXhLdT2riJiPrz7ddkB6j7
Pz+yGwlDw6+Mb2EHiJAz0knTUgfWIb2IWbyKdYIe8luUVeDeW7YBpeZmFX3ItblaNNU1BxRf75iH
ycfdsuXOjtzx5WZGD1bsytSCQUSF0gdZr4vUmmfOZWy/R1g8UUuA+V6XSPXJxSrTY/oeGUfKm7Gl
W33Dzf+s4i3lg+mn0wb2B/xth2hScVSKewIWtiAG8zHwRKvEvPeYTfxyQoCdBh5CT4VRG6gxIJQ4
fJQvHTWsIUpIkGpwjk7L5RyqBs1QJ3anYxbvI4wdVWFbTLO07KIDRChC6CCbkEgPbSCN98FZ0Pxb
htwQbKBWVybTZ8/gPthYcpLJfGsgrIhGmd7mlxoCF0p9NdLt+RNTGtjOEJxGqYqUjxgpx+suXBLK
Ly7bOKo+p0u22r1cAtmFzuXj0gpPx3WvmuDkaAmR0WWS0TuCc8U50IcwNEabGcj037L/aecK3HVo
YcFexmxUFT/AUa9pZftm3Y4QUSiTR6/958t+90hyLDdmnKAodOrR4dwFjpX450B5BoOsAPlGIL2E
W6hDQrt7HupJSj9k3mdKd1SoyuPEJjwvWvZsx4GB63G4aRX7XDz7l1EhDaEcda7fz2GNTDoPkr5H
Y9wDEJIA1nNb4jYHXttCf0bz5TiwGjFOunms0gDxAhKMumdKcaGa6O1yvtuTh4+yCWtoh8qPmkEC
RBMOW7UDIhoinawWpTBkGu9mqMOgN4DG691iwCfqdkr58nONTZPrpy9rVEPRjLiTGiVTzmGQFNbf
sf5JBSD1nYMEVMg/DJ8l/BhSDyzPVkfFzhY1HahBdxeXQfHM3ioraIvIn0jzTPycMUKMzUglc503
AN0cd2h1YW5QhQkp/tcW3NkUnijjBaq4XLCKk1MS9mKNtMlW1LBPjA3+kQ/29+A3RHPZKqOkDMnm
W409ET50jBZ3QMNaYSKsq9TW+47xWtmlPLmu46buHMwz7b7M7ow/1FG4vp/7f0kPPjnAI0HUG4g2
dUiNuOTk9BAT8wbFHjfjxTmAqc8nbhaWcdIOs3UYuz/CxVVU6xdTazyXrqeF7U0d6Lb+PO/3avHB
XUPdNT7zL6wC5TRe3sy6WHh10bipYyJeja1bpxNmwXb+aW4GSS9HHTp6rsB/VHdPrPbYNgvwIcSA
hE3BCPEh0KbBBCUeRfXKRRyf/tCJCMBGtiWCbtWkRBja8uQqtnZWwAxGOeZNZf+lqpwSe/fl/iVv
dff0HQCHTYTnyHTpV2tL/oDt4vMiFKhh7JKSgy3/YMOKZ0iA3RqWSrXA063eOIbFUjGk5TYRMbaq
DxhFk1YJZ6J9kNML1Y/X3nDHiehQKBsrWpOi+7xFXNEA0VZCQyA7irXiKnTKP86SW5VjQyKUIwwc
7IQUc0wqqzvqFzS38QEE4iudXFnOE5Ir4FzMKKIeY/7UrWCOe5IKVBXaikbNOTCsBVlInaECIk+O
RIDF4wMH9qEJOx5DPY2XAtUkuOOJn18CXVBTuChNI2VpWsoYDPd6NIHxzm1PJPJ5s2NDyCFdGd1o
1QJPKPNi2n92U/4hLVYR+Rcb992IcthamyVfEu9IGzlyBwvDUrTqvXjA/Y5y0/fHNJbx+QHxhrpd
E2kKbCg/MvUFlVTG//hmhO1ICniYYYrGdvJF9ovSetCwvysLfSpDJjUdb4a1ufnNahGR1nB10mJC
9A7SWeeDzJ2WHciE50TcD0XSiZEoQ2Y+aUc0d3HWm1TPErYBwvCTN3bO9mrmZHCmVg1u/KhLQ93E
F1SMrICe1nioEpvjJhFJCj7wapbHUeqp1NLz7HA8zY7tgWn0BWSD/ebfj469ybcvMIBvFdeqyMnm
m9zP+ktk/bbPnSNbmIobaw+CBqAZmTUa3Lquan5SQ+xsBHZWKZBuKy8bYvIs3iZVcu8eyARYbPlh
Xr+TZJtOjqzggExTRiTYkZ3h4lvHuTHo6eHbbjFTxQmDFoegStzOjJZhX/PJzgQbOjVYto9gqmig
TkQcQ5gWR6/nVaNoy8j2Rt0DxkLPEH2TErPqEyKIdGIak8EUqkT8PM60S5b2T4xRqKqfsGc7IUnK
js5p40ROfsJqt47eftscFuWOZVMqZZCHEzEVHit+b1yTacu1g9KQTj9tIk0W0J8VVXqNTj0VHygv
aOsplBh3UPW5GdnpM/kNqJEmUuEb2hMw+hzQVetG4tfNxX5e7ySLhvNt+a+7kUR2V7qLMIhDQHCn
9YadH5dTM3ePqyjxdAAHZf7tyGz3Z8XAJqbr3FQJnvOUPvdKADkUHYgPD+/H2Wdt1K64Of4eY0Xm
rUffXhapaQYug08U90WQAGV9T1f0oWC2gMRpom7PMMqvrZTegZt7DfvK3a6h4wQkD4ZvFwxBFRy6
vQeYJIWuBA2EUnrJWwReXn6I2fPVqgOdpn7e4Z42uEux2xsQWIOGUAEasnDzftVCxeshxnuSPTkS
W3vdh1FOVEzx+Wy43zTWTHlHAi9iNMiqHdquQ88latviooJMVdt7XUR1ikQvkYrphGfd1tYMJLg2
VFUh/IiwJbSbqeenpzFJ/2I+r2LSZKnVC7HZBPlqQUJfpRVqEYlt4MgJTZ9lw7TdX0Jfy4dK4PM+
FhaSuTQh5EhnUSAfRuvmvX6dxfpjw7dxxosBIYkLuUCkkTUSarZGjPFHmvLv1rVf0Iscq0w+xngb
2Lugcj3qp4RFVbMCvJH20J912BYOGYqInhDv3o9YH5DjJ4kelFEGuGBqN8qENmAwfRorFYHTsQSn
yq0/OHQ4tf10Ymiovj3f4yXu6Z2zRyhryuDWDvF6lE0f+mm7itOMXmpPNCZSswaC5Z/i+djYW32u
Qu6B+wRbn81axV/nZernUB08V/ZGJa3J2xoxKvGZsKmk3ZD5W6JCg5DgyyeYo7QB10tnKhkFBKb8
mt8c6cyY/opV5snOOdebMR2PTaqW51kamGeG1h+DX7ZipStuS04w49e0KgcRBBAgG3l8+NfC69sl
QoWDZ3L2VjOOftwbD+WMer85qzczyY+t7nGtBpYG3SWfrORe+JanIboZT8O5bwR5rpY7iONX5cAt
OXOYV9DwmdEc9GTFzTcVuTZ4jiubSWgphOHSOJwQrKZ9PM4ZLmvacSpZgMYT70e0iKNdv5QA5rp6
ysDGXIkLFNfLfAsbpCt4jzyUgFhkoN3t7fUc5ikwj6TSh79H3yjcpJFitLd1xQLsf+4zQsuGRqPp
Que7BXMzyxtX5dleeIYbScVzKHpkA2ITatkr5063xkMOyCf8ZGvoPBdj33YOA1fn5Kfzo29Ur2fW
zdeTEydDW/wJMbOTa6ITL6tILjKJ3g/EDLvNkp4GGTfkxqQuSQOQp4RIN+MWxXanGXQCV5ZR+5cN
XEv7Owv1O1Ii2d3oFo5KBH9/B9AHKLM0naW2/6bgqONI+QalOuyj5sgdzt8ugLB4mbj0597jbpkE
cHwdmEJnqHDh2D0dqiXuoSOZ0XSNsAp3ydghrK0y/b4Q1rI9ijVqfQeeiLE/9Icv0bsXmd2iSb7k
Q2TAAHFWu3rE71nFlxw+9ftD87DG18hP9loOyYY/YoZq3fYLwRze5uC4CJN8tcVV1TvmCxDMtgp7
kVUnYazwzv1KBj8S1mtRm2un0xr0Uk+y7/VaUjq2J0zOvfS09Ek5GY4qsZpBEK/8J45L3VlFTtOZ
g1yAtQFT+ePDY43aSVMyXs4Gsy6wXRquGcOcVDAZ6Fr7YvnjGX3GHcmo33cQwxxhNS1/1fZhjWrr
Y4kEpcY66GtNYhJGTWEmJmRSq5mIr/rsUs1AX7sBGW8j1EMsUNbgEoeqMcFuTp94x8J/h+nR3QUP
RbYom5HU6lUcsnOwQPTHSamVK/Phl4Vyoz4cHK8FcWDWYiGPt2JOk5QKv2TbjfvH5SvRdtUxzNl8
4FifBWNG36rlURJGbnLmsn9B5ShEQma5FuvizTxBpUtKcBNGagsXPxBm5Nw+hNkC3dvHTxYOXlT4
zYcBd/wnP9gtKd3F0+cDIwLAVA//Rm6exIDBJejVc4eb/1XAEnKxup+JdbH+aLvqmEKIRgchAHRD
m3D0KHkfXByR+GhZQrrXOJ2NpyUtxqddbA2QIzO98CbDrig3fHSvj5Tt5ASSkSXUHYNundFou8tF
/ov5SbWqfaf5N7ARpkIpkswQeoh3dTmkEzgy8TDmJrmb7EZie/Sv3KgEbecBgT1lXOdwqJqkvdY2
fa5FT0aid1RLp4b2lhH2i7CTv9S8PIQeTzDEbcWHa36XcclpfUoCSz659FFbwDLyynPkU2Y7TR3s
fGQ4Dr0fALdwCGAmZtTgB9s+TqAO52INpiFVB5W68cmoQDopYU1MLEe8aAglgFqBQho4Hc9RcG/v
yuPnud3mbkq4mMw7sEXpzJ79N6JfVQa3EB09paQinbFTyigMIvnPu9IgGg+HZcwZhwHCwUJ24uBQ
4LrthDeNXenqYmHot0IXvsRQRqoIIerE7Is0AfnYZ8cp43q2jqe1KxdusYrtAFyLaAuW7y6u245R
y1kFloFC/zooQCBXVYVCAQuHQVdc3J6JgNFk25ddnq0OcdWigNTslItKPhVgTqrfJb5nKq92YtwQ
HV7odGwEQ9uD3WMgmu48sjc9Ao4+0p+wHIjAopojsXrlx8s5RJnQ0VskicIcZbB7jOZXu/8AzzP9
AaMrimP9Jpyy2GDc843ZrI0qIEQuH31FKpR6uILt4d4PIKkkhY1xzn5GuDDko59evmUXNUwZhCUg
Y3FTMPFF6e2191kMrb6MBvIJeU6aR1Wc210gBuoWM9T8qHkGd/9nXd8uM1r/RHPC4Yv7n0z1+K35
qmIDhT/f0Dd+E+d04XzJEF5I2Q1PUqsEzruBFPr7C8SGwyk1E8MWiJLsBSiJ7AsOrFM3i6k4YN4Y
K32goqervw2NyuSsFk2sGaVFDIDlTe5oXjVu/JYA6/ItTGi+YTgjThhXxLJWvuIdxBtvb21FlXV0
PwgyAkKyZH/PEjiVTVkiAgjABzYvDDCHp1GjhtWPG38GLNA69UR3heG25QjgH7kunjPG6SQLO7b1
Bnf8ia8OmcRVMBo5lUl3gjJ5QLk06crWiin4MBJTq8vvBPUdwusiliMwU5WOSqAxAaVow7Gkzbf8
WJoMUs0vGpGjdysPMCVV5ektfQYwVTwKpqnXcCoDbBT0SSYRTTw6RkmYmWEh4/ivHcnJ1QuFKXT7
uDUc3PDeEwubh+/Wyq84Dl7HO60CiGX2AczAnnh+HHHuqKi8ROMrCn09+dPQ1usY99rCXSLDKZcv
quCARC+AS8nQARilQFlCMBci+3J7A5FkwYUD+uEH6cPGaanY+0QOZrsBRNcCtk6GqB5uKPHTBO8y
W8AVJx+XNGAKlb5Q4Hc1GCr4owNtWg/pfbNRrYgDd4lV7gCXzsTLhXe7LUW33wtFEOms7Kc9fIa2
2av6Lp+/rPFrhru66u346C6edMtwMS7s1eAJ7blGYZ9JSntZxy9YYCOCZ3gffTdZzvtLaVjAy1+r
SmryVLszU95wV5qoMLuyzuNOqrlqQ7OsvEQCasCI3VswVxLf7rg8+XlfuO+/ymIjuQxfBAfNXSF5
ii19uloPSKu0BWpMN4nXBRuW01KCuArqr0kXVb7ZwDAjF+ByMnNO65R02HbKiFRdLy6YiRKDcdmo
+rxSVdEP6OvY1QDkPR4Y7PBat1Ty11wjx5dzFvPpmyvpEDtpUHDLeyh/0lBydrR5X9H9tdA2mG1z
Fxt+e899aj1gqTKxaQ0JLyfW+Mshaj22j5fQVH5J12J9vbj2/EmhFB1mJMdhKrbquYfc4G+DBZpd
VKSOLBdww/3k6XoBJf1vDAW7xYyVwRCgiH+98O1M++EIhju3mGFsLOwCfeRW+wdkcdvqQThrzIJX
PdFr/P5MWPIcw2VT8jG1kRR2DoBnm4C10/e4dSeqAZOudAK/pbJQ+M0nB9wXj+9PJhHnZKaU1LJW
oGiALnypu/GlPe3m8UxaRgoqL1DtzBBJ+3z1h+iEvgsXAbaiHbAkZmstnej9RXdo386zytdmXM9c
UUfloaoEL1j9V3q7sJlS4BXgwpvm2odqfP3wwLV+liRx9DtiyqxvLU97yd2s+AZNq+pGdxffwvDX
HnpDROP7AstQuxE7mlldzd3+j20W9kxOM+d2FMMWFrnKAtWJKeuKyni7DMBl8eClNYg1nff0m6VN
mTldXwUGwC4c6D11sGqT6GuLwIpBtSAb6e7a187ONZaDqMzrIFhx7Y/Zv12TzxMhbs0wsNNuRjnz
2cBfRAnNXwFXnBf9LvWZDdlMcdwv+EKoyGMX1bx4w4GNJp4MY//lSHJroqARTnXUVomJEtHHDaUc
7gRQHuDy4XOkVrAeNvHOSxg+OTNGvGuYPjhJHNrGK1sxBNueDZ1E3WcAOhGtk9qeF9wstwqpmWGX
kmR8W1Ju9ddYjVAA47yHLoruyt3eRDDz1JLx1q3IyoH7fUud+GsVfNvvFW15LL7CSje6RE+gKKBS
c/8bVUJ01vHJ21hN1UmJwHFqobR0O8iD82/YsttJIwIochQeZIgZkualpAPNlbgUJ0B91FqioL3t
wtXjSx2IVOaoUOlYFFRsI1LxKWRhbmZpL026lU4e5HR601bWr/yYx2GSuhl5nroi2o8EjBcXFMaV
G0rhkulBq/d8xLCCLfk4nHBR0mRryRGmerix7FhLSv2ezHmyY7FeGulNMTwueqPCca3R6Us4XVnD
mWuG68IR1EFKezYZ6uOwAZXnEy7J2DSllBAmHe4sYmk1OL1Iyt5D3SyX61AU+DMXLzyhIobaY5VC
OtoYMjMMA9P8oW21EdLndK+7KL1CWKRw3jSrw1dAWNurAdME9zq+9bBN3cZPdt0M2egmTOJb34bo
2qB6awVa/WkUTgeGU0WkbmYlys8Oww+Di3oApvmUIoxk99V/sUZV7K8G/1pogpS0pr/g4W7PAPEp
Hbg2qiRd94QSo/SZhFgKP7RElR8vUHFhmYBSRkGSKUDtyg/u+VKPi16f0O7sRVipfoiG7czZofea
/25X1kihe4FpneFuIOtQx6P2SEJfbRXwLlr17v6+osn5CZCLmgGjBIk4GAFzJZWs5CGoeFjooKSu
rZfciUKBj5iv7+VulHyoLbeigVb5zFYX2pUIQxIsD0ujCg52usJ1tI1CwCtcTeulf7aQy5s3q2l1
aoAa+Wf8mUzIMAHsU0BZvf3SRnwjOlQYbH/Ul00vBYAsbmzO3kIR0H0unyGSA9YcAD2bbmqs7Ik4
Ka7SKrxD1tPsg/g6CEz2dGkDBJkzLPcDursMOzl0vz8UxZYcZI6XoqbTOacr1S/vTuR+gcWk04Kv
dAp3jasgv0ftCgBy7EeVQ1F1hCVqNY5GDazLXH9O+3g809qiu7vhr/cAb3tw5CvXku6MT0P26GJp
5GczwtnrGa5lMWd9lBJQCuHbM+p1OqBTp3oQVqf+zF5jAsNgOP4dub+nITB4hg8v7oJK7E3zLhFN
5YMeMerDDVBUSyqadN0WMrXmeyfbInXztoJFAMe7pddD/ywFWqA019KLeA0PPGedyPEexOq0SCHZ
DR+S+23ZvdUf5nXKwyA57j3H+uWmbFLRPHY6GLkawt/v9M4leF3EWDYBrLWuFwodiSamKuJwieQl
L4eWskFqTBqcGTlJ+eXcHxfBE/sp00NsGcmWFc490JjYwKuyYjNENqecwz3Kcaf13qtWFjESNRvu
LWN5wU3WFuBc/HXOJeFgxa4yAWaj2mrVRU/+asxAWbt0qAZ6u6TwK5KzD+1NqES+biCEMQUFOZHm
AEa/ovynHkz9JdUqnrnl6Bz2C9irgj0FPtnF+pAlMSHyPIqa3/q+jI7lMWwWZDKqXt3FHOlSWvhi
4k+NGAH2UN6xyXCk2dtRPYFmi7V5dRp8R+BIZuN+Oqa/svRvgPvImMu5LQvsQDWQ6IrQScHbQLjF
XqvHqMhmY1rnIISomhGChu8O323UDpAb1+MolO6cbrbbmajXe2zNV8XVVgmRapNCN0wBNaqrQrCY
GFFi+TiKVe0R7I1wE+9g4zRREOEMYQbQMtt+Z6QvQAnN4cvJCKKxU8B6b8va8uihAUcqEQ46Po2z
NIz1LangeEHjO266Naia3OqRufauIPXpGuWMUOvYRjKzZFptlOlJYlkyTcvcuGHatSxdkey35CB8
vcpnj3PgSPNfID67OX8VxRRpNv+kJeDehjSZqR6Man6d2JnQAAbwtRzU4vsUA0svCHfOzZkaKi3P
C/Blo+fYfRy0s2o/O8GeiMFLrOjEOKYP6dr08Ecgj3vdXVCellXQsNvoiL9XBvnp9rF/mQmyAPRT
2WLM4z5GVglorILBqb46Ow1vEogpTaiScsdfE8TMM/vceBFo3aVdFQJaSsrb+gCY1ww8I+bUNgCe
UBBQXnjR7Dm6+Zq/+3RhnMi6RvdA3Xk/RE9Dsei5rTOlrehJCWfEP5h2Gs7H5g/DkkdfSXZO10oP
FjXwMfTvNeTl0nbEFbPGARzhpyJycz+nMb42Md6BI6q3mmVQPSi98LvKj9h8ydEpRKrRjURQUHPs
Bwa93BD9h9cNSRq4QWd1Gb3Zxu3vgp6KNPaCZsS5SsnDwP3Zu++m9idPTBKGKn5p6Moo+GNXBWOT
jCuUj0cjdl5z6xhw4LaEHVq47PhzFANDTAR6Qdq/lvhDllqzLNHPtAGBdQ8EAdb7LvAeTBO26OyX
KSYyAGTo9kS5p2w47y0JEVxFxHeLlV2XKKRQjLbcFyuGpKivjKGUFFIttuT+1OmKgnTD/rgPlYDL
KMRBV5yEhwRiX/ItZRRJfu2ftCwl0gBgxIeNVSw7e9JEr/gRMKFVcTZqx+avxgwdaXl1eujmfWn4
IYHpShr/EwUeOWvSozcqUAEYQnnE3yq5qiO6qvw/NbagBeRYFR8TgVcWKoL1PxfQNABk10h5CNZx
0/44v6OgK9qkVTBKkco9ouqSDUvqb/6h2c5txMF2Ml5se7ejf5FTcKy+pfrM3MWTHU5QjEbTWs9o
m0VRZfqc9tQ23lBuW6hh8DYsicd87mZmqzjHXyzeiGPovba/+rQLoodLqFEdHRU63kDIfMWREGFD
JvB6EthtWkZHGW1R9nsSGcb2juEtYMktMiERCrn6Sr02azbvBCZSB5pN91AT/m05IllGqwv73UjE
IVKYwsBwaR4zvrIJMK/ITGmycqyoO8nUQvrMwlGIRXZ4t7awzXCRyReTOsW4qHhnCZcyw0Sxaihv
RvD9v9oHlnqPKX2dcS7Y+howl6L+LFurKjtXDPsfP4IS+/VHNRJK80avZb+c44BqFoQcUUHCzigs
sfTC3TFeqglzl5Xo+EpcIl+cs60Yj/nY9xXkkPRrrzWUea5QxZ7hA0tE9lPjJWpxDA6a/wv+cEpl
CXoK5sTbHtNP0VCAlxmsvC8GmMPdB9eD+U6t8RM9ALM4ywvh+JGRAWYDc2bQ3WUV9LFhdNP31Kvo
RMHyz7O+dwT6CwmMTA0RxI1if6RLRk/cAhoOzHdoNJt6rjXii4yxAfDORLZH9UK7OL8lktwDZj9T
YKrX71Qaw5vu49Q5RwkKzExxvX/2LlrmhPsYCzotMW/UI1YxaEYh/e+qVEuQxMYTKEQjexVqzeam
wRR4sGvkJp220plmiFens/ibgExpXuq7ooHzFNU/tK8GbWqoZkfQoyMTwqtRNOX6naB4d1iM1kt/
mTO0eDNiEmkHx9lD9MR4X+Urq6ejfLg8rfsQWV4hWcGAwrU6KJ9cK8rVwXdlghb2k9F2zrk7lwMg
1xxQQzLJuyzNG5vYSIU6LWTT5AMgHLm0mGcE5nppziNgaRGMSGuWhTVp8jeryewmGf2aXiqLj+ZN
oT4zupWO9VYal0LbVN3KuVWGBC21RgDqTaEQTKceKumyXmbWr5edIfp/G1MxhUOFoTkfSL6GM+kg
UpCip/ge/eU3lFjBAFjyh32rHXdJkTvcUksXjz924NF1fXxPgNqNk7d9bkMUiOL8f+jgK2dg9ZNI
qpiPJsMzUKF8mdu6GML7v9JyMjpEUviQYaP7L5D8yyYjb1r3azvZThaBo6tdeZAW68Vo0YsSQO+C
IYnaK8QAf90mPy065+1XnMASdLe3IJ4x1XiLXuIavqlfb3ywSm8+AHNWDrIqf6fqIqdd/ISFFxsT
+Vy1nQ9i77eRMqPCh+dgul5OQRnDda8HMH8C1Y3RDybTYVj0S2AwE7JTWLTnT5HSYW1k5Fw4ncyb
dV9mhWjNMCOS2N2Eu++E+kzjkyAMu7ucy6djCRYWTJSM8cbaLjZcjg7w5yLjBz6pFCo70v6YaKKI
Asoi6+Vyl0uE8wYurlIfs4oV6mQ2vlcWV3H5VUw6SgY/vzFe6wC5sHN6UCljCBoyO895kLzzHLQc
Ym6vlN2mEn85FYhJ2aONqVM2GyiuDKrAqYxvpWayNkGFkAZcchqyVokN/UoR4B0kUj+Djlrmkq3k
vi540SmMhAOoBEcBq6zn2XUxMmvIyzT8zNH4wdvWcmlvuImZoEYwCj5d7ZNGi8hATu2q3ncc1DgX
zy9svEuWXA9YCNJPT/Eg7kEA2Km3k98lKL4lHREq+TSW2cjlIABpeU8gOFZiktahTQzUeMdyEVPf
/LcKcUmaklVp+v6gyDvPEt7nOhhQvfoiPO0Zzd3foaeSe9Dhw7u8sm+DMwwBgkS3AOuTphoIqqmL
vKAGNdXV3wSGELGiX/5LXbC4Un12ieN162y9KVa4lppYdZ0fx4ukzw9J0/zFpP37t+J/PPbIsexP
7Z2I7r9m0Gi2wD1zheH/GULNNV0i9AWy2vJFAD3A7w4ffmp2ARCD2gxdxhDRg94CzE8tGKBBZ1bQ
kwJYHRHEouUwOqatL4PwG22m1UWGdNKAyF+quoUisU9EcuGiMjr2K43IoGjUbDep0HVrNLT7lcOb
RtFHILGfuFsVYmBz3te+z/eNelqomehi5b9oPOxdlJ6M+2i5kBWcO1NZPP/AiAiq7clvzxqTb8Y2
eoJvmwXimV0LVcMfSWbmcJTYXNRgw/LsXntVr+LGzZbm7whmAOXROH222L7snnDIYw2ubbdFZBk2
cG4y6emulCcx2jGt6qR5P2XFgV/ti9nSfahnubH8clMKmPXT4HuFAnADE/eRkJyCb7Q3aqfyp8hJ
WYyDtVTgRGsO3sFx9go9vWYo684LAgPZyABvdsxAB/Cah1bN+AwNFP1/PaczfKxvMZ4A0O/5z9HL
zePdIAElDAEf4EL/0JgeKp9L6ov7kyKJe1M596ySl//IaLXfSrDfGxeqdp4FMHjRFTiTPYK5cPC/
HaO0LkF4Lul3cskR5SvdtHoFSqN5RJ6vn/u+isc9xPLePTeaQ7IUDAqo/T82ASN5iZMUGj8WmsZ/
wgpXRsC0n7/LEwGNN2pTbty6yFy2JtTgO9VFPMCqhSf9iq9xo3d5UoYj5RytO1SpxFrN5+zBEYAG
A9gx+nDgxLzO3koBCon9RpX70QSjeRbw7ZtS/NFSCbWYhQT7l54ezTMxTUswtOmn2igsyV3p2DLp
h3SQfiQxK2tzhzOHPilhdRYvMJshw0ym0j6+/cg0jsJOiDTUZjz0gPHFZs7m7NFWjtoNAEbaT8nm
OgzAkR5aydJa4sRJteJ7/1HmBTln7JtFQqbeMXvRh4h6y/qzY79Vo+OIsj2cBb+g+e/1YV38YYu3
JWxRLsVU7z9mK1ykZ4np5FtWCr/b3jwZdiyKoC9zNIXcLv+54auejJPbt2BjlR6UKQSoQHo9MeJK
afkuONiqRTiS8c5R4mVRz3k072CtStjSM7zPIxF2Ru95kiD1FKXmcJWliImGUyH7HnrK7QXIuxJe
9cgf/k1c+H0Q5biR+vG2aexexdrt579zPrDUCtFMN/GDpGdWS3ve2kFqxM38HZEk+RdKZJkj5dSs
LiaBO/CkNyXj9Dya7nPqpoGS/3/R+NeuiUXjM+icU+JoZDoPttK+0DKQQfbTbflAdAh/RTs330dW
oORpNI29URA3BUT7P4G24BcysM/cInmPKgEYfoMvdlzdgVHKAG8N2CmfAd/PeTYr7dlieiMYVgcF
S54ZNFOSqyhX+pnMrd1gatiBuW+yU/FWZL3ERL9EpXRkAVgDHZd+dID3LQhvUP9cjFArWqZj6veX
LkzD5dg7Zxo495yxd9wELZcBPfbLO5Q2+lHtiVnHk+lxfTXq+PyrVwCIn0rd5SHeAmmQAiGWuOSv
83ik1gDvh5BxgxzFEyJHwmv6qgMghjx2LvNnR87XavsFiqVRtFxifYNsEgZkAzxRFBnwGvWU4tN6
ZiqJvmoOr/GQjUX2Wut1dODyLw0AjUMKNB9EkxkTp1oI0RAddEl2bqz6Wnh5xVKo/DtuANNn4uwc
dL0rerbcwY/d/Ia64wfc79Rv4/XIFi3OtzkZUS8lJZj05IujbuEq5uJPI+l3KyejsqHHL5PkcCvH
+vZWVoREmgIR3/nkfljJ18lUxb2UEyyazRWdqJiKSbw5aguhxYvVmhgkkaRl0xA4TRhLoSkF0BK6
PY8dIy1zDQ1UVPeKCGkuFeXXKhEnZfbz3d/ZTwd0ctJqkZodXB6xMN14qt2MtHiAsanj3YBntTtw
S4MPCgz/lCmtT4LalPpoq0ZGo0q9A9x7iO9pYLHhTx3Aobp3j8k4yZ3z0985n0Fa7ZCrccIPe19I
qDUAgqcToptPtpKbYIRKQfKraxmjwdDd4GTYYhEZsL8dC/f+D1NO2oyKSosnvYRcTr4ZxzttUNqY
LbAFtdIIZxIn3eRVn7GOKAeapssTCs5GevZqY1JiFMygD7B5jWPos1rKX+2qqNdgsFbJKDbB45zH
M3xWnS/cjS4pK0POyBgB65361Th3q9ERdeLpeumUZ6i+ocfbEYPTGEWlZGKkGhkurF16UJ/vm7xw
V2SqpdDmuVZiG3n5GJp5uZp5pmXyL3H3PtPH55qkiTVRVNRcH98zWMkZibjI+vgphmkk6mF/5V00
6yqE3bSxorCTuZdcWZOdakZDnIxCETPMOcAk8Bt58iPOKQ2eqRWVeXGwBKA6G39mAm4YS8pK7QWr
C5BrmTeFM/s1HVzD8cGUjZl3Xosnv83AM/6gAzJtdjOdgRzPxTqlBGnpW7JVOgaK2vGaiW97GZfj
OFOmZf7VHl5q9c94lo/867beEchuHwd2c1SbltDK7x58LWvFUsYLZ6eXaRKRlW7oSsUNVjUGvJbF
iLMTBl4D/dXFtO32+LyMyypBtgQ34ARKZf9DNusVcUkIuH4VfBJFVPJ5/PUiqSU8rpgQkS63CcBh
ZudJudFiBBW0OId49bd1320PhgTag/9eZwVEgyvH73MQME8B2BdXDoS8klUh1GqsVPF1a5SQTsTd
pPhD/+53gf5lCrXovs6b3zMwTkaDNcu8YXvV9KpHlnjDRdtI0cnNRf3s6pHOKB1wveMKaIwsxU4p
Sw3IvoyPtM9O620b0RoTIPppzD74aJrwbKP9GPiPhECqYay9p8q/tDh7MFqs8nLpsz2YBx/MXgnE
ik7igZTPdvyNjpvPMt7rx8Z2USvaxiuOn44AurFSvjRINgk6eJC93wlDEVhhR4Z28L9Bu5lse3CA
CS1rEp5JVIrs7VtyVPO/2UNn4uoeu90V6+KN/3HGhl0X3YNXzCkwSlnr106rq0ZtOvpEs4iBczSG
A2IDBQjHrPfK5FzUC5qJUEApfGyL1xMGEjskN8+4qAJsOko4/IwqA0gEitLB6s6ajwHCh7LrCJgN
vb2o07/RFkG2k4jgkjixkf1QprBpF5/HlVuMbLReN9ddjwQPA2QPiyMoIO1e8flHlxFxkbHrjvAR
l2Zz0RNEfvBGKPrrWRGNXsfMC4m788qO2kbyDfUWiUlzb/fpcR95ZbGel9edISPl3Ofjjep1/Hlk
X4R+Iw0JUu+glA0RSVOcU/vOI9NyKFdON42LbXfLJfxqvJ06hghKsoxj/1QgOHbNwe5uHKYa7b3J
uHreBrRVkMsc2uaTPFSqXyWybUz0dU5xIU/n4d4WqxbDTfPvDIDyzMxXH1vxJggx3tZqhb5O4BUJ
89A7X8+BOgDIKOtjQS2raKruO4VpXYaabpkzwcc49wsVMrRQKihq0CHoLekGLk6YRM2ynf4mob7/
khhT9gInHffWucg2PQDVoa306e1rqc7fei/2aj77pUpCCji2/xBsHqhUos+nu2zBAXxBYPXi1VW0
p8rfgH237Z3l76k0AOssLGNCrCMkvqOxlZfBWDyUe8VTJDWa9bhZaskxlysrDnvq60qKd5v1HhtJ
s1naJZjUpSIknSqaBqq+LWEH47OKN0rWmuLpAtSHHHo4x7UgLuRuDfD49Nv3SsnaY+wMM7p6myC2
w6eFFFsKYjvM2e/jK+5pqHRrrLn2tSFfP57KJMBYoQ5J1IfS5cW54TCNMppzuNwq1Xq4IdflVye1
MZc4O8eI57NRhThOBDX0OL0RuRmB8yqkiYCrImm0xC1bLOMFz2DaY1QVO07szIEAnBHAInCJK/77
RdlrdwFRG1xITTxgKjsoZdL5Cd7q7YjtRd4wetvfUeXaNWbRYA8a6Iiy1PvDrtPHjAXxbj3d3eFK
gRYRUK8/BoUTgzaSEeZrDbK2PMHwssfznXbCoGqWiZD6cPvnI82+PfgDxPazy5Fxj70EAv2FllTW
oYQtwYWGLg6Gyyv4Y0YforWUVkz7LSXiBw/kieWlT8069OUU2TltEX0iUtXKcCJZg+rLFd9zMGAG
GzQg/EKiPAvFpGQAbR4oq3MLqvfdREZzgxaUvSK/qKVp7ZL+neFaJweGA70r9cZuQlxkLNQ0cKaw
B0oSroebwMWRgQ2dkPxwx/4IQyockFFX2EgSKiQFP+462YQSYGAd0KL19lvShznegFdZJ7/cFu9r
Sj0LJ7z7VJzx2N7pWELFEMYiI0DZeKniABlh+e4Wexv6bD8JGOGDd3g/Om90znZCtcKSEQOehEpe
cPNJP1+DPQE9Ri+I4OrplimERbo6Ii93EpkwsGnFulB/Kd3JbdJAzlOQlvTltqRfk0vjwUUYgebN
0Q3N8YziHUPma1zmTnIh08FIxMz7mqEU76TU2RsHl2sjbgAif688KXqsknEb5bLrpczd9RA5qmOq
NKdW6ylokMCYgC/WJYwJq+PlBS26H4qCMNheCogmpHFTiIkQrBaysl2Ca0X7e/zA41MH94IGthEK
TWTjoRqfZfP6sOJZXhFh162pGTt8fGmwupEdvpqWRrgWrhxh3PObVQ7p03SUhw4zBZuwuWuKPFEo
P4BevMbBuGKV9yL+vA7qD8RUIzoXB/fX2mg6FjyrtdzIP1o3MC1Uqa4zOAO9960wnALlBzhYPDGY
hI+TI4QRABi0ylb9WXjEyFmYM3OqbZC2xhCSGUSkNso88A/ANOE6cpkc33IvYYRY+M+4vlpyK58y
fXzB8AZt0UTLN/UV9ocww5bZDt6WbXEOG97rhajrxnzehFTFGHRYv8Wn1cW1vSlRn7QBkCMVb9ZX
BM42eSKecJ37POptcTASvRXm4D7M0kv9FH5B2oBBOtDrl9SV0mRpMw5hQX86gtxkRayqdPVTtMrK
UQSGsN7QKhhofVl1ffl8/ynW8qFdvr9grz5hpeH9TElS7zfb1nALtFsl3UMJ3MByyPU6UFjSr9y9
IlZVYgeQlZIQFJriPGfUL0KqB0NnwQjcyU24ARgDbufQWRcfyDb5QvfGDM3K2YCoiHOF0T5R0NiG
WSfL8wjaeWKDy+7elJ0ASqFdSYTmSEAnmw6Sy8jugA1BMkHUupP9T+Algm33hBfiZb6kWY0Ff1tD
7BjMkMuDGMhjrXfrqicAi8I6OoMbv4iMzAFBx1eCn/IIlYZqD+WkoBYlwMBAGoZIsmLmDRfQITmm
nvUV24srwBWe2UXnUgQQlWjaYOcFNAkUZ/J9MCwx5Q8CNi4CKh5ovhYV6oQ97wYY0xhZAKW9XbpM
WkZlUGAB/zav/fFOWPxi9+m7elnGahvZKPY1pzpoDNKU29AdNyyAhAu8brcLfVJgRK2cGN8VCJgA
mImYjoWtsOqMh68GUBCkonC+yAwWdDYzHGC3b4N8bf5PF0OZSJy9rv0LhE8H65dz4f4VZaMF+6Ye
gzW9nWfO724UBD/ILEOkg92u442iICHnu0gcfgreByd0M0hacdnz9uVwyC6jO9IlOVUtLCTFj6ji
JgmE4/Aa8wS49M5FHPAuO3Mi6AR72hOzfew4K9aeP3CXVdQ73Ajq3K6Rk0OdtJLQHLUi7360Brim
PU1/A6CpvIUuuA47x9Wx0W+hzfOANy3np4ko9RXYIn5YzCWgbg9wX6FN1ei8bUupfC78lqvsDfaJ
RkBT1CiZJ1vn6qPpoWWIHtxEAOczFss3KtI0qRFdUq49W532K/E54kEcTjkp8IK056ay+tPJQeMj
SBre7yfKSA0XSE8pIMEsSXytslPCrD7gq/B7e4Q6Nfx0MDLdhnB6EKwHD+x+CiG4WyYrKLyxcj5F
Ty+6EGJ/ZJ0ZsPsUyBDmF+vF349dC5jgfqTkAvjQ0AD/hVU8+sK1CY5GQwwwSJtY3GprwpA6jlMZ
I9UFObN12OaYD4QGjmYDYqGV49p64Q5Et/iEZ9q+MYbbdaKkL1s7FofSQrTSnSlFrW9haaDVwgxc
036h/OZTMuc8rGft+SF0G7ZOS3g4yhga+QKVhOoh2tOuYRyDZdOTjfKbNFox++1tJzVn+44/xHES
x+GpZ4htr3MDRYv1mGM6bPXfngnzxOGM6N+I5lUru79IyArYmPY+qky7rRGXnuA9bV/m0v279UEX
2hfWFrggbFrKWLBMcajV8vX42bPwcR4gAGmP1tkMCYU8NZfBI83Td0oWzTo1IGoDBZXYqkICHwM8
ySM8RHvh+O1wGZ2xSycdYktAmeEq1yeOb/4cmaCcbeKlXXyBu8xzCXYKMo91/nOLJL4sp+2LMlcx
pciV/GLCzdaO0XyHjhGnEfGsLyh6qG5uKz0XkRz7gkFbaFfaChoK1t3PRZZ7Tg4NEe6LefukCA0e
Y4R+d+WUK7MPxE3Fx0dFrEQtQ+GrZjBf5R5PPMarIDvw6JCCNot3/34If4USRS4dCKdvCTHOvZfA
R3bl+9/qL4OYRac5THkPpRJ6x8UK47HXMhKzYxzfpn2Yv1N1RO/hJQ3cwYRqB13wS39vCc2F2O+I
67W62jPsh8DEQbjsKAFFmK+ErNB76wFmBfjMsrsh09YDW6K2yfH4fOKzBpeCCdHLUeNxThczirtT
OtZZE/5RcE6xmg/NkoGbineQvDl510g+mBTwzl+6rU4Nzs9Ez1misMSsF+t8SpNpUDtcJcPzMqMC
N/XFkEtHWyyO6RRdc4Rtm83nkITKilxyPIfLZf3b6AKxvaI7nsqRHFeYdjz6rb7LYv7PqEJIpHbs
XqvxfTg9OakOFqMq4668GWL6VrSeEXgLdhfRi+7UwOg276H0n1XhGmZb774vSYyPRg5L/nasy/nm
wCJDtEY244jZBdjNXBGp9/K5DZ6GV2EKaFzqznqc1xSmU7BDInOapNPX2GEfCkDQT6yjTkA7ZWyz
dEqTSqRVvNWHCgdcQer1r9L8TPpiVvczeaA+D9CPCF4D/TzNItLzqt8J3Dgb8PFwoLILGuuifSve
wvpKdy++1u/dteFs9+yFJ64Zk7YZQF/uRZtYkT0OAVD10vkHgHr2hIUkSV+7lPnEPoU6JPk0aiGZ
iSNa8/rX7m5WIf4KszXoiQ/8lA5LhGWTmTdaEaA2iuuTJxIeG7XsV1ddo2dqf0QbK8ssCWXnzM+V
UK7+JvBmd6XkSPHXYLtVG/K5D/IpheYdO/YNv+QFti824d7VFmMZ/Kb0PqWQVZFKvlPkncNQRUR7
hTO1IGvwNZBF1AKF5KZbFCcak/cLGUMwf95wMjn/SdYV3FQQ1wyWbZcgnxEATr3FFAk44lqdr5P2
WmIcM4ChMLrVxaAHftfzco7PvRBZQNlJWw6DQUjEvlUFtRIjxJezBkvb3tk3gP246eqXw8tAsWPN
W5W/SmLjuBX2pysrmeNeQV8EDkGeFuqK9otb6GutLMywegCgLHpBIScqE3HGZ+cA0r5Cb3KHJWUo
cZERUPNbpTSxcXOHssNNJTLz8SVf7J95vkCeTvVLR+RPxiaYxg/vt7e4rgddvi+VwhIzT3Kil+h6
DO5cJIoclkQfkX5v1GltQL4zifOAuwej0YY5fSuRdajggNlmur1IJJCYIqqI8NFC5YuqufIhCcfz
PoipfKFtJI4PiHGgX/IOOrVpC144ZD/EHghPrIzVYgoHy9AQwXJVexQQPGX7ms05rMZeoDaiLebc
pSy0CjKi0CMa3Evqer/ZlEtcqMVd9jAYo0jwCWof4IPt0OZ5MJpyjXQ9QXLt+inunwIffMHYlyK/
f1if003wFHLzzlPvkOD0g40OL16sb0RD/zcGjoH9w24dF91eHsVflb6zMMEwiXUCOI6D44PYXIjf
OHQkZ8ybKHQGeCEa9R3LSafReJCh5rkd1UIuceszbQe3d1SgpPs+tPNOSlWmdKkfWP71kgcI32xz
aslNd7MMw8Tx5Si+OCQxVLl+5SCOUdte4MCRjMMYik1p5MMB6a1ub5fuVBGuw4P9Vhoe4nI9b95p
j3SQPGe2hTVfuMOBZsYdUckc9bPTh7qCMb6BV8RHCs8iA80a/lr2SMETragM8LxXISRP2RqtgObp
eF97v3Jd/VN+hiMaaI1bg5/16EGsticvEvUIIdKTJA8OHVRjd5j5pL1ZsmioXnL47CvuF0m94N7X
wU6i5+q+ZeSG+CEeeGjMrqLAyak8oGXE2+V158b4i0affHVdXGiaFaMT5/+5LFIIX4lHAQgEIYbi
UU1t6wF3zP747Rgofo+5CXtPLgbapdOlhP51UDPrTc6DFwkEHtrAXr0OJOScPqlrdTRoEFRN+6WN
Z8qLAkKm2RIEkhPKvCr6FQ5X3aRBoB+J5D1qmod2UL6eH6AzI5UgyTT/2ytklEieNx5zndWGI24q
hqFpgwHCNksCL+137a2dmji6r6f9thrAk+/DkYDza5ezeY0Z1XOCLdoYaBTmlrm3yjrmwYxQD70S
hkVWTh3R+/mkkm308ueJsstRJRkuKKJAjMsyK3vsz65eC2uDRfwnGAbuo1iBr8AsutIxhvlqU4bO
Af/C1yDY7lTF83zPWvInW8osCYecSijYrXa3vwT/EcwrfubKdrbMYjzHZdjxdpxPz886yduCmVb5
zPrxiHilqVgXT3EK1mPN5Fey6lI0eettZtR6Ty3iYfROc/6iT5xmwRmGMNBP1GyKFmjEY+wqUmN1
bxMRVtsj6qKFCrGCYa28A9k27f8oeQ68MuNROkbbBJ09fb50RYYuY9ERz9GdCdNLTjECLQJyj13q
vFaH3kpoaYcYF/cnECkObOoBAOoHCMHaAwOpCIwknwsKsFy1I2msAvhrJ1PxaLn8nyCeENWtEULN
wy2fBn7Sj4yedSyr4RTFqkZJ1v7+yIk6e3M4RuRlZ0jkN7QLaXQyVFe//5PbCx2vYrjM3B8Twy4z
r9gToTAsk3ZmapMe08BSpiqv+EeZ2NaU/uNxiFEjogYG9GbssZNhkAWnSPBoJ8nm6UCtUVVtyQBQ
QEoR+1xRFNP683cVuBdfCjhaly0ox5Nlk2dygEIWTFJxSzvZndRiZCKUSFUckNmGtupuC5T4pJy0
M8PKYkcptRMxpKSeZ0GL+6oqUzMvWmNPvy3f+VGCJNPK30WmqAZ2GvKwZ9CyKQySUr2yD6MncF/a
zJHEyugs2k3Br1KG9hgAbyV+I2VCJPPHbdo1fWjZEID48cvNSLhn62ptAg2VYBSTynEoHsuT0iIR
2yveDZx6BUZ9Asw+4mJHylatjqIea9XuSidnjrwUUpe9wyl0abBUtkYnYRyePJp/3s2XktEEdp42
2UKV4R0HVC70S2wt5hX7eQ4ffYqVQXNsmFPymsfXIzcyPS0OJxH3LlwfDY2pkpfjTF1Wfyh8A59A
B4KrYgKr30KVhAJaT6PAf/o+t9yPYe+J/AtZirOfMkU5x6qk2+h6BiFnNRCZ2ULg2DLGS7+eJoM0
sK+CwZsLOfq57/4dY34CqPOeSCR543VZ4PLdomyXEkYr3M5z6MlJ0XuY8cj3GgSAMaKK7MB+mEkB
lOEvnOn+CiB1+/Ius7H7l+I3olN56fd8nVSDsi5AWGdz+MWSp9aQGN9e3Mw9YLFybmjx9fdwGzIn
qLU56kVDz75ZtZ+33vr3YOVhZxj4UZzWi3LCWRBY36ecs6YrvDxpEOZBGttDxqyPY02XajwSBdyj
fl48GU7g16WDwQFb1XTq6mc2uJs2o9W03daCHg5vzH/FDMisdwMgo/2vQDL1v1RftzHqa4+oN98y
wjgK8QzJ9AAV0X7QAwxXuIUaPxXB9tNddDY7u7KOBO/6sEuVLXw6cI1vVbxZLPqxc34fJ3v0e13w
n3eM6KvitsiFZ0tWZ8hV6K8FGrBWqZjbMRIKElkKEvbFGryw5ka4lDAL6OIG9Z+pGPZRQR1UdHdf
DoSzTBmbdgnWfeZ5+VYkKyIjyWgV5JQ+YHa7J2Af5lq5k/h5j6nCkCy2pTPib0gQMfp5prdEak0d
h3J9Fezks+mwcYVEzFo6hC59PH5pmNupbIRgmIDnIR4Fg0mnxzyzINzMkxb70tprdwvLCKhz65ie
zAh3nGZQ5wwInA+kNSlPglAKhS/L3x+q2c69JhAtPU7cNHbr75ABUmZu1amTbyZnbYqgTNFFWIQy
ZxZuL6GEjO1zbSa0Z/rVYLDGePsqnJ7oz8q0oIGdyRW2BYXXv52EDEIDGRNKxZ5Dp3dZZQQceqUo
6HCzWhlqQoi27y8JL587ABqcq+B8W/YZu9LnV1sqqrhTtbIu1Ju7cLy3LI+A9Yy+PrQPpK4V12W5
6gZqwHGXw8ZpzJ/vqo8/Jonlt3fZRsIhAOuE+2X4M9uQGhOX3cWxcHZZ0oiKA1b1EOSKcZm3mp1p
amoXx7qk9+2gbwxdgQzQJFsgZgnCRxp6xMHTmvVbJ4jRD/GjTIZC7uReIUZc8vr947utff+zYA/v
NEXJAj8Prk+E0R3tZvi95kuif6/3sKr7DvRUq/sjAyN4MYL8FfNrV/kY+6RXZqa+NFfRsip0qu52
j0Hw6HfOli3qfLBJVRuq/84f/K9B6nLS6mlQmbfSi4nHEE75LLuFj2Kfp6JVUXwSqO72Xf1b5RZi
YvrxZGy0pqnmeAy/TtrzbTywye8puHViHA04ofHrG9zuR59WTYZy4PjoKEOvX9OO1W7Tnyia2wYM
Fk2SdExU5fbbrmKePxSYyD6lQxPEMQ/t58QXEPjLxEfKv6jCHhkXUvsW4ZG50H5+ec2YOwPEQIBO
O1716xckfMT6bXE+EoxzDvC5lQ+tZjvV0+Kenv8yggcEuV0JMpiufvJdcXq5f1PdHi5qkjF9FVuu
nDWy9t/m6CZEDs2W1se621ETC1+xGoU//EOepn91xl4xg9OAKJFrk8On+Y9QWRu7NnWBZqQgaxXO
BfZ56T546AIAWLYLdrfKhmNSutphTn2RVTg/vNaIYjTfOEgNYkJb8hgvSttXmrJV3WlCil1kF/w4
IzsrB1NfIKEiF9LRohhulFdjGgdD9hWZR1eiFWwJ5xP2EEhuC8stPCCrWzv/XFOp5tlJvUeQl+rI
0iQUSwf3xZ5eVHsTXlrzQ/GyRaQzvPKZ6m9GNzurOMhRWUQrTJqi0O333GS43EtL78VRAz/wOUJ4
Ori5TyN3gBT/nqrIlcI4eOWolj10EJwZ+oAkK7yO07VCzq4hcLXGf4rG2P+MLXXO2EceY/kcKFOb
aQjhqd2M1+mPf9zvppftAjQknOCXEOLIcI8We8WGLHrgXBBlDTucLL4Dz1NmLgAc9UTi+AKQYAeF
uR1ZZfroRpkTVIXaz+ggOCqpSkk5E+ab4oms+NmPzHOXdFxOqSN2+pZXQWH9szEcQnto6MEicjOw
oml1DnSAJ5z2Jv6gJD6TsWTWnsKvBK98fr4HHxFe3GTXQPAA90BJSfCHjzvqXXLW+81MwWzbNjLq
QETFtOReC70jBPUcS7PNwc+1wCdXoU42bIYyx5qDCvgX7OlJn4f/m+R4JOl063Ide1HSh7I9Wzdv
kfPECYR38vITaTHypmFbpwDe8dPpAVjETjmhVkvSVHPyms1b1JTwFCTAP+d5znukGd7JJVbPCE1a
Xs5Pbl1xnJxQ8Oiwg3RQCznssEZ712xa0tcDOKn1gqK9GBLxhqd5iIR1wc6XuWtoEJahkUyJRm1j
H3AC3cusxWhImSQ+973dvxSOTN0tf8TjSzM2dQZNfLQviixjWap8OZ0fXVvrBHpXIoGjCnHrSO3w
heivZjWuyxCx2+7zdv5wgQfOQzpmUx8z4rrV+IZ/0jIR3dXx0CDEZt2PHw6yMJUC0tj632P6olfg
RbilBJhMAaaoCHgDr4obRoOwpoor9RWifGNjEqG1rs51fBGyBXtrAqKr9vy8ojY51Kmm8qFsQ2Vw
WCe2vASXgJGCQtKcxNKR+3Aoi8ylgCsX5KJM0d/4wALmzn9i5OTz2YBGa7RjNjMiFv8vE7QrLywX
9KnUD61vH41sZV8x73TNA07H44gW7WU3GGivrl+hNwCva5fWhP89sVn0Ji1X9ACV7muX8XXS6CD1
b90uRYReVqf1gm0CYMX8lT4EoZlOee3CAFm/GW1D/6ehBIdjWLE4BzJEkfc7wOuPI4xjc+4Q0Pfx
of/mMnMJWN93XZ6M/nQY4bjrZIsxGubte+gC2mx5vgwemZYeFvDhJjJHGzFX6qfkZsFvuII8z4Vs
uRDyJaF5Ad93UVB3K0TqpFEtuVUPVDc7thM82gTwRXsg3SiExPAvMLwIvwMvvjpwLu67OCDcQROY
nU5SGBehPUtBosoQVUfvp3iCByTUlMKYk0fC9FEUEY6uDN2g7aB/N0FJUiA0JHh97p+DkAoUAXjj
Ax9PCjZCkY5SJwfeO6FPq7d7tfmlXKTT+hQdFUzvF2uSIFJOK+SpBNIkctlWU5Ss4dPVLqs2zgNa
G3BlkBUsidsEXkvoNYhIp8fGFRd8PFE8B5q7ahRWyVOyin68c7ex17A9jhUkpQiV6Bz008D7kzPr
JKbEpslM6FgafGQ8uOjatAm4CamgdJM0EeuDh5OGEw8bqWj3abNFry9x/2o/SytKkFmWBC/ieT5R
9bTuvwqJ2S1+DUW2iRHBojTV26Ka/NYhVbxUKpBFw9HovzcClnSfbSTJsEezXo1tXvkdjU2dO+tu
cOck4BLDwDXcD5W3lRPAEifuTiPAGvENauijc59R05OTdqPlK98Qk3g9MngqytXmfPJgvmjtoPkQ
SnLfGXzfwQfY3ZPmoE5CN4y5J54HpDuNMyvs7ehjwKSRbL/eVCpeDtsiNMDZ2G9EUfW4M32ZU7Eo
3vtlYG9QMEbV9iOC+hYuWdG4sblPfhYwHSdoTolRpy4+wRX01Xddmmw1PZzADW6tBFr6GZf8hJ8V
o/CGDvmy2zc9UGbjb5SJ629nAU40n8GxUr2RCA3vyL1ZbQ+midpcsfcDo257m7PjPstb6FZnx2Sc
9QNrxIMjxgP09WiKd5dwh1avg0aUkbT9sI4gZjcQttJ5MM2zVslg8NMYHKs28/cxFrGppYrwk2i+
8VntO0zbgUxrVsXIS01U7eVbg2hd0TtwkwIWrDvlAEN++RVZ1gkyS3hkPwjjSk7PY70fEJ6puCTW
Ai4st3oPJuKccCV2cdIcelVB09ArdSOJLuCNEeJ/aJVJCePVXZohEU2zGDup7F4lOXN7Mr/lSof1
EiQHvefRPGXLrj6MG5g3KJ0FlqOIKMWYXKZ9LSZEhNaPI0CcDZ0rCMS2lGl0CptbbS581CvaTkwY
jDG+IH4brXvgOcqbNWV4aU+9DYlNh0f3SfSD/zb/SNyCy3oKDmwWG+SoJTxzdQqOtdZyTgnD462K
gJJ3KSIqO9uNvfvD/HGVLz/L27MtIUlhQ1+3KZ+Bqk4zGK5+D6fdW+o0MzfXWetZi1ary7v5h1SS
MLTwFTu1hbqprMXUMPagtyyXGyVm5g42bp1KKGcr1uXY+VaaMj1URfSuf5XpDKBVrrI5oU0hXf52
w1a4ss8wD4fgDPagQGxnOSrMobxx+PebAfryRPB1O5hPmOa4IfqMWea1+ecfShT2s3zxQD8zjOEp
712qduO+I49OVbEr6868qA33fFlJ3fJQctqko8oCyyIlCe9UOfvjoko4uUNBGLwAiyxwEfr3OY4t
b9h2kDGw2OWTJrlBzIl68ejGXN1w87ktaDDCAE/BJQAWHYHDwzOctJydRoeejbYJyaoyAswJvhU6
vqBMRUXEWmsa4uQ3tHMHtITkA+RT9UwKUyRyvOphu2gYa9JREc7jq84OmICOamvsQDtCuoDA70+a
l0hN3zsOOhvgFhwEciEhBpKczz6ZEt6aM4hfb/nL9sPpvGs8x0gOBXKdLy1+JVrVgqkyzpNSXMcS
cWoWT9ZYsISS+8eGRRpsJ5TaV/tx7io9EXSVZZ+9yhVxfW/Kv2ec4LsmjIgd7p/EowJQXR6ldKn9
cf+GkXHjveTEhqhZxJRzaxvBiUMh8g1lO9s+UQTAbYBM4onFT4BD1dUFTrzQAz/rPoBR9iFd/ati
l6P5I2rfzyKCz6hNWnskJPtp8IwBT2JPD3JK7ceGL38749NYfUZpxz3orUFCdT5rKIPjIUHil2Yi
W6LePH78ydP8Dl0t80K4Go+ukf9YuhlAN+CMU2HL9cLR+VvKgtVXMychEnTt5A3YqW1ym2mqneJc
JgWu4jPb0p2QhsSB9ZMYunaXwQOcEXBxlAgivRFGAOxp2QPD8LV/8sqKxTDKCCVZhw8DaYOLBDgU
YkeM8vHj7n+GeEGBpwqG/NJP8tdMTSj41xYy1lpCEk6QPAs9t74WaMUHU3WDx/K+1y/ujjQmaInm
75y9fnNv4/Eriwv8NckEM1/pl5XjWlJRWnb17BlaKx0tvkVWYknwgznTgfmeONwiNWx+2slkW9GJ
mD9GfGTunt73X3iOE7Ktnz7tzD0IOU7DNo/NtHq+kqFCni8D13dYGJlIQVmMgz2sxNkIxcovLsXw
4ZylpjxA2guDZcqEQ9S2wbdslxHoU8KGR8aOPT6XH2LFB/KtRY+jRQbZPJkAsjXhzIkeQdkaTY2n
RYXoOWzqlrp9oQENIF8yvjjDdpyVKp01/sMzJNRO2skCcMCDDj3LOZVwrpYe1ekRcCYW+TnCYDlK
1vkTHs1ohPm8AK4FlhCKODuJ1KOGB7ltcH3yU0h2Lkla6piOSGJCTMwEczzEHLB1Qt9n7Y8qtQub
qdvryzSbQi4EWZsbmwkXOUnSxYl2FMi3HojVaYqT1cNn4b+MamLhqgfSmmgbHcf5OJNQcOr5H45W
/cVVK/DW77cCI4hrkGWcOQ92iAzcC225jp2lk7Gz991KM7g6PKbX1gTDHvItILEoKsxfPoRH71Fo
aup49MnGcaRVooWuwY2yylNUaSsFPO9jUcv8NtfgCvO3iU9ai9y/yU/P8B4p7msEXCA5plc/nvZJ
HCBltLjqHy+7LR24BcatFGJS1MF580aVx+icpImVPBxdqav57GDIkhvBgGG2ng+pgwXtalx43uJl
57a/JnF8yFBCORF3ONhIPONgiJ4w5rgWMExMkVZRqOnQTKI2n6dDqa8+bSfAl+1vxlJRSCjJnj72
/S8T75wyMmpv4HVtKp5BwFMl3RThqnKb96rJjqaiSLVI1e/z1Dd5ByoSSTnFBR47xQ2yuiLnZuos
+HR/NJwqYfxkEbXyeriKY9/Q7e/gs+ilzSYA+AG0VsRHC+sbVoyCAsXrCeIsBNV9/ZAz/5gngxX6
p65RLcwkIwEzwzxxYILMPHCu1wtKCcg0TIJoYwrLfgKPJM3YL+gTQJxlud7wUfqdSL1qvmUDCHHm
nkQgp1jPUlymB5Gn5LkMLOZpG8Xf/UZ5aJ1HyRk8HfzK0oVU2Vkti5s8SVsk0DqhcGZMkiTY7yhL
GpzF2tikwapr6nEkGFPXqORI80srOEooBYq+5CPj6jLlMzQxlgRquSAuTFO6c8TmdZxsfEbx6TDO
a8ixWC/+lTf/oLl1E258Kp2ron5mTdnmq5xCLoIE7DfWRV/fzN/w6QGiip1xOqoztA9Vmbyj7wPx
Mg4X2T83OfLnRMJeQO5COaf9HJB182xunsj8cql8XYo5pGBs0AjUn4vvJDJYtxbdryKlu3RRU9TR
HEQ3ZMaRLAW9fgvCw0NlU8q/ps2bVkbK6FU4FBc8eh3j43T381+CJakrGzzfumuGUDX46J1kAo93
9lJYzkIiYf6MbkWSvI9kcSl6v1W9NVhEU6XxMQN0h2JNAqQcsisMcRw/HuqOqBkcd6mXkM0E1xuF
Q5ElB2/havrALU8tw2P2eZTz5VrjpJ1LVIIQOLaPlLcbbA9g2MFz8Iy0wY+Olc8hCBj7cGTyzT4l
8MrowFjlvI7JJGeJmKFbJ8FCFxCmH7hEF4k3UVmVO44pqdGlWSvdHP/lPfFu4eOwhSAQsjQI2UUu
QzRzgWtKSD/8frUJHPyiyZzx+g6gQUsGzjQo9reQZ3QzLpnugzN7uretYShu7F+nYSDC57lKR/Kd
Fibv6CXsk8ktEDHAxBqOWmTCpaa99LvV0898tIH0a20hb+6hN2wtN8bVXAzGlY2lBr5/X30BSe31
XxZU5WG73M5l70fxqTrJ1CLGzVOZ/y7zeYEn1HeVPM8xcySKN6bCSmj/edAgMgFsJv+Xm9LpMZgB
iEV1883JIo+Tx23M/xeYDokzEdULIXliiIDZ0iQ5vhxrU8i6bbju6O7RGj4Isro38qRvP/BRDibr
5iKhQ5I+mO8pXj5ta1ixQ+8WUNEfWqBwEDEcE7qyvvLNqCWwFH+M7GCvgLEkRMpInjTTi8rHSNPM
E7Px3NScB+UE3o2vH4ZVxwomzLYOprbId3nUBhelF5c0+WCPAqFWcC/m/Esx0c6RtcotNRxSqZv8
84IGlbfUnlN/VpBV1wQcwwzgNqTnkROsrRZn0Lf2UbrmltqTdM49Iq3Lr+8YSui9MbZN+HxEDXqN
fGeTB1grESl6gZZl2JZ4ve/Ahh7Z/+XLk4Pytl/ciFM6vK3uiULOzwJa5D34Np4H0wROWDmCcro7
gkA19Gl16ph15AQNU1IBV6eGFMxqD5VFHxmAsrkHbI/AM0s6p4KWAl1duk6bDrmjGbVuWg7gcVbY
pHvn3BwFCnoVTERF6/EpEwVora7XMj3Ro9S4h4uyZQkDbtgeAYm6lCx+EKkZRntFS0Q78LI2H7m4
OATcDBbczMNCuZc55P05C8WcndAxcJJXUkNqwOAVObRPERJx+m6QA13UedhNyN/sQCEDc6hlr9sp
GFrczGoL/7Af2INLcwKxxhO2CvZNwsy0gmDOr8eZvisd/HIhx2Z6VLPcvyEsxg9LRzsO6T2XyYdo
xOCgP7RfEDEpu4ZHzQmv4THbC/HyDNkLmNUChbeMx6L+MWBK6vpMos+uKDb26XQ+r1QGA+98R+i2
jekeSsWYBxMIHik7gC8gK80b3xi0nQ6XE38J5TwYc+FT3KPdDSYxYNewbYjNYIaVRfjXxFJRDjIi
atDYwQqPUpv+cJ67JTfHxBa/xC3QUpDL1Vh4G0N9/rWs3bDZ5uFjGd8JM6GtJGI7gPpgUGT1uXmX
hlxXmawWAVpI31fsPwqnAIOwFGo1JZrxNllPLWTXlYWURcIpHRIly3ZdL2ZTmVzHNHxUQoflwNnp
ukGQeCgDt56n1DunBu1gTLFbUnc08zKDDcRQ3bo3V1u/9DwKhgZMklGr8JghmFztxldTXLEZ/bFA
hJvtLZ6u9KfH5luv8h/kYxN5ePJk3QTTQ1Sdw+oMkMOnwyPor7vRGHPSDSJxc7nvk1ViVUEZJMuq
3zbUsFTLS9MKQcWNAVhlk6jGBj5eggr/pBm/VHBPF1ta1V7CV5MS0+ZzinENfyEqv5N6kv39wnlK
E+bQundjDITPmWTD2dDYWvsqAS8M1MAAqmjgmMbk2/QvzHMdUOqGG8MBOzYkVdevYMuYt1I3cQ2R
o3k3msTVmjitAztGwyinRb9CDHCXU/Nab5PMVtpJKanPFVo+fRc+gMlxLM93MRNrjbziPymBQkEa
g7OG3AWyUTH1an3YY1HgrjUnRoVH+1f06Y/l2ymcJQ56KLumbYjpNuvT1N99MxkKDbAO6jnIUrTj
e+jDCLnLUWFVfcjRAw7WqDY0Bo6kabDFMDVr9MIqGdNr1/3qJzaOuUhbD+kY2lC6b0v5wNIqcKA9
XL6Hn+/Qj1IRFFGHDDSca75wCSjBJ/aqnlYhx5NvSrC63ZvqVjOzdk4iP4zNK745uyvQWpSbP51o
SRLOFrGf34A62Bvd1FLnYov237RyvcAx0FjXGyTXJo/TSM3hRgPPVZK1Wsf2a08IhJR58DHFjFKl
qvyOdx4KIVROiZmWtvfe5ELlthNo7pXvB9+LNky1xytkFggpX8Y/o1iOg5nKXqlXJM1OKh7uUMZZ
JAsRTmcRg7Ui9nbnCgnu/Ex6LgnXRIx50v5zO6dVg6rIN7m9OAIG+u6EHrkd50o2+MYveCKWwfNQ
4G2MWpcQvOHPPtglMPPz5vGDvmBV08+PvHMB2V8a1NkZhVJwfv+S5soMHaqinwPtoOvW9BSfF2gP
yfJDnpNOFmajqmONlbpM3Z4IG0wr9rDUltQJcb1rBSI6sPRWp6qrp96rYnZdjeCjMcG8m+p38WBG
5mkV6XVMZkhjUhKYaD6pK/y2R/ovLy/B2H1mfgzDlBaiBvcrA+WRShq6/u/nCyd8icvYuKyPizpK
nmI3GtyOM6LG37VPc7hPBafrV0yfDbipIq9AAiginL+yEB7nnHhKHlboANL1wVwxrLORT4bafw4z
bPvRT39P0VU83N0Gxq384HY7rUA8tjqbg//K+Jb9Qhdo/aAbeLWNhqNaRo8UEwsq9lBG/dX/4/4y
jAocgEqMjiOkZw2hNCXjmYeVfTjsO6PtBrhdMouzfMjsHZUClKQw6/JXM3tgWrN49n6E1OMtilly
Jk38c889oCYMFdjVRl3g7sDdMpaSg7LNM19wQJ0eE8Zwbi4oCxyOKdrzfgKL/tqqtMZoJNtXG7Gz
8PrW0qqzZTtQS/oAWp58iaf4+VMbfVDbQcdxvTX683mghFhJaArhs0MpXp0NUQC/Vm2hfvN0/Wic
yiHyBhDb3mqn7sePvXqK4w5dwc9CrMElIV5Aspr9aa6E12EjINe+rSkjoe5mN+Q5UApaFLTYGCe8
6r2fzhcjva2loiarOPjNwQEbRnowBAh3+w2CpjAtqFEK/s9wY/VGS54IdSRddOqjFRxZm63jOzsN
2iPAw77KTnr4AyE2WI5NVZGOayFgt8Usss2pb3BW2SnC7WAs4T7s/rNTjBnBcRceVr5BdyNgPv9P
EphlYrXQmpLyL/vUAq8BmUq+b8eWdUCZkxHdNtUKSiAwEhgUwkWlEwcGfOOAZyG2kHyQU1CT7OPU
SGpdt7Ujov9WZ/C3nrCRAlur1sKVVBzbGLI2ua99U7LAO9flL13hfbzhD4JjiTU3XsiY9S3HJxhe
6+jBvv0EObixdvuFOGAmHGlHdUrYGHmiUk1HeIUjuNvLwt6Z8PUGfvxIFONvcikSp0cAz+4zlyrM
r67ySY66JchGgNW9g1dLKYnnhtm09siQf5N96KKNKQ4S3iXKmc68Vr3l4HBk6I/JaKnV58KTJm1X
k5J2uXmTswwCeDLm064vwUmL1U+aWGydHXM5GCnYJC9Pmo9Xg/EaH1nnR/ao/epgNvGTngL2vj2M
fv+7DqK3uTqhKw9boiQpU+6/0iHfAycK+8+U3ax5DjQqefX398RrXbgaNB9827BGmArhANR4ZifP
yCr5m47Yh7ecy3vsXdikTSnKwrF85YfYmycUJwMZyJFBUhQPHq8Io1I2fJYo2gNJ55Tv/MlLsf2A
3ODslg/QLgwbOjELByANUvTcm+Oy7E9stMLOvIMgfIAxp64OaJ586C6OLp+8eooeSd8762Ze8gvr
1rNP1ClB3IwVmAhokPXSvgRwAl5UNTKoXYO3XvWBRfjiwtc+Y1LGRA5z1K66uvO8up1OxNvo/Zy4
fWZnUatbQQ67iz2dsjfQcCvSfxq0LX/M7dkvZEWE/uUSjhpvJGqD/lX/+98YEs5ev/CS9ckloRc5
cU/ymd0cTdVn8jx7HKpDkJdhgaSuM4HdqAjddySwt1aSR1ghD5LJlIxh3cewUW4CW8vmjoSGIX6w
fTZIHSatXsIw9gkgUI353/2ShjSwrGSCNQAYU/oVr/7TUzP8BbtvS+XsASW59Eo+Px5zhT3dc5cs
QQnjDqs3bv45JTVU+LeC0yMGhEZpQhqpwvmOwAklDlbN4Jow7iMcj7xQqdSfBvBaX5nrlFUHCQS4
HLT6FBx9xMk91fpA1+09gMX+zw+E3BgbqHq4niaDzqqHxo0FwMj6VXN2MDOg7p4b9SUM+a6J/c4D
24W/YFcMYoj/OP5BcfKn4+kjiO8KzGuc2/Mzyr42TSgj3RvuUM3Oh2cd9p6OHFUbcTEb/PT3OxTe
HEky4G9fpWArzDVL75s2ZG73+Emt0gYEbWGU3hGxrHjwLV6HlJh2tbtZfQ0MtpcJPNFh7NhzA5YF
HE23+B6qGY8pFeUNCnQwe/+Azk2T7dZqCmAiVxYi1lVUcIe9CMst6yutswPVKkcYXux/uxskJFR5
A2h0co0BC9d0VHbRgYXOpzJ1+U5K2r36268Ezs0OID5MJCQzdh6SI3Aqcwc+xv5yxbuCQCqumgoO
uN0zxa5JOLs0+Q4VXFMHTw8bYC2+Q7qhiZxzU2R1l2NS7N0MJ8F7WarYoMKyBqVsXGDQD9uWpnfP
cbtcwehnCxh/PRcFtpLo4HiSigKqjb7LNkfOqZ4MrtB2bTTvQtBUo1N+kIjy1CgJtS0GAJh6Anqs
+zzB1bQ+Ba+9GJqR9y5De3pAgsv96Z4Wi0/s0oZv5zSvPu6Ceh6B8DTyV5eAGM6wcM3z7mEE8iy1
I/4+XF70NdHzqhtOrw3K/cgSocdkDS2d2YfXOrwHQEBVD/3VbqcAOwxWsOYEy4jK88CJ4+Lc17zi
glER7n4gRt9VRj0fUcqNvdBFnjJE6cN4zxB+lSHbydF7eMsVaEh7hV3mLyzbdQ/EbSv023O93YVx
nGDH48MjusF1CV1zHyeNetarbejwydUoocEs+6p65YPLk9YpQ2woyqDo3WOzsRTfEpfTMPEX0IeN
xk6leXF+bui7ElJYKOiUdgPabIzGXSER+ev4l91GELEcx58v0o//nVSR8d1Dm6qBlg0HCJZS7NYC
eqehSwA3SBpmIfr4nAL9MFjPKV7qLr61jzm4ClDFDQoagtWckIASsuYOp2dZ2Q3ypJOvNsROlhct
oLXDv2C5UWMhpdNceETlXPCKHr7r7GSG2znQZUoBGaH2rQ8gVIR9qqmM9qogWIZ2KzkeFZ7etSI5
I+8cOFYlVcQOrxGm5g5fhEHcE4rLR/twUdtFFWialuVafl5tGvC9UnyANkuSogr6VHY9X0XyX1bR
wVWIN+cr2sis58bhHBpF9sq+0eMj4pjBMaoAxrcDZIq2qnnSpNlMEQBFzxu7074hIWRGik/wxvKy
Lca1XzneKyfsh0ukxpMJC7dXOLTQyd6mNY6F4erY1Eo1hHS39ZDvqq4CdvBY/1GQKCmaAVkTMMN2
P3+uG10x43oWsMpA+wBRHWHf56lTaCpGoeJYr/anuHSqQcMPbrVFcNFiIFi9htyO9XBWiRuT4ok9
6rTKyCaxZeeghxkGYjlAewPFFk11a9vAxxMGFJUDS/YG/6nzq7I3Y6zSipmJ0Rxrzf9f9e/HzS8T
0HAVxAr2uq1KMW1tQR/Z13fZEf6e8K4V2D3cYxqa/5DgbksS2Z/kKYzxQ0PSP7/dmvM6P86lgV/j
07XLKkXcwBj+Q1iTYIqjZpExXPWlcfvkCd735sMfEWViCT2WHma1wrU7DMnzfiPbSey6mlvUYRgg
TFDmXNi6dNjoOHFWJL3eWGFy3wZZpflOGA6APPnrLQAsuoVxbyMBxhM7OU/Xbw7SpbUhDGU0v/83
pEKT6p/qkBdbrQ0YTPeheSsjg0/2TW6HgYauri0IA0xaFikid26Od76La7nlkcf2nnQsRBnMbFP2
ZdSu8V9yYrEIZ165Pnqb49H9sUpdisvKZwQDqqrgKYi392ygUYf64df0SteyvC6AFkBtj03xypRx
o7OtjYoYNnb3/CPL0L0NnrTyAoAUXL0aoF6mqayfyJluFdE4k+ZGM9txM9v+stDuDeT5K+TQGvex
Gw4S04M7nGjPLMZBei3CjYPss4aZIpo5ZdNnXQKrVjPNFqbbqcEY2mYTXPFXi6eI5M6DDAr3tPmK
itnAh64aulDnT3LVPf2bu5Ci8Aq3/1lQG8GEFMSHTfZdiT9vrjPlcB887oTTTYO5dUtxeI55yOTY
0RAw74UzTvp3DCv3TSX9Y0t8nclx8f320QR4Em2DynTq7pIpasTSyKN/QkoSe42t4vO/GkzKArTA
jtp9hXTardMxG7yfHiaCZFRsfjvCqj9H+rWQ9XstYWqWIGx2WpeS2DfwN0uMAK2N+83ceJKCCkXh
H2XPfKVrpd9NvKN+ov6zmbvOi0ZHGRYP59RBCIQ1hQEFiu72D0+w/62BRVHo89PsqDCgHsyZX/FL
R2kfDd8z24SDw9VVREKoolJnJ8/I7wxmxNH0P6gbhqKhO22/bwqimyhka88TshwXBlXDUjyjdT9J
T8Q8zkodw1FSQOgdZM/HAWcxQcUZdIf3rXVNfykBkFriRKGxfVN+N/deC0HQkXxov5urTgPbgl9I
nHKl2kXTnQ1bZveWKFlbi8+oAhueVAuW3+Q2KJvqzciW5DnlVQl4rH/n+dsoTwR6KaC2JGCnIQtf
aCnDZmiGZ6gq6M4QQ9NrOxMkz2Y39AHppbvPtsWwFUiTeaSe9q1E5SXLc3rTLqyBt6kk8CXJe/lx
1Us1FuLnAxC9e69it/L9m9IoHQniZap10VH+yY6+A1kCLtD0NdxQHRHS3Rdd+iysGNAfor6aqHsu
K0y2tjkpNsCh3Ju26Yto0m/1bB/nNsm18yEWL8MQo/+7GbxWD4dsOMRRDDAdGTmq/UUqBB5VgRco
qGV4xNHgkkBbDgHh99BfgLe/Vn84b9PrK8zjgoyOmHpl1emgqvAEkNY1fpFuBvyK4TzJ9SebC+/V
dFDZTDvqGklAQkFRKnm5gOVvmTGtnaYGGdJD+MwKQaKIxbaF2CPCWTsc0WeBTVfASTd/eYiGA2Yz
sQDS5WclByNYgflx8yUXLnwkUfS9adERQgY3hYlLknYe8tmADMOnf6BST8POb1iN6v3q3UVXNo9Y
8YU7nxyyvk1bjyIhXKTQ35lVT5e9YowSxuAKS9lHcqJBMp5cyB7aNsuWxpSpDW90vMBVbWb1QAWp
CalQcMi51bU315Nb4Hex7O6AdcJxbMGmHTgxpNLTYSobeRKhBNinpVAvgkL4bRQBbQIjHoLL4zvI
MUi4Y3ppdXNGIWQFLTwyRKp4B1e8gz+ifySrge6AxCnLGSQQ9FTwkeRM1JMx/+eDG1Y2oHE3jHP6
szoBH12Ykiml6Y2NQ9mNkGeTuAspYZ/9PiLFLxLYK5I1Xmt71cUNqNZ0XtWN+w9y7VwmoAiBN69Q
KGi8J+IecyhS4FrdS98LG6MLJain2i1gH4LSnuYd0Q7fcAmgLXne5QmNuFogEu1mgc/iyFeQ2aHu
C0sgfP4WYaeq3AO5ha2dni9yvnJBteBITnVPUHex5Gq1Rxk1IsZ+Fv+UV6Pmxqt3uU7GkgGX60mi
zhLs0QbbT3LmpB11lfUPIN5oCJiCA4MwtTUsFrShY2JqoOL1nMmiOTWDljkckg3khLZiaAeMkLuX
DzW/73kFCxP4EhaAqYXAcC6aYY+TCHh01Va2dbtuP6bqRNMx2DxR3aI0Y9A/uwFjPLUiyOIaGkVx
UChDkpyTwH9Kh2UlISkWbd2O3IxQECSJNtc8naYocLGx7BF12201TcyGqjimB5xBTEKoMifNnDZv
Ruj/Z8UIsLg7TUKpk/7dGHz3nASdplIawvHBnr1aZHDxsnWWmj1tC245eJ6vUifuOoCT8SoiCYrx
+fVdpRlY1M0D4zTyXvxfsKHJO2RNB1rlJRAIDSMPCD8/v5CqZRNRQplixYfzI0CdgY2yr1h/D3YA
nmMsWz3IJLk4OZSqVPTSumPN5SLaXLWJyYnVo3MysJajz5KWMfVRRuczmCuw0l3VazJbPmISy65q
E/MaiofS0Y4JkIfsUM/gQL+Le0Pa1n21hxn2P0Ff6c5h+LyiiYkjiaQ7YY7EqDh6IKS11bv+7C5+
U3CGzRTp1MNo411Wpl72nQeQyLqxt+0UyAFJlQf3BAw/xgJX24QoeWrJirda0DF2zngq5r7KKzlU
CTDn2rDq4OBcPmgzOOBlVr7m4LQPiENaSZTldqgN62zhX+hnkF/Bd7IEY3MnRwbcd/qBL6EcduXi
asXeH+6b1Pyt06QbHbDQvrljTo2cvBotkFPdltLGhlHvo6zF9HPUGTaV61b0sxgWXiD7Kw5Ms9f9
12MEF2cNZOyyhPxsz/f415rb+/1JymyriGMMzdGE8CbjxDXFAs7PRs9tRV/jC6Mlt2sJiKN0FH/C
a51qUx7dOAObn2QoriTv2mEqPT3+CS51GiAzP7sJwApJOqY27UbgJHlkc+Irh/kTqnB/um3Z1CYB
Wn5EVfKdW0jqGb3Y4j6pEf9+pEL2Am80f/0ZywFwtoP63XWx9YEq91GqdEnogfySfi6k3yi5E/xI
c2T4qqVnwa56+McwHqt6w5S6/BkxUtu7eU7cWfdmRZjXjeVGiBPEALMzXfd3oKs4AlGPdG8uic6J
AmKmhFxRvdzoFGP9C8IedjME/uBWsxEcJiMS4ccVsDhrS+4TLa4iBwN1eQttDvpOilBp4WHUNDk6
5AdgzOps8iIIEOUTMqRfnx1MHKia0ITstgtz32zDzP8YGpxGyLvlqChpqx9PM3XpzuV0fOsrsvaO
jwmlrTBscg41Z3r+Ez7nWZ12VvIFDUHYgNrkA7xZd3/bKW0S4XpIiEEoNEEZdPC8gIbkHOsMUUyD
AUJ8yoQ5+9a8pNlFhciftr8V2d48enZZHVDsm+cj0YBTnF4sbFm7ISMic60JJ5sSNVB6+3XmctTF
LPocAzxfHNMrEuoOJhF/i3Am8nX4PYbNn9BkE8l11UsDFjm9Mp9R8qmbIlsGmj1EvcmlzMzGiU0/
rMT8Ozq2N9kLQ4DxLPjZnnPV9WieRIZZ3e5iPZLBz7iUtLGYE0w1sUruvXUAS/jHTHCTvupld9fd
iJovmDX0gNciZ1wuyJ72QGSl0IRT03yJAlZaz4drT7TL/KWwgrEwV/8vnbY/cGZCJluH0n/L98AH
TgJGGDc9GpEQOL/yWW3aKOVYmxPLrQLPOkzVuCfz/xPs3hBlp5EijH8TAXCQGbSfAMtEhVnvZDfC
iVjEvxaLNR6aiEPRQCswc1k0YOqt6/0RzyPpRaRt5xndooksrTxDynMWvk+6AdEY7zO67Yo9sHCE
qSd/YnF2yQFnpO2iplnSilcd7OqsJQDqA8gcaiRskW9QK+7w0T4NCO7vNp+NiCdZJi/284jHzzWc
Lq1nFiGiuWi24xt2R56AHZpjGvqc2lumuwDv0CD+m46vumPwXJmzzpqATQ/lkffE2asMXW2b/j1k
Mse4aaFbFcXMOj3Yd2FUkb0CZAyXXw/0GAVK7DQKhEd0j56i15fVACDh1cLIuY7GwIXrD/rsMnTb
4zMZfHbDo+17kagrCEdzzR7zwEDO7W6m7YvUpZh75Ut8cBSlq93FKOoxg8j7Az/uKLtHJEE8qDFh
RyyZrPdZ0nUfGLNnd8t6auAmaIC51v5dFyitMwwHecJ/cKWBNSjv8cO20BJlzipv35k8EdG2H2SK
wvES8Wi/TsDgRcsbqbRFUxnJTVOMQSI9dsn+ARthDX64HENfmNVn7T1cjOZ6/N2/RZCvyxPE0GcP
8dbVM127S7c9r4PxzQbWyCuiVSW6oq/nRmSBINSq5HOmX0YhqMF7nM/mNOoxS4Yl/0+JFhxGZrMI
ZwkYz6oKtEBm2CvC8Okd32XLIwkkO+u+G3qhl9VhSu2vYvf7Dd0p3zy6y+kc9toSslHvwcwoDjf8
E5XFYPiIzIYXk0LowuMx6C5ojwH6ldCfQpsXoqA9+PkSWKdmrqp8g46aUPxhtS+pwXrGAx5aVHJ5
IgBH8Sm5BXkwarstiHZU6RkE4yXDNlZQdbDqadychEQWH+6PN7kyT3+iGAh53AqdfgPSXnnUEtoD
pRSdxiUD7xYuMI5fgPRMnAkrWLMgyBG2xFNJeaZJ9t5lClnaNHcO5PesD7+a3UcrFY3OgyxeFeOY
piVrNaTAN3L+x5KeokV1QzxPXHQBOGdkD6FVTiNrYyNu6b4CG6fGk2qDpASymM7xV19/KncCWZSf
W2czr1xI/Ulym+BCZSFXFXQT1Jfiz3Pkrw3AbN4YgiR/WIuQrJ9BcuMdv06wG+JxE/Co0t0fjLXm
Li8LoOLfIRFQ+mxvDkkJemXFJRBVNMLZBY5C7Xlhht+qks5Cj3KWOJSo8Y50KH7cxf1vAd+Lkg6d
oF4tGtUV30tW2PIimtJN/dV0/qukZvdBQXRujR65MtQZqXcGgo1s9wifUfI1R9K+RlpQa5P/0mPt
Fsz6biEVp0j2tNMf6MpouDYgvojGLXxEgK7agWji8Ev9nM2IgJZheSSD3ty/x/H6oVJUmO80zvbW
jekNPQmNzBZUtQ8A6LTT11F0RU/ldJZOFf6pF5/TYSXj67X3umvriyKtas0dj80GwvCEpLcL0mFE
ER7l4CiS9sooVG0CnEJhI6ceWsuSciPltOJ7g3V+mje/oIw0BAjCXzI6zuAz9I1w6llV7vtlRRkz
lUTrClvnzTottKMjXEXst9ENlQlnkbPeZu4dJ6mg9xCwvc8/kX8hUZd7ggsjA02c37dpoi7O/Yw6
nObbiK1FXcPS55VYQBf9FPL1IjSG9fg9OHMhgnkYFg3tJ3b4dK+sEnkDpCJEQaNQwDE+OEXGaSnW
38bANeC+e68rtxOYyiHZp3JZ9vUwLpMBMQ8S2fL1qPq7E2o5NbstRASThNkdykSFFW7GK1caVmTn
sJbEzSzPSzktcJZCLV/rxR1cW4yFDl0LKAnEE/eBddQXpIZYBH+0f8GSF0p2tO8ue7ST1RfhJrfI
YHTZzyeBav/4yXbjK9X69o2JDq2SjA/NZeDYfNCNmRG6cwwOAHgMsOEFZM0+7Hhy2pAnubTt04XH
0+N4K14lHFN1d9jWa+UGmn7Pe+GbgcDxgLAbMZfYPdYbwdYAyhciVfLF0iROA3FNNQXPl4FIqDt4
6VeUK2ejT7+HhAJ5yqTB1UXB5QQk3lZ0AibfhJFupznCBJAYOrR/HkLthpuqSfI7imn6aSTkn87h
ZckIqvlHEvnXe7PQLAUcY+TqZJKy9i+0430lPsOqGMWFtox7PpjHdXrGgvzMVqYrFny3Aku83ZNE
o374yeGejlGRswoIwHaO2/h4hJkoot9GQsqxpe3HqOAQEhRzlAaWKEo3WQwcCWprBTbz02MjLO4W
dTHz+Y5GrofI9t91Nh2u+ELF3VkoFX4CmqhLXKEXrLRcmq9r6OnAktSya5mB+f75xA2wOqRtsP3u
+CP1Kki6exnYrDr09MOhyfA11YeBzgj2v7M001DZPFACOeRwc38rjJCuyBiw11Q7N32yb1CxMVKj
Hwu3pvd3tweIWaw2cP2zhE17mv7Tm9Jec8PS3HKW39Kj5jXoJFA1Mu7fxQmlJu5LsJ17d6IRC33R
dcrj+2Qyij1CGBU8qLFSDiySREqA2hftqqklcvR/ZyBaTBw4yzYtiRLcOKSh9RU8syzXcrgziAGJ
bFmpPPkR+SozkPJiNljZ5mZOj6EnnT74tdNXljatKSs4yrIeyYxCax0oKGCNm0MuY4U53gn0mxQj
XeqYaYnPYYJCVczgcO29z9gS9hMhxV5TU9Oi53eqn6lIL0IZpQpVEuLsuwK/DXT0ZB4suWpKgyO3
FACB6IDeadghgcJFRoZgxU/Fix50si1a9H99wRq8Bd/XjnU/s4ZM/jFNVUFPc/KAi+TpHJCE/lu2
hYcXqAtIbyKHSuHg88cB7EkSBpSwwWUeTtNrTWBXjIRBIe9ew+4N+Fk2dUcppSAYl3h+6/W3JOKh
x3iLccsFzHWPgmW0anbYDVhecZ8NM3OmNygXkSmqORsDdSQ/VUD120vdirPwRSKpxkyEHAlAoRuh
2gPOKnqJFRi7cFs4ORWCNpTVVebUWiKHBBu5wULS/74STxBRavRCNW+lc3YPTBwY2jauDB9KwUsl
1t1b+IlCTf91Ej6RghwbSKGAcOsq9hD2Tr354A5vdtLl8g8PjG1oWp16l8SNbV2+fWcC1M6B5LAv
sIB6C+2uSnuIHQ4F3mjxwh1qFt9B3Vs4VP7FsaF8Xc9V0CdbaztedQQizAMctXnXBHVUCO7jJJwQ
POruKXAMBuG0pOjFLZv3EnoM4q6ErkymhTt8kEimA5RAZchGzXTeQn6IZLbkMc57KA9npqTU8qC7
hjPmIG9PiCQQjTAUIALLy7BBajulHZntB3NXKy2m0YDAYTiOU2RpWmQqVM2wMdmG6ncq6roOW+fM
a28mpq33hcTgEgAlLh4bP1uwo0FuhZVC28PZupkYiMtqxDNEyyg8OqjcuP1POPKnx3MKeA9goWkG
YVJMw6VHClOHKSHxtaaZG+q2YoeGJVB+9T6NBMWtwhXiEcOls2774bd3/EHDzfzNinz+pvvAlVl7
aztok01ktKlpbre4HLC37Sh2SyeGvijAdXdWhKs2Xsy2dWIFT2S5o4OsrWYthh/TmBNWEARpDLuT
YvUft4gWiirpgzuf+hJbG5LEyKcBAxeda1fnRzUdxC1YnTA86kfm7KYcC9tdJ3Tr7VZNyOUaFdci
bN6+wW3OgnwWY9v6M2FTAKAyNdHNHyAGt2I+jq6mCp8T3DJ8biPqRnjhskv6MuVQSqATA5WyMQEu
i62g382em1upQ3SzbxrPKtv21LdNjIKQ4OxCGUvNgEYDLADuyVKusUn+WTlAEVO9dT7biHfgB9th
D1hJQYJb/Z1Y4NjOzgSkVhN1Kx8Xm0LWYLrzCEVPlG4MC34BqAul/PC4rl+NvjgBDMGynid3RSzH
We9RDvMIy+4Xl4jRV4WDLGL1qJpEJbB7MP3dQ7T/Xl6UsYvD2bPqikeFbT2hdtCnErDoVBuRU4Xm
JHMhiv9hiuucIcIVs09qgWDfN6RgqjaVotZHfzTTcdHe/6in+BplAzrH7tD2JpAH3EtqoxJXElJO
GhyAWdUgf6Ixpyo1d+wz3xBvdPogBuwA/vlMrYUGaxu//5ipdppSO38N36LinhD9DqGwdt70mjO7
Bp2XOFJzTqdRic9uLhpXlGvpy8vOhyqAqyFPt3yzC8QO47ls/krKDNj/dgtxU4eQe/oQ+qvn9qOv
i5I4F8DcCb93gU5ddUFJ5e+K07PvDDKJh6xpPo5g1LgAlf68MdzLTxFG0cygNDSNxdj9VAxfbYkI
/HVV7sucirbeFxdcmfjh9mtoKHbnHN/G8DB+yvuOURVeoDa0yw98k+gXG4qDQ+r4e02tyMixZqFi
lGmFtVG9h/vl0H7sUvymppf8ldnTleL8xFe5M1CBdeHnZTP+X39hPZYrxrqyW7NV1Ms5aweZ/sK0
Yhwk+7UocA55XMbMWJfI5HFAIrJkk9OfHmh7qA8ygeCB73yE/7Zi9w4RJuPNrOPfeSFbmY5+bqYe
ebqWh8vxQ9byyuzfsvIFfDfm3bzWfYRyOTplwJ1mK4EF3J7HspXaVkH9Z+Ec8cNDmpk0i6B+cON0
W30ffdQeXEE0wi9ULnYPMJ080F/3XFgnBzQmkY3IM0VvpGzJ1W8+VJ4AVzvhCxUxzY0u9qEM9xUf
smE6zYt65ESMpFSwljfEG+KxZ4V/+jCxSV++dLxkclhZAvY023h5vcXmKkPcezohpxBUVaMksteU
qrMzC2DdPjinx6Y7PVWts74R4frOXY9IgkjjlwDjE+Oi91+vYuEqCZ6VDIncLOzXixw07qr+zxHk
ycoWMIugVxrtBsWa4naOuNqle25CgtuhsN5VqRkii1XBSgSXwyhRJCLfDEx7QOmHHI4A/herSWD0
L6fcPy5hV66ge+w7kmjd86NUZ1gbfITRJD7k7SyK+0Txc7iJ0CzoQIUtbqnJPLWzIz6d44lx9F4a
Z5x26enGSprGyNAuZDCRUr/fISn2uHI6k7U1R/EcjhYlVE94u9gdS8Ncg/jJ88gz3Hg8TnZGCRPj
tatc1xu2yAK3bKVXXhzSUMct1WrcBEOvH+8GZBBWB4tNKuOGTQa0JdbXBFt80aO/2FHzZROLA9As
s73KfSTlhKyB+1kbMftUT2Pkj8GrOYtd1mP9BncH/KSpqno7Kmz3L20tduyrXxIvSdhlMK6lMokF
jqK0z/apL99Q0kUtp8EQGPAseJgaIM9U+Y/rF6s6JRmIh4PnuvguHfoVKByKmnwYPf2zehH6+7H5
wjBc+B/7BVSuoZQbJFCCW+jXEvcgCZoDm8LyUIljv2XdlL7LXPLTeg8Q3T+IXGnyC0D7LtBw22HO
s6rcufTLW95BFdJgioY4XGtt7s/jvs76qqoOSM3ohDSXyJf2LiOQqH3sG/gJJM1UwJzgncOcuvX5
hcYWUdUeyAg5ZsPG/OPS9HhL08hvzR1bb7dwWyNIL51Y+fzTXWUaWEdgMNP+O0uZiG0QtC8pxUmL
jtzXg4yRoMyNhsjPwOrD+OmuufVriI7SdEMzHdtpenP2Ngni1Jf+dRDkcCTgPguDiqqsaZ3+if4a
4Km/PdZRis2FpjfJ8zzrg6cbdzV9g5sSofaS9hvr5dciRGQx83TZwVt/hpLUBueNFCHd/UmURNEp
vgQO+Ab3MzUUNlU+EKmYRrqvH/AA7yGc8TXKRb3BtMykwKsLXc/g2kae/IlZXkf8lrL7SNAx0k+M
C3z1TDd+tWc0zpilpu9UuhU+mFal7XwnqTBgRh3mIzVQwxA1K8UcpDZ1InotlmOMZPYVPrMxYgBg
v4/TWEpBvY3d4WJLdGnAJQG6iKByAUIo73QM6hzKM2j5Bko5G4yxvHCkiyh7DSQPzGvyOaQ3WgXJ
66tws5G7pdRqxD/8XkjK9cIns4dxj5JYfTS28Fzw8h+eDfCmK6FlpiHm6O2jLpWq/cJu7u1u0o4n
E2t/whk7vnvW/oXM4wngXsuZglGLs3vZ25issidsBZ7w1B/BnccjQh4rl6ldw4c2WKhjFaZnv+dY
6iEgcDrW8q2mdXyH76TruEHGA+wy5A9LNAuRiq/dHjeCiryb13dhyUToTvUj644SkSfNw3GDPy6P
TotctXhblpLl5s2AOHFJPH3yjuqatuE6pNYmbF6kGvzzru0DAow4+Dl92RLUQmpcZDY6+ZhUUMSI
8b+Kelo6LBOePuCtkMWwCifAba8VmLwy5P8W+I9L33Zb9hPJ1B0e89v72oenmHagmpSSPhFG+pZF
i9feSeci05zW0EalmeB5SVFdwTRrv5O4S5GC+Zdu7Sb6WNKxEi5z11zfetFOhXQ0mqpVhtJiRQ9v
Xgu+AsvFkoA7qMmr3Yn2Iim08CL6CKt1IuCqW4DSTa9vwBierFW0sCgcRE0rlJHzrVjlROftyd01
vck5mSCmdfpOZcBAQPRgVZF3DhRjfeWTzwddH3gW7se6udr7To2e4kvD9Wci9EvN0efq2Kuu5DS/
OJGLK2vgrsgOIOMgkuzHB+Da75Tj47vit6el6WfJVwtlx6CH582lGcC0lXdxh+trlEs57GKBTydC
5Pxy1gaTOAYqEOyfq3nR4fJrpjOHKc9e68XxdqXpFwgHdkiOZQPdJDAWzWuUbt7vSVeS05PlBv+7
N3thayswNL95XeUPc8HWHTm3uiHkTb1h3n6RmuN2nqKY20kZPoLV+GHDi3SUVT02v5v3i5IfYiPL
hZs0Nzaxr+8hRwKaWGyrjppJtkdWoOktkhUWoI/tZ2As+eJcHWl3O2Z59vNDuqPUC2nf5eqenHH1
B0Ifcx6tWzZgeCsXxDIwDwWAA+VTO15f/Wog8CypKfHF9o3WmKAcwmFQRgIwPe41zt/uta4eKH9K
tRepWJ8MCYbLsr/Z0duTOvKJCAdODzBmJkcvcJrdEDU2vCYPMo/lCCGxJCkXTEuhGCl6VZqQ1Uyx
75MhyT8IltoUOBRhBQPPZ7bgGwgQfi9/wPzJ9zWzDB6cBXOU/3vsWxwgfmpW2M6HrxsOiRkZ82vv
ED+Qj5Slt6SUSeSLmDk9Hay1vSHvLIty1Be5qP4VUYY6YizLghab1BXPck2H9IAKEdqyGMeuCdBj
19JZDbM2dJXM6Teib5tcUAGoPH9Y7mcybE7X0hN+KCdh7JSFFK7hDRU9Ju8t1T5EpNoKKH7lra54
TctFZUgFjCpzFQLQ3cwzn7C+Ic45vd1BjSsEiWO2vLmF4TfM/qx+6hUD016izRu8G21r1RTapKZY
yKTEyxC53BPEyEh+BvLawbTBeSooFOpYQpBqWUQG7bGCcAfUdLXggs1AJPt5Dr39PxrVeNarrA8h
vLh27dwU00g06MMCnxzshxXCYI9SxdvLDFRFYokcSr5o5d3U1H6ujWG7tVBWqtLNmkrH6AwaN5ON
AQ6vGlZYkIGmjkiZ9hw7fHGN/oLwZZMR09Md0BrlZfbX+eQApHCXk77hLy4SRnPLXTbeFkMxe0cK
rspZHHdUs/RILF5vHRhTHD8tCX3CnzSiXoxfkT/6KQCiiqIJoxYn5BLEBojYXqBd7QZ3r3IAgBtS
elG1Eb3JDXBRa0UC/6OG0p8h+2hBKShFVmzoLUs6mOTNwB0hdeZZFSGN6XXlF1SSFUmMZcMIdufq
WMZyd9NqzWRipMzBuDfE5agw7k+z+D0c5IjoyBhcpUMQNYJ+017OZHS00yjLT/RoiNxPg5H0FGGa
0O16fQMN7D7Rpbs1nD5HqY3Rn8ILSi1MyiXO9GPYCHBe2JA2XR9m6XCNKwVtmvdd0LJJ03LuhY+r
+0tkAYSp2+Y8r+jQntBgHISnzO7ZqP4VJaHw3OMsoFF/v27EVzUVaI5rVo4nsC4de1Px7BZ7m1/r
/Ed/QaVskopIzvo0GWRTffy+/G1vhUzcF1IuEHyKzmnfpuNSyaz7usGWKXheT1vMzSDMwXzh4GfN
UB87izXHFICKrYbpfPqnFutJEekL+hg/kSQZW5utKRIXbRDz9QLaYeruCDPCtJA56wyJ1DVBxFlb
N5h1oXdGir6S0uMybu+fKm+ViOED4UHZ7XJo14f9/a0k+tyC3inAsgkte55ZFh3wReLQr30fqUCj
0PrFbOUxIWPr9GIpAZL6Y1i+PKWqJUVdjg0BSeYNQr2jn+L95wknBB29J3A6O/uoaAfpXuPdxg/3
RMTMeFw1Hia5BBjEskphYR24FGTAT3fPFyQ031XGCkLQ6eWUZg8omXDhGoXnnC1/npZX0L+yPZP6
Ogj5EFrh5HuBS4gwrdBEu37QhRzrEykn4OAh8dBVmIo5H0m46S1E58vWNKhrM9OC6x6dHkmuU+CP
DeNl0hYRGcSl0vpiB47JgSz0jscyeZZun2GTooYdTKtlyMonNFIdP0mmjCh0DDRhLqjGfphjBCaH
jdMf4aDooxhAG83m2CGC0ihb0wmRVuylvF14C6JDDdhfW9p0aK/lhPP8KzsydPO5qk1bszjEezDt
E3fAu84i7fsvKu1OVUApxVFu7B4xMqU5f0hrVs6dbeIWBSi76lfLuySrK2yEiw8q7a1SfRLkPDzn
KuZ/XaG8/ou0otCQgQvHQ/gCyWcCgjEMqvc4ApMf3bf4E2tQgzAAxvSmDKAowE0Y99gpPkYyd6Ga
KA2DAqu0FoU/pacNL/gLookCgwQgkM3e5F+9i4uP0OQ/yC1Xvpqt+L6Tk5YfW7ZdIzkwAdVAj3Lw
MKPf5SJB2ZX06y7MMgJz8p+8wwMxWQ2rfksTO/yVkJT/yAGhJ/mg9EujqsOKxGszLVRVXzZEUoPT
kkdWr7fe/iA/1Fn+qCOf9Qgc1mq9UTH/67VG2BxmjtCQQXdQTH9lF19swrjxc8VozQ13DZ2u+DoV
+02uSdyCJXARk5foc9xvshrclwY9iKY/XqeUIONmXST0NYLIlJfcBhMd0+uKYhlR+WASdh2WPM7k
EtaH+N7I31jCFeXypWn61OC2iqn063SYZDKZzJdheDm0VW+7tUWkQAVGjpxjNSfIQBXmEQ8MCQ8m
ZZzkxp68PNGZ7rNdTsQpWI0oJ1YAAJRfw2tLTh+dG2gex8YCfxcbxODlQnQBeIbZ4CmYvd4YapXq
EWNR0i5O0VrVOVj3AnMBS92af3pOeSkMTWnbjFEoLeFMK7Con6jy2p9KrSIeCzTXT2UfkJdenEta
ZYsrKWjF+sjd6xnw4XTy/0v2cuhRRGhvxkvv4xe156hNXP6Z1IshZ9iTNtgleoO55QfqpbEorDD9
bs+3BwMu5S6cBfBLHsRu30/zP5MgSXe0BVD0raqYHJjUMQcZNr+hj1FrKC9Fat+HNEdoJZEgY24v
Yz8rIWf0b+0EFfojZXh8O9S9D7qVLitbPxN9WAQ3J3UJoXP12Fh/v11wBvImEw+lZnFQ6MH3aubQ
/JbZVn5AAHDWPGpPryZS99B5kzYAJS7GvjhltPTCpokwYGKRL0Nvl2JddcQgud8/HVWp6wSkBDaY
c6TtRt9ZWE/IjV0KGyDdXNGS+GM8E5DbwC2d7Lg2xLoBGaWM4T2iPZ6U21+m3El7DVFZiDNUpw+i
4vG/CrFmqntcws1RgVOCEonzlsTRmO+nXj3RJKMQIDyh+zhqH8cP4Y+9xzoZQUpa/J3HCh8BJuRC
ZfsHHySsP/2tc9dM4XYQOgIZcpCais5vQ8474/0bnwTrUS1xjXouCmmE+C9QsukiFpxHvOVu5Ss2
I0c2vy4nxuupyuZn6+sCxN1jjCKFX160aCzrNeSP5y4jz+izmSONugyAWgvyvo1h2kSZEWbzs3zn
f5gur5FoT05ZJnWSaCy/CJMK2hLZ1RJo7TWqDKiqB5zFunL+OHyTO5BeRGFOKaTW5X86Y1myPkFn
bMZm6I87RLS7xPoFwbrfMdES1Hn4h37C0pyqgGifr3hV/UWm+I9yNCZYfNhkRCZr3n6bbT0Gt7E6
PupLqI/Tkl1ZKJcFRZFW6e6zD/lkYGebHSNrgmCf7HJOyY8VRVzN8LOIwrf42IB+HU2vc121BTDh
ZfkiAwmbBdgDlV4cUG53BOEiR4qszuLzD4PtGPTNeKluFjUndL5wyNJ8BNBmZ/3akp3sqLAIQLz9
UBuh/uKZS5UBrpnA9ic8AtNo0GCyxkDOLwjlpz+ZEar6UxyDppzC0KBRJH9FZSwCTVgQjf55T8UP
00sdg57qOm6epM2NaOCmEWZudIZsN52sr0QLF/DOrFGwVkiKA9jaUskv3Z8faKpS0lpyThXJT7ke
3MT6P6W51duTizyqQHAuwt86rw0YNoyH6N0lPdRPDKUlZByeGEZpkndwV3tIOTQuGZRWTS17vOpx
yCuzVGu/2BcwP6KH7Gzz3euZdE44cRu7T2CcK/IgsIfCIcVrYEnEnYhBQWN3xHC6HiyOk3FRP1bb
D+mL1vqa/iG3eMjs+oHDEszbV3xVH/eZOfvyETUI1H5LFznW86zJMx7bgZ1VYDy1ooxI9oGLXDPz
a62reziZzZFHWqJmdIayT1/bzlW4GjDflfsxW93arRSVXR1Feztf8/lMPXvHJqxuY2v9z8kArCGl
PNFhNoBCPy+9y5+j/4mqr2tsBe1V+jioze5d3yfLRT7wJA7XF5DOReTpONsRCZAgj+7vqJ0iC7hA
ye8JoE6g6fIt/kYghUbh6rZaJqy9sX5KZ9yAZ+yRUm1ME0spLp9oNdT3x3h0IZ3BAWr0GpKbilqU
ZBEB2dyqCfMjv8NJyBPVTt97X3y5MGnzuc97q4mVsFwxGp70j8gtWRPMRzgSH3xzEYAXE8KESaRO
wfHzFoi+cDU4RfNoUVE5Yg5F1/6zadmNMtibkx8p3qI/J3ClbhOm9UtIPzFuwPJwxTiAqFU2G+vu
eRRjAIWYcdNTvXsm3xvLzR0Lhiu1b5+WauilOc/JqnfvOaEl6I9iqLsnkcu4j+RBh7ysum6RjPDf
uEgWZ1jy5pQJnL6l5jHF79SsuD1bo+wNoaXPO6hkEMhbF/YmuFhIC+jxlR7CFO0g8fv1bwZ8IMha
4Yr7L8ge2RgFoy01Bq0ma5H1FQBA0imYKTXWSpugAIMYtn4fKATpZlpQanCfQbanv7MMKHYQM/UQ
iucpecQlsCVMefhIktNo9YgK9ernGZif99F2WtWGv17sIRrYzd6b6QPSaenAX6mZD8Yp3nH4Xr5D
Q2N+YUjKWwL6glc2jKALQ145TXXT/hohFVkVYaiJeG0UtGBOOy3LNAEc0L0zRsAtEeRawssiIVbi
OyhnbwYly0OadfcJA8IUwhg3GdtIABKhBycKxkYH9zUvoNlIGUy269WtOxBLNefrtkM2IAWsaMLR
xh3a8tizIbTGHRcCQWe6wxHY0hfwAE6P4MRb7W3v36m0A7i+eoE5j4VwdUVJZ/MHxz1QO+4Ncayd
icZX3WYfIVu0P2vTwaHXgDfOw3PHdpzBC6B+JHxo4FasDdZl1r4YZD8K3Ro6ZB0IFZULbbz6YQfe
1GUYwqTyU8JdstAy+JDuzKWRd1SRRUWqGbqcG+zLYt2qCusUkcg6kQ+snbhGdIdcxN1dNthFHWrI
vDBQPMOof9QglOmj6NobNj/uVuKH73OkeAqEYnFwdMzDoHS00sJkUjFdef03TxpAF2USr9YibstA
zpIQU/Axnca0SokQEFTPcJFtdT0/qKvJwJOhuZxZhbSNMLdgnYPRT1WPU6MJHIx6HayyITz0SRjp
t9bBAYIoPxO7oo/P/Ya1pE9WvAYZf1gvHoNKtWetksjT1mrwz1yD+hWiflsatTW2ibd5YPmr+Rgy
0VU7QR9KAK5Lxd13ZUimTGDU1cGMzCJoDMIXYukFii7SJmgW99LPjPhUBlvpwLpHb71tAtX12hEI
3Rw82ZnBDaEeHWM9f93Oh+jqNH7XL4Pa8gfkhhUsfXY9sNEpD+lI4Yc6YDWELH0MQ3HO5v1zo4sE
0xb08j633buF70AZycun8wBzyLQp9CBBZODLFeWrbUu+Uy8pLMhPBtU9mWTwkyl4MG4Wq3WpQgf7
6GjeyqlIiDc3sVQXJeu0P4zXrNI153AKioVxpYm02Zj6P+niMQjtcnWtHa46R4ArewTfCFrfeyl0
vZV6BR3PYd9BHeSqIVr2pA1bSBbzitUPSoF37r0VbKXs7DnE8hr3+Q64OsKxgN1084T8AM16u1pj
WzqMwgYbmYY6JcuAl/UwVHSQhvfA3ar0rKmZT5mvhXufpG6ek8Xm43iogakLVgzCO0CPGwZe0T5P
vUXEdo18PLMKQRmZFTPalhsXxN7LE8l/TrLDuDTxPeBi6FHbAOFr4tLFxgPMOiJ7ZaYpsk1DrKb/
RxMpa2OP2MVRIXInVVav5xMwGGTJquXHIWL7MI/2LptXboV8qae1idZs0TsqJNF8RyY898XD7iXD
Eu2WVSBgBmD8MjbytI+0TzO/ikWvE/STlc37AOUvbN70magZQbdysK68xdFhevSNHBi9kvkTK3aZ
wWUTZaBEXugdcYj1kQx0OPj7go7q5Xq2kOY1JgsM/vz890C2BmhxtlSVPab5MwTTIfU5l9UIXCfP
9tGjX5d1WnUcobbhK81sgZAbE7CWgjhrfEXKG+lh6HIJWPajjXlLkhiT/Q7hMLjkCtQgnknbfd88
+v/SRevq4v6sV46T3LA/gnOSeAzHPMj6xhA1rg/aD8pkDifU44bFSvq71yvhbt7giBsBmGl0kMoB
KKeTngQW+Cd+Ka2K4NhoBXWzr0vphAsaEEz1jjIPefFY2U2B/qtEeeI1V7R06LZh2ObKZ0dv/kTj
+v/LvdzQ7xz3L9wn1TLosPU18NcYJHOXh4tL2//RNiO3mU8hiB0vcljCzqd4oNWcCR4bZUUnMed8
Y0wol2u1EckIeANoxPneWPUnf97YdsqDlqrd5iKeJLS5+3gF3ZPnZQn2Mtceu2U6hj4U3829Rb1A
6GolOjKXSmevc9rz+MBUxmAf5au28XW9/GFqJfXeOE34V8i0E64IqXtWaSDWiQwZG3qgotWZ1H7W
EzeTEZyFbySU9dYw5AW2ljsKOAK6DIyRGnH8Ns/eYK2aos8qcRsoU0vqkyemxQwxyGZMykeg3DBw
Tz44Z/4q7ltSzLf+EX3377GGRRXVSJzpV742CMe/+M22GMSHtHkpQbgauT7AHnJfdvIVMeqhKb6V
/mk+uIgFjHgqBbkLWClPXsW4W/vh3NIuqmCyx+1wgbJyLFyfQ+JNIs3nOpDY6YHFhl/g/jxQIYeg
XMAV4EzP+MZjPdCyHQGy2SKd8EaM57BPslhAEMnZdXt6V6xCkpw7O4Lr6AC6ujBDwXYpl52zQD/y
KLhR91dqSBWfLQ1oF0bJpx4ryHQFtgr/DdHIApMmo2GixZFl7TIm2xk7i3gs93GmrdP96swMlUs4
+VSaLy0hneiryzijR1uhO1l0glnPcoS1HcKenCcvPMn1fvOI9FMmo2Epek+u5xchCpm8r7H0/ABz
plnHKgggn9v+nYjMZEbxqSDRhd8rDRRzsuRP/N/Amf7a+WQXnFEcMc/mIYkXnj+yXjrclYqFmE2V
l1iPSHTMT3Cwky5j1Hcd3AAOHuL30hbTeGwIH+QKl21POvoeZOcERGkU9029CQzkK0rqYlqDuIdr
l4hN8cXg19ofL109CKX6W2RSxbOWbg0HxuhjPW4CAu+SVC1oB17FOTsyWAL1OS1FXi9xBBLJXC3R
PdYL4cchZ7ns/IW+QJT+e1jMXgpb4GVuoddMhR8i1QhcR2PV5c2bgqFyoIUUlUxWJjJeIMhlhhAB
xD4wDRMgWMBU9+q68SThMemv0LMzCrZWHecMcJt+mlFQB8kZUFIONlb9fOeJbXaTcQ4X0reuuQGS
cP9WUX5Ob6jtt2pAytoKUxKqDtlFMl27JCwHUO6LZ0IkCcZuS2MgvuvJ63RVHQpkCVoL98zNhoW0
o1ghte9nDzJnRVjN44EeMDsU933Y8bQUFK7EzprjtDxfWMRLvWCvPXuRlByjjkGhnCxlA8ndtW4T
Jq3js0mc49DxyFbAwzTs/5RWIpLxOb2ywb+GH+Oq83LbBQRVzp2wyHbYvl8RdTXB+pdYU8TErdkp
roqyv4cd6EwHh4h5w7BuX00e3CzFB3ZGi+1D2R2okV+4tFaG5D4ay9aX1TNE0lmr5pTTjMRhX3Ol
QtalsUvbTLDO+lXM7JwORJylf7aP9yA0CvlVoigilXb15xDJfw3bmgBcqJCFF6vsBVw2g1GWYDnF
U5frlmDlbKOvyid7s/I3jT4odkx3jvpYIBpimmVFbVZZZu/Gl4Iv39UtVKojiOqdb3eVjL9J9LDR
iyBuJMlMIy2PZRS/e2U5WeWKmH79CZeHzp+/GDdDUvMB/6v8LWfQPdXf7x04uEZjRT5ighVeQq7a
6x4pl/rnXaQ5QSj/g/DD6dv+WLKkUjWm6/Gd0BneNdYxyitbhmCEDEfIHJv/EDHHUDGfTPXflEgu
PoygqASZnCBZQ0ggniXxXvFkoWn2s03yapcV5CusjDRq7/DKnmCm5Eu5WENNEnklFVQpALfylQ2G
r82xu4/xz3IPJokKEitsxe0eJSANlHG8KTl8Sqy+locGJSQX/v2iZWzMwfE0unfnE/gbE6jtR2Fc
MYGip4SgaVLekhBTLCM4z2tm5uo/7PF1J6ExkfAY6WUv5M5ZM6RiR8koZO5zRrFSUeGdT3+gYUFk
hsCf+6x4nbXg/L97cN4OHOcK/tCJwxtCs/b450f7qNyHReFr/Og2viqSGl6lkLorc/kN3NJGMu+O
qKuAxcW6pnquEYG3pOeh0kCaabkTBsbxVGQTwexredKlblNXeGMNpxrTXXv444rxoc+dZACMt/Ld
Ghz/nPD5VJZrp26WD927ahDHPTjcIUzE7t/cB9/XRLISgX3JeaMfhmfz1mFpfS9MLIQwMJ1QOFE/
l12QP5sWMFAaqRHdFAN1PT6T0wrNmFM6b6KQrx2pfu2HRoI0RdMj5zHj8llbZ2mGidNXtV0pR6qs
b7DtKFe7dvg1Wbggf8wxfhY/Y9Y1Jnmf8teCPnK+xxfkYvR/jHwxup3nTQQAdaOuwlINmr4MgMc7
N5ev4OgA34lAHxGUvWgRhkIOF0o/IEhsTBxgUl2PBB2eAx0g/+CQiQ0wx2wua32GqhQ2woOA/mDs
3fNAAA1V3f9gh1i71ArJ79+H66OiYIfSR5eJOrOP5VIm16/A2Qq1vhMGRefjvbPn6tJy6CZCV6iH
qDYyL1+THdW+T6DGgxJRcdKM5txo8U8Oy90niW6+h0620L5AFFxHT9235XFqmjlXpQtuPDjGsLRH
RNlSutc+vAQdxSZJL28Scu6+uLYT3LP7qU5nRo9O67b+0ZHmIlwengbgkklUogsk9xQ5kWYOjand
jXZWzCAlweImvMCxsx1zuIDSuvOrhpM+6VtsSSHlqbH2PGewBIDjZY3jAKyAUbJZGxzzkAM7xyu5
AJU5XEii3MzoTClS3vgaRyTIrztykc9k0vT8OBGgCpXbQiBU0ELs8lN1KgW3gxNKRkxxoOOxV+ws
DidsV4P60Occzg8i8A4vD/WMKV2VCKQoMIODoN+/5f7vGNgu+auGUlG41j8YuoAYo4xXP64zeRvh
AmU2y93wHGa7ALC/bw5G+OSeCw2tlTQ+FJNqnG5Q/LsGwqNBiXVEUKft9JaUTFiH0aHGDX0jQOVA
LILViyE9GngEIRoxkoHIGicwWuaelfVrzRVfjZ+HHKld7O2cf9kH7aKkSwZK3v4BO/FkVAFQbbvx
X8t5tqMEzdkulfatLdjKVpuYJor2X9yp37DkBvgRq+c3OBVHJUhGC1zCoFne4L3jkSRMvldO25ox
WbbchsLSWxJQGkCoHWcxwigyLyWR/NPnfo2P6epv/VXQKg8y812VgaCj2NUAjwXO/6/Spnwa26cb
8SvYxidr03Cw7gOc5B4WVlhPFEISof2d9O8Udv+nr8a249usq4/H6RLGHKQyqX3QyFWmPU2ttrQy
PM8Z7Y7rmquFeGbf49gdTJwC/Ugc6HopNHZNc2g1rQdASeNJOiOLwe0VI3Jd/6KCQTRpLvykejke
xW72kCF01WjjjWx5OZ/Bn55uY+eThKBgy+bqyrw81ntJ4yFthSShDSCd5oywSipxJtDMnSGcyj/W
/pIFTLZkClA5+HOajI+VL1hmbfVe+ejTxHrTH5WzX+RyXHvF3CHUZIk1NMEVTx8NKGE3mO/EDLaP
ypKVP9Tl7CKBOaNJp4ns3sS3Abao+FjLSD3XkOpfJOPw32jJp152fGCyS/letL4jQKaw1GbivEWy
Rs4jgsEbuXDU70cFU/IDpw+5Gsl3fEDrI2wfnSwwBDfrzGsy7/MZpk/GoBUu6ixOgeFu4Pk3wppl
JOzXzh9Aqe0Jg+8yjRSLtpeTga8hzyLr6I3RRFvg3jz56XEeZoAd5Kt7N56ufzV5yQRo6FYfhIA4
xHMpiR5l3Sl+B5LiStR7s6XE/EgfajsxgI8tdl3SomJqwM9lG/Ba7oddqLy/fnHGLZ4NiSUp4oAB
W4AQkVlOC4aW2FPW3mO40Z+YzqPD8sbn7lklhhvRtQQUFHHdU7u+jCTE2yTR+vMHeVg9eKYKbHCO
+zI+4nQsHc6kBo9Cnm7mB0X+qsJ1ah9LSC6a718hPkzXBXxQkavcEKcimtnZep+wXpACVkU1njc/
Bdsb8+gprs69lfgrDa5FN3Mgu5C4tUT473Evr0GfF7dK7DlkXha++rXaKrMqiAwog/AaXWBlcMdi
5BNiRPqdD+Cx8IhSkUVIso4gCsVfETtmuKdxssxRqaitfbSzQcrXl+eW81ZbgBn8ysJ+DX5HADbQ
Dnpy0NmI0jhArHQZYoH0awfM5KATntWrHIeC0LTB8ZAcknSeWRxDJGen5cfwE95OEdmCTgMMQjfX
WAYrHOV35JlcGhx6GiKcRcVO/iEO2qW6MnYhW2CtNiZGwuxMrZxuw5UQ8VNNK7AkNgYEo7qOFoB/
GQgYX2o+sO9f0nu5IgezyC8TAoOhLRneW9jfjPQjirfXBQsdSpL1ILN6SpK5QtYvFgtECkOIRM3z
v9wvpVPKJziFpOWQ5T/+Cl3Slp/LSlrEfsk3SmuVyBA9QrX+/l3bGQ73StCFxnZnzMP0uaOVuy7P
B+WPgnXhdsCom6odWI5eOMmuv+DnJHttQHciEZHePCfjOrsfRlqnH0ceaxIhE8nnlSGbEKNI9hXr
IdvBrIWtcqiYqrE/aSN5gJwJi4odvbt/R5ffrrRd/Umd9bSdUt7JZDu8ANXYciLTMcrOuQS80HqM
CwS7ticqKeP55X1+ucgNY48M3pnF3n1+qKVG+rbwiadtp1Ysf746THwuJcTjl4Da1jno7hRlw2/8
Ig2s6RRj+AWTQ6O7uvbnTUJnSLbEZedGnj6PzmAV7t9kEfZUTv6wlxd8rRKlsAGt5Z57FdOApNl0
9/iLVJem77voGwsVq7hhigAM5ERnF/FyPLNUhjj4XFZJ5ppIxeqvmyPoAra2afMuZ5+xNcuJp11a
gVw5JisqG327Ew1Jvrl08wjeISOeQZIA5TYnvjAZwye3TV6evhyQ6ezoZ80fKUzdx//1H0If5wlQ
RRn5lHL0wB252bMfCPdj1ydq9/v5ntowoQOg09Dp6zFr83b6UqJhLSeEUp+//3xkxpWEEEJ28TG4
BiG32OWFy3SnWgD0qqZ2RDip2bvj4NMBClJ0jrRKyg79Lx536qiw1UKot8I7/ZXAefWOFo1PUlcU
A3btw+G0ADerJjjN2zjKDSFLiMo41H5kyENI6740ORBt86RRV36p6QmLVFVMuYDs24Y98c29S6kM
9mcBuVrs/5YehJVWlncMRhQXIEZZwmAp2EF51RrgXoQXRQAOJ3sUDFs2778U46P4etBzMvShfJ7w
u2wIy/5p1b8LJW1v3f7ZNlZHTCTXkXyYe9lA5RA6o2e/hRysLAU4tE83Et6wy525p0o40hm3ZE9m
yQP2KpUJHVNhD+wwseQoefu3J4LAxWkhoB4zOaGP9VX8//DdC55CaBQjJfupWu4ayjsuBXoyjVMx
dSweAVIpRY79nIoEK3vUzE9RgkoE8gYs5C6o+IhKAhgi6DPI8njydAsO5RYBl+NbekpS+HzRgvyu
NzYpZdCqatC7DSoc37YAGMlKr6EcDPdIiJzCsgYXzaivfqlLi00j8/SZzJWuRJYe3oRMC4NVftKd
h8yD5GT6tCi25y3LBuf1i0SmlncleS2JQ+FmmLvtpfIbUhzQe4MxCFPIRIsAlqBNseq/gIoxAknN
j7gEm42pGAkJfPe9bwa3TIU0zr6mLPf6O0lX8ICyUsWONYPNi8EKGDwnW59UD7k1U6NdUrIs4F9y
AcIot1qbTn/P5r9/esh3rPcu0eWdgaKuVINpkOgnS8jJQj2rcBgsNr1tvkzXb7NJSMtrpFuC3i+w
6otFrrvwgvfhfzkxWrgBG6VCopOdx4dn0UlvW0kZ5ceg8vYBwZI1HmM24g/XJr9H08trJ5OSxoQH
1J4i1DG0i6eBzfsp2PRAZRo8ftP6mT7nf+TO00dRibiya89s/UpIu+h4ARKsnv1R2Cl1HxouvhKg
xHAzYWicC6t8pMWFJct4gJtzG37memNkTAwTcmVJ1kASa87Vqqjs0MxhNl3JQucBcAdRfwfX1ojt
jOlMCLfJHe/2GnhbfhXhRw8pMtpq3Z4r/L7dWmLpVZSysC6Z9qePW5ifohAhv6X8KL+mHmwSsENx
twjttlxMWuZ0XJloKg5kpEj/aAlz6vdMOOql0zRd2wcjmiHxlGTIBef+13nS6BwVj52CloYrp197
/+/5xVU/P1TvfDoK9T0LfqJJ4kVJa7AIiT3v6gMKw/b3z9WeybAE4KqHjMCV2OpwkF9NZdfhzYIX
Ups5fRjhiNDiPF55rdgzjIV22iD4F3FaLY6Du6V19QHhZqX6zQnM6wezOjM0imhwcBO6rCl2hnwI
oyjd4gW4yyzgaZwcodRk4h62TJ0stpjLTBbjNMvspavT8GPm6DOtNRfpeikhp1cdcASs3op/B0Hm
4aeE8qJLDnnvW3B7X02g08IRGYv3kv4Vw9pRJB9knYG+3Jx8TOr2eVTdbv7MOr4ZD9wwTZsMfNnR
MXiS4uqre3eiOt/aR/fFRVK2mozirvhGWvllrOD1uCjCy0jNlp0yubt5fMMq19CqfhLgEgR1BvQT
bIXje/Iy4TkN7Sx6yuuyNUtDxHdlRbIbirEyHPT1KVsQBSim49MMOC3TZ6BIHnbGxOGvS851+Oqk
2VTRdqKxY68CFWnRgX8L9qaL9q0/HYxK6CecIGFemXsE9PQzyH1gqiCSRnkUIQWTmYsngv1twx5N
3pwY6Vix9brRnjaeiDGo04exyR7/3lGVoAHgZok180vPJPPXZ81bGa1aubw2T2mLDCtTR7j3FsnP
4t6bOzBtdqkUrFSGu86vwpVxJ47gI/lYcAENA19sGt4v5O32oEjZ/aSW93ieV6hZIXvZZYVa+DFF
Cd/fdfgiOjDqv+wxhkm8PfMy5hFVAU0rJXcp09+iFsCf33rrR4zKIW1sIkFVkG8cK97En6r1He1I
36hHQzffXCS4z0hsjYT3bXy+ZcPR6LYyCrrU+QK24Y77sArfw/AcHLfHIhgVbFmMekyprQpWZg/h
eeLi692DsjWPO1649t4qfsrPmH9FfRA5/Kok3RAhoH6JKBxTyuWhdT/TQwNBIjtAovISMCEz5KEW
verxfxqvmCAPNdWrqmMCDqRkG1XLOtN3UTdcd1IXpqSR1P8FbTdK0g6ooDvVxQgHJejR4g5B0+qX
vAKbonHUm3Isv/bUh/JVccp0cGwXxJmY7AUG1+8IY/rmTjU/NiH8iQmHYkSuDEzdGAAEexmCnCQ9
HPyV3jhkJQN5R2ekTH+iHRFOY1tmOdt+VJOFrFquXbeiJu3gE6jOh9o0FeSvu0odna31cHsYh/qs
BrdadyWDulqFPpbDgylmWnv/GL2QnEzDXJfQmehZqxjY2PS5OlwXHhw35bY7d3DW0MdArY2VnorU
6ymLtNRce3mWbEQUtgMlLTIDIrM397klDByj3m1BWCeQCUvb8HRXXYQ1lw/FSpI9z5Js+Ggv/IUD
kIIJ4lBhtKqa+Skrv/f25mDLmuByezWnwJPmCJ1YOl3Ufxz7qQj9MtprDgfqDBj7CTkVUF10qzzi
SBer03ptj5my+bfoj0Lw4zZ9x0tJTEm2blEqOPc7k91Hs+23R17POJxpQU9fQXAjcS+6jc5spngw
K2mAumPKDZZiDouOpuiuW0vLGqZGQR7o924zIU5904OfxmP/yZ72dOcIWa21Z9wwDiye6tvvvhSU
RBCN6w+nOYWs6SXCU0M4acSVGPEcGTIzxJ1M1i+icPONjqArheaLM/KYvtKbHd5gNhRzMcsYg7Wd
/S/jW1yiJr659XD4gxeXvAnp9iOeeTQ0UOvySk8H3VteVTDE67bbmVF/uxkrivIFzCL/U10pA9G4
N9v7V/27dCFpwTDrcbjF2CqFCLmaC9f9M1gjqA/pPzOfKYqC36pGohvbtQGEVvz3Hs1+QgvNwS2G
LNJkGpPDKTCBkKfGKrnWnAWYrq3ZkXnwsM/Jc4iv0M2oVRS0hWUV/6p1Lgzz46a9Q9vor8jVk6Sj
PIqrOFtQgv3xSLDsFueb0imF9FHfS040uq/vWzVAqf4RTyFmrb6z3h8HXVvW1L+JX9QZvaOYWuVQ
ZlTM7/UDcv5EP4IjxiblDQ41YgrcA/HZEzc1bcgMZDD4rP1bhjPp8c3VNR79wTviBhybE6ETcilD
4cUMTVd75cE+siPLqFOTL3pQIpny0is8wTjRYnpqsW8cSbCMIqmggKAeWnLBRpZy1xcJNcUcDuD1
PQPwPsrVnaqFXpkgbZc431eoFp3vW8l1yC+d/LpZYu0hWEvMTH6uIU66cSzh7OA3ZZfYVkPfNAov
bpWzeI8iRtnNj5gdHhyWkuyr1DKKuIplwukGgmQx8/uyrvrCc1Ycla5Yi2dSainIKd8CD6TUueQt
LmfaBHcGciWgoFoPL3Q4neAATfKD7XddlgfkkiMYEId7E8EhpeyPriM59v+eagb8zKRVKyFfjW/C
1kLtuhow69RDxokzG19eefmGQui6I2AbKxqs/oQqZ1zrAw0cG6zvHgU7331CtWsxxND/R918qTm0
xDoMpa+iUqSrBK8zMAFrNx1Qtlm1RtBd9VaaoFsQutm2bvedqqJT1XGXmal5v8od1JVxOtk2ORaU
3zenwDwsgGPk5grU6iCWvpqzxYaFO6YByXNJ0NI2IH0PvshzSZdgrdr37Etb2m7ABNgYEMozi9DN
/RYAvBBvU/Pg6XQ41QA00s6Uwu99UTVtxq9I5SaNiG+ja6xO79mPrAKC3eIgg9APJJ6rhnAvh58t
pcL1zWF+fXXNXJmVMX9bu/Nz1ktfRRRG6ub4WPupVXzlnjRx8SfIwctnoFFzvfdgumwsifRWWFD1
I4g2h7259Qjdw5rYgLAhcVqT/QdqaYXpaP/vA+ZPddERtlPxPFPinpKsruMUQQ7ZfUlxwi1uJKY7
XIah7AxmF+7R9SZWc0xXmYpQ4LPUxRG/Q31sCrskF+53UNxxvjFUphM6nY/ihLnQR3GdnXGg69HW
P5pD5tW9Vdg89bz4y0fdALs+v7S68IPby3+RftVs5maUWUj/zjoLeMKNmZ3uuzuVjFVmGoL6eAOr
eKGDXOORLBlVFgNxUwicKpMLxLXFQURJ+JqnIF1tvCH4383+S/kqi4Hx89ogo/0DFC7E5brvoeIu
/Ip749p8GYSweJETvoSbhTCG4Rz7kELgdiiOjWvMH3gWYHTbcKNQX1g9XPmt2Vv35ew/a0UMDx7Q
A07sFF2k01g4VaC+0I1hD1Zlvqt2dq5hpw7rkZ1HyXWSJcZWhEK2BoO19zH5iVASURCUe11oy7IG
lUTHJnlzNpDd6o713bMakTQgd1NGXu5g6+e2i9X4Rz0ySsSvKStI0YDRHPDmTdDPcNKHkt1dzpeJ
nbo4cahua8t9tQE6YE/SB6NvjGtJFUIpbSXzuv5Vu2DpTkvVQmvUsyJhy9ixqRrFugq4THOpHWuA
Bv3ELO9i0Xo1i4oOPxaIL4pTXHi35Mg0JPyOouOxQJRz76DdhNVYSE8uE61hGhwecTF5Xjgs1eWB
oDr6RpXNQ6xlqzBqSfQyinucbaiEa3Z2nFNa028KTVF+fHbskZ1ydI/mJgFnM/IeMaNCQ40e/TGp
Ek5XshxyIMdKya3WuVit1nvD6F8aRRCPzMG61Yf83rRZ4v7LDeog6ZvKjfXu6K0q/jZL60DSL1OM
gnOl3C3DysjB1JGTtHVMGNmlPv5fNRfvimYVhcbBOiUugTGNoN8UdWpZH4+GR2bsVdm632qgpfU4
rCHMVdumy3IP1s5N2Rp5Bdevnal3ICiSUzWxiHu6iDQtzduyIGpdPT6zSkkQvpusHUWKwf6rGX0A
5wGwTUskQmgrtSz/XOMLFLcfexJff4TTXyZ8sj9DkrGs2XIxuL2jWD5M7nVRFqBi0BfMDki3YP5+
1CT0DsFO22hooqCzT04Wpf2OeyMy68mA/8Bp6BB9vur0IVUn+TIZQnFPiEl9ZVejX9l/+jZEvQhz
NW4zAmlkanUiYnxqzI0tbQ+SJykChsVZLt/ohnKm8M2HxvVJulh9Qn6O9X5wMZgYU16Jzj0eKq9P
F7UIGwd66ndN8xjUHN6A59i0Xx4UGxwn6INiadV8petgUiR49JOzHvbKJOLAqUma95YwphtAjy3z
lV6dqSETiNtO5Oxdu5Jb2blS4+eodfdk3YNAL/4vTb3/YvFa3zXxJdSMFOF2yzlaeXCbG8SmfamP
oIFLuzkTrRAXbeEVZCU4lCjTFbvYyhbvyxSjtJymeuPYhHWL4rgHlxwK1lG+B7L6F0paJfizVQDM
uSsgI7fRuhhlekDT+HCu5qyvC2MPHzpfJqA9JBqgU3bltPaeq0wp3Q3J93nfS62kVkpY73RN43i6
XiMQKwrI0ZwFyN3e+Rksxdt69DInVcSnT6wBhWGFruH1XL+6K6T7YUPIhwSoHabC8KqdjIccxh5m
ExYhmrZ0GJ5njraTRUNTSxwG7+B3+GZZ8S2dgFcYIUvLKiQZYd0fcC8YZdO6QKFsblDW3RuSn7Er
c/gBF2AmjFjsvBEsQPt4AapRMx/m07xsKwQhVpE8X1Ffaqm4yhHILGIdoF3TLwr6MMYUUOJMRYDw
vQAnBwPD/mDfqRRiCMrbMwvaR48fwnOQXe754e5J5c6d6M20d2d56MFvRCd1sq7eY1FUPfRrSQmm
uUgD9sJyfN4jPyf+vI4gqmwqzKsQwsBaUyGxkIsZIlduDztqjs5O6qrpla2Y4HdAHyd5VYkEi4cO
XqFtiPJe95QE4P3XBrv54CIi38HlEzK6AvObBqY8wxLt0jPdfalQTmS6LkeuktvghWqnd+CSZl5O
H+BJEbhuKAhRzlAhqoMEPKFSbozcVrTAtUQnK01SeG42mSdJGM3nGoG8Zdtud2Z4oVbd2ptlFepp
ISe3lIKy/wCJKLTi0/dgkl7Yjd7vxUMQ3pyoG0RVwX+feO6I7TNwmtGVM7F4dS7glxLTtF3gZhFa
Zv3FR3a2O73xdxX6KZrFD8JBwP9W8wTc9bXB34EMpZHLbOJpoukPgDznW9QFnQDHirquCOuX6w2L
Wc/xj6knh1aF0mx9ARHGV7TwfNCD+xLCTgbfziXSmvicFys2CAB2ARdZFlX1ygTJEXxCVkZqaiyY
LBE4zylevgh1FVCzBBNrUjSfVf6/2/6p73v16SlvUxMcE7NP6UUYce+KsI7yXx8rJTLPe3D8j37/
UuvaNMcSReaxSNqwoc+JfHXrysIkw0e78lK9lEtFlYLRLtEfZGgaHmI+tGCNAbtzVD6nzJHCaNu9
B3PM9WUEPaV3DpHipiq/sS/8ceMfKRDoeFe9P28gSFWP1QBH5C7tTw+MNzf0iezlATynnUj7jX+I
np6odph0DtR1DIp5mAbCoYKsCDQjJa+fu1QUp5FjcYaX7yXm6jsmqfKCeFAgxNWQhUIVjB40QRp1
BxERRp+Gb00qm6JhxH3Oc4e7LaP4yk7abbrlm6awuPP8s1Z8KSgVaIKQa9nKR12VUKMejzTIIhCv
7GfK0HBcbmti13Momi/xTjzOZ/leKeajUhvRcfAtPeMa6EKSTOUePu9bRE7WB40S+tu1MffY4/i2
auozxqeJlipYslA2eXhv4/HqtjJEugxL1cQI2OuRvfYpjiUs1FSZtrrGxNtk2f016K1SfVdLTYms
OdePJhU6EaLJVU0qOmagHFO5XCoSWPYprrKJRt3Oy+ACJGr5BG+XXK6zWQs+QMz+8/1JFrcxOd+l
cznvP8IAO66Zu9Q+OwKrLrVrNAs8vMihc9T6eZ5h4m9WcSPF/WlzGG5B+shqAYrtQUR2IRdYFLaK
FD4VudKb9y8yen+Af+E8V2e3i3TxyYowhwaOunSnD1lE0UA5S5ZF9qZoKqW9/NbYXlzFJFjw3Wto
NotUboLa+I0ZNmD6viTL9lQFerCsG/8pG99Dmx21owzwh1AcurHdeqqufdSHdZHV7SQf1P9MfoK+
0mSuhPyh9HitearxgnIW3MFhfTtweD0yQ58wVweP7A+9Tc/X6k/pTrlmTXIZMnHHV0e3rkFaJAfb
QC2Tett89e4Y2MpLKSJEl8oEvkcYdgah/KrD8ANXMpk2zselmUIbs6IrXbVoJyN6iFv5rnTIIAfo
sPUpTYuY/9lo8hyyWUdhs7L0YeHAjoaqncoCvWBHTdN531Iw8dLDZsyszpqy+JTG7o3W1KfEMhz8
5PalJJYyL5NeMs40Hus8dIbegUXF7AwrRZrZxKiEa9oKLcYEwErf0p4jeLXPHgrTvq2TqHoj2XA9
VbHaSvidAgQ4cf0ArsbajrgmUNF+CGa0+Y4jh/y8zd54bAQhH2YACmIwtODhYoefwx5sh9quBrLF
mhlRQdpr047x844AsFxPzwQQplLYuXXPD9MYgzHqlReyxvXmok2QsCY2oBxI9EpVpfPGG/u2IQ9B
W+11V89IaIiSQR+cU2cR5mN3U4METsTfb23U0/9PMQI6SGGNPuhVQSjlGwHOK1JDfdtY43jIMQo/
Z+w6GKaARlejKL3d8ME0BXsG39FvVpxqLYYjq4RAphry0onehJZVu3FYOzFz3YX6kTU7enyiZOZw
OfkUuZWiiC9qB/LJJrf8pUt5no78Yg/Ee7+icslcpVPvpY5+zSVMkh2+ZnOmxf9uLEQqsuClGc+x
jh5vJOMp3LxD2sc09fa4NVkWcsRlIddmDOSdIvBQ8H9QwFk17fIQSvO01kTk2FBbYD9GWLgzfVa0
UZkBH1KZSnW10g1xn7Ta2jIxRbI8IZ9fu5N6pHbCbGa/sJpPn31Gh+tBoJ6N2mEwMAd2WqYbm09x
acy6WbbjEmxdoTg4DDEirfS1v1tjAX6C/oaix4hB2p9Z6OJrCNT8eLebLaFKUkq+qpovnLJZexJj
+XrzqjBSepJu3HbAJzVNcqM79n0R7DvSblqFvZ6hpo53s6aXxXPJEnaaZu7acW2tVHbXJB//LBqZ
Sgi3EDmAGlrM1GuH3ISW6T3MZMEzhfSkuXO8s8L3qj8FbgQmktU0d0IYrbzJgNe7jjuP5L+ttbZy
NX83xuKyAP1Mf1ULCCzkhuqozjG2UNGQhCjxn4XpVMxlaZ51IE1C9C3+m7DvkPn0ZI3d38ad/Jc3
7eJ5v696kctDUHd2NCdTaJ16SjBnyf82Kw3NEqrYRSLdNXdPARB8oahWR6vU62Ji8N1PhK8KqzqS
Xourd72ikY3Xqvmz7fe50cZWZuBAWV9nOLSkXtIbs+Efj21Nm5iRh2QBUpE0uP2yLZXIY9j8team
aTI2lRYk0PksWBDwTAXQ/pn6kfFJZGle1eZdN40vgR33BwYmF2dU12O4bZfGlibfgRYMc2se0QOC
zV/hbtxw8IPgr4b58CIasCZoGiUJio9DzGpnHFw1Jc5qcHok0aDisJfFyucne7c4/1aUEeloS4ZM
IxDeTIhS+M95DQwstR1OCwjK+jm0HI6NNrv8MPwhIE47BxopyodzuMmJkrzj4gdATdE28jNVpWMu
5QwNlVxV0Vqc8qlJ4mnN4ysdnemmNHSDkPnih2O0JK+L3gRZX4rS2rY61jN7noIC/G2/fAXXlplm
FmQd7d/r33O2g1LNRzniTV/GDxKzpUSSfI7B4ecrHxqvQfMIrSUhjkOAvy0JnebLBH83krMjV9RN
DP3MacKg1C8/qRJRhd0ogFNHYixUKCJ8vl2FhhlmFCvKptsOmldUx2mLyonX8q7NPob+hYRoG7CC
1PAIrRpLvcJcnHstKHrAwt0uiR89AXXKADvvlgDb3ChUYgVacu197vWqxCPaQsIa7nLWTZlh2sit
6xQqK25f71uIRnVbJ2Mt1OYuevYU4iDDHlts44Nk7y/rReKPY9OUofEbAOJKDvP4pFbpFKA6+6yW
YbqA4gkeRehSSHd1YKooNoWlKwPPp7z24ZpUs1JGHwN8JnEtXsJ+Z0K/1u72vmrzexV1kqPvMLGa
4ZBtWMwCG3io9GbFoBDL6wZeORlAloP8WcCb+/Dp8MjN5fRXNvsjQMZAOrcUOHftlIdMzz13qIwj
Vct9m+p5M0SoP6/DtWKjcLSwLjplJoJ2RDsoS2/wYiG2VmNUfrjTg26llL0HLt+fPIKU0PYlTL/L
6EMZyhuchRLoL2gQkPTuxMUQJqSDtWAqsYYuzfKzGCckj0LxghxHHmfBCGGk7QqTzQKX0372dZDb
7E8l15ZkIj4vGy1p0b8ErmD0J7UN3rlurkcK1PNWUiadJsZZW2sYJp7VLsObc7ilIkEYKd7lPpE8
I0o7a+6Iuj5MDcE4D3T38SDrSHXdP0rxoPuZkaVvKvlZnOjf9+vPUdXweGnsuQvDP7Th/tPJZzfw
GXTKKHYkBjDW88gIdDIGOLC5e34Xitp3ExWI+EqCRqZJEpOmHdKeGHzlFCxxKlsIDED2XjT258fL
Z/6BpJe/h/2IoYX9RpQyA4+ddmbI75esmTXPNC4m01jglU+S89p06NMzXjYnwVV1FkspNEmcH83B
pyAr/6vPQLu6I45GtSNSTS2PJtE0c/s4EQ2J3C83LNRzl/2OSZ2bVZFhf0ud2HIRhkuA8aKxuguW
NbibrUtEA6yWB0/etE41bcm9L4zl9LIixncuzkjdLuqdzaj0orcC40TEYGBBBYj0E9cEbtMUy/Hq
1T+zGjHR1pGzZV9LetzLxM6WWDbadaTfI2zJIfcC5GFdJrsozo/vc/cpQquOYNklUKLLoHeDn2bu
lPI4VZjLyh9AWkppOYqVK6dhkBJ4jwgW6CElxUMjiJxpTOczHaq0lIK9kwiAPBQsE3TKHXUfIYOZ
POjO7ERZ0Ym/5hhJqovtTwSLaA/RR8D3EJcfUbcxHC4fIcJBNAjUxigr5CNuIQl2nzpRDvokjGHT
44SakmG0Czey/vPSyRDy/JcUEnKggeACGMUEe/mY3n0XAanwtT05PCISWxmS7dBDZQxazPVv4qjN
wxcXNFG6uP3652m8Zm5je8ZuNwSIIBsFDKn3hLs1sX+I7MlY9OOIsYLhzurMPDOwYaakyMu4PTF3
UgAV4d3ni5aKS0jqEhzC+sff2votjWT5IPjLOGXcUxqilzQpalwWLtbcTcOswPXojdjwBGTv8KBs
0ELIx74p0qE7m3aYHpaiwFpHwa5vemQyb9ZOOYWJkdkA1XUu//OQbqlFNMfPQfIoiNwGLgHsMsK7
yXk2qXw4yugZSCdGxi6Ptga82I7oyIL9lxD5OyKM0jZiFiMI+ISEUxhV4iWVT54L2V6G2LEDl6w5
nbEo5Myyx6UascE1im95yv+3/1gcGz4Mr84lH8XNvXu85fWN2Xxh3AF0HK0GU7vPUu9qiEl/14bh
jXGSMn8VHw9kpOuOIE2TJsFSIzFygBDaPyi4Uam+6RxEHzAMtrsZe7QOei8uKbC9A6McByVY922b
QkQHONnBedhV3gj6Uejb68aA1YxCjNKiCNCUgkVllDTZzm5hrmchB41M9EGeGQnUoIeJZYFFUrce
WGv2Q0Ts9mxWvCpAzX1JqQG1GEfsSd4Xuur47oLoCZels84sxmBPNC0Tu37aP1EYQ3LKnaj9/EuT
CT6nxayGLY5WD2OgOGu1QWNm0c5hsQ4JlhGYayId+RTTmtxBh8fKyamwPKehLvTj/1TZB0Iw3h9m
guoKU8TGKOPfPcDIg2UDVASkWmvIAXbqSenQU+9qH8ITayNL8pLNSR7iVAhOCFXGVBe9aYEzDF2p
JIo5au+pEGnTFJOnGiIY9OTDgg9ZyeHDTRmrLa7VWMHWdbEDv49KHMwRkHysj2Ztob/mL543Imjx
8BNiRQQ20rMhEonegzxavZZpNOH6aBWwdtZ1AGP6OE8sWDLPCA6HKTgCXfuYnnCPkSYN0bLxOrA+
PfkbXDtnxgccCP/u+Ly804Ap7qL8bp4Hes2eSEsq7ZhHKhPc6xHt8IQDEtdjNEqoZnJwAWkWId24
LcVjzS0QUEkwIRd9LjzNOJjObyVFeoU3ZLdGxCchXiYjOHa2cE1uTBzzX5qI6EDPnvxSHOSjqQaP
caoqNugy/LxFI2twC9iVf+o/8u/J/xd670Gi/vsU8pNJNw+r9gydcxHr7awSUK/nnoIsu8/KqWcC
btXyw56Yu5yOnbuP9hxbJ/C3emSlXhWQJh4e9zbzgXzoqb9bu/PctomTWzZjMJMWnyryiMRBUOss
6M1syAcflrfOqJVOfPjD4sBmKMNU/hXMN2T83CTT0jGiwA17LxnQe1QWgrONo6mUerh5p99LTEEP
semKyH+MFEpwo99nbUs6MDO6iQmhsQRcGDEDFaHROM3Nzbg4F57FP134d/jL+pnEsyivCd18MKvq
jXEya0ErBKeougIlDsx3zL3slqmo6u3eya6KQKL6d2OGi0AdIruW52VBWoGAJEqC1j7QzrsEmFCb
Z/HydXSR4ztuwr6tkY+3/BzU0NIDkQU+duLMsG7VG9hz4ux08L4XBd2T69hIoqhQFLaBH1sYJyNe
oUdUnI9lYCycrVj01N83JCGKbs9DZYctlRRYwN9Evdp0IoHQ6G84F+dneMTtSQqmmqk/nB+RuwJA
U3KbZnQvRPiemomu1ruyl5WNsGLU8kQNcBAsQ7ZflKP/kGKTMr3oFnQdNw3G+uifmANnp8Bp1HDR
ppWHel50YiPAqg6n63K/y4zFWPB2SUAxPSwOmMgMUqnc4lpHBSwTK77yUgXmP+MPMqeVDW4HBTNS
ZK3XEd2aiiqgUAITDdm4AaZxVTx0lakb2KaMV0MpxiZfx/zvukUcrdzQbFZRR9XOy+dS3Tk3HfQ/
iaqG7hHtwPhP6jXs59kYpFEbq6Aye3hqxiExSYcNDoz0j/8K4i7N9E7D3HvVstUlGQb9dctjSRJS
bm5HjLeY9kBv+0gQrY6VbDZ35xSw+hFDl+1jTq0BN9la7/QmGHbb6J/tRbbsBqjLsaiNXhL6RCMB
xsej/TtBlLVBTP8EF+9wRiqyrXMF2+kJhQumOYIXPihfabY0hA+K8XiiPovJqT75OlZM00F4PyAF
MWkToPPjnp2mZe+0SU8hdp0bf7kmd8IIdOLpHO6P/VicuU5sWsUF6tsSVCp9kRIm031Wyq1MU5hr
YorZAWLRhY4s7AY8yD0XmiaQrnZEehFjpZpBPSzwCGevUjdr4WeLVBTUAVWA0RUxwNYq/bcrSq5g
Ex5saLIdSGI/i8Zr/7/NBhDNXgM+ROHCQmenS9Rv94RLC5wxRj/sfB8l96797Ah6ftqSLRFmdKyw
BntDdIwT/ZP8c/8CWp2Cmo+a4UTlG92WXhR6e3L6qAglH9ylm8DVN/WSlzGbhYpOPwEpkrFUdXY7
Od3k05+hRRlyP4HbUMXYM8huajjwwgtYKJ8l5Wxmn2mQdgf57RKY7Gw1XwWWBU3qf0+VA3x5PFU4
QeSM40BgOldr0IuhcdL2F639sjzA+bw4Bj9YMkhnzAYAP2+6tItx6NlViv4ma6gYFb9JFGsqt7k/
OrH/EBfedn1VAFr8tX/0bamr29losLIcdVh2AWDoTIe/BEDpm1wbxqGT1203AA5z4pxtzE0zHHZ9
0ZOAUKzoKFKRoPipN6zQHKW94dRyojE7VS3/QAeUofi2bFSWPHmWsN60vLAg2qUDYh794UgIFDfq
cg8LwOKQrYP5Ju5I139O2Ju55Nhid+r/cn+uHgA60Pa1WGvuutzHKI0VZQ68+fSINM/HtEG8gW+7
7SSuxEa2TkyyL+goDGWkwcz7cMbkhkthMuhYCVEPr0EoYBSvOPMe4Fmwn3DWpMAiLDjdTEY9Q8+C
Kt8tuX04hlEv5jfCtY6zPiFSsS42MEM0twa2MXiUxoBn2HHYln56EiJ/oI8rVijYNSm4AbzZL7HN
pz4fS816oUQm6D56rspxtrW1YzZNdsvM7ZZ9RUn1WSvKeYJF5IYdfUZaJVMiIflOl2DYHzByNuuL
crL8fBQNtcp1DIear3U11usgGSSiYNBEUvyLEmGNw9JH+lCQ8YzccMTzNs4wSfNG7wVDjUnEBWjw
4S0kFbRHCP8aply12MNaWKSi7X/XFJMW1V2yzfT4lIVQ23xcNgF4MZVb2MtHBylCrufa2hKJ9MGB
2RiOYaE1EZ9s8mCS7tsYLnakrvxwn9oX0ZMM5OhKbpVNBX6yRRaPgtjkENiVwRIXvVzKeuMBAMLQ
PVvhzVgMGYtSIie5kg4pWepL6BwRZ9js9BhivNQ6ikaVNvuk+86cszWwRrTAKoNrHvSV7XSmiRPo
qp3gr6XfmnXypJD4xMr+jvc18EOaN4h8DZ4qY+325Q66466zItw44+/BvZAjGjHXKhG3z+mKiWo/
drQ+9iFLTy7GSljn7Wf/okIg//h0j+S08TIdfz6dDEXM0yVuI4QqSSwADSJbpaO8Bj/GFKKt5LC1
KrPDdAembkbzNYYdb5FdQEcwAMIwgR+8MK35vHRIhAuCSG5qAQ+KSMPQ/Floed16hFonUptncXBL
5nFMZxfyWYrmmmBphdM49YIqSYJbbG71mhygQ3kaJJSpyXsgoVHuwp/zpnvhHGWFmMJmcIyI+h2y
2++bvu/xKiythRnEhTFq8lKjjpSIj7UoHi35wG1hbUEkE4Un05pG6Tey6HzMdiF2GlTD6gfkUKcl
pbHVxnajq/ZEJEYNkNVDItMExIsl1UZTGxajPiuzclK3gnZoQxtrWvkyhciGMkXIwttP2wtea0Ex
oWawQnNfSRBb9PIxYubaU7xtigtl
`protect end_protected

