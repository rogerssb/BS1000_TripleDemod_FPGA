`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hNWJoYUKCMS3NKBPDEqpUN3/tM5SHTzbnFf0cXlS9O8wG5bapAVhnYo7WCbi5bZGepFHKmhoartg
GTGuMOCv0g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o/7RDO4wbWYzMH7PuJvAeLWF4d2YldLw4LiwgRv2KwngM+dtzgPoDX6Xlc7+tNZk7wN5pm9HVSJU
e1Z5WHJKuMWIWDThlSkp7Wyzj8nsoprneMVnZYb/RuPiMnC4wphkU5WYbqi0EXs8zElrQiz+n4AW
bAJcAfLBkGs9PdsanqQ=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mH5ZLcJWPKlcP63Kztre2q+RcW6YrCSHi7ZKOAxBNtcD9c/y+BEUrzt+9ECzaV8J0LEv5w1RLRrn
/ZCtyu0HnM63iFGpCpDLPxjPgQ29f959Ju9/ISOpc9fReaL9c8zNHrQxPwX1fw6dUq78YDc6M7XN
sMc7qNW6RQ/BOCAdaGlOieEXIwAO/2Sax6zccyCbfXiXC4Xm6dWIRazbF5OyPRd2o2c/Gk7xPiBM
SJnvVh5RFDBFthXnT6jR1LmTQhTIYA/ozDqjsI2ZNz0XLDKPMjvsYEXcBz2/fW+B1jn4ETTeBiaE
2cLUC8Blxwb2noQVT2naHav1YCnWxrQv5Jc3VQ==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k7qEpRV7lVsvRo45xpEsAw27hSHrKfLOebKwKQnVNusN1g88wfmd4eyitfZX8dVjb3vd4o49h/PF
RRmgH9roiY8MPeV+zsFuiy2PeQ795sIAgaDBljM4Gcewzl7MaBmLgd0c/5VATTmq1ufnObHs88kC
mb8f8+4Fd5tDCb6XCVc=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V0mxbyBT0xDddcX5XrI6T41qozITpFwgpZ3WqxRYSaEDZum2cGWMlqvYBeYiOts0Xsneo3+ATPEm
c3litnzywSdTeVoSWAt1ppn217g/wkAlZUzIAEiNGf9zxOpX7Gzp66vr/wRdBmyFruFS6+Vifpo2
WfnferF+WCG9nEsn1R34C9H81goFYOq2gRUYrpwgr+GfBZL8rh2zFLS8c2l0isEfciKctmmIn0Zv
BJOtitBfQyusNZmr2oQGDD9lCXnv0OVTvVQW7oP6+4qQADzHgtuz6c+PyBeY0x+jjI3FqtL9vhyo
0Ez/J4gMreBvZ2WbKSFuRq7XYLc4QZWkI+mauA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16896)
`protect data_block
riRx+I8DqrZY3BtxICLWXkjWiCEfp4q3UB+8Cqw0DtBKvkU0QSmN6L4EsGqHfbSSPx50B4ZBbnII
h+DSZS3o7dx4/62GeMDlzxeZQFQBW8fRQwnB9Mb7EZ/YxOjb0JBfpeHOddnkS4AkhdgTNbhrZD4I
6D0MrcDozlEvebfiwJ+Lx7X7xYjMMS8+oUZm7lEIxW7ql0pJQ99lCJfQTnG8cf+RAIf5bxSbdwn6
lJdoJrdkB5tr5WDxXfGmio9Ayuq1gPlivKbKvXuT29ERfNqAkmfMi2SHMZZrordVsQ4Bs/oEt8yj
B3lAH0b8kGQqtUN64kd9I2Fn979Xe4f/FAFHyVjudbTOTVGX8NKfc7lQsiHWMxAnUqnMUd2WGD6s
zmL+0EDjzIy2mz2A5q757hBgXmD0z7i1vAvPOPNjNN+ythgnEuneGYfpPthQeIva2MwgdFJ4Uyvg
kQZ56TDGuhDaHKEX/9RZSoMtrDmhBE7ESB+4WTFMGQXyXJEd3fF/6hF7gIBH2iWiwec27f2BBmJF
SZKwUYpitpi6I4X87onUlDF9I9J0/MCQeJ+qud7oQzi4juM1cqxYqbvlL3Bvi/FOWvftdk+kvli9
JZgF4yrF6tGjdgR6Asw0THF8Zz+IkrnJUFH/dFEivETPnjGEtpzlogZmcW7R5MAgJYmmRPgEUg7k
cwJzwd/4cwJI8tU+JERRDjI8u5/aZbe3HnN0bvTG3LD1l/dD22zMB46Pvl994BuqJZBQVO0sYvx2
xEOlmi2QSmjrJhgoaRZQ9siZ+Z8lNHA/iuk9JidwT1Ms96CsAZ1ydihNZuF7png3+GxA7760Rv4P
sboEGj2W4kiZaL2MNYyMdNX4joBwQI6hQQvrIUjftIFcY6FLp1i/z0SsuILrRIJeFxfKdxfQJMAI
OGMvmDhAiHQF5jrE56VMtazCakMzlwQ1lajIVN22DO8UG/niH4Kc804kcyGx7SzR8KU+QIU+DxYN
qnfihyYUBaRp27AbCiRzAyAimX3QCJv9dwruO+hqWtAykbz4NtSKLsHGgmNznxe6NzZw4ATPa0v+
qsWA6SznD+aH/0Qbv1YGhC0nm/nxvV0U3Ag1HcV0lRyE6pe1tGr/xKdmogLi3Tarbn6rwM1nxNPw
W1gBBkgmcaGUqkSkEFgYE0KSxK8zoxsNP+nbTzbDt/+1J+b/0xAcbkXnQm7Ep2QhKwCTwbEeaU30
q9VkCD/P/5Hgwt9Jkbu7mn/25nKxQBorvFV1zOF/bip0ST3A59NiZ1X6sGUOGEESBW+36pFHgVLO
fWsWCzSH4tfffMbZ8RTyeeCY/HqlGrawbPaUB86KoGix2fsYj6x5vAvZU+lKapX+1tNrRev53oOB
/QUpoRgqc5uC6Ol0wDwV1jJzJb4MCY3JZ0vVHFEVpODVFd9aHmivjjgpK9W3+iJwZl7RkNrlOPFW
lThm1frVLzup9VlUhEBKxZb7Z3JYd3xLIinLbZjx+xYwdP8RIa4J7P2fotsWjqjj7li8oBcHkHPi
cwgP4wSaS6o0fGkdcHrEwtnxScnyRxoVlHTXbKnT+FKKY0k+R0samQyIR2bVk6Aqv76cGMCAe5Tk
LAPuoo6qn5MO0UZMjc1r2EL/ziVu9qZHhRbLohYplOReQAoGWej26D07X8nDUn8G+n+bKipSGH/Z
4E3RnH1xKVCBlmXE06/HJT+qFy73PqUfLAxVyBrPUh6cKfe0rVwCgaOOqiLS1UvkMSNtvcvBrnvi
jOKiqVSJ1lp3cShy8vmvv3VtVX2fOyzgFfE15e7lbIuRjujnk8WPH56D7oFPyK+KkLJ/d/PDkmp0
4rr9UIoWn0nKYHnwYP4gKs6DqP68ZiDM5Wyt2JBXlCXDW6nhZ3dO2775tKoycSsbfHuP0ye+Lypx
jCx06BZr9PGmqYrKbgyvN2BGV53LaFwZ+E4kqqNdil7A8cX5fo7uSjSyW5Pz9zE63ojSyVOfxgW9
vB6aSmIyEHK9vBFHMA4G0cT6c/9TTBu95m4xcWSl2hrMD69ncUDJtNey+ZB1uRPKazEsewWBbZD/
EmSYXxl0cIl5UMokKRZTrCY76km5HH0Wz0P/vgEEvJB9SwfvcSkroXCVy9dL1pZ2W8eZoOW6jJi+
hRSMCwLiya1qMs430decxhLU/vaGuC+XUl6QcVqbgAGF4RzvaP5vrXkLxFkiojmUZ3yokTLNyPt/
75nVM9y4e2JkzHgna/Z3K5ezjCS3cDaH1bcTmcgpEHSOE1G82XdxWnWE+rSIem1nNNGHno7Ws946
dZT9LMrcMG5mQhnOrJjsNa9Axi9hgWIPiSdKrgZn0S1hevozuDmmk8QW4ox3/re9U/OSLQB7UtR5
YGspGuTbwlKveNqwxG6RXOnimSFPSlJu4TCt7y9kN7XDYX45BSdiLDCa/iMnlV6JU70+Lnd1Pqgs
EW0TjOwNsVMmB+GSYF3JIObtYKNwBPHSCeHXRousiI8cLFlaDz6L76uIWEp4NX20v/lXogJdU0Z9
GhHKO89///m9nn0DGR9cLd2w0U4v1/TVSu+Oh7oujdbonLdAOoHErxrsLbzlSjZn88Ql0zlDV1PH
peT6YAWYOZdqkpp0kjsoS/tcfpRAKZ0yCgmMDZL6zDZ2YRR8cSblJ1qEw5Lums+llF4US64LKyX/
L5W6YVZL9dMylP/Djd6kV+Za6ZvlmWBqu7nOVllSVR9v3+z4p0fPpWyY3E/eIgRNL36BnfgHrZ00
Zi7lYEVowYdWHZxO/VN1T6ifZAu6JaU/jrjXZaOVC31ox+wFqLhpt8tSMXjgzt/Oc0b6KspePCRi
oMlvjFyRlCRlCQksE2xGcN0I5SZOislg/Q7iy6lsY0MT9IWIgeOOY50Ht/T592nBzvM6GOaBfHFd
FVx/n/tqcReNiFigAOo0zkmX2Z4Ot6vxhZ63FZNhqvdL6lJ3g2LwTt7aZ3/qLZVCI062wC+aFw/P
4+0MTPG+GgO6U/Ws8HuxP5Gyzz/GbrFHw75clin7wAF0/+lT1GUX4R7YyDiifwd1tJzkC9xIjgyF
fSwsS9fvzYg4qXNg3Kc4S2cziq6DzWo3l7YrzNCAC6Kw5OdhPrIwsEExAwgwQnncARVt00DboGJI
Ot2/cZpZVVV4vLn9Tql7rmXVUl5X9xzEBOOPljhdyarF5D4A/dy6r3m3NpBAaNBnwKPl2sixRInN
xcbw+50XfBGikbiPdJqtWavExnUwDSVvCLN27Er28D7bxCpjg6xwMtVm9dhR9YGI/E+qays8fh11
6Tugr3xrG3ySavKBFcT0ynlMJEfJ21gJ0Qw+21CJ4luIwgLek+efp8xsTEcS684rA21VnxWpqQd4
M7G22QE3iqH34c5b0vp24LI226RPszFVcXgfQj66Nm3fIliEmq5/lXXSbg4YY/fqevC2asFFrWcs
UCjIqBt3w5YlCE/CJlZ/c1DHYMvm8SYbpYPHdXjQ67LxxWk6/mpXFLHqSNV4B4gmDovP3OUZZbYq
lZhNhK8Ln6JGPEVj66yi02xn0GSNT3PmRm1Nn4KtDXOkJJ/+9iqIygeqwlJJhiaOTc9+oAjsennV
buFmnnI5zPSf5OSvjJOlpRF7TECZE9s6heBbu7Asci9iQOJVObLS/7tS2ZNnGW5B4n0Tn8prVesC
lIVknIq9axC71KhkQM1v09ucvyFoQMSwO5oJsk8TCn1/4AJqiHDQway80iuVghlDv8cVCHZ2rJIS
lZaI/CW6gXuPT6uC+Dk091aT2JkDHlq58pCvdCbp6ykL06yxQT4VsJGZljK3ZgBuxLOCcPJKA1Nn
8d3RKwJm0KBMCZmZei9nXuDccRo1lmH/scC3j8uqNj9Iqe6fySooibTbttbB7kfoBCIKqVJ8bEQl
BmwKnRkTSEmi25ZXkHQiEiUhO7nrjRhy6LCyOL6IKCZ/Ygmj1nfO4O45qoAHhvvEPH5XNLB5VlSa
156fYU7KlfrtmnMgngouIMVwvxOoZErKiI0wwi7CQ4edt6+7uCdl/HSZh5oYF5p2gjSpYzOWC5qf
Yg8t5RVbe0/LauPsq56jw5zhEjtonWW8/Km2g+gI2CTQrdmWAtHKeJnpw4eBnPD4QkfCizSQ3zAC
aU5Ws+xJlEDVVp9SL+gyuFn6b390ZpoHyTRpi2d7qwWt+99XwZvlFLYZSe+g22PJcRC7tZ609iJy
eoZmNupydUnd5G25nUPAuj9hxgbMTEGid3JSlSfR42b+lgcdefm6/Pz4X3MeAmW1y/KcaQsBpEN3
+CL1tvXFzFRwJ1lBBMx6mZxMHJ3R40Y9ZrCUWDKy3T8KEAfs9mdnB6S5D2UY2uwgeGwJjxlfZHwl
zu/IBDBw/e1WQYm+JHH8TeXdPIcnpkt1m9R2JDHvxvaPbtM7aB/opmLy0sYebnIc54foaga7Iv64
7AbYjm9OsXFGI9B4QmaWR2Wf/FzH19/8wY+bc1lLgnfXQsfcXPS8UnaQIsPrUo37L4BtNAgShajp
RXh0JRH6SF92CKABTsI8ADtReWzlGozMjqT33ERNkifMqKQ9FGHXKoa307W+rxGMf+dFpbAhy2eV
vEuUxuzrlnbnsknMzQh6QiuWdWKwbSbsjNq77z0LNsv41y17C6CC37SduANzur9IFmG1S6dyOaYX
kCP38D5gsurojeHBizVY+2nLSNYMNndPJIlgIxXPEEDQ1fg7UWzRlxJuxqRVPYhh/bk3p54FyJpL
uHdV7HR1MpBryRuG9qVUwrEMpm2Wt5uDGvi6qeU8fnlV6feoQsEa2bhCvu+0kM36G0kkoF+Nohtf
MW22rAonsd/eC9/wPmDz0n5XC4va1GSm0+uzcFpVQtfMqD0jS/1dGO78iJiWytpZp4t5llmelqug
RbW6m9OSRvnUzqfDaQJOoKgMgKUnBuYFZqVzan4TeiygSThnnJ3EaxwmL1u0CPxiM67W6Oc/CY43
Lqmtpe0uVv8RxxERiRjG+sfb5GGETuxj9GxUu2RCE6SdyIbCNLFsmvc1jtl+2u0frmP5ui8gje9q
v2qUm4vKlHmUCaP8Cq+xcae9U5sTgqMJIYehorBmjPrJMI+HRyTVQzm5vP/44IT7TsXh0fY+bgzO
tSKiNq1Z0KyQzUdhbss94nwlgt0kdgWxzNLrN07vpMurO2q7c6+2dPPDkPxitHkMwzTz8fa8l4CP
6vmcIgCvVJKJsN/bzzUAsQUw/Ax2Ui7udMFSO+gmHpB4Dn1uR0bm61luxRL7iinaZTEL4TzoKpZA
i94dkWIKTco013CbjAXqcl7VtntprycIzohMjq06BJWf6XdJs6Y3lqnYKoB3D2h7U1LBzVVEFv+Y
1KL50wCP6NvG0dOVmgmuwDM8wE6Ppvinom04SEjRMZJLw3iB8KME46cGi6hP1V8r1/t+YC9PfXB2
3qneRwlQYWgLHQKAGjD5wvdsK0tggndiM/jkm4QowXp78Don8dNLUOI7OBCFKzktefXOSrji8R/M
kpCn1wP1IxPZSl2FOgi5opXdTRFg/Dy532ffe/rUEyxLbq9MFFOalEri68rpDh1z0Ddk7uyfRhNv
Rd4cQ1Yf0Wgx3jJEAijnVIvprgAaw1RDt/iqn7LqxucdXwpigIpmFyvpzaOaCB0ITOCFX65nEXdG
qgMNNouFSUPQE+Qmn+9Q3GAHxSdKWAWsZ/WsvBdITBDAmjn4YIY/y4AeVKdLUfrKQ2d65pCe4zpz
3dbXym6C7bBS1px9OTyf5RsiHH+32UJMg5657covDalilmQjz7sd8uo0wwvj8kRqLyOebtBYvWND
hpkeWvgjJSHO/5fuyBNEauiMGzZE3VtRj1wTEXT2X47mmA3c0CMMeADlqYu5ZjiuRRl7R9vOdfya
dAGglIyXoPhlxmCGdxafUNB1OpAgIj1/1mF2Vb7RXXrq5WW8IZOjQaAwqGjFLEDdF6ZpeMwY4R24
i1zMuLj65dfg0Psr+F1hztkIQl96wa0seLODDv27YPTHalmPcSXxpwo0HwnKFVty6DTehy+nanGx
wjiKRlYkF2Zpy3Tfb9rpDLD+P7P82hzHkrgd/CnXfHxCCnUJYr5aE4urgRuh5Z6ie3NieTKbwaID
TlmlBMXjcpahtFedBb/6QK6/EeUkzRSr1JCl7Oq0ApLhGmeNwDBl/Jk1uq9dPt9TRTUUcYt/Mee2
kyOsu2Mo00jQo/ZrUUnWLPqyLFbUs0JFFBHUeeWN0hsCq+cfvM9aWYZ/E/jp4Dsac9TsYxIuOxbF
XWYL0Uf/SMN9VDanjXPyW5wWSkEaiWMXLQ8VxnyPmVQGGMDDzIIP9ODZ9jQhUgXzpA4RbSWGH93M
+xqX4i6ObX2AllxNnY6GauxSGWiocrDflRZplKvYArK94OWfSi2pD984AK7JisRa1K1TZs8+GFyl
LOwAQuhbBgqzM0ddTAH5FykExeTEPdCKYe5n97EryFLOTpd4URH3jUZysKTMu/2z4awKCXVoZuk+
bBVS2uGHFHjVr0RY7lXrTfMWbmRvJbYcuoDD6+IbDTLe9A1+IC/UPYIkL57IpYP9pTQqF79EYYXB
SwRjw4v/8qbG/j1gddB74hanKs52bIk8XNNLi9uowc11XnJthYa12QRVCFI9JikNfXu4UFTZ/Gmp
M4EwFuNQv9Pafg1HfaaUp/kKAFxNI+mGt+AxnGC0ca6YSQn++agPB69VH92tmZ9yhzxFVsY97mxC
mGwTtkfLiLU7nxQXf5H0hX5Zt848RNLYpT+4tNndWx8jTxwOfWWisZc0s/V9yGgAn/hebCYdjA4p
VI4cTOuRDG8H/OrLXrx5E8SxWWuCIEFR8ulcuSDtwDSxOwur9EBabz94Ax4+fuUJtF7zNugA6Pxf
W/DJ2vc07R5dYlTvBYgP7wIl8HESRUnKFpXmCXvtZHIoVv2Ki/8TlvOSyBK2kwUohHPbuLlrNXyg
9SS2MkIFoax+26BWeB2CILq2ML1Q9+N85aa/1abgIvP287OHNkStcoCaRLoFPE+LUjbH5tuu98TF
Mt2T8Xod9fcvAU4c49xh2kIbHWr9LyjEh35qiVDJwl+yusz+yUsjS70g+wA3j2wOzQz9YKbe90cw
YUMQextZ0l6L4JncE0JIovtg5x3vtk0KhqoXWWjwL2Idj5/EVMC4llwhiNIYpFMOW6KvOaFmNJsM
d6blG/WEbkjaucfPTSdDnaPn9foML4/BZPtOTkVe5QtuwnXekdUpZXcN9mGqo+KA0kDmloPnBEal
7iAXoGh8AVw4TaJUrUjVOz4PxkeDH0Of/UIw+Dh1d4xf0TdOua/xILjewUs9z+YCFwOJs3K5Vnm9
crJFihEzlVNWYdQZ1T/282ouvJq2XeHq+kdlFwMz3427jYELil8CW22qKOX0S5YnWIenwe+hF4xn
ffTxxcz0s+J5OeNDHxFIYGvbtNc+DdO3AEQNQ+29a0npG9YmTRw3+qb7SWvt/G14ZP7FlmSpQW6J
VBQIOZrJS6BFzhTlim1vEc+cQZXnyt8iSE5PPPTfwOBgIOcuSZSJHWYRds8QImxOuxzsTVsif7tX
skTukDLVoA6OVr4NuI6JHJhhtVmHCIgyE3Ap03RpNeHmBF8tnR22Lbky5/LcMD4zvg58uXtvQ9lC
N6EdIuB3SnPaM2la5jVfProbR9wj8v2I53enkFDDxvgMVV9d43xpRV2UvRbKC6MIuWcrvmNlEr7c
olR3zgwK1Tz+9azdo+wmaqi1++221MPSupll11BuwfrTFdKeqRwCduMRFk0bZgyWfC9wQj1IlkLU
2BiaoqJ6CbKv3lPia3iGZ9LdOd6EbSydhYZ7ZtNN0Bwc9qqgIiIRpFp8My4JrD2Q8lL3ggsMgf2t
i42F85tmTy9t+wioFh/R9Imjmoutm8YS1v+UsYl6DFz1U+NijGoKFQ8FBITtVlZ8/Af2MPDOSQ1N
fByVAQN5BoPoDZ36ugo8PgYHpgA91GZ9dyOO/aG8D6RvEk0GNNQZdUxA4gnu5zGoZ9KysKeg6zMl
b/FS6jH2TeKZbr5p0f4TwtIJMk3IL+amdBR06k/tDVHr9LPKFbStmQ1/DBbosM4nZICXE53nxFVq
KGcAQk07IAQyB4cr30LvxWchJUkTPAqTM1K1NQsJVKlZ8IUDr6ptWh372IfTF6RiSC4b4rqfbGoI
jrT2i8MQa7F13iXc6qoqEaZwfT+cWISWbGQcKwcNaBsdQu+Jx6orC0pnPWJin7mUVO7Pt9GTafwd
kfPf7t4Q87x5v8slxPkfR7k8TH8iFQ2nVvr2h59lf+tLhKSTdWoDZMo7c4EyJqOQzNVo21+QcbDr
TgS97ifdpOCRFbSJowMbBP/Sl/gtypTVrI1GG6IsXxUEryIV0KOS/VzKMx1BMMC+yS8EoY+EEi8U
msT8E1bVXyT5KZVCtSThEZTJEpbElULexlOYsU2x1o79KB5LrDtqSXZjfzqAQDr+CmOX6YsSXw5p
nisfDdJhsL5KftUIpuF3cB2xLlJSNXZchfpeF330O3Ywy/5HRlrpzXzxJk8g34vACw+SG7IfNSav
3JIPwoXxvXacv6dxk7ae5+h/FQxc28hUIIajGmUmBw9LP2pChqHEz4CwtXmD/UjpzmZRATLu1oEM
TZ3DbVvoSECyEujSFK8irKryZ3nxnvKjk20yVzLA3RXzuxJRK4bRj6D9xlPGiMWpTpb6FeLcggT5
gawhomlmKF9cjiMgIjT3oDFX5aHZnoE3lpHACtxHQt400UKC9Isvrsuk08PkEwcYXkwzTW1ib4yr
+M4Zqas776jlYnuUh+wbwozePB7YQEo1CwDMFSy/ihDb1XOjsuQ10DIqkWdSC/7KNfCDov4gjuCk
Ga3igoXyIbfhQYhsh/CrTkax1kTTmcCwKijsGD6R1WorGWpQbe6G994T40NZKIat2RSR16+Pj7vT
jrr2UctN7JYmpj3fAaSHFHxyGoXVQmDDA7UMZJS/MDGaErRNaSpo60JhjnjX+ZfGmLVlHlUZbZMB
u3396CBXEkVqzRYo1KH+IwG1Wae9h/f1wjMkxKdLD1U+LbGDvPp6yZ/8cp6sX/xIMpbGSVBEr1Lw
87W1TLJH9iYHLDAlgYU9OW1fSlZEyyPxALAdfpaU27SF3iuAxZKXLDZqfRd6aqDaMgVIroptUiqK
+PtwdJ+h96xS1DPc0h9VPIfbZ8H/O5GdiTbzE8gO0WbJuoZlZMSHGrC5P9lGO36nyg6HLohEokqt
/NIs9x950UMUDRa8r+82gFcTVgpQ+c9PRSD3mvhwMHq5YjckBe4Bm0Yn+VdSbr2dkoznr6MjnPxg
hQcil5M13MY8P/ZTxA8pIUy1plMvwhNG+1qteI9sgtZCPKwlG7SEl1IJos30BuLfqrNUKYL0LgQ5
y0jSnOJyQvUoOE369TNFg/nH7R2TsuOi7rSOZrZfvPz+XwpSWIQJgL7z7ziS37RKR+z3/Vxug7cZ
TiWp5mekAsE2X0AUFxgfiXou0mpX21/zLKUk4Xth5MMbGQksHpJF2zKgxO/+e9AU2oHvU3Yo/J9+
WeQTcQxPxHdsVqPwy6Ya0VOTqRGU7KKFSyJuDmuyUj4W+Ox6w0s1hO5SDhvOhQ0KTC6q0jH96lN9
f4O2fF598CDTd77MPMl7d+tcktCNTsj/pKsBNaDncG58x7gV74JYX5UqKlmr/66erYt0vkdrteCZ
dEBzuq75FPZnfSGn5fb/A5ICGpFCaPwCjhi31wiPt3Ur1xrA8Q7m1kPnl4AtUYZ3ZduUJVUU9Ohi
Hm06fHyLDd37lrLdTLfeGP1SmWPZwIb5PiYuX/QvIq2OM6PfHMnfLpWvCzuVUtVW/DdXIP7VHxFx
0JZUUgzTHEfsZ49ote2BJFxVQRhRF2jkQt4rc+x7XzXjgPqLElkgborbQ4ZJX++87KJHj7EEhHyT
j4a01I11eQgYZRm8/AwT1biJgxucDraI+CakE8xfBV4YRnsGu/cTcnFqX41fUQLIF2V/N6k+Hgka
Y2AwBg81bH8rgomg0DQWrKhhM4O8cR9Wavmn6bleUS5c58AMGAM6Ef2+NTVPXub46cgCzhXzVk3a
P5uaCjGFJEnJaU83fwgLrM6lrpN+6NzfxtL5zIrhgQmt7MuPHX84F0DtJOFQLXvEyaNSqdZqHvCa
W/qF0GZn7N2DcHpG/yohPmKOGs4tN8Rs9feQEHhfXCyQty75s2rAgZSbJWI/5WaG5HkpL5RGvnRT
HmIRdfB9ltQ96Lj/UlsjlKfqqygXrQw0xVXvyMlPJpuX3T7i25jBPU5D2DbBNhPs0AjUn8JaGn9b
E5B79b0jetgf6xVNuQR2ctuQb7RblMMmFrlp3uYqx5w/YvCXMECUGIZnXTG6f+1L3m7Xhj0jrbTy
Q9o6+YyG/6U+uT+8m2sE3jmVbyu/a/sGwOd5L7xfbH2jxPAydcWwd7RZi7fenvQjT0PHFydj3V8+
p6BQ9gBohMWKChrjaL7DxHbc1JWr9y4ittgNnaw4vX5ImHKfdcX4++DG2HY/zM33XEdDJNY+IuqB
uSz2OTp0yo7IfB4Cs+SMJLA9NrmGcDS4ds57nVrYBdH5FdmBM/HvIGEP9q/YhxEL/BEL5UZPQ/aK
iwim/gX9luruI3YXlZH6qqQ+s06RtVSnwNqcHtgKrJWJb4c1cCYcZQqgAskPjudJGKyVGSJacfkQ
v9/fmh6bTEwI/IB1eams095AmFtjCVjbCqwC+g7Y3XEIZD0KI+/zNfWuexBqRkUz4nU5f52pZ6nz
0VWAY/7jHPTDtZyo+Lr+GaFzDxV5uuIn9rz/Bd53pVEo88edn/m7Ij4L6FXkpV1JbhuX7woCOXW/
loG2AHqJc3d7rBjjznuG94WpKN8tKs/xCovH4A8m4eWvx7UhZs1XGFgckD9oVi6AV76W/X6RRFNS
CFG8bdrvPW1ELm0cYGqv5t3Y7dDvDNckUHpvdirhT9VJkxSJEGwyEFy0q+zGSWZqgyx5Bw1/B6mc
tn8fIAPneXbx13cWYnF0ywFu6IIMIfFs0Fu1v/aHzGMHLK58ICoWDdNpiCdvGjwOUqETzlVUWfdX
b13V2lPGCw///NYncRX9SNFJj9pd8eVeOLGD/Rm/Jwu6fnKT7DNr7rgvgBGuoHntGzjcPPIo2CpP
x5p18Hb+p7rNt76Ij3kS1dO0cJB1GVMCb/eEonMmioqvHFR02yYX3RmeVdgcaUV04bsE/4V11daO
NrjgUi6QQRSx8viv28n1uBhcfVuKIPTKS4mXtHm7GTMj8CfHvrxyviscafbSrha6ScaAh3da+15T
uBjMZB5WpqBmrQIK+RzndltAUHsHInQBgdnOeTVHWbI+FGdaYbhV2f4eOjdaKhy6fYj/9yuvDZ6Y
hPSBZaAmrKcmCEGmbwkSTbwLb5FC793SyNrDpYHz5hRHV39caT2jT2ZtRtws+G69j2zf5m+ry1ic
FC4iQHUBbA/+Cn6nb2Jkx4PaB5I+2jZ2lXpwZ7fCkDK3gaEzzZU/LV8w0HtDiKuA91X8n/fnblv0
NddwKatEPwPx3LjMSx5mjbUfOAVtFSuREX2uRUZR9l3t87P/sF0QDmteQIbpYrKiV2Z+5K9e9WxA
lqZy7ZmEh7q81mMoO5ZOQrl4unWwcVKy+4UuLDH4S7LFEiTuJ8qWOxjAwMaCrhrTevQsSGeMgHU2
bM2GmiFsX77jBbxBeJg5iwhdp8IVlxFOfRFjFedpIUe/fl00Nb1p0fcSx42RH2mzmsvQBlJV3AS4
gkV1iaF5vBFDfWKDNS78rb35gglaTQCT4g62pn2JmWLxzE/inE/MIg7DCWKIyxSbkn7cTRkON61q
ACghec96ceLENVnG+hkyOsfATqS3F1hfxWaicMWgVDUsLJ+HtLYAiA84zxCbEeEb15JGewE2hzL1
Yf9h76fhd1wLNcTP/fWdymo2eU1rU2h1+0yaMByy2p0CfGJMEYEroaBrGdl5Dthf2APUW11VhuAX
Qt4Jbc7LTii2g5ZA9N9FFTdaUYwa5nKjwW3EdRgeUfCVXXBKFLoq9QQvhuOlg74D7H73X76aMA9d
wkmmekq2dDfT6noiBt0GtS89eHU8gZU5kSR7YrBefviHHtpJcdpkUHbN+SRqo8W7UEWYXfSkThzT
a1W6Q0+0GAn7UoqazoNj4ymeY/fOQKYuY6ZK+vKSaojlDjUsBJJGJ2t0Numh305ZUrYOJhwot2Hs
knB2BBl9nRP8YcuFRzlrQQ0IcKnp4HHE/5AHpoYikWz+6HpMk2QPKxTIqiqTBavszHYI4lB0tcYj
HJpZu8byWLGgBfzynwHaa2f7NSOr5z5lOHWE0n81ikzUmMg7458snaYsG9HOzIdKEQcWY5jMFtAJ
PAGVD7iGS5K98pf2ws/BwUQWBmMgNa7uo+tp3mYQVEl+nJbLtDY8kfsH9Wc2G3aD+3zlXYijKQkg
4N3UZi6Nofi0RJJ9TVIJtYWcTobgKGFrL3m/rWH/3Q28m3KF5c+mqb7gKxIPlEvb58aRBlWVQduu
TEB5oSpdAjuujDybbkVWv1M4zN+YuiVhZHGzX9a7eWF7TR0cs5uDIPnhmPqe1LWD+DKs075e5mt3
tbX5BQup/T7KaVDvzF9R5ZYdLhIIHBGH5zXu3+gaVFOuvOqNmv+MdsiZj4KkSQrft8f2eRAUYpag
lOO8Br8KuqhUI8zXWkk5sgDzV/sbhS54UnfoKHTeOMHW2OVprfaljvEuMU8a9zMHijOQ9+Tq/PrL
gNXDIr2EpusRqwg0xuX+yS7t+r86vR7DUP8hYkCkV6wIqA6yNCRTB5IyWDzcZYL+FZrWncbgov2y
JMUqy79qq7qIdPyAAbQpyPw8LZuBsvInn/Ewn1yrcHU38MaGbZHutunPqGuEtsg3S9W+xjiV9ZsP
bJoPh5BO4xJnJW9ZH3WP7CWbxhu3E2ZrkhycvZKOPlQZA9bA1epqQ46SPvVS3AsRksZ6h15IH3CV
/mFOJxC/Qr2IcwChbe5MzB7hpBpIRqMvKpSt9C4hcbTVUynsIhcUihx5tFayllgFCgXJVvRjEKI4
x+faBctU5CWliU1KH6WjgUwL4t1fkJdUkMWcBE1TxUU3P1JFSy3kRaE1iLoz0OPIZsHxoiHRYRIK
hwHcDVMSw+lARlrWRe3tvKRvvARvS48zh/TwdNR2vhbiXjvmlrEWk+LeLNWqgnAB/X2w+t11Ddeb
5vrfqBA6tix49wn6nPvsN+8I/KtGTR/FEmxwPawIg+qF5O4BbapL6Iem2NHqg8DKXXYunXV0WkWB
O4IuNtGc0t28Jc+Qo7HoOgNv0h4VFOgarmPxQZxEuCRyArRBdXb6AzyNBkUX5bhw31J77WBE01EH
kE9fRvHHTT9VhPsQIUJd1MsTYrhyrQmiogDIfRzEqZ0lOcvg2G1Rui3R0Vojj1teLy2z73T168sJ
1hMuTRuBVoh4Beu4Dn5IBGA7S4ehqsvYAwlQ6ACpSP4pRj6eUf7jGV9lREDsfrDvJGuHMo8JW3PT
NAPIc0hUffXaWE8HwQaYQsTz4lX91gfGoGHPcBWCDwOLT0lgUQH/aLOK5eD9JWeMquYfBH7TUFhW
B8VktefDTTtHKIqX1iqmuB/7OYUkyr9LInb+B4QGMxKjThlO1GkkRVGitQKvnDkoRpxVk7QN80Zn
UbLxuaU+xa7Y8ifzS2ohSVVLnRg7x815rToyvc5kywbtg2nuFJtVdzb/1dmg2jUDQVrROhwIZ9dA
hdeC7mz7A59A+KslUg4dFA/3g9R8kBkS9QyqBOyg2xLtKGPixSmkteBYyEEoUcYdpukB1iTpkved
jGxSVwhHUwqxB5Qlcju1QYkKYLMbok4fhe6ChNP3USQdnx/NkI8dW51YGeBauNCjPwM4P77hL+CN
h/+/jEBC5taJIquZcD4kXMYbL8L6YJfvAwhfCLhTsDhw7+AgXk+3B6tbfnKaRGh/5LsrNYVKqJyt
m6U8So7IxRljHZUcKFAtmxLacyO2HOe/Hr4Mretp0cnA+hi9iUy5bZ7TbP6Dk2UisiuCfx+pdDgP
AmNlweL/nBg60p1tVnzG8IF/2GRDGwb7GDNfAfb//AYxlfuYM/ZZfXYa+dPHudaTtEFgdid/q4z2
jC0PmhrRBM5WUFX4u5NM6ZEfvTXAl4q/Mc2/Yzwz2jQx0FGTw1R0cbQbhp1xwqp5YAruDl3s8qGv
tIJEkp756w3RgRfWVdLz4V7c/kwmECHdceuvpgdF1aG2TB2rXChVZ4Zyu4I6I4Dmuc8S7wbVo4im
O/WWr3Gtd/GYbLX6zPcvZDXSr2t/mEazsCPvqoDBxubWNwIgzU1lcjufc8SHTmNNscSshdnznIZ8
Urnb+RTCUm4H7gJotWyHrqtVrpjgayOWwSBCtiKrJQM9wtNdPUTuIopLQey/Ct2ejR6ByRlRZa4P
cw/7GA05mSqpXRJd4zWYByOPeMkhNnfz2CkRfecsTwjXd/wEnAPgDY1nMDcNzBb0D2nb2VrxiOzv
NfyuUeKQkuYhvaGZY+/z1oEzhzVwceSKNTj4bSQBkyQhZOMoYy/T+qHlCcW75jHLBeq3VNH44UGX
zbzNINLETN9/wV3wmCv1ctXlYhEqtoOn0Gtwbm/BeCqfz+9WNdPQN8/xTpnrNsDACirfHRKSK6DU
NrpHvfMIR75CJgF35CyA+vthEM9w37HX01Cy9IOoAr4aaOePnTwfGkj9NBoTkxs4MdGOYEYydN56
9s6xrzlZ5aMNJMnSxMPJrtRPC6jTKQqL+Llqb3gDjeen+N7CY8LOKw9if0K/YmP7ToK7c9h6P2Uz
iD2iwZmHHub9EsZOTJTuEMafpvguiUvnlq54t4wuSUl0hpEaRqmKszonAs+t80Ly3Gu27IHajl3u
1EQnmaE/x2/big21R61ynKpGFgNi8/jy7oBCYZSq7BiADMWy268MxBdv+kDW8NmGo2octY/fzqvx
v9dAQzQjzS32PbHMn2X+NEMOGdTuyD9L8maH0LncBiCLXxmR5ErT6c7E/EUXpdQvKmKA2qnG1x8j
U/eBx9weTuqjGlGCk41Q4SzGI2UEFj3aVdb/nBL2O1scUjAciF/rPgw0ex3ga0kkfnyKnUT1RAU3
l7e4PJYBQ9QZyNuwTJoL5ttTa5rqS1ZV1WcPFaIDnCXkF6XiX7cPv1WF/AOCsxgxY26T61rY0Xxs
6Z+HgE4XyDAptUwMFZdjCv8XOKQ8FCQKTWKsSA4/zR7bMkepgYCZNsSFZamb/zfj27PGn0Dlpp8U
Wr2c86YTUDN67K9itsD9sNx9fNP5lylL57Gy2rN4SmABN/HUwg8wna8JmiIV5cSEhRwFWmNWtNH8
cXn10UBYeRjoItsXQWtN7vwlrdZQVkE3tCfhWxjXc9qaQm4IchMM/2VgHr0ja5OfXtISXlAqOXAC
pb5YEmdAyRTd8d0+Rt9+Xol0TzaEExT/FoscpPgt81TxvQCGRDZoMeJJ9xCyynXb14AzAvJ5wX9Z
uwuQtmeyvIDxwuI4pqHmnQRyjCOOtooa1H6enpAVe9ZzKq10Q3uG7faPO5t62engo/BRdJ9qvVGJ
StON3SimRL4rZLgTByPlo2iu9IHjsZKFm6BH+5Azj+xXXriQ6Qie6IiN16wP7QCtHSp9nwUtnDTB
k8nsB/8EC2iRtUYO48Bpv0He2xHs27zedhFzrtN40vtSXd/KwjufrPq5G79ugBzeZ+P0DwsymgmJ
nDS//sNohKUhUWpuOMywLcaPATb+akTKLSlFVFGFFT/2WvEY21CZM1QAYeTYeJ3AHqvnhgWY5E6n
z3R13ruEdmCqnSNLRR0Vgn+PdtE0fz2bMYvQRrIQgxQqC8ha20TEQ1TRgKdAy7WpH8/PtuElEXNO
R9KTLkDWPUSY9yOvc5zcVPZzafw2jFlGoa/KiXR36f4jNOf2loBVkMHyOoHfXCZ2NHEDmkTviDw4
m2uJsYm5+UDumTfwPjRVDJttniiHpZ9FGCD37KnbvqfjnhvLI0Htp7J0F1ZuHL2BBjaMS/KivizH
kB7z6jDSsQGOh6ACQ6/uH1szkbYCc0c/HErRVR9YzWV5aqp6aO2rl4rUUkQUoNO5wQgX44V99ujn
E1CKTa8AVIcqjabddY7YwbkvXFb1Zpdj7NHWZBxSYq6MIcoJiTMlDRLbUMeEz3R5CAaIqW3otNdi
Uv7n/u9pu4lKRfi+czdk9apgmzt1kRAT3O2OF7n/bt/V3xlTGnzSxWfYrLXK4+MiHb80fWcw+On9
v6vLbIayirjETijsk13ELDlSJL/IiyaH6q57jphyPOgh5qIxH/5WK7myldIyBlN5ZZWtpBBtdkUj
FYQBycS6EmrAxWy54+jAjc8LryllNf73ek4jyOycrth7R10kjXX69OHUlfnUX21n+y4NJ7woRT+p
qf8NGzzWUuyR5x7dDB5/pC8fXnwkDYZ/VkAF0FARp+xXzCeQpwlLW4IBnUWLUc0IMwV9Yqn5wfwn
4anIL2Ne9/8AmyhA0kVUPL4UP+pTpzMmL/GXlCjld2KUdngqBz+O58NKnH88w62fSzfkh4hxZhvC
DGkk2YziFucmy2rUVA1uHhsUVdCnAHD3Hzu93mzGGSFzVL8gKFAxnIYqgM9G6804AN56qFUkpkR5
frkwHTReM7Ni4LOa+XsLK4mkuaEUAEe+aw3yv67gfOWVmLt58OeWEDHmsBSK1NzbKeCVINh1jnZH
jqO/ZPYgqhFIlsskpRcLbZCPDTDHeBYk0Jg+IrPbHC6M5qFBRBG0yOyiLArGDiNbYJgBDsx2nzdA
mIIDAubQoEQ/YcoNLCtEjnGGfuMvKKoGpONTW4MyXCIHrS/IRtspM95kXxPwntVT+5mYpNpSrcdT
7PxN+XcODQhB5ZSBr+NWnFXI4lil7SkmXRT1kbl4CHuBMD5sIJUDcUyep2BxyNg95YF/fr9+KIJ5
7NV3XYO++beg+wZX+Wkfkb2vEPklYOsEKauXUb7IxEQYUIUg1reMFuJVzV1RF/MErE81/Psae/bB
K5NoDZxnPsnamu+qFXazsZ8sYlvJgyDL9f0JAZnoJte7nFlbJqLc3XhXcac3jAo1SfrgsQHvsPLC
JwWyIl/ITPoKcCz6Md+3VYeuwyLcTUZH35M5k00ifnlO2M2bi71F0QsAApHBz9NbptgIaCOdxnhI
VHhGbGPzujBbRwngsHpDb53v4WDJMbtKjbMPapeO4vFFU8OzU8xvbSG7YWcAs7gevBeoUb2TWUqd
tJ2jKfTaKaCShu1VK9K4D1bGY6sjy+Re6+TnwjZxvr41RqQZM1bLT5IoH1xWjp0iefIjCmDglFiB
t2rcIhKFTDVZr3T0TuvvuR6S3XgxPuDTA5mue7Qb8lGSlkON6RQE7xVcylAtBXsTUNrpda5TlTSe
5es2wm26bnQ3HLYRRaeLHGookuXR6Ysw+meKLJ/zl/7pv5YoSntctVprwlO9kb3HV7nBfKQRflu0
Sd8TpfGzDokt2S+6p+R4cNP31+kmAckbeZqWv2Z66LZUKVyHDmEBmuqSYr4lMzk2y/kwFMaNR3m4
GF/VB/ia1bUjhZlC5sFzbhfyefUELLni6D3xraY0Y4PzvqZ4fPT9xMMj9hUJD8C6tMwqyfAmctzx
XBpF6VGQkGQa5bN85itiCgTqi7c+T6I37hmDaWGj+K8hn/SIaqLr8G6s1ZDpopbOVSq70ZCieZf6
5Jt7CLsrxczV6xeCYPJmr5XPYn5vSvVI5H8F2fLhEe1otxyemBL1tRgDOKwW23KvtZnc5uSIf65o
A0923YMuoqoFxVdE+FeLiy1UxLpvv5TyRrfarpKg5RwlpmPyWL5R3MsgdF6TCo65ZAy6hE/rZ7PA
rWOx5CAHviF57jUA6JtEfKJ2+spQqSg2x6ZM0tCAdSXfelzy1hXoAK975A2ExUzQkebVwOmZjVoj
d52QlAj2jbu3wK86SdZ0Ud5RGmLPYINExW9unYi/Tmok3w7ob/IgIFl0NEgpCMOq+IQ00w4vr2MX
hMGMGjWwOZsL0P3uFn+Gbf/i4K8AqGBC8tUZF06y6kSRugqTuKDL540n4nx1yhE2SUix3RNp5Qr7
Er0T2WgTmJIuaQgcl4KGxR0BAOGOHftSU7KDXR64tub1zSZ2H6KxAp9ATk4FL7K7k2/x8iiN4e28
cb7T/+u1PCVi08Ud1QbEfJn//pgKFO/r8K8fm91gdh0RW7p2DiaYKEIBGD5GSM4PNlYWocQ+wuWy
QP5p0qvnlCnKE9KQx/isrXoGxtPq0N7vIYEWNxmiCCzIzXNBFc/JC1eyNcwd1wnM54r4pmwrVWWw
w47DQ7lLmnzjOBqDV8igiF8Kw64mnkKbu6CgvynkiWxdp7kNN5P/qHAC3shFf7iFVBTymLnRcX3s
05QZFgPdO+zlWAr+mXiDhYiZ49wHRnK9WyIQjZi+D7XQSqw8ucbFKRqnBbh7HkHEyQjnj8vEsMMe
3ouPLXQZhMd2rijRh968LQXHm5tr9ajk+sbiPa4qdpiO+3mm1dS91FuWPwKpIRZs3ZkvAK/XUOqK
upt+uvhlJcNOycpLj7o58PEU2gect7C/nvqRXApMuywiz7uuyVcCO2p3aXrEaNGCgwUfRlfHkKOX
gE33f0EWQUlcAhI4PIOHC+SEcI/IRf9CVPskDPIXNBVzDBQlbGfnx3pJtBBZKGgnyVsbg4maeD8j
EXLZRzIHJQvLZ2yUlfXGYQ3RXORmRN/WQuE4T9RtLSSvSfsKad++ggSA0MrlEZBXCF/6ss+ctEn/
1sgYWDI3bKKgtrhSdwyUIKIIDQvAes2bsPi6/nTyoF7Med6KLOjBBgtqqInprbAZbhJQl3yF2HNG
0JTTA6LiWTbE2izsiUvldOFAEBZAvpOpWVCFmr1tWZO8yrrY8LH/x6u8J7KafUbCoKHgcrxi/seo
8vgGe2NfPzvZ2Ed5ajU3PMKqcKvX0MrCkOkJnufnwbXAbFUlMD5bde+mHGSiTPsh08pKZvCGpHmd
GDOWSEcJDtaY4n6Q5qzI1uWeeIpjiFjMwu8f/Pwy6I0RZGewdXcps0XJLZyM9NfcTRu34r73Sd5V
JHN1PCCimrbnZxhhv+T1n43314WYwb4zZi4iEzmb0jnBGUQsWgrtYKg50icjtlVKmyJNKbJyivr5
eVuqhv2utyAX3JE+Rv47a/cUyQVXqGW4oXO9hoNA9cLttgpEd6QqW3jcZr0XMZCi+u4XF7DlYXwk
zwCGhhzIEh6VQDJk5kKlCqlNIMlpdRKesKSB3DcshwKSbc7SqlpTtSt/H4veoAA+c2Em/j+ZUgf3
rmVAFV0rlfWYHgjK+fo6saPGy2QQ7Xitn6qb6LscQlup/Mkmt8xko7gyunDScTJozB7VFoD/Svid
jRAXHQQqTv/Kb360Nbwc8vA0CBB6F0ydYpztg3Hy87BsA3JqrhVuRnGTxk3P3nSNrGCI65RNaUJE
Fch+HlR7wk2Go/zUdhZYW42cVXMDWoO5J3AEHg63ZEPjlTdHaF/dQG1AkZr6SUL8V29Z2rWjSBLI
3T0o2XPXvhyyspmLM9CdYm9oNB/r/ufAgmFRHA2Q0yVauxV0ObovjhfVbKA63bFWsxdrNu0iDXBX
Jt02Q7QzZnYtBKRPA70rIF7z1IMswQZyQYGEbG11YtrKOeTHaWdM8ZauS0wA+Gy52g8YKUXckkmM
PDXkCoAHTafMGsbqBGE9VT6/0FYsvqb5+IVDAjyIFCRPXxVM/2LIZ/qrlexaU+H6W4pGHxw4PjuF
GOuYYw1vxMNuYAFVRGg6bIfJgX2xa0w+hmRbOk1rq5UelOabTGoHoG8lMm4cSkaFBCDV7+iZDwQy
XnUyY2Kul/VKsORSE6qQqeT0agNHo6vUuTyoKb9lBkwIw1dh/3348t0eVrkV9YPNtXnn7EWgRQfC
tg75pW2Od/U+0fKgWaVpcYC9MchsrjGXie9XLvpD3Ng9usorMuXVvISWjbpIa6RAIOoyM03yFGTu
b7GI3moHomMniRMjpxnt5c0Feia4vSGBr6lV/ZLGoR/hnrHXdUDjVaNxqAsG99X+741wnK0PAOHn
AdrW8bhMPZ3xehWOuB+Jzs13IV16ljZgvWJle63a0i6d0A2ci/1ojF2kEHBf9PiwqFFJIsyZGaBY
Y5w6AHWxRzOuezVAx/JHiYtLIMIjjjEcGKhsFE8JrI4MOgsoxlf7Qp3LpUGDg+kxRr/vVmDtt06u
A5wdG8GEDNEcE8JO9RZXaY2bj92+POD3RJb0Puh2hhekvzSAe1AEqyLwiwlqrmI5OrXb9DqJ3z/9
PLVjptml2G5xvrD2e73HGVR3g7TJVwokb5U9nWqKRkECcuZUN/eVLZG6Tjdcby3bHzsFj5pLB/fY
VdyECyt2ueNaZa4vJdeVJ3MFE96H9qQOLQJfPiTxQa5yrUHZelCFgxefajbkPpsEj7okvmLiTwug
0eIjb8ZM6B5LaP0jG456tSX/uATCFnx1XWljAsBuitPptdfhUx3sYILmQshYBNIhnxLDrwwEB8Qj
TI/VGZcCdtI10lKP4HkAtG5M5ii4YwYdMujyYaeObIIKkOVdsPfTOZZsfMq9j99MZViZ6qHh2pvs
CfuoG2IvAhWtYtJ8K572bBTneFWtrdSuCyItP0LiFBMdlsha0h3vDT0CLwElIZtxyXquZX8W/YJ+
VeJd0opRt9Yqdkaso2IsARJgjkZQN1gAuFnQ/jhXgQADVdSGAfTntwnZWWkWIqkD2z6Ps1boqjmP
mfUO4BlbyyQ6tCgTxBw2JIesuvrsBqJWTO74BG7le87PeVxr6hY5I8O0adF69HRwHg2YI+pV6hN4
azJiicUvD5VBv4RcM41TjNDNMn3Ip0auW6Se7hqXsADdaAuLs3iMMuiRWu/LBzcqOmvLt1fdt7Yq
6U+wI4h1lh/eOZH4wPQlkFdLPi5as/K99AHJHboHdABrGJT1GVnZhTa1KgYOjH1erxo4yxb4VlR+
49xNrPkQt2m/sjLScq/y8m2cNlVzELiGSGYrXIahM9gMUnA0HfM5GLwABOLIMIpqBIxVPqzZze8S
osyAunAGI9rp3ZXYadnBaP3yzULXBnvZGRDJ1theKaSBWrHZ/lWwqV5J0JX6nkS9MPy/UJohgW13
R6FUHpcUySPKeEXOBBwLqoZ3pQNSAAt1LVB0mmtDIZc2RtFrOIdL/a+mhR8YHOxIzu2fZjSkHLm7
3qLJJcDtAPXQdTJo3JiYYFsQx/PZ7qmT67ZhQL9Sw/joF9tA2qsd2KIn8gw/gXYL42rYJStU4MoI
AJouhhIE7nCWNk/DXZCXKQuAtpp7Sj9kDBLyr/8xJIf84/6ZtmCRqOclp4lX7U0OlrlUzx5IVaAl
R8nEfQ3LckcHCkGw5PcVqrqmdkgndut2/EbqSZ2peR8WcW3zFdHvryhDj69+m5uHe8zSAnq5YAPy
yxDnaonRRPHV4sXZgem4ErXkRhRM9ns7Lw8Rgm5D12YGLS8coGyVusFExhyMGWGZC9lZkvIWEPqn
Tj80GDe1QnPPvc+EhyHRvrgbPpiBbjMQeNn/D2+xsUg76uREW54UbL20fNjXBflc/nrp3I8PkBmp
t/6x2Ga5P2j/kR3Jyma4sq69fCdBzgfKOjIwOoniTCeW9krWDVkE8RhG+Tl5ifRpg/854mhk2lU5
KfXwy5lv/i8R7/O2OJSfTV/8Rd1jk9an+L0y+y6kB5WI2QxITy4eOZdohIhVCOqNXgccO4c8vWr5
5HUoBp6rZuzdJbAfU/Ui/I4f/1B3GFRjSBeJlXXfMHM3xObDJGZIbgdSHEmKGS/+iid4RUi4yUuL
Z+LvtJVouirLn2OXHFE6Nek2CWgo/L0+7fx0797J4H33AAr33eEaV++Z8jSwOaYjtWZuxuH1ZEPt
I97a+Tr78x0LddnAmDq3CTXJXpbIbbFYUf17T3fdQ6h6zXp34SZYeI1Qbl8Ht+sm2MfAn3DQ6ne4
LE4bnx1XI4TcQgetW05SxdDC5NxsGNnRYGatc46PVQYppLaw5EtAJeJmvpI01Fx9nfABFbdIPyhU
otVradvKaXg8QhrS82AN24wIcJ8laJtChiwHMhpZ82bYAGOHzUNJQ4npDGTQwR9AEPfuxiZRw8K8
v/OZBHiIGNKJczBCCGN1FHhtQ9M0UpvHh3tb1MV5DtEE0m0bFfG0TG8jjMyKeaD5ewQjgjDFlVfI
LBFomlM/6ESxPMlpegxFERLtHlefGNHiRAGg0U09Ts99BKWebXKkE+iMOSVhfP69mfjNnl0HjGqe
5oIszKtoaAbMN/c1aT0PRLqbh8oetyIhC8qacm258l4R3c09GeotgdTEra8T8E/FLj0oOdnQB+xr
GcpJdmodIFBqyKXkdOEi35bbg633BIE4S4RthrUsk7Z/NZ431fpp0bh8H1HfbHkfc9dNOM4AZ/8p
f/KfNRmuxdXXqlQSWO1OyFUvZEgE3afv27D3l9w9qRgXav/PWUVVmN7rwGjVN6HpV0Xez6KayoMr
jcsRYfZbq3eqtEmHI5SN+nLcApFhsPJNmVlv0jpaAmeNbF+vJe4z3CZajla3im2H3Y5wZ6tKiZ1I
1f/NTLwqZqyKBv6OqIVHMhNMStzRzRSx
`protect end_protected
