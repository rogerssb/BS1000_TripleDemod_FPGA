`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AwDI+6E45S75vKKEvOuKiNCGUnjcAdFkuM6E6m1Y7ezjfD/zgPII0U4sc8miTOWMxK0mIJuvTyTU
Zzq3+fA5kQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
npZjabM7SDLcFCyp6I23PUa9xjRVWDHdhmXMnrES+yAJ4oT6Y9odkCvU+a7/cT8V44nH+kWRxWDx
rdH2uOP/zudERcTt/r70hF966vYLRtPhvKp/cXQVfGmZDWkkOaaorRwN06BhbEl1yaA2mOxk/GAy
xWLhunf0S2eO2DpimQs=

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Pl7T5UyPUQKbhKcNRMa5ILHn2UNqQ1JEr15Uxk+jlnpfuXcau7be18L8zpuN8QR4OZrjERsSA1Ju
xknLzH9rRoc4dP6bxM3kt3T17wJfQITyp/Vdfr2n3UJKrc6Uac7/0Tfr6smkFfudQaBf0/kpVSr7
NU0hpfcblwEixRts6b53b2PnWHxJL6ifMcguh8OaNYysP3F7bi0M/wcR1d/IKbDkL7mVKsCb/uAY
WBeXwgVfTu8qz/WisPJy2FrvJybXm47zzMuNC9JNoETwO9QETwLdiknAd/33EO5qulz4iLckgSEO
PddI2w1bDw1v+X9b7KLc2QTpJbwg7iQmqe8gMw==

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
VC9ln0bAMHicx+9d66bD6spmugA+Y33XuK+8l3waH+TQ68B2cd/in1w2mYs4NOh7K+mjTuOKi8CT
uFtgV9KtzoxaJVHZCkf3ekgIds1AVfK7ncH61dTTXrcG9TYzQPG2fSkHz9NueedND1k0+v/6gVJO
L/Lsz2LXdO2MaJKpZtk=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dGe1zqiiD7t61jy9uUIJsD0e3Sv4S2Fol3ePJlc5lALxHKmWFcrDXAtrmjGolrGJEGqdl5eBG+Vg
1yKkSbCH4BNNDbavwqAGGOcm0X0dcvMBxQhq0eiOh6rvjld7rLcMe6Nh3mbSnGFJ/RPZywPzCxk1
61GXttW9UOWEAdzo6vgiHrkk8SmnT5S42a/eCqDfQj5cdByUMBrCnEhtuTRznwZlscMc87Su802z
6I+xsUxa5JmBU2i2IWM6xNXRBhPJYOPSIiIznqWCT+NYqNT9fnuFjb6ymIDWKdlwph4wnmE/TUgm
xpdTGm8Kql9oQNrJj7DK+tmXNxpfSCaFAP1WXw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12608)
`protect data_block
fO20heXQGRnFm7xtDka25uekSSD3Li+fAtCbyz/TVSR3shcldts2jg4Ecv76nWtv4QQTHYMK+04n
GhRNMiJyzbGosIrNw9YJB0a0DgotT5+6OwuP2WhPvct5u5Dv6XHBoSkevpkpnqHselS6WX0CAP+L
jT2p6tA/j4pgBILnBp4P7k+3uhIMjf0W/Aee2HB9wj4HbL4kAMh6PkymLVwuL3i1+mj/jbU3Cb2d
X1c2D/wisxk2Qr4xMIOwod1mfhkGw0CW1SSMvQfWQEmKj9UVIXspTvnDVKP8Ll4Bwtgdi0OxCMrh
s5R40uzZJeQUEaVzl0ga27M0/JdOA47+KJgb7rJBw2OhC1L67ZFTcGZVsQZ6lqqX7/vhAqWhCLT2
KkN47wj2cR5dB4ex4nIyhKb/clBX55N2vPWFhDZExcSXiVp+3mquKP53DDzA+eb17LjZ3U8BAFZR
h8O8HKP+mMOgiaTwP35GFBRq7tBewUcWS5oyuioyEwYGW3zaOVYaF0qPBrj7qNLw2TD3WURxvgWP
J4TefrHofSNbPR9D/CVLgzpsRDJkfRjhh3JyYlhKXyXCo3vgtkL6oVFp0P2RXscHO2ZDhewnjQjS
mx/M+uOMBL8FqJ5s5j5zA/zyDKTD1GHItVPIsiXGNpeShZ7BbF8p8VCkpO/TSdfYyUer+e/MaEJH
Z7e9JaD3r9z3QsAXkAHmB6BEBYvWlb2U3+vZOPgQqWhIH/gayHFYCRm/dElYIWVBNxrEp4jC3gak
m5LuVMiWowmVMVv81uoUJ+APwAQ9ZkpHQFDzjvvW6yKgfbUgdb6bXB6Lf9Y5byMGUzBX39/HxBRa
2hi5YF7IbaZcZB8CJngn6+vNG3CXEEa3lJi5DxPxTHdkynl9mAqaczJiFWfx9vM7u6Ti5Twrqj46
6pkY/mxmkNHRVTCDWMeQKh4cOQ9/TMca1GRM1IJHvbyB60hzPdmKG4F7b5FEpaPUEoXcG9dQgDkj
/IqWZGjRQuniEQhF3hWK9MKmgxAUf4fRqYjE2aVwH2mDLc67+kzKnIdvIHbRAd4q9IlxMOH5IiHy
uHICQpS1OuX9qCEG3tj7bb1wKbyebeiex6+sUyp98ZeQa17+0ktxPVBlEzUj9LPoF0OIopGys3dd
VB/JTNWQ2oIrKepa37FMZYQOpBgs4oaFgJDg2D8lGM3rCMtUFXARVEdQb91cAWeOsd6R6ZRP1bam
uyOropO83QA+eYetWkXctqRR89/VOglegz2bwobZJQ+yMulGpt3sCmgPTZQqbEKDnf2lvGisFTkT
PoLI7NAzz6Jencg0nqwkSaIg8OffAROoyl6rptxA137P1DCZtDWX3AEP67WrszDPR8JHf1En0QqO
Nt/lC0oH4L9nZwSRZqH1MFva8RR0rPrl+StWz6IV7JgROaBsfsfOda+mKNNoS8on1+6yhHRUpkAd
76tXQmIuvZTxFH6NwuYBRVsV+JZVJFxeXjOeJaW/i1xJ/KIlRVy/PQARh66sB3TQFHtKnf/72UKU
ctprsIvbN6U1qg5cGi+HWed7yK75jy0DOFIBPPcZVv9Z2bvh4tT47owyOGWPZd6X8SHhWRLzZNM6
C8YMSq81UgTdCQpTzALzYm1NHBhEXLejlAxYIuy/AKHVrXcbeK0229zxPlmgxFRnfXbUbPxCnOIp
elBy7fPQ8vf7B8XQ7TdQyaSp1c8wqmvlhJR2sWBB27oHDzhSUhiHGN6uEP+rOywiSLSL57VEFl3a
dBcZI2O/+S8kbTgQBEMKFZtxNEFh0rs5tLts9ckbytVg6aJiHpgYvQAuy64YzL7DEf43OapOGGw9
G7NTgpneKdP4ow9ssbrzLPdye6Sl0888DPmGm8IxVjhGESrKJNnohF5bYjOdW8teE8pQ/06lD5DN
4/VfwiuUPSJe6O07jvcAQ5k2ZLUddFN2b329mk6ib+WXTmRmW3QEk2b3dk2RxCaBTUDc5EW425vn
gres5iK2wUxM6u/ihps0Mk4Cez5ruqSzdpkoIftHOPOx8ZKlLMKP1YethP6i5C3LeTkF03PWESne
R9cBA2StWJOhGwwVEmj/T45Yimh25rsQh7Qn85gWVzoUnFrmLcwaJzr72HHaCMfSwOtLe5OdvrT8
Y5QE0zWB8SSIBEaZ0+VtmXmYmj05HpzwOO3X9gUrEDbEAyyz21lt/ST4Jqx+vNgIyDTLChN1bEUg
abNhsQJ0AqskHsYrvgbYNI2LdeI4btQIljdPkhjboZzJ3dZfjwjuwTqmpBh9FYiD0LEx9lGdrzA2
Oj0oyY2mCbplgX5Y3VxOcoayJxNiWvTppViPcrYCQ2Cs9g1oN3GSeq4nJ70sQ719lt4M7gJ5UFNF
b3QCE36l2o86JlkvMpGOuwmcgYWS6BL1ZKSPac0ntDNyGJSaAxOjZsieqZDZg2PqGl4SV1nMP81V
Wmc++dydvI7SkAOY3MepMUHe4hSbHFJ1948OqDR0+9sEJuvtxuWX2ZT3SycxbkbhHtpvLmwNBp3z
tqxnrT+Of8zn3tBA2LKVZpz1LiUzxBYw4bX9Xh7xkzX9fIHDUKhfUdT/14rBNbTrz8vV8W4lYnJt
HWSaMcEZDyg/JkDqCdqKUhgNguWqHucr8qDT9fQhf6rW0i432oyovTFRQ/fgj+OSk3qkgg9bLtJE
sjj+7DNJxBT2l4XMrvLnX2VLiK1zmAjBzxmNl9JRZoQgDcT6sQ6JE8HpSDoxDYugWEsRNPtuCCWR
KlsezcbNH5H4rI+k1R7vJXLKyB/VTCqMMlptKfzcqD4HeqH7WtvB0mawAra6T9MmUdVkOLbuEAtQ
R8Tia4dBp2PIrVlllyTULYn4VV4y+fGEo7JhByF/E8oBv7EINkG9pUJJU2/ZE50Og6+E3Tx87mHC
4z8YabA3TD7cW73YYX9JlpemNVFglqshSMMzfQxvd0ibhQ20YFWroxhLPlS7VXOrreiu96KeNuQo
b2FCqZixdlSrCv9FsvJGxQVizCUGky3PTvzv6OVEvyAa8G2dGLojAUfUG+CLtrcjgE/Hn+kwwtwg
oKlU+zv6qve/kTHrKxork+w1kWAkrbpXAHvtDUGu0rsACzfTT1x5fasqXQsYSWtRsFQqc9w8jrJl
Gg7SVjsECn7Aoamd70aQ/zvH3zmtiQEVpyo8CY3dDEp8M2JWlCfChT5f2YoREi271tplP6bMF0Dh
MCF1g8yoSTH6x5mAl2vMUme/aPT5mOpEc7p3JNhMfrjuGFGABSr3EF+gCbtq29W5QI4j7hjJwfWt
yFJSu4IBGkRDWuUvJYk9lD9Nc2X/vJoJERcBI7aJgR5qggErkTCCd0qKrz9UHEIi1vcdyew8kaTy
/yTmY7iVNGnUs3jDk5XFlktb1xhV8PFNbGMQ2idLpWCsFyeZaw3/dUI6KLvLT6YizSS75PwyAOvL
R/HGCNMmhwwfPX00iJUSJQHphj/nEqhOLlTP3hT4Ky3dV2wfCKZ9BsjJKD1LH12WcEt3MQuVfbCs
FR6ggef5r3A1zeyTsROAsF6mq4pR5UvR/ABBfMC0glGnknUmE7GrZQX89dNwnxSRLWYaG/xk2Zeu
0fIVP1PHPOqa667SIZF4iEIjnyM82wLd1rCTMDKxF1VtUG2VJCHf8yHwZ3kidvSQOk4vPZvJ8bSn
CeLzA+Tu9mUIytxvoYIOtD1llCGLvCV1fXoampGGtc210AnD4WNDm/XrvYbt5nEaC0mgjUzriGUb
kL09SjcRX+IRR+lxKsENGFIbwe9LKShdFMS7A2dAyp71d1Rfvqoj61AeQ5TAEMhIOrNg/bYpJHX0
6UsX4UId4tWERGpvW/b08TSibozP7mR8DltOZc7Cw4o6dIjXENtIbpUad2CqFfAzA9Yr6hPLcJho
qKm9Ixqf9LnIh4XLJBg8J2SQxY83Bujl4N3kBJTWPdZYb6veT89jJYdW+lxbCb6NQVOnLoo2CilI
5fVRraDXj3WrnpoJTJYAykOzs4TSxwCThKQj6W1xgJFJZZVm+9Lokd8Qscjy4VuSXNlENnBfV20V
GF/NMY8cYSo3frFzkR+WsHCad12UM1bC+SnQGYpr6rlAKRw6x1dQPEMgi1onxD3p3WodwuS8CYmP
XGSlpugbwaEtr4RREQc8fSHlm61jJ08r5zHTmtRwW9CMXtnr49u1csFTzCUEd6YTpvyWjK37rX7l
fNES1L4kPhatgY27la8Uq7Ty5VWCl2Gx04fPA3rx9lljuS3wCKYdJ4DI4cJ6ubQNdAvK92XyffDr
LOLCNFiMWU4SHNK6Lj1uO1x8dDoR9fZEe8SitQciJJLTulJ8PE6OQ5B0DFa61Z3+Fa9vGCMmnb2S
xFUs+hDs3GL6mrbqoe4JC0ieSz7IdI/uIfnpL/hT4dEiPvp+G2pyOUdL3yyg4nl0i+NxMWGOYWTP
3LxjyMX2DeFGegT1vRaA3Llj2cMY/1NIQmwtZY37WTgE2TuiebO2Sa9CynmUMr8+tIN6qXS4bDa5
xJo4U/sNX9ELYy/nWBFthIKAi0hVuhcK0F1Sau1KoUkMPqGIt5/aWwLbwiYy378J8Ki7Z3C2XKRA
IRGVbPPkAe68e9bhz4aplHQJtDAvTKRiHo7z5sGLooJ+BFpYkooyD9oWq8CNp3IeyKjtcL8Pu3oE
WAaFR7bcMxHkLCJbl5VR/qMa1pJooKbWq2yaamFhBJE08y6mEQ9c/lCLHThZp5vKW508WaF4Lgr5
AbnCBczau49FhIzb/7SOxJ5UlJpxQAfIP8TFPqqKXR/9N8UFIZ+S763HWYGx/SwuAGl8AGccZzlE
r7QCeMHpIMSqJ96/lHuzx/MuyifOBJDmpiqKAjMYlw+IP5TE9ge9XE4GGcRvRJDSSf/c+scmox89
/tt0wqe1dmxxDP3bDSbRtav2d+TGEEjrPrjaIR80GIQG3cPLabOCf9+9vJvuxkd+0aCp7iykMNUT
O7ogtAhtW0jgGqOr03y1cg+v8dJzmPC16BsEnqijDztcouNzutFE1d5Wj1jocJNX0AAkAoB7Fi0F
wC0+lIfkFv/byD4EtfVwGrgN3dvKVtCMQ1vzwl58jmxkMl/Z60ovHPq6lUo24Y0xTVNfAU8jRlYB
7f4xgmgHqIY2uoMYs/BVd5zwo5lNI3EHixna41RUmdJfwJpq8tMNxkGJzXpprCcwyWAiwpro8Nhi
y445kNdyrDTgVCzUU6djexJHNp1mbL0njTfxFNS0sGAZd8eC9IjOeTWCvIBMhvcQcW54O9ZiVhJo
hCvGdEp0VHOWLD4bQi1vn+KZ7Qtl0VQltYAKUA7BAEcQ0jn/DQCDEAa7Mvf/esvQtsZSCkfmESMA
DoV7x9GdgF6xGTDhmv6Tfz00noSngaOJj5/PBfQe6U2CriUsmhQO4sTZDHnzHYqL2NR4UOHemnCA
RyfVxt5UQa4a+X1f/RRxv8tokuDCz3Up5kp1fbJGa2D35GIFgRwKJF4uCYnLqy25fPlobQdFuCSq
T6D4Cb9UzMTvLgNV6pHFKAK2iaRUMFtMJNjd2DP+hwV2Al6osqF0KLC0Ex99RTztrIC/u6uTR0vA
yJtjTlwbZnNO6fyhXyJTTqSrc3dDYxJuF9T7E2+vgJFcXXjujsCi4Ew8KZl319VfrH0vd/9sKTiV
5VXjkisDPKuZla4FybR+XjVdoeLplJ7ssdkAhQlIGI2lglDNOd/vk/litkzgow2pflZ6ZrW6CHTW
2pXpJIMaqwJYmogBq17dBKphCX3HccY1Ng403JwOewRiUF/GnpaZiWvk0fuHtVOwOQAMKEwSCDHX
JgnoNbynd4c4Ycm/Ecf/tLfASh2MMCriF8FOReKUgzQsDy9pEcKT+Q4ExvhRByYMNbg2RhgqAifC
0V0szBnyy44vgZVUe+CPVAbAsFMln+f5KI8qfWbBWiRoOVSCll1m3IHfUZMg0xd47FjazvRMHnAY
BAjr4ERNJJ4DZn3WrKHr8Sfphu6IKbsexGz6+5oiAIeacl9kq1ubJb6Zm0uQxCiCUENd5+GXRQBL
rk0mvSsGSZzB2HmCiV8Aj9OVRWthihbyUX+wDOT3AOmvE1e1RWaxZlkwdNIo8UW0Fg2kwveK5Frs
uzQ7ZZQ3TZSLe28m/hAB0I8zllBJAU/cx703bDgIDSyFZqlY6yUzzL/hZXIy7rP3hC8VtSTNiNyn
wGeuuDqLJ8XjT4VJnmDkgrYLXnHdPKFDlA5iUXYp3cjZhBQLMZWpOadv8/rNWL/WVSDs83upl0wZ
Wgz5Jojr0KOmqH1pqhPdRftUhwq/Oyn64eRul4ZtcMudW8PHxiPqNqp97ql0UetREcfUDwmgWNUN
fjWdU+rdZ1x4QLwfE220usY+5SXjwDbn+n9JtrMmZQ6/GEiZzcrx6Apan7wStXwgmGhsPlwsX1Ma
A6rJ1rjLYTos+aw+URHBYfR1g3BouPqSbNF4rAwqqRjvq9LpwAxdDXaNSUGMq6aREXZDwJ8xMEjS
fpxcZ3vMXMDQatOCXvM7ZsfY+T6S1zPV/bLwfX/Y/SzCmC6dKnCchipQPH5ToQUmm2RpHhmJZwb8
M/GSTWeBBpDDXX4p6mbMzZlawubkH6ihdpB7GTAsv3jJ3K0Vihi1isG+aEqD23toktXIR2qkN1K5
qUSX8/qrooeOOWv4oINBMRbSKvQi0pAD5ZPgHvq2i2cGIh3SDRPdnqm9gUlvYdRQ/K45Tey5ujRA
YvU14OZzKuuJPWy0lGDRRRlnE3sSZ3HP2lRy4RuiNeLYyawiWiBDrd9o3Y7LpfdofE/Dd5Cadl/M
hGc6xYHf8R9PhR8FtbwCm+o9reV+wBgBmoSgkcmDYebk9UFHTJpgtII88YbzvWbqdOSpOFRXPGTL
d1bpCfTbx/8RrgKTtSJb7cVE/suBGAkX78F1ZL0hUHHTDA5IBVnmWKNSKO7ieV7N0mzxsM1f/m29
oeqCCKXD3pSwOlrae80S9lwzozInYShg1sWXn5STMZuzZM0hMoX0VvzbnIeJHtcdIBA1Sfk8mHEl
mLVwfK2h52V9vMidrlHJdgVxNeYHid7L5rlD/oURfH74qWd9sqXlMoS54nfnlUSunlWBdZukW8Vj
UdQTh+c+ijK4KVf4d0rQipZlA4lKbZSU1uqgROcGyg/uyXjDTRVzoevpNFe9F2gT7tpB1cXic1rz
oHSMpxEc1YTADPcx3qZ8yy+Uhc92OUNdMc2sjic8JZZjKtZXfGOFVYE9xhr/73fhYgxL2iL/MWJr
tDs9f7//uEs3V7jpE4HycNFcQMS4yg3tcyLWRsxwpqBF9UJsl+2S/uuSdu6R2SuzRVfr4V0A7XvS
JdOokYCJtNs0fWgFinPSwk9NWAjxA/KATSqa8Q+imiWxx8VaEX+yodze0337VCa53AHZxQRNfNm4
nf2S49P7mj0MjbKkeuxT3kF3NBpKBVEzzUsDH71KtyZCMwCku5t6VotGBbN0YvqthZ3J5maoaG37
ClEOV2mhoL4mmHxDfgrWbE6klXcoG6dbJyHyUi6cHW/AxVkhMNnX4nmwC9U5timlEMk8enkPHba7
WFspLZEqQR8ZvSSD5POMRk75B+sM66YEBz4U8hPB+GrCi7y9C+DYSS+eShN3CM6w/+wZBa11aOAy
nmyaBpdiyNmU78qTlBWQlAeHagxw7tEKbP/mbFUWj59ANJYR9vq8s9xToCY5DjUCqBPdUmkniOGN
10P0+WXLUIoTw1KvG3lYgfpEAkNWMMuGTOLJzAQso8IHwIiFwv6dqlFVYs2DKyXqrZJMIQ8anxo4
t/NbfpJ0q0+AWLaH/fDKd+ycoIrEIIVGi1l9Uw2wvbTaaO6j1ShRblqJtlS1LRx6CESx5dT3PDcl
q4O15xxKVaHolUfAIL417sNUADL4gojJLZGl/VBXpRtG/2e2wGo0F9bjmBqdfeYG/MATj/JKs+z1
pzRY2htZiJAatvuixn9Ux5RK8LcbRnkcpHEfp3Mh2uYHY7Q48ywhLdffxVfagLr1JJ9W2KyaBnpo
hhD+sW5sI8M2S3YaLKUzmaF3NjlKKAOIBq7pHH1yi4C6lQ6SSw/VTwR8EfOr9NzBDw6KMDqYuLy5
JnbUmUN11sIm4Rr2CKCyq4+HULuH8bDNthbgdCosJVAzNt6b7QJ/nEiH44hdByZVimrAF7huNGHq
iOPwK1zXcapIljsujWarHL9T8oHtZCxSOsCPzxcg49i6MN7utcqxT1HOhV+sDemaPBgzT9lW/1XT
JjuEyel8IMBvkDzFVZ/jae7eSTKlVso8wOasdFLUT6j8IdMiMRhsaa2WhXDX9wwWHCAaWeQ4uxqY
fAfnHPPWxmeRJo5o1EziGcXg5d/tzlN4sOVwqUyafWK8rPO8dhJ2H3DvMHOBzTKKkxGWPOg38GSv
odq8QMNBGBi32MXOArGokCCNZ+fbkMyDVSdlFnnAedGtQ9kZ+0lJvnINVbS5XinpThOgCzCsZZTp
bW2Fyb1KuNke1NcDxOXAZGpEqHYxtkAR48CkmrAhlRg/u/aMmawTSXMvfrh7BJJ3idY+PCR5mNML
YPEIV2KlTNwcUxQcPZcKhLKaQjxbNfQ9Q8UfJ3lLxkcXde6HT4Eov9BO192RiwXQcWEpxvJhHKC/
5mQdEXTdlpfKasWf8x+agOIxxwFFDS04hr6Ne7VwZ/xHAG/3UAwC5BFnVyDrtM1VbzHm9fHEroom
TpbgZ9E6vMYSW312Rd9GzCGImjoj2bwnjQZAz5f7iybdzXG48vzX4s4VEH67kgKJhhgsWNhpfxv/
jCsl/hnX8RbHQ0gsMpMwFw4UtRgW6TLLRl+GcG92+V+y7oUAkBqk1E9oN2z/hVcgmeSzgR0UXXsY
vOcSnuQwQ26l9JKr94RBSOb1Cm0kfaiImA/ZiScIZretQ5ySJoFOM5YcYyuop9KXr6ga/PRXd2Ge
/v74SokjEVrtwUS3rVZW8EUQfSS/UrOy70yGuTBqF06X4+rh2+KAdhXcQcV9hqSMZ+rLUiBKuP4B
HcduDAIIDcdPGnBuWSyMfEsAWcMTzTcHVH9/ajCKw4HAzeOfqvAXrtNJ+ibRUBIVmb1uxuF+RzRx
y74iMo69xoz3VlNKnERPLZkcTIk+ZDdOpa+rk1p4U2KYrjcMVx7yrkdaBzXpFxy/Xc1ZgcPJXIG+
lwFQSBT3pmGMy21gSMxUBaBECprIEE1X/r4txjPEm64DFLtITZUe1Lx2p8vHmHC92sMe7JTthvIS
Om30NPRKdheajJ3S2pczWNc3LHc3ccjlwATWAnd997wvg2SYdtJCJOzOJAT8zz8wNnyqwNxSfZ4F
t5OlLLoyfXRzCoXgfQxX7lAWmbfsM87zjYxIIF/rgVHuDEidcr914dRP6vaHTNI5fgtQyhJTcR/H
vLCHlGimPopGQhxjkFDoTvK8eVCdPgylUESn+wj/zOfR3orbN5TkbbGANDblD9k73HSL7gCDXIz2
fYBavPpBhUDUqE+P+LwP8hy93UZKpYPGK4Kqbu0fk8Ffjz8wFKRp7D5f4LyIX3m/rrFAQ1qTT4sm
4RJgxi9Ta3OmPiWVVqkIppYvYZp34cpSiAkNqpz5MoxlL1O3rKUgHN8mSoKh4qTivEakTZUKUO38
OJEDWx6d+EHkcibHF5MwdpFi8ut6T8e9AjxQb3bONQfLeCwzoPHkI7feXjJG9+D0WZgEk6zhhVXD
2u6WxgLA8L+EIkVr8uTLWMFj0y/BVzMzIroGjjzdmWhw+CuihgZzRCcGFJ9xMGTYw8rzvzH5g5DP
11kFbkh+APyBfAgXg36B+vmkQgPonIqxZ8heO5vFeFr4jOVv4nSwQppA7GXsBxFZlSai9azevjA0
hvzmsMxcH3QAmQWRtYE5Hlsac3z8FSoFsseMKjmyfb2CxYdUBhR3M5rL6LGfYyofi24SSLAFrQH7
r+eACHUX6QIFDAg1V5meEe8F17JMfK1krtr5LbxCokOKMw87PGUhrWn5P1AE1ttbHcg67weBm4I0
3SvDD+NVkw3HUr975caWCzq4t9k3nSA5B8+jIeqvlIGeI0exQe70c3W6Ph7kbzGAF2XScxzlyBon
zKSamH3wfbSzt2PAzx1cUzRJrSuSJ2rHO9i9G4H9LxFBZpzJWniSECNwbmhLZiLJxcn3QJ09BoAz
xgawvDm6Dsh/qrX4w7MxomBSplb0VB6n6B0qVGb3cZSsUMOKIdFqA0eE9xfYHyhpnZUPocegS34m
Lm5Mju+nQietE+W3uE3Whj6ZYOjCUELbVPodRUerq7U79m0r4MXa9+C8268Nqb9Wk4lZb3Xyfur5
ZqDGMkVaroScwJgghUGTHAyHETvSJK5dOrxe4/gJpBFe63Xbs3XK3D6nO8Pev9JwOhbiRlkZaDI7
+Xr8L2/aiN2eMi2DIg9uNWe5aNeVnkhB1x46CowFipD582zPjaeOSncUeUFzfl/CUhENl+Q6CVxb
yZoGbHL/ZQcgWtQTjZzOeauL1nwoQ/qPvGn1SiHPtvPet8jTfPa9mrjK/wl6cRZQE4q6YO5EsQl8
JSngd8vDIDlO36JVrSnZoqEN3+F6K1nwAJRZ28t8E1cUjC6MdvyiZAEephclxYxyWhwmhvU9jFgu
wafMZRYNJhjf2+npUpWUeuZon1ISp8D47cUaCWG5diU5HoWfAANkY6P3AbCyy3dwypQdRyPF/PDV
tHmIzG46mQ5QMyCHNjNsba6syxJOJ/GkZTuzPpC+9OufZRs137OiKUYRTvIMPnQ6Xvzn5B9QMQxO
ttYimdIzYorSnoZ3dMiNynUtqXqpir1GFEHAH/9/4UzYhVsg9U+JkeS2XDbddt+7em6OU9xZyQnt
3eqtH1l1ki0ATnJHvn06KJ2+mrImppkKQmAjALia2XNTdboZDCuyLRCcfs5DYccGWNmX42leSGw8
YOoxl4hhNffzzolAwRykGNQpBgeFWEmlxevzRqtW53ispFWuymar7HByIx0QIeZdPNesT21cF8rk
NxqmBhBohTNkLEHGUhEJR9ge1hapsFEc6jsJhzT3xaLwXRobItfvc5/w30YCPum+SmJPzsf+1MD/
qKzgjIFfoDsPSXkt6FN8oagY10PqyKcTGZqQV6ZKPmHQzCV5udRygWOvi1lrzHGY+R3lRujaaBm8
2a72Stn03I4ups5EO8a1GaySjFK/THnucO4yDnQ+lXPfRa4wdBDKrJIBp9hV+ZGgMeGj+7H9RFxz
1TP70fNMVsCsKvfDHTw6lBTgYfiyt2wSaLBMt4XcYhF9NsBRr6GBipcfc8ZUA/hNjkIA5Vpglzo8
NjmT/vPqNlhnorfCF3I6WfP5JuMUaoslZj44x8wshhleYIGAVwqMctck8Kh4DHjgIW8foyyQWkMR
lgQA9PTCnjYUpqCxwgqsaGUapZtOij3lecGSqPge3snIB74H8Butn00F1JmClPmwsBCMt+6PEBpI
y7DdTLddh+zx+cps7V+Jkk6IdvMYilEFtHxQbqP/EkmM7TqTKTe6QelAvfwKlIR5UjLvKPaAbXki
BczYOCgXAUlVpkDmHoCS5hBVyarmMyC8YP27rVGLMlQhFvaVr98EhYtj2r9hGXvEPRT5MTF7zyvQ
HhxSUBekC+FydF+9JVYi93saXByYCDOr2nm45H/xb0aRocuppgq3naR76UIE7v86tCwgzZfFMQwT
5mFmZ/INiNR+fBdyGVO1qAQHDHkgVUs6ymhjS2CSDxMe0yJfawIeo+qzXFaum0L6BU+Gz+uur61z
8Qfg1EstHm7TA1TiUWgX/95qHLBEOLc/Cb2SPqW9lBFuxMdPLWR12/1Ywea0Z+k+ZEDWa6r/XzZN
vDFNGAb05qLyFMGRkJPouSl2bC4Y8bb4c8Em2HQ5CTGSAvy+WZSegt5Tw95O9iWOaPhy6oKE2425
AR9X6Zy8sly2H1xymHr6Gi8gcArInzQxin84mfb91JxHihrwGZ4gQT6GLBBqjsGBJAaYgveIGTqu
EctBW5R3D7boYpdpLIooew3ZmsvQrKPRupikMGB4Mc7MwITfkPzrIZIfEnjzptPJgBckZ0Pg2N9l
GFw0pwyYxQYmhfc90+TVbcmDojHGIEesYnZAefaTjsAUrRhmhs5OSF6fpjJDji1XLNa0pS2o5gLU
jA8PiUH9A48HeEa+70Zfx7CIuHBuFTM7H8R1k+v455bCqknYtBH6gANTxQVLC5ogn0MT9T+xYHfO
J6HIIawa3vSBKmkPHt9vRSPppgmrcvyRvTWQ08PvOo0XudjCuLsl3WP3cd1MoXM8zhLkpvZ603ai
Y7oNiIYzgHTJnjfndBsZDH31dVT8wzFB7RgNbOZLG3+x/ZZZ6rjs0qE1EBqBa7jCtbkU6UxzEYJX
hQnEtH9WkLgnf3xHPKP3Iu/+OSKZpSNo32TkWMRdj5BWi5CN97urByJWYZBSzvZla0O4zQFjQZvB
r8NB6aPQoD8xP1p5JZYIR26GWFRV5Jd9EnSTx0PwaV0nkkYGs171+n+hQFXBK+nYq85PXr5FIAVz
/aNH3ObkSHrdcQ5DB1rg+wXJsMH9NuY4uoYrNBTv1SarG0k76UauiyNVawxc20FKRHEM7h+xU4nV
XGBBkeOMtv0hdpN7bnYexG1j7qltS0Td+VCVWxJD65PpHyhe3wKK6XK6yx25SGODKAQHtvDoJrnZ
1h0eCicaPltqruT2jGhRlZDtxKcBqCi3GYumWnsxLOAUCcTt5+BdDKuX+nljEmDBFMxsaMp8Cwhv
cACtZTU1GIv/aQ1iSZVq0kgi1GlBTEE4c0ud4fuGKgqoTPiI+RI5vr5AAh4vnxlObDyev5iYmt5v
cdJzj+q21rhulaeqo3uZfG9ON4aqtR9jQXdAcAjOLXjSjnGj6kDWrMZ0SU+Lz/ckmF06CPAAg+PY
JgEsRbNHDI7Zf4pjeirv02jyG7uw0d7/WXHngOR1pTeXOmDP2gsFnrtmIPUi0l+Jf4ZyHm6QGYF6
a4dGqeMxcMBt7BR2f1ibxAU21iQtUTvV4QkGKxizDuklmqDsr/XdgYEUOZ/nGQ05YXw0N1wn4KY3
Fb+yc7D7m3v/vO/jwBBcPQSeW+5QMU2fhP8dtSSvNik7Zc53AFnysH4HrjF40cUPOA/p/Ux9g028
+E9sx5ffNXy/9EkwlBYia0NYrpvqPATiiNvGiLg06LHWxZTbnxiv6SsKxe4XF4LuHJ17i4Sgls3s
Hn18QRWeJYVopkj7hppoWtYzCqG90+PFSc9lU6KHBVpothYfPI6dJdrqVVQbvz6WNZtcuENt1pZS
C6bnq9p8mNlb2kOJv/xSELCMt0/vi/ACur8VfjKu7UjulgCcn6D7CM4oRY2hYQ3h521RK7FeK9OV
DTz09Mb6j0f7wgz/dWF1WVOiPJzzPYxqs2SJ77CZNvGkprxvHVMvIUkdlG0esZVBr0AOx+8GR0Nb
sDsXnbnJHutE1zMOwl1NdN4D9ukxboLreVtYc9LvqsjSDHxL+nasHeRnyh3On0kap8oKB7CGqd7z
ueZUbiIjZ/JvVFFvAWFOO08dtB2UV39oHvWmUcwkrty4ic037hWxGugrQW2LFQa4o4Yo2S6bjBH8
ywTTtacBvWxdpI0b2wgQdBqvI93sqqVf3fqfKoqRY2x68UupbqUUktGerBcbOTdXApV7s4cyQBm2
nkCKO0hi69MKjkjSr0Thf6dwiSEbLhJrqJJPVAa5wzXaBqVj0LLNxm1a3XAyk1bxT5Ic8ZmoBndu
9GUkM29tfxTpJYFmFYqUUE7M5EE37Zorl2ahhiqOkd/h+a1lKqQT/w9NouLhJy0EIA3bQMXyEHlq
mLpVkUoveS1Rt+ljgVjDPX2s35OJtg+H47+9iwlj/3KwYoPfgyTcDpGeTEmCR7djnT2EdkFeLqjS
l1BOI/tCwdRUsb28Xu+VKH01HMfclqDBHJCXGpzJquQlWdLuxqAxOXT9RsgGukDmrnFsEnHMEMN/
IWIWCa7di2MGK5OqOoUji29RPbY0d8UFpW0f/Gc/AkZok06+F2S/jh90UGl3R58RJcPKuPbTN8zE
P31lXMS1FjI+iMejHub+DrsIpmjwbdJYt06VJ0dKJDwKIggPlvwQbbojKmfrEIvwjPrXtOlhHmlf
ZFLqGDFQtkh8Lz4P9y/lsVsuMVDPqWA3sMqwFL5k8eY+15UnNhdWzjRioAVT3ujNRfSejFsvDmR8
ekXJUmTwFF6VcBNgBuEZx8JRk5uOEK+gVpSC7uis/WgSH34NyfrovVn36biIbISrpOWe4HH8+2Cc
UV4VI/Hwily4SfQkH2JWCVqLzc9IVc6yVv2Nn0lfifh48I5LwIlCUB0QshrRJqM2G551xfUnlTYv
vAv/cvyF8kb6zOxZr43jA0uh0QOR7ojHFzpHRFBmIspWLSLFlm6PGOQ/5vYNAwzJIfUQiCX1ghVx
EBDU2o03CYgYdMHaAIJEEsiaiwOwXBXz+XmoMdXwm7mLm20VCgtu/5YrJWXS5itbOZ4Wg1GZH3aR
RgnPbCaNqdsTUwmP9F0rWoMMyjxxZzuuUWQMFtgR0qxKTv2g0ej1SAa9BwT9a89vSLMmbMpY+nxc
9HJxK758fo8Q5r9kvzLUQHh58vLtE/Bfx9ein1K4SqKlBHWSs4RKNgqqpEGH92j/xNBHE7gZ+Uz7
Ievsn1LIaTQHaJP1yDbZK5iyeWlL1vwoUS/3kRiwMPhb5mAPQoCWUa+9D/o7OeNBUG0ixNqct7XP
Tr2OvY5WnGKvTnHXylOStGNSjW7Y0OYiywiBki/Cc1jiGt1jlT8S15yP+dMm+XWJONqU4tYsiMFO
Zbv/t1T6g2hSnCad4/qbL/QjMZ/UUATV0iHdylhhJ5ksuM3XEzKmLTiUfPSKZ4tyLKI1KYKm+r+k
XsxwhldOWGq1MWTroBiNTz/4ZnOwcKg4LsrTxKAjpEpUf6rGvIS4sCIECZaC0WlUFtzeDq+5/Dj1
l+n5U9avFw+KAM8pX09vql45n7zkciUL05L3IVeyr+5h+I5lhEZlwXX3TRkGMjfHXt4pY1Ry5n/A
W5gmTO8ZJMi7hGys8U61/36bpaW8bRCCjXDL3jdLfADWl/l2Sy5QzXj7o5RV0GDtkmM1GNhnO6RS
TDggeC3nSPnhnScLYt0oHb7aYa5EKcBGy2xV/BkG8I8vldEioR8HFgcy2/AuA6t4K+gSJycgYByT
NBjmtBjBZGhRYFUkXeYbXgHUpOhkvpTUdqU9OAkLg8qxQZG1RJJ+3IjNthagFgC53zexDrQRgQ51
UurWBDMndNGjyWhMrvCJt2rtVq+9gylmz5XqzuzhwzhulQpdZ0g7WOyyTetAWrZMz9S0/39rXoXb
Wuqd5cUrJBQsPw+5wqKnuXOG48baUDneN/dm3EVwy4cPdbNbV7vHdcL7QyHC+SCe2bk5IXwGBHCP
jIM+6HMtlT3T/WoiAZCxFbjWk70+QH823mVQ7bjmKPO+ag3M83IEBGMWzjN6sPKjYB3/zA+8I5MH
hFQq9NxaBv4L+xhLC9UVZYLyWRRcclniOW+Cjdz+zKZs2AmRYc/GrPt0tFT+fcmSMGBUmBTeHs+D
dtM4+dKmrhVgSp35lssdYhIpqQjauzv5G05FCrHkmmcy2bj1Irfp9wMMUBgotCE+u8k23eKO2ul4
tinJXo2p9JPb98wYXM5+rCI/MnyLLrV1H8OyImfH1LvFfDKsEouMEzy05RrBPCKGInvu+5JnHHr2
VQ3fr67n7YCk28SR+ZaGpdVaSa77JOdsWcmqDHUHO2XIYYwKmlYrJMUATW/lJTu6lpgC78qBXVbs
MYDxmavRPAzWbbhfDjkcPDjQFE5LaVOEQuUYd7Hub1+vpgjd8DSMy9D+7O9jhpL3mQOD6YoquU8W
QboKbJv95EaAknahux85F+cxJ3SNrY4Re30SOfbayuWvVLuh1L9lHLeWW2Z3DfP4ZjUgJHx7Nn9U
WABtcpoYbxRSGDPPahoIZHNOTdyPpPYKfEb8Wf3nl1HVusm0f3wldCqiLNC6PifOSt5b/QKpUe4L
vVmFQ8/AbxvRYMaF6gkkp7q9thABEdTlO2csMvegrZ61vz3qO4NYgY39TkIjzJ9w5iFRUSoIEMTz
JqI6u3hUG0O0QBrUcTic5rUBBxL+t4IvxKRiCegbfSh5blaB4aGzzrga9Dqj8L3MBrTE6ObnhEmp
7HKaVgcALhdwow3g88J3PxnFaXQx04Dw0LnVU+BvbACDHm3DjBLcdn14KsR51Vafd/vY0OKUKWH5
UzNfdwhU0ZS8sgFM9DDq313WeokNdD3b1YZc8CyUijg29ukWgmJ6AbkdvyVigiZGx0iZafPa10xr
IBiTjZyBHQQdC1lxVYmGXTRCOkqRsgLO9HPDJZIbGh2p3OQ9nqkcX8thtFYa1n1dvjwon8GWX93H
YKpAV6FdmzB3glA2YTID4My20j+6/5k99u7ZjgmUg1ZzMQZSf2Bt2tFINY9LAM/c+q2NPZPiGwKE
5lXDHghWzT1cDGGoi3W6Qlu4ujHz3yOr7Fvep2NLLbOdEHPg1jZXfao/ut/ZSkLFTiE6iwgEnwIm
pDT4zINTDkMwaQV2XdXdg4gjvLbVYF++6zrVZkvuxWt3EwwdERbjrtMeb68OyV/GWVdMBEgMJ97v
GKF5RE+PBMq3c5m3tMYWklFIzZiI2Zygoo28ye2rdcnCpCAnUFNBGXhgCSof7vYTwgpRPj6tFMv5
M+gHjHi5XPer8Y8DniuJhnxtGTVvrXoReNEPXAVXCB0DUFzWHdzZMusVlEN5JJAKsI0DZB++wyD1
LdBGJ/BSbrH9hGjrSQhi/YqHqwZ3rxaJXdO8+4prxdb9j7ttYeoFNOdPhHkIZ6XSAXnY+F+d0aO6
s+KNswb/RbTRp0k=
`protect end_protected
