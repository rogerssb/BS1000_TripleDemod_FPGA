`timescale 1ns / 10 ps

module bert_counters (
  single_test_length,
  single_test_start,
  single_test_complete,
  single_test_count,
  single_test_errors,
  continuous_test_start,
  continuous_test_reset,
  continuous_test_errors_buffer,
  continuous_test_count_buffer,
  reset,
  clock,
  enable,
  data,
  data_enable
);

input [31:0] single_test_length;
input single_test_start;
output single_test_complete;
output [31:0] single_test_count;
output [31:0] single_test_errors;
input continuous_test_start;
input continuous_test_reset;
output [31:0] continuous_test_errors_buffer;
output [31:0] continuous_test_count_buffer;
input reset;
input clock;
input enable;
input data;
input data_enable;

/* or this?
wire [31:0] single_test_length = 32'd1**(power10);
*/

// free-running 'enable' is generated by the bert input sync logic
// gated 'data_enable' is generated by the slip detect logic

// this is a formal statement indicating the data bit is
// a summer input

wire [31:0] next_error = (data == 1'b1) ? 32'd1 : 32'd0;

//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
// Single Interval Test
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~

// The start command is asynchronous
// This is an edge detector and state machine to create a start pulse
// aligned with the count enable

reg [2:0] single_test_start_sync;

always @ (posedge clock) begin
  if (reset) begin
    single_test_start_sync <= 3'b000;
  end
  else begin
    single_test_start_sync <= {single_test_start, single_test_start_sync[2:1]};
  end
end

wire single_test_start_rise_edge = single_test_start_sync == 3'b110;
wire single_test_start_fall_edge = single_test_start_sync == 3'b001;

`define BERT_SM3_WAIT_ON_START_SET 2'd0
`define BERT_SM3_WAIT_ON_ENABLE 2'd1
`define BERT_SM3_WAIT_ON_START_CLEAR 2'd2

reg [1:0] single_test_state, single_test_next_state;

always @ (posedge clock) begin
  single_test_state <=  single_test_next_state;
end

always @* begin
  if (reset) begin
    single_test_next_state <=  `BERT_SM3_WAIT_ON_START_SET;
  end
  else begin
    case (single_test_state)
      `BERT_SM3_WAIT_ON_START_SET: begin
        if (single_test_start_rise_edge) begin
          single_test_next_state <= `BERT_SM3_WAIT_ON_ENABLE;
        end
        else begin
          single_test_next_state <= `BERT_SM3_WAIT_ON_START_SET;
        end
      end
      `BERT_SM3_WAIT_ON_ENABLE: begin
        if (enable) begin
          single_test_next_state <= `BERT_SM3_WAIT_ON_START_CLEAR;
        end
        else begin
          single_test_next_state <= `BERT_SM3_WAIT_ON_ENABLE;
        end
      end
      `BERT_SM3_WAIT_ON_START_CLEAR: begin
        if (single_test_start_fall_edge) begin
            single_test_next_state <= 2'd3;
        end
        else begin
          single_test_next_state <= `BERT_SM3_WAIT_ON_START_CLEAR;
        end
      end
      default: begin
        single_test_next_state <= single_test_state + 2'd1;
      end
    endcase
  end
end

wire single_test_start_enable = (single_test_state == `BERT_SM3_WAIT_ON_ENABLE) && enable;
reg [31:0] single_test_count, single_test_errors;
wire single_test_complete = single_test_count == single_test_length;

// count bits and sum errors until the bit count equals the test length value

always @ (posedge clock) begin
  if (reset || single_test_start_enable) begin
    single_test_count <= 32'd0;
    single_test_errors <= 32'd0;
  end
  else if (enable) begin
    if (single_test_start_enable) begin
      single_test_count <= 32'd0;
      single_test_errors <= 32'd0;
    end
    else if (data_enable && !single_test_complete) begin
      single_test_count <= (single_test_count + 32'd1);
      single_test_errors <= single_test_errors + next_error;
    end
  end
end

//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~
// Continuous Interval Test
//~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~

reg [2:0] continuous_test_start_sync;

always @ (posedge clock) begin
  if (reset) begin
    continuous_test_start_sync <= 3'b000;
  end
  else begin
    continuous_test_start_sync <= {continuous_test_start, continuous_test_start_sync[2:1]};
  end
end

wire continuous_test_start_rise_edge = continuous_test_start_sync == 3'b110;
wire continuous_test_start_fall_edge = continuous_test_start_sync == 3'b001;

`define BERT_SM4_WAIT_ON_START_SET 2'd0
`define BERT_SM4_WAIT_ON_ENABLE 2'd1
`define BERT_SM4_WAIT_ON_START_CLEAR 2'd2

reg [1:0] continuous_test_state, continuous_test_next_state;

always @ (posedge clock) begin
  continuous_test_state <=  continuous_test_next_state;
end

always @* begin
  if (reset) begin
    continuous_test_next_state <=  `BERT_SM4_WAIT_ON_START_SET;
  end
  else begin
    case (continuous_test_state)
      `BERT_SM4_WAIT_ON_START_SET: begin
        if (continuous_test_start_rise_edge) begin
          continuous_test_next_state <= `BERT_SM4_WAIT_ON_ENABLE;
        end
        else begin
          continuous_test_next_state <= `BERT_SM4_WAIT_ON_START_SET;
        end
      end
      `BERT_SM4_WAIT_ON_ENABLE: begin
        if (enable) begin
          continuous_test_next_state <= `BERT_SM4_WAIT_ON_START_CLEAR;
        end
        else begin
          continuous_test_next_state <= `BERT_SM4_WAIT_ON_ENABLE;
        end
      end
      `BERT_SM4_WAIT_ON_START_CLEAR: begin
        if (continuous_test_start_fall_edge) begin
          continuous_test_next_state <= 2'd3;
        end
        else begin
          continuous_test_next_state <= `BERT_SM4_WAIT_ON_START_CLEAR;
        end
      end
    default: begin
      continuous_test_next_state <= continuous_test_state + 2'd1;
      end
    endcase
  end
end

wire continuous_test_start_enable = (continuous_test_state == `BERT_SM4_WAIT_ON_ENABLE) && enable;

reg [31:0] continuous_test_count, continuous_test_count_buffer;
reg [31:0] continuous_test_errors, continuous_test_errors_buffer;

always @ (posedge clock) begin
  if (reset | continuous_test_reset) begin
    continuous_test_count <= 32'd0;
    continuous_test_count_buffer <= 32'd0;
    continuous_test_errors <= 32'd0;
    continuous_test_errors_buffer <= 32'd0;
  end
  else if (enable) begin
    if (continuous_test_start_enable) begin
      continuous_test_count <= 32'd0;
      continuous_test_errors <= 32'd0;
      continuous_test_count_buffer <= continuous_test_count;
      continuous_test_errors_buffer <= continuous_test_errors + next_error;
    end
    else if (data_enable) begin
      continuous_test_count <= (continuous_test_count + 32'd1);
      continuous_test_errors <= continuous_test_errors + next_error;
      continuous_test_count_buffer <= continuous_test_count_buffer;
      continuous_test_errors_buffer <= continuous_test_errors_buffer;
    end
  end
end

endmodule