

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
esfZMsYAfgXl5/1NVMN2HuBLk4mXIq9zMOJXIUmxxCM3ASB4oQAFnvlT0qQ4RqGCLuc6E4dp8YY2
YfiJ3qfTig==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
frxu3a0gIGzWZ457pzmi7vYKpjmibBj5oTp3Nm6xd6yFlKPuVeOksFAqb+1Vxk7jGbsjMJnyx9lO
2VKXV4xFQMpUDAQuLbkh4Vtlfy30FgH+DdYgyNlWu+/ODzAyTBwGnqBBJRWXNc9v+o6I4rmHj7/U
VClAoMEesC6jruAbbGM=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cbNyAAUaXpeCEE3+JUKhca5KQeGFeBJanH6xxovFyeGtuBoc0MuL7wNzVB+LMvIhz4ogjiNfjFOy
erJPWJYNTjakyBQ2KCH+8XKRfXaB/2Qfhk1ktmw/8Nf/WJvgEDtu2+L4gPKqwO93MNdWTVA+E/aE
EBCYg1ZfWdcg/UPLdBw=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PY+Z0RSXvpKLK3Zrkj++I7214EYh7xr2/e4Nl8Wk/RJ2J3KnTrEGzLus2Svl+SvhU/JJwR8/pRtk
Cxuqgb2MDrHXlSxD+P9HB5/J22qYyCqHMtGZdRsOcTsKGMCCesuCLjP9Hf79ZOFvMD5UMWNYTypd
SD5yDOXbQROe5no4bzSGxG4mwA7f8MsN6m+OxrKBkJB/2o17+ooK4Myvs0AD4AQlgduQYIwshad1
8ZE/VsRTh1mVu30q0wUgNPRWy8fj8p6JpaA8jV8hCsEd1RGRrh3u9yhhQMb28Yu83JzQB0LgB7ZB
gCnOhR+tZ+mwm+CIz89fakBsAJimu/a5OY6MKQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
dNcNGxdr//RTutUgFtbRa06+j0GA1Bd7CZ0/Mk8HTgXvP7VVhMJvKvhKuAbTr0+/BlPnahR6UpYE
24CESfI57v75X+wYHFYGhsX6tZbthCLib0Sl/VTasC+DsjOCPasfshwm3hfXJtHrXq+BsUAj2e+j
SqI2/OjpNly7duOdjFzqAXOFIdm4DPfjZ2jQcFNlbTakfh68WpouAv4QpD+GeJUHYkmBgyQKKgtl
kV3c3WXWtWPT6DNWrstlDYiptICqYAAarF9Vc8+xW7gOuASapokdaHPFVyRdYaG55LKcCbBoluiN
J36ka39JittR7uAN20t1F9SkIrGeDt2AOd/6wQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eBLWtB0cBWna58k7uCx8WeEcws/CCSVLQHDhus5dw5ZePa7yqWmtAPvzy3F0qB/J6Es6WuyvqRUL
eQ3fuCXQRyh2WJZ/Kvmg23btMGY42O+kURJL/q4m+kCBbHNX4N/4Tgod+6/h76nVmqHJ2tdXDXQ/
NyPjVMueCsIMEOgWo9XM2Ms0x8mfVwKpoAwo4XM+7wuieBHw+cV9rqJpcpV+YrXad3YbrR8+OPYL
LSjcbjQlXs+TxWG6Dg/fS0HI6HuXkMlNljKnltrG7PX95TytFSyszCrrivTmqPb9TX+lTOyPVegj
yyw5GA01VXWdd1hR2C7kl1PwHuL5GhOEDAzVIg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
iDAjpnwLA8zQvUWbPDHdmHtJGVhGAluaKgmhKPZwbz6l4zb109t9UUWZVW9SxmaSiRoijqtGONum
9JW22JfnbtLpv505Uk5wbcfsEmvapDumwednQm+iuxyG1RCvvIO46s8NKYCLjgNB7i9TgPCmdntW
OkwC6bPnNFondMq+hQZHa6wTsga4K76qnnJg8GrNhzL3WD/sffBs0Fv9C9umM1G1DoJwb6PvDw1k
eiudJAXR78G3HzVioiO1k/iX1JC9qJ+80Fzoh+pin8Jr7KAeLbSFmbbWyD3gVPJVMuvwJrlFtYLd
p9NfDkC1pQ3YZxxhDDABiNcqlD9yM8xRpOs4i0IeSOKEwFu8MbatjJHfOz4b6r19rxRpnNEYeQCu
QhTbUkDWQoVGy1S6/syBuuzMiWN+Gup4FLWXE5Oenspuz3PCXIipuRc5LuNdNfphkiFcjLly3r2a
2ikXEMSJgmVKH7d4ILM8N9C9+2ihnpM1WMi06Wa3+KSiedF+FCsASwroogoO2zDUL6OWh+N7sIvf
wYH7i1WlodgBv+5IC7ukwTzGXA4oRLl9nMnWOhn/iDqeM9A+0ZCJTk6ggDx7LAN3Y1kjLT+KpL/n
VxyIiX+G5B2B3Uf4MVJ8oudl6c562dx6xEyRroRnF+7tvXTY+ZWWecnyYNinCpKg28RX3VfLsX6f
9OsC2mG/JHysctTjrzBloaBMf9zIMHWvu11ypAYPDlXlQrPvQhHvytrAlp3dyMCPZ5pUL65jN8XU
VQchDIYaptzzdrT5UphFJvZlycVrsplMv1MoU0SAMjYyOi+pl93WKyls300lsxogSkJvzqviu6d1
CjMmuyPpzhGPumHNKhOdNdsccQVoelyOToFCNqZM/DTXVEYriA742qyAyuKkKxW0ZZl7bf+2Lqtv
YYoZ8d+M7Ff1Ho4RSpJ+h4XxPpqcY1LBXFcaT96U3tqpmQ7fkPo6GdrTfXsFKfH2Dpe87UMEXZW6
MGqSS/pShIPhzPSM8SsGlJHWoMqihRI71nSopxtgUrK+MFkYd6cOoRJjIpqD6TJTQ3HfDTWr6DPk
gzG6kTlvQtRnQtvaCDF8a9A5xfQI9LmObtTuOtPSIHFZ25XZo57oTIEt3NIqCXkNKEbPVQGCYfg+
2JEE8NBkuKeSrJU6Sdud5vkqe++vuczcrODw56yXzEYaBSswhdIHpUKqhwaKSx7PFl+uicYnTEBl
JyzzL+B+FloxZmDI1/oa+UR6t0nvnX5ZX7ItFB/iHrdOfrMxx2RZT3KW0reIDB4zeraG2qGk2kSC
84FaLuoIKOjrdla6SJ/ejZTMCsaqG1aTp2+YUWdnCG+6nXkGTtHHwrKRLKuAA34ILf7kn3nPgCTy
UNE4dqZ6nf6O4c4HgCZOLwXj84FXP1YLeu7kNuyzJFh9t8zG8dAgBtJ+geBbr7hyixQ37d3Hv1iV
qYN+EYhi8J3a6795U88lz8crBncyNov/VgRV0H0UMJGCYuc94Ysx4dngLAiUUmlOmpSNVEISoHep
dud1FEV+S2IJCRCfLD9Xv3mmB1/KRYyrXnSfvIXz8No3m/EHdZCnQ6Fwa7crBBNOwyEMTWD27WGp
HnKRKv+l8fOfmD7CqrkTDVJP6DAwDuJKPAc7EFET/C6zXPFsiYF04d/OvhhgnarRL3TePhrZy9YK
OrhZ98k9b0YzggP675f+ta7s+zn3ejjX6dDSPpe8OaMCuzsJyhJa4RPKtT2jtiMDbapHPcFYSXTE
W/kCrBSevIpAt1W/XGDlG5W1mmKgS0m72fmvcEEizMN6+wTpv85qnfjGCPHm12mTJcIU8eyL1f8q
UzcT1NJMBWTwiFHD0LOXWw+RRfmmcflZ3okrLLzcC9l4hrQlD/TFKhuFuqumk8Y1/kDnvnY08eDU
5j4gWgai9zZY7XLtiWZfqHB8fCoPJ9IEJmxZMTQfzJiedroiplse2zdD7AZndO+bFlrOmMHisNjP
vBZS8sLg2uXYQohg40qyOo3dOheTo7CD55WW7JC/XVTlUXv6upydyTcT4uVfRZWxkOZv4gY5abvI
Wh3GDmQOj8bHcpi0Y4+D9F7RaGL3OKFGOx+J5sBYt86U8epEsIrPoekoT5H7SbX1mqQbNuhXMJTt
AUky8gbNtac9VG5ihkFvuC/2zeJ+ke6/6uXnE8PJZVz+Hw2txSihEBtwbbRvOzjyAhWfG+AFLnj3
z1WksecAMUFDgE3jb39WNVPGAWY9sw7sJfcLazUDFeI07mIckVNSsYABzA2ebVnvcUThZmR5Qzzi
cpaCZc9zlFbjRT+GIy4gYDSyoqsVUb/AzO3QEAmJlRrMEvUj7iHIvWSHaaS1EaYoaFKKxxhh0ZCk
+EwCNZxIf7xPQfwSLAo3VjmFDbddKRe33DMiAwsFdXyF1vfwKPVUHmvO7AVJ42RIIXtwrK9NQBIF
P/u5Gr8QiDZ9iv2p7yRsgOT9qLVa36V/PhlHblt1l88fE2aYtYDT4khhRVG8+I3x9ieY/1f9qWKr
ySIqUAWrZukjUKMSdT7Is2ZJEAdLVOzBj6pSJdbqYKIFt2hycrcgo9dVnio+SJMf41pAItpVEe7n
/i90kH4lGaFGW0E4boa5xsGl5BnD/K5ClqW9GoZKtDxjdpJps4XXG3SOxPc+ggW+QLOwGneeYqUn
nCIH0GieAP6mawA9dFkkfhOIhvBrb50INg9F3fM4al7FgqhlszWEswtQNElMqPTjm2hKIthFEzIw
nVOulA6V3vNPpeb/JItU7CPMLTIdJX1aJcin4Htw2Dkq8CrNJ+YXP+nQnFoRNK6yjXgOwn8FAOFo
UVM1rSPN0foGudEE/R0bj+UbxVz+QGT37nBo6tdi+ZsR7ewpdgQeASBc3z5ruYOSLLjR2+7+dM5c
Srp2EoR3cq4sm5g8bsE+W6uHYv9rrJdVxZ2zr/Bgr1ZzX5ntyb9EyOik+iyA6rcsHidk7Z8wJoLY
FNT1s9V0pvCMydAhVXPEOYAwJx9ASD4Cs//PkovP05Mu3V7VjbC0aa9842e7b5KcUwwRElnYtenI
jN9GfqBccEe5MfKNStNiaRkakoZghTcpJSK4hSKpeIDmTW8brfR0ZfazvHJVWW+jUIPmnbW97FKA
mGzcDkENRdSHJBfjc/jGfmfDA/oihmtCp2msp1UG+IrRcwiLLB5WbxRLkwE4uUpE+fPx3LRm/xSv
tYoLuI6NmuERxue9IhVnvrJlE8aJj/iJXaf3J6HnYLIpYWwKLaHGzXepdyaF6bVq9gUv/HYmfc+u
Dw1vHc9lm0+PUIVS9oA6g/4qWAnr1QpZ570J+iF8v0cD5fv4WvffzFPQ57VG8P7rSvLz2JtOFWm7
uYxXqxgzhilZxpPDdu1LrhUWAld6PlBNBamYxPEcWWl+dg1WoA/XCd264E0W+lom9YZbyK8kgaIN
pgz5cYAk0fq+/7BQtBjh5gusfm9nceGHkUgx+TkJgSQhs4E0wfT+2r5IHTLrzuG9JcItpWOte1o7
4bS+383QRBDEOYCBtYY0DBuXOSMjO678bq+kiQJA4tuepd2cfL1exAJmyHjXQSZsvw+JI7eHwSqd
JLNuVP+qPZUDFQcNVdQA+IelSC6L5ztSsfKkWR+yDtpsNZ2MjwGjeZQN4a5jv2kV1DtJ5zqHJIPJ
eeKL05VS6TgQ0IKDqW6PwjyQbepY1yte3g1nvHh73NJKureQS0loI7xn/ab9wOnG5gSqUzqrRKoN
gn3sGdXIAkky2dBTcVqKKi3TimlPFkBa/tdKJVf7US54FuKbOMmYQmktJg7/FbB0Mf9wXOEmpTzO
b0/FIYEXoCqttrxvCAT/NrefF0kClmYvXRNfq2a7SpqC7IXw/eqzFCPYhk/e7P0CUwsxZoFUDqgI
n9y1BW5X6wk6Ib2b1YAnlDNe38xEnH12UTcr3yhC2upwc+WmYG8GqIhTT1GfFtXH5Q9/a3U0amNx
UA4URdo+RalLEqukk6FLkTxYrPdXMMDaops61bhsvaBnCMxqSSZhr0vYzsb4id2tz2CpTSGFMFW8
REYbmiwnbIZ4Z687mB+9/mXAntHLLXsVaJGaN4+tAjaMewm/Wezu3C8DAJCbbXDe4dueyorszsY3
F4J92xfgoSshLzzDmaW+smWvaat6Og89w/KcrEMkchHdyhCqNEoR4JJUcMYyIcfD9p+v621lh8gO
FLnBxqvuHa/WlEJAuGba3BCvvVyc+SZLmQa5bBlQhEjbIVrsr8nGzykkDIRv1tOv4QPeZxO1DgMU
qKAJiyhUBhqOl8yA+E2PmF35yh3ugHQ/vrc3zc7Ian0bZNnMVwdWw7jAw2JVdnnQKGUadnasdWNo
jVhbJAwpmi0liWQd+czhT6QmEZW4OaeEvogWBh2Vr88gKS5yVm30xZ3o+Fwpw9QgOyOpRDNdSohT
u6smejVp1edN33QcYeQ1ZqM+mxRu12KGCsPepaPcbTO1oViy3MU9WZ5LUTlDwqSXtKN75jUEVWRz
Dd8xPKUY0wOrr47da4WV/nEIC01qDiDznsVJeBff3fzYA39PGQ907Vgw9hdBQV1PoKl+2wswPsF9
0eMiIS5wXZu0uqmeuJ4BWj6nDD1fDyOb0WSO6zXQCG0W3YnGr1m7b57hxelPh8+AmZO+GKDPso0L
IuiClIAxfFUUYGYGLHrcTD7qbN0i+SUMsWtnvm+0dW5acyxknWKqqEPDfNRyU4ayXEBaIB4z6uVU
Ncj1mk63ESyRBZwP0VU25U2j1zCKIoSs7tHWGHtTHskHnsIaCkYD8e2UT7k2m5UnmtKdo0ZLE/KO
vwNFV/ZD502y3cxk2O5jZA6UwPn0Pm1hV9Ear/yuoAOOJJLJ3846CquHwHCbhoCLy1KvMdZUoTtL
mFAbqn5rzYOVX/Vi3QZl08phSQ5Sa+6/WpDGYNC0lNlZlQeJQoS1bXn7uwYiUHw79t4p3wTj8T8P
9KigoBKYcNtzdbL/5l1zCGRkJhkP4ECntYgFx34nzdXfeviKUZbvRTewe2dutyEIR5kKSkgaeViI
JX9pYohe4lnjjBsW1dpn4OBEStwTggOi2VWHYvnlDtyz/nM4iEUb1chsPj65uOYshijP7LpY7Rjf
QoDY61VaDsl7HG9EvMiP3xaZDPSZuoZkI6hDMtf+6myiunqX6VGsw8a0icpoulAlY8/GrQJ7u4Ek
hSYFo17XmI+k6pGTdczJmVGXCap61tLbnpJBf0hTpAkI5g3wqqWF4XMXNnF9KzPRbB7gALFUc41e
79isNVzUwGe57cTVX2ffvQLa9EAXK25vdNBoEP3NbOKzjjc8RFaDY79AnM1zkbboH/iWSNXTIIXY
qLJf8LBa+aehZgTTy10Qf0WTOs1hn3FYrPruf6ZlRan99toqZTh4Os9WLoW9zl+8TNlIyoUZ+Yfh
EE8HYuKYqW7D4w3jhko1z5QGHPtmIrmgnKIIj+YxC+Zd3mX/d/UpG/GD01Xf8+J9lOqjdVVs8f1T
+Lez3c5Pv4dzjaElAC4iGsKoke3KvdSs6i41uBc0vtrT86cRTAs6fFMD8+x9Yf2UuoAP4AEHGVha
ZDkmfTf1cVMFddUEWv5Z8qUmEA+bn8ZSIG+jti16w2TM+U9J9Fe0aWv02V3t8D3cMI8wjTp1wXqe
fNgejp02ax9A17HIe/0dz8ufk4ME88NHmUteSMRlcNyE17zUFwO5GRGSpdhApzNyB8dfM7xiyZol
PEfkku802lMpFG4faBY8lFp5E0oDJeGg91iDLXKpyCVEOvFq05RYo9GmBVa0RsCoc/ZfFVNl/rJk
d9PIDNPdYzKR5fRwfbwZpOvPX2wIUj+oosanhwn3RHmKtynKNGu1RVgvePyXHWRvtXwiGUDGk8r7
FuF6ap8p0f+ZXLYmnHPJSeRu4+hu1Ttkp+cgDuspGZEbzntRZGmMlbVyEBvz8BsQa9mLkw0CfADV
+qWdJEoVkIrIqcNYHrqW2qlue/y21c3rDhtjV7GBjYm9LiR7l1vHK3KFPFcHar8HYVBojd5R/xlI
+uv0bQX98sRGeTmMjsxxQjT5Zo4kO2iPiWr7eU3YA3PvugcZiT+pFCbexUFoKPBW/vCErPmBmLy9
AQMfBxAZsVpqtF2k7ZTeQiZfguFHFxQVHyHpkzTHPYQn3c0Ev6oejIhk1e7ebn83K3lytx1bIjSK
NCiL1lzD00gZYzC8jD+bAj8Gx/plhku+zYVaHkF/PJ7kaoGCjEQlAJ3nOp2k+bQAH1kNlo9S0Pa9
g7NVmcsS/iBVtLYl2HScI5IKmE54kz/iWUST0go+YCwPcJPF4sZQnUEakj1FZR8UXy7SnVSrI9Td
q74gUVKoGjsUJVVFM3ZJIoOQYX82G18ytp7igACdHoW7nEW6m6MCQt+eGD+P3z82s+Yna9n+unIN
rmYA1rSoPe3j8uAJJ61X85hiFO1iED3n3OBe7zXzsrEs2ZETE21eQ8AXE9SU61bM2tbt1s5IDIEW
LdkMKFTPS1LfLnApGPWKFc5c1lvj6wC3QyB5ZMIUB+CF9FxQdWeoRSiXJLArnoM2ncf4d4A53o51
VQORZ5KxpJwEYwjPzhDAZV1XpBAnxR9zkAYeR/qmJvDPYX1tYojS70xjaP7DInWfMwtwrr6C+AId
n8OQbTMuwP5AqwHsgtFROtcJnuRgivKfrnu+8badyKMHKkfD1dRnWQTnLro/Zfu5b5mrhJZJPaLx
tqAAfEOtQfh45/Z3THOw1hDdFwzMxdGOHl788XmfujPKeZVXLVIZajNhCYeTHRQr8D8X9pxrsod0
AUb+AKFxViZ3OAUD8HNRPXsqVXKPlVL/YNvKBp2dGDMc0yYqes4DzQVuRpaRlGGCQWAv7fQKzhuU
vtRch91GROwF0AX/VDq9dSB3jE+GIvvXuj9rDMJ5ZORnEwVS0O0pyi3PJkT9zlRyjWjiMQyBffnh
PzpGdGIBx11VbLvqNhSk2bNhLU4inJgzWIyrkI50b6Lx1HbMVqTz+3vNZiC0ms/NaFW10OD4dtvN
GIbOlCiXOmGu4QYEGlEF0xY4uuJFwY/OeQIPQZ/Ya41AiOWo4o4GeIGSEpK+iKP1ump1SoiG4FvP
Pr0h2HUYiKPz5F2p21kTgmDLu3+0TAgeUiKiKIlduRPfaFK02ibpxYiUg1Cjsw79C4zKmRqe7M4Y
2Pdbo+FDi4FiCJa+B2kg68B9IHlQJ2SlgOJmyrRoQCZVqUCnFnHD5dMqCwLEOSRsMGcozqFjWFVU
wwOJMt/ojdmtmpr4BXuno0fECGhCpkFJASxFcM+692hGPxy3GdixD9lPmN3qd/WobeXxFX1yxuqD
SqRx2yFt4mgHIdcf1BQUE48M+2VHgMS5tH9tDGyZve3cjORrYvDs8XViNSLuwJVx00cZFjPIC37F
DAaMMJQdkn6DA/FXAF/x4m5X8Cmv6zUE8paiJ4uKK8BSL+N0KMqzG1a6e3w1oM2TpbqfN/yOfkDO
m3KvcQNUpBSKhI7rpSm7csIgHv1AD/JysSgH9BBXxyZFb44ekmyW7NpteVW+vRIDDQpY1+ZqGZy+
EYrhPkFC5DNbnktDHf/sWQPA2DnJWz2boZ8+D1bwQPDDmcvLOF36Ga93xzGlyKyUQmtx28ds0fb8
pkLxGo1676sGRTyze4lkly8M/nUVLPU0/IHCWtvQijpC6ThJoxX/LFVjrvYqqJOr4xWXYURma4iV
vxEEaVhxTHJstn9jStkT5DOf1yW8wVVfAOdoDmUWLOcVmvEugBscEEXFzZ2r9GCcE2bw0Nk2hIT+
u1GV8BMvyHUhcCofPhJfKOV/g7wf7LPGNBJZ55BHjzUFhxmk/vt7JBB8xIVEfhl/324j0/Xp6a2x
J55Fu3/VKZiRnIpzb95QV/cupckgvvhLiIl0NThrv97EcaQPoLpjwU/5QYbEJONxnl7VltySpLNq
4BUeUpYap8bfV1cuo/5zGi0w96x97jQJVSpIAs8m2UzLmARyUZgFncund0h/H7tImHFmXJD+Lowg
U2Vaph6YBNKlTTCCORf7/xmT00ZAlJuIhDjzoAVBVjx308EQjELiax1eO2eXCrP+2ykRrU524zz6
O/cCH34g/XkM7LwNO45rwdTy3O1o8hSGjuWWPzgGW23Fn6ANCZ+8XbFMCU+xNrNXKK5xyXxeHFgE
7ej44fiA1hK4DnhEIrCASdqMqvurSiR62x7x9hn/4uNTcqSQKXuyPAnd2zs7SW636lJPOC0TjIeF
7D2UZZCnEhOBW76aAgCX2TZOvt2egDhH+zqYZTHDz0I9wAUXFY6QtOYlHAxIS3YScx9AI311j4vY
c1g6IrU1C6or5YIiNXfm4bXY5Kbfskqf3Cywpkqo0N8gbm0scZExs2K/WT6NvwFxEeOqQMb491b4
uNHdnzm94e35WEpGQNp64WavsOCFN0yyjirpSHiIPGL6N0rXgLw6n1MIe0MUllSRuwmfWiaqi1bd
EHh+FlXTtV4aIk7VdiwUY2HiSru/FtDN0iKoOUcrpJSkfzpSixzUnRYYjbs0oXJTgKZdJoUecZRK
4wRt7A9w3Ea8naCspQ1Rt1uLUSlN12dQmmDj4A5ioMRG5FooqX+RuP7MoBmSEvhSrGN7x0gQdJaH
/4OpE4IWolhbxsEEPO9ZFL6IXaqb8EeoFX4rRUH2o6pHe7yQBgDiryKR0/xoRJNBvZKBdg8ZgW5k
E0H4/GIG/Sylt5RDAEbcB/XFYCr0Y+6Q88L1+gQKoCwI8p1EXYGFv4WE6d9Zcc78i+4tdNOdQN28
hLnxpX6U/LjhZ+CuSIco9+ckARMCt5ISjbTIXvoTTMJ62bE6qDAVVwCGdl4ON/DGQ2lz9UEBt02C
M2zFrkTb7bH87Nwx0Zj/NkhiT8NzkOm1oMKcIp8Ki4IXVDFV8pf2nfnq3VS3hwEf59LObqGN7vnn
/vxWqVEP1NUcgdcLGsEJ0v4QsxJSkHytK9s22fyAn5USc6TwH0Q11NGexGTI5AeKq9XZaG//5Q5z
olgbtOBklRQOTop3XWnrkiOqxGZaUzPW/mWgjssCHf+Ig/0wkTC+yrlDM5fxOu+umZBnlohfmxJH
r6MjWS6VV2q5tH6+MUHDJcoay9FAqHMDLOIPnZPAI0kLv12geoqOJzIr8MEpj31aEWGzDTUvbMMT
r3uvCZJ/lNt+jEF240y1dhjzx5wvCMo9Z5/rXHsiiwdYmY0P0YZJgeBFDC0IpRL1hB9E4l226keT
7OWz4bA8QeNOHCH2bZOW43rctP7VmJl9M+g3nWm+IHYTb4CHY4/qzsYPmz0q51ngPww4x3a3Jg8V
B02c0Gf1kJykwEl5F0gXA90HwAU/kDOVQmXgWRvmo9V4emT9ZawOWYNwsKmGWzWKYM5KSZTmNCqx
xo+USOqMUgxdEd7QtJRKNt9xRcPuQD2NeeE0bVRarcELRcQ9kdvJTFmuUfZww/wc/5z9E4zT+PQZ
dtApCRckWuy9HDiC1z+HX39LJFKSo6Kk4l8Gfc2mtRib2wfVcMvsXOHmUZspSuvGhihEhcL7/roG
k+eU/rLYeWpCsyItJvhcya5Vf+0wP/wp8GCd3O1tQ3ofB3DgalSCgN3lfGtLYUGA9BVLROuWgSTT
twTlKsteq5hSsA8cNtC6BnHx0y9gXMZ2O01Hw8Py3+0Xctu7WeTSMSb5SZGgPTdUCYWydsaFbVYP
oUozWaxVcJXMfju+IuNkPLfLOZnB8ecbZvI08zvUrgC+6tU3jqPEL2YrPZZQ7YD1ReTQx2kaKkxC
SNC+iZcH2Vm1YK2ESJNzDQpoZ4ieMLSxF/qNq6GZvcsLmdzC98A8h3QkXXPeIwHl64mB9ROmgLfn
FFJeyjoiI/EQAR0tDAdaKcw3f08zwX2lSf/1tdgXWujF6o9UGAm67zOa6uzqh96IzIQDAD/YP/5v
hhaisAutOnNiyeUGpVJ54JDY2ra723PbUgJakXZZQ1Y2lg7B7wZZ62k/yvUBcp3qFEi0wCC/eEQ9
w84RLnMlan62WyQRTorp+CDkb5PT0A232HWMuZlDg3rMhQ1JsPP14wi6vXwKYArtzfQi3dbV5ibd
KHrXQmsrNYD2DO4zgQ78hkuJs36FX31LbidgSQT4zJlOqBaiEAU4pOhAxKqA3nuHJ/mft0EIKeLI
gXnSHbQ05+G5OLwClZ2rvIfaE8tNz56pBMeOw1XxL8S7f43e1CR+3xuuC5WC+6SMBS7hE2cFjCr5
Mp2cIDxWs7//i7bCUfMkBsXbg8FcOM2bKlkZnkQ4Rd1pYwGQLarmIYG6IkHWR6uMuqnnHKCTUR3A
DSf+J23yDghcnySWWNIlPK9nT3BiFdvTzG3UDqruj6lVb7MsEnQbSTnwWPdb92nIQ7jrVmR3U8Zg
wxy0IepIhmN7lExc6q8Lmc1/txy+OBBGve2NLu+XIQpiBSZTyJQlIPy60atb0kCiondJGCAK5BZm
JUfylcLTftEE45qp2pX2BrAA+d5qXdrPL7xFZJFofXVDhErU9HWPCW89s2WX8FhycqFL4v4zwxjT
5LTlj4fzM4xYAX4dYpdUvh9idoQqijqoRTXVDRPO5RyB34FTbhSCGSIn+AUrWZ/aLRJqi7JAxtJz
7Y8OawPjFcaUmRT8vaem7RZdhNMpRBvJbcrHf1lLvg/5/mCu5vIOD7HKa3sI00AxSqGqXVecFOi0
etiT05kGjNHcdyBlRoFdWZBPKRVWI2G9sWMs/H/DauQod8NHNSEgZlks8Q31KW/xZMQVhaakiJLZ
1l6jLrowT5rryZvrU5XtOwHpDR61mbY+i1bpRpMWrkOPj8dRLsSXXZuhH2pSCGo8urqrRWU4HkUt
0LbE3tRw2Hj/uGR7eaFiOYAJ5WxUwu8CqlKHEpXM61YS0wU9Ysbxp6+PhwFVNVHvi1ccnH82xlo5
X9xvcjLYIUNhy7O9nMoXXb/EK/BkJPp7A+GY6m7rgJxq+oG+zwucJkmzGbUWP5QTltPPIVWgsiKn
vanKP9NoFnv69IAxCEGVaBsbcFqrdLs8ZmkT+PUaEl+Jlgm1iWsaf3Olm0OIIectO1KrTJQ9nInj
u2j/daTUn5zveFVg93irSH81JlVicKbcWxwah6ncMzh4weaEV9VeQy/EesHqGWGupjz7om7fDvLH
hOwx28AGCNsIPJyGou4Xc+UqjG+4liFJm2IEzvAvLuCPVzjepnNRVOPnKtbXdXKZhYaFZUKKuZHd
41XxEaBVehZ37QoNEkidwXzzGdktDb+FqrJny36b49r+ad4WpPpbOkLWa4ZVvZGbqT0BB/FEHvjz
15C3ImqYmojWairfOBWbWKx/UJT7J29YSMBh0mXVrAl8+w2IDPo+CueYK7eZ+/VYUSurndN8tbpL
7b9liWVNpczt73FcPkIXr2VWVaisOccKiLPFwEOxx5irrqZKVlSDHeKfU1O1EHhurJGdV3Z1e7CI
B65n4dZmvxkatmbt7TzVU3wEAUYdHMT9JFUmS2ZqfAqSC5FsiQgFqUIwUKu+g0fdnNXwhoEtagzf
/6hvGQrRf9QhOYy6wqeGlvXmfspc/5qaKfQ6+MGlqReasq8w6RWpA9+axodXhZC/b+nGdu7kgr2b
m+kZexF+SbeVoIPUvJYOBifjC+qavRHBKNgd9C5NqW09CQQy6K5YAUF9TQpzjmdVpADLYMjeX81F
oyI3hTCErjGN3jD+y0VeMU2E68YiZk36Z7VlAc0fEkhwJkSKA6Yhy3Q64bqTxNUAO5/epfIU939H
DLe1jbrchnnoYpmVnoeWFTzvCZLLtraYMMAycWZkj+4fe1Y4SKRJ2lDU0UzFZCpWIuDyKeru3xqq
ALlbRgNwkbMkV56p8AwQ/Cn4iDKlg+txb/j9UyneX7jLYFJraHKMhy+0f2/UhaUxUww6Mum3xX7b
OKuOZHR4HA8y6nyqB9jpMN1aZUYzPLxV7yPfS9Pug42sdC5XUAY9Msb1aPABeeymZ0asAG94GoNz
BDlz9oTRzi92/rzu7OZVqVMAkDPEz2nLYN7KFpHwfxVVefG/4iMYc6XjR14K5T9/dCbLxBBRi7l8
EhmURL9p2TQC05b6nL50HO3wH7NA6PNeBTY1VN3E/+FNqVu7ItRN828otaGPiKcce4WYNmbJBTN0
fh83FgoPNCTSgOCvliN4zvM6sadyMHmklvsRmWAwd/RMDEyywA/vwvcNqI+eYkNvCc4mi9G3hJQK
Inry4/Y5q7t8NFrKDzHqGpnfhDrrdrylbcHFQ4CGyZy/lv3TOxMh7tGTIaFy9/4LkqmvISCENSEE
/LVs66JCjtNjWEhn+ik+BHAEc8DofAZzzjmUzJQRblnpz9m0iAv4oYyvNcGKFXLZST3G9SgqcXJp
4btJrthExMq3kICYAKRAssRS9mVG6qvZZkjxXRpPoddqZG90AzmSHt7kvJo2T4OodN9AtV0tTUMI
+bYQl+DxVJBnRbczcf/eTUdrCudFOzbibu+fXQVgl5TzMG4EL7PEKUb00/jmRaQidv1mOLYGaZkZ
RGd7UXxXe2DgjlkCBuOFwOQTcgbVC9wF4w/XqQd5WeoaSZztVlylgaz4GNBwJslM8tsRUh818G+v
Mj1xMvIvhimv3rIHZLrJ4WKppHv6RgPj1J/T6FnWV7IS//4Ik9NtQJrvhX3ISSzsfLkoOuPOLGJQ
c96s6qmMtJtmx3RIN7WsYmUoeBaFel8iuhtGEK8OSnpAxJaoEz70k4keRGsvWx0axXq7SBsC8icc
KgwQCksQqQkJB4mZ3zTQR4h6c31WQM2NEiToYcBPC5gStrjJhk1wjNptTLPJT8kb0hVVZ4xtTy2n
9R6ajZX0BRllP9kqO3dFp3PtX2BJVQy+30y9aIXpnUSONOLQIfScILaOLBv94XHdki5jwT/32sru
C48VKOhSKpxyF1J1Teyv0OXslzCqdpNVjJVnkkEnZgGQsG6slcbflVZBGhJ9xjzzqUUh2FQ/ROOU
7Bd9M6Zci8ajvQN5Tv84jSf0GYhhL2L3UtyJ3Qu23VfFe8Xo83Zd1Fz0WLtCHQNk3q7laHFIQllM
x6gMGo0qOcLgHmtCTtyQJGUt2z8fYmTeBer7gK3ggYbBO3grDZog16/AcsXKGTB8OINTevGNaff5
30hvzCGEbEGmeivw1acGxNkZ51T90gn9QnDgdlZMshgtrHWVv34jDlS7WG77qIInD1FYfvqD4oJd
yd/ZDOWbI8Z8nkOsrwn4GGSBb2iN/KXFGp7k3i+Lgcv699FmqHMUkSKjAwMkBZLZchqQfogQUfKf
ca1Fo2mLPGz4tb16lVtu8aEo1Vh+O1er9Ooq5O/zhBBV9l4frQs365qhxKMOdttH9JEhj/NjDkSv
AkChQidI0KLTSf/xExix0TPqovLffH93NPv49jIJM4ppK02hTqqrjiG9j9lldo0XM0hRU0D45GxJ
y9GAR0leT13RlShxWsWwAhT7DU5WB7giOO+3U2NPejDXI3Bsb3OdCVnMfEWvS2AQGliRHjZfnvY+
YexWyJ716cklzAJCSsJrOsXIL+iR1xdRzKqEeJnj9gq90T6OxddHxOroues6oLzqg1fasC5B8snh
ssvhKXppqaKI5Pcj7g9lxlywZmVsmtgtQy5vdqC631/PdypGZaPizjUrGvGzxWMfw2bHASh7GyXs
czvzcjA+k9T0rjn6ayCOyR9BIkChoxiMtPdi2hnqmmhvtYlTbWKQifyQARkuKM6jGSb+NYxo8acn
ntF8657hMmlfWCVknSla/hfJygzih4hXtpRbPzY47O3DPDbqCOA9BauclsAvrhmhKpThSGEyEBpa
I/hmEEe+F6VVcBsxjTj/TteDfTO+PhBHUIOeW48h1+3VmvbaEohyv1UstOYDqv/Uby10eP6UCh3l
m32Zw5Q0EM+zgylKVrIXT+8ADic3+fv59k2il1kkkM/4SjczfKqlKhzphmTXsSIZWQxnrt4VPUBq
cpLYzjaXA67i/zUSm8syhoE6mJVZRbSB4qEizzybv60fgE5dHrRp+3p8+4mmlyKqLIc+nmvHPoVv
0YPlsWASyg0s+rOkjsClBOt/yH6ZxeoaHUxeNWGZx9kpmG92TFuNDQchap+OfhRgrqOELOcPb2k4
LxH2IfxgIkyEUHEOxlOa1+5CDJYZIAB+4voaXm5qQAQhCEtClwQ8KneT2SW5Iep/4NlJxIGpE+NN
LGvY8xJMqwR6jcqpprIJfj/FgKgXeAEGcWFmPB1/VcowFpkzlkif9XKz7hYgQTJbTHN2ihg0HELL
rUQTLuK3UaM7gfxg002JlNTpQ6AZ7rU1yUASi4NQ79NjW6oGCgkzEfVef7C8AtHIsCbtPC8NGuXc
Ip2xBoicMrzHSeQYpTs0sABUa3rOiadElvD3j0Wpd6PKdy1YA4MhYUjICpFRjRt4bUpD5rA0XeLB
Vke4mhKSB/oh1fwWzA2/cxp2AZdm8aTeJFWAnU3ZR1hf45gg0/VTBsGkH7XgpaMpycDMGc973ICV
Ht6CWWlBjV+dkYhxLSOD/7tMYuozFfOyXC38fUznBSQOZbOhLpHF1cVTsfyGNBlLr4YL50VEUsSx
ocoukxJWFVNUpytW3Z/mApv4TKToROv8dCf7yVNQx/WS7Jm92P8Bxskjw+Xowvm4anEZ5ecPXYYl
Y5+FG4PD90z7N5/pSY9hWCwLkTSYl9xJL9OfFDkpIG3PFPxDoUzE4XIdzrgQxSxfIS3HDw2LxEKJ
TdQnI8OhAfxEeHjDnsd2gXFZfLBwTCQvIeltdvjEGPy4lr0sbwm2weGyOcBvtOBUKC7eHMmiGxHh
WlDr6BoCTiQ3W64N2UQ4cMPK6u7UJBA8/mZmKpZI8YroVpoFLdTvlZaC9hUczxnBQ/DtFo98x5BD
qg6Dibuih5PSbJ6iaLp70N2lc3xhFQKgATWR/2h69ineRKgXb+a4595ndJopcDhB+r+06OQOzhLA
f+CajqidkV92mq5XPnYZ3tpJaeOzpX+QlTnt32xKuRluWFfulXkE1Y4fQALLEXmVmBNZqXYo2z8r
VW+55vHJCfohAjrLfZEukWIyPGxO2v4/Eg/yq3tgvdSnNMcl1l9zb3n4xunYIIbUF7CyVJBFQhDd
S8KQo1E6qNJlVxbKRA0Z5k6272BZAWh4gWo2UreO+EaGWzt8gANBEDMvX1Bog8JLSPFpJBsxSJX/
c7ZmerWqOlRmZksZxi9xO2r5BRKTrdiKlhxEzN54XsPhA9wndO76Z/l+pc02DPjse1sqOWn/jxff
JHV9PDmvcBdy13kkGqFBHbKCUnyLC86ngHwm2sPHyK/HKh4Z/aSlwH2Lv92jeHu6f9Lnbgj2xqNB
45BABW9qZidsxqAMHTSjl7QADFtwWg7ilE/84hc5nvrP+GqCDuo8MReciW5XV26+FxK+LWXW4IAU
boz3P5Kw0SWkuCdpHnGCTP0ekGvzUdIQfwtKzaNbe2T3jbP5r1/dwdpb6pJ3wTDnX1TG5frZBgQS
I0kKrkv2GS4TDZGOAm1xIaef/sa6Rh4t3BbB9+j4sLWk+72ivzBjqsklOV27G/tcz+3NOqAveyrW
F05lptD3fe5U/V7/8JDmCB8v8NZ2jG23m/oCJt8ejke8H0xj2DI/6jrURvetA3Uhv13X0OWyQpKV
pLmdj3j1lP627KjQfR3h1k/j/gykAV8LQaancyoGdeZV81SZ5ApNuGQ9gmrJ+Ks2BPJrChjDb5ae
upwdrbBBjFsmoOnsregjL9D8RbFuQAdDsfdroLaFoG7GSoCr5eIL/wNEMY1jM8F9v33p+8DFSbos
hkeDH+NDqM1jWc/Bw2RezAVty3kQ1QkjDjb6HZNGCgs4gHsPe1M6NJLzMB3dsPFyyXiF8rbwOayK
zlGNCGHGWUwNyj3VXinfMuprNWW/1qG2puE6EmgsfhP05R0Qdsea7w9WVmhR9aPaWPxsnlPhfBtv
eu21Fxcm39Z7FYj/jlN6Wj3XcQvYAJqBZr8bz6dDaAlFOKfV3ogwabY0YVOoiT+VE0ss1KuPjeX5
ExiiubS7xY7y9noooQhL6Q3hv8P5Ov/aA7eb0NcNQ5H6gZ1GYhBw8D2qcid9ej3KlJ3hRvicyiah
pVSOr1SgJwhwiLh2iDgN6tmMkf+xk/hSU5QmR+eV1PsFJjqnSO4kil/E50dI6q1RPIhTsUGHcknd
NdO4RhOKVVFyz6AS3kAXIF6QYbAJSG0BugfpqA7W+ee1hov2xp1vmuDIYZGHGsHuCVfZO5OUHMnK
A80MTXBefhYRNoV+AKXo8G4+8veVDdPBsVOxzMlnRCsiUzTcl5nIbfaN/szY2wqSKvJu+/dnWrYc
azaAL0VhzCa0hFVCvmL7kaIix5Xihz11Xbfv8Vo4fm9jq4Y+1Z+OYIMi/v9qc+FN1xdMv3kWrmCD
Px6DP1f2hpmkNpyXpZpeKYD/TnCsYVZzXWii/hxhLf+gP5SDCv6sYJ2cgnRkhUPZrYRrkiUiwWum
/Rg93OovTt86E/biiOkRZiwELALF+L9yXOXAfNy0tfEZEnmS0fK0HwPOcaPWFcCDd7zac3G37YQM
Yd0EMxWjaEP3bG/NTlA6W10Rm1kkrHuBLOQQjNZYMrSp+bfbW1ZqOjz+dcpb1ZVd25NIjVs/WpIA
5i0R/hccJ5K2pnYgHuozsv8Icph8Y/N42EzpYNcj4C8stIzF/rq3UeJmK2VYwHg0W5UU36ZO6Yzg
XhEHeSZzVZX9lyjopPe2wmjpVg5+AvTPXVEwrG7sXkCoc1rGp87+zFaCBXeEfeKjP0X0qR0GHMdL
1OGJT9HjFg9MRDhlYWCxAF1JeneEcW05V52RzaRJW/OzcVkkopxKzTAB87KOBdh1xCObyAuv1LmY
kBn05YoxfR5Xu5q07O48AXB6ugtyjWhVxH2zOeIfDwv37tkSCCq9tikJZTRawEDk5gwWX+ChiUNs
PZVfVWcarqXzgAJstigjSXwqOpwppgwsQfeLs3Q3ppz/J4GNhjxuUddv6Gkhrta+Vn99bR670D2e
2EsuLGq365EqFFTcfl8sViV0M41OkkL1OXgrKu1qJSRWq11XLAVDg2FT38CyPpIPlSrY3hf/tirK
jErTsrT5NEz2Y2iuv0z7M/DQJWc8f4UbDTYJS6ICzqh9tUbxhgT+bNEGdIg5aGQ7JoTD1vfPDYee
6xKdPTEiGBdsXbtqHsWUOuWb7I4LF2L2A78u3KIeSpQW9OntK5/CJttQ7fgosJLXCyyJU+w6h45h
f+EvX3tQPdV4eaLtmehzJIlvAj9myKnyuqeqFpW/7HfDiIjqsD9qpLL37B/gpL2ybOE7wvM2Yajx
bGPayQL6r2ilUynvJfpvCFAMQBPh4jEHKtdHHzXQCMIiqdaEWC4zqejnADuhrOnntSBWEk9HzZWl
O4jwur1a/5QeZbwNlcySEcivBJXMOO99m0Be4EZv/OGgBlA91HGI6h7PbR/1GjlYKjWHVZsFaBEk
hGnBUn98+1gAjnb5xuUMsIJ3o4pug6GiyTKVsoX45cXHaFazs5FlNpyjnqZ0Y/UrxaKRThsRmerZ
+a90+HEAkKNEhgqrweIuYnw5ApyI9YDRzxzAOEKDWDNBZhl4jSfblX1SClajNmU11yKowd2sHwDu
B+XE2cI3okCi1rr/T+oCYqbMNmmZoEgCI3wV+GUQgJptIYhCAgnWycANYyVd1PuFfMUynouEsi+6
PDsjVdWBKAO0uC4F5Te+93u7s7kvFNzSNtgukwFv0AFyqzmpr/oBQpZfsOv56Hroy5+u39wcoix8
PMGPJSptlKuwMndEIW553LLnrE4AcEIq04JiUAZSEMe/kwIprwdh9h6EQNZ89eKYfKwZ0PNmuBrm
W2A1o7kbHsFWUCmUYyucRG9DKpbZu4ztFHivlub9xkdFd1PoEDz37UvNctWkp8brCOZ0mLhbznww
MPYiTjiO2+YFmFXuAQhZiOCY0SlmAKLFYhy4rUoBvqwaW/sRLdgl7dMoRtnwUtNXxxVyANiD87ll
UG1kz4Ds3LmFEgyZYbNU6/dXZdx1AnOBFT/ViQyam6vhyxxZn3QfZf1lLuiuZvHn1rtSL48auLu7
2LK4TuG3evFA/vKnGZcrIol4lPD0Z7oUnGeDlauqnByNTWALFVM6uRsgKfzVeHqMV0q1UtXgXj1j
uHUjlvYYgXsjAmt8WizrKHIGS1sJ0uwsJh5fFBOtxWQ1TBfr2c5UTmBU3iuIV+8AAt6up97f9OIw
VtdGZ2pk68NSwFj2ExF9INdXzslNuq5+RZHdkktnIYZ+jDOKaXBY+AChs5EoUEg+htLHiODW1KJg
Uoia1QAkyTlNblmFDw+pxoYi7sOviJyqxjSEYYw7670d93J/pZM+JTWOAX2+u7LxOxKxcZ5mKqud
7ImVlIcAvlx0RTpzqgpFyVhUSq3fbkmedRAUumS+qi9NEkVsxKYPx7ja4mtVOvH7Ot0e1a9bE5Ui
RHy0VDfXJwzunxERs+xWaHdG39fhD4Cz8rMxJAaso7+gx5sdoFJT2kEhdGhHY43xWUpQi7yfRoss
n7DNVHFdmwftLuNFTt4qOjhZrYnL++BQM+yM8QIqwzQpNp1DMDpnPNcnymYI5WPHl1z6uy4VG7RP
h4GkmmI6CtkkMv+OJ4z9aCBtICO4J7A+rhdN5uuadB/4nzSHJQxwaxHBdeSBLPuzxjAu2vKgDnYd
zaNGK+T3TcxYXFQNetTqjzB5JO+IjIT6IF4A7RcA34RUz30O7bERW5O4KHEMY5DXfiqxFhPco6hV
kd0hfZR/HzjLJcjZWRrhsLnVaJSjp8gapFLL6xb5ksHTBj7lOnDgV1u5isde52Y1N6hAXd9PIrNJ
Zq8CAIgoM2t8gus6h1YaxEx1ZdXkQOggh30DDWSXS1Uk7O4w5DS7yeKacD20lelHmv7kaV23Yb2c
YpHtvgYtKxlxDwqODDpXPL/KMy8h2mPIUADTc0/W5JW4Pzvxomz6n7exUM2rMeLwjFQlQmVQOm8z
MPBmhWIpYvtHV+FMCdRK/z8A5bzKmZjTTNIL/FYA+Syxd0Am8Qd85dsa2FL1srVzKxUJuSCCLqAE
VKYkH7gcAp+xNWo+FEJ8YAsfmACqW3jcoGT/Sl+oWhj8DH26a38Xr5WoOUZph+tsJaYX51LJsijP
v4YXN6+Je2bHYmMl4kjiLmTzpdV+pZn1AQ6Eg7jAPRIXU8ArBi2tWNAKo7JRoEhRLIPygCjZEbjF
pDOtFrMbm7h73GHX2+Fxe831zBdmN4BL3rKT4mitLrSlL5gllKS3LUbtfPeoxjJ3B7Myq9ktOEWU
jwK2M1gpP+sJWVNa5XS0EIlPT+NbMSUKPosKdHTK0PLaeyR78TmDiVN83MO9LjLFnkkE1VrxbyA0
rhvznIJiAujXWs9+gWQ/KyJMsJuKdyHnsDf5s3z/e7ZGl6CN6Jxxa08q9bxIDXVoqA8tAyD4KxKy
cyNMm4bnB37s1gCM1TS7LbLBSx+2ZI5a71CuovnyNhuUbswn4FqdwblZCce06sOlx12eenBByDaw
YUQhyzCaD+fSrZ8YwmozE0+KnGhTFprl6Pp5+RpHWC1CM7ty+IpeGDTZbzsyx4SeFv6k3LAy7fgA
0ZKj0rVCFXP9BP6b+Cn6SlA4sRvP/baWoeGARJLCXahnF9NZ6nPycbYDYDqF9iaQttvuS0AJvSD1
+IhBq1mbvjN4JVwujymYIVeGX3TBJGvBs9PLXfpRqGIJ9ZKsLnCa/qOcbeN0Dlmm7IopCSdAQ0Rg
GXszxyiB3MG7uWvNf1tIeil6P4F/FHzi5LE02fKjwLpWbydSCWxEL1R+FdVhLU5yXrneZhRxyqZU
4WvnM+MTXnJUxBtgMAYhkRzlIRPj/Wb4C40oAFdgYCqnHDiI9XJ9BHOqEjdys1peLtp4sDySri5X
FIaGLXs9ERPhI8yLKbEjCPMcDlBmVYQMtny4q+hvh7M1mS2O8ZoP0vMyR1EiFM6WLJyOChhRe55h
H4mTkonmkwfTps058LjqXevjxaOQBiMPLcNdnnkUFFgnqIL/MMAaFhb7cCcsMs0JgnyuPFarPJ1K
6mwvwkvPyQ+KcB7I0aUW8MO6lQGoU0OqpLHi7CQiXwTQvrUpmcYSNhhgKGgWd7206CHTXt25pt/V
60f38yr5aDDA3YTJCapiphmmRPZqsefHmjzAezZDV4Wwj/+6/AlpN1H0+EfZ4OyRPLSVGq+5IoGw
6RdUb+LAsEAvGqpoXIxbRTnOD36CYEbCBAmTFtyO6zaKgajbeCV/aHLOqh5uYi+mQMjT5xhNyjbJ
jN7xluJfmH9NGMoHNY+lP2Vnzh980bg9H+9jyPpkOAzr7/66wcen1ll4PEg5suJxjc0SYd9zbuep
l58/J6uh4Ap5puzIdQwWyW1nGFpJnpuc6SgvJzBQEBxik6WezNbzDNYQjEnICpJK4ZIMwr4QyvVG
y+SWSb5L1xspWRH3xAMD1J2f7H8oGz/c2Ylz58S9NAL0w0cNmpO2WhZKC3dhuVzTxG3O8g9NP5f7
opzDQjzUKpNlyolqavesiXbZsqHs5EydUNY5Rn/m+CPECorypnwGilJt79fwSL+08SFhk9iC5jWz
ZeiSBRtgRI7KVDSKCOoj8j3BuAX8ZUgHXoFYQfzTbCDxImt5WNu224GUXlJc+WNLxLiS6s677r1C
RP/RdM/9YCdNjNlGSPHDk8KYkr5UAubh54VhKsjoydN8S8rxV4Lhrvd8vPA4yT+VLi6Vt8gcWcc7
dXSehU0WOW+SbiBYF5+K/M0x1RzaT6CTmYXdXrNui8qhFoXKIVYx0xE24K4pnq0eXjhQlKbuM3RH
ysTovwiPa5QQL73xI1xAP4sajWW0SIvdRKbd75REYeWwmV+3cfQvvm2FsSep9JtuDPUVakqbloXX
0VKKbUhe/rJ0Ar3jzAemMCLMyzmhCw1MwHw8a6fjZiGKHdzPZRRhhOfIVeKENpy/PQTZpFN5pz+A
CRcS9ZOkSgo4QV3FmAmcjj/5cUYgbNYlzVuOQHu7AQMPxlzyZ53NBSjYIa2F6jqzq/+ESJd2EB0A
GZz/wiGdZ/96dtkjwHPGYH+kq6kd3RS8ijaR5ylJogBvzLQrXafY6lXNHLsTUE0XU6gp0NqCioWw
y/xY2gmzFJD0/yT2WiwEPZOQrA6vp1S8F+qGK43f+727fvrIkGaOuq/3udWaw2SN8wsqUqu8DKAm
sLZYZj6U5YBrJZVN5+53kWG0ro/OXdSR/MLPl9oj1HU3dW94xIu+trW1mJmYN2WiIOf5oyS0HcTB
0MRvvdN5afLk09tr2LZcWQwcPm1Zzu0Kl6lJo9OM/ILDOz/XQj1bMdSYoijnwClWrf0iJX+1e1Cg
Rw42XSIK/6N0tMKX7pv+OhGpBAnMIjVZKb6DT1jVQOfD2CayvdeimjNR+PBLDN66yQK86LnDNlub
9ZuKfh4NZrV17bwXMyaLrWTh21G0IoEWv5wklUQ3/r4qlJIwFQEZPMfi6nNfQgLgUHTwJfA0e03G
H1t9wccJWdrRuxggamBLZAM0LMjLyvfoWKA0MrA2xOAZCGF6sv78yHgR2BvyKruuj1tAw5nbn2b/
7u0DMzgavVcJpzeKpZbYE7rTFJaDn4Fxyc/ZlAVMdrKbWBRpNV6L7Dn1sEPMxKNB2ucVhYDtFne2
uHt6THx7wYQnR5LmKZCL299FUFTwIf0zXE5ZWDvdE8c/YuUuKD/43NNpe8x1xw4mbE0hABKXG2m2
OpjT0LfYckVYO896RzgPU1//wbi7LEUGeEh69WY5kCtSicmLmHDwRbFHkWmf3YDg5I8j6J1XX2WI
aX+W/27vdvH5WFo3pd7bn0q4SqyNyLdHh3X+z+CZ2tPQsEcCCH86A5iVbV/GbWSf0GiAVPVrL171
9s0dYWTE2Kvv/S6QRhd0FOWoPe47wzJPMmKjNSBngSG3iqm8X6chtg4ojmuKCxaRA9g08MHU0o6C
xygkAtnotK6no/uX8Z9r4IukGnNxGPRH9ZdA4dNlcTofhHLGkY0rE+80XesnWLqyRG/fS/IgEXvp
Pdi8k6PtuoZyOaSEYNmprQgPjvkRih+b4Qg5zEs+ISN/wPcwAdDzRSgNVigZuk4l8G0rfBvsV1yP
obXDcNsHBqt2t9Swm1L0ixjnNt40/63XeQtITJIiu93jyR6k5L/ZmoCoEZxkODtufHVeKzh9BwCy
FWLFJuH9lIuNNM7rXoerCfoFmyaScsyJNZRuhywpIlG3GCA6fQ/i8olRRTs7L7pX+rr0aIAUtgjX
fOc8kRN6QYlvD5H74h5HhKZrBkKSgtpC2nwec1fpZWmcCQU03yxQhB7Yp149ScNLlVcNHO6AO2Uh
96/VesdXWaTY0QvI457/dif/vXdtCkZCPuiNFUFOd7EjdGXcQQOSIsvt+Li/Yv3dAgBeOMOT0VsK
6LZ9WicLw0K+rOClHZjCDQAN7faNTr0G6rBez9z+KpTVcI1sjDD5/D0SExVKSBRwEWo3kDjdYsxT
AtrNywa74RmuDySb0uPDy4Zat6g8jVVL077KlxnxaOHGl7dyHKZIKY5fPxlYjmZ1iO6zCc03Lgl1
+L5igeOxV40YqKxGAVhJq33eMPgLT+MNT9RdYymC0w5+4S6zlcXv7QDLBA2XvS7gXQ4RUM2G6jhA
jRsYo2vvVYMmkVA+9+xYd1cVDlrGQ58VMDSZnVpnfCpGZ1FNUcQbP8TTUinxysjQ4t3J7ycVJeZc
/VJ5YbrGnt8wkQR8YZLfFlg5ly+0wFNAACKT28yCzCPeoPrA3CnLQs3hk98UvKJbtHT8bn941mSQ
HooSpV0WuFA9ubbElO/sd7hqo3i1OtIzwg7gUj1WrKjbO2yXsKrp8tL9wO7f6ZMNng0BaUXUwhI9
eAXiTW7PF322po/4etb3FvGzwEpLeRYwXESTMGv15bQH4sxGcuOP3vhBIzkXp2Usco/tNbUutRCE
26fpkRb/60nC8CXkKVALywrZDthSRRwLBWB+p5zIFQ9DyPTTwbnZAANe2ZgK6d9LiOdFrTSoC7MH
gYDJqoSW2xohjYfxWqN8BuQp61Goeu+WC1UXtFeADZIGhKtdMeV0ViI/NGNO8kWoduLHkqlmOCXn
nCpYLyVLc9jiU1D7NHdoWoumvjN7+M5k8VDaY0KAouTipb5TbL7FyvgGYvZcmbRgVWNoNicNJRDo
eyEIkh+dtRQC+m8NYAvqH4SHodJgL5KfYbTopz1CDS7ew39zUTlbxSyesLfxd6Csht8UgUNuttGg
VOfzZ3ANJd8z4jqLB4I1yqsPFoOOQn9juPb0H4BWqupZ6ThSqoHE5nbQU1T+r2O1iMsf7dCm5Hgb
6qQTJh55OevtThSafgf9jsBzfcn5C1tDpB48qh2vYNAQRVd+Y+1KZcKJeiI5SMrXPbHYtMAgPsda
vvPkVmRWM/mC56xKZjjhFA9qFA7slNU+IviDrgh1jBB9BcZTYSoD6mQ+QGZkegd6mjF82CvQ37/Z
urWDhICCe2sfA9U6JPxbCtoA9R1P2Y2IZLzhHqF9/srm4lsfdxbhDMwQgyA/KtCesVc6UUnKlPwU
+tWG91p6r1k8wpUJ9y9jHV/qKGi5aNSv3DDtNWp7oOt/yRZUKXUrxRXnMFy2gHJTWV5w8aIMiqpV
Stb6PfwGmFx/HY/XXPSTdn2O1eqWBiJ4DD3R6yrIn0ZkzaWhAhqAhNQF4kuCCP8/A67ZMmJsnK/3
BSLss+0dTNmf7AbYpj/0RnC+CNbYp5ysKpicFVkkYc6lvuk7Cbt2h7mpzPH7MUeOU/5le1Bn6ZSK
ouJE52iqlq//1PbsOByw5FBXLowmdq2WGC67VB/DySNxm6y7aZhA30oFV7qT9uDKcUyyCHWkeflI
WxL1uLtZnEdosKo1xNBiFumule3xoLQQBNXJPdDFJXYIsJogVz0xl2plqcxbi3IMJUooBQ8zeC6G
p9wsyIta7BG6yufNfgltDQiH+s7kCblJ37ukg86XD2VLDD0e8J1JOOAl42qD8Y9Y0Vrem2cu1yAE
KN2e4bTTlx0/cbedNuR/ey5ehVsj8K7mEkDMtxy5/ZUpVWLR3xHG72BQswaP/uDFaujG1J42rzzy
svWVMQxugH07CZS5hJnEcRtv6ksecX6QsrnwUbolYqrqpXtNCm3Q7JHzzlemCcK1433ciM3jeiwh
k9fuAzS979nA3yudymMoKu8D5KbTbSqmuAnEWvy6Gl7cGmMq5tGA9P6QyIs4cvFCBA2FZB0rBACG
k21fR0l+0hy4kolcaPB0vbydMhsdzwqqYz0IiXVsAuQ2D3+FRNY9q+pbVMloYtqfFohwL7ia9xVS
9IskPkaAPbG9L3Q41AICrIyX16h1OxA3uclNpVXxM0LX2kMG1wR8W+Qm+uKABZ6qTXyCUsAxuKZi
7z62cvLVlV/2PMK8CL2s0KggtDkiJ102t77jhTZOV2XRogleGmiUdR5g0/GvcGM5LBV+bujKn7Dk
Hc6lFwybgLv2LFr6e8KU9xUs2uTOnu2XZluvmOYbYwyX+lp4dI+C4v4gkXxUfsF53Z0iInNTc7JE
d8oqUJzzLkt1puXjwgzNdhAz0siBwNEH/DJiTELk2+GBDl9yN5yLdwaUw0nCd3OXyZQ5ON00OWqK
c6jktW448JTmum2rfTHYhCQDJZIj48m8sSFGpbwy9M+Xdk4oY1RXhRmVaT3Zo9hdauwM90Vn04Dy
/viO9BGjfky5ZBYYwcrgxBmK8uYkqljkl++qCbkTBW6Q7A7U38xxrFT1V8cGCh29quUsBVnJshV6
6ec5eUZh60tZ5pHxFf8uKbf710hr5euFth+W8yBJt8OYm0J77Gh6mCBJz2zplmNA/1Ty4Fb1tNFd
nwNf8bHFSmSFiOrnfCOUo9GDpENx0BfnWVd+py8PYVf+Le4ytc2IMq4pwe/AlUT3Su0h/T5bMkyY
uRdShlLE5xM3p/I5yMLf+y7SyXirKt0qLt0/xRVU/kA0Lc6TvaGZJRRypC2mET84R8IO/yslGYEU
8xMRqqmj2v6Rs7M8n/A8apwrQy2KxJUiOolT9gP/3E8LWZor7uor7UYwT4hXsRSt1Z/AcdhkygqO
Fajrg4hLTQZgPlSdDLyRMvR/mFxZ4FIxJAYteZxx4w7FJoms8YlbHOS7W3rthX6ZS29NGzoS6+Ol
EGcCIxzJ6nFrys1u1qMyDr0M/SkCzD96sexZ5ldqYmJdWock3HxcQL6NzG4pqS9eYHStI6Gmw41r
Fj8lXsLxhio17FequWzGVy3jWvV0eZl+NIWx4yDvm2jeXc8bizNoQIicYQenRPDFiC/WzJf4Hv0w
MEnB3h8QrQdYAx4ck8BXNhf4U34zVBdiax3pSGh945vNXPSy+CEIlCVyBoGaOYOF171m/xeLmyhy
R+YdcIdHkDFtXdO03doHD/myh20Tj1x7hqbT9Vkbcn/ylMWbfO5kUO1CAh4/+vHwmMw7fU8lGMUS
CBnnY0REM3TWixTmZbOY/pp3f+e+ymv/Swqf8gy4xhVLcmRuYTCaGG48D/+y49Sx/nNIgcPeCQZT
1UPMn6nJHlAwS/Tqh7Hf7pueiZdvrEm398Lxojfd6wsCUQb1mLpUTEGHy2oR2c1IzbaJRbhK2t+/
3NOCw2A59slkTxinMyT1Jrte9dFey9K+6I02bfGuOixqhiJ6gHYFL2Bg5t7BoFd2J4YI6S7+aswi
NCZzu3+dp+7UyycQOzwEFlN6WkxgXOmdZRoGl/FJ/DOYm3XoGn3YpEeR7b7ZBSkUUqXTH4R0Jc1E
nqil+vpy+wG2hj4ryBhkJR84IG+nip4Pa5exOYAcQ6U06dTZCIpX4jSbya3pp4XtTuepAMlhL7Qm
XLQGQ4XYIBJs4OeK/2JTsCJINKOfUdvAdxgmDSeCOrmQCVufoWrD0xZBa8BgdCA7mK8GQzLGZf+W
qpIwnYAxPXaXExJd26R/jyXljiEnKxlue5fFI07ZL/o0ABE3W8DHLkC+uNUoYNAlUoayY4o+uOwB
CQV3IhkzTBaYoV58v+XvX5dLhIBjHMJZbkj+nNs+ajqrMIyi4DxXlxcNdewHAHmeKYXn2Zs4wCLR
9HBqhCxzX8wS9RcqNn/8MLYxTtoymWe11tQ+F7KJ86RBDhwBpB1m0lVlYZX/2q+omgSFeZqxsZaP
fh79tE/42VWICnTzDGqCIe5cXkK8kAQBzYEZRUQtt92hqHV+0tttpbjHltZxCmOoEXXsnNqBgcX6
FONrEYbxnTwgbM1PR4r/whnNgcnCXNI4AthmjVYUhf4PVuZgXS9Hq71GNpE3C0ohNaf5GRYPrQqU
M2UHk8PB0FIjbfLBz8cBTpZOQ6cE4gopiZ+9oj+hykHH+82GP52ePSNfvNd6Ve7nS9+RSAK4Bs06
yxFm+FzJpgZ10Y20VI5F8p0lrPPdDG0vEb45cRXFVgvFV02VK+xb9g8GRJ3YDLGh1cWLHs6TtXBb
jY1znayYIfJb+TW8cuyvTS7ATPVQ4w9qmsrtB481e8edbAXFuVKdtYvhPrMAjQNz5yb9B2kL+szt
LQBWHx9xof/JNLSCyOiJ0gQkLsQnlnY6poqYpWuzazR5Ar6/gMjmI913U1XVM5XlR47K9n7rTeKh
hVQ9y+uzKjwOSY3M/58ftn7vFMwjMEKQqPgRDE/V+2U0e8iEkJDKWyp6+4/b5RpP0G+C4+qSuLiH
IJQjBIyZc/q2+3gs0vX1PJ4FzGgDqtzkGmRKZhzeUX6C8vzsKuL1duHogyw9fUiqJlAxyMZrpVgm
Lzh0Od3ZwnElUJ8pMhqoPa4/751RYhbLO6NXc5v6uObK6aUJ5FsUypPhj6Np1xAw0rBRMQQhGlm2
GoB+tcLo22wUQJT/V/cNxUUPjN9L7UCg3bY85GBeAdlbg3deRy0es3doaUUfJ/bOsXL2WU0SVq81
MCSvCsQ/v4d2ZqaZBPt2C3Mg1x0jWIIrD1hYkHKIYtdcpQkGTY7TVyyt7gtmoX76lDGDlAlIYJS4
1tVwfqC+zZNWvlmlH92HUBmsB+MfqCpcRZCU72f63ZGOZ4KyO+sOmXo+dtlDP0VTPskpQLIXrgfH
PpEaQ7Ayd/1gYg89u5BXdb7Kx4f4VVwVXukyYWjU4iKQ8M9tgOvcerTQ3sIjP3uA5miGrz9cT+pC
LbN9WiWkDx57rVElvOWXZQUZMWp5xbKngid94NHZMXp8Scv4HF3xDnSxqTomi/j7qrdrSxEAqQWE
JuMSJzRof4GdRdP7N6hKkICYgWFIxXQchOtnZ7C7guulZHnIKkEMBHmx189kPZTzihFFCBFSOrhT
e85/7b+P1n0UjwHlQQKR2JDclI1uDRx/FS59/Y4WHG43VfEulM0ZA6NXUGQAF/CyCK+F/GJ+6apF
CCwnz/V3buspsZsy3TsPfqrsmHxBvcCNcniEiLSa4oX+TeOhgtHotCU01D3qNEx38hZBXzAbcGBO
IKqiP9V/ROidAJLx6WIV2qOB8K+Gvhb2qBMIQHwdFafxYaPW8HhNlLIHjFXMkxQaM3tm+yhATbib
mJIPbcSlGtmS82duUN9iKl2Vj8cCRHiuYx3KGKjTtV7yTzq7H8z2RIWM4h8dNLYiI3CfafnyG7cf
+GDONuwFL62dEsohtds3/6kkk6Bv+B8BUJn9D9UE6cgEXpP9vxWc5+wkIVcI/MpiJ0kw0nh4CGR5
ILMf7zbEsmyr3z1z+nFoNkLWOBPl5SCDVmlIU1y5DaXlLESnChZYGBXaoRVtum7ZPk3/07viSq2Z
w6wUFrkmLALV4hAXFIe0f4kGTYtTRWGLN6I7zsnVnxOYgafPYdYL6BGi56MhPapeebql6U+geK2s
4lPp6f+MsGxOyFK0dSS5AF2S29OMAtyh6PireVWVeigIe94LY8bEG9rDBmYA+bn4C0OYXbSKFzM6
byq8tsIjZsCV2JzQfwah64Ar+1metdC4DeJZOlf/cWUoKHOXatBRu7tqoXKOu5PncW5sVvCPaHHa
uPoRYIYVsAQdABR6NFAtBr13BMeJBxItltZkSiSq2J44ReSQle2HZDL5O6SQYVlJCu6lpKNuIgWs
8fCoQ9Yf2y0anUGTQMrLXzfN5kqmqXeRja64so3qA9BSSFqlIkkX95IGNaC7ocmDLGpW6RJPEhbu
kEgLMWRBrIbhZnQZ7N6bVsHjjWic5L6q9sMHPsZfehkQoY+9cY6rly/NvjS2K6se9Uy61fEGhh1L
CSNSJrA5Kc+a8Kqkvloiw9iXfe/FMmhkxRw+ZnGRqDMnWx56nD5i5EmFeqeCp8BtzrJ80NGtbgvO
GgBTRozeEYMgNf5WPVuHfPr2dpaC0HZZdnneRTf/YbNSvz2S791A+KwhDscK6rEx1IeS2XGc0TyH
u6MlEiTSMknMKZvf/ANtUfqsMlnsBtdpZEdXu664KLfeSUAIuUzOqsRveguSRzOtXh6qH2l2p/Ji
Cbm/wEBg+Yz84ORAyNN2uSepH8NhzSGwgFWA7S77PXHQ+qNfkmcL+bAcm5T0/pgSlzHEhrmwgLmO
E+UA3D8v9IpaJOLE8SvJNHOo6v43MFvO0bq6xIb74xuUUTsyP4JV1zA9JWB7fKWvcUL9/K61qMGg
t3JJLo1GL/6Aysa93AuHD/Qig9ASV/qdIfAoDSl0jrXReF2q/qm2/s1La2QfCoR/gdRLVepFRttz
dQiOSNtwsipRCt70553vUOSFBkSga9wY7AmLOrLvcg/F71hfnRp0utLUqkgwdQslfN6FO9oZVjKj
QQCcHv2jMxv8y6DfcrFJxSpNzEi0aFz3dmywLOYDD+4xzbTLxJ3Y5nAVm216rWIWU0fkderFSqsw
znP8q918AUYysyCXS31top3ZG8rEoy83789JiAgJ711sHbLaOAfuZ7kBsB7IczIBhS0zWClr0i1+
NFmSYNVcPPuWYU8LviiA0frVGgDESVhWDHIZGiGrj5AtXie/jOxxTHfZ4VxxHcWuTaVuUkIC4nz3
WGTaPUcIa5J8eUINEnBOvmJsrv9LJTQEIQ9/4tdRsQtZKy/vxs1HSthmU2CfI3V4qKZ4QgqFYK6l
fnWfBd3bhni0WsbxWJyA6u0oZ0TGlZJ2RZYS3EjXWi7rj4lSztcxkQEXn9XxT0tARXMaRMj8dTCC
K7ZYD2luhtOqJho/HOMsZMdd1NxCdX30Asa15AqNMKfG9hD4WM4s7sGjCB3rj/0pLu48pa0Nirte
McBrTAwzXCP6FplE8CLE887/iyAW5NuQIoicWv4sg04l7a2uaPZWOaxqrLq/KgytrONPAMZLYKrI
09CEdrSjbpuWnkAwUReM15vy16ZXPVjZ9zWr2xz/GQFVpHmZmnbBBfaMtM5VfcX4U89dUGxn9HWm
TVX6zEVhw5ip/jP2MuFasWSxjf69WyEhss9DrizYMb2+b9PRb2scO3EyTiYOqWLRDSGQfJNqFrEH
FuUvE3Jwn6dKjuhx9t7DXsfNlCWDO/V4EKBmK7WhGa8CnrRmo6g8cxIGZAKuAc8mXcc9MZqRB8fP
qCycusFtpN3Pdrvyh1IgLHvIA2jn2tIQ9Gt2QQAgz4v9E0wDrIIN/dm6zdfmPny19Rlyx+pJFktY
yNpFjWNdzw2r3EJNzZt/QK4cDV7Sp6/Og+mDxVjBigptUyhMnNFmwR5FncuCgrgyzaye0fBeNlfm
R51az+q1QpmkSJX0174wdGhmSuvKS33Q6jqeDYd3QX4lthkDLCvN1FGt6yMqcaEQBuyHpp9bETzJ
yX9gzH7MnGdbcybA/d5Timl0JTWp6KhOcmoCe7BPn9xtom5ODnZHC3BW2ddxVr6xrBBXogsvISGX
YPzZkdxFMCWcU2+rbTr2gBY+x+WK8Pq8PhVWdlGAAh13R4CSrSrqgrnvnF7LXH6kK9a0rX9s+Jjv
vsGrfYJMFZxc9SlqbOwCfNgF51/kGui6X3flqjG6b1XkfaXG4ATTc0Nwn1+Bmm8yUFDBOpkYKn59
AujWALhFZyXEitI/5N/ym5b9msMtNPVBkubsjr9IdMNKXyqWlHZmGAB6pVMR69FIno9sE9o6dRby
nhx64GlmQIaHME44JmCtaiBo4wpnEiWirUud66LKmwtfJSIufYYZmeRNKIS+axammIuX69wVWMfb
12jYJMjjUMLjjdtZZ+BNgTobNt3i1yHYFiu3au19/aW8aYoRHRP9PvtuEWPWRh6pCPiH2ZUYZ9Lo
PreioMvTAnB9ffooqb+5f2Cs6yuLpM6OfQpz9lm6FfpxVlq5U8ZseLOxdsDDJWoh2S9KQow5p2HG
wf6EhayxNplboJzY0CZqRbi886qKGhgFVkiSYOtv1aBKq+c5cdzrqwk9P/28QSyyBkTlfyao6Oyf
6TVWcNpd4bfeWjeQW5vnsPjKyRB2zYPu/tDNb3L/Eglwr/y2hBc4htIVUtbPSHygMD9TseAH3j2k
JbfdPGOiQydBgUgIvG2DPel5kDq83foSe+QNRjdnoTYfatXuoueAEoASA7AMna7vy7KhDDartz89
zg2cINKq8SojnfMQtN1wrUXksG/GN9F3OjT+z2dYW0LVTsjZD+wJ7t07vF3F5KBQfv8WOUE4hA9f
NMVzfQAqpHNZnzDkfKUnHvy4cz4oWibZEOCZKavnM7eGSQK6Sp4m2FOXRDUQqysyJ913wO3s0JFT
FxQ0Bl3w8YOulblZp7erptI/TuO3x5VQB6QLubU9YjuLRsLr+oB5oSm/otPhE3B5Q3SnneNQ8mPr
Hbcv/DU3xY65b2hXl6xH57rg1XzoakMyt8Ua5tzhQ1pFJxLRjZp2AO9VoMQXC5mc9y+6Q3VIYaDG
jy7Yiectk7TDiUzNwomLQV1slrVClCr82iXWnZt6dRKNL8gB64yg05obMGoXtJX0iHTRw9KjBQv1
JQxTtMPAqBDKRtepWM0GPYstRd0dKFAURyUePG7xHHCWCW5d3ZY5Rh1RIN4EEZHb9gYcAPQqBcyH
VD0HUJQxn862LJDxLko22/Qkk8weX3kqaE+qTiPd4xcESX5pyYpTXTn5QP7jSKN8jX3hhMK3dMAD
3Ac28uQXrdHXBB1aPm8Z2/yHXzlxkklQ43CVdMtR/zdpflRb1hy14K4xhtsqp+qvyWqrT8p13flN
YjX2/VecLHEFE5kDJZ4gjbv05IdyNCMvFSRuBQ2KdyEdiYpfPXktyoCmgUxdZBakXgWH/V1oGlNn
KWFJJYGWE+C2Qo9bDPDH2UpvXI3qWmUwsrXtBeewqNY0pbue02fAU68Fz/CxdthoBQMriHCl3C80
emQ9m0bT2K6xdt+B4eo5MZmslMeIFDcg0nFyo4rRwVF2mQ6Fh2QS7AhpAwViStZKONBgFSsOOM7f
7H0IEgT4HUFuGG0xnVCn/xc0zzhpg565QAiSASX6jq0w0bTlqMUF9vImyEnCIFTW0w048eawrmiH
meFiE5X7NbWS5i+WxGMyngcTvbFI1hqhSrwxGiKIYG47P72QBEdYTZPd+QNX9K1oR38ooAozcziP
miWCdjkPg0K3XMA7iZfMNYK8DpI6CokB97+fKVB9sxnH7p7PLExHFh0T4bRTRv/hB/QNesT0bCiA
bEeosXYZbZm+1W1IgGkwCp0vbCmAfoDjmeUny8JwAOCAGJK3zj0azt2YJsdUzCvv4g3EV4xsysLb
f7xwWtsIyb3MyvwX5dRAUkuUdifA3eIdzKnqeStJO8UDrEG21oKe9aIhALd+tQJY0kAabBFNqdrc
NE0AmDlu4got6bYi3PtmdTwd7RbfQngbK7FPrGYdlVEUSm4vDIefrsea0Z8r0o55PF+mu3/zLdHL
Ar8+rGrU/ykg4BcgNM7F8MIlJiRcKMdIcMXsfNN9voMBiM0gPucvlpf/7ggSfJaAu7Au9pZf5ZqH
X8KDS645R9nWht54ed1oe9pJQ9G9dNyeP+FnKP5aE/+jAfQlBtiAt3AFajTngTC8nGTpDYMs2qQm
hI1MiIfFOuiOkEzjfDvCRcps4BvVE/LlW9yjiZnGzfdO+LYqP1aO7mlrITLZqtoKmJk85LG8odrJ
Xw1+wBxGgr/RifObG/wKJsQWd85kyRAfIQGchLPBw8xuw79EhsxQHq3fJlizZM8Wrwoo5e5Qi8ip
xmBnofAprCbQ2pjerc99xkFsJaYx9901ky/+qplaX2CQUzTeXqwd3NmzQ2kOpco4Ov9IjnPupxtU
QB2GAOuyelOne5F9bKqCXQpxeiOul06Dw29iH2ueAVKBUKSzWwbyVj2drK1VB3cSGlzw9WVE4xHD
NFrSZ68jawgfEP4ypnGH1yw5Rr/3zWoppw5eQLgoLpgAYBU7VevHeyk9oU0zme6yzsVDvx15ihHn
tVQJ8BR+WUslZiNDYRlPn7oQ3HMKx52lEuoJiEDMQlhcRQfz1Dt6jtFZtO3QSgASGFgRkYulSVsJ
SW1Z6ZQsdUk6AvwCZtjgb2J8mEv++lDn55svdTXYQ92iyNSs9t2utSMDAy0BDC3KBb693bxY7Hqt
svovB0D93aeqgvSQ7q8idGCFIZWnyxWprxZPUlHpAyfOmnrPFTy2DcHEBXGPDJN6TiOgQm2XBoN/
pqR1N0H+Z7orAg8HgyuJ48UvT5zUAsEY9D4Ckr+uZmu6ssTXMFZgoDBZfVmOGNQfXEDkqRU5xXr2
uPew8oakCFhl/1adMTmddyb/NFPEkqdmqanFQ191Aw6X9Ud8BA/DcrWeec5vX7/6QXA7Y0qeQqYk
as8a43TbMeo9HgiNE97iq1Gt6podXc/aVTt/30q6vYE3mgTzxs9vUGLRaPeGXYpl7kD/CShSmz7/
XVlSdoEGVf5Aya5PZVAOnQefC04Z6tNQIejX4+EYG0V1F2cwA9PC+OQZGEu2H6vjAxfx/U14TUAn
GB41eZs0KfZJZtoTr1svkSjNgYXIerjmV9UeE0kUQhiukjqiyMEGSP8/Q4sGraxzRpT0Ep4hAo62
eagXDSpKA4J3cclYc13xTsZeNX2LUPMkiNP+b9fP780V2GRTMpuxXj0wxm/W7BkrP8xA4Lr3fgVJ
PGNGT65M/sbLeyJ0+z9NZeHtbKHRb2OjJjwG6rh5b/U2QIDIzK5Hvjwp+3rQPp8frbj9sA7f933x
STI/9sPLIuBCArxHVspTubwiPS7m2YXIDRuzKiLE0zEm/BWaTuOSPhW0Yq8+HIKK+3hBVjL2DiQF
y2gh54J8dD+8CoJO7nZ1awzBHV1GvOZXt/9nzWAbCMcThX0YICQ3YxJEZGCHRt9c5LfVbAyuEGmu
1Wt6JbZytPsoD4yJHZuZsWLzPjH7G9FNQTdp++6+PXlyg/fm2hy8mTAZbUiJbIXztyPzd65J5tIc
0VkhHUT8/IhjaODqjQf4ldV5YQW0Tlt2SwIUicM0c0OKk84Pd9fbA8TP7n7ykTB03ABR/ypVAYts
B0YcaTF2stk21Anw6sXQcDcOWPBl6ulV6eSkjdJIcFB56xlX60aL9LhOtVnUB4h2+w0ytiPpbT58
quU5HkdY49YQKXVOMiis4XsYAsBxDiZGZbitYBKni47YAVvY37jZCyYM0axocStkHOFX1FU9k8UH
GRjIWI2ZaYI1MFyBJ324jZcMP6JveVphdYx+gOq4jxQKhdBHR+pEkGCZDffFwPoF/1t/nXg8gNLz
w9+pLDlS6ITjjdUty926a0TguGNf9EBhbRA0seR1Fvri0hHG/JpikJtFyWCK7xzAhSbPkVppAVk3
Yha/jznIS7S5u8kp4XU4M4+trIpmtcM3SmfJjbP4HUE88I7ER/KkfeelY47k6maDpq7PmuS2ykKV
7oYsDp1SgGNI5Ej1cWVp3k945qx55W2E22KxHP/uBpzmwmfOqiVt5BrxeRfi/CePyyKnF7sK9zoy
637b3pX54LMXqluV3IzpQMPz/TABckcEtPxIfO+tPLQ+SCwIhmtMlbakdOcw7GRnk8nT1RZstDKU
M4Le8QEwFtcgFVARV7h7kEx+7NceerOfQzzzvITFa4KzkXP/EMgZ55/kGsNewt42FSC4mjBT9CeM
7qoX3ByjiDtI+MUOdKnLyLJpdln/fX7EcIawHwg91/eeaNXwAn9ox7FugFsAyVqFyjXKtblHX6oH
blH18BhNy6AviE4SNnTUDEB85vlOIH4fGGSyiKt3NXJaDlG5EgjDQ4bxt8cbFo0kfKS7UzQrNVuL
yeE/nuqsT9RtZ62oZ2mab9Lerest/If9INNh4/AWyS9A2QvUlGF9KptSSAvE5gBB56Y39yJvqACz
qcFmPN0IAiIOkm6fYFhFpwKvOHfIae9uMYobh+3XrMoLbvmOy97r7YDplqRklwu9W88v71mNR1l8
Hh2Tpa2K6thA3rFdZu1CZQSzztgFYZskfm+jf/aTSDyBfkWQcJ+KsliloV13SAVZpmBsjtkG0jKH
OsKkkNAJ38YkEGtd7PHRDX5ixXvOu1WtYsCR/mEqMDX9oa/Uteya5A3Tga944jnPv+I2xsDAKvt9
VRq22rMMMgXg+2j+xenvsFq6TDvuQyaFn136f2ErJ4SyBUdbVMxvQObni2KhyLn/teB5o5wt1b5f
/IZDFqLPfqZ8W6bmoNLWta7MNagLE0OcqtMrFLxZWP91p+1VHz9H1TkHmqia+Czs1tk5IpomkOFj
LLY6YvU7qT/gFX7L0U+1N06Iwk5bELnpDEL8qH88jviq9UkPh1WR5vqYn7hZPPAzor3zZtLfLXgj
oElLo9uyn/Cc+vVXBJD+1j8ayjBdnvkA0lJA4Msgo6jjhQQhNnE8sFOMyf7LRMuQdh1EsbQnUBPV
I1JGhzRminXUbG0b6UmHOfGknNPWd4TQZjMrjKx6Ko7Hz/VuoX/h7xo3mOhRMHK8yBqmUcyMd5Wi
s/J/yuwPiILVvxtXzhemjZIs5scKK2gL3pJtUg8VapGbk9AzQNJFqSjD/p3+c9DseKKu0qbUcsCO
X77S3Q3wbie1vE0w9r7bS4InVl3NdJ80nYLllSNOtDVMZQQYUWTy+CLhL4kw0jfnc6WRGpnmcNZ6
xk3+sUfJgIYj2FVELKWzV51MTZwDcWvJxoUlg/AvgW7u660jpymO7+PgmrlZfqFhnkXopdZdY/rR
YZJz113R19vlnAaL7BGzTGxWVe+66f5AK+19Syu0G5SyiD6PBnjGxFxO10aTXYNO6aiXjewDovs8
W9coLp7neZ5bVGiI3u5LVBZAxNXaSlS56T6rfWzWGKkIkq5NAYA9Xzxw9uB5HmeOqooWXMXtsbFN
RQJ/YLrShMRVTGIR7htOgjuLmNxc+7bRh+32lHWprQLi/1IPJAG5ZzCASpIjY9dMq8tez8OkW3J0
zEhNpPYC3eqQKeAPcEjPvjOdF0VED0BbXmCOEPEPJtuDLG7oScoh3z99XMPmk+t2ipbS6Wd9qAJV
iy55hez8XituyoI3M9EPfUP4YSPAp5faaqh98jpkCmFs5R9vuHEGrH/uLjBtqK0hBLEWn4CMcpKJ
gLj2tFkbm+7mxRhxMwG57t9m3QCw/08nSjSEx6Eb4HLKcSyQA9nwqhyaK4ZsIfN5eBAw4Pmekcid
dfWfi47WBJheIB8IwRuDADyGr4VNrsOSli6pgFvaxXBdz0c6jgakGVO30b5bqKx2hC8ctSHJKt2d
I4/KMtSiQHjs/iSjMevG7q3fz+UBZahzx5IPtwphmWI0ekb3i3T6/KwWWSaf2tnKdcBk6tSlxa75
M79ocHQD1Csgz8EI
`protect end_protected

