

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
WL7bD6pbPqaR89V/S2FlNYnU4TVqryWuNsZvmZfyG4So7oZUWkx+PkfJLlz41bGI81EcFfaGw6LM
8o2iHiwkRA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y0rsKBYuOvwQrBstDYcyIsVKr5/7no2EdAEtH4RPd+GDMzK44r5BWYLlK0OcMn+a1crJSQYCzYMl
qmOWlOBf8ah3f8POgqEbdNPVaV9YYTipmqM4AjpCbGMi91/1QoRZMxajkqVZ8N48TGg4cP/TJjRi
4z2xO37DwjjjRJS8hXQ=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
odx6xN68VnStEA95qQ371eFjHiKmggjYaPuhvby95tCA7ggfuoEv7351+PKASqlPGeFvPABoRvXV
qVezpgZcyEuPWbWyTwJzg6LnXeWorKGgq39UF4gKNTjWOKClYfJSjSFxnMceEaXYU61VGXY3x4jL
2WGEMebnJIK4xkzoRYQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
X/YWLHPi3Jqkx8MFxH28553A/zDDHAl66wu696jynq8LDdGsP1jOBEnegUxOtIq0XPnmGGWfuZCM
vqqYP8qLAz2XIPBU+IUw/FRBBrgSORB8iH1szNI73ElZbQGxSDirBOGoX7TsoJYyRBxA5upyh1uv
HpqzgvcFV3B9zyMncS+LM2ikhWJ3nVyQX56yxZ019DKH38UTlOL3scdmX65rURjGj0RBwiq3cf6Y
Q4Vfz+P9XBW3rHBJ4YgfyNbFj4sWNtSCSgdh+opBLi+WCZwmS2/ighKiRznhmqv0g3/ndNE8dZGS
5FqK39Oeq+Od/+E4Kk9oEX34wcmUOvfTKMuICg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ve9WLWlb1h84Xh/gr+AY2Ny8lA24U/qVeWlgQDA5KV/atwKR7gW61PuYudBQTGl+gOvoctOBYQE6
67pi5EJm21rdxQffmdwk+TN6wg4egIHw3uazWcwbaL8kAaOh7ot5rgHN4olfcoHP9dUVpWkLzABa
I75VI8adqGPWckC/90YJ/wrJ8Pnwumpe3TqPtkIN0292SW1XfxfVtBqsebK8XCMgOmvU8sXB00TJ
wwlROknoSlSYyCMZs36en5PnLvjqDzFRRaM31mxFyogld2P0T3PXh+Vw5S9GR/iyQ2owQMWIjC7V
s/phIy4InpaIi0cD7gNvdXAzhjbLo3QpYFKfyw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Tjhd6B6bcZ/gaw2CE9cvppas8Kf7kdlRWjxcOefJLT7hqmFnwna6ZlwPxm4BYzIm5Nc5MmV4xaCq
qpsSxy9wrlMU5AfwQQvZve2SzGbUJ9uD8/24EPEQtibNMK5M8MZcXEfkx/294Tscngnkxrts8Ppj
UfgAiuO7BqcKHIkQQn0E1Mvc/SEE58m8pi7HE5lP48wwufDxYPcPDttvqxcY+OKAwoPQTbDLTTA8
ee/4xcIw7R+AhpOAs4ypOis3MMyghozPf5or9bRn7NnDNGacrsCuUpLlc0P95tBGvQPYCi/pwFrh
SJyUZAckQkV61xVr0GuCzls8rwKzVfMDqITHGg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 211312)
`protect data_block
j+rWJZE6lJDmFgTf0q9UQIkK91RY20+Cb0Kl2+HPnlt1A0+GcGdizX9r3JYPecXQHHpMLuVHXoyS
SN/4+S59X7/9WyNNZ32sUPDIF57Dw6ceQzF55h451zkZbh+peN1br35Oeiekb9+UWlDbs+PuscTM
xohvZWQnXeQIxi2MeBJFHUTqIouN6OQm71lfgeoq90Uzclyf2Em9K3mzlhCYkoOqA7FpcE3CniBP
YDGeMrukQhsidl2whuHislf7COMlleZVwXDGnfk2MsyFkOtgNrIQvGMFnyyVMH/bsISXWMHaNaJS
FmbEv35MExxDKsnRlgIQC8WfFUhONB14ubXEcuirGKbE6WUagzerwvVt2rmMrRe23SkJi4HjcLpc
TnVrYdwg06ldP6U1hblbfeI6vIewB45asec3+hBVszti/Lt6dHGsWR9JuopyK9G22+/Ntn/9diGJ
I/KDrmEXq9XcN3F3aOeovoDPQdxouP0LG6lNr6hyFvqt5uJ7lxBuf1xMNGOKO3QwQN/F0jeYocKh
mUAkRqoXnWivPXaGiHweHHv6FYfHMAHj9YQ0ImJRpELQz0hCIJh8ad1Rr1g3OHOPLLjOFzCoaq5V
EsdB7qK5Mb7A+yma/jcC5sOTNhxmu/P/kCGgQjZSi74Mdo+jijyxvZaMH5CbKyQNliL3JgCbl4/N
9NCk7LqrhLdHf+Nm/F095rpoEJPV5QQ3uxAmuEoqiy4SqUXs2VGJPxu0T1qBrEVu0miLh19GHuVX
J+NRn6biHqQOHxSqlW5yh4gGk2c6RlP5Ld5UjOoJcA8AkVIesmYUYhvoyzBp0JlJXa8V8dhf1u3T
hOxeVIHw2hvmZpTTiS8m/Q1mVQQuFmPwq73PhPcGRSYqa3yyF+egBJBTWkMAifPFxG3nhLB3/6ji
EBwQolh9jK78tH8dH1SAF2Pw5ndHaUDsoHDaBb5ZC62Ewfgt/PZTKs9h4EtUoHwJCtzTo07PQfzk
9njr8L6oss17XnBDl6PeMKLYdViTXoHjK21FtGb6CF2m88d0ec3Hbmvh65P9jSLkC60qRFZo3dKY
Gtg4ZoZ41dqJCSeZvs6we8x1dwFWcADNx79Vd58DREnngMhU9laBBIbMf2aSYQu/PpOOSlthxh6j
2QCbckl8ymf9WyDDeNYzG+41I5nXzGY63qWo0t7ragTzj9N8epSCzLIOdkntO9zwpXmde6mEm0rY
Y2Go6AohBtJJ/JoyD8hrUeutNTxjhLnxKiAA1ovapL4H3dG7XNYy7gWx3NT5xy4TTRjtXgGUsecO
y49+7/QbAlopeJ4qQrezlXb+JwPNra+LETL6yySjff2gBXFOf6Sskrc3ertFWavXsdN20ineiNnZ
RON40HufOAZZA9z5GfjP3HXpcxvq6rWZJT4ionfK8dVlAE7Zonqs70oJ0wEDIyQKAxizTST5mDpM
5nJw6lgU+ScZE+C/HWDxhzl0MMFa00UfhUg+xKQixEqdlr12oxyVkZ/+7y+IdT+QIPCwRMs5OvKR
gMvk9HtmXalKrOuC31O6+2xzYU5tgPvlq2toMZ2UFK5Tm/nF/zdgB2qlOi7rVm59exVndHzXzJ/O
m1x/EitH8NalTe6Bn+Rdq+Sz9Od143sGX6sZY/R8LhCp6QXS7bsu4iYO7yXTDwG9aG3M16/onPrF
Hw1z5KoMFiHpQHIrJD0tM7BSUPHQKDcPpudmzVHOLeiMRc03jxVNji6pW3AzeyCkjKLe8H3N9rjV
Ir8Rm6McX3Csq7hmRQIs8ZqxEF1mq1s5r5yr3OLx69o9ZG8ZFcbroQe+dTzZPSB189Si6P9MYMvn
zvA+diac7HMiUnjZgF3kPxk+o8Hw9D6leZksyoNjkBU7bYohUkOFBP358JpO+E9Hg9dUy7zEU1qi
0u5NClGYhk5aLSX868YQy5jwudMNB9LBC3kFSRGbL/MQhVXYvNNBg2lClByhP7zC7PPbfZ6HqSZw
SmrFRTWbD9Ek/+dPmL1Ci2/nV05uWMlyqOo1MJHu0qyhY9lvFhVsNc9ahssxo4/eaomYvIHUCJbi
J9Mok7Xrw9URDyC+BctoVYtn/jbnhhhgD1MtfzFOMjwZgMqJT9w7QLxC0trMouUh8lbDfSQLuykt
BvPXXZcBMIEccqvX5ecE67+EVdPbmw5CDuJGa7YA+OiA7tfpPN2TT7+AZxKFDMX0TPPJfmJW/ODB
xccJNcvw+CYmwQcPGqp+l763AskpimwhgbdBoy1mc/9TtI5J61aJtCDUB//VISxbDEMO8XccFasB
8V6lttILoAEPyLZZagqKJB52tEOfJIfQMiVxe8pz9++hvebE9kO3NTO77gr0OI2PFhqBZrMItp/x
QB+2XTyGD1APzqoQmz55rnnTW9mCNzfmpkrwd57d3C2tEjlYOw1rOxKmFUM8+8Sb714xwovVSbyE
ZIzg1MXHu7DFgF0kLolYH3sZQt2tHILad28W03rkoOmAzzakxTQOJzGIgCJ509ZMizGnJwCwm1Fs
X2Uk5/dK3ISt87TX6g9e5c6K5OGWJj6U5Pjgclb5cCvX/xxj5sQMbpyMXBM5aDjGTZmpin8vuxU0
VqBHQDFJ9sjm0yWXvl8eH2JXsbrM4w9qs2O6tBq5bA579KFVIvBw4PvJ8tOU4LUoGuszGon9yr+1
1B946aRxrDHuDLnQujz0sd9DVnZ5Y371LWWuKw1yKW6RLl+cwID11NjnY7sXvvCxHJmIvNXFs2i1
5HB13NS/YkTHLU8Xdi0KRK6EDFpa5LrsghCMraatuBs5JlB+LzhULklj2bSUuV5mZwuLCfQ5mvqa
k9RUYpdEAEZ7Yz6j+qMXkdUcOcOuOtCN2mFTggNZpGw5GApd2EkgAp+CNTnGAWBc+U8Go9tQaagF
LXN0ZNpYOs0eGKf/oxwLZ/TgRzpRiEEXyRLT9chdooLDIW0XGl5sNgkMTyOFTkDhnd/GnLdK6baF
W1guLjqeJHKpxichKe/2MacvIuelfXetjT3fyYf+xv6vZbUrDeB3UZb+57PNs7ErSIHSIEcyL27E
CkG8DeaR4PvcI3tG19+RJToScJH4e2EI8hHxARD5+gfe8Rs7VpJLV0VdqTpCyIWE6YWf9fNMkyeP
JBW9g+8hN8hjLOeMvsAoXQFeaSYYQ+GaUyNIAamgoLIAoe91N1HTcG0Jbl264qGjXLZxG/i6OXUv
7/WM7ir5COA7ihfXTL0BcfGOJ35tzIYKl5j50d2t+0+b3pO924kJvX/00czNGNWp4nFvtfHh9IGf
eO6xc4XObtCRDI8QLANdtPAxdIxgrJ9EORn+IGJW1GSoDXps5YxdpDX0CL42Xfe3yEQmToIhWled
GtX+FC4LvtXUIrbQY+rAZnxqdSpnXI7KCxniH2MnkGQ+N7gzE+fHIJImT7YIO31sHVkMxAZ+Wspd
3tIxfmk4vvY14STYFc8ZgYTBm18qnWBS5eKV19kRNcwToN9GZ/mlaSKOJ20bHhqJsGceREF2phg6
/Lif5Mo0Jiaik/nGPr7k0p9t13r0d6kJksqNV2wqnOYWZLNlkv4buEPN1EG6DR7HGCaqYJUMP4/Y
w8SjJBl0bq5SUCRdcUc7mNkdc+lQkHsgZm1XCaHZkC/Dyc57t4ot375Aubkpocni9O0v05j4XBKR
XR/nmv3TDqkRSdU61lyY4rxLDg6xZUbonKQKw19jz348V31HF20n3ddiH3Do7u8HAytiDgZPYXsa
l/Kw5UgADMyyW/bd2q6AotXmsI15uA/QI1+diFpHgCClPmXCbiRlpf6ITcVB2opEy7eLt2s0/xnZ
tXVXCWWo3TZJw5JAYrPZQp4dwY4LG0BnpIf7ZTtvxEZuAhwCOK+WGx5KFx9JYFsFGoyMi6v8aGq7
/RKrWHnjDgrLGysIb7wNjvGRNNzEs0pSF5vxj4GShTB4zL/WdXWKX5igM5bfC7eGlhu2qGkoyjjf
rUshN53o6cdj2QxqHrVrGPoMQlnhRYse8hhzGdzg6hP4EXr9n3rgHkThQTuTFOTGoIsb6F0uUruB
ZCA7GhREzlSe46H4iNKr8JpWqQF0wV0n4jKEmNPaD+4lnTToFqPMsesE1S4tHEaYQMwj/GwHUiEU
T8V3MqzDo86Sx1e674bZebIihS/0jqMT6n8L9OstTcGI1UCTya0pYWtngVeTUI6sri9xLpXTlGIL
au6IdDE7Go4gLz1Vy9v4Sp3zbxVfLCvsMoT8VQitRB3XWxF5hmmCVE7Ec+pi/yAHBPFmqCJTo+U+
tf09+Wh8dzkJNkQ6x0tGWpKOna6mPFA/Hiefw6Nsf3i/Sk2/jRPs4Slxi1Cu+cqG4Ie0FJdbHTJu
6XQuOeXux+eQS7Xr3v0QFYUjhcUbQPn4ykvweEUbjpavjvMHc66OGWlhl17C4jUMiP1cdoOSbsba
dXnA8DejI0D4CeEndYR7ug8gv8Iu5THTsNbP2YiGLefpfaNamNQRd46kabYww96RPebjAXACUNs8
I0j8hBy3k/NyeMWqmiLhCOenaXALjXyT4JMFb0Y2GEfwk8EAMtmsotS0rekqyiqimQPY30phMyz8
6P0YHTQLTssZqpBSVP8XEjoBn3A1dTi3crSFC7qr8zJ4Rx5iUKMQpa+cpjp4u42XUV6tJsVJvVPf
84g70BR3JgiwQVieKATXxGmjouDV+/X021Vb6z7Ftp+WlwQc/8Vinfa6c9nxJ9TE662sopBpSqwy
GkFDC+jGBk7ji3juQgBe3uBl1Ulx9UdZ45GjcfKfvvIpsx1pMuwr3NBP1xCyxhBJD2pAjgWL8sAA
6jM9364kppz7XtMyxgJ+aMGm7ilfzSYU5vDI+fPMEVyulMTufE6fJuq3OF77WmrU+Xhp/AB9f5tE
bZkwYarB+GFv4xhZewpp0l10T7ob5lG9Ko9Nl+Eni6D2UDe97aK1DEj/+yLvCBxV0qkL8hN7EhnK
85J2bddpYW8EyTjgcVJ6roZszxzVp2C8fa2piKDXXmFMWh7oQMmqKdQGAdOFiWoFkNT6jUQBp5ZU
gjNXUll6zV4dkWaZ779MQ172yvG2npG45/Bk15CcA4Bo3sMa+XYpNA2fxKlHETyEaO4jaNvRjFJK
URU3UUIWefov/2uJeJI4HC5+p0I4oCmPwCSq3Tgji0TYv/46IT8UCIgsKnwXz2ptxiTH3thY534X
qv0Dd0vMOuXtD5kNWqoAwQzIxNMeS+5RKRCyDolVGoNCyxCZPETVWon2ScId28Z7Wc2QRgXKZsqh
tVAfduRWClIKzWrhyb2oHL9subg44uIXdadJjxrRNQLleqznpqtxJFrPfvtPSXK9XbhYI5giqvKG
0Fh/KvcTtr1bOIp2t7Xtw4xmoRWiB2tqtRWg9VBgOu5J81UPgp4UFUqWNASN654GE5T04zG+8XX2
L+TJLwiJ8qCgMFZgE729nWtV3xd5PKCLFBgQtWKSCMy/ioHikoCpzIZOHj97rc3a4E3xN1iWlGc+
fYj7QRVBQj3uf+k0stqj0KGHJHiVC9jJ+eRoZYFF/EB96bKmXAKe40PLoqfBq1CuBvQ9cjFVsdFB
l0869C/regUr6jXLXdBoOVcWNRgIlXUvwesf2Z8IEe+qbsrKoG3PSChumn83veZb+huoZIn9mmL8
wozBaxaeT6DL1rj/Yg76F62efAv3ete4mGq6bJSSbnrhC2b2FEf2txgqLs0gwyK6CobrtJrRtiLB
Wkr2ZjbGQZdhsaOEHWm+pehSsxIhvNhYrusD0TA1GvTGNjIQwHmjCPUZfwPXdjllg/CYZ/xu6OUN
wo9xaVVaLOMtgZ771nxnt8oO6+vapSiaroE/jaDtz7yVantNpCnOtJ4jQmHXJmHQIAfg2KKI/mAW
pC1ISBTf8Rhd/Z6tmDUHlrXEjzLx6JhyzpL8CQK39x6BBhaQ7uYjZ364pjidF5n8cG/LukKCtWDr
62iQmmAw/bnyI5RardQupB8tYkjoFAikoUZxtqUGtSJmZDsGWcGFeN1E5J2H7VQJgCxksaXxsXbX
TbgfyrIR3UZ9D12HxKIS0jhe1AUJikDvsFYQm113YZJY2ts0kM0FlLlOt8xAoiOWFBJejUxZqsRy
i2aiuyGOu9v6BDXb0APZXc0sn0SDHefidP/tBEgoWE0rSWJsy4oetPQLPEq9IQUlgXYbvjCb5DBk
j+GF4NjmEHF7oghXiRLYAuMaPN4+5VOdgi/0NRBVviMDnk2jCJOQ6GDmkxb5SBZ4bqSv6GR4a6Sc
yQqJnPZW8EgVoxQN2v2gRznzJMiKLsX4x6qjN1HiCHZsMA3/SN7CNamNp1CjNncmKQiLgVNMaT6j
KpPAQCsCPPpCgf2Vm/lO2RIXBFE1YdVNOT7+F0XB6+fu87AMC1Z0iUFB79+AxRuXEf5j11p0Twim
7UwxIGzgleYjGoLOvF6Dj5DNuZyLV1q0nCNz/DkZLyGWw6hHNu2VkxxhA+U9cmHp5UrgrUOD9Sd1
k9mqCjxoyH65G8KSA9W4rCsUsE0nIqt1jYAYo4+vLG2Xmhvd3hhZbLlbQY0qBB6FrSX2JS8LLtD3
cuXL3EJufXq6PO1G/bHhPCPM6X3a7BZr5O+p1BT27FqhllTc5f8NHmUkM30yjV5KuDg8QiR5Wz6R
Gz3WTGxpFevI1Ewl5WMud2AtIHI6IneidzheP0hZI3uB9E3KlxYBR/SY3uN+oZ6xvMqkm9c1ctj7
HUGNYFqhPrRTUqSqtkuNvvlGygkpOgCXQn95q19SKqIdecAc+p0RpSH0i10hg7CyWOheQisC7z2W
Waec9dXZPdkeJgb42YqzX7orL4y+5SF9+/fUtbnMTXRhm8nJl9K/kHgeY1krehXb1TBGBsaitXeJ
Zs1Vugl9phNkr9dOPxNOcQqUdgk8fZUKNNtZrCtv0W/6O7OuARyn00WwThndPV7xEBlg/dmO9MK6
7PLJcZGqaTsxcJeibksj3ve4LXLaRGbPO0X7d31Ti8d09wYJU3d93bnjzsqMR34Q+aV7uJjK5fMi
Kpp4i3KFjYqmwdAcM8PMgScHfkhHbA/z2l2sKsicxE72Lg2NLhRit/zRieM5UsM1xE27dewuP+lN
3Nli1tYIRRZTjMjKa/zSk5MGG3JS51vjNZNRvtt2TeVVqrG6hpu0WXqdmwD2k8MHt4+Tt8envQnG
/zPVyC1h/Xhj3rQdasMdXOFmQisUywQmIz+RG2HMow3qt37LMQ4QSMioQmSbesvbFxT0RHqt26Gh
SUtMp5u1DXUcYKC3SdCTJe9SlZefOXlOZnaLeI1dXru9Pt+QHsx0JcYiiTnI109tuSpXvTq2Qs1+
fGhyhSEkdFRtpwdCIuGHgvQDU5C59P7h6+lgV3WUqyP/KC+Obj2bi0ckx4mUTcEm3cINiD4vQNuy
lDUD1cc4T9KDQRIIz0bJmFxPT+RRUkcvWsBTwmDl3QL0EDqAjkXqHjhIfh6Z1m2dgIfQvLHGaYY2
ZzjLvS87jo3nIJ3Rn2iZ9LO2B2oq5jc3NRcR/QmUzzMKiaw01Gdg/hDjDNvuEKm44Rs/9ZMr/AcN
VS2Q0iEWiG6HaJ7+4BLBXiBoGTqxv8NlGpb7mCH45nq6MNRTUmZG2ZNodeEALVJUZ+pLjC6jJsk6
MMBbSgdJ3p30gJD587ASwQIY6Nj5el0eyvJrR8kR97WYatfEyD6Bw9yESk0UvRlNUjckOMK6I1Kr
9QEcZmv5bOpXljp7yIkygiOQ3LkONQ2JMofAvHyt1gYaM+zHBriQzPdSS+RcYgJUJ6LpZcr9PQtV
/YbBYvF5VgwnfesiXVjNmDAp+v2oB6EXbpvrjoVaHcll3p4p3RtRIZlJXi8lzZtsYIVPYzhnVPAB
afM4nSguFvZBQN9XdZ2/bV7BXeobXzMGFzeUZzCFRd+8gle2oV4rbjQKG4GrLd4g8F56IbuHRa8n
KytdnrfOPfr8GDf087sdkDk472tVqT6171lasFZW4O/V74dgogSXJl5m7fL7f5l68iwEpi1kE8An
B1sbP6SBJOceSBYrUj8hyqy9CWY32kLznJwRtS6uaCJeAkaGCKAPxRFYLdaON1agnvfxZdPw0Vsp
oA1cbcn3VIe9jV26pK/g5ZaJPo5Y7pKBSz/1i9SjwpXpumyycSPRlTTNn+N6lByV46NPowc9kQW5
KZCrH1y2mgV1P9J1cSsB4N5DzvmMfZ7iK2Slts8GEw87Aa5r/Uw2AjImzt1KqKG08PyfvGZyIDh8
IUY4CqcCeCPqFdjmco7++aK7pdOHAhsMNnNqtEcO8MqfR1kDVoMQDYSUw2U7vul5f8Kiupr8InjP
YGDf5TeVqxCeTk0+bZxLPQbrzEvLr6jxDH3V163+G3iuXubCv/CWVbosJZI7PqNIByQc+7mHoDVA
BHKkj50fnbYGoFIGmKnxj9JTqlWABvjWzESNd9RqUL9DD9yTnKLcOUK9Yy43dbI40ERiEAIm4ZkZ
ri98bbO2nzqC4yhzdVKDy1knO0XAv/6umF4pASV7KraikSF0REoqNAgmubhfdgK8TgcZBmbRMFIA
81Gu0PImLKnrTnsGZBD9SiZasJ187g6k2b5AkB7Cuo9M6oU7LqgC2Hk7lXZM4RQNc+bS9DA1MW93
5EmqCXA1YeWYFhdaq7u35nbKdLmnHlJB+rRzPVmfskMyDdLz3D2tyHKF7QDm+KaRz4H/aAfXjvxj
jycDXIo2X+FYsKL7U55CNBCiCrj2nyBhnYZH4gaLW3ryeN1VMVLsGpbSeJIuc3o7BUgPlknUG9Iz
fSKtwz+EPP09FAdfzasu9Ib8u2cmfjYqcS7Rlp6xiLxVTD5Rzt8ydeO0oa5gWhgpiIORXRxtCik2
oBirhwbCb1ARQpBjG/rGt5SOsqGId2FEWQdzAI+8au83Uhn0crtSApMwJrodPeGxDAZefrQiIH/4
RHIFiHmDLEZjeMWG4qzCKq4tvwDDLFoDpzA3UHs9bFWS9UqW/SHXRqBvfLDw9P96tZwV+tYfdaL1
WTCy8/rtAwDBJcsOkl3HFR0ReHX/KY/P+fSRhm9oAp5eum9GVsTE4dSYXFxxoXkcuyLtEBqKrqbz
ijNTLxu8OYHThxfR4irK2SQso0DD3qu9kjTeTAeV8jJ2CkEB1saAdTy9JGZFFdMnqfmpmcns+v0/
DQ4ii3l1y5gk7Bu4RiyMf++kO6rG0mzvUMreiIhp7k+TYf2NqPk2QF4bsRapSm4TVWkJABlgICUt
GOYr4OnT2EOpYpJ8F5JdqQRcXSxwixcWmKtWRj8hOFDzAl4HqHMOdb3mwQUEhWu/5c/1Q7KMyMZZ
2diUqg29u7emzZt3vZ+2WYdRuAawyiXsLro75/9BMhX11ZyBBFscb/PhIUfa8nQfg8UeP76XLrpg
rI92Sdps1OSk8vweZ9A+9NuX8cb524VGdbGqh241Xw7aqAbNZ0qkRscG8GV2DkON+0W45stSqklW
qMWCDlMgvjQB6G/iKOyUnDyj/ijterMK6C7tDnFPB6wEibp7yJmch7vx0VE574vatanI6SC6i1Lw
JPVFvNhAwjWvMzw9MG9hsnrj2KcDGKTE/pnLyBgFGeFzJ5yZdg0mPyIYDX7cw8Zf9UEhPLLbyQAv
gsuubIomi4u9HKgnO1mN6UR86rlE+wd+Nk/VEyVFF1J1qhNKMijZbzjeWrKUpQ2sKq9Nbg6QtOOT
UYFmlIaSTbCfSJJybli/7SAIb3h0lMSv05NbiMx1GCCLp/JIHmjCcjR0mHJW06wUZd7UdEq2Bfsz
s6hJxXt4K56eJuoClv6lXWUcn8kLp5JdkbUX/NAtYG1hMOb5pLC3t/kwq9MOHKlTeM4OWaMJrOF0
bqfgF7UXwBA2rJGCK1ZiFAPUioUehcrm9XgIa2KJTXZ135ZaFGtYIbX+1JpF0r4q1f/v7fhGUOuE
8xYeb388cJFDLMk34aN472h++6F6Co7qW8aDg1vEy47hmKVh78ZG04nlcSeoyFIf0m/mCLgNXYDF
/OdYfnNmT1IHSHbumQZuI8Je4ZBjgJM0IoyT8dhcBRbLJLDpjxo6yALmca+CxWhcmhMWdebi4o8K
8EOv9pYKFMumOxQn1qZVq//c7jNZNVKuxVS0ErQiahkWOiECVtktlA5YhAMuaSXdvUFMC+XWH2RD
X8CdpgWk6/Zl0vxZr7lwwGvuaNRz26ZFlOa5VqhfLUnJ3m+nRi/8PaR4POX/gqI20Vl5KHCWCJtP
kFLSEtUWPaBrETJ0DAWqATPWx76YpaNHZrJpYFi9Ckl0fdiQI/O3azozPrfWpJwKPSgI9+TZvdKI
IVXgBxjY219WxvUl+Y4N5Vbuwb7yRNFHs9vjGjl1GueLcDpfbP2RClMQ0mF39umtXPH43vZlM3ZV
FsJEVaNH8DLBuf/H1/W0IIWbN2FNwwnFU029UmTswWqfc8160x1OdEeLfT6J6Jjy2wiwqPrfi/nO
lfUMKti9+vA5UcohtZ2stQBdFfmWpV/T4hf/sQS1/QD3/1MUQ3UTVd/jli2UeuRi6Qvgh7If7tw8
qA7sGRbyVCG7PEpy6OHzf9PHDEF8N1baV1xPxb4jVgWuaCnN7bqhF/Fy1+xIBptTSQ08fMGBOX48
JLSUbORkFDX88ut1D8sNxyywZPl6ObhVaTUeaWmvyeUeeRp45HOQTcyJ6K8/ChQFM2nTlBSR9Oqk
Fu+NrnKFPo53HNtY2MqnvMJ+g5t/xgwdPn+K3sfxi2HonIpXJEFtz2vs2hqetC8SplIPRWhNQlWv
eHF614WypAbY3c+VCzYweYy6EAdWv1gil5oORS/9qwmhH52pkI5NFSoj0Afy82nXseZeoYgaCP8A
fWhcHdIRZRbK0JW/+NhSBQX7FLn1eSjQ5wFXWfhPWI9cG+dib41E/+zw2r25h7zYFPqtTd/Zi7bj
zAxvOR+7YRmBME9w65PN9kmsqheSTxBoQdExdGWKIQE1Msw+YLwSYuGVFnvGJkzeoJi6l1La75Tv
xZ/zZrNiI1vQhNlh6zizrNQbmTfu1FG/6Br8o7Q9NIaIgNW8pmbupoTezE5pnDnWD4xiXPgDHUlj
FyOQlgHRjbBs6FZWi8Yy9pdf9aCRBP/iyZ7uQEd51PjgK9tzYK7Blsc0dG6CTaJDiBunEeNcDtQi
NHhGHxo7h8Izq5LJWMW6TFJiXEut8VwqnsZ3yWta2QfKeFcrXdTjbtFiASoR8QQXeeNj84L5exrE
NCjThHaB+E0pbV6Oyo6NzySGKDB3uxYXa8qATs/w/6G4o1H3DTTGAVqnfJRDiWZOJWtmOxRG3bUh
Ju+nlK5hKO59z14qz1QsE5QbcNB8uFRAij++OzzbNanWTC1OSQc6Fs1LuklCOQSiq7CzeaEE/8wf
d1/baCtJ9Kh2pv+UtQYfLobsk/ArXtGacjRdzA7Y7UZvDL9bosT4FS/vZPIlBJ1AxpTpJ3Mb+FB6
GXzMFIA5dpEu3LiS1CaWqC69ITLVkyQ1b1R9Jx8t0wPDOFngH8N69NnjT08Cn6SJwTPnuEsU1VYk
CNV3NDvzqWhvj2F30IiENkVyvQfGUE1OuRMBSSR7QBsLXVincQwdKlY8z0gj2UVxhXhXXOchnxPL
e2P8OVSEJY1T2HHQOCpFpwdJFv+hT5amlVi7KO86f8gnARU32o4TNxdbxqbF5b4/C/XBDFJhXp8n
Mvu309oKPDOHuDIMs0PNge0G3TJX+Egj6Tazkz1sxyXWP+uGFAC++56p4gK7vg/8Ar+VXM4qoE3F
KGtv4cBNIEmrad/mf0KVG7UAx5Rki2gBFdJeMssRVvtamwHtEAf3zhPJvy5mW7PgZ/EXcBYytpyy
NqW+Chcp/PWJLzr7xvyQP7Mb2cQCaIvRXMqt/VVZqkPWBwXlw2qTuKJJco9IS+z4Q7eMiVrpNusO
SPGrK9eXpfBhaCqgIHQumgs+Puqlz0WXouC+HSL6KRs3BMjSeqTWpa6PBtgcTPtFTIWp3tgEGn+2
QZFPd/l729wEyHyY0CZvDKal/Qf+n0uD0FxorLpRL60Ym4b6eg7W0HMuSQr1R9INK49/PaCf/HXI
I+ng8NShDXIPpW750XDNMdWEZXY0SDyAIoGTOMvAQNsimO/G+JCK7OEVcI14VG//9QcF//ZmtJhK
8pBNFpODIdHONP6ydWMCyHJ9op5doil19qNzD4AFVOiuLu+AoMbHdsfOi4ULaeijmr/W1bLiGYsF
uwr/BiH3l/TZKETk3BF4RemUpSaNuu8+xGzrQIpahUC85guHgrQTxRamCqWwlTuuJuba4ibS8MPp
3vw0fRXKJJCgcZ+Pu8RhUvssqMmFawHR2M5tLARDMvmx18w2tkVZNrOdRJO/mymVtlQw5ioRI+R1
/owBTdKUbgVl4WlKE5+Zz3uk13gqjyi2BdWsIJA9VZYYE0K2EDtzNMP5Fla5U3/VHVGU3YkkfRNz
anpdhkb+Vjh7FzjiGob+DmT/URfGkA6ev/PVM4ejEohRS56MX6QfL5eGfSr4sck8LjR1efSyeo6O
S18huTwhRbez2hARjAlt0/WkTJ30/6STVUI1qtxi/zhu26w8uv5fF1yLkXrPdBAWvt7o54gOvQVw
3OxCHCfsTuf7kY3tck9Ou9bzieY+oFan1Ykl0aZn5Sh4PoF5JSpWXxmBcLBwHjBhBsTaSFa3/cNx
VQHIAzuC36TqB3FV4JiNR2orKL35Pw4FzAp+I65WPbSuxzgmIl7jlX0KWhqGCKU/vtX9Axov4pM8
juZgJWTIg0iP4X5vXXeFcwYM9fqZiNKZpLtxHwUcgyZL2/FnS8InxbcZ0ZAMP/EZJwYDFReoRs+V
txiD8AtjWxbfRV5nLSon4lbKVcOY+o35eUmM327R2SbQtTaJCRyPM07BoqWg1LudCadLA7Y5JDDu
8pTSgZ3WrlviKgef3G+Xy/bznxRdCNq7dXaFl/zwKf+G1VouPm0OQnsA5/RsZqAp4Flshr/Tfb3V
TeJhlbmrNsMUo6ImcKy1IDQwr48YwrRuX0Fa8Ie/jm62duLnp+nKYxBTpZFCSCnoYYjn8szq7Juk
guSADQTrIeYmgv0AueDZZ64NbLQnO7mgNE3JP43aEUJyzXfpp5ybyVwMe1QYKvIGanJAWGLITxDs
3Iwbs4XIByM85+FqswlARwk4F1oSQ7n6vjdDtBBTwa9Qar5sTiQWRAffvLZRi9X0JPRjXz9Ig7/0
8tCP+wUO66bJCvt59kYK45ZS3GVfmyxVp0T2qvCuJIPULQynBMCRcX5b+57q4IzWM9/zRijvf90D
lOHy3XLmCXGeeGDotv15hB+5Ketioih/7N06gpJM/lsk9bnhcR/PtuqrkTAhwSVpOzDUWQ2k4dkK
wHWTrJC0iUg0iO7f3MnBofiD5uX1gllO+XOZuQOcnNXy9sKSrNTmQ+QD0GzhVeXRY2VfReCXMqwC
K1tILBS3bdHm86TLRtDStyrfWAjsWAs5qaDi+rjAiX+LKTApKaaXm1h4uy7oPClnQhgROo3A8fiO
RSqzWdzLj/8UGJSoROO7s50WMkjzLCuXRFtLWUXH1QPZ7na68rnsuNkoZFnxq8/0k78IX7bMDQ1d
KZrwKUK4EGuOPe+iB6HMRXS+fuW/VKGVZR1UJZVYQxFX9x08fw9w79DqAu1SvbbavX0j3bWxhzpl
xGGpPkhCrDoZJSWHpMHZ+5RmlUPnVPy5bmB+JREr1mLR1LWIHBAoiBoZ9aWtoUJiPWa8MEGF9GA9
4BWIJmzZc4gQW2Dx18NBR7XI4l4jlGwnmDbxUcL32AwdmCQZexlgxKhXW+btHBEVykezCQAKwUBW
oUp9EKbuHgtgQjNQAdaYQA7jurJ2vwqbGYNvVvR4ITjEmquMJkcS1oyV07Lch3YVyJ4jXxess3b2
MjrsYqCHdn8mwnyC3Tnc38NiOV0advvHT84WCbYBKs16oIAk4keqr3l7vnEN/eDDLfbSMGOjjdsM
WEdh/TU3o9RjJRcZ1bybEM5nnZRdcQjYoeK0m4HWQ8K0Zj9bv6kGaXsG3ydU3WbH1ZtC7FbVQthV
kA2t6VFa3MUVoO4OBvm+BKBH+qQTS6Fcx3WtZMVvp+s7/pcDBN6O5vA8vQVJzsNlbLn/640Idwma
JsvyihwA8nD4CZHa5XfbN5wMRb2oHlUv1mXKSYNhMQvBThSGX78Ag/bTWX8rreGkONUeDY42vKfh
5N2ZmMDefnNGTDLwfANpJ2wupM3VtG4WVjbF0vbXhu4ADv2fk/WXEyOcjvIvuUrVZH7rB9BLcZhR
rNYJ9XXu/mglLX5CfgWLx9Xj7LqWd4NERTT+KaTNzOgRMRoIGTH3fPlqg/MrNt6g0foEtmGQu8Os
4yij7pCJWBGrWwrl+CAcHAmv1Mg1WzLup0wfHbWLdH1IkybbOPzIkGFH7gNK3Sg4J3z+EIDph+or
Ai/VXiHUz1YAEwPcW4Z6xnuWyHZ6P7/wCNIzidPB2CU7obKRF7B4dA+zlLe8ruBBbdW3ufVOkSW+
uqGI1AamSf0IVruSgYVw1fXVc4jtrgF0k8A8YJdC/RSAlCoGyBjrcy9zm0BxUCYJAkvfA9RN4Txz
BcYzrEoY1JkWA0DsY2Vc6eDv6C9aWED90lg7QWcVeN5M6B8JyTqEB4gmK9jKjvXMEVnej+AGSgLm
pZoJ1czFewNQFLCdYZ1XO1hIyNME8UtDn1dXflXfSJL77cGCtzgXpzXTsnimSAGZoeQyzzQwhKL/
rAQVms9fDT2TevzPr2AEg71/RAPBq+Vk9FUyioW9Qtar6H30Jp7TbPxVSaOoGfq2LbfuisPcNaTN
xhfACebLA3v9WZWJ2GgyZz76u8WKpagG9W63nkSKyDxmOJjqMZlM5T4lzIY4OBFL0OcPPbTzmV49
6VpHUA2+xi37okZm6ktNKIw87eVvA5bpzRB7shEUcK++i8CyZE78EYRYRQ+JziYSGN2+4E6WvvRV
3o6V05fLZhwQVaTKUb+kZ7I/EjXkZv36IIj8s75aWpVh+UUc3u2ZrLetMqI0F1wm3b1VEhAkk0NS
MYcjnRgOACunc+yxYWWT4nGoPrF2yIvzg0UrdN+Rv0Xf5g6zyN+OAGJuC1OH/ZsRTL0eMhYrfKY8
P11nsR/pY2sbbiIXQiB7DLcxK4574CYzsjgzmc8iH+hlV+dW4gUAYq1S79uUsLxBhfVfry3oDhCu
IdlD6psu0sRm3VE1pMimfapIVjwGVh+4M882UhctttGVYcXHlvt96yPcdMglf+r7uQHTudxZB4Pq
iaPBeBWL1aOmeEvihkngWrW26FbmLZKlNj0El5S/hjs0REj74VryZXCuenBIlOK1P/lUisWvVFnB
aNB7iYgDQBH+gcQWNgzcUh4BzsOw6eyDrGdapJpVD73WI+F+XECnMb77b4hme26Eb+1qn1I3BIco
QUfS1j17Jf0U4w7B4dI2mYJ2JyAvtv+A8XwNXKCgaOiAE/DneFdbYvPcl/x6nGZp7PpmvXveqsTl
7fz+NZ0/N//8iJjSC+7kun9H1m7lAAEGZ6IU08Su7HreuFQm/zGJHxCNrOYLSGhhWE7RZO7EYEym
lMAL+TN1WfOEWoUhdsk23LbAQmW0EzAVoi3BmUeTosb1P1mf9xRiZNlTdzLXjnNud6wpHJ6r42yE
RRGM7/sioEIMq9jsioOWwMDpmJ4hlHFoEYjOLtTIL6+8tRn2IVQupzVR+BVaad8Ojvw1gFvvVHAE
9z46wuJyG6Uiao6MXzJ9XkpGyd4O7sjL0ZvjXsbP3s2fCtso0tvRSKvz4/2RWDtOTMna0jQkT6r3
6RcGZCrUX1PUMgYIYQEIJqAGfdMBjUqhBdAE7Y9TQoLhnIHAgMxiCCR679Q7CgG8upGaolN5oJF+
hLBU/KIi/TsUqT7AAPhI+DjLSEgkrcAk+kVVfMgmW8KPKHtOmX2GxlG+EpqZsYGc56NsAHDxmU7y
H0uzP9xNyQgz5U6k3HwPFUIUZbB/HinBidDnx8SdgK6ypoiiXh1em16JgMPlyfk5/N9y8k81q4sB
skICctC6JsNRkFTayPwpaHKeSzXaGi+fp0e4+XXxPzm9op4iaKmsonaebQkzW4bNDzQT6wAMqsd+
kGF3Ng3EhOnD1uAIKjeEktqhEgyuH7IhzHMaqfCYV+b2NPOX6e3RSK3z4B7K780bNnsYq0pnGQXf
cV6nhlvUPljMJqrvlUMwpuLJd5J/VydREteT4VVipB0whArDH5GabggF/0yBxPJ4NIAJaBFhNjjx
05q8igKuPz+TIjEtVJFZMU1Qp5veDeqmcMuQsOsR43H2Wo7CVwFc444UKTGWLoW28OKrDCPewe1p
9xuZli9SaD85M1LHnMRlYwkxPgxB4OGKuHgqOYJmqTMFPvvNtQIeFh8u9eHaVzd6WUJ6ZkbBSvh6
hlqty1HIkniLGZdsvkvlNhA5twQc7Ux/lS3ly8oTAwCWhFmAq/zuQMsNmJ2iQXKxK2vlkcIngFB7
JOuhDL0n+ZusfuZvI0Xc0F/+DTUkvKYluVy/IW6V7MFD718XvdZoLnX2/QxrG6DhqV49XWmcNFPw
xmFqT5WBtALVIv/Fo2TlkxF4bkmtSsDMRi5aoKFi7Mo74wOVF2L7Yh8mkHmoLdhhOskmKM1pZz2o
OTqRJGWAq7v5qxP5flrSA5J7ajcg2/IKT3mxCKhpmmG6JugVinQdUU5dOonWZ26FlITrlOJDrpqy
/GAPG6xY9sHhPZyqeVEhw2LdoIf37qTfENGbNofXQJhJ3MpOvem4d3jIsExWmn19H93Ycsw3ORhA
QF1DIfAfEYZarI3lypLXIHbRpFoQsD5pUsXt0YSAVHQx5livAzuCdoZDWWKgIrjRiSzqbUXWBl6P
6dJYg2ukPPuqAzRwQ8cvoQ7ZiMzftrRZjDIRn27T/hGs7v6P7UecRMjwdmVg8qfBeGckyMZ+qSQ1
vYDmXCcK9c1ximryVFbovabalJyVXmNyuIHUBymTF92f2hAJLoZK6p0fJR4yQbOZufRJ6CF+rmmC
eRMeuCKWYS/+pocYDDcUFmEVRpik3lUyvU2eYxnlBnY/wfDMni/M9egxHbcaE9zLEmMnqliu8O6j
/LIZk5OMaYCFMGxWFq7XPSjMlO6oUKzBoXpY6bAwnEyb4xkh/aUuFpOJlXfuMxQEthdwMEQUB5Ix
yLnnHEhoQQEcXQ+HLGMEdiSaq4ydpHkw0kH6VDFBCOOBrl1GcZIiGwzASOxb/8IYCfqPb7KwSAVs
8hjpq5MhqvyItW3UXk2Q7D0oIOHRCvymM9QaZAjy/w1CzXUxAiBe7aZkturivOPdiBXoQmsVzl2u
VaEnBV/EB1vz+jhXZN+JGo8ByjA73N9+LpG3pvCvbp98UFq1kKn5sYeQqC/ahutCMwmjXfVFexAc
HAOgIkUtQuFAbmx3/6EdqplrcfwHxlYOr1hKfZdlu88pIJsK6ZbIsS3cArciyUq2HhtAgYgVgKWo
pRHwvYUuGgeDr+2fNNVC4a6mrB8WnAIpsSIh6wqSDGFC3/TvA+zabJ4dEXCyT5T9evBx33f3RNMM
WDCNaF0zqmun4ztmIynOxkgPJOjyhmvrzzycdGROevAKNp7ZT+hynkOnNu9lkbvCIw6c07wEDOHc
lYJXttRBzJgjg6LCrQo/1BTaZ6UZCTcEq9SqUBMVechOczTXA8/2+CGY8nGo7cMt31+KZxhQ5nV0
9hV/zCgAk7vEtDUl9oSkz/DOOSdVvf9nn444/qbbNnGS4gLrYXp/jNFfkoVUf0l0rpMMdg58ubpQ
78Q8moadpIpKIGOdxasRpKjl9kpKbdlYS3rRBZPBusjluQQ/zpLaw5fBDHBW/xhpct/VxvyTXWJn
RZd+MPjl3AzIizY5CqcU5N/NiZuz/Eqs0RBDk0/jznmpoQwc0d5fvVwGYNpRWE2Kk3/eeBwMF9Yb
OJDICYdhMxk6liO03W1oogbrv5MEE8ocifS99UgrCrUM+Cpti27RuGprEjoM3XWBskUkE+mTwJ+9
ez5YY5YHphUOGzzA/0Qs/+fz5suXqFWFAsDBDDNR9PY/ldJKzo2SMe3MVwyXipYWyE/UIfcI3ZAJ
8ZhVor5OFQ14BalNPUBByDF9FooBFxF5TXaoCWloZEnQTopdS50r7EU300F7+BWDrhcK3m94IqxI
+imBALpc4SPl4DEYZc8WeYbJFzBY7UNY1o2R4uwfDCnNNt3O+EyDSdtb3PbJdJv6+QFilj3qYAR9
hzlzyp+u2KCPJRU5+gAK3MF9cqdc/oz1m3S34u1A5lFAGOUPjUYdslX/aJieiVHvw7AMh5p6ETCm
avRA5GCWtyhpgENo9xET67TRWCxLsMEVLm44XDmFGIVz1pnEsWOhax4ujFv2YQF1aMUjLUDLxcpx
aL4cxh39aOH/zJNdV2TSf3Ck7ySRrR0NgBCkA9w25sOi8ETcQucR4zRaH8//LfuYygTJtRJd7Rtv
jGLf4ruu5Al3Kw7bRospaxsxLwdac/Ku4qjgZsW9s+tq0oE3QVCpdaUvok+B9a/vCAzDE0z8TbpZ
5mGk6GQXQ6gmrwJ7emYQQ/9j/214WH7ZGI9R/W7aXBCLH5pfmagZtgHsT1rHy0qKLX1/KQCakN4N
v4bj9+uqeGfjrj2zW0n6N0P00TsZFsLi9yV9AkdmobRGDegG1K3yMJXoVON8yutNWcDGOKvkkvP0
2cWVmzfS8mAamazPTRcch65BnLkAnfSW2ZAifL0NIISY8Y5V7I8YwLw7bwCXFwT4Morg5LVl5jVW
E27I6DqtYco6i7ydzTcjZATy0jH51sn+jKcv3sbnXotRmHZ64J1W1CWOOq3EylA3zkxO3u3KnWqz
6kyX2In85KimLdjJbHgixincn8ybOwdKtBK5KlecVT9ZJtow1if3+rQMTEZ7+Tz+T5mps/8LnGUG
Yg828yK6cuyfB9CfUDVUzhGyxMIYvRuHvx99Bgee2e9lJ/jjWb4caxOHVm+H8tTxvTFMQTAHtMes
dpXKez8NfBeyflcxz9PAZK3DtvEpKBlxLVIxkFLVXaow9sollYG+xtuU1SGJ7himkrNzOYK7hi0T
QmghNHLcOam1qhZIYzvUhLg8lvawbLjdK6Qcab3THPSNfIIkKsUrD1cwThutDPrDZ2rKoEOYiT2E
URhXlu3B+bjc3hgVF75B6ElirbhR9AukidsHUMtujH0aJnzPc0xYZb8vcdJYb5I08jfguP7SulcW
VIuCH2ZuB9r+Dn4ED0cbluP7TGlr6jo7A0W4Cnfk+TMYO3+47VviAUL+J3SUBBIQ0RTfWGf8VHlW
2lssq8kej7+EjpPL1H1R2pZOv8VJO25AurI15XWGTjg0/lqAC2QQl8/LqUypo+U2eMDZBZt3pSRN
fdVVwiU/FaZKw9q1pmc+i64LOLSCR2AEgeAyConXlk6liseu1iS1xn1evupJ/oMagdKtUqkC48jF
S0L1Wx4XrDiCQ4T1qEQ4sVDtbwTMlrKj+GcRL9fhBiYUa4zI/FtCJp77THNUwXIfFcqk23BG87d9
mwbzKRG9EQGyfzd8HabDemvwXXSTbzc2OHdhMoN1t872qL1W973bWfqutXW0gD4zCRLl9rpnGfi0
zDWSNgU64985vOCoq8xGxB4fYf/rkD+Is10zzbdxzvkSpJjXdfuB2axwK8Dm3lueuYEC7X836w3C
IfFNFHMJwHqWEdyu8fRXZjw918mPnwcC+/2FJXqMKPDs9B8GbDPSWphO2wHaSTyvIkwiPOaxBdQB
xPs1ncWSbFzRrioVdjGQ3+0jrUJIN/Sd8D/H8zR/UF8nHOpi7B0UF9FynpIUCzuYyGo54UO2ThP5
pjkm6XF1marJza8Rn49g6iu94LH8ya2SkL1uuwoCtjsZumOhvUJ7szLpZTjnFFkop0G7nps53QYd
9IBfHpzVS64T0Srjup77TzgeTzlQvX0t69yW6XhhOnkJfhxhE/TPJ2xbv39+Km99/h7L2UWDH+Ea
VjmnzLSuwzQoacJVJI1XQm23ZjbocpIvybLixbcFjpYsAsI09qaBTPqC99J0jfAtYRd6NVqHJ+gn
ttSva4rsBx1GUuXicUCnTdPEsl8pC+kHW1Avt+4qdjNh1ecYouIx+gupHtHUY64jCrrBaNUX//tv
8ndzK1vAPVjIsa8NCGKpkAvalhonDz7Dnepzia4B6yserB1Wp7p9alfQTTTc6bBf+5/NjKHNrrNq
oa25sT7j6aAkbfx90FYd9m+zZlIAOY5goVexpYocTmadGm4kDKYo93xnEmAKXbWTuw3jOjGbTrZf
61VZl38KkCqals1o05w0izGTwqUaLBdoGMPEF5+fmMfTb76C7SEDPkyPDX7zVf/TQcd0+/0o5oEa
KAjoCMMtjfWgIaaOzEdJRzuBeXFQ7RNkFsd+MzQ668yPoXxp/JEeJxg3rsGxForV0nLLTovPWgQu
XJgx0t9sp7Rl2S4gz8FKzY8hTq5TJszG/+wvyaScs88gFMZ4HE2wB6/64OKy+7onOGfHdV0wGIps
tE7nzwuYo2NGz0irwnnpSefy66C7F7bNbH+IeXM11V9oReCkQN9i1ke8tQFHN+htc5wg0/PVSFJt
nGolT6utGTCnwedqGnFj004nBVPcbXhOUb6xvz++I6tU+YpxMxkdpbU0pf6eIMlNKAsRDV3Wmm3H
lTlPZoG/LNsKc9Q/Xwbqvy3q4iM4rFiAtsFzJqG2Pxrem9NeP/0isJBOWxHY3aXJ1pXpV1U1Tb5c
kGCo8XSMe+z13X4A7O+Efv83Lb5gDaWM9JXKSfwu2d3nphVKeTcBAxF2gSuTmeqqvOBhaIcnLszS
NMn8hBcYESoLGk8/cUpGwYKofW7GDKym0m3AJ5SmWvt3xzLPXwiLJPf9GeIBIFf72z+YtZ87ixDD
eSuJTNhv8d1vN6mxwdjusXwKmB6WeKJK0u097Th51VD346E2ZGp/KW+fhwxClcKM8SVppfM6YKJW
qROGZRDZjxlprTsxWZvnMC1knzJCfckAHShtbINcfG/fyd6pWF9DmW0zC273aLe/eJjFCYcEFBtL
ob0YKQuKN/rMk7K2N8+Gp7wPDp7HfyOuAeEO1iGO/vQ52QO+1SRiHvg3lzFGBtYlIbm3NQFCoRDi
WQObnuTTJSmPSf5gTAVcG2THUKEdgeg2S4/cm1BHf/SxA1QzuiZHfR9M55eeJvOFpj8X3FUdjzrt
JkuErulvYQb70o/C9NAxqO6bT6S8ZqQYIym5U4sJOU7AcfvgofSsnwCH2/sKDuUctAXuv4dM1wBQ
UXgNDJ1JD/vXtWgjSNdTJ4/0SvziVIDYRbjmqlC8QEfF78h0//H+gnSC4WAKKyNtjfGVbecWHSlf
dBlT9EA0ybpQcMyCd7ERZnBl3doDQ9UdheTfHlFGPbHuPj+5IlHWGH8824c0ymq+FzMlg7JdSkY8
f4oHSCN/ckMtyn7eBhC03eDacills2SIQVXpPbXeVXW0PUexE3wasBPYQhdjt4g5Pky6PmSWGiY2
rNW2CJhWsfz0XJszayucJ7dvvFxxNVRc/dA9m5a6U7cA8aRC5b5M3LA+k7m5nKa4M4UOOVqJxFTB
JIrSK1fOzsB1pGP6ttbhNZtakykumyXsPQ6GcG47U0O3Not7nqSTIyzW8zD4J1X9LQMDOZsbGBxq
ruQX54eZXp+dsh3/cMt2EdkP/qTL240+MHdjV3rjZCHCEhCjbEDYesoszzAMn3KPDd+wIXxg4A4a
/8V5CwHFRfe7AHzGIdw47sEt20OUYroouAtWS3KBRP1/2sDzXuu6zaV5vBI0010/+DoGnwBccS8J
NU3mEbKBCFd1u0BtjHszj6fmF14DCfrTh+vcMP/Tjuw94hUbGWQTaFenUrim4AKRtQ6rD1x5ePfO
LaVA1KOupYBWC68rscBQMEJXYn8z6ruqgw7Xntyp4NCkdrjvlZdkSR7h9yt402khgHHvdgwNn0fv
KnFPFG71JhkqICSq5B3/PzE7hWSnEM5lDW8EzpBB/OkXwPujHpEryZ+d2ze7bLy1ZVS23CM8XxjO
J23+KAQQ3sXjchjmIoMwv40d3ABVTa08PdI/kWnUe6DEZZpA0V4N5HneDydwOYy69PoijG0sFlbj
j4doI0CxqQM1ytha+uraR9+D2GMyg5LJM1/HVCPPDY4lM66oJq40a13qDf3w7/LdFODnY9cW6mpe
Vzz/E7k5HzwcrBZJ9AsxKB5fPVzs/l8mLnKMhqvvLUJod55UbtvTsuTABc48E4Edn6sijCGLbWFL
OJY29FLSTO9KmiFlpdW6HKi/7OP3ldbKJbglyxg/3CAcoTgmUGIsdeCwhji/BJ5VbNR+rQEKgeX3
oYm7Xgqwb4yY7uSY6V3v/UInS2SKbTvQaWfVlCP0h78Fc4xJC5oHmIlAcWcG99ZFnEUELGZthN2t
1tRiH/UoB6KphorHU8N2VRTxX+5LFZrEzouYaUw4znyreFm7yLNuxXiY6I78L6XsWHjTRRLM6Yse
/wQKNgIyI/ujrxsAJuU1ajIR33MznnS1abXZXH7hAk77jGR+s/viabPejJArEOVCazwtAm0s33mW
R2i7YQEJP/drR2jrilYVmD3F/HLWIZsz8YHk5H/M+XhGTioIjmE96MbUsFPudDu6gjrg7escfO/R
EwV1XvGgnnlzZL7fN+cAsttQOzZn7A3ugY28row6I9zCjPKLZoOdwivE6XLP0O7DvOW0miDkXEOK
vkz0kX7nXP4dmhNbBpunULR/oUu7rFo1TfFr6hYe8PEofOo+nKhg7IfJEQPzbo8/d4VHWnZnb4GP
Hn5zVnc2QzBvd/wZSEzbaTlsmUTddI997GxSomGLzklcwNIjCGVooQ/tfSLMHECpsTRh1nnQA30v
7MgVau3NA8astsTAGP6NEQ67XXGiLsfPFZ4RbCtEB/1NNUVmPVS6JI7QZQNsxcEW42MmbKGgJ/z3
M4lyvgXA2u1RZyqQKW/ob4kShH1SpqIJcJTQptLNTyWtFm8Vnhz7T9vU2fqWxd9Zs9cQBED1KA7P
muQkqj7PqrTFzO6PMMf0DpWpM6OdaerAnCTn6ZNWGYDcYkWYA5rYFbd7M8l262Jb4NJWlcZTkB9X
ISy1yZ82t9qGc5+DNDMCQDHfsnFOzdMnO6XBTNKO7cirUo2av9edZapQwhgTKaxnbzWW5AFwltIA
jeDBT3d5Sdh8wBFtRxwuJoBYx7ACAL/muUq+NCo3x3Ys2KLWmF2zk5G5z66NDkHsglhpzpOAPzBj
6Zddygcbd60w6xuPaTHVzP9fw0SCUL/+vaonXKMHr8HLBBCg4Mvu2qCoq3F6zn19o8XcipVkYboC
skP8lxYqyZfmiOnJtTeqxl22lOovFNft7LfFmpgLSGNN1Kh53M9UJdYSP2RMtD94vVgCtFy1WygM
lBXfKzbjk7c6mkC3EOO7+Fsvx/BzBx+3lwKHQ+ZcDcSCSsGDCzDhh4kqOshM6YPJkgZKUohWPOVd
zI6bJEYNxt4eLDa8oT16DbApsjQFiIQAVz32izjodLWgpsw637CLSD+FNtQoETXsly3jJ+hq7Lb3
dh1Xhka5kUnKioZB0OszTIBAuCzLIoSvffKBRqu5wo7tBA1rx1+lFHrb6rzNF8e8nhBcXMF0f2Bm
u6+GUuVJuOAxKlmZ5IYY+qmQ8WOCd7kAyzDKNwk5dY8PzWARcrX0KsB5F+6g2MWuMsPtvXoPIrey
rwNFid5n+ExL8ED/Qe3DOE7fwmiUkBYVI306jk5+jck+us3V+WWYeB3lSp7CB78a07OSHgH+fnkp
j0i+TWp46MDhqY/znDd9YwhjyZrxCEzDMa10V3FGM/wtUYA+Un9rX6qbUFp6eENkGNygN8RDZie+
IhxHrUUrXSbevIi7BkKf2otz5talrxL0IofqFK2HSUw+YsQHAJ5leQCuFiCLfsrPKFyJ1dlnb65w
h4jEuX7gLIpzuCjBLmpWmVU8gAq+7Y2lkiwIeMCEPelCtvIDdqjM/ESixdlm8EEsRKKCclNlo0dH
FeajMa7V6PwfahmYhby5j6NwkHcvt2pJqe/ZCgCH4muY+WFIddADDohxPhkJCP/Zuwgqhbyer166
5OVpuTuDUuLyImpC1AJZMkyaLcdb+4OuzOu1puVdK4SnIwD3cU5bvyIr9B3tTjWS5mBFA8P5uTbw
oVt7vStLhBUTkfUZ3vqyPuJ+JlC5fehTkhy82Wgf6q/5ditoq4h/+J2F0O5S79LanHFtFYwg+BIW
Gj9QymuXyPqOBCBH4hBUMDzKRhjw4nak6leuq049N4pAAUdOSnhi0QIuNXYd3GW3RBTR9G67T9lJ
sHqkL997Nh4IQtHtavDRBjTG1J1OeFPre7CBInx5zZ2V22mWRTjD1KzGlmSxnmUnmV/Y2R2SiCfg
V4qhvCv3PKGGn+tW13wscoiLUvtBN16g/rAj11M7eJHvpU3syJqtiYcdC4UDJbEcuq5k2pA0XpsU
R9nZmKtqSshg79SLBeXRGq6sphLURiN1+Syrb2vlsoxOJWIanyAR6+URCMVLE5UvwJv8rIIXlzzF
0YYzoI9mgbhR2SN1EJDnDowqUTxTMwB7Mtj9M95izIFGpgwNIJM5vf9ICbk7oBymhkp68YY5jN3f
SNPf5skCcHZf8arE9BkCHe8cxsp6UMsF0TtYuiCOD9hiz7toQnWCUtNdRgym56KhiTkNtunDhg9N
Gg9Jjt/cNqrsXrk0yRo2xP8Htl7ei+XVJsY3T7JivgmAEcT4XNLEkeD/berwCq6LQF8Pe9+tV+NE
xaaVI74YQdpwAHLioz12mkvJXPrPlQG6dmmpcQj8x6QXKyiehJpfvmRfd/ekAlHZ5IPhU9HvZ25l
3mpPQJMXVgUvqLNB23M1v9jC0n3lM24sUpWhJt6xtZPWc1iXtWpPP0Igfq2zXHzH0bbdtWt0OQJH
IJ93yOBwJprBMMFlR8xNPG8y/KNxX74eefoaqUW2/ZobPXV32tEipGjCX7TUaDhDj5MwMsQDr9Q2
WutoeSwxBuVCbha6t3ZX+MKGvUfXXovFIrw4YiZMQ2DeMXrfX+N9+C1x33rhl08xC/9T1t0E4+Yy
sA0tm2/1j8CM6bd1O/g+PH6lfZ0Mi/kNNe18b5TB57Zs9ve7nFeY0zzszTF2l+pmEoH8Rsg/4cVQ
D5CQd5lX5MUYrEvZ5jTDVjnJit5Fo1x0grSYDOMGb6pd1iFChXEVNqVcZABpTgrwOFzYQC3jwHLo
aOELzh+cECAUfooMyQ5G6amNAjLFGy2X9GTKAWkQmb0uZGpU65qBYMZvTNHXpP69MFcSGn8uA1IN
6Iv9mSQUCd2TRBzD3SjxXShYcpFGMzcH8oxK6DO2ILt2BJNUexrTAAz2vFRHtvKSJhqA60ndQ6dW
R/rqpVmvim22rqThxUP5O/5uuZHYXQ1CHxkIlGjZbI5Lk4v3p9b/WxJykFwTVeAsvbPEyTI5W+fx
neyicfSNg257MGUBueZeECAP2xWNqwo03EW6TxQJAjiGw4ciwIpTmR02j10ikG47Tg9N5pMHUd65
IPYwlg4kXotVXTnK5fo4Hr02dQkwdWaG+fY4Dbz/rtWSStInCBh6U1cwFz8RiuEmI7oj3jCaeiwk
iPclzhS8wXnFYhgWQnn0ZoBGCrCAPoTzcNIOtZonfMayWgebNRsHJwsXLflAhXdu9aX3cuNSqg9v
Q05wHZ59ADvrIoxEI5JWASlBZl+lU5aXlLDdfHD5rEtQMBAw1W+gaQpDKq8ftPQirGohDBPxJdwA
DNawo4dJIUyzT6q3vKnqIqW2hAF8YxdWAwSCW6RArACSd3B4RsyLVhZcidrPh1IVELbHSo4RET/t
j/Xf2+jY2U3OgQOf9OnnbIh9DNp0Fe4YhGQa06dihyQrVRI0tOBn17ASEBAJYcP72VI4rZURQNy4
ZCAeLlTulLF9QSXLI6QGkVbQGo5lp/qtZTeDpJzBNcDzQGzSCaYpsBfj8w9kdjKs/2jQPo2XEaVy
WlJot/KI8MPX8XuNT5Yarn8NC+72zy/RTRRe44nEdGImmluR+HG9aDB3FQGwOGZdf2q0BmGZA9QY
RFlAOnIzEXzf4ViIVrVOu+ZJ1iIe9sFidMzuOmCNJscpPT0DIjoa/wNhex5u0QQGxTIZ434WaxQA
ypYJd8o5oaNcag0w4udo5J9GqH6ePQsnbXCdBBMZwrs+03zUCTWRnneKuCXbYPcjoYYMypErFRLf
HoLAolroimzSQ6TmdRDaPonbUfoSopLWijEySp/6AQsIQ8YFO4pQ3hjVpItRXuDCX0Q4YgY8Gtrj
x2T4Ukputy8FJZT1Jb4gLdXSBDL+kT6rSwnjPTwDrT7ivmYkVQO7s5zGJoSvguykQ2h6fW5BdiMC
r2OHwBt14XbiWoAMqDhzJlWUoZJCzigmrGlBiiMRx3pYJfh6TWztI8JAWQJXFXBAaNbJ/GtR7eQO
WWdFuBWlpNe8JwAPCkD0RuBAPZyVy8AGRwm5c28rzWaz1iJIX9pC+QsgewMTDwImA7eIqqTC9KEW
j2XNoWPsA9Rmu17zG9osbw+CvziKnQ+ltY+bQx8mpwex7GhZBt/cuF66UzbS3cAsbH4rv4LdKZU8
9aIEX331D5ICxMt4SNOmfWVdUIzzUVMXXsrEh3ouCAPZywWj/fGIwZ08T5FWH8Eib5elrMloXy1b
bRTpUetDi23Vil/06vOcd3ZE2pO/ktbS12w8N3YSSKef7T2POdNc3fRdX9jpJ9BoWBfgUxtoS/2I
i6fJmlHWrpvF8B7pMyNgiW/PsSX1ZBereakP7xDPNAjuQmZ7lzHr7HEUwE4ejQGPfudGcsSCAdaa
8zJr5j2RdZhicpnT60YWh6NLKkQWVp2h9DgViA3ZcFGMPXrQIhjfn2ItcjpUbkWaF3kxyhLCP7ep
5KJLBddMEd2b6uxmRch/7tsUl0AakZX7o8xMiUqwzW3CFLpGBclG0aGLEm7JIRgEvzuZMtCnJ0FF
aM9Teu3GrUXuEkGFFeSja5ql7rlnY2ER7/5FLgY9tBFewIkFff29fU3ObriYCB5azRdgBETej6Tl
lDg1EIlUUPx3dGX7tZFFsfXZz2aAi95hl8nljo8O2YgiMLUpdySqhgsFsfmmGBDR6Mnhe0yGprye
wCuW00zE0TS3UGXykHlRKyT5tP69iYQozhAL/DWzvhR0vJOUHw7mt9Akq68iJEQsR4K4U3PBew2A
fP7EceRmftEes3A1lfmuOTjN/rhkQdRBZxol3QTTVmh0oauIw+Nm0f2mVNcECD79URr00ZhRMrc2
tPgRSeqy2mWsutcB/IvgvK7Hx8tot7gTtX+82lFeOWXGSGwtSHdxhSJcT6VvQji9Ljs6fAvMhadz
m9icrWG6lWoYVxscT/TJJun/cS1AI6Ij8rVmUhm4KcH0I1FGmowmROqQrPwDja+t+8OM028tBCae
XiM33YvLZNVMYB8tDY72zZI1g1eBCvrSMSIU8At4yVnwtpRlAgHM4AyF6fvwdLkn4cVfMpwFPDZu
E2JYx+CsZzXPx2t4yD/Sxdbdw06ILM/iB+RHh39J4tITdX/tkySFxTE59D2HCiw2MxoSFBAZaRlb
MY/4bp6mrh59qjkCOGAxHLez6HZlBY52Ziw1e/vRxVP23HdhJ91LfVqH1FTjJhEqC7XYZxd0oRga
uhYYu+Nht0J6HOi3Nqt8Qf+PR5xcjtfScUzqtI2wY5fpTwyWmGJrtkiBA0qKNqbSnfzxz3vadRo4
nLJHgAC7tS/hBGYDjlxKrO3EEw5fVS8hPbh0utuygeW3rzFPdaQfJznncd8CjemiINnieaM+9SHQ
x8gAOxSO8OB9hPh+aAbHnQEjgOPFMCYlwolgoibeyseJkga8p9pvBB2FjZPC+jZWZf8jxKsmFFEY
GOmfTinvxysPcETPOUbNHdBP3nLxcgx8W19mDgH4FxxmePjKstB8aujyXdDpWF6u0bl5tlk0jUJ2
380Mh6iou4PTVN3d574khU7AwpAajsZevuliqbcFiWOF7T2nafAezFJdUvoaTyWCBuQ0owCXgFif
VaULJEF4WOHSpyHbPAN+p/0GbB6npVP5n0OSfq62EhQAf32PYgawKHeyMxjylYeJJqgEqcQ2J2nY
klrMahIXGE8p9Yn7snzni72udBNidiscGnj3/52Ote8zkHdinMvjziht/Nl7VIS8bryibiKCMq8P
kYWOd5U1JBGdhS6FvrKCbyeG0BlT1a3Rz/Re4aWQX6S4rxioZnRR58UZclWZVS9jsh0+v5dVgx/d
p/4nPoXfVJ8QLHYOcC3QTMRZzGkVS1VOBAZcrLtBlXDEo++bep08aXt1VdTlj93XMAB/0e/jBLvO
YpEM9n5aBxIs703coDfHE+2dmnuOy/qOwEoarha0esROVQPeELJdbRg+cMIBWcMaljX4fBrXsQhh
LcPOK0uC/AeFHspCDzZEk/vW6M8K43l7lny24ov+GBI/IUuq8q0L+QkshfvGzHA/Gc3NHIWrc619
ErKStbBqFdvaML8FZS2G9JcjT9ujRqkb6bkWYaUVQXrsNbpgkmUgHafWSHtHWdzSpg15+GaDcCLK
fPHFkCbDwzaQYcpecL5zRTVnTzx5f1nMxY1EJOY2XYPGrAM+KlzV9pfFJKssHsFZCQUcCepiKggL
goegrs4yYJYc/cpCLpPK5YTkk2RxW/AHQX+OZeMD2aFk6wAZZ40WkpqV6K0gMirQ6kQqTZy0Bufm
aC/8IcTLoe6QK2cRRZsmQPTgCVB9Mun6fP4XOh/iGUj1rV2be7p0W7MJe0pdG96+Xent3eKffpEk
gATcu7f52jOvPraeyfRye67MYYW9y8/NkvOEnVI1b8mwT41l+Quaf7k48/OJ2p3a3DNPeGmd0sQA
eu2RxsCGbonbybtL/RmeXexbk9uhNCGryoIdUNhzeJrmE6f14P8V1Ue2JjVjHaL9LVv/zZmOYaOI
fA7bYu/CxQ7JOB9QaMXwylCdPlsBjvMQECauwgVeK3ZXToyFDLl/oi9kUp33BnFOx2wl4tYdIkdT
6rlE8h+GNDXnJM+ismFOszlTHxRibYU/6BENfc320qIuUQI+clMgln4pcahLVZHivSOD3qxmsWzY
eCNaBWdcFwJkExBfhxuygPchjzT2sXE40XlgCA73cweQb6k43B2OpzqiVw/ir8hFo6k7qS5xSQHp
k0io1roT4J0Mq+dpvpGWpQdxIlVc7y0DgNHi+dEZAEZAi/ymrAVSDNtMHVZpyOzCq0oIXOBxTdsg
RC93FoJLJzUKwgXjuY5LhB0gEBN3+C80LeTprlX/LTIhsfgzmf3sR+5vOCoER7wb+2wiCYKV4Xop
0VK3oXJ6WDRe+9VHQ4WsZwt/soSFjdnRqI6OabO9JMouZyXwVcKHWrF+Cy5hBGj8sk9G5duZZZU3
EimPyhiWqUcVDFtvuMnpj9sAdJ8Kcsc4ttYpO8da0UT8nuoyS4/zmd3gyNWMODJgeHcJ/WfwV9We
G0M0J1PiVlMK8lhO+AFlpd9rNRMhbPm8Hi4yIwPjN9oZpsnZxxPBc6WRMcYAqZdsWLoYweoAweXt
4CL/CjqzEphNci/ABOMk7QMgKl7KRCgAEiwKZMQp1uVOIe/c2Vg1VjHGMJ5BG1s+0zl+hXLrf+eb
Z1h7FA3obkOgDDpEG2l1bPZ9q0z1tj8JYDrvpSANu/uGCxhUKl1lGUCoABsitUa7rwNmZMI9Cjjf
hCQ1zvIrmqij94/jwnGBV5F3fIhUGY2dZMqCaZc3OWRM+8YRg5e+nHEAlITrhFcyqE/4qRHG7koz
7D31RmQjl7TtBd7G/sNqfR8X3TbQ2ZZ301K3QxQq+jAUxZQKafPXbMkO5OC+kahUEfMiyPjgbzfr
oEmVRxNPiobpJutJqqIh7hLtT46PB9+APbRbpUm142uD3wVK8/CYZMFiQHPV72CNQ3LSRe4OPYsK
1wzordIBVMgHECdhoIH6usGw929QzDJf9qAGNTEZRkLfmcBOrH8LUkr9H4N8Bta8vrgxZRM294lG
kxRqKCED8umhtlIE8y9n2PWjIWiZ4mKCrq5cxHU7HUVOzz6TByowu+uL5uvH7H0CRlOh25Z3cQbt
n0onScyquVmHdbNRhd7jvj29K25pUaaALYC6HO7jddHKRwHcapQGyS+acPXw6i+3zeYWeVuoAHkV
0OHiSYqyuZOn9nJCJFcZV6Q68Bx1eCpn/FIxHpJDMmPQBC3pWA4S+nGOHofaIotyrH02uuAObRTs
enbyL5qUzmuyMo8YnFFPAGvJf9hSndat7IP532AomccrObseDHe4Y7cTICzu98RUtZ6aKIlFuLnc
r+i2IyZdavH9BvCzCophg8Fb7UzImkQ8c8/D03o0gFdTFHm3mHhLde++2qsULRF8YmZKAsA8U8jj
IlRA5cgzMq3LnsuXL626V6QpKJ/9irfvfbel/6lmrUWw/zLRrBT8CoaPs22H+K/8on+QZrYNvt92
5qs4yGvjzCrMlFZTVNDuwlDg+xqSGHPcT1ylTB5MLBUKIaHnFn7VatBqgq5KPFosLqw6zV7k6FW8
B2n6fAihilFTjSf+F5GeF2w7gRlT0moNSMwyvhT8DQzh8qI/42P3BUUxfG+KKjBZ8yasKR4FDNMj
xWKrNmXlO23wc3/clBxYUN0NPAd/iyYgozYWqgWaN7EeyTJnqyAZk0onw3rKYZQnWcZKt3HMePoN
/3yE1pKiTZd4hRqJG2EhWlQd2y4JScpqLbO6GdVcQiIIoAtn5I1L/CsRj0rbE+SSf5nBEK347KNp
jqUI2n+ugGR2KkPDgK7226swASppC7n97T1h9DkN/JxWDfhLf7nFW07uOe1Jm9RV8iqNULNSayUn
9cd71CqS3UwZh7dcoaq7St1KeiE3OsMnaddhbTJ4ywOQpv64lYHNx3rvnSyeYYvcQPAiB2T+K/O8
riiTPM5S+73V+b55/qQtHDwjFpZTpMvtoACtlCtWmrn2z/tLeySiZ4xJf4vMa8G0ZWfECwRxXcO6
BOIy+oWB2NjMkdvcTXbCiwbuMoKsbz7IW/sSyw3n/dOvuM1EEMqjKon8Gcpzn5bDD8Wd2WCljzWm
wd2f2+Oz6i3fL//i9zeHuNO56+c3sn3Upow9hdo/6mXAVICQpwDUq3CjXauPIV2Wz2/l0DlxYRmo
WhtHfrOIB8he4ZJDZufNcwQUCZbsmeCGKpGr8mCO9yvmjQeugZpZA1PaRGQ4+RUZuz8ssrYU5loy
pv0ES6AIak19Tec0t2uma3B0kTlQjuB9k3Y23Pryg8bMkW4x7zGiKaQz87nVHmR2aGV3DCKjZhe1
OuuFOrEIHYlMv+eGW4ZgLzarvCzpkT0kr1MrpgFUEGAbG3Wr55MAgpueGYl/80MzwWRcCbd+Zocr
kSFV+khOB4uJs3gR12GicJWRqbw57H8i40wX7QJp/SIUTloZR/BnA+knctn6LLE9rEhM1vix97e4
XSxrYzih09QZ198zdb+lg2RW4bAeRwCGiLu9LkfbWgYzQ1FzSB35tzpf1QKs0zPOjm1X2zACdOc5
0Sq3A2vaup95lDFDb0dRlgYJmjgExVYZPlzkBKCwBdbdtMotvvhSYdUAB98N2SZk6CtNfU+xsYnV
mRC3DGNl8zvtdSjDIgeiZUrXTDygW7RRC+ddak21tgJtW2y5OvZgE0T4BnRZeZEDeZ3tXQRb9nxS
5Ql8ORTdHCiwAp/FSvSF+Pm4rpjEp/oLbUATKeCzFqoC3RNhHWLmSmMACnRHbZ6HqQaScV0lC8SX
4+MeACWXRWTRqM8HwqGJOOtA/ok4AxdRjeweRBC7FiKDGY/gl5rhf0uJHwcGBT7aIwFhQmY84u1c
iNMPyTUD2dU8DsGF404T6yIq6JAa1EMoZDMLInejpvOQohR7PX087Jvv+KngLoWsNP9A609k/xbP
4fvsTosCcZ0v1knrVDSdg0mJgbLQfS24o4rSzekfS7CSiCKHQNXQQBInzTHmG5Zpsi/g+u5kcZE1
B5wzxAE1aULvx3wyDFhy0UxOQ6n0mqZ68R51gzDfNQ1599uf3brBZ3eqidxYN+kIq1ePkGHAzqod
Jl32eVFPb9HznuGAuhYpbElDBIeLh8b/FSmRgm4/dE6i0O6i8XiwNvbAUf5CsDffU9Eyf/wA669U
yz1pWi2jRIlpGKXcJe8+UkKCRccAErAsGsvxNQB0nDwVPEVr06KK1OcZT/0K7G7pkpI8ExYPxZiH
WHMr+GC7/rFV9qHMbyFPAAAGKNjRksTwOUHBUXQqwt4RPGWeb8e+X0nphfPvNPE1aa5Ww1cJIQKL
tUeRzadwXMPvMcS+N6oXqHoP9MlboLkvCPQl27YM/sNkOfBle49oOsE58tWYlKYWme0Fhe2/6rPX
B1FgJ6Jmr8iYPSFUy8eoDNQIMd1xZRe1+hzgCmXBddNr4BvNRiDR8bfTKGTOMK8H0Ys4ZYEfKCsD
O3WIGc2YHRZhc0vKpGPtAueSigQLkwzpv2O3cgBZiUsfCH/fYOISgSHOwTh+B1zD2v+/kcB80l0l
lVuP8oPFsg7nFpwGTgmoJljiWKCGr5Aa7V3FnvH1o8nOZhbGqU98DMvdlexkHtur0l/fke/QgQfC
kQUskR3eSnRoVhLaFl6BWTVjntT6HdhdLR9iTHFF6p0ZVgjL3AxjLw+TX3plBZs7Dtgqe5UQ2Z95
XP+rgCsIf629ujhxSHY+/T52jvGHbeOoMuD01ipHZLHUR5Swza9+L0TMtZSrK7lPJDJPkpBA/9p9
mF0yVAFsjs7iunZ76xo4PHByG1KrrPmHhs7Y2GKxUcdUgjdQjWiJI6DiOcqBw5xf9SS/YinFv1Xb
S6mFcihMURG6csugy7xpRiNLCmYShyBJiWFHKe6sXVoB5s3XPaXZdmY7kXiPpAdiSN7Uy17XM4RL
J+qsJmFnoz+lTBCvyjT7ETwn4GWu8HrVMuNwT3qHfebRei8tqWKYP6zga6impSqQDgq0r3fH9lHc
q3BwUrwrNGAYCdhiMF8QzxsMcA2uaTUaJrHr8wJGg9VwXSLSR4ioFzDbeV9N0i/D7ILPBu2BHgId
SlV4VLMxFBLGiyrQ2kcnZHA2pTbqr+u8/3/SUUhQ/7v1ySEf9kgy6pjP7hmhTkklfBGP+T92Bspm
Y09RVVQ69pmjz5VcUWtlGaEISd4Dm/qDMKTDXHL/wNcJaEzKG4GiK9M0MzdP1BhL0RspH7tunCFe
rhYZEVmshQSWOIBNPvt9SmdUFf42gvHFtxhs0fwYGkR7Tn97IbaNAyJWAl+x7cAkod87/yPXAFMT
NMOIOEKk+NiSrnKo69Xq69AsixmTvXnVjet/CLzUOYYEGhQk35o5UBS8bMMXGyNg04SZemMyzWQq
lnEqvf4asX12ykFQBBGtRs5LIqlQFHVtgM4MVUax2wFf0KLv8qQxvdfS7Cnx1hHSeeAOJiJbw/dd
FoQcqkSvbHvn3CE8C6cyxLzbYjiG0jiHYJH7BDLccqSrLKdJAXNBfMDoIEtzBIeV61SZcSWCeNrX
A3ZfhFkUM2GcToTFjyHBMeU3ilOnPmhJ/03f+DIoCc05hwUQgg9AUEc+B8j90cK004NMU5VrpLtg
gJQJ1l25KOqBB5fkkfIeKdED18BVuaRlO/BhMY1zSzq+YDG/eV4U8/o4sH0FVAjKQPed25Fh5bTB
J1X5rsjr7PyNKpMX65G7qhx1B0H/y3WOBzMZwTiDg7+OY21Da78uMikpIk/Yrt88Rc0y3kZrMZSW
dIHMWval0rJIbhbzvdPR42bfMt5NoedX4ArzSJGvl/2kfHAMWBWod8sxKIyxIPbnFhQOrbeNxUek
zstWOlphLXq1SE6M7O287JWUY/JPxJdlQ6np1cKxU78jobBAuSOhtJjN1OsFg3eQhTnAkkPlUrHV
2tQRTHpgJuFZ3GodhcgZFNcU5bM8e6CTj5xSzsXETfKHnysUItvDZ/HzIyvY3+KXD4Z7mJrVslcG
rnmrYDeERHgnRvO23hH/0bwD7jl3ch1UPEYBfX4YsfvHSaKxZP2GvOrBolqweebNDOVR/VVOlZfT
dwimHhzQpa7NMMJQABGfjjIRyh7EcMTwzRu6xNcQsfJAnQVI2tTKgnIlUrcLFrd7epPsEmYPtE3F
lHrQ57oBJlbcowxrmH94KWBP+2jVfrgF2k4IkOIC7HbGkJg1w09gWUez6ub3JKIkFUkrvFIKnYXX
aM+7KhG+ftZAsu8g2YBn8Bdfac/igwNYRCwnnk5Nk09f/rQfBEHYooAkVjFqsdX5Hero/inWBpSf
K3JdUaeuUbBK68HQ30uV4Yrh2WPlo3t3bFG/Fbkq/WsdD0CCaFitCJCZ+1TFujNHK5o8d0kI5VoV
xE3iBFU2lvO9Aklo6tUaLl3OCv2ze+AtA6RbpnhC5tjnPBfQC961TBn8gD//xPh2Yp7a6lIUi4I6
BU4+vHOljQ4np/gFt7oz30XFxBBVOmK20hTuy0D5hBjoOB08+Cdf5thQESi4hfcZb/E8zvjtfFXL
7tzXMiADd3/WvMTDQGD2phlhgL9DnV11Q0jqAckdGfXlQnt5OT2p8UnhGUN0rjYRnxLRgVjUe1ix
jzP8JhsN12+rBuXLyrNC1ppQZlBJ8pPmeZL7jIr7Acvx4ftpMY0luPCYBtd5630hev2pMes9ieYv
xje4pHSpVgODr8rNC8A6cXRluLFzup1PJ6A8N2hQRV4NYl2MUzDpGrBLQqcwwahUE7usKWKZvo0i
9uybX9+0LYrX2rPiTtTDRAxuXfA4jTFitwz9wtxDaSGKfTjxl2SYr+MtKcyye21v9JqDC9FGmOZL
hprfLjqtf0DYWxsp6gQxWtX6cVJPr17Zpyhkzcz1T74eTi3cyl+2BK3mu0/kXMV/8YpHaZJrfXM9
dfHjhNuAV/qanzFkQPhQq+YMsDxdTJAlNNFw3pfjLQC+E/P5NNNSClDMrd9fuhQZw5p+yuNKuWfW
lihn6holWFHegQvw1TcGGFrGsfBT5hQ9oQCCLJTW7XKK/mW0sD5C57I2JSg2DMUx6iQhkxJn5fAS
l8fEgk9fSUFJre1jK82O1Y7/j8Fipp95brTWQneHjphCLroShVItuzuUPdVuG4JOvh7xhwjIBu9P
TvuRdWjzTJtVIcj1HCuRfC2G7BB6e8F/8n6Tre4psYHIys6uqpkq7GswYLTSAGmHo3hINUmUe00e
2VUSDlLjVnvaOAEReqBKZxUKKwpqJIdPtR4QlhE/Qz9WEiH3uFYMu3yPm42rYUZbimU6PHWteyug
9xgvbt18Zye6XJDgCvJryP429vRwN8pyICIcx05daDKK9m8yFzHYQ97w+cB6hcPY+ZXre5/dW4zd
YySuZXdbR4wwlsePQPoATZnSavBlduWoIy5feicZO6MoSbQOI/AOEIKBOWX0Gj9cl+aEaWLDedhz
MDHnrVz7ZZxOw2pjvWWqCACZShXikmyVfR08ufFa756cKbhM2/nO0BhxS0yLryKaOb4typnjARg6
6mmkFE5A0QnPWWC7eiy9d05VrIDem/M8kOBint1s5TjEbk44sgvcK+k5seNV/xApQZLliVW5JiY3
vR5zN6kp7z/BKqnBEMAX2DUTC4syQCAOFh20XrzbTUgcc9ZcoMIA34NpkHvrP1laTUvP6vOmglTz
us7xDakh1fNZk9KPJWc+zy+NO9WDsIhMsLyUF9zJXaGOb+0YgLlE7LlDSwXIHrhu4Cl1cI0hkLKX
NfG9dTYiO/qUjbw/8oW/Xlci50OoGEbc4m5rwbZigL2zWxmk8jAm1muwilCEsI8FOVHj/HNYFjD7
ZA4rcrnvXVwK2BDQXFevskfvjI51HSdUBVqTxO0r7XJ8s3OHD+nn+xRbOWGT1QvgIvh5vv8dF9ma
s6VsKNHDVoTQIKpRaas+ixcUIy1I3xSzBkgk0P6Ye9/AMB1tieaX62ShV/OupBhmkhKYkOT6mtGZ
JKhs5IAtoN6dsJvdps/+2nE5dx855uhC6o58tDuj8xsksHF4zMCOr19UzPNR/6NsKQiGML4FhPzX
1+YLltjZVBbqvrlXmQPF1xbHMZvNMt46Q1Ar7ZFSpwwquiwCpcvT+iFouNWifzUVr9AG/6vW8uyt
pg2L05oT8OGAcWSIsjQCYHAuy5iodpeD8cJsw6QlcbkXzaIYG/hw18XmEfwcfD989L8qzk167PsY
8/hjQ6EFeUEpWIlPeAif9s2pZflU0oev/uz8zi4ADhOcnHASLsXq5DM6BXyma2lEV6hEuvrmNP/y
FxIbkNgF7vI0+m1JYbDora7CcQkSFHa6rcZNGhAw7VrSjlZa/JT1V/qZ4Usckn+kKiIG0raa5BK2
JsWWTdOXa76o/1peDgxsUvPKnkouXqBZXNk0cbtnRvvHnCn3w97CRyGFKJkyve2X3HAP3RLzLanc
9OP1Ohnk1NDT2dkDdWID396u/j20z0lHlPPh/Uvzy4zgtKZjztrwzM60qNPeN2tDjdKJIjstMXLy
GTJsO55t90TLWEU2LS1nVDugZIzAGp/WbK8GogQKpbANlLA/4KzBT+aRYBrvYhJiYD7tu1PJOojc
H1FtdycieltlzogaI5tXvqNh4T411ohEvwM4rAsyAegqLY0A+l9T5n63/YAVuXfefUC+S5w9B/kz
ifnsg9LBQcFoANsw/MQEK0LU4d8v+fFk4YpaL45ddJP+DvtI8O89sxmg+3caXH78qH7H9vf2Qk1X
AChy57gW1XPI0MVS8qOoyZCGQXmjNRXkttySlQwWycZY/iNwYJwm4Zf34gT/vEPE8/29t+mWv2EW
G12E34x+DPAsLRn8Q1giT7yJuS0KHEmUCXRlNX1ZNd7PM3+j30c1zbuIHn+IeITlabCLufmjleLd
zHJbtWBD8QSppz/66YzJf54orStP/vFYZaLbATSZ+KvQSVaiC/LovMs58XkRwHyyNFwYaS2AvukU
GB2cgTTRMDCF++kl1O1LeDKWNocXc3kI+svQbEFtINqZbc55qoZMNlTBCOqgxcaYZGciW8Q360lt
YmX7933Nn4feA9DEWyviW6yN/+CwJQlrqp0qXkzHpGpC+dhDtJ2jv4OuizlkNwtK5412nHAWYMN8
4Uco8ziW4hxfvLjZR7z2J6tH6gaYrzqWL+KNNBOGduEVBH35VA4MMeZvSiNuw3c3jphgrWKpXXU9
Z3S939/hBD2PZBz3R/zsKmf4ZRqXZvCL08yFyiUcTD9/zVyaCBoh4V1VdVCmuzAJRcOJeaRy1muQ
F7d7wRd1IPGTLKcPhHfX+OwG7GHjYU90QHeK21S4bnea7xsiXoMoKu0u+YAbwjIeM+g0InafwkDr
lBHNgHCBr6etZAxpPWf+noNKpGMv3bLQEg6LAXAwEKNfdi2BPJ3ZBshsmI9aWPr6pzZ6i5SAXIaj
TgxlsD/afzQP4hDLS3iALhauFJuEnZIhe6R86/flAHBpZ4phDgsDdPQ7sAdBGW59HShvSmT0Gpyi
qWg/ph128TcC3459wp+1+2yhX2eW5HHvPkQIFTfK53nSEAEvBHE+Qs7Vosuigfw/2VlSJZoUPEjk
a8DA0/T5pWifKQv3+UnrAoumHQhV7QcYkTl3c8qiMREmqWno87/eNA3ZOqiQn1WlUT4n/PkedNhc
LACZrYlohCmpiwG7MMTjARSkxnwY+c+3LuYqV6tVOG20U7xzXUV4JYU8YNyDJSDo0WRwtRFj8mWd
wGq8lRMVRSPJxQlZfBc1H8LtG6wxsw4KSMt+4sLx9vojvALbxqkgkmf0ZBC+axmdHXI2amkr9d/s
VLqYy7/GJobE9XZ2x8p7Z2jgREOIWFnSMOP/DnM9105vKgabzNzU7FlFZ4AdOfbvH3NFKNmbqObJ
rO3p2WLvw8zsssjFdvWOghtiIDAlOVtN4hL2Ms1a5WaOn2tac2cb1hnpJlZCTL5R2mt4azHs5LIw
r05MRVTL/jNf2gqUmJCUUOkn/xIAOWZcrew9ZO+C8avdzkoGpu0gbDopC9KQMaeVqO7CeS7jwi1n
fZ2J27hRCc1xLXWaZcc0dP1NMHuoIQ2jmrQBIMLl9THMGvOsfvI3r88zhzbIRbBOJFPtU2vtXEft
U5u3xfy8411hPfvQEC7h9XaO26Y+IpRfzQtSycnn1P1JSSl6WeGXmSAwDSfT328C9X3IwW1mMQQH
xjIuLRwuKtEHQg7MLRwepLW1334dAYF+euhCs1F0rD7QULK3Bo/VFnMmCYvbomU8JbRR+jJzDcao
ecrGaCCeQC9EagU6c5siNz3UVcC+E4Gu7P3oxfMd0sPXwnkikXUxmVC9p1QHPp8F1/Ri0/vKinQc
U+T/QkExWZx5laBh4gGRlNcSGupK59gL2tkxFj+eELrEFe0QLX4WrusmcjaLI/lmm0lMEgBlKLQt
lSEn3qOAqnmSd39jiJF8OdjebjCxF4AWSJgFRDEvMhqNgAe00nRRsv2WZfKE182kyDgdsuXFdFQl
/Ut4wL2p/zm2f2+evkoXN3z4hZ8xMbLbYWvz007Uu/0W2E0VxY0T8Fwk/xR3dMWDZXrabqFxS876
tTVWp+N0Mqs1wxig4n3bk8yTMdNhQL/OFZ1AbYqSKE1ICwSvd8e0y7vhGO5SYgQeaim3JeKArSNN
u6VjphbbK3GxvopWmBhx8B8+PcEkDIgasjolh0n7Q7vhW0kMzXNAjwl8H0hFnedn+jLOK7QTgCKo
C0z4yyFjm3ORuvSNEji8OdQMG7YlxFoxoZuWyGHceMaqoTH0c0pFeNI2yj3TwiiyJ2yVvIyLsm0r
Pgs7IoO5iJSEdV4liYy8iLl0bhvoQwiaEfZHCglFJMMYJgV07UQfy8pltjNTBosEuNWS7MnvKMk8
FfRc1EEAklW1+XheHS50v9J0nrIKFsVQo+fnTSlaAnDWxmXCa/cYQ/mc6YVkfdZNHHTRufrbjFcl
NWdREgDcHHkTRxgYi7+5b0oX1pINawIhIFhWbZ293GXmtRlA3mD1XlX4F3k3hJHwnkaBzwU8WSdy
rDhGe9R6mH56OLeSSDaWQFyz2NyhYYpSpRCR90r2XshAy6ixoJg0MHlapSfIncbTUKYEkEMFFlgW
THkU5XAk8p+sgKNqQjiNcczlyQbJVOLNZse2e0a4P/qf6pagl9NGdUvFpDPVJo97aGmDNIQ3t/pw
RKAo8fQ5GnQhwoNYoI3XjA3bzDwgRyXUWvlPxmgT6fxw0Dd3yRIAFugw9BTuInpL/QAfO+CMzFX8
i9lGZ1lWy17AMgTsaqhlOh6QPSsFjb3gqAsYFjjvV54Uba6ViSVxGgHZfpiLY6HRIdHnfw3BxHPp
j0N+6ZOVrsKmi2+Zv/x7k3t2do3CofMEOwjZnF/1bRj9UyKn7z8Ap9ymCbWch6h49xFxbEBXQ+rb
Uid9X8AOEaG8kIcy94RDUcgQr5pvvB82G+hvJ2VtQrFSbjJPjCw3r3FaETwV+TMtV0hL9Wpuk/r2
18QGahr+QG2Jav/+TzvKDYIluRAPg2CXJTzWe7I9R38MDbzkkT+AKFGpk4m95EVJFR1CjvpkavGK
GB5hN4DVJGx7wyMBJM7JlUqeLFlw//48fWrSR4q7JeqAzfJ5k6POzWtto9dmKBoyU1kwRoD4nrXg
wjzdmuN/hi2PfSW7PpSLjP9wuCZJUExvMIqh6Lm0Gtu3dWdLZCC7Y4VrBOuZBBVX/lmFG7ZqtS12
iSdoqbDkc+kSemiGnFrPhjKGQgSk8y/jDOq0yYl0ZJiCIGE/DdUn/gVm68Z+IZ4Xtmnsmp/mGCHi
dusgbrV8T6BEzAH68MWs4gGB+DxsYiqbAQdrUYA0VgRBTr8o/mOYk1Fs/Dy58lex43+8MYqOFPxN
uhX9VxRtj1H6CeQ3vPkSOxBKU6gMNWsYdcN2dyVi4tg9UwehCLMlT6sOcvwe3yl6bUrU+ui6CtxA
tXZLOoiHwPtSsAO3DwxPMfx/gImPNIZJiSK+FOywFfWw0OXf4DdaHWaCcBHIHQU6H7cqnRRvAZFD
wvk84VrOGYql6U0BemeQpnfWV1JEMO+2WfGCaCCQAd6R+2LiDw7G/Yxsg9tqun71YaORRxB0CbKl
9DHYwqz2/xo0YRcBb+Wbl89Zku/uKbd/Nhbvy0rtvnNy5zujWJ74Fwno0TjiCm+yGL/Od8zRokOI
fEh6xQ3lYf+/NoWyI8aj376iAdfQtvt+EJuoroYScNPTnY1Ec40RZfCuecwrtUFfJffUmlOxQPzj
v4wEUuc4hRdS2Z5UBqo3/nYAUUjVJT8vtMU+0SqE+kjkL+JAhemOoK3d5v4e+hFOicff5fmKE2yQ
G9DNy7U/sRpehbBQDFUb0e2nyQDwFc2Vm/42+1AK2b1rA1z9bm3W+D6g0YsQuBUP1RhK424oTAez
sZ4O4wRcY3z/CpcKG2TCIpGZisjS9QuaRdZ4XsPALBeNZRIK1f2GKKrbTpKoawljMKcEtz5Aaq9R
9HF029JScWHcD1fap5UXpmldD+PrnuaVKl+CaPFwBqYjn1r1uIyOj3LRCaT7uaVtJtUk8mLK73SH
ZjJLdGdKcLOhi8lKZpfi6fNV5SMj4C8fcfyYecC23KNpfnzH9J5i8FsdTUzrR4GGHI84f6fPCmIa
KV9r21/I/TsSE664j7aTcbx2z9JhggClnmd6VpueI/Xp5ADQYU/sV9jvC9OKSOXCEQ8aB1qagcF6
hovyS2K+t7zfX0fIYlzYreb/mWJTYIa9UdxArEgEv39skE8JHi1qgaB7rt6Cq2kM4ZZaKcD/nVI9
01dBUfiXUevjZvD4ZpZ1PBUC9sWuNVQunPAAgbFqoQDRMfntcSXFRBWresIwK2Mw4zCpq/Stm0us
3TpwSeCI1jM/+lk0CRNeq3HPZDS8jglvtjr9Oren0/W5Py0u91FkAuRcsmil5iybrGJh/F5Xon2M
TZUcpbRx6L7Cdg3NjsBt4Ca93afFBLeA335xAEgITv1RHzzFK7xkEyCE6SVzNMU2T48KsqdFyh2P
RQB6fj/lXJPSTWRIVUogMT1yGHjdfJjerlZJbNgWDOXi8x9PApOA54wJ3OwmTcxwsvtoEf9Ur95f
CGmQsewDq8qvPiKwgZ7rS2LNUhIVdexrNQnDdiobVYIMrDiJ9MBKrgma1paBXMwHWHiqFFRWP6cp
cHbgWIZ8P6KAfpoYiVMf9xowT3WdH4zv6iEf1DlnxEgnqZYslFVe+kcMKt3cXwSh0aqZcqTUe7zC
DKSmWNEETGJOxZDwtFu0+UG1Xrclbp6zUmqIFyq8VuZfKfXpzOJ4QRZFjayHFVyU2wZtZW6mS5NR
ei1qd0W2OLmMYlYGkaeqw2ZxAxMcoS0vHqHXnS4LSmAByHXIL/fgJmxlfXkMBULKzodCCx2YBWjC
Ac3cxDgJW7pfAJ53NGEIQdazrf0B93aBlZAV7jzCpJlhF4Bfe6qZZnrvc+42jwGZrhPl9L/vAL2W
rZ1+sZg9uj1yapg37E4jz9mxksSr7uysw6++Dz/R3DC4h9Z6yt1iBvgnfFzYBfHD7VSuQ263AEcg
lxT1rryuOZf7kY0ev9q9/3RsmdNRElV0rzyvmEV7y59QhFf7N3nRyHGZ/PoshJyllSUcq7ntdPtW
0IguUHCZaGR1I4Mnxt4v4VAy1XKUs0lr3D8p24iQasZIJNOpyeenzXaHEsyoWKBAGDQUrQ5leU9a
G8bOWi3ZBw8dVLnoLRoVpJro7Uxql15Jb1rjhzKU1gLcuBOvLZjq2JJFduoNwe5P1p6FoD4JQf3v
SvwWAwl0FTiXGoqE3r5k4C3FPTwizp4VbM45ehBt31cFi7VHKMPOmAltR1OFYxs6wBYF1VnQ2mwU
xEegVxNJuJU2wAamwUfQZSF3KoolvSrQaEhYEl/+kAjkZEMXNCNhfhQOTxgSD9G0uSC0QWhetxMi
Yv9TFjX8hFaImvVs+G5aYO3lwhRBmuLru8nX/DB65sxinav8vFrlev6eD6f8hYehjQVqs8yQKJzv
I6prAxFkY9OPY0W0baPCJ9CDmr4jUy7nBTnFK89ZkacW+feJ0rvA9ZEvfL3eHXP1AqOJFtbTLPfn
+rKhm5+GNiVPHwzqubMWOZ4ltGocGiZjNnuUvAXb/CC+Fj3XVDUeHCWxrCyBPp0jcTWEo7VgrVFE
gWyRgfwXZUT9C7U99tdCk+xKibPCvDHyev0NgfQG3mSGKX3iPfsbnQ7WQek2GiEAXij6PULDDF1r
faLSM3p+Y2L5kpUiEpQ7sLSFcqW8bjnTYky25o61r8FGv+g+X2Hig9h0k/n+NPprB3wy7hRvWDQS
2gikomnu72J1C1bvMfykEqpC5ifuENbmg1Dh7muBahpn3F6dgngoM/95ijef528U6tRhmFY2WOAQ
jmR/05Md9Ypyg51C8Dq4sMHnmbzydxK4HWbDZa9KoTY8dhf6nYMLNWshzAlEKXAt3wGY0TLA/etV
8ffefIHvM1F/UdLklvKvr+W7IXfRYlUgJlT5Gs8qswPMnz/cwVkpVqKjtiMjnPBcxt+haYd//aqG
0ST9ijSwwYeM0tjiMh/ts1iApT9bNHoHCg/bmF3lx4Cuh3Hx0TvLLPNQV9choBv9wb9TwWtKhl/X
r2pPwZrKMMMrWRb3BUvMZu4kennNHXiNO+vIVuh1VvLLCHJ0x5dvAqUvKUYrOXg2Ykf+qJhEQQdu
kEHfo1tQKOpUlVYQ8kHa8hs0Z9mwOdVV5zyAW5UPrEpax7QydwCMdDiiWrRU1RKiuO0d8MWBXvYg
gDtvAbevSOkcED/PNWsqCnO698hpjpA9DmaJI8l2wZ63/dn+W5hLUOXgff4pZ9Q8zp09SMzA00JD
OlKRQGouL4bl5KbPlhZiDpj/CDW5tfv8Oe8EW2YaB8E3RZXNy52zVKDQN+qSpcr24f35W1cNoQe5
0GqBEtES8Zh8Y3Pzxy7QiUkXmsuJiZ8YfXa9G86UdntNb63Q2+lgOBopjgxLycIP4DwvdIY8F+YT
n3+PaDvG9DHHHLm5Kz7lGWCOvtm4rXB2UzGddSv5enTr0UJpysSEXh0cykuMiJvxW77Q3tTUIE+n
QXOQHE6oJhFV1WaMGRs2ub/fThyUEKw5EqcbI2KSoBBq29SG7cc7tYb+8XlLX1QcPkUWG+YQCs4Z
9peL6f0KONZjCDUGvfNku13laJAR1PpdnYaINQXIFWAJWQ9KKYBzgF/BwtNWpdjm7aoqonrYYbKT
3ahSY6fM8OzJjK0UW/frLCCTiykL7Qq0FUtqDfvEbNIVU5WuLVxuOCwTD4Zvo/O2ctBj+hzKtOMZ
8XZQsva+AmZNz8m4sGIMWT8C2jHF+B1Vkm3Ff4XIWVlbz4hLIX1yUXF3j3g7ufmZgLF0ZuWrREnJ
ikZbZbjk/+NJ74IVu60yX97p1i+K48zEszPr+8Uv6CxnLCHosCd0mc5Za1q/kyvsXNNO6O+14lSo
LryFPXGMzje6TKbIZAvvJNfoIg8oA3jIfY4gXT3ocwwC3HWI+yDv16e8qaw/0eN/m9VEkRqC5+Pw
lAK3CRDYsepa1ca+Z/dvuMh3LISZRLonXLV/mPg1IrhhKnNQxBVtWIlBnhcZrciUxS7vG1Axt1hG
+mTXpnpCAyHoO1DwXC21ecGnELoB1SEyPAliONPxkcFbWgLbRypjakovVIs43pddOlzwoHlSmTjG
QTnESGnLLo6DCm0o0QQE30k7YKEzzOAze+gx8wT3pR8U2d4xibiiZ540Z7en4noo8fc2mqDMo4ww
NwxKPkB/fGJA7P6SGWKZjbmB5fFejL2qCsLKQkP6AJEbxBnyYyJYZkOTGsJiQqDPC/t2d1e6/r1a
KuQ9LxjB2pFVcus1ZOi46atAAIUdBKGWKFpxi824AV7iOYJ5p87IF18EC2hrHL5IkXaxZIMEKgBs
/+oGG2fpJhk5yEjUKM7UOq9idUWrLtmvAUznK93GKjGDRNuAXPylGE63wyJQwOi4B1oEgyc8MAyn
vfl00vQoJGy/jVvma2+tq6pyXXHo3zc9kq8+h61kwZzuqWnazo6xOEVLIiOg/gXEh1i6QWpfO/Cu
5lyE2qRCBrR3JKDUSSv/rUGVCj+ciZbTGHUjZkUEsEqDpscbnoPSn9JOSzhhkBBR8oqSpW+lZDPG
L2/vJcEePcj4m8aIxZPyTeFNYgF7+Q01QjnnVVhCmcar+/TU17iKlgDscmnrayZWZNUpIKqY+1h3
pIcWLO7XZXHtHmFG2+aYKlD/jGRp3JRM82zPJiN5uQbuaLi0V+ACO+jRHI3dTVYOCAUem7TFS8Pw
44vcXzigHj5oBwcxciUgaepNSxkz3ti5oz3eUAwzmtQiccfxN0UQjGrwPbY4voSomK1CKONaLSUs
9Kep6Fp1nK7OWV3kwigHS+kiY0Ey/bonBpjRBr3OL2Htol4dBFokwrXKI7+RN3HpUkqptznxQqPP
0t3cTdGmJ/bGOXAet/3kfeSlRfe6rL0f72kS54d5LUIU4D/FEo79v6ii9rUroWHZwZ8KssStlCHO
TTahujXvDFupROJyRol3RDM44m23oCHvL4rkHWyQP0Mr7MC5zCZdxai7UGhyTU8oh4gu/wht0/Jv
DT1NPaDCGwTE/6vrvbsVYfVm4kg+IwM7w1DEAfBZyG0nd3j0SZp7xY/K8oixNI+edggOL40YreUX
vvmfa0xOudDfYoakJX4LcET7Kh74u1TlSbQKmety4FUP8gBbe0kMlm7Bly4guWenrlEpiXgDdjf+
mheGqZmQJPNAMTngUsu7Xa+DSpfCg4OuBlybSlg9Q0cKVrz+gA5Aty97QOTaLmZbI1NsKye2artF
Bh8AI3uIyWKjrDUd1mYzolM5vVNpofgIJGieAfxdhzF6vidYuzaZy5IgdzLw+A5OzA0x++0Qh7OW
Oqxsv7gIwDhvEiq9bWTdV3dJrfA/RL5cpjTc3UcVmdtYZkEX1gYm63RidBpxO6x9V9Y2CXnf4LMN
pqopjTBWn1Au1Hakw5+yOBve0QDyCYkLuB7d2SA4GyVR2PcH4ho+8ZN6gMjzBP5roMrTDkHPOX7U
G4lEEgQcYmZAME51Jc7Kor4L7RIXOPhMY3vs7zP0l39wpp/0LFSqP0sfS/1AZWUlb+nUrx4kNJVs
QqHzg/3t9Bb7dmQzjO0dqx+2jFP5FaBqcn3bTNjMSmyKEt23dMs17P9E0HLrs/Kfhl+0V8jsN2eG
ukZnpmQnnLAI6c9WfU5AuKCt9cVXSRKmzUfHKqXhd1ywCPgivMlD6trr0M/FUmx7j5zG9Bk4laYl
kGxj7nMrF9l1u15JlaBLlWOEmBMcLu2zvnqavS/A1GCMJZL2tbldLLxzBt93k+2/Q2k7DI5PdVPL
X5U7nCar8T+dR5KPFU78MKDcU0TE4ka3iSZD6csCIvhf+Iwy2pBETJNesIQEUXePp+VB/hQmiXfy
g6KDbGe7qQE2f+XEyAqBaWBsJroVD/ZpoSRIxnRUn29Vaeztaq6rF1kXlEC+taTJm1IruzmoyXn+
uCH8kuyWG6+lT/HCBEUB5JYOHdFnlo4usbGet2rpT7kRwXDa0G7a2GlP4JNQDPY0Bdyk0KD1BJ7K
Uj7BvoB2cZCaHUGOGo4kki6Q+AvELgEBGcTFPhSZQo/jSPSt93tCIwrttK4/a78wWztoQXI8DNt9
H3ioxSUzK3j59/PTMMUcF6r8UBEMJ94J8llNL8eNvAw9c7nECPs5rbBJXBJzh2dVkw+RH0MqmNBe
qyZb4+wrPpcH427gt1appJYDTgvzAfMNdQum9zGy8Jf/auqcoApNBI6fN9waDYydIR+u7qKumiIS
A571V0BDbUN60ghY8rHMD3inKISTdUBw6rDaI+XuIK9rjJN5JOJV5xGoSCgwwiQ7XZhhfpYftcze
N3G8046Q+xC8buzxX+ElYv4P4LuAvhJLtBVmT3rcYMChShS54/tk0aO6xXt4ORTHiJXHNaIEDx5h
4XRjNf+GhPdradXy6DvVyeaBTqgTn9NF6MlKb3ChK7WR0aFRRiBfMa61QnoVbURTvOO1FN6r3orq
XLIMC0XSx6q8PRQgjarQKRlqJ5Wwsr72hA7GnSwDTY9wFY3JnHETx8wNJfSj9My9M4k9YG2yr679
DeeiLTsYqT2pufFioCTaMNhZNonjHm8uc6izluPIpb82QRAvToeMXsUvV3riJXXaK8Eve876OMlR
wMfME5BvuI3V0MtBE4TCFV1SJelaHweHb6PZIcqUGnNNEqyOzq0Jqb9to33u+8ickqRcY/E9ZqUm
qb5BPTrxsFgpLH9pA8xg+j0Ey8RYnEWdVzCM7EBxaDXn8EhjpaG8H0GUgGtbmNE60dYktNI2Q/3l
DGiMy8hO3jzeEZKWbrCztmx5eeWfwGZ5ONs2PSTXo++t0FAaPAXGm4oxDDuwnlI5obpPLccmlUmM
3GfMd1edzWHHRu95M0f6DoHoegBwqLSCijogTr5lH3PJQC/+wSOg+BEEB3eaZ671Mf0DB3Mp/lpQ
JTsRsel0laOQLsXJ2haDb9YXLGG4SxYJejbOUHy4TZAxen/wI/zE23ezmLUlmR2Yt7DE+PjneyBh
fslt+7G0uQPA+vCRxUiFV3QmYE5ZX8mr7+hmQtx+DqdBJrV7SpFD/y3sOy8kEd7O37zeKBh3pJz4
cTJifez7yj8Vp3zRW76g3GUXoTyUBFEsIOm5450sMr67qZV/6Xr0OoMoQPszzO2Z+fghP/aChyW7
+MuJzDhk+oU45LuN8hJrUcQEjW4VsdQMGpSsUfwwXHteMguYywdKaBRsIsOvo0KRvsVKFy6hzOdH
eOmJd6HQDQqT5xa/tF1s5xlpmxJeuL2G/ta8qaQZ4VjXs/p3KRdQ0qgMjsUPd9I7ei0vL2SGm8A2
+KlHtPDiU3JUU4AqD1x7LpGOWptl2uvM+Et17nPemq4D0eF+daqY5u5lboKTbVqhYtoSDy2me/h0
H7Bb4IVB4HIJXqSWao/04aauetwxxTJZSN0bBnf1jiQ2ql8LNV7O3IdPsPr4Cy1d8IvWpHYLshlI
VYqTvQCRZZfZPK+ww82mg1oA80tT4ZdoSF072AndR2l2sa/VZIS3IZ2eaHR3zy3Q+EO7+TKmuaMO
BgRERCWB9pNT1bsYGsfWkQ4d7Zg43frCWsAn6an+Zn0LzFctqDj9COMpOiVlJ8aeY9atSRvWJ63C
PSDF89mTI1YZNvuwVZJIxowcH3TO6Kiq4sCpfiuOwEr+P1UDc38iYSBG5Fi2eeDHMTz/1gahIt8O
AJJoSIQpMZ68MFDPBo/apfNNPI7FXWqEhIUs4vVBXrwpJOPtaOCFdrcPrr2IhQigQTQJNuvJJUr4
dUdSJPSwKTbPbYoTS8zAU3xE5xXf+97GWzx7Z1JGXc1yCNXYoDFrpd5MhOFvnIIDCPpBR90kfcSW
2kaB56oQDta30aFXwUFm2SrI7xP1SoDT5MRbVPc2xOiwbar5cn6o+M8f23zqcH4Esu3bZgA9vjJ4
/4f+DJi0pcg7ZPe7P5OYJQR2VWgLimzIm9sjgL0VWBnNcBpvwZK5IIujmvEd9xRchPNvzutze1O5
I6khIfj9a2WNXMQmwby3V71KUd4SR9AvwsPc0R9sTLKa8bCSp9ZbKmf+BFG59+XgUS1m4SsXsO2O
kHwn63pbQw/4r+Rfm3+N/MXPbOF2+OBN+evB1URdnQu2kElwWIP58ht6himMA62M36hFiyHOnCXG
71JtM9BkB48Ry8lDP2iGZaWh4kVrUMFNqFuDS1jRhKm7dvWtXCZwbZ84Btpsu6c/t2N2sPXvsFYY
FCJ8ep295/mNlgG/u2s5gzfawJTIQLLhfucJUXTfA03yVJY0HHtyQQ4NEVUX0MVO5Lh1oKLDMm1J
uAaDioqjDUy5xJqLSLtynDEhFF46cZGImzc7trqQqRaJ2kZuDjFHwfyJWKNtIW3/QHBB31u8YgI+
gNRWZvvosAWQwQfVhlvBXfliXIwJtlvtxNM/sdVpmwiHUytU116cERAeSJB6R2HoSLg4Wdq2zSFv
rcIX2cYLTw1eI9r/fXL/fwk3SW+fc1GCLRTIVIjTtaKtjnKRZ6S7mmlDv72UTnEBZAXwpB7aaI88
plVynbUkRbVb/Ch/JSQRr0ma7aZukyXjVDd8HOhPDE1Igzz/No9L5GoA5I/bIObaJWNOnlDKZGJp
tJzlIhHOKCavfbq5nqDKTT6losohyy6f6cHrRMfqIMRQCf1I7LlRcbL+FyESb61QxQh0J6A0jslb
HvOV2gCZ/PQzxqLYRJg0yBydZng4E27ho5JQksqc8/RgYGt2RZbAW2AOa4pIh4ylz8DCsrN4L1rZ
OuqX8Ak/MNmBdYk/oC33aPEsqYRczyC1keWzLDRaoMOPATzgiuDuaVtDfGxvokSA6SXb9PTyMscE
wT+a6rSzdX8T8Ui3fMr+BKkZuTGhIi1S0zqPKhEY7ckq2PkrYhlS690nD87dRaAX2JUIJb56NebA
9zV2AJrszzBZGki1Ly7Vmcmuip0a3EUZmenBqFKThB80UwuB+0Br5ACIK5Q/F98JEd4JSNAKVbSZ
cVqQnfV2RyMThwpv9KJ4qStWakXHnwjP8DGBX424J/zgyLBnftqDpZjpb73dDU/XWJ3MbMe3ajmE
50PuLs7gOQh3gAx15eib8UWkgoukeWfbCC49gbvHCCPno+yzmFM0TugJIf5N++k+0or61NOwOp7w
+G9fUWY2YwSRfTKsyWe25Yz+D9famLjek/UlpozkWRY5/keJ6e5dNQKNAVv3PcH6Cpf05MHEnfsr
I321y2xbpMJdOzlXgsXqwtestZQmS6VpxapCjEl9DdHNgNX8u0De+ttuhB4kSkfkpB1aLjrzdnAg
piBbvo6L9TsJZVDKFQeedmwRKJt+rChTb4kRkeoiL8C3J7v0FNVtQBoAuPLqTrGZulohy9P012Kj
rYQbZbrpq1P7UIuaRbXMM9AieqBqDKhDZGJFozXnmq5kTb78m0nQzwUTLkqeGbcxxqouRADat3vU
cPw1m+49VWZo1oNOjOdCLJtNWMKjDHoCwFYuWia1mYLOlR3SNV9788lGtRl/ULDVKz1evYumQTgb
yWJB0X9DjGZdxseUixFRkPW8vgZSqGEUndu5SnRpjLhPtoC2h3fmrzTdVOl0w/SjdOYmEN0Lo089
7491pMRZkraKmGCXNtHyZGC4zQJ5S9sbv2gsnIaPZ6hlI5yjArFHn/V/tjtZ7eenTEQS7waEdu8L
hR6ZAUWonoIPNEKs+q8JN/EQ54pMcfrnTn3RLPJsPrAtXZgOjrPh0Mxszd61d4cKahsTyQB75PY6
PRtcSLPApyYdkgJ+xBGj8RIxhI3YiSXu/kqRL01M24ht4/CJOd2g4FjQWG/EzQA8ILQjyTs5pzVu
0UyXru1yuWnS49mi1g7EKPAtdvhXKyjZtDUmecm02mhmLuztG2lsFKILA6pS0p8m5P3KVOjKvE8Q
HiUD1cwV4E/4TGmJxZw/4u5ZF+12kH0op2Nj+kKjS+7XerqKSWcMCZ8fJj2t4Vpj51BTy7l7onEG
FDkEJx1sVFXr88YniJccojTB948BgD6Rhn0X7MF6keNrhF1vzoItPlNcrkWEtnwz5RMtiZCA9XPY
7D92XpsuWM/NJLOxbERqppctQUUQme0q2F5K3k1MtQ6hr2EEssJ8+1MBxA/hi+5Rjg+d5kxXBgN/
MxF6f1suDW+RF9s7Q0NibcjH+Negl8/VBWBk9bd7UdVdvrYTVntmQeNc6gjCafrQ83JExnmQ+P4Z
1DfNUIzVcZ3H6g7SuX513h4NQFLprRc2KF6QoMRaiDYKXyolSrTwubZNfWRuPA7dKF0vbVK+eBaJ
YkUSuDgFI8PbjEAyBpxq4I18wAchUZujcBoOkK3rP0baQM/RM8XPQCiJ/VKNIlORGAbZK2CzhFyx
/7u75EoUe3Y+CJY9jf/KEJnLDqHolikozPPg+0OSkphQg60HOKLd/umFvRFatB7iFcewDwZDgRQp
PiErjP2VzlPFA24HBzoRol67MEPZ5m+eOkKH1cepjoJ+AC8RFJdACPobVXLelMAqQ8pECswEKDI+
rRWBVvV9MA90ino8Twwpflc6bc8rO7cUuxjcwIGP0vdywZJLOGhvpgrn60m1dvUgEaUiCSBZ0Iox
DNi5lLy9efnRA7xsltvWQSR5kGbDk7ZN+dMUvaOohH0qAt5Pg+1UUDsr3l0KEuDHksa9yDaEjpm2
wLy4uDyULhK3ltyAjon8AGi8mdw6EDacLvuseD3jfpGcKOe6BZOG6eSXnDvKF2V3sMk7XmWyXEf4
6BXJm1YmRE0XXhjAodMQ9oO9W2NiJ1ct+XlX+sdPDW/KQiuNG51iMuwj9Z9sfvczQDQ4RKn6wD2O
A2/1zrLCTmsWdgZ7/rWVTOdUV5zahOPJbGfuxnaehQzOYusX6SIquCOZqWOQjbMm9tbSzJJkkWb7
YxUy/boxDFQbhOnbDg39kjtBfVEL1uuQfXkp5OtclxITOXWuJuLHHw2jb3oTppeBx+QZsQOFQFAN
asrePvQ+8SBlq3b/WrtstSOXQuex6Y55SxEZElyX5rvxzz73fjtIcGbHt4hHhJXUsBbye6IvXP77
KvNwlT4hrEaKNvqZaKYIxUO/0fRb6c0ldxaDkeLqgxmISssSe/a/Rg98cKSfF1JT0tZR/SPqJ71o
mFUYHs6lV6mkkvoGy0M00pdVg29tu8cMDTklFbpkVJjJ86WDt9dx9mI2HB6/SET7/ZR2JEI8z0wt
+CYboQMAwkGLeJgvZdqy/vslMBFmXrw80OFG54gDOd29WiIAvasRq4Dd3L7mL9OwMwXTnrq9YKSo
L5mV9yOyXQoF1EnAn/zADbAmppjwxbOh1rrgasxQ1ctqMeFgDKZnOdWREJf+sOtfcpWnRUswGTwW
UxvbJkcwiWAj4cSnVWrCK6QvmP9u7aeAYMNHS892z9k1bv4xXkpzc1ESbOpZxeN+Vm6FkxmUGR9U
JuzbUJpXkKHPjrGkyhwS8o4HSW3Q9QT3QqtCyaX80FQHkm7wtSpOYV6GeNyraaOgPXbP2w1bWHBl
DbqzSHW2lt17gqBYBbMEUEccGuWgn3CpQkePIy0rBjsNGh+DfwnwTah4brn4/saEtswB1FHvFPsm
AsJrN+XnmBqBtkTjtiE1XJKJyLG1nxgIX089hJ0rbycY/hV1reGxzwn4yVlCdNL/wwZGZzY1uB5V
Vf8feNmnlCj9kzBJ8kA7xxDCCMXk9kU2+ZZLtNKUrZGcPb8+higiCr6ZJnqqbscHWy++DwIrgIHq
7MteFKpEBY1M/iSNyPf94MBU/hfW8YB+bviVlB+zKXorH+vWB7sTLBL8ARMPfXxG5JE7S6b6F/2P
f/o9wf1+5jO7vEbrdco7Uww+1RJA/qqx6s76QcQ7Ser98LM4AxjyBDQhfQMUPIITOertYu7ydA51
tHkoQ3cH7xBpTaaEN0S3VhnmKt+t0XqygjZfC1xHegGa3CKRNp1Gh6PSIMKCebEplsLKrX6RBDED
RJboopEYCGdGGDdNx8VzzQ+Qm4ZV3ssM5OgXoTy60Q1uOPLmTFwWsNduPlZAgnKWy3F/RXz3a/Oi
NRsoQdMnk6sOrYp9jHYc+2XqiOOfX90qA8YbHc+u87bXv6i1FwMaBIQJbWXfHn6+QYMbOOsxSJ45
P5qOZgtsWot7NIVTmAEEpNXFuPkW4imgCPMCQkbt0JERzCP3kvVjvVim9p34PbnJdpS7eJLgQ5kS
rMt5txO7TSFXBiVdcor+tVll8Qo3YUZe2ib/yL+Zrm0IpkPnhhEydcXLRG24NfB2PXFA4fcT5KBN
lN6VhfWgOEdjAT67+yEexCp4sQMcEsVSeXbTJBlTa98zqOoh0WPUR7vzxBT8oTgjqPUOpDeGC+bb
7gQ1jKWBvLB/QUVM3BeN9jcmPA7psQbR/jpC9JiagdL9tt1Mz8G/I7s4xHfj7Ovmx4gyvafGy39I
aA3mjOjPMsdDhkOYGIEarkisNhUIPbgS7p0pFOUmr6OjGzPYlw4T6WqiY38szmu3EAJjt18sM041
OOzdFjz/X7zfQPxclttQW0rpvZv3H0m48PLaQu1/9pS4nvvlFjRWjh2twyRAxqzl+bn+2twdlsgL
7PJdeoBN6gqEsW293K6rudfEEe0CzmzuHix3x5vYJOg/lKo6WjLRvRrngucXyKT3wT78iUMWv0Xa
HS80rYVBshy5WQ3ixRowgfN7DfjFaOZY3fT3ieiCbpHnwKES8SzYMxpi+ysf3yG3CpTFLZVGK6fb
+x4MVneFE59N7lTIeCXTzGF3pNSQX2rTYtAB3oEzh4KtSgz48NuqntZ2Qp4Fgk1v1ttJYuR6yBB1
j8e5WTTnFxHueC7AMqZynSuMhDgaIsmN5gvDj/mbbkOs+xEsHFwJNlClqdOYwbih/f/sm0Xz6mNA
CnLzfosc0a4DhQw3w1v/3S3bgk5qMkFPPX+RiYj6fN2zyIwViS4zxQkDNkc9LwtaK7JZZ3rRnlQi
75IYgcj8rI2OchYxzqMl/bqrLEoKMzhuT88fd+vBTI9nrx5FMlYn08GGPGxwZ7dCvZYsqJWka0G9
CgPuWkP59Z4RUkOPPZt6HEYTgmYKZNfKLASn3g8YS7htgEzM8dVTxJhew4Bxt1OmiBKxyomYjnWh
dtsSrPwKKW1KUcNwuqgDAhRWiT752+sfth5A4R2jlGO3rz+g4CZPr1CrendU1/Cd9XG3JToBa0tb
qedUAAKe5oKoMeoQZ32PA2e+WR7WPwCmA/c5Q0d3q/PDWgmKPFUCeAo+NtjbA1agxDuLw9efKwbe
JPCRS/nRWB5f7DP2KYfSjhCZdTz3ImGRMSYAz6fs5ifoOh16jAcHvhvpGV8AKud3eOe125aaGJbH
cop0+dMVdv5E6x/Mepx6OLntl+jmfzsYfV/Vk/i1bbCkvj3HlP6dZp4ykjEE/TmZEq/X3ZtcVj+p
ENlAjdoiaiV5AI5jwyzjWwZjwhB3Tof9WHY6wFETvvgT5hID7Arttub5pbPHB+MSwA49qy6RK4dA
yz9fglgzH2dOpA+0Szn0EI9iDqtwRIRx5gQ/VgXWwl7xHEwcjWF9XiF4NS9m+TVOrmJkzkarWqyN
Ms5nSOpJAGRttx0gIgomHZ8U4Oo2zglvMwel0B2gdqCce+RFkcCtttrJIA+tmJNmSWMGraMCzjeJ
E0p4gmguGLS01pRi9pJhr1J9hITjfnXaOz5/Erv4mqyFXK4aoJONUk075BHPOQChR8ISGmADOCLR
E692WheAZC0DTxVVKPZPodn+CGo0ZRSP7nbNqXgPhwhC8l10FYT7Zbfz7hMI0rU9MVbgdfxP8DZI
yTzt753WNXfR8LAmwHvhoJBEp5Tky8qudI94PPzfOzzUb8yTAUldJ+W2itK4WhI7SqyhhX4lQKLg
JvGOEiplN3bS1y1TkwkYoBbGCVAV+3q0MCzadyw54A51vsigAbOorTgbp1za/Phovw+EH5LNpQ/c
Zgj1166asBvdBXgP+JUJWGnHK4HWqlSNPj+zyiPWgN48zpzpU/J5thtzmNZa3AuwEnE2Iw2RWD29
y7AGoGWgjdjYwQLxUKya2LUgMbzSOgEUIrbRXe0llJx5HZR/NjuHKPf9ouEgCdJR29DpJ3KaqFkz
PmOPtMcCw6BTd76ufvT5Ws/ZKCQvUxnv8DZ0SQQNN55eZ+G0aprdM79LjVUu6YWadYM04itTy2YL
bkFWyYKdTMX94VrtxY8YkY6/ux2TTrlFIJu/Xe3NElN+DdRoeQhiGRuEfI4dy92hCYSCcCyd9HY7
mLQog5089C4VdoS0ulS7L19ifakYhK05YYP/TOJqYqeU0+A3UTv3A92n53KjDEPvfRHBtdJUEav3
MEuiIGL9npkZZyIv23NGaFjNOCL2c5ZATTk8yG0LC5ChwKpYJHZGj1i6HOZ1ZxrAICWy/V7sHZU4
Nk7XflHuplK661WiOPbfs/tGn/NDJYK93quEByoL6yfp543wJOLTqdVJivy8aBnh2nOYGTv1FPef
oZOQXsf1F+ziRmhaTXrRlaNY5LpM8mNiZJBZ5ZZ1xFHFkeWjWY1vtgA7Azjg0A3G6qwXuSs5uEvB
r2/HQkPFn+2Yc9ciK+jUiRurYCTWV3e4AkFYvQ5/oDvZhlBvfoWGYxEuLRETSMumdlIq7g5jqsu3
XLtC7c3Pwfo6nszQ0WUhPHKciEgVad53RLSnLiO4E95kkNBVqAVcIZxYmEAXmwdj9pG+OAiFmwRs
eJMYG8wp/omyd3ECt/yknv5tDt0EsTsU8ne8WqB0+jFMRb/1Z8l8dIDOQanC1b9JsY2bFYYZc5SA
RwfcE7YxwEMJWSwTNwazJ62oUfoKNUAhiRtm+HegP8/rbqCeeK0kr4E0ZDNy9o2tV4YmlBagLG4e
WC+FTAn7us0NLlcZpiNx4/TUH9Tbd0NkuPxAt3hpzCoFVVZE9sISNsOFJU1tUhDIVEVmQNC5LY6Z
LkkORq9I9YoHkATjFJ8VEx8X3mA380oKugDqDfhKHHqwFc9o76XqlIAtX62waf773vR2PagT3Fjh
COCKY9UAcykOuzu5a7pMLjTaIdEV4VD6oRTitIA1Y8I4PIAdw3crR2ZiFtAcprWkfeZehPWf77nC
3EpvCF3BS4+zDlyw/6SNYUTUdDpcCvpnz6bc6DlUaY1LQKvyJY3kh/T7ShgGQRQWK5zCuZgsG77d
hkw0XU02XL7Fi/ANj08npBAQXs4x40BAszVRPKCfn1iAtl81KaVlvMqoNogY9pODx5hinfed4wL/
RhTx4x4Io16FnSUgMvvPWrZNmuyTCYKby0nlvpVof+oCISfUlQY1lgtM8umQHw4GpXIxj6zNbxA0
D9D5UxglCGMZtvYaBjE1Ot5PMkYCVFv7kMYPeEExmNB++71vuinR1c1C7fEkgxsM3T2UoD8k4zsA
It5G9ypu/3UKddRiXTcANXuEcAhJr4zeX5C/Ka5VyjPzK5uAmRTFq4Vu6jMEDvb1DyIt/8/s0XJM
3gUJ933oa+sCqrQuODv1RaGUT7Vrtmvz0APcXz0TDJFWqtqNGfW3bSWvHhaka49CrjraspbEhbis
zOIx4MrLGOK1fAoPTkKyWEb30leGja1urlOkgaK3tt00Yeh3mjjDX3LtF1waQrZlzW4sJ91iZR4Z
Zv+NWPL3Smsfh/ohLC+TLMikN6RQq8GxBlT+fQcnUIbtjY4SvQJo5ItEAqcWSux+SyciHTSnOC+n
NZKJtFtldUE5h+FROYyl3XC3CEOrgjVhauIS0BV0Z0cq/f2ZLGkaj9VgmqITGc3UPCrqh9JDy9Qt
cNWxylO80aj3N+y0geRcTTNca22d+D2e/oGc0P46fgSkzG4zaAYHr2yM23MMVhm6eDUlU35Ohsyq
whBGTav6XP+9y/uc+VfLcowJjqlJkNYIhGQdI7fDoD9LUa3BY9ohnjBfNGz+n8t7e12zMXt3BMm5
tagA8fBfLc69V87y3lva99IAykDbizNO3SmmOgAUImnlcBXY/J9TpUkncVUNXd7YwPQ57cqgm8Su
0IYTW7O/LnNgf6c4aWm1XvWAc1mICuxw19W2eO/WQcTv7tWOMmgT9FBg/Aoc/SuvQ6JNAnSv/q6l
mbhetLxeIiLoOr1wzr1fs+0X0GlPVSPveLU0PmtOWEMz8/BrSW91y2XKXQ+j8pc5tbkauEnyqG5d
goJxAOxRHs2PcacENv9rIQ4TDI5wYCLKJTnD+Pgr8ti4TD/tT0F5pKXbCgBZ8gkHHFjH3QmaHDvT
QO8vj4V8UDT5NXF1BBEQfjwpVaRaeEpaZzxHfe3bq1AUS/pMDSgtvV0z7u/1NKPJFvwKbjC1ZZ0W
/4Ftyc1qIoSiHv8HYITxyiP/unGZGdaTJ8UZTBxD8TYI4395KpR5BQD0D6f4GOxX02p0crFZlkbz
++DLkmQbw4WVFxaGND+GJ9ouuErRpYbuydL2R77P+vKHoIscwCyxXccw5jqkswpwbEtIdVzzDkDx
regEjCLI8dAmYD8FohVZoss3aXfj/Pz6ZMIYx7R1y7WuJ0LP2iPZ4DNdbSTNGMotV/AQjWnRNFAS
hmudg3+evotUsroMQcKW56jfQaEkubxa9cn7dIoUzTrvKshDZjkZkrFNDq/xs4BNFmmsCTUx05nY
2TuQJGpWSmf7S+/BGcEbITpnWBkuUKh+7elt+bP5ky99V1J3mIpv213gRqQhdjSdc+sBWQKC4CSS
tutqpQwuhsez3zxfZ8IWWFbsNq1QFwtAFNbo8HcZLVc1ZF/LxS/KT9MxbkeWfKbYG5i8SguD2OyD
qr5wf8ng43h8DJuqMXsGFw+7VziAz+8lxRDrsp4C3CqSCQu6A4oTgsqCayCOKTQjx53bLGFCErB6
n3QvuKWH5z3QDYXBk6VMlWtrS1CpVMTSCZkdvnEIDr+u9pnVcihkuMs7k+DhT2tymNExAuWo7OMv
ShZq0DCGAGtxTAEW5l5/CjIoFzenhXgAIusaZobytf/nOUb8hCzUC2FVNQIndTIst4+4lYnD3aBX
PQ0z/D2L/ETZ309R6fCTMOOw6aFAOh3usF7WwSLHTXt6cybhIdbOBUbNNS3+St+BWO0e82mh+XdR
2G97fxiXMctwn1KJ6wzcI93WEC5cIb9i9wBNigWWpeDIS3DlbZ0N0lJGA6j3q7t2j05V9Rh/oJFc
gTWDpKFCP/85ZmVS/8D4FC60PWmpJsNrZ75frYC3UtFVYOX9kboHx42fEjwz57RJ2LHk+yxxp9DJ
xyfoKFD+j8x2pUTHf96nWBOq8FnuY91B0IoCUsSN5em0uHUgMlZuhEZMOu7XhUS/wFOu0Q9IU622
oJruqyyvTSykf2n/cohi4zg2jHb3q9EpDCo2Dh0dh2Igk3y9jNOLcCFsgNcgl49Nc3OF40cuVDB2
L5L/5bA/HpKEHuHDef15Ogq2N+JG8B+YD35/49cbk8E9SIAOU/N/8TrdPZunu9msWgUJQzqfeAsd
uAl2pO1/0sz7Tt0bVoqrxNlMJixfFQ6P60v+oh8rAmC9ET6P/JOUzLAmL42aqFpMUq/UQqhWIP20
ZPXch6ehUAyqIceUTSnjyyWNWG0Fe1u0h6AOObykGACJiR0l+8VY4HG6ec/wN5e8XhcryREp0coq
pKk6u95Pa7bVnbeKnQcECb4D0ughVF44bp/EMc53M+sbCBFa2pVuhsSVatx9C2KD+i1J4ZiYAHR3
KP8SRJxR1Q3mFLei0VMZGHKfZtQ6qs8St2f7+EIo33c/bQtHB+xt0eECRrVyBNpySk1F3K0Y/h0x
doAfcw0jy0ThDz2qzZ9mywZ0P3OdQWIQM6QrHb1ALXGDuFwG74UL4nEvDEtT3y+wtAwv8hqaXg/A
HPkKRgqEMgqYZj03QTfvfpV133lwF3pjU1935JxfzHxxW5BMh8V0yD71yOoD5NEmhmhSMDakGFk8
a2TgDsBtIje4L9+V6eU1jb5Cn1Li3wHHpCwOpt/LgUeCqk62ZgD4q/vvwrkisD/aBi4zFS8B+GQU
INj8DtGFCsaviEmfPmVkknxV2ozWsGYk8XvkxcUz2AQcwcXFlhSMsJSk4n9UUY5bRkkQpAuywezt
JemsJvqD1na840AZnoPs3pkp7Cj7jvgLak2YinWB+B/i0WI4MXIZMAzZQZVyo44WANhIMowg/qHa
DOQjFvNXaKyZQWdBZQweslP9TAZbCpRFa+8HvHXWLxhhCsJivmijJvWVO4RC/Lh4HG3ENoml055F
MNnAx2V+vd7BatOHzMlPktK5Igjv1DMXMajmeTI0wM8JGIZZsZ35ekT5IDRk7aAq931xKi5QLpF0
xsJrl75uu+2Lbu9/h/Y71g8VZ37H6O4wrPuex8oYgZzCMhbalZarQVPkz0oH5ArehU34cW+VWeud
vl47kXwxu0Ga8vQZK6zPkwz0Mh7pB6cCxuFbtd77dWyXl7h+PgsRJNrIVGu/ESj4rHIpUBY3E0Xk
7pUES8R4DK5NZYe1OfLsfYUZ3VM0a/fUOA35EzTbD/K2N4l/nbVctXQ/ETtKRiyGXcTaS57410vt
K1rsBzRdbqWzC1tkfVKF/GASY7jvkaUKPSjNj9fPyC75OWzZxT7mlLPnLlKKH07vsYB48t5Tqwsd
Xqe9x0K6bkRc6U7Y6AXcy2VmW9AIThn+2wsYl49LFAo6mSZ+y/Toyedu54k1P3eRW1ReZ8Gfrb0o
Z35jbcKv1DRSfuBc0iTLtHwwKYHJG7C4m06myXGZAyJgGyIJzpyLDU7HRnAEn/yzZFhsnQ/9cqeX
DdSLIfKS55BCIHtdrGqLdaS6pE80AOsHlRvO+sgOmn62PhKiu4h7WiBovsK3fHnJYU0uXAbBZSvD
vrTrNXZZgookagoIxBoBhwSrFYzXwqa3yqGkEOlT3bqa4ZX58Wd+4jwr9DHanPt9OsNLXnwuGp0B
1YTeIwuN1Tvlq2tdVpommosHOpKTZZERcSBfhE92X3B2+SMs8CBjNKs44ua4e7Ojx1QRyqXgNMmF
8+KFnbm96Lqh51nkAuyVRFQ/3H+8joR6FPYJRpDqpbD+SEdBk9LZlju+wrlq6a6JLLEqWOdraWlR
6Ii7wM6yhAmFK1fbi2lfg1K27waZTFaesZ46plj0y6sFgAM59AeZhA/Z8KF4x9AKMly2GWC7V+Zg
exL7+mzU2fKEZp7xmeeYb4UdTJQ+QmC343P3pA/7tBlqbOa5Dv0/OwBb0KdKdyU9ij8xOhN4L+ht
ICsJmwnyG+ULhvkXwa9x9V6/R8f80zRLMk5hW4jYhcuI2qwD9fMNVvsUwm/NNulKpLUZW6KbCka/
KPynMizNPV4x8VwR42oiw8iz4k8mpuWUeuvs/IRTAirAwhRGDdd8AMsH7rUhP3Gaa2Xxy5ZqRrT1
ZwJMvtNXmGpdgVcf/lNwAEnbFnUJ3fy7nOGl3jan8QekUGhz/dRGVVHfeRtFkx5q/m9+bPNkXZhs
pXsCyrjrT1M8E8BoZ4UNiTc5PsArpANK3aslorWpHJcs302j50tAyyaYtZs55BgEkayZygkOqPsb
bfUkm976o4IPLSH/o2aStkN75Bldd2OayYOH3G9eylRktK8rwGgbmHMLS5/3hXe+lRkWn9hvuwd3
6BL4nSHChTbHfC4XACsN4+EdiSUTeAeMqYqkBZffKybNWZEXTMOdVqIcQTUQLG0r7sw7kB4olR6z
GE/QCG6gp0c4+mfKkOvx8hnBqZ5wM5AcP8+NHYaltvWJTqZQni4hEoUZP5PApoEJucytde+ICLMH
TIs/oDp1C9dE7Z2qpbkBrYNOrhc3NU6IUpwiRHQGliiKpscAMZQ5cBTWluOEqIhmQlfrCFz9Sw5K
C/EmyHol+o1kBaOeHaoCE/mmWejztT0Rs1fCNtNlepVlqAYvbrCTtimSsLBoulggOq+7vyXxYjsm
pARchVrSdbEBlJIIxskUWkpxEiQNJ40pl9uxmvBlj5j9L4qJ8Kak6J8leWnaGgHT2amKV2CcIf9S
glyhotiWrQksUlXA20NWqqwU1Ou+Jhg7KfPQuTIqEOhL5lSb4ZA7UrFOJonyzNnyyZeQPp9LRrBd
RxBZ4BrsoGhza5HsvHCa0PQKSsjqSEV3KQSCAilGO4zPPG1r5bGQkLkxDQrl18fTMpL4GNHP8gls
zqjdPVut2usobjIvkj2kYn3hqScRdGbEJ/YMCboxcsdjJEMKsLgYCgM6g/iGqMvSj9cR4DDAVuUO
FsBIJz8zY8wf68j0KVNSd0YtvcjCMGmYxkPMAX/wX+vJ7y7Xp1cKaO6Z3jn4oZ8Xq7ylZUqHXjdL
d7LrIezvJgT5PZDCy8dhOkKfyX/DOfVc2zPOs8sygjUjjG8PcSXUJRK+8ULM31ZFdmqCe8wmqOke
ZxWAAbm28n4mz4N/dRAi6+mzEpgrciI0LXWNcSihDsNzphhPI7xHQWscFUNX77ZWCCjYQW9E+NWl
81V9PYwDbWlJgrlApEi7OpL46Rk3cTXRT6ZNH79yVbCcT3Mi1VPI/WGFfx6pgOKwSMhk3qd/4xOq
EqjI+qKu04O1Zgdos91KH8vqRnnOBkVsPEn3Os2gufiv41hc5nI0C9WBPmEoSMclY5PuV9Y8Xijs
svAMPys4RXhlrdqg1z/zKAijvgNHuFkR5Nxu1KfaFcuaLq/IkepQ5m/OVokXZ019dVxYTV1roOJN
oYP+1fqyayNyD/rouTkY64gJkQtzF27C+fi8k4YDOJOsYPQSfofjd9E2JX2pjl7lwghue4V4ecox
2qA8Uo1OBhm7WeFDu3Aog4bsmXrW2JxDwJ0inekYSclYZcXMs0fOBigJsbUEhgf/X15P4S/MQEsx
8M6OAJgnaVe9ELL9lWE4/d4irtOxSnaWqt1RJwbQ7OzKW2FI4jaARfzX4MBrZlH0/yaZqVsZ4BWV
Ci1z/XZeyfu3bLLSKdM/KIfBwcFmiY2lWL/M+mjMcTVkZIGirFHlQtdwycQvLioW7ULDRf9Dur0H
HUZ8lhTOsiVu+BuiUjHafXLVOTQKGBWV9O73PrvnDfAH/+eC64bsTFiTZK6nZH+gDRkHu8R5CUmr
LbZ5RapTtW5X1ufdecVU+HNxYGL0oJXWGV+spBls8HSPxv/EBEfB9ZK5RC3WSOOC1Hq0ItimH4m5
LfbbOQB0+tQhsf4iiYW8XHVA1HdN6Uu1mNwtrV9ue5WoiAMwt3J5r1gmlB6TdQT5cZMkDQMecBpB
nezcSuaYePTgPhL3y9vb/rzVN/0eLZqp4U7JEhQV1sj0TdIRqTotzzoB028imazQlWf3uVr1yOLX
JDiZNwfQ6Gvp3yH0l+Wj3IGY9JIiJIp3i6p5KsLANbPshUzblG+z+WkKvtjaT4/9dNFlj1PPa+W1
cW09ZI+wmHxd1BqKWGfemktRKt6nacadnnl1PjPaaXqoGB4Xtr+s+wYn/szm6BWx+8oMpnhveJVW
+QDV19Tj9noCZ8jMW+t3KNoV5pjKvau7Ia59ZxZMhiZhzDJdTtIv/4vnGKb37iGpyWsIi+yzTviv
O7XccsjMYirtbSiJuxnA86H1y8/v0QMHBzSB0U26IvpFV1pHB8RuEwBIl2a+lP6nArl2XMqiNIGB
ZrbS1Y5QEWhkxj5W+3xhSbfPqlrH6cnbnpNJuP31Kg0/Qn8j86X45/pqVLf/vIi8n8/2dBXw7T9z
fGntcLJbRcX3eLgK6kX+U80s1z/gpRg4cnF2els8vh2hvelVTgMJnuHQ0kI4a6NDXol3NW55bmni
ul+YIfq8MzGQjm32/VGZOY3uObBs7WFPHNyEWSCsNVn6MIUl0pci9p6MU1XEY5ir1LC8rY26ulTP
r5cHy0EAMzS/qpSbE0TLlSWyrVJTNNDYa3RjIvEY6LrI3Mqr/jdz0e3ARv3tPOni6fp7CfF7H818
evewBojcX8RuYrlj5aZsLa+LHJttU/T4Zjwa4AjfFOpoQm0KckkydQ10KB4rHpZlpEDxmvsFOzmV
NSWA5LZCbYJnrdvNSb1WDdz8bSdk4hNW6Ry27XMsVYyqiRVlKEMyvSSuqQds5PHHsCjgE/q7mtsw
qkdS0iQoXGOvX7tt801ggUm5fUA9XHF9ZWkQc2q56wHVJbZo1bc0e9kFkT06rL4PTLeDUT+qXypn
OQzCzKuFdr6Pmzj9Pqml2dxYPlbtUZzYPDxZW+j8y+TKWrr2YagXXKtYXGkzHVLPRtnemUZhTs6+
w2jU8BKyLIsPwHjwWGy9PlYBBFcOKf/6CdnX252koFZT0rDRWU90OMzdjQLv+nS0hy7nDuUX76T0
+XyvHfLZYzb0M3pKpgaOIoDkr8pDda+qOQFoC5mVZMw4waN7XSIYE/XKN0T0G4wttS5aaGKsFtWK
7nVKtjThkRs6keujNWriYyqvajYtnecU1B14igNUGaSpW0AgmHUurROGvNfHgSt2y9Joi4v+a4SG
GKn+yO5+7wAWDeds/iN+o7U1v6CNplv9tA5Qig1sXPPqfsNWiJWEuyRVVM7Czq01+Z5OIdoFrgw9
DJPWgGB0m0fYK7pQGEycUrfaRmUDhrNpMszyFjzahk+WQMHMryfeSwBp5fd2gHhTBk0uey24+igo
Tl/DkURxfa6CCI3E2J66YctN2jKiJLeudfrAiQ0+HEBG/GgxY0dGFJRosgWfvKxqwFp9NGSkZOLW
f4Ds35pw3puX6PD9lG7S1NHlssgud3+7Upoua6AHozcJvIZOnX/ntAPUJe9Uz1yAcCzkyWOJVN2S
UOf9BAPCyPgCLG6koRY1uj6U1AKvs+z8seDBbVGg2vw3YgZcni2qtugMZxp1Oyjsw+jzBAqB1p4m
AR6Hs2KUNPDvrdsZBKDOVs1c/bwFlf2iomTd8XvqESiNzyKqApNkacVkA79zsHKOIOEQSfGsZfLq
RnrI8xOAO1ws9h6iura9cePeZvuLmD8WxhJO/hHJG04c2u0DRSzeDCZe/938+qEdO8I03KDVX24X
u1nbgmiBeFr1JXgdj5B1lgaozPRXj9jkCozDfsuoGUwKHQp9CPbUtKkIUupkGp/rHqArh8WhMF1o
ZX3vXBoOSB+3zQYi0smqDIXl2RaktmnLWzAmJ/fBe7NSbBhP2SpY14WDcYMV4EwZ6dgHGhP1i77y
gnMctj0CziyaRLoEaOhwxkytvZIMGj5rWvov+C6Bu9PwT4J9Hn1Fcm+vem4/x5PJYLfNhNwaPHmu
4r5AT3KCnFGH0Es53tuaW6+X9Lx+iVPkJg0kGwDvBg0kLwRkAbDjE2qJ7VKYMJFMSicSPdGQnTg/
cawxAYW3u+nnNrzf3cXUp1ieLS5p+ggrYBPJn1Ll+ld7+LOSkBWzJXHjG+fSAgP+X3MOi/ZVRmDx
Kie/9grMhphApIeK75J5hh+If4RjL+nE0LxPNYRp4AC1nyDdresew/AwYIcpPS8KcughkFEtvVAe
eEfglGLsHZMmJjrDrB/gLT3FRi0sdvO9vr5FR0f48ElNNXvphjgVWlTZ5B26ojlAnYR1Kxft3LhY
VtV89/rxo1QJnuU12011FKnTwfeXZZAvlQ8M7P0ZUdVpLGMz0o7f3zSDgw5TwDHTcFgByEZorm+8
D6uaq0vfrXTepV67CKrhYJmT0xcO9FJ4v4Y1KCZsPeKZm2HPqU/SGyJckC1ge8SoOsiKxdARbanr
1EDVpuftILYhaH4tefnMZLOq0WmUI06z8hHhh7ahvF2rSUi3zRHDGfnx/Y+TSDXokWPcCMLX6N2z
Jy4hFJMO5tC8HTEfyRTQNJ7lbAWCCwM9New3Svs/sRCmWF7SR/7qraav4ewTNBHKkuX+2SjJ2a8e
o1JyBcw9QA/fM6crM7KJCT/PaZwJqM9S3NA8J9+VYK5wQJ1ZvpA3A7AgI/h6ywGz82nkf2GFY2uG
d0Ph3oJ0sluQ+Su+Ssf3oIeir7YpGtnvhAKtLEpWE242hgVsNJV/y2gu/PwlUVRAmYggZjNtqFnS
OE4TlbGQ7n+p/W/2hS8fuIZxqGiwYsKwAD03OjxMEAVPBWu2a0PEAJbzBKEOsY5L0/nv2oQB/94I
IKVYaKq0m5NS4eKtFJERZU1R6A+yRfoGopJ3TaYsqz7iUtHm5hNQIP7uUFT+gqe0LlkWThXERiGe
5UUUZFQGGeE0mvqV+iJS+lBYzWA1j2CqK/rWfmqail2W7Uxa3m3E4TzSdoUbty4ZzpX5eVgz0WZS
fIgcO0qJKqiJbhvIfUuyzhhB0twROoCJXfWBDdjOYNIIfWEp7aaydLrzDb0AGi0lMz3tRkK3/QJb
BNWcd8pMqnmoCW6zaZ6KvlkVdZ2g+/QDbtt4i76HTnOPTo71wuDyivAO/+9Qu+u4jf4lagYRRZFh
HwfBfzcg2zirCF3tzyov+KBtobm6y50h5i9sfgovSzv2z88LHTjhpSWaFszQDOhWIc49FQDhYCNX
APfmSXFybfMkT4tAiLlc10ytHG3y3w+4f2YrEilDWeNa7jp6RD9BLeLqRrGel+m/+VIq86+cwi26
dP7mLzPgPw6X5sE0DOWMcLvocGGceh2/DpfgzYNWTuQiOulwnraru7QYmO5FV+7b0QNSYqGxMtbO
xAmdJyWp6PX01sQdkvv7wo67SWs5wvCrzSsx124gB5Hg5IDLTBwsnLC6xBgMAVMuxxBzbagXw4MY
EETouHYjQP994vAsmFt/vrIP61MJf8TtxdfSWbMltQsxflioswTc+cjy5qedB3ZViMgT/OSW2J9I
bJ/hgAbBmQVLyD1IMMX1l/ZX7W3mnB5Wwyf+75CUDaIF3/AvRxo6uSg8hGsUjQwxZTmyaF/GQhDt
8YGalg120+eRMun+z9x5pDZvNAeu3nj+hkj14x8j+q6jMrAkxskLNIlixJuUPmEFICXxrs/OJcqc
sqWkugYULsdVK0yCpCrYzK78OoQN5avYzASnq5thFzLQH/Chy/hHO1uWMMComBc/cTrSOcDM3WhI
XoCC+JyyZOzRRdinp2Sq5FLURjL0kk0b0raUIPV4kk6jfecNgWLBQsi4qWokARAEdCzmzM0CPV+k
qbOSy8udgNmPtZe2FFdqJ1rxAIvGWrH+TC3A/4nHMOe1Lxznw28Rgr5DocPJd/IkyNAgoj7yCDq0
DhQsQXGdP1pYvGNuGllSzuta+MY/OASVs4stbtBwq69U7Wn4B0P4pHJnd/6hfrNb8qXstuKRVq55
nqyknM6ky67d/t1nVCOUawCdPC/tYzHXKFxRBOWQgCboY7NoiXHxsHj0S1J5/teaaFXDeiomOH4L
Tc+Bj8oOByx4IECDp7Wu5jjXswd6pM3eRMe9GXkYe9itcEWdydm1Job3+AvqkqxRa01zWlu6ueB8
PGPhfY+ekbIcNijAEJlLlhHnIZoUX9oalbbvp5iwSP+Pr9GrAFNUYPR9h6jDeLUNva5rbUou19e3
OCE3EBwhBoOscUEqkSJFwP9QoqCl/ZZ7qTk396jyQ7k9OcZuV6N27A5yua9X1EcLd5EBhwtQK7+Y
Q+XyrwE5qL7iH1LSvvdf0xCSV4Y4Ha9/HnOYT72iI79m/uXutk7UL7cOohcC5bcLCDcCudvqGxeM
x23gU2rtDpkh870/zckw7axaN9vwDxUXuoos1zG+XFUudpVxp+zYOzr/bOtlaOWiW74DOR93Sq6o
yqKtN58onKts/gd2VXBlFqADYuHavidh+XbLgWNw8SJMNpTWR69FG0apiY9UJCDEEWT/4y6m76YI
utITGFIYCit7TjI+8e6aF8r1JmVcdbkOfjLe92ScRAozWovOVxce2cvhSnA2P1Yb2hguUkoZaFtB
fMutvbhSNhSWRFZRNTyzEsMLDD1+yY1VtA54HfQFPsjN+Kox84klPMxKtJegniWJBOYJPf4YHl5N
+a+UO5MRXNxclDkqoPCQy4g9wc9E9E2QrcXUMWLIE/LAkonMtG9c5zLYP6DB2FiZqLEroSrNC+jx
KFqiwhvoxomYMOraCqBQ9l2t2qBzpA3RIv20d6gut3mFROUABAKw9gOnjnpBNnT9gEZ48WI2oYwK
rE0qf3zpVKuaEk9azrCuS4MVZgZz/BKlxFA92QcZw2LNHDn2XC/hIDMvji0l8NmqFUKeSx3vRZJc
GefRTwtrdMH7QypKJfsfEz9UZmh6thRkRDcNyHcYRi6M2NRog3wY111j0EzJbeSdbRwHflQLwWzO
jKFwnTGO4/BYdEsY8103yOgvoVtmERVZB93FZwvWxh+k9n8UhZQEbZXatbExjjXtngzm4xi+Ehjb
qJjjylbFOiJnS/Atfe4mhcNJbFcsrOLehqyIMq7sk/rl3rdWY6WSCGV6OUVokQOJ4SSEdvI5QBCq
Htqq/TKKnSIU6k4kBZAOdwPwXj00QIZsdOv2GBh+++H16NNfweu7CxBT1gSVCRCtkbKDuhi4UMHa
nP+cLo41mrMZW+4sBQzcz/DeaEbQ+P6QI7PGoo3kmirpg2EILb6WAqyF4/f3n3YygBTdhjPTjTpW
pYwO9Fji1HYJ2K0TVbEYkpNANfXtz7ggCVYsrWNrWyKnEQuTjcliG3CTMY05LpScqeTqn6rue9oL
EmuPNg5/2yE+CFHgrFMPAozUjUKgp5J28W/qAhaphSSwfQkoH82H6N8OFcplrUZICmk7gg9yl3Ei
V/UpQNlJYFj+ywYDExKIpHdGIPhNgknsFtU6V15SitnHpGdjaa7ytL3kTFzP8qEmE83RZHpKdUWh
vJomK2PtU2sesv9hEUKTCohk2dEJu6DKSM3ojQMzp+w1yNuSyECuGCt7bePCjVnf9pl0Dcd1dVRG
jcYTxALLIKDo2MlitVGXEZAz1lYvA4mrNyo8sa2RLCf7qrnt6RxRueG+Ac6jBtTPF/qanRLAb74P
w2msguZ//rkq0aOtyzvr8Vcxu+5LHIOyh5i8AVKwB0hcF49k50pz1a85yn1JGWcdW+6M+oMfoPTf
fM7bDiCc3CoviQJt7vz0PmCSLOGTsgV9/TmJLzPHJRroayh0yNw4Mb7sX74KMmuJoqE9byijWItE
EkpOEWPWM6rFL77uwaToNT9DQMXU6ff8M2VXLwrDIULUeA7+s2EiomWMES/o3/Qw6zhdmUBSqomJ
TJqXuIjjT18uuf3SpHPhoUEbtFH8e5qOma6y1wnbWRk5ZKt3LkyrHr+c+5hvIGbAnv4vMkNfJu8e
l2YPgDC7X99Ab2QUdtMhO0P+NPrZ3stg2lIY4kMx1igVDNPK3DM2tEGVKMLFvGRP/Zht6AEKtvkt
jHZ230Zy1SCqKFmh+vHpkd6wSoOvJAVXDzfXgnfAvLZcvQSRr/5aCZvwYskwmrtBfqjAjap4iw6q
AEs74XoCYXYj8ajBZXzegz9XvD4+DflBO6xvn98uz3hwxBtbhs1FzNNJ1bXbTrP8p/aWJuqBf7DM
kNcn4PsYyJIQ43FCCnINkWSRIeG3OZXDyQpQqeDY+nG09zOwHpJamgEaqHVF6ynqhurV/p1qpLa4
PUXRHgRE5doJb33+afst3fOZpH+CcmvZFoZlG4ccDjDY3y2QoKIOlrIOhcm/QIKJore9ij05llDt
7tHr9Fwv1iYJyt+YfYD0p/51JDrNapA1t5IXkj0HiIo+fFUQHEEpDTVjYiE1wld6DKxR1CJq92F9
+YQRGIx5LJxKvHcmh+MEaDJBR4g4Q6my5y1o/SMGXj5LYBO0Ysiot72CZwu0Ik1i1z0lqkqNGHb9
Tx8PeTFqDRtH88AyeM1qfC65IpTQZUXUW+ig1GWXzFzxZ+4C4YuVNIqf7fnlXOAvrNKRpM17Vbvl
82Dhi3C9yVAVf3O9em7YC1zvs4Mp3sB6MgpMNJuqHHZMOuj7E7XqY+E4ydZTMbv7HpnXfNYnpihh
+XW7p1OOw1b0+Tbef1wdwjXk684lp3o0U6XmMmQVGs7xAE123uB+4qvZb0x/NetVL2XCZjtAqfho
/YtkPMP/DLnDJUCcUrwDtWCPClmk7wIQGKGO1CE5MPY3nMuRLcI8pejnx56Go9CFJsXy+ZOMTkVC
XPZE4YOEIGubZ77eAuxnmOEPaXm19W+sw8ldQHNi+nxmexnKjCHMPw7PjwBmnuo/4LK8I2GtGp0K
1MIvjCo5SJJ4Yy0Awec6XTA6TC393Ru8pF0j25j06fhNWK3vpJ1DnlXM1Z/r3H6Zbg0L7DeGEgeU
h/B7mZh3u6W2uaQ/wl99hUzShzk+jZ1PmxtM4AAVYqUnEaFfL4Yie/1LFc3Z90gyr98mowL0fqjT
bYLm51WQyPLZPUGSuOyyJccDman5BFD4JZeMF/XhYetUQMagHoAsFSEcUkEHiEtEET+HrVGz7nRQ
0Q6qZS/PH85GwLJerO1gGUEn3qE07VJcNcXfcz0dnBciQiXlflFC2F0Gjk2BtnDhhzntlP83vgsZ
yuN32f4RHIHmhWkJ41EsvTI6JEEYNkuRKWVbXBg6syAi+c5AoomeJKbsaYUybl6nZ9uvXMPhJegR
IgVeCNfhHJNnL6TBvtuG/1c+lirujhblTyogB9gHNrrII565iPTWtphu4UVC5+/35y74E/n9kluC
T82JUcztkH8xT7JZ4H61c1F3jj7z2jsNcAZ4+Xoq7vFqIV/vftJsgaJUbi974ESQjjyrR6qyqGe1
2Dax5XrNuvzSuRquUMNeCk3P4FXVCgXbDIMRQALkr77SbuNEoOu6n9+zf00sSWcM5tfhsFcOUjBY
AFOdDRysDtkjl1XfqmQVYV4jlY9OnAr7RPSFZkCv1xOCITmbpM5esXfWb4/7EsptPSjfXy235j5l
tF/yGg/AssF4fUZNbtpdIaAXWE5mzqrzpQZIxCBcyKWsAjFEburMov9nc51iCULtXwIAN/miMmCQ
7mUeFNS7ZtMN4Nho8psUuZhz46bI4R6fPfwUgGvzPHx3O+yeV9M6SklPv0318MEMm9kwaIvz7Dgg
WjiBi3B9VapGkARZ4h0NcQWbFyibrcnQ/GhyuyDkSscqqcyy6+v71t/bFquRUHNmJtSxB6s2OLDc
f0tsfbPeZVhpMiJqQcy+EgumK/EtnBHiiahtCfQ4vinnJJZ0ySWulPgqQxrZjv1FsadIakq4DLHU
NktP0XzjNWNIoVp+gGBLe+0OUXoJ/K5PVhgbhH8U0xswZqhOAX6fLVpRArEoNvbmzM0uNRksBE5x
CnuViDWBrt3i2w9FL2QVDV+gLokVGrr/MmkHloHw6OSIKyUz3e2YeQMz55UXtjjM/H7WfiuXaNYS
j8s+mlZpgpqnkoQJ7ptGpesw2ROjOYBjp/lzW7ql3OHDTqIr7NwAU67zhminyvYRi2obYWJ8Y460
Tgsnzt5gsTtfWtyTBf0yqqv8t+EAL/t1CngdD+PeCYstWMLR/N3xVlIB/3ZGlGiWzp3ltUHkXY9+
K1QNiYBZAwrM1g1XysfCMGlO4cXw4FW/58G30JO4bzQPHVzpSlsB5R+1G+Z8dvnOvWPfl6Tyvakm
7CvRj8xyX06l9neK3WonWUM3s0D57cunYwLNqcyIQxSjBfVSMpYf4+N72F6B8tPUdxLWXRldHFkV
QiaHAzMwDpKt7lbi7HGSWzuxx6HC3Ab0ksRkhVbTF6p5y50eVBxLUXNFfTvWkhGvUaZnjHNijK1C
4svNpn/4AQU9QyNc2ssoXlULrdvF+JryoZ+xUMQpzjG+98c5Oss+YUmv+dYM8Lfkm/FS4tZW2V5o
dQVF36hmh98mB6IxuZspTMGt/9GgaCqKMxLJZk+/yrA+QXOx/PjyCKUme3lX9RQ9AqD8VJLRlTUa
SMDAP5gXCTFR+6O9+8Zrj8cuXzibmlmQGBWzsoZWkUx5+5ld4F70DU7tTcH5lS9iVCMHiJ1CWx1i
zhAbVRyHX0jcrq4UDRjCh/goVpdrI+2gmzFQcmYglFwNKzzCIMu4K3qDAmh1tdRGYxX7aIWyPy1P
h7P7FpIx3nBhjf1UumcPAGkE92duXRHfl43xk171njHvgDdl0uMgH5HOUbFSFRvVyfwA5b6QwZsW
YqDlPjOgXE2wkRsXFsbPW/PvbfqC1f5aLoru3pMqfMea012Zik8ljInqI2NLK0OhtU+Y5e7AGVCy
dHrBcqx/IGIh9TVgriC/grdpym/nMs2oTfZUY5YvTen6n/MoV9AK8kGX50/IXZuAHekm+6Zytc60
c72I2lw8w2pmoynHLoe69FJ6K+m0anJ8DUXjvNgVxznIbDofNpsc1Y6hHF/NNGL0aBaRThl0Ko8a
L9FxMX+aZ0h1vmrS0qnj2dQke9hq/QetuVWAt1iK8VfGxQqWYRWOH5tQsNL/uCpGUtWSJYrcvGBr
2jT2fCFZLReodSCMREg0HEzGp7keYhPng+nc+kkCB9UBfcvdCq0NaD0ELoFEBUP71doB6z99ZNPU
OF9Ljr5AgpAUGLpJ13+rLHmC9Lzd0eOCq5Ab1rpV39XleEwcLQYi0Y6Zi7WA97zX1nkuIj5QMEkk
Lp/gUrzjaFLcN7GzrnG0oT+9UrCSzL+ZIeF7WXol/ATnoMFozsFVR5tbUZQp+Qjy5QPwxeF2cMTM
25JOzkfeXlDgPuHMm1aBZdZvlzQA9wINsyy4I4HfhucYWjGa47ETMMaJm3viQOroqMsursbT2LPJ
6VraBd3AV2pp6E52dO9guTL2EaoJdBdrBzkqOma4JAJl8azRj+t9KbFL6W7gHc1hHvllQcboVeuh
XSFvv1EmluDMSrDF7lAJW+lHdzWpOE5yttoPYQHMRPT6bUIDEs1CRLsDN/7zblwmMGJjVHG1hOn1
NGj/IgQEwRb0G5oxe37yaedRAoN9+H2TZI6CJmarVOu+k9zIUxi3TUZ3qQbsqpBTpTXQHfGrRgz6
WlW4m7sj/NL3FLwE4jQiuhAlwx/giKglPck5IM8VOvEDupzy1EUyrLMxBujkIEdyZY/iTmBH3K7o
11iEBEYmY+8u6sx2WIaH5h+J1PdnIlyDgMINTjnXNZQlIwseMMN/mMnqHLJtivnowU+o7N04U8Qg
4V3HSKK8qJD9wImnUISyo5Q1YQMVVVudPKeT8ZIKaY6TL+0pGy9BxvDWGLeow9Z03lTpKLbziOPG
kcL1aWwrbfsUt1hiFwnxC/ApgPwAmyU4TTmUrLIbsBfXmqmJ/rMkh067+EOR+f8/VBaX7Yg85XRZ
C5yxUIk6QUHfvKAZswRozv2QhWj2G5Y3Zg3FFZweY1cv/xH6uIi7vI+euyEJPNkQm2f+t+v2xRCC
mfAgxe1yQ+HL8UwEAh58Mrb77u2/ute3q7nzK+uSyCD+UJqo7m5iDc5MUvSnWZ2Z0nk7Gcj418W9
3KxiUOONlOqnFTobKt3PtAmQ+w2J1U9b3SnvRkUP2hsQ12iGly9cphB0ePDVTP3ZlEfjdXEH7H7n
7Ixvc1k9TonV6KY4FGq4YhDum1AYOy/iyjGvxsQvFv/quBtHouU+nGhU+nvzr8zwda1q0oSm/RAS
L4qz6BlS2a99ZztCA4pIrbt7TI6WTKK66Zwtar4IaG5ofNm5mg8rFKan7ASdCgnVjZKHY23d8/Hh
2/ktVqoTJzfRJy9fpQDpLiC833LhVrsQPSjb0BLSuPKgmmuREOQdfu5J2Z466t3a7Z/Ogm1p93Jv
NCuA1cM07uAdIVo+LIKWxPyr9BUimQxok4hj5LiZ/VAkEF7ncBBatzYVjHs00PLBEGC1HvqRq655
5SQnzZ5scHznmLruhGGrYyefkXB3uzlz/IGzVwSzrw0mT1Fh7RxyOjs/gQ9uXbjJARLTyYXNcEpO
8+NEwdxcte4KpZIAO9r293Rs/Ym5cL2EJQYoOgNrP/OdbBQYEJKdaMJhQfCzsoxiYLKXpSncbt4F
wVzeN/TZc/qfemy4wHxFPrU8T3zC+vHRiSA5sBUyyyTZ6bzamnWUW8MUmLg9sEqxMLVYfmqn1k2L
cSyvTe+rdKTV7xNe9v1iECfBjGX6rL7ZrYwLSOrXxbfDqcmFNtUrVZZxSYA1FN8LggPXDIyBwtHw
+fEWE1SiTj8ApDnqlSpv5En3ixZXgYoUHgWQuX/72sQwpYAe4/QoCahR6/hObERebNYy6ih24n4Z
AQOKfo7mM8qEbtHenPn2iwhWHGPGEhqQD5VX6ulfvg8z3PXwe+2w93U/CVB3aXZjEVpPQk5/x42J
GlLMqByJ1vZ6TGYGTTAeb03cdlJhRjqFI90hriiDAcpTVB/VZ/XhxKt2ymEz6LisKT6c86pxglne
boSbLJHfKDwwYEHHJp8/c9FG8AGDDT2rXiP3FC9BkT8gWlo8GndWMwFQpqDe4qfPdmzRJw3KiWVM
cik3GmAyJzxo8QhJrlhHsnUH9FPjDzIUhinolalYQcON+hj+pVUEgA8MEINPK195Fwt93yCGXW/q
3BwXfyWeoGV0iWpuyVkNGLAIP5iNWlpCqEDQF2pqzCxYnbvpCqs1Oy5i81Z8rFV8bN6M7wZYIaJj
APgouowToXb/h6AdP0hqwtdUKLziupHESBcCJrp9dnP1222KWpDhoGi2EX94RDn0tqeWNnGmEO2/
xm4vIGabOSn7Flq/rr/f+HWkx+DEdiz1UNL3OmfU55KQmsC9sMVCTc6wfga5febD38o/g/aBot2f
IFMqlGub7zAtc6a7dPTCJVdbwXYh3pRtTXnfYvELaAydDyF99drbgy+74u8FauBI97iTVSfRPo9P
Egw/BV3e9Txpc04A9yfSuhdO4qTcvCglEjKqlTNA+71FcElARvxFP56ahFD2NuLBKGtIM18nAnfS
RYKmNNJSjOSuEgyr8Z2WKXHXlnsjajQSt9f2hniW8v0/0OeT092TcORe31c25U0Dhc1hGkj6Y+IJ
Yp9rx76EBXeh4u5GLzxsO/Qpp/HOW13wY965Z0wmQdTlmLVwpPh87S2yJO99hEYOIkF2mt8mlmut
tXLF0VaE5BLhsHDrUuxFJdAXJLtzvQdcjCxVUhjmD8pNwaWGp2Yy1h8Jx/dJtjbR1Ii7K4Y7DqNy
JxKq/xUSRMyEyI0jn/krK/wvvgKEenfiXCabW2og6O+Tg/p/iqOmOua0Ccwk51CDI5Y0tw667Clv
ZkH5T//P34+lmPKgBMbkJC9HBhCLzSvlG4bWAR1tlbPX+2pHHWos3M6tI4kTDlJ8jK7kbK0SPbDz
KP4EDMj3L9Fs0OVPZf/DAWoxQZztjmIDUYfbtPbwOVSoNuffSqxhQPMvSDcFzHa/b3kgMFHaGjNg
LzTOZOhBda3mzGyaSR8+6w43QYERj7WNCx71/xI0GsHQ5+nanBxnu5ZNk0bDPWqO+7urbFyxBvHM
cDPL5vq83/dewST2O1plNzTvqXwGybflnHDgPzUe/nukkrKfo2zsT3nMSmgzzrGmACGpoSMxGhcC
2V1R9agcUYZAyC/CuUIqVtGCz11+1HeZrMt5BXIT5BpJS0vbLyH/KwoXBhBNCTZ9DhBVM67/BvKy
g7uvefuhfgRuXr8jBHLOKfP2N7VIu0Qwf3MtjQ4Gr1DbP01VLb2ApMCJJgH/bdne7w3FeYHTeyDY
HdHDdfIePI1t5ZT9yGuPpJcSNmCrU8zsIsBNPxPtLvVtP05615zZbpd5Yf54WUONurWix7WBybry
NIh0nlT/jupJ25Uo5/dx9BGxIaZ+OKH2NQ6/COjdQ7FNlnUTwN3O9Bih1dAT5GOrJy4MyyG0InEP
Cuuz4yZZ6xkHQv4HDE0+LiE/6iTpCPe9b+kLyN7Bgv3mWRhjQ9+95arDrxKv+mhc1wGbiBjdhpqd
r6QHIy7pkC1kO9uEIpb9LVXbNmRTAExa4/R1ICwonV9HNEcoy1/bgmQ2l5dQLwhrosfw4MW1O4XQ
KBotVjlcP1HM2I0UjRPBPSPdR8Mp4P/tcKXoESVNgP+JZhCq4UORUgXtSmSg49bZ82S272+0eppc
aEka9M93jMsx9V02SELk46QPLWytZdedr0j6nKYBxLcO0LxKT7S139//rvRJ+e/NTnE3ZncI/nKz
V9Yoeg8777Eh/iwVOCOwOezsay5wlrtgU2Zy404//530Dy3nzbsS79XJSu22hPgl3qV43a5uDXzj
b3jnZ+Ft6its1gchKa0tO1NvlKj1BgRJ0cdPfWiga5VQ8/Q+R5d9aXF/KnEgzUS+w+oWLkqyWJ7D
KZJVYBPQDXSIGrLiNI8ecMbTtYHFODvFX6lYdItweJ3PucWnDGB53rt3CKXyPY9G8fd4uLufumIj
P8TVZ3+RXMrT6m4DbUf28iJt11AYBDtxR4MNxIeNfTUmUDFfrfqecM+IQBNqBMNEzTZJWcoMfA2f
tZ42WOzacWIjmtLjy4bPmeMXTbnq1JMnoTbIh1+4LqVySnil7an0481MOsVWHGJDerKewwTogzRi
6FjkInTBAiwIHkGpF/tauRb83ZlpsiehMbkVk+vWk9cbmwI59j/NfPRtIhxHzvM9oaQ6cZODAkO0
/kx6XsRyZoCcu49RylbvlbgXW6VT3VzXur/Mmn4mY2rm4tbu37Pvo5rOE5DvMoj1EACV0F+ydwam
Wv+qUpE8pekdT64L7JNHpQlgZr9qoBeHKXFiU33Xm36Lq5nKmBQuPH6+vxhvwR/NPYZ2rLGzceee
Z19C8tobVCgOur+qyebEDi0C8hGxQ43ajx/kaC/WrsqSrafy4uMpk69QoQjnf1A3KPP8G26DAB1S
4lyBKAdFhFyGqXNtM1MEnkqv3E61klJ8MQmrxaXHX1DWIACHuTd9BdU3xFmIsuQNhHgYuQ9JGf9U
vnVGvpMbDz9cE/xFCz6Slk23AApOh4C4dBYEgcgSt7zgnch+nWJjb13IpIw4yaREhT9r95odKpNe
hnEnwByaeyRBBajancy9bzv6lHy8chlSIxgJtUCnvftAn3oGUPRjHmeIQazHs29xUPBURv1sVZ8I
03cNymXCCbbuDppAiocT6yCqY65LGrghbYEq9wo37BFC+4SGJfE2IbvUSu5sKc5Kyfbs5RyM1Vrf
8G6PPmkRUnV/eCwR3/Gxriq5DYzDUCjzhysZ4+DsAHK+Sa+krQj6HOtWfqcnTX6rI7vmTgXD9lyN
qSiZiVDDRbLOYJBdww48oE2jI+r5d9grsBVsCCpk/gnGz90BUQpwSuOqL4IGRPiKXBDsYkjbd4mw
fNFl8LyvjCcJ9NjjMF6NejkYIhQUQ/t/ZoknA7mRx6uftBbP3+rNVPXFE7KYz4bFUdd5yvkO0KiE
iMkRfbtz4pyHSmbbXwWgsArDDcNpHA5g1Fw5x4k1CJlX/rwcy+1xuykicGsoFR+r+CqGvdN9yXdq
Im2Ns7sBeColXwHc5k2G7bpDavIE0RKQy6L/pv6Va4QD7gf4WJ4QzYqIVbdT6O4o007UF8KcP5q5
PYIdoNretlCWUhOExWZWT6EUdAhZ9SSoSa5AUgtKdo6g99Inmv5cmGxAgUt8o1kCfeZd7sc/YbYq
X78wppZmH/bCD5iiyy8mwUk7Malxw97nuaWNbuXIO6cxn/VgO0oDd6OKl0p277WdWJuOQ/pozBeO
pqIeshjd3/LEgnDRkw89MzXXPBkFDYlqJr53sOfIviVgUPvDQD16NavR5luxH9NCkGuGrKjeRbrM
WqLOwtwZFKzM9dJGgBoMoiGgatB9KQvWEJXE2yR6Aq2qultxfvqIiYeQA+NFk1xzj4S7aeHThpVQ
luf1H1J+WLZGJBK/vWu/2KvCVKijTMXcWLVXGZqPo122j1LyB1UTBwVuJbRmYD++KgcKQ+OscElO
xlaU1qDZuSVhPg8pxJmAHzLlKtPzTGtRW3seJ/8kioSP5P66z/JXPeY63qccZQDxAMNz/aIoPquR
O/eT/RAjZrb2/tLa18AOOw31Bc2D2hH5GMuWd4tZaGPGfshAJ1HhRRkzpruNU9eR3vBtpJgDeNp6
5ovgFUy9Y9CXO3Gqx3sI8GJk1arnCnlPL4aYXRa4scMXpcCdYFCqZVi9zhG3676rdqfC8MhMixbm
kFjoEPdozaB1ffa2Vo9afDy+qagWvXwdl22eTyt0JkfmJjcqU93ZR02aAeu39QMXDLLlxn/wdWxK
EIXhH4L346fpLracCYau6zTolaxrspFbtGENSy4muCUUG6DrEoYAehMIfGK5lTMkU3FvM6J3zbSh
SXCjpayXvDgp+S9MaLPLjdREi7jKvNNPUSYTZQvy477pSfjaCCGPYhAfcerDP/GpKMYcYkYLn30X
NLbo3H4+DUhgXI0ckM1cjUG8gTXINRinF0HjXC0AkdNWQ/blAJ8j5av6P/HuaSOCMc3At4ZPfvBE
eZNfJ5PLwU/qSdVmKLm9EFK19oZOLmKoj2xryvXS0PkU6mIf/ftTizW1UJoaUiW3p8A3qdxBG8If
pdh8MDGcMhaI30cE5qMQrZpguqkBDsRr0U/YABltrsKKt7o6se3fKKdgW3HanyRvs+wZpgWmiOis
OLkK9DtlZRhyQDaXYP+CEOI6pR7JGfwG51gxZgK3edJBMyDSdaieXuE6de0niKcVgkTvlspll78A
qWc72oIZ2rCQNB8yqwtMvyEotXrbHbEu/gO1iVyU1Pt/sKcx+brJo+XDYyEiPeyBbAYI1saTunzI
RXp2mTL3hTg2VisecSpi8ieDG5z1LYww1gilN44ode3xqNSIKrrABezQVvnoIKaOPbeL9eV4spsJ
i95W/gelUgq4GUGV1Lm1Jl3xljxcJiG9aiwIxvGyTR2IMS+XpUaB0j71/+LVDjYKKi+nMF5Gsq9a
d1cJbhyW11aNPKX5uJWtuFdKMbEERl4+0PPhlAeJvIvQsas6VO6ozFp67jXyHzvTY7r7IYC2mtfW
Pd/QaRIRZLdL8G5txcJfb9xuhJZwoefqKSitsyueAH1gefwMdzsBRXUFbQbuaSac7WWkk93WWgp0
9eegZrEEyYhBrODgbZx8dZa5dgBbycwxYOrLI23JuesAQ7m2o+mt7tGhVrRZk3xL24byCqWkMflA
FOIIWziDppUBDRa9pvXccDm5UsdwuJGb3s5sfZCwwz1QtVDOcfTJM2ZyG5wNHUnfzS4Z/aWKjcza
8FnORHnU+djn8UBLR9brMinYjTIE2YPF4SNAHe0mdLWuc4sPZbxEvd48cSRfRGfsH7edMq6y7HSb
KGNtjzFqIRTmyWky1IRRv6SVfUpjvbatp+MIPwzKhWqhUfE4zEPBV34J7Ajo2qBrRjdgcwN5vxlm
w6W5bkYBp+1uUZDc8UUpUWsZP194CNrobZB1LKdIR8yWHYf2aMq02en3v7LsT6EzeQxbygtqdsKp
t3W5yZDj8rlQ9ivoN7g+hopk00Z/hbajRW9Zpo84IOte5RHq2a65OnAoP4ULfbYQPCqs2ZgBKtJK
18ksmMlKQ/LRZtoBY/w5OtdjV2BiBTpgEqHFbDBuaV36gvd9ZdKJO/24BRidFxVwY5ELaQQ9sH+g
n+v5bWtw2lH7qc6GNKmUqPSldWBi3eVbb9THyRjXaQ5ie/mX+evxjfNq3ZEg08HBmzUeXfAOVp5q
SOSiC/Z7t/uUgkLP6NPvBumo8R6Xph+/QcJO+PeQ6/xfvs2fAlrVun3eedo1U1XXX93zhVyQNVQF
P6lMyWx0BQlLODD/xe9x6YDvw1F6bbVGTsb+2Q5Kj3B394U05KvwgmdPf/Iqj4QiDOYk0LZZEBRA
qa5OPqQuJblSFco0R1kgMUUtw4Dx0GtQhyugSiQg3JaWFj93tAgEgtkei8iYVQFrS0NKoc8v9bNd
W24H+4AUxHNFixDkVJvNDSGi6HfxVWkrTQgVdROEbxedASdwHmIzleASP38S0Z9hPBXshTI8IHlw
gPj8QPQq6mDC3PVYSlrc8TaRdoy2sZEt06WkXTCNlYFM56Z0svS0/QqawcU+17LpMZzwQqwjRv5T
OggXTeRfmzLiFxl57RSvnTTFLdsVEIoYI7InMruP3zpS8ZWIzYQSppyou56QVBZAuA5JAL2roBRY
hzuJc4XCgmSpM35Gf9YujyGWQPbl0e91Kh0jXdzMdOUuv6g7fOcCnB0Y1Z5GEVD6MGJBlVOylccV
Z2D/hXT79j55Dvb6piKawsZRRrsou6P/SLLSgLvpPYdtclFSgsmEDdaxxBbnd8TXUFgxtUxifVqn
U0mzuTj4pR49dqRNpltZNuPQI0EgYzQPletD6SPsIQX/wd6I0HFJcma4Yudz8F2z4q+Vzhizp/CC
/J1SsSAxtRbkZx+3ciePRi4bbE9VWZ3zyCtvBjwa8RFj1K65DvABxsUo+aLtZrzmqJj7ex3ykMn0
xxzlvM89US+R9hOMviNc17/MoAIjvQ/cOV+P0ZzgeVJQ8YgwWHWX43p7ExEmbE9wFpjX+NGa24ya
amvjDgbM0xstYlAoX77VGJoZ/SI9dHNhcZZkqvwmRfUF9jhEQUNOCkJwWn0oUnQN+CzFnXWA4l0Y
YGG/ySlRUQOIK8b01MIuWlSZh++W6oJlNpuANYYDLKjDqNkVLoYffHhgFad6sFk4dgdCsTA2cUCC
YkWqaT4C+Z70/CbMpjyM4YtUKhbfPHad2BgImYjPhHABWPF0fq5lRPGFhDzEEbjPQ69Ir520qHNz
1eNZ2udxMHf/91DIyuMm4WnW9tAJhlRNXo4vNATykLgCG47qROGkUy/aZUXx6D5RyoOlN6sqoK8x
IkZQMg5hENrlOFbnB09zvBDfTlVt27qQUrDrEe8n6rxLiW6kPKmoC0wle5gtTqm892k+BvfAfkEE
KE+rxwLBpNhK3K/xBcLfLiL7QcTmpWttUWIfeKhHTpVzj1tVOQM2MCKDqav9S9JMx4ZUAQ4SuQ/9
Kz+QiSIEN7yw4W2U4fEUa0P2GQGwY48bjiD6daqnQMjPcwTDJu5XlypeBcNAyshs4zttUC3LrIvM
B5F7nTLF1jKQ64v3IwyLRo47MgnRnlUXopF+ygaXXp7T8YEdr0d8yNnYHNrR8A3cvCTEPrvnYXKn
NxLviBotJAx2FMs4NLpaPsXoeVzg7pJ4XoTsjE2moJ56B4WoNi43rT44xNE0V5oLkX7Pdms3ep5i
hPq3dcHiyYZ7izIoQC5pq4Xdina4RzLWpsFJZ6aOzJoxaZd6kJDewc346vFuifRXF02vYmuPXSDw
rGYyk43hgr8p4x03QIvCflMaeM1JjjWiawToB/oN75CTwJ3m64N5J/papBdmOT5e4/VSuwgX4rOG
YtbOlwtUGYecqMafUbsmhFsgzGGde4fe4dfnLI3trKGJQmMoREDUxz4NB1Y6FB6g4wSrOPJkEy8K
KsOlxWM4tqjtEyE1gxlDyHfS+2jaAhkN8rA6i8GWrspjr2B3QJaht2k45Ou0qb53v0GxmkqNs2n5
uOTsBgzxVuwq3+G6UycEukudKQra72uSZMb//B9XOBikVY1J+MO5MdsCR6osBZzyVCq/uLZWYdcm
wW9S8c4YuRReUER+Jnv9aeBAJQdfK3RzGwUoROh9+wmQLVYO5e+YCepFCw/HJSDJLPP4VlvSNCUw
CuswU8De5m6iqZAaExP501D6Ug7VULa39emGZcd8tJdqr4y5oE0lW250UVPrd5QzkojoPXbhV0xb
McxhRj/xao7EZVI4ZrFFrojVpEjd8TwP/PFyGl5jgMD24D/lkHNoA9T2ooO52CTwAvX/EKa0WSmn
dkcm0ZH23q3b4S6Q9gwq2bhDUxTLm7gcDLskKf+4JP3XPjFGVsllgvRbzEGIrxf+kE5ggHDzlpfL
dexHOckf8Y+qp3McUWlR4ZEc5B3MsR2NCdWOQKF8O4ZlLTkek2Kxes1K1qpVEfL8QHPHvR+uE/+V
Q92CU+gwkurUz9AqSxOh3l4viPe0kXsc9guR9FZXNJHD/ZBwOrDFxq7S17tYwQYXzW4YFBs1fDst
2NnYkR1B01VBtDx7olsef0EINi3EtZgh0xsCRURpu9tbbyjTTiJzOJuZytds/CUyAQwygDxigYM5
DjZ/M2luOyY8qwmL5h0Xk6A3aHGzZNsvrfPilD/v/0IhVF3b+GG7BxtoKGtxrZh2HqwqXGAQEtgz
CbFqHixr/nUQImzHe7oG05gTh/STuFgvNjerrJn4JtHBC0lYlxMLONk0ZFlAnfBiSJz2pUqcuZo9
C+FL04QKZQLPRNwRWNoe3vNYdBSlvvWmkDjvwhLJVR8NZ3E/N9InzpCbHYP2sXNeFKEUuwzLd1Wk
kxF3CH4B9SvS9mPV7ZmxCapmJ9a+N1ZUkGCIA4B8X2ZIKpQ0ZClg0Dd4xQLc9Sw7UiSpFxuRpcJa
Nyqn0+6En+GaAx68ouuXItl5UovgYgJJ8jXX0dxgqtiuvabg4ayTRNh3GsrMKsNadvs8rqTtD422
Iv4ZgY4pCnXzYZyqnohscXEr1OU2Q2HBcVsLITkHuM1fvnc0fAFmIJW0necSKYBUczoEWihIR+Gx
YXf89G7A5ClNdBNtk2HjWcm5/ba5H72KYq766yRDh2KyFgJaeUpwNr2YphoU7DDJoyRFHNlHW63X
4sXn/zNn33QF2vcprPg7x4Hr/rS7hoWSLJfz1luD0RamRENYYtsXyS2NWgyedoV777drLLsfQIpO
fITEWDw4FRJhIyPbc0xqeCcFL5C0iwiPUPDJLrYFB+nnWCPc6UDswTBuFg/xRpy+BP8G+PHZpDFA
Wwe9wwPKnX2chCBGYniQIH/hsHBfNwyjcYpdF/qmbXYs2LCgX0Nvhvl/EWp9qhm7SWN/Zks5HVxb
NXg6H2tIY3Z3jje4nbIMyVZ8Ta2HLarZzyE0jRYmMk3uJV8VpAYCH4pV7E9wv+ZFxksnAcljH3Ga
Ob3l7yOh0wInPS2pfvLrWUoaXkH5x3tc/laZ+5dNVsVfhkHpdEa4OUaqura/PFH7lEChGEwfZISU
0frnNlFI58ULCSGbzj+yrb3Ope1W5gMmGYldh9MwG4/JMMFQ9RtPs9CiBtsMSi0OrIxl0aIKQv+I
TV7oxUjIjaXG2TiQSRXdsdw74whNU5468VCcY0gZ+ncO7UMsITs7edBT7YSz9eG5Jgu/R90lhJ9J
d9cuz2FCoM6u/85cVGTEArr7qFxXkbUVNDpQN2s5SKPV30J35VQcursDl5SB/en6lxiwALPxFBrD
bxIWrCVaWPXhbrpboV+HHjdvSmqJZ419OtU42Kc18AaNx2gbspNvIPGiCcNHLzqB17yF3QASHziO
cAOKxLnViXZGAHrAD5KpLMloWvbhbtCTke1aPdXrDdPHA3aa98jMhJHUC6tuk8SBRZ7EfMKuTytt
16KR/PYRAzframcfMTkT/AluKuyVqG68JhpfJm9duZypRfpRw7xHUrt0baHQljw6qBtdr4UQQb/3
9e5D6ZDHbm800I7LKqGPWnxJ0XH8+iRUdmHA8pVmVIaL1LgSawCKm7LcX3De88Xvhw5Tf/pQ3Ceq
XefljDt81zTxQ/JtjR8c5Nbt7lEGOeiZpOxE+OpGnerN4tzrpgbPx81p4Hxamx2CkD0cemqLqY50
2pCse6SUbZT9LYJO47d4idnsAFQ69n3ReOsMCXa68V+fXwTgbwWCztpJIpob4kUBuKbg/hISZO6u
lXo6a6YDxzZlVXfuYYthQkZoUM9rQy1aJDLnlva66WErxt4BHac5H0oHc/P12q5gs+0Qb0BUnaHL
qFS868ptoTE6JAxHzJZK8RUb2zVeQnCFx8tjSzxj7HcphorKRqhLOV5h8GJ02WTVhF7vtgrJCkaV
gpY9Q6UzKWslPiHo6M9dSxftQZhK1cNzV9IHFuocRirktHlUFmN9V0x2dPaGjNqaGRV0zxtoS5IX
oui11OaH221/kHFy8NM331BMjdJ3AyJllJO0lgBOx3TCmOmjLq06cOKva2Qak0t4zWntkSdAPSqP
ZVT5Fxuj7dbwPiHWS2IquNIqh9TPZ6chgA9wI/9NWzCPe/uHePZlIQNq2JTonq7ouEbyc1rvYgz+
woXH7QDwCL9PeMf6eh6Nz1TZU88J/9wQ4WvPs6NZLU3HX4emMqgXJP48KDFS+Z5bhGNy6oh9NQ8i
CoT6BbpgLuJXOko/IOHkdbZbIDst4rt8HRsT6w3o4gvkjVqXbHkwaDtVxmAV9sn+gmcIV5RbkuHS
pq8IMigOGdp3T6DJ46Qt1WheJY21waYNAJi/fiheZwajp4opDNiABPEKDepHV48fGQ+FibahHIDd
QQp3GSiIsFu/QRHEl1+KmKwxetlyNlRJROdt3AmPCOHT0TjI7Zrjc0nD0qy57eJNx2FyoUr2VpO2
f+1/6DI2bCihvsv52VRPg886ssMi1+98GA3OLtufdFosMsX5Cn7YiEJI1c9IVay4NKQ8FVmNl96q
WQHp9VPT1t/VUrQDHZXtsrCqEimL4AkIwIWzI697WAL23q4xoGwa+fu3yC4LTac4xgAhTYHEi4u3
d6VIC4QVyUQMd/GDoNYCVrl0ew0NMmXxmG9/WtXXOKxAEe/QLYamakaf2t00eMQSmSNuhJB13kcK
jC/TTtsaYwkvYIhK60alPBSu/J/OEHjLfpYwMOCKaycwDuIJuBbsjFsMVObQAEPfJAPwt8E0xLjd
ON/awNAagbJcOY6NdfIbrNvq/DzyPTlmwR/Eu2yNRipFIrcnFn61jPYzFbm+CAbAbCmm4byeTPvM
sNPDTevBPCU0ShjXHy5U6uCMyYwtddNCvAoiNWgiKeADeMLMkwelOLSlJoaA6q4T6ZMrJzks/cAN
nmj70ndxq17XmvxOKfoG4Y47Zockx/rG8jN4Y3PdeFd2BVGSUIag68a2jGuUrFysqLEH3xE0WPpb
wfpoKkB4RPyopLvTfssJurMr9xlIM4M2PPZIJss9ODesJ8v7I/FCCY2toxqFaUn6c+3xcFyxUiCK
+waXcvm0Ics9Mrp1jgnJ/kAWXsTYzejqoT80aCklyLYA7VQbPSmwUuw8V7DiSId9byDqYnLdWuhw
iKvebR4i1DJ04lZEq8jDPA7Zve6YqgKpD95uz19RFR1hj0eo1gLZ800AiqKiFOAl2xDRcOVcT7B4
/C4cyhQEXxzC41v+WiMLrnKnduyVY/YtbWfXa3FA/1xOwS9g7ExNs+EMH44dwY19iMqjx4xmqBTm
geQ/vOfzTYJGowRn8Y+hFGqBwp7n7vjfuOa6510OwRrowKOBImnrwZti+H1BrVDnaeL5I8fX4o/Z
AgOn2eCwjvgUKze37/Ekpxf5YF0yOd0IVOSGkSotMqDJDY3Nf/BnC6tsHGycWpMFU1w4Ao7pUOe0
PAA+LMhbxqnrL63y2ACUqyaNkzbWK6tXgnzIZqejBeomtlbwHloz4w0gJW1gsEG2mGEndOeehKe0
y4s/Ub59zbtuSmsoosGXxXk5GDoR6GtFbuQ05o6cMQfwTRykXOKGsKJ1O6phWtByVHDxDaI/Hqdb
07wLHDakLlG5zB7jQrKS3LBdZlC5DsKr88wpEA2s3Fp7B6pi13l3gC+4Y4NCs2UZhaBcETxonmy4
SR82od+bYl1XM6XQ0a+TpTiTdqX+BrfjjP2wC3nNX9HTvtgfvbstMd7ysH7yH7heljkAdnwbJm54
8JIeRZuLs7QdtvhrfSHMhLTnAcvZ5wMsJ3DIIQNmllck0BGevRVEw1hG317q84Qha+fWKFm+5j0U
6DgbBbt8Ta2Wtqwj89wNJJU7mqn/PEFIN+zfWJ+4I7XxiFneEwTkao5VTpYeHRSLrUR8MkvWaIcA
dpUgyozmyRBktmfWhQmHv8DPGm297d8GaNUwGa/5qCpd7vGhlICVvDIKT7QGbDLivX5PvSngTmWQ
GlMCzOcTBqZQyY+mY5cNvfgOddfQ5S5crYrGURLHrPjb2SlGMuLRgjyhegjlHK3G0WswJ3IxnuIn
0rWpmCvR1t0mxtVg7h8ekk2KlbeEDIkLlsnEmfD08npMlWEDnCCzXTCNlKPnE2/2vmyyO56BUNOQ
Wg+6tag87Ii71lgQMLmkPmLFgoyVP0pkiwW3uBIiMTcLlpm/wlTnc14oF8IqAMKr4thbkj1wVfzI
SdjOaZG4bJ3lfKPPVID+UvSrsoIpvyaIuM4ABbQvTLEl8QWNgrn7rHbiPR4u7Tfdm6HRFQVM4ikP
6f9x71brv0BJkvhpTQBmpWvz0jwuZIwDj0Aa3D9ygdnF0X43TBBEkLN5obXbjRchq6R0lcGuLy2E
PLkEa8i1YYWpYw++JoCCf7Vzmtlgq/AP464AyNjp+KUW6uhasrq039lqpncVO8fFF79HeG+uNdUw
8EeP7gdihK+dUX1wjtDnBiTbd+9124I78Pbq++bJ0JKPdPSwoMmPMQRyxEwzTJrt9nC1q0Uggt7q
+a/NThU6nbpkKqcyfCgjypNsXwk/a86LABnpzmoUr9QOReMXg2JjCCU3+VwzSWO7rXHjBjrIFPPb
/DWn1XSwdoHwnfvJqLThtYzqt1rQ4M642cDNYAqfvYV+I4W7BeddQf4Vf07koB3ooYDMMWQBFG0I
wEc5PsJshjqlUAc+P+UNMkZH2jT59QAbcY9RG3WyBmTH9IHVWzebHc/TW9QUw0cYjVcg6nWmUo4m
y86tXSeLB5iSAgligGAxvPBx1X4iJJBBOfLU3a+eyZRD543tldnY/wQmRFwh3Lu/x7YY/0+Km39j
zZgcvPxJksa55+EQeOPR2cCMf6WRWTUamBdyXZ4pA6dGR4r2KUL8bn38mWa031zpY0b4300sRedM
1Lvzm5qSzstmehTbk18C7PpuEZo/5xxzm3newHITA5Cjm/ePHp2ZKHc1XVQgw1zkn5Rqg7mbcz7I
1vMBszOORUkAfbmxkegBPI1ivCq0BOek2so+WiHeNKLQuIcW34OW5LibeQp8Phg89IoBZl6tqmH5
2n2mI2Gm2A8EqZ/ptMRqqy7Dkr5J5bBbshAqothBta5QHcJRZRqgJAvGxdfGyPE6dQh7ZABQepUA
P6s7DtpZ2ncfgOVZE5Z8M3+Lr2RCLeoVWiCOCafZK3QkYessHbRu89US2I+Bs2ujow3LvD+yu0D0
FRSgklnW9LFNvw7C9zSoEoD0DG/18q3fAHGwpq6XJhxYLo4qm7HkXdG4TGcDHhqrhmGUCdKYb9sy
cxA7xYa6ON5TDg77ND4VHaX7MtVMXop5EQ7nTz0LSRQvRvG8C/GIdz0MqvboK/f2DJBZUWIEA8w6
F75cTEmpevITEyl4oOsjzbUga35OV8Ah2oDAFWCX1nKvEMgQ2ElUiD7obxASJkOq7UiOXXkwEsmZ
+4QI7YGoAwjOtozpzgKSvUgVKEMBB3rrS3sQzG8gd1l3EGooH1PKukom1/ZoTeY1gTudezYjkE5j
3RjrJ2EyapjwbIyzWKXU/V18/kA+jtVZRhORjS4vTQJzlt6hrserjnmgLB9ha0QXFusl7iFiau2O
24otBgln7mS/FrcsoSzmqe5otqts9xzLGJF985wWFpLOiPBXg9S1Lwt8u70GGbljKOpl35t0YPa/
cU68WJidx7iMDQIUQRFzydfzhKPSXG5nweikleKVgrO8a3Lfw7qO6Mg+LwxO8jTBMieqb6DakaaR
lV8uAgyymAOwJQZL9fCWOt//pIAryTTAQukMXinD4rs48T/L/uzYxBsjqlCNiNOWTp44HJtqDEws
t5b1OP95+TC/Y+fEd5vRSjEAlFA5xlqZBbSJsBLXF0QzTYtafrW8MTWtNuUVQshGlzXSKyx/FWWK
WqyPQSQXZtC+hx3mUbua5/RUZBBTRs16/Cr9pceRqP6U9zKhaoxXij/HC5jbVL59JcWisiUbqhK7
XB6IJPstxoDZBZLaDUTIw38QlpHTo5nnxuyQ1SXWna2s27OAbwvMNtlP+229s3g+10NXrHNxSkuX
sF0UcUfZRZ1Rx3ouXcicS0pgaQ9cucTKSBDbV7J5gQ+5T/NckecqL/KQP9ZjIw0H6Xy47LywbDJF
KO4FD7/HT3p53RMMSVZjFCL9m7VRBNNHPqycQ/PUBK5LXesunS66mJWgwBpfguuRsBlk2ACMbQx/
DcfyrlAs6YzVK4dZ/G9Mc4S8G6vCxsZSkPdJ3XxhLx1byb9qvhA0Yk37ikolegWJn77rvQJUuAg/
/XmVNobiGNq4Hxfc7iVYcpiriMkEYX5M1d94EV7V8PCXK5dHq/9HYx3meB3VGDCu/zPsKNTbCNeQ
XIcsTIIZjoNcGE2lwCWTrSEEOK99MxOjAnsJhNDdHSOREicJ0caXUxBDezAQqSXSo0Z1Z23WY3GJ
KWBerdQTpernLtxGETFeesfy1VT7j0mnUn0NbMnxOGKlu//Jqb8CUEZ3ajUofEin3L4uWHPr/qcf
wcSs66n7QfqE1zioM6LGGwKo8KWB5uKUeIanRoA4/Jc6LIUBDZmsSZOsE74hwnwmgAe3fUx8TIuO
RtWZ67wcNypu3pAUmiAMV2JdJdZoxSW4QBoFrfDzH/v7/84skqOgULMzIThy46Z7ObBjJdaYT/wV
yZjxjD/NST7liPSiImtvXciQXlht+Hb3RIJOirAnd1Ar7Qlxoj0iVxc3XYLUbSWmLjwkKeSLR9QW
uIFseHGnTqwd9tpSI1xjr7Z+wlsLNp4FmzZve9PWuQzChRo7B7fACmFP6q+/5fnsu76VE7tSpDzG
jIU13T+VwlC0bbS53FsvERp972HAneSdA+wJ37Cw+QxYWspJqVk86CuK/EAOnIRFqxf2GsaNu75h
S1m2xaG6dloowxuAu1Sj53G2e6i4h2XtGMr7ag8kmxtrQRemcjOALgje4L2a0GRaf1LtoAe0JZcX
iwDYYmCzoLZbDuc7Yl5TlBONbs7Y7/p31rBBJ4pVC8lVhHKe3OlXto1WP0yuVyN4yNNZo3Ai13LJ
exk9svJWAJAvDqckHZ+P9S8kRhHenchA71faW7iYsFwiIhDNQVtzWR1NjCXUbMfiqUBXlxjmvfcL
ISt+CdRsgaL71z7UrZewQZPOFs+RXufXbWrfML67RYdarJI2QzhPTgUcGMqkMv+BVRz3CtBjoRTT
nSAKCQjmTjgdLdjXpM3lYW6tuRMp+P5cLlD2wp8CnN8i0YkDaKXIhF+gRAht7ZARqVBks+e+Wf/9
l73oLYVO8jVsgocygrvoxHgt/gDFlhRdvucJbzBP3X5+sOyFd6kWpUaq2QLFKyGr1LHBoHFVWKwg
GrLeqs7yhwjVGDgxbGGQfOLQ6DanzTcInH0mvXFw34Ago+HHDvBPXYIdPG7mFLyCZxFtojfEBb7q
+beLaFyd/7HGj8oCToMNzbYmqs2M9BeomnHg8Aw/556pfhOQH4h/CAVtfhbQNzbD3E1laJw4CcT/
9f8k8woemMfd/DSjNopa7Xu9V6tFdqF7rRqtQQ7Ga51JBhiddTBoX5BqkJB6yE+V6uZB/i65/CTp
rm8NBbpyj80xt3SBNL7+syy6Iu9sKENj4YjbHAqsnKbN+tgbiu+zA+unSWEroZuJ48aXEx+oDa7p
Gz4y1OMAsfbk3wRcfTBUkrWiY4M6n/OKHEQTD5CsNYDqGgmRRrFHlra3hRT7jtrJNgwuHUg9JgKa
Gn61c2DxNTI+KCD33TyS79W8OV5bJRuR0Cc6VElE3cRXMJojSkaQt54s24zZC3QOBQa24d501mTV
aAlYEwJVPmKGrKT5X5bxfSS0V0O12pa447FjzMOcpXzDJJJbKo6HvOonJiFfWnvvR+rRYMejgDqb
WUHItnsEXODfwddKKRtbRZHhlxwQURMVft04gxGzgjTlyp9jgb3PdJbrZoAW5AjX7Cf1gVxKeMWz
dy7jrExsspK7srjlTsB8CCxVssU620acy+6cBTY2A9Wy3cndEUQR1LbzBjO1ViNbV5jBxhgdKp9v
wY0rhJXLKcCCxykDIN8ExNCXPDS9gQvSmEW0Tdcu1xKYESpTtjOb+epEqjNME5PP0p/33KpwR3s2
hp83c8E8fdJ4+7GU5UPG+PscIPK9hrup9RvUHJPEPD+ot7mrOsII/4+e8K9a+DG+y9ocp5yAag8W
7dG4rTxzExI/wnrSaeynUg4Krk1vDAIzLN+jqgNbhh956hVOLOuF7brwsU4yMPG4BzHSua9iFfcu
hraxC8BKNDnZKLjVhygdOI5Lbpvs8HwjKb+NCRrbeccDyUR3ONk1Vx178vEhzJm9ikThJT2plJfv
NAYF+1B7TTpO4PV5Fb5sUC3damqt5yijUyRb0HDey69Sxeth8EWbHuAD9SVbQK+OIM6+kxD99Mfs
NcpQZ/nDayohAx2PTVfU6F3LHzYebaMlqbzMdGAI9QIRe2+IAvlIKeqmOo6UP7AoDbyhiV+leGiZ
HfkGCon2aCHqNE8qVocS7C725ij+nZPdxF0adP7a7hFN59ML5GBG64Ytq2jBtgmoxrpWkxU8paGI
U+Tm9BLrVVJhoQZt48IVI/G7+jvLndlFUijsfQ7l9jdTtqlCrOiXfCcF/E2yxcBbaXC1XknRDMTK
4z8SaeKIZ6Shhp1lmz5YU1/m1tytJO0qVQysO33jMew+wNCb2t3cdC0vUyGDeBX85t5fIGrTdXW1
ffNcnvgEcnlz77DkNKQhYaeqAP8++TmFXfZE7DeGztG1m6bEm87FpWmOJmTzelFZHpNbWiumYcOl
JZRPXcKh1uIZQKi/Wz/+X4xB5Ddwc39+KSCeKLxfFaXlQm0JNeEdiMIRwtlXMYm6KV63tdxMQccL
rzRJAPOvychzCcnnndywzy5ATfgJmnsM8sr3zvU5v+eWM0tQBkVgMeq8Tu5QN6xoFhRlqEtLA1P0
pbB0yJVQPOg2j/P77JzAmU2IL9RrxOlFJqGVFq3P0j8KExMygCALix9/kbPDJd28x49u+t5B4gS0
PEhEMk0B+1bZtlSjxCpyW0nWCZFStwGACrPxnwDEdQYKWIXkpP4j1PLaxFp30zSUOw+KC3FxY5eZ
odDeNs/O5cMVo7fsvy4KnDuc1MDwbOMGWyKzMBk7H33ev3ZTXEju45Z3PvIROyjRTenknLgcaTJ6
PUk7M3WS1Nc/03KxPze6xovn/Ves5dr9muXnFVby91oejBc3dm5Ey3fLJJ7QWkzzKf8zAnDlNEkt
C3P/pQUFu/uSooKYl7bwHr0t2ZrWnn1oHEzqZ5Mj3Lzs47Py9Cq/F0DZvltqH1h6zPNs/YlniXe2
5nJlNBXtD8c+8RhuYZhA1eFQkiFDYB/6ARNRLJtFuuC71tCFCHrTdiNOB1yQoF6E1yAzSaDj7VQk
Tf0OY6N2oMtlDGkd2Y1g0Yg9folFvQlUWi4MS0ktiwfyd+uxZU7+HjL6Hx2YowP/LVbCFctrr3jz
iY4mikhanvoMU0/dxImXgKUiWdM9uCCo9ryoPgf0SX0Z4Zv2jlUUjMpb8rPi6nkgo0ZXMS3XAL3D
3w7whBXaCBy07U28T88DW+EkekDzEW6AnPMRkEhluJch9xqsuOhv4KzWrsoMXsysddVbQzaAPQIY
4JQ2Vk+h++pFGLEkBRecb0O6nDjDruIcvtTaZXx+8TZ+IDEAMdtwhpsCacNqnvGPknsBRPJAA5Gw
5NzUv1ZN15B9+f2wfm9acL0MPwePnxLPX+U3DtU+IouXIeIr2UBwVISZwtxGjrYBRk6CVQ5W+SHK
9MKCaeazeXxyEFwLnaxyxQ+taCZeYJmQ86qM3BVMCeUSrHwojheT2WpKR9GBQLowTc6PH+qjlRm/
T+e/vH51DEcE5ifsaiMU/CwNFBxcK2hqfnnOlBB6ctOf4A74DRmHjiQtk8JbgT3NPHjQ9UTQGE6t
7opEvo2NqqIpZLU6ykIQcCHGdUU2CfmR/VBPLRJ3r3Ba0rOhH4Wr0RaiKjjbK75fKW11+Lno+oWx
AkPFgcvjTBiKcFAq4I+L0LdnPkPNkndYNM5HD3PYvbmZCukxy6rzOkbet3n+apVD4iP4hPZl/sT/
0xx3k62ValG3tujIipC7jQCHjqRz8f0K4ltPdfuI9zWoYpxZm4IcoGG2lOWV9O/OPq/rImCulpml
JTBzlnDt8T1FtQdleITksF85BDPh9kiQKARjr/wKjpxYlGYPah3GUXEZX1G8U5WbaIcAewuHKUIz
mj2hci96QFE0oamsmBm6/u09H1EA+5Ivq7DkSK69biDm4jWzSy3z2sq7eVz3Do0itpZsQm4/Gz0Q
aou7MjX6GzEh+Ms2A7hygEGjpK+Dmn0HIFhKNWT30KAqQ1UaarHPpvrZl8su2vO1lNQxUiq7Oc/5
X/wl5DcXVnxfhL/XbH4+Z1dZkypmVNjTAZjzWlNqPhCdc5NXzI3zBfMnlCVCVitp7DpMRTGxutIk
LlnWtF8I8XFKj7DMpCTH9PeHFq3/yQ/7pgeRaiJ/O/iUuCx6IuOydLsfUzGRnLPN38/71L9muIYA
D83FDewXQWhh0TW2YSVJGmBaJ8kBBk94k0HjJYzUnMRkdRhj4orGIHGmGjOyH0iWu64Nk9UvLsCB
CrP9pA8hBCp9EhyzQQAFSalKSGmWboIQuDU189npLzIPx/86DzEij7rHEa0MEpOh9c41VeRPK3YA
NSvD2BOO3gg3WK7Dx6Mo3L26sO/EROvd+Qmp0kAdjomXW/1yMZAY8ic1+bVAAcV9RValgXkmWWv3
xcMUkHbQiZ826ObMle59zJRoSon+fiSmUSjUnKZFUH7K8n55xcd2Jh1bMGj0iloUR0RYpupywXkr
5Sqnx3no/IFqWlM/+WJOW5RhcKRFQB1fFAkc/vQ9Bxcx3nNt10WYthE+UzqJ2fHpo/E0izBbny7C
gpEZNi06/j76hc5LpMcvUKB5Tp0IkE63QxBWnpZDitkKmS6sZAgc/YiW7QagqlzoYVMMXrxv1Wvv
Yf2OmFwmTgCQ4qjdio0Lp3Emq8l7LrsLpDpRuMMPGSj4HPzbPIE1CZ2W5uzdENVk3sN8nxNchsr6
l9UTbrYlrwm9O4D9PBKys7h3jEhje1QN5haiNvIaoybEzQlkPtgPBV8XZgVd6keOG9BV1dznx3Cp
M8kM8ydl0qL/3532eAFMCfPEphwDdLJu5ucS2rbnC4poylhRFJXAY9OxcA/cVbGq61ptYuLYHlFg
A3fTh/HynIVbZ2OU7iwxe/gYn0893OJit1hh4k37eZ+0N7YiWK90F96aG6Cr2c96VXCQQMUI12ti
havRP1vXv5lLQPTJNiRBq4vj216Hbp5k7Tj3xqALoYJZJ+jst0+wrakzCGxS6WxEUoVyEGkGQV+Y
g2WjL3lBAJNOPTUrkdl+gqJ8s+sSinKOrceyXTyXIsXg4HRVkiidM2FVbdYPmhRsAHf+FjmMq30y
gqOS2JCuPBRJEFE+OfFNx3b6T9sm2syTV5X/pX1mp45mN1oU38eA21C0PYhGTJQFAuH1U7ZzzUlK
pJmS9v1KROVeKdvCYwpnnsTL0ivqOi98iP4S3vlbOCM4MxUK9U1InOgWFi3m8HzWvXRD2UFbI1ei
Av7HGJYRugVsCWFj1Cog9X0MY0GLsjKEK6Mc2ZPesPXZsgFh0kE91QGGMgCalFdnayJG/vWZLruu
HEgoW4kY7iyeHGvjlhUl5uhq/7gtxlqGRB8wx5vbXU3dK0vDMX/GYRs1Xeos1l4Ua2itLoqTK+V+
/BRoY7v5rbWiHk0xq6bKNCGiE5SufL5CxNkfiaJ8UBAsTLfctqmePBtaoXYCoAOe4nyAN2Wv9xhO
p3XlHfn97hzn4EWrmVgojBEsH0PwjA0uWJ0jkbUNaLPRXR1Q4bym4+BwmYkGRGpaA3GX4OsYGqL0
nsWwwOB9POj2O0wEqDfIHerosucEdpj33hb/4iCggWyKnX2PwnpDJuJQz+brMFcUTvssZSi+/NLw
6uzzomBztSWLHzPmYQ1t+5652Wqlx2yjUccuE3xGJjugVwfmb+GNwA5Xzuo80eWKfbnYtMklDj2G
Wezh6rC+k6W8u/97W4zEiqAOBb0QJmbAdvYvYh/jUCC3H5IvsVswcDTLym+nzClJ5MEhjFfPC/DK
03AnjuZitR9Rhuhx4QxhaBYBrlgCn+JfS9b03dmwKYoSvO0aUl2ltNJfFztV9ylLuG61DJlr51kt
zvJKxokLpRY3V2o/Gi89p47jUTsWq0OaJBeXcyI4osRWaCk8wZRi2R6VVkYshO3eHSfhQqS+3CdY
Cn6Q64RHHaJ0dhiut7I8XyEit09GWtliZhQ8ODP9IGo1nMNysb3utTSF6JHpT6pgfXg534dfoFko
rj/si+VRlwAbTY1yh1ELCL6Q6a4roVStGVMRJwDF6Lk/KcpMJGi5FP5jCrV8scxVKeBj1W5GQYEN
nmohBRTk28JoFKo91EvbqxnhUoBJpL8pw4lp3Dw5DvMtlYhH8wiF68wOQRKNkf3/9WufUoJSA72x
zlz+OJf6FYyyB03kMgKD6k9vZUu0qlG/Ak91Lz6HaBj3FbNrgtywBHUtpbWtFgVsEDT4RJlorJiA
Dlg1bXA/s1UKZ7Eek0CQNHEC/xxusX7sDZZf9e1lm3KncWkLfgCdeLaAwm5WsNoc3HLG2woU1SGG
CULvRyk7wWuE6XOkPwxdFki+2tcvzfEM1zAk7TiaKiqxoktrDq9br1NusqFDe1R3ZV3PgN8D7Qc5
cbAYcetV4mK1MWqvf9Baj4XpPvXujbGOZVkC/rngjCKE94MIdi4bwhrM+HsSlozMILl4XOcQV1bB
JSGY23FGNZQ+0/9uD6As9KED9CylFa1xCOx1e0vwdHYiUoo5SJ/bN1dpT65qMLAeMqq9jOddx2hB
JVB2KTeYW3L/N337rcHEB6brK2kOompZH/dMEaA24fKpBi//oO2pp5xKmoPX9ZcZen+hWXZSZIXk
1OM5aBBqPjymB/9wKnMElKZN5YEr4FO/f8LDhFQZ8GL3N/JS9J5V1WDx2R9DX0slDnou2GuTA51F
8xbtt4BM1U8dJqwLMFUy8R3Y3MYYP0lxNXv65wX+g/jH6J7iN1psg7e2Va/PR22kU7eqdGBxbzNH
iFmYC883IIMoT8SGZ6YUCDJFeWBtX9HSNoyxJNBQqoi3441dSGE+XDOODdczZ6vA5Te5TqPaUQUu
bUR66UQiZ79OwdQLNo/VNn9GwZGBud2z6AY4uImVhyhIFxuQ2SR1ffd3YFmAUd1LqvjylzBFVnzt
r6q/VheEz7VvhTRYDa8way6qTk3eaINoFALimiW5PKC5pB7szea9eiwqpHW6S0AJctW8/HcPKKTC
/qMxkWtdJ6WHKGMgjNUhyq87gJAbZXzCK17SJi7q++IRJrJ7NniQcSMuRx6X4JHYXb1356mM/CHn
4ywYATseHr7N9i10obLAN/Ekfooi55amV5Xyh49/Zow2Mm5iolJqAH4VkxgwxRsal7k7RwgWZhFz
WXWAzQ/ODsfM3/ImuHzqzoqM2g0CD447gordzz/RsxFmYms/fJMyIZNrO34tQIHYuRiYj25OkU3u
lylHISjLfdwzLXbFtsoLkgPfBAQhfn4F4hGqqkWwTEjtw6sgr1YyaFXwYisrsGBDhmw5TD1v65Il
gNXFetHRG7DGmiTKORUil/g4FBYngNXDDAguxzSh85+zJTTIrpY7k6bktP6ZhdirXpeWreFB8HjU
E6YC7zk5ml9ryLCesiEMMv1lOSX+H3dbaLvBdLhd3C/vXnaSyy51m+0hmH6sWGMgzdoV7bC7lNMY
RsMolAme6GXW2/cACIazFeaWoJOcvYmT9o0hl3ZnGzwE88ijKY04lLs3eeN17NW6VG0AT2sJJdf3
Vrp2hOiVbP+pZAioW5L9NcZ/JfUIzhjn8c0tRyE7xVLX1cACgA2ZdcMsADpCptjDT8Ld7RA9PGa5
d7BhJXoB4TZ1GUie3UwgRLBpUZR1Wc3JdRuf52MH/5FY8dbev0f0VGxUUe6xpf2g4fmiYQgYt3M+
wB4eSls0aGm+O8+wm9SVJ7acPWdefn/mcE7fHAtTl6yNxu0zzQrLuFZ/SHnjarGL1WKZYkMBNJgI
ZKT+YiSyMf8LMykW2VnKHYDXYHQ9aMOmSoEt53TKQu7xTrsglm9xDJHOFh4oQPJnvEfX3lS+nRzq
MujulVbTbrHhJI2YEWZRFGSvhx0LMAqB8xBufvFCKQAM08UKXZyIUcYfP6pS79KUzi0C9o903BCt
fwtc5ifNpHhdetdJPhTfcc5O3KSMlGzYUMqXKNblqybzIW0lOlUNbQumkz+3+zt2vI0OWDdSrkES
+xXPoQ+VFGY0pbKdQa5Q0bKLxnJWSASISSqiRw33V3xeiyF7v1LBIf+sZK8XfMgHOuu+esrWZOjS
i9eygvKAJ50ZTabW0IG24IQT/ARnN3J+B5s94V1RBxMJsQDxuCv4VJYgXv9gF2dsU9AIOOpmpU05
XL78XnkTbUp64ZFa7mB0Up0S+Clnrtb57LclmcT2y0SuGIUTaVIX2AgxwUOPXvQnWVogJTocy00p
zl5TLCuKND7BAJ1Tqt5qFOjQ9n8h2q1k44odnd03iMWbVkruvhL+GEYDCyqqBJbshPsF6B//h91J
457ONQSuARW/lFyVpSf/N6P8zbSMix3vw/pcDf9bYB7/AX8LmVUBvt3NBzP2tmHK+5bqESQzg8c+
g+G1hovmjjaHFD+Fi3alJtvLJq0f0yZ+NFCQmX08RYQ7c+bWofxxpwTncO15/uEAFfTGKHYatv+D
Iswaa1uBOUlZmKhDxKOVhdt2hgLabrX3RS4r549xjG6ol2hcb8fEEX7UXb5nDGDkc65cpf7tnPHr
al7etDEzqVxk1E6NUAsci3AyiiOHTtOjIebH0pSjNGnvRp6b6UfqF0OgWpIcNsHWpcelH7T+MoiW
S+3N56a02TmLoG50iftzzCFocLiypWRVCyHvKwegjxC6DCoUwYfmbcOmHFwBcspXgZ6XbCqFm0Kb
h1CVsdVyD1zH/LFf1fzWL+3yrjtniTzhlh8l20l6d5XhSSyqM04+r8Fy7sX3Tf6JBeGaQwoqLnIe
rRssNqzi7b/hViui0lcE2nLg6f++1FykcAakf0YBbcHPTY33x5jE2ly1jRmjzIMI2CGO9ro6dEU0
DYPp360uI/xN7trEXbsz+TME5XQkL/H5d5JgghhLLaRKee0eWFp8WFL6ueajrbcpTw/V6cManfst
OBZ73NfCsfkJUI3cx6h3fsk6dXGsFHv7uez+8/S2lTMYp6s2FAVbH/acUIQDCsANsxsGG/tMGXKG
7BXcAt/JADVy7KsBdvI9lg3+lfRlHXVe8kPux83thCvAUMeL1O2k9KYZD657DfEZElonc/rgWpxb
GCjFsv5chew/c+DhJ3QMNb8ajHnYD4N5qitt4eN+p1ll+rN6n+rv+x1+233LFnlWg88kZK5BXmhw
KUdycGpaCUIV2fxXEQi9wv97uUS3Z5vj/TUawDbwoiAzeE0ZTChF2jDCca8eS6F2uXdZ+V/NEqWP
AVuI1CD0Ld6HqtYxtxgKU0PIOfTqF+nLA/QDqfO6d8mX1ujt8L7YZOqzEjBlDZnVT9rc/guaV4WR
rYjmDXtT+PtJj4UT+fixF9XDBCjPOJ5gVD2DrbQkb1RyEonaHdsjtht7MUHe5/PU5PLpz6/XmAev
E+xJauNm8rW6w/ExVQswVzOF7e2X5rVTkHxbUIOfbfCMteawDtioFk6YrfrQEE+FWMNpsym5zgLM
4NUnEYBScNzaUAmwpgyDWbqQ6HlWNSkowimBDtrPNKy9T1b4ZpyxVvNLqHytXNCSejyOF4MvYz5k
bDD7I2kwIsKV+nOzC6kRELZANygxzZme+93ZFFVSydAQITd7ItghS8AJlKJxXkddIzCqahVfdgRI
495MITaF9QHeHRbJz3eH95Pk+VhX65Fn3yVw3g52gKwEkYZ4LToGqA7O5A5TroAhK1VzvwefHflT
Ctj1Hm1ulYLeuQZdGSk6MS7HsacDmVRVHQcy9bj8s5h73D5oosTlTCCkZ5DPSWbUxmgGJpAYWjwM
AL9twHVsDdxeM6cOCTEKAoFXJSDIyXHooQgB0+OxBJrNUa3h4J4h/USCERQc+XM+c2ZSj/3EDFkU
O9d4hPmjvUwPISYZaHcBGzy+JbBraBsg7Omweh8FhH946yOjiFVLodHZkaGE+8azqlzWVUaPKND3
zz8705DDEsUHbo2gBAr6kpMnEwZrwNsDoV+CG18jXl2JZzTsr+zSu3eluTbPbHm3/KXnQhoezjuE
WbslZMs2WkE8qwSEgEShikPrf378GJJ1VnXDmsfBbarkKQc/Rp4QCLsZ1cT6/voZtLlHeSWZgkBg
ycL6jvZ5ReiqGFT+TtZPyKBqenaSuGCLEjcjPQ7tKMUx9kZtA6qQb1EClXocIms1Gk+itNBkIFBu
wKv+46fjDDk5cLgvEZFXe4lkch07++l4NcQlMp3XRsqTAdGBKumITVepJdNJx+2B8BxN892RE+zS
nBDpFw+FnSxjYfqsbUrtxttgmzopUzgGvSDPsR7sJ/0B+S6pP7TUbp+wWibpT2NDbflKer1O91sP
LRRc+9MnV+NqAgPQg8oLg0nmxRPsH6XoIS/R4ILGO0jDuLcPMBzOA8pAOGULEV7ArBmFIG6eKs5e
MVRq7BTqqyg93eLQVgN2K6CVEhxAKy+OruqGI2GsxzgylsQYqIyebIz0efpcwS+6n1ThceBzpoD7
waWa6yx6hZgVlR3wRHg3fBSLAlkdwY6ucb958+uWCsGSu6hd5qhIph/TXD66DiqxeXeBMFGbbb5U
PcbmIst6rqc2xmnMISp+wQm0+6TT1B7aT/WykLRVPWQDQ3aW9UmGzLAnKUEYBHNv3XMnjjzYYFM9
OLnVOVCnNEXxlx/lRrjc8eHNjZEZrVna1753D2a/QixSr5yZ78FUBdaIulvkNKzwfMof+z6jtoQF
WOAu8K0OgGfLBficysqzgmaaRBaTiAesCtGXGGhDhxR7fhXCiVb7zd5FUQf9bm91UQlklwUUt+cm
Tn75ANOU05aK0dIXo7wnNvXab3sKQvNWZGkKf+2cYpFVvO/b6COIr91LbiwPKXrD4w+OevhyJ73C
dTg0/Ex/KpYnUBiE/H2Z01OHhm7tDQYWpjYeCt1I4Lfam4uBuWqHB4cpS+9+28aKyfFn0e3zKfIM
okdEEIn/6iMiKbvkxJqZp6OG6r6rd7DemkeqlBPxvCKv7fQyW5vtmf/qYzlDiKc/FYO9fOTAKkD5
r6N8zggh2IFMArFAzD2vNTX+D/fEhoAWUPX4nkoHHUW2fYU2lOuN8XwhFiUFxyltF04RwNZExVaD
wuwfug8EMxTlwIDv3vP2tRiYqUvT35Rez7srd8opCMQX73ecmmKspfPWQJit/FUJQxExTKMQg1xC
H6aqO3yzvAHCisEtXIS6xPYjsnWD1TImVruqcbMpT2DTdCFOZSwUU0ecnEeu36JUe4OlkoVOCESj
8Hjn4Wkh1BiK6y3qui9jg4G+0Iyz8tfe9dfgKsaYZDiL3uO/ZrAyIO8p5V3TuJ0Eg76arGGXF/Pm
jZr/SG0WHNz7FTwCNr8lCvuvP0ViUCk2kzvsKEP5bJsSQZI6jgce8VcT9RDZmywyiztcVfs84Hg8
KukcJJR3TTcQMaPtXiyS60EZEyPeUGFUhvGuD/qyYjfeF3gTj8rgzQlf9WxYnMOKyLBY2xqI8zHx
bRvZk42pw8jUZGn8gJ6BWp/p8oeG6bSeyqSxTc19C9+WZYPy7HJmUGLLnh2HBoAgk2qqSEkKBk/4
NyIAAKPQjilgbY4s1AzYpDcI+Qq8AORez2O1Tplo4kUMHkoDOF22dt6M1pK/N1cRFbivlsREDkNx
v2t6+CH9UrhnpGsrJGu+j6gq3yFzQThV3mHdeieluLhc3zuyRvi5v5yrIsDBkOZuumQbSUdUiFm+
I16r0itzQlSBDJFUmNs6yZ2GOEfgKK8iPqg1Pk1TuVdYoolrilJ25j00nOJ1k+WczY62oE92v6HW
MLtxf0Thy03ZX/loI/5TXoTh/fi7xv9J84nRskfVCcLcFR1nLa8AYs67H19NMQ35ki+1NfTpWlrg
3z0ABwXzLKNq0wTffDEMkfPQyOVhgrOUws3x7qmkzaiW3TMCJAx6dhIyBHjIXQuAeYDTacjysLsF
rF+uvLiisSEQOAGZZqbKAJajhOik9aYvse82eyxbGFByr8uV988qd8a7xEs/yRZ7Eox83LLaLnNR
4ZULv1CMME2tbIQYgRHMJJLzTSdpcZQmB33kmB4MVPJNJPhYoVWV1JSnpdJJLccYzE6p90Avz0Pa
CJnZ/7aWt93ZvVJgwDjjGin0wu76OYMN5KCfXR/yjcQjZTvj6dspQCPv2270kcP3njQLnusykVmA
Q+nPp3rliEoLMDh4ucKdZvCzSNx7AIeRzwvgVPXasmj1NEap0Ujh7+7vJH99f5MVhXTsuLYC+0Zh
QryPTjKaP4IwEOXqzWX6Fo//Xg1a2JM4EciicaUnIKfhB+cprQozxPcXRSsGBR7T2rkCBlMEbMZ2
zhj67aqTolLU65ctSFly/5ZjeafdtOK3H6QVMTprDBWAu3XK7ajmPEvvUoakuUs1SLvsR6Hp64vV
COMnHJm0ZzKyqa5X7nLUHzaCFchYuAbgExr9MGnxgO+mQYFv5kB84ZvbQo6TLVqv4qqF/6xEO8eg
pFvyTdbgNwuz46zNj4KiSe6a6PeZTeNRG7nvCY92F84CP0skblqLsMXhGjhV/wZHgxToBlmL5PhK
63LVAKgxjmDkpbD4W2Q5mQeBa7naTagXu83/t2huRH+gl/ZmtHWeTC1syOfz8biU0WKMjvy9+VO3
yw3bGlWgbuROEthCzipQCoVib9vU1JdTX8xGzh7TluxUuKSpIclupZOfOzjFi6GAvZA2x15u+B/v
OxFM9DjMfswCuWtVduVXT6pn9T+qcobPKixEjRKmZX8tGvJnDwz/xzHSIoePMzSeJfYMmpxZEVua
7clTBPNhLhOyiRTfgNO5UbdGgkQeNSxy9Jy+m/QqbIGplUE9HF8w/wdoV5RJ6mqt1RZS+QB5ci03
GBS1JOixqEolq+46NP/QTYg/BaKHNZn/sL8IIVCfNZga0lWaNRrnsVNeq1DlES2Y1IIB6HCpYO3N
logc2sQhzaK/Rk+2BNApVE5k65e7ymppuMrsSBb+0xkqg7XiYVa9bSk55w4yrYRYjQyodeA2sH03
VPYL6wbl3jWx0ywmDbyt8QbDEjWaB/Yemfv+PoNR2y0pHPVAi4Bj+U+DU1GvlZ1Aon0f+JtLSqJD
bnoO1QT9zvR9w8EEPuxZ4Uy7PR6o2mvAddREorKLoJWOQaagtHywZsdhg3FRiv2UoAbjIGh/W1+i
8hLK+vBvHX6GmOgaDpgsYQ+dX3RdJf86FQTQ4o+W4WL4FPOwqMXkMJn2ARopKyBizCwxPLnumj81
hp/6SHv1kx6x6wbsvrRL4xrY6DiqKUqlysx1ZL6xMpPcfaPurNFXG1cQNuGk7EURaAgXNvvfWYtE
+w8yWx4VEKJLnmUC6zeCBb0SlUOuP3nsgCxN87hfjyuuee64t3qyoCVFh3EmZeEZXxQWxvvWWD2x
lUbTHrnAe5l1ObmeIj2PUqYkDbYgmNHPXDLc3ptf5CVVTnm7j2cd7mg3stgYwuWJ56m4W+gU3Woy
wRWmyuVWlANdXQXz9qseKj1Jq9KyoFMfOo9BVPeZCupBnYkapKI2SN/E9uK/lthw5ImM7ynIg14b
DKPIDfS0qBJSzcpRDybUau6kPansE3ZvHZmt5HZ21Eb+RCul7P79ngPZkvil5bTktI/LeKwNa+0x
MJ5tynUAXWNNYRIghMryymvHhYQD4S0egGnr2/MD38h+k9SZeAuPBrycPMUsESXYKGF5VU2EYmHi
jhcWmJzVNgnLsPpqz7HT4OJe/357pUlt3SSjf1f9xeQBJusVrMW5pLP0ahFiLAUphR0cv/GwfEAz
EccQHkVfYEnNAP8W/QMf35DzcJDHRPRjm65w85U/bHZbBNtrWUg1/f8K71zpWiPX4O1S1Tz15T98
5CJkwvaQK/Z/ULitte1pvgWB2ew64dUXKAsAHvX+9RqAqEFPcGxKB9UO2hRto0SQOn9STHFaaxIk
mzI9tVVP/HD0Oj90kHf0bNpXQ9rj1aQ7VgBzodb0G3AEFCAXWjR+rUUVpLfLwHqcDnD6W6/o6NPT
BL1CvRoDvlynbD9vplGn99/nsZb+xu5ljf1MoLDvtfJN0+hVrewNYbXZC/DOH7X8DpxbRtbycjJK
rPpipM/Rj5kzlmdXm0j9nl3F3x8jPrwVryTObYjUNes23AIwB6lxLD1DmCiJpLupPbPYhQCyMJMh
+GsNqMA0Fk1C4mYRTqNWhtKf0I+Og5RFgFOdmLqjto6Ek1SoCBTtGD6q9HAxvNzk4p7YQH8ygGxp
r6Fo51KVw7FG6SWC0A0AV2xvKhQNFSSTjPjf8HngU+0tmWVJ6MdABtW/18an9RElIFttbeyvKe/d
/syB7gsxO8lJj4BcuuK9X75a2B8ujEb6pL91QDhoQiOd43ijgVxmx3H27ZQzMRJ3HylipuM8gJ3y
guz3ghS4ef+U71FOVFg9KtJMPsJre9IpPaBJU3P1vzU+gjXzHD9POij16wpYRJI8DFAK7cYFoBms
55EmKBsdLCU+ZfIq/TLCXcY1XtFUz3sun0l6rsZuDabJ2tl1M4N4hXvVhNAFNY9UgoiXfqcYUYJa
BhQq2d2MQ8k45fbc3DBRoVSOTpzzikcWOlCIn6brBCfXwJG2rjLzHDPZ6VNf1tZGe1UQ2sQPsQh5
Hl3eaHVCeeUE81mGRDmT194ffXqvh3zASzlmf9texLqLlUf0vEu2ae6qYw8nejTDWm5JqfhZyqUA
QsmGA7u40qX4v0ouOWMTQkPUNbkMTLzF6P9LWG/b6/DFJIVvQsfBkFl+1MyAFGPxLLEHRawdg3bD
cpX8Mxy52+UZaS3+Ars1wjds+X7iXSBjPdVIdcjFZnysAUidvnZ0BXuoEHAsXPmefzX6N9QVY1CR
XgGFHpkHu5uH/A5kPLoHqdRNgjHOEFT+zaCd9Z4fyYsdxz9zOB/eEktdWG7TfnDv+sYhbjTuwsPA
eHknhaV3akoa2hY2gRTOYTT/Vk8XcmCHHfqejc7cSGiaIFR3Y9q1rPUxH/KV5RTwitEQQKZq+O4R
VyXoUwx9dm1eEX5aDH2ddcv9rXaU4B5rBlPk4aj1Ix04rxpBs8OCrYxZ2ke0JgKwosjse9F6Uoil
vRSirC/zZlqzokwP6IqqIp/WGqAowT6JJ9Pbjm8z4lD6daE1FyPw3ZykITxhaLyymOh5nzUaEEq6
ksFEAKqNkTVp7fKesqBTXa4cbIG3y+cuSzkSOtj+ab+AImKZcIEyg6YLztpNYd/pcuNIQISNMWIN
6g8M6wIm0EOM7EoLiOoBFHV/tC7OJsN6xsRrg0//XXkEDk1ag6RJuhiNIJzjoOTV3HzqzkJl9xT0
3vUSkomBXk7Tv7nmGjsfWxPdhjCQQBNz6QKQATcwblR5YKadn/kiE+mG5vccaRr9UlUNwIkGyMUm
JTYXhUw/pvzNFG6B3AzCQg7I4Lad68G2EUGLefRJ9GiSw37Qn85dnkBWRk+98YBTrD9biD8QrJaB
j3QDL5MpuYZv3qYpn/rNq2RN9CY36QthzBBktRFVSD/vLQdeTN06eepY31v2AmtLYZy7XaHO/2vN
i6/6/KlBF0n+F6rxed4uMvqDf0c8RE7MfpvrsRhkjYcR9qiMnl4XMNbKfbEsGIFVip2JYGXebcBv
PUBKq5tzVH/Ra7vDQD5N5HBRFXu58UrCQtosA1nualOEJ2OZIupaczyNGY1nBxIFL1Ki4kapaoEX
KTR2gbDxipvkYYOFH1qsjdNbRPzG1psDQD2wHJiLchhh2y5Y1BmNiNCQKH6tZn/gyD567PTrXR+i
pCS3D12Xnfae1Rf3L7cE9nHRt4E5IfQgnAjEhuwBo0MuOWsKrVVrC/iehRF68VhW15/LlmZ7ax71
PWIAK1GXBoD1zbnbsEblqPRxThSo/OlBg+Rm+L4K9GIB31zZjGYX+rjjJQfoPlSVbldrGFG4UpSR
7oVdmNHBaqecfC9MNVYTecs4BXWUl+BlSgtoI9+f4XGXU0W/FcPtOT3KjitvZ3dXk04UCM3UOpO7
PeH3DhVWSDnL74obeVaF3OlnQL4gY6NreVWAwuH1kL8LKhDAGnqqmGxijWPiUQqHu7haHrNWbuif
6A+Uc8C84t4kJPdW0DwzYQZE3j4dt/t8IpsclJtniGBs/sIPMlW/IcZ3I9ce9ersB+MijxhtO7IK
q2xARmTgQskGhV/FE7CLijBUcB9tBJgD1KhFQaEobNMzoDnuI6sRjZIsB8R5ddymPsOghasBWLQx
YW4gm/Ihol51cpDhzdKfQQkJGOr3PmOzZCvVzbPApPvj+g5wWKoXiOKz3XLUQ2srpuVh7wpfg5gw
F94DrJYs2a3KXc8Y00ZpNeIFMwTr8JJdvXhevb6gAZM243+rvPlwsNTIGUOC/Mh+lFGr1DRpDsUR
6VSbLGxmsQPqhMsHvQyqPFQp1CeaGcWotdrRqDN+nhpKH4z//6gN9VfhjdRbLlgj5/o+P/p2JJPn
zzkn3nL//KrbFtxbeoJS2ti08opClffZsgGpuhxmOOL7FeXHTJH7lHWO1q2mkAiETqr0KJKPQmAa
2tWUt0tY0aCAVUzr73Skscsuyr5jiT1K4Qxji3Tqq637vtFq1BBjk8gYgOMg1lYYn0nX7M0zfLi2
gBgOR2RacaOARVHdSR2QlD8CCY3UUcKWRAGuP6nx0VWj6a7Q+9jSzeFOuzdypN3OZMlDMdQ78DGP
R0T3cGlXp0fSEu1zFTAjtntfZwijnI6IUipMG7o2lGdx69ZvdUHy5+9T0X947pClqF+tCj3jCtMU
MDh7nJ0bpH3mJDEaSaWjhMpzg8iwCiw8kBn6+YXciwGJRNL8+PfJWF87dhMZL7M6A0hcofmM2LVj
+zKRDrPq374PMkt0E3KyREevvgZINKDSiQ4pGhrAbZ/CD8aN7iauwmc4Vy58maTKXgyIojUKnrI7
4awTYZy4cOiAoRYHB9MSr9JIuC/wk9sQRLqHlKa3sPt4u7fNIdhutxbnP1eOR5OLL6fKFa8s2uTH
Q12/I1wF5XGZ9CRK3NULQPNU82txtvGEmNFYM1NKojiaKnSdVYcpux2UQaa1OTAzxru6LQttDfQ/
ZJbCXpyK7NzlVoHcLyq2IJW/tE23iABONpVU/4wYxapnm8la/Pc3aDrIVJ0JQ4x2DEx/1EIj7aDi
3GsJJdxJkZypu+twRJu1cK4/51g9GkyZufa1nYwQSoQmSYPC+hnf+lETuHwDWn/Vmh2Aoi3Taerl
4Nqo4AaUyAOibzbKQiLJKagKVt5A0rf6c3X/Ftm7DNG9G+NXFRzUyX3F5btlY1C5ApF55TAKEPFU
Q11wEDYySEOLklfvcr50ixdow3UjExcdD2q1CJGBmr5DlMDMhMhE0FEQAbs/1khuBBtIK3mvx2Po
uCBrKPmmL1C3tL2O+KxZTIlNtT0JcAxqVEvvqEjxCDhIyYNJpCeiM/59eq9VKuJS7GpnliTLYDl2
RBcvKd5y5e0Ia7W8VpnsORs6SkmzsTpfagFlWMic3dYPE3UNdVduLU+sOgVV0ZkkBGj8T+kKAwYi
axiR5KOS0L8RrRfpxGkSpwQAxJfRFeRKIGCigCnbA8tLZVHN2d+aUpm9BQAGuytQvAby1fk+W4xS
iagCv1egFhhMzO6WIFc9SkYW3GXsdeURI5++X7A0da3KPlE9J1AB+ruQqMdhCmMS7JM35Rn/kG6Q
v0pbx/jinMkfD89+OOwbxAtzOriHk9RTfXyQ/V4rR/zwmP/DCawANuiZzsy9xZt5LeOIVDhW8edf
CIUoIJA2jgnp7i4Wro56G5NTIf+WSvG31R0FMfi9MRSqtqzf6iNTf7xGaoYq+KN4gOMAIcUU3joT
Q21pJlLyn+Fa9B0l7E3+Va3vsRlOlg9mhU1sG8I4WzSarvL1WTQXw5ZKdu5ErAI+Oc9AQHvEZ36q
uTX4c4Y/IAPfr2WBUZeWp2Kj2ZEEVIDzhkcVMECpF4u1bke0PbZXDjkpxAGOflh8wa+cLsy1L53V
jFMAfIPZujUo5pZzsIfwPKrzXQo4CSuQ6CzShQkpBuJv1QuRiXAZCjCc9MpWXiDbM9bYuqxT46Ju
biHAqHTB/AJl7OUrlYRGOT5PQ60XIRL4JlR7O4sQcVSY/YMgFgJFYP0qLE2GP/3FdUkW6W/eyM5F
PsrnNfMyUH5OuzuHQRo4QR421EgbrCZalYEYoMOBuw5lTddGYDROBen8XFuB7t6IuaiRVdUPsxTK
Wo3pGgvAkfdEZ/R7HVAkuhHBlkddawhDdqXj6yxyMVu1iZXmiIei4T6E9a9J9v5N/w4FdLS1edLq
oEE9sggh7voF/Kr90ScWLN88CX0eiBCGBH9r+UfFz1OaY5nJuJ5S9puMJC4DUcc46RoIIUjhNmer
Ki1o2DSh22KwV5z7Cp77BQhge1EsH9Rss+5BeT8QRpngG/ypFKZR7XoKS8U7OcKtj0eDrRhC8lTz
lE/ZtjSc7CiP3lq5jp4Kv5p9/5R/l63C6T0bBxD3i/R0k/RUi1o9vKLecoeWiulHPxu6IAbhQ/kx
VQYiEktwSJZYSFgRrpQsDOavSQLSC/2jp5dPPpdW6iITLbMk+4ptUlzRQNp6qOWmXPJT3UZLEo3R
LhHJw8aRJLmCip44AOtanQHFWZw/zmpiVFdgHqPwCkJaiZDM7gMFNKBOkcE0ID5hh7qfWc43Uz33
KRJEtUWH4Mnv3wym/I4LtmyvUNX5XeYyOXTO9O2m79n2+MwU2aBrRGeHSJBg0plBrK9uX0hGmSXx
Qg3CNw2zYmITQ/SD5r35Rc4WavZYK5RTEihjV3ecYOUq7w94Xsx2byq4pe68MqtUCjZHHuvQTCKn
nbUCejgZV0bzZ2Cqd+TaUr2H0dPYDdbUpnX+/YHxYImWLfjpjaX4SveF4JPerB7LQOYcMF9Vpqra
aZqMP6FB6CBLfeubA9/h9LdWunyTye7gSz6i+1sIcwjZnlNNuJa1viQxGmdNFuYrNIT6g2hiVrl3
4wuz/T8BOHcA2HhzhdBeU54ZlLDNa6lN7zhCxdQKB22sMqyRiNmpUtKnbxwo/U97JVgqWc/OhQjF
al95awCQAppG886Cqq3yiRTrFWc7jQGAFTfCAHPB+2NzuCv9DawChXE5PYDFj23nIb7FAjbJUoh7
+iy1A/MZ4v57YYhO+M5wJDHGcsvz6n/MLadJTq0aSRqVmXSi69Iw3dc+H4Z0jW+MZml6u5gJJGSj
9gKfsrRj5tmmWhA419tYOJideax+0ci1oFJIVNPZhwcbo26IH6fnw20UX4aUkp/LfafgnGL0C9S/
Oy2XqduzW9Y6OKvw5YvpCVnwcOremF5KMnfgphfiQkDo149Ap5uQLHiEKz6G0hnUktxtaoXAmVC4
ARN3T1TOEYncK56biuiILNMv20vaug5ABHLmUWFNykB23VVW3o1FYWY21aArwlAjCZp7H/ehRiy0
Jr7cnVO6H2nZeY3fS/H167yRuvUt5eYMhE1HwXiRafSqdGbhSOItelNCw15eWbQWnrwbOwEhpHkF
zLXebbvfKmPwcdBRDMgksQGXnu7bbKOxK8RakLM+B6ahzvsLi9GO0D0amR0zfHl3RY7Hb3ifZnRd
ef3DXe14EzTLpdOrPliLyCzd3OSfZraGwnzRrEjReXwmaDzVENBihNA174faSYX3Fj0mJ/mOZjLH
84ixwFNttVP6r9YZplM6q6Ct0TXn5Vj9juTciGqLd2PdUcm5cNaRr29IN9+hdNhScIg4WBRS+QiD
S4ZY96iS+F7lSEvPX/+n2LLgzsAZASmVdn2EZYn25gYiym9ShhAkXcwSJNc5+qu0RzrBBrD3rhX+
NAT8Tl7pnYJgWhaz3PFweB7MhavsA5XqlyZiiRO1xjOR2r+JvMfaDY+lzu18iUDOJN4L10/d4YSk
rP8xwq8bLxwoaHHipzTjWoork0LISLAuGfXRgPa4OtpvV6RV7q5cUUkiEBJcO8NYyytEF6wR4xjU
P38CzuOzgmhFS5CwlFr9EUAn+Ku7I+fcM8g97u3FLWhDxz+I6LD4pjEcdgAygsTylDUVa82K8uRQ
wjKiS7zh1nnaNK/l+EbyPmeSpBUW5Uam7Q1zluUCFJ8U5GTOZ6f7tacBR1xn/zVM5m/bKdf3v2qO
Kd7eqfF/iLCmoAfsMiiZ7U3dKFkouLYguQMsat0Gbbqy2pzJLFxTkMi2t4KpeNCUaFC4KypAKmNF
utKEHOyjNzD9ayFtTkEV0rL3LZzOu0iPenCIAhvn+FVVGw8xhq0j8DoNShfvsjZ/D53sEGHZOfpJ
FaPDqgC1Lk/d1zG6wNubQmTJARyu8ZNE1C//PR5gQ4MxO6NrUoHfnwWz/csHee1jrRi3/WJClVOk
Cj3h6fU1eH2v5wU5I+8LM6XyFt4N/tas57Wofe0CMWmAE1ZqmRUSc9IKyC8j/v2qvqKGf4UpNaIQ
VtmAt7ea6sihJWGcp1aK6VbXgZY7jPbONGHbPrO1Kwl4uSEvh9DxAyDB16gx0F+LQCTrsQdHrEbD
WJF7QSgw4SLFbpfLPVa0d/gKMvSHUqVs0/m7ge2rqB7aFxjB/i9FdCyDDbeLM4vWKQc0uEa8eplA
tPmAAj21f4gJzAiGLLo4Hzv+NDraqJLdE6+Yjs6anEldxN42xvP6qIljEx6vaqfRdGQl9C8NvUOz
cRfLXuZYnzOtSW6tBOys3eHZ5Ua5RgNdVk05a3lF3L/mi0pLWB4vMvXv5eWODbFA/GTpAuxu+Oq4
V1Gc00B78y1sB4N/ExfWaJFA3nfPl0KWZA3ViEQPQOCkoTCGuap/ufu9aZB+ME5LWJJMot5LMFXl
VYMUmAsIsf871WIsfRlG0ZF2qn30RpknAI4AHf97ef58Rpq2YuyjMg8oILM7IMKltK9qxMGEow+l
1JiqasIVXvfzI1exF8xO+MVm3Su4Qz05KtKXQHa/3dSzkIfKLb6SgMHCHzj6Utivz14tQzUMGvpl
qnmKv4inGYvx2paX8wi/l/fCFGxY5E4LlbtQY7SkDdr6jVwmBGI7ehjNZON9Yjtg9kiNvbiyfP4c
rj0phHUQMTrbaU9Fw9fmaLLrOKyjpHRR42H9+dSkf53przWPTJe47lLp6RSSNUD4HpujD7W6aozO
rWrlQH6zoiifM3/rNgY94R4S0oisq+WT3xoXiPcJMcz0Co1Zw+pU/EWOXgEsAumPa/eRWRck7vBn
Pf3MjiZ8q6AOn5AfGwDmhNTFijYuMxKWCAuOJ2NKVsCDgh3Af286mrHlTuJ7O5aa9gbt1ZXF2Zui
Nk3XPhxK/FBrapjvMRzrtLV3x9wPJGNEfpVDQsoGTgr8GHO5lVU9w0cHRYepatUZa4P7ZYJnDTgn
CEB+XcHAu5FtSPzNonOA0hDpdgNFVKoRMNba7UOvWdNRTCQci13wAf7yFWXc/wvamiSmz4Un8XxP
7dLEbGKOLEDLlWfV162wAoezy+tOZaDAro5qhQFWnPB8yNMgD8moLKdo13AHGG+LwtVNF68ZM71u
BrtIsRjqs4sru1S1YLaQzC+qmZr+eenIDR5sXIX8XRnY5WC6S+kmO7spfP3ps4VCV0bOI1Xt3+e+
rIsMytUU+KbOMeRexh73jmF1fCvskG/1Ngf/u93OlabNFfHAyh/2n7X6Gsbm46n/sMwOXFs/O8ll
mwgrYjXHCBZG6+Tqj4ExQEdElzfEqABLYTrRRZvUHolJyWt0hfPisjPXlw4kdpwuWgxOsjVNrhCS
42DDPk8vJ0wLWwTyVTrKFveGEVVDvk7Nj2s6/WDsIOU2x+IERs9OHmCZh/A9+8hQiexgLf8W44lD
bZfmOBvGK2HLmiezHs4oWmurAgPKAsujzS6f3A1wscfbZTVcXC4lCnM5AbbUUl1qe4Zrr3E8G93Z
HAnZB0Y8GtSuVJJY2UNyZ9qG77OFHjyIvrsCzvmv3u37m7/eHuQQodpXf16yMrABuPchDyDF16Su
Ab9L6ln/kqQkPy0X11W1yueYnLypQGZ4QLjhhid9tEJGbchOGosIlFrpdOaA3SjgwUZtAsVMGQ+9
YAfpAzhhIMus67hBNvExMmzTPuoWqWM/SgE8pMy5ZZ0krh8WuAo5u9jS4LIVOevCaxA03B7ZYZbi
hSYoxrw30B5TEerrGSTsSiZlaEr+Z7siTzoexvW0JC8CsxnRDSPe0BjBpSE3Am7qsIrauOFqaMJw
svghmoo801MNAEIxKZalL+cvPMlC6TfOT9X7YMWNkyi3NP4SAKxxJlIyn+biI/cF+FtNl0cU2gge
E+OtzPjInsEmO5/s/VeG261BtVCU5qDZCWwVlrjJexFgqmXTRGnUPP5uZ/otJJoc7xexJJFCMYYk
xXjCGcuYESaIJgxOBpGt16Sxv/JmcRzR4JCdpl9sGSQ9G7iwqZFg/Dr570TtMIGjVdi7yYN4dI0g
fnMi2MI0doBAsupFHqGbl+6Xg/fdENaiqY5Hi79ClvfmjEo+ajljeQjDmqD4IwbtAtIBjzNoa10O
GbOcJgAp7DOtgq1PlTZjUY1AAojvmaT1HNb/ZIYlDDdxpX2k4usTp5AJy30+bJofCkjQSKSZkuY3
zYR4WV6TxJSgTfhAk0dQbocyBaVUFX1Z12cqZyfT5H7wEryAMN0BOZyuXySzY/6CvAs0SoWcY2++
+5NL84wx1v+IqtxqhJ6DvoClXcBH16ErDvL/qtsrTvIAQ+iGbYHVkclC7WN7jLslv3j31DqYuRfR
DY7NPYUq12B2HUAgYWfjhex0+uh1Xm5ob73/WZMtlhnt+WmZpBQrpBElTjIkSq+1SEt87CgtR2XA
Dm9YU+La4qlDFeQ41NXZdBeIHikFtHkH/ZqE1oiGj97tROq+tpJpdWdxXhxdZnYXZovg0v5dLFLo
jxfUxJndx2GVJ7iUxiL0o9GYDVB+wVpIhcmoJ1bJfrExN9CcLssFGPzZd6WQi9e+GONcyGwEIIsR
jnzLOTe9+3TQqKUE9QiwNPZd+/Qtzbs6pOWnhMIDglNvxaFKqAkr1T9w2Ztkkpi2KyDhkU+x1DT0
nr4FRbN0Fqt81ENh3ra5x6eTxkkEhDEW11yZxuAVUYdvZX0ihzeOSCjk2Axt816RU2kv0q+zOZ44
pf2DMeI7b5NV0cODJk00zkndI0OIOv8YxO0JDvyTQlVdmoLVU95oP1wc7Bt1pk/2UcoQXU8yaUzU
ufPYJ6MyiFKUgyJy2dfjNBWdnFdMqFRtZ4Wxp1kh6+klsVV+mTUjc4RSdJN4H5I2mXjASjnYpp9j
Uv56vps3ZofcQrwSNnTQ1XRv5pxGdb7fVVERlpF9FTmoT+lYm8Q1oVJH39dD8QXlXhidO2QmEQTK
zQF2oD8sspJVo4LIwKsIixtXWoqXoCnzC+Xbzz9s3g5LsWmAir/3++aDM8196idIsq3B/8er/Mg2
B9MyokA+UvEEBcPr8g7Oi07oNayQ5E1hiXUNjoI7zr0fcSSVHjslyUPJ21kukyvPt40pCQ263ApK
NhpVwFmasCuxqbzXmUqWBf9hDNjxfsrj9QsEaS/lpob0LNQWgapRMqK+GRTD5y4Vo127t3Z5Leq9
rUfGLWFVulhVCDPjyD6ark+YWgTP5hyx8iXetyXnpprRP/clYhrFpQfaRoTPtZIi0ID/2GV8hTKe
FJz49FxZ/szSjP/075+X15xkfSeCQ0euhDNCB+5XvrnQ7I6Sb6+pS/gwJ3LkH5WzRY0EvQxvysiV
xI2uYpVLm6qDat6ClCfDBqMI5yiIA5gm/SvflJo/7f7AXqXQEwQ0myISpBFsyL0v/9aBdlQKhspW
yi9p0+kA9gnoPgIdnzj60s7CyuvE3Oy5j/1qXGmwinmD9eMYOED/v20QDNBdK2Olg5/k75eB5mTT
6+KcMiso75VqsFnrw8hzJcHYWH+RlpQw6FgYk77XOUjHyOjVaODVDsMP2g0CvrKzL4PYeYQN97nk
R8vDmHqvQumogkG/DKIvjgVlin7F0Dsm0WevDJ2HGHxbRYrN09eHJASXkXuGWBJpLn4EJcKYl3L2
o+QdRI8/KI7OVh0Nc2pDe9Ww8YbzPCazvBmutfnpFhKlHmggFAIxKhZrj3qiAgH+P74vfZ6CqsBS
L+Zs5K7Vs88dX7Iq6/RVZFzl2k8yBUKaJ2INcvD7TM+IFcZZWWupHP8NkuvNc7FvNbBVANFOUaXv
ZglAY0BmkqbL6gS1SWquXmLgGgstlBWRYF18OjLjBzw9oxqXS9ql3x/CrktfhJ0JGV6rQnE67HYs
3Wo40RpWoOG2Xl8B3zwc767Nim2R/qyFMy3g8LTeOHNXHJt3XcjIpnci8hCy6cZWnm7M3Mh6Hr4r
zDbRrbhl7F8AmZD+Y353+AnoeOVrhdx/Lt2YISaF1tL9+PMDC3dKhVYI1clfjwLZUyvObzFnIoql
KosWzaTGKbrxYF7FqrQOgvwvorkqiBPektY16DPF8iSmRdvtoQsy/m6/17L5fGnrwTMdIZMZGnbK
zB+eH6KwYxHDY6qe3Z8uBlklXHo0yP5mkUurMAsOnXgTFGCwsvAxlMHgCR/QWBn8Q65njo+qvzlW
rhuOmAkPd/7bKBsd/ASiChk+nqPQx+ZUMRwa4e8is+gABJz1IKKzRt7b37jXb7JHqMKJ0LGuPqPL
J0JO38l2PaMiR0llciOJX4OKzz7Mqpg9+OWGmsNqV5HhL2OoXAL7XnCWIOVeHShlLvztCsIe2HZ3
wT/4M6FU9LvvcktgKmRZqULIDt7pp3sB/MmaKhSwdxTCwmU/C7iRiiHrAAMJP3PpdMsxBBLhzemo
886uAh+vob6XTmxEmgCuTgS8fDieWC8dPcFo02MZp+q028+hDfH1wbPYLJbaKEt9IsfFWIQFbQlw
2or8qkd2kQ8H2SwzMGqtomeciBD1oKuFEPgeuh6IXEBlM0HdksO16lax/K/HdxeRsqUZIqBwd9FL
7YqkWqDa8w2gnFAuZbl+JOj5Kr+lFNln7pxDHkXA61M/Jb9nFTHow9hRZWxTznTVQo5ROF2ROuCv
uNModNY+713Kbmz0uyJ6m3LemAB5HbJgmvKNczLkx5zewsqphCZ6MArLIMC6tW9dkaABiVqgW3fd
0LKWEQcBenAWg6MHOvaCkNvTft7y9Kn1GUjIwSuhz9gKOFMn4JapvGbjxv2RMgYLy0ILL3q9cw+r
m3wK8erGcMnR4BJuR5zD24bBQYbmtczSrHFnwQwlaOn+okmUwlOWtsgqIrYBwvGsvyGBAbO/p/Q0
1wy/YDcwhDOeri0CrSsuFsMOuoZrGdAN/h3wofGpMBczdg5fcNobU4y2tbgyMPRad3ZsmW7t1Vrn
UY6rT8/Ljbtn0G+6jcZ9jfHJsduKCE1J0Ztjtx6bieNHELGcK0xKvD5t4FzDAJ9wY5LeBFxUG9aS
HaZgeIbrN6jg0I75WXNKPyN/Uncz7Fh846FNGO6d8ZukMKojioj0UszBwi+pEbvFg86sqnqWuecK
xFK1omzrzSt7SilGL11ki+VGcWVZP+b5M7fQDaur+3Gca8rJ0W5HT+UZHWihUu4Ss2FgPuMPey7L
uEFcSCDb1rK5kXy+PgIwkSKgXoy8zeGIzCWULUdqJg2Dj8X0+N0XKaL3/iapb2RIKQo9PsTpt2+V
KJfMwLq/GUnjTzpowoNPxRr7N2iMYbQ8Bdu4RMGOltAZeeUbA/hQycYxIhABRUbmBEtVHy4NTbUn
Jo6aqhOLPBNWKErhbVz8rTZFFlFZ06A7w1hFYwODgC0JEQAFxnd8I5wS/j3erN2fZhtN4+CYZW1n
QLUCWplizeI3mCc0Fjt2+YXM9B/L8ZAgCPdacDwJi0PooUdF8YYQd/qA47Xc8iI4ZXLf+nkJrkFV
IeXeSgSOpFPln1OwSyNNs2AH2sfYReouV/8OR3pQT4rIKEW7e9MIEbCNmbNRFFr4i1aarnQ+Qnre
7ijMr+d2J4qzEvRYxm6qPYsgHfB9TcwoIO6WneowlWhkr9884XR0LrizfqoEdl7fYJvRPS665Qd4
mYMC8jZjb6W17Q/4f20WrRHeMAywCmw0TqqQ8flbRZC8uit7dEwTrSb57kmOOrWKoypTLlv6wbz7
RjysABe7uVou5S8XrHB8jgNsaDlbPP9WFo/MeLlvlr0CxueAqEqUk8ljW0TgfhJMN92YjkQ48AsG
Qp0GGOSVD5ofvNf5CD8BKZPekVNZSxyGtE2xG4ssFcEMCCK6eECHjeh10mrRJJy3uaw/dhisdCOn
41dx10rKlKELBt1E6Xyz6CMcPDqeUuX7CSeJPFaiXqzY+U/+1I58lY4rYRNC0uLyIP2XwRN0Yve0
oCRafWqKJIQkBvJf8j3l9casOYpDJEYrxKnAFVOcAHwCwBIoGhENYIwjpW/KysqRHli5dpoUcPnq
qnpxKAYDOLw/SjCnH4XWUJkosY9R78SL65MYY3DLtioGKcOpQdWKxq0htcF9rYMZowbqHeNiF26j
E7ZmSN6tYnUhwInWfRIBFuukKfaGxgIafZXzzPjH0l9GsKVZPh0ewE+eVKmFk4zPOIhn1O9fXAst
GANeft5Kx/gk01FiM0TVpQDIBriOp013OxtHYtaPIn9EnGWNHcmpirDZyuQxRkUfcCUvS7hjgYQY
znqQwt4Wt9qVlJ+qVtBfR1835LWFhRHHOq4x5s0tD83NkhBG4hREQUkgucymlQMfqkiqpx6BvXrY
wuDpm7/2o2C2I1BbI4rIZabFRwWfCapKJGPf5wjpOpVlzCSfKofDDvR8xA+9QQlj3SJGWfZsWvfu
C+v/mklmMXI5jDXDddEO+xsFkQ86Pz+xq/1HVTw6v1+Fb3TIch+ErYesOCgUIqNsmBSghRdTvkY9
pLYF/cogVZfgHIQHDDhk7uBQk81tR3k1LvS6mb+gYH6GbVUr9a11Lc0G4arR4FkrjtH/mNmCKQ5D
UUGh2dbYQ55m5IJfu5l0QB2LmsY8PIzxZyumSNNLDXkoIg8DVY6FEdGCz2V/ndjLtp8f4arwAZ1H
J6knP5uP585md9ZA4FrwZ+JrSeX6E7BDuPbh8imdzGxWLekHa/gZu4uXnbbvhmjhK3Rlk48GbayG
CV5Y9A5M7ZHVrWp1YmpDAIrH1YryuJt4iuurDB34dOJKotGjzL2cD/ZvNqrwSzh6xtIzdySeGOyN
f+WL1NJZyMVa1cKq+vtDKn+l4hQXug060riqqwETeHl16hrJ8uoIdiqDfA4FyloNwqzZUpl6qiTf
IC3JPbKVkZ3bGWtzUUhGHNDwlqYkFA8Yybh7p4DDgTQZtjZ6xxoSteKP0kpDpPIn8y4Mqoy1qE2R
QzzDElPxyWylPT6mFzeOnr+4B7vyHwaWpocfnMVK/q4CppXldTRv40ZHcftR0Yth36LrPMWIOf4+
yE9H+l39pShQ9dezrhtrJoeJZMbmvCw6J3GMCcajzMNFP3JfKIt5h0rPSRFrteRZemHZyk+fCL1a
k4uFtTe6mnxv/fUgJj1mRRoXAI4kSgQ7QxpZAlN8F0BZ+Uf+wbjBb33VaicARXOKMnmtfk3bqg/T
Mf10CuzaHjl1CiSC5GzvNcAq9XGrXk8ORMwwVASDXKqOZGV4mlLFPv1Grx9qGVsg9eI0qm01rTQ2
T35dkOT23kNgN9atglj3FPsEZwQ9vv9trWYp2xTZsv4wIM9bf4pSRW/A4m3RTtwmqamS3Krs9W6v
KzAKkMxL47KQb7giH7wlBZVOMQWpg/oSfz9N+5uPVwnhNbc+DSa3A0OIDz2XIM4DnGM8REwWqaZj
XX/tY5hG9m0WI3+CZ+X8DSjcIqtCk+zIwZxewKdnjTAdkhOK0UF9cjvAX/fDW1YnW8P2NHNWZf1N
BtzPYw5/5rQoyv7KulTaRft9dIeLgvm7kLqwcFe1pG7X7haxIDpQioTmufCPqLEGDhQMQ2AJJV+Z
IUAw9BoRFBtbM1DVo0eVhVKNaPTLnBf0+A3eEVjihB8ZDGcE6muOOrG/WG3OzNUsX/cv+qWBAzmz
e20weJuIWr+FOdG4w40SVhmfRS+hndXwkvz8qlRqX9pvxuGHM6wwKzczjpFbv2ZoqdisqhYV7nMR
JyAociS2IvbnmJUXNLHL8/M543w8qtC0qMVQjsntUT3/ISSIKC23i+o8bBOLyLAqhkjuD2vrntai
be23cdwjmvwOg2jE7Zsc1S2OId5blRT5zZTuEl46uKfGGppbG4vgol2Iz+AZ1pAjZmBXosGHIhhE
ndUx4Y9GR6dW/9z16PbetWDV8WOHRbsqFzdYbA7o9//tSbTAdAA6K6MLSlhrpmYBKlh/+yAfCRDP
hNOuDfAVrpjKrSGIbl3HjJtkFpwjXDp8JHdTqFB5FkP9m2/ctL39daB5YP29omAGUsqBEapQAa4f
UINnT7tS6hgtGy7oAioilYZdDHG/h3m+F4Kgvl1D9C2QSr8BoZnrkA83WrVIvMB+qk3YEuagLeDA
IxqaJ4hv+ucpFrJsb6SZ1Q7/wDV9J2QJJc1RHy6/sd5Ym30cO55Ot4LgLPgBw+8AXtIqq1YTBckP
SDtbcnNaBFGkIPF7tMrxrNYAZlKC6guxDdMLM0lpzO2uIXWGFnsy2qMOQcWyTtd3ofxTeRAmVbsA
2qlk+eHSe58PoXrF2XBEXIxZhYJkBcdk9kL38m2Uxth1PI9etS1hlZmSHmwF5RdQUzTH7PzW6YvP
NvgL6rICUb5Hxtct2ZLIUSgMaTT8RIoegwDAPjr3kdCB68gIzIyMV0kIGs9C68GZ4dJpbd3y3RXV
fvlXthXE6l3NBIaT4CMymDNRJwuYPi/nx1GPLA3rEsJEmGLFglZEscSVvUYc8tEwp4e5AId9AQi0
qVvyOBp69dGZTRNKHxNUglyRT9KTF56oZi0nAftPBkRpcKyFh3wJafSN0/tYQJ0U+D7al2ab00RB
MaIkNehrImXdHcnjzJGzmGwUCpdkK9hHPVpiugkXe+f2Z42/FQwnwpFRrxM62QFCt5AgaIGFMbc5
Z48v/2KIfWlUJPqPyZyT0dDy1uZAnBvtRkcrms2ceq5OnuR9JF4GcJ0NNd0vBDBPL6jt2GH97kfn
ja7CZ89FWO+eBPLkZXW+LzsV72QC1tsqSf/FMTQp8yt82U++1onDgBz/Js4J2LD8ggkuqlrkZdQt
Pm6dNQ362tpfKa9Vt2XARHE5zRpcRblYq0h6poUk/2N1nyunP/G2G0mghoa27lIayjLvTBeTc59F
qiiLfX7kCeeZzukAF2SzZAxmq9Yft8pxkGw5tzW9N01DwVEGY9LP4hvbPh/7e83ISXyEX3w8bQ+P
7kvX4uw+2SIl5OUVyMzaEOkej/hCCz80LLE8P7YlrEV+B+csr5dylwZfh5By1o0M/7lj80RoGZJX
mBIka9yKcMquDn93OyXnmTSzeA4A64t0KdzPc50k8pB7u+w+FPrYBVrnA+19WVMcoMgIzdnu4iNs
2JyzGcsYguVLOqpYdSOPHxcyZus+zkSrkQ9ul/jk33yN+F3nLVSProVuEuS494wNMev4sP7hRJxB
tndpYvV8OO7wfSGX92fyN1vHctyDOL/lUhO8uiWQT4b/1kHIWdkPBjxviw/GI8s10rU/5SeeaUEo
8tD57s7d43PmA0dM868fISkXRJdGNFL58z7A92UkHh89WKED5PhYBMMwvn0qoFMUuy7pHpVTkcgg
U9gEaINXSp772kmJe2rVOCgFLAN5Vt7jzrwOqiDeZ44JZOABlEH1C6PRaUFdnaBiQirwxcc5MM7r
bZR/01Os4cLUGLHApg4OuowBxF1VzH6EoxQQjchuGJaZ+taUxu1q+JvNMkcEGWGkf8LtAyyF8SLs
fNZr4SqdrFatP5yAielvlz8fRV4pUgoKE8zUOdVyIluC9acr6+SmEOnYHufAX266O/ZmhqtULs2a
xts+dRk8R7E35w2YInsUd2wbWYFRT0seEB7D5yt1ZKXH+3XmECfR065LTDMh7wpWKNQ+dl1lyHXL
HlFsr7NaIBN/wcagQj+2IFEp8ywCn+LLvdxV8Ke+89TfCQCSW8DaPz6jekCHtjf7sHNwIfj0dJIy
cNXk/Ei1PbByFSFCn++uChyvKVhd1SuNazuW8/GqO5RiBVn9joTfSQd+Q1z1k+qxOkdBlqA2tdot
Lk4cz555YrDrycI1RSqM7Ty5RQCQ523ZANfgMSggGeKJpjpMoKfFX2jnN9/dOhdfNvkphNrwD/I7
tt5pHvJrM0Y9FM3t+sUg/YP6b31T0eHFMCKtEg9svQsKIwO2pMktlRaSbC5XaUzN53ZQnuhyR410
TcTkDyBN8xHRUs7vBOBtjNpLRQGh6m3wmfhooJa3/TPXeHy7CXnbDdRkVFP9SAPA47nuv6k3jqn3
TCaZ/oyAb6UfQ1cE0jXhZxI9rK5zvNsPhjPHsAAOmwGtKHFsAcLZye4BtkR2la2PMoRH7kiS0FHd
F8cTPo+t+duGC60nNiYAycvi7SAoJ5bKetDh/QqaGOemJyDMo7adyDfS4gp8n3ZIDW6DV+LLrOSP
9FFTKpXT8dOva4Z1yNYXJVNaIIi9FX1z9PCRa3WyZ5sWpCl7Cb8NkuI6ePFTXaKTzg6qFmtk8ZQB
b/JgiQtbhXHTaqJ6LdtwtatLPPw0OYokRqlDxpkQLshq5YUCvMXISWAvAsSmdRg3jhCP5B4SlAM9
S7uhU1nrqIO+TSXCvDM8+b9ZNUjuQYd2EyFT8elv5DymMmWkc/5rzz3AT7BXPK+aeoXGZ98ajbpo
yWsGpL0KShcg4k+i1V2lO03cXYdH42rSFd8DdHlogePLnyoFb0O8gCzKDLzwcT+EXqYa8Y+jNzu9
mExc0TnNcbOFSbvKOOONfCl1CLFnttKHxP0B4TAL5VgvQrcPPwVy493NqfQq1fQ5XU07kh1GTGud
j5qjqGcahXaDAg9myByEjmmEBKjRinJxu8OW+YPEUAr0kHYiFBOcH1syRoYPhC2xRAK5XPYScxee
T4+jWlO2VWaoUKkTnLkzd72e1VgxXnT89sWjvWceuyWd84ph6hVsJOSjeRxTlwm4VI5EqCzAd3UQ
+DSLAe+wj3chRlRQOUKgKWyVUUg9LiimLaagBOOnvgoGA5eSIs8dTcWST55vzqvL5B4wE0CJUZIN
KZu9djpbiH4CO9ftiCMGsL0/i9JRZso7UjAmeNkx4rMqtnlpX3s7AY9p3U7BMlvzlNBt5ocTlI9L
YRdX5XjLH3K0hvufZ5WLyn+IpNYI+BmF7Qh4Vs0zgTvqY+911CVn4Z3Xq8fCDhqI5zjmJ2cGGFMW
A/0PrXS0CzoLVdEICXHfBZC+PF8MQClDmpimyd9FPtbvZGynCf+iwKudPGx6zAUdH0a1erA5ib4n
OzYR7ko/eMbJ9ca86umC0qXoAK49EgwXNBsAphhiLtnOl4B+E4cuEspw0t6/nikvz/egdA4ebjHU
9aFlHITEzBfLqki8ola0u2UtaXtqZIjmk0f2u8Ql4INrm6XDI3D8SWKZ/ZXZ6WXVr7bYrKlhdV9n
r1kA19pTBBjtTnbHYhEdh8N7AXcVXAvPBNx/e1CmKeVTEMgNAn0Kon0cDkCpOHxQNl9aZQl4Dz/4
UGhFhH1bbqYDp6NR5nSyfUSjHG2boBDJcnPUaXRTz9BlnEDizQ7Um964H/Gwi0+sW8VvtYZLogtz
dqhmPW1MJAvXsxoYk5kXgoCJRFacdLQmDD4xJBKyBRc+dJ0XOy4pX7p7AMmDBKqCgQdPO+dZokNO
gKvLtNrX1yQEJW4SstKt8GIBGdrG/EXpsfFC2t5lIg6LrnO+bYjTheZR/hlQiUCPs80bl3UKvgyS
eDlHNQE/euntLNGd0PpyRvaQSEa4CLuvVuirZKmAyGCRR7NH9evY+mUVAMy45lSGnsK5fII33L2S
wa6QrIXMvD8WWej7QbEReMzkDdW/A55uivmxmu4+c6krswiO4k730c+VYMiBCjJpZqZ8TGNRCB4Q
M66rk95gz4dwKKb8EyA4y5Uo0U0ymxRBIx/dpxcIYmEJFFSuBcPRBO1FeCCuSMXTq5GWUyDsk9Uc
vApp2VMnWblvfpiYhCe2r1GE0hvIfmTuxwxKN+soBk69ee29Ks13QUiFoInulPogMmudDpo3i5xj
5kHRIzG4pAv8fJXHMY7WPPtDXW18/EVyneT9T3U1BVVS4f2BLOxpsVfJ1Gip+VMPKS9LaHYz2W3i
k89PLf/GHYqPlGXYm0cZaRcY/mDhjP32wu38Mhek/e1UVOpRROLb90l9VXw6Z7pdAiTHzrClGK2H
G1tFrrFzgdwRJT48SzmF5h63D9rd+mwdv/FIeDThei+VRqFwPuE+eGDDDLOBLNt5H4qKUFL50nkl
Lj6SMGxXRpSxsKpyD+BzDVI5GoSoCSuzwfGJZfhKrRLDTsJNfAfXTPxMHwPQAJPeYlS6ZZUw2TNM
X76QNaOwX4CxxFJJSSLiDfiia0o9FCokCLwJSGlWcasYHLhFDlL9CQVrPIftqt9H+OmsuZRb2JY8
KdnodE/gGkk9hRG38lNNT8FnrDtxsdtvJXgzG2ThTPMeqIaRxklkpp/haM9juBWhbFglDehXShsw
D3BtTgOQ538zGlaiy5egb//RV6fCNWw3Mkqbci4Fyii2v3xIVHFOIMXwMgRJviha3ZHxRAE59cz8
s4KESgHKhMBegS6CpmtxSFaoA5JbDTtTNRg9VL7EGNnCffSy7tBUcpR8EPdoPe+maz3NeU3Ga74j
E1QolsyJf27+3vFmU05pRX+lzHvIWZ3ekfRwRUmo6tGfPTgFP5WloJDVOkBR0QucHN46j4QPxmja
ZJxcYTFdOIgPlVXzItZvb2HQsuSfoFwB6ikZvz357pRirXP/mZnHZ7bgbzmN7OC1LsCtvjl0/xSH
AbIk5Y9pKdZ/Ou86kmoF/kHcliq/gjrSIfyivZ9oLXb9DyqvVIaZzbBZr5vuzVQVMl6bwJAVGUkd
Dh2/NxufB6NRwkyRhAHMMKpUwCEB2mzMEh3w9fbBbKVXu69tu0Ybfo4EI8KUU49XVgwfVP0SF1IS
7oSRWoGdC1vyf/Nk3UrQwv8gmFr9+yeWE5K1Z/ySkydmKwRCPg2uvyca+F46zQHaAZixp6bZdk0m
oumFxY8m7VVb7YB1IvsZhlcfVYNjRAhMbJvewf+cpv7Bv0sZf4NdCUL+5BIH94ZzvnMN1w+gU/Nh
0h3sv2KRrA6L0EqioyBpB60xuzZKTAtP2WoUxbYVrGRMWqYpnbfNesTLnjjVJOywnQlKIJQ+09Kw
aq1BDNCZif57IG1sKWWkM5/eDOSMd4+7yYMkzfsbiaYIwf9kaPb13IhgDCDLK2PboMsOiyL8kQV0
7kEiEVIY6xtOf6rGLHq7yISWAh9HWd+6j9bn4JPQA2ycYhIfdZckeohyE21viawMaz+Xhpq2rr/7
p2ob4dep5q0SjUlPLJtFJRHzBSs5cpO4NTF/EHNxiX98gEBjksEVrgB3kIXmO1p6yVyWtOVmMXra
jZ76boLVooT/JA4slf0zP5YAdu7qfhlqHprW+fDBu8tUljA39iPd3Djn1XMeMcmFLrrG7yOn/Jwa
GfwYVIn6cO7EaZIJwafJmluyV5GDz1jyzR6C0/LNamlGFBgjRs5y3Ehz5uwOIpLnYrHFxCkxpNZU
tZIMzibdZIjawvDbLngY0Obk0zmQ9/rXXvnKTg7VBSmKMVQ/2hl2ZAL5Po6jxr7JdD5X5lhiAmNJ
gsb7+movoOEAy6vMJJd1OmrrbINp/whxt3ZecjteukhrtXmHxTMU3mTorztrlG9eb8e7NU5/ByVx
L5Yx4badkp5D4kcp5b489EV/HsA4WONVQlbc2w0ZpEfsf30eN/HeY6kU79vVMMC2qMZM39TW5IM6
SSzwYS3zIDgzG7PkuABLf4Fven04jK8+dW7mOWJEMbOdJFfigcw1BPACBTHqF+vnSLdFdVHCZs7D
QXSnZULzjPoo9TIrwqEOJDeRmUcIcpxhvFJV1Lxi6M7nDFqtEEzTr+dzKmV23SO1e20SCa/D/lcI
1oDU9v9+Ha5TKT2xN5eW2sEaokWO3xkBP22yfyJ1cf/Z2mW1fDa7bDPMcmWLJmAf6UoaW6osl5f7
MtgMov5eImOnnRVi4iXcrAhCFpHA9NoDGRCWDIZ2P4gwhhiKP4Ej/KHv8BB+D1qfobw6RdiYdn/x
5SVheplkW4RpwslEi+aaD2FGdTEBDiiWi4q6LTwOupUaWpSNUEscblKxGr7M1oV4rB9ArRIWVqtO
tWxAcxVlYzitgGSY9+B9lpaYjtO5dbWMIQMLuhvE69JGnL193P2wo1MNWQlyBhCACCPYVbtS9O3a
OeS8NY87ZZ74ZY6w+kAiZX0eu2TSbK7woIvTjJAo30GxBErUb5Cip5/c7rjvyJJkG1L2RbSM52Gu
Gsx4t2N9cTkYM/gPb8/tLsWewyEg3JUyFtc6V8weGcSB+dSKPfG2f5Fbd5XO/WTHRIP2vGkFDfra
JH90nj8M71t0zLf7q+s5Yuf8tyx//n/lOe+FHsAMbWDe25y+Aw/dgA7JV/dszCRN3d/Tp0JPtzxS
YgEBHKCNwd4TJib4Y9U2gfk4YGS5vk2n4zAHVS5UABy72gpGN4hAXOWJi4xEtcrm48yg8CY/Pj1J
V+aP/EDDX4VMA2syEClwgcnwlHuMKfnXW3KHOmNXYyvAgdX4HCp6Wo+2F7i3DTtxBYKweGQz/it/
L7y2NOzW55sShLibed7gSPMjh0tdLXYqU0SF4ME9BGgpOWdS8cxg3B47vmpoWuxqxX0iSmGgIkAb
rMNkM+wr8EU5oFpLOSO3oVmrH+3y6CjFkhV4J6WFq3giUR2rLdUo9YjCNQTrYTVlrHrBHjCx1VgN
y2KeeIetNJmMFXOb6Rey5zm+SyUClsxhH4akPL8iNJkbVZqR1bApt6ZeyqCHF09JXm5DvFWBhjPS
mmZ69NC1mUWv/LHocPDX48gnWnsFpKmsVNmmYN87q5CkonR40NXJDjDR6qOZljLLMOZC6jKfObA3
eyEy2kY54e3ySs1qCkswcnmSHzBBaQeYm33Y6vgi3/s/l8y8wWTHp/bj9XvCYT2DEkRDZfEu5NTj
k1z2W3pJ/l/azIf2gOl9khAogrB7wuaHWJpOZKSJLP38xS/0qNrJcWDWssd2ri07aJLahuShW1eB
PbIDnm2wH678U4V2IbdgTIYvkSkIMbdFUU+Z51Xn5KBD4r6vEXim4YDrnP/hlM5QyLqsaRPCC3XU
NRJOq81xafHx6fzqWPri+8Hw8UxpxcLnsBM885Gy5PD/hTTGvAlXc7bRd5SqJNE2H7zfCwpHkweA
V1+UR6zans21In4N3LnbuaZa7UT72gINOg092Qq0GLrd1XMXNIZZDps8P5n+h+BV2MECzqGJkV9y
apVVtg9hNXgcmzCvVLrnfjze0GX/FlvtP9sYV/aie39AUFUd+SbLcjvGhc4A2XjMMMXcGqOcRFPY
cePUFz30xC5cOzn5TJbek9Ixum4Wo2SCbXzhUloCFGSpHjDZB48RjSzrlEnNdjJ1BkikXU8tU482
8X2BkfxiN1ClPXaFRkuWJkONqoeSoriXYc77gVCicA2y12vLHWzvhAq+7hRhOqOZTJ54sERYgcsp
9hajX7xGEn6wa08eh/uUU3BRo66PlqvEogKD4Vy2OUWAZuvY+SmuiuVnPCm56bjKUTVkduA9bf6d
tIt0+8Bxl6g3VN7a5ZniDRo5b5aFof1AAHGGhPLn4/S6//b70iG+zTUeyEFI8Nfxg+r99dvlR1JX
CXWHJiOUxQ/m5p33aoUTUBlrK2WBMu/MlUSn0IO3gyQP13HFvpVxFqCphwKsyTwC/dc4OjXTo1Lb
YZGW5rXPG8kV8cGSV5R14YA0hFgWk5/ZBg+HE16sOL37TvM+tJpJ3BY8hOh5BJt0s4eeGNWsm+AF
GS39baLjutAHixQixQTvaaCaxhV821qfNCPPVAfPVGqefOzyjaJ6u+nJKzRjqGkgaMT4AZX63LVR
TnAgczEE/rcLa7aBxP5nnloDlhOLV/eIfNofCijbtyCoEFdTrY5048dCczNsGw0U0iWcicXy05nA
qLwp23C+1jM665ebZiPQoQ65MsDsQsWSYN/+xqnH4ZNeDtm3YGetditvjj7qgYRGb0iuyGMYp3K0
4iNP3BdRThVmUtRZEyigx73NekIXR2SWk1p2T2VvHn9lFU/HXu+LgjCettdEj25snvp7kXgRB7zJ
GBEep6Ds8Nr7vW+DG1bRcAmQzgU2wycbXjSA2kA/G5NralVxwWAHRLLc+P/Bh/u2MFs5pEmnomcM
KFqx6I+lFrvQOEfHihLIlD8U0k46NHJSixB7sSAK6LfE56IAMuGV4cIW53t5xUMEca1tBWdIvi+m
9i4FtFX/SrusnY4aR0Yy+XfQGkWds/DPSDJ+027b/FVQgrkGUNpf3X3L5lZ239O8eR0y7AsITeR8
gSHPw6elf7ye3xzg/v/CKodIic2ecmY4G/1tjDKmCpMFnjGuCetFdARAdhvE8ZFXHGIY88gE6ROb
Ta+jLm1AAM8oedO4j0E73t5H1KWBFDzUcDve+QN6og5Vx9CzTeci9nlvddTNNZCPWmXGUYya+n5Q
LkM7IRFCPKNFPYgwOVptwLkgD7j5W0vjSHUskza3C7fezLhWVMzlgW7EGOdMD2Fz6bnl9s1oHKzo
qCPqrYLnHzOe5bwB+t7UYkbdbUMxHS80IO7/+zjMFdVBV8kE1nIqzIQ59vkkWNmzQwcF8F4CG9u6
SFFoaOxumZUuhCJp96NsA3nhZOEwZQfltmTsTk6acmX4jiDMxLWQLzaGkB557P2Hokf1qIS38pnn
g2K47mNOWMEiFNBmhHSkvB4WYRYg8j1YfpW9ifAfUmVSFII+UBKXdWCp1Srwkcohj/P7MlTx9BfZ
1tOG5oOa9GkiM5FKq4CryUaBaFqQyEfbd8Y9AOs71ZOu4YDW2Zq7xm66OCZZmAejcTjLhfbjY9cQ
nyqPeHgGcGCy7PXaA+jVJSd6d8pv1yxZZ9vTFffsgtoI9gUmNs5IojBc9+R7GLXzutIQPwNgb+bk
K4HV01g/XLpTapMzpk2Bw3SlfcLrI/4g+0qlXsaORA0WPuBMsHKWsO9vdW0gTVwXWfpyn/oSrHnY
SeOK6nVTCLR0bYhbi3AUmihtWYcFbXI0O4bCjcBSusR86EL66Blmn2DrzyH0cNAUzeVU4hh3jLT4
/vsKdJxpYsfy+RjRDAM5+1LUVYzRJd27sE3GUhNYVjpGCcOC2h/f917e0fA1IeXcd3LycscecPc6
BAbvobpqV8jsfxIWmuWOBLnjw4Ut9EL6c2JcWqayqoeUKTG83YCk6dNmYrH4qKeIKfttp+lKeYdc
TI93barhqZIGX35gQnvlcDpkFtrX1Kz2JuUvCSi3cRYo5hRFLvxZiDOzqcfsLfo73KOYcIdDhkn3
QHIL21bMlmgBbt+iPoOWXsa+1JCBOVgSA/bMEtg9tee8WphQlpgwpbMN1yoRosNiOLvQ7GolACQY
qp7tl0gOGC+a3PE94MMsH5qoGCIqWDjKphJTOzZLTLpBbF+kThwEoIKGxsE4ofS7oWN9WKhO287L
wge1RutLRyWWNXInd1LrwXO1TtUICTBezT/RYSvKlYWQErsYzZ5kE4QE390lNGu5znsYOvYaUiFa
XxGqZZPC+SyVkrnizEG+YbPz2yN8uPrGxS8FEVXKZ4FxyLEt8V9A8vpr++U+ZPxPMH2iZwhbywra
oLcaOW+rjBLsJu40anufeGKzNXPMcnLWz0OTNT4AZveVctkRQt9g3VG4B9a+zxf0s5kG5z2spHsh
h9vUdPgUSPIwJPY0n5uxCldek99yG+GoEl8uwY6HRjHJU8rFgg9ppWcrzJ+ssa3wGkUEb2OtFQXO
XLwmlTsH2ZC0AdkTuLek2gznmWmaAJf4mSF33s5iDu9imYiKVQx4zupyLFSqoUvLcjXvcG4D+RdC
cuUHLFQ6/IlK3bf+Z7upxEjJdpQ60AZ3+xW/O7XId6lTJVoE9tM876p3zPso1AAMvCx8E+ISrl14
zR9xB/KgZUhKQ+XJ1Cnx8E/M9s/0TbUN6IqDXJRuEfr3O8VkWoywRd2DxAsTRH4sAzeKy0e7SQ2f
tAUKRqJcAIhWZymDnlqwINax4bafrktd8clZFsa8y3Nm1AvKYr2YqbXmX0QvWc7f943VgLCW+8Wx
k6pOAGmEu1w14arOYIDR1iZzaqQJ7+AvDoUT+YlAIokpHZzhd//w12cwRTFBG10J2D0Ewd3KrZ56
05CpbAiTVeKgyVSIpo5MdvbUoS9BwTr5th86LH0xR8pS2WKHTv0tJ2CMYhIqtb5d/r0ECaXCN5l3
b6MuOFLeCEnQ/RnjiVImJyLuq6M+EUJzuZM5iczMgvbkbVuyH53Z3ZKmdLNsqOE33UiArPfGor+6
CA7/JMZkxVCSowZ2HGfKtSfCr9+9zRs4eQI0/Pms5gaYl6tRQGO6MH/UgN+I57jb6m5mO4Uald17
eTij0xuttcpKgc1M0vBZuEptJUvT8h/ml8KX/JLZiTnPUEI+ddO6jGrqKpTCjDMdy64xVm+vVSKC
0C5koF1Mmn3COUXfUSJHq000HYGd4vi7F3SAhumJY6z/UMVSiPhI3UVZXC3KhBFa9Y011H3lisxX
uzttp0HJjiKovbrTKTRf+NVvPBueGIiAe/3gK5+Vibnod6+HB5mx7MONwaGkFzvCOxcB49aoCcSv
QGztDATI+hX7pIcXNBWjWHNFPPhaBLntrOFsSj+unbkv+ffvTm1KmoLuQDRDkBnfejNaSg6yROyD
NF8AL/dnp+IT9PhjQ8S2YKQKzgEAVTz2ebXeQZ/1tIzFYAyUfg4ZbPMoOdgaSQ4DVnB/AUaSyNHk
vLIxveRRgJTArI5LjKC63tZJbHrrTRQvg1l5WImRUoiQyW6uLJ9rI9oqrk9lFrvZCSBDUgTS5Pdw
iCUtXMFeG6r2WHa1xtlyFDNXZOF24rFsyN/Hy/7JC5ghsL6xj0Nt4bpOMLVTFOl1IQK2AP3X/tuz
ELkM9sDnA1XXISx2WNA1Ft7iPcSGAn0KuxyvJXssn1YqpPADOxBZXnSdPI05z0jzc721v2JQVvYj
ZG8SHVlH19NhQY9ZOz4z2o7SYh1nqHtvMTpxZJMUZLWjCYRsvu5GxjyKmdCA6W2QjBGGZUc8XZJg
NXC9XodMOYuKh1x48N7sjWJh23Dk1j/mp7aG4AC2qZrB0s6s20OIac7RzioT9oVu2xB+mnWnAgqe
5bmPndQSzRdb9UaQZmynY9yRCo4cTBpgK7OsuMLOUxoxA+sHL+0pH83piDTcrDLP0mbhqRT/dncM
iYdfzkRkaWAAzgpxNCv979rcwX53pypN7sJk4tB2/o/giPCiGt6w7c7Io1XkysBcOStSQCRTOW2q
mDUZnWUBmqFm39dTgScMLAwdDgyNQ/OflUuOlUOHoX1pfnGRNUmoywIWJpz2uRni3r2gRTlADXkU
orDGW+ZKTTD6YSnkH7zGdCYIGxojC+eiPZtSxOx956pR5pNoArm/9n0N8KoTDOLdRHyfFt+I6DKW
8D27SOO56uWa8sCdG425Ztvvmx32sG+jU1JMNZeXniz4NTqHFcHvdDFpG3dKHtw+1rUB1N5wP4s9
Ohzm5rykpNpKqi81lt4BXJefM/pGEPT95HIlrwOE9ORo0/xvHt9jAsBb2iOhRr7xGJJWKo5hfDE7
Euzml22rpEsxpFwcnUDCr3MF2eIOFY07b7YGXIlOelO/6Bj3nyF2y0wiWHiwz3BPBy/jNmA8vkb7
Xcdz0HR/P1ExAnM3Ljels79OvMqMvuiCG58q8i7vxuk4iy//mg95EtmJWsbQbQ8ZAbyN9S2ubQ6X
Hxpnl9B5YhQ5cMcPTi0d4rDn6iKG40rtcN3vUHGIDsK4D8PbKhUp9RGEqIDfjSZsDRXhzMswomsp
5sltaxpFYcIUZqs90HtsxQCJXHQra1Y7c5UolJSMpFs/jYoXNBAJ5u6NZrUHxzfgqtxiy03oE1bj
i2acQpQVPeSyuYC/qLB1a5P/taM0THvwWngbkq3t1nc9104ifm3YxnMYMxOHdRewC8qPFGINUJaD
SnTxYtN0gaSpquRtnWmdPTeqo141iF3rp+Z3AaM3hOSA/7ORe2JzEkQeBwnbf8WvX8LU/h3M/+UF
z8vaTUSqHkkc7G2ZQcw7lC4vTsn0o4EeSx3+Rtg1LmlTkxroUdB8nZB3jQrs+76mgD0iAMESSiKk
oXq8K5/IYu5NADxvYVg5AnWfJppURBrwmMOkXK7yGPaPT9djs6wqSGNqzm4ZrUlxGHt6D0aBr21a
/1fnhzMvca5EXwMryfrQC7lSAfYkDJlE2Hjf1JGEdOMWMkawvHJejbVa4rAreEYkpSAXDguC7x8R
rpTj0br/8HqdlFnEna7WjraJWtvdFacUaIPTMlsNizSXxIDZlhAz/5/II8cDx+jI5xk7rY9t1EkW
GS5Wb5DVQl7cxVkBcLYsYMIqFDjmT8OCp8/oPR5ZHjYznKTczRx9AQ+qqPZKeos2oxvaIkO7qW8O
nQIoK78CdVuXtv+ChDJ28JBTD2e9qIq42Wy/vy3h6ZJx4wG+NXWOAk9MG25shjtH4oJR0RE40qCa
xFH1oY6SntYndGm4MyYC2DPwLfe1jmAie9V5AmplDjLy82yaYEuy49O5ZNG/Sw/XBmn1WrvjusGc
0jPLqyc/SWpo9PwsDbJzNnzwIZXzpERfEumutmVkUwKAIg6ECOi0yk9f7H/BsgClZ0ygU+PV738D
L55fl3T7+ER88bFDKzLlpHyXyHqYWBx9tQF5+dWd22Vh/pnnNYBNoFUbcDS/lVtzy/nklisEv3jF
+keS2z3TCwYiSvhXFl4lX/+kQf5ALDLDP4Yrf83DzncWRT2Xl27wHEWWcTouSdrxO7pSbta9+9av
WJCBGq6uhZoxbi0BYKfMO5FA6RJwluqANG/fg8jBIWbelzaXKhT73slao7V/ZmSY+MoGsMNW8iQa
ShEcJleEimHxfMzgpvIm7C6CjXmTesfxFXK5QyKFjhwURmveDQnlfYdnJrEqcjZ/Ik9Mrg6AgVIc
raaZQzRFCGAd5uLF9ebNDeVV5kEEUNI3YitORQYsTxJyZL35qQRBy1gbu51t+cEdlFj8/UUWjOOb
WZCB3kpxd1FS7xWoNNcFyyl0pF7jMTSrH5JknAijDIhHeB2+hGh3Gr0+RPuj80kIE4MQ694VFixQ
vApO4puJGrUtRCkoxpK8hmvVcWxlJg3xKN/BAJCUkWt5nwv1kxe7tNdVKn8UYfxSzgatboTBwux/
GfxCvp1sjU8fLVYKRjss/I2SwbrIKbRglHjLhYfCvCjoUwesCYHh2o7m4hRbmRr5IkbHitx1Lxiv
QJYyqaDJumZDMEuxVqxaWNoP0XtBUnP9TVD1+LiEDVdBBfPzokcEkCXtWi0soJodrqG6pZgPcTqr
LGzrkYVSDwVrDk0fkl4nmfujBy0/Vu1LkPck429LQnRSyn3ie03BCJJfirMgo5ebaczObW85YZfN
mILKb7Vj7hBcVt7F51lqupGGvsb8OZMo9FuNaNdHIQnNqAchftVd/4IGeTXvMqwIzq89bqvSut7+
p2oUHO0fIClNrZMOdhkKjdm4eu9k73nOceu3ncpxl3X1l2r/gHqK72uVyrjMuyoos4nVZF4MqLV6
qPXS4Ml/28FSrdQFBCrSk17kxcu2N+9CPHgPrP5Wnep6foUU2furMex4O2anqJXGouo25zVSkTKt
fFdPeFntIW2IQx8DXCfSKxXNrQRRms569NVK1EtHPaWd8hlQQQZvDH7jtmiqdqNMMz0JW3GUq22m
X/6FP/oaAaRMYyFr2zFqCBnz+J7k8mvRMy70UCxEHPN4p1RtUVlKGGSh5L42Be5nDWGbXzJP4bhO
XJo5s11sc3qvY43T1XfeCcI4SchDAOtYe8hbZO1iJHE+Y67elWKVfQbF8E3+yXu3BKQOWCQsDQ+U
0hKWvi7wnajzj4xG2bbZm/7HQIuS1XVBdKfJSxaRpHKGMq4M3w3b2LHB29Qoo5OPvzvwr/A39tP3
xBEXtKNUlLydfmkb69ZtcNhOiT5bYjh4iBTIe4VUHnc8i5GlOoFnUbabQkAv2xiGgoJZblSdhaIk
oBgXXT+G4TRlWGEKv4dx3zKFVKx1q4MZmNqwprbxSccrpfmbpdeXdOglsf5mGss0dNaj8a0rikoN
iU3Wcx8jqAI+BO5KhMRtdYoLEa3zDm4KhtcLzKcyphy2dKGWR7BjxN8PsntxZ9TzAxI7OTnCN8SJ
fe3oAY/PUN2FGzAIpvng1g2MfMwbmpFJHw4hCac6Pj4NrYKhpHPclC6VXOMWtc6tkkxT5YRy0Aqb
Jxm/qwJmrBIUOWIo7jFdrlY14iVjXeKtFsMRZdXBan19qBn3ceKovl5qT5Ixp5ZZy9aUH2MacoPs
ft8iDYiUPqgojnKEHSMJ9/3B3xgjiG82CCIW+Rx4JIcgIFU8Tg70oEFctHSSBR9SZTe0ZwihkWAi
QCty8dWUO+Ep6B7hPAYCkgqMUjc8pq6bMNPZjJFJUmplz7+D4ygP+G5cEN1N6MAzNCgAFT7D8WxU
TP8AusXzdfj+DkXNLPMoi8p9AyLmkoO6XDC2tagX9/vopDFRr194SXgCU8TC+8R6CZ06Kd6+3RId
avhlhRZoG987zQV0OTN2/bZukG0LK+LKtOsWFk3obHn8FqClmPnmbQIIVanYjiwnwPvarZIg1DW/
E2KhQ+YscXDzoAddvHG0xHhq2zHhjGgZ67eufWgBbudrtWZoFoE6XWcDiwelxxESk5LnVOjj7miN
JJfWyAq7v+FlgEqWNdT5IKgYtXqxlczjXG6fyc7E7siNlMJ5tB9PLFVEDpp3m2wtYUJzzopSsOGj
twB09/mHsPQa0sLQodjKpRcCAd69TAZQQiK0yQxnYEajpNaqFsL0oQsJA0QawlqK8qrzNwaU0AYT
lDZ+Tvp4Ag7NPhzsCayc91cBKUKzu+lSuvKAzCvx7eeiSHt+l/pEzWnYoPCkysNaacA69frO96QK
DoGeNiRSW9bOEycHTr/XYJsP9wUhkTB5P8mAQPTwjNe8bq73qgYkqCdSmJloPZwPyoLChMdtl4yl
GoV52sLaOXCfSeyvqSgO1ayejkLtVCr1cvxeF3RSraaNh2Tq9dUr5UW0MlDDfh/HD8qzVsma0d+6
X7dF207EWlv/iy5zGKp7xlGePB+FZqCb5kjLodrUVc2NPxAkbA8q1ZYVx+NPpUUWTtfmt98ojS5j
2Ht+8TIcnQfCqHubjH0+kpaHfqGvWae39lEXuUfIOjKmNPz/hHsnNIrUSj3d59P2JUz6P26GBP2I
ZnWwSAfGbN+NlvvH8/UyeHQ+ov414c+jFRkTIQ8RZXm6P9XF5YaDCb3HsLYNEvzpc3XZHK3KXIEy
s6VRvxVLiOQHwksIEAPvFtBTxzx/zAplWaMiWr+PnZ/Sy/2aDdvqlDwW0V2oN2SuouhwUPS0Cjqs
V8O7Nx/rIiGlAjJv30mrMTMgkEW+7Hb/yetRxMB7llU+OJCf0yTVLL58uGR2IEyw8hYbK9hI+kwQ
ACl+Hm5jAQcsFo/ZU/jdVpvQCY4Sp8N4RoTInqPO2DdDlcbnDqE84vxPVBWIfGdEQw6qnvPHUx8q
Qi2UlG3voqSPqXLSXG4FVNMsZVyD2nzQIuWtjTlmNDCBjy/dNgWomvW6pIHsHgdo9O5Zvk7qXgze
8Rq5yfLcLV9Y0dbb0flKIZHO8Z2Bch04y4GBYE05TUfTPedfIm/FYLFBgRLpYkHQfipmaZpbhV0i
NcEGGIeuCYXtIrAZwJ0IkHTiGILYpEVTtR7/xkO8RHUsBJcz6sW5HjaiMNyJTs0mV7lhNjd4vsPl
o3dFBGII/tvClroRzZF5hhatknT3e2qrzJVd2uEqId6CcwnRmuezXbE2gTKxpNJV3b/rWw90jAS2
IOjYnt7WaN/rHp2CIfja0D/Kg3SvE4CWsB4UhkTkXPv2NNUomXnqZOB6UtxGzWe92WANKHwOYTkB
UGFC71TtYJsbYdsqTfKT7OJPtYF/HjHtT0WdDOmd6T5YDavFL/WgkHRZcBlPPMxZBY1RHUS9htce
1XZ3ZqkBwxpPQB8XNUMU9CRPiF1rM7scYLNK76V3xb7JjUg3CY/nZax4EJYp0rkm7cVnI7yhelnP
J7Rd8pMlPnWwnZp34zu+9vMZzbStDFcuPQWEn8TqmuRTtlobb90eyh2MqgO1Vx7uB9O9oqxYWocU
fPZoueer2QM7Ee9dZRu40/riPUsQ5Z0oeezw9UDtGuLOr20TcjVUgkxvTxLaGTBUGQ3eOxlyF/rj
UjWWqFfP2IYMy4jhs0IZsB6W7Hm1OMkJyNWcXZ1WmAftEL+T6ZS7kGFDUVidt4fQUZM+dbiV5/5e
/YD76bU5zVupaAl0j0VurbIC2PiZQ+lYZ1VnNt912gTo/LycpBCbAYuVXm/MHsGqj2lFexXL2pB2
VJ6BeO823J3ZaAbkbRvwLSdEn+QQwmZdlvRF5Z1KjoHx9JIvkLZKgxrYF/BnZK53D44oDkPtvHf5
7kifJ7CeO59ErkQVGTKInwa0Ytizpm3GfiYyRYywpabmELjhkf4bLFXykhXJ1mzBbYlyfOOsg+bf
Uq3iI5LbJ2zzuMdBJ8wj7S4K7tyyurNZ/Of6C1bi1DtRuwA72FviZZK43veO29NChwk0mUh4cVcF
6IQTH4/nsk2bndDcsl5GtKMyJLdwFZuKoPawxyM8Ej9bSLe5Movk+ELWKCzSkt5qqPQ5ta4tDcni
FucY4uQZ4g1Fa5jfAUg2zIz7NZvYf77CniB8wo4Fgmlma3CKbjeuDa+0JNuotCUzy5E++fAJqp8L
ErIKelMFuyVRECeE4ZcaKwnyu/skZ+tmWTOH1q5V3Vgfm2QgkHW6g1C26bteTfiCmpXGrw04e54F
JOJMKdaFeM0UuT3wlhD0gqFNjJaiXVMNp387oPDkmLd+yu8VG+lMNOhjCxIcrXoL/9bmnzQNiL4V
24dhuioZDP2fBlA2pmUvd76I/0D039KCLvnUZOMDTdn6iMNRyzG/Vz2ynCG63kyJcMhfteO9BEda
rw9IqBMQqW88j82SThGRIfmyCVevZM+NiA2iH1nIRZ0G0yrH428KDPnSLnbGMN8s3NlUjUJ4BEYu
8vkffCxAKHOjeard3oA0BE1Nzz0cHF0YwG3vm0yIDmefwHf1PgpgIwT5BkAUM9nFqddR8XkYa8Bo
O80thKslfOB4QOP89a/VyKGOJbUsvQ8EROUdksqdCYJuzjIYq0Xm4nDAbjH1VehsRVpNJqiSdHF+
sJNbK8Q/L7J+2efTglBvlDJJMjvd4bV6CifLHYgjLwWM4CSF9De8k9tGkYZfN/iVH7NjLcQeMMqx
xMoCpk7KM699YcCqjrRo+r2FsdfyuiUdwsnuFf3gstG8IRpTTBnAxlzBABVjCiNdREX1yDiEmlAr
Kysl+8uux+olPuIvHcCsLbYeac7e42fsk36iM/LN7t3Y0h3Kethl1F7PQ4Tl/L3wJoQodzOj4oML
zuNJAt6ZnTY0vqlXlXlGsjslkzUpJIYfRbqTjnkx/S61URxFWFeVwQSAHZ2CKSrNsZjNkj86159H
kg0AEvZfNC/gEDGFm0zeT3oKgh6GVrGM5mnU2eiOx33VV39+ReV9gG4DRLWVahetlAdvFRiUnmBz
fo3TXmlq/XTowscLNAGCTvEfOx59+OeS1OdWjz+kCs1X90DQ97Q94kFKHX/kJv10efLxNqh/hfu+
UQ+HPM7y6Ej9g+/V/qHIGA7aNIrG/oY9WhzOPGABVMwa2sFZ5HHnaNl43jPglodWhrHUO+ojW0Qj
TsHhvB037AqwTQkLqNOaTT+OM6otvGohURK3vz90tMuphZQS/VUe7j3ivjBIYNkzQI0fu+z1X0/g
VmD3Q+aMDtMVoAVh8Ds0qvQUYrg1/fGxhPzDdp1GbZuC5DWOpdNlAJnW08tURVtJYZB3xQ6thY8T
wOBZ/I3k+KHs0EvtCSLwxfpl4PRwInwEyXSlXMVWekWH+uSfMny8558jMrlAvXByc+QA4pc4Duwf
WH0zGP9nITJqaY5bw8q0WTYnxy42aCsKp0ri1vyvhVBSw2eGHbSRQZBXZwfmzSKlZ1iLw5Gh3f9+
/HVBIVnCUHyH4w8MyAVfFIy2U9DOi7xJcsqj66mdD7S+VV/ZOrneBVATt2GWgh8+AIrP0IvTdTrG
8fgOKzvoggA9REngOBy6zA3mDi/OyTzYil77j+sCRqeHdlkM3Icn70sJ4hkW/MkbybxOTau21h4P
wR7/KaorSFW4YZ5ZukugLrA4+ysgjkaLjpzQVHl9OTHQeZ2LPnQpqhTtg+QNxplxvhVn0PtzlC8+
1RhzLRHzl9i29SRQlfxtvCtVyHUPp6loGatgbQPn4bz1F8bbs1c5jYQ7H2/TTnpCXeYEUgWIOMJA
Z2GzqFgaJ88o2UQZFuj70QUF+ugCi5J1mmF2bmW8nAjPVBtvCia5nPC3nma8hGe1LPuzAPvrfIeW
SE/Gk/gZHGbZGtIBcseh/YzY6AH3nLXagVSKkWRjdCA+ls+v8CFinG3lzXbeDsoMgPujBY/JUSfT
xRvaoqvIP8UogtpeUxs3uqj1jy3hmLr/U0zm88Q+RHxVKmFbAVohfmpZ3ehK5U0KfPGpOv3jfW2K
Wfa1EK3U9DLKwAqw7PjQCKoO1AjCRT4TG9S4YEBKBnJK/oMe6Ddzg8j7GGVnGX2eqx3PBsuX9OVK
DsWHrBAO+dVmqoxZX6xQr+VBItvy9ydetKDZmmOzdSuT1tdJlu7MS/ENaNCzhA8LB2NezLnFSvff
Clhaz6EwxS3dsEvSOcA3mWBLDEJ5oZAKk/qzux6aYzNOGQyb7E/lLnmGA+/4go/ezJkQnPPO01s5
XVTRRzahBoeGinWYLjrsHMZtqvx+iFyAd9321cfNYseLBZFOzRHgBXcx0xhRs6W1DhMPtUj2NNWy
hYBJTStXuREQ7x8w0TkvLzXMNFZuHt1vo6nUH91iNLwe3KcjkCbWA0EoezjBZOXoIilBpg9Lt3CZ
bGkkl5G9choVWDwG/MEufV8nKVl+GHpDpg/DxFMAL2q110Iiq6R5wW4nRrMLtupNBrHzcKadF3I2
mnT36DjJoHe2MWQmxvpQ8XBDyMG0uQP8znJbPHYIy7soVFtHzbSjaDVip2z6wEJ9E0+KmhTh/cUJ
GP3GeLjLphxJirFq+7sb+It+w9KeuRD6iyJLzUVKLfbDtmOScU3OlznD2xRj4RcHcbtTorQrdLNS
dgH04bbbDPdVDcMg3gcwghFR5u8bdmgN/P+YdFUP7W6iB/5Mi35EIsGpvRTI+jBPaalaiDOI3HfJ
cEM+3MVYHMoHAo3rlxgyepBJoXjCAT8DCz65oQaE0Dllyx5SVV9dxOhFpZSJSSBQygPM6s/4oFta
p8+XTtvLQqAqQJ8y3m5WdBxeki081NGMKkjTZzix7NgJvpNHLtW7xfc1D8Qd2bW5IDjZSYmu0QM9
ru/cWmcp1Mz/bU9imsaFNGgc1vsKXxljGMcJ+QK+ySUuMqW1G28/yIdM+nQYiy4EWih/AeUezmJK
UjTljJWL0EPJQvnYDfX03A5NZvreQgeS73FIrfW+K+flCeAS9wKtiwLNXKvU4ZDmYY9AZ3Q7dst7
juHowyqZUN630hnl6yV7jI3RkX4P4SJpd4lm82dsIVYNKxw3upFeaYkdG3g64A+yTV+7+V72vLAP
Vwdqn1Ls8RFPf15zVFqYa0Zb4I7GBT+oycJktWnez0xqutriIx1ytqtvjbOMtvLafN4qBn13cgcm
C2fL+BDRceJGxJwj4t2K4zN42X9bWHsPjqKKn6qoYF5X3ONeCFztrNV/lUJD4h/DJK1WLZSzZH1D
T7SDq/pUSkQmaW89kL+AHvaIqGltlqkjHdGRmulzZIiKtBZ52QRI/9Vcz1a7kLy5ke417lHQEb0f
2XirX6MnBtq5GI2803X/gotNfIywARSPjgbyAzx8g62wIHjvFE0f1YUook+T+IhIUcyT85ZHgOqd
0UnDxrtqA4FWUI6Ul8jfKTh7F0LDnfjz1s4VhWevRIQ9SF4DKREYXV/dAD7XRxYdPdMzemmzQWpc
7RxSaL7Ay/wjAEeSO3GVYtDYr7tECmCHmcyI7EsD7R6EvYhbw7JwQ5b2YjSoqkcQqVvGMtDbItjd
zcWpbfrh5WDHEc5pYDmgG2MNEVFunV9t0CZl5f55aA3vyRaHmbNGy92BzoC2Bp6OyeYDEwDJP2IA
rQdM1KwzXtAaBTJEImU1fiaPjVgovnatbhhBhUF9WREFdkjfToXh+HkaMQgQK+zi5ZOu3o1NGEgv
4ZJVoUltTzaoqIqKpKBTDjs1FFF0IJsnoITsLdHRlQ1IY++QwKWzBES3oVKPKOeJVUdsbmukBv8r
wx9yV+ddi4q1EzYl6rqA2yI8ZuHJ2NhONMziXYDel830iLCa+c4KAgLFoZtWCh5gCvnf1Wz3r1tL
VyTNeBElB86UKEWp6iYIr6j1cxbWFsEO4gIR0dbbxTIgtTwYTM6TBnkmbON/jkT2lud+G+fcT62X
iwChkLsSTatG9MJ1LG4n2rL25VAbSw8WnN9NHR+5YazIMYfhWv2Z9ZZb0c47KNgHLa43X+p+j2tX
8WmHuFkirxCihrqPM02sCRya1KH5rpfRpbb/A9TXZsLYdkUovFQwwuyCJrBRGbOW4iimhvfBp5DQ
OTzZypmMudTW+TMyDiCuciDcmyX8PoA2h5jpqHVsOW9tiPdCn/iXNxHZDhjcFSMEBoCiZcXLDUJB
xB4c2sCn/5qg8/MLf4lnRXzhQdRi3lcnQn/fYJ3p9d5j16tnyK2vHwSFrDVMkKMkePb0ejHSeCio
lk9czb1UattSfzThr0hAYIa7uRlDuUtryK54MHA0i6j6sQarxxViqhhyVbZaviHPiHfZLzqWUZBa
p+C2q8IMJvCBFbYQrZSNu/CU/Qof8RRy6FsSVp+kbXuTeofY/e9Ibs3hUaVYwzKfrRaa1FYdmgNf
RoyzAupxYXpH/EHRxmjDrfzG7eLWqHvLl3IoclpW411caE3RA4SXF1JEJGryPEkEicouOimkZ9xr
jXQArazlStx3c044AxAREl1q8vr8EFJt7c6NVmycYcmsv5ZcCIGNHl8dte20zAWsB92PqruJuRr0
wNJe9wcu+smYuvXWdowwBX9ccr4fSCt6vvCl2dSA1u3605eTBHNupR/SXbkrmcdXDJao/JLCTO+N
BEW4h4SL7r5p0IhJUOmSjVVdbKZSWupLpEqj87onEhwUvqvixMtHk+p6khDaGAgt3wGoxTIwBe7C
pTFbG9jr4gz5Sx1O/w+BOWmJLmY/8o32ehXDSqaH89Vy+C3992Ktw08SbXiG5qsWGcRa943HATLh
8Z7DDuvR6FzEOWca6ghWpJ4bSvAYia1dXshZjFkTqCfXlEUEK/L3IevPDNjJN12OUJN/GgWQh7Js
tNoc5wX3g7UOaOWmKSbr9GoU5UHYCy1h9blo1duo7r8LZXFgU5+A70DebGWkBxMvV0nYviWOfoU3
pGqVOT95T3p7A6UkRwQW8Dk9JbK0nYUZqyeZ44p6cu9QBvOWKuenHg6KQeA1Pb8ywXZ5PfbKHrGA
8CxAy8Olh6yu1lJb4VWhPr/qGj0viWt17IS8Sjo3BgaFTMvWMzMHp5mwQuzd5xoWvMT2n7D726un
VnuUmmz5hUmyFUm5W4IhkaWX2S8EL4hwxThodMI0g61c7J5dVitG35BfrwD2R9LGoRfDZXrlInIv
+YV6zo0RVnB9/K9EQH6n7RKP20jzaAG6lAjKKi7IFVIgUmZA4xscC3WztJLlMF1H5DFVaF7nJfoX
+OrH3kY32dPQkaMpSiNlfQdSM/ByLcA8JWYm9QfPvk4gLxMCckqx0QgFPTjKm/gstg85JFRunzVF
Xio4Laok8mGl52vybfw0x38Gn3sNMe6VpJurcPEeSqN3CXTcBYcmsHFRQCo5n+T1nB37DaEbwJBD
/teSnXO8D1i356yjV0yYLWrtmCX0XR3zM8SCenqD9bcRka7R025UhHouIecFzuoZhcgfPrB/yPnT
WFtciZZP3SaKg0bYs66st3uv9WndV298WfSOLSQTLmhiG6dzdJatKtrWKnmrryzUN+erAT7A1OX2
utYY8qFzo/0zRBadz8yG+biJWVvJW7H/+opBH+kavevKHwPyo0rP+3OSR6iaLZCv9s1AJiWgLULf
lAbrfnAVLM0rppPRrJrdqlZ/vyleES5xR0+aeWBetOIdOietKUdQJ56wwceOtyOchSjzqSrWhKIR
jKTQNVpIABQMoKj0UEMDOwoGE8iGn+To1Eosc/JzTsd9+U1+qXhjbI8Ms5BurJXyJtBLtC4dx3jb
2mznKZeT1FGjLTI+MAxEzJY96v9sfIwBAX3Blh2FwwVAyJjyqsHwqPpKCOVetHrfifoRM+0XMH4Y
P61zBCCRhnIbVSezn2qHLjrr+bh7jVaPKzPqTw4kINZWNEEGJOc55EKE6AFslbhu9V2jyX0uquV/
/Z7sDLYhmF7UCrtG+vJe92VlsmkVBUld1w8SDXvrJ+iWk8u8+HHNqtSOvpBjABPmRB+LXNdMEBgV
K1NcLHuxA/ozQWe3nrSig3UAB+qfX/7khutYDSbnFta0zBQHggjlSZAif4yqcSqpohDHoq7l9Wbr
R13ICL1GjlY1jyl8lP4RreF3intuYqSZZIjl+CFuBBn/ZoAI3wG80Qbydwm7+wWza+u405SaARA4
9zT8L9/4iNA1Xx8yoY+3jGS6O+yzunt/zYJPix3lC40txrOHIzKcewQk3YTkmPK/2bXbDBA/uJhE
47zCYhgEprQktBOViy05YRv3gStLPFb6lczJBO/O68uMU8iLiNXK9zBWNqzU1FnNaD5BhvZe4xUe
0Xbgvnb8nNFNYkNFE1sEXL926gZpn63F3kX0lF85DrByKEAsCUNYa1T4svPlnRtNytPjg5s0lar8
BhsR1N3mWKK4v5Bf11MfMra70vXi5DsD6h5Oo3lmsMx/CYs2LK9FO7UiTJzzRvHIEggs2YHDNSft
LWZ7F4bx8tsKybpLCCv+nwaAUN3/x5kzotYPjU5YKsGmzzi/A+XdiOVL9wFSoV5041LiyArqaZjG
U1iiEIyHs0b1IrdeSOyAwNSpHloZJGB9lHcSa68EXjeY2wpmJhx0wMy1X54X8ap0CGcpFzwzKOPc
YOzE9ynqijUo9B7yJ2d5P950NttpQq3zkkGkL4eLdqMIgwdApyNidl88TKA0tiPknUR53yu1ALp8
hdKzGJ0KFLWAGlmRWPYogGKD/ON2QrKLv3sW8b2F5SSzWz7G3Nqai08lEPaS4OG2jNZCR6HhhMCa
QHuIRa69v6Sq06BAC0RnLKVwf67JZtDfVUfWvZR7qDLig2uWCXL7vZE2SOiuJbsavS7UePKbwwKw
yzoHMyyT0dluXG5Q8R+DSFhUOiCz1sEnoXLsua3Yw4HI9zVSBEKAou1fQe1+sjRC1ew2BlIH8tIG
80IAHyX1Ajz+1Md5+PodbAJAE1w8LpJaDRpTFmWtn1toIJLYu0mLQUjGtR7cEqf7yUHyVnQYQJ0w
Epj495f84VVL1fERVbkQLhT/R9xdbfjJsZgu+KlAlPOjllHKPmOYD0hXkD0hJmN9say05MBz7f+z
8cfrCNflGsMtxiLbI2EEM0tHQc1xbcqT1Cg7xo8bxWX5ug8kg4VunGPuywcHTz64+TnbUzdS8d06
1RMz1UUzFrFKMfa6nTNA/hlwBtFfKUQwD9tSe3JUN8IZzNDsJI8CZ/pAdLv30zyFjic+IghRV+Wm
YyRu7mFPJQZI3bdbE3+DPvZcgABU7Yb2WCSymjHedtMPoegmgYEfXivW8ffGntXMV8vj/Z7Ua4nz
AhVQmwCZpcyeoog35NVF25x33hVGrNUOKURzT3h+PRh+FY/3A40XdQ9hJVrc0dP9SSJ1A2AtbSVT
HFq3iv0G7+gdce4x0qus4cpe6+rJ0NIiDcCMfmpKn9frS9XFlIQouG+DUDiTxtsyteeJESa6/ZwJ
esUy2JKGxceFLqLVsq2WPLVwJvWHosAsDVf6PeiTmgM3wnaRhA4hqFB8RWSp0bAoEsNYDBXBkSMg
xlQFjxhSCSzpgqz4D/7j9V0rdyUPq0f9x217TRNlTw1f3CGqSMHukdZAu/40uev/A+V4wdNMmsMi
tkAT9/I9HUKzXL7zA7aQmTUfuCT++1idppmAtK3mQMk54riS6ol8T9gRASiyzY1cyDP/QbdwgxUF
BXFUtkDPwywRp835Kcj2q69NeTV8NOVjLlJTIdwm5Cugn0kjegI24WQC3AzYVe9S7hc/CTZAjZvm
GCfNjT5x/6lNM/l9gQ0ZxnvOOjx9AxCAZ80ypYxDdC9kNou8j/MZ4JpZHQwu1qzleWOasfFp4YGt
fISWawwBj4IjINlSXuPQLrQTTC7ogjSO53xq8DVMk67vDEBqyoX8c7oKFFkdRMpznE7CBTkANAWb
/4N+QQVZS/QsOqCQ0KxaoCvhZRmoa9WtkrWisHBcoLdKzA3fMxIylw5p00m9qLEVRg+kzHe8v6ia
HiXbinGiu7nwKwQKOxq1ZV8ioMJUJidihRyC3qDd3+QZv3K9frkokAfMo8zn48MODcKUjUodJxft
dgPnzrvOKs5HKtASOX5Y8wwj+iL+f7u4pNMHbsnb9npaX3ax3ySBnSl3L4UkgbU9Nv0iL4xnvKjf
c8m8NXt5F71kwjYRtTZzWY2RDMK4WWDJfFXvWphQohKfRN5kYU7UQObsASVyoH+2Ugnr5GhnycrH
HIOtazrnRYdsZ+JQqm6bNQX/zhAtHvABoS3swzume6Sx8R6F2HvxSSDyHa6GR6iFpHWkCCzIsXwX
DvTqMpiJf02sOFQVCB2P/NmCKLy3cSxWn6I4enlF+9VtfcWqe5QOTIlkNUBCGJz45s2JGGdkCSp+
c9IqX9QB1X6OA1RUKOCr0PPg4AyGLJ8yh9oABzbN0cSO4y3aMGyaqWEWMy2KOBvom56cDoG2ElcU
/dUY3ZgLXZnPdMgLVKGmoFY8bm+R8F/fJsucsfM4TXZXw5ily/oknjN6r2OI7+MiABzr5DF+7F6J
Cgz5Tjlia8OhebPNgL/luWnvi/faUIvY9/1Lg5awL3ZomlnAqNpjbJidhg6LYtgccoleeEMMyOrx
cJbW0KvCnmBAGOqHiuIyP8pkW8QcHKbWEXhlK2zJx3zNqR5PnO0ypyehHdW3iikqqABPt++FGcvW
hiYdYf74XtaycGzMj9+CDa7QsOBc113PVxDtiu7J8FnlwfLJvoLrgsTIfAO/rbmhyTWbmu6/jLro
UR6sWPHNI8SbmhJmlLwxNGGIoC3NCzd6GvHnOK5gLyamuFRVboyh+uQbJvRZlh7asbijnNiLQy44
LMnocfWBdSKFHDMAfn/vOiF0oh1l9SwiVRFVtAPn5gmREIM7ZvFpJ1qVzao53+vE3S6V1xShU7Yw
P4y6YUEnOSuUFDY/EMC3wTYxe27G7pzEvtw4DgzB2y6vedBU3bvYNEAEI+MDYMSGzN5x+Y0eX0QC
m0kmrw0UZ9KgPVfBhq5gGCTbvUfulL63BxqTVYlirhSeqaqTw6xjP0qOmO6A9n6UY+jP/Q3XcTQC
7suL4diiGn5fjS/TMcNKOErNKeUnv+fxOUSVfxRnaj+RvsKMfUvkyhu0ZQG0d7RItMJf4F5lw2sS
zIe7qamlub2AOXmaGNdDeC6b9Da290ieImb4g8A1yFs0nX8lOYDw2GdXDIYh8GjeYBbTda564/cL
7CA44Q8GvFVtlxuw6qzkNiDiWlUGtkiMdBKdD0fYX9SzYcyJyrLGLnf7yvt5/s40YySLOx78h4dH
17GIJkvlHzmo1WTOVjyh7QdvJ4XLXDG2rlVqL1+Uh6qwNV/PlE4JH9d/cLbwaAM3ceDs/tosk8+2
/xFAhOvDJBKDaqZ8RrA4ZSQGvq8XIAKyRE5HgO6epcpdWwTS4xItt5JfPyYBz6DbNeTGNlWKFoCA
oBdIrVtdCFFopU3vMkcoby/sqzGVRKqO+XJVKlp7/oenQhQm6/kW5vzu/sdn3Srm8rHjW60d097N
Of0cqZ9n7ZIsrDUpzljcyMLaj5pcCJdFZlnEaqebVkLZ6ILn6u6IPG2JOgc3od8RXuSB4cAFdKb8
IE1J7fnjArn9Y4k+uXTmxS5jRE/XaeHrvU3ee5wJ0596FVMNRdZ2kRGb0JA4y+nvhni9uM4/5f5h
oehWuDOCTqTXvt0BWH2O7zwXDaiduBsCGwWWH7I45LTYDTXZsOR2OY0BU/rsaMba5W1JhSfk7SD6
ruJrl24PrU7vSnwdkTXCf/GtcdhkUI++0LA1PTsPyMwsYTa5k4iCuLlffvaiEoRohRt+CMjKbyzY
r+MkUyAeLM57tIB75gONoeONXzhyMKsUVE0ARviVdvVG9APE99DErBlrw7sChuw4f09cvQlCvAjA
XYMUxQkY2Kpws5OZ11c0Z88P8qmALFrpoTewg41U//Hn83SQhDh4OUAP4aU7K+k6nD53rRp/ni5Q
jpGIfUJd1IKxrUnUt/CyA4Qa/0vUNaB042VPZsz02rC4nx/4Wj8SBXSG2z9E7isYD5EbWpJwOA7E
/iRv1VlHMlvaePQ3aZguoVGH1AblmLMjwo87tvcWnTwQ0mrzITWK3DAZB/yD5jM/Is3D75bQmAU3
mJwgqJ4b4JVOptCsfHhsu2lSLYbio+1ZQXx4Ln4vBAnyJDpWngzNiEplO+6l+zhUWQvUMZRHLWQH
0EnZz0YMVd088k1qnyBHhXJplfrKQfZX8ievwA648xONVl5RRtRGIZDmLo19yBhEsVZg7BkMpf+U
/JSvgt8Zvg5sx3C7fCtDVkrJhsBYztDu3miSA9YZnp/LJ3s6kCaSkqX31RYBV7coYMNwIjPKEHsG
sE5PzywSs4ssItaEWTxARlwIoV7wKJYzgyj/3tG9h8JD5G3DT30K4ach47nRmtzWpGGNcFDlljbG
O+CzsjEO30JW024yCgB8rO5HHBMR3TyLGlfqtZpb2IzA9Qp1u2XH6oNUurw0JEVP9BukuJ1i8PxE
sEmgkeoCIgls6L01G7zfS++ixLzde91X17F7oG1P80DCiNsQuMShuFB/JUHmpwtkoSaVsA538qYX
OzhEY7DZX38yhTmEwuKjX5U4Nae2r28IHaPokkT8VKcpnTaJ3uZyYa8+wx679/EQD4Yr9DScIh+I
AHANB1I2x7vH9KF80KJer2nblVFy/OobGlFsw4owQ7KFC3JCL8zuff8ZSY0cA8wOiK+WTyqJh9+z
CqFElKk6MZZWfNFk+hSrDmzGiAirOK4AHyJV0jRvLvcphy0C8uBpidJrdM0peZS5kz0iB6WnY/zK
iWyR1HRFahpgSKZsuZh4hk5QKgLV4k8FacgPS8MD1+rmIYlbP8IZ//rTLGS7FIx/5/AZs/pihmWw
+JpW+plczAOsHSVG3yrQlynCfoyBInTnLXz1PoC/pSb9TNV1GqphaKcvTHHuvCUVVr+Zewkw2+bG
wnFUt8D+8jDIyFtpyB2bCP91KJDVDZSNSkirTdxTq59VozuOr7sv62Q9JsoSwSSiFBaz6YL/0fHe
kq5dSFxKNuHUSksTXs2SEvHIkkgIAn0LWbElwUWYyNHG0Kf9R155x5qjGqCIlTqGWIoMo2/7DIGE
Le4Jo9DPyhLRQwZU7Et3XXMDDsJytJo2Lx/WWWdu97YPESNBgUj9swUtHnQg6KTTqd1gMyBN6n/M
WP9lBPfhuDPgcEIz0DYUrja2B4PiXUqLMcRzWYYZUH4bn0D+6bbLDU7+RuNw23g4dU8kPaXDh/XY
uDi4pKOAxWXyUJvlW0vMQrny/HOaZ0Ao2GAylMWb8ZrmbC/+S5K3nayY7jYH38HY4qWXGTA8WCO8
L3jSLXpM15fMPl9//Kat8yyqi+4OwOX2CM6UHoDYrVopcRQ8U1jvQC1e8y6Zriac3vJb8dz1X8Be
HueAdz0YDOLVQ6bDfg+ThiKZ2KbXf2uGLT5uBIPOFw4sogMXJOiieIA1i1ySMr7D31BiVMhGdvS4
LeAS64wspVJV0DR+5Kh/n0zoaXBZgpI+TorU4JmXFqvas6/qFZTJRZt8CijVoMTWxT1pm4sEW2W0
SjXefZH1Re4Hnst5s774JReagJRT0qlPBbhaXRmzsdcSAwV6q9ew8jy4axR4/gukSFYOEy8n0I7e
ChfxjFwHics0cF6K+afu6bD5T2d/0uPEHGGWbXiDKTM0rks4CkJYB63LWA97Ho23Fmkw258jjO3c
hltXkrKtITl+ralbS8BcQGJaszU17D8zUGtHs6VHUSM8JfGsdUzgLfBg9+mh6TB3AitMkxjEqG9Q
bScyKAYOIOsPjedNdosGHTPiiUlSpTqsv0v7QaRUPdZtWryz1zZcNo9TCX2SO5JXLHN5ODMyLq4n
9YSPb52Q0MvtAD7jXX/pLJES1A9Fkh3tCFUvVqvwy1DlDHaCoJLLX0/z85LgtcOH4UhWU8GGbJEw
MFc3xHdepGn5l/tj6RKqWE8nOZtU5tnULMES40N7pA5wa6jFTUFCnq5kISqYY4cmdQLw0vgTBAOM
QrNzPp2Up2Eizs7h/bw4puCQ0ox/Lo3a0BIrXcM+q3pEv0C3JFiMbrnGHdm4JZA/ibM0GqOo7MjR
mY6f2MDY5d1kCj3RRSCmYl5F7JPPIAL5W1XS3DKfFbjYD1GKvVYsSTIIvIpdyrXpF8fVK93/dRKZ
TU8BnD8Tn/YHaXAsOMVUg+dAGR4vhFpMmWMN/pkd6PFppyoeW/JiI3yFEBEfZzpanrsq3BQKcDWZ
j1qdHT3bLti0v47TzOUBWIHaMiy3VdTW86nkNJ1xcQoz0nXSGzNI5l/F6lAm0mS6a1RHbngHpk0u
0ytjF/P8Vi5Xb1jYhLMkVSN9KJ/9rU12r+lFO6AO7enwXCZw9EizO8qFbUHEKpn1oFm+ZKapEx+s
QXVlcubXJlfEwj34ZU4/idvCUaSdhkHMCTmS5zN+Nm8H1MJAbA0UZyDLKWyAsG0Pl0URBwPurDAP
msqAQj73EIihYtSuH/qGaFZzCVgLKGY/w9Qd+JsRv+m6/+Oh8zjzA8mk+KTodczzez6JjLnBdBk7
TJZh+zz/ep0+exIsw1+3mjdRYXV/NGpQMJC6YhThVjnXGb08UuoN4aVCd/m5iHN3SA5+iySHa1lD
Nm3ahxfTXi20wfpw2p438f35oLzMGfKCt1zbUDz8ns8dDrtBY1WXQLTnWYBwUP16LvDrwVYHd5Pa
vS2YPSjKNZEGj0jGB6FXyxoP275ijAQ5gpZvL/owlfZ2XY7N/uRePV0l3Nkm6l+hyFearlpw/PCg
I9BSbgCUmXk/SlxPcEx1tc/VYd9NO6Sk0JTulAMrdAdRyATmSkIKazO7ldouf7CNjZ5ayAKDYNZ5
cm8xNlwG83K985iEf99H8E8CBEmaKkg4CHI44gVahy1xm2GUGwhi4HFQIQxo26URZGmwXzQsBYxm
3fWe8vkiGCCRl3VaILW9jO9Iq2HzI3nJXrMV12I5q8eMfGULPMmZEUVZ0eSvw25NBReBLNPc1pFt
ykeOOvu3PnWQ+jcM/QDyd5PrHB6x0BPRxMeWP9FHCaefy8NDATHlzFd9bJJssgyMzaQiD8NMd1Rj
gjSz5PYJzAwvnaXPd1GMK+tEd2mifn4mnbk9e5errF1r8Opiewda7s2TTSDX7iAFOq6QblfC/wVk
lcK3Xl6WM5PjoezpOezLyZFSeu92FHleBtO3fQkmKFJf3reEJnfiX7oL6tE2PAqOmA75O/M7ZkTn
L6s3jdKo/E2lmmxAgagtteroHeavUaAS+3kTJ2RE6+Cp10NLm/zPRxbp8qcixBzh0qW3YCfA6ocR
DaJuEvtyhduOYyE4sYfMOCFY0kF7sS9JFmsfXJW9atbpl6m5DB2+5F13tqT3jioGLypJ7vLsgaDO
9EFNMDxASMrnfLk4NETdMPpBFDZLN5BSM1KWz9XKGK3AAi0GsVzXGovq62CoFFjyMV11WOlOcNSY
hmsODeQzgGqQP5gwFM7+mUI2JvFFClvFSWItGHBSleb4pLjd/vxPr/ArBs7dTvXVxLN+scLlpnGG
+3TvHIC/kF36jJO96n96Te8+gp3nMw3IJkZHWztoS+n4Z9pFiewX9f2dOEndt/vicjM4g6+tABl1
wmcAlpwzc4MKumwjtkO38QMDKsLnhfUfgdJrxY9JlMo0fWa0Jdjt4y9u4n6qPswBSwUSXhZkFpOv
o7Ex0vNrip1aPf5nn6P2+F1POyhp/awRZoLZ1iiCFczjqlyZK3dFmHbAucEExgF3Jzwzo43MVGgK
vxFW34xensDAViBYY/N0fCP9L5oqLeA4xkkIGIrlI+6tFIwwQr3qd4m724psw6YS9D/WIr1JzqvN
nGqIdKs+XUDGdUHYE//hMrLDMbCfLf8xMfCfnW9mqd8L8mmab2EoxUWzRpbkJUBErfOb8Ixs6CcI
ipOqFV3ZclWv7JV6KJbq6+n80xLdESUa1ax/6lhC9ECxUo9vMC3/uE3WGhCB3mCM1g4nfSqMErtk
ZBC9emcgXOYRMk3oQvGpOHBkD3nkhbxGzM5cmlCgE0ZBsPAd0y3Qu3UjIl62xVkVP5N2C22CxJid
h1iKam9CsIMy/N2J2Zq50mwWBALyhfZXEGChyy0lV3dpNK28uO6n20Etkfqm0Zs2Hsx3zCqrfdUQ
eY+oZEYJWxGoXzFCVz0sROs4e8kJeSM4qlVvlpR7tquWFW4+m1HX3HyCV39Kpqzp0peqgW/YDk4Y
rch0/Kea7bFQm58YrmwH04Q+63jehBklx2DztUyQvx0loMSqPdKIHPv8eucf6Lfe25p+XqK0XFVE
emfYmLDIBnJkFNaVpfttpETwIKpJ5mCi3imRC3WqcEBh5yJG4c5nAk4i7HU718xCdkxeQAOP/bMq
THA/rVaTTsykCYo9dlfSXLloXViPqPzAhirdKR7UpATHjrw+w0i2FZspFKD/XGGVU62iHU+XN/w7
LsVEWIyCYejoeBMJDLY7o1/mo0v50L0GzpLkcHSGpL7KMiABY8uxRShrZ1ENlHJrcj0OEGZuOsF8
OabIMeKy3LIAKtBfbrwc1auwJkmf+NoyfR6+aOyAAxJaIMMIYOefr1OCEHYgCcq91RYgH+X29y5I
sO/RT/SYX5BlfAN6wLun/bYEov0esyn19V1onYnyWTFh06ergp4Rk7+oGOZRlwcTutjq+h8BXkt2
p4iC9m5Bbg2ypvPb6cUeDlbuxvo7TVIGKA4/qe66YTVWEyrcA9iI/1Uuu44jq/0ZJ1IqIWejFafe
xLRKZRak+FDEEgAZUsIj9TKU1Osk9/RLS/mJ4FhTnwZkI0DWU/3eDlZlfrpIzxEXj64/0SlRoDZy
joj8zhgBa1U9w0ew6/bjj1hRaUqrS5X5QX75DtbuxdoPqdaayeWnrTNj4hGU9Q6cCS6HZzKd2Xtp
/rSkY18ICSBRAGRjbB5yl4vQmX/QdBZ0+CualKiRUSvwOyrVIPIQKituKe+GkMdu0InXFjqAQo8v
E6GoJu0GaT5JViZ0m1Lh42ITlxA4zu4b9mt3Y31kuwAeMoVBkm8kQ0NPAqmoWjWWuB9fQZgj7NLZ
B8oILA9lIJwxf8SnF1+jLp8PxS/trS6HyU6vWxZn6+sCtVqnTTlJthQJoHCKsVNKgDxuVfrg6Q46
SJPX9vz546JXdDJBp6BqTkeJUlL33hfaKgh7+hKOY8ToEMljhU//iEbupiz41/gU6nMhCCT3pUtI
wTCr/LBc4tLkr7WlL1sN3Ibzq9nNE1FM4eSgIC9NnC73fvSEKj2FG3Jl88+xuYFzj3yannIOBRCA
LvoWiEFKVdI8IiNC4OJO1kpcr6mPDUwVaifUzpjfWWDgf+MzrfrVCHacfvD7p9jjMJi3S038AChN
M/aRp+pwqoVKeLFwolfPrZBGqZUpqVyWMokDx0Mit69dqb/PoOwGEgGWEzXZ3t+NToyWF891ua8n
onswe20GMO9LfX0MbA5grrRUB8LShVZ34BAi+SOvEIk1eBdVZFIGfo36l3GBO8ISOAgAeh/bmrDX
EQSxuoZk7cRpsbHwzdVV19oAFOoFP1w4k+dKjRKutPJ3gMbb8QGd1lp1wjGri3TeKB9pU3J/APbf
GS3BrlIAk2Oa3tLdpIOdypKOu3fvTo20UP4rhxxxaCRenkQJtQomjnR7BNW2kqI6VCjETj7TvPKU
N6EHvsvuk4axt4CQDojL5+QM5RK/XLpVbHR0+afHDeVzuV/thu7ZCykIzQVnobrw/Nyed3jMTKYQ
rdbfCp3yQfVB49pCN21igcF6z7lUV6f/bgChU0vg2dnv1dnUg8aidLVWD04dQbC04KMOsMV3hDQM
nhkd8Rl76cEzi/nm42iB17aZq0KD8h/dms7if16iNoY0huyZj0pK4REYiG9U4JRXdSqymSpOb7rl
yxA+usKUxqBE5TWvzuH2oe86gIGmI0c0YdQ3GBxsq29d8BFUsmdBtrzUsbXasB/ecUfnwdKSt1MG
PK3UlLKQnKiwIQZHaoPA1+/iSW5Ca1OJhMRrfQC0BaUyLSToksT5rxFwQn7bGieCaCjRZybp8I2S
ZxEeR4vzr9ruqWsVX7CTr5p+1E4CwGnlWd9UZIBLIq5yWEI/MwgA9YDYf1WoJsBPIutbsq9YCHAX
0rdg433qt3qTMcsBWOdTpsmDA/fniZ0cV1EJzgyRcWVZJylOnop9mXoMjmTjDiHSwBd/copCAHRI
KHctwUeY4K8x5zmfzpVT0Bi+NG7SVGSWZDUe6C2g9jePanLik5dU0m3o6/2IjrT1tfL3rnuaTGiD
MAvwuYwwW0NBxMhJuPckRMFMaTPx3M8TIupASJPZ1iHAocTVih9iLhE5QYumLnD+brUatGBp2rgi
2GvWwc+ZUd6fE5zRV7xVetNMl/MJVjqCAObLHaUR1wuiKbzcc1CoMpgdhUj37H2Yz2D8qyX0FOA4
BlBAIRq9Z4AXoSUdNdLVhhXnWJyitBB9c7eHUM/6oxAhofFCmuKCRYVuCNl2EkZphdqqMYk0BDPr
Ay4vrAD9/yxiK1a53lPMSGnrdK4XLrT6HkyZ2fJBTCBeeMUAm28/jAaTCFn4HT0kQXvWPXdaD1Zq
JRq5DCmkUb0Qm2l33SbVoVOS13ktsLnx0GHI+PN0I/ZzN5Vz9G8YTuBcqFFc5ORkYKXlB3HWJHDd
GLCvNltXrQuvM44artP5x0KWRyncIvIUTTZ3ViZuZDzz7cBzSuvpWvYhEbxGPJj3bXXL6oSJ9JWf
RJl1o8NEK9CM0Au5Iv6QCLASHE6ZZIRbaKSuFdswuEHe7IYnyMn54Hd6N+un7z6bdafCRjtR8kXb
dwAd39+KENGMfJqJ3y76w8Tg4T1hm/U8rREbN2/QPsIMTE8QZ8CwRw7UiiGX5VMJrJnKv6MMuXTQ
ny90qM15GhH+5K0nfJe83UymM/q/KV7f9bBkDGh+0ziQB8P0ekE1RKy6fatW0IY1Z1CuwmAF4RS7
NzG6gxdV4bOHiapwlofGuEhBgADtoCbQzj5G/i3BZpUVZ4TBAyFgLYI0GcT3ydWFcd08VMng5zt/
NPmT/8Sc13H32ZAC0VN+WqLyc+kBEryZuA9tE2EM9IoL/QvFzINwbWTcQnAOClA156+PHGV+Cec6
/ariaBv9snXK/s9ovHxYGDiBFBdoKsxa+9t05o+yyPvKfP123UpWXzS4As4cXH0sVzLNQUFssMkP
f0O9Z152Nm7b5/1pO+Acw3qNigI/RlrdWUq6pJaIOOxFhhNyF3wT3nW1prFMvZAdopW7T1GkVzjU
c22xZ9L52KbggtdxLbEa6AS2GHupKW8K8hbGah5znEe6kYMVT2aVOHLm1j81DdJ+TgO0fHzuNaPF
7VlObLhbXDZE3eeszAjahttdIU+VKEw9EYBPgAeYb3sSy+jIXji9owZTHGzPlOm299VAzZ8eKrwf
J1KC19bqBpjYyMpze4HU585XlMJOw+7p2PFJbdWSkVbyV4y3BTagz+gs0T7vfP9SBRow/QIptxtX
vVpJXJiofmHE1o6WeIMI2Olspukimw5npUU8XT2NC5zaZ3/KNZue0YhmEVwLGg3k4wXnLKIUzh++
jThtEu8bDwRGYD8Hf7LI64UX24fT+Y9Lyci2rEkkrw97Qo6IoRgGDrtscZmfcj9xC1KijKimBHFk
JWtCZK0jE7cFiLjKLF4H2x2/tJAGludqyL43YCAM6mUNtS9HBe71fp1OTyg3fqdwZni5cJ/Zwg2D
MwM41oFWvI8mw6mFdkNOoObM6e98l+tdHnZMlhXjMPquaaiu/Altp94bT338r3Oh3+RzBsnRMR/f
vd5TEjj/N/fHfFaFEULjhLR++2xcRLjN3CvAXPksCLHNWic573cphLKGOruVwKG3WQh/Ka74/aXT
9SdsFy0oqF5lk4NI/gV1atWsCOgsQ9iMKCmRqmrl1s6OmhPVolv8QgO+CeEFmbJCGx5gdFOtbCLS
NeurcUXizDrdnZrmw43gSWbpF6yqCeV0xaiDDchAIF9XL34BCU4NBXQuECMgdO5jkTG1uvhdjxek
cQ3jKO9jMa/ovvyV4H6YKoIdNj1xbxLuRkYK5XJdsvQwRUi8kiySGftHU2VS5EPf2b1+9lhYl2Oe
Pj1VNm5XGiQh7/qACwxjrn0UNIWxiIUih1R54Rn1GPOBRfJfeQ9/wSSbSTEhLXYeAGqO7NHiJUES
Onp2PEoejZ5jCrsz2cV7nGxhYo9aLD5m9md0AdIHL3SbJYMKmasdyFPTBPRsp1QjFkxIKq7YS2e0
kSKU1Nj5xVSO83jeXrlc0K8Pj3rM+uBekH4AhJlwMTijB4JBpaokhDWDCQyddPQyL19t56UbG4+Z
b7kXc2luMWWC3/Kzg/m3OTVh572qF8hH8MzwikxA2867Zwj+0CMbgT9a9w3HKeRe6GTb6PqNes6u
VTeqdnsYcwCS+UzARgwN4ehQsdUDk5pB+vIl9FhoEyNVrFbWYnPssnSbOpDw0hZNgv5ODyBEJlPI
azOlcwxeGA0HaKqyf7XiAb7MbAAM/0++w8LMFaVyeVIeLOiPySr+PqiwXgpd7VI/DdAyPcQ4pAG4
8e/jMi5FNl3FOqHCRsRuSMTv+aheQVqTIB4SfNhTktMvVqCs0aNYFIoKuMHpQqzGIyZu1sd1iwGC
sw4OSZ7GaoV+5iLBXH1gwPOTC8kYntMvfoenvNS8DladPfTex3EKGM/BWn7gfSV64d2wJcGyNyXW
HyYdZpev/48u68CHWusVyLUmwZXrJyaM5UhAZGPClHeHk3pPJbwjFSX7Llq1kx0Rn+prR82RBtjF
+/PjtKHdA+FPYU7wM8z9oZWWWlpdl4eadm+a95Ab5jHKYavcrvwZ+aCZFzm8c5eVJEaE7If5HFPG
0cVNBzvZvzqHTbmGed5RiAJFzdGdRhY8ATcpIMOfRbAOw3Z9ca5+UbuJaPUEOnYjDEMfm73Jcs0P
PMvEcu0Kg0l8OBa7vRyd6U6lVdvUASBFlz+xDjbmMRKWJILw3/cI3CTFwyrpOj0g6dfdiiIeuJ4H
HXHbMe/Q1EBzr32LzJ9pzwkFsZA1wtm+7Kc+6A8uDs5GE8L5D7PD7ECEuPzH5ZerUCSxgFo4kqK/
HIfdb/MSnedMuNLdKdVMCuZvw+lbmrVSWhdcrLEOkbfdPjfmB9Z8coBTodQktzmphATaOlEYYEVQ
1E6zfTWMWrTaq2UJ8IZaEmJJ6fV39Krc7Ly7G5RMoSdFVH+575nDtHLqUhofoA5vK099Ll09mf3H
qKjHqXgPqTatp/hu4JggMZkGQmhdVgDGDQdyA80LJ4djvgQogpLtoSTvvIfrnSBkefE49HAggsvD
G6/TIsKBxQL7UPVBtXOYyW0icPU3u8mVhNvNyYEO5nBqh8zxsAyjzwydiZeQgbVcvT3rx1ZRhBDQ
LW2b3JkCeLw7nzC1EHnmJ7WHRssl6PT944TOLK+9FftZo5dSJGVLlkf/Gy4x59xj/etFss5dfGLI
9G7MJtA+j9uqRgUuhZTyZN8AvLH2RmdDBIp+Znhm5rhtYrc9EHmLLhz3wpYgEl/57cUcMwfhT4y2
HJID5g/VY+fLyErF6wAbSeaMNuuh3a9sCDw5o8dxNqbyq6ruyr6ZVl9S11sJj6axcrfF1nxlKcAH
2K53CGLFalXRkB6JWODdyXvNV3MUQzN4LY5Al6lAd1tNLkg7mUe3WVFh/KU6hi6rnKYJwfM5NOnn
Zs2QIU+VT7mWlTe5hWhoe6OdXZnoQSMhYyUCk3MhaZryMdnccFkMXSoJYjxt/ee60KgeirJU1KR5
yH6VBytxICR4V+0MUVHS4SPZvHRBpo+Bxq6sFVjLjixuy9WltzQLMBhVavkXSbSjJofpOLAqj/Sf
xb2yvG4A3RpQ7/+WNdI7OT1nM5AXnTXTFTBmlJOf58ZT8iCrqM+ld93Hgas/743pCI5m6MynZF8k
5RRIZLcccYZY7hS+d2ycEp4m4mVixaHgy6WxGLEr5nrHHRGCr08Vxy//q4xIesroOoqkmqpilX+b
1HtPZY7mWi5obgm9IADned4ldtTBdLlA3T+3M8wzAfDzflUxcws3ttK10SXqmxnLQpjiYeUqqEmN
1nWoE+3gEkk0teMEqBr67l0HQO0TujPnuM7wVml1nvX5rjq/pccvR98qNfw0LtHOsL2vphggf7Hg
chKt/XLhVtXnDF818d/yXkFmK1ilCT/h6R5VT5D4u0bLOGc6uhFTpy03Ie2GjYUs0eFhmusAzxzK
kogX3EgX052ZNfcmMzvdajnnljjTned32G/N1qPC/UuuE186BEb0EcT5nr0lWWxUsnlc1MnDCSRz
wIkWez4rzSeGm9gHktGW9/Vzr6lZZ1mjXWZ50p3DpxU0f5hMhJC/2G37VVM1Sd1tNbHEYlKCF7om
/EoYfDUrlJdsr6OHCSAW3l082NN1L8pB/VUebWVOCOk2o3sihJ1L8b83RTsksVfsmdXI2kPaojKV
sZ7nKXPotEQW+GE04wy8QHvxAsbSwUvdfsyicY1A6DgBL/ra+Zc/de9kUU/33JlrraXwqfvFmh+P
+WUsyFmLcVN6bL3xlp082L128dieSrFShqfo/qSIVok7Cy/lfdVYIv/CJ23pw1LhnonD384Pr02B
4Ifqc/Cmcu5drF3/Ig2KHO/IOuIa3t2ZO4/V+F3YD9UlpQVMjBtPShwIMIx+i9TtcaJfXVhiCvEi
pLJG1djB26jAmBrN5qolUCF5EjX1f0Op3+hNDHEFKahWbicOejfdRcGNlLSStg/zYvsCiBl/WEm4
+0NHqU1FrusfPOPWt7pF5d5UidDI7CDXBOcyRM/gISL9kxU8mRdLMwsZ4CdmIre9Q2fRXDJ484yb
Nfj1r2HuXg8g4ewOVeuzMZLnZUD7HEswgTYIthiI1Uxt4CPplhEO0q3MP3JelR9tMxt18dXEbFWz
AhjgzkEITRoskWAJagPf51CK3P4TbRRxMHJTGZ6NR2HuGIu7da4goUyslYKLgGHNpV2T19Ar49Wr
KHDQ501qG6t9dqvqHYlQyDyT2aR+6lb86W/qBFYeFlAwR83SR4ouxGC7V1urTv6Gfh9CVEuD6XKO
byOI1Fw9HYLNk6f9O4EbIej5CwJQyiKEsGExD9ywkFTfB4M9oFx26Y9nEV25AS2NspWwYYLmYAfB
kLzQy7T7aDTYr0tcd7bmhaqWqK2kfk8zAX8vYD7kRNthWkHsdiXXj6ULK6HB89FipfUpPwLe1jwy
3TI+fuaCFGQKTkER2+XFsKOly9omoQa2q1YVXIdexb3wcePlJHZjdHeV7Atq0pHycLTSjJLIj/bc
OcCWCGVbE4vzB1PZ04tMl4FeZajwPp21iNGvQ1VA2NcRDRAKPkA6n2k5lw8qINyUAksczFJqYUoP
2Vfcss+2ZfETDZsR/q3Uyk2tN4URmDWA57rEQPyBs5yazGafHgvsS+LNgYg29Zpt+uvdh2Wbrjq3
Zgxnx300zzQsyxN+pCvvat1MlsJYBve4YPMB+aMEXYHPYMcUABX6Xk2K52hJ6kBCPtX9y/zuHByP
7h4CLzK83Y8WRxa1qB1d2xlVFHDjAPUZi9c3JbI6hBUXAyA9hIDewvk3xPOhWVZ6C7t609pLZslc
xRaEC+jYlmQhDA36fKC3fGwsWzbxskMtaNIa6m5xPVpP4QPTScHPBV/M4CErktmt1RRZ6m/7iMiT
koZyOhdHuoFZjI4joKUX9uy3zvQlAHhN4UbKGC+Mh/lv4rtgiB636J5TtI/dAo43T0LCeqGDTDAO
5K7++dsB5DbzXoKNLP2KMpBvyDlLNwI99rjNR6bdH8nhV0z87enE3E4MeyXQbR9pY+rb1yydxCAR
jlMOz6qU/XuFqItcbC1ZY27uuvt0YWa6SNgp0g4aXOd/J8MjpCG2jSBzg/MHkP8JdEY4gMt7OEgh
+JFwzq8rwC64n/HQ4TvP6URUDqQS/MvIgUVSOMHrym5GfONgfz49dGE76KmqibNy/PK/eZFFH3Kg
qKhsHkZdw3YJQBdaMHa3U/Sh6brpkTSf7GHK6BxY+dQvAyVE8qTqOEH/oXz1dY3A41Q19MqlnhVe
yuNSpLtZ1pXMCK8SGLTLKiRyL9QRiRSlvGyxn0KWwZcTqiZI5V4QdkJIauwu/+UioDyFh2LlNel1
ohrhX2mfUUnMw6KJPztPCEbrp3rxBomkAwrhfGIPrlE6pEJuFsDozzIpnYkdQMz2Mh0Vr7pa8IBG
TJSLQOACwc8N5HzQ0gyfTPpfcr4PWfBQg2Hl1BpZSpEfxKXLedXn5AVBjriKkc4rKGKkadxjMdQU
wZ8kSPFOWjmSh1GFWhF7Otv3q8ynzxiPiVK52v/FNkH/d7NnvsbTCPT0NEg9/yoK5zMjGnGHf1EM
KvG9eKq8j0OozeRKhZdHYr1s+t2DkSaU2qcjAlVBv2IHPLqL9L3ffHjznklDSFAFwKY5Dzl+3a3V
3aVK6qhlsAvZBSojvyeztDTs0EGkLJmS5q7n9T5T5rUDWX2eqrd9pzly7o0sLYkdFlI+ABxzvbzq
LbYR9iZu3or6johsi39PXN/8Z9v3ZNEwBa7lPS8uefGP224Ci5Y0xg/GuUO+IcS87FJhHnHp5Tgt
MYXtUyhG1PM37ZrgGa609C9Bj4pdFGif8RTkJjZPtr7kxVQ/B9gCTGOU/wfbLFqS2VijmMREJgPB
vSdZ3ZElVgiHLQeHRF6KkkeYnR9md0MUT3SRNnT6jVDABYXEng1UYeXoxK1GpoB7nACLV1YOiNY8
2ytu2txFEunOcsiXtML5BYxFXa1PW+cIqZuhuPHGgLtOnRQ1lI+BTedoJLbG08L0anIIorvKK1Sk
6TEO3XRQym8BcgTA2Xdfoiey1DmLiyHPmAfO3R79jYmaeUpwTp37fR4MgUXg8NLtA2qthmWYmiXX
Ycz6Qv4eW9Q0MiRH1z+zPHPhsnAm4uG8YDitgKq2OF6XQxE9c0X8GgcYbhNe5NSZrhzc0dnIWGmG
dCTwvsI+NWMC807Bu/CbXS85SyP/fjuGQp9tPiq3OhEMcRhRz0xB0x+DTKSMo382mu6iETI3v+/H
YRCn5FkQN7zOlKm5Z0X9wtN5C7FFlEvSEMOa7KN3VakksXnBgL2Xe8n8faauCSeiqLdJCV+BmzSY
NLrA8A3rQkSVL//4LF+l41vkLMJZLv1W2ud71v327YBN9Vg0sx+mXQxNX6yLk2oEuMt4NImcRPfF
6WPkR4PPWxuMIPqBS2P2Wj/029VlF8husmP9jwhmxRvhnO1bAxN785lGrbDcooclE3HulWgBG29S
499xtN7sJfjNuTQGBv0IdK/vigelfxs2RtH7ZEa0/ouEfvDZXH0+3u6/SGrHaxlgX4Xx0xi+GFav
lDUUsPoxGvX8UrqynjmupgbnNhEKazRCOi6gO4zewoUVwaVFKZ/ChuKhkTTnKBwi3+AogzRIar8E
9EinhdYduzsYh+ijdyq8Nrs5bMYx4bAD42BNxJ3KmAm1550cxjGrZCd0XSe9qcwGRUQTwsW7zjSj
CVh3TZrTOTeX+m+XyBbKkQl5edUhJcYQez956IiU10UGxX5HY45FWz/ptuY0JXG6rl+ObTNA+xp6
czO5LC5px3QiRD9Pxi19ZnbO9VKrzAyEQ/nbiPew62VkslZYZMqLrJtwLmTMeyibiFVJ3iOxYYrw
WlEN5xuqBtF1pab7dvhAenbtDwT8VWhjS+BQGbrN8DKskjMXJrHrgzDQIXDsligecbYhk0cZ23OC
H95cotOlgidWqWxwj2sTCXPXYDIENwwDe16xTaIO4zImb194O7EKay2s9vvn3fhYo0hyiURmLg6r
VYvRsoFWV69e1anj7VhgpuDoIPUFtc1QD/XaNR/KO/YLL2k9myOoRwofyFqFlttpiGg4B3K1e0Mc
8AbwZSI8SzldCeMBJhkfbHpTGdPf2rVyfi4fA9yQK2E4iTQW4YuChLfdGrYiiqOZHuj1a0N8I0AJ
U+LhFGERWImHj1+hxkHphx0Szww7Ek7pnMOfOJRO3g17eyOsCrcLxdo8XxnsCVkzAdrXjp/qTOVq
XqaLlmGrfJVhsu+sb84dULmlwBYRBhz1C+8r0h6VxSote2fiBxtDrGFVjtMTed3Ck+jYigJgy7IL
TVzhiYzkLdAl3nWNB4KkmPkj6bQ0Uqe6SHsnjCu4NxEGFRHTFJmMFy5tHH9TrTfJcynWpseO3TM/
Fep1UB1IlOW18qwQVI5rm2O2sVurDYdxJdRVKI670An2jlNtekuksL1HSD87XLY8D5FaYHsUe1li
QEVOpKrTH1jftqJe490ytQv4n0dIR0XXEQRH3mZKH3lZvB3cnVoipAR5AVOyBi4s9JCWR2Cdh93A
F80MHwug53tNS+HOZ34+SxS8i9KWI8XHlA0ifZcKGmt8bcW5E8Iw29eHgvkYI/ip4UfrWgBWTbYB
wfzTS+sJq9sCDFjDrgeDtmrGfqf4sbqiN+5HNZZpu9rls9NK+P8Qn8afFK6ABrn5nKZ4LuTeNNx+
jeWlWjcswFGG0R64JqlqryBA6g872mD2CkFxRAFHHxvbyM4Ql53jGJf8X2tWXv7QcKL8S9EaHPy/
bqBGJzyKowF5+hZCTLuoatZmo+GN+TQMy4xOkoXkhWF1IQXdVq/2RRVpMptuK15Jqd2gKVFG0Gpu
JK+cNMMbvJ3K+QIxSFKU2WgMaVqyoNwsfEz/anwrQMVVRDa5Bgt1HGZeD/Vphg9C69aV0eKluGjF
1hLCHJ7WYVQOIjF64pT3jWAErU7lQQDV/WoHUWcfym8m+Iqes5Gad+Gpax36c2ePhL+31m7GiSCU
H/aNEHAwHpSL1i8CbPO+ThqOhFK3ts7CXepOfncoa2LUzdHVo+wEZ6lBAiCVQKpK2TmnX6iY2tSe
B3USFhyJRmbnxnZMQIxeCxQ8PTcQIOR6AEFoTynnRjmKuwS9pTGPSM+4S/5bLJ0oJHUn003EcERW
c20Ec9pfmVyCH2SvnE5ECRGV9UPOkClUu2cbqajHJWUL+kyFIySoqWXF+I2P4F8uocCdWKLwAtab
tBUdo1zY0RN5BoqA416t9y9eoiPn3os6g14pIQzZLso1yGNwlYOR4d87G9t9DCGQGJfCZwjznVss
NI4wpIkU/cBd8pdvV4yLkHENv5Jc2kkgUrD+fGDsNlkjHc0fNZdaAILt2AvBXqbpe0tkT1d+fUUT
gIVZfm9n7VrTZnYu+e61ZRV96iiUsWARKgoTaWnLerGXVXE/DigMZTJGUuPpXXqPq8vE92A/Li6H
K78GjMholIpybymqqjis0behCIkDpeLJXs3pV1oXHCBX1Jf68LxqGl72MVUE8G/9IDLXGIGKt8Th
LvDWzw6Y1m7rDL4GJqYED+TptT5NAdUjI9+Oq+BDP5FuOOOSipY2QCXqrw0M8cSDMQtVMxlP6zZl
U6Bo8BqtE6VR7upkx7EPiY6cmdd5Zg96ciomyAj5VjTaSWyhILJCd2RG4hQZ1yFhWrpyGVlanSE4
8x8vmZztHuRfmqplD3E6phrXc2dqUXa/Jf57ZhW2Hl3Ndkju7n8g7zVshCJbzBtOR5h9FItcX2Fz
aMMh68K7THfgrbyHKCZVWT2FkZ6JvOoW+/nCaQR+8g/cJUAfhVdR5Rz7Urb1lW8vfdhTMCnGGYOA
uZkgM/w9Vq/uTHTjDekHTtvOptO0VOc4l7lU6OikSYXiWtGlDPafCkqwrVvHm0MP8D6D4SScXqxT
s5eEELSqVHzecK3SsgqxZdJm4+aNhfuc3QmOtrr44dOQjZFUsqT7CqnMfgvt9GN6YPRxRAKNzXWH
LXXKbfMcHWMAtzJuPzuSFLuDW8wovj/GF2QrmEzwtxWN6W9reaKI+7tcqMYQ2jaPXyhk5jTu6gJd
dy0dDXE9FaRy1e1FoSvhxqtGdw1u7+8W4ugS+HYhG4+BiD1/R0u5Q8MgzLojMUS1kUd1fSgT2+L9
YUJbpssxakWdcvlve72h4Uykce1qhI/Ng/JlSEtGnmSg2xvGffLabzqje4R5mio2wuARnL9m/SQV
yDJfFGq7RUU5CszjmYa0cS+pohZ4GgZNJdC0juyQC02Zsjly3cH03wd+7x685vaVH69GKvV0KLpB
eznYT3rPbNRWPEfjI2utmCC1lgnJgL4ZKE0B6R941mKgHhRLfYqBlEcg3cAQgRspKgqX6gkeCZOG
2tIIjiRNkPyPstUep42R3qNhUnyf7l0EkAJ3DJhMgx3Dxl/YRyp55PYnfkE9TKtStZo0zu28qQGO
nIRDbl/yfYIozMy3wAoKEDNhCFeITIqQR3Ly+GunzHsxhj1SRNzbGWEsFWgp3SbAyrKLWUiuLzOh
gbMS7Z4PxCvaskm5RDA60F7bN85RLHWEjJa8FQ0qJWsWGk2IOYKmGSBSMKOcYIwZZpNDczksZyhW
Lf28UOxGIw6vdxSL3qRFgtcppQ4ZxLjAhd9Qbgw3k9CIQap+8Y/NxmL04fjGwraNtK8QfUR+tPIz
PcKZS514luU4lMA7aw9/8/QpPUjRogvNj8UlUo5pV2bggMbgvxw3wbU7/1cAvlc5z6KLCg2Ay5Y7
p98gh9/6mksgBVUYluqOjhtQWYtM42Q63AyY6842swVJzvmv9BDj3f6PP/ae7fZSq9q59POUbPpu
gd0pH1t8EmzFgF6NJb1EdwhF8X+2H4MSqoXIByZ7voVEfIHNm3LMIAz+PubM1zzKhqFjwAvH3SLn
01Gcu+qD9DuPkGMEXaoNkTIKdyG1fqNNPFUUAguKlfxZ6hWe4fz+ijiP92uVM745W+NpFZfaIIIm
f4bJDrjIT+1NNl1GnwIjBNRP+BqY2mEawTB6HGMSAyR1FZJnKy8mW+b0FIirEDQjUFk7nPwYNYR3
iOmGEOKTkHx7aspkXkA4TG2hjbtHMaN5m3hdXRZZzyMLCxjCYIKQTES4zYiAFC5HsXtKljAtuInU
VZbYq6joxn5ng9WBlnEhL4QO7/YKd2fWkx1oi1oXfG0hbB5BwNTHVxOSbRAJqM6r2f53QqckI9zz
yg7VvDEOCB7zPPfUxYPuH1zi53+VEsGe3WDleuPsN9lEHt0AUG/5R+YLqyX70JukcFxCOolWi2QZ
3iWGqRkWhnErD56Mwt8wYBE90gN+ebhxnwSzb1jyKVDLQCO2E/wE9SdgHMiuxgznVlbphhkrdoUQ
KP0rUDhhcz27Oo5PbuP6pBQA4f5XoOldR0K1uG3mHwZtu6AlZVKp0uAwy7Luhr8QZDuf9AJuvPi+
kBCAUHRgyJRHoA+lygg5oMZou/g1bL9YxY0JQP883O2y8OGQVGty3GrPa//Ql7tPTkdTxI7+9sU2
I3n65yGBABBuZzosNLP0xWKFhKHXt3UPUezFtLeSLzugXLvUxpHQz/r+9LXL1u/JARUQ3WQPnwyf
q1BJclnPVw3h/JOOOLgZd8c/JhPL+vOpGd5BdSuYecR5eQhccHTm3IJ3bU6aFqRqHvKJuatmsCst
sul9qGm/eTY48NWybdRhyl0GKGF9/xMDnquGXxsMK4/yOEKUtS9SXXbuzjqwnlc/0DmE+8WnylkD
fQjh4lTrk5YXvHEXi0yNrfFq9o/5E2jcLFJ4HJGwCXn5IAq1mLR6Ffe/rbpIJ5A6TBaAFa8twZc7
95swyVts9BmJucpkNcsTfjWiugK/2ul0HGpcC1oePmgeAdA7AlvUFIQHK6H+j3gGHr4Y2XS0uonA
DupemM7jiCO/VOWxmqL/+1IWzmQterazQIP3rJvRspvFAK5NaD17i4lt1nGnUMLubpai3RDw+3Gg
K8y+sMBJ3nk7EnzlPGwAILOeyBmat0HHWLLGQTYefbVMASj/FCJWOcrDP/1S6EK7TP2NLyU+ZmLy
r5k9C3qozO+IGJLx2HEjeyTonYH6tVEhBExwtFXN+WeZIrMnVmi1rM7Nr/4F5qPeLwfaqwmw77WB
wyPybjqqBlnJEestIrKrsQNITQ8cp70OU9Md1pTbXOmAY/rwdv+OYRZeLhS2fhjo1f/FL5Qu2ams
BJAFJzQ7lRp+IGlzCyoqu/A40EGk++Ps+AdP60anW7Cv9kwrrx7sGoDFrx56xfU8eJo2H38DDZbx
FTOoYS7eibnSrAzLbgiW+KOqfIVTb0XMcEJbLsvwvcPp4yU2D43XhsswOj8wNS/wgQRJbr310VXK
7fZZZL3qGZ9ABcvw1fMo48LEkhVNCI3meNwl+SPNACCNmj8W1XNUT/+tZar4eQR+2PzwByqCrPfY
5gZ+MsTNHpt2V1aFRdttPXzLVHOYd2ddPWpltkfvk6v7Al/XNkH7u2XGBGgzIgggGCQk3kTWb6V1
yGd/4Kqq2lVDkeMpn+I7uzYBOQ0daZVDnqXaNGIds6O8PKYXw7c96OrEIY46onqV1HKvRDx7lj66
Yhnm5WPEuMP7BU4RGLhyWwtqizMPQ5ggD26E6br5PdA0myI5Hv+yS6v2ArPj0+dn3X7OwsLBkspt
zbTdMDyp+kozDHk9cIALLqJkz36hrO1VvZwPKuYD6a0WD4HjPziU8rUUvN+NWQ+7Ma0IXFxJqr/2
XdDNWbxEEeUArD2ZQoTlLTAGT+icLN3gU4wWFvMqhzXCrJ25no7dDJdwo8vnygQ11JJ3ZOvaBrD5
Jjx4VS3VfjSYOebeaia0ILARTx0HaXtbsAEFqJK//f9yZV4o4Q7/50lSKc0hxXHMoc1aheTFeKHQ
ODCjf/1+srNNewTaIdvakmoQBinJNZBCniKtl7ebTd0MGvEZ8zbQcRuuTNHpkVG+O7W1F/EVHmg8
MhVYvHVjG/rtUnXsFUJgZujmj7u8YNkkESw3IU5Ku34r6KIJl6Bk2wdYFMKeCJWqIjKyFH6JOEZT
Catcd+xSXYfAGN506BAnNEFFaI3kO6s5aW3OhckRmcy1UYK/7fnQT3jk87bFyZrJ4/nsxZmOtAVv
0aOt2+EkBH8uGD8nD6Qr2oJUSUgQJKFIwdq2agSFYSJ2MmZ1TIYxJCw+8bLCCACFrbfsQxeBdmB/
f33JyJ46KxSOoEaNxN9qWiV90PaelBLn6zccbmpWaBEQX6Hn1v11g12C1JLYQw0Md/nkjh7BFwqW
3howlgtNWFjKYc43K29ZcayBLdeaOkb2Tmf75SEavETslzWXDsxpoLuYJJUPSfTsKmvFC41ssaWi
hnsU3Cs5dn2bqG+c9wg3b3pNR8LS3FHQ5Z0ROn1/1I5vyqebnKB/bybpDP5ckS92jDm7yXPbPKwE
HGOl2J++7b+gZk0Ur50qb1hm4ByodcTGU44CnVsob54wVyY3PLll8gLq+HuhF18f6e1B/OcWyTvu
Nsq4MeMrS9s+1lC2ozp5BySK8EBslTF6at61Zus1xIurwvS8xNwEPffpZ6nqKrRaBj0SSgL7LYss
8XibBR8Bi47YRIT71q2D40Z9P0FvQ67QfENk+rXSOswBDW+PLODBUMRKQrzH25mIO4aID2kCERwB
r6t/bsI9rwXGefmlNA1MV1BGNINRMe1XDVs/Rv81RYkUiMpSy705kgvpo9BF0Z0xy8XxnmG5Drk9
MLaO2uJYyJtBHP1867ZMg3VfZrR+akg7bnIbuybm0m+aRgFI2UDKhtKwWtxLQzTvtZdmowFewLKh
t9QTAzhUGsv8/cDQhiH+hmaeGwKCIaG899wRJgj8PH8zvdfRZ1w1eUPN9ZYECE6M8R+xiHPWhf/3
uAF31ybzZuabycztYTs1zQixDBYe26lOyRlahGWSQIJOK+PSPri8lqxGwrG7lzZ5W2VGY7WdEfje
KktNufoQUGpZ319NJQ4wAppaYm5bvS4Yw6diMmVWhoDr1t+5mPPDDv8g7ubsFxmR0Sp17UdUWiUt
ExD60SKJkwSQ6cn2O3lEscZcVb7rQ+ioYvvMszQTpcNLheoQV7IY5TPo6ed+UW/P7bLNbxZNJY4W
lnuD66WXQ317QFtBYtwrcKFFgBQ9+VhJIRz2ns/aEcEne2idvA2I/PcHohVuCPR1W3/YW9e0u8NK
dg/XXJuVEevnQxXPXw1Cpy4IT73yfOIR/esmgYjmkLQ5YoIv7MhxobYBKD4E87mzErHBDmcbVTWW
RYzUtlj+T+jjMSM9UW5yrqoVfeKXo3BfaW0nNYLCWo5DeUmogn1zXQ6o8t6sxgDzL6K7qQPhaeJO
fd5rPQruKtIaUW2zNCjmcq+DECW66xGnt1YurU+spqfojzxLB8tg58jF3R5Km3qxn+XvSy/dHnOT
B53IAvQxvyzZrgm8qWlIbNSKGloIRnWQyCOD/tI8lh23TuHhdr6WU7ZLc0jUS7dLs8/0tsqXNXHT
Ddyk9mOayTfri9/sK11mLxlFBHWb0VtjodHnHikKALZsZG6o084s583IiZvwoQGJmVdRuLbKngGt
GuOBt0vApcp7Gy+GW7F1KmK3jeZ66Ba5nH6ugK60h4rDbXHzQQ/oXjvL63pTH0B6OKQWWXDIBlm3
rvORAmVdokmMCT7TO9//HEVuL1xCWlCVlWGhgvihk4v+tU5xxeoIZMR1oWSbtzPk5ztQe/cHEGHt
S4h6i56T5yxM4QYKmct0lYug6ifS+OKZSsI+cDIi1bQ/eO2g3Y/0M25wHIxlLgAgQZjfzU5hO0Vl
QVwnL6gIQLriD5LMWwy7XyjewNxtApTumi1l4EQeSGgrqlvHNE0oZCqD4j+99yyjmBRznlr1AZDW
axEH9NYKIUKPfAJ8+w7jEh0YEFQ6t6udGwa8wudTccB22hg2tdpTDxpRaMJxjMCX6E+hZvCi8YbU
Ustmw/rUGCmnXFzabS03Mr03mwdJNT/ADb05SvcEIeB0Ea4qzzrtm2aj2BKY08idOKbsLEGpngT4
JNaZPT00vPymvBkUqGF57SvexgFi7W84uSTD8uDrGOfo+ryhhk6SCMg8SY1IH0PloCmHM+GyhF6u
tzcU31124TdqNymht93O8fc+BOh33eJKBa7Yz8Fem9KxjkpoTuGkEGja+TSlHfV3bXS1yKq6GgAR
JD871/ER17ChX6IWLSK6cMrk8/Vxcfc1NB8ivSXy/kheU4pMjwiinMLDA2hu8xNtSpfwR+ddOR4q
xLKc5suCNXxoLYuNfGtWikpOBLO593FpcdZglD0zhJ3dqPxYMK0tjb7k5FpQgRn3wEa69i0JjEq5
rViF1TcaH2bA0OWeEKIuW41MzDijsJt820zAVlBVHLCXqA/X2zBQu0pPG6oWh1QtwNzEkuoswhcR
6K+zWdxDzkAN0LknlK/0/0wfXF54fHsMdOPMHSKsWMAYF+rKfDauZRJ1d5cfTOT3IdRbIoHFg9jL
Q+U98aOnCILZjK9ed79WO3bTvIWyIrNYTK+hq+jDJ7E4Uv7QtVw432lnQSC5a6quO24TkTvZpY+y
1Ek4iZq9h+P0qY1WU/ZzixQ1tBof+o9216yJSDr/fjk+TGm/Sotis40BINYQpifRvrRUiv0cLGR/
TPCoaKvRXZvGEfdCaUBjO+XQ82ZO/+6qbbu0Eg2sy/jAeB/5EJ71FghyJeWzaTIYX7IAa6PMoWtz
U0uj+7wR+4fhOyiaxfdqmtOm+D2QCTAc7Zk6ZZ3pO72FJzXtW3lIlHkcaFpZWVPfyD4WlmI3YHGw
R9GOypAjb+Z3/ydvQOKFYUb92kXp7I+I3ekc+3kQ+JLw6UaQSLOEVLvcHqbL0uUuq4k8d2eype8f
S1YcGMlHi9ej95Z9CdMAB5ODLlZ4L6NdLhvIszzv63ik35LbwFNZguHVRmcy/TTrMoGntsqETmVJ
xPmZiKW0Ikx01dvbuNMrHat3+Qs7DngjM71KymksU9Ml4HU6XIkPi0sqII9GSXoJ7aLG7EkGN7xW
Hgr58uEZbL5zpjr6clBStxgSg5TFi68oNzXoGQtZVN51aYrT/mRco7735UMMa1HlH0NH/tkGzCGb
g3nHL4a4XrEItzMasCaYgQYkCH49m28bur1nlHZiWRoUqyPf7pOv9Ie2qr1sTWuu9L35FdqKtwlZ
pvY+5knytcah7PfnJmWrrUSn+UZ7hJD7QFOxo3YbwpXY+A3vtk7K/yECMfvlo4v2dQ0Z4UsJgeBo
XTfxIkHP77Hup4V8eKoXgyizrni8tTwo0Onm+w+IyVb0BWyZfgYnLLK6RcvutN7wci1UZ+gsL4JM
eW2CI+Wd2ZZr51MGyhl53FzcfspTsGKEc37OkeJ9I0qpzg9EbutANmFH7wH2DERPUWGK1D+H6ziL
sPKBR14ejIvjVY4Jvf+KfS36bguqOsewhfk+1MzpthIdvy0biJu46gQ2TNH0T+USOs7m6njiHwTm
cRXsF9SG059XE3PWj1eS3jGY4CgpNAWQ/xdSuL4iMtaPnJD2hbNC1fjUzxSihxYtJT9LxQtmIY/i
2AW1qyzBulLnAepdha0xw+Mf2PXQinS08AZdqPSUVkLRKIcp3msjxHImW25ZH/HmXjv7ow3QeLVn
w249iTwUFxcY5B/6buAQfyT1RPf8+7fNhYKzDPX84jTY7kUb0xoILUlgpDXeYAy6mT5V3bPF8yZq
anRkL0qIYY8DcpOnQk0gpRc6lhn0ZO31toZA74KS7lQ7TdtRoICOrloC6csRpg6Yb91vH/FjDoSQ
WBg9OhefPh+QoUlmk9DPMoikpAH8mlFfNJuXWsD/P/MNdlPhoHI7azM9uGajKK1yhoq757Ntl0NM
8X6pCpCK2nQdQ7Q4JeCGveAll+dyiRhUqgjc2HJm35q5k04bAsiCoPFhCqkzO9chDb8BRHeDl3Ye
JvMgAKFh+qeo/3DZ8uYMmpxf7QtYyeMRnXH1+KKQCb0yEesaR05wx6XUyxZ0w4PvKu9cvLfkdJVG
Rqc7XAbhmShjsV+KjRp5kN0AJ2X8pguMkhJlDxskXru0QGu1tm1xUW+vZ3s542mPAvdKvbBqZdwr
HZpoWkK4b9zzCdImrvsfiRm1EzXSjYZd6eH9E7LtT2IySt3QLGgj/s1/TniE8FtSwo7b1nIRx7+u
PBN5gHdOQJ0kiIOqT9jLqC1be90/HR11hYAPCf1ViPqmUaKRKEUj8RNsNOhiP8P4KVnf60mPc0ht
odYF32VjQMi7KjcH1m3ZzklY6ViqysgXXEw22CjmUpJYqyc9RzSq5ETpBl1o4LG5j7Es3h3NeXYT
M5DbWw27PG9knDT8BFeG351jaKeiK41lHdCYzhObZ3ag53RF6g9vup5Qv451LGxqDhzRuxlCM7uO
fqzUh9TC2eZrFYep8MBdai//TLsOHqMtbkrzK7NmJgw8QL+FcOnCOgIRGKItShDASZ3IekxXbZtk
+/ndT3K38uifq0jf4ROtjAsgsgVM7aPLC61oR1IZcXbWwWvBRG3ygQxLwmomgyMK6WpwFB/FPdvK
m5Ujw7OYEmjdAENxoyYiJVNRxKVWjkU1NTRifaICdZuimVWxHK57ORH+Wrrgx9E+7Ajl/abu7SBK
BjJXYOEO7pejgmm9J4ulBpEJ+R6I74gcCEFpCFkiJqSalYRU9+oOs+jCmyNdrRVkcd1Bskz/X91V
wEnqECEHJU67uwmX3STPjipdpd7QZ63UY6Q1r86U6wYyMU0puvSaSEy2ga3IyUOE7Ql9M7AqQNgD
nfjwPHyRgfsM8JzTn7pf18G8u/Ij2dVdRqqtzjTan6NP06YANIDq5vEuZkylkaLkXLCvU45OlJq4
bFAhDJU36fn5kbue7yqMfSdJuhjqaCIQ6YyyCUrH9JYNGNZLr8V/FPbJ371HY+Kt3BXLAu/yiUwi
4uKnk2RIokD/FL1MbHfATWh4q70vsVST32cH/MDWzEbV1bH//b4foijVb/2/6UvW/HtxLYGlvgFO
i4RDqHeRuziSrAYybXJ1o8+9aDexsCAAFoJciSwxH7cDpKc0q/IOuMXaUwYjY0bIvHPHCCP8efjR
RlucsGxLcz9XrIdWPCse0+i6ZrDLRhza16r+rxHIgRODNljmfTziz29lJafm1xaHJx3diKLQWuhO
8tCqJWQWEqczL68dAxK8oVH+EE1/Dklzk8qcLvzVQSmOc6VY2OKhS4CermnYzCD/1YJIbWuqJz8R
Dh/wjnDdND4vZb7fhBiMGGlFYxngqvZK+oi5rbCXaa6ltLGmhZNIb4UN+Eecqcf45/M2OE0qzw5f
bx/ZdMz4UlECKTFrKA12TX6iK3mI7G212e4Ml4RCdmyNHHaAlF+X9AFi4eE8QMuMqgQ7mPCDbBbf
UNGQQ3X1NosGbEKsvRIQLDFCfIuW4yRf+2nbjmw1Zvwl6CBeRAYOkrNGsjGWvMNfsyXjCztxwFVE
y5SKOzABJhC7mRnFfD6u4mkK47YqSJJP/e1ojlUtdjRDWU/LcZzpnt5LYnnCGa1qU8q9det24/kg
2rGNO564ff3V5nBJcNE+xQ4y1mVLPUZakMaV3+i5HTGzZ9+mj9WbGn4j2F4c1/5g7LBGZb93PZDa
QTOD0dwLr95yE2oIIvmGQyVnplT7CQ1FBDarV3X5iCfZ9dvzH7WwHg2pOHVdZeEd2quSjWKyRKdP
EzgWVVypELdMDqLuScFaAcfKu7/rV4lJJQ9ohRiCwcFZNn7Nz2JFmR/YuyAFwFNlv+pUp4EivK7H
sbPI3lh+o0HG0ZeNsc+DcaayGlqeZ4BP3IhONvsk6tmijTSrrdNcroiMk2EIogv4UNFzsDD8OrIW
G4EnGRjqfB1Ie+UCF4s5x1y+pI/D/y5munA6ab5JYbZCwr8areVQmrsv67JCHAd9EkKQTuG2tvMG
q1ehhCRcQcVTbjOB7HYCKi6vdNB9SUTfAooaoBxWlDPDH53mjSJ+Fa5EOn3KSk6opHChwz+GswuP
ESn7KtQx0Lk+piKL6un0BbZ81rWB/+OPnFx6YpJYts6hE+njya0YGOoolenYJepowSBOghWiDM3R
uUGvSKtNCsRN8P+3Ynil21AasTO07yLqCFHUuuWHjA6IvibVblxxaR0BTyQpsHYyyAqTXjnmc6hN
QXJ2RN4/R4exzAsVomTw22lGI7aChRlJ0kvTGK2GNWvHmbP2y50wga/eyaqJ2RDlW97iH/dXJhhu
Hv6Tnz/V6wbBgdMcPNmt5A0xUw/H5UEcmxqVM58Wf538c1AVyZMLjL3jj3jzKeR3GDfRYD2oDj+Z
k8gcUVCh1XO0C9R1rs5vMCRdMgNZhitCU5bMFE49Kh4ZfMaIqQACiRlJOt+Izzszx/8zHXva81Cy
MUv/8wqfnVJ6QTkJ2Vu5GiXJx18ZKUdyGC/AwHmTfbtQ0dOyBaooVx/dlmyPi63OsF5cgdtQ5PYD
tvpOPJJ/vbGVTp63qyJdhung5ETfnqxijKgEvBSVMBZfZC/kh9yHzg5/2TM2nhNBEO/lYtMT25j+
Heci1Jn4jwIquejykecZn3Mk2Mrc/XqYkJkcxUjj+EreRVu/nPghEuU/y1766de/NHNGus30lIF0
T5uLZy9C+aNdSE1PRoNFO87Tjb3vtVtDWOciIRgsd/o79RPyCmL8HsDWrRTOG4N+lKO93GPFTGVV
Z0l1YYdAYpr4Lam1zotaOg7Bbfy8ss89nxCIA7eif1NI61Gw9V673pU1JqtH80g/zrecY6nS2U+I
zgFgWI8wfVBHyG/dax4kWCtt4tdRCl7vmhXMUhBL/wt5Qw2oncl1zgm2XIXWXaJ7VAB7kdES1OBf
FcwChAMVMXqm4PX9iKa2oMSKnzaQ9CfLvLzOPAytqzgMhzYmmC+B4TQ05FXNo7y2XsJxiSA0OsuJ
kVOdUQWCdjZdKfkbQDHRKVvDFq/c3ErUIkmViz0lpmcj7HO4At1gRwPJ8HzYCekHOAd5QUpa/0iw
kwQ7Xxd4EO0cjI4x/fhO1HdcosuPL58TJGrfnuS/316XIiBNTUsrj1Ebyqc44FulxVeXC3ebo1Io
ik19YQs3bb4JZpB46qT3MMuaqFXohQrMOqGJ0RD0ILsEjgy/2HL37y/VdVXdmOTKqpnZBPAOZIxJ
23COALLzn5aHXoOgX06ztW9akvzaCzhMkYUXNiR9k/FMmnl1I/3DImwENCzrM0lP5s5fxD7hdvYW
2yTYj4qUNEDRDZfua8RZ9bAFkHvZ6j5xUppwtmRHpbW163EBvsSn3PTZep/jp1vGStsE/8NSELqb
fmBn4b5Udss8qp8Bf58leoyEtQx7P2K0Pdzu0PV2vdjU0dVqEexHeAkPSo4SN31OEKSiugBAtyUB
m4sHeEM41LnXLv5ztp3EqFglHuZyo2t6JCKkJszl3WT7Gbmh59f8OVrQQ8x1/eyvDHFEJ94agpvh
aBkMVmfYjNOPjCIZC+hG8w7+XQUngt3cGrombt5nzi41ubQ01xk6FpbAHYtMVY38LVOwqpa+CTQ8
wQe35RiY0OTF94cwdfFHhvB2ofUeBXndH/SrplKqtk+oNqlo4x70/wHVJEsPDmNAbFCR8FCSaOSE
LQjE9VDIthjut3z/sNmDtcQ6TCWAXrxPknEMfUObWPfR0STSQf2clxpO1oKLQbMjb0X6DXXdPULC
9hgl0+UPn77Ac/hwUmjrN7nJy0/NRxc2NDIaAQe7M2cTi325fOPguNtM/1ToagMQC85X/Onj8X91
OhZ0FyGxL0K0x10DofsHFLrqC7mfVMfWJV8oONTroJ7CoE1meCH/FtXnOzvzrTWJGf1WLHXCrnzU
iGEq8O0/2Vs3q4b7enLNHpjOC6Wkf16Sm4fybxLISUDN8BhA/JZC5Am2WXED4CH1sTCmGrXeQ8Vq
/U9u61Y024zjUab1STN9PyeZKRe24hswJ9YTT3Smm4gmNGBPguztXEcrxjRAQ0W9lkSrC42Z3Ozb
flvqqUFdu87J47TwS3Xd4gS1JU4y4ZY+JAlJbC6Jn6oPFpa23n4EFeG5MKsh4aVO1f8Wrz+MzgWm
kWda/WaGtxhSqU/DZBDFw/g1jUU7WpJOEiwHOjomZv/DVGji6El12dvkuMK2uHjEC0CbvVlH4Ha1
IWayAFCJVoyCuLGwOKMNRtgNvc15bAnDSjp4A+5aDljCtkNfh5jxklSoJ2SZIFlaR18TzkzUrmq5
eODQzsEODmbYCQGEzA+FYVB5iqeBFKMboSWVqRrNw/1hOlyCB8tQ+CC4Zrb+TlfcxkT/x6y3vDNx
0USflvK0ROgJet4u9oZqQa66ev7igEscBr993G9DKuCrCJ94MEAJzVEpvczKP3SePQ5ryPbUQjCo
zpmbCSZCY850WW1NEgpsJ9PXyC94nt2igGmMz7FXe2aFEdL5OIT52xY/1+zfMEHqdOmWfWdnYS/h
Hngd9Rlv3gUHm/kt18v/fH50WAqsxhaEK1IF1f/cGHXvsiB7XDKVP6CPK7PPwx5VNx9nvcJ/Xjmi
U+ap1QANUB4Bf6VBi5Zh+7vhHud1t2NL4VptaNFQ3CZ9Z1uftbhL7rOJGvFdM7Xtuo0A30Jtf4jA
xZBmyOuraGSK4OZXyY7p9pTO4iER9Sy4pS687Of3n65Yuhptt/mL3HmuDWhaMIpEYiUoKi+9tQ/g
OuoFpZkfvXUXLathR0fTTW5illVwjhV9ulYHIa4YVgKgZ0PGgrrofRX0ThhvhmKs9Qf2nciCGtht
49JmdAHRyp6lv/oHbWB9lB71dM/sm8TK16M9/EoAJDzWFflLc8OdR8rB4xJzzGGegeka4g6axIiE
U/rg6d+bD/XmqdhWunkUy5xSvgmDgn72QnJP2zHrMaRLm1daiIKrcZie1eT0ZtrxqOvesvowjVcw
sKdsLRtg9+3SEcyRNvs6M5VFHNkERxXG4lCSkT6WZV1HXYz1LKFGkxxMLYaPdHTWVRkxO7ZKiho3
4aA2SsGcVc9EW0vwqHDAqRsPtpUsRT/u59PCMPdDwbOu1bZdhcwAxueTnIl9IMebgmJ7QyPl0FxU
tGGfzrxN8zsoc+NaSdsIUu1Yn5T3Ochl/wL0vDGIaLGvZQTwCR0ppq0YPLavu/S8NUzAy0g3zqak
CKd5Fo39fi2+Ma75o9f9Zh82uhZJ461i8XhMTaFLjUn6AZnb+BVNSM8KrAmONd6I0ODG2kNLbx7U
sEw6bwvBB05dVrwBwyEpRk3bQwG19Y/FBLmkWe/dJzViqMry1IG7vFrT/DUYb93QxiEfe1GPB8Tu
OlpiwFXan07oeklVkB76WUsldSjzzwEqx1Z1o4G1PyNljR9bgndGXeeBZUy6ntTGNtyE/NTUwaaQ
MVzDo93wYetw6hRWVWMWc3NFHdnKrwdgBRB3WKsaqKAZAmD/RrOY80TKLeB2d8h5OFBUV87Z503p
d955coOU5gKWJS+PYOpEm74L5bC7ppwSn1p+38MCc/DhOdW7Kdtk4jRyNk33kB2rhMKOCcUwVk18
pyAj9VB1LtClgZPyIYddLDWTiIYQnjybnRSM2A4KdUvp0PSRMLAdSOKoRPreivzord7HEthEiI+a
6AeN5FmNZtQWZ/LrQ4Pk7S8DFXkmSrD5CBqUgtLoZXW3VWtWYc9ocHow+qboLXpRgd7nXEyMeWvG
Vy3PZUzFcKszwK6f+crg8KnvXuvalVFBfGbHhk+XXCI96CG6aSjHLzLwcCk0XB7wnB0c1XozLRr3
dgi8878h2FVEccAjGrQ3672mHj6HjCWLWcjeOL5gkzu+sIq6a2HWzFxVoPGDPOgS7yJIbCK0Gvo6
Fl7XVQ4e7wJl5DEu6IJc1kb0aC8eWAJx5iOkXxvkN81aYC3HmVqfIpRqtyDHV62rPGJXPtTaoKOw
voCPdOGpCdWYSgtcSqZN4ipzdZMb6DoKqAeBN/OpclyUfmjrDlvsmD2YKTREglIr8TMk0Oub4Gsu
TpJCaVCDhP/j9QbB76yaur0ST9zQpEu1n6F8VzKUCk5xlApaGAeGd+BqRyU3RM1hTL3lIzCV9txC
GwHJLHAD+YYH2Bu9WAv1p9PLXgo59uDMasZ6aFyLecWV/a4zuwQu2WQGg7GipUL7nqydonil0UJl
F7XVq2VPdqZe5dNoNvqGVxN1XxRpLbeJaU3fuzj7TwUaS7w6NL0cjIkwaAucaejC5NXLCqEoTHsW
GibioIX1idxZ0fOLsU1fPyItWCDOBeVKrGiVotJYEkreUC+NEFqIQfM71U/sJrcg0lPqQ1H7HSZx
9ZbWXQ7iO8ic6XcvmIYNZEXLBVeuwUxuzC8vL0zcLxx3f9ncgiL2INSKrzw4SMW/iWXnXqSTpnto
B6m43bSO5TkBQuWW2OlHcKlJvuVZ2FDMThQPkeg39dfFMrKjoXBBrqKMCCSDP7gZaUqFtFAabWVm
O6E7Y6xgzZPdOQ7buTVQV4oqK6I/RCdJNWi/9W11OMTjYEm99/6hXPyIFzpHfgwoqs0ZXyH1Falv
+5gGkky5RQHqxmMxjyXPtgb09mFC/4SuLlCK9DQkbnkNEDfwwpKy8DVenDAqQ9Q38e0yF0bcIPml
9dz7CVzI103/iHYCCYlPufYcgaDLaY/fzAcKUsNohR7qb5w9Q8MFvumJrAbTsXp+hb5/SBDL9f10
gTLfsxijUW6NV0iwxWM693oAwLgDFCz73481lqLfs9vftqLPKBMFZTM+1TQf0KkgXNV8+f3MwXCQ
yXvCzCeH9HXOqS3bNURK6PF0S1CIg33ql8s6EblAF//0BbbPwlFt8xTB3hqFFYlqp1aiw7sgZH64
Ru5sp50aQUeW7faZ4dr8azmbeYp3o6GVn6WtCCaE5uQcIiTibiSwCo9vTagJxMWBB5g/uG/7WTfe
2ctgYAvPyiJquOx+r+SbPSxxSePli7mDmodRM+++JTCEpqRHOoqgfnHS34Y3gmfZ8RdT5u7TI6Tw
+Zs3z0m7GXezjYt7sAmbDv3B+L+OPEYQt6hdGy8J3X0A5GqQ6RMSGMx/EGpD6mNBcTtPWd5b22fS
oEX9XDMYHCQKgRiYJP5HTPNUdfS4bYNT2XbMx6mkPC23ekJey0pV0O4Zv7zm6xDkYRMBocIy04OQ
1wp2uSR/0Ere7Vi2+gZ0jleLDMQlbJ8soVpV4rHPAVXDG+SM92PUmtdjX/4kFrwfqCWbISr2xPpe
bkUOA9Z9xx9n+SgaH+tm6g7/F6D8TSorGUcqixSoqydF0MHTd17cqQrMBdgkz0O3atEtpoLoVUHy
muNkYnCg9pwbKNCB657fegRQ0guxXe9Cii6zAb66Pb9UuAaJcvFBMvdmwjuSBLLtvc88paDJucom
l8T9AfiNl91XJtqGR097Rly83k3iYS/haYRe3oXj/Kp/a8UT/VX+BtyBSpabq/r/zn5P8GKjQ30k
FWGy3zzYmJTbEwESuWIXz11xnkx9vF1Py2LWmUEKptJxdcerLYwwKD1NVCZMU0nHp2DBFgvU/Kmq
18OMrfDViwbJrQtBtgOA4iShg+H1xXZXwmI21EIWeER8qROBo9VSer53P+3bd78qxTxuA44otswz
SPvUrKA6rVgXT0SZZ3YXuXxS305isFtfqiKPHzgM7xibKBYNgM/ruvN8cNT+EBfoffyh72B402h9
JfUm73L0JiHludyzz2VZqwtsRhrKPh1H5OsH5IY7H5MzDNPrCGl8oA+rRzHU0dth3+90WlVsuKrC
z6WT0MSdX0S28IpowxAhf/BoOWQa1ZDioizF9jU/qM9wgbfcAWw9pPNmDnJZDuRYCzkN/uOODIwi
cm/s3RnNkCVeY6x6w5wDlqv/qT0WFHI6n56OEV3jV4qaGxUIOhqz104Ara4srB7QXFg22BKrvsfx
rQgfbPbU9cJrB0GrzKaYQnq8GMrpLppveNsI8W0os6iSsxWsofb1nzwfjWpMJnNZo5npJtAi31UX
s5LhdPWwj8o2tlmf21g9boPvX41Oj1UMXp/LzOiLfmoH76FUn+unFdhAgpBt0+fkPcwdZfVrOnyO
JAcJ4Lu+vrGWd69JiT8YCmdNoJOjlMiS41zR6sjxbzzBpaoucX9k2td8zd/ppcYYihczeTPT8AkI
ABOHDp7SugOLdMSkDizViJlgIEcmNLWwrdSzdDQD5ul5XTUxfNt6QxOWC1JKLmN/eVrpC2MIOFqo
yDzOPyryIJYu3BhCq6Lloit31JVXCw4p++rj923p9fMLbcSIlbmR1fTOXmwkIpXZ9C/cuznFN+GL
5tzY2vghfnq9PFfn1KNQ4LlT8l2pW5u43RWa6mWKEuUkAYFJXeFg2sS4wfeDeNvRIRbjYyZjprIv
MQ4kcRYf/KZK4Oq3TA/tcrqwPUflMAObRRcvFk2Dx7yG+/EPCw7WQAq6jFIGnfEI/p5rOeU8cP2t
XrUqREbT4cepBNjOqHg7sCZd2UYoxTK75B7fMyE8qUYjbmsSR7II2EhB0bUUfSVRJdF+9cXftMIb
tUXFSsSwG9RX4REOP51btziEQ72XdC/JVTGAN1Qs1g/7+R9/fQoo4+dWlbThFKOlXhuWRTRIgZQv
tajTckYmSU7eRlHSdksok93WbrsoSpOSio3ntFyrfrY3Yzsvy/Q56UxQuWSEko0XRAs4aTcONW3u
6eEPhIcGpDj+/n2g2QYrJo1S0EHcRyhB8XxCqWEWf8ISs2oz+OvbK7LG/E+FanvZWRltfeuAU87B
vGEGg0z4JdDCROTIWC2bW4qBXxx7QqK5XGhnAluvOVnAR6enNSvAhDiyTaYtQF0BpxqYpluHH1Uw
lx1fogh3sXuyeWPACUylsdZ3nBMPiOUDm6cBC6Vb+zoK30i5l9w/pc4/Qjp6RUKzyHCGKzXqb0/o
PooBbtfOBLGDuGTD3Ge8AcyIwY0SQKUPIbqJIY8ri9TGGpB04nMChKwt/0AurXRb0GoNchh5DimZ
vBlM7TcC0c7Q/UvoiQnaavbPOqN8aSyQjNN+ALg4gRKPABYjIfTJ9rP5h6FoxCv/6gF8WvYZi31j
kdHsFclV1EPFjlEIgNjtBjqoXcfwARGEIpcbE+bJ9qOZ5V6CrS4N6b5SOHltlB8KCcu//Bn9UQIp
13Uj0XRjkVhqqm3bEF9QpIlWpc0rx5HFHHemxgBkHUl21QP8w7/0PkHMWiueD2XkMg22fkP84W8k
3VSk/S9B+NsjjPHIxo424o0RcrUWPCwBULC7hvFn+93EQanANfRwyvul52d3KAzN96qWi93i7YFH
FGPQgGVhNRq7x7invnWYnD/pOwBgozpc9LLt9F9y0wbIjx680sp4ALmqCDDZ3FW5Yt548Rwy9/C2
6wzEfucUXAbamGWEdEQUEp00Ob7wpfLnbmXsVXfTONKR7RqTM/yuWTSQhN9Z8Hi6OWvEnQLuGW6q
6P4qvhx4aKxqDQVFNLwIDxzng6kqav1E2bfII6YqChiCoudbXEVs3+SRtVOZ0yrvsFH8QCMUVuqo
2LrKefraEWVI1+BwW3B1j5Ks4bknl6oV5/XzuKvbq5uXLUH/WzGv0wQv1wJzJChwcZykUVM9X+g7
YQPMpxIXI7+/TyWtCDlQHxw1c0nDiZ5YPf4vkWTuHYVxXoDT9G6K5qKCwoB8zYoso2z+/b3a61aL
qFY0gsnNesSZReQChC7LQfxwZuQYbsb9QlWbygQN8Obn0VERQPX8J+x8WPXYiN+MeDWK5HiS4lCJ
RHWt237NitRFCQXbbyMzuezwZlvSHQGP/vQ+ENT9W8RwPhG2rNOWpb0+zZgnxbIusy26D5TVvV8S
UcofXZf6FLgANoj5HGOIJSYy98RkDUd6OuqJQK1Vs7F9YzgFL0J6mke44ufvYvqZOKDk9c6Vf6UX
2H3ukCW25fPcLHwv+44ssrVAoKPFp7za9bLcE0xPWYbvv8IuOt9zEer8Q3ut8Ugoox5sdpZ8HBKW
9+/LftQfYKJ1EAzkUS33N6xdMryLoWzlr2RhaHdl1vdVtkGs9K1Vjyo0EW6vmn4N6J2X+BOrF22W
EdvyNHf84mddRhbmWmI1K2coxzLR2s0Uy5XLObIoPWNLvt4Lw5k7hViCugNT1Tyy8pyU0VzFfSzv
LAOqKQZkwOQoyh2rKAp/Xkl/0XfwBOqFbntnEVJID6SANdjZGlMk7okY+E/TOkcdFlCnoQbW7Psq
j38lIYGYV0fq3XN+AnIc5TtVYXr+di3er3z4apobO/O5iyyeJhXpCuRUZ2eluX1ellmfSlAjcc6I
v/L27fr3vin34+nqy4mdF5KEer6xzAmBKon5mOUAx1GKVfrmzKaFOSJ7/Qrov+N6m1Qx64GXdH7I
WWOGksaGXbuhsUgcdQRoh9KugTXCAPktKKZQ8tC+vyaghpwW4b0GjH7d2f9Zvn4WjKHpi9gZI9+2
JskS+QwEvO9hulFzBtDnggjGc5shr/Im8xeCbONWntGkEHRjkoU7cFj/m/GydUlBrl8Xim7RbLtL
hsSYL+1QfVfDWaRzdvp8CgKM3nsuxE0wszmudTw0EyKFpvwYQ+3MBymn+AdWrHW6tUpD5ANAad24
v4uSW5sqDUcBL3RYrVDMfxfrG6LvRzj6UdXZm60KjGx+IwIZ91ihL0AiMMqZa0PNwyr0aTWQe2sk
NLDoP6ebe4JBMnYR6bL6u2DwOBvDBivOvaMMkTE+yPEqPGanNCv5ah9nRWCnJAW/h7GrIQUs9k3Z
hdTgo9+MMAOugjwBL5/VZsr+Zg48Bx0SPNFzm5QBAM8eNZoddQKDyozLVxaZb2SxiW9KnEl779NW
Crc+NZhtiAcr3cgjOPyQHuMLxv0Lsk6RL0uyYuUoUak1OllJPCeErjGqqBzDU93GU4sdJq/6Y0Ej
KAjGuTLBM+wVWtP1U3GvJQ51rVdksnIx08dXQg8m3P9ZeKQDPvIQd+DjkIKtvq5CCPJyCLSESBqj
u6OK/s5SO+x/btL10OO1Er1Bx/oIl7Nrypq5Fpq0SqrWEZN9j5gUjgNlzuswVjzVGzMpe+o14sVt
9+UBj4TnYm+afvLrmjV1RT6UVqn2KxkZk7ojgt4erIgponYSq3IHzYgZOhCtJihYIfIf0lDd6zyG
C5fwn3Cy3IV9FXCMgJIUCJxf1GmTX3yuCy57N7r6WP/zR3fM0wW3DZNGXmuuyiubfU6M6t0vzV48
dfociooexat+vzUnWM560w9olVaoSlKkx6zN+zU6oPZ5iNyEgGXyrMpEyCUBMMwwvcv0d0ZpEF6A
Yq0U1lZU3SdefMaGVZ7gO4e24jL4kJ7e6Gl6hl2dxPnOSGbh25RRsxasKCSOJRdLaASXNablZM5z
NH58fZedeP9VZ17h0SBnCFAMqSe50UK20kOvxROxM00RQIYDSTGDL0JncbpAsNjt9j3MOyy7lYJ1
1a5IlcwGQr62W6HmSXTupL/9ETpe8vVFIkddEazwNXKmb/nJIVcH8gatRl3cGX8YO1yURb5tpQho
RHMmO1vS21zRNeiLkfd1d276fvoS6MmgM7p67Yd22w3k16uNBCVzXzlvjgH2KzOP7WB6E4tt7kJW
Lfq26Gu4bM7RPhcpImCei8MahrkwZSTxao4uKwaKOM8GdYmV1EsCW8adrFnyC1t08PgfB2+zq5Rh
j8rFNhv5gdxq7G7fOBwJO0ck15Q5pIHMvK4HgI/7+gd14qRVeMpmtRZQpMg6kgzIJx5xxCWCh3+G
v0ZZ/xrIki0CcoBdDeh0hbTI8YipJphl/W59mgcvRkkPZAJCw0jlSlfvrjJmxPNs2NGh+q8Y5VBh
0lkeC7s7W1nFREQR2Z8CzCWx8CLnNVpsf9UW2Wy4tyDtsHmODBONiLVmALhq+IuG3wlW3zHD0TOz
AqfZfCGEjP2BxNHtN0soUro6RmhOTpGWysu2Und2IJmZkoRUHOMDxw7w55s02TJlYaViiB71VtGh
Z56A/Vmp1WbnZBB+0QIvEDtefF09pgbZ6JzY/x6m20TOGHgS6OptfD7VJLamKhj/cPSHJsV2JZd4
xa5Emuei7EzHjcaBV9KwqchV1ly13g8I0HLUf0vko8dFLAT5m3dWGv71ZbtbLN10EcZDup/sorGi
/q4MhhyAo2+FF0zzmNnK5D/0WP6Q6KCuYkzRI7Q5dh9Fw3XK9FBlJie7eNMIiKvCSxhdo9ZC3iLo
hG6LjVaPE3xiLQ1yxPySsaPIFa99gKGs+L7GhtPiub+lGV4WLhY9XmETZizCgSXpOpqjBX319/GX
En9oeK3xdU8NyE2R1noQYnwqyazYhYcJ3DfKamGNb5VVaZtDA//mUSnNgGPgyvLoCLu+r471JMRg
KVVCdbgbQfWIumm4Tp4Jna6wB+0jjqICE1pMOiycg2qt2K9iQaI6JSwsCDTG098xXAnNMnBJWtFc
6i09Lw8+c1cPFGw11KaOsypJVya9qSgPrPujxvNiFzpA5DumeIpVm0e0gE1/XDQtQnte4/kxokB9
X9ScR4VV4F9Jcx7IVSfeJ2ptaa3LS2Z6CsKTecB9/1iCCwskPF1woqC2ABgggOiCiYbvDgmzbTAl
Lv8fHa3bRxYE+29fjWiqy6DreEmPVRTVSUWcNVm3i/PQo2TLzzbL+u9RaBPHXKTWJN9xWXCOqCpD
Uz2qUkJrLj3K5yvax3nyIS+KxqosHbFItiNBW8hivOPgjvyn1vH0tbpLf3O731uccWiosrwxYZE9
SVe+XDFndtrblpVWaj1Q21G2PM9Spe0Act1PRbzsJdf/ksxr9qNQryu2Jo7lbz2A4Af4JxrD5BHJ
hQ8Sp/nX6d3+UZKEmb05GLBRir08IBwzs+3jkZZtJBv89v+heN+qonSI/eWWpL+FrtNK6tK7Wl/2
fG8Uvl76MKjSzBMLoCucblnlrnYjqf8kfRUtNfc657Xnd59w14Xb3rMlYbqDtYRqga2ek9Au2XC+
rxOoJRfl1NF5H7Iuzyz6Nr+7yctVPjy/tjUoFqCO4qhS8T0KpEHGBID2S3bSj3uEX6ZpAsPjcgH3
Nf96mRDgyM3PJ1jnmjLuOxzVWNZpqOF8dK6yTmn5tqnoA+d7MBLcEBXMVyvR9CrjRxY69JO+FBU0
/X1JhXztJcx3yfrclRLBFAg3xD3b+djUx9+UNAhi1kHVn8yA9F0VwbjK/bWw3qWIKBCkbpFjflRC
1oTzaIRZnfQfWEOw5E/2gSnUdDpKvNWJVE+99M0uq+X9EhekoP18/orJmffiC1ThSInXw2YzvnvG
SSrRCwNVYWfNYgTa0uT/RvqCgMJ/k4pn/esTVL+rSEaWWDsnIJB+Sxkec0k7HETLcGi1qs/E66SO
9IcqcqlXGjH2ep/yKUuZ/3fVH9lTFQw75wLZ7PcKJNoeNTEjJNNUfyu3lgQarsG2l7YsJmINM4Ik
ZeLezXqWyZQ7ci01DFvWjKPEaAAvqkO7mEGJPc/X+qFD3lXl0QpcwqAHyoFlTH652QNoay8+Xl7C
obGWM3/P3Xuds5k+/nby7I+I9tgrR3N4sP4gFfF9wZjJOyEF2OW0MIEACfSY0rYUAu+ye6snr0U8
z0/4yc0ida7G7srUuFEvW8Q6VMtaL1V6dPNSZ8kcwlpJ1LajOD68NnwLXGk0U/OP4C1AKJJpVyUb
F4yUg5ga626q27jwpXbM+l2TKTQ9421OBRQ4K86OJ4toonaVsPDad/ddcba32dIHPyvpokNroNyu
IdS3Tsj13K/+irqow9cglgaD8GHaNlU7xI4mjrREPckV3gko1cDSxx+NBPwrAavO6KzlU0JnKn3+
3v3ZSSasF6XUVoAFH4GBiGa/MuTlHvdEm/jBbUS9NlFCjtduA5cVpK7sz65rYx6nY5DQvLreLPh2
C61GKsolQ7V1q29OfUvTr5ZilZpM2hv2j0RthHFOH+XM5zw9nuSX4wablDmOerJRpUX4yAbA8Sib
aeFyTgcqF7HznxwSRaOAUvqBa2rCHXDFV6N77CcK28cqfpy9PcqJRId26jIOiTP2mFFonmAQBYY0
9//s/e1s2l/eNZceBO+ihktmDHo8wSYN64NnwQZSNH5dDoOmzGMe+o1rcTST3BJR/A7jwMIvo0yl
cVi5bsS6jf7QLDjKgJNdFn6YVherYlVIBa2IFR6zX8Et0/ksZBLbqS7bfKz7YQyG0UZSFIFCZYbu
vur7fgw6mPEeoQb/yIl/nh08M0EM6rTJpfj1tOFdlSE1JHwsi4Fjkx3AwQPC0ym/LmHPi6/TzxAB
0ctYPv0LIGfele2Rue5ginH/t1IEQk9jRqGY6qyR4UmG1Ov6Co9kYATSFpIuCuvAEWPLmWwqg6ZY
tSAyQmEDitVR2ONXdxO0xgkjltBLoDNT6yqhrB9tkvR5esxXPufhDgSyieIwjfbVSFmzTZdSJLuL
U+3Cj6ZGnnsHUmg1/7xvv3FlakbIM0kzkyO+DHy+r9AqgOU84PuzhSBPmMCovvXSxVJRIsJ3ohEG
104tW94xd2vE+9atobM1+U/SE+gUX8uYXyk65YXLHagMDgHnysfna2Lx9lQdQYIOlNuQDnHTMwEO
KhElEYzzoHwzGcaV6MxjIzktTaugs50mNpbutw13HgVU/ajt6qrHKTXgkzcZ9wxHpDYPucfwbbtU
hWiUMw8Xnv15oxDBktYXlS1G9ND9wdvhBFIZL7shNpmzKqzsYhcZ+Os7slUEVnclKXGnyoA2DAgh
9O2pGKrytzEZMjqYuScKeT5gLcZG+vR3IdFmGaFmanN3pemsRPvNyIwpMKNsVaHrbrO/DOMsYf+V
hLvpzTUzlN20IpMyYdA2lc0Cg+FLwECOtfUMCpOcO+ZLhZ3+WUDn+IQ7uV/yeMnzWev2ZIY8lf27
7ij7nTygSV1KTqjILC/hIOzdrJel0gYOOWzM73QoWt/qImEl7aGr1uBd5uVv6UljfcOrbe8KIX8A
B302id4jWcAFQ8i+6agbzmRLH2ge5fBi8RZDSXlJeYE7TvOzUS1cws2PsP+kwML9QXhy28Av0UpJ
A3LUJ22hDQ0sUG0PTjeq7fLFrNZdBm5knS13KI4cryPox1l0jdbz9ToHcTzAI3Nvf4Bgq7wTFMtR
1O5NIRoscuj3IPkRMdv3RHEg3uZi4FXes/PQMZv5ReY1E555GKYrsDiJVh8n4/dOfDuSIG8LYgKt
WYO+Beu1fx2CekjIiFXZ6dCD2JcE3atdboB+eS6d5X0/HSD9DY2ceGQPjT4hr5vyCWbIWSUptiZf
ePShoT/xcVn3GYCeIwQqYsyBtmwYmb0EuSLuIRgCoTVjn+dWhjtQWJqxo3EkUkwG9izcwcS9h9MW
g/yhs6jzWThmcfUCr59ZM0a2uZxlEkPZLuX34NKdGnoJi7AAs6RUr24I7yW/Pm8wusTuvUmGkcTJ
PehbfbK4lUYWwx/vjxMfdlijeCLUCt2gApHNa1VmbZMJyN1AJcNlevxIcb3f9GPKtU7bpv1X1U2K
TvcmUA83EO4P8aCK5Tsu75mnDrjFlgSK8FVIHP6qSVX3CcxIVqu8CSB7HvhdsKn4WxLbdufWQqg5
iKjlpSfDkFlS8fe6s91qhYDir776YvXxYBRAJGwv2FUggC88VMF3lSHkWiGDXWFeJ9iv2d6yi46c
qUo1hiKJ2dnLOfGtxwpGZNr0+/Gq9jGv3++GIutbHLva1ngtoQn7FVLiOl9ndrJVdJoApxPR72Ez
Waxl9Ej73UeXMrZINGiUgOPDTzHmYnhZHlBKfmWaM78b6LzMwZz9j3fGCabthqPNchI6CiaB19ni
RfT0rHZB5/0VRZ7m7n32cZzX9yjIent+9XP3g54/XDLBXUClntWF8RpPQLxq7cLk46tfPZ3I9Bfq
iQiPOlUjcesWe7s4MC8P0MADxABN2g0zW/RoNSt2gcKM/3Glei61ovtDfUkC9h9QDLA1h6WHQwY4
okuBwqx8LPmGdfqz39M8I5I+Pqr2ulyGDfXaUiD9jV91Y+QN3ijcSFqzVZfUopYhDcJx574wE6PI
Tug54xaAEi+MvpIxDVCc366UIImANLCr7cghOKb/pa4xtwMWeE/F2CpArJnAmDB1k65GjFAt3Z8W
JjRxMbZOm7ljynqKMQa2/0+ijcBSHt9UgzfkRr9qBbs/wHgENhl5qBZlU2tLcGCP16JyNtVoIVQo
vfHRh5rXZ/ixGx5oQL3kc+Oyt0a8TOZMETwD2TGWVvnAhS7NF328JEWDsav6yijMnn02q9ar0ky1
LIyQa2p+RP9oZcomPCYsY5sv5iY8gRjZv2FsJOQ+UbF4qRQFnYtE5633DVVwlWqylaowLbKp0dBb
pQQm9WWGF2J4QjfNwTcmB2k/EFX2yDWpZvR6ogGiFsy//XddvN43oS/1NVKUuaOVqv7/Qa/MbSqL
AZeldET6+QoRFFHaGQK6I/jiwWkSkD4R9bJ2vuYL18jUcHqnDvHUZ9AEr+V8ZfWPZB9DFlxkHdm1
MuMqe03MkT7PfVud8jtLBOagsoFWu0ik6EriBj05Oben5VyPs9O2QKOJvi702zbCWsCPS3/ea7zr
zC8yhPBAkbNP+FAwGmsWL8cGSDOLJ1zztJ7YbxaBUOgrDyJUTA9BVycqwSwil8PBv6jZHrf/0rxp
R8LsIuPb885NJYSF9sec5LqINRHxnpRup+6AWiBo1l1OkG8rhQNO8cwSTCRHIbLmRSt8p050MGa9
yOyZR8z9cFtQvUJ/2xGVHAbdM5wMMSY/Llo0mip+lTR8Xl4ADcOBG9iQbDQ1miJCsJJ2tgPKaiSW
PU4vyaupxXG88RusQn9OMBj6xQZZrKcNvKSE/ETr5+3HbAxYOAKe17JegHPAobUSWzNzf7MNifxG
30Z+v/ptiT2JMU7LOo0v3sMg73oPxrYs9oynAl9jcyeUg+fUxrP2UeVC0l4luV/x1nI9kj58AJJE
CNkPvM+Q474F+Hi+oiK1ntVsabYlOlmSJaai97uR+GscM2E0wuUwS9FVon90zFytLGe7DYa84JiR
5ScbHIRoh4iSJgpUBZnWiPTlF2V7B0z08bHR30iZWvIuAYRXQa/Bl0gk4/7oi8QJHCN8zCeFFM3y
a+3xluRrM0oL8nk6/GfXNw6+sZQ2UxDIkxRuOSnr8tfTbyfyunU1RcgxNqV6x7SC0hhgH7rtSBsJ
co/BGGYA/ghpjGz5Bb95Vle3zwfffHbTrIfRnEH+OqccTMghCs76ddbwYZsF9FRwj5cFR/jahpvs
/TdPhWu9mED0i9G05EKPCkDoHQTPABkzXbXLeuyqpIzJc6oGjSW6fu0W0zX8PzefNH9Dyc4fCUuo
Bjn6vy3GYEMgk8B8cLG1inis7r/FfOqr+JvvmzZgueNkWIBqilxy+O58gyIVg6Q/eY3d1shG53mJ
l6hc0FutdLMS8zobnQbjqNykJzn8Ww4kJJWfA3aGuJ68PpbyuXABAt095/Z8Olvb+3r1wOwsmndx
HIDlDubalu1Cw9GBzSQBXrbrf6829dviwBrYk03ZJlZIu9AzbR9MMct+Tp0EXjfvG4bnirnYX9cs
NUVij+98QOxapCE/aRtqeS0KTl94ILWXtpuDwhFoQ0eW+elK+r/jNRyVnfAL9csVZlRqFGdwgGrX
/nbTrUIBIsZ66rysknyfMUEfpHANwIWHcA+bCufUPye6Nii3bYx2TrQ0GMf3XBM0v3qFf4EEgqF9
ZfB5nC3fFOqRjgETd3lodkXB495A5AS6NY6oIvXGC+/GaDSgS8mJMU2dUEnHBkEBbFlizeNbK8f7
xuCf97jrieEGK8C6DqT3UNY965cT8W/Y05/9d/6ZJDoBajQ6GA6xaqbRFtc/9d3CW8i2FZ2mpKr4
hRkEoIvELPL5AqBvpwRfspqfDqNax0vA7pangMuNG1Jc9hvbIo+Ko4kGaN9g8UfbbxC9GMVzCimn
6dLhEEmSuSCyIuqmZzabDvOD54A+TDfn39h2cnMoPZQp4eX2trsIv8R2Lo3Gpk4+4cIkT9WMkyva
ZIOLI39c2igOAesqTJsXtnElWX1f9jdrOmYhTjYwD3s2JzC1YPUrhNRlRoO0eTuO44f2EfnM3RZ1
HAehivApu72iB5kDi57fGEm4BeWX4O30+4JU8VL0l9cz+OwAEWo0CfTEnfiHC37W9b3ZDSizVBsW
K3mJ+sa5e3TmOaRpGOp4tmzU7YIwpFzOEBX/iNu8fuLO01xjBXeWcDchwzLn0YAgCNk12fEJ1zYw
EVgR3ZUxuyZc9chgtvkiU+W/phHyKMxQ1hkdxAOuUfuTViCpD33sR29QcQwc8GB7shcxAeZyNpew
kxXr/vMlQQycqpElpvuADdijP8WMtPJ917BrAk6HnmJP5K2wzYvztVE8S+K+BweVpjDfe6eFG5ZQ
xx6eVp4sssJemzK6vfxmGL0C1NEs91JzuubeNHxNYpqT2s0XnZWeJnbJepQ43aMTIThgv+AOo1dP
Rg+uBXJ1kg14azQlTXb48W1o5Ghtf48vEInmD+sisqztbfnN5kqk+PxSOq7h8qLFrmhBJ/qf6yvv
O0gx12GWuMSMhQcfmJhkdDMm/kUZxEmK87CYfk+vw7S9aVQozetJ4PfbmDGcp7ffMImMH0LGcMn8
jMcR1hh6X5pmQarRwxu3m3YrDPcVNFeSX2iUEBgke3euStjNxQPRKBEe1Qsfxom23Xn0VLmCiqNe
E5QoN54bONfxFZMPjQlD7Xmng5IThfaoMYSJVeKCTJw0nfNBunp8JcHfQdEhKdFWhbpU+PrzYRfl
qV1HLrGqHn3bcZszenV/xrRIDosVaqSkEXM+RnpiqumNBMkVOoL0Pkph4YbVa+wozS2PvVTd55B6
Zckwb1jJN6liL5h2c4QdrGVlt3NZqpILyOaIf83HtnTsHJtvIvntkxYj+ePwy6nDfxYtoOCwzaF3
+Wl96J/7DuBsB7zNr7Ny+qIqv3iisurwRUXWuqJY7yBBSWkkfucaFgckV5kxC7mwP6uSlJO0rubS
qIGmdB+cGYLWuYOpB7TAb7vRxRA8v74bxMkvSSee5Lu/6CTUtVu5tzW7vsqIT2jlxwAhyM5ovJmM
3GlD7k1PFTVlYzOZKB362AETtz7D9gTNHuDeoKdN2S9mOeihneoyFlBkNRd+66te8kU0lPYpZDBM
tk1X6nghZFmZk9McKivXOFvHkUjQ8TtfM6qjA1RTp6plw2e9XMUCCUsuWrueXgNEqubID10nMcNk
yKxe724Z2+EgpyQ7q4Xay1GMNAJIsu7KAhDOkR1wLoXJ8FbotgLgKm5aXpxTypyweNO5fVenKJos
UidXosqxxvoHNUf63J6+dZA12ifjta8Ci8I/7hpfRAa2PKo/cL9GSIhhEiETnJp7u6TjSPR/boBe
4YANeapdTYgrlDmIle7Kkj9MyhvaluQg+yk154ZpLgOonb8M1lx/FJq1i7wtpYuMk9D4/mFa7BvA
aiVjgnB0FAPKfGQmvvdTZ/8wAIdaXRHbPU1XPUm5KpouTu4KWUHerdBcxvKlITLhyoLZySOmRbBb
W26eSqi9jKgjzRUADS0nVx4miatTKV54e7pf1ooz8My1tTg0ekMcqQenpGrfwF5rZncte8orLg3L
lzkTcApmRjeCZTEUdAAesewgY0qqjJCUq/Dor0KnKJwS8sgdatAZpyw7ZqdQF8BOI/uYRXviAW10
RLtxNW4lrJLY7E3WhAHr9tRwUmCxPxBYCZ4rVjQuTq08peuRActBtltZiXc6DcXJJAeNWnJqAlwF
Rek/VAMpvn8bg1xXb5jvilY+dKNwno0L+cSeRvHIlHK8O1w1ZB05rDKcwAXsOx/dK6tF97xTTkhi
YMfs3LGCfoGC6d4QUaJrI9DcjNYiJTpg3hJwwdLjE+RrEMSrtgtVHIxZuyF5yy8P18tJsW0h3KDe
v3M2Dn8VFWcgz7ycaSXUiLqBDG56ius90WMMdlKAlHE12zyRUAXIDYqpEcPygXlUVKO9e+Y5Cwob
1TGDElQ2v81g8GEIMpRpJsQknunhL5wB8W/M1miKOiBBiivxapoq3aWeStA1rvqtEKvXYYSdcbD+
3/+wek9znVeOyn5aKMhkvNcdg+16LPQMUeE3PiOJCFCDZgWXe5ezZYLcH8uOqRoFluMTZyViTNuc
2oxI/E9Mo0xeXxmrBVdfqoD+hYHKQ8JW4LsuteKp2FLdsibTHOpy9tLSqbLm3BqKc59oP1COxyow
NViyTCKr8gmzZjWtytmp/FqbVrWiUtI/GWEr79OZz4u/GWKa7ezU5px3wN85TSqRMLNqIgp72ni8
UveDvLA+geiQQ/6Ne79xeuWvyO0KVeVRCUs0taVdzGlRbRk8ijoDAQsdd+rJCsMgc21Jp9ttyGEQ
LWdx7X8ssIH2faJZPkP3HVAN3VfyfmS3Kzmamxeax9wdzyR/UXLPBE8xzB/WoSUBqAf21lzHOfy3
qv3zs+2TiLVGKO2MTzlKO5I0jnxaXeq7lGX+WyQPYBHodtbgDO3OaQDAh5a/FKF1/mr+wA2YkVWa
SlIjm4m3K0JjHGq3mPrwUdkRBXtVizPe9KbiF0t3VMjFbvo8i/OTrkyyfLJeJH87sNdDxDDlRSXv
S95PSj3amKt3U3F5Opw20HA08NIVdeqaTe6zgeLO1phtnn5s1Yf36zFhTZGGJ3xcMTcFFuQhxlLr
8cLqc6zy0cEssB1qvv1IkUgySJsQudOo+690EY6RmNWG9xlGpWm4l48RKbzXP2IJZLKsd1bK6Mrk
oqxHE4vr0hhlEL6gUz1VCS7EOS2VZ5tJ3f8VHXpccqfbdRyD0Z1vh8MlLafbwHjSoabMgbhmw+gz
e9ZGnv9DuvKtsLMQACGlVWGpZK09dkFYg176YW11BpOwp/v9nM6Mz1/nEH4VNysXMHRAjMN2dmkn
4ebEvLd1j4OV89C06tgf1mnUWpxWRyaHC0Bm7ZP5G0i+bSWDeIO7TcKlPeEw4KmLXIR5TbhF42Jk
qftHxX3fNfGOyV65yQLxMJxzESiubHiczhFIiz6qyGZR3PB6q2jtxcbmp+6xED4PycejXZQb6Pow
vc5f9/3zoPnwuX3Ofl89NXOJ99ge55mOxN9GSV/kCyb+e8QMXE/dgXBlR1wiv69rmarRPjeaXDYu
tN6we1vFsLM6oCjVQlrsLgjQ3y2KVZHUQIbJakAr+ACoozuyXhmk9q7gO/T1B3aBKpG5mXcxvZBl
P/WxfdZroyQUlxhJWVAcldHg0wMJ5HwqXbMwTlYDZg/FZfyPfQoHHQDrEUdckjN4R4B5lw0+YJN8
NO7vaqeH/Kz6mdcyODb7e+dlRG1SvbuOSyz3B5r3qDqdpAP159I5otCrIN5EC68s5FObpq/IhfZf
SWN+5969mVbGEDwlmW8Tj0rLjqLpKPb1DtUzgofFEUqachIqfjl8j/E6P7L2RuW9FwPhXkI1+Use
74TFTC7PHdMhGZ69R5oNGKwNW2UWtVFST7P4EfazgDBxAHFseeSwnN/W9Eurde/DKGpWBDw5rerV
AS0eE21Jq1gdxXpjMlq27kYJE3cHAQyGkn4zvsDmAim7awapzxqeXSfDC3mvtuuJQrbycRPhrkJ2
kDcsdXA6Gf40WC/n1paZ1rEKeQXsmTAb48wUAJU4d8JJhbwKOvmCmJ2AaSNuBrYtTcLdk0u+FnCI
HmJfclEHcQQappocEHZ1jI1f+hpuKjl47Vr8buq4wCkiyYsA51m5KwBJ6JBgHvKeEu0MyQK834ii
gu7ybTIQhiqgwuFvM2rjNg0Go7LD934FF53BM/kZsxB17f0LklgEVwlbPCmhG6ocPihcv3uoXy7m
qmOp7qBYz/F5hYCWAx28Nt7OGn0bAIbkarrwUrKqo73BHaCy0IsDlZcMJZAsMIzzwnk+iuGAmrBS
CWm39OEbOfYF8paiZciESgfHJXDu12rh+Y+J7f0vpru4wdXJe0R13sPmslyJ9CMVgysccGZ4xDQY
6AMmI6F1Kt0MnSvhFFhXxvOWr8kqS4aIsSnXbjobSc+5Y+Q1rLdLlDwow3PqPOAkCUt+qh5JMsYG
/T5iHv/aMQzEw/Q78oY8h7V1pxxXExyWP1vuBcCkl/C6zQacH8Z8tHAbjXRW9iQ3Y6GFYmzIGb8d
di9tHo16L1ZbZdHtziFi5TAMePH6xf1J50pc6zDpHraGXTu+IXRm1ZUYUGNg9NGdS5b6v0lyu0Ao
LEP2O1RNs8VDqOd5VXDMCqVTwcGciYtyrOd/gOyl42mwM1vNcfsZ1NLXuethgE2MODZK3lrDE5pP
+G832V8J4xyRGZYli7TUyyWjOuUqSL4BgfIvbLOMfTMj4a8A59ArijCkGhJololhcvMvUuiWcaoO
PACNET91saz6KxFNGiwFuzcizk11F105X33h2erPLIDAqTPgoAe0BTkdDYa4wkrKh+740H2jb+w/
y+VwTqLLSR3tr1Y3i0oJRIv6XZlBKZJSwCQzLHnYAqm6/v5ga3AtGTULGuB7IoQb/lYXCYwKvB+J
HtTMdKwZPa2Gd//3ZB2J7RJz1MQ+ig3Vy4DTY3Hg7m/YiWww91ZXmZVCQyDoJNIA4sJ4ExXHOaZn
uvDHOMeN34WGwb6ivkB9NJ9naMuJ1sq2P0xhVO0ndr6f1nJNgFIYxTpzEfWZTCAKhSzJ8by+Vy3u
RjvnZy42xmTaA2CybFC+sBh4XVBhLN8IRjjVg7yjvDHdJlO5kLn6K4FTDJExjA9LsGLXly72I1JH
vURUbhZKULDxEb2EgKY/dXgSebK8WnYjVnFIn9qiCbWvu+Sowf8gQzwDfunjQNV5JmzmN0fASft5
+3giEjAahVCaf3Nqj5n+2p/ez+i1LG4eVxdIsV6YxoM8EB33440dybSvfbM+YDaUKrt1lcIzjCs+
uAE8T4yyNCjsUWJoLYopwkIK/sOuf7hsdGm1bIIe1ZlIo6b6PXIZGXIK6/y25kk/f/rSDBmwxJq1
5HLbRaQWMnfBwePLlGuE12RMsi28BFXKferULU8OJg2jRjmXjEg9b0twD8XbEODLcyrytRFSrakl
yJMjpT1pMkjWmV/BiwuWEJCVpwYohtxiKTDCgv1Oul5m4WksmWZ/dh1x5OGwnUhTk2V/2OsAhbXk
ACMUz8j/SEin3dTA668dNFEQJioGhOaiO6/WazlOslKU2y/30pz2sFlvStS6+yPZGS72qd9UYyHU
zCtTnUrfsFDMUJHg+uvO4AWu6Jcv40vsUmVaoX0xNdnhOUXALjU7UZRVUvGXM+NiQViatqDcs+We
TD3K9MMWE/LQfBZ1HeFgt9moY3LrpX4MYre5eOnkpirbH2Dc9V3Jynhx1zfBwUImEIFI2+6aVJmt
YcPT+EFWfFE02qMkoBl2b+L/cw2H0cXkUrqVq27/oC/+4vJUnrjs5wWg4a0ZI2YyiLGj4pKJVwgW
5/5a8bmdC1Rd7niXn3cT8ZJYu0oGgGTtQkQX9ctDwcjMX9a3DBqaUboFt5R0loaPatdTb+dctwxa
viHR1aRr1KDmkH7rEtuJ3CRN+1DT91yrRakZclyz1RHrd7mq1oSxR8JMs2Iao/kqnTCqnDjdmHsR
+pecAuaBQsnK+MsRxTn5Kg+zJLQMIU5gWOsyp2v619Bau5q5F09/GMX892JJqox33XWJh3nwKtxo
q4gaORLqtmCTs+gZ4QhOxH38pMZtWA2VlDpPWFLzCZbRu3aQBMmjNith97rQ7s21bDDl6lSw5kyf
3cDMFMkK7RME9wWRvYlYYXKho9Hmwuw6MjJPSZBbJqYxaJA8/tSsB4P8wPY6lO36yf8vZY2u53d9
8K147l3sufcOgmuQhPit1vDriOVpTydsyOkEBcqCN+m2NvmIYD6Ky1SEA1FvocC3HObDfAk6+qOu
vIzCKfD/HJ51UviQrnsByTdYRw9aexgcmWoVSaKBWU/aBJ8aVj6BXbGtmydBP0kVneDnMhiQQ3W2
SXRJTYLrxv9wltJIx6LQ3W6W37Yi46Ay3zPcXWYHTuO6pzTEySVwmpydKQ86Y0NwwO7RGfu+ySwi
b7xzA5BdJ1E05QSQrq8+ZcE4qr4aY4rR5OnSSMU9tIikS2uqmp/5kqf7JpyIJigpQ+RWZOblIWkn
CJFO7PLSLK2ROTLqKcrxCmgTMT+Aadtmkwc1kg7WwEn7tgFuzVVWXFNB96dtYjQ+7NItsXoECeTo
XDla1m3nzS5RgcWeIp84MHT9bX0PyY4j9AIRImMVjJjx9woSdWp3W8qrOk/giR1z8sKEmA4UwaEL
BMKuURs6VguoNivs39b+lpg5KFoLYCLgyyFfAycQIg3dBlOuPhKZPismGawdf18mUvKI4dfluUwF
C0U7KIKibk10igQ74/cV/7aElB1D78Y++DwkbvNSEdDBgrIEDAWtSyRrKlmYABTncVY/Xb4kitgN
RKcX7oMkwr84w74wCKmOeVT6Dr/Kzjdm3W860uTuceAGXUSXJugEALwSaBNIZdgYa8Vji8/9pysu
GFfbrIFlz4wnJL9r40/3IYsMUTCOqlFyTNlPTULRpona+IUxp+6PzhxtMNZCpH4GDokmXap+R/h4
lIyxZidG57J2JrXktCbY2lIQyK8YhoU46c2zdrR/BGFP3PyDzVtFFHosc0MDK25fELQQQNzr3+m1
VqjPEWU3pihdKzIB6LPrMODQgx5qvgjFxndEzTek+2Qfjws3Ie05T+YJWKg4K4gycBnYry7KPg39
LWWJmef1wIPKrC87PuakAC2nFLSfVZ5m542yF1TUJ2brMUpcZoMJsqOj9k2pIdw9uL5HCtMJTvp8
NW9QSZptSUVaHkdGgcocKzHy82Ro6lav7OOqyHzd3EsN48XgWUZnpjGjNczAIsXoaicGcLE1SJIf
Lp/a8cVmNGoViExkgaHCrCVyxnuFOwqjc6I2ZmIaoavyq73Vftg4YF+xSxAc2aEHTwl9aKKaQfpC
IRV5rAxSKUQC/Z1l9S45REl4sQrOFkAyxtJZKRuTWQ/QwUiEDSKIHn+BBRVmNV2+wiCmygecicRV
x0a8v+wEPDFGMuWctMFsj7gaf6oMEe9Gbfhxy8sTxwU6Qp+jMTUOLR8ZUSrcK6IKhW++VFI8d4uW
2TCgdEAyx/HljEHH1c1qOenEwYgS7dOprknmlCeqQkS7S4uclSESr/WhLq5d75kKRA4l+CapGD3a
9pBoe9ohmYodC7FeDQCAde4hHYY68vnwwc0Jb3DKXpSdf5KqK8bbG1Krko/Om8a+ES/32GsQsRYt
6iHDKKTRnP9Pk3P2kd7+r5vnLELaJEKpstRTpEaQratZBHGYuBEr8pOzWQaLf0oD6UxjKOaZAyds
X3X7pls7k0glrB5Ms/vYtiXha67DCl9VnU/KTci7pJnf8U68+JjzoOCPk8w6GjK2T+gxnsNPCVF+
s0YNfXaIdg1o5tLvGZFYjrAu0szS6BVTOizAgXiv38EUqHsUYG9O07DqZAsH8H4a1c0HgNg83yc9
yzqgXq35TGsW86d0AwWiwxnB1kJQUWwLqKdOeEz0/8eXXFuBT8mTG49EEWzJEJX8OpXgS6ZpHluf
zuC40soeH+csfBJ3k0AZmTr380BETgBgfuYtral1IijnMSu5unJSoxk16CsaXL2ipxBu3MZc9Ick
rngKlO1fiTlfnxJCkoPWvOkqM939a6tynMBwRpd5WRZ1y3oAj2do8tBT0cTC/GUr288s3azaMX5I
mUdtB9O1jJEyRKqAHnMunPWA74APTB62EnESVUirO5m7eEXJJVFnHUB2m8eg60L3SAFHe4cqE01c
rUGoOtYojrJJ3xbSa9qxO0Se9by4vOxqpM09VW+qWDBcuVfc/ZZrADDtULxF2sWPcNSmvW8xlkPT
GRk3k2ajrMXSWCEuMlf+NHcH1HFeFNythKNeAc8kOEjbVQm9YTCeJ+/4EHrsHm4YtVghByo1I3zO
RQfcg3L3+bt9VTytZJ8HlCcPnHX6AGdVh+FpmZT+NhYg5ovQQRbrmqnrixyIchTHz5Hk8AwldtG4
T8vxuHq2xj3Md9aAU8pMvKkn9Fiz7mWTx5fm+QYib0wVQ8Wv9eqN3tkLH5paMinZrYd4nakBETsQ
nz3Fc6ulnRS+pOGuBf9U/zsnTM4JVHKUQqrqdm8547D8uPPOd3cNXiF39YTTugSN4FT8dYRM60M+
Snu3sW0R98AzelB/oQ0o4UkdDRubPVShKog3zOjt3++iuZkg7CWCy+7067rQiiA2fHYC7a+kywP2
YVSMJsxFgkAAYcqV8YvROusT1d/TgK4qaDs4J0Xz2GOLYlNE3TmYjgHQAylJB0qZ+qndcvvPCI1a
jDDaCkI8C8KHbdm+OAXh/aKDJ+pwV7JSSlCXA7XJvF1owZVqCCsT/fYFaKx1L4UuBWxJKtxveqm2
aPGF+edeP4QR3Fo51X8TLeIUXwANj96t1xmWlz+7O9/ljBwi0VOocc5qtvJ1NiPnSONRTaMOzdAy
TCPHxGIKQixmWx83Eai9bMduzUQJyhmO++9oc7tj8eZTxRwJxFMUJfmMUhsnVjtJSAbbteGZaRal
+2p3VbxhT55x0SsLN7n77KTcS/KOlgGjpdcmh7q20cpRrRRWTPeFS2hpUALPSLZf1ymhO1Zhati8
aXDQ7J/8AtAU4EFC+HzPtmPPD/ZdcwCNWu2pkylh3mTMSWOBvJmbdUw6dAod2U2jyGH1q35TQkgZ
i1IHLIZeXfyzGCDIldWCzVGSTUZ7ey8731fUB1s0GUKS8N6USJauFxJMo+Gv20HXNIFyo7NKveTO
C69An87hN73x4aNNVHAZRbqF2VfyUnB0eBuoBnNPZNRL8l9aVS7fjm2wulBebrKS6/d7h0GxKn0N
6MUGakQYSHfRMd7szMw4iSE67nVqIpKTz2TaEpec0Oh1qpcsRHaR3iXp1Rs9J/hCDiyHx6bEvQlt
3O4MGKtFkaz/DdxZMXAQib5c8yE4rVQeE6ISRk4812kmFH1pVy88HzUHRzfLcsxk4a4dFg9pMg1i
7NrcFcP1+/5fUbCBXMfW7Fku4bHJKJ/Iu9o7laaIrg7c91wVX2u7tVYcHbcfbyo5LdJ00yyj8tB+
K5AcmuIkEL/NhuRj0sk6T4+fC0GF0Yi+wU6xDJJBWlwyqysQ4bgRTkRSGeOccZ6/zuYDkTYJfNtd
HibspfKBj1fSksACRyaj7BfP3yKteS15ddFpar2Izb114yys8n4ch4gRvbMhMVc1uavNu/u/KEa9
jT107sgt4XYwqqzjv4rNZkx3MNiFrHUMrt07V8ZQofgsW+12APLZhLl/fsQjzLspJz/JF5ZzVfzW
rQBVZmdcLTcTUwDAwnBO7v1XDGAcV8GQQDlHw6a2wLyzfbNp5VROS5ocNrGy7ImpfXNgJOz+49Ot
DabRB1z1u/dxF2E0i0MUSrOlBOi3CAfKPxfo4I8yU/x62IIA68G6VAfuwLu6EFjtnIs3FZP677wG
OE8SgpyDwV1MPGef4awLDMv0YBlyyAdwisq9r+3uf9MMDFZooCEndAyPll+Zn24mfirwpcvdgtdG
4yU50mjRa3vCSbGqfPCy+YETxgm4EgkYtULyFKiOIOt7DJ6MrWrlTKaRAvu5TBEPVZ7K2Kn5Z7bc
O5d8ZaBkE/8sBJ8KQ4JQQyzCPDg4eMHUhKdaoJkUYonka+KnFhgZyv8DqVbYWSeOJIUDnkSUdNtz
O4FeAtapzPFW2EHWSfdgJgABD/Y0SCMnbL9rTotsDN+HmNPCcVgQDmGu79gotJLWP5SvBQMm5vmY
Qin/uG+IbEdHjg0fS2TfnuQqel+Dz0PH8c6JOKEZg9/6nFiX80e5Jz77ySEfmZrnOOwGZYwMeVbA
NqbG1aqRlwnWIjOLyxqfiJqZmTRtiP8RRMeoiZTPPEYd1p9PKcXzwJ/qWlQ1rvy/wPYnRsoT4FOk
E94dp51QsxFfd0PjVqy/Aixfgi1ReLxJ9n1a3vvT99zKkPXaqwZDpnK72tIzTN0uE1kzM8OHi4KJ
rDqzdcCNTVH/fW7PtdEiUR7isYqqCqyLpEmTK9g784f9rqBQwodT3Ro87p09rCcN/ZgwsvDF8e7t
3Nqm/TZobe8Jti59ZI1B85zbE3bWvyE1tbMfUcQhBt1Tnydb00ECBBcl/LWNwCeFVZ5dm/xn0wZx
vxudJlRuadL6Tlt+tKlAhQ8qa7bZKYDdhUWL3sr0QQVVUaAw86HOKToYPAvRFwaO31GPnNSt4CQu
O6j7SCxf5xybS/rU+xtQ3IMzt/kj1uuTX9X57M6hhSsy/ZzpLWP35Sy1Ix/MqUBdKiT5zZmpLQTD
t73F8RjblHKxoGMH5zrLvbOPzVZk7VEBMLZcbuo7D+P4aiJtSoCFhpW7gjREQvnxDtdtTsE+YsWt
ca4AKju7AKYblqz3m49WtldAmn00v8ARBtC9OqeCAqLvby7e3TNSgLFMuNmB6UB8vZsximz4egEx
NZX9G1t5asCZFXugk79EAwFqklMQXrl3BGWoUzEz6xuBxMFfSBsvPHS4Lh9mqKxzcfUtVLA/aC4L
o45tGjoEBFODZbyWS2FlokLOneC28WkT5dOzEeES6NfGLbltPk4cFE/gNlyFsE7ot9KjJGVMnKbi
wktZwfnSTBE54MGM6/TnhV4KCZ3e+KgJW2kjneZp79haRWpcMiurMb0tB6COOMZLmedKjAzSwqVQ
OE5+JV1RZZQEIiwldZHoBPIipd+kz4NxWHjccb5Tu7kDmcqULghQx/nyEhlBB0QF1m78tfCPidza
ZffoNyXYTNqtucvukUAIkts5m/QLVs1QiI4HP1RtO+I+VNPULkGqFdx2loidFd+IJTssUwjpc2jN
o1PhriPzxruBhK0CCY0lJBScOf/Z05Mk/ZG1TMcC21OikszLJLTql+RMrGQSxx5a52e4WQGaAoBT
Is65UXXeZ4mILfwPPhdoXydmEaUBD4Io0qV7paWabFdH/fkXLDP1W/+mmffyn98dfLoFbjzszP5J
SJj6jwsmkqFPRpTJlJO1YtQSdarY3U4IQf21arFcoVHUjCQQbGt4OIxqtWQ1Z/Rz+nGQaU5Arel6
90Cx7lRFVgrVme//ezABoTgN/ibqVqsEqOPgXUo/aKBam8xrorT1S2/FtlCfBmLolY+fDvWb4Zmk
PcwK+eQRvW3WmGyPn+SNFojD6A9watVu1BM2DkTF54AP2EIV4TYFU6rWD8VoZ0KMWIM3ko1JahI8
nHyXFmBJK+4++eQ7XWSPTyxLXgow9hUqQYVVCFgGai86tuiT9Nv2Qtc9vqfy5dQJrIyeqEzo7WuD
bC56sNd6oQUKeZXKSzqCUi3S2YmPxJrnX76sjkpUTyNB4PJECMTVLhf5I1CRBXFMpc1TWyllEL4j
ismM33cdrm4ylVWvMlDX1BmYetE8V6cdFPz43Q+wumoVMfUEDzsvKcRaoAQFj8f8sRKNDnnHbZwz
zqLMrjpbfFSMdhKccFaMX1UfduJQZheyNji7Vk3qG/QSURWX6H/rIC5HEJD1RK5QxVdsjFHL+/f9
5uvTZk199eF+9wHrPbCcTqSJhSbzbNOg6gjG0A+I3IJ3lIb09rBfDN9o4LP9Ko1wHAGHF85RKK9q
9kFvak1TigEX7KeyQIvTF2VZYP/qzkc9lqkp4mCxvlxdBbbP+63DmA+9088BIszjfJBG+LAOWTBd
ay5y6/8/5WvQYwK9HmBfxDOKXorpejXafYVrZwuuiD9r+DMBeyPgqIwtdUL7VmSHXliOxiu8kTWN
+3/eiaTbM8axZ+ai+VhoHrtPJ8WzxYTBMqGTRqnvfTif8Evh6aMLLjuMRCRcD0ctyQKKu2P5yys+
616Y/I28+8xq9npuE0rkQKOrzUwnPDsWyvRfizVTK2XDnwg9s861UgvZDkHoN24YjFWnT/ZZqSH5
rEGwq6ACy/5QJ8VSWXS7Tt4zNeH+qve0a0p9HLHnCm2HZMOZGSsDb9tLC3B3McK6Bo/bFy3tWXOp
NEFugtXjW97inYoFmfE80Af3GUsEr2FDppZSRFKY8y5oWhnEGFPJ3Nx6suNU5O4cmkUWdjGgIw6+
c1SaybF8epo834kOKvCm+DilD4qYU9xq25SLdEbVG6mJG/XuC4qVg79G6+l/4GNFdP2+TJNP/os5
8ofQH0rBLyALw5Lrr+UVcfck0jHcM5Zegv1jOpa+7+LpyX/P3ZRmxfPacenChjIpSBsJU+kmYCO1
YxvNB19vS6kYgQodbD97IQDc323LBfhLWMap/MVpk1UcaCOTcLD+ozrDQ+U3hhTrqcxUWTYSoWBy
INp5pjP3TerKbuzaNfS16dwiBl08woJl5XQzp8cFAQn/m9YP0WYCKeYLaQniqe8pXjnKvGKsYyne
S2hv7dC1BHXgcXnkI83jyAeL5oeVs2C3h6Wk6g2OpElLTleDyRb0lFhYi2FBY2UrbVVpF1GVzSO+
hMDVdeCa/O+KhTHo7o6+O3/PxJ7Ah1mB5h9J8AbRDwxaaOxuxZMrcjp78yRrqFGEQnf4qElqaISZ
UvUIvUD01KISMeUdevwR4aCl9JdQ+gx6eazMxIqBDhP6FAt4rkLz6dU48FrN+dKBxF8+uqhjhwyD
RNFjPVvSMxQ3gvGRe37KDVSEhBwYiEyHIuyrc+c9NLVRSgOg7UTICvCMJTiDdPqYDsyLranU0961
lZ0UZ/mPOvTHc8OpxGIMInEL8fRDVe1MbQV7CRxzEpgytr366pJFuBL9ATgRjOXxiJoPGNxgRSNh
ZnW1Tv0LNX9na/WjWd7ROYXprETpXpk90SFHw1iustTS5ejW9dh6H1L/OcUbHCDp6rNlAxeyaHQK
ob7X4BGctm+/7aeje1bN9+xsZrgKyvQVd5JGgun4XYDyQda+VOgd75LoAXYEVDLkn9RpLe81vcfn
fUas2X9CbYRLrXH7ByhMJ8JmqkPvHyulcQbcTJj5uVCCZZbDbzdtPQ4gDjWn8MzSVMK9Hk+Lyp0e
VD9JptkEQ0ECShxsQ+5JQxJwPfj1ySWtqB1gO1oz6fBsm3+HR9bOx37sgskt2g8wtIfGThlIXkMP
hzGkUQLJ3uZz/OHD5TFcD6sxG5tWzqJOZ6vG6lNGH7yAtFmPKzC6HF9E6vVCDnbWX4GmyTwS/auu
pmXdDrxYIx9yhqr/qC5flZzYU69KcTRS7yaS8NUWFiem5tF+h0A4EzjQ1ls3DPFfquchRxi4YrVt
wLiATTCAotSeuUkCibdAC2T2daFllEhTW2Ws5OJKfJoiJ/TshxbItrtLHtWnJLaAEsJ2hMEV4+Jb
QdlDEwaKxzI0lxhDYr53H1rgisjsP+Yxo2dk5b/hIuXo6SDnnUHBN1uGoIofpLcoT5HqHVmK4826
7QiZkkZOMc9zmdn8HLic4aTTjTUZ922/c3rx/Cb97bXVDhkIYIowSYvhUhZPMfKXNdu7FFFebR/b
Rr0jJO4lInZdvJGyh03QBkq93oQaoXXMaItasmDnVmPk8+hoKicqemA9BzuWQt+OZqxY/bZH0M8a
gNqqBKOUFnt+AA4oTozsHCNhFxdOfKKO1tTAxG4MAmby44Ie+bcGHzmxVqaFrPHr76HasNNmdqGH
4eMz6rq6ZlhAtct2Vex7VNYm9BEjpLjpntfQ1GQ12sHNgFOREl92iVjO3mvpj7fz5yRkNdMDtLhl
+Ul5Xx8pHkh9jykv5OrDyW8vfjV4FGWIT8is+H4Qet8nyPRGdNZLh4EzofA/d6eyI5wlN5GZVU1O
GX9htLy4MASRpvGIYAqfeMA0Ykf+Qcr2eeS50AUIQoHWRTQimOvkZHrj8n+yBIbovOXruOsaCwYR
SsZvjrWiEG6Ubi52Rmwm/nnlMf7njErppsAU1gVUWocHquq0eYOXYKg8fZ8UmHj60VG/YLpX/skm
SR5cMruMNVm+8tNsIYv6GsIiz3Mj8NOSHT8VuODDdWCJ/upHLVaxF6X4T+76TNQYabyh87WCkpTo
xbpmMWzhQyZaGMMt5SNd6eySCQtTSEOiTjRfnnarMK6syC9PBTVdLrcddPQ1jGB02HMkw4ahrsQ3
C6SP06oPJ8daIzpPPpGg+OEQAsK1kD7H9PrnWLyMogTqf+bAZZyWmvjzYd6A39VrWp2SwyuoNsUO
K/PTCkb7Bp4ZkFWh/sdJ6zUDmH+azJ2m4hEtrygIDyxcEcTBBF9K2itM8ISBXtg/RG1ujE0wIlze
EXBoxH0sXdFgxhpWVfhJcHlJ2jt3UuoL+x3fMeVUEQNHI2wHUDXsmlbSasvjGQBLVXxmDijl7uO1
zUGGnoczPRDt5PeydJER3eH/H5sBO5K2K2eEnwXuM7PQbvCTZfcjnFYHDm0S0BI6WTd+UZjQUCG8
ZmqHSar1PCwLankrSAI8PoOu5nT+NSmxN27H3ySq0Wrfx1O8kniilpaV39tglfd3zm7RiX4MWE+K
rKu7twAf/Phy3g89K48pK/NpQNbYEUHUgX8MdJU8g/dUbgg1aw/kpbqGNYHqPe0m4FN6lSAEXN8w
dN0DGMc6TK7NiPBbXTVeHoRRsG0YkXUKTYhs69//vkEHdVr5xWjORtzlM0RvAU9frHqXH9/vVQRy
S0oQuto+nPBFRV0jlX6vJ5F0P3bGcommMxCrLQUqBkvDpAhbM5qFSYjfW9CvGWLyqnsgZN2ezPjo
Jq5SVqRvBxUz4Dcx3evRIdrY666LN6mtnoJ5hC1oCemNMGkZ7ggAGF7mfUEvxwTUUnB2Aq0JhWIW
oTgsVfHVRmvXg4FqQL5+JhXlgAbOlM3eQbQXsTs170Yaax/Ywo5aMiQU2vER8/PfKd6M8TnbjmvS
Fqb1wM+SBuLBx6a/UaTuuSWf+1u9kI5ugum/ZH+ZvVVsot8vDBnJGVMXM0SSul0HXlHburm5r3vv
Na5rrtUVZKmfRhzVtgqK1IinGZ3Z6bsIhrGU1MPdBX5e2qJGA7lLkuMppJp5WKMEpm2ODWiTBjez
lCTB+danyy8ZTWc/2p2ZRDgVpHFGoGbyPbErgSjnGcngrg44GL6U26onEeIYUksXB8UHque1yBbb
UoQCFimyRDYjSs6VfzjkCcIk1IY/dcfepkmleLowvlBqyo1yi+ixX8mdeHcywWCy31jGSLDnkv0X
9ro8jU/eApl4EhRcYvf2cG5uy0Lr3aE1tkr7WrMfzdeeGH8LS0hxNdn9cqGJdpUbgRWLMlEFB9Kx
obVA7GKC3HJ92LQeceT4Hap3SQpe5/tmXWCjRW9XViNokBRZHp/UJaKTUsP2GYW8u1IB7Dki/cRj
jg/HGfEPfGV+4i9VxxfpJvlnZUD7utjTJjBomNKydI88fuyt4T5QTn7t1RPiM6Uxw+LAlcGyLVU4
bjM5+pK23rh6cqe9OaFnWJOiYeKG2xrK/LKgtlNpVs1To/9oZxQJYlkYxDRg52i3/gvZleahxBmT
iUsBtWTULvUMuf8ZEBHcKQiI+LffMqg3XTzSZRN7in7l9bk8kGJMiOVVhhmSRd2tr89T4hebwtG+
rHYirJNz5+Oplh266KS0ROQ4P8GQL+pyYF0dT5DA+34KHmtZoy5lWdMLWzc7gX+RqNtYMAN/Gp/p
grZ2Koa9RapkAM8ZtNmnVrJWrGI1V6v4zE6q9SRyVIi6obkQeUSWT14FYfHg18xXia7TY8J4d2Gp
u65RfM3jmtuugBmJfc32CxtNPSMlAkl/6BmtXjJV17StVspiO2eENPaHSkHkVxxYTD8B62DZSX7G
cSBfI8gvaLI2Jr5msKJHP8xUswnhm0KGR02jcCApSkoJEuPlapxL0RXYs62Gwchfn5lX2oYaN6Ll
TsZSqPJMxCfkckXCQ0omMESVTgfCx2hT4PR1byqAIX3NGPWFYSaAHVWzQiv7hG6/SXW/X4nd7fKH
Jj7HW4/pmAPo5ahrAN0NdQH4RkKZFFX+Z1kquIvaDZXZAOR89hsftxSbs8yEoIdzmKOGU8ATZzQP
IXBP5CuOmAR7jXCgU07DOb1zlUSCE+k88PExaanGF9E+sjeR9BTCdX05g4VrAdvYdAtsQFh0l3Qh
vL9nJMTlnBHzjc33ZxkHSl5T6Csa1vRIsrDLreFU1Bp/Qd/HGN6ufL8yJ+LGhKFhidUhLlsJwxxz
IydTefBBnvKhVZcbyDUOliV5HayxGbrxDsmJfkWbA6yLQDNvA9Yci8gSi2clnUfiOm5xBjfOiXzY
8ZwnvQbOFdaeFrloVcoG4ZqR4RfPXkKMu5dSekINOYiQgn6BIZuqjtIl24ndkk0fo/2IcEsMnsoC
Z41flRZIJnlOSTl0wxLtsBLnF+IZ9eaYETqBrYPy7zSvBCGFdC2l7ZjcOHxzPiN3IU619T5inLDl
B/63/3+/M9g2A8B6xm90C4gF5rFeHCz436EegebvM4LfFwsaQq2l3bDtH5aNVyF1uwEB4M/DemUP
K2/7B/ZIPA5uBsq/8Dem9be1UCuNQI2I2xE8DIp39gTKqLrqagyx8JNuebPDJGeZOd3p2+gxzgfG
T3XqA1dW82uC57eeZlMEOAkO4492pi5/wrHJWvlMn0WOm9wKi+6AIWociPFuj1z2D2DNVHf7aNdr
mlyDL73P210d7dDKgmiehWC/QP6BMyJ5s14fwL9IGq8KZ54KYmxMXnFNG4GjeHhoU6i6YGNRgspA
/K79uYsCdcjbEWBktun1lCAnH6m9aQAyUY4aCjucQW4/WOTc/9TJ0z7BTOBT04CMGj0z/xl9oYWE
EpARkHPSdhNsQ03v0snjDkjWgtNtZnwUILntNeMSonq13FVAwbaqd+2MZ3kNJE0nJe8GGFu/uca0
1P1kyp1DuG6oo3NHl2/HIq5hkFGfDVK4cXis8TJoDGe/e4eXMT9k14gsX3kLc9p10xP3rebw4yjc
+qwgd027DlxybhDgVG3y23kKiaB64vcGNueyJCDLplUEU8g6DPUhC9EWVBkZc3q7gOXccCe+iGbn
c5WcTKUUl3otBNqhbx5MJMjcByCjlzHg0uMGgxY21826StF3jVmox33LWrHYwfg/LR/OMMKO/e/A
sD4vxQ++0+02NfpYCmV7aS8VkiNJZYeatNYqTAv3aRRl3AkURp09DApGbAAzO0NfiPTb4t/JWxzD
4QwrK1gO435V/EFS4mj2UPZnNcqzu95gZdWlOPzDHeg15WWA+Os7YdV/G7Oky5taPP8vTn6zu47O
Dsanl6J2Xe8XTe0AHW+HhnQyLyQK93nr0IQuGcJLFIR9VA2vi9+0YZh/SMIAo4yBebTkcG6KDBQ/
ovnn/UyohBdioLhjLy31t+UDwawh5w/ZpKIzeHFb5EKmdK1dpsG7tpNGpO/rw3eifF0bqtaDEDOk
aBY03DZKLtkpM3pFj+VxiKe+m11oC3OsG84sJxTCKBUiYep80sg1NU9a7PtfDFCsNTnc0qt4zLDj
m7BtSU4+R/xdFsY7zt1VMqemQMa0KF2s7yD6fCgu+qn7qkSORWYlSgZAzL97EQ6DjcutzYKu9FwD
5+KaxNINzCXnvZpRs2Mh8xowcZAuZdldTV4c+WBnoj9EpZDrntIJZU93xXA/klD0Kdz6ny/E5Uby
BpMsIrIsUMI+RrY3XDQux5HE3ue6iuQVbC4f3QWLc+uGoTKwiNZug2+OILcO+UChf2WBg97NAAkU
sRFwp5WIB/FT0TIrb55AZKmsb82DzzcjNyfOAKx/BD37/tXvhGpf5s1h7dDQ2481fXLTYx7DGxkw
mfTdoUdRz6NN0ZmfKlSzZHFYqmIKhDrMphAXjbFnB50W0eK4FXrl1yR46AhKKZB0AfyEOlxmztCE
VtcT7gaVcari6EtqhZ7XaLYiCaIb96iWcUIdRyeMhumtaJj8pCsuWY1KIeUUYYb+UAjRJKpidOFd
msB0SqjxwjMxuwxAOWycLjcc7G83nxmo8w1AiRVCEdTbitkr1L8Seh9ON36Rahbf7ZIaXNfj9CGa
uZKhAj1KwnRe+VvXxMa8gdfahH/JSvioliLr/m/D19+a0R7EkxfeTrO9RY67re/tF2MlBPQxbLqo
4DHPxFEPZl6iaO15kqr7py1scpBFs8HeVEi33aOBNFi+A9/PpHRKdQeDb49LgLkKlFRSyVzYjqqb
4Jj85Dze26wxNxZCzfinUiIh6s1raFZQQNYvmIgFGBBu6nzrLO0D6EHVbo5z15yrIjdeSoODSS4/
5USwbOL5dZofK/3j66cBHu5uxJENgKazoabwnaKrBn0CRGjVj2q73e1FOXFYJFCKHfys+0e6THwM
uaWSRoPKV9QQKk1ASYuzP+e72XzQBwe72Qdqk9O7U0wZhLKNPIOysh+ipvPmPFZvb9cl4Jd7AFOj
O4clpUnlT1UT7SjHbyB19vkkchziB0QZoHketRGIiW5JWyCzPXIM67kOgPDcEmUEjK08cF0vhueg
EnEb3OA1lMFUsm444jvWA7JZF7NKnB0/8oV0EmS7fNqUXcP4in+tbrrNQqII+rrtTlCbulAgLnDN
RgV5Mgr4fwtwBWCJXEGd8l2FbeQAs5RCt+8HE7T10YeLTGO6+37r8IbaixIZjdkJlxyzUWjd9r4o
BoQbHtFUuCcBNzEu9srsWfUls79QWpuLCbgNVDh5sthAW/U41SUraxpys85j2J+LzPk1NAr8vB8Q
5I0MQwjKdBZX1uWmVhBcHFJQl3s6Ljw00iZ98vSMzXOBWEWBt+VE3UMUmHmwl0Y2xTvtKGZZyaMY
8i6m1EeCwe4FMo4ZggiWnuY0vU3Gkeaambz2KR2hADJORCvmhc2nN7eJ2pOROHfETl2KOZZjaaj0
mg8rc35HnklKHQT2xWCVUcwN+518i/7nvxEbIyAFmoAbFV2IuiaarlJ+v1oOIyAo+DRhQgUam5sG
3WStqkihP+N5xqek5FXWkKhh8V2n2qmx1kB9s8CDmQpppL39n0u8HfR1zhXkxubabbLCuzAFJkOU
izUylUiF+Kp6jYSLQJdJRBUZgXYdBsojAgPP/ia+VbK/WQ6jjeEGmkf9LRMuVcOBN5at7XoJIRqd
La3oBpDnPcAVwM7/LHW6hgXZAA2J2mRpBPVEV5mMLuN4eOUeNNVF3k5aZiUzO5Wcj/SqE/OmpNLc
G/IYzyVIl9y3gk+SMUcjeVrhgK9AOffuFZ/LsnHm2tWjtJ/r3SQYgHA40rSBUoeLsVGWV8Sx93dH
y8b3iBHjblfj7xmMh0vAd+BOQlsHBQDPdjWUKE+nmqSVwsXvvmdDInu8SyUx5jYUBe/k3f4mkhDl
2xAl0aCsWvJFUhxgOCrMBUo+UZaGpOpiPEF3cCgQnK4+bDsOWhAvdJV9J7z6jgRKc/yVFTnlzxmh
F48LK4/QXOmGqfWhdIhfM4s3d0w8x8LcGrSPDAp8t77thMZJ5D5TCKbri8p0ISQQLniUq0w0AuMJ
/uEAL+g6feCUSIr62+LL+rRA6Q5xiMqhDl3ei78GU2jsQMMdxYuPXlxNF2Gm8N/lydSMrTSfiZYC
TVCCVS6t3h4/6bgeY1oEJc7KhFm5jlQKbpLEhfM/CckdcgHFcwCHwVsXa6VzUoy9SyzJDjtE4ZgR
BlvWy2e9BZzKQlr8L4LSIaAVj6Dy98WOfFgnj/AiHyS5Uj30kOolc+Kfi2w5TpdVulDGQqrUK1ti
gNrXfPBqwt7lSdz0KqI+VlC1MuzDx+/vVX1sFGWm2wRrLZrNEPkfZJfIscNRymS3vHiPtweIzaSK
ncuFsFn8HFgf/KB2uc89cRIuhd163nbSqWl/jbM87raucbH3LTPJSVxkz+HoZC9KzxN5NlFqVf8v
BngBPs5eTfZapmoYSn9EYBBh8G9NSU5/PZRsIAC/0zcgFncVLAQbYtL4FRJ40MsMmSJYyLTkTGox
pbmkatsDi6KYJHHdF+vGJCOZkINS/zNvq4jCBVBp9Zc1o4Gyh7UCvdv0ODHjjET7YXEsnK/xEhWP
pOeJnVNlzUUrgR4ow5Az2uvIEEUzrOIOHGx1sx/gdFbsCwhGe6dzVGMNzozdx3BEPQAetVV23hGH
fcxR8uc4xXdBJaFzMivIGaYUkLLYQ8e16pDW9A4aGGeCTMPyyJ8VL64jSYAh+Hgzzgg8laqJ8d+8
KpA5ISNbkEKrv5rgTtqYtchaFD+cSHSTxr02PUcGEJh+Ly3EZ0PNnx1D/XUJ9TQmH07D5rXlTlpE
W5rdSrtUVjU+6GRh/5pKxL4w3FROmLEzjxgwOg82SOYv3p7mCEsuQwO0+rPGNENvhtsJ7jcBc1I0
kVo/vD6kcuU7XpAP8XaJP7GAmE9x/4VSxuC7PsCNwCA6L0QeyrfNWFN8/+vItFv/GY5XL8n9b6kd
TPW2UN2JGxu9FJj6+Z5lZvso12aEI2nuhvtgjdiRjYW/ZPDftyoVni7Y+RbWfW9LGzwu1JzYi6oF
kqjkF7EbfHrhMA9XPCuOTFucVlf7XyY0aAjNq/r/EwLnrOpSlE5MeIBri1Wqi7+UmrY38YnkXSmZ
9Hy+/y2PhTincyAVEd+lxkfw/E7O/jEJi+hlWG9AloI3mK32+e4uhJcGIlrKmWwyQ+ohjafGcFry
0RBUG1xbC5ND50iLEgobvlzJLe6S4nNw/ESs+w12zX5mqB/NU5TZLdVdS+4pi83qm8jMjWzoSW3g
PfyTNWE0+WDTGLDVZEG1iiHX7hZztoG9QoV64kVDtYKT+U2aIf752wycHwLuEzEPs/fB4KV8ymOv
z5Dd+t90quKaD5v30lnh/Phzmh9QDcTpFxbID8F3Lv0oF6Ta9qfJv8anxpBCXst4TPSqxt3Ija+P
6AqB0FyNwE19uB2BcaeXh25WC4EvHjNMQY0qJyTVInjZ3GvjB1o6v24TYW+tq2//yv2A23OxRxL8
KgKoC1E6dLS4/jMN+diPWCcJni2pqjEzzch7OlJET1/LOz/ir9U/vLwSo9ic6JUEnoTt/+QXoeJe
2u+4un5/2C2mpwxevzBgco3aZxtEclQppOWtC2a9mo3uVNiulsHuH7cMcr918p89yUV898efySPh
T3xo3xDogCsHagaArtvR1EAFChs3+IHIkZ1oiD1yO7AhRss93GG7vRe9mMFTlxpiiIa81DEvMFZx
pJiUyDBdneI/3Nzx0fFnY84HPJ50nXrUGm6hMXaWbdbgQInRSSDj7J5FIBCtxeM3OuAbHMipZG5h
VXquCu/b2e83U7fRounGslQyXAFFHWIOfV9V3MII73TK6jtLNbS7uy7dwwoWT83JaghQgH2dUar8
TJnmnPbzkxkdSeTDwnlB7uyesweUeLT+nkRT1ybORr0y5kfO26onxKhSaa0/ZJPDWLl0QbSRmL6f
b8mXs/eElpI1UIr9U5bZ3hDk9TWNCDurWSo2NJJXFTWDss5ibKs3za0NipRM2HJLelk+/7thg5AD
n3SGxWuY+aO/HMKXy+Ce3OQkn0xynRqISgYjUeQQmZZploo6zK88ri2MZdo4sbSpVyBLIRLiM7yK
rJ+5/ps8wj3pVzXzzpBsF7KZOkBpyZfH7aVoBwlYLs1vFv9n1CkWVDYMCGvsxTA+KuvWC9DWhg6s
QxuFQposoPdW625FkZGKF7H9UKcJezVMqlMbtWAuX4VHG47CpKzbDW168+kIkA5bjj6LzAnrd0u/
ehq1hK4opSBXGBn/0kpU8oIRGPBMCT69J42XhdtGhIbgR1KUG/o8q21Kwf8VOOHpTSZBff+xGN0K
j1iXokPp7PkboVeSvXtNvZoxyReTdAbAjFXkh8oOqBODOa3XuXCBYzpx3eEY3RfUeAFOjEsWmaz4
AG+cQpriRtaNDr54q9zUeld+UGoswGwoWaSB6QqEi3G20Z1JAXSDtKqn30OlbZ51JLSh4N1YMiup
V3NMT5+LI1RZ3jZIV6Ww/SVLzhlGc6jNGqk/MGq/AXNecSpqcelPRU/JyJnGdJJ9xdh/iEpHRFnp
JOV6Fq+atmTOpLtIdCx0M7C3eXgJbV6djiskkurPZwKVvwUVOKE4SScEvT7f7p8KmM/LMoOg0b+O
6DXzDYTOdSvARFGkn4uhwHadnvX1kjstlJr5XDRWox7qgSRo+FhxtUaVj8KHHTp4d1tSuSLqmJM7
ZrMCvbwLY9FaPslxRYc1GiGENm5GyCGrM6Em6LdEyxlGKy1H1BdL3UrUt53VY7AOOWL81PIVV7k6
HfX2u7zvwxoEB2N4eaUppkEsGWHw/3tkXxY83Y6Q4kC5F3ILoeczAnp62cZ6dV1Aqafe8IA82zh6
Nou6N9exmitbcdplud/zobX4api6EDT09V7v3eCQrir1MBY9g15jVPMyISOgZRbzLBDq/CnaUHb4
AKBzU5S9EtGW5NhsCcf5snaMJbWpBC2V9Ridh1zup+vPA6ttdJHFv7eUlgcc7TdyfU5FuaESdiTr
s2m9LubhijUYIAcEGe+ODwTzcDJs27q4ElA42SgA0uREVGvwvs1zpKP9izWMrc+vqbcw5ub4aDlM
9fO7Wmi0xeWedcilzXq46NoQIe7MvzEQeTPihSL2918i3L3uI+0rLlJUC8SCK7Ud1mBlz4O1YeV8
uirJ/35085xOuRpSYCKJBEAFDM+P3gctfae6suKFuL4ROXo+dkMGRk0cEkoyPjeXIlhkFZbAcR7S
t7IVSuPyksyajrUitxxPk2KH2VDLkfJQXZ74KzjhY9o2BiUtKKHfEX1fzY0CSF/9LlOA5Du4KqCw
kJFGJwnOf7GnLIQ1OqlegpNsu+BBHuo2e0rQzdLmmSUBtGKNmSFGgh9Q9luSPMgxnJEx+kfdAk1p
ODWk5ROmztP2c7h93+fuK1YmZnOzVOhmewtrRu0QF40hTewdLSiR9p7tt5uDre4JKrTKadrXdJP8
MYEab9x7H408I4uLohws1E2iRyFwapP6BhCRsl7kJgNvXBIx6jqw0cV9RNvuZPOom9hkjuMGlzW2
ZviwUUGFvxFRokTSttOVJFmw/8fNBxF2Gyx4EDwxHjpkAqxWBxKRoKjkQZJ0m0871IuXkrPc+EHx
+IBvJDWVUZPxATYVB11JjSvRaNZkDV/L5/3UDhw30DuOnhkQXBczQwAPVsKrmyxZ2TICG/kkAiLJ
ZZZl+8E3NCi6Vc6Lef+OjJGvCU6rHa2XSKFphXcQtqVsR+mf55Na0Xzpm0agYyq9r1YGgmTqPGd+
R4wcDNPg4X5FtseOnx2wX72yrckbFKyfJe1l1exAP3aVFfljBCC5Cb/cR/hV1gsRTsh/bfldq9dT
5D4DSviiRnZuDQvLojVj9sDgPCc28uhYcoEgsfh6Cdx9L/A1VIMzWN6iAUEK7HCnXds5HxLrVAQN
VmkDfVqwEYJ0ZrAly+CIfw/E7qgEh7QoD9i5o6xsMzNtKp8g3uaVD7Y71oij2oWdVw5itoIkAWNQ
1rWXT1yZm7zq/5c2e5nhKZwtLqrVojcd1CLAITt/UfGkSs3DAZpd1Iw+W2zsVG7fm3OXHZnoULqa
FPPSgFezpyVSI1SctcGHUzIsmdEtC/bGJFJqFOdwqNRMbnnWdUdVNzWppu5LI4LEwrrIqrTH3dTS
WDvhRHpSyVTlBCmKhpTqBIwdb/9mPEtFUNtRX+hKr5S/3yZuk8VgnXURoUH6PcM2WZPXpQRanLkw
iMObHBQG4t90DNXHDAxe/bod7NknZX2yo8MNDEEXk2URdHidawrAYJrKXS/iRqo5nu7QonAyOEiG
SJDDmEyNC9hmOrJK7q5Zy/uXQPte4i4104e2C7ya2bj5hnVMTj4r1/v1RIjnmnLw8H24N0sqeSHa
BS2bD/dNCdDykZcuolISwDOILyC46KohBWbCtMiQRHPAKt21zoVXcU2j5k9FwDCb/30ZsNEl2f5Q
uJNPZwj/f8sm7r3ee38xM7s13WlFNIVGc1aGcPt7F4H4BhOmohVrmKMpPYU7TFkvajd9dilhHJ8v
3DmLbLg5gooR65prZdWH+ED4Z3WQvHZm3pYTE/gwuJRNIj+m/Jz8r1L5PmbUL3oorC+4odg7BT8S
XJL/UQhINDe5SoZphOxktyl1Cu6IWPdmWl3B5xCKI4A15we5cXoaqbDUbcFp2JRfKR98nW/qCcwt
CiA5sdF4mduiHfv6Ah9k12G0p3pKLtA6MiqzN9e8WfYgSKCtwb1B9NMaS2N0Ob+gENby/FAuVjGT
kj7ruozulI9BnD8IK6ZGKuEOOKZAfGBTyelFdYkGZZyYkpX6IJuGDT3vcWRzYCWvDjVmDzFPijjj
vJXMVXVWn/21amgXUPmrcaeBDE74YHCIbAhBCosOMXeY+I4xPjRYGL/9PwIF6W+LxZmRJ4l1chZl
teX0WTvnu+akhQZs12Y5AJLt6yty+t8I7K7/c7sWcELpvtwwtYI3diNyR3weAckKVwOrlKP6BLrf
xwvht44+Wxx39Z4tRGDNFUqCvdkqikjx1xLMNiNdO767LbuGrEN6sYja8JtDzcb7Zdj8y4NVhN7/
dHd/cd0bObPcIKPoQdzvBs+N3riJypmk/rA6Vz+7ucUpxgFKtFTRtBRsPqJkOIDTcWiiRhuDbGKm
IwAV6Wh5xRyvl4G1UO0VBPBv/VSw7u4ZRyEdUIRTEINuHu/Mwh0+53wiJERSVyTEgcbkOjPeDSGO
JeE9q+le19A1GCdBqMf5Z3eWqw3HlzB3M4ndF7nL858C4qPxiT7eNcD6AUTQ/cIdvqW+41oFCabw
FnNvxWY3QnvKL6B+z78cgI+lk/J5WarqDWRvpgWoWfiar4mDxAWUO4/utS2xrKDTj1peHNbPtg0h
sETgRGyTpWxyE8oBwraAsGg7iG8n+P9oRHQGeoVUgPzgUFUSTCkUuDyfpR+OlYmWypSCv51jwA+n
cRIwXb4bdNuhgyyt4/DMZCInjp+QbQlbPItCx3AyBbDgxC1MtKiCSENYzdoYNPKYdrSJoo67NV+W
McMtK2FtM6mrYxxpR2+TNlHV5sRqY90Ka0wKWn03dGh1wkw62U3sp4iT+UH2kdyP2UW3sJ+1ARTM
ZEze4jhEL2JUEynoHCUM9RuOlQRdxFH4B1bts3xVzvgWTpO+ys0uGsu2GAoHqIglgk/OE00rTI0i
LKyIzdKaizA37ujC0dXzn0hGYEZuKfZyB/Dx9k0GjKv2oEBsDqLUhC4u+1KAzOVeOM0zBTxC0gFH
rAHFfQr7n39lW/AJnwlWZP/n2sgEh0bSpFvnVonzutIRVgNnUeBfLXTPzHzyrW3O7KFaa2SCDPZ7
Egkb3X8swf7hOMPNbv1qlSDYjn7QRajYi7AWaZ2sm8wrVM5UMqxiOiLnGWa2XWf8eVqLIa+wGOvI
7kc39Tpm7yb8MxFvrkgDPTQAuKfkrHYpWwkhbVpGzK5iOvW8RLTDyGrvwy2uA7UJPRNeJIYiDE3l
EF3c3uzO3TTMNAglsNBLGQckyhrtPoWqgzQ8KXiZulqHngOUVskK0GYnrcrvXpgQEMptf/Jr7ZMU
8LWO4NOe0zmnDG+Ex18hrv9nR3cmTj3ztnFGwjHF07lGqm/i9rbXbiTWgbWtnGPUV6ARlonTnx7S
GSPMstUoa/ZvyG9iagnlEUmts+17g9NMMbs/RAIPYQYfe3qHgZpCW41icpLsLslOmS1PBfuPm9gg
EN8VF3K4fplucb6U1VfgObzN3JhvGYafqBewuzvBY/TlBe1WSbaiZ4xWEFHc2H8LS1y97AC/fpqQ
5cDaBv8MGbNLtQ6x3v7mtIWo3ZO01FGzx/0rxKHpkFH858SAfkoOg7/apDNfy5bfWv2QmOoDBy2M
CTeqlXF/g5m1L+jfHUPSonL5FP9F2D23yJAWmXrs40BVN0298PHqccM+K6DEFOt+K8cMTBOPYer/
yyoJcua/hPfmGqnyC5Jy/MaZz+0u63denrUDzk+6IjjaHnX/L+MFd62ZVwBKZqt/9jhHlI+NHeIK
lIKFtMxhm+n79XQ9jODZbnRbjYsxilnZMUoRk3LrYC2MrjJuvlRdu0syR49azPH7ym8FdwVG3YTA
pdeWau3uVNDNh9kZHkwRCZmexuO8Zw7W828NHx201l7N6xbBRbo+3qvSXflp2Q2HSyGk90k69+vB
05/3EhQI3Pbm3d3jrL7dFkRfxr9SeE8Q4EnGf4l4MXKWyR9prSS46iZTcflQJKJPShusVEjGs6d9
9vXj4WS+pSAOSBIOJZOsI8BZt7tb13n/WNSqlvvsjhgV9JmvVm6zjK8p4qsreIopb177XdigX9nP
bqfVE4Dn4vHFid56g6Hls6TXS5XKEjCjoT6Xtfes8YmZfbbKSt19MdK3FKu413EphPkfMTbq37R9
rb4bbhPPMEH1ozOKkgWotwOMUw/BtrHw7wKGDNxioEAdDypAZQEu+04CdsgvFLsZa5P7N+FG0E9y
R8RV1gJuQAw5QUkA4TmLc4xMe2pKnL7RzelylVFzLA0OgkAnFNFuetJM5DeDqAwO0hvvLH7pG25D
QXyjnwqrGslllDKIVQymh+7Q4DaztUjbSBW5ez/TMYduJ8DO84PyplTbhFxwAlC6RccfmfFrJOUw
yvpLRrz9/Gw9ovB/OllOjoSogwp9Y0U2hDzF3tw5WKoJ2Uhbwcq99Y+XE0RRiIiCagZ2P97I1z8F
qysbDZBOK9no+kmUmSZ9zlha9qsGFWY6gidQs/9B2XCLD65jUsRuTH38hdtegpUsD4OnrzQVtt8N
D015f7u5uGkm5hOmGdESjEdc9eNPF106xvUvMTHpEfCYwysBR3IDnZhHiQaAIe2eqEjWzpbeN/FK
ic1feX3WJFx9LUbxhmou9fNxC5iKrLpPkVQ6EBLWxCnYujQPG6JMOArrIckV1AgpFB7vN4oK++S/
BjZ4QJfswphSmXEcEGb4GJaeLJeSGnPIweRrHktG0l4ynIhuf5JSpN2AiamvtCMiOvIVQ1MeFECh
NU0sfs71EowW/HbhhNjSb975QMjGDqSOcmrj2vscxNbRUfKVJLtiyzrGVvc0Z/TtP8Ty+kLnNRfF
eWb5qwCJd5Cnun2j3yZzag8qsA140kZ6pgwSelv098K3gdq0P6jsBTCbKiQR1sUr1OWEg73BGL5O
VqNsOU1B2lZmgxUgr+UMi38OYPcHD79/2buD9Bmc1GxcQ9EeQpZHtCbiXTzw1loH62qoG2uEcHt2
tFkpl8EQuNKYQU2gNdJjb4/GQlDqLcs/DyqNrzeZEpmHl5l002TBc2VMbDSPf48ICFFzOBpb+Ffp
N4CvtzYG8mAPUWBR5r5eIUjfr98Js9rmRHJzYrHtTINh3S4aYEHLvARp7/ddP4f7eDit2+jfBM4X
lzpZYtzvgXifvwqr0SS0mo9ZsJyTjKhHu2SAFfb1otMBsSSeDCaonyROa8mcEyWEQvAzGcRhgRiI
ejK+kPVJlK2I2KqXlC2Ir9VzFdv+kjLtED9tV7XqjAXHpPEaXsecC+Gp3I2iDqyRBe9dLtmqck8t
KMFfScaOls7701DBuoqoa9WYxLfvp7peA/iCdW6DP4acAcqnH5kZlkxCtHYMUz7bP7FCXZjVUIGU
7SbtdlPbTnzKNYlX6fWm3+rZp7IJaoDmCCEB3Nff/PLpQYjMf24rNquJ1VQLEnaNQDcFIntL0NO9
L7ar/gbcfvM9x4PWM38EWfLhFmWlenWLWyVBCsstHreO9Bpj4Dy4PVHJC7vkI/LkluvEjHxsi9o4
4qrxaosuKQi5FKFlEbutIh6gpSwZgc0fQlxwvbSn/mgbzv9xsspElCMiEQFUVoT7jQcL4R1ivwau
1FOFAlSsUXtIaoFU/KLUM3nmLcNx85myG6OZFfdJk+j2sZrN+dI3N9gesldu4/D+LIEL/1GoLuAM
9OdodaUFic62imJzutOFxIomU57wzVjNdWjhwxh/UjCFB3Uy1s+TTKWRY+NsokgjCjBSvmes6rbe
PYOisS4DwJ/RPbowDnfqJUyk2q4VuLkEGu6w57SfqPBF+6pE0LgSzcVCiVwe2utoKj94Fa8FkQPz
9MXyoE3M6I9sJDXlzNrlnnicCQmlr/YXa9eztlyu+o4I6ZiBImw2KN7dy2MGti5+3oAwBRHdmbjI
fkYSI1NXuN8w3Y6KRqL6c2/6mf8Xy6cEuv4GyQe6RcXQ6J6Vcul7PA2bSsg7POg8uX/82cjt2mia
D8AD4TxNj7d5eRhgTep05WpZdJRDGqDj7dyTHikVWQkcXEDE0zVdZzaC1S45Y7uBDhA9DnvyQHIt
TuWaVzjuXoVK8wkxTA/u0ti9fEB36/Dn53dmYl7S2TbdIOSYlkV4LeDquPR0DDfaJceJJ8H1AmQY
ZHlWwSwJEiVHkd+f2ZeDzpEFDseJWzTZCo+I8b1eW1aw1V8QXnf/VYvOIXCbi/eb9+t4gwbBgYq/
itc3azvdbAn0k/C8XDUIvH55nUbwtYW4hJD72FxrLG4/bGO0Pu0dAIMfDhXDbvJ9k8xT3WY3M92O
oXZLNGd1G9Xo3VCbZvlJeZVmEX7qMZpw7LE+1TXmSGGPUD12bTm6EjlrUiAJrJ5+IqrnidNp7amH
j1tp0bda0ReBIpzhQN87mOnk0+E/+1hvQXig02kbOAn8h0iqjo459/+VvsD91GWN5fi+j89F1+YV
qDwxBthWu2Ax2lKq1Rmb7NpJeHsRINzF5qUcWYqv7Vo0/DO45/ndP4ZAUixVptEY18+0/sRPqtCi
h9xYYSADJCZ2ZWl5QjeRI1IU0kpYK5BNNbiQSHOhHu37qK0T59lQGEZufhDS5wvUze04/Z5tDnFn
vH7dN19DJ20QZeM8MMchJ/wTJVdqlWbgSaaasF9cae/l2fgxMrPPjb6Ds8jySOeDcl8JHQbg+/uC
knvgN1LiP2JpHRyGKXgN4Wa2lJAEwLnFRWqVVZAHvqadKQsPpP5RC4Jrjbpv2raHYqTZIVq/RkJv
4klisrxQXcFdb+Ezd16LACeoYHhjNBlG9eqh+7ltkTh/T6rF7qpKs04HygTrAIUskigz2/3qWijH
ddNxVl1Q9FoqI/WmdPThcO6ndNghrQ7FPisXg23mpUJ3KdBS8kO1EFAI6BJOyiH9vON4xDTx3Ql7
f3dK395R8gM+HGWK1aygsfjC0mhJodzabpAO/op2JMwVFXS+dgM+OVkl8h94OzmzVISLoPEm8+Ri
rNhalkcanUk1CxR5Fdr8FisaSlpFScUBJ12WNvxjWngy9r6GQHdyWam+PowM404v1kk7xXQMFNI2
gCxI/Mt+IaB0M4uoYEkR4P9ghrD97oLI1JtJ734+Mg/gDwl0seAg78DAtK+hPBGQZaDJgeBv/vbb
1vBcjO0TS4N5YvUanFHcWJMSBb7s0Wtd/MAzHwWHjJZyfe/P/iv9b4lxS4itsiR3QpgpDu0eqsfQ
7aqrmbtbQPa+NBx6koRZscRsyfNAZsianPn+Y2pQGy/b5L+/4yDBv4+Jk7MnTLE2TqwJn2HNAKb+
me7LyFfgG0Vn+NlM5LepQxibG7BtJyYyWmb7HxMMS1PPEo0je5EqdaSHr+UHJDOiUuOu2pGVi0n0
z7/f7Iurs5rr56r5/HQ/Zsa1JzoYlHGvI4H3/irgW5oOxchKzaBHkkmT3cJeqol9nngkGS5I3y9i
gupciOSN1hgkc1dGU68nNEmhfIFzWBJFGkToopusOaBoRYgwa8taj85HXXTvyvAyN+YYBdwT+WEY
XOCuuCMF8lsB5N3yov7sAhAZSSA83a3CWhPNv9Ap0j7oPpmUsYFN4hXpRI5Dtfmay8SusQqxwZg7
aMGPrlTIrBjYPQmnnDQODZhwEpf+OQLA09gZLDeexQek3F2KDJVtWPDiZ9VY0hj2fcBiLwWCPpwd
8cTVCs31tlCxzW979aClHuGEu3ep6tXooBSWXzcSnjnOXQOcrMBNxtGY6w6Q6CyU8DPdR2mRO9rM
Qkme7w4VWTfAPs6AZTgQQaxPNdjuEHTTGU6zmvooO6cnC3oXUUYQAsa1SI4+ZS1yHI8jqXXG81Du
GByPTRqyqPZZE1CaDfRpx7WZqTwoH7q5638uWfpodDuHZK4N9zssHAxWr3o9TJHZvr8c339CTd7h
rgOK3nK02H8syqO6dzAxhxRSaCvcLLHpxO+BhYjuu9sZa14yjkeo3yXzAysA5maMmoJyQ3zz8e1N
8E3du5CmzgG/tfASKKBj5wV1BqJRLM2CKw6CzfYWnC/eU3ko1L45ZWuCkm1YNvvlm4YHanift+TX
Jg7hEEp0m6xuw0LOBVVLu0vS0ul0vN8s4vMPjmfubCyaZD/t5OLJJaKyBPsxchuVZlENcVRBCRpW
2NXEt4UmGbkaSUUSj2rcjpt+lvMRsPyrMFIKzlz133cV5SlLVFVFHM0ueBte5NzMoZ04E98NB+cb
uJ1FNgV8aQz4eXCIqxJxyOu71dv/O5Rq8Zvfoki0KWjT9fm3rVZQhsE1lTrZ8DxcqUgrZQsX0aBN
feki3CYyBL9yO1Nd0KMR0oUaa5hBjIj2qVuG0otlR8ENI5+vB9UvgJclU4jPhC2QsOfw2E085Ts8
pWLDfA76FFrmzMvpSzagzIWoYRms7PVEK4/fKjNN3C9QflncdpovH7wEkVyh99BLUkHgBitPHLQv
ER/8Xn5xbtZ/9NyzaywCsT2Eiqsupag85ceUA/eZLkDjJWVrnpgvF9sXkabeH9j0hk/67O8exRKa
ZSk2SSa3gQ8Q8nxXusD9jXMuTMquaKBYdrcOFdRD4t62vJ0wBSBd/72HqyAKAnyJWePagGLjL7hy
bQwnlSRcflJXeFlQfi11HkvsYR293H2U68eVxAgROpUw6pdoaEFJRz2SDJOmx4a1n98VDD+eJ0Wj
GyK7+E3OVrWMaBrxsV6BYgny1MzSPwARrxgK0l3JwoUddqwpkiFoP6Vx3+PC+Kz511kgX/AFKPA9
KTrVmwc1iJvG7hLpsC640mAkEQbVRfUA1vjGdXgAIVlj0iGcYC61Ab/3/hzG1HSFdv9kSonK8erO
Tz9apm21/0cFwSorREp7UGZnWIm57myhdU7D4RxxZgGl15q5soU2I4l+CDRKP9jm7VUkaEgrAa/1
Lvb7sZUBysTwv6L9klD2ttkcr18tXvQ2J6MCpArbYgLbSem0UrbhrduyE48hdHNHrpcxls7aHJra
X0zOCNtvuT686VlP4eplWiNT/l0ckvSQzbXayXcMqsfAPhw0yi5Svkeem60hGDeyDd3zJTQwDrob
h8g23DlTx6082ezikLD0UokS+xD90RDEH9YTz91a93i0CZeA1WwIrI5LyuwSovPFCktz4ic+P1l2
kdRVArj26y7H/7YozpbrLdofvMTFNOZt16UVF2yo96s2uwblqBd1z1JUwIRYRt5PG5OdeWK5+6Gw
KVdQ4t3DfWzU/yHh12UpsGOq7beGDDX+XhFqhanpIciGJb1Zb8r4xeURpOSL8zkflILfw4V3okIr
9L/snpxA19oYec1+uNzzR2R0Zge2CeNIcSF3c/pIolWMVuCdTLriZ5Nt0thZGNA5KoyZDwlQ8gz3
F7JKdnfzJekAFNUNwfWQUWmGhHlyxj5b0yKhP7EaO3AluLuQOyY7Uce2CrPYTxxP+ra8qPJAvqVR
8Q+NmKmv9Kaj3wcYeYOpKpxQtEnGKoefaIaLaKD0HiOzonEXdRXRDuEzJqu57MhDFssjWScASnSA
RYeQOv4be/m1N/tKQsqOUS4CZbRRPcn585mKK2hmtKy9z/unNn6mdH7gjkRkPAnp31fAJyQJCyNl
h45milUWP9xLZYEgd8fsxehnhOSh5/HNnwZ9s+NulcLb4oprjvaLr9yjFN9FqJI5F4Fb+Z+uLHV3
Bb4W2X3ONYVHHIuUdJgLjYpqvf2l4jofAFa7vepi+Um8V8xVfIquk1lix3WjqFwmRQtjgcKWPnz6
2K9T4i99xiqvkFtk/tEaWGV169ojHHqnvEWC4PfwBbO95yV6guiMo/IH3K6S4S53fV3Jdwt+0C8c
mVKsvrWhVzIVswblOgpYKJ5bFur8a54UDM4fy0d9FHOCO5NUJj1tnGdYwM+Kaalb+2Ebxc8f+7FO
mQHqnIOFbBY1PLkFcqAXgo0kQubSzx65OMUbKsvAyOHtd8l5/Ee2QDlCje4CGw/SACw/FxXBvHNN
RgrGOjylvzVMbyJN8DSxNR6wY43y943MBumQV1HaxZ1AXvX3ivgRDEd8C423MHOkk1uDyH3bJzez
TuAXHOwv78sv9V2IMa6nQud2IvCgewmoN4e5TFMiDH4xdxcxdR//4SJgULDWv+4tuG2vuYhaSulS
1Erf6/+o9ysk0EuhVAinJKMExrCKQpXUYYYVWIAeqcwVEZgTeTuSk9raYMw8zl3I3HqU9UzpuiEu
jcDH4xnGyOabtEZNXMtNLsxJXhI2H4f081VrRZXwhYO5/9LH1zBXpoQvzYHb5ZA99hgtsRXU55Jj
AdJaqUklJulOssjyRy9n6wd4Bfmka+p8zXpgRa/DWQPt5iTusal809fUA8fCpB4HIXzuj5HMBvjh
Xnt8rQbKxwDAo3heR3NVaY4MYw5ezLsgul4c+G2IOUI5nhlsrgd6BrmGk8Zqbp+aTEhJ5+NT8/D0
0wvn1dYiMzR3e9A9PGSswghNRgKIrjgCNbOmgSpdV0idqTKHbLRgEpECZGtJoysL8DjRWloea5SG
7x5/wFO6d9+V4iPxU8BpNkeeZDC90rZisr/zm3zCtVreOJOSXmP5swgUqr83hAq0nw6KDtrx8a5T
k2fcqW6BOAP5ARnzOGIYPCRse/gZulL9FSCrJ5vsC3iO8WxJNjj+OS93bm6JCVkXAVG7NLV1JoMU
pKP0hEBSgYvN9PQQV9baWASIF09nQhlsf1ZZnww4xaqphYrKgwGDTfrkxnIGdjv21v0B+Uf48seh
sH59OgZiHnfENv6pv3D3dEdge8/TB80zo0jq2eAC67DLqjqMSMDALAZiWo7iHNzGlTiMJCQ+U7Q5
xz6n2i0xQiIm+/zDrMOqwwy7SbmCeXiuqwFN1NZeO0C3zrJc7Q0ACxFSLowrDwKvHSzzpXnAsPXS
8lNcFDEUE/jnPJG5kK7ekJcWIhqk/xCT++adGsY07Rego21uPLh+7B1U53ki+gNmykku7Hg73Nn9
LeQzU+PxnWW/eHTf2GjoZyaoKJHJv1z60Hah/m8pcmjcVwiZT8KjQAoiq2wMuvjACoqBOpGE15DF
ZMXlLw9b0uN3l73/jQen3o4QTRwYycaooGhzhc2Bi3zwYzmRPpJTLwPPfvOoSKnMYPtS9YQ8v2LE
Kgldvi/MCQtYSehDMNk4Ri/nm5R1XSwYG/yNBpzRUB8452kjL5jBly/wGDrLJkPItKbYaW0DQQhe
Q4OMgEyys2twQWa4jMTrhZ8nZUILtdG3pKvPgq/xVYyR1FJ3hapbfSNXwFTrkkQOlTCoaD/9q5sV
jd/NFgCzwHY3PpWnZ8HaU9E85Ro1gncigble0O6c1nFkFa6OLT4B5CNJHPU6ujRXFFbn1b9ckJ8e
KQtPp7Mjf//cPgqJ/dEBKEWEmu++SneqW2uR2DDoMjAn90MAVdYChRR2dbZcdOZOkHPB6ZB3/idV
4dDznSZaNEDksk/yy1BEL2Yw0KP7cA3xpKdM1r7jNYvjYry+kF4Hjg8poJ7eSdd0La6ZxjMUrNX3
ilL+rquBzYBoO4Q9w06iat06X1YeQKj2/FZ+TSaYI9DuaWGJ/9cmaM0Oq2E9QKhkK7Zsis5BoODE
CZ1/H5+soCYNFol4wNstJRypdjVIsv0lhlqcV9+ZiKOZaOZsKFzCgS6Doq4Z1JmWDOj/YtTqGV13
hCls9dRWaJOfMVGKiI5PexXuKutSewiFOWTad49UfmUVb/VOrXcdZgTBpZVMZrWl+aX1RsxwLm+b
LGWb61O8fMnMeS1diudMZ9EucWwSy8G4v440K7jM7XWoOYrRS7BAAxOKirJNV92qjBaDqYil0QOn
2m5U2gKYQjc3ln9r/yxz8oVC8xcy/Lu3sOum4incWVGAp/c9jSmHGzADxwmYhS7iAJFJPT86pSCf
jU91WbrxAmkLi6NB+8VDWMpUDZJ29dDjBdVz0IAwvv4nn26+wZqz2RbfARKhfTE+GMBkXn4Bgkhr
LZS0YGtgrLLRe34/5ksu4LdLhi0FTDozIpz0JVJG2DUPA9nWcC55mqivuwewUaeyGdIa6RVZKGyB
PwQuZlldcQKbim2nQ718+VWhag/8fdsnjeqlTdsu7cpwFCwT5EKWWZj/wTynoir4uOJJdmk5RVfk
L6oMUMBA0oYbVcoLgdJfX3+0M1zzKvHtvZ+Nw9azfHWNtGi2BSsQAZ9fcIThcfQ1JPYVVec0XAac
I8dwMGEUDD1TYRqMZBYgvCwps/C1Kc+VL5mDcnHM3HnBcT+gLKcCOvhf86GjY1IZk5tafOYWvIEQ
yC3HKHR8aRqfNXpmIKnD2IZJB6NGp6A9Sl+MEfEApYKEH2uMiGVvHPnlfL6oSHg8pC3HtpabWV3v
IXcDzBkCKXhuQa0gm6AEgsqabIkqMXptx27afjNLziMIzuyWtzeDZS/g+7HtgL5/lOo4nrbXyBuv
XWxiOFbr0KBrhUa8lXVVCoq7bqdly7Pvn7W82aZ0kRxBbNcAEEtS+QwZGuXrMWRirxETrEBhkMGH
xewaeKQvquEQMAXvc7wKCL2+TvIgfDuVSeIrtbud9nFP7rXIdO5/9r9ng0CKO32ea4bOyg5s+L4G
EKrOWop41yqvDof6Y9ICyx0J7pNSfZVgMwcOAFOBCRaxWHBFlBsU6aTaFGu3l/lELQLWKYWqFk50
W7oKCyb4+6tl7GlQOQU4vudUVg6qRZTTMtxpe9+0bDfv2esbiogGdycPTb4EtWm5mFbfrkyCuunu
gll35Yi9gfxGk3lPLXhPwrgdDbFbs9t8IauGnZqvYzwUrkVJr9RpF9ziUxLa00McBp07esUg8Ufg
Kn03kPB4TGBaXq2/F160Qpf9Dt/u8jpzVVGE3X9UGJS8aMTgDtsnyljQ88Sjo6snhLzVbJQOxOZW
ljBDNAawyEoZ6Jn8nDe0oPWUtcnH/Nni/5dfK8EMMOFTaN5H2FV221MI0vvoKylwSuAH2PCkVjU7
ZAG7ChWjLVCKZwP7vfQu8fxL4rf86L4z5GLtWSTTg9tikveU6M9u+s2xdVQcg/XmHgm3ZAogcDQ5
E3mYdrHCIvkb4zeVPqseWMwX6j+h+CM+B+AcO0kE4M8dOwoAhjCuHla0bmeGRMYoJnA/S5zoGARm
AuvyNhpmvhpCuNHQeQx+FUl9/NFFgq72sWFQ4EI3ZjJC9BI738EZiKwkcgXRHSGhrndyG9MltXhQ
4BILRgpB7tC8xyDMF9vXfsUVGtT7BJNrAHXF5opGkyKoHqa48I9V2VRRJlqInFgilRetSBGARRyR
jakUFpOW6tPMfcG0NehnAyHSsfJfYCl1wqDQxmyZ7Z6SzCn3W9i5b55I2PV0dZY4jStYvbk/K7a8
HiBA1g8eADn24LQI+BGaC1rOV7GedkHfsfH5rkTAtPIAZtGO+xS8g3UIzH9/bIHm//ILxJ6M+jh9
rf8B7ntHBvDXeQnZE1CADhNGhXm+Ydzh2LKGnMPZy8vhiRRxrS6FAHShqnzKm+k9laiA8cMhHZhS
eIpTjwfO5E4R+JspJW7HaLzyFZXUJyRtDdpxNtWhhD4eF4fAmRSYHxM5IsYR2VDAQIHl7VEN8SVe
skGesff8xDnX08/9l1yMTAYg0H8EZda5xvClSo48++19GQpI1N3Ej5zvL+z13vB69M4kwvKWHxNe
T72HOxpb2+1Ez4Xfot7Gb5YIxbmRfdRGfI1ZtlYTPONmZ2xa5+7Zekjy5RcXAb8tf2/S/DojfJOz
jadW0c3N8dTk5Tsnnw+kwMU1TzoXN9d4eV09i/PgIx2ZVvZj1QV8d44uPVoq7YjygxqIpi2yA/9a
MMTWEHvqDeVfP6qypuV6kfLK2XD59lh9D9Hcc9faCThxEvbiyk1zMYQRSKwL3PzjH9y537AmpqdI
gUiGpZenSVbQZhzJlutfHK36McbWT/OIBMDvmNz5XHXHi5s3cGkjo9eWmba7NWo2AZ8XF0TCxPtu
EhcaeUiTZqTaiHgdDxwULw0m4o2W7WWvsbJbw8JiPEL9rOsPYz/SmlIEn/oUzzVx0fA0J0m5zPn6
pBoHPs7QsNWNriVAwcHmv079grOrHENH7nHUTYRxFQZxVo/0z47DuA9ihOK6SRjKKsmFaSI+whGl
vb8aCQtk3jh5MzNLByJloc1Q4hxwn+cOLomj/R7IOy8g7q3KUeCCar9yaTx4JlsNHN7jPWgMucBG
Z1H93yLdUp9Nq8iDDsB026KleIdUIFigv3bFYtzyiAvFs9gi96vkx1nsKVP8bK7ATNhFVACXce4D
00sEfK3l5lI1OHs85tJ7xMdbfpZ9aGGv2zyTV8JhHBmygAW+Fes/jXCBGgczpP5uYFhJopveG0yc
Z3D67TsZRMMVYZNoWvgDtZ6SqhUvtNj7f+t1RrAttLwx2ZfO2QrIN8TB8f8w03Q9D5ysrr+jMwCV
/lQ3G32N383kS8cyV5h+bxHDyaxCB80uhV/Z8FNHHwDlQI0kIQqV4+v21VNv5n1t2WHFYchEbDCt
fa0fFMBc0ATryEytr7tqTKH3Ib8R8yUxYHD5AuKlVwIfJA4oxCTQh4jxhqZ9WVfnDeIdf2tlo9mm
hJuHit3lsu7Qjttlu47ylQY8/e7uXgnx3OnaxSVTerpGJw6iCD2Z7CBvF95CyYtdmO3wxStWr+XP
4wGQ4/Tz6N6sYGqYBThf5IdCCHikLQz2JAd00IM656oCDiRg5iffNO262deXEyQENVC1Rx0hnNQL
xes3+zeU2TAz6Nr/qrJIG/F3Xpg3XYVQj6wPRbWmcIPhQ23R4h/qIuYO8v/RAqGHCRfr4gninHMX
YNK20iCH/IUeSvAFNOKAvxsg/io1x86sT/dQKufEQ0PUBa0bBG3r445V/Sh7d7QojjamhowskZRr
CDxevvzarqh0oI0/nZKeYChnX8v5HU1qXmQJG4ByzkXyxd/EIxKGu17xHJANzOuEyRiVschfj5hN
tFJWpY/q2KOwUeldsxSLNAbJJAbbNCgPxMyiQ2z7ZLXVpx9ktFViLgGV2rnKe0l5sL6Bkby6g7Ym
WcJSA3TYDMzD0NuaRv1zTTGkOHOm15HWWcvhhxhZ3FC4A61kDYONxFZ2N2P8p7Vg1pNSkZ+4yCKL
xkMAWw+Pf9AGXf/7kOSRCcYqjvb1cJmsHOPZqcT04KWeSiO0yQx7/U1YhfdAlIJ67rtPoCWf11UB
5x3eJzQT5b1bbnJpslzrpYqKd03b6bELDIQrb8TjR6G6G+13cIhyGSZe8HqPoqS0tz5EcUik6F4Z
etZSKKi3pyuB9s7Ff9OFTepqZ25ozoFMJVMy6qG33km7HN0FRLWZMYflPhwfeVRL7/w4Fs8CnsNO
ACgWL+WnD+nJFubQXX0FlHX7jt/jIJXFNdy0FBEyZhkBxSFFs5p5FLiY4n7VDp8D5F4uooVCG4Id
379rouiZNn0DO44MaMgp8sp3nDaBEQqq0UIbU7fgl1pB+qdNsjmwYwm8QyW7yEToriYYFTo9lXx4
vss95kd2/uaHTDIrm71h+/qtWFa2hG04acdcbaPKr6T/lmqhKLH/kymUEsKPCw5lM5yhdV6O4/RS
oN9Y2m6TreCXtpxaVRSX14fz9TCt3KTohzVEMKOnMC6UqH0PICBxww/VZ/tKHjNMZ3TCXACEf6xF
JjZ/3p3ILyZTKDjN/BIrwWWr+FLRJuNml972Ef/71ZU5nVtVgGP44kYr0bGZr8qVv6RCFgh5Ekld
spGmjksNsz1f4b9/OA6OUGUHq8cQ+ZdasDCUJZnyBZuleX3i7TyhhODSjt+UZApG4KzHe6+ESPRZ
NCNXIp+E5cbHwy48OR0nuNhY4/lLNWZtJOtzHsmnYeKbEytyNqxLbvQ4K7NnJnBMSYcl362otwYV
hS3TBdAnxMRI86NtnXwQNuy+er8JTJUJmnnnMJXp532J/s8XHEdn6S1ZjvSb5hxtePgL2ajt9yME
5Bjkaf5U7vnI4Qga/NSScnyMoiW5GtlpQxrRRAeKgcwwVSjjtSBlPVIrZOGjbhLybtYPfs8dolcW
LhwjLPUSovSrUiErWRvSYZXRAKZxjieR9NklgN/RAUzY/wIPmB5fzw7Vz24dpWKYjcSWFGK/b0so
GylfCfeGmAJ8lro233mkZI41EDWCxOqZlKOh+2HIDNrs062yX1N/Z1A9abPeFMc9fdJhNCpMSu9u
XL7NYlAC0Ou0+BBIFy4QEk+OAOTRwOUoZHwsaudJb+U9lq8Tk/v2TUOZqBuTMuP+Des/tUBQ68Bx
/ZOMwM/s7FTkNpDZ4V8Qqf8IWq8dYCy7fuLTij4e00uTRYyRndYH04RZA4Uq95jZKx5Ciz5QXMCT
r2Eqcff2VYMGNKn1Prw6vMRlZQFm8NYDIFshC8RMw91L18zcq0ceOKCFwNG2j9GZtIzBK4mR0Kza
PA1ueKkohlLgvXwBOsdm7cVZ8Yku5HyoqUUCPKPmfTXkA5uK6Oy27BwuZ+zcuTpWO/TorgG0Yc+O
gWqYggTusMDIBnlgklpKQ2CRbkY7cciKV02/ZyhTBodf2TcBS6sjuV9nKVRQIxPIF+w5vDuo1kQJ
YpmqC2zbud3IzR0d08LGHkoxS+TfnNeiRa73aZ9wgrry0mzHA95lanVuCqjqnrLKakWuLCYHzQPc
cPx6d4E6sJ4ixhVEnEPHHHGlLjxeJe+ZL2bjAAQaACvGWKs4AAQJTrUw/oiYUed7+d8CCSUAaih5
IhoZWWl2bkpWa7rXk8laf2GvV/N4DXCWRRCRaLPGqIqagbEEqKgLPFvRNoCAAB3GWjcSsC2ODfTY
5p/xGJhS7NI1Yr4E4KbN6UgMRFZqMvHLyRb7M+gtUaDZd4quFnh2ysgOuqoKtFndiGsBalh0VCoI
fzPIYsxRQ0ZfY4sneCY13X8r1UgDi4QFQT1erE58kCWGw/FYylVKiimwbQzuQnOrSESlc/35WkJ+
XClNl8L3k1QqcNKJOcaNZY1ZS8aDB1xhLFvvQW7UKDQ1VGa/DNu6LIAy338P9twf8xYkEYX6CI8D
Ln25S9s8WBmKPv05+OaJtF8yYyZxaiSLDsqBnwxrN2qTPocceJiakE2sInl9CFSGGaVL6KiT1bhD
Xuqc9th4TCSXyG1YXAcit28rgMvn33GVCfeAjLCGIlH8AYLPeXFR42hpgsAOgGexQlmDvSjIh0Oa
SCzb4L5fBl7x02LQw3zW/rH1CRkAicGk6gyZH6qRDqioJnQB1dmlSOffhwgIYHaV5jFzSYG08BJY
EmarjrlckqPE9//75DozdKhLbTRVugwjAVR0TyWe98r1JLW1wzPqHl8cKaKeKZ9MhGDhBfg54O4J
+J6dp1UgcGI55W7+cWeW09eOlQ5h2w15kL8jAH6+6p46c/M+itZUlWOC1nThj67VnrClGrsSa0jy
zg8zS9AmQgf4fhkL53PNTc9UyuW9RMq+0gk9MjTa4t6CYdXAyTeyUpPk8tcjNTQteZY9rx7gY51c
KE15jDaiVePmSpgzE6qF/uylbT+XVSbWaQvGdu42CnzjI0VpHKw0dS5qack3qZP9OYlzBqkRrTfK
+ubzEKk4IQc5Z3Nm9yfcWql0SXdQLqdUhwIZij3vlCzr/vt7hi1Bi22Hh54e/LYEVjdbyhEtZ56+
C4sSH0TUY6c/B1XC1JvhVnxwe7CTH4AbuEcJVP/1ArosThXeT4OSB/HQR+nYV6SGl6/LAHA11RUV
6TAkGVhoLmBlv237cqlLEasA/8qPax10U7FlXdp0rBs9z7sgBshIP24QGIyiGdDgadrJtWst50ji
flsvt1nSi2sgp8+b41tb7iIM5jmgzp4IVuz5C2GaseBYa4lPEOQF/ZrLLpEwQcCpt2Y8Bj6XOOip
CkICOzJvfMRwm61HFnVew5c6VcT9HNRjZeqA1LbrSmPyT6KC//HrU9dFtsh5h+P29beQvYeNXCKT
jeL8VgzPO+4/ztFz6u5oRn1Wql3cJQouXA4yUt2IjTnySMwCd8NSsBr8RH05Fb0XIdcxmgUvYZmm
GU88jU1xUCZMSR4G6ouhsXdpgt0Rv2mvaHlFNi1czyvrW/nPfnZdQ+rb9OilaqOqZapa587FDzMl
RBKYd9SxmTsf5fECw6d3JAOW+va5Zo3NAPAtskj/quINfGM4rlL6GCA48SHBitn/qjaA9y2491Zu
4P/5V10e8Do2jjHS8IAs4ZjYmHVgtxSmaw8JhIfqFjjRDoaDdN+0708Al6XWX6Q0L1yDUXfaAhI9
xWE0QpCiaCnDeEquHLVtogOzl5DtJyo6dVqxl0fwlZJybWRhqsZHzWApC9X2ha7gU63/R6lAPYYk
Lz+ZwJmOT+ynr6qLstmzkAEAhsYmMeaTy/XWulRyAGb75XFqQ4M9HM9cnhiTS6nVI6XpCCVrwsHo
ufSbGtTNvRBgHJ35Wv1YrfFEQq/uaGdaSGTo9pFdrhASpmnzGQ+sxnglA29K98Psu5BH2jwP+afP
7QIaznCwPqg+OhhuYiZPfv8wypM6xMR/zf8dHXDAgDlx0thKrDRuYpAvEjQpRD4n8nSCOYaE2FH2
rXgtVakIcpHfkdROe49Re0+YS900CkZWLKBUVWwZoQ50s/FeZ3+GftTvg9tYJiy0apd//yvppZYX
iIgu4k7RBCC6ZRmrnnlqg66Ms+rkak0xQdPUo61D/Oo+htwpxvJ4sATDeAE72VQhMotEVR1WFm8v
ZwUiRJvuPBTLYw5d+1p48iStrHIhnT9D+OZ3JRuuZL04CfPvejZ1QjM5tX79nJP3SMmGfhpU++Zq
t/YRzj5kVG/fv5mSGR3Lw0N1oeyjKfx95GB9j3lEQ7+tor+uJLj8y2wheZa7JcFyYypQA+j9ugKx
ahCB5o67zv9OBTni6Tx6RwZFXRE+AlX0oiNwoNGvS9A447nQNL7i88JvjP5lJqF1nTnpziy/rEWr
b4zuBlNeT2J/DcWTeftfOLC+Srs9rHWT8eUQEIC8w8kLgwFq5AS9vlD4ucHuxJdtdA4YANivRUZA
G1UzPe+03OgxXeyn1x/qBWR9HjGzlZtCdGN0wMCtoQbudYVRDMBRVt70esWkj5yk+4bemc4crag9
EGv/cX6j5IytIJ9ypaoNsMsv+8/edDIvL6oUkDZgW0BEQU1CUlwFoSRyDI0pxDMYzMmFLZbIfWKd
SspwFU99Gpqb/GYCFv+4aSsXoRtgEIAFlRg/+OOtRFi3ncIjD5N5hjUQ2BGbluaLOvhKg37giZEK
/VqQu8gJqDqiHEc+bIUYBJ9vTnEJqh19TrljxX05v1XJepGpuew2VFlKnqpVgqQgteXBimMrO3ix
jM5JEQOe7KNmidOXNP68CuLrvLN5N2iVkf8fwL75zauyxIkh4CIuFLrGw7HFd3DPchZUWSrBqypV
xsG54uiY6U8JvkTcCRZknJOPsrtTzXH6pF5A3YC9RsQjf88V2AaX343eYf0l514QtrISmdjuLIfD
RR3PtWSRY8I0OYIxLr9saENdFmq9YmJoAWwuINCwTLCbe/3ETEmH1ysaZryDka/TaXz3Exfpv3M9
IH16HhQM+qCaizG7CEpvmxDpYSM2HlwgwdLz9x/Y3Eips9wpCczRZ3Q/VJCQknoP3ww60vuhHZdN
GDP7oZFeZ53LtlmIq/iNs8kgFzc6LhOu883jufDfq6W8RuADK4JEHopM4j+iXjYXMliWqBuGrJSR
cIKu0i7C01yf0lxQvGCMCPwDmYECW0sD9mhhewqcPmoy7N+gGfi9Xbs404dlUxsYusw7s+vFgSVU
pNGk0qsxmOisdBkY6JoG3JlUwxRJztEbPLCqEy19Cx2tmFMK0JSP+l12ju7mvPiPDkkQc5g9fWE9
L43x7yrgqmnpg/HG8KWrPpgDLvCoCqDeNbpTkvio8mASWjflNfhbFKicXhg2XkuCmQV1E/sIeKJJ
odNoPVS3N3bvzpymECOwp8nMxwiuaqhbk3iAIaDSV1qC5VkxmNywhaRHg6WoYi9qylaAwQGl6P4T
lPti4M8ElhXBozkWg7XDDKYmdgYqaGlGeSdyyXIq14Jz63qEf61YA11CSlocRf9jZMaXaBrfzFkH
rYDkwE7skLS6h2KVPwDYgMh3iuL8IuV6W7tLzkVT3F1gATrJLcVxtMEXqRcITn/1MClE6h/tx6JW
moDYWbaqh5sYVtVdl6GGhgZQybBBaRFRNW3Y40pijK9hDiRxpzOcdf3so+kvqfMrL63ticgPNvHi
EVBfEC3iGo4LAchNl38S1FCtIhOrsPvNCZ0Vlf3AKx22PZgwRIc/rE9OZ4XcrqBaHd1EwxiRcxpM
f+VxUEaPrnrm6euw9/BHR1jkSGDvH5Wi3mtfKav17MJ+dHkGeDW5PJixuutjGNfzSBKyRJiBMrFA
KrcxM5uLRiocXJcD9r89fMMkVYTEjjG0K6U4uTXQC0enzBmBZskU6qCnHCcfl8vi9VdiHRJvC4Zp
4oPb8/GxKeas56mrQtMq3tR10SL4uacIQHAOl/x0gj7cDY7z1trD0Im6A4qcstvJgb4lnk5sSeYL
WoeRv7vaFYqZcb1B6BqsGJwOq9V+YInA0/tS0N9+qTanpgQbAUrzuJk25ZaYutq5fXcxkTUMyJyr
h7/1QO7N7+ZN6ybt3fdt6KQ5eeUQomm43kWBmJjRjDi7WH1S1aZi0uvPmjEre8krbhHHuvga+FCd
g1DlL8kz4jB9O4EGTFK7TWPwCL88H7g5IEIzCBKQXXetE2p+MjbzbqrKvvWnqPLQtqiw15+KgTkq
olVxh8LhZY/icZb5IsEvQuC5RHZe/Zo9N1nL9ay3luFSKSum2Qf9OhfqhfnlxZiosQSgHdDt7eq8
c5ellovfSQDHMXId03wL7gKCDpv8j2G0D1PtcU8J0aRwUL/oSeawRUL7qh7MJS72pdiAQe9wSSaJ
Ztp50wslFEO+bldmXLzOSUbUUNum8DPco11lFjNvrBf9clFZSWYJBSJi53WK9bjn3F9Z9kpOsEtT
aUKtmAUinDVITorJz9ziuY+LSr+38GsM33AlMJzxWiQgvNA6n4jI5i4GtItK0sJTQ9sgv9Sg/njE
mRxUsEYKbBSiK+Dt8TWj4k7dZ+QXGiTosjmtjje8Q2VnBDOlp5Ii3BOKLN+JTpb28YLUpAa12N+h
Xp3B1QxC0LPIvq0ERlz4GBsuU9mU3SBaMUGOKv0brwidwiQuGUAjaMe1TB+5Y6RvHHy2B9rtTXIN
797ty1qD9stM/C5VcJ7BngyD6+Ha94zrDdMMPPosBoBPRFeLaXyJ2rZ2xiqmRZKtYM3Xh9MVZCzN
FiPOhEfTsumdBDVODsrNhd6ubmCvL1WdJIWZCwCJglYEhE+FLJVPYtlgxVi5aam4PPdmzRxXp6bV
ERfazKKgyEShX0r23njthDCmdhn9cYKrVy5yJBV8gpLcb7ySmxsvHDKUlVgeKR7pk4oVUPKjtDFy
01CFMCELa6HsNbxder1gv2bmYkT1QozIrgYtCzO4ZyYn43y+N0mfgTv2An/cqFeciDlLi2lPzhNS
2riw9k0VjS/C7fyrYLvwHNfE2btx6/K3AwuHqFhkXcw/hawqcyjWDDmf89qOvArA3ihC+vGp6vRd
OpKVbHFmjx/hrfUct7jpLgz9Dz6tVu9dXzXPfZa2fF3xiVFzYfXn04HuUhJUO6ge2I9QzU2Mcpgg
KIIYH5mFBBfP1MSVwNKrDq1eT4TFp+654092rpLqbUJyFlTdS3ipqJ2GWx46Kgaoe3qdU7H0wMWd
XHg7c5mDlE9/x+VVt1OYP7FbKb5mu+s3A1coSWZEpZbX0SyUVHIkorJa0qqpo08CIMcTycsAiHyV
poLXwOh4EDJWlFdgVRnR4gM4TZkZCAo5Y5W4I70n4kZiBtJJPI75Kcd7wOByV0doCtpWownRWIwM
OOGzrwBbBj/c5VcmMiRbpE568bcaVL18+YY83EncxCMG0QJtX3mxTlT3EqDnunqL2XCpF8bj2K2F
sGGj2331GUohKmEYv5lduE/X1vhfEBvkEfd8w8UOnfaPJXcVJzTlQINJHzCkmXnlZIAcw8zTx5J0
jsxFbTISodaTSTTorh27sYXEsuoVC6fDvO0ld2WXipm35RPcGjTzMmVyaeuYLKkkmFQmI118qqjX
yijJVvzCxeVYqZ8xxbfjwrdJfXkVELIHS760knj7MwT+kH0veR/ySxadFkKP92y+Aj3jWitWewEs
VgQLdmBXL9OGfc8kSxtNaFjCFklz7uLEQo6prIEM5KYaNV1WRiqNIV1j4vxnB4mo8A64PWgfE3C8
i0VCYQzCzdFuH5v8g1GmaafmN3SCcHfUVTQ4pTDNpF1jD6KyP5VQhYVnBPJNgUGqgIRd3HUVKnyy
TnQjYn6btAheZJNlnId9Jb6tvlDRzRBhY4IDhTf8ybZSLVcbzWdOJyyQAkLyV1UpsTbVb2jYUD1Q
gJt39H0WUmHbis+kV9PrG6FqOV2722MbgZThwA9mOpkpc5Z62RRFRo6kSAHnwRZWgMercL45hKCO
9uptzZdsjpBnltk0liGndI/WnPEnW6AqY2lKKbsdyenQKURkVMGPurotDRsH0u/4oaYxvW7hIDwF
CFNM+h8eNWXc4nkrA2ttNYhCvo+hKJAihb9RuPwHYERW3qiQAXioeYK3S0EqljUaUVzglA8+Jpqv
K8zMdp7LPuSTR+62GeB4vamTg2hqZgLxh/mcPI5g6tMLOV8HlC4nDtHEyQ3+Y87zW2A38hcAeIWF
rjVvjD9Fzb669BpHlK3H02P+ERu5Rr5c/eIi64+HCpx9HQvng9m4CL3N0mx+xTfONAK+1SY2A9bY
9ecWmd9L4mt6eBujQlKmFrn1Nmngi6mpYCriFzbIJXBPUx7etiYQmXEK4LBNVEtIXVWvLQR3Dn1w
rEHh2t48xUhVHqrdJ6dmItGnfreHIB5r9bVnTIKID7d5tz6rhXvNciL1XvsgeiOqkTTF3jLuLqsm
n1LYpIBw90MIg7aaAZHcFU2tuRzhI7hhh3VSbPSBMtixhjobIYBY1H/3kYjQo6E8HkXwaLPNH1pu
0GKqFpGKSrBV0f1OWeLQ9JHyZNabseHxldZd3BCt8dnqnQ3Q+eHYYwMYAqNHpIQPIiZk/nVJv8xN
oM0vruBhAKyRyDjXFnOYluUlAPCKFQAsLRx0LwBvy8TjPPPLEA0WKs0KZS+2ZiR0Uoy7HyMnZaUl
LubyGzu1VmLAv8CeMSwn+AteI/pZODL6Ua8nlKXMEyN3NFhZGCjKgMqi2unSqBCQkgNKKPaIeggW
GG+0Hy7UQn8sYRzkM9s2bgvE1Frsh20c+FW0PJM/QmPAA9b92GLLk3OhhemAe0pToA7aSmQ2WoyV
7RbXzhNU74ymXZxiXSUA9Rl52MySR4hyRq7a7DZYdfMNXHR/lEsz0iJdySy14eC2AUWfv492e7Qg
YOnRZjibJNCTZsfUr4HRQ6nFtW2kqjePHhu5UVTLESRWJMuvFW3+uXefEZnjndEmXouy28RI33hN
AK7gKfmbV887SJ2Qpz9xYVx9exrDKlSg+yEfiPEMRwke32QWSi0bUb78DI1wNX2yHghBT1CDS5fb
g1Fi7ZuGvDgzAmG3jSmGUkZX8fgjqJghqOduyJyTKHCRAWaDnp8wJznHTvlHiwbLhE19AmpOU4cF
J4et7/OisoZB2fhrakQYkM0W7ourWre+Y8/beiSzcKFqD1MrSUzbHHaS7SQu+offZDL6NT5/r44R
V8VoBtmFBDsVHnQWPpBHUZaT1Wewy51i0dYY/qPr8Tg+np9I/voKsjapTaexsoxOSZrOIxfV2acn
//zSVy8mFftrErjM7xASwW4o6takXkG31HXQkwURo14M6S2MsX9YJuX548FTBKTSfwJFL5gGgIU8
4nxEtUjmgxB+1kFGUVB+fnsEQfjRgRpo7OD49mE7k5SWIWhJOLNJcbSQBqWiEof0RDRUZ83z7g6U
rqpFURPHa5LPjvgoLY+q7ogZRd9pzimrNYTgTvBaKubgMaMRx3epmHA8q8WB/yakTIWwOkQQAciS
w6+bp9zB95KJKzYARPQdgQbmItdRj1PNA++2R3twXycTu9c0B4ltKrGDV+FneunCmJ4s/i7bFVwi
ZsxYSFDr8bwJLxXYjJhDm+fu/PGs0t553zcaScCPuLO+42iHBLWBFUIT1hdOuhs26vkViqWKhSaU
JuoImn1j6GFjpulNaVghCJJ64opEXu3KRzqzNcDGXSzwf7zophVueY5OjwHMH5ih5STyXM6+QNp/
RM6SUNm31K94ZCKAsJ8nBUzhjDh5UkQvTltqh482slqnki8zmHSSV47faxuA0HvECgIfaddPGsY4
zsj2kbxo+Jey3igV98jzLDeZTKruKyR7SIcCxtTi0CQTNIV8KKOXyiEjpdI/W1CT7I0XF9qMk1bO
pnnj9SigAIryZ5N7J5oaEQ7KvL6tny+Kwr4vJt8nZb6rjnMLfTdZUJQ9QtpUbDUk3yj4i6o+hxCa
84zhjPJxUt3UWFyPReHuRd7AdYuY4dN7yXeebjqZUfirh5T14Y5yC5J5EG/iGbGFgNoiG7KaqlH3
Oi0cp8yDUoqcYVlRGiYzb7poTBkrE6lM2zu6KLYR8AtON0ictu+92YNZeLcAmeCRyRGYnbkiyOUt
OltMOZbgxtiFHpKCBIObFVDH1ANx/HaElVDHjrvkD5gyS1A34rAPNh/d/SzvC3boezDl1R55RC7C
Ji+axSDsXgvRsNtDrJg79VTZD23j+F2eYpoS1RRv9FPdr7WApWOwY1DbPVij1POPylLX/lKqmsqx
7tR7lRqEOnxsq9MGdZoh5G+Et8YoPSSMaSzu9XO+t4N0V9lyp8532m7x30D5tKIIh+h2UTeNnwhp
h2WlBUx5z562cHxAKKr84DgYDk9a8F7gEDzspYQHJ1Yzh6b4DUrYlbyMeulEt5Nz4xKkLfNYi1Mz
aViKZfKwWj2PmihaqQtJS9yRsM3e08Wjk0v3lCcgCTjp51sAFqNo9QfSTvvU9VcHAsbHe0b7Gvdn
WW+kQimw20r4S8EOAj3Cz9LvvW6WlAvVA8kf+O4yyYEZBsN1Y0ng11AH6xEIAAzZlIB/+JB5s7Ke
jM3r4qtB/hDWaCEuBVdnD9vcgxFEzvpavBXrcKBNjbxtAtchOI2Hc9+MybX02jcm8g7rjg4cWzIs
KZ4Vd0Vh/7Zer0RKlv63ku+4hsvDfeNDro6+g/YcfyZMMmh2DUfg6juLiQnS7iw+OodQyu2yrF/R
bALIwoIvoKG7DG4I/H3nD8JrdKqQgmBmq/qLXPnmww+Y+wQ4PHE/gecH0DxSoAwCCDQoVMW1PL7H
+1hlHyP7MYpXcF4t8LocTZTY2mLa4JF+UA+2OmxkS0JgvJYP23bQBO6c87WYE8wybgRkM0AHAlJ7
0icn9+Z41h4kYt0WXACQWNuKTsHgM6DE6odLoPjWTd3i0dhBkv6gdF2nbOgnVi8jOMlfc03Awh5M
OFw0OLHJTqh2ZPyzXFvMF6+9mQQvT8iRrgwBRKKLfppiU3MmfXuaHTvvNp5QSaZvEjiOEqsZhU5p
KrGJEKqLTIwFaO6GLRkf/ETr/fIwc79aJ8Rk80DT83LTCCs/+dh3zrsmkikPxIOkklUvKY3lpxk0
65Lh190usKbdwr0oolJLqLnTCDmwyTXVs/0vR21ncT8b0gx0xVHH5Sbobe+lfUgVkR7kXDKGRdFC
B/9ybBBhrVrLiAmFTHrjnfLd6VBW4Cc8I2oNCZamNT8SF/3RLRhtkg0cvYoHFvTwr/tD1bnNJP/M
1Bpljy2r7X9LBExzppT1yxNmy4re5t/lwDKIALSGZR76/3QrkB9jsRl/DyjFkkGfHSu6ET69bF1P
92MIiYvb/+j0htDHLKY3lAzCHMHYQeOBkmF1aUKlBcvg9gvbI2rTyn04zto6IY35qAlNR3Iqh/p3
Vbo72pwjt6u+MoPQClVLpqm132+mL89qFFKiqLkoVwGTO+u/9nnqVPIjbGNpzdpzKi356uWhfFtJ
OWqA15M2Z4WCvF19FH/IObAB9sQI4xlTE73lAXoTgI8zhkSl4VPMmDZAm0uw0Sy6VVCXDTqE+cky
T7834eSwPv4nB/45qFuGNywrwIoCCj85msbnjy9rCk3FtAy34GbUQhPpIwo7N4BEhnRXuFQWKZUI
jTt+OqRSkjdNvSTvzVSeRrBmtJELQHMFbR5SmUnLasQU0fObpDpj93PDlOUBr3g9GUzbVBLaTEol
wOF++w/1lgOMSDJ4lJvBz3uX0eA/vqjB7oA/o822u9lW57LGQSQbjipvKO4fhmN01JyCiqihmKV6
OpBz3QoBNHwd3ffChfa0xXZo1EUaUl4wBpwCcdct7tJth5nmeNmKb7DgTFWzTit8zcugh6GSsfht
dDDYDrVnvbrjMotFgl8T7L5rwZpGdvAPyj+yrmnQU+oIeUdd+JPDvLNJjtSxloBXtkQnWHNrx/uf
SPv+s6PRa1A5yRSjHl5msQlq0tdvsPpNps7sYrRA9k0Sd3LOPcX9O/lCSgIfuFCzbn2i4eNUze+k
EuQFBA51Eyn53tbDHovx260lBLA9s8RkjaSEHYo7W8M3tiazYSdwRCYJfAU+R88cyT4RsTFobU8h
RDe3CsjqwcfNeiw+r6OwRG7A34/dAfT2v4lLqe61eL/MrrcIyHqP8uf5wKgqfnOY3szrQT2nks8A
Kc7rxDNr9V2R0fWAyKjFU8RRpUh7Idzolw3Rm9FAGGn8bA1oupgsYjACDK0MzeTHUZMEr25dh23R
Gz8JO4s2aYa1KJOfnxtbGHyHF4HKOSvQOXFzuETgIlYvz60SBn+jJMIP9piQiVPnj+oCdgkfv1c3
Qm0I4kEW1Syspxz1ePd25+raaH+UG003fxmzcA/hiIHYtoywx7/Jg+zVH9I1bxpl02mjLbq62xcA
PzHP1Nor2eADg67exBDhPfeA2TJv0qbQkFXgUj7Ah6kdVplG2p2udwL+W5u7twPX+BWRkS9FtftM
lzJNT47e28fU9/S7jXa8nGPxfnqj3nklVLq6dXrSRtgoaNvHsWg+Tc0vqQ3h9LdbOEV03g6sZfoO
HUbkKVYV1rJpSYXPvlJtcEO/oxHrZG/TH9oPcJUvCO+P7uXEgSW1SzfTlXg48o90aK5Oec/Y4B1T
vLE8Vs+EvcSzwhf500FdRJFVR/MZ0oc4rYvX+KKYpUpAqCR9uPph/RSiBxo4E/+gqLICxi7j2Xl+
Qrste1vngSX1mq4TchhaXsfEJkh5w3wqgMOgkaMsBSD40Zrkqh+zXclesUsD2+mdCjS50wZ/lOju
7FYP2UP5nXiDi+/5yaa/poLwKlhQEp5YdAyI7ceOP+G+pJES40BJWNHSe7oyO5e3B+mqCLx+tiZj
bK1GQByW3jPleRN3s0uoeb6ju9lkom9xsToTMmItmagFN9Qqk5ZU/8DYaYNEBryZKeXXHRyf0lHv
nbymc2+OLjzdUZpvdqmGTNSqRlfC2iiYvwTvRlek2/Ru3to8DUYJw0YRqJXKgqEaIbDXeMhRYJNO
gL4k5zAM/nUtufJLe8DGkOaBk7e8ZZhIv1JSnYscN6HwSz66/YDTBhmiokzFfDOpLyG6PX3jMEGr
diGgWO/ziUwu5me4R4x0nY0x0bY8jJbrpORULIxL25e2/156U5JGlXuIy1mHRPXlXJX5hH8qPe3b
248krcwAIkvlWO6C2CAYqHuuW+bBJlm/YcO5xs37EZSOwp/plic5vxVlYcoIpF+E+HVPEQfCu4wu
tdJgLiTOZ4VVHUajN0Lxqyw3zXwUzAb+jLpqBCXu4W8h3Lc875p71JK8KFYggoewdVink6q0v1S1
PV05FY9fvAHacRN8TysDUHP5flg+Uui9dVNCo07t7JAIqCKG774W3ucLyphgSWAE6Qp80X/8J7zJ
DldnDAo7x99Ez4WUGyE/ECBvxkdhJEzhFO0wPMdEfZBuAmfq0t4Ja4Nn49ELgk0F0xraQaNchEz4
vXGcv+c7gZljwVlQHFTmZY4EKOhIYpuelf98kPefpGLK1Cog+tCJPgFLy3je146lDjStRRuZpygz
QCynfhxHQD/C99r7bHRLXW2qblLarfkwCmIpfamgxxYQa0URZrOaLXk91Q68/T+smhbX84nJSrCr
VqKeHC+wmju3wmDsfc+ElT1qtqyhvHP6ZMqBdkCfMIA+VQMOGYym/dRlcDMLDkU0g/dawhja4rrO
3nntbUY+mUVKtrGF7O3gsXJOWZb0+eDsaDccN8bTbrr0PTmV25oyPPBjTUOqLaXwK+eOJw1EIYM8
6ys7mxjw4HZ+SPbvvLY28dVgV1RrfczDEWcyLfVW7XyazWi94baMwgsP08YLhaY57Ugjf0YNwGnQ
7uqvEexFPpKPoHuEkfD04Q4M+Sxby2yjUinBw0kPIqMZ3rqTqnzQ/Tm7h6CLY3khcSQQJfC+ZP6H
YMNy6N3jDd3Tps1W1HtYy81yy0xTP18r4DyQPkf59MfwuGJ4ZircbLxgSxV87kFYTI2OQlF+83r1
+LPH+b7tZvHR9jtfuKMquGUp2pahVsKNTZGlm9oY80qtZ6P4rHgEXmd3WxNLKcat8TwOy7ZtycQI
yIhCZ1QLH3l8S/IsZDTD0XkomcBkMv+RR/O8x+mbS4gVTmjLZKS0VidkppOzYZ6IJBJDmSeJWs8a
5st7QaXG4u9ryAPC2sUiQI8nTzxCDHuYh+C/jxl/I4SL/9r3uns5R7ROM6VkwdkCVeKKKZxmludC
GZdAtifhXV+fkXz3mYuVG3QiBMTRPKt99CgC7ZLVC6IWTkNin3BesxYtdXtn6eufWYwSRyY4qIs8
fl0b2HiVviKPWfM1BrAKKvFB+01BM1iIovTErRJ+q+LYVxKctVvqoDnsmJotNWakzc9CWJSn4BA2
X6dJVNfXdiaRJit68jGbKDS/rhL6omA36ZAZT3opMCBeEFUb45OgwQ4R9SIGEImAMhJhKXyi1+YM
ZC5pCYtiJItwRJUJPWwdlMzNNpNEBGOibaELvbzUYIsg1JzJCtX338gqKYawBiWY5yB7cz+hqyx0
6HD4I9qXZoN3Gc8uMmQpNu7oMbQz+FZNeGWBcvGSoOkKY8P0Rh2NNo9d+c50LACNVpX4gqIckwXt
rUGcazDg40laJQKuOXXOtpaD0JqmYnp4AX6Oa/23ZVgOzbZBI5NTTmR+X9i0IxvRJiXbYqOp1hAW
ms3Jej1ssFwHBF3wS0RbIKkNVUXvSaJoEc2nr6nS7FZ4iskttztvPy72bMzrgh1wD3S2ECmDL2YT
RnPR+IS/QofjY2gxPi437+mhxLdM8AaM8mxFnae8XNiKzXI54ixjPVIW/4ytUNw98OPGe/z7V3d6
AcVzmz4FX5goOCbu1EdSD95h53u1zyqs0oEFrWUbLiOdiRmXvoCyqX+Q/sl6O+H1mRU7lxoAiKp7
yg/rWmWWJepdQtBqMabL5Q+VFvfNUn2ieLO18YhoXBAIQk/tZo+4J4lm0SWqivOg1kb7VXRpdtrT
sQPe3+NyR6xReKoTPGkssbTLM9gvNM11wphc4qT6YVk/zJSAHEmxbZVtStLzQBN/1Y4bDnutqUiX
L3NAJoNGVm1iiUzFnevPlKg/8rwZUiIYfgszCl4Lc2dELFTCzc+OlX5b77nnd/Z5BEBE5X7HQJkh
8CWStZRyP60sMR7XDnXejgbKz45OhXuYBDDeLCqszXYaF+Rj4idwuyACnO5EhI76gAOoK8iBI9r0
OZ+lXA4MMZrSndYfHR70I1YmXR4vewX2Y87o8SX3NpXBfsrM9ZIFc8HzXhdoc3bzjEaaPnRcIpV3
fxzOBFczKCSHT3YDYGc7h8G1NyAm64lE0Rx/zWLIoc8nItiAmW2PWiPgYJ6SysEmsfIlXyTxQT91
VljCQnSUmjaPXewuIr85z0hGev5EVMpgwBqRp7ftiVhlAcuIM78Epy44W5UyXAE00fzgLnIg3wt4
kguXgAOJBJ8KlTNtxTbPhtucEdD2PrFBg/MFY+WGPEg19SFlLo5QSNerarB0XcT+S8ACj4NUq+QF
UQgGnPZixvKyGA6k5qHYL7l1QUf6fmY+RhJUowMqtwXYvBFyAES4i7Do3TJEVgNIZfRQiHIYHbNv
nfuDM0UyoCORB46cgo/0G85yE3+LoaSLqzvqwou2RCCkR3Ft2Z/1zMxZpwmUq5OaqxAJv5SBPvNr
QyqcxKKQ8Dv3HSq+DFqZ3TnNNNWx71F4d5CmX09qno5psWVXJk39pPTZBEpZ9VwFSmfnYcjI/pyC
mAxygjjP98HA9HoKSiJqPVkTEOpcm69Xob/CLB6mFhHmtDmUCH7B1wlS/fnOwd1w+z3kmm4UmIS+
R4nx6M/xP4pVo0kwkdoS3v00AnLzHeLh/End9Bp7z6JuY2hfiu2hkdPua76hQq3dZfjMuw0xXUa7
4o1mYhfargVYc+7+NKIQyRqC06/ajVXToDPHmDdGWQpz4aM+n4IJvVHeuWTOTUrZ3Ob2yg6jiW12
q30LdCefgDsOI9MoXBMCddrjcmOu3kLeX0vDxEYY3y/tGZTTI+mtMTXnWQ4eU26RErIoXFpzSbA6
fZUmnhS16dbofZy0ISiqkZ1BReg+pzmEpZExU6IDZb1LJuIECGOFiOikqXRt3gJVfEfSbBBr/SWY
/RTbgBharBmsLv0I2FHCtnwk4j+q56w9IiA6YtQszff8lNa9a2JdlvU9HsqACkFZwZBax/jNZtXb
yDisME4f4wS1Tmj9Kwq4IxdjgD5m8GRmPXsWKK6bIzM5Nz3bamnnvZaosIaQ8L6wXc3kDcYFYkEQ
MHhJAe1Ut0hxuJi1AtR+4sVnSDH9ZDHp2gEtshq1k5RNErbjsP0VQWQfVdWyHS/XnF6nJ312Kf8J
PqHeMZWYJogovImxF7x0w8W7rESkEZqQsr5Auvu+b5PazosHtLzBjDdwGiWphodZfdC29CyASF/n
1KNqsmLxdhkHQ92NkiEucUVuyA3AU5p49b0eOh97rrn2np9GoUQOH43gj7UHfxm8Zw4LZvE3iCbz
sZviVpigyg7DgaeEv3J7PRj2cRj/rODqsHW1q8qL4nQ3Q5D5+uNZRYDShnwo0r/y1y+8h93FRA2X
MmLYim6+DwBvkDMtsVmC2qKd/s7K5TU7o1Cdco0+cofOeeEnnSueUqpYYRFYJyrkx412Js/9dBz2
2BqGAZoeqfZli5BgIeBPutJwtXufzdOj6qF19DTax8XFEgUOrSXeYHmRq68mj5ejqCr7aRFxl1Za
qiHUX+uqa2I3FGo/EU7jayYTIxWPH+HwaXK/uZWOYCaXHDKn6MMwcdAcPB4XYMNB1HD6v1PQGsGY
pJx8RukNrmqLakar84ISmcbc6k3Uh/GBy/h5HLofF5hDOBPY68CxwGizeDYYSZGJPdvVQ43/FxmK
+7Ina9j6aXDYdtpiOfeV6htz/PGP/PjNwF7oWkc183OkcsuBTZyTdjlcwhN+DPs1tFoDVGf05cUm
0Tf6HFInKc679Psxd4/lkm3uKVf5Arj+dsCXmJHfyNiqaz/0ggvM6+maUpADRkFqIdgBf/dfTF+T
hpO5wcH9TWpjdArMgk0xAWhEk/rrfOv5qGvc/PHqIHKocKiQKV1WADtKNQ1krPVOw75SkuTO31Mw
Jc3/a19apBn1/49EfX/5umaqQCizkZ51RhCeOA4igl1R6J+3MUE/GiBm6KRzvat8k1EQXiyUFPaA
k13Zpannfp/xZJw0sEwDhEm0qhWgQEtJ4l89x7pvyEy+SIZp40thriWoqUnPu7wd2RnNzy6+l3mp
n3dQbsgGWvYoLH0l4pEPkKw1kFw3jFkIm0Px496rCstKWSjn2TbIGa9RyI7Iafgb28Vi/QpTMAKw
L17W1StFk5jcbH/WVMam/FZLogusFB0Vk+celEvur9e4VqsQi0QmW1602uF9f0OB6nho9Vu6MJmD
ejTyWFF/W5NdPGUTLCFxQhmMvZTNjr3ezrh4pwOsvrP8/PIDJ4zJkxWsdhV30Tu/Fm1lTmQ4JcPq
UGDH9YmPE88vuLXCgqL///31O+9RADITAZPCvqSMyyanL5ygEw9CS/mepupErgDZ+y2o/wzhSsVa
2ODJeIXnLtWScDqFJ4XYNT54xONmq/9hnrwMExal006HrEa8Kt3erC3/tVNiLePsDcXVwLXDNIFd
eyguSmC0TKcXwDbnvbWZYxIJwJjqsL416KV60bEvGCKkXW5BIiX/FLfoqrEkGu3M/6uHwNpf5cv8
fYHK7w7gYfHIoC3abpMuUjbS5lICdcX2BTaxqqoaqKorX7P9rI3H1qxldsVdBXkI5wai3nyFv0Xs
fYnoI1I0UH10Bt3T3bVHktyPxiaKdh8yO2JqNsXxVykmCChVNrqH1xSBkAR9wOec450J1XIOlS41
N4pQJPhWefYKXtsuC38YbryDWiapid8nLlYsztmoTMjz5OlFpuFc52uzqtxGoLahM6E8s8sIg8ve
6V6U5fr7fi+p8kVEjak9aJ6ToO0La2I0r/Yz+PF+kfumw6nZhi8TRfEfqVqgiCdbg1PhR3Kcs42s
VqSwzGz+dW5lj5s0ovsujiHzLTONCjE0QhaZTsxZu7fOMvnvvXhP2riaR9hPMS+6PSyliP2z0PXz
GM7gHR/udDQqlTSjhgfWTFyqknuCr+v9IzCv/RJRTet9S8+0wyMAjC551QkmZqXP19EdaZUv8UZL
AgFA7tOBxsIA2bilpVDCazfA9k84KxV1HEwU9Xvc7SUnzyqkwQ09iocfj7h7H5yh8RhH5gih+VhI
Y63WBlthBGKh+06ziUiwgp4ysWwReSN3XIX3AlOHqsbV8X4Owra5bQ31i4aAh9kkeIi6IdStaBnN
t6MPOUi8WSRJzRD0K6nbRqrGwx6oFdw5VUi/URWBhGG1cGpJ/qgiEXibfz9KGUKj146cfIkIieFX
ZhFIGOo89CN2wWwSRcxILevtZ4aWOZFa+Q69vTIqBSnvEPRmFXZs6XNQYdXqToNfN4Ochp7yKcOF
4fWf+hsoc8TY1hNNCnuD0KS4mS/k44zup8w7kiv03cxtYBZ265qqw5H+/7FTqEoPPls8A3uYtVfu
D0cU7xcfCf0WMscrkiwIgos8natM7NSTy33mHquhrs+RZxtb3RCjn/gwAmg41dSlLJ1rn3CZ5W1E
9Zjv0inThjKhbf3qqZq3GC6SLoPxaIYSxpZxBxgdSqmn7UElpwuC8pigFnVgFDGEskbrKaUyY+sr
mQCBlZpsvw3kXcM/QbCNpVzL6mDX2NtOYEtP4fkNGvCWMh5rvSPFXzilgBRvog/J4ucu3aI6PtKK
GXfiR70s+7c14JQRPvhQglxXDAdOOFH60cZmxgN8oty4K9ykMzx3QB8ZNAqkE9c7GYT+fGNjBn0Q
LpWZ3Aaj+qU7sBIdOr+nzHdFqET/ZFsJSe/UIcfrDKNzYRZDQjjCnF0lFbaF3k6z1FYOCxXG4l+8
xOKjFGUgYLBBlsLO74GKdhFBqWfdKIs6/wI4VDgnTsmL1dLOxFQn3cwBHVQu6dGwb080zjwCFB28
7uK52vWI1OO0itP4lUWHY0mliHUhM9NNh2chvFIoI7A9JVfRU4O5daJMUcO55B4rIhv2sn7RpisY
obygMsnMg+auA5Jof7F5/huDMhkTxQ3JL0H/mIjkezS71lPXvjsr51a9ETKpL7wm5fT4G1E3XDoE
80MV+m+DoQqoBYAyH++nsSXV1W2MpEVh6IOgF8pvRNmU74GxKqCTiG3B1u39IG31qgJPBSYNFqDb
KWZeqOvDBLQ0w1Rk4+zXRkpP5FlVcYBVtRW7nQN1yEd22Ixp7PmoMqHE10SGRw54q9ftd+mmE3aP
izFzyh4VJHw44jmH33I+UVusoUyQAS1voK4pEmJvt5oCLBNyK7XhWt3PJN0trNwhL7D8C/IT7Ijx
QcD1e0dvvNZrIcfw4nlcX8UHAVtSfhE3IzfdByh1f1aER6bWahNyOmMEX9vy8SVP/rSx1ksK19OR
Ua8JFCEtXTJ1tD3Q4fraBWdQ9W3z2YtzqKfoQv43cMXayyfhx7LwHWx0C5P4uLEBVFA1J96s3HkS
fDKIhE8iGEMgmdIn4Xbxi+igzThLJJGcO19AKb6J6cd6cvd0ca9jTp9oK3YXrh9uTNXtzdMh6KIk
a2tcPKCC2c6HYLYAYjKcwvqJdF/O6/8zNLkpr64z5DR/NzaQM3bI8vKNknSRM5LKE6YDb68j/prS
VZOoZkhxMw04kcPgzGGyXV4TZC2EhG6W2N+t0gvCsj99N9QwjyeTgJQePCYGksb3bhtBf79NTZSG
6m3wK+fA6OgeMi8fvzdC9MTwQSDSVqpAC9pF71b625Y2v6HPYyo01skK3jOnp16bKRlU2Qt+lyfR
yE+oQbZzd8KonqtYUl/vEqaQZzbwRiOG1Gf0BnZMROxW7Pn5ZOAUOcC8m7bNO3ZQHK44mGw8ephm
g/+UpAOzpOSO5aboe2VSyTBTC2q8XDIjSpAPojrxpLT5OpziLBT/qiof2ueKYjswj4AIV8zR8L5R
crZqvWsO+ncnlGhORDo/EI8cZrILqACSQPIyJuG5YI0PqOaYPE2c3vLCPf73WPnqK6xae6am7NhY
zk/H3Bcw3fFXh0a8PmaCq1Jt5HoFEBnrG/PGOE/JwJBfRt+75IqKTCZPq4OSlG0HLFNkfErVD2DF
fTo0Y/VVumVFDY2k3oWLRFWktHAUy+W84w0UMKuS22C8/6Jkou7JAvt2n1i/wVHFG1xR/jVKBCv7
8q3OdPeT3ssBz+L3dxkb6mPmu4WwyMevggVn+Eqam12hcnRCxYo3IROTmxj/YJPvmOk1e1ENAUMp
grNrsJMKpIqJ6hWD3Vw67S2uDoN/NWctq1gEf7VCiz0yVzKhA0795yX5GmFI/NpD9G9cuI+xooH4
DpyRuLxLabyeWeDROPTZHTJfi4fupzbUk9GT56z4HE9Rfrw47arVNr9+apKnVw3fu2zqnUeCnEat
/W0rB/LnS6CbaWyRPZLuvae9OmPZIIJqYBsE1svTR1xzub6+4S8SU80niAMUa8PkRiSorGKKpuVe
GqZzT7xBjreV0AE99txyrZF/BvGNOmQbrJnrZlRmJKtmVvXFysAcJXq/ve/wTBE2Gdsq4uqKjAPd
COvjJFDfn5HX1WI3v63E2bxwExFwGz3XSw3QQqDgXkGQ67Xjz0tYjZhgDTXw7iWaPnB8aqt8Yawg
0KvcFlzs3kpXIw8SLIUP0urLpouF6ZWr0KIJ4F0W2gtWkDJKAb89dN30LqlNTg9H0BE1vhnBI3zp
tJR4Ps7qr4s+zbZ7WctvP/Rd/MCe1WJULnp6AkpA8Ks74RqHqYzrBldYfy4SJ/6k1VznqhRHaPgX
MRvI88P99v/A9KIBMlISHprU+apw+22BujW803k4tBjREdAA94bne/MSVYCLQnfwXoFSGMzrIRjq
LEXeJ7H4jm0MKObeht7XBkie/7Yu6SkAZAU/Ge0th+ULdEDSpbGt7xol1bt0Mkkiuy1wsutCFR/N
gqXBXhVrZo6UdxTlBUALnXNVPqRwK1A2Ha52tZ53ga0C2qvvqIwAueOKbl03o+EOyYjgybM4wT84
MO0kVkXAw0ZcREgqHPrkD5mbwgTGq5z0Gq3h9oibNBuf2VJ5uXo4hF5V7Dy+OlgtiMLOIOr+IRGx
MvJVu5SDhRZ+BN/a9RB/V5c1KM0E9mjJSosQcEth0s6oB0rOl+OLiWAl295nkafyU406CwQJVJgW
1z8BVsFRe6OfSOT1OKfmEnoya+L9dmP2vwndYcKpWax047feBJ20rCTR6vr4y0USBZ7fQ7UEXnmH
ATHoHBhxoUqliB81wyXGE52Jh+03vDljghG9Et2YWfKyMC/RBejzrPsjTd5wrn5hOHBwcPjkam9S
ObdTxyDKvuj4u+3handdLvBV9UuJXJyW1fLYIrbjyo8vRYVMBIfachV8tEE1T6vmPfHt99cHNM96
H7PTjLdec5IWVV+XdBn7PWoe75NMnvqvCURuZ9BvUSdbCnEzvUenbhk8jokm1nEM52Oii6diBHAo
czNHQQEfwbe/gMndaTGUmQSFZpJevNBsg5ZIiNLT0ZwHyFKHLPEf/zOzZ2OC3MPa5xg0/ED0rYrN
rPASFcubJbjAe2W/Dzccn0G9HJ/fDL/b2NlAwj7uC2qLi5K7XJqpFjaP9SizdmpDj9RWA3skvEvK
UnWV3KIcJB75ew2pCIGoiaTK0u3YPMsBnLE+l+8mpucIBMYdDGo6E9WQedqF8qRBEUhj1K/v7sN1
bbF1ER2XIoa62O2dtp4VXJlfs8TLt7Otz4aEAWCVGw6q3yWSlO2Ua7PK3eC5RrfK41jKPfsRF7B2
zbfvJaiZvF091HhM5Ec9CAcudXPYieSyyWbLiG0tUECUUQsd35PLODvf+CVNTuE/+AA6mL/ATSN9
cpAqalZ8d+Ru4t9M5jOEC+RvpjqGtSRzwpy7hH6K3XYVq0MkaoTkLiZ6GvDMUy1U9MLs2+bGal3h
XDijAj3dPsPFRzhw0dFiwY2qzzPXl5ZU57J/UXfn+cbtd2Q2RR+fcEtgQqDRXSBK56cvQjleglG3
sDzUDdUZscrYwJK4qeUArXIB1eFIUbKFWzZLnJpFDJp8GY3FFle7785LqKEy8Y0SVUQsGRI9N85g
Ns07xiX8UkD5jPZUrvD0buXx+bn4ZjtZCmxwYtvyA/YO14IbWI6mYQJSNx/bsq6zLM5/k/0PebYh
pbY/1D1Q2MSlR4J3R7UeCOEKG65FOjP11hi0yr2jDrWfqdZqnlp99Q1xkuRe9I01cKKWYA/PFU+m
iGQbA1q05qTiqKu9A7AfPx6QIl4515b1DiMDliKkErbNvRXsGdA8EGNxYjuDwq+8bRqxPYKQPPZN
YrV2CQzvCPKPGinVDUYWj5GEnsL7t9P4vETdHd7nlQ51OGdt3IizTdaKPkpFi71HYzMHZzkCl+eL
7NApyiCWkzYeK2Yfy37GQHlGnYfT7vsfcMcYVTe1BgqlhQp5GsRW8bSDYu9NZH2GDT5JFHle+Plc
zPCcmbz+XFvHwgwsgGjbD4zWd23CdRA2Kk3dSOnoMLgczHqr9Hh1dXKGORXNiV0ukWoJkcunT+mP
pHIW2fnqNhe2BR8M0FR42atMIaD4Kq689WN+/fKW2o+L5FYhhxnJqgSKm7UqEv2I1yg1RtoQcKbe
VMyP084x74+g1KDkvEhZQJ9yStESODexJO/Db/xZBjfbSwXfdp3+CSzQtRJLBpacLnilLKmMKVLZ
1ZrBZWw3arqfMWK8OXPQHK2VHZMnoTM2/Eusroo1aWoQTs/fikq4Z+eTgJQe7vCEls9qoCGvqVa7
9woVdPjp5Qk3hf/q3mP7xuwaAK0Xi6Eoi9Awsi9BMAVRAkOqr96YQUdcLhn2qf70xkQKxquOaeyN
vlVE8RGiDeOoYYwpBaC7PVJE1ertMLtxn194A7R4DLYzk24oTkzDCKrw6/zRbelvXulQVoxVIsdC
vuBclIPCw43SCdaznkgForYYuumSzlBjmFIBRuLmimKCH9zEjXEpHCGUKGpnE4IwJYxGrOKKiAvj
BBMuW5ck3neRs9+uGcz/b3a0d13jPYNecATEwyiJg1600aV1N4eL8QA6UgocAPXwSeSif1355+d9
b9XB3dGkRibwNi6MGtnou4dhloOT8rdcwjALTKILvy9dgUIZypan1m4Ld2AfLmMuWar+89aSDWnn
DIOJGwzDzdgyV+7a//0KcRuUbJ/wC45oDRGNkodeCVaoRD5FZokEBUkopo7BDlbWERHHJorSbc0E
4I1tfbD/wKYGCmEbObODgRXKvOd0TokcWF0+JP5Rcf72yvBrY2JSv8e7TFaPNF1RPoPKPm6O2u0f
ugQd7F+od7HlKS/SBZIGTC4FKcgey2Vdef6W8otXPgo3Djk1LSpsH99z5I2JfAFAwD4JtCd6BFSL
5O7Xr59Na13B9onb06ryFrfb0kSqkOGvSI1nLys56DP7lZLA2GlHARYQu34PK+fpWEJzRar5lOk1
nmWxrqMcCfK9/xTI8P+4n+zcHWOo6DdumW7sD5ERybIjOMivqxbMcIslhKUqybnlgPrf+V3aOtSC
k6m+Yw4WN2JcWFmGvCgmmecY9/mk5iCC8xk56yDhqvA+kRrRKASBRrsCVdEVaDj4zsRfvamNX2KL
OlVuqopdV9Hc1W9b2eTSZLr19s1Q5elIfo2wPzp9D38QFrSRDfC8GYbQfB80qDEkBdIAKZCiRBOs
+uSgE5MXVYhv3R02LJtAxSvZ1qjoovoUBLGjHGFw39NRdBDVLFxzqzj8/titoAfCkflIEK1Jn/WT
m5wc2dDmRtAN5PU4Gu2sTozje89VT7QYCILYajuAzyCmMGT6dIRtWpLTRjkiZiG/Z7GO2dRDPkkR
ECnd0BtCKHG6KGNXVxxXxTL3YxoLgDqNjCvBaZ80u+kPs5iMM5qzNQqcJyo6Nzw81yq6yYRpLsta
yS3iGzpdDbN+AUm70s1pHnHxmzqtdmImcUTjrWKivJCT5l9g4nfCKbHRjBUMqitXKCnX0Z2wWciu
KdA438K1xJKNYn8ozYedMHJs9++R+AVXzifA9t4kuMGZl3SEZq/oi9GtRRvFcikX3jtwp+H5Qq/K
XUstL8eDgYxZG1Bmp7GQMgZnr+VHjARd56lY/I6XgZt78qWaX012mKS9wg6lpoY6Ehhw4rfQoQDY
MGFU9mUUT1qqw/96n8ZvFAJrqs9eM+v2nrAZ+i8gp2kT+IveAD7VBoa6zSkyprCcj8KyPryKpMCn
DQlpwd2hXlqV4saMdwztgNMCUHvjtRpcOqUL4YJeJePovWOllF4WW/TpkZSMYflgPFTS976IDQji
u1CWwQZip0KsjJxpAhZ41HH6o1kOntlsl0dMsqrr/9vyW64qE33J6pNJed05WqdIVKDXNg/XSCrQ
78YeTpUC6h3JAZoF45K4YlpcHk7n/big3lnRpBx8mwHYz0oHYWBs+jwYN4mbCiDZexiY0vylSt+s
QY1nWg3WSSxQUCQw/FYZfzHw1AU2hzTvi2wS4ZOBBpvHGWMhxLo/Fjsk5KtpteE5HjStFXP+qVf4
7IUod2d7W8DwqrZBUW53VjaW1tQwSNSVBxXExzFnFJ943b0NBhy/w7oMNpaf9H1AMxZlCurZ3yPk
2MWyRc65TVN0Ve6hjk3BmpuoWK0e/ANmkt1feHqslaDSpO5opsiHB3PKvyrvuoHYyZgsFjqwS4yr
6m6048kdxdD8ASpo3UO29/ajCPVn8HmgqwuK+I1PiN06ewO+RNRMoA7k7EDm12qvBMwSyQ8PS7vf
fJr4U2HkBLCvec8pJVh6PVce0Bz7p98iYYPhyxF3WjammowkQliy+uHsg/BoUvw8DwUlOjDyb/zJ
ZTKfsRQqR9JwEeKEwcFO06ROC6WT+kFaj1xhRpNfuWOCSt1J3HDaX3VfFiYZG55uAWlHtXcVPzns
QpysqfM4vWsRDFD5sjr4h9HPAfA6d52mltHO0iYFQiGD61dKKKCkL96GIxF768bNkhznIaY3L59n
HRk9EUIKzcfkF0TkZR6WmgUAR9vnHwzsrXYPG7Yw2cWY+fio+hcQcBfNUF6omLXqbNYUki3L6WuV
7omt0CTMMiUhBwuH6FcC2p9TSKniGzwkTOgd5bJsjqAKh3ATfJyJyAgDtYhQw7Hc4BL3HfMMEezW
VqVNO6i11s4cB8BMQyEPxdxECVp21iHc7FLFp8u9xvWpQa3PdrHBZ8pOfch3fteN8T82ggGk/vo3
S9LHQJc3Fyy1wW+TcYypl4uNpTD1n5k8P9AC3QWNDa25DOsaN0x6RtIuawyOmoyk4Wnd6gJ2rbDp
sZaSA/9esR3mK6zyzqEKJ8mC2iRpOlP7qmo9X8+KgDMvPIxJhnD7s5hri/pPflB213SJFV6xS8XD
mMoIpbyFNti/LiaoU4wEpk6scl95qx5H/PHjSCBcxbVz6dS0QYYw0sm9oM+Tbz+9CThGf3a6LVqu
TYMPVURq6wnQeWWhjL5gKrUroSZo8Neay5yKjrAh4gfnupWAAS7YLckUyhIQxn08moR9uL4f4SQH
F1VCdgX1pXTN/mmHX3wKcVa0CCX12D8QyuPchKzVIZciq/27osraTk6PPdt1OpMDp7hH+wbuzIhz
O8OJnrQnoHD/tO5kZjSbi+t8IogzPGa1+1RloOCBV+idRgTPszXAWrwHuwXPdnVh3CKD7qf3SB8U
Z9rEUphPxYo7/m/YQdipnqpcFSnVUc1v9zPkoNl1vvqp2X/aY2bXLFT/NG2X2t6xRwAGqIF7P4Bg
KBD2We3wyr2sRF3ZA+fz0elqtXtHY10rXdtCW1MtukFhwU9kLcHiWbsMCk8QhIKch4Tz42UmBxih
CYZSEZfdGsk53ZH8cl3otO5dgAw79nxp7lVaYentqf+Yl/ZSJsrTZ4WfyfEEjX3yh5BicoflHadR
NgeER/rGMlo8vMXlpb8zAaIrnvwi2WZhdW5X3zSwMVOqSkAOK3JJSVdL9uMeoyx7SMvzd7MaBCZa
pAPMAwAXoWfOkG6QXZqptN0iVShEtJXBLPlcsa1e+r/16PZr2w67uAjCQ4Ns6BoZedRWToXylzfe
AD9VA7OSJrdZmqneJmmmTodADb4fZsmBsmnovXiIGZTkTNnWfQB4OPB4pkdee+vM9ziqq5ryM/+R
n1l099ByPFsoAQYb2CRKIB8fg6II/5deeshhaLZHPTS8uPviZXRZVJfy0gKYRk1PogR2dsi500s7
NVTXNbK+NL0hfbhmdmYXg0kiQ8NyeHTgW9Ylhug6fDCghGw8fmpmFBeMkXLFKIkhSAd6fcXh0ZEn
5tHrWHjTS7mkbEv1Lzg73RmOMdWg2PoNsEYNI7qz0viStxGm5PDcRLvp02zpwHpzFMuZ4oY8d5qx
N93CJin+9egRVLqDKUmYKoI1YaRA9sTHEbwmzcIC3tKlpQvp80xmX07Uvb0loPtNxQ33dQw/mjlC
C3K7BEA8yUV7ri+uWhQu9Hvl2rXEmLrtkQkJgi+vwNpZ17zpwsbMzRjf1jee80VQbndGg4fLAkBs
OsGByr2Bfmf8XvhcBpeVV/C0fJtiVo6motFj+GlygGZLfxD5472It+eaqpjC6ENxtDHH3841rbdO
RWL0P/1hOS9gZdw/rVcZOEc6P+42//9cqN2/w0bCez6r9S29bkSspjnhXgNn7xkyGiN5vUbs5rc9
YY57PHqh8r2Y3AEEz4ZpK19sBRk7XXFnKw/8P+r7RIq+s5mzQQTJpf/lpJ3rOoACFW7+2Ngf2hNv
gfq6GwjZGbeN05ejHptUsAo7DfFWG/0azSmTZsfQ5QqAdtBBfZgf6Ax0ekSeuwQSlE6EBFtzLkpu
tjjO5RrFPwHQ29lO8t93t031S+Rt1yzbz8I/wLvTB9JlW3QHl58+DqDL40Sb6wp9nB88K1COuVOW
w8HJpo7/kFMXllPAXAhVQsBKu3Yh+269pamZ/xy/7NSh6wKxXvVL8YZJ0OF9kf5o7jemLCkLDzZc
XZL4WgHLYhAmZm1Zp9WWluRrgOdhiOW86q4pRO7+seCtOMUvLuMF6dBFHJvXHb1JLgJsqqrTo/MD
CNIcKNS3aqAdwqB8z5+HnQ3HMUGww/Ins9lbfFHCp+sAZYqJ/H3L6qU3fYjOU9+Zlkzu7JRxMnvJ
KQ8sx/wE0ylL6QPlb0gIest6239XgWeoNEWblJgsvo3eCPM4xjTeb9WxBpXl0JolMcze/nJhT4la
6sQTcAzT7BgRkynPs79gnLgDXbiX1yI6PgindFxGN2Ezi9lqVTEF6aDoPfWDA7rmP08J6UyXQdY0
/UGOrjTPojl/pdYMaX8noCXpmYsSvj3CQg9UfQylDdHhgoD0xtcvwycTqW0YCArMGcNXOIEDx+d9
CWtVkCGwW+X9AiKo8DgslLHG50enQLQulhiis3Ybrqq63Ua+Gmr1h6tqKnadp7GtFE6IpdSdMT0W
EiLINPpa6o/5TT18tInPjg01cg92dMttaFnWpIR1XEc33EHNoruuDMS0V4WXSuj+/kJtXDvl65Tp
m2+SUYbxbEsxaHbJMMWBQLSGWEkdlyOQAW/uySk1THCB5AIHCrHnqdp+ZyrB6obMJ3dM7Z6AkUv+
5VJLl0pT9hoRg4PGB0DEP5yotK2TJPWG6VoI2V6A9hbySCsTg+GvLmqHY0Hc1tKJXm0iFzqzaHSv
2HGMpxhNDAiaLk983iuDvDNnzLJJZ/qK3w9a0dYxCAH7IHoKpQxlk8Mxsyt52AsaBC9WWxyyT/ZS
8ieIUjSeU9aG7ey51gSEzSy8VTH5dDd/Rx8BoIanCAfg5kynDmk0K5aTQHAmG5aKrye1z6hbo22/
/rgVuPzK8Rmf4oOTAYhebnJ9wuAhzo3vigIcH5VRReZMipor9Xt2R7YBtKmg//JM73fqg2s1TKvZ
kPG1a5sO9dBOfYAckbo5frwoVHzjklRZkiQHZ2NT/sy6KF/IX89+QTYMFMSdG9F/luO8tS22le7S
PU9kx5zZ5XYTuor64s2yzvNRJ3MCdL9ipmS6YmXzZkd9PulwT4+MDDWaFM66jXxgm0N/q0RsBfIF
0OpaWO/8m51NU0IeHBodl5jMnZ6RbP0LHVkwgkfPCspI25ZsxATvBQ4oS0UYN8IBu1f55QeN0iqA
egMZyZJrZJGFr8yekoz5UID2RrsvYpFqm0UCjiBV3TW960FxtQXVWmjneUSmK+himDNXEI7Kkxte
HPh52yDeUuG3eN053ledSuRW31oCEv6mk8mulfol/iyFqtNzKdF7PXiGWBhU4hT2V0zKZy6C3Fuw
1KCE6f8Yb4iXESW+PHjnIAI77sjzLdARut0V5xYVAC6bQcoujFKm/f5DjJDuTBwQNgtpCCxlQMNR
YkwqAyAopdaRz1F0Lm1TOHAsS5beGa314SPUQFkuaiYX+Cs6GZ3w105ZTR892hzCuoF/31tm8+Mx
Ufs6WXjhETdJKQxwx6inDrIAClJYsqkGRGIOgcyzusw29xLG3/6rq3b9GKYObah5E0vdmi8k8LOw
OtIkKaETrBbQj7Q1ppxtNp8MWIJa6RU/jXw0ZRVhGkKxsdloWIveHqoYFsW5x1rGSWPm1GslLlAI
7vcWZJgdFTo91wOgMjS/VojvNCPnhVMA0tGLuU6jPwYGzHwMs4nG/xLn+AgMf3l+mW8WnuLt/ukQ
4vjl+Q7D9zBvgblF74h/GC0yoPGerWcxvBmO2VPtywyyzDtuEhh9cj2ReWsW6HbGaahgiVerqmQ9
lydAwR1Qwg++sITQkRMI40FFP1B6Tri2IRa9xH8p3XLVjDGhHuPFpgomF4s3kQGcqT4G+niG8gqh
ryFKzlpVeVd4eSfHeeJE3XeLIhRWAMYvJb96Jjhj0jUAjI8olWx5jrQ7RvVxMo1V5Y6sJG1mTNtK
bfh1cVtBxzG6ibhpIFZYALaTwjLUAwG/VUr0D4qsmWilPS27ZEV+BetY0hJ3vRe1AxGIitEU3EPS
efadQjN0yYQGKYNeeN/e/pgBAA1rJPq8JZZOXruQSTkt5mqskN4Ez2ezv86tMYY75yEgXY7Dp2NJ
EbJAj1m2H91lPnaruQCGNDjBn2dKbekii/5m3YqnuZRNBBUcf8SP7IhJK2k/LLblwrdqV6JrToWR
xTFh8i8vI6Ts4xudxkrfdyuEK8ys/zB+QVwPuagx+v7NOHsGlkkzr5Ar5cat5XsjLyZQfpe+1Eif
sNG8K7Pw+tR7Azy9vPR8rBBBtwjLj4m7N4sN92ngbtmaWQAGVzgHqnAH4X4ZdK0PKPHs+UVS/NLT
SnX6sBVXOayOa00BBjciTq4nVwy/ZXotnI6PSflMY1F2En+nEFUHIuuSUr+jA8F8BmRPC2XCIGda
aUSp+hEPx/BxARFEM5/p4MRaTHoAFbpmoTGHrjOhIG0ICy8X92yHZjOYep00aC1y95pg9Nv9nWik
PhoT6lNkCkgbicSU9Vsi7YW/76PBtOfui6AyE+Kh8jloYooYA1MAtbAfn9fgYpw/AmLw1iIF7SwC
LF1LJqiM1CleSBLCY9EAsFrhOWUQxP0n9oTvbb3tKQng8Gjgs0PYHC3mOGCqxrAfaRjwSQZSqN3P
w4i7MLoKlhh68O3A3eXRd+hM2C3mnKP9ODXEkKclVSYxNgADRwrXNi2SgTYlZ0vv5tF7ndBHn4VG
YuyUZV2urJcGaZ3aWFoyVnjohkAhkPi8eFct1FpTQOMIYV4JLHN/xSFvYLFCn9nb8u58p9c3B6MK
5RdL/X6LDX9AfhScvSoqHHg3zlod3hnRaRBSsA5mmfIbcJlCvdKrPTJcA67iQTscU3Oj4LEuHAwv
a96GZYcnV8jo1mLUM9lR05eAXzsO/yr9U2i7gjLeY7iDlSQb7zNWqzPPmdQ72RFYtRQKMbpEb3Cy
XXwaCuuEF/J+4CvqOfRCP0tNPiereTeiwGMQoddm4C4whlpSu0gi+M3gMCArFow/XhFaWIox6pLm
xLmpU02rZbJb75vBBV8E8d7QeVoBGRsFfhc9tquWcLkoy4QhbsgJzNu+Zo4/eLR6qq7J5YhmddZ6
f9vfJPgVWhJndKWTLv6WRPJck0/S6+2Cc2HhBhJCp31LFtDqV6xAK7fyGsZnaTCI2sbMVlyu3ALA
iVnrq3r0mp614W6axSmXNw8/Fwscag53Qx2A29tUK/Nc4RhKzKN6kka1n+onwxxzRPjzr6PDQn65
T2I29u99jEGGcI5qbG/VExO4orkpgLKKplZV6QwGA2/iqKB/rfgXlRZ4NXvAqWX/MEpus6zjKUOy
Is8mTQ5xqeleWbrYH4LUOXu/Jiwl3nBckoqmRjbooiTm4GZ3faqSLsMPEctcfYFCD8fjVn/lUZbb
chBnvslKnElMiPooSAYthpCT/A/a32PbVmeniyrqU0BhFe9Ste3CfF4Ci4wYbSMLeHmHHc55boIk
UhFXG6c5NlLBlaLLCraY6E08ojxaw4Iu1ZlQFpbI2ToQsWJXMkdLg+yg+lIg9fajEj0LInOIYSHA
KZ0Gsn6Mj3tx5TPX7KAr7jJi2LQxuANuSt5WA03mwj0AZvWFvk+ou8iT+V7Q4yOZbsJeriJZRJhA
GKImDgBEG7z2L4vu3C159EnFxQQa9p2H3QC5FIMMvnn7nZJNFgMg0gpcSNxB0ZvB/9SonHBrkbT3
gDxVB1SsLdsDg9D+d5ThZ5QiOS+6998U+6fC/Io1VtR1YV6X3n97y9SAO5P+mDzenuKTz/msFO3/
Ku1lu7d84EvUonxS/ceivJC6rR4jOcQJFydA5D21iBlLoX5oM2WuV2r0Yom+0B+TkM/I2kDw9gZR
eUOtIkOThJeoT9so8Hxp1mwGGYFB5P0CWGNtr2juta2WMEGy+ONvwlzyo/MIs3IJwFy9gYTeT6/I
01lWVOuI/c1LYfWypUwrmEnbzAK/+am/4XDoklxBMf6s8GddNRRiglel9Nf6HkuWH3o8bkTdRLZb
FARgRpImk+73ZyxHa3dPOawt+9WN2yR/IC9/rWcxOuPZaPxRbB0WVqvEGroMFLe5A7UbDtOzQqB4
9vyodCmyGPrxHB6zFko68WoF2WAY274lLmwIKayvJFjTHs9Oe4fygYl4CuVB52LD4ze44xmF0cbG
6BzxfVO25hKxDLnMJI5qHSyPGCzCiwoIyOzKWVwYcE9HpfYseGnC1Qu/rkazxdL3kMr6nrlAetdC
Zrz51Xebc2ZkB3UptssdPeFCOUAoSzoR02hfopddk/G3OU14aTULD6GcJ0kWXk/NPgmO6LbI2wpB
VgN9jsLxtHmQktU8mPeTSq96l+tHeIbIsWm9Zk04THDqdxbv4B8fxV+Os/cessz5rCIbmA39UXtd
QwLmFz58jbaC7IBqJ4nWq5/hVj7eYg8yKdMN8JFqye0xT3KF+0nKC002Y+VAGJOUwtPxw9w9hRQ/
iCEaifw1QF8XMvaJYQUFP7Y42wbdZi824aBiABtO2Y1GtYtGpta2+r5lc3gQbB/Og7PvU81EsPCt
669E1Ot6cjlSc+SSPo+OkXzUZlSCUc90a22GEy0MM9TIn9Uj1wrFfOH7vliTQbevaZc1pWHnNs/9
N+ArfqJMtlfRAp1EvKvltAMVyZSOGru8Olm809OApaff+rhywCcluRPBJPSgkb33fMy8qWaNbOFh
FXNPZb58yGpFF/Pqp2jlib8TxzTKNsFDT+fcjxtKiulRzq/U5t/kqKhp3m3tz2BT+G4LUiKEVHcW
ScO0SCxkc0l8KY6udDsTHkfGkV5+NX01m0KUXj889rA4uX1h/vSH0/gIGjdWtKdUSkZhlWI6v2Q7
PtRHtP5A5oxtCzyj5atBC9pojzer4uqMTh5i3qCuzHfC+zsm1y4e5QWRkMxw14hZ4NEf3/0EzInf
5yvOA+FcqcPmgXZ55DJRuMgcnYHaqrGHrXJpdMIdOFZZyFEsBa+6O8DwRqKao58klaxqAms26Hgo
EP0OGaid7C7u8go7KcwZX1uByjPHc5Lm23xHsvgciYcaizkASL96AQHA6Nh4bUqNdQTvQCzJf3xU
xB6Sz/aym3a1s8gnXwBAclwOdMoT3OQI8v88RD7hpNxLIrbEbxUuRutBAJdFLhhXAznhae2nnZBt
sVE4e4X1YZdCXA4q9bKjX9+TvpgB5Y9GsC+sB7GjIbl/bAosO3oXmx8OywL0qUcTvIIa56Yrafti
XK0u9AQsoy73xFd4ANwrpeSQH0WT/hyXU1pGVxHjo41AthYzBAjbXFm3BZYr6vW2RVCzEnXB3tNi
d4RjQB76w2ShWsKit9rOXY7CHfteiwS3/bvikWTorVv5DHlzxMGDVYuxveb05s9Af9gFURg11rII
OGNBfsoyRQDgYXpGzPdRY1NLA7+Ka6smFVxKy+5tCcjNmXk5IW8kgqyX84pqHR2FOPVCDNuIEeXn
JGVkhHpAeUCK+srAk8lhsemfmyHiTouu4NjAzzLYVf2lDtXVtA4RkxFH+Efduk/poE7LKchHm6RC
miyuadVzWWFBe1ODwpIJhmtojXzzj1ec0y2CqEl/zLjqdhyjzRbsn8/eiHHsgFt/6Cx+JtdHQWSJ
RWC06kMJDhw5U786ZBpLFln2GZgyk46X8oylfgfhmBnWd7fRgtBlzOLBfAykW1Viv4ygjpbOVT6p
1GyiyOZDQ4NkgA2sPUBAUvJvvZIQhQmQudBQowb0/HCWVNqA/+wx5BYtoSsPaiwWiT9emkHchMQ5
KfXenwDHHKQrzI69KPz8THbgATwt1mmXyhvafRD4LUAN/c4A0sp54G5fhs9f+YJbn6BGipO3iQE0
WhjUdJVKRJ48Tse2194LBY4ALzIzmFcGUe3MreUPxMQWsloKfAOw9UNmP1g+EJj7HkXixlU9nzVJ
K4lQgRyksBMidLTrCyawoKffSEtm827GZ813gXAC7Lc62RfEkLTxRdPNUjt3c8WgMcCPfpe3As2Z
cnY54h/fyvjb2LhjGKICv+UofA3inYQJelUcnWUTFkDaB4cJTe4C8bLF9dgHmBLPIV8jApTQQRJz
tzjR5h2DFl4dk0S1tV2Vn19shrrbhGJpXPk9XZZ3FF2tdLK3lVrQXAqdoM3vjNOzp4jG6jOKF6AO
cdpLe6eqVqWZm+sEz22/RxeQYnvZx1mOmTBRyZmQrMTjPkiM2kjctfTcGPqlqx7eA2znwnZU8hKr
GKpviW0lKBJJzOjCsh2LMlK/ha1r1A6H6QlcsfbfxVCK6f8idpFAjVtRu4x4YtlRBfY+qF5+Qyfp
QUZnOrL2K+sHXPdbpNcNiUk1fKp+TPz3kJPYONhdDJU0Y8+QF/GbXTvpD4VURrbAas2W3T7QixSE
IyYUh85wuYQTHq7MuCTo6TVhDzK+/IYjl0EC5lqsOu8Zcr/62V2Qbr9SRFo8rWhK6NqSeAj2cLr7
6t5wPaU8CqR9nKI7D4hUTzbuPlpW9+ClqGzmM7+e0BH61Li2WRVguApxj7ecKVFc7JobL4AKbSt+
iuoQ4vxIQjX8E4GQBUbQtnSSFa5ne7yqYBBQXPt6QZC5qsDKMFlTJSFXJ3O8rxoIVHg7HSqIjE+X
EUdnEM1lvZENe/IZnVuOfxSNpMNUm5n739Dxlufetjoy+0ovV7q8HoSXw4lctChV+tpSVLDfiyLG
rgoAQ5OSqC16hXokDRAHJW/VUG0qT8vYdzuDHq0kVfwJPYZyOXTML8Eb+2KJznnx8xYW+u5IIYjt
yLYuVVejTFlqzFHhz6K8VfDZlPxjKLM7PWmeTIhC9Z4NssDZ3HwCPE4tJj8pLynCJEJi5tBUSwg5
DNV1YC+hHNTN5yZaQtdXZjW1qnRIb/CHFhXWw1NSEh7ekIYp1jOnBTUVRmBHnevkFZST11S7MdS+
M6QtAsI0r4lgVyosfwOfVQu+eev5yF7USKrnToWufmgRtogL8ncV51Jgh0MUeVgu1JpED/+qhTEE
LZYmLDnnxPpfQA86n/JKm1r0zXsKTMwjQhmxWaUvDGV76A15CimwJLulWGiMZMD57tteYMzi7tZ4
FRotGjz2pvlBxIAOtPXHLzVBeQprRXpWesG4It576VeznVwinKP8IUgBZve4jj3D78y5h9IDtk2N
9J31Hje3IhRRlZ3/gXa04SFFkdGsZFtU3SPVLAdTKdn4CCuBnbnpbCogkg1nSM6D5uHckSPF6U+o
N9sxqlSxCEthv2oRnP+/uRkQJ2jl+wBHBvYWxSUxmVjLBST4U2alJ/bPado6T6OhOba0uwsR2W/R
07lM9QoxBIqQO5o/DdsW+EQK1ke8n6xPOY5tzAoJ4K0Ggtk5Th0DUiUW0W/bNWYLCYKy7/PIj5OR
y2sFtBm5xm1HCOYo7ndqDC4tbowLQlj0x6I7HQXEbjIaFonYs7tljvMtRVkwl64MHx3bauHal1Og
423/TrXJv/zwH03xPfhY9BfVcJqFMGUa03ZRprYeYJn5nOpyiFfkAOBujmI7ZbVMyy0a19oM3x88
eiyE+pk/HOzJgyzDSdhyuYF2xGWOc22d2JKlnRTyJAsqFcxYC0GjtLxpUxl4xqKThVKWAaNY7glq
mtd7rk74bi3G7s0RF+zDsUpMP/usXKE0o7+9bYyvll+QmytAXZwXkCJKBOpzq8aiWXBhkYf9q3X5
s8XSRUROmZ7LxIaDyE4YTHr4/5ESDqQAC/yshPBjwDUtikwEkT0Gvhb4zN6ZPc8F9Q1iRqrCKdsJ
Fk2ILXfk35BE+fBGgu2rYOQ+2dMr/p5IFbduo9YQB3CDUOYg1NT+gsd8i4GxadUf71nOpepxgz4+
u8lwYFu2NGCcGVu20QWn17ugApljVobTY93VcC0f53vBVo7TUFQstiD3XBGQypKWUJ2GqYaZw+Jq
q8Rm+QUq4F94u7hGa8v25P8nQHfaRRZ/Bcn28RXHbkrdVCfSav2bPNO8yKFniXikJkyOyliyuavL
ul6QJhrcMYWoR/pDMG3bu3hMc9E5OzLI3i0VVUjmsfWpK650eg45V24SnAiKtnif4eZfDnEq4J+8
iz+WxSwhx78GCKMh4sC7XDjyzIpz0rDSIhWOTnwUbyNvEVs/5bIO/AYBMIVh/TeFR6oWLrKDRiW4
7bzaELHKuqvidV7m/rV18CNNMGKqNTsBmJBBwudvOZtZfzcs+k5tVOYV4iR+7wnmh52gVaPqeCem
c3splICFe3H7+eP4JihFxShzX/1pp4kqGHJPy9YNtGX6epOUbOlmDHE3h/R7BKMmNRnF8zHeL4X5
SpitSd+ducZNU4YZveNhkJJxwGBLBzbtEhjWBqd+Fc26uSYhmEt12D/xsqOAcOY2uLoZ+Pn406u1
T3YtuM3bZL3uI9gKfkBTVM0OECiRBzhunwzj13sP8mOvi3VG1rBRyvphmh+jMNBI3lulFLmyMYOi
TIrXvfxFdOtfFB46z9HC86pygGtRwGfLmBzrRRs/st/NiEr9if3rETLX93f97gJWCycyX4A6jgJR
Y+QfykdKp8hlzBHbC+s79GXQomzSXC+5RmBJd7Bx02eTiIypogHuxIfHdqOamb8RjucEG325tEiN
BK/Cmldy5xvN8Uas5aAhhnlCtMKRI6Q+UlNnS+FoXQjS41KNLAPfp2Oc1YVYb4hwLU1VqIsHbGhs
x8W7Nm4O96CG2cmKMI6605ReakjUxypBmSvU0inT/1vVT+AsKCKTM6+VEGgx73Swz3BK2UwpUNcx
CJYV+YSdJ0ovVaaeA8D69fS3pjKgxooHmekR4jseL0KzE0sN2u0GxxkYP68TZl86nVwuuhCIndhL
z5+ptEt2yWkIIog1be3K74W1AiGdhLKjYpt1w6mq9ggWyWGjbvrwqUhSvCrEar1r6eokCD2S5Ijl
Yggn0BMf7S+rHowDFijbQx+v/Z6BC1FeKknQ3Xissm1p+BtalPy4Fuwt9/JcFR6/DrKXrfV4q78/
IitZUXgR1n1J+mIJYegQh0QFEPPrajqHKg1ogYn1z7frU9d+ucZHUzjDxOxWj3QVc5irnm5JVoNm
bnIikcZONuhZGOaQEZGVQTAPoqCundkNiecmlD3CTZFehahTH7oGA+nYMI9OkRATaRCehTe+HqdK
50qnNkH595lhV9aquyyjEgnpOFljC5IUWrMnltQ2bPV0nqlCRiDZpxZbrDkIBqwrTIsYhI8w7Yz+
w37BDorQ8fDvMwodEXptNUzx4gy1r0hdWUQoFBL6kOYt/ey2fPx5/aF6S6Afvf4QtwExurgvOW9h
mtqzDfMok6PJQWqusOEkx00iYh1qDiGgh9y+qCDs7ReSoWhgjysudSymmtR+sAjg1nNF5WMVfN4J
yccabLm+RwSCiCzijmJl6KGvK3u8zIwpjcUb+tad9AqCBrgdSW4x+y4amxjX8ydiAVCA4dY7ZR8U
+bXL8O8RriFuK7WQfNi2IEW22CfECVOsJqY+wN+/OnCJH5ByIsSDUZ4p6r5w4XP6FJT0WjmpzSJS
wvFwKq+jtVbyLAOcOAVoFVilxxVPK1f3hgGe5B6pWCorW4LdMfnkyv1NorE1A7HvzxNfWkhZuQct
6NWzoU6jUnMnEa4OpL5G0uJM95dNuwNgay1C2Kl2/wfJCVv1zGsU4oG5L2Abpct5ZcMs5ks16gwc
ndj6K+CcP6wuQdSyZBKQH/nGTgtm8QEBH7yGC4YmHk9OrSWROsf2imYOjgXFmtK9kQ/aqMH4QfQt
2kR3FMxOgCphllzbnAbuxufQn6v/igEKOD/LpVQRr6eu7mRGMI/9kzifwl1OE0JaD5tc0wiolBpS
IfGLfbpGGFpzw8F1/MCdqmmE9lLWC4sFOmUDcexvS9o9k13EtCE3uhlj0Epy50auU6lwDQNO5lnJ
0HeZkrDTGczRmKVzrbKKawOvNvyzxsP2yiuRNh4pC8YbtkfdxIpwJMsca4cgs9HT389hkKPDBnZR
c2m/irKZCWdhmgrbYDBS0EfK9AkfLovgOhQVsbUAy0P54wvO97t/B8p9jFob4IMbYdJ48YsZ0w5g
yDUZezWC7XZMPJ/UH6lrIiyk+do1uPJ2CCxuu3Am6F+EsRmJ/dNyNspU57LMRCNZ8Qx1vHBjOw7J
r23a7d+QA+yFe7YdmiU840vc0GkaAD6hKTNWw7G0VaUxXt3E84s79H5PpfifEpp2mNeGYnKOCQ+4
7gbnQTi+NJdOeNer7ON2ZtR0OLdvVYEi51jBrAcChJtj3sBAswxWLoaxuozzmcdrCd2IQ6rrT1tE
Q9tr65rx4GTxw9HzvKl+D8HR/MqfGZkOgsfZ1PYLRRUbs5ogcCPr9lw2diVQWpvkckrQeIgWfwno
cWhbes1uYnU4h/uRqHvBEZ6y5V1FtDO4WYMdBk+oFefvxaceHxLIbcu+m9XNSEiIg9t3ZRR//FnI
d0wQZDj3ibOKnfX+iPSnKtfcWaaXkVQkQ05OdzIrggcsrEh9oXIv2CqvvEnScAchJUirsYLHOvfm
ts3qIQA75Dwzn+xXKVCbWHGhVssXCy9He/mnpejOC4/gM1gwGUq1RdmMRByxGvcsg48suAPFtNfi
2yzyz/myxkUkOOnNHiorOTHk40erxxKSmTvSXMwNSC6fjHksx1eUGIqUTa42F7BPeU7zwGLoimu9
GRGy/SVpwWDUl/LClM1ZEzLCLjizjwsbHyrIEEcbR7IcKeYvf8//JAoDy44aU3D3gOJ48y2ePojg
9KTK5sUSfQ1w0HBGgUIpU2nuEBKhwspw/m/Vv20LYYXJw3GS9iO95cNfFGcu6YcqCg1fWdPLJV+Z
zvcFmtPnOCPIFDJ791ddxHMnd2h89U0gXrFyxRUeNhTHlIac6oRSRB8GRRvdxXeYhqZWwEMZQ393
6nT+CaFv3kbkz5mJlHgmXuAqGIdHxvdD8KEILJNe67EdA1pkHpnVVoLGmTAjD3F6D/EoYJq7NkYV
ZDuI2Whgsk+mJXRsCVgnh/66X8D2vH/1SuCu8q/tVHuXW3qTWHSqiVT6FAbz81nCI1zOJAL3CqIQ
X0YdwcSStbVdgCgjbQkeszy/xGpfNnaGZX7gWs94u8IN86scsTh0lItWXNtB+7GpI/m0vamQwhlL
pq2Stg+N0YPuaRdaQcp4a6U8y2y79VImQ6qxrdTd/zAaKEnRKjL/SPsYTo7H4p9WvjzSs4dIBzFV
PrYulpjm3rrNw6Apc0NVNsBbWLcmUtwkU9qOKT5BF0PSI4pUyIS3s9z4wagRJTu3jmGa6GgO9tCs
PFASYQyYDju/lBcA4HwIcHBjgsnHEUIINa6QowPEfADe3hdpNebYB3YkMGLKMUbtb0M7RD3S1hhW
skfA46dwgdDG2gfGNDnKvaQOK+Y/GMGDeqU0L+VnM5MxLaz+Jd8yx9DbX3ItBiETABnd4v/ty+iv
bNbUKJWzkTlP8gRf1Dmync0O+lIsi3MQHjsD7y10oj88W/9QXe9qCoriyaE+ifbdA0hy/donrglp
TvKMehr2QwTcICoYsa+L7CFrVzRRWxlcXcWB7C4ijfmrynWJLbUsDQXfqIr98lrPmJw5NF/WSxpz
ruCebMZPuNe6vZzkEurNqjiuj4/Mp6Em423IFOb3YoB0HkwGSIdOTM2WjUvrCyozYDI1W246Z+W8
kICIKQzcQLEs+qC9qsT8scN/5nuwGzVItezzPUMaJL21EJr3v2yz0GTr9iMJvWfi6VbxESCtdfjX
mlCWTvKlGvEsN0Hl2Ci4lt5qxMf6HgPm9lTG+72QYyLReq+l1lCg4FZ4L6VqmsSuoPbN8/6IjxGA
snDKg1Rw8lUznr5XCWtS2gXeVPC1dygCd//CUbYX1IW8YRnhYS87iEeMbqqL4CiLECnr/KopvCxL
owoo9lT7eyhMnjrdSbUYIfCxHDAqaHeI0SXGTcjEpj+U2KS0WRhmRKCSwZdrsglEzM00uyKBuoE4
CbBkYLZX8ZpzaE1GkbwmP35IIDQ6CDKapP+D1Uyr1xgZgyRzKdaxxgqQoiQlzdtzc153p6jiJIit
/twC6pYWsmttV4RGmtyHbmzAaL9KrFhTo7RtNl5SRDpQRCnWzeGtnbdU00c/XLe5AQ57MjviFRMw
F5v5JKLyqhkgLU7ZH7G/GFVies15LV9qQ/+kMFhJgXw7XHlJd35IO8zN8Mjxe4Q4FbUE+tSajxYV
NFHc6ZKVUhN6oDI96FI5FxUYkzHuzgDbdjlBNf79z1hufoe1E8NYuEeOb56K8hmSsha0/F39NGIp
DBSSCVBhO1NAnGFuS0Myp4Crj7lXqWQ/b4KOiwVrg34fh48Bd5SJ96dLRovBxL5IFszqqfKJqL8z
lxmxfNaIR1uoHEWhPb57elqo1HT1e6s+DRjtjz6uwh/KESJKvi8ToJfq/TlX6FrbdSZnurdvUd4X
NrYyn8gSizjpo5XI/KbThbahncZ+mhGEqbVoxVz9V9xmwFHLR0CZNjni70/pt/azl9pd6u30NsMU
5dB6QAjFIjyRsvyPGz+URoWF8wjZyEM4a3CDbD/izoWjP9hC6bttQvdnBUj+00Mha/XV5nR6OIy3
OgA7lwOa+NbCa3nRejTMupEtGo39gPVRo+dfk1SEFlqlJPbGYNT7/FJ+9i9jBzspZyfc3Fue7Oov
GgtujWkh+Gb/B4HKPHE8UrOpCr1XKcWyrYP08ucD/rbs7OxPLSlLilgRy2ZcIhTuRPfzTFAtvP/s
ECwGsnBKhBXyv4ZQZnOmspKupTa68M7LL4F7nvUAzWSX0cc8dYBqB6YfXHDoyxb5/AeTQV1GYe3S
JkiuDpdQrIfH3eqUOIHX970Bb3x0mQIXEXggMU3LMmTF8n2xiRLP3mj5cjahm1Ylt9AWnCogi8HY
T1XoJ4oYJbbFYfWWSnbJ9+3al/n+xwxSjckQmnlrEkMzJVtcOdG2gIc46xwwdAxFbDggTzRadyls
cJ28E5mdXOPup71yVF5MOlRJoWBGCsJ6+a3fbDkWQTXieOPWrqWm08ewmFdlD+t6HbBJlwbvJ6ui
vrBJ7wApOWIAM39kxjAc93KhRmTtAyVsm5fuE++4LBqCukrpmhlEBrRc06te5s8IkkPzzMV1z4qM
1qYTu0hS72SZDxbCZVzKA7HgkYZ6RpcCjjiLLulAWeQYKvfF0sEDw9bzKrmVuzVxGPFYh7Df+x9/
otJiBArvW6Zwxm6TRl8oQqak+neBkmodyxfdBcNkD0h30e+82hnQPTLwxOKWnbFyColLedjBIqaF
RV6yRwAR/+6aiTJywDlaW8QOcEFWpHoaQfa2erTOyk9NHS4Cn2M3/n7lbBJwGeoOF3y6ZXNR3d13
Mpeay5Vj6q+NMmmFygoSazMOZog2IDfC44QOLOAeVWAzLfK/YglhJysgaQa6r93HGdJD3WdDKm+0
XbFNI/hahpBzJtXLl6xR+TWkQAsMAJQ9+x8dQxBBobvj+CaGrbRvatij2VjTEx8hoJ/fYrtnsqxu
dusGL8UCI59KPp/jSt0X/HBnR3iNnkKt8SSC1BGZnmxOT1H4A8oMBYwQWKweWO1BsXZ76KZNQ3W+
MOSgf784PxcK7soAXx3LYzGwB2JR9ASbO29wGEBhhiFQhu4fIS22ShBlQmNiZyJXPzriB6LUAfir
dH9lO85h5uIgIk+rc3r8YE6aFqgHr8Ib7YvJ2V3pNsOkLmnfJSxmu36+NAnUUo5hr5VNUkbx6l99
zFnQQgufjuDBG+Rn1kL1kprz7bI0MnO9B1Do6mtAoDyWro7ooEz1rlp0uez851D92K1/FSYqbwcP
D/1muavm5D0kOmC+rUuoFmyC2UeHqZ5WgFj6kvyVfxLbbFPJX5tiE57VXqnOGOBc2ijclTa1yoVZ
PuLXacpxhgVcICSRLPCgSLAUsiad3xVnemnJy6O6BNM3TUrrCtP7vouaSs9uJK8jWRPFlUdJStMx
aDZyuzwB3Ny0kKszpgMG6dnNEnvkgD0ucm4Wr1NrQiMCdroVFhgXrNDF7gcaUN/dsDH9YHAZbnaC
mdj9hhOTqQhr6Rw8dhfo/LhZ9kQqwFwWmGB8zlE4gPY0UqyFHLSu1+7JH3ltx6Q3HL1vmdbyBjak
2kRnCH2Bu7470VCKNr9u2KXZPiYKvHQfdYUIg13YYoq8TWpxaR3IeKfTYlwwj+mzpFa/8dB3o2lI
xTK0WyasTyj+q2TxUsRoQ0Ny4YYJMt2ejcKCaMfbNDDQgErli7zJ0LkyC8I8SKFeWRiUNzb0ks66
PW3ayAnbC8SojzrnXEZIO88Ezyh9hEr+Fe68vJBlyUjWF7d5zOZJJLofXO4BDT7toyPzsAUGcig+
8/+yVWQSM50FbES+GLvtfq8JVWL1CTdkemcEHc0ERn0EPvdpv7W3taDKhwWrqiJx4I4NOJdtZrq+
Mty/XgfgBFb0YOf01km/YGwn1iRgQf2h6NEP4JSuLriCOW6OxI2nRS3+T/UPzGhElOzOweZ7lVJ7
Vqa6SdzzxKTuPv2Q1miPKKlzzR8DRu/P1fM8U1veISYsFCPd5p4XUrvJd/bKPAa2YGO+6omvytcD
7UoCRu+6+7WHWmDnZQuLL7bNB/W7xQ27kXRpSWKX/vc0XXhE0CXzp5nBqP9nYBQx5eJ1F5M1Srfl
NbRoBQrdKz/5KTdJEwq+I5j6ZAF6uaq2vD1mNtbPdDp3rIjk+w1xqzOgv0R3R2hlPpihotIKq+st
9KfdC37gmTairHgOolLHrVMok62QyG/Kli3VJd7xPiMlsKsPqx+puBj/NU4CN89q/bItgXiF4b+0
TVBcMy0Di/fRfPLqHsjAxJVCrkg7mJQrRdLTM/6Lez9ebNfl31jx4/FDuYnN9I47WJ1xI3wtu2HT
FAl/iJMCHybvVluBAXQN3bv4DIk7xgisbBJjZsH3/HyugWMqrmJMFVfyCN4ZulHDDD9r17gIvYWp
0jAjWRx6TGi9WgPhCMWXUX3S6CIn3wqTDw4xl1pEP7vIUSa27a+UeWEPMPhz6qfu26qbPfTAZSnf
FK2Tcytnmp8rT321k21A24IiRFvfgpTUD3C9lT6+WUU5IZ2uBQiiN5DTO4tv1QionUx5R3huA0Bf
n7vylaoxC4c0fHp36a8pmzkFV08XpqEyXtLRfY+pW1JNILupd4lFk82+GKYN6GG1ZCLpkzy7RrHt
0PSt/9IVhHxK8GEE/tqxTM+V8yieAKWTscz35k2ux58Cfye6J+yNG/JRGP1gAsZAORMEBZWYrQ1i
6Nj79KN/mvhxZm7rHb2YPPml6upEU9oDmbzQ1UHy3nz38YiWGNtomkdUGQv+j9xp7xNd4z5uhwpV
P2GQ9yqJVPzMfrK8s0pGvbJgNhfSAJqIEYA3TYYVKZLeVm0RReSI/KQ6vy41aJ8a4WKfJPkFmgiz
yBsnFFBuB4nZtVUJFLdta3/2+AKH60Qp80JqPaepcwZojawUET4FyOdwYjOG9MZ8AroyYoDrSOpH
DZsdABeqPRPdMNev0nXbjsCup1O4R4mDtZYOPXLXa4n/hvTOWkvtIvi7KIRfdxnd7E2ULJNtaPvr
mNbK5obCk+zpdKpfXTPZavDj+FpbcE0POD93wibUxJp0+GFC0h9izUp9dSzVvjXDRnLXUeGT3yEb
rD6Htjc/rBFkyEffRWH+OWYG/tsbh4aQ+uIFDeiLlf8UtxTd/81U4KELUhJW5CAJgUPX+MN4qJr3
JgZMWyKv93H8Dzjq02mQYRF6gX0aUa6SW7BSZOUF3B2ZpPcLaQiJq7MmLIP6TzySKCtJWibFWnNJ
wu4pqQdPZOQ5YcHpXV+68llqF//DSWNT4iorwiEZ2W1s13ONsgzVNz2bkjaijDKjOFcd8xB98KwX
bjFraNSju1xDyqc9ff3qwuiZrY3VuuPvqg+k84OGotlmsdEGtreRU9mmIKRuxU1ImL6BhC8RWgp1
n2gDfVFOO8vlGRbn1jiLeMWvWUaFa/lwpWc1T8NbKZFgcmdnQr3dKfiYLF3/SjaRNcrX1eibonUX
iH5hqr0LWy5lWvQAKkeh22orbG903LHqOgR4uDSJYsRpjJINC6I0yJHHGI6oQkNehKxRz63TLT5V
PTVtYxamDhIqGGdwJXRCqhAMd7PX27Qkk6glKS6QRivL+2GEMpwRG2qm81aPiIO8AkmOcFGzngT4
suUUPNNiMzLIqA9iCUxnsv1jhV9qS+6+gTTXfPY3UutIp5cZi/9eRQM61PjmCRFnX8utE+fEWtX4
CRFOYxdfscueb3kpo0R6UTLTF1DQcxCTbN4829LuTuJe/92jcJkcAl5FmkTBpgPQYz+5gIgzWsrE
Hrp8nJbbgLvSiWGH3l+M4Dk0ztMK6oLN8NiOJCeTKEMl7aJzM1i5TzhRWCZDBQsX4fqlZ1tt2EGC
JPz4Q/pgi5YhflJosA0T1GAYt46gCbQWO4w5bk2rYXuM1xv+mhSQoWhf+RbqkA34saL/1Q97Crjj
JClXP81xeb/oyEi0hUeIFo0tCoJqBkIr7oUG7eXEsyfCHt+jwdc6t0HpDiewcccg2q8h/LxMOVqR
oJriLWGCWbusLTJkWtaqPCu4WPmjK+36o1SwcAouGqi/ifZsHxW0THAHukX2HQEgNhkwf+xWCd/e
06Km110sQDvAF3u/ajDoyrv8xyPZzd1jIrZ3Dz0UZy383TmyYFkBGzgcykMv/X5VEDL9mRhc0YEj
dc0f/r13IseehzqgEU36hzaqLQQRI15ffb3Jf2UefH/EAVbCA/E8or2mLUjJpJnXHxA38mBZDayH
Sn5NyOscsXrq60iOlEGkw58NyjqMACR8JSkcoV/r54wRckYeYJqjamCyvioVJnL3iq09xXzVcVwd
vbfo0ZX+FHj9NUoNixzYo1Pk2Gx5xTx3PdDKRwTZ7zf5zWLiPuW3Wq2AtgOZthT7ATaNFrtKFkug
ou2THkC2aQIgcSNE8koPDrDfhqIJ9Uf7iY5lRoiavCnJFTFtAeWtpnMIvOQKbJVBDKEhZ6DAp2O1
g3mA+Wx9RW1ocQMjL0xJR++jUCO1FCmO+usBgg9D4nWCiFfkiHMJHux5EaHKcbTzy9JoHp17JefZ
xtIkonea4w8sE4ZKO02r3Ute9kviiiySm3IdDu4c/13IGhBaMZkhZ2B86ySgsFZzzwcdFx3fWFCi
OXPEwypuGJ2nfpintP3oWf1luGcymPraDUL627QdJLu0rJF9XpBDRKX93xqb42cKZgN8bYxHNJIZ
QKY/KKfQ4PFLgJh+GIFid5p+xdS6p03jcjnYDPQ4DVnG1lPjTIkhiKT7YO2txduXT7FYmaHSTHnU
66ZxSriOPIIWRpsPUqqYrre4kIxNdcuTm+A+4YX9nn6eZbGFDQ5S5TQnY/Fpu3uzptwcSqoGMmQw
yj/f9ByM82PKnRHFdCxXWWItHUJMgXLk2vQcr5KwbrfnVu4B0zAnKtcEYZEn94pL1+0KEN63jtTS
zwM4b75CDQ4TqO6icdz44GcASUDRbr33l8u3x/7oxd78ZFluPOih7zcH3yGvXeSgMrvI8o36bjYS
eu8iuSKB6OMJoXYWUnhAPfA43yl6GgYnNevnEV06PG2XT1Ycf3vah+asZ75IxT5juHrf/8aJVZzq
51X4uFaH6h6Ro3yqqq6EVmkUaOJfYnmIAQUDJe7FJX7z3X3Y5nkQDQNlxuiuTAL4XyiHya03MWJX
wlpkJ0NnFgQC3zxudjxc9eyH8pXRP88TSbLkw63omemFe8XguaINkPcUeG9Meh7nUJyT7b8LdaQR
AW7BBmuiwrP/GL29YjbLYJQ0aThIr5oGECSzkNQONWUyc9tdoxJrApn3WbrkVkFcS23i81iJZIsE
KUtzO6wFq2aRzVgXlG+BaQkoQ/dAYL2OWRO30+oft5DWT8jhypRRgdNk7fMk3BIJ3Wy3tySRP+V8
6H+2JBUiln5qpJIiAaUDOmkl5fktzVCyMbkqFWl9VoPauylFgqtqEeaaK1WLz6vE7nMAZfddEfB5
uxTW22KkybjZmAqGshgd3uccruYygkNYrPDW/NwWcgpacpB7cCVtL9c8wHp2hyVP3L4e90yn4PCr
wARreKnOsdpxfLasFca+JPsVrtWgtgSK36Xs4DCL/Y193RZuT/4fKvHtu+UuI0a0pegsWrVdrSbi
4n+2A3SLYIuHEMRhIAyFF7P0C9+bqaYPGcoV/Dg5rCeJJfsckOQNYzARoHgNXk2H6skuOf6sSor5
nDp+DeROZLSTIN6hRUlgrKXTuPAIjDWSQbmaodT6zZwxB8FUeV41RMAt93oEl1oD/ZIFRP5w3UN/
SzomppIE6SduKxu9KxxoOZpcVPgTvMBqG/AdAR5STwVNAn/b3OfYrC8WX6uksrtV1LH9vHJUWx7V
jUthCwWq0z5peYRO8pQIgH3Rv4JIrUWhTisA620CeLoljZ7YKv0Qvw43t+jxRpCVXSO2cXLQ+uev
1bk1s4thw2pObAk8PEmwVffGPQdvIFr90fBfbYmy92hA1CP3btLizb8qPHwob6vkvf7970Fod/0g
9aVefiiIL5rpp7Pf++f/Sr6DrgWzAvvnApCw7Ima5KMaf/b5o/p80ATjkeeNdxaQp7oaOJfu6mU9
RnXdmCemwJmcogSek9aaEvIMjn3G++P0ruRcWFezs1lZrj9UEZfEzY5K39POilWdXKIo3QnDAmnA
fAK+cNah2ZD784pGVssJ58r/NZJaPeU78i0/Q3GJqLJJ/cYuRlAdCO5OHJX0xKXSQG9IDe2QijdO
NJ+yOu/yUSOWGHuDw57OHJ69uwVISp24pgVY2ebjprrjSEtQ/fstsZkArnH3v/D1FlaxD1beSWlY
0in6fd/+DprTOa8Zn5ndGRL9g16e8Ei8gJ6x6nsfbQMcFQLzZETHpgySJJR+CIStdOF6WdIPpomQ
8D36xQ4ujaTPj50b9yHUu96yBGd6G42XbwHK+Ypo23RpKhW74j9Hc7sw+AfqyheIl4M4m7Fv8uzm
cJvla7YBaitQeaFWP+ReScW6NEc7HFgQYcOBd5mzcC4BrGEpuENrgKaOsAG8P3F0GkETQrToAQsH
HlZIalgYI/Mqy2UM91CN32OP2M9YojCuX98KqjP7IQRapFOurjw4DU2KRFC+N20hny09wjAJgFjp
S9mTXJ8uf2r39AZEjt3SmVsoowdbvFMhtnho5xwBap+UiVBXmGLaqIn/DF83xQFdMSUoD4K3M3s3
SbHavjQpymn7fW5YcW2UEmyoKRKICFR7TakjZDQaYGNkVX58SbEfNpqB2PLOxDivEr1X/v47IJFK
jgB1ohdjj+HusF91kVAcOb8dQhnXpXbQqjfbU1g8Xgc3Hy0lzwTNfxuyDWB48BrzIV8mNxSrZ5iy
jUQ7QqyjcfDJycyxUQsUnqAhKjjaU3CcrXt/W9uqNaK5kduqd4EJaVvp58qtzfvYMFoAhVvQOPVG
KRUVJUEWHXqvMH9c+4VhFycljnKmsxo49QOTJfPGYN/Cj56ShRresl00QxEhZCPQdrooETxZJO0u
fe6e2zT+HQxZBmKfmwNq4MlbeTI8qTzADmTEm01tGtpTWNgGX7jbP/ajaO3daWFUJo/6YjiOMK+A
BCiP4jYlLUeeqH62Bbwn2hZvo2kxNszeDyaRHDqCzz5tYk00PksL6xTyXKum2SrR9MI/0tUyxDiL
VHlBZnPogwVZYIR9ASfjwKeEEMtpfeXydYrfPIl3gjEZxfCxHqnDfecw9YdIRytEXWRSFaNH8WPJ
5ZCwQbUHOG+4lznxEWZQVv1hkiZc5iWpefxECaW8hfbIifODExgCH8hJIGXX+HCV9Yb0ejpkfuqT
lrnLY8AwQVWw2mOqdjwtrJ733cRzI3vhD599mJ9+e+WJ1Fd3izQelo0YiW5TXfLCUGMjZdWkWCYt
CK/PXk8G1NO4fIoL6Wxpnan/tuW11ea8/eWqn5KZyrSha6Oqty/eHc0reIu7LQ4HTTQ68ct19mJe
R0Kr9xwThnsYfNrKLCy+FLg9chlw1jhPAYJ7S9UJ/9VXB7sYFgruZpQLRV+Y4/h2HOzBC3PsTgAp
a0ZKyx7qoo9vfD8aOqg1y9c05cefmORPpFJni5a+YGw8/PAYuZ/oChW6XXEQCW2B1FUU4AKJ06rp
jzUtmMFCKN8e5L8kQho7J2Lo3tXKUW1ANEWAlxPsq9cKC1byCqDv89mNKnB2Qynr57yl3QoBR4a6
MB9eGZlhSVZkrhbVAYMJNpJE2L5bwA4clw3Djy7/1hjjkZvJ91Ig4pcB4N4McEgGWl5pYMTQZ25x
0IOijUfvG+zQWK24TPhngQ796Cnm5D2yVzR9ne7wrP1XLIG5vQAv4Fjq9DNNAD0XF6UEq5XoCnuX
t/KJGao8dvaaoqiVB7pcdWJDZ71V23AFfew6vFxVV4Qv2GlzgjI/X4nlEUggidcJpYPSS5Ai6ph5
LHJQaidOe0m4zJ6plhNh5v9WFxhWHJDh2g5qTVnaY3H1C+hoQcDhxmb8eTQ361kpLaX9mnOBkY1f
AlKr8c00nhSgdXJeWaZ/Is/W4eGxf8f4SLN0sT8xvR1czNNlC1LS3Ow0Fw8Yy+M4lOpH0foSO2O0
XYznpbVK8Xt/8ajY/Sn5YriGmBYQ2kTy3UYB6bPsT3jZlV4bRQcjpYfjSnYQoln2N4TeiT0ITDTs
k1JbOBQDsIPmfFkcZxalIZ9hayiLE7o9zJkeDpSeUBY1SrBzzEGSrv9132AzU4uVJqDekSJUSdeG
WGFxO3XZfu6Vt8Det9sYUc3MLyCB5zJAbe9Xznkhc8DD5vVAAHF4G6Fw+aUx5ms5NDW2SIJViqpo
XPUOVL3ARc5SscSpjQ7SRFXJd8bRHtrt+kw8XM6Al0gA4Z8ch5+XlLudPoTte/y+AjC0xLAQYUTS
NLf48S0WPbvK+JxkbjVWK+aGfZW1DqHHdAf/Uahlfa0UHRwlvXJu+/E/mX3j30n1rxV+LIJQmLM7
x4Rnt63SIoCQmNBsB5bJ68T4dyNPuVOFB6tvi36C+PLiySNPREzutXOxTQ2l89ItZJ9vQTPM4cg2
iF72v7xYCdM9ALJgJPhB+Dqd+u/NTJWMMS0+y6qurnpdBMNz+oGRwjOg2iF++o0mMI97bJk0VFjT
aVbZ383YlKX86PZ7K5NMRE+9xMtUTJ/ISMt+GJQrpEjDkAwXbEDJWji+/i6kIEm/29/ZZNUHL8Lt
qfi0q96HSnIWQVzBO0V8fXab6JiXyv6cWtvat/KDigtY+tmmWY/ybqMpH/L6TQXQiIEhA0h3vb0V
UnEpguwqV95Kf3NbanKO5bhoA8OaDWl/f3eyZxRExumuLSXY6+/7bQP2Ht9rgI22EvNPiw6336Wj
y5LkSFCSe4qQVEEoiM/IxreDCiaZ4bAohzsiNwpZ/X9lvB8yARBrwXcGLSGYNTmiN0COOapy035K
Ef3TKSD8WislJOdyH8wWmXE1ALrcMo7LfVLW/t8gaGMMzgJ3dPkni9etXfAhayw5GCTxM7UCIAZ3
yRA8hz5sS7Pv5JAj1xmEzhNmwQaVP7LFEZH6cGbJnobZldRMhgi/Vk1W22MtzRREFOaXy4Eetn1I
tUiO4q+LQ2AaAL+WNHh7nCYEJVwQkKPSV4Qi5Y0Wxj/a9igocfFvqIkMulVQHDXbvSeIp3Vm/KJv
5h4D/r5nstlezxIGAJUth7EyaGEEaAw3OMPPMW3pcRnw6nNQ2oHQXqa9/2Ta93jc386TiqRNdSwZ
VKauDSgZ3aFPJfpIFa3swUvtiwK1MJRMBCDMItqvNQKQSmwpNsj0FNjlzhmy/GOcsw4vg0idOAVk
Gw3ZAHRzChN/wV2T8NFYrM+hIQOC09uBdX0henHLDQ4u/94L06O/ixajyJMq9puG1pmmghLkWZ0a
r9lYB4V1vGL72LbWlY5Qy7A7m5ZLWgB6c0H4iiuLda9wxH60w/5SlFfeWqy3aOkq9izdsQx1hP7P
w5JB1UCO//8uJ0pHHZKyVRED4smwzHc92Rcecr6zuwKVvdHQ8SqRIkPZpkoaz4+3cg5YAMzaNcem
Br5i/1UrCrLhI4BK8P+vwl2LrzYKAJf6kUS2xya3lrcz5yfLi5/wwkIHWwX+LlLQclHFrRoEWE8C
A659WBMYViJYpuXXGsfDtNlFBMDD2D5+7+CUrcmbxqh/ujnKgISUTcUWMQLzAd5C+PlaATW2SGoc
wzY0i5S+rMCeCZmH+Hhq4sgC9IlT33kXVDRt5p2dyaS2XlQE1O7FpFTxMiOo6uuUgj4pRXa7h0hZ
CjH6yzDUNo0wOrtl+3KHGuq4eO1wbX039UBZiolHD61ZyqEHk6VRt0fBZBh5RxVywn3YHFZV1AD7
Pok1kmpXRXP7xE0Ic+b+oE90fYqOmSih5BybPs1hgzhz1L0MN1gN59FfkNVDQy/L+mFfoeBNFa4z
b+NElnFV643i//e2bWC635WYT+6PofpEiMRjXe6DMAzLXumLfKtIai+BAWRfsR8lJPNV84ZkW4Cl
oGPyjGI8QxT+GGijTtHQYDnxP0ywLoStcNtEXT/houy86eMjf8atq/d5iYzLjaZwLRkc2oFOaz7E
ycRIz7PUWB+qa6XGJntTAyWG/r+qKM3bX/N+PV5YoivrcE+xLelCmerL2VXxKNHnoC1bnQZ+COkL
0e84lNAWh9sPxAObwmdqMiRyYPoYaCO7+iYfBXnbBhxRFPb+ZIkj63Eap3LAS7RJCXVdbbsGVgE6
fwwfyIn/zoyBSSPHWRh6ZzcfTyeldU2i0/0KlZrm7IxqMIzJB1TueOBZswgPNMCJ0+s7782K9Jn1
2pxT/yc/lIY7zCeImsLozVhCRr17W+qAMLravTLbq6V/U+RHeyCqtTyxp4ctKdvZ9V4ZPc500D6h
ZRuIjVTdkRRdxp8SJa4Hcsl/+OQmYDN02Mii+xeJSNWK/xh+YJRCAJi4PuzObSRVhS1246pXsx27
v/Gf4kteueLdhlqxCbqKpkBEbjeFrqN/shSueryL8Mi3iict0NRXoVvORFwS32JyDQr+ZdVAaJYV
+D97NWK0CPgCqC3SLAcQTPcxSlAOw7no9b+YSno2zOZTvrhqWsCIgE8p0HwUhRn85hHQ3Cs7GmKm
5JX2prSxPecex2JTxW53f8J4LSJZcUZApeMzqzuBlmbwzgbZVTMnY5/59da1GDQlem2TqLbJG121
NBgeJ/lvIcGisTRkTfMuLcR9B64vW51BmyRkNQG3Ed5z3hgIPA8uTMQDYSOexblqustIQ6Dsbfpg
o+WFUIqfAgk0qkoONE8ISMHWY2J3CCyz7F3ozLkBG3+/dyzFJ3eBoyeTZE4uXi+KL7WtZp6nj4T8
MW5kEl36mWD+6Jj/SlR/NV4amqVOBNb9Qq8Oxy2+YoHfiY3Ps517R0u/jzuP6sFAF3Fva9O3O9i4
+8Gu5Cna+6ZTEYcKyoChGgjWoRkT5u2B6lMG13Qj4q74H0DLH6Kp0jTqSUbFaLjjyweeruNu3s2q
+qdbAuzvjiLjHnh7CKYZP/iy1xHQk8bLBdxlUOS9BhGXJb2632pEtolrdqzErY+DVowa5ypuP88E
Vf1e4IYQ0ZMFZmg2nUAL5A1IQ9V30lzKX3C52R2pm9tIeEB2QA4M1V79E8Y1Q92N4VcPhDI0FTak
CCiR6R3sPtlPJBmeYCWW6sKmeu7TWujE66A6E9BYOtOoSOSaVtbj92bUUZ9hU7liebEUme5QJ0sl
PwDsMrUHmNw7jtEEuq2pQTMHhLXN8ub+FvhFMDsr97krLeF310X4iqx7fv4pnY6Q0/Hseg0dCpM+
WsAgcEiJp4FOTi5a0ZzRQdibCqUQbZJK/Fyg7T6TeLt6fhG5qm/rbmurIkwKK8vOt2jvknMxOlVx
4oqJKCrObnhSpHwjDa61NVwIMHNYcvKej6LZcciMqUUxQv8DCCjWy9Ar5XQwbBdSGTarvcsnpBgr
KUbWulp0baE7HvDXPynp4KoGWNYXz2g0WBJFurp+XmcwBG+9aUk3sm5/CEfJ9EONp02fRNjG01Ev
YsHqu0aMtqIysar8nTlaSPAlT4iEMtRoktSVsSjp61VKylFFb1eEOAT+RT6L/DkAlx7LZkcVZvdw
wawP1NlGaDce8iJriyqHBhMYoIBZ/ZzyN38iTn9Vt1vEzYj/zTBVQEcflOEGnF2+y49bqD4xjuuE
DD7g/3eRsvZLmJYxIGbmZmOipTj7F9FO9vI64XQcGSeKeREVSdKv36vzRW8lqCO5BdRciG9KtRju
dQAaAg93j2cixm3bFEawwHjV39kyb8x212y5bhA3F5vTEMXqp/XLRsS7qYm1SV/6u7+r/5f00epF
aOA2Dx+VtC90Ja8hMVH8OGWZ4LLuVPHdTA/075j4l35YmjzYbHeimQEhoRYXlkjpN2aKH8RdkPor
JH7yLT4h8phx3YuVNqF9iRcoOIWSbKnxPpDCtxg1FMzWmtSkkikaWx1N0R/B9PYuaT/03KtfxhQZ
MbFNv0/b80lzgKhL/l9aLKcvvMfVoMxQYtKSKgEsT9f0GCZGSVoxcXnMrwLAhgr6pk/6nq6UA5jh
X9Qx9km+4x0nHo52sGv25bY4+SPLbJmvyc/lEM3NAaBB3BVEzgIpu7tom9fD+hR1fOJUYaKquE4i
AYjEPCzLukKq7KsfvbJ2a/WKCHKTB+dDGlXcEA1gDSwGa2jRfLymlCLk81gnrvbX0Wg0bAVsMHl0
XpRwoYb0FGKVCZXbGS+ilRWYAGPBLRMNW8XUXIJYCzqo6jA0RBB65V1UoYwSUhMQtygVHAEksFcQ
87C/otIFzu6su6+huPFfXlmeJ0DP/cRrrKvGzVEn0KpX7Rwmspm3rl418PR4FDQovxr/ODgPNpKn
9hLmCHLWNcnh86rxkkxu9KbcHnVOo3vKPOLrhgDrkHx+e9WmVG5qQ8JDeTOhx2bOlFEMW81qbGl8
AEPA9ZG7qsahSGyufb+LSy9wsi8/jnTAybbh72AcRmsSaNadUtCvpUJndYxwshn4uYuURTWq7N2w
zmCcOBH9X3oQ63msRx0ireBqWJFQaxZ3HE2U9RzqHl9roaKncRmS8OHMvYln5G5lYbX2Wip1EzIu
lzfkSRxfYOmHR5IqtcZkychIYzmwLWmJ64QBkGl99GeG33QKjlGbZkzWXy1/Yxt7ZP3IaiZuhE3w
1GA3q50NX41PXPA1fLsNjiPfuXY9qjgZ4lAEbYGqc1u+o7NTa9tZ4HfuxEpCiqLKs8J9isOM+nYa
747seRpS4+F51OjPmr+NYgDaQndkqR8zGbw7gW4o/6L41gWj46iKUzylz00UHtzBDH5l00i5jpKR
whBhyaHcNnoL5GB2W7UvSuz0Kx7S909tLtc48/Ub8L1gb6iNwaL1n1PsBa3+DqZ6+uWKYCqbxLRP
Z52t741fg6R5E7M6S1qCPkmREaFM12LZKvfZDebQgDceTYFwK/SeeDBFQhyFYMiFVcgQltOS+2q6
rRmKIgTPs2Gcnotal7/P3O97QUPONfPnnhJ/jzvJ1d0WLAToERmGKmf7ioShdtwaBqKxIfwMo5uL
Sf7uIbR9HCH6BzbeEmKpjy7geldJVCZ3o+NC7+zbyyysUvaHSr30SWAyea7C6ZfON1uwJdN21I5k
mF/OeFZowulnxct9d21D7cN8PvRT2WJjci8LAIC7VZtEL9+qVbUjAcg3QWwkHwQkpNxOlaeUV2xj
JzmP7ZaMKV4Az21lJus2B0jvK5ZVsekVaXsertOhimCtEguzb5uSUh9tJo3uz26EDgd0hufrRmh7
seZOx1XL46mUBTMtUBWiJQ+aXBQnnYvSe7JQu+ZWws1H/AshBzyVTBA58EG1Kkq3x3Br6eVcIreS
BTpFLtxKDU7vfpnHrLiEucKMyxsVNKa6+jXK2RSfRSwCiuDALT29nsndagG7njpyfd182f1X1tG6
Bl3CRBYmd6Bi2K4F67fLBTMgta1r/LDTqkkXCfRodYkHEecwXeyGRQ5P+3bHm5zmB/UY9ElqgRQM
BiRoBODXzomech1mxTE/onhcjlQfoYJvHs8FbVfcbzlA36ISZ3t0MIADYIeexNkH1jeGrYvtZX9B
fLJds36+ezQGkT/fWaH/91R4iPnAkmbkM0J1Na23YSUPXkeAm02Eh+S0iuGP3cW51X/kxsb+P3eH
i/2C96KxFnMbQ2KO1RRiXS1/Px56Hd4tfxlVijoVaQS4NRwOmYjkMG06iE3UQihvbu5r3UZ81AvY
vIEPViH/HiDNs50HfuE1T0p1pqpj6GE1R7d4kJjYwkrovrLnpc5kZpux7JNJJTeMisAXBC1OviDC
Xj9p+GIuJ8cjkeab2WMPP0SfCjUDiXdkEw2ICI/X7B/J9hieHmOfuPAgzC3waahzyV9dQH7dagOV
PMzwPm8lj0U69+Ak7FMf2OZiD2H25IiRTIjfpsVoJh5GGUp85l0V8AOqEsu4ON24N7ddiEGTmzMx
GnrEi0Oy/2lFxX2E1s07flyr+E7jx5CHtcZoDasSd79rjjdBmunSO3geKf2R2UFxRMN3d55zBZIe
kK78aDOE6vCYxXZUrBmxbAIpy/cTHWX72snLxlIhUs7WDQWRPUVGG0uKbJxEtXqPkVOkeMlKkkFM
vGFLyiwo63w9/Fcumbrk+8i/RxwKS3+A7cex4xJ3IlVAhHdnkM8tf6zQTqZuPU7WAk4g2jsAfwey
UBFmu6UbtyPLQys09+kw5r7MHvInu0D8vPmYmIRFcn23xtugvZwbhZNPf5I2phcM7SgtLlsiJhyK
IcTjVTdzc8um+1g4X9oQKb79TvJRz3bW37S5cJ/6Ny3CNdaA3It+M/eh/CkSsZw3v+xIq1v80hnE
BesuPEP+ys8XoV7NrWGEpr1eslFDlPBJ+XwABObqKcIvwgE5UcixlsA2kc/9hLyB+3p2fZDRVAOi
p0lAT24/F4DYoCCA6x+zwGzJJm3mfddU1zD9YBOonLah+mmLrD0nJQLrsThcBCU980dXePp+2yRC
1mZr1usGLesJbHFb6Yy1Yqdnj7r2FmC4Uavxfwp+WcuLjxZg2e3HDshP7/6CholK9QPHhdHmE6k4
3JvTDzTmWTUhSq9SWLZ1JzD3hakdkJR3Oa1RlAUGl0tawz7vjkm4PX6A/w4PN7fZOSS5eUBlw1XH
ERCsDpvFaVXH+BVO++YetmiYmNXoUj1rOjXgHaV3QFGII/b7HbVn+FcZViG+EFe/lwH6dRNpnpQ5
KhJO2fLpElhrWhP8zyL42FH5r8RQ1P7FO/nmErHYH7U+Pjk92qAVvzK53bX9DsdflsbIAvEIOPG4
IMypwGhsNazoOxN0UwNJJzorwS6RWV/9tmSsHCeFHhLt36VvDG0A2pH01GeXKNbA0EGWPwG2xX7O
HClMqKmMde0V/t5esEZY4CJz8GTNumGZr3uMBxnx4yDz0v31yQvY16FWM7dR1peDEql5Vc3jxMEA
VfEqmVdFIMVs/5l2Zx147z99APMMWsE4qQrzNpCqpa+Lwp77ee2rRu4CnJeYMIaLBF06Gx0her2S
5N0G10d3fTlR029YGw8scTjoBGtIgT2IwlBo+PqdgGnUjLOEMZlbUfX8T8O+MYf93rnjKYrA4aRE
SAHmU8gGGkG35rSZaOp60ms3Txt/HBE50LjfepOqqrHwl7pSlPvLCzh9xqgwLzaz/PbegE1OJzYF
Qe/XFsZWLkSy8ScDoSk0+MwlM+SLT8AbPmlLIr3dxz6LrOpuVQtaohaE1vVn5Q7ByyOGJ8kzuRwk
4a9b1gcb6MOccWvfYAtNnr2mUpU/OL+j7cKnT13aJcr4jxNDX6gU97CI1+bXuhTmrwZ/1o++FagH
ieUXkxJwsBvtdh/6zE/qBFqF0jkfz+HYzmXJx2Jrk8tkdnDDTepNa+ZEgD5GqzJkixf4520WntbG
FHyhPaNTCdc521Redh8tXP8eSmFWSbO0XlHVxexU9lbdbVNiMWZfnK+BjL9LgHGhUK4M0Ycw13op
m4rRyRNGp98nH/LDobrgtI5YmxcuCdBcBqOkdj1IUn304ulq/YS1mYrSOiN5/8WDb0lT8zLJYu+8
3iMwif/OtRwylSAZQp+lKygYVXiu2C9SA9F8V17LIfxKy1wbPguu1PfA3xUt53JRfv3Geme6pveM
o04Kwwu6BdTgYwgADhjWbHRTKjcfUtJvmWEkdDsfGxVFYFbOUGbyoTBA4gKvEZiAw9+sPLEmVqYk
/YsqGwNYrShWs+0eqKzLaefhBF7hYTFn4Vw+E1HnIPl8MWJupuvJTdV76vgrZFYAYk3pBfSIBfpx
Oe7rPEojRvPQ4elJX85Dw4s8R2cKW39ZKdnWJjyEuENMhVf/0qLOHdUlG8wsrETOk5haY2Fr938e
rBionQCJ9QO9TvMiDSdhrfvgSTdCXINHj21hdrPA848N5ZDBKtGyaRd5fC9FXbOIZOtuVEXmp30W
thTejI/Bzy96BAweD7jgb1e/wsJ3Nd+5mk0I8REeF7vm5xdnGWUnQ1RAF4WC9xMMcqImGOlR2K+E
V/ZxVVXFCeXP84d8bCuQRd8lPam+AwOCcvdRH4oY6r6i+LTJf8JwGadZuW0AUQjbRFidj+j0aeXN
to4UhAbL1jrKfBHpi9292JBeEoMxY1uBYAPBzwx4n5Ip483EIefZIitKBxBLmJjyBmdY4SrYQgfL
4jBaQYhHCsp63Fy9FJVBw+ImC7IB2QqX/9maJapNpS/j9G4oDA7QEQcxrKV2EoY1ZsNLwKUEZQCp
+Vzu9/pFvLXKXEW24hWYoDWKi0QYw/aAsXvqqGV8tfGoeJ7Icb0FuiBX6BBZTCKyF9Tb6CvBGLPu
AOEt72AsUyDu8QUzeWRBQsvALc1fhvagBUcb3C3gBfp/eZ8EDjGiUvnUN0qT6EmSq2Att9maCj+w
puOqoIrFD7IDhssoYGPpJqnoDdIk9GIYVPmqyohFqMJB71TqNU3tDqn/5wnvPWFr12v3cv2YWvte
IDPB7PWjVn8nIxYcHnmQEcQY8UB+w4FNOC6Bt1F95KA+JLiGOPmoXVFQ//GQAEOCKS5I5AEmg3ov
kmOrKN1Zdk6wTe66udej8uQEkvKfK/2bcQjZAxtzf/ctSuDpUxQYREnFn2DBdA6rNWxQZRQPhy7s
qT5yH+KlhpBr8FSWJUgoAHRMswj4i6MDm6VCOzdsh1iFWzLoB/WgqS3uSBumIcnVpBXWeJBPZpDP
UiN/zMtuCmFty3+xI4WhOx5z9o8DuVi2V0vJVv4KoYRLeEDKxvqmE6uWq09Xvz6UZKQrfT/I5Y3K
oNAQQtf8Xx3r74w4LAnUBZHY9dGnzD0hd+0MdLb1FSxf/JJEdfYPq9ILsgq1K9q0widNRvw/d/JF
JZzcGx71T2YE6vVMgh+giDrnw7etc3gIzg61X2Q72+YcBgjPBOpSwtbcuDOBZfG4KnyQ12VLjWSE
yjYRQ/oQiuRr1O3Z7aW7qT+N+aZiBLJX5PyTr8UfWAskSEbDbNQOGd0jXTo3q3rTiEeeGTzuEQ0p
0WXZuR7sC9dMYPJRZLByE7W+GtkX+4sL5d2wWlnS7o78mIasXs70+zdl2HF2NWWFsdy8yaFEn5H8
FxulhBcfpO55XsfwertwSUgs/E4GdAcmavPJJNAaqQJBN814+Oy0DgT2m7Q3ZDL34JHy0IRPCpDk
d/93JPt9AUCtOEBuIYBZULsgplJuntClbY9RVdZYkzvBRypY61ZcZzgWF1WbHiihAEhoaCDrgYZ3
i5JlEHw7ikF378CZw6QJvsio/JypfYs+Z0pDbk5e6KDAIYYftrx7ASZP0pIbS0FtpszUalN8HGz6
5hIKRBl4RopV0lPln3AmMVatj4PllWFmjZ03g+S8782XEi2uTTyIuVIsKbaOpYpZgnHWfFEgtapy
2JMf2+nv6TsGXMkslOGCYHizyyQC267n6dEDoZa9wqbWV04pDB3d5ZwP62RUXcfv9DM0B5mr08me
JwImfr5w/d5lFN7Pu2i/0sQeFVMjAnP3b/P9/khwCZk9UyTh7J0M0r8tyd3GxWpxL70N59wHZtoU
mEYI89/A18kU9MyCW+kNFmy3oy30hhl6HL8M2zE4InhCOBsAcrjh8WZWYVbNXTTfMUlAHZ8KmAzL
yzhJlENl6HGmPgDMVDwA9x1AM7Y0FozIYK0B0HOlPaKd5hXYsF3142iiPNuw8XRRQY0oi6NwUFVm
IJsH1S2s74XSUwPVKkDWPqQ94s/M/ySlTPgTBRNHxp5k0xQVo1WQlBdCGhtdYyZVyWsRa2IyuWv8
eB+75SpfQTI5XlgH3+HppGc50Yn2vgMC2+HMLrbj34YyY8dkY9bmFuFvwRCjDEe7gHvG/dMUVauz
ppK23S6j49+U2PRrBnJIr3KCraNMWZw1x07K3tj5Qsc43OXDENdGfXIlusK7JiBnxg+rowFlwoCC
ZqVRMNF+xJdsZMmaQpxYcWR/Cu3jessrfIMJry9OOw8yck5z0ukZs2MigX00LX9fYX9ttevkl9CG
ABxCR4y/t7TRIg9yOsPmSVx4+dstkWR0jZJmPr94odECYNP0sN+EF2OUCo9mSeYfU26gmkuTNQiT
j6LIbYu1Hpc6FsYZQKMLwgJEeSIb3rqx1YFgqHwanSP0aTC7ipxTqmlHjcOf3ljR/98yw1jtKgOK
IT9/QBmOcTKEdO54qYQ+P2FUreqMJdKS+v4tYsDqiSXqlSHFuvnm6NtrbhbSJ06HYlm2jK5OTrXg
TpornNx/CJBltFii2fXfjnO+uGPFQy4Z4K6G8ulkIkjldJFGnwuxvW9boyHyppdnZe8XjcoF+v53
cZ8GtzQ5Gud3ebWNAmzK/FleiXP0eNr4k562Pe5gmtvfzQZgQKv1DEjbBOB1IukTjzp2gFuTzI1D
cwgHlzQT7NBrkRAAnptmYNnRunutF6GVzb5TaylIif32fau5kNpyaSU6ZBmvF0Qc2x9HbGyZbgpS
7+WwFAOvy+maA25imOE8loL05+HSTZfYVFTe8R81Rld/UPB8SRWWMjlqT3GEkb2ZewYyzVxrCMS5
/zjBCAFqNuWvYO7G5ss0c9R/vc3k4NluHV8BDeLwejo5lUQ5E3RkL/fPP2R/KXjgp0z44X1bwESN
TNsMSqxMlNRpNoCA57+GwtphLILius+eMcfEbLdi1egbU5HX1QkqMF0t3M4FzRAmPamiW/Xy+frh
GkWr6pxV6wJh6YR+yMMmwO8JjRGiiXmAGROKcv6mn1oK5xOkARzGnpYv0JapF27AAzLNBJhiPqK+
BgJg/0AL5QpjmdKHsON8WAbCW89PL98NAJs4cp1khk1nclGt3Im3NJzJemr6iZGFda8Q48V1deG+
AhcI9T+HCCEkJ9XB0CT2PR0DjK+gjQT09N8zvimZUPToVv3DPUryDvF9pasJ6j+oIQ8gn0YTPqrF
NYQH3EO/BBaZKk9TCfnA0V7GYKTJqPYattczzjypcssLNoXzfoINFcLN/Ntf7EQgcdOZpGL99W8F
PDx5Bx6lqUp6YTsKSD5r90fnZEnZ3zDFyHvHRrvLI6iYZDRAu+syosDwEMSh0X58tuKROcLh+MtK
sH7KK7t0PHza2rxQZYQJBPh6OExkZ/L8NZktnq+WLESQM2LQGLHojY+9+ku24uZ8Zub4tDjdFxIK
XpWaoHdGg6xa1FlQ5W+b9rQ5nA+IslAHM/Hfed3crHoueroMCRyTeEN35pf/BB8dYjnohgzugtMI
JvSQG1SPtcH9noVPxczsmeWQtE1ZQ4P04+/uA888d1xJAs1lXZtanJAOp6oVaYMBj7Hjt04mmzQ1
ACI4eyPHF3j6i9d+4k/gv7S8CquDxrILLmhkXKHKaPQvqd80PEve3jLy0uVhOVcQOg/PJ3f0Mpi7
FJmH1G8lph4tuCGEKLTwG9SkSdc7jplkug8dmTL5O4R9+KNjcrO6SA5of5iYeDrovsAuGxGnTuYF
zn2mqTKW2uuLknUiU30gL361r0XHJ4W8Ldt553tNFw66LYPhqOBul+say0pj9Fjv4Nj2J2lcKVSx
ZG4BGiY8iEs5BLQbroGXlT257YyrJWH7QxRbCBx2UY53+OjgAQVNCR+pvutuG0w9RHlBuiJFTUK6
eo4vq7UBOKiKGkvRj2oNRbgsmerGrFCcKsKSeD4EYBw6ogcZZDnzzrrH53Abv7213K+1UzLZ2a6s
fU9ReRC/gK0hj4Barh8J/+4QpjN8AxbrsR1PnXf2scTT1AwXgcSumB8EZILGWyP6FABKLdmopQRO
CLiVoaoZH9LpjIw7sz1E4LxGO8A3PjBk7kAeaLxnqavAfqTXTyIYqx5a11AR0O1gfljdTrxvztRz
O0nfX20Zt16Gd5izDQ8DzpgdDaSS+mYAAHf/d7UwZv/H/Eof+dFF6WiYyB90MG+jlzxJCfviDve9
DcUOyVn8x6If5QJwGckdOZJhF+VR3FsGDQnsBC9OyLuMfObfCqnQHXUlMJBApDYISFdnFw6+q+YW
a1i4o0S5zyug3BPs7I5N7GHYLhx5VHj8mTYK9cGRGF38QTfNZGrjyKDk/eoK4ZzBrV/G5X4SzGgX
ACscc+BwUIj2CmDYsLwpIu8+mB8pVcUhacxywddQHN4u5NMf50r3V71Bu9p8Iu3hOpEMZkt93PWC
c0/DoywD1iaIrXf8YvG5itDpLnThBgnW8Q15Ibc9oVW2/uSJydLb2HRUOvHrkiJrJUf/0TYfrZXo
fhEXxPRf2tpXPRco8EbXrDigqanrHqENqkyNXEn7bKSx2WLKdBzyhribnMKoVtW3G+YG1mQWDJiX
GnEhnlty8ogrKxT5UImtfPd6T/F0qFeBss3+M1aKanLUkBOn6RmcduBSRVVPzvqhdkHWsHV7i7Qp
Rw9U3I7teLhyiBaWZR9O5XJAeTPanPG7UcIhKvVFIDh3qp3fThyfaPCzhK4x8gUY+ZHY+3QRlmYg
xRgvQhVwn+qNsdbnzFIPHYk8rW0C3BVOVNLNmFqhwp+Uyh9zlKFAZSaUjcex1CdU38CC57cKZc5C
UWR9iUMR3RH1kweKgnaMX5vxYdNBXXljPioMbpKD1HQIsrl6ErLcPzDpwsr+MbGkzL5Cfi8aSG6P
sSTesseZBbpiZdLKU4K1EGZ5MCo219Y4MmAaKymRMQlDHSEZ7xuX/+/WMeWM7IfV5CYR5NhY2Tkw
OGeuOx7yXbtGIBa+AL/0CotZEPvU0eib+eNqkG+64ezl6EHz3Dt8ErPKlazKx3RWwLMCMlTODXBH
4a3JpyjodEcHL/rFEGqKbCuVfH9Bd2w8WP2o3OGK//if7e93HZG2YADyh9JgvIpSsoq/RHvu63J5
yRJ4x/THki9lMEH1aInWjUfWPaYNodJz2LIxmpGHCGComBj3GgFdrXbwikTEnQE4f5OoNQDBECpS
gc2z32RR+Z/7k1xJVDuarnOYl84pxofCtdIToApPUqSnB9COvKDYuVuqYGjaNJ95bUuBg9qEOsxO
Ad+ErZpHbo/9ychlSVcetXjCaCXX0g/RKMKAmIPVd81K2h2wB2BCEd05QdjzGUg/8i+NAT3nD29/
ASp9VZ2Md5R9kulM1EyVX88QUWGGIGKh2IBlaTTOO/ls7jYixdxW8HZZNkKda68vbx/OYxH/lmge
Q3P5h7Ymr70wEHVhEds0a6y56alUa96UucMBZZvRVkEGnuwf/8hBlfKfcD5Z5W9UtFFDOki0svtz
OoVxjnIkIkG2JlPT744ViuQLWsCnbBdnAF4wVQzstbVst0vPFg2HiQjHiGwMLw3/3X08MyiF21Vz
FIFEirGp3zVtpU3D5qzxD/cqjpjSd8GHWh33jNrdn+CZ/RGOw29vk48iEK1zwiiICQZM+HeJ+R7U
Zb3S7Az80xQAD3ywhaV46rATbLglyy6LJfaXnT6srhZ97rbzGlFCnCFyE4uq8a2IXfccNiHkWnMf
Aw8RvpQpPqYaoZ+ek42muAtp6MDxPgWOrjznY5IZPzvtq9TrtMk8wFY6YhVAw5uLeUyJOuGHyMek
yNIQ+VzKehOOL0CSUHZq6s/zpiLt8URJWW3T28oA+fLT31kMSagwfJtltgJ4oUJpXPM7eZW4vknY
qfKtmXHnTSCG9EapWOjfXjFO2FPMIJKh615C/tROyj8eVLXkx+n8y4l4c0mpqq+hSC0SSUSzZmHw
vJpRyBJLEqEVx08j/mICBnT2A0Ez06cosT3jOIUOf8PmCljnXD+AVcDGXLKXfUYj/DXX7Mqo0rI5
9HHOoc5iB1B26G4VHDKAiLFGrgwwXz7iPYaiREGXYm9kBE/zNoe25BCP0fQijH3YPa80kLNaAW3k
y31hztKE54OPH7pVFeQCopr5hc2tOS0HfIuA0Qip2wXn8pP1JO0S+DVtSRMspxCDkF74wdPPFxOB
0E1lptb00+khqC2lIqoZx0vRwB2treyrjBvk8NEu2+QmeEJaSRVwjRNa6E/0l07nElflQEJHamUI
RC/oeoTrpl1nCv/1qznPN0CdStwspgn/SvGFjXvBSQSG2vd6empoFnKyubgqw7JFg3LqnLfJxz9Y
QsawYBcLJSilTN4lMfZt4GgsCpmZLyMYrLu/u0fI1lJjMYSOzO6qOIUhiSA6mT3SLu+Qz2Ep8hVM
DZ5R6Ye5ADZy65QIr59R7zfG3+WSkrI/yTgnhpATZpylBmyt1edL4cyNuhGBC4UIZ/+ZWyNAsi6U
m2xlt8catI17BB+yD1Ag7YLPa5Dy7TXCZaLy/qDixaPRs6cYep7E6ibQuJETEqjSOKsF1WqGwitF
k/v4mHNTyIOmqhY6hPg2wSZEnYnYfL9i8tAqvPojOkPGrj12WTZu23H28qGkIQxw5k5XjicRrOgm
MACKXkMmEeMaEWEt0rSGmucxHFK+lUsdOEG/AvsqNL9R5AwdC1BSZI+hwOpLSjWE2dZX0t6t2NmA
RhM3fJObI8xNHZNCCyZHcrBWL/16DH6BSUUoZ/eeq83rbyuoJOMdp452jQG6cz5RrCE5fKyyAN9F
OOUY4yEkNUljaQolRj6skdEgXA5BEX5RpRkTjkyDrpfE4SgWSzbJfLMBHEg0sNfS+2UGNL9bI05M
5iNrKYpc9Jw7FjfoqeCgFwOmLgw7PHsZ3/vlpepxW9tgtZSg+6JJBMN1DjLudSzWe7X7WQH7OOxo
V+1Awrhcotxn8C/jdYejSHbr3H2tXZZePwo1mGOUuYzE+cn2rB/RsVBB5pHXCaI7TRLymVcHeeqn
RYylhx3XT07N7hTN2Nn9+C0waHmCFxAHJ154wCMq/W4BT5uAVAQz+Bz8Qccqw+OGZQayQVQCZzR/
Gnk3sD+Konb1FaoNJu3rOf8v5m2gjUXOby3KxaiLh5sFp+n8N9yRaVSYiUECl3BOWg/KTRnbG6kp
0xAHdtFXEvFelFb6FE0dMLb7MsPHBw8l/Cdft0fu0S3YcOUJL3MKga7OnyVcrRQnlzIiPUidN7DK
KKRUbC7OztfM91HUUhk965UQ1u5WKRJGe4Wl+Wp/q/PBpNNJFFAA/F3rJtxMcfWcM4rRs+IpDyq6
tyXwX7s19sGBOT/rr5lstzPaCskrGrc/WcxhQRNFXFXAGuBlQhX1rugXRn+tGqn5ZaJf66sH/EI0
xCsEoV/Z/1ENt9Jv5I/wefImAzCYUD3TVusaAhM2jYQ5LMeqcFock3/4J2SD51HWVM/ZfdHxxLwr
LvISs/sURp9JrKzjltXkHjb9ChK92bk3QbySdFwGy9Pi57IHgH/OY0CpZbVoPBBelodFCq+qxzAk
Th8JuXiKwqSOV3FXQW20PfTby8JD3554hZITY8KOAdi/ae3ASKXukMEp7rcyOZa59Vn1/IMeARe9
rZHX8S3TV3nMn1PcdxaLff2mKQ9Sazg9I6trgACpRxvX6r4dQJqF2QPzGY3wFWOFWUFyo5Apof9q
JfbXcNjQlql8M/J6/pb7fyKhbwD75hYazwmTibcAQqua5E7W327ncWF9kUQIu41juQ6r36h3Ylcp
eXvukQYoAlW9UhaXIF+TNlArU9gZByoC3bSDQOiDdvrpOan0m8yDJbdfhcrz6izt/fNFzfm7hGuk
OpPLGTH5Zl8ZBhxR31txE0C+mqeDLsME7FzY1BZn8YvRkWVwlBYwVt6AEdQ56behn3nPO4fcJT6c
XCWF0LaLycVagYssgzLQFbZtnc/nKgLsOn8edsAG2ezpJ40UlqakRb9HdWGH17/L0yiRj4YXg9vs
ghBRRD1Vx0qimqVZJLH2VB5sLHeOPNGdRRPtXwjH3vJb+GAphmn1vpj3yrJTkb76xItIEDuKw2vt
8FVe0eGRTMvWNxJIuNxUFb+D7TkLzGPehQotBqgBx1z2GqR/g8mf9MZlexhj6n3cn2dusWIXxwOr
cXqaoHCHRSKSwvrMuLhi/zN7uFu04lXKImexH9yh7fT6SW1AWsSqszSUvGUxxxOXfKVrIKKIBWY3
8qeRcoNMVbFcAscuZcRBPQd+1Wz1zTOHmXxfu2a0zpnz5I0pd7FaOrSemrnJCAJwxKlMxqCOSAch
L8rG1WsSDJaIhNrTAZyBESYD4x4Oi3hrXVMw12GhkWlqUMRyP99GTlOb0BKXCvfiBd9l8/7hXjpM
OX0LikkkP7j9vT1Mo6QBzvF5aLySoYzqYAiz5RG03OwvtDmYOkXef+bnlip8B+gqtGSAvek/dtdw
E4/k4Em/luR2ieB/hnMCYgfYxfRjWDHu872J5j0d5tyZ2uR7g3Hi4gGV6ZAPNXV2CHMYS3UGXpE0
hwUe6UVGTN0L+x9fGc8Hq74PohFIkZ+C7wxej1NJOkYAtlPZO72r6DjDiVzMCdA/LdTiPImzIjpg
r52pXenZQLMpy35KU0EzuPg6bNK1bNe0UF3ct2AINn0McRmq3TrbbKNyz1LWAiICZEzUKRDZKWpr
/iMv8c7sreck2m2GG40BPXHPHeOAtN8ZVjhVNnXEhJsHdE6Uty/xCR4bI/zWoocL09vEb0moAYGb
ksPeyQwL5DRtXenhgC+5wIib6qtF8xOJKCO81gjFVZNqMZir9DpGAzf3c+1aSwM2SVCOW/BpEBnW
WiJZPecOBGc3bTIn5WsDBN+kUwqmSLCIs8xbZOg/f5wXs3jQ+9i/22Cu4N9lai7VgBV8PzK7miJa
wfirC17YxQo5WVVmk/bZNtKDuT8CX0W2MsEzkpKRLzXTQ8owpVzHYD0TdCb599FoQLaskYW2eR8F
EgxA/CIh52DMvhufYRXVmEZ6YkMPSEaLHnsVnHz8fjI2i5c8TZCZgVDOPjx16nlw3uBaHGa4Wgyr
U/I8pfAXpykN90mwJrzLZQmoptDYFp/QoNKgMCaD2SSkMaNTph8xT8JcMOOtLS6/W7M/Ek6VBuv9
tY+W9ffFxmsPuIccWZia31DKRVBVDAR+vrhuPP3NPSuwbUFSWwuSs+jSkDjXbfLwF8m2pm5PPfe3
+XrihhjDIf28rDRf/I3qcSIPTbVEt6/t30EaVEbUGKKn57AT4sqxdb7T8YZPl6Q9OSv6epigzKei
v+0hsIObbQRskAz+az/D0OLbrkN2tPSCa8u8A96Nywo7ns7qh6Gdm5s/7u0Ml9RQ1M7GgUzFvXaP
YFCxFqf8t4eEEdei4sdtBFEV5fDj10qoew6oHvtAxKwjKXCIGoiPKK/5koP4yyxjwSDDD9kCuF3g
NtSE4iaWSIBnIZtr1m5TqBawPLJ7UTJcAbUJOXxWFbKTF/ngYbMehg0IRlfXJ2/WSDg5pZgmjlrp
9BAoOq4DDybg242Zf9nTM9CnyxJ9mr4Hjhw86EuJLTc2O59gYUwAPT5SGkoTCUn/kweUJ+wFhs9q
kAgIDuoee2yWcS4VCt6to/hkcXUGTw+grk1Zp71ZIeUPTk/oaKB1CzTr+ihQz/1+GIM24W5qQ4dF
ufJ3uxHIvFa1LE3j5lu4DHQBD4tOYtRyochapcrYHlFWUQ0eqwtx+eDl7/b2cN+vxbTlfXdVnCi3
tN3waoMiH8IPepePG4WsQD8X4Fx3kByzJ/b4Aip7Kf2KxCzlYLTk6FRfNMeM6GDN8G6m8ReqbTJZ
/UGn0BZB7t02/47MSHInGX8DO/hnyMRUWRIzNS55u4kbrDKER/ySUhFKqLyrnr/Ez/oI2/6oY2Vv
PcHpQ1Dmh0NM/hgMLQ==
`protect end_protected

