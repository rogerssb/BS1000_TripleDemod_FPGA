--  Module : ldpc_encoder_pkg.vhd
--
--  Description :
--    This package defines constants and types used by the low-density parity
--  check (LDPC) encoder.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ldpc_encoder_pkg_1k_12 is

  -- constants
  constant C_ASM_LENGTH : natural := 64;     -- attached sync marker length
  constant C_LC_k       : natural := 1024;    -- k = information block size
  constant C_UC_K       : natural := 2;       -- rate = K/(K+2)

                                              -- n = code block size
  constant C_LC_n       : natural := (C_LC_k * (C_UC_K + 2)) / C_UC_K;
                                              -- M = submatrix size
  constant C_UC_M       : natural := C_LC_k / C_UC_K;
                                              -- m = circulant size
  constant C_LC_m       : natural := C_UC_M / 4;

  constant C_SHIFT_REGS : natural := 2 * C_UC_M / C_LC_m;
  constant C_CIRC_ROWS  : natural := C_LC_k / C_LC_m;

  --subtype asm_t is std_logic_vector(0 to C_ASM_LENGTH - 1);

  -- hard-coded attached sync marker for length = 256
  --constant C_ASM : asm_t :=
  --(
  --  x"FCB88938D8D76A4F_FCB88938D8D76A4F_034776C7272895B0_FCB88938D8D76A4F"
  --);

  subtype circulant_row_t is std_logic_vector(0 to C_SHIFT_REGS * C_LC_m - 1);
  type circulant_matrix_t is array (0 to C_CIRC_ROWS - 1) of circulant_row_t;

  -- hard-coded generator matrix for (n, k) = (2048, 1024) code
  constant C_G : circulant_matrix_t :=
  (
   "1100111110100111100101001111010010011111101001011010000011011000100010111011001100011101100011111100101001111110101010001011101110100111101011100111111011101000101001101000010110000000111000111110100100100010111110011110000100110011010110011011001010000100100100011111011100101010111010001111001011010110101111110111100000110000101000011111100000111011001111001101101111010100011000111100111010010101110000001110110000011111011000001001001101110000110101111110011110010001110010000111000000100010100111000001111001110001111011110011111111011111011000001110001010000111100001000111100010010011010011011011001010000101110111101100100111011100000011101001010111000001000000110000000010001011011010111100110111010010110110101111100001011100101011100111001100100010000100001000001100100110111011101000001111000001111110111010010101101111110111010001010110110010110111011011001100011111111001111111001000111011101000001011101101000011111110000011110001100111101111011010000111110110101011101110010001101010111011110100111001100010",
   "0101011001010000100000110111100000001100101010001001101011001010101001110000110011001111101101001010100010001000101011100011010100010010000100001111101011010000111011001001011000000010110011001000110010010110101100001010100001101101001110011001011010100011110000001011000001111111110111011010011100110100010101001100001001010010100101011111011100101011110101010000000001001110100000001010110011001111100101110011111111000011000000100110000111001001100100000101001001011010101000001100101110100000000001101011110110011111000001111001111100001001101001000000010111110111111110000111101011011001100001000010100100001001011011110010101001111110111010111000110010011011000100111011100001001100000001101110010000101000010000111010010001110110100010011010100111000101001010001101101010101010000110100001011101011111010110011000110111001111110110111010110101000010011011001010010000111010110101000111100100011011101001111000001100100110111001110101111100111000111010110110111011010000100110100100010100110000001110100110010000100101",
   "0100100011110100001000000011001110110111101110011010000001010001010010011101110010000011100111001001000000101001000111101001100010011011001011001110101111100101000010100111110000101100001001100100111111000110111001111101011001110100000001100011010110001001111101011011011011011110101011101011111101110010000100000110101110101001111001100110011101100101011001001100000101110001001101000110110101011001010101000101010110001101001000110101000110010001010100001010101011111000100011010111000000001000111001100011010000011111101010010110001011111011101010111000011001001010010111111000011001111100100111010110110011110100111000001000011110101010010111010111101010100110011101001011101001001011000111011000110011010111101011101001000110000110111100011101001110110010001110110000010001111111000100010010011110010001111011101001011110110110001111111011011110110101100011111111001110111001010011101001010110010011101111100011100110100110001101100101110001100110101110000111011110101101001100010110100101100101101001110010111101011011",
   "0001101101011000111110001000111001001001110000000000110111000110101100110101100001010101101111111111001000101000101000001000100001011100100011101101010001111011011000011110111011000110011010110101000000000100111110110110111001100101110010111110110011110011011101110111100010011001100110001111111010000000100100100101111000000010001101111111010101110000111000000100110001011111010110111110110101100111011101100110000111101011011111111100001110000010010110101011010111010101110110010110100011000000100000001000110000101011110110111000001010001011000110010101100100111111010000010110011100011011100011010000110101000001110111110001001101101100110010110100011101010101001111001001101100111111000011101010000000010110110011000001010101010100110000110101111001101010011111011001011101011000011111111110101010010001110100100000100110001110000100100110111010100111001111001100011110000110010110001010011010101101111000011001011100010001001000001000000110000110110010101001010111000111010000010111101000010101011010010000110001000101",
   "1011111010011100000101101001110110001000100100110011100111011001011001010100110010010111011010101000010111001111110110011111011101000111110001000001010010001110001110110100011100010010110110101010001110111010110100011010110101110001100001110011110100111010000111001101011000110000110000110100001011000101111010111011100100011000001110101101111010011011111011110010100101001110100011100111000000010100110000000111011110100101111110010110111101110101101111100101011001101100100001100110100101100100110100000001110011100111001010101100010000111010001101011010110100100001011001100111001011101011101100110010010110011011011101111111100110111011000110001101101010001011000010010001100101001111101000011111000011101000011101101010000010000000110010011101011010100011100111111000000010011011000101101000101000111101100010001110100011101001001111011001100101011100111001010010001100101100001011011100001011000111110011111010010001001010001101100011111101100010100010100110011010001101010001101100001110011000110010101111100101101111",
   "1101010101111101101110110010010010101110001001111010110010100001011100010110111110001110101000011011100010101010000100001000011001111011011101111001011011110100101010000110111100011111110101010100110001110101011101101010110100000001110001101000100101010011111001110101101111100111100110010000001001000100100000100011011010001111000001101001011001011000111101111010101010101111101100001001011101011111001110101111011110010101111001111000110100100101010110000111000111000111000110110100111101001011011101111111011001100101110011011001110000110101100110111011001010101000001011010101001101010011111000000000011100010110011010111101110101000001001011000101010001000111001100010100110110110000001001111011000100001011000100110000000001110001101011010000001110011000110100011101111000011001101111000111101001101011101111001111011010100000111111110000001000011010101010111111000100101001001000001010010101011000101110101110110101001000010010101111100010011110001010011101010011011011110000010111000011001110111100011101001101101001",
   "0100110000110011000010110010110100010001111000010101101101011100101100111000000101011110000010010110000001010011001110001010011001110101111000111101000110100011010101000001111000001110001010000100111101100101010101101101011010001101001111001000101010011110111001011011101100111011001010010111110110110110001011001101001010010000011111110000100110011001011010010110011110100000111101001111111100110011101011101110111000101100100010100100101001010010111111001100111101011100001110011101001101010101110000111001110001011111111001011111000010011010101110100110101111001100111000000010101001110011010000000001111001011111100001111110101011000010110101110101011100000010111101001111010101110110011100001101111110100111000010110001110000000000001011110101001000111110111010100110110011100001110011100010111000000101110101000010000011001011100001100111111011000000000101100110101110001110010100111010100110011101111110011000000000011010000111000011001100000101100011011101000100010110101000001010111001110010011110001011101110111001",
   "0100110011110000101100001100011110010010110111011000111111011011001111101100111010101110011011110010101101111111011001100011110100010000011010100001110000101001011011100100011111000001010011000001010010011000101100000100010111010101011111011110111110110101100101101000111101101101100011000111100100000010011000111100001101010011110011110011000001111110111110010000110000011111001000010110011011100110101101100011001011110110011000010100111001011000001001100111111011110000100101101100001101110111000110001010001100111101010001101110010111010001000011101001100100111110101101101101111110000001010100011000111110001000010111101101101000011011011011111111010100011000111111010100100010111011100011101001110111011011111011010100101011000000111101001111010111101011100010011011110011000110010011010010000110100110010111011011001101111001101010111110001011100100110111000010000111110001000010011111111100101110110000001100111001111011010111010100000010010111001111010001001111101100111101110001001110110000000111000110111100010000"
	);
  
  -- functions


end ldpc_encoder_pkg_1k_12;
