--  Module : ldpc_encoder_pkg.vhd
--
--  Description :
--    This package defines constants and types used by the low-density parity
--  check (LDPC) encoder.
--
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ldpc_encoder_pkg_4k_12 is

  -- constants
  constant C_ASM_LENGTH : natural := 256;     -- attached sync marker length
  constant C_LC_k       : natural := 4096;    -- k = information block size
  constant C_UC_K       : natural := 2;       -- rate = K/(K+2)

                                              -- n = code block size
  constant C_LC_n       : natural := (C_LC_k * (C_UC_K + 2)) / C_UC_K;
                                              -- M = submatrix size
  constant C_UC_M       : natural := C_LC_k / C_UC_K;
                                              -- m = circulant size
  constant C_LC_m       : natural := C_UC_M / 4;

  constant C_SHIFT_REGS : natural := 2 * C_UC_M / C_LC_m;
  constant C_CIRC_ROWS  : natural := C_LC_k / C_LC_m;

  --subtype asm_t is std_logic_vector(0 to C_ASM_LENGTH - 1);

  -- hard-coded attached sync marker for length = 256
  --constant C_ASM : asm_t :=
  --(
  --  x"FCB88938D8D76A4F_FCB88938D8D76A4F_034776C7272895B0_FCB88938D8D76A4F"
  --);

  subtype circulant_row_t is std_logic_vector(0 to C_SHIFT_REGS * C_LC_m - 1);
  type circulant_matrix_t is array (0 to C_CIRC_ROWS - 1) of circulant_row_t;

  -- hard-coded generator matrix for (n, k) = (8192, 4096) code
  constant C_G : circulant_matrix_t :=
  (  
  "0110000101101101101101011000001100000000011011011011100110011001010101000111100000001100110101101101111111001001100100001000011101110010110110000010011000001101001110010000101100011101010001100010101010001111011000101101111010001000000010010010000101100001100101001011111000000101001100011110111001000000100010101110101011110010011111110101000011110011101011010111000110000110010110101100011110010001000011101110111110001000001001001010100001011000110010100111101100010011111111001000010000111101101011111011000110111010001111100000101100000001000010000110000011010000100100000110011010101000011000110010111000101011001001110011110110101011110111111001000011000010011011111100110111011001100010011100001010000011000110000111010011101010011111111011101000100011110110010100000010100010100101000001000100011100000110110000110000011100111101100010111101010110101000110111011010111001010011001111011001001111101001011001010010111001100001111011000110010010001001101110010100100101011100000100110101111111001010111100011001101110001000100110110001100111000111000010001010100101100110101100000001100010010010010000010110010110111010110001010100110110110010011111011001101010111001111001100111000010010010001001111110101101001011000001001100011110001010011110110101100100101000100101110010110000101011011100100010001101000001001100010111101100100011111110110011010111111101111000101100111000001001011110011000100110100001011000110011111010101000001101111001110111011101110010110011101000100000100010110001111010101000111001011000101000101000000001001000111011000111000100001001101110001010101001001100110110011011010000011001111101001001101101111001010001001101100010111010100000101110101001000101101110101111010001001000101001010100100001101100011011000001000100010001011001101100110010010101111000010111110011111100111110001001000001100110011011001001000110000000010101000111100100110010101010100111111101001001101010010111011100010001101011111000001101011011011010100100000111111011111010111100111000111101000001001101100100001011110111000000101111010100110010010010101111110101011101011000101111010011001100001001010001111111110101110000001111110110010101110111100000111110101011000001100001111100001100100100101100101001011011110010010111111110010111011000010001100010101101100001001110000001100110001110100011101111110001101101001111000001111101000111001100110011000010110111111001111000001001110101010000011010110000011100111101111011011000011111001100000001100101001111001001010001001111110001111101010000111000001000100011110000001101111100111110101101100111111001100010101011100001001111111000110101000000000000001101011000010110111010000001010000000100010101001001010111110110111010010110100111000100011100111011000001011001001110000110111101011101110110111100110000100101111101000000000000101110101100010011001011010111001110101001100001000001010011011000010100110100011011110101010111011110101111111111100001110101111101111100101110011101001001000110011010100100000100101101000110000000111000001010000110101101101000011000110100101000000100110111011010100110011100011000111010110000111110110110101110110111101110011010110100101010001000010011001000000001000001010001000100000111011111110110101111010100001001001011011011110101101101010111100011000001000111010000000001110110101101111000000110010011000011110111010101011110101110110111001011000100000111101101000101110101000110010100011101101100001001010111110000110001110000110001010110011011111100110001111110101101101000100111010101011111000110111000101000100011101100100010110101101010010000101000101010100010100100001110001001010100110011000111001111000111010110011001101010110110011111000110100000000111110001000010100001101011111011001111100001000010001111110011001000010110111011110000010011100001101101101101111001100001001101001001110111011011001000111110001110100000111010110000111011110111000011000101101111100001101011011001000111010011000110110000101110110101001100101100000100001001100011011100011000011001101111111000000011110011100001010011111011101010001101010111000010010001110000000101110110010101000101110000101001111110",	
"0101111001100011100000011010011100011000110000001010100000010111111110000001000000011110110011011100110110111111100000100101111001110011001011100100001101010110110011101100010000101100001000100010110110111100010001110110101111010111000001001000001101111100001110000010101101111111101111110010100000101011011100111001111011011100001000101011010111101110101000101001000010011111000011101011001110101100101110011110010000011111111000101010110001111001000100010011000010100011011010101001110010111111110000011101100111010100111110001101111000101000111110100111011111110011011111100100101001101011010110101000001010100101100011001110100100010111110010100111010011001000001110010111111010011101101110001110110111001011001010111111011001011101101110010001100101010100010001010111011100000111111111101000011101101101111111111000000100101101010010111001100101000110011011011111010001111001101000000000000100010100111100100111111001110000001000100100100111011011001111101001001100010001001100000001111010011100111010011000011100000011011101001111111010101101000000000001001111111101100001100001110101100111110101111100111001101001110100110110001101011110110011000110001001100110111010000110001011010000100010110110001100000111011110110100010111010011000010011000001100000110111010100111010000010101100111011010111010100010001001100011111001011000011100000101111010100101101010111110010110001011011111111101010000011000011000101011100111101100000111010000111100011011110101000111110011010110110010110100001001110011100111000010010011110111111111100111101011001111111101101101011001001100100011101000111110010100101111101010101111100010100000001100111111011100111111001111101100100110101011000111001100110000000001110011110000100101111000000011000100111101110010110111010111100110110001010010011000011111000101011101100000101010111110100110011001011111011100111010010010110100110110100100111001011101000101100100100011101010101100000101000111101101111010111001100001010111110000010011110000101111000000011001111111001011101110100100111110011101111100101110000110011100111011111111000100010100011111010111100100101100000101001010101000101110001000010001110000111011100110111001010010110010110010011111001001001111010010011011000010110001111011010110111000100000000011001000100011010111010000111111010110101100000111101110001010000011110000111010000010101100011110011011100111110001111101001001011010111101111001110100101000101010101001011001000110101100111100101111010100100110111110110010010001000001001110100101100010110100100101011111100100011001000001011111010110010110110110001111000101000110100110111100101010011100110001010000010000011100010100001111000111111011010001111001110011110010011010000000010100000011101011011000010110111010001011000000110001101101000000011101001011010111001110011111001100010010100100110001010111100100100110101001111101010111001000110110110110010101100001011100110000001011100010101001101101001011111111101001101011011100110110010111101111101101100100000000011011000011001110010111011010101100110000000000010001101000011010010011110101010110111110100001111011100110011000110111000110110000111010100110110001001110000111100001011100101100001011000101110101110110100000000110110010110111001101110110101110001100110111101010110110010110101100010100101000011110110000101011011001010110001010011000101110010100001001011110101000101111000001100111000100001000001011010111000010101010001000111100001001100111110100011111001000010101110001011001001000111001101011101011010000000001100001101101111100001010101100101000010001100010010111011100011010111010111101000101111011111011111110111110001001101011111011011001100010111011001110110110100101110111011001001010011011111000001011001001010000000011100111001011111100010100110010110101001110001010011111011000011110000000000110101100101111010011101001000100010010101000010110001011101101110100111100001010010001110000011101011001001011101110011010110111110111000110110100100001101110001111011010110100101000011000010010110101011001111100100010101010010011001101100000100101111010111111011111110001111011011100111000000001010110100101",
"0010010101000101001101100111000001100100011111010010001111000101111001000100010110100111000001011001010100111111001110111111010010100101101011110000001011100111101111000100011011001001011010011100100000010100000111011000011110000010111100010111000111001001110011111111011111101011101100100000100101000101110111100101110100110110001110101101001101101101001110111101010110100000101110100000100000011100000001111001110011011101000001001011011011100101100101101000000110000111110010001010011001100101001101000100101000100011111010011011000110001001011110100110111111011111010000100111101101011110100100010000101010101000110101110001111110011100110001100011010100010100011101001011110001000101011000111100001000001111110100111000100101010011001010010101110100111011101000010101111001111101000100000001000001010000001110110111101110100001110000010100100000100101000111011011100010101000100010101100011001001110011010101111100011000001110011000000010101101110010011101110111100011100100100100111111111101100010000001100001101011101010101110001010000001001011010010100100000111101100111100011001101000010100111111010111111010001011101111101000000110001101001000011101101110010011111001111100000110010110010001101111111111110100011011000100101100000110010110101010110111110010010111110001001111011011010011100110000100110111100101111101101110011000110110101001100100101000011010110111110001110111001111101111111011010100110001000000100101011100110101010111010011100000000101010111000101111111011011110101001011001100011010110101101101110001011110010001010110110110011001010010100000101010000011011110110011111010111010100100001010110010111100101010100011011001100010000111000010000101000001101111111001011100000000011010110100101111011001000011011101011100111001101100011001000000100011100110111001011110011001100111011000011011100110010111011111001001111101110100011001001010000011000111000100101110010100101011101000100111000000111110001000101111110011011000101100001111000100111011110111100111011001110001110001000101110011011100001001010101011101100010011011010001101111111111000100111011111000111001011001011010111001011000110111110100100101010110100110111001110000110011101000000001111100100011010110011010100110101000101011001011010000111101011011100011110011100001110011101111011110111000000000101110000011111000100011111000111001011110101011111100010000111011111011010011001101010101011000001010101101110111100100111101110111000100100111111010111110001000100110010001100110110110101010010111010001010111010110110000011101010110011111001101111101011001111001111110100100000010011011001001011011111101001001001011011011010111101010110010000100111001011100011111111101100010100011100111001010011110010001111001011011111011010101100101100011001000111100110000011100001010011001101111010100010100011111101010111101101000011101011111000001001011001110010111011010001000110100011111101100100011001101111111000111010100101100111101001001110110010000011100100000011000000110000010110011010111000000000110111011000001100010000001010101001111100110011101100101001010000111110010011100110111001010110100100101000111001111111111011100011001100110011101000110110111111110011111011100111010110011000011101000100110011110111110000101001100011111110111100111110101011001100011111001100110000001111001101101101110010111010011011011000011110111101110101000100000100001000000100010110001110100110010111100010011111001001010110001010111101111001110000110011101010011000101110000001100000010100000000010101111001110111111110000010111011110101000100100000111110111101101010110101010000001000100100111011010001111011111010110110100011001100001101111111001000111000001101011100100100011111010111010011011011010110101110100110111100001010010111100110100011111110101110110110111001101010001011110010010001111110101101011100111101010111011010000100110100000111011100000010010010010100011000000111100010001101111111011100010010100001001000011000011001010010101111111000100000011011010010111011000001100011000010001110111110000110010010000100111001110000011100001010101011001100011100101101001110010111011111001111010111010000",  
	"0110001000110000110111101111000110101100110101000100001001011111011110110001010101011010001010100010100001011100101100101010001100101100101110011101010001101101101000001001101100101000000101100111100000100110111001110111101011101011110110000101111100001100010000010110010110010101111000010011011000011000010010000100000101000101000111110101101100111110000111110001011111010000001011000011110110110011001011000010101011110101000000001001000111010110001101110110010000000110110110001100101101111000101010011110001111010011101100011001100100010001101011001100010001010000011001111001111010101110001001011011000011110010100100001111111100110111001000110000000011110001101001001011110010010001101001000011110010110111100111011011001001110000000100110011110101000001110111000100100101110000111100010100001000001110011100011100000011111000000101101110111110010011100011000011110000010111111100001111110010111011011011101001001000001110110110000101001111101010111101101101001011011100011001111001001010111111100001110000100110001010101110010100110000101110010111011101111001111000110010010111010010101101011011110100001000111100110101011010110010100000000111101100100101000010000010101010111100111111111010000011101111101100001100011101010001111010101011001101001111010110001011111010001001000111011011000011100001011001010110111101011001100110001110010011011010000001100000011110011101011011010001001011101010100111101011011011110000101011010000101110000111011000001011010111101001011001001100010010101110111001101000010110111101111101001101010000101100010011101101000100110110000010100000000111000111100110100111011101100100001101110011011001101101110001001110100000010111111101100011000010000110101010010111100110111001101101100011011010010010011010010111000011101100110100111110011000101001001110010111101000001000100101000100111111000011011010001000000000001000110101110001100101101111111100101000011101110000101100111001001010101100100001110100010100011010110111011110001111011010000000011001101000000010111000101011000111010100101000010101110110000011111110111101100110101110000110000110101010011001111100011101101000101001110110110101011000010111011111101011011100100011101011011001010101011010101101100001000001110111101010100111110100010010101100101101000010101101100000000101100001010000101011011010110110100111110001100000110011010001110100111110101101111010110000010000000000110011100100110110011111001110111101011000101010110110010110111001010111111100111110100100111101110100100010100100011000000011110010110101001011010111100111011111010000100110001111111011101011111000101101111110100100110101001101100001101110110010110000011111101110111010010101011001011111101101011000100110000101010111100001111101010011101110100001101110010111100001001010100011010001100101011010000011100011011100100001010101010001001001110000000010001001110001010011010100100001011001100011011011111011111010110100110110011110010100001010100111101010110000111101110010110010011110001001000110100111000000000101101000101010110110000111010000100111111001101011100000110010011011110110101100111100101000100010010111000111101100101010100111101010101111111111110111011101101111000001001100001011010100110100001010010001011110000100100010110000001010011001000101111011101010011000111111111101011011101111001000111000100100000000011010100110101101000001011111110110011110001100011000010100010110001110111101100010010111001001011011000000110100111101000001111001010001011010101110111001100000110110110011111000000010000010001111101011011000100100010011011000011011010001000101001100110001011101110000101011000110010100111101011101010101011100001110011000101100010110101001110001010010010111110001001100111100010000001011000010111100010000001101011100000110011101010111011111110010001010001100000001101110001101111000110011110101000001110110010000100111000001010110100011000010010011101100001001111001110100100010011100111001101010101000010100101100110011000110110111000011100111011001100011011111111110011011011101111111111111101001101101110001001100010100010000001101110001110010110000110100101010011011101010001111011010",
	"1010110001011111100001100110110111010111010111001101010011000010110101011001010110011010110000110111110111100100111000011110100001110000001100010011101001011011001010010000001011110010001101001100110110010011100111111110001110011111001100011111111010111111100010110100011011011010110010010000011011100011111010111010100111000011101001110100110111100100011011100111101010010001010000001101001101110001011001100110011110111011000111101100001000101010100001111101010111111000110100000100100010111101110001011011101001010111101101100000001001000011001001111100110111011111111100110010100101101011111001100101000010001100010010000000010001011011011100011111101001010001100100010101011011111000110000010010010111110100111000111011011100110101011001010111011011110011001011000110001110111100010110001000100100001000110001001110100010110011111110011111001011010001001010101001111010001111001101011011011011111100111100101001011011000001011111111101100011101000110100000111011001000000011011111010000100011101000101100001011101011111110011000100010110101110100000101101011001110010100101111001111010001010000010100011010110011011001000110010100011000111100110101110011000011111100001111110101111100000010011011010110010010011010000110000001100000101010010000110010110010111001100100000000000001100111001100010011101000001011110110011111110001100111111010100101010011001001011100111111100101011011010000000001000010110101011110111011100110011100001011011100100110011011111100001011101000011110101000011111111011001011001010010100000101100111101011010111001110001101100001100101011111110101101001101101000111110000010111001010111110001001101000001011001100111110001010001100111111011100111111000100111010111110011101100011100010001111001010111010010000101111100000100101010010110010111001101110010000011001011001011111011000000101111100001101100101010001111100010001110110101111010101111010011000101110110101101100001110110011111100000010101001011001000100010010110100110000010111000100010111110000111011011011010100011010111100000101110101110101100100011011110100010000001101011110001110010000110110010010100101101010100101110101000011111100011100011000100010010000000111101111111110000101011101000110101100101101111010001100110000110000001010101011100000001101000111100011111111110101100101101110111101101110100101101010101111100001110111011101001101010001010111100010101101010100100010101011101100111011111010111101101001000101011010010100100000111100100100111000101110110111101101011001000101110100010101001001011110110111010011000011000111100100111100001011011011001000100011011011000100000100111100000011011101111111001101010110010111011101110100010001000010100111011110101101011101010101110011101011101100110010001010100011101101011001011000001011010111000110100010100111000011010111000111111001110101000010100011000100010000011010110010010001010111001000101001101001111110011001011111110000001011011011110011000011110100010010100010110101100111101001111001000100110000011101011100001011101101101111111010000010000110100100110100100010100110101100110110100001000101110000111100000000111001100001000100110011011110010101101101000101001000011001000111111100010010011000111010111101010100011011110110001110010111101011100001101110000101111111011101001000101011001001000110010011100100000011110101010011000010010000101111001010100010101000010100000110111001001000110000111000001001010000110100010100100110111011110001111111001110101101010011001111111011100111001110111111010000010000011010000100100000101111011110111101011000111001010100110100000101111001001001000011110100110111000001111111000000011111101000010110110010100111111011110000111000001001111111001010110001101111101100001000100010010110110110100101000100111101010001010100011101111001101010000100001111111110100001000100101110010100111110000100001100100110000100111000001101100110010110010101101101100101111011001000110101001101001111011011110110011000111100000100011101010001101010111000010100110111000011011111011010100100101011111110010000100111110101100110110000010100111110011001000110100101100011101000111011100010101110100101101100111",
	"1001000000001010101001001001011001000011001010010101100100010100000101111001010111000110000101011100101110101110101010011000000000000010010001000000101000001101010001000111111011111001100100000100001101011110010001010010110011000110100100000010000000111011110111101011110010111010001111101110111111000111101001111100111001110001111010110101010010110001011100101000101011101010100111101101111001110000101001111110011010100001101010001010111010000110000101101000011100001001101010001001100101110011100011001100101111000101101101111010000010010100101011101011111010101000111011001001010110100100000101001010100011011110010111010011110110111110011001110100010111001011000011010011001100001011011110000100001101011010110000101011101101100110011001101011101100101101010000111010000110011110101011010011101100111101100101010011011011010000101110111001001011011011100101001001010101110000100110000001110000100010100000000101111001111101111010100100010100101111101001100100100111001000010011101101110001000011001001001010011111111011111001101010100111001010111101001110111001001000010000000000011100100000101110001111100001001100101011000011101001000010010010000011101101111110010101110001100001000110111000101010010111110111011110101001100000111110111000110001000100010111100111001110110000101101100110011000011110001111111101011010101000000110101011001010000011001011101110100110001110110011011010011000010111100000100101110000011101100001111001111111100000110111011001010000101111000100011011001001101000101110101100011010111011111010100101011010110001001101100010101010010111001001011100001011101101010101111111011111001101000000100000110101011011001001111010110010011010000011101101101111111011100101100100110111001101101011011001101011010010011100000001010101101111010110010100000011111011101111001111000111110010101101110100010101110010011011100001101101110010100110001001101110000110101011111101001011100101110001110100000100110000001010100110100101101011101111100000110000010111000011110100001110010011001100000000101100001100101111101010010001111011011000100101001001111011111000111111101010110111110111110110100011100111010011100101011011010100101101001001110111100110100000101100110000010111000100111111010001000011000011001110100100001101001000011110001001011001111101100100110010000110110100100000110101110000000011010111001010010110000000001011000011011111110110110111000001111000111001101011000011000000110011011100100101001100010001010000010111011010111011101100100110010101110110001100010111110001110010111010010101010010001111000101111001101001011010101000100000000011111100001101011011011010100000100100110100110101010111010101000011101001100000111101100001000101001011011110110000110101111000110110001101110110001001001100100101001110001110010101000101110110000000011010100001110110011110010001110011100100001111000010010010010100000001111101001010010001110000110011110111101100011111100100010100010011010000101010001111000110110000110000111101011000000111100100110000101001110101111001011010000101010000001000110011110111001110111011011011010011000001000010110010000101111100100011101011001110001101010011010010101000001110111100010010010101010111001100100001110101010000010011101100101001100111000010110100000111100100100101100100010000011111110111100011010000011111000000100011001000010000000111010100111000111111010000010101100011111111011011110100111010101110110011000000011100111010101010000001000111011101010001010000111101010010100010111100011000001001010110000110100010110111101111111001010100111001001001100000010101101011110101000000100111100101111111100011011010111000001010000011000110110001010100001011100000001010011100110110110101101100111101111011000101100110011000001010110111001101010111100001111101001101101110010110111000110110111000110011110111001100001011110001010100000110110001111011100010110000111100101010010011101100001101100010111110110000110011110111101110001011001110110000100011010110110011010001101011110111010001000000011100101001110101001100001111000000001001100010011110101101100001110011001110100000110010010100101100101110101110101111010100100110",
	"1111110110110100010001100011111001101111100011111011101011110101011001011011000111000011001100100000111101010111000001001010100001110011000010011110010100101001100001000010001101111000111011001011011100110011011110000100111100011100101111011000010111110100111110000111111110110000010100100101110001111100010011010011000001110000011000011111011101001101111000101111101100111011110111111011110001110111111000000100111010101011011101011010011001001111111111100101000100100000001110101011100100100101111010000000011100011101000100010000000110100001011010100010110001000001110110111101110010101001010011000001001010000101011000001011111011111101101001001110110010100110111100100010101101000100110001101110010100001000010110100010001111111000010000010000011011100100111111011000011100001111101010100111100010011110000000111111110000110111000010000110111001100111101101101001111111001000111010110110010000100001101010100101011111111011101000100111100001100110110111111111011100010010110101011111111011011010001000011111110001010001011101101110111000111100101100101100010010101000011000101001110000100000111111000110010001101010011110101101111100101010010010111110011100111101110011101111010100111111110010010010011000000110011111101011100110010110010010011001011010111100111011100100000000111100010101100100001011001101001011111000000010000100111000001100000101001101001101100010011111111010110110011111000000011000000011011010110111110000011100110011000100100100011011000000000001111111001110101111100101011100110010011011010001010001110011000011011000111000100010000111111010110100100100111111010111101110001100110110000111110000011111100000000011110001000101011011110000000100101011110100000001001011111001101011101000110100011001110011001000101011001101111010100011100110101010111111010001110111000100001101010101101100001110111100011101010001100010010010110011111101000100101111001010011100110001000011000110011101000001010110001000000000010101010110001011010000010100100110000111010011100111111101111101010010100010100001000111100110010110111011111010100000101111110000011111000101001011101001101010011110110101111010110000111111000011111011100100011001011010100100010100001110000101100010000000001001010100001001111100100000101111101110011101001111110011000110001100010110101111000100100000100100110110010011110010111010110000100101111001000111000010100111010001101000101001100010100111101011010100100000111010011000000011011110001100011111100011001000100001110011111101001110110100100001101101010111101010101110101111110100001110100101011101010100001101011001110011010000100010011010101111100101010010001001011101010110011110001100001000010010001100100010001111001111001111110011010001011010111000001100111011001111000010100011011100100110101111111011101100010011000011100011010000010110100110101000011101001011011011000100110011011110111111000000101000000101110101111101101000011110111001000111010111100101010000000111111100010101001101010011100110010000100001100111000000001000011101001100000100110000000000001110001011101110001000011101111100111110111011111011011001010100101111101111011011110010101101000001001101111101110001101110111100011001011111010101000101001110100100000100101110001111001100011011101011010110110010000100011011010110101111010111110101110100100000001111010010000001100011000011110001010111101101001100011111110101001111110001011010001110010010000000001000000010011100110111000000100000011100011110111001001000111011000101001101000010001011000111000111001001000010101010000000100110001010011000001010111000001010111011011011111111001100010000000011011000101011101011001111101000111100000011001111011010011100111111101010000010101100111011100100111110010100001100011000001110010110010011011010100000011111010011001000011000100101000110010110001000110100001110111110110011100111100001101001010101110000001111101110011101101110101000011111011010010100001100010001101001011111101110001011101101011100101011000000000100001100000001000000011001111001011001010110111001001010100010111101010101111101111111000110110011011111000010000000110000101101111001000001010111111101010010",		
	"0101100111001010000100110011010110011110000101101011000100001010011111111000011101111000101110111010111101011101010001011110001100101100011001000011101101010010010000000010001011111110011101110111101010001111010101010111110000010100000101000001110101100011100011101000010010111100010011011011101100011100111001011000011001101100110100001011100010011100000111001100010111000110111101111011111101111110001001011101001010110100111111000010100010100001011011100110011111001111100010111111101011000100111101001011110110100110000100101111001100000000011001110111000000000100100001111011011001011000010010110001101011010101011110000110010110011111110000101011011101000100001100100010100010110010101101111011010001000011100010000010110110101011101111110101010101110011100111001011100101100110000011110101001100000110001100011010001011001111110111001011111010010100110100100001011010010010110010101100000000011101101010011110101101010000010010001111111111110001011110111100010011111011010110010101011111101000110010011101111100011111001010011110000001010111001111011000010100110101100111111011011110010010010010101010101110111101110111011100110100100110111101010111010000001111111110100110100000100100111111001111110010111101010100111011111100011101111110110101100001111110000001100110011101100100000111011101001111111000001010010110001011110101111001101110101000100110010001100001001001111001101100001111011010010100011110010110010001010100011000101001100000111101101110111011110011000101010001001101101010010000001001010101000100100001111010101010100101111100011110110111000110010010001111110000001110000010110111110110000011001001111000110100110110000100110010101100001010001001101101010111100010001001100111101011110011111001001001001111010000110000010010111000000001011000000111001001100010000111101100010001100110001111000001110100000101000011110111001100010000110010010011010111110111110011000000010100011001101010110010010111100100000011111001101000100011011101001011101001000110000110111011011101001011011001000011000011010000100000001010101010001110010000100000010101110101001000100110110111000101011111111101100000010001111000100011110011001101010011001000101101111101011100100010000101011011111101100001011111011101010011011110000101101010010110111101001011001001010110000110011001000011110100010110001100011010011101001111111001100110101000111011010001101111101001100111000011111101011010000101001011000110011011001101111010110001110010100110110011111100110101101010111111010100100000000001101110100000010100101101011001011100010100010111111010001111111101100001101010010110100010000000111000101110110110011111001111100000100010010110111100110011110111101001011000011111100000110100001001101101000111110100100110101111000100110110110000000101111111011010100111011110110110110111101100010110101111010110110001000101111110001110011001110110001010001100110110001101011000110101001010101010111110100111001000111001111110101010101111011001000100011101100011100011110010110111000110011011101111011001011100000100000000110100000110111011100010000000100000000100110000010000101010110110000100010110100100001111010010001111100110011011111011101001110010110110011101010101100100010101111101011001101100011111100100010011011001100011101101000111100101111100011101000001100011101001011101000000010000010000111001001100001110100111000010111011011110110110001011101010011101111011100101111110011101111111111001000111001101100010000111111100001001011110111001101000101101111100000000100110011110001001111000110000100101001111100000101001010100100111000111101000101101100000010000011110001100011001101000000001010110011011101010011110100001111001110010010010101001100110110101110101110000100110011010111011010010011110001010001100000110010110111011110001100100101111101101010001000001000101010100110111001101001101000110110100111000110010010111011100010110010010001101010101010110010101101011000101101100111100000001001011010000110001101110110010001111011000010110110100111011011101011000000010001001101010000001010001111101011100110001101011100000011101111101010101010111001000000100001001010110111110010011"
  );
  
  -- functions


end ldpc_encoder_pkg_4k_12;
