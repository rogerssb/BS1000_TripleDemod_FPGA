`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
rA5X0qXbvnchdGvwkC7BLwL0xgsutDscHGewYRLrE0wPUav5YNWyeLFp7cG89dWIvhTxLRuqVINg
qgbMFWowoA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q/XfOsgfrfXHqICez3cQRnLbb7fFt9pwvWssHAdAJRCU0pDVbiiNciCUcSB4MjBPH7zFjJNvMljJ
FRug1GHh+3Oqtk7b9/imIg0NUHDuzpqXAt/vNeewoG6f/f8LdzHYFn9VI99ouK+tZAY69GUxm8/x
hM0A6LIVgAbehMz2FHo=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wDn0LliG/9RUsRYVHZ+BhgTKKNYUa1z/Wdg5isyTtebv+qekFNF4qr8zcP82znisQ8wk72OKuOxi
4jpqxgS69ekyBqbL80q4THc0sMGbWHFMJw/3gGWhE/m2vrdmiUJW07woqko8UqYBBrM4m+MpTRKa
WFAk01Z1Ppy8SR/BymY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rCjM0DrXgYJvcXbZP3O6VXbKJg81UldnK7jNokL2Z5f7fP+aOkInB/rcyQufxHALCZMFyH6eofqo
X0nGeYM6AZpljtXco98yrLoXQgnZUeFDraqqHOKP4Pv2SXgRcRQqfolVnvxm4bNupqHzK8oo11+L
+rJOSmEbl8UAQvzqGYYThU/E+4Bf3qdGaataIgaVDWn6HNwcyorqxF8rEgOh34E+kdZc4+L+oumN
6DPFerPqTPChSosFwyUQnHKsMHL1jQe7Ms0GnSS1vp/qXbCuz1LN2ntxCDUTEOgWkpfi+e12+bo+
8BMAhg3wryWVRKH8VN5N8zINuxLnOeS3aSNRgg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vJ04Z2uqYe5dsOdfBl1B1ZpOu1u2Rdhugg1O7xJzUTVVUlh6RUo3pyvpZp5eBr6KNzsrsfp3NtXf
lghOIhxTkpb9+sXm+SYfpQVBqCG+1LANsZbDDlNdBmo3+Z5iqTHT6WmukttD4m1V9sh7tpAxNPmN
LToWpTLgTeSaU3U9guGjCHAdG/9eUoqQwwhpiD1HvfLoHZgRBfleigGtrAQhSxCT9kG/Z+VZUp68
52m4abNwjH3CR8PSQS95RzqZVCb+gGm+g6KuirFiyzGiqMOy18gbmaOUnMmdJsimzyfx6fPQ6ffW
peUBcfD7OhQwy4TSP8HJT+FOHY+lG7f6icenkQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TeOUCy4oivxfpE9i+LrnEp3zTm7pKagAVD8jNi+kzqrWSrIruutUYzPLzUZsDyqIXF1QuGJNJerr
8QQnVUKALiqEUFkMwJD4M8WSmnPjrPLZVlzhAa6s6gIQk8n108y7YILuOjiMcJ0YWpj/epJl73Uz
VsRSPwnVVFsJZ1jR6gy5JoG/VVx02JtGloBh4AspKkR7g1RUKQ/g8zwkNkrBBPvhX/IKsZfIJMuy
35gDTNKwZdy3LjajQvfrhHBg6pRl+c102EGVfOnbkKZARKtX/kHa73bNtpYCvmdKt/a9sby2gHqg
2NXnGAKCt99ahn3MByK1yu/wZqtYbFM/SOOLUA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 57632)
`protect data_block
5afvtweQGx6Tb2DD4FgYra0mRBBREbtb7SB5CmnFXHHJJObLhEtyzmeq2JoJdtor/5zvKggIdSg2
O1pzfVDrRQUjiIOrIGuv4N3XgEGry2yu+fbkDODFm6CrSG8SJpk/CZFY/w5qrWXLICjj7ROy4gFw
2Vuz9ajEkU6f1E1vpa4FWOV0HYPDZ4HVdQ2+dKaPUyT/uLT/WbTSym8vPBGLWHL93SkwcYYOlH8e
4FOkNmUqqBeqPdRiahAXvSGoGNRNve1IInQub2EJutrlDSpwuhyAVcnnfjRC+Cfbp7GBeEyToRaw
FlKn7+Xu+p7U+EQSS7599h6eRGGR++S8SJiscgeqwiYG333ErTuglNXOcbqH72Yd4H+pDBvzXRQF
+YQNrMgAqP1LU4rjFWzWVRFdU9BTT5w1kBYGIWW760idbANxv909M5PpcdApNrAGZGT+mBLljiKU
quxEZ1oEHtr29g/6vlXvEcVSm0xG0cPSBKR1HSEM0ziWw0kuNEEKei5DmZ5RWukkWkZlk9zwGNwn
obpG3PHyYZOwkrrnmhxlrwwj/d1fkmhkL+p/lhUNl7dpS7gDM+5p+6nbUVE38rN8qZC/8z9Lrbkr
91/FQ5crEO0uK/z7mkqFY0Q1rzW/97TV6gmVhoJ1LQdQQ+1RUIq1GIvq+V/3LIumNQnV0WNN5L62
y5ujQuWFMw+cDG6v+xkZXODbogAQrZVTz+ogOH122QZtk2PSqjg5XT0X5bDdZ5faNT6/LaqvXoci
/xzCHY7Mr43CmF7XRrhKo91HUI7z1AoT43Rzwb09qtS7grfjJjv2++7XpGP/5p9AQWa9VidMs27j
OEZFn1wOoCeOmLnrlcCcT1htjFvSS0cV4pxJSGrsABaYDsmIEyFvuUiko+yeNF15xRWH3/NjKRnO
0GHFfJ7tTDQD+iw1r8wVE/xbhFtVoaeW77J7RcEKGoTz+q61Uls2CFLlbirQitJWm/4DcW9S4soV
DU22lwXrFk3//e+15fvCf+p+Vy2Xx3oUP57oTdLHWE/fMF2/V2CTM9TV8v8fQFfFEKfCQxXv+jBD
Ynlu/afdNQ4LtimWtPw0U+nlKGMhP0rBSM/LnQq1qgkWCsar+Qyux64sL1IARFsKbuvd3kOy3QA/
xXFhzDhD5BioDqcNzxLejOVmFCXNKKbemeRM1oEVcufYaSuBC2pXaC9XSwZTjkWFE0tJ/w2pkCaa
6pSbdVW3JIhf0PHdIDe274uoaJTGDlSljhKAjQGr8yjTIM0CNSrA7SDlGyoptPvy+ldb2HZRl0TC
KinKCbnWvFXema7UHmiOGVdhU97BjKTtDxjE349pBXuTt5ZGKEQgjqY2Q8V6F5hCy5SXq08fe7zV
AnzBMJwH6ZtJeX8GF2V0UiFhgDMLQBWfKKWQEEcf8+IgV0J3oNTOtgmZzZnpwWqfRnVW/Zu1Tia/
XeHilZkoQ2QXW5xmUUoUWYl10PV75K2VdL2OWm1/MuxVBpyl2SJvTHtU1LVRjZ2YLid69Id0HgbH
h1QdfeMOpGVwf/gJ5cPaGGsp0jj7YP4NxSMRXsb3U6XHKw2zsjtdEhoOd42TYvew+WbpQHntijIk
QhpLeBQpdWMwnT4BBbsD71PvEI3hjHRPYTE6bAmaRnc8YR8A3yjdsCi5lsRQ/XmKfA2v8zL+8VGP
jGuzpNBDEzYVjMqUE+6+5E7vX59FiyVOlQYR9Or/0mjxhUe/AW8Msz2BEV/+V4CWlauFZ/htwZ5d
cm1b3THDvu3k8K9pyd8AFOUhEcBKn4928ml7Ka1bBVfytMiU8pvO/5bCwVnfxb6Eb8GCm351+5SR
9Z56UYJV5nrG5LZWaYy07MaDRM4wY+ErANjL8/G8jZTZ4NeakLrP+gGFL/zVVTOacvMbiVljrIJx
hpY+olShf9TA26aYRxQ0bVLLCODffT5N9WXadvkVNwIH0lhhV+z8H4Gdm6JEmp/OsoUTVJ6e8b4Z
rI35LvotgASPHgGRehK9vy/180VoegytXVu5haI9C8K5mOw8sn9iW/0DsHC5haqMhK2Qs49NUpSh
uTy37M+Ez2DaKKELebaW8iRaVEDnaDxTN+/FVski0YNi0NEWLB8/3UF0DUO8fx09PRfRi0ZZzQ+8
sdoWzM2Y+bAg44mWHlnkq0kzkeRDQvd36OSuIurJvMsyZqwaW5FEF2aMuY8ZTyeE45Rn6ZPVNltQ
0GVU6H0FA+mh1Y5vjtANOLjEvYWYo/m/C77Dk6KMD8ru2Q0UMvIpGEwgKk3BlT5MJlYmF8Znbdk4
fuDrxnOgRMWr7etoyiK0DR87QCT3CHak0wTpwvQYrXBaaYYOwJCx1atVBRw41HraFwI6uCM2wYCz
P11WONVHBnqtBxoEAuKDxBSF9Ac4SryFkdD6Z1dTVG0+TcdTeyAN/HtbXsj1a8RIFW7N3tf5M2wu
82czq2qSuYvL5dzx0y36R2Nv04JExMs8Vm+WQq8Zs8kBpyW7J+wqMLzQTo1Ml5ijbTbGWuOCmDdR
tpWqP8eeeXJ47Db2LwCU8uvhAKNdpzF5iR64KTUUfPeoBLI2g35sztUgKBLli8OEkshq5QR4gRb1
WDU6Sw5OauHfA7pIf8+eQCJquxIwpKoRbp714eLb0kVTBoJuyhmS2MzBsjZjJTOT+1EKuAnNoG8Y
x/rF315UfoCwmGQpKsdVfSqMoyPlSekzsi5eHR6M/aG4m1P97XLfMpcuBT4JlV8XZ93vZt8kcHdW
Ycfh6Sroz1DK5IkG01PN/Ypv1r6iVJDLQQ7/7nmq8JdDzsm5OICPqkZSUq8/bB3oc0kvD4+g3ip4
34FW13t5WJRl1HSAEZoa+4Dzs00OF9zhBik2jvn/A9vwQqL1G4n3ranPHmbokPGaHVwauWV0Tqu8
GNBqbwC8e23t3RsJacLKs+yXD8yp3kaeqjFFSBzPGBIFw7lrAKXHnkmzla47OneCEAj9hbOT2Ph0
ydvCNHFdEzyd45S4mr7Y3e8IePOtzQQq+62B46CLLGDsxUtW2nhC0GLIxiZ8VewO2ZMoMPdaiC/g
yKFv/dwXpM/Jbxphits9Y53iCT6UPCHgazk78njJrX0GXvWOL82AahsWdpLkG9VOAB7Cxj2CF+l7
Y2hgyW55KZuem5moRUZeHLsPxGa6KxeL2OsQJBoGJZiI8955Y8bbDPAHhNT+ztPjcEEONCskc0np
M4BX9mvC34FPuewCcHe8G+PaiY95E2i2LsTdeRSvjXJY/YVoDitkPJMe7OBR7cO4zufnQbIkwFDU
JU8WLSrt6m8Z+TpiXY59CAY/4CrirasJYd/CQchteCbnqqTC9/xchYjPEMFhi3IpaBonISEySDiG
/2bwTK0cEGoLuP7J5pj7ro0eeS5qCHPiUXghNn77tZn4wqtydvSmJADyA3uqZUJFJajqjwNTggXo
4eS+UbNdOP8YhIyROzZJMgl3sLtL3p3A01/SWVB3da7pGKRsURipgK3FECNfpcL59Ghjim7ke0B+
/D6P+ivdWavfDf58XaEsN5cVFfa/GXLW3Y23dLX8lR6aozlUlmsdpeudmWTdjEUP9Uef4/526Id/
ASDtv7OlXWiAq/qSaodwNPfxjTYobA4kAL7cqaxWO1fQHWjr/9KXvpsANd0bp3G96Mu+XyVII6gk
4jETA/ok8S9l/KH/Tthdc90v8gKpXBG6AxmsLudGXqbTYE1DTZwrXJI/IqK3a4AYYnTe329WC2BE
ooU2emt2UF0h9pAAYYzBao9MESPJ7KrIii7kwLcCn68MuhaOLewbMVhosyNorA8s8kfQY3z9TtYI
eervKtaYba48RepnYyhJct/t8ScrYxNrKubY5GZTWNqNADkAU0r8MCajuJIDGvtnA1OFnR1rgepP
w4e8Ldtk/mJglSCJLjQETzBEY/jSMWtsvdwfrsjnCGOwCUom8BHd/EsetUPx1AU4vVeTxVeYGS0C
36ii/0yt6SuTDocy76e2q9tOMH9kOsvRQUAELUWiSyZIdMZezusrppb3Zf4rds5SI3roNIcRHjU4
juVyD7FFDk38yJHyZI5WO+576BH+2Krm3ZwImGtXpDMouXvdR8yHzdn8hASNkiPR7wVktquTXjG7
9kzdOTywUTB1KeJG4bh1HBaEwE9irjQHnChR0p4IriR14Sp6Dcx2U2lnZfaKeTp+jMv0rAFsQNM2
6ydE0h+gr0Pje5ECxl8uJyg2DnY5TZu3q2ccHKnZaC0FJ9pxlK5SmJqZBUVCcLtNHE/EDgDzN6sX
D2wItzqPlDuOm+BJNkvXQsR+lAgJd82HdIeBF9hYvmcDbvZA81ueS1G0xdaK753t3E3fCmJyp25H
vGJ+aOzTewm4XAqMOCKLaDNkE0uqm7yUmFZYxgN/Fqv613hu3V4QRuD50wdLXK38LKCRCnWCQ3kC
85y6IirnKkqqFxM5R06K1VHSQPBNFMFmBnjQR7g/J/NXv89WI9zde8MRpv+f2c/iIFZ9AON5mOA4
56NKIvQmPx5I2YtSP/4qmvN3ijYdvjby/ZDh0xlJdSkbUYi9rwVOUXzCd2XL0Gv+TY/lUNxlHzfB
ZWWPbj1r3J50e4/HasXUHs04BDDFK36+22zd09HNKNgivv2jFYfE4cyXiut9WrtifS3zg9JUsEIp
7SqZlVcQdUrJqxI6khbsFDtdUYVu7xdJIaWW2eOXJlUYZsmP+YHytZy2MD2eYP4Xm4uNEt+w8qCK
Ah0C1UgBZdgGi2HRuUzVDVKHH3MBlRFKbTPZZ47C914JcW8yNXNBewrjRFrZ5T4l5oBtAnrjAdgf
QoU+0KASei77paOuUGvUcxPn4Xb6BuBrimq64LU0RHmycBOHI40VpwmxgEbAfkwVNw0Y4Y9iplNH
60yQ9t5OeAQ8RJzxO9MY+BxfSnPEC/rGmKhbNvEG4UY8sFci3XlF/aBaC9+lk5OIINZ5kFU7Zl6P
mOYzDPo7IZaqmWN342HtlY+MoRyHf06khFM5RaBDFNohbjkyC/hMs2D4NRF3cG/Y3jPNF2qeJFDR
WqJUdzG+VGpCmjQWoAjzATOeZtZot+oXYRhoOwDR6FSI7zi5+i0ZWW3+YwVkYHwGjhOnThB1VUp1
AJ8+A5kuObdjlJ05u0WedfxDuDmEgWC4ylWPmXVc1/7pMO9ztcOIumz2UuCCBb82/SWGiHABD0SI
lufkS4uvdtQZDFYpDoNGJ4E0uaq7VYqmOMvAW05A/kzoXtrS7McESK0AVkB1N9qf1XxQrXf4s5s/
hrDNWNNlajHiL+9jfQkWv3HzrojUOa61uAXxWzOBONTyI36HqPn0brCl5sVWxoCGmRfYWmFvJIpI
adRDA8zAljBWDpsgiKsYCMh6n0jvy25TOlLoZeEebJJ4N2/9azfSKnam0hsRNw+onusbW/8Q9PB1
pUfzEHc0XRQCPjyoDnL2J8BxUcDDt+eqP/7LhVGi3Yj/sm08wVolIXxuMLwIRM1tpzzXyGJkSLuQ
Ls7GuOGvQ67GLgeQUoPjEkQPxnUFX7mzBxeE6JsTkbw0xpGJogMRRX2Rf3gUwrXm804LmWm5jQTw
c1YGlJvSBWrrElwD3ODrvpvcB6gVygXMDp2SEuVDPrZC6pC1Ke1FuEn2NohazyU8ZO2zaELrp+Km
d0O4MsBlELHsPE5cO/66ipIjbKcOTUWgjr1BErBetOimd/i6zJE323jNl4B5qK3vLw6W+Rku3MUl
YKvbERUivWk7HTpTmzWwsB+0JkEuP08vW/8PHtIZrBCfX7jYeudcVJp3BadQZ9G085mZWCYwnlyw
p5Sgwzw39HCp+F9GmIbymI0kTiYYeQg0TAzR4zbHosToXi54t2zLRJwCWBFzUfUpprVqpzvsgT5m
2GomrYNR7A3R3E9aWOgA21lriEr7F1vuun1IvRnxjsJ3dJhX9jC3rkUZIQozGTzw6c+q1QWESW7v
JETKCCTYHIHb7JYuVjcxvFFdwBDJ/IxkNy8h9hJMvuuv05LN9Bz47MLq39HqSkRwoStVvTKfmpnJ
QlrmEHHapj9KgekX1FnM/+DAVzzQsoH4Ej/MwN+0+ZYeSK8e1DzrkBCof5p9a2pYXhfmxR5XHb/v
1V37Kc4CxZFFmmafm467A/zq2uKOSpFMpFCEsFF42IYysCPKm0fYBRU9TMZXdvD6oVhR3n1cm/vG
NAtPlxNZsNywLveAegVG1P7UbASulNuAiPfkkuN2aca2oxRz9PI8X6Jk6j1EWiS0/somjBW6gt4i
lzY8dV3zp7zMaCpIQbsZp7knEhvYq9f6bHl5qFCsF2HSsPc3hQ4itMzOPsUhNzAozCuwOqaQKCCp
VviWctTfAKGYqhHJNO093JOleIhVU1SKDE4+89uNvlHwtzomNTzPzkv4KUvnvV65Cwce7a5TfQDU
w4EiyVhAezDbGEJiW8jeHQMmHnm0fRbZh/B6L2AJUp6tFGqKcufq+xXKe7QKC21cPzu/c9ibEjQW
AJ2CpUARlGCpysXUqEUMW2M9mXHoYGPYU79wQrhvMBdwpjdrcLX6TzBrWWGSX1HU92mwK9L30X/9
L2hxezfNNPTFVExtlmwdO77+jSFObem8an4nZAaLIqHkFKhfsnSm50NAM8bmlu974AUWVktZsx1k
JN5pifpbSaW+WMTUrvvay6nn23We6CDV2iKR3jzn2QIbF/kYtN7kEcT3q7sKFkgYLlZK+pKFG6hB
BgqsqV8+D6hAkyR1IDDASuyZNeenpGvQ/PpiMmfPIPfWugaJ0+Zw1aIDIOdE2FJ9sPJ/iVQJwrz/
6C/JSkfhqAHj1DFwDFZaYVg2kdGrLqhxRV/8Cl3GoJqC+K0EyAhplLpvyHqHD3yWsShOh3NKMZK5
31ictioDVEhD4dbut9AoNhBCAHRFfQp5oBfAiD4AP5+iHBuFDCGOrQYLdU/CyBXHtKp38TXk6xMT
qh9Iug2glfVMWUIGsqlVBhjfBpWY7rfKEKUiHQZgNx8DVo1oLThKluXHoY1ELZMSCx3b38eKlNrw
s1nhi8B1/4B2qhgntw+jFlVh46a7hk1jHtNZnQdEIIm7jLADuqllpDB4woPoFUfxFd5LGZKdc+Ex
YIMkrYuBjNfBXypZLV0plQOdSlosAC/Xf975dC+AwPXGFzAnnO5q1DM6jkFNSoLm+e2wU0URh6pf
sY0GcfHmmf+DdFORqUM/VkKKlu4g35NbZ3wjdiYao86ccZSBVMFxCA84I3ycTHtTE8ItwLDPmOZE
DzR8yCVbItcHiVI3sHXlGhtvqXWd72/JrcZkrHR7NH6+D2WiGdkdTvGQRXAEoOskYsJu+gOD1j1t
8mRLA467DX1dWlhW2bjQ0zip0TFiyaayVXu7HazEG4Lt7u9i1oHlXr/KWdC87QWV8yXLzujnKjnr
rR7gRadbNhH3HlNGVzitKb9hrvKgtPQrH4h02gRgl/p+t7qvdYewUUiiJ4UB8AHGyxjTkctkkHes
A0CiwC78jdtrQVfMDQcsNWjOqRz71QiGJcHVlLI0l9VmFlxFdg2ESxdj0vPG2ttr3kOjQGdTMrIJ
8megGsfXXUZWtkzV2AO2TaH2yEcg7aItMdJjREa/P6jksQPSbVX5douavLzBORbTJtIGJu/bTrKO
nMO3gYiaERGT5wBUse9CuAX4vaJXfvCIwpxjJT56PmIfoIWSv6xCTmxyxiXHEL2QVAUjmCzQM1x/
qaZzMJYTFExEhCndl8dbn4vZiujwRoYe1uhwszQLaFZKOTLeyPh33Fw1RyMDQpWVTpNBJDREp2sc
UpDVo1zU1w2GM2UMWE7tP1Rm3ePLVIio/k0udUv2+/ez36qma4jqz+5l4jOjPBlwoEHPG4X507pJ
LNMx/C38OMZeII53WCzBebiZRuc0nw/aguVM8uwUBReDLIGUKRb9IRM/Z4kpI7RSgz7w8LJYbttM
j0ufLaa152SFGuL7Tnu4EtCa1IKSGpLU2kAbW6fzH7oBWnwQiGfrQwHSsASOXV8i0yoT+sqs57hg
cM+opR57PbmdhxpQBLYM2Di2sRrwmjPk0Zj97Qt1xCxHEmqeK7nHCEdyAccbp78ggzk1F9rxLRNC
oZIuCCWIMMwddch76AkueCAfLv+VkwTmxgzv1uTZanipwE58PfRb+bXuWjLrPIonce6mCkCy1nQ4
HZPKyUAgwcbA8euK3eX/ISIf/G/NXsKjrGJgnfIwCBg/Wr/il4o5XVmYDds+1yOiw7LTp1Iggc61
YDf3YOuUOS4HmhBzUtQnvYzz+IrTQKgYLpJKncNpCtxgDmRrffvtcmlkxUzcIZuR41UwZE27rCkb
UvwxRiLqS/XeYtTslNcbxh6gf7zXvDCk3GC1YWko14ZuDPZU5hsNI5JzqbAOgxddYOKiUuczaLCq
zQLEVMS0g10+QVYbRw2c3mGC74+bpoZdtMuPt/xUjzv06p/tKdc3z2eOezrnZZPIPL4bIYYQ8ghw
p84DBRNvm2nLc02rOURKX/NGNeQxJOKK1ryq9iuzCP4hKOZmBJKus+XBOwkH6ie6HLrNVhMaE2Uo
Ya8PCSefdQoTKZ0JaW/Rari1QfVbPhOEWyKQbzG4OJsjTjlP1/a5AHYDzSo94ygXsMdEH6VbDrLQ
MTSkpgtB0wjEsgqh2R7LwIvdkX+iGnIAf3AAle7W8eztiBXXIGxDXCaFO9wmEEn7DixZT8sNySPt
AkOpt0K/biEFaplg+FU7zr1rb1aZ73UjBPRwoqmVF/EQ1sVpkj6+shkfVgLEyFcGbqJXvLDGTfYI
iWLCxeG+8326SLlzw3hMaZdeMjIGc5+4XZ1+/jvYzzA5NPZeZgO3pSUWOk62h7GljhUYpx4RaAUm
3JqKImqpPoatDFJQDDOSH3prqIn8/bxhpoTcWQsoOpT/ChSwAw+3a7LV8gC3xjkujgKj/uvKaGau
rQF6VtVCQJV9mOpSFJfJKh3eka703fETXdq3O+KDYNwux7z8q63K0guTvRqkWZnIByyf6voveF+h
eo5MBo2HrRfPMVL6R2pjaxMj/UAAo6UbZF3Lt1HevX2Igtu/ZqqPkzXvAODUIi5VADFdixjrkHlI
PdopcljON4/9xnhaeMo2ILDAvi02NGXAeYI9wXQucniHy+d2l0LAWcXW/wgYCAOKH5pSomzg/g2h
49wnCykN/xrusapiGVCX+9Dr8Hbdkpbb8Ml6NVQX38RK/q71j/dKqvbGvpOFffZdXr6av+tSzUyw
RPmMa+xHGqz6RMHP4AjWzC2G/KXrFxQXzQa2V7dA6U/JC53finvuzCDQeze1uelofw/glB11Bofx
EJ2fInf/FytmMUTri5mpU5eqBL7/SboGtD7mRSh7sYuAt9jsGdxNWDTAjFzLgHEkBAEEHplHuT+b
dDkscZTASajhIQfadalCrXkmdFEOqLNeFY61AHWPP5+1aMMod/WqEWDnu/LlQi2r/Q5MKhXYLaem
SOrT+95kLwWgkcRi3rG6b6Zab2POxGozu/Z1bXi5/Gq33MLnltM54yk7kgY6qBxTnLP8Ii9lS82S
yKXQotAlryE259lpZSnjoZ+b6U4xQyd+GRFFv74aPBplJOAiCDyH1tyEJj7keZuaAMTrwqPzLtBO
B8+dQTmMj9GeZtVqGkLVWI+A07SailnqBUPbhm4/NwDYsC2cB3+KKAGOtm8oPirmcEZLH/5WGyaF
6IGA1Jf4d52WRjWE+s0OFvoEZIDUi0tY81R9zURYY3lEKlIW9yhaHl0RiLSo3QKI27kvf3+3hpTc
C3/a4vL4ve4L7xa7anFHgXo3un0vFto+I4EEc1j4ZsJTIVbCyTUJImbb7CJHynDx/utYAghxmnYR
yySOIeOnhMmjLiUDfU695D8cNTGFV/YDY8nnjWHVHPLq3yipEMVY6OLDDVdvzeS+aIDTx/jFjB4O
pLpqoMn3MGMn1JmatFYZ8ZilbtVWV7jLZu9MdwCwDCWLiT+n9SD6/77yf8c939oAulTxMXKyxB6U
4ZOJfUqEC0Dt0wP9QY5gnqrDG3Qpmof3rkSSnatLFK4Zb8uxnYUC/B/OZA9LGbaZkY6vcnGNWfB4
2oTm86/yCb4FZa+P/8ybRVKjuT25DgYKH/L5iWKU7eddAUN35rf43kMYY3RA+OH8KvKtok/TCYcM
+gNDzqqWNHHhswYOURyt+DBeqIQPOoF9b+7CeR0aam8yDChWNcQ5WKkBdGwvv1FbBfm6CM13wa/b
ivwc9fnfWI2ZqNi2/i5ZeATpJzegN7w3gakism7QQtXw8gDw2Y9VMILKvPkln7iwDk2auG7p/Dfs
xbAuRr83C446X7w6jzfWDr9IDfG9gZazWj/gdhJX0eGEyxV5QTPUbq2UwcBjToh11+RDjDc/QbUS
Vk6q76qPhYMLtaSA8Zxjd0CUWKy70aI1T/DtHkHh4cvbalM3LY+OJlmaLrZQjVK3Vk5/G6tYgPOx
QEiQrfnqMk3qb8e8B4mXNFvG/pzEVlPHIKiu9pFBAD5Xe0yQiVksnlcaQgtx78BK2Hf9aP6RC+kb
OYKNdMWHQUgUQ4w+KYG1MXUUrCHNCKDollQ6UGCLtdki9gDprCy71aX2BUm5clM/i3VInAGfdHke
RR7VgReGWJ0kiOvf7icgCrAwyLiSquEIRx613bdOxAhtxNICLmFriQ2pzpJSxGg7d+oK8zDE/rpK
UPOGH3X1ITRxyOPj99w9vAsFkN5O3LST/+mQAJ0lW5Vb5dI81XQbvUO1y5otrus++mvRLgwi5gnp
WID6kuYGl1AcPlDYBSQxDwcIltw9W8UJ75K6ULJdX731y6QNozXFIdXViSSBYsxou/S3K4J8J0Ig
4M6USj/rJtvgZ3FbJC+B2rYaqeRacOhugI/lwvQr4Fkqq0UBSC0gqdL8aB0IIBT5nwhMQrKn2ENZ
3a4lZJguM0LRWd7ai7OX9+Wtzodf2g1whaYEPgBSxYtNvIoeHtc5R9l+elZlFvyurOh5QhH0SJ8Z
lsuNnPyRLIRev9L0mH4vAMXNQy7q6Oy6FuVoyietXNXRwyHWXt1ALmoryDfTYfrUBqvCwFly68Gn
3jO/ymrBL2pRY29MgfTYMvPwdun0Ox/qSej+BkBQbZBcn4pqX0mptBqX8q4BSPiedE6f4+OZB58w
8WbNp2rqbj/Mi4j3yMrEF4vsQyyNukaRrVDCEyrOsgF1CsFJiMR7BxQ3jRCekaEhHbZSiqDfSVkj
bBgekjfqH+Wl/hzecz5mAuYJ4TkZ1NP1dFtTM1QOxiTvwe86aR23ByGSzguaw4bPxbvan8GdM9GH
xMGLwleZVFcnXjoU58IPfhEOVqdG/Wil29a9Jwp0C2Tf1K0uP7op+HaePInzSis6uLjPf8QU0dnK
NpWN8KO3wBWqVZ7CazEtPgdkRYQvZp9LOHwCedYQx6bNKUnU8cxm/1OSKNFXKyp/ixEPwa+gZAdU
zUz+gXIG8jwPdeemt/2QJfH0SBy4pLR0fL6PXJETV/+tovVEICnw/mU8gs49ubMRRJvJW5cez0CB
C3+1mW76voU0pcIBGdRCXnrWOlGh9FOzpSjdt/4/gvVqcPdLNOR3Eye0V/zlDvx/8/kwRt9IrXPU
8EhQmmreXNCgvYxsuxqg5oE0E11pc6GhoRuIHP5k6WomATGLckKE146ON82BOgPM2yioCvfpN5MX
O/5SS50lVHfmHmDw1qA3dxG5FPRO79WO686onOh2khY1uDfS3c6gZ/xGGabPizQGsfAbyyHJF+4Z
BlpseqB/TFBHb/+y7rtdztMWfPgz1JKAc73mg6XFqpU/kO/g7OzZ0lTJ+pxpQcOXScyvv2faxy3H
ekM5ZDOFU88KfAV24TiB6uV1sSl+ua3XDdm/UOvM423xxpB0qnS2pPuWq89D6nImE1vSSkxmws+b
iW3+mpjJBbLSw9VJMKlucN5jOwcamz8iec/k4m2wb35Vdv5EGov5dFWYwgb0w3HS5MwlhTpPlnxC
jL5DYXnQOU380MkBa7AQTpSnDG837AlEr4u0oJDRoUsoxjNuaKPKp0yg8Ob48r6auQ6smj9J3q8S
bw1L/XHQyULn2GExK8sQgTyb+bbHgwzQQDqejMLWCnB9kA/NAAyf6pzJ/kREpBBPFRuHccb+M1Dj
xSYvWNU+a66HqQlaal1c89DkcOnSS3k4uDpx6uDcEft9uJZUeumJGHO63vPZENRg7PZptFsG4sir
Sa+GX2bpYTqPc4ya68yj++kegPRG+r91UxxPCLmiu+vRvIshOGNC13eY/ix6fh2JomgmfHTi1Is9
TSfpUZnWKOZvV1tKQsxUeeOfqv7zjWZLCs3CwmeBe8b2m/uozHdcSvOXZzhTzPg4n4+OlGgBxUdV
1jEIlHBD3yYC26WHSIuLwty9gfUk7gogkEn61RFa78UiM6QMpyAsM4szF2TnPIsjViKWjBUqqC1l
AJbkIEQqOKdkEIwKU7QqL1LGwdgwFl9hs6O7Jzh1sXgEdMAEeYVe00ueDdxImKaDaG9pg98D6SB+
28NUhnBu1klv5Ut05GPMuOHNaRP5t+1WU+nreJVdU8No4qqkZ/FSg8kx7LHxtMghtii8M8PdRGAO
g6japx/xEfit1wAzXn4YbFd/QsdU3shhD6De/2xjVTHo1evscJngwwvgRi8j/fNsDIKwSR4OlpDJ
KS1V/r4SIIdTuyZijmnAnu3DPur42Z6TKvjzxDsSI0maIlOvP6MQQkj1avBe3I9pKfAewHNE24tl
42gLZfMD7npgvSjPd/yc+mci1g+kRzNCBrk0LhCW6oMIF+tZBj9XgKYRV/t4gvmNxp7hx08iz71w
A740Od5ZKukoKC+zySUjpqra2HV3c0pCoo50f7IKgyhGGhx+O8zsgVrrKyWT+Pzbq+kJl8RkPoIj
TTEysRc3vRYtX2RqUWPFSooXKsSCqEXX3irQw8JOWMR1a95u2sFl6tSW6iLVqSOziPjhbK0+xnHE
j9O1H9yo0UNmgb+q15op0pvLjV7j1Fjjk2tYfdcFquKcZNYKkAyqHq9vRgHr+MWi9Ti//8Cq+Yev
fWXCFmTv1ePWBwk+kXV3I7fYQclshkqYDOnRvq6ffWIWfHTYOb9/sKb3g+DM/J5tOtdz/r9k9hTb
LktTfU6/TRBPziaCjZTX5GWTJUxVUU/GqeCiFkSTH+RGl2+82THu/Uob77MYBnU7yuQOetTsPCGu
FgEJUtF1b+rpKn0SrI+itvu8wvuWOcJfQOO6v7IxY/9LUhcuZaNO2uan1S7yaPRj9yCubA+wPDp5
yP6i85XxC70nkUVrdOh4D8PdN0UKRtT7IPwf+L1wlScw4StRuDHfNOcW6r6Z/Aha2wJlXX+B4qEK
ekQDqioHVFGiI/N0xTMBKOlkdidjJHbrnz9nKha2nava53JoWOYgI+uJ2En1fMpyqJ075TEzGx7a
PGn8+6yUpEcxvDz627R32kDuKc4AvwbIpYzOqyXcCJQVmf0ZXHWdba4NCWEXugCUtaITceRWgTm/
qz8UY6stMuECsIWwS7qBxcN4rKT4mPjYmXMt0T+vmnEonBLCgeWaP0aCFbFjHfVkrBfRm0RLnAw9
bqb1Xx27PTxVdyqFB4hXKjNRcJlWgEQ6SbrCVeY9d1LhwbhCnFv+Xf9cnJDZJr01UZTeZ/nwq/lp
ms4mOQUPBxb43cYiLarRCgKN3T/ZfLxqJ6yNegEDsoAKOIfvhtgQZJfZTk/wAB1tCZvFrD9BLnwk
stAL8KfMHLL97vG1tJbouB9CTbQWwsW28O8BRGOSZLOQa5ENA8ZVooJ736IzfKUM01ZYCudT95OW
5cPG7qhvtoB5lf1o7eR2/RFG6qXiBO656TcIwL9s50SW0G1fVRNIeKvsJwmUMPpCzujfHN4zlyvf
TbUWCvIwzJbvbh5oVQv31rhvGHEOFlQPUo3Jc+jQ5CJDegIaaJAOqJsOBZf/gtC8+Tr8o7TKm+hw
MH22XL/TFgIt1a+R5msu8BlsQCucHou4fIFj7LwWrVEoeN3+t0prK+jRIo6sz0dCeSGzrZKWjkKQ
Bb8IdEulwYouhSt4x1fX8y1+8dybfD2BbC9sT3/oxjfcIePFOJh2XkfznydGQajdhHBz06OcSjFm
yu5NvmKZ749qeU5vsFQEjulQMnBcR4v8a7Mj77XuG6pwADnOcmRThqQlP1u+3uVJbpuljaJydETK
YaBmIn12t5wnimDSgxnDInzQwysbN7R5X8W9agScyVFa2Nj9CtIIlnYZvT/kUXuqt8m7kfyZm3gD
Hv9fyhH3eoINSuGK3jHGm1r6j1wsDqfwZCtjKnyr/r+3KsQM/ABO2UTvSfe4UOXVmZRBl2byRZeo
n6/4R9YZi7JNgLDBM5h4iYRMon66W76/0805VaT+Ce70Wf7N4hA0bs46JtoGeK3rxnO5/x23iG3p
L9niD5IEjpTPcJSpl6FFmo1FuDHY84VLwErSLwDAzIPpW8yvTRPveMHXv/R6hjCpdwBckLYHlpbk
+njSoAeBPP6IBob6ejl8sGDwjyVW66InUD7aydbT6VFbDQqtBqJPl5miskHP2rrawNhPkkf2XZIh
A7TIFrBLXSGUrKwHk5R/Tkge6Vz06XjXtNYjVAlPPtXsNzDjnvrN+i1JodfijySAmMCd+77ZCH91
Tw7F3mSrJ9Qy42ZraCCHtm1ajBPWj//J98v7e04WL1GrSxVWq6Bafqqp8EA5XObO24+DZvVwL2D7
UDap3QMFFBGSpV2H6xF9wQv+JNmfRUkLjkBD1E0cBK4DlgMbz9Np+xpyiY+RGrHm+MK0MyPwF0wN
zRk2VmgVkhmpmxtV0YuaXw8jsOeE2+JJiA5bHyI+s+U8qkAlyC31rCPbi9iAt9gG2+Q0AjddO3XB
aZlyhixtvE46nsz25H/7cmlGP7fdPDpauFfcR8RlrLPt9u9fKppxVz1oY03DDS8o3kcDOeW18LVR
v8ZoA1FxJKB8uofbXk40/y17gtlyJn8BHmwnT3tRVXnXiAhNN/xwmhpO/RSkuMWNWx3qfmwrh42O
dUjKc4PeKcHCbiRoS9SX82a+8ME626nRNaARz6Avs6GkgU43LViCHi1xuY4dZ2tCDklV/EeRKHVN
FpqBvPp7bvNTyFrJOJN2lfjTDWiq3nBbht3N4T7bsr82Vpbp7Xdpf9kFWQPMWUXAyUz8mY4d4OOp
ssOhQL5+QbprvgfNT44KuvoxVW0RstF3Ribi7LjqrjuqELs5kvgTQpxh2qRwtXlL2BICXWH8V2aC
JuIGMbjavamju7ObgqzVlTIUp3+nf90dCJBooO0pBekKneQGVSQ3+F6Un3/Eod6ERft39re2HR23
BYf4M/7fdw8DM6KDiGwDyNmLHXCgJJybyoODH2bGZN0+p3LgUcNCZJhEJMc4ocj1juyqNPmP0X0c
Z2yLSBqUAsP+YTlhog32ZGm2IZPNMNRi/lUtSECDq1Ul4zxh13sTw0uMKME1MIkjIhQlvB+gYKib
9rjA0f+5c3PLzZCfUP18y3oewz3dakkC8+3WZwgJq87jib0GPN6V6wGc0wn71OYy12UvO+fZB/c2
9YJPVfyuVQV4BDjzC0gJ9DrruSJxedgbUImFKa5+UlrFR7btF0Ma4S5+eI4PnPEHaY1Mew3KlQ2v
ynYQO2ArPU8af2O2JxrJjUMLX/1MWdEy3TeYJjG0TuH5AmyJrQb+PcmV5HvmbVARwvhoYx3sZwQC
dp49V0u50eUl5o6tLEzV1YorLCACkAol4AwRRGnlK8wydso7ZJ0liodsFGET/Ezf3XmmuR5AVtls
7q95qkeMomKg1Ux/r2LCuubnxdNCqZo1g/9xlHoeFvdXunpuGWrCHchABiVy9UL9yJygWMZVsJtx
jT7oZAMYUNpl1+vyKpJMjn8X9wdZniPz17nl4QO1Kb9zv43uz+GYQ9phagdow8FBwJWQoS128HqO
cbYHaG/O0ruLDPiPgGWZRF0J3b6Cl7EM56wWQvL4QlwTmPlrX3TWVhIb2UWkd0i4BoaAkE0V4v2l
z89RDN34TYiNy1GdC9woXEUa8d/gB4JPMk8iqgcPJe57hY7+M/v7Nn0Sv3jh+KNkCHw0Aha3F1Ty
Bi/wmY5+e9YGAhI+Euj/yStyVEOqDEicnV4jsNkCE+DDD7DqLisHsXiQyiHe/F42G6oxOJunBQQU
SSPI72yw5qWO1mW5p2Jx4Xo+BMUB1rW5EPmxUbidQazB171HWS6BRijd5zzq2Nt//KbQI89FcZ4i
PIc7Z37lpQlnu/Mtc5rtZsXd3fwaAAlC9eFv0w3WBGwJ3PsEXJ2TApdG94aR354CapCGTMBK1yWd
oTLWw5Z0Tr1VLDsNUpEWUhNZSQatWkxftgS30qqleScpyTt9j5B1zt36xlWeRd1BsEMUgJtesNGx
gbxCeDqguMe4hxi3JjfXlreegZjBidSGjG0epgT2mPvtLf/ebH0jOZ1Enooj3wYIRGqBU7P5NqCy
RYWk3tU6WqRsU9swlIwrhnyzTpfaACWUQUiCGj2VX2pT98WcE5Jkaw8XijcebTqrh5LL7g/aBcC7
ACyTXWxL3On1U7xgW13ssR4ilddrZQWPN4X5qZxx7epZ8YYu8SWY6eQEgGhhYNEZWWu2PD0eWuHO
WhdRbbzbyaR9XOyGolzS2Xg/ZLs9gU947gToKFaf4JHvDDL9yi7JTAcLITaYAgBwEugQaAUyDYsD
NYQoYmxVcvVghbpwFaeVzEbZ5awRb3xMSQTR6eAPUhcv4um7nsdbmIL/mNm0jo5UcKp8XjtsMlaq
CY+ekKmXn6dG5L+mlkXc5s/ZiFNnFh9mISs/cEz31gJoLZZcHaOTx7y/R30iTNb68jKGXgXxt6wb
apdasdGmZGDLN5a5iHv+EwozvixJbDjJrRafjrPIMIoNwsdQCYu7PfAUCk4pe8DPG+b6gJnrB7Bc
KwaKStcwyGNZZDnma9CrRk1H409KXSWRpgHyr/JXBCKXCqTxXA8H+PSfpN2tMopHS8glYHY4k7F1
811R74Pq02utmjJh/XSQi7TsHhhGkBwjIgaePZwsW3L8Hd62/iwO3y0kt3XTvlGL8l1oRM+zTebU
dR+gAOq/MF8V9fTb5oDMrT4Jtd65xgmW3n132OXZthpvXGDHKH05MeGRxc/YmW+Sa8YqWDXBUJ3+
McIvnxOVRfxdKxueW2ZH+/cgdoQDLpuhB2nqdBj1yhO+jmAwNnDj1cBhGpyF09jTZib2chjr8VA+
Z3TpbRYvn9ybvtwuqMoTgrv/25DBSNVvaruyhpgYknNq4vRIUnQDohk2Wg4afWCXXeTYMT6Mz3i6
KVp19JumsqPjAbksshfMFmjSGGvAPczArV8s/LDOv4cSM02c3Ftabx+PD0ILNaRIEvfGMzkV63VO
whvNALG2MWhFkBYuXCufbkUE+H9Xf5R1jOkLAX4Ur0FFbCA+F9gRZ6kS8SIhDAtncTxlQnqYbj0G
dMERFvbl2jMNUSOjtG0bLY0DBlbNHdlZ99zblfSZHsgD871HxaQLtm57bDpVPKneyK6/I/u2C2Zw
MQlULLPAHeeV/lnYyVozo/9hOdOCf/8HXQeBs9bzSQz+mEHyV5+LVDlSYT6gzO/NLOXNGo5b0lJD
wilZBCoOeJhnyvrI55YKVe7Razk8SNRLSNFhswFkMsNnkx+AvfLkQtklndCPfXx8CnSufTTOXbyy
xgfjPLNVCSWvBXjc2R8MTyh+qn2PIPZiOYfZBc03RTuxVMpSUNeWoSgjOPbjFrstm1SwR8bzDZhN
EgaqsAkUVvGfSOx8j4IW2+k4/JP0CMtJhqXWkS5aJrnlcCvnH4rUq1imRs1JkIJOIsFAD2QfG/5S
rJebnvDWYUFXyqvBivY3bFQ/EP1PcSZ4HH+2ZTEC7dChXjlkItS8eHHQoYL/hFd6cHlCeo7ITN6N
yyfI1OnyenGT8rfou+wTRyH5Wxp972IPAAAd6C4qkHPtBGnntvaud4ARZ9VUAMmLsLVmldcHx+g5
skdN7xaro9r4mWFYsOTGXsH2i5GVjAl/18zoxxjFbHYO+KTMNm5IqVPSV3kLjqcR697gnjY+52Xp
6rL6xXLEdHW3z/V7AQuots9lrXnOrbfIasIT3YjX+QQaO124jAXAKJhV0XrM1weoE0guA2vpQAQO
znifE4Ey0OF4Oxfyt4JPZQCILmDI4wBTm9Ye7uXggm0t4cf7sFL7WsI0+cXRwsfpQvmHBi6jx4TV
tYZnbg/LUuaWMJXrPEX+rfHoeM9BeAYVvoRxvGC9hs6AW/iSAU1gq/6OM1LXMwedk11ye14wMFs2
NfB8+65d1Cj1hTPY95DDAAhcU2eGLpEZKuaKWNZ0lRQcrWw56lHwg+ZAE5LUyTBh8TF+cZ7BsTes
he3NZFSIsZjz28JCaHiA29CVicep1MdV9t28ROjuj1AV7+PGGcXCV8vqYdNsQ0VQcUTCV7GNiTqT
1LsU16xUrtU9nu/rjPG9ZY7hnlNDLdItd60p14XvvbtpJjj8KpWkfR4oMKxUI9NtsyOsT7zGHXXs
wZJOxM3JcGI8q2otXzkat9cLgHULS2Fz3bIxr7G6qbJqCh69O1JU1AvOvud8zKTq0aIGiVEZLzKt
Dk2MUU7x6B1JA4ZrmroFbu6fTt3PxD8l/PvidDiG+XVRaQ6uEbArAmrItDb9E44I+OnuihCpLpMT
z068tGRz2rYnd/OKaZ5vG7cI/quCLch/JJRx8O7CQR7E3J0jCJDf12582DHb1tUIKSMQ1q+4Bsd5
VFLC6zGH6oVxDBJOuj8o2MOLLZSumy05X3NtTjjqM6Eb05wFSkgfukwRrwcUa1+cPU+2D1AlElJC
RASDe/bWv0SeuhJL0X8xP/fx3gVjf9a6q5SGGc6fDIyG+J7Vp9/Zc/6aBsmXKxRSBSaKmx8JYZnm
dNU8bFFEd8Im7fZO5+2DR3lFdq2KHJ8VxK8GUrUwQv5SDUcICsVBM8RL4VSuvRnmT61iRZA4Rr9h
nUJhCE6bOjsPL1FSwGR/spXqryVmK0jpsVySc8Dvay/vvAAzw2SF+eu9QTeBMCN7QVSZpNlp+Dkg
tRaDdtFUQWEqx420E2N0cSeRS8O4YiQoSZG0FmkR/TMUNOFExwAov5m8Y+6Y4KAmHAYmfVdJoHl9
jX4eKF8HWB7I8dkKt+Dfs1+7VaTax2X6HFlAaYuP1qTKcPjEszqNHR6+Geeu7hJlgJigb1teIWBO
V4SS6UzmodHNb/i8r0CX0iM++FVHQG5ZOUzBhCTrrlxPtup2314dK8JFH2Ro1uIW6pBl11OuwkEj
pzeUvQRQcVZAbn+nSMvc7gQMeSJCf9aqpP+HnNQ7Nj61BOGh+adCYNmJyv2WTT3GXby67FtCQTf4
AsfW1QWWTvboHb6p2WzhZusnfPuHSQZYOBnNqRbV8ehrJe/sL1SLbDcQopOVDWxcJ/mEkmZedsxP
H4M1bH4BWpW69Fx6hINPryfzJB9d46Ee1LKTPlU5vYKcu07Vvg6fB6G3iP0RDpPZdy7ebpqFf3ST
ll8jJa/KClTrYT9P1bfICwrNGadiy/RaX6rfwCAMKsZsxxQS3o6yIZtbZKZUgIe6/csdMLlcCmxb
FP0YoIBej8Xx0Gn4lLeliaeSffKlMtaBozkNnLS/Cw1wWty5wWQlvAdd+rvM6Zb5hozFgYzB0+zU
rHZFviwxVnlh5GEt23fW4JU6a3mg+g/onnxD5NSU1TISGdC+KBcpvq338r/7ZPnYY2CRbcjNL3MF
XoD/KSSVCJg1whgD7JAE6nubzAff/1EDx5f+feLWSxlimN1ax4n0PG5/vg5OQHXokFN5pSXSTm0W
V6EpO9d69+Yl2GZCTy1AxLpHmlp67tpGhA6WnZaTrSSrse6wGlSDH7naIY8t5G0N9T1v9MaXCDaH
dMxP0+fXNNfkcGq0aiaHAFEEwBQDuipovYyYepztE+NSemkYkyLtk2DEt2PrZk9xo1IyRZ8eP3Li
uTLfBFZMa7QIB09uEp2LY6afnBM49UCB6WgdF7dsLfbF7hHGC7aH9LY6bFfekPHPSsJba35tjamQ
EJaeX2R8pZv6Jf114cMpWuTvH/TiZsOkJyE7Q71yLK5/yNgIOK0Q+r5dcxdFoG9vObrBM2eXYiU6
uteAs8bLRCi+pXceLr8c2OJbk0O50jmEdClgsrQ18aJLjYEi37RO3P0iLdXm92Lxq8fcD7wAp5hR
Mgz9e4NYqE/5zCvzRtzc44TuEeO61gp1iBY2OGFXnmmVbjBbGNp3Ua+WrsTF7vuXyz9K+D2UrMqG
MBA/RDJAiYaeWsJK5/gCNhWNvtZo6pSa9ufi5QS5gFVEAjxthZF9Vu45mCPdobjLxggqEp6kBv6u
hevt7/LXGhANDa4c3H+aAPLwFEQD1UPEnO/U2+jmpUfmCwRAKluljiSMdyVRtWJYe4LX51Eq0KH2
6myU+9ioRj7R1On/+DxJdj3KLVgDGSJJOxSHHhZK3YssIVUJZtYnuc99sH4Z+yT7qBVSVXN8xDzI
KjqB6aBgFJGdo9IWZc3HAaBEkiiB1Dibjys2/PgB/LmU/S41J4d54Oui3G7UXsMfjeonnppOxFwP
APqmN6I9zLx7FlKDezULID2WNQ2v01yS3OGEL7zuG76DNpEpCul7pTdho/WYPwtUt0RKRNE7xhtY
ECwKxn7bkcgcx9QqNwOgkpR6ffQt5C4m5Y9OfesWNAFWjvVgcLFhV2hi9l6kcTwN8i6+P9UVB5yP
JQHzcVoDEBtyQnZwhNKSHx3K1LT9qDVUZ2CkeTqYtcnK7xijHVHy25vZ5r/m/7UUFo0feA1A44HI
L4PDs0vnm/hAbO1XFciKjtdrWg824wv4f4ptXudBKGgld6/C52IqZ8UC8nR0ORW/RLrFqe4/18B0
U0VEOk2FMRTP23NyuCv+p7VpBtqcSnyChkoF4X1YffhKGIQwaWxSnTkP8OuDV1ChVL7kXc1ygOiF
doejd9B2MvwaVQqnyzJ7vKkgFeopjep9F0srZLfZeFwlFN3Ic8c1quNXXHuAVawCyR6m3ZJ9jlyX
L88w+LsOy17BIylFtRiYh2XomvFiIMDL9WSKI+I+vkzSnbmhQG1HB5DDaG0HPXoTmNSx6tWV63iA
qCdxs8pxmQq2OcI/oJSl+3PT9RejReR2+xOw1/fLc4z8lJX9jZ11QlfDAaTNcarsQpBBcAxIM6me
YbA8LqR5ECeMFHmg20tvDtUZIxuaC5e8XQC6qSQh91JG1UTK3m7xDSix0TcJbaEVawyV3cf++s0I
UpO6/R7HnRq1rT96hCov+ISX3qNd2Swnz918yCgssqRzkWDaYUeispN/3/wcpTQ//iVmnB5qILxn
u/Iuoq7a1uTaEDAzSGj6/oxR+5AcwAgCEPfj6HuKbkk17gzYM87rO+uhl/3xpPOmL8Te1aki815g
lQkjRAEVFhrSW3b3yRB+ukPn83XFFbLH5IfKvDlVpUecRJ/0PpPx5H3MXkHx9CqBZhlFCh/FaNwC
KQEellohLyXs/defcswaCNIeTmcdmZ55DewPplwzpGolZ+ZQa6XrjWNnNJZG+DOAQ3TL903pkwAo
4Wl+tTlUr9NcEjkwPcWjoygbsBDGb6hMzsGcNYqXKpwTjRIzqUc852YBNhoNaJlpkzMBd14qKO+C
upmmwvug1X9ZIR9skbUgLfKOh4/Ia8VANKzxNUcYDhzCqWjY/VcLtKeoLoSKe5pHNxvfCC5QQply
Lo4MIt1g9Pnh3GzV2r68tuHfXYx7N5mQtXc2xp0PUFL95lcW+ydzuvQFRn8/DHFuhfQYB5vMFLNz
kgbs3ILPMsKn+jrX1mwmT1fpHbdKb2lq0cfa3OIuLjMcugTED1MytOQ27/6R7+2In5ODQxOsiEB0
DmBza+2LwYwhU+iSzF7FPFois2R4qyArC70aOczMoEvQuT/ZpIyhBb8vP7eCb7ePWaJz6fZ7QI47
zXVYIom3Fk/y6IVa3sMlHBPy320rhYtQ5x7UOcKxo4iAsrh4783AkeptHHUKSW+OTfbPoij3BF7W
okf7zO6oo1JxcQab4xFv1UsTVXL3VqnVFDYURYEiJvavN8v1OKaDBIm6Rqyx0ReVAZC4QiZcXf/S
SFRJPDeXOAEp+FeW8IjUrp5Dvy6rhsRaYb2v6fPa7Ga62j3SvxD92HHdNpmjnRLHKDOGOU9MFyvH
EtVKSauN0u9LpZr6bsQusE93pLbx4AeXxKq5/bEF0zDvU+lEDNQUMd3kybGfkrB7fOoV/40PPOJv
1pg0kSkl47bv08Uc1jHTj9rSSXrSkyn5oIf03gpWCI5WrccmiR+Eja4hbM4YhXD3hhFnWul3nZYV
V1dBmmSx6iS88VIEATr7STXMx50+WCuQRBkvgxZP1OltMN5fnqDP71o8o8xf0IiJGHPs9ZLzVzKQ
mVUkelyZ8dHBVdgDzJKut3R8MyZwo5l9Wnzwe8yCmZmbBLeeIYbfljH0/Xzm+Gtzl1mCPHEQf7TX
AwY+yWMo/V5uWVV6skcvqKC+gaYhKqyClBTkjvW8DefqIt8ReOk5iEnSxZDqBMQfzCOziaSN5Ib6
hY4429fRTq8Ll2r+jjtkL3LYBLfd+X3O4qe22tyOKj4kNL1uJBUk4PYSWeHjODEDA3og9iggHf/3
qkU5awBw7luRLoIsr8fnlaFnCVkDx+pPJc/CELvITn+vuPtKWQmkYCJUGOPMoX8lcok98I9N9HJ7
GFbf2lnQayJOfTr1NJyvvKr1YxbWvxQ2nyUd4ifhamnL/03IgSuVxY/D2+7jicRS7Wl9kp9b2yN9
Gr4DPXYQJXtu8wYJT4jppa+/2LLXw/jB/Yeb11U14mXNXyXHLTQqiW8K6zj/xKoLC8y4YJZR/FdY
ty3G3JI8BMq2oDxXK840H5wuRj8I+6f3DvyOKnTWOr9BAVX5WiALfQfSekNr2dxbdL9hwz/Sb8SH
QU6P4bor2iyfqmi3imrrA1i0gYX33E1fqYAWPlUBTjLJsZOARpcOl84I8KmhF0jyHRgTOP7esj3e
buA3QR3gtN04WuEYu201O0LGt0WaHzHWUafHKCmXTCgTEq2r4lhQrT9rKLxuf6QGYy+bxbhtu9JQ
3L0dqDjwt5nYsY33HxbZQfG8TBN8eNtpNbeeNz684A7LaL4vAEIblkO0FLFanpWVAgeIT4hTG3sO
tn1X2oZoyxnRqOw3vvcuYsybUynKkRH4k0dotol1+ZdfySjRS6qsYNy7W+wGzI2Lrci5fs17r22X
BA8Vy1jufNS6s/YqSG98aOWGhP0JJrVAg59Sf6Hc8KydBKYWvmil1vf8nQqox9wPrFlmE3s/XEun
upaqsm2Qdc/AI07xtV+vIgGd2s0R6dtXX95p7gIKhJnUA9udDr9sbfWto3/Y98Qm3DbKirdKqMSg
fiGkCpoq4edClQKlTMxXfxdqeeCyz5bB3rWZJo4bBryBcza4W3G07E8RZUDMBgyWI6YY2+t4J6Gg
sU/fv51Lm0Yu/qFCVmiD1yB1Lr762mN0Khbud5JNMCy1Q0+Vrrd0Vc/vRwKi8M8wFFUMfGntNSes
f1mwDzLQZ9FATgnxyaqJn/iDJPWPrpXCaHWd48+5CCHrUpzYXdrDHxynu4IwggETmeHcB2TRUtIi
c76KIOi4q1zVY40rmFcC5I4oeV5Vwymz60Cq8eZNR4OG3gpwjRfymOIaUNcdOSYq+NeZAPzuKhAm
tnSWp4wYtJCXF3/JHJTJ5fgZWnWpPU3Pw5ZeYONomi/dESUjTiakYVOA3JeMXezEyWjiH7v4EIwJ
QuOEn1vz2+x41zd8aU/MX4LpBmdERRQXrXvumpTdhot0TDtEOY8UHta/gIjPaTrUsULDc1Jn0Lqn
uQ4mimzFynqC655qivVz86O1P49vnV8wLkUuxzhLi18bkTSfnIcdOS/PaGcM2+ghpE3Hsy14ZEji
pli7VDPRkF444U0TJBcRcYIiGpI8QPxDFfgojDKi/wV/Tdm3644o2lFRmoa+cI0kc1kNkc4ZK3NU
MiqfVjq8ltjvUi0uB/RQ0C1B9GdHBXp+bYXvBrW+XFW+RTTbjJDMARAEwnwEM/1HqNALmjFBf3WD
l0zlYpv076nvlVuiWs65YvEjRsoD8i7wcfsy04gtBdt9z403QcpBoDyp6C+Mg/peUoDQnOFYOZ71
TIfqs+cFamICa34EQr+7r+GZS6I4itZ+XMUxJmRW7KbnoN3y+om6LGv6CEhD4X32epmZCgtSPRGc
1VzdNMDIsskecTBVwrSwfvReGipZb8KDxglOipqnQTiAUe+WAs+uBHYtXwW9DTG6qdLYnIkF0jjr
5LOldLuWTKWk/zRTuHuCuPoChGLk+7c4xHQNE8KAbkprHLJJ+I02qaqhfhhU0WM1eGkmHT+HPxLu
GG98a/3qUFvhi/0h33ThSyhgA5b9uiSAMSm8DA4JhO+VjKzMbzpR90w558r2ziQLZ2m18sVQCZxh
yUyKJVqzbnEeijS5CHymEliI3zuVcqujn0EyWiMbfOERrcqMfyc59HaQ5tj4XSTVNlFoO47bFbNl
leTIERCb3z3VUtZK4y0k2iWbSEpgmSXbk17t9UGaxhBvul8bUVPZJ5MvTkx9pGBs1PPjYP7N3JqT
6XCkDAPnS0eWe2xRSt3Io2MQ4bNKV/Z3gyjR0pZfXVcOw4crNNlJfcURvnHPotBiuZIxjb72aU0G
xXfpamxPA9y02qHWYtoImSGr4nqryC8MqU5dp3dBTqpEuTzDPW0OLEOHVYMFSY+H+YheynW2Ip8H
TXTMenE9wNy+SPwUVnvyfWzmeJyvQSHivqGCsHOQ+UOOhBg8ppqA0I94E2K1bBjCZcSGQ5I6X3mp
kalhXJH2pTroiiOsPp3v3jkP3+5uGmOxsq30p+/VeGONqD0k+9soR+pENvBBGii+ZDlZTKvdxBsk
fs8wXCbrVeWSI2eJI2qzIovOe1n4tSldfAhtY2CbBmUDlPOIgAI7xeKYcJSHpA8uAp5lUe3T6M81
n2wwynOEAVOHB7mYClCAar9h8YZ6LLsEmu+5O9HWGmbwCZrgk+VNQIVL1oWx9X0LzYccf1rxg39j
VJOHI5Moqww3i3x9Dxw6hBrff90UmVghRRnE50L+aksiLnVRpZOb1jOdmyjSEbBMhX4UEoufOYUn
0Mh5mk09PB7W2HFC26PaKi2dQVeXj2Em4Lx/wDNZ8o/ibDEB/oksAaH7GQvuoUazCfGWvKJ5yN2O
a7IjLH4ihlcXSfo4k1+NEfzNnCvlFxuoproFK47Kxsz7Jjch8Pr2BF2Ax/pZ5SGYuO9y6rnOoiPM
FdUH7J1+xupaZlBX7UeaJNojlWE3r1WS+eDdcwMBouEhzBkLcBmTg/zgvHWGQRKmpuVZ2f4Be1Bt
zuapFHM2Iod2UVNpSIxhs3YiXJje+dt7hSOOn6U4VKLbC6yee6hulz8Qi4KO2aFmWWo2iF0r6f1Z
YjPw6OuPaa4ay1EBC+Vrnl2XV3nLe1wtEtUUegS36ozv3EoVWqdAIfH08+iP9frsip99ViAtrjOZ
DoKDbpHhTmAGHmj9n8ZeNdTtK6NDRIx84VnUcqWVCCaVu8yNpCWgfaiNyEoxChwRoO/5Bo0nMqvK
z/AwUArQCkwKATdrqWuan5DRdgPoa+RGGW7+X9XyJPJLTrLMQF4moaqKlBKOVNHmGOIyhV2xa143
ETfWWd5fo8qdTCVcI9fPmzoMOf4AwjR985Vsl0/6TEAuoV0xbxni5hTGu2VoE5IohJsJlnyqqxRs
3nRgV7W+vRXmw5zA3h5/LUeer/Ku5zz5EEmjmPAT9wcuOumXghzcH1xFacQkSGOboFldT732lgq9
fJ3DbRzc6J2OWShdEXaWPD6XGYlgFTZEhBmydixxhOuqTnZqmkE1c+U74A8jigqCHGp5JEP3OqAA
jqLEEhHlwmVjy/c6Qj+dREEGU0tgwZJsJ8w2s8zmwdIpweyOnyMNk2WWPkSz+incWXD5KznLU4QC
xXo/5Wbmb5E4xtvJyBhFWbszJ69FrU6xTPB/bX1FYgkks593Y1we/7pBkxNektlkRKL/MTyVhniP
BZudikyHLQvtF5NvkUP6Dco3OSc6UAyUEPCPpXtVhU0/ciVyuPWAM0JeArPo6YMg7FT2i1iaNFE5
VAoD+g1uYBlrNbf3n8qqlPp07BH1gpc7VKyZMMdYeHabRgXuDyRpjsrBT1NULh8gxNFwu9NEavB/
4FVkLIlIzccvQC78i1OGVePv8fJphG+JIy8zwhkUyVY9K6PzWTB6R7/e6MayDH6U7q5Fibs3r5L8
0t6XatIggElVyDGR5whlWmwOtzxWLkAlZTwKzsgn0gHjjDrVwZb7VP/EY1VPyAF9Hcmsxe6N+Ctm
TOIye4t9H18diBK2ka/P8+Mlmti2InZR8Ylrk6IU202msUNdtRU9i+zisSu/rKqJLsszmzEvqSsQ
JjE8EpyrK6E2PXXf/EBJMMDmlrhLAfG50NFS+xWIuIOzC9sfM496J6/PMs2QScxFrvYSl1pBMa3h
bMKDwrmfNi3Vfm1PJL/2Q5uvhb/mqvSzfi9bWsqnLLpniPy2/YU31xDdTJSmLjmzTzWU2gjKrvct
y5g9Zxmzq/mWy7jalbeOyHYz4LHtEJHk5tykvm7EC9D7VazTdajzu/2R198gdMiU9NzEkwz0Pgbw
nNAI87Mc9o3MKp2td4/s+8LzG8HxAczAIq+81yJ90qVO+bZDfUPAa+ZF1x12yMHoptxWWygeiIHO
3Y9FR8wwjSc4rPb8jVVhugpCijQF6FmOpJoQx8pvfPoO7TttI9Jrjoub1u34TBRPBQEpxH9Tkt9R
TCsMQ5JhEbK1HKOzFSCjtIELtW8PN9h8hejTzH864NaVVTP9FsJaaMj+cKxADCgMyvhedg7zahTQ
PAufcnSBwYf7xjPfwNhvqxVbgLQ5+8PbjkbXAl+kaTmDjEvsjpGJaRxfyQAm+tGzaOBuu1JwZ49U
/s1wHo7db1F2c3iU4n/SzEKpIayyCySX+Iuv+ybtP27zhoYbwL0XwCPLa1q7nuK7Vznq4sQpOldY
z3YAG1Y50jeVQ5UDwSRwxbGWE/cuH5XlymIJBgWUcEi+DwMZT5BkHhUkHS8smUVcVUJEv56Oue2F
cNDPR8KSeBKen7LC/CX52Hdg2bLgJuQlMHNaC33TAUJmHmCVgPH2MZHknrgprJslEAC6k6iqB6NM
7nSjBCKkQ7nVdEN7tBOCiCBv7CvS8V/OTtnPPW5QsNXJWCtW1zMMjXAhVqhoCg//ZgVK9nIbNbGj
CFSPbV+TOxYWgdYcLEYt1rysywT2nFXTsKyBTWZQJnpOzMzYDzunT/IVZ98mJHFrX0kdkEEEemzb
iNol/JtbAhAHyamZZJV6MV2wWs+YVQZKbVD5Y/gCwHtYwyMTtb1VsCx61ujCTSWKpfzzuZ3Jf5UT
XQYz7xd4pwFcV1JUJi6sO/tzb0+oX/rC3XW9IdW/k314bDADK+uFBV8c8iAj464FuO5sIeYscBgc
1r0zYiWvvsRqxTTpE4tO0jiqMooblVfbVQMuRZBAGyfiWv0Fef/F91K+frV7YGaOpQ8HTn1539/u
WqcqiYEDOWNyxacbni/FnWWWjx8i6l0cY8yQuS1DGEFpuHuqad0dQ1oXTzHPlOqEIOCdfMeJ1G5Q
YJzxDM+ZPQjPop/yFYqIDh8+BIu1PDvM9PX3+wxMdATAryI2SHzu9tL3DPiCrfJ7p1+/AXTCmGKc
OF7r/2y5iZ8pXHLl4aXm6RmBFjWTNbYIRxRu+oxV44OtzL9pMLCZ28BiBiXaNpWF4KFtNO7H+lnQ
Z5Vzrllh8BpjwUlR72c7tbsbnmsDubZhzJiZAMAhxllx+37y7yhtqC4MDR039g2vHQa7pkgGMI2Q
pUsoHqHMfOQUMB68iK9Q3ct6+CPkSAGIS1jsuP/oksEVpt8O8WWhhMosLGBJlmqWFQ4Uk2KED8U4
+Xw/V7dM2VMWmo4ksUkfLPm9o7BTbZlSGocRy70znyTcvFkdGadutBteU3lAr6iNR4DtJXS5OgNI
FBtw+qJGUVpk37EoGTHgojMFy+KleP/btoyNKh5Y7xwCXhvZx+fouf8pIP0+RHpSbVcAVzJz0zhg
NMjn/N8U1zuVXFmlFH2Mdi1T/5fCZZRxzHjJ8FKvxgq98ghN643LJS0UCr/5M7xiTEHpfSb+Re4z
YXx3mxzIQOf0A9Ymeg4xSozhxErl6jxzqJgzL/minzZyC++xblSbNOhiWbLU66ZFHUPT6HGrvCDi
t5TC3VYqBBU0n6DScKJoi/ivGQN56ZSqxg7mIECVOq8tvXr2SCzzDuHG7SsK4zq3A8efnb+RTqAK
zQP0Eg7qV9b2G9X+GF8VNtQuBKeuARB4N/kTlFdsdQ7IQe/zaFz0XVsGlkI0+9ySBBY8i8Fl7RKv
S7nHx3St01Ifiz9o+mzyq8l87ruOqc+6cyQxWlKVi9P+9djU4MqtLce9OBS1ZjjzgH6xcNfBOMGd
EwU8F+Ax4wCilcCT/epleS41qGl653xKPolkgntfFOatPaAToO2Ly1KfPF5A2Jj5j+nWK4Whrmmu
ZVf2pAOqZXet+47MGHmYhfD6sh+f0eTNQgBbNLJeCiUPKcR6ypGqePKDTpRErFmbIqpsXTMvk1Mb
zcFdTz4GgLjVyFjFor+HAxVM0wrzRuzOSi9+3gU4tpPwDR4Lc6TjIcbFEpFYFOxT0Cfb6/q/Uybb
FFYE2YSTGARlzQk8hM9ftTet0cVQeLhD4UWfxlvkB0u8eppgSRPOCOUDqxmD8/+x55W2YXauyqQ9
PVUl55MNPBk6GQU48CwaJ3ykyaE6TSgVRUFcD6aeVyHFcIG8oIJzWumb7aSbnyGoBdek/JOxf411
xAM662F4LG1eoNwSh22TfGvNvoD5NjDHHNlsn4MijY24NLFGyanymZ7l9AuFCilEu1ffo/x7KZfm
ppc7494F7tpd210qeUGvLlr90IFMDGtd55bk0204/2bo0L6BHLvN3p4DO0vc6JWQPUTBqb2lghYH
XoCtvEs/8lnPJwq5W0f/eK48D1YO96G45y2F1yjK2UvXLdfJVFhzzByMLpfT+D3xs6k6hbNy/YtV
mthARqJF4lUL4qbIPmwWNiaOPIBluGE/prZCcTEw9P4wznxu1A9Y205VagR6QAgJQlESNmUpVzaU
qxRoxHuOm6w0dwnRhaAg8mgbCvCpat/i4fimB2QSXkD4uSjaypUWMK4AMxGlCXSJfV9fNtoIieBl
WtMrnOzcq2deKnsIIZfaWNLBpC91pg9CSxwBueFo5LFRB9LPucUjRPj7KFg5OYMma081k7P1nMrU
R2r9f2zDudlU7BjZ9SDg55dSCYopQFvgjEYdSxTAP6B4NxNUf6swD9l5AK/QQdCuLEMfP7n6zv/m
DgEP87a8l4zua9mmI1Y6sq0HnsteekvwSc2av7lyl/rEWIw1o+IfyJaTQQlkoHgZgFhIe3X3LVf/
8e8r+meCmjkGjSljFUQfUJ5g7HhRp9KR79VjCTiyA8UQuhCFjQgoK0rcbjTxDHb2EwvH27d0S1tu
zz+BZpEL3dcFjUY47Vb1iIj/V6Q8j9uv4RuutFX9wcWz7k/niz3Dx2pXWrMbUFkxRKNxxcGO7kiU
zh081S814q7WCVOeKHNd+xs2CCUTxLkTTJ9RINoNs14pD4JWtNt1wR0NXNkUS7OxVzHKVo7+j4G0
/UBWh5TVlHoXcgbd3TEYwiAGQ5gQAay8zFJQsFpgY9nOLtQtE69Xklr4fCETnVbKw0J7Jy/Twyyy
mwBLouL+bBeJw/z7j4o19L+Lf0aS62BUta5Hv4ylFwy+XDmSsMb/sMjyQSrT9LEqxakQkOJu3wMV
TtO1XFEBZ+8DfGW0f/ZwAUk8XNkxPHPJcP4PYeCR0uNwbxM+DqGUsNd2P1reMh/ySsngYh9s7mls
PPGgUHPOmd2sE/rSICQtCdehX9BQK91gNgr1O2sCWiONSbO8P85FY9sPB5AGWNeieQuwI8sFW+2r
UZOHTM5rCgzDa1TvvOqSkMy3Ncx+mystzjg6hDtSH8bjZmGr39kuRIdFwdaD/Bf+4pAawxLLaZb9
UkJpYSqPFS1DTiqndKjQsEJWsL39RDME5Mr56lW2MP6V2yyX9Zv39JFBi5XDxXblOdPhd8GhLyo8
NgY3LFqeGE2e94hZWtAgjzfFvW0FZOQO/zXylzwC+K8yXvrBPSaAp9Vn5oGeU177DLLbxJRPJoZn
tqp2uyNgswO0x9yOuQi/l18Xa81kqbTIKVzyTfGZ6b5X0orGJjGPL2cdDLTYOj5j5IJUz7GlTprN
QgpOkFfKLi5bS/gHF/8TlOYXusLgpv2pm64pm7N7JUgAdwinofadxFVYmvg96FRMbEOziVNU3H47
knNCrKqVdpapKc6wNkCjcwKC9FQaaX6KlxSo2PKWTKocgtUCM+qdKVCvoqY5++4QRi7n2shPlIUl
OgCHE5JplH9UdzNZX35d8wejDbmsQ332iXKe+a+mw2oTswjznolxuG3bhzXaLDlLCGxtp/svGMfM
52A0j5DBefot3K5DbtrYsXePzlJgXaafr4RRAO90t3NyYaCTFkESfGtStnyGmpTHtgCGgn1PvpKx
bclMSrqWCfiGyRSwZ1kPFs3eofCBus1Z9zx0rTYY5g6x5ju35ebn0Wum8hbcoBjQaQ4m9avqdbCR
2xWWfgI9rQKIEWDY2pEo4pgnlod/m7DEUHAyZcplI6tJDWIu+CbIk20nGQTCDBCGJUARnQz7nNZq
i6TQA7tNJHPYla0OV/r5ONcKrER7Np6QpIPhI5klZ48sKLePI4UsXezSGxhY/EiuAzH/V1x1Ie7a
1vLpfSAWsadKvVTYHNYJQ4Sy+npnAsgBrIAYSJg+JHOzzVKIHZM7VF6tNIx6NUYZoRG07aAlrJrI
ptIQJ9y/0VEhtHMHkcX+f2/XIf/mfD9fKBUQ+8y39xTOUXAj3MLAXUczQf2/nJPU+yPzjY4agLLQ
itZOYBVx25R+ox1zbrmpYkuDHcoXftW2z0o8ptjerhoeJZcf1lse8Y+8m2y1UNgp1LZE/wjl7mMH
UgpzRnUd2+fF3HWpLIq6ic906YcLiWEPrQU1D8xT5b8eqU6Ph8EahgjBOabW2XJKiEv2GcAh5uX4
u4+fMqOqlIUm6H2KB271T2gQ0NuDwGtI0Kxu1X17VVP6OUdjBchFPI0QhP/hSk5NIrhaENMgt3fP
wQE6ryVvxEv9W2SpGDB2gufwmiTt+dVXVYRic7q9XF438zKwjennqkq3v4ntHuJwW9S5H/OQ6cBL
OjD2HrK8UFkzzZ5l3Rv41OnPMSBWHysQRqacDz/+8tiN/sIMMFiQ/Lzoynqnpdga7ul/WihU35TC
HDATNPqLZgiYX29q7EbWbaAZp5c2dW3WOj6jqeL6QKCis9aQwvr0y+7rWJhPgBTZ2Nq92LDM4PBa
S110Ne/BgqTBUZQzDOqazMfCAgY2RnLic0CmR1nolVfxpKqNJS4g7LExA944DnsizJkIFu5ATsnC
R0uen7UVBGAvYHyszQMIx9CTD2PwmDeEQTNnn3HAbV7ZCCBncNJVOw/6LoHQryhlx61YDUxZT4BN
y4sBYe/x6qY4+bmHGJubm4Q64wzbIfWfd1tXHrKKaa+UA6gPr2LzkwztN2I/Siyn61EbNPxuXGr6
6aAkVr3xOL/b9YtWgJAUuxyzkDyZIbsBlDIzIFj0ki1dB5C1VBYn7nqz4/T21RsIwsmNG3wZI9KF
aLso7MgfQA1UbmTRGcjYv3nddN3B9ig5+aIna3pEftZ+5idkpLloNUeaLnWbqnqgQKIYJStsNziF
IGrwDI8wgJwTc/TtrH4VqKU91rnbZctmr28bIQFNEF8CLUbYrvGgH7VvvJtOsHssOHG6r5OgSNKc
xVDl3lyzjQf67jS2ka2ZydXOEyC3PG/DmwHC+PLz/oPCYMDk84bpQnlt8ppCnWa3xAUiYt0DWQzX
zHuFa+yAReOrl4Cvuqgha2vY9Ma0QKV70WbdNzmiMVg2WprTE4epr8FQP+WOXv1Htn0Evfx+ZIzI
s0YMbLFCFHsOrDqEHKIZS3Zvt1ZO3cPxNk/XTbBMqrNFqBss6zPV2iRLimo6tV0/S7qIqm3spEjB
NWB5VFW8tmdasw072DYqAs/PrG4HgvHjEjuIfX3/TAI4xQ8IJT0WHvU/cisYkjXLREI+secnmDV0
UzcJrm83sKsxfWy/Xrt22vpGsy1KgOKUdR0NSf/QxSGflXIs6D/AUEtIPo5RanQ3cjCbEEEv3R0i
cDsoeXXmfsX0w+zcFmPn+zUjFm8Vzd7DOEafckMlSql7TnW7CFaLNe13eFbmI820oRVkI2Jhk7bv
ZPNzZarhG0t5EccLyRpTkUrKEaxDVmLcYbRQi2zsV210O2bXxaMh00VrtbqX2hQLTs3hRoitMwMV
dy+gcYUfV+HfeaOLf+mVERjE30lVjJsC3ab6xQW7hUBhTUkmOFzJYFLFoK98FzpIJW2V6V4/IOOg
N1xF6gr8Gs65P61sbjR8Po2Mc5du04gxTwWVfDZRtACx/AvqxnjwRPZh76ZNa+1c8V2qZ6b/LM78
WAndEtyS7TBaWSuUrShzKXZT9oIzgffzhWaKIG76oJxQaYVtQSVf6h/PVtHzjB/fcf0usFbJL0R9
oMqJa9D7FL/5eokoV274eZ+OoiHGeEBHWhWuqIeeyeVv3vSBZd7vY7RPLxpklxR1Lub6yhF386bb
U41zVhecf5fRbaqVatFUaN6jCzqqxN8PTLwc5oFCrLpTX2N6lJjs/5DhB7kfgG9asPPgoF8fiWrF
gGFr6ssFCyBHbwej589iLwzKjTnduXAGItxx4IYIH+H8V9629lXMdD1gKtWh1iLaOdHfym8F0hKa
z+24FYlpVe0YW5Q/LJCucPW28aQA9biTfNyBM4DMWmbwrFMGxsvyRhJ/JLTTHA+p0+3aazKLFzg3
/5nf1Rww1RY48tQ3I33VMa9yc2lOmNIt3GgAOvtNdoRHVet4v1bAbEFtaZ+BKMhuy+PyjebBwJ8h
29PIx85v6txQApYq9I0Ei33qIryBwU7xslQ6Qc5xWSnfqwuCtnPxzB/z2Ys206sLVGQ3xvUUElw+
32OhoIIZ0Oe/uzM1CNBS1e4j4jnjSTOqG0s7t+npmvhDaF9MAT+3eiz7lIN/NNH09C6bkLfrJVdu
m8gqXCx0cABpX62a5SlkxqRcwloNE4k3nHKfyDvMX/LazwQHY1pk2ykBXKILzxmNF8K62OHUCL2E
NJ4g/QomGnNfoMk0hyuF0+AeS8gSCmjma+nrwMt2mysy+8uMa/xZ1FmSg59LBHyjyNKAoUyhVQOC
sEZoyoVq5pM2kDXY0j6//nbis/iuCHIctPt0QSVFZyX6QDzOtCURiPKhHpQ1ovbsDEC2g5vmysG9
ZJnVo2Zkbr3V+omFD0nMTzArqIhsvPaUQFFUfce6bVKDkHuISiMWFkHyPN5akxLcCBV1eVSc2490
0rJkWcevTpxItMqlrO5M+MDm+PwWlom+PcV2GgEooxXFDJmm+dmmnfQwzy5IrIgwkeEr2TIzCMm/
rWx33A1RFmjaGu7xuZUk/HL4zi917ASxryNoQ+SjxrJzyRqdcN/RHTCOgLBSWjg6RMEFREy9OoU+
bNkMQB3ynvLS/fJ8xm/GFRjJYCC2VTMX4JnQH9j1FaGf+WzQmWudP8e8nzM5PC9PKQhSQd/g7894
EdajpTQ7k2iYs9wHYsiY00MbuLaLU7mRcwJk9M1Ft+O1XccflaWWMLiMuQEMkktplJx5PBoyU62E
/MKngABuoBb3j2mRDV/BlS/CpBhhHRXXDaNtirqf7R+vqVos+ov1eiHMEmNdUImuK8c5tUl233Ei
3KKUMrQfg3MWT4AW1AINoPAEVrmgbKsTCf+fK/YnW4uS2V8jSXAuwJcLdnN4Ylf7awFQLiPINnJt
kCrYOJZ8TqilTOfYH3VytXWzSOAXUi4+bO/0gdJ4ZvhQlUYU5CbfmDZqqpFA15+SsR3M1K2BvAmJ
7RdRk1334eaf/jn7Iq/7K6SBLQx9v8FatWKEN3E7eGNi07ZDA/p1I0p/UluzKpykBNSBijkFGd9F
W0b9OnzHfm2WPjDuaVgE0wgCn6ka34MjXn1zYQdrvezr+XdVcMc6ASlOZh7pYni0XQRf7BKsWY7i
ea9fEAnIDt+a+G3bgujjbvlvcOPH6nqaUAx6cubOeHZW+tVUuW9UpmH2t9OoPZ2+40bBYnrl/1yF
yOty3txzgaHwVz40p4oGTRROMqBF0l565Bfr0t4N7hCE581k7/ei9x0yGV53qwYdaiO4vFZb9TgK
8pRzjee35fcqE2nIgG1Mv+xSDbUTt2fyjko34HkoUK6LtH9llYfYZXQ8QisfdCMKLDGI+aw9Hyok
oiCdrSs0dpjJhTSWRjIgwu8k7ZcYF+VJ3nSPC8T9+3nbiy3hFle2Aec11tLIcLGvOGkkfyT/czYG
VOrZHzzLI0tF6rdg2Yd/MNuv/U4HWxd2GUyCwQVmeYsOU8QmnITVU1cqU/Uzz7MkVxfGIZemxDJ9
z2J1VJxlmz56Y4SwPNBCnjP8sdaNP+vYAAjf46GJb3o5d+s2ViD+ZGZlmOlin8bG1QlUJInB1Oea
tzH7Odz0to/Jhj9tGb7pLACLQdLuTiS8zVVdtTsXc0wmuwGcldDMGwi9YyY/CA24SW1S+9ERLR7W
n3cx/6LYUKYGS5KhgZ8l062siGSNnbE1qNvvI+vMFAHRaVr+tlyUfzEJybuRJbAtbgMOsTj76DJa
qpedF1aC6Lk7nFayt0OqUI1siRmPGwAqYZSnUmCNljG0JWHqULbgqDfyDuSQLmEZi0xrqKwS0ttg
YGHP0hwTZ6rqgae7hgyCizt+NW8ZSjYfPDlmhTITkCdaJgfAWSCUXBUTqtFuklqyVCd0pLAN8SGM
p0T3r3JuyMGLOu9USrJP7Z39ZPbNEvOgNv7z8EDz34d8aa0pyS2oqy5EDWEJotOFAwaYaiKi2+3E
3bVemJjPGaxSqlW2z9TUF3x5cGkJSUCo9QoQHpz0rk54rJHUWSWu86tI9pv8whBoSaXxFwxqjk0A
fyF+lIpi8hjrZiWtzPJcgVfat+0xGJei38MJi5O1PFuVkItwKQwAPhn7JTBf/Mh1WysX1U5wpyf2
6RL47EarZvqEr7LH+1JcziiZUMN+/8mMPeSuFrN6e1E4rH7jObUAcp4/IUi7iu5l7/UoZ3sLvPzN
rxAqImG5Qw9nimUTZ4GcYeErAR5XZEsBFdwMU2D6erQLj1LTdCm7FRQ+wZSVWbpoQdyZc1oXPNG+
vCtlYJo+AP4x5fIFhY7ElD07HOVqIRP+YIzkHqEvVHMUdJSquaycjL6EowbiJQi9+3hUgBmC4SbT
9UO6vM19kQxM7zIYFSuSAcheAlRuAiuYontRlfcdSzZbhOi6tjLbmuv3YCbcGUEkX3XYIOCclIdl
3yOtCluwTKtbqOFmh4sfnAX1hSfOFC3rcfUkW7ONDchLKLP3OM/wi17oG2V6HBY7CBmoP4n5M+7u
+GrKFliGZ9or+tavBrYFYyR6I6ks8zh5arP/UCZ07mOJv7fcGLrwgXkYz8Aw4GPLYrut7rUuBJ/s
w+5Z0WPU1fJSU1pjzXQ/rxeIjfkFzwZAMWkkWQ0GXlMjPvsDwKSiG1kVJlPYC/Sq27iHtYS66GHq
Orrrwo2KtrYgAg1MgzOSPP/RlXO5RZ1wCmgwKeSH15BISx5b0qwTB0VsX2Df/X+TN/SO5Kvwv6eq
6tRdYCmc7fnV31ISMdiyjsAdpf3K/ZqeFUAUO/Ya0bh+reXgNhQFjB4+Gk2+wmVHP5E9Ia9XtT2w
tSQuKoGXASyWThQvy1ib26QBLcr0+MASZMkOzKuKrE3/ixi3ikEoBfbXDHuIBJhs4fQ9CQwHn88G
yg/lRfsYOoj+Kv1v04AzONQpeKMly0iWXKKmCRkf7fZ77+6XUu5fSR9JJft0CQ80Kqo5QXAu/ISi
7I1O5yDSKxD8D2+mTTEsiXGVGPOCt346PFIocI8emHrn+HUJkk/+KT2jjzxVF9J8Tph+uubC/6Lh
U8dlWpBruKgnfVJiZWhbq+wium4mkun/BUcbG42Po8iQ/BKTI7IKcy1NMD543/GERUF9l+V1TQvT
0ztO+4u7mlK50mOBDxelyKlRWek2C5oEJ7JC5yCR9DivpD296F3V9NbD2E+4Gu1p7vjg1FV2Ef32
XXnaN76r140viDov59sxQLFyV2Fr3BpIXRAtk9trwfVQwo5Euh82DGxevLFWSccHYnu5yVEmekWc
lAz0JXh9xi8KtbB145NmlD2Hldsm3NuvbCIrfVFtF0PO3JiNryrk2qMw1J2WlEMg2ftbbT1Q84Hj
eQ5JvWc6UrdYpZAhs+9fudmMA78vNsK9+Bva429zWbn+3SEjc8+fKQCojs8upKvyBA4JVuhZ7m7u
dgXTVhp/rEzpH717mODFcSRp5gQDxhUU4HlAKZsnoDYlLjhcnC5IsYhAGVSbvwNoh8b6cpyugtXb
lorHvkzV2rVfID87BphaChozju+KrmfHgM4iJAzf3jQ4Rwk/VgIGHNCKWgn94KEb1mzDzFb4sfnk
FhlIpxOTWRHwTV5VowmbTNACQeeRdmro/VKEm/fuEcERUR3l8SuSIxXPHYBoIxy/HS5WShABAAsv
u7Wv0fbx5ZdaIWF57j4CP0yPy5aUp0twULLw+OL0x+pZjf6LaDx/iENdypuBZF4IaMfn/L2vflCO
ccsgplIkIcTsoPMEjNq9slr1e3yZ+hqVlZgmugyu1d5Yng5Q2ToVs9WxDRy8dOP3yQPOaYRCnjFt
3BwG+RNWR+5KsVejWDaFl0udOLbnD8tCw9wKHJJPS5Im8Sf4Td9+VOrVhhQKFGpQbeHZ9uDMGQn7
GaWImOVfRsxO2bVpxr3Z00OtH2aLacMoBExtVUneQ1WvAXn1VOuK18MqHm9ravAGbEY3BJm715vR
VVoGh8rNXoBbaB5nTbZQQrv4sJ2KD3GqDAgd9JVdqHZjp3kZ3yUttYGUuYx+hC8gSuR9jeYXTXLy
m8wyDd7tHnTFX/HY4UkohMbtiVM7RipH3oNt/OmphNonqe+2BeOizs/z3KpkXmfTOapjUIS2juTm
QiH5GfzLAytNePF1F+RgMsfxa+Uq2AUiWVtMe02JljRe3lIjCkBC/pjau/BkKZNs/9PAmAbYjShH
LW82PdpL+qNztJCvEh2thXKP4ubADoL41D/7MvsCX2Dw5yW1J5YqDKrvliOAiR7i6pYFCnaPljtS
rs41m3j1tGq/e1tAeEsqghs2MU8Vr5iUFeRqXbmoHr+iabO12gPDmbwO2Y8UYNNuSEFjyGrvVEvL
6RH0tsDYYtoiwgCPEDCRwNRAW1CklSPf7lWnZ1XLSHRC4dL3FHJaNDNU4OWt9QDgQZIEVbjhkaKg
oRqShBRnIsEAZ9NuzrHXYWx4tabB7wm+2jDTr9PryYhfDReQz449H3ANcAJ8kn9UvxcycCn35xnn
IX7Y7qkfvqxF51LJSD5B/hVzKwQD64MI3WJw5JTcoqzAw4aU4Ac8ZM2I8X68dHeem65/kVqrsBwc
ce93YjrvZ7lhFReKkY+Qr/a4P6qD4Y9AiJaGND2jj4axsGEEW+E15GAfq98kcSU/t1eY2Mn/H65f
hEnDQX1x46c48gbQSzbdQq3IaPV/rLQk0x9u+hEQB94om9Y/hipNPFb71AUH5QT4R3BUzAZeYwsA
vkAPTCwSocQsGrR4hHcCwcZEcmC3NO4QcLWfmHB/v+K1ZNRCVxV1VSw9vXrV4Qfs70bf0A1TbPn/
jR1UVkYSNEKgfoKcRB02hJl220Nt9vp1lXpl2cAtYsbL1xf4kdhD1kYTGBl53w8HuM+M94ihUPDE
YOrQIfL1vhIyNYZxGFKIb4sA/vs/wI667GhWZ9F3p+qbBxqnGx6Q8gbDvCqdHcnmnrihqTYAI6Mj
MotGltf+sVNVWBhytibatEPMAs4yFFm6VcxPI5qeOHzOsOLRpAngsr2q24+tVr2rktxBr2PbZv6N
ZYnrR4jjR+IwnfGsNbQ/pq9Gw5O/+YqteGxfaWkXpeMsZRzbayUhr7qr46JhJu2UbXTlmHAPOLaj
jZ3f+NiO4xWHeLQlFHyQa8oXxVzSSxkr69f1Bt8OUaK3hcn/+pDSIf1k7j0UClNU/iqt5jNnTtbS
Y+gdqQG8RUtKzPfBVhjmMfOfW1iJSR2ubdXGWYRJjSHxLOL8ApcWi0gX7gSgYd4oqeqH2tYLRE44
3J9EkLDVMf0m/Ig3WJCXTQizapHf9gfiWJMMWMmSHG1SrZbWut4Z02AbibcoHl7ntODAMn0S35Z9
nSYAmMshDgaAWMwxPmeysUeofu8eWiGTo7d4nyR9KIJcXjblKbwZoVClMxC6f3v4lH11On4FrJfx
JgIf1Uzr1XD1F7TYZzX7Sgp2z/3VGtsazKdGOhXDtJFsMNmt4xWi6Yjt8jpU3Tf27WBivV3H0dDo
46oZL2JAaIB4HXJKRn4J5dps9phn7U259Z7+XdUphy2LEuqulTWTXpBofuY1XmZHMgcaQz9m6++N
Mof+D4T83mTURxquTXktp3VE1AKUdMT9scqyYadTP5PhhW56LG/Mmtcog/ppnN6s8KuZLtF6mbnp
Y7cGkP5FMIRIVPavPuq4oqGGyMNxGn4RzdHe8yNrW7frigBs/vVG7RjZUzYgtXeMtdSg0/NVYRIc
wmalmuiEcxSNRBRi/O9VWNty3pEFP80L4t/uiQKKgpTaZ9F2HyMw427ALifZMppz305Uhd6Aihdq
W3qqBNzEDglJIrLmadVNbgWQ2Yp3FTbiDbTc4c7HY99CMTphnvLYM2AwAz/G5fthFfCsJSOKIr+y
xZqc1qIMF8Ws9Lt/AjL/v0PKUzARzLA+yKnlo5nEE1RbRaJRC0lbVm3L94/+w6prP4jaafR6e1Gd
6oP6dP6/w+Whd6dFX7RJXWfGpHkfCN0hgGZNGmb2IUVaD9U/vKPtosi4f2dGJRKDXVTtghxjBZRv
UFic8vHvM0UFRDCyjORr74Tb0uL3+UPnTsUKKSyTUocAHzwYvP7O3QKHL8V49ezLKCV9XTcQVhuu
xF6bo4htSnEwKrC3RKcvq+XrCxqlDZwJgmc5CZtB6NrAD2qA4Y1c9/M9yfZ42V47J1q2C2rX4qAC
Kjo/U4brqjr2eoerJ4tv0DZJMhNZKTmotlJYMWq+ddpFRV4zlJTygwHyYkytWwxRtcpTb8UxDG/N
Q8B4o9/UF4f7a9p7YQqsAgm8w/HAlgwgX0cb+pT2OaN+lItzjQJNuNgjmuC1oVf4RX8m1eJSEkpJ
67T7kiQb3RdBunCxGW01+9pePoSHmiG+26D92xkW/BjbaWjevoxekRIXKRKaYGOUahxo04hkuUd8
n5vbHv7Ohjg17m4s7KwbQDa8kr9lCszsgHxH2oj7ZJg22YJkZHQzohqZOoFVgzTGNS2H6VrBARID
TNt/pk8BroixFjkPRfL2qTgc/nOhTaziaF4+KhRGU9GTdIoyeIOBSgvkEjfAtNVNBMg6QROR/bJt
I+bRQVz8DHFlTdr02k+n4cLwdXpHxBG4vHxip2mXEbQcr+OL/p1yVuOVb0373K8jYGT1mCfZQHK8
Eg4aQ0WONe+1PtYJaT3N5ATvEKsU5vmQAo5GFHDRFisvqSXHFW1GN2uu8H+7oR7Ee1/tuId3JztF
3hwTE50s8Wx2IihkqYq0UzD3QI1WEPCXD+VF1mmLtaJaqzaGrBCHh1zowzgiFb+XXe74gmtMl9HI
QgFUbzhtNvWbFXjCcgDdVHg2FThV0eOuvyi5EErFE2pYyXWlDj+up7P2meG71tkmepkhL8dKo/+i
yqjFkl/vDOnVr12RPjk00HXyqtTEiVbAM81sHm7d93onMOJ5mPsvJ09e5liNzDATgGWH2ToqsFoH
gywm4EL3RZDf4UbMy4Pz9cd9mpbaIkYUvV2ALBwKcrLqHHHWsn7BtwFEXTihSicBtBPoh0M9mZOB
5ENnXuxL36s1zQYtty8s+VjAnXNYKNGjIIaoJQdQShsvVQ6gSSy1RmKSxDg8S3B6euOBz1gXnYc1
6TFkmfv/HNCjW1rlWqLIpD7YGeJEE59Drx3QbJ9sPi6yrMsPvwYTb6q3hsSNFu4MJVbah19ns3I2
ADQukDoS31J1ryiwWoTMhIGJJTwjvAAQu71Y5dSifVb8KGNv/BgkpagNGkhOQTPhed3R6jslol/D
XUfRA2Pi2+tCNi5jt4cYtd8q0ryPKjRGxtzT+45FhiQPBiKhyxd1kNMRywi4HACftbbn98nUyBcx
LvWFyzlVPSd59NoQrFD+7i64qFe/66RcrwaeA9BXuuNamsrW8tt8s+uwlwZ5cFodQjXJTDRzwhWn
uN5EtfM9RqttH5xEoOmmGjWgX+8PIF0/aqCRCp50ryoUPGw0AyYoJV5f777379UTx32cbQKKMoSZ
22cirqukeP1Slf8t4P/Xg8YZR+DbIc+1Imszqk+x3cC36gienZZY0eN+JE0UrFZYeR8gJaJkYXWk
G7JfHjxyN9isWkmM2TqH+s+B6ZFosxZh2lvxXceYqmgU7jS7lYq0ZUqfPQVwOCU6vyD5aWgGi3BX
aKvTFFWzGycEv1SGnr4/wSq4MYrb3NvutD+H5CXOoDn46kXJztAHGAhVOKZHm4WBR+1NLVw7l4vD
cHGuCZWXnmfCKqTxB11HYP3J67eNhbDZX0nschhjA65K2+garFLu5dAgP/OKb+WD3UI064ZlIwSl
9jxQ+jqtligv+gCS/g4NZ/FogETYhQ4eYzIViC903afO5+oq9TADSCiJisFV8I0Sw7cWM8bcwy3Y
twnO4sEaI27YZdK6U7OKnQdshOil7vK5EZvMr95Ja5eNdGLQzjeU2jhH1ZEsLg4f+uDMyaBCcfbo
gCTNBP/ga4/gmSySVcQQdbc7QAXUYtKn+P/BAjY7TvjobZAEHsNO0kowC2S/ERUqtqz3NSLSM/US
XrN4RUbGEOvt2hJK2aBNB1GlkYi9oUKAjUwKPQUamWUO1p152jIh2EZiEHb9eDBQGPOgie7IiXZW
c8WD6Z95byTSp9yhesRJ+8EPWxbDA13En78M85gIixsJBUNVQOHC9Y5lO9ESlcWzl3n1DJiEiULK
MWZJhSP/TgjEQEdqDKvXZXjM0nDLnMr2yOTRcsX9AS0BkFGnImPyMeCyWXqL4meCVGMrSCu+hFat
UrTuAIgKug89iFKumoIqO0+tA86nqU4EtsjEwZ6XERScJo/ckPCXEcMaHQZ4GCIgX/CCsE5jJ0Tx
4Ty1lIJUaa1978g2Uc6F6AMo4xuy2sKmE5Zx/SmiM8x1LoWUk4MkMA6DI1g13uo2gLXmKeFtpOQ8
Zlxx8hfzloi6ZCnjuUvrhTRdmPunWof+jyWsIu3U1eovKO2G37O2vHfZfmTshOIoLcR7z7nE+zol
CL4Z+0CMmRHUJSrVSqB7kbHG0eHkIOEqy1AMogCS8BtRxnRjc/gSYu2g2HvUvcq+OJOEeVPAait/
e7h738eGj2697x7+fHkGPUSO4wqLOYjyy7pgLSADMoCLqWuMnPEEP5swZ2OcayKZvJXmPBWKnSpq
+1SbdG+S6FRHTSsJTkL2CKZv4jBwWRYUqzDpeuTByYagFeCpZW/l6go36toPvmN+LeXnC9L4z295
BnaxPhpQKbdh5rW5s6OmGgyX+0JMYZzaND6vMD9VbDCqDVDlhJJjNBszl9WFifEKqKWsmDh1AB7o
kvFeE1djYpzc3j5QVChQuOdR/eNlLyRPcdPs7A0oI+SDqv50KUwOZbh8bs6gMtogQCKnxLVSIKFH
dT2dut/n9hKAkc/uIuTKmZ33mFMfmaAf49LJ3piy0+UU/dm0RE+iz7gFm6E5HO5vFEO/RiTyp6MO
KCHyYc2nspStwHwSKp1EvvKdO9fF20xHDopsb7bBAqLCoGkn7MYTfKg5VVt9fBwlK5zFGz8Gcar2
pBHqlZ9Ykhul7k3BgNDB09iCLtPlzjS+TJoxKHPVWRUaBmAQ6E6P4XOH69Ese9UPnO7UhEdS8FFo
I7ZFgnD/mGWI5xR29GFmQjF4VQDAlAq1CYvCMiuLTPl0X+rcgJ0pPvmMPkt0s/DmuTmnTa72ofiq
QwaseEy0KBak+o4iNxthJK2CFCS44KnlFarE66GLXy0lyXV3dtG+RWGfLZsTqK1kEJ53xzAxm72Y
Otlts825/ifS3Nxcnb3dwRpiEXw6QC9+C8a6K2ifg997xSU0KnggB+WGQjYQMbhC7Gqa6Pxwl5q5
gQNTBB++s5tgjzaMhVz8Ql0624s44RVTpym3XXOnIZx1BL49ysC6twMsUVQ2sE6ciiInYo+BW5Yj
tuG4jXnOlq8bvyNb08BdHnKVtI/DgQZbGdYkBRnBoOp3I8KVGlIfAUe832JjGPb6QdUt2w8gPVtA
fuzR2tbauS0/iX269BR/OVX1Ous2iOy1AEnJss/AG78ahHiZZWiOsfSyRkfYsoUOXaFuMLy7vzJf
i+H+MEhGUR/z8ypa9KavR8VEo/OP8/Af+VfAk2ESpvGKDUT6PxOvvcqffGdP83Vn6Wqdi4HDIWvj
uJBPCfH9G//eoHcitSqnp5LBUx2JD+nV3x/jctZRZ1sK5EYFeQUT01ShIkuE86hDqy7+cpIZOADn
fT4A/4+GpYUFCHtTVTTwdY1/uoVdZeVxmKV9Pa2uXvX2LFE7a7jtS8uC6T+YU1/FO+mG8GqpEEJS
h9cyd19KyBuxghMnhA69Loof5KViIbeAQuNkSRsMUzWbsTYh6OymEcxK45rN8aLv9fb7eA/SW5rP
v6bzO6RMomHjS9Hoih/HsasRclo0OIKN4K1RtwCjWepVVfpAGU0fAXllxf1Bz5fQiJuFgWQvqWVT
N1Nhtxhf1PKX0KlGU87pvGhhxyBVA6kSOQshBz5RpWOQ2D/oce4vltiE4UcuvuD+Qxuu44WhEC4R
L0+RgJcY88DpZOJ8jmZuMkWlstGRqNf9ihhAwNqlaeoUjU8xu9yfsjfSINdKrKQ8lsNBTYHJ4h0o
gVp3KzJZ0zcmde1t7L5q62QYZ5pHfVqux/Tsdv9/Wv4mAjKCnpMr4YU/3lJE6lZxseIitI+hKAWJ
c6jAQkyUwe99tlbKhQWkrEZYYTEOW00/zVwspf4jo6DE+D8ftBe6pi3Qe4A0alcFNCco3CPYo6+L
5USXlN0HHa1dfc7HH8Qz1Fwktxhsr6bfksowMkSrnqcsmtqzw3LPLKZFDTr4v+HaK9hzLL6MRbPi
iQwmOnVsgadlyz9yCRb1NjCYK6O+5eQ7UXWmwAUwzNCmd09zd92FLVzHM5Nmqaz0G8Jz8IyFk6rU
m0vD6mpZHVkouQfdq7tCU1jYMZsTIDe/H92zlx+B1HJekVgD5Yuv9Dcgymz5KzlKLPyKnMdq1dvV
67tDH/G18P/uZEjKlHZ4cRC4myik9AP8R7tUF984KGFHVu5tDQW+mXoJ+6dijI1edZ2VPnrtjqDu
vIv/L/K8knXI0MJccE8u3O1pdQObgP/k6WflJAAw1B2f2u8ez4RXcwS3sMImoQavIDLQtKaqOEgc
iFG8GLdni8dNxDgRWahM81wwidrGPJelRmUXxI7Rv3NdrWTqAgGiBOaC3mJ1r6EpufWOnwC63K9A
DKZQwBtvxXZUMGx8x01HzhxYjD1UGDQi+z0TLyKlRdQgrYMtKKDk9136tvFtu4GT+E0vQCv/jslp
lbQq6S13Qsi4Ojp8q0MKJcsdtgCbhhqjYyvhh2dYMxKq6FAyOhIakidWwwTMvogyzMPkQn+0JxMs
+trLmhZad+wHeY5pjbwlYcXKk4ALbPcRs1ZE4DmMVyEBVFOYqhfTcp1QvHC8oqvCic0clL0QnswK
4yhF5JwriXJ2ENDHPu/lZ7OwQbzp1hjhqHZdr1qqXOczDcFOxq+E0uVFvJUbS13nR1sO1xDWPFW/
DT6jhzs41WvWqZqxpMIgF+EBlt28h8a/7rdT9pSWC+zfzbn6srMzoySIpiN+t+TABWkgtw5AWPm2
YxzsHRUutO8FDjAyijFA1WXY1QnopYQrYJ48Ms3aNnD0KVUVp90d5gOcKuVjbNI64lA+kn0U/N+X
JXOidZvqgQORJUO4rUkqTgW0NDwsQgEkL1JLQhOsyL/RySkDn39NV9wxF0fpWBkVTdzH5OPgApQ2
0dOeoQ0GL48SHmabZTYPyQ9Yu8RidIBcNJ0Gj4TinCnJaMA/M36KUz3iSvBJPPJU5loFN49h+8Oh
4eqpvol1fnUEWSnT0q4nGDJxUdPairIvicqOMVIAcY+MBGmeVDTH+g1HAZsloJvB9oUpztxxZZIW
Wdnv2OldANaNwEP8qHfPn0WjcHu18KVjaW/S0f/UsfSz2evFy1v02ly9VsIvO6MdwyzmkgMjGGJ2
BMhF6fyb5dcSGHBFqX/qWVxGkHZEQL7FkKDCaTtq95/OhDjRuvpuGrtcfyBn16sFNCwOgxVUEgPx
np+V5pA+Z6VPQvy7MRvCRv0iCwJTTqrGykF4n7JTg3/do6R7Z5KWPQvYMZdHcGZuFezWikOILsYP
Cit+vpDVBm5m75w45islKHsX4mIbDGyGgxnFwnNraKfg4FMBuBoffpKTKtzuMlLPDvSl+BL2AOrK
mUl3y9PAA24l7E78QT651KtmMUVH+ojrquY2On+qBXUVJn51evrpUgddX0+KAczh1Xqu0eILxozY
PjKYglsw50uqEnUQ8aQnGNUGtk5k7waJk4vlOL9yLRSsYJo3n/HhzQBmHUJJaT/htCybPMrzoXgO
eS806p10GmWrNMzbJQEq396jgA8jQ9kfseWWX2KRojK8k+FM5712VR8HgthIpUuIdkomwB1ti64B
HOwVvObt02TYOjNhPkb9bg7ByfzgO1VhgC/rEmnNLU0OZ1JKkWH2bO9/oxaA2PcXiogRBlG+ecfs
Y4suglAAC8wvIWTwRWeWLs7mKT+MgtXS+KPiVwwJqTdJwz8f5EG/8F62g+oKma2IAGDJwhg5TmdF
QTuPkG7KrFhi4eZoRGizdC6TQ6FdXA4z5WZLMUPmPPNcHe64MyrWcYuCNqiBuRNvU3smr6SJvR6k
KumZ7tF7MeaP86V2BZ+j+t3FuqQMOR3LjQlr8yEQD6NBlJKJqAjdApbOysRKN3KLvAb+nTv/B18Z
ipRnyLzvRy8xYTzgfyUGmwbezgJzB3n88TanHo5oCWyAl3Ga6RfcVnsypcpJ2H40KHg/TBw1IYzK
YeOKk1YDCyYl7cgLLvWeYXRwBMUWy+5XIG7PLzUGdSO+eF6jb3q1AVGYpiPgQ/aJvRMZ6SGnEgOx
IjvxAE5rR+KnzZPSQHPbNFvX4Svvmgmr+Rp4ZdPdteA4mSNzZ2DYzWNL+00PPADqy91LPIRU1wmn
mMeA81Z3oGtZe1xZLhOj8ynN0Go/vnvadoZIwFog1HA/vGE0AqNEAC3belTxozEu4HUP9fCj2rIG
bEfunRNRbu0utD27WEJa0+raqRqRpJEb4+/+Fu5nKWlpbeIaBkb9eh4WuRaON5i1S6ZtzcLrjff5
0ujspr2zf8hu/ODLhMmKwGKQw4f12Z/H3zGEH9DdT5q+T4kUx/z6MU/23MESovce5Tp/bDYEcfxr
zUj6+psJgHX2piqhoiLGlZ5NsadEV9xZFhRk0nRRyH1aBk0HHBV8yq7Wrh59rivt6w3JmjD/dvz6
EjsHj3UtK4Nvc9GZHiYK0ftUbTSLDVoUbqboJdmSSjwpg10hwB7AJ0RwG2ez7fkK+qJekMvO9XDB
uD4M0jHu/8WgU8X2Zx72KgJhrLpMyI0g4J1/j5sLL8/TuNBlJhVtqRfk3nAWKrAQIUgU6D8lRrCs
yWikCqU4Vom/ZaIqgJNqnWy71vDNeFTiGuUW3FsJeOYCHBD0cMiLT0eiqSMt/YbIy/gcRgz1/kei
YLCGg2Ebp49Li0rJYEEZPrmBVD5rsO4i0GomYUjFfNef3F3cevgQX2SsHZ4QcaUWqKou4bQSe9gw
m1Z21Irx6q187C+LzCOgG3lozIyUZdKiPiu/SP71PrEd4yJLL1F76Jwfj8K5hKAMr/AxuiFyoVXN
fpGFaO0PDHeOZcAK9M5DcfCxXg7ky/He+kqJxmpMjmR0D4A3rV2X5xpBTsN8NdR5CTZKrHOYWzN2
P1eBxGGOgZNseuz7Z9PC17SbSmXfv6y0HgNYSh7KmiINCannMmmOr+GUvUXTiIIEF1umu9tFZu+z
y93Wm7ruvAg+veHoVWh6zBPg5DbaWE8qyc4qzifZ+zgfJi5HXAUaWAVsGYAag2I2IZqv/L4O5G20
TGaE/9y9gMwRdKodEhd56iyRUOfMlXWSE0cHhVONoiELsGNYxGQ5SXRZtA6WcCy8H0ZB9Y+C9AW8
LUfGY7Y1kFv4obGEEO4zQaBm9h3QjiDDAW4ukiFRoYvf+3X4UHrpcyMZUdJaXGaBFfYgNozbrdFx
NkMO7XxrYYTzW1AprfcOs0e9E2NimrSmTRJy0snF3TrmoZgxBhPoNNKuhRmVMpVwtczpoMfMqC0h
gKnPzCv2pvufz0CD7vSRq/aN7LC5amD8faEKRIBFdzACD6DLe/RVMO5kUugo6xrZAIhU1OZ4jC6f
ftwXfAu6DdWv+WqD+jW6xoffzlHvOaFygv5xIEMIRdyIMUTFBXUKLFLFV9ZjF9v4bCjvI8booQdr
76cCyXfBzrECYSphFUf9sTdYvL4uMR+SmQ4mPgjaHkAJFRl9fImQZXyPy+tE0LIsYE8nHEoGB3EY
s0K7raFipTCFX01N++996OsCQSDQF6qtMjY7flBZgbqo7WXJHouzsgQNc4t0y04SfkPpYpZYt3ZN
cyGPuALNDhNPAxzb35zFK+OSVPXqjX/9R/yF3CZGnNwDEp88loDGNeMAKRYq8bxotg9417rkSD2Z
Ypnbe4/Tm0AF3yzRb7wpm+elUHGl52zWsB5HU//QJKZLmThSaBrg7U258EWP3croIb17IUnGRPCC
DIcbYFlpJZ0OCOLqA65eo+LBkcI3Ug9mzTn784QBEQHcyQhDGBxfw2RrKEg0Q8QED3Y/dLs4dsAD
X8GPXvXNibIM8laN+yt89fB+iqz3TE0nMej+v8XaUnKWiHxjDWzktSvk5x1sxwjMjemcvctfC9av
eAdqjWEIY/Ji7vowufqLsKSllJsi3iCcYG/Csngmr0ZtslxAXVWWv1Q3Ut4tfOKBG5dLPNqFFCdv
gIK7nNw2MM2u7mlyOBa2s4ULOr6ioEvNPn7m3xFsKfgackPfDuultOp+hAiUPR7+ajPF2lACXJaz
QNhNDPQ3LP7uCpWmr80tEtMy50mFz1RmK1PA9Svs2vSoeFzz/NuyPvYA2U4OTeTY2rnHGZmAbuIg
7/42Kkj1IS51Fmb27Mq1Shxeaa14DT8MoCd4oej3H9ThAVGtyHCqq6jnLDCqw3d2plbDpAaKd9Z8
7lUtQoCMI3TVb0BWFB5f9dLZK4tU/3esTmq/tvZOdhTO0xRjiOwFBR7fpOFgzK2MXXKs7+9sS+in
AgvD3S9gImQr2oHF/mIVylgqZiunvtHN5P1do6uOtM9G4uV+XUTBU6+WoMWmPLdnvXByzYK7jvOw
znNzZam+bSakbzLV9rFcgsyXlYrKbLRZoN0L3ZzXsRSDYmCouvInxm2kCVvDCHqEkxfy0eq1Fc2m
KpwENIhz767DtN9iXW1sfO2LFNIC3ioQeQS0c9rAjn8BX57JgekwljTQZpxR8AyDOi+5c43l3jS2
XbkLcxNlrN+w+kGmJos+F10DVGBwJBdRIM02Mn1o14Vh1PfxNQoFNn8DMBm63dhPWhDM+KN7fdHU
JsC6pQWYp8dhIMRJZaHVMYp2H7jsA7W5F+rL9Jlw3O9IlRWRhSbE5JPxDM2f8gXwB2FEloX5NJaf
s6iSCeQff1JfHErtfi5o7O1wFvE7sAYJCYq+6qt4zs+cMUwVF4Pb4Qz6EZQSgPU2wp+rq9l9nw00
yQqAPvaL8fGA98mfEspF36GOuWIAJDoqzghnphC02svZX7LnZWWLVB5g+4jNHc0rmq3igiVNHlJL
f8+sUrDcOAPc0fEyMWSJaaXMww/E/ZmtRDm5MlMyibKxnmZUgrTUkBFyckKsMa9sdv1JIIVKh6yw
DIzEE7UV1INSI7tlM7+qRxxHgvjtbJN6jkZX1Vbcgk50DLLYkKtzOkUeujx/nSwNsCCt8jlMPBbj
gpRvUSipi+FLJHO50azTPPTgCFkzSsBnB56XOJdXzcLJtzq4QWdcTrN+jqM5IUIr/X4udTOKp61A
haoibAi/VCRZ4geyTUqC1cNWFFXWG3SPQD/UjOBx4BeSJxI61zAY7qJbWqQfKMZrq2vI2Q+Mds6F
KSxZVxpNBwUKnTGJKFPFVFvxgz0ZGxlmbRqBwG2Aoxf/6987QlwBD7U9+t/6jgrLR0uvSMrt15Fr
Jh/9OvvY/SDDWaKxC0GWTYlp8Du5pYldn6yBshLo378jiVpIm0mOG7HLfZcQHCcE4/soaB+ntker
svsWHT1GZLpR0C6TJq1DrOhj6ms9Jh+YDAeinpmIwuEh5AhO99/4JcDKizHJGgPf5ZfRV4Z1rd8y
pWpNjzgyLBDATsqJEWn4Uwe9soR/b4GZVmuSTBZaZvnH/rQqsYPE12o0F+TFs3pUci7l1lNTGieZ
sNVDPEtBg6KGwMUG5Hd1m2s3pbVwLk7HQ95nhwRp1Y63Ak7eSeCYJSMcbZu3nBd4w3Fpdb7DAfbg
kPVwUV7dRNOSMdSidzaLhIOciEVkuFC+KrF+WqxFfjVfmQX8hZwtpeRKUUzthofVT39WlAJVe2L4
9S4r2Jn/WG4WN0g/TsUY60Pyaxt14D4Z7O50bcq4USeQqjz3wx5CJsNN2QgKePI4Gigqd1iJksBO
nnvhfIxm16PF9y4E2LPG0yZVJpN7ciR+GBAIRX6dQnUJV/+4hQlfhnP7ASRwfATcyoHRCLUMv5lG
1sUGf/G+cx5iw36tjwNAx4EnoPekAkMKykOPWyLGlLASv85T16e+GuLkcB0G5ZvfObMSB1HX38iF
YPrri8jofJpTAutieVRx1fTK4AgH5lbNLNxfsLatTBLM3P1/qBIalevr2mTV6v5Fy/pcCxNS3y03
LUROYwvA/sd2X4OFU9gaz7KAP8M5VpKoZN0Dc2TJw0rwKPAVPz5p+X40RulVC/P3WmLrKRYQyg++
JSodMLbelCxGvol7vdkrIy0trAciIQ7IFPtHYEX38N9o7BJQid8445p/8liISP4VWNoMXjscPK3Q
PtG+yYBd1LAeDXM4tmGNQYwLTUv/3bkpur/baNIsVOGQivq7+M1/JCGgbLS8620bS3N4Vmn3U/9B
r/SdQCsBMdu+sWgR6NMNA0ETqoxbY28DHR2Rsdc9hxaPqLVwOXtp2LP6Ec+Eit4jBGNv+lVnBVAw
avVP8HNnLkLgWzp9LVE80rbLLLnGc2mR6KEwVh2/IrDlTfqVS16/YM5FMAzwhW0knh8Ne4769Zk+
j9e43tBhl7CUgcqVr4JXG4o+fMcw64FcQXI9/6om3odU5OTdMQn/2viCx8zFVdvxir6oWUW+m+q1
B1pVlABB8odPd9HMnQXMC+ZzQKQbU9pNIazjf2Bt5j6cYPoNksU6gF/v/H8OBmjigIXu8q62EIxO
XFYK1XjJcdQ6sQTzolUIdOVTSsGs1wfjFBws3W8EYXStZN6y5CBhTr/9AL/XfpU060sk+4yFW2Sh
f4cwTG/TDaqXDkzSjrmEDq72k/od4p8M0hh1li+cWieSlTYHL8cIGjQLfG2/y8CLp3n5zr5MWKSq
iffhr3kfufoqGD5wf51ZhdlUqFPT/KFfJSkb5iy+Tzbrz5s4+SuqOpSoy7q3MVbrpuC0DC8TmynQ
Do5ii7zBogwIBT1PMIRTdV6uTCQf6rB9lt4fPQ73xhzv9P86dSi08yRVCQbVuDV99tZ4ov9ZbKdh
3F7Pl4+It1HIwa04ymI9bZRJDt02TPvqQZHEgu/bonFcspmVFmHtDG9dI6606nI3a/ip92AWQFaT
h7UMThFs9sBFsYFNFHmQjEzDrSNWtdBKjcBvymvoD/4eR5O1KrFuiPE8ZiFUYiCiQuEhdUsEkt9P
OTkKXX+1Kjhc9JzX/KFNGFfY6w2Yluv/vAm/3NQiJNZaWI3enNMBLZDaXZe2BxEupC6XgSVmlt/C
fLYwiPY/HUFS2+yzEBzs2IOlYIVmFwNXM7XaCJIfVr+lEF5VkaN7zuK8zZyS/QWSieWufmVXdFHJ
IlVJhLDUhU9V/dRzNt/Ixy0kn9PObwOsbAPnXg2FEA9m15iDiApo5Fenu2jWJyH4ZD7bMyVdj1yy
Y5vFfO+6Sj/fr5+Z5pUt/x00qJiTF/NB+vcc/KE9Pa5aDLaLXoU4GviZ6EGRfxMsoX62bQ9zhmdA
KVe/HQCiyRdrZ500yCHN6U4deXzW0HW3//EeOMehcUdq9FXdM2o3OZU9JSvOq9JvedaEVczcpsiC
k+ffFqC4/q8KEUI7Mrl4PV+TVCg592GophgZj6g7Ll1fET4Kx0QUw8gqKm/Qow0e43buTFcxh2gM
RFjoS3HaGELSyHvdKNVuAGSK/B/7YGWNAbHYJMcleO1ave7MT9Da7Iy3+EEwquB/I1LNWQEI7ttL
0cuMM9q6ixtMqsSBXo/Coa/dI31YxrSr5coByvuuNQJK4xZEn6HH+SPaIaTJI3xy3uezohhgtGl+
7b73pLlp75rIwd26ZHZYCx1ALOI/zTX/GdjiMdXgeC3Z2OYwfh4C2A9OywSccgV2TtVbQsoJ5Nlu
Q9BIm/fMJGQNFltzoqNdDgGQpbB8d3MDTw1ry9KvZlZsfbqPuKyjFr4b8Vi2Z/cPjZCvGiV17OdP
UztTN76QazwDa8lQhouYtW50knS5DbNAqBGs2rGknfP2N3bogEr+kJKE2OF6qiz7WFsyB/JysQyG
hnOGKV2PWAisoMJDHfrer5E6BSEtp2KjnRe1NOkfHBTmffb81Vze6RFreF3AMr54m8iX4dVdqqz1
6LmnTeJ/hBAT+OIhyhQpq0q8uvW0PXKBq63klFny9UCKs3xQzt1s4TEnsU+d2BTykAKX8sdmwz1N
NGthv1jlgD8ctwu8fEAbgLdTjiotWAxnXh6wyHQuBWgoRhNH2eajJSgkTC3oJvScntoUVJ0sPDwU
P3C0qQLFkkMDJOhUY+7I3fcy3//EpgHuK6K+lVJulHWXxlD9TeyBYcFR5dbtGM4R8fz8uYn2gLcG
GyIER+LBc/RohWzZ+4gN52iYioQ8xFWqF85O7BHwRq2//OU0IpEhFTQc/K4W9YcuiOoEc1RXrioi
CPpOA/75JH21OkXP7zmFZDyYd+9IkypQyEZLO9qkr788WYLMP0twRnNGp3EpBzjepCui/2ea/FNz
ICMjAEBep29OrAI6gbyZxeiVkQwzTcLoKV9JPHLOkJO/Q1CMXJHopPkmroz5uXNuA8RotEjL+E9/
+yj20zCYHq8wwtYp6PbGiHkvocT35Ez0F2Ib6fCPPTB4X5OaPCHYvowhU6HnQcTD/zyxQiwH3Crq
il4oR4V6cObIM8y9bDqU6P5Otoo2k+LjnAUjeFTPHzZ7NDzTXqWRa2XHZ4YMUOyJN24OsM6jBcbS
Kc6pJCQEzIAeO98IwankKUJt4byI9VmfQRuYBtBKdAax1B00zLah0h4PKFwbAle9myNThmVQqykr
4BH16dZEcIF0SgBq6Kb3mG3OVZgcofUb66h+5hHPxGahkmlEJv3z+bbyZ1PmjmUHzfsfF+pv/YEJ
rwosOATs1kFA9Otf1DpSyK/HlvI3Xwdof8UK4N+WkKCYRuCedS7DQwIDULbPJvfSFUfMQth6DrkO
XvjTjScnYiv7jwe+KFPBiWx8RU4IsOV+mISrie7DfWoved5WubVwpBLGwrEOF25Pr+fZpxD5IOZC
1Ss+z4V3Iu4gYIVtCS31CmoNw72ZjunMM89MwTKHFdj51lcFl2r6ez/ByM8gLyrigxQdpm92H7bf
tmryhl2xWB/Lv8CeeoK1P21+P4ilEjHYVwW1p3b/Vvi1F+6LfzVgm4dltplkT9q3wZgSSLGwrwjj
w0Tvs+sWixIOsJq0fLgjpqv66zJ/S7CepRyOj1Ltt0DXvW6ZZvsAxYJeI0V9fXVVvcoNq+ZnlRNy
6VSbYP0vZxgSNC+evoq4dLVvP8zhlhEmlc65SYiWWJIy+mJOmvDmutr5qvfXLU8X0sipWRm5ojkL
6zhAHeO+EyiwvL9kYoWbUcOvzsKPyrq4ddTkQ5jG43eauAua1TWhzkhS2cMv/FsAoTEoBOZ/rhcM
3gwY1BQ4umWus8oAYnYMvXBrzqyYELZYhiJQzMDuBgGn3FvTCjHoz5XDU/tnpAycaznaKPWkBbdY
Z1itTIUemygFEuNwxwRbuFZtU9TLkbEvR3vG0X74gx/ERP+/ynFv9H7DyMvg2/ei7uKjafDYp4Xi
23Cp2RNkfdzhL2mj0aYGfEgcWk0P1Mt2Dbe8IUmQQC1OECDkjMukIoPbABh6S3Rx9qR9pnE6EFiq
VkKdKUbjy4lR652aBYp2/7Xtgh//cqFmdkRQ0vGQB4l8T3iGfE/N4r6chbBdt4b6nORd3t7r7AjJ
MoOIHRawuHwFWCl0TNZ7lWHLoALONqfcztKd3/8kC1c0npQ6mEbe+mXbA8FBE6dsZnZOxBBjQphy
tkk9W3v9QjkOMzPOhhsq1PQYCAKF7714bKPO/8gHDD84CkStuOYqpCgaWFCCLtZcU4aT5H/xdcI7
T5LhxZT2pyde0KrtC4VETAXMrOLnmXxWAg25grlJl6K28WdD7+kII+cYp3gtKN4ftBO9Qy7zg7BC
4zW1DqiMEOfkJKtlIzNoU1rAy/3RVbTqzBBsJ8OSraaEsxMOZnaeppusp/Snwl+cFzvxW6DQp4qS
KCYWCAT5LWJ1nEt//NuQ5VIZkUxvp1yhYexedF54Gq/N+dnrOCAcSdzKD6nYTmkzagJvEpCtDFhj
fxlF/sSV/9fy/BWILsqgthHjcV27fEhi26qpNgsPz0L4dQ752bzVv6C4VWsU62BSO/hD6lndpaog
sXwsM43Kfaf0sCb1v0Pc1q9rnSmK7SsyC4k7hfvilsycWdSElj3qAxmRHnQzlbDRZIWxBJGy4Ped
22PunPZIYkAOKSn2jkxuk7dFaDcerjYnu5Nv6EBkEh49LJgb7O/b+vB2T43VsPeIodt5mn6WLEe5
nuiiFUpgcUMvwCuHp92jEw5rljOQnWa/eMrK5UR7+/8zBjUAylQl/fxl8CUAa1iotkh1NyUl4pqh
w2sPKGBShZMEjBG7Bv0/bFfNzMxVrgpvFS7NI+2s087rR4V7GfKtanJcx86ysGKNk2NAs7vFiuP7
sF62xs8h11CCn7UMYzssDBSehU7Cieu1PJm6ebGXRbbyZzKwzaZq//BB8GGj2nExfs2fTKUWw6t6
ztnV0Jf7u/JO08FJzErY2yre9dyasXjBh32fhf92cOfPJyrY+YaRuBFHhcKwjcziP5k5XFI5j892
0u9GmzM+76xOCWFbJfUru9Dx8lYk6aQY2zU/uui7+OduiRZK85Fo9ZnEzyFsyZ+TzzMBH3lj/Ahc
qOgWFimyp1EFiXHz0xNiQkTW/xt0bbKdWMaV01JycOZoAFlEjOHNTd3hItlUbhjHWjmsUqD2FT/Z
XFpTsYJpsRFX8b/KQFuTEluaD/lOBiVUiU01IRLjGsEwmkkblfFgqMKWJYB6vrDhyjOUJLRuuGlw
DgkMcXZCe+6bKmLqF8IYenUbl0HZrhQqc8Y4ZV9lXScSZvwzMq1j8R5aICg3p1PZKajL5WUFCq04
haQMJtH8E4NSPq9tSuCEXMe7sIiLWmv33l48vMNgfgFo5Rb4WsJvP4QWs5JbH7YXA6XQZB49SfkG
Cv/cZa3gXNItgKEq80US3kXbtEZK1zDIQyvFh4qb+VuTL+hBiaPKTTgFRhtUgFoYIk/u6LIi3S60
cmflM0t1ya3KW0FusIgv0fR18dT0ZzO3AA2ralCUhh0CsSyqtbRjuLZrWaVG9oVfK0cTtNEuAFMr
P3rAeLUXFXgCo5NCcBelmjvlM/WCIbF0EXPo0kMvV1SEzHwR4p6T6l+KlwErjJdsGp45E9k0W9Hk
YDL/Cdm6pP/crWYneHhizB3mO1MPK+DcXZ63vy8v5bSx5LrlfWY164E0f20435HpR6NlBtns3KfH
GGdu/oY/cx91q8vXlQpY4ORHlBdVHC+VLN6zgLSuGyZe/CXNrg+JR1UazH1C7gJ2BnfcKFZHxvnE
TvPdoul6uqF0g58O07dY2iMPTGZuNSTqybEtUC8y1RdiW3cgZeov/SrAMQ8HKL3FG+J0WolBENaK
jIfdojLm4KW1UKrGYGDVVHRUV/lbHSTiUAk3qRVhRKyRSQovJAPG3YKPLr9LMCqy32Kr8g8ZzbO3
0UJDqWXzwIygw7sTGhi+E5TBgwx1+F/7bt7K4d0z7xdagkThXTiyUa1mEHnS57jWECuvyqMV3s8e
VVmRy9/qHCuqvJWL/joqGXVrfbR5oGc0a9/gresHl0920I0TTX3+sf278gbvJsO5vgOyk+o0sDRx
mtmTWTZnR0GR4jlmjcFzslp0lm9vGgxQn8jDYaFHpiVC9FEp/bS3+VEe373WArwqriy5ox1pbpcd
fcX9L+0VzvPMIA+aWTtPpYG/tm1FJ2u9sP1BTlKakp/5IxEpN5m3BrzfUMAq5cZCxUjX/PGhrq5+
z317GL40aCm+w7JYXwRivFdJs0jYOWgeWPWzm/yXu8x4ofin3bBRbRlDq+CPz8PjOy6gIfBghEZU
75ljjoTgHrCuR8MNTEUUaI+IbloMkqK5K7+nxNgy3zOdxc9ljL5v/3zc3CT2fbLTUdmXiM3bZ7Th
Wx44Zv46JAzntM8SyLCPg3qLOymahXqseNpp+pLIZu27eApYDiBkUHWcYEzztw7qeM1Z0+8cBxF1
lc4EBFOsO5GEw+LTrgbOAxjqpsJn6Rg0sE/TlqzNdyr/fQIiS/Lu7EoZ3u7biwAmJpi5CuMqVYbV
FES8ZWjRYox81hEfcZAg732jqaQiVJtZ7z/yq7jMncZ/V4IwtIpJMuZZ327eDISt8rmTWUNflEo5
ctDhdbw2a00LtbFOQQlJ/zevV6pr69VYXMN1fRPX1wds2HWzTkRKlr6du9VF1itSvrlvAfIvUw2R
xELpv5zUdG2tM+t6Ld+M79C1SvfeiYG+eIDnsxT6aG1UnXWMS6Hu/0eL6RuSrvLbcL78zEWO9AcB
T15dFFyYSYVOYXFcd1NdTVBerR7ICNtcSy2MT41d7z6pki1741Xl1kKneZZlPiB5a4YsfoLwZNTM
RgSChgzYJRY/xAWgV4yk3XZeEutwJxl5ihBXcV/QdfwUBQdpRGmKAiv77O+qPmmqRPFBDJsnhKis
EuwyxyZSr+bIG2t5py6rNCH1kbg98HgbE8BMi3bKxuAyHOb+HnYdlbvmvBIAQIMLxieGCi1kUE6Z
fH5BIRs5txlQ8Jsk8U3ZmHRVjk5NIv/PMnuG0QrezWYqPnLSq/XpMPk2a4P4k8IUyDc0HNBdRUwk
GeaksV451hLUo8fyrtTAoW7BEugf9xVz82wLhfxhORKRUpdPtWNUQaM8rdLe2wSWQYKpJYHR1YT8
d+pGtW4w0xgeZa9CkxNgDYESbxrJ8fdGSgbpvXk7r97yoyiOYyRpNFunM2YbA1lJulvuabYjQisr
kQjcwUCR+VbBuBhPzYm+62Rqc/j7h1B5aeDBkSa7qqisVH/HymvmKbmwDTIW7zZVja9WepThBPvk
tdNNaZfAc9XbFBjagc3eS5EfH7YlvtahKo2HxSJQYGMv6copV0iaYmop9Xjv+B5IYdYkJO0QMOGs
HnsMGtku8I8X78prfIc+XMfpr/enuUvi9HrbdUOVm6vWVKGyBXD0vnjrbYXjqxgj+n3pFSsb01PV
EGr/SDq9WoNOnH/34r9jYSrjpg/sVA7jycFPuYzXUqAhO2hloWppN0SFGky3VjElLz1f0R7v8+I1
3qX1bFiFDJnelcc5IaQDnkfvmZEBWZTJuKvPmlmgws8QUKsOxTJWQYyIgy0x6ExU/VKBbkxqW1ly
fcJT7vBLxq4HxRbibq/5H8SVxpVTZACDTTCGZZ3XrLAl9B0LG6OoKMKpTLAlk8BtT3U17EGyWKN9
ui907lIK6rIM9phZbENx1c0qB7NOzbZKNV+/4VH9UopNlu9uNkk3ioySYloRKzxFZFyws7bTRPLT
VBgrGiKlSr1NNuvRoH7RH0kPw5WErsvPEQHWS60xx348awggHNvR2fd6Kzze+n3xgM0G1Y5wW9nt
LBrQxxKXh8SQtvluHta+RQJcVFUZ+bDI4/Kx3y0kBBAceC+3DdG7gUcDVKBE88q0ISviMNFhBJit
nc8Qy6MN3jh2fSZ8sOcdZgvsueQa6pjEuxBX2vD8kjrHBnt6XTZ6zwTtOo4Z4jSyxPsWH7Y6/pO2
UhVckQuBT+vOcdJRVj203upLelwHvKYdthMjnXus4dGGNrBV833DztkAkot84I1ieXoJjmbTsxpu
aDmjOz8ewBCqe+d1L3MuNKLb1M+ppUh6mrihJOeASZTVbQ+WZNwYkh1nOwOUs6muVxssMssbCXTz
pblmW2fGg2gdJi8U/d/UwO7BMh9SDjgCPTDU+futl5mPDbQD/EVcJjd3UFF5cCfIntJY+Ml6J9Kg
TreVUxD9BuZGyKr2m7ZF3+XbMtk56y4X2EErO569zG/5kU/KAXN1No0u4Nl65fpU7P+AR3lqcLsb
Ip0HIKawLuRxSxmZ7fr8daWxPXDn/wJNcq0FxJyIqt9fLIMWzLH6BlfjUHX6rtSKh8WFiNwtPDYO
Ddu14yzW7I+W9MdFzeS+LI2oEtEt6NBF8tAFQVgfdPHUfwYypy0ZDltCDOYYvR3ts75NGxU10098
vhUm6vKXB3wg50qdvchfrUtqv511aY99h4+jrvMrLiinHuJfHIPrqoY777A0FtwtVpGNM8k7JZgF
Dimmg0Do2A4y1pA8G4wj5Xv2xeE3o/FK9YTMK/sQzQa6tF2UYg2zfRxTykc4ykKhuitzscufGAZZ
8AnmsqxbqG1lYv+/pxZiv/K17tl/p8T3HKhKsfVIyJ3b4TBYIasDUN8DUHM/vox5Y5snIVV/0YR+
JL3AnNppC+mrKO+cKNS/d81VMNpi0qzO3V5c+wIFOiKp/1WY9iHCkQRVkJURyXNrwJNkLbtK5EYA
ebdWV8TWPuKTQdiCda4wbfpLZl7gRg8+kK2bKU3XGlCLprSf8pnySwrHALm1D2whjK9URwBmrjZC
SiG9maFfcu4OQn7hEtcnpmWMOtcz9DYtg7V1uLC1gwl5QeiU7VdetNLqMdn/V2ahlJ8eaKCICiP4
mPEI0cSv8Nwhz0ZExiSBipdMKczXQ8YcH/rMrsUTUR+PyEH3CpZlud9aY3U/lnk3+/Fp3aULHrKr
DSYRuC9vDMC0X7lAweav9ERi+X2tOHadhOfjM8ptEit5PmYn0V14K2GNJxAwFvQD2UbK+MJsVVE5
sa5kkQdCAe89Wwz1EHsINqmEgzlkZBh3QhLRy91gXGtOiELoe5W69ovrjqFAaaukSpUYLrkzW2F+
ysuF8kH73yqhD8V+Z+fMMWHQolWP/7KidDwfVpYSIpa1b4FzlUbNkdSxW566OYneMjfMIo9BqgoY
U6Pc4jmzihsDIaCySlldJEhmebM/BN3qtQfBaLuwy4qmUyELDTUWaTV7v3n4kDBwMvHdIWDFWzd3
SkpxXCWjO258u+jwEuZCwEWUVzUrco7bfsklFcY04cZgGZadFju7gC+ZbnD/JzvDLBXyI/Sj9Xas
nJ7+tH2G165qeWrue/kDCVr7OLADSwluasoAtISYy/++gLZWRaHwCzkPBJn1A3YNDncnENEWKWzc
kaYp2WGHYhjtcdr2WsCPp0Kob9ffh6q3cG72r8c7ttxElKTZXqxdcXLse0XhsOQRlu2DaqR7J3U9
Nrdcv5sLuQQ++becAS9DDH190cBlaKMUO6s56UB3trbQNY/UGt+XbdYv0P24aW+1lqECxiFS+yRE
SpDXPFUwkamFEVFFk3blmp0BwtaLfiTWh+c86zmb9b7ygxVdqSphe+XNtfugvzh6OCk+s80CvC36
G25pCLjqWAv4LR3X+8KudP8yGsGnLvhe0QXexv8UgQPnpFM7aaH/T2eGDgoy61cTZNflAEWwNCR9
VBCnMJ32g6euG4Per/cbXmHrVsggG0wwEYKY373iEvqVD0SVFY2le8kYl5O7D/UjTeOgyqWxdmgg
WGMr574oH+mxNKBHJJYkHmMk795QuaCKT+sAPk9t4Dtvz4g0r8I7SBcG6VAmtiNi34Nsr+8YkaHQ
iIiP1AUK+L3+pqm/k8P9Y98KJhLz+kvB1HC5Z/jp/fSl9O+rIsIspTq9kL37NMisAPpDV6jCOtNq
Wn5PRMx1Ikr4PEKmKTyop/xHtbm7qaPwcAbQonSLIY0HNpSyE6m9bj/frzHmuWyvUG/qQSCgycbd
jQTcd6OhCUTPl1cChTX94bV9EReR32aNsCoQn1BA3riB/HpPPS2ELJgkBM1hJhBnYGs2NhQ5dQdm
NtZAIrkmrFB/by8kR6suoQTP3Fo5pZ7TKaGo8s88os24itvOEq4nwQ/w+aBNGk1kWxO7oAh7G0DA
hqs2/kTD0JQjjZaqghOt6HIoJ4Vq72AQa0XjddJ8NKyjPXw1pGwVLJm5Qa4gUQx6qT4G9ibFvr9C
JkM6O/bJtmWidQI28p/jXsPCCcthXIUH+u7UhiunHdsoaDivD05W2D5KaoaJM1wAiqetu5g0Oq5H
0I2EdjgTJOukc58l1vkfUrHGyRdLtt3CM3Kd0/sPk/pNwd15Nb2tEngPvKNaq3nDJ/PAFA1gwjtp
h4ID8+xUht4G4RL/Pbyz6N4Hzbf31UFcHzWA2wMe+iuukWFl83mIPLiHuuuMYG0OShqSsLUlNy5J
CWgDLgVCgVautMKOzSg+senwcx6+fcaevKarkgaudh/HgG9V4K19sMyOr+g98HjdiYM2AQ4oywZF
IDyUM+Laa7kCm8WPewy/TOs64smWl7p0k4lkUEt8cYD434N0tJolHWgeJZCzb1HUGVckgZxL4LgO
LuV7M79ZOcenclAc2ZAZYq90XlFQ7xg4C3Viq1zwx/JQ0BoEEwcdLIm8rTmd67hSMkac4ijnyTfA
DC1WdENzpjYPLAi+3OWTyWtMtC9c5UB2COpLFEah6+yWkydpZQ71D8xdCtT48c5aO8kSOUtYV0+4
Cf4QBdbxiruIZebhs1Wex/OKdvn2SYSaRRzc5hWwBAeU+AaNGmRmGa7S6GGdcxJh5oOEHQs4AEG6
fTbD7aqZAQWnfSBU7KWeP2fexFiDNJHd9IT3l1HO7o8Ruxin7I97gwC8fhyV9i9alUH7+awiNx2X
VV4yLF5qyUhqAQb+PnKySIBy+YUvWi4dicz9aWIpg0Pri3V4TQrhL4H4+9+QVaOeftgydnYzrHo8
And9vXWcqw4VrQo7dUy5n4XUO4XJFvwEagh4kbN6gAxz0OTvuVBZU822Ec3hlIWx9mQxDCvPHd6z
lXiXfVVG1e+XfO8EGnUn06b1n3sUWkt7Zh2sRtMitCElTWYOsmhnDcBrtda7STRPlLmTEeP7DGX0
fZj97HoztJaLC3aJOS011FWAzey6KZXtcgqfM5JWCrGwC/eXlRF9XrwfxKDa772FBloNcen9MpgT
PjisupFIdzV+aEv32IH/52bPKhy+JML3Y2KsxUZ4El5syeFpe0r11qyj1pYCZmZLp2FrYfVM9lAU
9k7F7557sp6kUdr1H/OAAktFD+FQZaPLuO3fAO6SfICG0ymrprCkB7WV7SH7LNQ0fKhQcE5WV2EN
6oQ97fjiRSHIAqODp7+wk0OcDuYP2eWkaFI83cLA/AX/81bWR6BdjBMOOL5rhqbvD1eNU3Op/7Ed
BbPB53maNcVyfT/h5MlpttAEn+aFr5M20QMq5iBFH5prY4vygE/l4CSp2YHd5DoR8WPbQU/hRusg
oE4BFP043HXNWNvufvBGoInmVGxyet31tYbUQPwD0rTK/IhnFczneApn3+FzoIflQi3w80pDEH79
+3YyCY4NpecYg8oC979b2XIN+Wy5yWH+mkNbkeJyQjLYOQzEBFu1xF2dJr7et5qbuoGhI74VkG7C
7nMGXyj4LPGJPU8PT5XJEfJrAUqns2cJS8Rs3p5USwocPLNshfpDMK19l8arbwAlwX6c+yhPVurp
YlAMMwcRTewqym67ndl70TNRVYnpAvriLLwWJbFt1nGm6r0/lXmGCxxSvbc2KPhF9QBM9lxa0YQQ
GyI+ObY9CzEdBXJln8LIJoEgF8g+toq+RWhu5htvQZvqHOtDckIds/k0tpHGsIjZZe2SjszoY09p
KQANz5MZxUpirOBNlNMEPeKq9JVkUo9b95iwWOOxFF5F0DjuFLTlre6XoBMvVWKswv/CnIUHRfPG
rooWlLDK78ZgZlFhNGCjJMtOnkd4N4vP9vcHTNS7DXVAAaf9ZQY6iq9GwON5Amd2VVSxRrvqqwWU
pqExpO0OtqKh5vauP1MD5QU1LP9mk9sjIbrifWuqo9q6NJoKpYP0cResz8mnOAQCctTDqUtL20za
5l1xSAwegExqBhgMj7CBzLiX2GZP0juodQmbzJ3XKXns/sG8rKDx6vw4I+8y/+Cbwa0QNveICvPP
8QXFY/mMZnvA98tPM1S3kK5JkL+Y/pdsyM39a9uVTnDNW96B06zn/IH4R7qPp6L9hK2ZrjT4OWDE
JXtJXulZPQS+zr1O9IXCJq2KQJdyYVWFcr55wBaR1ZH07IEZLAfh9xRukpGOx24D8SmWgMEL+gfA
41Ua8lEystn+iaS2EEjU3iR5MCY2jEXwSrPwlJ/bYGIDb8tfapR1Kpx4MLVuJ/854+Qn9Pbc+Pkd
weBEyaO6hws8hoXunb6N/9pBi9XxqKejj/Oz0/m9fSh+shCV1+2mg9KkZTXADBE4lDKcfaQeowMs
Oq9ALpSHXr539evy7aUkHPnac2YHgHLw+mBOYf4cqyMOZLUTHHyNJ4KJPn6PHWOmT4rEG6RjNn55
ThDHw3D73NoKkmLbBJSC83ndWmgGnnE+YIRMDn44cXt0FU6kXoQ5DuXaqx3GbLzdeSBZ/gOR9pU8
x9JAy6tF+nFztVtQ2FmGjnjeI8NtpB2MbSHo9tshlJg6FbhVqELzWlUdaWUdifbftMKG6qBH822b
tEPBAG6NhlI3R55ko2TT4pLia6d1ZcgynlWUQbqk5G34UYO89CrhlqYHRNgU8eEx26wyYem8OTT5
sBcWZgLqsY9/f+AZSzdYkyvBIQgWXfTkK4zHEQY4QRedgAA/HNxUGcDhVAHYwMqgnbdcNo5RPfv2
XBMonzhkoBUEtF1BN5jKNUOnjODAhDOqmvkgWqu5abl6wyLhITFyuiJPVpSZ20HOhY1NkYPu1zkR
3UUQdIuFCdWNasQZCD6ETkU2Q8pzNpnHIHkd4p6trxc4Ji+Fe3ta8jJGeBTsvyIEvPsi4asAAkv+
wtMGbRBe7aIpUzxZLbrLok/0y3Y4x4AEwEPNzbktsh1fMR33455jvD0R3EnIsbGKsnp3+FxRsFa9
7JJk6sEbv6G5QsTmsn/tAd4t/qU9o27XQdNbkc9G3cUpkKlhd/22FXTEfycDcBI325ZfZs3qUPTx
JrG8yKxoPQRi5mNkM2FKOiM5BhrpJF5Yx2GRv+ZAYO+Hg2Whxmed3PmxBJkSOtOmvrW86HwocHmO
8ZV2QNmkJ33EjGd+LVJYvS7XierfiHDGOqohZOzPsGWcKKueCttYvgwPeCirSvRBpa3KsJOemiTB
AXKi2/oroqFIWIKTSSuDN5y+bf4Sh38ee4YCOzVflPc7YIMA6CWd6tXKhEVtDJfj1i1eThOkkGru
PPc1zNcZljZ3+xz8W1lUlzBdDQBcCWehRkkkXSK79ZxYE0f+xMcyXeGMYfwcviTiJaJttc38xcQJ
E8HXDbKxsG1rsnzvGFUK0StqYNBrtQsA/lGSPoFuTOClbs226uihQIsWDrSzIVSXkacipwWocsZ3
6vWJHSvyjPlPgxSw9JBvgO/BQI4BfZFMeSwUaAr3gTDrI//o4cOl47x7dfN6CMFjpHdZ1U+DBhkL
q16X4mdUy8v9RgikpPMi7QWGtdGIwgyP/7V7vVHEe2qYFGWVL/yI3yxa/8ig6QcgwreZeQEaLb3Q
lUhvfA5gZHTye+CN/mQL0xza7hqNKWhWc/mXoc6qgRseYw/K/AU/2K9hFW0HUnKO9jxQ0Sa11ViY
IuSae0oL3d3DHt1DxzA6LzZvdcfaT/VPYuylxMo4kxcRixjDhXOFjRC8s7/p2QTG5hBAdtQyPIpE
h+1FLB0w/+ydiHbqRDMUkB1+mNaN+iNPc3l7nbkj2OigEltVl62fQjxHwsZqD745HejSMTP8U33q
3r/qcvTx7qspK7F1/KfoELTqWHwpae33m21v+pLopW2Dh5YvNuMWv3bPrdooZA01AgIopCrDFrRq
XrKfbNHGeJzM0tzDUUKwADuAuaCZ0zKLiKinquaGlnyqVxKbY8mEgxJIjSnV5xGsrr5Yfe/CCNLW
r5JHkHDq9WX/kMQc4vB1RvIq1DbITadTzgnmSaSyvkZwfpv+PgEYUu2Ry9e/lBydDIIyK61S4HpC
i3sahGmgQLHpX8G+7lC3ip0nJ9wLUGGSL1sEoIzysdG/BEc10Lk8XK1VcgNMuUlDCdOL4P7VjNhr
Eb2YcSJtlFrmDleOE2ZEfjsJL4Huaoobccw8ZwpVZneAaHoqUGYBoXxSV4/J6kKb5xd75XGRNQFK
zdsta1WWgLrhNZddiHfbS7lH6YaSnNIGsMrUrwr1AfH9kujMh8z0FH1zvOn3/P1edrlu3JS0JP3f
gKUwzPh4aKF/uUQb5MUvuHJl+8YlsKXuzTl52YF8Y/WdK1N4W9ItiOM37pot2pKk1eFDsg1bqXk7
JRSegqaqzTpzugOKdZpfHWp5jPnXlDQBI0mB1707mpbFhuBsmXsSDmjF4KNulhZZsFqrO8IZ5wTa
FAovr9j5vO7yB9v1lGPouQRet4zGx6BOYmSkUzun2Qcg0JeEUZ1U97nHwmT1gOXoEpPDah8gu3ee
efH+c+R5ChYszqEme0HuHYN4Rf2ajvMaQZV/kntjf9TVKcFwu010vKUkCySXGXS5O0yNsqEZdvO/
Sj1IngNhkfnSXBUQgbwhNnWd01RSZAMpk2wbGetCyjWXH9DwwvOZ4r8AStDPNgln0TfnIJu1pFs8
dCQg8oM9djhP1BrP3ue/GPfNdrsOLfpjz6/947p6l4VLMFUZQwcTA2dnb6YDQm4J48SRoRhWelc6
QSSss8xcO1APTpkljLLiwooLEDV01OdoTt6WEtYa1PyMWI1Fmv+dQaq3b8/1BXO9at0CnOA5qTiJ
vQYuaFDycjNjJYPwpxDbJkOktTPE4MLU2q3R5ywYNXITnDPde8FVzNheQ8h//2GL7eihR9VvyJ1Q
u4S90WEwVA4HfjpTSsB92ekv2ZudxMb+srWaePD74xyWrmfROYPh7TWvtWtPGhXjgu2PPPfKxoDn
ZjdC1PkAcrhy92NcqZoNdnYqex8JH+Y3NTr2Sr1d9bWKj+LxeL4uojxYqRaeQqKaD3l4wR5L76yh
ob4675FTXCi1upQ2alww24Geqsnwsb4LuW9jX4WLWispF4IWr+SWFtlPzZK4lGuzNZfS4JJFZwup
BRaRNzAkAgOu2fL3V/PGJ9M7L8zeHPf+ED+54xgE0FTrp8z059JLkQUEf/cw+Jh1INxj+rqEaZ8a
w3hb23uBRaU3tzha4QRXHXjB/LA+QnPmbn6jmJP3GMnitwvfb6vyyF7jwHE3ulbxyVZycjo4qyNn
b5cYqoRHbp5IFB3w7O+ghkjtmvpYwM0gKWICGPGj+8hE+FzjD+m8F5AFotn/y0TC1CDKGZutfhfk
DppuEL4+PbmT5QEAb7DeCKs2Kb8ytz/+eS94a20gVbA8zjTmNzq3ed1Y0oDof9eA3/FlSm8Tjvrs
s2iT7VlJ+eWZIpbDfZa3tkI+gkzHQ5oDmSr/KMA1rlk85nNJ+5KlMagMJnoqOo6Odoajv1BTzyDi
6X6jlvd7zu9Iun/SYtOeTXK1ViR1oFc5sxmLHCJezMKoaxY6vKTKXT3Q01dhbzfeGZLkoAPoiCR5
0vBLDQfAPxaFq1vT3A0K62DfVMRtzeE5MjwTVeNBa/cvwYns47BeI5r+Tl2LS9BmTC/5NkMSetJx
XXs8zosYODD9d9HAOSj0QmtyNmeXw3ya7Df1ZtRTgWeNqcHdAXEQNSmB831Fb23fIhkikUd8qhTe
HeRBRd6cvW56c0So90ociVrEhqlm3lsIk3nItXm9tmT1pnNPDRJaqPatpCOBqt7OSm4IKozIRUuo
ZfEmH09FSVpNpt3ntcqavr+d34sDXwAGpqRoHAes82bNZUMY14LTJwaGS3+kU8vrkJFKkwnyNwjZ
rElPicp/SFBRcY0XJEk4ClyjuHjJyHcIXvaWSmD1EokQe3AndGgEp+IFD+AQtAXUgbc8ix4I3VDs
5ycxjgLwPOv+D+ULiAbqrjWAIaRNyDwIZif+FexnjyX4EbmqNUOSuY0egtxXAS55I6VwAYOUewVm
DO3sb2AfCyu1d+JIJ/stEnQb/uH8lU1RXfIMQGs8Z7L8UTUS0XJ8oihBgGKKbE4pr4uEZ1m0U+qF
k/gqMQekl9dAyMz8A/KwNw6xg7D7IhaVw/lMjMicGFq1JKoCjnPf2XBuknlTelrmaq3lSm2GW6eD
hUGX56CtB9uVRQkWon63YnW+vuTC+akiA6NOqhGd7U99I3ybkBpLqZMwxMZ0g4s1WClLJiuuSE2R
jS1Kjd2pmmLz/36JmRTFZ/NzKqVA2UXz0Ju22TrrZDslV0i02yNBpdPfRYkpCF4vDhG4op+yc27k
Rmjr6H+FO68WX0p5+XKR4XZx1YF8eFE/h75n7BoGc6qnX10+JGt+EmQF29d4f4s8qsV/X1P7vAZx
Ysj+NuD/0RUGiApjRxm4Rv4S1h1q8grAf8hn9WVof9xwmCD+7lNhNz1PQKpHFwK9AO3iD9+vWxKU
coWTW3AwagaQGlgZ9oaO62x+yKKhzddgFrqznLcJ5GBy9+LXAip+dCYB9bQ92RNjLiJn3jwxSdRW
1N6jjFqdWLUWvb20ayS0mPmuq24ESdSsVsyMD5t0E3SQfe3u16D+nbCo4R1IpzHO/sW50lc1n1nJ
6R5sxBK5vdpd+PVJKdAGQFu7dGFXqqAij0RC2TTHRpxh/5WkgAwcKVDJEdF2mgQT+K2nABPkTzM3
Dodu/xdiTgYdTRZf2wJmX+nCw2Z40gCWn9XvQsL2oHDdwa8UMMSNGBGYNgBcdf23LSsUrh8LjV3J
L8jCVcU3qF4LfNig33UCpIRIjlg2xWazryYwdjjpGWrAu5yq548dPxtrcWV9VCjw5qlv9RAsXn+Y
MZLvtqmJ1pZSZ7rxRdFADUf4vWpg3zppJSf+N3udmA7IoyHR9VM1OIlsuS9w4AMj+jBnnAMJF3i8
t3gs7CyLYmKkEb7ObYU9BjtTIkUxo2ymnXVHLOs6/rRRRCM7P2WpQGpnqxcxdOSxB2OauNJaZkVt
Kq6sdwfHwWGRMR8k7QnaOGcJyO091KVaz5MIpYJNNSy0KhUymMqGSgOISiaoXy48bqmvRMYIOnWU
N/fxv8pEveLZm65EAuGONVXQmiX5aoxSZanTyuva4GuwBaCNyvnyNPrPevK8TcYpIZUA9QG0iCJn
5zK6nxsi/v9e5l82+z674f2XB5q77kg03tuxQkzvGpEHkDnpwU8MPw59RUZ6jqnjU7wH+x1/1dmC
oTNbwueygPQlWgdCeGkVtNCsuMoFr6grdkJFhrmvo5gsc9OKMgcuduXjdRsGkS12/Py5V0siWyGX
hQaGDDwE0jO8UcObP7nD6Vq6yYXD6R2Fb5f5TnThJG9pT9JhHfZ+2wzz5pcQR0N1Jufxyyn3K2HW
uMx4x6IM1FSx5a6IHUhD7frXtrS7K7o6qffxag3wTP4clRq0uBQdkN0BtGXz9O6bfZ3zTEgdMwqQ
FuAZz71Iqb8YKOGcZ++TL0ff0jpYxTZLD9glDPcPe2KdtLgwsrcEtMSReAdxbAIePUEnMyJURKrt
BufIZMhBElWeLYfQsOpkdQuCdbJJmWYLhE+FVeYhBI2go1lQ/sFx+OkO6Zkn5X5TemvUC9+Zlt4b
YPdikk+7TmhFHr8HyV9X3c8t7vPnBH1EHu+IawnTUWP4azR34r3DVUazlE1doW2Jz56T+yd4vLdn
qXvrmB0b5Pa9UfQgq11lZQZcLtB1/qRzW5cGnIErGmQs9uY5Sc/Ck+L8KfYUppHvkyRQY6gvAt1b
xSYgMEXQzBoWpM7nF9kGLJZ+Ia/BT6Em6dIWYmjXnmE6a0eCurqCW24woSOjMagSFaGTtaZtp8vP
2OECn5COurmlloW8WvZ2gZUu2jPMkB6z0tG1XtJ3ZmPmoifAdagZiPLu0gta7h2GZmIMjVK37g4p
EY/qGXuATlxAJhngm4sbWamrG/AD3tw6kZk865jwZqsmNZOZ4UTrNSIGxNYgGmXCSIOC4wgtvIsG
uDkty0KeOvBF9AFTmx94TroV0ROFAN5lzX7b/ajpDIdHjk8Z6gV78xcKUOvXmiDJxt+XCdYuoTbP
Wsm1tj2/LdM3jxoP+ZMiCyOFTje/DlRw5bWE+u6+CxTTnEQRr02ueq8mSckjpgHvr+BqGhnlV2aN
hWdEzeulhIoR+aB0UiBWUHFDbXbPsI1pQortqE7OTM2aPQdPr+lzugKp85Ixjrv7aqcPWJzh2HOs
kQ6PmTaGJngR45PKoaMsF2X7Rr7AVrenWP0ks6/cVpLYUy/AoTQQ15jPhTXYDe/IsCbaK6R+npL4
ksSRl3EItUwRENJTogxv7c1y65dKZxMGSi/IzhNZYw6wBrFnm899AQGsurN3cUy3frsKzkC1JcM/
lAR9PW+yWEl9YbCgluQEd0+MVATZR5e48QFm+ZREIzhWV9HJERgbGVX4s+8lueK+tmMCtFh3a8Nr
unTO1uG2H7j1/bHKfvyStvfRMirJd1hoTA3Z+UY9u4SieDxQWUo8p6EeiSCVTfhAn3OPNbtijBMs
eanc7xcWinhPsybbexJl/OxhSvqaB9woF5hE/rbZpqeZc4KD7XmeaCbZtqR6xLwP5vKEkSLFIEMX
3OPcbK1KdoVRd4Hr9iHsNqHrM0B4RVQptQ+/ncTRzFM4WYlxdX3wtI1bED3ZtzuG5mvYgVgizvlH
1YK0+xTCFmA0SkuQAGndLV8MA/qUh14qXGsyd8BvKRk2N2hkNoJdqQrlnEQjJ/S87YLt11mT2myy
PcdSf69YZwSbDQwMTjrpWKdVcRkp5Srtkwd8fjICJRXvTa0aFa2Ji0NJA2Blqas3lXjM8PKmOZAO
RMZbYm1bzbSRuhu6/xWcA5eV/lcqB5fMPVtC45zrXVSMVXI7IfvZPjLE+lOPGvetZ+Jj446DRYv1
YhNvhmwUMnaOC7Rc8rBlt9fNCAlY78RcbgxeRpWVzQvcQztfrisvbpS74WlIjzUFcH4Y87Z4F9Hx
mHAWYkhKwjVVA6M6IeshNWJwtZcAL/dZnr9lYx6KrZAQiNxvbmh2a/34HslJrA098NE+yr+pPrve
I5hcHbZQQgBlqMtn8XemvtDgIzPyxLFbnAtQD4q+37oWmuR3VEMKYhU5tju0p+FA2jSDn4Jw/Agw
ZPWPkzLL3CBAyyx/N8x9JGofcCVMyjD1bZZFtcgoT5lizHBGlVB0LdQ7NRTb7ULm0R4hJTPBTKWd
QLuE7WQMzaIOKuKgRYiRSf3jjq1bRkcCUdl6pfbVFXOoSnATzDjtftAXKxJGaoCeuBCTzqJoj2wA
tnaYznL5cKjTzQzbKN7/rDnh5Wdjztw2/BFMFK2rCokfYdnaeXSdGdv6cz3QKxhRweQ+R9vXp+nk
4zmtj1z91eDCEJX6umG3FFadwRzakGnzgI+35Mv7Mshq2Jqzihj06showblbcZ+oHTsWbuRfmkbo
p1TZ8efI+I6bRJSCrvAVD/0s0KNz96IF72cz73wGLQcl3sCwpc3mDxmggV3zrPcnFhdlPhbbEpFi
mh9TsXzRkTHYsjFWf03sxZOHOpVofAbMhOZl6bX5r2KIFA+e+zep7OrmKqZlyc3T0ZjNiti+1OF4
ElBYgx9gC/ZfSd34N05KyvK+rzVFigWzE3u1+L6dDnvB29qkCfOPdUbKoRYj6uOjbnHwQ46pFBYk
llpv3vTkF9HzsWoXq556Fwc1C6/K/tmC9kxNY67TcYvtmsuNzSC2YeJyetaLZySKOYNM6fhx+Lv1
EP8g3QAUwmYOvQ+F67NgQvTMeZC/7ewXGXUGl9NOakTtbGkdJ3HiOLaTD34CjNfbezUMfPLcmCgE
h9NpxiIowNguHuosm7X04IE8NBmC2M8AK1cKyGlG/wbhSm4q2e/yj4ds//HYvbgwV7e4Kh9dQ0BH
3ILtL+pfqxXomaqY4jqiY+dOqOp6C1TURRrGgE7l0/ylYjWbPhWxDM//lij7H+8uUA7xvFejWyAv
N1UUbAwBf+AD8hBU8qbD+TjAmRRc2Vn1+GvWZcScv2zn9YTUJWHxfFb4vJQdVRO3knUl9eztZEX3
6yNSWM8OSHOGPyzEzpY1iGOXoyuOLwdBJTvC+4hf7kkd+geuS9ggBTld2n7ZeJML/pxqYoTeNJ93
1hl6VUsV5W+Jd7NQcX2G7LsEH6wNdkPts/gRfHaaIXV9McL2Qvg1IPU5AySy22FCxjgzAlN6ANMq
QQWBPdT/mD+3jDD0sGv6TLeNGb1HWJUX5NaUJBL2uBeEII7N9hDQdWGU4D3hW6xCVSJERyimvNYG
HxzZuxHwQVqioYvEZ5M2vNOzTnGtOmKatCeuT3sSEjxidqYXsl4csjQqz9l1e+bLNDvguOE8IyyP
hVhUU7eJxPgjl+SDRDz0cXiYHq1ZpE4lY6QL1dq4ndlHhEmTRSGGYMdfkMPP3O6AuVihyzapNxJw
AliQ1Ndway89SHku64oY6e+hT7HYOVHVysekDKJogGil6DD+ZyiDl1jvYXIQZUubATFTld42CkRt
qUE4LFzg0ZAiAXnnZ9s6AgomwVQBv6Es97NVv+ONWvS+mM/59q0tYZX3AFPv4EgTFRKjWUvUOzHY
mIrMWQdr99xAHqJhUOeRay0Iz2gWq5MyDQJYUCmfTp2hqJ3ZoSRT/y7XEGivbdScJNIFPARoU/4w
sXGeuKYj8fN4qM4Tyh7C0eqqw7ZpMU7tUVgTDLDnIFWGdx8c3MHpCaLqEOnrqI4cwnDvAn5EmxEX
3pKo9f7pfbrqJ8sghvL9uRLKk169OvX3zrPT7Pr6SHnPhVeXVLzmWGOzJJZABNpdnkE2Z2fyV7yg
NlGrY/45mT+q4f/mg+fOTDhRZFau8qywh3E2KlYO1o6j71RUYeihZuDNIkbcEnjoL4bRSzojd3bb
sU5ksWIm5eyusMzvizvLav7OPvdSWtTKylAgxaYN/oc0O5ywyc81pOEJX9U3y7OckiiYUlehUW21
KM8Z0CI3/FEVNK6HzOOFAEEZT5i9QVIPctRlVmDzn51K4fOl2M8U/UsBQO5dSVgxXATVDKlQz7Fh
kWBfeeJui7wzxC0yAEWYYgS5BshxoDhq06La8rz/pIVGQdDuyKceI1HtNrIvQu0jP2yfhredTH6Y
rIMmJIdQLziCD4ZuSZAzyB0/4tRgHqDvQXR2RYZFkBU17uRbhnS7AT8aUbweZRc5PDNPbo7d28My
x27jCoWn6siuvB8vetOdTcRvNQCUdePUPVbbkgvfQ6XtxIlBi6m8a0QAMtf4P0PMBWqRFBCfsXFG
C+ldDx2LJnScFXEls3/OFS7CmKtLtxPKjBr7kl8qtz12NqAyxq/D6gGgXaQk4viNqLYEmX+zl44p
5ZqxPmq0GdvSqUmc10qYfPbbHlZYdLZK05YIBxr5AuotTEttXF9DzHCNnPuMG7GXwlLWveS5wF2N
jHT4W/XSHNApCXtb8RlaVfimpFsjdU9z2z0wQNZhq4PyFOq1KGPxPM3qAS17rTcLQbzY8bM/IWwP
69STL7A+xgxeKw+yLSuNOvcl8qqulxPFFB64HW71uM8Gg19/wSbyQiBXkfQ+9W2ksMiyUfQYbvH/
2sT9swBxfHYykvnF4YmPdYo+5k2jppwAEqcoG3csFJl41AE0VyigPk9o9xUuR6ZYrY6B1jDWffQV
sM4lE/2bU8fuZBBbCtFCMRkUdHPE2tJrV+99YVhQX5HuS0IClci0J8tyXrSQ58LRbb4UMqF0X8dP
ZWzCvwjeiVvlAYJac92ZrSuK+IHdsOz+NjrtV1BEndlXbYwbexVHUTSmGl5HZRUVbDACO1ZIvMJu
5uWZ8Igu/hLfoUmbrqgfwwTazrkWBbIUoOxzszjiWLZwEVp7bOEgUrTF7KjoBbiE+OURzDsvHSxp
aXBZfZ4kf5dt6yVnAEN8mz7cHNme6/lWfBRysNNw13ly4YUxjLfN82Zq1nTf3YaQxbSzLS5dnKaj
VCtT6Z65WNzsnY/xj6lb5p6MgNDptK4OCi5WWlJd0xPcijS4arT2T5Xtdyv4Y/jkY4P9yOrbNZqM
3fKPZdNCq8Pj9PL6jJZcOP1GXy90QLIi9PvvzZZ4K4gOXKJtn5Qv0Vd2ocq11P9QRylen5KOQvdX
IZlSxwYfabuB7VcxX0IeX2yIKbNq7JisyK9MXkwFeAUIh6JRCDTrBPVpHYZDazt1OfIPY4cwU0fb
wq16o8GHYUJs1KeRPlyVJsbnbbLwsaQDMIhjqbwmqGMKNELCEYhLLNDxUkcoa9aVzJ0WdFb8HMvp
a3LIS7cxMBbT74JwZqwWDtHBf7ItLmnA+25zwqqk8vzyWba3LyoC23vnmFda1Xl3Cc4fTTM4wjR7
eaQUCMwdYe4hSvIduWlkaqqmf4uHerowbsd2SV1Lm5K5I//gwU6h67Lc48gNXIs4J5FoxLbR7G84
86YObAh5txR/lceOOC30k1nk6nSbNSmXy7+r7F4EaeIlZcfE6F+XO22O79PJNVmTYVhB6B5MUspB
u/XF82r02oZeFyUHa0gLxDeW/08dG//KjKmIyZOYsToRIsyE6HKJlB7miuV00cM4XSmxt3t6UKK7
ahttxu6j+EnVQLRbjL5SYf2SQ9yO2WSuYF9Grs0IZSPiNNk1lAsC8/cO1FhRLFHzfjtbi9WV1f04
QaTf0vXS/E/IT5cnYO+KkurI/aVYVD9GFL+eQups43Cyr1NOKVjnBxuLF31ePOoCGmIPN3ROPn9g
CIJC74eyUYRM3ocHHJoaQZOOsoBz2vxlvCirIVVdTiLCAAQuARxy203KLETlkWL9vnvHGsx19HVA
ADkU9zO57fwlz9Qp1bbAKsdvON4OK4p8MjNOcYzR3EACZjA5WV438Fz+E1vIKkJ5uuo4DeXgBkTn
ZBeSPVm9Fgg7BEKILWubB41rOG1DUtA8QuKDhekREAWjGyXqaeUBpWcRgMmEx4OcMfeuH+d04k7X
uVd4TGC5Tt9W2hMsj7MVatWdF9iOiO+ERksVrtLrUpFJKalEZLe7+yJRozblKEkhRzSMXCtSf7Wv
ud1oyDGyZkuTZ/1RDOzNxMr+CBk7wC1wcC0Iod6Ndwozv7qkZ2aeCGWiQCMgRo7GNLltgDdk0tOS
0ZtG+lkxDlVlMI6NXy6+QHLjoHHXd8ypHA2Smbl+tSbvPkfdO4UoAsWFEq0VTyRfDHYSP+HpPjSX
TzI4Zz5dBjr17YdRQlUqOsP0/ze+HgvOYWFInxSjxCnQGryJM5aJFWSXgFnkwrQD3o8TcJ+5U0GV
wOL/ada3wS1z7TM4wDeeiezlPbUBvHkziVwf6Hl/tcYzfgVVptXnXihdAA++awAkhYrmdfZnMmmO
YfzRuBkztzjvMC4o19TXKQiqX0B1fMcJkQTdq89EhHF8oxCXLGCQX2BlyrDO/3y6E1edn0JIEthW
NgmhchNPtEN2gcPvJ0PaQr1ULxb3gbin4ssuQ/GhxdMsDq359B4PaomYdpF/Dpo7WvZ/527DEv52
eKRWy5MwIpfO1FRPg1SgTLZW4DNr+F11hpJDp+K0fio83po1yWNbZb/03p4fpKKOMk9rSBUjcZJl
132CKJOjJx1kfSQvRAqPa4SuXedwWeQf8UTWgRD14So1XgYQcLiTyVAVuTos1UJN1sZ4nh1J78hd
aAOkTuNbiR3GrgyvJlVAN20qAwVUsogGpaLkCHzjGXJN65/hLGnM3o79RBCbYqq/lh7JPJ5Pxl65
ZiTculGojnmy/0/Ng8vaNjYDwdzkynqhiAYUZ8rBA3+97bvSduMpTIZI5NUJye6rAI/YtzVVXrG5
7viVpvJvsau/F8Bj71dextX9wfZgmp7RMzl2X2SK6p5+aQEZv30YOfpyPkGn2pwck+V+IIFo4XSQ
YFtU2FYrNS4N0SC8LoNtCZyZmEysCvhMBxWwNPUQoMvnIjLZUqWvhuj9sn8/HBfizyipU9y5dOem
Ph/UJsHAXeCOTIYI1jT/DVLHEGtwAZ4/XBaBoqX2mzye+PZzdmr0CyrzkbzynkK/NRP8DMwHQYEe
mDuIGQIuKVLwoVK5Yy+ld0nv++YiAGZVRiVwemOoacsso0XkgUJlP4e/6oh5ZmDdK1+a8ySh5xcs
G0JuZxxpw9vzi0UKr3LNhjcYeFlpq0crylpR4u4r9kPSEpli8sp9SObPD8gu4b8s4ZP1Y3mdsvN1
e9lQjxmCldyAzpBx0QWvjvarCHl3srpKTemepVSmK0l82Wj1hT5GQ5yr8DhBEWpvQuF7VUl9attp
iuRjKdtewglkwDNoc3iTjiyJJSQPNLnuelEoKGTZEC1zrgVaLTLtOodSqA3gZIq+SpC5dzTXv0Lt
Wx+5dwJuZ05wffK0OMfXzkm0RrrUMxnCqkomR4wzwMTs+YzmnXhfZNTXXLdR6Faw6nY+rmqUREoI
0VcpS3pA8Quf1b8IHuNujXLRYF7NcEEmY3unMf1IAFvwCJ3wf8qz0dLhpQSdKu3mUmrfBJTwigAG
hkCk3VFxQ5r/xS6iHFrJCujvA/H0/hjVrwXJSwSSJUuOFZzebyQVI/rCK4A2e4GRNa5S7i8X/tVc
MRq0Auedr6da/X/rb3VaxanAnl2dZc1Pdlk47bajWPiHYlJ9SWUJwiC1a4402C+j+Uv1YbA8UnLQ
Aj2Ui6Fhn2pe6M+RPNVueBy2uCWuOoyubu7yPC5p2z1nof+pyb5vp7lGSiaHfS63SHezs5i0cOKZ
hH+egb6rcCnqdwSPJXpNeTbQG3HkQcJ9j/4LDyxb89A5a0HuXK2yq3zYsBIPqW7/BCOkU+gM/i1E
bH0Qmd4zSUBnFVOb1YvUI/YLdcUMFHiaXEnJZraw5fNYo6tFXa575T2iiW/ZaICLIkOO9kUNkTj1
xk5SMKdWLee/vTGFoPU+fvDbYYqGVGAEcXLnYsS12/YTbyeG3E49aR9tutPvxU/j2GoZm9kEYgsP
M+vRnqYtJtQRPhGSoevaVKZzQcK1auldPi00WQELMWCwSC/p+Sx51BzGy4KgcxE4cd0gXzUGbZif
YJ+NiHgLU//ljWxbn0dHGMDzlaKXqCMomlsrYhQ/H0EH/BahEnR0K5B6OPyaLqsFk7sdOco9jmaV
RCVRjUJmlYOJHmvRQLTk/OfBBdywmqRjWI4v9L+3Jh3y602vk0t/uh4lj3YS/RY/+mzIxWUCqylz
BgLsrUrfeHFcs7AjHyn7/yK3o7SLUTIMIJOf6zZVDy9/IzP8ToALGlAsm4jkpeN0qncEhaJ024SD
ixOWIv2QnxP1R4zPGmQ5HUrrV2dkSaKRzC4dT0caaQFeHaFyjCyXDYtzCnah0Zz2rk+utOIuVWOe
PfeytGaYTnThSDLi9/cvnGUjLldyCQAdDAP9BSN/rbJyOaYqhh3NNTpTKT21mR6P3QH0tYB/N7t5
PnwaWLDxCuUJPv/lMQJD7QMk9Ly1xF+FWXXAww/3EViSPh7T6vluTnFEoDleEubMMGRgyIyem1KD
FgIm46AQpFI1btktyqmTTFQ4Guz/12txfYGbGEwghn7qm2JMMl8MjkKeVpn7UgJVkjbbu5e+487o
40GXoJB32QhXGeRA+1GPJvuEopria7goNlsCYp+wNGsRi4i348SG5GEYKVz6zg/J8l4spxl+wvbQ
1rxZBJLMfTlSa/41wKWBuyeh67V0W+LZrG3pjPSREWdA4EAIy78p+NC6I5Wq3OwokvYj1KNKLQos
e2s+JK+gBItS6ocKwQG2Tb0sFZGzJFxBW24pMA8A1dler3kZiDwhYHmls+RAW5yV6LytZ12oiOsV
7D8OHnfGgrThOB2SimZetTFbakbPHWEKpx04k21NF5uu2jYlpn81VIUU31H2vUQr0YdMURNoD8vv
cYc9/F4FeQndR2sq6Cym9wb5qf3dBvyy15nuMv9ntEoQEAnkdz3fw/dOWeNFDztKJj5YjWZZA3f7
SLB/tNVvolYdzccFRktTJF3EESarg+aGHE+ymJnhriAzYIN8b+PmvfzJAHYOZXz2NH+0frMZ7OK1
6YrFdM+nhbwMAqWbbdyrMjga20gURxCYCdAoaxT9yZ6en08rMdxSTp5NftF5X2kClmQbsWWAgWzu
NCqFnaYQkX25JnCytHqnHpQcw66u2pG9MC+80R4fKmyp3WXlyIWOTnTyh+I0Oeu1eVxxWE+jlxpi
ZAigMkn2+A5yua2PYWLCa1Om9grCJdsvjvGia8yDhn6nb+DbgIZDV2MRB8VII7QBlLVp3FQpm/qv
T8qo7i7ZuBklaIsHjnjuZ08yt7CI62CeXpKMtSbHNQ72xMtKNoUbckgsL1MxHKvXRdAPIfxjGXZ8
xmZuZaGf4onEehJmoJK75d+uRjq8DrOvq4q6083Z/ish229g+/tEL5QhkHju7R/jVvJPBPeJkblD
ezIwTwOP0LsXeq5iIWhMm7V0dBVfRtoxxFu2VWFR+iY+4B8MGECVKlA2H1d9Ss2ayYy6I6sQdCEz
yaBCA0t3dZmaIitV9S3cmPy+nfpo/uxyMcV9ImQvBggi7t2nPCMwnPrWMpKSkYMf9YggZ8gaQtqH
dOwAhVJdGiCAmKi3li8kk+vhIT9FLzhSrjdrYRDChpP6wG0VN9hAK1fjw07OUxQZ2tiqnhbEaPN0
2vbcWGet3NlrA3yOz6l8Z+t4/MBoUs8qaiQeaDmDbyTrkT6JXDjffQsNTr0jydRcfUL3iLcebYpa
eQ0gi+/A+DgKJM2Vq7XgfwXOpcgjcK6x7K5dOaJhJT//m60NTEEbaAzcjlXygM1e5lUsgoC9fVoZ
WCnrRd+P4cNMxV//zhHc+/3W9WnTjxau3BvNkwDR37HFTWU2PsSI7G7OsS5+ShHwaqTvAr9jEPNf
UrbPldDpTmGpw1cSJJdG3cZ+ruYot2gfVhu1Wr/nE58nlr8IO2lCObQXwBmJlCqoIe2ulWyPACnA
9hWtXzfeqz8k8JlmYo32sn04jWEBm4AR3kAV+FjJbJpxL2SErVzR2ifj5spqA8u23/GT3lzXgnsH
+5iAz4k8KnlIeGXsze+/7lN2b1RASA7by3oGANwfKWm1KJvAX5SaTvH8HICCjUrd8yQy3nxuYaLi
QnoiERvhBxs7+sr1ZHb8nxvWUfCrcH3ek8t0i5MyV3qwLClt9mKLEP3zPNocyVuuA10hjUSHy4fU
zW3HC6hePBdQQRjbEvrNsau64g0DC3xEQMVvyk5pWbi+UZ+6erUV6QBWyFjjfz5heWWTIA6eSr62
ChpaOU060ujIbYKsI+tt3aPSf4X90gKt+GRezliZBJuIPJCbMWM2kbZo4A4ZOyLI+7sHDEQpjIEv
iQ0ZFrMSP9APK/cweYnCB7Jz2w3/df7QzLPmtndkn955Zl8pL34Sf5Zm3Cg3Yqp3Fh0EhRN4twWP
kqIRl8dcEIsMZzpPYVA7PpQAYRq7H9U6rMoYuKY4WO1TS8sDmY2RBROXpXKY4w/j1i7iZa6iSTQU
rQdc2MEswyle3JN8uppeAERoDtNRiqV7LMRW7j9hurFaCQQAhTy4G23yOaNl383m9OSoICVrXQPX
422GINiPSYOMu1zYKIMh2WlNqPUOlrrE66v4IYMCAHmzxJTgBqTWrdJsWk8lxgbRbduuOohJ8kW5
dn+HIC8H6HaSFM1x7OAIS8I5ILVSnsJy+wmQasWrqYuoW8zSyrCoYCJu9oh5oTQWARGugW3t67ba
EThnbhfeQyxgKxsryPzqDpk5ZZY5sqM4nlPX+Fpwmyk0YUaJ5gY2mnduzSBxqpau/5XTTs+xu1+3
TYxlFv4UIjRc1sisO7hShuuYu4qG7BcNNCjgw6DmDJ4Nmhw9/3JxHj7BPpL183qtx3yQqaLTs2RJ
6HxyyibZ0ZDDVuiVtP16Y6zle41qpG7wy+T5yMYkqc7uugXnZq3awi6pE+mp9wuACQ+bBsCv1dgd
Nd/gOFIcGkGVZAw8SunsrkFzDmNHceVY/M9LhxDJzEN8QH0Jg6pAvgRVC2PPILlj7KE/ruMg1bBj
5Ut5cZNdBel0byPjrJ02doJqm7gj1fw1zleyvRkDuxsfXiSLjIWglinRO8ZWj2dy3VoOOx9PjAwU
zH0c+xQazc1t83SSSyi5zQuW4rFpWfNqj2xSSB0dmtR6JfGapF/26Qz4p/EbUICb+Y1A2bmyu0Va
h3ltmITxT2w5Fi2vCiQBn0s5iaNueCVfOTg+M1ijwOI2D9cDPkG+Uzbi9UTt9zXf9W/yD0TLAU4r
nKHZHyI=
`protect end_protected
