

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
k/BYGcITVzkj19j2HCuCh1wA+/VTFblj2MFzTMZNbTSHTj4w+cHpukw11MhMCn+1VpaV4XPk+KCT
F60iuGPAiw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
E46yTwoXeRY46I4q0sknAG1i6oVD9Fby9HJTDGmhPLYly5mCC8LOLeoAWOb2MChDrPQjbs0lo0pV
f+CFyY+5CIt4nvyaK6ks4bOkktm8k4x8SdlR0YtaVdd64mBwZuzP2CDguB2f6VrE7ugyB9Pv/D+y
PzNO42OY0KKracv7T9s=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
yaX0EGpfIrjKDq88PFxDkQ1Ih5gVPzjdX7cjvCAtwWOJixqSt4eknB4pThz4Sb76SURO4/kG72IJ
X4MEkZS7pR18pfDUs0oncDNZ/lhY8qySVVP5KvSvSGJvuEd4y4JWUPlS4pg+mBSQkD3ynhwRO+7t
/q5f+vhDl8ABSWnlKqs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Lea0NTFYyEg+GckCXsxSFBANfLYogm0qN5YvRb8u3w8ZQu4vVwMbl4/WN0QXKfZy2k3ZxNQKz7Dh
oFdjoeGsDLzMnKSnrBT1pHIi9PGOiLLrg6Lvgcg2TM5HrK3jIayh/Y5AnjoZLBttQ1q5cMiS8QeY
cX1MV+cTx4ovtKU+NIUTJbPutsdS59oWDtjR8DpN2LnfIJ6nXUntisb48CVYqNKGn3QZ5Q9SeW3b
xwlvAgIsUXzx0rXauLfH/BSPN91Ja9JgI+cb4+D8D9y/xpsjpMIE8qGKkKZT9w3gDP0xfprRY/mz
eayiSfKIPy4P1XQfBdDuTHG6udNxb3Gn/xvQ7w==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BRgljJEeP6z6vVvDwBuXh9cKW6awpue+BLUABGrJ/7mchmbRYCpvdol/LFGVHX7yiQwqBDAClMv5
xJ8KbMro6CvlKPYH3A6NBuEbPnBfCSjWwn6p89wdQeA3stqsOw19i2oiIX9DAX1HNpBtiJCNKdOK
0nLwya3/SE2z1/VR2GIcR+tak40u+wRkQbZKx6m0GiWFvcZRKPbiTLTFnTT+MDqgRgoAjaUHaAVw
tP3miNiSXswdta959DVvVuH/uQeXipnpEKpytKyq9/QSzS8wsRDdWG0SzDLLITnXMD7C3/ZfGirJ
+MwqxM9f/pD0A3k7376qqv6kz6YBPfyVcNMy9A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
t96cw5VHs31F0QSbsQRgm/N4gTp03rujgsz0kvvkpIXlRIuQQZQ2TMZI+9F0Kqm9UYCsHzsucT1R
e9dnnzUZ1azv6XAhIozJmAJx9JNqEKctF0ycLby0+bxLRoIts8dWX+wrK8RjAivYtKbYVfImpn6A
04qoiobCCJh9Yq2eE1Mw5yELVbAtnkGGTfEezmcsny4L1DIRf4A1ISPYemouvYdZ0B5OrtXZDX4/
+6fMrKMr0hHxqHGqmi6lHskRbI7/T78PFj6oG5Hoaw1F78As5mttBqvaoC5ux5GCrNuIkguMTWNE
sRdfJrMxL0sNJdDNsC2po3KppjTuemj+5sPkTg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 125824)
`protect data_block
mMTJCVKRxQaQvXdhsM+8mstWEJYMOBMa5RLxfD6UVPp05oNAIQ/F9t6KwgH3qvMp69vx16WIDzwW
0zvsEDzpho5IUbjluJpT5fr+Mx2+3qVKcmuAMx3e3+iYBhmrvoNAXqRg8i2Ugotqmn4lir7J9Iqi
NCheBwIYJ8VecI5jnd7J5+Xvjgyw3r0ZOeRu+EKvuAzWTAUfSgjrPBdbrPvzcPaoFyjvMtV0WPvs
b9G/Zoo2Rrw5DRxFkno/yLdxre8ozPtfdAMNEUR2DhGpCy8MCzkTd7eDEr8kfRl8m13ELZyBOYF/
0UlB8TwWQIi49oy72CDLO1xRJrpM2hpIbgCJzP1knP+GvfZwQV7WWMRPdoAGikxni9i5SfNMs0cj
o4P6K57tKee9fDjYl4NL30R2TotUltdxuQyGxPrseP0/Cbb96k4wFrUMgKUz2wcrEo6UiIpAALvn
vlsXiDhCyqRvbUmzEamTe8/qBCRkHBenLSKzVzf7cg93QCRbBe/0l0X+tJxDLguAkZUJEaK6r6Sq
KxvdkBTRiKspbugjXbT0387KSxcBfU8W7O5j6pEv6fEL0gPCVWgXGll8zEhIKk2bKPnyiefOcmTV
h8cy/7kqaqHHHrqWVSr1nxugOr/MEN1oS3VY5MXA53vCx49CSTRv3m2B3GTAeUHZK0QoCLrFYWQ0
+aiv5YIH6ljRflr0G1u+/EPJbCoWeb/ORvaRIADZ+G/ZibnuqgwmwusGUoqKv4ouQlI3t7xZtXE4
vbwYAJbB41OfG2GIqf7QpVsDIyo04mOKyJ7lxeQgaqipnthcPCJCZ5aUyZfGTgFm6oVo5ht5Ynih
IIFkz4FssGZmKxeEfRpdLdbxOIePK0x10tR60DCqb1hFpM2rFlVzwtO69tg62UT2Osj8apGKAZVR
f+ZWWyGGUVjbMTdPI4hNbQLVpOVqS1Bgz9U/SL3JziMEKTKS6/hZ30RXDSKR/ruL3sOTNxr2VqUT
Z29NzcqnGUlogrcJ6Wxw3XqcIN50uG5cA5vhmFlj4DsMy1EdKYC7TqtWU2DkaQg820cvYLIw4pUl
jrHhXGaK+EYGlDLMLmVAocZ0UG3xeGhdmDeGaeCUXi8gdg4DiXUci3Wfe28nRS33PWuRr6RD/7QT
8OTuRO8Uei+7UY3b2FF1lIHmwQuGjyXeASD8ivH4n4vTsCQiQAiuHLjZjpBXyUSqNE55Sa4ZNT/a
/VfwG8oWDyDKCo/c26pXM5IiMJvImaBTTAAWG8Z4sTzwvOpi7WDHLN2qcyxCRgytJ6I9Wn++++e/
3l3YVX3J1Abkba7c/EAeKvy14rEs9NtLzfA0RzuLDLcqDGLLPFjz/9ySd9J2Og1LF49SGmTFo5I6
iw3+mKaM8Aow2w8BDUR6Yjdo//5za1kKI/XhqDmHNZdIW5eeZowdqCfRADYA32+hMUBKyp9yl0OO
TTbHdGObWWyGv7ud44b1lAWRF79/iudTjnXdbfXKYk/DPoNbYBfH1TmXU9Rt1DWroLNkEKuH0/BE
zg2U9CCsJ1e7ZSEGe8Uu/C6KTjuhYIkYF4StJmvN0SRr5qtfDkgG/x0yFzxMCDy/EcUfUyHgocgZ
N6KAgoNyBbqzUKItNIrIepjVexja5M4zIWZZIiJ+HpXZxl337Z6Lb1idblGktXISwOGb+QUj4DJD
7UQkUD05v2cZQ2/Zc3Waz4hTDOa5Ervo+oxsfqfOhP6mMeYpGIOzLhykVpTcoGq7rHssYjnGWnBr
xFSxt/7UDrctAX/SYsgQ7s7vFBF7+yM0zzfmN+griNV87Ud1ODmVoU81lreJvASG3qOxpH1OIFun
r3CZRwCTA3V6idtdXRu3YmlpLgrVVwcWWaebUpk+Dch3hK4QryN/Sen5NHsptYxkQWy2vOyErl/0
PdSr3E2KcgW9BbjbHHZ1uHou7QVbZawUD7svuPL9nnQP6U2OnAibi06Lcb6xKpaWOYiEvp1ckrpk
Ub0mPsOeoGt9X7qFedH+o9azJ/gdIKoub7cVV0vBiPTw6TqXWR1ezKG4NGALByIDp1NtA7HL+Q7Z
Yk26Y6fhkxdVE9sTm10XYUjqfiKlTCriuhxy5DHGn1qhI2gdxtOFL24ngdOkx1bRkwso9BiUi39G
XIpRqd82HVSXpB238+2HubKhP88ygtRvRubiSpxXw6XM1wh2HdOxz3qbx2hlGFr4ZcygJBZTkk2p
rYuFPaggjrsb1TX1pXmKXKgj4zsgtcbjzZsVuBAqRTBtt5CcAkVuPLpAmgLwM7ucMpzcB2vqzV3D
7yViqy/Is9viX9bYz6cWoKWuOiVtZpoYVYcnaGXC/66DmmCyAX9otaq1BA43LFGMeC93dEIT4ogs
xdh0ENfuEaRNYi+mLTnythq+FKwkVvuB4wg0WwgvNYR4Y/GFeTsPZAAt3iPBZNTNBJgUIKyWNQaz
0ErKHw9RR3naA4d2E3DfsvZVzrSG+h4Og8TOAYx5EQl4IYL/JgDCzeEk3w/YVNdvdMrUWP8mLFyz
AgWG0kxEAu6BACj1zwP7hTKkOguggllkd+8cnXmCmzKNqLJnjvyXGgeWR8oKwcBD3f2CJuvko5Bs
rDuvOjOBb+PqQ/2UpctnDAWRIxAtANBrJpFBvkjO+wfxw2pc94FdY1pLn1WMi4B+cd009sK/Jv5k
iaXaGtgwXkBPnk5Lx640bt8lWhQjMVZmI/xPZLylT9tO22rPxF1uuf3K/c60QCrH8Xh1r8vhFLMp
LKDyEgs68MIew5YCaWLcXMhwSVf2k3nagtLot/zvFdzzv8ujZ6T3KdePDYKdV3ZFoqOTXXZ8rnUY
ZEPc0S1YhGjeEMXdvor9FQ/hkLH5GoNR60pEK1dir/HQS/sWdpxPM4Th5IjyHD9Q7Mi3Boe4I9gQ
1fOcF71g8gowfJ6kq83tDSCdrlebR/rK6tClzF/kjdsj6Ngl8uCxG1LLIp7vT8a6EhyskYvI9kuA
sGi9+SvXv1r0EUkHnPDaNX5aS9JvL/6PIzZSRscLCoUz2v+Il+kHSYWWb7OWttedBdVgo59Db8vR
M//VYAXrYSIi8m+/5Ji+oLHnct5GK7bFVUkImCrqRsHrsJdGqhTXsg3vvOBwjQOIooTtp15Z3ueO
Tm+LnqY2j2SQwpj0ejuR2ItaW+dO2pjH1vZuryF3YSyqXGv6QFjzVCnUGr06L9PHiryHzan+zYVc
jn04KZP5PouuT+dsmrztorZkqKZ2q2bhwlONf4O3oBlmrCa+QYYmqJl1iviYnQXoutKbF3BwgWTF
DZy18qIYxa/AyU1EnyAfzdzvFyS40ML7BmjvPGIoueRjwuBICum55yoi+/ZIL2NvYp5Pf6vjDlGa
cdRlNAVunAFd06kPm27+pHEuheH5ihDvhH7ta75lh4uXjLHTEna9tpV2LqRNO6WOAQytA+2WUZym
ZZG+pZs7kVQTPnjupJogktCXmPBoRTwcg7zRmdU7mQAY8HVvyXQ9grdPBup0rbFi0dwhxPnyi4au
qzC956PRRiXXYSEmQACE1BRFA4noB2gKamGVzPte65hjdbRe7WLffLEHpolbCvNr4YljoTNMdqJO
giIylaMo4dsUy7m4nXaRw1egI3BLCfkC9pi1cAn3LznETJkCcVnowqv9q3LuJgoR/ZIMkf22nW0b
xayb/N8TUHleDzELjJGuYlXvMgvJoc366TWDBJpcVuQYzbUGsvX201Wqv5ffQ2aArWK1Lsaxae8w
3Z1Y1Q/A1kSanHR7B/SDuslgpP1UCbObSl2JGb9AiNaljaXTTFyuNIOrd+VMsmEjxCuH7BMHvzQJ
DLCQSqBxuPD6Uvv4vONB3YWDX1jqnXUyvtOQ8CIwQvL+VlrTVbqenQGFyqhyXftDPKs/abiFs+vH
poPS176dJbYn+Bc+aeYySUAnEA57jlq71zAYPDOzVi41vf5dCddDPja+f+wmJHFDHExQQ7chEdQm
+4nzbiyOGv2IRtgxt+x702VXx3fDHkkPVmgisP25aRUQ3IywdDI6TFU5m17miV9iXDsR0lyOsgcs
VmLdUFVp3/K29KG2z7QpEnDb6unIHq+rQf124rP6vGXaH4bbmCcbEKiLbfwJ7gHmALo2ZhJXwxo9
JM5w+XQomvQRu8a529/oUdQOGEgNDyBJHSBB4cXg2IiIbHqlSeW+WjJNbAsVoyJWoxiPw6iZzYbb
guyjckeF+EBblALEiqcgS9GHgnqmzWisdB8yT0e86NoNYtVW0eUG8EOfIGuYwkQVeIB6WkMKX0HJ
TyPSxq+s8kpDDwKKnA1ATxr0PKBYhBUKbM9vo56KehcKbSRPRTDZsjKVEvtRjGRhKBR7RaV5wbT9
azHpZSxhKsfIis13rcHIF8Iwsd09OlKlHFgXgUhurIjfaCq3RBqc4BoUMdbd4M54Z7QaXRvc6GUM
ihmG4kSOEP9MiXIXiDA4V2jQ4qLehKQw+qbnB2P4PJ3dEBO4Apsltt+QtmCErE8APtOHfPBX/HAq
JeD7FT099Nzt5HfPntiXAZA6JOYeFdCcU3cKDw/lb1bhD0bzc45alnF37x512U5EjhQ4pZNuwx4H
0SVsGvhhlv6VrgCZeZsyRjOG2D5SsKTz7y2gCXKO/OhY/scbsqLDRRY+ll72uxe2xPTElrUdN/o4
nT6I7SoMyUkvjAXAG/rGbvirP67w+n3HNhOiVlEaYqsVAr3stbj6jezY5WG9CQXYyMR1zdM+Fgkv
IhoXJSM8R9TXvLP83p+49qLuMoxUJH8jHn2am7VCuCsVPk6Vv166MS6EXv6z3tNlG0TK/gjYGg7+
jVXpqp8n7PViU2jGeoLrzDk9cbNVKY5hdkyUFF+1wDbirs2A2fA8AkT6jAADTHeQJU9K4Gk3d5j3
exSPwYX189fRHD9d/fzYVFe9dC3TvU/rLmnvv86nY2aJhgDHuT52NXm6n1MzqW9383/AaM8TMwnm
3E2Bs66zAGipaziHmzMr9/a5BFd/L3ZJwciNKzUgPJhh4qyJo29AU9aERcnNNzTs9QdinIRG1oMQ
EXKWKc8QuZQ7uvQy9Oqit74HrGkhMri9Cbb/szN+RdnwmizIm+QvMSeOfxwvfzVxKBk8+usLf3KC
YRQ7Unr845NhY6av9xBATZxGW74+ij0GRIroDjOMgFVh/0hK4Ae9PZE/vOFmSNSq4o9YhHWuo0LW
uqWUIvXtYHM7qFZKorQd6UF96aAucS/PuWuD7WsTWU6g1BduLpGy7jSDpPmeBJchnRuoRzDfIJC0
djExIl3Fzk9jigtICNQj1hZLQaNZlDg9EIdMCZ0QKyOx4ykg/NrBX3efjnwWl2dtBpD04JLCPurO
zsv5S8haJCGnhu0FrcaKdrbH9jj3FTpj4VsvfqeghpkucN3h6HAZJFliPDwsXBX+dEKvS13Xz7z3
H4Tp8cVVyzkYllVJTzyB887GvVl8o24jwzYB4VjqoH/MHgtMD2m9wCGL1AQiZh5Y9dRJmr2Mgw8L
Qhczll5mn08H5YQRnJ4LvmXgRvuRYNem9lqNsidQjR/furHT0rjIVtI1McF0DY7TCpCPF1WwQ7Hc
7TRhD14ib94IljcabmqHrSVwI+LyJGKZivGyTZKXkxvwR4jbAi2IhzXHG7GfxaPV4J0KuInx5ncd
B2pPacU4eqKhbomE/XrjtvPS9JUVIdSWNdc0SW0VkswwJo8BIktSqQitMbYAA/UjlUfb2n1RuULa
TstRhuRPiXzZudZw+OSZfMMrgZUx3SafzwgLzc+d065oT9jHXTMuu2wSn94ZMy99Y9QGmdgikgSo
jydQ9e/xRWl9qQ53dJK+klxXZNajeImFyzu0yuNFVbjHtlB7V5VdjVaXqfsRrJ/X6L48TDuWTLl7
rSuGdMTLLkGm2+qIv25wPf0AKmaiU5gDaeCcq5yP+2bLMhxEbxUE3tct1P7gfyMj+gdA1Rj+pIg2
e7wNu8RfPc0XUpjDcMqnO+G5wx12iDnJ9aAXskXXzGc18VdvFkeiTYrvBx2oWMTMstkbePv15WGg
1Rm+Yhmy0mDz+0YBw27LAPI+/wJ/WMnbZb/bwbHs+A+pXsm0rvdQkELoJYA0jlGUGNFQJa/ko3yy
9PTDdOhaEdYlsTTdSselFB9ldJ8S7rIY9dinYLH5sKGHyXjTis8RazmJ7ITOnbACBS71h5V4z9og
4naEcCOEecjzNFLsxpiZ3qv3T8/SQVkMrqwKKe1ZS6fwfHCzq9+sxxHMCazLrp0sj/ZbmXhoooFt
ghns1yRR2etaHgoBQTAhiT6yOrzw+bhwBfaM04X8hZRKB9IR8z5c7eq+TgOuLyfMooi07pu6VTFc
bffGEFZYaCLhBIRuXw15e7k5bGVtlCuYzEc9qDLJDSRDTVY+SHZPIDikZJBPVds+dJVDHZZ/gqCM
vwOfbj3M3j2+bH0AhI2lXPQ1rJQqv2g+ZTsA/SjLVCfmbxTqz2Q69nE8KWM4t7LUWzDjl9zQALYw
YDT4X/1IM6hOGNSulyoMUOuqENidVScoOGaUN7G4ejKxThjO9WE7YeWsUl/XRDayhxsMBwvragjN
GvgxPfJTrBJXqaVW/rQEeYv7yf1rdV5xBLrEui98Gwyfgbr+s/Wn9rYjSP/YRyvZF/0Vul3g+U8q
jo4TfIn7bgiyHBC0VWPBiqYPjFLnhpKwZO3N3QcOhQkrbxEnBZQAUCo0mSd0g/iOg/ElEdQYfFRz
CWxjxxpUm2tKB5YYTYxNDb+0FvlQS39EoV4xIAL/rMxd0xRoTghYIIvtNke1nn76sKSBLz2AKhD9
+bNLbdLWPgivaPFbHiDdkUfhKFyLHNShD8c+g87si0Xjg9s40uJgpJOxi/ih+bKfOL1TKPaMh/Yd
g1R8mAKhLZohSQ35NxELBtFeWVuDtfoZ7f+LfCjDINRUedrhdr/GGVxm0sjNgNKmstPO/Lvnxev+
ECkyAR0BK0+OWqhKUWZ1Yt32JM+N2l8EtJhuGWbD7wwyQ/43yh27KXaViic0TD1lprlSirps59xj
wsEZKBa98yQyQkrllU+gpsP88F8RtCvkm1ifEx0TdzyrYozZyTibkPIPTMVWFaZu4BjlljUxxCfN
GxXCldDMRxMKd2W1HdK1Hx5VTPzkjAloxoUnSNkvD7D7eyGagvhXrSSx6o7iKRXtFTv5SLfvqlL4
fZQ8yHN8yM4YCZ2wopiRb4lfedvD8G4dW6HMpyTYZlMOIQJstMAmnOgRr8Vrbr8Oe0NHUdF4iOyK
pQodnDsTgwC3RWG8D8+w2FO7MS5wk3Pf9oWKdyBiJQHpn/MTPYPj+DKpxOMQuqE9iV0xl9B9a29N
2TwezguCIuUu/ZrrrFXZorze4ytnSAAXjqt6TmhCrpAAB6MiDqn/KnUK12czdewLQGvJ8s00GFuS
4PNiqeNIFpSUGluaUnX/BSOKPoUh39mgMOjZrg4m4wFoihBl3enwqR040SWXwsPgcL6t9XEP85Uz
ZXiqbYBF1Xicflpn3wgeYUsN84VyyFuLWyK2G2i99zNsTvuWWgghFgyXp3ssG3/l6414mFo4Amv0
YPkPyrRswK7oEDe94JE0QcZkFoo5nyiaoboIY0DyTxamVAb/Rse/66Kc++zRnIB8zZo4VIdPXQB1
LLAoUAKF9Kcp92JAmBgamE5Hd7Z9f61ilGq/VLHQr5NM+bMdaUAxaadhz4AHesSzTCOhIImRb7Rs
/JsITCi3nbE3PboIOjUz5XlZ6eUEevFzAp1ruYwBSBo3K37tdbvje2uaJWKHRak2VchxWf/FzeID
hFS5Y6SyxIvWd4MGff7pcERhpwaamIrm5Dk7YDqWkrSNPPyOoUFwZtBLLZXiaF56pKA1PtlcqUpl
3tPyrgbMAsCeUitypiwgrpnNDyaD/Ig8znzavawhLBW9W0Yn6xyxCNzmtbUbKTMUkTo5Th75QdBz
b49sa26cZR0lMOsqBHKFloBiguIl8RXIEJg0LhLGPb9yKjA2t0bNOceRaypas7pBDWTrko9smUj6
UzS8cIdnYS8WIcawibdyhcB0WrsmcaDhyQmaCsYBYLw5+tfkIbqc9sh6g0Z9YCQIYNxKVoA6CBJH
MT8ez82EdXVThf1gl99ceLKsx1TaBICTeh8zmumuSvJezHJ5Gyh5OP3avu82SpodYwvseYE+2V0Q
ntjAdfjYERP8ZaLm8zy3YROvUZrac3gXf4S3D0zPs2/qPCtnW6/funBIGvC3CCDv6y4dyqLD4RSS
fP76yueeXwi8XT20kS8yURk+6zOhwcTox6kQ7MNVZB972Gh9gumEtYpjoJV+HVk3RrHX3fcjfzrT
6mSJYcaHViJ+y6mcEvBHjBkX48UGRJ2vl0ry70IIZkCDrWeaTZBJ+Nm7mPKZ5RiGzUr6raHQF1nH
MIirZOTHspGHCskwfVoSPuWZ0DzzMZjbBd9bjNcNkkyouTpkuTfC8w1CIhpGyXnyUZ/CYdq+Ip/y
9RFeSMtMI02JMFnzuAtOarVRo6hmqMXQcPqrRmk4B3rou2hoTljNwM0kTeFKBIwZoRLvpAkV6HQz
fAf8X7DueeMaemRLgnL6JB6IJhpuGAnaUahAxyWPxkMOqDyNTKFxwXu2IRpv8xvnoaQ+kIO1JUJH
RGWbcViUvfBn2BxBpgLuRX3e5bwdyzLlrRkZ3/91L3fD3LevMi6uMAv4EAZyJceaSbOCpHSGDl+j
wtHSB7LbdncYB41R5DCVLaKtvjrG9NdktD++BMkl3aDFGOyM5UX2LZgHwFfShox9la6hKXcuHJUP
UM1Q5I0tU6rrhr+2hAlodeKTq8sMrS/n2YsL05xOLiEPg6KblNRrzZ3Ns5DkOviS/iLyp7l9QjbR
qzPtAc3et02kTJ28qoFvt/cgmF1Y6B6DXM2qNEsCIoMJE1xqX+Wy3/kR4zsGGKl/KEHi04L5u9eQ
Xc4Yx/lTRBqN+HpeBn+3AOSM2s8dIdnMVGVs4K1klWQMxB6bfEqwVbyeZ2gG++hqRZX/7PsxlSb7
o7beCD6tOngR7uhE5HJV9vf2uOhUn/jneS68+v3nolXQq0XGPapxE+pW27GmBGmVG0WGO/hSA97M
tNXwyCHBmtMKs5yjuZAvMTF59SLwnTrr15FQdr6vK8t/jWuRhHGi8PuFm3hCgaII/gKEh/tXc07E
Q+pOTsgLXEwXIvOND9ZtL4Z2+gKzyX7NiBujq+2SXJ1C7lYc6Uf7gyrTCfwVdAncVPI5egN5kDcH
kn3kYWwiwHSoE/RYsaiES1fcU2uA9JJOsG354k85iNkMJaGbYtQHltqp+K5SmDIb+EfNB7Eb68jR
YVz4jwB0VFPLbyfogsHPcvLr52s5K/PQ50FKXwfNkHdT92Er2c2pKoe0XlMbi0BCRwoePB3syaFh
qiHI79WIkJxzFIPvmmRgryKEITJ/n9ALJDwQLRPdCL62rbblbP1uU+oek8Ewt5CjGC7l57j1Ax4i
XDEZzH2934RMaiO+TumgtuQCd/ioqH6TyLxpBiDZ0+CsoZ/fbcSYbz92Zm5rOccTdeNYBUqGRD9l
MOpMMstfV5yX0zkh11vqxfhKbqCAjR/VHlvf9SOXPP3ctVjgjBpnyAv0BdZYIUeyFT+QxI3/UkbS
rjXFGd30lKc5BWWWfzys6/vdrRLdJJX7YAb1KgjAJg3UW5r5kj0nk56+AzAXx0usANBvCiOyRRM6
RxNEc6niYAanrSp8bwDIdo9HCclb99wpATdIB+tA4S9iBzGw7Npb10z233EoiFCJK0Fw3QuvsXpy
9dUm6XKI+QDHOFA5SWAP8x7L0gUv183Q+3y1oeuMerPTWon772T0j5mU/frWC87eNPj1+7dVhRjv
b8jxm+9tl7Kj7R1WBdPp1QXdr5hNlBtmDN7DHElGsFokGGrK/2snnayTre0b4jM751wF7Eq+mG3W
Xc3ueX4wDuQ6wGNuUL8hTWpY4mBdlVOheT121enyLElVcaTIW5sQcLrcN0QdSO9O3pvNoERdDgUP
o0h+CQuRiKLYZPaCrKscT6gejDBul2BmnoprRuCN/4L469FFAYXNNacqbDCUD1AIhqwphgfyJmZH
8onhmwPQVUbmDHAIBZ69Zz4QmGHKrYXmO8ArXWxebAQgDJkCD3rLAEz8UzB7hMgqr9pUuRM0Zg0R
vMGXclwtYGD57oXGpNDka4lwgZVLGOgwy+KUUSUUPrlfpHUpDBoKwNiaCjAUaqEekK4T9FyIH6An
8/HD2hKXluKZtul8y5zRjadSF8HoMfqpDoGCtF949u4HdYRpE4M7o94zLWKqIjWob+yeyHx10cjn
DmzWw+MC0WmD/vgxuwo9wJlRoxbcVIDkuvPUpb3UDrwKzKvcwHtsxIzFdyke03sSpJ6Sgp9hkDxv
6/NPINiO5O38IL7IM53xrirrfkQbgBwj4Vr3wbMW4of5XqeUaNES4eqbE+Q3qbnRpv3Kj8gECY2d
ECACX8PNM0zxoxLhvGEzJneoccoD/jBNNQB/Za1s9bIgiv/EwyF4FKwsj0H+GCFbPkkHO1I+iq8y
LUu9zM0FYjVVTgjnICh6YFxOdBKOHEDt8qTtmnjeyqErZsMWI5S1e4g17suTuN4w8GIFgDkooo98
cdgWIg7amtJWZFOPxM2IU4fH0CV2NElPIQtCsv8N9DQmqRkxy0j0wrnh3Q9h4rnJbyxFCMpPuX85
M6HDEi2/IJ1n4NQF1ESPPKy+NyT2az8cyLKh5cGUkLmIPu50kzt58BCWm/0mEtbH8YErbdZ52pU+
zbZdXoo2kY/Rvnt2E4i48V5bmBoOG5QMEuXaRFmky/7sNSh1EN3nwfoU93DtMdrjVYFyYiEd0nUo
YHdWWBmNjtIUgATKWkMlXvlVwT42rvP6p8H8TyOTQuCAvLM5B3FQTWkF/Gs9MqZdjJuJaX/kzMy2
mGlkikxXL7GYlbQl9eippjcGx8zw2Y4Hcbpxefra+NImJy68vkLJyfX84Xo19RIqxOU+jP6kq8EU
jZvkV0ccP9xayn2H1BhDY7/RDwvhBxw7egIoCG4Oj1UpwLA6oTEVn3SQKnX2Iug3mazDvR/NlfrP
GDhFIJi3VnDPGqS/FXi5U17sKDnKuaAGAUGCGP1/10DN1hABbeDMGsIVxNgSI02almpWL3yseXcy
aOn/RoaYMX6PgvsC3jmTzyMJQIZPQyweCMFRvOYPgCx6Ear/xqKNLaUHEaDhFeskgwxxBlCB5XXC
kM8GhIkUBD9paLf0p+y3izS/goWWrExX4s5O5dvn1ZwAUN9INIlmQRQGVmnDAQQo7nDiUTZnKbUP
vzSbW4yEyW4UFFPDKMou2W2bjBuz3Gjv518NAmS5EJdkGI1uweWq5er0R6QEGXFtBhNWws2u9/bV
G7I8ipG8giNlMXPK2i4CqwBcaLkfwBdbFqzIsM3P2Z+qxQqjJ1DlZp+KEouO6ZtpDvE8i7D9un+m
1Mcir5dlb5RD4Y/nomMw98GmqbEiHva2jbMux0fahzCChYjVEWWrzYbYqY9vC/LlPCyeS6vibd3A
8mFGrpwz29GOEECZ3thwtb9+okBkjx0upqssRU8PjEXc7uat5tbPolk0P5AzSorLMANZgRik6tR0
QZ3TNGo57FNXsV4KDukX28Z5sY5kVDSXbPIFHUUBnJCleNGtwHKgcTFNTi5PAgr2X56YayDLBDDA
G0SON5efQxfqrZMSNIhqQ6aNfSGurKdNTQWwVu45xzsBMxbk5p+6fcQaictpr+rclKbt+HzOwaCC
Qw60iokeJEc3CCmFcJfe3X/RuSNvBjKcw856WlF5w7bIiSfLkin96ZVeb+Q+ia2+GITHgFlAoLHX
FOV+W0v/0hLDg0O+SBmU9nuF6hgOCLCATwTaIxA/hWebhimpacgZZS5wtzg0CE3G5s3m3gvvmWBm
YBCAhHFn7+GYfMjnqtmIbUQzjJ9/q2wL/CJm69iEwxHmbD7Ttc/Xid4fuZsdvM80UqZWVGdFCez8
uuRmGY6/0WrmB4YzwkYGe8UeAOPT3B8Rb6rCvehSU7x9p4h5Rdo0MZEF8ALiXDIbO4gbi4AKZJTQ
ZT4DsgtD/GlThZwZGK6xXpkw9l7xN8wULhIxOMcuPvu2g3dUA2zLaEHr+keFIs5A5Uvex/G4umYZ
X23j81U3Rwt/gecePRIiS30yS2+Y+sTB3DoAf9A2TrK6xNhhz5Urbf8JlcO/8eyosnGldYnn6Ybq
U5hC05lVPlMXk+UhkZK2V6I8CKqdQq0s7upbPpB/daG1/dSL9HB/yHvB6uaYTxaG4eVhBui5mwqL
i2QhrBVx1bS2LC0x+A3dEObiJWmEJnzn+A1xu0pZLi+odA5RV867ScQ9id1x84dUztmY+sCq3AP/
9/9jbW/ZTfzXhi5b3afz3l5zVVglEBLTx4npSwEVBk5p6prAJJr/7cgDmL4pUXpreqToWVA7dYx5
FZIdUNywk0YUyynS7j9ufeKZ1EIXqsY8r008RFW92WUJ5OFftQcCJrsTHbn7/alxOnNiuONFxouB
KLCEwf8YDz4rr32niuPeObgfyBgaqvuoAzrQWRwQckezFhNoPznQ/AcNL3yxN58N/qo/HLplu8LM
Eiq2ZjU6lyzTWicItuvAIzOIaPbFttAqfojGKXqky5OYXTuKfUaWxTz9bgzX8f+iGi09NFnlSRi3
3twDOvPYz2AMmNqvE7kaUP5LGMS7iXFDFxp5bpcG6SbCVaLKmdYO0WZMfGHXrv6XahJ7JsiA9rS7
YdpwE10etz4ngOS46S72u0N6LZTXnNbbuh6KEwglH7v19LowlEyf0dQNzdhs+xO+08u/uPzXRGTo
faxnSYl06LeFXexiBCkxsEB+PhBNRQeQi/LhqMJ0fawWCSC5LeCcSDyjktpPIZvuUt6nFXylBxNu
xwEuR7QZkJEFzBkEdvhHQfhf8QVktF5tNTNf/wITPPvVwADcAOHHwM8o5O8kMj7+LSolpMQBgCJ3
L3aU/0VVl0JzawJ+me6MHQ41p7SYhe5noflxsIk86Lww2SFN8+PC3ohbF2SrbGQeGd3B1oen4oHR
HE+9YcNozY3yIhUZL5vGXGXE5qZRRu5BtcyEyPWr49uacV5idBLWfAneG4hlLVgeQeyu6O/eT2eA
pUIFegeaxJre+kJG+LzjcBP6hjzG86e+/+NafPCtJvODUXhVArQctbxhYClPWq49Akcp5Y3QB75s
36T5JgQ79WT1YA1+9oBLRooQ9Z7GHErZR8E53J/gWfs6NhUZbr/Pf3Nw1V4oOShQC7NPdkDWh6+P
7exAc+SX0xolEtOwtvwkVG+PM9F4tvC4AkyDhKSa8sUIjXkRZKbsvl9OXrgUL7HOrYrf1kIPFUcg
xIJqWt3rZvx/MKb397b+dsUvlyfoWMqaWPK3UnwNTS/AbCxhAm+i+fmk5TyP0PwxylD4bZjmPiU5
rTIMjIT5RL/DRSz7zCJzCAejUCu4wtX7ojUiPmmUFZrdTeMTxt56GPGDgijTklm5BnaEGRIDmKLU
kzeTCUdrz/cloUHC46M+fLIbBkifzGHhNuR+L5RhtPQDQU3kyHbyyxHa7Gok0om1k5SjbPU0q7o4
m71/dzF5aD5w56nmfLkDnWVSx6m//aV0PTm88mYFKkWLro/Qk6JvtkI+gBxUs1/U22HcPvdXDdAr
/6Fh71dBssh+ZUqiz5kwpqc5LeCc4fvLU76QKMWe+iY7qd63PTwqIPH9+o2/QqMa9jgJGWJcbO6W
HfaLFSEkohaebf82lRdGNlvd45q3K67l6zjrpN43uVTXpzJkxkrkG7ynRVCr90vT4RD3T69HCKJ+
9CjeLFKFMdn31/QDrQhA8c1qYKi7lyrmwI19+99/rM/pH0QvMZtLAkSQPfpjrRc18QTop0r/XCNi
uONh9kSY1aWqCKz8BvYix3Zn5JVumxz43mwzAicGNdSkWWYb3T3vpCjbiCrj/X5K/7RiGyGzrkP1
eQVhsX23vWVKz+uKS6uFthZXU9qxhDzD5lSUeDyLqakPNo77g6UgGUX30mt8adjgA2ljGOGNuJnh
OJe68UUtoCN9BlwfpkFWrXLNdu5sbKcp4bTJpd5HvARMhaCqbnRverwCl0qIYz4aiKsYXfbcd03+
BixaF7ikZGZyRN6jqBklrss3hr+Dzxvog1zB20vawnRViS6YKnQngTFkrWowvDurYNGEZXopyxrc
OGdyZfEXMPZNSRJLIW4RdrqWN9aa8JIG8wW3fAEA6qKBfV1KSm9AYsePB4n9P214gQggseHnxM8J
CS484kPeW7pNY2q0IYSzOWSTEo0tJu0Zo7VafRK1Azh8AJSY5SsuFai7kz92nuiyrh9kgLe2Tva+
ec3bR26+id6ypyX2PuRSs4BMeu60s2xbWtDZdukx4UkAXsPdYaFwI7ZsvJzXCJc2yJelfny4IUzp
ja7L72cr2aT87SZEMOxQFmRRli6WozNsik7vbyglbpPLp2EMfQxyM23T72e9wtTMKjjPrOaO/tLy
1+eoHO331rJaZtpGITiBlTnMwih7TjB1mKGYkPce+mizl8YLhCPhxer4mJYHEJtrGEiRx5jjnYK7
hWkmTf4pJxXe2Ods8LKwh85BZO1VyGLarah9KavoNOlX6a+Me/gF1DaHQ2exLApWPG7SUZo/U0a9
YJ/3Ysq6JiCTwhJ9OA46TNtiJFpMSQfgA5DaOWqhrWesS+OeareipOqAt2LZD5Vs6UW7375nbPcG
VVr7HTyu+qKuEZcEKsTccAployC5rllgjadj7dbw3dRe+CsLuZ3LPRWy9peU/1S1AM4YWdNkCooI
OgQudA8UpP8NkuS/7w7/seywxQS/gAXAIx3tHtgL193kAh6PRkNwV8cGxGbcziZFIAlgywHxVCiR
4JWGh9HnpX6wL8lHEBcsmoqxHg2cPb3rZ8rOiSbj4FhBr5b/C6eJEbIwaCdjBlqMiyoIdnouzXFH
ooApMUie6uHdcVkOMEur7jS5D7jtDoTVURCG85JNfUQ/vtq0U9uKZiGJAuL9VoII1yiW16zkKXGZ
ld0I4gmF5wo77Lu2VJk9qUjIYBUgu3Hhb6pgdMz3SuMzETUR+iATJtDBhFZQDbwt0BrOOpeHdioU
MQ9cHnfNoe23N9oNJBEjITJ2fgTVlr/mD71uB3zrsBlvG3AlzssPCotgeY2rTnsw817+mJ8qJ89H
5XIa+eFb/Hhiy66jXanyYFS83T+1ivnho5FYRtKgesn4GL2QyA5gSpud8rpZoX9UiEhnUu+OuZwd
gfzgTgCTVshlE19JA4zBTocIZxF0G/krOANZrDmR5NAbE2vWB0xj+ULNJKKk7cFTyjp4LOcB3Rrh
P+UlC/Qe3pWJxP77dpeFRr0Ia38MDBFHolaiUtmxZYeRMI6PQ+10Epz0lh4/3yrUUmUa5wCr8aIP
H98i9ifPEfUFghi4vttehOPYOUiU3zUBQz76EdsrC4B8Ft+rtFh13AKuIDjue9pZjIu6RISa9V8C
uOaODQyI9PXeI5p1Ig59Meua3f01b8GGMREeFxnCdZXiXUYTjmqhJlRyIL008YOF7Uey6pjYdH//
51UJ85k4OqTBUIZuSa+FMsBt/icfqlFW8yLOB/ppxZXb2KM0WCT79zNEwhPBP3itthK/6ARhBWVq
NOX5263Z4Hq+dWBBd01a0DLveOwXWI4Ryk8WSmCI3op7J+7HmS2fTxoYtKIxxouaDBLIqDaF9mlM
wTWWfHgYIN5hqRXVvygZfAFWYLBN/LJv22UTXV5OIQmp4PhbYZ7BlqNBmKwuCJUy71QMXqKQSmko
DLujum2Jk3ZYVozav66BTHiV5WNaiWusdGU9svuqvtjCow9/OYuXtW92aeVN5m5ei2Ir6FCUfvyO
dxXZxx1dvsirF27SpX+0Epo7qStAygMSL4HU96NWz7CfbQfjb+uVHpYEHgwDNJsJ4Jm/yVFiXW+z
9AhruxARSYcqP5ZOCLT90mB00tz3rHHkaHIjW6mDtouoNkfQAouBF+lBIY7hGsSVbsb/1b/gQirT
IjOv7/3nKedattUVKynYXrnpDPyrUaBkyUOOdB7Jw/4UO1bcxWG9Pf7h/8JIEO4BBB+t8k6Q1bPQ
Ht/PTwXz5GO+M+Nyqi2a8uxJgikUmj85zI9aitKLmf5SMa1w2FuMIqYGuC2jb6kZp9GxH3Ue7f4q
UiPfTT4maHCAPo2RnXXJc56svyu6V9aXolGkyb+JdiS+ZtxQ1HkRBZb6ewQhYPad8/L3rYidwwVC
VqwWjqhKfrgVpAgz+aWz2b0bkd1zm+9fCTSa4dxl7z+vQ6Tdm+faYEKpWfJqqxUmDxZ5GIBiOb0J
YDncTw6e7xGNiqNIxh+ZdkbgoYlKfWsoiSNGX8Wm54pUVIxIj+ALz4/bGiv+Ms8dZ+jRFdkT9vgq
dZQ94t+K+Itymq/0dFZ8U3zgoc40igD5KHycDzoMqz1s8zXHCk15L9ve87N3hg8butrsGFXaMdC4
jbS5vwo5d8oXt6WKKDZm/oSVr4PkElqLmL/m61MXMR3Y21n/Ow8Ek7DjfiABlk0lEq2CyTjKPk7x
0Sdhs82FlOSYafefuY0P9BMh2sd4hZPKqevDFfXD5F4z6XYI1XwkMI9+mGNEwcBrhQRQpV4vOhV0
HTdQrvv7NvFyeLxxesQ41FK5RugD0tQMlRG+TO2EHP2GfV6wZUL0uxOkqFwqM0tNAptjAp7L5Xty
bb1uAVyL4/ITrRdGKNzS5XJV/qrxljHEpMDVdr3COUf8InVWLlEpOFFk7vCaACnlzP1lCTXZIEQC
J17weXlooA74p2iKsLBq6IsRrjetNjy/cxsskwskSRhhwmvln5RCq0tcphS6LivDtjTU6X02cvM2
HDbMYrch54ol25t45Fq3tJzvtTC4aKUUrclC/jv9doIYdy2Zz4YrfKg3hUqhNCLaWXCZPo/K7pJt
DXcOyx96DiZgAbR4vYV/oV77AANi4zqIA2siIcdQTm+IgcLxMKY/wzyzL2/RX/UV5S1BNzigGFHu
UTvJoe9O6iWSZYd+1enRcrr/Wns/8mg1KzwwVqbzR6M8Q+sYytuNdYsXubbs4H/wuVrWDsRxtZ0g
pf4431lAI52MZHp8YwVMySFlzZaiq2oz9NjqM47t0vL4khJck9nfI2mkXFzZ5ITd9Y2TX7/ZeU8H
QqLZgcQOdEn2/H34s7XiUQMwaKOQioNUE8VdRHpD+Xfd7jX0PNVW0Yn3hNL7m71IvxUeJgTjpIWY
T3KGomnfU9uzNx1LES6rlKqKDhlX1W6058GLgBFq/YSWidKXrEiWi7ZUeweeWVpEs0G0e7uyenAD
tRwz9eU4a+OGm+i9lrdk2NU7B1q05qnv2Ic58kezW7qLi9weJJQmeq8+x4WMkn2eVux3h9t0TXBo
JesHX4RfHBVSbHhE20fHOJPFrFha15dsiT/mUS1Ia+d9HJZbvfI8g2KBEVC0WHYftCchl+8ik/D4
Qk4NucY+0c6coP6YmyeApO2uNKZ4BgzqTp/ZdzYawfpEqZL9TgoUxr/BG0WtRpPeY4EUzWMqpvhk
NFAXKRS8tVSLMfZkczzTxdcPEQQNUz2h2FF2ysecSPztiRTavmC6Ftn6L7EcN+l8uA3HaGwcRrMJ
FcORrYFHpnrjffLkhM5lSF3Ow39jsIu5psoqw7ILerZ0OuKo/TvIUTn7IG/oUADemU9GBQ8oVzRO
KeVx0vXnOXq595SzYPPivFITNRFpQ25Zziw664fbKyvIdksiAbk3bFz7dibw6GdFyo3hWK2K2Zfq
PGH/uOQGLBx2Iu3hXdZPAQovb1Aoz5zedhaLZ/BPx7OT6WnecL7wQY3yc6ZRNAJidxXVraZCzYOE
8ckVeKLlboQFNjADHldI+G+AFrncRbXQEfRQOxeOA+hpaGEwbhdpe6zmyfwSGTFLmYu3/X6buCOs
ZNe+om6bk5W5g/IXbAmR8k3P0Hf+OwTGs2VUskPrxfu5SdcohCR5AD9GU536jXGCmqs9W732koGk
s6hc5cOhI9+sOk/HUy33NtVVGerQV5UrxczV+0sAurIWZkGNm1wFNf3OPlENtQa2zT14H/VM8HxB
2zR4TifUB0bTL1dpTYB1hUEoHZKfEMnJn9E0ooUhWh6pjuJ7zlWF2EndQ01Kp9Qiqa3vJI+LCI2V
wK45EXYbE0AwB5jOgzI06OEMHKqElKmoJf5RX2qmNiVv1s0F6GVw5FLInvlYOKP6oXzz3h89gz5k
slFP2wWtbpfsCNPcjGMQhYIQYTmTCfAvq8LpDU6xrOTAxm4FxqtumHUB+9FfFcx/Uqp1t9kUGNFU
FbsSDe6fYdt+bckfsRqYQwiKmzweeQ/x1KYNL0mqKluHa6wmHVjTr5v2HlQovUQV1pl6Z3tqcLxC
LXhk4Hdguf3dC7A0bMqbdDL9x+a1risSUVwy7E4IgpaEg4NbPlkastatnz/n4okCxzvs/8ov4kzC
JYBOzb/gfDPfbZz3Y+uBUxbqrAIDnPqJx2uawMjUIxOtq0IIXk5sRbSP2BS3UFMvBYOCcXGjiwXN
LRbr7XjK6VT0jvCLnYV5BxAB/GN/OlZe8hFKmL5lv2SzC6cMdFKSG3R3dn0GPTjhnoxhV0LwFAZW
WibgTrW974Wlrc7gIXtpQZNNCIalJWOdVC4fOGNd/fC/h1U7fbdzYDhBpnsxerqZvL7hrvzBIHc1
zxTPPgU9ayNWtPgFupqAL//GHm+2a/0/NFPc79RgJF53CSdTVR82cys1u70MDvOBwmoIf2bm7//N
eVsyxxm0l9RxvZgNhVTYA5UsHkjVK9P3c4GATHLgnO1pk7wjIA9fB5lTSaBylmD46HjAIb1aqfrK
n2wFqZYrXrBWVwDY70pngz0oXzImfx3qwB+/vL3IE+VHeKSFm5OVd6A7X2FFQqzIaZhdIHP3PMjt
fWvgY8GwtW3LSW5C8Czj8GTSQIHmqltplzJr2a1qSt3gkvg7xDiFYilZQl63iD/Z5kvrbL/arzA+
FAJSaAhXfAxTwGOSn6cVKLahNaiAbum/RNuBAHrw0oJlL10DmO956ILSq5qzIF0kQJ8TMzjUSL2c
ebzGOjCuqXkKgARz4NIK7a8sDiL6dp9oNDDgTLgCLurzvjVreKyK+rC3soOxq2OGnJjh915165Oy
0hh58yPvwaRjn2vKUxzkTXwK8yTFOEdDtVKQspNZDcpGAPlNA8F4h9l/6qiIaDAKZYIwbx/zYblI
4h/cmieKDyPSxLyCbawxtV0GjCDlu5syOVdxNh/3/llpBzKN9CFFNTdThJYadqBSt/HKRvFiLFHr
Qg/q+Vi1/kEg5QkbiCLKFuTcJATcgyTa0ua6IucQtuVmZqP0NTAO1MkI9vKQAqUHjqIOC5NDepJi
PcZBjedC5ujh+pgbzPCRyiHKsSSpoOex3y3BDjdY8fyYuuq5jIz4kE7OaOlSdIDisF9V12PVyd9/
batNZYTBO2jtt0LYPo6Y2uaZwPE20IcKCvbv4in10vjoukYKyG5ETwlqlJ7drJKBvvu7NwrOtUim
2t2ahU5pSf8Y02zxHMiKn0yEIfQ5/BR/chNu+7auNQs3XxrRHE7vBePhJfTF40JCJmiD6V/ZLg0p
IVBHoELs4UdzaJMP6L9Z420yfX/35fvNtEA3taXEKp0kRnporYHn6rpCgkOlbCo1FChz0/LetMIQ
QVLnisa2JAoia9an4keO6B1DHm6zlNnJv/XWIZGQKgubEWxXXKiAywKn4wddFkXc3pAfF3skgB6h
N++aGLEkxb/qoCprVkIoQ/tmKGK2p8VcAU1wa+1ZoNHQgIICTGhy/R3W7QA8dMiZRHwNJL8WZ607
QqgTwb28UcpVt7fjrX95JI6MQw4MSarsP+ng3gTnjgGTWIX+dwqzGasnpe3qPIuwr8aB28FzkMvF
+aJLAfXmtEaB/m+HVMc3vJ5CvXLeOA7j9SiSDRkI6zj8Hv72me45KistQdTpcKp6UTPoFVXfcWoe
nPEd828cIDZ4jjv0J91hhi2JeuGVrPmq1Kd7IOvjEpBWa5zWDqB5i1KNlMdkCG9oN4/ibLi4ESJF
s76fCTzQ4lsvi7FFbdK1xiiTIuE5hwABnrsr4lbhBCtstIM59F2gxk3MnStmD0JVp9w/OAgZD69X
AroRcLosHdjjwOn6NlaxZdy7a4KB+Yzn4X688ydOu4vTMTJt/KUR4ovMXS/P8QFXx5TFp7jdoLD3
HmBNmB73N21MH1kMB0i+rWVO6z7J8MoKxEX9usK2Wlg/MHP1wI+ZLnapT0OgpV2cYcFzAkFTU86D
QvfbbWDvgWiRyJxIB0WAlGr/qtUboVn8zhrIEZqzgjFhoSp8ILfGsmBrGUfgkZBriwPq10G8HKQh
G5DLOGduMYuW4w1SJayX+Y2tKk68TrMt24WOUaAwDJDPxUTwuHemPtVN0567eoByylpg3FW54mzE
mBHxWVJ76YEusEB5PtezAKBILCyXFh1nCBtY1VlrfVOmkyeG1M/lHprLlElxbG92DNx2MC2/vtfx
wJa1ROdhEQdTs8ln7vy25ddK74eTzMMmWdEsyLuh6QQ6n9uhiutDJG9vIDvFE65EFus96OeGf53s
HUzy4jA35SfSD/SWmhWCnj02rYrZQuwUuUkhSbqEODw5c4hfE0Mh4rZj3Zd4Ojy12v2RFDkt63CG
BUvOmX1a9Zuz6VGU7YM22yNUALAZsQa+c2I6xd/Ba4crsuU+SDuCySOUN0QJOW6VkxMt8oe5gWVI
eZ1+pkR7S7JzVwxpEoEJ2qFTukoGSAFah8nuIkqTcqUiKPS9uiueURPN4pxhBWwaf8F63qsVqCHg
f6f+7veKWARLvCryuSJFArjVmp8uElDT1no6aevDp4fpyTfJvMc+kM605xbiYUH2cw6aFul5Wk4+
k8wHfppX/LJ5eAG4z8WkPGK8P5IDSfG5MoyK4cN9zz8cVz4t5JhKXRS7TKMqyLQH6RgKfUUAN3FR
Ly5k18VQNaI/3jGsO/Bnv9xhjO4Rns++MdLbdgORgMy9A9bykAL/cwI81Vremnn61v5uPeZ46PH0
vAzv6CAfYJDJ5oKYiH/NsTNVWVNv8rnKBzeV98c2HKITGQHri43Ce6Qa4Huq+YqJhqUCnhpK0+yr
Dsa7sYWO3mDmFOynizg9PPb8QV6E23mCKNVD37adFKc2m3bLS38614ft4nD5XyIMSQXsSdHsc8Lq
NbY+9o+pEfBPentg6VAO6siywtoWKJMG+40cpTwpjbXr6q14SdeIt65bLyK9UuRt9D0GZzT8dbLq
WtWvQwznhPlzuPsy6I4M4dnv7EHokkVCnjtYl0hjn6RHqn+XqzIner9MXs5pGYzDRYpH+P/V1y8C
GUlEMjCoVf1yR+DWFDC4Kp8Ci1mn1j0WWtpcmt4H1cp4exVrmD54nQw7fey0Rw3C50LJiLH2MS5u
qcNlcuIfrYh456ER+7OZNl78xp1YO7jpPwNyxYQD3id8hllbrXYGLjnfoJL2woUNxig4/RoT6mJf
scHGY+HAIkn73FAqxQdHPGYtgxGCANUluI6QDkPg5jAaCwPrgnCljyEny+K6CPXKA/zKE34kWgM4
gfhJ2z3TmIk4v0wCwwXJf+f7R5Tb1kvV+8iGFqj38I7MEByTddS1qxCvxGxbHtsKqi0gtTkZpNcP
8nP6DKap3suogjNgCaDR0z/lPHOQ6UuH/WgwzJE00DdvNxa2PQSE3qvGGCElhwez2SYxQBnkh+yu
DEJiPxuqNXNO/82aBBA6H5zFFHehq6YaiNrrqy+nAdk6lDQ4lWzqrHiI2h4fFv2SsoZcu9WiBa+I
YNtifi7n7Yxku7ssdWJEb9RihBYo/6Ugljic91FqnoUMTICdCsDZNowjSyO3pTMuHGdDBtLzg8td
uHbROxq8dXTksHjQQBjMlMU2nG4pwf61I1tVzSO4jURzpqDWUPFGDZixhJ6Zh+7mdvkAV8p6DCnG
0ZdZYeUVn8QmUlTtmiNEN8ykfOF+DXTGJwXY26kSRMhpdLXucOet8wfcZk6d1Vul12IIH+mjAKGj
ZuemPSb0C+4A+c0YaqpuWQ9ChkDRxcpCKh/o1bhNVX/nGG0W4FB3dAG18GciYKoBBxeCZMnzIA9O
FB0L14Qs8OC+mi2orAXVVQsonZWrinmceq5qMYDTxQwn4P3+CEyRY4mtQ0KVKxDWwYarF48IHtHr
FkAtvjs3JQ+iLlECiuoNc/FwHKo2jidpH7JmHWfNlFFLoQWGDpU0ppeLzs74KjEP2oqcydP2FWrr
kWwHx0cpysuc/DdCsHKi5LA1aS0WpNpzGfGUiaHoyfSa9jK0anlfnFD4kUn8AqF5Bllpf0WjwsIk
PKY1HmPqkdrAi+302LvjjiAetE2cbrzGlizLuSyBYVQokcS0k216EnJkj+Y3OnUOM9igtOoOU5wo
a6mTQGHi1XfEyn5G9hb+jIz3fjIZRjk6A3r0n8umr2J4By9lOCklt+sQ3W4Dn8OQKc95xlU2Y21L
oRw1LzQ+d3erb4GSD+SE9U3SMuZrLLXsKFp8IA3U5YvMwWiNWsRoSb574bBbrTQElbsFXsJWDmwy
ucmfg6YrECSZ/sqGtR9s1/hWyq8Lh5SHm8vQ/amne6ORDMpIsgdroXdqrq7ezbOFlZOW9cyS5vz5
NC0LcRUvaddzgf5k6iwDd1lngEuoXiv4WdUNgU/3D1NYC8CnPXwh3Bxo4SauyVtPNT6ZLi/lB7ZE
MWLNCOMxgLdvsTFyfRVchWU8ng52ADxcbIKxcDLoLSBaaE5f2rCjNzK95S5RCalP630SmQhgeA89
UC/bqx23cZqMIqof/2LR3QO3Yu1AY9sybvU9q+j1xHbw93bu1+R2HvSk5cJm9WcW8icUv6hnmLfM
XAMpyVlHxuLtX34jYAidiIPnovpwV1dXgkyAp5SpNc2ZYiFS9mNdHSnyS+hSlLDHNqeePZpMVP6y
Q5mHK/SjhlbZ6OqG+40fDRRuPtLmniECXq64YfUxrBTNHuMPuR6ttIOnN3m2g7W1FRQamWha4p1C
jdbHA7rAdyuSva/jvqrGUCKAhvaq2DKPTpd6dfCKd1E+OFGLqqYx3ITLm0kpMtzFi8KAzsqH7Pvx
V90lSYvNGjsmcifNE0Oj1QO/qnOm20E/oLLJKjRyuO6OcDL0kzsKqp5jBETd3x4mWqkRQEjbOArS
iWgfpc1dSPx6quq8wJm0Sd7biCmMxFceFiBlxWKzhVn83gA28u+QdivfiFIA7X6xer3c5TbiI/Yd
rSrPG32jYZxMmpdkxagpFxGgoTTt62W9B9cDheKX5T9x5+fkmH9gyP6KeIANYizhuA1bMcOiDo0A
MXqPHoAdrxOIx6+JYmcidqJYbhBopXQw2/e2rE/iZTPxZ0pEoK/Yw6uXNlRk25pcOhsuoNcYplOo
DOZdPXmG+RuZK9F7IGWyB5SkIAy5t+yIqtCSqbLGjpSmhae5BmrmGHz2IDQ7cJKCZEGYu5j0aVk5
8HbKLo3Z7ORLfPcrq0OI1QhQItXDEccxPo7VqtvwNzVf47KlLRo3EdAO6LGLeU1olU+Cy7Iz8OXR
tzCsZaJSrvkBGosoGlHDVkfyfSzY0MD0IQZQJXF9J0gkVqXRX6iCEQiO99+cuc/MjXoloBuRpXaF
2anaQ6PIgAr16xDgpYzYBV2PfFx/PT1PKxdqO82DiA/rLb7onJGfyco56gI2O40lVRclFzzXBewQ
CArdroECrcJtBTOk5D4q0+49iuSIJGDRYZ5bVMPays7xFpiWPD/eRj7YLQNnDiqOIg/8kgVjqBUD
cGrbbKUnW7KuNUMDEZ7bvQsLs7Dmv2HlmLd8nd4jHipQC0op7MhfL0sZkwH7+B8eDzT1Ihb2AqCS
gi0NZiO4cXs5KGBe3ItMWR9czrt8IbCpUVy+KohheqOYSpfSpQHwBJffyZzNNcDNEKIb2IPNARG3
Oku0YXbck9HVPkS1Ej3wOlgUdrtC+/w4RB5x61zXcrMIaxZc5zrLRzP5ouVLUFG/g0Pq5uQRzWHo
k4uNcHotkmLjIciUVmLEeQXwpYHxtfDbZ9suLYqyEKhYVLNnD2Bhckuib4kbT+U0d7mMvuYS2tyE
DqX1uEz37F4KOcIwuE2ijTZ6kdW+xqFcuqumAoWmRf7rIvNqPKoNdktbits3fzIghpFtPpZ+L3v9
3toIyjp708LRvus5YG95I08cFMMGSol/bKORel9EbX5eX55PipoiGQCNO44K7XHrR0XZ8olcF3yD
XhsXKuhpmCGH9n7h4r7Knb/UL6XLJVwAar0AbmlU3qy8TYUegpa3DeRA+kmTH6h1XLaYl3kL9yqi
cES6Kvqewq/GDhp2cjXfUqU4AUWfqrzp/7DASYTkg/H45dHvHLGBRJQM+twoaGd3xxqX4mY1QyGX
a57fLvdjsLd26kEY3DQLm0ft66mtpSYCb5DhM42+PQz9fjj1Vo7/UvlRabGTa548orvx9vOjxuuP
XV4VXX+vjLQcTT3bL15CuCX0FNxV2ChU+m7R9ev4wrTxVVlOEfZ/XAqOL2U/z1xB7DlMue06LDRs
8Qt+0XPJ4KaKbTLC2KhHEGGvBOmvhcDth8ggSneeKulLVE6EE+BzKPG7eKqjyxg49ITlcYQdWt7+
avDZkQEBsFxuYc9PrvAAaqWhlRkSxl88EzL+IBZUOhr3/OwoJpLZubwiP4P7yrGUrTHkJTTelzm4
Wa6tx4lMgAc9B8pMLI+kvZnhnGAbktDN6Wrs0IA+OIVliUIfKnMOvrMRJ10JnAz+hIeCRITVZgvM
ItZ/139u+SFho/kK1LTblz7XePBeCX3pGU8Ug0blN2oshRPfphb4W5My3wCOn2estOJf2GfZQWnq
B3i6JisUYu+Qegydj5pVj3hS/aateT+DLSAyCCSckrIyhFTMy/9rGhixbnIo5QU/1JU2ekG4+/Pg
JLGiP4LJhHUqv9EFV+ta30d3DnvcZnyUKCJLp4Vm85umKyg6S0KtG06f+ou89KJNw/5dcC7BwFFY
u2ouvcTRcTKOs0Ue/bBu3vOZ6TX0p4ZMRCTo/PGgHscbBGH/p+QFo6WNUgQBTwDOL+2h+J+hSGY3
f87r1c2g5BW3UsW2KNJJZVt2IXR/QilUdvufqSpJTZ9If8TCBGJMM5yJglOgzHgokgIznTUny/ti
HMcoTdxpecjrL802vUidvUmBUbE0GSA/WptPymKkvE8Y5dqHn7kZUqzwZOi0Thj+u7eFtJMYmUa3
c/aHEM535VNEtLYJcUj4+XhDx4OnXM/ZvpJ4ATKFfmbPYQF4dyNUVQuA3tV3kU7Sl2apz6hOEr41
YQ5nziJUEmJSuO1Igl4uMrlsuT2keb9yv3E+xDzfZujk9zvtI1hWcmp+2mXexJZrsWRGpvfJhGqu
3w/bnGUQBePnadY0p4BQFgG2nAcNr71z8l4i/F8jJXDOS51KIw+Wbt1EcUYOwIMQv+Iqnn7LAtqx
e5cdhfB2tduAhaRxFVBRcl/U6ey7RaMP9GGIxcbuUO/3t2WuMsNZRekp4HxUsYxHYkTY69Jmetqx
xXKOMO/za59z6+8Rdv7Y7M7xNlzg8WSmRyH5cVh4bpeIA+N7D4QPymmnbCCLiIYutjVBR1iQXwXo
I7l9WnZeVLSZto3Cx/68EKy2F0qtAmeXKZxCVBOm6OTy3LBJX7V47kdFqEvr7wuW1NHGSu+SjdH4
9z4VtUvHh92+FhQTfyhekSe8vGPTZcby3egu0K4bXbNZJgR3tNUgxrlfwgcKGC84HMLveXvoLW45
kutD50osXbyOCfm5qL/h8Ljqh2M+4JmNJsa2cSxFOdIa4TfdtUs1XEIDHXtmoUsBErlqOqKIKjEb
D4qHbjCj1QvQ+sQKNl1D4vSvOZZki3hISQRtpstsgbyb3ezvUtAZRvgSXwXwjWuqtK0G82PZVrgB
zrWAZgOnwx/JnBmcwg0VRvFOWfQG8kJOuX11hgqJaGx7reWogPK+pPDVOLc/e05mjbx81Ox1UCrY
/vp+Q4H4PK/XzAd7As7ajmkgHKu3tn0ywU09KVi7xFf6Ixyj6w0QVdvpKFm2EQMIK6GO3GAh3j7F
uMvWd87tBYAe1m1NNGpFSG9MqT2TU5TzG3bEiAqkj2deh2FtPJ/jHETLRAelVYujXWE4bfNgOSSS
eJHg9OQi0J1Hn0Y7o+Pkgj+eGbZ34yUpHn409NWC5D0QA74ubYlcR8PICE3RfwQ9FHA0xrGZmzc9
BKH46cC1k4GUVMUvL6uwpIMfl1nhnT9BXMi+b3yaxg2UA0m0xuHhBrXwkmNqd99STaztv3bBfZcn
FBN0dgjtgnTd6FJCcGIphO7EPA3qi6guNdQbw4ujYNAk+Bw6QrLBcoHw8PxkiQ4OyF5acF+nsQc5
gC1olOhFHiYiXj0o47I6EOPzT22PlpqzSIzyYwt23NZeFxdantcImwj6TiXY5XM9niEdGn/2q8zl
FT048Xt5tcdG1ABB8DWxCXxmBaVRNw6f+TGwgJ2+YgrWgKTM96ALPW1xsoFnSc/6qsqjLbCwKJHV
1CAMS0Fbz8kZ8ZKLg/uNBEmYbp8iQddhEvtDPZTTHMG65O1RomV6R6G11nbgiucYi8muCN9I6zXa
H0gLtc9lAZ7XjUAAN3LT2eTgRmZRh+zUJiFNgkpBcWGCK0bGZ6ObIsUn2xsC/webCBUlfpC4TfWw
j3k4lezlhDO3RATJ8N5ObtQ5DsATLJfNBx62XBwU6eK1bQjnzOhlhdc26BKxgsNRk81FtEWm/3XF
SLZx51Jbzq+UEerUFkf/Pw+iUBBNPd8Dc7En//DFeiJVGiEZJH09rmoHlICwe6GaAwxYOrkwmqed
4pIWMrXctjLsb7kIAuCzS9xA6CBLEPE0vxBt+CU1lFOB/78CUtxycKIvGSYHzhxo/3OsIe/ioz9U
bQilCrXX+SSuAUGS5u7+rejf1QUD7o6WqlRbHo+lMnDURle8ssABVb9+k0knkn+eUhPNBf2aVhMs
qFrUrrPHdDgDFgIxa2HBOW8j1PSKr5CD9qAz8fC6dS1YzVmN52fxr1pIAAEslYSqZcpsLsUJpXu+
WEY9iQx2Y+9F65X0nRqJNU1xqHVm22lfGsEox19hiEFSIO4cfW46WAgtg2ASk5t8IG0GA5CsEt40
2r5P3ETtyqA/MZ97aTjvAO6HYUiO5E9Lx84KSCBn+FLtrpvfXrYNdUxc2fRaFWMAnaE/Oo2Vamhu
1t4JpXvkSSRyXxUdZZnxJfZqkrgJuW6tgeRzMpAPNkyB3BHbkJD6HFLXWDqlVuXY7aG7m0zR11+S
X57G9yMVms3oUedLG2CDnuBQoDxn2DHss0UZtZSkgNC891dYzUIvkMxlOoJF2j33Dh1HXvbKnrRx
jgCFVOIUt582d6RZ55IPaqs3kIprH/lZDKZurvEcGlxpr18JNqBBkRIGKzKWVaBBRMJc8fWCNgRS
/8FCFbyGwdYnRACjH3s0rGIkVtV6dSR7xGe1tTtDtwXy9WZaLKic72sHkRd4uPnzDhliu7IWidYX
z6M/hqoI62K1Of9nmfsNU3mY0xsj6jkHxdmEyoAgT878vneGrqKGQTk6O/rB7jv0cx2WuWM0Krrt
EaU1pQX3kvwY3JFLX5SObg3xrc50H6M/YMw7OLvBEuozW6wO15NJ3jyORL0ikLi4TBTOgWQhjUzG
pDiRdgH9HnUXRYEFc0NoG3Yr0YH9IR8pksoPGW9jS3KbYS81H1VctYXg+CdufrZNkurZEGT783DI
FxG8Ha06r1iIMiXgUfR9Jw8AL8+qZqFR1x0uA9uj2g02uPxlA8cXjxOLIX51zaQUqeE/C8OXYggy
THqYWK2u1AQndfp31JQ4oj6qNqmammulE+ZgobFy2uYD88OdDp+q47UmnwMqFEOTzHYaSOlTQM9P
wEou14rd0QO5hPY4pve6mrWGcdi1hgHm9o0MH+5a5kxW4ByzBMIKxJnyDQu7wYmRFR1+Bat9mZAl
OTCky0ViNbvxKFVg3yB5ZlzKeGg77rvp36T8atgcSb9acdyxdmD9yTrWS+CpxsTl//Dy/IVLjmKR
CF4m94HUmIQ1ZT9lJAfjZ9rX3USNpSPrH9Vm/s77Jj0DgBM1k+rW1AxiepoHoZKsCewxWQsYCWCG
6hwTP3S9hiQyKBZ6hz83h8tO90Dm1W8x1brLi3+Yc0ymSduc1oINZzyVzOsO8wGFHP3y7+GaerTw
xqKx7zw376lTz55iyCrFeldTCcCELu3cv4uEZB/6jrhd+y6oD9w0vbMlXbspJZI41jRd0eZ53oVv
3wVXV15AyySXbGZF3113Lod78RCI8EgMMCC2Usdo5QvrGMWnTfU6Wxf8HIg0tBZ8UshvGdp/KreS
pKVFF/OlUcsRv4BLUj5Lx0wMKd05qW6ICa1mhNKpfB7Fj6IfOXSHmdqJIZhOGA30yCOh4oq6pxrb
SYG3xGt7gDqx1mJkw64gXO4Lrrn2LMBUfujKgff9JzYtu/3GvA7c8ZS63hO6N8wM4NNcnryY33wc
LkV/ezTkpUr9ubZ/IHdbor6AV8jMk2rONzlKtmTiF7aLhxZO+i38xtX/RynZsQvPbE3ii5obIjJa
3kqw866FWHx7khfxxu3tN2Z8KNUN2twjrQSPHRm/D+Y+Yr7M4hpk2V3Xsh3gSlgUCF6lYEipy3ig
TDfuEpaZuQAMUa2LbHbGYmNnY/ymsZcZodAj+aUqFzrd1vhvahw9ScLwRdDDNgO0d7Kig7UQnVw/
gYITT5eKY3bG3ulwTQ4XfqB2ZHqU+vQx8KdqFJF6tPoiMOD/vqNOQC3T4n5ahQ53t9npCATcKfAo
5bNDwVU0MXJjayFAGKdrQjka2Q3j0uRrwgNh9fjILVldGPhK+N1lseZWKcRykrR+76X0ZqldyVli
8efz+fNyVXVf/IIx/yJwDJjfadfB59/Q3/CQuFt3WWA6yaUfkpMMFGm+S8dqKWlh+FMXGMOTWN0O
3gAg/iusKTdFVureer7Ja5XdlHTYv3+dy7sh7UXb81sIYv7f2wWgEudVJOhElFEd4LKxF9c88xvJ
+FqB9dhwvzLmAocTNCm+NAd3AIFSWo2YHuoG7pJrBDgAVhndQhh6orRTNLLrXcdL1PN0FkGDMoBy
P3zICYy/ATJ2u8jZISI4bZClFX8ukUyjIo1VoBPPx02N7juXHTxdDqFsrvjRl+74UX5/XCnE3rQd
gNH5hsfDX3w5LIGnxIcj72pAA5KiCdiY7FROLfQdEtr1fDbJjl9kg7OKN4ZbmaAKin38qSolEKjA
kTjzU2l2sUPdecxK8AJfaycBxYQ0CTzN4YGbagOag+ke3tD8lH61ZTzLo4S5TBwMNddyWqs20185
DOA4/b5YnCsa+4gru2d4XhipqKZDyC3qApWHCbJCXR5bpQfHGEIXPkgHhvFvBBhI7jkyEJgCE8UJ
4k9IotlvOoLi7yR2jUe1DzmTs7UuBZ/S6oY3mCkuQuBKltEVVDFbsuD04olk3SLimcR7tsDuM+yo
f8rLKt3Y6pgUuWmKNJIPx9b9ER+L9I3UHilQ9vLPKT+85M+Fqbqc5s48PiVsdq+RF8M6hlc5FeL/
UgBJ3vNZpnAYdKI6pKlP21VTRuzkMAfoV+Nvjee4mDSN7p24w4+VedFskdVzHfuz+B/IauSX3vXY
vWwhuO1J+jT32GrLOa+tsADrhugqQIfEBhggeGq05YntGr7PMgsdhwC2P1SH05oLm+K+JJNJdFBf
QGCDhxfYnEYW40nFaMj1hf4+lKMnYflvu1tBSVaw6yaYTPnwvD5ZKgsd3omT0CrXk3ovPafL/F0k
YooqSBvfPHw5/p7MVEXOfB0p5UzcYu3Oqgawhvy8/d8yGMw5LUcW/TprCewoUFSTrhvsfzwDf5df
pM1Z2h2+RcMaQ/eQTqhM8Ekt6qGB9e4J+XyH4Hoo+EZaCH6RXMv4GLYscU6u7971v9SRtEZIT714
jPpxfAd+n27jj2A30gDto/n1GrcQ3oJECycImeSE2soL/4fwae7INm6Z0GWkg7BaSr49FY3KxNm5
alfoT1OZm0m3Lz7hZ0GQIOOE5CwMOvlmmdoV0grlHWIEydGCRbb0crlWVXtwpdCKs4Dr43DuIdKm
7jqT878VgUoMQ7mYU3LmJ8R3fJpr1lZdnK8wDZJt9xdzHcdMPHGMQ5BxWe3QPq/4CyPbi7JQC6yG
R/U1GOZNANStdVYOKcI9za4MweY9rfFVHoRfxAaRahjeVCC4OBWRyvqdNJrJqj394OEdtE5E7Qjs
vq4O6SS7X8JJerXAkLQtKTRRiruPc3wkE4iKXSTwbIybEzM0FLBzMTyM+8w+elA7IOfyhTeUL3Q0
j02CdqSxp5AUn/PYx15hwv93PTB0abQGTqEBLz5bmyh4TxFDAYFRbP6wgH2g36Bv0tOBaP9B1nA4
OUrrrWtqSHwvtY7giyaHDK23ipmc6ZjN3fTAPC1SFx93RpTILWT4G4fNOa5xm+oE8XB4pXBa0zNT
J2jNW+e6b1FdTsAs9sJisV3s60Ve4L+7FkU27pZaSeZza1uqoPKhTAH41PHlk/TvxdT8SkpGAmkE
WXP3VvvTUrybS00xyTyppg28U0Z6Q9XjFa/sty6zx6tMpk6w+XrnVF3En3LZgdY61Mq6PDd9ENMS
GCXurD42WB3zcDr7J1xJSaubIYrNpQcV0JJcaKXKRlNUS+lYn8pqu2K9nqD3QDylOB1kU4ats4Jw
KgTqvmGYMHBLm0zKTUKK6zHrrGb0+HCIIr/S9Wr3vZaj3tmZ6vn7Gs3VmqGfwKbrf5NbpOqEYWUX
xSM+OsyUDLujYO4+VVjtQZ5TUIu+zVcRbQhAHAzR2nb5NQtPRhZFrjGtNtYpxWz3c/3xZpteFmR0
SexkEdYMtyZp9PIPpc5pn4sRnjq31DFCASm+oIC/RtcYEUoM022sR9h1bnAXW13zmUkI6zblMJRT
LofVN2D7+vFxbFODQak0UHkQDH3oNkixPV/9pAKOmMywKU7AXJW8jpan+4LRFZVhNNjSReNWGpOU
ELbDF07zARqGx0ncSMo+WoXC9bTOYDkUbrE73EqtC8kX6s6EQcY+ElERWcgZ0cksscvQBYuaQ+U4
o9mJjphuggouO4m4DFsFq4BS6VuJK6p+loYoZ87+p62s6fHw4PDz+QLFqiFFPeD2BMAw19i+hkSP
lAVSLKT9T6+YKoV+MJ4TFGbb47SpaTcZtMq6/UlnatmYQyiwv1G4TbrJedw92PH72zYXAivmUYfe
3HK81+juPBUjCX5aZdfJlFCvVAsX1jV2UFqwi9CL38nG1xbUS6xmEoK13+L4sviIDXPhecptjecc
t1nJ5hrZGv17FUQDpZSvP0pZGDbTH13P+ZS6R8mmrMPu+1Dw8wjB5d5m8nGR1AsNo0XDbn0CikTV
oOI4sXFTHq3YqgRo0Z5gbC9MAR7d9JRNCs6oaECW0NsO6MjwTy8AOxu/li398nSiw/0ZaRAIojvW
BpgIBB0Dwkf+MIjoy/0oFWtzOLab1NdsFf9VFzs0Tk9QSfH6OMH8ckux0zDDwy/ShrQW5SyDYe3Q
NQfEGvhLFytiHf8zaCLihRE6rLywMyUA8wbN1CJlyONpZOVz9rFrMyZpxKlq1XAYnUyGnghqf+qj
dW2gDTNetnRBbmJ/qYAM4OxU1DIoOJIKV/h63xRXFD2D3MuiQNk7osEcIMKEDMH7LlngXSBuwZ/c
CbHXqnHut/NMihoIx6yiESV5QZuYWXnBmWmlgcZpR6iNsUGGSAtI3REIpdshzflH0mDzF5YkvEhB
YSfcSl9hdpOfmaTe1d2N+ti46pPQ8a7EdKpo4Usp4/nqix7DuoumrHaEkxKx1eeyx66Mt0/7Ofsj
SUOzIAIndYrJ15HaiPiDnfuWeGbqT6E0Bo9pKYhqjIzrlX3iV+c31rycmDEk59elerX5r8+CneDh
uE5hpjtY5h5jjq7ux/PDXns1fhXjbx95ELNfTv6HZhH7vfXEKZtpMW/RabiswIpm4xTR6BmhJ+/W
x5cVk5WLyIadDLnzsyJmwmJRzgOQlrUhvETqBPHqUp6MvsfdmGEasOHK0zBk+k7hGjMGsN/GynXZ
ou+kY9q4u95v79IZCi8Ifcv3KRkIZb5iDF/+JJWIJCjV1ebH17D+RF7KqZhtv4lEYV9d3D4pw9Yn
Lw6Ie7fO7UnfjuJktEfyybx09oJxgEao/sWXbjIE6WE9OxwUpMgiI4t7kILTbBgVxhFsol85Edze
vNC7eSIjGvnZoiDNrgbv8kKSHVlb7lWH2MCl7vsed+Tz9lxt7QqIX5+I58rK7skh/lmv6QvIFFX1
RMbl5GcWnr3s3u5c2ucsyFcFPZclLl2mCB2oe8Mq+X/wQax4auCAoHx07fc4coeuYidRtry444tN
QeWSTNLnQWoEDFdZHtrxuv5fUeq8wd43Cl4ZospDXQqB8hRnje96h1G2vd8kvWNiEMFtSMQ9s+Qe
26g8NIYitIuiYS8yRLRx15n1XLMjt2E98JIpUN50nPZXsK4Pas1mbV4DsplWWBqw40c63d3nf+lD
MlTdiVvii6xAohvC75B16sU1L8Gt3as0nIXkuiJcnRFKRNjmFqRHdG0zojWbWHIqPkrB5qma9UuT
/2cdz5DXXzgfYYEbzEfJFx0emuk5Z6reUhzn4lhJEIEuzsyHZ3tUeuycLOSkuxyayL8+UIbGJgER
4FTvKciI24fYyXig/i1KAWGlyzaRSrcH3EanNotmVjPOzMM8D2tRZGJxLBNPeSaCuZlmfDqYYSgW
lsKxVGysADrzkDPfCHPYXyOZKMKWN5w0CpdyqUS4Is/gHKlaxNznnxSPcDbu4PNdD4l7TjPh+p2U
7X+FOmHd+xhR+wtQ8QUWf8IJiR6TZl3FxX4ivBHcnUFqg3ChfFsyoB1HDijzIYxJK8DxyUmEUAdZ
CjlkpLdcW0a+5kr44WIEq+sCSDks4y0hzCnHDYOuUZqyYNOOsI+ujN9p34HNmE43isGMpjiRIdYE
WPdLscvcLqrnqCWvHEEDs+hZ4H/JQU08iuB08KN40ipypHKyMFxdf6oLTQYGQXRvKNSOIxEZiLC7
jTALKj+mvijKqnFdoBDGIpXGwfXWuz7NorVvdNtxzw3JvIbJ48Zzgzl+bjJtx/gZDhHrpyJsabjF
wVXWtOoj2MIpiPrmkXD2lD07ohbF3LsRyynJHchz5X/if9JVF8UInFhE28yrEW5A6aNhMoeVhwmD
hrd9yY5P6aHkO8Gj+YEsl1SOtMfFYd60m1SoQX7gqrTqlBZErXlPdUNTG/1yPu9N/UE73YbS8Jg1
VuPDulX5pQ6iGmU9CjZt6sdwwkcxJKCYbZuKODtBl7a8k1LJkoz6Xk4bDY6W+EklANc2Di/r/FMB
Yjq164JygZCoqNVh+kCdE4jNG8wVWMvJfzYPDlgxoRNZV2L4me1Vtxvi/ODVfXsV0USzjQgrkazX
7fgAZCUk0njkIjtK5bbrKf5XnwhFEPpdimJXtFeyGvrx8BSq0+E10M+SGd12ExwF4xXTt+IfYFSb
kJSJGDoBgEXnY0rKAUE1YTIUv0kLOhizX+/i67IgHUE3plnCNng1PDFalzpT4LrvvGGyXEVWJILl
+YEOVRB52kRPGqglKHgronhF1BcL8CA+IMNO0jdoe3sx23p/squshpaa4lMfAwhYY3HHWG3224gb
ykPdmWYueww5mFor30hhqd+yMUYDwSZwTbgYTJ2DSJ/XqItEAG6I4J5M9QWxUmXDrepxk93F1BUD
x5W55Lz1sRAE1/GXpnWfM9Zxfd+6mGa2OlNiZ2U5fZ4c/BAanLLGo1Y3f+njTN05YDnTJ/G3gbXU
7UctLZ9cZw1BxXU7FDqU+eG286SrB0V/ZwTEgI3opQ/TNKyoSsaPqBcq6U9Q4F0MWKs7LukBAe2I
CqUt1GDkiTal+fiEW1293Uq+Gb9sLU3gcQeoGYgd18WsnNRWGRCfzsiIdGjDMSnO9/vP/nv3/VpW
hqAYGhxqE0+RNdPDyRKH2wkwAp0oU/JCRwT+l51perNvzyMF0Tlj/UYwnqU8HV6fCbDqm6PuTkfW
rH5SKI4YCNapy4Ov1GhpvQfYCsQH4ehEc7TOJlSVo/gBaC2SqW1nPCHrtCvWv+UR3hhfKn54JGDa
NTqhOlzptKXDShevDPmKLQ3fIPCZGThw/90yWf9H8ojOeeXJbSXjSR2IUA0jXcH9GwKWTxfjtl5p
wRP1aqYpIoeSxa+cVPuRJMf1yc2Rpz7/kW6jq1043W0xaU0tGIJOX3pYptOesCeBfT7hdlRGI7dy
ebyISeb4IrJlLrmGKrtuSGUXVSi7fGHNhHbf3NVHuM8a116PI4omruPFyI9n2i2Ymiq9RI/G5Lvm
BxlYqjWvDd9iXeF2dnQDTT6putrBDZiZ8LQbeO9C95NHHA/B+j+rgOamiVvgrlNsN87XLSkG7iws
tmhVsAw64gp4e3EdkH4tGR3Y6WD2AJztEm6Exl0kBmUNp0ugF4eQXW+oETQ9dGFrMz8hihyj5tba
JMYAFrlV+2h4yQQvtnucR7PzuweYvm7n2WmUhXj098C652JbLFZcuXqGs93aALvrXGZFBq6rUPmH
Ni1oTZJ6sY0S1Dp5EZM17G81AdpJe/WLtTVPxxvqshIuPShKAu4mZSugWiJiYIJMqQcCJrWtHw5c
ixwr9lxXs8QRSB8NJyrY5u6NuemufG1WNILHmnvIndK36hg+nYyrYptj3snuAVXqsGGej3G7EQvN
z8hSLPKmQtZDlsIRMirr76C8/ar3JxyMP2/Gyqoa87DlGg/R3JzpD+NSRDHWK5o/pO+tVNgVKFlA
/l/JijkaO0bHNcs6hA7spShfNj0YQ3pN6ZuPKuwFigzA8ScZ4gRKPbAXUdl9DPJA8TVMYPzfDSI/
Yo54T9V6jsIXUU5WwPWGTQmBIrxLD77OjVdlF+dfm6iZgGLssoPYPindBz6T5AOPdth5Y9hu5NX1
fOeeK0QMuaWzecNJcEQURcAZpd48OyFdrBWcUmFMceP5TGTK9h2q6BjteVjpRjHCPehxQWllBz5G
EMFyodt2DoFkf0yZmxhvLvbTOqGf8i16A65ARTh4MZ6gD39YXWx3a1CdlyoUN3XfqDG//3VdDt65
y1qRd21An7YAsNSGhnGgCWvFPPJsjivPizrXZnfvMM2dRmNnHsVX8a1Fx0ZMkKdFLtHpLV0pv4Z4
xhM0w3z9QLGJYXMwbgbFCsCQArIjExZ0fXE7ztcCTzZe6GswdAMPGLRAaFHpoqHCF+YRkI9WkMVV
SBwKLQIX1+B4G6aF4dmiRaXdK3LcvphqQPNmWL7eA73ihqT9EPMO+pOXClbfY8Se7yo/69b4oQ58
1HjLJW4BW7Y8yxezsyvUq586+y5FPDVLdt0yhg+052EPGmi8GXcek7tRMz5n1G2MYdDTNYZi+p5D
2qoALCvS3f8vIKluSjOKKeklTEuKKFYd38dB9l4jRF2myb59BRgo/B7K1ufh2bznoVWBVM0wbJfF
sMWKCV/7kjUrixc0MyCFPS0V/kOvbWXvv6ZdhTSjkGagRdtZAXBO3rp0QR0yMEDgWRI9G5l39bdk
KD0YRxtIksf62/3Z53i63EAxaqJtMmPqBSiwie2NmE2Ns86oPpwVGagvtvZEQuFPeP0AI72RfoQA
Jrdk2reyJ8vhnirD2tyouwoGSp3utfDSUuvBFNGh5CfasRjiPJl2mzS7F48n3+5E88XaA0ZrXgUS
2KZy1zAaaPnzuGsk8Wf080rdYOlrxeNpHT0CNmux/BhomeKwwwcjadsDcBTNQi4R5srkaqa+5Q+Q
gem2EfnSDw6B8po8rKUge/F4lye2S+oiy/JB4Hd26As8vA40el4wq/DEfNPjq7MHTlmo23knsQyG
WqxyVVEMRQ4YrylVr1ZC6nflK9jyKcbJstcJlEGrsO/coaWqyyXRgouV802Cf7qkMKPQcV/h5FhW
MFcHVJwQjzDXRBeMtzhcln+XdmsTLzVT01m9h3rZrKZNSWKyOK/plv1cNu/OSfG41L5sS9n5cgF6
HxLoJbsR0gR9M759GWVNJ/2vjbQqV1vPV+Tx6cpxq6YIO9qpVKKzdXXzZPnb8JgWZ9Z870QCJngK
ypyWkWCH5IdorJeC+LqV96yTDsxJG1Ylm1u7sel0O3tJeBcpXdmzPkQ5O4D80NMrZlUB8pHi2JgO
ZV8anC+c5FUAwqmS/Qp+N7ZeoHTf2sMooPGDlaLtUmjIixnpuHt6T69F8R9ychenL3vTPFTKDEbc
dDfhuRjZ/gsZAo8sNKrRjANXwQ652/w5N8+0jzHxgrs8jZku2OD42st5pQeMetGf8j7DfE73ZPoV
Aa9xIP3m4doxlVdNC0qXk4ltlH3+zx/fNU/CpOiUTORejfHXqzH0K4egdASxGg4dssjvHeUsoL6s
6faT9o/QYBS84Q1U0xFGLcFEkHzPJ4bGQhIw05FH4k/dMbH/XM1suMPFeTANXM+Iuj9Hl2u/lNYU
B8DpbY3/EVO7Ecw5UONYZK0NFujpptPgWWRSdMRf/d1Qmu49O7l8FwzcCHIB41zO3ftAC0KZqc8A
borQ41J7Sy20OVHnnAMWnsAg3KUIEUoPH1/Fa7zSACfqTF67jvtck4tis5nKSrXGlv+WbAnoumSm
I4rZSuuWmSws9Bk9mVqqHTqUpTwtC4NRJHH0zLQcQkgHEI/2+zV1ksG1M2OxaReeRjmiY+UClzVO
v/TazABU7hIcsN1yIJ5HvCtGJr98KEgXQEngY7i4ABss8WSdEyGRAYS7IOgtXG/CzVfuIwHQLMCH
B0OiSdsLqSkJ7hAHMsM83AQ2+Cf6sTFjWXO2Hx347ta80Qw5D1Kzzs9EBPo3/FAadBkMpto9Trsr
xxdqRspI6+QrpAF7NejAa42eJWj30PGiJzJ9MmoY0MZ3AAFx4J+J8n5UBZik+6FXrtwgh79hLop1
Ed8ql6ZRlRs+XK/iP2sQI77SptDIc+4eTE15bc6kogFPlG9XD+DPMR9jfZcUbS4MCa6aFyOjbZqp
T8gesYLRqGxe9KY7oXucyPpBktNKFsKrfuZuIVQm4tldFiiIYp1jsyFpb4wpOEehpYuLz8Ea0BHm
Aqac4kcA67OaAdLlhAvr/RXBKQ/868AhqWooaiqsnI8C4o07e4FcJhAI6zXfofvDMj2TqhYxAHDY
h/9blnveWfuPG/MjHxwRliP6B3YFq3FT8tBlULN16PvSFl+lp2PEj36DP5k5+G+RUyH1GVw2dFZc
5M9tPf6Z3DmbiLu19Qs7Pa14cxeUySNhuKHDH2zcWKFwhr1lp9F6v8xm/+2sMmg08qlV71Tx2BRh
VdtU2DxE3vczXOoA1z0plC3/J0KAi8ZH9SF8LTKfahOqPSbSZS6NguZ5/8QySkHMgVqTCdQb5/tM
tmRKKZjsfN1UodsGObZkppux6lcKW1TUIoRdOEE1/VWSE0H7kM/w1f5qCgqpYgkUjhoZQ2MBo8bT
8gj/Xxpi/GtWN9T/2RqhkMlcMJI3gJI5f+66pgpNLsdgtTWGIg0vbOioM/XqGU7pPP1VBqgvq59G
kB5n/OBBBXmSnz6ssMoYP0SXpSDOmfm3v9kR1fhlpmZ9V1GVUwkaGeFm4AL83QISrjiN0RBDllgf
TEBXSS3VZJd/cguFqJCXVJIS4sBoIvyhJMcTgtT7GK5xeyJ2IklFECbSkFbMdCWMBI/XxDAOqHdV
GMSbaarLH0ukBRJ4WhiFB2LxF19vLgKwyveUbrkLRBsciDQ1zVnV6676okWbfBhjv8yRSvJivsbu
g6UWmUdNvGi82BtKHaf0zHPbxWDy4M+PfWarwW4kFy23Xkxkcgz/IEl75AtDKZOCmJTA9fbuhK0D
7ir9+XSHBcw9XXHwInm0r0ScMWYAV1lFJfSg7BFXfnhPqtVSooTroh9g8IYDtoSO3fpvkF754DJl
p+N8RV0hN020zltjLt54yBXK4FXT3qrQDFdtESrh8gjY9MTVz+sLJevtuMoA7ycinfSiNx0TZ+Ym
xPyJnHLirL5oZwtDICn0ZvVoaqMvj2CqcgBsTKmbYPePTO0XNLuqzy6vkMuMpQNm5jxUbGuNQ6Yu
+hrQVcee4Cc2CllHky73fQ8AxLnduyYpMD52R0l2oG6RcQjKNS4OAWHeLJFUoPKhoom3EbXzMI2Y
I8XAZ/EiBxrJYTnSvty2CdHdukXAVSLgodPWGcDcI/E2THZfLJAIHsMUKWJSga5hzsf1tFk23ctS
8d1ERXcChTuVXl9+K+hGVaeijudSmUz6tzc2jXTuXKgE2s9lYuDXwdo2TXxva6HxrtpzIN8cVRVK
qZMrVXukNl9xr4cjTdO8mQia9LLWJwHSNkfZi3iMZQpSu6HqlWfFd6Zc4nPEiapPSMP3pw4+86po
kF7muBf1dvNZ6J6CdGMuzYT7c3RUxkD69ZM3luPxUBQ4mjlL8fAQao/HF7qLjOurmyrUBnfl5xiz
rbEdIW0bW75WRFOcECfFJ6YlrOfedEYwv/9K0icO3QTqUshzjz7iAJ3WS6FfYzoxQC53hzXi87OT
7wCNsEkyhcpDCk9O/+AvJGzNQLzqPOwkQzK0LLooTc1rDaHQglynfHLMDdUr7u/pn1Lq6d/jUKh7
3gkYN5bwDcn30aqN46qX87+fjQ9bqs86qYJ194/yrONqU6W6k4rxF9jril+I5qLUNGSC+qEy14NU
3UnlWyIqyZpnC6d1vBUACkqd7eFi3wNj1RZSHHErhzrBnNOgxmPfjoK/+AP2BH7dseBV9m3eicte
0dNijxU3SPI25QJoJDZJzH+G2LuOWuTVvGWUvOhe24mLulqQI++eqs/vQzxIi0iNcAU/d45m9wVC
xk5kp3EGDsk39XQCK9XcoPx+gPGdASK3StSdE8MMz7levXYN1KrqGEYXtp9DRdVemQdMWFHy8QLx
rNiKsbaH0kZ6HSSPIKQUtTo9nH2sCorVXASdBiL9u5w5ZRfL/rX2Jw//r+gLK+yULkhZpY/R0xg4
8K8xPlWy61ek67NHU4/Vu4OeTqvcqfG4Ck6hDuMUD+lRpS6rpnrcFYafU/yIVeqaGLfYpIdZqLuw
72z/j3aJPeJ+OUTYVZp80MKoG/2Cqcev0mTH7zNHLRVawpmXyP1pqgg0mGGmioD52JvDdV4ucbvs
rWFhYnv8WBce2WRoT673DegEt5mCVX12cNv81nylGBh92Va8CkCHyIecu7kXFMp9QLJe6mHkcBXc
9OMFQhm4DSuz1AI1tWC2oP9OdCPI1zDHHlRKuitPAU+qlUt+GWqPoTnGuw4/0ZzCkKoN8EJkxJSm
RWyNk9Q2SnJks1iO08KsyUqq2kHnVEe63nincObQ8yXlcAO54s/84xyRw4BuFpRkINK9JJS2+mKT
WC4UIY006YM5mWGkhsDXHxRgJiSmW3ApfBeNwa5TSQmhAlCY3Bcl5+b+/CIpZJ8XO3G5KghvFndM
/ak0Iny/QwHrK9686kHk2wDvwgH7JaFD3CbUjor5H5TnE55WmU7Ut6VCoKYbxv92mXyRWwG5SSvw
t90Etu91inmUMZLk+3vVb84t0bTrVxOO8ZVGSD41aXZn2KRhtCXU06qpFpBHrpdqxIJSaXvXtywK
6n2Dfm+REM16UXQRi7nqOKvFiNyJNMb6FhIcgegJw13jZmv3Myuk2oyn1iEfQsn/y0URIfMj6Q1V
GEt1AQkGx4EOkTu5tDyFajKexlY1jP5L6a7MXgVosRYAh2oJDy/Nfzd/uYV9pd7k7oVhv9wWwQvB
x51NaUyiu5teu0W6Xm2akKitn+vDqKsLz+prsvQdiZaHK6O4yp4S7VMI3S5dGGq0XCOAtzgNLci2
7ATRaTtIXUI3y+kAHas1imKlTZyS0cXRYLlZ3St7mxsay3SLyXi3LeSylDv6hsUchVaFX2ASTkUm
sRvcJfagbggOZ5e4UwMlKXy6vQg/pE1hJZ5VwniytM+mOIltyU+XGmfmpVIcmqhH2ssv/NMa/EkX
jOJCqfF0uQa2hqf5/2nAJ9wzT+eEToVw7QPqUicTr+E+s9wPSWYWURhmvaJiv72HnRuNa7rBG6yu
ycF+7YoOxGz4N3y9q8TEgmFym46VKULvxEaE44kgrQ2mlHfoMNBUpfHJyx0yKkGh8FC4A/eH7TBL
a7+LZyjum28br5lAtWPEF8k846rhPbkFs3nW2ArW0WSbRe62PCcc5fYP7uDEq5kUs2Qz6Y3G/fR2
jaZmGFCvqcihwBLKdWJkq0b9gyazQ3t51cH0XZ35BwsWpBM6qXG27PakuPeHUfJbZ2X5Fb9jaiw8
vOPFAHMrgYBgQDwtjpHLzAaP8vm/5ou57qP4+bHr+Mf53brCVSTS+7a3A87Xs+kNIygms+ArPjOM
PXgNvd+qrnv84QHDc26On57i59hPWZQD+C0UZaWCZhuYmHC6upUJVxYba/DCuAa/iApKb81mLq97
2yUI+ZC6x+obnH0TDzypSuw5BTl2JxirAe2IqPQqHxnHwK6ov3rSgNjTay7Di0P0gWFEr+1RNp62
1sF/9iLCe/JjAIX7tRwfAuSLrN/zaGkNx/W8mDmJhCW7NOSGvTjZil1Mc0l19UbpaF8sBKdAbiZ6
G8rhSH5IARK4X1e75PdKPXVK7HL6zMOwDQtcSeWuSnLjTs5A34MvtqKcB01yQMlDB5cjDmr3KsMw
xtP9qsxcqipxM78zbbzGgKtN9pmXnh51aKt1qg3lc2NUD6n0KfZ9fz0gL0H1VCTj3FiIJ3gJfSKL
0PanXSyhPhGZ/t4BklFFjjGtxn6ot7Zpg68rVSGSw9B2gRWbl1BaGimT1bUNfNs/Jmxa7YMI/Xc2
VIsltw8gp653r3UJarzdt6FwiygYLslajz2iQkhWcuntUlAKgfyEaw6zmiKRI+NwN4Gq0Z/ME1VC
3UbeHseWpQWOaBzZ+/aTd9nzxdy6Fm67wZiyJXPGK8snStLHdX0TPuKxEQ2h8WARPsR3AaT7XFsg
WKZJds249n/Bl1Y3dwZAZ5hR4S29uIyLtk9XEM8TFZBO5+L6sx7wQrA90ZcnZbwOeEOXVKvExB+Z
VuYUYOwFX3cwaubuMJq3QWVN1AhdNtRrPM9kxU2FFp08P3F8gLJhzEzE2RmmVHW5IVfa1RRd4xjt
QcbFpdjBvsYVZbvC/dYCHjphnCZQJAl8aDJ40CI2bCFOJY7/eIjF/aUvn72c+PX4KW8HBlAQUZN6
l6zhNNL3rdJ/3mZxC2dtAIYzyjBoNTjnc/h0tCVuLwiN/0ae1t6uefoC79I8vcz9AT2E/3ETqAq7
mTGJT5xKT7lWFXTtamQbv9T+5zIY2Ysiy2I25lisUo423prhHnCK2zZuHWElpOI0XSu1UMajluVl
c/rL9tUPpwyOvqvmqlLC4Hltg9xiyBXgTcbYL7Ez9O2U4bv/TblGIfJFfAa6c+dHOoAa5YOLeuRh
mLSZlvIKSZKSrIeP2VAeL7l6C/l7YycoNk8lN/p7zAIRVMD3NRFx0y/I8D/KUVrWO3KQh0PVtHle
66UwX6YvDc9D4KydkiGVWUMNVaMwcmrurFLuh1Hpw/YGqc8WkbLKsrvcUNjWyyHu6Q50TxYRODMf
PDA8gEjJkm4jjNKwGukB+swQVeciimAy1vrID2zOgMuq33MXgapkYSysMZGFFh+em28U1HkusYNf
o6NV6AjKq7NtUqALrH1b/w5pGsKk9kTPwc+nlNrUWrp1ow67ebz1mJ9wN6Wkf97q9BU+qxIbt67H
QcVCTNgdq1bWrfOwArCMRUJWQiKDCSF0OxBoK7igaBKAyg8F5v9e52xZOjYNKnoHaP2VSiNLFhrX
JYfIYBXhBvhnnVutM65Gw0PR8HksPhgiIN9hzidkFl6R8vMfUGqvga6+85t07rk2Mb7lB6jz1a8h
nDwZwTu++a9uARyfcdoCU6q+R1tjgzXQpH4Qq+bhjyCyG+vWspgFEclH6TU0IdZ5MSBV1N47Z9kT
OJIqkfXBD+r0ccUSduuyMdmFrpgykSHPSYSPbGHNV4ftYIBYcbAnAVCy9p87NuVGZ7MGPAh6eFo/
gofCiUaMKwyw/hLQYN83gvf3dU5GXodOl34V0G07ldKrgau1o/RovgOrOb+FdbHCs7ydQ6tox/8c
85QuWRsG2taIfo+6wtYV+0qPjziXnrkxc0sGQlDKeYkFt2x0iTj6SB7riccemamYbezub6LASJP6
706blLkqMhYMnP6q+5NCevK3TVshIplsrQYJsCi22Rf46taVWTU1g0Wpq1Uq/dIYGgrwWst9ci41
pilSU6xKg5HmSP6z3gowQBRWTKStXXfNdHwBXz60MFEYqEgV4L3EBSalQ1jLfS4GZJvgvSCw6Gic
bSi6pZadlpDLqq0dmrDKZiJLs2h1YLtjkmXOIKD64K/bcaQoKGss0LAKZD0H9fXkZyXuwNQ9MbNN
b3kCfL2zCm8qXVWbQOxw2DT8JhKB+C9gJJBtE0ikUUNef0I2FxsfgMzfNHvVIqWLM1Srblz/bpxa
ldKzohohPZPJas+g32R5tekvBP/r1ZdviXw5zyCConk9tOquiongF+9mi9mBvBJZCgIucAEJbWwt
asRRudgoYaE6RugeyF1ArZGqOxOxrJWJVyUDXCbRadbxlYABxzUXev9yd1gJGxmwS6pO+HrUAgrl
Sue7oBm3bSdXfnNFnYkZtZh0vhb7m7lQYexqjuQlsbZ10UWOy6GMDIqnYWDB79vCgnhpo00PJ+1O
y7S2f/XtoJyY9OJ0VJWUxTjZg/i4+thZHqA8qEwrYF0lHkYjxh54YC2BpzXNK0+GeYf0DMNQRi5K
0k2SoNLRMtYv75JMEjHhlDfRMz8CYN1QpkkG34GFoeesdBQ88/Gm/nJwwZL36S1p+Ht/KQJY4BLy
bncs/Cv58zHAdYL8qJcHWwMqgMd0HU3sWZEvjZKEMSVeMkj5AL7uKFCBFsyI4nLeDp0WG+ibJtWh
Bu5f6gbQubK33qKyMuFx3UOSmVbT7MNjzP1gDV/h9QYHioWhcFX/bWcR5gas2p3OKuaSZHGYgKfi
PK6qXQmdjVXWnQybps2WMnsVwmVOU9+P8NKQCmVS/+xBz3r/jdqZWLpUba+OzJ1I3RLrvVxN2OdI
5sPCplSG8Ye5zan+SrRkhgl99+V4tXHyroYv5IqKahmkE2ldA/5HjFwnJak/sTa6JvXYs/T6+XVs
j5inBC7JH+DRXRaL9zFTlzn3qSos2uJ/uKtqrHGxP5dogtyBcEOgefcoXlWbpPk5iNF4tlD9JaO7
Z3sBbmxsrxuxa0I1enz4LK1cBavU1oLUfF77KCLlID4Wz5+qxDwP3mlzQK4bz9xFkYUOY+S9X7xw
2y/mb9GrkwDdd4i3/yBxCdIKyBFqkW1TPy6kOP7fX6WK2+8mmDYioE2GWXpklL3U6/ZmTGKm5dIg
tdo5gJRI8+wWvkoBlQMvzARRHNGZHFYfbQTD0/dGJTeh3vTk3qugU0WvKf0gfwVKXk3I0BWEq1ae
0z45+KiIHoZItZmlX1cgMCxLSbMs5y6MfK5L+TTo/H+GXX8a/xWZN+ciGGCH2fFzG3Cf32Ujrii5
HFr9enPUoDQMTKzrYaC3hUlNTq2lNE6X85xMcOqFV3O8zGm0Xfvm6FPSOtXVI8/WKE3PQ15GaKBx
zQMvUCnSsaa4gniy/4oHDGKAco0NTMqBoazYGWMIG+IQs7fvVZRI4bVXow/TxLHQDXXtT6Xy2L2F
UL5wiNWTPMId3UcDitURLk3KJjqDPR6RpuGFEy5Wh+O9Ot2DTYGfZPvDU17cMllsPov0ZvxELD44
avOZ6HbZZBcRtM7Z3besnFn5nnet+NRpjeuCJ0Pf+idV/+uJ+d9tQ6IFfuWyoZZEDnqZdBu8913b
oyqKvdP+eOdCKKQigfUJAhsPc6yrR5VJssdShzMs6CVBZYCJrasyrUYR1NKpTTyBREy8EWtI4ybK
ZFIKKfLhcajqDNQ7k4yH55XRqKyFLna8MTb6bfHBwmp8+/aiwfFA714YpgsK23Td5eAgXq5QRI1P
P8t++x3v7tduuDhXqt/THw+rc2YbY0xhK41XhHpJvk8jXbGzYmhtkwPqW4qEbN080BZXifKLH1bi
GLfhChYDxKdzjVU9/APuQ3wipeHsEAASKd8Bzkt6IucGmY012yKnX9py2sPHBgnUY5WaVnYVePpB
RT2jYnQ1xN27DPnGOYpvBu+XTLk3qMmYBySgcRkWpWE4YSPGowP1xDLdf1lkjYoFI5Q5iphrd2HD
mmai0f+ZaLCSmVZUqtsbMQn5DKIm1ZTm/986GSMqu8Qv0UvHl1k4QoLaWxqSZ4ZzL5J/CFyX4RJz
EETk/kP4Dt1pIqGx7Djx8GJuFdDIhAgjZEyqGRKGHGn6jO++i1fqg3oWQPNCmcoH6lt44WgAfhbl
4zmHk8BTMl8t7F7Wb7bjkI9RKPGHQiBYWfLFiX+8joJh4kpHFo4z3/1/OiKBPcP0TiPTWZaaSSEb
8wnUD2fMa9O9I1ofEjqKFLM/mLEWTOBFStVQ11zj/c5W9pLMqoqrrjnLdP4+q+c90GprAmaDFE+g
/OVNTiSvd1qV76X8ySelO2IpbswqQOJrjIt8R5q5oZSaWTLRlH2YoFmTdcaTXPqA8MZp1FKZ9XlC
MxGBpWZq0jS0TmZqsZwxkU1HO908GPSdMkIBa1d1Cl8Neg437yJw4o9dSIj0NRVZqbPEKNgOcq47
8YqIUaBJ53LsfCfGJ/FZ8WJT6p4eaucB4e0w89zs7LWJ919vh9ZB/DfVe54uz/Kto6mEy8xRwiib
Qa5gRiB9XBJMcPAMn8b3jDfzevGaHyqfEiM74JzxTAucpQwSlI3uXUYhUcXTJes0rQuS1nsXJYGX
XcpxuWbTG5QTx/4RxBUKTKGBdJ0VNvfsApJLKLB/zdHBsntzl87/r5F00qy2DR5x/QVr71HwpGpY
GZiL/ntc7p/VZbLvSnkZiKV/wyT66O5FbvHqf31aWq9Cu0fPzNvfAJb3HIdpKU2wRLYISPvpx0MH
kiET2V4lMBTC9GIYIEK3hGbrYn8qzjGCnUPPG/7A2sdwlApaE6ijt8lxb/KYOUgdcCSLITHkRUZS
hLo/9P25UWs1J4NJKK2ELpf+7wdiDOwprKH7FkMx7GgxSfGRptz2QK+gRKScoGeNGB/WKg5pRRCO
RaBNqqHuz6WbIVRuynpdyn+PQJGkKfHrmFamrEcxRIUPKqE7CB7qz62gWwigyXOICwypaRupHCNI
rLNEkJkW86ebbd3PAKTRe2XGmZ4QMYhL2rjK1FHbzghfqxXPj+cxYBGuodclRzJfS90q73b5oZI+
KRj3sviyiWvErPgdZFlyh7qeMYUyDdqndbgj43hEEs8xJOrQe8vnPgE9QQwk+KOeys5baj3+obft
JzUJ7nGer/mIgf/P/wx7jE8MlS/FViG/C/qZ76QKG00VV1Ej/I7Le5oHVoDgDnCOkoqHBsxRZ799
pUGcb0I8SfhWwodZnsbDKogLW7b1bn2Iw9YqIen9RleiVw6TaX99OOoXqtuQNpY3pZVQ/vmU3msN
paOrszPvIyuHAo7XU7oCkJD+6XhJd+689ZwBz2WYE/5Mywu9qsK80KsJTexAshLju3h+OrFledb3
djIwK3wag+v4CKhXal4mDDK8imJyHrrdbvyPWzlIkd9oQb2nUKveRyNC5V/7YTTMqltzwVNdmFMl
vvpFmGd1wU/KufPCY5/K/Z7Tx39CRnoFZ9iJes6UDbchIO78SNDM6cabBxvTNkB2631PgWgf8nC/
QbpGJo0mX6z2G/KfHjCwPIuGSc3+PpMOh/dyFTTtAGG6DZYr3gUlj2Bj1+7hD0T0HVvcgcfaKz4F
lbmgnwTl7F9f7Q9hZ1dUf8zPhhpWJK+Yo7TWuNeLVhIo1r8OewGO3Gf6eUxQrx4q4ahABHGLgsCO
JuhSgsd4kYkutA+EgTiBSbE1riIJL9ULgDn2vUbVt4VAhS2y5HL2oqmUgTFzol1/n4uBsdNctFke
oAONRXjlJvObAuW5rpI8e6P259Kcx0A5FnTjROkd53ni5mRQXwXu6vIXAiRgpAIG3bjrK+d0uRxb
nVLi52PImF1aY3gF/Y2PNwaLoWbNik7KDdg1AifrZ6CNSGwIoYmplJvaqGbtnGzSp8LoBLZWt0pd
3FSSo3O2tTuukd8aOp+UFe9M57hrQOisdUCvHqJexod1g97tco1yolKGn03TN+/D/W9PDkucrhxz
W86NEQQFj2L3HPvHwF7iZmV901A4wvz+RQZOt8Bt751TtcsDSC6Xv3a6vAl+i5fGpWZIKPaVhH+O
CuZkyLoNwU2vvqiaVKNuYM9xL4mdJc9Jm1CPzettUHl0UXPS8zCmEWBsDQL6mlLLf7ThhsFLKYyo
7UaAtPgL5VXoCK0EJ/TJg7vyQ+5AefMYXGX963KaSZNjT7o4m6V4xyKEjLGs0reqye8NKpeYOj+C
D/Zf5sDxgn+WRN3SPPM4krlXcHsYjXTD7h8MKkY7iH4hUqLUgnRDBSem6idKWIoqC4VcooyYn5Bq
s5euqa3/Lfy6QqjfGTljflKjK+7Y+ntmVXRtW/4SssolyOZYvcS0AZqwN+0nguWiUHYw/mlKUiSS
TD06s2EvhwK7IAK366xW2RzwGNUL3xG5lV65vL5yp/jAQZEPazO4R5mb74OUxk9+07vUWs7ODbea
Ri+UB8VfTYXOJcZZuwJY9+uKBBSS6Wdfo7n9zPDuhHBi/V1CTpE3k2XKDqoEpWbBcl2FmzDGzSUC
BSWXsoWz3H9nd7wN5wMTiEC/RGsXMZ96e7MPI7ja+dNZVG4kD3zDReL7e4qTr7mnyPAf0Nb0xxk8
j6Hfk1zYPVZq+J0OGf0DWnfR+vMmiJjHlqgtMP8o36iw2crQv6etZtiNx3Q0SSZ5n6zWBrj93bmy
+TySYtYLK3EKF+R6yr+IIfs7BgiMi9JfNrCNdV97pJM3vUl+Alx/FK9cPYmxvv5o7oR3/+n6ULIf
WsV4RGEu9Zfhfq2M2M40EHeBx8U0NtfoW7sXZiPWilugnnhHahChvuejv6OTBh1qUNid58eaC9Us
bOsAOvaSN2gEyH8gpFxcrFMDgqQRMXXNNVMYclYrRJ0E9eUXx10VeGw9H7zE8wyxUpV1J6lfBkzD
elRU0SGNOMkZmxWZWAaKQn3xjZiZP2d4fFG4rTcYYHVG++C8PYElcm533AFz7g6UC+FLjvMjfG6F
SXTLNue9As2Fucdfjn0apW96zWILFIARGRgaUKrJIrzVUH2uyhVARSdYHnCAyrkk40Wk8p01NBCk
W6QrmEfmncyqUt+IHIX66WFnfkd88i/PRkeuRls0r9qqi35UDjBnItFF9quduaoe4ae+58z7MQQv
qqFLP3Ag6k8GcuHXHwt8166b+1onjpAe2O6ZhOGQ5pmyUZZyY2ixBDHzSxwwqwCBp27j80E6dm9Q
rS3FW6Olk0vvOrEFfMEAAOi3J64EP+OIZ8rJk9n0n5JoL/q09RSn6VWt9HHdEfhyN0hBvinBgWDa
wn4u/tadHPK7ZlUgZBxWqHtEMS/K1z4ZGIUG3kSqz1BVR/TcVJ+r/nXdssZndJX5kPz5CfxjMeTs
f84yUa9hxZROp7NdYjfb21amvh9L/phyinHXWCRS58DDxjFKM0nQpipkLPS4+iCFP/hXOFpior0o
zkrmg69JWatE/I7fmZnMIgItzHCeBmg/80S5KR+eoo0eEMEDNh0NVRnC5VwHHaskM+pFyqB5pzLJ
Rb8CgeeV0948V3CPHvloXa+o1EqYJT90fg4pmeLvl7qQ8nCZlSpxnP4TUiKesqQY8zSJlq42v6CL
VTgStRtr1VNTPRnMqiev+sSodfTiwcBiHhjJO7pKFVhHZuVbvjlNWQRLJiV6vU6/fxhQGT031HjJ
JhKbxurwPmcgZ+k1izHrPImxNjioOR6CF7lQLeCS0ce+WU8Zw6tRPEPU5Rrvig993/NveDVsNXNK
Cc817m9iPf/59V5ML/Jm5Z2JGugAFhD4fdAI6/67XY1Jgp90h4MCsWssmymQsLhRpKomJihfavcy
DL4gDScTH8C1XBEHLSDmwR0OcxQdGMOzMX3vyA6TruW9h23eB1bz6a7TUFkYz+K2xMEDjWXiVHGF
NZJZbax24+6p4CCVVVv407zjPP2m34MyFQFbbrVOUrSeMBIz+lr1rgVuR5LB7NVv3wKwpRzV/Pd1
xoimz48r1FBaIOx1nn3kY2IkFLFSCTXWBlEnGPDRZf9qGxn1pWBpgK93ZzU/no2pmYjp4YWNZ93y
hD8v7dq7uzsakHKo1mJZibAt2tnjJdbMnx9vJ0PircsFJe5jypnBLc74r+a38mlt9hD4I5O4GWCd
rVp4nYoqIAmcCoea7tvqPj9l2PG8KzC6aG/NWu8M3QbylVQhnJUbirncTQTwCnvfGfv6UOBuWhSN
sF5h22d7ZsTEb+jYWlnMAY/jOJVf3seksypg/rbNDNkr8YozuAHYL0oVRqKwGzSFNfNyoB9e4HGa
6o6tGvz82JV2PCef+dOCKmguMEz7LZqDqbq3VVwWIowsC+rOQcVuPTcQeAJKX45lNQyQwIxnFbuq
9Ck/B+TTHMw+ktP1d3OhXfBExXtSS00U56YxErOX9Jh+mrnTvVmyTUEvzlulzeVl7DsFfLb78xZr
0iLRu2TrxJsaFKyQgRy4n9KQQOTEsq0o8PS8YNKfWkMKw1FSrqZcFQquiME0nh5uNkN3ztFUXfvU
mow4DG3fplfa3rDxGkZRRTZ/4x8EISr5ReY+f/gn/7DTvKy872mJZS+ob8K8IAEoyinGMqLrX2pH
D9b7SXMZktBqErwBeYKj4XHehO6vG1hctjl4Mm9Qb2z1h5NY0c2AyZm55oMjplIpPUEQFRExZDH9
i05Gb/mYYJMhkBUSQhSF19HpjUC8nbPcpHCoCAaRlUGUpvM0/hCEn6jq3K0elUq5s60YrL9LntUD
TJlDeyGJyxC6rPP4Lk+a0CobirGlkxlW3CQ7mIN0bJzGC0MxmiiXO4nwZ/Z2InkjSbw146vZBaKP
UtW/nMq9KbybMIn7icpzlQqHVOJeaqsx6kgatQC6N1rwCEU87p3EXNojqZaKhzPLugGtv8U/1boX
A6ZB/IPIatxcQnEFgsLoNNs8oidGHbBh5Y6tA5lRgEVLNJyjDVOUvucen81Hv86EbQ4OUx1QGSFJ
JJtcpMah6tJx6wNdl6sI3pNtbGuLxsvj5QFYhGdx3APwJWqdh0vsH8wZtQZMnwyLN9XJAvgeV9iB
vwxfOeAJYxK68O4aKYZ+mx1mrU0H+MyHbseCpPSl5HuTJRekXcUGjYRCGrsa0VW4/6+aWnHhMTXY
DfxqCkW3zQZeqINEHQrpGQuBQ79lJP9/RmFGcjKIWLlg6taxfMh/X2VVlyduBT9RFv61vDDcaS0l
fZ9ADstlX687f2M9yv8xyNiCrftsTw+4gRuyXz6jM/pBKZwEwr4/tXiQmlzrWRFqLX4Fx/04koec
XZF3Kq28m51zqmIHfav7AtpbY+OYOhLKSa3+F5gVjiAl6cgPkKzSIghpZEUNlARzrif5K5k/lPoJ
WWU4TLpkSjQnnVADrv36TgFAPEX+UbLNwzz6fdXDRIWzFjzyS3mXs42qeTdT1+0ZqT9wc1jOmr3l
C7zNDTjcBTgQimuAGsL8HpY7cEcR3eGTd+kCNPfojx8MqccUcVjcu1RR6DGDKXcDDK364HEqTE7V
J2v2RylTM2ZGoCuUdfeT0v2UUpxnYf5gWS0qfp1nwSgYZH5LHH3JNkf0DkScOR27tZT4XKbZA5BC
Xct6YSlgFllCzmYJ48JAQIm94trItdzmgbySpkFd1YLXlftvtwjDvYN2k/wwDmQZ6+HZTeZeDLwe
yVkfBPlPT+9U8PiGOExTe1ZUoPGzi7CzlG3a5xI0Qc1OMFvTXQBY8jqLPBmasLj94c0snkKk1iyT
3Jbj7Y3pQ6MI9XwbVF+1vzk/YPBZsqSdltv0BF2lfr1maebaX7gwbD1zUg0E/dT1pWZcNmUhY3G9
p1HGKlhM2DBk8iILu83uxTFBDXyux7FlnSqszqkcfrL/8ncL0FqTH3ZvMwpGdcW65zKCJhKKLslb
6VSy+3nC2N2VMhpoZYtBPMLCjQ6C9lB9ezqqgzGgPf+EJWjVpWxm5IXgwgynNN69YXJHnFXNDOR8
u0LUxURK1gTFoEUNN5qaActy3JVsPCC/QXkTiytkKdE7sISrxfdWZ17+cP7iQVJSQgKfsDcrMxpb
u8vdEgF/6DGjvzGn77WqeUAJP5DcJecYLhz157We25qQ/t0u7W2/+ATJwACHpUsKlcAhVuhoiTrW
ZR15oZmC6nNs8/dm6ugUPRlMvdnmpWMXYuvxDKUa6M0ubASLgmDivsNbyy4meguURFB78XDf3gSG
1EtTLxZz5n+Q/zIfCZ+oSeTXeExDXBDYyxmgo7T8/yVKOlSIT7Pt8j943p1tZGKkmMlmyM0JfSlb
V2ecoqTv+F0SREFe/SObRv1NwA3KHHjMCur8NLse9mzY169jWv28k/ilJrCgArFxJ2vox5cDjWKu
9oM04yUH4rwrigv/tr4TlFYDoowv3C2pq4oAi7UynmuI44R5ERx6hlbK03Yx3u38+LuKlOlz6w5N
57UdMvxuh0NF2z4GlfbVa7L//v5jDWwjWIe1FfUBxJCG2CBRCfFIgLjR7w7AMv6sPo9Q0pJLil4C
on2EOEzLMsN30ZfIkuxaKh4b48w44rHmC/8aDvUTTwvhwE3gk6/rAYkxJP+FtvCyKSeluTjg4n9q
cZ6Wq9At1U//adXqYfEPpADaYmXNG8dEgGrWh7CkBsAzsdMep22EC2ERH1kUeVwi8cbi/+TUPgE2
kwHAelyziTZ7eavZouiw7MicnBhV3rEzfAunbSUdU7CKTlzkIGrCPgMgHi1qCjo6M3okepGO+aOZ
nWPlPbbik4ODx+1CCnmFdFUv5kiYrALjceTQHCip0jQIeMUac7LCYqvSMxBkhmCInASlFdY+Aaum
wnOOUhK64XjeJ7iqvYyfK3wyqedr1oiEKmNmc46Uet1SDmUJSlaq2x2aKuURsja5LYuAJEAFRn83
6JcCC5JE328qwK41kujFSVtG2WqHgkfM6u1njRjG4vKkQ7XJ1i+RBbvjMNXpqDV0SPKigKuC7rHy
iMjAsl53iJcyxfSJy7zlet8AlZqnIvTfdVhtfmo8kzeA9s9Tdwrt+Z66ikrqWMnAdczmSDkbVgyk
npvGI0AlNJYelt0DWMOxlCMYLD50OUeFY1XXk+E1i6wMRvFuabe79d8Rm6oBR7ZRD5nnCPaSG4aw
rhsh6FMKUhchr5txPN0Fh3cxchlCvdJnAURsaXcQUhJ0ET4yXXHxFBxCSdPUWZRt5rYmugojvqNz
XX5HupThsQU2nHiT8u6uh7GEAu5HvpeYe4pJn5RRZJ09q3d5ungHnRQDO90mkWPTTMGRuaLHtN/m
2iKV8gqT/DqwbV7wgSmiLwbx9YSbZbQMEJNXGKyit97etDJ8BJ+mR9LfeZKgHjk3nEsDLaBSTh48
n9UJyA8HqIp0+eEJP65MhSw8PY93xh0lA17KaNRGAERUv759wEnRs0cPcKtFQXE+FYAUFqjucPle
pT0+WmJjtFjQzP5g4CgInqa/4pug9epBeVlKSkz/IevzCbYuC+FHw593Df8gzzg40ygfO9D3iomf
s694vZV43vfXBvxe3Xvos3jq8ochs3AWtLtAMyvPnij5Xdudb6HVGmK6Dg1AYfWQdRORr4U6TE4N
ze/w46YMb5Dx5rZvFHZ3i73yDhuTyE/45CmTVHE20u4Sjj1rovkXfGRaW+EUYp0Tazav4ELx4uQW
KuXNGsLS27XKcsEIg0569WLG3H1Va6Nh1g19eukaddKOARQWhoyE2evhuwxlYlg4Lu0Yf5GU48KW
BAc2IeOjYNTTS2WGi2xE2TPB9or/YT6Kan8g7aVSkUJAZqW27w/RnIhMW40myjpRZ1LdMJlHx7Wa
DATtip9CDA9Kxt3tJwhpDkQvC5UK2xA1DyznnXi8Xu6jifN6G69OrcG8zQxLGckUa+iyDEa4dg8J
cgbwqYrhOaNl6TQeLedEYCxuhy7JZLdjTEog45pLha2B4tGiieMHL+GIJxbHAMAG6CB5uIuhuYTE
CipSigEdeN/1mqcYQAWqRTE566Oi/Swbml8+eqTtmMWeyWTb7F85xsIZOb9XTDDVfRXt2wWKjKrM
WpuDHy0G7VJrhVT2rsQ0eIY8r9eJnoEbLM1cN8F8MzZuKPyHkqvVmNG+w7g+EWok6di74cTJSiY9
l8GMpLb1YQhBPCYW0LAHVtswFh71i3kajopnCvSOtZNuBNP1FJFN8fdFLTaf5AD2BKtcJvO5ab8B
oypHR1OTuhO8hwWfrkyz/jStE1F9HTfmuNzk+ckoe+coy4HVAnU+O7EBaYnSFqF3ShFzbVqcqCPO
d83+gvw0+9tBSsKbgB91Z0i4qLoViGPAPpJtJV9mjJjRPwX5pwZ8WJnZPxpzmMnaJl9vDsfTZ5km
G+37E5VSwQpN8XNDoGUhWzGnb5k8/yNy/6As6I3zCKUWfiAqUVb7FXoj3iZT1MSiKqgYjnyiNP3f
tbHNSuHlt9GYLw8c9S66vJ17ouSceDs7V/aKF73EL5nV07afNUAwYrQgwKqMCXywowlbR3gI6krZ
EFHfeMzMeB/7mKFgsQPwMgRCZw5Si6cHaNDuKJGW7YYTEqRMCfNF6sGGg8u/1crfYGCw+PXOF7vr
pJNPGoDkMEp5+o61EV/XboMfNMe8X/e5QhL7N6FSH06fl/Nx8ITQF/AfHHExhkz/vx92g+hZvj33
BNYfiUFVEVoUbNET9Y/9w60HWFLOXSdoDGlfbk0scHX4dDNu4lWR28A4XuHJdmSu0K5nRAJECnSR
DS6vPJYhISW+AW4llrfxCO1wwRP8HlWR86YzEZyyhRtLUBW1DfcF2j7QhlOxsXTgC4wpr/9IMV5P
Btz7ozmu2FhVDTPyIdIP9DVEvaXDSOBJcGl1oZDYx9k1C79Dk+sXBWzdBT0wz/jiqlBI2I86+/n2
oj+JX0mZmJDOJnEpXWp+GceesLhGa07PBVzSJ5k7jMxnswLMdPxznTlHiEbIQxPJIOXma+2K3TDk
QUOq0kkKdDN/+TJfB4+xp75HBte8XU5tSJZnYw2X4ZIl1U9NzBldBKBwi+pTTroM+HhYbGGIIVi0
hydIG253HVvGI5gQLCYGrq1b0786JguyPfs5TK2iXabRAUvBSgI2DtIIvPkjFuVlxQoBFqTi8PZ+
kvGimyfqT3dSjL2pLoet7v8+yM9tC9WNP0XPvh017A91eXseRJyyo+LqNGgXf8Lu+mDO/NC9veU2
baSkwuT218U35rz5YCVfCVZg+Vg3bNqSmqa3KCpU/tA6MgMmq3W/69xYSs6WPgdAYLZMIRarKx1F
cFxVkugLU8ze6knoTqs9gGtWVuOkDp5x182yC4sJ0BRjKpSDttZFa2FgnMT60uPshB09wwkCK1au
3g0PLP+4zcjggJoMZ7tDUjo5k1EzSDnUbMYFC+qtxBU9oBKv7pQnCmYrArAmHmITHeQevQQAZ7jh
mKk89mxO6IFQMKwJcSdCvYfQISElF2gW0tkHNhDc8HmmI0MLF6xrgr+EBKD42J05DtxCRHrxk/pl
cM1NCdODRu8hc3dDavu5vNQnYAZGAxn8+g9V6UNA1rKyxG5sZI2+iM+rrE6RpBZStPJhCiYLfhcX
4KMM3z5Dkc1YAVrAdiHTf6519GYwgTu9XzrV8KQD3s4/0KZvUiA9Dut9YKzTSM0amk/EWXJEjzYS
lq7ObCGFp7JymG6J2cmF1DiRNFJkwcq3Uf0jSO+xH++G8UHLZCPWePyvZfbVwToYuQ62BVLj6LaC
3j9i9CwJ+HuVnTiaKtlhHv3HWyb4RjxlSqyr/+dEgQtsYHBWd2qPF2vNvToFoKNLvwdrbgDdvMeW
Ly/Nthfiku9w5ZG7L35VCU3G53wDaj7IAuFsvLdEst/EiubPtF6LHaqr5bWOTp8nSI02XwaXy+DC
DqmphdVpf8Tk1yuoB4bRMov+qBHz1ECgVha474E7LIA+wk/N0MCuVnOVn4bB4WioyHadXEnOhsNF
2layQOMfGpG/T83HVv+FPEIDepVoYiyW96yA51x/whyzR9EHrPjXlGfjdOgG6OaXDxUrX7/FVCy/
XaNXjahVS4WdXt4wYEECS8tsmdlyjtmqpE4zrN313bA2ZaCEJtoD9P9oU08saS1QZaXJfIOt415i
piFH3TNm2WbR6AoEupk3Um4tBrP7Ezew2HpqgeClBsvuFBQ8UD+xTewWvHbKSP1bQjbXFyWDQwmN
VKAVdPDqTuhNPiX77spoKS6oZJ51w1L4uFoyt+vpum5Y7Leu8VkmNbm9n3ujFNmWwIBxwnUM/rNS
BwzCehyeyyz6Sbi3W2AKnuDk7NnnfwSiZYydl12dIauuQu8dH3WEvg8CTpgZn+EoaXt0vYl6HiLH
lp2NbJssZxi8JnbfoeuKA2EQDd/zy2Ueu6dmyhrxfQSA8sZtliJgZQbxZCl0Lz5M2es40j560Eni
bLkGfuiovmCat3/kmZBkLB9/UvslxaZ48Fj2VHZwFcqYnYhsw0XkzRNClUin0il5QCgXoqJMW76p
dek6tkY1MGF4hYgKeFA6OV/78qxVRS+sx20SKr4ZPBr5yKXrX1iv4Cx5ZH8p9Kur6l2vrQIApPeb
hQvGxNex2qcR8Ne2sbT+W1mv1PSXnrERGWyhy25BR0vQLfQrfelebugR8nqvLkH3rjyz4XxcyFh+
MB2R3leDrG/CRfSiD6ZSEwf8SQWX2EN35vaf6oB/qRdL8TzPIoKBX1TnD9Dk2/ZYBYXas3/2eLej
BFaLsI30v+LWW9FShnn/dSVwbrp2sniCFYjN9ocYNCl5hZvGzoQi5AXM65D/sAW/08a0/raSNYYC
dT7rb1EGXhiMTOIk8now0PuxQLryDUISERKUwTTp/f5ThfIK1hhBDwoNDKZwx2EUkGX4YMhH1L9H
oCREZe1250zSOJ+4+BOI+nBNC/w+n/0vv528XHjUcc70ic3GXt2WW/l4QI9oK9iYbpul77Sm1HAR
QqHbjsNvknpgDotZs4iLqyeFX23ww347ggOLbQtFx1KzS/jOl7MCcTQ0rzLY33zf6WGAfsuV5+JD
yNBC7D17nJqAzfSV7cW+DBBnkgOvHxtgU0emHVQNKOYuCSkezyhbuVvQ4OTjo7duFozf6s4ceqgk
+KOWP6m+jIqxmfOV8vMiCJ/BqIww8Qwu47aZqp1rd1GlkmoDBoC1ahEVFmzFNCraCc8aWt4Epw8q
1ZYO0YpzPvBizp8cnoM1tRqxLlUjCLnd2JIUv2hoNGepx3OiO5CgW1QgTQ2B5x6l7Zv9cwWxy3KQ
J1xASDFwqeXhwqBufQWrCtcxU2JJ6KcDdyEW7Wk/plFUnf13gnB8DXlMLjm4dmol7n4sSgoleDvN
z1ewOiInLSl2dhEjahDDm33zstKct6+youGmsIeT8Tqz0ZOd1+McWkqzPAjzxreg1IaR4Y8Z88Hr
NBaBt7Ss4nyThemnTf8nm/bd2gaVdWfeoSeZAkHRQAA0S+v12ZRnLh1juJPHvICpF8hLzcen+XN+
IXBqzzoOKMRBLEFu8VeSMiERpa1S0DMogtBg4iU5lrsXsdMP1huDQohpnKtyTK4L7XjB12Ze19ns
UOqvb7KCRSQqEXJZ12xS9sj9QclCabVB74M+9+CgRBvMCvYsZKePJZRSD6FrKYusX+08bBFF3RdE
npWarQi72szkGe2P8Qj+46qtwlh5NwuwKZcHE9y9a6Y8Bbh3YLZF12If0C50T6B9Ovx39u0B8pg3
CDjib+KHhMYm+CSLrpW/NUjEhV5LwNs3bXOEY4i/D7PWYn2CbMfB36ypi5eeohWfAl/KtcUFPpAg
zf6LAeMpuRDGedSd6HS3f1FYFNwJ+m8XpLX9kkll9IJTfJ5JUw1x4r8VE79SRTte7R8lWSfxxjBu
fj52oLXh1rse2UuJw1hXH/7Ipo25IYHKvSf6GuRaIUUmHWAzD4qNuhEQL+jIZY6K9zU/RUCWX4Ly
Dsry/HY7r6sxm4iPxehgFboi5qk+WVVxtzQBgEYg7lVqC8aY1wuY0Pz7nhTe8ZZD4ohDJhMDHjuc
AF61IDhlnOOuotzDdG3fWMR4CXFBeTPbiOLKNn+H3LwsJioZq5F8rz208bhHmGVgR2KI1HTB5EPm
HevLyTZDwj1ar7SnSb9C64FfMqpByKkSG8FOxrjKICKf4qnZS8QAbxhfK024FYjybBj1t74CD+1z
D+uOtKjeubbwh0GN5UgQHsyyFQTo5uarzQwk9N2bAVu9QoQ3ncqi1OkQstwSbhg8fhldg3FQVM7x
wL0ItdGs0MC3qdIGmJ+Lgq6rMHESZ7Ah5zq4drraxWL3ipXwL7TyUgm6NbV/j+4jl7LtNlDUM7wE
gzRyfN+vOY3qtjHxoiIkqrtZTw1kA6RJeemyJ7Eg216wk9X0zAelLcuhy+x0Y5gu4StYiSYFbrgN
ViimthcjRHuq3bR7fJz9+HBSSe2mM6A6lQncVIHhfn+y+I+o05F5Maiq/Fj0LCKMAi4jdH24cJ1G
bugu27G4I7B0VBIWGxMMUaiDlSk/GSOeIisvgp8CZfltdf5qunBUUTGwSjOWzUeoUgcv/qsgCvRl
ofyWHuHZNn32dedM9+vGM4QW5PJt8NH/fHcHYoGUbRxlOKfVVdfEnr9ErFx15OaDvsz/EawVWta+
ssKOGKric9h/c59kp8aM/25u0c3G3mu4LeHnMjbtvJsWxpslzV8q5ieXSKxZfmClCTJoRPrIiF7e
EYHwz9BHmrDKbzgCwDC44O2o/+IBjm6FG0QXiJSk1snF0Mxch2XzPHLSm89kjE1PUG3XNhUDGMwN
Bpk11UxxCExH2+T6FXyV2sfmoH2loaAAYSkIjVvKMlhnV0RvFYYTAzTeoSaf5uh92zQEl9AMPPgZ
STQlro4snI9iifHu31w1MoFu/v17mYmmUAm3eqeGYY46ZokOYNMoISEl5U2jQT5FUcODuDXeXxYy
ReYkFvMih2zYAUzd1n9lbUAfp3szOV5V+Gj7UmQ+Sqmpg5wAh4nqGRLNXDixD9W6kLRvW7ia+lt+
yvjPyxuEq2T5cABBSqjoPMXKgeBIyd6Ie8YzcJjJaSNDW26au4Y3une+roLatPKY9F+ckqLVvVmk
y2CpRRXPUGBPhukWTLQ2aq/dkbmcVHQLhAqbA8MWQ6OyobhvDGi7+9kVBlgLBMVYF/uJnpU22kGp
3Lb5kuBuNXtaIwRFr8otP4TjOc600SmlsPCZkQbXAFcNb46QObvYtN99ei1RWgtfTS20wOHnzyPB
O6HiPPHVuL/VnYNEVrIM2GevgnBh+ahcapCWcbQepDOfl3Nn9ElYUkX+/QvdZ5aS5l3QeAbXE8qo
OCp1/l3SWGc124DFsR7Gk1+ySEWEiwtuMwdOyJK//5jJp9JticITGyptG01EZ5J3yW+H/uvE1cHk
32mzzyVy8hAjTXzBY4U1atBU6kUhRWR/DN1sLWIBrSerkUjEbwfNGQnaIfweynLvmiB2sag2WCQ6
cf14xptH/07VaBeE5r812JIIWtPzwOSNDx8KqkoXpEDNHM9/T9mqI80aEBj4txb78C6Fn2qtzMZh
ool44KWaQfI04t+j5nyb/6EfHWU4rfgobXbXBlyOEzEyeDUyo9g0iA13YW4rv8sVqtIXiM4wpaWa
J1GgJxp2wTq5U3KAGA9pnevaOqtouXG9XN4v/theZX/biQhmQcBC6/ShfK4AcX0ZIXAOlI19HvFd
IRWOLdMHFeLUu4cROkVg1tqJ1oWewEtOGQ7cDNdDj0tGm9pm5J7iCf770QFMBmjCsOSgSfFvVzUj
rCY3KvC2kl7SxCLf0V6SYR+6q9VgMZODqBtEIpkwjpWCoH9m8AETryGEuTfi+PFiQFQ0Ch46++xI
0+Zzm0QbBQtzEC1mxA/FGW7RmI4/0tlfi9Jk+FpDTFgOFovhjT6yrxkTjSLKT2kt22II9MLrEZCo
GYnIYnuRNTGzszbKOOHUOZMi570SxVqavI4T6WZuRzzP966wsfAZjI03LJMIYj08FpKG7BC2B7fg
ZiX2IVfhuiWoO3wTAMpq7zWngMSSZVlpf5FtPaqsxW+Vmdo5rw7MdHgasjTZh1Ctw6CCJPcHjF2m
qODGNgNy82MO+AbIzXHgSjmcvgMkMZ09Jna98ajmOfmpmjgDa2CPiD1QIYlj2x8r3WB0D3oYqSdJ
cXKbpwG+A1sEHv9t2smq0u4Irz14vlalRnaBjvjhM9GzAuw5gF7ZW5fgBEXC5Q8yfWE/JieSVVuU
8PEJsPI3vdBWSfHIrhleXpVGf0mTwBl4a3Qd1CsyEkpKFgAHYRdyNtuQg6X8EHPYG1C/sObvdFkP
6kBmTUhbemE865Oori5Z7O9PUNMPlaCLzlu4WdTutW2L0EE1dWMzf2eZlfaklWb96MLTyyAa5oNY
YvxkMLWIj1sjCXZmP4bAOCtw/G/DHjO4MbcJPXSuNGW2TskjQspVtN1vh5BDo4K6MsYqzgaBIqFc
LHG3++mIUFzcZ6Wwoj/f1HsQilmZYGlZhJmVA+XenI1lqRFmGF6fZq8JoidCkJBqkdXbcLGzGbC3
mgSyLBaGB9ExW28Za7+bU7HfCY70TrlJHPhHWncmdH3LyHHenT8gdx5XO+eba826mmmaeerx4oOO
EyP9pCoZXyYux+7noyeFsSSthwKKNsaWRWvjJmk6raCufN4H8ucBOrCeO133Qo2SgBpnA6WolgVW
pWpp976z9L715XOyuCm2mHWVTRF8HjqJWY5PU+6gaVmH7s0pMyE9iM40tPHm76yH5kar8dty0whs
vtg5d667XzuQsYCspz+4eJxTpGfv47gwJKR6u0N7JBzr6Tp9xw1FV1TS77k4SBJ71b3biDSVSAwD
SajEK9gqGxTK2pce4AWkvc56B74/CLhZGjF4J2Ii9uUIlIqAMkBRJJIaGOt4FXTWxZD04DppQyYU
GsP5jUTTcg6nB536qXa9ZGw8yPr89d3LCWaXtwWIXFTmePLDG+0k/BRA+p4FfYw4LaLIdeI30zw3
wwY/dFDZdffK624O588fsQYl8LLzOUHKy4LkJyYmf3SOqQeFXlpryGorjOuOoarLbUW29yRxYKvW
CSGwMG+ixu7ev0DUYwEfbWludFrziweXma0WRWPUCVK1ExbW0bDFUSXdtuRriQvkFUmAuBAwKs0f
xZwTb6xRfrZXtBZzwT8AT4Qxw6qq3NU4XBeXERwPysbHJh8C5CoqitI5nnavfydm/v1HisjnCsA7
0tLsQrtK4KyAg+/A0fzcLGdP3DcNtVaxSJSfIEO2o/ChC7FW3ZMrg1ramPW+d4gvGyL6b72TD5at
P4y3Gip3+TjUNIJvRgW8mqPy4X1MAzKMMq0+I5fyiwo5zxHHBkhiQo7nPOgdQQg1DNlwf4bTxU/g
G/+nnAZ+K+I/e67Xeag/0mvITBeja2JvBrTtyhpCQb4p5mmxxrXXUrk9Zr5R+4tVF3KPA+AfXGry
yi9ausB2A8LQBxbp9eDqHY1+DtFjirdS/Q5Hx6ItlCPI55821DhFAMKEw+03oQ07mxqfLBxrLADw
ODqiAsUrMPNxSTPOJperdra7RMo6I/aUh6WTt3NduVhNix3Eeekq+xX4MGlGza6vQ1jJb0lWbQbo
oN/balzyr+vtKBt1Lef8hUCZKHK68UXUK7eua6Sa6hL3Y+/TWy0bUZESE6tATCpH2bnBVHXYQNUa
bvoatMRVjay5/GDvPkmhgIYxGOZqJG+47yhnNYTsxlAol2fd4hTJev9bqTthAx66wT1uLdtbytCo
gDf672WxVRpreUwvehNO1vIZpJIVniBPYdN5TN7lOVvo/TSqmx4gykeqwksVULIebZ5wBJQgSDJv
gYssVBn6bz9VXDoKO3R6brf4rbWzrJZuQwP0dyM3BXVJveEgLg04BbFVvcaCCyvn/3pgqOlFbzpC
HLVq0d7/5m4Or929B2ZfC+RuVO79K/OEkGNZne5eXo6dyO3AoBchHFWUtDYTsoP0gVOyvs5HcMpJ
kt02F1wMJgLMZIiFsY/sUsLrSXLTxOJ712WilspQiaqJek4qncUWGQ9JsrrjXjsO3S9TvFzJWAdV
PtMnIMXUotuYB6VyL9886xHX9KVSAK6rO8QZiBIqoyn+qMmBRzgDdBGXPiq3smy7n19dACXk7h0T
u/7Xhgcj1i9BZkcftaA+6lJKUII67B2ziJG8V0p3QAO8tVlKnbTVssVGQIVkvHY6TNfK6tSHIB4p
3w5BWHcDuYHnAhoN7F4B4MNvDEPVTjaMevD8PojiGsBtc/h6ukk68rDbTU5sT7SxCnLq47xhsmR3
t/5SJshDHgxZEx28XGBIGpzlUKL9DtOdwKz2QZb+qIYzMtPnObE7r09ujWdoknkLmACir+ca0a6G
m2dB/W+/sgPgoxtQiSV/giX0N+sFVoN1JP8muz/pGBodjdDriUphp/rbeeGcVkCsSX1GJAi7aOSA
K5Bq3PfQ8eII6bfsqz7TtNvWKuoWcqjQvbSFU2CfcFgmcotmQX0ZhMeWpFfqRA0y/oUZNlxPY/MF
YqaolqDRBtj89LQhV5UEfi6bsn2EPkmjLbPNyiw5lC9SjI4hMJjrc8cOOlpHmRC8MjhmQxQ5Q2XK
ax54Y2gsBQXJvLD9sRYleFiKhM0SihV+OuKjOL3HgTt7+1/F2kwqQ7HMMkPRJveDvrFWgKoCMJzr
onajh0ZNwpO4ct5OO6UvMNntwPXFuFgPzZxoKZ0mSJsD6JyXZ5cMqpH3KJp3bCe2+2Y8oR5YFZn8
plVKQD9WbajmSGxihKv4xxP3UE6Dle1rdmyVEW7/Fys7ybIIK8Lnes5h2PfUfAOmIgRXduh1nYd0
nZJ9GSkHvXqZjuablk+KmdDMKDM/9b7SlHU0NyATLuSMOA4mq4JGCUtfcT1/k78Onodb0/Hf7ECE
jqzVl/hIVzLiRvF4DFomok+DZqaULvKVNDinacllEpiqzPu/WGVLNMQNSJolFNZlYFOIj8pFmIC3
56gcIxh0bc9vZzqREHh2vrme9RcOh1Dphvl52qihOgYMzGTLILNIkxevHNYnXGpU6ugps0qSADpU
b0drxTWG6DXa5D0oif0+oXozG9L3jK4WeiofQuzxBFP0z1Q2BMG0AfY1jOBjvqm/LzBkumMqG5T0
cA+bbcfJQtMNm1LSu6FdRUW+eV/JDVtHJrg3ucEZpQMMGmK0yEPkVRO/JY140zQWc8k6wkwu/uX5
owo/wlchHRIGnEdj7UqJnKmP8x5c0RtwAQHltktH7qH2oN1wfiAi6kKRY+Jk7vbwsEFcwBbniCOk
3Mgq6gDnd403nNltc3smvOoQgo4Tc6MnR8tJhlkwx0TkCALyDpVnlRUr0lEtOjBL/VUI0qU4bry/
SkuUmpDiiT9x+MQh76ZdTjhkaM9n4JBA6c4Ojn7BrAnX7QOas1YQ5zyCuEL7i3kFX8TF5qF9ZCS2
Rx4kg7gIKnkyAsXIsiP+wdf+vjORdkiz4x22IdS8URzXJDo6fQtEACs/vLzZ07Qd7Sw3KTVAkQg/
1TvzQDgkAe46okwgSqKdgv7jwMOcFPm29alCmHr2+a3AvjVmBLyTogL7Ip2vcBtEr2IGLz8G+tk+
KtsoDQ7JjEsH3+EPiyw2YFtfRVAOJLnpVGfN6y4lAsniligxL0vRw9COHN2VV5GGz9oGNZX13Znq
DsqyAdTNtvFbpttalA4rwZPQAyBRhDUrUtNgFsj5uI3pIsRKTNs8J9B9NHm7V/0aNGfiw13D6BCt
hs496/j0E8gMVONtUspK0Ub25RBzHqn0/YRGQc9+oByVf6HzxWuLu+cO7wkTHyIu+Ym25Neg4vdd
JgaiqnhHg6lc17bl+M0EJsXJ64Efo/ruZb5kcfgWklY4ssJp9w68DRa/KOnMw5GegDmJOLLBdvjF
j6SbuAsNF6oCZzTiSEoVbhvxcJ0w6AyhSUmNWI2LcpiBDPZe5bk8Wu8M0BuhSkzox36PzMvRtrMK
CRV4emCpWtIMl5sx68TZcRpDAO8xKPAKhiUPy/Yosb/czmdsI0MDRTh9ugXTjuPhcPN3OMIA+cZq
A/OMWQbVSGp71Q9eYKHBoEMMaMZgjTzwNwxCH+RPXN5ojphG5R2KO8/iuhCUxwE46XIjt+A9VsDz
S2QKZFBrSBJDLSSL9fu2Yi2hM8sG0ex93OVGghvVNNtrxcONu3N7QBU/LtLWIM/oUuna0svqmU3U
Rk94oBwqFyJIzM6TRbBaEbre9+GmX4THk6uXSoAnrrWsKdmhs86sEP+k9GAaXEE79+iqhJBWovo6
czHTrafI9T1TS6xk5hjgEcIyV3/Cl1TXQsYDXtJ28bHD8TLItqOyQVHTw+M+JsGzGwTL4YrYrVOm
DW4UiPHajQOwWSc/N6+GyJo7GV/rYB6JUeHAze1fS4JXtrN9xc50btKmYMrAgE7EgeIigMiDlwbi
2nzAR+6sLnTS1cpHVs8fQlxrjk+5W16tmFbYSlbl36hAu7QKcjlt07Crt3zP6BGwzh8txuwbtIHD
oVtdhc+8r3Zhh0aCuwpKgC/sGCkcZuR8mYIwPGaMsrGiRxZYc/pISz/uijNa3+QA+DKL5q41Ai5d
K3103QTNZ3ofnZ48yFf8FTEkO6i4x7X8wiZurjQKObE+s42wzjy/wMY3P1B2ZGTUALnKovlAEAV4
jCPJXg35mu+xUl01AH79SHQhFtRxFiqjToO2H0xMUCGld7w4SkneusU5ddFKyMH57cJiyKy91Shj
DSF6gnWIIelLzGzJSnQxcPTkb6q5OJkJ4Db+wMNs3e72cijTi+PzAP6PUtEukN4xWIuuRtFdzApU
X6v72tqn6jRWEEf+LeqxX1A4gZJjPuWXFtEGa+mG0eSKXCMQ6uLlj9LvhJEnPeqTaug89uiJIBKW
QUmQMCz5vEH+CftWdMq1LzQ5jilURcjKSrxGOSZdlfwW0QfH4AgMkymbk3Yfr8TxABclw0a4jKfO
+qgkzZvxzKRwBUt018lMJTERAwQTLlRvIQ7jQEEr8ctrG0neOyFIE3V4ddAZ/mayot+vUqWpHWov
dXzyWCrzca3gaaKCpKiv8EJb6wWaAvh0muq/tqfPymWVboMXxu9bmvcae/AIwHU1Qs+NLcTPv8/L
RztT/jodypyFrWfTOTS8tJbdsGtKOukVHf6cqFlqNEtLbxyTHG4Z+cVgepoFe4qCAPzSlAJwLb3t
xTg5/uOtgeTvCR3AHUsSCHwro3a8JMGBrloghD75Wj6dz1AcpwZFiNrTQYzhL7dbr8LN5CCnYP93
/8y2YKiwtQlJCJuCDVQQbmXUN7z8qjoHn/NKqcmR9YNOjahgGuSsckl0/CADDC6rp4rEP2oCBB3U
8ag16kNqLdeZTMEN53WQ4dmiL7r7ZT3kTQjPItaqPMsUomP4zq2o6wmFZJFuO4jKlMX+1D2FRlvE
vJtoMOFRulOHUQwKpc+6ACob0uAZGTVjcJpqdrfVTfDXZ4eh4oPmZLvCrW+r87fBDVhsIhdIxYTN
6B8LVBfh/5I20kJUcRC+/ZK9Gins5GwFQg1MUwImkcs+aE7LckV+Lq714UNfb3ODEnbwG9VSEGOP
ff0S7usf7cPcXi1vK09oyyvQRqq6ipCQ8pBuhAYRWSgmE1LnQFKXDB2g0tntwB6eQZ8TGRsD/lJv
CtK7cv+Ow2dQogbVOTip0Li2gKUTWLbobHXqbkNSooNuUWlBzsDQYCIx6kLKq69POAkvrXtSdMdm
BvDkbRy84bZQC4ILsyVU5JB2tA5mNagH0TJkm+kXVCL7De6X5mbjtlopnXGcLwsEd0iRGujm/f7i
9xFFNaEVoXblUOoGSh33veFExu95B1TIuIFXmCJmHFjzNtjqPB7si/AccFJsQ/xP37zGw/eubjxY
OoNTbm4cNDEL9NnlgidccVlZGJwfPkhmtbCfYlkI1JraYREiS3/BEym6g+6reYKioPToktLe9/Ee
DLiYgoLX+fn+pJ+V8NPM1G+YOCm9eT5qu0AcshVkp+VII6FQ40LIXNJCDgpfN0iH81bEnDGHs6UY
xnofm3x0UCbPuX+EKuylrv46fSYA87LMu3CwOcCdGyelvVxEu27fmbvdk4kc9ThYBpvXigjtcB7V
vPArCiQoN/81cP3FzazkkVKwBfua34jSJcnqR2RATXj9jbgfRLA7WddcOcvsPBFZwVlZHUoBENnd
zqFFBztM4qWUeC7O2j2q/0g7gd1hrTQkSfohD4dJz7yeeWEx4WF7jAJd4PORqSMGSmnNjUT6EfUJ
0bJ36Te0TGuhEK6tis3PtJySpxNYdNJuLay2bLlFgJWa69BpA2UbJb4DA3zTSnhskPqHN7gGO9lB
+4xkL7ho5jK30os91kzCdSOJ/Q9iPWA+3i3rx6SWOVWq8uFELKlK+sjDxFsVYTwvynL+7gE6Zfdq
2fxuJEkl/gMIIVkNNDbmcpCcTzg33x39jnkWIsZBhFejNbM38pDw/Rx7Cx45C5ZcFTaxj9YdV3P1
xty6Ks4SAm6u+pcHQUdA3yeew0ZxWmS4RKbG9baXQ0u+ubRnq2WJmT4M803QYc/oX5X5I/P1MG9i
zhIhBKtiTC9KGxZfur7pSkZxCImJZphKs8eDj7HulRCPXLgsCDzebxQOCDwB6fHr5nyYGxSciiiU
yti1pdydZQ49PetVkeTtVUN2HpJrIGFMHeqEZo2kMkWUxGERkR+KyPacXgvOBRPk8Yobwdo4JpTC
bCTm8yfyfIefXSWwxoOQi0gmtBPicbNGOBmseTkUWmHrKsLGgaJrdVSxSVekE6dNUdVdY7ID5DiS
lwTN2mZGbC/+pOjnr3E0LuT8hbEl57jJR7XD30zt3iS2/wz3UEka5/8i9WrnsbGYvqFGCDpPA55T
Ozt2afpDURbxVa2kEqFriNQ59AeEsS7LaIQmMeRqOBC+jkWV7wv42pG95xgpP2O0GLHN30VPLAOm
V7Djnm4mpPxYitWfuOVtsrsuy8GkYaTxwuZo5IcWJUNuSThR+ININnGdMeW3llRh9xkF62P0lHg5
x2jtBLQyeTbSd5zPkd+cpbRIuZj21g10MmlqPsPZBVHy0pEZWD1ZnF3xseH79fNAze5Edf9ZSF83
xLJf5mR2Cen0tydDbszWnlcQY2zbAS/1YECkhRzgh7un29MBsqe3Sp24u+yFQPGgJIFEdpbm8w12
YUkaOgCtI0AhPnf8lFwNUR5tU0WikmfMi2Rem1O8IKGzskK6hoqQNqntNxum5jhOJuCSHGE/Eyc3
DlID/3XK8AIRRZAzFjtXHsgOa5crlwCHyoXuEImQyDS7UhJXKjzR6m7nkXwxluHwNoIl8OiFZqGk
Nx8HddQYwLazQ61IKthSD1LUXu4Qv2FtKLOw1CaB7s6kp3Uy2kqDDlSSBSd38lmDBz72XIglxAJm
03SwEH2mGYs00a04+ya2jsv7gl8EYYI+SYcaLvUyJhnqntQ0081RcrK0HLDnxjSDtbegjQCBPq68
SLIU8MG5tzmpVJ66LKmXeqg24Gm/jXzs1piFiSUQMGLVwJXmahWHz55o52vtAOqOEKwsvrjYXAZB
PzVJ+I360/fSn10udsee7CQhugF56zbDvyXYs1sJ5M9N5kom7LOq2U/gFun+ynp4EE3MGeZ+yhuD
AhzrJJG4GD2r8vufZxd2lumQt3UPKzSifuE9yOxuiTuAvF929CCiyXnvmVdbvseKw/2Nd+/mmfv5
ombkacy60DDY+rY4OldpBEV9k9mpNoCrytYrs57o3V9k+VnZfiN8WVcbfgPAnW8oNWzV0686gfVk
hzrmAksMrJxXq7qFlWuEh+OXHB3gO5MaSFQ3LELzudQrQumz0CkoiOPS20dt5MMBpzSOowfdLyGI
XLt2+zqAlOHvtfTZAhHoYZLb9FMj0XdXVTIVVV0vIfP5dX3dqCQvEnbsFrrrcRUqE0aXmfmkcnYj
BnKVkXEguTn66WdCgVK4+4hXh/1QXdQxgohRsFpK9VwvPqiJRBdKflfxde8HFH8QzdC8m3/iiv3b
rTg7t14i1EVxbVwEgqHI3LKQRd7pZQHW/QgfW/DywH/n6yQpkn1tRy9BXxeuZyeB4HANt453gc1i
66WrIdqgAYQlXi1N2enuYkmKydPur+0OayaNMtb8K3Qa3Q4ofHI4nxlgytqxCskqs/EWAjrr+Pws
NLvmyQezS8Yfmn+ifNcCCJ5xLkpI5rWciv1OovYfM19eZvq+D7xZO1HivAz/XhMACtXmvpeM3nLn
EIEmHwdL+tFuxwaPql1rqJ/sgEZV4gE+shiJ9YUXK2XE8Dq9we/DIWKh5WJ7YxYgl26kYvvvdYCT
0t/J1QGlg6zXKUjEdTr2ka2xY2CFAV7Ihj59O5+MrBphdwS+Qggnq8hzEsp7X42SxKwqO/PFpJe4
ko9ZnmcG0kot5JRiWPljsk8xe1S77jXgRpepr+wBL9OxC8OrRIBfTo1RWv7YIuL8Bs7e+rER3bFj
GUW7fn+lxfLpGyaazqjxMKSQmueBu8dgkqTspv9HJ610FAKFw1a7RTifmvCgnTHK35jMnrz9DHmA
yorvRs2CSnxlqswRS99aMi2MsNpBKYgs57aXZbIcI3sVCSgkV6AALjQ5/ZFw3uvMPGvLxJ/Ig1xg
BKmuqVgyit5fkjyd29ASvIqtmI/5jclXIFJ4bQWfo1d8sSt5332b4R7hxkfjIn2BC7nYOiN7R7Aq
fTyQ+9FFf/gBofidJkVepIff8iJG94hfEXbUKcAJ+QQf4CdD76S5ed6YmMP6NtulbQbvKtADP//u
km0k1FyVwVYowrv0zkUmhmX1pl1X4DkPbkulmnlX21vTmnRCB8UeG/7/XAK0lld3MGCRZvw7SKH0
mSXP566awtygEfrOae5bS4pey9YHocfeC+XAqkZO8jko5Gc9AzJR83hhCsTtd2gjOVRx0CCMmQQG
q1R544v2YEjdi64zPUIen4oX/NDo+C7m9MZk8lg3DlAYcwWAClnz+NzJ9mERPjl4qUjZVIdfRTb2
lgV2wtjP7A3aubfNKMX1KQrOOszLNAVuEc4KpiGVkBD9Yop5y8LKEKceQ2VflRZkrWVz051DTc5t
gUKWxLJGThGw8EwtgyL8xT+bpEoYHCuPPMkHD4OkfafZUjjJnM9+cFSW29zJIKfVEjzG4iair+XT
LR2TDMY4v5LjCURwpWQV5z196i2mLQblCna2KY3lepKzEJWULHcFj3tkhS/juXvvXGW6RVV0Zloz
AaB2vTAhXCnZ3Y74Z/sX7fJ3/8EFcSjzawhMMbFHJLfWaSsGqJvFWGqbDREbHslHusJjn/8kTatt
qwfTvzHqgPaKqySGcFLySI/geDjqneaEExpvkJdMwf8+vhuRKGn2ilK/mveIuXzU+YteX9T+GR/t
uwDsAjrsMx9qkifGDl+hUtrhUwwNpV1XIB4cZ9rALlA4MM0Nq6/RQiaQ4mpCO2B+H1x0UxnkLyN0
Wa+AbLJWwYspZd3F5jkIzK9M28DE7TPGjmqC9L+LhHodB+mmhjlflzf0bDKyW0R4Odn3dYjl0Qqt
C1sCLtyzysWRE38R5zhrqdXdXKwfhRuncErDKKVw8VfWrGdlbTxeQbG5gZshQoia1Or1B3p/9bN8
i4v5M3yLWiU7Pgkf4SSKMXR8gOymhXw9WHUGWZnb17vBr/LX2fwE9PheBcftmNEev5d+9jxOWaoT
d3QwqpkXSQmDoRu10bGjYyp5G7pEFBBpHOXCviFTVDwX+8SE7x+ULnP0twK/zR+NV7tTR5Y6fSzw
VyqU7yGbLk9sSGYZC5RNgOXbk71jc0EDApD2XL6xs0T1mobHSRzi/7C36+Tbg3NQSkb+sYH//ksu
Us4t+QC/u0OPZD0/oQo3pD639O3kteng3jnUIIC8mWSvVlWC8VebsJ3F/iVlBu5Boh2beZI0GAoA
y211j1yWz3T2uEQI5P38qTd92F9ypi3/wCF8rCnvzvYtpoUuUpxptEM3PVEiLSWzVSx43gH9CRrG
jwqzn5lHvhz6k4MF+uzW+cIBTxf0mu4ees4r3qZt9ka1D30X1QG8AL2KXcbjBBmZcjDuBSf6o04K
SaVJYQboXsglEcNeHGqa2tPBGgP/FDCOQPVNDGS2PNWhhxtkmKxYNqXYHX2TJE8qKnTJSsybG8oP
xnKt8IhV++BSI6ntlknWou37gew9XAGUN2lVgsd25JwyTrLS4lSw32VCVbrc1eH5WrejeCjBPONC
XfNV8YzNZkjBTF2meTMpCeaQFtzhKonTitf/j5nW7ebbSwtjrPdnjMJWaV6OHBJ/rKKkbur9eCYJ
bB6RdguCY7hHP/AIWRY67mj9JZrHufVQDkwwlzI7ytcuQN/mkKNKONWDd3lybLe9hTx2lRFnRdU4
MjwP0dsq3VefiYC/BKbCmw8T+2carpPnUrMX9JUw7t1ktMe2KgiO9XgZK39zVp6uvk631eeoxkWK
nkz/FrTyrT3sud7WTCyQ4GZXUFZBom4HL+W/PHgTwUL5Jv2sSHIuVlJvvRuu3yWCzxPg2CfpY8Pj
JjD7vAo1fKkhCkq38uZa2Hx5NpwUwN+Hbj9ch3eimoiDHM6TbFMFvp5ZEJbYvMdP7478NhkcGIrs
mwmkyVctj4VEJ1UqbLi2rt18QqAVWQo/pR1wjTLKsJJpl6uy+rP0AJ054kwCYXx93ezs2sVu3KqU
8zsAXuWxmbLAb61hRXNwtT4XvXEBpMxsU7wL/JCVK9/1/kjhJco8mNtXn6KImaK2NGAi50dKQs6z
gaccVwtqSgEJEUTHDnO1PYWKLEK9Npn0sjr/o4lTReDsxwIw35c8OoFRikbIz2mDL8mdMmXToT1U
BB2ktgxm1lLfFBGegDpTVEV3GKe7wdjVIVuAeS2Sh+coGnm3obU3TGyw/lBmUxQgQ/r68rJWk0M8
PMOWwcXooT9Lb+px7n/by257xT4oGdHEVvMlL5A4bPf1/CXvkkyRIf4BXkr6vhLO2jlTtK6/9JDe
3Y0mmb+CA8lMVe4Br700mH4N27c2lI9Qou+pc3ZtvMSOzVH8XGOUbV4X6bvOPSFJchK9tXd1WLih
d/XXlfLCZf8rmM5c+Fy1YQhJr2Cjq0ShWQ/dTVKw3f/PY+DIJiwSZiHr6vfbMyyC7DOo4vqpr9Kf
26pq6x6GLPDC5NB1t+FcmfMJiTspItEhZs8Wqs4OZxCGf+PyNQJjPeEBEhOoxaSyAmaf/kSJ02QD
QBw78fgvDm8mv0wQ6yiYIcD4uWrbsVHmUlyNku+XQ/u2VwPN9PSCgUQrpbz9JsATa6hQb79X6eEB
tjCy0pV6mqxcqhPBasda77VShDtyaBPKKMcSsHcIdybZbjXRXC7HpW9vE4FRjCpkM+eoMpw4iPx6
ym4rIVBhkPUPLvJeWVhZh22ihRr4ZGkIC69cipjicFcq6yunKGgFmd/yXONUk8fGBZe11Ys3BlPX
93DVvD3ujFCzBPmBcozv435b+VYXEuIPBoKsfaYO9uAxYr30rD8bkZhmVDRPS6niu+SReOP2shGl
CcGPlyqj0KBy5IO+btA/3WGxJfXbOcyOSPiHlvkG5XmYZDqr+rZ3vAHyqqNsE5DyCacaOHD74mxe
4qaSaiTyda2fg4UFpg//+0OYTkBM/AAakeRPH2WqIDK9ZL/jE9vNp7zex8Ddo85/a+CxC7IgOG0N
iYI1koxXvGWAIkwCiDdEBqLb4BRchsIcm8q2khFOC8MkGymUP+YTPYRDXG73jRYZg9aSoFNmE+69
ExWI5l7NgtaVIzeeZM6Zu/Uf3yvXI7sT2f1L7RnyzTGPdwcHl+3kDoPPQ2S25l4S8C7KMmYbfchi
4fntLSg8MxbZS3JyBcFu7+5ah1HI4joOZvUqer0Tt40wau0D8i1tXCYdIDPBzrFpiFGowTAVS2/O
I9E16xkx4K/8WaQ9U3aOGm7/kMI0FYvJte2k0BEdi42BAdgD/BslDg1RxzmsNxYWCK8A8i1LjxXw
pWEWMBLuD4Nj9zQCFDnzHv5ExVbuOi1dDie4gofQMxwbqIIxwnSVhlFWk/0dz5sCCutjGVys+rXV
S87HfQSjXIqFm8bLs4bbZHUZa8AqEJvZELQ4o+qDMSHL8bVDY1VTYVefYZG3EEWx2LiEfZl7TfKq
OW8qrqb3uksFv+8EsGQ3XSIl7jEuhOAVxDVuTV1hpwangfwBVuVM7YXa45cZZZ6/in762xIcXc4d
KrBZWuxmqEz6rRawq1TA5Ca46t6gVF55/03pDXHmnLvX0rO9/mpMaQlJDAGMHMZxLG7wbm29RA0d
M+sUW1L8BFsCPpJZSIvGZja+f+9pGtxRxGAU29fYzetgyVgN/1e8GxDicBZz/qdxXaMWlS4CR7LQ
X5uAWkz+i9cCNUb3y3NL0yBiuGKrAkfctwU8h2TwTtr4VyLBm5RrLTeStjTnKIfCtUM2z1XL/KE/
vhSXanpRT3h0Ox51+x0i74R6h/2a10YPRhNxOwLoERjK2yuyL3x3GyHE7S3kzvFoQxOxAjtqjdj3
FOTnIx728x1Qj7/VCHKUZNi8Mb9Jrel6FlkgH9IdhoTlAOHkrLroJrEAraCd6TBSoPnVne3wo5Jp
j2jScjvJWx3gaqRBBV4mqVcLMhcciUmLIQItTZYPTy/AiHYsW4c+JE5o3hyk3c4j2kh5QAIeTnNk
pVTOzDw4M9p3iE1+xSjqehSszoEHuzqbx09uGrX3By5jJIM2b3cxrHM6epgiUf2xLeQY8/BAVUqe
3r1keJA1igEwTI0xxNlf0EilKPBHV9l8K2gn/mid+xoW7d0rNAIJKxdojxsUDb+DO2hKPydHtrzA
eRPvSaWCsTBPQIUYl/UCHre/bDBJLkRUKAui9AjwEmCnG7lGNcBwvNVWEugyQvZgK78ZaS8muwrQ
U124yF2Y/MWnWtmDWzdo31FVxdIhQ/anZ2I4nwsAzHBjgq+B8L39TwNfdSOsOJuT0LPNbLC+2hb3
SxTSUgi/p0xGe9sKXNIQMa1Znuq8KpxrvFr8h2Ovgezve39Xi2gQnQykWeRPcjYZxOp2RWoD35eo
akWU9fjizw1ePdG0VDzagVQ40LdreCH/ci8KWtRgFIEhxbuZkTY7L7dmDnLQ5TMioT8bbK8+nBxN
hKb/mVXF+/4xHYzPH167EKv/DDC5vyjvP/smxkmuylCmaC4LLy5/Q2jurLAwFzFAtmMlLbVdlJbj
CSavlkyroki17vWRol7i2/5lWgXsTCqQhaMUn91qq7ULb4ZkfT3H9JobsmxPydmZvLWrv99W728O
vkX7Q0DJBuQcDX+NBMh+EgQsdKGt5C/Vbb5NMtkhs+D2El8DVNtbREQIkRTQdwiOTyMDOVRZ61bM
pFyVMDms0k0vbykUjVlfW7miGdqMSg/JiOfUEUX1YlvO2wh7nZXtfQohX/81y5EqQLkUpGhUsE/V
9orGF4nrW7GwS30wYNM7B5aj/rCNMPG5pG1H2qXasCcL5dCLOYnqzGZ5CdqLtYvLsoJHb5ovrMq3
9q3VqNCGViT140quJLBfqUbL3b0qKcw9M0Gkeuk0hnGnTBSZj3oQmpNwyjh4pOiUeR/e7nUTgLM5
6TKbQ/h3g3S0RcYX1UoaMkMSHG5ASQwB+lmnLZF/gQZRE/dLSvFOtgxY1bN77Y8m3VyaWD8fcX5N
F+1PUJiaFqJ9zuuiM7ev0Iw3O0y9veodcHgj7CZgtZCAu13ZerpF4riif4GskTIrw+rBkaIGz/qV
witBWzlqUrPQiQQcx56hVUnvTVTLrcA0qPX1NhQ9tR1JaXuTIk6m1Lf6fhKTAw5IIltCJ3E9LMgd
FlztVJujBZj2zgY2BPRQlhVfoEWlpglUx+tEflX8ka6zCM9lMtyz4ee1r8jLjVaZTTm1eekR+gcV
Ooeehfsrl9tDzDsgY4V/jpjW4TyhmQ1q3wIeQyjWCOhQWC5L/R9BIXw88v7OgVj2IlT23hwFs3XU
tsE/GGWM6UtXBM7heYyow6Cp7ylEK4RjR7ZQiLjoDVywa5WbaBbGtD7Jle7ttwNSNJsOzaoWYigU
xlXjA0TjaQVRzqFmhrh58i+BAHXjwD/9OLF3LPSvIvZmpIiOoQXkazrzbjDu9JCZVSVWSqoQ1CMy
AIgq0uXj+auCYdD/upCPR6OHlFMlMEtGHyM1Hec5skTcmrEJKHzU4GVpOvqxJv6T2ZWBdaSi8k70
5ztqY7hZlqtN3ZQCpjV4nAhCRw80kTSu4P+FREpuxnXsEDCpxwWPRyABmWiNN6CWlmk9FZu2+brE
LkNbHsGvo+8IGQP1eiG9JE2Tw9kOasKMx7MFVR7CyljggreU3ahrcn4zfHpvssUiQh3PaUMWxpes
LZG+F3fJPU+IHntOBC832DKaXN7otQBb0JLy9tsGKZWadP+U6gRMlcuxGsvRDkbOu0/ANfvGIwHj
JiRXwl6i5n2JwggZzNPHcUFgjhWL5+2Ew5cglVl8NWvW9FjJJSoYyrF6wUI/zkiw47hcyB6YtbCb
MxuqcVySl4bikgN7i7KnWMHwsMRp7d0jlE1gYJHs676Ost20erY3izJvqRYG1Up5/acsZnCYew6G
TGLLa9lTfyxU8zhdz1eSHQ/YdPeoO4V75tvufqbM12mgi2g0Y7dFgT5PJ5bwJ8gD3Yks6HkMg40j
7Cazy5ZRQSEXjQ0HvIZSv+nhI43JVu8+GswBohPJVB+mgWUVq5TBrA4TtG+kG2Lz16cNsJUDJ3eR
A0F2vu/yF3F1DVKxioU6esmkPAshjL5bQIpnHOAFEwKC+cTI0RtgNLHEml6YOnipjZ0huMnXe2gs
EGU0ssYTjAN9CwLHtzyaChAFYGulnvEKjINdAwd7wyb12yDjYKuqLL9PUHLHkwAL+tp2fJMmfAW7
gB9owWNkILy1JjWOTR0zSFiWcqjKuiKiYRb3OC6Y38GzPTUkd8H7wA/UkEJHKBC4wG7ks+QCCbGL
WzPKvbVi0riks9lG/Y7wAi3OrgYUKTfav6Mt0eb8hDQZXBK9valzTI7YK0KwbUr+1aws4mt9QMn9
CBazv2VNcFudEOiZvZ19MZxffi3z1I+pQUmig9sihBRNCsE9PUGQBuqs2r8iHGVm6s5yJnknOYId
caYtoZgfF44CkFbtFSrDmi3PT9MNLfy/G3W4RctZECI3vyVYgtgABNDsJ++t9IJyzT7eYw9HKNXr
tRNiEZjIpYlLUdCXb+tGiS8uPvW4W3WsC1GriG8sD5kybLubkW7n+8GDkBJNyZvqBvuSAx9T8tGu
wRlccR6SH7lTE8LGDXho76ngZ+G9sw8Ibno1LSplK1pZ6UuZBPHHFnVtngvVUrsTg3kwH4LcTRXW
4ztoM7kIiWMlaCPxAYXYJWJBjo1ssCVFGBW32LGdwWN/NY4O6X01md50Du096xz9vbU+eL3Ynu+y
QaPfwy9+++6eDMjKnRuXGsmlSDioqOyueD8wmR5Vw1NxYD+S27OzJ1hfRoWMok8e37zflEan1YjJ
qzvyiDlzjub2ETEMZoRM/eCbhjK533FmSZduB9AHuu8n29qXblLXfCZNEo4aZ+9gPrqsSyOS8XZJ
V2YxABqkI6jtiiIGauc1oKXjxeS/myC1gMY23GKw9CFT8P8WBakUh+ac2MzMajHNyrdxR/nl2jQi
k5wgYh+J4hoJRl2i9VaKaXBtVNewF+lgIUseZgKnznVqMYESzD9F2Yfl2T85uFQXn5d3VIBACQHH
53Vt45qn/XZbwYDCdyD0JLbierVI+GZZfNaoGbm2U/4HRZHArXx+EV3TG5EQApslbElupcHPV6kh
e6Eqab4YbWTqeDwVzUW1kpvM+T5ouQqFHEWlNIJG3chqcGisL/eW88BOpj0ritwiA8L/OqpmFACB
hwpWCzNGNOiNDlabC7n3XAmCFO9OsxsnNVu5AzHjYU8M7x25izmleAZNSRb/Kij6sl6fUXGlK8nP
3tiw6tTNYWD1U+tPcM/1VutLsELeF3b3P/W/2lwiTrAVD6yBa2/cSJe0K1vhZZOYtXEdWaJi+0FX
THtl8YDYC/1MxwOpK7zJ7DvmK/gehb+t9LFpGqtaSvYx5mahC/WiAVejL787ZiKprIPUDZdMjK99
Hyt3v9rW9tNmfw+ICbIzA+rHNiI33LtWeJPz1wNpxeFJA/h7NiZUf2S1bElh9m4PP32IxIhBIrKM
BiaUbcWcqUnFR22mT3rxYdpwythzgkRRr48vneJAkKtV4Rc90JTLsYrh1VJcbtyqMoEjsOecml8z
KEYu22EPPoioXGnDVwgVG6G4j3rVd4mNxeNGjxVUqwivmgHDaf+yIhKU7VVGo6Ilr0EA2fw5xIq9
pYDnxxI0vsxHgKKF7GLq8dbUUMU+6Ber2GUMUdDiFTkhlfPQVjJlLTJUM69UsbI2c06OiXDopIs9
eTB9EUttDsAZ1YeRsl2kILz//hvQliJB9E3rW5+rWoLSAWoKVTVyAtZychYI4YoTZOL5uESWCf0X
XQOHGZqxJqzB6PK/lMUKdfBHsO2A2UKDLWlp80NpgNLkwbY0i++x/Fh37ouUJg2fi/EsZKR03dM2
Is7infpfZFob32DSq7Nw0y0rhaRZk6HTjYi5M5p1uZERS1vrhUSV/b49xIYJzXs4xOFbqT4FOVNi
V5e9eTwgNm38cZex5sGZdMv8ucvC3wbkals8ZSYV6WB4X/gu4/AFVWzXE7t1UAVbrpKrDsDCu4at
RR2/fI8sq3OAXNGugSSmUTySaWA2/IMmi60gdIYGRbHJKWSjq/iyIjLJpr3X75NYH/Gwcb2yJx59
pbkFeLrFDEID7irZx8TCQjRBKOHaNS0LYK9E/9Sgo/QjjCmv8JTrBjLXvJWZrj+raTlkWrQSBHPc
Q2MA4bXF+iMy/ibmsMuh8wWdqBvt3j68kPTGEeIxFVNV51intxAH5C24sktLc02GJuT0NFSJGGEa
m06AZTcmdTnXNL2g+cvGrKG6h4UsbpwlimqIBG4TZ1nxCmVh9RLCCIVgSHbBepoV265d/hnuNdqU
0SYZf62R5gAlyuewURk5tEiWVe+jY/1oW6hnOlcJFMV0/PHkIJELZzLa829KBz3LMh90pUq+EfAz
WoCmZF+7uhdmedrB4jIHs6d7+YSGIi2C8kEXsbbwXSEP9dnxSjJOOOoCW3ZEii+QOezLpCQqtVD3
Agyni6Vbnoq9xhcEksKawlOv/eDoQm8nYaeg5lzVpnFt4HYxVbHYIXd+5thprhmMDio5zIGvwBfx
6cvgzvBzRCyldHxG03BztHlxOev5shj/yxDzFFVk+OvKj/bYPhDJdPtocES1OG688dpxyyW98SmB
XkknUm46ygDgORsls20oe8ch85CZpXFuzSGHFhcC1ud44pL/gAv8l9mQ9LmfKZy93Yri5K3yWZhG
fCakF64p/mc7FYm3GMhCnBbKtMmNQjo5/wClGoMeQETFe3+lLIzj7zNYWgu6U+olm9e6yL0sJ/eO
3/UBQisy2F37q4rZ7XA0BJ7GmFoym4kSQqQw/pSuoxJneaptJyitj/3riewQx99byaJTiwAI3/u2
IZ/3IaqLMVnHXIq+dCNSEgJJKyCyWoBwf/qgaRBn5vTeuYwiYFVsM1RWRyPhNWYTDEeDGovcKKjX
v26HBEFl/V+mqeSPid/TD8t9813ZILvMslTsPXuw4DmZrqXSvPOxLaeHPmy4M0LFaH5OKfuwYCED
9xcuYDGb1GaAQmZ6kiYM1sjIYDi1FEGwsFeOl8/6zSJAr72axdSWirjRtE0MbKhe8fZpzuxHs/t8
Vpw891KWHMTjbto+nRy9s1rWEZrdZ8G/aabSfJdeYqBovau5oxYQgjdc04Er3UgNnVPqTq2MWEpP
m2JZxnDbe4OM6nz5Esg+F+wosT/qwwT/IRvbFq4UmlLEZVe2ycLe+3qH8ZwMshMlp3IuQuQ6n8Kk
zjBNrSEndG4iN9xCRqEF0NjYMYl9RfbtcQsZWwDDNji8ZpyIpN7180aDBMjaRWavxuoVCFl4edDt
gkM+DgeNiHnGkRQycPd5FTRORRMzBr1TjUBoAjbsOYjeRm/2ZlqWNVfll6Fu2Y85G5GZbflZimwR
UFkd1ysh+i8212axQ5ly6T4KT6uSUHlaBGPd/6BLgGsRZ9i4O1482ObNFT9S7/cTcx3lSS94a3y/
MGqUwwTsAQdL6dGP1NIvTalYx3/cJaMr2gHoAcrSKH6r5S+7Ip3XHAIRN0CBJg7M7TGD/y7NSe5y
2AikUhCVBK9TUw3qWZlt21gMAMw8A6n+1K7D2vMzolPaX147mFMe3jHJ/22ZrdUDQ3kCi5hnClRv
juaBH2h9qvSs3omAMr4W0ldX2iZEoSL1j470IivkXaFv1n/O3yXp8Xftut/2rWdEkBZpEhN1BfPj
9zuQydU94p4RPqeeMMpfPYAyYS6J68esN420XSfId7eowqrOGbiZgqYCIMXYZuJMix7g12ptmz9n
A2hxWAbhW7OJ2DPZDm6mfxdRoHHf+K4R4pIHtqwPradpLoaQtFyIEiftdfyJFZL2IcWz2xDdzFsd
Rcf4vSlmCTzxpi5asEhgqKXgNOtexwo+fKb1x5EMcykZ8jnxHkSsSMArG0XqLjpMAWMsNDW8RjaK
DCRAF/3KRwu37KXSFgotFMCR2w1yXm26SrJ7BfZmqoSeXxZ1uVUMV65g9nrRKetEdq/h8l7IQEEb
afmDPjgJO/6g0Yp6b0BwnQqk1CTOa3gDsMDsdKhLhlQDE94nYchAEgS0yeHiD88IOIArEFk4UpUI
y1FCVBRx+Z/QDg+bkUPtCipOiJLWqMxeILXnMDYWadbkaEBOS9JvyIZVkWoNidYCPVEAhfdsyTLZ
0xqmx9NFm8xg4kZLQI6CYdb4hXjc7eldU0CuM1po9kwbnwn+Y2PnaJQj/hKS7pAQQe0OHniYChpb
Ltaz4mgMMj+aZuHrvDpnxBydzoQtwWL29mNrEobSnViKm/ybzli18nh9l56LoGh/giAwmo/sQSel
Ftq6BJMza1ur1bcTm0oUPzNjPIKm5jyXUtmKguKY2p4k5q3rYr1F1+PcMnuCKzTDl3nafDgI9TIY
JVjoPYqYM7w4Cmxu4rWm7qIXxAxyqNiV3JITLN/Ak0W6UiZrXWlaC2GoAffpsUW1SPdRBNkONQEa
8OYhzLDIWGJwHQU9QtWTfUJuzbhKSnCxMI1p1kvM9zsV0aYBBfPhHIynWAbN33E9kAGtitAvWrlh
RzxLxPmHQrpr/2DoDLlMaaOz+0d1t5wipYdMIjTNZGC8ScPCqDGOpA4OdrbYGQkceJtJ3kR8G3UK
qhllre+kfc1u9IR69mwBBBZoxeY9UEdyoxxpzsKujpKlged2EXptFZYrOrWantyQkUP+Bo3TkAVH
nddk53nrdBU4Z+53clEUC8wFh4RUVT514UOmNKDuqTymcuanMHbw44F1LIl4jUyaqRy8aIHHZMtu
W5SIpQMrm946fPV7V4pxU4Y3QPIrGVL9SDEi5NGt4ibCJyn9EkWkSCyBVPfKXxNRxYIuKHQdBN/k
MM+NbygijBGRr7llGhLHitGJCIwvZ2v38pqvSyyiQdR0W7PG5m0whEmuQVFbql4C7LMaIgFrSZlG
kgXKaURnmMV8sYrFd16f2evCdfLSG0ttwxEneC/Wd7flvlqrjJkmPd3dyTUuK8rqywWSLDDknv3Q
F/nHFpRxdO+kF0USd4+W37CCKgtd08OpOjfHgHSnw99SGJjvUuwZ8Ygpz4gv0j5sQinHc62Mgth9
lI1doKJVLTrCDtnKXOMC/JFJ8cVygHY3kRk5ihBDV8RNqcrBSLJBZUrHn2K7YZxuwq06uqMlF+Qs
uujFsjYgK79GRmr0MQMT8nlnWMx0tfhltJiqr9Gi2mHoDZONk3DR9aFcts3nDPXf47LBJqaVkkvq
DmJV11i24QmYZTScEUrK62TiOlrNosIalu537Iea0iRUgepS51YdC8x+zG7r9QwtzYIBrJ+3w5nl
qWoBclVmrGYvxjtGsGKSC/V3dhNsRN4AzeujvSMaDFGXym+2FjPqOz15iQEaaFTerw4Wbg6gwJc0
uuvHMUd9JKvceoAzKBAG6jC7LLde14CZqYikJCyMrYYcFN0ftQlc35xRgXTwwBiHQ6qVeadcS+85
1tIfjWujVRIxvU5Emg2knAd0zn/Cy1Wm0+9fe40IiSnx3G2Eo3tgzIwbBMtpcRIHNVIzTxKnT9n4
7NxQPHkmdomOWuzptGVTxFpu83Xfn/+g3Bar6K6qoLg0MhNKhZB9b+Cpb02J5oNm7XSA9npPGSzJ
o9risUWvvDgpPxCKqpZyN+BkJw7oWOwYguL6Rw9P+4miUn81QKxtCDaBlL/IFx/COWz4MXo4pADy
x8B7DPNRte4v/9urNH/9u7v388uWRa5Ck19ud6RFCjEfMYE1C07QvE6UuETdV1ox779PNyZbhjaP
bIfMLOX77TNWAFnehHOxmZiYnjAGrmkDTDyVc2yodSTFCFMII+Clv85TtPcnZd5GPJwmPxEF3o0u
cTx6xCUHBlhBrUvlR5ARAZqNCOWS3ppVkS5N/wUfsGdtCmtUE1KcDonbJ5O5vrzWmSxudSp0nYC6
ZD8uz8VmEFSUrDrFltteZsvPKMc7YhvINvt+tnL3/veifI45ShaMUHCvtRcdgkvaY1BlKoTRNaS5
NAcwEbqT3ZQQSRNSszOoEivLpYW2MNXnDkHY5z5PYOjz/k6l/Ic6vYpCl4wtC++Gga6sAkaf+kRX
7dUl8CaIWmmHGbpo3yMHokVaawezRwc3+4IQ2B6n/x7sLiKGKg2/daQMlNJIfG5GJURgJxiAjb7x
YW17NYZFMTPejXYkXmgPW7JT26GpXaS45pWa3b3bhpfDtDReHR69Adhv6sxEK/SNMf4wYUCnCblk
eZy+t1F0zlLetRwMi+tc9MOBoWtggRB1j3x2/vR69cf+WOxoH3a6BGZRiGma2uUcs0YLl5KCZQOt
KdWsPtSpvdae7yfbE2+tTEIPj/FrMAlR4+dcv6P03UsNLppUi7aVHmBT0JM7cYsfPb83RSESrWNl
RpiJBFr8ay2tAMCrEDF2semrdwWg6jL1AJwGMEFsxP10h81FBTmagQw5emF5ve3UR8IOqjkFXzZC
UPhdVMfIXnD1jI1ILSkSrICU+uBtfLpswCXPM0D4qSLTloy7v4xN1fXwHskwa2ZfP3GySbLi0Vee
jPSHO4+UzDBXZXDM5nK03b198QqXz3imumfIBl9+69RKYfKRGYRLd0ueFRyT1kKExygpj4WzHm/C
2ANl2KzSFzfll1A9s9cNki8ovGaJfYGMGmMNShut8iayu6lhAg2cUKmaGwwtGVRepEZWAYokzaYr
oV6DcaSFCA5tU3D2JQrrfb384rnGjtuAAB2Hsp3nNdFnae+IoWjF23JE+Igyh/Hj+2iqBu6WxROF
gAgeHu28MFeFpQXWmeoXq0w5RCKhgOdq3WaOZw9tP8IiMxR7qVJooyTIdUm7V8gv9bYTgJ3bTpyF
IuQZVWruOjIc9HpFrY4RDWISDPb7HbOjwqzMLZadH3cTkLOlDvixsZgHNrVM8BDi1o4j+1PaAi9q
jTDQSZfxv/tQxhN+u8GIZhaZozfx5iiLVCCV8kh2qqXgvg2O820rZgW95DMAebJ5eLsW6eG2Inhe
/kvXUN7sdL7HD3FXhLBUZH7eJmXYzBJ122abxD3nzoFPgGPTPBnyazIO2SThJheclSddQyhqsePK
/fpqIAwEyf+rpJw5va10vJDzC23jF2KtOOnFySG6ekpHaHdqlJCEUSedebb5YoOytXy+tf6FoD6I
jcbjfSV6ObYogUnvxzWQDtn2ZRfms/OaVRCXh5iISTSbKMDUPJeyzvT1TmdMeAxT20qas4oKSO4X
BqhbkR+fQaZL7brdOabJ3cQN0ZTdU29JVQcxSvRLFAM3kH018FplCHnHGWNWb+NUvzv/qm6JjXK+
DwCqFAY2md8GNLA/DpHCVmiryIMxcIvOQxmYuJm0h+Z3V+TGGgm7SKvDtWNqD3jXHHARRLWCE1Dd
ksF/vC3XpwL8+E/gO6riDQLhi5VUY1smSSaLvqLEBSuHNzRuWslcLrTMHyFAje5ZCe09Hyu+isEv
4m7BDsQYi2hl++8rYmsfboWfU0BXyWlRJeInrhyMZczfC6IaXzONsP1IODmUfuzIpYOqB2dVCXIs
YanssQloEybeUq5Rex4UK5HoOcInZC0dcslBeQaa1l+mVraGm4vPQO1ccD5yW6E13HskG5P0ikn9
5TjCigVrrGk1XJD28Nk1kAyZPKpqMVfhOCkO5o9cbVVUjCgUPVV2GcY3NEKnRkOY6P7MhNiKmUrK
a4A3eUkehJMRO+Hc/kGgBoie9gXWk3cYpBVPfdIsl6YPs+O6B4W+HFiz9ytH9WdIyp2Ghhlmdk4B
cEdtpYJjUxskqoIe/F+XVukRaFbMQaQM1tMzvbotFE2VhgdV0hvKxjog68HYDnom/JKvMyZkn97p
2I4tnQj9Axk4fKeTlUhpqHLnYS7dIq83nuw5rJUyAPkl+vCYiUZkL8wMVGqttQqwmmbsQuYw6Fvx
7YeEu3sueT5P1PTF51ICZfh/4N+vTMb1V6vZY8Mp1fcJoi8TlIQXKiEDhBiiA5rcvkeD57HZi0/h
yONVx4lEuUL4F8HCYsrxqX1RYt8E+qXXBpCwnZj8hICIwwCM05kd0oIKAww6AXo2aKxnIpinLD+7
fAnGFidns+uRDWnYuI/us9yOp6ITrNlSiM52kh1R1HlIv0It9NcPglbdAegbInMHsOB1gBTfkc51
1LBaDe8EI9CC4ACBtyG+XNnhS0Xfy3iJt+qjK32K69kSmtzwLeIsVFQb/UU4E95tTe6Y+FKVWLQA
nWMXqRCsDCJyJRBzDzRvrbfAwacebY3IFY2+P9M8znYXski/UEa7sn6BZmBSHipAi4wclXdcpFeK
8kFAWqmxXGKFkOrgSmoq5ZvlXajX0Tn8imBlTlYaKqHdVHxCu9c4LAWwDrFh139CNBeEvodVpkny
eo6zWG6dRQzSzO4s7d1BB3J1NPnIPeDMbkOXP2JOimucyzTlv8wHscoZJdTCgeylZryG53xIQ5Vc
ocUCtd1AgXjhjF8f2W75VCEmIej+gKcdw9tvck+bGCbbSlpm0y26CXUVbAnXuP4TYrQHImTaZ0k+
vMUdBcUUOoJjflSMSbZhQQ+x5nq+pEvHUiZoxiQsd2Y15rdSk+P2CdW/QgVYjAUVNyYmNZqZp9PW
gez9vGGImVr8z47PSC1rS1WWiWf1NppjD0p59xOl5UOwx6vSQhlWR/ZEQe7Ch1UGdfCfS3ry/PqU
q3rbrgWakQhwLd9jZD1iVS8PdK6F66gxQwxEZVcW2ZWwlLPfAMXLK52D+RzZQrSegXn7xXfYI5wm
wk32N4yPfsuJF8cZNgZtrvYT8axROemk+JeSQ6Ow/aFY8A0reDaIM9HVCiQVkX8qu5+krJ25Ja97
+C7NsgiWSff7Q6+YC+HyC4y6IpKUcv+YQv+1bg+lvJl99kWZcxUGmndQXFd0yaZbyLusMy7o9YNu
GCqpolGZxBs8TiRFZjJZuqsSwgaWbXnwjm5Vy+zTNWrNqSAVycEghypbK7z0W8hqN1Dxa1IPibee
Gjw7QGyLi71ioVEO1MA24ZXp++V4pAdOb4GakUmKchzSJzIm9pcDKb80GLH61QvH8Bq2f9YlV67i
ibImBpp1IHQnMi0otzVyYES9JkLXYLzrdavyD8r9rBr0Dph/Hzax/W4o0y+BBSJ6i6hYqsqAmMo6
pflT+CuBVStP+RdX1g59bOUci1JItfvfrHGp0wcFGNEQKU/WBZDhe8OPu2B8TXg0ylRLZQpu87LM
GBHij2QpXiqscRGDiYZBc8i9QSMCk5kC7/WVzUIYwMLqEyU4Fqj1PY1rXX8IOb8Uas+5kH4IrJmS
zVJiwW1cNEalIZ2YD+IsA8krOR5MFod04kdnzg7KqclpWk9uUuzLtMr/6FGmaGcNxN5CNKKZufih
yGBBSUoYUxR+sTOq6DsaRSOH2NO8AB/Bbh/MQQ75rGJtYOjYx28c/YEpn4rsWB3g1LmXwB4/7FPz
XcaxRdrXqmys1jAT/AjFna/wn/YSqn+p5WkqAFOK0ignuvS26h4FBimpth4IFVlMzjiDaCQx7hqZ
FzpAMLW90EL9662rDPdMv3D46PbUwYSV3y1F+FrnetOPOVasDXJ1gAXymsjN01ld2Yu45QP8ijzz
m4yNlGBepYBU68PXe/lDsN2NVf0lz/pkYTI6huOiYyaK24TzgrUz2kjiymsEmokbgreJqu+j/A7j
IkFgWWwE23QK9Kl9//IBn/TLzZQ8SS3qogSDwyNlJSmcnKkhcutZLjFd0oSf6tw84cQI32J/nP4e
eun9WwvYEnN1KLASjk+xyNJDPb9knOIwCXcVQrchUSBkhAtdVXysT6DVDx9PBTCERdDSagZuiD+3
qXGmWEEX2hlg3sBCuAFsH63rmLuLUdgZYQFWFGzS0UWosRNyfYotQ1KL/Wk2g2uogS01oii1ryRm
Tx4loJDY0ASNkNNp2IFr8aEcYDVkuSBqXfCxgJVwi9C/DLvRBGXCN0Svt3NdLNnSL/pZX+aMXS9b
zbfD0vswgDtoyEhwMwuItG5NYg3GzI8ZwAyGvO+C6qFJkz1yZHWHgenzpWsRH7qfGde9BWuxJRWf
dyNf4mk5+UNYpsj7QJu9gXENjYnsv/KibKfS5BJhyVMgwjFxgFcE2Hg34FBmKK1FfoSAi7OprzOW
8sc/bp83vuxo9fuxjQ7Fu+1KZY9XiMxFcCU1yGRhIWhZtCTLDZz+/OkWzCYmWYEmrCRNcMHlOvFu
75FeRmy7NFgBO5tkL+Z+o3Lxefg7sfTdCVVaX9M/eEzI9npXLc5braaPV1tXepAUONxNABhgxVnF
nJxyMrN9H9xvXbEl5BO3iUgCDYCGcd5aMj5vgU8NZtnh8ZA0pJkxedtEgoJe8BqjLyjC4qhHlr0h
8Ig5DKoBHZtipH0ndxXBAqA1tenvNsOGbNH98NU7yoxzW0d8AxZFdnqVy5AqVKRhKgHw5upkjJb8
jVCBEVOUG9JT3VYmio8liqCY5gK7jlziBmPRNNVmJlrRvhhGJTwXgeUYX/Unzs1djO+/jr3KZckS
v4qhQDrzjzyijduHNBRTOM3XC7QhCHHVyXGlqqqdojeLWrae6czwWA//0vOLbZhG40Sj8C674JOU
doH0GozvLAmfSr2WNFPfLkaq/tVqtL297Z4rehFJaftZWL0mkQdpUZFd0WearpdAfl31eiq8U0Qt
1By/lGmicblHnnsSqW39DLhhOgWvRHt0MH43z8aapZGfXgLFSiN8WcxniR2bQE8/635EajAnj+mn
CMMULBxzlrxQJ8d4WaLmfIbVdpVCwOE/FQCDlvx69+4YmbzPKS60x4LJiENtyi+r4vsGig0Owbia
F1bI82xaDMPNEqeggDiQ1R5sflCEfWz3v9tyHH3eUlJwvM1aGNXqcoty9bt4n+jd8Q8BEz5EBePT
+3f3d2eVNUVQVPJ8esI47W+ap+OSIMKOEAy1LGMpJLOVSdBcDJ5qlG8KzutkbUL02zQGSq7137ej
r0a40UDvrRsWbOVFWzSxWamJ14ma3m88Ip+e2xJo+FBhyjj2Z34g41OH/BjvcxyUlEoW8LljQan8
7b9t6sM6X+952XmZW4W+GLd7BN/TJvnKv5k1n5jksr97S1M5QPsyB71G7Qe4429FNJm3OdJHjsvF
Yl9phakRG6CprRI4CJ96csXpmoW0Gf6qGRCbsT9xPXskUaOO6aLjMBx9Dvz3XwULadDROBbRJyCE
8ToMW3aQyAgI2PJqYtOxdinBTiIAmRKGkikvT2KsZ+2CSGQQCKyVhh4LcjyJRFfTvZW+7Ob+cok5
t9fCHhvCPFxUChlWmUuecR5NDGcmjHHF0DgD778aQ+xwoGVTxUfsC3wSoI9mUfHPLkM0XMSyx/VN
Jce6dlQFPm4MHv+Zn4SHDo55MB/RrioMItXsxVBraZJ80h/4D/ZEfKONJxh4+zY6ecGwiTA2QQyQ
bNDsbNzku7xjQX0Q1h/OOclAI0icbDCGYT7HZps2/YzZdmcHVyIqpmvngQbp+/+qZgzSANyHeNpu
jBnG4epKUXHEICKa8gbBcRGnKPOpYoaZSWJMMsfSfX0sdiupb5yknSLBLgZcO/eTN+SQwxSQV22W
3tnrQlNCmsER/2N4reYi1CTDhvWz5gts0Dkg5AUeXpA1+mV9ZBHx+6rKsgPRp2K9FAmLzXNkgS3I
2ObwlwjY05qrz+nF7E52pSCMKSgSmYfsSn2QAETUkmInXh0Fbn53H6B9YYx7vgN9k518xoa1jT0s
pbAR9jQNgSjpveCwPe9OCSe1/bdwnQxzTY7DSlIlFqVGrCxpMr2GUXE9ygr7Z2PKWQqChUb3o9Ku
KQTlTdXJnI5gRQGtK3a+a27lGyxn5wE2GUZm6CH8ELmuSyeeETCrD1jVySNYwH1DGbXsJsGSESBJ
Pz/q2WkH+USlinp9QEqo1poXM49/7qMS5b/8KByPLgpj3goHgTvxY8pnO7aUyWxCJRSxSRHNBnS5
BWaGtyflWv4iSLBghAop+JRt7wr50uFERO0Jpko/S64GowPDbOOFpxEEFWci+dEgg1uPzSF5Yynw
ccH20QNZwkLMqWdRisQC1hu8QCsPeaBUbj5QKwc7W097q6DOjp5Pk+ZHYQdHvBMzMpCYmPRqEYO2
V7bOcp1FjJrWtSLNdri3WtVQ7B8YUMjlnGbzKvHQnoKxRRKTkrrUZaO0rGfCuqUa3O/SDEgSgtAz
1Qj8ZoR4NB60nZXpxSKJQJNMhxYF3hbN0DpPeqgW1/9Vx4yf8oLN9V6b83/pqk5dYC41G30DtqAM
r2f9mNRwsSzmzUTpY3qZuqi0fIFLihOl33DS5Xrm9sO9C5I0JY+7ifzCWyE5RyMOqtq0d4eHZGpX
mKI5y9JFIPg65MRJ2xemnCRBRkNhuseYE+bMCVFqotOXrDuzrbEh7JbR5NzsNBLPEIGcvdJiQccF
dBRHHqHsgzCSMl8t3Q9UpFsRcxdkdat2rypp04oOcDBfCfmx5o3Vr7ueI+7OgYRfOUrNBLv+MouO
ZEOPKsIfPIHOdT70YJhF+e7zPzNNp0tw7yolr1nhlwGaiPivss3Ic7/iK+FJiBVNsaTzdugPUfPh
mNHd1Sc+vDEYTgcyLUfRjY8gfR++HWx1+8LLG7oYeWGV3UkgGc7qc4vOqkAXbAURoY9aVjNh9UzS
C3AiNTOcISUT4SMZbgeyEmCfEXEIs1AFKKTUjeyWhmfb5eEixXdG3RHNy0icj45twz17BASrZc9s
s4Fpm/SJw76p+cVYS/UY7uch2EDspE8x1p8Mqw/prWzvuonht6JQDFf9XnSoY7jhS9ZFnxmS8AOC
KqPiw7nmCYwPn4eWl9COLCjdczi325VjxuazPWG/UUdWLrV8tNYZUhw2m90Mft+rAIzeAaI8CmRd
d12bYfb8ukPv3XrYQm+7QM2M3cuzvW7XJM7uPmX5nffWd8duydVcxVCFODJIQzyhBCScD6ygFyps
nnjeI8EVLIxC9pDZQtpAYL2aY4avmEDjMr9vZnWAowvENxCt84DXL6tW7pV08TKmBj0++p2oxH/u
r10M7BcgCE3ykfDXvqgc5THxkmIQd9GNxyp8nNUWUspWujvkdkQTXGDeJRc/HsbkgIsD+mzbxlR/
vXOynWghMYVw8N/zIbKJ3qAgggYXBkvkXWyTBYYHdMt+lE/HfJZm6ECe6kR9y6XI9GZUJziYmplt
lRtlO487+yD3vSxpTvj1xtbYn6BOZzReSlbHn9GRR9H2kUrvYhFlqoibmBlgpj70yMEAAslSYV8U
s7+bkPotFoupuqftsvm5Z9ybSgjIulr2GY/5ONQukgxzyniZYDhdBmRfbNciw2NlNLenXKLv0+Ha
deVPZjZpede2BWzZNbrOpezcOGy92QFFpowTnEFGxbjZ/nRpSyVLjDJOtxQR+vn1oXjF+K3SRpQu
GDOHrpMqk7JO5Cj9xzyizZml/G/aVpv3N3sJCRhePV0wEkUVFZmPxM45q8yRdeGtbNyPNwV9ylrP
5aNKi+hjfYgcKvYVExasZiXimoZtizwHpq0tTmDGLZvYzRZGgic3HdqU4v88G0t9b+7muzoXGlNI
P4Z9ej8fdWBkIqRVnIz8A17WLueMp2db3uNkoH8MYaDHjjjcogEv93jU/BEQCdK2klZiD4vYs0AQ
qn9osJajB5/ZJtXBCUZhv9gu6y82LW7ovoB3cjpw2yWdA8HP1CNu4N3Dul6morDauKGq/nMT1YbF
OMvZ1YXN5qbtjaYIkrDQEjsLXUulyH2Cx/AXmjPQimtRnN7Gfm8BsPM7+Plf/VmAWCmmXZwTElbx
RWmzHxPbzoghJIEn1IAZMvE82COjAv0auewlsLCPFtIWf+5SWTbGfvGpAwXtYdEk3O/r4wt3G4tB
4QO4zj6mBauGU8OE/V4wxGHr1twxVvIPXPsolmnfhiXqIhi9ikQvu0j+AgiDg1y2sADOgdbrlZ0z
HI/iG0BWk9oAs5wK6ymY6z3i+JpreQPjHfWnUx8JT7YkrrbHPbq+DBPFH+fjiJpifggYAXnjmwLv
1uo1aVXZArHDjN+apoIGQ5AQxWvchpBmQNyZx+juKKR7478uG9pJT7+7lzPAYhXZZKV8WGLhQ9qq
lKYqT2OQcDuGOvAJzF6K+1a93lXXhUU+IGfH07z30fsYle4jvL6kNbpPw9RAuB/+/Qw8nURiPagj
gVGxgf9iG5rfPiwpWSnzsvxqn0/yukeM0mCT50THPW3PC0jE1Dkuhbo1swnTYdky/l5CH4NYM3aE
w+oqSXiJeb6c1VYVtte84xs1NtrtjXZ90/lHwmNOz7zVYc8E/535UOdIeRDs0AUXtUJ0XkWOsPAp
VAKeXfVJBGG1mJ35QF8j+pwHBqhbrpepdacE5yzBbzL76vsh7eLiCY4oLM5ORN0ZizCFtb2WToUo
UnTIN74o3XkCta3dErZhYh52kUKuyZxOfIKEd0SYTmCnybh7HCKt0kH2quWZdrWgmSIM+0PziYOl
jgC1Ul2xcCH0DPVnqEZeiO/bhKNGdOWVBGctks7nZdAfNGW4NIKczIXzUAKTS+OjamfFIxFuuICN
eK/Xxdh23jXfElxprNTDKKH1MOXolpuHQZakgHPgyUyM3ndzv+fcJLxgWDSI8I9SAQuJdWCkv0xB
m4U+n4gOt4vZXfT3lGyui4POivCpoVAxpZSFYsYIr8Ky0mBy1Lf+2AbUo1b7/WND7yJ8XuYF+euj
Qe/CTWFIfUJgvtzVpSsOC3WvmC+CTZ/m9e1j/4vE5qcbyo2GPFMUgIfxViZn05I6oFcsYbkkj7ZW
Qi2xPOWZ9L2dyLtuQwo0SZbMyycAwKnyA2osm5P3u8UPKlX/tT9zNOKlBiOfVbf1zElxvvhZX34L
5ybR3kEr3rYAi5T3QXI3Y0TEDE3boBabdpO6M24mcDlj0UAXNoLfmvBKYEBT31RL2qCvIDvUos58
nZXBhzJpJ9gAg/mrTNZW/fkwrbrZSxT8repNL1SrH/QzPaE7xdIxZhEFdk9kGbqzGEAj+x0JwUQz
jN0pH1IFg0JiKzdd7Mm2kdE2qYvkWTHhFIOAt/kE173cHWP/GzdUDsmuTNw7Ljng4xsqxWsggmAH
LXuv9CKk/gQH/6P47DOHVM1MAkxn4KZOpvjsieN5+FLx0VIYwz6Xp/yzPH1Yp8DqNgiruL9331xT
4cBr3jGjV4JtnZciaJRhn2tD1QVbWTd4ZW5z1tPbG257PU1GOiofdb05D6UFN+AfW+6LAJER7at3
F7ZWdsW7Xv2soSziOwghHmbk/QCCyuDB/PiCZ8eeCVnW1k/uxNHO07VQiZ3aIo1N1Z6qivAhYnut
SK2rYusmPUnUiqn4dN6CZT7hm/fTEI47yGHZiujOtAJtW1WaUa2EFVLWGEPxg1fCpd529Nb81sHf
tlj5TRKQVuuPUYK44mX5DSN1MFBkpdlzuZqdiiIh9Wlud9YzYK+OhiYgULz0+jC3S2qB1ta5lrsD
CM0wVJf+HsUKYIu5aYGOnf46gDsuHdkFgiB4B/BfiBLEeHVyz+2Q7eqIomb5Wh0sojJFb0Ds+FTy
tGgWadE3iEUFyCR4u2WGIASfTMLoG7OxFOuP8hmyVmfVMJejoxaR1Ha3TYZ71rzdXOJVlCcn143U
yj25jFVomVdFmDFyasSU/hR7RsFkaHeJIyZuNcukiOI9WwiWpt2IRvl7Vz6bJu4g/jSt4wfYgMW/
AU7V2bX5Jj4P6hG5LUk5fvYElBWQb7DrGa/pg0IpMCG0HT2xzMClZYGDCHN8RaQTQ1P3jZCQ25Lh
DXm1j7irqoLFs3LyvcTlAOCj5AB2auEtLj9G2xgIWkn9hbYIFQ1H2WBCr8g6xr4kE+7R7dvKlFh4
vniFdpdZ2j2g6Y94QQPpEwM9NebEYejGDErPnPnoPMj5ym8Q0jeAA+y3Ce5kY5SUvZTs1EW75bfB
p5KVoQgu3hTFITYgwWCBe5pNFMDQueH9THMvGzP071GUqUPpwS+0DbxYOtZlmM6m34pjrZPIviTB
oAIrL08ZmdnID1UtkqVaJO2w17POjvDHGuj5O0bJHfG5y/YZC/O0qWzgzlLQjr7glENnOg3xtFzc
L7ErslnunYdNZATvjdESVbsbGKecQWE8Bln7d5nO6TK+nwDHgJK+rry2Ucvy7/8NZt181UkiGIoz
AiIsXSMcYjy49uyjb3vQA8RO6+f+6wXOB5I45I+52SzuvJ7ey3YZN/FqStW6d3/rZVoehctURYQk
uzf150OyWSV51WhKgsqpYee0ujduJF0rTqBRRnsB1iUjcL223x2PwCIugh1sSpsocVlUdiZJ4AEw
GG5eLthWzu+DG9XGv9S0kyB93JVsxRge2ijhec80Kp9TB75+BnVP2/5Nmqw6Sl3n5EwSRThjQUyA
OsXW5ZI9rCgcgfbRXo72Fhk/LN+wYEa7b8cZlYtDXj/NHiMHQh+qvWeQoHP5PsmRAnprMO3TqU66
4Dfb22k7be+icLHum5pks3167lNDVLiTAlK7bnaRytJPogt/EYxiPcxCWytL8CadCJabHiurz6yM
SD46EMhHMt4lc3fcJ8m+1+tK5IfmCLdji28GywJJENQClxPYGTAYVZEyiVUFeC5sSnpvjrg+4A8R
tz2RV9CXqkOSzkV/rCdlxkWBYUQxTFvt2uFwIkKDtr1QUkyDLO8JCDu7s3vTF8EuXX6ARl8UOSLU
2g3jItH93fPlGsyAlGkOLxr9DkPTFFc4pR5AvgOZ49QnpanfRUxjZNQNoj0TSV9HxsInmXjrhxAa
rUQgGoq3t8tVoOqpd7wBqijKE/Dml0S1wDgdf5IwPEM4+sKGqS409+/MJaAH/HIgfBOwnu+x9fPo
UxRfmV8oIf1NH2Lq+I/RuUVEYa8B9BBxBB9tgEz0PoamXDbEBkVO5xuhIvh9rA0rmwEKJjJ48Ra9
KRuDzuF/WvHpnyPYuWr//9LyIkOidI04yyGBmdsXVscvLe6+n1zR3bNdLS6v0OOSYRr94oQuAKIe
fdopFlVZkuivld85fmtMBrR9r0WSZQiNC34jkeGaDepb2gSzFFqvGx/IDO8Eztw8RVonCe7FZQfO
PLNUyc/elOTsnmf1CmVHjlUybDyu1HISj603nr/ketJr0rLi+1LVtE8rJLaYqc8rfSZ3ZVve+940
acxnNFyU3jydevkCEIvj6Jdnxmn+96b+YQHXGYBbYzAW5mcG3WeAx7P/HjUHL8iaVxeLfyzIALDf
STSSQbxARiRyQTfygcuhFwlGOCJ6vZvi25xHj3RhNX1xg47ufpE63ILa5dmoXEsSU2foIISK166L
uTGyzc8dbO4/lJR1zqmkxh4xe9CZ/JAcr3jKTlLd8DxzUuoK1bZO3NCTPAYBujhD6PgVIoa2KBJW
JiT3b0qX3C7YUEs/JHv/pRI6QobE/6/FQ2J8Rai2ENc6lsZ6Qc8tx8Q+wA0olKidTFRnkpOxPsBN
M1hk69rkZahAPso6iVakPdRoISdeXL5PRkBhshd7NvJlC5W/4IKmzvKa7hR7z1o9YFa0gJqI5l+3
yZJ3SWWdcWrbfwWQxHo3u/tTj397qMQc2d2Cm0U4ttsIMowe2WL21rO4kg+QIHOkvkY9t7yXY1HH
u0cV54hRUIs3bC5JgHiCBNLLO0u66ncTZ2w8tlWJvLtNJhK6RcE7pXrKMHczlv2aJ214UAW6jkgs
lQq5YX6QabwO32ookIjDrtI+mkKO7s4SBRPzUipGPo0RJtal05mtxR7HX9ubzm7Fwnxkdv3v5sqd
rbShUUTisMBiBDpK7P2gXDAzAE2avrZlhbTt3vYdOePgSn9luwIotB9/lvitWbW3dDWh0Q4qTds1
MfzFt+bjvuq+SnXAtkDVOR4fF5RzETij52da7hQSxIzot9pmD8MONfFJEs4z92d6xlHaLNhWT8AQ
nl9pONqSsCJKfeh2C9QKVJmZiubxAEQbX5lzOhpD1d2OGWqfcs0+/C8aDSx+rtW6T24SaEU/Nbj7
wSEbHczeQlZWgUY4bgRY0wGulam8uPWkYanCdu9BJhYJOn3VK0YJ7CaQx615aJVdSXDFGXaQHsr3
3LBtyn2Unmeys+TOlTHLZKIWE8JPYcf88Hp3bzrOh0zF6J+fh9hRmwUYX6ifSuSfU739CdAePJ7x
WojajU0lFd8Di9slcBRmOq16UXygO1nDRg5tk6uOGtobcCZpk7VqVngB8evijSeq/p++C3O2CbKe
XfMldZ9Ly19ONoLd596bMJ2SKQU0tXpLb1sM+/M+9uLZTQy96WHwQR8NWgIrBLOVKmj8Y6q2UQFN
3zuoTAwgYnsfuB6Z9caG/prAlK/ndRq7CDZkYkTBccBiR9s2sCxI2rkw8RB21jaT4NKYh7DvAlsz
i/Npb0UEnsDhf+fkzt0PzWyq0oorfNNzvOqpfhrl9FfgkwO4oUF0JVXBcOSDev06ihkbEFMWJwhA
F24teQpQ8nUfQDdAIUhHQiBG+1uOxX1sxZmwYjaysOaX9CXuMwm04LZ/t/ITeAhGOgWqFbxlOMs/
sTWLo0D9FrIqJl5L6s139r2QRlqCxiESH3tpG6KEoiRj+62NQ7cPun+V+jh6IuozbnWBo/yx8Hq9
xLdwt6To1iUqKKAZk0aGGReFT10P0lWL6UF9ZzAR0kJPH7Oml5LBmI/rP3FKt4niY/G32YHap+p4
i3qxzpBrKt1AqBx0a8uwF5J934Q4g/OSml28bxmSYASjcAxv7MFhLY3XMILat04zkKZ66G/SQlUA
JNP83xe+6SPXcRs0jH0xgUn7yEmVIWIe+AX2pqbkFNplnEXTGcFTWZd2+7cPk3spI5mC+GIZPpQ3
AHFDm9U7w3n/Q7bA5aHv6ZWoG4F1SOrmcRwQ6g8o3OnStlT8EXgKUH/Al2NWqA0UHLteGcw7CcNe
ZlS8jV2chphhPI10RkZgkdsiYMVmg1omyksPHTHWdjEQnW7o4f53fqkjHTeR8uWU60srq7SZQOQL
n/q5pSCf+0ZbRaKumBtQbWyPJaBDhcv8EmdFvpR1OGbLkr0C3vJQ16vHMGL/mNUiMzPoxbQZMWrR
lSmXvuafWAzoWJVnlo6OvkzMwN7nAsPYHGFRf0Dnj/xIKh/X39vK1G+pMS0qEJZktIeWm+/0oeUV
XPrF4cp7RJMUzjOgDRudDsVtdR+rDO8ydydxHjbsPH+1/OMSzytOMdUzddXKnmQ2cvfS0lQPDYOF
PrsxEWYPgAE4hMFDY5bADTUe1YLN//bCTPYFkRptsOkYTbLl8iJ9UsH1JhpoXfhH9atsOEQBdGOT
OnvlyyJUAjzubV6/DYsLJIngjv2qNA0Fwfe46Sp06kh5q5eMlUipGwrIrHmGB+4a042eGUjCZvCA
sjgNhVPoMnlNIJm4fcxiDedJzVy4H7i5EmdIofEZZl6LrxgIIwfADxWWGfQ31SgR0cb2nghzPNjI
pbGOfNOQRvVf0BOiIzMkSOeaue3qpDcUd/MAE9wnEWtomlT+bUwLyY3uW6UzfgaT6kzpUFqcEFXr
I/+wVxuBurdCraaw8TOlh89lO7gF3uMzxObDYIzmAXalzHjlg2+fLfjU7GHjlwLtpP5XUc6/TuPp
YmL5+/DpZsREMoFowZR6hwmMN0ngUGCmYw7ChhnWyZ9rmIxmipeLe8rBIL+qIjiROv8XUJxUrA/K
ADK401cjsZ83AK6dV9rIB1vowRCze9CZQPlL4601mgxSfDPuAHXjBWqkpom6oakrCDB457qpsNIC
bnwcYbqBZNw46BZ6IqFvZnHfowOv/DKxA+l6qKXXCpR5rJbERi2L9oD/hN8qP2ACc5GdupLIM7cL
04p9gKA0eMMQZ+98+G5GLd+sIPnpl4NwmiqrB8zJC6rwU//Ngt0BWKYCi0hs0j376z3S/+Sj8dgz
9/9W5y9JALgIfTwd5nfKWpPTvih1om24ahIw1DWneaxXzy0Ta3e/QBma0D2X/6/PdsL8Y+QYgeuv
j47ihtBr9N/xbjSlNXoxPLgOVWlZ9BxiWWTR/ILatjIf4IoF+8zRvaaBLwix763voRQQ0wwtHMUe
tkQJhxxfUjaw7/4ixZpd77P2A3UC01qfwKd5VeaEXfokiNFEyozkR0Zmx+45cmWnAacR2TXd+zZh
zvoIwoxXSwFie4VpeXn1TIDlEvetXlg9zL9Im1UtKd4EeKdw+ImaerxGnR0JRct/6BcF21kmWdkt
GRsCbjLLCXoiYncwTHu/d/s/PzHm+U84N06G8T9DX2LeXY8+Y+ScJTqanuXMQxHK57AZuNIbdUeH
IGfTItaxYXvtmRalaravcYIZ65hjuUjMNUKvcKS1ZQO7jx5EWLWIIhpND81UqbbMz+2pMb3//tDu
lHyrQJS4LCZvTr2BconN4rYZ37R/LWAWS5zowpOjZ5idUiuCTs/mYzOozi4pvT4bntxxhaQgAuYy
k1oZk+2uDBS4A8blmujM/nnjuQARVrGYI40bKD4JUKEn3K3zWIydQwi4IXj/yvMG9FvwbCISzg15
w3ebnZsiAAV4hE/QfoxGWyAiNuKe2QWKpIsFMcD96kAFeEn0LNqQNIrhC8elDzOrhK/V1aY/EEam
Kgvvm/3juQzD6LXzRtr47EbHO0xNqTN97pfi/kw/+ZENUDkPhASNVX1xswT1YtyNxbZ7SOjK9AKt
m3V/zcbOkkcva+ByLKAFOjxWUqeNtAHfNW9JgGBI3S6CN2xRy8PxO84uHdI2dwcpHvmmow5BdDjO
C1llDgWC+/RHmM9cl98rZ4greWClD0hGLUa9BNec4kmuJ5bX66HADVuGhnaO5k7lov68tSynhUPm
ws1wvy73ZECV3SFxzbEu9kPLQdWO9zWgPKvpmVRvtjHgVgDLCJmVzrfr75lLzO7wBya0eOHUjXO7
vrkJzqqWefHlUwgoJX9xnLZu23FuwStCpqxaauR64Q1tEGRSUg77gnJ3Ixb+nHiCMlcvsWWvk3EF
SWuvlsjpmj7P57ywisBZWE9hjXEUhowtWBiAVZhwovHGqCjc11cVdZrn8x0yv9P8A7Ripqt9jzQn
WR40CeKBR0EZbndcEPrUe9cC3PxArzrfe7/tQMRwxiA5ssBk/0ndYsxrd0Wv/CfwwpDw+ghp6CYE
qOlUlIJeKDqmDH8Cx4uyfE1TTv6KFYDEa4sqyVyqg4X9+5Zju+Wjj1LXxszqhz7+bZlmvBvjBx9d
Fx9AtAiaaniUr6K/p1AREgFJIsCmEfOR7SZMzPK9cO1kthhzBwRqS0+68SZc+kA9Lfq5PEnPArZM
lU4Ja/m78RylN34HjRXw5HqLKCtsCXwkkG+VL5Tk6AdmFOgXF7UxczB65Brq9t0pSEidUP4gPK2z
paeeCo3Vz2BK+PQjtxzisagPOCGld3LoOC+B+5Mkqzn6WLK02mDgVmgHqn/zRCSrF3wcTg66HxhW
+aS692/tNcdfEAwES8KQJI570tjiVjoMw+TTW2pshaSokBW2HbBj4br07DD3EYR+sjmH7R3+KmcH
UUaadDHRT0vRuch5m7S+HMrqOSlpe+Ej4TZ8xUsi1HqjBp2rHD3qRy0iwJrpgKu+DiZHp7qDuAQu
D3/nllMZL3/nJeuiO4Fj8rSVwFh6SiX4OMM8uIQ4DLLyTSolz+D6QzeE5FG8hNSf+JLfyMhQYhaj
+ljaxzga4Kd9Are4ufvmZMSYn1fkP/dFmbDnSLwtZJ8Cm8p9cHr4vR++Z+cIIDFUv5ovHP7gtfKi
jZeZROBCnKSAmVLwATPLCDjy9AIrGtfjUdRFtLcjL3NAutmeNH++X8HfIsjxTEXjIGuywgzmc+Us
YQzx0oc0oy7lfQmM1xUP1bvzWLUlZIuk6yNiMKBwDtEAseNz3fcaFHhjy4zcScoTp0NterCG5Xo1
TaYD+5VyiDoqiHPJ0JxMvbQqIzSzs1FGkYxJsIYld4k0vaZBRrwAcQJx1JJaGKRPcHbu7zslLXFd
izBlszGHAkw5pf5f0i4Vx5UX1OFuobhlltU5cQ5nIYDpPEyC8xiCzIO9GjFDx+OGq7l8qnk+7dTQ
6nMmQz/35YtoeZ+uDnXBMf+ydVcjfzoWurNmJh41oSQiy58j+6vymjOl11Mrwd1kkAEW+ymCg2nO
KPN/JUy57IjxFtELevv+uUn7qeC+IDZX6OheKD6sz7A0OphZRR+kigeUZie0MpGcE934kv+kv7A8
r6NPx9cHquA0QezeH3H4RacQITURPq0YOINC5DakET97bjA/PKFGrNGdLk/u1FcpunJhNfli8RMJ
Ytel56G00vTKiquzS3Ul6GU5UmNQBcUXfnuS1T1+TTgW3x9Jp1dicW7QlK4+6zu7T19wqsbejA4i
Di/H3jWEDzTw6KdGOoekDSQG3Hc11h/tM5awRuET+05CGekvjeu4K/W5aUOt+wLhSg/pEZX8NkpB
EKkLMiUIQqpA3K45985ctguUe+hDTmlUZgqaQTV7iPTUbtVQPMN+1buT3Sqb4ZOnd8KAkn5RA0Lz
wkdlm4HJhbVlBuHIQ/zJe8ONoAk1qbRaA+vEgzMbv5Iq/JIOuSnhtxHXonZBmBvw32yp6gTo4ctR
1oKuILMpn4CVLerOZ3VZ5qZxk3LTee0Normqjrq6dvSxTOgFTvreB/eKYmi5N5tsaWPZCgK1qUKm
F1N/uxiW/gLLkb4d6SrvQTjy6tjnhzAyIf9lUg1xry34t/S9VrWzVKcm4WlN+gKaS0H/v9SJ/k3r
ED8PmnK2gPHWQkk4Qp0PssnaT6MH8fDENjXQ7LmCdq+/SVspfzAmdKY9ITNV3jq+Z5JK9ampP4pF
YECCEPPscv/2iGp0uvBDhdci09uwnQhlRcTfmU4HWqZAX5NBX/QsXnQnC1UarrmZyVsEJeJsSTCn
lbC8Wd+kW5F4ZRzozKeGHa3uFA5Q9STIPqkBSglpLH4xiwg9gTPe2NckjIepWElklUggEsVaevWD
FmIikYHGF9qCpYcCzI4XFxKrE5jr2XhGGEbPyjvYCKej9v02Nu7w2n6HUTd5XM4PwNb6u1aTQRwF
yQi1tSAJGh+95SvRv0oNNHdfNwtIrJbO7wEr78nxB1XTrZRVFSbTesz06uOiVBN/s7F0qukzVD7m
e/QNvhTG3BAlufXpndzjuy9Dw4hegpH/xNcGHfbkZjgvZpZMXCYyhlpI56agO0bdg0YACk02nWhG
0wiEFHjvmIe05P0QDytjhtZ4BUj8PiwH/zPHtjrxdNfyyE4IsWBKQ7wsly1vEMXnP/ExnBeZguGY
br5/soBNf23rwZ3gyZAZZ0yi/sNGnWJ9+tDi2hPeftXZVl1AdrSmoj8dYxN762W06nBQX6AOAC4P
sLEtKaa2UihbZ/7nbso8uyaxXrocVGi5p5IMDTnLPTYwNn4lpWigYkB+yDAhHFMThWe52xRLmWGf
mkQM51SLzrH8zjAxMGq1p+tuI2gmXiXyOWY3s1aPCtMLzl9KMyU7oGlVYMsPCGtUD5rmj4tyomwE
t1nHoGX93AIwQ7INX4st6ZkBdgTa0RMl8iTIfqOejYLlQjISsmuLHjtY5USyNBBpAPdTq3Sfwyoh
ua8U2cvgtRfZbpk9CQVa1E1uKb3DpwiGfpe/poz7+LY7ZE7K03ySmrot5yf0bIkmxsbVxaj0YnTG
OHxKig1CA5gyXSF58LH1ZP2MxratpoIEbyVdL+IOc3s8dKz9mq8NdBULL0FFTAAEfBY0Q2FWxIYm
2rSX7o7k/fXvnseC4sQ7FuoZTDZN0ldjl5tKOwdBTFLTI7jVPG2NTsMO6PRRmYMJ0ytIm9RFz67J
c66p4McpXF7O9ywupJWHqHaR3PagsqVz08YkX6zWSy68RuwOilNTK0g0taLFey+V/A8e+4Kg5/m3
KI71if8MgLxBhrW2LRn3msij4kx+As/DWdy0uy9gRfPSZvjgKNk/V1CPDgGskxDPi7WgZ7xneGHT
A8KHnI80ORr2Ve5JY/gJcV04hlKHHGEu4wnmyz25KkrEph0qoVNOdLe93xj77ELWVFrYp/qwzlUE
w7L1ZYmeIL920fydPs1+UnrXR9xJM5+jZH9MIMAzJhRzoJbX12mo6VeLWEl3vG1rxPNKvb0V5vJw
yo4ns2v28Dk/k47sM6MePhFIgmP3zt0VnTutpySiH5i4T947mO2FA4KhyibP1MDXx9LcXRLtAibJ
Uhc4U9xrKR9S/dd6jmwEnP7EawaB9dEW979TjydA2p50x24CSnGd9uAgofRGY2PjATqo7AWbrqes
0TU7XuyollGAvk7g85Q62of0zSTvkSLX15kQIh+WUnkVVAh6L7KhE2xtVeaIRnRAx9p7EmxKIePD
9JvNDZHlJD3k2Vdz0ULofeKKIaNxjYOCO2ELHgXpVHD5FXAe7yYTTaHCjx1l46AL03oFrkVhEiDQ
Y0Fvk5RylV+ydzyOUgm5J2TEbAfnU0nS3SiHldbDMq1yECsPjQAXQ9OBhJZe4OhIu0rzSfxOGf2C
Ep+MM5BSKOVvc963piROXcDCzpzuB/EkpbVc+qj6rQ8YkA+MbIk79WEeUoZ/Pcnl1DJHP030UaZx
DpkVKrlFXuAg6NFtUENk4K3x816pBb+70ism2aSYJOjBbZJelc+BMZTtfQMyhNZ6ch1x0F4xZT+B
dWK8LP+oB4F8Gi6tL9Bd1M7j/kajR4PBXU0rlPF0PKGnIC4TZ68qZmMsJGi7kKzKYHn5QS2/OGIp
wV5JylYba+SdnWSh9SUOIKcdECA4HOw6KeDE+tPEjPx2esQj2BAeE7n4Z+CIUi9b+lUoBy9lC6zJ
SbhMSjDhYYzv1ndVIBa9wbXP//30ZIxm2WUaNZf9rPi95A7qdl5h3C9EOPbM1BF+7NhppeQr8vZV
oF0UW2lo8V2SU0uB8SA0mrCDfBSJXclI6s4SnbK1TCPzKgdzxj1KqcyGtxDyN8ltFOR0YY8eiwjl
vukwo8oeDhACqRSrG720CoDvOX6DaVsxSQixFw2liednBYcXIBTpXl0/R8Z4Xj2uKpE5pVdz4LD5
+N2Y6HMCkpsyGpcrjdlt96WjKdyYe3gXNAYdjC9DkoxxN7DBMjym4yzq/5SOoBC9UxEtxa63dTRK
lftZ+J9daqph5MyXLzvA+AmjMRMtZg8ERaG2x3fb3V3c633VcgVYzUqYuLI6SZ+S+NlE/nF7Qlp4
0mAfIDhar4ZZUS+seBKoXMv2ZwG0CPK3ixVBEYl3LPjfUN/NhKyMw/aMN08CTqX0q5IjitY2lhQW
EhYMZfAddx+zilv4VJcRvlllmxSlHQqLvjNzIXXsp5bIT//E4zIdWFsu+85A2q3YGYRpi0j9VxAb
u45KGeXCz0tLgjIIHPxbXFnkv5Sz7ZSgJLUhGg/WWdjOz4UhBNO5Sip3om0/sAl+sMwxxMR+FgUY
bKXnRDcz0Qch7OFZarmw7WekI/XCrQ1BUDq4QFzHwktfEeoqRkUrjCB4HQqdu4v6IssVf9POOnqE
9zo43i0jgTInl88WYR7W4GJLTJh7J+u4bdEptLB+QCx+6Qo+/2UnPdzOT+j3iKocDUT34cFPXSzW
rXAA4FIrHJZRFca1V21M6I1OvqDXaaMiuWYec5IQguIJUmtKu5N0pAKbGcAMWGKRAb6ZUzwsmBOv
J+wSqzGz8bSoFxEzfX32OzXv9tNXRRfrHySazamHE9lZrgXJGcEl9tRUk9nueCN/iq5Ab8xlwlLz
bpvpNtcn5+X4eeXOtW1zomMwMzjpOb3ZyAFPyBmY8ubsiVfdG1W/8DxYXibqOyHGscdx9MqqdXVD
0CnBuDyMMzyjuJGQqn+2cJuLuQOb7FdH6Og18IOZrowgrYkzrqc4ANI6wvdErGd+2+r7i4Y8ydjY
HvSCQJzEYkWYTdmM8L/FHayvvQWa3ApAmkpLG7IIPMm5J/mBFKSyBh1WuAJb+xbnlHJHd4dHYDyT
rwzNt+/8tERZ+lqaxiD5hLBpIL9tQi6FR18WtAJDpPSjuWHFEuIlEVoZAZq+TCVcRyPMHDRtRD+i
gFg/oZDOgE+ydn/bcTNgOp06017Tc50kzff2UHLjd3XLTLXEnuLenyVAQta86aG2cL9BO8Bc056k
rk60pzhUp9+FMZAHauSH+Q20kYT5iEN5qpL45BKAvUahX6BZIVPrb7TxL5HPGMiQJnbznrT74aqz
1phwfuzZnfvcr6NHopXjOaWgTxgjLWhZ55LgYFLuhpTYwOZHwIZUPYM/MYrl0ejqjH1wa4eNV2YR
moEhxQehGDcvjhVnZqL7m6Hjln+GU7Mfw1vpVLWRXqnKgUINkDUSmBfjxhyrT+srp2BwI3j4Ygi5
n2bgohqdl3e5u/UEeqzVNWXhrzvj0TKyaSr3rzQUP+UllffGeBB2M/Gsb6NiMpLvPY9ieQ7QNNXX
avwxzAcbyoDhmdPVG2shmI00m+e8N37XYWjEn7XNR4OvhCPqt/SzN2nUM4KfLvdQB7kZqfPo2edx
g3d8+41CF8XjieiK3zWCp7KUMq2nlSYULxa2t3T6l4eo71DSqpVrMkV+aQgFwrgqSmHVxxFdE0Qh
C2xWHa4S/Z255e9KzWmHr/qSQ6LZ5yLFFt3Xtp/QjPYd6XZUsbTKBdRfXrdkD8IMM2F54TUFaxjh
2YKDdz40AjKVv6J2eDUL3lgfHiXvXfD4HMR7Ur+CU5FOBsCh2ShfLqKT0fPZLfmRZONBEFGfE8dH
249DWmMLs56j1bjJNvlx9VSPM5HPiiahfh68IADZDltx/mMobhV/cNpxwIJLm8E5r2mmKqHYXyNr
eEdO//PZ3kLmu2Fvl1X+p/K0YLtFF5b2cCRYC4KmI3ggPUTkFfZLhdDjJs8G+RgyRKaPDSMU34w6
R8+tr2K5hfwxB8teHGhlT1yTx08Pv8UrUWckBj4dMymaM7JkRFIDpZZyfOZZeTRzmxSUOzRP5kdw
lsKGlPVK9kT58v/4lrJS2eHGMyN8sgeKAvuk04snV5D3cPQ/+UBrN0A9/hSlIn5ayIfWM+G8fLGP
2OeGZZihNM1FgTM67Arp5/lCRb1Uv6V/+/fGTBedBko/E1TgsSZ/MNVGy6J9q1rmmnNO7T+b2qF/
AGhwgbMkS7sF+7aYYb7x15fuG96oVCLTthEcKkRKw0sooUnwAZzZQ87fJbjqRu3zJXVu5YyCBar1
mUPStz7+kFWMBCqSegclyzB4P621BO6sXkgK2xMskKqRdqjd5Yi5yASLDW5VK0CekbZqHqKzmQb1
qk7L+03WsbQGU7WhkMH8XEw2jybEFhgo27Oz4O82K8M8g+94RnFWi+0DHisRXBierAsUZbrWx/0s
Hi1YKrayoMkmbiDDDipeg652v6HagfIYTXf4MqaTQp9e8dKbLF97nuienxVt6P9/cB48sFiB8tam
DNSs/ghCxb50eVOg215JD4K9d27aB7HGOmR6FM8FwQqI5jihv6bEq+9dbo9sIV86/FieY9GvdOyR
Wd1kIDQf17ltjG/XLz8qvMyQIzZvLuQ2v4vxYSEDL38zOKI+lpqoOQpAHTodIo5uV/Y8+sl1ffcr
cSbn27W4SQIpwTuYkh21O5Xvo3YHPkGPCK1ERlFCmCMaRAz6VUVnRWlfhNh00hiFt+RwcZfRhgwz
Qo3uGrnUmBQQLdJ5UluxbBwztQvZo6OFPVdYHNv/nYWBh7v+EiEeB501cLHjzk8Vt2+AWMtmXRsg
L5024as6f6uzasKhQEMnG50x0bxEuo3jexvatnim+4aclttXSNqwV47GnAgDHc0dK6lntfoeGEbD
fraei7LRKAlfRO3oLvalLSHlUUO4n6Re9ca7YGm7gBVGOSycjdAHl2amaL7UCrDIFxyi2uLQIOHq
K+lSn8hiCp+cnkgwMuVkQ6et4LHUFT4SBXX4MVhGfWiZt+9qJ+wta8i3fn/BO4UFB6N6BaRtmHl2
oVRwp4J5TSFy3fC6uhrNX9OSASCzQIsJj2OZpbRdS7BqPJLzP1eRz+9YaMEuuAfs9TeYDtfOjdy1
a5GnEyuEL6Qo46vpTw+PIoRCYnXgOxnEG62fSwbtyDuLCzk9kS3zo8kGd6tx6hVvN38AJrSubgC6
vWPJ3P5PNMoP7oihFiuKeWM96V891OOQWrAkaBODoNNEY5tXeHxGSBVU8RXko7tzBV0kYR1Kqrce
ceBlQm3nSeCCg+MExduHNyxGpunlpNxaCr4ARy0ZvON8uLQ4eiytjL0AhOXAC76rIWC7lO92DZUI
7aiOXGK69TT7rKug2GgG++hUro167wNGAJD7WeCFLtOWjOYOWyRhnxlrkH+kEz4oTYw8UCAg3V18
Z5+q5dm7pMS8GCRYg2qYFboOaMSUivPtsz1f7oFoTdVXzk37ObItupph53dXUz314HZ1g6PGi6zM
x7B5xC1+kURax4vFabY933SnJ/oNVbcIdyBWN+EaLAeImsQw7kSVOoSOimeFu2oicov5Vk4jpJ5n
J2SlYYoade7XwuImjcLQAUDabR9a4A27N2czW1vsSPWwEoP8mAqy9uZAFKRzL+EudILIUPQmrJvD
/kokjNQR8N5cqGeu+rTNfBIlFUObAJz2Ye1Cl5oSFtIE/Q5YGqNJthoN0mrPFWT2XNc3lKbaQ2jg
kxT0052xqMoBPGRjgn/lGGy1q8ovLp53vs/u+RaV8j8UhQoWWDSxZMDN3RZXAlc/7RtnRqi9Pg53
OI/V94k0rg9383LUABH6LEY5q37/kY3b1rdAOfWq2MfbOjdnJLvL13VXQXpSW1ZoOcHV1/EABbus
3ZmO/wCOdga/a3JRFuiLuF/ZrQUU/spBFimOpD32QCi4i5dZMVgrEM83Wi/eystmRV6+1E4Umf2b
6jgE8VAtlLmyH613hdMopmJKN4aBohJT3iy0urjcTLXA6H3VaOiEUGIU16pNjkn2SLMIRlLNf1NL
znqsQ7yk6LEBaXfkmqCHkNwZLbWFYamOQSjnANQXRwNMr5XUfodMoNVvrhX1GfXu3VGXHXSKkpFl
IHhwTAjkBMxEA+FmNYohdflTmKIlA3h1QEAKEUPbkZrlebEqqVaXfCMzQAefsOxg+t41y6tB5rT5
Y/7tSQVBORSPDjhRaDm81w4rB/BoLWwTAIFU2NM5uwHbqC+PkI4kUb+veRziJNaa3eMN53WOyawA
4VBO0RVnBVNOtUQybsgdxirdKJK911a/HguNFvMJloBBr9GrnczbHuMsFrk5mCWovaF9oTHML4x5
l6JTJ55I2kiSYt7IWT0DMPBtjWziBZgv+F2l3Xvtfg4fPqGsjLG5Uusgw3NvY32XUNA5p9d4mLhJ
cdAHMdY7/k3xQEXQGKqyW+F8SNfcc6uJbI/bXDWBFsm92LdtI+FnqAj2kzvR3YbB8/32srdbS3XM
e74HEmOJFifXayFSgpR8poxK4dQmpMXoQ/pMH7Zzqgtps96KyLxtccFlut31KYFYiiXHtu9d4Ooz
T2qw9I2YJJhjJ9EKNskI33GzlqTMkYMwDeJyQX71HlTr8ofTg8qGD4nECkp6R4lBhKNhM7s9cgSt
jEfbP4ldtbaHUSGZZM2/ye8iZFrD6m0dpwigUXV5C0MR7QDldkWTrwv/epqEzTVHNwTftR47smJn
zrdxLnatQc4G5S+8KcA4OtZK+BiD3VZRX9e9730HHlz3gGgpFDMkq0IRO6okNoMubwCpOD2WWyQ/
nk8ZyERAw8zTMYX1UwvvYyk+7oXoqrT6oYu5zc+3gjf0WWNcob9jlFDJjqKzt4g4XScEiVKcXF+j
npZI38m8K1ShiKrTvdvmddOZgeR4AFD8BE+yxmtTbLBEqlIheMyJTYeqI6GGY4FNDtB28xUfIj9B
zLv1iDrXLp+Y4J60bFk6bVfoEkHQgMClJzvGIHktSpWd4EpCFI+808BO9BUEqohnBlhjOoMET0rt
Jb102l2NGjT34MHwioPh6w6RhivUjV+Q2x1MpejUyd5bfKKwd9plY/M1LFEb6wyDhQpu+7RemyIX
xLX/MGaAGqWKnhysyXEan7P9ICwucU5DjDCA4pMstCtj2ska+9gmDs7RR+7ByUwpBvVE53irhzwI
nz+iNiCDWQTzT1FUZW22VUy+mCNKhCK8Y89enxUT+8EUogtwvg8DBZLojV39e7ASqP6QEWzujrao
8dZa3Z3krbVUAczgXzvMiUTGR8dOATteCcoG1pc/5t8UQBgAzO6uH8o5qaIuwZnSG0Ix6eH86S8y
J7UO24pMlr8QDKzWLx/bGQtWBFw5NMigbcGWlMYt70J1L2Y2JxYQ2Tp98gYZ3XuP01EToyYIhpDZ
/sF1/YPDHOoIUB16EyBu4ffrfVntpz8fLLRcTnrbVQLOq8XI98g5dsWyCsV7IpBsXKnxvwHFMH2O
oaTqSHbdTE60SiLsadr+5f8y3P2JlSIGYRjjxXBDfMx/SaeqImicbqwRF3WPWGEjsABbID9y4mch
v04c1rmB66kdmhVJsrWCiKPzN9Yc38VZ9hLdra9JGgiowROiFWz+oxitIufHXTnkexfy9hd0uCNE
mSxzY6Q3LYpCOLCU0WhmNeviHdtSbsxKloOarDC9Q1egUD4aG/iGvNYYo+KQCTP2aQwT3hXHpNMP
RkoCLuI7IlL4N+G5aKFBllQlheiMnn7IiTvTXlbkaJBe5pC8c1StF2w+chixyf/rKgyHL1WluL4b
hTSBlY5bOn+i0gC1+6Wui8crWQ1aBjBcw21uI561vRo6LNu8aStE4bCS+6e7XvJtV2PbGGb+csLB
SwIAStPCrVTrimY0Q3Mk/nTdjm3EBkJ8a9pNSocfndPSrAMDdwRIp7lzQh9INdpilhYklqkDC+EL
tD2lxqrcJIEVAcG7/cYP3l9VMyVesNvmi4Y0xeomtxsnr+/LOIHSoxocEysuU/2xcLL3Fyu+ufi9
Z2Ptvh5TEkOjgRb3XvDQA1ZNoPZM5GvVfIrq0RgfAAtelQVeOVUIOHVIJsgx6ULDKeoYyvZxPOZj
8hlP7Y3oVtagOwo6HCHFeSqlmnUBS0ToWBJLAHZlE162rgdWLmSpr+86hUJkkW3/Xy1m2+IuM2m6
SgybTHhqpX9apJdbJ/51zFl8SoW4bGLrR+sMWwWenYF4g0r4zqZd7i2m1UwFX9FgugTdXn2KVlWy
TWa1C7yowccL5VIq2ZjNOq0lwrBsG5NEvFQSaNed5h7CnJ4OuIvM8IGXnqgMwbB9Hwks5svGFG/o
A9ckkzVNgCK8dAi5WBi65ifdC3oGr7ChTPdm/X6InLuBoye/Xo1jYRXkIXcUuJD1wF66wb4NZAdT
K+Veo38Hu8GIcwwxhHSvFm8cfBGx+gx7YPUOw7QAoOXwtyqmOEHGNPX6vANIotqHNw1CVRswsjDr
ED15Vdh4pLjAMlVuvCabSFrRgRxAgDNk6GAk3k/N3pRvJtPIUUYGGnC9j0g3afS4xEIqDImfe8Aj
+jtDN1szS6p0ZUHMxymq5/x4o1cZTfC2CB57X0q2J2oCqGEwODriIVeI3yMX8mfUCef0VbYSfiVr
pR3M1WK5kXOhIVTCE6fDAYvK0wqyAVFM4yGOqy5Z1uV4EJorWbyMcSbvz/3B+pPiOIcsM0mvCxU1
VvZ3TbqlDEKVCcRqJC13mgljwnMb2BkzlDk0lSYuyQuM+ro5fgxMSOkJLXjqb3IFVjNTfSOWM6qg
u17VkSKEOI8fpFqX2CoyRoai259eyC+7xvWfG5h/qVKwb44CnnsYqL7BaDLP9Sgpw2dhGnjUXVdK
/l3dlf+E4aDUNiHhP1etiFVovulQ0OCBmQVHCCEkHM9cpmxkI4X7qyK+8Qcc6M8VNu5DZrPvbeqW
tZhCBu7mSVyTUOKAvHIOBCpBHwEXU/A3UVfQqTIedygJzYxhyYUWH8Jhcg3s79zQK24XsuSjwi6H
F47Je9XvT1gqYcQMhlcL/R+3lMeLJrufVK8l8VsV8khx4XbsvjEy8yNear3uYaQRWuRigX6xLZ7X
kklx6QqCOnlmzIWPtgpC6yp9RIF5WsxnN6z89vDFIvKMW1hwiMczQLDuONhefTwrgoSpNU2TKb3x
uED0j4fb7/iMQRKgq9HM0S5ZC8a3oBCzlymDMneFMYErhNO61GXLCbJWi9jbQy/ShwDLjPrn/yyX
jBDlVFxbHFlQ6zppB1+SnZYUYZU8A1SNiFVfP4u8DarWItmW45bavJkJF2WT529bHVPfehIYM/f6
TsYpH1ndEvD1LnbrN9Q0wB81KQe77X17aZg6ldC1WNdH1tWtNL7WBBO2b6I9U3jPUPuFryfB40Ll
SfH/X/aysxNoXQwwj7cltBukvp5MCBvUMw5aM2z7RwKTNuvmYCKoj+JrWzGt74u30lf82AEy1Ciq
c7grroSH0QhOslrde5rR+yIz8qABX6C2yV6/+jJfeBPTugvhN39KmVHz9Wr9xlrvwWM++Mz+sCEf
3gxQ+Gt83G7HUAUKugQNDb8pZtrH5WyrFy5p0nB0pgnkywrFAHrDOT0YinQUeVT+7YpVGQlDBFx1
nANjs8FfpJgIaUF5/XrpUPiQcwc8dtgdpYOzmfN2K2Vt1kSCihRLcrWYKz/VU5cdG1cTySDS8qmI
AUuZWpg4lcww/0IA6ONsh2eMGTYfHbtsrsIdjthE9p6rFgT4HcfjWgz/jh17UicIaKkVlgBBzSMY
iJ8QUASnC+ScpEYz9JrPToYLFpCiQ+Xf9CQ739Bxn+JhKfz23czb3WPo3RqxQ6hb6etdc45LkQXt
d3AyFsI18aXiXu1YS5+hTXOezbJvo5ZAk02+Ixlcw5RFtE/cB5j77WOXzN0NKGyHwHdCSZijYEbm
BVNkUJQSdD49ZkkPGVzI42r20tiZiDF8DN064iinlgxPQYdoORAiVt8Hp8Xtb/pLJoL07HqOiV9W
v7PRZaAl9NUYqjnhVHKdmfvQYWVTaT2RmqJmmkg3Bx6UMpeawqMcuguf9ODrySmNhbs2CXpNRVIb
Ik+c51M1eq0foYae76uFjjpVlKMygJR6rEbIIg+MiqAfyOCoVkxRyoXCf0UmlMHwaVRjI+aFTV5H
MPN4RAN2pjXC0bpOW4JzV0tLHAUUnsv/Dq+71rNOZxQcLOY7Te3Xc3EzyM3P5fuV8XNcPEbWphKy
7YFEDS+VR6JvA2VsZT3sFd8Rf5KP5muWQI3EFLEfVI2d1Duds+UX0iJB/1ANewB4KUlS9trDwplc
4cghLIFpzXuf810Wz0xJJNiAYZoLmC4/UCaiAIFuZTJo7tYC5jEi60VfQ34zJHW6XmEIdXR6MwD7
4r0eifmYCEi00ehUgEgXBvXkriq7Q21wCtfli1JqS3fdfErmPI7rxJSzMgLkVilEWiVnuwm7343i
1n7tfUrtyWzZMfkGI598mYDLBlb7dzm0RFetHsgZQiWDeHUCQZ9Qlwy55jZ0tW+eSNRf8H6PkSD4
n0mySsPop47D9Pmjkc2ZRRh1m5pgnnm/d2EWkdQpDUAZY3Lk6TqA/gOs64ktQQAwuKPmehbaHA51
iG4wvo/ftL2riJgNtETS1d8jxDc0O7W4bUVLkGcUG3rmqtuHdFYjWiCAEKWK/jHzGWWaiMLHILK4
Y18eYb1wrq/gNcA1ediWnKu7ymuVFWEAt9IGYDTVQ17RbIx/wSuM+3G5aQJxDP8JVJfuLh4chuhp
I4F+eVy3QCASLAZaSq7mrVI/+Nxn7CmLT6CJt75h9np/icKjgmVjJLW1BJFkf5sOPugytgUa9BLb
Yv5cGBONl3CqIZlwi8FL+9dAa/EFuhIMrJiqzhQseZAlgLONxbO+pN2sIXj3GP8GNKx8QYqSbyha
LiOJdUTkWliwIPD0rEwWah1DiFLY7jzXf3Ykg+HmjS5MOEWyKhGTAtSIpi//E9Ds9k4Ct4+veksX
1qmIxyUCP3gzp77fbj8g9FwEDPz8bkhqjwf/CHw8H9+EOWn7mrCX4fdQMoTer1Jk6+CWlpy14+wd
9xP+7z+YZUyJAqR167TGQ9Hu5hK7vUFfnRJfjMRpSluRFY4/36dRuI3R0ZVBCSZ3J6aJrNoDcTdF
S0N+E4KN8/Y3CVeC3gBHph1d+Z+SnyE5ddihdD+isXR7BuB0ZeN+wJ7g1Or/3rAO7eDDoapXNgXD
hZFqX5xJ421lDVV8KH8CWtv1lQ6Y0Q5Vg+xhazmd2lvaClp6TStGbRhdfePn8vgPHz1hikaXNNHz
gTkUdkIiLi9vtp5TbnDUWG0DBWVIjzwCK/KhVct2lnXOdcp9MRFLXc45Y4yANvSwOzOnCd0GOuoK
4f7V7lsifYQtsUR3zqFBNs+gKRdDGsQlyZLHZg9aFWfUituOYF3brul946Rb1BNftkJJn2xSfGVS
U6uPhPlb65WYtDb6tfqmWTe4H6MwMs8mJiVQ1YYyNb+nEkVMuvXTAGdyBHk0mdqD12lYixe90uqX
WL8B6LaTLv/9CYTPdCu9q6LiMV+q/9B0udvaIxXTsCFvhdAYH+5Is/jNrDssR1FMwI5KYQoUUOtW
xqp8LYdcxfaO87TEjK4qDs/xT+Zp9JhFKZHP87/HmMRgLB45gwx8PF9AphVI9JVT97qEXPcpJ6HG
Mpq4+5WN9sykn+8608y3OgvSwdVMTc+RrirtFrDB5/3yZueiF0Pl3QkRJ46G89GEXLNs4Mz1hyGD
zJc8XZAvhwevpDjz4NOW/mg2dsaF5hYiraD1VjmXj+4pQZ2J8kSN/hrI9AuQEX3czU1AZQ9E5q8j
mJYeHA89mBTiOodBB067mAHgJKcRrSsveV6cd7231OQd1SewUtG2MPWk05BAdTi7yk7xPDTrujO1
F1deMdzv2g6pH3eJH7nkTr1XZzI9/CgARs7F16M9qQ/eVIBw7H9MTFFhocB9aU6Tu+oNV8R8SdN9
/mc3AjZxsTCG3K05MN/Jy57u+k8NVg/3KKGE9wSTw0bt3oXdXVoolHhCmWwRAlo37/mtAVmUSah7
abN500cG9jnLgAbdeCefb6ukleJNf+PN/AqqoYNErWTE6Tcrr3Qhal4zSHLHu//PUeS+eBR8eQ1g
4F2ItXu5GgJ+FUXrq+dYITI7FCrMdpZk8z/RSv3uc1Kz4G1KD2U92mta5dw5scAHrc/cKzi7qcFX
ICBPXjc3zqgX8z5wPNiAKD6CzscTAJrNoa39xKWwJYxvVdc2IBjaxoti8lR7ULfUB5+NiCaY7tp+
Bhm3Ml6zhd/zxFYUVdApFXRd8Hi5f7cuQ9fp8c0i/ldLVnhPFi+GkHag+mR3JF0SBpVA4+XoXM4j
/z6kx4dOtXBzQMMEsYlCETfVEXF3jTx4VMkTf9W2HxPuzcYJg0TVnP+SwJWbSdOAh6fjOWlrGQVz
I/+jXv+ZsucVw7G8EKic5y4vTLV3zcEt9bLyAkPfwa5Pj45RWQpLdTWPghmUmfZAfQjrVDgHvMNp
vYoGcjiSofg79nUTuRfCIS5ktnwmESo4okeIzVZ+NIz3Qpcr4wKzHuMc5OyTNeRM5QPEQ4/MhgpJ
3/pczXNEbUiXgBUpjkcyXpXWAdGhRGcPCvbE5EVJ9F7A/GWVtPwYlTM9Du+AvBQji3nvqiAvLSZA
tAn29IHzIQTvo3/9nxLFJVEaw6XVmA00kgHLOlQmWpUxlnusYFEcGpU3/OufSc7koSPs7o/drAFH
1XAN92FRKBb7IrdGl1ZKciDKPlC7WeCsN2OExJ/qK/oEAL3mqs+xa30cNRQuK/xdACyHz5alaWuM
ZsTL6wHBbVFX5IUEl9zS2GmBsO3YSih9E9ZgFMOL5N6ERYU3/b9FFaYqi0EbTCANV7o/6axcl/XG
9kNWs1y7tFmGALmp21lZldYGc9qWzsG7qjqRTVc+omMPjUIvQxQao2m5XzD1wmFBwFTb/GYKRxTs
jt7ALafkkk59Q9f3HXrF7/YSmIRrbzIDjIA/0qFs1LN+fBSEamxl2iJSaTI4wM7eyimtHxDA81me
DQDHxZoVF8MaeRW9RSCDyTxgc1ofsT85kPeBYaM2K5rUDufY0l4DXnlaS8JNxsFRZVHjHICZNqQg
eq0SYMvwNZ500EmqKydrOMNetgbB/P1pjzRZ5jW0xMzyud+3x4pqyYYETvSq2h4YfjB4lP+NK8Kn
Ht2KHoAEkktuwgedony15Q4cahirm+S/l4fhsKW0t6Aln7dTNU+d2EA2bYUb67xZVHf6/W0mWOkM
bPI12zMNUc0ItfUvYsMtk0YxdTodcKHDxxqqDgNqvI7XMmS6vpRpD65qcAXFWwxZP9z/h0FnbIqx
SJr/ZpNzPJlIgwZm50zcqP8KmyJB2YSswQ2vNXeJxxrdITZ/+HKKDQKR2UQSOlA9tmet9toa1DVl
zZGkLzLvj1bGagZ0QTKCVBmmS7ApMbJsjd1b4CFhAuRoi1vAqXuc7ebAMYv6s/ZGIX4l+GAxS9zY
GNXrR8oUuiy5Gku0qn0uPBi/0ksSwXYpurGU823OzvGPUPdauteBrZLvQkDhZ61pF2xePQ2+M7lb
22EGeUtYCdt8Gw7mt/VN+ysfRzmb+VMsCJ4jUIuS6636OCIQKD+5/bsSeXpnZ4pLcPxswEpxLWum
AfgNLQi52OYtRn5Z+e8akkoOyKuytU+3PGj+GxEkCeQdTVMgR565OVnoq84fIa6DTXlfzjXeNlJZ
OvCaESA+IPi/Ke8DnsfeeEuNtlZWqC0rthVTeHgz99M7tYS8qW7UQqYaTsdksjjEaklu1TTcFub3
wYWpK96sa1CopuN9Ph3P/5xi+FawAMJBjm9rZzYWdMUaHGi39fJIFdqREt13JB7Zbb7FX1ZQS62J
vZY3Qpg/3iobkQxrK3GDpterjLNQhmSw7vcz6dV4CTwmBzIROs24ZSodTex+Pcs1kgdAPGgDTpbT
BfQMOeCNlS5fto+rEMTZL/HodxQ5j/Gm6qgcRCpom3v93qIQbGIc/BEwXlmy2LaYc0Z4W3+9fpbX
yMTE3G46YIDNpAmEiQtUlCkvlPQIJ167EMYBcCzLmWro1FCpRlr9l9sLv4opjqis9v4m0/1xTvx6
lpy52cu/DZACbjUC5LF8uA4BedZoYzcDz+Qiz40bGy3pgVpK2qffyfgG0cLADVCQdBsXH2VDUCO5
CZvyYOJL1qBgJCGSaVqberr+o/6zk4GebNkW/JO03qKbwm+6V83SKGFKkBNwhGpWj8YnZAdBV+A+
Bfvvn4x6UrTVjbP03grVlGrq/xt60A1GrNIsISeAfRPWFbtATfQQUtFwJZEtS91wjBof08zj0v+6
qvyXW+A5xkHSY16Zee4PqqfkALpuQd8cg/zvxB8z8rFlMc90RAD9ulP+R0pg8n/uI7NAj/S8LHhF
+GKkg6JKGG/qydFLkK0lkwsFWjGx7FGJTq1gwyaT/jdi1IFxWBJI2ixmHVC6KZO0eExOm7l/1D/l
JqE/LM3wZMR8pPDP1aXmBw4g+ZvvWjWgpbC+ksO5HFJLcN9Hlu1VlhFjP01mxOMUcAmtmMVZFi+n
LvxdMtaCCbBmJktIv2mcgx2RqRP5QFqV5SNkYo+t0SGdrUtTKtVoRQx/CRtrl9UtgPlVoTBfC5zS
B4VeY8zaDAp8yY4n9BMYNg6/W5eDP739g0CmtShQb/v4AKUxxQ7MpyYAW7TgAtn/LGCx+IYSQIKh
Aw9aku2RSvFyGiHUajhC77XQoQpec5UF5XcABRsJBInnFYbHVQKh+48U4z0PjhqVAwkvT0mZaP0F
1aCEfoJUVuCjn25yjslTeE2kDhaHo/otVeoxOKeJlqkJ/pRBDA6/h8OFw+fbJCLplVq2fy0b5Vrt
/BBKvQyUPsTCqB+p8UZaNXO6zPK5/0tBc+uAutou4E45KkQdbQ76EQZQqAEyynuVqEyIDUvT5A2M
S7bimhX4GCBbvTj1IZI5MjPUW4JjE8wVNIcwMRFIeB+992sJeAuXB1uy8crrSp4jeAVEJatyGWDg
05ar2plM+K8R5YjF6+dAboXeqxEa7f1CR4yMkdKTnFbyrDCZf0Xst4iXMuEK++Vq16WCk7XK+4/e
oiCFVKROaJS1Uyjeau9ssQ0V5nkKIaQ86OcslxKZxbfBOC8Y3zRQVTWpXHF2uFL05Z88Ke3JpMyR
W7NDNE0dBm3Y5vXj+XOzQt+Vx76s6pi8BcNRY83cENieXaujuxI8xwwe+951o+64dYlBFyWQW3l2
hTRfpDiTLKXZEJUefvs/gVCMqboE73JmNRvnLuPDOmHmo20ZPjWlfmKqMPoaq+vEthnud2krObO5
txJm2c0DetD2zz2ocBVWb5/xqvAxAm0fWOV94ouQx5thAVIlPcmy599BphJc4iMmrzXqUbUDOj6t
pG9wzxPZTeBd05FKKftbwdcPDcrpMPoMB/aYmcWYr6S8751DNd/rm41Mdxq9ekJfaf+nZ3KqvUoM
UObc6ZBPoxsklkSAt/dt9G9sgShSpSwUXjw64LAn3KWP8dc5SqnOV2e8f2ShjvPhW1aH3fjLNuoQ
Ky9+YqqAHqGsHBXw098FO230m/VUUCrNZ+ndqp4T6sutCkZYfUzu4y5EsPs8Gj82VEn11sbkPQPr
Rh+PMy//NeRBOacbAN1RyuqTgTyEEVPg5GRd22o6ZdgjecJOp7BwvSBD6Ek2GzlHGrGdePBSd4nY
wySrxlVh90iD1CiJuzVTgEm9/C9j5kuubb71Chs/bNORUz8Y5fgQJsGigu4kdhiLDbZY+vy222rw
G1ePBgQl3/ldSEvwyaX5uCFSQKQfRzUANEMppBgprvbwFYZ9ve7+cSCR0FdWuoVlHpfPyb0pUiRl
5zCGuYCsvFa1x1eFm4sJ4ZA4KOF50S63kju4hVwi0syeORDi7jz3ZtuW7lih7SlBMOrsKFzLG9JT
YxLYDAcEYXTbOT1v6ejIU5rL2onOCvERFwj8PRatFwp9yoz1Vvzm0/zqVGNOYdltQMfAzMUbzImy
mRjZ2a7ep+2OK9QWDu7G0nQGT+PumRhlJK4JfqwhWw50oWn5QZT9BgEANcSbinz7W3a8e4M3JoNd
ZIPgfI053GerBp7XlBKcUwTWDcbuwoBla4NXKG4Bp8QjtIxS0w4upDsJCXYDcaKf4H2wts/r3Ko8
dXxpWcayFideliAheE/welzaMRrlinAKapi7AHbmWukJsHhT1oPMstbEEniHa66SQKVmvUZhNTWA
Nq1q5UxhbSmDlqd5W6D/E9AukmPaYgRDSL045fFovNZZeFcagQdMQw784jtLQ+zE6G02GyCCmwq/
FQYJlD8MINj4YcCmZ+ryCoNPxVT9dsWLwfaRmLXO4B6bYsXasH3HXij8lmgPutasTZaW/85UJXqc
tQFuvec0q2xolBQf9vsPGEQqK0duT2GoA7yRDUD91E3elGU/2XoQQ6YNcDo0/XjxD6QT7ryNaZe/
NNZigRx7+XEJ0X4NjH+qj1sOKz0LNXqQS0BqtU/FYLqHXDGY3E4NdSlfkq+4w+9D/YvPCgoYW9xe
dslXHzFdm390Rtf+fUKoK6vYRR8eS2g5uuLUKWGRsIiHufQzz7A1P/vda+zYyO6yGQ9wlj8/Ysff
WHrOVHcgYdbkB0s3eL5LJATl17FDac1VB6SZiwE9vfF5GnzpTXg/jwfdmWcc9pWFhpxGBq8tzAZ3
/YxrueYxLxqUYbuZG4UW58PhMNLslqmENTTJX3rXLfSFfAP/nu2+X0Mm550cKlCPKMCWvFal2GY/
Sq3GcuyVYIdcpD0TY3c8i79w0nyAhRwPGFyWhyGnHQeXZKvUHW9aFNYW2wwFWlJO+tS4+vqHX5sL
HEspx4yzKEGMSfuyCH3Cs3laUID5jNTwu54xCDb3FtN1bURf/rl3vm4y4ryUsKUjetK4L//IJBF0
s5gGs90RYrv7/GhJb5OT2Dn2UsPi2djtBEZXwjGRQihQ/3AhK7jH2ILrIWFE+xhDu2PkiRY+2Qoq
BRqKWW7Ca66us5iPHeFdIf1e4aaFVVdoR8XtsJH7FbAViTRRoWmVoZTXzui6DvjQ60PRAh+K4cxs
MbChfCPL9ZkCtFQBYd4N/epfXynm3N5IiYG0qjTkN3XR5FRZ/eslIY/FwgCRGGnQ5giaUageaa3s
X8elapZ5dt/0NUui4srVByS6m4fa23My1AF0IudhOK9h/KeY0qvuwtM2WKCgZi3HMeXPxwzJKUY6
LkDOJ9UvfWbWxBpbwaPKK0mJxN5jN8jIlWPVpxNQbAZqK3d2nq6WIpGpeXCCSba7DGOOTQhg8Z3B
zQ6gAtdIyCjmfANELk6d+OLo8V7jQFe509kog+s9AsfhMDgmEwdnTnyor0/B5izeDTFw/BTh91rS
gT8r018vCTSTs2zMz4RqC/qMwizzHqMpmdI89oHKKvZqUUPvA+NpUWPmpaGnawylV/kjQ1T8MpRn
ZnVhhdFGs3mU8xH+ZKtQtj8ySwFTo/Ltj/Q7Q8GXI68epUoO1pJmcvrkDfZE8mPOqsaIjv4nSDyp
DG6gMHihnJdQfoJ3eXGynanZ4QB5Fud4RCgQPhYVtBpjWz6x/CGYcz5/9Aqf+FLIDyrxJlVM8kNw
PxjHSmIAICm/WCQGPdH8vlWtYBuDkbm5i1/qcj+dI9GhuiAdGabwy47L3/N8L4bJgUfCGvd8PdVq
fbjVIfaRNVGqrA78eBRSa9/MFX5ifdvV6o/aZaV1j6k75Ix3y+ETspeN9ZNfMZ+QSKnKc1/lpXe1
l7S8oegrxVK2JC7TpO0eABADRKEaARxWtxmNVcNUi0ZMa4N+oT75IU3ST/y3jbViTh2+aqvhAbNc
+xCq48pYpkmMVxq/crklLbc+iJNcpIDdk3/igIWckG0N+v0nsQWJPFOo/rAa91/rT6cMqeSMBbn3
Y6NyevyDX4Xuf3A/sJ3LKh3ZTKKoi4lH52icYxrlIw+DEtMDyDfSz32eSDcydadSUJntxogyvTqm
CXKbGOd8JiCbhBLiefjifBvHhkOdsS2OXbcO333GD+AcTs9v3PsgO03tWEGga+NrZppvvTpwRrJD
mS2t7VbcrItWTQslPlKIKNVso2/3JWNRukFbV3BIUgqh69W/tqrGMG1rOhapUsxREtTqji2sfGi1
uN7m6wXXKz6J5OYlrFKMsRxGTOulxw4vX79zbrKCsPnURl7FMxD0tyGaal8j+wQteyhvSwPXppPq
4JXT7OyrwGNkx/9hKi0kPTZ85+yumdtKsHCPt5Ow2de8MAy6PJ7kuqnOqfQiidgH24DnHKx7aS7Z
MK/Lz3XKzNBFHuns74p1H4zDsNrTlGRROazFjOfxg10yNv3NjiQJ2xQVn+eSkG66XaM4cHt7ZaTs
mqlCCrrqsIshXFpl85kQ0+Q+F3WUatbr84MjsU+ZpQKvuprxppAVe+X/89lbIn8uUiCgyx3NA0r0
hz4KjI7qmcPsH4GdJReuBTjXEsqvcEdtFnlPkZp8sw9rHZSUA7gLroONoKsSLZolnz60Ad1LMYQp
aR8a0INNrJGSFMR+TxyHh9PdysMsqW9xISD3JSjf6MAm+EX70lum+Q+zhpdaJPBfqOyWOOzXePav
QF4U3y+PtvEh8KL56Zc4bL+kOeb4erV+hWqqDfu8b5nzaZmsg7LAip72jZXT8HJqg5Rn8VhooUkn
/cKvRiYXjvYdw0darOIIzRGhaTpacKVKkTRMdODJOGR2P0Tsoy8QhGXRoBbl9ZzGWFdzqoyVgcWR
m3DjclxW+kh0+pKPL3nvvmqI6NEZEEbKApSA5QZLAG+2TQjdosDiEgRZgTqRZKFu5EG/7ZOuBe5J
ZbvlttxXMVhZU4p8LR/3vS+JYOh3gqs9RGT7OuSKPnNruYTsMurcKwxCeFuYr7FWkqleCkz7yjYK
1DVkn588O6sNjOg0Dc4B153kHBCbrUszgEPLCxGKbGgGGTBUjW+Ch+7rwLlPhzxKe68FLgrAj/3/
/aaDsImJbwgxnWteox+Mxvrn5aMh+BG52gBzFzo/UNz7NGvDzahVuvL2ADI5JA41K2c5J+qq+WoA
g9SrUhARy6CvAsnm65cmILbZyh6jw8BeDeARECh/ghru9yE0yfOafnrHHZbRlWa9uxXvn8pvgmWG
VhsnI2XKWDZqS1u7AbDsgrEcYqLuNbU1H/dfsQgYv+ugWo3I85qIGxWdsq1v8ScqIu+MyuKjUmZB
EDpYnm/Ezkat3Gtq/3N7MqylacwKwdGBQh6hnXizBChGUCzt85Uht+/1UxA2Hw8aQgWbsHIW/qcR
nApJjO1DO5smnG5JumMjw9N1EB0JTa6+6P+c/7mmhYgxCnuaMumLDxaPB6IGf5XMAvwinSlwZd2x
ROJvGHKL032qSW+rJCmGKPWwg6zLJeXfZNxdT32qzP55R+e+4iR3UhiMiHyRc7eRXTgrXvSvMvZA
JNlCCkTJ+vaCtYhxtrHN7qTG4jeM92ZLu4bA2JVjqU2s9b7iL48lUKCPPdJRq4TglP0ExVmNx7Jv
Kg0IHHgMOomE3C8Z/wb9jZlLfQFvrnlkCiJ9j6rZZ1SpKwqomAwZnQI7bhh/No/oKYoubqfPpje2
gyIG3n0xVjaqm8tR/4jSvJNMcJ1lslTA8rWppjeOfLe3bxud/N7TLbqjvEtsyXMYAlhRLBY8Ac6T
P08PWxkXM34n+orO9sKd07FsQorn+vQ7WnBhfY0EZc2iMZh+Ohz3t/H72cDt8yJMXZDTli/ISidw
6ZZpb1Np1YDk/qHsv34onrFTwNYsggGxF8m+yPBTW7r80gwBRgYdv3RB/GYCtCsZ1VPVJAa09fRB
O20vx0OUzFdC6jzuVVDZUDiwLr0D2lPiHPAdMTbsY29myDoQzGK6SyMpG6SQmljwJemqIcwHaBA4
lYOhjkIFlhgcQF3CPk7W8s9tFRYu24oE6kvcncr7mIBQZDaMy+jZQcTm0AleV+r86GIsEQAA9QWg
ylH/EnHqsN74TLStb6f3+WEJyQB8gHCiMKmwgo+/Q4U5RB+vuV8XyzKPCalOnahE+dZKcrxBHbQQ
HFYgKQpsGkrFmR43or0e6FgMhd1478dQRBaE08Cxn44+bP+jYzm9g8A6alcOMy06t8+1YeA8myaQ
d1i9DL2Z5Bg9dBTRgWjohO26tCc5gS3qKTkaEWTxsuD5JoCEqRANVThRIP9bEVJ5LQUAYzEUxavd
Dc8VYHoFof6VW3pY0ML+sqgVWVkGIq9jdtHaXR+64HDUUdXWUlLyZV53G9Nqb/SoR8hzph5HQnqK
Op6Wyhqwa9eQFcnfblf4XhPuKFQsY449K05v2wuALTZuS/iVldN6wzd7ts+XUCy95b8YA74vy8SA
j7ylmgIWco1gtsdlG6QUH/i/p56HXWt3YDSTpeXZFVADUfiAK6zknspBq11IEBF4xplaFtKFczrS
5qCjCWbtmFV+7rmPF+hbX/1RKQyCzHW0wmjz607qhoayIDH9DwGakQblX8e7D0iwa4a4Portepu2
DQQeamrNanQWL91Jbik9ZMJwcUxIczacoCsPgJc3LD3b7Uw49P9/HAhJUn9DRMAubu/IG7OK29uo
JzY/z0w0otaMa74P58LP4szwalE1WJjgBF4UYImek5FURZm6Smfdbkb1rzqQ88Aw2NOXzd9ND61U
QdLM+gum/2j3w+j6ZV9lSm9v0Zvvv6oRaXGum73dUbfRiOXjg5tndp0ES0/d6YDAdKN40rlX/zSa
ILpQ3va/iVuUrNRqWy1dz/ci0LFA17Fm6jSfpZSfWg877IRO7CwgLkOTiNmnglDKVrHi/KRL1l4a
GXlDKIvsd+Zlr7SwlgMKpvVUtSZfDagqrajaOXTyORwJBnOcWPHDWDIYYhYLn+nw94G7zbPbCxSw
h8wossTf8lX2VJdhPjYYllZlcAbR0KZvHZn8AbuGZf9mKDoDfAH7PV812JzcmI0Y2LAennDIaVQm
EVz/ANsdTPyJkbQKk8dnhkBCVUrCke5l4j0lbDgcqMVAfhJl55GbuXrqYvaXuw6aZqxC8gdd9IjO
buh7A6kZU1b/UrVb3uWdbJe3VdXkGEac7UBs+Bza+Sku50Nz/dPugaof5+kvC7xH/UDu5jpa1xrq
O+ZsrZ3usYdfV6Oyo5zPMHKamZDxuJcKrKBbWDWoSlfjYAapcQItZYG2TKieTQfVn5dD6VG5Z9l/
0QjFbAzJ7HlJX+TLdjF8LiEUGlleFN8D40qqrvK7e6q+rM5uvW9tC8K4CQnB9w172nZHzYfyFSGh
Sd3vBu2WkuetQgpw0urA/zslcAZRiRk7xEJp3XtoZxk2ve+zLINUNtKmwzvL2QvKvqDn8ECyuNp9
EukcgBQ7hViUezdUcm2ioJiR4uFUSWyukT7ELTAmO+KFcbzBI5ZyDTcFGNgVxUvqmVUWvl0JZ5IK
i0Nj8dXo40Qww9WUbleHHpNCY427oaPhl3EKYrQfoy8oq8n/VRtu4Q44TKLMgoeWV2dAM30cI0OB
DJspz3LKuac4Dly9BkDJxX4o5rMOQSaTdOjVSOKyYO1B8+cFjfSRs2qj0GvFr2ubG/nqWn/M5ZY5
e4/UF8/adfsPZHgSDnq+3ONomWo4CcQtJHXg03LpOOuDxAae/jRqjtPZmkyRW2wzX8gqN2HUTJLJ
zEkh68qfvSXgfibw/V3SOrgzAIJkdQ9G7hsYP36ifRX3nvuMIS56fJ1TVLscuQc1PNG7CUPHni6h
vlmx1iOR5LmK7tu2xJ8jLGpHE2eCl63yOnF+1Hi4FGGjLLMS0PREhZwn7ZnslOS2cRKhMNOE055u
Bmq9wIpqCGRz3vFfCFTCcDnOeurSXIRifdH6JBc9Gh/Im3e6INGsEQJCkBdAwb3w6r2uiSSDx11U
i6FypPknAR284Szg67GBNQ/C2G7nWSvbeFdrVi/41akv4qMQGqss/t9EobiuleTboIjLd5/jjDa9
W5ws6SIAfbYINRwd8mWxELneiA9s+FUZfPiJsC9T6LhWYjCeRPV3+z+Z9jG884K6kwUO3cLNZ3vL
dQ6OiQLTv6OifPwe0gTEC3AqYBbwSQwhWZlkvZTYC7IgG9hkjmKvZQ+bX6i57rb14xkolKQmNuFJ
7+FkOcKnmR0TNRL8rbbEN2kr39k5c0lAfhD2Xo+4nwU1sMPdgWkc/XKj4AZ9zg3r5jzMuZBFfyCX
uZusKSJ9TZieYrIXGCnbimZhzdtf3/+OXZEPJzzhYsfZAhhaV6tcA6mFbQC/ZaB+WmpZk3vWp3a2
pPb8V2mk9Kl68XA48Wt9oovVXyatUBgpzRt73xLkkdEgqqZsINc2q1+B3CuMR8WYL1cvxMA1cOcs
fN6vPS0I2zxQRMyfdrO5rnXYY+k7jcwm0qkLtMY+e9F4uUHiVODWnVPQCELH2/VVyISWiGjBxOZV
X7QIwZKpfPVNFlmzF7Kp9f7lnX1nE0aHPa0OzR9X6VICpdeW+GRId9xMfcmA103mGxfA71lU6jt5
7cA8dsEM1V5Y8u7yYmCjFOEWj49NXh+t7fsDMNx45f7EBXvOr7xZyG6PKQvB3swu2kKsKEDhTSYk
P9iEQ0huhJJ+K6dqJRSRlqbs8rbZMWlsoBGjmQa7I+U+fAA5lifHu0LwupSLcYGckPKi//mOio0j
aV3kchrOZ7qg2jneZFxJZjXSu6x8K3gDdUWBiYSnypm3qLGgcVLmzLOGhKdSimYdAXogS76sm0lQ
6hG/ZBUOTSlDGhFKbc09F2CpLA+y1n/gvzY7KrfJp8f2sc45ICYylPAEC9vY73e2X+ifb6fhvBxh
De4Awwb3jZisxt+hWSg3Ue+rlJwSHQ4DiimZCRZ8EnCY7DCSBVfp+72BKjdMHcm6C77tbmzsOqPj
gCLvxjrJsG1cvIeWNT0eG4/Mh9mdkVyremsBDDmRSPoaGWRhK57MwJ3GDifzDR7nWyRoU7PBiDhA
LEvssLAJVRk36cGgjlNok37H1+qTeSdV0CQ+vzRd5ywhlvvVx4M/blYF7Nd9431/sRQvlIuiKyFj
OeL6jXq8pIh5AqY9eQzWq4C9zhNRlDMnWcWTJvdzAeIJrKMCDW/OEWZ9Evv3eppqHroXKTBkVwow
Jm9BxZ9LLi9vMLgI2gmZ5Nj9Dj9BxCJjcQ2LacEu989H4a/ZRimS5EHRlhBIYwkvPD9jeCPf5QvH
lDQ4GR5d8hmIBKKQQNYlqJENq8u+v+QtET3g17Zb8VlgxgQysz6PrPm46n74LzQeDn15OIh1/OO6
lTDz3CtIrlztZC7knc9589ajPHEkt2ESEVpAiuJp3ANF7pu3JE68qCl13otGvBSJvgeGxmgrnZqA
5BJ1YjZ2wiJwovbExNvQW8Qlgsh975zAA9VKDK5IIakYW66eJjq62F1jIlAbj3t4cXa2kMQXKz8v
FLCTiJHgxPtgKYFnHVD/uvr/jY3F9USffxBM62ZNGqOOiTever8jBSx8lujVhZ5gNfGpXQJhiGho
pLCpI4GTp1B0kFa5bBdQPS9Fod+5KnjWMJkkTTPS72fkwGBtrZj0FlyyygwPh5u2PVtpd9eCUiXx
23iEJ4PTHXoqnFBlL2FdjpkVGwykVpNbpj5/7HopOYQLaSit2pqsllbAYRTJkRTZzn21QBH+PKsh
e+4cCOpBglJPPi32UJDPD7pY7h+LYY6tgxjv0Q3/cH53DyqESKPNyeRjt1YHseA9pmxBMfSQKts1
8ZLNpbKcllo3CqdYMztf2h2BPgfbUk0gTkDOjgS4gLJLmQMbDGkZitMPR1lIROAgDEl4hmu6Wsjt
4x1aUBNNlvmmDuUyL4co+k9ZMd5mnTMA9uBIno1tu593/MYLO9Jrc9+IHR+MYR9jo055GEBu5yad
+CgO2hBEkJAgDgtPBP9LFNWU4X/2qq3HPpt0+X7Kf9dC7ZMIBrA3MqKAdVq0o0AkOM9U1DyTside
iJQsUlh2KD/PPdbFkieauoZ0wDWbsS3uK7pmBm0Rn9oAZiiU4yfZMWWLSGALExRykCSSG+FkMvvz
4YBC/jaJ3TLsdZQc0N5aFgNTVR5+OpM+lOmIiWprkekUQvtQp3jzeDvjq5WbaAM0yktSr2tPx53f
Ph6npN5ST6hJAieZhapdH9zbRj8X6tBHe/nPpOGgvnk7Qf4QmD9EuwG+Wc1Xmkofv8eZAX+RcxpI
mnI2lF35IZmHrKxxNXDt0SOIb0FRvDuHKo6IqUiX6bN0Nm/LByGaT1LOHoLhxfLdEyDLj6kzqOad
3IICycCzQOaPegW+EKo6+QHj2Fh1m5OuTl/1tIzdHVHpd4f0utwWylNYRsJfy5QmAUGtUugEXo4D
0SBwTgBcKzG1jKM3GZwkJWHFx1XFjZH0+cGguEDSinN8cSKeWILr/A4BjJ7M7imWXJSf3KtUXp+F
podI6M8D3A57T7FZ8jVnA7l0IvRmf+C7VeJOf3GHKIFutNgLH6881N+IoDnvWL/Yjdmyy8IDEn7J
Tsbrd9qzubeyQYQtC4kSsu6gnSiP9/HNTGP8LXBRQNvaqQ+bKEEblrRvJ+DpstnmH66w17VBfyJk
jA30lQJ52oNw6HT30FM+cXt0NHzdE/ozbQ27KheJsQ2DuvDUMaEDy7qnC6pP8fMqKC0xTjLCOz54
ym9xRXA7hxp0WxNWRuXboAjvM9IcMWtfYso96DxbPHwGtjETZvjysN3GKRoGaEjhWL0we415f7tX
SeLmqUdajS5VdaNrCbZBhNLAae4gDQheF/6i66/340NXR2TV3+JBCzMLm6SiBUAP6DdPH8zEtEAy
8E7vDArAqobicRh/2ohQ8ePFJ86RgkBQ6yQ6XcOSgqbUQg2mD5Cht+FPhcKy1Hg9r9tx1CJvEcOL
Toh/PF/fey0+blXU9aMmM1Z8xR9E/gjh5SazO6QFfa42rSMaJ9Q7tcTIbrfJiaUDCWtmknlfGgJV
Vsswr06sIrauDdtJ1SbCm+Gi+SjHs+U840uPz1YgjLxxEFYzLEBwth10EkScQQPlKj7KMCouuXPw
n3b6wTZbwL4VZhOSCfe676HlMrOv+Cv+hmitrjqNr/ZdVJ3IblA37LLunYF60awiSmhrdaBAs1cA
MqMh3uIVkbWvM4m8N1k3YiMWGG5SWrYAY11AT44nsk1d1kb8AiG4NRqsCS+3ioq6Kj2jsjDgrhXb
77huWvQHMcnqrbi2AUvPgweqGpCifbrHsWAHT2lXeHsxu0dvY0IpqMdcTGj6tMTUJ74V7Ra/oXdm
8OS6f7yzWS0VixHu3UwMNsFQpXNG7aXsem/AgDQK8e4zhR36cwJKRalE3lC98XsPoLvaHCr256ie
Ez9sb75TrUQVGJBkgtCBx7Ej3PuC/8u7NnR/A8aeweEWXZy2W5L7dMu+UglH8GgLBp7JVZBajP6N
eUATGMYBc5TZD3ozPqQvVXudhZraRHu3n4Ow8O9NsgyUCP1mDWffFiyK4QFqVDjHcIfBXLFsQYSy
tvchhbafOXZmwD2dCB1cqVgrZZvLKdck0jAnhbjRdVJV8tmK6BGr55Kqm+uU4wWGNy4ZXNIt/iJ6
NY3El01+KwZqLYl4xfNs/1ay6Ln+fcu71zEvlne1wGs2yO40JP9tcmSMgktnB+b7OZDJegHudz5R
1PNehNxF0bQNLcO1XqHvLhbHvnZDenItz8AZCpqajdoSz9EgINLm5EwFrr1DXItuI2P9s5uK4t4Q
TvU9WW79dIVRQkaYlwpQGmJlEA37pUjlFUgvVP3GvESYxhe8qz7FrndiO5zt3T0zckMvIfrYWKiD
HeFw1M/ZQnPZ8+JYBHn5Lvexet3+ntwTE+7HKVnma2T5sp6WLaEsofW+2/yaraQn+hWBi8+NGV5E
sa/7tYs9xbSwfPrvyGwRIXNX2fx/LZ4AQo13pCB4JtRRc+3YPXpM+LtV5Kd5vderNLBEd8G33jCl
g04ZAtYKk0sIE5j3EK0GxS6cr/YUGObYRqYVUaFQvVXMoKEIlpxmvx6eoOKCPFmGOg68QXPC9mIq
YskNvi2OUFw3FqFV/IA554U9/o4jgUVxB0/w27FZDwICQSIHyT2hOcgc8jU/1gkuMfk9nOIeYNF5
Urx/Pu3Q5K1MrYTmZiA336y/QF1O9rKzLtusQeEMvYBFCPLA46xLAluCEy4zVJJq2RzXg13ror/x
vYY+LKaiELu5VIO4G8t/fetDZWajuRZRZ+TouWdWDJHJtLewAsBgN2fpeB7uRnohLnetRQJFBvGU
fV5LeeutvV6oeRfntU3KDx6eweJlxABJqaodnRgVDWjBz4nDzVTO9CUgZa1Rvd8hmOXIj5H78gMf
sDHOU2tCYwrMGb5qGQmnVjjGzrhLAZHOcat0RZoTvBrWjL4kp4vPBSmqi5Z83ksYhOarWRY3wQkM
KBCKM+jrIxsOfD604r1iFkjaLVG11+SpCTijKmPlmfEuT6Mp9ziNvI9AZktHxRP0OtmaGENv5KrS
fHghTCU33NR/086JnDLDcLBqCgb2wYLnEnCe0iXtl4cz1ShU5Pj1dLzXLDVO3MnHqJil25A5qPLA
+mDxrJ0K4gJW9F8MGc7GPBMIcR4KgGaZMJzWpIKF4TuNYizrZR+56jhPBc+NOYsBrcrtmQ6FLN4C
MgVswTOvlGlFRUqbLDbLPYDotsrzU+aWHFKstVglp7dmj786akT1zydUBu7y7JeN/yR/9rVpzdWy
jLw/pb4TFX21loqKjfSrpUA8CunVbnEq1WjPcppA0GjeCNsQ2q0Xc02PBt66wUkhyekHm1gc7uF/
gn8k8fsqPc13w2wXT/QwiuR6prJLx5WAwuLIx89KiwUBhZKWqc5YKEks2xEYbVVfYZiTt+aQzKv0
jUBPLJSDWOHA7dwiLXqi8zxnES17K7Hb9mLupfVdzUJ2p3vj5hhPEID1HTLqjgPieQ0P7qX+Z3Yw
rmXje613XBIoFNhBjBT3EU4VroF80zaIXu2vOQ1A53AW+NoqG848AfSPnhQ5OWELQbZ3ogl4BY3g
PAniONZ93w+vYg/1PmeHVXuwHxHMTv/+J+3YBEXDpv3wOFrAk6+K/mWDKQls6/teTlinfYO9FjEL
nQKUUJyv5pba2g4QtjZlPBuO56/DIZ9pWtllP8e1j8ju3fq3j/nWE/76AfXO+pa43qr9mN0FoIt9
TPIvmXrdGeqjK83S55X8YHWj/OAfs2sqKaYoXbHl82/r4aY1bc0OLf6+qX94S5yAxjlajuuUy+lc
OfNT2hfh7osExLjFH/tVkurpPAxJlZLAhYbZgGU9n5KmaUx47lJa5MakOwglLXLs46pXyk9jzDra
q2w5kPLi+nib/jyK2o17rnXYvgI3sWtex7daW7AqPDkPYoRA8vqKpkt4dSDzRzMNgpFhaEntYRTu
B0T/vrEVy+g5R726w47r5jnqdkQk6ImAPMX7os10tWmZPhIdjm25wwfdIBDLgFEFs5oqvCEwItS7
I6sXLyWbfAzW4xQy7nu3r9XwPpqfZy2CNXjbjfe9rN9s9uq49RdXaD3IPU1eokGUCLop8o6vBM1V
wZ1brQ8pZ44Kz1/Jjj7a0bIjSNgiQ8Wf2MBPN1CKSUtBJxqISGsUb71Gw2X9DtWxuLbXC9ARi1x7
yusKuDzP4dv5EUQGGW8450hJsvywHsmrXHJxD93XO+G6FLJ6919W/sS5SP0UhxGxGNrPSbWkJD8w
fRC1vuuT74dAn1LK1RtQIC2mYuiuNzDZ0ygmm9pzQD6cO0+QbIToDUR7xWdt+ls3W7ekFhj9DVgm
ONRfqlyIniK1OKJe+T42jLyc8gtIJLrZHyQU5Jkj+k0eyss9jbe41lADEx7y2GkCFTTPGs8jEkop
bFXRuZHb7NMSKBOcYh+hspZ4WGxDku5kSCNVGl9DCSYdtR9QA7SldKmZZa59XR4yQ+1NG8D/rTwr
pBI2B6bBoSNhzeselzBb9H00BuIeQEmRyyxDL+d9iNqkAPRzMxrKHWvBFHKHgkCU7tYqFldRgHeW
mXaf+G+6dAT47NodAQULmlfIfMFQ0f62hw+FC7ZaU28AoUEkl8D1mY9CSCM08EZhRPrO54TjqL1w
n2EgBuYF4XH2Ffy9W232pL+MLXC1FblhkM45Ui6pXZ6KyQGoAOV68xRKshF4YT3o4WY552F49ekG
fwBOz//PoPxOJgdJve7eoRb5M6BxloeYPpmlMzf0RdhLRG7QOLDy/ICukGHiwCew1H0DAReWAArJ
jZ5Jz7Hc9NFlEn7aHpa533SowdRfC6HnKyEyAIOs9MvroadwM46cGUXKcpas0JIpPSBL7Vn4kDOL
7OZnoRr/4ti5lrT1slkSGTuoSystodMJAiteEMN1cVNpYIoXk3Y4olz7eojOxSR4+8Oi6RUw912N
XjFEdZf6eiH/33mtvaWxPcCWYFOW3wnuY+b2oCoX0l6OEjEoFj7kVS7qFDtsiswaEKHNibdVvzFA
V7ixLvSZW9v6nMl7xp5WRT6Z1HXapypKSI8J8WFgJoXMv/aNJkRMYA1HcN4CBKK4wFznUUeTIIvK
7BhLHYWJlDE8SUIUjk827reHTVbses7QtUACt4BuuU5Ne2OnZvafhjszWWNxZKs5zNgk0CR8BVyK
wTQAFXVkxI6ljGcZRopk+OXuC/rOxVIWh/uJIS/7AqRQsuUezxWihAmKORx/qsj/gxHK7ExFN4xc
lByO0BdeBGu1qZ+Y7CkaqyLfXg2X0fCJuz2/J9aZZwx34fDeWpFNJ4yTsp70fH3O7tfCtVIDiLpK
dolSno6FBqydxNMRgGDl4fKj6VH9nMAbMTuw6fZ97/SNUPw9/ZX6TW8osIgIE7x0n/zsT9qqnl6r
nXIRbuhaJC0ai4ko/BpzVV6Ly7StzjWl951SCPCp97dtNRayEeLS7SelM+piIU78cYndlGoojem8
PfdlvKdwjqX8jgPBp8Z2WclL6Lnzw1c3/mHmF03eBm3NTeyqNaiO4YBgQkvJRrnBnAmObHPYfW9u
yEEQqtcjdM1aXFxhO6B7yjCI7ZLcj5PQD0VoxlAqT8yBREsqyB8JS9ujx/DoUZaQMnokrkvvaRI6
HM5dFKKu/vzy14RTTUvcz0xStqYb9lIFbe2h2RQkL752bylA7NS3KYaAryCALgRmJX2lhquQsF9W
DTdqaYL4egIXHEod00PCXkRRBvVkvEa0eIIWiWiKH3T+saEnekLeeTOzUFzguXLsYWrQFq3i2t5S
zevDhNysgZYknXb18XNMbptU+xieZu1UgclXtwsKMWLk65CrfXU/WvoduodstfFHz35vfEg8AGp+
8XyRIYY4BmHmQVA/TmUBKyh1qfqf68mkUFigD+Iuv+NTfc+g2Hz5qJ9p1VY9L1vsxwHqFbj5t1Rl
bV7kUq3fS9jhA44FGMn1wgLrqB2Ag0EtGkFNTMyxaK8MknUGSSjeSfBAh4jSnX0qprVBXCBoySiK
OmHQsxgAP5Ca6tOzsFikik4BsH2Z6GTmbJWof4We600jaLzJ5eTH6byOk3vRd/DdTzaHR1v8yOHg
wTci/Q06QdLzVbNsUrku3JqTkA/RonB4E63YLV0mMJPj+KwDpKqfnnQtdBfOlTF3BQX1P8SRPtQt
N1a8XITRXUNfkepqnScZb6HAepQZQbjD9BYJcMc/9X+7ziTcgFOIobLZRtTO9w5M779A3R30Ux00
relmrNDa9Yt3Xhu++jz5Y7KImsIBVxgvmKrXX67KmvBeXSzcQNfAJjVQjJA6LwvJRxNSQqvqh6lp
JiIjcLtD4FU67vuXo9qcMyB+4//I5Zl669Q7lYtZFG5sUWBiVjHZcOzmZJ2KdkE+fBqutzFE0fsG
eWWU5W5ZK78v12rMyCONPOaRViVhR9FX46ceogsYVKWtAWLMK/JpCfuKJnK4KHNjhQLdOK68DnqA
mtCVqtbrnyqAV2qWemXzRn+KdN4sXCYeutgPgevtIxucKMpCnDS5wmNblnztYjXzM9i4DJ5GakI8
fP76Wbgy1PEtD32tUWvYX4vqcn9PvIXgLLmvJsb2d6zDG6xGb7DXkAjWPbN7BIMXXAyI8uPMf0qA
NjtFW2PsTN7YN+kTL3Z+mQ4Ya0GZ5FlSY67K2xWHc73Ac/ZIb40omtCxeYQn5+ydNTX9YkOJSzFT
+RkmgHdxRFdqO+f9vJLOW1+qvFzJdswEDsCKQYXZ5umvOPLl3VuLYvDZsE85xQnngV34A2jdtnMS
aQr5S2o1eAgA+D1CB1FuLCaFc9sywsDaeCzjgerKKAUwvyG00jp69hsXqXjAl5QU53ZAcgqaVf2d
opOZcWqRDwlz/5tUxkDX9un+tzEdav5h7KdTgqj0kSWTzNw1nHlCvkfiCQWAFo/Lu8FPBTI6XBWe
RmuKlcSKcSAjE+No3zZRHLX71pyKsM3XKKtUqLk2/eKLMpYkQyBTixplzefUonzn6UUZ/hNkVZfP
iaqs2brzIOhOeUXB4+IJre2U4GCSw8t7/JrWPAVrzamPCdWtC3S5V7ypum/XV7BtsKsUD8JWbMwV
dQ8fx9bGsu6TPPs3Ikx0JZLpzwknNkzLD7Wf7RkKUGbPGqSL0peuhIqNMDz+OH3lrTj13b/q53fd
SVSoI0dwTBHfkH/RnCmenk14CRVoEFvLzIVdshCa4GVNQ7hzmmdKzkJomGlQRnVItSY3J5smyJFE
pRGJmC8JCXLKq184CoX08tp0oJRdk2cgQ5fn4yFcgMpMykKP0IA/Yg8rMain5aBMG/NNJfq/OuyQ
M7j6VBV91YPic2k+Bbd65jGGxM07hsaFY1YEl8rpk6Picf1zxmuNJWeIFZ/ZJVk548LO3ZemQ46E
lRaeFD7Ms4r9eKeUxZUuI3Kg+T3Am1zr+g0KgxYFQ6+yTV/8cvJ5RsEUHBooXZYJAc6NzSEfKDYi
DlVYmJINKf+uk0t16mtx56PA7+pylVL86qUhX1JD3Ny0nGMD7E5p9W5HC+P4Zuog7ZcSweAT7cqU
gHSFSUKd9tuA9z4LbKQo/zKPHq/3972dZ9Aj9EvxMkaeEddFmI4iyH/zrXSl/4JQY1d3AbXywRvz
IWjleLhMvwmjj55ef2tkLFPGjA3SUp/e18RkTJNTSojoUsZC81uAYx1W5LXcTEZbTcNgw+Ig2J6L
/M+L6pUi4YZgWUndUOB1q3IL/fAfSTZ9a+sr5VhpLtr1pD/UiX0oobA0kYtB1nSYmsvEAzioDEB4
YhRymQ1VsAArF21wHQ2bxitzOAn0pmeMqQomysrKb2SIwAMdjMFPcWLTgfWanFokSvqdB5d5m3yl
J+3mK0WXFAr16kPa/RjFlztYt8seJoZAHK7mu+n8QOI3DxWetDVSyAsfSiU6EFuj5Wm+Yp3uaPek
+LzqRuKsYQ8oIM+JEptLn1xMx1DYyRVcOhd9Dzs+bFfiL8LYv7VK98uEEm3a0CWjuQZJGQVAN87l
O4KIxT6znAQD+Uhyvw6Rym1GzNm+onpyKUwKd2VrkqjHm3u6I11C3NW6nXvkwZv1RLVg/yKw0ZXH
BzagD0QUu0pjIl7BB+HwSebHD0OJX3JeLL66NZD5S+c0YxINFdoHjB/ClVU2WwTQkNp1MgYU8mMV
2msZGw4sUu/7xmwCn9yKBDPb3jxUuzBtxLHZPfdnBcmaVE0oRHVDfFxJvT7fgTv8dAD8JwSnt3Hb
g2GSVGiwF57XmK7pNGZ5UfI/WCX+w5tD6CyBqq4Sir6rV+nWiiilu18qKFCHKHmXAZLcJ3BZtvzq
/UlQ24I0UpDkx1XlgKcgqkp+pmLXGNxiPD/yc4UdxIIGTHr0TM8CzedSspUDTFW7c1mUlobQpFSD
+AWX9DWimvYXaxvb0TIzBYwRRQRjYPHWUiO30w5HOJttVltSvlyd8x4IouHIi+z6QHhuQW//8nPQ
62nj13Gfzg788IKirUF3upMquSWWBSM5beogh9tm0jJB9hTrD2veFhhjEFtdYLVgHoCSHAOLG93w
GFeXGRmG0rd0/C025yQ2kpYzEi09vkXQJGc4RMlVNIW6qWclPKuEzdKZ1ALOLcpzEphWNyhjGyuP
PtXpfmBOXpEo8BMfFL3xuYpUJgd0qmU+KlNVtotku9B5eS0pG3IyDOizvXlVO+sq8HGxJ2yVtYYM
iXrmSY3NHPI5z7cMFweWOusW/1HanYlu8nqmR6zsZgsydwCtrHsCcq9O25vaPpYcIUFdzDo9LtQb
XoB4dbUdqNMgllPO4LLJ2ZBbwex1zAajAtySwhmJPjpiGo2aM/OM4Vqa4FNGKABhGI9SfJxXxqoj
cAyj8FU+kLrugP6EhQktsy6ddHowpGkfkgvahDqc8jO3shNBy00fPv/IIBu4piQ9se217LUqTY56
OZJA7/XktcGrESYkNlejoMWx3GtYf+r9IRDERziMsz//CxPnKjrD/E0R0z16BpGqI77PzqXeDZTd
B2Od0VpczAmeyM8HVSRtNEyo6C+lrQ5cFuisUfDjFTtTiB/e4Trj9O9pgjbBJ9J3GrqRjL8gVgNQ
n2igcttMVmxdwKDGnqfWumiPT1bdlCBjZDwHUcpRgG+VKJ2ZoRgiU161iLB3PfYprGi1w4pcJIjF
TSXzlzeEnD1E/DdiCW37+nyUem+52dtvbiipLsGeIG2sjqNjC5qA9/t6R+Ym8dU/pOmagEwbvWDZ
ky9CEq2uOxhsYXLuNe4INej+ULR8WU4jPtyPSV5ARpnNfQMqD8YpTBcCIaWT29KkTN7U1eAYRp69
UQ0MKsv/EuToNcv17ifIpUYfcxOreEChQkXPptBauIEl0qEI7WF0GP6SAxeqhmjBoVXI6R547tXi
kc6xQsdYAL3W9n2G75Dyv3dmz4D5VfoiUTsaQmuwXE+DbBLEOILjVV/jmEh6WNO5zqfKS+3DzkZ9
/W19lLEFU4sFxmg63OLWP/gMhJtKT4UK3OkFxztW8Iz4fuhN75Fp8+N1e+dvpmZ9YSFd5C4GTVwn
QxFgAa6PspEiqBlqpaIkN1lcVUZBFkNLsgx2FIO5sT5CsDSP6W6ysfc6lOEp4IRInji0mqeHiA/0
SpSElgsaWc5Yw9tNC4z7BZNmIkKsPRkzFniQ8rJZibQbf5OvasUUQMPGH8dAwwILeNAEpVQzPrAr
WdS5KbLoQeftvA89Sq4tEPOvm2DAbvMFFmiwfjkbWT7RBwwFYayox234GNIiP0uBic4HiY8olASp
GAcJHGtczGibv764uRv08dhZEx2Q1DEhkGqrErffiogR9nlbHz1wmHdvajJdEHdlFnJGBCjHEqAk
jehK6oRBHjwdodGMo9dE0W+f0y/BGSY/dAYu67TjRMzRAdtlHLtNx3F/Mo3yUZV+ElOnIiJwsL/r
xqTDYTDSP1p8jmiZusIUU+JrbV2JKSGb/X3rBzhmQ+Tc146fsBsXJFJACcoWauj6KwPbCK3i90WF
LrtHFWdlnWS/73abST6bJ40SO8OeGa3HH8R+ueP90hTNzKDWqz7KcmRrWm+qpxd+MWgSV/76dlXg
G6L9QKcNsSU92RSstmn1J+XTBec3ltzKOHZEVAUqDKCLv3IDdyPUXf7gjhbPlgKviV4o/IBSAN1b
YU/00lh2twOtF77K6wOunmB6thmSL9PL+zGy9p3lN+Pn+cercQWJfzFCEXSUAMJkCy1oMJvKdLGA
WS6oHI/eBIiG/Efw9dw0vGIFiZC9tQJSjYtvffXTUPkv2RCjZHhaeOqv0NWfniUpxXkxzJ04Ncuz
n4RW0oFn3/5QwqsTFrAT/jUmbTGmABkicrdbPdMK0vvINnd4N+3rQmNWbatdbpAx/iANs8Id+RZh
1Sr4RgoqrD1vB/pmXohX6mwkUdhKY70p6ZSSSbMHze6k7nS9puaE5iRN6MmlCA9eBNsPqWVER2/C
nl5bulX4jyYs9+93q+BVudRHEvBmkwWy1fYMiNmfgnAw2mMoR0gFBloRiDTpctxhimyL4ddLvM/C
WkVp6NNHA6O14nQdY+xOkUdlTaH3wqowatsC46pRM+ovuSNaKivMtQym12yd2sEUTyV4bjAdzd/H
LI+oljBKE0odqjfctUwOwY6FGiiQ/iiw+4TG26Ffrtyad4Z0nyEsLY/8U/7xD80qqucpfJPQmMPC
F7rI0dJRUo9BMBmYeU58Ss15N04xhumfQAPA1iSrpWK24KhP993pE5aumz2QBwiM8mv4VsJT4p2+
8Q3YmIKTASd1AVA0FwCnhnxWBx1Il8L5+1EwnA3WtJqirl3KgrHw3hOTket68+Bk4tFazHQf3Pz9
fJGW9PpBnHzBi8F0rDVavfzgpTxlp4A68FOmTXmWy38Vbx+4wnhJJHYlyjDDQpyr95PyTGLU8pve
JAPUoQxpIEB5QfMbKpUqMziWAJtXkMjB0XdoqOLgfCLWbTMgTJQdqyvbatse08JP6YIGlFce29Wo
QTUGv+ydYSCn57K5wQCAmkha9ZCNVwWR29VEfwifGDGWdNH4pmjlKUS2Ph4u5JV8kr1+VmGHWCUS
+BBasd0gX440l6TdqFk5DnsBfxeHyTWgPKYBziARVH04j5Xc1X4rhQ6aKVnU0VUsRzLekPGdRDin
aV6+XgDxrFSGUupS6sCm59apCoRKLW8ks6Ru4t08dfkz0M5DoueE55l/zVardcRBM4KsW8TKRgGR
rfiYLnX/Bv8dnlXmTSh4Fx9XXQ7BcHxMaeVZd0f7b6qbEPEjUvTxdoZE1utw7kzXFYIVQYbJ2/Dy
ttDu6bGupOG0yFuiA24HQlFN3bPhA8W5lBMWY2mguWJOJZW1OTaxJdLbNe36O9DI/l9a1M1GmkZx
IsHK4NRoa8Ui2CUdTqWuNuHC59KqrF4m2m4BSC3HTagaWrcz7zEMdIK6hswmQCAaihDjDltdaLqs
sPEd0xLJwg91ymUZlYQ+Z50y53Dtt04p8qCgLgb0Drub/DSyS2F+ikhfS3upMkDrxg3uEYqtX4gZ
p/yqPhM5DBAHfgw20ZK8VlJ9YW1f3saOtXZCirorXNjHDUJfB25bt97wQuwkZESVyOdGYuDvN8ST
Qr1MOEAwyyDCXtekKkhCUwVtCrJZkBtJoJFTJINwUhkqwr3ycnjJ7ZOhPMGWmMx64oK0y2XgZd8T
AXpZXN2pgPW1rdd5N2yTxglaYLweJRJX90gAqdxR2SavZA+/vvtHNb0f8jsyGVaP0E9pWFvUsxmA
6hhtu5untZlXvYIgu1SwwAhbvYgskndL3DT8PQF/DdUb0pRXRlAF1ImhUr41JsDIa8rGVtJUXxbM
wk+uyP8YXE+OCv4skoZOVmEEzMM/7acpDn9xEF/ilytHKu3skbvQ2DXfli5syaz+paAdUhDYzTRa
wPKKV3cIKL7SZP8l3sT8BCHZi6yZMFv/IdrK4QKGnwRyJkZ/Gla1L2pC6KKT0OB58Z4RwoGBPrI6
47dqDSTZ6S61ug4ccK9Jjz10atpx/X4fQyJaC5MhEct1SgjIPew1Wz4Muap/zBsYy9uQexVGJl+X
56/udWUve3fZow+wv6qZl/3ACO9aK9IrRGSwUR3rTakMhrJEMuSH/YEd9J4ipnUFfOMBx/Rp/Jw/
+rxSAEiQUxXYz8EApcClqgmdGWGTf803AbAExI33LVK7hGWSfJabVK1QK0BT+Gem9kFhJdOoxZvB
TedizCoCPcw09KubfPteT9tsClWzdZoLyo+JH6+F3ssxdM2X5jpcBhag6NmhYcqnXv1lHdVB4as9
X5gwG5SLECYQsCOq37F1jkrGbLE5jlTkAWpvI3BrK6pYflXu5jUQEiildLlx8zW+3Zif4k2dgTHg
3Anpmzg2lQWUkqrNdjAzrBTLiYa21hnTdkboWaDfPispPWw3+flOQoXQIIIrOM1bMbLKB0lE5UCt
TsnjZRepQv4rHFCzlbXk7ZZqxpdzzACjXRyWhwZZ2OnyuVqTm1wsOmA9OvQ7Q1hi4TtV0ApaC1Du
knDpp3yCj7UMiliPYCBaBOoiYSJqj1cgNwXcJ/n7Yu4pa7yUG8BQvthZzX++j4c/X1rklurvBdlP
EZc5n7rSciX6+O9CSYX0I0k94wGS3VUEn3nfL+pvNcVzx7TLkObGfS4hoRwptOsDhDyrKOzXiqFr
pwDukO/KTK4D+7lsbAXoAYnwtuz6kh3pgngbXO7or/pWFKmFYQTtblh6VmwoQuzAdgPnWG4kRdDZ
Uhi9LEHFbn3uFppLu/cMl8lLNh2pWBu1CNl8Tk7iq/zhhmrCFW/qBgU2k/15pLlntVKAq2uVfOoF
tVKkdgPylqhWH1dnx56xea3ZteLc0jPzPzF1gb5A7R8shrLnGpVB3NFidSuyDJV/fuwtgHd5rSXa
wpwJu2L/+yvprCYoze/UvlKp0ACbLClUXA864nTe/l/TZiLKJdW3S290cuoim2U5lC8aMZWMbpdC
+Cj9hPMOASTLc9+6xJ9kKMF+zm/vC6rAL9JZWoUOng9rgOAiityhjqrn5sZ4uwYNepdEaUx8nMXk
Rg+mm0G2GtX3PDm3BiG/GqVdPXozTITc0YU4ubOk6jF8PhvNRXHQBaNz6//BDg3WK8e8Zlahm60F
ybzDQDYKg7fI6PjbW5rWYp4ePXt0chDb72XiUbEtkKygJiuxEx0hNEI2k6WkE4VgUjESSgAAa/sB
4PbQxAXJHyPuYcb6fcFSdYbMHQtOr3xYHLRuRp0bHAV2eI8G2zv5MjZyHRsG6BkQ4ZQjkSxDXVSQ
LVp1nTGn+5TV8VYfRXF3bRvU+WSD8IEHwIK99asTGgXkPJJXYNN8p99WpLk69N0FUZsh3uFqPToM
7RpaAiG6sKTiFilagYeHKuk6uu3121aiHCJX3uRYYNoSOFshC6rTyOM3U83Q7D+G6Odinp32pO9n
VqD9h48nY+lG2CQPYcmfLzuso8/XqsAZNDk20GSThaRh6VTQhdxKI0/9Wn85nH52KopiUj0DtepZ
UMGSLk/xxJ6DoKTHZEAUpC2DFt6rV0ANlCLBGkZS3WCXbUFkmv5E5pxwnQ2KgFk3oUhZfa86VHlC
HvQnPP5qvh69O5VEsn79r+sIKYwGrvDANgTDKPTd9X+r6UUiIs06sZnXvUkrKfcLodxel/7iGS62
uJZGw3cx1HM6o0P9FcDUsMiwv2tg8NHoG5THROo340Zrx9slyDOdkxcp+hkbBrv7MaZuibAIEPu+
GB9k4vnD3QSdf+lxKzHWdz1ye33IN2e9jBORuz8qgaHwOIrjZiYShdTPSW2o2slAjyTbQbqLnsj4
SCwlpRZ4MWDFcPW0xQ0S3xL6rc/9zCTvKhrQJRWCtTGjH6PwpbcMeLd9RK4/Hg2SVfVJlP6hmWLZ
LZVl+1tqPhZPz5LAlr8Otu36ge7tJWx+RNw2iBJ5l+BrB9QcjtcoOVExHy87/rt3OQv1vxbJx7aQ
UHEmqkz3p0267axx5u3yU+1/m1vfJY5ORslHgEPX8HbvZXtDDNkyyJ4LoywG1EOTO83EKkEz6SsA
3fmWVmOutgdEIE4fi+YhQM9FuWZRSuhgn2us5gMUnV3B45PDajphec99FtPKiB7DIUWeeoU7zvoS
/tcF1qofTOpWQ5OFh9GrYytoGatlppUp8I9SRggTxVirFuySqbEPO2kTnkBrE/1hLjyaq/3pWhUq
QhPvoOJLPJskRL3itk87WyMcRPmFxLDw5vS56Tzz0OIp8gUN210sNMHl9NwXXvKcQCa7j26uNn/s
ctWMqLDvrem/bZb97VAwxH5mJTcwYvu17sTBafNiZJL2PnYEXR+6b5rnmZH5znD/ryoBUCyrTE7z
C4HWuFcoJLpBTX4SpvkgSFAhtecNZnG1Er1medcQaO6HGGq2O1p+lIcvIH+KQdFXdobk+9xFiiFR
1D9jB2qXUGoxJdnjc9n9/ZQB4qzoVP4cIYdRAwCSncTKdkN26AmT6USYcD14LPC3UG6/wQXbzeH0
91U44l6H0TQAdrIr9jgumtQF4U+YNSo7ErmERGQGCHhxeXeI/9eenhMT6PewCSzOGieNS0N0svDp
AB4Xd0MpiKJzyBNq4ORDPkMCIz/6xOyMZfq9FHIUXxQEQ4Fbdhr8+jHw8LOIww8cK9hA1mE5PYPm
KEnDJsPyrSQxujoueeMoR3+0rOqj2OkcnEvXs4M5zxE34c1Tb5a6mqARO9i0+Q+l7S6knFl6+NJh
6cK9Xy82asZDP4Bs2yiM7sYVSENiuJ34e1c/S4KJm8C0Y6sWV8KuaaD/4gsB050Ump7cKHodntn8
NQzN36dICyK4QntyP+sa8N0tjdwP+xKQCNYpN3ODC0ZsY4aQCx8g+dVuhmj/3OClrPKb0PeHUK7k
OMv9l8a+KxzSlNw0e6l8sxa0OYWcLx664VJpvHNjgFeDne+Vsvn3oKbxXjcJnqTWdM7faj2JQjwQ
e9sji1busUjP48TonYgY6TC78Oqwc6YN3ubkAE/42jzbzNCj8fKvg0IchqJcXo2wH/nG2vlouLPJ
vVlzUG4c6MWWeEyE8YiF5HOTUUpZ9UePDXDQ+wQTEpt7R0Zq0yNznHChpme6Sb4t7Rc4gODRV386
kINzA0+tUcrk4w8qz7QHKW876gzAGjyHPpkKnj4ktDbmVXuFim6mjbro4u7pPB7boyLNjjOLcLBQ
KKZCWLnQp2HaJlvrFWtfUdvnyoyrGRC5ET+r+FFgrGa63ggQnsmcYFDxNBQQcU1ZYue8ykBmOjkR
tcNHNTFkN8bHcinUC1TmqaBnIsgaX1DaURIhDIPLlmV5b/nu8ZI0eTqUpivo2099KjWjoU5TeL0P
T+/QPZJFlIgZ/J5c+cR7SHIGqQa3UWEFx+REAScmiVkfeo+Xzg9aYRlO6UWjvejSzWnIXCFBwiQi
up4ZKppAomEMqJwcEF5nUSRi6BM1EG3RXjfq1PMmsu/HwGzeBRSF4wJTXcar/5v9A0u1hmqAtCSJ
vSkDtB3pynpA6ZzvLyqSQ7zD2+4y+tDAutSUIXx3kWHERUeu443JTazdHgFEF4QjCM6sg/prB4PA
2JAEnSssQf6kldARSGw6dRf6/BjJAaHBYrrrqhan60Hvva8EZvuhuQouudYLQY+kuG82H1fk5ZUQ
HyjW7he0tCQe59RQ9IbTzvkxr1cpVwleNFqquI/wLuslKPI3uQzDS3QhMRJ/JxyZb/NxZGesXfO3
DLxRArGilGgPcMAUfApM9tdF2unxFZIJaf2yqD95AMvoaj90U+9yNcdyHTZv/XYswhHI2EEkmlbS
hXyKSqukfWp6zypDJy6UpA/0ib4b/wian/+hvSjn9k2cta53Zkl2KGje0RM8upTCk6eJbI2nToaU
mHzBemTetewENrmcRRZDlkGyHvXtFwE8keBb2Vp4uUZBlXxTnw3YLZpFWL+Zyn3Y723y9REkH6t/
z2GvszXtV0B44BoVO+3nJwzhc424mqDcHLOtZ4zTWOxqSRHr08HDMXURre8jf5JvDBKG8G90GfiO
lmH6eflCzG7yyH5Lq3SwZJspTcH2Fnl6tBzopsvlJbFqVORT7Rmpwjm6wRZwvMyQ3yCDYTE6w8/3
rjr9NTgqDTxvJZC4KYetYcfGkOjcDHrovg/8Y9lI1JfLwGLZPcrWtNRAaD5Y9UN+oZ+cys+3embw
273er2bAYeHn9cb45NT+npYlN0iNuns/jLoGwwuHiZdYKKO+Nnp2ra3QuhYttpM8Vk98vqmCCTXY
Y23dv2Mz2ld44WO8so6v+lCRXN8X2mJrGbshE66WQzsEVTb0kyWnMJvZs5JaMIm8HBBBtlXLbXV6
+InlW5P/yCbzsJTV/68r3q+8DBORHHa2pCZbZxDhQzFB61NikzgbUFMEWJQ6svp8FoMiNecgmKNu
Ix+KpQoTLrfP+S+QMucPcrABn7eA1FwvFiUS0o+hNbhgYWPQ9KZMj3jCk7nLO5EivrQJqZxDQdPv
RPa+J6juKsCm7SiRf23rtI9ElCWcBzqtVcXsUgk7d/w/4ajmWvkXzvSJNFVCcVD3Jz0s0vZv63Q5
gWFExclcoU2YULXxM6hdvkDN1bPJrJunBslyzPkIPz4TBuuCLhCbjF8q9XGksWHWNHzRKQfC3evR
vLQyjJYoP6dsQ4liId1hGpuLvDi7UhJraUOK4UEovaScTZIwwGYAJIN35f5PbBtuCuVG7P5S2Upc
AulBs8EFVZ2JCwZa3SkwWw881SxcJFkTI7xnz4FMmGqgQgYdRQ2MVaQPFl9BR6aIu5W4IGRXMEeD
yDJ5vi8i8tmgfg98I8e3Tz0sINkxXj4t3hG2jFWgzYOXTFOk+C7pHku8hN0isZonJTLcll5IwDgn
xBmIEVCaTGawmQcx/SHSHt8g/8VgUKe83cq/U5VjPM4mdeymMTrL2P/CLEcylzsCGmNYj2P31Suv
6Yl6nTqpo5qMHyO4m0liOxRfGAn06+zBLFdfjbmejYwMTW0MbpoWkTfucJfbM7Bc3EpIyJTC6Z4d
C1rbBWdBuDRjQJzALW+QSZyvKqDglwSp/dTxsrXegj9MOGOe8c0bvw7uGbALeWK1UuCmWGPfoVQr
ZfvbIyuswJ6JY/XBNPy0PMWcUzp1NJDW2I3rY2Arhplz1OaxNJRlO07wKCtddf2dNuSXINkLjnK4
KfazLXmHtJ0VuPUrbxk0PCo2SI0HnSouujOLT/Bi8mj0mn69SwvHOZnXpv80WrywdAANUhZVuqlo
PpW2RnNzt9xQnEc3V/2l9s+i4tR7IFNzoSZqENnY2KjtdC9rvo1yKHAOKMLfinCH5ndxiL7MStZL
kCflSo6ZrVLd7HO4KJbhJhPmsCI+h5KT6hiWJFKPT2mqGNu4nDBKsIv5VOzow/mdwV/kNCW5ddnB
ess3tN3CHrEP2kGQTsHWpegcwSBsCcW/XafLY/Vxp9SHxKehqLaqvNNPB5rqTsneRAAJuhUDppkj
FjlOIR8IesBtJvsY6e7xfMDFvYMkq0zBha74qXMMYtt9GsxdIOmN6L3odayNZQoki+GdsK8WOuf/
dmh7ZsD+Ldtg2Wz5PaeYqJYHxdTusN+2TfdOvQwmP2/VILjjLbI++VQjQsQNsuY5EYsZk1n7UFxk
vn808EUIHLFGIttT2xtULUYoDa1HzgdVO+SHzhuJGZrJP3rGxG3Z55n0TlSuKllHXLngXvNLS1iT
M1BANpmHaQ3VoWHvrMRxASpId5WCm486I+DVxYvqGeXNk+UWf7Z6wC4Slqcd/qn630m+/GBw2CIC
AO8xO1jmx/mv+BZhXNzNfftSxhLjy7vZ9ylTSYlR/H2AgUc63ZbxjuovMvFGYCnBkBNL0DTaf8Yh
e9R122WCU8ECuupQlkiQRu+kWgvp5E4DgZSYZ/oNXJLfZhCjsVHjiehIMnuo3WH6aAGmgSksFCMb
IA5bT1dY+EKTNx53OQYbFNqNhHgXQZ3VFlJuU1Vl6H2f6LWpZHgsQldpgAR+Yx/PRni2XUf3GHvS
C+7OlNo6TtFeK+HactCKB/Y0BonjR9z0BUNSonpbltKfWt9ZbfVFCRdcYbO2Y3jzvZKhv/Qm8OIn
aaOr5Cj2tviWKQPOF/nWI4TX1z6jgnkrZE5Zpb7MzsWjRgQESlJgY4RLIuPV+6K917ojyr0dudzn
ZVcEmUDGrt0X1qeoiClWhvswlWgvti3BMa2FGB5F635MHfB2JS/g8mWJeYSSgArafYa+1q/NaeR1
imH9VU6hWjcfRGmu1GPEVlIsobDLUHP9FrpwCAtUohW4FaAQKlY14SaZObBKin54pNl6jqlFGlQE
Ae1kXJftsa3czF43JmgWkHR1FJKfeBs5bR4YFbIyGfsb3cX4M5nuSZNGBymFz19/95mBMfSJR2Vg
k2EkUxvoMbkfDjlFwNWjEOvTI7t5EtlIlfDOopNlq9P3wF8cHH/b6sOVRM+kP1ggaJgHo42SwtOG
COZGLzaTYvo2imGsurRkqdCShV0VkYFSFC/iS57RpEoFf7H474iUEKkVUC+ZaObEpC4sBz6Zf5gh
iAwSRtWeHtN2blJaU9TBPOaF3sGPHdwKEjM8lSjJHUtYAZ83ST/qAUDsk+q5LKz5khVsm75jKv9w
P+6ncD3nko0r27Y1eEBPK3/crT5SWVGAnA8XgS0I/ZloQaQnJ8PKPIKWi3ViwmBSkPqPAL77obop
Egf/9OUF9O1QcNDFhCuQ1Z6omHfJkfoermkYJzAS3Layn9JFM02iWySpCwwQ2wd8ZCjPFb6qZrBD
XCUY+Sv7i1BIJ1u8zShdLai+x2SS1ozOfwuIJaDtuEIuZczJJnU7u3cfOO5cGJLQrD+lIQxRlUWS
eWiuHQANsoIyMTx7yi5wHDnlVhHL4rLyXNP5rj5iNgfGasObll6sauywq4wSgVbJ/O27vYElRCX2
7guQiMDpX5h6uGlFPL0h3I7dvZnONr3MMG+bKpVSK6gPd7QXJ+S1vr2IBJQSqHtgR2atweYxQrCX
mY5Yi3ZMUaP/0zJ62vMtl49rS7aJE7TkWLiRQ3vHDpOaO+DFufpt/0Zw1ktO53uE+7+vAwHet2dd
p6EkCSBAeggttSwc91ra7fDZ5BjGFzuO2crdt7yndOO3N0vh9gkcXiu9XTW4HL5S+oOwivH2Plas
1YgKt9vAiAZwo2VCljtDLUs+PBiGRDBBW4ORP7m6rhxNmpj5SSATXe1gbcYd4i9vapIjQxDuRRsb
LL/YzxSSuu0xVi6ymOwNcJCOV6pK7l0GRedQvepKqaYFkTujE8Ag1w5gMiXhZjlS1zNjV5dUpkOV
Ccd62hO0Bzz3ytTkiDO3tAAvrJoA1PKTNrlAfg3kO2rNMzOsMv87YWsGIOyC1wFhnP8vAvYnn7Pa
ttXqbVTQRuBI3WRZLd05hLodLfyLklW8CHKI2dM4Pb64q1aN1dBO7SVDPT0bkdlZbC82HcCuSSqH
UATFLjwHwZmePfTFrZatNLNFSqjSF5plOvzRDS8N92k8O0sYEQ7II30klW4fn2IYzsxvR6qJTR7J
OHnzM/x4hWSDrwaDu4Wlr63kBi6R6br+hAAQk5b1BZnjBrpnTnthcHHSh96rl7phw0JP8+ZWMRvJ
uTjXUCTPwPn42Tij2saps11jepdrxjoPzf4ENO9L0SJTzMMsWm6rEogL+oFIVUQzJobHVbisMQXM
Gj8QzGEGEZHCTr5UCb5W3mdHvYNEDWl8JSBfdSebs4FHjOIZnhxwzwXI4cEduY1z9+LXw7JK0/S4
2Pm868d5AsNKEDR9mpHXqep7Sq8CwhKUX/FtkRFciVlV3QsOjsmWvMjD2pJ4VstW3kotnLsdWWX3
fmlVYXpoqOr+aVgKHozcFMendeslT7Ka3Salsw9osrIs/1uB+4NClOZhXt0HRQAg2JLZmsGQbqrQ
YzhIFmLQQLTKKnKagYh1ohV4SXa/zgj0aKfSvmjRlUyJvFlq7JwwZIOpdOO1r8jOpQpona280bUB
uyYp2UYtEZBhFsG9XfMEOYDWxshStZtBbQ0R+keTGvsziTw4RCmcYj6ElPXmM3KgiINB+pCY0YPP
XCEXHsZD4J0lIaTWpENfoRFSqGzQAMfZ0PaX5yQnqpbieOWO7Tk2K0fdGnfkpJLVQeuxgBv4lOfc
8RCJ1W/Po/A/5TSu8ACIACzUbhOwex1U0sVYMcCT30h28xAPxmDEzxKYm+tFnqV/M3byHfVy7X2g
DRGJmTbXP1z7pGT1AFtqVBZhtcmerSZYetGDPSbReql8ZqDMDqoOaeVNv1eWnv9fGNFl40umB/1/
H5hcMw9ANoWGHsnuiAybaNkbYSwmaEmyfkeB62iJIXJnO103NqiS9hSS9dwWSWd3vF17rmdcMn1O
kxdwYuuPlgPUOzJ6f5tITHcuec5kK99ygDngDPtDeVxVbu0xmVbAUCqXndVnf9NjTAvaYbQ5/khn
3x40Bk7W5OUv9mxtmzrpnZ4b9dC8Se8WjjWpxVGYwFdMtYrzPEz09Uy2zu5F0KbBDR1qsXMAsRV5
qTs0QFET5IEoV7xL5h11N944rvohj2EoKVmaEwz5xjdWpeFP4tWkgmV2SKSYx0iA2lxGKaPp+dce
1sQwM+4hOeqncZHg1WAD0WuzJ0ViRLsP6lz/Qf4DSPpWkf0L8Q5dxj1TW7csCRVEghakEsYEHmzJ
O4ApMsOlM3EcaKG55iprpn4tD2nag7s/CEwgQBG7Gk2B6ZBoK9sI4iwfdNqMI2fcGolD/lRPskuP
lPPeNqMUBapqmGH2V/MUxUzT46G671uP0QfcVNFwFGckr+4Iz/VkcPlK3PhanzEcx4L3cCIQ9HKi
ff5Guyj2WpchkBj6LhOtGLBOPz8JUUOJMfKu6LRE3ymDMnx4+BeWlQPZb5dv54tfnjFfN2BQs5t4
bw9HejPrzSbRewmZMnQySgCyIpw9OE6BGP7s4jRxqRjVXRrEnmNh8H7/1oPoY/2V2Ia6Ejycxodg
eaXWAg/HuN2Tp2oJmTashmR5U8+NMvQCxQi3mCugJa+8uKZN30NGTlJxdm8b3Igo794MfkxQRdAQ
sMdUedH2EKGSOoWw/bd7qAK5qjN9v8+rgsWp+/ZfY4BxEOGt1sA8lX4/nwZWtdQFwnl49eNXukKC
kzUE982dqIh+GcDgQbqcJ8mIfO99M+PPz64pPJ4dVu/xsdcmlZpE2nJPeRH36ZQ8ec/4PJ/DZUks
6UMwvPugbg42sk4K+fupqehTOYGHSKYyzcEQrBFYQdjdBGPoZuq8YRCySajEyZ4Jfd6OZ+vV2IvJ
tu5B/SCYH7NRRHg5e32StNMUv1fAWA5R+Oy+4iL/mrusIc+xW2i2aZrUQIjTz9fV/DHw523PdKgY
bgo5+geC+W4P9wxm0RJH1r7uLw5dVJJrOmYXyMgOXG3yGMhningNHB1Mw1vOddBC+OqDgh9HrNBj
4QUNzxeJAdh6Rr1MksPofeXysjnGbWv1MlC+gcs8u5ZI1Mcgj/K26gqKBhk6RqdV2LpipVVYBJSW
K/+uGJdZLixQm0TnWB3o+FQpm653vKilW9Q40707b9PWSc8xu2Y/OKjKemRbdeqChzwakz/XPaLg
J6RhGfCnYd5d+ExSRtqVIHkiq+GHFmvLqOmCHgbiVGs/E93uhof2bGmcfJkHhMRcA5vSGqTmsre1
9dV1vxeewgMaep3eLz+4+SdbBXqy2dq0QkdwIoCrbMLpQ5udb73MGa+rmOXIlrIoWAlLGw73W8Kp
EDt20TMyBN/S2aBPslY6UiPnitWwg9JofB2248pBEZ68+uiW3gs6xEWTlWWIcx8258RXnzwtXs4q
h2+Gb1IQd1kJ3K9LwtDd51V/umbF1X1Qi00HA2UYxo1XwMUIn3UVmbhiRnokeP/0l95Urf94UJvW
I9dCwvIRR9VYyYXQztBB85zozKZxIdhUZpTcgv6ahoz27ksSLPMKQWuP4diquE7IcbdXs3JFBjI4
P0u07ZeYClFlOdP9lQWb88H83XW8hCQoclUjZsWED6dewtwYulH1MPLvD0DF8EVDCcks6Szbx5ap
yNFK8YOOGu0xu6mwPZFBMXO+MFqzYXykt3bSxfMznXvlA/yfpfWu9SmwYBGB7wjPNMNQNTnX8a9V
fGjJmI5Ane9kKOATqDtHx24fqB+d6smOcwZhn2b5DKEj804hE4LhJLbsTohohfC2oCDqixtjtW2R
ZJPVimfNszipz1/MJgLW9f1jvzMwYWF3RPeiKalSkJYPGak0DNkG3Gxn/FNBIq6f2bCJTN+H3fwL
QEeUQkOyZLcXqAbkLq5MlwxLJeihm082fcft19Oj4nS8I2siM2dI6wEYCPUcnZYc+6hOX0LmFBGO
eAokJqq3TiPge48Oo0neMkQzvzi6fOnzLom+zzgy/WFVsDO7yCWObQNbzaPoE+cdMJvHJvDhnduw
GB1qX0yKTuBHpAgqHtVB2HF4/5tXpnCJbLwaMT6DpZ1oNzzQtsou2SxcJTQDm4FrFHOChrt9z1wz
bEJ+Q3cDZIW9B5KOw9ZrzAqK2uNjjmPfqJo498q+5S0znxBmJCg418sP1QZDCOGcP+skZxS1tXEm
Qh/IpYm0qm+qarXkGfzIs7hqqZeMX99SB5A7zYEK3H0Ha3vvr/vYSaXKzxyj8tOd15URuJ9YmdaH
kdQBCgQ9R8KIwnDDMjqk4o1RJoJ5PahwgjxLYUT4yn6OIT/1B8Gc/UrsRo4miskgjhrWu0GS3l9t
OyepkWRjFBm5sozb7mXzAMOOLHncxMO6uhWQqFgZ9llOP1ilpwkdNINlAyrPJC8HOfY2BrrwLznj
yfcDQtrt24pFuZ6BlZrG5oLCvdI0s/c7XzqWPbjEIllVmSmos58NMWtXwfATBxMfxQRCcoAjUG8C
tqQ6Q0hCun9R/vr8uH3dgdYutZ/Vk5byeGTCDTMj1PFc0+8HbwZrmyWcK/EF8b7gDZ70nhPqC1G/
/m1RedvXvaLoUM2B72D7AYdAp7jvMo8ioiIBQtmW9744r6w6afGfK+qlXgiKBebI5V5UBJc+oEmr
qaw1qqUqQJpJuRr0slQ+dZFViNYAPVOkvPgTh8n3oR36SxhJH1VZScSei2zlLw1K3D+4BTLhVUlh
STmfABpnPou0jxp/fyNpGj21bU3rJSXU8Mo8TpstxyyGlYHsT+FaG26oGm7oFfeLX0WQTm7uEP4p
88JEXZcXe03d5lhg1LYGSJD4tQzsEni3NwsVTX0sgpXMDJaB5m6z3DbyUl+PZoNEl5Ftz+an5MXQ
Iv21IuXVNQtZO2sJp0Z6ehOXWv8Y+PryTQfMDdybYqUDm47+Tt4RDFpnDKLc8Km6OC+d7pXOjHPc
/5XmZh4ZwpUBwdVQPAdwsJO10KfpLhEdZLTIqz3WdE7Bq7YsHjuyXNKHBAY8eJo6OwqG6B0TA7za
zU/rhGUlPYU8BPACQrvUeOMYiXzsM8/7CEcv9lrgY6K1Fc/Gs0ZKECZCsQ+YiHzFgi8s79AoHsN6
xJ9XVkTHi1ULHgLrIsIU7Hukz0Zm780OxH6qiUy/Zx78GkjVOXBS5EOFIiMrjHEV21E7C2Lz3CH+
9UI0FX48Mf+WSnk5L3QQIgniIQ2SOgpv3Y+mm8RcTtJG7ciTRFsC4+STCCAn0s85qKYwybwkEco/
aaa2sKNuSwGeQC9Uc6Gsx6slEHKhtT/NvvoBRISf18X5oMdN8scQlYb6MuVGSoM2tyVFI3dwf3xm
Qow0soNfzkoqDtHjepIBa7uCwUWaP++mXrz4VZ81veUPIB87guchJelBy/8l5yBcli01D+b9Rpuu
OIQOU/XiXL/Fs0Jw2630s2+/Fuc9v31Nj0aJ2XB9rRHTWdNjtGwcmSCnTNX9zOnOwL5EC+TPB9Vc
HPSgNKWeTSYbWLaDC93sqhPAeLJj957XASQCWrTxwZLJvm3U6U9ycLL2GK0sg6/QOLEvaEVTs+V1
KgeBxgVQBMo1ysCTVVoB7KIusijbLA3EcLl3UhYHngRBOywMMVjx7NzNUE7DRjTd++0ofT7jGArR
cYiipWul3glt9ue6cYRBJRSPF/4wN1grtHE15CW0X2tKuAW//vRjd07LNQ+P58fDD1b3OZxczxLy
R8cwf0czKA2S7WJ2ZaLMfCIWuaCHsUS2Tu+NvWuu4CDwUZq15c8jkWJQEnnONGuYpcWQVf9SejcU
tNZj01fR9NsHgRGgb9YuFWm5ACWdOry6jt2OYWIKdnriZuF4zYsuRi95mrK2dlIGN3inJzTfGhS3
KC9iwBEHnCCtVHWlwIobDYPlo0An2u0GbliILVLO8TNkBFzkgjogHJ4abFzoYjNsNRzveg+0rd+m
1h8UOlE25w4AVGAio/+7zeedOaqS8JMZZzRvQAEZw1GstpUPVF1RthUNjxKG93/qLxO//tbH9sGJ
gLCBbYq914y2A/ehiQ1naM1BYO1ZDqzAd9GcplHwynv3RIgl2q5IVBWhl0S/I5eXUCD6CZVQ6fyb
+9n6u7YgVSMslAj7ThOIvdLgxFEM9e4ibD2Jck4yJPwt96Fich6/eNRhUJJ2+/PKomqNmLYT+HfV
HSB8VzHeFsgcpL63jExW/B6C0Aad9J8xHWV52KipUG4poliH7Gud6KHcqFIP0hEkyDBpo9mMdOTr
ZCc8AM66r68n2ykGnp3RsyeaoHS4b5QsWQ96IHuOvWI0ZidV6uy/KFIT8BhO2S7Mrp4kYo4BFIgl
MjV9q4+A13ShznwcmQGiYVDamOgD0zZFVEDMICAaLn7o6f+/ORTvM+D8M1w3m/pvbyklZudF2ndj
5Wmda4pq0RzmrwEQZxDqKLL5xQn9N4Ed/RZlycKodYMfbLyqP+kO3ogolIHKv8S3et75et3nNbjF
p2lTVr3Qj8KHPK4gmoYAa5w98UGJzuIaRWXwHoit74uxAqM+NwoMJFJ1eEcd0+IbzcAwRtTciXIj
WuIogICpRBV7mQ4vd7PctjnJ38foZHePhlaNx6skjQNFMW4ogU+N7ElgJ04/FUwcgMbCNycUFI8k
mQa3QhhdYhZcIkf9uW3nB0iQ8Rc0h4e98n5AtKjp/1Pv6hYVuciH7kq7UNki7hJEM6Yzv13ud7O/
qJUztLASIPIzRlzJxgh3wK52ZOUDgQ2r676+atRnyb5cQnS4FriA+aHhRVure1xStBLdqepWktcL
xOl5E98ig/CtWqbvsSVKcon33wbr/DPmeQaM+d3IsEWICGgR7xLClJONbUM1mrmMO0SeucP+jheb
S1sTKzkW7UNX3VtzFV6x5Ar+Zt3ojR5W7NNez/ONflQmrjdi/EsN/eRC3Dr3SMlm9Yeme16pw88q
y0I0xOHI3QbCN4CIII+v+dLJx1XLPyDkBkf9P8Jmy+paVrC0bQscDxJSOgap2m4jjFpw/Jn72KU/
fagL26sbHnKTH+RdC/fB8dOnviKFJyQI+0sagxKX8cJtz/hlKOA9nhrRenUoin7+m+kqgjPO5HEC
QA1iIzfCBPfj1eLihTBCn7N6UXbxerrciEtSB81z2Jx7CxtBwuRmR59pTM6DSJP2QSld1dKckFuc
W/O0cMkEV5O70uBTuquGT1aenXPAppyQryT1ZQdJfQQ2Sk5j9uINyh0loDUMDCGDZCDohUR/i7RK
X6Tdf8Pyo0VCA/DdaogUrBmZ3EWwcwOWIN/z37uu0pJ619x0wIDPlukypSnxmHRfsyOWOsh+0deD
aW8WNUj3SD8HomCjVEfaPZDaK23qDwAst1kaGTYAmKQoXRHvH2rVr3ThkYdxzFiCF2BVXDa9XW48
XRCel525JAdAzDS99k6xAOyxGPWgm4536mQb4i2pEanUGgjghCJUwWHegd9/r1d5Ttd8gOvcGdEy
V/9+mhPcL14Y4pV+3E9WX4cRRSBb61EZMM3up/SWiwaGgvvvJDI5aEyvq+MSuP5tEbCkp7GBWUR/
bhfAjzawlw3wTLULqMGGwy36Xs8LPBCgzD/Oun1aBwJWMla7EnWpGBKrfns5HyuUV28v0ZBW2RNa
m0uooXIjaSmzGSEFt3ww92V2S9OVTc9N36WJr09y8lRu1kTbpPwVpEqbBPRBlaWz4tcXgqTF2Smh
wL2xY0R+F4TPfashs4vCqT7FoVBXcelGtpTjmU5kZJmBs2VF2ZcpP+n3jSsjt3wNNx0Q86moyhLE
fa0/Gvw+zRzaSAWlXg7lMou/dBHEtGpL3M7AeXTB6SGWfZi0+0w+ID+fcP9MxZcMpFolUcgBmMgq
EuZoOJvMrKL+Ni1ToiFk7cSeNwYLvUkFKOHRhic7BXIqeCtzfm+Hqc4DYkFEaYyII06ksHPMVgyF
KMXwBlTsV94GD3LO8S5IXJ2mKy0rCS6Ed4cOVZtPeEqYWhShSjCiJwp14hVEym36z5ySwr/e4Hw1
cCcefmwmQPbb7rAHTQ5hnjyvNiJfOyJhhtzrz4MNeM/0b1//vcP0yHQnIGDh7RZH7abHizk6o/E9
yrFzlnC83YW1zk5amx6Pi+8/dLgTARS649/TLHSXj2QpX3iv5kSThNaUWGU6OaFXgJ7y0EHles9k
+JHchdL03butNHXY1Q6ukfR4Vb4P9nnCGM61feDC/uYCyDQPGM6TsiYh5OaN2ZYiZdviHJ7yhz6S
qYD6N1m13RQTVUSJaYow4lwail4fSrRe5OPMFEhwJxaByxkSrl9r45k/kV2/kAE1hyEMqCMxnYx0
3OBJOWqiBDRbkncehfjO53b0JXDI+WOwa4d0IF/8Mfr4tiRmc2gg2mVIc65Nos1KbCWm0LpRlfWg
XcV+6ZLSh+E7b0bm/7Pt2hf8GzaLPUS3Rh92MEY2Q+MCOJf8CYLri+hrhJaXbM8jOoYNLorfDMsq
p3/UwhPHKXhfRKTbbPldvTyohn4jKf9t1jjoPePRg0PX1as0pyMT6TpaDOO1FdGVS2cDORI0rfUT
sFYsHvJuadGkkGKP+VnVDnTdNyYyGXDjcYIJqDGeLk/oWzDC8j+Vpc5ImqWHwmvTcLuQ7xfTZZ0+
Y8h9cQ/x7KX5sKY/PAZaDOVuOcjFY0pOIqbR8w4fd1rGJ3UAow86+cV3s2sKO8SYjyIZ9uE7z6eO
3nvNp3NfxdE6Re0PR/6yC6PA9cABY7g16cyr1VwlmcNxgWseJ1dj7ueLSRUHyECTCYluINBPhMQZ
AGMBzSRwqm5MuUTCZi9cjrS9EiF/8RJJ/bhVUqGr5ZhMxcxO/RfT65FJtIoQXue/ZYI7BxRsUI7Q
gO7YHdMUMtEo4T367f1AhZzO361P/709HD3CjNt7bLA1XwyvZZ09IRYZj/2DyUPTvyr4KMKX85KP
AH7IM0Oqk8m0L/R8vm0EYLuMyzSzEzCn9U86guJkrYdx8e6q1R90nBtODXocIJhWuO2NaetJbQ6n
yvjbGsWIEOWl6tBP6cirYt7Szhk6jTCnLgZetGHWx57GAyCvCZrYab+o5fRB8BV+IDNh7jtTXURS
93o6sA7y9zPxIUga/HiKD+oaxuqICv4yora6l/7EnaLxaU5DFpLo8KM8r0/lVCNvgAYLpTZhB2Rc
7Mbemmeb4kbbPpfwS3pcNWtq39L9/oW27W6irVFEd9PWyt6DPQdGk3uvvIvcw2s3npW5xP09BJIG
I9hA8jSvKJqan2z0NzKv0C9QdTWhS2aBFRASJFf8pmStjiuqaKhBHJ69LQal10ULqjCRHwsApeUP
vpw04g/kEWfT2gRctnvKqGjQHofNWhMeRyIKV1neOypt3DD2uyuCk3H3w4V03hnVi367F8riLmBa
QvTZ9NxlGb6ALb+lfzqU8mG/kD2R+Lgntaz+XEAr+erkNmTyNeDS8h8YmbgRtj66w/bOM9T0lOjq
0s66bu4sqAlMSXn372SQtPZahSmHzk4mu66HiKj0O3dRuYXP/nAFc2cNb61cJ9Dm3XbvjmRS1SM7
2yqKSh/RAaToIpeSewLSD/c4hamX+OytpcrJTGF8mkq4P0Kwvv5PIMhyxw1SViqp1M9NhNwix+fR
cinEhAZy0YD8taHaekSjJNrV2yAwGzV2QLEcRW57fS6X2Y01eL0xdRBTJSwWgSfR3EE18ji46tgk
2en1aoR0rqnGmRG9I/Pj8+fFqSNhpYOhIOM3kFaaBIp/T/WgUCBdgpDu6nxjI4KEnV/1Ch5Fhb6H
CwDScvk+oEMA25qLGxQNncMwpup4zUovREQiIU87rwBGY3VbsUr60EkCFlrQt6KNLsdTPNRwStyB
xJmdtBwlpiaXPp4QbI/Re9VROIQj8o7+yT41j84aULJ0U5XSa16X2YyXlARYSoHgZu4FjC2gL+yF
7lFv0IDoJQlXs3s/hUWKmsQ6QTVWWOIJD7Uh/TMKGVmAew90z9zoCBitWQJ/TVZG/MmRo/+0PJkD
ABVuuK8Tx1PQKwvsyQr9igWoLuy33QpiHM/lHSPJWFlY9LzgKxCmxZVpy+XJT3gpipqqo2NlUdtC
LPKoXvUM8Y+S50azCFshVkja9nxG5mJT9YOxhTDmJFQiUtbAj3s/WEAbQIPF1C4FmsVogfEA5b6E
y6hw1cuSZt8rkpu8Ef7v0pCR//Tsa3NtVmDGuIgfv+NgBdi35AfmSdxV0t315LbBtmsHAeah7FNi
YPeXPuD2TV5g43CnrEA3goiujGhmJb46vB5LUwFRAa7snwLdYh1XYMN6GTSHpR3f4Tt2FOfgeLd8
/TkG0K/A6oNlocZU3mTL3ezWTJPiJqOTbjC3cRhYAze5DFUuVDYsrLEjG7skQCJG810j8ImuhUGy
+r7RFtSPhvMLVhziIZz7tQehiNaSaPKpCcKZN2TBxGeAuw8JYRJFMexMfIuwLDBLpZTAYo2vXkbQ
igvjkejAerwDUhQglArR++YJiF8J5Lh2fkMz+erfWAiji9692K6+Rek6wfN5U2YFE7AiJj8M2Qnx
kmZBUIC7zBtvf2TDBeTtUTJ+25YBCukRRu5ZkEje0o/sWbWyaShPltHmPrG1DXQXsvv00pmLbEea
/MKqyFevzBtH9QIiW3K1JgG1kyz2Zl9D0+y2DU7DaoGfVjlQiKfwaYIgpXS0msJT7fwi4IaFof6l
PkITKKO8t9XQLh3skOuvz6fdoRLjGGvpF6/ndDWkF+eLcjY0GC5RDOx3AlNsAyklQmRDuND9Y4Ia
wlVGef/PLwF/1xr+DQ9ezAusszcDy0e91K9LqBnHpc42GnBPLT3+qFf5YaDlQAt4vE9Ipi9PSif+
8DDfjKQS3ZWu7x5S0FF5q81lXajndH/Bj5eyCeX8QGSrxRIdVVRuOUUxRLJhHbVDa2E3FTjjpxbg
nTBayZY41pBVwQGQaaTXzcVDUPq/yAsywQRMmM+FG3bM3/Nf28tZ2KZ8ZCbqVaVnoapwhSd47kFb
d6vgIjMQ0CbSZGqL0RClqOsFU5nIfWPvAQV2PIhSydyu+7hYBovVKmWxoxIbuRgtvCE9vpmvXT04
U9bCxf9PZ+FqPNJWwF7xXvmawdOHXEP6Hio0LbcOunI8CEWeFzlBEolzBZ7ShzSxnYFVWckIhPr9
genkLhpkfAOdJxXG11WTFCZLM7qKlYomy4O8aV5jOaHdqsLoreu4UNo2KOBzIyAF083bbzMm7fMD
vSvqbmXLB1MlJ7lhhdDb2NESYY0LY+qQjWH2jsu8FeEW7wVV+Pa5kFKajXX1y9+Jp+VZ/SUST6Ud
sgDXNkUKC4OtpIUWQYjMwUSi03HtzpYz8MYZ9ewJKgTAdxZ0Ubfsi40CFcwMzq1t1JOBrixf8gDS
LnzATqWsP7Ui5VG2BnQYCFpPnFV4HUT19qLkxLT9UURM0aoS8OzvITN5eXhk9fYvW7TgUw1gDPu5
HvbWRXzKNnNVQzpifuhFAhh4RSDZp7e+QfR4BKG1ujM3fjJrKbAtgd1H5jDddZvTOBrSg1Hz9Hkr
2ESRlZm1q10V+vVgUMKCrB4qFrh364A0lLAsWWv7GSrxQa+zqgU0E7e8hvLOkowbJvsa5sa4+PD9
dkN++QRvBc1xZay/Nw9zfDTbLlVs7sAVRxdIg/8mg2XX4Cns3vXE8JOdT2Z7o8cQr2LPGfKM6MjI
TCYkz8GGrbDX4zeBr+LGBapLJcwF0qnED4p30w1t5vRdJAPv/t8NnVa86jPKnchRW1O0pdYRfD+N
Ww5vqBPtdpKzh7jAhX4qkGBcXmbS8lGCDy+z01wF40QghAtrm575vI2XsKDTFc7Sfo/00guo84ez
Q7ZNaKY5kxWm/sWktOECAxB3jmA2uPPxzZbZCZtR2xAjVB14fG3oVMunirNU6SFFlS0NFQjorEZH
zZ1oQfu3vnLWXzgszCMdHsCwKDl+FkhwszIs8ft+dI2Y96SwN9tivBgLB0+l//CozBL3xmLt3cGZ
x/q6LMl2MQunqsChCuMpziZo1eYG1ihlsUedBAhQFCOyoN5qQ+EK5cH+JVz1IjZBcZgTvkaj4le0
+fYamNHmuJw+s8Tt19E5EuKkF9JP7XtD/HvKRw+n/RQVRyzn1F03+aB2LOE7JGUScqCNzi4Gldrv
BS/J1kkEx64IgrPgbZiLFLIi0GdQ9FEvrlP0kFp1kXSdV4WMvg6zIbsjLEgpPcucviCVIgwTry4t
m3d6EzUwsTOAoKTvtiY5FMWXawSmG4b7PumIg+uMmwT4Fd2gzxZ6Y/33WHyyNnSqz1LsKEdM0voF
PPKbuVqimVfbAT/x13dcdgugG1FG/9HKkn4JWZ50CrY1U81JHOBfu92y7JnlVE/tSp725xU3k8UN
bokv0Pr9MVg8U/f+7g+0NoyiqnbHYPH7Hx0wM0MjfLR2ocuEuPGlGMcYDehjWs65K0xMPNLCd1tt
LKVskDStYbbznEeGrLJ9U5wvDKIdNqbeN+gGPBwDw/7887kvYKDPk/j7Yeg7yAyhb/+AJvTD+NYz
w8II7l5dxXgXtl8XtJ7nPiqx0qzqn52AWyrWLlcQdsiy/HjHcHhaC/093pJby/VQ5CeyFWvN7SMH
Sj3oD8XDroQxueafyDCdsekDCBZGHJcV3CtXqtp8ugvK+pRMi3Rz1M95fw2y76ufB0a8Cdk1+/0s
lAQhpkKVr4p+8g+jvIJzu7MnqEo5imZ2X1SM0zhw1pn5RhhNhjI+o9rQdha2WCBNFW+kABePRrRz
s2FMuwocOCx250h4tXHjlampVQtevntbAn4dwHT2PUnlxcABobwFHSJ2CwvfYuh13cuUg7mBGisz
uigw1nG/3Ok9AMvK/YbOWMlooH6VbMwsDEOO8cAjyGRBTz4MtRmvF3/b0pQvdCeab8H4cRZ97iNf
b7/E7mCMnvC9RPelFfW49Qd5GpbJIlD9MnhtHd++j0pT8mJ9N4yDDg1Gd4mvwi3rjFQpRepeb5R+
NcRJOPvzfK6z8iwNEiO3ESigQURcbrwxiGaYSoN8zBBgIUO3KHqenJjR2alpt6x63WlZ8kyqvrHs
NqcYAE3/BRqCbY/kZsNGRAqSjKkMDFtbFhwa+VxO1GAz8yOVp0+TyKIh88cqG4AVxaA6eMl/zbz6
dXWDZ8ABeTLrca9NG5ktdMjUAuV932jYJ+yQPJbFhDXVpZiqPnWBIGYJn7AjLTrcOL8BQDgEQaPl
c5KFXLsKNgiTuBWpqUi8OhYfEOXWmA9pwMFoQCWBs4nOUd+m1CGU+w8RdYR6jD6GtkmGiAahA1pg
IDP8s1Ecw3/xD7MIKeWLgpm8oZdvDgFz7wtQD2t8FdLNvuxZAA8+va9qxh0xcxgfVw9Bj7xQHtA5
1ySqKxVLTnjlhw1QkYRsaeeDRU3segXJJAMQ16SAegSLL/3+Wrm6tV0doVlSoz9Nub4KrH3zIrFS
3OrYpSoGuau6c/SNNYG7zQR93ZYHduYBBsTB4PdBT2nl/InhdykeGbmBwfhGmXWSz+1PSSw/DsXs
39lcLgijvbuojtWKeaTSqTnZpIITkElFJjuVmemX6+YrdFYK1M48YERGUuS2gnUJdjFjFG5tdLgU
bGNVdbNfbCjrvdsuwqgBzEFZ0Ht6JcnuUSbMbyKc+IFN2d2vm1NBdtB2pzruOe3xZp4fgGNGP+Hp
5/JV6nXVYuX2HJFp0ed+EaFklffdiRSJY+6E1LNWYsQ8MErOtaicj67KhB0FBmkABxOsHLq9/RHm
QZ0Si6+ah/1SFJ2lp1p4ZogyotXM2MSOXVW+Md29kP2/vDXVSQPPChnNa0HSmsnnoPVHk01/beVB
FRw2THnC313XxoRSoJ3/sA7ZjzeAY2Luq3QZaty89tnaBtQwk5/W1wsolzTp9j55ZcydyEuJmmdi
TPTFm/eNlOGwjV5wEPje/MAYxPbKkSe7tbMhAbGxvUgJlrpPJE2EVoz4ffRHcwtdLQVXw9RMdrl9
/Df79JOy4D/lJ/y+wz2G9BeqSj37Yzb/3k4SvFec/N/ATxgAHM+CmKnit3Ty2IeVCAHkuG9ZL5qM
omAMPRedgzu05C0hm1YVrRnuHfYe7DVEUWCRbHnZ24h9TwjeGnXXn1HEi8U1h9ZM8hfzwrHv+DZB
WekQWdA6HQx9DtjTwNGjNidKxWE4A7EBU6qVTfNXZGql3F4fDOkw5e5zUdhMlUEdm0Xd9XoG2Ei3
bqpFb/8pEgdSaQuGJcSv+EYRKXy0B95Dgdvs7gKUSlwH0Lne76JtBemmuNX0JeYKBUFPDPnt/lQ/
BvEWvde53PFNgZRnshAtrU66KOpd6RPpbFLj81HEBd9RcZkjEJXyu2fEtQ1ZI34B8JN/eS/OwN0M
bYFQnOc+WgilR5xXadWkCHvpl3qkmgCpkr+TFTAnXNpCEOuBfmStrFyGIkItitDnuWSxSQNAU3oB
48rk6wbW5L0bdpT6spap/o0nHmTEUd+/YFhwTXP0PYFOzlOBQa5O6pXjzg3gD2ISqeC3JpgoRUuu
2ERI+/QCBoASTVSCoZPpyEsfElQMOvwn4OhgYq81w86ZWZkBNSVWF6mq3ntOCb3Rahf5OsHxYh6/
ak1enawkwJ4Nq7IxSzmb+TgW5ZRJb6cA124vxBzlwQb00OuQJ/m1ZmhDHcFx+GpGmwqv55V62aPC
csebuzzYmlvdzBJyFC9OyRQ+2Yf/yFzcFOZB1Amou8BWUDhl0j/ecEKqHo16sl2OK6Ef5Fvu7UMJ
mY66tJvGZRJbRlNDKTFmPYYsQsk2K07+lM/HkOhYGdpcckeYrHbxOOPXOHr5UPDcorY2x3sO7+Nb
qx8lFf2L+BJGELAf3cY+S1yloeIvQzftC1ob6z8wm+dOIbf0g/TJFxtuZ3jUX28APV/UxTwlwZsO
iRsSx62DGYYPyUs2LXN/2Ub6bhae7kH0AX6zxV9fBVrpRVF/pDjL9g9g0rK0SAhB0ScFCQ+vqgBU
2BaG7QdT3C4nNidWYQW9MFxbyP/3aiGaLJ+H6Z4UNyrjaLuzsXdT/Rsbx3vvH5Y9ExYWTmyoqelI
A2gxevDyXm/L0Xevg2BFlc/BCUVjaWinr4CG5tnmRs9tfTC5iAMMR9eOUelRx/fSvauoKOmuqRsT
8aYsgF/8klOGldU+/7UXR16DEkXTpkNb3NHjfx8CccbtL5iYUBjdnw9NcMdZ2njJqQ31S/3r7hU0
/BqcvegtYPGUnEugjQcNATMv1j7odkjUBOB/lDBdFkv3jPPTSnQbSpLTKnYgm8VP9Csp5Z0SsHuw
W3MrG0c8AO6362HvEPeG2QwLTfQQ3SRsgu5k8NBcyKzTRTU1Mob4CFdNJKNg+2vLyDjiEv09OKU+
iEZeBmz3b3Cld5U120vVfreDzqR3yLIOjci0aTvn+5nKcHMOrqLCJhUquCCPH9Qyvo5UcMKd5wg7
cwGUzw/DK6o5DX5VLi3y8vM3pHWrqLAvUpJdqzXM+D9ix8iYcgpReBtRpAUX2+wLGROtjP1x+PWF
4AyaHg4cNfyFQA0fis3LSI4m4Pu1OoP9Am2BzfaEqcu2ntCjRlqi0HgxBKuvcI+40EhpVYnJpx66
dYmGPkjOzpSdJUgzHssV8yM+jpBYYtpPnTMZxhC/bGhf2L7X4DLX5mjVbXCdMx/jU1c8rL96ynOJ
IM+rxUTkFVO7WBmcgkatQkXDrT6ColQo6wTxrSANLCyws8bv38Mc9jj5atr0ckSmIEtx9Fh9CGkC
RVtgMJgICI/WdWHlQI+IP9XMk04jaePlKIL5eAV3byzysyO9//uWiGpWIH9Z4364AI0VnXHsQ/b2
Lr1tsmnjDyZppEg+BluF/23u32N117qt8ZX43zWgk823pOe0G2q9fHtF6Zs1a2a+TejPymBxjxyB
Xvqm5J5Zb0k6B1A7bcipValdRlPsmrutUrx7Y8jxk4gW8YntxaZoMI45F9sGRtgvDOiN825EJone
SZF5DN1FXgZG7Xs9z+wpfXm7UftKTyGjjGJzNj0q178tgig6Di+bRYSQTS7Nfu+C6AyR1GqFqhr+
QrWUcjvRwVAEgWBmLTi7S1KhTFt/bz6SSIlw0JohG8E8WJd1JTTtJPcTZTSNDsvb+wlpylBDrMl5
xroqoFXNvhhTUiz1I9+XIagoMfZ1xhgCD0loF8gTNwSwIGdMN8COFXkM/bAiUjxN9fncE6nsRgUn
+E+EOQeqEr46RWLaxwqvtNI9OVo7wo8VknbhqQkQ1Ps5S9hwQYmjmQRfYjA0JiYckcenqPgJ4AG9
trXVyYDxkHdXGR7cfKhTVpUGFcUAkq10MW42fwlfvvqtD15efzztrcyWYbQro4J3yRsj21agEb0t
KJV0OfFooBgN+Qa7sn6WdrqeFBP+1S4FAB9ygX/8D78d3lfkLJdZbAvDAVEz03dqkb24O+5OmXGs
HrUxEYT0aynxzKi5dYukBUtWFAtAZJyCfQkYnoQtgpQoFgLCAoS0uVNzPe04bTCkHLkanWCTp8SR
hry/knCyQIrJFGh46V3Vr+DHyIbeihNsHfSKHq3veSYxwoXDP7FvVrloq2kMLcYM4CdkNLZ7PmcG
NSatsG2gBwM5vnNclePumruocD988/+yPSu2HRQt46jwKhqBc8+3g+PgSY0RUi+cEFzLUn8J54zU
pR7R0oaYo3cVnCbRi7H4fZd/QVXsnz2FmXgopCP9Qx/jGo0pTXc5CAJ4kY6+d0dGFv9ViIgTuxl5
h8aeE9H1wv7sfjWjVI5CX1jhFnDK+tktCcirbkLQ7E9ZOklKEFCN+MBROCRplScvovzLBhKgHGAk
MmlXb912642CP7OZQ/sKvNgSV+7KU7T8NCQkcKbe4w0AcaLcztPQJm2HRAv1VU5LDNJKj5x1BxEg
y1eXDUJbDVw0T2r2RF4m/rJH9JS/OvpzqVwR20b/BbEcytE0/0mlel3TuMZc79tYRgzLY3hOM5oL
c9Tud5/YMr6yD8u8SmVQLctk2Oq5iJp8RJcufuFXKIvL4RqtMSorOLCBqUuLuSN+8lPyhnXvYSUC
tkpkZyOxFpG6Q/qq6BjabmlVf3SBAA7GYKNXG+lDXz4X/CS4pe+2VGfMk5vNF09CsrzcwP+6fjd/
7c1w9O5DczjKJrmz8Oux21Y/2WHWLZB67X16F5XSjPhVTRBzX5zyEFyQcQmYRlTDe53SO/lV+6mA
ldA98O8zQURk/jf377RS0rEoqCRnRIqWIUFosEQukIYqsPuypwUoDyAIGNSjDBQKw2meOnhw8G9y
m4x5zCEIHY41kqYYxJMtz04U8bnblcH/a0mQ/d7geKCYC7ie5tGRYnxXoRkycSBkMAyIUd/hBRc9
rjSmp2cxf7fVv+MCrFV1Mc6BcHeYeGeUeygZlznS/9MBpYkr0S9SA7eo5A5yHDJMzbPW3BqTcSJn
Sd2LE8PqaqYSm8goPYIBBHPwYRJkMVcUp5H+wJLKCCC4ZP9ylh9m7lC0IT9u3rxxmT1UTPEesopW
W5D63H9r+SLMAnE3L3XAnoswwuUj+EPxwjzt+ShFSHWSzfgPHdvjZDJmEpo6imaDY8qaIdjpME6j
kv7MRXC1u0qkHTtHLlZAuGCrkFBp/1Q9PzR8XavmOHqrNsMerOb7xMtrrXQJXqIzltSDxfizakBo
/CMYwkZ1/Jf6tUd9uP2hbaEUnynd8SOb8xd8wBh02K8g4VsmqQdLAnS+LbR8syGz1rVk54RqMpOe
v/zhlwA7YzeShvhOgflCCXQSXrN6gU9ITfLAx+VZxwpB7i4F7+1RjekWPB9Y1Y5mTpAJ1HOe2IzZ
vgmQvSLg99iXWPWcjuRGPHyJZhjdVE9YocOxJTdRHK86cSXS6FI7EoAoTlfONoCKlO1FJninMkZg
IF1qlCJTKh3hcmoHE+fAKMQxGtz+0n5rG/3A9ZGx0HQkLllpueii2XLF7yauWpEILXDYZfZkN+uA
7xHAn87kkqENgEdZmnLvcjWdwp1UY4RnXP125pttWDgXFcNmuIwf0iIa24BdYUijVMFnTSSX0JDt
T3J8Kc5WBNwzj25Ylx5xyfMDQKPAdlFJwBGWEyRXiJXluZoPxHyPogDhgazSuXEpx3fCJDN00FB7
9hjSipSE3HXWgG5LwOgbR0zJDZB4UCWA9J/w3bXKPE9iVWAAQmHbxCg2IGcDxQFcNu6Q8QkWi7x7
xIoQL8U5HZVmyW6V2X0bH5mMV7UQ2jfD9igYiyZLA/IT9NHwLP/zwRa1XaHPo7ULa68KTAeVfuHh
SoplfeQ2lM+RfitIuW6d+Y43mYQ07DYMGKvyUB4TwK1W93692Eb5p6ZQdsIWVxlzZsYjfhCLJA4S
STrgZ98D4RNRwcyB03GlSqSdeAIaYPQHnohS1/hvHNpLBpM5p9ivvBfDuVPNPFrn4MXOGjJS/EEz
rVBsPWmN013BVMbcoi9F3AQaObP53iFsfftxpOVbUUcCVXQ0p2hiLgnptzDm8bdO1A6xeEJbNMRY
abjeIlR8i8quOoUqAa59dlkt1BrBq2eCpUB6Tn+kvp+U4rK/SnP3OAu88DfttnLjugFdlOIoWjB1
VZg/yL24H+3cbFX9Zm6ESiMHtU4KU8z0NSmnf7FgV+Ml84xGTx7I7Wr64QYjNAEeF0suTeRaZ3lc
VxGLZ+N84r50ZUbmkUGIcXDs+hrBu5bLxvJkOwetWeIwj55DjOoihIPXp1cON8Y5IxbxwhElPGsQ
M0xLIk06Nm3mrjTRbvzGbCHej0FsMf2F7i472ui8xtHJqg2jNihNPVukN9TZsriUJdyTVztDGw1/
vwBeYyvnc8tIf5Yct+Hq5RE13E5Z0HeqxEmQa98P9dMVubrUJtzHVOcQRZ+705HDRswLwYO/6w16
7HOYOrhgvmvDn/Spc0+i/e7FMdyVWau1TGGBoHpzzQrEEGp4kCG9yApKYYXdOzhFtFr3MDUbQ1c2
1YgjYjO4XeR3FRC17ier95Kl+zlSWSSD0XHBhlwIxuxceSjlkqypEtCJXRt5VA4vLKjw2T9j3DIc
+SC+Vi/O83O/CX6dB0LXjQulLqdm8FZMQlooBG/aqBqn3aaAPBwaMRrrFpgKJx9WE6oviFw2stNB
lwwtK3DhfZHwO2cDZeX2z8fkvmod+5ydHAXHvdTT+OKHXsL/SSVQ8IyIv3N4jeom8s788Nx7lg5h
+FgnFhCom4TVaPDB5P3MhoA7gdEYlIrBj+vsrYa6Sl6appltGPlJLf8rD/8UmslPsHlkfDTNalfQ
8jN92X6zRXp+dpan2x19SbpCVGvLLesm6TaJkxF16kUEClNMo6O+N1I4cTyTZlqqf90dDKenDyLl
9fNvf+KpGm7Pzpems/rmOcj+vYfVQULXnzKktSo/Gaw5dqaCWPGAmU6kIEwzYcbotzir7BgGOyoG
SdC5Iz/eNN+GrJs9FHMwXBejFOLuFH2hClosw7rv5Tnpj6HOnrX9yw9otOxxC2C2nBZ146DNYVg7
IJv6KzBLUIEyNcuD73u0y5u8b/przdYTBmH8kPDHxPVKDZ6BjQ38sqW8JXXSKGHvbuXUiBtICSD9
tBlteIRjE4+Pqazlj9Sx3McUxz3xHpHspbRVT0ijKa4uWdNMzHWH9tWteMITxQH3kblinjvcxAbX
23B2N8KaRGglM7t8OMl3dRjTb6Q28tm1LHcevAEQjmGbhZ5nS6PIJrMPCIpOszvBUMx6IZTTxTVY
fPI8HFGaZs+2W/Qwp94VTVLDvNBm2myfZ7jztjdY8BhvqBzTS4nwWmMMaMW6DYY7bhrLd89v12bO
isddeQKu3CPk2R5Gs5QO6dboDsYb58lJuWGYj0e41Xz3E7ShjGiuenMvk/la8lfDsJFEtRuzGi1D
e+jn4qvP93BuFqrykNqVcTCLBTg+rm1PXGq2rTuHxXQY0q9qOOgcXqTk+L+qp8VDAsiYxbCdOsCd
eRTm1UedxA8u33fOXjVfV3kezwoBRdNSidHMSaDWAJN/4kyCaB+b02Jv3cgCnLtcRDvGwHHEp2rN
//LJG9JdUjw/0S/MpQIu563i6sAlFnIwyRkXRvzDPc4Y1mIUanAjPcKt8ICcT/jkwzTD/3BENPBk
GXFxyPBzsbGhuH0ZTPHrejnndPMCRz6tBsHks6Ytbm01HrhUnoe6nPdI7wD5gG3AtRe7p9w4g4Ye
w0sLyaBai/KUNT80IiVWaTTXH3k4l177CTObJIPpKFP6Y5gHSdlozmX6QTSGMPIgLHKPGS2eiTQd
s9ew/rOdQRgtSpZ89UtpVL2UFXj7jZvp3IImz7x5yPj3Y5ethvRZ/aff6ldFZb6kvM11PXqfRkNx
m9hLvF44IasN2qRVx2bZKUL/CBrRlhyzEtGWdYIx9v2bnbCVz/dzXl5SRobjOYQcqeFFDrI9S0n8
EQoENaWNU2zBxH1XZ+s4l3Z5HDX4D1iDwlcngziz/TJJVc1nrhKFajWVUQKs2GRa8OwAVqXlKg0H
kIHShnsok14ZeNnjWWJVd0LXiRb0gAbd9LSkObB1TdWR7RDPNg59HL1WeXKvu3425C+8083eJvUs
xXbCtU0n38sp0CkXFfmLtanoiPgG0mg7PdYInbgRxxgMmosn7NF0ZPm0vcqmv2pO9GJpvLqNYpYz
A6VE5zWpqHsLmQ7ItK3yxhYr/ymqgatGMT9pN3fvXJ+AXzTemdvfSGx1Q/+zHb8QRzaCmDfRDp7N
K62UWiobDo/Gi/ooacSMDzTVc7R9wDpE3DidUaeJdOi0vSW9l5BS6OtcaDKGV/T/huFtiHNx9niY
rP8Lvke0QOWERtgsF3xs848FLzU7fzuHIioigS5qE4EKtw0+SI3HlpSZRU9L8dSofY8Sg++Vag0s
Eb2W7X8fDT5ME2aDW4SbAzuxNLe0ZELHiGR6fJZAyG8EQazxxbU/n7+otarsdjwc4QD8mjBkBU1w
Lpq+1HVyZ8lIBEGHeblg2rznvH2yaSBllxR/l9V54AalOocveqdjx9ZQ/qxyxnkyEH2fT/xxc5cq
YMyCc3jQ/D5GoiMWPrN8khw3Ok2x2sJxY3ajwERG1qcLM4XpFsMWPFY4nIHO6vZjGEyW9nH+DlwT
JIMmiLa4m7MzntlwoTl00UuQVMO5CQ1453Cqh7m2UqZNZJiptqurP6RLGQ28Ky9eaLlxJYbAkHsh
X8DIoIL3ZUMgSsgY3oEj3ZWXHf8Mj4T6t/hFwoVzrPzTDaCugCNfQb1HCdwdszZxG1ZSypC+b5Yu
c5x1l+fhhxZvxLx6dkofCv9kuzM7Ya9PbPM6BpwfNt+bUT6WizcPwPuswT1s+fj2zqz/o0KHtcWm
dA8Mm1Uc+kLfHORiVBViNbfloe/JBJhMMr5uOHRAI52Aq2wKw3IC1aHhZSL45NMFCmk+xP0BS/+Z
pJmmfrYFSWZXuddAOaW4e8q0kC9ofanidhXfdu+MTo2ul3dBeU/Gdg2Pcf2pLeoMi8fYd9aWhumF
rW2BI9NMkDHE3d5R+ESlRVGSuLZvSKteZBbV2FOjjPyVlQZJgAdAhuwUbWGlAVw76CE7fkdbsZWR
te3Z09hHVhRFtN6rusW+9GDOVj1P451mAL1R+5xzgBn9Azpqcos6/snyqyDabcDDUQhxTt11+RTe
fVkK4G1Ih/f3njUjROmwggsvH9FZnZqwtrE0scxppi9FjFa4HZP67k9jpCrXh8h3duy87/HnO0xD
oECLVEZPfkp5U+6zVYWlvA4WlfoCLQPY8+1ZN5rtRGK5VkKiKLLaJVfJtH6UefmycI+I+hdqKU8W
pA25K0s/u4QtKSiwE4pokGb5jHNUf/KZmOBTT6x0G5HZBEMwEzLcr4pYjerIdZDB6tsOrdONb5hJ
kStwEf223Ns4Z0lZeMToWGv0F0+yBJJO1LQ1uqT5S+xy3qSangXCNQgdWVFHwruCwLGvCYlbNDuf
AF8nblHw0kPwtSOs3/mwiUhNmgjjY1VIJxEo5TmReJrXINwA3Kh8Yv42FqZ95oSPyHcseSWrHGWR
Fu3fQPXtUVqAknGOQ6QDGylKplu+VVdNP7yiNa/pgL5+wUVnTsWfYAlKnxao8i0dVIlRtIPcA2Ne
JcTx5EExsc+DlQ3YeVG0T9TT4N7E0OWfKp9x06V44hfokJbNGcUHoqRx5+wr547gpl3sXd1MRxjG
BH83xb8mgJkeK3ZjCpgJfOMMpL2mMdN8Tjo9kMqTLV2IQbvce4fLgyWacz8IHrRnd2OUai5CY8Gn
MC7eRv2pwBLHnjmu/8lhGaMdeuB2XmZxkhzjSLbkLY8Bji2J/1qbl4bJUjubi3QIB1rW3X4sm+ii
PgoP9OZQkGZ+pej7hgbjlxhW6hse18q8f6qAlvjAIdVbsV75tK9yGIc7bIRywRUQYJ3eBXglElwU
vpnXHFaLbo97W2NY5aN2+64Sm57anLsBqhYwlrGZBNtFqWsVmQXLf7bkYtbPumJpbq36T0jdUDFw
IIY64Sz+Ji6eR7zYLNhjuv/RhHxv7RPQ2haXEkvMtJbE89mAvKLFsiyKElI/nCn1gzKUyW5RYa4T
xE8OHpAV8R8m6c2aX03pih66dinkL56tSF+707+0cBoaPP0ben6dEU8y8lC/5/DKivoF3ooOrtsJ
VB+XhER6FGCttMzC7XZCREP+YVtsehqG7jfrI7ZVNeeJPF48qBiaGQ21DfexibACWcaMzRGHrBJb
G3pcHl/xhYplXLBu1vl6Hnrp9H0QwP9WaF+7R5h/31K4iiibw1jcy5r4waSb/H0xsguJO8UEuk9b
MoarhtT+zkCfPoyBETK3YhTUW5/X5HBua+34LBSUECQnx5yJfTEqFoXqj2NS75lPQwVfhrpXwN74
zqDJF0RsrUXbwi7GSk12lJ7+1GphzOFfMUc7MCJt1ceKt0tXRLlXmp2iIUN+jVFU6KsCcTgZvgRR
mzZH8nwI/rvGGG/LGbOOCAxZghmk3egDUIEDKd/bHVj6ZoHPlaf4JAr18eJ07N5K5GVdkPUS6C3O
4cX5kDJgdTRDyWBKT8zNwTccOxn1NfggjTBiBwlHRd4C2FE9hW1sBWCywRC64rWDRKG4MT/eS4CE
qh39QDD6o6rotHp7JJYtUJMX17URHRtB4EyMeOE5Jbn9xbpp5xbViI84U1IAynaA67BALxFyAuSU
wEWQNDTWa0MokSsJf8N7F8jllVWxFhi6iptQEedszpQhpXvRxoWFUxMzuryo91dQi0w9B81VcNcq
R0IMJK/VYDsv9K8M+AZxtgYOai2Wbgie+zQUcxHOHtMmZXVcp8e2wpK2+zvgW5kC91siQEi5QtCf
ldWaKa3DDt9OV/qVto1v4FrUV58g/7AISRP80LoRxz+tNop8DlM3UuS2hdvzCZt0sut+SFsrHVTg
Z5njTyNCcePOR+S0D/IxJ4yk3PDlE3YFF283MJxOktdOl6MS/UTKFJDp1ZwOLvAbPE99rdxrjEWg
koIGRm6+15FpawQttdluzfNkLP/TQ4Tn6mx41ILln1RKqFy4Xj2kuSRIfQBLqLW7hZolq3+XGZY1
lw72DJ2W8NtoEgpvsUhVfdwaAYV/SXBQxl+Awg+fwDQ8PIkmLA1J3dqv2WW1P9oEEB+7znwmDSbd
fwAR0u0gDIsjhkevxkUg968JMpxWkNXo6Nbi+8JmPsGMIwiMoipmRtKxn1wLv1cROwv4QNkFxNCD
nMdNIqO3fyuH8sbF1n2d3E2F+smjBMQtakIJJBgOKpM3ctbR6fRY3y5mpUDen9wYFSGPNDzw+svX
UINRdQTiHEkwaKzpcj++bGkWdPQ1jn2fFEA85qkarctod3W4h8r0Y+NbVcj0/Q6Fu9P1raXqwpn5
n64wpcqpun5ka+wYrRvL7xpb0TgalXmAvU9L00SvfZuGR9EpP9YP00VSQRgnPnCEavSyNeVWvaoo
a+tC2neNH1n+AFHhApS4jH1ovOGY85lqO5O278SkzTTXKrcsH7n/bj5i3oAUL/lDuWfipolu3/Op
xU3b80VT8Zv8+pJPLMFja9oD0+0YdJDXapLM/wcslq7mvsqlKd29HjrTU/q6PgHovMl03ZVK4S+c
0fFKahqdXT/NnAy5X5molLNWdgvshnqFKihWrdmcaEOZ1WiEQs0M4B6q7bSpXwj1Ir+TXNM4Hflw
6VGgCYUF/jFsaZyWctGnygp27Lcje54pnpurcPko7cYNcAJlYkb2smO7pZ5xEGrHMjCvntluPDr1
Bpc8CbkZuoZTdpaHhaONDTeqDAEk2OQ6jN1gfW4DAKJSBC/ilQjDTiRxCRCOJiGkw/ACzqe9bd3G
/cpRt1stLq07pQgCtRR4B5l/IlSDYv+6lHVVgAG50bjZj8+b35SXlWAtsVdyRy8N5vnJ74ZVif0P
0dw4Jbv/4PbfC6hiB1WN5KRJzYFaOZZcHAUSCO0ihi3RZft/T+CZaTTUE7zC6wmiWdEdFoU9aotb
1d1vDV51BVQ019IzA7nlGMbZ8TwzqZ9r6ey9L5jpzm282cLrl8OXdDYuGzkVJFwIq8EvgR2zk75+
OmY7yxc6Wq9ZG88ogt9C3XQqyMx7hR7tvY8NHlj4VU3HJ+GLXyo+o5ss0kay60alQQAShZuv6twR
6f1C7A/kvYrzxbz9WhVP7GRCVmx4DYafZhFGuFVFUMk3upU5WQ2sveb9QteTaJqTRYMnoR2KpIUC
YbzWHBak8fn2TvJB71PmhBAyc/T9Y1ijVkhUzSgyZ5eSgfgSIKA1qgCb7+B2Y3VntSrP7AApi3S5
TL7RWKaNu5REkhAx2qB3P9EkBakMKDHavCWDbsPjXso7ERqvoN7R+pvhexXXozT0Ff5zXe6pnZ+k
gF9IYESMSkxU5B4Or4NNgFVDOjar2+VjXH7insQUoBP5xRi17UoTo6ROjqn09riIENx+alhi6f08
YGVgPfBZNQ/Ije795g2gEKadKDz41T4pF66eOJrBsGRDTzWlarZ2MyZBxXZgUiBA5mjqM0FxXHxJ
3JjLpUeTZ3ZFM99k/1XxegTESdLEcybKtSNiZuJOmf3ltSHyLuDCAglu7TQhOQZxTTZZLAOW9xxq
clBtznv1MutbUcaMFlA+rBYeSsUczH47Sr4JcoKiAu7PkD7dbTz9XyMcMxi90h7cad5da5rNhGcz
U+HN4D6A7qHZ8T0FkNNP1Ynd6mMgoOWMDrQLlS+H6KX7/LNUD0C8c3+j9CytUoO3mv5/j4O5WE/g
4kIkxu4+VmSl27DIapxd7Kc7oS/HHFcnWl4xO3tQy244PC1N0q3X4g0eW/LSbVfb8BY0k4Zs38CC
aYdLC178wGPMyFBQLuHRaydT4/cDgH8bnGcpvwQbhVgLEjQDo3ZpwKi8o9WTr+c/XsVC7d/EE4bh
FiI+fGE5VAwT16LDfHFHsVVJJEGqJfhs/6o6ICuWUFWbTWe0U93Ybcx7MMHt2cC7eAs98JQoZJZ4
PJPiVsLSha3ALP0oBGlweMgB44YbaJfLZmL/Orxtlj1C/ZNJd0CyDue/satqgUWhMU3t4BqpOZHX
rBXQ9KfvJ2Xop6u5/8BX+VI8yp0l2Kuxhwxzcy0TLvF/KDrdRUeskQjs8Reh3KwnFyQqvvh9036/
FitR2g0xSwavJUA1Hym3HyKTSOyeaCDoiMc03KTbYpMX9Be4CRGA/khO2uGQCIFFZn5pLAyJt1Yl
WA+3ZFjgtAx/K9Y0z9v1EnpHrhb/iIy9m9KISblECxTQUgS8u8mhOKZMKNwX/FOfyrT/ys+Rodqt
Cnw6Cy9aD9YjhWief3B7b/7aFqYIYmwztgxsZW4KsZgO31UIVbmbS/CyZgvZWUwKW7K1yFAkjDSd
9pCbqvYVm/1INu7hqyEnsjdE65wNey+V+7N2sSbHyngI7312TRzA1XgYs4YZmsdweDpg0tf43sT9
QHiMyA84jKQaMyyDsnq39SZu9CBMudA8HaG0S6VrF9SJJcjlnafcgvb8wFhrynuu9TrmiBCfAalv
GxoLGqOEqmqotru9Rw4zDuxqor+FZP+YVWVg3/XXI5CGrIfoGWDsfRnk5detYcdwMZehqj4Ifu36
FBIu/BTE92AD/nNv+fnkUVFwPuxo3lz4cDZr5R1il/Leds5thtXo7yhYOKgg/9TtYeyvaQ7HeSv9
VbJhwvrKy2TSSPL7TLuu2YhXuZGatSDdNlU0kvPqPR2HYQ6JF/GEMMwjCzNgm8SWlOyDmC0ICLQv
zO9ltzgO8I76ojqSh4lcRZlRMBAOeNTebeWaPtUs8HK/IEelHX8CTob7FTNldn0X5b7qo5bWifBh
Zn3oxkgyQiNdM5B6Jlf7qmjbWRS9o3Elg13XzqvW5Ppq8bRTBfM5tsq6QOmcrRDfsN+2OtwWH5/l
xLe2B20w2DaqYI3KtBnFyodQVfsNvcpNUhVnxrEbotGYkd2fdcqNUG0igBYjLhtoD9KrhbytzwNF
QDEsmLAx4bRG4oGmD1pa0mqAV3luAuF2oJ73W20c5DQ2xBJg4ihDtqGNsKKeHSxVgI7AJU7OoWkE
41hu2O57qhBgbxEYjjBT9v7HLZHX7IAVfJB+KEJthJehfVWLEjwHDERx8AIMunTL85uOi+QJNvbU
5/c2LzD9Ovy58X6ohDcjp3jKjIIyvXL0UY/HUEo0/zMfnB39mjpeK8KCHnvc467GfzvL4iVS9/zc
/l+zX2uio8427oBD1bAd71V4juXau2/r1faNnphEwi1boetrPd3Ft6dPDgdXTMZVZv3Ymo6YOrIk
NqTT/2FCdw3zGtpCxEZGMsCmTOIWsORSLAfbAqd/4/ajVdwBE5v0bpCcjmUE9mKB3fnplyJWQO53
exakGQoFOnI0OCAq+7aWW+jsSREC6gd94E0vXbw4WJjHBudGXUGr09A3qMzWpX1fZoFFNBsNp0Cq
AbLSK32w1WNbSE/LWMB9VpiG25ucHXvRcidAk4bVqwJ6S0D416FWaP4jYKWE41bys8Uo2wD0eQuB
j//4X956J5xZzS4nkwDcLshCWaMb5cLO2N+rxzSV29cGO/ZlYSdk6JhqxfUW57+TM/QBOqsUChPW
pgOmwd9zn6DcmyuFC87XIPTho7K3RvXTnNX9pVO6/eyAntMiCJb8RJ4u3k0V+0VqUp975qqvrdS/
zKPM5Kd3noqoBG9jxoFYrfELWR0igY8S34TIX7vP6/K1QH902CAYaYEM0Y6XrNqHDhlCKPyscCGk
8MDR2d4tDVGjnm5a2bRte0gYPq0/c+6A3hfOadhAR/WKlWhVBvqJmhrj1/ENDQagDn3Nc5trYrBY
VFfnpr6EU2GtggEb8TCgSAid6biEqqyozr/sGoqSa8WAjxpaAC1qRRiI3a7hAEu3MfxxCYlgcAdt
T4KeBPVlzDe6NbCftrdyu2yDUsj1mzzmjSOb8UsGzgDGyO+dvbsQJbdzA9S7bC52IKtjplPH6aHr
KMScT/PJ55HuJdmDVjTkjGU/gS3eNb0WgFxJr3sxmhx1PmGWpA19foRsBPTfIfl/56H2rgbSQPYN
lIc9b0Gs5oJIJT4ZSxtcb6+suFpo/pRO3oIe0p8BuuPoNez7Swa9QTLnbUTJozBl1wU/nRvG475X
Vh8IY3YUGuBzt/4sFnuQNm7St8cjMiAHdZYvrqdDd89BBPl1jdiTz0tCzhBuKVaoe057sEAiMzRX
6aFeVuxmEyLL0Oiu3UvsXIg/K8coy1z7S0EcpAi7EY8S6ROQPOR/qBh30EZveX95LHXS9HBoqurC
ySL2AvYgjZgHpV5y9su5lLlb/L0cvcmuabHJV0zc/YsNfjJGdvh1mkUp/FTFjLieAjaFnEaYUHac
ztFijfsjMLaoueJae1Dcw9yR+VgOZ7+vWDOUeUbhVml9j8KagqpCkOJ7xfIzb6G/VkUSZA6CZFnP
tpM+hIXIzAqQ38OZADDVEfF6vrJb+C0iKn2AxCi54P6op2S1IS8RW22O4bCIVTPkp0mYEV9Rv66g
grc/quxUNr0Y2wIHylU2I8eqB0dNHEtqJxrNo7G8GAV+5VCIz6rfv6wJ+rMz0Y/VdTlpTjtMnP+L
m5oRdZvB6WvDI47YH+vsNZiXDAwjVxzDRS44ux9ZM1qKDztis6ym93S+e9jEEsCp5U5BQY8t+gfQ
L+MntktVPbyKhFyQ0sky3PsHopQuPD81prKqRkxMVnDzaZflSK9znWu+ELyLtw5Z3E9YJz2lstws
usTgK/TkLMMlQRUlpopLRhDiLMZrET30/OwMOy36QFLjKfAu64SvEwe8govAjUnOIDduuZWg6hk1
T1pNDk13GubwcodbCzySTf49HQiwXIm+gskwiFZLMKA/VaZjGkvOrR5cAaJNDGN05shFmzWVP/JW
wdForEykKFlxEYx6Ud1O+GVN8vBs2F2tSC3PChfKDORZtO9mvvMfRLN2smr8uhg6ZSpJ+SLaUqmh
YYG1oDTUK+bYLGrPuNNKaFRGudTrsk8CDbepMuVZI2xUCkn2uBIirH1/0oy/myeBHitwTYK6DNXD
IxQyBbF0141m87+ePp8YKa1Le1drYNE5nnMBMp2R4Ocr4uxBwbgjr1mtDSB5zT7GSkpZZKsUYC+4
recQdCD6Y/a2/eIaV14SGeSVaLmbWjBovLPjZfA+qOPVzs1Qegz6emxUcC4gPeVQ+LIwewUcunTG
5lRjHQGZ1yb9YgjCBhDqTVEkAVQVO1Re93Nx3VaPAGMavsO0GfDm3llV4BeUEVYxIGRtgiI1K9bN
WE0QxB20ihn9hay0oyxTekilgCbOO7lLpLbCzch7buv+GrJ293UXU/owVz19VZX+8aKgoirEAnhH
nfpAKrSYQbIy3F6xS00OqCYZXYC3oBcXmUP6TbLjd4WEDbL5AaS9PrI+ZAjmvbucBopMXTEobFrm
EI/xsjG4C8AwaP3cu0MR/Qfjzyho9LxqvQRpswA4KzcRCrmY0EM4pQYFODmc2JuJ/OF8D4Ks1vzZ
YWARbX3XtUUGdM4Y7SiAHNR4Umc1oOPlN1R+ADuoHTFvLfqSGKfy04FkduIts7bVDVQksAJDMxUu
f68Pjs/8UkBaD6k+vMWW/DfvjQDAF8CAhjrGBIXcxd8tLHWiEszPU6hQ2PUzkN6JSCYIAimexfqq
mHF3mZJCAIQwdL876b8ydASAiOzKU49UOjL+57Luml4Yyl4DwLR2/VZ4dRgBVU1R8kndvCU4WCuk
GLKcD4eo8sU4TQTcVbigE26B1g5OhoF3AHclQhaa6HlOCKBZziv0GtpZvC8zKV9aohie/gBZ4h53
/gnJgdzJwJbwe8dT4DjuWJq9/1FfXGYU6oA7er81xSRGEyI/lDgmRCjar5s+E6Tdlo2+F8C48DCT
ac3iMF4lMp+LXMgEHFdRuNTw/dJ6Va+WFnN/sd+dT3IAnRjJmE3YyHmE9mpB9gJeiB7yhjh40UXP
7MnyDRz/mipwl2EmN4S6EXhEMAcfy+Qq1W2VrnYYD1FqrefFnPGF2XrD11GJExZarXN10+zb280f
8gkRGJTZDs44K64EGAZevOX2NCnYUO5WIEGMaV+nHrPdWdLIuOKn1+IH2gAGe2xGRYdWegiVeXCn
+y6kozocXo/i8FwEO9r7yLlPJMSMFHnkwkPSpS7W2vvpfMyEPq2tMuohSbu+uo6DFLx6GSN6O58R
53llM0Kh7JPRHKHxUAEugWSUA1EZqFMILHjMkjbiVU0kYgRh+VapFW+VPTwXw2qSwrJbWY520f+X
oUNdmI0K1gGu+eKZKBf4Inehkx9k9BM23SYvDaWxOlRw5PCUSSUSoftaznoaGXAfmoGw7cHXoFtA
PICMKZe8EUdcurtKFt8F3LL47bVCA8n51Xm2EsNDf/q9kF7HClQLYj9WZWk72/UoK7Qwhj41OpWS
WtwP3RqymznhCAIyNPSTMaqS/YYbH5+84uXt7WHEgueTYJ1lslHCdxfn+gc14ab2D+say9bsPiEX
yz7Te5VO3ylobRoGcsbzCjo3P3DGJnzW7c6hbVdHvQhWwTmCYrd/l7WCc7Ne5JNj0IF/JN/0UaTF
0KZjKYGu5pwCtT4abCeI8F+LTWAp3TOdqFy8BIxGG5G3ptYmwltbqaudvTgiNGl7NmY3XJK1HH3v
vmpHzLnIDEbVtRmnPZDmVcGhNqarxi7Itj8QmSWD38FfRE+uFonu9hbtByyNuu0bQTE2IlSg4Efv
M88H3yPw+VPy5SIiBrs2WROCZZCVr6WauRgtbOwMfysL8qUhqf8VkRCgbwAshvkzB3NFrnfEDOyY
CEqnVm0nxb9sUrGDRpsrykSmfMnocnYZxUCAng4dX2Zy8wArkt3ZNBONy3hZVQ3UEJ0kPCjpk4K6
gu7leTBmEZotrD1iIlHAKV28xvsU1B4SMDiELn1eH+++IcTvcjUVY8lkoXfUM+l3YRqv9uIU+sbJ
7DyPf0Q7zS/CWgxe/Vv6zCALbvFhB49uW24slHc72Wfp/lSvlWWH2S9rZ+dgkkuHYj5LifrYXXkN
+NK4/tI/DkPQzRgX1Bok5UAcSODR3xNwsUOegGi7LmWK1AlvmOoXaAV5etDJb5eK4UiylxxW6+Xq
xY3c/522JvjoCmpAVGKealjrV3NEr6DwkAPkUNP3+hyBIStPnzfEdxne39Oq1VB6oss+twatqJ40
daD6T+7faheTvcsOloHr5bW3fY7PT6265H3j0eMKMi5Oe/Kbb6qzdnoC6O8OpNQ5hjRfEcWLkEDv
uWOcBzSIpWsJ8RcZSkq6aLNsfVu83vpmFPJEScqMNMbb1UYXsdfAg3/4CEprk1lIXvrYn4m9AoQ1
xjAeXNVaPvyRDjkZJ155rIis4ES+eElfGw==
`protect end_protected

